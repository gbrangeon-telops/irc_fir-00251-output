

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OHeaBmhw2WWXga/8pOVTMIzcYutI6Mhna2kzvZmeKvttg8GRcsMBDXpogvkdmdxp1KLLzWXMAKSV
fUAOBPVAvg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ao3tKAmGrk9jDIJ5tmEl5p3MIRphIc7Vg/SqO4TER/rFDRMS3J83CwQ2b9YFrnde65FSvizCvsTV
0Knxkw8zoIma+TSgIxOnivhI3WBhgKeA2uGkUI4h7aI3JKyXt+ar8rATgfMIjtkwwZmXnAQdFAm/
DhnKD9KmESp1ihQZWxM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tIRCJBwrqw861TllYkYZisN+3Hf+P2JXRGH4rS3/mIyKaeRa8ciKvXh+DuDwE0CQ8FK1JKt0o7Wy
5niCab0pNdgMIWoeJTN4M3Yv3mIYHhxe/uhUY+qL9dbTdi1peu0ypGwB+pCVAaCMnYsMP87ovoxG
mFxz/aWHoq6z5hUiOqs/8QctFGTu5uGrqo/fDpwnQByfUDzc5kOGUXom+7Ix+u0CBnUzxUPMVE8H
FW15FWlEhZ2/WOv5odw8POvTaQir1St/I4TCBaM8Ne779Z1F4E4v1nyrImWHcYGt30Ex/kdASWup
x0rIb4g/F4zfpMwk2F9PI0IRzfsxsXBx1PSZmQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vDR9iZfmcKoc03DxzsUkjAUcoXZpLGp+jz9oB+bhIzk9fA1B+YkBJ4B6wGhxOSVsIGzj0A/2+sve
cYv4/y/PnMWoVJu5GAXMXsNWS0+yhRlFm65eqZTnif9T4BQLUfDB3Poe8t8+8qJraoiNha1dShh9
FtnafnjfaWlgFCK4DSo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P5OVsGiC3k02pbA8zjICborh5BXFBySD3cMhIIsNr8DZdx+UrjbiVbqZMU9Ry3hJ/1iX0Q8zDyFo
F6W3nmvV82n8xeQJN36fxUpz69izOLDYVC7B/XqC5I6fwrewIKThxTuK9lZtFdQHHrzj3T2ZDLDy
Z1+PK2wQ4cNjjft1DSS07aO+6gcWXb8X25cWmNGk/P6Hl0pzIcfFFHwO6Oq+bJ671kKmsX3jUKAg
DTTCgxx1Ex2XG0j8cWCnhZjmetyd9o4fKBdb10goxmIXB8/8Sn+4BcUJVLUQkMnRwy0YJGGtpiHs
ZxxUU5IU2sy5csUBb6rGbP4ap8jLGVFhtMQgiA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16944)
`protect data_block
5Ut8NcwLbNigFVJABwwpFfb9GH5WLaU9rx63KeF/GdSK01J+1lY+wXoyQhTzRCsU7Hf/J40uM/ha
2D5e7rKbbo6Wmu1SeR3tJNzmTtGy6/1o195cWniKDEsQGf2+t3Ibp6rw9/TKewwp3mJya/k6Ynw5
1ADav3CMQa9opfaufH6mFBoK3HB1flV6u41xsIfDlWISgFQ8tahRqUQkrZcOPL+PJ4BIUCX7ExEb
ZfdmTyetxlVH8ZSisl3VTgfoIz0wuk67oEu0FYJoVcflhVqMqBjJ61H1r9mtWjhFx24/kg/jV+4o
Y628LfqjFvQ1GaeuO2LXAIyc0lgF/EDg7IF9olchdpebQrGvWK+AtsbS3jKPt5IV8nSyrW2DUSFF
7ZDN/odWLoqfQXZCYgjA0tFsz5aU1JzHx5w2wy3WWBxDXCCQ9brERbukV+Gf3oHjp+SAo88TUMxW
8kC/5KBlUr/SIksm56cgBbdwM0cAfYxi/zuxZ3FRzYQDBQ1/fQXCVH8pwIwWAihgla25IvTnK304
FPMNa6OVmcqcmxSCdrxZGJbb4yX8RBZ6gl4hr0h5J+HZMsq7M20rHE/A9ZzDUHZ+nozMlRzBVPMw
XKUU8FHtDsyfTh8GUNe2nONBHButy20x/8PBKn72ofYPxIUNQKtoUNnP7GhXdsD8lHFSU/7P/Q9j
E69/Sg20g//Pcziz61qOw2vhje1XgUyh341CxPhCs16rEiCQz0iScyXYUSGJ8t3IuW62JJAuvaxI
4AY0J2XU8o1tJk98wVesBhmynl49AbKh7xMjBcX4aNH1jIMjOWG9r+v6UNGuVoen2MyhcOi5osGf
12NwAg+7LE8XoDvYsB7Dvix57aL9f//J1zNLZxxklPK3yIIhI+7opgebohHzB0l8n2zADi5c5M2g
ADkJtE+cGCO46cc3I5ochDQt34PosgBSAmdD1TPrdag3FqY31d+dnOvlxJ8+hL6JKyMw7KSv4A2X
z5S/eoNzMGdi2hADWlEKTk8/m15Els7esrhXeuD/nup+4aq+JfDFF0beoqTQINqqfC9Oa4YibyBQ
ayQMJjIa5dvLucgoe/haU4wrcUKTH94Q/pjbxhiDzJSP8UwQCZC9njJSIO1y0j0F0+OY7mHM21+2
gRKjb193SCDpP+axw01r3x1M1qpC2wNBy/npoNdDlRHT6yq+/zW7rgSpWxTLJA73TTLLNuSWKcg0
GJdq8/POVirEaONSS1bqfeJO8G3A38uonfUj93DgawKELM8yNnkN8l97DlEeJ46BaPTMvTClkkGC
0+Ut47tEHGSmhRn3kiIDuhRwWE5qHYpRxrzr2T/nLup0g14oc0QlouE5nLmv1zOdfv7/NBIXSuzf
ZMbVkgzeBf3ubDpQspVyeXunbgCTFRNY3u+yoDovS4BF9WrkNoZEQNvTk/qYsFY0B8B9EG+7d3Ru
wV8Kfx1BJYUq9XhtjheMdloRh1nAaThZy93VR6Ta0L8RGDbLmuO+pmXWkucCpgdC0C2+ZleMyqPQ
oZE785W3dybx7m5u9BbCnjRO/zWiNT2g2k65slE/fRaUcDef13dt+yeLVU1svrwkluYHBc5eIsrv
671+PmDgJd2MAfU3ct+BSdO+/RsjrwkI0V0occ6tV0YFQY8ZtQZT3JPGwAL0u6ZAP2z3CP+LWqlK
H/0aOLND5nWEtaSsQY8YC37uIcbMxIYNkWNIQvLSXgFuR+tI16EZJqwYBQsHpPUGBCkrf1nWTI+m
0AWkwtqsIWcEVnblOeH6f5WVnekCrehBvsd3MViMhDP0scXUbY4kq/klTf+dL9JLsLMwXRhD8dlk
r7SC2AUBicFJaaAOOK9iPfzRbk2zq5IlD54EGSxnDwH3uKQB5eyV4GvjZmxzAlPz3KHD71834SJt
YZO6QbsQB2eJnMhVqoekDgxzKBICofXxxIRpt54j/Z7/4YVXZuaXLI0W5VGBj6oD+7qc/AW6JIS9
2dUiorsrPfljjVAFpaPKPTAKPZOKUGnSbAyrxjWUgG6Mh/PtIrxfqqHiSA8KOA3gnoDB2jUGvUOf
XuFMTq2UqZvCnCS4bpuNmO3kunVSVXDIhUrDaYzMZ6Lw7E93/tbPlEbouk8lW39u3icXnKMmSYHR
KvgglIeGfq+1DDMZYcYbZDcwmS4KPdpZzuCctc2WkL4zY9h9kfro45yAWdVp8fSh2hwyg7xUaw4t
ZB+EzA9TPTNXG9kx1IgZH57Zwp05F+oAfKLQufayzzTU8j98HGnuTMdi09t5EEMDbBNILabtyuIJ
c7dF9seSdo+2C38Ss0gM3HJ5dJLa45DevAiUouGvBzDuHrvPnfq6uiH9+fBOGSST7nKzk1jROgnt
LtCc8MS21QJW4c7rc7LDMUCEzc66Xju1c+hUcEFtwwbbVOeisnmuAUEv+bFF9OOwYhphWRRj22VK
L7FCzuo/ZbaHHoU4VWNEu001mKdCDmndanypIZNXF7qsVZEX+aoUQBaAAySHYbGXZ6N+xTkePr7I
KTp720anaFmfvqIAehjShVIdGyPAoOXKxv/96Y96EL7oqy0JXXdwJoxD+J/n/GlPpNAoJygvtWoi
7gKeaNTodRRrNaCypVipruaV30FSP+HpKuMs1Xi2Rxg+fduh6OzdPQic5WNwxUKGa/A1v5JX6/G9
F0PjIRTOuJnIVqHhVJwiQlcy3cI18df7eK9YZnpSm3o1dSwyBTXFlMA5YmUHeWa6mIeu78q3g+3b
oLKd72wb1Hul6DRfWHrgiwr0IylEfvrIw3X0uLkSRf/7rEr2++twyj3jZZQufJ1NGTHDidPm2e1y
0e2k241JRnexhB0Hik3IWnfdVVYHr5YG3zj8LmrfIzuruWLGezdZ64UufZ2MuatClMHUlJLEhO3j
YqTGGjb54OT4ta3BM1NlxxAUhVYUX9E8dRZIIg3wrf5HscVfOp9ynJlzZyLo5ay+8UQIr7ZGWKdx
i9uE1kMLndh4QXjbL0CTrC8jbV7CXLAzkqFeZDUKNwvjvRSgJwlHzz5VkdIZ8vZSD+iAEXK2zD1U
lUReY5swhjVH0g2t+mFLQ8xOGFxQO7zksec9X3Cq6RiMH1mr9rlSiCJazq82KnwdmpDqJW5L1hJu
0Njzd/ykPCgpcyirqu93UcaOhh4+l4e6kJ7oo492TnWnVOfMvfRD+vNlJ0p0BIcZ8C7Vmvnr3fBR
5OBhrgM23WH4GH5yvSL/6QLH7NBD872fK3qA0/6VXj9P1t8PBZ6awFN0/w1XXkLFuwqqHfzVr0NM
J6NY+joZSyeFGF7+HSYQ1X7DkS3ftALWtWYwHBQId6stEG9ujxGNINoKSeMtDZ59cYun3tHyqkvK
Kt4dPOrJ11LyFiGAHUnqZ0lA2/s/oCq5eHqWYe+3U38vjdMI4J7LOfClyzZAqJTHxY2ycoZCkhkr
pLxMjlFrHCKahwl/sPKv+i+48w5flZjOui7RX9j2S40eYaF+ECmdXr9GF/fZo1pembITgL9lDSaC
o5W99B/6YZA5exj8JcEV7P9iefYC/Dg1KXlQWK1mLfSVPVmklmLfCMFNI2QDcVBkZB7Wd2YQasix
V9+May2tFSKkhNOmPQwpZH0qp0p9YnxWv0077MVaiGFMBOGNtpEQdMGJcwUt0JA9evL9KUSfBXJH
iTEXuCwaeADF7DZqQTn68ltCnY2Gf171Y61OQscfY+x8zzQr6nBN0KO8Q0vCvnnRKUcNtVBqtDqh
b9RNyNp/KhW9pf3eww5+lnpudbGwIpOqoRUPd5SjWAy6B56tWtEMGi2fLJ+6W5SKngl4AQHIzLhy
Uq+GkUxLoXzbzDdILYt0UOa5aZPg5R2C1VvwupnXReQ6w2lWNRQs3cTJWQebnmUJuM8WjIv5Igv4
j2XCbeOWk4KswzC0YribfQ4WwR7FFlzZEOwH37GHT5z2Qpo2XCbl44J93Fdv4i8lCeBQvmnJZVXc
ozOwLW1Uk0kHl2adnEK+F6mwbOs3iVfkZnuwNJ/AAIWo4RngW5UuuMPd3mJpkEoiVpvMM3bVx/Jw
etfuYWEblKLG7jDgwkO3JCEzpxGIND6MuZIt0zFdzjIGTTOf9LkWalDgGdBsktxn7NBoTbFBqPXb
//oT2DQQQU6ZVXSI37Y0XvPaZtjqolQVxuDuKWJHeSqHps0/1me7cnlkioVOZb6CkORalGcAaUUk
Bq9VZ2I/hAPaPWBz1CYhKOJURkcXU1XNdtSgQjjbiraUcf0oh2NZRR/cPzHw9MVTonYLDdCo0BfF
k53AzGoSk2OpWjw/Irrp2vP6Q9jatvmAF4/pGT0culnCWKaOvmDaD+EBr7HBdzuf6bS9SEaiEAiU
p2KVZpKNi0+Upi9VK0+wb5BS7P9sVdgzlttyAaF7x+qk7vosr2vfNC4nAZDjtctkV8KYwMDeXRqJ
pHkh1m3OkIOP7nQfPYQQaANLUC0dPXC5UqcozJbGxx0/wc09aw+4CyiRCe1it3i/V7PlI4lHjsAV
bsZjCElcWe7Ix9xDo6WYC8MxxIuXRH02Xg1g6Rn4d/FCimSL/2id23qW8gz6rTro5q0gBnRTYIcD
DH8utQ5XnB5TsKXkZKXgdwIl8MytVBF439otxtMtfVsbZ+Ws6EqJTwhyLp850QLvfzEjIubU3AeU
dWukfX10ZOYZr4w0eRAenJ+t6fDHJcgHU69QOyl3ahsnxEFuJvHcJbXUhGw/HUVQtnhC1Vn4ZMfW
vCuIw9D8gP5L2wc+SRGJTjy7hv0vMUGhZNlwoKkAiHlnBT6/LrbhSWXsMNNvd/BnCkBWinEiNqOI
fRAnwLDxoMqwvjoR6/jYEV69pEH6E1Hm6zmO269dVTTBvACVPIZ2f35mMaAXWMTk3HYy7NMb8/eE
d+276xVif+ViMNAwO7Kg4E+pLaBHGPIrvaRa9nqiwWwtw5+R6++ybet9PjEiLp3iMwA7Pm/Zvw6c
tJX3J+yVqDvoq+BajtdFEtrvUzpWMOS0QPQTudDsGPaPS664s7U7sO6owexp0Wirq7KxFszrCgvW
1ZsTHuroj8mn16sePWHdS/2YPX8KJ0riGcUoshCf+t1Kjoff+SqUNccqI0O4RTXNrylYYVYv2S8k
giBdjS8XUUUfGXZt3+44Z+uGeKjIeQFAsdWS+a8YBR3OZ3VxYNFJBZuJuO565b/wb/Ujlg8PgWE+
pnt/c/PaeZb7Ffgd/VtovRlznSdYGk1LHKzOEF2t7nSY1I3Ajw0qYU4sXA3OlmqYWaPnfE56+9q/
doV0zB8GIAJGDTGri1jxvs0yMKzeHgBaU5qBgRHYtHTJD/9py9w5cBz+VFuSduJLZkpgMyvnmQuL
MJ74qBWEqWCxvfUAjkh2/YupXPfQZqdPc9aSwrVzWecDZPPujqmmfP6PDSdjVC+wZ4Zx9AEApXMh
ijrLnEEJMDBDxccvdD2KNVj1pe8R+OxVt8o+ffZHYErsBX1wO7uJkzDRxLeBu+SCRmYhLm+DjoSZ
YWoZNcEtUFi7HwEAW1W7o6r3z5zwi7DdgW/nkBaO3JL0aHHT2CpwppEZ6b7/6H/FM5HgdoF3+rZI
uXw9I7G22QSWiuq00bDm6SqQVxNAYJegdT0eFK2raCPqyMlXQRcWi/B6Yk8DiDInH7WyvZESQYQ6
JKhIoy4xu/igk7OqeAFxXBMakDOdPPXpW/pZ1nITnkQoqCTty5TW3BNhuBsiy25uNVs1H9tm0rCa
OfCcJxEWnQLLTmnvYy9V3Nz+yYH8oEo2wVZ9SBF6K/IuKzjO4bHWPXWaD0o9OswwNeVMe2NSTKHa
WZy5hER+lDeEL0siWTCuG4RBL8gzD1PwW8wrijoVyyr/QY7FfwC1vz5yTRdoBM5ZOdHizk75ymBe
C7ttTgJDTql9ZPcURBT4ogMuHyXkLqV6XfxFWKFltPUFDT8IvGSYhmrNVrniieKXcgmJifXyaK7I
DPSPIg9l4fOtOnH9HoN3SAn9EKLu39QUca5oap3MlBVJplLS3cfpDVgQilYsfJUp0lXuD1XK25y4
gsFiWRY/3Q7h1XjKoBFv+4W7wzhXLPa3+eY49tr08yjQIc7m0fkX8kfhBUI5RSCQNLummVThn6sX
NDoXpCmOxxhTGd49Ov6KQqzjlJjl9QctzWNQuhfR6ed7claVjkAt8QBvIw1TW4BvK1tBi0DnlSVm
/mSFrNpkzWByrO3H25t+KPcJHKVahhlWF0IQTPKwXW9enzPkBXSwA8efRRJNURqPqNvfE8in2Pym
OyVIF2r26tG73OIm4jcPYZ8aqmcETLVF4DTDqPrNK+YMipiH8lHNmo8RqtWvI42gTRJHR2+rHfO6
1OaKcIGWqr/xat67c8K1QUMM6i7qR5SSrjKtnyqULXauaPFCyw5XUoStEQ8Nu/fR7opwk8jmexcx
UNzTs50IRd4ejqfmZIotM/NBuefgdg1ylhSfcEpgi5TH8Lg7bWgRxpNBr8FrB8b7MH0tA6bWiANu
xM0H++w+4Bvld4XISfUgdcvbUvdgo3WYSLh34rm4bloyPaJpqcuv5g9+zuIIQ/kQAp2xVBQw0te2
9ZVz1dzJ4LtMZndrsqnfrxF1ti2Sayzad8J5Fr98u5/eDk2HNG3vqjN1FoYas9ftiC8MtVacb6km
DT7Ly9TVLXFk5dMeYM6viaT/mx61TbF8iEG7AGU/GsZ97sxd2SiXz1QltT2mWnKaR9fd+zOxunqu
JhJ78G7hAG6wJnvD5gn0823v4zbsNZVxyWYGMhQ23GhOXFr4P+ZmQ6Odd7Gg5FXFnWVhMGkBboTV
WHbePoNr+irJz//8mCkk2dMlapvQXvxwOmuhy6dS+7Ut+CRiY0ng7oGlFhKX2SleMZZDX5Un18aF
rcaLhd8RWEqwUP0Z2wUIUh6g30iRbNoW/eUJ8eIJguxKGCopB22WXNnrkP3PsOteaK3UB60hJWC4
vfNCFNc3vRC/7k787PY9hUXGHAyCQ6E366fqPwbUYL/2xdVXBOnOg7WhiXqhw+ndoKryYFxlEVN9
xyJD7wWnkB90vUI9Q6bLmwB27RdW3Mmvf5bc7P5obpECtHvE5Peay0MoV5e+pYPKF/uhx3GAGuty
VcyD+o7pkZpDyNXh8mU8Lm97h6GkjgcrAXNGyrEJW1VyIzNAcP5DNwEludSnIzApxEs0rF32LMRx
3ZeJ21GdfGsEhiympXycZrjrS6xeH95jbNkcVQ4LwyevfBtS6mTMRoUmORaBX1zxovDZpLTUwaqP
Hg9mYo454/HUgV1VLeB3yRn4FYDnTUPxIayswFmv3UMsgTJUwarjAcBZTCubWb8rGYoqv/fDyuua
LqzvMUveeOXwaRzzXqJm8sUju66ZDdNx2qBeklXSL+exhbDkuFxfaY81QRf7dbsDsrWp0fqLSz1e
haimqN8BlAD9JCdBeujW5txNDKYlYCexZRraWdIGQNJE1s6NlrxaNr2CY1V/QHbLNlyVUsOfiUGG
7KKbVq4kC7NX/QeAQVhbuypJ/QGUr2DKvPT8irQrN1Fakdc33nDw10CFgTvYKHUYZ65KA2DbpNdf
uTG0LScPJkyCCjQPygkqajdHHTC3yOP2twt5CHwXGMDzybme0hFlx4Q5ub++742A46t19mEpmA7+
26XSAiTa/aj8qf7d7k2wBoAaShKG3dACBm4eB0Zc3Z2/iFgxurysPiafIh2/cxvRqYTaxexwRXZD
IorvPYbhG2KaBP0QE8Uxz0qAFwfNAxE5+0z25Aqou1VDeB6A+GvQFc2YP4sDRcRTHh9r4YPuNBgH
AYrCkvDJ78HEgnM/9NwBBeXvf8hL/7u+EPwgR/e7trBHevfcp0gEtsbH1rNok7icP5+PRRdeMyHb
8n3Rw1UeIqFC6qrnloXSvjYa+5oFcyZCPbdpRlkvCaw3IouzhehnXxnbvyNrrs21HHeL4V20Xduq
sasJYHjJ93gcpyysYLM0YjxskxFXknrmOuuQRwiprvWaowW7RE8GwChJWXWIrieJg1ap6FH+Msoc
M2OSPtpP9Pyo/YwtJa8BEYqC9OfsrDy5B/1W8csjOhkmjmEk7tR2voyMULDcsxkcRjJi5903fhkc
p+Z7fLC8NzSrtIqZ7teKuBhJG+nl4XrdXFFfsNTQ2TLDqDzinPxVAc7MWrSluUJN6P2BDqxfNlAg
CiZkJbWBvhxQK11uP2X/+eXfQGu/wk9CmwMVMmF7q6i5IkLEgsNa93s7QLnoARdv3xw6nKRTl6V7
SIojjLij7u6o8wUSML+ksW+98Z0oDvxIzgWX1Q9Rht+G3k9O8QTy9j9wogDYog7y1XHvrB5c1R3P
bowFNEGCC38EelY8A/AfsowjRJxn7iDScXyZpBU0dFiUshsp70OfqAZoK6/kfusZhVIdQml7kdOR
gHIB/Qz7bfqSN3ncruaui3fLkYEcR8Kq4KDk8JFXiOEGefGug+sq1VaiPkj6QzzexB/UpP62Yz+q
JJSobTScJLIHABxwY8tObCQ4WQx304inIbfdJnRyvNV7wt5lIaOaHnlyjdBnq7JKJ4ZUFkra4mYv
kGS5v7DFDcGVItKbzgRRYZssTNcBfcrJ8JO95aCU2uphhYqeWSGGxXY3L7IAjrUjwhw7s14mO0L9
olBTaD3PO8bcz77I6654mzlsyhaqmEoAn7ocAC1fRpwIB/qy6NWhZIk2A9g/MS/cZy1+IiYYr+Tt
pv5vdAzpsilC+XW8Yut3xPukQLV0fG2+R5bglW7yjEidrSAOuJxpfS8zk/e+/uSHNXFaUf+cYfbO
vB+1RWmbZeceuR7400T++SSCGOVYx3efVsLOAdJVLA+GyJ/5YMTzFpyOOCNUT9st3feTQGIS8e1y
dwn8rEwg9yZo1vWEhntCbBCJD/uLxJotMq4f7AeYIeJ9ZkfES2O6uSRETZtH+Gk2uIo9uPJdKub3
kilp+vhSVTrMGRZ02mRWwl6tDUo3ZEyE+7YlImNeuZzjTs1OLfmbyJA1DxB7sqMoc3kkR1JFpjV6
GzLAcLASUHEsiePasvbe5xzDqlsmOq+14Qys1dQX3+nk5BANhQhsyGjkEqaIpqAfYuW0H5qrMkco
RScvu+mPqoKVUQ1y+osFnSyqFSBDu5CI98W6s5SfYfmmySdavoB4r/t5ZbPLO2a9nd1USmFmV721
0Fir4KwW/1E4FnZTJ04V8/Xizc9vp0GbSXfrRLcT3pyj3/nHE0Ql5TXwTeJjktQ3DfFcGn07brQX
nZ2tgVsFnnwOmxLGftgpdqjc9Jm2yZCU5HoiZuD0itSe5jrxQsaTd90quwoO22M7JIu9DphtMOtJ
a3eJGi/Rcr5fB1Z77rATCtkdzn7uo4+mdqLyH+YsyOGSWlU230vHgoFHRTs7NoOIjJzfA+7lOrK+
fsalHNtqNgQcFX1qsHVOYGqgJFAWrKtQrRUZ5BjarMyW6QyBLHNWE3FQ4N4tVoxlviYM0HNQkAlh
g6KPAQPzU25DfdcU/DvAT7cU8j9BIpZPuRt+gh+DJG5S6p9KrRFKAID7nLGg0rC1vX2Ea4q3zvn7
p8XtnJlJWnBb8kaLeb6KAzHIRKdsHVmY8pm+Em0I/mdBDl4LQ9QWEj7o7NANJmo9e4Rok6q7o9SH
pEFBBdoM96498x7oGJPajbLL1vi6LpRj+R28Zu9HrEhU7G6DYEYNaHthAGTSRmxNx3DYLbA0kYfn
3L+7XvqK2wSDKDrvyKD3910Ecb3rW7r3ZRQc+3rOsgdF/ppxXmyUzcKs3sftnp2khJnHHz9Zu4YJ
75PNVGo23hU0F9rrt5y/z0E+OMIlQ2/K9y260EZn3Qrr+OlE90Xm38mp6LkV56ZJmYZQMLr3jjw4
3kGWYfHB8dYXXiGT62Mb3URXbWfUnZ47rQruVBQ1FPl4evvo3i0RscJTNM29TgqfDJqwKO4rODNX
9k/ra7AXxzMz7djsvn4ZsRZjcAh9vV9eIpCvXFyTt6g4XuAYbf3HHGIzEJaKbwnieOUFYsXUOPEr
MbHWT6X1nuEKoXqnNJ5Y42wuRgKUh3UL0OaGqwQrdoH5aOlv4Rsg16w5vD5LdBN5xRjGSkr/ZjFy
zOEsibzclNwweLdRLr2phgswlLbUeWA/zbhxskgkunlOe7cMAfASuYBK0pQzC4VPT7iX1avX8/4M
1IG496MSf9bB0p/MfkuT4c4o+fUl7oGL2chfvnMZs1+tdIITzXIcMfsystzBOwtaUkzKl0o0wFDH
GM28zZZWccqev0VEVacaCcDhsLLEBU/nnneIxaGVWOvZGkyMPJZwwJ9JALccD/E2E3sh41bFLsDx
yHimFyk8EKvoF/lHtwxKKt9YujCIRKx58b58E8eNf4/euot9Nok9dyBALhMr6tdoBu0DSQ7nQ2Eg
EbrP+HMVXqOBXbXoBojSiIu/kiOf/QV05wHP/gEtnYlNa0eADsc6AGvddE0DtZLMx3o82fRYmBcX
IBKZA17a0oZyBAGTicLCyP/EyFIROA2OqbjbkMTf3usM4vis5gmj7Ae1RW/awp2JZnkg7Qh3JFQ5
ZxgP4ZDOhShV5DdQxPgjLCO5Mh2wt0rFaF8zqWB5RUWaQxNjXbPSUY2+cH9kzLoRVcvG30cTfF4R
HfUor4QTUwzhLEFIS4BSJwG6+JGj8WLbBwXJqRxjcQvZQ6wNQ1virwUoeFV+aCeSqE2nWbV+rhAY
YfGtWb+iS+8ABCjgKXRmCkc11CmqyfLYbGiQy42WucQ0TanNv+G/WBXRSMRXqlsjqDDdgQy+9trS
63fR0ML63t/rnir1q7TIQe28wsUF9PDU1xi+r4xCwvxXKSnCUcu8wTWldnA+uoaEbidrhOcRBJxm
NMM16qNkmas6t0lS3iri8DbgD3zipGgP6l7vnN1BNMQw5FervralTPARm0Tdq2HQA8iT2hhTLLCM
ndIzJj/2MFv872t7DpVyz/q/lxjJBDW8MM5Sdc7enitjK7p+cbs5yDUuueCcQe1QFuAMwue3V7uy
MHk9lttycErz8BYZQtr7anQ3LjBp8kngrf8GP3Fep6+K7pzlmuHFlfrXArBRreOEtuSHAXRrBSP+
P5mXFgFd7qEopelolc2Hn2HG7jBdaVgk50ykCRvVHjnAGO2WB2YMIonqOYt6gG+zfA8VNFRIQNKa
T38iV/Qm04gkE5gVAvqM08+OcJiEuXj60lpVC0zUTxx76rmjoMBUlgEuIptYBxNWEMd9RudJvk9f
d8u/PhkH31Vn9VnIMS0ePO3swWEDoIYPlHIC5D8k0ZWpwkrVKD2VGlmH2+LJZLAzcmCAvdfv13lf
fYkD1WeBOm0EXjpigMlaqjtjrUQXQgiyBI/36NbnxKsWkF1fVger2gdsvQLt6qvdld1bluGh4eGC
FvlGjn1EXvEeEFHUGDAqi82Y6RlpuaTy7tGESDEsJUJc5hjYAkzyJGh4tvc+UK+TjaTlkxMvOC3k
AHYcwxT0HAw6rBVcM8sSm/MrJ/opwNywGS7MrrdBQ3kcQG1vW6G6GfhJPzAtLTXDayMNkpSigahm
HZYXkv39TqJa5dBMNtU4gYrSbMFkG/th96+9IqSYqldUfkg9KQYxaun4mlLHIaezPGqJZUkSGGnd
OpdzEoa/lcS2v+d80uKs/CDMkoIgfIBfZriqO1CkldBL3jjpxeELdoVnrhBXd+PJPsoCr+rqLMGb
HzjPs0m9W/lKnPYEAG8/tJOKdtYaod85ffHm3mjbVUgINU+Lm5+zUomroic2EFjmN83GRXaMEb9a
2/dIn6+MeQHoEn7x32JiYFRkU76gcO1BOh8iFFfk+Pu9o3FODdFe+E5d7coiPTtxn/IqfIHQf9Xy
BdVKMU6qfq2Gn9uYnyFTPJw58zGTkZmcgYVJ6zJEZCPhePd30U0WrqOaQeFzfDsvBmkyVofRl3lg
HR77MTkMyP+6kNEYrVgEXZa/oHwM5ewcXn0NsyXNOcvxcJDOgAYm0RSlsItueZmjwIBD9Xo9r/yh
yrrdCBU1ZQ7+BPcrObvW0Gc+tNVlxU1lBKOos7FpTkIH3nfojF1YJmmSgdbFQkGo1sCWakxCGVuk
YIa4InY9PDuxafzWHX89zOG+j2elzMEIzjA8DOajF5MJ39aqyN5cGNnnT/1Y09xX/vDLLHfDrNh/
Ay2tq0efqu2wb6kru9PAkmDU4aBsBlSk/yhMTwZXF7XH9aE5apQRLRS/StxGYFB83eRIPpZiu7XI
hHwU5rOZAp7J4qymYetZed+dlKRrMKphjPkYnf0zSImvxw/B2hBRCGRLVeTHC0Z9gfHirnn5a4K+
Cq0uag5OhS9I2LxYmpQYtP/nn5zwvdtTPXCrSCTo3bUqnCug6AKeeoMytgFWj0ohZdyvJguQRWCY
BUjzSIhb+XY/QmzZaTGrvm36PtUr2WUlSzVeC7U2oZMY7THbEVSsisCBXkOaPI22XLPs+GYeN6xL
qsdidQ1HUQyF6hafa6sNAZ+db+TpHOeqZoEf6AvuoCzxRJfXV/SN+omDz1VXAaHVvhM4KGRzC2cz
YYkmoKj9oMhI9VPx2WIb9+iUsZwQoxMvkqQijkt1mbZdd4ae2OVs7XsotNld5IwNIzQTlW8uoN3m
JYfBMHCM1dg8r/C247ZMo88pfVyv0w6lULiVrWVe1Suw+gnlqcA4OfOwmSDD/I82wzMxaok0ngxy
elwx1FltfHbqWvNa7fi9EX8LYcY2r5RRyC3JNPmFYCMZHUEn4/MGuN187t1cFwEnqOShjqikuxz9
jM6b/fqZuuuvM/M9eu1MT0wxJnYDXnyw/096PAczXoQIkVISXa8lmkkpquio5FSddwq6eA201Av7
tF8iSVonQkjQqh3GCUiX7G2qtf4j4kyCSD/Z7VzdcQtFfDWDRchMfOrS1NrO5udXambo6cUubklw
4JFe0zXboVwwC1KzJrJlUWYbwkse7pWbfVKLAmhgNA7M/VWDv+fXYj/e4N/HELWao1vjsS79kAH6
VqNQ0wjUfLxIQqKA1cBkjYifEinglN9xEEth3mNmFKaU0LOYuK5cAa8QrJDnUny5h1oKXLtMgY8F
n+p+lcm0w6LanqgenlZ9YcF0GF/WovsSE2fvMZ+idoN2nfRubCqJNF6z+GxqfxATUMK9dhxSghBo
Kmen6ymQ1OtFKESaxr7qfpmQTwY1kz7FB5Lc+6T+lAYxSmhYN+Kj0jfUKT6PFHfAqQZg4WYN8gCd
adBnqnT8g1H3coY4fKL0Qv6vRjUFqt5lBHfGa6u6YYUxEVXq86IltS6xMJh7W+qj6OMLh3KZyJlh
y3plXVbOnrBS6Q0MXBmj4LFg7wqgrX1Re4ZIZ+f1E0vEGtF9lC80p2tM/zKTvNC4tqUD9KccvaIv
gwRCzHoFi5a2+ObZG2TscKmdKlRJTcZ5/mO28Mt450p6GauaADgT7f1YkW0OU2fQCLMSOdpEwQFG
XuZkzr3X2ZfNS7MxLLLLQ90szxwPwDfFmyDKdYWJoRfaE27lCt3rjxk5vLkzT8I7J+zS9oLLawgP
tL/lvRQq5h0Dh48Nfy75ZSO1Wk7kwukfKgxpURTM34JrS0b0hCBotehp6RAI4LWgX+/hRL2paNGm
HGb1/JYWhftVfzZexVCH6mQ7zZjBy2Sk6yt5U0QBjBFPr+7ID831/685pxh2n69sB1QuEkAA5WkU
e9HatlOpbwnfQVBtezqB4Z34OBpqGOzgtUphWe3zFEydtWXDH2k5Oa7IWCGci3rUjpTTTEXlzLVi
RPCY6czJ/Ze+WKbWfHjv5RhstGk8lJKXfcBrm5mprj3haVyuHSPjKKICj3RDZTjb+tCJl17qn+oG
+vlJzzXnhkL/zcW8kOdFVBnsrw612MfHmtPs2ySM2CvVSPYFkCRZTrvD1LVuT6jL6Y0ao/L5DTTB
jMZfb449NNzVJy/tUkJR0EplNS1vW56O+9VEtBCSZrgA41SUUlvQIghAe4widnGRou9FbBi+G1mW
3cNtGRc0a5cDx0gtWh9pi2+6Ml+Nec3ao2j3VumDj7P6wpmA3BHip6cpGSz96XQfyoG4yH0Y1xK6
q2YfJDZVEIzU+ucUh96jOL2fpGOMTWmDAA4v0XHAWPmYgnzZTo13f6PhnkIBS9Dq+jtacwxUfBeG
Hm7tNUQbPDgAu4mUAMMitcPmqO56vWT4lo9+AW3QEz3e11apBCDMYxiZZyrps7scvvR1YRypDwSe
b78vf2wtTRVk66mD38AWwsO3/CI3JS4daYRvzP0hL2qO6ON3xw1oaUUxhbEL7m/KM1Dx+6cP6ajf
jJkBMg9lK153ZP92uHRLwSnWWbN5G5oYWVcpyVfXUe8HTGabmQzDXxrB1QR+cvVfpp6p1J8kDuIE
7Cvl6Y7NH4A/uIjN+2zkz8o3KYVtrS3YFKAVmHjX1uQ/c5pY46vmycV3mUPsROTB7kve5/MUhGsj
j4hMmAAyfkdBqB5m4YP+Mq6ekXVMX9O1nQtbbOFjrzZKTJcHRQdkkeas5lCYs1ZjUZIpm0rAIMW3
79sZPzUijUVA9ez4C2y4U5I7QyC4/DkSl1ImJQayjZz/Hvup/IxPKjZB2nd2rdLXRJmvMa9BxEMT
TKvHYDcIW/qPeXDRtXlIEJBY4eED3chYFeCFdl5pQHycekuckCuotrSg3juyAgk5FdO9+PTzOqHh
QKH4whtZ2rbdK18BxNOqAo/eoUjQ987M2z2B3zbrWuAsMI8oV6jVlgbZwKC74reOBjyuKF0+YbaG
OaXKi1nBhNmafC7y1XFKPW9rZCQ1/YojNyyEXOL2xskObiGRJsuUmhCi7d8BlK0tXVuWNpXtRv3i
AoFcqvfQge/BF61IMcKS/0IbKKypDPUCijdmhp3IRTOeXNl2BYHk7huopzni4VBNsOvIdMXT/1se
vcvVNvJ20f4SRqc7lPZC/cRgJsIR3UQy9I+SsZ9oqqmDoX7Sky7E8riRJvvi/xfSh+01wH6/HdGu
WyiLqr4kTmnOu5UhOMLwvLlatkkgS0EPp2yDSKvXLI8+pTYqaCQwSmhN4vIBFIfM4lLdeAuE96qT
TWQ7r7AG2fD7Em9btFgqviw77LeIVsbGiTJiKeSTjzng/Zn0AIxfLxbY3Rg8cB77w2RbJRzyw9we
iOKDxQPO9tRjxdtk/QntCf4C8iso0jjxagcEgC9gkI2YfDS4+xjj/h4QxKWlxqfSrx4Rt2uW2N7G
6D8KRXMU0x/3l2gBri+b0suOSXDERqc9D55T7Y0fKpnW4Yj06qdxO24qJl+9Ee81ZGMrhlK8+OFc
11h8xOb1wT2TIjbmuDdoNuGvR5S+rIuJJmGIvqauj2SOgCc07wql5H39WhoPm9oDOu1HTvbs+OeI
gONodBMLpgOFL6gNW/dO9wmtKn9005chq1Ci1YeUfSSRS42nFRqHpPUELctogSfiKeEEHbnAdtQP
mGizTyIF+UCZFwkf1wDZ6ql0Tyf6ex/sgmwktItALEvSlKN3MM4ZH7SBT6fOau+RmR+3Li/RkYnu
BE9QGhPrhU57F9KnO4Jz5GublmWQN4+YGkJJQK9EW88Nkkn9LCwn+mOooFuh6QwfXMNIG/QNLDGL
psbJEMwbyEzI+yOZIkhz+Wt1eewmWMdH5FQkZtQwc1VoGTasf4cz+ZJcUtzA78gb4H0L6vVWJiOd
LfqoDUbaTWKxqAm0/sFZ09o+VGn2o7jWwX4W51kZKBebXyaUGytna7Qx41quUFbdGH2aKxca1xFJ
nwoG47v2eYIZ/64nYEDyMryK5xIBqUjM5hr8cVb/+20bQD6I8BvhRF8kJOsQPitOrqrVMPf0VcCz
p+D5kCyiypvyKBD5TGMzSY6KqhZQInQAM+aSU55glpdn6pcemgmkG5DnQb4wIwVKBtLK/9ekCfMH
15pZ8PjQSyTqbAe2URmTCBtNG6hQvMmL9zKRjJy+BlTFj3qk7D/NFUqdmc3pU6VBLltNm9IOiIUT
oMh6wAGh1qvyCIHOgIFpd+yBPbVH4U7+zLVsbRvERy2SgNnKcI6Tq93fnQM6oo/4gSuIf0GYKqx0
AZIkfM/Ske71myhxUiKCinTacBZ3LW5RWeyadzBKAJa+L8kpu8hsNnGuUbpcJx635WAOT+E1IsMz
4dzejdrS8VQsYWgXeQV95xLM+6sfjKarX0F9GvRsGpnNAaLfT6SjvyH4AEMax9SK1mTJDQoThyMI
z2QpEneJjnk9BN0KCS1rZKOGRXHLo0PbfZ87JnqkopM6Xp6SXpxLYipphwA96MkaDXA8ixK51hmj
gmdHGvc4v4IieGp8+xg2Xd3xsvWcZK+S46fyuQHCjeWfH9izBeuFAxC/Nu4+RBRgkQa8f+6TEGUD
W0h9dBDfPeLXnDlAvTD7kH0r7IKVfoq4nSii/2DVO/YsoxpZGw/Llmph/uWAzaozwVeLCsYga1HM
oXrVU5mvnRREyIdRJ3uZFY1+DK29tLJt1E2OCOqn851QYxkvWSkRCoLe7zb2GYa5n0ah4H1T8fsy
b3HVhyuvz0Vy9rXUC8lZSu9TLiJiaLQImm0z5hCikrfHVc5y2W+V/8+Ooo3L3nisgsTQtwCc23Nl
esZuz01ZvzXn1n+Ccc/saPDXajL+bKKGMATQ6jidRVNssDeEJJbQZbz/TMSCS7LrGeofqZBCGnf/
AlJvkouxgZZVabYgSQTlIXQy7WFsj3O/QzS/GwvCQu7m5O4sget9+C4kJZrsRuvyYeN/V57Gdt5M
/kvr3lI+udaT4uVvQNCkFttkwDjkw7YJV32pOi5C3wO+IXx0N7wC0BfDBe9fOJSQ7cP+Eq2BoiHK
pVQQvswXgHZRNO44f0NhmJwkPt0HvHhFCNiucarW+M9tFRbS+fYUnsy7kg6u5jchd9+nHzJO4yWd
ii7HVGE8mYiNYYnkaAJMgdLDhD+X2lRZ8FrXVmbg4KSElk0ECIrJKKAE3xeY8IZtmqwc1FNiPJew
bGllFggPd//CTEC7PnUaOk4Gu9n1sbKi2DtH7yU6/xASTjXXvqBtwHtdtSubFq8wlM0DhqwSqBU+
PwpORorswbmYWEFtNnKm8rRyygrGmPybqh80izPwCfbMZy6f9N6IF2El9iUdmmqhDBqQ8RFlNN17
r7b6cZx8dYChfpyJrs9iNl0lG17dBGANF0GePhdogSLJGKBvhIxs38xrNdTct4nt5DcnmhXKhdZv
7YEcN9MuXRCeQImrYeoQMwi5QlPs02c2dsl3V9sNx/+Fs6HuO/nTQrDKuarbI6QF17n+TO9VrrKJ
tQtkIUpbk56eDW12o7VXjnftQFhQfv1njsRv/7IbaCmAXU09xGjUelHJv0SGXWxRRenN3gF5K+gz
Nk1UsbGWK6L491REJjZBw8eSdCdPjotfEWREIDQh6011ur3Os3d+zso8JWD7zVB51rwfE1G+kWKq
NpfhcCtgZ+CPfkIOsNMA7dwdea6RThNOQtLqxTjBqbCeMMuxgt5boe0G0sJnYRlfT+zQvHgDloUW
ptNaALZIk2OHt6M4SoUpWGolKHW8g9cAxXY5zbfnYwwhgPXKRVyLG4mGSq7HHCPyvcBdUiOVkm/h
tGAcSFLZnsL7z9933fpvZduZeQG0xLZZ+y2UkQv4M/+62oAPDFuBpWMfjIIIODus8gIuZwdFq53D
1c1sFhjd9oN2Qp9H9dnTM8CUZjF64hWBD/N2UtdCfjsPHNMrmWRfzEonThQF1W991sRE1/tkFkWa
U1f0GHC6lLFTg7kWtCfiWGAqiwVQFBR7T6MCgQ5LFhC4AGbwItuUmmW97JoFY8Eljzpk2GxmCkfJ
jFNpCSJNNVlI8xfXbKStFSPPGA/sr1nDjq6EgufbzDZaZYwktWfbejxsuq2meack0UjpYdDm3Vw2
rJd7gF0NuviWlS7kIhmRg34Dj4uTwG0i917hiolPPKosEAn/waUta2pWUuUBxvfGQ5oNPEd0BIa3
GAgs7LDrbNqiQ+A6ChVbmProfA1S+YmJb8GALooDLwKFFRZ1IW3CRi5+mmexi58p9u77uasv9eiJ
3C23l1YYpiWhnlvzmBAHN1Ka8ZVa4Wp6SH8HrG8wLLmg/W5dO3OREAJghmYX6AslGjHWDE+ZEsgY
ONFXxBYu6kwJ7yDa/kWlVFl7zqQY+CkVuPUxwXywkjSJseGWGWO2uZZwASioHlET0CHY7Tq28XYu
+q+3NtY8Gvbq++KAKIZT/qUkvmBssGoDCM+lGK1c5xfxh0ii3w2M/1Q2sDCgu4igNhK7+7LgFjjc
jN8pwiUWijr2Cf8gQ8wiTCi++M6fwhcki1X6zeFP6U6bpelZPB04+CFv71Zz8HFHdXSfw9//eq6h
YMvjigtZ3LyA91UdMpg7MVaVNiUOzR1QRaQFQA1kA1vxGYv34UrJ6Fddb4nE8SvuPjj2Q3JstwzG
tu8TeRO0MB2jSwqd2JokidTGNkXDUlHjTBewR8QdeEmNTGsGoTqI+G0AWz9gSRTw/dqSiu5H14mo
rSnldLzvbpLmt8OJ5OuD84f7+1QgR+xm/nTQi7iPMCCXTiaYcGV1OA/d3A7fM27HSfGtOnJSObXa
Otn/mEHBu80MMD29R4WxUzVLsU2I38B/mEZyR0GQj4nfzhAAyl3NYy+IJWaL7xXXFiUEDwADHxRp
TTrhaBHBkaK1aZwFIdgOu/aBTuhOtJyjWXeeI3gbi4FYDo9unMonCTFAtc4wKkL1PQ9omARM6aIR
J7IxzvJGts6my4yA0t28q5UzAFEY5In3UtDc8VrdLU0CYPrOHmHC7XSCMUw5c8JxcBJyJCY33X23
ReC2e4+zLjyi9bZ9kCvMF3gdoGK7ZCstvEVD9Ms6luhqgzYoKkJ7Ctq9ZoPzo0UgQmEm6wiykPri
mBMg4+VAtQdsk2WvAZ3PlrcHGd04G/jptWnvLL8lNbin73+GD0qdU792N0dqlAWmM3aR3KofxBuy
fuvIEvs1Ku0F/SRyPhH9BcEbp1LrmluQ8YH8/uej9HNNW94Dsx1MXM9z5AeAzH/w6GvJu/VnnmQM
lARpSBwxRikap7WqqIF+rDzlt9zecfBuNO4slOhZdu8rUje7/tclg0SgzGrOJtr/QjURKUu3FDyz
6IW+HFusO+1HEOwgvkSJ3ZZi1OW4eUsGo8NkfyV+mYwTIP+mRWnAGVdNpxBwYKaRFrxuHqFcc6N7
ycbIyFFzJahrPnKpJvmgQkyHq4M4hYZ1oP7vMSp7LqhaBWHAHAiymFHrsM+lr5ieqmgWmBdbVV5m
FfMemSNH1aSQyyIfUfzaWCVCz3BIDX6b1p3h/BenvwlwN+wPsdo/RV5Wc62SDbmVrlH/JW1kNkgD
6UmCvP7kYwvE6zIgUj/mAXUgvGq3RL0nifoqdO6IoeZheQTZ1LCStiCZ/81nyhmH5Kjkn5M+q6iB
h5fRoo3mzRZExiLm9G+IUb9u0pt2ll1HiyuYVPdMU92FPxPkVYsp86QBO9ear1vpbCMqSDHp/RGZ
QsufkG1L/0PG1aLQhqG3LHyPZslUKoCe8J/qpGiRAyVJB/Zkfrw+ruP8WlsRKF7aNVZ4P1k+0Cv5
3glvxvfEr4h1raCryStVSBfSWbYozOqIAJ7BsIeyY8j14jJhsrVI8WU5qTW3Tw11un+KTT+WjzCC
fEjlt4RHFlLzE4eEu5oYzFuH8tMGJPVCtkFV7twSm36el8PpKlKPOuf6TdVxcNfr4k6PhcvPgXBC
bhr6nE7JJ7xwmj4NqxWqpk37b3cFdMrRjs+xkdSOjBE5A6aynirCayyd8lwP8phTo2j9VqDn2x61
JKmK+SsxCLlIiceDKs3iM7oJIhZgtanyZxwjsG7ez7HDj5+C0Nch3jW3tATf+UMK7i2DEkcAQzG8
kaFTKvUhQV4/ye3L9kI2vP/KoxtDKIdiwTYccepbL4ISVFTZTl559wjFcnqj59KXVrINFYdjfagB
PiHGKKo1V+6YWXFCZVe22sl5V8eoMu2pXPYIf8htBbf4PdJtzqL25EabiHz9jKWnB+9orLBB0csA
EbtHgiXZasI4CWL3nCd7eAKu+lp6GYk1xeNqma1zH7db0YPbyaZ3l9ylgVvHzeHbRP3KO2wkEqqE
3CBHxnpeg1Fq9xW6ILgqwy51fNtY38+UQDtA4O7bfJ5XsumM/xD5pMRxPAj17lUyYfmDHhcBdCE6
kZXJ4gLuzzGKmMlWdr3GW2tXVaOkYW7oVkKiqxGv6V74cyuf05BzwpPlGHFHOdbkstZWM/AKEe53
lOIJDno4ZToYY+XJUpEvfzWxlYBiDTbZ8z45gM78RKH6ETTW2Pz155QbcTTgdPvHNroujlEzwNUG
h5ey7YLI+CSCN3TrDWJAZ0iC45xPn1UwCoLMMqdJLj+/hM9fPF8ybfLjesMzbk164WOuuPWsmwQt
7CqE/FWW+17tegvzLaO2x2AuQ4o8gp10CvMRLcqNkiNu9+p0V2S+1j46QeJdO7XEjFfom/NocV2W
J/ZWJtwJn2caLdPKgp/94pn85DhCkGdjdxvQivgxLEuJ+WELUBJV40lpO30C9xtxUzBdeOwcF54p
lzFOKpGyi71NNnakTTbhrTRYZolnAaJ08cu6Fckt83s6lDFEfBy4jZsqFHeMAWMwaZ/nyacq/Nwc
f78EWNedWjF4vXfLquPbRDJMqQlwZS4xp1ImTCRpam6siPq7RsOZyABU3dfhrMlqbBTeHhwWmV79
T7KNGdI1xaKhptw5UveTyRvtHm0YUYhY2yoVqFgtRfN386cqwn/23dUvzVrfk6psS2+8BEU+dvcc
azsdFfpMPHM7aVHn6Tw0PdsV+UitShUemCEKt+X0AnHM3vYeu8NzB3PpItsuiPcKzbTVwUxDCEBk
JrgU0YLvVCO+vRfO7GYq0r2B6i80ZSFmqTIfy9hV/fwTI++LJFywjyjVRgQnTKykD9ApbV+38s2t
SpJZE5HlEXNQd7mXGeDAspKfsnxpXyDQZZOATTJU2Q9mCDXeyscOcHweV6QtIg8Iv4x44d4LHO7D
UElFnv/WypAm+thERWTJvbtk6W0PsA/ViGjTB8Dgq6Jh3rhS4pYnZ7P6aBuW/0cEEgSZtyMf0OsM
tLVtmQRQVkEj0qAxHb5Y8T8ptQ4H81ILAThXCNJxAzcF+/xk0flmQiB1dYW9PMb6t7b1DYLfNCt8
Izz1x+TBR1I7Czv9/5/zzuZM4p636DsjdEG227ySOi8J8bDooGk/WRnv9vMoabqH1caPsTfqU9qc
v0t6hdlAvaztbAp1DNhQXC+y40O+mi9buMbRlGu9S6hNfnv1S5mrbrMlonJpn3q7oTnvPJWuFDwv
/T956yeSAMNV/yZ3NddzPF/hTSCDODlIT/+ajymgDK4Rfbz/QiztDLNmIbSxfVUdiLvsCK1+oc80
L2k4eoeiFWevr1dB9klbB4hNrnOBJpbnIAhDu+BtdUD4gfqbFdEq+Bex2X4RAV8pDpARVN/yjB76
JwRbpLftQ6eXWPPglDJINv9AcjsEmXjNvmn9v7MKddrAAoeC3DlQAaBfTiIzqDSMDWGK8kDYWmFV
KljxmAvWw6HCyxx2Ndw6qIt2vCYWT7GNa20ttjz+JVn87qf0eTMbhmKI26BAVode+DDuik6QRCJZ
0WTtFvFC1zWr5sH8ddVy51B7Or3c19eTKU/PIfrMGCAemqlWyHIRGu7Y148VqGqeAiFi5nj/0fV2
3SiQ9Om2AGCO/UT3bevKFEgkT9YjSfAZ+H8QfD2MUiXdHj0CESyzwTB9ZNwTK7d63rsGUPM1F+5B
hg+W2OcE0c71gbmcDMeoMR5KdpcciL9rz/X0UknuXh7izmYBPkd9ib/bGbXmMui8rgOGTWVTFYS6
Aqj2u/ZlOGwmNBfHIdweSLVUJw2U2vHC5oeI4G/MigVzuLrP68yg9TnBp5lIGGjuv5SeklhwR4Oq
pczSKn6C+v9ZeUrOdTROc9ZOnD+8yxKS9CrLYmvdz3WeT9kY6+0HLyWNXoSryt2EPO5pD5fSSLTV
URppkR20pPxmb8atNWTVsJ3rZzxr0Oq51ROH0wKtMgmkyp7v03Zr2G+XAfqscybXWih3/MEEUv39
fRCScNlARyoYlZ+bnqXbtLJKt9qenBrtQys9KIJSEcELWax2YfHkmjnsCcl1molwmHXO3u7pXdEz
rUbQCgR2PMVj3P87fURZYf3/L9TL7y4I+GvaD4C1DgMK9Yp/thS2B6/G8rpBFPanliNSbdqGpuOy
uXyvvTRC2CddxiXxn4MHyPt46Wnjt/AZIMvi17isSXliqaPFDg9CyOaTQkYmxJQwsmB3o5w71JQB
dvPFRVixjHmqU0LXYe5aMVY+h6Hz3w6xfUBUB8dKwTsYRV5627wYHIDIfhmMmxLLnevEWImoBk/k
6nfJe+pcdKAFFPBhxkXPA+4SjbdTvLmWfKoDCB4+XwUNBfquYN406aQgZr6yOmZQntNeBEHN6zde
lbJkPg49wEfUhwYh4geTGwO2tCzVNRufbuyZ7COsJn4zuXFFwtiiKe4Ie0u4iG/LdrSKPvkpDSX8
Hqii0rla6lonyjZBKihIJYxQH8Dq+U7AxTHti6vhnvTf2kXvA6m1zEZ4AogM6jTqCVly/XCsBodZ
fGyYrQ9dHTzJMHaAcV05JyDoexkPqMziKV7w9u8n+Uv1vOzScHbpbNJs6JrWbdryQB6ydZI+o8jW
uDv55mMdGNUKFzrIUZho
`protect end_protected

