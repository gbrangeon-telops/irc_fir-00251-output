

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rLWvNa4xmaUmUmTsHaZZpmf+vdo1ZTZAwtQ7nnw7ufjv5GWZXhLdNQy5Q06lrQkoXFZkjYTdRiP3
F6m6R2KGJg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hpohmRSyxraB2TfGOSuLyUSGGabJEMublC4fhU+HZ7LC068YGUgk2aE7EHkl1WtDE9Bb6v5v3Qg9
2I0FD8nMKFfSIsem6wrqx6FPpal5aJB28sq90dkao5/Iru4xYelKhv5oyEvq5w9fsErMuciA6N4Y
mVn0CtqFHil9PLQizOk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e2qQeTSxab1fevbjz90nhYXx0vSvMvWBAXsx6NPtcQGmGbeJ/S+FZG17TXPSmNs8pJl+7MKHcPRl
s4fPkRF2q+UUqzkqGrUfIOlc9iDcSV3G1jvuqC/KwL75+As0dV2zHDw3g6spyRgrF/QyMSev2EDX
wNjTOD0D7tDHqk1b7PsRTM/m5LabqbFbAoaZk3OIm0Vx4hjx1H+Kj+5LKlzym1OWRKYofd9Pxrcb
EMUCk84oHB+E99UNC1xkjUMB3ggxmGGz+tj2pQbz0ixGcWE5awa9i3czC6zJ21Sph72Xl+p+aRC5
JcGtcY8i/+JbJchaWispPX8x4NW4FjK9r8JxKw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vltTKSM8a/zRJ1QJ/9B9ijVL2/YbgBrtsRTG74WarkSfaW1TYFA90LAMjfijw4Dh6V3t9bzMVLiX
18WW94nb3vnRj+WAyEjiDaLRKxJmoyxgwsVe3baoS8c9YLsCvI4C+2FRQmKh6kD8j1o6xfJUhYAE
QHwYAw6Gh1Fc1rWYuMM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jeozeC2hZr+0l/LK5n/W7u82KI9P5tCxn4L5QInLhVBS1ZXkJv19EUcHMrHeYhgivoQ0MQ86TEXP
Iah9T/vQMV+h0mk/ZiG6XOYby7qUUR5Ipu6A3NdkCDCZw1M+w2At4X13RPUlLeERzh2uCLeznee9
UbtfGUHB0e0CGrBNEj1LzA1bbcGeOcLXMz/DrWLUmi+Iv7nTaL15UXhNNoh+XY7m46jwFf+dQiLA
SkppMG/4vt/EhyL+TyDlc4FcuyPEIIJCq1gQ6KO1U+4QL61Qp9FOEA7sAw8XZEnuD8uyPmi6wlXt
gqJWUq4qR9zExL8yZmy88nYYAn2YB3+3OVd4ug==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 123472)
`protect data_block
sC29W943LmQRahKceKC9oz49s+eBMYWXOYB/RMvMmgtO4QJaBd1vDBt3txxBiZqP5IUxXo6Wso7v
rFnOzoX/EvOa0G0ulGXf2I9dJdJas2wMY514D2lvWyoEkd9MbGTxBSecI1h+8pwfX1kF6VjuE+iV
xxRz1L9etcdCzqH8U2eG13pdJc7St+YvWnwhjQzp+ELyiuOgP3QfnLtYWvFcF2CQI0EeTHceAMWi
316fFeUlLM4qk6W+H/tQSR2MaqODBhRmCf2401l1BoPwMlQfsyr431xqMd5YpeXInYYI/yT8S4kJ
aXDUrVxTR3MYDDl2vO5xlNYWSIaWbFpk5xdUp/wGOg4NmUVxjJ7KF8kTTaC4qLau+fXRmvssMtva
8faaekNuYEH7IaHodY/nZ4u4hrULt5Bw7T1VUvh16Km/vbcVqzfhRJDP8JWR9ZfrVUo8BZ1mQn6h
vVGumteJXkLWnWQ79tjM2I1ATtbqk/FquSPp2iVJdAvAlFbc0FbdqtNuehRZCNOKMMnFU74Jqh3o
0jWLWoF0lJI/49M/6E23J1Rk6E7ljQLfe+ZuxBMN1sHfJHLBnnqIZBLWQdkk/9C7Kcs3IV2lmc9d
1zg3OEcej4NC8ViwhhNUwGEVW7ut/gzXr1Q7g25CbNrWiCsr7WKOctO8eAAd7l5ZwdqpWeivFAg0
khJOD0C5Gb6j/rHvKmM1W3wAmegLn9yig8wkeMK7BJgWA8PmVaAtrfM0Lr3/0Olcs7YN63h957Js
Af4207t48ysY/wnjIeNwsuAvUtv7eyz2awyZ8V2Jci2wgsChLNKAVSBwwm3MlU4+bFuK8bOZOvYG
R5P6mU5d/Xavl/+M3LKKO1kfG1PcfHVSI6wHnD7J8GRYAGCF5dgzTb4sdLTn35uJGDm/io5wtqB5
GQOdewfw9n5FUpnP+2TUEAKzxu/ua231ODwQJhBLHWYIJy1jIcwv2VhQPhGsegqZID/7lj9tZgrX
Edz54bcaTG9AfFsY93Ma6YVjhwVON1iWM2s9cjs8+O54Zl/OtsVwlJgWS5CTNdZMV0/uwwSiAJNW
eCu9Cz/Xsc42xi/ZKp3OhFpS4bQwyYTSObs01JkbBVEa0P4yxscxrXNdelc83/guOfGlEnkbAN/q
VEwXN5fPROxgvdJL2oZi2d/goLUyN2RJDindlTEMdT/P01YAPP1Ci+DKv9c5+jl1CEeP/6Zr+Lgt
JKV7ns5DpgZzk1hTN9WdFQEK2kAhHVLFi6y26RpSuBF0S05/Z0RhAR9BtuamLyxa7UZ0CxJcHdKX
jUr8cyhbhh9QMLxnfdILgl00uDDN07JRhaQPt5WsOFyV3cmvxQxwAqTD6ppfn2fem9GGkG42VogW
DFWHk2ukkpJD2fQOVaiY1LJX8LVNTqudUOFSf9ziDgq4ZzZ9Q/Q/QWErBxuqZYyWdRxTH3E7V6ng
0vZrvwR/bvsJpkpSMB7PmX6ONGgJG+N4fqLuWPbqqlN5mWUJVbxXx3UswBbQUFYR22X8QQeBFmK/
JBibZkgjPArDyD80o+IOhgFqE4DLsARhQOOTPxBIbGfhq5tLskY9HH8YRsgOczmnkBzNGLi/ULky
sSxt74G289VGd12fJ1F1M8svI4vmXRGx2QwrUjRYimwc/KGzGNbBMNms4DMYwzUSTcnrhqCV2ESu
6ubbGKs9UGR0qML2rxmvewlgiGpBFZHl9o35xRv6RN6Kn3fPvGwZ2cxZ0GsX0cA0OMQgEZ/SjeUP
gVA0h73xRhetLHh3mUgfk4dTMygohzezxyCRR+s8s+zwS9CjL0HzJnbwmdgXVFlUgNEYp31dmebr
CZW+3rkTzQJU+B5IKGK/mFOzVTwjwvcCHVs3W8MR/bDF93vuaDFiDTV/gatxInktY1SZomZQkyrw
7eVTcVkyn85dh9bgbuz9z1PUDZTtgJu/CgL3krpyVp4BLKpIWd5z1lk2CF+VUTa/VSVgOmv5DIHn
z/UXFQkQmUdhbZHym/YIQ0ZawGhiBvBr0Ca/GyAA8W3lMOROUhC7BPbq9z2ys57bIMZ3/lun04jS
kwqGQ+pMdfdQhFvNpZBU854RyJrx7RAPVwSGs5DTOXfXqTcIsSveIcx/6BBW3Z9p8zCKibnS32E6
8z5kdjQ/UzvGtPejKGGGtt+CBm2w0Gq8RNbcFt/vxYeE9E1kA9Mr40s7000FAqh6mmKl1xcf1ayh
PhWh6MH05UmB9t6kZozH3P53MmZJKxtGVk4VeUTaiO7j4ovOWI3RlESx/LLy/m3rdmoTDL0gH1aS
VrqCzjmZauXlrqztevcg7nLMFcceLBgFD9xfZT7oUY7y57BbldqzpEJXYFB2bSt222QMraviTN5i
10cdBfERrmC3x1e3PqQfaziBUwfcjUFH+/QCU5lK2lr0OBaEgxyis0RdGjTizkI98o3lfLiy0gM4
ns8RirFvYbj9gm/95oH23JAYMwwr0OMvBGHpjGYjpcVZAnMbeyQZvO81f/wRmMx+euhh4xxbBH18
TDvYH6eT6AgT7WxfxBHhwv6eaJMzwT7AfDVlgHlA1TMRVLrbT6A5z7dlEP03jfkESgbRlRatOx9A
FImfJP5+M9Q77uj92kR/ip/plP5nPgZUgOBPrMLQOVIwJuFU0J+5DO2FdJbN7gh9EaCyYQd58vix
LRdZ6pkL+m9sKymR+xVWL3nlMbn5ZAAiUuoH7OkHIwDaJwdGQrT/pgfja7gc4/MF10L7C7+ZiNkm
2JYowfpiWBJflkYgiON9c9U1CbTdiKcuhHsuB3tMjx2bV07XRx8cxjkKuY27cLhuL+efGWk1SXsr
uFQ3USd0ZZ2CGTMTvjvEHCbrlSGRMQCvQjEd0bs//G18HgKlJj1798FE+FurN58ADCwZWQqkAdDS
qI+JEO3OBVKrHtWCYNV1KkyULFU0gwMPNv7rWxDkeUhMAZoyCro2scQJXLXIxx/fUlZbdLI/rt8r
YbLttERZeDd1ytHwM/Tqtnukh98JqEBIOiJfKLsutK71bKAwsJwkM6JfxSESt2SvvsEGMOPzzCy9
opWQIPEK/9Y1H+LwCKMxRa4G7YM5ydeh91Fh13YzykCBSzt5nWHLEM8P8xSnfcSmyQMuHO3fbx+z
z4fWQtT2hqRKgXcZAwGFN/Oy68qRwdXnOsXnKP9/uxfPeHPiBKVp2pYZo2CIhGN6Lwp5dlZ/CCuN
6viiD+9TmnSnsvHgZGTcBZtKQjgi0RsDobxVMN5zOJCwrJIBrTcvh5F/QaQ8Y27qqnlHeNWlKPPY
6POo1yar+rYHBbfNPunJ9MvLL2w9EG4sBq9ltDzdsXHYxnmNnnpkUnNKGEiDd3gf3MbjJbK6i1gy
wFdgiBZz6+g/JfUw++MYsQ8KzY7iN1Y2Q+/+Jc4Pl33ZQvF57wjD3ynnrsTGBw0gNLrvGtbEy3OZ
LRSYq7y+GqHLWbhBEwgOFOEgVC6AjHkOHJwJ+sLkgM7W6m3o5Py1QTjv0oEETzcNlzI2YECchgyj
oG8t9rHZXrmmgjBCnAvtcaa/Z2URvdMLuEHnG4zwW63Vx9CMj+2qkOmeipu/Fubpk0FqpBUVFe2g
np45feBxNqvhTw1MX40hv40pq3HzyRBaNt6DCR3fR7jWbB0Lh9rV75TwbJTGe1SbWOW5JYqHpmiD
mwcV6lMuy4zaFful2FS1jn0M+nqN8SUMSOrDYKX86MIe/MPxCyc54VCpVfU3W88kW/1/5picLNfd
4MJL+bma/sxlk7cYt2DKntGiUh6l9s1Ox/VrZmUaL0dIlL8plYdtwdV1gpVCEZfbWPzbdzRBDqs8
VK7Tj6bf9gCU3Wtinktz8vxUuf5sStVPiWPMLWuokufDLNdKNMby8IumP34QkQO37PIOLIAJ7anN
xw/P0zcPJau9VvaHI1i+l3FwOtpCCdb+D2tvstc3y8xjv5JMlQhpeKLJWaUk4N/HHqf41mIzTZD1
A0oeWHQf66Ig3jSQKYXT3hy3qMsHsRZ16k9+T+9xDvrNRqQLGFU0zfscUpu32nOlw8iWiVscMy3E
5bbHsgiaUdwA7tthxYGzI5aPUK7z+7EhiI+P8FLCVcYIV86aLPpUod318sjPs4Gb20Va8sCigNc+
P2lSR806PISKcC9N5PjudJK8XzCzjsVvwxbQ9OxVSFQ4mhev0IL3xarA1rMWTF5SLWninqtGAHfz
9iOp1NIbswvJ2XniAVEK42uHHfdxGP3EPxrpSPTq/h8EBpurE9/lU/x6eEALgYatlJODRmx4qQ/D
+gDohVLUDHT+O5UpBKCnrsDiJ4BAn7IGooKyWcPKsBdgMmA/3idTFcaEwV8yvE+I+EzAJwPKUV/O
BuutjUhsyd3jEI/+4nY3PpUZWsmV663adU7xDcFoYmA0MzvWct6g8iSaNxRSqeuj22cogu9Mai0R
Y2oPNhFU3CeOemDfQlhx/PqSqwlOxcDjUB1pk6v9u+kZt00lPCooAfq+/IyPd/AeJYx3HcApGSLl
4B+9W6BTYUfdPk4PsSy8TF9c556pS9djn1J7syUAps5Ln+Dt0fKS6LqekplPNrZGyVcdAF2plb2b
Zz6exN3AbuFYq4dpGbJ1K0VsF1jVf+bHP5r6M3bh+oArUSD0KAMUaKgaYBzS+/J/EBSFomW4hW5D
Aev/gpdLgUnp0D4tzMqCZwyPJeURalOGZvWFBt3D4usheNM9187JL1UhOh45nm3CpEALBLoef1q+
bYlB20IJANtcW1888xQ+RcvOXw8MuILuWlz6ZKdSe4TFGghTarLsEuO4yBhdo0loDEh94VaYABnO
tbXNe59+havLucB2K0OYF5U7Moljk1cs1QGm0UcvR8FH4TmU2slabS23PixLv1d1Famv1vjdcuaQ
/vK2A5ptm1TpBY5+XJq0ynrLgZncu34UFJDYunH3o2NFkrgoxI9Rl4xhAgFFQZpA/HwqFRtgqi20
yH0fMC92vQE9/R+mgdQJtpKUkySgzlhKBswveJ+DoMLN3oH+yS9wNQi2ruN8DL7j31/G1Jeqf+om
t9g6CSwFF2Q6t4mRwCrUH2rAl/9/7VnH9jq3orinx+hE6UiILaZ9kCHTMIuldeRt3EFCmOW4qqGI
zUc0NJf7sakFBSNUqQelAUazdFvdj57UXfmk0pQsN7DL+XT0HhdZGSZ/t6KsGIP2r6UKvk5wpEu4
DicxxfFP6k29xZJXPbEuCwdZRIj2gdwKZoFc00wlqAzbzpw83PSgTdQH//zLhWOpaCQPzOKMW8FA
XlSv456Ehvh0mMnECBr1wW96Jj6k2B9jzcBad92byOoOPIuAFcrhaPIRNsURUh2Qm50P6i0S/fI7
sdi2k9T3xZ/Yh3P+tesN6XaYMzFd7P7TMYNnyLScY8q1sU35qPSDyamW21UbpatM3XYPG9ddUJeq
AkdXq7sq1af8xaMwjfho/CTDH3nmOoifUu30wSS4oEkBSf1CiUKWhScGihWmFp0sJQRkKPrG1LWM
Z4SMUfs+PjCw5PD4Hs2xNelD2GCh6/cYjJz3z70CxizPm9AVTU8wlrWUjVusvX5fKaiYBnZUw7kR
dneGDRD+cg6/sbJcEAE0kbxl/qOr6fKJYdynoDrKYm5huETyob5GZxYSTNyafv5Ks0GtfKXH5OAJ
cF369QehSbypuYFbBz79I0zkKo95jNtl66obtX9eC+y+DDPecL8WogM/JnQJwWPVDNFkAD+Vw68O
YN7np/sV7srMBUGtdAkJvBPNFCtCMvLM+H1wIH9YK2rUy9hlOUBtp9K7VnarXzfIwEDG3N+tQU4o
ilFfteMzYSGFGjBViBa/krouD7OtGoneesubbs0w3AuSHOdvaR0VMkMwl3kEG4T+q9ptUDbpfRJX
cMBFVIFq6XFSQqNIJVLHAvh0hX1bBUtSwOmr7QWYyF+qDN0lXX7QnsDVzYveZb8f49t4taQhSTdc
jjsegU41RhhMX9TcBolF2A/rgyezrGkjb7m4qsQBT06PtpwFX/8Qp8Uy8yk+ql3b2tK6YDV60eTG
BxIi2BkkQqJCYy1yskskyWFdBkp6efrwpIKpoyfOrKi9kcFLSUCwjvA5C9KeLrX9wJwfqk8OYCiy
Gl6ZPjkJMajwgZiCh6XiYmooluZjBOYkhkro7zyg5v4bY0sCbD9ceGj51uC8VSLhApy8nvSkKBWF
k5Dbh5VST0F57XzSghddIIR9J+v2kt4tyyiy9v0LFfMpDiaO+A6diQ84r5szwQCH9YMpzY2Q9BHb
2SUnIWa+lbQdREssHk+qLfJS7i6RGSpk98jMcAI1ZaG1KNJQP4pgBLqzqblfTRTeQwRoIpLzJ55S
0vcggxN2sa+l51S0uvhb71hwZjPuT/M4XpEZ3MtBibvkqBYJ7UvL3+/hHxmPf9KZACC31Ug7UGDn
Yh7N6Gj2SobpNMv18R4gvW+MJVgwetqkIVBb4vEx0DpBdEEad0v9Ho2ncOJnMqN9r/QF66W+4S6N
qkndtnzkLBrEtNMAWec65cIVsHavc/iM9LpLaGYJc4EpZYWEGqDI4EyC+xRkxSity2aMNCNJaVw0
xrZ4Pvgra3dh2rO9npM91JT/veLqUq8Cacp4cdiu8tSgEcG0k42ff7k1uNL9U2AJ+M9Rx/z/uQza
e9TSs5Q28uKFRQ3NHBMX8EYFH1DfCtC6FEW6q9BQIzI8cutb27M2jaY3eJ63hSM4iN5lfRb6fUOR
5xt4D/LGgGSegciZ8QpNvpybarklbyiubwjqsdQ58dQxs7g/VhjorebQ7jWgq3z/qCbGaAfTdTTC
G44hh9Nbek2pCvkIHPCAYCJmFF3/A5gM934/IIr0jvpRbbeIsNNwJxfcLmAbkdM8X1+06j6RddIl
CfV7y+SeeWZJPGTngvB9hmkcpU7muRBN+7VHK73zwyrhlDpnds3xY00aQXBqc9kPakiPFnuKJg9w
tak8eP27aEkUhzWP2F1eLSQPS/bjQktc5163Ezq2IaxnorNodf/k9NOVwf6KAxzoLbsTNst1gZHp
Pu0kjDKiqpp5w1oXheuySEhIJH2yjoqGV8K4B7FQ6nRjRoyCpjKS5+sgfAQpq+RGmbwo6+xZYeqA
DLkOWhKZYXyebDIAImPHnU1bGwLw+YBPgAqy7CbMVZb2Y3NK6xclZ9NMKJmQ6TReqI11gix5valF
XFF0Vfgm4DFjDf2T8GtFqJCZXSB9AQc6cflMf1J6AkptsvbP4HQmZJ+NgADTpS9dltPLLREp+hfC
fDPEyqFkTruvryHiWAvZ4eQXHoP3vnlKzPRPRPw1+B4Br7soVqC1NAxMuMRYpxIk1ZpGFgarcvie
1fxF9c6ERiUApT/t8gqigEKpbioIqL8EXGkQW2UjsromWUuRYsNlAsrCv3109yhvuKHGJw8Qu4dT
3AnsjQd1u8Snz1QvHpj63JhhAgZvq1QuFmd+zzZ0OIvwD+ku/06/ZShzMveJTQjnKZ/WpjNhYIuZ
0TiRBRqOwIVUKTQBjK3LKyNpN27vxq+SDmXyZ44ljDjA9q4Dv5Ch2d9bvB0a+Tuz3Vh5rOk7P0WH
1P9CD5Kkb5XtasGRnvXsmeMtg7U6tsNNgwBMId4TCfwK4AvfCAQjAZ+rt7eDAf3hbpcVnN+2Xrdw
qqBnhp7dKC8bwheDJK+62lnVVjLs3XRSuZhKC01d29UQqnBrsxQfjuIAAJuhOVvJ1jKT/RGWgZss
h0EVRkn7vtkzDy5Ulagnob6XA0SeQOmkCpM1wGbBojSPhI+BxeQXfvotwRyh1OgVNodznx/Jbfg8
T6QTsNWa0c/teT3fc4sBsIKxWa4Cum7BVdgBQtS6N6D5iM4NfTmdlnhBnU5XOarOeCsVJ8fynM5a
YK+NEdnt26dtDcLUvE70i1yrV5nctba7ON4ubdfYfi/CQZVn486hcBgS9T/vwaCbAcxu9nls9BdY
wBGRxfD78/ix1Cy7KnMgK52In9zQawqByT1ooeaK+lWHLV5iT0QMJ4Thr9DGHllTMMkmW3GSmQm9
TXW2dOmboCsm8tepzMmyPb8slNUNQUg9gRprFHV6f8RK5ZMsbPchp79xZzFEpd25pyV8IlPJwza6
VDrZ8h1cvCSuXXC/7Xxpba9W4f6eSwtYXkjUxi0cFuTM/6F0PT6zi3cOYnVJoP8mSc7zwZjBotOw
ZA4Hld/bEBW+liKg9MJj9Zkq7zy5iPCZE9y1Ju3mY67pNfTHR4/OBaBGrsHnrvXFDwaCKUZVG9am
abUPemddRsZbZOchPEWi2TiAFznzaNcbnlyK4CvqHk9eubs3Tg7E3qAVRiiOPHTlc2Sguih1T+Zi
amo+1Ni+vQubH4yCjW7f+2xfhj7/owWhw8D3osf9oHvS00tEH2VbuBsDfiCqTg4A/m1cJQV1734D
xTzxosUoT75/h2Fc07VMVMYSHJgnIJHQ7qlFOHuqcqJIA2kA2b9K6IX5Qy/EkAgK2P4kq2c6lFQ9
Zeshrn379oYiMBYjVhr0/QKgU/siAddX5a73K5g+5C9lTbS9rzwzYAo6h5IbOu2KkuH812SWRzuX
jRyN8jraF4lpuWzQz6mnwR4TBWQM7E1So4hS54atnnZduX/JFlfH7itwUGBBdgZuEonT7WIwvJgZ
dAwSYZtH/mhLY6FMufpM+cezpNCOfFlBTGaVO5UUa/2w84WRabHkDobO5Ftjg6Ki7iJ35lj3GQSa
LEa3v596HYbzCi8hOItut0tuAARUJhtaiaFXSZIgJsAjmnULJT011GKKM21wHV3em5F7oN2hkHgB
q6ZlA5GyJWyupgpAq1rHyrKMKSmRJZqsJcBeip1aQ82fgnxnsVG3+0RW3hmPf0iWT+vnqIUsz+wW
H2lFMnKlV3bz4ub6aHhfS8c+LVRMYUNVzQ/LIh/MiznCqh9DKon7qxVBakmxvqU6TQWynwVls02E
7Nn5jo3A7B1Gbzki2GmPIClsDsQFLlly52WrwJkgXsh+3qAdQwxJt72iGjo1ivSZ7XMU73FsfPpa
aKV23BLQf69tO2jAaUreMSLf2vc7BiQKllgBTxIlHB7I+H5MB6uWzrRFgdYB0+bO1HjZQ5PhBW+Q
mtbVPOx6xLw6lpv2L/HpUaPc77C2EkljQw8Hz4iGd/t4R8y0vuMscgFMQt2YX4n0MMc3+xf/VfIv
WGrlxZmU/pVe9kqCpdYIjKWf6UsDboVL3tqRq350dvB3ZR6K96jcnZ4sWiEfVCJIsyrnEZnuu0Um
G+WC3UR+DZKNMGCfqIypol6LPsoY0/a0ZLX5clJN+1XG1qX7V0kESxrpWuRt2PflMpD89Dy6+zFM
Sd5TUDgA8gaX1kO3wv4QcsY1FrT2jAnIlH6aELY9+BSCbOjNGcCFZ+ttURBklfvpymY2NgKEs8YC
O8FCdinAo4Cr+ef70xp/2N+hC2VJ26NTYBRzM/w4DosavL6SVu28yERreXEnZg1rOzTUiQwkO10F
6jgutwErz9BmzUxmkP5EBeYdroM2FAEKz0nR2/qIgU20TuKrLSrq76maum3lDTOUEa5GNFu9TFPE
mw20bp0Cy1qPiTweiOb3s57YBZTfWFYQr5pKf2jZM59bIwZ76Up+uh+WxN3qTVVQ508YlMZXu+fG
3Mh2GmwK3eHjhVjesGy2+c7FvQkAW3o+pbJ1szuxEl0fW4zKP+6zxbgNChlBLf8oESrL6X+LGw+L
XmOfsNX6oowlqMzoWhLvyrePzRfKLTclDQrCzScYmEKteQu2GKemk7uoDD5U94Rc7yqJjA4UZsLl
SN8ukRugA2LVxUInXmdlLglqk/39VWI0SLeeGX6pm4ShuuzhjQPgAj4rgrrGfxu7aKmcb7GpqAnN
42bjOyMH/0yMurX81v72FsBWjAxipLHkm/zSL7Pr+eg4NzXqUUtKYc2bg5kQ0iU2BwvXrF2lZfw3
aNobvxW/GL2VDFMUnLbBQibjf9CRGJ8ugMCBofSbNSHjBM33AVAjHBzOjFTvbfKcLIQjqCRXivs6
Qee94JNzmRI1r2Am/AbKeZAnBSpVjW42YgPLtnKoqRzqtk3sFqe8YpZ+mxtN604Gz/4uYudSthWv
r6lPx6C06uF/+XPheL+DnmtB0/meNyPUgGinqEoKQI17YBUiHCd7JKFXQdig9myrEEiy8v+53Ejj
suDm54NJmSJvwiSkQzZsa4QmzrJfp1aGf/oGT16RFMhCoJovwU+7JAeBh2wY2bBNLf2DWdprdZD0
WGtJrd+s5g5uTwlYonINvTuYt37xHgX4/fq7iSBG4DVjsi6gkYDj1DqupgvLfSVXqxburO9J29aF
6gnK44NhbxPVkr6RDgUsE/BW1i/ZoLpllrCRIsxyblEbTh3g3AjPgz/hf2jnQjA/ltMhNk3seUdL
FAuognOqo2Z99/ef5NeaCpxDLY4D1Q5+fOtVe9dZzG8CoO9nxV8EN8Jp/xUCDwWwlc1EilQVY9Uw
nPsZnY4Knz8gERGGARzSgpl3hxJYSKyGrEo4FOppI26plnOQhNpkB4xpoff4HHv8g3muSKuw8VGo
45+CdzEOOqrUkvo5nBL7ey0y10eShzwcdq+4m4oBL2yjw6r1tpk/ufwCVQv+2Xs6qCaKVdTCeBoF
hShg68/Ynd0kjY2Q9oqWXb8gZnqGcMJaTQrG+BEjwodDLxLM4ls/aW7pmTl5H64xTCiNkdSRcUiY
q2DNnAqv9O0+do+oKA4SAGY9JLk+uGVrs5SktDbMipzu1f7dg2oQACcZr6hv77nxOL7fxNbT/gLY
3hiC3CXz7fTmOr8bae9TrWoHWoxktFbIYiNHdggnpXvKs1qlzWIMzYmMGSkTpBKuIXomiNVT5/7Y
ZLB7/nE43xqcirvivcuk+hB/hiByk5LuRjDw+BqXX1+J+Q3r9NAaS9WgFkfQNPENrOwKEA1mNBNj
Dxm89d67roKtOOqzOWgr/O/udJ2hM5q0jkmZW0r0kmZ86SfSTzb9kgfEqRz2DFugt3SV9yDf4bpL
ZiYIk5gQEYJiK6SBdssGE/C0+ak7G4t+qcqT9sc/MXD37gZwDKUloEU/huikqaJM2gXWK6/fyr0Y
oqYQiP6QvWDFJDhNr3fb67EwL5dV730YUiUyk/T3C2nKtVz9Je0zHKNx9CWIrgmco8JCSy0T/g7j
0otcBB7bFB8FxiSfM/KYQ73h+jBII/nnU40cd6pj/hpehaGK0mfco8ZMZyaYS3pA6ZHbLIMxqWGi
XYQmz1JC5ySiWOKX2HeZap6yVObB/6lGXuaWbn3WX/mGeWwnryzoKwSQWmGXjZ9hZxchbQKNK4y9
Bqoh8rjEl/OK2JPS9kpVDzNz7fjA+0NbIk2LQCQPA/aojUcyPrLBil+L8xu/bVuvKzAYSZv2N3Gh
xmIJNL6/s93z/IRvCK/DNLsEOpcVtEeayBQ+z4bmpSER5ZUU8an1f4F/oKNdzrWBo+rRDXw+t5EF
LZE9UVu7g4VD+EMJVBloCwdYLQSCh/EjRpSZq4lkh4yu00+/NJ1G0d1hq5hyNBuVLSyCv8+r//JL
Qym89ySu09FH5P3FDae1Z+nbSsN/wgdyG0UcTLQUr8ZoPIw2V4BnUnF5r9vYYgxjsiKRaFmwOdI9
OkkuYRCFUZHGTwo4oOju2JpIc+tVO5mq2OzTXRjil7ptUGiMODk86CuvbDM/K+snejEBUyCl2TJ4
uRj5GDVlRmUtc6N6NSLMDEaJPlCs3wTjWjCho9stPOgwrkvLcX5OZ03qYGaDX8Ri0rMRZ1yBJ/+d
mUwwkKyT8JVBVswCaGioz6lgQAWUBJGNr8ZWaFYYxQDeLnWKy15psLHsOnJyycSn/x85dRNJHSDw
eZwT4AUcAUGZdzvb/zSCrsQjOid3g7lUNhBdXJXyLODoT5BW8TT8faqtmeo3I09jHbJtRSfSg7lX
7TsGNxf5sxVRjBdCSOFeaQFQdUh2PY9jNqEj+Kn9aSK1kyknc/J1lDZVIDwAuFukMnAj28zDH61t
vsVrMXAqX4V+/TLk5dTlXlmNJz1wxy7uNjrqbe35LEpuRVnbhw2L/2kmbPBtWc3AC58+Tqqnt7sJ
04YhIX+C6o6iN5VE1pctfRBob4mio5zz4FqW6CvyDTllux1gaDbnqubz9qp35ADPfkW10smXKAvA
2ODWJZTF9I3au3VvDYvFURNX6WCOT7VOKLSdfdgPYswEli/zpgWDMxEBvDETvFpGr3fiUv9Da6Rp
vtdlo1grhMOV7FsRql/5/qNHmtJqq5jfkmxAAOUh6SmO25j1vGcLSfql6x7Lcd5/8Dod0t6O6lVm
Tab9PZUEtFvXqJJyynXNgaNYPHkAlSZtnc+mRMs4VtpOUulcOn9GaMJBJqkEle7dao7vUsk480xG
HqiUp6+cZ+aSRPt0Uo2IpCLLVIrrLTPSeGop6Y6bDhVeWx+Jaf4VRmgIdGL7c3XnCwOOTU3bxPSG
dAZMp3PlBVytirkcAFPVqBe0NhjnC111Ki9WQ7owm13e3tZxtcMFsRAIYs967kgrRN8kCoZfEKdk
ebq7QbYxkRnbGBGtVRpnxhHYuqpH4RIVzJrhCjO/i62fB9aP1UOj+RmCWbAV4uHMVdiRf4aWpNF2
Ez2xkfaSI65zMmzufkOzinlL0Rk9Ng2yr3Rayn6AOtadF/ayS4fTAmJPOL060feGokY51M4NuyDM
65A0AfyYhOdwAV557LxK9wieuJ7t+7i5O8O5TP7py0aBahZzdfW2bgQXLKkuSaMa6ejdSuNSm+4L
cX1j5xVvJMIP3wvzTw8AxP0Rzd1LXcSJPmWbpZve00SWSBwrP6F2ghRnOdm+2llsNvP1s3IERiB+
2XWdWBlRrL3N6tQ+taIsJQLotz2QzfpvFQmZNyvHi2qLkay7gIwtLwWAxC5FewIDJeBGoFW9clt/
gK1GVoDbGhEPeK96EHovWO/QRjw8amer7/DkuCh35APJPc6MCVDfVGvNRcanSBDkHZtwQnrw6Ayh
l0X5GdjEB8ZBLLYj/PUQ0cqpGKfBrSul9Y9lZh4FDYezSOZTUkyXRH7WgT8SJpIQCU/G5pBQ4jwg
P5dXLXGx0wqypfSeR0ngm5BEF+LmpUbcJ5I9vTnJ43eFiJ+ThHYPJ6PvFm1LACgcQJhD+8gEsOTz
PVCPFq2sZaygfxJkt9LXBCXmZxO+FfTjJ7gOA89WnZziGZigpTKig9inrgXtj94LsVTnH3T23nsG
mNRTHkf3ZSUgzVj0wct1hZ7LcxHxLdrZo6XiM41S91JICM8xU5wH4om+SQmceFbYJEXtuQ2FF9Kp
iZL6rVFjDyn9ljK8NOAm5sYP1XiSUafkNQ4Ns52K/A7V0Nbbahcyf3DMcTp3D172nxDhLIvZP4CN
N/anHTEuaLOkyOmuy7A/1V80EbAIPm/ldmmmNRj3Wv8/PmOktUvrFKnrMrqRDfgP4+qZqBi8TOZv
jTC2oW2DMVxIxRkfiLu3zS2FlSlUjvkwWAgHYFcW/qHlbDCaUoE/GaaaLYVVAUq6rB4Lzw+120H9
qT7teL4kzhZbOTpv+KNgAQ5ioz9yLwDM+Wz1RQ7UCKach3yut9Jte37HENA3zi4hl4v4Fi0fJdq+
gaaGAL2ySAc9fG+Rtxbd0UUn/ehfzBpTFx5Eqb9cYxPHA+wo9bklTXiDDXrS600jCb5GmY32Ra+l
hUa63UWnxLA3kXt+3bXJ+yvrQiG+0cqaimV9dsUocqAHYpl86eoVVbkgSEhfdFRzMFHnlbP8Ownz
tY6lG++JgxZqdzl9GJRPikImEsNRaGfUZaEmPCFXAfmbzXd274ott/TsJlsENU+2Y7Ot6cYSQE6X
tSxOSve51vNE3yTW1/xFzxPC2KHet7T0DnGJUhZuBDOehwdmkRbKJxvcLayhy05nwuq3hYcnhuVe
1ltyVzHn7/dldXlJRmtoX5S2QalB/lkmF7MCi4CK9IVg+b1Hl3gaHxV67iWmz0aZbjEc5+wvgqcF
lU2tZthNv7ornxvZzmxMZosbxPWntl5ND7UUlXu4klJRpBSc249B7NdzEFtLRECDgtd8eo8HXiYW
1zWf+Nsv0nm0CXtwa/UpMAFqJSB+qbkCqBN3PSmSzY/60EcA18Kkn2r2WD3nbyogSKxiJokZSqsB
hGAtI8hEoJjgmP0gy6XKdQ38Dc+TQ0hHrnE9u/Gt8sdwZHxUiFER79ct0R1Xk8AFR8uPI1uVW/k9
eO7783uohm3eBAR56tHWqfViIHaNecmk/f+ZLM33b2erWhxYEhKiYfZN3fk+R0SpszYw7NfAmov5
sgeCjsb8m45dRuZFqBj7VynzNIOG4ke84wlhsNx8Qy/bgttnrHenRf0tII5rIwSzbIMM0pXiQKsv
prMJ2wiV7ZPFfiN80an4MUmdoUphhgzopzSIBFG4hI5/dT53JUjA1r0s1qHopY86iITxu4ZWQ54H
bTueqiqNFatZZzTMAbq3QhnLN5KeqaO4Ig0sppFEQqscTuVfHsrLlVORENthRRqsh6qNvBf+yxYK
RwugWC+H0n63TIO8QAqcIfmanSFriCvs53OaBLWFwuuuwIQqkPKN7JeriYWUuv01Th8xIHzup0Iu
4jjp5HtiS87+t3QlxHt+9RiSZ4vaq4kPRoefrrG0bPcusVSDqGRMNkEdqxpFxpFSQ2wP503R8Exa
anzSV9avCrL6vS5P97/UKPSJR9fz4/dIpTxy3bmT81VNkwa09zv66Wi4K+ka66KaxVfpnmIR0dLl
oRuqW2GF8m+GsdbmCu8Riom9qwU5WvNgVhBiWcmr14Yx17Sv8+MHqhkjpwK93PxZh543RleZWOmp
KWmOs20jTSGqtw3XdtR30XMuunhu4d9yTxGcegpECJO3hjqHX8/vxOmZXX5pRJZVL0EexeSrKmid
UpxA3zwrT7e0opMx1Rh+LqM5HXU4j20JbPunKKt27hvR2VKdkDG8CORrXAigBIjXXcY4ADd+EU+b
7udNsUinBXnPe79NwubBkO03PCKaWdiDlwrFZ+hAK22B2nx7pymc/1tzKWrMs6+sdgJIhEmlnl94
EQh0ynHwPX9ItRWQxyYRGg03Ir1c5XVCgX3SVurBAf3O96mgNQNVn7yWD3gcaw9e2ApELM2gYXWf
0n2Kk1XtUV7Avo2ZREd3BrV5tGohf4aaP8K+5FYCLBcjJPtaFIS7zEr0BjEVMK5E8mmq9aLlScq9
l2cTRdTpi34q8BvFwk6/YHhLTei3JVERX9311c3ZejbmydYjNe/hDrkxRCQZfqP+r7V7T2Jw5SXc
1maXBcaiz/wH/zci9CMk7xZujL4SHEsiX/Xdfj4JwtFrAngrR4e13tMEmv3ftDsiHMlcwoyfzwup
D8LPgMNBov8snEKuubdW5ik+BviBNRF1kInjavuq/bzQT5jVMwgGBWR/blFjIX+kBlp05F1HkLwO
Kyz72KKFDIWYGDih2Y54E/k2EK++2piO/yxgpeu8tK+lrUi30solFqFIqa4s7Fqzjl5adkew1M7P
Xc2gG+4cBl4THEMd0gvpa0ZScO5WAZyksEqUn8V+pvRfSew3gd6BZCeGeS82DoymxdFZeaJ2++1n
u2rl7pvoputmPysi5Z/5qx2nEQIU6uh7xx8Sd2/VrTiGxu/LbslzvPpKB5uKP/NxCf9fuUEMZSYT
F9oKvEeRWJaB7mbeLCmiM9in8catuot1lXMR4k5WMp486VmR08nas1OUxoIRT7KMqBGStJ/t4rge
hcaQVaY9JPtKdFcxijdZga+pawB9/HSTJ0sAcbScUqpMn8hoT9zTyUnInCVF/1WQHuB7Kkq7NAtg
rNKHwOzEYILD9VwN4Q30nXL7lEE79fqsMLN7tLZOqKam8mHH87RJzX6ROCFJXpGxmxRBbl8lBbuB
1Xq2MCoAHK312uhHmWUdHx9FbjcOfmEswCiJRrX8hIjJV5bL5CujHCSCwea+1Jy0IV/MaMNJQg2h
XWN+yIh4X+SkXX6BoqbWLirlUCOz1BI/A2JsVG+dxgV10JBZLcq1jAjOEUvnJeDn4FHR00qw4X58
V77/Vg/i6uDwxrJjlwpooGw7jI7Xb1C30XOwyBZtlcLwJ2nnNlsXqAhlxOm6skVzkFQx4Rpy+CLh
kPX2Vr7twWxMIlgBrSDcZlPAu2JyKnpnWTM2hOl5JA2SgPAw2AY3SxX2ARcC1PF3X+Q6WJlAeOoe
WnWWtYRhkuib3PIfu3zYYlAcZM+LMonijD4oWj5JhW1uC+A/WCaAu0ylitjRj5+RD5EChgco1RhQ
L9KX5v6Hr+3vCZLOlszgfxQKfZlD6SUu9TAwsFaGjAJdqoIc0CvfCGKfDp1W/qN8M/ILjGCMiiOm
ZftjHz84nwcjYKr3B92N9u5LRBHNmHs+0FgBbJI+RBbiGfqhbIH5xB6wgUF0tnVCwxiB217aldZc
+/YbNFygUt0Nm4733wB0jvtg8xNO2KFv233PfbDoCuJjxSPHb7Fq4tF84p8OhywQfbBmxwYT48uc
zTlVG9FRtM8R3sp/YWpo8aNbcwBqLnMWeiW5YvaoIjcx9MS4qDpOaGg5y+UBN0F4prUXyCnIGJOr
IYKkkmG6JjTqo2VkVseTxJjGlE+Uq3JkmywtguDtOVH/7USlFc8DaW5D+6prT36U41JZeXTob+5X
vYleHSxLeVWJ7gnu+nd0T0Rmkm1Ga2da2DBuAIb57Te1DDuSpyJOaGJy/K1oZ2rVegfpVdi4DZNR
0NYytUNLe5dzPbAQaxH1aV37Uf5+7G8TOsjKhwQdzi/s1dh/bHrtKvh6RYdQGXXfHO5rBSRxxuJp
DN6WWhPT/nOAFzdGp98ifp0CjeIqyOZofkuFIrH8QwxIjn3la6PMuC9Q1gfDCYVGBGJ0lFTSvge1
6YFEt0LK8Lv2ufVEJswNConNrJeSU7QsQr45y6RZzoOn37D6pkvyf5jk2PF+v2/aW90yKZD34c31
Iei5pBIWiSY7YRSQWK0ULZ87GN/Rx1tvVjmAgc8b7XOm5YsnEpXE7vtg1WqsH88GP9Rv/u1mI0KD
fnupC1yE16VfXu5pCWs0+UtG8OoSytGjPbQh4KcyGTdI4jZjDyIZZ+oRVMIBkERYfygKOF435bx/
VtWhorKhWBwGOrxL8ZHx7DZgh4mpzOGet6wYg3BraC/9klkorl59IhM8KoS0T1eXh9EiN5/mQnDw
4vndONJC3AQLgfz6ozvbmaXHCRsWj+IA5GQfMTVYnbME1yZv013c1go2WCaSp3VpgDBiaHp154Bw
X0NXyHmox24eDtddKyrMCqKUszEN0bWE1ckyQh2YzyKOq7sEZciW0PVrsIVDKCGHy0Ct9XsX1+kl
Kz3vkuNj++jf+InA5kymH16GFOfxobGJK6x9KRb3/WvoiuWrRi2rhwiUppiMhMkR6rRN5cbjT7xg
LIuOW2KKS0pTEe2gI0ldB7avM1Pah/lJuKnF8dtczV8Exjw1ncR5sERi8VZTcyfnmdyJTb+6Tr41
2oEdhcbYmxP/3jDqcfi08pWEiNfdYXB1oux5QNHiqB5xjP7LRc1aeLs8+qjfhuXSDXSI6Q6JfNVU
MbVelC94WkSurQOHQIzJFU3OthHZb4zXyn2RWlyGOCsiRPmXqreHBB/i/RV1/vaqJzIxIHTgF5tw
ipGvb+J+BKU1ZCLpgZL3KOpAYtHAXigDIlTWeF5WLruDOlRmMI+5+EvvvjgFR5OwJZ74dJuk0Oz6
l2+ITfu4t64HCt3NnA5qjhQW0bdJ+1pAkhQY+E+5ZYaftJHkeKKSnCMOH1y2WhdKeghX4BvDRhWk
pMBAqk+GD8qIhEkhHcmXgq4byMI+OvVzV7H9v8Hqp4S1fj1nXMUBeUX8KlYukDivtB0LnA3wAWvP
idAfEc4b+5YordGm5usB7lbSsdotp8+7zhyKjN6AKjwUNgFydxH23c/tz0nCEFl7YzIf+yVL1tdE
rXgH4G9B+Z1Vdfabq6JSKsi3sDAPGpy9rXk7UZ9n2YSHDa1Wm6z66V/JZBEhTMEo6k7Iu6VtAuJ1
//oe9qSvUoILXiUXfxS8v/i67NF3DoTvt6NEORss3Nn9zuHEnDXdb3l1LqWYhL+aXvyiARPrI8KU
OC6MXRHfr0JULYCgJiwmBZpPjtAGzH4jQv4yWulrqQZXkHAMsfqxt6spScTrGdc3al2irY6xwaDp
4+iUIMh2YDp2y0eQGZtOEEr/R31oV+00IyE4P84GsQAMUWQaKSRrg7M4vv+JkGeGOFVlHgwDSvd/
qC9WjUnTA45/DdpRRQ5vJvuisGZCsXhwgUA/kRmuJGm6kEwlSKKNJTJkG/OKRhwF5Gy7pl1Zik64
zJWoKi9BDUjjb66BcJxPLhghI09RyFmSADAHGpoIiZLHlpbn4+nFNsGCnwEtbk2g6LrxNDbDfAYa
/ittwilxjS3dh86tNj++PzkIjnACOpVOzhVf6Vg3oX9HPi3OvmWi3LZcS/mpnaGGl1Hm6M9A0OMx
6nYYnEm+lXmtDrIYABgTWAqDHhgP53gZS5wnf7IkOamfeu8221u2VYdT7O3IkMfMtAvg15DXE1Z1
6DfDY0FPFVZzdibbPhdXuJmLBgsTTAtWuKsmvxxPystNiOgZRsoR+R666GHpjBM7BVPzeRd2tGhA
22V+gTxI9os9XuJ2hT+y4Qxl0pylR/HKCEAtm9TB7YpDimgwuN2bxo/40KR8FevciGJC4nT5A9DS
vgpfWzBeogQX24HlJXrxIN23bNEj4BRy8Wgzc1LeVL4B962Dy2Btp9eWlLRMEU1X9Z9KQI1xrdLv
pgi0rT4+rSfP2EPsk+E04r4kAfNrBzpuNOMDoJizqYFxj9aOwTgp+t8TeS6xVW7Yq0CpSGWcm54+
r/z/IXAFVdkS2pDEZAp0FMiQPmGKGf3hOeDTxw14b6f2N7AkLJ03ezKjrHBeXEwbzMUm1tu7A9H/
hh20psaMUE7nvw0hGrP1yTLo0+5VroycQ4i5MZQn9XGgi0mt+CyMiPqTzM2XD0EEUoZUe+Q8ti7t
+QBPGrTbRwdeLMaPuYWdwe+YL4MS0TJRXRu3F54/ocAwPbNMBxrTbBFob3LEhDim8i+VvlvCjSoB
P4H0V7bJJadW5WCVcqo872PKTvB7lyhN0ObkkA6iYyl0hMfsBbYkaiY7A7mDag2HnP8+HhAi6Jjz
3qZ2Ljpr/LfGXwqpLyD7snTZ4CfP2hqZuyKv+VDneS/y19kd0R9S2sWgSsRYDuDMwJ2ybaPXGEql
lwCASYghaVq79XEo3tp/YWKW6PkKUIE8JE1vgLSlj2QFYxaN2FpjxPRTymbR6mZ41O6YP5iFYUNg
qN3Al3XphhN6byEM/mI3xyFxQ4P1JV8V8EWwmL/eP6sdmrl/vHz3o4rTPTgwbY+3jrrMdQpG4lRl
RL63AvLrnP8PqmVTiRZC/8cr0l8KVtV2H7RBdzKsaJdLZaX+T1YGeMLIVupyhZzzDjIRqN76ElDE
4p4RHjpZNc1KI/o9QzKxOvhfi6+ZgMcH/9lf5nh5qPWCpqwbUDtFjeBrBYYawydNisFN/Ri6v/2B
KG815QNEshh+NIfZuOni3H2qYVdiq330tgNAU6fDHnjkj30pWzu9xuWxEQf+Tbi53lrCpvwz93Ov
YLbnJoJt0mPR65YPcYnnFj9QL5Y1XmnL8SY/VsRCW5vsdtUs8EeQ8scY/oCNepN7BFQt6PLxQURf
/lnCsfqiixzAJC2qnAb1YEq3Cdn6LC3RxjD2VMYC9cXc/OnYsO1SJxk3ebHhyOBBKIfcs0oHQa2b
lUxEcI2zwN3ysoKmO4hq6UsKIqGmF+zwL/0AYfMTK7TXyajW0Ilgm5TEYHFcK0YU04n02Ck1FsWX
YbNseuKbnDeD3bPlfdSLX53L+RfbRReaAVwApj5PLtXAF5yZC9TWm1wdrybEMx6klbV3VJkaH/6H
H5DCB09erTXyIbfGl7edp5o82kq1wNyy29qPsXZoZxmw04keYa0i+0v2K7SETdiXjJ7MgWwitaoe
GDLcGQq5o9NOEDWHE8ARU+Z/3mqa7yVTeJVHMGq5G4W85MKfW2Rc9HJv9NtQUUBHHQgYph331ZLH
J7Q8pAo4M5Db+p/8NUXeL/z0SlZdtc6ZsySb2Q+cBF0jgkHelAGpjPR8YYkMUr3qwJIvDB68p94Q
QYBDEmVQrUJD72AOegC1GNnwsH8GaRAWGU5+31GWO1Gu9obUtdAX8L80opuaZvpJO4HmYjenPt4n
rjQN5Ry/PD+fJR7eRuoJuQm4ogv95AYDtlzzbl2RceT97wtnEih57OmpROb2a0TyNksWtf+dIQ2Z
G/2lqLzxndJCvfvLZSA684TfH7qdSzuCia91WPoxxlt+ySlDWyXPHclPk5BS4yUoeyk3lV0zyoeh
H+AoNqnUGz/JfqiAJFSDv8piayqHSNtvlnuxBKxWrlU7BuLF32xMxM5EO5H/pW5giOSAr+Sc0S+P
XY5w2pTPsTYB+h29pOZgjPudaVGcDtxZSblqd/8joVgJvfaPqZan3lvegTdUCcGFV5b5QaqvLf+r
zVQT4RTZwTBWRDBxRpvD3DmICuwMKNSMEdLb0vQdmteXjYSo0KhKlIpsVdIAgXlRAyHFcVj9IIAK
7E+3S0/QUdYmULNLUbgkuu6bcKRIe2Fn+zhW+THNo1KtNatVXMhLxdj8E8h+lbKPOLNUwr2zrQd8
A/Ffb4fpCuL7P21wSI83saAz4Ch7D1tgKOGWq+N7PpMJwFaMqG4NHn9HWrTDeOLcp8WiLZg+8Zt7
Uj8br90jlyFyheZ5De2murcGtqmhl0QgLfVDG7XaozhSqnBE1dLIoajhiyAiUSccUDQwX93amGsM
9r/7AbIvBagSbY57WGg7ISiTuG9+/qWWuAHbeGbgEhYGD/njxlVLMDL1M0RQRbVsS+yXka9gIHw1
mdH27d4CH4bsWsx4JuDywPeBr/jey/RJgo9edwb2Kxz8HV0Ai987ShDXvMtb2641DniycY0LipfI
uuvbxXhzL59clM9DVD7ToHRAEfSDZyOw/PcZ3pwEU9vs/wrWHz4wWZMWjpVSsthGuMPRAbQgTn9R
v/jotW5GDO9gWnrVjSKOi6INiKNVK2LsbXt58OsoPb556thL75Xlm+L8LneH02SgwxkLXdMaxtQ2
saGQuEgX5aBO4oOlEySGeBujtv4gt/xk8vRDqsux5kFwCWiXb7PER/3B9fhPhRNLELhbifDS0h9Y
qmSF0aQp+wAlxYtkLOY5el3+mFA94PkB60Yzo0Ut8KE6m78GV2wtMmpwWfJiJbD3sZVvG8PoUFWv
reXtkvti9aIZWJuqq1bjFRzpvMNgFlEatx6MRcnDvUB5Lt6ummWrW0NxskUF9JkzPRE5ed3zxB31
lnUAFwOxRfocwkQb0Goy890bhIA1rCrR464kcbEnhQXHWyae/j0hulY2AW6YEw8XTuDoXWIUBfSj
vFQ0Yw+e7uLdPYM4OXg57tXDJbDVbN4sBcbdpwMD13PAkpIvgxWN/D3jBK/LicU17cWvZ8GrPU2Q
VYQXrEOdzHNjOSw6nbpyaHrmuEw4Sw6TJnZuj8q8MvsbLQdjcBqh+ItZYw5QErJKaRO81jjN9pl+
zbAkgnbLcowfcu0M/UBkMgvJLzGNep8Rv00VvNq+A1EvGOuawOwHM922WCSJl2yzdaLbLEgODvpG
ybu68yDif5VD555JZGSSODqOEZPomPTZmaD1QZbAICoTskdtt5JoHCPD10YqhyCMWw5lux5FnXSQ
0LZcQYI4J2RXsPqeBJ0mOlAml9GRNMKY4yrNUq5uBLXfSz62minfU4eO7sBDPwHYXrHFVx1HpjfV
gIxNCO3sD6xuw3rNK6OfNO64N//CisC9oLTC0+gYPKwNz+2Pqeh5L3rtaEPh5smcSSt3swpbFesW
EN/rVXS0RcOOE0HZ5ciXXIXWZh/ReaAca+d3cnWcfz2ALssyoMtvUuooP6CTyfimh1hfFWLiuM9f
by14LC1fHYtq5Nm7kGr1NBWAdlTVJ8nv4ZZaNLObMXFwKTACNuwdpEKvVXToIQle0f1F04vtMdGH
ZlhZ/4II/MW50ZaJvRZph5BCyE+5lIU4qYtnEHHcdzo4ixCawcI4HxFIKlROUn745L/xCCYKLv6O
LuNeQDP2ket1GSYFdO1VWj+trN+QEgqu1qZ0b9RBNk5pOsk7UlKREuAokY4AFFuLEJKQWQYYWvbM
AFrbtwt+x2KpTphhFwEpbbdBokwVd6vzQQqze0ylFci+d8izWv7OtbTjxvy6NBc6G79hFSVfrgFk
3I1cVMT91M6NAh5s+w63MdKedVP0N1QVJ8PAV3k0r/AZ4DdWy0akkxb7c4V6pV3omAa2y/F1A3ca
kElIHadh7ke1SdHkpTdn7VP/ReJWJBRFoWG4PqeMQP90EsRdXXuWWMmJ5WCscQEjQPZodA77kdq4
rW3HSrQjilrG0ZtTRhpcKH5aZH+J7do6jN0RFDw9VJlCvYDVPA+LJL8fQA6OUzERCPFaDLjLeoFk
rl4zC6pvL7Zeuhl+rhfmXs9VC5+ImPV2Opyr4VNoVnwXen7j8NZszgJtPWgMdxu+RJesH6lgEIrF
oSVWcWSI63WR5dFS6COtnk2rYYfoePjoXb5XP6jCNiY4qv+vIs+eVHmpPVLbLkiOiysGMftHskGr
Tdtm+19kKTaKcgOT4PXwRD4xAbwpvlzS1uS/OGQ7qPMDejJfzcOWaeY0rIFOCqs4ZMUdjw21k2ro
CqjVDm2ED/pHBDRXZtnU93L4YYbJqHkDfXKt8RwiM3DUyEyRVZUsYwxJebeH2I13IRgKyBAKpB6C
KT1HZNuj6N8v8sJk6sl/IbJvin2BfBCGhQdgTRtDJ43AyADaq6hXKOELNq3UeAU8iU4TWT/yz710
q+louyIXMwn2stEXkmnN6WASJPlvJgdOGwreLL5L35SNNJ6bsCfr+surezJmQ8bEXUKsEDkM76WI
oocdRCOe0LcYAatrf2K/G5X2OQypwCVcDOj/ObAVH71RZhmtkGqLyNe4PBVgzoIs98TAheDCsVVM
KK8RzgLw3dzXgFklRV1PVsA+QZuajMJB5moro5qUtxQXQewcOyd3EUmU7eHTgL8/BgvXclSXcNC0
wNZ8B18lSEAypyKIokUrrtozlT9P2R1l7kEcVOSTElz0rxrQZoBl1tU7TNbIid++KU3n5MFyq5Fj
kjrQ3GzRvfnRZxPDSqOcHUQWkNJ4KuFKkhQOPTwcBAeK3f1zx+LzWn9abBQPtI40VmqDJuZhWnt3
nJI2LoHSLLsDdU4+NgjH6kh0RTW5+aOjWVCxm6TgB6SAC9yIHIYI/J70kc6qMKpP5hI8oGpTGK1+
tnXrTeYHXFnziGVjV8dfrwVoiqEhYpHLkORPiU2a1RyAlDF52wi0KL/9iDh5t6aJ/fvIvZCzoUWd
IrgnOKL5RkT5eHYKyNoTFQkKCUiIPgLEO/adqBZriP0vJsYkO35EEff2aZ97xG1h9Jf6RLVqLA8d
i3voB5IjYnRJ9KMqvJo5HC6PlKASygh+0GVmMzGLy3jCYfZiRHE1+pJdnZmGluSxi0qJot2mvZz+
6eTpNDDL5SBrixkrNROUGgLwLJnGjIiVdbHSXrm8XDh6mHMN8COvsDvVjWpeY0e4/yQJRVtEVLZL
rXOsgjfihXagzqE2ILYKt76xo/sgattTzL/f9BGuxv0ORrYKTVUw2NZMBdJP8+MjAg6o+nhZ78E4
bmr2J/2I6h3hccf1hiZXmyJx784LK+XVUyowIFo1kXbbxFbuly00Dqg01AN5nSKDNMtOV/gGeD9P
8i3Im//35r4Lo1F1ajps3kH95D27R6hAZ1yhcOjMCoPpCXXAZKlFTRYtoEkpvcgWsq44UYNcRyNk
8SBv0l9hNfG5vxQlTdbamSw+OBCv1mft6x4iKwp9SNPTEnr953hxJ0oCHBb+bXr9bJGHPE9TefH+
C14+eh7aBvy1LjqTo/8h3dxmmfGP+D+sjN2OlcB6LNwHVjj1tj3h/MBqsmEBEOCm7ihbMIR7pa0A
dn2w5hhlojTwF6aqbqbfITaieT1c+12OP5L3nIg8g2n9nqDfE7+4qq/sxKoJwo8GndzPrQPgFnge
gFP2nugl3DKJn8q5Av0A2u5+5WEkQPj3LXEroV8THRrbKw1oY6tXniXURXacC0G6C5PS/hLvXOlj
rhtYGzr8Vtt/+W/31SLNnLzqLO1epNDh++8RONYp75K19Ju+T9LWzuIVNm4dg3gBEm7MCoKjF8r2
wVkbuBxnfJUscpggOAS81ciMtXN+X7P9zffKfpWy6MDvzRTn3huTDqMCKUC0AnG9b/YHpsFC7GGT
A0lKkE66wD0g5ct3a/77Grh1N8a5YKDOhOGhXzRv9LLJA43IBPxktkSlOSLlLScbspGakZy8xAsp
GfpBtZY5YIrhHl5T0bjsxBQj5HhyEIkk84Ru6dcIC7ZYu+oSYBG/W0Pv4G9709Pf1itZAI1Y3QOP
PHTX5UmUo8kvAjVafZr2QPOINUUbx745SNvI5/AvwzrzcDX8UaLfSJER8KSt+8Lcf+d0DSHAaSMC
YiT4nSWsAj1X8946fagd8jY/L8G8yjIczCqJL3lIf+Qch1kn2KNSjG+YgmtsKGKFk5a+q4LRnarb
DQXItaFYqWriweB1rdNO9kBNUmb+8JuJHBLRuE8dlgr6blHIGPaBokIPon8yZK5+2hUomSGWPmuF
1T/Bl04RrPwRkTwhmjANfVHOr+CN+wKJ1Y+mtn4gy8G+0LMtl+AjzqeR/zjKCZLsjFdGML/SAG8J
UjqOW0WOxORGHWAlSjpHnKd9P1DmU5IFiNNZSHshd/E3RYsw8ij1P6aqXUj+AsF8TA4K+wirJXEU
kpqSPeBFpKbTBqVc6joB8ZVIKk2wJH+sf+Y6P4cEL8cluSc0cu8B8IkxBsD5UQ4Unslb0fPBVBTI
GwYT6QugTxhXwX23yBHL/n4anU5vNg/oNFg+HmL3VY3OO+dnxpHpRPeIqEFeaKfHE+PQ20g91+9E
cAq+5ErxIsQgoduzRypvQh8Exw/2PsfVp1uViMWgQW3/bi5fWYCWiIvTnyZTnWRJ2aNLR0JmIz0m
agZDND2RWsE3HHELxU95KQd7OcUUjdCI1b7Z0J0hV9cOrDUTgBy4fPh3zzQfd6cXhApTWQ6i1XSU
VPaQgZUMYM38QkPXGxt40FOItjlg7p1FarRdFZ8xO6jETbLKKWKOckK6hjk7ZBD9iGPes6TVl949
e0lWEe/NK7zTt2MbWpZiWiU0myJpY1iOT0Vm+5gStysZ9V/tZAq1b/Eb8r/KN+vGHfIyCly6GSa7
xXLRRrsNQcCxTj20ssilYv4R7Ag/Idip6losYOfAJfTW4nSPytx+zWZdOY/vfTqO9okpzJcSqp/a
Mm/MFnpgojMVbTyHfBYMWzXudsZjkGupL3XhJ5n3cumAhGWXZXFcP8cbVlyxTauRqOWACxonIrPX
+EOjecABnda+Ackfpeu6QAGwThGLNkdcXco6tABXWKeuEqo1Qkl68Ocj5cD2+GfBB9uP4/GVWuxw
Js9jbZNRSvWKB7TlI7Z4v/FtA1f8A/4ibvQKyULjBd6iqmRFIKmQdB6ZKhN1GhsHlHhhmLVhWB+V
Maz2MICOPVufx6UrMTYDWvf/tXUcpafG9Rg4SL93HIapnzw7RwyhS+SvhOoFIs8eolK5Etx++QvL
b7v/oQv7E6tJcqwX2wzllv3gqgk8AMheLV8P/0OTHYZbNt23h/+qYUGibEzU7lXObB2Jo6KtxAU9
s5faTPLnVzPP3jNzYHq1nMZ5wI9qTEfIdVcf4x08i+fPLuaeLIt+Z0gFoZeqrMfkiMCzd+vodBVL
FjyEbv2FXtZTc6uaF28ysr0sxvOSlzgqA4nEHyEzzW8rVTJkbTj7AAIYMmk4C5IuAGbsKI4vg5IA
lPkYDUoeQoj3JmJQhFQtxYAtd0jsCQ9oEIxl8oEfUzuSv1SaKYg1y1lvbuTCYyqZBvSJw8MjnLUw
j3wP3TQMQ1862O0806cyuZPhAmoljfYMennS28soVmIAaIvHOR2nrsvvwHVEV8b4il/omGYffAjW
GKYciY5ycCmB6U0zBplkmLw3nNKWF8Dwc2ZkQlth5p9O5xv5QPo47N3NL5Qc0DV5HoMdkuzsjmZL
TD7dTq5aI6RBK0oxaaAlmF0grnnZnHqrPpGqMPNl66ltDHhlD3V4iVz8avXfL8u0nN5p1H8anu0l
w8cV2vIZVK/vugVWms66+Toy10LIuJ7KTg2lMfDHq3NhrzspbY9L071urxzLLd/L3SPpM3yQmoab
FPjioEoS0Mw3EsgpABDq3RuMBTvZIlF6os/CVVsAMjwkaAq973GAz3+FogxndnIKrclhzYDy7CWE
44FhUFWals6mHTMMn6vKA+POBuS/eF1Vf6nd8zEmkJP7a/w8LDzuNJjaNkg2A/uzQRACa+QMhEd4
NxY+ap5wHYofCtZqjp+JuTdjxmlols0lFSkkXOOsKz2OwDyypOIbaGknF37yeOjzM+CYgMIpatqV
QzOjWBgZgwHVKJtsCofIIOxQ3Oq8a+GpBlx5j97hlbAa8oSAyLMUzakVOuTFsuieVjhKpMHycWGv
Bbdxo6dOXw9Qhu8X8soY/9p1ReUCI1YTE8eDwYQmS5b+m1f2Q7pa4JKmXkZBVEzbWZZ7c2YkyNs1
YLlFuP+7mPLc+mXm00y/nO9GLBf6Ny8ofh/tpmhsdVFjVTZ2QvhRFldhXqSB1ZowKm8siTq+gTvw
PEUl8jft0EdnE++DrTLyykanIfrkTGP+hwhHlTLRTbDViXOo/Mo8GKGK5O7sHWetlHcUA4IcbFQ8
mrdN4p5qsfZDtlxJ1OtJWX7DBUVfJZ7sJdgcV+sTNTvEiJEKX7ZJn5ooxL3CjtcbY5WaGSGxwkIM
+bLzmUx7rWdSDbpSXEqpn+0ni32vOjRLr1y9gRkyHH1bze5ca0O6qfMtTLEks1Z80ulSZCY4wnu9
2CnqUaCPxihhszdVDk2a9UQbvCJpMj6t5B4p+tSF9sENmQbIRx2Maa9IiJPei43mb3cHYoeIGE2w
06r5YSLKFEgRMpQ3th2s+6vxR11Rkx6PnlvzjadLKWn64HvmIClEq6UiWMr0QBfeTp6JyuSr4rql
eOSZMZInyMpyQRQmsVnsaauQvfWjfsrZkJvGwbf0XaTc45Pijmh6hePQYNa9Qsl41aLUGVUWQF3f
QOP4JUPaK4UV4AzPrFmtXRxk4sCr3BLUKxmgrQWSdZ856CzbR/Sxo9C/cHn5aobz3zOYnjUhAhYJ
+kvmazGF5wV42ypqC0U/qlQjkDo/5ql5Wh/507i/4S29E75JSHpZKabS11ivm5cc2DQyUY3zHH06
yeDGXC+ciF5jX3OJBA85xGNy6EqmZ+RgB1wFSqRs/JXT9Wdk+EOCjwnzwCsDlxOOEdpmFlIm9q8r
jzbcq/ymzVzAIQoBmO46g6+bUDHRMVnUjn9nR3r+Wkvbxt0nTQ3uod9ae89qyqX014ZBLmWNaacp
J3cNgnE28YrCulK9Ftk7Txl+Cbl0Mzn3yb+WY36ao48LYCdOa83qHzqOep8+YpeDGLs7ZcustRxH
hWdWVRXvuNzgb6Dhk2/thrTaZweJq8lXCU+R9TeXSUwa64Xsfb2440yn1/JDBBt08cb1Sgq5/el6
LTh06Hpzle45LmdlG3wiBPe6T6rcZsUJCyhe6kkEK+KNtNDRNZ174CqBu9e0+GflhOaGd/+2KMJS
qCqevTkkmNjJCcCspr5aMk8KSM2xVARKDlMfKkq9JAYF62zAzoCSOF5ihTPiTVWk+hwIw8lI8lUf
ujPWRP0KSxLY+OOHn0r+IvsTZ0cyhJnHEuIspJfbPR6MG8jY4E0rH4AamlAr2B0pN+AwSfTftRf6
Mxg7lya/bt7mzhG0ml0dHd8hjXmhxTbI9Uq4hAy14Ur3lJgAsAFjsoRJdyJf38dZWyRSUNhx3g+q
qGIHVV+bo5nN59iIqSA5pcsIMHKCPWF/aIWq5iObeZha2YH3ETRW+sjbP4NUQNxIW/T/KHDXqXCM
B/KhJwt0ictphXPDgL7XtLY5Xqwx0UNkfBVH4skv8diORX7asitAS4DaKhKipQR9ZEY4gwwCMAvN
5+vQIaUFESTGzMQynucgXX1fHk0x/Dd+Cixh/YQrhMvZ9xV117MEUZF/tnFUDY9bY7N0KI6K0Y9j
FucEoRC576aj6wRGU2nYlIgVN8K17Q7pdmIN5QPxWO9QPhSJs8GofmDCUhWZ2B/iKhX7WPp/Rkva
s6qJ45YG+znlnjRTmStx50TcBAgzFqNMr2FcUrrcpbBAF1RuSKym2+BKMqLYwtvxGBfUrNPfvbWF
qRKma3vdkb35as8/KyrOdgxY6rkBvG6OQmlXM6gIJ335re771jnMy/6PoF6s5jq9IZJsoavpZQpt
z/aNVn/ECkwE1LMMNlG3nudkFO5ZVSEhGzADEIr9ypnvh03krEMgb2wn7eofq1v8EFzwZWZ6KFm1
6wsXk9cldpbiZ8QWkoBd+EraQjKgEhotMf7k1oDVerzsQqM8ThgvBq5EozgcO/gSGKir/d4ZonJY
Fnc3Ko/WnqbeKQGWVy/4GE6CcX1hpnGMvW7lVkHpIpCuPsyapIpdelfkuOzRR5iDiHMgDFw+jAm9
bG3p7cx2PIGuyhFcOnTGwJ9iYheb1HepOfWDac4bChrJZ7BgfZ9+ccjcaLNihjSjHGFKKFaSn4V4
tYXePEgQ8dzW8JVsLhQbkGym+j/UfWh4mvmlKmkpt7J6r2UoiaAReZL+S9usQUFY9TLuZPE6zKn1
jKcVrleJlXi37E5Lvg4Re+R3fahwkxqhtrBgnPSk+WEV949KRgOZtNlvSf85RqDMtIX0Qpb6dgo6
1XHrK/89CPjD/EuGHm9xeLnuI8oOcT/sJtudc72VBOm5h6FKurP0SKCwSThXk+XtYSzo9PYa5Iyc
fWRoW59CMFNoH16eVLTHM74z6O7cbhZBm92Nn0ddOLZGzFfxdOl+WBUQrhE9WV9UXu62YlumfjVT
Sw/Qybqk9C5Q9GNA6tNmMhFTy0yj0WTiZ7Dav7nmH9Hgu9OdoiYMta1QwG57vJLnnzHk5KYf5DP2
dAf4C7Q5WnqSbj8aJmi7DLjnXmmrrdYIJPZU1iecHaLThaiv5T0BKd2WZkmmlEoeIDuBbRJ6h3nf
34heQ7/EMEhh7OGENmXuKDKPOPlS5NhuHyVxxQWbJYnyegfYnmWLusbr/lHjwBdTJy1PDPncJjBr
5WBJ7mJ7JAiD8wt5MRaMmRFf3ZwZppf+Njh4hI3kuIjaARkBgonqCorwH0G/2WoHKI1T152wEcOj
bShUbiv46K+3KnnFZFj/e0I1L0+mosUTs0Oy42GeSK2HI+EhVXC/3ia/KbD3Q+DT4Lu+6NF2RJIw
l4YkohzHB+kO/7eOKTh0G5CbV7CPhYSQaLCfQFAWNySIWhnst329P8OG9cgEI8HpSdoCdA/MZHbf
jzlXqx17lD7HPnyVllHf17T2vg6h6ZRntpnC5PULr7J2BB8ltBWtHYWrNXakR5t4pAB0vlledobv
jPlIUdPViTIG1+qC1/LL7o5YhwfhwwUHUVra2TTCL0cYWhrHWQhp/VjaBFwXDghPHWqTvMStCDRD
Ar9eJpNvHsKr+vlS5ExAdb0u2JQ3V7H1fSRGTiGl6fRjf6mc1tLbudW+UMoiPorqBcpk6AWEaHgQ
HVQLjTzd6fIX07RYv1j4iW38Scm27SyKJNrerNoRKkUfGVv0eVxNGoLT0TDhPCPSQhnXGlJZEwJt
e2DV08f8UBrOMHKGsGnfYDuFmBahKFqp33QA/zdk5UvUCqxNQK2Oz5ZGyNV/z8ztmS8Ioeo+ZPwX
ZAAr1w64jcNiwqBBdz+44oBaOUO3CN8GuTsWN66iX/G2XrTkIORBeMHgpgoesjr6x6/L8ibZBAnl
n4lQytOsNajAKP6g7mbvaInf4HIypP9Qu0zXXRB9Wt9eA+kJVdUeiYRu553c4m6EehbrAwP/RY12
VowcsMX61T4ZLjRHoMr+zdfY00+OnNdjEtsnZ0lh9P1xDBiaSfaiKvIzPQirVHqF7AHkN0dttNSr
AC/9nhr/kUWihAt0gUvH6CrL57fm5saFWg13BhbmaEx6m+3NfUefRyUC+s7U71ThpEvvLhNduFQw
AP96jF+aEoNeZveiqyRJbMfnlCrg/XaXzUvO4tcH8XZxg/Q29y3M9jdODkjTxQ8VVoVeM1A2YPmG
lR0YvQQorm9Ww6LmnE+37kRfueLIVLDH/UueYA9OPn92llHc+vmJxoYHTIcwoFaRqECRj2AF7RF/
i9FoAN3d9A2HFGBJwUeeWGJOtx4Jgo0axgsrVTxsiVTUcwtDj2lcqZXilr5vLVOrbNntjEtSkQgW
J0sTRjlyiEY/v2xFt88mRQVGbEWlnkrjkX4hFldajb/t3kBA+pLMnIuzXvyfsIYvhB+vZNHE0ueF
OTY6trdY70tXyA2ugvxsyjjjVoVVR9tU5OlrcELcEwiHWjUnDM4ax38mF9h/nhi8jHUxAxQUelZm
ugzS+LoeWx3o2m7BJ5t+QBl7GzyrYXNSRBOpMDaSqispXixc7uabmsLgXNKXh+ocIf8wjDn6bMN8
fDY3yvkdZTyOWYZMrwiX/OlXUA3lzcH3m7flqfJIjRniY3n5c0FIyHh4SdU4P7eth+SLW9OAuf9M
Thwc8mHcV+UYFa+mzZLoc3vMbMmuii3Oodtng7/zxiMSB6QRhlh6DZYjwfO7fvV8LAswCBx85OtY
MNSgzFCRcC6cOkD8NPBLWEgo0ULJlOke2k5pV0UIEsjr5VhAFh5tKhTR6Q3zSlZeUOffLUOEFoqE
ZTrjWSUORda3Q1hZTH3isoCt2tKo+UXt0X8K77zZWqXh/UL0mDYCkzSHQRUx2+HuJqbhzamQIQUj
SRpLyRiLOXbkcgtiv4VfFajIGUkYXhyu0RH7X+5KhcQcbw3ye6aEPZvsTAer43hY+Ksxyilc0kHR
XMj0AA3u5by2DajTKquR2DOKE42cj/woojUL+lcOdfO4NqCwQlN5sXT2hK0yl0gvyvAZqiQnLZ3D
S5Ii/wIZVcq0WFCVZufA+PtrRazt+fDO5jVmFtVGB4y/d1MLUJBsJzjJ6I/07EQw9tb1UYZ8619h
HDNahz87L/48MXxfDqKKaVq+kk3g/3AW7GreXFgsxEHMK9iIf1N+YSz3wpka+Xg2guSm0WiUHGm8
umuYpdeL09xGcdeDuarDrnuPECmXMPQLbJX2t7uRtLYMnauXe8RUP3f7AJeQLvVsmJezflvxgPsN
pzESYOXtZVhHIvd1J3j8bK4JOseUsj5uIWTEsX1+HZmRhYK0o6D2o6BCvGUQC4lKOV16yKQpMy/Q
1nrzf6pj0UbnYs9QbMqoCoxXNd/S/H/oLLWRUhRID2qN29z8lDAOrGliuEqQXvgtXpH2NaufUl5e
KZ8fl95l/a/5roLGBbhn5yVKAzctz+3RrYpwR2DD64mdRXLnIJLAcG/gydk03jGvsTzSP/54EDvO
IcANgEcWD6zc60LFn9bm0z8qwd/wFrI1iRvBJZnhsmJ7luSxWxiGHuu1fSZguYbQtDoQSM6XwS5u
mlMhAkPeT38Ht6RQWG4zEqklNB9FUWtKUiIhOYHs9DWHcU4bnTfwDMQaDOrBfJEFlWdljtTji5Cc
WVzjZZRLEXYI68nYaP10ovhs4DUPKa64mebISyEPGmX3lZIT+kPWaXLRVBM8UpGcNK4FBEqEBySZ
qB/+FUORi2LtEn8/rBAoxm5RpqZrzZXTL/NaMZHWnLdu/tEXNXVWL0lvIUs19wc4lLwl9uI4If+E
9cEeLcuSjXqevmznyu6BVN+wIjH6iV7KZnVZtNLycIseVmeymwwzCjRH0iL2cHnGs8FLFi/4JSEZ
Og3Gdlyw0EneZLo9jrJTpbX6h++NXFi0dcDSbCZrbNUTTcXK3pGq8fAr0TUl9Sc5eW3G35+/uWQt
IkqFusACYv42sVJwWXOmyr61jeBD6P7Eup1D3P/ffIn12QSoxH0g/Awl/o6BwXFr4zO/yh86lH2/
LPHF6wYaIeJBc+a5OrZ7kXKa4uyNUQw4APzEeYbKfGIYC5itymRIel7zIo03lNr4C6edtHAfgjhS
fZT1igmSKTEcAlvXp0pkhCSVj3V6+hyrKuPQ/kM3A1l8HP3pJ2sVQsiK62rCTxAR3jzFe2WO3tdX
IBNqE2Y6NTgdKnya8P4+aV9u+fYXZE84aVNLGE0TaHJooLcmxPaar/rtMoh7cp7nIAaijROhoPPo
TupvT8G1QjEaiHb0gYu/r3WpjbNfkqZa5pSvKuSbKmcwAFfmPAXo/1CkA93svCVvcW+G7FHAyiNS
woHAJY60OGd///Ratx21t13RD5JmxHpwKJ1LmAXaFY9htwbP3KPcEg3SzOfT7U+Yxil/IwxnAc2Y
bRXfQ2e69E/iOn+XisjCLYGlK9KQIjoMcEV0Tt6+9FuHSsMhSSYf6YMWTWzaFp1/M8yYqc3hKNKA
vMOReEtROIHY7snOatF/iiYuFUeQ3Co5MlhVDGccF/MVACs2ISRjzgVHY9cPl+w8WVgZ17rrN6BB
8H8qKuENyzdLCeO5yTJ+o8Rkd9NB2qHJlAxFwCKJUtfcfjIIkGFCBBI+QxwxTrmxIgIoNoBULP9E
ukJkZe2jWYa95lW+A6T7nt2weC4p9WPkyJU70bbMlwA80KA75SjL/CDXQmcGb2veQQ66z9i5lxl8
4cwndHOeZiGhFxjCVhdT3mieUf2lAJYIfNyknoZW2AhUMGPL5AXMITyI4JrQKUjbafY9VRe+H8PR
HJg4lW7S4c19nmRNcADHezeOcSaUkC56eaZsvrfh8AwNafob6kf/lAvnMmJPDoBXRggpGIo14q5Q
hBNoxxMeZxNUXxVZcFDMiouIbxbi+ILkL8/hrtgnj+Wa+wNdvXacOKLcDJEaBs1+fo4MsrlHAkT6
5flRCYNsHERkd5sihTag8Xp/f6c/vyCARKGXfswVgAufJ/uoRXjFEIMqMCZksdPlWURo4rYekr5k
JIWOCR2maldhbT5OEzWXJUJBd1fATYjKCG0x7gKCN9nCo3u7AsJYzEI07kCfnNHlplYznFlaNTvZ
ikjkSn/YZ86J6qaYxVuQf/tCsfT1/wOxDk1tmyoCIYx6SeupSJRkwNs8VUhcWahu+qV37DT25EFs
2ZrVU9ieDKaB/T33hDgkU63ZanJHe81emuAApaOmJu6YrzxrMfsZzWBYINHQHRMBG24WiYhDltxX
KK8aWJb3mEyCtf0O3+0Era4koeiNbtxxFR+rYE4nGZw2qypALfp0ajF3Bj7WtZhuCmePJYu+XkiO
GNckO0+QoHNvDAGefpCqTalPyN1YV8hNDldwVmld6DNCzhrPaozuBjMHU0JerYuO9luRsipq2Lim
FCNBgn0xrUMMxDB3iVlRDGkkHaHXOqJhI8bepJkM7WUjz99PCeZG4IprKjJbtcUqz35e0c8gOGHB
gXzvbGG91fYOEeQK1x1bj5I0D1Wi5CiIWRtjEb430hnBiMXX9xWbuTOgL1WuzhtZTylIJgyyYoi7
algdr22vvGvLkPiQJowGiVebVThjqoORqN+aVxVuzryP1zyWDk619NFdk8V2uIOK8CGuNP6adpHo
6avBMs8G/avEYohXm5U3UvzYyveXQbfAVP2zqBPVCQSfsvIfoNexFonKtglReJre0iwIVVbgC5MP
07r+MarAAe9J5SZht+CR/sd2OqYJbEopU/DxvSOj24cUm5hnqIVhgrg4bPvNMsG/IRcBGa/7NF8F
cqRG0ZS9Smu8FnXcOub+PaofQdkdLgbTIDn3RK87eRLsRvOSQ65FGfdETDls2LIo+5JPxsZqx/J9
Fli9/1fuN0YRe0vmnZDmd9q8WHzTYxWLD9w0IGWReg38omaEZPiaQV259cJyQnKgXu7t35+GRv+U
0fl80iPnpbjavcMYvkp9LWWIxlN4LKacx1WNmzeIVFSbLLZP1vVUSCjStDOlMJyhJILk3HkHmugZ
HMZqfNviT0n9KWkdGXvbPGgCCihv48IFczUKc+QRabXlL3L66scz2aIc6A9VMjjvLskzFVyu2zjT
U10fA+i3Afl9ZAJBjyokamxrmMMPq8m8b5APDUmK++rEm89jlPMTz8lhhoHhZWTWKA2D33J+eEXt
zcj9of2i/FZRjIHqBKx+aegGJgCsrEOH0gSUf1WzSfylpyaixDG8xi1GBXtxqzRCNyG5ScTUZ1oh
oCmhT9+rvxcQHurIso3VmPhzWiGFJ/iTT/eIHrhVKISf4gxJspaA3wkR8R/lkRrAJCiQig7hpXt5
REEtl+3TDJ4gpJjQi4QrtHqYZX6qK36QslA94oVg8hq99BousVudcREOmEQOPG/eQyc2uikN8qgZ
IuA/Nl7dEmOaVuLI8yaSbfdfLEf/kNJS4yTk0AvGG0RCUawVWj0ziPWRiczmBigUGaCdbp6Vgs2c
hOc87g120dxvhf5BtwXPs1ohwwdIG4d4rBpvzR2QUyuAnQopKhesc+Xg47O4Gtuoz6j4QRWXIe1J
DhA7wgeXZIWG8pWykXTtWEnloxGbpB4SdtYfe9Ssl+YHAh8xRBBpH/ua++sBppOm1kdVQ59Q0aws
MeFwbDmda6kEI3ZyacfIV8CtxXWhSll127K4pCG8x07PaKC92WzvtcBginHLRk8KAN/cIOJG5T7f
7jbYnJfQnWmaQjuWFn0r/hX4nw7WcqXYWTMWO2y/Ck/mP1/1/e1tUbRpitQOXuYnT6NRQ8eSTkae
ZPKlDuq7Rft6ecFFUgmfIjoYN4piZlHu7kBq4qpNgiFbnX5jmWnbxQdcuEeEwYvcR6zhlBWaWOXi
qusEZA7tJx1Kyj1YhLfJUfyenmNK/ZKzjuy5mpDyH9uPVvtuSYmoGSAJ9ShmAFM8ubAleVZZDBJy
VTv2uWsl9CSV+zXUTrqjZ2ZJgI9RAvHisBxX+ZG862mg2bwCe9jTV0Xs+WRYSsPETwCdaEy5/0Ef
Om0rxFNaCFpAqEjhSSRSV5z/0JL/RKmXXxZ3BoP9tpe2gDAyW3ZUaGx2zLf0K+sWp4Ju1/X2jaGs
iTMBcJYWXZxzBcwWnAsaQjGgPAYkfzYpr8H9BTUzy+zEG0Lzy3gU/Tzvcsopl03yOTVTPvCzMqCy
yFUHFnSIAIGJUGO/kUsWHUg8H6Q8WGyte3vJLNdEvXwh7GjJ2m9NTCtEQ7WIyygaAyVUnPQVkwe5
e9tS9JcAuf01L53s6X/ImrRCx4zOC8HaTvUM9YQf9ePCFMVx1trjnOiRaJh7sXa5Qq7HFtF8K66t
xMYMMavvrwTL46V7s3Z2vrcNHPslhr14aCJAQtJM7d+vJme42cw25obOl9EvSd0mBpDxjrw+Ye69
GGK5a6FaniGKIlWTdn66XDHCaPoVi7+cac+D7XksmKtSrAfLqd3nfmkl5TGWykpEP2yX85LQT/F8
lUc8Ijsa1GHvfwo2M2zN365N6DH+viLYAl95T8o5+v8DEILwWOznzHx7mTtgQ0+/MaxFzyAcQIc7
SFDYholvgAvZZRmj6BhAMBN5R0o4GfkyEAOVQzBhugBAFlES6X9DkDuld8r7OUD0oNoC9+ulXf7u
PCAuxdzxUcHFqoKUS6GJG3ZI9uK/Zyhnfwp5VDAA4vhTOtFm1d78FyruK9OIcty4vpZ/sML/p3W5
5VgddngUY4CaB0KKW8PEafDkuI8V73h3LTb+yzPQtDFstduG4asW2NIgYjALNemLtF9uadVHWXHO
FdG130ER3qj770r//4bS/FF0Yvm0nlyX9xIomr48lkqvMAHk8oYN+MgNwFIYpaoMy8Hknr/x3ZqA
r8PyIvoYIkriIWnmUybTSfUXgGmyrCvRMdsW5gbccxHdjJUeUrDPW6ZVVQWhIiCWOSynJH/cUoME
q+pkOgDUS0h5AwGCvAHC0IvNKPeDYv2gCPp5BAj/r4I77EvReZX+kpwWM5HAnKapLJ2mrAfLPmHo
fr5k5RVhD28dHmtQVk4dViWfbVJM4EXTHenuYrmJrk73H2CA1Jl7EhL/FiIHOaLQW9h12YHd/beG
nzS0Wi7UVYPNIGytiHUGjYtpmg3/1IL66x+V/BahfNBEZZ4v247d4qBvaexDSiJ4ic/YVf+hpHkH
JBxQwH+OPoSW5KSrPWFKYh3S7GR0HLeVB3XbtYh6iFRDHrPDtyU7kKC61/rLkIXk/Da5+FiuS+1+
j6aNseoBPfNKFSoqNw5UApLiaXSX9kTKlKb5uRLxFdTeYI6PJimAp7GHYo0wb0TSHR5FkJ92Ps7I
FDutXv+MQJw2opUy9IyNSU8V6Vpv7stqRIvLlaL1d7Ev+dEXiIqdc2HPOvfivJgnQmq0R0teR8ok
FeFxdRGGm/oXwGbcxUgZfuMAwtyuZFTtlGSiQiSplt7YAqIWKUPGgNP1l/jBc+Ub9bgqmJgM7k0j
wkImtj5GEON/FhWdY/JvMii4Gzaf60vPBOuRgMdM6fP7+mGdBCfsK4l+J2bS3G/Bdm+N8a6l+eKH
uOVrQPHZrwpsEFOIs8quYUS3UBeDRd1YMj5WJKC7U8dh64kxtWZabrDL45VkU6LUC8VIVORtmHeW
VdS4kEl2hTgLIMIeVgKJgyB5l3LX6lvWtZXAmUJ/By6ShZk66SW6HFUGZcazGfaISlqdehEJFhgq
g5W/2Z+PZORT9sobsjJU9Rk/WYpSwizalE/xXA+YBKDZMmRVrG7HgqLOfVDkHdHft8H0GtXWEzQs
VIV64L+mu8/uU76CAMBKpD1SoqxXpMxJXx8FybPsVnk7H9XyId2DENFEWhxIxhZnqGNR8cjev0Ht
fx0A3y8aRZlXrw0nYpPPx/npTuQa6iB1yLFEpCIkzfcZ9FSXj6Ztu6NcVZQXob/lDBhOAJPYLR7K
z9a2QxZTJQwDcvSl1hva8JEjHDIoUsxw6NyHvQcSchOISiI1p+mkheO0R8KeSWg3ET4fc7vWBj9f
GdiovTjTK6vhLI9CDAvOgn4ofU9x8LdPLlUbCbQTEzEPSszdbbtI4cFWw7aL2gszzhJFdtU9jK1e
Yr0L7MF5k3RqtIlH0DQq/iks9BdoaBx8O++iP/oejlBp5cGJ5MET8MI0DZ5neMLYaSI1CR4Jx8fM
tYXvr2KG1I6X4EXKHWsnYUxbyPLaj+cIdgFZyWLeed9REC6mdZfDXr/0eF+PEXl15iwXgbARUrCX
iq4Bg9M1dMoUDn2+Zmc+B2FBmml1Qq+/mobJwHGMYCQzNZtCbruEDeZDOoXyuvw+wPK53XrlwYh9
2twFRhaM3rpjzBmlWV2zrSZQB197R81r2aHswtTp71M4OYss+dU4GoAyZ3jP00BDEh+mbU8pqUC4
4hJKsjmv8rMzY+GoHAbxpld4+neZoMTFKBxvD61D79tJUSVaSD+iySsaxnCY1zFCEwY8xuk30w46
77HQReAGQ5okrpywo10M0NMOKKkcKpkV1cks6VrSo6mleDXz/hvoqa0F7RGu46CG3ipAcoF2Waek
/9JmW4y+gn28y8rLGF18HnZaF8drdPWWi5wURImECbA929CpMheTBTsMTJiBzEMGCidTdttBXRSF
l7ttwxhYjUsYw+SlPAzwZFs3ZBMNdi4MbUg4GYSWE+HlgnDVEthOv+ZZUeJYebgd/49Zia5KsJ2E
WI/kb0bHkwLZ5kT+xz1KmIh9s9DUjfc7h40RFGowJktD2igKH9eqSAsrlcAq0VG+4Z1PaR7e6UGy
yfAY62Cq6co/ns+a0rjrb/v2UH5i9mxROf+EtjHyD//nEgJoDYO+2dEXGpIqaWOe5a5KVxkKMkHw
mpeAD22lhO18zKGIu5fYSigabF3zNBJFBFAUJr3LhqRsAbpypVrpPJqGp68+uaRE4EYzz1NIMu35
ThvlgFRzXcJ6VdgthgrQ7/HUHycamYeaYGBr8/kEy4sPetKq4IyVXYov1q4jfs6B8ALqjI2f8+qX
5fF3q6ydz1KYSwQC/4xDAlLR9yIp4r/Vky/dsjYw4cBSaAVjYcroVvyHQNeXovcyqnt+pgFFBEdU
435qgY+NUsRj1tmtq4oW3l+0KwcvkSDLyWb0stFh0ADMEx4N9n+cXyVuuATSD61MiHpJzXMp5Aeq
++WvLAixlz6HuDiDM7s+Tvr9qNhoVXSgcWekGoMo7KEsDxw/iqiAVYFlVjQOkru5mcy36FtOKaaB
2q1Ow3kvCTkww1fRKCTV/DufWGsy1PEEvjEgtAVhJhRLLfWqmUdu1FVNJ5scCpbjo8lUoX+zFd+d
GP9XH9truMIQfu11blEOkNh3iYFMOmcVQRKLgm0zPRwfomH2zy02ajFuUkxGJu3Gk2YE37rAhnH/
90RhY9WE7AINT14xhh1iFqK2jT9ZDV7kqFq/jQYPHFZlfNyoliLpZl75kHwxTPCDWlgMkJ0ZSfTD
Q+r/Z2ROD7I57EtQqhowax4tFc5EpeIo65qxlCq7KSuk+AKmWrcqvWC0H5/xyFSKek01cLH46QPX
1IbiWnKrxSUnQSHGkclqhWoetL1/x+41Xd7qXcnG5O7rH4sf0d8bpWPnrW2aUj0lNEjvm8ohQGrQ
Fw1Vi2z4llpcBzFkBn8XmccUGfW68eK56Lak7Jmjnni81gjoDr/OWhQRFxlbmEDc1Z6y2Ine3G2n
0puIrypVacQVrZkfLdCk6AnsLM7kemQK8QxVuEkm5ZP4L35gJOBQsLk2qNqZHxKPmfTuL29H9OJu
Q1S9nnQL+PJrIaqoVeziLW4C7czo6Ch5ephrN05l6TPbK7cy4ebqW2bjDVVasHs4ximTA0LUpuln
E5G1iZAER9bSarFZYOaiq3L8NcvSO+DpZNaTQH4jFpqoVA0Mm/HN7WnH+iafwve3vEefFPf6qgwM
CIx1S+2AbcvnGRba+2ZMNYj90b8CkH0PIb81x+Wxi2cLxz/ZBnmemXuAW8ubi1i7trodIquixHcH
oajeTD/stvtcxTbupS9w2l4cg8CsPqUjtMQ73McsLFTWEuRNTjMNhumgcvDrvTNu2dW8znh82bgk
P0viC82GpAT9DbYLBjR3fK8fVMgGMjpDgMKrJ3U6ZNqzu6Uf4puR3z50Z0KnFSJEBHDANOmwru3h
QcuE0shPtqPAHFuAEoQhicJADCbyl1r8jAg5RWsqvrb42CJEygq1HNINFmQxFinh3yHeGifQFnEw
uc0bXUlzqwIphP6N/t890P+VWQm6ffHhhWVPwF1nb73btJUdu5FBbGi9MmN7xe09cdtje64XYBq1
r6supelAegxKZxjQVhRq4XvvfEeu7fTgd5jZvor7x6A21EgAPp5DBH57T8t6oJn68p4oFC5YcaNj
+2juoEGUyfj/UnT/+vdHK5SVToZ/5jQekdfwtvTH+GPL9b/AOh/SSz50PHA2ONcXd0BoxiY0ue2z
LZMxEYTsDoJJXwBQBC442zGzwNUoPfF3S/xbIA/SM8GRDjSrs49qlKGULd7Qeojka5cc5hL9Yay6
rvIfXq1f157s5JkNBVoKxGcZDQta9+fllkxiDq+hK7WAMUM8/VESr105EvW8mez7KIfUCjPO2oCe
gOG5IzS60T2y6zX/LONH+DE/7oiHoM5KFFFOGOlOHuyVe7if8KoQPA7qd0EplEg+e3QJcxSYzV/3
Jy+/GHvdXgKXOGJU7siM+spdaDOgQc91DGUqB9GHxGR0BESxa9ONvrH4N4iGtpKZRjEFy7wAfvgg
voF9DGxjKGDrUVMQEsuHAVOsbP18APLIkh80BMtXZ4hP4ooAm3WVldjx3Z2Xf/XvHQxIoKVgKOpB
1pnCnNtMjpVj1DDhLP7oMmM+DaV++iLAyGmX5dp9nsbV92H28WhPbGEh5FzbxHupdWO1wBxPBEUz
HV5Le647UhzRqNFHW4Uwy7H7NJ7D7RfrDnzUtNr6inB5FLLt46mR6Y3zGYTuRyRM5soTy4yiPGrT
6SK9iY6bZqgro5PpByuYDx6oocgRbmL8UnW8vAIUI5d+QVaYeVTA/KG8VUirXJ+1Jx9gXsvpnKOG
f/XKjunue8S0OiYsyON6ACFUfpxcF/caIBE51YA2cPTuSBiKMo4H5xLXs8evdrgz6A82vo131wcq
5En2P3faRByXnWvIrIJEGoPxbwszXCQ2tf/77dmx53AIg9yr1K7DLEmP6Tq1Ds+iiknnnk4owXqU
wZjmvAyk9WzqM2D5zB4868QI/oRIGbU4d0VyH3aLegWlb0ulHQnLxdHefukfGAdDXK8tCrDcoIgZ
FVwIrEk1FR0F7MXmwurov87z5pgEIxWCcXNz89s3VAOJiSVi5qe+5dW8LRnpyTtUAXItzs8+4Bts
fkiYAKz8+k1D2jpe+BEwhnh/Z/xYk7I/djU1tcZVmagAEezq9OnepZPc9dpQRk4KYkOzggnzlH1Y
F14jRzUme/nSZkjXFdW7a2zYoGMf7kiGwZf67ecvSwZ1AqD5rHwK9vZQYV+HL+E/YHdxSrNd5iZ8
Do4o9aCi8x1xhCgepY3AXBHxDkatV0W7toftUF1i2ZpIKZR9DyAhb2FpdzzilDroysDtNPD2GCs/
i9g+RnF6JgMzjsuxJ262LHCdG6ICrPdpOJAEbOQj1g+sBpD7eV04+GV2R2WFGz5yr8EErgJzxmp7
OL1XeP0FOvGwB1vjOkFJDxl0M1VDwIovtI0Xgel4hfCJAZrRB2xshpv8Adoaa8RdbWc/wAkNsdZX
H4dBHXltj7dK5WlDdODN38gZJy91VSNbYS/BrWK2VsAZ58weB+uerF+grlotQf6zEMO2UHj6fG79
nR6kSCUAlMocaNh4Dt+AqzRoHfD2TKtnpD4F6+R+zKDb7mT0T4nyRDI2d3CnpE2ZdqVBT4gvhOJo
eZMO/Jl6TQWtKurvs9QcYdKyMLGlAP9ouLaUyitn/YfmL3Vau2PIME7WHp3odhh7KzUVzrXOU4yj
f3TL4J90yeeNijiUJC60n2601kEWXult2SYdbvE/2tFrrL4ik+wX5ArHTGkjGLhF1G/A5GMsa9YN
E6Bo0rKlbYC6nsrFrIA18xT2hXt/Ie33i0vvwf9FkjGjyAWpHSGV3zk+Z2zAdVgrw4NYyzhoGXgd
Wltyb9e8Ty0dKzN5G7ccfPVOorjU/xA/11cwyfWGDII5tbNxvtuTzP2cLmMRJe6LI/8W1QPPjVoK
h4AVmxiESb6sT8OTUv2ZMLn7aWMbIV5tCZqIEx7BJBj6RTssPMQHD6KLOaUdyOyf++mcwByuQaLr
hv6oZi1SFkP0CDhyN5IE53IWnusHhUSHwLsKzJeYZ+FK+gf0++/77jQctEjdhcB1/Uf6+oPHy00r
03hwhfCoaOSHaJTpsLJTr8UkxBzMDJKlnkY2gsCDxxNNKidSKd2sShrWfQFs45WZWq1fFnAprBl5
dCG+uoGdBD7jeVs8hWsVEU34qltQGZci3PQNRF3NTPYvFsF3zGr+FXquIxSxikqu2ZZPKWzj4CVy
WSvBCONhJQQnmBYnkAwGk6QZ+inuVVrYM0Wi5ioRVkPxnund5Cjtp6qq4TAC2O6qp6jyeAgcTEBh
ELCH5og9StFCV0Hp3JQotyPizcXyLeUuPb9IwIVm9s4Hl9uFzVpgOvRYHMTydUbaR1Y5/aEJtEXh
RWJk0msT99w5pAwjXcjW4/qDd2VjtxTM0gMWP12Wp4jF/zrhVjUgbB7k+aTrnQuE50J2j7I/0uLq
prH3PCsSo+CKjJlvoiWfWj6PgtYqwZ9u3QLV988QpaQNG42HNZdzTk/HIexjL69ReCOvH5AZskGm
yq6lnPvjbhmHklwsIOjgSB9uEYu46tpgaOpSVunh5Fc88b0IKrPNagkwIrC7GQOCNdpHtBtd5U+h
mvhfy0eefsbdNsfG9O01KsxdqtBgtQZ7gWbzAiZ+Hr6JJwyyMNThxPU08Ac3l6NJjMjIRtfU6RbD
h3mwJK6zs9IPOc25Tj9se9Px7Ectf6e7SSkVb8s/ENdJQt6Dh32j0TX8D+BWFg7GES6JR7giCxqE
J1DKw3VGFhX5VUigTIUjjwJJnoiqsHMsyIQ6vjlqa7vNM3moGc+qRYyOvB5CU9C/HZj4za5kg2s8
FeI+JtPTcIgPEMxocVX9kHvPirkjeNfl6cytyIqIc715p0HWq+ntxwxyeL2np4GnkQTrPWmnM7SP
rze+t5Pbb7nSmYBvyeDaEfno/RIMtDW0D6mx2Q6kUqul07Z1jWEGwlpI4oB5ykPzrotr/2QHpjaG
XoPiRF27lVUiN39rtylL3PIlaQrFg3y+utvo1EjR9mGy7YppsgrEnseMuBaQ+T0TubPh4WkdXLBY
iXON1EcmyA2SegzPkOXea/6LcF15kH1kBzQy234Pi3eqeQR9VnXpATbiPHAirqGC458AqkSrDgSM
I1WPSc4B79oBwKYukucs87WsD5Z9HbYdhVzL2ygioGpHF6+uY7n/8AmdTjX5om5BAXZjJAO045wt
/5A+xnpMSA9+oEOtjGySoddTlYPKLZakiD26XCxQmDg504wk+qDglVCiwttjgafb9hBe1jZtJFMf
Z8h0gOxvmE3aey9l00tDbCjvtUV+dYNWR4beDdCgnk6ife01tDhkXlNAKs5K1CspAnD47iLA9w2F
vQAQ5/pVnSOCLuuwzgJa5YZTftZxxgas1EwRZGlel9CyKMVTuv/C6ruHC2tFGYWGM0clCGb3zAEJ
9L2XTU6LLeBWTL1nOX3uOJlAs9a8xAYwIZG9ORE9hBxDwvtOyqCZZw8jTI6hsOgty50qFEpxFjcU
CwgASGolrbbs5Y3+1Sqx7mZt50Hv+Fdqy40PbE/chzpx+16mebKy0AvicMhhLwVDAsC/LOen3vvG
JtD89pfVOYQZ7suoPRI2uV4KkVOt2HvKF2b50Y6JZtofFVeVyAFb7xdU9O0XGRJ7F3kvfbFYktQf
xjfTxCQ2vFAAsFk6Zh0ifC/jJWxIg9L1v/NkvggKP77VCKCrvJXc5Yo9wuoubnl//mGnxXrFwVTp
GwXJyA6koO9NdQ0KAXhEu6Yek/e9cCt+9FOJ0g5B8+l7bMsHpEVq2TyvJKXJgumqVRTaKBXHElR4
dkvFGsLJFgv81UcO1u6MFCPj4krujbz2F4lo9LIa+ZIdyClUaTsFgk5gV4QxdZElK+cs6ATZsUr7
JOwPaTk9iwyAao7tJeciQo0eNhcmHjtFvL267w0/Oyw84lJELj9nJvM5ncfRyTDvnNZZStcolkrS
FHSKIHiN3yYgvWJb0S3Ejv+YQZxORxP8+JxQESigfUxbzRsby679q/xufbDN5woYNCbfn1sPMNfY
57ix7wDIseqoIBaZNRB3E2SCPglzsAxBv9E+TcDpOSbm9Sgr2jolEgBcHdyPkaoXCy0LwYg74kqu
7tGXlfmh1iQJB2mVS9uf8DxfAjBpUYhf6THflq05fZLvHPetC7Cy/BoNMSJsbavcfZKBB2LKIRz0
YoHluG+JzfRYTrh1kKUd4nqVZ9QxV1YcC110jvcqOmqr35zd2bbQW709A5xBQngxl4NilFdUInt/
4pWiN/w2x1Z98ZXJO9L0QjIlVpuYcS7qPEJFgZCmuIalC7oXVtPhIeOjbr2ZxTuUFwWuNXswu9YS
96p/4/6r156jSfXnHwsFlkt0QbzX0qYtrkgnWDvjgFdUEi6UaB2UwR4sPkyzbzZbU1cilX9XEJTy
xk8xkaIcu43LM9++3nrozu5I8FJB3Ja9vWTYBbc7AUTNC1cQFF3vrKN4Cvp+JojkZ8VgXGVkIp5d
bpmlID0Xucy9prQupTtT6zR0n15ovLJ7yuxeUbAH+1nWKB347OmQjkYtJWysJlSE8iMQYt5FUNzf
YQWbz7+XSUYmTGmhh7kaD2A/80gXynCgsnTqO44hQVFl2+sFmGYe5wqolKk+BWUj515msaYj+V4D
8ycAOAJYDZljP3d0qYiQX2VCfkDdZToyp8WM9zZpqtdW3iwLF3pPolpg5QqSjXm1f+vT1hO5ctaP
G7sKs1dknxL+ZpA1WhKbaxFZq4CsAyfgDRAR5GM/AJRPn84YpM+J0VKLlu7xOcTJZGBNIGQ2VFlu
oRdoflmTG/yVxU2V+4UE5J5/cWvU4+f8ZRQtr/YmjHTYRpg8xYD6ouMNKGhTrAJCXDpx4Zc4qmYQ
+uYPB3GUQFQIZf+h1HEN73BJVf9oWg1P/MpwGB3kv2e+Nsjk+/co77tzvANptKpBm2sR/kaQ/2Xf
6PTasjuWFo7/Gab47ZDOEAtUez07OhPpQYwJLDWQwVzq1R3bZcxIUaI7228sZyfc0iRzkV0YHUGg
RvtXIAFlEtrjPRMCSK1fy6YqH5RyS/5LxARJzKZoLwM2kiOJywXet9gSoL+6oUGvXqF4pfZNbJul
t5qUWMDIo30M0DWR6IeMWM97dZTEFvj1qO9kwQvUffA6aMymr7WJHrskrdn3045UljA8/wTL9Fvu
OhEmfulj7LZpcbFAQwAAasU06XWry4Ewk9PoqAVJwiAD77O2GwL8/he8u/RoWHxgq3WD3LCE1t5S
jRBlCrOu8RLSTRtK+t1fCSQEHMmKzobDNbgOezIjMUqsvPDDlLpVc5HpR4UL4bhFMo3a3s53K361
U8Ce8rdKpycKsTKIOxykci2UH9WxDM1HowgvQZlQOW3dPG8XWeyv6K880iwX/DJtGTxCoUhxZh3v
sGORt7cNAzUbpccdjr5wJzLvNdDd1qFKlELZdvDF4jTIquSNTwGbosR5qVaOaiLEgk+2/9QUEY66
pmzEYPjinReKPgfVqeCDZWqQ4dVH4MUiqym5wlhA4Yz/d2ZH1l72M2tm5g9Rwwl2VO+Z9hc/4Hj5
Nb5Y+fwcK/ATqcBpZbgNPLgqUcY1e0jeeAOGxG+bvtddPB4AeYwdHs2vfyvzx5Rjj8zsTx9k5s4U
ZG7ftSZ1xw169w9yPzpLz3WZP/c1ZyW+7s4bm8fGmUjyixon3RqSQIn3juR1OOGmUPUjZjA/iQYF
U1d4OiE9BUcfOWwe/ZB+JaJUecs4+ZDhbUmUiqD0lW3a+ZLCfmU3TTrUJdE73WmEnSRallDFwilU
YSiUYeExCJw530AiOupAtIQ6fOfW2qLGpeyqP94OYs0nZ2VyeNtI3HdZiVnjp1l1A/d/oEgz0yFx
WfX9K1U02tyVCH6nHpfe09zyS47neMx9E5xsygwpse7c4sP6YrFyw679gtnI5B0dFhSnq/w+ga1k
xA88KjjImW8phKl7VuRJfs1iqq31tj/lXnHe7LUgRZ0NKz3x7F9XrqONsXAaCHuD+wcZsPAQ+6DX
8024z06Bm6N+/xeAkl5nOsHmbOjfm3giDiXWGUi2aVNoPhXlvRwE/dh2pRvsi0DnY8RKJDH4XUlk
tO8cT6IfPL+OyU1uycJMcWt4cW0Tq+GaYmnzRrbrd2Q8KF2D6OtS/QkXxb5f3MfaTl5dSd/lS1Jo
kAvNhXQshVjq3GPbRh8e0oYuHDD09nCq655F1pkd2QGVQEhCyEARSRiADIGj6t/EP2tlMm36IGE4
J5b4ZhrLSgJhg0IBIvg/+hRkskK6y70eQ/NYKN6t6Y07NOhEEPV7AyJIPvvMIPjylULO2sJZiEsU
eeyzeHu47GICWN0U/f/DJkFy1vGQleeXPxdNnKFtdc26U3YFiP5OQlCWC5ArsuUFnIhV60XY1KrJ
d8n1Hhmw5RKA/3RtlQdNfAeqoK3VP7iMn/7I+37tBktgmbZrZDBarU1zJhLByZIhl8bO50O5cNQK
NjfIydUjyTxuWlr5a+MpJ//4V/BxtbsjCuPaaVWK7Bo+wDUjToajnCmyZg4fyhRePds3YfUCw89i
hBmwlHiQ7X+6CIv41h1lhAsLbFeXPrCiPmp5KvC/Dng8YPTSkceuwNd0zjkWbtTcT05KoObJozGN
thMpyIcZi+NBxEo+h1lbNWLqQUnxijRFeiMluVXKVm4InfhkKRvEn68EGu41RHEKyDvebd1YCuGd
Kv1hFqT9Bb8AN32GeLBdkUpR3jya8oPNXw45Lj1F0JMs7HuKMQbBQdYLtTz7WQ+G88BjJh+m7xm1
Xm0fSC/5gMe5sSWLKcpQAHN6OTWIrKP8Xj2LSzfMwCmIySXY00pGGTYjgfudr/T67FtUyo4wk2Wo
b7Dg7BMDlnrNUGr/Kd48Xd3ADX38jRK7fyqDK9wCMGw+pXMtS/LJVYUsKh4lbeVumKuodKiDLzV+
FAGH49I/cwoYBafPX8YDS/p6WPMAYMa3fcMsU5Lk81HHl6Yc0VulUSgbVvOw8/7MIvfmA8yDc2w0
DiYS53kYIev4AgfldbbbYQaWxeQl21lvtVBBihuwiU6sXF6idecfbw648dy38r8LcdSzBFhGzviQ
hsb9Mjj5ScszXlokKFyaFZY5MgDJ5JLg+VNJWX+Q8/XsNCcQHb+FB3SmxxVU0E8qqFG17aBkmzU0
resXdJgN9wLxn4anyZOaIv23fuVpqDAsd/Xk5L5o7pVlWDtACRt/Pv3pq4iHs7bLu/dCtBCVEAs8
ZjdG+1SoVxB9eyUqyTjj6ps5iDzu8028dG+6B68m+URZ7wgd9MKZSJApTV0PkKfapzS+5j4U0gVj
JtVHt4cSTuX36RGyQ4f5OlbBNbKDtP18Sp3xAHYWtr1noE2afGe1aMG/3Xg1yv5dZYbDDrtbDxiL
mj8f7jU8lluPzG0NqVIlcMy2vwOR5mCP6vywOX5Pdb7OqhBvYhqV7+6vaDCEsvC7Eqd4r050NjaE
JFmSp/bgJErxdF2RILZ9Abshm/65CuMItoQQydfEHioyEahRlN5JsWzD1UCNtNU/dzLlaMNy1KOA
n0qkYeP1j+4Bu0l/utEBqJygZahkoDpBWDX4mHTMzFmXSGeM5xG2ql9HQ3klS8oAIpmhuSLoO7I2
22eVV+P3TcRtVPmoqmxIiNEuKFqjdMTGMA5v4qMKqCsluuw+wmB7u2vxX+FTV5wDV2QnyiY6Be/a
lOd3s9iuJOMfZe/iPsDbDkba+x+YwRN/zQXB9bLysooOKnurCUTDPJRr2IO9L/ikfn0ONvKrpe9E
yaD74WMN8OyJL0encun0/xAiXKsiwERN6XazKHLBafHTl3/+UTOy6c4ZxfcpVPEcUoh/NNWAWmWi
IhRxJFdzjtBig182vWiKHOgEXgX7slprns5J3ggscGZMbj57G74Fkfu/M+6EFZb5L6NnJnFa/Zug
ra2nnDk/eq+Sp6u7HcP8e6llTQMzSkBar93GHjryDH7pJDFuMNxacye9Zwcjv53vXO6i8szHYg5w
c9ibZUk67vRFXyujCRQ9bx5fmRFnerLylUNdc8N2mrghFGFfZ1MhCNuvTpyGDLgA6iXwZEPm1UmL
g5bQUYhdxjniqwyV1O3lYlEXt1y4U+Soqzs6DqKoWS58FawReNj4ooigXvhKYDDQj86EJXDXwmQi
TCHKEeZUeDsoe8z1hRAXIdg3B8JJPdmBOWamakYi13x6Jy2fKCSstqlWGddtnOnSZkl19KOu2GnY
BpPYvOKZPULQe9fI4XSg8+DF+GvKMtHr1jJlseFr9wfAYl72YxsosB4nEJtkF6PqXYh/I1zmEWX6
EeFcYbmAfVb9K6nERzFe1hbKI8D5AwpovpO5c8eDwU7ZpU6w9PHZSMRiHdqJ1rWXfyTaXtoqSBel
ACHel0LDUnBmP6idmAdtqMO/JDWTrsVN1AbQnQVmY9j8OPV7jqzp42/jvWdWL/UQdcdQRhLbCdVn
tjAN8fYTC6eEGeVM0yq1SfxlUX/jpDi/Qf37cQ03ZvN1IXPagQ3tTbjjWxwvhMTpaQYxEUQ8zzMq
Su7A77iafJlA2ng/LW2odwAp9wIABG1xZOdZHpIOvSMP/UJCe1LJy0pbvAt3PfP6mDFzjDn49hsu
jDe18YKkXJEgJCDJmmVNIf8+re7MhBH5J1Bx2a4xGTn07HI6GRE8mvnnoc2jFPPYEZQQxClrwwkC
Ws2yIaTfTnK/BXkWKIqh2cefzvzZ9pdt21ekwdOgacyJjsjBHgIoovPilTd21fgwXMpxXpNtUWeC
u7TbpD/Isw5rP6v6H+SCk2ID9YloHOxSgcFVJstq/qRtjFmJGJ37FT88ZC9pbPmYzFmW+zEo+354
5/3Hrq3wVUymJ9k2dxzR/C2POnJa/WZktYPgtcji7WIgwm5LwsPzqf2fk+yOlk1QzmUSn1R3imZq
8thrzAHIHK6J/3gob46rTpaEr/1SwScQrgl16FvFuDx/LSX/+UJrF/0JQWuBjRfhPO4deXXmFWno
NiceJyPO44yP59D/CqntNed06p9JM3VX1wZ6HGNkP9U1CwnDOBQ0JNAhwP37UZaKU9H2pf5/A1IA
a5Wwa2SE4LUuug3qy5Lwe2oKeSQh3GC7rE/TpAw9J4md6rqYjw40a8yrEXkQUnuaSRMu/S2Kfn5d
omMjhpQQsdr8M0jmvEks7kt2gvYg4fk0IHB8CpRSPgOvc7TjkW6xiJjRbLaGJ7O69nTXDfaTLbMn
ck1s5PIng4c+4jZej8zfO+vpoTJt3mHNtSGDrPjyB0KJhPrxbpPOFB2pNp4qQjfXXSajZkiwx8wv
pIn1tUt4Cjxmm148jTjKC0ICuYbrIaOMHg3j9tIN9qEUN8U1hodXQ29OqM0C3KTeqz6UNDo4ga6D
ubK3/9W7ucuxwgCCVHj8QwT5EHNf1dtkxEOrOYlHEd9t7yKZDf523RwSR45/9sfwMs1hPLAv5KLU
iL/2eABOKSIrcMWrMbCPxuNQ1+wh5NC5Bh/4WKE/f35Yj9d7YyTOETOxDKsRNA5iofAlJKMrtRPF
zfurEeDWsWR3iUDFqzBLjn09FnJX5irCx1b291fNTHAoS5oCyuN7MG0ANmRcKXU5PSxwSTwmWuJx
ECVb/r8QHLxw4kzmY4EecPvI6msdxcyt02WJMGB3+N2gsjB+6ogwn4Rpxgvy9LCv3ivh36sZUaC+
stSH6FhHkWU5wt6231WATsUndkeSrIhu6n/elYg3jz5vMtMhaoKMYGWArSCdkViuN1XTWsV6Oinu
+IXQMGoohB2lUUTP4mvEDG3at7Z/bXsIVJ+zSV05NhHOl1ONz18weQqC4O2St1TroEejpduA/oO7
oAFWP38DuN3/Fld39iA2NX/zRkTE2l1i9NU4O1w14g7dMnIKzTfNggFVpkPHEOmXcbQJktpv19vR
qEe6rPAtXkaM2ciCsx7U2pGoP0sA+W3pihnJDKhPbFcswSXh29lrmwwAWCRnDNUQhtx0N+i52YbJ
e1N5R/t3R+psVIu1Kxv+3ZFpE/NTCVhlWM21S67Fubvrlu4tZf9LofCfIuqy7ipTRnJilTZ5qgli
t+kemQuabpoqe3a984M1neZIcbTlv1OtfZdrjHzLVtbY9bHQsqkpOAC514Bg5MOHi6E6P6Tzl73E
tSQuREbyjmqFGFKkzFhv6b7rQQINxjcnxERMeH9dJIEYoLmO15Vlrp22g1RJPDVBhkMgY0lv3c5m
APXweig2zSaRyGQyXYyUTxabBAxtLA22liB/qimPU7MoWEIGNWSnDWswVEt4Z6EvCTQrl4Ebk97K
hMx+qG5FyfmQeax8eh7FpNiaoWZ4FrQeTOy0dAIxcVWnMeIsAQMHn7L0gaQa3Sz/FhQy6fHffP8c
FPCid35xxDWrcJycxWYbKNHSyfr6n3VMhmeZXEMmV2z+b1IJjQOZqhkiZ9EjWeW7Nou1nvdD0Vtm
4LH9mBtQkZ4JtIGqZDXfxvv8QnzI4E58CujuBvZk/EYbehXNIjbHis/nxsyU3VbQTE++F/jVQdzI
I4wMvec8QfeowU1DHdy4Lo7w9VsUqIeg4ER0BnpDPwbm7I3cZcNxEpHXnFTkWZuON4njQ4nCXF5V
zvelieYaPJn5OLz+8xV7Osmzsz4onlx9AfGlIwpN+0PL7B4+vWt4mD4LQa0u6jWOjwxz67CxtWMw
hgvIMZ/74X8hpzPQ3VeLS3Wy2WoCoj9T0iWX1tydObBhNNRAFiz3fyv+2gBLD5v1dBedp78yrkCE
a1PLvi+111sTJkYWb1r2EEzHlW2Rqb+vCZ9gb4x8UNXURJpXuhOZIdNImpSnFJ5auIDg2U5RH5VA
xIhybUki222xiJCgYZ+XluyrRu9csbJkIzZHrD6V/k5nCVw9g7qYWY+CU8aN98/lrFUvEbL8r8QW
pSBSaX3MPyimL30jCzCWSv4KHgrBlx1fgS5uNe/iCiwOvONiDffmn16U6TGcNFKHXitVSsW2eWXq
UTSZi5Fkfzb3MqmJauyEBeviiR5VPK4WaMcWs+fHvOE9y3NW2ku8AfMk0m43clRZbsooxySBCp+N
K4ajThZTKuc7K1jDj8i4yzZ03z9etod8Ne5y6aHHOCLBqOj5n4GLtYxLYFjrVmgpfT9bNdkDI0KL
qUI2Bc25kXT8NR5QptKc5+EMOmm2A1orWCT13Ke/wrPh6QjS4byfEIaiho8n3soEKR0RKieNLvyF
eUg2BQyz7iJ/c0TTnCuwmM4KeLVAvpXMLRjX7PyA9mvJKei1T6xBU8MzpbZOHR0JLvhCeaBq7wvl
BEBCVv53YmzUGMvOCwOaUOPkIabBBQ5zDQDLWnJZ8/3znkfrVKeLK1ySX2c3YREkuJOrgSt9whBh
Ds1cD8ufbML/nNZRuzolHWXastt6lZZqdQj8nj9V/ipy1o5YzbRPgYqLSyA+2GAWuCrxuu6DAgwZ
srfUKF7Nbh7RMqbnZSDUAANTCq4RcCe40DW40YIXutFy0sK8aWoiMm/vypYVtJV91XQSIoIvMuSt
jYYwlXK8ikRcFMZLQnZt1QBJxUFzRKCB8ETnGBLBX+8FGZIuwiyyJpXfyvPc2ujsUqWmkkxtAOX7
hQ8DJRupixujxSXHjmYgGNMKZ+AVvP2NgAjQ70ItuAIC+HJu8gBpsOwmUfp6ajAMKa8A/9YB47jc
za9t8ACLxFFLhijl4x0kn875s+G3/tt/VBlFrsOXb/O3uowhhsKg1PLL6KY6WPFm4lI2Z5HNJ5KD
vsz9ORj1dnPTir6pAsfRI7n01Jyi2ARCI5nM7uzSMZvNF5rOYyXAsvLq22SyucC/5TjHyhTT63Nk
yNlyoqXYN86uFeFbjlmiSMpW86g5nsPZVTcxYzBVVrYRBEdIHHeu5GwbepskyxBuKlfMrDF++O1G
yYUsWX6RavjWaoILkcGrpc6AauVo+uSh5E4Rm8B07JL7kJsSMGzP0KBdN0dpAMskmPSLji9A+4sZ
+CCXcIvo4fjMzfOf57w8zrZ46GYIEy5VanXcxiOUzvKhOqHAgPjOMXE07ki9FYS7Mg2MkVXH2o7N
FIg0csxa8yVKce4EWzkQ07uSL18VBKEFcXVv4+k9muOr9EWr8paKEd8eaT4TCG7JsemZBNihHzvk
31mMWi8vh9iSnw+8BRKkOjAxlcCjzdzsB/uIU1OtFCboZ0FCtWK9sS7T+RdAdgwNW0GJi6Acth14
gOCADF1jeSBSewW086zsZL59jKrxRE3549pMJjFtxryzgfFgA+3JwRdE8/OTZOsWz/Gp/elm+SOU
XdtZ39mSAvT5Uv9EQIJwyiU/EUXkqBDrn/r8TYn3zzp0QVaz0IvocV4n2Gk/b8KBLCVkXjD3BFLY
ZzSPyZbZVzgQI0qr+T8nt7o8ZcE0PcrJfD1/RkQX5XtSgMUMPE5SEgh1D7Xlh0kD7CQn9S7OAREv
KRzOe99rMHXqJSKusr+wN++FoPQlQJatT99P/iqEmhe1YxF8tilsQL5vWNTYaBzdeeszUIKh9vRJ
sIYIzc/L/6ZmGVWOPhNqIkc0xsaLZgfQDLJctBnXZeEdYYp9XtuQo+3GqYO+eXZNO2B9S9+RfG5q
0tXZFfY7PGi0w6hYpAe6pMp3CNLLzvZtaSlf+FWs6fd3YXP+P8VaM4iR5OzKNviYgRTQGi25i1Od
WVMN5gtmdag3Ti2LQPPaRUetKRISSlhmYA+0Z690oJzKcqo8r8pYIYBnFAzo5NtwSrcjmY5K53UO
UaN7BzojF/LyeuKANhFVFqel9ezq1JPAAaeeVD4tSBsj2b5Ipd8OyW4Ogjk2+6tQILG7xFTGgkJL
vbRPMefvuu51HW9pH7Dt94frsYa8q0c1L+pQIJfoi3d5xaoaR4RCxSQVzrBKwsYClYfDsyFRlxKJ
Bp+zfoPDd1hw8J9q2v+SJcuv8Y/HBeu4dRB/x/uUI1RanQ9j7EF42x6sTlMLhuzGq0Sl0lZL+kZu
RVEfd1WLyjVKibKi/CvOgqXd35pNcftamD18LWyEMOLDRKF7NdqrdQpGE+EuWuBPI5TAE0wJSI0z
7NtKuAi6KwEnegKRX/CB8WRoSPHiAxtHknkh3I6jXaAhgzEyEKYoJWpDZOsnPxf+0654IVj2eLhM
N+zzp9Y95+7roLBNesE5agH7e9XWusJwe70VeOmF6B51lEFv+5o/rL1JP3UrzvzglvJilbfguAMy
YMAOl9DixEhzYFxzdObvdRGGudAkNZYXpSEQDOdiXRjU51hw2QM+rrauCvJUIOXZmBLqTm9LecPx
KJv4ULmTHFKNMSMiU/RAU6cOa0RfBIEIvEa7+Q36yGb8qCUF28D8dq9bTnEEMUDHY6nGD6vTIkVO
gOmK9vXaFMGuLYODHfVONWzL9UPw6RIe0j2GJ0rLC/xSaCAxmQ+erb7WbA2D3P5exOFXoNS9kuwr
NDCglYPR7Ybgtsn4Rjyd3QQTxMHj6Jp5DjJqfD79FXQ3RDOny/Muf3wGl7bmHTJT4yb9f4AurpaR
V8fwQEnzRJTTa0f10MtHF/xlr4MIEeStw48RTgMtfNwP//i5isrDIpzyf7iqYGVnrYqOtb2PENi0
z0UUVITqCY4F+chM4OzNqjoYlQPdor4o0dZHe8K6Cjs7vczJiXTtc7sMqr7JWo0IfaAHDJS81S2B
OqkNXonOtSebEPCjqFkFN6Pe3glHBwlwrItklgBya0XzsBvGNIdKP9cpGhG169Z6aZs2KF+Hrbrv
+T1uZigcYEGud7JmcseMkPp+Q2+nLVknByfviJ1xFwDr5sKfg2YqXtAhAcGS17h1PR40auNth4UR
1+6P+p/o2si1V6f5LwUpwGKlwvR+RYEOXF2j0ZVSTUhp79yDCNzTT4SF7IdNYLJlu29Ro7BUVIY7
USNOiDfYC7AocdznbNlnw9Cw8eAcm2PurRdftzrjoqpm9sr7Te80u0SE37ks8Er+1Oo5xdpSF8DD
KfiqlWS3a4ZN+Wim/sDotbtxn8PgnqHpcVBsYLm6mk+fN2Ure8y9kgZ58+AuGKyoYzfcZ2ckmjH2
0LotqzDWtbpRfe1Riwk+oFWan0vwi1malKKsRXnPOJmXA8tjOU+bZ0WeDMkcXH1DZ3ler2pUBrWo
r/0RP+ld6oUawCJQMYcXjGYPhlmBcrDqnX5jMEi0sEjR1eIR1pWuUNyx0oPOOJyFBjbM1O8eBRaX
zl3SoIWHxurFCkU8cw8KexjQIwWarv5Sx4Qhjz+Wxx1l55GDLrMbKlrTdoDKSOpsM1/zlrviJ8Pf
6t/KUhMm7Km3+jULtR+zu2DXkxrgYOM+gAsG7mZKcyJaWEA33+JaO2/55pwENNBnnfDKBsPOi+Tm
f+pMrLqed6mdd+1y53z8RT0kUfmyFvZxLYHgl86BZi8Ct31p2Iw8Nivq4/9LC2dQL0eHoY6s+yaZ
QgVbUQaCAGDJF11HpyvdNNJI1pS2/X6i98a1cAyXycCSXWI7dcKDHpoBJEU7PLz4Le4VUtipKMuK
pvn1byqJM3uoZnT1EMBBFnD0mHvCVRcHh5vB7KGJuJEXwxIXcFzpwzk2FtLnrXXSS9D9Sn2t4dWo
HyrU68diSGVHwLn4B7rzePgVXqNweab2F+XvjmpF3zQAKQhfC0B6SHCBDPbp8TWVW1sKPH0Cevr1
1nusr/ABCHZpcG9nkfiC7+B/ox73dpMYFoIQle+LIOz+DW9oxqsgSxelxPh79rj6aX6PnPpGcNou
ofj9Qs7wCrlOKxV91xnNYqrSWbYr37NdPnJ6F8ayFOjTVuZnOIaKI4gDLryUgoIdQ9Ud0WdpM4RS
iYhK2vWkErvPVSzK3HzzRaFlyIRy+unm72lv43eZoNT7TczCk+YkxKLorspRQMZ8nhYHAdAQjx6W
6JceFXJId22PzMYOsHyg34Xsw81xI3kcP4cA7g7ZWmbFnSapEyR7OPW1fEq3YICJpbNJ8uAmgVaN
b5mtf1KwqOJmX7y/dJH/bj1q89NPLCUwYeqgseeBj3hvkgXETJbecoqWY6Fkdxj/myroq1FjoqI0
Pav+s32HjMV29vYbaua1agd1xeuToqi07ptB3OWfzwF72V5KRaUxM6vDjlb5RaTT6VtQ8q1i86Sl
wdoKDxoIwZcrhpY6ep8a7tIMFtS7K6qqiSRfBD6k3df7YKNJ5sMB0xerso6O2dpk4t7wgUMUyUrT
00Ydd6wFywd/Z6auqytJrPnNaGt7cLIi82dTcAnvVwg4qfKwuYvRZWYqj2aJjYX3f+L9QKtLPxnE
o6K6nMoINsucEZEk/B/wwj2/Hv9UjTVK3YWF10O9FMmARom0Kle1kUiAridCmzdnHmS5JYNsXFhd
dIMGPomyJr42Nv5SRaHyOYOTixdjarQbF9I5fedtVd5KBysM29eswADQMWvZelckhhmZe0Ybeu9b
08va3IXm9ymZBwe+Ht40dAs6Px/ScXzY+2ndKzs9KKJXrE0ICGPFpS+bb9E8j9cabPo/yR+VIB31
Z5qzlSvkPNi/PfhtxQcz63xDBedczjPe2g/iJrV/u9qCnWi3TMWpTPyYc8HZxutLk1jOFxGU5Egg
wPC7jwXOxO0ciOk8tX6IzUCUjuD1kSdfxLl4gNmOUajeYWWy9Ihn5d+sOYh0TNVERbRFv4NjJG9z
BKps5wUK8nDHvTZHmkCbyGdgSkKj7PuKRhkERdz6/oFw+lUsVjz3mlifL3NVpJ/R9SomwOh4D/Wd
cPWuhNYL18LeoGL3QAV6VOOycJ6zlFgWf0TjiR6y+tzRjmdZQrsSRGhv8MTszJ27IS6nQCvQ2F0I
gNuj1aM89EHJIGYcj0Q2aaZ3FxKQTu3lBvcQjPvtlMK5yyXbeCD1VjCUww0dYelylbc87KHuhsgr
6VoYqIyhk+xqgTtAHMyTwWpiy91mFBImStTR3z8QX8KCKVxniT6fr9YpX5y5hXCVk3RhuI/h7WmP
cRcE5HWEzZufBN5wVkyGpjGophbTCrqF0sVoaMmFDQv0yVV8ZwPgAia7EohTzryERXX5D7u6wAOd
DXDO7RlckUHzNzhyaewDaaxeDOhSQYI0Pp0Zi55sO8vu3takaWrhD5nsWU0y//ZFNukAPMTdVHAD
vSKDbBHrbycxSMgWq6lY2rFEegP8yaRBczUerS0xfxrLUBtk8fzlLLhZaAJFu41nUfoTHMFiOlhH
RwN8r/O8Ubul+zMXd6Vnko08z2n+i0mYU36RkaEPL6WC1yrAIZrkCjVQKkt/GwfFhb10EETvxczg
xD4aop879nW3blIYz20h10vHhacPt4ojYtEHk9n0Ti2K2AHxiVPVUhtOnnqMhWqOzIeS4AAhMgGX
fcnFokqEj+fJtwcXBIi5aVbKSZGXLuXaXUTeg6F5C/xsHL8VR5+TFWpb81YvUJyN8zwoXXxi/baF
8wzeeiQANO03nSvP5sgPrjz58Z1lSruTDdQGpXjnO5JrLEgY0f1/wap5fRq1hpmqTQhDmH1QdZkv
HRKWqEFXKSbrsmIbTWeVRZrEN53XPJprudFMZ41ca2sqxFFHzjEuQa7/hVS6WCsbkJZogVFq/7Ul
pAGe3cXYOWNhrWl2Ew3eCBEW2ftoeWiQEJcqyxwkpu3xhWYqBQSlz4thXiKMAh8xTmJH6gzXbJ1p
m7zLtzJwIUYEYVzIQAeId3cAkAWXpOci0Gi6DcoDJzZyLrwkzmo0yw5NQ8XXz2kwKVWhE3/dohKJ
2WZviupxo5dKkb84Eijjr01egOFZjR/xdIFlDlNRPRqcvxfINhdbxKn2KX4z8KhnIoBoNn/p4sWB
g5qAF8vi6Ko7aqnBmPA1Zff3ju8x6hqr7qPsRLZEBfkgDOvbIyzzERYe9l5HAQhLetv7pQSno0e1
ao7BRKciEYDaureBQ6nWNPJSggVdqsPI6K2x9ceo+jUYP2qOGdY8Hf+O454jwmVr2scgxMi07yWW
JZ8YoPYFjMku9F49GtohSWWv7SC11+ZraEEuqDNMqSePVm4re92VzQncPkSi8jOw2QElWXzmY5Gr
/rvtWctF5d0ORzVThNCzlv+xmndDehQT3QBI2uHXYSQaugUq8PrEPsN8JtZoI06XY5quCjj89AO7
HZNRKRIx7L6zDjnVxFkbtzJoJRpOsZ7qHu+QX8+h5zOsc/UhYUX1bfImJI2pBbRtmZb5HnTW4XtC
jIpK7gTE/KS0h/FWsnbcilHbcKFHYENpNtBNafObSYpv9EWPend+o2KUc9ETKphHerURotpNqr6d
tEn/x3qFo6wWuPe89LcaaauKY83Vd2LAh9m4Arnb37vOMnfg+1zFdse7XtYwXToc+PgDfHngF6/v
BfvfoL6ba6Hct0+fze33E7Vao/27CwbNWPfsKw+ROcsgQeam/O6R7RzQyrH82P1m2JmytloAQ4Mz
0je7Quq2qjROhbmTyGW0bCmSkCdpV1HR31QbJmYcz42p5bQdZrE2vD0r1hp5ysGO6EwsLXdyLPP3
om2wKeuqGzIlb1Ql1AlUCRb0UnI5iWg2OEMZQQ0kF8oOsZl67xfZUp8N88FOAtrfK94/1C0B0rsA
jIXz52hQtgO8JjUTgF6u6sCxpAJqRedc76oIs08IhTLoG33zGLQLMep58A71+sko0ncItVUCIqnq
k0ivwTIxsJayarJHbkpCvDG7rIqcAVqaOHDjp8HP5eCQuQtCm+TX2E6KwPFrn8YM04HJ5KbuXaM7
f93VSTjORvSLblVSZ6hYIOQPmEH3/9D+Erh4SosnDkhp3/Z28jKVapLVoA8o65+s8Cbq4qIRtW3/
fgQbgX9E21Ii1HQ5AXWXXX87sYwc2TJgdHQtBT+FvWYd6bA9wmEfeqUYmKvfv3eDovmluUFPiQqh
tyrFWNzvp7A44zjAgV5xIqQMkRDWxpDT8otcMtfMj1/eha+5Sn4bWZ+EgCjqqG56sA82EWJp64JT
eNAIRC/1q8feoTmSwUdnXThMhSX29gXUYnjYOt1vWExyG8HSMiBGGkqUMwmc3JAaD5OUXn636yxn
/7+K9tfsbvvoLpJ7poQL2o8Amr785yHauycKpSfhsjH6y2vFhqfP7KJFrdsizPI8A1H8qRTpzzmd
M1L+3+oH8KdhbO3ziKbeJaubXkiyXJ8/H6DhbjNtMgrFNTLNhnUIXCYoItVjEu/juEAgpC1ab4wa
dIIH9mCHE1Utfb+LDecXUcCke5ba36eiksThutMFhAUZLu9do3VeAJ9SRoA9wb1vV9JCPBswolQe
MjD8mEvqANKF7bC7vRSyn/8Qnu2Mun2FdmKtQzwC1Bfhiq967zcSPWXNU8Cq8KR48c0Y1VEp4YaV
VP7JVrxFrQ3LXFOjDoa5wRJXvtOQcj16ryNhkrfkmYRMdPkf5i1dVGYm97VsB/QLsP33Ja0CZtiG
fEzrll5dyZ37qlEQ8uhA1lBoRjfDNCguvMjFFZ8DbbAITZ1ofDJXQfH+AYxWXHpB25QxuzA0gKqn
HlQDiRJogULdB5Da2OgV0+9gq+R1Q6A24g7shmGhN8BxexxJ+ddBvgRiH38Q7XK+1vTsWPlNORhy
cv1S6LKtsuheackK0n8i+mwao4o1zuquLm/bDiaiAEVi0ma/MFC5gaQUO0iY3BXV729UaqSNSYTz
UIEZw+WGNXPIHXEViQG6vWEsiRRswSXVMMOIGHCF8Gat9/pj+7WCFiL6d+eIuM+J3DKYzWxnonEV
Cs6YmP3UNTpqD2gwp/teeMkEEKCcmtGWFY0zIomMRDdqADzqcQzHTwGtBgPTYYcdTSt44wMJKbdJ
lHTR+U+6ddFEfeAkCegHNUjkRfYktPd5aHqoHKZRUv8hYaRsmUvMBjWb3cz1UYzwmF6kPMn57CyI
aGpL3DDfDw859NppVLxD7uHVfyXCIK5BiEQ94BM3QDLzdPOn+4bvCrb8qoiZpypEfK31vBw2Add5
7U9bInVC6er9cLEhCE0fPm4KvlTWRlXT8ovGcDtW7fJb9mDntALw/ZUCIxPJ3PYVN3cnVTYg1JV0
jDjzkT7dpMCn3S1J2Xge6uyahqbj4QclOnoW+JLVknaw/BNwaSuxYz+D1tvQNwOiMSMkJ8FexvtY
gdj/harwplUY78V+7/9dHiL7DiWrQ5GRW86utQ8TRwGctnETN2qUC4DIHNfHz8EE4AXLJKyEo3RY
5J4UQgPUGJveqM3bzvNtzqNTwYnezCnMytcBcDYffHLHNaFo83/YjeR9+d7iF54pDlXaEAJaEbwD
Gfhd4a9a8SCuW7GWuqPSW4OgJzVvHmK3UP3O44pHOhAKT1NMIbb2QYR9ww3Rdqh+iLRi2VTTB2bE
roD64tdDw2tgsRxPmuzQRSpTW7M5ykNFRVmaVgLksaHgUtDRLUURLTjFWHW3amJwLhwXEZe97EAY
uAxOGDZkRBkk94B06nAgOo7EiD+pLnBUDgmFBaAHmJ4HP6Vqzc1gpXCfT72YtvxOdXHbQupwKgpE
wXeCutsQmhPsgcrYySY26VLYx5BzxCzvBxFm1CvdAVoYdt1a/YAELS/Uq2M8WiQeQhmq5bytL45G
cHOmC2SSo8h8yTyZ53Q1i7Iu++W82uGUuAaHHYWP3vtn4sNwPiJGNymagbvzO2jspZYeyZkw7qKN
8+T6CymOaep0Ydk07d1VwgXlZCosqJgRPLGVIwwWGHGO2hMErdGdEd2I9FRnRnCf3PoEr+0Q40Wk
elZM/EYTCbas2Ha1tBCWTrwjsBdOt4L6ctFw0rScF9bmYDPVjhKeQdY1jYTR0yQmZWOK24ofHWcz
4fyaTXu/GELwa0nB8VIMNEIK9BB2Q0R7mqfMyUItQLFsLMh/ev3USD2d77AX27xikf9URsYOsugt
69fV+f0IuMThU4DeTFk/kq6+AGMEAbDa1QAccZimJEfykkDVr2iLUFj850J79WtYH8EEqrXEoATh
73KvnS62sXG+QMJBEANhryR5S59k/iWqbv/SUcVXdz9sWtG2KrNXGOrvb8c9DKzPvzUS++gAwhJ+
H0Fo8+lArgCp1U9h3nMTPCZ3ZElpmI/abHD83m9ctxBBTtK8O3it+PjDLsfSmYOGFkP7QQhKrql8
SgTMK0zXbguIFiDh+SfDK5rqbfQf3pexbcFETIczU4fmMc04t0cLZUPfOicapS0yOe52xWtYURoH
KLUtKiA8odKQ/0FLT3TkTKsVsS2kTNbLS/nTs03QJ2ugP5nyozkVzRojooCt6zZw+C02uAg8l5x+
3R13FXTw+VSyn18w5sVOzZkJpCO9CmZtS8cP0Dk75h6xIvOhbGIWtJjB/LbhMZ9CAqf2f994EsX0
awFDz3Y/T773MVhSiYstJlDzFzebOfxhYP+s8VE9oD9esCHmZiDj/vqW2zRm+HkJgsLehC6nQuIV
fLBU/9NEvMp1+L0bX32G5cGWS76+EajRuoP/oa3ZsDW5jREbFYp108vv0p48lcgObh/Ki8xOGRZJ
v5uGNARwaK0oPAM68hAzPZqXlwgG5AV50Yo++R7wb5tbnWcFmeRNocoEQwLnJ/r/nQrJ3QTyzaSM
Vs2HUDD+n9gvoSQmUWQ1WdNfyTEai4+54wNPIrUmlRGqOs1E6/SEuos0MTk+kMLqt5pD+ELVI0HK
/tzPopBE7SccfGxeHYPA9oO2p/E9SayvvFhQeKwkKI5iBBhbsD72agrOArJVnSa1wbcHPaLu2Uz3
ZBe/8PuAB/A7EVIzuDt0J0EUNV1XCJAWhWxnTfj/ptf/D3rZ4Gt0ghjnVsrjpFDudnEwlei1NWGb
jBbogi9ka9pA4oF+C/HPWnR+ot5d7OlCHHfRrO+TWHliqhSYZpTUpqCYf+yjSSHG4l/jB/nDXV8M
lDpPbHdIIMR9/ahg2QRpF2SEi29X7jxRgDqmdAAYOgKY51LkdyqmZRHbpa3ivG9lNwfifUmT7FEU
Z/mpEFS8xViDteWCxACgdcHIfE8ZvAjDUdCjLKAnNb6KxiAZaORrlXW7y7g6W52UPSQPfU+p+49t
xrJFWfjXogglSfNHB73sr1w/B3znc79VWq2fr5UcWKJaFOSHr3Fp5IpeLy901NJfd2zV3ZVGY1Qa
sum41iW/E4iUBVrQ4p+bQPlo5xh1xI7M6Blj88pQ1N9zMZHw9xuBEVr3xcTo9og47xaX5VcJ7rjq
IqM8Xk/Y7DzresSFaGq5kuCQGvT5HRw9OMO/OVbRrndFEpQSDg56oeob+w+TEBux+zyCbldjCJqz
iMAAiRCX6IsXViiUVS8dWSeYe1AMXh/L4yiE1LvgwYijDZFFLKicUuDtL6pmDRSjvKIFJtzGOzW3
vwOPzP8Cr/sy9WnD7l3+y+fuJNQOiXgKH823ZAEI/Y9u2GxWdhESUvaIVuHzd/vu5iTdjUnslJk4
VjwNQztqXfTXdwPsuP2fHacC/W9WZ8ajyIW+O1DxoCbgHqWl7iCokReWMXgenwrity65H2eoU3In
idtZ+JVyztzS9z6gmvVa3gcb/YUasnI/k6cBT+CK7oMK5pSpU48wUvXQxtBEDMlrWTZWDn0Uhg6q
wGJxTmV52MDm1dSu9bGQfUytjHH8+zhvqGDfrQhyqYtvMkPLYWaF9s2ynaeBzx2JyYhEBddgbjfm
gpEqLAKe09uOIlAUSo6fN74A1RKX/PBNDvFbuFqUrLnwzkiFQdsxKmCeyW+7ZYqlXsRh8d1ADX43
AUguU/yOVpFAKd9t/LqZ2Rr2gNjjXdUOJzQYMNARIT+cqF76dws/5scOjnmFTYQwCAxEZBDd9jfM
ejp7MT2P0oqExL5tU8f9/KzBeMKxvhc+FAh3akD7jPWdUixj7tZpNnU8D6v7S54bbIiU40jk/Ig8
DCNPtZ8KzXlH/6V958EVfPmRc0JTdHZIjlH3DdVrzvEKN3XaCvUQVc+7fw4DoPKYJ/HeTlXjQaLX
imjoF7Pz9RZG6CzhohwmMtw3GYrQtyYVbpGFiYEahmtBUKhnBZEzqvSl3gHqiWYD2QRp4ACZLC0i
RwTIKtx8a8jDsSga4NpnlF9oOl1MvgZvHw38IsysRKplnjoONhnoK46jZGOUs5wlFugW51NA4t6y
idMN7e9qatHHkS9sksluCaQKT89lPg9uPEfPMveJfd6aQNX6qBWQxVSTSDWsgqgcG/IE0pxj1SZl
6Od743KpGw3Lvnespo5/9ofuXB1HMcXTRxtcryr7+fsL3H4Du6RkTslPe2rvaxdID4ivJJGagByj
tFOM/MVnZs39RTWu0tnSPgCa+XKgBuD15YH6tHQAcZb2psIx8Dy89GYp8d/EFT+Fr8Sf7hR8dbui
ywJmVg8ZUmHG5C9UdDqryiNr3UqidX+JFUjH8UgBKSLW/I06pljuNmqN4yU7Uw22x5E1BzXCHAum
IJDLZhzOeTgOjDN6tvZl8NyJGSPFr8RouGNXTIlyuHBW+dcl+8EaBu4QulG3fLat6e9iO8AlbxJt
ltjuRfvuizJJsnZrkbJSLOUQOF5q0porevjwK51ekHmdHMdxJ/mueUpFH781l9cCME5C4cqKbCN7
kF2+UdPHCYc1G87ck6nYz9yzCsOjjZTlBbBTq/eCyXDfsaBd1WuCPrs4YpMa0tcAZ5llR9kEDc9M
EqLwCVQpYH5/vyyd6lsRqqz2xEdpP9MnrLd8Eqi92CY5fgxxrm+IEH4mTdxBfDMetBSZym7kMjUl
huTGo0yGtWgE47H6akGt8euba99BSS7TYCWudIGoTJVWM7w3QV5aQFB9OBO7MGkrthg6blT6cdiI
6eJq1txGveuppReSJ281k3wsevj6ny5/1wUCVzKNe1p07BEO4AtG628MH6H0hcIBiOYu2IjxBJvd
vxoHDS1CYo1viGYbN0Sf68mtNWCU/8hTNn0jt4rIwhIXm/hFwQXLBn4lmBMrOjE8zF9JsBFAxwot
rME5ZNmQGXDxhrvUMg6njKoWQeI+9T8gvJbjYAn4c+CplWskySAiibB97s7bhFoQMFgCVR2ep35v
dgxPMAUXNmFQPSgYc7hmXtnqlTks6skq/+IFi22Ns/l+NpJ52/ypNgxgyBUXMdRUU8c9f/SJ2iCO
MZYLCX0WcQTptO03+qLMbgVWlKnCymw6MrJrWG9yTf/odeWDDxVC48pTSQIWjZ57+vKC32JnQYlh
8sTAy43R8r57Ha/AQcBv0VECBgbCqajjTppUP7wdRyYUKPxomxKydEcwqaGIpkiI19w1IOoxcg1k
VEa0hAqbQNEsT2jV8mX3Apitf5FexJGynMqsAw88wf1fGLBvMjB9sjbYXddraNwFsHQ+l8IkA8yH
5iswQ842ST1dnc/y6CZV4otkhtqk5hytps2FrHlXnzHH/loRp5xUMkdjzIGVaE83uEhIXcFXRfjC
5QIJiWgmh89ep8ybGPogsxrsos4hFbUgUrkopkXdDQRn/xRq6s41a6DrIkjfD+Cfj6nPQgc/2QRj
N1eRjwyTE9X+aSc2V6UW+Ht61qgKfALgWs7v2v+mS6B5ro4F3MFB0Ixdj/YrRTTTbIZQmItzstvs
Svi+VUSJ+FRCloNRonoEzLk6WcmFg6tDie2EvL/wsx7Gfs6aWZYAGuEkKUchJo8jxLmD4rcB69bO
lp+ofHE4b/J6tOfnhlKZgOhUixCWYSwCKzunX84ZxXx0SQWXdhR/7+QbEQp6pr84oob8jz/vV30Q
QESLL7lNAPglfTrMux/RKe/MY++m8vRrrVcIvTG3twCRSpV2CYTMYiTZvpLORMSgGWzPaL70dmeT
ICx0w9Ctn/pqMAsb/qx7PqKjZLJFQKgOmC5xnAxczVzpqkgMqBkqrXWeba9DzWfJ0zWjVnKgbdHc
zgvZJJBLsuy8lLnQzPe0dD6/MiVxxdiojt9k/X2DsQ+lul9mdJu6qMNBwEKXDsqlLppu/N76aT4E
xwSh4MuzNyWo2IKmqowys7K6nV+NA7l5gh7S6VYg/pOlzYQjTeb/DYEw7iaHavUgPK8I+BrMhq8h
CRaX419uTwOowpjNIbNvooDWlmdxA2oprZJu7HyUrrYGDjAJiiP26Uz164Z9WsxUIUyVKmdwwSa7
tBrf7shfy0G3JIV7D/SHs+StD074rjG5zxh6Bagh2KdnuNqUgk2XaaH9gG4sdJhuuLS20ZGf0Jdn
rqpvOAEo5NyepN37gfUoajCExw9ub8SRhXYUseBCwo8yPhGYDAD9DYXw52b7T1Ucy9EO2+Xer8Vg
KeUG+p8SR7+k/UUWcQy733Nt3zWQOKbdsodo/3rCnyz4QVnixdwW5l5x/t49Ecf4qakA8CXolQVH
CkqIOqyCDUTlxLlMj9jIJ8YtQh+ZDrSR5uGK8SMJE6cAY8hrhdpn3yIwT+NPaiMp+IaN3u0kW3yH
SMU2hCuy/+H9K9yxOExjJeWwY2+1sWtaO9YS1YUlaLqHR2n7/OstLGqt07Cz4wyqdbmygel36iJ+
B27TQ2fhkrUzTaaf1mumeLt87SP6ArHNqek0yPQy7FPQxxXHXh6kok6+tuQHO0MKZ3fO89H6SSXz
XYqg4GjtyTvoW8nt4nFtpzqDfz0r40vKcJNEKQQlkeMIfEgiJbrjILnpO/px0MKp+omGjj7RE92G
x56bShIhyvEpHz7Z10mKweQjPPWizYFtAgP6K/9Pr0cVVhk3ulKO5NGo0yV4y+QzmOLvOWhz7ezD
mPRqw9perico1aQZS+0wEezMMOihsuJGE99SQ0mLynRNWmXj4i7aSvXFkC1NE3XGzlpLfjARAnkN
O1s54JG2c0iNVYSD9Ro6ODWmJPSUv/eENQUvp2TLlB/zlZ5kivqJcJTncWvj4WzijaoO0eFpESIO
GPfa6gvcErkSsMNF3V7R66tw/Ns0sdGzYeCEmRsD9q4uFSlp17rdqKSks3huJ8Trrff4DqpuppCO
6CiAbCXPNTXTYibUnMGPjadfWZ5hN2Ktntg8kAzkHVSeYClZp3KPCf9vIuQake5ZToy0XbbnxDHm
01v8B5rgHs7ikxPQWi0lpvq2+yMhivJmBQmjiRPFIYYFMOKPdPjcLz160VeQjmTZNTRs0n/WKvxR
+WowlG54BaNjn1Wux56hk+BMk39AKziz6HGUOQjM+2P1IXFZFUCc/otACu0J2aXWeWUZomNaYJSd
WPHXoyStnOteQ4YrpewQhjII4qHhbvuOHvMhnG++bvggW1csqMeoJe5hMlP2dvNSZM7kM6Vim59F
jNFxqmQcwSIIBbtzHIWPPGC5/Rc0d0FIP+BmUBzqGdPpGafDCTTDjsym7hcIfMPA+9vylP+CxloD
5bG+dDgZU68mnQgwCIqScUH6WcSkwHm55vr2bihBHitHDiXd/jWT+vXXgtXvyAJYZaSelIYgPqAh
gZopdT4qHkEJaihVHygGOt1b3tZ3bHN4h0noUmP4HdNrE5lZePcieAp2pk7f+7AcizCoidtmmJpw
qTUML3sLxW+ksHYaA5kuuwc85H7oFyDPmZHys2dQCGHY4dcHO8LR6sTy26RO0big1A6rSvTyvIKk
bcp1M6bcfU3fAiJmVLc0kiD7VTi4Ilq/q+8QzbwOmuEoKLEC4FKMmAtfCA+liTp0NS/5tBvNgqfM
pZ+eQNxsDElDrb44CQGp8/26uYZbHFJsEr2hZyWloQsO8bmxB6DvVmduhUsW1ItdbJEk3UU+6TO+
xfPJdiWBcetUTiN5pNsP4ofHP3trLqt3G1L2/MrGop3ms23IpcD4hnD5y6cjF5rlrgqRg6J3rcGi
M+rbo/f9l6Ut483pomDonEgmWHsWDtrEGFuRjgMsGVw30GenlgAmpLsZQ97VZfW5hUvc1Ml1oxxg
UtaP/USTMpJLGRb+h56d2XIBJOlwJa52F/4JuHyaFEFeWLrluN/I0I4ULDAmGoX8dxQui8meP7yX
kxPkB+weyhsjYFFAsX/aIhcl8cHTER3j/J5ABsgPVderjyee6MTIAX6sxHmpgSllmEBRVdK8D1k+
KnR52o+xvExVm6JZCDyggUCNzNjJqBKQyC/C5n20ceLvl4YhPDPkwnhXFXyU7TgNTtjozVHRK7W3
sT5AxypbQqsdA11D8Dv/1liAQSOhWsNCG+s449t9ok7WujZtv/4iHxGD2DPOdkoi6P3jGtjsOzRd
qBN45hgu/nmIExP6q/0vdLmqkJTAUUgvlqRzirPRGSinjXeef2bzEciktDYPb+UfADiA4/GAlgac
DVtyERFtknECFf/siFUZ53Zg239vVed8Wuiol1Oqt8HMu1TqnetDoZt7AbXBaUSrUZ1C5heNnHl6
/99uAJp4ueGwAohhoBtUNCqa818HQCgrjrhS5UQdknWFmlkSZpDM+0d1Y/sTA9WTv6XR4SdCnfiv
RpqRhnRjU+MqP+1GteyqFUKvVbICDkGGOTSZu063G4abjXslSvQqYaqM4nZTe5iU3Wk3R+Xv6oOZ
dQYM8T1HI1j3J/QhtF390pSMw+GPK59WQ2+3gFqcDIy60B+HShP1/Ei7p6ygt8FUSqfOwoM4ejs1
S3NEbXijGzH8MGt0NSjbrH29YYvP0cm1fS6F7LnGn+UWkS0Rz+GYbSrliO5ED9DbOikKeQvXKTqK
alcJwmG4Cxnrc+Stu7kRSc2YzVLNnX/wjdo/b22K/xd4w/sRwr1WcekO8T/V3+FNjzBAVXBoEhRS
LLDmQPAiTEekzn8aYZ1KCfcwm+d6dFp/GjCKgTvetDJzKlhVOjojnDO6GBgfi/YyMbhyArC8W3Az
Dw+Qdc7Fc2G8n/uX1cE9SEAlIe2CEV2QbcPK9+Luk0TaQIhpTsrtNLa9PhvVgsF9vDWCBEtVf57f
YqwvwHBQVECrXkm7G7sL3DNqBb5fbczcZ+TGhySIw1d/d4HW3iAYc2qvubaZjWuMyNmVeIMtFzD3
k5XaPDg90hG3MIALsjuK7rs1PG9K2h0LcwjeG6ik+33Etus4u3FAy1rsrv+KS7kWt24dO9g1+aMg
NcKuBG096e3w5CMaeDvPrPHIA9pIM4FFXClTja1TEtvjA7DGnt3kl3rFAU5t622bHeWimuqZckZH
h1veGdAAXwHl/10zCdDZMHznncm2+g8FVRMzxlIpRUekhisGsGWndklqVLJzn0S5LQAD70uQ0m8m
XxapFxG6pKDaVVIj4A+BBwcDYZ3/FTh2pdkJinLQxIhwt9OjaNeKebzOmFQuV/O978i4kZC8yegY
Y8FDqBf9N0MyMFIRdMQxnj3ywo/6HKSYW72HGdto2kJaTA/SMS1QKiiahytG2kZwGJ3LbEpm6wqB
0Zr+gdyL+uoA/OI8Y4ScrUFNl8EBF98cIxFJjSG/t97ac50qq7XyzGXo1W9L6KAxebEdayZ72cxK
6NiqTKquF4WebtK45wzZ29XvAjIJa6pzDGSHPzVzmrWJ9kPEaOHN/GM8HYdp2d+5dKqxgS2gJNEW
IPfAhNtv5+oMwZBQJq+EmO0uxX6lZTDzj3uboGeT0dHizkFontVhj7AEoRLrh9EiF5UJLeTpc6RM
jKDDzPILbd5el1EblhYbJqr3JWlXwSh65q+ftzOG7LjZYNwkotjoHzkQpNZ46+myLYgAZsK4LD1e
LHY3F5d0cHKBPPM4+rYPgJeSlgw2VCBX37Gp1hEgSMWO3LGLIe8FNZpT1pGCPqkCNQ06Gv0Kcy/0
iGLJAuYel7sFTjYTp/I9gLIs3CHvgHjaaMqZVDPXtRGlertlsCrw6whrMB/mQGZahI7ogxHTXNE2
+BDIrBQml8pNAGvYzfFTzc+8EJHZqHJ+MQ2qWkW/KAe7ZfCMAl5Xp4Uryc0eosJ7EnDrfYPN0Of9
1GoWNbA08kFI/MjVEwHsqVzvFMBJKMdId8CIeBLyW+pUjtwA6lB/VTmS4Y2251Dl6Ah/7rc9Y7fp
blAf9rEVYmWQubQ4lE0AAuJGHb6tg15FJzWqCkSL1GLL+a0Jg94lzz785NsapiO6skZ2mTKIJiwE
MxAFR8meVzT7vKR7qtGigCsd/93+PEjIxu313u14DIimwJHhA8VYITIV06gij4TZiEBMtR3nIvWo
R7qAtW51i0qOFtw3n/XoyGH+OfNKkMV2DJByTJj2tKD5zFk0eHnlalFVgGy3wDYwtZlWOcg5+tNZ
aHWhqDJkDLcus/FTtL1KIULkaCnPrCUl6l52OG7KCiRpB4tV18s7Icao18ewvuKJX+oUhzqeHx/z
VQHpFGDc/HTooWs3cvZYDI5hk2EYXQ3nM+NsEUFzDmpAwPIQBc8cEQi0ppK8f9h+vVEIkZQzhHq+
tRkuHqyV55931jIk7hGdVHZKjAlltwiLrvFA+tajP4Hs6r4O9M/ipgH+ROhmFzQ9QER5QZwx+lmm
/2+qUOmdoE3o0mnW0aASI84yPJHYx16XtrJPM71+BJJRBQgzv/ikWdNd4lFxzw25J9bcPdC04tFf
RlMvyZjjc5zY1dAl+vzhs3IxSO8ffO7ywxzliUoNzRBCRR5gIZsEJkRSVr8JhDZwjeZmL+DH0MT0
+ghQLvt34JLPBXCbWhWuR2HYOBX6F9cOr4fFF4vIhxfhJpwBrttSydZBsUZd5L9YHj9AxHW4AEnz
hbBc+77lxiv3uIIArtAYM7qMsQCWbZhNkNBacBBV/YowP4KjAUJ5CpkzJyZfXndPYl02WSuTc9n5
FN4KFenpSLdtk+wbvE+L277jYrK8v12mm9T/+Y6puICL7rjD5OWECR/VHpsw4yBSSzr4hKz1VMNU
QLiR1gcGA6hWTDb7h5RZiV+x8Mo8wlUQ74VYYo05T9JHKcTHAtWAFxH+BVMMXU3U1p3h0A2Y0LH7
re3uv2I0wGoAmJM4yNowVR4UXCBwjyk6q5lqAlnQpcEk9212h6y7unGjq9Fs0Eqq8/iokimXbGcf
tmsgJP99692Xi1N7SpILJeEodo55UQ0eeRwrePdHg5LRWAsp9MLoY1EOLuat/M0cqgZmL0dgS0sQ
3/xuL7bUrr8P3g2//8QKW+On70niZdgXnsAbPm0HDJxJxnaFU856lWR03cIYkIXFpEs6AoqTAGyU
mDFrkMlg1WdtNExlr+fXgDqvbm655BCoJL925Lo7d9RDIYgWOnbcwKkn3lmwaI+C3amu/ZakF6z2
fdW+gyCFlgoxtFNsThRDZsIKqjiZ47EDeoW49N5VxViJ/csUybcL633Hb4M+SEutE1g4NC5rWbsM
Yo76fRpfPu3tPRMpUzeKrBkSAC7y8sPF/927QGWH0GT8Ymjy3uI98A1AEClkdQz1uxK8WB+Nteun
EFQiHK6UtCH5kNGrtvu2GWR58ya4eWyqjQci6aA8T3r45zm++Yyxj0qorEPleeiZ+VB+KJbRFujN
a+HbPF3Wo+PJCLxWp17OBwvFOLpkF2NWXkSxp8zilLsLXXZd1bA86a+7M1iwhW8n7DKqRf0sqAsv
+2bv2o2DZC2NgTFxPAV/DrpUCbxb0J63YXEjEbM3qIM9nWN18fPJg67hFilG9oGV9cPJj59DQF5o
5rjQUh5TSKGMEyPzlxbHiCGll4KC31kQWKcQzKjuFrQRnkxIoybvfLvGqI8aI9DqeT3yT/n4fj2U
RUPuCU+bwHy3M/e5ZF7alMzVVXQ+YDjKiPrRhW8m92e8tJOixkEmGeuWpchPIQRLUX5nUBoS0J8c
WeaaDpiWWOjwrh0OfWN96w/YGbU3mocCuuEsO43LGYcf3W8exW3tqYlqljtusVk9m3hELVRfL8cK
+yVO4lh9Jd3uC9PKNPT6UgaNwXc7IwNmBBPKgcKlWMRUDCERFUP7FOqndZU46mWZCSLq4+jA4Fd1
TfZeEyig5u+qNoP1/DD4qXHm2IEZfhMyvBH4y6Z0CGpF90w8A91jXERKQaZF5FSp2Wcp/1+EI2Vb
WPXkK2z5Xkdvgj/6EGblG0B2sT0n9sAq5UZQZ1Am11yqnn79mjd8uMzp6bLqlayWr5Huu7ouwBSG
O/8Kmyef+BBspyWA72eEIvELpGNvZMmNrNR8gfN0X6vGD+hIJU7r5VV75DcTrKU1Do1JEABN7cG0
kxd1wwsFMQYegwIMrBrXNgrORMZLimAWRNhHdVD5kc56pST/OBUmBg6Gh2c8nklxZeKpJGuAoRtR
r4eCxbnLzUGBkPnRKWomEV1Zj4flFTgvxnnU4pwH4hAEzz8oisyszT2rxMOzF5jetWUiDSalxUOu
j0uFIJCM6zLG4Pz44Co8ZUiAtIiEh2RM0F26jeNNPkvnIdvk2BgXnTG1dhK4pzNWwMYsvVow590y
poKtZ0R/5YMhdk1KHlZbxRLeVkrZXLcVYLZm2cPxVlAplfD1532zlQDaOZlckHINZf29iMDOC3H9
THNGtZoEJOEBVxKPEe+jJf2pOLJt/avaQVvwGBaxkaO4UxpINXTOR+ufOQzbxD5dfoY6oFxNeW+N
tl6b0zCRWoZH0CJomrMGLGUWO9UfyA4XEEOZtX1YBAGZ2Khsz9fs6Kg68kxreLdaSCbBV3g41TU/
X5eTsk0g0iTXVFwRb4cbIyCVN/y7CcK3Y284n7KhxN8zI64ChstvRJXeFIDSy7QYTlvss5hI6ont
EYDJxh1mOOa3gpm2ijjssOqwhP5NTCb29YOvJX8zm+qk9BnKnMeLvOatGwI2WNSNrnR6K4+5UidP
F1x7EFJKEozQo6mHcVYY/Zq8H2k1SvsPEjqhfhUHAmCwnJea5oPulbQlk8rUQLKWU0Hbi8vzAh1s
lA9mPmLapApi07al7PGrOo0crs6DaZwFPbI0R9+lkfhJeAu0vESfk1nEwL9Hx2U2d3euZ4k+KNKv
nkGFCCN2LhpsV4dRfp3FgRtv+fcCKEg1vMT8/JejSPumbAXvN/YFtZkucEfk4Ce+qahDCbHFpkOW
UhSgToVrKbX5d9zi8bow64awkFv1ZP4WFB0XYjSKqmAjJve67ZVtoXGqsZ+nwtzwj+qrOwFh6d1u
r3q/+ufjb4jcJ8Kcd1y3g7aInX9nAcxhCZhw8ovDOpsqb7dlK7RU9DSqQrOFVBLNGlRxTYLS/C7Y
3Acpi6cFhsuuPNUnHkQbGM5/P+tuh91EjxM8FpCqAm+h567hz5IGyY6fX/Z66WFTc3IKpw5jbCjx
XbtbQ6/OeJxSCrw1jxfw8ZNFhVgX1toyf7JU0lXz5YCS6x744Gedr0TSxE/Am9m3EWx2Aj59O8n8
0L8T38vX2UZWubtJua6kvRQ9MBnpqR59Z8gp1bAXz2/li2jHEikJp5TeKfjmQ6rujQAcZ5sbNQN4
hm+tqEKZnx0Gr/0uH6WJvt6BUJPK4sQMz44PISzXwz1glrO6S8UGXooCvhvEK1ZA7/HLmBOeqQNF
QsK8NqiIm1nWYmQRZUaTQ+zvfeOmYhSH79hT8em/4VtPQOLnECpfOeGG2b2PB6mXfz6zhMGisTxP
9JaFsF4ToC+as6VaIUatKJymVTiohlvWLosda8CrrHJLZzubS8WIW6BOL6xQa8IVeJRn/nSMalk6
bUAYW0/K5LeY3tCzra5D0Z357h3rVbpUpxxtSCw+xR+FL5ISpyJZDOMQcg/lI3BD8dw9eMwzEihO
R1f/QBaVAak17Q41wX8xRTKo5iOcphtESCHN24hfJ6dC4pCNoq3Ku5s1CFrLB+uQTO2f8y+rE/xD
X+yHdJ+hPPYehvQVuH/kVb+6KPiDx1gd75Hc4UMlfbfZY4Pws1rFBP0lPsdYW+n3nQOtQGRHiM+7
B8tniJtI7iV2AJbXGDpz3N4Q5zoSvYGfHy0KN+2YiWEMIQ4uUzyae1QintmoehzFxodRRfRLx3qN
A5+brt7S2jLs4KxI7/LqLT8ZhpqXEegTzCKV4ypvITcqlDCQChDaSdPXcuTGDMXs+2y/91zOTXpL
sDy938cWbjcISHTb7P1f5al2mfXAp5MPxrwv0mnskg9ZcXfMqU6JJSZ5NWAKAy9MX//KT6WJ83Zh
i4jNJnUnDpIp6jTh33RK68DluOPsLf5YLYyWpX4/izdzZD3KRh+v2dgeV3PHDYiF7xyVB8+iLxuz
cKY2ta+x5WWUwFLovbLImuAryxr2UzhodlD0ABDJZHy7ZYITY/LKuTgP93GBwJ+0wqYyXp7+MnYN
AMIO2HmB4gA/g1Ix88ra1lMTIJvDC2HwkWr1sxfI/+yLnAQy/CK/ry6JsqU966HMt7wlaiU133R9
hSSydS0Rw+mIY49JXBqKV1YQupCyckDbWJafE5V2MQ7sCCY53q/BhDpzd2e+5BdS8Mj0+mQLWTnO
eMnvpU36SYFnXE8hZnKM0mtVen2qro/eLn9+Rq16XPAl48H87mSO4Tl7jVCZcKv5gju/xgvul24b
Kmg3DZqE7S5XfXGmOn0vRzwNuTWjQDicAmYsSVxpxyvTuVF22i44IWINzwNKJM8D9KQmmrkTTJS5
vwUBLMhPq0bRpPGEHsLgsZFmPVuQUrQ7ANrtIGVfCgQ6zUtHrD/Q3/m7uK1/sNLljcad49PJmpeW
blbj3FAMp0DsgHJRnu0XyMr7bv+oWO0egYcjLySAglcZzCUU5wCHVoTsplhksbbzU0617ENTSZJo
ZxGNDijTB+5kZhjII7Jhj8IhUQ9uW+wnZbtQgXHnL1RPtpjJJtisFmK/TC4Argkoeg+hqIclI7p7
oRJLOmrmbyjrMtLgI8NfKfARPEHtYEiQCqjpTr/XfXb3+u46tY5Rcpffnj4V3niPPCTfi42pcTuV
NIvM0WCtK3g7oMr97Ug8tJ2exJvfChJQ6vNOmZGdrDnZVi8E4+cra0FING6Rl6d9LK7i+ypiSde6
K+5Jzfyo7ojAHcH21iPhlbc+oSVCR8ZdIxBKjsVeOyZ677OENh52tABK2TWauJOULwrdpNGIUlgP
lNrwJfmrrRhvf5359ab49LASslfo7JXbYE1Kp1hvZXf+3VWIYsP6gcxNs/eOxyV2VQaRlJ85BmZI
WxoNoFSEHgZHC4Bpqhvn3Kul1rDEY0r1AFqlQfIP4pPvUptqH3BrerDIvCzhAnPi7jaR79JuHh7j
NB26OslXS/zr+o5z12wJNyxvIob5N5VwDLndeMZPr9fZxNhkhdteQOZZMDl7h3jUJM84b9tPpaZC
o9Q4ePGiWUuYomxTD2p/DMZVxSt3LNZjB0bnensaSS78WydNXV1EGG15x689RZZW9pzIyM8bkb6D
d72iUm7OTSgL2TdEDuHui0o/bWZ2wY9UEbMv2syD6qahujgySY63yUEgL7cktKzPX8BIdxiBHHUs
5V471uPZsa7zrBXgceNVFwWeLW981/UI1YtUOEy65U+dUxFyruTzY2eRzDP7cIwaygPgBKtI3cud
1Npg2YaM2JPLR1qBi+L87wIQcXCN8IYqGMOjdRTcwCdDfnLxjy4RHkpw3frosxMmlISUVaJRJ8MP
irEc8IVQAVMqByGN2PbtmhlQw8dgsr1yB5we3qI7ENhvhpxm5rNj12W2hqGKqR6O/txes2SLfS0c
N17nWShQ09bCACukEurzLZfIbOW13XNl3JrWCqhC6I7CI+KIpzPNEWTlWUSkNidcY5+NyILey6Ic
NR21HKJIlLDDZpIXoCIYroDRBf1ZY0Py/VTS4agPqpMFPJICegyOY+fqNQMKK/h5lIhlCnA44esO
mNCM/w0XgqTj3EPC8pxof2bmORPORl+/IY328ZDvCfKsGthGk70EloP08gv8ej/N8GQG23b98jaB
Gy1Ne320mhZ0u6rL7XngY7OyZNTk6cGVYYTEG4bzFyBVOpBAxSEO54+rKOm6s3VJKmqw/cx2srrp
aP/vyuI5RJ6H6aICQV3njeYdsXNGwV9ZGiFs55/lxwhbTtOZXILFstJNKTal3/b+w4FaQ3ZDpOiB
VBVl1X53AVyXPk2G2l/a1EQuwbJDG4cuJinG8LjgPzz4u28c9tMsPTV9a2dtWNFkQTyXkOc3AfEd
koZIolKT9b1ntJ+WZD3FTMoiPmLcdqAA1Iy7EiYrl0dCc2r/ke0NJHQKcEOb5P8NFxNwbCyH4yPz
H+kI9V+Q0wsTyqIdtTmW/Exu0San8k52EVo6UdjsycI0M1cte5e6bEtPyFVsPwgcQqty0PXtgw0V
g+LmmO6CHitY9/65fi8VX8aaQAe6Yrhx31jCninDGLtNw0LqSFYuEOADnEdEnUrA9zmBFKCWHd2m
pnCnKwncGLv7K0tBIePCqTaji5iFdb84b6sqzqCdMrNCySX4FaUu3FQ5u2tryegPdv+LHxWCOX8y
eAT2Ioo9a2ksMNjAR1EgNLrqiXCD5Hl7Z4CF33AAK1vm/4c+Rump9dLJ/MENrNQZLHnGBg7FzCqd
EAc09ACzsyWpMqKrVut1kLp3Hv0spFo6PSEcMgRxMIH/PLhuwztiwW2YgRcYS3uYZDbijm6QUCQo
+NJUqnPshzTNOOrU+GHxvEjqHUUW15/0WwLeM5BXwgxiAuCEoKIf0ZiWWguZGWRWw6crz9AyRWxw
omTSc3KMWGsVtgin6M98EsbC2HExR/6SuDCJ22FwqXJC8oCacu6TR6NahrNVSh3pBRM+nPAD5Dpv
5/7BbQ24G9Hvp+YQ9mmNp3KIKeYnypITWT/OQq4RJBSeliBzbN92N+T0AOrsU0XoE/L7QQRrV8Fg
aBLZp3wwJ2uI9x5i/6Pa6N8zLRtr63fwJ5fVrEzMMVe/ZhuwGqboE7UtjKPUZQ2VQqYZUU6Y3/45
715dixC+MNOL5nVjEiG5DJT++yr+tvAEpAUXIOGU5D94gCGS2hsRfB1BQDixKaj2LWTjTpUV5/Ho
QB9G3YOCEcaPxPNCs1w3JoOQHS1haLarnWEeFg7V62Jchmno+IUQAqaehtKOr10yA3pUG4D8ialU
2pHngyXwwqctDYw2NSUeaL0Q7uzJ1/ImHtEKFuAtT6mzXh1m027uJpB8XkKCqM6EeFyrt40y2wF1
NukuUPbFkl/kdu0WjwpoFfbo5L0bwHs2OrW14IRqeV/j5L6UENFhCszNa5Ya7bwvXN5Ns7TFxBfn
s9BL4TfaheUk1arBlviUsmrvfO0D8DH6IwEcxSMtoRhUW8q7M+0rGPPgF59nV5vltzXTZnN8vj73
UTtlCZXjSWm5SJymEpZFtxZvi0g12UvtWAv8F0y+16wqUj5WXpS89GD2eKNJQDWto+0CNq8YKBGp
0jDf88YJ7IF/YRnBaOeBix8JY3VbrQzgwfxNr4Cb6O0hfgFqtI9qSS83eEGHihNmWw47/HPmVFJC
NXnKeKi3u5fAzQTJyE5WXZNwiwHNrCKaXwdgJUV/8KG3Eo5A2Qw3BndHGy8AWFy/t8x39ICTCyon
Ebfyr0ykRuxKgCAyKmpFv4WBQV8pZjyj98tFShTKcdJRNbimRqip3ZgPQcFYzuvIQ/ron6DHJKyi
TAk8DchaiC8uBFxerNszBqFe/6CwPseXGE/1GRs5jZXkq8x3FmJcFitzumHpmBClibJOR1AQ8zXM
jf9S2t8zmtm/v3bV0FQaRz9unZCmEou1kPw0qkCwWZqf5+MAXMRNyAFC8vTFqpx9mlvvJ6+kdO2n
YznLwvkkYVYNPG9X80rb5DCxzD0WkI9urZZMfAPW4/rzLrKXj/7emOWVFzhyKHl/eyNMJyGqjFpN
BjCM3b3z4jB83O8i0VdAeWuNUvH10HQvmWHiRwsC4BjEX29spRSzDZHjAfCxwLC7wH80bs/JI7yJ
Q1qZKXaiRKugQqQ8NIJnkVWh0biWxvhOHd+1PwUuqaYxmLS5UvKHtX8FQ1RpYdCilTXR6KWHABWu
wjNis7WLXwt3N6YAJcTbaxg3/Yl8vQV8LXzfoS9NbZh13pSk4xzb+WGlW4tiQP6fuRoL/rhCe5jF
9uCsMXStbl+j9B8vH6lWJCTVDD23r/itIWNBTQ6sByNdFNuV4wKIcYrcl5713ue6IbSLFyRq26gU
jFTuY2LE3wowdySTXjIw3dAtQqhv7PyA3IAnOwsw5qs6G0+hjcK8yG4pdOwMiA6p9iglu7954Mm/
F5FzW4orqi32Vuj+qHy/uecxad1BWZd7RX7lA39dskUAdFlGCOnWfXJemOF0Q09GAvPp1zlFwci9
dIW6iPz+bhS0aezextU7czstyGwguA9FvU5OMT7WoUZydwurF/R3fJUFCRCu+itWMOGh0s9Z6vyr
Ua1svXe/CqIzIJG2oSpRDOBYaV+FHlYL8ZSeDqPA3niQvImI25EiHD2D6UgbQU4x5glOXB5zY4Vr
EohPPUUZbyf8Xv05MJ2EGJISnogWgJ2VmFcz5oDHvhJThPzf0OFACNdEwdS12X0yg4aZ23wJcTW+
A7Qw2z8hezxCmjIeIF6srLQEcV9lCoPlk10C5TdvtbB3l5WvWCqe2EHKqDJ/ebj6PNFGgeI+H3B3
9yJgY79cWxM0ysMPhuRDscnmof0ITzcm0zRhyyQs2frnjcrjjfsOa9sFiglsKajJxbCtEIh/sjK0
LwMN11woDg9zidlIQGOy2KKvez8Pb6pzqzJL+szk/P/vCsbiBotKNYfUnkJRcqogeDV0Wn0ZJT0A
0nyi+uGg0ex5hNE8+jZTFZI+cNgObBqPFi8uJwVNU95RPfofkaKyaWW5k19FJ7hxvelOrv06VsX6
wiP3mdkn+P0WvEFibCenDDLCy52faeIbjAkf296fve3e1T+x6bCPZFjhRXcrYGKZBPyIX3FOh1uv
QB9lRqsAQzhgw+I6YheYVWj9xZBRTGcrliX1eEy/cW3H8GXcdr2gGi2WKsQKZSyVbZ9c41UVI9mN
p7E8pFLyI5Ngt4w/jJTWy+NxRC2+e8DppveEykTuKfd5xCo3yF0wyBIg2KbS55GeXdpjKC/EuK8W
NBGbSYAa9/UAAQaT1cO11R6Nw0VVVedXoh6xRT2i4FlfVtg3alytmLxZUnwR7DD4a2LpnS0tCUkw
c4kMXrnMhxvl73WaaMY2sTSONe/eXPIkYgdwhqhRSM79BCEOtYKRqqffGkiSP6uTLMOLqvX45IUI
5dZkEWZn+cYdkzBV/ot3hWtqsJP4mnlKczPy8ODQdAq1/Qm64V4xmBrnMQNJ4qI7vUa2dZe3xuQk
OpCeXRsPOUigkdySffaXd3xq4srLnXoN+NQ3BOg4cvkDN5LNK8lu2dkPDnYlxAjn37Ged8XveI/T
l4XcRh9qHECs4hDE8wWIs3EqSsWR47cm99ib8rGS2HtuzB+b2pnjYjOtEfNtEq5g+Gz9GE5vKjWa
URdJUWL+SC4MbfPIiUp+f+SIvlUbRAJAFT3oBHQDeXeIK8ob3nuNZSkJL9kLRYPCPIW2TJwUt1hk
yGCH6j2yVN47g/3NjDguMsZKORmRBMlHyoU80TBtXJLJobB7cKbNVUJz0RB8zThd2KtTx7IIQOgD
0MAjr7D5R4L4GcIw9S4p8nbriSLDfNNG+XUmbDLKk491WH60Owb+RMtydb70UIqLpprNSah6LRAK
th/oME8wAuSu85Y6cW9CYuBizhse7/L7t4yenDjlQjnS6X1JXvMe99fQglI5YdVenhC+jLgEakFT
U0ChlBaQefYkM4j8ZkT95AGfshwM8BzCCxFwyTbi59Eem2Z+7aOoYk1e4fZhlGQ96TTQmjAfeKxK
nONyScc1Wh1BDGZAZP4+JvlcAmyL1nLveEVgjW5zbs4KuXftiXd7t/U3FEdPtY8C9nxbahO1e6NH
l/vvv2tgXP7Ug46QfpobLtHaWUXDQWH7QcUiXQKmB5/cXFI2Vmo1TTPCZyB6qE0gabUo0Hm0h57F
C77ixb48GQprC3Cu2XmgvCuwPH18+EIUjy6dlMP6JTbUN1yTV9O7C2ndG9z2QkTkLg7/vmI/NL2A
NeBi3pGlKNEt1PMo5LZ+lRZFZB3Ogt7lwjU9KjZ1xjyMZE8F/7qqcA4HiouRI3DcwNXGh7v5z5np
Tv6hmQILx4EmC087N/hRatACtn9F8jtVWjniej7LFwNNUZnp3rT+Z/nmAhU3U/crknuPoDIpbdHO
dLU1zJBkPXJDeQdSgVBWF0kCi3mDeHHLnhcUHFH2HERx43d2/dmz1FUC0kyvbQmu9AVgl1RcLlWh
INqkrraeBNJ0rHXk31u4kEk7yq/BllhxNt35ZJticScHFUCUhBGEWO9FGC+FUwm1ifo2vyAZuAvf
jL5iyTnfZ5V+Xxc++3GcMHZXIFQHITCT3CDjDH1d+nTuOw+VWh0BJGGlRPxzdP3IzsR282AFXwr2
YV5P0c4SwKreCNKhVys4MlhP0Bb/BHb1uAT11BqYVTvSHwHBMWU/vdSnuynzOtAuZY9X1GMiPUPh
8DXOMxdpbqNlZMVAxyWOfxJidZMrAx8bA4KsebGWcB2MklwJ9Em5qQkb4PoiPUJT9yKaJstO7avt
adBhm4ax32xMHibVn2a6vmO9lXmk0n5VeD4hiVihDDKHiSGNbhrymjy27UlVBXPFuGKL1xO6P+Cy
PHk5WoKDOO525rxAmc9AsYpeC1gvTcMY62tE4YTDuwHzw+FBc3vgOzc0zpxqh1JGxwwE044WaTgh
KnAJ7OATOZwaweHqYRRaa8LUez7PB/CmU6wjApeNEXCln4ndenCO5STHUAjQzR2emJH92ad+gRIT
j9Zje1RcYopyJYBZrZZGuKF7knr8m4Fs7Qrn2s2aOpwesgLyJVHXBs5+CoNUifLtgSXZiKGS9WCO
CIoe1W6ZLoEkPsx6e3SSanyMdGywkeWZS673XqJxMUPdPuzU3B2/O9tmZEXYHT6OhptYo2p0aC4D
8Pr2hnZgv0AVM9DJJTE4EYb4d55JHQhgZ7N8USC6Rw1PvkooAwbvnTbkMrOnhxzrC/Yw6yhoyVx1
v3UUlwO63pYHEUsDQ+++nF5q5fus8pHHNBZfb4K40pKIaCUTosp8FbySDkE5Bz6PFxXwyh9QX81/
TbT2caWYotHUeA9+nozoh7EtRig3C2LnI3uW7lpmLvEKxJ6rAPTmmv64oh7ITPglThYu9fQ698wM
OongiT1BVW4cU0rZWinHkv5DvYhz+9HBsEtUdK7vYZeo4nmyA1vwVh6cPGwc60ng7PhlPQzwxB7P
FQB0muQ08Ua5qJQ1LWZ2UTSvqPF9BDPzDuVIhdhX0Ykn89bwWV76CCNZlsSEk2DDFOWOcAQUVD1s
ZVYIrhEHjQ6aOs43j7IV6VRbJD5VhBbNt2n2op1qA94/IF5ztRvx9U7JyDLgdRe8Ih/rAB85q2z5
XzW5AIDD1x1IX3rDgg6kyLudbAoH2vOHsfBKymYAZN9JgLz2nqteIvKuV/qY3kW9cTsDKIMZPYIf
vqqOhIvhtGZFreY3zI7Dsf0oC8j2U07SLidGKv4bYhzrvlQjnemxHOQmM+ZTaL6EghPCzkshoUnB
draqvjWFcPon37GUK1iybvvWg4vIDYs+idg1whhotXOb3UYxWEAs7NebVXHChaMcAKNhpAv/sTU6
TPs0aDOOEN9zbNryKs8cyaEVf18ORkWHLina0t6cCczuLZowMHvi75hj632qrQ51taffcUWXG0T0
HuSCNBSujlmW6lWatQoPKVuFNnia/Jnhg+lAZqVnahDZffbiJbCMAULrXJA9a90WnTQLlIRkQHbt
gae1FtYzPFuz6ME65MxRBT/V9U8nUtS4Ww6TomdjytZFBUWRTzqpabU7RBow07sgE8SzLgVgp+Tr
7KG03Pfvav1BkIDiJHeG/68sQIweoTqt7d718dViVsFSJgRqZJPoQhOFtt6kDYG6Ze0O68qjgFXM
EaApbTuZy3F3w94N/Lfj3uTNtUPZtV2Nv4NTWnOSkvQIFCOgK//9sxeUUkEdp7BaZmGFaGnQg8QR
g/QwSPSEg2S9M3Gb96EAlOIVCkozddgn3q8VbiAjpe52k+5KxyRtAWHYkQ04VhvSnSGgmOM6yVCU
GDvQACFZy66oktjxuT6f+NQIv3s6GTg+wtnoHH8e4syNs8RSNY3OqwzWbqKjBwB4oeREwJra9Wq0
2xDvbhdWPEPiw+e5hqFpRrNsD43q0e1N32fgK3DauU62ONEhF3Xm/WeMwX1vmzeGsChiu6U8ODL2
tVu57IDAHBbQ1xoIL1qvfBncAR5xZXC+yxgiqMcKTEnk/JTMWIg3Hlt40VMxVB1TZ+LZ9IP8VbWZ
ml7xyC96w4kCiA749AhAILeq1bY0+CYxI2u/AxoT8YWoFqDTCS/XN287om2egyDVRHxQ1g4LL0Y/
Xfoxtw6xN+CKaf9a4xiWOeFQvOP6ODdLVvp5OS/RSo8Y/gV109yjjUrmC71dcBkgygaBvp6UdE35
eXEg2DD1E6nuotLMGEmX3XyXWOjoJIn8KFlMNyVzPNfFcGnbOP2g3oJeY9cJQV31Hn1jNe6WxhYg
fQOSy5pBUq/10IQmYZgCujHRKfC1BQlG+29g5NGpoLjZcwNYsdzyp8FidaeO9Ofhw4tIOG5kM+Iw
paKfcckt2fdE+ApKeWhuHSBkZMjOUpeLtbqC/Nz8K18X8JOONAKj0I1OUOkZOaFUXs6M8YUXsfDC
CWFsweX4Yg8ZbZFtIlKN155fksYnGmXsuuQPcW0F2lvwQIB1jVeayPsqSMV0pN49rQYORZg4EJ/7
GxEvr43JOD6Uw1ceR67j4qci/skih26tf6vKi3CzT5GQRzv/E3+7wOXVj89h04950GYdmjcG6k+H
m6zO2Yj4DhOVcO63sfoLDyvBvGyzDx/yKU2VjWkrJwwL/2v7djLaEiNTlCNBSNjLvRtBVO6a9kao
PkQHPvHY8vnSSUsUj6Wy9Fa23jCK41IWuir4BWkBQIBOsucyUZA+EeYKXHloXg4kgxpiGN2ESSH5
1gX0luwKPSfC3qdN/K+N+Mt33DWBjK8KkJRBwF1JTH+X6M3XA9jlegh+OTbQ2x1FuvdC5HnKNa1k
u3i6jQlves6VyABm1KY5vLIj8VUwexJB5FXlRqUJDr9iLbT3dDjvP5k7btW7tbCFy+7DLNkKBEFZ
DeN0bXTGFkCCbuWQyL3qHWiNMlKHVf2PZc8mOnyHwr4esDBc6tYaANeTDuLuZG9xm4CDRUcrkm0z
je8QMDpsNWzd6GyCbFD/ZN7ZRNbExT5bVKQ9/+oOcQ3NnOBkx9c+zWHBizGDU0pN7+dq9BF5FfdH
5mw4bAR8QV8lQarbXi5pvN7fqp7MGmqqb1ZuCod/j+i16w0ZgPQjtxyNzTZXIcwcZaz/ZK6/Y4+g
owhPEmVENS/jH7jL7yQ51fNkM5NkygQ/u2NCSVRdWLRHwUgza1gmg/VN5ljyLMtOt0DM1bE3Qrhv
wdMbwsAzhQ2DK8zVxUoTJbdaCkSK1LCci3iL+ba5BkMV9Jk8TQxDH2GAVjU2MzpSUonzK0jV2QjB
7iyajo7CdeKnooUYq3Zkad6vACORJylfGFguxivTV3L+/0c3E2ib3OQn0scCcU5Bu0Au0QbU4y+i
4iSVUtoigMIs6/o6Mp1SpS0+lu4rGtlzSqDNC3bX0IajtbaD/Fs7/oAmhpQyeqvP3OopcPo+5aeh
+oritQjFLGxUi7CDZj5QEw7920Dgvkd2cDud8hAzfnrvDQfzygwC5axBNEbEOvmN9XGB9cKLnN/6
iSxEaoTpEWMqHzS2plFVo8EWtz2ekDw2Q3n8tW21ifKkvm6M2+efRfigPdu2l1CeeKtv5L7SjzlA
URg8M0M7iJ25gq3qkLhVgGUnktw1bNRYj/VnFqCzWJRlN8/m33Sgi2y2BNGp86zMAhkLsi+ubJVB
LQoNh4Fu7mwP8Bf/1ZrfP1JCJsoqfZTZqko+bZglCtzdesOGbHlmDgrXin4qZjKUFPDg4+uGKr5q
9d0Mbpl2T7Pf7sGAqBfkiaEdZ9bclxGESy47j2sGri7gt7r9fF5uuYVSkjOJdZWQYQl7cBxWv8c1
8Vc4i9sMsyOaqGiCB5JqQXzrbZPAfnYSLgitJOjNIemGotim9k/oJJdiAJ/9aZjIUgVR98Y9XAY7
koVluX3OqmlGy704ZQAuhrYROFQCO6Vwi4z4tnK0932L+6hxi/EOvVCKMiqSDvouwqT1o6Ic6sfU
yqMpNrpCNbxVAK1pgH3J6l7EsXt1uBOm7pj9FV0ILpv5MK4i+/7y7fu1iKzc+ZDAzIm91FMyxw9w
fxICFIRfOQ1MoscQ1pRK6P0YrljJQDl33re3C3Hai6whUuaMaCZl4qjydfaJo+J2/Fr0oBjrHoqY
0CuDkGOzaS7fcXoyAv+BK2bz1z8gVRh0z+k5lxhmvgKNAd3mNzyoVWE7qdZh96Sr9s23WCi6RHKz
d9KqBoD8kP5lNqWV5apjUThFSOQ/UeIB5sBbg7hSKo9RQzzUN9yeqZnColFdQgatFjS9TqYAT/ct
NS1wxMwoT/xgg533Ci/KdLA7v9x0FRwH0qFaTxSg/nqN71aOI7vwuHqTUGIZ1w9AbHdyh9siGe7j
Ud23l7LoRJFU7b/kKKV/cTMkJHA2x9M/n+WNRZ5mCt47VMJQsX1Dkj2MiqMSK586rH5IvQ5Xt+bA
KiOio4+bBP6ZBraMGBiv02hgUTMaDRAVOyLBsnJFmeGwkD8Oc1x2vz4+csuosp2Zf/cW1S7SCi33
YMtrkq50etfL/cK3DiiZqRIfSzUmlFbWno8bXUj9/epkdcQdNJAN5SMfhWUPZeIBwJsO/nRqw0yg
OOr6+evtB5fCwkponVDuSB/QyPv+Oui1nyO1O/SL28rafFqQQ98txnvSApbV2EKdPK6MHNgsKW8p
hamUk7Ez9u6dtvFGVme/BiDJtAkVc6C0J2wDfPbCOVmN5mD2bIEgzcvJlMv1vXzECB8ESbXYrnSR
YPa+eM5WBa3vu++B22t5JJtwEdRvNbg9DtZxhlqfOUIE1uJuAA2+3ZhPRgoDRB9BgLu7pqazLHWW
qo+LDFDywc7/JnqIQWdFoZ6hU/oVr1LrnrypNG7h2hB6+DMTjs41afP+g+t+4IK3/C/daawFDxpl
ok7vIUMAQhdKa5d1UFd/f6YHJ33IoNzBR7DqOHnGlolanZ5KWAn+XLooSGTP/OFeHCWQ79QfUb26
Rgfqmo6i1FKMViMsSFy6ZWiXb3+WfaDEI9S90FNWybzojJEYHfHvtqDju6OvP3nsKp5O/kKCxY88
okd/FdWe+V6D7zxIC0g+bdzbR0z2uaHqFydyarhwyipdAH4kiwTC0mu+2e4FFzuiuJfxzrAi8Nux
YB+n9jPaNLN1UiORr+WwVkXrGekKLmqgFi+01FvL6JZgKbvMXOGTPn9fddUfuKzzwfd1OJqrAbfK
2UV+8Bgutrj1tEBYCTbAnkRSwWUc/BlNitU1KaDIB6GhmyxGVRX7YA349wm3WJhH4G/ntP3vH9iC
UP44fz5FNtpg5qxJ5KFhj4AARqWCp2VWna/TyjjuhACtMxz/lmt7/mw/zB+xKdi962Tv94pnZB4t
pWCIvxKSt2LviNOot3Ufl1JWadWZFPSfMqFujU24ViTSFDNaF4OXJ6xv94yxeU6cLMWuoqDOf4eh
Vwj4p1ZrED/zLmtUVT5nHiX6q3WHznD0E+NqS0OGGm1pnmcJk0sjRum6o9wr36BZhyIRH68jCvXz
4ic03EkQdr6iHXuVwuJMpe3QYk3vuWNcR9APQ+U9cDbr0LpMEYsC2pPUVNYnp7ifuOvDVb6sWeJT
mjIOJkDWD05Gt0QJParXzqVB2DvEYCkesVUnOtWn4OZI/gYGbOjmo9JJ0ggJsQ1Yua6zItTxckU9
cu/jPqSSRB+mv3OPy21xpkYg2YCY1QSoVJVYnVMYt6Qx/7cbpHDA67zKx5pVIVxEH2BomDK5Jerx
aFVk5Nz3CfAP4FDjtqP4+h74EITt14LsKT/ptrqUuzE5INd4oCZr33t8Q6vO9ZNsrOMROsOq6Yvz
zPu1wH7iHFmc0MkomQusbjwkgrOFBSJ/nboHDNKketbBS8lXomFD8MyHzoF3IDlNHPWs6GxeazJI
Tw5VsuXGzMmmIo1wLYnk5yiZEfAzrIfkaJh86YbHeW7g4DN42nNpIrJaktp5sWXRP38+3X8f9UmG
8+L7DsOEJU95vDsL6KkRDoe/Mj+j7LyKtYCwhADZPcO2Cc6Ku08OC7PHgaSYni6g3HDIEU+hSkdT
iw5QgTyid4+gXNxhe+TtHMidU9FW0XveVVamRTL5WgMPb+pCou2vpuDjka5mrC4ldj1GqEJyU7X6
KB2/swh3iD8UrVu7Bg9+aHvHNISCWDtZVNB6XZrQLH4Pql1QfP5GBlM50/bUwnlPphY/QiYUiJJ0
X/NssdqaKcZ1LqstCObk1+YLsRYnHs9utzHSFZJjuGO5eDTOjf/JybcCy/5wU20NrM6Jzvy6LzPq
6vin7TRla3Fl0MoU5RqtC5H5kyeiaS46QB0YPi7a/Ify1tSs6YFVTSXgu7ve3edMbEgkIz2UAuKc
WLsnjd7td4yVde1laCegy2LaXrPtWhEhhVYjwoyhfCHe9g8UWRpBaItmyEqbqMnZHDVv5iWINQPn
CH9YEbq5NCn6tOfdv0d0ImQnH3Jvt0Q7rlPRBr20mTECG0KB3ei92GdI6kU2Lk8el0ZGDAPzrlHB
Y5HPepBG/tMsmD/Y3Gp9QnNjX6isrhvMNRHsqCkvE0Zin0ApHu5BeSI1RJOYp7syctKy88TbrZ3a
XRO8q8z+gzmf0EE4+12HNM8o88GeqWIE4YukcZYqpyAq1kPGktOQPOlBv3CfkMRonBcN3D4DNqZq
O66yEr/XqFbmcfra2IO2UN1HRrbQn9EOd1eWlFIgc4M8lH3gkJhgBAUmRNOCH3Tm3qAH/wmHucya
uvCZ63rlrcpmaApGB8uZw05slK6c5SbARDf7wL8VNF2TP7F5SPyC684uszJ35AMMKm0JoJK3D8cv
qYX0fuiA04tIurDHAvXuEsXxlB689ZTmOEbBbnk1j6FkbyA8MAXsvR2BMJK5gJB8Uhrau58JIjAK
1CgZ4zsPCSACryGBkOecQGBk9kxEdqEx0ldFwRQUfCZbov0AKuDlO1TIFQyHcj39cPEDq7SQwl/E
JK7Lae5TrI+B9WVcrEvDYDknMU73E/ZvG2AqOg8CnaYguu6gxr5ifLT5G30KXnST754y5YQSwaU8
b+yg1qNdu6j5zTfw7COB/WgE0I5doji3kDfXk0Xd6ahbBCoDJmeWBo1W7f7itdgq1oOz9TyIlb/h
1MNLhwxjgv1icjyEcUZ7Me0w4xKeo5yVPQXDWiauNo0kXxJeIJla0Mcyf2ybEF9EKl7EldnTFxev
ADIwNe3KR0KJdQ0MS54tg/BFkrOoyL5NJyRYv7rYBie46MdaqsjjTXKNbhDNrwO+R7CyxV1FSBv0
0paYMEBdMzxy2P8wG/rTDw5WcJNxdJ2XNvZv/AJrl7+pUKnalfxIFdm2VAFlU1bB6IpGubZsOT7C
5C/WxpCMDjH2PV+PK4V94JYudtJoiXkmrI3O1GG2rjs0uaReX2hYOloeRh2ocVyLzWn2iLOG/ka/
05Ig7KvdHHn/sBmHFOEgBjA41otIRvXCvO9NK+7JD+thYWC8zREe/CyNu/DjyfY0ITHSXJMeu9CD
sF6aS/olIvQFn72US5rH7clLSY7LscteYBvOnWNIulhWcNqBhAUPJFa49oLZJfudqcMmd09xKaCx
QGioQMqfsKuGsOaUcre/5gmYZIRth+8f1MKpIaA+XJH2traUzoht4YaTRQ0qoaBWFz4EqXu2F9qc
bK+9F0JtRw2xMIsuMqUbaCDLNZ4pjaQQ33oEY9PQcHPRDUHy3jpa0HHD/b7fqIjO7jkxUtz88GY+
4Mm+LmnwW6vY6knHcUwlbEKV2IEpR6Z9m7jLvJqApHwRfS7SZXfHA6m89EtHb6XF991I1e/yioF0
GZMAZate39+NAaOaM2W/o2dkGMc+t6fSy2/UZuapEOU9YNPNgtqI0o2bmutT5JW3+SnNymR9BhLX
oRfp6UswWad4TDt2lMk2EgBnteR91WlQnJi+faE7pmOP6FgYwI+4+rMHQ1RNQjTwk1aKPRVCOrbk
2snYogweIX+1AuyLOtMwe8sLPt+kS/jpCaKX7puJmcWAkZkgUQoN/Jz5jvs2i/0fR4V6fZX0dK/a
bVxn1irdePNqsRZVM+60uTjuznZxJoJakjOTQck63anQZbWGu+BFDagDbDW7Gg+HSXy9A9pjtqhr
4MdOk819qqSTILyw+s4hfq7eJV2DAeSBLzjB1EZRLsXJTPX+UqZ42STQJjzECIOvVcUJsfOtaJZI
Zhx6icpXkjRu8uzDOoDzBUl9kR9OtVTyUGA/ejF3fHIOjFGPm3vJsD+5lmUpBt0xVmYfDZ1Mw7bO
ZUY4YSxcdFHKC3X8GKvA+K4hfLhVM2Cd7O93b3P1LjF3zJOmvcsWhen+qH8Q24nTLmw22DyZPc4W
wXlfYudL/NbEaLzkxK2h7vrjwvzNph5c1CffiYz2CcgCGsMPiQ7MFx+clnwDfkl5OBK78O917OU+
CbmTHVAarEmBKJ6zi1ObqJUgjUsQnJiRBXRPZbYX1OHPISELy1TVKUK/2QVajkbu6FgPNXp/LRxr
vbldbCcDRfwUqJxvkPGi0jCPJ+NBwAzmisoFRg+qhpHUCooNjLIiV6gEbvKFe+dSmt/ZM/MsAoBf
//4xF0d607uemo+eGOAYV7LlLEtq+1UN8Ha3Z7a3dclca/2J7T0Wy4LJiAgMjVFAFPKOLFOi44yh
FIXrvmQEvjqa6ESk8HYRrLNXzqq+Y8qlGUKkd9yB+Po6QwUUQ/dbZrigV5jAxzCZWIWXfydNlqcA
g311h4qu/HuSugw+My4fkhd0oNhMC/0fLSIIDik1SeaNgvU3pIvkrDB1KLcyMeAswLNE7LLqn05P
3Kc/BHgcLlxr7cRPUTFDoLGpgi7ik2B5JXZ8fCCiQBvBWeku27B0kHNFpo743F6eARNZ11HBZbzB
gj4GHlgNMb+l0H+1YKPuEV0CKvCSdNzVbsWjhTITigIbuW6TfBJ0RXBwPErk8rCpfrjie4JjJ607
8tEozg+mKFugOiLw8JZw73Pm4/3Fg0HxjOxoRVFJ+1pgfTU7njRN5BSDfjxei5i1HJmh6YfNVkS+
t3CpuB71NkcNLmS/nzZ4OSGcy04m3d65B4e9pQaIOSAEv6Hfs2kc8P6jRWLVKokeKI9NmDQeeM6I
0gkyK7mYiXtjzdr2dyva2bySXTONEsCgf7A9m4UTo0KKDR6bECwZJb8m7+XAzMxb5HLPQt8pyf7g
VflAldxAgq0TUsuRM8ZpzViqqYMMMEeWymxLsjRIIQDCHeWYofhuV3quoE7YEEX3a/RE+B/xPP2h
e1ALhGftKeaRXZr9svBiOgQeaSxqf4oCk4LLA8QhrmPuWlCMYPlQ5sOIuiGkzCvUnm2dJdAhHMnh
v8QJNJEBkTonUrA9LPmDc85OOcj9gXZen7/+1yXMe5zSCL7BGDVbH+6GMf0vhuK/X2LxBU7sQe/x
5FpKA9Y99IpFs4WywPCpNOSu6OeK5OYn2KSitNsxVn9hQVrO/HCSJa9PWcq9SwrNszzhtXiGZboh
3o1vW0+4uhaza4IvkwLlvKCjEVTFaeweMN7QYNCR34dcYWUi3Mzrp/bSZ66aiSHkjBJAYFPDTMya
HhBgHtcVB7/ZZBEIlBKoSei/iKJbeJNYR3OK7t2fnkRajOKZ637Eozn3NwCt/hsj6Ld/ugS7GgfE
I5BIvQGWnZ5Vt/jDgINISVHHvQVF05wxAI47jYVjgMhE9Whzy4ILPqC+7fCizxXrDOTCtefxreAU
2JLYk5M4mwYGdz6Tbm3pxrtkGsrbuADfsbq5XPaSwf5AVB3rYw5hSR82PTgza02lOK+xXzQNlGSi
oAJn85x1bl7j2IzcrtIWWYekP+i+87oVu3PLua4QCwTImvUQfg5iV4f23YCznMul7OS3arIJilWN
L80tML5mxeHmGTFUfS7uVUYwm7c+0jimf36vq834HDxqCllwuPwTj9YAGuIea+mc7mrb1YoJoykd
IzKf2arD0wXfdEoO18XSm5umRRS+GM2BrocKzL3r4H235eGwqCmFQsyMF2EwB0+TWEQa+1MJ2/Cy
e6qP8obfdlszySZtZq4Zpj0jgAE1AGi7v3hlrxXjWfOgiBaLqH+XZcGQKYxKmHMVjf96WcNadReO
eGXPPOCYM7TSeuEsbm8ltIc2VDVPx0N/sW1AgYVxjhf9aD03sYqOv/mnSel/RAnrLsExLXUTSR+F
ZME629AXW1YF7hvxEtQjcrkZsr2i+1EHZ1QlI1ZwbfzaXsEELe07Nt0S116eI7bJVocm903OixKF
om9wt7hHNP060eZ5388IY/nVllAWSyRu5vagKxeVXi5pXrhV4+QCsrvMmcWgumqgCCOpPt8+qT63
+HHgso6KzXHAQbivyf6UAoD/KuLM1++6kCN19nRrXCnByc7Qta8lgnYgUE5QUlIK14/vnT/zNgKz
6hrn7eBxE21SJl7CKfUeVhSQ7kSbHPwdDbxztm/6VifDHcrV+3iwBQFM6lkF4dl6DUqUf6Qyc6bQ
xDjFVrR/XqNlp4B3LT5mDUxZuC2zJ4VP2zISzNCdMtivUSegdE8xRYyn0M5qBPvUpmHCqNWA49xl
q2H9yhE6u6FPgCkLStA1Fmff257q9RxwVUKkO+c7uFm1sgVaEbl4YkwCPFemesuXyOXZ64fV6Tfm
mpltFzdIGXiXJCWf8ezT/YBZojfpZXV/bVvU5pQWIxmJZyGQLynDGW4FPc5WE07F7Fs/N9h0fN4E
mGhNkrZpeAVSPF+aVTqDrI3smlO0hVrDKptJgj/rT5bEY0S3gSw49LQNvO9DuLWEnyssEL8HLOMn
PsmirMrZyLjh122t1lGofzrSC7ZU72It4Pq/6DsDL3K3kXrYNUUBMbxd3oHx9QB6DoG0+PfoDOn9
g1/PzGPlbExJMV81hr3whUbpeBDfsFMtfuAtxOHZFleP89WIMMBpT4ouzCbC9IwJMZX81l41RJ+q
2Fu68QjUJ/8defs5RySfRwlEESDjz0L3kYrz6cRg11HvAbtZit2GpQwN7EyfOXu08BWxgZbWpLlS
EzAbmiq/1y18k8eOo5rmiJTpjAIizl+Sv9/VJZNXzIhrjQ3blzjB/zrev3P8G/RyBiUsR0H/8PlT
hmouLevkXnaspCpH0En91UUI7K1SPg4iyIi0NidzGqyOeiRSWjrgTKRJ/JwicrwyNntS062iT0Lg
QjdO5vWHBOgCVXNximzJLqXo1q0VQYE5s0Qnl/SxE/PRaepe8Aj5koEYCrl5SI6ARwMPw7Vuk69X
M8mLytkphuow+ZkdXFE9eW/A9sKbsfPMO4c6NrIhuOTtPi+9Nio1LvVgfTJy3CSvVUX68RM5TZpl
g7n+faCGmrFFxNQnNRP8vWfZjBS8qnEA+HAv+yjCJYdlZb8B5I3ri61CZMSHnXywUBvVD0ABlkmx
tGd45+BhjBH91VG4nwe3SMTCg3yWBIEvCyPyd3ixlRXvn4b9HcNWNC4gt8C7mMMvEszmlaxkQ1XX
WTx14+iWtMAitLpKGGRKELRAYnGjbqd0V6ICchudZyLkMquJfE/oSDEJbWDyIktNE44F+ZHw8dGy
kwufN7vHya+qrtGTXaWeafYX6bNxnFz45aG2ZCR1qZgoblOvzFZ6hpmyAbT5qQ9LqLzHDYV2XvGD
7tYCktcHe9cgcen7nTSVjxXMYe7U83rl9Gxxy/oOXaiDaC2gy8tCdWEqsq/OUgz31OUKnXWD5UGN
4DAFppZQrhnr2OIffrRVRTHFhoPeCU9DanendskqmDy56KdnS8R1bAUBS7tkbpl5POu2TWOIi8L3
w/egjLJfIMuTInPJdlFwrb5yYX1PS6ig/f2OhJ2Gr85Li+nNcibniG1cr2Y9mLKBX5iQ2F1xZRQZ
0mdDPz+XWBIq94tFMyz+f3TJpXSIqN8ILw77VWA3M7FOPOgdcCR8af6jomvbmWNM9lSo7I/Oi7Nu
jAaLz9lIr4rZt3DPAPPL7RzLdyVOI3wfOmlEf6fnilzk8iuUrzk1jHHGulCUmrocgzOvB/XLkLPb
TMjIS3uEvsDU7QOots/1abUhAjBqk2V+VfCXE/Jygb/WxMSesRgYCGLNBgWAAfaRWxAwvTrrx6sE
pgBjl/D2f2t6Odolyg9Nc9T9hDNOS2VcSejiEhR5pKODWkdEGLIdJeJCKOJY2xU8TtEThCxYYl7k
0r0gTyfJnP0f3iRPbxrTN90ageXiFatiClaPHGdKNzA/EoyDTzfWCv7kwqWikfSw5/hWafYOIkpb
668dSdHOUoyvkJPQ6ajZbiTw+YfXks/9qPDGDssd1CNHLzMYEGztO7fvfFFEtNN3ipwMlliFIys6
ywq68laSv+WKRVLB1k08+AZ12q0DixDjq1qMhxuzE6/4xJnLyZbDFxVgvrfptem8/dd/aSd6Mhz3
NJDjRu4WCiigYgag1Nd9tKWVWqxdI2gITAj/CIA6H4S4ZYspz8g+K1AKVGOQvp8AGtut6zsX+arQ
t1V2F3jEvdtGnTGktL09reMvgOW6VjgxrD5HkrdqTEOLG74DDUJVRoJhrHEmeNe7qpsCWkuJzQnU
VLLy6YhBMcCYfngwoPVPjgvvn1dpTMZuNtQsMTzmAU3KvJ+hdBG7q13WPozaMlhfUCylN/S7wfBw
MecqQTIVgKMwLL0h1bvzc54C3OxeoKO4jYOwbyzcJTshYjlK2f0gEFwGPGSzt/j9UiJNK/woa4W8
BY5+6QFlodxCUoy6ucK4Aav6Fpryf58eXwOm6uBIiswEsi236dEf9ZPEJQYyVL4uFIrwqG/6H5tw
2VpEIbtBP5uVVMt5tZma7G6q5CUYEE1SJ27MHXrASsO9+o8x2tN931NqNi2PGGQyG7ybCbu3PPcM
ZRirdsUmMXtvBLXWZkDhHn5A5vqWlnLD6qg3DO8MWXy9to6J2Wc+H6zstyO2tFkIWB8KTdAzCqLI
5Owv6LmLc5T8ZBl86NGFLVqmySxZOD1BuQ9q0zjqpuxQhvtftCxFyjSvK2UHrfxTdGZaysQKDELJ
YcszbmmVLU8a13jJY63NDP670YzidnOeCM7ZlbYOYMyq4UZ/OQG4RLmb3NFyPHmRrvRxmex1KcFB
UMXYCmiOeSGCjiBP3TkH1A82DJut0dR4OK7eFJF4qkMsmZICHGTG0GyUvG0gzzpRVOc76YG8bZ8a
RtBYgDwMRxkmiP9sC2puNntzO6YyKhCJATQn5dtmkTNTdNcDpvCS1s/K44ev2KKaT2sVPsNpAlo/
E8WYkYdIX4OMZv8I4CsajrXRFfhudFQNGDpv2yx0oPQWtlqxRkEkKElOkLZfsQwv4jkfbaWEhaAY
62PvIp0Khmn1gZ96UxV4VipWXsvtuD5OM/6tRZGINrwgI6wb9fF8qSJeSdv5CLhdZyvqvr701IoW
coIxL4uSgYwj75uFYkWr8m2I2lmzuhw+Cs5775dYSdfI/BtSYBr11eqdmpdECR6kcNWx/Z1Lmn4U
Q5rGqrlNSQ2cb4E8zT8xKrtUcHPfPD0FVLkICFZKCHfNRAKCSj9YxezYXt1SbqYU9Ci1EB2MXu4d
nFFRLd2r0JPWEt30oLaVbZLWPOMxICKsDDKQ5pem+1GPTx/E4F5/OUCD2hHBfDz/HwmCceNFkRLY
FeuIPhnJvlhFqx0tnzW+svqzvhz7BjXOQN0aSF8o4VsX74n0AEoimK29KI0D3h60dKazdiNlRsL7
1HirmyVmWP2cMWbhVPcgPUU68yCEVadLaQcg+4KWPMtrfQVOwZcy+DXzpWhfd8Z+NTKXcIRfqRXB
TTCN3QNUGM9n5RCyrR3Iy9WbCE2nnGX7LWQBl8tTDOlVcRfSKNsmVgEBufVaqzFkyzIIRrsAbNuE
zJA9dqA2iFRcRbMsWwUtb/A9kAecLRHKsP4s1hQA8JXeHMTjpJBU5cTYpRB7pHt31sWLN9G12mcY
gIGmMfp9aJx2rKJK48ykobnffhGOKhUG4WbpWX/DAQpmv9QYuhIxzlqYVATBvpxvYJteTDJ/cHqy
7qV5CmyU+3dfI56CAIYQvvmmBp7QXW9GLTBS9xmWvfRjK3KMgJc4SBBzLrNUtScY86dfXfIECFug
uc7FiLEolRUSF+PNjamG6xyj+ObvCU5VYdpqjrC8s8KK9NHfS4eyWGIq/phY+72GzZrlLDPiEL2F
Bz67o4fvdviRA+K+6OgcINe5QAmg8XST+O3bBBkwNxoMrkiJjJZ/38G9dvu0Ip7AI1n97aaqAgwP
J9tiXUuW6AI8loxI6SIiboyVQEtoWoRfaRoMgi9jOgJ4+jAncwvsA/vFYif/gHWhys46V1QtX5CL
GSWbdTWIVijP/mROozlcNqfGwGwe9TbuyDM+pd9D526KnDFSaoPTIx5yyYOWzz5gLXdHwTS6o08H
2C/lw85WyM6VffJ8br7C7t9qETx4E/tLWduxggnJiY0cnRVEdJrwTk/Cyrv2jF0nHYi+poy18zlQ
8wdpck+p3AITs2aSd3q08gMTaz683BGh/X+Ne/tcFod/RRERzfGUxWAvIfrtw97cfz3pZqdE54VJ
XHHbCRe5edq8AeRqm5VNwpH0iT/vmt09Hq/5WuDvljcOZgYLDx91qLvD+mAvjTKMmNWBvtZ8PzDY
5CXWfd3a16vIJUbbBRFHyloMIITQO/nq0ZLslZ6pF9TLb3DmmEgju3VceQC5PaHDVbXfobPyZqmA
RFz20r2vHlQEpIJDfo82IdMpM3XUh+gzu1B7CTOhD2FROxVRmciFdDZFc2mnidxthat9ntK/Mm2f
QRLu8kNeAC5jsPe8hpOS+8vJCOyVjtuql8rYVyW/CByndst9cXoY+YCqYtKYS6vQtuBaPL89QwA+
wXOhB26Snyga2FOF8WIjJpOhw/Yx/UaeQilW/27Mh8PwvRWcJseSAH2JcRm98qtDkSESkSUQRFaH
YCpn/CYrIatFCusZQMgqZTBUpgPdempULrilW320fIyULCLxz9xzOUqvTGYyuaE+eCBxW1YpMA9j
a+BjdY6lVtihb3PSl2mOvQrYLdhwwU1lNEhO3vSN+NclLf0Mmc/8t+bd8SC0KqKoMLMqK8USDV3/
n5Y1zbIyxEv7dwcJpzKpthTpPi0yVAD45NwI0qu1kMJGedcLLBAlspVyImRAO7/SwYH1Mpcf3XVa
b2ZVtc9P7sgk1QSw2VvPiUWD5ANquJ/x0pMDNX009t+pJI6eaE2dNaov9CTSYofHYGHntcsu6HXb
LoWA1fjWkmRIMUg5ASViDnP+xNSoGG12P//dNUl5VmN5/5w29OPFB7mKar6Ajlx0cBRQu/8K8qzC
c1x0+soe5mrL3vofNkeNTFEW3oGMXvkj2xcISwjwzgB8t3azucQEPDZXm93MO1IqLRSooQRmBczY
HUXQCZl3LLWNbGH5dmyS3VJvMjf2OpkD24FLFGWjWf3z5tqrM+FYQZiuHC1oVLFA5fg0FJc5Ci2o
5d9cffZB0p2+0r7RHMgoCNb4nDlS3XU1MSwI8RVFpFe7FFJBp/ATf/mUSi2jkLQvX7A8P5Dodnob
62MTh3Y8aqE52gBIBrJGTSoIAFRhKmGXYM7N7L9S6Bumw0PjAnDG9fptUIxqtOB2j06VI/gvSiAL
QBIwEOktnLsMTA5E5u7HGwR/o3eIYPLeOpLn6521QQsCd/sFpa+L1xFclpSRym1gnTSbxMLjiNlL
U8hOOC4iNKTKW78/8hFbRKG9bfQ4n70MKGC064Z9hunAPn+cJBFkz2wTSAlvtlwd9TWqZ1RJ/D4y
wSdjI2zUey03CJDFdEd65UPZehzP7VlLKL0C5sbrtYEe5ZYeBFL0sEDYaVMtIZsGMBWkBszplDq2
0iexF8jOBzj8TFYX1c7wvVPkM100arJ1cQ2tytjIPlE9Z16JsaSPGr03QWzooDOdsdrssmF+1GoD
2x3sqlCC1ZAjx5htNE/R7lg4yteRdh8Hle3oaRyN4fLjT34SXxKJRxJ+6lhosVXdth4LmQpkDz/z
LzYW+u+xVRpKx1JyfE3z0D9SMjMOXRnkuScqGXuW6ntNZ2EyYpCKzpl/JwCyGaeswXY89lp4rsIu
3mpblaTXzXFo5Y38LPbI5yGyDRymUfiaI9hPapiKgxsjdxgIqie6waEFpRnC5qXvmxqdp6gwBzTM
mGXOsfzEwNZCXBaAU8nC7y+TB8Iu5LGp1uypQUrZ2tbpxV20HFu49XJEbEdSOmE0UQ+YRRcrvKQp
WHT/WjoI4sOiWnPcr6BxNcpfURCnXEcAUNNoGR1cFCpWJsMqXeU2pXg9FHgCkpYparUe4e6gtCOX
f13Shdj3rRTkveJ/dLuVy8ffJT4AzBRxBlAJslkC0/VGSyku5cpSKtHGM8namMOmRg2sYQTPMSVP
JtSJrFsdUO42ZSSx2D9Qa90uyMAfNtPedWm2mx32y2BwULyUwgiN1tLcBzlZIiGlhbDQui+b/fmH
5g3Fj1Y42brI8IeahKtxfpCQ2e6wHtNoV8ArXTbfPm1MoQP33UyYnjDpRPfiolzHB9WYWJHvceKq
g3H9x+T+/2Zr9+vuPl5+nlxlgRF0BSwB01eYoRsml8FfuW1VBmSv8zwOMmx/qDvDWHSWMM8UCa9h
NC5j6OrJcBXYcuWcezQKQJS6gKtJZgy+aiqmC1QX3pfiUwwYHDaBcPd+tYLYm4asJank/cItfNaE
i9BwXZyohHbay501AK2jsIFynDRoA5FFaI/uwkZKBPYLloIurArkU5S/EzBlTZU9rOBKUq9LzUi5
uDUvKLbt7YQv1eW/0X60ncQRjCVq98D/OTpNV22Xk9Ftj/6PQGMPiA7+tii/r04ZwxXNEuHiwc2n
q+ruYorbNF7JxJW85MerJ5X2mKeyP5JbDiA2f1tV1ajurI2hYEcgeMAPYcx9tblMmWTbpLqL/pmt
uUzaDlOcAOkL4z7Uqhclo2LVgNLUojFs93Hm5waCMeRIh1lVPl/B4m8m9o3511Xea3EmSszAGpP5
VbqgJtGO5P3ewTZBdU3Ahfx/bzgnJHWPwwyhXk0V/anW36TNV6YJ5wBReMp9x/y5vH7XVhvpoD+9
WeB9xnzCixBUw8ulYj3weHEsza1C44dIeJycovmWflbPU9uXcbU7frBlWmmraivHZhifBb6S1/MP
keaPxofxYWGBTQ2aSXv9lYdPDoW8kOkzva7qZAAOLhkRUFvEzFVb0YeXQuLMrnqiDTNydau7BWeG
rJkmf/Vsdfx5mxzpaxAWBkn6xWBqiOBPID5aVBsa7KwGA6IaWQmgN5B3LqOQe5llJsAm+cWRTORp
Qw/UbRCGPz7Jo/f+k8XC7vvdxVPSsI0Z8xkmLVjstYSYb8umdG7yCDt411Sxb76DQyDf0vCJzYPD
GQ+VDONVV2h2AJEpmXrkHLb7EdBV9acEhv8pyGfcgVdBNjf+EK8JZXvItd6NLNPZdr5CHQlnTUrM
er8V2hOAhM9ru4YwkhCBv/uc/Pukwjqg2baus4Hr4JHMHAjR6mFsQ1C64e1LaXxu5Z3V6x6JT5rS
da0oqf8ijMdLGxX5Vm36UO8svcNkFmZWVX2dAOnSai/9e6Gj6lklfjoAFTPn5iV6tz0D6KjVVq7u
XwsAEejk3EnX5L7mNUeekdntW1DObdBpycL6A2qSOHXdf7HuT0AfTzYakvhBM3pOz0vQ3rrRmtEV
3ctBzI5qtNohIa2Aakpfms2xrzqAU6+pE5ZTthu+ifIEgr68QHM98Wg5gWP1i+lg9YNhgQ8Oqj9E
WH1kVkFyHq7iV3aaue2HdnBYF3njVGo8lPBAf/Mp2yYk2M/5ROtnTCx9yMbRHaYMh3HKskNpo1Js
NQ1Do6to82YShBc/i0+4sv3m/yarr5YjfdXFMBmRywgNZX9LvM4IwPlzpV3f1wM7QvSdarS4oN15
g6ngMhv9eHLd7R6zU6uIZ7F6I0F6nbQSR2/vtNdxj3ivKUpb1jPFoFClMYASpRe4Bdae7TCHsZkN
xZFN7GfAM2Mix5GQXS09MjyMgUxYW2nyL3k9l1IhLdiupXPa+T2Sn/L4QxiwrEn4EO6xOngvgO+1
r8ClD+PtAaFJwsJ9AIGD4QfKh4ZqyEdhHJi2jNl3+OsV/0pED2TtaF212V65Y6/O00m2snNThikL
A71P0i7rW2im2ujGBPr7xap2iKl9veOyLqVsUJfUC06H+vsdyoPAGKRAyrQsgT6Imokda/8EEL7S
xXwF1UKVBB9awylNnXs/BzUxxfvZ4VB7CcIeGVk2Pn7sDVRLG1/r7D++u6tmrnUkwuhwC2t4khOm
ke2ER8oEST2szf7RSCaxW7Yg0xePsDroPwMK6NdJgOjBwnB/ii760KiH8zFdEZ60iCZy2NvQxpQC
L9mGdDXEEA5XaF7t+MzzOh8N9VbQaO0K7GKzVBsIIdtIDPbBj2sbYYX27hh0NbU41EPWh7HT/XQ0
57t37tbvpYIyMEdnRIGmGbwziAoQ8LwwNIlONRbedCS2P++QPlBH4o64ZGEANo2oBRZqvEdTOYKI
cNuirHYjT76q0rNh24F+OJ4QXr1k18Rbbd7Y6p8MBJ5+WGBWQtPmwI0bqysF/95QjfGdEciTZO/5
irVnGk48+AWBolUCfyDtq1TKG8LYn2oYDfewZ8tN9WUSAlltGwD7MW1W/RbLHDEAnT4tARPpYliY
4bXvS0zpWv0GkrTwdIN5ShEovA9nLI13ORNlNe51/JLb5x+/hFGXeyyAYq6Ow0zmfoXEq2S5/WqQ
MSctU1KDscIRVKpJtfPNMhKqP6uYHkmM6SXUl8iI8Ni+vRXSmhUxKRpKlEzv6liSDBfZHHmT9q7k
PoTdwaGpin5ZdDu8DTMfuzKv5BskRNaUiWJJLT8XvdnEZWwxnqhqtdkEyx+L94W87tLw6hi33H33
EUMmhGYpRI03AyMhPjXfT2eSHXzAWUlBsQ+N1CM3/8Vk08fiedyIlvxMO27+ovDBVcmMqsHgRdgC
RvgmUO0Rxv1Oj12VfvoW+ZakbbZDm/Blo18Km7psHENznt89kfPqsm5NSICBfYERCYJBRWF4dinI
6foz5+hHsvKXZUwf/de4UKMmfb6pKzL/w3g5cWygOceL6jZS5VfYOucVdmCvLfG/Mehf4+kO/bei
NTIz63tC1Yvs78yJopQurHSSOLQV2xWNt83phK7QzcoBKjN1gevu61DMCRAXGfZJIQZa522Qzrqx
oPH3XMNWu5M6t2+HHTov96d/YKN6qU8H9BSS45kSz7ZtLpAW6TsuVG20GBj5YsRvIX+bvZHRJR2p
kR9e3TR3fnLWkKqxyuLvBDZGG7A3VBXDfi+FQGYsX4Kgf1ti0Mw8nbosgog+Hprgw7SdCmDtsw5F
772RKUrLd6QUUzNFnfzvUE9vq2kMNu+c2u3s2G5zYFyX6zyNRGDn2kMSNmwmr/ndHf0ivJYn4jVc
CQzp03Y+B05blMhFQrjeXVh8bGB5LUbYffUhRT+/R5DNvYd0yNVOS56DF+nOgxy7PGcXBs5Lgraa
I8lpQxQyXNm/vxNqtLN1bRuZ49lNZmY70CHsUCEQWn3tpL1ygP7T39OJ1L813Jj1ln9IXLtMqNw5
qNKUiN3ZNUSJnLNOGdLFwy9jQFVHE/UFnnnoYbe7bTdq2TRFW/n66/nqSf9nHNl0tpi3JJ2jxWDg
dchjAKNhYBl4XZX2LRRKtsEBpwNWOaiwuxr7R6Kgd1dqJD6sRB+qOyo/dt5BwG3SIJttkXZyllaz
1+cIULiJ3CFzlRyhS4OSySJbBSazWJhCilZB+vEHUet6H7UQeEVxPE98CkrM4Ejqsf4eKANDb2Tj
Rn9mI9SN81ShfKYmp0Cw78yybWbrY8luBvuLyEsN2jwFnK7POuerZuwNANG/5a2mX5Z9xQTF0+py
uqbMGHJUhl8WpWZNSP3V9Tmgve0wUNhqknOmJb1f+f7umWT0dAKnlpYmGRrU7l7LdeFSn5p0OlTF
qtVbtIJdJuz3w3aWmODEdtQtBJuYxo2yX2gFt8cWxK8IyY7WrpfMV/la+AlVCCYeBJ4Jn1a5x8QE
ObZ5m+LjK2bKHPK/jJTDig/Z6uJoB8eGcwP53ekHzYrUDVZ2flG250+yBPyOg++gbC6zW/UqIMuJ
92/hnEKPDLSTFPqF6G0q9AWAD2q7qlVbI+znqO/jmETCb++hrMQ4GZtVX33QIbHL5O6J46JBC9jZ
jpTYXc6PiesZJcGzb3oXk0QkDiUJhAmaJj7bv9Zs/oxB7BFzngYK6QTKbsxs5t8dTFbPpg4hhP2I
aDPOidGYz5lzBU3QK942Y+jc9Car8NoY2vj7aaqO3VZkOJCfYRFcYyo7B846QPZmRv7LijMOnzHr
pUvdcVyu+CwK502DvouBrd7ohUEMagfTNQ9twjguFbQKmV6N1g/B0xpTyR7DeWhnKERWq5tsLoTz
qwxPnC1Xrt8Q1vSUu3rFFgj7cJGTVLYb/aE17OTV5zxnhwNsKtq+pE62mwiKU1Lofwp90kBV0qFy
aBW5W9qL3o8ubWS6atB0OMbVPZavBUC9NhilFjrsx8H0ganVR2ZezDwQadYzvcFoPXHLYYFYlNAH
4h5iVJ+0fToM/YI46ghpv8vR2/FvcSp0ZjAHTbeXaNg6JxZ7QfWNgOvr1I6EI19+JRkD97UnWAiI
hd/mVU+mz2QXGeFC6Do/OCuyio06a3Bz6UORCcoCurzDyt4J6fhAckbNThiqxP1NONNheUvrc91Z
yt8npgSTJmIkrzz/B9++kE0cP7MHYl/AYy1Xk5ns33JkyqtFcVuGuiVrbhSozZ4BJQNtGywzsWl7
Fhk8N8ZsLJYePPSPODbyS/XyJ8I8HoMP6c7i9tkJGDklI23ibLAXEdwikz2y24zFg+/WtqgtIALb
h1oZazabDl3T8HHgvvNAHaWVIbSCEXjSUehxtSblKNw/vV2YtBIn7FZq8kcy4Zryn1l3oUwUVfwq
b/eJjRzsYg+G1PyPunEGiKHXbDR0apfpXg9gDysKr7mM3/klfjJHJxmv+/S2/Pu481C5/4GRIq2K
bfrats/mEk6wnhf9ZK+ZIzFkdNP3kcGq7S6dYdoGX7RbrQAFUtohU1Zg7E+dEIA//dL7QeY2nj69
xOHg7ZtJ8iVvamGWB2dZZ9zJ0kNYfBnus/MHr7ow+kDL4RoBWQCx62ageb7vDONIPDZXZbZXeydu
Rtf66xJkRSb5bcaqkt8EUJIM7MfcJg9S+QqSSKvgaoYowFYKmhmc3BMwJhd5G+nOCEg0hWqIQytC
yDTcqDTtBLVU3WYN46S9hTIMrq1pjXZQ/FOGAr0NS4fdtCwxSb2FikJiQM2JGAxXzyoZeXmkU++R
/S19tY9qtuT8u2etuaxKvn0rL6DdE/Iiy3ie5liTObh/CWlZacEb2n05SuwplWrDyw4B5wvn94rk
CinjxvoWQurcLH+7cYLL9RAZQyZ72k+nW+jwAsPHq4MNC/hda5MS32tCH+NqYUnAJJohujiXV6Ae
nv9Z3XhC3sxk04SW8OSWEakDPPISd8ZXiW8qWbWbtQZeEqTIkaOQUMvfPwOlvfk8bNiCu3ki+iVs
hVDMA6BrbyVgGub98D6Opx5QI59I7BcfdGB98BR+D/9EAv79G6JxAm8mhJ0qhxE9qGxLJ8HRE9UB
+97u7xfbs3TCCnepmnMOl1dE5G2MDR/msc5H6rUMhUPGNE81Bs5kZEkDpEE4zmIAqQp3pAE3ShIT
Njw4CZ8EEN61kc/MQ7c6vQii4bUBskXM+7lY1FGgkrALvt3xrZKHL5NQOyMadu7PESgUX0Us4sI3
EX4WYyLarasoQ+ybQiqpaN4D2/NiVX4+dXwp6MwPt5MDJ+kM3p/VceMI31rAiaMwo1jy8LdaKW2L
hVRigCs59VL3ykGzGeVsDnZ0zToHuRIMRd3Wji4H2l6gkvfqhm/1XwERAbLAaEES2O+RHVohjn8T
A2I5qBVScFtZsHeYviCDTxOH5ItVAOxfBWJuwLet73HZQDc3TblsDPUTqE+s6bRSqRb62pUawnt1
hLQmvS9qCIw0G4zH3RfP7X/TkSZGLYX00WdIHZTVQKxKdmBvDMc5zsQeK54tQPGHz7g4yPSQfDp8
vFRU4Vf/TztD5sKxGtEc0lnU77cQcgeP5LJV1KQ06GDdLuGZUWaZFHoMDm20lPKM2asccn2snSvR
8CUtMODX1/LayeEtdB2uBkq1kgzO6zCugv6y3wABiGxmZghady2cl0fcLWY7N1rS40TRLfcEMJCA
1T0c3SctdmoLh9RZWQkjbep1nx98vyeoYiqoFdfV0MmGZtmQCnIz5oy/Jiux2v4ZwN0Vmj4sv7i+
RzYlETbjZLqb9s5XA28Tpd19L1qTUxkXT8MFUR1fAFYSYzBJd9l2HSRxApNqBLYFVmBxTCUdYe/c
QgJ/YQjLUj0Ze34PZMx5McjBjLVjnkUx1/f0CgH7flVkoFSAl5KowaqwKb1NgsIsqRcKA2lbE9JH
fwkDNhcdx1PREpgW1xey7EFX3scXlrTQ7ZGNmT461yGsmA5lJOBHG7+03/xsbkC8F34KAh2pls8p
HA+0pNaT93oQeRycDYDYXk5cb+fF7lbB5L0UQ8TkMNtqkGX+qBIVf03iZKPYJ3JHR3DKkmQ/epax
hYh6KP729/r5Eoa/0HPDGBswlMquebHNtP3I6UxCFE/kkwyDbLzqN+C5tEnzMQK0Pn7WNzsX8Xpd
IXe08e1l3JWhoVSAY5K+WuocEkDEmpOmFaMVOQhFQEIIYgbFFiZmH49TmN4jC4ijVIpFEHMolqzh
Knj/SpXYzhJ3sdPa1QhRoZ8sHZ2XD8vOa5TEvorTBsCZjKRmtOEshM6kE84utH3il+cOe8/1LkgV
xxAOpX2ORUVWpjfXARunP0EMX5ZJOBgxOdE9GtrRYJcbdabxLeG7LpSMiAnyNcmeMHyh6yxqra1Z
vzPY11L0Qj2oQ+8BvWegOU324E9P0NaVIOdh9FwLmm1wWWtFj9nmWZwvK7OhMr84dnVp6eBU2uyi
COwRZOHokJtfyZz0/8m/nLBP/5EzRhBxwkIeaGZm8Fbg/2bjwT1ZAG2vVZ3jVxA4XyPns4/rC5hS
LfsqWC4xczgeDFkkNs/mmG7AfEHUErpptnd6wGLHU+cXUmFoxWp+pHWnHaNuoYsaYYYiaaxcHuAK
EzwxcY4t8qLCHOh654u56oKaQ6GdbRnyx9diLRy8aA+oBW54llk3ykEWg/04CKRDDLwKVUCPKH/n
w6Vbdr6l5GUalVscOa7SQjK4ZKUlGiI8tRm3253TblFzi2s61vO2TiTjkoQSg8Ad+Tpdj/6XopGl
8d9s8p3i1dZ9c8JSGpPMmGna790mmHXHMK3nNv+FFDdZStYykkgGpAaV5mt6weUexx9CwJnXHQuW
iKJ/PgIm10jakUdAIo7CzJTMynod0bzelrVwhXXmVFzCAi5YP3Kul5p1ymO6yRoXPJumiwkRyigz
dGbhYCwpJZLIMci9hFw99oPJ3PHz6vVUX6HxNHTza+xYGSq+PK0VuDZF2BVj39hLFXTFkn9iZqLn
aPGDqhmpKGuNA2SvUKVQVdJxNOuMq9JYHZYlO65Odi86E0d5oAk/ndBrdgNWunVfHfardLtVIdyL
fNTaAh9xb2V9RjWZjWZtIVpgBHf/xqhDDmCOb2t/n43rAgyjgMama7H1aAukpxJvlvki6nyIckJR
BDXovjOlpgZJxU7Yn9tgyJAUVGCWjingRYnuodzT4WklwoAlUb3Rjht9cpa5qgKDvU9oyTlq5oDb
cmWqpGhzAPXbH9Ab1cXPh5LacthDnVzrCATeCrNsLEDtK3EDr51mmOt7H2VxTlLJKtCXCtG2SGAW
RUQpW2eY7GrL7y3CoqenEEmAHFHo6utoH42smZpQs/bko+f59JcijvLdbOD5pgmUEMKnM0ctvwgq
Lm0NsxHBZfmD/kW2dvOvLd/CDh+UX71ncErZziq0VPVvbKYadEivlTv//s9Luf4x9D6ylrEr7Zi+
p1W8nwdMgJ10M5oyxpvHZZNjvxlhG/SBlW4cpP92uR0DCf/daT3tAb7NVupzQQdOvHMkDSP9rBPq
IP76hkFDMa+B79G8sJNHNxCaAXbTl7tbODKQYn2FBgpoOLD4PKKOg/dovkr9M0XVoQr0M+BeDxRS
Td12cxtTkbUcSw79y2F+ihbl5G9dd8OYH+g0/21ZhIpp+PSfkSnOfc6WlfzQLz2oHNZvtY7ausW9
tBKj35TgJqwcdI9Tc4ANVYtsJFONtCPNgZM3pXvfgFLHV4ESkXDDkF+QrVA6xUUvVWV01Seta85Q
X1GftZ30W4Vzy8HqewuYesneAjnMcGkdAjIgf9h5zzZ6lnQmAzt7GOTUn9g4cl7tFvb1+lWsVC7M
o6QRwdZnJIX1gXb6HGFBaFYP+egKPBu+/6mujB2DhzHGpQhHsGaUOF4oGdoE4f30FSivGkyfTkbQ
zgzGx19r85rha/l1kJlLqurqa5XMOuVgwjLlk/r4CtcfQkwVMVTdzqkiknJKH5akQik/a5MOS4G6
agslG2bLqxvZPuBy8rlEFZzZFgAEV4nRJ04WpnyG/jb+bCgnqYJpt1y2kbiPq88WN/bcn9wJVfuu
QANJ4dkDbkSnYDFH4zdgAM7Zb1tGKxgao3B0gZvJntP5RHz2hj4+TF0NcsdeY+rSAxSChFyAlGVw
zuM/Re7M9/kNqRg4E8/tWRJVglwYy2TQcCcb/R88HaDh+m/38fbGumtkSL1nuxLC8CMGodvfwaGV
fPUMndaoAhyRoky12gEtrHU3wPxtH+9S3P5JTZw4h0HV99/WIh2RifUdFYG6Ku+keV2uUK102x5B
Y4xl7IZ3ahB+M5f/omOvkj9mGKrPQRP9x9Qg8UB0Hf8ApxeHp73p/HCm+Uc7KvLaYCutdXxNpeW/
/gKYJGNU2Mjn2orNX3nf8/V8RIVIdwwFpl8IRxMVP2PbP2jIcpKG+BCFYDlJJ0dFFOVx8OUulFGq
AsZw39Zlffd+wyJLP0kCIYFudxksW+Ju+7FLtubltx15FY+AQFQ/dMpim/C59eUPB0a1ZKf/QSHu
0+qIMhcEbuMi02Q/j45AR6CzOGvkzr1E/vtWir26qDUKZreW3yDFSwicpar/6FMvZ3YhsQnkPnyl
5wE24NzOMDQf1qrJZRtdl0+0sWrKbTkRtfbV5iwZJoaJYOF0yc24JX2u6RXM7hPX5sx1dgZJH9tG
UYZUClhfataoXcmwstS5ZUOvIJzj2ge/QHu4VOTQJvq/2UU08cZqgMO/yyWg00VZGWz2fIx6kEK1
693VVEZ2lDCh9yNowmzssBgnVXL6mjXibbqhv4FcwEEolYZIIVfwV1ov1u7Hz4zXkcwi+3i3B2Lz
AxTpmk6UexHqHVf2xgWG5aWAa8gOUYNJVvpxD/4aXI6+8tH6w8Dgy/n2YzdOcD8Qu95ihMdHHgr8
AnqdT7tteks0j0e8TWufqzje+yok9Yx+ldNwky9joME0AOhTVyIGS2tmXlzLXO4EtMba9fZFKBmB
vbo/mkFhhIiYCcYnixYkAQq9MFGx1MfTpvNl0Tpx75WIB3SnbSS9oVIu3jrzcpwQuk2A1hKjnR/V
i/E8V3aTSmOmE8XXhlMKuRrM7HXamU4S6du3Ue3bwsbXJ3WaMYtckcE9bCdue3/KAJhUMY6/P54M
E1xNCC+DD6BFuSuc36wcaPQx7bik9/PrA/H9XQuNifYRj0AvZUlAaUWFCD7DHmRo8w21R3Dvlyk6
qpnCtvXkbmwHJvVPL0RScCDXM4sUCGlVLqulw/GQ4kQuTufiyAIiweAR3VuhmDpWDYX+xXqWVbcv
nvAz/LgtVLrOI2ErIoR/1TFx2oGL3oTidEu+0+WP2/+aniKiczvGUZen/L9yB2JJ11LwDcpmfa4Q
BStI30iWjZl8rQUu6HSDe+TcUFgA8fJ1XVV5rjOYnPM4jTfjXRI6TiN7nMPZkQsYtrOtfFBgmJFA
XyCvafOh7gYbxy3bLbL0r1XgdnPL5pS9P23kLK1XOyZvTlbaB+iE0lvybrmmmckoFshArQKutRsY
4mn6LgNV5Ojez7SZuuznlx8ggkAxWBkGoax3c3bIjc7zbyFRKCSqiZZVKg9PtyHglwbCaTlh2+ip
jbcKOis6xFMQVO+kZvsMlG+FyQMwm4xwIjlLwEEXVHsFfxhqwbqC7MgdL049pwKZCHFtmEUCYtFP
dzNx1SLIffIbiBk7eu+XVAIa3qQmTgSxFl2ShCQeuVv8r7EDrpdeaC7aJhEi7MKopUIlmywoo1dK
sT3wiNjDDDbxU/0ni/zI6m4Vy7h3QIc679Xy49zcCkxz06cWSrHbhziT92QjrZBEEcl7TkbEd7xJ
CtFysH1WaqLt3UFijs20+0LUcrWXwiwwQmoM638NaDB8//hklJBx1ZtpULLU0fzy5M6fjFCKJ6WB
7l6zT2mRRbuRPLNO7t67cms6BjCUrOmwEEyU+/otk0yMj9v+MiVBtm18EfrpmEqHs8VnOEmce00J
d50yOH8+14iNrbbkmbV7U7sQZWazoTyqQxAsSjW1HUQTfnEg68UczYxinl9uziQhL/oiHiZceYRp
g70nUlk/jiEHlkwfylULK8jSUMUGj8Mbw4hC6plMRqq3TZZ05MtLmalqimkYzRd23CftLTHjQm0G
3PeNG3cSXNI8sHZGWJRLDwsLS3MFVldOpVMpvzir2BmYCj8RFQrGJgHn+iWm0fbNHdzvjBpYi4vL
tlboboeLWR/2vJ2wSmFMODtw9S92opF+hWVcjcoTw4sGc1jUxU93UlLBFaMKvf5G2AU4BmyZ/gQO
RngCaD/q5xJvgCYbtBVdWd8tAirfpSJNivoJGQFuUukJ6nmYX19jdJ6UX3Qt7mzSrDTLzCuA/dAo
XZZuciLE0Ic9cm6pl7K0VC39EWyqxzfYh/KbJ9ID6TYP8bftEFBB9IamfNPSetdofLAZqlyrO051
SmisaNBschpt8ZQeUolW94pWOB9hDYlKvogaGe5p1r5aWzQBi1nAu6uEcy+iIQYE5/fe73qq5PxV
x+ttBeEDu4m9BkcwC9LrlHhtsFZE3EQQAPOU7A8xbVxb4WNWuE8TsljJjvatQQoXqXB1yLdPEDrL
2wRI0u3H5vhh1iZ9GF/XgrFSnrD34Ce53yDUOdjyChTOW9Zf2bK+5TD1csJSNGxOsXmZ2m/NGC1d
rxLo8C6r7H1a4h19BRcnd5214V+VChdoervVVYUUKicZK6CM7sEHOpoXtb45VNFn3ISxDyEvbBmA
tw/Ey8wb+E5aRrIl6PUNTo1z5De9ssb6PZV9tpXIjcYfl8zPGuvTWeKMygl8076VkMCtzZaanyoH
64A03jIIUKcrlMMlG4DOmoHo4CwhBzSULNN/3yYZZYdkejf/WoTDzSBZmwTDbMoXIGJ+5v5hbC5S
3QexgkBWnAStKGKqV+k9Gq2yEh4DcdeCRJKnf3qxv0GGxT79YedQEuFvXipUcx9/mmmJezPrm/d3
Pgzt1BaGDU2QAQdNw9fmjVc6ArhMJMf7el3EhiqBxm82xqqLrFbBjLD7+ZdjAErDkD9yd/Y7ZzBa
tuBQOujIibMCLCbSFTJt7J//jg42iUYyFCHcBTrO+dIj/1b+CQbrbaPDTLBSlHXNtteOhOJimK+M
VK8NuUtfxtfqSkqJnNRjzULy+w50iLWg5t8joTdI/shEukSQjc+sTDtFNrWqofv+IvoYsNgFuiHS
B2Jv1d4NoUmXwDKvLDklgeLQKuB9bboG7ElSybasggMxzT3cntFIheQy1Y7Vz/scc4rYqebU05OY
8iCohljiX63iL/AB1pF1kkELdJSJ1yGfxL3UtrbUByYjvVJQtSUkF+ymLGNqcmDOUcaEXG2RcLcx
aUt9/mVslOfcAtqmsFQ+JZOutsFe0Cm7CndMXrAvhYX2UEINvVoj9/aaDp7J2g9OJ5iPGd1v66Qo
0PGCLHNhSji+1QrkPQO4/9pafNBVod3ObFEd8qzft2X/DL0Pe6svlTMywRaV6OvPmJ7+RpTYZQGf
rYuc8hg4b/iySgotfkA1/5ZaBU58VMFxuxaApUMktfgfIk8E77U9m6dlOXprdGhgil6SCdMsUcW/
8vDUhhMmj3yJzsQvM8MY40IfF8vVm1/dOB/BtBpydki0Qy6DQIswyxGBOTL5vs+qHSJybjtZJxvE
PNv676Rxe/6PHxZZNEthxh2NiVMjLCI4YUYJqkxf3yBN0aXa/cGYW7k4vhIQgk85On57OAQ08WC+
kTOJvnBlEL8d8ODg4fMIdxEN5pIWdgDMGmWhCEAnY/ovVTYqhnDd65QXnI0SJcidwa0Zd/ZwQpAT
BOUd/ITgHzO9eE/qprlAO6UoKuV5GGnF7A5KMC1PHsRDVhWpCO65MDhjEyASwQ/0EcADu2P1nJeU
bFFLCJ1mlIO8w9be4sD55CTxXJZHRKoOodg3riFWr59jZaEmBaI7ygwHMx+0HUgAbfdGrRITcjZT
MEKnOA/47g716OYGek1KM9PyuiqUIE1jjASCtE1WNEp1iRT10yigWxZT+UiO41iDYUWKnMJM02JN
vSEdsLxo5BahFfDX9eTgJiPlOgQqBB1GHi/T8FX0uOGVO2raV0EOBikAKi999JZyEIU819wpPghl
eO8LcsYCwvWDwv07ltQHLfQvZ3pl1yegkoCZ/2umROtL7zdi/US7mVMA/tIcQoWnUp9qGBwa8ISD
AYpkP3c0dWQM+mJzWHv0QASLIfSNFkF9oVXpPgV3da9+RqXoDqsqs/j3LZvIVlPS/uWNZcBnUN3x
FKMc9DpRPiGMX2GNfgF2BXLJFZ+XcIVZ4nDOvC0ziFPPyDrN8mPgJRWhEsUbN96IS13wYKeeTJdk
55YkxkD+DuHyald6Ac2SguZd0phOO9lenVkVHVwqKeyEzvacwzG12fIxiAovXveHaw3dcMke5ZVR
WE3vO2TmaTsHEdmXedEVNHK42I2wi1XpUbyqXZH4iuVBeuXXflI4nWwhZFdXZIfxveZp45nxqnw7
bF9JDW4CPNvTZ0bTI8nM5FCCuB416GlcdSapfNfj4D4hUJ1NrLF3dUqiTxPuvwHx9taOJ6s+NMTq
wrpnqPUtf7e4SMRJdh72mq+1pOr8hf9AttjRqI2YeDtLXaZ5f521D/PbHGvtV+mcyL/JQCcI3h1j
azFfIHIbR7TEgr6/vQfKGkyuZ3i1IyTV18ujqegKPCZ99Xnm7CKyyhJJvLaQe84co1QAeJH0C8hX
rMobE4ppLJ+0BZH/HmRosat2Rei9ma+NMU+8IpYxEYK/1poRwdet5oyAfURy0eOdZZd2zXhEwuhj
UPVEubJty1PRPsghL8r11+56u46V4BgsGw0uFjEJgAKuugwTzCjfd5mnjZqPkF22nT+KXSWXLmzB
a240kLW9uBKfxqm3xozYkhyRS0LFtlxQI8k49/0M+HgmkIJ3j6n/ZQpbadaz5mQu/ikTnzkFpWyX
jSC5zUDShQSKHJQZ73heOPSHHzWo4zA5ikbASzo2tRhMZ5J/lePEeIvwOQVsFMYneZ0HfjZpBKxO
9mdaK3iY7MXW8j1Mu8EQ+Kr7Hsb9LJ8nwFs7wCIW6PgF1uONscZ4HTUpt6PibjDNC3Tpjfk7IaKZ
wmK5wz0dib9jonXO921awK8bbr84Ho3xygl8F5p6/OPqu/2TF6WwqmlrorV3GzjVBwuxIKqddyv/
4bu0pNyK2nt/KYeiuSEvNIM31LTOQvEv1ODVo+D7cJb6cHXIrf4oSWIQt/pxTn6/FsaA86wYpjH4
yrSdYI3tFSXzmjQs2DkV2NZPMSph5VoBlftw8uGRPl1d6ba7qkU+H2e8BqI0zv+0lDaUaOLzaNaH
hSpDNXaIVN6thprrENGrr+41OsvyfnGFRNq6vKnaguXQ4f7oJV/dkYtH7u7yr231MQNLUXEpavP/
c/SH5vsmhZVL/pIx5TSKhgZD4QWgwffknovouBVf6q1NI+JZw+1Os2oq/M8KYugR08Uocje5aGyM
+b7CbU18i0pfAHbkj5iqr/ZwYTdtuV6rcihHZudtZrVFa/a6XxpY8/xsZubkWKSpEo8/L036OfcC
TfvI77Yt5CKjOVwFcpV0Ho2wGrZ0J9aUAfCYAsQISElivDpMaigCRuut+yjqhbFmvanOi+TGpsJm
jT3YUJCxSyxwQ+seIuAip++e2W6Vi4Es5LEhefOiIZy1D3oQeC6RZ04+KiYSb60QAj9rebHKTode
Uk5go5fnH91ofves56zD4VRD8XQYf1iHoYaP/uAiEUUof8Yebb4OW0BII5WkEARQpzTrBw8wCWlc
R1SC+ADDNaaP7otozmLGJzsZpRV6LUmW3OUGf8Hb3ZDd2vnKWZg9WHxB+K7T/WLIiYKrCdIJL+ad
6uybBIxvLAwiu0QS3G3fX4eYzWlMsYOwpAVwPrQQNkGABGeieE6QTLEHNIxMFam57Kp3KphCtwOy
g8hDbhnP5Q2q9EZ+p8pFsdtTHOaRtHzeW+ZCa21U7/3Aw5NhupeASO+hS2Mb+YUjcRyN2sN7D1v0
jsGeTmDxw4aNLVz7np+gtwzubzH+yGwUPbNEC0TNT0qHjtdVBz142bb2vqBhp/eidXVOhLp2r6/c
yp3KTfNUqJBD7KUR2CJiqbgxcTLqyeB2YsgCBsjbiicxWVuH5E1GKNGJQqi2bzv1gZWOfZpCGHqE
wnpE1jMAkcxHcUVNkx0XBiOdGGUppddUrpNG4RFTZjZHvS02zoeW0PSUm7cMffujM0dmrERTrfE/
WouryZo6q3E8Wymu5+dUMxhYTflMu3IpLUiNr+NnPVa7ps82/f660HQC9OkjOJ2PNkRBS7lSgDfF
QuD0TNlueAfdclhm6nNJQ9GeTsZarPSiNkfJ3+X786auNNG1IKrBhyPTSGlyKjbIysB2VCHMGahL
yausQuPNeMvBp6iXM38HTNjTC8u6EqRK8yWw5u4puZjEKmqe5jX5eh5okVAk3xy+hrF4IGvV2asT
3EFKvRAyMSLplZxCcU8AOterj/qwRcXbhjU6E4sfkJDshB1+D3wDYuI3IJCt1Ob66BChrx/XmA1i
BZS3MtuqwWJSda7OhFX2blcZvo7eK0qbqwWsJIBxyF+pI8Y23ilHo7bNziwRG63i6u6UpfgQ8V/4
0V85JqjnhCEXwxF0gaVzVXG6J1dVIBxMcMoWfDYSG2Myv54eFqZiOYen0Ke6Lh+WckmN8cyas7T4
Ei+6oqaDvkMQlTLyEhsi0blifuBkC2rO4s+u52yIqHstSrAkWVnvfiVaBhvi7QKKEunFQOhSvoMx
Nyu2K2Y8v9ZiWFP5T6lsIsncZTS3TIxwlm52gaoCWcfVKR0tLX9DEgpauu9zqAB5c2qqtiQCFtSI
BZxJkJN7fYk0UHKZAQfDkt31Nc9Si8E5Ug64ntT03c9lJ4FmEiVN/6YWdCEjI0pxjfRL52wO72yS
mBNtMtCvqKaJUTVIjb3TXaAVEE2EI1Xh97G3l+1LgfQHyrqBtZs25MWlOoF1D7xVJ8jcaTwHlkvR
WmKZv5EvSO/grGDtOuawLDKcXbS1ARg8lHNI3HsPIbzw+TrqLuVkPuhDKQwkVdTFzbPdQM89sA+V
2ufHQjmuvH0Z9+OyQDtl8mZ+UMrCKbn7nlWvG/nRveKqPf9Jv7S2MRHzOpXwDdE1JFgpneGCbgY+
ugXEvgG9j/oLifBDTKkGE9tIBRvlzTSNkSIcyjPcOpgnq2CDWzClzqNtWGVr2/hC+o3Kup76ejsB
F9AzTK2L5+OoNoL+N/atw6u64Nc70SkpshLvqofUGKXi/TfdJCWaCuFu5VOYd/q2ZLsqmGNETw96
3pFrJ9lDmca8hQZlQ5eoEvKRrHGHxBVHgNxqLAfZZLkcYhdqpAjxUvlPVTcCwewaQO81Yllq2hri
QtKsiOkQFdeNkLibLXJMkVolhTGHCY7ke+2Jf0TSFgxlHFH+n4Mg0mGX20zeLX8zig1RI7iUDCs5
jIZiwUn+E8O32ZW+72VkRCz8QHdr8vpLc0njiHpyV0sbBKZmjDhdmLGbSC0RJf1NE7YS1oxvAPQ4
Bc5LuWz/2kTjAz59xEiu5tU2QSfMa6iBwwfHsz30h/UTbktB2ifV4fBEjgg0Q/e0FCTnscEMz0DX
iZaA9MBqtjenEraCmfhSEDLvz+rme7P9Szl8ao4wjZWE5M8rrTf0uSllLLqClMUcSSk19dSNzFhg
jlYZv6+UZ1JbZY55nB/Mn7zMmv6Utfwn3ZIitKLKF6eflnIyruUJqp/uTpvScWqMS1q5X87q3BLO
ccTtQJatuTJcBy4K+UskmoFVx3DU7vzUGhEotuHdygXUadtL9d+FbXmFg7Ctp9K/GN8V8imLGUxn
IOr9qv2/CLXb2PnEsyPqxU1xQAZ5qp7HveYNQxHv1GW/WBmt81o2jx8zcP1aypsVAd/RXXaCcLhl
L6XlTE32t50VorphA9Z/lYqAVGzMvKOHWe39QOg5bEmIM50DeVeRNy+V+8IG+Gy7cZKFF+WP0Z9f
XZczCL7U1XIAbgSMAyqpPQ/KSbDrRxy8GUvIlzBiXJ2k4gHGSuysWocXCxAjIURu0azos2o8SBGN
ccnedWDvcER5z7FJ7gHsR925oLrzKxONsld4l1uDqtntdqSqDRuhsPOk2q7FLZ0PoQLM5DvNuWuG
yYQUKzVgTDV5Us4lOwv4oalQ0DEOYTUQ5m4xpMUvICaCYYkULtYsMzJo+n8PoaHCY1t+YVWRplgT
EgenrGUnK0mQEedxG69sygPjsUDJuGv/1IA2He/KkBqvkO1Pe6weHh1dTrqc8reAMl5GFFt8dWro
Njk4YaidYfrMRwvobrDQMIG2lg0viujHAR/0eY0xtkHwAWA6NLvebUNyHIFDWL98yc6RFE0zpU2c
0xi8t/lVMmQWlKPZv0mb4PM+Ul2x7w+HlMXfZqDCGR9jDJnPVkWCBVXxAMis5wwUlp2f0lvnoLcb
91t2O0q6njkj7dE7CscgQ+euOg0Lx0GtAn3tCJdzULM+MHNmUCR3t+hhYhZ+CtB1UR4KO0M/Ik4X
d4utryWldqRXQ5hKBT3/EEeprOtxswkUw5TdDJufDORZVDgWigO4hiuPXjZ/aYDB4JFULFdyU313
8GJZ8USV3UZH+GGlvHUuFKwqqegCNia7OVwyD8aMmhnhyxIM2hYluzpxe6cjbHcHbNoRNh7c8qAl
woxL/ljV7Y36PDG9z7lT4uh2OaPO8p/DOUi/vW028ymZu/vPn3fuObxtFFaJasivEkCI2NFufdUe
uE+o+gYSqADLqXN+f7DL/s7nILo1b9ddSB2zDG1okogqg44RoFwAoRUQBN8jzcPLZgk2rqoux/LL
gY3BFb4+uTEeMm1jdUWylgPvM2Gv/2/SY7vGD6RcFe5N++rW6ytuMLysc0g92kUG55hcSH4Hm0Fr
eCdRuqI1KAYWb2KNZHvw1ErAPHreHHRxfyIdiDjjFwKdkHmjuwAQ4eFR0yafwijGFJVp/DQx6b25
y+duABv1L6QtydEu5+CwUbsv+ia+Gp1HlvavZO2JpGVAPrdjZw98mPklhs7iM8/eNCIuFLPMcsG5
DqsiApkFIiDu8SuvbYkd2Cl2++NTCv76eLOeBJW9BLLbVzoYKge5u64bKtHGibTvYovqJmbEALZL
bNc465zjZVSJ4DRiJNxrijajk+IURiZJqElZxpmPRq8kTa7rruoZ8Dc41HMsn55foBswAfFOQuZE
llmehtz9juBKkitlPsJdDHuL+32KPiDy3MaGApF3aNTpmOrovTXaqEfQ4dih2exbxY2g6oUlp0s+
b6/orW4YT1vNM8x5H8NA+0z66bfDImxZhDFajSLyqXyvIrRVhRkxynqDm5isQJ4XBQ84RnYe2TYW
IA1ImGOJKeUMqwFRdJ9QX1qDU99jQibmJSfVe/P62vqln8r4/9Anyf4KZv00/nyogh/gLerd1xX0
54PezUgzaGulF/x72+lUSFJiAXdrBAtYoKaClrapg1mX1w36qM/UBKvVOf6amx2Ug95sl6cBlxqJ
iGxCHk3ttLPOgjPB8K+ysaKICH2LTVdqukW9tqbGqSCB/nPWIBikl1yNkAOA15kPuBlMFWXzSiL3
JRDbfqX215BYkgPFV7CW8XkLcsVyoAOqfH5zfVEhDw+au3v21fL03QVxGuafR2rrKfoRSXT77mFc
5BuAY1FGdjvMDHXn5Jk8JdaRGBG8wqQByL87NOoj4EP89Xmx6vGzzuqPpztM0/UGsfRopAbkPc0u
vVErcb66EZ2rrI0D+NkCXAkG6YcfETImGQzZAMzHG+I35hn/d2AU0hujjZWl4HXCES/zmy1qy6Hr
UEYuRxj3XEk01hXQvPM1fn9UqeD7MsBMNNjDfhNBXGec2aGhtDVR3vR0QKGw4XEOHLnbnphEjlyT
0z2Byvj1BFNJQMuLCWHevviyPrVdAYOvnlqaDKutllH1mjRWqSXpeSWQOpku4gytQXuTDDas5p6h
Ameq0MMGoQsEzNfQSGrNb+3Hc1VLbG82mUdiHD1pGntw7oMquuEFQaft9sitK9k+0nZ3u9PNCm0i
dV37/cV24CzrxsXoAvk7xfZqexfwlcMGGfm8PK32Nx/mQKaWPGyfE9rOMmbD79F1X/VsKqO4btKa
IB4ENUBAaMCiAhhrMK5XCi/Nsq5XyQweAPA35hseIvsI9e/8lDJyrMTFVLnoNsnwyQ5X4AzGJSk4
+ov7b44tytp78mZ0/x6+p9H3Drj27HPIX/WaYNuRcI02J0CymSbFN8hrflaE3RXNcGxvPdOc0fN0
StMNOyhAy0s8k9qx1JoHMCQ9ijA83w/l50ltRnGjLbrR42bY55EnEzusBdMSv395XI+A8/IWS5MR
mnk3W2NgrGRW0Kwkkdgff7gsTREzHQPweowyRF+pwK6g+2dSyqMosM/0KCNCE8r7KfgLKo6pSgil
IgySJ4H3/6kIspocWeNwSObBRWi59rPo3qXPuDsm1P97xKYXdQMOQbHrOuaiFFNUZA2wx/FQj90s
N1pD/L6w4YDtJEHFeD15U7W2mUCW05U7NeSIX3liiry/bQxFTASqGSGkCaK3f/Up9/fFGJd4ZiT3
ruSW17dKNZ6ywOZAIQqntnsDRRZ5HMXyqrj38dBtOhlMV4j24cF6PiKe7YtERBNoxEldytEWgGJy
AWvHKjyPgaTA43Exy8tkeF3I+IqIMRGMrpeP3B1YaDQ+WK+/SXV7qP2UR0bz7/JlZke1Asg85Nl/
bXiQ1RruaF9vGG6RgYZOdHOoCUU/d6IGBU7XSBhT58kDznOepMA/mTkyb0h24huls2cMp2lSZgyA
2xmyovtXYDUsRDukV+5wMifYG7iFoNFGlzhESOsYrU8dPdmnWhu8/X9YNpqBZ8UESuzJ5L0g2/Xs
qodE1Os93ki6qJA4M9Wph9oA8xV8mTFRuQMrV2FmhiSvvuGNbL2u7Btlxu9nf60vNZXt4sBgE8hA
2f5I8SCWLZfzUr92Jb4kL7lInljfZD3MA+RLpaD58Fkr6ktLhdLr+dp43Qo/6PnkdpnbsHa9ZLax
r3RdrkfOBOmz4As3axvHM5iCUd2RR4U6l35KDKxC6vwhKnO5Gc4LX0VNG2gkbnh1ULLxtewFG88L
Aa1sMoSIEz1/91IAddqDGAIh8y3FvuHNuCBTgIoKX7tW0BFqTVRoxf2D8lXNbwVduE3O0BIM5GZ4
2Sz3XmeC0qYvbQLCrfLzE10ye/4RW5URgIr2rNd27/eHb/Px19ChcSljASJbUEt5BwJAxkoeUIaV
kR62OPIMySqBIZT7FgfuT3lPr9lm2S93HxaqZvrbIlKW9VLCfQ1DYR+Te8Nn7a47QLupmiVLUeC9
TT0l16TKozqr3y4tf6EerIwgPC/iR6MMqaJEuF2367ZwcDrDRngaWVz3KI4MktEpwiJznUgjVugl
Q5ivP0dpXNjmJia/JD9IZ1QjsDdckEJJmKmSfAXRnxMOPsxVPbk0BcSO7lVwlmI5/xm6tZmEPv6b
lUSoFJsdHKzCz/x3/SpgwDlyl+v5DfVvU3yv+/gLCoOEBbcKTR/OT2OOIzMh/m2RYrb+0sCoRfFe
rcCIs7+S+MjWKl/CjGj23ncJI+LRvm5KHYl4GdZ/g+DSvARONTqP1zJ7u9UZCgM9Uy68iDHbI26A
ZUb7WXP4SlIPwhHJ3as22E7t0vR3dS492EANdEfHjrnNedIBbHp8xiO+CeR53tqjnA9UIkybRBj6
+EeB0u6Tt+H+Kcoaww2CjfJKw5R/1qgl4m6/kO7V2XeUKf8SI92ml48zYkuqA752OJB/Q7N5SVy5
waMcU2wqaqsF8K0VzxGQGrOUeHYG6+wPQARoOPmhYz41HxfMx6ux2aQsygCLnV0jx2hByPDa6OTx
q0eSPMo9SkKRMeqVAn/ybO2YBdo9v76SjtVgz+BXMSlz/wP8jAqxDv/niJ6rOOazEuBMgypZN/l6
1Y/LoLFCXNwoPSN1G5kXYMU6R1NCXwqqeiWqZlVpjH3kjFmQ0lI1HQo/vQJ5GqrRZe4feiFhMzep
gej7Sd6ICHo0Di/J3YCGpwqcS1PAws4NPac2tci3HABddLLX+tX+M1FYDQ7+BoXl/nqof4a4mR8S
f84vTEYrx1JlC/rk6ZbDPDOKfn04v8vsZCKOc39sXcefNY6eJApt/2i92Ft/me5Q7tBkjdZ6XqL9
2X+vpvKteOCVAM5FphZkfHYcnbvaHbEl+Hh/DYTHNPwwa2yERL4GWbKbEVE+LDi3co6PuHDC0Be2
Mbuk13JGxK229juRAOE4kooZn5EF13Oafl0IWpv/OabBx4jx3+RMxJUl93mbzEyF1eJLy3LK/RIQ
kD7FcjY5tZ7y7QSTnC5y6X2yR3RijL1MmM5x0mLJ3VhJLp6Enl8Acup3XLAklzyA4Rh8exqp07Ye
3Pr+aJG0UCuJh+0PRyiIfJTAwCXK1amPddTE+9vIKR51qmUyF44rXez7/0AXSGTkIlFqDkfsNPbC
SuVikApDxqTFFJ7FJQpxCh646q4w8l5cotqPfHcKvl5dvGdQKuqpIHCxISjmKjJUd8eXnuO4J34t
yJeDBq75rhh8PCqKQzxrr6XZaTIku/LJSkf5hpB5LiMgScyVnHB2fB7Ril/SGAv4U5D0HwkHUWY4
/XivbdKmZ7eYCu+r1D7Tv+PWijOGc2dMV71YUEO1EEY0LlBv/vB4dSxqE6PTVSAK5iqgfGe7usJP
CzzcwfJY2xTQ4bvWniWa5mm2sI5e+UjGBPAkL/te0s0krENQTpqeGXN94jjquDoBGQD8tgsy53A4
9iBv9QXGf6PUJLycSFSyYZFSgm02wXWl6FUvTq0ebgb4i0svbjN2GQFPwYgUcjS66XVZ7952U1mo
ThMFWaeN05ACZOCZKn/12kLTJJlO8vU7aBE7i/ccHkWKKL+2bbHyyUkpnK1lubchOfFT1zUgzKhS
c4V2HGY/JIicnJokcV/RhaOU8G76Z36fx4Lb3pMqXlK5n2ZiWq8bo/90C9gt39w0BqagOApHkY0S
LHlJRYVbDKGm53j19kQA8jbtOC/kviU93tRwWAsPaRtrQ6oE49y1of5wTgaMxmrRCZeMmetDXs4b
vCV5F2FLLDM+Xcc7JEXNzJN0Svb5YOdYf8hFSqA0JZoo4DLXhXIX4oBw0gRLHLeOSiik9lBEc54F
PzCShIPCs6lcWo74LajTO+Ax5Xe/1T4IWzwFgpxwiZF5bmX4fVptJ2Zvwsqm1mGN9Scgr9mzymVM
kYn6Nmu9QTCsrzpKw/KfMM0o44pPIeYUzdCzVgik5HH10wIKlI8MVn2z1oar4B8Hq7msF7vkATvU
ccjLMRZB14/Vf4PXFle4YFMibISAGhE+Eq/IcPupybDNBc3qK6XZ7mP2xXBMNxp4BthvhQQTBB2S
INb0QmprLJP5pF2zam/ELE24dXIODFo15GD9jWIMoHzELsQFOkLmtY46rNi31VErbYMW5PqFw+IH
5zp2tt7EJUaAAU9xbsaIgmUYqiQ81VcTjKaIQHtSyQ3sow8q/GjSVkWz/FHU2h07+bl4hUD6nK6F
3GN7zibJDnAuPd0AByFv7Zc1IHWMFHeQJ6fJScFK/VH7Ur3Eymn/lkAtUbNh9Xw/kVhugmeF7xw6
+NcdMkth4QEAmoVmJesARqZVLU+ypx+BZpJvV0A8uz9f9XVD41t80t3XxA1yqVetbJyDbNrO9MBA
+CTr0YB5EMTva6d1DD6KfuYmTnEemmoTWlcJ/lJOzrYnEUSPrw9qr+UUnVaZUxrtIrI1opmaHwXd
6aC3LzhdIkzkrE0R/mqBNChgjGfvDpfqrP7xjtn/lV/o/5A/nWuj14OtNmHaekAxhRfSQ+6BiiZG
cYov8bZ7LI0Zqr/1CDAtGwcE+lFHF21hdm7RuAq1072+mwCQTyIe5MSbUd2eG0mQh7SOWP2d+YJt
7CpdvqdGnfuWCteTPWK4B2/6B2APSG/i66a/a3+++kPC0MqLabws4hdineoy5pJE+wK4HaNOBlxF
UISNCv7VLPIHsYd/iQHq0e2F9sro1lxNmVMLfYAbQ1eElKAeTq1KUA3oLCNd8rWUolv/8Xk0p7la
YZp3yaVKecxQh35J6iMttW4mmseCYVdendvjdLct/Hxpypd2XrPuVCoyxMIS0NpILq3of3ZjJ3N+
6Cy+1AJOqptBjuhDCiJ8YDzu6MSmFgYiljnOlOad8hx7tz5SJoQI5HSbvTGDc6G+agO8WlZ7ccTL
js6Zdm+dydKF/CO+NCvXXdqZwqSxjnrPiaNkBH6BIeeD4gK+PAPuAQgd8O41EgmssTPZDhk1LWI7
SA0yDk5Z0uTulkKghCY2qaz0s5Owl4hEiDDgORqAmvCAJi4e45Vp6Oy8/fBysTnpORAqqMrW5jJ3
j3HDrRfPrlufevfJFY/Bug3fmI2FSrGzJIOMR31YeOsPVk1SlQhVU3vAYadajHF9J4HyUfSAwqIb
1dHLJi0BkljyR/4twk3myJpYpHcvNv/eYzD8LKPBEFgKjRzJ9uvks+GZ8YoZpmcYugG0POY2iuCd
mCIJK9zTI+ggxpvICBBkt/D/YD/boJoaLCKlUmdG17Ru53SARBoJc9uaeUBJLPmdnC5RthhH6t6j
6brvBKru8F7amDQc9VPl4qxsheXvUa73BNiBrbrG1H0RWQY0jIQKrlYBedus5y6CFN1t/GDRZ2uC
4m8boBA8Cp/jI0Ou/bJPvq+55mSz7Aap6HmPnGZeaWtJwrXQWrpkjvn1JYK/ZCOa4QN0tOunloMG
CJlCE7pdrl+e7/05n5jDWUohOkA+NCTZACL+WB95OcWYfUhoJTnpzJ8Cn4ZQLOsKeRdthmdNvOvL
bpXEbujSUbOoF68xAOeVnDHMJh4AoPFFwiPqMc1jD+yR18rdfcYv4rpRhej91gfzFKcHED78ecRr
yCt8hUAh7lz2pqfIvyNOLJvk/f7ZKuj03KaebP1fpyXvxBpxngu4PaJvHdQ6uajdNhWQWuNA42On
hvDuAKWobtsN86Lf6CqM1WngFwoJvJDRHznx5Qo1PkW2kbXh8wUTgbRmYwG+b4hnnKAqqHNsVASf
ySUtPEt3sSy2rltoDz8cBLXVPYqfmOtvIwsj7vXHg0Lwn81H3mTwCoAKkQ13jBdxwYBF3DLzCj0V
1MumVPlpqv2p2YDgNt9klqrgGbQEib6i5qQZJdN4PU1rEkNM6PzyFOqJ3pps6y8MxHykyOc2Lf7E
8m6PNGPEJ8BeevR41JuWqG7WajQjdBJLskQ1fSvOE/UIjrynVRnLF0osHSmUGr/rcFca2w+oZ5NE
l8St0Gzl4vutqqD83R9Y2Fv0E5iBPJJhUgozGOCdAhSw5Gm/8norCf7iFK/HHZVuyjBa9tJlY0FQ
a+NDuF1BEZXddVFpNqHkmnmuhxOHr8ZrEe1naVhXRFtDEtQ51SwqRVHJ9kCPxWb8B9I72+GQjk0R
oldDmNXpIwz2Q/k9pgXUw6OFmPEi8lYAje/6PPpl/qllLI9tbJpfwLtwVqKd3I8P2gj2FGzkuaXc
XYUQQgltKl8wX+MhlttPLEI414OinXhJO8lCegqx2HRNMnEHeCC+Ou6fTSvcHu6+S//9wvUVskOp
UqGprPWjgSJVN8WYJx5g1c5diBWc+Jhb5NDfRwYnWxUZX2xWD4c4Ll7bKGlLhfnS8QsFleqSZQEh
CDzeS/fr+BMTFwJiFQzOGAA3++AUPH+Xg7wyOPp97PpZ77ByXacANiVd9leSfQtoMbVl5dYhAwbE
ekM/GoPN4H/91xUHY0Hb9tWtqn9Q10jSrHqdcrpnGoYfKtkDIPL0iPYbn1nKJjteTD7tNyMsCKzb
fyZuUTqA/cd1A+P1FkTwdPbpptS1Ac+UVtV+B2p1C4KT7+y7TsmGEFO/tAHgy0JT7lE6lztV5On5
3sOa0Cvr4VVnCcZSFM5WVtqATtQC7YANpgtP/kA/cJhxqCm5je51SaBQd0/SsuSnGa1TnM1I7OZH
EwINv1odGYSjGhJmy1ZG3oqkb09cHx5NiXlptYhD2DjM8hQNFL/KoFNsrDihbcZzVV5GSSMP4CVR
UMU9gO6OewEMrOTXP2FvaD8iGN2ops1OyqRl4JdzEONohHm9s7DFFNyk5hgmf55GyTAMQqLJQzXJ
hzYKvm3QBfan6w2D123CTyCn9OPEhFPOEzvnBhPvPmAkX3AFPD3P4SR3LOgdGredL7/IaVfHnUFo
Eq6DxcQCbvlg67GHeQXwyJVFM0yrO7R2psWWd13niIO18XdY0OUiwxOuNopN5KmMKWAoaYyLluZ0
DD5uGJyNaNuD4npUH/QU+dfFcipoSklZRPlUg3uaQQOhDFJK2IyQllApCyo1YRKsJ+XNJjNNJkzS
AX7OjhE5dbhD9SF13giCekN4xv+8ZiC+NLUqr3V9EzifylN96KLidsZEYh7hhd3jv9fTt+/CXQSi
pnUxywIcMiyx5F8BAuuhELf3ceOLf99Yz1+Pos1CVYOIwwzCtAk4RFHjuOdBUjaXE57ftg2uv7mN
p60zeZ0Y4V+b/tDX0SBVquXoburZoz2Ld7Sk586a8qEqGbyH/+zLuz7GMCQ1lcGnyCaWEX9mjd4P
W+T0r/nXc3L2K+/J+y9324FGSN1G3vWkYScZkokXss/dqYMsqc8g4viBwshgFimDHVPkPRt6cifl
CFHW6+1PyYN3jiZSoqzJ3MZZfSSz18CwGS3aVoblc2obp0XhI/eY0LKXW+1875Dvlr9SVKkBO0M2
ajMBdy+KLSdSnE7HzDlHhk4BbjHJoSGY+I1UOshP5Y6etZaVs9KaGViJ2oP44WS7dxDO47/pJMFJ
9XPOI5KfJ3BTc6NtRJwagCIOUh5APAcv1opaP+Ahyrlfc3ENzdh0KqEhUvuJuSyiN3Y7wSS0VgjA
QFgkxzgX1xicwjisZRPsdEEyf0dqG4D6y4YqCWcySSiSpZBX4ZU1QgK1D+icaSZMN3csSxSV81Zn
zKc0M/cpQc+ERR4qJbglRWRMo5Cu8f9QNO6DvMaZSyambhJUP4FvVXhD2oI+e7SDXQECG9fV0TXW
6XN2ZXw0rx+OHsgQC5tKhKrfJRqFx9QsGRgsWfmtxZU9q5+6COKHCLs8A03jbi2qsMRFinxCg8Bl
cvqj088C8D0FAmSma4z34xFUQ4kL9VI/bHp4SpxPj56yrt3GD2BW4/GjewJDrM/AcFWK+H+3uqDX
zHzMLieKsYo/0FS7F7DmOuEz9c/U9viuBQmakv5I8ttzepSAavJxHk4xeHghTxZbvpqq1JFQ3+6Q
6Xn7bHtExnKcbgvA65FhLremO+R2jUf+4gUqxb81YdeY2Nzb68rfita83kV7gh+chxOuTqvpmBt7
ZfJbFWNDn80VUwRsGh9tHeVqYNAllWNTtBGIM7Meopu7JuB+4PeFddePzpPzJKNfNFj8T95x/Fbh
XJxNMjqrjNR2uB64t6y5+RMSvJ2njJ5my8eeuEwTlhFTEXbWzNfAeCnhmb/OUKWk52JBds7TJp72
aL4SuEjFoZPdU/W+YdEyEcCAZntKwHfxUossVq7lvVP7dQJBSoZCwxvyCh+7FrP/9o1hMYpX8JcU
c17iF0G+ekXIqigJ2ZxlapmkWxZLcPcC85vZiR0JDLe/WwCt9aSJoqky1q1/DQw94MXduTgM9Ktz
BuciV6BgaSl9nF7VWDZwfHtwkqOTFl5Cc9dL4VT0YUHfMm/og2Xgz4OTTIW54v3X7YkYFQKz9WfF
aiT/zQvg2gyfL71KHAegrs+Gir24h6aViXj9QyM+Lm8mACAXQ9BUzpbbGhrut7IwUoXe4K2tFm5N
tm+++7xp9CfJJ+sA+G6shgY+kdmd9sRzn/pZGvlCcJ60nNRjN5lmljzQVh4RokZ5Lb4sGuV2IyWi
Nbpdk6OsHhursVIgNz74WEcLMw33F8pH5pw69b9c3izz5wmJ1GrCntd2WGyivyaSKQxJ5QyN8/i/
xeaBEyZmBmx2WC6d92Ckqpasa/tXqKQnccxigqDntw2kBEUawqG04jsNXY8uaexLWApRmXhLmjHl
9nfrvaGd9tJYtcCI7OM3PByKtGftt8I77ZA+OSy7Lv0BXltpbJpbXmCsbzuLOwrZzM8mis7nJCaX
+wFADFXAA6mrpgDWgn+N5IwbeWvog5Q5B0BiboQrbSjg8hE8oUk9sFDHox4EbukIGMY0oc2iSyKo
Xd4JkQwYKVrTtKhYpLXwVZww/YkRDN00FLV8BVt918B9RLK7q2YGt2wSWtuVKhS/2blS29LA2s+E
uQ82syZau/8adJhYmIIBEXYxTYHSMF9Tgfk4gc9D11ETf5ElYu/pY+mGyfN6nR81yLCXX1dKL0da
Y6BzNH8DOFrQNVNDXIevB1/6/IpnN1xWhYuwpVwPYw8P0b7F2NnPlS1Ir9BX74Qu+RbPUmUChcWg
rv2zUw50xXRnpM5pzlYVRisz7lFuV4VdhSMMZlPpwqc+ebcLMlAvOWwTgM5jEuXNTyletdM+3P+t
5uIo69i8mw7nU6p9Le+RfDYeQSmVSZmWDWHYiSmXjSsdqiwrSBde76277stpNPjR1o0Yd08Ep1Ny
WYwgT40wuAkZ1pvw5wBHf6Bne1ejJdWLDSUAO5OefJGXVnAgnakTkoSOAq3/6bvQfeleDI2zvNzY
vwlsfpzBdguIqBLU3i+BbmpqXwE6ckecP7c2MRhI+IaLEUXP2DQ7p3Zd3ZOrXPF9jANfngPLT+25
sXAboj0fTK1ObYGZgUOqLDVY7mbf8BQZcQ0RCTsA9ntd/zdrqWi7pLTgJp40mkM7vcmeXQSOArIr
I7YAJ8MT1V1UU0yjgN+iXGLBLW1U4OLMAvSmoSUZva7Kz36lb1WWuMqP7lE0KZ9V9GitmH5gwz7D
oD4v7TnQe8yUelaodSrKd1qyzUDzcFnxGvoUtTQQHeslYIg5BVOWLWejSSVVQhgqa0p3MgFVtEr/
Yiq+FnSLSng4ed5212wO7Y9ZsL6HK0ncs9WXTLxhV5JFvjNZPiLjvzzhuJfEHUM41CRPxF5fJaOF
9o8arC67ZAuhoFWDX4WvMTSW3UJg1ehTUpj6Ner/p2xABvzTTZQIHGDWDN0mjrH7vzgPpqTpQxf+
vSRxn06kSlPym7xsbQEDOGOCpeQFHcuHNUJCo+oqLeZDhglM6y946ost8YOKr5Ri6QM2TsDTmqYh
OwbhyaK/zcg///UQhZCFxr58VmTH2JWvzPN7dFbQcFwBCHJItfpQ0gA9bLPZJ1UY7duvQ6HCOePV
1a+4GSHEtLO18eLkORCKU1Cljx4/YMjv64YbcBPFdOynb0t8CXzAHwBNAQLxf3WU2cOPs/9Mar/d
QNf/H1OrqYhEK2Dgf18L0vDaa+7G04uXlX4Ji8nrwDyR4xh25MSUTSjnxmKxmulDTlxD6mOeJZgu
qilyuKGtdghOBplkiDuS6JkM6c3sDT5yBb2yF5oheqc2AVNmTBbroxT6l+d8sEDp8XygOuZxbE0L
3R8fJ7kVS1w8cY0fs3QuSjI7VnApPoKBh7mqUskOjSou5dgqKaHNxFDTiR63Mu7eL3BBGQj+p2sG
9zm3PKF9DxHZ3g0+CI/iK4nQ1blnaSK6bUU5OQ3IgiTDc/w4ymtmm1tiyOkAMfhLlDtKvp4zHtTg
MyotV1Dj+kciS9Q17qLU5CK6ffPIU5KxUjod7ZmeS6uiLtdKDGCk0bptSrC3cC+bOdqTOKsiRf3N
XKm+IWKoNNmZtWYkgCijfLORdJDTyBF2ZS+YZkawWuBQSHp6qcln3+L5oqFhhvWyukr+w5iaZSLU
Q2QclWM9L51kDX3llc2icIFiGl4vn/0xc4l7CPyKN8ubiVNg/5CyP+tl/5YCOdCdP3r1p1oVT9bV
H/DZCMQxvqJSqhppl+dd8EnXaH+us+wPNWuWF1gtVcjMWhUPEIgSQX14f8FzvGShCGNFV/ND2PrQ
YcR9QtvlKmz2uRnduYPQ2Cx/jcG3vfOwyRkK2rKS4Jzvj6AJ9SDczYwhV6Kko8LNvwIstEM9Wb3G
ukHPwpeqGZaIazai7+2JEclPKi3JMQCfPrwtTk/qI3XZUQEKEUSEN6VEpB3Krpflc/lhO5xDSa8j
NMfEK024GvbYC2jPRp9588RepH+GT6F8LhBIeAleaAIkvsYa0jaYmeItVMf7Yq7YHdY6UBbP63wF
IpxaXJa9B+cMqnVt0PUeo2UuPjKiActfmtKLgSqM8Djw0J2sfvQ1EMas7o0ZtYLaIg6CYXzTs+Bp
vNFSRJPwEcVPz3uLrc3Xf+MHfrz8NTIOucqTcE6nbL/8eak9LxWJgWKMztzqrWLzRBkiI6+kVlpL
RvMaL0ICYPWBrFqFWil+YfcPlDiEyHcikQ0uEfCPlJJrwSxjBvoWwhu9LZfkxDIjJjk7odETFAka
o2xXZiLzyqneZShf4oE7imi4YVFSwlcZShAA3AFNCDUHOfJPJc1lmm5wqXNOoLQqGyGzrz0SGT0D
4nEZ+X0/by3baL0hPLk+yuB3LfV+2yK73nIie+OTy6nrTn57XdMDn7+RZefubt5xNgpHJuIjKnH5
IqlyOJEB5ye2e6oTtWKPr6yDIoZMbw/UEt6JirXSwMspQbriBAeYmKqy6cle3CBPvucwc1zHH8e4
c50Pzip2pqLrK5dFJz5YgLVBAq8C/4XpUkHeg1BcXvQeSoJP0fN+NQtqoJnlQQMuOmu/olwHqsck
BZPF8n/polLS5DxE/09dM6NLulHEbOXp2ZpUBTbPN+qcAvv8cngXWC3Wo/PNYBDiAFfxWrE3oPVG
OpKpvvyotK4VXAcKvskLs57hy1WubLFmrVDe8IXryjam7lnhkzv1Tu3sVevgVq+0Za8rVq1dWTNZ
ThxIC84D58pURyS0EkGaV+Orq38QgZsiqJqOBnrCeeIf/XD/vvi92/+MF2J47wR0TDSUO9+/xk/L
9ruWSB9Wpl2B2Jmsn1/0cKwoGjJ3uZ7xK91+xOtEDOiVZupCAJqUC0ZM7SEF40AuuD9xsNKPP1v1
fIjW3q1z5HRkSM3O+SvEaXAYzhB/MqBbQ1tGrSJyO9UUzZVbghGe12Uqx8wrPJQ5uKk2uRNa6Kss
gJ/GN3sE6jkueJ+CF+ju3lolkNOqlVTDIhQXuPNW/mMp54Eu3FGe/Ppfr40t+oHtFbjwo0kCrvRF
6dqYyuQR+cSCmJuXjh1ImxoNX7RHHiZGMv6SSCMw6FoG+/zjj+lG9bQzUlPOQkXPSEsrgw+OEIaJ
39OA39mXrfxHk7RVZP0LTH7mC2G84bRgxZA7fyL/3X4m6t+WTDjzabnGTzC+EMOTmct3jkKjAVBU
3ngpv71GsCpf02d4/EKJIVqMyUuTL2dj5N7abV5ztXmEi03NCIvo2DLXrpIVMvRdyn8fgau45BwZ
XZsgIPav5CUHB4l492X7fq/2LjdgSIyh39n0AmDz2ApXWCmifn/WilmsNDExMi7Pq62FoW7wyrUX
JoWRboB6+7bZI1I8bxtSPjApz+7nRoWHeMQJ0f9h8XQmyo4FYGCsdPzznFr4dq0ZR/pGXkIPjHOg
Z1qLT7i8BRwmr7gCS24RTVRn8vdFpWYI7GudHXSyoTHMuzlTps/qeo+sdpfirgPs3YaZd2iv/C9+
6suKGSYfraos1qtbzaPiLxk25S6WSeg9uA3mzOLdHzT7uT8gmqdqwD83We6C41+rWo773oMJe+cp
reUEywGRhlO8tOBlhs5WPLMYzGscOrAohJP0P7+tA6VWcZaYWVLZxZFdal6rnqvmxXucDAE/XRyw
UEfqkrVwNlCCDx7teWx9HNT7aYceqOY4UnWXD0+Ilw4pLUl5XmhCdwcY6/THKn+4c51yavJJEJBs
eTk0aljaFWET4NMYEcrIIdQqgn89/qTiUpX8mBtmSxfRYyxpbOJeBOZMRTMUe1oj0HMCg5FD0r25
QTIKZs75gnLiDR81a0GMSXHCPwWjQGKzCSzmSqixja3OgEpfwA8VryMNxtYM1TsqXbwHUwGxq3Vq
bf++92HiVROUqPc7SdYVbMmGGcDVR5OXGAp90NvUqB53nI5iT+LkWFCnf0Hp2Vr3Q2W6lgX1QrOI
E6zApdCiWfHuRHNMasBQwWtOPKSU3LZlUGygsz9qDBLo/8iwxgzFJA05J0MYObD8CQ83Bupq2EJf
H62aeCb7cXDAZstR0FsbnAtiy+X5BIHV89f8iQQkTQNorsSK+lai2zi75M9TC6fyWb7t/SgnaHXh
YGP9yv8O00HirWccu8kRvTOyIEz5xn7fek0xANYSpRP6obsV1ZMrdai80wcupg3aiM45dIFDJicn
yDBZloyheo3Abyv0HhX5x5BoDfT6S+lFhTv3PzbsYubnofBtj0FKGFvZkXX4F+PA1o/haZcrB+gI
ZxoJITeCTdSm5BCS+Se/JJGGhcjHCW2MAAf5OCEW+z4ypL1Eyo1kfK3zu7/3d6s4g9FiVs/axxwR
8czZSbW3TAV3xPcheidEfT6j9Y18+V9AxgfneHp1L5MNreHQ1EyVC5HmZWMi8d4KS/d4YTvcz1Zz
siNu0x6Bm87PUFZHiUAzXtsm/KjAPMPNHnYPJD/aFMD7OLxJJrig1ob3+FEW4QcVDYuNRhb6YOhl
Av3RFfL64pNGxiz9TLCBUXfHwLDGOyY9wQjTYUA4X8VCk6K4pOE7I6/2moXNbJXIdYGlXPGDTrOC
NT+wviYtI5S+VHgrORkfuKqLC4wz0s9c8ZFmbJKhEbiteUZQFL60XIjZmkj3X3xBO+saygx4j5Rh
m8WTkNv/AL2dD9nKq0RreE2Gx6EKXU9dZ5ZkGV3cbGZ0w8v96t/aqfwY+954bjfh9utsYpj0CFzc
p/u0AxgvTYsfieovQZ6kxDLks8dW3OiIQQeieLkpYLKBT/TWzpxBl3qxVcZ+lIkaCiobb2wV7HjJ
SZ11Z9wnYYdRB36TlGyQjWJPenC16pqqq71rGf21+u+ER7aRR/xiYX5NR8z391STZO9MDsgABRLT
mTnxPVfjizoXKnfnFGuGdR+RyghBsk5ijo1hP3r7kAHGShZTFrij0rOXUPzAXU3mLqAup8VwwjZf
+Bj+JZM9kj97+MuXzZAnEAUdoO3IiJWiKppVFKjF5PYA8o4m0EZq6aRYwiqKZ2jSRZzSj46VoyW6
vxY6jcL3TtkZJrIQpFAaGtSpZI8ADcuSwOUJs9Dp+g94UoEXkMocSTABLaBdWurBRYKBAbHl98GQ
NRBcv0HmVhi3V8froR220pLtzVo1Oc1J94rCCYVniFrvSrpUYoofkskGp7gOOBjIJJnVImJ2mFcD
jIoeFdquhpsqs9rse2HFL6bzKwGKxiaOVkEXMPBVbK44XqKSnPb7EC842gT+/DkfE+z58/rIN3Qr
I0VuqFwjYBDkWnPu1dLB4TmaLPV3v8uy6ywXDxGbDmh2/EShsogyb/k4gg5OtMxUTN6ao/qE2CYd
6fqvgudXHwTkYlugY48cQM119yad/pA/ZFARXza2R8S5H+m9zox96HvLTlyA5ru4jiR/9q8I6h5A
CFXM5aOAljZ5IRNOIN2FhuGMk4fvsWIC1/gUTNtk7JOfm0bC5jWqyhXPUW1IgPrh39Vu63l9+Kp5
HHxAZ2wAXm5wvVsdeRhvmQHLYUUiziIjrPu/kjCgj3z0Y/TJhKs27FUJwDZi/f8+7o9cEWyBs4qa
OJ1q1E56XX+leYJaESvdCwsNRdBKp0CgLEGHp2ivaR0yEQTqjgkEpTuB6yiZ7/bGPXX91Uin/502
6Mo53eUmIUBN4bhpFVgFWlEY4yLwOI8z4CEiGRKAK9Aeu1LbyYfX7Sr/IKLR2GKvySpSvHNB7i9K
5ki6E9/7aqdr2wZUESDJtztarS8WNF9PEkDVBwipNppPC0FvAAiNki+mFXfd1JBxmdZC2uMI2AAl
AW1Yi76IZTlRkSUlSI60fwuuoX7weR93puKn4sfs+oouWakvCQerS0D2xvEW2PV70GVv2JIziHqE
j2CA685FRW6grZFJn5hppAWI7fHq7JO0FJ7hcKdba8u3Mx8Y6o8UBTiUkSzeplLAIqF7By8vX9sf
aHJ4s+Vfqz3jMhyZNFV8Es//FMIuQQ5D568SzgxIZWqgpye6az3toxLq36Rc964s+nW7PnPHEdCB
IJSZ40FlEP5fsLRvZylwd/JMCgUouXljPwfA6Lzg9qUXx4oSRzCPLVDosxpusdYw9m3mrl1IOJhs
tdrJskJ0DSEbAt2zz2Ucp2op5wkpe7u1KlJEkqki5JTZ4jeSHs//yjhTr5VTzh6suLdEEHuJuuR5
Nov93M/4Pvp5yyvYPA4ezPy0wT4oJsbPfzHQYZM3NdAIAEafRRvmwMANQALW1wQpm24xWbC+Nbso
24g+Cl1ScVnwm1MbME2/3kdHjO2vCbKzuWvEze0da3g3Wd1g8SSB2BxYuYskI4uG/pbOnJvDUbZU
oTDh9UkuagnP8kgSNJs0BfHRfDVQl2m4qKzYvGCce9dwU9YbwEdBIxnmZhowbH4OPZEOukzlbUBy
+IqLyLWqV59C/6pIlZP+4/kB9BweHl2SFagGWCcEU4QVba7Sk7ZEpHQdEAh/h3Kf0icLopJDke90
zjyea7F1+9p84uXTbFN5xDdHu4PLfKJ5dpyWT6TVWuV2vKkXRgwDpkX+uxz7fPl3hnttELkKhi/9
X0tnrVcYFbVleryBg74HcUEGgot0vXklRdzlz/oCFMSIFXRpNm5BWheSRNxrzHAPF8HMWQd796ot
v5holR2wEfw3iK/RUdC2Bf0DMk2sqBWZo+8Zyt03CkV37RIAVZquzYYGz2uHPcaA4nF6A+h9gqtL
PlzvmUBKThNdYeTeLkXXoRB8b5UdNJPXJdc+dNgt3EOicCnXuXPIEVAKQYTtxru4fHP0QIwZzujC
toiPdHxA/jNS09F56/Ve0U+BDyDRfar2IcTq55GaB3BRtWqJEIyZFIXJJnRwFzk3PXCYnDnkK1lV
ER+IFYfS+yPl2FQflq57MaOgzPQ7NUobVKh60P+RFekoFRihpL27EOrnEhhdUlcEswXibgZvlmS0
rYZYVzPeWhJAnIhOS2E16x9q/uGVbGlyAxNFXGtxk9Js8/GMNCuTi5rhrc/wmCHooqKxsLeQBNNZ
IHJukLVYfQNN/j0zQM8d1CCRyUddbLWWjSgjH6KICbLzCE+KEhtEDybm7DPrU8OGNgAotLY0Zbqu
N8J4aNVpIV1zJJ3N0Lvu7nLSO5DN6IVmaX38EXTmB39zr1tEuti9XVy3uyRhAWoLmALMK4hr/cXj
iOAi9DpI4K60KB0iKkFt0wI36kRhd7RENL5rw3o91Owkr3fYq3xvvL7yX+ykMcNTarB/csQ+xotp
a/dnr2u7wQy2iJUlDJJUXbTZdNvRQvX1ZN6dprW3Fjl9n2pyMGGFovNpQ51REijQ0tbc5wtN2Hxa
N1MJUIw86sbk7tcRDJTCW66JrUdwL3cdpCXtjMih2hFRMWDOYXXUxTYx9OBk/ZW+ueZv2PjzFp50
at1/+Ca00bScg2RX/G/DhrImJMk6azEEW2mfBS+RZrMEkm5ltjK0gsggOr0gDGNJG8A1NRR90BzK
v5WamfD6WmfnexNl3czJIpW9ApLeuBfoTetAYG52zlmu73+/cLrUlpZfnChVeCO6egZ4RvlPFexK
t+ixw4PmGOpVdQhP+/8NNiRlc2TRBkSLLkXmIpKgmIggAb0QvnwaHsx47b/L2bqY8az0IpHRJ3q7
fw1hPUP6M6OBWRERAT/EwxfRJ0SIfGd8j2tGdpYVWc71Wn7pGg2tTj/1DRS8TSYB2sGzKwiX+bqS
BxSb2kyn1Onlhh7iCr2YeBlz215REVws4cWfYqExEXI5LWDQdWfzqdfDFTZK30hakaXB+Z9wYg9a
1/DyC0htXzKuuwLqG1YjmAxA/9WdWKJ3ROis6byDVQT/tmMwTqRiUGqVgxWUEC1aPbWaQnExEgGp
vmPWoSNoe+mR2m64udfgJvUCRlg+6u+OrHX7eieCOM891l7REcA3GCWvEppQXY/KWYp27kEbFQ0Q
1aoemR88+lKFGIfYYJfEXuz53Uxii/HtfDKIyOrKuY7dsxaaoImLENPt+brMnVI+3ZnqmnDTtK/y
gvllcfFls/4Nf6/R5NHTZZKekkfrBYFWa9U+CMioypD3I0fSqbuxooiUinRLk9bi/wS9Gz+oeYwm
ElRqwU5JE9FsYiJVLzdzzupjY3udqNl1Q33EaCqsFK3CZcDx/CUKmaVYwf6nOgrYrMdaJ8ECIiBA
k0xbcmyx5s+90fwHkdGypre2YW8Ick5D68lEfOHMr4XffXi30s1ASIdsoG8He1T76NMedR47wfSI
J7rRoYgkzY+2zC+0bdOss33OEnjzi/MO+m0DK9ML8vtUr+3/R6jJl5EE5WhGBXXcp+N6BJsobivM
jW6XyFXzdUk8BFHz6t0D42YGlmVO/8fuQmSNO8ndcmBXSAJs5ioS1r4+ukSK6Nc8lgszWQgTlz9f
7p1oC7ZHXTD4ifcyBc+yAFmhjSR7v4ZbL8sXi+HqntStrHsW3ImuW78lqBnXOMQ9L+vxZTeKeqDw
f8ERWOzZ4UkV4C6KrD7IHXw7nOFjA7uSCKJD4OyFzg7V+FP0HtxEUTt8RAUIsZ4kFZFqrdrFW4mu
eHxjGLOZgBZqe6SALboVFlu1MKmhAELJxeO3B4vEsRRwOcXDeJ/xWFPfUty5OeZQaNbU2KxGDJLC
Dqhf84iAkAHVHmKdaJ3Z63i/1SzI8JoKmvM4Sm9MZ7librywiMxqOFCkDGSBsWe/ixHnQYUXT5jI
gJmA4cDMv0YQJ23pq5OQruuBZ8FPx4ODet8EejiGgAe5n71qX0MuCkdzAsxz8FMGp/uvnTgziQo6
ATkyoZQ6C/DpPjhj0zwDZy5SKks1M0jBfk8IO+9ntRPW6wkaUZqPxRWWdoYwxxgnltYJS7Zqm2SE
8Wt4cWe5in0Pg1KEyXXxNiep4sUyTzl5n0vcJMcQuzTJwrY5IL5x12hH394UP1V3fIRdTnC+Kgo0
1iLwFSQPzlCQfVtoo771TvcpUPUh4UpDm+Ch4xAOhA7JG19rhW7HlLeXNLJclfa81N1/wXn4yyW9
Hh8+WjuDyF1r5ye6MOh7bVkD3xHD+f7jHgkjpn3uiHRPYZs/CgH3NpgkvLaVnkqY0GdRwev0n742
b0H5+Z03/ISYUF5UaY9N6Sd6qiy7awcz5EPac7h9mwIn/itC9Ha5Bk3eozqvYwTcJQqGNdlxN2T+
0Ce8bPhjefDBUvUh3YtSUpMVGfTq++dXepGLVNRsManuajBbacR/OZneNLCtnIwwKssiiaC2TkqO
Yww6pILTD+l1VwOWMH1kv6eeoQe1LX0Kn2hrw3gpk2EqtFokPnZhnwDX9D2LvYOc09pKuSOblrB5
QeEaqxXOEss44agZd8H9pO3wg9QFJVcA8MGNx+tfW+gMLpqc0IJ037xLGe3t83fLoDnJgystpAQR
Izrq/Ag0uRZheJgRpvCVoxEVD4z//0MXM1EqHeIwGAin8XaLhzlTF0nlhl4HtkVyyQNS+2zmNy/R
GQVHuEDIhQqpwhqw49lQAeyX6u6UegQNAYzw5f6O8vhFmhw7Gc2fllip0rOJEthkULRf6Qg1tITM
IEtI8+tP2O65jdKGAZzo1LIQRUL5nqzSpVQnR2xXUnFayUXhdCK8IQ+2xpNdIT1FpN3cEEiF6XeO
HB1xhESeUVIN1AIjox9Rnq9kAMlMxOw2F2q9tOzGMr1DudXShhFQNfEfYrUlVpdvrzl0IMLDGMb6
BfVxNzxcGjPUGEJQTFm2OjjhESANgTERDPcsI8IamnmoXWvtWH+ByPOlMOiu3hcoIYs64ODd9yh+
G+hZAWFJC1Lk+zFE4cf9yqv6qihAD67CENZnGoa5fzs+FBhSSy5ZN8sHQYyM4K1VzAHpOW9vu6Lh
zVPrPkshK3+uBid4tp8CBbRWa9CENjKJ1PRerSSagkk9lWMkVncH0bHHZ6bk28xtiurQ7ELJx+Xv
e4W3I6hPwEg2aAtpIZKsOwyUFfZorHid/cni6sUIxVjiJ9WYhJxVL9M+NVDHfd/LDekFqAqzcFcV
uV084Q7KpfTG03KWWYw4plKTdkEiPMhUQVFWzIx2SrI3nqpylf3l/eh1vBVDn6brujy7NqMiSk4x
vhTS1IZ4lng14SaLVHnyN+vjZzhE/86JxmS0ckcNJLW7+8o+UAnnJxBjy5y53cY4MZnUKT9DqEXL
G3u/UZTCWUSXXWIlqwHvLoJd3uJjH+TC71tFBQeEWAiKVr7q3EqZ3mgO4KAU4R7dOMk4Ybu/S511
N0qEPXPo7/iiWNSfaKupjMBHAg63cRp1HCrE+YuCjWNKPU9QK/X/eRdchQHe+GaHVJTbGGHc4s6b
0F6LaY5ecQWqWw91a5wc21zcME+ruOrP9DmSiA8XxzOWdZ2fFT9US9Nyxsy8Wjt/kxpXL+Vq4Bjb
D8hYpFlZmYWzHNetyNh5QlQORJMI9aP/uTgH83M5CyEphN0jsga+zvjFLByTnnCtfexEbEyVmvk+
BxjfeA59GUzWBb+U4G7bZBZ2EFdPL85sT9mu0rjLmHx0LzgKy80ACOK8tgiPuCOvYxbI/jX9bmtZ
DO/L3QJhKE+bBhlkMB6JvEuvPmiJGQy+AXSLyDLFK5gv4U44SVg5Mw5l+IOr26zvEIyvb5kpSK4+
ae2bPNBnX/tfefxAoXfYk6XkREaszPhDX3503MTnFl/1rvaiEByLoLVkEapO7577fUReJ0m+pYs5
FJR3o65VXM4h8/JPW/Ld1z3Eo0smh2s6f+eB/uu0zk4dflAYhmIotZuWE3NnDI1kKN+QDobnt6cm
qOV30E99USH2Ac7atPa7+OlTA1kNeldMWkTG9o1xDwr8s3uc5YClDh+IV7Y4Q4U1RHySPIyRAu6Z
Gq2fZqHZHLryno7DAtziPIUM7MJoJtI+n91YZt8rp4+/3V8dHNUThu0SrwrUoFZzxQ3LAHMsZGuJ
DVPWNgej88GMuUYcBmtfL5eeUyRBUC7ejQJTsxnJSfEpllyTbTB5umOlnzLXyBA0GmNISz4Anw+z
03wAJH9YknxpZrCpmK1+ZGdeEt9DYhwo0Nb5TrW/+CMimR6QJMExGsJwg5rWAKZ2SRhK4bKlqydg
HgQniRw+5Wg5mUpBr77K6niZdWg8MUMpUg6Yix+I2VEtGZpNQn/vkhvP+T4KEMVkDF1+K7B/oV59
fLRy4qz9i7ayU7vpCVV+pz2eK56duEylZgUf7OK/9y10HaQNcU6QbMmqdQZMf+zaek1F4JaB8Hmx
n6QivmHX4yMUjiWEACEpp0l/RyAaHNDxbTrEEK/PFfH+JBxtH9rAPW5H1cBm5QEkZDnrB64qoppH
jlzGmwWwfUhUWOHbvQSWsUd6WEVrQSgqkCkdC3VczvIkSe02/qibx+RLnLXGoW4K8o0+hYFtvkjP
9BbfGRmYJ4GrT+8K8fiy1lb4yieXOH7tLhlI0dsZGAzSd6hHzSXNgyKwdluHKZTLos4pg4dWpT3G
WG6o0Yv05LMB6pWcuxAbjil5qlO59VosMNaqy96/1XKqXCMf4bkLKC030Fq6u7XehgbMMccEvv2a
O7ZD8jKJWk++zwUIEPMLPwFdy1A7Nm+77wRq6dO4rbWKf3XIoK+EdChvEDDrOCS0a5NEAvkF1T6K
iq/x/XU+8L7zbth25wQVOBM5yMsCxM2bw+DVZpQFKcBHnKfo1mjeeeCiEUuEg9tzkiqBcOMx4wRA
rscHu3bjbGaMhEf4zEhMcSjNu3qgPkqs1nrVTKhSrAmffmZG3McZ464XGRaxl8kcJ/VLkp1/Brsn
daejL2erLD9iq5lvSvLlpAUz9GERVI0Xfs/dHtiAXavvIGp6mbwTkItOvWG3y0bc+8H9kWDpSRBx
n6pWMDqAo8yhP21HkCtXzdKfp3O1fEgPnL2kn2ODWveRNk0ZToYWmVIBwufEa9BFvFGMHv9JzYqS
FMCmtGiuKDFlNoce4THq/f5kWrhvx24kx4fKQcX4Ivcb/LsraKrLbbU273FyfHkP0Al+tOmgL/QN
yvaxq6LtpPl1XsJGfsn9QZkRo6Lc5P8cVcYERdJjegG1h/z3TBS0DPllkPuVDDW6ezt3xwdw2unR
e+TFrgHy7MoIigqSNSEhWItsmYvk5xC4c+pv6canqDea1XtCPh3Hr3eFrEFa9OlzDFgxLstKJM8N
+gH3hPkP546uT62JQFzEj2vccxhx6c33euhaztu8YGOqNkYQaOsPLOn1/jf3oRxS00fOmGPFedtt
sQoaaw91S64E5F2s/xicz2SbrnKYd3yKK0cZ7/P0xmV3ICHQvgX874XMxMQzPIFxZEKZ6Hn1++9Q
PeamnRo0acF8zzl0/l68frdomexKKZhGjHJVXs4tpM5vGyAxDplLyJJwIF/URvcoJWLVFuTc8Uw+
hq5iDbjqZUj/zQj5wxCfOCqfMMZCyOnFbNwEwcIYrwLlCVukJNbsvDkRaotaJWM46B2mEHJ3fBXu
QuLwGG+IvHfnISH9kITmzDu3qRvcRK9u62xNibHy1QmO9DCd1ogAqq6BwIS+sffKWy0q05XvzMH8
Lp4RIsi1f3RjpZbuf0k9zVs8ZaKlXHWjJp0KRXsVF5Tgjs4cbpreNFatTveZR8DUSHMbjr1K0am7
reLCYwHxvXlUZHZPte0wgXAIIwgxHe6/2apcpKhGk8CD53Mw567wpTPN5+MTBhVmUFjo/MDPnWnn
jqv4UTZA2OyOg05uzdP10Cnr9eojSQldcRXvNhNSz2VC4sQGFoan4USDWeG7R0cWw6rP/p8ZsE02
pB3PNjIwhu6Luqztlq3jluadR5Ur9CzZK5TUa1VABRlsKv4EuOTnx/5U464Ur8Mr0E/fsl9p+H6+
IalSek6UOag56/N1Mavb4i+hrR3Jdc4WoeLJApyUYqEhA5nFBtQGbsekO3JX7UlXVAszIxkn3Zsd
wovanOdWDNLmJnpfIX1vTDHfflanjBC+tAWfmPGWirRm86Zs2804Rb4EcyzlDpGvDM7NO+goWa4G
iRQs6Nlm/JpRKx5WQczW2vwZIf20xmYVZII00ovYypaTTMOQpe9FPcOh862Sd1KxKXI38p68VNix
dsd4i3qKXC+C8CSq1FY6hRblQA8YjwRb9iqUPZMBpFI1ujcYW9SYgik3tz6e3z4MYqORdM1uzyz2
L32ekUJctiAy/PBhz5r1hQIzDgROrbIZ7DKlIZmRnPodsByI7Gqi2uZDNLXEzXexGKGvxwxXjPuh
30vuT/63vw6jF8zsMvsAIlkJG8O134mMwoyO3+RPkaqd4fd9ogcgR0MQo1+/dZcmQhmhKhYAlwIr
QAab5cZBWODHXsZrZp/P7DcVPPqWbdYccJtpJD4uYHBv8SlqUBvd4K/fif08oMGc8FfLuxq7U3Mb
pJGVgXPj48ssMYaNYA6CnxySfMWVq+KkBMjUaGB/WMWum5iTtEFWnW/s5XEGibNyMNkORSpd8JN/
FB2QbrWOTTz6wJWdEjNc4DK5brgJDLBu3la0PRxP6HQ3OduJoksYk77qI+juaW4hF/fVRgTZFhZw
Zu50du1CuOX6ntXTJk/nYOLruP5x+C1k+6uwpJaByjryTNLEp5eNQ2DcGggoJeEINamEa5Ya0O6j
RsO+ymRhcUYRNJv5clxD0MPW67Lu90h4c77uxbjSd8HFk5FbZxtyS5DD+Lgzle5mGNlkdnqUuCgT
Z7YwJihkyYb13+GKeRkp3VR1/dr3qQ1IHszU9NbCivze2Pt7M25TBfBVv+PY1IR+GIp6c6Ox7Enk
yQOll/FO7ErCCp3zeO3grlAtNZQcwuWaOKYJe3SND7YuQlSKxLFpdDQBNy2vZLxSXhuFxpoIDpR1
tdh7xoI8fUFhTxzqqjS9OWYCAN54FtIRS1mN7Uylr4mxdyHKdxhH6xQWMsNYdFCYaWkLFO73KRAP
hk4NY4Tkzwp8H2P4VrMHZ8d5Os9GIYuasYXtosnMT2zBC0PYl4UzQj41t0eIUm+BcI3RhV44yAxO
bjRM7Xzas5SX4SxBeapYki7LMC5BttJI+77/Om0h3Jq4Oc5//sjZ836ZGVGF3fy6xgYnL+2lCKFH
48nswKkwSruLKvhMJtHh/7FKedOEXxXLflQ+OuAh3UeKDRGpswaX+oA6WlZC3e5GeSxjO4gW6pe+
ZngXCOgC9uraXrmMDyPr8iWTlaNjjQYPYAwfJUYw/yV0OD0afhSi1COwz8JBZbK3HVNpqy5miqzs
THXa+8AX8xDC0thfDntDegUDhdWGBERFv/GnpFBek/86Lmp6bFZf8o25RqzFpjSmRzABhjFXaP6Y
J1W9OG1IkY8gA06udx5xG4FEWwA68xyD2YYq4iSL7eEvVvpqwdk/Q4Ev/cB0qKbR1VVMHc+OnZxU
cO0YK7G95eNC4eG1pu0qm/CnG1nO0YMJBjDF4wQuMQ3GLkXjEw/AjSpf9GkttUjmu1M+yc3X6fVn
GTG2XxtUnViMr9aQ2Su0kviyq2pTHiPh0T3TlQG7sjHpWoIvLHwCiVDvChfAZkKBjgQw7/UnwKtt
qSHnc9TDn6dlLqHUWo8OSmrZxqLDB3EjeBUfsjIlV1QnzUdyskxNYhYDQAH3f3M5K+NJMW7KsI4A
onCRMX8jZ6YOBS5DbQSxIvVFb5qniYncm2eCWbZmXOMhQuvDw7niX/Y+ghNquOrTkemfba9NLzFD
bZLfUAAHmpVuJ6LuB9wvfbcTdx6Ssr2yykJz1e90V4FDVrxrJBEMNpyCIVmnkcJkNcAwyXU+pmoM
ZvA54P8Q/ny2s1UG7cJP7V91RD6Y0mRCjLay6B5bWFajsvGvTWvCA0Z3L+ZwJssP78J9mmT93Szn
OtTC/f8MwXdv+aVZnOZU4RTOkNSMiDPnhCMy1HE/hx3O/SKFsyyN+C3u81/yLWFga7Ohhh9sqgeg
PwoS8HrXkwCOrJUnuTO1XZ807QvlfPe1Snn5PIwOR5xpiH3rklbZwRIADTIxy82YynZsluEdIE9n
Up6eUh5wadTlhIIO8aNQznRGDXqEPKefEXUSTWQyDC4fQKLxNovcBORr4oDVFD91CjV2jigEPEwi
RO5qKgr6WW6QmccBkveNQw5/bL+ycWjtT04ixHchNS+MW66DH6rLts5KId99ITuZQaunYYagdyKc
Fbr1BE0RrRM+YgAj/I75ls1LjN+8Laa04hIl8ig1rJKSLNAAM4mOGoTpTZQafsspw/RgNtr7qc0J
JB2b4Oj/Cyxpz9DlHRxNcnaKrSg0Qb/nPOhrIRjiY5hOVsVO20+OVD9PImzWgFtTogjvbOubETVe
JEoSfQXynI7Ep1g1CT+Es8zfwAVusJZ2gGuJm1GVIQw40xFcLm5YdGsayO7jg9b/5ayVrAh+V1QA
eidUCbjVyHjwlenTR+eBuVyS2v6vTpx9G7dPJczeq/fY8rI2SLf9VLejEb04vo+2c+ouVEBIsx9H
amO6nYpvAl/ik1Nz1eHcodscMSkvSIocl2C74GKHZ+jENSbb5N91aCWY1mXdp459NaY1FSe+sJ2j
aqZDFTRB7XIhYACIO4Gb/TvwECl/5KAeIGzHT0meLGOl+g9Lo3bpev9v3a6VHzkVRSas1rUJKxpy
5v1h8QcMW6tR1K7xmIfTnuLVcuNjQhHiafEAggBwcFasacXG6kBj3UmPLrEWwTLh0cxkTWSlvtVx
mZgm5wIh/S9hwuDsKUEPT1uMhRRyj2iVAnmAr73Lumg3wFnBTRYt9bYFOMJEORw1+kwH0QcUyaRs
OBCM4LMTga7D5Z1vYC1RMcoeDbzZDpUCk2pkbtNH6ZlJdeLh2HjDrO3mZ7wXPbGEb25Yeo4Ow2FA
eXXG86mQGQMCVFLvNjr4GmGUDJXbTT06Q7boXYdVAcj3ndDChGnfOT+v26MEeCByQhca58y6DD77
oW4coRaOJiwNydmx02sCnK/SPNTQZ3/4V9SSWmYk7PEdLcRcoD5hsA9WcQK324YW91erzBN66oFn
reyfBzEHrfJ32uR5ZsTknskVOQtGHzyhbwnwelvXD5UfXaauC6H/XJ57ZxUQjHoUcNdQ/83PUsm4
DRYj4Y6YYtZV3pgjfO3lTpti7cnc3ZZQVFLd7oIcdC/HdUtn/XdIrOz3sf5px5r586FS4W4ybjlQ
i78al6g9RL5Vt4tgBXEMNEdT9W0TxiMghkZWlyHKgwMcjSRYE1gYcAcxx2MI7zc5cxYQkb5Kgi/T
dw9JRApwOWb9p7MKHJu3KUf/JNSdzRcoTyoaBUFU1cDjx5CWKX8Qvsbvd5PRSG2WU0ru0GT7k5w1
KlVql//zXZ0EKKt8kXkOUZh+XSbEYzdBtWSagvUxnJ65qJcQ3mm2V0l6eYeqPxMZAXY+84Kc6wlV
sQU+juHXRjuUsObAk+s86aB+5i3+XfpLKHj381ULc2an/MCGU2nY11OktRYQ9v6kwc5hXc/H1Y/I
9rExkgWywEihfuZ+GKbVWwvZEGjZ9d2bTk+IBLtTPTCxo8U0iocYEXfwygr1uXXe1p5b+APoQvg5
Q+Pnhft/AyUlggP7gxoj6CJK3NldvMQWD3v3K5jo9KEKJLKUJvTCHvzN6r5xT21V20V15W2mSbTQ
KjWBS6FefSEQPYsws+YWZsFNGpXP3/Mai7F4aXcfLb3CNzajkXcF3+rMJiQ/EmTzdrkp8glabQMf
wpeuoDV9hEX2p3BxmQVtHWemW//ZMRndyiF4SGmMqJi5Di114A7/pGqqy49Ia0/msdCObda/pGBX
3WRYqmxDRSDe19D197ogzJLjotntAKwiJOzOrNG9hbs67WhRNp5x9Gpiev5LqKumTFA8RI2SnRCI
gbQ1q5KNiO7GTR2ca+l+rJSsIC2zb//8pVtuMwNP9FSEu/0TtuJs4EO3cInkDHxNUoBRsSP/XXIK
UV99KAYK5kgL3egsn903KXUaQ399cKFa6sflxWeagx2awRRfToBCs9za4KdLjcxSeHaKl+odkw8k
tUnZE6ZgKzYGo4bWPETJgJzokpJL0gsyonIJbOIipIHOe+CFJQZxyyhc4qbEhdO8s/8LmX1ZwHs6
IXhlKnWSJnPdkUgUgmy73vY1D2XJxW+g8RvQpI5ny90+y8qZiFi7auFSKdkMNhnQqpn6jyCefMMY
dVKNbfaBSgsAa0hJCc1bJhqDgWu7gF7eDt8OAAIPXtxYBSOydv/nwgmt022HNQk0IMj7xQSk9aZx
XgFN6O7APQo5YXU10y7CKcsrkFRGMg7RVDVRxHDg6oNmxW3q8eidA6sq2Rlyxq3losb6pJu1AWuP
f2yWaTI8QtkKfHfjuDlKqnXRZGh1/ol70kqzHgAKyS9uzGg2yI7eFRtAPxAYD8uht0vBiLHId6wL
d96J90ViHmAhYJ4ZT+GMPZ0rJKPJdRBDIBMp1vjj0EHNAqNakZtZg3/4b73hjEWipvATk5RVLkwK
C+UJG6IDA1nadMA/1lqbkupOEtFq6Lbd8Iu/3brk9q31cGzVIhnlBCArhdUNyQhLuuOc8IxaQVSr
1HkarvhYrcDNQqL3h8J9J0/XuAcYQ7Mvjj6oI5fetD9HZblpja/3805qXP4v7AXEGK39/gEJAdd6
wsdF5EFx1/k+SwIgLNbUJCTcC5axAQ68ZOm5zy3rT84d2t+udwwUoBCQyAfCoyeH5frm7DbLHqMf
MGiRlpitYlk4eIcTTlvwobg8ZOUDsJB9iI4hpGwH7a+1RWXMpPmW0YWnSY/02epeSElbrGDvy0jI
GkQR6XBypN6J+PTPuxMWMTW5aHt5O9KUMLiKmVh5hHrRKijABjdn0gH6tkrJsIyfAPH5kcj1sXsd
Jp+12DhE3E26uBH4P4AQNSDu+qBYRl/E2u600YSOYKNH0CXOdYhVcdTWuy/OaNTW0FBUzjbFIyxc
bFVhoFx4RQk/VdXXPl7DDiLdOWuDx/TuJtWTxWfdI+tjUUMFdEWDH2NF6D4rw6dANmbEw3hZNy8s
KuE9hcUC4LIFY17NbN4izoB5WjWZuLTHW3XQ9myeA2akMQuWCgI9jR9GhE/K+5wxxCgOx+PC1PNC
JvoCaul2IvvW0k1col/9ReHJwi2wasYOWYx/p8imgBzmENHc2U02nkcMskLMvOBL0qKFRYjsxiQE
vx5xTtKvQfNEYzmlQz2gn6K4vZ9TOS36ssVs9R2EtePVnYEcXrRD5piTv5jj9ywrhQ0KJF0JiCH0
SuIkdGVBwHOYAKCiGEA7nhgbChfvfdhHpzK5PNb2aXIjUUMGu3dS0YwW17clJiGmZVNBR/i9+ay+
q+RHIaH9N1d28f583fuf8URtOTasrioIWM77ovl08L3UKk7dygctyccIgiWuw5L7Qq4IGVACX646
FT93NivefGUJ7a9ctv43SzEI5/qDwQeLceRDEdJlVlO9sok4SPa1vIinI0Xafu+vw+4/DlSLM4f7
lhcHrFvckxChXORraWO/xHCVqj/9AcS4E3ngOH0Kv+Iu7BvruqT2nI5PfobzlyxAwJ/dNekEBuCV
8JBaa4ONIPN8OryAORlE54c46OBSE6e3Ea1D9z884BClivmg/LTv+0WRas3uheU79Zdn0qVc50bl
i31gClEtO/msdnjlmIUwUiqO0DtKX1REXM7s6pNS/14v3ctiYe3YUw8cJNNX7XGdFU+IYr3H28tm
kWP1kUgya+Rc/2mCKobvD+q0uRl4VDGdjTX1fsXSLlwZacoMVYZA/pS3srq/AzixjZ93/V90rf3h
61Rp8PUWo+wrFi94ALWyiWs9wBNcn8JmCEKmMdSa+bCIeHChIRYafyJwWP1Cl7VAZwDwBU7VInbX
0IeKl0oXMZFdXPfTvX9KUaJoHRILHbB0oJMouqJ/ke30BxvhxxJc2BFOWYUpJWNJ3hP1/ki/hlVU
R40H2P2WbVgNMA6sT1OCg5CV4/yi177/USQVhowFpQ2F0KoVNUZGnr8M8Rp5oFA0RQ+0gUDcpWZO
kqTRL3rGHKSg4zZX+K6YMwzumoA6uIR0LM0hTU011LVmo1xRttNUyaByHmkTW+d/tuTjkbWrJwcn
xtiMcxpCZLzrcrJADaIvirNZqS+8DNo5UHeP9t7FOV1A3RZ1R2mk7ubzn9WZXY+h281On/Dk1mFV
LeKaCxoIa3P8MBXFjZU3sRy5DPQz4EZ9tU4GevRGB4oaas5v0ruPjSi1whKIwXY0IqngIc3SR0Z5
h7fREYNPGO9ov87J4JlNN9ie1Y8FcgXyYmNCNuF5hKiibzK4aXWpGE7yH6SVymV/oODpD9OBu2eV
11msUegOq9fv6wittUukoadyrqR7qRljun9tTZ3M3KZugVq9107A8rV4oNOEBm8FmYm66hvapUq7
RA4vocIAV3DXozOadW8iAo9zcA/SuV1ONFwd4eVL3w72Pe3/wBnzfwltUyBgCC6SU4Ae0nSR+oDj
wJwVR95Q9ZRXGJK5j42S7CGF8UrNuX1Kdq5I8Ekd3DnzzLwyvVs8skuAPPR+Lcchh1nCIIrwbv2p
i/7ZFpji+t+cJXv6tEQL0vmuCQgM391Tg3rYsXcQIZLZfATO/X03OaO2eRFLUMukYzy64lDf1Ol5
ZRhKFOZrF58/j0l4NZVfGywsszNaKSCISNPfFeECcJ615sZI0gCgyYc2ZGrpArCvPdDEGKP9g3KF
Xv0zzSCF8R0yZUaiCDFl0s0KfLJwLaXiQa03otwqWyywUHXrg0/4m9JM0T1lVhW4yKr7tZ2h24WZ
vhx0XByTytgK5B0J5V3wnwaz8KqPZkyO+0HCu6p6b42pQsdYFrCWvO66xSluWXdzgJimHUjvoagT
W7t0zAJtU77FpM4iYBIHg+EkyJmzRa49Z9VJAzas+s8qgsUQFFfbqndgLZzjw4rwievXsnSdfKx/
/H9JkO8WI0i/HxzjjHkCxp7oOLfEGxCXEQwVrjR+zlJQaVk7oH0cZWkNzzySgMUWpDqdmL6YDSWh
hNA2Vq5oLU6trLF7ScY1Im8iP9owCic0HFjkNRy8eEaSHL6OA8NfFrfIDf6b+DTFFrb3tmQPt0zo
AwpwAVPWyOidS4DEn25ARFZMvlnn4Hsd74g4r/k0JKSOAng4fMBf17XaeIETykvxNCEuqIgmESwX
iiF3UHZWBcA9IjkwrvGK9Cl15C4G1iiJsAG/zl1jAKRzk1+CX4XHc/NPQ/6Q3FsnJ7Epn+oCrcMI
HgLfr8Rv7XtRnq/u/4gvVxzbeFO3RkVEDf00Nse8VJMBSenafjSRandQXzD7+qIWzJEnkFUBNPdO
VXdseGec3hBaGXdVzbypB8zhOMdyALJHkYSeHYGQCB0l2i9j4RiNZuQeHS6JHy5C+2p3gokSqlnG
kZzuPjvWvbrXkgzrQ4/OMrFHUkyxPrDapsEsxQlM1MpQObb5roJ1HNwj2YnlUnzP4uU85+REd4zv
cAURdr2RZ/w4L/dsvaSc99NDLuqEAh6xYs/F6ZB7ruIQQj9v18mHQdcjlTgQoUpqBzPBzihS3Phu
9YVDB7gs9c3QJ6KbywD31WclxOssN1ALcbKkAipFmMaR0YXNq1uRK4DlTJcCxA1NEvmXlEjHDDOw
7sYlvEOJFC9ZJitpwLv4xuu+m6wg4/9kQ2j+aZ+vgCffWCDWajfV+TbS+EYBiYRfyaeWPzbLXEjy
hQAjoRsusDRBb7L9dPuzwgadYOC7lEonoirPrs1Y14ms5iiApBmnHRMUJKgCcOCWlnSO8oAWA/vT
3tQkREGBrcZ+kJhMBCBMqvX2bUo2pipc+xQ8mieHsvUDBdRsB+ek93uXGUFzkdYUoPpJ8a0a1sQ8
1M1UOjmgXbtTkWBGTY+s4QVGXQo+gWKlqNHzyrBp5k46oYs3xYITvhDvZPWOJv3wEdyqrL32F2K5
DhfIIxNRGtbrMFntBB3G3YNA9j3pvLOYMpZh6nPAzBl0eeddD2oiyT4062y7W1GffegwmBc5wf0k
TY1GsgepH90k3gJv/wolr12tlUCeW6l7Nu1o9fliOwG8BXpIbiIk6Ehf/aEMGqSw9d2c+1TDwTUC
f9kHNEGAgIbrFWuAwBoOg3DHEGreMAZNNz7CKSC4fUzuOux/guXEzkmcJY7MEVNrNiXvunlFxvv6
Tnyzmljyd/1ODlTke9iUtmlWPwyd1688NlyXFbKs1oeNPMIa/8i1jvhBcG0gZLKAd79qA7URLcUX
i3Iox/0UFujShKp/pkPeSDW9aWFh9WQcG0+Do6DaVsXFhKrF6U/uKxcmCrPSeQ4vO3QQ0oL7nbY3
6lc6X/OUxVKl1T4eEaPg1G2t+3URpPZmXjLGzr2ob/i57aJ4U5xpOi2JY3D/Nld2hZqRYNgwHHuS
5T5xtoR5kGWWrrbbLJ+g4ReofIH/ZsrBhM2G7kMAdJnn+Wyhehxl4WKoj2oMCtR8BOt1eK/aKBXy
T1SWWp3ZLMiSEcVKENjhR3mtg5yeuo7w7u6Uou8cQmgEBEfpzCLjGiJO5J6PGPMvLP9JEomORFQA
yM7gjewOXTsTfBj3F8notYSvxtMBj1RexELl4hcabQUAa6zSCbv7M25vx5sMB5FFVTkceX7Dsbu7
z5TONeUCMuqa9NrBp/kxPJid1MjzXWndzsQM36nKfdWHKj0AkG52V0o+3EYq22FK8UArtt9sORIF
y1SeEqztvrtdq03NF6ZHCZVAcQFX830GFBg4GWPR8tpmHMXK2e5lnyLEXqprF94s0JNCm5qhtwPN
uF7QFTenG2I3KRNpKjMv76xZBZCQ9HVLsONAb9UU2wNYx0HlD/5hkpmn+PRqnZ+4wL4L1j6Xd40L
oVlzYggZt0ADAhrQWMHOM1gLywimIjTR0HUm9yaebpgPM1da8jua9pq6rkD1PWQQavm6KwCnFP4C
DnIcaPhXRbp2zP2smGELaWeThXDEK3ndgbP+NGcgQ5S96xV0IQgHOnQgNwwN59Gsr2QgLhIGTt6L
nKHSLbSanrXfCwq8uHs6LsFwQ6P0+SjnbUYQzvM/irFVkq3KE8IcOrYZhzfwogt9b97v3h/4jNAg
Ey4Uxvbk9nwuz8t5vP3Wsg+slsojbQSJhyQizRzjaEio8p/vRnqtSFFoYEmHn7L5Wb9pcWWijJsE
WWZtlFSpjjeWDfNj2Sf3VItf1M592w6RQyi6g+G6GQg0x/jtGkCMfKrOnOfxr3xelRUTKrbhCCLs
ESsVZvz4/aBj5+SB6KC+m1p42XTeAy4k720IyNIkcvOHluEadNWXnfpgxDM3jHz66FftQSnK+x4X
N53pguNGD9/4vB6WXWWZ2fe3soJey+CRfI4Juk47TFHdg+RG3wrXlDWzgemtwOt+HhZ0Yk0hEAal
EJp0e1gIhPiEZMIWkNybRmrHWm3OoK9gJsyI6YHPGClNwMHYeCDjUDIyPfDJE6+heBPL1RamFA07
kcLyTtlJL+1LwamNnmAmeboujwx7Xwi62Dl8ccyoZkrgW3SIZb9ssr45G+x0dpE4QEACwSXlZmFN
/8QjTMIj9l/ebi601HKpu2sLxjwjyQK8fUhAMz27sfkbG+tJt9Rh1ihS5o9TJeWX1r/NIXCzPThW
8l+Ne+KAQeIS7a6GJ4t4o2Sf2UUF++OnVZ6obmUZWuVLRDQNaD+ZLCCPMy57fs9okAgbu6d9Zj+A
hlHUU5HvfykZnXrl+AB9V9nJW4EvaX6BUPUjr1EYka8Jy3oslgUHtu3xUsKSiPU/CHPV4xQXZoGn
sHV3ujULfp3RNBykOj0+3vnPvGuwgsUtDX0E9IXI6Vs59mAj03Wm4x8XCNYIuh1uOj0jT0Q1qiqi
hQP5beJ8FCN1GxlDaYx0fBityAa+YzEM3tO4t+KHghRf6tnj8g9mM716dLmeGfOGtiYipVKMPAhx
DaQpiXETHQUnzTw2v225pUo6vLaXraT2A+og9YsyYZS9U4PPefiqycVYNc541sLiPZB6TLtWIi4U
+CdKM1g8H16+QjDTRBQSBeY5hDMqLE68U3SeoeTKqBWvhPxSYxwzDrBs++9ijdO/pS76ltuTXzHJ
tlWXbDID0YZFvo3tzRvY7mEQVeAIOuo5IIGBE0USILUWXiKCK/7jDrp5xC/m6A9zh6lY/IrEmtcL
MPSTq2km2vbDaBE9xdDIkBOuFLyoGQpbryYdygNb9GJ3EUw0Erw9EiEAkC8iFPQlAm+kCCv69Ium
rDU3jjwvc2sFyziPhetygZVP7molKvEaMyUXd8IUsDUOkrzx6kzyYHHyTZMCILmPtqkP0f3h8K3A
hMmTN6F9w9p87AT0mUFV+VRA0UrK3jb3lNPX6TGEFMOBVrD3mO4+6lXNLGDdSOtb1lWoekXnma21
mzYdSxEKV3Ym4qerRtyZL7KrImwphRTtbsRIAdog5MUAalE99sGg8Ffhl+5iAJZ6li2Q4sbAfVch
pOkt96R8Dm5eyT0YKiDWntl4spnSUPZn7K9GnBv/yvmBDz0mrfiB+UunM4M+hA9b1L+8d2nC+Ld1
i6EwKZ1DlaSunBIUbZfo+zk9MQ9mu2sI1ym9rD2FamfQvDsDsEfBd62XjWwPS2GiwMiialGf26BV
F3icQbA+txB3Rz6qfqFFvUzIi+F8LyMXiQlCzh4WmX1Dav5qbs8cdWnIZdzub3P+CiLsPBEnqvKm
1kwMNO0Gafb1We7AgRdSvX/bUlF+gPI/NZKmRsSIthUlLkYQCNqEYxE/qwrtOo/1hELm3N33Nl8v
sqFEopw3EoqrNeUgQUOnyAwChaBEV+DwXATqATkwpb2lwS4NYy8kcvdSwmeJhz0272VSSNUfnUWJ
+mj9F3yt2NJs7stRp9yif2WAkys05DaaYpwwUKNTf8JhrSZxdATxMlYoJsMF60BAP8/w5lOXI02v
uthA4qSlbk/QpiHlvi/fpGmgCl41/9FlrXmJBbUyrJER6FcrIlDMT03LCcvdcIYA8cCNdBLtdhan
vTJ85i0yydyULY11go0EehRFpwZU5keGnl3kXtFgaczhSJ3l1Zh0SHinvoVM7hbT5SasgvfNxref
Nj30+vwra55L7zZiQlO6dnF8MjjgVKa1/fKtIe9WLbI32RGiNiCwMIKBGXw16QoGWBRcqPuXsjnk
5MpXdMbgtXWidh5r2ahlgJPppqAiRVMv/+XAhqa7szfx1A0JHTVWu1nt8v9zU57wNuI/cGEc7vSA
7XPv0Ix7/BeodauxyZ0T2VvsQrP7Np9C8XWLgQxZB3113/9wFA2XywJdfjC/VSr3K+CZP6HRh1s2
fpYZgFTKdLFWo+ShPD6vbph304QRWmdkQVJcPzCQvHcMP21peLmOYNJfQcfGyi3OqvAQY9FpExp6
4epsQb06V7sViJfmtdBvXeFkG7Qxo18szQB4q9St9NQod9N6+6FznyQGhRGP5U9OP91TqBqbFNAU
0D0c3p0JbQzDydo3Xbcf1Vn7/dIbcZ9rdL3IyBgik+CQ5j188GqpzrDcV/JDxEE4OayZIxjBk+V1
HZ75TeBy+SNgYmEOXrwwuEqGPUpOaxBlXrASwvZlMdAMC+NdqdqzUlyIpBeq6xyFzloeKT//gY5v
tyWxaFLhxpCk0HjAoPuCYNWM5PnCN3ghuiI1xnYfmPbJ2faTKsD2Cca0/zFD2opGCmctlndfhGXr
/xxJtEYQoOO6OvqnIOluM2AdyNLRzl3MfWIRNtQqbYP2qihO+4LfLsz/LtFQZ5dFY8J6jGCO+bGr
tb+P+vO37zo8Bw9VEDqOT+W1Z1ATvkoBuvIQaGB4R57NNYMYphEbbKHyzJC3R3WT/JhAsW82Y4py
TposXb9zHnaVWarLocMuj7Tu4GYyZXPpiKltyFT7k1NX8YADA6S2sqsi6YU4zMJNEFuYNYwAk7Vf
jOSeqIpupXEtVuOlZiHcv3EJpKZxS3AV5+OkxpCd0a6uh/gbUicnzUyP1AcsFP4zI/KtHIKC0256
ABDoAVS9pWFAqBsdUk7JhXxjCLm3rO1lQ4NHoEWiiC70fzYXnJAMdciSexMfjIYBk2nM5aFqqw9q
ADvqMOXMnglLUBHV1oWPx+ubOoBm/N0VPwnfwIsZ0sCP7873WbuW0BaNu3t5P+Vzl1Tf+FWtVt6R
+tM1RkYcdSKaZCW3OHQQnb1nRNV8BExC9XRMs36X/Iv2gH6taCM30ryOQwRbhN0RvezilDwdA16A
tCfLjbzJaPVEwUeZda0zwA3p/yIQz7oZ4w9azVa+O3atFUh0piu85Ta6EG10QW0BHsQDdcYgq3aw
/HiRgVyrFDyrJxVgAwFqc8NhGHTXw4OtfUZ22QhNgi9eTcfhESI+BYoiPiUY5PYYaxKhaeUeJnKh
tDYaHM5ROmSxkw5/9+YFgchjJVlVwRMmttKypfBulnUaEfAvoBOG1PoJinWF7qWMUKhYznRkklpD
dd3jdWExM59X8nUVLGmUNuWeGRGyXmrvowHXvnS5WWsqQZxpGASQ9xU9rgz2l6AA01505PHYyCdr
rk7q+zIoekYAH0nY6oiJgOTG/ghiN1MftzjESIsjJdeYCbEoZW0tbXjnl+jNQ7i1kL9c8CjtZyL2
OlLgG1RGRQcoW7KK28q5rMOCPCgderfldDxIr1jTDpH1U1MXu7r27ghwVqug+DgwW4IByXt4ZH1Q
jOgKu71sdmFGWrQL+FwEDgdzNfLPsObPcVX8LLI8zJP57OF0G2O5CODJyI1O0GW6f5EibrztYUsH
G7t44UfNlJchDfdGmCiy7Mgfxdc04fi8li9ww4eaDKgLbe34WDkYPOAvmeM5Rc9oU9yl9C8eKnXc
VlqwqDVW6AS7m4C3931wMkJKN+QolxSd+6DzWg7s24pYtqhrIKzoxFdR/KS/OqgypCMWQ24lMtBt
l9RuwcqTLSlsGrOuqdSOiY5vx4a4J7akx19lUGE3ChnYy2J7MCqJBi0ZFIDjbBbeFSFw/xMMlKEh
VQtkd9uRUlipxvEAHrVFj81VCFSwbU+KQNM01q4HyYh/c3pyF44OHftViJfJkE1XgUm9keRoO4EC
LQUc3HnLyspsE4Je6qMFR/tX/1Agz+RhzHB1TA8QPTPlUXgZYQukFeBGoVFscTPck5SPyfrCTuFe
gyVZ6DFvCISe4Aw1enRE1Mn10qiMWnBk+IOmjG17i5t2GYBhbKVI1+d6DUDXw4Q5nrcfmhGzicCy
TIRu5RC+8f4Bo8WZxl6yiCgkA3et9S3GlXdepZLHOl1SsbGCK7xFHhqoG2WBGgZDmv6nPfoTZJju
TK/Oq+ZNA6NOm1d1qO3O4SBW6IWJHuYCq5aNQ3yg0UFJE9AtcaZQhK40bYJOikkRL4E1ZeU32yen
4eqDyMtDudFjUwRtZ6WlzRM8ujLOAShTd/g2v0VpY65BApkum311t5auff1+7tXnMO0A5y82/wve
oUAe253PjkuksnL4deXJ108Ni/mUOkOak/l5BSLEtauLM9Ybh85z+UBYWxAC3Q+UZvavAZOxRDtz
EzJ6dG8byqsLtpbGFsbuRsUvH57VslHYNzFlhcxtO0T104qspzngZyBsrkEbmrA0YN37h/5OsVp1
15EDgeLW5B5RWfTSEixaGhoIyRrXwrONUUHH101PE1xWn5jYZSgqEdSWYXCgufhkT9rJJT3MtMe1
tWb4HvgAli1+hAlp1/ieWAgjI2/RVMUcdmA91at0u7GrvEO+g5fRotNNku1FwYwGEDIgEBE2oww9
f2pc0/Psl6/08fmQK+xPy6rIBS8LREVQ1MZQf1voAU2+ETMA2i+C0ePnJNqqjdFoDhamc+8UEbj2
GHRYZwc9avEoqh7ULCFue8WdZtBh8iaF5lJsnuokBSexTLXeS+PvAWkZAjpkZgS8uj6xs2r16Og4
4hvx8I9mNm4HklS9aCqWJmkFm01MibmGaLdZqJSj428wofBX0nIpNP3SMBqI1pG+XlryNzCvfcvH
J4dSye4C0pnbmWInQpqmJBX+jQuHOqt/+WmRydwi+5MBWVRbzid646wzt0/Jvjh/HEjWUzojfW9f
/XBSexOXIb5YoS0XUgRYRC48ZCrAGyAVRn+JrE8VmSfx20myboN9L9WadP2R2DaIcSXPIVUJNhT/
wt+3PSRQ3GevyER71P8YqyZTa57M1ogTWUssYI2uoJoAxRE1X8890VGQBuE3UnIZe6lJN6IIvnjt
yagB9h0aeYlVBG/wbh39MoL+CWzDF0f0UTxfVZ1WEBpwoCJt2gPqRs5KK9ZmnAVyYeq4dOyAnxoJ
FBi+ZRhFiYNanLEQZ2PJxFfU0mrJfD3mlVyTNzyeIgLfmVHsYQSHvE+8wjMKie++gU9BCjgXzqs+
aRqnbnLjNQH+yzFjcBh1i/HiTvbyoCeJBC+4JTzU4kfBdwBuFJQrY2HbF95IDyU8BgI64FuccwDm
SG38R1X1AtWFkjdy28f17dlDz9p44QfgbZ2ZTgpbceJ5HcEGNIseD0k3xMMn2LTBa4WAjcco2JT7
YlNm4kNBdlcuHMMBOM5A5eChYBBaxXjyN8+enp5JSDlz11KVkIT51xTIf4FOJp/OpUKVo6S9Jdmr
f/Rp8Caq92geYP1peobbR/IwM81nNxQVXfcI/nIUduYLnL7kvXnjd37GxyQvSENBZptQaFKf1DsK
SN/TAwG05+FkGNhpqX5Ca9cxSGpO/xVr3PCUnK62zAFbyCMXU0E/lByv4wxSZuLrzg7fZUm6TUHD
txXv3xhVubVdtq0EbpkMSHC3LADP5pKzIcXnicmb+yOyoIsFfChXFam9a6zsjG9o0TQiBTrISARz
+iEKdEvqN4jxHrxEjkJASDkN5e8PTLBae2ED+HDx89f5q5INr9VUagku1I4Fq2OYmQexkBqbvi0Y
aXiVNSDwXFdr497mRuM4MBtaSARzej8tNWvg2OmvBh+6JH5Rt7q2XqZPxWOhz8BTlemY45WYhqjK
aArgE4iensxz6AXIeumZzG1D51cjh3aCFvqyi+gTLOk+tR5hCGMGtgqDnJb43/fCp0OhOZFoiXLm
NXNs8Yw/nWG7Yj0GPirgQLwzzg3cb+sgFR4uuPN1Yn1CksThrQMPKHWm+I3Kebyf1AWyt/O19cCO
HCmAyKx40K8MhbzlxX/nJdG9QqC4ei45KjfrVffPHC2hW7mWEHkSPzHXunfMsLo1zP8iG/Q7UCs9
JoH/FHC6BziQcMecUYFnZcTJC5CDvZNlMkl2WTbxD7Bh94iaf45WIgzUtWsjFJ+Qn6E68YQITKVS
vJrCWgr/r174/d62EoL3Lb3uqDkYPu0ytKP2MQBXZkwtFUpx8QX5h0nQh+H8fJAtHHr4NGHHC447
T/IwLxmh4V8mY8l+KXTe6ahWOrl9ldhOi9Bubm1J4vgT2ex3Czv8ReJl79zlvpVI5QKqrLpbr+Td
pfMQmA0WWJeT5KOYpy68pSBOAnW21o41n+uxZoL7GOSSRnM8S6vYbHD9kSO/rzjE2NVXe0TtWGBj
vjbUF1peLsbPfk8lMTakJDkZ0HPgCUvpzntkplYnrJxeww9L/QaCYSzKMCeY6OeonuIh918St13b
qS2JZmgADNmvWIIWSrRGlJRTm1N8x5vKs65Zu6DS08x/GdJr4urS9TOh2pZr1Nwj4mhD2b3EY0eZ
RwvTfZcr74Wd1QpaJxwpKJbERnIXF9pDAFZve9H+foMv7wjXQR7UyIK4cjOaFH4GhDXWz68fOalR
8E327I0s1p7Yt7TLuXGePpFXmVY2Wr6sn92BBvz6PARZ6Z4yijUCdR0vVgQ/InOyYWhHWPcPvbSm
EeGgrPF7qVNvOmKUYKmDKKIKH7q8dI8cnB37yFPAhinEMKLLGHvIQsmZMiRDa0zXxNiSJ5yD1VIa
Qhsi0onPJ1iP4lIbhT+Ix+Yfb5mVat62KLwKzOI5P9G0+R+epTMwm91tFZR9FQE2W/unSXPlMcrN
5JagSSZEFGRaCyoW2aJ8J+8EMap38nhQNLI+KFiZmLHWWCU7f60m4tpu4YgCFE9WY6v3h9K9Vezv
4fq0wGisdYUEf0K3LMk8/zfcUy5Hd7AKbWkC/OrDIlJuNqd88dp374rB25NUkiAWu8TDcMgPlw6K
4leDUfrtYAjNp8kPVBIKviHn2LQ9HE2ToVJAYf2RS+x23OsSMYXbfBY5EnKDn9PbV0XHon0SOTQX
q13D2v27ZHR0TO/Ov3Zacek1lcEjYCgWnvgYm/kSNNYbrn5tz9ndM7KIvuSZlD9K0bWxBBBA0W8E
KqZwo5NYajzpxq3tYuV2apBAsd8rzLaVMwFKSWhAK2VIt1UHYxuqUwYw25m37o3VWNvo5GlNhu3Z
hC48/YHaL4uI9dBUVSUPJ0v9BVyBsVlhZLFP50fHOOcLZaWA5eaaBZbvNV2Z+pDpSDUWPlN7YvSL
gSw3EfwoO96ICIOnMGhTZXxxXil/qfJs4kXsYCeGG1wUOH7uiYPIcC3BtYEbFN4tIhnsDpO3trX3
Gchk8ZYSUYCuO0ELd7GEV9c44Plh+9GTyTneQbKjlGkE1yg3AyuhWY8M3IftM6UXvhE9kzUaZ5fV
a1og2YjGaJaFOjS58mOzHhTVZ6P59QNoCa/RMdN9PqYAHHMxGAxlBaD+6o/OIkemLuPkK5cyFPHi
j0fSDMErZQ3TOa/+K0iJuE+oEIYRnA/s02/5+zemHMoGgoVrLu+cKfYic/CAqlhdqQ5ve73EiWT+
15WWXITZOOoWIerIzfWR45hg/ItznTx0Dxvp2q/ChpSxER2dfPTjoGC5HHKqwfzD6Vp0aGvd8//Z
Ep1sR6Iwlt1UrfPF6Cd/o1JGJblTUFP7vHiYR6AhaVt/tP1axF2Xfu/+bRt02MNhZFksxdCtJDrW
Ar/dEQmDUhazKYDtLDDIVdUU5PDgMxHghK5q11LApfUBmm3as+brw1n6PZoF8r+HYfF5MxeU0aGq
UKKMWz2XNo3eFg6jiH9y2wf5iYetlLsf8Zhss2XcDBNSpW2CvXLZrutX8pM5gCI6y/qE9KHe3foB
w6Fok84gVGQ2+R9BjTBe2DP0xZ6NS0G1OeH4lY7tYBXKTz868IhOlQWT9qKXC5uGH7QFY6ZFQsrP
kLLvr4DoYkH/PYA6Zk0lc9kSDdlRgNotT2Xn3GI703afERd+27/icT9ZYAhre52mm2m+8yOGYEXB
xGQValUVtf674e/6QVupwpzGfOkOhJmATezGfunwSXEq5mVAtKa9MCW5c8f7hBCsLiDJ4TNzHqee
FH3OHWE9tq92hPGuUg37Q1v8gaaAx/s2Lpp8z55+79PIJ85LD4dHe7XiXgviwokAVw0RrmNpoOR3
1sZkQfkoGRgh2y42tsbiaHeaD5vFJi2d8IThXTGTFhcrJd2A0OZv821tHYp6qdWdJPAuH5Nnur7N
01GAMR+J1UDD+0p8p1ttrzK1IstmwVNIe/uJjwZGHsMS3A/FX71iOjMeXJDqdHip7j81uKXHrFc0
gDbxPjh47gOnaQZlQpqMGaDwW+XGJBjrMms/uKiV6tlAqB3tjngchU7wmQvjKAywQ+ayv48n1H/X
ZpmI2stRF8cDUf4CpizODgLHDG4XL74Uu0ok9aosVtJ5TLWr5Xr9zeRMlTEaN4MBtyQ32GO9vL1L
HbxttRLBPKj3sRPG9rbM5UHFP+ChR0fkF/nPAYFxWc5PtvO5dqGAF3SQFr89ZVLgDBKA4mZ/v9p5
6HPEcLy03shfVgzIQdiJDLKJHAsMWr9vC5rbHzKK/SPZ4KPFd+r3QSzOkLwiUuZ5c1ra7H8AFepJ
AxPl9dEJ9krIqzMt3EBTU8DRXgb/XahMbsJii0+NFiLCWZd/XCV4qOUAQdCio/LrkrumXmN/tm72
ugFXrFQ1//Xx75ua7WqVn+PzYbFtMiMz0kqY3IbDjJyMwGc6phE4+5sqpAisTLlpzA2TdzjVhdFw
b9nvC/nw+ld1rWiOttiO+h4cJ8dKHJd04Cw07Ql+BatLO/noTlrq48xl5BOKKTSoaNn1JYe2BtwV
mGaHlcgprtcHXkEoebttL3jsDdarEc9cdiddsuDx8mpTxdMKGQ3pwRJOsbanf+5OTF4x5Hn8Tceb
GY1C/v+KUYSYFgUD/n8J/SH1e2r2urh26dFhwwNZbcIESRIQ+vdsIzHxEozQd7flRJl/7a5wIx9z
SBPAzCmQNhN8pCUWkZsD+0DE5A1syG8R93Et2iDzGRYchjkjTx0Ib+xAmjg+Kns45Ncoiyi23LHs
cH89kLAh+j86Rb0syXjUcx0a79L1XvUNX1PHLJsSZvwvc8R/0gsiuQDN+K3RkYdClPj6sHw1nP6c
NLi0RFnKam7waOhjvlSZXFS1nzzRibgoGSRYXYMB/fJ6j4WxfdI88a+2Sy4gsco7tYzZ4hrkAfEA
VQXBEurdv1N5P2hVwQYnpcNdOUR2aV7aZPbmOkdIG8hiaubn17jjBiBxGFZkVfin9g+qLcYnfibw
RAufC3WjTlrUk+wiJu1aSdt6Q9+pG7fa/PREqrXjmMMu1TTry1kn05JhOLwC7gfRPqYesgFRWvz9
i3WEcoqhdkT2uym2P+mFJvlPQG7uku9sPXJ9aFrKyLQ/ueoORgbOnp7+pb4hIuR0Efu+cS9Z/EVz
No3V+yljLElP/5f8vlvYR/w4xgYim1XnCZ5bYv95f1A6DtZJ/l3KBHRclfBK9VeYl2RqJ4rbmloT
18fVzRAxZFq4Gtvw87pWa9abh6brrbuPJFroiMksHI2zhYehEstWh4MLm5KzMX8loGGA3p9HfI2C
AfeYfkhg6pWgAtcFAl9aZXG0sr43UKgSMgmXUVFtSohAnWhVIsre7/xbOeTXQUWEDePB4xmIPujK
BYM6Rj1BviO3r/55c28tqfYLSaGHpRA57wxKaMfmGYK4aAoCxfI3WrrzmwHGW8udpmAEqfkqTOOC
dMl5JL5rztZUUjn9L8yxMnQTTynyg9k+EXGDUjAHExKCtl8Uezwaofp/qBjo41NeMApdGzKd0GFo
Xyb5XW+hn5QxVLjJvjZJZ5ojEDho/TnaFm1BwN/CzPVtJC26KNTIzU8i+mMG2D17HGyiu7gls8wq
X15TCO1fJeKUkFWLKMWAI9ZfATuqnRZkduZWCKVdTEaWzvZjSnfHaC/9kByqE/2YXM9A+edROahT
0rV2g3VSPSpuI+M2lAoX8eayOFXXJXMOoFZLPlWsMpbchqlVm+AU9PKWsTR/iXntnIpa4kcRZ6eX
IsqVUlTlSoV4wAb83pYl1jLWHeJ58BvGmCR+yDhg2YvlQmRnw7Z/hwy4DR3o83RpZUpg9Si3ufRb
IwBqNPjqOu/OSe0KAUpMjdr1M5U45WDUMJJIinwNbg2frbovTtVNDA9esLw/y2RULBuNiWw4U3Xf
QoQsew5B7amkR0Om3R67RdjNY+DCSXhl31UBAC236WBPdbWaZFf1LIducBWQgF2pRHUznpy5Oq3j
8/PU/oKjB67TOOJzKUBmp9Tdy9oW7ZJTUGMxNqEErLFKDnZ/sWMiZguOb4Y7/9ferBCVJzcvnXvu
FJZSj+EKJ+8DEZ50s2gbKqT+Jp28o3DkUyn7CSYHnkqmGBbO+ompA28y0t32IhdOk1nROU2cQMgi
zF9fqBdoQWOJ2rm4a7V0nedHgK+ZRQ9F3V08eIz0vbxMJ3Ak3OC2IaMUxPoOzR8HGHWalyHlfAHf
Ukbt/aZaVDUZumj60IhwLYRiVD8JN+fb0taRB5bIz1xX5zp9A3+nDRYhF6ChE7Slgjdd8DI+wI3W
SWGKpqdSQO/xN2a4dk9PF7ELZEvJVcGCVt7wH1+Eg07HPGRZBEAxEtDWwywYn6UJkpNBVajFy4TQ
owbWZFXPwvgPEF2bDYbwq54XblSv43m7e4XbEMIRnCyDQK40kMdeOFNb3rUDsFgsjRByOQ+2OZg+
27u95aUs7uEJCmEsNkKIIZuN10ZqwNtmNKj4c7gCsyCbw1+DWzuEUtSl+LCEFBIVkFEEMoNDQl/S
PV174vOzpX+tXwHq3uF1a/zl9gAx2OKpL11Hlb/17tpy6QaaobiOSbN1i8FVw9eYpIiPSLh+sF+r
mf12YB+yswY/sDlpuA8UjUTI6VhzCGABH4BQrNkPmV9ysv6WcaQuVN9+IwKjlZJ1VxM+/X5RZfWp
RD3wHAaHIVWztqRQvCkELoGdyo9IuyKRA2SuNLTsQkqvCVemHamLY+umpzUhAnFnBACZbMTzFWjT
sM+GlZ8PbmnBBi0Q2z2ZjlvQ9uF5fDOvFceSRhF7Sf9SwhmcqvjNgXlLz7XERCpJ7G31lk+CpNpS
zLHGoq6KcmwF2mYCZMXOJtiEt+looI8oqVYknLBR4nkvgvWfq6fHt2bYkJl1c+T1I9pBME/lSjf0
dqWIgluMnHaQ5EHET5949eS/6oRl+sxqVk6rIXzrvbZW1Nrcbb/ByrawK9N/CD7r8Pnb8DK2kzeS
zLabzTSB+CBRL+GIUPreSvjNU5ECyprA/1I7QZHd1NnvRbtMNSeL5MwCwEkH22MBqNF24xpKQbZb
szlSu932awNa94SmpjQNBrGsYiKvVSLEQrZh5EZsxf8OGRnUEgcMnjUK2x/OgkGAQqUXGzLv/GMp
4SVS1hn1LB002uT1XETdWhCTs7Sa6qQGoD46ZdXVMh2PcyPUMsU5fhQUubst6diJP51iGUfCOhTI
PGjuKuRBQKwnLQRDNt2enItYWaVpUemgwobqQ51C6Sv/4j/SsvzdOEkgAMH5DvjlSd9teKAp0dxs
e6IvBaXl482Yi9jScolzuAhJKzt5InK2SzdHuMgn0nzBN/1w4Hxr1R7vFv3aCh2DmgVhPdLynunR
IE3ztvljDU8GpgD9qdNfmq3c3vpaOwGKEoM8NJPtQJbbxmoNkUNmLRXzxgXgpnwrbXb8yYW4VZAo
knmUPLjKYi6ROn0kD0p02EqF1xDXZr3D/VpSnAwllRzE2CVfoxQyKUmGRHhIfrJisjdl2w4SwE7+
UG2r+4hHobnoXPfK6zpJmsIHUhpcGMlsb4TP8vCecLoic5nwJ1Ze++5/t70gpyjFwuZ8a4gXD7jL
vwJDz97CKJCZHs/VovU539TTNL8AORVoU/gbX6YBOsxkeIBUSX3mNTqm3VoyB1rMHv+UqQfHLjoW
3S+NCwFFbD0pSnfeCEnT1Q57+NHauUdpMNewf4HpL27PT8QA1FZ7ypzZe3m1Hn3ZE4RCp+ydOAhl
48vVBO12uA0+HlvDDtnmNempMOOCc63sVL9Y2fUjBBoJrvUWuGlN+Z6bvo7qrxnWfkOwrxPIaJBc
7ijFCc73ZVtZblFbFR0vr9Nz4Ggs9H+J/mnjloLUcyenlq/M9BWArN3WP32i8jcgoYZArBQrVMLB
ucR4V3U40knNFVHmFfxckBZZvxJRGZt4VOEvAYvTjoOlU2huU0Q8n6OpxAtS9wd8R/LDfGSs7O//
9FKMf6MPg1N5q3EYbwhqfk2jYTkI/NlZ3g6dlG5vaz84qTSuZIkRbpVoDow9rtWv/EHOqolCXhrv
0hdt9Tw6g+WEw2IeYFUKCJGRhR5mjmpfeat+ttcJrGBR6hzq4uPAaH08jZbgFFJ5nsyoYAGI/b2I
rCrnaTaoWTANrR9c5Pt3xGqdZCKWtIV/b4BZqEgkHSmWhHpHevSY/PC8oMU1z5j2wKfgwQmKg09u
x24Q1Gdnle6aHZ3JnkHR194TLe1dgCiuYP4fSJll0ABicKH1SGHUil/dHtqtAYQZbL201Cv/c1Mu
Yox2c9GvtuqgjuMRebaA7/ro1sxQMtZsC9KhJ0QYWiXm5Z9j4aIdzzt+e8HO+/gmYlkaK+1nV7hw
4cWlbEhom1Tc7C5QQkNRHu3MzaSpHmNk97paZwupEGf7LaYZYtQ9fcE1mFThzm904GNXOqUMcCuE
rKdlQ2VzasRFCgiDXaZrRLyKZIcIYp7cYSsZiRlOT6VxyleE/HwAz9vwiAV3qB8BmI+iP0TFDnPv
MawSUskjioKzvsNY+2sLlna7novI+DHFoetuFaQ5L1W/CvLqx4NZGpcyGgT+oStLAWsbV0xO8Kff
cvvXkX9KU7xxWClM4LmpUVSGpfigL4M+LqBaVkFj+FBX/irTm3zLR1tc1MzGph67AMau51SW4J6S
dByR5hi38YR4kUEIoPcFrwZ7k+JSrie8wSxmcHjDqvnKyx22jsI6Z4G4BPEILAsxd59K9YzvUf+N
Jg3ASMac9JOoommSX1C1qKSMP5l0zj2M2aUSrhjU3iiFdn2ffflODxyBrhK2XIuAmGVCI4wVwe1l
+OaGl7nA3t99Z4cCWTNjPLfVAV9YUuL8ZJoB+aMzKBkLhUGgGxF4jIqeZiXxm8GmdELGy2tJOu0e
0EycNkkmttowiRopPH1XrdaGUhO8nR1WkyvkUvrsJbgxjRIPCQPF/5KQNjzewKuQ8TKG9jigUKXJ
YTmZ/CRVj/nGhKz1aa54I1V5hLY8FbmgqU3Mkiopz3nF9yU7bhXAn3TJphD6a/OmsShidWLIlXQM
AGYqCBUw9fjecBrLTtbdQnWrHmXBECCeofKdEuDotjM0nB1LuS2vB/Se2vbei5qwWvuLpRzw98jz
rMnrKuzKnxJkdjfQ5FfBE1YrH5o3ocY5d2t2Ue27zy5EQsmXObZxHesrfYfiVaiaCwTFk7xji9sB
hdjgMpnzHU22/WwedCOdPkWvJbVNLbTPfHxNz/k23oDJj+vfF/3jJXcj0zonXZJYqsYR1dKCz7u7
9g94V82pXZPdyV08sNsWA7/SN2gYg2a3aNA487eXcGgAg+coxUfdd8Yf84AGJ7tlTdVebjlOiXmf
+8CqjJO9bABE2bzpO0mH+Yr2IHj3c0BlGk7v57WcfpXsglzLCqeAZor2Pkey0Qa6w0k4BSEnhDEC
j96Zxevzk+b+R/KS+SNGzCqYPAhlZGBydrt6BGfyhPuPIM1/uSW+2ZTHHBanNwfH1Lw3bOCS4T2r
2CGpAfWP7M6bvKNRa+29C89HPBuiWCLZczXaHfz6m/gFaSoAUJhaZ5bCzd+Y/poNFHSD+SJUJLk5
yqJN4XbnnvjoJ8nuP96MdOPNYzbVutI02OHsBRdP6tFOj9hQQG/F3+MF+HsjfZ1CsjnD8V1dpDa1
NW73V56fcZL55OU6kF3KzOktjzsqHxdATgbiijbTCT1dIe0SKoscIwRpgXxBz/htfO7xGYz8NTJf
3oPzgYOG/UrVVNd9scK07euFf24GrjPEgzwCl00Nb0dXirsfq2XPKNnDKjJAYHV48SeUyZ5lgj5q
nRnzi+7XQVvalv7DLBayOMNJ055zwJ3Q+lhImFBa/duU0qRQij0iu5Ay6GdESqkATAx8e0dFdljo
pJ+B2lLy+NIMMjqSL5wiF+S/+BpdY9NfswcWvkUBKemYkUK6n7MLHIJ8A/6KjY8DINN6j3OqJiiq
SR2QVmuCA4FtqduDkawuSqGi+K6tY4nGIW7mSIx58ZEBfjaAlsAcFECm7b15kgnWxbwVuFMl2TLR
MjYjrTDfggEPEMF7ln39/VlPpaHuH/csMhAQ97X8e/L24fyJjSoJFGt3izUY/uwCYsF/9zmhM3QN
+HT2OsVs/wIYayEkY9w62DPpnbJz+umw1APbAGHcovFRIhsmQP91GOOE+Z0noaEZPJvUgZWCDwpo
Thv+/EyxCwhVCewlHU36Eh889t8GxmyCW9K/p1EWzPP8X3MU35UkKvUtHjUt+RfiMO60dF94yBv9
gS6XKtdh9bis0R02to2f8y1HRqLWSrYwdzANXkWLrqz1h3PPGz+euW5ua62f01i6rcckGWdcF9eE
JKNgnv/RvazyKuv5Ql6fLOboMgBFWT+gymI64576mx3fOlQEOtNA8Bk6n6+4MvUWuSpNXNsiin8k
HuK5cOC8TpXyHV4UJOzOXKzGTVS0CxZ1xGfK06Fc2AJmr8NxdpAn84Ugs2SboPIzWzTUajtff1ja
kuzO7DMjWHiHdWeF6Chh82ggxQkPy58PpqKGakbb1CdDl0ovK65vNO8g45c7b4Z1lyfrtlikuy3I
MTTqPuEHNGy7ImIS9KCqPK4vXBuAEUwCv6oZs9p9z5h+vgRsXrED3bomVsU0oAUn9/1tFQew3E3t
G8eDZeDzbUvJjT3MS6LZM0FxPSpvxJ1q1JEKrLit3QWTtCtbubjWk+e2ywszjjVvFuUi4U+eVPaX
4Z629bQ+tdbegk6VuzCJ3PORCefc2SVC1U7VjnfNO6fxbLTK4PQh0lCejwn1tQ4BeZClOcKLxx0O
UMYw0jte4zDFXhb6wRd/0LDEwO+UTe6j6y1kiVkGLTDlnkB7tKqiGLDw/dxBkrdZ/pem11BcOs95
PAbbcS20+I0n06AqIPcAYbQ/vgp5/Q4ygae1VMKJv3+HGxLJvrLGpxauoaMbpQJKmyHa3c5WqijF
YitX/ln/ikBU2/ea16+dyz6teJmftWjuLd6tCWj9Ca0sy92pooRyRTl/CnCfiA+/y8iajCzLoSv1
Yyj7KkwQdsJcobTFG1L9+vS7jf6ZKFPK+7OOtaQU+IaXBjR7YSeD5flGbuIaLBmB+cIrW5rVDdGL
K+pmreDsL2PqOwsnC5Z/J2z8oIXhujo6g7dKGS5g3dKT/AkRL8F1zznTOWnOCuvUJpgrcI5j/i7Z
nCDuhgAFsMhV8V+NSzVLlmnBGH5OEBdrnRPHeFdqGUaSIr3Zg5KwJ24VngcL6N/tkGOCsdTrTnio
7deuBDKMPtYtRF+G5FxDXV/c/hQQGskWKEZS8PDwGNGOijgQJO9Zne3Nxngjy6SgZewjWRPk5wzv
kt4JsDJFzpuKCPE7+vZFd++c/6rSo1TOW8GrmUSdlotgNwTaz2Ky2Hs6788XHEfvzB0+Yg97Mp5H
mMOtzfSJ0lpIyJMUEE+cysHVvEZ5EUuwLIjusySRAbUg8Jy9y/ZfCzMOb/QJdNFqu6eYKObtZerd
v4iTZq8pBbmY/ve9+Z2I8g/ZR4SK6pC7+xt0LRvxnvpMBcEVg6AxjqU8iyqsLxpr3ZqEV2U2crNj
AoAsL41SCBhBZ837i2W+iaAVoTpNOAfNEiAqW4cK7x4eOSKLqBvDj/IEU8vqc7NoYs96sH5bT/9j
XysMMq3KcomhyuviSFPyYqOUwncUxnKvJYUS7wnmiQEg5jvaKr6PhzZid85hYWRZ1m7Irymr3qUr
vbTV2AGgv/PBbvLJHUgxO0OZ3YbDYNFmDhTO/8T170c4t2rCnpZVN3TVLuOUT1+z2lpw81usMPoV
V6s4/YxgP5E2f0kfAjsKhhZF8JZLMv49xuaFtZFW8BUIKnIbwroifgbnevajGKUBwIJD/BAYg0aA
btl1Y91BblV0jiWodMVogRDWTca098Uik8lsoQV/TAyJot4bBSP75Fyk4jFNshP/sQLEPIQClxCY
u1JJax2ajufnoLDHpX4D+bLEsWY978klHiMirIXQCZYe1jrpMNAkNLcqADp4D+Rc4j7wWezmAtn6
KdZsrFg3k8FISzAa5/OpDqjqYjxVtcbkaOeFyCowkATPvbCibzOlPE08pXuqDQap45BtUmEMxZ1+
IOk5ZBtsIQZKRW8bTDrz9vBIxYTDDqJRrovQDkfmkScY7V2xiXaunO4d66GdEYdyIJ4nxmOJPdYv
LFh1cMrT4yiW14B4z/Io63LPUzfohtKsZlxgEvY7+avqzkiFVqsx0I3jzw3bAEjyo+qa+uAMEmXr
KiUO6aVikz1VyZ/3DRTB8Jqd8QAwFGhvaHVK8hW44DXTeDRx5uYIosDyrasDJyR4Ocm90xEc3C6o
czRil6zz3alTNgAwv8V0v5xGsf458bZRD0JHcMeKog1QmLbmZUASAQgRUOFC6RjdvflLNiCwVBvP
f5vHwCsc7nWQSPIcvJIcxxqNrCHn9cF89J09vAm1PN7osrSCDv9Kf35IioxZNUpcNukmKpUEAPb+
WLwtLhfcXfxART9IGpE/2KDElp6+IbOug0lOeFdI08cnZzOz7+DVx3awhYKplbf56xUrThovxo48
XkZHDp3wivEEo3QQzwZPay4TTmJIFx+ma4ezD1sYygmJbgvHHjm1PWoeCa5corzrmG7JYclgXXWy
5HQ/d4XM0bnuMDAJNBPO1h8iWhsWS7iEx0TzltLosiyA1pBaqFZiuleY2Gd1SMZRIXLBUj+sJSfe
o0xx0sjv2Y0Xdp3SHjRkfDAPgtpEOLjTexxGpRv3/x47WkzSIEbaVGIKX9felpCjJWUPgSJNFpw2
4Fp/Nb1Cx1cVa3tyTvvwdbAlzNBDtgRze/gdSy2ZhQYZqigKL1L3vPopWyWRxtUWRjvyrflteu5P
FMeuzTk9w4BadBb9KrLCzOVbdJawLCYFzugf1lpgQ08REbKzA/Wb23NLtet5/k9h/F6v1ZZnXtc2
9fYmiOiAXfcijmZb4LqayEgOt8BIRziFdIMAupxP6I1oqjItjsFz+UlJvICAt+HUj2pZh8nYiA0n
sRMpfHx8gmxnqw4rxCEMrZQCFDJPRzm8qyZ0ZsTjk4hFpbBHnAdzgIpriynTt1X/aEWRbL2+E8mR
8AdrRDLHzIhTjkdtcfHIa5RK+006UcbMiNtzTTgz2/I6FSYOK3wgOBLDT4mRmYGO5ra6Hg02Nhz5
NJWbGjY+IKFg0Ho5CLX4alKF6WL3RbZnEjcVaMtBp1NLBSstrgL6ney9vdSm/1nJO+On46wHoa6H
q3qQQc8tZpBXLaMyRN5M9PkFK2DjYUTzIuHyMACx3q9v14lnnFAtAmEKaKjBFXdwoOOwbspX8eba
jCEm8FDhUG8lhD/JpT3JiDVqUF3qGBvhtbALhSIvbp1lGsYjpz1rqW6PFgQ+NiZ7c67Hufl4ZAd7
P7kngib86SSmv4yOEe51u56kLZP6pdXNfFKrCfkkBnSCy/rwbBKxPoN07PL/ZuYbdi+apaYB7gT1
+Yzl+B6CIvr6B3IvXincHnTOyvxxT+M2o9CuieRNazaSrUY/+jeMr/KQnDddxohWigh29BsDkK5r
8CHWkbqIv0jkubnbJcwF2VmV2ATqPXW5LklE6iKOxOm3g980AernYS+gaoegcnF6e4ll9kBckTiH
UgJpUWS3UfGAkcowDurYDYLwURu3WvcOLYSTWUouTVtUj992bflMe6Toe2f7JMtb47DLsYfRWYJu
6pK9G1CqPR+2GfElrfdJwI5fME0ftU/3Nk4PxdTp1y7ZYfZyykhkYhfr1eZj24lD/j9+8Ve5cntn
nZtZamCEbTC/Eb8J+Y6wK/ZEx5km4yZc069+Lv2M95YzwzyYq5JD7Napk9buKzhFZyEzBqm0Ne9Y
9mzMKM/QxhXSVryXacE9e2v8neRFbCs6SdoBWe+ozOrWV1e1X5hCKdaNjNgDlAuCHBIwgHx+23yQ
OmeFTdB6ZqlT0yS+ieUM46BQwO7cBBqfrRxWuNYdsR3q8iRPdB3nYw9aXdjyUV81zbbRPaKZXkrk
RYp9yhQn1IF8i3sXmzZ/qMCPtnczpKencEYbBebjHR1FCyjqGg6rID85Q8QZFrXIjZuMhzGAsCMv
dTpRZ12oW7L/3B37kHUxlsOS9ERSoqsXXxMsIp3ekIaDfkEdsFb36O1VokCczQCGSl2EIbtAX1p+
HeWtMnvY0HmDJo3ZNxRw0VLVWldJWm0Bu/pjiG2nJLGycFxpn0WTui0NyszDtpjFMSijAKlD7Pfz
70d3c7wEnikv9E+BdWZP5YtyEOjqUmpWn7qXVSZCpZyisH48iCi3RC22Vyu6XJ6wtuw+eEBIBiv2
3JeQXYyoPrqC3yRe1LgXSlFztujyWsN11k+0i4jtBfrfQbO+RbiaTy9qyFz0zaL0RZmH9IktJDgM
55hb0yY+pODclUIfe8js5OO3re5t/+4PhIuhMrZhoZNlBQKGT2odAOuy0SJuGc6qOqudVRLlrq6F
+Af8NdoNJ3PngsH7dyLkPEsWwocBEUOUFKPihTRoynU7pyT/TTH04ma/Clhflgr5027MhwNaJH8y
IEBlBg+dhhGZknhbMbXRD38eMD3mFmR0W+u79bg9+o3IuB42gW49zUFw0sVJ8HiBqhTUzYz3zkth
NebYb5I7S/NAd82DM1dw7JlQHxmExMwE66wSd+4k4Q1AoMmovmOsQ/fRG0bLDN/ThaXSKaIjBEDS
vw+O7Cn/6mfZj+WDXAKGCGQMNr3exXSYNaorTfQ5P/gDfkxbSRBokbAFDy8EiwbetqDLhpwnIaZ4
K4yPDGF08jqx1Z0tYHF4SMyXW6+jpodBVpncgXaCdubB4McmNam7SeEi04HfrLmpAydbtFuIUbQ0
b033eZrOHCHkzMFCvWtJMRJfciq0gOPoWv0QZynMlRJ5zkP/SEwAld9KBDW1ZLxP1lx9QnHO8O7y
r6gTDqrC03qrP/9pUPs3JgNHK1iCZchMOjOuc0Y296sHyDyezLg95d0rTXx3B8jqWezsM32iq1ca
QD74WKL9mF+sP7ftJvxxaJgDsIpDIeBcye8eko0dQwVMvNvE4s3tcHlApW7H0TwGgEM9LuBxli9R
err1hQE2CIZRfr7LjbGc2WBI1iwziPrVFoXYMvlIFeHWO3D99VeQleKIMj8ByxiHvmlXwvQ621f7
qZH8vY1NuDxI+n1NkPziwdoQYfBxaqZBWBWzksfRQvTmJFveV8MPCiVyQw1u7J+WhwoP/UyDq/wO
XRGemAh7pweq11ik9Emd3ji9yGhXPL2i+gmGOIqumeKkyUs1L9PcujLw+kGMJ7qXMSxvaC1X5+h5
7nB+62Ivf6beN6ZeKDbuslVeQee22GHiJJV5b7FVjCDuo37ABEihVhZgHNLGqDVEq2u3tdAxLJbl
95MmBM4orGI2dzg0zo6g5wD3LeOWTNq0Jk9a5vXfB6lx6xfe5ns1/yMqHaz/e9zcEh6ZVG0iz63w
tpzgo6t9CmP+eHm6c3acVVWBgg8TN/hMwRiAQNPm+OARbzf5D+CadqsTc1hqx9SAFZOuLgF6Lu43
J4iDnI7KxBucmXxqbq7CGssH+ofIcIh04qylZBSiU5pTmR82KrJ64GHp/gHbK3q3v59bcS2kBovx
d51Ejiwvx3I8Rrpi+AJRVHH6Zr1JwE7jvoXzGLyPfZz1ZgqAobW8+lHLJkd4yMrxJFO/yyDzgYfI
kcu3WwUX3sowjPw+KMBFDVZs0KuNoKEtNfED8wlHh4//FOzn5chgAgQWIfgfpy/noAiFv9VWuRJS
BK15TxhvTOPCEXDpjd0lf4ne8AkE6AAOMZtb5+E3oeh2FcsOjRUzKrGC6FxMyQeqfMAY25Jsh138
rqMIDULH+WONX0EeDiUkhIJLYdQVm9hmG8vtpbyki9aSrW+gr7So/ELO9S597vTtbsl+PX+6iGhg
epuyC8NNePu0aPFU+qRDuEHVJwFNPDDdpzTw1xyDfMh/tOIt5fRo++127bDGoRCx5RKDMahuzLQg
uAk6mRaihwAFk0ODuE2yXtd50d/R4KKoe5yJwHKiV+5+G72ATkVvNpRzEOiMTyogEqRKRYHH57aN
8z2JsxNwwZY0R5fvrCWjlxAY9LIWGV2W9KouW/3PV5tMQqKYx5djkhovbgSWsU+vtvM17eQ/j86I
lYpK7Dd5bYxmKD/jSl99FRT40lcb+iHUd9g2NtTwvC5rhRkFGndEwQH9be+WIP9kgrfY87FFbp4X
7gJVeRAhpzC9o2TrUvc1rvX9kL0UJJkF87JdCXoOiW6RXWW0cMpxpriJagNEl6HhjZqRGz10kdaE
Qpm1i/bLzAEBBFUjcPV0q8sEWczB3wltlImCDfFwGeJA1fmfeuveODC3siNuqKJ3BD6rrwFrG07R
nxQlJWZiGosJzD2P7ascgpEXPL5sNL49GpyLQQuDcl/FwYyobrCp8f0PNaE6AO3BjiHOHTJdV1yD
0eEwwVjb+EPawzz6gciem71hFyZeVxCPGsHcX3Z/L1xsq6rPEkd5mkGJm8MKDifbpNax1FRBHeql
/o9J2WT0PTmOFYifHDAnToaBBpUwYgW5c2NIAaKQA4bjlA1sXapqXi6ch07APeWTmik2tnuc9RIN
PJCzy3kK9WJo02O5Bz0g6NvSoWS8RpRYSgC13AfDxqElPElDWaf/nmE7PVI3rSb5mPCzYXLuuW6h
B3Y9dkj2jtb8qAech27r5YUWSCEkkbdw36IGDW8pBj17TXU4FXLuVb1QlsmYjfSvEMr3k5u+78cd
0WCEFl96BmN80NSzjvj5396g5MJwctm5fBFPiOPdCUAMX3XMtTlRszizU7MKiVWlJ72dznkPclhf
ui78rRtgdvJNagdO06Yx36fgYfX1Kuc4nIMye3ckn+0pr4oRIwO7okAyqrqjNARX29O1Y3mQF+7k
aOpFNGf/cHSBQ30j9kL8JzjHg3xGag3hYpVrkyU8W0WouuSpMtjyQ2WCmgf5T8ikKYhqum9Msf9P
WWnOBD1izHgyonux+rG96ZKr7P6Dt8pctTizvnd79J1yQi0HtX+mggd2rkjI/mYJuQanV89oB7wM
mRnHFVO31VtCGrvKvaBoFkqEyS4Iiio9Nb/BBxP7Ymflzx3x6m7FdKGlWVBV4vMyybZiSfSBEv7y
Zjxd5/U5vstZFZaIugtEcomYGoMlwDbm16T8F5SHVe+z57UYLXL5zZY4zo7iKUtbfxVoOhCxKYra
PfOHSNEOwF9ikgKMAaHu+1t3igg6+l0NhGdlPWYBJloyiETK5xLI7PZGSX/sIcnxGh8uRN1f4MrY
sOn0BJU826lJHmg5c4ZsXExF1bz77/hRge6CZ3sok4Vzad7cJAjaQJNCTGtYQ6x/k5OESPOV3s0G
NTG9aGi48dTwH0w44Z/KiLMK6zUTOomGuR96LgC0jzUXK/SRT92rbmqVXCUW9pdwGBtdxMGWUPW9
viDxCj8gSUeS1p2VdIC6HyDy2HmU6PEqdo6D22mREI3Dzr+1NvIJVpChcy7ZkZnqeylRRBxfCZvl
RmLZsDFUoesJzdf8ardYBktsu/b6im6n5KtiReHqdjT8MNiW0MD5f3k2MMNcOIvgTxi61GnAzP8g
VYlR+J9zFu3Lw6rPmVrJ70sykitH8wMCL1xczCQ9fGirExvoWFSGuHmFHYflZZ4s2V3qEU96rcaR
+0zdWKlBst/bZSnN+9ZP+e9/r6BI+4j8MwSZLizIgdqSyyCQNoJtDeSa2fELYNvbiMqyPhQd4B8w
5+C+/N46LQ8U+tRdAYCVwz8GvcY+J/Ani6+7Fx9nmTIDZFlElrKJSxDc/EP5QCcnLYRLyyssyd7u
372emMXeFGStJfrC146Z802ZBDu+wVErls0c7tWDGkAGvgezyALgsY8HMoBpYKZ92eChwCv85Mrd
zmnovNMRk9yeTWDJTHUz2wqvI2j4ka/+xilIeEhBIXCnowYFDZy3fjqIeuaMbWHEA8P99Z59gcS2
nDBNmEypT6dR+HDxqvzBKFqH5WkDEcXQF9hxoc0+Gb2nofxMwpY0vHzMPLISpjKpGPXRxz3OAN2f
tbjTnoNAwXD7yksNlHzlfNfUSac3BbMUoaUVXjXR2sbURbR2t73Zgqmm8J/wWrrWOk83kEJa0Qoh
ci4yvqcfg8b9nvO7bAqURGNNEOVhf0rj8y7/yq6Whm0cwKDI+L6HXoPQkR0dugZcJjlnImGcPIPW
hWoo6S+QaoJu6cTeKoMF/zt7dDgENlQ5RzVhn/HDy/uZByq7jxwLfpc3nWGJ0ENxx+flQ3FsuzGx
R+TKgpVBLER6FB0JeWZdrB2YAJYc4s2WpU1W6mVw2OGpFz/Je1pl5GDriT/L8cYm+kjx5t4LS4ue
Be5OWKgD+iyCGtCX9Dq3RRkosvbSQWP52AR9G88F5HXMCOzeFtJ22WgoarrZKMfjqrCdDFFRPMlw
6bJZJow37o8JLmsqOWiQCoFtM/sacWDWN3GTTpyMchWBgFTNA6kEJUYuaLXA/6VEXJkVt1SS42Av
gb7RIkJc/JCf9+paNjVzGJlP39AuxnogQXJw0MX4er1yuCNx7JS//XLxD6AJdDkCxh942tpHs0K4
5bOGOzdu1HiJ0xh9qZE7ObrdbpuUGnQUtsEMchLgMqyqed0eef13QU1m8KTAfVes9fZ/CFu3Ssxu
/jwALzFgrjXbKWcNmSEPDtO4V/06sg/EJaONOVzI0fOAwcMG5lO40slhCsXojoZPYhmuI47tdwrz
+kOqHy92ogKaN5AJ3eO4jtOLjD8EYLOvMSvBng6lOcD5iHDY6+p07Dtet/L4rf6JsXxXpqvPeRFI
KQSRyoLb9wnSuc9StZsKUi+vWLmC/SHVzs9QLjjr8pPmt/Jnr8gN2zqNu09Zl+U7DPogoi5Ry9po
g/qHzZ88d2daEQ==
`protect end_protected

