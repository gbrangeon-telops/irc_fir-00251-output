

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
To/0Y2C4coh8VFh6WzI2wbA/wXer17nunFaUIFXEvO3kBprRAlXyefibFdeqGdMCN/jPnm1lnQge
X/HG5CdHuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nnkNk6e3rHUR8DaNj0C7aWkCs5LBgvWhHhtsF0DtIcgM1egO9JMHLS9VXFoTsIgw40ekMylMZAif
7Mz04TLeS83J8LIkLQIVFCxUoXkTdVbP2vwAOIuzbV0fNimpIIdRDB4Qyrb5oJF0cClV9EVhM+PP
xrslkcRoMPftZWbNXzc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fa9acIf/jWyoTf/ZQQ2RdBUZgeC1x0Ej+f6KiTiJLxfGAO1lB8jxkDwdqife8FqrZb9GuA0CC+35
3eXgFQAQNKjhv24q1nYDvGkg1xQe+JaS1IiyitufBE9Oqujx03ehRV4B4wJ5uK9qxFjJm3WBZQeA
cWZiPDwrU8E27DqZYUHGXiufRSfFhYToep6g7NhnZGCmAfAD7Cg9pLa/AvxaXAS9nnGeBo/RPlyk
G/XXEB6YF86+MUOkeRMAxi86Vcag14njI42hNh7J8Lfa4beMq2Avi5tz5eGJq8y6uRjal6wz33O+
m0Nk9SOLFKAmJ/ib8Fpq77uCjrQp1T7Cl70Ebg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h4sQ6/cKFAjr6toNt8WCtcnxvbT2RbQqvunqru/ZMP069wFljAWXbbabme1u0tsoVT7hQ/OZYU4t
+qXe0sbPKDx8M0x1MxaKDasoQ543qKQAHxR7Bn28bTi4sQCu/+YxH72mTMVFjRAGH6M6e+MhTnGO
FYX19oeiewDQZSakDrY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
C8DUdaX7Hd0diH5RVXOZCPD1GItaWr9F/mVcGAwJsPm7j/BsnnF1JwcYxytFDkPy0E+fcaWYKz9u
7/hZwJ449yH3vkp0VWbVjDe3BqRjhnTwAc32kEGR+a+f8HB/6hGM+mJkcuw5DhoveoZqvYIICYqz
iQAjheEs1g2k4DBWxSdaCPNW8fXVd3J/pZQSuvaNRnCtPGOVMt3rO5k/WAzjiaWwDL0KdanM3fU6
uD93ZtkLZCLilGdf0EAax4p+pGVd1C8GYV4+XW66vJmZoT9LNfQ7rG/mL7dKp2aZ5DJPqw3W/O9c
HVwQSloSjbmiN1Fhr9Mdj7iCZycwuy9BYtMK3g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24720)
`protect data_block
kzhemROg2wfutZ9pBt4pPLOGPTo4qIUWER99009/DBYmGMn+bzI5YGvv296s2sE9hn6c+0yMfF7B
0NbdP/oA2tJUyO8YRCyFDypTznJxCTLMaaUM7U/VbBhtkrDg9lbls6oh4noMkD+/Ey88GXcDP9Uv
Y5dk6nKFvmTR6GEWSnQAPLyrfhZIWFCZcSoYwAoDHc8OVum3uPbiPnvpj0+9jiSjNthpqYQIipsy
1ywXfweNHfCDPOt7daYl86v2Nagd3HwdIYR9FJHf3iMgEQnB6z/Ixty9XpRbP/DTVrGBuZxG0ubU
5/mwH1YaQBp7lB98XZvSXipajMW3Q8k678kIkL1qDc91h/AS5UAqP4QMKxhsOtBpuS/6VhzJmYEy
8qhLig/RIllMJYKbWkQ4hlweNTkMZL/VUXlHZj3xGJDF8N0wozKb8fECPiVxoW1mG6BLam6d6/Mr
SMrnXuu/v5Yn10RvyKP8iMJpTh7z3NeIpi1NqPNO5nkEI+cTmFiOy38QDsysANaZsVTMgJtj6qr/
AujLyAhrurvttWGiUxn7TrKVLcaYYVbJThbrrSU2OYvEE5rFtDwgGLvb71woPjbncDN8LOJMDuup
ZaoRTwZRtIIEx1rlxjqzGOdqBYcyeC57ch0t6lYVXQRqKlX7rz9IWHJDDJeF5Yho6QmX7/jAL+oV
OjboW2cLInPYIHhuXIT0FVNQ4po0tSIrxIxZBex3qtvnbiw0hlKoZU0z643njFJ/tmxG/XZo4syy
wnPIXMCYo1nCex60vMkPh0YhAM4oWps9Qll5VnzwmYN/taq6A5KQtIQRQAGdVIzvZLa2i6Si54hm
IbM57ozTLL1PVFk1BxZKx1a0+4+6ImRwOtlteeYCjKIviKU4xc2QHFTPitnYFz5tuW/SdGSBFqCR
1r3lZyoQ/5eGIugHWM/i3ZpzA7LhliKq4UoBXFUdYd7wgnQ8vzkX5xoZY/IRjnmz0H3uU/HX+WW6
xDJTNRlE8+1GsfFjgETvZqrd564Q6X72ePx2/M/c/GuPOgNTknamkVJet+DYdEnq8qmnKcS0PB70
kKAx/zRW1OqgVv/ruTA5WN4O+Tr/2s4PmORJTP5Q4mE76Cz4CaITfDbzg+WbaJNN/ZqGlP+Ts4kY
IQrg79cThBItAxltKxXjS3vZcfcktnNgUzLDOUclSmGrn/MNpiNyZ0I0pc6EfylqdED6hOveE2D9
9ra3meLiKZ57WG5Bx+/J88WZnr4dYqnp7hAM/sgDwfGNv5oN/mlvQxEfbyD7ubLjZZcqXr88geKL
KMUlKtzaZMVrUiRspaExcDtesxDeLwGB4eh27Vw1wZVydQDdvOyyOnp1PmZGa+8BIB7cGt2JuRfJ
2oSh8TZfGqGh1ytIHY5m8GuX7yu4++fP4Fepoo2tt22M8An5zhaVHQJsfyVCZzVbBHHF6m8gbVap
rBeYS5rosTZcEzjEPoQ8iWhQwbDP2VORi6WWLjfUEsKB6qKTBDzc2fBR5YgMvOYY3mRV7YUo0fM1
ZIZcY9NCROiZgjS17u0Ylvy/LpHMKYP5ILvSTQkYVWZUiP4gK0JbHtqGRSi2xpz6veldq7z4GYqv
2P1PoGBAirWHBgfYuDP08TWNjpApcV6slgLYsoBA9McN0XEhkCDfgK2b3cQbIBIm7J2f3X7V9hg8
WnKEDvgNuekrZtTvRvxLzg9goLoLoMMAuetxyjQ2u+ANoeIiAjHjliZ1dSoW1u88VRvK7UiDcXHj
IPO2GzgGHwCdwolC/8Xe+rnfNziMYcPSw3QJsMrVo9QzLylRQaPG8EH10gb/+xgMrU211lhRf2fF
aniae7dqXq9yDs7iqsc9TOqbaGRXyQTnJu05kAZPG5GGmF0EG+6Rqo6E5whbEihePer8lEDBhSuz
iDZQFisB+BCYbQoxMr96GN36O2X37OeKSJGt+jTI8v+d6vsuM6qD/qV2Vqwogq0FTZrsxvVU5P07
JJ6uuAemfqxexlA1Z+tnBjr/5zbMHAOC7/c0FBcldNeyxlIfD0V2vjsfaw80w+G1Jp9dZaY81k+R
IbxXuUmBUf0WQEDytMBfM/RzWJ8CuTEaSBH+Dif7GQMC6+XN9m5FYlA7lKDvd0KFeMPSvbo2IJ3a
EuVTzFCsFOK648yQGjLwNApuxciJyPO6ffNBVJonbn5Mc5tjlVQzk1CA4vI0LMdIwktCDimQ99Oq
zt55ZMLxJilNyt1atVfjcN6/aY0Tp/9kVEyMVLxSswt51hdM48elE9yE5fVu2cb325qeVDi69XDx
advxv4jxpPjAp25SmVLjoSUT37YtZdGSS7KMDLezPQ22KQ5cQl9pFuHYgU8IIy07ccM2tTNZ0+k0
shLPFErX1d6gQpA1viLpaROAA8iRFPY+idWF8t645ccedqeEO6nP3JY+ofYhtvdCVgdqHuyse8y6
z3xxkOUsud2CHC9lEZ41gdH8ebbvc2xgbJwy6ijziuB5SziL01RhkwNH3CYLOtx4ypugv8vXca3W
RA64jeGleZb5OPE8/4/onamchpYlpZubiZ7v5Qw3V18SF5YoNIXCaHK+2mT12YaMufncwwyYLoih
uXAMZCKM/rLnr9tEH0jKa96hy3aZrwslNc833ntsFX81lM9WlqLEhlWa7VI84rYRqKbcRMZetxjV
ek5X6ScvfXc7W1uXBQpRRioVkNbl+NQ3F2LeQ4zYSSCv7Elv9CGJCkdNaLIVcwsUcMfuVWsGl5fd
G0a3jTV5RzDecsN3VByUWjIh9eMzu4B1RUxBAs7ASfgXuZQWgovrVJVQWbcv/7Duh7AQjXMqn4/9
Ouj1zNMfiWeHt2yVqL11dn/m/taVF6KDNSoq11SApohq1TX+ZORVz5r5LSO7L+w1+3nEQcunN9Zg
Jl2hF5gCddavrybETN1okpM15UjpW26jlz4PhCtXONnsbKRn4OcUj0Z8D3iYJweclqWASlttDsfI
tMayN+3yA/QF29sKc8jREgRyitsEC7bPnAWNzk1A3vVZrebPiGDfpDm4DDt98mWMhhSblRSuafld
iR52PjRk9vIj3IwA9iyReyB867bXTWZhs3Q7z/9pxKd9sYtdsg4VGpNVjvek57XShb3ruOuLYOFu
PBPDR1fN9eiWuniwwuJUsxW0IP7CTWQAVIq4WSZzyQqYKrO1sk2YilKi4ydbmSBkQcaAihfatXt5
6RiD5eE6r0ELUpfaEka2Be519u+QrjtoY/m3c7vYfKSbIk7nwFDjWdqaaouFA82s9RZoYjU6dgde
qKbB/wc1p0zzzlm68YFycr/PM/oiyR5nGPNhGRfYuetHuK7oXYgp/kPsmK8XML/8wj6LVffOuzXN
ZJ56RtLaVcFmQpLX74AIFcp9/iIhk552T9jAGQ5unEFVCnmI7r1OiSXXmIqv59q8BX6CgYSrFWCC
eZB0ykS2Xq1/V+NuesSZUPf9umwOvpjOanZOTmOiKJysR12PsGlNpY959pkU0vGeNhiXN6f0sDkA
/bVSPIzgqphy4dF5B1LF3zvSzuNYEcQ7KdEz5IurSIpo7sRef8msSqMbsRr+uf9koS+ymKeqDjHf
cz/X01YeFRasIvUFG5BGHO0yM9Ms+dF8tMUQ+hH4g3s95mE43Ui+Bj+alp2nrWO9UdMHKl+2ZmlB
V11RIEL0q9h/O3W1gdFMEvJPgyBCA1S2laUe9k6RwXdPbuNDc+AGWC8FvRbp8/iSP1RUYFZZsqkg
awXB4Y1ckhSPWpSPawkUaOoCho/X/BJJWiXu3GrZLE45Tqgg/O80ZK7YEyEmAnINR1gx/Pl9XssN
IphF9h9oj36JmEnzfOT7Pq9G4L8COQ2nPRw62M1Nt+HTD03Nwx7IpLeQFUhWZ08VqzjpKA6e7QJb
+VjJyLHG1AxfdXuGm49IFpQkrVW74nzaIvZrRgBliMdg8Vik+jOq23DJvy9uRR7QCpTbT4WVQ7GZ
FKvvniUvErPLRoJZWNPe2GrEA66OXSW9P9b7Jj5ptRBcgLCiXkmKBNs2Ym63ezS47yAdJjwzN3I/
zKYdg9UPX1FhgaEOYg5Bkt4bV9g7VjeZirT7xDgq1SMQ7wb7TXzfzli5clzE+pvcoG//e7mPRAwS
xvrZkDcLsjJHCOH5Hr031r+PjK61F/jYQyyGIzeexXQCEY7d1Dg25N6lp5UOcTrTrF3DbXx/+XZb
yCwjBSXTG/0d72YUxYSVvb+x0VrAt+14SL8CT8BvYXIJBJe+nAVjXe5aLcOMKy416p56D+SaIEJp
tW//Q4Xbry+Ki6oqZJPLiuo6qI5g9WoGfVZVb9E1wN2D+WWKC+19Uo+9ymc5sjvQN3/L30xf+wpl
Feq0oOvw4X/baO7XiFF9BNzJWylpmYUtCG8q3ewbKtzJY8E5BVVgBKoZ+WcwAVseQL+Vc6kNcska
VcnoEBNR028we0gBQbGsBAkjNg584ybgkclVCfD25o7OG29AOnmMH8Tua7A0YcN61qdToa9id34d
ugGRXAU04/yApOzcb0KQAUouNIRQvW9GTA8jcHTAhuhfzq8ja10vzfFmTwmq7vPLTHho1TMc+G5S
PSRG+LIegdAISkZoSo09ZjOOxA54xnzjvdv1gg6iXAitA9mM8ynrxigWr5HhbqvKHV/nqJ0KlsrC
EfShEbMVYkLPGCUm56BmxZuQTczJMWAKOZ4km5gdtuvUEzdqWP6ioJlWSfxXJiqr5mXM4zF5HNpG
Ed/z47a3cwNVWxmLs8pc9LpUp2Qm+am3ulgDH/79VRsbLy4l/4jvWuPFK3bn5zoyopwqgYlgif3A
IhrQkV1JXweZSWUqjMaDggW0dqjnUcsi0G32qEuCBCQsUjxmPi1/BapZ8j7gCl71mvAS3IEn4CL6
apOAVQzj/HLVFO6hD1syc8dDGgvfuTacZy2goKt/HFPe8/zX/eB7epiqU+v8/1NkeUw5xEZWjL5L
9/RSy3ac+4NryCSgBFVDDW/Rtxfxl6moNNhjd6kkj+bS/dkLZKSXIynE2qAWDdytOqkYVycEsXxY
d3VtM9wQCJjC/Ac6NAHsefYSxSCfHo3s3bLtY+goiCmBo83uSwFP3WDFz3TnY14avV9ZQ+R3uFH7
YkO+4Idt4BYCqvu9tdHtwSXGA3DXyvYNbDD0qS0nUbEspubuzf4Ddk6GUNVMDPOX2oVS3/6jajLY
FiKDPU1cp9R4wMVzwVvxiGhRFkSGr25yzONdIUESijkahhJCNC5NV59druvl9o/Y5xEHtbkTIbAj
jQUX9WLNjR82Z2TnRrKkC/eNMv+6SSxdYaD2IgBiGG/jd8ReWb+i8Dp2MNYgakuSAZPoM96vc6Yn
Pr96K+v4ZYTcX3JURoHHN3C7mCtIOxny9gQVzx8p2jSq8Zw2bfLmFP9f25yW8iBpPbyc8qMo3/hb
v7lGkvEHhJbNQqdFIlYHw70Q861PfTTItkZVg/2mrTo2PW2Lsb+KPhegv1fZOL3yf2i3ruZHUEMu
CciEa9BZqfFe9f0huBPHjwFUePOV0oxEh6D0ck8+DgcOcEkdvHZEmaSoJmzz8Dor80tyyDrLHZ/h
T2LFtacNPODP6mnzB585Sy5xSP9kW6WIR+vU8h0epzAgF4kriK7ySyRBnixd4Wbb4e12jZCxvqqY
OmYjuDlD/3Vsr4Pprng1TakQB0EXPxRKpwSiINg6bbSt7jtmoVay7a8UifPThuO1e4ggd/YI7D2j
6rog//UEGsI04rR2xURqeELsp6l7UZXaFT4+mAXnZNgE5DHUtz1C9s7Z9AtnVZ9mJ8gfEob6y6ns
5w7Ozpk1Sn3AerJh4cC33yvif7oXlQupcIQJ3mIu1F/2BAkHWa0PcPMDKn+Ol5mNfbZHg4KQNwTW
Ox+EtzPwdKu/faOsf/KGTqMQzKSDgMUZUJ6YTxP7Mc6VMzf/Fgw2SNfIsrYTLGHic03F/cbvAHr6
XHr3sZdb2eCJ78dxZQhPrCPq4V/36OMzNjC8ujyuSq//1Y3fmgMOMXB23huFQuMdrVw2APwVsQE5
sSPy4IcWK1zGGNnH5YtjtjlYFvYDKiCGNuh/AuohxvVRdEHA3Ef+DQ3uBmEj3IeyZuydXuQko9sK
XTxaKlZbcvLeLlmdpQ9mUzAStHQx2YLNfxawNsU6Kyn80wQshpZNJiQYTP6KdFSWE3AMOGS7PJz3
oHryE7GDXZkgzzY+4c2z3utHyTvNUommBis1ieHFziLKfEkGfwx5WfTJslyFCLzcOH+C8NIpPa5W
3oMMk+gEQLcN6bAEuB2vgz5YXwPGNc20/E5xnxy5i1sUUeplthqV4z6DQ7biWg8caS9gqpTC5ijg
wasFD1A+wxu/D0OKNj/6RKG8sTFkEpIZY6E0ZcXY28vkl/J/AsvQKfRGj49Er4m6Ti+Epu7NDlLJ
7Pi5PvlaJ8eovsVuaAiYogEOgx39k8/y09CcFFph7Xw9Q13eB40hDcyuRFB7sGZbUSm1YDv14tql
tCKoR9K1MmJ0rbBT4G+3h/ZC0aLTD2TKtUqXof8jUtgZcfYqfcAuwDzJfFq5zP1TOcyr3HkDiZ80
mtd6U/oJtxKTJ/C0qZueF0Y4jyjxbzVOzK9U3umgzO2Ql+LmpYmJ+mntayXQx8HuaPUnY2Ujgh+n
SduR5TZo3egBljM+D7//jkkpfpOJpTQq+Ll9qiiMtArpG4XFZF2K4ToGtD4wReuWQ6F2pxMTauN0
Ef0UpyeDVl9xtpejQDBRXgL6X7LEIc0JnBvJBgZeiVXpN2JSGE0yRqx3+Sbudtih/B2HUCtCqQ3k
DS2IY7KUYRGE0PAeiOvl59iIoWOZwXs0K2s/h3z+Zn05YOc4wcEZoXsizmtj4EZl/dUzW/I+nUvS
EUgXqP4zXUu5ldLst3hQkKd8B5aqq882wFYnhwmtJKfEprfATEnsaSyNNd5TPBysDw7UJV3XUJOq
S8K2xNoa3wECif0Rpkjoz93YTQNdv02wvHDCWBCx/fWpH/L9cMaekAfHSNblp5GtZ80dqqYq2Cde
/p/i2+89c622b32gjc4EmjuIyx12FAtj0ayJAa/Bhr5oD70e6Q7MaYFtl26iZdkKQPI1S5qoZJah
VytzsNlwh1YK1tgGl4TUJB3pBUQWk+o15JkS9WdfY1q0eSSZPczSTuIYOwlfiAAiTuFFI0OKct/Z
o0m00OLhKsG+6XNxJ7rNvvlRq7dP5YVMG1R71IZ7CTDARJYyuPFcWkPdOAELBnmjk5hOU1U0ZxC8
VKeYUMrhqM95wQVlyAUdSRmllmvxWt1rOQRXC/l3J5LbwNBaNxTFDfNK2Oax3iCp64c0PJVeE6m3
aJ5A/Cc/iCyF1jJtBYzYYJlUGOmxNe8V//P5x3XxaReuW8NJ5kmBf1IgVuqdsgvmyE13rE+Wx/mJ
XREXcJV7mfXE67MxOgnimtfjvHvoJCtz1FY7/L1oYY6DgvIig5gGO3MeWbqbocOQEI87MIGJjYwv
KjnF9ds5RE6cMCKdnmXrFOGEy/WrlLvXo9CKIuGPVDfbV6xqiLqtD/BiElxe8giRgrDou5JWaY76
uRd9GPBB5ML2DOs1Cy1Lxr+q5B2OfySvGkdThBeLSfWBOHLxexuE581b94sPP2GKmQGok5Gghu07
83qPXYOf8Qz+/ept7DjAzObJmcInu+4KWfiwP3ZjuFNei04FKu42HbvyS4zFiLr6IBF4mc/ApZyG
h18vXQYgv3JYwy3RqPChLm3RmGsFoxmBVaTmSemIOUud+CoUySIZjEwLT2mYZu++ouUEAr8OJNyN
pdSXNk3O2DeUK1EBvaZMZsL0b+g2HRUiZt+mfDKjI3G1Ox4OQwmY1c8lDsLILHZL5mYsvixna2wF
wXqWQqMC3T8BQWaIpWgJHVXc/0nN+r+wpWnpqlfqoy9Axsii6woeDP3SVQqbLa3oMVDEgtYBqAmV
T669sSzihvWiQUx2O42fdUGKOZAWpFKHEkO16FSnwGITlT8jPCe9bieE89b+JnDeRJNgPrsVASxI
mM+c4cZSKytqwQDjIiNfCqRw8U2wVM4f9aZ3O212wzgjx/bQRkSC2QD40iqv/ObX9HgV0Wqn9SGf
uef2LnVbR0W6wVJZ4nwzL7Gx3+esX0UbQO9RNfFObG6DcYh31VpGxZgSLNKKcpo4Wubi7mys95N4
cWEdQWCXrkEj2aYzhhzyLTyIJ0jBJ/uD2OzxadaIEcBlQwSwPds1cyXXHCXRfXEw1oa9pEVfpQoj
9AFiZ0xZH3QKQ2SS8iOPL3JsgrcIV13+CCYIg0Ru0GHDzS0FFhePYJ8LMyeGr0ynaye3vw5Lk8on
QuZ91afwgboJCpCXH/0LRHPLgy7VYsAZXRkKENZoHvTJZvQzowjCp/WMBvisabhlnZDrSICu14I3
rEZ/bTAVQ0GuWVP6fw6t1DYWm0VNtpNt1UQIjeZ4rH7KcssSwgAtMvkpT4mDxDxnef/sAMSDh2Xp
9tNbVzlToVJm6DQMLhLzpT6NflAGD12+aA1oeVuWJ+4ydXRIE9BLuNzlniIHtP7fbcvPfkw+QJnK
No7qGR3aoy5ynUPFbcOKL9pcoe5bXSyRBHMnAeKWJw+UIKOSnBfT20zoTTSkW9EgBDS5zJ75uyqf
LOCyo77zLJrxGObO6oDCPWivasICJEKoFlVj/5IwxGKp30B4mEjyu3+i7qeSHeUCuL5EHJf4A4Wh
4H2LSxvhXOUEwhT3O/36sZXHFCv1RORoHxm2HF1LrP3UcOvj0P1u9adjlMAF0W5ko97S902yDrrZ
hQjIVl4QCAzl/FtZRWhfczZ4xRrXvJVuc8+2IK6VZklDHTKWc0asBT6W5CXcZOZwOMOXY+n9/1Gb
N7EqHbyJAArv1TiuTZMcxL6vdLHycRE8egKOCLVlk+MjKke+Xyk1wlq8YQun4xaVMJt3jAL4O1KB
91dJomERuqpKDfIF40eMQDE0Ce4USIyjwKxHB22+aG/WBUyXlf7GRNrbqGyaynSj+u7nmPG6hhu/
HGyee7a/4BHzqBrvn2vOdqT1zDgd25GOfuQXTPcBEIMeIpCUGjnGbrCEz4/dl7dJM+/NIVjrg9TW
Szwjx9xEtzb5iEB8e+UjMS7CHcMZUlFo5aXF3gAfi6xSFPATzHmyrSSRnx96izjBqbZAz3saZd3m
iw+gdW+KUNm4zchw/zecA2YnA+cDc0v5/64e2Ss7MPBTQ00Szy1VAqDdE3mgOka+EXRtK2pbB/o7
Q9zQkotymGhpFcDk3UkK8jNkodF0Rwy5AmwvmLuK7OK7TRd530/6KgA82N9eHWmCOjhcugK7p4aJ
cbjxemdlR6jj+UiKdiNreFos8EYbJ1ronxL72HpC6dha00GxqXhJpdSCGLfsf2BbhaBNgURBbb/u
aoALPsaxrR9anyniHws7RWb50oUJEr9wkNyWzosHwCh6P73Kne0fGP6IV8C+i7P+5dNYJohkJCNi
ZK1z47u3rdggxo+dbLu5jJucdMZj3MpqCCJi1A4JyL+Ryftsci4k2O+91aBoLS0vILG/nJbgI6pE
Cj9z+3bBi3LTeDdtVqblrfgE8Sc9Bt78B8QsmehFF9kQFEkKwlN2ZxWZcn7FqEOt84Wh16dva5nx
1ccspTPOJXJ+Say3dq1pidtTKFy3Vt2uSxdOMs9dIBBNOvAGVZsnHVN+7pLb9v0dvL89Fj7lDgYn
H8mJk0U8w0bHqwugnApyh5H5S7eHPKjXB6/WsvciKrXDHEhadk1X94K04eNayQNJyUd5gv8FUzPo
AXBz7BqHGtr0kGDXNkwAd+56mLFZSB1UG1de983Go8KLPILxhXiwEJNE+KjDb4G5VPU9UC2hR9b4
5ftg7fb3MtoXm7ZXYXSjUVeT3ujwsdsTn2wziQYLdGJXbQMhueiXXI+o9NA2ycnnDyy5yqrxhi9D
19iP2xXUmRHBmJygAXpxrHbXNm5X6E3a9C0GjKuok4bSFEX7fxM7lDfgGo5jv/OOFBhi2Q0aEW5c
0nio11R86cLd/maKjMFgQSJup4yGHjbLiUty8uHpFAo66znrJdFr8PVDGaaNkUvyIGaYWkw4NiGK
RUYwTzVPi4EVepTtq+cVF56IXkZjwj0gjKHFVDhXXZYCWV13UNqLraaOu8nhagUIvgC/UtqtZaMx
eZRusbfSLC1dShN045pieJkQqmfRh0g9E4hbmifOeilQh8jIf85yAECQP5SgRNWbh4Vg3f5M1+BJ
OUx4DmMFVqZsK+Pai7WJPQD+LO6g9HxDFJL3nETo574UVZ61uzJQZQ3w6YlKKEXwZnqnuHdsWCSS
rdIBRSMRq/phfcLipuYGLxaYziph4LiKubIlqOZh0OR+Tf1Utm2SkHiCPGbjOmyQlKFKzQwPkRBx
RQuybEVRZ06tR8quSbyD4/iApcivyPt4ZeTCz0oVaxkEERr5aXEMSEfYa6zWaWq4mSqcm75t92sA
Hjp7k7Y3XABKxVL8mGmWZfHgP2J1qkOjFD6gRhR06NR176zBbCfJ1pmvQC+chTBIFPpxDkdaKFGb
ECpq1lB016qi9MCyFiahpor4hYl7cA2jtOQILE58dYyoFZoQXYygXnbDsg9DePoI5lgmrsQ9G2mn
Le6WE3U018xO8WKgxOUDcP8JD1uTwVH1wUi6OB7ZY+7PUAFuCtZD7Q0uGDTN3CEF3UL6LQWgXVvU
jfSxYOyVXAy2lBqV78X6cOnSOE7Mj9CWTRZW6u9DLHBmViVaEx0JtE9aYquPEGF/abPYuOVGdGjf
NAgI3x6tI+BXWk0B3qSIoLSjM9WD+q9PJiZeRIVnvCt0SGhTVXxmMkihJ9ld512aYStMme94wGvR
srcqm24nJo7W/LbuxTS2sIQfOweGxf8BFdgykbnATHsTnwayhXXIJbQcPDhyIK46gSeO4Y0XatTT
GAmiTF6JcyBNi2BEcqEYqNqEALUG6oR+CEMnFbEeBjQIjzeir+yDYoE2pzJT/ypPyRslAZop2eNy
zg7KwQsZxApiuAzJL9TQG6602T+jW7gk0F/xd8U1B8Nimqu17QFlAtNvnp9FzukTCo/tWUEtFIw8
89PQh3GXNppCba+RF+E4AUId6Mp5ghm8VCaCn/li6UwBHMiV3Z/JYUH2Gvl2HyEeTMaEESHRbPNB
eAJq84AzJ2w5rycx0oHYCy6UqHCGB81yB/YtT+ZGX+BTduRD/mlQbeyNlkuzYXOEEqyCLUTv7QQ3
eLNaZf+5Httn02JM9fg7CoKYV159vfA4ofK17AOZ4GHdAk4ymdw2fm7zuzXB7agzNU2KNJdIJ8eS
hrcJsA+Hjrr3E8qy4Ec3XqZdLU/cB9a1tp8F8EBLBYJtqo4veVN/GaILhrbZy1CHE8/ince26mm8
nwWZj8FH64inGKnRDAyE/BVezzH+XS/zWTP+vHzAAcBDfj3RMi00RxyrlYyEt6RI5s5nkJMAqgRW
5H9MZHJk1Ld6WdI8+CDbT3kdPsvw8nW1JHZSV38DEVIc+AOBAOY9teqcc+QabRYleVfzcUIOPhOm
4J3m7Om8i6WVJn8nNIazQDP7Vs2oy5U1cKVP2IEhSjjvj8Zd5QoXxEEzqBvafKlaaOO6mQuwI111
L+hDe6ROVtEKlhl7tRpDRnF0M4EjZi9rC2BUKm0ltumlUzYTh2eEy6XvEDclcfwrZxyoE9uYu+k5
NTlPaQWFpflK3Imj36Y8k92PDLPoeHG6KOEvgScJlZrCYbHabrznuu6m/HkarjDBNh/qKhstb6Xn
a2SjdWSw2yp1KYmiGZv3Kno5tqMFmwT6bfTd7jXw+c+4Ei9joeOia0+U1otjQxX6++lfqLyzh704
BmtCIsnMFx3LE9XOWoz4uWIPvxKn+t2vM1/9mCO7Lc0c2XCEdxg5V4+d2mPrkBVuOtH8TUDm//fg
LtHOyPTG719IagqB/MPfm/cXd4sKGDJIHAmXsgJNupnI+L9Rr/tTRYw9oleqp+A027x4kfFOvByb
V/DAzTjkIsyY1pKiW4VayBi3j6u3c3rctIKwLmCBV95F83uxvwuWRkAgkqBi9ZjVB+5TUZN6WxxL
yAAHaWZPYLmqiwTYrvCVsexJLedQHXX6qm1mNAzlqjIUjgdQYwaovOIIV21HxHwkZ90SBOA2ssrr
lZxyD5RJK0qsiqJ5BUmaE85hldzCuDjsRGToLP4o1DclBd3vH/XQSSVH5NYHXplY+5rDp+i2tsEN
5XKK1EcLGOYDJJJjcZL2vwXo2p3kc+nInqR8peLPukuXMm+4YxM6PfrMu2y8cRf4bJIuATp09iXb
d4eOCaeHTcIbtxU79qaBF7eb5abgxOnxvCXCGYDrpEj42Y9rzMbd924F825atxXVNDYIoVYlxvHP
QM7jDeRyLJcR9na6EsVMMGTn8kRn36Fs75EL2GqL6wXU2gBHuhI+KyWbmQvESrBrZzFtkCl4H8/7
RahxCy9HflUxcUQiHfQ+W5boo5mpGA3f7Z5uQi1CLVETwN5lcSMAV6jxHtbcHSgxHjN63W4yG836
2n/JK/LxaYWPjp/9OuxFWo2UW5J1cOlms9kGvIghXdTQwTYfc5TMpjQWAUrwyQ/5xRtxCVyRgFQB
UiTahOPuYIPEt++613uGvhIa5MR48ywtpdFsQtR5OrMTGUNQEczkz/F4VmPCDVHzXPiiwzcTVgs2
qgq2ZabN3pVG0CwqsQXJB7QZM2g0fwGEGIPkg92zMkL4CJJw7wMlzmAJsjQBsknwvLLbP+BJe+jt
Uu34YHal291ViZkz/KVG/QkyD+NiE+tqK/eKA+MMH/qtBqyXdDFSErG9LygpJq7aqwucqKnjwi+J
S3HqWWcx5XqQySRY0Ef3G56RJsEa0CRPz7JTdQn6Hr1PCJnkJfYoT7vZ0B6xEQk3itoL1b7xq3wV
j2Uyeyd/t0UD331iWNnT3A+EUXW2jSXIhS/FrcsnAjsKe5b1FCbT8s1j+zn7WhoLU2mcQPwbyFW4
11PJBLHSQwE652A32hpUxsrx21gV8ogzaNN9+Xmg/nH9FoTSKvtTDG3cZJ9aJpRq0qC5sEEzOxan
RFwye/hhBjB2J1eTkKn84k3jhtz8UWNbRaKUHVXjuj5INIGvrORvSuUcfoXeUzxoj6JzHTD+Xwfo
jlM8yJ7+m1MWiQ1og0zWcMp1wDOx7n2gC+x8/itMOHLp4fR0WNh+5ZpyZ4e2T9fzhixi6B75oRQ3
9n8K2I3Y54ogoS/YhHb8noqy7u9F6Krg948VcBHF1D4z/KOXCfz0HOL7+esPDJMJwpwT2C2YnHZ/
SCD4nHYXm9HSuf3rRGvF9x0fyby5Yjd2HjB4w2jwj8MmWkb+bvtDZhGPKSisXIMBUEbqHHfpD8wJ
fnRbQMehHNCWGftdy8pEiW7S69MZjBCiHBmLVjw1Nsr/anPJWgcDz4i/0NB9QeFvhJv0oPdasQaz
jtsMfGgVuQcIc7K7S/MRhNTWVOtisRci/npcTPNlpL7U2iNjuyIo/XKVTMZ3eTg7v2pm6Ogsnm/O
krFpj+P7w4oyp/28E9yMnfiwFWpMkl75EM5u5exegshZrsBqjsNUDd2PzCL22k9em/bKioxIS9mz
xpSo9rw5CEMExdBcjrd7ylgaNYXx28ztYHD7n90C0dgLVw1fI/v48O7xZAgC6zliNDCW283/SGpo
811AepN3l5BKa7Tp57Hkv9n+zQCNvyuApAl4vY2JMIzyz4/AJpbbN/WUJV5FTdnekt+3ripWSNjZ
rcvYYz9Hkal5t8dTJlHU5RkYPeiez2JVDt9PzpVAXIkkbVw5AWtFcuukrL5QfniamvDFocKE7JIg
m4UkMlnZhRR6viRDIzvyAHLexPeLyPK7Fdu71/PUIt0z7uCV7tPeidN2gzTpqnhFuvj/DDQ00JX1
6xYt69GhqSFYg7qqCakFDVy7+1yLXh0xBBT4DyfggpynJbRHRsyeTZ4MawELDZoRFaZrfzdQK3AR
vETmXKMGktJP/9WS1T8T1wuKr4sNw1GuaOzWp8iBZ6jURzy6thBe+sE1Z5npvci78BQb3+nPHf+e
j7C3aBKFT/Ee0Tzi5lCtmg93AUBlXq1iYw9Dydyz1zWKW09R0iDJx455YWUiBWBPdQPQOvKrrz1V
bd6M3Q3slg0E9PmZTUU0KZaTJXlMoiDZxA2SZ/weGo9zEzai7oYwMu2Zmuukzupa5B5dA/L47KH6
7KmMYYtPJpJLjiTSPvr01px/VgHYielMebvjPoP0zozQQhP8fCYq5SY+LRq/g3KdeMuA0cJHAeUW
VwXCftX3aek7yYcdpTDJTalP3AHhZFc3zpJRXOuBf2M9dkBflatvn9WYnAviIAYi3JZ4PgW/uDtW
O0YmnTdZIIcrEI+CDXS1H4kNM7Ud4NF4DKKYbqUsJst1OnLssunnvoUXqEqiqhGOt6BoPaWxFF8C
yz4XhVD4DTZpfrZJGP60svpPkydp1zz2VGAUZTpFJfW4Uj8HganbuK7MiCtLFk/KfNZnixETfwVY
uSNeX2wOrqUGgzP11WmwmuknIJFcQYoKmBj1NytkcBI9nWGBu4vUgQyt9spUEvbo7O0XPCtRlHle
YtBZjhEb5PpbpJo2bYQrtyOweKVYuTo7XwfRpoiRGb/IJVnBDiDLX9url1kd5JI6wDoRcxRif+Jw
gGqD+ZzUQ/fVnBWC8wsYPjBLw/lNYsd+1hYmIIdx8XVX1Mw5vDuy/TSKdMLF6YYIH+lelfZ3Tbpe
J+HTmjHdufZA74dB/d4RMsfP0etcCu8MWtD+8xLs4/MxyymEusuLlqSwkW/5zja++FEXhKAFaCxD
+HcgaLiLyiDI2GTTBnKtWR2OqZIWL4265KEDomUAxlhT5WL+zetMH7ZB0Ef6d4/I1jISC7VaaKCv
03825dTs2h2V1CAo48K5eikh13P1B/0xdLNDmTiJWlgDaQpBY1Pb5Ni5j8xI3cB3j3k8NDayGv4z
Y7oCKmqIyCaJzGQJxrhKE0WQ7p9QE4wJWPVeLFMHCEOfyVBNrsfStJ/opDGND+vVJaiDqInDBus6
KANxXMe77kANu7zrYlpQuqc4uPnLKt3A3v7swulaIiPkMVXLr+7XEmlH7JG/PYvU3/UiYeAWxoP6
wz0xLAtLrOcfw/nuUCz6ZldwjIa7b98XartRe1FtB9x+NeZX5D/KJ3RNnRQZgusEHtCkJynB6K+M
1Qmy7iJ/2rHyf52rzQ+vooiCoPLgpUvtdFSPeje7TUrTTfH7Tcd2FHS7qZL7fX4T+b6BTwP+5Nd+
BJDWvZWD0rQbHXBc8PIY8vkQPYB8LeQuBj7EeI5ALbNfB6WADiAZa+B2LztaZsj+2r/STBxupeEY
uD1Hqd3MjLE/v1lDQVo4+qqKyh83IZX5JhptZh8HrVrnq1PjkW57H6/XOEFXGW1RRB2630PZKaWT
thDPEvH//qFKtDBfv7W+5DXauO6nePTaCYPm9UQrn/zrVBspRI9aPbhMnQXgVZNGRA5CAJumHHQe
UY3aFpNyYKcKAfgn31RI1fznMZxMKNwP/jCWjr9YBL9Vdb/4nhl2AE1BmFkQZDTlteWrd4+NKxtn
TiWyxOZLcojzC4EPmC+AfLD3cqZ4XjAtS+FOkK1mD0Ncvh06EgT31zhxC/8tlDBa5tSVrodvt2kM
HVlOvc7cdcKZXO7eC/uL5mfnTeZM2pcycU7Rw6ydjpEXO8Z4GLQE5SSez+Fwc1EmmJKOZ3IGKpcl
lxkqq8gYk/H8SO+BNUhtqNQ4MxLu2xqsjpYO81g9LnGud4SHGERzYhk6y+5NH5eVQEg1aoW4WnEy
Xkut2g+/JwJGQLFw9zMRFxkAXhbsaWdOUhZZ6gd0J9ZeaCVfAqbjwL4wZ+I4+T1Vv5G5bJj81WT+
yFo9ucxmW62R1hk15j2xKDQVzDkK0lQvLBuNnMTwzKY5mT5ON3hEzQ2LqCzNuFrjDXrxlHaJ8wLH
4xRfpJJ1DMCcCbj3ALIk6I9i5HZ8byDGNZXAU/CghvxRbu8gV+X72toL8kDRjYwe9uVh0qf+apE0
j4PgghmYL49NX81s99gQW0z3OtGFgqz8GYiCreCZgbEs+FGPmCLO24bgGNwxyj8OKyZOwnv0bL3M
wRAfXjwREx5o3IlZRMBZk0H9jTscTMIivFUgMw9SlkFnUqsfYZ+CuEBuPq/Jmux6rica2xQPOv1n
R413acOQjIdZSsWRENy+98yIQiue4AwrthlVqTUAXRnAaEe5tYG/OcFD4lEJziVRMRKX3cFbLVJ0
VPmKKh8q63q5p/94FHS2OpVKsxGjf5Fz0AkPxs0MaPfDtL2ue3isLQcSDd2v1Hrk2cJ3VOi/kypp
W+81BfFCGrOCLZXWqaPseSdoSdzXne6l8Yy0fhY/AHwoNI4iLA8m8q3iTU365eO9AexsbW699i6P
NxMGXpbvNg7EBF5Bw6JEZau9Ty9WokgwXBy0v0C7pXlN2Ic9CLEyNooW+Yq+rwn44t9mXJCXDAQC
fbEsuakoSbTlwSjZC6n2svzkTr5JtlIu2eNNXxLUlZQhada5QijjPmwvPun7FKvGR1ndh/QrfTLN
Ueie5b+6TgxDwwfxjNH0uVxbk7nSb4w9nbeeLUep4csikuwU7FY5w/5oVygRItdPD71MBZ8M7FeT
OGDuBr18bz9tJSbqkZVOR/ihAQInYTWGGyEA0CZR0LipNVEWF00dggu6cJJ/e4GZlsS4ZYG2nqSh
LkocKxfhxlwvvJuAbbNxS6YizJS2Hk0K8N0VQZO1/rhtte8v+Z2S3dk4A8646wwI+a/wtln88KTG
+lgw52GgFgLqc7xfjycO4aQJYzH1lKxvqV9y26+F1fo7hK+fHAvoNWTDA74A9Gcjebixl/qXStfE
AfBz0n4i3LFXzjO2nlMgm/heBmUpxJ/BXGFdt2NLiYJMU7M6VAJG7+tB/5EfHJinjn5yL1/V9mCX
NT8nhIxXkvbyqhByfwIjn/3tEN5LyVTdTLk7Nc09ysrRmpaE9kvgOYU9h8auhSP5U3BM9c13h2i6
kgW5fTaoAhY3dlsamqrOGT/Giq6o6I9P7RK52FIc/FSVAZ8IfbMlyZtRYsc3evgxUYR282RvLJwG
wxS00+DRFdZ3keN2UmAyzmciHIEW5/T7Lyj4ovWWtr/5WGjQw4RRG0QAGo9NSEYNuF9/8x3ZfcDd
BSo3u85TwYPIGNMsAj2ovWlh4DIVjSFVbTCpL0IyYuao/zOSgeD8CIZkh5TuwCbQNi3eOgP1+wbV
pUuN0WSvpvkwPiPC1wTWPdhMrLdfJg1CFIUb/ownNgA8lSRH8IE/cyroBIqEyZ/0AZFFBFYnCNGq
+7MQeNB3erO8rSz8ZRWVTnGh0/EVtwdG4NupAff33JmX0mgh3h6rtxs1xASxBgdjh5nj+MUAVgxS
P36k2HNeJJUoWau49gRBDdVNNDBJskCABf+LXUPXrfRerpv/Bs+guh+W5ctK0KHZLJATpFrbfGLP
TdRUiX0phUu/TVrFg+FXFjGHJ9P2P6yaHZwVQqs1zv3jEYjbzsR6rYR2vLx74RyzhdaqX8w/V5jV
7LCH/U+IdLP+W59h1mbW+EZ88AXpmGjPiMsDsOv3Xk818zu2jQzcBamKA58yRS+G/tDBpCWlS6DH
wHHW2+5FYx628mJDzr/OfwOvUie5AoKNj9mPblwSv3czaxJf971Av4dK4vAWeQ7vfnJc+DBcqSP2
YEERs6dpt5Dbhjm5SqdMVim/BWuJukHsy4UWhXeTnusrA2R2SRk8tB2TJVTJk03J9ruFz0vaR4bU
8taTAN9ToHIRxYu5jsy+YESKG8o3itrHl8wVBmj9WhI6BeJpZUUOiVKkgXqzAHr3FsyhwWvdnD5k
T3R2OFLTEfVboWqNwhuK6AkbW++Vtek48JNAnOVh8rT0b90grtlnc8TzS4umqaYpjiUjZw2GF6oQ
x76Wrf8tcLzlgEEIt4zwJyhqnQnuuo+RyTQGB8RWrEOQ7BCxcnPJdO1Ngwy6qFAASjisrBUDkmo1
vuOTEtR4BxkpgNzDaGrLPI+xRLxdomH1ttfRG6cu/0oQqix7iv4nnzVeSDb03IdEYm9coy8Jgn4c
pnGbdQqEmen5U1+CXtCmihsHKtTjyak0R99UOFVZiAoIwkxZROkFE9Vknt3XDqjVk5/RV5nUi0sJ
tpdOs1R4V+nE6hjOucoOdgodWmzXn/E0I6TovXej69Jcypv+BjHr5GdZp60ZXvttDFX4jP/FgUN7
X0g98y7X3eb5pteH9s+x4j/Z78OvMRntwkaGHKsWBJgWl/rwu5a7JHTTwXZwnC3F2OQxSUZX14FG
Zdqrnnipw7X6e438zOZyGNxkHG9PGzLNTHh1A3PFrplITGNUQKuv+GG7KIcFlcHMS8J/3SCJ5SmN
S1DfzIwms9NsCwNLK2wOBKOxdVIO2CD2pslzyhRFmwSZqo2uz9BNw7QaCVSkbYgsIzU87Dc2UPST
coSo2VcNbT6embk/7dArgZ71ybKsgI1kzDJMGlzWX3ubRRBKriAvLZ/coqhdkbRt8x9hT3fjOJ4e
LqPxqo57qs2ReAe0CrTgHm9hIMDBrhlYIm6qlr5zX91rmc+Xe21TGVHkYQYj8fkXNHLYgBcVSe+5
B0wYS9nnb8dpv76oXbZIsXCbELXBDIiHGz6GsRmjWFiBJXwaAJWZ4BA84uqxRcuMA2Mv6MPIjwN8
2acutz2x3q+gFtQ99ntxjTsdZtg5C8/73dvrQ0KwKRohpt9zb17GClcGLuN8PYuueikFjPdsol/P
mlCr4wdkeAKztjUcZsIlrs2zqE1OWIcNQT8MznlionPX4Zl7q5NFzz+5+Kjp4PO/8HcIBovn4RS8
5rMhuR3G3gYDjDThBVCEG2yby9nF+/CdVC45E9JogpivYZ0QFKKBUbyBl7Ur7Y41qM8J8+fdBX9U
L+I7FMi5J0LDXuZFS0P9wsH7Mv8NURrDUHiilsAV7K5OHWAViTdWyXLcWAD6A8RUkjQzYzuhhGpR
rzjihOFuMueMoxza0tb9FltA2Nah62oNoj0E8z+3CPj5zAhvqlrLwxPZFeNLb0gU44oeSKnEY56x
tKd478iJ7cSiL5Bc3tie7+4sEYUWA6KeVHt/Dc/JUU4eJrYSMi6L7/ZXD07SJtGOuh0aS7sBt4gf
V1fP+lWLZkZpKR2ijgqPx2jKa9okOCbWxCN74HPw2mPiY7pvgCOmqAGUC62XkQxpdD2tpkvfP3sM
MDJQQ2Z42O9M/aNN0eJkrMghWq2LGAvqekF6poh/NyZmLZpHCB6A9pQjE/9clogM6ganp5d/SzB6
JbxlqzfsgkTkiR4g9Yro5wt9+W48jPWWxm5k/yTpu4EMdhE63NaP4Q20fIrb3ezao+A4xOvNL6/r
IF/9K+EuOeVhLBDq+AqoU9SwewJv0H7uQKCkHmVfS0RtLPH2hPfZqSlmCA1QPVgzs3qvtPP+iRlK
Qdd8lmj2vrx0ko+0ld/1zcGHuzyHy4U8IqA5B65vGdkEaaBCgibPf7o00nEWUNR0F0QVss0nT4py
FKXmNoVrEUptnLLu/PvzwL22zNPAdt/MHYP4VKqBafRKkgfXwEtduoOZsaKG5W4gjo3inSmqH4Ko
vJxrEmHJRrsAthSP1FyJFHuFQr7S+5gAP/7PI5mO7xcWjZ/ospBBWWBUCuynWd11FVj9TzVKfi5g
BveXJU682qTQzn4gDHZBoIBgeaPDFDcwAXgGEx1PIxW4nGKRa0dICrAE2e/8fHYe1mGG1/U24ykS
fUu2rRpdz798tqMaSDVhbyGMEvWloK9J8dvE47PL78YQ5mOsUAVhRVFjmkHpRA/9k3UgqUaAtlLj
izNLpPAoIXqstgwKJbJTP4+WP6b51iCDO5wDssqU0+1yhZXIl61KyyQIUExAUm+f+BFxb2YfZODl
XFAOedMAwk4iVB0YWQsdoU/hKTt4CfTulB3vWpC22CkBe2m88dqbInEDCU8KxVo223eO07cvflFT
mESls6W4SeoCEXpqiUvbfqt+qVcIb0lDbE0PKz7WtlwcI64EP7eGD2fSyOHC9UJ8wVTMuY8wgdrS
DEPOqyBlDLnlxJRdHAWYrfiwxuFomNO5DU60dou0SgpF/McUXbQ7WbdXUDZQl7oXiAA0jgbHCzxv
EX9AqyL33mcQDtFbbILF3p/ZxXCIYWVGyASKIW2AAYiBhnBCY4hfB/EUAnD62YYh4afqtrL3qS+c
bucy1A/9EaNmdmBpODbtCy9w6D+i3bkNy6zc6FzeV+3x1N/mVt3pGkRf6o6h6M0NXl2g0NZAwVwW
G7AvTxh7RhsA4rGAvaLxsUjT/qQLXQ7OVw+1QTbK5mMuMWDvGvOdvugVWFh1fpV2ZsOn0nv7zjxL
Ea2cjtKZTzYVHSaT1ziIIwKBrxTSHbZ6toOVa6YWgyKdTgOsHMYxsPRnBdIgkxp6sAzF+8mnBVIG
UMpNCas0N9hv/oXVxzJZGiHkJB56wel7lcFHL8LQ1KRHFdFo1Vqo2HI/9hxmp//IQko4bdFAXWtc
y+/v3lggB8X10W6bgqsc2AgwXjwupRukEKUOL55dfVreeaHdtsNiocCqK4kcFiInhSxqfY5EOE9h
KoJSztY0tm9B/7Y4b6te3m48Z/xO3jKAEXZoQ5NFuNzAwhiwl3bxZ5gRIEhzV3wPLIdokB/Ghhkp
Tcg2Q24tSebCgMrZ3UnmrRmiS2MfoPWiZx0GZaxQ1K+zCTxLgD9VvjkYcLr5GINSplXKoiZO/M+F
0RsGMCQtJeuvdH47A/WxGk2poeWwvJzuwhep8DqtConEr2gQ62Szh2RbhR/Zh0iqXmuPVuUhMGOy
wsCHGoYPHdSkrTioVuevqiN5sfLkRA4IP6zy4CX+uhRd19JAOYSo4pJWwKVw209uZekqBT+6H1Iq
/FcgdhLcdqkS/WpB6Woat6gRy8tfskzifTEefrt1V6tY9gF4oBsNuyu6fwBtD9qEJvsfJ9mnhKYx
gtlTUKd20zTcteUE9z7dpnLa1OndsoNb0AYSb6gKLKJ23fphWZYpyVl5RbuB9Rs6MGv8sBJMoOAM
O/GCaEKq3upY/mLX0IJoDipGNYRJdJ1cPiay2GwtnslQ6ZzKWOePtJg7iLhMlGDJPBycRf5Dtmic
xlCOjx6ulmcCMZbZSjUDsdxtYbthz7sMMtHJVizDB+LoEVcTlaTmjAIz9Yz1d5lL0PfDKunrYUUY
XNYBMDxbmZooKItkZoN8ByZ5hLUahujkdQrLMQqcrMPgwQGXVquNRBBSqrfEQHYWtrGsiEL3WiS8
/JKMJkrsHOuugjY0mJ3mwrivL6cKYq7rWFpb7eHlB/M1gk8fw0+ya9WstXkdauIxcef9p1U885+8
yaXFd6dSXu3Y27OBJ8qXpIhlAFbNIHh/2/V6I2HOD5yqR8HDt2mTqCbcGgHZT3jvIAWYTfeEJSlK
PsHV77cDW+hov/I0zBzZtL1SmuIIPa0b9iUQXLNSuP+ejXYZdwn5KmVyT2CCXlzjZUWCVolo3kBe
+b3UKGJG92sPiyjDIcpnK1lyxkRvpNQXVp/rp2zgMojqazy2xfF58015vQOBWBDYa9rM52t6D/XQ
vSC9f+6t7aSzLfD4C4M4exbvzqCSFJXd481u2To7BnXCsF8/NKu7mKQ3/1bcY/uwU0f40eAlo0h3
xnoWxjiusOjlnunUhuDXYiq57Mxastmkjy9l8TyH9GXC2z7DLecR5P2TxfEpfN7E8G3GVVfB1CbG
bqu8ltIkuusCcx+a2EjANfXRiX7JDOVpxmoknYfrqDMwKFJ9aBvfdwUwGEBrpGziTsSwjGvbtbtt
jXfyUrsiAR4vC0ShzPVM5esBTyU/Cdqmte7zuATHboxNLYmzWNbiXcU9MSoinjkWC0v6ybmjh3E3
ZgDE3SAChbAZQmamkKa0uxfUsUqiU/R/BDwdoE2WvgzXQN0MDija9aTufDP0zi6AjgKDygw+UTYs
r6Wjk9ebqioSdkL3im3cxbesHw+Ii5DbZhE7fXiFXb4w1Qaujp8AJ4jcoHA/kLl5w7Wpsq0QvBjk
b76OcQxlGbHbxQ51fGjH5cQtkyQMbVHEPdANzTdDkBy2wByxnbYV1A6BMUVMSNzMzFDtyeM5EnBG
HrSY1WW9ivxTHfzlKij+ar97TGTAjpSVLVHNfwKl+/rpgI67oDtQXNAhfsduBQ/C52KKN2KwRYll
jT93KD1EcjUTdtUMpl1931yRqMCDUVyNE9H8Z9HMJXiyOzfbdP/nvCOxWIB28YoDgY6ZllsCFGvZ
PBYpehKkt/9sFa9l3cyOsOw7jWQDUc56OT43ut7wENlE/lNHC56SK0SAtauU2CQnDsFBeAdlPwe7
8uuYjakDWY/T6SZRg3csyYwZzfqXrAHl2joDnl6EGeYZqThBhLVoKhhmDcE74C4TIg7GJbMCVniZ
P0D5abeE+hyYQjqwWLPWyGfG9KsZ2pXYg5LwzLoAzJ7VROqb7uZu9iOBUdsxndvqn9HlsZXw6sbi
yPP0BUKpr9Is9hR9MCYkkZ+2okxGdy3BsWpYAyyoLIUtIAAegIwaUDaehdCdTtShCIFPZ8EAQX6V
v//ZI/gtMG5fr9SuB1kbJfKyuneqvUQCuGQU9vX/ySn707fOYvmfyv3ac2xlfk67xrZezWbDf+fh
SW5wziJhRxrNYLTqY3eIQXWkjgmWRwa4e6Z0JKuVBs4FAeeeTKd0TqeNj9DnqE4bcTmtncd701iI
fJxzaQYDLDWoM8+4ySLpIfZGNrya3z2QV1CvbxS02k2mDskPmN52sO0xOeOh28ESJQHa21JYnpI9
UZ/nRZwPTLnpZDL1KITK2IILWl7K8fgnkR5n8OuQuiHv0KLQuYYpVpYSARztD460QAGFHdbsHe6r
HWr+ZA+643JCYdFZwBQ9hdMcGCz5GqTyE0ZLMNMvw15TU5lQaX2IDa0XQ0Px6ZsPH+ZxFOaQ6Mzq
qI+VZ9OxNMqJFOg9vuBWMsE71kWFEI8Jt65BFD1RJnldRXYDEomxLheXhpPRoVF1FkahX0Fy6BT9
a3McIkaiVSmJTA5Mb2pqJ73/uGmWGdLOPbZRb5dSJ19flbK7TAsDpAISywOplqeeJMgnaHylcSqF
/oHHHOBHTXYfV/Y6lVShigIhebZxp4i1Iys7w7k34r1UbGBcUrIo/sY9sx1tgmnDIQ/J9CZPOAim
410O+zjn760X8XO9xs9+Xwafdoq8sAcntXIJIFZCwFH8fpNlNhpSNJK/AkKceRE3GnMTQlJkz6ao
ATY8NKQNf/XNBCSGMI2JbvSvKvpVxOGFWqTRqbZZ9KgyRKmUZJSnrwUOPCj8mpi7q0UMQ3AlPc4p
BeHseXwXsE2cRrieMmsISrYx67aWhA6yW52XTJPBxN5clzqNxnsDRpZj7a0N5fi3SiKu7GiVQaxR
8cdc9dxBnB5SjD05rNf17MEiBog+D132QjPwHW2C+mWGVL+oqqGlNYtl3QghPXdoRvc4WzVkRzhO
XqRzH0PLTIquhFigJIfOIWzyzTJIyMjGYbPGHeZNF2QxQpDdKq5bEAA2lB18xRK3mW7k9688gJBV
MWarWO8MF7tUfPxD1Ht+xq4a3CjwCKaNgR9sZQn6dVlmB3Kb/9d+B5DvioNR8fYoo6syp9s7Q4hz
1zdQd+WNgzjycR0+bERu/qZFg2tkW4JgvMgPeTqDcPNHcg+ZCGds40nmA5YcDVEK3lzes4wHF3jU
bE1aPF80bKX8uCX6zJN5cwWhHJMDTk0Z7lFhiBFU2528+GUsVYDIuw/+hEfcC8skqY50SbyHUlB0
w6iAU0w8lptEIUQe+79UrXXFJMbjdgu5MlkXvxz3ZixEGfJW7RV00Dq6R+x2oMxtGsZX2M0Rf7jM
6+dDWuAR0Rk3DlO/eCPdBXyZNTOKxM3TFIppkvMMJxS4Afz2hvM0+I4AH4ZNDq6i6fTbaiSXPRG8
1kE5UwvO+hAsMmWeAvfk66rOGk9gnBb4JCgheF0Ug43/+oBTwZt+05JvrRqB0hep1QzLiIV49NyG
IAcSCiz5X771K7EDiTy1g6ae5LaXCn0NNR+/FlV5oOrFM9wCsA7n/qMLtFh2Rrd/Oqen4mu4l6s6
LyZS6P+/RaILstDaiJKHEmAESRILeBfwRsj0DigW6+/ZlSjUHfY0D+d9a8Ya1E+59xFCmYyhbxhT
pTSDLpM/8DwKsaTLY+7vHbpgyrdPVjezOYkRoiu1fIpDrOv0P14TG2W7FT97dq08Uo2ofs+NL61F
avwkPvqlJrUYm6QTc1RF7IdWlaWVRsBrJRisLv2UEm+HSUD0e1Rt/yCLKvLgmKbDSIV+QNKjTIa1
ztLFCJtQIJLY7YA5EIJ8noUKKyfqoSgPDE8gsMmijmh6L8VY0OF3kLAnPe6ZxFMSUESDql8xjUP2
aW3aqJ+rmP0KAmJbfLkzwOFLF+oZhjrJkkGk26QepTbYj+QviMj54n8ttb7ullS81ieQgefQgBCR
UGvxHr5EJHRSnbIkjtX35xC7Cpu75TbpzWYplt+tORTZp9W2wMSc2jP07hhg5UWuYgUwMTv8eGG6
r4qZ49gUCCoK3VFoLOAeC94MgSPrfZeev1vZI6Od+X1R5saM7ZK/52Hsl4kgYD9rjZGIyYUWByPg
zXcNs7x94KJb+i6flKn2L07foqJ1GtSSCSIS8T8a9dhyW4wbI52iArh6OKWMfzXpVcYNvljcGAZo
joume4Q3m2r+wwHmfM8Fpuzo70O2j8fKWYkwTAV4PDuZjrUlw87e8l5R6N4PNZLKaeBbi3Zo/c0i
OJ+88E7ns6X5yw/d+P/dQZd0ClrO22/DyNDpLEr+1V81hmuHXx2b/aaxfdClIkIBGrPiQbdyh4qw
dR1bfTpP60SQPs5YGk5MFov5Fm3y+F+2hYq6txTYfdXAXgc4z3kWxqzlpngZYcCYiSk5O+aDQ0wi
nQsnq9sQ89N8xAp8HbxLs7xbSGn3RcP8cL/NnNtVTeRTUh9cG3bfAzQPJddbf/3jiv8J2YQ+Zwjz
KI+D2gAWgByDPhIv1HYV8+Q4YNSNgNQYd6dAxTpJMXPsA4tuie2CflMY2zujxTh2A4GsOsHCJpVX
dkU8fxdn0wpMnQoHapDvzQp0X+AFfEOwXAUX/cavNH5R7Ab5Y0DZgUWjMexDqAdtUD2dw0hZXUSV
ayyiWork5zkkwgY23err17OotXmERG+CjaEiZk/Ei10Bf8gpS2CV0dlH2uybCol+ncHPJ/MGYE6E
Bt2G10pZbm0+/S7LKktPBiLMW8tmhF8pHGiNM89Zjxu7bBKZ6lkHunwGr0pBQmzAzC3P3Fm1rBq/
OmY699CnHDqvZW2vLWl3+zGZx/Lv40xlXs+P1V3dX5zZiqokp+Za3yCFVux3KIVQC2ktyMTzRx1m
xW8zT1c1W60XLXK2r9ERqdmBRWStehtKKuTVDVCDY8aUIDt4zAP6mgdLgBSCB8/0dZoSnKHcrcZ2
ygRh3qnwygtnrX+M9MZTQd9wYNHm+xXB6OSGYSxxL0PZEvkrb/4yLZIJs0h6eS213liFjyFGGBH+
7OnolB8q1/Dyv8/xXXty1+2NKkOUX065XdNZCYkz0gABGsDzie9ud9Rwf3vOKZgtCTdywEUf+Rag
PWELnUyIictbtDhO2bVXb0fnPMsb2go9XMoGzcRrmSU212hd6jsbD4TWaOnenMIxEqZ8p9h+mTL0
0S2QF866xnmSdU0QX/hXJLG67JyojnBVF2JPylW45vKjdnA6oTtqhnDLLUagkxRTkR3iit+hrBQI
mGOzDd8NzMTUZW/2DYPvNqlJCBaXUS5CJCmkM9eWNXmYlJWyHtS3Q62/1ImAk6NXYCk9kc0A8bjZ
nHNACmSMOs46w2tmPrj4nMip0UvMzZqdB1xStPlCrfV8ZJspm8zttUW9z9oT0BPjFs9DlRmOnwoV
NyTwAn7jroJKMI79vefySaMx5CFKf62ULhX21qOjx1DuBVP7NAZwW/mnTq5qJl7BMJg9RYo0n5Q2
lSsg9DlBr14amhIPnCfGKLx5hIJqknm+EjiBwiO1UvBl3yrSsDRdF4z+IoOt8ikkYBQiPtIrGVqy
VU+Z01vgdkGI6oVMPxwF2ehfCoo3WyzLtrD5jb8bhhevJZ9Exl3WK0cyE1XVfQO+3TWE9Uo/DWkT
w8KiUt6ZlJkai+7yZovZrvyR61FUeQtZQNwJx/ksP+Id8uMmXcdwo1LMvMTCSLs916awV2a2d8vV
fZ2Aga4bbHK49rdRm8xPZsSuQBnZURaWuwWiF5u/hxHSV+6OlVgu5tPRaWWcMtyHM346jTa0HRlj
xpVkyV0PZgkwcg/922IlQYUIJZXwu0dOl3RjS6UN93QK6a6lCBwnwlwmDPrVos1n1VV1SFJPitwh
DjsKvBlgObULa9a/aHOwjxk4yvUM7NbaR8AR5n4r/7lhAEwi4UwAZv1FxIIMr88Njcxlo69vQQYG
jB0T3tpW3KB/f+L++3m/qgfvcmIipTWz0ZtIuMiZXdXLYHSDKqOVzGxf0uFumgPbxHaSuN7L6zgZ
97bnx+3pza1w0AGtRdZH6WpW5iCXwEK/wFX0VrTrupfYq+v+dgWvSgMIG2sqWeK/LOUG+t9liOVo
HchegMKMh7K8mBSUCu/LbyLhE1o570Lkhz7/eJkW02jGcIq2IYMgW4IHU+IAtvH8DowaAMROwFmG
o7GxQgodSjS+imsY3XjWipd4S0LGbhXie2nCTzPSdR+L+at1zMhR6JPRmppNrqi55hpqobILyeG0
RS11adI6WuBrhMQdvKLZ4X057IOsVRbjDcZU69CWqdMWbD1HVxeD+BrewogYHfCH696wJN6a9lQa
7VqJyf4kohCpsdzNjX8PVQ+KX5LOVeAKGnI6cVxvL0VibSQS2mbT+WKTRVjMay+1eRkaYLy1+kWT
fdskqPCRTqPgVRBUbno2ZSCR/v+SG3Q8fZ3SheSfjWurfPFnvQ7dXs47NPPL7vZmrnvgUwAmqbaO
Nb9dkmGYMh5gA0A0N443G9Utzxhc5pPeoe9VC90b/n/cSlTDB/zfwy+xMPOM0VKtAP2cMC/0+iub
kxPbssAX3fVtD0p51pYGpCWUvFSQIsHbBjA5HXoKsS1h21mD1PbEjKT9l18ZM8t+XQS96DRmqpzK
KX+gV2N3O3YUP+dpjOx1dpjO5vsbthXomEytaufD+xFi/32rtmtjL4wxl+HxtH1320JwVluoa4nD
iIRvY7qQH0ZflcbUyh7MRaLJaNwnX5fb4u2OydLmyW8tJc1yaTtQMjIPYV/Cf/b6JLA1DmHEb/F6
+UpEazxmQK+nwC8ej9CI6rgQaWoD54+slZBUfYplpCgsDcIu/UpO62ROVL+4lTidtaBQdSnMd8aP
e3FbelnXZW5AZ/mgjcaZd5N+Ph9wFgE9flwqchX0jBDbEYb8thC9G/kxUMYhFf4HsbdZ9md+dcVR
CdlMFGGaC5gaGXZxw6hVCIKgCyWXqwuevY3AKQGRNzrckJSjBstrQSR35eFQVvzSGYcZhqkHDvNY
jSifFAOI2ZRPAdGbMm3SBuequZ/1Yc3XXC7I20rWSUVE3jPlF+DQj0PiLWzH77kj6dcuhU1xGblp
SP1vkU4PTk4oczn9qc8dktdSJtv80+TvgraoR3SrBXBg/B2PMrjgIYFtNvkfqIUeCaJHGuuELT3i
hEv+JJCUNJavcvQblvyR9YCdR77qokbNCOZzmko7qiLUmDNQuR65q87pSs1oSehFIrAn/+3LJEum
KQx1hRO2iJvMRvAc4nEZvue3IitKtoKMb+RIBfCuAlerkhzY/XPk/rjGZ39ohM/Mdmrtnh/NgH8u
NQhFyCfD7ZABU6qtYP1Z6UL0XiIdz8Sam+4mYSXRk0w4aYCMtbg40ddyH5sdgA1pohPiP8rukovY
TT1YULOuZM+voNUwK4ooxJVyyvHOqSc6CPn/wnlNlgfjhZJB3DVOT/pwUAMHICq+nIiGsqxVg7pV
LGgWomiANUKQZ80tqzFLx/jNREN0ZNKGzsBzoHUu+aVnf0Ze5xL2i3Ju9302wZqiU3RQY1RHc1xn
+xPnkxcp4Eh9B723NXGNgVCcuJEuCPgAMCK9VLl2h28h0bJ+XznWyeXMRfIS7OnIsJjBwdDEPWPE
Faj8YSx9syg5fMbxdzqBQEmOd3mgD183/YPxYHaehuEm2EFdnuwGHzTUbtnnJSfFn4McNYdQqZMd
x3wah4hOGzZdbQWfhnCMJWfpU02DkCXmlbLBrITIqQplyQYzptoDIP0UJaVHS32vjzpEzMB35PDY
FId/3bTrXebqN4NdtxLX0GiLoTMtYNOlxSGG0Ip7VxiZtqQ4e9lf5bGTrrtT/A+8J4liX7MeZgRQ
0G04wA5C/8N31MGy9NJDm19jOz7U09WLxTOXrt2EX+5Se/Kb1Z4aQYyG910Kn9Zy2tUbkTeMoffL
JJn6qiA1s/CTqoxWb6BccUORE+0xM7UEalJiW9J/ix+5jNsjNgQLf540GgB/xN0rdYCWhDeuZCTu
PqtauPZJPLTPrynxfmQ9UcE6ZgciCcposBb+JHcP3V8V3sdA6LeFHAuBUE7NFBZOoe72kMHDBmSE
pD2NflcngyWtatZ3pfAd8BjLKedKAn8P+1cbLkcNkVtho1XYe9zDiARB0sORNGl2cwO+yyQ1nlw/
pRj4rHVjvg6AQLGZzK791BouD/EKnnV7LQqHAc+5I3TjPv2D47NU/4gkNnwlbFNfe0EiKMWRcScE
V/qvYlelnvqUghhq+NWa3Sm6B93DlpgpdH/nE9MiVkyDU5HftZ3u4G0ATggL2uCxB+owuBRm/IrO
ud0RYq7zIzn+SLlkIsH0hYDqjweEiLpfAc9BY35rOhzLIskUEkF7HfWz7KZx/1fqLeubh0NWpP4n
sA6pFVB/wvWSJsG3MwXhmYJ7EJyVfIxMxu6X6xh+1BaZpv2i76Bu/P1gvVvydPLUDB2Jxs6BNKE1
3exx589h06isvNx+4ABa6RPWDgPpGCXpwqxzwE5f3uanPSSNtcX6R5pso4XPNJavCWZwqAsDSSHU
8ZrRxRdXuEgoQU+pKHkBxv0DpAcK7PABZIRX3tJ6ukAi7bgAVDaaOSvmOJmtIv08mdrx9hqHD4Qo
O0+x/M/kkZ+Ki40o3AMTqZL4ZuENadUL5IfW+olXj5E6b9v3Vb3Egpl6TJQbimDwpuGnFm+bYCPT
kvnzMkkWGqX0b5EIlANx1ybWP8+gJbyxa53j6hu29ILRf42ek8cXBoWzgjgUKS4we2Irl4qWV/AN
mKf97mgogn3gcV3wE3TLhI/PR3i4wqD9yEBb2rG9vA6BM3633Ssb7wGKQRpzKOYDHUrDLfGEhz+R
bZGpYAkHRNQwekA0iZlW03EcdW+0kIEuU5XBNQmVyCFyVsjlE3nuHgLg5v5xwiVThLPfZaKU7N9S
BVVLRQoYZ8VURzlBvhFXfJH7LSsnjSMUku+Fe+llEYL/dPuUb1b/66sYWDIQil6o1gcsUxVkhbNx
S4ecZYFnACW5+KcWkcP+HpzAgV0lYPYb4b1iOQKQ/0q/B5aIsdqZ7HeqvDwm+a6i0xZ7KIY9zWqh
zGgDGeCn4vDPVBH4nZqdFmxDjE4y8xplBeKuAalhNj9iFv+d+yKYKf1dmtDQUpOvek/1yujlrzZr
MJlzFSrhffKsEfagn6yRTQ9n//tdICnQXE3N16SxegfIZZTe5Oos/cDW8iM4efRQS2Q6V4eblLcD
4HiQV1vFL7/squdxzuMZFKwwsvACiYlmF7CNHFJJ7KrWTyDeizCeks8cKZf7pZOBkqavnIAnfWi+
o5AjDqRuOvTGe6eubKN62sZq+SAB7AVu2k1+MQ3lsDkyqgdfMb8QT63JDHdszRfnqcXafyA+pBbN
cL+rTq2FBeUKO+JK5nfFDHTFkBdetRmCmeYDaOHHdgJR4P9bi9JfwhSAi9u3Jctn1ufx1nw41GTM
w2RzOHPAlXP3EQlI2Evg5n6KaEdJVhphFYZb4JJ6g1sJXbSCTg1v6E2X08+wbkVRPyeb7DflV11j
utQ7NfwSqFsMQrFy6Yx9BmIVLJA1bMXCYFe2vUx3496ndoakjfN1XyXRC3+r1eKCqMEM8xgCGLst
jeW/hQghe2CpBxrDhEhmNpjRW4ZJ8BmMY/DMrUjM7Jk0t+Vq9A3DWw5QvDDml65XlGtqYjV8iKSW
5aGx4sls6vPmY82/waTcjADe/Veb61Iis1mnrHPDUvwAjv6m570okupvVHclzELCaNGL8L3vv2pR
HIeTZIEoTe94tcathMxIB53u09OhOe7skgHWTy/xvX+wQSGLEZ8Xg2eCPPcB0kXfyxBUU0QbuvR7
yjdrzXxDdsH000vfGIP/zwVf3b5CAEf+4J1pEF9fjAN7eEKN94JTBLEPJKdr+RDQal+fMAtZPRGW
1Mw2sT1pJ4Ulvj3QRXjk/cIgU+p9i8LkW74r9jrBWb3YxedFblrC52z9RaBBA6kSmwwipS2U2I59
Dq5aHrdWNzZPh3ethlBVUn0uJDIlBoEioGpskK+m4C5NBUFXuQfk6FldIVZ+QZHy7QdXIucnnAv3
QEiwQfW7HwYL/s/zBh1BtpiA7UzElEbPgn4hoJOlYwIMcV/0D4scccJTxQy3LSbx02ptGCoAs/0p
7dEKN64RgenKmRKQeW4LauKi3papd1useCbv9YWxj2mFINTzV6wogSq3FcnTsGyX8HbjEerDW2+g
naJXFG2CWDu8xusGaGdkoL1YlZlvFMCre2PmFBydnboqKq+F+NQyQsziCwQK4GXcFmmCafvk46r7
6tZfeXi4VHCaP2lumUzPKOb/5kQOLyaBj67jsGWqxw40a1OdKUEznHpqjUOSIwOw1kJrp54oU1Xu
MsLGLJnkUDMQXvIwmSpB+yIDXUEcBg/vh9xxLzyBEBdSmyh+XFge11O/pGXQVMDagoptNhV6xvl/
i9wJg7Z0X3hMzmej1ymBM3FZ/uDZDchGu8ZqkFGG6m73oh5c2627K1eoFliqdiRhnc9G4zO+YX06
QoENq+Qm3ZT3h3YA8hOB17BZUXuECXnk69jmBcSwYXhvDd5lsbz6RzTQy3dyr7znEHmRZsh6Outt
LMZj15sIRWzURkYtxGEL8FC+X5YBbTU5OfCBuDegGct1CxmBCib5f9BfBPgXxozXZhykRHWkYdNg
Chr+X6/avnfX+cudmhaqi9ny7w97Tz+iEmcfkRQ3k+kRKtjcekUNLqmbJYrv2GygwdiD9Nphcr2F
NEabR8N7UmF2UJA3xpTjk0FFt6dhqkqUcetADqtN2reBv+AvD+MKZ3pGZXsdsge0cPC9UzrTnjGb
VehJvHlzWhlkk1653kGpoKH6EJPv4zY+qH1ObrOT7PDwI2C6+KrcBieF/Y0E2F7DM55rWchYlxyb
/UAgpSn6Yvx2sx7hy3j02oMnvWWfX1P3Dy8b3KLEkFseD0c5CjBnX2ZgDyzhiERmtiSQdHPGHokW
n08MnQYAGMqwcjKZBrK6PVSPMz21KrheppX3iBTIVjHd+YytiKUyNhsHmCzzzFnYgwB8YpkuhZI3
gKtyQD4oYob2a3Wxi8Fw2olYUTE6VracX6pIH/I8rRP4MUVBs0eR9viXcUZSAqMbN0NV1eD8igaR
n2gsyigw6Oiw+p+Ace/L5dwvT9XISp0Y/PCCmCUsiRz76zMWZ4shoDykRoyzUlFyMO35wuLGUgmf
jYMf+TPSPqLi0LpU6nWO9KBFfD4dfpkEfvGTEvqKTpQEbzmgsrYHrWpWxzB4OQOpiO83THmb6GQ7
IIwX3n8glaWnyiQcVPstrDdezFOonWxnLt2wDddB2ESZJ3dFp7DsUPVaUphtcUQJ2DaQ7A8OliZK
YcBIYSCEYm1w4Fp5cMHjI/NnelSSU1lZXhRlAxnh8Xt1p3Wvc13O+rXwj187ji0bjoOB2QIGROHR
g/GilA9ay0C8NtYPsmLx710EJpk7tPr3vzkmBJxLEAZhOD7r/DGanPl6Yb1I5Vl18Pfyrhdq0rCP
ILkI89nuCSnBwZVTT1yasguJFnkROlPvIRlqmCE8fLl3N88jnESKjJpn9sZulo4QPJYJ0nrDuA6v
sr1r7efclPZJ9LX782XYFlJ423ZuMmkCkD92pNWmwyjhBVF+9S/bSuy6CrVG6jrM4jUekS5EdnLL
mH4j5Vcn5mtkI4F6kbZClREmKUXY6uC0k1gaQRf63ut+PSlU5QWJXXdljrCfmayBuQzSFZX+DRPB
yBFL6N3NtXMkFxa2rLBFX5wNknD3bnmjNMIFkPbW9kjTZ28bKri3fjKkgbkWgZsljwl3SU3zCyrC
Yg5yeQT0JDGG62DYp8q0XyolMlWhpAI/A8R0m1W+4yfz1Lv18ELcielqn6Bz8UuHT+j0pNnoPufd
Bnd19aXAHllVw3CeigTV2tsim8d/2w8SRSK4Ewix/RK9qUB21gV9NHZ44KamrObi605Qx2pb7OxZ
84RQraX7i0RhgaoVL65aExjLtOZoX5r7Y2i3ZCgEflvsVNZu7z0tcYE6vRkh0/j//9G7iN9vR5HX
S29Kdomki6u7hCMQayYmKJDGqnqllrA/KeDmM5iXnh7aKly3xkplCh+wyAVBOrxJvpkl/rlOU9R3
lg41mXsScCn9v5nVeU6geII0/oqAjksVllhK+NznSA43Zps8fhKgRUCI0md6+PQyNxszPpryVnB+
l3/zNM16Jtt77iuzCjvqwzHQHYtCWeqAwuBciH8ubstcGDOJ2M1IlSbJui4dWyNcfi1dkpf/H2Xe
A6LisLSpnhkgWzdx4A7sAenM+97OMSPd8P4zDdgagsuB476wFlX4WtMIhcrBNGE76lUNZrMM9b21
muue4MUJCk7BEOE30JhMknC5kcoIPz/aBa9wSMFSp159UPMXH0YbPuzuS+RaUt3JZTJxsoFuRDs2
t1aUuyS1bQ5AcsSUTB8qCYlDSfi982HW1VW0G0JtZc2cJrfSk1/e8hhKXbklm+PMnCLsfbRdv1c/
LbxukZZPJxOMJstrVcjyxhTYohsQGnLcM1LdO5lt6Jqm0AsOwzyt
`protect end_protected

