

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pTeL3lbzyXpg3zBlG8xXBsi5mPcSaOx7zOxONTRBSW321/dGdDH2TpaC43BqFdYZqpUNj4ng67vZ
qArBG995Sg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I0+MKhxg9FScVNavGFQn2xkzaE4/JyCe16C1b5v3ObJwo9nXDzI72pLgwgIfWMASSmFXtaAAw0ml
3uLnAPMYr1dgB/uJGeAtmT326qa5BMsAV4vQ1Yunxch6eAaFBVMMeEWawv99YiJK9jkH7yDAOpb6
smI54SxBdohXuGVE7bs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bDMpPv/P03hJ26zOMeRntjG40FHNolyY3dG2sIAWSb+A/C9vMJYUZduiM8NsMGgn92oqltQI8itf
kfh0mxfLeub+eu7+DutH/IonvZFuvU5PDOu5gXDe5IZcX7PKYSeWlg23QrTg/K5l+bblhZE0trh8
gSCxX9Y5M/tKkk3Ah7QmsxFm+D2iD3pm82WCrtLPh7JqPCGwGw7ZkIH+rqgZe/fQHahkffxj0VdF
wp7Pe3wFKtUoiMTg7uNHWsoKi6g7a0GVmS4unE3L9HQtqDdu8p186XHZQqxkv2iNX9KutOONjQNy
x1JPQknSlGZ+dd8WmzTlL9rwhQHGdMhFcdrMGQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CqlfcKpSPaBiicqGT47t9PnrRSQ8njMbqaZWYqvnT67KXQ7fxmLQJl9EXGvFoMEq5tU8J3rLbBm4
9pWLf80+KgxXgS9WPEn1zRTKt1wiye9VOUHfewp3QYM+B5lPR0EENtCdssVC8DxPUBy9Aythtbty
2YxNBkGFMjMRSnj+A14=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jiVIVHHI1er6oSZsM5uji5FpVlbZFUX1C20PfTXKPYBzpAjDWZhROWc8xFgszwvy5guzSmUMWOgw
XoJ7z9N2ElsO0s1NH9ojznzy4rNB66tyJa27TZfjI9UYZ/9rfTzXHnlr6WpUX3IChRrS6x5LI1mY
orERQz81jyLKT8cB3O8KkjO3g1Ks65ZIeY+E+7T5cJHzOHJQcoiTTtwLajrQktJS0RpyUJr3VZHu
CSADq9QNuiNkf73BoFHvperz6rZhWbdV5MnpWKfmllMNlSqFwzZuWbMdZs7ZNbssXYmUZlJVjM52
JpTXdo1N5lXyKjXVvDlv7kCHkBmnfQZM3rMXlw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17184)
`protect data_block
DnjljC+5xX1DFYNkRGxZQqdKsGlJ9HkHwKjDL7mMdrbGaOj5JzeOTbKd2uf51gCk65yBF4n2Vr3s
ggQi4Vx+WJqsERGEtu3tByLyupP4irA6QpVP7tjhTDYMftOeClqw5Icuz6X9DxcYMZXGMQY2O1U0
kX3H7XErQXjMazKHX19O7vRdFdkTnuQtyR68WaOn5SE743GYtWoJurskVExO6ABsBWX5VV3hypVN
yMjiM7fdaEG8ygH5KZDnSe6bhbHqEJhQv9wJXcclIkKyT0mORDJvAM1gy9sZxECw1Ifegj5NZ3hQ
WLswjhiPtCFieEXvLgM1W8iTFOHlY2+T4B265csTY6Wc0rXh1N5uTO1yaEzBAj2Dh7Xcp7dOrLOc
6E4Y6cazYaKuUHx7fWNpO1qhglOQ4S4QaT8Zsrxh6nHJxV/TQizYuhQQ52cURQFT4SzfXD9oLeeP
R42URllv4GilsDIK4KL0Jc4NAyMHBvRYLRrmOlzHk01GUd6sr0QlINll3nwf9YJaFXubQUelGA03
0pmcENRM0DYyl55D7/qKpZuoLNcrzNnJ/ePEJOd+HaBvHjOdrpn941NpN2/SHLjdUFdnvx2RpIDx
fxFGx7rDUmiLurhXQ6g2UTxD/JyIsC65RTfRu6mpDCKKxcMI0YWP1EN28pOf/0Ym7Ku4qFC1PAUf
jpDciK3sn92Oakp5FFXaQGD1wAzke6FAc2GR8USGZRjEQoA9CeekShzxVZTDUd8PGxsj0h6M3H29
k6bdc3/HmUpQL/db8qSSjPA3RtgaKlGDmtksUgMXbDBp1OiHmpVRUAwGhoWH57MxUkmQnBoF5r7h
aQM9m/xKLPCVBNbZwuB+6HFAPjvMShcBHW8FZGuGN1pddjNCPNbX4/GFZvdkQa/HXBD2dwAOmg8o
o0uIgJEhra1k+l5WGLtZs74amtopT3MApfA/mGeh2iV3b0jSvoFlQHGgKrR/4xQyunILLgQENUZO
c00bDx6j7mrQeBnlAir29tJMji2VtAKQshXcoNJxaW1xkA92/wOzSlr0aR1+vDT320hdY0thLF4z
p41vTEh54rYkCq/KNSdn+cvz01AseqR/akUv2FX7oBT9SEyJL/ozvzfF6KbES9G8WWXdToL/wKlI
urcVtZZXm470fDaSwrI6+Rx09IjgWFwj4QS6YJPt6+NHClD+j8jYqX1AP4fobvtchjfergusc1Jt
OLxCvMoeEXJVuZWV0jOlydL1snKc2uD3Bs0vT2pOD3HHbwTnuMazVA1Q9EzD80AyWrGiC+oRGkyz
Ki//E8Zb0tRrc8XQ60m9JAE31wG9MN7/8OPJjwo7+5J66UjnkiLJokO074aKsiOhV6FkBoz0nraW
KpTZ66NaWDA6y9HM9jFxv2kMK3UdlRbAVgdsHvHILoIoewV8PpFSR/VVMY4Jh0YKAMPaU/h7nxMg
g7L8zrJZ8cpegJSqPEWwyVhXVT0fD6tPcqvqgPFzl2yRg+JAVEuKsdCF4oGfQiW2KBr9i78suEm3
tFaTJTBk5PmnE/NqIbeaDr4mxeeyN1fV65E6lI9oJkw0irHeaVFiNPFB6SDVLtUUZgD3Wjq/31mI
WYOORGnwuatR3AGm2VU80KEI84PRBwMNgPy9SjCHl0yH4OpFhgvFbq7rMdzo7SNqwSXVaXPy7j77
CIFvmRvcF90YWnnqPO9ByC5sGBc0b7XhIGAR9nBcvreCDJNn8ODqXq/hNyD90o7Wym6F7ByPNZTK
BU5kX7zU3YBehi6mSEeaa9ImkyWRNOJyuy9wxbOad0JM4lLpwN89tgz33giI6tJsuplDd1/jveWk
RRxJA3YI4csGxlYng6L/TEsxRTeJOmCV/i4goi5rRHXW7BfVGniNXl/YKyc8E1CPGqSpyDG6l8i3
CknRInX3Ka2P5XkHHuGuJM2E9nv1WABW+6idgj8lFRscn6A9Qeeqv5T6qG4osN5Xq0i3EVviYba0
2HEF9+J9zffMjl5B3jKdm+jFCBhYU7h2RxYBlmad0lBkFllMXsbPRS9UsXB3RVGkYczZEtZDBWj1
C742evt2XOx1ej9nkEwo1/iawxEHK6bP8D7WE4YxHYNr56i57FtHHX22JFTochaJny06rVVaMsEj
ojJCbtK3kAh0U1/1JtKvOP7FLta/8uR7dhkwyL15PlrhSUsU53URywaLaG8yI+9kXCBBIqGT/oDh
wlxbOcDYwmE3sLJVxTgytA/pKQwVxcLWnE/EscP054ilTUV7n3i6tcw+x/aQn5mE2uliFTxIDqQY
y/YkZQr3cucfIEoX4a4ZYge7KlXjPYDTLpf/PBNoVzO0xz8xIjNT9NwNpFnQZ8cEVMlDaMXieq18
KT87XvtTo1wFbmVwAr6IvligDpinTZu5EwptCdB8AU4z1HXBmTUs46i8fLAyvo/vyhSuNLZB1tAV
FFAnXIAVQdRGrjYspKU5KrELGo4B5CenbmKyFnfkEGvg8as+UWiUz68aJNa5A/6vAfIFjYx+LuwB
TT9cCCQJcPOGAHXUEZo7KrjU5rb1ofyZz68NlqF4geZ0uC+Zfw/PvQSPDURqNtk0Wtd7OLYjujc8
fSYktP55n+MO0ChVuDIBmk0AlDVTTGwer0dJ6A9m+WEso1fs1F1qXkq0ebxf/Y76J2aXWnepPFjV
Pc5OGKZXCeWP4heEJzAoubmDIR0U9qfu5KB2rDtnm6h0PfFFdv9oGb1BeKzcyjtKGCX2GVjAlCPx
Xvir/4wmGU9WpYR1C4u38hKYqxPeRcbFz4raD33jG0vvTssJoQABjgroK2r++UKS2PtTE8nLmKgA
Gi8ahestRZufXuIT8NSM78NsHQZm2aYxRoPIZt4x3OavPSsg4MViZX4Bfcm4uPvacVafoTsYOfM9
KAxFFVHUOCZctZ97jZsC3OZN/+9ECpThEtB7cOX8un+4+gCI1CPwYte2yOb0dbJd5EZmvqUMVaEk
oGSqKj07EG/Y3QIc7kb+RmkGYOyNVWAbTL0hx65KxkCMIKuUAGrbwpDKmUxPMbTzui7nCEZJMwr6
RKO7VubF0c5kG3d/6oJpy0jkIrIsPwKbBpdQsb30RCdRKEs3ZYXImNZUhoHAS3/GQUc1dyW2kcco
ljsAjI1NMmLFaQ3nZLwJkldjPKI6mGDz7Wp82fte0IhgxkHNRvtE6E8MlQNBRlMyL0GPkHNJjvsO
sWbsCJ0AcLLNU5+FbVJx/vWV7l5hawa6rfXm6/BLYAoxI+nVFezCiS48ZPKyC4m1+Q793LXzo2Xd
4J9ta2a4bfScFxEgxvZdyyvxPczFQH4FPsnauKmCUpD6kP6LGhJRUlRm8gCq+2Niu9jlef6ZZIWK
4OR9KDebSXQwaSzL5UXB/0ojcBbPpFz3a+lgMvKE7+jgZKw56ZXeDDG3yTAlkjCUkbZCKw/K1yeO
qb93BGp1S48QObl71JOTAC+0WNPPwLWjH6mHI6p9chnt3MWFj+L1wOz/hvBR1Qqfsk9/AzVfjaqt
1fyLAANF9fFdmBJFHD4AmwfPxuGoq7GULs40I2IWahSihgKGP0EWLlErlteVjZUH3vovZT3Af9h3
fqgxKrOAAgEnklzhwLybVIlaxEJqIO4ehA//bg9coZ7EnqWtUIUVpUqDodVMVc44Y94wWoV6TpbZ
Ncl6SMBCoDK3xquYm2OYr2sCVy/bnK667FYe9o7tQ62UUobd8/mfgfTWFIJsDaDrBKH7XQg5rQYJ
kmMacXXHgOJwylKa6EerNEaov9xa/MQqZDkl9BayvZCv2I/MWHWdEDaiS0DT34T+jfxEwYGqXmyt
KIMrCNSnVvIyA348YNBpXOKZiLs0I5gyO4VJUSVfGl0Lt0SUZMJwGxO3myNYpQOT7NROUOCpNp5h
nGAN0SzMYq/LwLc9jNS/iEJoCmSZn7HhZ5oCAp1g/POANRnw13aC6sVFO5TaGCMr4Ao9I4TvE4l7
jSiGpYY1xzRZwqEmrY1HO60q6r+CWrGH45GJ/Xm9sN1bdWNylf1ekTlWgo6T4oip7CW/lGz7y86K
JwBHzCBZTbqKUvl2MnRi0OirO8/uuHtYveWUhmt5K3LiSDS+eBK/I+7ztFg/xhxF49EMlm2uG8kS
WEM3uQ51huSh/ebpE82450VZVq3llinXiSNzjVDlwQccD7Ms38y4hkIXzGSvDfVKst8ctyeyGGAY
/tWDo76DfZVUFCNyhLxUjSYlQRXV1ccKUHhLjpk3fjD/rZrI7Rr11fU4lFlN54WgLcURLfpUkhY6
dHDSwh5DLbQGmqj32tJ4w5ogc5o9C2s/2vLQ5pH/S9P48Am0COHhZbCyyMmdBgLl9xY81ncMns+s
qpcfqyjbbcbV2lG4QIg9ut3QH7ZQpP+XjjVvomgxKfOVp5MQFm+U4FEtknCTfc6jr9WlL3ztt4g+
q7se/vmCizNmJGEDyuulTEhixKTuczNL8MPXMk2A2bOZnxXcVh6xH8vSX4W4roo+eB0A3xng0act
Q738Hfq7WLua0hzoc7wbK3OmHgwgB4ekUrHpnNP4jZf+ahqm/cgQcEt95QT4br930pxU+Zv/nO0l
dEfeI/JWdvSoy7lZwAuhCx42a2j+AMvj5YvrSmT44k17/BtlDiC9r8xFlbrFj47q9GvysTsvkkyY
CD2HY5RJCjIp0nKo8IMOYR9pV3Ixdysnb2mCg33WXoby4+8QiA3Au41T82+dPcBjYPvNLuWdathj
uLSmzFFtRCBBvC1NEYohEHT6mwRHuGxT3smP84TMmdUxNW6xxXI77zwtXznIPHpQl4OwETTuWpT8
uhqwTuUvQz0/Uwr7Bl8Nl7IqpIGj/dzYAWCH0M98RzxMJmmoOtaeRmnLcD3QGiRwzSQBttWsZH9T
bX/g7tQN3eozXp5X/TNGeKl/jNx5yXWYbIisNRHz9xIZGxFncngj2VrsItyB8KdtuWJYxMEHHpKk
FkRQKuBHa0Lb3kBtRR8FCRJOCuIfYjz+G6Alx2nX6PxK74vIECPcF/v9SR/2A+nQSoNvc5g9R16o
MfuGmyd4RvnWMEAhNMwrGMUrLltoMW3EJhS4CiIkguaBN5uv4eWYww/2UZ77IVQUq/Wo+aQedpTZ
DlETXUS5fsz1cYSb9oxCo7n2auLCpLDmwwklRxqwH5AMgWA3Tx0SjEVh6Iib2XYa71tzhXNtLM3z
o0pvqxcnPeyTusRuOdJQ4ynwIr1va5jsgw2EiCatxQiLh6/xhdstel1zca5JNtNY4MvPlwsuKHGk
4X+3h04lCwHHyTvZuFHlregI17+KWjT1/w0upal4o7qUZPFejbZt5T5VUSZTCHSE11IXGNdB9QVK
gNpZc03Zu71SJTSoC/uA+vEeS8Hh54M1/3qZc5k7zpwQaQqT1V0OZGCH/Qn4p8Ylvv0+fGS0PPIl
aL/aoZyueykclxq9zkmBhM6f/NBsxf+Tm27bSXKS63ckmDe5YUN4CZ3pD9OFjkSjRz1YJ5RiLttc
5k5YkG7gkrPzfI9eNn+7Da9uxJg24IgIblrEaxbwpFp7CDgDjX+vh5zWDSWkJwDDGZKu3HcIb8Dt
uVy6+A62Qg9QEwN5i1jo9oqt1+tumREKwaJT4CFTfNUydQ1xT8opbnzKsu84Lffr5KPoOoL9BNXa
YPI9qjVPkrao3Ea9Kt27DtJp/uIjukWVHTgrEbSq5usxtL3v0uH4L1gpTN+QEDBRN+eoFtjetWqa
CXDfSoVpsugcvkNeHdILDiWtAX+FZHx+XifkJfW4Z63fDDMRnf+yzT9o77KPbkP8mgwOyxxL7zbT
Oceu/EYeoCBR7LzKJfOCqjK0Ax7qMuTMcWJ4lfqHT4cd77yJdryR7c0G42HU9bffKE1aDxVi9diC
mgJ0E5pt5WUCTWyqr+psn25ZM7LfZ0Kersi12IaCaRy5nV2DuS4Y++yI362O8pUL8uXXtI2j7lDs
TFuNWPX0wNlDjfm+L7kduFRFbJai6WJY5bCqby7zrfId13jAvqfDA2kpS9W2C7TQ5k0fGS+Raih0
9gXJNdNXG189E7aIqYC0WPsPjN5GIRygMPIME9O3mlgQs/01xAUAI4B0u17EIBsUkEw42yURWDMd
xA1R/ZBPL7F27sSsjsGitomrb14dC5PXR4awTZ89x+CbAY5eaPRQ7OEG7NPRSRXoegv/aBkHhqxL
Fb/VFChSlm+NAipBZe/hPXiGPiO1IeCWi0F2uAW58kR2C6f1o/oLP7h16n44MexzbKbDkx25jam6
WlzD1YIyEcar7YL+OzZywBWj2GdYugFKte9zmR1o2kwJspNV6OCnynbivU0eqLLeZ/gxB6S31B/c
VHHVchB1TqS+W5bnYn85FIby97hH7E6BsMFRGZsP7n9RFep6BhMy7dyVKaWgfq8UWEPqDGX2CbNx
pqS2aDTMvyEpCSN4aBEEwJ6D2TND1nDoRVKylaIN4HbdPM1wL6yy5R75u1yQWPnfOuBKONRtHT6H
eYPrUMsfMGnoPaiRAOLhy2TatlUzSyT3aj0B/2aLC2tT1dP+pYn/pZus6lwsSuMMEjIR8sX/kF2R
3s2Mz7Gzvzey4uYstOU9DdQxk02EnX7OYibpmG3jcO3S7dcUu2VhCGT7hrFt5ZYfbGE/Kks8lmpT
TPq319VkY7F+UjQH/1vELlvcaXJ612iLbRkIvHwcZ3NBS8Y+pTJhMaLWb1P3KzoHm0rkE72FTyj6
iVpBhA9p1mNKq4iaLtNC9v7vC46YuLdZbkA8k0njJ42/9BNYlTFwya5x7vBTpk/SdURdEPH4v4Zv
aGQUIAQTbAnqs+hPgG75ft5DrhhbMBIZ+x41OBURTVKFvb/FiSMhXDRkMh4I+HBJPdct4J5cpUdz
7mUBoocvfM2xGPLh3N6s9HgGG1Df/0NBW9qyUdgWABBos7jqCJILOD7jrQPCJEnrTfgFhmde/5Id
LYZSpm2HmEuvKEQAPGNyq2BUDxNML1xKxh1rnHGcTOfJidTH8AS1XyQWgYlU3Jf+uUYzSRKfvgLt
Og32nEO9CgNZHsqFLLOLBFJnNpWkySdexE5ExtwJvKTD2l9qxIShPCeoCGw2LIQ29nGm+dQaQ645
4jWscxEj7AnN+NA4MiyuuQei15tgBjvyghp1HZyHcWwcsAkuzE5zHJOtkkN85/Idbv8XWJpA+qDS
Qgo/n8yNkysbC3lDSPq1nQbqYzXgczDTFJYmakLimG/3fI7Lpu1bzuBP2mKPKI1XodD+FPEr/5oK
RiyrCCmcqO1C++sXy1nNGxupwowRpSCLCAlechpO1jqWHXXYpSXBNRPKr1iKKpERzCYBLzj2Qzwp
7FS2tDFBCPHBayRyexYdIMlDSFkayIf9H/8K7uOVZZcxKBDxHTuuM4cbeM6YNwZ3cex/P5p1W20L
RcEl/IpsBpcuqxhHPbmGSQ6IthTO3i2pKxtv6citgy+a7ERS8BD74uNNV2q8LA/74sX3j5kOb7Fl
qF1yLtZTxr9UCVSbgC1Ej7JhZEVHZhz7UO6WRJGnNYMOQhCAfZrBLu/a1EuBxl/fu5VceEt0W+7l
DDrjE9ulTJgTnjjAT2wSFoNP0hkUTl+2QLixNF2jJSAvC9vxZmakrNsNiEj5DlgCD7vdxdXEhACh
h09ln7rNLGI0dUiBXMkE9XY9c6R/4O4FELFBAlxrhrqxBLZCpj4W0l67s38pDUf2YtkEhyXB+G/k
wG3cH86ieegePI0I/C2aKJ40wX/W/A1Nd2OQI07jnFOORbVSAbC9kvJVWuhDaxbvdqVnvUegfRwC
Z/QFRQTl0wAUhubLCLnxxMB20VCGiMIuK4WzM5dktvOcwP/TcDYVSvPkYB1q57fqbePrsUGpsI7O
fLn41/wHTZw8QO9YjSDXQR3nof2ef/mgpM8efPlkVZmeZr9ZHkFyoQMIYCcVK4ByX5cvZ5yypMmZ
/l5YRuf5pTC2zQJy0zdyX+3dj+68GdBCDMhP8I73DLxtDIKoprfsPRLNmCTwQhKXVdGcrbGBJshw
r9dHJV0sjhbBnLw5uHSjjOQn0KCp0Xo5oJCM1GRT3yaK6aB882kgoxwbt7hcUHAaILQ7HExj1bZu
axBOuUSx4+ExvY6Si7XUnQCQgg02G96ntq0cvtdJ6aY/CfstvtbYurhkRZnky76KdCIYwmeKjoyS
79OF255fo1tKemQVZ8Gh1w9H+CRHd9fQzY2i7zvgf3UsjS7GHo2xoOCWiFJ8nsmV6bgWgM6vk5Kg
FSWIqfY3Xhoq6b1sEujciCDs6+BkyEhtGmFfHsqrUXUzOrA8wT9QpMgAZxbnryMpLAH44CM+XD9h
69hIyOSvmFbc0ma3XmX/hdb73oWebefkqKxlwk+TZaajg2eb9TJgKpr/sLqiTbm32KZBACCA6Jp9
M03TZGlFSUJlNZpJvY6MVs10WbulQycXbayJ4kMF73zuNxzSI0opfB7wsJF69EaUtWcROXwoEaoj
+KlzBUinZsK+u36i8n1OdHFzjTlnrxX18bP7gijjBo+KNo8dn5jQri3bNMgF5mH1FoEK82QiodAW
DkSi3dGy6i+A9OQtee/pLqy4fkoUBztsNslGrSB/jNVEdoclrlD1fEhegy1+BdKtknuTcty22pOf
JrZrlXDhSyKLtPx1eFTR1877my1/+PUQew8CaB6dTlSMJBn7Bu/+eBDkGjqdaqsOXtY3wHhOWLCT
+M6ROabLd6t8M87J9sOOg/0vAWw8eRCiVYn3DTL0ALWN4MlpnW7VTEXu+0iib+NJzvefu1xlRoDz
ggXSiUPU8zuI2KsDgtBPheJGsL1CS1Gl1dztwY4wpS98PBv+frvBiq810iJz0nH4yAKXHyWTGQlQ
LnapXfSOz9OPwJSeuEtOFGdcizUEyW+emqMZFxzcSIBwXDfi82y5FrMaqbVn8HkuQDtT/f1sZHLJ
Z9rqTww74FKKJP6Yrva9/uCCSeFlKXRDmPIdzGcdwZgIFJczEMdGsZ/GRe03ildS0fRHSYuUdr1T
oCdHfVTjbRi4+hTg8SpLSTo/iyCLsa4dMQLyyHkUGF52w5plRAWOlFxP4xmPk0j2qdboWmriIJng
fgDES46g5wSJjz6btcuLGGcaCMeQWQc596mObPDT78Akw/eUhjtvDra2oqra69Y1JvyEg4Et/SOB
UpGqBMruJ0g2NC27aDu6GOTcn5uZaFMJUGGWyQAK6n7twcrd9IXOzXdURzQU/2kNxUB3typKQJd+
mLQtrh3G5XIzW2nJLmUwyAh0ZDcW4/0Po3uHXKjeW3Cn8ryYTUC/iYco4PEQD0jPqISH3o5kmCtB
d/rwBP0BC1dg38LiKskCs6QpTeVjoan7o4lH/zYi/qsAOAS3wLbrqD6pIrC5s5l0yIJwNiWeTqo5
yH8CQ3Op0o/yac/NMu02sC30AGRpoDuRjGGIu+oCb2MsTTMm3f0Zrit1KPYwiDtAEr9KiQQQUFrw
LFO1SdPrP2kXJsVnsMtJLvHEzWloMisVop7lozgO0MOy86b3SsgmeZAU92quvX/tPAAS6JVpmFaZ
qu13cpPrikbHbtLMsaamQuwAnnuZrqPn29tV6sYumPuZzTSgwitJR90Zk1SPnQoB12zH4vsRBV5s
Yn2Vl40F+aJAHw6Uu+Ul/RKZSchQHByAf5pWyr93Zhd8Iq4iVPJgaGCG1iVZsiw/A8cmLdRBwhrE
lX+jbfm9YbJsC70Y1C2JbvNS72ebje1CxwSZYYpE11TqejQKDsJVdRU9h+KgMN8YSSbUGZNiAGWa
lsW5/KYFPGx/NK/P67DsnX1qVKgMcedOD0PJh3P3Ny7DOtaEj3iG7y7+Axm5BVbtttIwkYGTZXq8
vdmuPd8+gSAVq+7dZDvSLWacVaSoNZaOKSeQOiyDg7IPy5RHilLV1tUxuFDkzqfRN4CBYXe5Edtj
tQJB96nZBAPivh640XS0Nq70mCU9TKQ0SRGpS/LPMb969C/eW0GvFkG+fwB0AE5bu60K2qUBYx1M
5W+CSWYyQR6KSMOttmXCmya/3pDE2P8TXll7mXEn4VRi4h4dG683/8fHvPE19Tg3Z+PWvKSqX6qe
mDtN3WpC7l7ymlrjgULqS9hkrxAPbQke++ZXJYP4OkoWMk4TCJaaQXVzdXJfz0Kejbg+dGLFZoS8
tf/zKNohT1cvcLpwVcmB3fraedMXpM4RTqg7OhwgKT5jyWH/pQCeolEOwrrLf3KQNFNBbJnBqVIX
uvvI8JC5NQYvuke0HF7ncMzm3Jm1oIgcF7dObW/FWNMsi+YpktA/+g3PQSHXymtwsH1lCpKtBTgg
ewC6OdEM3IjYIOY745JCsyLw+rXzjZQkY68QKJ7GWZleuUnYH5QmdSTcdrcwJ515cTiOrHWHkuN5
AWFHq0sIcIaqAOdv9FsA9ppLpIUZW7PPbZjB6v1Bvu1nlH+xhCt0F9sDmKDcXqDz5W34u1yrqOYn
ZShANFQoe0cGUaRmfCZIaI6bBZjTFIRzZTVgRBXnBVvQ6cCFaqmu/HkJsNDayqXp0KFVVQ7/5zCE
9Ted0qilM2J9PDFFZvel/tpPkzuaVjsbZsOVxF4/zBaTZOq+oYqa24jNaPfYf2iqxKuAbmNOFjuW
zKuM/Q+0feEiQU1VSEJE3jE3APO/r6lTxBBoyecfCwnxbUepqbRyzrSzvJyspythrtG898Qnkr+Q
u1UYGxb+Y7VeaZhx8utCOH3TX0ISyj3MYDBndaYYgIQEhOPKIwEaHHU8Iph8rCiNuXwo5bTI8WBb
OAWDVvpehCi4NPRdzn9jQPKu1WqqwMecfR2thEoVkHV/vt77Lmj4nXe5zEuBgsW55cBW1njELxQ7
rcjxpLdUsP+8zJIWxNuQZJNiuFu1Dy5WTWEX6+YEXamGL71R76nNRzZ3fe+RJpdcYvjx/BLqfTJ6
qQ4y1xSQQAjxin/z2Q9K9liBIqFJTg9gRnzR21GHE9mfDoXBZc4vk/i+nUz39QSiS+NbFtTEsRBk
mzIfo8d5hUC4uG1WxUdc+MicF3aq/zid+o3ZU3FfBVUEE/lE4pLZYOOWwoJwe33UOGd/9EtIGR2N
t1yXDlno68sPyE+AK8K1L0usJm1wrmGuKNigrHj3nj8E2QC9bbW5Xi7F0stx205SDOdvAqVIb/hn
z4tvPdqCHSX48q6o6dVoZFuUfth+01lF7YeFxYRodXFLEnA4nazCwZoGISxOqRjteL5qe07fL3b4
RysndyrIc9ZUbA66C7pCk5DaXht0q9u+sOlBy2xCRetd4pUFyJKEedOxMetfKN9T0rbk7VNHfJQ4
Uw/VBuY2+qRxqATJKBaPv2JNU+OCJnMcNxQw9kvWB2XMxlulH4DLztG/fLIe8ghweqXQlKcY30pW
2DuN4YrVfD38MESM7lZo6finaJ6FmAeuTbHmT4ZoXVIpJxhCEMGFAV1FHKcyEpHViFtMWdzx5k7b
l3d1WnTgXtXzutbj0mR+F4RtdtJApmF5aTRNSPlTIaSF4BS2gKB0tEaKU1lASSikFTteaL6MwBYR
7Kf2AI0MOXzbTxb2WWXYyLqlr0ZfB5B5oKyG2MDN+5udbc6uU31p6RYvSyqgst3Xe+UNMIom9njD
QTDROHYIz7G4fDfh1WTlQGafZzF5srEkhXcbR+TxR57FZYxswnS6nzvmpch2lqNx93ElyczfJE7Z
R9gkTQOSLN0kjFRXx0G9wL7nB/Lttmoh8YpcxGydOwHMW+4Iza6KMP/M7IwXhUdLDXc3da3DLrPZ
Vn9NQO6EMJa6uGWB6mgr1kNSMAbh5uSHgAqQqZrcUU3Owf6a3IHQtPV9rBFjEEIn2AcRJhze8FN/
/aEynF3oJexwuk4rCWqQzi3npwdBSNMQ5Vi11Nn/D4GKM7dSccEmIJJ51Amh9//GOYV6x3wrrgax
DemPSrUnNq9YGJYX8dFh4Hao3ROVDd/1gJYeYu3yD9WzAH1jiYkiYKs5lu2+SHn9v3vsRPAAcIzX
CKeVwy4GmoI4qcEwYMhdsORAVg0B5yFomlSxw2/yVDZ3jNYJ7REqNclB+8gbHEz57gfrRX+hH3ZB
Q29QgOXnE6sZzBCfkFNoEoKqK0IvmVu3V7kCW8CEBlg9YYYb8YwTf2mkQNpYuP85XZhP4/xUCjvM
XEW7wO77uPLmQHdircpMXD9x2CtRs8E9w2L363Cch7ToK2s1ddzKhfL3Aop8WkbCefokAj2vf+pr
j0IkCb4R9VUBZCndkhkUXNDnDPuRwHnz2hDzu0i3qDvUMRwfVaETg9n1tGHgIjm24uHGTL22qQmu
41tFqsJ2ZKaEa2dod8vzP1gL9K/wNKcH18DrQWIFvCR8dVDScyRivVseohBVSIMj6UU04qbNLkH5
Wp7X0um2Vg1HV+2UvtA1JSLs7VYfP8oAWJB2opLqkxmdaYtXRRtJnMygdYPgV/4w27WHfXboWAaq
UzFu9yQX84HR7ppe3XU2d1qNY4tr+75GP/JJBLK5W9aC7Xvl7o4YVjNE7+HZnSqvVKy1J6C3azQ4
l1x3WSDEYKd57ryp+BX9shyl6Vxs4d2QJ7qZFRBlaLYsZ+SkoAVbgNnEoNiIbNvGnRj1gLV9d0py
HJwGYsB6IMkLRsuF+Rt6uLPaGRWbm7uizpAn8wzKoB2ugb1qeZRcAeuPikxJYKFjzC6meGIh3ltz
sE2b7EbIZcAXlsvWbTQiE8wsTA5H7CDz78gYFMAOluTEoOa/DwhrwHlPChZ898fgkfqqUqL99H/O
Ew1A4/psI4FR42F0TDrdhC7KmhGsyYuwzh6RgjlP4O8iED2w9VDKrWkyZD0ghpQEoBNjpNDcRlLy
O58Yn2PNFpfajHebHWjAUxNUFGPMhQBuEZqonhZ/36fZZxnhQX1kXqBm+FiJkeBeIbeVrz473lRj
nQQPZNDVdqISRtHi/R34GO7IYtVaX6OwH+Dg4mcTyKUh1DjqQGzYfUbcoYv/tUtmhAzp1zC2CHYc
Y4umlU25soY3ENV3F4UoVX+ElkZFzobp2XmfsEVx9UmugAsovxq1vo7+9WjuNf9vs+khMvMwxLYa
ig2yX824/yrMC1J8DVLx/W3eDcSJu+Naw16UBag6ctNuLxbvp6HygrFZtypx3GF6D1d5swOjYJyh
K5qP/FFYAspuDIH2eRqlHEADlIk7sRBjHR27+kOeTboXf4yHE/8Cj5Z0dId3eIPOcffTRAB+JkwC
hHW6KNzWPRgsYdVNJVeXUrQHC1Evs8JAoYlxBvP/bMPLvpOJxsNEXGiBtHiW++reiFXf26aBzGrs
UI7YHXdMRGlg84vSxYr9BfZajNAfnOo47raPCLVHv/0MEk6UlikPtwXLVzNRhn1VxtKgOSgLwISg
tk+N+E6e1nRG/GmIuNGWsDLUEIG2kYHgbCzs6ycEvBXmbz0EHmn4Hn1GBuewFZo1yNONnIy2Pq/q
fDkwjTYfv+xK/ZH70oim3UiMW9G6Qz6qhr6Wq+FqjeKTJXeq+e8fY3KpItufbH0L6juNQR+DzQTF
MIKtx0hG+5ZAjkEgIh33l0WybBBZI74MmQnNzCSKJ2TcY4WQInAe+WMmrZ++1Iasmj2vRXkVg4h8
0LXtIzV8kO2f6px+Xrod67juB8cEvfFjU+ikXkFHsxldmyTBAFzb1uwL9U1cEnuQHEEsohBMfh4H
xfs1zlJwqTDYvHnT6dSGA+KE5yMaSb+tGMLdtUuiKfaKwH7Ucsz9BKFk1p+ZpI9XXGqkccKJJVOI
L8vjbBMQgNqt4e6TGNK2Hsahhj1ElcAeoYFzwTVp9kpx6k0ZTis46SsD0ii2xfOZWLwlQ2IiAvlb
7wuiP1ZD+8d9CGeGsMg8uet/jpHgrYQG9TW/h1dR3nK6/EoZOL+Cww2BO2nsuFedI5PXZUciS1LI
aRsdCxQzJZ/XvDPtCbJvCwLrEaOEObnM2ZFi8z4RhG8iJoEOtEwF/s9clzvQ/FiJgOq2g8FBxqZn
CgxIgxRpjFCjbJmaSgLsWC2UXFl+rOlw+M6qkDxsa2CDcT1Lq6bhsbxslOtVCEfRdAlwdVqBSgw7
SFyguMundvitZG+ZBC0Abnd2VHE6v/WHtnMmiS8FeqkWsYcCPLwf9RLNFmSmvNJ5MDYjyrMtWWMU
/9wigkB1eJg9k0pGrDif7jVv3gBORXbE/dIWxWC9y+8Kdms1YLFCGy4RLj9GdXH/sY9XfPs64Ibd
lYkEHhAnUN+JgVFk12Nc0hdIiV2Rms7q6uV/ljn13CKD5Z3Aa4WccNdA+kvGP//vivSEHQ8j/9hG
db05MgfXZlQZOO7pY6DCK2P9ctjsrKK8QHyveZ7MtGRZaAu4Bz/Jz5CuzdsgwPFxVQtPqiTLd0VG
tQFOwxNl5BWPcUIpC6jSA9hHXjLL7IbEG2ICeLeKPRSngFEzm0S0HIe2Vcw+m8XsEcVsPcoiGsDM
wXKVn1nRNtJmX9lUsS+8CwKNMwtVfW3R9XzxZ54q67flY0ghjAV+gnwqgBUCLykSCqct4kRAWVgF
rEIZCKl162GupFyY8eAn5frmXI/POJvhX5d/QYBwHgh2QEvZrchC93FNn8SNVSBM2yshn652cvsM
cnUR6XT4LmxVNvBzgVY4iLyfW6iZyiQiP5YlR7cjPGJyzIpqNOxVBUh96sqWqSRrlnuU4rGaWeap
5EZl8f7uBue7F2pqaScMLbiLgC1UDRX8B3qWBifyiAYfEQeBBpkKQMTuOpmrc8ua9yBxAjZFEY3B
wySSNVMXen9SqvHnUq50m7cz7uftDEWY9QpupO13hL/WRpjy8wtQ26stcB+liE3kMy2vVyO9HLDC
WjLJlXnpAaHCDjAABRVzBa8bjTvDT3yxu0X1caefOaCcD5k5smhCF350JWQJTJmIDwjHFLZAbUjP
W6uyfNoOi8KjlZ0taeOEkovR5n9VzNX5qNkrw4YCb7MkmhmuDUl9WYLF9fuL97hA3ZYstNz9GdrI
hyXTMeEi3OeSIePsQf2Wfqx9f+Ida9F0yhrm0Y+TcAPwz4Yjf87sOTakzSQhm1sQMqPvV12u4ndl
TIXqYvfC5527FAl40wfzdA0ZHfKLA6c7b8jnqHQ7l79ZX+RabqqCA7eOGrMPRVf0JEqvo7U7ZOqk
vkmL9cMYEVKKxNiP/GoqN6GKUgZ3w8uoME+GolwN/pJ0MPekNeBzQFYS0xqG78z8HT0eHTVf2bUW
18g69VjaUxeGWfX4bQqkMcGZHIfE1K2eVHWv+wIJX7lTIStXl9cNLJW4nF5wZOp9p67kUBCkSt5h
JnVysWS3OO/uM3RmTf1FL/FkUfuYJawrGCb9yEXig1ZayFbyccNpq7/Gzu3IoCrLQcwVUHeVIIbG
xg9PQlYo3kSSneVlRXKwPXFJ6xXkhFZOhgKe8Ew1EUg03ZGvtyvPzN12481LrqJHkGFgCQdclfwV
sDAmyJxH8dtuxwzgJqZG+dMe8MtKmWP/xrkMiWW2thjRFUARUs/rR6qEcrAc+PDeddvORrQQAx0J
3cAoJ2fXGs7m5iNJX8+TVf6eUm9rTRmlhI2ZZh+oIpWC8H2oHjRfTXyDnmO4YLDnPhO5jFsBqp5i
dvHED7WUWgpLvvLaJ9jYoz1nafgU/z7ZKpLU8/jScb6d0Btr/2RRO0gG9n30kXzlLnFa2sGMIdsE
C53mKHj8IsTLuMET/Vmxo2IwHR/ruDN259we4qw7OqkZHAr4BtTQ0lHmJYweaQdSwshj8NrQ7NHP
YjCnMQYbp6BsxMHEQ7pvXunEsRJQ684PhXE4SzeXWI+omRTGNgdUz51r16vkNYi92ogrnGDpd58n
WetszZnrUvMeyQNu64WeoajtwctQRPCXVRuni4BSBjuoya9Gk8p968RN8eiqKrn1OQILwpGfhur4
8NMMhB0d3tn7b4i50ydJioRO85wPSvjpRWB4VdwG6A9aNqOXbiSNu20JylWwfxz9HOaW2fgg6aGN
2DkGwQU7t+LUaOArbIG2FUrunMCflpApxXHVmqpHvNp/LyCRvEYmU3psMIwtxCnnNYD8IktEoj00
CWPMbDgwYl9fO+kOXEnMjrK8P5jSq2lcRNFKbhUyIjr2wcv7ueIKRLQkKJO9hbCIl9cleg86cKgi
SVUyoyC4X+xncQ6LHhbEvpUAnxHKr47mPggbGebx3morxfXrAYpz2fO1xaD+DmqxwmF6Gs542NVO
KhvUKMlBvkwY9Z/NaNwTB8QdPQQdBLxHx1lT0iO3Qm5wxUdM+oKNxrXuYehwYK1ZSjC+0dQ7ETM3
DjxcNciiK4fFtay8n3g9Z5yJL0YANUrNqRQ5KFBBqWafdtOx+JyGb03Z3XwdXIRfexcpTk0ucvU+
77YpulrFGeTCeVhrc5Re5eIZhLGLmAMxUM1we4B4rwUckFtcJmtuNbfCgpST/bt8ezz+jejU1ifE
IXiV3Khi4NHDIjw5aUz4KGz2zcEAfvReVEg9YhA02iSQB6X3irkPw251dx/b4YYOd+GMNd0aad9Y
cvX6vQBpabiuovvVZZdEb0m8gYk21pZ3CVrps0hD2ad0Kd9w+YFQPbjcxhCkjNNfqHFcgwOh+nwv
XoycZd7o2/1snCHXcY+EIQbVCAJfpOq8xvgcg4J/L/b4zVjazfnagvKl3ik6mu65E6KYykPr3MdY
MX2QGbUxIWuI0LuQlFyIJJ1+ydGDlMvKMArUMaGwdUAF3m9UCHfztYAfKC7tCkCQ23kaEKrCLF9C
ZtlkrUvJkAfK8raey1zzqYBJ4+XnY6DssqV+UKJbhkfm2RFVLp43zgONxqpUYr4/d9lb98RqInlN
GACnWFYMSTTWe2z0Enlf2UpJncbabpTUo8MrO83yh74LTlsvXtd9y5JqZG82/or4YAasHTnKccoI
tmFqbrQV2bH0dDZWUjJrs1Ks6DXBprQ3yuGdQLIdwpBy38iPyh8nmoi/UrC2sZuF3IhkF9QrudN4
sAofC3d6CQPe7z3tZZg4gw5ohBEOUuviWLPaBiw1iH+GpjNdvrEu+AER9X/WdCFtRmTXs+S/T3N4
NlpVVUkHG5j+B/svGI8PuUdFjCBbtMKDkbtdC+sIEayujCxz/Gsns3zaZeog0NewAocg5dz+3zKi
lT/xy0ZK2uRpDRfy237hWI4FT/LLagDNwaduDPTMmjIV6ab26tMNYjEFrk1Arj2ye/wSokWFpcnT
iK8yhjpPBH/MKvxp7tepMXQFZzlsue03TRPfA1+AZd6f3F50bmzKAnwR0AcB5FZSPsgJ23vPvgGO
88/JvBM/CIoyXUSztOBQksLvY0jde8RMJmCtg1SNvQU/PAhYI3vovm+ZYRn5ZkUMIrAPRbcltINz
t7QoQIl6BWf+ewbwlMwwjU9hYe8N5Ps/4x3q/+mYbqnoVJM69AgpyO+/XAiy92gPngfbdkDM2HNr
eo4veqoTXZN/CfkXf+ZL+QVnylTHapy5/rMHzQtZAZ5+Df7jkl0kFfO2N2V8LvvvetIh1zKMQav0
VEbQbg/fzFIbUK9zceJE5xHfzHnrlHevK6qRP3UJsbgeOCwM4OCpQDF9OWHRnW9ICODxzEh/tRd4
SX8qlcUDaNDNzwP/mlX0FHBVCWu+v4XhQuveg6J+cdhUGwkxH68EF87JfYy3531uSDpOfYcqcuMW
261DhuSc5fMWBAc68QRJIAmW+68Qlk/gKH6fuPpSad8LrAfe3Ri6bEMk/hvbfPQZaSKBQPo8tjdh
g0PnCTIlovlyOrp+lOIOuelziA+yNBsrvVPsnihQ5TdWLqtuASYxFUNv2xjnqHxYzj/DFc9ggxUJ
A/a4HsjH5Lsb2LlZJEppHRi/GwyumlhPLF5JBqdoCLN18d1pSO2VFVL6TYuMkrEg2krCM0QibO1+
K2ClvcbH4qYZJBodV16oDiza7w5dndyFwaAIlUnCxWct8LSxOY0xHrThYo8+QYICT+QVEILauJek
Ib2N7LbBNzWp66Ru91FM9Qk+3dCtTYbDAULdvIjXl9ezFN7fc3M9oHC0OsZ/t7Lx6aFXk2UgGivT
do0egW1ceqWOQ0py8cpvPGoDT1z/+Ym8Ze9jT+trAd3SE65xYzbG2nVfFCM9urIaP4N1o115Iylw
t/TbZOF2uDomrbf3Z60etrh5h5AzeGc0AWQDHUcoKoj6tEwlt2DRxUXQU5iSnLWl2cs8TFnNPD33
DapgAyIVkSFwDO9Cc9ZGazXR1S9NiFfRtsKSGNVGDkhBgL/vZHJWxrF+Edm1M20Jeo0NB38XrENZ
VJSZ/eFNIH/w9doDCBwpMy19j7n+RB4ZRP6+hXXkFTPmUHoT6EmIhNrnjqAlHSe1jS932qjzpXBe
gy9d3Mni5aEohYj0UAwf0N3jtb7lGUf/M+fEuJHGpRO8FNEriTeFfG4bKwXXoRlXAgU/JPdOZ64K
Jd/iGWCt4D8sW9lYf5e9cl7REiCjDM+OtPGKb0QM2KAy1h0m6lm2SO7guloJuRJU1tlLAkwbFl8/
295/uN5Lowaj5gHMrw16jA+8pgcEXhE8bx3ABlcxYwJ64F/5lAQA80RIR4ykq9jTwNnhgmlhtjqK
V+6Y5aHfCuH+Xj4xI5o3UHYKAXh9jnkbhPVYP3XwwLO8BW2Ybt+j8kqr2qiRkq6hwGXaOuQjW5xq
yn8OQ4u/j6Tn1Oj2mABj6qDyAz3p6Qbl6rj8VUHZ9vW3Gx6Pvungt2iwfdWaAwTgsAg5zl8M74Io
t95D057UOd5IoqAADwdnI0ms3TdDaMRU3ZYObDyASlZzlU+7wp9hlcNEIBfq58WHZ9WHzBbpjj3g
gED0Hv/Xm1WU9kSKeyVFyLAuh4mvLP9sJM0OQk9Tq8fRTtp3BcRUl03TRQcJg0mq0botAcM9WfzY
ddt0PJzCLNseLlvE6mlYmjWe1eJKh5P/6fdaG7e48jJYUmmUkSl7OfsAmNMstI1PEAiTKAo4+c8R
YKGXn8hw4IOS/gGok/+FvdWTDv8oYgs00kHnmAIpkUK6ooC+cTNnhXsGXePQ8t46E/PWZmpMnBZ3
MbJoI7LTYV4b9NV+FK0K66impf7Q0hzFPq1HAXmXz8LKAZbZohdVCJ9okzrBhLJL6VcRdhcYhtuV
8uDsjOFLTMsGYRsj51UcEOorBEOY2uml1qvSE6hBcST3oiFmY3zj9x14QHEQBkC0kS+pDB3D04cW
aKQ4fC2DmKiI6YGYkU7lShPBT2WFyuPqaliBhaV9Mg029JcSgxuBhN+DZ9eR4QCmkou/bcDdeb3H
ctXW4UPT4xWleIHuBMNSUjyGYh7WwQhnZ5a6/upaesKjR43PiDOO05wToot0jjLrHvIwOBQJtNei
jvHL3OLUpE9gyfGYSRW/6IWQv1mmBl9mgxFPQ+QPPmyrgQnztyd2o/rpqmFeHa5pZUVI4IFzkXu0
V2ikY6NYZ1Eynsui/MWG+OdzG1yQ+EzJ5T0ZVbJI69YHPdWhGPwR+8XkI96ypKM2aVDp31+HZ3Aw
+WMtvw7CvsmPAkwCwz26sYKwGlkDPZ5pz91b8pvLxXcoaAnYdxYIDUvEE02ic9qg/zU/vSIHddKF
l1k1KeBPOKtqe9VUkNA1+pmOYrGCDxi0lBy3VC0qmKfiJi+D87sNj/WqJoRUA33Q4D5UDjN9Uxls
9q23tkPOdIcsZO7PPjqF5HQdZrGZeQFcIsnrX1NbxZQPi5s1tf4xnmgv2s1N29HJf9OCexhxqULA
B4DErHsEte2isd2YrC3XtWKKLhyDFAIWUyX0k0Em7J2+6GeKuAIKyrxoXc8zRtCdFh3hk6SKumJA
y6GyL+kHWuZwHRptU3xcSVSf3syhDZ0MVGd+eM3+blh+HDOrDgJY5gpcFbbC0qO/jKr0oxDh2XB2
CbpkC9L3k5z+r9K/Ch+GAoDckl7TElmvg4GqrTN914qvtIG8Ikaq5QWD8TVH/xmR5pB5g1GUYVxr
IpzvtoOxaJYgSmN58TJpqKUR2O6bmHwz61wGiK74d0RzOa5m3dbimbOh/UrMeqrFV5gGKfthYFr1
vhEFDy+ifWaIh5pA6dy6V40A2cqVIS4zQd1NCrVrTmeg9A7qfTCv/KAiWddobhfWMl2D93N+48cV
3VfvGw+ait/MH6GTWebBD9Eg43nyiVSssTbg/tMKuZFtMOwFojyk+G3NrMlXnyqa9Cz4jWzlJKIl
yVZJDJ7gqaASiAsfFPs/LTIq/VFlwvYuP2qODk0vOOoj8eoPzA1DeU0ikjP2SkbePUTJm8wBtuqg
Y9kDWpwfLfgot2oMXTbTyX3BwAnYZ/K2oGILbAvl4HRCu6VjzZM8RURysJ1wzjGyvyYpXaLdnjmn
wORZa1G0RW1ZvhEEUk3emIDYPc8XRirBOn57vhxPop1V2tjel1vNHUOnSWbPUidgA7ulVNWTpuJ3
q3bn6wInVJRs1alqRut/rwA6d2Nua8qM3BeHygIlMgNBWkTMBnfhZyG1WBYlp3+v1KsEj5J9CWTO
W71buiut94e4P5pM2uy8OyPBHHoZR1Rzeqsv8NPpMXQLgqb8+z14Y9EwO4VAeTRq6TS74KmyA9X3
uFHuu55uSpbvUZmP1OqKm8V9VhzXHbzZTuTh0NSu4tpLWtd56Twf9KyatvOlFICp8WGEi8oEKmlI
6PlcqGJRv6ag0XLrJb4orE023FQ4A2ktiSTjRL0KRGL5EVHWd6o7yoBTaSy+T/uR1SBMY7Xnc8Zh
LD7fM0MuAztsd0UHdWjqSjkF4vsH3yePtS5Uze+UeZorepKQGp/+B5TH4OYOfVSj6FOb18YbdI+t
V+nHV8OzROg6M04I8LLYf+9cBcAsP1mG9ZYFVWIrRfwZTmVdmdTHIdV4GJpaDdT+Xc8t6lAnokvk
0WpgaReqzFogjpj0rgyHk5UOiAgdE2tumBz4HKfbTlcbvshEvHOPxVbsQJPP4MnRrfTfANUMcyqO
3BMRQqWE6+ruYA9TbA5PI7I2RGPo78Vit9N4vNHeGNBDpRsmUHr8K+utrJ//ZDNhPjH08oZh42Nu
9FtU4RV14UHPyeUO1Xmu20NN4BW8aoNEIm5lpkl4ZPrKFRZZ5XUbtM5Yt/d34Zt8WU+8wRCb/P9H
jhQAGitMEnuJD15iZEbWLILGTik9fg+JY8a69/9eTzKMaiWfIwjVCNW4nR5jFgTbawJQIEKoo+Cr
Jh06R6+J8nNv4R2wFFHhkUwAA0tOOSFE/BaMd1DlERj3JDneckImcVsVVS0zid/TWe3EDXHULu8X
Y91biopG8gu8/vIjbznj8NIN5DYNN60QHzl85xhnq/xxgo6jeFcZvzw/oGwN3GDcgBEpnSnYpKkL
bq7B17r+T6+UoHLLO0Px8vw5X6I45k6209lF9wRfof5tCxpqEtPEiCwhmE5XzZBA6Wr/vF9Ke+ch
kQJPQv2t9zCn9tIFYSi7N7wAV+o4lYLjrw9RBrxVQWDbO+4qCxHW+o5U81eKO+Jzmu7TwIpHrVTt
QBpTj5KYTh1+HHlKP5FZMp4XCj1DKdhyRRqJxhoU7nNdh2s/Okb55p784YvQCT5xKcxbQP+sv0wz
NnLoIBkd3SmlMs8lV6/l0DtSHQ0brs+AeiUikihXIV0JskVwrf1ltGkcp3wIzZmwQR4r1SMTSRED
H2GsmB8s+bCc0NEjLIjFS68C0gmVnGgI6QYg9GRzlJIdUdzX1LtjcPRhUcPNeHrMXVQIidYQ4VLz
ODqL6illb+QABcELaFCq9AYvcMT0vmZwgXLGgIK08AtmeBk3nVOyEDzonQxOTNSQfCz1keJauph5
DT4kF0IMeJ+SAD7Kea3FS1do0sTF/F1RYBrffwGrYzNOwhgGwz1rHN8CmV36igzIk8DZ5LdlYkC1
dmCYjFK45DXsSxkdgrm8+AE0FtzkYNp0z+9+5XmNzO3c9Ovw4HkdwktidX3AiCSitxeDYXWW9T+k
mSuso7T3zbJ3R7lQ7CuLSIsdXIXi4XUCqZFUO9Df7OAzYFOxFNgFTGpX4Jf/RXO6Ifr3HirgvB8f
Ey4FXYAen1W6Ny/nggq9UAmAQjwrPFhqE7P+j4/HkDAViOZA02LkYHlKekmUjOHw5nT+y1RcC2Lz
c3Y8rWwhP1uOBwl6faie0DSKcVNRGmkADKaO+rd6IE9p2U1hOiCMzTn5sv1MkTh2L09rIk10mkYp
SR9liRAj9A49xVM6J8CvLnE+O3t2vdHls0VsMifC+ETIZ/RNo1+1GSa/nj4gbhxFEAveEnXWX0/j
sbNgxk+rpX1o3T0PQqirC/geyGP0uF2fc4fm+G9QAcJU2ULKP7pwTpjXU3JZ7E7khFjx7kWhF6T7
mzZMyD0D5V9o/IpGnBSOXg281ke3fII+p9YWbMMQKlpuIPLiwXnQ424sJzMGJm5QOk8FdXmxFOIs
9KZEwaSF5mQqnj2D9kmR8eBDO81o23tyAfiBHbZ2y+DlCzJMEI42rabC/UVOVFRhs9+RmrZkO0pz
WPpO/IPt2FF25QdMFkDrWL6X3dfTGnJRwgB/2I6RCOuFNQgfewnGsq5BmrjVW09TkIRrDOcbBW0o
MRcNaPM53xuvVXsoNYEBPa4/gg7TIczAmSHptW5fJM9nQWT7oCJjaraVIkp63bzE5xWTs5uEXyxD
aBAoowJrwpG1B8jcNy1gjLqdg10PT0aGYRICF8HB6hYFe5zqwPrEdXiIYjZYbchaOsNfxZY99ME5
AnFwIKAxmNnN+nboP4V2zNvoZ3q8f0VVu6e3Rx9dm0RiZq7HYAvu3aXOy6+WG3xOf2bdKvkUNEwq
Kbnca9TEXBK6khBQ1KTXObObCBKAgKzO7kqbfYJnSudXzlowkEUWobSNoeDRjGcRgJszDdUBJRA/
mTahKSpS/ZdJgJalTCeTYW62QgMAhHqVzsXm/nmZTsow1Bxc5+GRfhPDULNckc3mKs+ijVvzggxN
riWICFfRP0lVuWpxbJr1yP5d148ryN6/o5Wib41IGAusUQvafb1eixNJupLuYOvCJ6vMUddfDaBr
T8pil2yFpXykp4phyN8fika+sMEq59YzNVMD
`protect end_protected

