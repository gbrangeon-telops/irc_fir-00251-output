

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HpfjZK6WG7sYhkvMgAngy3z+9zzwD77820wau9oTTb6dakSkVNELcmI1vCDbEcS/48D2LFxL/qT8
BNFOIZ2d3w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VPnG2AZhAX4ivH+F+USmM4TuIe2lYrNUq3Xx5puxPaV5guza4OeVGJP6pYRxsBYzj3S4OGH7b6n8
K0l2LCX8eil1TGx7VbJh+Wd7uUD2r86y3rluWkRdWUlHXjFOxoCZGO3zP09eR4IRsG+JxbSDSiqj
FoMAGfR2zks5CEu7dtk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1IQ6dlJ53C6R12Hzl/XoBaoEA3n6gOO0fxU9jZJvCev68EW7XPnj0pNHAKpShucryAUuc2FQgbE
BwIwQ+0yjh3dOW/yrG6sHXOI8NvAIzuE1LMkRT00JCNCjyt9JL0PrhVhWC3cY50b1mAkSZBVfMWL
G4c5aMtB6wF50NpvOm20Ptquu8OAMlN0E+mHAN8qvWTR+CwIDUV/kvH/83yRaRonCOBULUP7XzwI
uAjFnciSf/F9eC2blbPxLHlWXLQDQaZnUw7NGNc2Ufyh7lsh0GoZzefU/JIhthv3ktn09r568XNe
kk/w7iRo/w4FLMicA3dbzrMyZkiVt8z4I74KAw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
x5ctSMYno/7jD9HwXtHguBvqXjqGDToxuRubQZySJLeTm3iuHlQTdlRRlvw3jNvFx8WWN4nEmWap
sLwuJFUESklgDZc8wPsu9plvibxKvIUprit+FQWsTY564IYlM9a003tG4rrtM7zZ9yfolbWe2MY7
qJFpoVf6XAxMMDrPtP0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JhbANRgOr9SOBKZDRGJGrZPWNKSEG3awknWUR+2QiYueCqJ0p8+Oq42E9W+XtOMQqS7h6dt4lJzf
s2rJvfuxWWYMk0rVRoGeqNzUfiVHbjHTaPdjhGKzIm4Kgu/QJ5ooRwBflBurdW1+74PtPtKpfjcs
79ijwPcRU18IbRTlWf2wzAlLDLkDUewye6if9pFfqGP8EVIxQIb2A7LmwWnM+VpfHc6KRQhcdZbj
LsxdBzKwdjN9Cdt40472gpQEnBtaoqRMW+4LW5rSmhm7vTXSum0cU3Afl+AWq9hUcVWPcrWeYdm+
aNrNDk+A5wRHt64iDTF82GsVuvkYpCi38y+ffQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12144)
`protect data_block
JQGM+dJHYw5FWO7+JjvhcEqafCFIjR7bTZLQBRiXHdF6LveaJ9h7ONpf0svbOObpYjoSvK9EzoLu
wz3HJtnrdAK8t9kkONRnfOP6QNBJJTsqqeG17iLTs6bJP//hBCbfRVRT8m/U8adS7Wr8KqSfFrxb
g8Aj94H4AzB2ywGFx+Hqou2sNwZ41yfJAcN1d3MqhTZOM5p6oY+OG/X000R4DYKc+AoJ5R0g98Kl
qTx3EJcvHL6NRMiakiy8MIXR64kd18G8r0+so5hDO/GJYv165YCt4YBWAdJ6E/ExrRQHuO4uXZUk
w/majJNQSa6+PgNldR6ZUfaDNttnnLC8SN15tUv/dNnxnYuUz/d/m+Bi7dZrpUYKcmSxu123dxI2
E2NmR2cALsRFoyCdQBFnoBcy0veOIlKuhhno/qdpUhDzx679AtiP1IDFnxqeJk7jUpLKoYYfp7sF
0zo4IhUiF2OfwoI7DsebaNfcCJxxOPHcG0m5ibZR5bxBv4b/xPYmMEfa7HcCv5MwnC2PaSQhm+TH
J/GJvK3bRThYnfYeEbjNOGqujWr9RYMDWob1vtJ0rnJSdTzr1mHdzAKtf8juJBHTV0oNVUYVYlBM
dnvPDf6cgaxhHRrUYNUYP4c70+GRdafImvPSFVHZkzTuLK2gAAjpLTmfR79iSIp03zni1StlMvek
dGW+OoYlod2jJN+RCT8Zi/Ol7+ToTcnKnTJIxFBmjcift0QVrO6zudFuijY7fbMWppWhSZFTW8ER
qcHB5utKWSmGgiMnJ6f9DEddMDNK0rs6GhTkF+1E1WUHZ5L2xuNaVtc1qfBvVVgkj15NHdGnwnmP
FxeuQLVeVDGNW59Cjex7xrYLv5sWkASmssgwd3ahzz6oZaW7H9bdhjs/dyZx5CNIqvdeaF1W/nzI
ebx3NM7RbwWDHiQOa1utY54hSQClEF8HnBmS+9tDF9hlP/4ovsxPe6jZzSdzLePlgdDVmxR8QhbA
yhd9FuxQ+7RSlwlezvuB5GjRlV/tzCrOURSCblF08lZKpSRRbeZJq2pDi6GELelMn8xvvYA7P+Ks
raVppWUNepiyKNOhOYVjaTs09C04SSCXMQ8aECuWXGhlA2Dy8CtF3jqiSYVVFDrigc/zzGPXO+Rl
S4NnmDIHUzmbNTxjulfc/CdlXTp1QTKb03BGi78tYuYPFMQ0MRasBTAIK6SeAUguYQ9oowk1MagP
YL2HzQ2MCnGtmPMPiLiKacTnKfOnhjQacIcketpYAeFwejiXvTb9AHRqhznml8MLyIicEEK5uA4O
JMzp/BveajYmZ+QakbNrh43GXZipgS24NtSBvngFpCGhWLTb6rlAX8rbkfbbwTThj0wZV2eOPSfq
SjVu/AFlfaror5ofTJ43uyvQphkn/Ybb/z0O9Ri5XDB3KTJfH6FcL4LEg7FQeb0wzrUOhTcM0T4+
4PMT0ENgpm+fE3s0Xr+tvtRa/VGjM9wFn/ySnYy9AdYo8WGsSxaWiPwURAhGrJP+5xqlj+0UIvD3
FXek7M+x3a3Sx4C4PLgRqL0JSBHGJ4KNdSueCCLIu7s7EQRpd9KXl5pTZU3Nx8ImIumq7KjLWJYq
iFkNlcR/yq332vgQh8Om0vMWmyxG9KYx6SHf1bs/k1MErKfifvCHZW137m2jZ9ueFgJWqshn05GY
yJfU6xlLe8w5wfArNCJFzwhWKUwsL5vBEYy8J1h6agHEturG9nRSeefw+4baI+etbefHbf0BtRKy
GrBpJDWVwGLtEMw0TMJGLG7ECXFHWtpF9BjO53UXef0N2dvh4hkoP+xXc9TXFkvYPoennyqXjzR9
5PuE/AQDN3riL1mXyeK7Z1DoziDL5WfocLDRrAxGZtkXupnfVkmWL5QuSlWFjTjjVYTZCSBL9CEE
J9oR8Rx9DbDAQYq8+Sc/vTOPOxmBAN+8OVSpR/D0cTW1JcfdWDfgWERF59Gq0WFm1CVDUTd7guay
bl0AWdyV8CGjhdP0K1/xZGPcKKkE6qqtitObjODLi9OPaVheWdj8lorVx4QvFegKfwxbE5bS64xH
c5DXuQcblJm9ChNmQORjdzPrev8dYKduHXYoyg0jdTnFOEDHE+nBJXq3wCZedv4BYirUAazdkctk
GEaWo1v7eC0Qh55nERSRAMy07sKZC3iqeg80zl4D8XXvMu2EKOJvpNNEAo6imMiqlvIpUGjn8rzL
a+PFc64tCZRoEpwxIRtSGRmN422zTkhKmQ1JjLNLly0vFwGzyH3qVjtVA85Uu7xXZooGyy9xWDbb
vog3ZPgONUhn2NAvoFKuNREV9A9ksRJd2SH0FsSw+oZ/TGA/hhggZ+KSHIacbejZqMdnw/P5Qd5N
8Bp/0nfxby5grGjwG6a9W8z5FwaKu3xIeOQasXrS4WF5cTya8bGSiw3jXG9/q+bpDAKISfQ12gnk
J8JKLzR3KrPmFANzUxXQjmoXyBuK2VFqmDlaqg4TNWf24LNwE4e7+ga+TVK8Ocq1E3vBrNAfODT6
okmDR4rCB7jeR5FFSdV5cJ/HLtZFYwGHndPJm5BfbvEpVLhdbaZSAcwZRUsM+oFbJopJUT7+tPxb
qCePL6hpOAsaHh+SJ3GR0zQ4OvmTZoNF0AS2miK8nLwyVKNZmNcMnqwB9PJO29TpOMKN+zPjIFQA
z43IOxumipio0np31VK5DF/GUgYcMZOiC715r41VhRguKLj/zBeNUgGG5Eh4XC7ULwW5NiMGVYNp
tRlHtsEKMR8dWvmHHiJa3ElCcYcLzL7YKUnpPiqocaY+It3BCRTHdmmxaB2b4d/wfBK9LpImP50k
ng3sNAXcC+4zASys1uqey220c8ee7v4PbjjOQBwHRhQvvG5oOkGo2dQ6QUGMPxl+82rM3K02o25K
HJ4noRwKCAaIMCRYMoE+fHwlE0d+SVuXL7P241CQzMEGxc8QDYFnWC0GpnbYIEV1v7zvmbEUl/mI
VwQdlRl9KdFqoOhOWq+ZNscUxrciQDmsh3naXBZKe5Hgbgc+1wc4F2EJipWLok3fTrm386ySdyFG
k+DnyK5aJXwFE4lZtM+43WOfr9nXRAw9uFksMAbIyERSI0TabeJyd0SOGYxGhwovvnq8EzgufIRC
Sd4oRX0inWzHl1vEbvVfNpx5z2HtB19mIYDTNzFHxOCxTVP5UxbZNik2MOg/HOAWNdc3+e6anM7s
ZuAnuieFq4m2gYTPSdPDU5jMbjyDsaN2paIY+d5/gdtMZUGH6REtUHq8uHTz9hkfh1afDWEQWPNU
2A7uqE6F4hYNnPeMJ9IO7J8xshcz0UnmE7RcuH+4127vee+gioZthR3SIJ+cZilP/qu+V38vRwFh
SYShv/FsHGP9gbA7vEpfK3uedO5SOnRD6hMpjucFWGlEkKVJ3iH2t+CUzHERoVZErbUjRiJAT1BS
EjxCtyPfr0VF2AHcS/DnAbg9pZSTdlQKbkYIZAvdm7i18ZqVHWemv8/xq8UiQhCv8looi8fytLpB
HI4Eb0EnhuT31rv8tI8g39/mOTwH/vtVU4c50kJfLMl0pqLQo9e47qbMghLfQzfJ3o6Ne6p8289g
PwyjCtJKR3UaS+mU3e4yzT7Hx50SBKGpK5gEvGKCyOD934fAVEUiuol+a7/uTwvCPrGBAEKSR6qo
XZNBnV6U7rKdIlJlDk1Tt6cbY1OSG4hgOk1wyBpJ2O5GU9kouxPDkeksro2sXY4q95isjoLq7wx+
34aWIexGwG1DQFvuP4wzy77yhkcK+rD2ohSuC0bnwt964joG76UhitnORjfyWY7S5+MjsAqYPfY7
21gWJAq+XXt2NwMA1OqVlFzGg0IFzNXa1PDHBRXEhOsISmXHb5LbbDfXqTW20aYLXU465It8pflE
N2rfz6VLtc1Pkt3D74dxExkCtu2u4vWKODiQiYTmLbxgSRwABzcSFpxckQf5BsOlp9eJ7FKtmBQP
fSXvWzZybAmLU/hw3Lznr3TDseTGBbiCdpjzVM7oByh52716wMEXFvYLzCU4pnDNPF4hQZSp5vlM
UYp6JWBWc/eeo3TECEKF+pY52F89oEg5CMov+4waVuXG51uLVa4w84bubrd72VdGS+zk+6ZMUSyf
hMsEUTSj8rPBAZAPr+A7kj3kM92J/l+JPuuSjXaEbD8QblInwZ4UbQmLq01/nFy5SEW6XlhtKpf8
2rGM+uSTtjOLpZET54G2rqa5GByYTR2w9jKHHFZh3IX6rcU5ilWqZtQW2X9xrN0tfNYaa8K0P5dG
YT6/TJcCXWLd5JEPCXIPeFlqssa3nnI/azu4rt5oIS1MuC1eoWjl7WWnZHLr9Hyr5b3OpMdisvFt
9M0PgaqC9bFJFTZQdKK2+pwx1G0ymnxaBWy6QXweVC3MIo+WXaQUimi9EYQLsZVJUnfCyw0oWP//
vqItTcqQi+jSk0yv8oBnjb493NJ4ij0Tsu/ZdLpY3YSIJzATVjow+vRrx+Ons7bYZkr2bZ8eNMMG
KSwuxbN2HBEIaS2fyh8sEh4Ru4f7EXyalCs1cQ3QVB6EdFcywdgZ/u1i0WpxGajeGbbTWvEdOE6F
ET7DMft+2UESyBi/q1CCccm5HZdU3AxUsZhSebiLaDfey4PddHPlss/1fpaGntEY2eIR5uTBxi7T
E2nozqj+P5Az1g9rEiOvkqu59stFoAainy48xbJKrzdo1AmZ1xkHIvSVSmQAfukDu/O0fRenRX0I
MjJTKR1czDUXiNrLlpw7ADZ5jQbcy9Nas0S5gpa3lB4A+M3Mqv+PJcn3yN9Hk6lZUPnj6ACKTNzZ
QZz34yv/u0lhDaddJJsZg9PnhKkSUME3v1CMkP9TR26sUeVwlbPGp4HmkBKAWpx3LRrdkdM3YsXG
RqF15fw/xP9BEiAIT7OvhPAETrTIBibbJ7K8q9HdWtjs5dWBHc0D6k3QXiDnB+QflPSJuwjEu07E
9EmpndCuMKiY3jCUBMtMv+6BeZmU18TWmvr7bxveRcreqD5adaeKo+FdZEw/KWr/fh5nPfm14srX
s3p8ZZW86BXFDp/ROhUkzRhCRkcnLLuPNPxA7NCd+QryyU1UopF2E0+Sh8QA8XLb5cX+4Zn9XxHC
SHf0D8DJ+2kl6KuR1lOkA/SioW+2ksYYh72SRt6863A8zt8VfVKYk7N2Ra1mOG5UcUTL82ruJAxf
Rn0vL2jy9w5eGLSuhdqIU72zasj/y6UX1DO0S6Ek6EYjBy9Th0Uw8TeN0gO8G5B2Xna3Fx2lOMXF
g+ZBHsVYUbReSvsXqOmyWBagg8bsU14PZUd65nid7QRLJmYc4hIZ3rIfF9qTcmmFHsMWGBHI3TTO
Yw78zfCw85CjyM34ar8Yx3OxE87tka/A2pQFtUfXG5poXg968zegiCsDwObilVlR1q1NFQlE0Bcm
y+06UbuMlbiKTf1nR67IiyDFF2fIoz8GyNS/ft+c/uFwnZwhfTvjF5r4c55HEej1EhagOAyNYqLQ
9CZrIU+J/li1BMuYNTLQtiGq//VMv/32ZYqXF1ZitKhlXKY1DvNWF7mMcN5eZXqWjX41rJQ2/XOC
VG42OWZnYN3SL/kqHOlNXVmdWg8SU4de2q8E+BHmKbqQpRLqb4ZrrE597V+DcbjPxOXEFo2TB5Yw
Fn4dQsFWsmLPtfAmvnsBLgL11Bi8Jy96Izhl0M9k1L69wHZ4JUAjh2rnAtOx/x2h85xNS34AKcdc
1Lx03UgLd0wuv+1eNwksiZ9yKeP5CtHrhCOf6jVAK0yczZECSmS72x7TMBdHSs8pSUHpDlNqAKlX
BGfWoXM1UNO5YYdSwTKst66sOjsoFWVrTtq5S5TeI/hRF5783mJIpKrTewiuE0cmPVpS8t2Nrqby
4nt8gC+pBaFR+XJ2q/KSUDdGvhEYoBc/P4k+bvHUl1t6U3SkAP+NQVweYVjWoVN6fUz6Et0h22uO
DD5bzhQtGO03uUYq2UXsQKyNA7NB3HZQO0MU9R0cxmTGGXqAny57NLg6HuBsBKBxCQ3DETB+b5BY
WjRRCk3qej3aNHl4LQZXmnlmmrJmnR5+tDHgM7tkGyo4FRSUCVZSkLKCH5UMlW1cQsktx3u/ll0o
evWh6GvfcxnwbtZaB97vULiL375GKd3MCratDnM5tLxY26lmArxboZT33kNx9xgXhcDA1fRcoffQ
FCG7n9rUA87zbX1wDLZkX8kNS3SYx76CUO27typmqwbbjUOSnQrkQ3Z+D2XuPcG2vo7BJyX5OY/2
WuCuqFFWL8gjyliu9xjj6DMmbZ7Js/jGfHls/fW9Ar3fkro7R7L83xIBs/GW6nhxq4mOuWYXbdsK
MOLCX5Qcj3cu96oh6Zc8fmp0Gm/wjKrE74cwW6263jdwP7VMx7Fqwy1F77RACz2XeuaRC5E6SgYf
VYuFFM1Xz+cNIWS5967nzi/BrgX2DVQcoGZI4Z5VVcBm6Hx/gV3WXVhvjDL8Yn9kg5JIvWiXyvLY
xLm1azflSuj88DUNxBCA0jIVJPWSaBW+XnWQprtBUebDjBilREnBJSDzYT9XtRWwPTlivyMU4vKQ
+M3w3sa9RImOmPtekGyxpZ/NbW49FHV7Sy5t62NLZ9lYUSnXNxDPvKp5tXN3yJpLO9pXZwVtucaV
R0NBSKJO2t4tWb5EU+cS7GkvrYxMb+uBQsVQ5nR7ZYyQifArTc+3N+12BLSakK0rfWJPix8aebzj
rThGGM42TvpiIX8OgeIO83h8j0uo21jm8eNvWXQcgFq5WaXOV7jc9SOyophTgtgDiO1+xEO+TEDQ
2y/V08IVHm5trYJdjZmYp3DtBnE+JmeAV3RuLKaG+efsO6kfg7Ttkvi0PW3yliFKWJ/56iDDGfv7
OByD4Lo5In2cejqgaaQTeA25FfdWlWcmTnpIjq5RaefHjWOmAXRUOFCVRmDi4pACg6LI9rxV3IAc
M2em0/SLnteES2zxYar/t01DPc4HJNkEuc5zp0ysc51E9WOobbQC64FIcvHlcI8x3pl33PcoVZTj
iqDK6V9J6s1UVa7rBToU2hsRhLrxDCEW8Tsq4XDnfL7InOR1syoMKBc96GG7fgojhUyGzKxjXVsO
NJGDQnxyo/5n/i+DPlo6vLs5Mqmkfj4k5IwAANL9FzP7CzKywG6Txx7hWYu9Db9f0NM/p9RG6Vd+
W2XVU1x8C3+AlnaQ/+OhLeNMLLA9alszNSnjIu6ajwYdJv4QJlXFfOq/M/MZSidoPGfCJRK9Xon7
k7lGbIpr1IoY49N/NRKVE8XJyjYw27P57GvMxCOnH72rH4c1KvYncjHLDmr1qkTveXhI02Hf3fV6
QcQ+zqp7CMeazaCghAlzU38d8yUvkbcbK9WHifB6OaCp8CKWjEZAtMrVkY85h3x7i218tsPLI1lT
/WYCicXSwMJtaMcEE+ZShmbTfgcNhar8ymAj1ewGiDeh3fYHl/W9k4aenl88zUXrcvlHhaZaGB1s
Uq2i3gscITojhvaxOJuQCgjpsjpjTgZK0GxOMXykAqpFeN52Q+SmWqYbQdm76npdp8Np+LCyL6Fk
a9wAfN57Ba9YIVo95orm0viLh4rQcFEmXmeyVpfy1/+4FGBz4Jm08rNkhszeu0qeD3p1lsVG7sS2
eiWSJtGqusGKFVd9nc2vubr1khCscMUIpB4N8mQI8ArKhZf8X/GTTA2n/934OJczpodv7adCLq3c
DpTkzWsNIsaUPqv/0Dy23PesDILaXzm9D4MBozNqR5JMxB9AMCv/3cJXMXj9fTbB/aVMO31vYo4T
+PWLGa0vi2FoOQgrddSov6ZCmtMOgSFQuKMb8Kr+F25WzNslqviNNJjsjKp9VKvIbYETeTkrhnav
dFTT922swLwOxUPZs9j+rgLVd0uwUNVG07NieupuAjabWv/pGnvswI1NUTiflnEiLLkK7DxVWNiN
zyDIr+46shNoeUd83ZJLsg4AkTSM7eBKw2QH/78+BI6KdXW/OxSymqKnkQxhuk5cGsnGYxEx9tCI
y0U+cvohrewVnzZ68tNvRNtVYhWH71ou4gtAc4RRZcQkTS+r3ScY+0fOSTFo0YAlgJXL6FaY1vYr
Rn2LAeVdAzFpEwxawRclb6HdGjeYhUUnIJ5Ml7TaGhyzMB+TgZqXNgjC4Tb/dfRge7UXwf0S86Au
tj9N18+jt1/eLQiwZIQGiMNja+i+Te3UfwHM4IqSq1K/Rmv3ebCGVBijqXdg3PSBpf5c3vCVoE6v
FqJTGE5qSTw7roj/zkQ+Pm9LloLvO6WXJJ0gDUFkqYqFlLxqEEc7U1wM6UCUgElMNVshDqLSgjOy
hhBawXXG2+sdHWP+U2fGE+r+fQFqQssWu0qnDgHMh9HepyxW4SR9hrRUfGQLrG4etSb3PRZvaZv8
AiAn8Bk67WWgrRFq8nhiMFqsCxgjFg6M2lL8hxkDJE/g5pE3IUbGEZ8zoJqCCpOah0f6xbzikGkq
jlHKOPtubfcyLYWAtSU4HaTpm9cGyFandFxEITbM3125bomRazee8rOrLLGZ0pvkhWffDmcmDabi
EhwfIdy0/+H05QfJdhBt5GyFLmCRiRLt2Fafmnzx3gDOWKasFvYqIZ7nwQ2XSCeoOveKf/8dEwcg
dfsiLs3fv074gzewZa1lHi6vvfQc5MaA9/Hz7e0wy/flwFngda640i0oHGeRI+PVNRF3hlPY2guP
fDuGSVJbFle8T0AE+NWs90v+3Ontx50LISyuMgwrl1pfzo217rsp+2HAiVVqA0m47LXu4d3oats+
IDVqpbMmET5wgRBUQryHtsvaDlO14PhTlEEuUbPKniCbNa9AMW8gMijY9r+8gtiAdnDN7wElicDU
K+8BQa74zalnFzic3TQQeMNu7tDQ615OvGqSpSYfb1T310338bk452j6C6OPPfMdmwZeuQLjTHKO
/R3gYtuq8jrBslZXmSDtyqkSjaeTUMnryF4pc0SBun3BB/e+law9hoX3epTLoFkQy5DKLhOA581z
8UMmAR8iFo5YVZfvRbRWoS9VQx/MJlS9nacLnQqlH1kFUMzE2cnwsHInnrNEbvnyIkOd2fJMIjvT
MvOIBLWJprvZAgz/cU+revWOn3YFsFbEKTlNQQm9adl3eZqpOxGFFW10GRML/ZeVsB0F1oup7Fnv
sC/X7jnbAHZ9Um2XqmgZv4/JS9vCx3S6BwJkDnK60TIFaQDQEzemi7uSZ3zN6pUQKqP4OFa2pZhi
LpMQcKFrescrBqAcuGTouIMxQhgfq4Jeb8o/XPrX5hq/dFrT28Ay7PtX2XqafDfjFXGg6tKiJZA4
3jmfbxFAd/thZkpqjdPZ6ups3JPkq6uokl56FCPVIl8AUv9ynLkIPCZ6PUTCBD8RtmTIQlLDx49y
3TQc1qDFq7XWv1L7pIF/M+sWHPbJnaFon1bF/cTPodfheX4qUA3sy+GKbb5SSOIAEmX0qfcSPpkO
tHk9pMgj9kt/6xOxhUIS7I1/jaZhe5G4/v8sQLx9LEPMUUubsWMpN3Pvqt1mMwLpK1rA5LYpcSBR
/00NFvlTfoy14yBhIt42rxrz5FcTGLRMa5BAmoLGOz7QyEr3Jf66wOM2yfFRh4azyjy3kEYsEiED
JOaK5l6og9no6+Ia3Bs8SGdKxt6GgxKrKAGB+rf9Ztw8AP4ILyywcHZEIWHPwFB+wx8kl1wSgCWb
mOZAfVtPQj20/DSc3/aslDFfg5MrwoQr/+Iu4zj+h0P5uAP1jq64rQywvcsOajyVUmXfUjqGLHzX
h262gFEzSp7jRZ2lnAaV4Pb6SQCkavVejo4NcfH3LJlamdr4ST6OToP4XkovQ/1ozVchOjIWub7D
gS++96ObZr+UFmzZsKDLmp9u4rYUNKQKfSYcG6kjPz5yj+S1N1IIjpD6bIpMk1SOy/+ljJYZj8ZH
Zl2La6AAFezr6MacLIHnE3Jfk/IJHoVi9iRVBeD9pU9SN5xlqYFTr9pMQ9Xs7ayrOFjideJZvRLz
jg0uHHPSXpE2pGa0TFZeTLh+oBhXW1oieIhP5Z80X7vqAAVFdvpI9+9G2aq/U8ym7GRvYCOIHJ6+
NRprV7o1vX1gU8oERBu2sIr9TLV4AXOjoV/MkYu9nL3ZA15Nrppn3HIKRG0g2XzVcFyBSxNaalyi
ZP3AjZ5tXI8FtJjWrNs/SKNVRRmcSRo9QA4+32J/SYnh/JO4/RUn2A7tuM0xsh4fxcbOuU6eIJkU
SxugSy8/blfBL8CPz7FA+IkL93hNZ761UCqVlFj+f3X52DiZJKS2sA9wozqPW8PLL4oSF4OcRntX
BMsuKVSFN8qBkYXHlBQhPZyhOYwu0C8FElPlOlMP2fYNm0inmuasxhRuZivTvq4PkM9m5pdMzMI2
CvzF4U8ms7S/KdQYIhe0Oh5HNuuav4hxHKzltHvBPj2uyJPfzdZaWGForSrrGrqunnX+C0DsMw5k
lPGzzKwj3otRKX9B/8COiRZb+S98t2WyqXGqzsANBcZgjf1fQK1UBes2tCQwc9ONBwBjjpmfutMr
Db+QTVTQaO/hCPP3GszUtnSZGhuuBCOKphnXUBuzl7SW1xf0zqXCliA2fl61e7XkqZQdaUZ+2B9o
FnIJeAOja6UlYzPusaACQdy1wdUY4GM+yK7zNnYP8MBUMHteFyqB19hrDikLiiRkrj+Cl5qrz8ZT
xQwpRtcX7BZRjzXtY4CwSrBNW5V6iBKrv9/ZrN3wSX54xZI5PtYFtkmGYEi0ghan0E6yPlgDXxsd
xRYju+8k+YrgPJSokvnyoKCzkw6YW8yXXOt/C61AkqxUq+J6Lh3neDFMhr/yQn0MGohY6gdZISH5
3m82jmcF91R4sT+NGEwcCrEFILgIGX7yoU6lr15c80F1diXi79gXEunHQC8JXnW4Y6dOrLABtoKo
j5QzWrx7ea67Ko89k+y4xJD3m9GHs451hkWQB2YOAHAOIBTu7qy2lajtswSIMCjbXnQVashCHKQz
Sj/fftwimfjNNjNmFWv3A37AKVJOqZJv57pcryQcBPOuYTiJyuV8EF0O4rDiNaJScCrg6PVl3ZWU
uzyWquyTOcie9Z8nlTyujLjik8FrJ3sOpW8oL1+M8KyqiS4x4PHjdPFYVekugCo2cw8JH4WEbcME
n3RR1FJ+XwentdEBOnWHarz3/ybue2gF1nMTGCurjOGzdiwBD2GfqalWojBKfj/rQiZe8rKgjfAM
NzRzWfscr24g2Pf1uF1kdDm9STAJt9nwcaCZChM230se9GOPxdSOIayD99Hh8R+TzdBqKZmCEfYX
baBVy+nhJ07PSSB4HA1mkz6QdLsbT7ck5IMTCCHc0LeRlSpyMx6fRpM9DH+ZNSMH3NXDTAmGvcI9
tQeU8cNddgkDYf6zGC253CqH69WZ58kVL8TZAx4jtYvDkeS5hq94yi0kxgAfr/5eRMejWVlPutqL
sd3G0wSfs3LU4b7drHSLsw04Vm4BcFhvRtzcx7tQwBjzOgEgcD/5MnBhj5Htb3H0JEJbLD/qSJb7
lOU2LU1RD3JOOsiTe111x7BTZE6Hl+PMtJQ+ItmSRxrj7IWVyY/FhqyjjkqK498K2Mo82xryMkBq
PZ5c/38OZeYbji06Qs5tvx6NtER1vPGNETVwx+TLDvXL1Xec26M9CP0JPvHYl6FqaHHnMYco3012
yO/8TIGEG0Z/tTGSDMqsFMzWSRJP6BfvhcvRFNgnH74F3dBc5IXK/hkyFFK+NqwmeruRoAjkeT43
qPGd9CsJG1QWqX2x+saP9sqxkIBjPiWZDIFMgjyLyc9Wvnq9Qkte94X6rXEheOLxWTAqtNv30YpY
fGmvcySk14EuUFsH+tVvx8tcY25W1WrYoEJo0cXLU+e0OEgpaT5uXJx6Wn+4H24+3jCEuGeZnueZ
38PIGMucIZloXF4FMOFqKsO1+9OSr7xMu01nxfZB8LJv8RAq4A8PTThH+v6+GZBuZKVUpRD1gidP
JKkAnbEPgUfSMF1hsMPhD5vHIVp931tfF1bsP16aQXF7eVxz6fTnxTHu+ijwfa6+EoLSpVSyeNaJ
VXWWeUwk0sNGrJUDUCc7eILFceknmyPuDKsQKuMmAMEhReB8SXQ3RrjefzsXfxch5BBvqDwsDMPi
+8p+g25XYgKuBgB9amEE3RlL+Dz/QDvkIKZvQiuHNIjdPAGC1Sa62KoxaqFgXy2NjIdZXuosPu+S
HbjbNaC0hkxPNI0Mf7AW6fSpTxvmLyu0GN5mxzhhoZsy2e+lHyItBhYXz/sl/wYnL2KUFpMgQSQD
/5i59GOtKu/WgzLwmBLhE7KrlkPxjTc14UBQ8YqJvV6AKEHo9iHDG0w/NPPU3J5HCCRa58qk+oHx
ncgMM7lroKjiQkZSgye3z5/ZJc+tJQW8obN0jlIVRsUCe/dRb6g45zdGLwQ74ZfjEScLqPI27aQY
huaGmFvA7sHD2rLiVo9zDK4i97od4Zq4a2UWXaQqTL7+2vCVgIkZGH//azxagkyHMoLhN9wirj5A
7IpZta+M3Io1yjEwhhX9d5QnmJn+jWVVCoZlKh5CozvJtH4FB9X9tJcTiCQQaVIR5abI4NL+NX1s
TuVZAshfdmgW/VIDx2sAJdseGxTs3Bg6F2jV9SPT8/x4imQYOhJMxNIsEnS7C5GWSIuG5W9PY3in
G2XM9AKDss3thPMkF8nQwHlwRBNf3JCnIi2re4ndr+9nrEqvdRnTDA6rqVzrNJAIq9fohMUibyUT
DRtt6ltPqPHFkhcJMlfNXY/9oO6U1L5Iu1xxBkGmYev5kEwFyM21VT5zDvrZn20Uz8gYg1c76POc
ECHcwUeVD3gtBlmz6alWz9usitu1B3Gvz9CYCcyjOj9DPKSthXvahiByqUpNiR195B71gmFjqWM8
EdgZHA7jaHHjdt32eRhKMxOWPmClBGcKca3GhSkxT3GYtxgTCvIG3XRIm1vm7XPblJkT4frLLer6
5R/CJKgM7i/N5QhBOOqwW0A/IYExe/aqkctZHW4EKD30T8yHNbVksh00qDrXkreazP9hz2Glwdwl
gj4rqCDmqzBYgPOngltRpBr5p1sVl/bwTVn+A93jKvZzd2pqBlyfEH3wlq+r/shwh6tlVkljSogd
x2YNbTdfG4lnIuixf6DqrzzTHwWVCe2L5LCOwARSl+4zGvGoSUqhAkl3On29tWbuuBVm54YzBLWX
PNmfOSDDG3z/vv82JThJANF+HxNhRLRUHxrf6qQIJ5kjtf5zM+YtBu/2lZ3bv2fC436CwjW5FS/b
bQNt13yK8oVFLs4JHTF9eC2WgomFxkW4Tk1S85aMOr1HDT/I29PRb3j8gND17YvDLXsxJqA+wPAv
YJrf+LmWv5gs8zrp/mRQo7qTG94NOLmDrs8GTaUjdLWEmA6APR8K7poxC/KXY3o2E94oLXY58Qo5
/45TtuGZrklrusqcjSzwU//+n6Y8wjXGobn7hZmUpoJ+aqGGkE0RdsjZ41Y0Q5liM5fJxbevKTsw
CGqzD+TpqYFyRlkCuJXPKdCaHUx424KSOnJ6DUdjkYer0TXtetOj3LkUDJZxuqVQYy6dS+NATmoR
bG+zG3krpF+vp9EWMedp7CtqiKOJcBTJrAdTcoUUoAeQnewb/Tc0q0iHoV2VbpdS74d3v0e6HRue
rhbbUL+CaxVFaFhf1/SD6tqLXqCV9SLCBBd3ohW2kQlTm67OFKlGKxdyTcL0+6eWrzPKoeiV7JUA
RAn/GnSq6Ngfvga6oaNub6szY9QLblZDI+dyzpYQtfH4Sy4aE/hO3Ke3pNu0q40WhlRsT6fagh+y
/riw2WPfkeF8Vbkt9KzAs+rKO7JsdQmEjzFq2Hl2IX6QEkLGVpBnzG+39xByHgmeRxrMcgn3XhRv
nVIFwTYwoJ70OcCa69FdvY/bgoGCTLjPI+e24oz3b85HKgv5j+O/blnsXNjXzd/Y3XsSGXMB0d7N
mxCsYlzgavpriQhko1Bmvl2pkGQxSxtCJaMscGvNVXk/XY6v2Q4yN0DtdNGROze0rgWa3dkdk7jf
gyomDRDiEtSeWM8zqyyk+84CKCE9QofHdYRRgy9OUg9KWMYT86XQrvfIsdlay3NSY2bZVp79oYJ0
35RO5fHIur/cNb2kk2OiWLn6e4r8VmnBj/5NDiQcnkMzDMTaNFtatKlw2tBE3OzwC64xrZUdIqFh
dp4+CLlsoy3hfQFyMTCD0VoneC6LTjmuQMDVc+Sd5UZXho11v4EDLONboL3hOynZYeeK5+GrIKdp
i4taCZ5ENtTXQmNAa6/k0jelpReGo89kOgQhEclaLkzTWiRe5motzc7paUXcmMYXabIRbhLRiu9f
7ebvkF/oWGV2YLCHJSJx1EBlLNZie4COX0dFGzRo/ZeylE4Wiy2EtHe0Wvdgnebxbn+65jfMgZOX
0bDHriqyf0sFJz2sLh2ErwsQra4+01laL6qTZXoIIRu99lMYcEkhsVH0efyxi/wDCNAF563iyYjd
fdUHWIoPXEoXqY9k/twrICx0YlVIWn/00nXi8L+aImjXQXt7SwBQdEEuAV92EtkMHyAk2UtuvZtJ
EapLJ9abHvvRk7Vf+j2SMTL5BEYzqItBo2ZmexxlgoXoPgGmcg/u/buWA5L0aXzIBJV4hDSu8vEo
sQ1St/NhnvJwEEgTKPcFAhi2xOGGDWKDnIeLdigKL/Y5NFKTuRPNzu9qYmy9oOJvIYw9FlAheQyP
Hz/utyRr7oIJbITPNRf2MmmCn4xtKDlAmyDhc45FcMv8i95WISzsw75Adx9EmFCr8aKVlV04Dyzq
DTcMRtuZ/yWIJ+BbpX8M24xqX9syKEnKdRamiXtb2RP9r1qDPEGf4f7KwDyoDm7wjvzRWhVfqhre
ynXP7xlrSqrAxOmP2VaBKIbwqhagOS+AaxSBVXK1o1NzEQ0RvckborpV2/5o1N92DG0UVhSNHfVi
NQGd9jheMWwM5t3TM1Zf0VysILnn1XS+9viVaS/fZ0Oj9qYuHk45pS9vB8RcMKyUO/mD0jxgiyLg
/XZLEl0LyRFlCCjc4ObgCe6VYW1N8jy7mD1FcSEIPGe1EvyLjXnDZKnlo4g0+aYdu4uxI4aL0Hja
BNUPH5b81m9jNP7xiOfusVgFvm2h2v5tEL5GNEPISAm9DlMr9ftP3ge7lq16rEP6tVHuvCOW1yON
VAVU7d0uPm0eCv6LcLdYQzqrQBJbRqDTcinf04l/DnoYcWvSMI1jS+4VbcQG0/nwxBCLHDgXRs9E
0yrUX/htwuFSvqnIPgOfXWluasIuVSvJuklJjL6+ORPw4YONqrrnb8g73w//LRplyy65Nk2/1cJ7
FYgf8RpxbPioj7CJG8uP1XVMQ66wENE9cDpqm0RcsyyO+y7118gwgfjlsDuPKz3ZFW6EAh8RSU8l
ojO3P6RFF26Sng5xUBEW75O+Jo1w4P9xiQ9iGFwE0QvHUvkxh6XaXQqfZwSkecp55RPPT+jCIP3W
zYz5D9SVaRsVkzQwN8j9f7LFMGXEySnAnFuo4gSHP8qGIf7N+TqxJAlCncbYDr97LaDRoKEoq+Ye
8KRr+X5ev1ozUUsIsUXC9tNm6KQieyZ+60fGDu0oMdc5bhEyvOBAMc+5P4FpVsDGcMZcnWqkuXjd
rLG5+useLuLf30p+nCgpBCO0STmm6aCyWlPhhbBC9z/lpL9YPZlKaubiNx3hTIcQihFcbgFrbyNd
f9jgTOmPybqoVkc2AImiKjhTB6qmPaLwQWmmsCswk1fdlD6T9+SQulo4auL+jxn/5VND7dmgLS2I
AaIs4XkqCZZSU0Pj1CxywKURBZ2p8QisOrhh1kHTjQRVdJ6arM2HM9bdP79iNSGKWGkeymNPa+fj
dCGzQ8UdBaMefsBtDhNey54IzQZsbrEIRI2VjpOF011y5zlicOocmCNGOWxeNYbGCbpWTfDtEcjg
4gBvJqVeRiX/xl7EVvi3oX0/VyvSlUI8TBlv0xzziNUdwNUyZNX5EFSIYoNuQznzrkgYdMftx3i8
cCb3qy5baeMzRqr1B4bEYW3xfQU1j/+35q4gYctDcsN7HC8y4F0dNLndlNxwXzL2vaq2ewe0aBiG
qBudg6dIFiy3eUPnwvXHqG2pqOa6EJNIhJUzTLkAgp2wYFqRa13eIwXd7Z28EI+sOJvvd33vhBD+
oCUa+Pj1Xxuirl1kjK2vWUY4ntyOAh9zNRK6/UkofvjuctVD3hyf23LrMJKPPhk3Nx28kWWwBfuQ
ZQUu
`protect end_protected

