

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iisr0ydwFOm3eepmhOYSaxO3flYpViRsLN97vKyw+ai+x1TubmaH8qRRwK/QFeVsjlGTFdxookcr
olQwv0bmdw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dJvTzz+PoD3n2Ot9SgKfpEhIshJxklhDhS1tYcrcmprfs5wN+lN+5Y+o9jEEql61IqDkJEIGu0xp
zaDWEeMqwkFuovmZnp/AnbrHb7R/19zPRtwSyZ8+VQRLsRMgscwutXu29fTUST6Ribitutae85tQ
1okc5mYK0mcSMIggcMg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZijKIWnBSOuwn6R4ZrzJp1qaSPGZMrP8GTp+SV+Sn9xEivGxLJtGM40xMLXxiYuxIopDD/A1usG6
HkSoNT6OzxHJWKkUEyyVzrZuJdNHJ5q3s3y5LSNY7eMxN9lY4/gygh7aVIBAO9YWzsWu3HLtrHA5
2vsUFQxQdkG5OTLVP1rH68P4j/dhqr/LVHw+9H76c/knGyalpHLRC7tnHQcfuezFJWlkzaNGHfUo
b5cE1YTvtdlZVmw2sVG/GbXIRi5fq3+Okdy+JgckZ4dVWbI20rfa9LkI09/kwD3anyrnovVQVx9h
F0AxolVKVVyWNAaSu1fvXllqzrdJiRLbdnsq0Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LUajPw/jRTLlmEKb+9YylQ2jxw4jlSx/1GGaY1wFfWFdMwK2p0xvQMjui8K3EqJF0fnb3QNWuQDl
1vTtf04vcOAHkfRCeW7Mbp8qeUTtAsflGIPJDxHfVU8ZKprwANsENc8LVrpJ0WnjDFQIzJw7LDqc
Jj2TofWjKprdxXsMnu4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KG6kiSPrd66zvVpG96eKD+783ebVLVFNF7pXgq+rCyBBRoa0N9Hp3DIWK5125mkICodI82zuSq6k
C8aCiPbDiv4tiuIn19WDNNPL4ncknL0KLZTLAkq0BIQIsnFNRaZegM9aXOdMYGKYLpnjSD9KRWRt
WPXPZfwprSu2D7PeDZMiij3MY+cixttgVmNfcx9Kkmvg+1B5sTSDTVs3fqpJBBO1YslTmxyJAIC6
uDuGqvQ1138z6f4f+f8vMXratK1Ypo3jPPb4FTNLYJio5Vd1Nbpl9kRRtj801Ie0GGhbggK6IXJx
785o6wX6g3tRyoHXGJ4DGUmWlIHATg0KIAflYw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13424)
`protect data_block
OHE+bFqKhYn509LfSse2jYP/MV2PSFqs4kVnMU2LGTrYmwMdpqdxGqBqn1hsa29YYA7FJXVUQvVw
OOhlY09AQttcGGu+gAj4qF/Ngz0qT0moN9OpxP6AxjXZhS/L1KRZUbklHM7FMvzUaQqxVFb0Dfcn
X+aaXo11UyuE00X3v/WEmTxRIC1Gg/C8MZmzTxxMY+q7ROO5pchiDpQRfFBbYJNkbTVsAyCNtqvi
TdsBRrVIMY0yQxKGUrzBf0FtCaB+uGW5H0oHC/hVXBoFvNRagd7sOY1Cr4fuSI0PLaEt/dwEWMlT
lWnod8tVZeJ1lKx795gmNQwl1ggjTIKGTcH5D+UjvXNbDXFozXNBKi25396qew4oKXYP4DZ0HFoI
JQRmElJdwNKxD7GXqavGRV7FC2dQncAMNqRoKQoeyxWiBzbIrcYqbPYF8m+8F+HSGsMy9PzLLdkP
JL0SHh58uJrc/OcK9Khs3f3nzI4+VxWjwoKOT9h1b3+9wDW4gHcGzRLwvHRzXXWkn6hTvXT6waaR
QHhFyISeq/F8KTaqr4A7BKlwdrLHPMHoXCxunM47VZpsCTJXf+lwG5QRrpl/tScw9Eioh7KbJZ63
ul08Sa8ZxuyuEJGPk458i8/DygsRNGUEUwil1mXbLWfKCWZYvxp5arqgd8qs+/0UtO0SvlnP7WaC
O3BG3Wwug4j1HMga7X47MzEGvCnGGrxg1QnEPuJhNSQAipOWGqWHK3veFKyE396CbpFs7aZqkH8o
+nzC40BMAm4RNi7EV9iFucrhBynykfiH4pgVbGoqMfJVAg3KU4lIoGjxGHIWBBI5h1/48hAq+MR2
2Kch0/mAhYYq+EbLcUNtunbVstNIpaqljaQ/EV89n9SOrXrDhmdpm0sCLnsK9XiuacehVlxZlcNK
v9rjqwjcpoti2lE1eed31Kb7CtAzUkKsADRjsKKZLWVopZhy7m7t0ytYnUnsNynJCmRxJo0xXuMM
gVeXu+pvqb0dUArrN84i6gXeLHNC+FpY9iAZmVcfAFmR30YPbxhoFGVTs0vBtqDSFl1xODTLsahH
rGUo/8fiEIId8iF8p+I8o1+aq8q1TadnyLgpSCmUhZztijJLJUd7ZuBIIohh25TBCzExUOSe0uW2
46Fyf+WG3eph8fWuVj2GgvJe97PrxH1EswP8clWqRjJ8ChkkNgC2Nl1OELcIwBOYBioj9vUgK03I
WmV2vlUWX0rlvInSBswQ4aC1cSRyJ74nS+tGXdBpM7PduClJXOGVavD5oMPRPpz/iITy2CZbwi+/
dkWGkbeBOjRDXBIwZk2EFlygLkNNFRoLqpfSmwEbhTLBCI0Hao1J6xdhJK6FResd3L/teGaLoLT8
7dDPIDgs5ufXaSGnwbGB5iSB6mrefNn5I9sgWNWliH7m6RzGv0F/Bxq4dBNen00fxVl5aQ9s8W0V
kuozm2UQfwDG63nTGHzKSn73eIc77O8PMGGkYYQdMjgpIp31UnW3J1H+U+OOq27G88HmHHTxsDwl
8nM1VHThqHXvzkOmiu7774aHQI+6VDN2OMj29M2IR54/Z7V7C9ORBfo3o3++shqboSQxYQw0oSLF
YwHykFrFmJpe+C13Z+kP7iHSFHboBMKelX7ws+O4SkBi/R3nQQXbLr3dz4h1DM70RRaA6QWgZTUH
bmH2EHTFpkxLpkB8w5l0bCpXgLhMX8xZilYljdPQpSx9JAmPBUShr4yL3f9851rGe4HXylDIlLkv
ocQz1vNb/q5loSgDBKFFn+S0kT70GwP4ZX/Mnbhvufr3zCRiDLw2D/5mPWHg3WtCeZuoxypYGPLV
DPTT9Y28/ixT+U196Jz3w00nahjqIT5HAmjSGmgxWKleNtq+H22OM2M6xbGH192y2qrvvWqIIYRz
901uOh/PyEa83+qwbaTT6o8sFL57oV139uXXl8wS0D8DZlHUEfrUUwjrwm+BMgB7Kp/nbfZ9rVOT
GbEjVSsrDRgRb0P967Fgix+nVNAHyMu0YjImgXnfo8VpcSUcsrytINyrb3Zg/MEn1R4eG5T5O6tt
LkD1Ao3SM4sZD05tFAuCTp4Vjm8jjNVx0xCkMHSI7VLf7fXRCato2wtWkOdN6M42tcVjRbohAUCq
Resrfr2HHm+XvnNuAe6CTIzJ/prjqzyOQkxJum4JQdgkM3hddabMqbmz9tPF4EnfT+nUP2KSlPsf
gtOVtIChzNlpF2MllxXmCqBe7ev2gCFYltv1VvbgvVN78PKznZUWOBBwGKEQvd7wysbbQhRdOkgx
WwS+cewsi+MUU4CVhfs8NV9dpexmL+SuNv/AlGpp9BAkih4R4hFRwRWdyz8HFu85ioNaTEIH8eJc
YDUOgAotj9i/7WB9DhpJXrK8j3ege1WEjrfFHlr/8OiiPgviZVFqLWHCBv1/Vwd8EDsHrHpSBORT
Bd13YLMUqws5qmy0ecJKT0y6BzKAz8TsxRYiSD3QADo+Cah/M+E3tDin8KfKcNk01dT2Qay3ZDcA
bzv4lYnka6dNDao/TO9mQilV0NDbrjDhe9GJa2DC4JMZ4Y+auCvP6T0pPkP3oW5abUwqtlMBfT4t
yfzInUI2gZSHTrVKKzVutGAVkT7InVBAMvaecCdP9SbS/hgiklwCHLvaP31rjIeTrjQmv4J67zDD
UFShnxXK+vcXAlBqkFHFODgFH04GHa26HX90jRZwO0MDmPsCyCGwhn8L3dep85qt4a52J1p4R30R
jLOkhF1D3ddCzfHSM2OEYHJ2tS6uJ88A7gHbjuOh9++Hwy90MS9mCsMu0UP7TY+DfZXu1pZUEzYE
73WEpjmMfrwCDu+PnxVRM5OzNIvKt4bVnQd3A5QVTH1z+OIIrnCxRuygkq6JxNpH1RGWSeGG+Yuf
AarUXyfxKVjn6otCPAgw/vDVyxoDVOcFz5zWz4PF4FFNbHu9o93vhOlGTIJIgW2BLmaRNbSelWla
g7Nu7vlymswZWpemuusVGnS7V8l3eCMjCBa1ymyhBvIveeBlVPv1FhJxt5amEiZQ1NKcunYvVc7Y
+H4hsWloBfYWcfQcLfffOD/pEJ1YRQRQKittkaZA5R8nxXCJygeUM3tAalprhmxl3CzMAhV87IGN
e504G2b1OSvuW4ODQA79Snb0afom9V0na6RmITQ7TxcKeQU2loIJkuBtBqYUb+edItUrAPlyaXum
cpEA6yrYQUNQS0OQ6x8QcofhUz8X3TJNZtAjefTsi0+c+HkRrRdIwvISH43XC0x3Qbss5NheA6vk
hCgQttG+yxhTQpLVqTJd9CLCz7JIVRvlaQCndKq1XDafXrcaidJhI4exzu9YGRn5YN0S5r95e5/U
i9jRWjVM+wqTo/3lEop2i9Q2K5UrDEEl8uxwgK/3CqiVH1QAoYgPQhXdzkg8lDfqyDW8+VipiBBi
MMYo0cOHCM8nQ9OJZzAl4NKBoE/bU/1WJVqibj1n5h/cWMBx7WcdaKqR7OcxQwUCc+HVssMwFw77
dlPJJxtozO8zpGd7iw01wBpjI3xCNoOtBRDmayvGKuy7ROormQyX/J97u5iYmS26nC2kjtJW0YIV
9VDiS4sA8AbAHlA+/0Eip1g6DDyVTWYaCw6BESYQzdI+ezSNJ05mseENI25RqpsGuGjYEbkzOvdH
kaZZPOIldDTGs+P1z+TDDSe5FvVyHm7ukH24lly3Gg17+sq6JNtt1ickBmqwbUEOlxBpyLrsyORh
C/62Wt023YHrYPmovYJ90iv37ohsFoQuovYH5YebuIfbYNkWPAZ3ZisVxSKk5QqMCqz/THtM7QEb
8kckqcFXf4x8eELJAGACCCWqRp4YIgtJkgzZnZGYKrAl/fBzarqnKrz68PoN6K34J0L21UARTxIB
CAbEINR36ILH0xg7h67Sf/HoXq+vPgBZuyEH31kCLyIi0p/xY10A6mYv8FXEZnS9gagAJMlogdX+
HQlYA+JWLhuKfPtQ5Ss/s8YEEY9phDBVS28hkiNVsh9BZKq4hdYV0ZAYnHylWPadYned9k83Dsb4
qdzEHKQh3qInodnDpmf9weMtgBwGbto/8/YiNARjdJjUF68wEvrhTu4vLduAamECq3kjmz0ZoKxN
kRRhoqbgbJd+tPfia6ADS+rzRzdFWzc0QCkbHZWAnqXbauLRafY0mn2iM78CZpZ1KhKZkRcJyaT4
LwA2rAJlSxGZMXJpAmIA8UYUQQfraohxxpv+ZguQrFJkzM+Bfeyd7wMHHFKYEO/OqxvbQ9CfICdp
V+jw7dsLz9wWGtDaMAx5qFR+nJsAh3cKoanubYMQU4ShAfaToYHI5y7JVPDyN3hKUyg0f7ce7ert
BvS6h5YndADgOixHkyl3ShjMTddkHsdrJZ3NeS3eQRmZ6defG/nR9Q3856m9NI6j2IjG+po5g8Bf
CvgFLNvuNqsT/B9GCCbZ8E2Rj77Oy2U5jxactLywe2flFD1+m41ezKCfDAEJQ185yDhxCty3g8lv
bg5JuRkRkvTSEyxYr/Fhm3JkFugvc6ImYsvjNa8l2KFHiDzrMsnj+WrSf2hA7nKk1BKISRenW8l8
gYUavuY+hig/L1Ij4LcYeBES8gQ4B1PWgk96R1kJICPBmSBEnJJftfn93DK0pZ4V4IY84Ris/bf2
Gbo/qXghWJznbNmaWFyYTQQaq5ymtV7Fb+Scj/4rg1B4KtUvW1A7XIo3dssBvLyAqAhI/fynWGhw
5vGzoLjgA725pKqU3BQSM4XHGdhUCYOP20Lpl9wJ/YiaFnS3s/+dg8K98oEoQgSOW+9Ua5ugncUx
OJAh4NmPck/ovE3O9TZvtTGTL2xKm/QoAWQ6Su8cSonogvvb454A7TwmYSVrbjvpRbCC56sK1qLs
CAJ8DkNNDpAfj1sbSULkDpYNSn1V2qfyVk4LKMbvblf8yShgwRjEvcj40bhabQ2AzU9tIy9uvTR0
zwOx6ADADCfAyd+t/EIpXLQRKRkFRUXdEYW6Ts+zdIQYqanJjLWWdpwoOzve1ImtAT3z5hhu9Xef
GbjI1uDlDjcDEFn2YRhyPn09njdWY5VpZRpAWBCMHHk1rARupfVESz7s4+v8u4vZWxvg6bleS0rn
bX6Z7YdyxnSrdbk8SrlctAuuKTHa33rd1pgxxtTBjkfTZ6P6n1l3yzDP4uA2VvsFO1famgNxHUpp
982L5aKYEiBCmxM26I7dz1cg0KS0QAmzTEeE6xir9Z7CaW6peHr7zRZKpHrbyD4Z4cudEYeUM36D
XIrHyeOJOENohydUo9hQ/g/xIcBocgP8UXr9DKpvvfKE70ODWgv+iuofquoSn9SB1kAR4rRLynzH
1DU141gmaGqsl/gWy9EGhUZSEuOXPoaEH40c3Htl9Mim4BnRBBOzXrdU/pCczFV1jLWD75HGifdm
pOdNVcEp7wcCvJ2BSF9GytKttZwfx3CITEcV4R4nXiZvkYvNV+z6H7By3IxK34DyXlG1a4R9rXBR
9R3+SAST5IYhiSrC08okRA7HuIExScr+GwYnxmbTBkx0/5RUmXJ52f3jafTmJ5OSZ8ippag7dt+k
Fe95NjcniIAUHi9M/bdwMy4icIq7fBPX99h9mH7rhHbXasLTuFRzRtIHAI5ERs8BWCbfj7BoeJOh
q0PFh6SLmvFwqSCC6AqeoMpiNutHrOXz3KXVakvdb1zOfy/GLK4C7jo0qPJBe2vChTvsf0vD6FEN
8x7w8WqzdQ8yO8hD4Fn8D4jXdIU3Bs1mzfVvhc6ZDqhuF731TpdQ+d9Kbwrt6Mr1+nDDQCGdZASn
BkKN0+qUEoti8oG1/07SGcJQjnzgmTa8x2O4PcVBUzfVp3MhXG7fnenzsJrBRMxSNJ4QmUbMZ4zS
COsBGFGst2Ja5JUYwVqu0ovhi2GljpD4mN4F78u2Bq7hLj62xfoDCzcGeGoAfsg9JAWX1KHhfxiJ
6VV+cSmRM0mOpxq8FT2O7g6jpACvx3iIQjVQ9BuPPg6eQXXh8G3jU9XnbW0FYqi3UQYvPwsqsKzo
xJCXHx1qDUzrzRoODe+KiaXMF8zXy96/T/lUj4wHVvQNFuZGolmC2zGj+RyVSltY6b4uqQ0mOPA0
en4Mdevi6GM5KnpjDLkzY4DKXGPjl+r2gsiuixyBt7MgDVS5Xvrl6d+K0a52UsfdPqbm9xU/r/KQ
6FLjeVwMH7TL8GIHb0EQsMMNk1NaxtwEATlCh8sDNPc8iH0/K4kkJNzmmm8S2iH1JJOLtKzJ0l/X
xoob4pU4s/fso3nY+ZpwWQPMeT1wi1XX8SwGtCf7HXP5oLpo7ky1Y4Z1BpNpTPvVKyWUzxlznfRH
ry+AYRjnLmjm7fOD2jgcnFfzhUSIiOqiLioy76ea4pzqz400LGdYL7auxioTjFFdxhn0voqO9Bli
Aq0DCqsiRp5SSJLF/KbeU5a8zCqGqEsyqw9EQ3nBMVe8i4VT3elmjPHmKryQI3GaWMF7x/NYRh0I
lop36ipgdUsDR13N03aD+Fr6U3ahHP9Av2f4UNOKUoMS3I7OZU7tH1+xkfYJ56ZNno3lCWiWooHw
RYoDecHi9VizYOoUw1YEOuDagctwW7IvfWyKWUMOEvOifDPd+sfRXS6KC6GxR7zcYqoiu8Oyk55u
hBlEvJN3rAuEYIG4Z5DAp+Q5fGS7K6YRvfDteQ0XDW8IX4Ny/xIoWca+UuEAkP6lB/ZUNQ+I9Ca0
+McI/J2c5i6jzxSmGPzk3pNtVlx6mlkO2CbcfbFrY1WPn8ZxLVwwNvw2YG06SGEKrIaG16rtkTnF
B3sqDklCxyF90ZthhOIG/I4dNfZtDFYifYVdmwhU/IV2k47OTNcS769HXi4H5Y2dOo5LR6ZkUwfE
pcS2RRYMrCyCBY7szGrY9UCeDbyGDOincxIZIFSvieoHSCqIQl+SnC2G/7CW157b/3/8RKbvoI4m
QKBriH8thVcxj4+F1pXa8hHcxqHnot7oo7qU7criYCqTorqj5NqvYjdv5g55w6BZWPgUBluTDEzI
RIdokqmg+gF4BJZPTDMwnTx+wOHKVqhy0NEoKLkGfd7KWt6uUzsr/Z8BmOJszj5ic5SL6YpQ2KpR
KYFmrRAFVRrYEcIiQ4PuNQWLuj1Oa6rt+0XpmDa+X9weEb4ArMqbmCsVqtB0KCIXHl8oYx5lp4M0
j1kDkZ/bp1k3Npk1jCrDJTYv43ZvZue88YJAl5VoB00BdVkdFpYZI6Y/La8V3is16JXQtu63xXbR
DVJgbT97ywHDWsmIsNKNyrWwG7OTfzAF4sbOkuAtIKyb6bgix1xIZBIFlsmtvwapEZfSsRZFzL0C
JQbYODQ2orEPW6M+cvH0P+akuNyfXkLyt/79H9mUd+WaJKO7pCyQ5o6zEMNA4lAmh5bSt/PCjiLe
A0Z8nYV89GOkUgkJNLNteEwNHT7rFnblQHMdKvLS9+4ElMJ9F+fwpnzLhX4WSpOQ+rghzM6cV63n
dLBzyAwq6oxMieP5+OTiWOHGAdR+dKevPsQJiaxgRkt71VRLyKtSArLZt4n+I+409ukrUd2kPPHe
IIQL4M9y/61HWDbOIjcqCH9SUb6pVDybjG6py49QtApN/aM7ssjfUaJ3G/fVYiBEIvg5jPMX31Hn
4kWgghN2CiqC0S01d3jf4XFoy4/ZFV6YAoJtjq2YtbbZxMPJY5yAo9zwZOYdNhuZafs+lSWbY6hr
sfumblV3owBJGZrmkQI7FZdT+wMSAEotSvzGFidKaVJ/mCUXQxaA0KKvLOKBtWonUfYAnxLAkRXD
tRmyMur+Wv519x2OW1wuRD//i53XeOY91rQLmaOMr19UQ3Eq1miapUrF/bq0mQ/RPhMtSQBglf21
YNswU97ilXyG1jAiuav+wmqTAw4PiP3xLjhGMKSc7ZxpSFJI84VaUf/3IUp/Kz498PupdMO3mut5
Nh1UH+0kaezbIxfGXoQoUprczaQi4u7eSYiODP1Z2kAThjapU3jCKhbeGivIgqusxOCuPtOjFPh9
W4MvUTQ6A2CDpOqD3SoDJPJ1tsJZJCHMXEvelTSKTkDs4PBMeS3O8rAhOjncAtny4l6Ml57GI8K0
aJ99brXAZ0/52v1Rpx6e2RwJ2jNHxwhBZhVgL4yXp1TiB2cpTNbpbSxx4qyY8rfmdq9dPzLAzxK1
6/zOcCOzW+/SVkA/kz/eyqt5xNw3Io6QeMQd+mXDKcGDlwG1rWfPz80YQ8Oyci9Za4lbv/Zj3Hkz
RSGYI9+qHxhKvs6BZyG1+KC4kALuHbGBIkPgMJNZqgPCCOgElnV4fbjGJ5RbS7l2+zrJ1oV8FOWZ
Q4mlfbFRcJz+SaQGFBxcJmFoSJPInrKtEefXuTdH6JwSBaKRn+pS38KGPHz676EAAvl4STbOs0BA
vNkxwS6erd4+VVE4YahX5efUyQGIEC5PF8F9eEDCi9pda0yT9GVd50d0GVBauXCG4E4SxLFW1LBF
pdG3v50bheEDw/rgv9437kJubX1uo3xSwio3YDlXQ1JMz59q6WzBMl7R8vOnXByTA9W8oGVXTgdF
SPxTSx0gIbQe7i4eQPx/U1AVerXH5Unp3NwBB8TMWTrPoQHNZVLWAhrDQRDWUF+/eiaGftq/iglp
JzSs4CeUUnMDggpwfBjRJHunoccPXzPfnq3oRMjBAMZa6gBYu2/Gkqh7ANr8eByXuRVVolhLRcmN
lPBmcnGnD1yPMl/QBd/DimuC5v10XiOUM+WwhIof1cMqQkO6lkCV7hSgYk7n3NUX50yt+dbW4Hea
N3nD/sLrcA5IRRe/dPhJcAT8ApJUW3N+Sz8EFwqSnf8uuOhyt+KixYGR+G4taQJrXAKkfy7eawQU
jhhW8OWPFhOB+JcTnzDXr8rgNugLiCBPNWb1bB1eUtR1CWwsof0aMEZOrFfhmRxRIjU+4Hvoqz7N
kFwnoFt2Qw3R9gvzoaYVIO5TLK5p3Mn3U6t/+aomylixNP3KOBOhao3ThzpQwtBA2Ww//g9HLU+x
XchO7vyx+bU643858CMI4g81JnySDFnfXH/tWTPDATqy4wSyt42ty5PGcmRKXBa/cET6Co+LqPar
ASxsoj+Gidw4FVml9HPQ5zei5mU3ExBeEXyzqAHiaySeI6ux+FmaCFYTeVUbt77gYZ3WPAHl4o3/
tRSFeJYKwXn8xPzRy1pPkPVj2FYD8BI73Ob+tx5NeL60OcxNWqMFkhL37F94CL/eDomUZRR7ZR7O
fxIVku3ZUmRv5dEcd+1GUQ9bT3+8heoPrQtmgEbF4s/kQMKsn4q4KU8bJ5L0iuEruRiSf6JAPKMP
3hKAzeBFA9Ekb8jcirvplyeoluKrIlj/fG8+HZ70TYMkq0/48n2eJ2Q/vkTpZQGR9UlK8cD7HIO+
pADZCRweYq+8XAsbD9A1kE/0Mj3Bd/UD0SVmC8jvyEoIiRtDabFn+K6PRXxef3JZz8eMMbyryWuQ
jX92dX7pe14120jYtlRSlhCxEyJr42CsmkHOYlxTdx41CpifUD1iuOY2tEDXS9fP+8i4MEUJxQd3
7nJnhpxG8LbfGgVP2V/M2FJ4+OFj2u4NpkhGoDhWOnDzkBwn07BppOHaeM9h/SfJCYnK+yNf/SdB
efBScnTT0PUygV4lp/FkLo1P4q9AkeFOZ0mzjmhp3i+ttmN5ICjnu8gWlnBNnruejd/yzK+F+4B+
uZQZRioOvnQ32N4IDf2SYlHGOs6BFMkPT1qJinKGYOhXf0qiL2aA5/jg9NmPAAnmJudwco2E+dGN
gR+xi+tAm33gA0/RNfdg863T61VO7wMcZZs7bHVzz9kY1tNmpNXmOmbV8oM3POt8w4QS93TlOLc+
a6DqvveXHmQNuXLxLKY45NeBiIatQNBgL2UNHyIUQ9fT3K4h8Uq0wdyzCpY7Esli1MXw6c3tLQ0c
8wH/phPLXt6VSbvh57gQYASaZWXcj60B+0ThJlKnESpVn9SHa2nw4xkVzo22pZ2z4qbXQNMhaY0M
5YX4pIE4sAiLNP80Obr081miek49Azlln2EpK+dcFEaxGkMETqB3eADebgZDbcnWTgOydSvm6/i+
vkNvfDBeclDBS1loEAOBrP1mh31hnZ+3E2bQe3xx+jPuroUVV614mKBjAfGyVo/xomUf8xAz3q7a
1pn8ZQzjIWB7zKROKcnIwvcZt6TDo4E2mBKGstVyfTVbMTr1y3PtIAuVDiGsV2pjCpKoo1l483MD
0QU3AWungLxAZRQA8kjANNThPOP9oYc2dLgCWI5mN/iDiipeui6xfKtIdhw6PUd10KrzBzDhwaXk
PNaZwf6PC9koqbregdYbFolqex7fFuhVe4W13SRE3IrKaq9i5WRe3XuCyNnrnXKuL/AHHRTxDGTK
fN/MoD44qFE1+NSlHWCSb3xYW6bmYNhFcnSUDAE4tvI8iK55uXl+t2m3aulFCf55SEE582D5oJWT
8407HmiyU0sd7ozG1d9GuBBgoBG8ZumjiWKof0HEb/ypUwjVwT7p5KEEd/4SFjgBSP9c7RvE6Yyt
bKuxjCWJeltMid7oo2CX0ozF52dlXP26MYLXCAoshcAkwmCV8Kb7KUnFmQs4TBV/ctY+XqwGxIk1
mcONfa4Zz396lRAYtt9kCrmv28tyzkXNia8aaT5Gf5oL6tFBLxtX+ebPmLgTWFO0RF2+Vnlymnem
YdTVZBGxJGTy75m28i6/VACOomDVdYRBDIAGNsxAERQCghUx/p5dAU/MkRViJ+isTtz8SzzMBdw0
1uBq2ZjPNZOxJrIhxgyDBAaDSQyXPsTL6GyzDJm/x47EtA0GoweOeBJgfn/4Xj0KqPNInkP3Nps3
Bzw46Vs0QXABOgdWDyy8Cwd1OBE0RaOyPtm+gtd+dNyYP3iQX4UdIxIOb8vq+78+SXxWNTWS2XAb
cvd6Zl3HBDu15BoZ4lvw6BRx2Gs6XpG7Zr+w1R5IGhwX4224Wyxppc/LId54V2OM70bEo7MoG0bK
qARo0FybgfTOVtZs5+DsRPf4FLnbyNT0WkheogHtY86DbiWREB70krtWhIJymYQYATMBq04X7Lka
CnDFwkELOkYkkUQgON9LGaFbkMw5DoP6cZg5Ab/b2QPBNQVAgy/bxKhhS5UbX7A581BryRzzxDy/
30CvSiVIa6penI0W49DMpsH/S6N9BZuUkFteabuhpTGPBeaBWaRb9G+1G03u/l9BRp83ASmZ0E7n
1zofX5zu3W+io3htY8dtk4HjagTtvXreaAb8QCASWOHGeGVBIczRbaXpFIxJqjh0XKKRkveJqxZ7
Tdeu116tFAVjJVoHLhrqI5Sx3VkXhuhZcKofYx6XKyM3aQsacrQfXxxpReBNqnZmb2wTBrm8jCPF
R2ZSee/1+M5cMO6fvIwQepG+VTmm+eIsePQrRRSs115EkDtY2B4WLjjOWQJzyzPerTP3K4Is2P1b
Sa61qDzju0lILe7azrxH0gkiXLp36SHS8jtagMpIBoSeX6n0yXO+JER3X+x79YM4nqnctECAXMAZ
ItgqWAeC7E09yWfa63M332+sOtpjA6YXHxBnB14IQb+kIT4npQZHBX7fA6fzuWlG+WryEyamqQ+t
YBI6uCSKhH6MejMsYX4BT1z5X8Ra+YYyLN1q9V69mroxCtJQ+oTogRpERD+7n3XOTtaSP6ui6efY
9nlo0wBryw+HsXjQOjjLcritIud9kSeAdAVszhOa73nXDTE7APJj7D8IuwYEhDSNHjjnV4xJspdm
P1CTSvhjY2Uq2i+0rNP0l+WJsrMzKt7TNlLukKgVW6S+ck8RLgIuzpSdzHsh/9vvgKjMVLS1kuQS
3qt1HqYV8ONMrYvILRhx+La1rHlZhpKeY6khwZSV3YjjJSwglRESfhH+YGP+ZnoCDQgyudYDamTK
p15/LCXUcE070nrvxXYjlQI08tKyVK7YdCGOLlkXfvHqEM2/g7pabqxWWUMkFfT9FVLukdBPsQtT
VeBmfrYBYQdtgRN0EjBP7Sn4vY5xU5BKg6GtVwLi6Gu+IagYQAB0ecCN2GOQgGbsy/QCa1angdFW
+KLD9J70fQUm8ZKxGPIND6Rkr4274H6S3MnogHROYZmtWhdT2/H6dw86OkKOe2ycUDmQegH0StPO
9prulE0MNyRbce3ghT0/mJS5LVVDmBQ4tFR/cCvIXhka2Lf4fShNJmvuH4y2ONqoG6P2pjfZeyMh
Rc2M01zIOlgDiZLh50ABKh1vfpmxyMnmHFgiYCeEPJ3rTT+NEIDuAJ9vRhxMWVJBEAXZOmO0pzzb
sFXTOCccm8yzrqxv1QJ7wBsysg7aTkKE1w3H4RHfrD9z4m1kqNHlIPWje/uk7ETIaHYWcK4Z8CKH
l9hAnQy5XcSU+lmMehp004uIX+RO0dPWZjEasiqVlP1R/F3cM6PIu4hWLIQWVsesc3H4NZnfBYf1
X1WFMhwW7uSvrGCjuFaspaAy5wCiVkAEwz51YJwLxSjynKlWLMktjUltHVwk3hUKfPDvdGxF6SRG
ms9rLG9ffYzRrIOINCALO+D8oVagTAET+Us5XvnJgenNbRfF/qw+kTi1OubpENDMpzcENghulC4O
J+oDkRb5bQwMjfGmNYTsKmCHeuV7cQHn1bUBi9lXLdZ84Zc7uavrx/V+1BuB7AGJeFFId8bkzbn9
WIxLW7LuNRmMoStAyCr+sxUZeAVQyPiqmjDI7s/KhyTb88uNp4MNqgYek7b3KpqRqiTMXqZSX3bU
Cxk5/IGcDgVq3CFlGkZc1mjt4Q1xYYzGUVFw+8gn92zAhSLQnUvzG9nL4IBqxuuGCuKkul8+jwhT
j8GQGKqYIndYagSumHhGGysMxPBZ1nXUUTDbfdzY1c6LxHEAXHpm1nhAZ9LjgXfu1Aq1nLGiCTLp
wxyKa7Y9dywaWGsTrvK3rkF4BVuqSOoIMtIt+FK915aF/qRoCY55iUfribBW+Kztjq5hiMeP1ZzK
VyVnibLAJHWiOfUGVpWFiOxP8Afx8rhXBKbxRdYnXymydLWT502G301J6tTcVwdrc4gEqDAxvVBU
/GKTw5ruLQM+6hiJROAxy1/9v2r9mT0SP5PG07JpD0et9a+jVvfhZt1a+zeV8kM+VkaYZ5sqz0TY
GoBMDxcE5+mzrwpbR2l/9mcUdRhJl0ViN+DFknecMgGEpf1BrpOw1lXFFm5nWoeQZZQ79rn9gdjt
1wGwHEmQyNJ+fqgcMujybcJo8SdHq54rPQjyk71RvgsIikgMC2Ff3EXggKNjZp5N095mN5fN6LV6
MgVIQIgDc9o5Tu715Q+kCXwWp65wOKD0yKfUk9HUoWMRs6eKpawH4TSHR6qj0p7EAQRTDJBbpyzy
zSveS68MDEwSEx76IRdM3CtOXlb4sh7o4mlLZ164WJJ1bu95dSs3xsE5H2qDIeSGRMr/VW8Q97o0
auTQX/iDxgLLBM5LVoJyLa5gsF8Ki1l05ROKaQhWBTUqqw2QzyOCY1Ay0kcuhLf+MW2ij2VgJVJt
jtRNW2WLJvHOTs4dgkWCidzAqVTiWcN/CThkZzkeVAONZlY9vh3Q9D/EHh02cZglaBxFz5XDHAos
yuR1128RrwnbHujXerotZuZ/hiatLDba7L4ZJvgTZ97znPGEg64C6qj6it4eSYjXJ8wioJx0F6f6
lipAR6boIKgEUN/aaHyeXa95jj2DEy+RA9ClfMm+NbV3BHRrxW/rWymDxIU3k+NoZZ4LGawZ2FBM
PZW3S+6TUsPNbGx2klL2FcZO84tRdh1+586NAR+wcqUZs6AMcYYDDGTBIUATAP2dROqVWdo5GbDo
Z6UIqTaRbTHx1ubriKWPnPBzp4ImUlDkiV3tteH/fvvHG6J5RubpLC8qUuAZ0YGy6OmYgrofbFyf
kTIpljDZ9rGWoFzqq9igol4o3euL2kf1nh6EutM2pyzv5UWYNXABEYe2NiWYLQMJDLsU9+lj9o79
1/3jQ5eTYRhgQ2QDpYIfD5NWtGp70Q7c3K98nBXgou8bEH7cnH2WXUe9x86L9261bxPNX1WnKz0T
+wSi3aHnKUPwD1/gBBhfHMoeXbLqTDmIJiw78ivMX7VNrEqXvvt1xxm0EjUv3f+/4gmyX80VG6Ap
/8lCA0mon4lUvSGf/U2tP5vHAM0caHUmZhV63QnR0MF4WciSmSJvJ0Z8swJLqRJE2ex6CJt5wkWv
vfakptEXws1f5Bx6z8ZLDIVVeL03h5a85IP76Y4c5uI7i4hmNeRVf9oATGrBtAIkJZAvqwErd52m
1z1hFKW6dZXKQOID2YYgoTD91OHyDe0KqPDA+FiWz55ob1KPWVu+st3ema+1zZ90KTaIoY/iN/ZK
dvJBFs5/0STIGHACwUY8a3k0Y0mc3T2Bgl2U0krSDh1zcVv9VGE6EBsqEqZdiWyr/5cHpaX6Q3qP
d3+dEDWAhvwwq66Ux0svHFAONG7hMawx+k3xmWy93ZZZYvIVo6Z2hnsTDu4v1mPndRRobFCa2lVg
LSZJHU0nKD+SJQcasDdbRqdh3JT7NLq6/CMq/oMymF9jie+5JKEi420Ip9iJsN4g08a12N+qKFOe
JsR/KYPwxpIbO1PAjd1gbau6ubk8iw9tqpjBegmP8IbFPcEWpV4JSmW61V7pyR5CAUlrn8mvDbzF
1myw7XXViA0bAEb5vigfjBr6cipZ0rFNVR+pJ57SX8rKffi2hSzVW/aTvBvFUCYG2OhnlF9t2Uvz
BfI4njsSFU6ee8KWDgkRkM8lS+50i8oPt5We2j0ta6LDTxgcXd53Co9EPhYBDPVTRHeinrgpAhS3
2TMm1Kc/PU8ik8c4u6g/DaX8tXjl3pI40ojAerh4k/mXuFprau5wVMt+pJFId9aX2pi9MFEfVXUL
aCbcuVadTzgxWw1YL7a2uudVwdThmE44CFB8KP/bRJrrk42qjTnHwr49m8ZyPc+3tADkSelC7u2A
hLOGfQRginGjtbb3Swn42Y7GSMwtun+dk8WpxMyOhUnYRpIvAU2tBCc0sqlbAdz/wrWsm+SFTnUf
1cvyS8a03J/av8z6wotIDHJHUOwgHSwB0eRjTVNRTVfwKm2Ly1vEEWBG8oI1co0ohQaw4sCeDRVB
JgMmyp/lPrPotOUEcQ8evXLu2gy/GaiYIF9ydp9e1xdfcHZu4nWSqqwg4e7x8UnY8U1sCHmMR3kx
8AAFAk92rex9T2DdnBW7QP4qiZ6r6fNWviyhPbjNgXaSJGF+l2aUTOqJnV82YOIGdT0n5jpivgOb
HDkCXHiOw96zLvO53Z8Bm4KSIJq9a1iMMB3naEaa42v9EBwQ0+bmNFpOEEMev3LRnOZ78zAkkbWk
N9e6tgKwAO8FihA0E9xb1M/08Cme5Vq0G+7gQ6R0g7obOB3Lm0gqYP1y5mebK/tvSg70Dt1b1Y2j
6xPEht5xru87/KYoU3DK7oqSwgHJY8xRlBQ5dh4G0lx4XBTV8P5xMAH1FQYOSmaoIZZ4ZCBv6OQE
Hl7Bqjft0MviJhiZD1gt6sYlLvisPr+TZGgJSqq2hfZhZ7lmWSZIJQ9lMo/Eh3TeDiPDf8vQOWlN
nt+zdTVVCw32hLLRgHy/FvmIvGGMNlZHEhEE7qBI3zXsWAve7p+vJYfDoHoKLlp9YSiT79xhFAOR
KG0VOeGcj/lzRSb5XHDKm0V6jqtFWjbTz6HPxReBqu/Q4axTKFsP/0P/7+xxHymBB8Kvmgpjkka9
K8MkMC8Khmes6TWvXJgdGhN5WaUXXl3Hxvwmh11c3NNkEN1V0amAVpUV1ip12FCBUHSHyj3+1656
g8nXRFtz1fo59Tov2lbMaJxpbhZJMjLlNJOeARN8oAbnHRXOZsc+6l+cjykIQRazi5fGWJ1lrgiC
43osqxttQo0CEFWWxh0ucuoqrGF4pT+aZX5ganqTXDmq1udVFQnhuz9h5ER7g5VPJ0bCrEuvosd3
kY4eVjA7fDqOW2BURiBrRvWzh3dEk9vmYVnn8OTxwJTQz7c0T2do+Xk/GpSLfrllynoQ/44fl9ht
EOWsR1npq1Ye+p4LpzpHFgg9VG7GrESR9H+xTYI6COclkDVK3+oWRHaReE9ZpodRf2m3XKwru49v
v3UalmN7Srj6lwW/92rIxBxWUHQRF2bFf8g/HE3aA33mXekQ8I75Ejy63IUPPwZo1ZqY9qZLPWib
RMfsFf1Hxb3CBSYGDaT+cnJN/wD9IOD+ehD4skX/0RkZamQ5ws2r1vU0Opbp9mDyCXYyr0K2GCjJ
6go+e5Lk2liKj8XWg3iTCYokfyNcakyqjzR1r5PilGM4sseHkr9vxXk5nuQPD0XWDua/ALjrsM+d
iligsEjdBWDzZvjjYOEfGGuM4Pgsg5JGRxsNODSOcar2mpIZD6tCu/7+zbcTD5eTxTGsisblJy+j
NY6w632Rw3j6Bxzn4PqLX/qlgXxcAAgdalnM2hWDruyHJQcYRaLx04Fx256zrYE4tHFpDbEVFKST
TatulQPa1+qTSx38dseYABt0AHx7/APpJpH3KpO+d10z9mWjtI/4/P0cXZJVlyQ+8uqxDylqKv2Y
XCTo5L7nUmJvQtr4xrVjTFT3LuyMzO/YL24R4HDX/HiOO5QYf3hUNxqvDPwMpfjnbggqkJUmkowG
/XP7RJ54MPeaHciety2szHw9lQFK7rVwtqu3eDdw5XfT7JeuHm/0tGPUesh+igIukSt683aDFuxC
vCieW88kLLa8OGFOQfKlnralFqqY/PPGZJaPOe58HAoRhJy0pPdhaVpdf2ZwOTjFkckOHz6SoBz7
PJoSUm7LYXwgGWS/Ij3DMtfhGcqm/rEu3tjQaNfgl/8TakAmwn7BnXOpRjKMBx+Xpmfam2wSHOm4
Qs2qVHIC09CU6mea4sT8x8YdOy0nU6zk8knguUM14zIdJ1w7ey9GlJq1zft/SqZVE/1sik6vyqT8
w7BlRCsLMUngsuQis5O2C3wDN5K5THxVuCsGQsP86lLGv3MhjKxICRjtmD2ul8LYxnX2Y0Ia3GnK
W1bAxPUne1DqAY+3040/xk1D5F1h4xofzHNExUl04AWznIUJHzE9E0JCtI0tdK/lxq0U2AHSHrLo
fjMq0PzfhbnFBZzL7N1HEwH1u/GVEwceDHtoY41YY1ySL6pkWnj8/Dziwjlp8nKLdp6Wikhe/T6r
2ygwaX5KMsy6gIRQgnXaxZv+7qK2yhZJC6OYQZwfK3Uugdx4Z9vK2hYQ54ih5wLa1x1YtiwUOpGD
BITKDP4JVTPaje0r7lyZJ1iQ/L9QSjaqH4lr3yuz1B0YQrZo5pjk3mVh3hrxDxwb0HbM29ogjZLz
R+VqQfEoHtbqBnXwSwwkT6amm3wwe+yj+kpsVr6ZlBAOj2eJ76n7wxBBlMUnnlHkq6eMOsLm0nmX
xoyGX7hQAhqhL4iM968CjIyXF8dv7mSS686iF0mRAcTVjl1tf2xYm9BwqhMupX2g43xOxM5zKJ83
G1JO+Mls8K0RFuA1vjJS9FtaHSP4XBfhWcRINtqOnBDT8bzOtFc6uytCQMKv8LOGhD5JJoo+xjsY
sfMahVthd6k/fF3RjFgTBPm3CtKownL1BD93UjtEAmCJzG39EPPPSDSuqYDLQ++nQXZnL1Qp4kKO
k7V6ZFEvSm2inxspMd6tLXLnUgUpZtnn+qcdkH7CMZ8gGzQuM+LBSIB2iz3QTxcu4ZkyUXNOIQXe
UhqdkmNeUxDHfK3mZoeCSPQsjWJB29oo+D6TvXwePv1k0TBrGuoly40dPxiuLSaKZ6ncC7nnUT/5
Avh8ooqoAWJ7WboOZPj8VpeAzse3V6AFfneXgrnqTQurXrm23j9v9IxUais94qQeu+VjvMVopuNE
BsPxRLbDfHsEOhRXLT25fcX9xdNo9CyTMCIbJ89lxCZwkhcjxEPpUl9xx45RpMna/CRxuvVd0pGn
LmQr7jeGZMnsVUWVead5wrvYPGoe6XNF8jObn7I=
`protect end_protected

