

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XZtM4bLmkglBewlWavfkobXOIMkrnElgJo+k4jE78ykb7oIZp/SGV6Fmfr/ogrusY/kHxxmgAde8
wVKEHfi+cw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qj5OXRmuDbyb7tXOe/IIP9hVzpHdYEdnGFMGPum5TPAz9WJzfNr2HnR7yYGe719tx6wYAvdRlfH7
1KYaZqML4WollrpclochLq72pgPwbtC9iEEWlamVuKdvYSw0+IzNRBHdKqTykxKbBvXaQ7+UOUjw
UnhOWIyi6vA2XCWBMhs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wc/9BtL9LkvfKqZJg7KOk8nPkSL5jxvAGfC0RV814LDUHBZcOVMBTQdouKf45+uYbzuqQuzhrFia
FyTrOU0b+Dpp/D8a4O6aOPezhZlqDF7SuDaIsbNJNkVeEPTzKN3+pib+HJ+07zD5sgOQyBLQtobI
4fQy7ggQ0o0bOrWPzlXO7kD45yraaLu2CaLqYlQzcDjqnvaWtdvg8Q6aRiloz0plB7OdNZ9a1tRM
Nl6v3ocdKRatScwi+YnBgJn5ewXMvGYuuBOXAkUmcc+AFWML9u7RnCLEmrft5oAR19N3inWP9hTR
9sdW8LGJ406SdzZiv/gZpUV5t/AFjTB8Nihgew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RuHNUBMTP+a4VfkYIP3nKug+Q6Ygohn4DcPwrCybnrM/u1NLZNct3nJM51Ftp2uYn4LtBCAEFd4j
J1ykZQnUjNHc8Om8TkpAk8Xoe4lNd9c07VFQ/PdNEPsRZobFbRhtaTn5kYtwFZszGT2+NVjW60i2
zzHWmeNAYn4vMcnLRnc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M1UhZ+OMYDjkT/STr81dVx9PmVVG5A+2IqAmn0405vupx6bbRZIy5mB6w+gLHolhJXN5SjXXAhWo
hTPhhYqRE6WXBSt+aNme9SGwhhYQCQHfdP7l6de6Oriyjp0GyOVTMXW7th225i4gd1/MFzrJY7uC
eTxBA69zF+OCz0UpsBa0iiqA6SmkbUtST66y3rCQ2iRlo3MqgxqTXadwVQPjyKh+YrZv8hSoGQfZ
859BObwRsVOuARh2h2mJuicqAywYo8mWCsE9MJAhCYkJvjGEbdjUCSpq6KjZZuBtdg5UMkBgdSnW
7odTSYiZWcCz00u/B4xtOP+tFTZhOrGrUTKipA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 81744)
`protect data_block
H55iSGIOLuGsbPX2EawsVup66LdTYUN8fFpsycEpf3FjebrKyUHxko6c8SUEk2Hw7/MuBQEIRW37
1NmwTNWRhEp2BZb7RI3taA2DHk6uWt/QXmNCV2iSKVv231nSb3LI4UcEOGWKNXh4I9eCz0jba8bK
lvYfLA9zABG7b/M3x7xVnreNFMGej34Hqir21tWngpb7Cja7SgKfDqufEgNt1ost31cD/AEsMvgj
UZEzurXZyp6wyjIdjbthPpIkNt3fth720/6JNDPhAhHOq7uDloIx9kzy1QsRsN1lBNfIHOgppy+2
HwYzteNQJ1s+F/n1rlqp5ZMvUcyXz+XY5UU5jUfMW41Db5n2NGm4YcCFz5to6iIJWEV39RUQ7tbO
/7TaPl06QsiFUas7/wm7m7ZtTWXGDXQJ5iYAm4u4T/+nRX6oomvFMbq//mjKf6gmTHzxL20XFh/A
1x/gpZti8uVS3Xx7fhMyDthmzhvIeXJyLDgrob1nm0aLbgvWxsNTjyIaH2LQhyw8kIjFs53UqkaX
RQ5yq+Yc8T7/UwjT3Qu2mNylmkVqVEUeVWy3W1QN954+L1+s7dWcuNPfLCW/U4nKVgSSYdo6FFvP
pygiXGibStF4PilJ4z9twAcMKzU6fQyzHaPUrdHL6QXGHwZnzrtasxvZn1wG3ksYSWXd32NBmwAq
tErQ9Tf/iW2xtxAlw+/9hReFXdRJjSP1pBH5sAicvh1GEkQZmT5+AYHymjUhygMJ8uJZ7kSaXnEh
oEuFEwaSeXIm3s9oWuu2WxdrP7pbcuqMIOqmSDNaSym0jdukvTEfylE9IambGB3pJHAjVho2+FE1
P/iqJ7jlgw9pJKmXGQ8PFyQkoq6I7bcL7EKwtE9Ktsyv8skv/c14JsWjrkRNa6VaxKSzD5Juo7re
q+FlJ9Z5CNUyOAbyIern1tO4tBkKuoZvxy4FcYxrTjH+MkxTmZ4J4OqS1gCDsrRIZ9m65Gi7zri8
d09ehKxFaqDTKA5kURMi6kn781kg9xJTFeUVq4iKoz7W1TWgVgWYoXt5Iluuw05jL7yQXJuDJgk4
9gp6Xew+Bmck4VqUKKQru9ky5d2DFROYI03mcUoGaEE2BVa+KYuvgVNHlNOgZaseNFirqHjRb1TF
N/MUBWUzo0x20lKAu7NCmAWQnG7rhNtC9+AjzHALmaTXyzQ6QO+wjbE/71JmbHet1U95H2RJ4yKF
JifcikSMAcB+WH1nWzQFZrI8Mme8xebLJA8ZdgyVtnCYRQGp12zzaqMqHlwi07nfyoOfIFCMCS+/
jzgDWkfFn6LuzaSyipmbuuJ49f296vYuMI1j1lHyGeDvpBlHebKkp4oy+dl5Du02IAjVNlYJsELA
ABi5Bo0X4rHDvhSzkXWC8eP/kxfUdCPXW0h6ScR8pMjNkJcLxVXptLZpvtF22jwJRtMxybldLH+o
zh+jnuyz+T/ErSFYJtodV994PJEg40vxcteGey9vc0RMtO0jOpRvJnXg3t02KVLMEdNoi6ZxFZRB
XcT4enFAtp70g3xNczK/xZUSqwF8Fx2FsmHvuQv9nBz4ff5LTNdQbcWZ1TOVcyFgfiPi4MfUWmmx
v/CmfE/zgG0bVnpWxB04Oyo5nPQxbZIb/GGzRFAL+wDHsVBtcMzP7YVJaUU8Tgb8lIqk0U8Mklzg
OhMdTkbuf0BEX60eHBxGVr7RG/4mREdHS7QikSGhvh4zaSK6imC1uggaYFaOqKm6rFM+wA7hbiFx
FyHitZra3mNWI/Rp2ZlMfVpBZzd/7U2b5NN2xIXN2Ab7uvnSyLCouoqGEzNN/O6CZEWAoH0HGdEK
2RKlbklbmRwxb24MV3siJia8hJAtlsCfY5ApnnqaGANpjotuHzGueROEZoRi5305h/wrQbDNO/qD
NsQ5hAEYqtRDz7tAjmbpGGYx26gN+qTQSe4Ei1S62wl9ExML1HxBGI1y6DwTHVLDQRSp+G6g+PzJ
N8kyjeEFmdl09ipMhXqz3NaawX10e/TcDjMvZuY9MGQ6MiTp/aWRZcOnMOWAL1smi77+NvCACg4c
tqYgDDMvJH1Rkw6N7SlffP6nsvXjGvWUvh6HqsdwoSolWXxGO9Tg7r9+c6ipocarhf1xb+XPcTqX
9hKxGgdaeMuCdyyhi7nPupzxlZ9Yz/mPFmyt7q1t0k53OUFaOP0d9s+5K/k5UcyZcQbSw+BDi9yn
9ToR3Ug/YMzMrdhx+elZZQ87FcB7LR8cGd4zpvIU1A1MPSxY4J+Y8oIN/rkBIxibJxMB2agC6a/Y
svuelZoJHVoDbtnEp6viWPq7YvXJNoUkwH0yWJvJNcHllDZf0ugJ8vyjn3+BryGL5e6uXUlR+PeA
zW1/ht/fnDfwbpDBW9FsWJIIacC4Byo22B3ZBz2sMB3wyrqsKg7cd0ueU8mPPRb5+ysaUQV6jWTj
+sYXfldkD3nf+ThrFk2P8N+9gMUEGrC7k4H7PVbp0xWVKlw/PFKUOsdT/OsmBccJDoUGC5rNnA5+
Ry1/tVmJUwDpmuy9HGpep1ggC5Ga1/wDdI/ejI2kvryabjz5KS/IPyuiL/PyTODvBpOYOJm6A2L3
+5CS4VezgHFLe5V/etrs6sdl6JFnormVu2+/fHbvNXaogWm6QIyIbbegNhMhcUbABuLYbPlfRO+Z
n7IgdtJNNymtWjw15cepVyKvK5MhqF3mHZeB9TXAAArgXe4rPUOzJ84WSoDgIGtuyH/olARWmiam
ZHW9eQpw+E5mTQ9wvH3/1Yk2E3DO91roBXMSgyU8zzII43+QAtVyailm9i/SXIdOEVd6HajPbRUc
IC4d+rm2s/lokcJPrUzibpacBhtURfiaSm1lyeh2x0UkutJpxX7y0sjGY83F6Vq264PxKXQOt5Ta
MgRPmy6ys48hJuI1sqcjyu1Bt+lTtWN3DGudMeD5wnLD2fLSbdXs1+/aVTE/FawZrhO0pz2MMLQB
Inohg8tG9frkzjuQIQ9gs8VAsqL16J6sk4pyNib+ovGs2nZxyvnWPVN57TKSlpWDuLMXH3qsZ65V
IV/P7oymhZuBvIFCXR/EBB3l2LjSgL5DorRoRNYWqf/gGFAC6GTk7WoPAulgAXa+NBze06aJn+Vo
tDQowxdC4E2GujxC1Wra9XwAjCioCskp1x5gi7PaY+x0uf0NlIgDxaUBeDJpHnc+L7Pw4PwpSrNb
sTIEsbsTrIcrLhFxQlmBpsVdlc6xtQq1ynHLqV6KMy4K3phe7BsyNeJ98tnJFpFW5uEMmYJoeh8R
u23yAresXw4ETKqVtxy5LzkxgTLD3Twrj2fFtlxufLEKZxfYEMZJiwK59LKzXVPs96vy77LGu7l1
QOkWk+VOIsfNHqFzVK0O2Ur3mVNH7c8z3TRiVE63lqn2cQhqCiAI4P5JcsJKmHxRHvHG4W/NaWpR
E6uD6Kb1C0pYbrccb6vvbSv2Fn9u70bBqiEHt7J8eu9B5wuWc7wTZcmcTBZCKSalhLy9dPRRzZO4
JLLS1yXGmSlE3Kwz097JB8v0iOjShxqT1ku5c2XLuXW+pc3yGDmMr/bYPKEmIPBlWpOZNhjppplx
ceblK1XrSHFpjESXOacbvmi0Kg4GeG4xBIi5VA9i9rvBSQEOKXj99LtqvVmbS8onjLDcuQ1qxFOu
vD7seO7lLpHxs/WaqEFB+HIla3DrtmrGRyxnYp6THco02BBcc7iFGIJUi7UroCEoTGsH/P7lXCoz
o6o+5+8A4SIk78vbmbr+fdG4piXFGM913SX1TlaWj5gQDseoQNVQZnI41kuDMzMylYf4N16fUQzh
NQMuAB9ZmrdX1xjUZ7BIhxVqIQujAXS20klrlHIKUci9GyYGYXaIcktOBPL9yIUbPj1HoaA7Tm1k
7q/ctj/2eusnkd/FkqSjXeJnf2uoZ+EhutoNpKzYpTtGieSpQrjZSejsDF+5eFWeDjqSIoi/fErN
Ah9GbmCrL/nGLYY0MmD+LubysYeJ16/3QUIN2zNP4eabQgiadp5j4N3BLLPHm8rHHZeyYimbxIlg
R58dyGaFogKE0pETF6PspuDklJENwmnJNU7NzxADDQG7TAG9QEuX9cxuPcKEUEC0MkISAJLsUoXD
hiTtl6O8pJwYDRLSbhN86nFkg8A2ezVZyjataZ3xO+69YpJS1he1ShIizSL3i/NAGELIlseXuGpA
D6lZ8XDAukTY0jkk/cgbcaxuARY2RAkYH0edliUHoJigu89JNhdLO2vnqDyEeZWP4lQkb2C8kNVm
Dw4z/R5xPssjehzEo9foORNShlFaqCPiJ0WpZPGleZjzGGUMmR5lQq993/SNA2VFwHZnVawplqCE
nSFZRQr70tnY04dYEnWUEZ4vhEO+thUkfiAnklHhXTD/NXwCRiUiQR7/hhNv0ZNfsFP7dXz3rzRB
FKMwslDwTzSJab34rw1FRU/yakaPeC37W7uzcAlh0ajY5eMeY0tR96RpSmA4Q0dGV3JGPaJPuVcT
X3LWfJPRNNc4Z/c0VYHEYSLpB349bUtbU+Fk29qBzEqfcNFbYt8IlRjfp/s8CoapAYCOn0hwngzX
Ra7e9cg2mHtWunb3VqF3N9ciYybZsUGNimjwBI6E3zjFXxOzmZKNF3HAoaLF3g4LpH1AeWHAVR6f
0EBFyeUr2Lv7Gq0gSUIReVWZtdnNaZEh+cMlcUzoiZSp5yHhTPjf+63wJJSzQbkjEiHhtTBOoTrX
4yCD9nN8zhp7yT9nIop3RH2xeLNTNMVGOnMmgkTcK6w6cMOsxATWSWVxMWd3yRl1Ly0eMVKQhZ3J
n6J7iWXc55+ULqJGeFnYkoKIddIYKCiYC7qZ/LOu9zV6Md/MjT4iQe9FAt7uRJU9sH/MZkZW0F7q
9Ah0svxDHPu4TePqLtr5MOkHEu2R0wliXDIQfc92Yr+aK/e+yYvaIWmMv2tzdxjdenA9MVoraqDl
vcczrR9YOei0TBwWwg3wOchDZnXbCSDsEOmA1I5gq8FO0bYGy0Kz6PN1jF6klp296AlnwjqxtWza
EwjT7chprHfhe96v72nbCWwYm3yEmqDWwjudOXIFUQ/AzpOcPXOv3EvRoHo+OGO2FDJ/vka4KvOu
mEjyo6fIzPbOP6cazNzO7LdKxSQ1AVGtmoECL0bE86ItJCec2Uk2x5pNQH/CxTH7iiDf/oddoZJK
56nhJ1egnlahN9erH6hcpl0ivo9k8migRNycLq5TvBsXKmqYyg2TY7YGlvTvePV3wLvKzP51KfzB
AJ8C7FjAADMnrNvFVDhx6Ca/RRstDe3VSsumHSvyXXqj/B2gh6Tf/wP2SyE11SiAsPE/0wM5QR7+
hiqiipURUUSZysvYLjIyfA2L81dm3o/B/Rj928jGzhlByM3CWmJ/OVJqmY8KqCWXM7A/YIAKHIjR
JEOzhaLuCnVCI/lEcuJDs0jkt5pUUyX5YdYcJkVb49p3+TgsLrcUpJ8M3NhM669dh24cEi8J9FLX
BbGGBlE/eEX/eyjRA2Zm4rDYU71/wMZb21O0T+nFr1u1H+joehhwGxS2ph1rbcKfFD7pCjdFBChP
zTYO7OVTXPOYMfZ8ApAFPb9t49G3P7E20der9Xef1eS/A2avxTSJDHLAJa/n98qsWCHidEs21pK0
FkvlD1/Yg5vWo4Y9nbmsKF+ll/q2alvO+22H5Yzj3I0NguKjqhInizuZ9Ojy8i9a8HCG7P/kkSqu
Hj4VDqw/ZTbMjQHUS2GH3Haf0F/6TH4XE3jIj4oX08J8m7aNUHZU5bsAXJcL1stO5OB9HsH2X7RQ
5Ifo5Hd3p8l3tvCjdbEkT+4xq07W1IL48tsHPmkuOgozubGWdhqd9ZopuzawqPISrQm4ktACv1Ak
meZpLpEnCuFHgSxO5PXsmCSMTtbxCdEPw9T619rT8bqonnimUCKpEo5qijgaOyqkicNmKm8rGj3o
YNwHsKAViRpfvrkxNLVAigE3UK6ElER5CjHr2F6ipzu2aUa07OGZgbyi0YORpOmX/EwZam4pp4v5
2xsnyn7WqA57A82/MV9VVd6XMkeERKVypGcqJRWSJjPJmdI/0BTjMGwpCu0rm5SmvjaXulWew6Ws
e3+V1eMKypINjSrKE4IUKA2uT7ISazejBSYARNB8xUq/i/dZGcM2hhVM5bPOQ7CnGuYVgpY8gXl+
U43RiOoTDyK7sUllE7ZW7+dUG+D5M5XMkTkyZx7BIA08OTDIw7AzOVZG+nDgXd9fAvTk93NP5Ryq
Y0p+w6PVNBgEek07GqF3Q5HvaL5idI29PXNNlg/xagrbwDNuy5dVjY9MJm8ytCAE1tR2fxG1vw5C
lfPnb7lXRjKG2VqpIu1NbBeliddNQ0QLKlQoXGsXvY47q5zS8R7rCCFGaiL0mHzaQVFpjiDLDN1z
O8Gbwg5VnpCD3HqkdVTpSDcTdJzxMhpwoiER4USuYuk58QN13mytWe/a/r/ik1V6PiBQ4g0RQkFo
IacTYxgi2U6csnPub3CzTovlLz0rL6okYOt+dNm51NUcbrinYkjAyqYGigWtbe5xWVHlW/3L48Fw
0cud4pTfuoMH2qgcamzVr2UOIgRs2y8gRFDY8TMU7Z2f3t2gfx3wEY5nhsAAQo0oXmBwOL1VKKgG
gBGznqymD5/1S6taAtHkn61PXuv7JwAEGRGXy3xY8CBxA4ze+NhIhON9KJRdDOvclIqEDo8+I+7R
2YYcbnKqM769UnbYXd2UHQ87y/PuyVlmO5yQAggHqp+HN7inKFCtg7g7LpzIo/16JqjT2HvxR2MN
cJqk1Bw5WYoSFzmoYLcv+umGJwsI3MmArvvPEiCovVmxiQB/L1nl06uMu8uzIHFTXoOxYALBksuz
yoX0Qio5DdfzmIjnqm/tcT6c01RHXi2SCX4INI+Xg/GpzTwko+INDSU+bdC+6WZFiWAIjHLnZC1p
1zq0jRcudpjPDiU0NUDzYszoA0On2FG0HBcfeNYiXIvOyRp432VGsd3gW7rUTe8oUQ5nXcbxCghS
1vEiau1zUb+K6rk4l5EsJb0UUg6S7pjpZN2CJpamVG5vSIyFcESCC07wNB9di9WoWrdLlyYB/BzN
sSUkIDPgCRj5pWa4Vpy56sYD7mjB50VXpF1tdKq1cTo7eYZiBE534zwK1Oboy6U5wDUROlAxBt+V
0uSixWd+bPl6h885wrdvCSDlUmXCauB+uFRsA+mZlZ2bMwBr0yD/kIn0oiNrvD6n4Dw7DWhKzrII
o64MFVuUYHl2B0XS8tsZVAgMMrJRF8OEzJPHir7qaEE49sv8JD5V1K3M9SG4u+y3xljl9yqNgQUg
L86MX0GvcGp7X9IEfq+Upo4jVoUczZ7aROZKv0dYXSI8t63nUmmgwXiM40a0sL2Cv4Qs+1UhcgwH
utMOxvzv+y/F3+OxQsTiyRx5ftFa8hvbXuJK3IR5fOYQX/Fz5aQjtMrcdo5akz4BOgABr0B4fu0U
72SmUf82U9HzUlRQy9E3hfXd/qP/qLfN67S7JmbPt963XY/VZcQdA9+kpPRU+N7wsaGNdDPUazwG
mcaHwVHN22oEEcGTtckbu3ISRlydGyOmwq9z3wrKB1zlst5aXCAgX6nBlT8+OmSJCv9m0tgtpcZ+
AZ/+PFcAkv5gxpTBHZnPnz84X0Eu8ogtvdhYyGF4zFrTLHoxVY34LBayMqDEmFuj/rJS4KggDYgD
CiePqXlJHmsHRt8LSjX0oYzUL1VF9IFGCIafeDwdP+JZPDtobp1+Ko2pG8sFI1FcT7WOt01wMwqB
VRhdmTYPoRYcM6WJVAmGqsmp6hyS/hAr4LJlre3f01ALHdtcc+G3fFm996KcrxSjpJMiwtFIVvHs
mL0M8p8AHBGlVlrc5z0Qx9KXB2pEeXNU2yXiOGk2YfPQNVVRXkCJlMnmlOUgNKHUFutzzQIZLVFP
BHoSGqnNsRSCXdhk4A6cbTf00AixKqPZOQpga6fYyaHrRz91Flgm3fZ06hexqzZD+VhZBjq781N1
sONlnx7WuuYwhPCwtLH94PzAiCmaf47hHJmxUEIOmcQgkZ7eemZmBa6h7niFAc0Y+uu/8wHq/8ia
gQnB4NzvHd5ALaHYQ/3gR3PD2atXdLf6rhzwxTXgY4DTtSWV3fiGVaVrbpue0zT/m+/rptIH/+zO
eLFHCg8yGJTazzA8QYys7U0KocdkWho86vOF3211cAVeOQFYAEykXu8sbQ2NNHmu8r+29QqpcBH3
lfsKad+dwjibTr/CTY4CuXsWftmEen6qgYXUNffDYhE+uxq0zYpOtJ0AhFtOGs+WGa5JgQaQ2AeT
LxeIZ0n92L7015F1j6wx0sMW20lAomWDYpCbhxLmOXqmok7nEnKBN5722VaGA1FxNV+Fbbnfg6q1
bkJV8pbyiAHoZ88QUnn9KistzcrriVbK8ozt13EIUJrXcm1RaId7b3trZkG6Tj1EKL4s1tdn5HLm
kEqdteLS8moXqBAfuRFt8ErG4Im1vkcpfvce6eDtF2L+Mq7/xbE97k14ZACI+2lYS0KElZOP640/
c8Et+NWYoYe+NtUp4T/wB8y4v2cho6aC/BiHEWvLv1BFK2tEWX2HGC53GRHKcvkABkOxTDCfWoAI
dwKnbinzeSlfbuAN1o+rqr5827cBTIUXggm+Pu8RonFz4QmenCwTHXEWWcyEpthmrpqM/d305nu3
H3pPLLTyzUpKStY9anEtyJMB2TUFgPL0lJVZiUNnDV6ILgQ+txFxeIzNyZk83mJKKTtsQ9QjRitH
VQLLhCcnJBTcZRhfep2caQuxGs4nnRDhdw2phEhiS1bWcVvZuEezrBQglYCvZRrr1zjFIS59E/8U
owPnBBXM3ukjgQccu46YaYWFXdlaxJLvx6gOqcfMGyRaH/0cPEJQTDSsw/qxkbD/TNdoqXblcbkQ
0hWMduc2IOgmxMlwVXDxirEUUtJWsiMtYsnE0d9hEUtrA+NBE9vAKbzD3DPtGD6jtRL75eBpP8E7
3WDtWCQCqb0ipA+I9TicyXccwKwGCqKnrZQYaS5t62ENP9PokelcdiMQL6ig+8dSH/wVtykwagCr
GcUYGRnLB7q4ma9FejSOqtSmPYTdcLavWI3k0La6xrd16u4revDrnraceiT6A2ivd1R5dm+bYiiR
FfJ2oAK/AGdAFHgQk63GoGV6k5dL3sR5vUapGdwSYuP4WNKFs22psgvGRSC2p1KIRQBEoF/2F/rq
X/LnYdmbAiSzS1FFAo4nF5peTWLOZgTG8gnmptPpyaneoOaMN9LaVuJ9BcAHpTatcapQrDC2AxpV
tbsgKM5iMvflfpBK/7hV2SmYQRjO/OcyjXa1vy+mbH1rAoxf/me6cxi9FvT22++Iqe2lCkysK1d2
zv0l1XX2eEKiFQl/60ReglP56t3hy8ZBxcFOuh84F1gjHI6bvgaSuSIJYDhlnEObEEph7qtfGV4O
lIKHPiWVUX42YaiRMDd2zjYZuTQtSpO3R+6BxZ26w6Cme3Gf45oRz0DicggxCZWQU0kmpblJlhML
Lrq5yD43P+oZVlyvaykMO0OHhMy9+DN2i3w2hryp9kTWep0H9h55ZVSZJna0A49cPg0EcpSWnsF8
Qy/xnZI3i00io77Pi28ZylzhpuQ/d4XAHoNsGPgpBQ6iCydxn8x+0MqvVSdJHeGKmeSBBzEmNLZl
RYpiMOZ5bmOmKAQkwPu8s4LefqOLVzRgoHjhDYxDK57UjgGqaeXPD6xZdr+i/WusHY2kiGJPOz0Z
hMtZsO90i9v6wEFVO5sGw42zHMWHk7GFJzQ9vXm66AU2eNpmvj7VxE4atKpvSoBvIVQOnhsq6OZc
9Gf7SYxFFzWNdK8G+oxtRGZEUVU6QgnrtcDGqqp3ush1otB2urXXPKKhD5VUklA+7qCs5VDMTfl3
+1hWExPstT3WH2WyzjkJZhlL+oHkukZ2p70vV1/PTpudH7/GiTzg2mvb7u5xK23+IK+WAJOYOWT5
x/rYZqxoOZJ22qFu+O77EQTcZnsBWIjymHSBiKwt4acK86HSBgbpMo3AeiMjjet1uGZW9Ms9/Acx
lZ7IjGkBoSVre6S7rqkil2wBk6OqDWXAdjFZOM7KoYDazKUR363akAc09FqcqY1O9CwnAHQkYL33
FzqkiQUjmE9YF4GVPBB0/dsPaa7sfV1dItfLPO5Ufc6JWzD9Uc9f7ZuiyRrxGm/pZ7qHLvistGAb
XutSJQ1rJWgp5ltkO0OIpvnxDyqx0BXru2XQc9aO2KJfohA0pnLBCJiP16JpjJ/A4tWzPnmaxZsi
dxd/CAflUDZ85Giza//kEbOfrCf0l4VpCX5FleiY28f6rJoATu+/1AKbDJPI9FayfmmhG3GXvB8l
uNibga756+npa0QhOF7Yiacjrw9YcvJSoQYtmHmqCwcJOSzNM3NqZ/4LH8Us1r0hammgZ3cHsJRv
Tf+MgwjNIRmdEfaPVrExs8F38hRUMzXfv99QoRrgVP5ntjonc5+vq7ZVe6eJNDgwG9CSflqyWjQw
WEwfCgdv9OxbVdMDyAVeE1f06wHTOOiejcpT6sEv9FTKlVVtBIymdjedXrHj5Yips0rggolEwMu6
EQs78r84GK1IMKoL9W9ZGLCTgoLcuKAoErAHt9dH192YtUPaho6fVBnLLpR4XEsbd5OPJrK3WRG1
NvWcpV+/XHuHThqNTnAWtYmM7gwvW5lmsvLlVYpz/x2xXwYf3q7SZiAuwIMY5HUU+8SRW6pDHEGd
Ft4ndQm5ndPt0eLVCAEXpifpO/4lFHomTdmEUbqVfg38nXQq2+IQ5QNLGyTr2k/vOuesQhk2dkix
LlYRjmjwct5VCuEqEXO9eFlD5OVfWaOmoWmnBWUZx9Tjb9XQjGy7mk9U8XsRe5+yCUPD3Am9G+Un
EKa8DC0e9kuyRiOESTTR+IbYS0s82ofx2nvobhLvnVRL3YFFSsyLexdJ1xfozwxpIBr7NFG1XJt7
CmKPEGUbtplJXfpHv47taPsZloTIeCzHK4wUzGqLGiRNVG6KEnUSGSlXqiJQTEIW3Dh92obvJCBM
jWEosf6JSsIbP5p+3KF+Ge8y6TnF5cPUVlWVQw1dBbpwUMtq8RhMvtD05mjAjspm+rMhr/NgJRmV
pDHQD34TF6nqn00idjxqLqqRP1GICoo6fyiPLNCE+JgQzTEYZeJabPzsTkXj3FPpIgn/2bYuQY/I
zaGtSKeW1pZhAeQ+VeL84qMKPS4MvJHVTBS6mnWiPn4IB1gI8nUOV3R6rp33kD4nD/7RxLuXLMXl
0XxCp4HZZMz53XXZbc/INReNOgv5ctbTOmyXUIqnJGyKvFhY+4DkkcqiBi18h5e56NUAF3RFNTLj
nYs4/MsSau2uagS06WrHGerjrk2WDS4Z8sWLu/pK0oV7Y4xlhad4FVvJtAfMFmn4im21ym8V1wQX
T8tf9x8OeoFjbeCE2oMLLrl+VJjNHUI9C/FPs0cZuVzwiPQ65Ndt96OCZYtxTwF0mMHGTCyB8pAY
Xk0OThIn4XqWyKpVJhdRUP4HnijeWFIuhZftWN6NeKFkugv6npB4X4zcuZqDopNjzzdhNkotMfb8
5lp3BOKOYmCECQB4CT7pkEvOMHb4XkbBIFByscgFXNh3+JEQNkuJR84CnytOZMQw74xmxU73cgLc
3gpJtuIz656t1pqTnpOEwBVScSFHPYnulLU7HX3gemakmJ5Oj7JvoGvpAiFeGBWFMnFWayB1Ku/7
IFAkiKK2yepKXDCUYeSXQiSjfzMStNIhFUoVqWKD8iMgHXAvh5g6cv2NhZsq2H3EW1hihlRCpLhE
J6K8R2u3U3DOwnqlQbTlipgV5ntR6wbmOqNhVutscywN/Se5jZuvxhXBJVdgYP4UWd6GAWek2lfW
kdPF92c8+C/DK6B3hhOX7QYQKsMDbNnPsK2ofj92yjTUO2GQjjTLUYyG5S0iIW7sp4Y9N3R8KaF5
Tl6DdNGvPrEuAKbvPvZbBLogn61InwpOvYiOmk7iF3KPCDDqEwZDG4loWoCXKcOBW5AX6ddgQZ7o
PdWMWf2aSnGBiK7kPytesxc0usZE1vRe8h8HY0XDHJUYacDbpV7nVmWWcUQp2enWVtgrtAfHb2vf
TUlooAQ4gWkMkfqoK49q51z/ja+ucZtxggp+A7p97wwTU9mkVQe3LL31+bOzVZjIm2gcHJr8d3Su
C3xWYeDyEiBzs0U8gnZEkt8SKdUozUHhmvNS3Hw8ePLBYNv0bIAXzpk7gVsBkdqA1eycO0Y8LmIu
9l+xR1sU+e8Vimdy/UKj31Mnj7vrbLu1mfJep83II9ptbaIFfpvJN8UuPImRztIUYFEb87va1CbP
Tj0RpvvinlNTMFclygeI+UECpkms0sFFKTrlNqbv1K4rOSOxEqP4n205lxo0R7yIYa8ONKzl/goS
xCS5/33DU10V25Ov5ND5or1cfJzVzbQgjKOVoWdl6v3iKmTkTPh8Z6Y/wZ0pkIHjhHuyFfcA+s5l
pcK0BCv4/UtpI1kXVwUyc+Owl/p7XwQgeq2fWHpq8u1Q6TU7vVyXW9GCIwx4vh6yWEcWu2vbJLC6
yyIsHwJurfBWyJvo1/si/9P+BeZCsmALRh4VLW4GKl6Akk+eKRkxXNgGxpFQ9BjptpiOAma0loKo
1IL3eYz1zuHrmE6pCd+DtbXtIkpvj/HIerKiC/VuIAXPhaflYRbSkM47jQCEx/jA8lSAoMZeW9oq
fI1Hp9VgF/2IAJI2eyqPLrf5lbULnG9Ur0bMxxM8UPgGj6PzwaSNWA9co1chS+tA3Q1fExr4PFsu
1x5+BLr6xzo7TsM3Fj5v+qV/o28n5PaIonSBi91LVAe+/j0IWrNmS2tXqLbtsholS89bIK4j/gec
jbWIjB8Zw1rgOMyycAJdF8ofxhimSD1tLLDmtQ0Q1yUWr1jh9ZNtclVzkTbjISzscQ5pBGvtW1IU
XGR1UXa+OAHr7lxTJIv9iCsH1Hzv5hpenWGibHf15qyTKeK9nNdvdo3oCK/RLBpvUaIJ4Fk8Fq9z
mbmBPr2w3BkPFFQuRAw/lcCtA7y0UKwVe71wFt+G1v37ZzthpmE2BqZ8eixl/x7ZiuhX4CQyQxbV
6lDHDoqazRffoqZJOI4p6SzkpTGE5rcVnTqhLvWxnMPpi/boL0qEbkyLlZ+ZND4JkwhzFqhFUuQh
A+TCCbjC+fMOHe1vFtCr7GDBWr3LRZRLHFhXXpLeZkIK2hCe8SJ1dgOI/us2uVDHpmon8VT3qTC9
Rc05sr/fiS4wxRJCkYWT0+wqugYmu37DlTTBk3SksNZZv1uik/dGbHBCxC7EJVICWoLuopqZJvPQ
6fcPTWQDB0FyciD6ZOtA6bSYOHNK2JgRi7xiL9Hd2EfRcm9HtdphcpThwg1aDjl/wzCPE83jnZ3L
Opx4T9UpDLU/dPpwQmkoRzgemG9epte/5+V7tqIKkqAotUOxFMU+uO7GpEPQk96oHdLthuo7ThQd
a1v9XkznwU+Z/8Wu4OLBh17HPvCPe2qA2r1LjTTJBRNSSU8NAcvPsqpjVv3t1I96TIznqgvB4Wqc
mZ+3jLfdCuSMvzvl+oi8adPT2SAvG+058MHwWDRYoWH6zp5UIA86tSoSqA3pTKrqsseo1waNhxO9
73GL37YqndNsHHIFI9ITQVsAYDAs0xViDv7XsxWBkAfx+cuHpSgz7JLe8y1U8GMYKJK/bHNUQYtq
Z/t21Ei+DxFR/Aj3yxnIOq6oyQwUrtT2wTt5aybqYP086ocW944tDN5CLhk+X8Yr3v7OUXYLh07L
dDmpF9YaPqxDipUp4OVSAdEEnYk07r4pvtNr/V8F6CUP0G8eI+RdzbJK4VVjyn6/rdPtp56hLNSq
waDExMmLeiXBAUtCFTbyQk6eZRLfWTlObvdu0ZhLXfm9pr7cfXsv6HbivUT1D+ak4nw4in3AWC2M
AlbrSVLBvGIMR1JkOCPn/rUHUoD/LEZbz+FP+HqPcpF+xYA0FjkfDtGI/BnSD+dowbFrqCsWHnxT
BiWsDcfpkgPc3c6Ws8Ez1bBoHNHGAqc8G2+xNAfZMgyfKC9goT7RRATi8j7Y1b5R30OShqSo/84u
wFUFh7b8ppnENRpyS7c9j91aVllHlTe5uuNonKuJ7MePEqFT1O9NprXkUJVo7kX8gd3NosiOymzc
js6sinjRqsOwP6wxc7OP4LYY9Xnljb5ng4FhRfM5yItkkcKm1Y4cw0rE4NCPAhBsqjn5/yKTmW5s
b+/EYFZ1+tAyAbk4yqOp+pYMyEtSc8oZ2pl6v/ri2Dt7VNJZe/y4c8TUr21/eEWK0+GasVyUukBs
fEBqTJH1oincbldfW9Yz2yHZNWtxfkBvMZTfg3RmaEOhuvA/T4t6UJPCRvp6w2Jhw+5GVd2mcGWc
m2GqfoKuBcqAFKycP+4FeQi2VYUyi8HJ8ZHMZlQqgr1OMEZAhgUcWGoQEqdJVxre08vFoUblG10O
jhxvXL4GFkJM1WuBCG7ofE0RH+ayAUumfkh6lAV6Ts5cYFAHGlO6grTw28ly0XE083t2QuUJLXp2
79Rpz3DmRT5bH9K3cxroUns6Xd+Xi70pm/dpTDzzBP3s1V/mkbUV4I9iDXirerWiP6aHxgP63VfA
NoqN5phIMNktQ0MXkRlikDp65GKYVNkaCl8446UfnUQvKNYsmJ537vItyfltyRyfJQWiowkUHu54
JELpM2O/jX+VAFAV1H5Cm718UXoRUXymXKnA4TlXh/dlJqJIJjlena2PWztl9quMrPeuwJSliACA
lUkkgc4c7NVHq+YOKlSSgTAUDViqo44JuqBzA/FGdyA4UOqQYQa9ihge+RSuP1ihXkA0XGJtEFNP
cBNITIbFlGo1n68ZrFgu5NkPn34/5/fiRKiBV/c5dnvnrdit6sF89m+oh2SdtuypUFZyTR/WY7II
VLwEcSJCw6o/tjtFTziGln443KxXnck08ELP0knwXLDQzbzBVVbwhbWkbABAVFJ+ARGxMvMwk8QE
HPc4rw/N3KSAHkF0Dd0J2mbjoKAoyKafWaF0jjFvpXOJvji/L1xoDkCReCKtUaC3hMYCpH0s9Lxp
0Aw9LYiNUYQHkeQ+P3OgtdH7YdhsjlowY5y22tVljnhU0El0Sbzb/CBofp/eZv2dOn4ZWZDSnzIi
FlwENPVJjL5FnJhlZQwDMRqNL4nRIMX5/QSL7Zf1ZL9Enl9Ezd6J3qtDCI5708U3CyVFvGnKe7Y1
sDGDTR5zpgHyEbPIA9eg+Ur5cBpzgzGPT4CQy3uNUOEwHok96hUZZQf9DQ5fBZcHPLVO0Ct+ae8T
WuXzhaviYVSFpqaITijutgdnrN635c2Xt3tdBxQZ9LCHY0VZnUmbchCJ4YwXfNUutnDf3m0H8PUX
BLJgC4aUw9Nj7YBJFe4y/4PPETRvevEuvca9dMxDnrB8lyLojeI3xayrCmMIgCWamfzR5xCtN4m6
xlmElE8/qoyCIP8u4DGqnFDbNX8qjbH3fSUPRhtrqVBdIEAJJs5OUDjDscc92Gp9ymJ4thdwDwUl
iEVyrbIoxqNWg3FeA1E22nOoJFJgYcmDAp1ifn6W8q+3bK3UQsVqSoR5mR4N8JMc2UXfEEUCID3g
QdH7iKRAHnvx+3MI4P1qPxYVJetn8qrw/Tje9jL8ODAEOQUiOC1Rft5sfnW6SKkJdqexpWeDTwnq
M7IryJ5Hd0Xr4aik3MTTSDwWWFM4ZcqaydZatp0iG1FhQtoYayaDb+0a1SixFudEiKy7J3shf94i
uhge4qTQPNwkIlZ4p4s4rdPPuI+7K/4Vuz7trPam8qUNmhZ+0ndRhHSunf3eYB3horGSwKaaSgEl
M9tZBuS2G/S0KdXrjm9RJWEzjra6b5l0+DQa4cnkKhyI6q0rbn9N5iZac1IbHcc4UYcL4amfTrD6
PpFJQxo0GHzfyYZ1z/hos9KfdPm5uhJzFJ5yF1J+eu+C+BYjyTqIoYeCHXgKJzs8lhN4CumSJiuH
fF/rlXNrwrFQXxdAsIW9WKLHb8xEzRvns46FVji6sGfmYuozbYT2hwPfMNgWsIk/GCGnqe2CAQ6p
7Lyecwr9whrbCXVVXx6z43+TyeoDU7dBtVPYy7FlmW+hpfeXIk05vVZS56UH7Rv5ar+WSW8UfcWD
57SYHe//bt5Xp0feyMnf/O5hdFy+FxorHBIc4TDbbZeZxvNjJ78so0GqYqnk6ofsRdx6slWmfh1d
PNvBp7YHIcPu21WTXpxPxlfsdVPuZjJ4OiUHIjG4N13XEuWQ+3+yFW0R30+W6suUhrJMSTs1im2d
/47c0gxO8TI1Anyam8yBZU9vWGbNl8OxTRyb46ywzRMQ//LdQ69rSJuoUEiCl0g9OXDmLwCYYWOc
0+IRuD8NEOSuKMWAfvCcFHWciplJK/gaVS4O1ZNsKdY25VniSs0cvOUO1q93MCt+AxvzpHaaRqfn
ZnAY7d2Jwht7GC7mYausNWzquu7uZ4zNzCG0Dyux7loah0+hPkE7z1+akOG0pydmcX9GOV0cfwEO
kLPWu9z8uI4fTDncjpvGAgrRMEPGOFLDxJnmvm/eD0PGnELIV8qhI9rwbAcsRRZj/ZWJpMVH3Jaa
0bB4zKvJbjTmOyOzcxjP4WtNBqkEgJ7C342xoeli6CBQ1YqZ8UEU2AQ7Um4NyRAu22FkKkcNKbQy
uefYVJIJSyBY89ik9JBCaLFp5opFhT37pyWcd0y96GfkLa6JM5Mn0bfe/6lCDEO//zOgJhmdZr6J
6KrgNXFfswxCtlFjr97H5KMN+e5dDceur2oSo4wJdiqVtFJpRdhaDKheE/xVXx+h+NeskVmnGUF8
xHGHStN8C0r/owE1SbMAcz3++8KwNDt6QY4WUq8v5QvfVNzV7L+QVkV/X2i5TQc5CqSm3euawr5l
L29YC8Er4fzb75DIiPI+IZGhvjiOu5LIXfB0rcgaTU4pIWMbbcEf2RFq/eP2eqpderdFluzl2ReO
G9k6q7h8oJV2DrHfkUj088jxMg3KaUAbcHN6P6Li9mHu8HFK3baMMGW8uc0R8FrzUwiK0hcnur8O
WAWOBY4heC2aqijZeSDrTLnWeDQmoI0wbf62rJ4ai3ZBhzZnG3kibfkYuGHE7qPMG5W2PQC3V4nO
X15SuoXuzRl1znzPcxWW9wjZv3R8KAitIpD+Sc+Gatx75ucSOlb43s+MsL64lXBVf3bUC/91D/H0
XmkAdAXFx7Wz+vWXOyztf6Y4SvADy2BIuAqNp0ztaHGpqXHIElO73t3cGvUFqDuSaiffHms2Xjez
QQ6pXCntNCRz8pvQ8JUNqyRl2vKhRpuEe6PrLVZ4VIP3EYu30mmEIGhNPOLozpolVvzsNLU5APPV
0AHQJPhOHI6NfKMo6ua9i389W2ZIZ+hdQRfXpAuenRVV1BeLo8zxRkpdBlEBa4dgqXPkNf8TUruO
8tztOQzuVrwKDNJJUl4nTpvfLsCdhZBxdsAejbL1yOAG53Ey2bDgYxD3MOTyBt3F6D8WK+VZ4BPf
iW09UwBcP6kAhbvE6/8U3GIouhIuDdzMVDb2EPo1wObe3UjOoYALroEfR1C7So0Ea7+7d0TI2IJb
SRa61afpngUSuykRKw7vAD2C+tf3bBj+gGFqi9C3mjVEwFYrqKrMDfnH53TZSmUKE9C2MZLJXkAr
bzUV5+YI6N6niFITzaDn9infwuotWSWnZzlbTYEwbleYbh5DtzK+uVgB+Ajs7xIg2hYgQOU5PYWY
O6mqrtUX5yb8eUhm1EldFuYmoL7CMWIAxkZArpzwASxKvULMXbIh9uZXwQ3/1PFs2YCpgBNZbrDE
ZAnrsg0S03/G4/rYZhJcTJ9RZFmY+5OPy+2NPmeHj9asdW5CDEXN9Lk9sq99Rc+ZGI5vpOUijeGm
OT1GD2KveNG1Xnlne2VYsqb47KUkcGa5xpYGYvj+AZ9HggMGdzQnP05YzHCilO5BvCrqDKEOY4n3
KlFpO49qO0ckULA2o2gQT5u99rvLtifFDX1YkII/HRQVwXuloYzUEpNv5kc3QhVR0/2zlxEXHgKO
AMsvfH7ZbsfCZwnvkHL8hhxzAgqiZ5sO+1RMzbHOyiA6zVut64CP0qfp2WqSUJwUAOFBtsvvON3E
wFQMYccSCfYpIUkTFcNkLTkYdpnYxrxH9VGhcuhuPLpbg5UOMKmLdh9r5oZfBTRKc5L3ecqUdxqS
nYdiixwfTK/vhjaa941JUs2NYpp5M3oLMxISrwYdKKNzuELV7/pOLM230rE4fbQ3eCwSpaoRRdU9
b4ZWeR/wVuLyYr4jlav4ytZyDzuwsvKdNa3Nc6g+Gg95uOSWxG4nts37wc/e2ih6BcmXkeHf+ja2
kSY7XvTxogTcLOESj+bDZY32QaUOUqEiQuMEkWHWv1QLr+BRfV8zexgyAXBOsUrlTAVgwAifRTDT
A9oTEJDGLhjKUwvhgTIcUBRpEebFzqA+Gg585TtOuf8WGJkKAUsDI1W6emsTMDVOWHwEVpmkdlpa
RhaX33ZggL3i2meuCs1NonwZfQ7sPmyUHZ2fxNtWCLlt7slahQTW3pdIRQpcfrzlPusJ2BTqN062
I8Q5GV53kUm2CzBEnCc4wScXsh1eH59op3u28vDU+cXzrHj1u43D9AinNNo/1cIQ+Xspjfn1FMg/
MH9tPFwmn5xR4EJehOGziFoO98sw/Yg8LI49c6AsKLXBvg5uENKxwVW2/4F3v4PbpCtWSHvyKAJ1
sEux7pPZk8Bgv655L2L2+d25J8s+hbfP8BBaTr5YO9rijO1fQUAT6NtuhSRrWS61wH/eeSGRf3nN
0087Pt77tC7kzYy+Q5hDnOOHFDyhLBzx0+s5bB3iJKICzzYuWrQRAH6gLB1HweaoEU9DE9dtFhPf
CLYSvkk1Olp8NggIb0ln/FRdq8zx6fIQcJGp0qh6ylqQrgWz298gTR4JqqBtjZa/7GITgmwLxE6W
qrgGuTv96k7tYF/u9JXYSqJA735m2Z4EH+PLUfDvXY9nx84O/y/6BrYMlpamJknHVy9CES0Ly+o2
xtmzbQVH48xrJjnB8GJxJuQEEI0Y49Gl9n5fylL/WfiSY8DIaGhARgsI60y//4xm4l464hgBcDpq
rkqgcnm+VIfoIxa08RcJ2NQylCSt60ioJN0QaGJGLR8tSa+oz2OJuDge3D/JbeUpLHlkwfRasK9O
pVfAi8+SCmfLwN5f4sjUYf45XD4fAHDwS8AUHOGaEt0XzrTnjLN0aUKDT1bQ9qPe1pKlcWicKZSZ
h9tfw0vEXEfR1sTNFi6IPPL6MFbT86jEGo/Kv7FGM/mQAS/Rbn8yHuOpkQdK8QZOTcbv/Fk4Djhb
69fVWCko6O4SVXoRkil9BSRBjfRNq+nhiUhLVq0mJvEG7s7XzGVVbmt037UF+YrSYFeyVLOd0u82
Gms1tgFIbzqgFjBYxhzUaie+n7y5068KXi6cmAieSjFeytLBPTGoZ5/PzrVXJxpzut6jSbwUbwMQ
Bswo1pSWt1+tbUbmOPsm8ipIofocySPKjD3TpiV/RyEdLO8BqKuD+wYip8Ii41l/Mcp8tm9Fkdte
lapH4Vc9qqSp8CjRM0AjHu/VXrbWM1jLGkXpZ1+HKSR0A/HGWVU5ZKl04GvAW2DtTDl/rjIKnKlv
txm2bV8r9PcY26zIYdO8yIleHbAglP50jyIT/PmpZwydbGp/kX7JA0+jfK7eko1bE7MGJVIh/Qst
aLS0GOaUC2l5yZNtw41BJjX+x+cl9/HA1zoEgdefTnp219B61hKrBBl5x9d37xGpqpItt/aSpYcy
97px1gUiwDgACHb4KPPtl86mJZcQKc6mZMHPARSGfNs+aG3tZl5gTl6yBdBeaTUvg8l1Zot0CRc+
/VOARa92LfljTb03eSZWzoSwn+S7JtVQ9wn1Q5nbQvnHxa1/uZefchNZtzYlA3mgW0Ex2b7TjjHl
MVETN/gYYCJ0qeH4U7OGOMz4NJFEDhfYQ8KKW4LeYamemGrkvb54xhjRA6VXAh2gr68Fn++ZjYT+
55dRtX2m2HXeRbaUbYGWLMw7EBQPK9XsmduPi/TSed4JhlxihT/Uht8O9BvrofNdyNY8peTcXtWJ
Jyn4UULuAvklxtuid7JXdlXbLt5QNTjawM39CGma3F2lA8c54M/vkpC1qHhTb5FHcdQgWZCgJyhc
hApRp7OSmGOTKl39JVLc9kffLSY9sqtQFIqnmnzd4N5m99x/J/xglSkApjNpvV5Hi9zw42LjuWMQ
s44H//qeWtzteSVyPwXfhA3bdbwEp9nKN96n9TXQE+iiOyCxtejAb1TofTXfsYYIh/FZSECh5HLi
I753kzW4KErLrrkGxbx/9EQRY3DjtBN93bKIXRuvDljCu9vEx9TJJcPNPzoZ3rtGo2yAMR5FTE5d
K9n7XD1uFDo0vVvo/LEVWEzBcfdUNIR35aBZ88AxIPs3upHRs+vSdaIkQKvliUzmStJRQH7iq6Uc
67cPb7bz40HibFZiwfpgEv3xWzEZJEYjDqqYmFpnQvsR4nLd948DcdaSss1ZxxvAK0tIP3uqTkmi
0oD6eQdzE29r0caSCRzUE9H/e+KaIhULv9BVC3xCYA7pvVHJVGbxwjQXqAdSND1vqJQThPrQznMg
jeHh723Pt1bLkbXSIdo7aRM5GPuvw+6XOw0cHYRUVvfflxCkcOdIpQ3/Wj91SlU1od1hsFIuG7iZ
RRrVUSC3wcfTbcaBmmcBJgikiAE+wLNRUzseh/e9JNjjOJ8TG4xu8GOMIlHr7P5wjfXldCckqcOF
2YM9w1sxGxNNRSnWW5UrNeyIzw94TCc4lAb1DEqRfT3777LjetWaqgocetG0vzpzR7rzLSFlVa0+
od2N7qxQk+r2bYrOrpmTZamYYpbw3x5yBSuyoAd7CDn6XKc3kjEkU/G/YwVxMwsdeW3uNVl1Bezk
KqIHs70ltGfSzfJBbXm1KUi9f2qPMEHBS4heTqrooPr2VopEVdE2N3bo4SpCV2MH5mUUNhFYP3ab
hx3z5KmgZb8/MnM0gdEV76qFdw8fF5M3ofZaZ2UGYv2f8E0pqB01IrB/fRGiIjR/VvyCLJ+gW7a7
c4XmfpKx2lduHY2Q3vsd18Lipxm75j4pc8MCdBnRlN/ifXW1odro+tQjlCreGdPfiT1YI+Qo78Xq
sO1lPq+aXT3piJPZ8/hc/8RjYFvKHJ7KXTXHszpfgEwNNNkWhVjznsG6RaoAntdwQZ8t2RaXuX/W
Q8dS/dsMmGj9wCx5zXVFA+r9zOcT+hOoJMDSIw1YqidCqJs6WVrnPtpzrxCeovcRJrIyWme1gx3+
57Sj+2/vNZYhQlCduC31J2WHcwsGex8qfUCwX/frjWcS4OdVwsiNC8smD0TNQxAhwI3wnMWQ5vwM
eY6MjtTlvFBzSQvdgnClFC1iFh/tHrm0JPQdH+43vipNdRqANYfNqQ9j/nwIctD2GS5fouoeVmFC
3zy4CMZMh+PdxVl8yq/d+5qRYKWmz+izQ7f+IS0KUPcQ8qmGCN0lMOKL0YvPM+L2piVK46AV4Wdc
bUsc7tcSTUlOjYOcsMTnRGKoi2V+gJw49M0sL+sZjnNh/bwVX5PjZuAYN6XHEOcuHRgNP4Bh/mI8
UcDJhSGIiV0Bm83fYqEc+wQK9fn5KxT5EFxL3GtoCmCj6BNO80fOziQx2QEbGvg7nfnAEVbBIrSv
+fRnTIYd5kBBY8gvvi6SEFMrqRqjuG8tqK5gpzwb2Fnm9f8w8qAra5vMBX5VNf334vKHc/RVWiG2
UM0d1kIXvLxeXW21dz4FlG1dZsAK3XCZDLDLvl11E3x/57+Il/iRc0cU+cmzsvWliPpbAQ2pgNYx
53hvJ8TNgzOtjOCl7q7iqEOcJ8l1qUrEN2JKOHCPMOnKuxqiJyzw0QC7FlepEoqEqD7blmrOKm/p
lOu6Rmji8VtPbIrurBObZxh07wxDMfP1WR9tmqxTHo2bNnQn2xBGrAhrwt8yTtoFcXN4kIvn8MGQ
+pUQbsNV4VXzpptUeEArf2o7T0cBgpYXX5XPkePOVPDB690RubggWnet4tsqsvx3bt51kqZpr847
n7eXfMvCUiAS+c+DpMwSu56ToS0Dh9So6SdsdkfSTf9eujpY3B0Pgrw53uoRr5gId4yWA/xEKNpd
IGpAnF3H4aGh8owt/5qNVqTTTzt7OFKMno6+bQs86SGWyr3eTepQEIatEggaLZiTivIK8TBq4j+4
ZX113ZgItZjlLkzbAMZSJsDMkfkVWJFFL9oOq/gQikIFiy2vD2H4+Dd92UE41oRCXfLkFRNcE8Yr
1Uieyit0E4saimu3X9UruOHPhKZNHhdlRndeoz7KDy6NjJe458BFcb4ggogeKtxA5URZoXvchkpn
kwDHjlvevZLaCqBXusMEYRL1LHEWPTE++ZRURfRTm49WSW21KQMvaNmnXxoDiV8TSYBJdCfGfntg
KPiDcr5WVtxdfmXeijylt6DCh3BBKWBPy24uXurklUhc6OA0GXBM4zCXS0lKwaDMtcjoCIsC3gqq
pGvIAqNo2+WJq2keKgwSXSk71F4AdYSS8Y0eGrrQvqYWz+4UUnBTOZqyJH/XsszxHSZa42AnyLrQ
s/p2f3jZAudhWN2eTq2YNpxfmJHl7m9sdOMpuTO32y2b9coKplgNkHnY+aDGbxwjmwnAtZ9DPj64
Ko1dshySVWM8EU0XflX5R7dnhdBefAVD910SyEtDpqcmIPkL/wp2bDOmInErxGmNSWT1h5MWdcGe
K7ZG7GVjoaWNttcArk0iFYnRyqF4KQT8251QAbmBUV3Bn64jfz6N1aiHSZHndBEYq+r9sWil2eeb
bqcxVx07ggekdRExtFMBbbkRshMy8iscUDPJELa/Eu3LZ4yzAArGZju3MEf3JBaX1IC2mDq4irJj
43DzmOrx63DuZEpzvNvXmqUPOH8L6ygE0381R1jkdDa5FIGzVhl9HRuQw/7fbFt7+qaPCd23I0VM
Tt70sTw6fChGUD25xe4Sr9qouFOrT0AbZ3xcZgKOC21HhMRHFagovDIMt+ciS5RL0ovDzBwagt+R
0zTIzNzjBfdKmpB5mO5fcDbXepJaQhN2RKS6OY3kxmYsCcUX6Vst04jBI0aAUwCQxRlmIlSfVHTj
Z8hoSqKHUmdVlqe/QS+2ztkSHojLQWVbSqR3EV33AaYQKxIVFX9BHzBT2NIeJgFlXpbcy1IhX7XQ
LU/x/BZPow4boyFHSwR216dFFBejxpvK9lo5HY8kKtM3TtADgPmKJpYRASOP+0XBIFJXh00xB1rF
K9pNf7+XQavSxPyNL6griL9oPB9tA9Oe6pPeVIDztrHnHHIV1+JsYUtItiLtH9SHmbRAxXy458jU
ML2zuIiFrUchXosmiBxshaCLdRWDublcK5oNs379eee9t4qT8qlY2t7aPKNLAf2YHpmL2ENPspz1
OnuxdqhlC1Zu47KZE8FnLl1wgqIqKVBsX8CRCBbLxsVihhapwHpZne96jvhDYCe01q5HCGog1z5Q
TCEkibugEFDC2mB9XNeMiaWuFyNwL3JZ2juGYm5uRPrEYq+14ynjO/PVoyewZ6Ps36b1ISAkdwVG
O42q3cW3jvILkQnY3uHqx3SsQDxge3HgeiC1qx4zlTW6F6FsaLh6eLdn3CCGfEWNAEtAUWNLpko7
EcpLbDHJjNF8IJtvV4PX6YQWvBsvoXC5ovgV+iRJrMC2ulV42QqTUAinAbQzULKW1qe8e2Ion9ql
6MKWvdOUf/ArltUjYppNXFGRJlUSiuQKYWZBURlFvQ5rfUE3+3YrDO+898rGKT3OilhfZ1vLBd/m
UIlAeivv5WT15nIBSDZQ7+k8hgWmJI90I+RAMWimm4hnfEAEv+BAMmaDWl1r85sdey85QP7OjOpz
JjZDkJivkIIPKwZ2rcl56cLMOX3Xp9zRPtvDi8nQqqhMOR5fF3VX8bGj7YbAbsiepN4YiNozhLpK
xdDQBVBXYXvbNe49okThvrsXZ84P+iMdYXEdmfX3P/XT56pT5jKP3X+f5VImPECMAZuD0M0rASEM
hJ2HKHVCLNV0TKB1ArDMY/wULMW4kGg1wHQJTP/Qbx/AeA/ByGxJyHQZ81XNZzvmgz+q6SvkLDs0
iBIqmi59QNCL5dLJHN/aog+EsEjD6BgxF95CABqf1hDJnGwsac3tiOESeG/qhRe5Q1dtl+IhgWtq
qvt6wwwcZnnABCABbfgLSHpjC3ymyPFvdhH3TGE7iIrTcAtofnfPzfo0dD3gqdW5BOQ1Um4Rkv0Y
FbAkKsZWzQszUtMooWR5f6S5i0waB9alUis/i1AiVjSAtIExeOq9rLAeyTdUsBzxg3IxPOs4J/vi
NAfAeq6kYq2cbPTc45cbJl5ZaAHWszdhDgewdkXC+dLk3JIrHsaJY2VE8Sdx836M5G+l0suXBF2p
a7KNuW1yC1/vtG/PO/4i7cnPPvlI8kSCUCOekVJWo7AlwrDdoR1da7wQCKGIv9vLo+N4ObAh6NUT
8Trm2guQj/GEc8DG6F8oag+7iBUwxMlKYitKi0wP+Q4dxVInHM8D0vxcpiS18ftHO9IikKAr4c0+
lvSmaqPilG1Z6f43cz92Lo7v/lopfF17jBYv7sz0OE/8zVbgv0i4C89ozoA8rCXoSe/i4pftBODH
19hGdlcih7fbQAmplacKP5fhMSrnfx7v/DQ6q5uXN8xNwL0I8/TgY8S5OIYkhiVMYlec5GzuemQP
BpGwNL2n6PKaPzzoA5AT6x8yPg8+rZ/7kku2Io6svNjqS7cztR4voKNyW5hElBqtK3dVsbjAh8yf
pi+n5IvWUDdsCowpGw3M5PlmdPLWqi36OR/DQQFFuKP6SZq+QpX/pTbM2b64x74LwvlftEBdjACA
BZ+lG59l4kKC1C7QwPMnOTr4BMQ056/RDKozYuMUF6vd0g2jY+rpzgu9YX7jv3jFRlFAXM+J9+so
Qat5fGEqbyxrSNlrz8dYIEdv0nBpp8JDnQrXoLvNJFq7Eqaer+kMOIBRE4PzJJqTB3V58Na4V1tS
bDUKPOCbydgvMrfkciWlazp0mvj+k5WrrHkFoZFmGwhOAPCNi5rPOrVKm8p4FkTOuTINH38yq8A4
ln/1vN+VBZfPkqMFmLQTmL4Fen1B6qKCVCZx5uA6Pd0ZaC3vWzvmkX3fB8b/FbnjcTwrH73FwSj1
KXBt9ISxDUgIPHuA1NYblY95N8kSf4FsBbTU2CI5i1dpG9pBbpal/l9x6tW/xF00F00kwx2Y4hG+
cEHj+AXRGAFhYn6m/AU9MNB4JOZI9Cak7/QMaJeh58+y0fzYXWVdzZL3wfyfpeY5db760a7LLKTs
8OjalXlaQAlLfUGaycgwqbJc3ByD7B1YU7h6vOZe9hBUXpbu5DWO7QOt+USb8rXWVR+zl60Xhv6+
fSJ6Vgkg+rRuxDoJ3cDVnBRRRoKb7BFP9AwPdZnH8G9B+Q1HIHLp5ThAnU/EQa76w0JDNl1k77G0
kmTIwNwjUPUJUUMN1OPWli9Ificj4vFtiwh7bN+zwQBwwjIXW8ZzfeH9ONhtTOxnDLwzX533U2Ru
RS5WKQMl3y1AvdNGwYJfPxs1tUBhoA1vN/SCceSASww5joO77SSoCsYTbPcf1J10aQ7EviK2r4in
NcPpngjLMYleCcLNNWRabY8L+jUhvvUy7k7RIep+au77Vd6lLyakR+Ae7wwKn4DQLzF58oqVy8d3
AD3+/xm8Q9Y5iBCiK5QBownX/5cREZk4oqpBEcM8PjZiokwcw3iYjiyAPsWos35RXjL1olLwKgW2
tRKLD6lnQXcwnqC8oCkRKyWmAotvqBFdLDgD1iqTgEZZL3aCcQAKUp6gQTnvXCo60QjwZn+4aeNp
eP4kFLat29a+6b2bQtPc2BfjTw7fBlbm51znTj42O9gqqzUPAKhkbxzg7Nek18HcQfh057uYQbrZ
aZksRNlKh1CPxIG8yR217gE3TTbyjgvjYIS8QKJC1vcFfqvLfU0eZZcXaNAxW8t6GIHNOjJtkfo1
re7NW5sTNhILMtykYfR3LBXkpEC1+iVjCoix9dkxFPezRTNg7LQCmmTEWKGCgwJo7rCeOPR1S2qp
Ig3ASUSuEjF6U4Y4IYztDXV5MpqJ5whGfppmKamsi/G/WLctWkJ9IGIMikb9jWBiEjdSfcGpnm/g
G2pUF55dxmwaZyW2L78AtdinmWnnlg36yYYSknJd2bk08a9Lh6Rbas/tide8PqwU3CFUAq00DipG
vB2ZujkBvxI826d5cnI5dljtTbZea09WE0wuYPL0D+T0umqC0vK6w29kq+y0cwjvmoPijxb/Bb2L
Fpe+Vphg1fhlDJFCVasdkQtMMnqWmSVgfVd99bmOBDDxfB7WsR5/6pk+WOuQUoqiRFcfBBZdaU3V
IF1SMAiH3lEJe5cxA9mOyA7hrqj7vw5JfYXGUA2Y95xEyMdupkO5KeYdCye93CDdx7HKz3nJ1t+k
+vqin0QcRlRldvHxBT5N2bSlMs4ME9v3kWroXug6KP1UOlW0zwS7m2pP8stpPQjT1hbqHqgXaUtu
INn866zmTzBfKXuRVY03ewsm4fM5JCbO0CJENBMUZKGp3TJeTNRGZZ+DAZVoP/9OX6maNDSZigDt
P4naCETMAKc9nzhPzZiWkkYpsFFC+xh7W9QxxGNEuPrtfE8XV9Lu/xTOdvx+r8DmgY/zpYb0OfXz
+R6H81+h94DVTDjpOk0Mqk1V//kSzZ8rq1/9PeiDAYyJTQJr5ItbIB0sixDlRGJMGf99OYO2DDdD
7GYcFZFVInHdLgrgBNp8M5aec8tNzuTERfT99zMtpQv72iKhLCZb1B2pdCQPzMBcOlPMkdi73ATd
RdsYrx7hd/LuxQ5DcK8gUSuw37G3YS1ilS+XkGj/oIKJcSoaS0RaVEycblNubqX6W6Vn9K5ZfVHv
zUw6FmWPX4IV0jKIT6Y8XGoW0ICCRKKmtmt6wRHQds6nWzjK45YrzwePgTkQESuEbPvet5vqOmuC
NmW4Nmdo3gQrnTWx3+EzqyBoAVGVa378pyVAGqkrnc9xr4gBBHOlNQT4qcwhwV4Sihxj9NBNDIH6
dXHYHRdborxW/1sibWWRF5qyzRox0geeUx8xHcVYTuvbS/OyxmTHLNij0p+92Pg5cLVhCLaWyhY0
gozUCfzB034JWkvB/o8L6MzI1GnvCQP5yLLGZyhixkQxnJebanaH5VzumRoQZo9EaPYs6jTlyWdK
DqFrpXJoM1VzyCI/84OEQNPpEgwylP8lIpDsNGw1KSzHJiaEcCttBoPdbgi13Z2PIGh0t2ftlFMp
050avolxlsw58PLtKshTG8dQgeoTLODJjTCSapDFE4nQNl+3yTUDaoxYhJVidnpdgDmsauRfr6KK
7nywj4Q6kFW6BB374EuHUe75aMqmeXDJ3sz02JfBpLMV2xdwts9qmMYbKz/1TcYK2o2TsEFJ0hif
dV76HlkI45lY43PgVFur1lrk9oBG6wekn1jRshLDI7sajGhH0743Ysf10NWLl2+3bWVrpvHc5peJ
HWfhrLaBNhCcLx2UAJxB9YiVIj1GzNWwzHVyQKlzXG8P909UzRUDVpy5029dWtJyt8UepAe90fwX
wSfC3Rshmg50jBGNdHlr/LA9qAg+Kepe3ORYHbi74AzCbljtDti0ykmbPt3YYwzo2k6qUHE7nJkj
PaMyBrTjIxD8dCmas2zVWCRitlZeA7n4kKZYz5xt0hwda/0VfBlsjkTwIuhqe7qaDmZ/lJ9ferYE
8Lo2LpTTrlE/KwkFksJQ1qWeOcRVmq2uhQWWUGVxDv5fIawB9233ZhZlCkL99lyeYoXlu5aUFYYR
olCcNxHi1yR9Rl36bhF7CrW5JoVeVF+tOmQD+3eZZmk2/a2xEL5pEW+uehR4Vn855ZJPdC0nSazZ
hsMpi9QdIfpkPGVxlp7f5qUSxw3nJ7TOZCqm+gyWET2cm33oiSx6qy3zReEwtH5LXprtLu92P+N3
04yOcNvtgCB3vVM/Nzxy8lWjwamBpo7xKTcTl37oj/YgyVy5IlJWVE1v1kV4ly1AK2bcgwp9Zdal
aSG68+CAsb+DOYidkyYQbtF7/RElEjgSx1ibVp/ORfY4Ne57RAK4eRoZBMTUkfjhIvrm1+rITgvp
mJWlbMN0alGuMzGpoO2oMKnF6ws8cqBbPobi+p5vcAt9WDolWEfa/i0QAYKDZ9SFUDeZrpDB3d24
EJ5uGhse+fuPKgUrxAT5m2P7QTTI1KPYLlDTn+iy71+jRzL430bDTniSc1NaeLZLfsmD4rCZaRmb
SXQNeptPqw34PcECLII3R1fmTVa/ZgdWtDE7s97fjyeAAiCR1sBBM6X8Zh7dPVnwQPmecn8j0cHj
2Ws4S2+pAjKBXAkLNXba2EWXOkIz1MlsgUAD//7FbvRTTgA1SQ/uE3q1rvlbS9k0fZ/qit7tXjVU
T5rzkFcXwrhYb0Z9sCHtgs28he7Kqq37T89mqvjIlcydYk8777RoYgnGCilsQNpmjHBR2lt2s+PR
MI4Cs5AfToZZzs+s9uuZrOpvx7W+bfPx2NGYk0orKXwO+PE8nzDXjwUe2uoh2S55KkUcq8Qqry8W
QbyeYFRRpX7uqY4wtG2rw7L6+Zk+7U1FbYQ6wzuZqKPGe5DF/thsjstIIZ7SEQdnyN4dJaGZJd6n
e2CfI53tBuJEuRv/a5IROFwWo+a8QZKDzRQb6c06uzS+ERdNhq0Og64hcoo/C3QF+hNVJCXsbDN5
8HpRAehxrekDh8zfeXv3v7YSu6p3xnB9tufe6MA0wM3DsF3YSUCJvGTyDoOQoSyKN9adD7Vmtn3I
9CI8NwLTBc938WRM4ML6TJyI+UX11rxRfGmehbAbAK5HR5gUT6TkIU6A1PMJQqVtmM/zGnoan765
64Qaq4MPuKkH7uad8qH+X7RXdC5LcyKKQTR2pedkufbkSHoXeSlyy0T4EQiL1TalmXc3ZN/AuwGy
rtTBkR9aqTtK/EVLp3zKWd08U9Yel0wxyLPwzhC+FidCQvDLT18G48aTDSKT2TTmin37rq5/r0Wh
I4dWWxdJD5hUF+6c3UuJ/BKtqscQbsNOmfKD57md4i9a7t7NywNfFvXfHOLhWm7I9YK5T24q6mOY
AuEtk87Wv4MUkHFxNGdhPcWF+uoG000V4PG+szHr7C6DjM3QqN0boFfxpxidUv+3DfaPlJLjx+Th
blUM2hJ76I2tT8v1s2i/DYGBBdZh/mWyS0pk4OnCql4nndApqtIPc/7j3CFwChQoaOC8fxw996BI
LZywV+pH/pJMfA6BQWrUwqEzvswmW64ar/etQHvQGkerb6+czlyzAafEAmde2vgHIQiWIKViMdwQ
FdMtIDLvPrtHfVrFIkmuOzCXTJxSgMr3mmyhNyzVNXUoXJT5gIerS+I8v8FbLrKfkvX+vn/1N7Dm
nvLzFmb0EolCbXxc6kPrKf6pNpyeCvquF/Uq0KnC5fGFbjtfksR54q+iZ06OLhcXidG0km3DvLwO
clUHI26LeR9rE/q/1EPTtNjfAJ6LfKYBxgSdWeXtH4WnjYieGQVYT70D/yEoKQ+ZosBhafiWLbTM
Y3IguaW3fZIIglse6yUDNYC6rJ+OfSy8jodbsDZkhElOd2DDd9S5dMsKlcOxwohZEx67YsEAI+bU
OfZ13spbtTP3PgsLdxcTB1DPEm3stWE8fmDzofXZr/7KP6iest2xGZdCL0+pQsBQU5uWtIiCmDvF
CrRYraLGH0kojiwBkev4UhR8IBryqUq2fZrBY0UulS/UUvNsMaExz6QlHPg3cxvqvfpq3C5gbP1D
OMDw60PZGX5sM03BKa18YhYYlR8UKiITmggYWygtWL6ZSQUXiEd0IqOveGOBryXkRAO/+vp3RQ1w
AleL2/6Jw62DiS53BQTysjEABjXrfgFUScKg/mNKIshgBOeAfQIVHpDhT93n9CHPH/QDzTNyOH43
caFWJxhymHWSrIowSnlNk3W5t9x+dCTwlDH0sgNT1EdX6Tff9hKSzOX4N8n5c5WjexWohxdgVhdo
NIa/sAUKvdtT/+akR0/5XTnngUK743dDNSwNE8SCt9OprTYXPHCT/Ea3Tjg75JE58BsoAXcBsefC
plpgvGqZigBx9GCXhuNKOTvQ32DODjrLCQbEVJdY2UYJSlnSgghvjhYuLcCQHVqoPXLnW8ovSGEo
ByUYJgxGSaoou21cnEF7vp9utAFjNUTIOAZH9IW603dxeRVqKCua1Ilc/vQrImJM2ZNeRGeFjFEL
LJv3UbRqABsgNcrhqf8Yui5ayVulOhr2zGmSZWyRuVJFK77286Rx3X0os26gAgQWzpTbNQyPfXd5
xDJHpJd0bN+S6MYnxh8PiswkamO5Hdoh5IqWLQrIlphgTcBnUwlNX0bPUw/N6uABQ7tCUlnJu+Rw
lBc/WHahFsNLEU5GU5qLTxqTPwlSW7Fz+4JhiRJwhuy2pza6C9K2EVeN7iU3HwJkSPJ1Ysoxqeul
ZqSgxT1jOFj8VXpyUqPCKxbA+dyb3Ty0RxRJO+Tmt0FcdwqYd5a/nGx9KNMu4SGccnGRCgDAJHaG
K5qg+rFwYUrAjjtu5vWF2L78Cj2P68ogDRTGEISLbFZLLVdjlz6m77UcYgwmEPfvFQVoyY4NQGNh
MNDeK2eXzYsj6De9C2E2wI82Vf6GmwGp+3Oan5M7O+stxX2gdXfRt3Y4wovnqkRXAKKf/kJFIKeb
aqI6lgMZtVZ8d6tlzBWLn8ja5jQ+uv5/Z0MSiekivWSzhpL1mxnf+OPfygfXe4msxQNHWkJ9jqzr
tCdKQIzmWljs+az1IbLT57ZwWT7QNJ8KfviSbmaB9kh2WCFaaTGvYamsTZI/LK2NNVjBEszm8KEO
MeFpKzlP/mOwWedb4NTpjaIb0LXnTaVpDFeRI/Qk+BzsLcOcGvRdxN7UHowZxzUbAAaOy8aMYl/t
iMNYFOC3sk78/6WMNFI2NPnXkZL/QlzIwSuEZAFPHZ6qxj+ZxvMhIIRkH0YVsS4bHdOt9zmXpdRe
SrATNwxhGfJQ3/Q7vAMZBzwYPJyWKjTIpo/rzJFdyi6w1aTpitVpENBb/3Drca0LAsIe6+zf6Q+/
O6IIlDedFZ+3w3/X4mtVIm67Bnas+U2p3piAXU19Nk/OvXdytYmNvz2EVjJnpvp2fEm9KqSQ3O4m
x67eHBIzL48KFKbZ4/dNGrrbHvQi4QwiYelTu96DVs/cvhod8VSMf9qIFInqe04g+ecSnBt28e0j
NQSk6ya/KTvEI+z2KmL96WRU3PAYLfR6PJrXVb4FCdsZ7mG2ycxCqhRJvTL+KvmntWiRTsbxbEzY
pZZMfDGverXlcOoAb4+BnTbXkKAAFPpCKapBUDDqTWj1eYklbzrZcj+51UPrVhsm0muDW9ndBGQN
HyJAn/dvRNu7z4088HkvwvqjtgG/T6t+WWpeKVsTn/VqIm5mpDSWtWtSKNFmtTxsxPYHInuZP/L+
5uFWMZ0cCLXWtET9Cj0wMMEDCwHBH4ACBSR7uw6kNrAoefjrdFvz5MYv5Suef1DUWmInI4hoLmtg
vzVRwFTcnRMy1B5Lcty6iJi0zU9Itt/2KCRbnEIIeOixnAX2I+cGPARLKIaZ+jmA+xzbgCvqrhm7
n2N0zZMuYpjnEvd/1A1l+chIZSC3GCdD3nW2R7cLRyJAufQMmHZFDGK+h81+Y5lpDgzrZue6S2qc
M2f9VVUri4cXruFFRmRqU8/5WqYX2h85qNDZcXeZx0SbFxzW2oraOYo6AhOrD+H+ejt1IdGXiLbN
OYsGFI0HP1IZ7ZHB7ZWgq3MQj2N9oKkQGKKFn+CrepIhn6H41XqHsUjCHEa5Wgav7ZbzqhOwSyuw
gSVYuAzr0Xqd4OK5pgIK6Bh5s4OVEsa/PdycSEqrWs7QJn9RL9EM6ckD4lomF2AZWRRdhTZDrBsY
iFDH8q4u/QPQ0+qzt9TwmCG0LmM+nmjNEoEAwYuyuumdcOD8F8EQjEvm5HoErM5HMBY2o4Ja7tMK
nlgYDFHhYVU+LQHs3lrbuI3MaCqNTXT0JC8cupTVMWaAANO/RmRBepSTcfo/09nu2KNMHETbfNzf
YjaJY6xIku2BMIGuj9aNjBM+G8DHakhJQoDv4O4pJhk5x2akwvLiR5egEmZXt1xd1Al0wTWXnkKS
XJR4jRkyYakf4YcD5FXYgTrHx8l0IMA8vSwBjJSYSIe40lox4IKQWWaGSup144qtw0U1QVDHGFd3
r+1Xk7WFkwSnoxcN6vw07/yimHXk3u2py6vUEbDWGByiGmuWoMr8rL1sC2rJzPLahX1WDtAWtqky
Wxodq3C/DMaRqrfoTnG/e663Es00LnUGJGTHse8T89bxwABRUKjf7csh+rsyJqe3AK2AP6add+IM
aiUWNdE078hrZBvR49B1t4vdaPklcOn4ID1cOvo8fc5Ral3CdsM1xRQ87k5w+j39tQRdP76upeQ8
L3BDjjW94H/wwYRX9o6K9pBazLtwkSqigr9iK0gQl5DYEXnlHYfIbSrCvaC7BZ6Szn24Oit489gL
udsca0swZSf6K6zGGEYYPZj82nga1QgWItC71x6CRkdkWfg+3gcyPASo6drsy8FQZ2BEERIQGhiF
toMEjofzRk8JSNyJvp9BvFy3OCUToZP/1hYCzFD4LfVFDbjy3lm5ipJufaP8iBBabfqZfX4YLs0+
5jPIdELiWR6zu+yZpSkFA8mrd9mk9wCIOdv4K7ufIruO7gIET+d7R7EoD0cYSWOCVGcppXqWZ203
7bnWoV6BC4L+EJZxPJ+22RkQjI+nj9gjTHg98rJiTmRZx8EQtsSlfCoKRG3lF8OC22plGhsVMSs4
3h8VA02AqSYG1zDpmq6AGLgDtULEKLfzJ1IbdCR1CzyQStz+BhZxHvFeAAVP3WMlxBWiDyYGcJ3W
zh6p9svIbLshsU4lcfE71O1avLzyhT/P3o4fnsJU8hPY9WT/fSo4speCLlBc+nJbpjUJ4F/gEEuo
HnEOl4xdLDcww48IRMWhr33RaFSLuHuk91DfjQ+1ycZSYWwFF43mbIUJwK8/02NCFvb9RhQ1Lnzx
65lGLVL1dnvcbl/daRJ3m2AI52yHLV379xu7vspEk70g2WNZELKOIVpjgGz3bvcSD6NcmEkKpp9i
XERCvDkPqieX7R8iLpa/TH+Lr2i9B72iJReyL6Unp/yY8j6HEtGXeOxoKMUycRGDwOdTzKBMhsdM
wUKFiK9He1t1MVzJL8m6qsNH/nsBgBPJcOgV9Qj/zM0xZtevGXtmQTdMNc3OjmEJlC8YVWTeFVhP
mfhnAVSZMdmT2RYnaEcHtqd9ELqVkiEIM2BXCc1IvZ9Q5XY2lra2jhZUpcSvIBH7c54HrjJg9oRz
E6uFS5wC8fTq4iIos6nbmFhY/20k0s9cj3PFaS+HNjbKALkehC4SLINCG9SDq+eGtQFJ4XiJ2oOt
3K2QpbDbw8eiOvnJkCuIFGr0TVQe1qMgMP0juSm62pQEy7DKloOHYSlBiFdDgVU3XVDU//z0xby+
LhIl4vYU4ZFmtrRB8FyGVYbjPxHVebV4n5YwUbmPFhCews8xGP0SL3hN19TRPX9xyANXffe7suds
h6iUXcwe56HziYokdthdIZEOleP8hnF5e5ZII5mReElaUmvm5H80MbvV6WEq8reaHGSv4bQgw+Hh
oKGEfg9+YP743T9hkY3rF6fvObUIjuThHlh7iCTQPsFUUVGsJkmShFEwy2DjA5ovE58q6fGEGmgH
Js+0jl+7j5BUrd1VLw3+ia0mL4r4Um/rzhGP1mCIymnnDVjVwemvT5Zf7HKXk5nNHGWCYspOVAKX
vV8lJDfjNOE/qJ6o2sve3hAXGITaZSNxd8iwBS2YFgcUKpVPI8iFN6NLml3B0RlcLxoWMyxAtJRk
V4UTQp8nDPIKe30Rxhz6ZOL2KyV4+Uz7RPOOqyKmvbUQn0h92+gzuNVLH7ErWEkYDvRiH7y40161
fxrSBefOk3U+wzaCFdRdRPHwq1BG3DZ9Kug2gJqORDIzDQd75XZxSeD7bMYQqrHkIIDHiAF1Aw/y
5DFArOJ6d/UzrPTy2AXHg2x8kVYcDdVxB8MlQIF3HDpfXWp7b+hoZl1S4Qyr3vZzAg3MjAHJG8x2
9o+IuGNz68tcO1B1aCesqcukNbVVKg8HH/yb6I+JU24GLVv7T8DOLbObTpIbRVQoyfAXjXzepI/q
dMjc5Sdjlp4Xq6v8BFamOR3lDVD+VmzCe32NP2AmXvk168FeVnO+faU07COTY7e3cEcnt3qoCefZ
GLMIK0pErgIb6Eck49URM80evbReyePcNxZXxZ1J5z9qo7a1jSZJSVfAnxlBcxm6aGKNmFgFsCBX
Y8ELHNg6D/FwZCpkxd8sNcMMDrAX4HL4r890mfPQiG41tQe/eGO3voToZuzY8dgZwS4nOtIctOQH
f/EO5O200NPtcaT4U8jS1Gyu1BNdR+LQbpzAy2E9TOlgb0lAHDlB8vIalEOcATx7RiOmCChGJwiY
CiWIjC4g0vvOfbUpQEugcV39VIroTJOiQiEz/Ij1TlWzkQ1ONOX8oNrDctiZrhzRH5H+12eMY3BE
MfjNxTcH/ZHNbblrZk7rL8zeijpFzJ511IrpaJpRth1VfujghBfC1BKkUYObWuExlFo/MtxGu2QJ
42cQUhQKnJaRMLFA+WklPxREdt+mlIKTnfmQXulQ/cbVqI3Uuwog1gMnSVDnZc7nXrby7vuLf321
UPRSJCiqdse3SEr264Z3jipNiTtkJJ9OuzPsnphPAnEdPt8CQhoZFrZJxE7z40ZzSNtxW5N9bGy0
02xG5WrMvHZVu6d0md66UpMS05DPzUUN3LhEz8osUJPXjh90j6oG47vYlet6FpopQpoV1VXXcUsm
XN6oUyIef2MH85COkzvjPc4/xXgkzSkaoC7YiOPK+T+q7cXi+iPpV+lGxATgbOS396G6PiRI6hTW
qD3XoWYK9GWJFTARSqMfmjEiLTZfZQHO4eOs1KiRfHd5+hixiZkbh6uLGrH1RAHVnsdGLTyogpxC
eDdTk3ftN3cTS8qYxX6dTEGnUpkgie6JMOWnxU1h/8ReI3HQJnOS77IigNhKZEOtVoD4H3yxD7BB
LbX/G19ZR0G3JgnM+pi+iLJnp6H7AITZqjGy/zmOdzSVTIyRS36kjR5XvNfl9Ck4zaklA9nEL/Pw
OtJZR5h/4grcj8gmDrzoOhctPov2Pzybnpms0cRCrotKPm38HjC0B7gBhESrM4ohTcf4DYQBi0Fh
SK1PADCSq4i9G1x6rijMEbW5y4Lq+gXhk6kRNH6H9l5ran20HiHa8GlqgzcUDWUbRvqQJVSFb1tQ
7c3RdP9bgo5n0TDLw0MqpdRE/ic4sKRmtc6xzZPJlzP5RK5ASO765y1JxW/cpVf0tVrDqEKE6CaM
LzZodUg7IfQV/ROy9r51gmRYc9qODw4Y9nQHppIy0I+MPDsLL8SDePmxrVp7S9j3sNaEzeziv9Ym
l6WUhMPMHA/XJefTC6fDPpSIGS5wdbyGoorb5dsmeaA5If6USre3+Sp3I+I7mzBd5B4VH2z4MSky
gI/jYXMqWE+sQvKWLn177wBGoE1w+THQfL/edhlu+EDpko0tNMfunQW8tFONVI0BThe7cNKRp7CN
8dx8xqDZfUMH35By4qxm44NDNRvdSgviephqYBWyPD1MN/wqfQwAp4DejXEK1if3sllA3KcOWS/h
sUvbc2cRo/1ZSZ5PQHomGWCPlt9fifJfb1BdC4EG34WNPXgtv8v5vo3xCy55Yy5N4hnXZgmuaI9m
yBT4+LWElxKr03WtOXkmwl3gHvP/05o/wjOy3B3tXvd1jPx1WNXPu9kXIEpRcBJbkh7Y/ktbutxu
GeFQQBeE0Sj7PeZNjk/wxlmeF9rgtI2cevtsnZS2soO24SxlNq2IB9r/xxOgd2iaPg0IwSba3SkX
HVQbgr1W8a1YfYqg3UyD/ngriaQR0qJIZR3yYB6uTvoCKl5ZaP4CNxbom281ihL1iem8eZ/0zpvk
ctQDE+5sb4yWAIQZQ5qafbml8tSooscDeCjbrVmFavgdYZ8jYlAqInT4R0qjTxx4PPnlP5cFUSoG
5trf3l0jX3YqVQPCZV+2/tlAiyPg72fQRtXjDGTcrWGgOdznTQKe7YKXW/o4BhVT9iQObiQYUxjY
T179R4Fp3gl8JnZvyINmQHl+L5uU/B86EZR5lON3WnjQIJlvRywpRl83dlwZU4qKZpB8u53gyK2V
SwN6Vgxyyzbg/UGiBaPwRd9hTAmIl5DY6g+6UnMZ0M3MbLBUUWn13/dsM0WvKPmOd0Wd8aqixztp
XWNOcmJbge6tWlkHEVD2ss105maB7GcFdZYflzjy3pGdECd/+Rr+hqrhN37vh0iJ2GpLCGFQ60XY
yEOSzI9I+xuHAUpd9jlWj+r1k0e3xvhRk3ZV5gpQ/0X9nfxDH3NjeV4Q3i4t7NYKNhkcpYZhY+fN
L3vR9dA6aCUfPz3uQA+xSbXZ8pLc7m3ayQcc0nrubQgmlV2tg7FU9ezmcfpS8a1W1XQtf0dSvwEe
hBWWlUN9AMHXHTWDdNaDAPfuM3oOWt2jmrV0yRgMe653+vVEn4IENMQ0vwgtsxMadchdJonik+ht
7BfvMXmt6a5Qw3CLqi8pvPSbkoWE8RT/OXRQ3USK2zqFeSkQStsBKxhMRfZq+n3RcqgmfUxJp9jJ
+YeLzvca5HCb9XB/pBJ3xTXmMLzjhm0PsxtlMNH5rgs0RZzIZKGh7TNH2+yWBAWNfo8/TKPN5B9i
opu1/naoRIO2wSRvAfzmzY7V/z9WXDCJmlXp3FM/gKEPxUdDNvfeTbfkFntyUnh+fK4VkgDCrVVO
JmbLVhqcQ9+v4J2LPF6s244dGd4MvNAuT8M7AAw+SpIPtqdSDsWMVs5vcXUHgjcZRKkCwXXmfJIl
I7IyQfvx6esGWO+R9KJuXUICq2L2dyYv6TVDAmdETXo2IwERzxkkqx8oCFrbYpiXlT+gcqX8uLku
T3wuIYLQrv+6YKdQq98DU0Qadn8aS/hr7Mqtu4YbJkVvdUfc3zhkFTeMDFYigGDbyVAi2n0v384C
hSmt0jYGS1gm7FEc9Hc83JPJfGAiiaMk4/LHWWr322GJEgf90uAggXc73PZKRfhqZwrHYmZ8XMFs
f2MtW2ysUyvWz/HgTn1juAqiYlvFQL7uKN3sfiwaeQWpjdIhlU8+W7/jaA2S4SGeRSig9TAbRG0R
u/nmryyKvTCl4udMmGO49BXZQDOf+A4nHZEv4koCHmAR/ISMBGV0n0fw+5CSEehQdS27X///DCUB
/j5ezIWC/bUiyQ2aK9m4x5OAKwD13N+TdBqNqL1gI34lVm0z3/B3yy8PxPrWYGFlkTMgGR9Ed1Z/
lA+vIW+4yD2a3ZWtQZ1eNsMjmDONcuYDtrQWQmdLMolTr3T82FQ2rgvZRyacbnklTwAyKMvPi6JI
SKOImaeOYZsHPl4K6ezLVfjpFJLG5hPYdDMaLVcy/Td5527Ydx8yNx8iGzYa4k7Pd+F4sQ/EGCHH
9V19v+eWT81acml3yPiLmRWmN2mKNCefr+zeeGHCdZfNpCRuiEh3LQHw04OebBiih1UGLPWLt2sU
dZk11oA7VzUOI6zBj5n0xc5HgIwii8YWtrL9ARSP/R9z1BfIAD50Ey3pFN5oEZqOM4CWg60OOu6G
kZ9YeizNF+upM5RhevUiv5jrx6Rb9qQTlYXR9wDjGXSeZykGjC82RqwbtP0WNYTaj9apx1y5U6iP
RwwxI9OdYGaOO4ztGlu7srK0756JP9BY7xWA6SH/M+vHreTCH/LyUq3hJ76ACgr4eIohn+n2Wn9u
/MBv8jxlkEBLyEYEPph2HTlhJ3EU3f0Y/gZa5HX8vY6GQXyiadyfgsNd9lkg9rLpUrXp/JJE8JGq
LfihiSrwgAmJ0lgllv7oJYokdJoSXH7h4WKKO7A4d0tRlLAcu7Li0XDlUScXfBlE1S+MpRPzdbS5
sm3wqaVbZXzEIuK0RnAtjBAXE1DZlY0VT5MiprHTxoaq9iX2ysVoH6RT+psoGyMBDhTvUmTnPEHs
Pi7rKBGlvhSdTOEWsZxSZ2HKoCYf4kbMUtrITri9DB4xxk7SuiEhmBHG11cVGFac/78OhYWnXsCJ
WvzLuGJP/4aesoQJgONfVPtywnNRmItQf8eifxlTqSRCbM7UY1oNt6KJ53vlDOYqLwPdjMMylFCu
qnhACqf/F/i0CuhgPfGU/C3mgDRG2KmjABmYmIh/No6Thu9BSmJriuskEL5i02d2ohNZcNKYOp/I
mzrV9eF/IxEXThJjtOO++gFsctmHrx/39OhJ7Yz8+Rvl4ZAPDoyQVXMDXJEfAHLDJnHxJfiGRbZB
DktA60maIskgufajn5TqHbQY48IzADmO4B+vSPuduRVR3Ke9GZ7bowzf7XLDpUajlz1m7IVdDzvN
Yypb48CKm9eNOgrBWZRuzQYyyDBa+RIsL6fjOyjEhOpKFCt5yYxgVB5ZxOddXFyCyXjR7lyCgOS+
LERRnV0KmONCe7SoOwornM16tsrDwLqoi8A0/1SnEZSOvuwM0GOkyVqdT3rQEKA4vxYhM+FYsDVp
6oUwjPZ0Z48sHhwWUeQo/dVc/xarVnwGBpf3GG44LGJt7sT7++naX3kl0jxCqAVn83RqVVEeMF8I
GImAPaqgZ0s1m2U7/IdEdYpk2bC8GG0aLm0BhEhK6qn3AZgDfl3F0XfnP1I5XvI9kYzo1/RzfqbQ
H/ZElwWG0qgDUTpCb2MBFJURP8Qa3dPscbiVEP4hf9deIt2UUTK4YwM7sRAeK/9IPHc9AEyQMhKu
Vz2h8/mDCJ/cIrRPJjxmfiYPK+t5kqD1WxO/TbMnGZbMYelG6l8V0ENVNi3iMl8pAbx2ZXKEivGv
XlLfQ8pQYWgaTu2B5N14xdiAqxunueho6a5iEw/qojsad9DGU0SxZdqN8/CRy0gAMz35YS7QmNSP
jTm1usNUweNMXr7NVURBZ1F/iLhsL65TiHwmA1qWcsbPPdkbVxPsa63S8QrhZPV5+r0FzywX9Z3F
14jaRi5imoi7Sk8TNu6QlbgLBXTVG8JZhBFQDSk8kHbTn7E2s/KrUMfdnoMJ3RNKMXeZtWtnMISp
qlYOTKpS+8vBGAjE1/Q48cI5yhUqGAiPDm86UI1MeWLvbHii89MmBYKSwNLVE3LTx3OP6YP2vThe
gNgSvhZEpTYPjqVLHZR7cTpzz3gOXFTdsErCiUSy/TcM1u/pZ6Z8tJ7dlQJw4i0oWgPvy20nEaC2
x5csAQFdkjmDciHfrBP9P8aJ2IE+HIzUhAs9hEZEMhE9wa2FBdgib1t89ZS+eqsiaVV4ZnVbWbJL
C2xXFC5t0Qf7pQRH/PE2U+IQmn8e57/Fe827fhD6KK3kGwfEfTcFgVLpbestDGT0rpVEgXpG//xC
tawtgpC4fcC3VmSAZv+lM4m3cCjFnuBtM3jVbH0Pguk/n773DPRHp0ADemlLe1rRbSx2UuVLW8ul
H3+72qiDv11RfNGrS8lEOJBaGTyA7+zDIb0GwnhGevFUYTBFPsQe+OPzl6eO/tU8JG/cAS1Gd8Xz
k9MpGTgo2Sh34SoVNXHvdH43Vc+9R5kjPXOtfflcErUH0me0tqWxG3gHWOkenpNyhEeOKXn6yc25
TgOt6879sXHXSx24/xWAKV2D6/TwuJN1FB03T3sewwWXrwcvyExKPjWB0qabSVgIiznu+/UUc7xx
bloJN57H+63gpccg1aw+aCZgR4n3WKo7MIJ2Lrdzgho/AgIQ0ujf8H54t0nMTduR+mFm/WKSNp5y
WuncziNc+Ihcqa5eVBFuIXtoWGkahjUJhQYs4SB0LtoVvY5gEmuDkU4AHjmahdyt5+5oMRDoids5
DtIJeJI95YYjsMkJuSeEzABvMu6Hy/jf31KnJo/bvH/oFlGFM9LFUHtVE2TQSx6biGquzY6bDiky
MzA96ACGOuYC7UCQAunYUOUK1B/gN8Qgg8JqEj2fMlzsSZYHCTNkS8NusLxe6L7xTLJQe2CHGbYD
wo8V8swzcesi7dwRwEWceVjClD8H+16e6Lj7f5gnRqGNb9dkVCUYbQcQSk3VVgy39UF9kwjHF9p1
jmpX4YbQ0ZtzVC02jIG0kwtf/xpJf659pok8ZIC0wUgYDCNzcA9j9VrpzkPj+1/gD4CwRxbid7Kg
oXQAa5m7aLWrybAqXAu4CmV4cxMu4VaKn/odc9TltrMNBMWpBuLDDB4Qt5COYzc3hfHegSsatqGc
P5bLQMcB/5dTHG/k8KmAehDt23EiK8hFsdIToUcJDigNWFNImRe8x4YDxWlAl9GJLJ3O/o7oz1Rf
Q0fEGxBHOm1/jpliZBA+w4Z5NiHzBIl3zRWlZPKmbWg+Gyq+pZWZKf/0LuFyIYGXqWS8srBOonJv
oE2KvAdCmxQCKx7hbB1KRuesu1VzX6Lvlg92peMyqxuFPtrWJ6gwIEGOLfrFz5nx9yEZpRnmFoRd
eehca6wPWTK4tIYZYczns8HzYSbuCEBcNZK3mu7zPAIH3uLdQsOOIv25iOWxB/JKeuhJZFap2xOi
lHt4tDbuHoKyClzW6mHJAZT/7KJg599OSb+HI5OXzUvtlqIK0+RFw0myTEisEjtpr4mpX5eoIi+n
qv1stoWJp7Nj/u9xyhg0Y5xqk048QThk3KkV+D6j5TA5RGfmogAKS7IVtql11YlTtrDXK87uzC8s
r05CtL8dQCfD5887R8G3ozzL1dRJSHCJIUmQVzLYMFca7EOW6ssAjy8BMGTnnB6S/T0mvGpa/801
FynOkS21QoCKbu3Q9zuf0ppYUYzXeNEblsxcOiaa25T8EVqjGKLg7Gz3HCIrYcotxnSb2gq19kOL
jlk+UHND9hZCx8vtG0yS+Q0K5q6zJOQJO2x5w6egN7QuYoPTUgZRw2exrc9gH74YL4PX8Hi6Xlcm
xY4QIjtkbPEWLIC3vIpxjRnfC6+0mQGMiov/A044lJpL6MBa734jtCVch1udnmffUZ9wGPmg6nmo
On2xkvVwmGpMs8rqpKAA1D+tmL6kQfjc00z/SkutA2G5mx00bQHtlV2W3dFQ7Cu2V3MrjUO1dL1J
vDmzdBshnH7Hj5IyRJympwLpXcvlBsnsnObXGD+uU+ryWolZp3QU2nLiKvNkBxbegiKWveTGvK+P
kJq/d3pGubzeZmJYenmdF70YQecMPQZV8ZlaZuRLM2b3ullwlcVtg8YvktrjSJmMSt8FkNIQbc+6
jSk2sYmju7uR40IbXdoDZp9VcWZtGsMYBerdwN2kRuY5cY2QI/p/SeMkePlhBJ8Hy9zjOQlz9yz9
7zdcVolu9Hx6BGjWOYvTzpPNlHRY+zuIZxEjosRL7wuBcommkYLlH5pHc8bPf0BOx6rd/fkcSIJv
sgK5gj0L2h+bnN83Fd7P58Chl7gpYsXqDGXqDRysU+y6sEF+kGSCTAcinwVGfJETcGzw+13qP4aF
7zo50xGyYtxAcMNRxHutapSmWWipJrIm4xRkjkwXVzuZdRburR//ihnYx7urTwM1/i4HqlbjABJj
mymMtxdhhPkK4VULpjWCVNjKkr2/LE2bpbKMyos+gnustyR74gGUk9p0YC7bTSnwgvJoBC/maIO5
9AhdK/+xsO18WPU96xhQ2lQcDOWZcgjBQji/mc8dz1GLx5PJ4IgibncJkPHFhBtIA1jnWeFv61J2
o/VWJxzKWIFS8dqpRhlRei8d7z8Cz2wOVl25cNu1GLkKwjjNWdvQ2IcGGJ/HeIRt4U7JzIaD8WGr
7kNS7V7LRZh88OYrGQS6BuP94mt/oZjPVPiv/uTtQZTqI0kHnus/EinuelxBQBTHkFkKNG7EvpHH
m9SNoZEzezkP3KXwtWYH+DALdyMTtPLnI186f9gUqcrwuuxqbpH7qx3MK1C4sbJY+H1/fFhk8EY0
DUgpVBqX97Uoo0xxFF6EzQ+kPkQG9nLVABQ4erB4CjmUHAvWfnB6GQyFhZlup8PSElNr/r1LX48N
wcz9e6KkZc+AIaIX9a9OR670cUla+ORzrTb6p6tlLTc3NAtSgQFNR7KHhJwmnVKorWbB2CgpSHPl
rAw/GpEw67mGXhjE0aSBxSZlB1+JvTwFOw63f3nk/BCRVIyBs7bQbp4A9k3zmi2JuzlDClU4jNPJ
97vR+i4SgaK1et2CafwQ0IVNo7QuDnaUAXqQzoTHLQhUeDJF/BW+d73vxri2xMfCjI1NDZENkwjg
RQU2JMfR3JDLpTDjn77rcT0ptFsCu3Og15wkHMmaMJcsmtyUhNxI2tDR27QjCgGLsqKiPd+4m8iV
21lu9se6l6zxk3MxmbdmYgYetb6RTbl32I0QnxPs/OI77W3KifwyrUoqYT7uXgWGO/+r/y//1BNi
JkHV35G+mAs9aB+BFI5D145MTsvTK0X87YDf14kXG+qdNAeeMnNgXodFX29J8HY5G2w/7Vfs0but
hIj81rNHYn0BZjN9WeViawaEf2TdccF0955zo0CFlQa9F6eloSNJrLW7KHNP8J1+ulcxpKLzdvKc
ScckWvaRSqsxO8kRWWerUK1OKZ9PIM5m41DmMKtBSrseyRaaVGEvumO11miARCeQdmJDIstGZ5Sz
64Fd02RYIf+UiBOTf7xnKXh18srsvRGrcFcO24djCkUrGC4O8HiRNM5BYFqUy0cecqQfBBCHX1pK
erIfwywj+/VNlyIZfP56mHoeSrdjwCw8HMsOYquQJSGB1lgAcD2yi1y9Av2CGj7j5qI9hrnPdyCz
o2g4GSixJSGYUmTWhWm2piCqLNIAICU4DqR1bsVpOhKqi9HPtwClIHIv3gfXpjzUJm2ylVw3m36a
06+CmFRfgFWybWaWGiPtYhSdrj2tdZFChn9/6moH5LGcBMj++FySAe2ec8b8qCDzywIanJfg9ziu
GX5Z3SLqq99awSEm66kDXCw8seb1yZmRrxfYb9JNsdUQepuKYBefdMD9c+Zt4sNtXJLvRaBP8/2+
H/zF8T7ZECox+vM1nln7qC5IbYqSWzx3boy8UP7DnZQyFeE4QpQ++DsAC6HbqSNj7KR1OWKunYhg
x1PNcgPwnzucfEJaDdpr5GKxv38R1rEm5Ip1VbABvbGqbyiqKeykFm4W68a+d67Ni4Zh4s83fEJq
kKCZlB1HLy4jbG842CBBTFDg3DewWpmK+ku9Pl24cxa2vZYCvv2J2bhbCdRwue6dCFuQCmarDNBw
GC2sc+JCKyT/GUWdPF9bbGJ3isaZ1CytZz4OoWOsvlcL6PUnuwugqPshpSrwqYKYwj7zkfrqfVkW
uWA2EbsF8I+d3DJR+O0n03J0fTbUggUJJEwvVAawYH9aJt/RGS1ShmLBLZKmORPAsf2OZvo3Qiyh
F/Y6c2ijLiU/Nj2+iSY6wTAxUeglIl7CbLBca/JVmDZc/gz/pbNcfH+bwq9yQxcpnOOTTmFLjbJa
HT3KpDr8m16BkuwvwGLBjeK0MN4xKiiAzY4L5StXYGhBaiek/js2AljsRjiAqpQTA04aX2OT1RD3
nVraJV2SYHrUBBfBX0Z5hSXUwmea4LiGIliWT9Heup9We0guzmr7E079gf3w0OqMH4cf9qovP4jB
a+ceeffsDSVqal7TY9sA4BkW+aIV6MK0PJa6yK4+MsnKZ2D0vCW5HGQfLOkbk+ZybpWdjggSSLdT
0XjzYzOifupKNt2pubI63lU2b1Wl3qzKj+gJoTwMudYyqT8Vshxf6Rfc5Xua0IV+ZVlCWBj8GA75
3qH5k5M+Tym+36Q3QvLQYtjWrwxUHWYVKQxgGsYMo6DD516FCcy2IcP65kbGBoq5yWM1jQ7J55QU
EpEvAIPc3nXTprzSP+/tgd+iOrs133LX/Bq4UjDanIZzDAyCqsJJNkNCOke+wmnNVfXGUs407IJu
kb3KgovjZWdlXht3ACnH8jZG1y6q+AR/nRGHhs1TykbCSu7bJTqeCFXvMc8pgNsVnMpa3rINrcDF
wRlflbTl7DaSF/7t+lyt073BG+88TDHr72ILc1IbFtZz6KmbNEQzpxBsPIJ+bulJX9NX7hSaYtkq
BmQo4b/cB8N8BlVUaDpdY3bDsJZhXN6Oohm0sPD1xDmq4oUPckj1thRChJtq9Z6dx1RfNphR6vF0
4thdSZFj3ngva31uQF6cWBUGn74CMZYpNnYVXqrzDejuzndaT+owsV7lvc2pNugjkgUgf8G6hIyf
ZYD1FSqBL8SWgAfML0aRG+WVGbdVnKiVCItbxg1CHwcBC66fLCiDXSHKqlkMjABWFdhxFZl8WIXq
uB8VAP3teASPljdkoqfJjLjv5PJCSfp2kZbMcmkeA68Yz+7nOrXVzLp80pw1AjNzoM3oWT8gm1IC
R4J9289YlzuKp53oar4Gsh9UA80j7beSj1IW7itsfqWq4wVhWaJjSsQ8v9+jQSbv6uu4Y94BMDWl
wVeJd9hLeEmt7UN91uTcrCR4bdQDocv8yqVa+BqcCENG40Zrx5b+ezZ6KT6KR5xjLGe+BuYrc6xc
ZroogFgu7ZCXMwyTs9nbS7P2CYaTNafg43L16uKA4nUBaY03U610WWH7dsuN7qVLoE71FCgM+wxR
9XZW/qHMhWpDYtXmJejZK1uUGwOEjZHsyj8zJoJH1E23CT3qnDh+0pJYadx6pmtzq1Wr3QSN8LsR
N4fzjtBtbWUQq67batun5JmodOgNotJ0ia+WMeII/T+Ch4wVXoK0yAQeLw4M71ZWhYqZ9oqnR2J0
q2wPYlWpquyb6DtqN1rjJL+Uh4v5UzCjbItJUK5JjHkAY06YsVXnTcTaIYnB2O9EuGbr5K0naYJN
boECT8QVw8QqW+DkxUBUciTA+BsEnzcCNmhoh4qof3Nb0dd/j5qcDUVq7PP2r9DQOXEXg9y95pz8
/hyJzRJk84PJf+P4pkq5OiC0mRsiK1JWa0k0v2Sqj4EkYhdXxXEsBanF5onVr+VNHrpqq+RSJQeN
PetFgqRfdpcCpE0HCODHhTHhINDLcqxt/ZLHZhfLiJgNXkGp8Iwr3iUwaDj5/z/9hi6/g6U028VV
c9w/yccKhszW1aEF3RrEMqa/x5u3UcuA+TgoAvG2HrRM7IGxj9m4U5LBkbCo3LqJD/KvG2zYQpfd
r40mPdvytca8j64V3Vft6P97i4S1YGDZ+zvaU13yBtXXdU4G9I7do3dT2gvVK2x5edxrZ4/4hCJQ
qDH+iMRGK1gzgWw9e9HhxA3stDL4FTWXuJ84OlT3l+XvBiefVfTfVW+7f0G6mcV4a/J8NGXSKi5T
oQOf+agv+6WyQaVqqxnPpadClX7W+fWQ7Wg2eOWNQ+HR8EZTjz7fD8aox5wPTpBl3BO06XOjvWDJ
hmTdw7fAobRbr0cUI3RKuswOpaQwhLEMHjvpUgA1X+h9PXjnU2N4lDF0ynQVHCTcmE8BBsTkft73
NuSxGltswah6D+0ft5qCA7k0KhuJwP/HekIi24EnU1SZ/aviSK/VthdHn34JJRf1m14ipApP/9D5
VM7yK/N//jUW4ih/RAEZ5feD8O1mKE5QZTSjG3oadcbX0eURGCs8ospbF0y7kdHd1042qszEJgzV
u3IJJB40pIuB8Z7fv20LFgBVjHbBgC2FwfacTXXzew8OCBxqsMcs1yC/VHBbZ55EYonAZiEvDQyM
UgJf+86PV1nJiHvHMMfd7pUGMec+XV/gwipE1snl2fMAoc6hiENXISJ3dVty+tmRpWElibNmq5me
05cKFKsMl0ncfi52juhCvdS3poUZ+4mC0FOWQZj5Ft3cyXKHzah//KcwVY+WUbeF3jfzcyIDIx/r
GNRToKrbqhNR7U8T9ax4nBCIYkeQLuEIIpWkOJWXGHwN3AU6tFjmQfXREQ3AlcH9/K57szOUpkGj
SAEZ7GFaY0GdSi3625gYTB4m0oOxYGkZjWlf67UNfnFqwOI+OX1jlJaaWYHka7ZTxR+xLcaRcneq
eRp4x7rXGebx3ZHZRb5eaemVUsbIhDofhAEYqqZVxRKeB8MgSsgnpSmfSEfYGEA1VwZTAZzZzu+t
rhIavNjMELSSJTEpPjrCovYUg4asbHo7nFhGn00LydtzJosZOR0d11pidV/skuDhjbRa5ycT6Xdh
YtWCIJH00bn6QlRIct9rLVxShHJk3EByEy9hfkD4uGbujkb5qtuQMNbPws3rvC/vG6sovXCu2+dL
bBDpDwv+vc5XxhRL/CroQuwD/gDR27osZRmcvmqjqT7wDOEGWSTYtFqh6bGtkEvb4lZv4pk+0ncD
osWuYXakoo7Rw7ISNIsEOKC9/fdWJ7oSGquD6iUO9ozKrg+BoSfIZB2ft9avQiCalWmH8+dPH9Ec
nB+V2oALvp1WaY/cqgU6KhRnClAYFDnXY1FVD4besq4t7qt/H22Q9NKQUyi5O3XZ8ReTzTi9RNaZ
I/hh1p+q6E+LmzhkmdTG2L1AE0Z/ZD4hukPsTog7YumTcx2N1MsryIIWVc/kwguT8IgCOGBcy5P1
CYP7Z0YI9FWdvP7Z0xh6r+FB3ltPuNAnJ3giyKTte+n2fUk+lXeXcE/yHpnLWIbD6y2dsoqd2Pa1
Zee+ie5PI265zyG/Gj88H1ka0S9VTLHzKDm6oFJw6zkns+JdAjSQZWySp05+K1xEwvbqpNTnbVlq
QagNTt/vemOl9NtLjRUbbMC2JwMjwoMPqLMALU0mV7VNMCQ6jYc7Uk3BYRgqWz4QOtlMmykgL7LI
ioxCyZwc4o5EQU68R1Tt2FieUeSpF8ZvEv0G/85P8r1AdK5zOwoYrzj/8n40XD65kTEz99+5VM9C
ulaKuAy5CsJx9jUirCe3m+BFZpbDtoypyYy8ln+l+BAe+tAXyITZotpkmpF+uPeXubi9pVc4yi67
IvFD16EFb4oy21nNSGU9AHyLZRhRJ/sizV4nu2gnOVqVqRYKC3wL9sO3BAvbvFXSmvzO6FA7aXc/
Npx0nBm2KrnCvmoEAR/fhPSavSoafckL6M15cDCPj/7CmfBi7ZYDmThdeeE7RGWTswRfZGhW7Xsx
JwoUO90B+dK/dKPnmMP11tuLDFIwAVNjC4ymecQKFnhPAI0khm0dGQpmlS+7krtVNw8UTnOLn9rs
r6cY8Ulj3gizkxFczan468L/riLV2vIWriYWIrnzQm111ruhg45JJrTepbnyhG1N3IRDm8dKjPOi
cV2TeFQK8RSHQzRbm2niCWrKUgxuWiC4GwjTj/vPFJgTjFz2afKUvbC2vMcvOwVIkx5hnKtlzHa1
yUre97Gdr83LjeChKqNUM+PVceKUFtm4UBCq81ZJCMQTW7FpfCw2Ln5PKMbUnqmSANJU8ZE/K4Ce
qdG29YWsANNe6aKYFrph0wfF4cILfOGS/Xu6PxwydsoC3L/1kXrAsotmjw5YkB7nKtHe2imQydnz
GrPyz9aLf+vus430Kf4Tvbjg/3QGf+uYbHnwuiUqECS9sUREKto4MA8tUGmY4sihDkjtl5xGROPo
uOXvxA07PXDvGqrs74lp3VVzAYQ+L7S572I8rAXoT7BpBoWRaBK/JVGxudLCTvYZvZR8e19bV9el
8Jw3zT1ChyawaZ7ccuO59NOPLNiyq1M6/rcBCnj9rct5VyWvI4gF/r41a/FHX/zliV76ycDlxTwT
bru2LZbUf7AYQLh/mUhp+t7QT8mGVk6YeB7gL8r/2A5tRtUT5ZSX67fPrKn/Vb4jcpZdBjNBVzrM
Iqr30ionQwN2P+BX/M5E2vuIGoJhHeQhKLmSwe1IdipkQel1IAAz0M3BB4+fsNKyEJZfpxIeXisB
sFGsb6Rg5wVIHaWcuze1Al6y63eDWsLXmnDmZkKx/UNotAnx64fy4sCCE9zyjZzyUzP6dOosqinG
/ZGTDEMNrJkEjcEdk942SOQBx0ChKJ73bUR0bgP07XB7skFVTBukVg+k3jQbQgnh01JZLI8jMX4w
vqDlHrEHm2G5v/CiDzRmG43ZGFVCUMPPQyxMug6XmJVKClrZopFoT2IWyUuS+rCRTh5DFWbOuOaw
DhhB55zwbibL86DF/HfKaA5KYCjrbzXfsEXMIyBXKC+MMR/YsIMPvkOlIkdaLX+Gt2qCHeRqyYSN
95i/4G//q9VFELeZA8sf1Icuwht6Km1cgNJZFdHIHoXZM96ecVRdyEJgi+pTf5I2y01ZcT3PwQDK
2JJ2fnDhdgbGx9HCvOiXLuLbANo0ye+FXpqvo13DYu5o2APKuzHDqROHFfuObjMpcD2Tdid69Hks
eHXK2NFtU/YOrXUq1qfgP8tK9aopR4Kl2HE1GE8uhYvOIuo2teynuZRyG37UMzhuwk6zpJwJrmSP
tj9SXPs8mJhUQA86AKJgwAaArl+dDdGBMbAnPCymC0wL2kvgwaA7fBesuxPHzYkYgerK43tX326Z
f+nXp7s0BNfwrFlWXj8tGjSAQnrF4BC47xgidq9mg4uy04Ca2oskTn6DYPuwUdAR22DjnymR7H0T
rvcZbRLWGH+Sx4/Az+qjfYtM+a/h+7fhroZhGheRc2DaQX8+OV0gJjrgmCLtoup9ipf1wbUWy/m6
W55LmQK9bGLeQVE5/mh80ZI2O3G5RzZHUa173iZcC1xAYumyAAQygcNF9cgtv3poR7TINMlQN42g
NlTkN8SL8+u7k2fI9yR8q77O5Dy28vZphOU+psm8ZYpkydvc4JIWDUFWcSHRIryGCzKkIAlC2n9y
cXILqS53jkYA6xW4VacI8UgPfsl5OyI5eIo3GNOepXjXqsJYq8hrlJyp+fpfsCVHBULE41ZHkTeN
BTCRDKhJ+Fk7EG+5PX/eVtY/TBgFFddY8bZ1/SRFyR0Lhebbte8oFl83XBWBgcdvkbE2dj0SfL/2
fTitEjNASs+Y175v4ZHY6aKvZ5vYrMNUaDPPk5sLBYGf/HzE+4t01VvMAouCSjbaIrFK5jKl7+m/
3KolNUBmBP8KiyFsgjL9IDmeNGIPvE+CbNldoOgY1ovDQMQ/nQMeV1Wss47qazqSbOOhXs2LiKYD
r1VzvnvbODrypNs4gHKkxeFF+UtwEPvAykicxoCjpdN+GazUKxhyo8JVNazJyUcFvrDw/R9Qyz+U
e5B3mmeicFrkn76aKWLQJk8L4B4JNsxytsuwraz9yONblPD0GmZxSbkBSxArkiSeRrsqnr4cT6tp
2bn8uL+A/k6iCNVgpRLTaUbngHUKRA5yMXsPPGBq3aRFQKSvWH96bd3zdzzRGIi9qYBGO0VvIDZh
p2pe5LbBKOsiIL21puC7uOXyIqga9ocq38duIGUBk/bwO3/Tktwydfd0F0de0ES7e+d35PmZSoyM
s1K8e7mwX4CbA8/5K59VeNR797bJy+HqZZtAUBbigHqNGcwTmF0H9maiWPJ/e9i2E+7lqi+HokPL
6mjICF48+ka8fxNbr6b+PAErXUySqVZpWeubPAw2QVZ74XSPqktmV8+ih6f1c53O3yUC+sp0hSWt
jbsvPOHMQiaroyL+dO2TPaLxgzEp6YRza6thD9Ysldl9j/CA6p2WW0fevucvW+bATqjckVIddtvN
bHYma3Hinvts0MkZgsUV4gzpXFZa+pGtZvy+CDqwF1Vy19EAIngjRq6FInNNKciI8xcfdaFEKzJ9
az8CqcIsMhDHe3fNNkIOVOCvNANsPSnKt6V9V5tYOjGfBf3a87/B1sBNMnn3975bZmHuIOqHA0zB
5zbB+EvX6P6BgwzlhMI7gOclauw5Sw6u12b7VKd0aCfvnMOSKD0+ZxTvnEIvmLKWxjfjiKuJd+VG
Gy7ytzEpm6DKBQla2CT+j8VVi6tYKHEFYg2d8GeDD9S/ptST8LbloHN4lCOVk25vYbWLclbjXWLT
fcfdoOO2k2P3H8Bn3byaAeGrs6tHeg7UXO+zPoc62CUkHgLg0H9TOlub0Vwskg157Sq5xHtTq7tK
BDyPzrJ4nyKYIgiKjtODtmPgc1JlIU/UYprQ57B2uY+gqmhovi7u7pz/NhNwbWg4pAKoLZjDi3K5
ttEA3CaOinKYpkvQ96Ruf9ZnWAvXouLpwIN9nRK7UB1poYgNQIG2R9N0bNt44J3e8IFVHOsWwXOz
L42IWYsjar9PmoOSWvBFRzyyjmpWLP0HgK9PvR051+o771RFQCLmZw+orJiXpi+hQjywFlBEnpDk
HkZ/AOxn635YLVep9Y+BIuvBJi8HdthCsI7BN0GufNpL5bmtU430X5ILb78i2buPu94Y9DkWywqY
UleoXRG+XFqsOpJOgoBuRvypHweCRtVOiw89gcxKrGO4HbVUDWRQiDV9kcteONyR/eO/J3NGjDcu
nMQmihKJ4Yqnj+chSJw2Gf86UakiUSXP1IgKMfTbWGt80LBFzdzR+6jQeKVMz9GloxWs2avsWQvD
golXBDDSAV1MAibxyrZZtMvG8kSIoLCuEYjp62+68MKFQ9bucnLl5eTV3uXDqDfvxUT79f3KqzmG
jlZGhjghZRpQShvTuk40nFsSsSzXIeCsYZtMLKNO6hqFyiVvK7h5VEPzPyKBUlP5jR+zB63muea3
1R6gjISUSBrGxdN3VnLL+LrN4pMwLKqimKiiAPzvjO+S40B/XjV6ApMlZ+GYjj9cm6PRqkn5qUA6
h33QVjPVupVnNjnwgP/Gtr+doZnwgABnKwtd0It02rH6qYoVWjutMPoYHkIcF5UejhqFRLsaotN9
Xu3gjQEdO34hJGx6GhSq/5mJTLZhnPu6vbmrfsSx6uDsHOr0yOEmkSRL8HsB8Qx7E5Ba4ifRnhk+
1R5DQIumumF4gwgYX3FdoVeGeVrCIlh4MXqs5OrE+ZFV8yXNuR0cmA/Z9oEMn6cg/z/spuh+EIvo
kgQmHUbl0eqwU2YLOy+N68fL8xFqLWQfJ+6ofdbfbSJCe8j92gfPokpUqmOrS65EnVezWgEYImno
mLUUtWwAo18s7IX1xBq2X9o5tlptVsstrCqVQguA+dKAqn/sligQIZRzab/Mxa5Y4P5PHay8uS0b
+KRAIgMpgW6alPSM6GP5E+0HVU5ioGqwo+vFHRpVDTFebvyTjFt6MpvAm0Ps+TPaKO8WApV5Skff
MLD8WtHwXfeWQbjs2VnaOm/r4P1Hn6Y+HXhHq9WtODNR5Bbu5uhuqTbWiOt0aOZiMV93YqmOx4bn
OQltv/3v7bu62ZoDUbJGWZX1+GplUC5OjK8hh0J4CdBBppEyoqRPGUPseGXBklR4mPJk4QXGJCl7
1k47mNowduz51ZFFGJQVkT+EENUqiQc+xzLkAKMs3W8mSVQo+nnDn7Lp3KCQEBJUWJR8cm9IummS
e/WnQbcEIN6omrJUjdeOnsZOAwCitpOXTT3z0L9CaZKx5FXWB3Z+R55r/ccOyS1lFNLYMt/GStBg
zZ6EnN3zzg0ww3LOo18SySUsCYfMlZJ4MEigKFeGuqxotTkMqvUOZlvlIqdezVP8wKyJFAggiwlq
o/Y1UVk9Xmz37Vcp9LphDYLenVrTr6myu8vT+ZggQu7Ptdeff1G6u5X2gtqOBJOfQKuIRKmuMH4v
AjKNouIEtqm8KLrdzBMijaazvVfssn96cCzME/4K3rB7vugRcCSOXB0GR9z7QkxID/jHTuDH14LK
ur041nvk4EXfbTrd2Cc9n3/FslwczfP/bYZtRQfzYDnjxWECaiCwQ9chbHaliuWaYIbnccZZHfdk
hvWNH9wUShWV+6//v52EcjAgJMD+hM5CGQ/rJKgg+A9jgoKARbdcBTQcIJbf/aECcyCLj4sXbeYA
6r/kVuw2NsrDksbGyzyCDoWFyVUtfPgHfxRCR2Au9aHynJlmxN+sC8Cz/oeHN2bgtnupIR7rXBHA
2D1hDHWfhrw7HEavOUsrKaniqQmDFmePsbgR7O0P6bm4ZZMPHKTvwqw3B3OvGm9RnWBJ0R7iGT9P
m6SMZdQFUvUZ9m5dVIk3XIeiiMuvu2QQdj3xo1GshunEgr6AIVwuVI0LgRT1zRgt25Z3nId1FXO6
suXQlDosQmbsENU0WvRHCgRV0F44YpU0K6ZkEWuMnYt1Bpb9wTHs1+yNwtvqNeK7MMmlxa6C2Dlq
89Go8opf0iByFEApXZzDvagZi7kiDlXH+CG8M7FjV3jigJ2J3QaouSvz6f3ea6oj8Nm84RE1CKPK
d+z6kk9+S0BEimlNlYcRhVDqKV1U+ORFALtEzHLPcv1esHalCw3tJi26RYSzIekaA9uPCNLy0LQ2
oa1xxKmdR9CQ23cwvSUBWThfu47idFzKHKE6LhGIugr9c1zVB9W6xx8jOkERsDFjQ9W9nOBWBkFp
Mo3Uw1bsH1oMYlx8jTOEBwmDr1C43r0vjxXMsWPseVydVMjS5qQMunGU8iuv+XnPiu5GO3C1tmZi
Nd/KZgeDspRdG+MMzckIQkWdOvWe8FObYxQKbowTxfQrPa6v+hbclec4PLG2zO3eGMNqgXu1ZCF5
FLaLpVBmV3uzd4ilOfn2eoJc9qmufOCuG4L6s9dMBaDMxEbUxhBJvPqoIL3MV29gkVbJY1RT661U
NeTk4f9Abga1V/e0gtMrgrXurej7TenI6ScQfdqZTCazFYYP6zm2MKmESFh7keA3oWR8sfLXVd4r
rrCeI814zqr2O5V4mpST5DTQhLDnJqidrjQJepNC3Sdjt0T+dNGX3sIrAf13dE4Ie3+Yvr8+/BJf
btI5L2I1OvVH8sGvlgFE8WuAL14EL+P3CYS9mDynE0gNl0ZByqesOYs6/Ll2icJXYtDstTAo98c0
RQwhNLW4VWYardNbWrlzrjZmYdHBM3HQ3dcdbsadz73CsG2ucgS42ojt8tKIB7G0nJWCnCt7r+Ub
aylcDflrTFuyLFydlqKRZuOEFysHer5IKGWFHKGZvOr8JXDvPSY6IoLEE9xZJ2ySATuSv8qdNLSK
rKO0ADJNjwZvXKrFZXu3Ntzz742nWUrf/Q8spAiKyaBTS+dBRsug+R5U3IyBDrMVC1V1OyqezcOo
rlTxjusNPWZU/ydlCyqK+xEyPaSRo8sXmpv9V4V6ebdj4MM0wfJa+K8Qb9wpGlDYDBm0gJ3gvLb4
kYtwk+lqHbAZhO+w57/LyAUNpQ7qDwQQZpznBjolQjHDfrlK6TWkKqzqmjKu4YL0UyPX2S1FilWr
ew1ajTQa2tdp/omdfrTjJxeASPLAJW4UUMzVn5BLYYjveTQ486FTvQ2WH/1onVvXkJbc6SPRwy+3
V1W7Lg75+AOGaZxyeMY9rXSjZ9fv2gqzHnVhIryMQRRVW8HVOVsfyqGzfilkR5C4grD1cHB771OU
flh7GNvYcG8eEnTLp9GBSSzDD8IgbOXQykCYVdZ+yzi3+l3ugOIcoyO8tk20JTFDhXdydbP14PdT
GGmARobGVg1DEF4bUtsPaJ0VM0HtM+Dek90qE+neHax1XvaqyzJPbkoBbinhujGsTyPjcvMjnlDd
+2vvrJ/Tb8Igk3Y9q5oTrCwdMH3XZE43gksnXAwrnf34WrkNOnr85VylK9bhNoLcTc+iwQDf5tmr
UkcrVb5LPTbRHCYPMyGQNInCrCG8yKCWs7qLhyNjAsac9Dj/uL6eaEutyVd7nhNKdcGjE8vfw6li
hA4EvMJDVR5MOehaL0Nuxdrc2XkqKnm/rk/EQWiOTQuBOKLW1RXNQ+xappNvV4RVtvy5LOijZ8g/
w6s1hd1ydRTqjHvSutznfTfYTM/dj09Ay5ENmBzxW8W2eWTKEZwWp80ch6Yq/alC5F6fMTa+lOh0
wpREF1MsIP4Ie7svlf73vfGpJEyoTzwUGxNYw8QUjqQQ2TJx0fBBLRnd7OSz6PQudXoyzIWvj4kX
mQKpqPjWVo09YranSIvTpGGmJnZpSHuTQ5feTbJ1ziXv8/fP34KH9Uq8N7Tumt/K4X4AtNmFejbU
/i8yOQixS3YBQAday9MRgcHlFifHPnivnu7jMaFQorH4VFKAIluH45zO5ytthbIvIhUBFuDHTk8i
jbwDjtv6gVcOAgnzW5Kp1ZXgbhxnEmQF1IAiMeJ/LpoChfDNh1h0j8b3XasWvu/eKgcQjojHzL+h
kTpu8AJIOcPZ/lR69CHUJ53yDKVsvrVyVTkpXzZliVeA+yDBvLbePYqbxfpJDIkGMOIOlDvuVaGe
FTx3Ab4AyGrFSzv5YnCSNnIPbElmGgbQ2YYwDC7PK9a5JGULeh1HENySyiZ2MQyMiABFOZEa1SXv
2HYLC+E3aDLjDjtstalW53ny5CFFQAqG1toW6SkaTaFsSl461bReoWOGBFuFVaG5ToVeNWOvOdKS
0SsbdU3QdUEbgx8vR+WuCzFUkiVpepIJjsN5hQ5kyWrE/qz+aYt6pxFjnZo6MieVTcZSptFPyb56
YiuYY30QCbwJojuN0g46kSdRRgQU1Wr1uwmjrdsID2WStQpsVUNqF7OOqd/iox/L3p8tVyr6piIM
JjbEGkFeUWqSp5DJMFHiJkkwaxPmq/EPPAAnhfCcLhQnPDffIZfn1/tNKiF3t17cW0H6WN3Q7bTJ
8cC4XZRi3aVH9ffhvX6a7eJVASCzQYwMNJCUPXcklvvhFYZ6pSEN36O/3pMstWlGhLgPF9e5sBCe
F0rJYbiBAvidrrGCQyMgfp7TMklxKzp9K5VdP3t7Gzg/DnUEYdOF197ucGbWJ7vVQf+yGZ53rgTQ
Ii0RRq6Ets2u318OgommtOJREpkzyghR+QQjKvhrFbNO7R4bh8kaScMfC4BgpOzYTbiCzzGQ35B9
x1APIAD7VSXeDIrkrrMaVuRj2SKVuOXgxHhiAP+kFOjll3Gpi7fe146EDa2akPcGAlOWSyOVEwc9
oEg0L8bSR+RLwz+Ewspix/yBygYXlTIYwKyPR4Z/v7i2OCX1I7NA0AWlOoRRiTch440kk/GH+LB6
BePyiLv9urCBidGMnCIZyhWnflovgdokpeW9USwl0MrHBQ103I94aqYYcPEHBRdB9UpgCgXlE2bS
d/DQ714zn7sbY6MpUyft56N7aS2WzEuNLSfcWTAqBXW+jKaBpTzDQHUwYtE7DJ7oywmuEZ1am13A
JEr8GwvmzTeLPMRsQKidaRStB8VY2TRCq8mwDOb8F0VauYM7s1/I2HnefjyXkzmh70d8DH3so0n0
+CN3prcz9rsMIU12MxvrhRzPZNd7re2OYxJS+6Xj9t+JXcN+pYMzeKHVw4a/zNExbOKQ7REwDApx
pU+aBsaISrKCchyLuMYJ0/y+aIJK9SH92pRIZRolVKC4q4BeSgs0vAEeQELrWS5h3BimrgQjJ2IF
14fjmhUl+hDvWV08zULhL2sTkwXT2kXv7nWkaQfPbLDKVSGAnp6229LQcm7HYl21aaaGL8XZ3ptH
KkLKwQ4jcaezDff8nnMneAA9rHw/nZxeTVRkSiYnBzu6JMSWDK6ZycTv1et6A9f2MfCP6VZ+qQ9B
pwWL/QARp5QcR6XKa3jz404CgNFEme0UbQClLV0ADqhNJjOF4mT3XZL5490Rh4yHP4zwwHlwcyrd
098HR7p7RnFoBq+RDtJus8bdrtC5aR+yVbEq9Qt9fyEsaO+d0u0lMKgK5dXsD2aNkL3/Rz/yr3Ml
Cq0gZNv8S25a7C7PAa/pWY5yRkDEZ8J4QlikLJe883VqwQnts2T2ZkbRhiD1E39KVTMiYutJhLme
aihn7O/wy9jzjxyqOip86C/cNUCI/ZVVxiF4ml712df24tPE5KA6eW0iw7vWjJBbqPPvxhIVC5+W
7X7njxn9ijHq0OTbw+7NrJIbxy1TfbJqrdpONZ0wUWoac8TzvPXj9jXOLuumfQFUPCk+2CtwDit1
bSI6XAdyO+unhBnFaiAXsaH8fIe5TPsYARsPNWtjCo9lHHIb10J2uX81iEsHgZijt4cNN1ywjK7u
REo5/GDtGXuHrkPNPH9oimNZ7qfapYPBjU/MiU0eDSPBx93Qj3M2MvwXOHprVZOB0glDNl2C1Z1E
H74W7mJicFiGtZchBlyELvF9No4NQEKbUxvRMXJm8e4hF677hhrmnKYXyBZY5er1NqahRR6avXLI
fGYcwQUvIzh4yPqqloMeiJojKbfjUz8nLPDpvdgCEtWWCrNFXRmZPFWeeuXJh/FpO3UTpElSz0py
ZF3ozt4BUlpogvFF/6moF6QJzc44Gev/vYgbrNJE8ongGj5JugNHnzZnBLxcAB8VT47K2PQXRJ4O
9g4ej4JgwJX5J7CD7OmsBn89yUoIEahGysn8/HqTZm0gzOx2J4W82PkRFYZJCHrWK4UM9M+sOIxz
GAnE6JKrhdiu/v3rhFbu/vaNV+4CNnUaoISsEu0leCidxl/VS4mgeYvZgo2BxfApaHKLndgiLBu0
Hmzq1NFOr9okEod7DNtIMLNBjqnzPvZZa62alch3Bj+YdVvI+nlI3iNgFBOQVJ5lJKvfC1cjsC0Q
bHsjCSsugZNRM+zZm8HClXF4T06VYtWheZFDzaEAwIk5tWMAKovK6RKCDVRSeVbnUlJyYYVuqHms
umwURpCdv2EPUKyhC9D379zvX68z0rm+BRTHFEVXnaVmSRI1mSbkw/i+ibBQf1/5kOBM3IgIL296
KjoOb24rZdPeT+GA0024UvyuWzQmFXD+ih17I7Xn8hKZXA8kWOhim2aS2SoXuI5uDxvhD+fdeQda
/RQyNJcTBcXC3MLLxiVU0u4435NaSdEieAeakd5oCpgsWBDV9neC8RHT3F/iSv0Kq151urgXEiDa
cmy6LyZ3y3tq5QP/XM8WrtcYrTfY/pEsQxopYloiyRf3kPYvjUhn8eeJe923jYkCXhH7sIAVYQ55
w6CcLmfRSDDr9WJ+mZTOd+O9uJaix5WlwcHB/US/ClWeE7mqoZv7HSiTwL0G5Lm7hdxyZahpLdOQ
vUwNhbNHqOKckNgpQ/grUp52VwlxnvPfb0rRcj8lbnbyeBRaaCYSpze0a0hOYci5xMH5oBV+90Vh
C4QRQpMAV9n5FWSeT4m9Tk59Raw5imm3xKmON0kR53V3rVNbSQdY/tB6jF2k/0dKEUzZi/pzZuf9
5l6BalElEvdynQPtnn1g7aW5HMkMQm2hiAbpi6YbQAg4709GwyRcHPLQtI8eU5AmQM2f/ju37oCZ
4FTpfAs5kQ4n6Q7LsUyMOt/kDpc1RZJyg+n2GBI71sacGRDtsdBxhbQtPHpNc2jDm5/R3Oy61P6U
mWSpee1TtaWQD8oCdlE28jXh4bijj34XR5ld2Cbxh8zxSXq1F/DykipnhDXc0euKqG7JoXjZcZVh
kND8kl+QW0qW1NUV3ADQ9Yy4nEwGbsyJe+IYGxaH2xKJcTtL4g6nTUIWHi2O5McA95eZrDmTK9v2
xCDDdqVGG9fXDixvy1icgYT2WstKXt5HFXKn1yZ6iwFSIXr2zW6CDHpYFK08hjYKhdQ5ZZtzHHLB
A+VXfCDGYWYE/UmUCjvMp07Mpdc9tsenaX5EdOWxiMdu0KI6rmGMqO8im/yncem3ttKLYgieuVwt
p3x+y4j+5JxxzvRObXlCKmTGPt+vMbmxut9hlBWQpAiOtFM3hYwWRL0gmT7K8YBwYzGj8W0VOP7v
AAjPUzsqvdN5BNrF1I0PwXWGiYf9lu91lvBI/ws5Iwa+7hwbl9bRnmDcgj/NlAtSayaQzfBGb7LN
x3spjNpO6tlYwfTubS1sUQwC90h86A4IDk6q3KuClaf07NhmNRECQFoME9f3a/N8ZW6uh8ErDqxr
syv2l+BBLwmvYcFaNREIPOxbKF1A+trTPsUpVEZ5QxF4n1UrSKk5uMgaR4bwU1bs56Z6H7FnqU3G
IxM+wyAFWnAkrBvgXwGItyJyQn5VNz73nHrrdiaGhdGzfGXzJi8qgOIW8WSV0fr/9mNGzBXtje6G
BBLJIejeFJ4IuU6RqLAQy18sMWjKyGOrqDLGFBTVpwffW7aeTRrW6s1O0oEvZk4kVsgL9sP6tipV
srGtCvYnsm/8vb0eE7r0lWjcCk1z9flXOe8d/Bz5BVfRUkFaTNJDNDx4qz9EdpJgnu9kAhQGG+AR
EUY+NR48qpTpQMAxjF4b3GZ3dAhzq3XpYdEPj4LCsJ4/af3oE8A49iu9wXiT1Ac9WHQQZimwPEaI
nye4Za+0PTXr8s9MN7LoFBV+L57o3Opxpz7XNV43isu/L2W2KYSCrFcUCf9+7zFTlG2gM3pqLSMp
JKwPUkz+HFvSA568pSEqhbeTEiUwkQweD+NJtyfUy3ixZoDua5zpwiLyS9AFfcAS2ZQc2JXGdZUr
u2INfUls1doCrRX0B8X+vwey9B0+KbMd+Bj5IT/PKIlS06lg4MXQyNSUPh/tDA9kBCD43vIAevPD
D6hxXhZhf4E1csIXhOhBB/FHj7K56RJwiaiijy4FZ3YhWr/P9zIcoyJe/mO3/yUu+jnEuDHSuG9s
5153iEVSwayaOXbelx+Lih4dnP4dfO8dz9P15dEsRoX6WmXRqQQIhCFKiGKbXhPFBFI694iYNUJg
MOyKRvseknTxlpkRaA8kN4Vo20/fIWQg+wMH8YnBgeRQT0a4GZqBidNvUCnu8HnJ0JRf8lppGk39
MnjWiDZHj7pv5hXfznLbD6Dez27rrVtsAcUcJ9UWkkZC34PI0Tr+2PHMvEhWPriopYpPGd3sgKrG
q+HKCea3vlVyEsYKVi2SG/R1vkJ1E6DfglS3NlQphPmAyywGrY10EH61n2m9cOgDLSmn55NXrHKs
9WqbXTQOqXKEaL4tWG1Uox+Y39osu76LF1vkfid931xnwuPZmdbjiRfLl1MTM/fGBYWVIKD9uyin
qI6C+5wEX/8H4xw9EnLN9+HfASgdL/QYOvJGssGeRGdE4BdLSjYPFe3C/mekJg9rD3HJGaU23zNR
MlwpnzGrXy9fN4sB5F+sweZphALwQMIdqZfazRR81b4iZmOSeT4Ih67+UgZTLPHQamrE3w8RAfDD
A69wBrdu+Nwe2146Z8NiAc7LyhXkX40ILoSp2uElCx5jOx2zDs09wZ2PWnypNGrWNVKrZqwJLH87
TSOpffxZV1nCL3mryAzhks1fgzrmQNOZRVgjgjwYNGl1vHwAP6fXhKnTMTymPM+23mrQ4If7jeWX
bEnq6cSiw97NLQyOgJjDA+Zt6HYHOExn0ogWMZl5o5XpG4h+eSaMKlfca/dx2+Dy6zaYuG6Q1/uT
QiVF1CUBWsNTpVg8LyqCsNuQ7V05q1A+ms4a+EF8esWKE4a0yK+l7ZDZ+31qXLTdz5L7FdUh5trC
hf+7SJ2WZPjQB9TE7HqCiKpjxDmMVm0o0PLOW8lXwsrn1MMqst0oRKt0774h0RIBHznlQwCf4HvG
YzN/FexWNQeQh4xIept7mffLYz4S0QQNjypZje/xo3oqScerz5QHI852Dp4ThIW5f+T5LX5x8taa
VR3jOWw8Z2Z9pVbEeAbfqWR0eh+LIjORfEk+mwOlFhWLxwBMn8wsVhaVMxcDk7H6ANhEEUze4qGu
bUg1R10+a9koznVYIYmxy2JaYpdtL1SYV+9kyW8YwiL10gYk3MTJRULax6/2zW+O56Ys0/FS2f2K
Kw+22Zk8rlweq9fpt+uTBEep16M3xsDg6bDp4VpiWzUCEEUGIaFY6+k7gkhhbrhE2PuCUGHToQQw
1SwVAN6s9IiELwMV+vKOWXibkc0pfcvt5L/eyox5423R4rEGuukwVg97keRIXCH+INNIlg8AvpW5
zBHjddOzyOaeSPsCti6xiFbwnAuFO5cVdS+3KU5/vHtLEAn7V1yJfKvhizXj2zoqbzIkfS7o+pXP
MgRgqvdBaxP9kAWGNiZRRcS3eyJu6Zh/8tX1HoQ065lCQbhBbSMGCOTldIzZ+yHsS3j0r1vV8/LZ
ce5/ff1WanrzCkq+gTyUjLu5PPFqoZM0tHgd/TnwjFpLDJ1F5M44it+6Cmm0KGQgr/3sU0fUyowh
pkymx/Cb5n8JaNH6kV0Z8+Xgqjy/Q7APgLQTVytRNzTSSX1PvuuQv7EBbX7BA8dh3YMGl0YWy9ks
aIEIytaEqNMQ/b85BPVQLYwd7ZQJ+IpFZ2lHYoxZc7x5BMe/lMtY9fvGyjVC2I+5Aq7kdxKefG6R
Llv2HvuRcUJCoLsiWhJ+/Y107qbjqBzVVZjYroO1b1wKq0qVxYoLS8ZEzu0a0VK6+3t8ZrXUW94l
VBtlqEIGxfqfnfrmV/eCCAuNQ0IKGBGOWEBvEFFkUe04imHYfzVVvXCtwtPgV3UMYer7YcY8w95k
A8wS1wFaUzf2UTc4ZOiEus8oNuDF8YEpqDT7wyQfDVerqBrMAjZymGn2Lbu8Ezb5FCbB48X5l8dp
uy4CArTv/kPYn15vFKU6agzXQkIR8dIdBjfkE1jFz3FeE/Z3Cg7ZkD0SEwgxXrH2F9NBts/QDtLe
dqVR2SLQr2k8l/ZMMC2PcyZtj7lRaXFpWVo/32qRLBj8aDO6mn7F/dHEVHLSLSWKMsmi2tgkF4MT
hesV2pGDjp2AzeV5hyZEZj+w7hZhjGXIMBUmjRdq+iP+eSweN97iRvvqO3rGjPAV5yDcnteZB0U1
rZYcQsHEeaX1tPEoCPtWBIoTwtCpEn4O9mf0y012LySA6otjCZpDx+4eqFcnE0Zw9WmwPZGGnyi/
831Ttn7JB+KUB0MpwEdjl89MjZRRiDpDEO2IjOQCV1ix/JMajSi7tEz7fZdPnUdY+RLxK5nW7jlz
pLCsP0zpyeH9icMWyJIQRjQwbV398OQjveq+GOYIHaIbXkCS2rI0X60im59e46XzTaT2jZC5+nMc
Yfalfn0Dp7Ag0N12xQ370Q6oEjJh7OjVEWoBal1cZc3AI2SfP9Jcgwj/zJZxOS2IxAHiBC/G4xLr
x0FqDTpLc7aEjpR2wLMY27WmA4qz0qLy8Wf8Wz5RsiUVrvtgrv+IIHvHQUFfaD9P1CjPtUtVsTBM
OkRvSax+laRA0SMyQARopWKlXrsRAxu8dv54+ufjEGaQOjyb1MuYa/djTtkXP9Mo2Mtpe/jajQIR
oDYXsTPS+JuuHSGIAV3Yf0e9MKOHgNlyOwl75+tImyfffCXDgOPhFAXUmKhRcSXFe1wc4IGQpQat
/tmxc8djKU2Yy+rAIk27JezGSjepilirYi1cezSOH6005F1bbAn4vbGvwg0rRn3QBxi+f5v8/Ipz
odAIyYutPh0YzmFpqPPYJV7WXkxCwTbMhow6ejV/ceT7cd91xLKA9pYWZOnTjk52FfCkV3J4nkRx
rOKDIab8EaFZqKxRXm6sH0cxIY2K6XERHqgrrrNbJFpidEVmGRogPs5BaBY96g9373sKtCB6oBSZ
6Xrj0/Ga0p3BRm5JK8sdi1VILxuowjia2VRDJS43OeA3lbjYlCJmtYbAQ0ux5EvCx1sKPik1fZ5a
YVpr+HqXn0cRmS/j1tUPiSxFe/3Y3F//gJEMzgBznTCPMQp1PtKLM0Uhn7c/rSYul1F+BQUxTwf7
MQihWV8Yu0Ez9MVxV42uVaTOCNEjJeOVuGAhyfYt/LmShfo2loT+HpcplxrAoZmZ7WDTivlRJoP8
F+Cx9NQjkX437hHaNhjJAOC7n7uQll8XCFCgGiyDuK2+uMfg7Y5g+dB9lWfgxBWfsxKTbhjgnAaP
QmzB4IEVLn/1yUVMOWGVFPNy5fR75Aay/7cHN7f2RRUgxLaC3CJTGZ4Gow0jcJTIPQ5odgZE5o8y
wPxBK7tdjee9I9k+VQDiF+bRgZ7DfUzo5CU908IJDNVB8jQLABLCegc0KPntT+qRY3YU6jZySJ3f
pLYazA6t8+LCYimfzNV051f/YC4IEaQY1SxIouikT3PDp4B8XOcVjOGMuWi1kr1wa5yLw8rDBxzt
FA4i5PEVVq5bpGBKzOMNm36TfqMdeqYNNDpwUJf1MCAXm1ODG0cZeKEo04ijFUJzeYl4LCJk8RAU
0wkaeaJJNloyw48e/+R4kV+jhgAa1r748syr8NESsb4rqb0InpbjCCoSRQFCzPGW88s2xzV/Q0Uc
a1T0WJp994VZzM/RFPdDjGqLQmpcwxIvreyIVGIjs8IbqBrc3lmueqW9nJ97fJIBJodEFfoBUy3X
fzT9NcLF6Phk1KKUbEtbaryWck+E3sa6GEFauUxVBqpgRbrVVAzwDYznL7/N5JaOouWDu0Yd1qDz
Pqs1bN/rUFcMBuTsgy74NhIbTaWNgO1AGw+gyrBfK+4bny/b0/fs0zAyBUvjN5sx8zQLnGe8qHRB
xKxYy2/tJxXvSVi/TynSniEk7B90gG+rn/6DWDLOwHoYK1m0Ij9NIwPTrUblTsNuVfi3UyRikSAm
yaZRdl4NZB/Uwr8U/PTXeukOSrgvujIXCPkr08QpLYS1ZF1R4DMQNNo0WDiRgRSbPkwpwf44UvoV
hW5hyPyrqeLHL/UH9krv/gOwjoc4A/FjtE9dOMb9HDOwEnrbvhBszMVPmDOKsPAEXCJvwJMPQ5/4
oVqjEKZspsO+hEabTLiCgLdX/+CCFWZoUk0U5pJTbbXvfJpZUOLaKBu6Q6211KO3+IlFTsigmXM9
LPZNW0+fjQU4uDh2XCfEMexQ0M6VoA2rhSiAQnxZYC/QZNKiJ1JNaAjwH14SZgSwVO5E0G8JnH1m
8RRmEC+OVHiSagZtDzxQlEBwk9TZ4XdfhQF1Yb3CmpFrR9zaQyvRt/VRy+0FEu/dBKHCsEq0nVih
H2E/RqAuggdk0q8dqMc+2i6LAFtUy8nIxbVRHN23ZpNrwrywxTgwwQhnRMeNIvVwrbJqFAvaudX2
n56jhr/FveHmJXDlR8E0evr/8UaG/eKT7poqK9ECY8NHZCZN4o9Revd7EeGZhXSO+Tpr3rujvd4L
YbeIbHbrc5pqPrlz4mXZgKdjwZHFFGmRF7BxrFMFxA74AsloX0IyWJtKpUXUE31MkWp4r0W4ZUjw
aRekSimJ8tA4WmRGWgf7LKefqBviwCFNRPN2oZysIc76ouxo6LMP6sBNAcvVkX8WUgSy8PFKDUXm
b8IAZqI5YMlN+CyadoDFNgb0dQ5iX565iur/yI0U3gt7QMJM+coGQ/WDCPZXqdshCuw8nIA5in57
Ihx8yUIIpbKy3HcLarbXlEQ2s3E9OPV84BedInmsfWDlPJXbv4Ty0DjVw+OIPAF7C2AKFo2Vb+IX
RSDx/1kU2peOoXxMFwC5XtPHjEAMtNanrnYl4TtG2ualLGc+mq0qjO2wf2OMTDdWHo9Hqlf+jFse
9WucmD86y/N3eEpNydgI6JARIU+6poW/1x0ux4BONf7NYoYMVzc8Go83dsl6bHIvEIEOME1Cgw+7
mCVKMtEaqPO5XgtiRWcyH9YJb51XgtFpQrboqPyQ2S9zZgQ/VBSpqlRyGSf6qksinVFg72Hqk6SR
AmyBTBWH/ZoNgczk6Nc0Hy69Ftq+TPOVhVt1DCVGLv0OZlzUSYsRuOQvmuKqzVWGSXu/I0AWxRkW
OfgUAAnLHNmdmQvP+CfrEGWYK6MOLVWFuGwPwd2H5pzqc1RZ8gOoxVeLR2BtQKh1RbwMNH6MnuxI
qAg3BAdRsJNPd49K62m7Mwtp8Efc1/WS3OdxQX8pmNhM4JJWw14XzJqIHOpPJ1phTixlc5UFmbP6
2MylYwEGeblT9Y9L96Esq5wPnYQZvtdoO6NhC85wYF3GyFTkUOCzvSvvFFzOYcNUL9B7kkQOtEAC
oK1S8rH67jOxx2kbKRgRdplhs8WeG/KbR0tbLdR4FPfhSub5ogZmAW9AzjwM9gOqBu6Q6KyaWDo3
HxlLPXqn3vwgMd0UT2OAcSGvoV7CJVntezPe+gP5K36OpDpcTtoxe4rQW4TB/oJw+zUE1Ry7p704
GTOhNaJk3KZFmr36p6vjvMjZaIYLK1xvU5G8tmCubm5BDkC1yeSFA1MReMgpRSdlCbzlvcE3nsPt
W8aj9rm0ma7pGfBUtCdeDviQ2VL/yWHy6hIZtdmItapBMmkTT3F3k+ny0Nkbo4x3CdIg9oCV4IXM
DWD0L1DO1fHY9hb0YEDjxc8vaW1NeJ/wtHJ8594HzN62CIi1RJG3mhwmhzb0o73z3bMhaZcjkmZ/
9ri/KQ901QgIZ8s+23+6hlOJGp3RPRoW4ni1ahZzmDQKthJ7fqccWm4194F80Mcr8UK+RR0iwdH5
s77ERsfpXCjIarrvDgTPTwRcoO8bYs32RqiS4o1aPJgN3BMIhgRZXSgLA4bHttn7qIRwdJTNgD16
xO2KQilrGjRxUXJe4ScnK43HSaZEllcE0Rs/CZm9Jd0OV87LkC43BogX5P2UXVYJeKAUkz0i0zC0
BXqA8vl3RaOz+ClPQvBuzP+oGn7gdc5JwjqiHdbZGP0kbfHyNCh7oPEXZ8aNlmToZEnM7+zbWWnp
KwbN/vsJSB+AyCauJbOfHVa8NBd4RvIQZZ/U0zGIuWBchYdSWJR8/ja0EpIJJ6xf1UYx/VU4UwHN
M+wLCXuFyx2e3HJRztFV/tdzbfR/ht3UbuRI07F5BONXf4ylGIy0ZENt0LbeVUyg0/so9R1hTOt+
Cf0oQOG3hUV5Dul09OMh5HIKr/yR33WfyiwvkUwRKaxRnX2xlF+mi/34C0EpDPdaqfwUIMbN5FCf
D1upoDH7nC5KesbUVwjw9+VToQBaqukaen4XWuNiY5gTMkFCnE7Z/uN45HvRnp7yrnicNIHOO3lm
MXQtCZ7aCpaVi6WNBBltjx/uCOvTiI2AoQQHLe+yi6iN7JF39t6aj7j3SNGUL4vo+hn823M9oZVW
/ztto51SJT+qamVIm4e3z6oHFXw9iYdTqYNbjiGI5qQiZQbWFzYdq9KjNMhfeUR6xh/uNPHQZByC
VcH8rX03QUaDVnt/yBH87DjuNAuyMiun+AN1fLZvXSn5LhQ8v7OkhXUZeIMbihiWnckYGYEKg8R4
bDTjTeDAEH9wVOs63GRcX4woFG3mQfXYdWupUKaN050hZFvL1OZ3Vkz/IIGfE+410a1NG5d7Redy
K4STu8+vLRG5DRvHRXi4DF6ENHb+oFgLqwDwE61z2rEfo5ciF8xncsTi1fJRGurpZCaVMOmrErZf
Hp4cyXeJZTzNXr+CvQb/3aJ1Aj03Me4irH7Bz9OIpsysDaXVS0Foyxxj3AX2h5vyx9I5IA7U1fAh
bF/FKLXPk27xeFh8JnikSppHyQALUeYaAPb+czzxbLuDTzGU3IqCob6jOA6fcDPChy+CcvRiEeV2
TluOz6bE8n62WSbu7hRFeMS5jdQrDU7g/xPD5ibcptIhWQsRYCT8ITTAtWgnp3zlhC0llNdbbbxN
WUiKebF9lG0gdo49CsgPIxY6sUMxHChaio6odXsY5jUO39mU0mtAyhFZlcU4bNIS094PhVuv1Vq9
tgmOi1g9f97018mS+FSjjO9UIMZeRjt3XRwL9SGVdW36spUK+QAjGs0PKmcPthdTraLrL914ZMdC
35grtz9v7CflhJwjdX9T8mOU9WVfVxG+xS+tNQg7gdmhYvDfDmy+HNasF8qHnjHqSvwzMllTF7oD
qlVHWdnT81RlNyGDp8HzJ1H1ZngjgHJx606LtoHabFunntccYCuW+r0MJ2x1Odl0h+/y9qYTeZgl
ftIy3ppDfxb962ZUchl2ywrQag+rf0xfY9qgN3bOPjEV8Xo6illLxHYg0HzLB9Me1c0r4qrardvL
cvZkNxWwsEYokRGJBwRNO10/9dPLuMinSssSKYyf/c2N5ewGXI1m+d6ienZCqvxa90gNPaB8qvv8
9Fbd4sqwWvxe0OUorhYWlWqj+W4MrzyzV9ZSd5S2jV6hN5ZoO/Po3bhd7RRDIYZ8r+stLHkxEPi9
XLNiVfaRREd0nW1+OEViMwkvtiW1JVtvnvRbOtCOnNmfU7BoUaRc12UvWp7esGpLojmohfqOg2GP
+8yYFpAImiNUrorSx3OcVP3HOOkISV4IzhDKtAb6YGQuNd2q8/wK3n2xyXcAOuFi2Y66ywsf54cj
QIRcmuzuWkJ1u/5gFBhfAaGLp8YY8K3IURP478lBrL0PSyfgbmqowMuZfBSLlKCYQbxLlQDrcsqw
7EajgvkEmIRursi4FBRNtss29aq4tqR+NbfGevlvV+2FTPLEMmAuLtGQ+r223JLMKRzN5fnkVK36
FXSxL/fDIOZB/PoFcmn8y95jgwUQT4cOkBGffRO9rBHC8wXf7WoDVQiUOWmA2AmzGUbtv//XRUnd
9OVkhW+S3cQDBWq9XH/Ljwbnvgiu0MvU31aK3Lf+FOqi9+u+oz7Z+AdxPXRI+aqLZSHyHVNM3hrb
nMajDAU7LL4bzbc5CA4DRHTJmoNx1wchU2rkInazDbH+iMcsCHeaCOYpRLchUZBeiMp5BFC4+GQL
D4iOhSGzjE6A5IfO4yLpj6JHUZmjMN2QjM9WnBsikUMzY1LsKygOulXtWL6ZwdMZ1qciHfntcz3+
zx+o+lFEfxNDbDuAv85EV8aR5vcCfg4Hc1meV9k19ZepFQHmxsvxClIAt/QCKe+ROCGZUI/fJSNN
zy0y6qnfLD4XJ3mkSk1oXED6VqCLIVJKuSi2t2X3S18KcGfWD9wkXxYhlZR27WyuyLz6Ql4yeaS5
3zIqjVpdVrrjUhOrzgizTk0he1gMflOamrvrmdbLLMcoDPr1D6l/CVrdA4PNQMegPsOgmXn8ZYzK
dPXu9No7AXRTVvoE8YrXMz20gHUDR79DjAKR+lzxFu1fRwNeijNJgQz2/vZHlJk4weIoR844Oon3
zr0ulDwXv8eivmDeXDu3sMsqNKi9/Zrbzq5ZVcqGa6GCviw0yJAdFCCWkvcYC0tI8tYtLcVEdbm+
fu0ft30sQNQdFFinybAVdshYjPso01gI6Vm774+Yeu6m3a0rOhXN6HQ8zE++h1STxOli5C82SVyY
kTBKRpaYtOQ8CCCJed6PO6REB7yPYDtK6uV9yKY5pbGeoUTT2O+qS30iSoZ1Sy1/BOMzNzIBbBQ6
AmsxRbcGIiOZbCPQbzM1l9ecz5AxO3YCvGWI1ZOzZzozB4rX4R24ByPeMz/j/hEHF9jWLlir0wX5
oYjwx8yH/x3JHRQKVnhd6l685F8TzdqRD0uRsEh1eW5PmndtXYiZo77g5O8OSQQ7nqXOEYQfUxNm
SCRDcX8SwPmLerJ5a4j9wK1pJyP8accsE2UqRvRRmJcOmWmUP7YQ0w15LL/oeyMjcZNcYC3a5JGJ
YnRUeLNWw8olwOL2Q3MlbZBdGo23oiR41lEeIZeIHlyeOof4ZfGfZqxjP8gMti51CRepk+jEFdGM
bCgjcVRnTOrd9/y6jx0BtixnZ/QgS5RzKx2GNpxvni6roAKrURvP2F3bPjFwc5UpEQyryScnVDjg
+2PKltpxykkJxdMvj9DnT162iVRW++xUpcTFYRloG2F8i+hIRI2xyQqxGzg945wJc9axrxI+2FBH
DSM0hSsmufMsbOnPUrRE+Q3PuxHjPAtgtMGCLtBhsWn1KWWk+F4vfpMTQIixg8ehYnjYUMKc71CD
8WoJhWCdDhxFNrAU8vxgN51M3ebYpF06qetAiC7CD1gveBpOAqiI8biqNq17UTqEdaWlSdTFKTRM
T4Q6cPnKZcSsPiVI2jDq/YGMwsZrMeXrGSuH+c6I2tpHCKoXuz2ScbVoF4/0DmsPfcHmvSwaTS+x
Ay1FsqT1kOM8mf1x6Dv9aYd9rcZEF7uSzgD5oPQb0qZAMtauosGXJKC5miUA+kadWgQCL3+w5Ubd
rdQh019px7R9qonRI7w9fG+VJ3CRfUh7kT+zhvdzD0+JvWYZdeQNTjkioucaDHljwr/RzeCjf4vV
31Nfxavd55lUZl9C1LvH7L+FQtkgKPazFdR3uX88nV2SQRMyTgmZV899U1FK/8yUcV+21/RdSEgI
uq5xQNaHqiEo2oFD2qRtzL8wdPXpME/omPVNe3/uOG/EQg49zlFmxM6mXTQjk4PpWduz8toiy25b
Y/+WP6grQSZIE8SDqFXzSdqN2Xs4w3girCHdn1Ln006Z4e4fHKo677FFyv4Djx4EBt/CKdFaNV/X
jLBkkXtp4uAuXPMCa8vxBH2K5CZRmDqlFPkA6K26+h1wN+6VRjfTUy57lgmsetbKmEF8kqUAdmgd
6wINbS4PcC/KlJWCEuANsOQA2VOXY8CpaS4oAGXe8iL+ZcdFetAInrCmjQAXg8kEcoIIFPQqc/3r
19BAWqQCrVXgYPM/E9e6gi6dBybOH+Qq4hVtDzk2dip9G+xxCMSjoqaYaEsES6IAwnbbVN5VpGC6
u7gA6naWYTOA0jVyqF6AnpH6IgpVni3HsfQjM830hjBZlm1Gu7thR2EUD9kvqCFQ+qHjPIlpkGdi
6R1eNjxzGP4sd9adLdVAPA7mgghyyeWw4WA38ALA3tVyWdtJuOXY8CAk4zQaAZw4koxaJnTNQCRt
yWIgEWICgQnPliv7VrVrpCRSOLY9mu/68TLJMDI+po4V4GivxPlPzR8g3x6VfURnHlEtDz/aGtcb
offlBahk3uMMSW1f0R3adjiQxoLssr//d5qFvj3/Cq2MJswbC0KTFFJ8bqVHqC2DGO2VvX9eFlYE
GItCHSqCerDv4holWG/WGcgR73VnuIp1zU84EZXvM0uIJwKXNq09uFfbE+nqBb4g20T3zWwQ4JT0
aEaoqiUgeTCO3C7uJgHzegCKqbBArmIODWm+FinayGCMBdxE9xupadIo7GPxlyKW6I7nXTdMrsz3
mJ43CZ6MyNGpH6xJBRNFkfQye19Nf1F0lGbAmFqtZre5lxu9qcayU1XQJ1DFQ7XBbqay7T10HjW2
hwqVc3nk7r/q5fTNZTslgRwK7C5qasOsB8C6ayzZPjI7Yon51z16hUp47QRYMQOvBiZ0CEkV8hDi
qpCYhzys2mAVgtHqCBI1hf0RGJ8JB3dy3ka3MRpTUZo+Eb9aIqw37qzYWa1S9sB7Wk6MmwbvSlgW
QyXqm8BB+SkXZQVQpMzHzaZGubL7cFYSCxNzaXNJJw5TJOCeprp757Xt+DSigRo4pfOU/VU7skVO
UBIKlNW23CqniHRq3INOmB3eI1XCuIvZxTFHVxKX1hfSPbT1iQkzLCbwAOJsVPUY23OY/ghkth2K
HdwrZ88oBI7RjZtEPHtVgo7F53p8mORP2INEIMGEjKXqx1YTRmC5zRMzEYMQETSvo8tq1wAg0FZP
yyf8zZmuU7/BRLrxDtav9dO5rqvzuWjDqbgTW1ygNzuc2v38BL24IC8TlL/KzXCmoYZlxoUWdw+O
BL1Mk5sHAYjjPWJgN3jgRSbFja3agqfjK2zrg80ALENNQEOIbcyxPa6d+M1BzIlaW5UOgBnMuo8l
YrPVhkLEj01gmtDltvOVtxbPOw5N5Khqr5E63LDqBYpsV2JaGcL82dKwLqg0f7Ub59q5OU02PHqZ
fbQR7U02ZhFO57fUmD1/bQ/zFcni+o2oe/h9oas4hyrBWpZx3yGIBmelzQQ0L1lTXMqa9ZPdg+W4
YRHZGuoq3UtAnz0EPIYHwaaleUx7WaDjF6FHaWviz3hxJPvNS8chAUtGSSUt36upvkyfW4+pbci+
aX/eA8o5IQyg3mDJcpQSVmvanrxxINSmYHOteF0ftr5ewAfEc8zNA6Z7BIQeLv93oyHCvGOVhIFA
CNGjMtDr0vIg/wQE23Ecf80G+/x8wCbfcjCeU3XDY3bHe4bvijbIjxuLDqEhbRJEg91Gx3XlWrty
PBYPOxJsDYYXYoVxYcDPK1LyCSIfiqkbEl1Sde4Z67GgCLjZ9idptWbOungw6pepCgCAXrDgZLQz
DWGyZjvSU/YFnHeRgEdW9m8vKACV5fPqbZqC7fUJ9YDuqaLsrDC6HS2wndbtNDj+r0wYZUbMb13/
rHI06T4kuAnmU2hcpBdVkE/RHB2BTUNvLFZbHZqHoz30qXIgn/Gs88IP0rWwSUJmcnTb3lB0uee8
bsSgjsm5/IdtxwsxWVquxW9Jujq6sMt3UvrSoYEY6uo5WyMd375jc71M5hEfxFefuFMMAP9t494r
FHSxDL0kO+McgtmwO1bwFKQh5mgwKSnSMJF7I/oAbAwfdY8yffADR0KFIQC4iU7VU8BdzuXwa+Tb
69+4p016lY+tXmf/PZr2uWj84rwf0l2A+K4fKMfA8KE83JxZAyCQMnwX1/Ti4WnAXE8ldosuxGcY
6AwMwcW9EbUJ+bbmnYYP+fDM5tQn4JGAW3gM8enFWD9U0BFvhvbtjgBOzCamCY3cmsrqFwO5vlxr
5GAqJvAFocZQjILEoI7mFSpU0c+vuzfOdW1YByVzKVLxdxaeVGYago5/blvyhkZ6IDgXqQdp5roW
dTEQK9jMQ2b45wFUUMoxP0lolkKR7nKAnJTbssI5wFDibWGjxU7bbGwvOZpD7cvWZMHQV4mnef7d
VqkT9TFHLIU0BPhk41NNlxddglNOTiRqSSpWlWhQhsVqQmLy1CVndP0u+/iO7BeG6mp4oQBwYkWn
qgd3ZNmxOg9cc3nsXIgMr2nhtsbCBaVSbdBzToCadDm929Khn8lpILRL1WteXqTeCkZc7XVph+3b
nXsluVQivxiaTZpFE4oBOH3oIUunyjdp7asxkrKtTq0tbHTWuaDk2JqBFoX2hsOql1RwlGOe9BbW
KupIsLLY4dIK8ElBN/87IBi3IQ+fIvowsfSIOYOTGnfoBu5CrtaB2d5Mpa9eBMg6EtwZh38v4kcq
zicmNUMNd/WJo9kTQvyo4AqbGNK2x1otcc1MkZk7lcWRiQhOOBmAqcyb1EnlHWrmOz7/KpO1D2PV
pzXYOD9R4gxUCiKpqvQzC8go36Cw5a3cEbTcD6WGiSsoaAlxjH4UCr5/sRHbF3+99cuYNK37upML
p8CQKwUcBnWPTijji39uqOqDOYW5Nwc6PLRKodCuWY0xREAfk1pDx/MI36Wxlc7jZQoVPufTysg9
+iB0Xu+WmBxBDlFKStiryWrrEnUmWjejqj2NAiTTUDhnog7GuAhSiPkTyn4MHy/oCus9hrbfWYmn
sBB5JQ9lgxFr2p5rt4t+XOr6LqpU2NafulLum38RDrX7YSbnh5gqAT8x+UWGfP88Ok0PZg52y8f/
iRUQPp/d4SS8LzTwN3vQl+2RzRaE7ucHlc+KAzX0RymyMK56bGjbNplbtpOf5rT1ZECF66ImUwn7
1nELrB89FW9aPOLgwPjvlml9QKzPSIDh+oe/s5Kx54jSW2BJUCdsy8Q8RG0qcya8IDyRAHDw579G
UiPwELhIu4OYKPH0hJjsZIhU/xB6Bm20SMyqDr1sb9yTKzs6iIJ3wXfWyksT4Fm/U8boKL+xzNwP
vNujnMfIMJdtLz7jXNUWpOChlJxTDeLlulCBodppn8lYY/+o4szG1Cb223S6QLMo2inbJvxiWT89
FAOWbQdLXlYtany6Ue5+IAzh5c6Qqp41JA9aDWZiY0foUKm5Kc1cx843RO2L+3lvfNoK3YNFE09v
LaKugAqTbJV6ANoiYw3N+xRhs8qLU8x3Q2xJdkoxYhlUTi/+i5TQuHVVfLES12GIS7r5Oc3JcUAG
0GBN1bihhzxpRIWVyIXojs+WmpokMNW1VxPKFZQCYSz57a+as+0fbuyclZPyYH1cuO0IdqjcFfnJ
QwsSpU9IjJnoZBrZXs+CeoVPFAmqxiokjf6G1W4t8j8g5dPPO4WIuvElxKrn5j/sK239wwF8M6r8
bZzuqEZpU+Zjar7Slg1iVnFnSTNQVmmcBijr+MonkanJVLqltPpWMDF2GC7UBuwxqInP3spyM2gA
s9scQA4zyFcd9Ps26aP093nQ7euniseaIYQNgd7gZipWJ5k2QXLiXKQEOE4wxPgUb5g5sz4dST0y
+uoE4KN3GsNaQfrbdXGos5C5kMegKv9VnHyfsnQ+g7f3aDeTAhLywJBZVjhdvu2DW46cg2PwNyAl
w+ZXo9soTMmez5K9sWdnMtWvcA8TceMWGNiq/I6TqsvJ+voxfulRuZIh9plryGtAJG1zajfs55P9
chDiWgS3ZB1tqc1dIy/C44yuNYQUHpTyQq9IZuetwBv/1qem9KXKZvyjz7Z/NRrakKMssFWbqU6b
/JE9iJJheODRdhr/YohcU5YS5VQWen1omQWLte55OaH+y619TMjn5wWj65FKliLqYWNv3cICG9On
DAf7/2TRWk7oWNAlB9cXxrdp4bE+FQZ/c4avECcm6SbAiLwAmB1V3V7go/jpHYXRz4SqQ1x/KUv8
8BH9za9dlBW3lZCnL+wSxllvDgVpa7QMn0gqbgTUtuI3JHN4aDLzhAstAYBy2d4wULIS/LUDrbnT
0HCy3TfGqPF6k3ckpnbHmuwmoNERq0OYXtuG/WBO82zUL1OLBGmmPtmiG+Qz7tbpRTzI+GFBq3lk
QEmOAgm/0EyOSKIC9GYsDe6nM7GaTs8Tj49zrJ7oEXbFvj9rTORMxSgMkqaDU7SjQnqy/xOcl9IR
AYHQ6r1XbyuTapxMJh1kJFKOUiHWKTS3pSDOOmU3k/465Z3ZQBGeH13evSrO/7osAxCih+vy/YoU
Sc2xlNjXHNAezp0CbsgGb7tQiIcmLeBHqDDmIVK1HFMKEK0HXUESgI6NbwhhrlReeXwXnzydsAyt
sc4jz+Teo0oc3X1d/Bra9yrTtmDzoQHbHdnbrZNtcmUGu8Y9qi55Jb+buixkh8Bb5nYyQZK4C5cl
05Zgmk7RhXjUAu6K/ygOjp9L6Cg7v705wOH1BBA3KPB6jGRkqf2RKKWutLqcp1EF1UzPu5OdH2AR
bg/RCPPi5JrdqNje8MfDqYj7Mdp+h8BWJYCVYqFc3mlQDIV/wfqnBEFIKbZHv7uwIjV48n5aKd/l
uXFV5XFZOKV0cvVWBHQH/jTrryDnDNSxE3c+tkVLEJ7/STdLBt/HPXFIGpDnART208J5XrLzuFL6
yImUruVtj+ZmiXqQVHhesVBhfXBVzAmCFrrm6qC9eXTCZK+StLAa9m7kAkYFPx57P0Lch+T7FcTO
+YEAaVebndUGeicdDH7EKmD6+TJ84wVgdZ0nenLemawFSK0CHAm8GRm1R1psDf2JC/XsME5o4MGZ
XkMkzdfu9fUq+xD9AsSTKfc8stmDJlEv4KXrqPJvOOrVxK06cKBKzQCCg2n01eNd2sXR/xNQA9YC
Is50/8pJDnwn49w20hApHZGxdBPaaefpn+FlHvdG1dgDNJE01HyQYCV5dq/bRXI9snDFdO1W5qGo
5ikmyYrCuF3Nax7ufKXFnY7t7SDCBEJ+cEBVGp6V7Qwj9LS+hTBJx1WwBMQkC4i2CgPZmE7OupUT
iWKb/zS5yAKmFeztWd9+ejtOGc3suut4iZAIZMNTYio1/53hSx+q/soCHE4pD0mYJ5zcH+9eAKcc
u32E3FIvdo/3Q4qdMMo7ajoXDr3DAZDgfLCs1561VdQMoBbAghEddPX6DWT/W7rhMzMt4LQ5lI/k
HL2HzEX1rG+S5ZW0jymyzL2XOiub86NjmkLxjuh0QtKO0msDyS5hfSPiczHZMl+JrfAh9X+EIfcx
pd0wQx6qmysN2bVzt1MqmKtprbS0p8e6jclD993CABVjRfpjih6tvp6GGzJt/BUL5+llc0BQNpyA
SYrtO141FMoSApXpfnptybZkshclSSasdDCfHD6ZUhLzG9DIGnWTR2tYp9sDp8q7DMlxcWtK117i
jB3qTJlx/ondDrz6H/R8iIVA9gshkWPogyTt9KIpa/+84WRHUvlIAJJllFzTfRg2b4Sk2bekTHLF
TbfoAp72vRwsA7vkd0FOXO8E4/dj4RLfARc+e+o0DVby1vaxStqtgfZWWLg41neaG7JhJlTPXqnj
ZbdTKiy6HvGstC/Ipg2XbUMN8ZDSyQUFZ1cIAZCGDc6juTxPZj9S4SB/Gpe/nFyihA697gPZO9kK
jNp3ub6h5KirP+AdNWAJLckJBH9elSXbNWZjwZAlFLAy5kh54vtLYpETmFGGSUrtVPPi2VGg+06Z
dJe0zcuhSKU5YhmCLOB31AkmW7niB23P0fJHMlGD4W/fHZoU3C6Lkc+0y6LvNbqAmVzd6COiu1Ml
cnRCacYJuErnLIiQiXFjGi55QEep5wXZoHgOWNi3yiRLyEhN14ksL0rSjlI1GfzWg0k7QHVMXelg
Qg2TtIaisVkrPHZ4Mn2PvnA+f3dfPWkgHyoYXj1y53DLTLZTQmDvPGv0tdNTgIvTL+ZqEa3S3bcp
W9hwKoJ5csWGyfYEOJ3xn82PtimduPmliDKAjVfkSpwx8Q/Y+r8B1QxsH6j3VyStBl7Bp+C6CfO7
afA7cBaWNjcyy12eaXLAqel0LSu1sG4flkMkSvxUNbNI2t3znZPQLrzQ8JgbBSBBp0vsy+wflUP8
7E5/G0Vtc7CGgg/TP4EsxqsSGhVKquWTGuGEzz8fy6CxXR2MYlqPn6UPI2c4pQ/qgec/ZUVccsvQ
PTfZb8gtMB3PUAxx6RBMus82WBLexudOwwfTKITXthCBnNDGfpXRnl6CU2D8sw6IZTGvfIHtz8D9
A78+xSc6JmoGRt9WyGiVhZS08aEVo9I4nmsglgR8heP4INL3CtosuWV5RbOuwJKFQWLaC12FlvIG
tH3ZaOLMZQGFWXbtsy1A/Ae5iAJU4G6o2BRFgZ8Y1uaSf5aIOCgK7D3IL/QlzVhK9dDRPuZ/bjwp
GLAsGyJUnNw1PAfto41sqb4fiSEX846hL0gmokYNlpzjhBMM0YCRc5GxfN8swvmwOGL5aEDw2TT0
xRE0Q2EcWx0guioTiMtOLznQNB3KCxo2LZdJawAGdd36MuM3A7lZiV+VnD3sKeQ/H48O85taG5lf
4VV3q1EcIlg9ylWq/zjnzJDhQyitn9MX2fqY86efSlybAAfcqS/8FyyWt3ovSwVQf/jNg/S1NKPT
SIwKNRn/GgRSu3N5r4aMfd1n9BozgV+3BKp/k3VmMMfsqB9wURurWOe5yAUsa8sUMCr9lUljHKww
UQnIEt4ya2lDkZJLGjFOMEuLsKpcaOwcoYr660VZ3nexykMwTIfZAxpOP52jy6V/rErQK8Jz+H9Y
wU+rl7Y2sK3l0lSP6BA2W4kmERXOVxE6JwWeQG/0dVu37aCslYHDQBNrAl53QHChwOpYvklOlc5B
f9FaSvKTKQUovYQaqbMhmH3KgwhnDGx9Jw6yGT1XKx4qWWbZAnfoXTbzxTD46Dvo5c1ntl7oD/fW
+7To87Kbrt4aFShPoh/SYzsqAHQ5SPoTkxNaTLgm9B6l0aEPRNW2p8rRg7xwsCi28nql8wXeHGgY
TXmg+IFJGE18KgskbgBndzqT4gscSFYGnnYQNlNxg0Bhjf8lRIkAKodyODvl91tG6eHCweCnsrPg
3d5Gmix+QaNLleUqFl+WNOC/kNUhM91jgNTzVgJ7am2fwbLyrbkwcFzNfm60eyIEJNIezY19LkNv
XCjUkVvIay2zcuT89FBYn/CubfKdeYsHrZxVOJIrm47T+V9cPIcrNI9Khg4fOcnu03TPQnpiq3xZ
3eAUUQbSlByZ1BozR04mQBQX5isWTReiaitfXdt6TqtfXKvbcxtjB8croxRDqjD8nMdf0M/skaq3
dO2TWH7EPGiHyk6a/I1UqTSOCN5PdDt3UHfjNz4xIPFYE/fa+akSaa7wZrPN6RLTuooDxnW3Fc+w
tfWQ6nh4t71IDNAHgApgSZBtAs4K+2F3YfuVlHz4H/pgnRqN7sGyzYjN+cTXFw0y4+gScBXVv+Ij
4ZMuGLs8gjMe176U+n2RluPhBZi32ndJGs2UnpVmDOQ9a3TUqNrNCtRQHkG0AiLLyzz1pT6J9oJA
GWNaPI0OpKc0SAVG/qkUSoz8LHheCbkQL2Op6/U9/B3WCkr90NrKru/VNxIpgGT2MtqjsS41Nb8C
fkJ9iLImjXKfvq6fEvDquZK/RfDyYDhlL35Ea/+k41Vtb+XCdewqmSZoteGBmNvfa88v8ZsJ+t+Y
bCD1tMo8dpdRtQgyUSEZsRTwdRLBqQaW6o4193bxWWVm3mLqgOd41GpBp3pL28MEfzSJQAeS/L5p
xYt96BRDyLDW+cRpcUsJxpI55G6vv7WwmDj2Q8gUw0hJiU2Pmeam3JHNmjJ1gBa5ZSCUeTdCDw2b
50ygakKJtsduGlS+C7paJulLVN7NuwILWmAe6zhmQwPhJYx4Jv6OQGSAkcYU0zdOXsAptkpHhy3R
BCAH2/U14u08zIuY1slCO2SoKxIpXDUqfgy8UxKn+XNc6+mkGz/O1ablEk2Zs3pxmd0JbGyQOotL
pQnk1GISrYMBpcDHKmqSGHTPA5LD83oEoRy2QHyptZRR8eMHz/4o6dfmS8xXUlYqvyQsaMomGE2g
dv7tSHMahHIDF4//76yoOsh4JlbqTTxtotCeeTx68M4ty6qS3BcVzyaqLvtpBkkiqt0hRDRxeWp+
M3WVDcB6rmefOh4ah+9vZ71uysemvHYanYJuIGGtpnWGbHUdLtwQV79mD54zolWiAHQvk6yz22oK
OrD42IwVe0kvcBbG5rLKgPOTGDjURWinUMeq1CJtFWE84kNTbT8N9+5VhDH4ShSlKO4pJmMhCEGT
69oURk6jlzaiKftNOm4IIxqUx4iBA6NN9bbNLEIxgxiOuVw6SUlEW6eQqFdTlFF0pDFhXEAOeINq
Iv+vH4km9jkC7bA93vOOf2X2buEGw088QjhruIjJ8CjH/xH2zhziMnCgvB1rYJ85Jzur0Q8egmQf
Kfra0gDTr5s4dC9ZWMSbjyH1LXr9KONNbRjtle8+bs1SjNF+ZN4Xuj4Jk+dHNfj6MYgzvoh3cRdv
VQfogNICz4QW5ZiapAGXChmVbmhdjrD91uGjCIAYy6SNhypvJoDUSQ62kKe9jLOAavhvxAh1jKwG
VAfb0NtgjPmPc7z1ct6Ub70Bk1/ZEjdtawRPsyt1Bm0z3Ul16sRNZqubvWWDz5/T3PVYwk/NoBti
PAiXPPShO6TBsAQU+037mijNg/4t80PXiovc8gbWR+ZXfLtKstt4+vXRqXmzyNvZthHqWw+2SB6J
Q2+fF+ck2QzxhpOQ6YQ2H2DV2ps+n6+5+SeW4sakgx+vX+X54IbUQTNmtJL1Bk6QMGHhqup5ZWJT
SJGaVLVDscIPyg/NjGbNYG9EblEikiPtkAfknelAQAugr/v+isKjIqfk73Haha0+z4tIl/Q+SZzd
Kz5/7E3AhvFAQDk1SgNnk5esxM0BY4g0ZhlnlgO/ltWGyvaePL1zk4T/yvEY+OwJq/FGAzYOSJNn
ujFc3mnqoIKUA9gjdx5+PIPh9l//0xMtioWXjdCRnrBqQO566dnFC8ROhNhcsUuDaFPslYr0hhVw
ct7x1AasoP3CV+3WXEhRsDYYkFQw+TuaD3mzzthjvCUxJ5Y5dTlijWDuc8mVnjk7X4/FNekeKWpE
yyxT/jmrwIHHjrkHEkeSerTo1cF6NbX3ys+0MRXI9OgVVeykfPEcPmdMTEee+d3I/BiFypGs3QHg
6EolQfaGGaYR3EmGFa98FOQsj6//MHO9UzC5kRdGc4bpB6nsTl6YaL2+6/XkXQIQM6F/qWjKut14
AWf2f3bx7XtK7Dvlv7zjH5CDwWc39hCT8Av4G7vD7Ap8qcsCeRM/xoNwvTOmpxE4+JPjXxkLakTg
LKFth+GZKiC3XC3MeHEyzYihLICCtijO+UV/HxIJ1FiJ+wN4czguj2mA8pj+IceD2SGibuHmpCJb
Gb+ymAwoFLeoI9WRh7S0GgsaWvqrFKTGfA96mOaLVeP97fhpqElMbJ5j84wpUuQ7pNmIJlMcqLzg
cZSjwMAL8HGKMvWh2Oq9uxceaNGw69BVcBBNeNDP+f4gA0x1C8jDj2ey9fhrNngl5oIlRAxlK0de
ZLGiPnjvvk9P5akqU89N23JHGST4qcJoSAiKb/v9TTpGQOZhJrFkzhnL4+3fWnBrhbk/YQ5LXKNw
HMRdJcll+e+CYmX1kQo7x97F82WDGX1cQCjWdoAilBq/9F4jCcxthAKvB9mshzXgYK236BtHdtXM
vqNmMLSxpbf5XQ1TFeCv9HlyxQhLmRmLOnVWYUQfF4oDBoksf+YDxm/mWVVl+7DkMFFkAIrc1+RC
RaUkf842PsbTBhKP4HoN3dzTThDvmrl1vLCFSIc8botecR4g7kUJ7PafuC0Px8LMqzdabvO491Uz
XRroMEiVXKpX3LCtYlmUPPbfpGo73qCiAv20/YwjhRa9J9U+RuvdlIRcqyHsvySlF8rEABPq6Ipn
cqHqG5M9pZYZu7c02Em1lFoODId/vp/DcJBSIR4cWFxvSdoUDgvzvxmjRx6Uio/RKf4DFdqDKHMq
JkXX1T8ufIW4dwe4TsRlsU1bav23nZREQXiT7TfPUF/3Jx7EAes3cfzhcyOIC505jo8zVG5dw6k2
cxJuQ04ZrKrPoOttA/UvjIwY5sS55xphwKYDG10GsKsuzSXKSvr/hjwhYYoIrjwLgWqQsj8OUSD6
xFgRI8ubT7B0bjHrLVAi6aTlfDdwn5xCrRckCJiZKU2o3LcW2Rmxv3awiWNWoGrpNqvvxqoOtQEB
azTLRh4eHRJJiF56p0JynvrKm3RQ76VO5BXMtJKEYqBV80frv3x6+nbWkbG/MptxQjLhsFh8sib6
6sr53Lyx/DSU4qOF52t/Kc0RK9r7FTnDSl7XSRtk54ischQ/NRO0KRmzHEJ1weh5xbFwvlDtgEZE
cPgGXF1pIxekCEy4WhLVBrTk/KAHNHpsRCPQ6xssN42HUD3VfBeP0St/2qK/G9BCHU7LPcX+/nSn
hwSuHVzobl3TdsY5OKCi32xmSdtB/um06AZJnADiJkEJSlwXCOJXOIKmPp0Q1THVjEWT2hKBRobL
qABK4atfQn8o1cWj8li9q4wI/lIYM0tBwfDHgfCBrnLruS4gwaCEt+sviUV9rGsOG1lEZOLtCg+s
IInuW4AxLwnKpxn8+oKoH8Fv0/6f44wesn5XImDKxyESZTQ+XqvGaL6STV5Sh+MFl816sqOTA6DG
QTaAHk2V59YmUDWy/uJ05Xr9uPVKrSf6A5XdfNP+G28X0j3Lolui1QurQ79WOuaH9y04pC6DNTkB
R/J6A/TWWFbh3s5I+OOQXoEogJcLFWVMubsJmzFpWT7poQ34H4Kap2lgX+SFk5jT7fFejMhTcGkb
GH10jLda8l4w4uhcApKxwFV0ozQIRIUTnQeZaCrv87Lj60lB18y+x2v0hePcIgG3nm8v09YuCYyQ
s9yv0rec4h6miEnwOqZIOMoeawU8tF4ysCA4XNLWe2sdsCVI4SjygujNTZPGLccQJsdHBW1JCHm+
eWtuj2iH22zk5/GVGnEvELXnsJdXEIE+EJD4xukRUNDyKs6rLKdR0BI0QFjKEjbl7TBR4e85JsYS
l52AuSmbUXVllTuJuw5YCCRh+ckHMx/vxEg1BtHkPKlUDkKIRscYIM3lgOGnBqvFeNzyhguLtVcb
XeoVkUbb+/kETXyeHbAyAKKsQL1Yw7lItzwRgacprR4v4/We2L63Vamt068WG9G/l7bKWuoYLLOq
mbGXbVO6Og1WJAzfH5ldoUuJsLLjtUqoeKf/GGrAR6wCfrE1JJnaeM1P4AL4LOD5N7JHknKiwwr2
gthBABDHFmASKj6wXxKbIb8WMcaiYegVyfdas7ksiTiI9pKd4jK5JprKpSYsKu7RtjUNSnLswjHX
933lxyqdPsSR3W6RzkCccoP2wu96QdHWaD1SM4ed8+2JbS1b4SvRqJsb+D4qkG3Q6RJDFAoqhUtm
MOWYOSP2x9tglyDhBCDjPv5XpDyMLwgidg0gzVNnO/rNl+rYB0o3NcBYWw5/Eyasrwq3W1Db5+i5
J1cZxUriX8JBoeQvRJdVcvaGqrx6PeaA+FPKdADLgUjMUQ3+29efyVh95VVZ1IZlD5KSooZV2y2E
pE9a40QrHe0fO3TASxX4g+h888bVs6E7EoPu+YYInny+v3hip//Y/CTdtkNrXwP6dYtjHG2MYqkk
l7Tr8LS358GXaQfzgel8Xf+9fS11WGwia5DRBHPOq1ZCsePUnuFVLV0CLyDPh+U9ahV9QIH3v+Kn
vmg/uNX5BFdZmIZ/mpzAGye8jSUWHkDhJ38HaZQQDo6q5BmjnJrjvqmzY8fTvWBjkM464Yu6/2O+
YzbFJ5qdAlg57COhWhM0C122z5VbMszqqC8CeuTMhK2GW5neyj2X8p0VHzXRoKupNyYJSFxFbwl7
lNtpuvrELG2ecqLXhFKEk2rnvzysRoz8DOfV3FGQAFftATqLy3b91N6ZNLPjAn8o1l2ihTHb09u+
AUigyPp52CDalIWiy5yEHnbsBH9UUBY5FEoi4EJN1g+Qm7cIIu/n3xzPbdtUf61TTAM+mB+CNUQ7
AnF6hTydpkU6m0FLieGFon1Bb0uaCz6hHySA3qVXML1bkuj23OgBTNxNEygRU1KqdwC7Y7in2q8V
h7rvmhKMof0Sn/Wkf4Yj3vkddI/U///C1tV6sL8S+NO5vT7Y07FKAGx0SzV84aKQ8y9I0Y9LQij2
GfvzVVVZcLanqBQPIHPPNEq5UMGFMf+PCaUe9QTAhH064pPDQW2KKyvz/iM7NSbNSDXR+yS2SGMb
wlU40lLrLmHStGol9mSohqZ872rHoQhaCHHaZd8U7WYprJRpDmk6dFg6ud79NojokIxgAL9THR04
oi6SIHPgZFUwX8FWrHsUTpo3UuOZ2dnszaAuwpu1TFsvI7iNWej/FBNXoi7KGgD1sDwJakBi9+b8
LTH/Vr0XxttThljWJrqQwksLheNnApHoKHkmVbzUCyNMWuia6aIivMGEycU2yPbrVXKqECdKrKnV
sAU79/DCtznY2V9ejg5qzRBZA5sd1RUSRXan6Pah3xgyaJNZN2FjdURWzYMhx03kPHOW5BudG1q+
HAdn9FeXAHOZMJ+8bQrwDF4T4zOib8w41WFxZZi3EB0O57WOgl9chIOwXg1qqv5K6i55+5z3BpAY
LOvON3eGAmUBmtv/J6KJFJYAGudZnTKfSObZogPcVON5IGP1R2ZXk4pf2MNdJF4Ne4PdVAi9n01t
kD/IxkIDxNSK3MAq6ZQvU66bfl9KKCfTrgrXyhNqoKczqcCefoe3AOOwGeWi90FwEKzmkbRMnjj7
APiBKnk0R62o1cTAF8Hu59PpSWyjJE1FObpFwywmCA399MOmNohQYHBuiHoALNQxMhl787EyHy/p
l4kNr4ZHyY7pQqWOuVSDmwXPFbes+pP4pXYJ1l992b01vGxLdXVB58pcBm7khUMdEohcBkwiEY2w
rPyCqIB/04jI4jxDy+zWC/644qFU49qdk/gyWkH3d3BPxC3bZnFEf/jxdvzxW0b4HtDgBWVqux8x
xBTPssZv1GcPElOYiEact0PQ5WU/yH4qnrQIgK8PU2Et5km2bbvO7Eusw6ZNZu8IqnA4U5rT+5Da
rbndmtYqMOlrOfDvFOk9DP2uQE+RpzKjuqo8ptkBn71iO5sv0oGmfMfbPZXO7nGTNl4QkTl2bABn
V0AwWwc8R3WtgDzvJ3adFaiY02w2QoMpkD/aFj9VKekl214BtGeuXegWr6EoI69zgrBsSIh8wJbo
iomaVzJfbCj3Rcx0lcG0qM2cn3xwknSD7QhL2jt3Lyh0rLbjZau911Zz/sL7dfHk/ynIlRXqsXqT
hUf+YRpHNmMenSueaK1yDCma4Il4ZoscufPkIolOGyCrfQDgaZwDLqJtbKiMgNaaPwwedLL+MC8c
/flbW6rMvedP+CgBL+dfW+sTRDRRxXDHdoEw1mBA7upWfv3d7rjNr8ws4qdRAY54C1rYKwzCo45n
UnrV1CU/nDs3H8DFRUTzXCuyb4yYnEUyamyw3YFpSP6Nhj7/SSmqpByPEgnsxJwnk/olAWeyRYkY
SA+hK3Hi31nR06bQwZ6neKSVOdCPF+QkvtRAk4KIJulCt7A9EyOcS4MrfS3L64M9WwTaR+9pVjAJ
w8V+Nj5buZ04CmuPzHMec+zcCxm0iyHuM1BTLviEN6qKVscRyRoHDNQ5X6LzYVZbc+gmUapY50zl
dCTJ1OcHLwtHDFuQ7UVIMIadAUujTU48CO5fuL2J9TH3WpFtTUpXH8HIEmv16aYTBaCxDlKRO2Rj
BpKTTUh4LgWvTeLEuJPIsEYJOdkzhy/tCooE86/ZIMAqufuq2D54abGNVlnHLPN6+C+0kfxq9oxC
1IRX+DHu4ZmhUI1wIG+r9vh1I1NWT2lMyrkjwpi9hTF9dSbvOzJQjpc0H5Kkf3zNp5BJnJ9tH7pe
0qCIUqJ5E2E2Zj3wQD45tV01s0OaXBTranJKIAefeptjCu2R2wW9lHC3fwklKHoWoylULTQ/t6M/
nfDbFTjQ7pAKK0DbK1kjfl3soT+Bf1naAWv9leXaK/Vmrrx23Mgp2IIDSLv/E2nWKH+bddcZ1kcj
bgol3WKKA4GPKPE1jMgnos7fgkzxitW14ahNTB0EKWFWVIATvg4KX1g5oy90cPqe2HSi4gH6Av73
kkVyBcoAjTc7eUnT7udQ9Au45HV6VZUfWf/6cAD79xSQWpRArHLxExeV/wm9kPEG1IAoQTaJWdOw
Nre+jkrX3A//q2hScDCrvRKOfUPzGBB9pwGdyW38KX+krEU/gUvcwFfjbBhSRIQZOXY5inwPX06s
PrOL2KUkWtXezJcGo4E7YhEuSnT5iPhBtWnfXb1MHPLVEma2EaFDRru8zq2ssXvhdnj75n5K6Cvb
uoE91utPjTKkvabVNfmacshHHcxmc361e0LDyQZ78Lw926n/p8FTVvbTehV4AxfeGUNEF3wSxtml
U58ui4dx4ig2UUk+bv4i4CtpcltZvgegz6k/c+Mb24X6KAlsW2sRKKuD2epEES9b+O/gYc6vCTo2
RsAk5tb1OJ/SOeSdXhXfh3uOfpJc54ksYW/M9D5Be48I66x/tShtxpfsLbdQyBX8AH+SbWFfwquc
mkoqkemBBL0VHzbrK8Ik24yZXdOxB69YUN2SwszWpzHdwLIM4eIXIciAK5QIvkzZtyoLYyMFyQP/
XeXyHmFihl9W71+18pS4HpTOuYPU0TxAObepXfeUESUfMASoSn26FDYSEW2DdEThrHOL5OIe1wv8
cpNv7fif/iS7+sGnUGBQtLeC+Pg6HD8eF/XesSMxm1IdXPeexqOJhdFe09O3FK9m/p3Jxsvm8Git
kt8BBunLwzAnWNuDiTtIFup2jnCEYMTs8u2siaNPNmGixMQIAVr+eWmHfixLSA3cokwHRUNmVSSU
5/M0SNVbEZMHX2/WC+o1qrGXXk3Cq+Jv3f4BcSpOxKI+s/Hpe4CB2wv+cYk7nmdjYmSpYDpJOhqQ
C1IeUODlbPLMgmDUh/f5k00EsVMYMIKf/nJuAhgMTQeLecUArRk9CePXGhFWhcEPMdSQaWtnufCj
T/mbFEKrpILm1MLn01JmThgyYYlC8w9DUBJWV+hdCb202Q8HEJ/P6PRrQjEusg6CDk+0oZUX/MRs
XO0SNTd0dFesVVw8OECUP2yrPJWfBcDmg9WfVrAckO4nN2WuzlROWJ8bCrbHfa2pf3Zk1OP7cCWe
OE1HHEyZ/6wl15gJM5Qo5YWmmZPpuh58I6AjiP05DP/ydMwNHXPNAyiZ5EyQt2yxLrbwsQpZls3K
3r2QOf5hep02M3CHMsu1n8n8W85TezNHiraUSymuhUKzoLY4EOLRgxIiLDaqZLw8JrH5eBeL0V+J
2Ymw5/G0d9K0xp9p668qknHI4rMLUU3kRFRHqpwl57YKNHr0hshNqu9rcWEjDXobO0nwCDlSqfjO
S4qP4fUe99XnOE7GiD76jrLooDkC0y8H+HZP+Bq70cNa5kHd4227MvLLkzquWpG+caCVJyiiXANo
DChzu0Pn4IBS4o2w82xTeuFfmZrMbJelKFKXvQ3zl/vzZwBrBLlQvCAigt+m0I3ky5LxJrRxuWnw
diV9N9u0jcAhdxyzZXNIZrGTskmU4guqp3Au6OqkHKl/6NFBdowwi/8xnYL2aAox5PO9a0DNxpKN
wTHk61VJOqItP0rfrb2sxMVFzgIUoVNipYnd24zfo09y5B1GOfxBUKtWrZqyqq9zj1FldZ1ATDkg
XCF5KL7Qbt8F3hG9mzJdZY93oo2EBMsuI0aBW4xkLzDwzC6QahNX31RKTz1Oh8Ns5x5oEbTwlITC
FGxNykneoJb8UokQDNBnRiXkLt9x8sgF5uP8D4CIdKhmpRfwEMLLA8IxPycXKTHcOGXfQ8oZsBWK
nj5FNl4XZAnGWOE0dLL0Og/FgMxGCKeRCHtm3xSpMK75+0dUj3iLcN00Ub4lU87dSL+OKbAeHEzD
ENp3FgVS0yPKlL0S6AXIGG6E7azCbxcbsMklfmvcSs5AsaESXS+R3zbL7R8Gsn8yNrMOJc5kY+wr
z72YCX6wX5JeqzRuvhOzzmep6EH4Oi7ndVGF6pTmnANAbHzVJzozCqNxiXEgumZo8myQeec79y73
jVr6/wp1LfnR5nlp30G1iCersoOSEIZZFf5Xm3Tr7KQLllZRcDdo709C4bvxV8CJonph+/CRkNam
b3bz3yFyWomAm0hXBsuvzi+vz3IIwwcz4xrF7mIQ66tkTlOVFey/JKYs8eEpIpQvtqc7z6kt5Dma
AdOo+8z+rZQ5zHKcNJ18RuaZqvZZpSS3s6kEax2OSeqgHgBxVzz1ga86msV67v/6cbbrRLsy2dnZ
ok4RMsmUZInPRxP5nVMjuhjooQoyjw6vpwUl/IAsphpPTuUBhjBTRunVC3+SQu/39KCnYhh2T0m+
nz/wu/zVzIBNE5JNMNf72iTu8B7ualT0kRAo4Uq4rhAI16rkxIjGJsgTgEfiEj5nuqx2vZnjffBV
f0AleMf3e4dwaE8qMV4nAI4H/1KrZ9SQKq5xI3K5zwSSa6r6c/u673h0oMofi4FLaAV8PU/FRg5Q
pcQ7VEi8LdcYPjGCE7CPGYKds+ZdN1UIUd4GD8tLQJEAtL/3dlXtxCnSEVX4wNiM82/8rsrOulVl
J1scQ0JfxtXX5Tiirb3v63XCrO7Dt6Dx3kF+0IBBiUqN+cQHtmxZ1cnitBo3xM9CGXlWA3C2WMK6
CnujyFWxvDZtHvYoyiqTaLiGASHsiwaNdtmgZdd8i/aV9pFEqE5FRSZeMzJox3rz1Mh9f5gRhdJ5
4snkHMPDbSSoGlMVEEwwSDmRAPooGTEDSiHwpRlcE+rJdg3PqHfLAFNLxPMP3sry5aUREyiYHb9r
Zfu0Ds47AlRTmawOjIuYQ5Tr41dVrpftb6AokA98P8dX6orYprtkxmRO3Raa+qsl6OZ1eg8UgRSH
AFtH0Z1g2pE7DEC5Zu8cdf0vIEagHJldHJj+g3k5ABsstDBOFeYsI9FvOBYByN0sxCtIiOy/YvMM
C5Hk+HQKIWFmOF9WnBNDwSSRQxKd6Y00KU3bz7ogem3/cz1GCZ2MR3sLLJtIDVAdo7+ndEjB2+Gv
/8beSQGdhZoQ822tZMSSrf9eZ2LcmFXesFAM8g5z6TQ1wxQbHcknZcF2c0ITqLAoJGJe0kGzbR1J
Pzu0cuwFgHH9Ozh1WfhZr/RiFrAHL/KgtIN/WjJUhz0WsInl3/YZ+X/0FftuPkaGVEnaWgiCZ5G7
fTmUS2uqq1ZcawG2Znvj0W73sU/59W8d7weDJaFo1QHzHR2tLgR7SunnOeAs8pigFdenDY00FwuY
Oq0HDc4gGQRg9Uwmx6BV07eluRMbFzpfElOBh4z55bW1FBU/e7iQ0GF8j5kJcMO4RP6gCjrDhKlP
qRliqrIgvpj6Wg6pFlmVc95wtvRVr6VWl0qoW2v8uJy13P7GsGRRz+RB2cnRV6wewpPKdlMnK283
9/kHvB/LyVJixyqtMYbLV8GEKdfMJyMCwwEsW4t9+lkj/awFIDY5zgC/iuGgXoJ0AS29Jd/8EFHf
xj5gXr0AI4JFuRV1nZzC9mgtJxcrZWj03wGVlns+VgX6EWhJt8L+TYZG/LvS5HYNCsdE49fhYqb/
76YGXSc16PBCYRLT2zQ3k4hoAv6qX8UY/qk6EMEp4Oh7rRDMRgEPgK805gde6W4ky6rVoW7QVbkb
zDykWrq6TgnHjb0fTW/r2Zu1ppLDQVJdwK/Vr8jsSfOlNGOvd8Ds/yafC7V4JuyQuDk0Zp22pnO2
55z3gidA9ITpzl8fKHWPXMwPXSMBkcUrGIj/HP7gOBV7DooONCacd4Wc0fm3JyWfMInjbsRxRjmH
NPxJImiTo+o/BxBnJdufVwgCPV6a8J0vM5sE3XUvDxev8EMJohp0axAFhOmxoOyuUogbXn9E8bHo
dFBvoH5IDulHNjWu0UbrLghGvXQ72yroURcvBfn7rtQ+jEJTgNaY/rczQ8A+eG/nTRaxYJaZhVp3
tgGTf+cWBYMMSeS9hGbB/q4YmLXZi1+8e/6We+x7252602RwVzbzVUELUz6PqK/rAf7itOcF7BXS
TukOur8PmiH6x3XntpDad5XPkavkf8FURPUwKhiOg55R5yH0MMH81rPxllkjCUQGD6MZnsaNnyCS
LScOaub1oDgysuAU0/RduIbJtxncU9Xc72WbTgfBHNtGewOmJkVNjDgusqejpODXsnxQyaLCsqzp
Xm1pOmYY3wj0Uk3JbTahaywJVXyE5FGGtSw3k4KlUepuyjq/lIhO2kpOiKqgN0V63XWxfHGkXMnJ
gLRi7EzC5yziReJQDGAkroM+9fpm4N0Yyo8yC5PbXU/clmuvPwG4ZYd1pKU/f1Ab7RnENA7jd/4H
wsp3LQR26gTandSoQgcCmZIIp2+kDMy11Mcw8zcry2GxK8IyWh/NOUcaaivBm4Jwe/1HyXkdPf1z
ujX2h6IM2ayzpHzjzUYOU3wzkZiCGzK99NZ5v9OxnvLNKb6X+Yg+oxwEIEu0P2a84xJS6Btdsc/K
noIRTL+E/6vfwvnRxzB/jQEg/HsQnawYtvcYpDuHqoZYsqVgMaIlZowOTbItgTVfnyqQIRzk2+tL
MUWe2naLAM+Aec6o7q2u3R6db8ZWZzmu3yQgefYbxIHf7O4Jff+YG7QrqvrXWySoEBvQ1DE5DNeD
XLZZUQpTToK8tpYJmKpJPLvGQa2UwUuzJr4vFXslDCQ99yu7Hqz8YZZYfftMeDvsys0j91jvnMA7
Er7r7FiQw01zu7+rW6E0QF15EoNwMsGulVI3KviCAWkyfcvrt/kWxFSx7XEiWPOWf5CY/8qhOOfF
UdjCsWn7oqZUNWBL0IY5oW2nG98J3AI6tZoWFcUQaw1Vn5cSP3jyN/NGaBZJ/4vqmSVNsfVfu+DC
DUKqbgoeDMwfuwR47Et77iXGZrwmigIusD7Et+rPW1MuCIW+tJygb0pw1l8JMxWa7Yqp4qVO6Fd0
6mzApiPQJYxj2g8CDywJBJ8iO/5ki15/aM8POa3tZA6NMY2Bk1zVYMYPw+GZIufLT3GNEveHityE
k91KAddaIwbvZ0aPlO7Ey7nyn9EjXW9N9owzxdOGPfgXbhtKArS6QPAepwdB2USVDTnHohrnDvfg
hTPx8aKkDdguU+4s/zqksg6NOgV1OVzKJSwExHNrTF/V58YxTbxnPmT+/KDYxTzO3DtJk5BzYWeu
4xtPFLRBxDHMdueSQIcdZ02wcF3Mu7Pz09sDWXvdkzOp/FtODXUdy9vv7rcopEUY59EQPbTVbVmm
Aj5Y8Ui6SupCbLC0sYHlB8WdIy2Yu2rDn6s0tzI2VRLOwXt1GtWFVhL2AvGZJ63RQJDwl1M1sAkl
r2gqvqIknOLcyJLvcLXNhrcysjBO0lKJ53YM/nwjBh1NQ844/CsC8AY/VOIbzFFVUETtSbAdtozJ
eZB/U1ZO2Eh0oJGOKBxb8iL0Kp0u+qd3esbb+FfuZ0W0xGXpBewtF8PXpmuBl1AECoCvmlx4iIN9
nJf0PnnRlMJdGNHR3k5loRLqYIgFejh/faEhUByG2Zjvjvfame3peVR3y4tB5C+YD4UgfdRbwzIV
AB9TTTX30P6bxZ+LZa/KVRq3aqeXd5p4c5y1+mwHuToFHDJGd8TCTQx93OACeT0Wz91wZaDoWzdb
2GHCIuaeOw24PlgRQ6KxnR1jMW/J+30icwGbc4EP2Zd+DXc8gA0pf1ZOc8sL8I8JuV6vIcuyTCQi
RkT0azTppfOn1JCbgqdpGoEUy68nx4QiuUR8m3ksoFqL8gih+bNPJXhHlKCAzqJ16p8Bw4sHzRyi
EQdmms+jhiLO/T13E4xnfcdMbvrh63Bd3aX3VuFVOkITcKNqbLeXZ3ODYWfTii4G+nv7F6AS08AL
sAlCasHil2rM6i3Z/aZwDXZSLF+/leMB5XXnvfR/yTEmcvp1lxfIYSDrFhxP4M1AWmYlu/yxlPCC
1Ok/z733ysZcxnKmfO/Vo5wLS8xVFmB+yF8TIfm7OzxOblByhwHGA2BpBKI4n+ktt1AyZneI/wsg
oLl0M3zRpCFCRaUes5mPFVUGOIb7Guw7R9+nzywj2zim1BpZXylMbxK89eEhJYZ8aLWoWh8g8tjp
Qn0nfCzLVaaATeYykssm+hPxJloRj/I8Vbv4rjD5h4nbN47sxuQsbfl7isOWswy6g/Ixw73kIsVA
QBgBFdzdQbvgguNkEQGS+HBFamauZofAsLJiJNJUSLvKS4j415qkjtlZiWJHlb9SFpkHBDcmGdzn
OZqdD978kNwiMSdlljNQoNw/K7fHYdWu+JJyHa7D0FELCutuFsUK4Fv6Qkk+Wn7ObK2XYn7dnXw6
RWTpUT0mWBRwwtRIolDBeNh5GjOs4Y6/xESe+mB1es64RVYOyvOREs1XrjKX82domrlmmv4RYTR+
HvfahEHwPtfzGg5xS7mgwsgDOyv8YZeC2u05QxBMxvOJpkiNFxC+uRN1hHEkGRxmEjtSs31Ee3s0
ChOL0qDNWDFueZ7aNu8hvEoRa8u1f/ZfBFJ07nFmQISORsmVz17WxNEq543VluelnX+OPEqKVJek
1maLb/aXLBo6MQifVOoWgj/17/BmjaK5WlW4kL9oW+k/QfeDzPZRXWiM6Dor5VV/G8P8h3x5O2Mz
BoDmFpmzMDY4MkXw6bkM8NfzoA1xSV7BcZKWTy1hJd6f6A4s1g4FKYfRWmOB6oTMJNPEmONFEzf+
MmQl0yZSB5yeVTxQVtQvUN1o8i1I4s3dm7eCn+9UYmwZsmKf0883hrCXvcZDIseusYxXVjbUdJZ9
UOn4IdtRUzgqH7bY4SXKlw4nwzwwWZDN4giy1pMWTdES15+tI69Io0ckpXfW1r2zWF1DJG9j93co
SbkPcvYMhpgMrXElJTPpES91OBvizKmbWGJp2B8CR02RiBuY6p3pKie0Jzjtoy8uC/ej4NkaZ5Gm
XJ0m5vU+KdC5m82xcJpFT7Cg6AxdFuXCY98+cHoSRBzLh7rSCBLncqRJpBlWDkyqaInJl5vvmLGM
zGxB2ZdLoDWxz+hkZ+3l0jTDBvi6hpbc4RuSifL7YT9qOne02exvgB9JPv1stqrvwE3aLcqv4su1
Jn3zUCP3TqLXMCP/mq0Y18Xf/Fztf9uwzVB+8Sf5IvBnoc0Xg5KeIny+jVP51+WWtEedUI4gdPjF
xt06C+OHhbJVDgh3geZk4KurwDCmzDjbssg8ifho9tgyjnZMHUW7qCjdyY9kA2Q4iX3siHUnbz+r
VwQWsre+/pSE/kawEnSkv3mM62XMdukyTWCmZlcZy+34U67G1HLcQr3ItsEmUkfJeMSjj+Jb6Q2z
DAWkhben7XQLJpjcvx5Ay7IkH1dUXL+aaWpYhgqyYB7GTeR94LJo2ONIDyoPG8X9/6jzi4s3PrLT
YQtnDzk2cECD/Cz15YNqZn39QlqhqAsA3zMO7O4lDEq5MKziJ2WJpsEM1jaysQQXTMNX2LR7hU9T
HjhZRIIhcTR0nDoPL+XhgjXMK0/DK+3Ke/Am0ne3PJnuHqGqZcs+lnx4Jtn69S81VZhoDQ4rIVw+
R4fHXbMhVyXjkNqtNP2D/uu1WgHSjykyJbH25hGc3XCD8NbMSbije1Cs3EkcLZVi4kTxL7XV6wAF
bwVcE/pwe5LsrkSVrmj9gAlUTW44XIS+k9sJTuaZVeDOOZBavVR3m1syPC6+y0FiRGgt1/4Cx+cL
H/RHPqS8zOyrkxf5J91p5nl+JveY1Cd49MOUQHHahkbMYH8CHKzbXnXfjfPcq3fpRmZG7PTu3Or1
jY7+ue9qUSqayS/ont3ICkXrWJ2M9zJm9REZYdquLdmuwv6yTT65kwL86cwwW5mRVOpeviz36nHo
tLPqRRdP1IT1PBZHe1aUTDmcAIB3HB5poT+0O+DWMukwyDE7JK1XsBCT1Qdw5qJU5EdnHXK+poHO
FCfKR73twj8oVDlejf2FFmxGKJIfsyuQy0xVHtjcm50FkGv0yio1rNw+77doOlu7efriO6M4e633
ge/vrL7CNQaC/AekOI/xLmjXWtu2BPwQKyXZOkZSG4HTOn/o9mDpUlI8X66c2+LrU6yc7rKMllFR
6JwBpK1UfEMzaUSlTJdTe7tHUJo4W2gEhDHa7Yyp8bTKNzl0SMlanRqTaRexCZX+L1SE2NRwI0+i
LcsGj1m+7ibZWeQXVnXQoEg9YVX+xPC/MM0DWtVUjAQh2/M6Bvm6YpriAefL2zkNDZ7JLjCXVGDi
dQtkOTHJIU2/tyIzsftuXVUNhNpXCQuSef1U4Q7PbUdqwRFGxDC4Z2fpV2zxAZLq7Qgkok+QNQYb
Phjdl1aKV9JiubK90WTMAJkwfwIEL/++dv0pf4b4WFLXfyGr0AaMty5XKnZQNChD9EPFqvbKWkRO
3DvKubz4TDKx4XR7rWTahsQZCz7mZn2FiAGLI9KE2fBoUzW49QaHyCb8FhHu/vA283mwmLLxPsH0
vY71s3MkRw3n/xRH3rW+O8nbo9fUm2Ukl78mJEWXJvKpKDF1U34ucqkyKf4jA7E6LZJyTSwRcDir
oKKDzFf/ZMPOhAOVXsI1KXi5bm3WO+P/Nr/4sgpwkcMWzTGrOKxj9qvPPZg+ksH06gaC7s2cRqWz
eL7nrRBJKJBMpcCERkLXi0WuAAUS2g/niRTMnCNxxAuWHdTjA4dzzQK1wosnd7ODdP/3SFa/HAOA
vdy+qvNDHZWj815ARvKCaSatRjHZFJkN3sHPf6vI6Cy2yB02C4MrGk6IO8gqV4unXT6fxQzOzonE
siyAJsPHXnvOEKFWpmFVt7KmBPHgBNWgLjm438uXQAS42qDI5LbhFjmoP3U6J56HCwFSdatFsccF
t/gPEUOIbyvjhuzFSCIqtFT7eYa4EtuK8HwKNst41EoEoWJCYttYxhF6SJfyvbsqRlmI7lPbrQud
xSPVfpjOt4Y4IMHDAGc8eYxOI/S/QqDVdKqW30aZSNNMaFRmgHeJpPYb2TYXdny1bo0CT17cXJea
z+Z9AGt00Zdu9+23oqZsj48FX6edkuEuSrMIEiw1edFxpWOHbMIfpIRlGI1k5R6//YgaHfZkWFch
nVub/HR1HSYyErqXkGIoxIB7Zw4PqKU+xJ95KPsrsrKg9ZGPV0pfcMH8AYJddmnNSYIwYEiMQP//
aBGzP0Ls/080C07jx9IskZN9qLk+Bj/6+aI+f5qGGLFdVFHCULv6ponLJH9yTqoxTUV3sACa3Oeh
ksW/BD6ldmp5RT/CBE/RHMpCcAzxtX5y+j+zVaUC27VcsH63ZrXLvKed21LG2NcNFyL/VI9FViIy
3wI8ACMTpkCTwHAVBavn9jJeZKQ7tdd9QEfU+BSPLyw/7ou4FQTSUKrY7X939/AeiGDGf3deN8oH
rFhd+Y7hSSN5ra7/BPt0IK0cqgkbxmoq4gpEKfGmpnHm0CM2KrqdeoAonRL9/5zYt7t8bBEqxJPn
tmcZanJUYQli7IqJInXWSYBiA2P8aXpE5eRHxJfjPP5ZPI5KzTO3H/A5em+Uzs3SYxDE137tWXkW
iYmmyYXV/Uucofls37QB7J6+uPtunCh/oMVnCHw6otRt7RKsa4b6pD8dL90+mk5p8U4gwtADhFgJ
jpkIj7sgD/3bt08dQkI6mUFZ/HTj9MhObk7BWf5qwBBTpZyIE2KW9eaKs4JEUCcaChjzjUpbpj9Z
7d/FeBMX+RVHTGdMtQfCN2T/bh0/0rF2uVAaU5KOiqVoU4uxsKTP5ulK1i6dZ4YVfwb6514ow5Md
NoC0TqSQT60vhYVrnOQLuYw5ISn3l4N6WPhmGaGxpJnEsiGeZDaLqgIV1Iphp4IUDCMdfhY9or3x
FJg94R/WLkOcWsXXo/oKYh1QzVI51fIz5A1NqHkJ18/e7lgKnXtdRqfnDWSz6VMUm81CxWegWdUj
KAJaASycLpQXI8W7hMosarYXvGsSywHqSu04ffGRtn50SrT04QjFlGtGt003PZzrfoLy3Sf73iFx
dho8HM/A3FPb/vMXl3Qp8oAzAwxX45cURbjrMDfa7L+2SqMxtC3Dcxhs46yDXD7zkY47+IYd/EAM
JDNvua9iVA3WAMvdN16oJK8f+aj2ffNSMiiB1frS3ey/OCCgT2a8DKYoM3BHIB8MsXvhGHp8mlVC
dk2Tgv8uuc0FiouHgMoMzXmioA4wDT/Ym/lhOMlKvCeH/ybLMxpLMmTWrYRtExo7bzKq5odKjFEV
vjsuuY4iOsMWtsEUNLhGCdj6pDX++JejmRW/w5cYpAdKFwZln+1jsBNOuAa1lFYvEmC9swCZ2/ST
OFZ3d92cgSAc2PhyEAPFZTiRWGesHNzxt9cDo/pEVWsxC1mMB3HerxmNGcXEw208MqQ07glp3sO3
QerWTw8s5Vgi5/Dd9G0ENFj5boK9P6ofYETHbjYjN2iA8zTi5Tuj/6yzVWemrkkrgQFCbpDWztmq
d+trn+jmTICgDQHehL7jReTjt75km1vXbqzT1pk8vEpbTSkNb1IEJ5T9UIe9CN3xAMkMkwWG5ZtD
HDDqGSmoE1F9CeFA1Ru746enyFAwor4lt3gFvCG2ul7Yr47UtoZ83+q7MIAqhg+Rljtl7+OF6nVk
UV5eg6k1a8/UnNLLmjAohqgOeZV+pW4zmztJLCV0hv/yfFIMSQICEIs+kBO07mGfBBTSnq8R7FDj
ziCa1CPHPbDvob25uZJdHuv70FrcFiUyPMetmZ+rVUKK4WUWd8tyI666t2QvudEms2ljGbq2sKbH
sl5/Vy0Z88BMPopf36MSHmK0ogIj+h8goAXOIM6g4EnreRQ8ZhhGIXMuYGU3bI3GXNCBFAKsOzOf
vs4kIBvxLjIqoO1Tq27EXc3iALJaM0QUP8O5sge9s2uiktqgstiuY7DEtFSfGfqd9sJbtMrAeXCs
Zl+q6hDgVUBBni16hYUvDgpAOpsTVgKxmUpJKLlpVsYVD961mttkNXqq/KltkcclPXdU226aX6NH
rhb/0aMKLc7u6ZlfCznS5goQR3c9alqkjMuWZSGhutUdbRB0wZBYCQXZc2E+1RdXnBHRkbrmh74N
Fbq4u9FkEwLihR9xfbrLVJl/1WCFIX+yucVHOGiQRSV11XkVveIjF10MRZQnQoFvFAtB9vWoruwJ
OQ2rRnPJ2eTcmGL/lUUU/tsyoiLnruKI7YONjV4EbCl125kieqk7ehQXlIEITCO0s9zIqyI1OKjE
BManKoB/CTUg045BNGT/xXqWlrJIH3dtY3EZscQjf/W2p1xc4huMw3OxMX9ndgbr+56rpvrTpnYp
Gxi/cJNcAeyHp5kI0YdVBfhaIWPC2oRdsxDJG5CY7rSVmgP5zbs5TOn6ovIC0nf8ypH8zpwmpiHR
+QFo4b1Q+YOQBQMsGbaiMd/1N6y8GzsfXDWmKtwanLmRfiPli1C/TUDf71R/vNe9x4Pva3EOaVbs
VdGObezvJ6IEwxMihgUwbh8ue4Ekaiz7RJ4mkJSWLjEoMjSBuQLOnwjyGFdO4yGddJI91/KzV8Nn
IN60Ne9coGoOpUmn3ztR/Fq45Z8iRHq/vyvuFezND52WLrCt3jjjdKag4TQ/ub2PtvO4HczqJxEv
TRRJDH71CYupUcJltSSXTxRdotTZO/YdsOlJTPMrvl9l6ffqXKEk7awS65cI/1FqOJseaJNlr1QP
Y/dwFS4A8RYyO/F2iUFRGDcQe65YByA6rXV/b40NRqdYs5vngndYRIMRt8jawEF07xa6p49WXx5V
YyS4J4KFF6Sd6WHJoVWkdlugZoQTt1ZnJJrg/s2nuV/QowVPTOHLkXY90EMPgx5SN5YDU7hy2RCM
pTV7d/iC8/HIq735TuxkMQfm/ejRw9SKf6QogFIsKhnY3wPBXn4+DQkWv6ggAPQsioOXHsbY738f
cczBvyfFg1pT5oCn2PX99J5NC8WWSv480tvaEev9H1DAYACAgxUOPCWsBEu+/QsFN5UQ48UFK1mV
hMJoZzBul26ktESHI4GqjKtnlTGgUMmZb1rNBbdhonESODZGk8D7gaYmDD9+/OdxbK5wWdiM8h2K
jarWISAAoi9EuFdacTITRlR5/+MvGvEEunX73wx0NjRvY4QY2OXt31sFGPFz5VmqlhJ+G3RIkOH/
3NMEB2ls6RIY5QROup/8CgyHZyqYP0GKoEK6n2s0N5yQ+Yg5R8aiTuUW4crJnKVhqO9EDFzjiD/O
yFRPsSRK9ZopIZKC9NFYsjehZlXCElSHoPXfNc+i0/wzYGMDL5jy6/OYyYBR8XZtl6nMsElUhf6w
jPVbHEog7JqGJnPnA8V6f+e+etnZJkui9RFBeQgCREI0LPfgg8Cs30/Zf/oe80j7gYQttmx28++r
qMPkAoJqmsz1mXS55ExjxVHi07zid4XJk4v9mrRyYiCgkhnDU98PoNNhDSyz2WS1OUPBTQPm3EQW
NX9vO6m6oFhS2qLxIsQFS+lQpJbNhdjqiKhXqAt5b53mYwjn6kkTnW2RwofNH3+RXVA15FLv2wPd
2cSdnLXk+TBSRypY6ZPWq3LhAszJXCrtmNIcU/pBvlX3wFEP6bVe8U/7yK8Atm+kr5ljkRcU3qFQ
g16iYZG3/pmDY5zar/lucqGFUfSb5MIGzWRIpVINorOZGWUGE//ZvXuk/ACmKEeNYYh5BHcOrLmk
UkW8/DaYiN8QE66WRfbMWejOqF1IZ3LWww3lxIh6RCKZzfZ2wKEhwP5Je7xx2k7Iz3am0sGeXDjh
VjF9Fsgq4Zuj4+tMZX7aRcWRFo9OEccbV3LqX2HOAqtVfHZawEioT2ZGzttTBMXC42cuQyNKqOOc
fIQDqhTbcb6KnDtkGufZS9S+CgaR2i+SOqQO7NCfW7rAvcaqAA2jOmXuK7JBoJvDTTly+tkhwOQS
frnXv5gHaqbnRQptlGQIQEZqz/vdMFF67OmnG+O0Dy/cvpraDPevMm1xJn2ybqIm/IrcQDyYm4fx
tlXTWcMKYW+D+oolLInQsBOmmmXGgKcQ21tsPHy59juCzjwJxHlEZ2PJVOp72o9lIYCcNndqTzaG
lIUEqzn8cqvDzeNH/I8uZqXOY+0wGGM1zIO6k7sN+b1mYEp5NowmzUWSWgp3HX426C0K2+GCRs60
5wiq5pBDEPfVB8udQbHCW6rxg82tZ2y+ajs6sY25pjX1PQs+A1vPiLklZh9EAsdG4ObnMVyhyllF
tbEamBKKMSk3z2zuZSnKsOhifbuIfz5rZZSsSTz08TPuKKx2s0WA79aXJd2Crl9v2ipFvqx+intv
p274vZ5hSJYctFxTDw3UzMs+ULI373Q0z0yo/e768036ThRMQDZplPPMi4eqh59zWMXXkDKmfKI7
5VtxeRmXEV930gOQN1Wt85qqYFQGVqjH8DP+iSZajT5R24poc+jNPPFq1xMDawZ6SS8Wf1PpRQyk
kRi2M2cyOGd4V9x/kE4+8GLfeA4nY97BOT3FipXsVPCTlF6PsUAjF0HnhoNekp8XnE15xsvBfVH/
0UfMsBHTFzejt59RNfCQQ4Y9psphncRnvuUBfQl63fdiZ0hLdnLSpbHnBTsLhUtfd2G3QsTju3pv
c7zIRPkC5ajrymytiow9Cv8Zxgit8erqfaKhglUzeHW+2tXmEWh8jywNNiL2yvfd7ecIIXynsIEh
LRtVYZuWKJxZy1t9KPYtuDr+CZ/xol8iUnWw/bBI3tL/Wsd/PjMMlwIEBO5Gk/HHacYXunNPNxbP
1F0+1w+DgOXxlhwKFYjXqMvAK51dm0qFAgKuwRVZHS1wQFb/DhQ4seyTsEzbobqq0e+cRnrdnned
agUGIKl/hghzgBRffO/2iT3eSBNiDtt6rvNjtwgo/85rcQfP9LHe0oP0eynR3cPmki2Ovys39+TD
kYB6MGfiAgN5Kj7PATFPhQD2n/3T1RpBJCjFYmKw6BnDk1Y0VDjJ24/dLf8QTRcgHXUdS/xz/46a
o/OTw1t7addWT15p0kqf3D2oyloFTvl91ts2O2bN6BTmZJR5OyLYGGIWtfkgkYJQssNHTVC5w4L6
m0SDgGfDq7DeH/b5QRM05YG6e8SC+qMSIiCNdPghgxSgRX4hUu7/pN7P5wQHrCDV+D3z35Z7ydE0
pCIEduxlzwU/PA2YZlvopz2EeERaUdckdFe6JYUgPwhJRi3eiAmlnSGzoGqiwu9oo9w3Eg1ebu4Q
Xh2eDBRigaMU92x8c9nP5C8/KQDaNnIwCofa2cFODaKvWzj4e+wqZNRP8OZS4mdCQfsFZqkNK4oo
xOLC4bDeJEN5aHH1wf5elxtfHuiBAh/Zl7gVHQan9rFgc4p1j5MCjYU/fkalTJxwYWcd9cQf8Z43
FbCXCJ0TKcw46z13WzX8FEAbpboIGZXCckUNcgFebzI6HJk3iLFQuyQRcT9xj8qXvJyiVkVM49ik
WRJRqiQxc1dkQbHKyv9l2YvuEvNc973j8o2RT0UcT7+ReBH8zaNzjd6bf8KzZ6g6Faa6YGpRvmdy
TCcm8+RXPbGwra7tMNQ9HZrFv3GmuoPDUmsSUDieJ0nWo323YMDIXv55fQ8D0UlX2UmFLeS4mpI1
1+PuWi+TyV4711cJ2vp1ayPzcwtuq8jj6hBkpdnecOun/8un5rnIivJ1HR9Qv83EoV8qDsV/t7Ci
NMCclYSt54B77aGl4WJeKgFHUM9EbUhIWYzMvWnRG3TuMRK7eshqM/aBylRSEcp0FdmxZuicQkuU
Y4Cp/6lEkCr0fcZ/kRIRnpoeTaWcGp/uUgmEKhM3wkgu8q5mW9qrlY6ektYG6FAfftosr1TZK9Au
OeDTYcjB7ruBVLFR90nFl6SWSAv9j1MzQfQwZyk9KE+9q4Ighk1tGkWV/ARzw+YQYCU/DNKjmZsc
9MrpQD+q/nqGdsW3pILv/cP4AFZvhkpwSKxAPaE3QinXisxUHLujz70tTqpSaxWXihpHUPuuXe9g
hcxeLRlJF4w9hOoCMFjQ1yH1NvojjMjDKdFf+2kii9w+1+xAi6aW1WwxQAp4/4oxDNsUr6S85xV3
HcuVDyT3OtHH3tV7LRmoZ4U+Mv3/wYr+WIpKH+HQtgeTy7IhYgSLrcqEbnb8huqHvdB+YpEd1Tmz
Sr+JtMyo/oyMm9IvBaNxid8yD4P4zLbsD1ipCnI2Y+tJaAgO/eWAuQpfF3jBy2PBVPndV4vAjBZD
L0rGMS7gqZkvNduigO9iLNrLdZcVszFNMK/My+7+OhYiN0HLddg1JkZtmZOyc1EQCFLHINqnJQ0D
8iLXfijJa6NmQgDwPAKcMZAzxYSO2UoHogyJXWd9/gZV6W8fr8E4SHHbced9tLlEgynx3GPwK9wg
MsC5CMXr73bSEK0SOa0CO4RTub+60k2AGFSSu2ZudtM93+MOD1LvYYXH0y3M7y1CpykOpDa0f8T9
UGdE6c3n7GrQjiO+mEfunh98/rx/VbqBDFgIA7uoZdWzJBjj3+tD21P/WO3hX/zESrkQkEDAwF79
C4813/OOzZZ2xrkfQZoVUb4y9XGTdHQdFLpAdcn+NHHVT6eYRDpH+g9zMzFjQmcyz9qnqdc9kk+q
a9No6IumB8FKL1KK+rQkG83aIjA1FtoF3aH/jnkgsRi+TvICAlhPtJiAMF7+X9Z9EFp6d53rI2fg
zo1Qwxwqv5wkNNnPmdabEQnP+Js/VYp4zACqTNL7OJaSPQHw9wwOCt9ba8QIzlEt2As7tnaibaQa
erRwx2bvSzZF1i7UvfEasW36BxOxQMFpdR4QPBTzWnv9fqlbdI3ANZurophJ0QFipzDp8lcTSPeu
6NXaVw2XoYPL6VGtzpBR0oAgfJ5jToOrknqbRFzG4dZfB3tR8QGmEeHe2ph3ouG1A0rDqb5eSgfP
ZlXboEe+QyvJUR3n86TJ4zTs1okmG/n3In1v0OziZvncxBeQ48wZkAXLVEYBJ87mbS1Sjh0atriA
1i1x9kATSrEiieAXsmgYLi0S+st3NRQpRjKd1wtWq2OzBjXuh93ylRiZFr45dQrDmEUHNvUOx2IR
j6zX91j7Q+sP/f/siGN1K7gTZbfsMsR8Llli+3gw73FJhqZ+gT/qo5+OSB5UIpbwvsk9QsRUOuQy
sFmuqUSMnhS/F9EeN7Y/nMf6QnwN6ebeQf4/EcEXAXktYXCheKX9Gv6F0+1PKjFkv9hkSo/fucA2
RIbjz6f2m6a18qCICSbUQvX+jZY1v+NzuyyIxXYWB2/XY0j3mtmoReUCUU0zZCvZt8mUHa/VQeKw
0bNY/cKw+TjcjcijH23+QuVx4yXcqDxUYKghQaka2pDqvRPu/cOKtFjFHOzwp0P0LKleH5faNA9f
quR0wNdO9Y0ZkoCmuml+cbM088lRQQiGJ6+srguinnQ+uSGYy4mvWriCEOVzqFiQmZ8PZqxqQ3gj
rgFO/3AlW5aQ/zfKckIw/CODelQvpA2By20dAzzi9Qwc/FHseeggIpbSmu5VdvERy5DWcVWvyECJ
ge0pjCOcpAwCfVpWqw0r5sR6yA296n2nVwQ4oH4XjGcm+wlyXloKYMsL5UPseBa0w4/ZB6zqDC5x
yqkOL+5HZcL+U5gjSA57P7tv1hJOiLUrv0lGxVdDUOnR9xxUIwYkg96d0s1fZZFPUG0/SZ+BmNnv
1PX5A0VQ/pn/gmeNY1Hs2V0mQKmeaKPtk/Fo1H2MYmIHWY6JCvZKpKHPZK+HU117CeGb/E8xVepW
ZE4hiMxU84ko7RWhIcMEfJORdOtUzKRT+SaFCxW/b6QEU/3okmrXW5u/b3eQIrnwbtoJIMlE6gg/
M+p8HF2sGNGmM9fcZc4S8nJ2NcqZeETqyESNGgSSzifxxLpIuKDT5CDytBAnmG5H6Rt/7ejOLkL6
vRJqIMGLB5luOvpFSOVbevVphymDIVTIcC95bOMOveH9QoBFzBKlXlw0rH1xxrkjm9zvJkjklw5y
0HJpVTVfDZ+S3tL+Py/TJjWRHzqt4GCApo+8QaxUSRI0OHV8N2lvReWto2LXvuJpeSl87x4deezC
Z10Zh+xuhyQLm4QjDVwJdEPlyMefcyfobox9EFGz/2HXAnx/phkbVWM22npYOE0lTQqNrnDgEvUp
vQOlbVTsMJLOorypDYrJaW43E6CIIQM9AOO9ekf9upQatS9Pd2vE4BQoMxIFtJWlkJVLt0fhivX9
TLSKpJlhmoY+SrtxcI6NJQkRMkXS0PQ3B8BroDWwJv1tM0HnmAh9jieDBSKRTopDCc1c9I2asjXp
bbA6qeyKpLItgMAGM7r6vnbPw9V5zGPUfTi2u+pN5jDBVBp5e4x9Cg/scwH0KMw0tZpVOOzq4vSh
cXZ49/G19ADJpJdVGB7oNvi4o/AJBl0dmiUa0VttaXXCakcIX3B/vlgYVAvPX4h4qTmf3a9yNxs8
NTcgTDd5QmQEbAagchtH846U0x/VjT/EteF9I92HvO5wra65fb4Lhidm8dIUtigD3emCV0J57yrX
O+Ovn4FjGgFR+EvMYQRSxj4hQYZDTiHQVSnP05VmwmVvtUJvCCvt6eElbfPPW8pIp44kWwm3/H+P
0vZ02B5E2TbwfmWBVTdgEzK5KYYMq+/Emeu2Zc+YOo2NdwyC/rLCPjnBmlxjPCdSmFlwkgt2337j
NQ4921ePC1YfqumwMOlOaDu2DRv7GRC/k8z7sMt6VdfVhyFlLrFuCcxhcjDFZc1ouGQsJ+242icr
W4DIJRVlH8vXo5QMKRo4MTgnaRk1apEmSu08axnPyiLYYa38F6xvlpsp/cFj8FCZEsDd6JlAxwCz
V2fIMagqlsX9IL16+nVMdBMU6dnQwygAQT+sc1joOrtnuhL7jaNBjwADypUsZj1nZroMmZ8EZrI3
EhAHmV1aFtaWofrFActh37j79fLL8sPpb4AMBESftjeeYsEKbtO6qJ4z3MvbFmpW1zrtsaqQwh6T
rkvsvvoVk/nmfb2Iafoyx/FOKUcV/GJWFInaCEiHTi7XgSC9fS3R6zzSNLuUakI7/GsyOq99vGKs
WUOthrUqio8O1IcDjzPH8Rr/Wlq7Rt+XrI+SaTJdh80RUYz+EBieO6A6NSN5xtC7yJD6bkSuS8SL
Xw9QbSaIOgRPaS+F96vA6Wm20A2HbBjecb29OQGcBvJaPJBsBkS76Xl3IP4k2NUm4lXjZM22VOJG
eI1SvpBj6rwMTw/Iv+WY8pshaoTHsTROTOPfoNHUXmCAJIJho+9Uk4XsP/mI7dUD4cdtTm/8F1GZ
i9EfoVtpFGVRjjtItQejVBvatiWqgL8qssu4pIMc4VRwR+4dTuXB4F/VsDsoCLwJSO5dww9m1TBS
Iie0kmwygqP88IK+WmRL1T6e4QV090j6Yx+RcAxf49pIVreE54rp35kGwQptIXCpkopjC1OYO/je
DRY/bNSXnT4HAwAURz6QdWMmOFuoVmC+gkxt6Qow9prrmULGw9v+ZirmG2EIAwTAIqt3hny0vroi
IIUy6P8hdza5JQV5Xz/41T+tsvl7SPpMZpr3c9NfkVzxYtuT04/uZaHGwHyKsPM8IDNExq47GEEF
uXNP8PUsFeqmLnjlBtMz0keBaR2aJ7978i6qTt8I3L6api+aD+Rb9HMZZb2nvjvWJHLu93xcBuDM
cLg9GB/ZDBjy8dPuRiu9lyv1ybt6Ujz9NarX/W7VNWKGzTDtUhEtTBPveBYInTXBAqV05TX3+Mg4
7bHg2XFxZgsg1j/pImQlE5HpU8E1CP4LowMZL5KmXmvbAJDrfo/MTGp5qOAF2sIFu6PpRxzZ5Qii
4oMrcTcdmBnJoeaLu69ZTzobDNbz3mlecUtar1crM01au6nbo5KLSfBZ2aKNpSm5YqN7/Nn0ZHaZ
1j0vYnB3ZG5fN8tyfCE2NWef3817K1UOSMgJkQ4XuxuzmSYB+2h5k4e7NHgJzRhV7WkucHROtr3g
QTdjXFufIES3ddanh+Hqqf6tZxnOFx6QCKOV96OCWicRgyM1s48yY17pgT3oviRXjtbV9oAngXZT
dJyY36drvddm/5Z27i9+vHGAfM16B742O/VkQ7gcSruMSLcTrteF/kGUgP2U1trlgKRWvvwk+sZL
mBTlJpzvfQ6Dp6lPD3cxgwpBbfn/howdbIKtRYKqpbbNDeJ92nr+fY6DcE5PKIfL8X2jgXa8aO7S
WcgtNcD+0j5yghOIx3JtWIVwmO5YE52/J0LSplkWHWb5kIIjfb544i0Oi/xYR1iGAQcjs6adTTl9
jJhFpy16Bywx9GwyHgAUrxNcQkOivSU/1x44m5Mb13dZlMXu3PgCyGw7s/kbUy5V9T9NeCeVe1OZ
VtO9ey05WdYOKRpYnoV3M8/cfPPassOTLKY6rtVfRPDXAH+22VwTFsOuGoa+NtInNhZMOcV73zpW
zR4s6JxmwTeO4lBeAulVm5lxtgR0rPv4ExI3G4rOr8uhjCJQTC73b5M9hQEtXw6ZLNDpHBUqJNeo
5hzqpNCSAicmaK4pgMOYv3+ChojFuda3vRBtgZnMUl1Yza9qB6u/8AnwgDW1ZnZjn7KuKv3G/n6D
FlG+tW2rlAxJJ6j3U4PvQmvKEh8XkIUxWucJXTgYrwfHQDj69YT0yTu5huQ3KNimYsaSZPpn9nWf
odECCphT3Am/ETupn9uLKSzEDT2I0gpgJEya1JFnAuwNN3qGDlT//FZ6ToxZ5HirPuarbuv+ZJoK
KouI7pt9ePuBHua5FRGyZ8kXCeyL+GgcoNJwkGpW/7Je55gFTNLXgzXZrhwEudllDwYpbVY08Yod
8BwmQ+r3LuexnsecCNYIS6EsO0dcPq8x+buKheD/705ZTsT8aKzPqBoaEBZfvsreoAgNzo5EC0lX
ZBz2SCo6XfTi3IOmrpg5Kn8UKGH2SxZuIgCDJB+/L6SUGeZM7Teo5k/gqxYwMOhJeb5pProbLa3V
aYVvYWNR6v73icMbEEJFP3K6bTwl5uRpCnxJZ/WE9ewkNxVrmWPLfFoErPBW92VXarsEn2ebT/0h
uOL8ifYbhWhOuiislrktCCaV/Dw9hivjzTQmEfoc6HIFtXi2OZ+piQDUt4mZ8AUx7+fdszZdedhU
3j7wZhBxGm/VDW1W7mCG1lt4j8wAcgF2Jweg2OIG9HLEKgTHqlnAP/DD32+DiWwh4wcNBaJ6hVHV
y4iOqQBO915hFNO49jtqQBHSnBYbYdZT9vtrsXSUHAqNLUp5Gy3sAuSdPfA/b41N7MZPk+yfFkzT
N9YsG/8PunPESqI2OHitoDJ53LENuqI7qONb7DMSAirI8ylIG+XPCi2hlYh2tm7gsS1/7DxOYit8
Ctcl0fSNxHvKfZrqYog51r2qQokVuJrls7g6I0a7y7LGZVJpW4TdArxYeoBl5J9GBHXShNtSypHW
9+lYsJ426DE6GTTI8PWMcJz4UHc5T/E+V6TRDcIhpexAwaiTmqZOzpuV3Ayxp0qJJrtJf+Ee+cdn
46pD+rQA2aFAkpX5BofnZgjMU+lQQO5YlfvdYWx49XNV0SYYq3wPSXc5wfTybp7+iCcmoOTGm5Z7
BxyvAGC/bITk8GJ6SE7e7GtK63fuXgQ7H50HzrkSSSTJrBwYzn+INl0Wr223szFxn1UVS6m6K6dX
ptY799UHTrTTkbdGUI69Tqyh1ZUCHNoG9AHQ7sCJLjHiF9uNaArNZlGkCy2F8CH4d2OuPYtNkbWj
LTC4AHHkutqOyuDxe0FMdMSD4Wc4KLcsgSbsYs5//ynPaMORMs6+MwlzWjVP0O5Z19UW5DY1AbB4
GAz/VH+bumDgsEv0VmbsfHwN35aus4m00iopfp4+OixUEW7nA8iQKZ+Ncif7h57CbK5VvLoN1ULi
13oXUTdfUK0nYc+sXlmMJUTaN5ascvMg44NcX1Llfx8Gp4LaK3/d3nzJb5Y9gcmXsmB2aB8ZHjia
mpGc2mqVDOILEtW8NuDPisBjniGQOgdTXx5dtbrVCYM17zbwDG7Jk66Ja+Vx5ulJRW8RQv99i0NY
yet8Tn2j0GQ83ddUEPuw1LZ80ldQcbeFrdXBtJz2eim9DZtjrDz7SzjAAPy8lkMGDdIePzEYfli/
wRuWv5+dUm+m0LIRtUfnte11U1d43pqaLI4Rui3AKnxNArzqA5UOrWiFoL0TusBLfqHnEHWZEHXW
oJQf5yAVcy0/6koE+1kgm635lu5ssLcPHRdslMCAXfL37mjABhxoIGpNuLkqKG5lL1g1Y3U0o6fc
JFSBGJeEvGWUYs7JEc2hkgJoPMeeIUfsB0tXnKh4PSAgEtHHRFpUZI7HBgUjx5hE5RfyQd2dCI1C
Y7NETWTJZT8n6UG2jpGSS8ju76xNQ6Vy4VsDUqKzURwWlmOAPR+wTFm+sKeQQ1j51m7mKCecUliO
Tn+UaR6IeBuO3PGhdBPQ3lF5mlmGvrZLlKpY81SW0eVj1TjlfeYcm782qUUAqGXSkf+djUmfQOKm
EkdBey0zyJsO75d7Cta2TJptE27bU3ivw7iAjwDNgME9ydUqIL3SMUiz2zcjxE9nTsBEEf5EuDdV
UGvEvmvwKP9PH2VyCK3L0E2RmTiSbYSsnAWUVLUCfXSknCoOeTlbt+/36LIaye9fnnve0QQCbdCY
WFBaWHpVmZkSk3KaaFq4o1GPbrT/NKCbSuBGXq/qBFCA3rUrhnnYGccU7n+pgmRPRppBpjjV6mBq
5SqHRreXKfjttG5+kTI128QcaXSm/qY4iS2qOJJOxOTXCzuynrJTBP2boBHxHswVY8pLb8dK6qil
BfOL4AwznE3pe9OIoEuTeB+v8YPiJDNfwXlIOZGpY4obqWRR/5PqILR7Dbj/7nMxNhFSVxZL3Tq1
JmxCSCToa1pKUQMBWbgVxZdl08raa+r0pNftsVk8G78epkx2/u5DgpLbmuj/dG8wWivxd2j97icp
aeqxWdltQ0y0CbNfesDsBj5/EQAowGCqFWaEikpFpNTszOu8J6hIA3se984BYdSCu/8lWPF2g+xE
i2LyfGTARlgSmgj5MjWzkPjSCSs3fZlHKGQZHM/mbIsPEPEUGD0Vkdk0hN3BfMJW/6h+kMs8BNov
NvHW//MUBhTtpL57eWnFW0VdfMDNykI+BqM6Ua+FoWt1FE5K/PG2ibCMPGWLW1BMvv02WWVBa+Wm
SjNAT5FGLflVS/HMP2Ge1cBESTjMB4hYB3yvZaWhtPkhx4ISc4tPppEzDi8lUmJD30nbsZ38HVz/
Ch1yRK/2ypvKnQDv2ZNdxFZ9rCD8TpcuEiWq4N3ozxcQtoXXX8AYzlCcqtniMJOZ6QaOiYSgfCsI
ozJr1I9GcR7BDWBxnzqw8KMqLgyplBcWhws0Awpy9Z8puzBuQQkmb8Pbj8AElP8wP+vbQYehZZdz
MsMFg7neNCZbC3DGqZKmOpmUxtVSciRyNm59yIWdwx7tOeu5eS4N+ai4sm/pPR3G0R5J8AM8DkTQ
YqbiO8833jW2WLog5sntuwzVXE9C0KNlsVRNTcBqtsgTFyWg6ZMsS0ynthvYqiF/dmy9QJ6wAlwQ
UPcGUntnoEOpSyPU5Nz14qiY2wfwvcGORZrm8fNS5WfliZci45h42clpPdk+9oCS3qaphEmeiQel
8pYZ53xX60hIseCV2DP/NbD/MBDHv8g7q8QuVqwzlV/CNBG/mlfCSI0cudZrPKQv2L4WXb/iWwUw
npZ+rfyHqUfU3ATo0LmrBpOJ5qqT9NSFzh/JUYdj95fxPod88rwycbN9oD2thIpWPh9nii8Po23w
VMb6XTTWgEhaXfGBy5UVpm9IlW/MSo0nNZA8AKGNNliY9ZmGwRxko8RvbzElSheoDF56XN/D6xYc
bmB3xfnMZzZf1n/V23jBbuuwDvoD/N0gST5wo6aREr0mvPdACQZZyIMNtTYiLMrG1bCy86G7mDoS
36O8Eo36yYdAUSs6XtdIurrddc7dYrD/85rOXqgyD5WQ9DbNm29QFEvb+QlslyxqAim+1HTo8HtG
X23E0H7K3kVOazJ+txJh3Z9WLpt9snaEgyhWwnmWbI0yfRz9M4wOrRNiU8Nq7PSB2U/iwnZOTL7X
5dTWUWG/9QhTQvZQBMHGS9xgbb5p4/PDoZ9Hd2332anA4x8apg+xXj7H4pbs/CNtcUlG1QY5yLp8
WIMqeMHbuUfBRJ6BnLb0RKFmyV52qou71Wf5kGFFlz2qIqK0/H5eu8kWSoW8LtOSPYjx0GZVHDtg
O9UP1RnR2xgw4nSCmuIZx5rmJXuCBDPorBowLT2aCiWFuexDAtWzxNg82xqHfaxhNJVz6T/7feCP
ugBoMxvGv01g5PWrdHYb587tm4lQ4ROIPX0onkM6rk3VWkXv/5jz726A1Q4Eq4M46Kl6xwJmomBy
WGAAnDi4KTufx954kxq6uGjjJlRlI5fWHJsakCsitM70oUAuUYdL9o2riegKyDT1bFrcAdEH4eh5
RH0KvGJYfIa65HDLYkyDhlzfeMK34b2W0EfBE3/0fyNEoYr/X782ipxIFEZmMYo94OZ6IowDv0DT
AQDqkPtCzSGg/x9okwWBxdoRLGG03MXXN2xDNB1GTtAFb2TXfn8lb+GBND4n0esfVMWEvAHt6fsL
haCUmDa+ubLhqU9C6riDxLfE+Y1d1/YNbpJbB1seIqg080LJemAOU1syP9POjRlHQK3F7Wcu0OyZ
IpMYPRyLMCf2LYmVSMhZkLEZdJKmhQnD/+JJk9pIL8gZLGPjoiQoqgXRfVXsWFs9hsThu7bwQjDp
ntsneaUfztiqJqrPA1K97XFZsTAWZPjXY035rpfw+of3DKjBzeGYL8D15SsKQdCaGut7Uda2f/Of
0BL7rMpi4LGWyDrowR0OMKKkgfn2vrNMj4rzjXbeTaX24H+pvKgqsOxCqMXf0VZsepAstS+njaFz
4V/0LMvlYgRQJCon5XSPLdwGPM7qn6FADYb96PUoaZ5WXZ8KTTo2NfJnSLtGfC5gs1kESS7HsPzI
tW/Css8ws7yA53e5kdIgITZOUTsDtbZ4qK6kZ3G0qbHJUDcc1BOTubA0+3DftBr1V5PbIObS+c/M
wo2e9qdZc4Xdi6cvAo/PJG9ifV4BhrffiRigLygKIx0vMsmG3XOD5z+LfLxP2zLtlJUMlgupsb+6
jXLs3UkZIJTOhYv+Yubbf3srmYgpn5T0MiKwK+H7mvG2NgoHohlpr6oTnYMWg+mfTTQFcIohKYF4
XPp5Vq2gVlCDRUeYGmcw0xdRx4vLfmUmIV8nCofyoIl8wDb+fe/tKIIMXmYtz8VBDsk+p6KaZq4T
LkXlRiRFMJLeE4ebTAzalDMjc8dGvxP7ZHpok64PLDfZ41/jamL3ZkJyVYgZeXEYkH1qlHkC28wn
eUWaBplQFkkpncWXWdiF1dx/VasscN67hqSzqjhP5rqfAvS3vdzlDfCO5pVU4v0BM96ZJbUY5NMr
2vjJzJK0csFJU1v1SjDS0GQdaFK74viaPadMv1uyWOIC/2+EwTH4IxzkNMZ6N6AM5SHdiWxLOEII
aMdlhsWH1e7CzwQkyfS8pT4qV6Jpz+Sgb5TQNNvkkTrITIXPFzIFQJ2NFS9gZqK2BMC2ZZGL6brG
2gTTijQtP//IeweCVSH406F/nRjS0ezUGebzQ85zPhHOijSM92Ze5d/Nkfmb46OnT2YK865fzy7J
/VuhObGo/gk6+4mnhRMnMlAyvecjItiVCfC1MLFWrnaBcUiJo5ixgRBHWOry40TkEPsJ3YqgFMme
0nyqdJ92ynt+dVrXRTohkTcczYOFhKLbpEefxnzJrtlMOWRGFz/DQT2FtQI0XYnvBjCmSxddnJYs
0O1gVxXwisscyf4TJYSwOhhRVBUGKHS81C05ObcoUnnrXs9aDjP1rLXIUJuiD3RAG9wigRXEFDka
M+179INiMqJSJxDBfcXmyARcbVUvxSNqfm5D0Py2f25DOgW6La2XzfIBSVd+7hxqT9HEObbDrlMQ
btVwmWQvW3xkzjnZrDgby2u3rrGn9CmIcgRBLHCpBtjUxt10SDuqh48sf9rln/in7OkGT3n8j0iO
PJog8HVyC3TaIVhBF8FcnzAZniuMeXc566w9hKuUlNZKq0hUEEgBstjZIABBS2xYf4Co7r3EIDu9
gnVcdOjRSJbmlyK7oNuWKuetzRpOj3RBsJ3Y4fhUoG4goDew3VhQVWtVRIQM8TZFtG6Y/Kq4FAxy
4HfBIc1llmgItAR9khuu6aT1RgHzC2ZFZWYXQccMpDEy4314vU6vQMJJGDH5XjnPL6qeSl8IVdtg
4/gJILO34jhBx58e12eSoesGdowLz8Ikqz3b1sDpMS3Z18Tom6mAhpTKHFJ7eRGTlQv6OA/Z08zq
TmEm05ZMkK2b6pzqmLy8/d7w110Iy/uBXayBGstFMfpCfMxyrr/leYiX2/f2Hme23+7dJp99tETv
urE1rbRRoXDhNCj+n9PkylfhOWEHyu8PUg2U07Gh1yZ8V4i1Z6beIaChu4iiSqxJzseJS9hbu8Ps
m4dt1i1QhvWUosZr277q9IodOEeOG/1P7w8nyKsoDlRRWtlPR+wyktbpAyi3vP3PYq2i0ATghUKT
YWjaljOanXGs629cNGuAk8do9exxlsfb2DNYEk4p5hiK1flmyaNbNtkLEBtYoReLoi9dnb9S47o7
JwYdnmHnSvBQDPvadiSa+w8liA7GICFvrG2ixFBU7ykqrUoTIbX/srIu9grsiKkwDpH5C6gjWPG0
bJZkfPd0CDohgNKujwtg7G2YvE7XQJptXHZ4NPUzKw0ZjEP9F5eP2vAo1q3F6womufvuu/u+oAAf
5xeDMvRDviq0ciluW92Ewj3g1/5S7HcVs/ltyqP/Ru0tONYXnuVeDBf51rAAa/tV64uu1uXuVs2x
zQVR3vI8V+2+QeKQSA3WawMH4vWPu89hdhVXJIR72D2pSlIaWhsT2e1Yph1lpI4f1LSUO/6fNHwn
SrSUUmMnXnxkoZS0KjKtvHQYA3WqGk8mmNLrTuByZ3Y39nYuCUsDPN16jPBxFvJ+92s2O3S4vdGk
V6Hg0DOsvdwXq8weAN2/FrFZdbBFSqfKUdcn9xldulc9vU1Rn8xHwQ9KESgG7gp3sO9FiebaLppO
HD8a8LCDZrWME4K7tbzjEpP4SzZutKOXdJ936EN5QJTflNE/wYbVUPkCPWmrC4qONuDdtaj3Po1c
mpRLYkcm2GPmRXECzXdWaAEq1hwj+18Np/kqXSlf3RZI+fmlEY28Je62ifON8+bYTP/3VShiWE1K
I4sVM8nsss29HiXxq9mgwKUmJS7Cxke4d7tR++jynkH1xuKd3DrEBLbQE80E7WmcxDNRneF+lBGp
n/bwmbNINMidQCXT8nKcU29Bze4OJNJSdOZ26y4qu6O5MqJqlXZVDdRh3K4TzPLG6iNvy+wyZ005
4mTixPZFbNi12ng5XEjl5RB8sL1GknvIGmLRhwrUPsE5NeWpxrDldH7Vyj+bf0ArTeQ3gAVQlmBh
D7Se2jJYp57uRYxBydaO/F8byww//EXrIwoZeCxDWo+EpJQwGYYwcPHKSapTOk9l3rjTm88lPG7S
ANyMAEodvXyx1m6bZXbS8v7jSzoVn3Q2BLcIe4An3bkP8moU+q7yiAiHaLBdUONai8KwH+uObPYR
/2Ri2mwKi6mzDPQvLS0D7zA4ivEJNcgpy2WTDW3hBxSw5XciVnG6de9pIR+XMBn8PF3rGn6Jny/A
2x7BYLF3qTyBGoeyS/BRBWufRJp5UAGGR6Cp0+wurUIL/ZkNnHEZlPxSlTR4Wq+G+WToP9e2P50u
iGOhgVCD
`protect end_protected

