

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hajT1eUvtcpbI2tr2ZpQ+yt3wRoxz10Ck0HI/Kzj20i705g6DeZcP+FvEeRZMeE3iSuhECQss2IC
TSZjW2KB+w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
i/I1IeDYXVmyWoncZmW1nYLxm0OqNFHolb3NRcBcmjKOMCITsjC1Wrr+uKyOyNEAzg8LAt8SApGl
0BkTt3hGlwT5vH5JpMyxisp39DIoQ/2rHyhelRgIJSLTMOjHU/hpeFRg/8m17ioym3ZBfIcVRSy/
8YqL+H+Sd5EIN7orPrU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZwMv3uHNJwRn2Ww5TFfON6zTPNrPAlVNsMdpIyHdq6Uz+3GTAES373CyUHUP+cjDCtRwMjqRzGuk
B23rvW/CpivFPlGt/mLvn2R/n+PRdHgtaqKJEYqkidXp8VZscndj5Jsns7Mg2gtWutKvoptc7/8f
8ZVlv3hAdKdz/jYv3JFkYYsQYs/9EMmUObpsbPxhccaLaqAcMcp2DPumqvxQeqn7235qfdKNrMcr
c6uFXng8fnfR9emT//lppNqdkpAUWD93PhLZYTwVVXcjV4e16eyGLhyZTZ2QS7WZbPAkj35kG18o
nJcfgFC/GO+Ysd8/MvmMgbWhQocjtlk9D4Q++g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F+8QLMkCmxgohq3I7y+DAO2INd7sZ10O4AWi5yw/qOjlH+MDCzvNaVws6hhgvB6On1+CWzlrQ+vz
8M+w5LD4ga5aEaF2/H5jzH7q3vP0dvfZN4yRMhZ4TVDJv5PjxyVU6bHIlNhOrXl3MF1oGoVIjZ6h
IEpVBqdC2ShJgsN6O40=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Nc2OtpFQZFg8m9MEwwFrTSX7PqIQjLT0ImG8RPKmLuLlbhKyDcq1HH6KjYM6DTZXkQahd7sF4tka
CU4JtMixX4Y8KRzlmswh0FCLw/Aoh3nJlGD/KZ3QsZu5KBZUxKy0A3ntWjfTg1NNZ+tsdv0ZU17t
6SODHMUk49BioUo7eB0yCXF8PR27Zd7koQvLbFKTXZjGgj0ayut3GjrNM8A+4/o3G/elRT5WscCO
qhmVtlygfHoMk7BWSkupTlNlfF4owb4C7/AqdxneLzHPlGWymyNm6olzMM4lJP0A39+MtJZjtTaU
VxxrhX4xVaQG4Msik48gN+qH3ORiExl++4Wttw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25536)
`protect data_block
3HwGgNcLtmr5PHt0/F8xLYWFkflHha6Wz5i12FZrTCz7Pn7xvx/JvBxlhcSmeoTF4+p+SBml8G/n
gjgfQDhteEQIN30BO3GnNXmXrT7RRAQXHk6WbX9x0x+uC5lq7UFGVLxlHwoaBsmsbO0LVGd6Uzxf
ieZkf0PwFJWl40iMbtDCKIy1NHc6OouQxWQKienTC4KNgSVurHNwVNoDP/MdMaDvwE+ZAo4PP6Cy
Js+WatMFMbjLVeq9dWAgAv6quTRFCiod63FrB19u8f6Jjj+aGkjKkAUGxupiKllk3n3y6jJ/s30A
M8dXY1kxqyt7DfXLL45N+Xmur8XRr73oF3yomnUxqBk9a/ag6vZkLphW0UYQPSUNqd/VMeqe89xh
spDJHse3xuIllCklavgkCDudf0D4ul+MnWH/5tB9+rFkNO3ygx+vWRuLcrjLKNsb5o9zFm5aBuqs
7v8B9VI3Z5W0QkNsw0u+XZrdx8d2tRdIr9t7L3DuEkaYUon/lSqq4tpuQJPt6sXXNGc/oS8pqjBh
kg528Hfpb+iZsfxzEdfOavCK62OAD7/wlcgBMSMWFMoevM7UHdp2CLfbxvuGmDv5Zc9pexbaSD3r
6dZfeuV6UX/cQYNGcCSu3ggD/4LzbzI/hkq2qTLXy9gITAL2cJv9Gqcc8BfoJK8NEkQYvM09NQNr
JkH/j9l+nMtXnnI+rh85m3XuMFI4mhtrM+IO9unGX782jzqq8rJPG+QXq6jOb8Ctp2XjZgIOzHhm
NgPCjaiqu6Yb89vqj3eQntRxf0C6O9molblWrfRTLUGozK+4iV4DmcCt3RL9VRSsKj2B4K1ZTBiw
GoUyJSojf8dF8VCcxUD5UBhOGC8ktKZyj4DQbato+moDL8wsncotxv0xaERrA/l2RetYS45EnKWJ
XBBJGybV9dCuVSgG3eBnJ6nV7h22k1iopil9QE0R2nb6pQJ/6e+GV2vxAVL+wwF8az6qfeZ+TPAo
9g5euCEMrqZOGPoY8/bNdHr0xdDy7Sa3RyjIUw4VzwbuEW/I8RvnXMAZwaUQuTOzlAqx7swJJJsO
dXLiAtwLLpDaAXiOErnol9Uorgna9OFsSoKY8pwBmIw7mYmKruXaQdUtj8QssNHSXK3P07MDcT0O
Occ6dC95YGsJqEaYHEbcebAzug+IPrHpAFvszs60DKcCkiRKCSLoKena6x1C7UgrEyd0DidsSxqg
z8g3wp2Hz8hI3+mZzy2E3vqDIqR55gUjONAWysyHk29vjbWruNVbriu/ZfJAnNK5bmcV/i9L0La8
9kisZWRrqAGJOren4D4KaNidEWlqKGln3+lLw95Q4o8CrFUuFkaQY8cMMbWNdf2mlyYPbDJX23xD
GT40BxtaBIHUx5594+Ln/rt3msf0KKGYA8hefI/njJJ8HA4XjWyfL8T+05Q4lHBalBK3Exx8FIiK
tJGOaeeSvBIj/tNUMpENYUCEkQg9lTmNjY4DmSReQBv9ArBzZtOY9MfoWA8PEVN5ipRJ1v//YLui
1pINvEhf2BslcO1FlDW12l4+mKAWws0pfiBX4OgolR4nDNTewPs6GkDBjRF/q+AcLBkd+upqyUOh
TymHruA4Sz7hr5h+kjErC7gNnBkwh07xn674WeDAEeXx/SzwDzj6e21xPhliGhVKwItA51vsrf2f
haHi7cgJAGW/KJdqBcexV8FXt2hfQDsXOXQt/ZMIjSW1KLtfWIJ6a8wmaMohkWPF6N/ENhTGsrwe
7dgQxEkkrDZkYnkUVgsIL9r2Q+RqbOPSwhv4BV60lVQD+qWzmrB41C58tscTJeP+NMW61VY1BS4Y
yC+5ilm6zPvJctOcws+tXNZSNkTBp8KubOpyLbPdwbFzg8i8Yid95sGShxqC4xFCE9Rn7NndzxlQ
/aWzwDvOfmsz89QtVmOQhBut3WQrzQiypArvu1CE8Zymfi8KS/dDTbaIbcEN5okdngxPS1J8WTHd
c3B6dZLS/+EeuWjkYVaE74UO0pyfyVz75hkmRtEovWxrAyxCQfmnr6F+x3jnjvNhn1rtcaI3k7Eh
6QeZKJg+2sdMOP1iiLq/Wf7EzRAkYkVyhn+z7wvnyNSt34Z2EpHoJaJHDfGxMmxQQ5/bFYK7Zrpn
W/HPjwyo30qM3m5ak9DxMovtHWoc5hSgaRUYG4aMtLP51eLrhIr4j2vA63vPrZ5Edtca1+RE5vGn
/vj2jrmDUBLXInTJSDBYJ5e1ahf37XAUyesG1XN2hupTnSnS4HvMaVPiYwcO3B3qzlcEP3nh02PV
FZeE3nA3usPGsdEvPeKiYniA/Bk6AiWw/PMlnvIK3c1gqDhcMBKi70TBj3AvxvoDHNj31viAuv1E
Tj5W/Qsh1mT2XSMSO1LJIVFbLvhpugrf3VPzcwJD37rOPlWvujWwhm1g1I0klz/llBbUCZIrp1HV
qbjO1F3MjZ02xVr+2NXSvklXzN3KEjm28MvaD0/ysDyR3+n5JBu3Fh50N7n9P2LBzH3dTvpCxByO
I0GF5oH+PGZ3cgcCsVParkcJ59aCn0qGGe6ANWvjeuG2hV28MVc0JR64eV9/dsGjvomDc7Xg1Q+3
zMd/0dNFYVPWDbzBGB14BWh77BlBw67e2Fc574Gza9iA1ohSDdsDazUdBIJh0BQoB7PPh3kuOKZV
8PQqtQMDo1VQZPPJFIPmOiEx8nlJTpW4OyMWmbsD0Q3pW4oLGVkkltBh+DhfmBTFDGRm+7kjPdVW
0CwGZK0mvVv1fqt4JTxVElp/X0nvkcSNR+1CL/xcFPYsvMqlZhioEKodwoQhFzAX7L8HT4DSYprG
DM6Fkwq7mb0TWnK9B86vZQkviYtyIxX5ekCBWmzAeyBcv8cHoKyi/FDlY8vhk5ruAGFAAM6bg+BI
ltZpGeEVHVY5XruV8sh4VnBmUyUBfBDzU/JdEcsduYMsS82D1XfUe6Dbgam36OxcZq/wIvggzGDd
+3h4vbFq5L3F2BN2oZ9P08oDKR1PElv9UQR5r48UKK/08lWAJEdEtSWZ5yGcCO83N0WQ6MwfNhUJ
KJipildfkaeRFdoVCpt/rRuGTxwygyZRAhK1R19idmzlmnIXj0kBv632Pww9PnMwYbZgLaSJAeeH
WhaC95ySVmF/1PBXQh2EVdTXnnlMqbPHw0h9kDdm00pNlqPvQvpP8By2bjs9oMIV0x5Uk7R4iQ9c
4ItQ29lHaRjCYQimakxRuJMHGKDePkkn8PaYNDZp/rUQDhvxRV5/OVdqAooNVvBDawahNK+lcO3S
qXJ6encqCyrmEXFogIPhiuNdshDA9n9dKMxEkyqIQX3IzIm4pxnsLx9WTqzwDHwuMNWrmCxqHUWq
ELrHwSbBM3c97M4dq6niEzMGb/QZsvR8OTGmWxSS4mWIr//+quaiJCjTwmsT7C2wW1lobb4K2AfB
zZEvQZNHyPpPj/z1lggKLiL8C4FzZxQlkVb8U60bLK0HU/XDt4YKEhD5dgqAHkwRs1DkhtvJtSRO
w35CVD3QKhlbwPH/CXkg9IEbxmYpUS2ylRDjvxmWZ76BVV1mV04iirYUWahudlycRE6aUCkN0JCl
QUhQJ2rZo9IkdSa2Q0aycbDse7+yoia4N+RcqMpWiBji/mJDNSaPHzrU9lZ7h1GVO5z8hDLZsyyy
m3NabQ33uyM5eljR8JqlJH5piG/fFcb/09KQ/OZPW5cYDPabp8XIpgKjurZDh86mlhZZn7Ryn8f4
UEiZuJrRq+Q89xJL9J/p0IXkKEVqs9YSqf5BSN1AB1jYGNpXCkLGA4sqJys0b4eV6lXokI4OSZxa
D203xK6AiYlX6ZlTaEAjeH4XlEBYVMXAlc6jY3U2iDGZil326k292yoQ9XzzbaT/nCBv3t6jxkeD
QJ6vVYhSJRoTa+N1FpC6kaqnXkaqg5UMoglzL34QKR91zM4U+Il6xqvAzKMdV2q12xVIjtUd1BBA
nTI6vlAryFt+62oz+mpePRcq2EuWnxD0HuXMZ5rwz8eoj9MTbyv1BEMSvBD7ZmXiYDnfwLAIiEyg
mOXKA9c5/20NiUvs9htgdXq12ON1y6QotOnrNWVZZQyUeoNXaP9RoE0ipWSKxwTpALWlpqIsyafz
plZMxGL95wig9heeQpoDMJ/Cg3jxsIetad/s7r0jsn4G2b4/QtjWfX0egFcFfyiJqf/ei7DuQ+Ft
P5yqMSeRM5V+O6GZlD+TTjuZxZOK56uEoF3lRd8NhQhPnYsg2SeHGdak3DL94X2ixbDbg5027/8f
YWhj0m0/8TrL2Xgm5XmS8B3VDTkqs97SuTIIxPcSeqk5W8uFXeHktSYejQEK83UyHe+TlVQ7ZiQi
5GbFu26hXgwP+SDxwXLdX6fTScGEISl2yono5nBSLgcgBHHswKFjQfLlSs2XNHnYWuQQiuTR/SUR
bKIuTLuv/A1eLkR0Bvnk2M97g+UGH+o1AniSHkMH9dHbu5ZfTkR9qq9dv8CNubYYNqfqM7lsYl15
zuCY1WRqaPS98U2tUx9FiFgXx3kwK4t5zqQk3lk8aWwHl5aCSFxwy3w6vvJBIs5zElPyZyLKNQ4l
ZQ9O2ulEyugMXN6U6TFDkCvynSYdoTQqrs848hEr8Eb3Bs3QQ/CrI6fTTF+fmZL8Ntllk8z+cXFQ
qOHLO8lshxMCpTcuStGDNpWu8cU1/DJWNpG3Xr7jpdUKWdisFX6RhzFwu1YYIqL9TPlrgECeN9hV
a7hEwKkX9NLiqVFfi3Vp+8Cq5tM+An/ej+a3afqKd6HSU9VMSNS4oOJFMwm0V2+nOF7fsGrdxuta
TpLvY+7OwgQR/0ZEvu7mjZtV0OAUuOLxJJeoTiwe4bq3CuqTOag6SrlnNywyLGODZFU66Tz2TdeE
HEwzMwmdSF+b/3QC3eYxTTqVWiTjXjw/us4XjQLO6stxqXDBez+93OO5RwciC3ObpjEM8mYssiyF
VW61Ml/EqBIgbsagDxuGXqO4nMXOssUy5YAcXabT5Bl4sdC0UiFLFNNoL+a/sh4q440xitW8r0H0
tYjpziX0+9OTQB6vjzqfsCq55XGRCMaGtovzNQAtv00lnKsdDvb8g3BSmwbUwR8lS1tCpkL6QriO
6V/obA8L4fgk61bW/nqqVv90IwUU4Zoo4h/ZKxqFj+TXLDoNWFZXBl0i/TriML5MBSxkFsuSsk2b
Yo4otjtQvzBza5ysDPayP308V7IcnIsabpD3I+BbZZE/gS/lRd/nyMxTixUdwoQnY55t0E/do3pD
eAW3RpqqLaoM20RKHRP+XA4AUrjBao0RJC/CYhti0NIhKxsZ709/3XME9IgGztFAW+mjjSyNX7N2
u8OihFw07jW1Y5SbtasnmR/23UA14UYzgOxoTo95CqKwIVH6iHyJb63kAobjy/sSbTg+5C8Lk1IF
SXBps46b35r3q8LgPEoYbYI4O/TgWR8d0rCsK0t1VfAuK41Qh0F5W/auE48W3XCege7SxvUdGmVY
2cL23KxJoM+C0RsXSQAPCuihv/nCC8daWnomcYGK5q54aZNhISFsdtLv2/xb8NaLH70H8fhtxZUD
LaXpNkSya4uOhnYaH5YbfmcemoM9Q185vikw5Y0+FNJvHcrW6Ry56KLFi7EkvVDR6DiNaI60050L
+6O+Si0ge4tAHFQdhY+T5Tqf04yuQOP2s0VHkvmsbk+lsdWBwUhxgi3iZM/RAXNGVGqb4/6sWpkh
7f9CycnSQ5RcsfnqhF8BkdRbFFsOC2PqHYrhipYVFQr6VA2N5/rVTBw/ZqfjPiO7Nwn6+UgkaH65
R6Et8I8sXwDaaKq0CsE0KidJnWJHwPnmEpSnGx1pw+yDXHE498g7VEJL3OAJfpl9rgraGfL9n9km
YMnsa60u8FfahvVAItTuwPbkX6AEJBWNiT+nKTpHkOClWDqyurKNqsWQsJF+KES/cNrRXC1RiCnT
Tff1Kwj71r7Wpd4pezWy7XaPaig51OgpI+mcN4aRYxMzF75pDq5iuMdkZr7Qyvn/70RrxScJRLCx
MOp1p/D7JOOAae3CM1kAf/VnjqQqoKEQoVI+bHII2tFlubpm/L2iP/ir0WMjMOJ8+lm7NY+veJSy
uvsZGl22d7zdB1VeNPHMnJhXA4ZZgdkbG2sp02EOw+f1T6hJY7UQKF2QoXwMfWhnXm9al1XWBdcr
DhPtWWfuNUygWknRFNN74OnVod2TNiTZsuiT4qQGhZeebH6txDVOzEG0f5bJT5WiBE76mRxqIO7o
dTagg6BjclxkQQcVmrUYe+cyGjney3btSypev6LunHfP3qelEY22DZogjtMaRZwodrit692bB0Mv
gu9liB1XVdbdMu2lSDVVonBUWoWTChkH/gqG0rGztMUO1jt609Giujguwpu55uo6meFrL6Grlxf/
jAVRe0YSis41bhtHRecDv++nk0AH8d5YrMh2wzGAVldi+CRF2aDHqef+MxF8ZsTOOOe1QBoF/Tzg
TTB1RGXthMhwiRoCFbZTbuLy0eojm9UeIEk2nl2ApFBbVMMo9Ptl6BupMmypWTR4h8SzMr7qtf+k
sBzuYSGMV2qG5tYV2IlPBnMQT0HzPGES5hnhyHe8fd9mE8ZfA+FSAY0lWvrQ9jD65kVTHfUw7Bp4
44R87t3Z+hLNgGiP3GprtALrggGp+FYYJV0HXfo6GkHQtE1bEI3dNyILc9l4CtwROtFowLGdNrl2
jGMkTR7cIRFjX3Qhbe55uPgPoUYBLBGATsq7VukTHZB3UIrqhOxQI4WoEl85lYIniyF5ZpKkA3b8
NK+0VAOU2/hPFYGAfh9/02+gVwosSxCsU2vcidrJeU6MSd7nTTbRU+k/0s9JwQFTE+UtlVI1xT23
bKChi1T3yvL7f2gU92Xan/xBmEiuBpxu6cs/Wzs+OQW5zhpZDjG1vO39EaFXEEWUIanJWsKKniu0
jD7L09FHMPAFSIVb4QiGAKnHipZcN+R3+EJvi4QXC0mHN8JqZCVUfUrp6VyIipcqPj9GNhQrgJXC
dZJ1KUBTKs+F3U60OTVABYfHDUSBAm/3u5qw2wuDFwp65IMFkFODs5zqbTj5OdwV0H0FoxNIYuIK
dz0OewMibf2jCcXBydMuEFt3xHQ7BWE1wud0I7R2ZRuwtM4tfLxXdvOjHjtP8tew52SQfNqPDZZM
kV1lHHRI3g7HsQEQgY9t9QhZV3y2I22n8RUrRLUftFqaxPxbl2ruotK7gS9DavP8Sr0sAxUX9IKQ
4qRgxvvfswOu0g84qc438sdLCLJ5QHk5vc/TR32iBfeHgRutCHdK3R9Rlun2D2SWluYddplrJh9b
hraZaYY0KP42sf/lukSWKGI8AFSErG56KfPZvEaogJXvHu8b1iMNbJ1YWoFbislNNtNWoZ6JUzHB
E3R2mFrpiFcTbvYBIk07LzMc/jy+ToNveNOZZhO9G7Dzd9Rq+tPEA389FT6BRvTnFnZ0r7e/uitR
cqrNX0zkhPiC+GKL2zeAJyTL3cXDScAKQB338mla94y6023fj2ltbB3ddlQcLxW0nVdbrHJAHAY6
PEk+WaRF/L4Bd9tuslyYLI06eHjG4BgGV12vnbyHlbHGOZD2xP/eqoRmf8+SCJpz0pop9jYOKzDa
uK8qc5ZmxP177L9DpPoJ+/o15NhlsRO9mIWDf4sEPUhia3vHYqJGzvyeR9UwbqGc30s4XgBclBTQ
mNoVdD7FZei+lKBqqZprDWeOptfzFP8lArAD3CFpAm0wXezqn6oDyuMv4U8Vbp2D2wvvZbo/i4tM
czVk4kJ3Mhkj3ztDrUoT0KeYjACqQyGYyBKbwjc0RAb2AjefqvzU4PbwGfQ2P5WXqFnwM/uyZKdD
UTPDwKIZ/URnemb5/hnVS+DmydTnmTpazClrwcx3STZ9JSx/QWBQ8IUdQYMtAQkqSdtwk77IMQWu
DrUT8iqok4Ry6u9E0/rT9FQGUtKDopCFFlWT8FFAl2CsVopB7EjQVOZwlCoRgPCAaJEZ1Z3k3J7B
/RTUgKkUoFfeQzJTETkzmNuBc/85qt1tr/+11i2Opa8DWbvAx0HyMLOxYO3AipcI4M27AeaB8rK2
mLwTGLf69cBbCzSdbqtK1cME8M7kTYuN/g+OJR66GnfMuvhnqJkj5LKZqXymbKjLdDWEbFhhMJXl
3j+YjdUe8WNBU99Qyk2/qq04MGt/WXo4+zCp8SXDDGjviBqXO6wDY0o04m2RBhO2i/lpsYmXslO7
yecjjgF6iltOp4vZoTtwcnXkR+nsjgiHK8LN3XE8sSAC/fapnbjHDzxdqg793aMajFljBXbArUCg
e16O6e946NzKz9k7MoOoYhytxNgJnMw+ihZrKD4HunMBi3NyGMncEwJXXavOtwKLDTqWfUIkQG0S
9K/Xp/M/yCVWP6Db8Rw6PQTdT5f1TRx29UuqKuJI4ZBIeSaZGOcecF/Z/ph7bMDfBfKDfclv0P5u
kmBXOP+rEy3zsMVVB/2YjJ69811OnUT2I0dQ5y929TfEL1DlqWDhf++GOKXDlQORoE7ppzjTSJYw
XkPCxKOvfgj88l97xJjXjUMjCb1NlJ+TbVOfOriE15pSRAD5QFJf8MOGVArsKIJHqHqHbx/AuDSq
UyAMRICFDbUn9NsUbEbI+BeGg1izwNmaLQoN0WR1ZmoDud8a6YIszMo1RW0+L0RAZ9CNyCsi1Tyi
5oXf1AzONRYpGpLg1YmlHpbOjUMsagLabCQ04gjt1+DZTnksmzlzb8lP+zpuRYTkt7SnpxJkEcMb
OGMBiy4DEKVHSR87u1ZPXbw3c1+xVtjhrKpEM7y4KapL9VLqwgOgxfYhnOyih80eQrMgQfAWTjGF
ZGYRcOSi5SODAnFPlmJex5n9i+ya4HpNdPlVx+DG53hsme2c+zjZhVdvZoFftjcPKL4UVUfOJ+sp
8g+y+lS2s3YYT0ijOA05L7yKmULNz2qM+8erf6rAgo3kia4+J2MY0K0sZXmKO5dO1JhP8L5iG4IN
9m65j3meIRrJLwE+i5GWQA5d3eMU7pJlMeW+0kBpO4oaAAvdB8cdlhGgTjMz8SbINmKNfgzrl98t
XZnppzzd1Aiu7CahR+e7qzjfQBJGm7y/ox/RwNv1+XbioZ6Hfc6gIMILHNzHHwlcrOTCxh/NcaL0
hPWfpYEJcw+fDnatN0RxYaqPddcmqKHYETyPCFpLfEOrTUl7BeL9gsGOjHnfG2EwARU9u/cH87yR
hZIDGNYt6X5yfd6ictSA4IGZdLXjM17R+bNkq+NodAbNRDThOudGIXKGkMB06vpwz7b8nS1TMBoz
8eZ3csFXvgtin0DliJ4k9GuzqJCVVUFsDHLbMfATyBAeQSd9ZsQfuf1+cvDvV70SvpCaYQxxPJqV
chETbnJGCfWKuAQWkU4+ILmNKAQX1qI+qkRIntTj3/xUzx7bx9q9a7Fi3fANYkp8JEMYn6rw+87u
ku/dSb4QGLUJQjN9cKpm5XAmTbo9abquNJfJTeWIH9loPrONNRuoXFR+n/+ORcgz+yYsUudSmRNx
BhVxINKfkk8JfU5mmoNuXEnuripKgkPSFkekWxv88QlKpxjZ+MmO3oePq/aWpRpqrVO1XTbbWnyL
V6pMggtZAslyjJ3BscBGhf/DVZJEOC8bqHvJtLi2dgHNYrIKSxDwuRXDQiVJ3Byh/pyheRg9Wzon
7CIMp9TIaB5tzznzu8YJ9KonnpURU0WIGnFvB3Nr3iCH6WIgTEsQNEyXJUazVMnSEJclXue2yTgz
7jY0ZbngAQlaTCSjVIoBs6wJldtGDllCdd5/El3tLiGp/L6vicyWN8zfoiONXWX3+YFDTHhTVjRm
/9+fxX4TKaobs/cgFi75z6F1dY1JPj5mzJq9ImQpQ8H/Z1J1ZZOWXW+hjD77W/sHYsUeOBAdUz2f
SnvNjxuDgvl+HzctfQ8UrUQXKhFyMzLKkL8ZGXyDQPVJ3EOjNBOsVhZjD00S2YiwIVSo8jFARhAI
E8u2ahrKyAwWENVWsK2yjnMttedspzIhJK6IUIpEO5p2L7d8wcb9jyPygyj9QO/rMb7YJ0fknLxX
2kQt+m+CYCxYsj0YYvs9vza2I5Xpbd75RpKKYJbjbk4p2iNXLjeMTPxbDNCdIvLXaU3LDw0SbbCY
doIc3T6SrG8fgGM3fc1zAhjptRQX3ho25dyvJPKG8skFX5oJEc1FfLhoGYpScSzCLwEc5jaH8ceP
egFWkxyv8gtHgUh/Gr+7J+HZ/iSEepcbQt2I+Feu55zHt8E+EmbN06A2DHhMUf8KPS5f2ELobRRf
9HQVlD3mEFqDBnG8TEpRypuKHHW0n7JltOMltNbMfNa5rbKR6xVo1hfrlBhqrWxeIxC2er/JdMOX
mcezLpi7dCt1g8fgBK9LCn3rWW5GnkPzsGJ0jZgPWzyr/R9XdJWXhLwikOji1vnYTfVGN0DkO6TC
xmEbP4uiWGVk4U2mFLclRBsjC4Y4Kd1KQEKPEvrCdHSqtc2K2c+H1STElS/OzysS3k4fW6XEl4DH
vjM+mgqWG6rjEkrw7Eg70OV0fgoYyw9TAFUSMIx9E5ZYiq+Wf9In1zIZTOCK8Jj+WU+9RMs91QeB
yEA6XHmPLbrnh+1jehlNnVGM++n9TCyH3byYazKDkuKjtF4Ic5lSz4ouNmvBhnOx49uM+EtnES7q
BSv5xXFoTYXuXDvPrq9azV5vw0FWCshsIO/FnhBCd2gKaFJeEgYmbi51qDOViFOP+adEawc5gIyz
b6/6zPdH4xEwKP/uEXtBtWamIGRVg9hPKYx6hQA4b8p1x11zklU6SErXUiW6EM7PX+iXRUkgHx9N
7cuDvG1OwnnlBXlQ+NyHcSRbZBkj26GSM6uWpKBdRpQxO+tFQcxjE4TTU4mJ2zS4ZxJ5/15Oi+DB
w+MAKhg3vYErTho3K0PvhP210EAMjDyXx98y18xcpfS9epDD7jJa/PEb9N/60vhJ5SEna0sBbNrl
7PkWe1B9vbWB/u1ULWQ7IweloIbPAs5R2UXKhOUccv45smEc6mppcJWR4ELYkAYpI7lJMA4Kamtv
PK/yasSSoVaWAzFaO1aV+jtiU7fr1QqBk6Odq4RqLPkOJQkxqLk9bNhIy5KNV0uh8+GE6Rehn7gB
04Jywdk85tz11y3qAjiq2WVE7nbbazpe0kzlC9oUIJmcTuTxxhW5o7Ffy/K2e2oObK0QX9nz5XFz
cJPLGDW+hU887qdKrvhHLbQ17VJykDbviP8D/PjTLOhjR1U5ApyB4KeOnVWDncV6rLLcLnueebAz
ip7WUHiUJKs6JgaDp89Uryb/VqpTXmYzpfaLJkJLBRiyylEhir1enL876Cg1ZTfdMgoNiDaAnErU
iz0Vv5B+2DNNPXezbxXlZK4siQ5uHc7SGm40ol4dMsDzwdLmS2/UYLWN+JilOe+ZV/FD7A1scmQa
WYYOycY0tRSzLSeopHvMg05O8ioZuDz6MgJ9vM/AFgnbX7w9yigy7HRhbITP/NxxrgYaj9Hb3cQ8
eTouyn2IVn3NRCbUVrGC6rs0I86BCMXogLiwxp0c+UdfKbIFqrNq4Kz9xS2JygKo/MvsX1RVm5Vi
Wp1Z//7jW+XpmkfL3rUXX5ToRfS72M9CFvuHtdHVjA+btSWExdWWFGvlmjHBemGLNG2MZUgNIejR
P+pkglfSXfvyCVkDolxE/6s2Tm0Wm0fPVOOURB3NOUHpXEP/C3djcwuZWSF+8iWK9WNQKkOldO1M
OH1rdCu+OkldGBc3G5VOpZQuNDadyROGE3oWASnoGb2YVc7quqv1CvmHQdO2IxtsO9lwzSj410o0
MDGPpsSQ6l8mvvNbMjJ6yprFrZdAThLEl02Iz8avMC64+D/48By+4Qt4GxIYdEz8v1OFaAWEw7xK
XOXEt8nOyfkKEwsoYV/eL70KN/QWJScLqM7FY2ArCT1c3wB9oB+3voUNBihI9utyoZ6Qvjcz3raF
WqhzlQdHmaVV0zxaq1HEalF0SDGN2ThiR9yBa0n7LwdYSYyeQLd3gYZHvY+7A9WGYGrkdOoFifua
BddKUI/siRLvfBF2c22BkNnZCKiw7Rz1TcBGQjLJR1kxX88ZBhYO6osFX8eOHyahLesA9cHL+/M/
djq0os5XZovdMHwulqTSrd/kf9CfFlhhyVFu/R+Ro38JbzmxHITPBkbRRNEUNIlxZl1RlKTwU60U
S48/RAm1NFz07eJw63ZMIdWNtMAnJDy0dz7vhH8PZ6RmdsQXL/h+ozZkURAzSfMARB3762pl7gcU
KTdd1rIvaCnUSYRotfVuKTipH/FCj07GCp5sK7lfS4sfc/wLfmGoeEwJqj6tAAIYe5LyLodKZcYg
J08Qwf1BIr5a7qZg18ESVgg8YDjuYwOKaIDgjLxyvCqFbkooPClrWxQOxkWl4d9kjwMWJ+bg3xnU
4N9ph/hPN55NZQAwnh8bTcVhr4/GjTMgEDKuMq75qwd4ISc0aNSzebQOdSK7defKAGYPzXiUGrbl
Ar/9pYRVWVevyWPg03GpEhYGzgMpWHg376jma8RbwjuHKD6GaU1sEPXcGGJbB+XTRlKH3TE2JtT9
ovBBmE8zeDGG8D9VYY9fqn/U9Po2TdrWtXKu8bc9NmSp4/s1DkWjdOg9cjWbMctwbI3qJh0cUXb2
93ENj2ynAVYOEvQ2NbIwNtET6oR4AQ0fSNX34KfbfamUeS0nHsCmBZHNQhxcfwKlHe7sOtvxV/Lp
q/kiF351tXm+m+Q6pRkPiJBlr78Uxpx0mjXACN9NdPag+IOa9QPk78GHT4RxaRh8AQiLbfqXj68k
3akN3vMdtDSgcu5F2Lnbn883r97TnEk26XYnRpJ7UAWc6rxtgi5HabrCQlC+TVH+v+TKecL2EIF3
dnourt0hnRU1njtZOAuRmpcUNH2iTaXEi0YqFYAutu7so6wU+WmoU8GuSOwLEhwP85KMe2DkvcqW
xeiMgThNcMCNMq6Hpijkqwr7BCz8ncqOy76p/rC3lD3pSrMDrg4N33N5L9YuVi0DXPvBwWudoi7D
OLKuAbpuFrumwbsus+VWjoqayRA9kruqV3dMqml5Ca8y/V5ft3XE5ADdHLBRu9goYZwk3SSClu7q
nVHO8DAZm80jhyJ/3JxJeLhMYz1t2gUP8EAFASI0HIFSf21Sc8fgIoKbN4zRSkictCVReQbItiP4
D+EpMzatbY2xQ9zmr5E56hd69qR8f5sWMwB26XaW2IENMvsznvjoeAqq1kPs/XjZHoS/zKsVTSUH
2piEzwI+M6UuxIpfqDf5XAncrTKPxC7hv8sCfYLUWQ9p4VBTCb8PHOz0QlyIyETJrRKi/U7qfd6d
574YKn2mF/M50s6thkEbrgtkQe53c6eKVztJ4JJA8AOcgufPm3VC4A9oslXtz67I3bECrXPT6Q1I
Cot/VMWYNVwvqMMNQ/0b1R1HVpH0j/EqhZ88Q+Hv7rviCNo7gkOc6MI9lDRA7z1sysfQOFXo1sEG
JQanujL/cZSFNQZO8fvwftR5k8WD+DcK0r7gpxkraCmCRGcEyyO9lS9QHKzwYQT14oTTz/FxMJQd
G+SOlBwOqnnSguhF8f8Hongf9B5bHkEsjXvjMF3WgCvSP8hDK/dU7dCnNYBGTGCv07wb1BDPBAOC
vH6wKw+Zod1vvcYvJv0hToUOGqzq320Trj1DUdHOTojpzfvdW1QjvXALtwCsxq7EbFPkadtSreJX
56nihm+wagZ6L86pzQVpiNgeSaQXJZpZz9dvp9kReNVBX/vuh/6tMew0+HXiL7Pf2Pc67KFGF4tG
xP29miCNJsvoxNSnmnr1E/x7C0nKIxXRhr4FzHjJjpHXv8ebj1gx+u5b8XdoiZZ0NXSw/Mdy6xYI
MtWjbn7xp8qEDz0RX6bU46e4hVmTThQSL0PYeD5pcvns9fR1cL04bWLW0b8AoIloP3Vh3QOgrWUL
ByKU+OsOAAQPAf/dZemcOiuvrIgvqW8jhA35vUpUwf8mrrXh3HxLKMa6SqLmDZ8u/kYsGIeN0jm6
ecYOcQq+iQkJCEF4mhodwiTSTVj8K6WcR4RALhPZzQZqwazaOhqbsBzccwfe0veTW7l1ur51kXMx
d6bmccmV/c9vSwK/9qDNOlXKjzpgenDQTl7nJy9RJm2IDQWTI9L0EUJpiijKhPMf2nDCudoxEc0A
PW76dG7JaMcZRC8I5mWM3JwZocXe/4bxKYNb7SzIj3GoUlPw5oABnTL6zuM6qPF0uYxpuLs5oCEb
yxtqYAio9O+UgV2CUtC5XpoJlMOeSjHfJQYVTvYx/04DW2ViEevn6vZ6sMfbnPQ3+o9hQwy9/aOJ
zr1YJfZ7KWJhQXh3ceJWV8tLL77agvopw2ADlqvxGiEA0bLqux3lKvpNaWDXnUhv4h3yU0VEpFOL
cz+SKjzCTV6Uw73h0PD9hq2civfyfG/DlFQVP55JeP7nBJfc7JeyGOyposzSRSdBKi+grAq5pZLB
X5uGjb/FRF0xbeqfmevh2YveOFJQRUwhrh5hgtDT9UusQ4UokLPFbY2j6TtU7eTuVGuvNfi2ocSu
KG41GQYl55z6B93QREgkpdErpeUsL9b08FvbyoYZ1Z5ZqlBPqW4r7zCsddqrsedwnALaWn0t2Bh2
ljqB0OxBamKpm+6CZcJBsCM1IcBsWdg4+t5QESTqT6vol8Y9oGr5K1bHibaxYV2ctly4Aj53uX8q
aarOShUZz91Eb8XnCrcE4/0ptqwk+zLYryStmzm6jgPzr9PruYwH3CMdQL3yd+S+UHDvISKhoFOV
IRG35Dw0i+jgcUNHMDbWk1Hgc+N+jfuFyRPhROj6AlA3dK8fYBfBa8LHex0lI/yGtlD5q2F8mkSr
2xfIo5Nn9jpXQU9LCkLDm+iKuiV89bI90EtU/geFyGUCbxqQmpgROxd4xJn1PxuiUqsosQT52DRN
8jd/ryPdwWRaKoHGznXQo/miGD1WUayFXVUEKEK0ryRn/pp+OWEnK0soidZuv3FPw+rbC6gFYzNl
GXsBRCQn82tQnULJgfx4ydzsfR48YbQKhONm6L9gQQ55UCNjFJrvqdlYAByW7kIoXDXdVCdAfqB1
jmtGqr2IXCadr8xtf71y1H7ku9zXmIX6WVRw/MbYFFsfV6oUZ3WTAL1FnbW9CnYT0pNQatb40vrx
V+7q+v29loq/D6JgpvpQb1Aoc0X78/mg7fBNWBBA7pc/gHIScS8w4TIyPk5fjlcm8jhT+KP4tybs
msNTYlUdI/yTBKbAHYm0+FFyLCX1agpxyhxoJYBK/T2rYNe1SPmnbhacwh+M2zhtQLp/d4juWxKV
JpI/0SRrvU7VVgTRjTJgQqSyhQOF2NwB6cg2zlCEpFeAWjU4yt+RmErFA3eUxzEFg78VQEqgGi4K
3WOT68oSgjGojtTeCq0kpPb7Jwrw8jJyA260lm1Bxhb4B25GxBaAij6mBxs6iHh0L/1tcDCYbn6l
fXjFlxNYLcUxnqaY0/dcPfgzKqBL9gGY3ElipIDGui+iR7HojFSIHna+0s2/Q842M0FtBbugg/ST
euVV7K52wsnE9ADLkgc+veAoRsY3ZAdGKMg8wkaVAI0LPADB0jxk/x8Roex9hl3wl96IL4mGZ7IS
TxJ0PREelZFygS99LgrgAHrBapgtYflw1O6rcUl7MDDNgYvVEG93LzX3FpKoZYhEvxvwfSnWfGDs
xf2w7FoCJhHMZDC3CbLh/KHbEpIOoHRFAjx73rL0WgqLHrMLVn3AZgg0OmunaafvlDNnRztxy01m
qnvNySQr7K7cDxnQ+4UjasiAtT386Fv3FdiLYe7FJgMB9C+ky4L4+YDg5Lznoy/FLNlJQp1XAc4k
wHBoVPnLt5TOoY7aHT+hkDgXvae711FME3uoYq92MpEX+rvSu0BTPvtpWhDG5JSOaLZsG3RfhfVO
xUrOyz+4hD8A5xgTnNX5npchSF962ocJWFAD9s2be8/7Icy66d0oBfqlSCpfsRVuiVL9fUZfjD5d
FbeazAD6yGxo+uDpJn0byKZkkZpZ2mejtFLnYJSYpAsWHMeE6hh+1ZQpVKcp2aCRXsdQhcoKAVXQ
kTsG7ZlvfNVNHaeQnZkxx1Sd+OvkNqBPnUJFFvtAtHhD9PBUzJCHpaz6epdVH824uv4AfNgiHry/
FuhDXz6Xd3CJJ0HP8pe7QZ9M7KdRG6gsR3X0RHQdW2LijOtS05quUF9FWYBbmDdEGA8MfZfUrbS5
Ewbo3b/hGNXLnMp8/PpAh6TOjgZ0dsRKEu7JbDkcsBhCLWOiM8i/8JviVGbizCFQRJemisIiwRGR
kxmr7Z0RM/kQ+8CIAoSf5sClX/xWP2HxjMt6YK1Q4JCE7P/SVHsrdAm4x8tTQREF1RPskbrN2sBb
O1CnWTAwY1ga6DyGdk+HzfwhksJe6C0PRhJK48EiTAiaHnefPg0mFsSczjpOubgjXbo+cpz45KSV
OVc9eOSxEox/mli7RM7u0ARMAXl18Eqos3cd2kduV5QRnGrfJsR3sasrJ5xY6KsOdndQu+KZ8wtg
KTuIF5DQOhsEM59j7Xg/ajLUpSPm1bhwYGMN1spw6/TW0jFzmNc+MBvmUMDACiVnie/nXI7PBEFw
Uy8M1He62bINvlfTNzfZjCxltXdL4IO6+fiQGwPYk8f3ldrTCcERgjvlpiHDXEOEv1/SRiPGp/5c
4xb0b6XQhS7qCHHm5PZe0SRhd5685VI46eMTP2LMjcKhve5veCsR2ck6S5Ve/5rTuZpE8qZ5GUxH
y1/U6ZSYWVOMKP/1/w+6Pxx4zrRuAqr2jYMqJsxxXA3d8+ezPoM7C3Ww6N5l5WOPJTqzUi7yGas1
a0d9XckNmQYKge6g3D0F5FE1eDtyjB9+9doSmq088fX7hA2FkMeSOXN763fE1ufm1KaJT94O5sPb
DWyyLpaFGmOgfnz0Kq62Fm4ppUZBqyWaOeOAEMdtzbtwzcDKT6bZK0lUpKwktFNjQk6wh6qtO40K
UVYJJjNEqznMF1/HIdblA0mJEUOqeWpQznti2ha2qas3G9Q+M2oQAydoAjgonx12BalMTEheVwx3
KkATmByFak/q1GRCYxWwepIwUVSL5OpM+hqtAmsU8q5RRHTgiJYujjv32zSL61uboWftuM6K8wGG
YvWHhiw9+j1lixYRlrcDcHyA8Fq4+IvS52/S5qM4Dt4xJ0UIRCSWj10vOvcgqeT7cDXQmDII93cF
LT0gdDzY4rmiEeCvGzIQu60ZmlK76ti4DB6sWPnsMEXT6SDR5y+Ee+mu3NkYo6uOsY/0zhmPm7eq
UarJalR5601pPDcIqSzmGSrjDV1ouQq5ruV12WJfVNAqBmE2bO3LN92J09cGKnUxii4FnYvatM8s
pAPaUAotVsXqtsNw6xVLwGGXuTDm+ZJFrwWK/dP1ZvJTxFPRCBQhduM7Hn5dP5t+N9OAnrLuswNP
nhaLvNqCP3Jkr9yM/4UOUuLklYJT9WTEAOxRSjW6tT6oZafiT5KMsqbJzOQanewMWO63L0eQU6J/
/xgxjcR3sjpKRRKe58c5Q3RyZHEcvxvYKf8wc1yM1mrD5ndjzq1rbhQa8Kp4uaDxnjsu5cYONm5b
83vK30wYgzOn/gGYPN5Q43f0eLEIIZCndZkPAegJTCrhQWpF1V5momEajMUHVRQEoePlc0NfRD7i
OtIENW2NlGmG71ci2ePtfPq4+8ih8Ou7vl4unoAGzn8waq3zJTs7eH183u5NsQxwSoRuz+Qycs8+
ZdNHrzhQn2dWTatpyk1KVANCm+nPAomrtaTUNt+ka4uveWULIDeQt/e5Y38MVMpt2yYxvZRRtNJB
sZDz9R8pvwgfixdjKUy+mAiauSGfJYhI5TvXqdPa6IfYb7lrSqZGoHD3BzRrgCkQ6cLOiU3/ePS1
9Uj8ULmjeJ5/7dPHemdNszGBeWO2U2AHnZKvEL25sFlI34TSocVQPZuwg2UZOgyHMCPZbkNkSJ68
swbPUG6w/kAcO3JXr7+OxSr4ObmvTdA3CwFdeiu3ulzHlKF03RZGz/CL+8fMlxBDoqLJTYEWF2G+
NcKVNqZEOfyAb4AQ33cbMTR9cy8CXXKSIHCFsBwAYWs3r8ckBoRD7UAZCuTpqQOUPpYSRp9DVlxb
Nikt4e8+vUcltchiR5BV6DJnmSfdfI+75mq03Na5u+1mn/FHTyFWgD9o/RB0d/m+B+brMDKD03sN
8YDVAme6xOMQjqTyc4HBD79Mi3E9N6ZnVfZId4I3JfvUUHwjUmUvfYeJDOcTnSkkcd6xO3P7UgQB
0+hOaPfukjDJMmVEedBLSFvT1zeLsBHcsIL39ex5K0xNg9i96vNZsJh+xsEz7kmiOU8aWGVxB1kr
7Wpl8aUDOZeMkPYGPcWl/Qtk2k7sU+XSv9xMkzzD86i2K0IJd4jdxf9CiVXCUH3dR+fxsRqZKBoW
lrXL1r+agICQhFLd6t7SgC0hr4uyuRBSFU9BfO64GLTJP+hrYQYzypOR7ymPbngX9jjoEpvcYSU4
rrma0eRIR/3qRs+efWmVgui+Hp23rW+lTjIq4JpC3X7VHOJUxyuBx99eusO+BGUkUm+I2e2uXw8O
ldtAlboCWO6hSCXVlAwFI6IhBLy3Qk4xL7M+37e9O1k/J08nH9LxUVPLk2JxEO0pHFW7UDoiWP+R
vdBpvcMKklTaTveJDqGM+p6J+qDKbt/58KBl28xT+ZhmQGlnxjaLLRgt1400bLCJrnnwQJTtAlSV
RosIoq8AsVH5qjQW1XifJImBG4pNfSPAnCpO8Zy8x1/GW7l6TRs7IYazy3Ida5EwEZOfPGdc8MWV
Nfu+nJz+Z7fh1Kl0q4N7PLmRso8Mu8W3KYVLHU2eVQ/hnK0yI/Af4NhPzz8ReTjX0AAhYs9rNbpk
F6kfZSb9Z1MFYo5ZlDnQPQhVq3V6L7OFxi6ZewzkB3PHmNMwlooN7YMVlFPs6PsCrExgxdixvxEI
pdrmomQ8z4ug23jIOE/WHgJUGx3PEGrjCqr9uk9vBxvq4s4lj2IlcaDPvVK3J/ErKduxXwxjR0GW
hgB2pvVwZDT7dqka1gnurIMvWdn6XxZG74GUctqtkxfMZXva+DcA96m9kYZDYr8WsbWRXvXCpsdW
un1VQjbYHVhKfurG4snEWIdgjrjCLIP+TdhmFKyHotguwu+ZQZsT+dXKN5TjgHr93zTDhU1U1CkE
fezLK62OW1aC62Tqenm6hm2RRGhSr1yAODcesPeMoCrRdx0uTZHVUGmpnwtb8skp0uldPD65JOng
SHK1FyP6I2OrXgtZESksDSnZtOt3smA++dADE/BCyROs/otHP9c5QwB+ZVltd5NcZqugTsuF57Nw
sOtwqQoHo5mWW0OEV4+3JRbgN/iED0fJN0z9CYLPauFrir4+wJnMkVod9YFSXqSBOzoD0hePCI6P
/pZ2srCk9bQE+RiHKUN5mLXaxgSPD1Z3ZBjJu8HvWnIBaIgLO+FDw6xsg3GDH19m4F0E7j6nM3Um
al4+DxJpkZEfDCrpnnqsocKSYa/Etdvg4ZRJOU07AlWEAc2xW17gHbfVfckHoQJ6DIUnQlHtBsnG
os4xIWTVKhvSFDoZYzGD04C/GfWS0YauPw8z/LYpPNz+/7un/z4q2nmjfSFVSEe6/YnW4MsGSVdj
9VBtAuC5ryBiFoqOseR2lPQtg0D9zXDlD03OKRM6LM7Q+CGO0C4XWd0fmhRWY5GpYf0xPSvCXAVf
rSoLbgsPtPhi7RWPD3+4odyUtb0VdLBdOsZMjZycP24TcTKw3Ls2Oq2Dn7yqIJ1VWnBHBtEfhcpw
bPsm2Dt0DNNFsokIr9OopzD2b2I+PQS0AWcj3ag/y1zOQoayi6hsKON7AEoRuqtGAPEQ7SLmV4wW
Fstu/OHwttjZeqv8Fd+fOe9YVtM1HGiabRP/3CRmRr9Jhzg8TrMHi1Qr7JcQtihAAZFooxqtLxA6
gCNS6tKHr2EOgyNd9l83EBQk2X32XXlVC8VOo9mTS5ogCY7Lm56p3vrXAtnhp7L/FjySLqUbgB4Q
ek8ubOUmqQuMS2JYJE5Wrot8c43C+48d2K/7OMblYBGE4+35hcqQRaZquZUCSDUgbFyGHyh6L9xw
iX8dahTknZQXsZosGG0QPuSyC06blxjoZ3usiYvpWsC9MeU1g7HHULZ4gVDQrLbwTBgH2nHdk2Gq
ya+Ln/ChsgSPvDa6XAVs34JOQzGd/UyRrXRuY2nmM+PdqDAivr2ehkoSpplpREPemrvWyChH4a2G
OgBMNY1GrbahBkUMcVDMesgS6Fx1havxdArId+yCDmFKWdE/zOREr9YR8YhX+6q1R0MLQ5qdkrm5
aDa3Q/7MabO1y3ye7O8oH9uqejWxLg6wYUoWhRzUJh7PwDB47g+wtzCWaPKMXVsYIDB4OpLFTtlZ
mC3SAqovNAy4snQqqPL96Df2y7bqkzR3Ab7R2Z++1bwwTA2OJzTuxGFKqmVX9/BB6Zdc5IOOd0tl
gD6VR1Q+CIOExQ7+H4Qa7yBBfD68d0sIcEYcNVHd1zmDoyUYn+cqh51isuGV1fpbnHKOBF4ajV+k
SE+I8Ay+fRjAIfI31BvVBa/EmSWuBCd7IHOqy+BksuZ/OmLtEhu2jgmoNKabioAREutY28q4Hn18
ANIX2Sr3pdmCqh+PDEHxymkahU+HGMzu0sKW8OMHNo/P+vtt13I6r7a4U8SQmy0/sybLXe8LK5H8
A/d5xS0RRiDxhwMGjcsixcpK8nPwXGrz4XvfWeF1lxu389aycLu0+OFOG1YdY1mFh69fnZvSWhiF
s8nfZM9L8MAlw+dmSkRihU/xu+9efinpbbj2U12B6Whk3TmEaLhIKMaRKBYYx9vpUG5xsBBZ7x6n
CbEfLhrFlcjJiSug+W4Fl2z+uBF3lfkh9uZfdk7G8U6Lb4ITJ1D9s/E2ZBq+FoXoKib9cK9zF8Rw
/no2m0paKj1nx7KKKRvopwPC2apoivW7ltVQKgkUdAzrpEeiqE98fx3fofi3VYDRcoVdlbEs0a47
CyJc9e0APdqJie3HZCuNdY8HZgz1VTQg8pHjfHDmH5on9D/7oA+XL9RMiPYswCtdYfi86q5qYyyk
jsbGekDu1u9Drs1EnhgxIZN9LSipaqICD5rLCFhrXPkLubftVRlgR7E+jalXYNrgTa7X1OZgffxG
kZx2DmsXMK3ufD2DlrHitJ/kNEXgGJW2F0CVR8bAMkM9BBT8Y7gKnV+357E/Ptiam97GDPRwFn+Z
pdLzyGfkJVNtH0XfSfKLTedv8vJDTQnFt85q/aDVC5EWR+neDsSzMD29hOvYddALCyucpTvBk9QN
TSZMEIJkrGhDxORR7GmGfvP/2IDyS8HvTpzPhVn1seA0mm5N2WcvbIBhs7gJP7RdLJIx7m0bYoM4
Ca1u1Y/Vh7LZC7Fcm/oRCVI5rO4vIm/m6WLf69/zmwqzcRI/rKrILtat2V4egK3nDSvQ8X8jN+D4
F0vgYPzr6nRKLe8isiyqfj1Qh1g5ZCXyHc/WwFixG0w0JIAiZQYN15rOipOcI7Et+nHMS7X4Pj5d
GJcNR7NnNUDKGn8GYxXljGOmtzr3S4m6tsYn1ebW7ZiF2MrkhQ7EgcUOjtQRnjB7pAYpOuUgRpLo
D7eOAa5/gquUeD39ds19WoYeYaMkVvTaHNEO5xXaFvxXys8oMRwL6u8qu/jIsvOzQPx9EdwvJbJm
BvJdVqtAMva6XPxfeIkcbJljJhOk3gfpMfAMWPHdGwyFuAs05sn/lHczm9C2IVUoKEaPswCuPZGY
Aiv9ep25X4nO4W8OrMhGVEUMF0V06i/B8g1AUvkTDgG3QJQV89KrW+q3kNLRJL75VZQGNFtcarJ2
aewn0MhKYROcFD3JC5jMZC1Nt4g7CpykMM058YYZJLH09E+Az0CigNlL1pCVvnVl2gQF1QOZHU44
9Mnbh1gaMb3J44M9xlq6Zyz7H0UMx4gcCJ5EuqD+EGGVua1bqi1sLwrWxphg8fapIWMIANiaQyKp
ig7QczFenWI0fSCanHlX9FO0Sre+ucqhLEkSWX3bgf8XL2mr1VCfE4dJzM43Dqd6d1l8+kLWfz+2
h0hJXu/DO9YBFaoIkYl9aVAZzeONlUBIHAAiMhISE8jN9GrgKjJwEZHSzIUaF0HdF9h072mbDO0R
URJXwYSq0O4YMS4jo+/gbK1MG5QcM7efEmSdBQQSBrzn7FQVwaOt8AV5QCZO+f/C9Mu9Vo/F+sAR
e1gGjFWeYaoSDGkpTY+KCCIVW1GogpSRu4VZ8J3W64Y2rIYxDkv/KdsChAXbRm+WUXZX6iS+zzKb
eb8NFMxSWRRVdgPogAS+jgfevbI7JyBxIdL3wJzF8Q4HquQD8ruwQHZpT5wboG6v578XKW8i6IwT
fSXI5c3MOjzZxbptepnSRqQNlU39oA1uc+3eM4/lL+iIUJJslV0M5oGyG9StiQMgvVEltl7Ux65n
vbrR7XEcVFMHRmh6oukm7Py3wb7idI7hilNhKA1ub3MHbIRdD4W/N0PyR+njWaaUWDmOtUySBI/J
z0NVleAi2x+bF4DFTuMIl13uy0miTFEBIw48uzGED+tt62NXuTMbqA6CAKOuGwqYa+/7yLOAwHeN
B5WtJ4zZL7Xawuc86lLQbJZK5VOGoZeDyamRME9uCAyHWUOwW1UR0/XtKLKaIO+bihf8XzjS6SO+
2R1FmRQr4iup7bQxNLodwrxfVbJAaQOWFWvFHsl1BQrD3fqtGeDQIgd2tiB2C7EBbg3zhOlyy1fV
bT2BhcKy/QnQntgHzMWiqrWjlfcVyttGVsIlIfmYkLrRBtDJSdZ1zXMHGVXKwTbIcr3ch24UDNnP
5LPebsIB6+K02AgqGKBYVXkjHx6DBU0cgUXNb8zSMREEaFfMUubguKIZY/Bwx0ELVhGf5P6bHht6
VmvBzcIoq7Gl4rXRI0/tYNaVKcEhDhQ+NVolj4C06yrGib6+Rx6ri/raagDMXQTFj6C1zx6PiFzf
yWeRb+eS+QDbKYfCXZCSHU7lC1mgN9cZHf0tQTxVR8e0vStrZ4WfFfa8lvEJaIIyFMFzUuvTiVSx
5fFwe0riDO7rj4LYF959kTC6EKTh/at0+hC3qeul6U9xIiDNVc6S52HbFRsx2hbPGh5ffO6o3V2i
qYVqfYozQH3bV73762VirHAA/hEJd4PIlJfIxbOLFyFE88tpoXxhGCKTGIdSI9L4Q1WWCNj7oIxf
USxEgiaFHvYwAguNz1Fp5aiaugl6b6iHoNp244ImUfREkSZRGvB+yCwOAhsV8mgRFbKj0CDc9JNn
n4kpDpaoehP/l/J2b/E4oMm1LIjX3YMjBAJMOsQdDBJjWtBrva2KHFXW7tH3a7pCErjWM8dFWx3C
cMKpqiNbvjh5m0sqhVxTN5dYpZPrXIlf5SWcLUl2wk62Y/P0eufuQqfvbnXGM6Und4G0GkJRpC8T
hvgOnONskogu3hEK3ZRUhArGa6pRWX25bk0HYelsylRW8gns/rKEPQUOVRt2YdaCdwTANeZfC/Pm
ehmyD4HGrZtpTmq7GYkoQXjIzCdSxxFC/1NkfwXiHHIc0bIScXdZRd9Id+m0zFjoE9l5MCHIJRRF
zhndNnalk2km3ABZN0JPIJtQrLb0T7syhYRFCMj9a6DKvnciQ7GLxmOcX7Lx3M8QfECOG6Ee8WOL
4dlC58SswPlPJ3Yx4Sljs88R6SVR4+EwQofU5NV6zMrliCqUiSe3fa4SJD0grA4UgaepfrUVRbQl
tIXpOuI3/7aRTvAKVjfdDJw5SWF7lzmDzyNsg4LaQUJaskM7ud85iqjxxv7F0BpwtEgL7cek4MTe
FLaJQwiDOMetFhsfTJhOXDkYcxfdQluN8sr3kcoHpr8x6Q2ADWiGltZpHwbEiWe+44V82EKbvLlT
TmHg3xHsnDWrtgUtkUa+BSTIZWyG2qSrw3G0ZoXkJLIzDRBfU6fORWs11nZ+phaZN8wpEMRd1ZUG
vo1tbpqK71LV6A0UoLYzlxR5E4V3YoruGgzugDwi+Q09Jpz0+Iyhmel3NcEhr3xqmGtC7PyZriWF
vNiarYyzKQWYd2OoDEWIjkY3u8nASWbSj5YnMnSfJJio1TAA0L/r3/BSJhLLboLGS9YxxkAepGz0
UMsq+D0ylMVK+Fq5Taiz/pYO6dX59Jj0gz9MZm9h7XD4Kx/SeVfpqfz9k21+I3B4FnWAh8C0uMaP
OkiwKVRe7MEDzY9SSlqO+fOProo4d2GJd+wqG3Wr0QCge+5l83cbCUnBEbDONQPOM+nqkPwoP7Rs
1SKdjSJA/hOBwQ4qIERJ9hQ9kVI0I8XLq6JmUkNZ14YE/zuCJqP+TtBNb4evMuVxzHDSK/wcPumF
4JzeJLSq1by/y+PBxMuh8WZM8R35ANawBUVU+r9x8oGoA54zQr2HCr+J5wuXVPeV4IqXmfGtVJsY
XlsflwNFCfyNe0zV/p4J6fQBcpdgbKYobjDHsArdbqz32LbLgBNHbOCiEtMTkACR5WYNmw5sknbF
IBshhoNyIAm+4IL6c2W84GtdiAVN3Dax15xVWSyvao+SE2JYxZ2fWyM5z9aYLJZ41icImQiQ+SmQ
JGRpc1k4RwmRGe3fl9hgqEXz7Dzemsu+ZOPfFp2vX4Oh2ayC/oLqBrBg7iJ3W4oB7cYZ0t/YMbSz
EfqjGtdHGbFVOPv1jqJp3+B3OvkLuKnJ8J7RYYPTTtVTl772yv01ZTmBjbSyyPOgtyqdocoF0SaR
Nvutzb/mSei8OQLJ/Zya7gOy6l96FWmbKCLbkpjFmMaqd0NzyHKmGbivefyBVAirtzuwmtOM4et1
i8hna3Fi7Yq6T+M4YpePUzUaPukTBJDsZFXpDa6L7zSXr/7NiVA9YJUnxE0dZf7KCprgp4egzQai
5HRzofveRq2dkNQXgwUZKeyWTafOhUeKOUZmjfRnUbBBFk7yXOOHAs4aDJRsjR9mIDZRF1UK979M
6qurchCsTvmSqcha6Nb3m16YmB3CW+dl3rxR8pkPV/LX707HCtUcfncjeNTe4NT+J1G7TmwrvmkM
w3Tse3lazmC5J8pbh1t7cizfFduLjfHeE48C0J46Kau7hVd7oxWvTu+NmeJ4iTwzomNIfZWd1aHV
icaJtinLACuDenDFq/lPnOcZ6PaWaMlcHvpjzPyJCZNVG72RV9oQYkCQwWt1up0TWxzjjda4C1jY
Z272EbIF+TFRdALl12tnAvzmMg1LIkyHOLhiaoDux65K2O/NZTcMELH4WYGarL9IbNtlyWdxH870
J2cZi9PiB6fRrP/FBl3Gxzf2vhIu30/kAyVkhLWhUqNcSG8j7g85xP8QxMScXUgqaWqX09lHSSD8
tJPnlrwZ0kR0ZaT1/OrRkkwp7Q7eFMS5JyUzfT3YAWnOZlhZuR2zZI+1rIQGA1kCTz4sWr0LLW+1
sB48MrFI2QBr4S5uerygl7UlIDs+RJ+g75oDgZ8vzjxyVsJXF/1lfDvhnCLIoaY7kTHK4NOUE84D
PbTwKXveb4AUIzJV/EVyMQnS/Em243EsJdhAQKjV2VvKzs3nwXYj0I1pk8olvEJhSifoZ2BbLnCA
okk5UgNbCCFEtJDtLRQ0z4z4wo2a4YQ/u47PITGeVhrKCYk99OOyEVjUOIe0loaB4nIws3urlpeX
O+FXZz/AEAv6ojjLkTmiZzQdMQ3pyMmzwdfnhC9KhbQrcyU3jN0jfpMHN+bmEeL3WDCxv30Oh0C0
gIZV3K3J8RwNgkuRg07zlBzzr82kFZCw1SvGUVK4PXhCPoKHHLM/2SN7E8FIwCFk0GZM09fpueMV
7p1vVNzya3gbaWKfu3hHTwwTIB7125ZdVsuCXZUcAkEVi/qJGPgu3pL5Que+4hQVp/MiB5tSxyrV
qbDJeG9VjI7HJYOB8Pp4QD4rwiATiISMDajIQn+lFv6398hQOGc5TKb0gY7oLy8hnjcOLSZ9VS0T
jSzaZkzPz2rN9Zt1vnHqNykFX/I2ljsoZ9tiNUep4FS91fRzPs+5iBn/O5w6YgEF+0ZjrLAYkvGN
wS8h7cz2XytIxPpCkdjbXzoowPjNh53xvG4OTYafIhS2YFzkRdyP+dnNy8pwTzQMdTgRaqBLJSL1
PNHxq2mUwKYHpsSmS5SrbfTZcIzi2vj6oodm/ke6dHcnoIFhl6qlRTk8qu0JCOAd876NuuwWHqMG
ZHrUM/wbWay+LscPx0Mg4n6PT0A80sQlXBg2BAGd0FnenB0kwzcvUJ2XRhZgzBPJ9q+fSTjVRInA
OCbjaox/o/e6O3LE01j7GgIkqIGDaiPRJd35Wg7vCRP/Bv4gwr87uH2C0KRAxX7w5g9sa2NtevCd
DBy8iuuMGT5etiGe0h5gxBVpSvC8L36EVwS2erwfaH3liMuH/QJT/uBu3wXZ5lxIX9/YLHkVDh/L
Jg3vsSz0aK9rWod2UIAOmzQD1ASpKP0XrYSlUBz2dddVvUOYncfXN1gmSodjFIJkn6gwfmdmvs/k
Ol486mHRsNnmL6bW6Dpt5atisPVUTmBfPRFl57Tx55flxAbx0q+zvjjWO5bdDdJDPd9oTVOMf5RU
R4H3P7si7Fml3ZRAR9RYX0uWPwfi2Rr352XFi8lOEDVCKe8fdbAi0+k6uHZK/38tzXk1iL40ielS
eQIPuVhhYQAwAK7Tuv/Q7xlBrcSNwQ7DdsMjXeWu5SYmHqclDcSeb5jzPG4yNVfsGuRz1HVoNgt6
YpptQBwj32vWP9sstD74vx0JGX9zwUrk9f83wFX/NRfRnmVJR5Y4cDt7oPcvZsHjbs4DdN7EzDkD
afSdXxfo6iHHXcd27xR2rlhapGLgavzuaaBJJGqVwBsOxvqF/YaHQkDyflmWvneHAivhM9UdHHg7
7M0t9ZfvitQUXY+crYWAhuRKew+uNeYLQW3TOrkxoNOGn0y7s8NHcfnFCdo1/29JcnqdIu8756s3
iDK/peIEKDv1SzLCqH9Z1w7R5A1IGcTV5Rl02wpurazb/MG4hQbgcXSN8wJePOh8HHux9X+rtenO
FsUv7VillVkJcC4QNKtHbYNIKEZzS9FhugElVXnX1iqSez3RUyYWR6u/QxsIf8rPDGb/7XAZXlm8
fTLH3ld3D5S8RQpzoLco6lJFnf7Wol6hj1r1/qWON9JbhWFetF4SXn2qMQaL4xvu9ht82NDkHgvz
GsWQo2UYvxrQKsBfDBpw9r1IKlUVegNuzm87Wv6MNMz+W9bXsl6mE1DtcBHdPgQtKUUDzWhVQWH1
m6YF8meEyDSN3Zcj/IjvkVLmUW1+ThgtvHcSW5A1NKueUW50pWtJ+BzSJF3ngLUrgNBDAFwtDTUs
PqIE56YpFEaDRQ9F+Y/9ILwud9TcgU5eyil7DndPijRnLwyfPrCRsG6L9AUNGOgr/1/ead2KiPH3
l0+vrV/mVE+XAy0nwEP3FQuYIyV9Cp8Qv9+9Y5G9r3w+4KFnDe2PR2Z36RO7EdJcljHbQ7b0X2j4
wQlZkP87VcBoPDBBdcGxJuFfe5phRlhD00WSUTeejM7ZodUEFD/N6B5+2vEcONqxQOqYcrU9L/rQ
u9GpBEPSj7u/Pif9JBJ1c4E8M3Hk19PUjobIZsAxapLnQMcREKFY+5tjhTnzC931t5AAeagcFd2Q
k2qNQCgxflF59bo7CXFCkh2RsB7hItupiCtSVRMrU9KjMVY4EaKI+bUh/lwA0S8PVwU4iMjFoo5r
RGyW6zKMjm0y259Vdj7wfLy0se95R4MNc41IirDgmFkvX1Kv3abQBEl1r+3MeqZl1kXlUbfeN2fj
ArYwvczzGEO213eK74rlcAC0/CqeBFV6h6Nfel8bxEE8Hv8dZNeUs5LD7ICmDvXyx4P/YVs3FoDF
2Aw8B1/kiaS/SJmThG1WfR9HIdypBgW7L02gaAGvXt2F+i1KIMoCRPpR1V5QDT5MHE5+S5VYYypu
9NmLcyUp/ue1rFUcryoFaftraAA0DGiXx75H6EcodH/4DFdBToA3F8VCcwvoOlD6N7RbDslpvMWS
sLJJcq+dlslk+gwVCVr77C985IgbtJE0XEPBklHwR7LpNMABJxudljAwMAJ5ukDLKb3aQqlTmz/a
8PPK0hL7Hhg0KHTrWphWT8YSdxQtY3mr04evXax1NRLfo4iyZ84mcXgbxFxlbyTrgR0NgXKZSNYF
brJsIECeONX6vHHie5g/9vIEJ6wtNLDzjnhCZljTv5ByHmJz039PM0dBzrhibIOZklcy+PbTPi7e
F0JLMfyqLgXpPva/h16vWvofvZGAtbSZe7O6uQUhroHYhQNiUScD6XGXWCpQqlI+BB4BJMI1seIg
5VgCpzijwZ9awpWWslf1PRdTM4jGenzjz1+kSYRM7oDIvyMsTVStoQbTdwA3OiaflJDYmUghxhn8
9E2u3fHt0uAC8aKEVM8gQsiyS91vp5TlMu+tfg89okXqjCOzJnE0LXMhdJzsTim405E5xBbfdeIY
c+M13vZKgUVP+tsypzmzmfGaYChn/3yArhzZJjzbMtMTQ2Ql/AYOKO45aHfqMhkJw5wEuoVU5O1r
3mVZzJ2dVk0cjpsw8KOFdbRt7RV+3zDbqOZVFunhUnfdZHaxTONJj+81BXUgeMNN765R2oHNTbMc
ewQHV9Oanb/OWJ00x63ixl5I0GDbgf8mkICvxpEZtSI7oZwHSHHdQG45WA6Or9/2ygRX44KMQTbp
4X47WtoSWVUIwUIe+jRDp2Rx3k9+qt0F2HP+A/N3FFi3WuuY1yG6KRz9y+mU3yuFt3thgE6V8srv
DgL3ndYFmqIT1JqWkdfmVgG1BhjZrh/eMkRLd6EL9BFsoxs15W7753XwFA/cZQ7LKfUJQNKdWtxR
kZQHLAoynQUaaggr+LUIjrv/3rr19Zwxssn0Q07iF8Lr/VNhpm63LtZzP2Ag7niW6sPdwthi4p94
jCfZurH4ROn6MdQmdJrqGsLP4hZF6bWbJnyhJC7VhwueB9h0XNBq8lsg3exSmlcfxeFeoc7NZH6f
d19V5ZEojL8+Tz2tJvlyKwsbYbQmPwLLD/dKCkECyF/jADgYCWy3zOizCPjsPhwicV+QIOuY5/NU
zjYzwRJdXfVo6r11zCSyn/vJbvsYOAgdaFB5bTdeAAIOugfVWIDmhTS9huq4jQPmtvgTV1TBYABV
fkBxcGl438tHqtxQnWFxpfq7/pKaEF2sbrjD5d2pXnLMKAxDCHMpWlp2SyT0Uz1FGUHGcyE8MfqG
S+CpUy9/ec6NmQXvymgR7TAyPYfwz8QAX2+sufOa5GIFjGNsR8oTbCaSqeiO/dkGtgzheUuP39YY
XD3WJ3JbtpjLgMiLUxfrF1C6TLjRSsMPlkZD9SyCI5KwpYaoRouHhMu9W31izvR/ZKeIFXgKxBuf
z6jSDwWHZkJ95j77rLOBxzBO4BU1jz1XhXGS+v47ZQFhf2xO5zuXBHm4tdjXyUHmfJ7eSdHaC7ri
JoDZr4a1+880Ij5Z8AnHEiqF7sz6pbH5PW6aNLnpo8ef7xcD3J67MJxJ+6Y8LT3+1hSsN3agUc84
bd0lN61Jj1chEQAwE6t4M9RsyOUt9sh1ndPU5Lqc22nV044Nu7Nzds4LBQ0E/OG/i9FSm/vNExeW
HX16bqIIP6JhNA8OEqAr26XSuZMLhPPRtSXlK37IX2TbnMZbFGxfOP/fFEUCRaRKL675/Fc0s4oi
SxVUCRJuuq37UeepZ9SkrqQkhzZg9pGEHsRlAKiWSA8vrU9vNUiwXct82jyeBi0JBwwDLRCRRltF
Py9JwnhamSCujOr+yHLBqgIWsLPnPoYVOyl6d8kqR2+aCe8JCGJcVruMZl35ZGy/kQTjDXRtidkv
U7TyizBZEuPJMZOqWj1yh58yM/bPahvhVCxnryDRKaqfLAPYWeyRU/S4n7m/i33bG7AOWn1M/ne2
4k0raMc+kIt9kWDKwLJSb09iI8ymApYF8kfO63UJpN7g3lEJVqKSy6mOnwETuS7C4n/ge1n8bLjw
ScrLxX1h/JI7PdYcEFJZPRUipL3SMiI1I8VrpD6iM/xSfaknnSgP5tqW/6FrT2cj5C2fWfXZVHwj
BZu9fGE1nnIN/Ul6daCgoxtaO7yrDVBBf6J5tNsj5R28J0Qf8TzqBLDEaA0kIJw3kXGcKa7UmVYr
UgiqSLJrThoUrOgoE//mFIXtaAwgNSI3G50HwtpG8x14A5ohvet1Yw9dsRoGJ09Hb1HxGO9rTiE0
rttlJKoALq0Vqxd6QX9yum0SYjFRFywctLWsHlF4BZLU2p/wL6lgmtlf4fK8veg2ofajQFJr8v1v
ebbBVRFYfSWboAYQV9KCpYVeZowhWKsq3W+ZyOl2iLgzpKUiXQWKYOpU4F4fjmyPMIP2tw7unrtL
FPTNkj49ZgRC1wlZMd1JTvuppLdnSPtr6JlMyGQTcT5Q2X6zaenbk6hGB3vamFMyjwiQJt8QDq/M
XfUVEPMp98K7sngx0p5DZZ9txTw0lC0G9RVEkKdkeVH9/GL07aq066BdYsyVCqU+clKKDD0YZoiN
XQ97lyg4KrEQSjOhB2yHKSyy2VW2Wm7ESWj49Sz+eQiaeGoR5n15z1Yov5OUQn6rguqtqNIteJUT
657oQs/ddvXQXlOcYfaZ1B1COwHMHt5JJslbHdCqruEmPxhax3s1b9JU97DZetKJStC/AA8QJZEt
5EEZFADidiOeZ5+xoNjOxgD0fBclT/nL9y/dHMH64o+FQWYlNP+lkP63UBB/dUatXoz8SaP0BIrr
wPvdvl6jP2aWKOfCE2Tv5yC9knUQOfRbGL7tLioj3SNjQtycQySdiFK0BfEsODAxFnS5Rf/d0sOG
PknNsh61kqdl2FLbJKhWF6x+Lxppge12ZjE1SUBDYYHhYPbZZGVNDw5E71DdpyErIyNiFivNs4K9
LaRG8m/1N12GbOkq7/lRkZeye87EFHZ9bTD5yM8rjHjNbegYw2K6CVr5zjMOSDgSWpuScjq1jE1j
J1TJECFH09TmkpHwZBnhsaQMW39OG0Jjz4chJdVhRq9dLbJ0Fv4PgBDKaZGxurhvsvPmVcrw2cw1
WxrB2HToVszWgm/w+FsHvxU8377X/iD52e04hcfh0QEvdHiUfgxA89BHG2Id5skBkWY5j1o5n+pS
VPoN72W3iLcW1iIjpZ1SJWq0u4vjd8pPs58sk+BwrV6kr60iy8l23IqCaOqEc4zBo9U83Cw7HLqm
/xBdjaniRGDIxSXKde3cMEMaGgl1iqLWu1pkIS50t1ADTa7E7e0DudcXDZLCjHO+YvtXIP0Igk6U
wa9uw50LZa8OCf2ZO8pjiUz2YLach6Un5CnzmeCBpAsxvqjYhrmh8AwKCwKOtEMEQ50Utu4DO5fl
YbEbnXYobGMWBUfTdjuxemwWwfusnThXNWkl381rpO6VCLUSmpO0a74A2ryFKpWnjHKzijnCYipF
E8tKCzHrjAVmtA7y15O869qrBPeqg7DzQLw82Bu6bTlrSUCoGkY1uFIRIFE1/2wyFFfkNN0kTq52
iulxqIRE9+cIy/vBoBtpBVfrTWYShqLMv+hFR/JUSLyHwdNkKMZ0M78DCezNeVgSYIYGlzubuW1n
3MIXzrqlDCPoWzRq7RScQpH6sVvBci1OApGlxH4wyYBPzkKEcv/8nOFpzzL7DGnFCw8hmh5Za4da
Q0iBzH09yELddU7T6gTOlKTeP64DOLEUXNx4l39h043DVB5adDq44xOGzS3DevKkP36MPC8cXlAl
Sr633GOdcQjo9rAJCOXJlEcMPKursk0vrCSE6seNCeNPEn7ow02DSsLT15D74YRunswWzFFeksnl
BN3rLerR3ihc2qrvxQ8ZSWNwMZhjVWnrvNimG97sc328lKR0dwBJ3fuvhi0l8fxj1KnnvenKR2KA
2DPe0/CbqE3RLg5MgIJ+ryok/qpYionARFIQFy+OFy9KF+2bfV7QtXeDtdG4GAaCPG2bnMaPTlxo
K2S72UL0lZq3kMybwSihxEo62X5yguie4ID7kpTcXlE/IoUFMJLV1/glDehr9JMEuaBTzOp6N756
9pJ+3io+iG7Te4S+6sNyKFdEQtObv0VSSyv85ViUL6S2IazasAkwPrdDCyvoOYbZXHQdWgBopLLr
1DJ66+dJy/bGKzVRaO/3QCggELsqIJ225kqOWvfNWAlfARWxBvQ9c8gKE7weS2GqkF05AVZrrVgj
sjVC0yLMwy1a7Rz+6RTU/44dEcTjbiZTK2RcHx2XIMUXASgjxUD73VdGDEiwqfcEKZY+fT9YJySD
R6li5T8ULiy1Y0I41UpXDoPvpOSQLuRCckP6rbOa9Re7MMcI5XFgJ26lWdMDFg6bmBpBaX3abNGM
u1oaH+jubTQBealndQIW+CJNHIoUJxnuCZnleL6rlwH7THTzRXGhXH5xeRsKdaMcZlSsXO+hPgmf
aaTA4CQOw7OMbWILT4WjLhgiXZesKLqTdhkB2at/1nNvaB+zF2w2rEZgNqdaH2AF0NBSsUefq1zb
z31NqXrJDslvFybWtpkcvkoAQuz8VNaXq940gzpxmgt+IqPa5uLeyw6TTwWJXQoleS9J5+Y2ONtK
Hcx2kGUBhBQ1NN2bT9x349KS9A/517dQQ0xwzUgoYJ8JmJTkHs3fQWFNEF3YU9nrJU9z4MMli5GD
qVCVaRUw1NgtrRYyNGwXxKRWtzDEghL2MH7b8SFjMvUrLxmbt/ojJ4avQXM/oXVx6NerrN4nJT3U
m/569a4sUNj4OFJ+nfGXQWBdziuAPR98Y8Z0IqzwwXCgQp5CVIuHTJ+zm9ulyOutbPVwpH4gJhaf
gDJ53IAT152YmSepXqx8yxjlsBeGODDqC92qbkIqQ0s3tfLMD4/nM4mQa6bptTDsMaLHwjYbmDE/
Sx+Rtvlkd1xl+Y3quObZEfl5bf8tSTYn+PCZHtAP2VTpkaUvEjfOwEgqIJmc3LsAFO/3AuiBS4Ma
ZyjnNahhDsgDEGV9m/Ux04PMJmmeQP41csi968y/WybL0UTWp6Oup+FcmjCVRl7TKNdPfsNA9ZS1
tZBtDG1E+xFRKDZ/aJORPRoi9RuIVAusnoIweUz+9f0ydOE35QsMnBFtOT5rBDEti/zkjVdOXtYX
lCkwAl+0nIsDvWtE+mCQGWff8IjXlit51ssXRpJQRkW0taWh31fiG5UJZxZSmNFP2LDECMjM8u6u
wtnm090pxdc8X1NNWTsm2rnQfRCTrrplaAphnNeHikJV45CnFos89sxdCuO5x0caKPnHVH06iEa6
/X/IcMpMJ4/SlIAXJKHQD9vu49xjjMPWErh2nZAWk1p8BzPs7YqsKAeIAF6Lxpt1enlhY7OlNX8p
FkjUK+ZfjC8pfdPrfZnyk6jW4iZoqhgYjUyNIBzf2aio1ad6XDarDEEXodiujfEOArWSLNh3CTJT
De3gwyWRUXYDQSRaCmD6Lnu4s0oMr8FZL7CqUyhIb1j+T8nBteedpGWzYlIQttqCX3WYh6wYV9cx
b0k3bHWDiGMMVI4vpP2Ion3pqTQowvmp3GXBLAS4mnts+ZV+t9nrDs4F0x8bV20ri7kzftQtZyV2
QFDx3ylFp/r4Xo3YWUOjrfy9Hi/2Tf7ubT3hotQ0oIZcydyOFRCQMOMGxb3BZz+8b+qFQXw1Y6Sj
ppLP/oPyYyGCw+q6C1sRHeNcNHOxfAmL+7Wt+FECSNHokE+cFLjl70XhmAUabLaUAFl6Atvbid+s
n1mXDq6ELvImnDbcu2XCIH6COSOxcMvutecl2n713B8cAp4Yv4RsrQ1Imf3PK55YuxcVTyGHzJSv
P1JF+eBl/4MSY2Ngdrh8a+baVNogERq47MClFJBIF0xC5uQVpwH546pF/5WvB3Jax7nJHd8Enb12
HviWLJeG/Sa2s8+X0tvXy1351TYZ/OtNr/qYLCO6WpRTUjI9DV0ICJZnA+lU514cWdB6HHjEE2MV
xZNSCiFEQp/jxm2abK4crczLQRPqtRaQ8UsddhkPOsUVunAc3i3lOSUrvlHcAeaieMEjC36HDEvm
2M2csJJ0xhj+WXlSZZtk1FN9es6CPQJH+SDqxfIXSE3z75f7RybtxoQE/ho5IqsXqeDirVWJAKpL
`protect end_protected

