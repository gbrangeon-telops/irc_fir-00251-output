

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qCd+mYB+5ZYTiHGVPy4TJGVU+1xhFKOwciEzku8LKPbRfJOghBFppfv5cFbq1oB+i1BSYIHhjBHe
eBlHNZ1Z7Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U42W2uzowOkwk+UQGZB3li5Wu+ZZMdyVhWtZ56tkrk6iW89qDlhJBbms676mTh2iLt20rMAIN2QI
nrgBsluV4yEsobcfFOejzkUO7m425YrH0cSwookeI2lEA6QsTIAcBHaB/5shcOjOwrXurevqKKI1
D75XL20Mu1iceA3triU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Nn+1VEi9KmQsJsZi+aKtcGLlFmSquXhfukwVLZNoicIm0aMjF4ddZCMvsg6rFcVwB/qfiEbWhQta
pSDRK+xrjxFlcTBesAmRjUBiW3/wICtAFebLqkLpSTW2uzkYDkrpfNE5IjiANv3SGir2AFafH3k0
HfjDFe0WiziIlRflhOF0bV/y0LPPvcdBpjP9raAJY0w7hoeg+e9PIbHp/PMxlJRxsOwGTLR7XK0o
em6r0lXpVib2l0JQy4vnsZ8th3GiX0bt/UuR0caCktJupeOBsRztdB3gkPhiKQLg0696Wa/3XX9l
8h+H5UXqQy9EN5D0ZK0mIS8tAdwDRw6O0hbAiA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2LRSSTguNLx2WvUvcdH5BTmA+6dHxBZj3mWZxmBysCd90ElOkYpPTP1RgJPbqjpN9tofDDFDarkq
+qbG4SV9hnaX8iB79Zk1+LwdXefyq97462WHnxaG3I/Bff3hJd5X0rJVBnbVgHIqHzt/V8g0jC8o
7m7eoWRXpC5NpNek3W8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MM8YGg7IvNumb+k802doh47T9OSqo/qSgWEpWTgYva1SqSP4phIChk0ewsR6o7XTxZAD05syyzDH
Qfzl5t+Blxw1Jl5F2WrihR2G4uVbXDgvFSouhPopV4gzzwlFtcYs8jnovuVf94AiRDosYHN8WPZW
68LlNRF7Ti2drGO+AuUCHhYE6L1qXzzHwb4c9QJYmemT5/44a67UOyG5CnTiIpfQTpVHSTGdVMr6
z6vPgkB/8JeX7+R+UD1AQWqiV2w63od+aHRP7gt7KRL+kgJ6qCMGiaLr3Wj2C9mfPy61ebJocomY
5wy3s56g63xqQQnm665jsZbjTUelVxQyQI2r1g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9984)
`protect data_block
ipFz3hj4v2obBB41xC93eM2GsQIIGyVIOXEBfjxePLqcfxbAx5Ut8tC7zfb6KIn8Q+rhsNwO/z/i
lKHJcke9TMiYFUNJMsjYhMZMmgGUQ5ig62XfxnfL9kbR+U63Z4BL7LdklOeXqnkcJpPMxaAqayE5
B6mve9jyPgCMjg4w9LXlyW3/cpax2m5QUNfpW5UE77JefSRFoYQ7bxrMqbAwGSscjJ9h14SUBrx4
wJqjDU+PO09b4s9gQavQ7Qc2b/MJa/e/LCAMANLuAs2EzFBrhGVcVvYksrEWqC+e8eUuU0DG/ouk
8xVeiCfHpxU1VrtuTenFIAlteuip8aNL4mH6P39/O4QJEUnhLLStXFsF55LNlMoz3iKSB9k+zs3x
U4fjHF3MJI/Im+lpyz0l4vH4VcBvIA5WN4QWzmMZBYgU38wMfan6qDuYyAM/83CGRqAnGDrTz0nF
3Vv41wJsdHnBxcRzYok8fQZxW4GB49ERBrkumGntO65roua7dFueJzr7T7Vve336oPWiEnua3TCf
XjM/1XEkLdfde7ZTFD8Wq0sHMQDXDWfGMtL14Xp/2QUT0P2A/e5eifZv0ZS3FWX7u/swICJ2crIk
UZxL2ZVSHjzQwTBF3HiqrExoRGQMPf33E2nr+6vnvoK7UoBgQGPvA23qDKHh0j6prWfd1sMhg7gv
rgYL6Jl5NKVbL1KsgsRL1k/5lSdt5765OMkmzLOADWDOx6oacKJqGaEDot9ahUT7S0J9kPPq1Eni
wWJ98ub8Tbw4bmC0SyXbWxtj62K3+wMLYRJ4yoDEigt09xRaxTbG/lrc4HCVVvjJ+628Idd15kNB
guvkAMw/IGK6gxOim15UVPb3+hQnK8xijYdvSq1jkUqf4CShiIQaPIkUB4npA9E/mKm3ctBm+4mr
vj/Gu2EnVsVRYBc041hyinX0ikMnBFZvQ9FGb99z6/M8tHOHCqqRZLmkDhxRBEFgi9zXQs3GKqw+
BL9jwcqhU5vhX6n1R1UXXDF5nxX0RI+lYxnTtcc0rf9MUaYQFkv3zPxd0aGV3yiZJAWILVr7SzlQ
BfcohVqDVBD16EySQyoz4PHwS6ld2SQcGUKkfr+wwZJybWZZCrzmWBcmOgdWYqSenWZlyRfsnASV
c2ZbSJEBJTrLcvAS3hU5lqPRAIl9howxaQ2sz9TNcv2rlMni8dreEQyHDbxz0KvmzfiaVGmsUZsP
7w3S2OySc4r9nid4BE3wV6JdFMJeKKqbtN4b5W5sGCzhbZFNtlHWz6p4amYsZvOKUb/k9MIAMlh2
l70bflr1/knjrE49P9FLTSBLYNsMONbeJBBuGhQiKtvU/bNQUNCw0rdsRzqABSDqEqIuSLbN472S
ONx9NvnmrPDmBk6XkSMzJN84HAIyVR0eQTHa/JaRjic6M/wY4CciIvVaaBZn3EayozFUBXlA7Idn
TRTGmW2kTo4j14vCESVK0aD4AVh+JaiwQRmcVYBbf63/sZ4adgOo+t/0iYQAeUifFkRAVPOltznC
G1uBvn5iZnHe8i+RzgcKFRRWIuiu3zYt+4f1iSZwapQd8AEgF2KB4xqysnfCzNstHQj/4v5xPY5l
Pkh59RYM2dVzoE0qL+ySExsx3pIdR4yKrucEKaucdrFHLzoFErMZLs5Q7ogKeWAOtCLEDF8tP34Y
L487ZlgqDz2cQVgtcUEZ54WO97QHOPRpBeANKVs7c5xX2pTNvNgnq5UpFaki7sE1k6eFUvlK7Sj3
thypgZ+QEYySaER0q8tDk5Uufx+5ORnwohiayJLB8K/ZTgnz74l5exVhzHtKnTCzzkPHYZXsnt1B
nCgCz35j6SnohRpy6M4vqnHqnoO+gNt3xiHsv2+qB+049KfBByKw7WZIoZKgRMq3cyeQTYG22n1z
piLp6rlqoK8kUpvNfDP78CzCwqq41+vLvhx9EYV5zdg4Xcz4ncnZGFvPbTtrxFdk1+Eq6y376V1i
kP3/X05DJ5tX/E2FQNzP/EWjrxvTSXM3nDGx8GSb2Nr3aLLLPLwdcGHIMTdFUBETXgx6ee7xgh7U
uQjWmvWIuXcWf1H/R3R9gAgpqEWBQnSaSWV1GjNbW2DBxffT8Kkw+bvgMPlaDXkB1eQPpQm2MHRv
PS+Wgf8Cp2WUGR/+FffUCLyLwrapylnl6sy+qIox3ZeQKJx5iKMSAJZ4O1EljSDSZqqZn0a3DKhQ
lV6V1QxstnN+5+v9hGHM8oivna5HmDWfFInCqTBT4SneOPYZvA377hbp7pQPER+KnLBSKFCIB5Gt
X+l4UxIAfO9QHbzGEAjsL7MBbBxezKq6iAoBWQZ0Eb88q2dbtOLO9DvSvwyE7aFDAOJX2BDIlu74
6sNKUQpR4iCrGVG4BMfwiuonEag9ERpgLdhJVo1r0gETrZ59pQXDZOEG812UFVq0XN+tKjkiBxXv
eFYvoTwDAtKlG/Mw78meINUwWKma5HzZxXua6eo7eCrFzQu8z3GKeLHlNVUgsUkBD+twIwKwvrxi
grPmtLVwF8VRKoKkDCEsdf2pq1Po+/Ejxp0YsZOVyIPYugNphignjZ4LN4fatmMuGsO69h2AkDMp
W27UL7t6TKga+1Ezqk020timBmI5MxVIDZRR1OWYbQZA0n7nLtlhtiQTaU5ns/UfX6tXhzJok6lj
OzW8KtjPNrYc57RPqiCpD587D0F2aRk52m12PWvkD2l9mWqmsXanRNBWec662vhlMB5SSXJc6fUU
aEltjKal109zp251Kd6Kyb+oQUAj21azTHy1Dyvp/D0EqJL+BSuxAVjXKcIyltx+ssSjyTZIcWYh
Yc03RA9PM+kc6ojEeQ9x/BZxKWySG+XgFbJFIdfKgD1Ft44OZXAJ3hzNAjOFtwCgUmHtfj8JtgvW
P06PuLtB1ZK5Ibws6pFnUI6Jz9FajTiWgwWKdmAdq0RMKv35OhPeCZm8h3RbxHpjTRibgVG6Lo7r
769WvMUjsaH4SSJqziIXTA4RDJoXPjgPuudBpjUTGLexxQ/mzcJKbX7N7zNS68KIhVLpJmkJVStw
4ZcDZzPUsKpftAnNYhD8vMKGAr1LPX+KxydzzPLHMsrb7zJmdt2wkJbidG9jgxGAYd09BvLZM9tn
H25UHgOdQ7RcMSePkAZIPa5yxCnGPErsJVKjSuGF+XaRRjSFKvOt84ABGtD8wr0UA4o4oBxy5KNr
gJl81fvYG+Ax6ctvjNerzhi8VpzGhKSIiqh+A0tVnadxjeyXnrCU4QHApk1wFZzwlOw5+D3Uuutz
YIq50+2by8KUEy1UQbePYB8QibQTCjzE5CJofGvJ5/rDp1kax4qH9Lx7xAaMUoSgNVK1E4+YxQ/l
6KJp0dDZopTHbPPI0g9kwBv5TVRXUI6VfSsqNbIbsJbliDf+PjMA2H7PaFLshlMvWuAPzVL54Mk6
tGLKks5bKBAWGzUrZWCecVC7s40qxI1/N1o9d3tpNmibwRyWsdJpHsesjkMIfLjPkMMr4vzPlXO0
zoHPN/+Ofiko3mHTvfJQnx8wz+7ZYGHNB5CABbVQ3eVxqDYJ8+EiYAC2QmwIc6oXRgkV4trfawAq
qKgvPwccGZIhkX4UPWWLyAchlQqlbdSQsXD5hwemqZ+0vbf7oM7apY6/zaQ8zRS2jlAC+Oux7P/k
Q9HCc3bpFbbaLgjop0TohQj69B+h6iaAnMnnH9+iG9jNpwTzi45sIclcUdpeCpdL72y0q5HuEp74
lawS0oRKogO6Ngpc3fc+LvAh50f7Z2hllKUxVWaDVW3X2iYPOiMqysFmb/9Q698Eo0BwNbeIJ7W9
1cxU0iLt2jujXVyycLQavrkzjEMl5HHCnC8vjFUZkCCYyWjoHLrcpFHF7AGzPlvuyokCrbFMsBe3
KIzO9klGr4caaocEG3add6x4zcEgoyPKrF/W6vgU2rS4prPDeKnDXdbtV5eB+5IB1gUQrcIbcVCs
wnz3Zf8WTAnftqUG2kXAz0CdD/5nivdp+JN11q3vpHqsdk3oiq9JqbJwvHwnkREpEVcuHaFOBAOk
6/5pg7Tdl4cJ/5OSoQheqp9YHpqqYNvyDcQAsKLjPI4xUm4YCeoaaKipXjquYJtuObwiNPPwMELg
Y6y4RPnoicsVKacdr0DatS3udOTUFf0Iiv8WtalSOVU6Voeq53PWAgakV8NUgWY2krjAXMSjzZ8P
bV9n95bk1zFxNExWYTs8M/w4Kf8VTRfmxlo8byERhTVcsgB5/m6jSpnOq0erON8A+x1KaUDsvMoL
Nq1rkMAKHi8RAvho1LG34ZcIp/AHO9BX1L4HpbKalwsxYQhQsHjcHI94vFz6hd9O9AAXjQcnaKpk
eXJ8FT7s1UxSvW1pnCEjviWCe7ffFnmCRAe9tLqmWm4N0MXignzDkQG/lW6Tohvtk4lBdrLmKxxF
e/m73C5px6qfUDhyaPNT5Kba8+z/aIsvthEslEa1KSE5LWc3j1bl8iyDaNJPg11xqIFIr6rmfbFa
/nfX3NLMMKXJEVIo4OHMAAMNfQoMnzo7i/MBOzMwBfBC2A7NimChGuEU55alVv2b/TwpN3PAgys5
NxoM60KgdguYqCRIPW7jfrIm3aJ/5x1VXW78juMdRYJY00a1CBtRFGP4uByGxiREBa332qpCZ3vq
1ToWqjWSrfgwDqbwhui2Ja2g1KLZcROqqz27g1zsPi4pPcUSbo0Xv5iPOF72yhBVLqYOcaGHcVvo
dSNlkEMuxEQhO6E10ZGtB3QcR1W5JXBySpLQTfelyPup4jaxi2nUGMTbWNeLb9Y62gfwj7I093OL
/vgDQAwevr4meP+RdYKXyKD9wDMRnsQ0GMAYM9EX6tXGy3jIuJhXe47p2RS5mq80LSAJXrzWEaLR
Hw2kgXkgWMA8BBMvED2TGJo1VBJd+FNNHBybuKSdJRvCJ6nYyv+OJjYYqikrJv9x9+me4Jub8Bcv
qmJc0KBXhI0Asl6wFVfaiqp4dzkpAh9c4ZPjU90qxiDp8HCEQc6sEwYLRsvaeRQcEpYGbIrkDxwM
XZL2CHaZjnQyHEk3OA6KM9/kgDwhiteRPMBs/LtLr1KzHODi7u1U118FN0oJ2G8VE/DLjnQbWLD5
3MgbHQuCu+stW65dUmVXjVqD7XZsGPrZY6qJoiqO7cD7ADeSp6Kyc7U5ZzrJ4wj/yJc0X6768DuG
rA9JkKnlfzuA9KFxovLQrX4SC2I5XdDJI5FdH0LbLGRTZ/XHo8+yX/HHx4lPmcKvNeGB1th4ILGu
Z0/tetiZrdKwmJUrsLg0bp3F2UUeJAtmwIFqI0gU/+v8ssBBI/YXlRV5Wd0sZx2PK41OfhqlG+kh
EdUrJ9TIsJxwlZ2TLmy6/+JbAkCPe3cRqdGg4D8J7oCYTljKQZXhhyeaxqjGijNd3YI3JRuaLCsH
xF5U0V0tZUB3foyTPtrxu2F9mBTfIDKE5I6waVLHvWdhBzlFV0QNz+56pD851GuIMsGu7gEhxAoM
/dgq+38SJxsEJ6wpm09v+C/MMDGvLHI2FEOsb24Wi0nalHFOFipzrFRJtlIAXkRIptHPVxpD3jhr
fCOL0Sx5fvL5OgCZgEoyj9mE8WM6ZwAIUxSo5wONFLsZ2v/mOiRmaJCyAGPSoDckfh2oiRwYexME
fz0dIsVsGCqQvss+Hd3/WZMtLW+D2427JG75q41+5VNXRfAkf2bKPRoyIe7MHUkvcPV5X8Bx5qkt
dLAesLKmI3Pk8EZ7Op7/S/viBIsyTj6slu2J6p1/vDK+2q1WK/k/XVdp3oHTV/jL0n8GFi6zk7Ip
gc8htz58SMwZb4WaDA4ErNEDSuXsO/NoCD1fU5Faz2dLsTLG6RFVDopaxI4eXLUbro6LT7m9ATzK
LdimvPyfVBd5/XucNXgDjLlIbVCfZmEJaWF2XjDlDzYsJRGulzKESZYnuUuIiSUIBHGDgfhHiCnj
EdSlT5zeVw3KTo4d+jBuT8NGaKYp/276d4w7k1IRqWbzWth2qB5haOdtlg14Ct2iS01+zaPO902/
UiRYI07u57z0gS6aMcdoHmELMnFQCRHNwWirG/+zk+H4xtfdEPvsxxmejjvigz5s8SOBwMWCui2/
HcgoTzpP+k/+mmQokRBcFiwYomEOChO8yoxv9QvdbM9Wiq5/XHRJLgxWDJvyxuB7+iZXU7VEgRzS
y/JWEYt5hhh8Xpf3fkXkKvk7VHY7ii/6k6UvfQb5IGy8EzFxB5rC9fl4kBU6TYavvJxGhIloW2Xl
/k4m2DMYPRGWE+N5ZUogv/u3bxqFPer4Tu9X4KHS9yhmwMjAM+2VKeSjVILBQIPuGiq5jtKfLKOM
/qns6xb1u74cg1LZ62j71yKnqcye1slhT9+ddA2gJLiu1RdSkzwijXmaAfT/b4uvsZqFBsq/qxAm
JN160ZqMN3mWr2ZjYcYhqQsz8JNCUjEQPbPVqOK1Tj1IuMbe4niTpILMO2zhSQ9dZT6pPTo9hkja
gyBf9F3g6sCUaz0Jay++EHXijzbYYLA02lV5B8htvowiGTG63LofNPginUQS2GjiPaOvYBL4ccx7
7wVnXuZcKTrey3Oov8hNYOd2A7n3kUoyYnai4W6JlANxT8G1n3E044xfjAXNB4z8l0sOSigYvh8+
T9mxRIztXsyTRnTemJqmfK16iuC72dpRXyFQTpv9IVB/uG64tUWF5Oh+2TC5dzTY9ou4vNau4Jmd
1J0cNP1CiEoXXsVyuIBplhtjt4J83MM6MSQ+isUe0UAIh5GUWjcXgHk2y1qM/HpKt1wOnZ0o4Jmo
60BdtX3ZuPRTD86tM2OLoE/zany52ya+Gao5OE0BHqbSQdDj41SHUaxPlRwg4I3NHOdbqkjlGcHf
bHCdGQI176ytp7+2nFBnn1pu39TFQX2rohx+h1EqMvYDB/WtJI8KKZ73KdCrqcJnGqh7tYo7Sin1
Ae9lje3VubzElqmuwhE247rtDyqM4u4epLwKJhFBeWtg/3+RZLTAL6H3HKDgVo6/v4BjfHDjzXBO
NCWmrphY9hdYklK6ZwwFovXsUlUeS6oWI+UBaoB9YqElJbx4XyLqbAsFICAkvCNlHWw57o8s5Xc4
E5b3cezhDhbMgRE1GpDG3sFziaqgvBGIHQAjCjxURDAsmecFJ2MHKwYX4LW6FE0LkSORmdimQNjj
xsU8Ir2hd5oJAVHgUNs2tykgWqf3IKnNUf6M7/qjpKSQOJgm3ZxeQRFXejMhD/gxcl/YpQ8189si
I9aDSEuFpxR9nhL+81LgH26rz9En8JIhomSEZAcGcmSNBWamYcx0StCDw81HRg/aQT2QOKPd8Kfx
fX17SlYSfYiKoYEYW9SbcMZSilxaiFr6K9YsyRbZQdgO12OPQEhcW4pT5OKeqHlemAaohL6/thaN
lPKC19beFv9AEwaC3+oxLhiG+l9+Pqt2i53UpiYSLu1Aoxa1ylDvBqymFigmLfRyNR0WYZNbf+3S
OzoHV/nn9uOZugvvPE8H1eYUn/auPHx5b2hoWk5lsxYAWc/m0qDewl+/XM+3eMtNk8SZCjalG5u2
sw9909jD5O1/K+oeK242TJ9Q57LMnOpI60mI8kRnrydnxRNYq1Ul08Q3RpGnhyMjE2cBV10UsWBs
pd2xoMdQR4eSba4+UhGgDJS/nqlFFvkvuEbroAOXPFxH8xBEt4Xr6o8YeTzjqIxgevmZ8hpLweoV
3OlKBKKudwo+5x24BJH/zw3pxkR7/tln1kRGAVLvvONNT8+sZ+lOY4WaO0BN9EE+JLBYlBErVLfB
UZ+7xa9KOP2ECxfHjFnZKmg7h43i/9Hjvil/wJWh6nHa1Gr1jCPFNzBWsxxkND87pKbgJ81w4pky
JBnylpzE+tOhxJShB9IRcDnX/gJUex8ToyhrJGrhka2pxcNQyHfUhl4deHaLHBNMS81ZLGoI3meU
acu0X1uAhljcEemTHJbS5tjbQx/kpe01lfDDT3ELdUCyxXmSaPqQEyguWdLIqY4U2iLd/h5qiqCK
V1dsVPoDkWuNDtBvPeaDz9iBu/qSHtSMEvWyTfv+oSUHCmFteusaeNdUGwP8KX9MOiCxP1iONjf2
EvpnnQHzcD1Hms0Z+RIUghHqd0s3h8DSopMG8dOiEcwfpwRTUU5J8TOUcXtmYwd4tpN5rJYaw+Ae
IsODlbPVzI2NW5Sh/21SuwO009Tt+ySm6x9FCv3Ti6ICQnfM7sWGaSh+W+BlYYR/qfyw/F1neusl
3s72YG7ay2NbLUJgA+N3T+moF3pBP/3Ol5as5c8t6wSJkVvbjdhBW9blIM3UqoIFT/614onarMxf
U33k8CZJ+1hD4X0xTYL0TThG3U1jfjfzHU9Uj5d1Dtz2fmxpyfcyY7VbsRfAqEOy+3SfMpqPqJPq
DfUI3lfp0v4VVwgVpKiwL8oudxAbYOQBIbY3yikggP4KVBlYPc5Q0TDK/KJDWvrO96q7vZ7LE8mg
tCQjNuREg8lTFHHHOYgA+oL9O8Dqwp4Y7o5gfRPG3/dqwEcM3sm1UbaQ8djH8oi4G/ktSu9mQroJ
SUjY9HSflQbu56WaXSsQFVkqkbqEmt21u0Zh7vGNT4VxOYaWnf+pDvuFMEn084ijxAko8UKRFHAx
A3k6aVBhxbaIVUJyUMNGpdH8fvhFF5twEeF+OfeLUnyvLSDXFoakCmu9YQnXGp6+5qgfTajFlPct
wBd3WNVdJ9KyHuN48Fqri5OShBSHIWMyIofBJ97OXNS1/GouTj0YuvlyiTTjH+El0+SfUccqvyQr
wVeY2ssCi6J9KPW8WzFg8FCCyFrmEbRpx/IIfB8kTrFkiSDcG/nRiRjnEZa3AFrvv0TYChURUwGy
IAYH3E4rVvvs/YbRNXlrpk9dlAN8VyMGymTGCl//eWoxgGuzA+0drPG+Gv87eT4+Xo7u07qwuqj8
OSt1B8NqtULvqhmF9A1u8uAlvIcXXhXy+3+DGIuPWGwOFmxIb+ZVkerM0rxkk70epMT8LAHdTPTl
EwHeEMQ0e7G8zgJItQH8EFU/0H9JYH/dkWAAMPtDIDiyVnmCz3qUVGB4Tj/SP3ephUYm7arCVU47
Ogq/4cJz+PDFhyJrA7vuLhDUq4sCaty/Sh3S0xKjqr/SqPgBFXZa+oR5lpkdj4iGEgZVDj0Kjv2u
sjNSIF34C8o84Co8Oi2E57V4DM9lUed9Jb95WDV16qjN1hsMxKcC3r4P4Bb/Wd8obXHH2QZuiAGy
a3Xq2L9wFX1kmt7Uj39WiHI5LevE4yJEej2PAp/8yWkIbe5gu0ox7gEQoY/blX43GtJWWgiplGSH
fJr3MqtqIJqUIkjHLpbbLhH3rILIWqWbpi8FG1jvqnKwntszx3UY5QbC/2cA22GZrFjVa6lCMt7i
r1MhE/FX7r5ditnPINuABpOz1LfK0QU/DOxXPN/dtCCExFdXBBuLNlOovkfdbyEaknw4eJJIDZqG
ivO+advmoIMqZ2UEPHmNqWCEN8pXvD8/S1Er3GHzb0jBGKs0Ydf7rlIWXBtnBkGLt5fkVDO9ao1n
0LwYe25P1jxn7NqPlBdNnoWoco4AvqCtj2CihL69CR+9XLP2+yw6zsyWMBu5TbLZNx59M3ogowq0
w7IBinr6ZqKXtp2inFwf9iPAkeHx7OoMlPKNj2nGtpGOwitLxa4s7My6NE8/gzLOqbqOPpkFabog
blFFyR18gf/yi1x62tAGdTW0oS8eHKzAlCt918GyVX4yesNqu4Xdc49ZUWpLJ3p04KM33paetb4i
dGmjVtWLeRXijTeUq/JqH+q0VgxSUhNPXyNNEirVWJDvaHyX7jJCk5ObLqwJKr1eHfdzvFKw71ek
HBFMLDL7hI+6y6R+FQndwFpV85DlPFCXHl61YAQBq1PeULKMKnNa4c9604R9MYYYcCfBxR86FH07
837zDBuUhrqx4//sbYVAKFcrDo5PgbmmayJdHiqFvyKC13/STfxQQjvF+F3/lkSBctzsvAVrykR2
lHR2iv4iRp5kw0xcpdPtYkU8HIKBl0PJtdJT22SD6l5kshb7oChiY3lftt1UVGADUTbQJqGbVob6
mqR3ikB8mPyWzG8l5owQGLe+4Gv87XcFWZ8Weiklhxd8sTuqIqG4XTV0EGI5rHUqo6RAXf2oDX6U
kRRb78lDNn2sB6sMKpfoE89ow54aUtIK1qbks27VsjNQvWUQ6ANjqEwoia/fB0wOK1wbndQlQ3af
Xt3FP7pDnKETSEQe5tVs97C7HVIikjZimShoKjDdNY/lPZTYJt7ZeMJ/DaZR8Sir2CCO5rkskPwd
LFvphji2X9/NmTJ++NXk5KC8ZKjNDiWgw4O5CaYtzTQgWp4/vizNqeoIs6dn8xLRFAtykuhbXgg4
XkJcgEhwzDOxKVOmbrGGPTdgC5Rr+J/MB32xCGeC/Hv6Qs3loQ0zzkB+L7e/OOWWc154hLE+KlBC
2+rQnLy2I6xW6fiE1G/KGf/lYLr+cSSoVTDgtzdh+ug3VyKWF1BmF+Ny4IgfV4wY3S0KOhC3maIi
Qvrd6XcBVIztiq6BhCGHca4aWGNpyWOYLlPYXIjiJDP9xb3LS1U94B0jNvPiFltFpN5GUkGSk3Og
48f/uTnSTAEsgwtQ34PSFLMkf0olKDy13GS/Ns58UnakXLTmjrOIttNJh89J2yKPAc9/pNco2jH/
CnqB+i4Syf+kWj3Jp68GL22At7awN3XpGJ51P5WWjt6qYzQR39CD6ZpU1tj1dQAhBazHBCcrv4Y5
61aGhzOaS4L8hS4JHFid95ZP9YY//6/HVOozPa24lam4I33oL0V2CBFt/KMQWjPnnJ5OQd955RsA
q+7jlI+CPVuNMi4xBocXGYo2Y+yBQ5OobCi4TPomsMZelluDCBeOq/aIlTLmU7hz5OtYls3e9GeN
PZpgZlvtvOduHIEHV8CGQKrRhiCKID8pmRO1+3t17ec13B5pRqXiEXRA75XDmndgX6xoNKdgvvD7
J7E+Wb4giKdiSp9TokHD36gDc7mS5Q+0+GLdHq/HMg3G09m3BsY7Ke9x1WPyqSOorlxuR5wgamdb
x5M33nnb2by4iZIvyyliMujDRG7O8MWwUJg4vbDywFenyOA9MWBhyhsj3vXi/IQTEh61a5VAVrVB
ZwykO7sPylaGY5hgAHUI98ZfvC5jmlog+XG7rGeQHHuL3ewvQT2wLWw2CyP45fGVnv/I+GPsIG27
nASt16y3TDVdfbMOZcjM4MTaGwGAdW0J5SR5yF/nK/XY379jA4mbRmYjWnKjPOzbUmX4UA5bme2m
t0UyIQZqZeOWvEMPV20IEotstxjKWIg1rBexX6VdUl2NC0FHf7Vb9sOjGUjtIZnZMJyP27bAGdDg
PlsCjsMBFZH/qmQHwdDUar2LZf9CTDU4YsJ8zoOQa8nzf6UXgJi0MvcFRhoIyr/1RbQ7UrFvH5Fd
eBeR8uOdBS//7nRxYQ07+hXQ/nRB9E4uWS1cx1l2LzJ6Nr2iuPRDrpXreX9d/yFZ954XiISiK/xh
Gxxmt44Ow0Ul1VZ92EX3C0lj0fqXVKXqs6e2VbUaQQZPFeyXxU8+/uujcKf+mxbKwbi1YkXy9alz
a5VpNughhkyEEbArhBHe9hZtLNv4klocgpKpUiE3FKakiTG+uNtPJJSBCw8ANtyQYC+o1vbs0FGY
BNkxriaAgRlMB86a2iIgooZZ3PTRM4KN5j2RHlzyWfQrnzHkLQQCGUyfElWrXWcR0Y+o3ur0CpY7
D3Pckuw4Ez609bUxXLRXweAQylH+jwYcbBZkSf4PhLMgjMM1JQEcuo/XsFfdyxZ8XxsMlrvj/4xD
ckVK/qnM8Gx1LO0NcWEs1yg+aij+URd2ruVLk1g7dShvaCNcyclm6tCDB2uH5VHRom4gzhchor8B
WGO9uDbXETMk+kV+LEVdr/WwaTuT/MbaKUYljGN0dbrKRSxXmfkIWR2raqSK9czD7gMHiPB+umxV
rJ0HFOc7/VQrjjXzznFc9/Z/WCcq2eh5d0PyZOlZB9Ad0BNZr1Btiq+ndOtO6mrWh3ASIW78ABvt
uvIGTZ4WFMSDKUtye2+zu8zvngpnWysqIt+a32cn1ngSlzDH4nT7jgX4+w+mvKhH89jcV+pGnIgv
XBP0g5A0t8+hmHMTe+q1bMs7Lu6ykNSDFCvzACBXcXhz4i1ZHUXYRqa/Skcjy6i5IvVBp9AEE9+B
x1inGGJ/XX2V3pGyg5IOhrSbTvk5ynIB6ReKQJlBm6auh7mEDpcvJYhkDiI2RZYfM5VdS8fo00Al
EFLOGUwfJ9KsHPlL9vZB3M/Y5vh0GdP5Dt4q54UFYDfFxrKc2ylgamVSytDFvhdg1v0Zdzoj2A4A
69z5kpQBnerYgN6ykk+9TtKom0GuD94RBSZDl9FPN3qPOwspO+BhHd/tBn7XVUffMtBR2U9tESzz
K44KV1TjPXTiGN+JjuIKQrRF9cmXbIQFyBTrM6gTghykQFKItbJMQejckzdj9LkfldA1mbr9njI/
gWHY+8MhUi1WrPeMsOI2Z6DzM20bRywqGo0wkeMGsAj/9YQQBQtSqTmqyeFViyCDbFZ+kV3JWAjO
j1Tyn0IK+dbhuYtkWn3t6grPZqW8c4jesiFhI2rIvSeocDZLvpltufj3O/OoNRQPXZofh30QFtaM
TTjWBqAq6NTb9EcUzCFPkFY+Egb5lJDakgWfIWZOcv0OSTeRNWsLDM7EdaYxpNLMrdvwT+NePhml
+4LmAmne24M4J6U8pqfdYqY57mJFuMbmj4o+Srvp/EEeDs3fx3DVE/0Xkdar6S6RJEjPa3UZIYBd
SZ4wz+4rnEBSWGh/lAdGE0XvdR4/DsZqSrnA58XfM57RJb3yJhLl7lo5oGbMv4FshVG0P5pCt7u3
nSaXACXtdCZGWH4DtlTEgCweKkIDLwG+GsxDZhY/dBJJ0vav05v0jB7trmURlqCzSzFglswWVetP
90GesJskr3AhHxDG/RM0FleQnLSJ2ot12m0x0D5QyAZZ7aaFdtiCwbyDy7gI3OgNdTq/Ig95S6wA
DzSWM6WBZveANpIadlyiARsVBGgnc7U+W1YzpOm/LAagxEUIMnjAhKjPwrxBrbSf7g8o8Rh9f/AG
J24T8Am58qFRDF/ZrTif+vNytfm+Oo0cJCvfr/kcz3lhXb0xiNa+jKyj8rjWZ3CpQj5lVmkgta5X
5WKmrqLixOcj042/QwNA+VOP4kNsVQ8bjKlSHBWXUr4Mvu2cL1T5Bxs3Ocy4FGAjPZs6scBuKuC1
rlS7/k47la+5vQxlXiSWl45iGOe/MPrAgd7GpIdz1rgkn3HmYxq4oLyOTJFvKzaMfj3+NNYWDkoj
2L+1+5K03oKx
`protect end_protected

