

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nnA1LvIFtXuhnEgnrDveU5DQhO4oCdS4/TzHWVjuSWRiJTWamPLe1zKRcIJ3OgsD949QJsbaygaN
jpuk7BYNZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cfy8I58fHjYLB4BFaw/VxzidETwabyuF6c2nxAde+hbLnyzOfkymKdOr4Pk5oDTY4htTgTDRWzMe
dytGdfmZXjp6SJIGysindi/Logxabu2rWzFmbsNC3Q0gro5se9+3qoriCL3M82gnhvX/joJNLiXg
rsFmmSylhS6v32W24xg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gu3bZVKL/oo3WMbeK5OSi9dLiGmyQy2yONRw6Nst9yei3DenlP6wnhfHYdkStFXi/uvWUBEeZ7hN
0Bmqlib8vQ0eJP09mki40prhGAwrKuqYt+2JunlvLYMjlmKGJOXPgQJfoYTNzbZDTWMAPlUaZkK1
oZkHNa3Wtk5m49sk7N6rE0lY6V2L8UfgTL/MmCwu7DKHNfTBd2W2KricGJ6ICGb/eh21T7mo+KTw
su5JPh2xN6VOnDqK2JFdz2Fe2UsNNdpq35qIZsc5dRna+xfhp64zhbzGUq3oNeTCYYFL7/rkWyjk
xMfq+Y7aGpW1qrNdKLCLUa3C0oRubzA+yEUHPg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CjIoJO7bPG0vgefcLg3HndCtGBfDCnGBCSVZItM/kv6K6ZpvJnvEpEF/v7GEKszxgiutC8bTrPRk
/jMI//klbN/ln/AMlW7lDqpJ5wXp83c77tloVq04bnPwc3DaApr08oK3Bf1H6JgBuFfaRFUfxoRB
6anIIq6YC6xrV65+910=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D/ZhWxzQ+2vaiYn3/fV/u9o/WEb/ogG/V9KccsPCOCWeaD6JXzbX1wTvk2mHL3gwIIjopxpeK8ct
Dd/kho1WYC462ZEZ1ijvlrdcQ6jRucbVeVK20vWFMC1CO9YW54zFCdUIFDYoBjMQnJ6IU90guAMg
K2P3LVnqKNh7XA5585Xm34QBVEtkbFVGa/nBjX2k27AaOcjv8CeFc7ihUp4B6D6YzM34GhHkOxNj
NyMvVJlZ5HBA7JHakPw8PSgdpMIr12xEOrEcLpR4AR6H6hPW9blh2XXVPneGey+XXrhV6WAB7P2G
TGbniILS+ojY57htkmkMwgWfAakIRm5HfiYkdw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4720)
`protect data_block
5FGlaXEFvYTGVz9xDfJA5t91Qu5jK7nAWJkiLHqEPXyK9E8wssLlGBIrhnS3Tz2F9fNVTDvO9MHp
z3sNSpA52ZxCbRJbiJk2djZ8rhq+6F6ixa5sMmQWWPQs79mMmFJQBK5goBhR53llhar3pUh07wVU
Pxf2d4t+npAqDYPVKjO6l2IEKQEvFi7G0RfCCyWJ6Eq+fRqZFFNHkofWSvLbdI15I4wr9eujwGjP
30khv9IbUAEX+0BX4zdpjpKOUSb3c7o/oAodWxLIUHPTZlmu8M4gXVBexNmg+3hBgcRa3+4DwB6P
4gHtwlbpqu2WsjFVWHA1IqJv1QxhGkI/XWJxtpERQrZU0EFhLwwpsbgQotltrHC0qcp5TLkXGuKk
vkgH4Il9vSITmV0ieGTdHTMjOxjsiDtv2abdntSQVkBOgx7yYoU8f6WNgCO/TFXjjPu0rthU7otd
OQ+l6euKmzJporlOQcIQXo52MfHiqnZQ+tIYw7TnrwEVG/932ofNRpcqCftQYcXOtI3gpKvWq0yw
LKTEDlBTVrv4vCUR8VqCNsIBSY9NEpoNVutPD6+YYOnuVquwqXBiU0EzghaZlmz1cGT9ZlmP6Lnd
23yRMH/6MY9PJAAlXtdXE7Xh9VmHJAHcC9PCI/EdL57MRiBn+DTgSpBRKBEwyRV8mO9LXfDExZs3
bmQfTeHrBiRhSp31IZwhe1gCq/G3KzHErj35zb8ygeF4EBPOl+Y8ftmFYYhGddKG3jUfKlT67QAH
/acUgbRB3VvMRC9JgsB0U2XI0QAbHeKDSyOlu6Q1+DA+wSrfGpsjXiKmbiSvc7co4g75ykoNfIhB
VhHJXsJ8Ihn0Vu5Ld1T/nfm6b/O9S2FZQ+iOTN5hN89nBv7r3+jAE5fL/WChDyfNMH2Gz4we5hXb
4ztXIOxc31/fMZgtbyuN25tjlQsHHqDh9Sn1QW2sx6RSmCWxQ7GbU+0N2KvqRTlMOOvA5Bo/2cLk
kLKcFqByIZcZPNYbT2HAXG4SfzMVr41Xm3+/VzIkuX/7O+yHDspPcra/pylKqvH4vTNjeU7sF55t
9fphTBQo9bLtapO+2OaqsqoejMSg6zyQrGVInxXA0UKHYvLbknht5LxJNwlllNXG5hNZjJNv5z5Z
whU4lMZVSGKnYlfhkeUgLGTgapag+BJxOP3O+3YLvOT3AIz3dvPOdgaI8ACrRDTrrVs6GGRdq0ZI
JoP/cEGsgh101OlC9OYxqwNYRfpljwV9lIX2nkZchvnIDTLog1cyGEBWMDZFAWfZ2G/Kobz55kBh
eBslmU2NNXS8qRg9jHU0leMMnRxcisktK4Bgos7FUKDXvN7UC3a0tv4Gol4yGzEtEGMnrqME6+rz
4CLowJw+84Vc7n2HQWRpcRNlaD1r4Jw1zUOaD6m7/xCBZmi0RWemqUOtDGsziWrLjNgMkXhMQI6C
FeDbiPS68Pqo+2L6UsOn3DRqqgYZuwfLbMEDQVmFAdVTAJ6VIhFzpuSmnuWhbbyKtFYNpI6ZiCxd
7EXlBcmtKb7VoK904c7FSl9tULs5VrF7JEjEXIuwZthMIZRNhw0YFsRmBSYNSrqNl/3batPrsNXh
2ZgKzvqimZ5TL+FGw8UibX8DLWRnptMjsNGTSUSenzF1oa7/x/yqEoX250Xa5SbgVXklNh9jxNFk
QCWaWCd4ly8IIP6AsphI7kab5BzuHNwyyNscm0CCfmF8BAID9kouoCMxgWjBYmUyafuOtAj2RiS+
VlAdQOg1aMcfI3L3yEQ/JGS5ffgmaE8cFCCgdgJug7K+UqC8z8Gd8D0Z/j0IsCq18BFti+9Q5t9h
5R/+uE++EqaN4QTpNRJTcqcFGuJiX7j4kJbxqfhPgXIwwneM7HlcHL4eWVSATHVCQMx6lVKZ2V6h
YuBYPqSL4UqtG56yXPJwglU85ofw/Tw0GFG9ClUuIMLNB9HHVV0dwImUqH0FLWjQ1cyN7fkTBTwl
uhuXF0WxByS2JDZRg6I4kiBSOkAl9OcmI+tWv0JYRv8PCretQJamNNCP1rXTw1AJPsLe1EsPpzAW
w+CH4MZMxQz+XesjSdtlIuBErNMOWCF93n7vBit1Cfw7+XIi4ahG9U8QHpVINFn8pnPwgBYzCM4c
ofFyeU4cdGZvWhyyFiIipbZ31gu8M/AjpR8CfGceUpsq1x9gaRwpxT7W1zWG9juBA0FonxAcJkHD
kTK4JyNU7qpcNpMtcyMw+1Mde4Ov8bXLHMqLOtnt4rp/AjolXuWbfSYU/XFfb1VdsQK25kk/7dJy
HhW7On+NzkxJX0I26Komn6BRyEW3Q+9jRa/sKq5pxeDrBUohqBkjWkI9dqr1Tqhh7ann5aXjh5Gv
NnduCxCwFfXHxyCD9iS5yiYKSlXFWUCblOOiW81TnZRCGbpVW1E9B2VXvVDgvgERe4DkCROo8Ycl
eBEvBtOtPV9za8D+CNHhdd4RUb3LQKABWhSbMg28CLXuuAGs4x+G1VesEsa710lPgDIerlZUn+i9
MKOG8w99nr/N2MZZEURnSSgOlIdXOsi7JpnNKwSBORKRkFOmE+9QVOwJwtvu9fGKI8jEfjE6oh/c
ZXRFTPeoxEnDQ+bE1LOtyqzDzECQ0Ghw/b1KOXEpdjI7c286aJWhoKabj4k36NPwmWev0Telkk3M
RvqhivoxGtXat1fHJbRKuRNHZ9E73K/iZIUMq1UnPa4bF/FykUyFNKFNNWHt97soKqcMCqDS9ugx
Bqyi2mdbszIxv1eIAFEhI3LTPEdPhWNU2ZIL0/luVQBXQfY41+UW7OeLrWRwNG1jepx3VIryT+79
P4Ho5WU1YiH0yH3f4UVbec9GUWTQm3DJh3hs78q6D+d0Y0+c/xsfzMAyiPrPtP0b8D8NZKbgxTd9
RaVjllerB4gan1WFYcu2VQy8JTsAqZnwhxVYjneuKAbwJqh8vklKcvz41uo5pIbAlmXYn4OrFT/i
FOIn3g6J9QI9Vx40KOqdhw7c3aepBwzud342bfwDjFyIgzl4abFLctqlDI0VjiV4SKVUX4iMGZZr
NQd8abV4DlyOI5pel6JxQZRqII+EXFMBVostfazaBs51tTy0zLxwS1LMY0SeUlJ4mm+jhqcs6RR3
tEOTamPQvcn2JVEHiqHx23PpynmHQbZoUGVimXgCY3QEGqTD+I/Fnj4YVHAJpgcwmJUqsu30273F
z8Vtb0KRr77f6YRz2RBTvYU1yJzk9NPtuQcTqw3NGyiFsqqAGK1SjGHQToP3ADR0UXlzw25AiFDd
YVBS0dwEvuA8wBcz7X+HCRLmdXMym4f+zPsTCHVShLqaQsHMYTIAY2fXnCYRKHHon+qnUOBLCt5B
8w2DcV4JEZ1lakwHz68Yfb9rnahAzbVtiWkCJjn7ounT7lA8FsG1AmypDwXB98Pu+MNBaTm/pzvN
2PsK7gBC+IIRi+g0JuXMVpOHMIxxPdiEVyfoRqfOasRtDuZIL4zNJLk3YYDTYeNnLMG976cZFblm
U/9NL+ebaw+hnkKcw0nIu5USHwbaNBN73rqXCJCW4iTF5rTPDFKzLcrm9LXZ7hFaZkNkdAcGMlPa
XENFUR+Ow1f7ANx5Xvt3aYmsJRP1dAMK1piMr+PhHkuDbdcr8+eHKl57ceDdZiPqM4W73n9giMJd
Gv332IxfVFHDUAfhEZKLxLRrbGVlhO/nqDjGb5XjGM0JZz+jVmqbZuVwzQQo92UGw7yt1TzZCkMg
gnfg0F7T2qVz7wF1xzZ2fTIvMws/ByWWflIn7JuW+oH84qff5yo3rxnpxA94AFToMQ3tP1etnCxe
IUYbPXPTVOrS81ete3zbvuX3OIpXRjvYixK55BWlyCzhi8XJfZFrjvFT//kLJ7gRuiI3YKhl9Yxz
aNqmEYQSjX577GLMI10NXKpWYabR/xvArs76u9M+FQGANuijGjO06B9eEbKyW9qvkbb3xOhGOF3s
6x07PbqUQGE0v9yo+H0YzaZ0dTUp/cBMgsevOlCkffJj/IpUO4QMntz2EFsqnG9593MxG3f1+9iS
wmmhNxWAOPq3tuvzC6K6fPp/ekbE38bRpofN6KojEKplUs791eobI66HwivpjdTiLSajuurxycd+
M0qqRJCFIpFAkzvPrkuUrUDGTM/Kh7FxCng0A4qJzD+w9qbSlgKWCWwTwhWlL8Ws9dOLXJPv3SeX
ilw1IOn4ocgNdclYDjWRrDpGe4IZMa9QKvk5zIRef0R+/qZWwWZC070zZ8r/nR4LxB8V9N6IY4Pc
L4E4x7hbwkhzaTWuVKO4g1qOfs9dwvor24LUD+EFHI1G5ut+MjzLPvzVfz6c3Q+5K1gTpORXuCYw
Je0SxeMk/XDbteIVJ4A9gGgGW0jLkf63FrogQvqVq/8B/z0dEW3msu9RVnycgwEpeIgFVIwxGTBT
WKM6WfHBofXG7LKi6ypTfPWsnAjmWrx7XxIi+zqU0yXWCuVTkkSKXZ0E22Nel1Rhppgw+TwvO2BY
EXWzpocJkcbaOs7oAQs/cwvzmWHqMAPTnxYHk4zgP4tbkRKZD+a/1nzmRnDGtUHG+BUKSHdSff0L
KtY6r8AEuDq2rDNoN8OXTY5oDgEOlXU05+QPkeZyezHvOKk+Aw1/89IJ1OBABqYYWttt/6Ctebk1
DD1WZtTdqix7KI31Np5+3d6W7Yo1ZReL383/wsNy7+WiwlWQQtRy3tA4LcT5fxLmsVQbHtTPdGyy
/zNij40mV4LIjPWxfcOCfTq6ozJe7LuPVUSzFqG8BpPsbwmRVFfOJC4NXm/BtuVrEIsgoorU3Il2
UuomcYxG6Fm39n5SGQz4C4VMdoc1JNJ3KZkq4RE+YcfmIM8+1G7hntpPXVSvX0z13EhLEvhZcSc+
BbEZx1OcfJIfKi/2P5Knvun0cOaDiHD2RCZayMxRWp1+v+xYGIfW0nZ6creghlHupdSXaioHBP8I
MyXBu4/n3kUJk4jjQWI0Fpvk5LWGW4uZmcdHcQm+whmUdGnHJZFBniG6kUxDj4a3QAg5/7aNUo9k
l/4nCoP9zJOMnqYtpYDBSm33iwuy/Fu65A2A09UKVImzXN4E1FZ2jkzAWuZjRUkkjlyz59tbUBTt
/9KIapQ2tQs4j5rFLr4/opONqz9f9e0U65ydhmvNPQz55u+Aub10oMfTb+mNC5rREfY6B/tHwcMz
I5epGZbYpd+T/EIPBQUQQmBN24UdVwfDS8dU79LFxEOuAe8CDTkFgdud/yQgUosNyR8hL0roXgn8
2Ywvg5aYu6uwPSqiP9lGz8cQU8JUM2/X+/opTHZdoj+FuX6muArTQtGR6ikEqqDyNsGPzY5zyF2Q
4eRrcOTdjSUe5qQ4RoAi74aq72atTwfWFKmcBpysL4azbGEgATGBikmElAy4ize07j+AdAEUv8gG
uydfH7wtejz96JdKBzYHdiWKNNDs7PdnUOyZWbH4fIwHVSQ06ln0+j2HZJKB0x9RSxZqKRtRB3KP
E2cqPpb3b2hj95nflyo6fBsbCTtLTUhd8qb27Hc1b8VYRehfLxKq1AwchLqq72rcxKNYErmwQ+yF
YdmIg2GgplimGIK82bErpjCKvQVtyAWTbEcGCveSXgzOowusNv5Of+K/i8SX/TS0NZnqlUwX51NV
twOfWk7crxOu6JMcxfiR9WHDtcKV6d0w95uFZEPkZZ7VWJkV7dec2L3GfCHKTiAeaQZyAmVdSRnY
F2LuWJeJgwcuEOUhUYiW4JOTcT9oRWgvUqZBWp/QS6+0Z3BseZOpuGhMwB71v+3/gJ8pCnRNOcS9
uFX3+XEQw0vxB/rrj+EdagL4IgbiLfcHOfXSJAqeTgqeAumBXQbcRmodo6CNw/f0NNDqkyuoE7ws
0sTtXL7DgquS4JHVCdhhoGCux/VYq8XgsibCMZC1bqy7xIkUGGvwURuK5xlzVT3ESa9wquEIA6kf
K7Bxwn8S4rTGrXqfz6bAr3+pKeRcnYIuXbIrF22dW9adMfhhh4d3E6o7/Osdy/52M3bfr2NaG1IJ
p8affE5aDKG5wbvE0Vlu3vIHTcIRfctzLo3kuY9HtZorozUqgGsipm9uxxLy4233PvAHrgVZlMZh
Ip+lI5yLvqCN0EVjjnjpepnbfYouevy7k1Df4N40Sh8oq3CBABJ3Nz7sjpCrNuGyke6Yl35gPyv5
2vv4VS9XTwNw3NjeL5c1MGak+Uc6Au3ka482yEoXd5plGsRgtXwg5VIpk/SDjV6YaqFSVnSqFI4V
puCZYQU5u17f9Xii3uhkUg4+vN7zPzXMagv6OFbQtc4iW2CZxiNOKVXirJBuqA==
`protect end_protected

