

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IkKQ7UnyfG/i0Gz2KESfn5rIa2XG6JjMuNzaLweotYfssoXFPRW5MF9/SJXIBGc5jwrrtn7ZIvXw
ZMKFyJ3FzA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A7z8fuAKplZhDCneI9mNA3lof0N+J7iQN1H5R3Mj6yF0lZ6gCWQLLnnmsEoxkSX05NXSzlh4gcEg
7rRfO6LtEEhf+XGNB65vpBYpfhGyoq59NAHhGVo4SvBM+mv7uMxOGdpTeOCZ4JbHV0AkjL28mjov
93MegfTkvdkm8J0Lvdk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xuMQUwo0GDzI3cOEq+tu/2nUcDmn/7fhQTHPWWNseJwSS2v3l/iZo4evCcnhY45ESTueA+ZpjAko
WVoSIubelzbNSlntY2uMGs5oczMZtiztniKkMtgrjy3EW9dfGbHhtmNrOHGIHH4IdMr3kAy4Vh74
ZigAJ9A6+7kI6MsJi8v3mT1ARZHCR6MWsQMcVGsi2drnsGRWoYryCO5xQR7B/cwBGzMymTal23NM
pQKOm5sZ3P6n60ZuBiOsJmbRp0+LVYxKNhFdxlNXd0mwyAZQT/UOuOuVbjlNnKY3+syFmjH1X2jU
BRKqD7PfkYIVMVQ6XvOwQSNLyki/t/1FG9LntQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2lTj0FQ90PRwxkOhP58Pis/0pnBIhVIOGqxXo4lWUDsJI5sRS1Q5L+Q6i9o+BNlX2LRPYus/9Dnq
5ATglZxA4PDv34H6B5xWMxj6PrHSWzf271mNIoMFrjsSBdzp3H4BqkwksoU2N0BujU4mvFktBj6s
VuYwP8rZjGtZ8cTr2i8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WKc7lQN7TOvrS4DJ7NNUxP98rrzfIQuz4DIZ8eAY+GKFx6NuoyinV7kCt4N2qBg8IRnkz00LUdTl
h4FZuBrLJJyfOOGbqIiZNIhgdqVi7fXcxV2ef2SWPHLvr6kIV0N1TmRIBZht7FPZCej+/BNW8QYG
B1Rd/mmsAB7hXx6GfVQ5u7NRsVDyxlcEghLjiM7GAdTaOWl/F6pDM3aRwjjOmid8Gt7xmiYfPT0B
Gzk510O+OqDJRqmdMvwBmv3K/y+M1RxYsLOpwIle5lGrJoXR6zj5dZS3g0EOtylaiuYJczAHSe89
8ncn00hUVfz/5JZCkfgcxZH1LxGTI+Ly2xY+5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8544)
`protect data_block
59F/ViWjedIxI4Ck3JhQ+CJYtriITYtu8ajvs31mswJjEjugSHbmhxVRHO7TVJGu5ch4yY1DohTS
Kq8n9NYTH1oQFCdm5gUDPvIDPPswYwC0qfbzDK8TWx9WQ43eZCNMmPxvBpvIS1b/tKzDzwf8d2j4
bj0M4uj3B/KAJi1l5eVJqIgygLLdzpX1FPIkarKe0UH5KB5ARvlrrdqhUbuADhmEgmvq3A3zb352
GxefIIJ2pAFjrc+gx2LHzWiq6qhbsNGu3dq53R0BUGKaCP08fLohTagryE7eTvYvJeL4SF5IH5oE
iMpjDPaJA4uaII4tboh5cSQRspV4aSakHNlgHFNfmWVng3g5KedN3Nc3Sn88iXh4luDV5dj/MwnQ
BHjeXAzf0IIq/vO4k0F1XZVaEXC7LCIcpOlFPliafOHT4pu3R9kKjHJIAHSoqKuaAuBaDmM2Khma
vftoMAna+rCviV2j9PQU2xH2TJs7CnO1G+FvbO2L3HDQ1xAd3Ss8SybX5Hnoxa9lvoh1Vz7hD1F+
MXKSgcVvkJ+hupxvuou5i+lJYcPDfVjMP6ZDZoAZ9pfLBqxAl73I99V7CY+nGjWRgt9JdrPduUYI
pgN1OwkNbDP6aOAdhpiG3lw3bdWEItat/dWbYF8cLfMAGePIw6C+3d9w9BcDPxdnxX1XCYawoLl4
F0TWjUOBcGsHSBPr2BAWyvIWnXM/Quu4Qiyyl2kYHv2HnakMf2Y53MtdeKR2CV2z6xIgGyM9Nwp7
owhuX/TuFzwz17zQl+n4eu+YRbQQ2yegfqiOXsfmU+gdf40M0yGc7oetR72lPiUlMqQatOZG/kmy
89WatXy+XcZOhPe4iCv33AQzsOXKgZZA0y4k/ADepr83ldI0dtOeWyvtABJdgrbGiScCRLSPoaP+
hX5bevKmmYe6xF4ujrBKOXCZuz73OMG2KwP0ws6JjaxlH774JsUOvoHAvqaGMXzst08jC41lNnSM
XmhQB30jVpLeSDQCN/5YKp5o+//YYDTaYmjaXTIseceLTwqD7qiVYwY3S1/TI7qlBTmCwKZ42IHW
sx5L9GWCjDxpDwCQzVSoVRqxjdLu6mso74X+OvtFWl1WcXgkiNlE/g2lI3OyQW+/2Lfbya49Hbjd
RvgpL/VPWcl7mnJS7aUWGQWnWldx+pIhr1ZGu4Suq6Wi/8WZx8FpDt+RVO09IL47rQEW4hIoEVgR
VQBdmwinrG5XypifUK/YtK8eSbrwYMJR64jkTtPGUy3LSGUWlwrslvbuGeurKDBaEFvIDMfJF52N
SlpUum+UptqEbc5M3QFVqc3ZBk/5GSUauHHCjwHOOfmVK3WDWS8EYw2XMKFy6ODtxak9yCYDyeae
rwvOt7w9XBNKUESf3laZZcVbigZzkT5S8gPqJ08ZHsEoJoQCzaaLHCmwRMunVVY821bySdYoyjYX
UV7gyDnPLOgsdeSsO1j+YWV/YvdrXilb5Tej1tdfklxLHpgS0rSC0QmboYlKzPYo9aj7X5pPz/2D
kEFAFqwXsVXkAoYPTRDdt32adAIWwC4tprEBSXbAs6eORIJOL/ju/d6WCt6Vd4cgsxniZt7szgKR
qppncBYDqvEnMipfyUeEMwCazFNuBZe/do4nxZfMTIL6O4cSrCXemXI3Aw7NhmgnUnzxBa3BRMyY
Q0cdmOWI/FwEn5F6C73B3dADrx9DSXZygVg3piZOTMaE+ujLxE+dKzmkYalYz3w50OrseRmm3MMv
E88qPMtmqrPqx4p2aQ/CPpIXXHpI8ExYus6j+Qy2hSqbQi+V0Ne6+3MCTbWIWJQRZwtHgc+oLoyL
l0xdTputvXriyKwaOvxXtkhp4w1d2RyNKqfRQkrkFSJXKF7i3Blt2CCFus1+YYdAChaLtyM0RIbt
9abC+8ONFJpSMJcc8iE4QzXiTMy0LBYD8sq7COmiB7XAd1zj2ns/Is6V9M6gxx/81r3NjwqzqMs0
xRLzrmf5TmtOPepNDdSZ0KzustXQ2wdPRmJsXZHLGemRI7Gv/CjvkCn8ChlRHyKNOEEwNePHt6Qm
e2C2tYFKUbts93VbrJf92bZWostvcjdMK2ocokWXTFqsYF81exVsYfa5kPzO8pg0w68cZ5XXLh6z
f+r8YdHwrawpNzlExwCWpGZOASfrVbvL3vdEuqUm/1N3+pU3dujAia6Zj1RDq9a+/rUUR2j2yP0r
r99CVBGVp5/bk20QrbshHhM79Ic/fYGv+snS3JsMSMqsE8fsLCydXl2A4Psk47zLCHhGDOolpM+9
FF12rDxWNo8TqDGo4tyAFtM+NWknZj0+V2e+Fke1IgVVQAL0WQlA9QWMItX+AfBNs4eq1q3bezzG
MahUOcl5tvfyEmnpaz670TiUNveWR5m3urNIIQImyqUlmI7K5YA1tzxgp4RZVXOXYw5DKmpuHqwr
/Rs3uMBI9mAUcSPwYikzLlQLwQMLQ/BItuOlFjRxrc5gDvYzaVXMMGR0JMX3zE0//s6KVQ4n/3Bl
DDpHN3tI8wbIkI7o6cg2irXDqtU4Mz8XYnUycBtYqebRQuabCx4LKQgqEmwS7EQ6iIdUMLsfVMxJ
6S/cgiEgCdMHq28ryUygSHOm0agH43C5o03hljeQpHutIxe+skdh7XhrHt3+lA9vihWWM10qeyVa
1kRCQ3AJShgdwripgAe2Hx1bOV51tgLbQGap9pDy0XUJgxOrbNrPoLk57x/N4kweRopsfSL9yGL9
Z8ahN/GS3cebsotEt9e0qTL6rAaXaiySMo/QIjwvS1BxC5vjhnOysukri2VR7qtorb1kIJtc4knL
iDKmHvQGP+s4P7i0OSRe/JzbOyON7q0J1DdNWfq2tEatN9yYkXJUZP4GpKWF1+6egffUuEVi33Fv
2R4P9ZyVpyL1pMuScmHhvDVCtlrrQNLUOmAahbXlx+x7Zg+XzeivaTl+26zVzUh9asgOQrJZI0tV
5KpzmuFV2LqrR2lb91SX5tp8OyR7zqnM2R2rPhBzJAjeB/JMbX5rnkUpB7FtUr+t7ap6XzpmawAR
J3GZ3PUuqdhgaGRyPpBnCSnKAczIJg6UYVilSzY+sSdy8A8CVHBefvc2l/YvPaXx6bKtSssv26I+
EKE4TQAiHyhXh1veaiR4U0wKp2a+DrNNlAspNkZVrlhSaPf+ZhHsV7sunbH2Zq4M65rDxhRWmefl
64fHf8Z56dEvaLczaFvvkHyxk/rPUs2ev2vGN2ngHsRxn0YG+PJIEDNLRCXyMUIa+YfnOSZZ4tJB
2kl0euE4Iu6f8hI3Eh+xAQuqHOJw5zjIM3rinKOVNUmRf4E6zjuX0dg8kz9W29x720M+Osi47TTr
6KX7eT44KEKnzThzwVzFQef5TUTVnaKGibcqiW4nwK39eWpvaIDDqKaxAVXuFFmbXvpmFqrxQupE
p0wHz3itwkedXfYUlrB/8OzcMhgttKef2V3Fvtg9bx6wUtEAyDwdBPNSIkcVdaoWls/mCF5DZjuO
JPKH8rFklfx9UrCn2KNZEIWHDhxhCtCVI4WWXvWl2HSdrpDFe5cm2WzsUlrRu8mLEU8j5SyPxSxz
pxGUCIdC9QVAoQ0ILjWhLvXb7ZNAFS0nvOB5phg2JlVzYMCi4NZ22m44H2YpWvtJs3ncAgd2kgpe
ucdouWmK4j3RxvFSd37yqELhqNE/F9m2rBHSCBu4H2hBXfes2KjKOb5PMMySIXvBW0s831ATaE6Q
AUmjNxO41Bktr+vZAVLA3xgMAGdCmQ9nar9XdILTV4BUPf4tj3Zc7p6QPMFLDgPpbuoDs9JM3X5c
zAGK4ZAsEYKZ/bkIK23OO4OZ4kVULadZ4BniLQDECEPr9rJNImbnVSrYCkk4UABZMP0o4t3Ww2gj
Ap6LSgf3A7qtyN5fTjXoTncsFIXk18VRhPWQT9x3twjmfZmoe3uHsTxAjlYcaLFbwpUqlM6MCHlo
7mahqneIv/7c7lADoLxOxtTTmkXDF29Qaug71DL41DaVRrZt+INCBtlGCwLvhSgNqokZay0JuuCv
ucuskXQ62MxbHl6AeQNP/8Tw+Fb6Nj638r5jDRgw6IoQyiKfRPA2O1grZOJNU8OMYzrVArdWszb7
+ciwGhGLja/rS/xc0/Wc2iKKzpdyZZZ1Jdd8NIElTpQ6SBMBPm6RV6PfSPZ2WwfErNJiyv5ICQud
EfnpEPiBXj8kOm2JsT5ypQoeBpgMz/G6FYjsp0QhIOKWERgIgOT33tpBXud73mhcXmX8/XOzr8An
Du+tBPH9/bWcXL73EVm4T1WSGJAC3fKB1/Dik3uymh+SwJpOXa3yyIcuE957BG2hOTRl9lGNPmvD
dMonV8zlq3WAki2JT2JwXDlvbk6yiqgpTeI1Ko2Lcpg2fftopqolGOv+0bOcEVpibT517mSTVMdR
FiXTWXRXaYeM88bgg9GIIdtwVzDi7Ub8eJ7g7piyGVta8A9YcNgrSV502bjHMfp2CGLW4hKSIKsk
tooQZMC8OJBEgAoZommzmrqKes75lBhUCkeqOYW8q3hfTEciDrF6UNGvdUP0sQU01Qyxb7/iKVlw
Eh7eeB3B0owHXsxyvxCwXveBW8kDrUQFyTHdyucRi6kU/PKVh05T4o4n5ioFjEoodEADn2Dl5/ci
YC4mfMHz/WWptQ2rWAe3cTo6rAfvayW6EY1+Q6iKH6YURkXZYgz462Xz+un0IgsQM3o7ksom6Z3P
g+4SU/dKnF7v2DqNRGGBgAoeYdrem333uLhSOoTF0bIax6NPRhoruVS7nBhF05ZaKm2nD4/0yoGi
PSfeRmQCKv/1CqJhaK7MW6Qm+lU18tAo+75mLBlmvsrT4B4v3nLxU0qRezi7yrwCvbcahHeegyvl
5LWhtrfeAdDgHv8hmPXcQqKeeOMT8wq4zn4zstdwXT2wIRaOjZHNoHkSyse1Au/DcnPHRs6WIP8Q
MT0jwEypTNjDJDeQVnFI08zyWT5P8+HmeBYnZOVLKVq1Lqhma2aNnI28wL9aN4zzgrHmPrINBrg6
DtK40xN8xkrJvyeMc2V6Y4CfhgwI6KsDX5cs/LmnhidGwSWLifde/tCMlmQBnx1RvZU5Vx4TbKE0
rFf47yqU7F35EtDIzeQ7puWGyYdZxtlHX5WuDwUlU+ROKafFShxPXj38EwJ21BWuFggDhp68bYFh
TKogsqmnmklvkN0JXnBqOcB0DYWOFIsRbcCfe8xj1EGJLOFEs+JyfguzHAXpnBbxlBsv9e6dHX9o
KWme2o8PegFr9zG25XXGgGwVoiSyNIXlKEToHia0eENfAdat2EmZdVsaHHNhORzZe2VOYlsscXMc
Vj097jsYKzO6O4fX7jUCmkT0i3Q+LqJNfW21qEF2zv/7YMFvb8qeZ/7GyKJdl91NGlggExejQi/k
Y+FHgwMeTE0S3j/G61d4t5QNrxntIaQSPiCIelCH7rBnT6Re7YYZL3Tz9B/T6xIjPxvMueUBkFpy
FGWuvWiS8uzMAt6D44j0K2trfj0W3vD2OtNcpXPpidoomXK047NmhwPk8cwPi/exhJ/8DGYthjxr
KxyrBDaBXY2eg7Mu7LHul1dr/bS/b8GRqvj1IWa1e0asl9ty3EMuSHZz/N4WWnNjz6ATKQ0j/KSh
TI0uA/kJYPHSJSm047x+T0aQjUvCAiapN4jtE5i5Jee1P7Ypb1+HKqdIuJrRKfNlVAD8CxqdftWw
wYb06HD7Xs/QyJwuFXbKDoLK2vFstDuN+PATYcuddIBhZhFZPz/Rax0fk5rlsccIL6HsOdICHfs8
6xZvDefrBMZCSavEEbv5R1UQfLP2MVpRAcXxToYq/aUTboOvSFmwEBWBl2yIrOfSJ5sQqV9KpMjm
dJDPo696vS1iUeFSWlVLiXx3fHgxolYvV+f177i9cluqFAII8/YXHFDcfYlcr/JkFgERi4fj/vST
4xmPnXLB4e8mET7UnlB7UlGKg7aUy3kjzx6huLOFh9s2mSwH7ECSERNP8O67VF+CQ99bJBAYBCd0
JNceH7c9lhGcesAzCdZEIR9hnRsirjv4Zl/1c/8ssk/OhWmjETrSvGdmzkGvu2y97fQvJcZ+GuXj
qke2kivcCdMepXqxO139I/x3u6JODA/p9K6sKkN+TpGCcPSRjyTiy/JMwhDnqWefPYmfIjDv6eQG
8CWS3Wk1QHQqHQTKUerFxTGpUCNJXbjI1D3mFQ7y0+BexbixT1L0/ydxpyUMhIaFLgqVQk/XX03S
MdLIHNnggCcGxTcazFaoC8qWfEKQXWH+XtyGDK3Sic6136vC7gbXWr3ecpWm5R8x69P43j/6H+v5
22rfMhNUgGsJHfAB2Sdb76/hDnbIHVyz2hAps6+zGJ47mdbEw3phpIPlakZS2MsM2YnV+9pbsdR/
vBYkanJ1lB9YOPnps+POPGSk6LgFFOIfRj1pYBmxdhCfduGwOQlUApx6Qzri9UqnIJMKhhd2PUGh
iILPfVqOXqkzFuHGaYViQg+8UpPK74qPosjQuastzjVGPyiiKLnRnzQN1jJIRHs1mYy3PR3eE7K9
TePgH3sKv3U1Zqvjw9uKrinoAs4zZcpxzA4nG0Msq7CCfEm4jA90iDNwi/TXbytLQmPABpOwoT97
CO+N2ukjaUimYkkqQhCa6VEadnU/Mw+/KBcY+BOAQYd60NmIEHmnc6XOlurvAn7RX/HEqnAd99uk
0E/wNn0Wz0pOqgW2tbnT1Rtqq8MEw54uWfCMZXyu3jMuslOZalT9qjCI6DdiWGN81mhssPfNmbKi
EhxFpRXvxVbd1gCoGxQ2jrTvRx+thjE32hZwtYjIsKASUY5h9ZKRpgAWWAr/8SkJUMa79JCvmb8E
GZTjWSrlwKkSg60GVSq7+CScP48BoLAM/h2eOo+KX99GG3fUG38pTX7IABYDw/zMsWaWp4sydP4w
vPWLRoPOE+EHkpz3rTLQCyhnYvzcStgc6NTGiK3TY/SVU20dJL6gDVEiV+c5xQOekeHKF8PLkKdJ
dvSLp8R81nbgKCLsoEn/FIwLy7RYTGG9KP1mvsumfBSAL3wK6Df8Gx9zgkhnb5l7kLO6cU3cI91y
uWuCXNJb42J57+gldBzKOUVvF0usq9G9kbb9mgGLcM+tlcSobEcGpKoyatBlsl7kbJ86xCrKr+g+
6R5EQ7PIIMNdMyLogTZtedJ+5ffNrflo4IRd6fNJMEN+e2eH62q8inMkXC0Z44re+nDRLfqRjCNx
hJF6NIBT98dWkXTnxI1rcL3TkNRTxkMEqtjUJi2varcgfTOpomxGESa9CjC4Z8EGwfJIYZ/uzIXo
bWe6MPAokSuPrZuAORF+XJiCSKjPVCbqN3qfKFZ+y1q90XLmAZi220NakLxda3DslutknQo1SBcE
HS02Ucd/T2jTqRUtrL+qd9GjFHNQcqBQQ6HHMZ9ljO34BCeYeDxcEbtGGyKynebaWZUsVK6Pqgli
QJPPmjVzh5zrLrVa3FrWmyNNiBEkCPukXQMTJGAjwhM9Jd8TNxLGDeQHC+XajYcMcphyb6hcSdRs
lrt+tKGmTqH5x+DMbJRzgS38SAUkgqKvG5XLBIgfHxvsnXFJ9JBcuVtErQ8vL0X43dn1Elr68qg1
1xqWd15IGhdEjc3mMoJR4fJjFO1r0xXzHgbjLE645Xi5xQm5b8VxmivvF5iXHH0RYQpnkH0/hK0Z
hKOXMAhqHmMlRM+DEpvLyuQY4lvd6ARIIvLuZBCkwpKUOGEuNYY0wNv9m/GeURx7pq0PBSU6S3f8
/ifGxdxF8b3BrQ+68dqIuxWv0EidduOVmy11tuDM4SAbUJta9El6AfjpnFSmHPHw6DZZ70gJPgYY
4bF8+hD4G1fS++txfHb22iVoYiOxisHqN81DOE/2dj948W9+fulx9+0EEFoh5bKh2qTvS5z/YgrK
RcAkDNxCqvVYRgf+aR+2libmyIAqyqfI+R8ct6HdCTacGPNqyMDEmC+5gLOmlI3ZWYzkWI3JvRpv
nqo2II/u/39lfhXagjPnbgvDsgs1keR/JoS4ul3GZuDHBjWqUJ/0vr9laGoBQZ3w58JYjlF3u7mR
epCs7MMPr9KyFWNPrETp+Qrn4axjX58yF2n4mbe3Lo7fAtueUZgJtHvQZujGz7Rrf3ZKifh4Qx6j
tXqc8VvZ+sj7CoKhJy6+FHrMDiiYrroZvV06jFH5ZsXI1X0+j8/bASODJeoHAy9Ptgq06JZpOP5M
kU/2aKgxMuNaxemFdY5bX9hmYonRvr6jrIHdHhv51/Hjg/84Quu7GPqw+NMd8sSJKRnv7DndWUuL
bs+4wAircxaO1rbqSWYPzMYQoHHxNRwXsXtUIaYXK1aaBUmOmtRYRHU0uAgadYnnwgwSc+rRDGOx
ULgapak1eY9ts8EaNn0xqqPabxvvxLrGMbhx5v1SMeZ0+YR5FFdr50yflx5UtT0Ljo1Cy9gWzGZ2
rAWZIXUEuzhSj+oFaKj6y4GwKANhsSqAUm7DdCY3yGzHapyZFIpRolz9BFF9BlKs4tJGYQZ+cy+R
UNMCT0V96VDQenzfZmM1zMSXab64hmq7X334YnyN7BOG0CMacU619AT+V2ehBF9yU5q6BP96i5Nl
k7ucjm+2XiayiaFk7EB7rpLRBC1X19WbG86eVgn7ImLd0eZHZV8xFgHeEuz2WtXzi4rY1SUMpAUL
w/L1bsnNzyF6XiHtcATPV0FSsjbARBMpOdNXM5V8GIPMQPKgGqWVKQeHWaZKqiPKfNlNZcYIFq6r
5hLF9OL/9zQhfzZPHEVr+ZJyOwyajNIs8Bu2IH6rqbUcALWnWfWrs6ZhL4Cn7Uaq02P75QL54PA5
hgktZSH0xkrLjb9GwO/4zagB9moxLDurQvDwND0Cm/qtWX6pkH+8Qr5uqimHdBsuixJCYkm9fkcd
xCYKjqaJNq/MnEcSAeZrKWs10dptBeBx63z7YmDDM/UFnqhUbew7KE8EOEUDFn1djSLl7x8nBCg3
nkjmI7SNH2agJID93ESswUPbZxtx6cNLMDeVDsKosY3sguGNWwTP2TrnrtNbpRj3alBwzrbj0xGN
wuIBMrAL+KeJF5am4cgbG7WSOAW8RsphgA5jtYtw2CZiRajZc17ciRysbJRZuJWPpRlec9xxcOSh
uO3lXKiGDO0Tf+H6RCMuJCKPIiMz58udhf0CgvHdQxOpc0ZIE3xcnTgtdcrTRnop4lVre+j6TqM5
2++AQKhYRJmHk3wPBNzd6xsg4vvBfUWpucpzmbA5rxvL0WfNlH3s5EJuhavj0443cQDoMtnPFyZB
lKv5hVYiZZ9kfSxo08Spp7PUkH9rQHKh9cRGxwGeEwzIb6BWRQ1e75TN2F4SwrrVn1Oh71Zkx9zj
tSf0Xq24ygj6EYBWRG2dncpM+HuxxRcKdra1N6l4zsKokiSGv95f739S8dEcfS/b2Rth81u0Nz1f
fGgjM00ZB5HUmcCkYjK2j/NrssQkBydt3cM9InlnVhdN6C1twRe90AxadNm5bmUGoio+NoWZmCgW
sRboH9S1wXvkdpN2wN56f5iUad4b4a6e6VmauCBX++BdrhJ7kiZMqvsO+ZbP8nC+AJ5Iv6l49y4X
Q83K9BlLLmVkTaL/RTee35mckbAW+42GrAEef2aFFta2r2Y7Pkm6dBBPZjBYoEFgNEUldaHCNo7c
WzWf7JqsC5uLudg/uZnp8/wKVJ7ZCUxMIvHiK/IqeGOi/N7XsYxlXPCqs2cWW/c98treijHK0FBA
G7YUSic2c9DNziKXsWML8TSvELbZv1lWW0wiQsSte3Fhsy2WZHMNSHoD/5/8vlrM6hIli033sTfl
ncsC+GwAIGmwOi6v+ws9Hdz3048uCxgj4SAk3OkrLrFcbBGqpQM2oeJI3tWqlfuinp3jhDfVNmi0
VHyrCQJqkwuDuF38eCApXGJH8oKp7ieK+nobq9NRYBp/JCzbSOLHFWu1iG1n4yrHhCvf1OzakPm3
7RV4kBlOFIZvaLpiSnuLPXhFtQSJvOYml2qFVyztJPcIao0vaAlPsWdOqVdgZUCKl1C1lYhd15iU
r30qFKAUCHHr/5kGJ1uhAEq46MuHPC5DYZm/A0jdRpUd64ZXLgCGhO92WFc4vQWptaYPX9BQuCvn
KsTUS4GLkvQlcaTgUY7WIDtotlo/f0TQhv8ubeCjofHEXvZ6sYDAG+aeXJyu8HOFd5NuilwVsyR8
ip6Z45XZc76uiilBxMFQQODrqw+zgR37nOs2bhrYed6Ppd8uwX9HW65dD5RLkTiKAb15yiZA2M38
BTN3iPyyVpmEG9HpUplCSHNakfAHp8b/zZUKO7R4VQGe2lOCMVphucgeW+7tfLSbKtg/kfEbQIoP
L7xO14FzpW//KYF3ucf5p9K/IHPfL5vHMEveQAAVGhgjx0Rt51isWuTE7O/RZUIymp/0hnIrnvNo
4/jhhsPOCrjaHUblT4gOllYkroNr4E6heMeEMvmcMaZIIAg/emx0Uz/fzpFvIFNd29EHNnmFEQee
F68Z6R+7dbwQTa0L8RqHYHXygd/CcOAQ79IL9Ii4g6bMpWy9tPppTJ8VOxWha1HNfAwLcrZxZQex
R7Z/bV4POxzerufs5+vPyetAU/ajZw3N3cuZA7stJYLyiwapkNLnqC4AOOmrl3ol4CBF7TJFzE+U
9jYUvwJ8GilJumglSPVA4xw+DymX6Q34EW47/ijuu6QWyV99G2tRKKuvmZ+3dnwneLLfdtxfCYDM
OxgMXY/sFOmjVxtpTgVVwa3BNWkg1ox6Fp5Xliinl5WHZzg+fWAk90q970T4CAAQ+Mabm9NN0Ydc
dAF7Fa9W1XI5WueEw45ctpdLT+h0odSl5Qel+7P/aFksX9abyISPrEJdMPh//9b0RT/DW7zXmybq
xDzpfa+4rUtTqLFDiSS5en7kZDtm9Q+aoUCDMsn5q1wbintLotUYt/57erfPEqJUIYKSx1rXPRpj
l+DshQfnu+c8e5PSpjlqw8pxoA7/5O8sgOF/Sv5v2XthcSS5UlzGdlm3EZmX677ZMyaSGthN/Kva
ncca71bwNpZRt+TaeQmOwEVCqlUoY/jSNc6372I2VMpPYnTzADCfvI6lP3PIlVqVeaACFjekpPnH
h9RiTTG/nIP9nlG/Znk074HWDCEXDlBZJ+vNog+wAnA9Vvg/DWXFxgieX7nxYvYw66P0ybv5z9uP
skHnEzBsBAqgSI4Sdd5dpWgFCF+a8AQrT3O3DHfTc/alSn8wB8Ts6WMUTwIxU0Q6MAEoAS0+p1ir
Fv2IdhGNY5sp7FlMERHk4QNlWTFxZrgONS1ODyVr0/mXFqaeu3helNxCr3FsofW2KFxtDJlBynPR
No698z4+oBNjKMDttX1IPP+DTSMSWEaWv/jX1AZwDsPAYcQRE/J+kCXG0pAAWWQxlvS8
`protect end_protected

