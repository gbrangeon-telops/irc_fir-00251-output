

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FAkw7gRmEwDx0cT0lLfFXgH94E+u7pXWs5ahSt/pzljIAtlVd5PhOu9ztNGUELVfoO4Gol+zPLUh
TN9yRctY4Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OsI56UKE4Z4O4++RpLw+Gr7y1Sd3eUkdDGmGZYBu0aWjoj+iDwzKGBcBG0rF5D+4LwCAgnpAGiys
xLyYTz/ObATK7L0zNe+Mx/H+/j5j5SXpNvpcXkGCWx3Mtg6EpqxneRyrD34svh6fn9QBg9AkFvdb
eTcam3dZU+Gacfm2Ivg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qc1VB803xD7sVBXVT5KuCy+daGAjeSNtMgViDKH2bpJoW4aexvjdVOFa9Cn3ZQUudsfzbRtbOfND
3qwRkfwGKGa/rWJp/b4u168LG7R497q3mKgxz4wZrw5VVWth06zATVCPkvVwwcP1aVCYV0wxe3+F
BcZo/LoE5dzRftELWM1hbxUlZMlSl/apI9c5DLD1ZPtssPXqyfH8yGBCJ6IwpqThHkCcKlxPWOFY
XBErOYYrcO+fou4DBovYWIgQB0ZKOhCR4cvN3q6rg5XOYT99xP70Y8jdZqXKRq3PuDDZEya4uwav
9zgp9xA7sRjUN5/fcIvFMcfDutvNPIc7IvkzWQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xeydwtnivo2IBZhciZFfy3r1qoKk43zuwlyfDAWr7E6QmSwqVQF5VHmc7oNu8/L6oqsi8CW2guof
n3LQZ6J8fPLN7CBNStOEImWoOU09vnECk8Bwe5gJEo2CSwnqojJJlM/jtH5jKtWnMb5YecjpsAkT
3bnS2U0oIgAvNLFItdk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QglgmN/aSMz0M17AlWb9oRKStkdBh5nVOwe4/WnjlbCHuTNXWcMIzqLlv5JcAmIdzL/13EAMS4W+
LbXaFXFMcWHAzC/5AZxX+CZbwE46qfB6uGUmUBTFEckk+Ba1aO38uKX6EDual9TqDkiz6OPrjmC5
MifvdDzh7mlaB+rYqb5sjxUWUfJCpXIOgO6lavL3535AS2e2hAYpmi1PB/ejGTuva2r1NRmDkiUk
Uq0oiyBI4sQwmU7gFF9pADJRyzpgRQuSICfI5NAGRTR3by64/5TeOArBdjuY9arezL4gMGXoOIu4
E5vrAQOLZikLF7X3/wpaihrUarYdJnuPPVXNaA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 48992)
`protect data_block
Edpm4EfN7BdHb/yaj1XEqcJOAo4F6QcJgfN7G5O2dnO143Hw9iGB+GLBQ5EJ9QPLATPn9LedWCwT
Qbg2CkOXvmAkVxb/CAs63obiqOpnRFu/gPxnv16D5By+QDZZq+QaZ9iV3nWidl5xvBFXiPhwwYsh
SlHIzSVhZjEy7lcxJIbhj7CAU2cOx9Ar9Yh2vC2sgjtlAUS/4GvRIriiyWWl0u3i4iC9brTQFSIg
0ZGq7ltUHvkHKL0LRKYhS0kfpZXDPiJhrEam2/EiIn7B7UIZ8y2CFpx/OUd/k4SSIzra2mY8F33b
wciAyolRpBdRBNKIVHJEaFtTjR0PcNy/ZgD1sUk5rylNTmNGA5iAWa27LcccVDnS4M87mNSmctGR
d5SoLqWZDP0KpwWa49kzozgpx7gx2KojXfQ9JSrd9xiUv9SI7Of8zIWDJwkZovXDYl9bcJmq/nJC
YBfpPhla8/y2HoIZyuRYwqMbqvKfF1DDWH94L4ditZ6jB2BMNb5XlrM0SUU5ZKSuk+PjiiF1LBh8
TgRHC6e6Lqx3eV7DoYhhYljXhiFbD7eYtOPErBVQH0n6AvvO4/u68blfT72VHfkrMjrtRgcv+Qzb
+PXJmz+12+mc295WMvd1J5y1o7lB9mBQPOvQ5OOvHxFSVRW0Ur29tMjKuM2GHuDAaglcjgKfCehF
zBNrnCKYlfrwxfW5p2aDiv2cQg5yFhcK3GvBkGWtTkcZ5+TXuKmnopGRm3vECL6JAjbNk1ImAG9b
CA4em7/jQQCjL9SKhiCD5Tdq7mNMXpKMEAjMhYwuc0X+vtsONR4UiRZpk4zsNRi7eoxO9TzqtUg/
XLDMahWqISrqV+IHNRdCBuXlwjl8h67yL0Q5nn/scD5W221rUReGI62JX7rBc+scIUnpqrMfBI41
Ohh49iVWdm/qhKTlf3eyOLRW4Ncy8guwVFc9e4EY/jEsX7W9LvHkoZNpbWta6f8MqEEQGaQCu3Ye
R+f5ea/zDdJniKQDq58lV/S//U1rXWX7vYxEodk6AcGkwOxjio2ff/+M+pvy7qTmUFYMbqlLKfzY
sKIEoMNf6ewynFEY4sIAVaXBXergdN0g4Izc/E/1gjPa9sHZ6AwHhU3uMCp6Az1C1ooYYECYmPSX
/Te7WJtgtGg/xSsgHDFcSF8YXwjs4ZtsELT5RySWwIDiDANQbboPbBA0B3RxDEFiyvoihce08Ib0
fc2E85sM9tWYa3wiUL0MpERZEiB8o7qzi7uqZsoch9oOm0FqtacnVrDYbRK3VP3ir2IJg1lPQaUE
N6YkRWusYFgs9u5SOuxt38obusQvB60TP3tCW7tCJYwPFaPXHMfudnur8zp6dzDnrpqtp4xj+zWw
QmJZmRdjxl1/cYtT4y0qVHS4dR9Sx5TFisdxMcDb3LLwF7/JLcFlfD0tmWk1D2QMLQU8vomyxv6A
9knBjm9OvxqBsBXRyPLSp/PtuH68ujtttFP+OQZCTnLKnRhs1njC7+tw1sx5oaVjAxls9TegaG8C
EopKsBdORzpFExAjS4NK6/ENqZ2JCsOAMsCN1ei2TNAKFfmE+/3TzeAtPe4zD7faSg6dlj0hsuTv
zHfqOk0bxLWmDX0i6pBAg+ngIYkdpE2746p0HzXDkoXnrjYPdsKNqAffUL4JwDdGIhFUHjlmK1gw
zFWkwwZAYdAQez6gW+GYvHOblg2wHN/6PgQKL9LHoCwAlEDAaWuXD5ApScLJHydYmCI2TnJsx7lZ
ya9ajCtXJFPUojO1rJBhR1Be2xSaE5kjTWqBDndW5VnJNeBktKMeW4r9LxS13DRGFXCy5v/YS3Pl
vivYv0L4mTbadopQMcOCZNcQIutjlRlGA/illUDNW+2kidXO7q8p6+SIVLpKLNZQyXFgYSJy9/Px
Q6iJrfcF8LR9m5Tgxt0bwxmizzTm4TJ2D6PmSgQszUezihGz9w5RM+gid2sUqq1eqTQoc4nMVMTK
cQteE0Ph/JHRDQTkPV4OWDtByb0dNFrc6WcSHDgPbXaCUKA/XY4xrtuzvf6YvQl31g91nF/sqXqV
Ko1ToBKWcZTD3mRzDOH7tb+O0UhiR4tXLFVlXZTu04/6xCPHclbu0QSIp132kJ5E/YB+lUlRPfq3
rHFsQQiGg35ZkNUsxnOB/ZozSRiztb/78W3qWRaId+fYb5ZHJlHYfWLxNtb27Aab5SOLlCb0LXbJ
75oUxFqbJFOEB0Rhf+fTteAfOAeM713MtpGhBOatbA5tEBGJY+Vxs16Mp2Vv5I0HuPS3I9umlRjq
oWDu1ArDauY5dVMFDmXwcSWVRcOUfYGvbBJQUzGdfW3cu8diVch5ck8Qqoazm13u/sMhctYZla2P
rpAsKhCvls7zw9t+Z9GVJueluz8IA+SXF3I+MKvoiqJAx2KIPpR3mgkNdJbTBzGPpRLrBer+6D1u
vaFZe0J6p5iSLhmE2gbfv5RYmQ+bGBPfNccMyFO9rPmVUeFKu9oV2wyBsSgeCU8YrxMMHJmwwn3g
yEi4NX8CkwAnIyv+qZ0sP1wg2VhW7ldeteZI2wvsZ8FnDlU20NEmaw6+X95eVEDAP8/XZNcrcR+j
r5St5mSCjGmlVtRd5UdpDSV05r+HPGIWEKHs2s0UpUN2iOWUxbPmmfQuUmS7q4rXDnSAGz0TJ1vU
W7MzNgmHCgjLlL/+1p80mK0x5kHlVn5M+4KB7ZIfPuDmcqBh2ToTLaJCqwZdZOYsarUPnoES6Atu
ISDjnK9big4KNzgs/FTOFNRSE1kZNXFMFXplWl0lrb1Q2yxNlUwKy9uELOGzbFHtTuJJ8Jf85sYi
UFZLZYYLDEeWk/Sxi1xfLedwYMdTDTNs953j2pJ9fL25TheghvT7r+//KQVtfAfqJqUVb94sgoEX
rc6ahyYCwmTgtyVKeDkcvDE6Xju8Lmygbu9s0GWcsL+XtnIci4ZzYOe1ZE5VU8pPh+Ni8gALTuVc
7fyLbWU0/ISBpLp89ISvcZudYBEsNx9as22nbEM+0pUXoRzCvfBhG1SQhi/xGDnzhVcYmRZ5+Zzk
5h5/WGg6SOPhC+EFUpCPNn9lcUSytoGIKY+3UyfB989BXa7hrlt1JI3FpYJ8JrELoOHj2heuMlJ/
cTHtaMjdEIp6KoWwcsON0AN09J2eK6n/UuluiJuE2eZVC48VCgANhuGuwJeYiBttBuacreV4WZZ+
kAV9POLQUmVj9DxFk7PW0nBcKwbrnn4at1YDTlFFem/52kyRhNAf3IxNuLQE2tXD0X8smVdDtv22
xqjhmxCoawHD/TmpCEtes29Vv++4dNJz2VfpVicwjKB32HqvZbmyxdgO0uyert7RzQXz17KXskYU
KQJXmRX1RHmOxKY4SUVC8a0aTveTjGUC7/2YEYs947+9SiFwTqc7lgwdsp72m+MPR+uw9Lejs87D
EafAIAXVs6Y8Z79lFP4UG+Rc9a5f03W9pPN72QeqT+fbe0UhHxTopFdhXn0H36p+/M6O9S/FOLfR
WfKQy9WeAXMOjpovaMQwqD6WxMx4g1JtFoYnjbi/2AtRhHNP6ooDsBXwEhN4Xy8ETfjP8AlHfVLK
Psw3P1DOeJkb2MF+Ds+Re+AX1KBkLuqUBeniqsqiBup8Qh/YSr4ji93Hz+I7OZYshsf2aSkpu2kH
K3a1XYKcDAWpztc8XlpowvRNWoxI+OxAJEoWCW++9fys4oMbRom2msI6sS5l8LhV028BthbJvLK3
bTTWctHjePKhC+m5t690e2qKO0FIDHQK1Ler8tdb26VA5dZ7rDx/mFeGoR3SNYob76KyqfoK44Ri
LH1UIM0dm/K0KNV99HJ89Z2jlb3n9CEgHY5wKP5mhqCEsY+P73c3+5qb4GNynQUAxQf74BEvGZVg
w+HHYfw6ZyfKdSGMktf5glLu8ki2Sur83gqiXhdR265PagSI6S+qq90rJYrirT+Ry7qtq0DwsQrO
bN1E1uO7OY4HtrW9EF7sRcwbdxP0xWA8r8HR1WRVMI8wrwpQdVZZsyz4XCjaxiBzhMlgt9jkc93B
9Ldr/x5DSsnbX+qM71itCduQnVVFyxehD6Cp007LN64cEp5610+FevrbG8PMWr0Duzwt5YNHu/B7
f8lGy5LC9cm8pGEuceKAPsp0kMzWwveoiZyRrRR/OqZ7nbgJGf6PK2DDF/yeJ7uqjnw3JddKw4Aw
V2XRmEOWgyBUQOUZCun2TLY6/3m65FHh4557wyiyn1ZJm4rln+PIz/cfJcEKU1387WAM6nRJY+DB
qR+wQRIVBD5epRrvjdYyb98YGA+uOR6p2BZd8sS07h/CtFARuFioz2t1N+C4+1sieI0H0Yvqd1EI
VXoN+tw1c4BpE/LX0vr/vhvCWA/tDKoDGaX26ReS3FpydROGltQPk1DIMKEFfxA/RKLkLgYZwS/G
2YJm286+lQ638x6TrRbk/WTRYwJKRvwNWphuVPOOTf9SddhGzncNZEHLeoy2FfkBKeQ6KUwL1qY7
ABEtO3RaJiiLJtJVr2FDNcOYNJHXSH+IwQ6yctVO91Lq9Mq0oRwKXk0uonSkks+IHfqX34mjxaTk
SQl+eK2sWR/5M0FK5ihtJMlezhHIHDctAwhHiUtO5LvS2GaCcoYUFUzJmFdvp6IwLMayWGF5FvLa
u80v/NwuytZt/6KRQJ5+hMqwveLNsd2H+0p6ZbiyHiUrQE8N1OCysiKYwJYobCuT1bYXKedtSVov
n1R5zMWBeQfOnNKQ0gAyaHy2Wn0Ex7eaekAYyTI8xcEraGgzAMYkd4VB+W48Bfb4k8Yg097Upnco
Atl3fvyr3Xhpwlo5DXDhgMTvFbX20C029Y7vVO9IKXyj/h/kwnPRe60VPTg+vA5cc7rUEjpSUlAt
bWPZiTr7TLPWKqwYebjDQ7G4SDKj9/Oijs/CXz93XVydqm2B7QASlApN7hWpaCk0B1ORV7SKsCGJ
ZKATORwvK7FDDvldC09hRt6DxyJehGYKTOX6Ev9E1/w08GxYTyexxiTSMIXL3b5hdxfI1f1JCbIA
6bvI9esvdtVLUIvD9okJMZf4SD43PK505OBBardfgZ2qIk4u5Y3kcNZl6JB9SipkUFSBHvIQjOaP
uzi/iBG8vQnaRmM43h03Ixi4k835kR8mghID7RCzcdiC5N/f39Y7Wu5Z/nvOC9g5/Yig5E3w5xts
nwbNcF9yIdNc1zsG1/qO7joE22T5u9eq6sw2EjXdYuPnoM5kzyqAtmxtgeGm+/nJ06tyo/1u07Zu
e7TDbGISoRA/z/AAi4WEmgIWz/BW35Q5AVOEXzn9kSyLvyy98TmPUWdMNn0ArZXqdsoe7qrwruvp
VTpxo0angYED0PK2zGixG7VPN6pI+rOvp2zlUojBhWQJRiJg88EzAhHkyraKtCS6rM3rrOApG1eM
Wv/JtPjpFIuB9Kuy5ofkbMxBgpS8CJS3HpzV1QJfcAhio+D/fimxYKzNDBZgb9DFFT+o3SjFRCoq
5M5o7FIwm4HsAoWozAAJuXaeXgJewBduRhBud/AD3g3OIuqUTYuA05B3bjfnInbTwQ7Y6kCPTbP8
Arjz7au+Uyb009k2Z+MvXtvyDQ2KbCTPJo/EVIlcDZT5BIPRJEKbO40kHlOQj91zTli4sNApBRTB
A/0I5K6TusN8tAuqPx9rtuQlyTk8Lducj8IYlUpfcJIPWeyHfWBjqEaygDoNItkLRIdq1RtsLp5N
BSEL+SYMDTLFgDNFzIZBWy89JuNXDxitv964s1ehlEge95KoKVb96ZitkPaGlopCm90Vu/+gSFLx
8dbEyfPgWg2baM32J8u+slCW/o8nqXrFsIPWjmwSU9ByL1VnevK5yBsE6eHam/5+sE/t9d4Jcgnr
Fzcod2f57dU8mN+r28Xh4yIqVFGv2cKCMylz+gq52P9RWjsckfS2Wa3UoAjisdgb1BolUq6z+nHl
iQAZOr2l0IVP85SLWsPoym3zgxjEYM3igvnkySNj30NuNIymlMIRZuZZktH1lAGVmAjclTqFDksa
my4FqimSxfrVpci9wXCTLlKpXISiUdkBlsavgs4uYg9PhwZ5kL4dcCEWWFiaP1GuFipPwCoSUajw
jClkhO6/4YOzzZ1v0Frfs55VcyjipJQmhJyld2UjeukPojBUJDxylUboLlApme36mkYdz5mnrU7N
vBz5ZDAkGQutvg/gVPpL68ZX4F+pr0Q3OIK74lnsuno42pSJlJuikHY4+LefB61akMXxAf0Hp3p2
R/e0EigiiACMqbP9wwZyUlkHohGMoQBr5Obo8UFEbq0Iw82yYVi6FBvRHDi89RoswiT5oNgLuIVt
ExQlvMlpTMmYjHHbMoH3LRULYBBGJpob/dSR7jy/a1zPXsTCnoxmCGnBkEXzsdnDowJSl/HPodpZ
g6NwEpgRlyPXRGm6zGUyg3fAzdeiSQiZvzYT7+aLZ5B9du+YocPXv4ywaqnAFxgLHN18jeb2Obha
8uCgSJbfdc8//jNZKxIsw527OfqcjrF47qNZlg+SkhB94nIB+Ri+spigH1M2RJ0qmDCnqc7jdOkh
4lhKiFe5039wZ+X09nrA64gKRbLcxJot6jXwmzPXQjG6lWH7njcoR7fgJMOIb2idAI23rPkjn6sQ
LNUjojPIXweMobPPXZzChi3vJTFNpUZ42CnRL2Vo2SaRSekuKI5l7b6ePvYLOj6yx9G18r52KU8Y
XOnK3IWKo75Y7WQ/+4INZFAR67l8TURTHH14rkhu05sM0Zcf0N6LMa57AM3FiJjODxVkDQBEVMQB
UZWN3FQh4t+GcfZ0Sl3HBjDKu3b3tW6DYUsE3MJfHDfkUyBmK/PQv/AvtRYkC14ifT0D8zlAuiq0
L4Bc2q9aQMxDWq+D+rWQPf6p8caFlM/dqpN73wuvTXziOimUfnGwjybb4zR6hM27hVC5NJg15sCk
6elz+xMH7MGqj9LkAzqjGLVnwt6IG2Ho4IYx6utwtnFEbDuFuiQoTSOaBFA6KDVAp4tKVFBO3/5F
FUUnDMdLmlmFXFRtU+4zFnRxAEss9CQ0xIuHtPSdNS4oOcVBNDJ6HJviXLSzZbnMO9TQDYph5/5Z
LRWHjbVjOUZAFJymQk8qXM3lTvUM86wxZQIkH3M3la0Vwka/7VkhZZ9hQAh3OBQ6w/QryY8VgMAS
kdRCw4nQFT7UG7snQzSS/ryOdYcb2CV7PT7HUfIzfyHqgCEY0Q9wavCevt2IuSBXQxOFBg0F62C2
aKY5/RpiDHrD/0ybiLS3XxwksXU7or87ou3FEp6YTRm4IbpIN6Iv5QrO0HxZcRRXb1s2UgjruGfl
lh3idnHanE/G7W/WKgWVvKuLffiMW7ZI4sagay/UxFADB5Urt7ckIHc5ka5ojbewfrBYe1hF8I+Z
3QD4AmHgd4NB9I0cVVTWYgQ4G5Ol5vJkflNgqik6YS0zyCCPDyM4ouDsWrIzJyrvMcviTQKefoBE
uLTAQVtqwSXEeErYkJpTQWfhm/f9JaDHa42NT8MESlHYHS6RWq6DNkQRah6dtmYdur6TIUfXjHdQ
YZfpUe3NWyMB0Mo7Vek7eRUOgsIPOpEwEOIgZDfsJBdvkzL5s4k3RffrggeakwYCVJ7Rfzj8AuEk
YGnGO4x2Hteo5AT4hCH0+SPLHFfYOhscYEwAHLpoJSk9oDCF7IKm1mssQ1hZBYJ5dsuemmVUQ+Ge
n6Eoc7DXuiXK2vq4EqDuqNO9y0pCzSJvpA7Zxol3Mw+F+V9qnX0Z5q8M5XrMl2JLno6HU0qlf+WD
r9qTgkm54PYymSRoFpxs/znzKYpLmNTOjpS6YT0inz3n3DogLtx2orN+mIwPN0Eda1rNKxJMiI+A
icbEAM1CQqVIzfM/XTebblHcyUoa3e4M+BrWSJubOnMbhveAOOquR2zpHpdh5FsPAGDLZXPnr9qH
JFQVEkioNEaoCp2oR8ZAaFg85r+Oq+kfBxoufvd7IyrklMBaSZxKMNPe74BBLElR13xFu1bukvEX
bVias2eiGPgrfvkEU8cXxsQYvSgOeAdTyU4QK7UpbhgSlOd76W2X2ykTa+ZfvvsbwxqlsVJjbbN8
m8sXetFIjkKdsETg76dFcAnYrVrxWOaaCu8hxHW/JvuAH3dTW1pn+2zSvmBnJnABh0jw6+tJW+GS
16C8I+iOyMhcYNf09WWsrQ64gqGXyuadpPMsOnf1x9M0U3EhnVB4nNDYsQh2KDjJKcmUboI7SyBV
6DBdChtCXQDyswexpdfD1THZAKgB9nACg1n+kOuX2/9Nealz44GCROvAcvDzCQRmnE59LCofzptt
3HhTlv9T2Psp86iQ6/nzTyx6FuLsRn4HJQ8EkisLORrJ5FtVwtSMYm3ZqsizAbOPwLTnE9e/Tkbg
W041Xagd6PZIrF53srdRs/pWf8Bv7HpHaAOk7WVcbB9CU2RhIKZ+Bai/D2CXfyLvgHyuYnXMh2kk
reBwSrt9kw/BoOgK7axkzTZd0tZovTAS6+z94PKNezY/LXnIOWp7LhCAvyy3U52RCu+RxFjDLOAq
Yrt0sCQnQNb8kBkwABRhzpEIaGqmd2ivmb2dBHrbJ6l17cceQqpzmWqNiY15bkAjWXPrbbfi4KCE
csEVeTVXQer/8IlqvS3NFm/SnaWiRIvLmDAqy82Z0kOS6/zw1pq0cnd2CGt7EUrIS0EuCltEdX74
eROPxUi5nxS6h7X7MRQou+AjbJRRIuxxdB5Xx5VVVFk8HiZtB+9DzCchvGR/8yRZJm+NaWWUi4oX
mIwPqzOr8lyLyAiHgvxz9nfJqGdXml8/koDCiT4nx5VvBeQGoYLELlYFQEXA0sW/mXk4Xi5qM+sf
VNM2GrsAZu32Y4iABVnK4xEyCb4Ge8A0SDcCHCwFqlxDrJUKL4WstQwDqsyaldDzh0L9ExTtoHJa
iuuBAsWnejfDcmI7XSPbdxCsirdWccF8JmHXEXmzoe/SKIY21Sn3+aL4/Blgw6aLWD9mIcNshSwa
//Qy4U0BebTWhDY7yQMMPng9A5KFB38mYLVwLbnEkZ3mzUGAFgUPjCy9bBynCw0K+i0mJaMH2JWn
BJ3ntuMuxrkJ7Qn2PqihlIuO4QzNaK0SmxfUaq8kblNEniBY0BphVYSmJGA8z4jMW0g2bTmD6SQo
MLdfKtfpZfoMJsqc9bAF4W3zKbHpL10O1N/IeKCWOvQwaSFEhUwKRCead64PMOXk93JILCCbAduq
g4i/5jFbVfaackulSzCyRna3St0wOmzM+SugxZfMm5yKm2cXGHYgdWkjuklqBSrdjq2Yjxd0u+9m
5AKcV6+s8EUVE8ZImvnQYujl4NEyWURKfK2y1MNkxAHngo8kWPxoCTfGxBYipP1CEJOZHh9tHAb8
C+Z7oQaN/JDpe/vA/gR8ohu+1+t1t4qw0U7vo2z/3ZMc/8cJqZL/+48u0Ksla5TXJZF9ybDHVr/W
K2usnitMp+tvY8YL40jF4IzdBa4jPCewak7lxmiT50/3neW0JRH8nodSH5xoGoKUNhHqipZyhldv
XQ+qmM+HjiFFIXN0Kfj98VSgEJ8gWoMLn0xAFkSuDbTw77zLNu+z2+wZtW9Suavv2NwNk6dcbPb/
jhO3y3S0eSvN4OaJpIiijoWW9h3CLmPa0ZXdh+HbZLnGzh4G8/XwWdSyOXEmF5rmebd/vk1l8F8o
4rIL2LeU7eZFY/b+njw6dU2McQgVqJyyW4LZdhkQ3wHHJfYlBN7ER+qPZeIvRtGcK9UR9YEtEfVx
z6Nj/vdoJyMKp0p/o4+fF5vNNn/eLKJGAH7QvzcIOle2vvxsKUkAJX0raRIOtAXtuKtxfu45/dO3
J3a5ItCSkVPtXf01UEYzhB45FxFIqwQTia59sDBtyQ//lzzPb+db7kMDUhRzNR+bDCsKSwWD8a3w
xoIIdCJ36u7lTdICcOEI18SZQvqZ14s49fvK4bP6jhT4zlRt6XnX4DXBAdCZR+7ICTs+KqY24iMg
gh0bp548N2K/fjtL0XWSjxtp7FBx9rks3iYxtphRTeC8YgToNeBsWZOltRsDYw1afDYwVooJ2VyO
4hN0nyheTJNPhcSCacq3oUojxUVV7KOv80yn7Ao/Zdo4ckhvnFTUXr+dqEh2XPeSz9/r+2b/TnxK
H4RFNSRlEH2yMDnqau/TkU4bxR8lrywxEm5OaK2F6ySibWh7OcV8FMnpFpaQktba3XdVTdC0RhEV
5FzlmBhEvCCC0oNZIG+mOByFArXdQpvItTM47/v/epELb8irrUGGyrxMvL375aAA+zUY59xdJD/l
WjTKSG3hfPc7Hm1mKt03H5xT9SVZfhzeDm8PR8ghRN6qK9ORJ5zwV0LuaioeK6XkfGQwmu63Teb9
0cXnd3FQElTL99cBm51HpSNIRzH/uPbRbTkYfQNSsxLBNmmxLCjPJ30tlOFsVDMABNrTjYOSZ8hN
JPjKH1DvYJthV3ZsGjkRC/NcUxB4uywzeTsyLTvoC6M07UEeO80a0fIxdcuqADKU6YTEVNvRO8/i
oVZ8E9C23nNucBCCBEKXd2NKduOUargOmpz5lj12BbMwdpTAShdRsKGhRSgskjRJya2PG/0QK+Z4
FWqDg4n3wdxhtxbeC/YvqzLJD0r6JXNbAJO3SKVxBuCB6kbe/cHxflOjxLimrbi1Rj66XeDgSvmY
CnkTW+4tpeR7LYWbHTovZUkgC+wvFUAhjBv1YDYdowbyEynREIQkeikZvEj7tt+hD1agAvv9ioGp
3F8YraMF3EQSCSF1qgZTLGx1RapYzvJ6oxfRxU+ni8KxB3evYNDOxwp0dNLpqE9uIleEDCCwXpnK
NmlTmGbpHBUbAi0tNlzMgWgwBv2i4ryNfz0e1AF6LZvuOs+6bl72JH9351wRTlpsZs/u9OcW85mb
WrsDpDlnkkDLyQmsio6+HWzxqjswSm84d37c5E5N3XM51oGZam5QQd/yoFgb8xGds0Y9Lpgjgf27
B8XtTb06G4O8OzIZTK1b5ipN5GljZ3HRaNjkjTmOGfDavjQ+8yH/ouTeA+aEhjouPRX2WOQgh25u
byaL3SO+kgj9tBHrGg+pwQz2QerNGpmQR+KMjNqDnkRQO52JXP9UCtdy+TyTLWe2M4nEMaBRz/bh
9EBhP8GSNNSjWrisNK1RbPKuIfPFOV5GgVkbGzHVsfs7cYP7jHyDZQEFIPoXzjLBJppiImImq/xN
J0QcwQrs/OUk8NmtCyifWXY6tQTm1a9zeSBzVR77VM6elrSmNMN0YcDUe4xbHexVoB6ir7ac9pee
lZlaRhoL+TTRxVYoC1604RW4ZjsO3se7BnUsmgMslUNTJswo1oPGGjipW1FYXz0t103UGjyIvMTe
VWWreFNvzDuFH3RuoZGS80VTowV58o8BFw/JrWmHTMOrBAukdJXnQ0cZ04xlrAoGyYB3YmCx7NN1
ZmYMWvfcg1cSeKUYrf7yr379d4A3B5B1guiXn1eLaqPa1JCuDBfn35amOlTXOdFjhdcRLcMS8LM9
lb8Tuc9L2A7IpXjQQjiVCdsOY5gSPig8wE/SuTSyVhUL4CCyTZBonf6Ln+DbdaFdMSRWJm/7XJrI
UMzsvSCaGZRFpvP09+C4NhjL996Dxu4Pn3fsrY0bW87hpd43lrRYwyVocJPi49DS7oX/+ZOw1pQg
UgqyylDfJ+HoMqXin/Qv4EjQKKZScsRmsOdiEdoIlv7WCP9KavuhfjvW++LqvTzuXgssH1ete7zK
W3HTN9Fr4G/fz/elr+ZLRMK95StdPzc0IzSLp24jbhfGrrCebCkJZVCXpRYgGooTja94OYkpH155
hmxOuSz8e2kUrFswJmOoOfT3D95zuVe0HkKqoagV/+ZyK2f+s5BbjglhNsDTjQ8IJ6pabNdY7nZa
tN/81P8CXSWm5qy8/xB96lqooLGexMdoZ4ETAy4v2lfxkL8nSyIj3hSS3AH+5BMjdd9T7QNz0XGI
L4yjz62gGzV0uBAaC2OrxSG2Neupts+Cjkjw7hrDz9PPAPv+jCbnxDb9bjzbSuCEAvkv8IqfPzMP
AN4c2u9yhquZOAHQ+yLeG5zmfTymKWU2eEGmosQzgPHe1Md7pE/WsNfZh7NKSp7mGt0kR7trZ0Na
vZ2yOOvYDuIEUSUjPFQrl9vQZ98l+H6pEahlDkl2Wyl0cVnzjkVMznVym7EviNisBHJVdE9qFcGk
qsBGn0TFG3GFSa0EmOV7RDLl/IHINDlKDWTLDLE0qOroXkKj4FltPd/T2a+Z6uaDYR2q+hwnwn0Q
gA8uymnXv26rf9tle1EL0FsS6evbq6hX3onn7GbRrUQNF9IpqZEsj+Hr5v1/s75O5itkK4a2j2mJ
gsLv2D6Rio2iUZDsMFOWRuX9JGAHhVtQqdMJzWYIJ9fYjmjBSh9iw5jHa2L16iYSVIo6KGpvAsjT
wZCnLALiQn7mxsProWP+iM5f/WyFSU/+AAhm+myqwZVhHeOmb41HhN2DdA0xcDKv2YEYhoeOk8dF
oQ65U2UVjl6F70R0oKzNTRvkbgKCM9ul1oz8bUS9sZi3RkWjxEhIRg8+9bVxjQgoBnhGWJ90s4ez
PjH/jKfyxu013lAfvHIl8E7EOHyZ50zPlKbA6IV1stmYm57tRzghOcm2vPv3nNP03P48eg6+KGv4
KZ7qcx4SBwi/q1RGvs5J4cSlrXjcCrjMnHLG/k39fcgPCYaJpnYgk6yBevdQ/ebXUX0LGQK1XyHb
iA/JFwXEXTr0ajQ10zzn5Ecw7WPqkKMvvMh75hhUCG9OcokIURPfJFuUQBttp5ZcrVy/Tn/2QCB9
S515bDTYdc20fNU6bP3esHV/XHF0aVH6WFLqtzDER8ROOpjMRSztIt5huKLdnYAkp1OSBvgOm4p6
PUz4rFS6Luq+AgfZ+J7GFLLx1ZowkFFyz1NFlgeIWQ60IYYJ33iIKyYA/SxzmwC+i/s24Y75XqLn
/1YPr3EQPjdce273Ad7h/KJyiY1j3pk3p/od5YeBvtXgTDBAeaU8cSLqVhQiw+sYj/RntWGWP5Ne
nWkzKgBV3psl6lWLnGyZfr/GHvl9HlpLxJz5BcCQWBv/hRqoXNZ0ovxSQDmdRC2lgN9MdFRcXZ75
P/QUIX1HcQyz9INIWhbAgL2Fxm0jbEzPN4CyzcATSs9uqG3TOio/pw0aRUIbOdA7asoGkqV8LV7B
g+XWyZTWi4mva9U/us3tRm9fkufM6+F3un++OQV/wHQGLoBmksaka8G4tQPHSieaVVVAG6ea/4ip
U/2tLWVTUWlD53eDnqvbdjldjzmObitEJPRrFy9ShZf0Z4v/2UZJMZ/BHGT9baYKUjv13vePQ22J
xK5MSy+tDL8WXyeqlazFsTNajwzpNsjZwuVQeDLfrkoUHwWPhJRLxzAHQlOxghPrnTbbWcqX8fMH
taCJTItFbFvMldYwuDV5NVCXjZwIMKMSU+Mh8HUsk+6suPeDisoD1WOdq7A2tA3Mg5ZAc+QgZ303
NTDXP5s2wFqV4E0cQtLmvNfzkxFU6kJNtjpUBAvigZQKH8dgeVl/U4wF2yXsbHnRZan7hW3eWRf4
pvd5Q8cbDdHp0yQjgcG08DDo54w48MXdJWRvCRGAK9jaeCJustL1E66srURGwhD98Qku5Y+df1uj
b3WRd7MEtDTeFyJbxqnTC14U9o/X6xL9Eg6/kJG8OrZxRUOBE1FleDnZq8pTp/DTbh2wTmjxhQYN
k8lfIu5sUeWIcQVMRmzTpqdvVlIb9Mlirrrhi8O4emQQ/wBanA9QlaLRKReuOLrmxAcRj3wPM3l5
rSP9+O2ishvr9yoXLBtn32U9c7h6owreHTCIGTwIFe+8eHcwsnyKWrAYtuwN2SwM9j3QcHk1qNZg
JVXBDhtpNFzDvNiMD7r+8JFuCgjr7NPSu5tYVbSCOVYx4osgcVEwQb97s/77qEepaMunX5hW0gne
XVtV47EeR9XTlFDeeg05HQHHiMQZDx4yn+BbOPaE61ihctefFamuNw1MgM4jpUDBSS+U87C0Cl+N
ipK/yphW5xy1u46hLmtmRWUUL1QuVZ9eXTmBC7T7oGvl8UqHT/Wprb8CmyySsXopUP27NkwIUjPo
HX0syo8ikFiavxTBpvNYFf/qO+Sf4/u3+DaXgsENJnijpuOUmw4BeCMNjXJmwiaDytpd4tGqBMJU
G930QdbCtHsdmC8loquk8hJ1+EfUvp1ePZ4/fBAJcwt8mN8idRaD4KnVp0ovqzCVEk4eCKPnP7wn
H5ZrVb2GJNqnNrirEAvyxeiRdO+MNt3vJaGASrHQitulV8HCVjurvZrW3eSlqMb7jLs0LzBzmVSN
fagIFCrJB0kV1hJ7Gki0DFTqeIP8nkts4QeA6SnhqTxw1lLwXdZMzMuZjWP60ZLVugotKfDLd9BW
QEHGT+46f2RHUUnlMxyIxXWWGiiXrcNrOpGQTXZvDom9AzcEzVLEmpCemJUxA36rx8at+17KtWEn
bbmq5+sfTBg3xxfe0ICynYbgxGn7b2N5r1kE5Gu3OatA0dPN372dx8t4jvY9ILQQ2xX/gQo+SI6z
LIYNh9h6L64wgKsdMHlQjikBoWLaYTC+vpIpTMUO1wM+I2Q9wGJqks1XEEHoNazAO2053ta9U7/4
u0rhj9dPIPSEbAPJw2NrKj2p6qD9qFA6f+j97O2AFG2m4X8iQK8qH7DBLUmZ+cp6u1RVLscso0+R
8xKb2P9vbXh+QQTnF8jgY4FUpNK4P1dIYfcAVEj0HgBEj1pB5JTL5JJL4QK+EoVp8cpC9w7vSsQN
kwgI1f9Fop5Ppc5JNoqTcRP9qzxGULHj21J4f934twjSX38oBGldmIzTkJY995T2h7D+QLPXIi3Y
uJ25PO1MIts6b2xMnT6Z9QbfhdpPXzJla13UAjs+cuAm+no6lRBqCW/snBvUY4CTq/oTVt+WYWaz
YRNAZturEr3vUKQZ5jCPrmE1dFJLmWCZuBIPbK3juEpT7jeO2EBhY/tEwlSH65JbsF9H7UBXwbTs
3Rjes34mfCTSKvetwbr3vgeN4+O9Opwz7tdDPs2R10VjljPXazKDNktnXmwcyt4vH2lfhXO+RqTN
5qLIkTe6SzsZIiobAIUTRoa/flLHbnh/jcRlIc/7iPu0gcunPcyvU6i94/IodZ81LqGp6Yy1Z8ud
fP7QspeSIiHTs5ipipz0pdS6vvKCdt1UoL+27RV6wx64rVyME1++h58IftUO+hDLcXBeA184VfaV
f6d1B5Bmapq89P4kWDfk22aqyzhIYRozLiL4S8WPCMRZT1+zSk1F7hXzcRHAr4pS48UjYgbDlLTL
DokvKvx6UZ1mdwcPB99zZJRYFpgtdojFdErziwjn3xEAU2aqgOB9KgMl6nS4lLnsXtR98tTxaI5g
8SZxC2sDgtzh0ilF04A9SjiYuyq+71W6c/UHJ+tSMR7Yckr0mOGSggwMj4Ga+CB9RHR9D+PmQpM+
KVwCmd3+sR5m7s8B2gUvrWWpWEN1/qjvCmX+WRjxY4b3xa2aFvtSbmQNxeVMSXiNgLCY3KMm0Zup
WR/BvNMjukIGKWRH4OyHDjev56sWJw0BGiOk5EM3IxgZ8fsthOLrMYx+i5jS/Z5oFOV/67/R4bOX
KalF0FC5DTKG6L7Yiv+qQxwLbsk6pDQ2G/OAac9qvMb+fGLf9fLLvMMXv90xh8belAbhcadHW/um
x1SYhTTbjNG0hhqMZXGNLR/By+FsJnZ3+7Mt6sIcnlwb02vu6fqPkzg4McS7OUSzvYSkuqZOywKs
zqPfP0CctTuhMEtDcHghiD9W1qfrgmCdkPC61JWdLCBILS/eBQZDP0gwVB4lVnMVTUWYYMVyX0VH
w+PeS2fTJ05kwCtdq798pgwzAFvj19U8vY24+/wii2w6hxr+rrlETk4x7GSrCw7V1BmDiboB+gmT
nFbC959D5hZih6VGaYvvGLvYqSkcl2fObCAmKWvUzrKsWBicsRqBHhhVJL0BC2JWQkm7AO39ipLM
rivsldwJppbENe8WNB7PFE4rHwT5eMrDOjY5ZHhnoRir1OgtMlBJpBPGqrwEr381upV/XV41jAy5
Ej1yryw9IgMg09kKtrwtvTTW4Rekn9Y0LAHIl9QJiAerixUZbQ06qPbeo7y04dmbGS1IysCc+cWe
2Kd6N9auPKkYXeBK0jUGvO4+2wo1aXWdfxaHhUGJfRdeOR04eG8M0yD7KRhjapvS7YyiI2UPmiym
bicqtYGF+f1AvflWVTNBCi+GNvNvzWbqoforaGy3ziH1+6zJM28qlW/UKMFIYuXvpeUyhnx87Cys
Pl8+V3jYCtU/crZwzR1RnquKRPBCYt/ORGQECb4KSHx+dDufiohpeqc52KIFKnqNTH9co3iIGE/e
iNSYo7M7UJZ/WSbuOesAhk85WZ8gp5z6RXT9XIBeDqEqR8+AR5biamheGThVFlnkOG0CDU2XeP8b
5PYkwo4rzxwCYWIvVUAKEPrnhGhRsPs50ApdLwFpD8M0ASO0nkkLro3ZVdaftGIWlHOeJ6hjHBbc
25sXYJ7+V3HxXhP2Ig1jJlBfirrhvf28Gop3v+1WnP+vycSS6GBib5hAU+14NW+wCVeHxBcMHPS+
zpduUETVMOkvrjymzmEkI4BTOrPEj5Z7i83byg2XNzQtSjNx6aQeRerZOxgMwKxHyzaBNgv1F+8f
27pkAZ/Bz5+qw+Bo+UHL+R4aphDYpl/NPqgm6CS+a/bMEds2TDOY6cnGfmUO1x4oqZIWi4YjKTcL
Ah6L9rK04lrm04+PZ2/4LYAAeOxlCyvdjOSmZv+VifG3wiI6w10xDAaG47BYeD5L2uJwBt/YZjbG
Ut24NJL2ogIlKFIHKYjE9/mAHFbl04NdI1tHln/2Xf4aNyRIWos8Uq8RNM1RbcSwPqBm6pGzDNoG
DfCYsHSGXGObanvsFrbfJPCQ9KPxDzglXrTXxmK/MokSS1qUVkxVGCGnlMdPsCWPzKaRN5p4ANoc
CB6bsoSnpmISTMR3ttTM/l9zQ7nX3NV+WI2opA7FpZtmYNKK1iiQgsk05pP6yh7LMrvTfA1RUqHF
PoKWHRF3WmxgopUdI0yB6ZmcauMum+UuaPSr4y4sJ+10nMa2m9aaJc2dVVBfGSIJZ/TtBLyjobmf
QiJ0Vqk0iykCCfsuGbKeYT6IlktJUVeIZOaZfeO8hr1M1yQW6eFG18LvYoaSljxu7V+Wql4XewIi
e8OvECXTsijNH2lg+SPtEvYbcoRFkCMLAlEPTbuwulY0HyovtsecuHHYTlAP0vV9fPTBYguICpZ6
pOmK2pMCnfnloWxcRAlpFBUqpkPySYIvpaz0OEq/Q+TJrZ/KpsrH2npUimusqqCNM+ovWr1/Bzuu
FgzINAifa5SI7Kn41icw2o+GxLH4eQvSDhnzXD5kX2LZqNgghWijfwVDJP6c6kkG5XWHwmXkN5pc
frfqLbHi1DPM7p6Ybw5ACGTTdeCeYUpgTJ1I7nPCM9i1URvRI2Wm7/aMJNN+7sQSzIIBJH3M8eQP
kHuuZd/80sbdG/vzFFXIO4S8nhP3APjD0Vzj7Lo0+7zM/Ya+Bu+ZgjFWhp+mUTU4Lo+IetK+B/YQ
IGJZq+6rh3JKl7oV0vT84x9xxVXeLb3PAsexmDrpQ3KeufRf828NyYbzdntlJwprcAXuu38nVIM4
uCOwuTrYkGORWjmG5qruZF3tIdeHBnW3NHqtOcd6LOKNIAzFXeQlwkjNFwM9n0EGSd6uLOjx6SKd
LlvjtwCdWZDJ5JtFVAaN5sE/LPM6vpwFW1dAilXCepYgghYo7jKLD664odG5kjwoNGgEonR0KGno
Bz7MO+Z2CKv3GfJxrgsAmkDthDncx4MLUR+eug+su/4BfIbAofPNePBF9lxxp31oELK43DtNEdRC
/D3uoaI6m+ABtOW9qOeYW/UVUpfxwCGB3WUF5R4PI8zpIl+G4nD0iusdtxhlF/KQ+a+5C/HpStlC
7dgX8HryAFR2aynaJ4aEVng96jT5A9l/ajlT1921QAgk+PRTsMXTrIr6UgHitImKmR/KvuI65zvp
2IYVoO7Itn/KD42znG8qnLfvkdSUCGJ0NDqav8fE94EivbWpTSuW5Enud/5ox/fnnaqTmaBpxZQa
NyfZLdwivzU9+tn3ke749yvaaobqNlKI/krJFtr8b7JVyDVqNTdarqedNWviQufsc9Sc0GsujgJG
bh+HCRQ22a6Vr1NAJsAMC0N0U0TcwmP6x+3Pp18STC76cot7hBt7rrYb8y4GAaskdbFuZIivF0cq
I5ufA3AZ9bVtmv03Fx1qgsKyqI8z1WR9x/qkAhMRPwtbOHYX6JvC6b1DY7T3qncM7XZPrGz09KGi
xhw6HQX+5+veb9eV1tmU3xRjmqz5Qsbq7YLMzVDv8hstsJUuvuiAACR5O3UdiSGcbLvp60lKFJW8
VFrXszccK1BMd1UBqpElyyuac7BAuUf8UhF7bK+2T0orkakvuGdKhlhNecen9Ghu8H6Yv/ZV4thW
NThRE2Vro/WmaEHDxjLRKjrnHm0WhlpwnB0Z5vvzACsGNXtguigEgHsTl5LELorOJX5YTmIXw4Fw
UOrkeplBV7PLvuIjlHAzJ57LNjj3zcRu7MkUCaIkfOky4AnIeSIkTyw4Mzk0HRpJU37u5F3JcA4w
1Ses9w61K5hIApPSe3Onu+eGqeCRHbDDPOxIaAAICqK7TY1P+AxBABfkFxxgDEOR6X1j/SoIRwTC
9yXzo5mhkJWxuJeX8y0MKmG/32eBu95tMrS7lKTr1GaB3isu4TSbXChKQNv/AjVrnbpamjG9IP/l
y0CKZJL0zRI53geJZFEugTgMf+OM6ZXTyayVvvLCvrBEJ3utyWsWSmHUVxFT+/I4Ts/bkwnyI15K
OMtEG176de78UvsL45HFVHIFiUL29fkW809cHSSZ5RL/EG32txydRyDwWMRP4q3vTLFFlUMZSjYk
KP6eGD5eEcr8/GgtfEtNlctMl7xkmrjp4Mavy1XmCv7on9uDnESz8ZBkqWiXxaXA7PPiedFDIYWP
dLO9AC6P9+80Wm/epK8Z9wfMr9l/zNiNF9/GBzDugiizT4XlJP0uwQ36ibOfXJ2fa4Bawwkdxu5/
oe4k5mFBA2+Na5FQiu59ZDoDW7TClrhUGcCphOuIjPfUImz++HaNr7P1Ov0Y6ed49XvyYVT/dw1d
CM7MNFRbt5LX0Uwvn2a6n2rV2EXMwKmppoml4uuy6YEeA0EWFDT384/k6PZI1orN0+0XdGR2o5qd
+xv/CKGAqV9tCXUJuSEMDKJ76MvjgUBnyCTNiHLOa/O4WOJil1vXNmiMTK4M69KkgXZ7rgt6K5NF
r45GMii2nn96YbDmk2HMX9Cc5dcrPh97tNGNQUP/d4GZt1xKG1jBjhxQGrTWEM5WGZCc90SuLMZn
GiGQpseUMdRmcuqqv4uHK6+Jvk0Z+Dy1GcNj8gmgXWOSsFB08qyx5Vf8fRTRbatZNMHZIdJzcVyy
XBZ16j4sgxvCJXFUDO893ZrezwBvOCOurSZ9s40+2DWi01kiBgQAzcV1VT3bicL2dMruiYHby08h
UatgcMan8/U7RTZpsfpdKDNXBOQp+jBWfW/+i6zX8BdFnh/YpxXhs0nBAx3TyUzgaosr5O4OBq3H
CSPIakRJHmblG3qWQ3FyymrxNZC+CrJcYEFVDNf6lBM8/oivHQXjQFHnyN661YnZj+DpUM6nfgwE
sXjbCSzURQaIOeVlMoeSK6dwyyc+NA9/Y+8GDmHgWOlejRkOJ2fv66Hnlh0iprpKwUrNWcCKS/9d
Yw+H848BLfLT29i4/Z7eGC0QE7PgWe37SCv4RIFEdz+UgLldRqfwbLnxw99N0pC6zodq2UJYXtIx
2ha0/4QzBtQqFkq7l87qjCwaaSbPFevlSnewWBSSzkqurz5YkyxPBXmu6vp0QAdwmXquberzBRK3
Rcqht4T9NJNQ3JHsrStmk+RWCM8S8mDTyM8DrLGucjayzssHS/iZxdxBPhQEpO8NJUkqTgDroqja
k8+k2WgdnnPNJjiBN+VI4AR+b3wFlIeAe8uHs5MAcwJn5FSFCixB9niYnOBN1UZW55r1XnN18xaT
lKKG0wWsUA2ySxc9oTZeVbmTT37dS+kIX0MZllGWQNeYgyQ1f+JBAmiqotk/fVCDp7wTBq28alBh
+zeVubyEHVRC8MZd/UfOyKdNxAs4zCglCdTOj832wn0MTB1tT/zTw3qBGvf1+gZ+ptayJWXgLsKh
BZ2Gs6QKWTnEAiOU9OHXJnlCaABiss55S8HdZUBY8vnpV1hW/8iIiyE564PtrUnEvou6SFz9mKey
Ng5kP93o/Kg5akg6BlNs2nbiQKXXWH4xP6zDMLhtBwFfZwHcr/OPCkrwPimyB2gPajvmSFK/wJ0j
p0WTULh/+RqT4GKeRnDZGcIPU2jvD+aGJPlVS/D8U4nUioEWO5sLMQ47hB90ufAAbJJInEE8Nl7f
0GmwhyrV2RXZgb3Vyb7lsJp4pwqwdTY1ELhTt0U+wrpkNSseBQJ/p+9lZtWo8vq1vdb02EJU0QLP
IlksPhevvERcExBb2Jk0oNJpammemozKpwBOBr8nLDKWnLxT+xpGAXcqL4tSXWqal/Nev7KEwz+9
km2Xd43MIHs0JrUosRhaQ1CczXX+uQT1JbPpM/0N/cZ5UYn/JPBWKM+MghXsIrU9E2xdA4+/aq32
dOAoZY0STrMHXU7uZ8Rs8E+7i2kLSGC0Xzq3OgdKB1R8ye2kHJe2/T/GirwVnmWdnWIRG8ziDDpW
KSVOkXduJEIVgFWkC3+T2urd7edtnXNTsXHTxH1owA7MLPW4pBX7/lnFiIcRho43nJFH3CE8bl0f
x6tSHUQXH7VUFBCcvc9Fubq6BfYtAp1DiUr+lhZqzftUctcQVkRggSwPubSH5qcmtjJXaXuwABuC
YLGdjP/48bUbGwNTTjmvmkWLTqOOSGzoxvOHAcZ9sEwpUB0cEwNvYyCfMdVoQYUljNONcNNCjr8U
FTt73izGmTwDKH51y0M6c32sWd+U5Q6l0vADxTOKmptBhdrez0PLW554d3f8hKjEqCvpp2piKdsz
36mCGQTr8wRBs3ef0rJ6qr+P4c8F4Ju5MwADjECZB7swcZMbhnq5G7UcwZt6JTOo3JDDiKLfSRs1
+bDY2UiHiTrfSyVLGHdAvQd3XaugF4t79ywbse3RuoGDIEYy8v9AXvuKqJJU4emcC6WCRmdG0KH+
HA19Pq9hFCBzpR1GoVrNZYoTTKbrEXOY5AjFlM5i8Zg6WdPgsTvKYIjX9DFNNi3ApiDoAY40Xuo6
ROLZYxVR348ZIZWyD5LO1uPskQ7GtRTKGIHbNA7psT/iYT/MBEz+9hvEQjSw7yoIibdm90qtEQMe
p6j119g0ysd/NnNxlaRKeLePrsFnHRyXco8euu7h9Gyug9nZME1qqCec5sGHapy+yNXLEszOLFHB
yFdI/ruirNzSm3fO21aZM9WD2Q16rs/siJOa+SS8oepaogrEu4i1YGe24ATEJkiKFEnI/soc9W3o
6TXk8vHHln3gpe/CcRsE0aWRbsJ/EjmrrjnFoKBAov4kXFPBYt7EXOnk9k1OF3Dvt+zdt+isUynP
QeLftQcVixOO+AL/FYAacQkwqtbrb7EOeMxypHW2uyybetpUIrmjsyoFEsZn7MO5+bahIExJ7Eak
DtJ695zJAkPuV8ISd/P1kVVWvpQIwA9KPhMvNNaIEm3ajAPv7rRV2U1BGvrCoXik1F2aA2YSm9Sl
enHn8TeCdFNpkmVWctxBTr62O4VpwtxgSEdGUEcodCoeLXthyPwNo4QboZo63G49LzBMgsZVggvY
ajQfxHZpg9OOZKNf3WYz2RBawCVKEb1u3P8nyqeLn4dmveHGkC2DIMBx2i1p5l57f9YwEffq7wXB
BYWcENxCS4ckZIIxF2QWRNbz7uoAOwyBNVCm1UF0f0VdLOLOzJd30SZqEFDysJSVGpK1CU6cfCyF
QjG6ZDeDqd0fGOmYopopQetBelyIMXaXXX+Wxc4LQxYLlu5vgjpSrsT6az7i6PdeZD0Olp/mRGLt
099JUI3cWFIcrchmFTndbz/jNbu82BjnJlvLEK0qqXupw6wSHxDLOMyVpKPldqCa5V2BXRq8Na3k
TTlbofJZ1+2pJJGQZe8ypx8DhSJZAm48b6NxwiayW7KkcCrwn1h2X9rDQ2mlpL6xoESQLM7T9l55
/d8orUSdh6sdYn7s8xdxEoPkNMPekgsJFAzYUAIWCAqlKRi3WtI2uwqbYqTv4WZDycedk3Ljg1FK
3Y3ZiT7/Exunvn3hxq/0Gerq+21K9kGOPMjYr3mkQpMcxb8CDHyKPOySPKopUpPy2JvvGd1C8wWn
o9ARqr8ojMH87Ev0Lm7iwWQviGJsd8aaAZ3h05fXbPc4IyOmGMAw3t59vCtl6d3u4SfmM43dA93g
SatkpiqtvtIZL8brwwyJG3HSlJXKY+Ky5taGftRZSNbq2ixiOYVJCYGZ0c6yv3ItxEe8TBVaz+dj
/wb0rSRuOjMr9JKIw5hTs//VlA2Ga4/4PohYzfKBEW5rnYecrTfO4i3hi/wkYYI2LF4k5ED+O/tS
S/h1U0KaU91Rcjfm+ulz7IWqPcVxcI5LazGo0QE1OYKS76RjE2vKqVSXIzcNtPGkprqegTzU0byP
olea4mXNNAVZMQ6Ju+SXFiFWnUCtrdHErC26vUSnHp/JqstUmT9XEB08emtAYPvuxOSpiPF56wYG
xzBQSsQZdpMh2+XCq+1WXyvHZ9NzC2zgMsIHtm2UtiSk/ssFqI2R3AfpeaI/o8K8B4+9mLVCbl9/
qUyvyQCll1detPHPgqFnM8XIqnCoFl0n/W+DGlg2K1oTAWosWUzJnenKUEuTlo7+ZckvpkvT6iRN
yjppd6t7anOvcXd9kwbBfzODYaYZ69IzWT30eJThc/pK9kZ3keEzEKlejSQMd1PLBhWI0QT5pENc
FO1VriTDvlhhKBVrgESsoXB5fFvFeciPvrYuK9kKKaZgLl/oDWk+V7HCp1SOGbmoee9W22O/2Fpr
QDSGhrYi3+7b5///KvIA1wHwyIvggyh+x7KrVsC+CggbqLBwyWv267BBZgFRIFBUMBBsC0aZCznP
1hhw4LmSDP+0XoVv0lUeITkDL4TJ2EaWdRctwJDyZholLA6NQhHFQlbFT5lHeCvSucYvJU/S6+Wg
4yNqD/HsM5xAuIrGyQfsTff2PU8lIesbmIfgige7SyMRsoHFOttzOIvvM9BEUQls4PViXfCq+Y4I
BgdojNLQ5qeZPUxpBE7L/ebjEuKakN5ig+1X9NghRbVrOqBGbYZjiG06QCGPXQD7ltwzNYsF23xY
29EDDc+Dh3Ubz3PTDAAte+uI1FEmDGM7hcJn9ZAYc6OJ/VEibJ7+Q+779UiqY/ca02VlJ27ay/lx
3V68RF46xINQGUPY31M5t/mgAiaYAQsFWpsm57WjJZCgGO9TiqBDofRCiJJXU6GZf2UkJFEBY8/a
/g+U13y7HBfvY5BS4+Sx3jm3f7nzk6wG0cCCRMIPVUvUn7PrB3I+tu/22zOPF1/m2+DSXPflPap1
uwAZbk7dp6xB2GcRj/SjZasfd5i96fV8T39qYgzuyY3wa6G9BWYka6WTtTmqctcj7GHHTzqpNgiz
p0xg8JBaFU7nWOSTSBLRP0sVN4VordPz2MIC5IYIraZksCpXKSdpOcMsXu5w5KH8KzpS7C5Rice3
YeF5GKqZmSfMU3wZfCC0sN9B4p4UTyiGeeVjBse4G27qNn6thF08iO6rcaV6DHiU3HTtReivG/9Q
hfWhbMbf/snTw0/PKxFwOiRCecJSTeJpbEwF0rcb2UHoT82vmKOBHIA7arZI850TbTFgqLpBATGM
QUHjBzUiEPyvwynN6CX6FwT9YpMSi4CzrKG2KLE0s3xrhvCgpYParM0jsnWuc0UjG1DwyYsCvqaD
7Ok9guWVGaEvGrBnM/VOuD8HMsShJjRXzd87H+/1jYBhSDlJY+4zZUO9+T4FL2uxlJSxcjJeSWLG
GNG7hrbJuLXS0XQlnWSeOWDrkztkJ2cotmODk7QaJNZZ24gLa68z9Up5PRAl/MY+25CEuhC3eUun
dBP0wQKZ+dbFktewloZZ1iuCO3pPzrTc3qJS5YoA1/hCjga4WgZCAnW2ZZKXwU81TqAENdv/RkbF
CFw8/fZlaqW4SQZvAxKe7ZHgMw/XpWfZymIFNa58JcZXdVakjRK+JOZGhfYtNrleFN1oQhV2b2GQ
70NcsK95H7SjNMpOYhpOOqTFPqiP20fi0IS7mUmzFNuAdyqm67Au9pAE3FGWaIo1yCpm0f5Z5x38
SLpWQjK4WflN0OMXe1IS9tt3V2F4J6H8gaclerkM9WdLKBOLS/zrl4jBWsUerDpEFGyi1iSzZcO8
OVZTdXUXLPkxWV6l5XEbZikPey+OVWyEyr3PMKKT7jMILAeROaz+NsbRY88Uj8Nd9Jy7VssbUS3T
YfgkmvGRS/z1li08zPrz49kE3uu7PcZuDkTlxrYRzwS19owSx7QabZPnTGWT5U5msE7DctPBFism
iotVIJ8qApZJ1wEOMVK4U4IoUvutoBzOWRD66U0nC1xDVHLkBGkmtCtrMt0boi8uIwrNChDIKv94
AKQQDn0TmSoFxrUTP18cdjvtq/hH1S6IE+uW27uTSoG3/HrvA4A6yiuFBiallWJ4+5DyX34kVq7u
9oB96Am+0NuArkuRX/AxLqjUG0Njo/W0PBcxZ2ABUR/LU4RdRLa2/kfedR0hteWy2xsFu7WWuJYZ
AD5js1tHDV1jkOzPdn7SANhvEKYNUtxtUimv7UhRtgkS1d/Vl/58eqyuStoN6gKh1HSo8Aqgr4W+
nfcHZp6/uyh0cBgr3Joot5FO9NyMzLeV3f9lpjz2OBvs0+xu0YlZnH8nBkpG1X1xnVfLY+JI8Fz+
D1pw912jl+azT6SECVAq7rGpcgc8DNUY9fSj0tjIkk375WLqmufvegY8P8GdyTR3QEUamCULi/bJ
2+Sj2vBRs6T7NYVJEUUl1Ak9F5k7cHkceFcj4GO60FiKeOQb9sWNEl7T7jUMsYGviCwH7D5zPJ6+
u6PHxmdZmMT4Th+qTs82pbb1W2eZZ5b8aso43rnuSYffu1xbtrig28Lgtt6EbA+UZ81qlnhQYg6Q
y3DfiGye+hXOfddHtkVsmjHELO46ZtkT0uxTmNnbmvitxrwJ9NSk30HpaWTF+djB6aMrpF9TXPwB
cRlUZPhHgSFixwv8F7LGgeFezkdcmD/KdxYsqpCWzEw9LMm6VnucY0FrCoHvpc9AuGnyxD0NwzuX
qRD/WtG6g3BLrKsdqv/k1HczhBWjgiEtnID7wVXzDI38wKLwUDudq5yGjopWQPQhY/n31XzU3QJJ
5eSL9zlBmwk+4+gfJXrFn5pvBI6B2qzMgMQ+j9xPBzE2qfJgqBuFZX0RQNrjwPu8Wm7JOsvq116W
btIg6YQ5k+lB/Khx2nriWztJ+N/jnvilx59vaJBBs+I9TyIzM8KTdJUQC7kztVrMPP8CAuTRRLK6
Rn7mzyP7FPaktKArMswlCwi2U9Q8CULHh/5TP40+BalCoK545Fs2GNwfUX0OUcL+jgMy0/8htSlM
xyfztQNulo774RaCHdwdpvWHq6XLdFAybnkSp7c837d4K93v0qmLPnpzurtrXfH8NPH4cj2vaecO
X8U64wfSGEiJMYobBFRISX3xq02GGvFJjrF9yAdB/gDJTWFqBLvBSu+ZbjiFZyWbminJZvNeCwvp
2orcLC8/cyPUYmOIXFAF3TTnDxJ93gbH0uqykd4837FNTO1nXoNYZAuLMPjW6MZYWNGbVFkHFm2s
e1iQ3Lw30ZcToqCfPUYWOkE7fI1mfGuhPkr2Pe0cT2IQSxf64BJFUDiwGo3R1dQIms9PRnt3xy1C
XR/SiIhHbeYZ1ghcsgPGOlZ7wQK6w2zOw3+Mf13/RSPkrj8BUctf6Dd6Wa7eT7KQSE+7gfzJcZZO
IE6E9D3OzxPUZVuQYWtTLX+XMN79hn4BN+4zeBWN/dOY5vuKWAmWdq+HNT2iZaVkQEqbfIOmvwBO
K1UFnUkObzdSiQOKIYE/OTp85JV0IWX5LQxkHkKBpIMaCwx0XCxQ7yPWWGVLxe7tLnlWKT9C6/pq
wnaYoZ1uK4oR3zCVwm5ClT84C8OMARiyFV4xePanzcK6PP/1B2aLYaAX2Af2r3sIJ+6Locd2u0zB
POzm2Lu3QSynG7jdVllAnEwtn3pfGpVORYXToiptBGT/hSdsV+sC3RRQmWU+9CbEbLVgzrc92cAj
hUve4JVO6ntJhaGglgoezmDyw3sZc5r/HjRvAf9ADzfyrxb7/8gV66Ki5O+deK7FCkFvmJ1WHmGH
pzQYhPRXZEygleP3xoqPbZf6GIRObJKOZjlowQ79sCSOpFwhn37l3Y4H7tVveRGrH+pHmtCwLY3H
L9N6KQM6mi95O4AxoIHGiSxEyJpSCnY+q6m07mNjVRLoh/Uma7k1wiecb3jGVPfv+ZZ//9jlBZUt
f+g5ED9ztYJp1CyPSX7nZSyRdcVuY1MrNIPorkCIiFL9Xfgi7tKtijQ7gjsj9cDLb9UYfb0CNFlX
W4UHm/ptlMdvWJt5PRqLCNOarpoEa+dvkNOx7G1gNuh+pfDEBJjIRlpc5FKcKox68eele+x7qj3D
y0hPk19grMPvSAEnaMcLtnEmDqcWxdta1HyDqI91ZkbR7Jk3zOynaNzke5m8UrQVSyBdmtSFJwpu
HMCx5VgdIUIDiTUmr5cprEN4fUYvn7oR7D8kZgp6bN5rPc/g9IxFeI/05/gv4xPj5hRBjAWRBUu4
2jJ6IUsSa8OnIRw+Yg8YbfBEYOMg19B+LHt3eEz2tTIwIiP9hXaMD53G8OaKL6wzkoSuzEZJzY3e
S7XrmFoXFiWv3F1Afo57JyPtFNwGg2gF2ne8FQbyvrpR4FzYt7UbUVcri/OQ1ZH66XwAqCnL3i75
YeNHmKp3hWMA+NH3+nEjacUDeyx34CGXpNjVA5T7+8NIAif5VvbhIEO04w7jFt6kuehZQZB76YC3
/2aTKaIaJSngrCbkhd8mGWlsSgQ8OFvBKx6rkzWRFNlQ6gn6pBT1XQw9a2X9zazPtmrhg9eQedoe
+SP0/oB8kPyACBRGlsUyjqoeRLl490LYcGfGQHuHEjcPNahEj38599fgykzaDF5tYC/A46VGBbWb
RCPIUr2UFrXTfIBv9VvxSTC++/SoczB19Cv6k8pBKAfbo1G/zZaBwz5Q4QYz/sYgCJWiy8rfWdvJ
KdGCylnmHre5pDmubSsUDSsV4mWuzNTg3sQp3yiCd7vV2q5YzCZPgQ7O7vw4TC98tixITypGKpwJ
zJzwmvYpmk7b22aZqYM0Zc0M/HPxr1XfZ8aVptrsqIO/W/PmNT9mouYtKRIxPh2wxJQLLk8Ubxqz
uPWlgg0PiRS882rb75SVNcsRpwQx+C5WRPOkCEjmQ91yLf191d52tRDZuWLKd8xoyJ9E4+oPzRPQ
auB+Blg+KPUzhN8rncfIX652YFojCuf3eotsBR3yb/jpT4x3NWua/k7eXwcVyecuqGY7AQRw8YdM
RidFmakEVdBc73TP9wfgXfSFYcTpMegkzoQf8B1PlCLcGPgZf+FTe3yv794RNNRpBiHniZmPBAve
NcMzNpdyCrcnWnd1zS0jlLkDP/cZaq6PXEpg3Ds0EM6OzuNONgSxl2NAhEk4zJLMQ0ipREwaRwb2
RJVnyMAxDZrwGerNAzJo6wodz4TUckGo1Oq17DD1SGOHANN+id+W7aY0zIZSJ+m/tsZcUVih9KoL
FGOfjDZojyr85vaVWa8G6kECx4IfpKsBt5jocd4nRgA9iL12syqmKOL6UtPgPCfmaIlSWHgE94sr
Fe6T+GZWK+V/GavwrVtWYVZGMLdXPjgcw08VGGtNW2e5wbHiS6Ef055Nqb77fMe8sVcANVdvNNwu
mq1j9IJtAYHMdZ1NvXWC6Fk5IAaWaujq/829hF/XAPyM/QnGS0uAGTlS+xj2GmCKvsJrPogAwope
Fwx+lStjliqZCPCzINzAfuDGJLgJ/z3tPqQY+xxGan1WMXVOebvpta1TmL18Ru4Tc6g4x/vLw5K+
Yy+dSXWrrcCj94qX8D+tuxhwXOYyPuQo19hGUs9+YwWxvms8qu0YMWZKmoKbtI9ECvEB7cUBeofh
vnB/W2BsMchN4gKsoPbyZcI3WX51a0G2WRJMy7DNpLO98aKszbqkyxquNJZ68Hs/MtjkG30gJjO3
u3UQNF0/QVdC8sxz4dBfp0ZGcwSSpPByXb9XIXJHqgqejeaShvs2U926+xhl7r4gbwSfwBELtZvr
Eh05mO4QV0EY7RpipX82s/OMg5Q6BSOBfvgswfJQKt+7IvAwbISwtFDsliPQNL8bfcfJOJO1ppwZ
Bf93rKizkgsWr4uTpQilXFBEXjWV1tHhGOP8SsTZUsX80xI90ktYnCQwN33J3jqKLkXx9E9wxnDe
cGoLQcodpzzOYZ3YcYjD3FAIyhqHJAzYp0Kb2awuCFBBNAJQVLaDUk1FsnojGTjy3OW7I0h+rcpm
4DP98Cli3Tl3QaeKqwEGMMEL/OY9CEUluSlPrvTv9A5C+FjLKD7K6B0K9b9CWTFRFWkzfLFqMpbV
tRo2jGKRVxGtUDtGRlPOe8l4klPGicgbdxGt4f0rcQFQ1Z2vW/l9aYK+IPFtviDjxzDWYcuD0rdj
CwzGxlTdAc54mtAwyU7EogSVqowSBY70rrDg4523ynVLfN0REpNd1CYM4LR6nvXK7v2yNkrn7KWr
SruoSfi1sKGEgT4xfmaa8XHRh3vBLN0A+kRRFN/9WCuE27uB6TiaHJecQ8bbI7aWZ7QKKxDGdRIS
NO8O9zo8zHF73VlIME9hUjOTY66V4F7QFy6ZYLmI7M018UjgAPdTNcpYc0j9GfVn8vUq4W+Vjl6a
orw/kwulHq15J4JPmtA+00REcf8CEMa0rKlHzkOeG48Pr0BXUa491v0a4T3zIw85ybPId5ArHGF1
AbslHzoxK0aK4dYcpeDj4FNKFGvACd/4pFfw94M397TqArErZPY74oeP9n6OnQdp/W3ZiH8BSzrZ
00Htz8KN4nTlftnaJZY8HrQbi/JQOPMHlPNviS+x3q9iBV6WkgF9S2/OcE1RYjyJfcaaScMQzpJR
mAoaNNbcKshdtOdMTaihDZWjVi4+NlC4L+P/klq8mSkW8umjZicA7ME5pL7+80TcWu5GLNPWttlO
YP6oGprtBVf/umo302nQQLqmQUuZKNKinVz5mJoxiArOKQrWSM7Y3n/A/zPcWsq9sgA2VMTt5QW9
uZSz9KyXbWphGDmgs0hdc/PHNNW4nFmGAYYFZHV1tLWPwPvByQakRIvEkVlS5NzcRdhxP2p7gixh
XioR1HryaSVmrZ6u9B4axLNz1Iyis0fQrOymh7chw9XwMeRKnZJ1wbHE+S6FDajYb5qyau5lku5B
amfCjMdBD2XLhJ6HdLF/eCd1eTHLKOb5mGGX1Ywm5r2LS9En+xRMzebO3mcadccrG862I9veKv7k
dFoldpcff8Q1qDf+QKGptVQmj9RxmLJmnpSF8Z8Fn8Lai0nLe9weqAr2Leea+hNQQGOkpMnk3feF
e6CvVGmDiWOXE0gZdJTGML3RQc6oBvGBpiHAE5I3LZF2oo6Tyh1H9nFQYAs1eeH0G1PHeL1ASCCP
0GD+phy91UIf+bmgFZ4WlmB2gM8+odJVM1z5n/7HatCPtwCUQ+TYPJT32ZXzDPWTZLpJCY6S18z6
yfihdVx7SjRXwobCP901azDPIfCQTYvAm98uceC71KL1eRrs/F0wDEBG0U8peHknm8WVfxXKJpCc
4DhsX3IYnKxyPk4xZfet5n7TXUI7//LkABlKPz/fEuI5RGuPLU8GH7G3gs0dMJueNgtBK1VNls5Q
zQK6GmvVnDmTNkofNEYALoB8mNIH6QZwKyxzi+7/j7cQsYQ+O/Co/JoIv2pJCNfNVFujrHFECpxR
EHCtZPSIc+vw+JDWrTiIAZZLWGgdgbeZRAEgL2zYJlU7Os1BTsjZwZmAw6FeTbBr94O8ZdDJ20wR
tx5FhYTYOzIkPNed9LbSsIfza3w4wsPaoCmAMpQJFsbnVhHS8J7LGe+1/y1LsbhthzWroSdWjWZt
p7zRmux/PhAN8L6bEAGSW+VwB6Dd94SmeaaipUvQ7b035C6tZmwtklcCh4fLOBzLBzpYNxl+BHkV
WZioGkaM8+c4JEkBMc7I0v1L3/1tCrUDDm+r7ousEkU4xHgBxLja2PHRbQfh7yhZzCT4e93Q9B5f
+O0wHdTI+Jx9cEBNS5lcAKKJ9Y4ysr1PbJwOi0VP31Qo6/dBPBK/0fi3w/8c4mVnzYBkuz+TNiJ/
Hx4oumQBGyBCoByzwD5HZHg/FcBv2cFJq7RiLslrQp8yDqtqzixTQQ0uCf9DEIUUkZn0QenHwjvG
2on+Nwut8LcRCMW9+9yfr8GcVKAcnnwTkeTvRrlYNOl3wd6yw7+BUO8SSLc9QkrkQlPS+DUnLH1z
DQQATseV35In62qqolxwA6G2smU7vsDpzLtUpNSt0kUthLDN3+mBmMNl0nPQk3Po/8/rEMvvUzRE
SPFCrU3gDblS6bUjUZkUbSuoJSw9fJymobSatvJ/R/DN3Fb3/s9cKu+fXR2YUgqevMlkYWwCQaUN
PT2IqP+Vh1pS7goeLunzLVixP+drrGurTrPZyObSX3bZlE8+j+AFQA1Y/l9S96SC8z/vHQDJKQwa
/dt8FvzWEI+5qLypDPP66DK8rqYGsis0aXCo9xznk9HspqtoJCcw80C8Dpqr0zlquT9gchBKH/xv
QOFgelqnof+LuADDiqQNAVnbgoJuLOkramfTJ99q2S0yxxyz1fxhpA6Tz3XxQgpgELKb31C56nb8
TRQdOgKu+UrkY/A2fNgM6Azw3mE1nfdu5zIDvMa6AP2y0lK9hSU6SFqJKVqIv6BBDO/UHSIYG2F+
F53Wd9bWSfiUrF/bY6a6AkNfcfnm4CC6xkjQ5d5NnhCDV++2nzlq2ZSJhxrrqCKS5jkwxWqBoPHf
uqYtgqANF0uN80rFQPR9xEhBNp7imIdMKVFdiC3IOLIHKoFbwkXiLwc9J/AlZv1cI1Xm1OJlkV+J
8ARfzlmctMUGyLFi5z14QjJ4j9N+DVNz9H40ywutHyu+WHj4S/2GkZp7a1epIBVdjFaruKbWNx/d
L4vhC7+0205PBFW4hV57x8KRwvxLR/hvmWpdgDfTGGc4axtDZVjnIXOSwIz+ZIuaar3b0EFgrObb
TAZTxv1D0DGelIa3NpPoT4ZhWpR5YqQRV4nRb766LUUpQkYpfaJmxWvdKwZBC+GMijmoKiGPC2Sf
wlHFLqIq61sJSTV6oQKZ/hEHvKjcwxMViFPTJydRU1iMK+/G0Z8c5GHyVoLepsLXn/ObnsRTgm+n
cOsWBsLd3V+HVElM3MeB4hHaaxNVI0QfTdcbmNuWNpGp4ElxyjXcqSIRwiCkmpTZi5329FtrE+lX
GrXDd8jxUCQd4T74mBddjqpLbGxX69/ZteastzxjBgV2zwTN8PN2/MQlShlmLUKFhHx73TtLERQU
Cl8iyb54jdVN5VtHRzTCpOGoXJEuuWd9/tlPvxarAD07Gb+szz2J6XN8Yn6tf2iFY7gDDSFfuxYA
5rJKZOSJUlxeikdN8w6qMQ1do4qTeGNgw6NHzXwG1O4PrmL0ZjchJg1bSrIhTH8XwDJIIlqfmW9p
ZmfHtAvwRAzw76PvD7a/WGH3a+Vp6c5xccDBoANozt4CINJWkHMIKl+LLfqatzoNQA5zTTcWUauS
05MGVDCG0hs3N+ItOKCjbBf5QGRwB3NkzsbFdmbl4A+GsLfqQo+6/febz000+F6Rd7G4OKqDe0+b
RbMSTtM9mvkTDv43QOmI7qn8ZDlGegLxNT/Nh8yMnjWyAy3B79ZXvxRIrgJvH5yG10EMq/CI9JkC
TIFU8pO3pLSRmhFm61HkxpoH1zGHxkmuGK0QtMv4GMlZsnOrzHUeKTPCUyXoPC6568jZOcs2WV0P
LPUD/cdb9oQs/Pi/8vLPoRbtlWrckSwgNIVU49NDrA7XE65+kx8lHnYQp4Bt7xdIGOQv7oqSd3vw
2Z9nmgO2hGv6OKOlXrnFrit6r51sDt8GPoYK5DECabYmno/2qE/NxG9A6prVRolmEtbkOKBl815w
VGbY24b56RhRegb+5o9SwT8QUmjlgf9a63F8Hbkg7Ktp3QGTKQ7oJOmrz8dBBu4dNGnaCnjZsjN6
4Lt3XX9lMHCO4DIPuABt4qCTBH29fLPlkR3TP2EpcPJYLxkNxHkiT5WZg7ll/0CtoP9TLkuak4Ii
ytnVFYd8N25xGB3B74GAz/0PpN5oziT7meYTAIvtCb8BeEPukfmiDkrkoo6H6+MLypPe1izs1CNV
K/q3dkbSqyp+geENgXmim4wE6rLoO+2Z5sAZwEPfQaJOrJ7mYVsDfbfa0Bxo5hsLcieS9PB1YuH7
yuvqbW9sokjwhH+YrKLNzUHBQ1hdN4Edn3tzmRSNhFZaK91PR9WwxYnWeWOBr6jvxtqSNzH62SSQ
sBJRX0w2ooaeEqfB0qjVLpAFW9aITHLN9YWwMrqFNqjMyKT+6JJ3dhxUUl3CAwWPQRlO36gepBgR
69/NfLBBTMqkk2v4iVv1GJWBbg2GxAgr3aHmXmwDeuiVnrONGSb69AMFf12hv++dUWDTNGj2q+js
eEs6NZyD7nrCRIqjM6oNu3+JDQ/7s2E2dKuqJgPT+iVr3adZwSedoV30gvDahp54lBiHP1/x4YRm
CkXY9GsyWqnasPS4e5lCFHrAIzhI3HNB3rPm74LEfwcVqWmjNrKf6wfOIP266U9oMJ4HdwLIFsUk
5r/BBYvUubx0GZ8uBDSgxP86fVz5t8obq/h0W8Pa6M8b+4CzK9jWHeWPqV2b2FeZp3Vxrk9taHfT
KJI95zGJiu4UL6EWJIdxSqxA0P0zOdKEh/9iuqC6/etRshS7Ipuo4ERW+ydtkAOgwutxDFBV+Go/
D5QEY2uQoU4Z+plABySmzVilQYVrH6m8Y9vbLiS5/G9lIv5selEWLzp5wo2L/VuuX3fduyQ98s9S
ex3V79OIfUayimCgMKwsOBwlv2WOUvLPN8Or+Lz08eN2QEEA1zm1XI1u8QuLvc8uV7aVwu7l0yXR
+A09lWjWEX5oyVoAFAqtjkUczfOItXzkhtpl41HDcobI4L36tVsiT726uATmIJmG20HCjFeDSf8y
u1a6nT2j1qqkEZhy8rIosQBY+1Yj4nC0eLpaPbP9xPK+WLyU+v0PX9xKaCy2sWiUagz9tvQwm5UG
Wbf2aNur86rsukRKSBRoum5/r/7OPvEJacTNVXqaM1KKMJBVZjt+Amu50DUoflJzA7X+usF/AgJh
cy/HpUcuJJ3qECvxHZRkDVDmr/HY5dWy0chV9K0AVrQqtFBirugvO1zsGu+Ogp88D1TerWyXiu/j
Waj35O7xCyNK8ymao8vGenCn4FgG7OEOcL0Rvu7qOZ/HPSRu67YZMGAhozhRy0VHLviCDNzqpu4p
CMAiX/XF4dHrypJfFDBlp3fLzavJ7BaD5+h6vp3B+lYHStMKE1mbJ2OINdFU5qD4ov4oVnZ93iu+
kVP4lsHdBbzAj4AFrSVKwyBHnPrlTIZIhmAr4JM9lCT76Gf7O0aDtRqzQnKozS327XQEy2JDoa72
AzylerTq/DVNc9+kqM/TdguOgTNSqEy2lVEz+U0OkhNiSv6fWnfYJ4OqZLneYPTMnlVaEdyfdAXe
WVAXIR9/fs5NHZQE/y1+FhylzepJjGzNRqaws6YUnQnmDlu3mXKg7p8lzLEhCaVHWmcojT5WSB6A
adiSgOWPMkc41ehrJ2U4uJQJ9PwHv7mwW2xRy92MNI2Q/yl4MkcRc1CqEAVuWMA2fvTQqKQPfmxu
rF0IKXy26Syw5cCbzqBkIS+rlPsf5+fKTfLesTVGzp2vaSqWFG8jjcb0FPYAHgEHGymLgiKE3g8M
DlMEPeuSgtrZpe5Cd+ujwBoeizx6joMtY3ZlnGktocE6tcVUFoK+xe12esZ4w99LQJUELp7gStkw
0BcsGIsTtrRcLjPj8SJAJgz0Rqg+hNqDe6J7ilduyZi875l6ErTkJgyZSNWFUTRjMl1vhfA1tb6N
MY61xZFvdJOoyj62GD3X8UDcQi2hkNoPi94mzn3UgbGr6OsJnygJNLgIcIsdCvvLNKQgq8LI9hL9
fB63zGON0hiF3ygqQzM2EakmLEs0TYf96wW5mM48Y3LxZmxme38aTaJ/UquSCJVeuD+SJSjiyErk
cOunV3AFVO1EjCq6Z5ddV85UsTm/OLeJDge7lAoOierZR6yeFi9oY6LQ2aIP22vxBr/1hh/MxY56
VcATgbYgNJEVLC8IrDQ/Cp8YKMeQztmlUQL5rychoc6vifRRwgRteDNBixgXAGsUwd8OxsMEK/u4
1NEP3x//fXM2+EPHwFXem/thyfwyZniw5CAiHcN2ISgzI7EDmmA3LHV21fiNCYA4TiMce5k9vLbe
DjeZLP0xReAoXfDr/UkyFJ374AxPH/jY0PbXgbKAJvXUKod6Gt1Niu/Nx2OtJU88lS0ZrFvMnd39
eE1rtGI7tBIsOB/YIesgpao2Sfww2b5v9gN+TcwMJSDYjAXoAirxHdd692bU4BlMZO1o9DVlmJkb
ojpotysfNhPj44aW62yHS3Whd3lFGVUQh3jF9OwUavFEvJ0i8XGz51RpijySsqRnK0tPGGTyEHzr
GVCj/dlkMUgXNe3e2wBvJmE33NuHrMS3zVf01A9XjvvZa4hlk88dYBR5grWXUfrvAXQC5V2aS5YT
BL+R8/BGJzkJgJbb1xtI706GaJLLOEMZ0ARv4mO2hyUWrD62F3b++6pN3UfuLevPRoAMY3DbJVII
XDYwn3sqn+ZfUddRbCODJ99M44OJt75TehOCin/JajT1lGgUNPbrETRVTEY+nqBmvbvrMNHNL4Wh
TjQU85Yn9SKesA85ZfJ32r0QSw8f2kg+a79VoazdhFDjL3AJZq+ta2N2oes1gxuHK7WfGF3ZMRkU
3q+AvG3ClVvB373OC+9ODobEpc7YQM5O5PdmwXb2xGB959qFBS5mIHlSJWXzrFvvsSUWp9OXSb0v
MIF9q7Ix13Syf9VC0b3jDmt212X0ZmEqm0n+Be5lh/cuPcnO1DZo1TUxNX2meTH7cDcG70UduKQp
xxGglL5OdzrxGZ/emKxXnLy0SXWuvCnamZUdV8hkPAoMCtR1buAQLroCIUCjHsn5RfvAkDZm0/Nd
t0UfMAla9Bu72/jww2pOh1Mi9R/Yq3rEZdSCm8ihMRGWt4mB/09JTqFYDqO1DTs/MZTpLKCSc283
UVyCoC3TSdLxo/luv2j6b5Q9COkmQkF6IB49IY1dCGkv5u8Iv59XfzQIT9Cbhl1Y5pAWnOJwiI4b
cP+27h0M+o2Z+Xj4ooeEl6MusqgitN/JnqdClTSrVNmnO92PltHV8bVeAV9tSP7Lc4v87ioOfpKD
wR1mFn3sPndV1eRraVIzH9LmuYCKVA+NisnYHVcmAlqkyUVg717F9hme1rd9Caw4q6krlFUEMb5y
ugMZAVyAKR+yHItKrdyIGBSC58PFdR36USvgHxsM+bz3i7AYWyJJLf7oQ0JinvtX2vnjWj8tTmhn
49Ao6LGJ79/LvaJ2r6wqpYg7EoqA+SdKgbxYptgck/pgJCLFIyEUIBIFTSK6tQHBowDSfinVS71A
jZ/kV7qmuacvmj6cnCTe2YDP5gECdjDzXfm5xR/fCsZQJO8fQR9S6nUF7A958wCIP5EYU4Qc5Ojw
+2F+/strQJdfcQbq8qTrnCFDzuLwyC2KlOxWL3OQOoXHg9g4VLXE7oYqJnuAwNKgV0nuJCVel0Pp
69oaCAjSYLn3wlaNLvzUUYxeZhMToS1W4I2Sf4C73IOoOBPFJz3417347/R9PGEMT2aXG80VNWRz
TE/oRUojPc+eEGvclCdY/875ilSE+C7/uizbRdk7LzASxMqZWOAxG81vF1EL+TrDNzvwL7onSbRR
WHv9/hE6W516VcpgbscLhElU+MXeJTm9eMACPjoCrKNyQA6CBflkvnDeFLacAsf7SxXcFA8nKNbs
VOAt10BfZQcGqWxzpiIId9F5fjHKV+7vShRa+XIFnXNKU/kt4FW5oj1Jecz3Oc8dRDI2E09ElUjB
AlDTJCGCzEr0nyXuAMqXUzmyA33c34eZToPmsn9ek/TudxElFUBAmnnd8g0l3Ye5M3l8lOYmqJde
absH/0HvLerDnk8fMQDPLJ+W+pzswxK29nCBW0gHvibbo4zFyknq4Nw5EcleqyMwddGRZ/oNx57u
ft89YhZoUg4wG4FllGkgq0ar+9bjiV5Q++S1C1DU0xqOq2DCadNyasG/5rqsKck00TcCPCRjmads
h0ceJdEF0tHLsUH/6y4IC7MGHp9fPO6QZUilv+1TRJG6vk6JGMNsUXjRC9h5j5/vxk5ebuQyU6ag
hPqNv8NsmINdeJhZ/2JCUXXDN0WbGrCQbHJmw+qlBmMjgbOG8dBEDqymNkqensq+hFTS38SoA7sv
W14axhrDhXa6I3CekLPsgfUHe03p3o+ebsFg7w6s7Wg4eA68kJ913G5pd4pgMxjx4lC3nMiXoEW9
sciMXJSpiKXcbfqR5PrZ17DZQuQWa0UPySq2ELcNXZg5asdTZysADx/QWestqPDsQEn1Y34v9lPy
pT8YCb35Ks3R83ZVibubGj4Rrm90CmDQ4biNCtxiiBaPFg+tZy5Aq1QpsLQYUlS8IDvGIIfo7MXp
8UO7eRaNerJ6IJg0ahlmqew4wSgfrK44IImQ1nvpoWCnooKJ5oNg2kh9edv6ZWXxHRMaRxdFlPZf
3l25jRWjaHLAX7c45dAJ3wcBnnnFGbQMHF/iHz6e3nIjJ3qtwttGptb52gVL/ucXZlbCGKaoioWF
jdH7OtR3mcIvrEVjHJWruAX+l/X/4PglH1LUQDGf/DenR2QmyoC3oKdoORzzHEpkXtXgGhjxSKyA
C4E6z1nSDQn+a4jcJlfV3FWk/4+nV6mFQkXCDTsSdjoVjNQJPbbE5W4vgmffaWCgCyPSBQv3K1mL
fj4RTlhN177W78vjZeDJbeM01RYEcVyrBGYULKxqv4WBqHCgNKrOtITZcekVrlhtEjsM8hUk7Yrj
S2PNVOkpDoBJJ7YOycWvCN0Tl1snKKa2BVjfIPPsPxLYhS8FSriJWQESuxMbX3bp3qt3sbIyulRU
gR8fnfnSM8MmJ3WJ+G2WKJLgbWeVbGG+TvXl6VgSdgXcO7TyW1ZIPuazqtdU1gFKX6r3XhqobncA
99AFsv49iqxQPXxjxycR6XRjTgMJ9fKMUvoXmQpJHEgPp24bRv/sxUrMyonSeBVcjwffMSdoyEAz
dHuvoewNszhAO+Eg8JWxyfgqT5In40QJZJjtpN00lABHQtg0o+rXkOTmXPCgM5oFa+B9jPK03Llj
tU/9QjZTV6TC81fVREZsn4pAx9PKw6fNkXVngBxTTqYqLduxZdA0sNKttRYUX7pji8opwYEu/bTq
YIKGEDfqV+GaASk/xe9/VIQxfD3o/TQJVb9q71pfLP64i11jmqvaIEsq7tGA6I318yGtD1jAKgMt
BvzLd3KNLGQbUooc5KMQvPWq4v7yoWHTjM2ij+fyOLaOceqRF3UwKGus5pbBTDnFMFCzzgEdtirt
B93Kua8ZPOQrmpKiQSCcYLJs4FWf11M1yq82j7Qb2OIdRXbPJyi5zmf/7AT1s0NK7919ybwMCKo+
6R76j2hDhZCCOj3pLCgaQeNc5jTmZD9MDUM8POdVtDLEB2P2pSmwGfN9kBUYQAUUGhheYPkms3Rg
ncokjClNxu4gYzAkRlK5RYRN0K90U1DMEh8tbuYHS0dkF+jG30eEQOWATlZAZletQxM4l4U22MX+
CMGGpmN0s/eOkxmzotRUbLofBWRYIYUBV9rIEvL46sNAo4X7G1V8k7ZxEFmDJ5Ej7IALu66reUuE
IqSvdy/lJfARQcpfyhLWBr80RktE8hoNCOCsxpXn2myZzVl0dG2OAIjccgXiR0fEBLLZDBsjY4qJ
Ed1mFMLXkO1dPhPO1d+yZpvtAMjGbaH93EAkn4TG+BBF8/zxpg823bUEeY6a0rrE3fAbUXR8E1ya
XD39bUqkpyGk5YK7Lcp/1bF9sh/PFGWEl9/Nex24rKGRg9Jhu3mzDiigY/665jCj7bLJf8e/bN+H
FptZyCoewCYioz1OfFC//xCujINTSL0L597hF4uUAObzkaoYzkB+wl8rmZ3Ii+p/lqUBFLQc9Gzr
evwBEuLUyaGfuqARFkvXUQSBMckCrHuLM+ojqn+6x13iUidoG+U/mtuRq6+nj/bFmGW5ecD6nibQ
QjIxq7wFkO8ShXfI1cs+8OnP76tPA0LU2I3FtzKKOnju5P3mQFYbOvYO8+8Jkf/YnU6K9zlOoozN
WW5HhwyK/CgHaQtlacWvFSx0x/G3E8Suaj71d+Zg32Qa1RiVXxiMZ/SheoK8tkiKqEIqP0eP9wFI
u9mm6BCGvbunTsgAyQ/VV+n5nSVzCMfoHkI5CSCJE91i98ghO/lob3nZAm2UUGNkdRBbXaPbxmyy
PrDPbI3Ev7fAJ1v8DCm/WvuCs1p752+uRluebAu8eUiX4Aa+5DBcAJ2OqkURrFGcokRURZsEYMrh
mx+SeviZcv6cFpFiAujLBCMVKiy3wkIchDsVuBgmclefiUqG7RKy3U/c/Ac2qu5cJR7byO+XNCbQ
qNsLsIUGXHt/Hu3Mo8QtvXMwtITZw3vd9xpVTrLi5jpaBTFbTUu6BhqqVEunyXC+AnLRFdUdYQB7
F8kTvb8iLlR7aO5qqUgDzazf75m+R5Bvp2OSMnUVJZmNHIqyYbIgx6F4YxGzUO251QY6FWyizJUY
95AtuEiwXuIbkpEAXfomsUYj1Tl9Aiu5M02Bp9vkwfB4J5xVaLjIjNWP5xvYTesrmX7IrIEAKDrQ
3dc/kHUJstZ89umKw7KRv7N8EDj3BKZkwPX3jFYzth8ZNFtVnPHmlz7gVkpfb3LhUz+kcrAbWaDE
8FbjQaj2EVFIieh7Xvl4YWII9TCMlgt3dAinSEOHZmTW4MwJ2ssIRTAa5lQ5AfUTftPETFTdKS3D
id9DxMc3AyarRwt74rguESGIRv4u+zniv1VtQUp7bmf+zDT3dgxcwtKOwzL7GCHD1/3r6Mny+ILU
y83NEOQZiScQKXlrLpqJlXorXIK7GY/eh0QKo6yCkiDUyjoAeLTeInp5CYmQ8naugAsEy/wh9aSQ
QDAVOPbvM2Iip0tdjfh43O81BEe85DY+8LySF8D9mGSt/jmGHamozMR+n403Y3tLhvEMbxk2zNNz
OkEmfahdh1NFQJhUyCWHGUmh2QafnYSuKnwm9BKFHW1Tm3arkopGUGHnIZhtGjSbmL+2NCr+oJik
iIdnQR9U/nXvvMZromn8af8uPAFmeoJqEnrPyaYqs1IyqB82hcR00RQHZ98XRvk/E7KqeVgg5Sz+
lhtTnMxdSufIRN52lZ+/veysEwzBJsz/KtVSzqNdncgTiT8h+IQ/ABef2HtPml1Xy+aYFAhajARQ
OclVdO8tM8OgsAZ8O8kduISLF08ukfDRwIdNiWUmIbxc5Kaqc/MXI16pf/6vms605bir0VnKaqv7
HnB7XxIzdGAbaSEoZhlK0H0cgpq8VEmhjXcWd1pykL5wjB6//tK8MTjG3gPV+taCiyv3/sNauxc3
qcDcdyCc+cRqKzhaVSPpK7MkPoYqQ5PPKIyjtSvXt6SZJvKkOVPN+fV8/wTV65oX7pllxNtL9wj9
Ip5VVGpWOY85fb3m52XJesDFQG67l9N7aebDllRgkh2KOoMe6AAqiTrT9a0Ux5Zv1WMtwHTj281C
ZZoAhbT9ZAvJISuVYzjoWu/FbK7Nlu0RBtJBKtd8j/ECDbF10rt7UBDNwd91esW9lrl6rtzlKfLL
/D2uwxZVEI9Bah0ocZGW+DjC59Qiq9sla4B44SVrwA/P9WUZZibDlv3wwAhlWgAexCI8pobaLJxz
yqkskSd6IIjZVNNZ3DQ10NSmRYNbMrglpHZ0V/kvIbTaabMo6v599jNHqxLVhgMZl0IW3ay/sjl/
PfwhdfcMWzONeifxD7cYJQHidpjN7hi2A9M31a0ywB3BB6yUQse7nguTFR9GS53o61Kt4EolCN5/
CmRHnMbRssoRO1tdk3Q7h6SI09y/D1ac/ujX+aRlEdIROYL+svUhMrJ5EE1ujxVtbBOhtmN8po+M
sJCqF2sIVemY2qS1wwD1nyA9xa1u4kgclOJXgvbFmhlqD+jaoX1QPRW6tX4s2peDOnyc/+06dEfn
7/bC/ORYKAyGmKLOVhelaFOhMEnRvNArhf6DKsCYSNc3tFA554aeQD9BA7LQB4KG6kZigQoTb7ka
1OXs+aXXVXpKRjYtxAFZJVT6F+QnZpRBtVbI6swPDkiNFZgqJvVMJec/kBL3IK4ujP0xXs02+J/4
oRRjyOFiYUPzqiC3vJg8wuEAzowdtMLbzEreySWwBXDe/X5suHG6X6Mnqf3b2kWVHb53PRXaSUYa
igYieOa69yxDiE8Y7ZQZziHA0VhtHKx8Bto/Eznr79p7bsHpjDFJfVSIeBTCyWH8KZ7Ino5BeCGC
pX45BH/Zh2yZFTnq9/5euYPvRx1huCcHmNfJbEEGgkxB0CzYBzENFOuKZxWK7xnbiR85kZy3M+ZS
FK4OT9aAbtI/9UDjzyL6w9cpDF6Ka3iC5VjZkgTa0TKtzkVqZeU9u+KJvDxG+eytvRiNMSnhC+N2
6iKbWC9luH1eOV7lu7FzOGJFbpZecTsQ2XwdKFDNka0N6lqeQAoDo44KMH1fFKMY2SygotHghCMi
jKRYWFQwJROuo9oeMW+LISzCX1IRCChf+UB4bglNeJeQmF8DyS7ZRxn2kXyL9uN6ejRO+KedIpYr
/70RVAFeunlO1pb5tWPZ0fa2WQgXu3ztz3BhtzZiEdFJ+tBV1HbFBmKGCvxKwN3lrXH8dgHtAJ4A
HM8hY6/4AriEb0VU79hvAzyTTEPdOlFgLl9lhC4JMhsZZNG5NajOJQEfn+HEuJvjj8oSIf4duIPp
xIcgEKe4SSM9+8odgjhl/mRzOVxQf2u9qUq8tqB9b7ak5vSDuwBooeqczoDHzt/aq1UZLPfIjLXt
mKEUB/M4L63/zXB7N0+Aq6BaJ4DVe5/vvIY+tQAlF7s6/0roTncC7ZeSsJBjlwARPTqFbF6VCYvl
sq+6PFM7+ZtZHMwVE+k+g3U/St+xGIDLQDW9cWtsdHprwc6WkizQwGsfeYDbuHwp5VgtMVtICAGG
Fgl+6ZgfOfjVnurPFb7jPFVssi1Ly2uOe105BRjqP0SPw5IHqr4HXzdyQkUJp5fiafJH2feGyXCE
MC6OZ0gwa77a0vG0LY4fjH6q0jBHiTHP/WA0/y+naQFZeXrxdZvVwf3uk3vs8dHKS0SgP8rRctm0
kJJGb9FbuD2eBJfWi0qlNNN0jBOEXec48rJmf5xdeogd1dUurcX7jatC+fkoF+TUBUMXT1qTjBjZ
P+cGgimIwx6MQxf700mbGOj8u3aD2xetGzKbUMOTClkfjrZAPrIBzpJgWFQ6Sa5BdqClb+SWx0HV
FcPAtW/wyq16Zr+WUMxVBAmeMiVn26zoInmXQNPmi8v0/8rhh2X+wiFbtlCNd+TyuKUsW+R2XOQ6
qGWQw3VWqxq0LkKErXtHDpXnZIpJLeVQZvsHykJjR0FLW3q86ZdtcB0/9bF87ftHSCPRh3+ISi3/
feiesmH5yl7J2Ay5Vj471zAPsjyT7pSOWj21EvfRIbLM0H1dd1O59c+4VkuzeYFii3W+Rf9anu7J
0s/qEP+F92dzKC+N12++k75CrGTC5NdK7jXUGb3zjLmWhQtAJST0TfHww4WwRdfNKFZegUHqN98w
5HqLHHHuKHRSXkb/Nb2DxublJJ8A5DWBx4dJezexbWTlFh7409Pua2Wdu+XIZeTwnD0HojVEw4wO
BWywS0Ed4uoPUy+C7WiX5s4y3aAN7qz/8J/rZ+drqd43l6jH8f80v1AZ+GhJFYDsDxD3jhXbc/DD
1IjUh8VT04whOffcwrCbAYgecICuXCay3pqgChshrCPB2wsRjJdCZWND80pLScG9sJeZasSBXHJk
XmXDwyFT8smIaDWqj+/HnPU4eiqFTWNWCGREvVlFkRXgZ1kWzyBjGPLcXhQhu9JibAl+wxGEzhhd
hVqq7iOAwDKeZ4Ay/gEQlhXrMhRwdIihOygao+D8+v3k1hlpK2NWW3uOhqShHKq+kxbOoTmAHpPn
6FLodct+lE1IgK4wmiiWJFyHcbuv6zH7HEWsa0VOkrGPWadH6v0mcr/g0TkLj9awZ5hbPzc+e5ZW
0ZlnQ3s/I+pQMplolENnPkosXdOjWWQj3CMqlnZ17LBopQ6sELbHDC9S14Atz3Kf3pOxDsv4jtF0
kUAXtfysjmFa6KPtTjKRaTGS2fDjJ/yQ/LSDl861Jnj4MT+wbMR8HrKOtRYNJSqzU4VixUENT+nl
p12GiCM+xlVzz36T2rFYKylXO8/xS+3SHWCVIMhenTL1sGrbjZUluELgWPcpaTmNu3NUjGzCodZT
FFZJNz4KreusviWdv1JBD24qy6ZSQjBeYtuiQtz+16IC/SwUnNdg7nTNVhwsFzMsXmer5/DRpfFi
26CvXQ56A5/TgOCFgq/tiAkmrBqBwvqS4+YRQxNe3rC0TMUvVVQa5oQysxXJgakUl+FbPPX2dZad
jbu6mOxFoicCeGm+PvXeWFUspowr6V7KF//XXXiFHaTPKIrs2D/7HhSkKxNYUU3kgcXdKZ8LHkZu
Nv/A4NTeebnqw39aAyk8sDFeYYlmdgT8GI/rehO7gLXg4g9lFxwIx6VXJfqQUX/L1nOhjEmhWUBT
1nvsIkJvMZcoU6KEcVLpVsE5yLfyej+7Zbi4QxwRdLQ/6R9OU9/GwiAzvytNQM6zWRlFDF6I8BIm
LdGDsEWLtEvu64VrdrrPEQDILwqX1ypcvxXeuGytQ9AWwhOGkYSa5CAHe/EMu05p0G98Kpk1RR6T
kwVpdS1zvjoIro0HSfbR5b//Dh2shbulqPo0eOgdPEPwx8WoKKXbZ9xXOtbmyJvf0JAxO1PrjFTh
LkxzwU+dAE1B/z9RKQZ/jyWsHGqQCkqsqNrLPr/frGxDICl/+gV8LYbUJt9IJEAG6pD+nR8qZwUV
s7ZgMXi0UkI82rG0y38OQwNtv2v8C7fRGi5VuX6aImRN8nfotrmWY1QoIwnksS3l4zO9gxgds/Hu
S/fB0iA9fp9ac8svRFxP3bjvmGkc7BPoLuPXjK8g/Jc9xRRYEENgihbuoWBKIXpEPI3/xOwwJPvd
34zzg6ao9IbxPJRETlS3MYCUGedwQStA3mRThpnqJRkjBijgm2irHico/3/0PuxDu0WbkMA+mIIG
zuh1iqNb7n7ORxovqc06DnLWZh6AD1PMeU0LLN5xskBNO+ErnphOEeCzrGNnhBogKERGvKg+pVOp
T87B54gRAhHQ+ixOkvcA23z/8yqmv9T6q0lcL8TTtH386//MlDVew+6mxVACTJlFc0Ekk0JHjd0I
e5wC9O2lslCgt/C3Rdt+r9EdxJ34FK2mCnMWb+H9hqE4EyuUXwYQb1pjnZIVxNWJtqJl/2S+er4Q
Liu72EIxZCeAwnxYHY7JxxBN04YzzazJNht+evuHmwIntTtVzZIRV9ei5oBm+Gf8/hQYwvzybavo
7CANrNO4+k4KAJdbWd4MzdG9ct9+b5GRpmAfsCVVRayubMcmr/vz8hW80/Z8rQYYuxBdKOj58nAf
wc3bbS52G55KKTsuTuHdNk/y3rZV5J5hpMh/uNPJsv+v+BxS1iSU7IgBnyE7UvSj+ETBq0cs7O+9
deZlelTGBVPPQMktN5K8uj5OcjC+WLvIzZw0XGm9y+sHFqNZHlGDUJTr3QDc2jIt+a8DHLtqfrJ0
SVxaDNi2F16zcM3IhTUbStQ6Aj+Yn427AaEXoeZNlKQ0BeSvrWA2STD4CDs9u1fZpbfxfI642F4V
AjumKfKQLNgW/ZBO2+gfqodu/WvcwQ6SbhzwS9Dhq0mV3OzZlgYDTT8XxZSaRsCPJrwsLusXHMW4
yIYff7lKM39wAZ9vxZzr56DTOr1J0C3nRiYc5HiXa3g0g3gybigfjzNN9X382Me0ILhNp7jjHtAf
9eLnULJwar2vZjK6KfyDAUXxCf5DrvZ1nDsoka0fKzKxZN9vSZ43RGnaL8ULOHpPTRrxn6pk2/jh
uWvytyQtM+RTm1mYgRO7tJFFIhWc/wWIY2tUmP6xES+EIC8fDrsyXz8/+ZEtqnEIpkZRAa+nOPuI
69XqS9mgkfyE/Wbn+hpk0eLyNN4jV50pCWeWOlRi7FlBN4ot6lSIr8ir3vzd46epSUtfl+mBk+wz
zk5Fl0ncS9Ca6ywMFsktnuWQk+todS/Z1ZBjEV8f9qFVkV3yAt574Xmk1dS8APVuBYMLFydAtHR6
18xaa9YDyR8sGLJb7ptgu3+UywpsZ4DBCPi4KjNDrer+vilxjc7ujnwCGnVBI4RxCG2ZFOG2C84D
cEx7YTpuPmj8NeR9Yl2X7nwj43YDfgi9Tev2G0RSmDniyMe65oGtnrRnleCTuL5NrqvB9ec9unEb
/pGHRNpmIcAUor16k7dpxveuHJZkcnfb5MEXlczFOjd+M1C4aX0VbNNhFd9g47WcANeSXZJY6RcU
wS6kNKy5d4bDQeVbYAbkSYuPCnrsUA1vR51nBATvnkEsLiydPVMQ941PjSn+OAH/XIVAdquLkHD2
YQM72Ajqabvliw5eLeW3q9bQTSC52otLszqTw9/mzjWVMPTC0kTVdZ1w7zTUjnE9yGcRwjCSrAd7
0RJufnHxpksmxLh6M28hyAuNBY80KswNUD9JfZS0feRWcWo3cFZErig81uR43wi9BGVh8/N3Woq3
8qmM5JSeMU7TcsJIhFw8/K/U2zV53W7pLzef2qoPOhwZs4ghzMX9DPWFzdhoAFmeQrkpyI1b/aRz
siLRJEjcOxuG0nfCwWlhI5GMJ2nZ+Pte61e/eWyUG8hLixhajebYO3J0r3Q56J7BMQlRo0aFp8i2
nAfi5hsL1HJIJ8Pf0oOOl2PuYz84S2MgVCiBYR7qeSiTLMMs9lCIshpw/Pm6HyOqcDximrpuapYP
73AlO3nvEfpTSTmHPsxDZHthJxFT63nl4VglnREQuiefYK3Zmexqi6Uf+0HQzuDomclHQI+Id2Kp
PzB4bhYJgU5JQteUKu0Yz0FE9D1e22k3cBGf/P4fiqWoTBRg98r57nGrn1M3DTvNtWEevRtxD8wI
T+iILwqHMySzpOkU47sZoQ1Z1RDYpK/oGj/ukaGGjTCQ7Bd2Qtc3hYyw2M74f9BnXemzLeGtLG/S
VM7rWMVEb+lJbS0RYahHGHpAtkO91mZUPcoN/X5GD7f9oU4aRWwmL9F1Vv3vvfamhoERiF7Afjw7
zTR03GxYNYtiT3DXpfINogFAP5QSvzjSPo9m5HRsk/dtQ0evRpNBuBIlMtBzsNEB8fOZepKMUAsl
8s2BGJxR2tyFFEU8HbIKaODGWDmeFw9+ic06xc/WcabmeMC7RSUt4kBTkPYJ2MnreA/EUQ8X1snI
im+cvGNjwb6nYvhIuFQN+aaSFZ4oyCf48OxkeVH8Cd+OtlrQHMX4lZPa2+crawFyjsz4i2/QqPT8
d++ghD5Glg61fQG0eUA9cjufL8bvFRVdO1/kYRd090piDLxq2LbRNPIP74EzuH4NxPP4kzATlF2N
dEEqb9t3GvcqzmSik7rxl/5izR6O6XtsuHJXu6jfHECB/48afJ5UGrCYqFc+RpbjtZjPAxDtARcs
ZZb0y/UmItk9dtQM4JA3oYGZdzukuFUHIGM06w0jd3S8Dk49XV531zqrzMLaYinguVOFfvOFGzFy
cZLrs4njoRhbwlCHLhcqxg13qbkmaKpqQIrkrcF9C7vT/wS943QKz9cbBBW//9RyPa4ZkxzTE/x6
s2LwbCDxQxivEpX6sbEMzxrA1RBAWUaxdvjj+eyU985JePyCxemIGKzuMHfiPCtMVmmWqmz/LOum
IOyrGH2kEuhL3lp8lMCCH4lQmU4v91SbjojxQtm/nwjVGXIqB3OCxj34aCndwzLLhiW0u7u8xNZq
LZzDZ28H9zhw2IWwJPjcE33lxaBlPPntSbJbgXXkjFxCZAOdZY4MjUNIM9zsg5LJN1EtiQ4jhggg
dbtj6wy5ztx4PmCeB30aDvXclOs23nS5P5z7ASGD8Qn8JcR7deLHT+Z3Mx6uhaNJA26Thbbm7/zh
ldXrLtF8FzJdnk7YFoQjrOdT1VJU2OKJOWb8D4ZrvYfyIQ7Y/xVAh4NH/UJU+T9xKEmlyRJE6hm2
Yt7jDr6lq5rmWMQ4LMDj21Kwx7NSND2Na4Z2dHmX6LmuRez+fg+8EQMJRus8ixOZXwdqOSrcSrxw
umh6GJf2NWKvd/98dgX5xI24TlLeKKdC2C1KUT80kC6TkOGpYlxPBkPew8cIwNNSho9C+d+8VIgl
/55xghpvIHzJvVgbLrbNgu9dradmGdsvgqywKEL8BK5lzik7HxkSFWyKZEHDbzkBjpuIuC48/7g5
SS2T6fSQEfbipZBFbhSltFcl76q/cCI1uF1dqkSeqMdBXr3Dbgm/t6ah8G0c6LvPGeaehxGzi1Rp
59xQTm5I9izEWf7quCBCUCRNcHkk0Wof2w4THfcn7GQyaijChyh3mjdL3RZS4cFG2sJhdhIXEFQ2
cfvUWZ56/Wjf80xf/zqtRXwsG4aHiZYx2HnifOdn648NO7zBaHvahYG3KjTai9itiA0Pap97Rmuq
BShytW6mwtVJRzH82ZJiqttVvj/JLvYzVhFY536zaUB3mWtx3+TLcqry4ZZy1HLicu3oiJR1vx2v
SwWhg0AoS/lM56nmjupiLRn0nO0ZUMrGOz4mTl3In5gNVLzRp+iovQK91y0teyhX/0c/h5AhDrb5
9UBgqkU1L0XLjkai0ZlvrAMdEJlxWPHA7LvKcnaMPz8j9XCHmVXTPTA8v5Jpju+pKUEk8FgX6kpB
cLGsAB3E3Iqz0ryGyNUJNBTQAT26fHQPRcdWkJ13zNd7VU0l820b8+Rzul5vnnItmFHAV2BzIr3a
ke4iEmi+i756vhuCbTIQkU5vTqubF/L8vxXOK2oESbjZueWgK27benm2s1yoLv0Mn9F4340vyzOV
zLX5s9BGrq6lRr2pkGDuON7CUzrsCY5+FPZ97MvL7Tp5kn25YgDcCx3KcQnKBZgRu+KwRNtsQcKX
Xh+RPjdb1+rXi/pFESxu8UYuyLNNLs+syM7wogsBTX03s3xn+ieUstU1eWgxHLy+j8V4j+DPOzT1
+ixNmo8GQEb3WL+RlhA8WjuHzpRVcqUdgT7buHnZTiwc/8JolTdAN1ln3TWJBP3DUHTH0MwZeSjg
nz1rZtejSr56LI4bWjej/nYZPK1D77OmfbOkg2T8/yMQQ1oZglr/LccpUz3nOQu12ZZeHm62xFU6
yvzgpCjEIsJh2DN0ZzicIhvg9ihr4tIPD0JFFA1h52hZTet9ioUR8yVa8zJhGHSQaNlzW8dtMLpt
Fw1ItHKlikibgnJ2d4+LU2LMRze6pg5obljT5KO94EJQO3Zd2o+O00HBFAxJWbSKXQiZes9zz2Ok
hP6ZDrsi7taCHHZLhH4vEF6EcX/3FLnHvPgvUzNKqppHIPAawygZH1n7NNYGh8vA57YwlvqOj+Ab
8ZB1wzfnYoBo4y3fM3PM1GppWeSpM3OOdAwBOxoivn+vR0QERwtxlV/6MBUPHsqQwZgzAfEXGwcu
bMN4oErrq4PkZ/xKGS+BqEJMlgTpN43IUTMkNn5fQJ3h9aACGquhEofNc4xWyweCClCw4QqPW7rS
sVBxVQ8lMD4uN8ucTpeVrcFoNUD+QgW/saUd4Dww1zZDWuskpmV5TmfjI2oOrdmG+1i2+chsSSRc
0KjHXCRNfakjKyXxte71jw4jsAGnZ8Wwoq+yEmx4WozOhbuFfKxHkFX2+s2jgQXIquJosRa8wG+H
sXIt6Lr3WXhN7olnu3KtZJMwQ0EzZjJ9WEF+yWJYasGMmQZR5PEKZTr6dLP+lRMmu5D4043VOOOW
d9OiHul5hjS71OmI8MR0vgV9fgBemqzdAsDWnF73i/2MdmUJrNChx0lgXTs8Lk3xFywHaQRVTpN7
1xyyJTZFqCIMXSGEtZd90PPzHSwwpmiY5NmRATJABpIgH4BEqYmybVzvhpgZvfLmOC3KBLRV3QmM
oXblmQ7bRFwEAT2/XaEF6VNHmSCAy7EGfqlN7lxvb2Hzwo/fFTsUCSqDEwv3d9IKLaf/x1eEA/xD
16kcn8IU80gGpRzavUlceo9bhpvVc7yzvC3az8dhLs/qCdLfrjxWJS1rWaJKFVGOXWg9ietAdzNy
ulW9cMPv3DNOTuK68l03F+ww2yxaBBm3f0rd2qfgLlun0rb3MYqv98ba6tvrIZtG/AGtS6gJ2Y4r
TvcZWkjeFFHWsDyde6nMvsiPxitUD+1S0By4Z8KBazH6h3rWd4bncJJUnXsXpbm4UwavV4VYAv4J
kxONaiDKsMJFRyqS18kzAnPCwr+msUQLuLIPmGCRhO7DzlkmcPraMtLTSjBu7DsWVlusvq2e4AwW
kAJuloonpIMG91v1FZ4Bt+HEFCX+ogvOi2gLbno7bzguo8BOAb9fk7Yoa9qbcYM9V3yyec6Vl9Do
0C+wHDWGqGWT5fJT3m953SvT2fdjzlp/gsM2cz6ksDVFEzSVt0BvbAulZrsqqWEtygmCLNicdwbC
kS2m9ghQ2QtwPSPG5M0BRaXajz+Q+tq+Fms0OChvCpRQgEjrecsQHEKqh1aSsXbSFMvxBMTgrW/s
0uaF3IweWRXS+HkSueIZpC72EC1kUKkoIskKt/8s34zvy+G/DKy2xvi9QA3WK57OC3IujL2eDfDX
GDiy3CHj2MjFp6QBjlD3VIf9dsSIIOvPPc91OaYZyQxeNdmxjIEGwLbO7KfVCZmp7GrDh8O22GrU
s4EtCXZNmEWj5TSFrCgRhJVdHrwGVM3o09BjnRm4LyI/JfMw1aBbKAZi7tXtBSY6e/iOMHCMUBYx
jAvqCXn7rEF49dkxhHdLEbiPizm1tPF1uAE+Yn0iV+M+ZvChrXUOea+tZR97eGcS6A4aI9Vp13wc
MjfVrDSGr/XIpmGF12lLjBW5eE0ODPTqK1gfLRQe7CQpkp7CyRYbq8tQa2UWSVW3awTMQAZDEEJ9
o48uHfCYcJwdq3p4KDQrjKhDEiFakRsxA/SBANqf3MGVY+M/HpOl3dflUpPXsMLF3CR41JAwU43I
rOWSkTJbb6Xhry0199hlzl8ZLT0kTPElL4BrMpKXjcuOPhAxL4a3oveWIeirpW+iYqXF8RNv16jC
MMu30D4Nrp0CeGfdXuigSoklGym9s3ieYzz1bxk2LEA4ClCv1DhaajyLThF3z4iIZzoGTVPHpddF
LaPjiAXDxKHe5YEVG06c9HFzCOBfeY1m6G62/YGMpwvE278dQ4jFdvwXHiKuAflxzo7HlUb6xio3
kuGjnv7GAIwEDIAlhT+tOpmYt4zfm/h3iDid61DlI96p3Lmw4cR8+pEYgBmLtJ6/KOJUq5I/h+W6
xkQ3/K9W7JQKET532bOSpomrRtP9pf2YKTJuUcLZLGGabACmJO2CF8x6SqtAI6NYpCIt+TjQEOM7
XhtcdiHdiodjksVu7EsgqawEpclggh9C/AJZTltVMS0rODUGk0ahdzsbD84eDn4g5Tkbgf9nDS0n
6XeY6pMUX44HCYAK6ujfq1bpx7qg+WUzfI4sWcc0I/3zlxP7iV0TlDfzvNY7mcwt98xszsNIaqa2
3foaUAkKX7bDBeLbFxJek88XKh6EjsViZPhRFXhwrvRNbgpODG34mgY79QJGgN8fSNF8o/lfsOOv
xYSIPxk62PS9BgaMEs8+WiVRofpJnri3aekdYd3DKKTBVRCly6WSKG6uAUnsK6aq112cFYqz7Li2
dm3QkA633MMH0GQr7i4HL2QSG93JBnOMvVYcQ7WN/0Uh4aewirIHpcuXJUDB16Pin8FynemsLhpI
vfZzzUPhF2WHQc9O0B7+b3SYoTHQE9sBze58060WeO2zXwv7oBM7jLh6Z1BmlRK+Mt9yR6b1viLi
KcfokLKPAhWFEBqWt9C/S4B78NiCpxF20zB1g2ZatCT0r1ToCHBPtBb8jybwKfSoQph9114ZIooN
wuNbNY9s3w14kVud4j+hQ+0ovAg4QXzBr3Ny+jylfbQGPCZFkpaQN1NM/2IbuvHc0B9ISf8uKjJr
fWOkjrYVpsJKXlwZlZTwu6J++xza0/l/ThO61uVMQDaQbJZZmXGfz5ICYn3yUOCkOHfEY4X3vJnm
zFp163uOE/fYXJ3fsBq3miGsCvxXuV6EV0mujFBKlCSF2dv/vycGmTJANHWpk/rH4SS1YMhKAY1w
QuKkh8RC29Q4fONWL7NSHac6tjtRWnKEQdarV54TflfH4Mof2Xffqiotim+sQVCg8MfhuOR3ggDM
BEbS/Gyce5MD95IkvVyirO1+ECiiUDgXiDicw/tx+UbN0RxFwW7YD1zz9Q/lqzi8OliKEXQcLbe3
jwZDxdcvWJE/HsKrApafJY4Tcqzxm60SAs3+QpIAlw+I9fODe0yQdtX13wVb0+sKtsFKENbzhCai
DP0DELZ0ex1ceswnf8skkretZt7Aq03YShSoOHxTnf4fP+8UOuC+brHUZt6Ob5PQZ55tSm4QzAl1
eu3vJ2T0m+8YnAXe4i9Bv+OjOaQHUHIAY1pxgO5UQV+F0JcVbtePWVWD37OdOu1nb3K/uAlIEQgR
KA25PhDR+ogOzT4c7Q4kOjaXm4trI2MERpdlH5EHe+WTmkGlEaplyYaVhCbrfSn/jue0pvi+pk/a
YCtOcQ6ry8JqBI9WRY2lSqHvV3sDImiTVUG+7dAvODvrHs0zAXVn3eLLoXbb0aeNmlG0X54fHK+E
dGN+Jk76gBWlkkH8QkvC0DNTSmnOye9lt+tMBqjWiQkHcNhMXK9hbmll3zopBfwTvCyOb9z+BW8L
3IBDzj0O9UvkGSwhO7mRl+h1l+7FlxaTwY4RVGOVrOMldMDrLnhOO6txb7wR6Wghnf1yw9Ne5BMa
FeBfKHtJL9mNjP6ayr8jDSNyaJ/Xm7I16C+09IgGXhV2konatc6NoCPcPrIgVUfm6/y34+Z3P5rF
nCdaYalB0PeimToSSnPAapQMD9RDV2HLPdOe9sDpEkW4LxpolwIsdgGJvVt2UAz3+wQA8dnFPbSt
5gCo8QGNP2QKihhLwFZmwZUEJIKMLb7xCleXSFQ3Usm82Rz6LiG2mpwKVAShXjBRVAXCIAK0B/iw
DtQN4YjOmI6bQsjXih7AaUhfhOxBmcb/oWQ8gy8ncKVcgT6pWyJ4FJ8cnfdCXLH+dx6uHwCnPHaC
exBfl2cQlEQFcRBHSgcDoN4c1QYKm8YFH4+hLX8TCQm6IWBTBh8PZ6dEuzHPOLHfo6xhKIIThhrC
sAFogjMXPYTc4iFv3NsPCOug+CiNiKkU7lbOLOYYInXiikJUnmaqPuIfYGFb9/SwBQmpqsLByoLR
NV+8NWAJ4egRbIAqfYnV9lYWWJckt6ru1LciN0+PSEMlk3cpA6BHi+ufcfq6XBspEoZ/DmM9g5xd
EJmcFWBsOio1c/BgjQQTW+bRlv4ogn1V7kIPu5+RVi7XK9sYl2hPyvXvBPNCOwYkGx5hc59XLaT0
akeKNffhi9kNLVVy03fFW0UU02sx9oYNkV3yH5fXbs2Gr+Hl9AIvM5muZcLT9wHdaaXL5RELq4i/
R7Kj3T0C7AN0uMvVjpaZcFrj4MQLTXIkG1ceTiSxx0kzIGnzG8LfXPIanTANeiawmudTNwEuu0/m
pEWlXKi+Rc/KUsNwXWOpE/MSuiFx7VX3NCq+DpqSGBwtD9Zan+xNmN1QW08WbFxSoHKwK7meSkmd
x76iTv2qkSkhBkONttw9WIz79evAGXshW4vFqMirgTL4YR+ovmbC1tmJq5F52kOeC+a/vlBuHC9Q
O55VUd1jZX9CmBupAD/H0Af/zeSUcCzJFss7O6fueBDdYVKjFd054E51DAWf5YS5W/Qp1cVhQIK3
++2YuplOkoAvuJijZ9g/Y08D2t4ScuxUGNf8SjNSMpV0xmkRLVb5jaF+mgf7qJ6dVc+LYNt50k22
c+1pWJ+PnJzWqeaDeeO1lXn1E9k1EBXWE5ChkEuEKTIEerHurxOiujXAzhZWe4l3mJj/lXmCnY7m
QqBn5JcR+SdK5q7TEjNd9hnnCsvWYFbW/Xpv7WSp6gwxxHaT4l+VtzBh/dkLsm06DUllVtEcE0fL
SExqqWh6SufJStty3FIvv41UYQKOslIskSeZ6oIX1k8CxyCp0xqhg6zzkKkOAf6pdD5Ws8dsVsl3
z7Bop8c9rA0YLg04KO5lfXiis5aHqrLEJzerommvAzoVmTBjrpndZwJEh60O5b1oTwhi5gHiVl7S
ol0hxk4S6Vls2HR3pyqhdBLqSXDAeeKTp+BTawZjegc2MufmsAx2KfOcHGFfaohF67gPPU6VwmzB
pKBgqc9ivZmUFBghLsgaAR8P3O/fkE2KqOXqiC3fUb7fLoSPqHU86IgT2R/Trx2xUgwhqYLLLRco
TGZdqwjOBPa/4u5ICL5bXKwegFl9s+zSlgTYTS+Wt4VFsiI6BSqwOy3n3EMHkDxNqNlhJUOJMDlL
bOtrg0yIQkt9e2ZMfQdeQ+7FM56dw8rhQQHRnc1mHSIaZE0XlTwHnW2lZCSkyV247SAtO7OOSHJU
yXpCIWX56qFRCbOSTLuMZAPdF5u3/HJC8lqlNmd/CEmwIgv3Hf7iATAFTt1izNNMM/QwpbuIeWWd
pmBK+Vgt2ENOwysWYSP8K73XBKatzeSJlkXI5hioZjqgs4ZyO55Qpv1mnTSEd+vwVM83oqpfj648
RJP5tpJOoR/ksBgM3UNKc9mCCCueZ1DcJ3JDvzAumArMyjnzmmuHGINHlSiaVh0O+PbiSKu2LakL
+kr2R3Pk+z8w5RxbAJ91ziSRaEfQZTz+mlOjgwsx+QUAkw++w7B3785QlcFmdxHpdmmr0kaor6Wl
WjjBXYuyV3xZ6oLFPBQM4JEQbLKv8wHRcW70cVmJ2JnENlnmHAhGKhRj0QaeSHLdeuQbP6DhrfCt
8qtYSty9cPwPMIPk5FS5krfB3IXfW7W2RVIZa6lQxYW9twIbaqiurWPX52jzwVYJx/DY/XwLlmju
DnhktQhMT/findtT15k6KovS0ltLyOv46tRTIrw08lNLQ3nDtn7z+2YpU62iFqe+MZSC+eN7j+Yo
k2DPyltBYa0QgUWBuWYLObSoyromolZmjADTRlA8Yb+PSmnldFul/jNuXBV/pBWdXlZl1/VBggQv
yA7tNqxsVzhGQAB9Cv4MJhXHOsTZ5VMyTPxG0fIxJbyYwR570c925aATBVM7FxeVIDW2gTpTXchZ
Jq1kr3lnXeQk49PURVyOgl/jisuH+xr+f1w7kiFNYQcorBgPS5Nvmbbi5tdWSp4L7Hp8Y2/nIeQy
ipqZhHP4iBzRwWt0IVL8p3PNGTS23BYszyIFApa7tPQBssdHY6TBjZehVsU+/lxc6KQmetskS34x
M5ziXk4hbHo4ZMOXISv61aGxUzgA/TwjDq8urjW8MPTKJ1vF2Nr4zT+f1S3j7FjRzzKJ451sPujw
PrsTFSs5A1VFy3Rb4PDQCqrljNl1DyVfEOEId2KIl17GOdNfmpr8ebNQRP+6JpgR0zWngxwesAl+
FT/W+3gF4zQ+qKiKdwAmPKm+uGgj01l1//8Q8spPxnLrX/0O0k+GAvhbNl0LIu947ojOpEeKfaEs
Gg1GDcyvcL3ElFSLCdbJFGFPsZUcUc7pe0HCVpidANnbrE0+N2JxaNGIxxpRoUplxvuReaW9KIqq
GYIwVvEW+KpOHGOcObc39Jc5Aj719pGCXcpD1Sb8IYry9vwHSvkRqYNzZwUQdIJVngoKbAFxm4nq
KzsAbT0Du3i/bj4nG9Gi4SG+ACXKlacKOqJCdOiuJqj5fkJZBdM8b8bRQMVrVgaeBE75iKjQDHvx
E+tTRXtC27rpOBEvtq9eVePJP6joE4VdRhnVpJcCMXbQkD4WbcnMrQWQDTnbiaeoN4OufZsG/4HH
GEyttaBzCOekEUWiQIh7prquNkD7OY1P5cgzeUGlhs/BJmJhhsNxuzWE1YcuaElWgLWyoMa86HOb
7AIdUQxYeqqqfJqdFEpyF5pHAco7UH8+X54h1lfoF1sfM7chBU2GHBRuvOA/ZD/5gVKCjtvISFPC
L3JjGhPAhhwxtfZe/X6u0mNOMIJyJeCOKt34cO0NdwWZqi6omv7as0BuHzTj3MvhMcRjjFp3WeN9
qYcMT3D2zd797gaBxwwSbrZVUsxGovNfQT6yGDxCRCHATZQchulqO2/J86LY8TyLIZHczuJewFbx
v94tCqzDry7Zla8Aesi5QghIdUUfv4o655/+itOTJgwL9SyUMOc1Sfutt48pmijkprhqa+GN0rtl
aMHnZNrNdYR0/dlklm8CRmb1/lZoj9nvmhVVOAiRAyTcJLbnNIM/ioj3aYjwhINq3NhG8H7Poot5
OH5dfXM2Yy8LbugSD50U5VO9pmmNl2sH/8Vrk/ySp4vY0nKRymJpb9o0ABmpRABd3w9iymCjS/nW
FhtU5nytkBykFgAvnt6woqKKZK+X3QahGvP96Ubhwz1HrONYnpFctzJn8vERZs2YtMsvdiSPwvyl
OdCYfOZsCon/EXSba2HTilAFO+mBAkULUusZTGWRYUL7e6XriMfyNUI6E0pRUJjaaOPeechc5rn5
oPINz8IvAbf8EQFvNTZtRNVm0G6iwZadEo6xS29Pam0eHZiRwfPwyydei1ZE436V5M+4kGTApvKQ
Yesr7Ry/vw3X9XTOOPTaqzn1THf18jFiiH6sOecbtX2JV1bUQUjf96GhobHCh7mjB8vftV3dCoaw
VdrfpvU2Y124+iY07H6bXXys/FJKJT16hPrP/ag3YqaEdvfkQ9lfN0kPNdC7zyftt1XC2mj6o0mM
K7o2lYna4vH/wGJCQtPcsrnJHGYVVDkbZtKa1sVG3WQq6gJgbm3Or10FK4pt/ANto7sj39AvcwQ0
1ZO1aZylJa0gI7KgwVTkqdvQHQCx/plxGbvYVR4WSUVhWyvMaoa9vuwl5+7eNR+D0M4qOqXLkgud
+6W8ph6DoPt8swzX5iDF8Rk8zYdPV/AV56zCXRMRkraFkTUPK88Aao/hzMtKrRA2aOM5VrbX0L+s
KW5YEMKxIU4f9E8eikjbCQZIfgYcs1DrPn/DFUQ1BX6kcBOXKKS6TCnAQ4bV4pkM6Q/60yU7GD6K
O2v4W4Ngb7KCPF3EcHyBVzq2+bG7oE9FW8w+IsnYWiBUb7JW6oaYfIeKTG73XBrnTzoRMUGvGMYQ
H/DLSKqxXEthk9tRaHjaitHaNXQQ99YO8h1ZiI9jbSkL6+FPEvYFkSv0lFw23Go+m/M/6vw/wGNZ
n2UQo/K57qdemhAmEQuBdWCknC+XidRuWeApzTS5HtCXTzlf9oRXne/liwOe+oir0h4J20cBAoID
mAmBLt6H8cnqBZm8goqgIsbXSIxIbMGhOJab5F8Ntc2rE1ovkHAP1rwRsQ5pFEw5MbW31sgUxwGC
MDBhYEhCEXnUeA2g0MT8cNa9xGETo7iagXqUESkbYEic+FwCmxId0fHMjMbzJRESrPQGgnJZCNfJ
Yjwzjbs2l8woSi2toeoiaDjgkH/jkIq4ZYU+zZGYqAFLB0ScM4pFjIPdXyb/n+ASZ95lrHOzf6Bt
OaWAX38hNYXGBH96Xisr5Pe1TRjFxxJ/I1QXHKsoesT0QHdxW6lz/rkMI14ETYrw3twulHCp351J
RxyJ2U59bY/9a+kiJSkPed4YgkNB3L7qMQsBvQCIhxI+Ksp5Aye+e75zd1d0oR5lCdYbqMMdCve3
eztgScCzMiY6N94ChqqskUYDz+qE88qYMxxPwM8t9HnWPIFbAp5Qu5aI3uUdEEzIizZ6haej1HZd
GTOqEN3Km89jUhx/KMh4b3wNcZmHpCYtDFadDreTEkUx6kJOGiicNgVZOb4Xby1YKw4gnW3AJcm/
XzJEkiNhUbWBYBi2XCTFKONwKa4O6eO7I/Xff6tK7+epcCioA6w516uRp9Q7KKp9iTNn8IH81t2C
UKbJyDDMEXtAZbvGBc6+U/T8t5bubMa6ZXbv1kobhVQ7c6Mh//nEBGNWU+eBo+KH7EuGZBRJ3oeQ
WaDoYtR03y/OVVkdL3T96FyWn+9XaeIypum/WoYCx18tsB+5cd5cPBSkePqruv9eyFjeeIZFK7S0
/JlP+grXpZ5MzQK1hJlm7cHFRNupefrDGcia55E4MjbJxnbBxhcLVchuWP7dJKNota0Fgo2G73JF
RT+eFNkj5eyQmDWlD3xiZcTJiY7nHzg68S99bB0zAXCtNdmdpQEBa0TGVLylvfuAWax7NxZltIXG
9Yy9/LHCQ1C3/CBNBXRUaWFdDLEZDbsJNTzOMXRwyd8217WEnLScuwgt9P7AAwqnaOEhRGtpO7Cy
NftDS24gfAWQoDmS0K2TzGhM3eKFVYC4cvFJQdXZZISQDXITmX3ISmJ5uBiBCh5bzSuYvd0CXjQZ
NXchgGsvbqDj2jKbbI7Rbz2+pvhL7nV2TuHhdMnICBPFssfrPj3W+WPC2dE9XRUDnb6Wu2LY9kAn
yqdi0+waJ/wY/0Ie5qkaIPlwWJQHZwQFVgVT1WO//Dcu2JaIDgCB/62//D2T6Vt+IXZ5/Zy5BBfk
B4pmZF47oklIf7A/2xqjfoajA3MvZIFl01EuZP1K689BNWK+k0H7+WPJCCk79qIG/zpwHqQ/P/Md
03SeRcJzU5E0Vvs3OfZgYWlHdsITBmGkFe1jeGwwoLdtI2RTmr1yOM3EVoLWDJqHZYcjmr2+Mr+7
tOO6zwG7nWmN+bF56+kJzosJ+l+LrvVAZ0BzFH6bgt17n73VFYVyVfvgs2935imV6bsW8LhrSmea
xSKFkMCxD4z2oDklAbStStFs1zpZlCzthWaS9EC24lq951KRlySXL+x3Bk9Xr/8YiVu4fxPxoYjy
p4O3rpN6/oNrcw8k9kIxesv6K3RJFctY6PYrujU0fbg3FlcxYlSNlScFsq8X9hYPejItsxROKint
WxhXcyPwUmPSpQwC5M5Wt9q5LgnqFM22m5nOqVQgc++D8qKyMyrGNzNBOFejkCQw7b/LJsgfZZG5
hT3/vNxbcsc9N13AEDQ2UdZtKgkGqLV8o0Kx6VtvvCQzP8Q6Vg1fxSTpxkYbXs+HfLsrt33l69KS
u4mjOtW+R19/N/ZWsCfQzNgsxe1geG6eUxJ5QvOjAx/whTS4RgymxeEFOh4kLUts7yjt/XEermhZ
Qpk/9l9Ld4Ggmh1LVuc+/dE118WFVykWIUAlaxRKZ/7zMQYiO+VwtOVCdFNP7V/9PSXrVKKruyX6
+8lJsZQpj2+4qduBgyCSFdBDarwYK2tfS7xLxstvJ7s/wWvJ7dnQoZEA9L3xvbSslTCJtIsPOgTP
tN/fqtvtF4rK40yy0DtTjAuNXlvguDyWRcXLnz8biWswhOy4D+1mNWkPGhdW48jbHH7b901wli4p
uEWnvmdknYZfEebaFWex/g+TTcdyYwxj5nn9DpecPT30dC2a/kxf8u9d8nsr703keEZJRdOiwH5Y
C7s4oTuNWErsgIuHoQIoPoBNtZOjryKqfgeSPtDtaK4wRCt+Ji8vae0toDmIlOOAWp48Pk7RkrvH
nKn1V2bmROUybaus9tcB3NdITB9brsDoX2amlasAlssWd0tucvHrteByJSvCO+BNyOH+oMygFVdY
JLWc3lN6LONmHerXpQi8PeDdJAqERCU/LOY8Hqgrf6hmnjypdcIWb7WcwmpqMFOy1OQbYIL2mmGn
Rdo4LJBSF/ejKkwQXgmFIg4BVPB3f1rSwm5e+8I2RW0+Jlc2t8V7gcNO9uH4zmLeR59FEgrC5Nxy
JRbZjnOhQK8dXv/DqQHss/RT2NyBJ3KyRLyxxJXgnqkvCdN4Zp1YETMVLdwwgJawPrq8uRCh9sKT
NMlhLO5V4qS9rV54Lw5C1ADor5cXXX2DErTUtohrjkxfkc3Cxaq5snDIJmRO29ZlLd0HPRBODWxz
sLNosL97Jl5ZdjizzjMvS9f2+rPl9H1GEvLN18FM7rmhXyj6fYJ9FdVJe8PeY3h/6sPcC9WEh3Fp
nozx6m3ZKLozjNF18FFZzUmuxHny2emHnTDV75/fbZQA2XghfSZ0pXzwNqJhHVecApLUuCziWTKx
EnpLn9XuNbhEVrnwUO1F5olFiNnTP/KIr2UrEjb6cCd51k3F9fmXqIqzvNpEb8NcEzWyrf8Zip3I
aff/Q7Cv/pj0952FCsy6tyzLf8Y19XB830AwxeHpYm9qkPxtiRYjevZ1BeCsHVRZSB8LW/RAFJV7
Brrxi+PPkwcU7rPdmqzU747hBv1Jb8nwlIDRnhIqEbzThtRA+EZI4JqgUxgHAzxYWbb8AUiIjIyn
rn5iY3+60JmUSv8LmQQVd2HSKWPA5h9ZM2haUq5I0X+SWwiVWdVcLAT34me7YiwlqjgKFMEVDHtj
KGOD5h5JIWkgBtKFFdoXq1cM+C2bZLwr6f4DnLWKaYbmSSCqQuGvdlPxzWpw866Ozv6l4ZsUB/+d
WQQ4Mzc3KOW3KBT+c0BME1CXZRO4vP2NBWSJCGR/N9kq5K84W4X/Uh3rmC/GbaLttO3R7R1AZqVZ
plp0x0ClTqPNWKWBClSzGZtU0BEx1TSoLs9iMFUAS9riMmqHXQxIGVgODj2QmuXIAH/Wfzirep6t
zp7HQhyIqb6G61cv5+KWIrqs88n7jJTvLeXZeM8mbyCGxFHjFDrVf//tVbkL+vmvaNWUm8IBj2We
KXfFm2DHhDAKWkmxx/xBqFv2j4XFcI9ZWb2GRluJaxN1dcOHTb2p8dl5q1iDNOVa+6zOal+limck
9nu/PdTJNDCIPfrVPwNj2uMJgBAH2tWV2LwKawh5bYkASE31e5G2et+vn9bF/qbdu2ZWSNbTwMXo
rBeCNuvUrWV9Z4afnUUoH5LoK9JWRtyYOrDnHC1zcsEmI7rUDapm3XFVBKZtbINSE+lxz3OZlnm1
/DP8J7vKYju9dScDCgBYZfXTW+cx85r1yERXYr5n0CBzgk8GTHg67JT20pBHyLE4jSsg6DB+9si3
+Mc2XQu2CwyWA0lELh7CZ5U/+nyK4OGQOyJviaeCN2/TalFl6uBR9ATntG8WoGG6++Ahtm8oM1U2
1m/A7JCjM+Msk2gbY4QRtz0lANIkG51NdGb7/59+LlZK45KIuNj/PZtrQVjtYy/kfPcJQnXlH2bE
miBrSg4E6Adpx/8nLmw1Kafa1FEqKnc9O6WwqWga14ldmhVE1WGE2MoNM0ecOcxMS74xkaE6gyMy
QJSyBAXESl/hnyn8nkUQfUna1a9vgledSZBhsIQ6a0QTKX15l/UNYMgu2Nhte44XySzZ+QOe/mTa
ICWUbVKhVz1geNVUz6mkoEslVFrvnmXb/0yaINZl8sDHn9deen/thDcFGdKyca3EEndc4CB1EYCd
JI2N8JjvDWfFEEm52u5qkJ9l/79cIMBS2TfLit9eAqhY3yaf0O7wmYgKB6wJFsv9Fi/rjQ3N1uJ8
kmIoEfQnXlpMzXv8L5aT8Ey/w3ySX/n53BMH/tcjQf+0sGNSoi3c5h2GqwvV8rr3zBZiGN0BKdjk
rvtYzc6GaZGe/YrzYFTq3rTy93Tdja9/bZb/4wb8gS12uhgl6ymucwXOM8BetjolfTUQ9fm7CM4I
ptPu79yj5UNrm+yMn0BrxKiXR7juITQKUGaKBiP03bpdGowom+IHY9vakWtdbWJnt+jJr/xZi8Yp
4Nxdd8awPpWMt1TjMBf95Jr9o1RoJJcSgmaJ40gXKPPeopjIQCXFn9rDWly0+zItwJ7DZw1YjDio
JRRLYoVtcKoCbYu3vxRinn8yaLRhFyFysWnIVAWcm9KcArYgL9TYDYkvF7eZrVmXmMAu3IqE4WFm
oOGcfdKftpguH6F+r2AdmVAwkwq4toX8qyo4WSgyPOgv5oLIJyiB3z4wqcC4KhxVHs5K9Cr0cN1B
dnmOU3iwLB9zrj4ktpconyMCm4wDsDBAEAYXvU/a0i4yrYQkiKYaiSi4glUL9Hzql6arxEugpMq7
GExLfCbUXq1g7eEqelF4WEIIAJjXmwvYfxCJxzn98XSBRc+gyHnIJpHGIR+IklcDnirHwizpzNg7
DkM7x7VFigfiWLvHX53h1lAiz1h1YxDBJoIymgWI3uQdIutBN1GGoCnkIMN1jLnYWSY0hN5tioQn
PumPtKY3u6xsl3yfx+ipmNQr6MkigxtFpLT0dGFjf5GenNiSvduW8yz8n3JSj2ZxCXE0VSbrv/aV
OOqGtBGxHqWADzT2ZEYTCdVK19L/SzY+pG7FHOtvxX0sLVF2By7AfWNrQCArZBrxipKG3+6l3lKU
R51S9G/V1G48idT2iIrtsAy5JuFOhfVZyP9M2dYA62RFxGpJDkz1HDgFvTBn8WbVOiiycZ8Cw8tt
+iNNPQ+7roV6rPzslxl+qbKG7KH/Wu0T80EOM7ihv9wfIVCTCvKQc4MRhjcZ41gXcrD9uTH6BnQY
Fc6I3ZazV95KhHW52h+f8NZ+macgOvOlykmnpvXtzwAEKhodeGWGgIbhUXPVI3GxzN/ih6HL5vZG
kA0iSHc4Sez1AB8g0y/RaPq7Vsq5aAODIEKREVldp90q8vwoywFbFL8hHEZ9h2+riFZioFwssxaG
0xY4X1P8kkiBeFaskwGjVRXJJZUCxaf1+bFKo7uUgrCaj/ZDVyLfskrm20DTdLmpgVMGTpvR9mh8
0c7mBCxfLcb9ap+TOurTe+SKlW4lFd32dsj9P2SUl+1Valz24M6zhir3pPpkzYOE9jYV2grcXtqP
6jhWZAqV9x0JMBo1IZjBUEwy80k9oooyXWdtNRzZVyUU/OXN2bSx3rPGH7GH9jToBKu48XuOLzfY
3JfcMlqWqwCulmVWeT41+Bsy1hOvKcoHRa03zE3J6rn0xXf8ATqUFmLdLrutXTLZS2ZlNjDdSl+d
1CN8mwxwT79+qdhM6zEkBMOVNkhJEGGXae64bZRTUsT3V1iStjOtmmIRqGJxT0LFQaXJdI7i1R9T
56EMA2DesXDFudcI59w8nt+lFk1vj5YH3HEXgpQHUg5zNl0r92V8OsLPI/yP2C4soR1ZYlDZHpk2
y+Ug1ujaUPktyGoXrVycWWe/jHbiaCLc0r3IGiaRrsyWAy+Uz0oq8iKd5TGAUKG0dv6aCL7zBBqS
/edJokWQT2r1vH/raN8ZonaLeb9GEyEdizSr2WexhAXRZ+LR57euEVEJFFd4Vs8BXqeA0sbv1J9i
3mgHwQjayaZNcH6Tv3TUcbkQKco99ZK0ntaqe30lLCYQD9Mdl1yp8L7FC/RJ01xO0cndogFAdqJ1
hh53J2vHsGqJxA/WbnjVXtBDfN6EWYjxiueFai/ATdmGKV/PMdUwyLfIQZ/nckce+LnR4OFCOaZY
E4QTfdR9LSw8YiAyOd1QPar+vwlp64bNWbVemQeEreofN9XA2j0SXus1+4Gy1OVhm0R2U2L7IJgn
pMvOAA6lkO/cwosAXFl38Rsg4HAJbTyMXdwBcoqm/J77P3xiCDzcQRMJCyHvaLb3085CTXUK39U5
pYnaNhemE3Lx+ex6AVwupu9DN1NMb1DIoMijmOxAU36S0zVLyGlbaP8u8a6TRDZ34vU9XV6/CloO
FgTi81Sx0vRnMVPa1XW7vNPbhqsGnV1OGwD5m1pwvELqDyIsKtVxuMLucYAfdVS++HJelC53/z3N
wbREiDXwaA929sCjLE9NrkXtEXAzMJDet74j28vFnDzVi0jpCESvVbavwNwHn601vBZcK0O2aTX2
ByVqSon/pYhqGOxFSRcUaS/SJ4hTb4HV1N8ZA4dLizjx+myDhfgeX4YcA1JwQV6SGps3TIKwUbD3
wO5KX7hgHs14c3xpkZu+4z96cxrS7dezMVqDcRsCwvAnOVhce2IWxzAh66ihJkPEv+G9l5uonS1d
4woQvdNnCpesiwcFbYCdf7RXGF++W63690PWVLXdN+exADtJmmnuV+ZYPcUvieUuotN0ALabNOT5
ZUFkkIzRonCzfHltdpNsGlgCQrS7pLnTW5iSffetk5CrHlCdDg0+wnd7vo5MWiQ0NVnYT44znmij
ZTx8yE9/fodUwA06Q2nk4yZ+y2ciQ9g+TSGbLGSoaAjvZd+iReRf1dJaOL3gY7xJ9fL5+L6dEycB
zbsUqKnlZe/ECsJbZDIF/9NPgt6cPpeEiSxBpIB6gqhd78IPNG9gQTqo/s8Bxx+nHmDT9PuH1uoL
iHqs727Ov8bZbLOkalgMY0qVDQVK8y/uObdIMwv8umP8GykKIohxic5deFx+ymcw5G3a/tNHdS1i
f+LVGNNsumGRFLtBDwvD5ML21MeesPcNVn+AQM3M1L2vqgRm9GGjtuYxyNwbagkCElpiYGoIvh9m
3RlOBI8kK/TYjmA0aGij2fYTAodpGHUCMGy9DeOORT91fkMvlPcVPWtInSrIOsne622DOE8Kp4sf
JNzwn2XKnNfwbgtZQFmhVjVmUSfB4mzTfySW6uNOtcejBlfAqMPcu+zVzugJScHMPf+Veespxa2w
6YSGPpCWT/D8DN/UxE9Ww95TkJ9yhr6uRj83iQo9gFT2ePx3Ioux3JHWEcaYa/vg5JPkT8cqcPM3
ZQpufDAgkjhvFHOljx++gp7oRTX47Pel6sjhsAT+qQGi+s88O//3qxuyRbsbdbmzbN/0ceuMPJvG
AkzZwIvFQRDQGLs1hdPA8jhyD19tjIkJT1dPSz7W51gpDNqFdJVO6SSrFB23iOPakP3xlRkZywM0
dWGOYr8fxQhlGBn9Gy3+2ZMFUnPD3beHZsaWHvhALu8RW7OBmEQHKpmtM5+7hYxMFZ3R+swwScJA
MQZ6Ajm2DX4hGZ/cIqNEwu1CMZiM+bHgRM++FXwebU28L39f4ke1jw+bKUTJHRX+wCansswt80o3
meBidRAfWhVqIPvqE9hsMMRXU+xwnWUhTfGddaeb9tlGhLg5TyVv5FqfIx3GHGdQlL4PKmfCSuXJ
dA4c2CN00yFLvKtbct55NLDDgKRdpS1lqDJUApP+rP8bE5mR+VeH8CT3i53dIeY+rz4Sr6cJ20cY
3injoqS+z3FFaDtb2S2ahCfcPQwQpD2YEPFxq+d2Bhm9sjljy2/yBmOnDPQXc5mk9C4zyVHadtnc
7Bf9oao5yGOUU/fo3BO9MaEshhCq6/w52z/PvdjF+/yhiFD8TPB/c/rbmNwkyIMKC1VlSkrc3B1W
PRp6t9R+DC6y63CXlUIY8ik6XZptqXuD0it47wm/Up5fu09sCukTcBr92sEyutd91TzhpYcffe//
nvcAEqiUvnWDappdTSMXplYnmtsnG/LCv13n13qWE8fc8mGb5uBfloNtX0tAwvqUtbV2Bu3b3mvm
59rarrGVI6SSI65HW857uPvk3ugBvk00qwHsSw0LXyuOCIt0Uq4UNU04Tm1GOVyfe36SWRVUW2nr
EQLiSVCL9gWJVG9fNK5Yw+ZtTgJ83Bd4Hpu7xX+tE4uZgPXnVfiLsVC7bFb0V3G7sOI7s/r6LKJE
aySToi3ogs/ygNf7IbgqK+pCQw0Ifx11viQabaaF7wJRCvikxm2jAfwqiORXUrgBmpcFuj60p565
qb8tZOZ6/M09L3CPmDe/f5BPwedKfUop9mARExvhAjugxGXH4Aca8RSO76tkJq6kSFsKeEgkw1yA
nm+zNpmP40DMxyjnlv4h/GmmLnRAMlYQCfRPiteCNtyQcg2NrEUw00tryg3RRizmXegI/LFgiuSN
OzdJxBnA3g/EElClPZIOpjw8DpryAuK6s20nCs05ySyVlqChU073dxifeNRNrCXPSP2ldsMT9Veo
zEDOF+fewUCqqw3weVWDc2DAObXXELlvDIywivhxbKdLCHyYVPsbc8KDD2fNmwbCuSfoZoP4Bzrz
SS1vcr83kfuqd6Ah+xLMGpo6ECCbJCNmeDD4Rwrj0jycFScVj3nuGw39aE6RLYKYXGkEFA1dxMF2
3ItlRQNoEDfWnBkfaK/89jQ0ESyOTVFPL8IVMIkc3bufqa41ZXLtGaCwjNF1zIAouTTniNe5pzv5
D+cQvbzMpGc7v7l7A1bdFZwg8kpGsdsgB6d/B7PEE/ZPlfp9syZIFX+aRqnkKXlRpBs8aa2f28gk
04sq7Bv92i8Mk2rJiKd22UA+FOMcULQClIYChthyyLFQIVFR1VBZeQhi1wOzN7kof0VUTc0g3rQe
LbqIHSlWioClGhu9D3j/dw6wlbbBoI0Cwj8AYBxCVhtbDPA8SuOAsVN5VwDXWvQaGNLra+VoZDOo
O/X2crDIiB2FKXCQC1IHbUzCnTIa/VaUMs56Dq4fnLLKsjLB4U+9hd1ChFNCg1NFokY9NOwwTYBE
2jD6OKcF3JMPA78gNmSOCLur9O0k7EvGM40kGLjogcuAdi2pvUy/Ht0WcvQQ0Urye6EkQ6aBa80q
RPjbcCbstSUsqPZlyhmEAUAv+noWnhvS1RUe2ibFUlx6gxQZVawm3/ZwooXTLRtz7UqaHL1oZ8F5
UioXySrG8+fn1phhMszexnAa4qxQhmTgshkNcEGrkR1btTa9xllbWhbVeruWPtqQqmN0wC0noJ20
h/Av/X4nXELyBe6dr1evlkonBCWBjUpz3Lawy8ueEltnECUZVuRRR8HeeLkSyzkuvbvnIqZ3U93b
ta/aczGckraUgXOBKhWNwoJ8EssxX7CUAB/qBwvvfjhec7k9c2mdU0BZvOuXxW3k+HmwDzqiNwbs
ryi/MVHF3A6vqYnqClCLJ7+ou8t/fyTiQj5DYPZtMEoK/omg6kEAD48AzKkJ61neNWYWm5sTYJ6v
0ee/aTZ+NNgKJAddkHWcLkd4TkNYmun2VppKnEQvEjLb7Mhi8BA5dm4FfC1g9eMhmNs8shAhGh5o
tf5dBNYqiZh8sCLTCjeWjkh5Zsp7VcPn9QMYZjw=
`protect end_protected

