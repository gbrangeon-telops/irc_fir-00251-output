

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VqgplFNkI2rH3rP35CdiLJAesBBzx3ahYCWVov2QY8pnSpbbPHZzKXALTXuf8Lg9RV/60SesvL5+
Tx0kf3Xi2A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YpVJ/AkbT/7j7nP1FpW0u/1drBu1Ym0xSQcZVVNR2BH9CeGHgikyUixQxXpCsKnhOEb3pzk2wV6b
2udOCqgzaZfDIjjaxTt9/C6XIY+oMyWDycOTnGwR4Bf/A6rFEzTLA91kxNt5/tS1PVy+wjb7FCsa
mgkYj9eNUdtmSsLezko=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pSdvSF3+OBx+pmFIuKYX+lTRtc2CK1xqA/WmTxOA/9c1xuF8tv0giSEc/96tBGsFFqc25YHyYiXZ
gYsCabVJMk2jc2XaKW+XFrRUGrQYLd+QPrzsIggnGqpN1i2vEJ2/57QIQEt4pR4jX78IzCIP9B1I
Mief83M338G9aIgdzONBxsD1Z3XK2M1fqZBI+UT4b8E2guDKnWsCC9f6WqxH/+ijAu2o7kXfkz/w
wH4eaCjn38eBIq4U5maYpwbVxvzCRoB69hlCwEEVDievRmXHouMD407mzOTwKaIkf/tAbFyB6i0D
s5Boa+TiBtHShhLBGBRqGoq+2UpGEaVgj8o3hg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HVe+dxCY+VHrZ/rUbzyWsz5ix04KcDyyUrFaCcS4yZ4GTBKi9GYUFVfTsXMpSX8pxXieZIsbIrAR
8ATsmu7QwmViHDzOMuS6sHzr6e8dC4A3UKQC6xKKwbJdSWPz/il1AOb6t1CcrpGMLBXMZTBj00R6
KptQtwRx2C4sHo/bHEs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gr9tWfnRHlUz7X9jwun0huNacy2IvVfab84T3X/BBntsyGpCEQL6hR0/eLuvmgsVt+peH9UtRKIo
Mx38RlMVlftuoIDUnixeoGaAc4c+4+tb16q3/5V7og6YvplXdBH8LQEEDNM3+H5ouvTLLeMul2Yk
sNNMGtkGcvzxpzj7QTVn+eSHg5B5sba+LhJuLxq02/5r329tzFZy8dtsa4HltD5DQbMsj44UHU8g
J84rl4f5z2tzAq3mdpwIqfhK2vn+BHZu8UlcbrIJKEkQpY9EPDhgx0vX44IIfHNFCmG2MgNy3yn4
3WNmBdtLjzwOjBTyBBtqdvJWbuTYLVDhGJrWQQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4656)
`protect data_block
L+2JzGz4J7etEj3+YPP2cYj+JEVlESZm7Oa36Rh0m4HkpqOZAT36k/CFwytmNFWGVzvxsN+Ddby3
8vcVEBI8YNAHDqnBGdpmlB7SMSahEHYDm4lOkkjlvjO6cLyxqa4ELSnIKg5sr08Jc5AUhFfru1tb
0O3tpmcCe8tFzMI22qMxC5p93PF/kdSObEUugjNJnI22GCsc6i6qrtaFaj1zKbWLlC7VMZOtk6Bh
R6l7uoP4X8EAQDbmP+/2ywWrVjSKV6kBIIMfpKGDTAGoh7SXIkADH0QWSamMuwx/RYRHVD/R1IfA
iNBQrIUpKJBey4zHeLjfrTzgNusK03dZGXTsizEduuxI86CI7UpEjZVxAOvzEkR31TihUD9H3bo6
eGbgCLuJ59AuqGLIjJ2AqWuzI499EjeZwY8t6Aeg+hmiFdkshMxowk5h83sGyjg7PVA1/AkmUyuw
UyXVYmAkXWh/J3ktEy+48J17hlkG5NfsbiY8mhn7lgjNEFV6w6m/D4YTR1IGdZoXrr2rq34g++WQ
ttNV6ml736DsQvtO59IEANNPw5/DZnlIDZYu6fulE3rmsSnu10UEWIgmkWqO3q8uLv3+Pbjp8BLV
fw4wkVwXdNyk5I3JK08Dou2u3OkHdFknI6SQSipBW8w5IaqIWXbRbLokM1baHLfIkoUy6H0AM7Ep
gqF50aJEu+x66w6jqEYLZ5hUzXtj6QG0fSsDfnQGQ1V1AY/t8eS+VL1dmCSMea8nv1sGun/2LDUc
qg0AIjdCYrgHtqY5UHPFh6tgEZreuiHBi9a/xto4/hggD7pL1pEySCQunoETt9hwG5KUS5fXyS5V
nmb1oqHjkgLg9gtgBVqa9TCSEMVqB2nxAAls8SXCyUd/h3l7bj01Ph0l7F3vM4lDcLVcUIaBLozc
ZIZXGKZCPTBl+b87SH9NcHh9QvQ5dFtEkFF7jzwx5z/YfMkIBMJXZ/WghKJNxCQKY4H8P8TJjFLG
bZ/LJxm1UJ/oPNOURG3EwP3bcFi3h887kWYVjSzeFyTboqGsKBT1YjvbMIKdJBl1UEIqRp5W8prC
kXT3QRMqRtDxcP6ddpI6qc2hWBi2+9/aaCtK8QBALBc7Eg/TXBmT5bVgA5H0aFMQycWkP+Mc4R1l
/hJqIpscRY0tu3GRTFJPqqKMjHMo9ib+C4sVyoktd/nutFls0rPvWa+0+wbBBgIlHD8w0WMauGxk
uZYeHTXTxOZ16kQRyxScWLG9ulAvJTcDQkpiK/Q6ca+UOuGCOkBU2q74+YhPo7Hc8Qg2A2qlWD1U
mxDCy9JJldESWY2V6pfKSj7yfFXxcnG6DyMPBY34wF1FTUI3tBkETvXL26aFxbySCFvGYhO+Cx9/
CY75MJCmMOePSQowgkefGRupyDAZH0UgE30dKuL/l4pof2FJHReFmWdF54kp5ohQwCK88XbWbr7K
F86dEvqSsd40zsAe83YQD2ZOEJfMC8g/NKqma+WiEyIv3faPej4B4cyORd4kxGoyaxVZ/tFB7bKO
3hKSU26tw+77VRlnWyBUJAEcC7bkSK5XXA0/t1OZmnV15kaDHyZVbOdlZpJsSevzDLGesCWuFKki
5fv8k10gWckxhyuasJ26LYi4P9qI8O1qhXy24ygros/a2coPO3Wx+YZd0fW96fucplSCVxLxrh45
g6HP8LaslipduuRB6WytiR8c44rBdhyfndwoZKB32gmKQaLrFM029CaoYSTFUDicbBcX+oPtEH5Y
keHTfSUfFaFgiQ0dSKK+/b+iESlc2WnsuF+6vs/C3YWXIs8XwJcmJ94xItjtMuSmhPjeMuZmAt89
5SAwtHXUFh0Pc9PbJbVQfoIH6+adjPcnAkwsYbxhPZ36cKHw3ygyoV5dzeM5Y5lnGQSudGNKe8K/
oNw8UeC4SSm/nmjRve/YYh15xz3h28b1AgxnBqtj0b8T6Rp9hNvKIgz6z3EFZ9gv3JyI3XFNjgoX
aq8R6dK4lDmwr2zeoM2a+lBOjWsQpU8GxcDD3BE38IsYr/MntZXz0rlVQsaYnXWc/SKfZjWNPD+r
JuQUhjs4UQpE5ur0gvOaIXD31Y8abqlBo982uQWF/2jWtq/ketwLSMCANysxouW9jjjhCnSus1p/
0DlbJs2UOanpSefsqa+sDElSNk968fvmkY9Fa0Vl6B54yH6E9xjnE0QGsX5F0Vn+wePg283aA6qu
SdzjcAcJjufbwZPLbCuRF38/DHQm7IIyYtow1YN6vy9MVOpsX4KUwK1usHc2iKwnE8U8o5iYpJ5G
NOvFXaQ6kogYKHTmJSsi6XW3GKjv2uZAXK9SmyEE5C7RiH2a7w7PgsrUSDDH3kmAgs6KHFwHyzdB
qsDXiTpfnpZgL4+dsvj4nG+ztLfjneShJYuamre9PWU6SfDk82DigoThSIFqlCrwoH1tMccJR/pL
T9xKE7d/L8GlIMeIXyyJ2/fm1qkHKcBAJJFm4VFsE3dnKpAEFa/ce7rq1t7t0N4Oiark+BXHCgOo
V87bxEvQpNETSIVyzf/KYYkwjLpiLb0gvxpiMBpsSdqNS+46nf+P5Z5HPClOyfOBRy6MlKMb2BSa
08P6Ms7Z9NBHrHUwVQvwBYzB/6owfVTh7pHrMSjQU2eAjtqSIKaZ96J9akU52xWi6d2E3fnajn01
hnftk8DdZsmnNFNVEvPpahrCC5tUWm0MlSUMhDyiImMD8lT3sulBIidYdElbkmL3yVCBy3JTAWef
lJSt4wjCcgtefL+WACu2KBKIs9ES0mgIypBD8SoyNZB7j2RAcQc24Pc/F4LFq+zaH/naHoqlR1oi
ClBcvI2UvnENmKfxRbu45j93ZlojHjbBbd+Q5b2Pk3NzhFBWqm4fuKQ3Ah5Wcejc+gOZBn/DeOty
7wPYsAk6Jd0vsxGHRvFM6vTNHLKDpDs63+0177+svjpo999u/CbAKl03UI4QP0QZEm9srfiPYNiB
PyquutBPqLHjc6t7SXWZvUgUmMEu9OY1kA/HFMc77yb/8xKTV/YLyq9LJrMefzrhkawldZYPOLeq
rHLFnJ2SYGwn6VzfjriewdcFQtob0dnSwLZMHyqZRKCm6A7vcHPYizd6sdBmswto2vf59OuFNFbU
rjC0CMz3PMizwDxu+ziNqptptNf3YiTs7KV9nzernD6A+wDfeY3OODUwQkKIzfCnu/bMvHejJRnu
YIE0sViza1s5gL7gMmHwzAi4O9FpG9e9dJuYD1vA6NIjtlbiPZiiu3yXtFIzCXfRZYRw4wQRwcq2
9fWYNWiW1Rwa+xMy/NLpX3ez/ZU+7wFT2jzDOSpdvC+sYlHZbCQH0613vlqlZckJanP3EGDYiwkh
1NujUjuMD4VS53ybAITV7XQFGwb9WknnpDH7S8Qs3vZ3vofQn26oD5DQVBVIjT8330Z3RYtSX777
Kndnw55SkDyw34PE2xXVvCKUhpAoeksVhoDh1+qWCIknCBhCCgEvyQALHkyV/50H5tlfL1w28/u4
BAbdUwbO4hiEans1QCRYHm34RrrwBSSIAkIcpBhfBTZYI68tZ6pIDwGsfvFlhoFRJhzAhEXt+5ag
qD0C7e6yqZTP79XZaPoPtRqpns9oeXXPMogLYVGXkWabmUx0b4UHLum99R/WVAMNNGJpVgkBhlY2
Qela4QlAVklGU4fAGAF4rubLYHcbCwkQDhviT60bpTtIXEyHhkuNbwwD75S5cpGaK3xY4DQLUI0X
qZnE3Gde3getaEyAJkZDIkNDe2D2AFNHd92kxktBlF9drv/0wTP2NB469alBgp8/5GMr0vfqC+MI
4vgxoEMvqBjuIN1CWNo/wAvh04Fiuvo+qlq81Qu0sWNI4T+6on1n1NJxA5duvdgPUue7VUnfOr14
jsw0gYX1NTZ9aRBw9yuqcvbNt0UrMltR1/6lZoREN1SRY1cX8UvbU3B1YPkfauOHU2uOzLOUQ5dh
alC4i7XZHp14p4YwlBWK+R08FYkymKInuTipE9Xl+FXO/5Sq15XQxeK7CQ/tvQyR7kCNGqgpX5+P
+VTC/t/zJQ6eavnCrM/v4V89of0W0L4jD8OxFQPwWGPg/PJiOsLYk9KgUoMf26ZwLXdmYWGhO6v3
uPcRuoprOvYSOynFitwQ8pXPzVZgfgt+Cg6hRiezrd3ABIhLmDwo9/fd+Jgmjk6IdkuMgjDwns23
dKmdYWbbMAz6RFb+iARq0SPM+mnbL2MmIJYvNJ0pl5MLqyRFAWlYEYwc4JDEO3BDjSSqGzhX/Zbh
LUlGJl/Sq5BCJ9pPY/o44LgyykK87GJ+l2dFzz9oA1xPoI3gvMIs8RPAhA6d+HcD0eTs5NphqWFN
WiS39+hjwgllQlP305mWpSCPdlZOH7DGUQXQi2c5AWabOPF32ReHYE/ldH/hGbipoODY8Pdw7Qh8
JFHP42qKebBW8A/k7ou8gYF9gzVITFcvg8BZd5vTvuPQ77tYTFjk3j0hXGlVLgzuqTKvI1i2u6TO
+N128JsE6hQYe8uzkb8uUKffoj+e+q47amzcF1GpXIeKt+5/v7ZZtFrrUCSI/5PKLUI8/bs/u2eY
CqP3jROaXFSULpMxXtWTwz3iio0KdltkQEx/zRqPHckl6toQBxE1J1dr3c5cK9FN4OnabTsCFjO+
HplMl8wee8CVZ479HyCKw6DDnd3Z3k+U6HXr5fKIHGOUb64e4KUg8Zo83KarvSafjCpWnDtdy1kI
4sRhQluhJ69zflJTWb3XNw4NPxXCCQ8XRUbHoH8lMix1ci6qsTmNeGY/zpa0mE2fhavh0TmG4yJX
zV0ih5KvhLPnP5qhGOcxBNzsLxJVzw175Q890X+k3SgE3mXkqyHibkIwNMR83W7LUX4XXCW1JAcW
z3K9VkCnS6r2Ufdebwyw+x12BkQu9xamMN2Mdr70GUvm/c+73tliYWk+u13Tam6ktbUcgZIb0aPK
5MrD8hk3aDGvE93B+8RJKGaGkWK/eDs98dmLGQnxn9RrA/4tNdQVl95bDZgcfD4H3iLIEHRSLxW9
N11w7cFHWYPasTTDBwKBHGxLQRE/ih7E0QhlfNqs8SrLdZO1GUUhrCtMUyEkY4eRVyqmKg/peg4O
xxsKwHAMMVR4XdKCwKjzRoQpSX2nmiVszIKcPNnb9iajTBVP7uaP0UvQYVuiIuY87EiUmlzWil1e
0lZqDz1zinCF7+0KPLMfFR3Xau4MyYbaxQ8WCWRbzcgYIsoTIimmEHmHawMOElbsMkKfeIswBBmO
AfUQQU00M/a6odXpcACmcz7dfkj1+V0FA5cdg3VEk+1ZQcao5rFZYKyN/WNzzJCrTvEi4hsePKl/
TZUf6ccvDJBQG7GELlavnZkzSplU7nytluF4INouObp3AQfbYCvwbDJG2Xoy01mMz7BmFDXbErH0
4/Qp5pdo+Af/V+sDyDXipfSwdgwtPNPLVP9p/7X3R10/jukXwgE6ONL4wVC56PNqJDG5ZsX1dnT+
jp921tyIU1th5UJULOObIaeBFGYW5NP4s48K/z98R+Wcvnv42tm8sjEbqJJuWG8WGj5N1UbpS3NZ
FP9z33gz9CA+x1KpDqz2wY+pSf+BKZ+LzUqdCoZL7QMG3Ifcs9sDsHVR+ABrrx9KwU7iywzYnbHq
LOqcMzx10/1DqmTW/lMH0+LAv+nwTASqrMloSSIlKyfECvAfuQMyCUA10qFUEtwvL1Qz+SXm5RlI
1yYQ1SrITbB+JNfvl4x8NslEgcAOjx5WXII1A1whABnxPeKIuOcNOMNi0z+TX8WjqmFHqodumJDV
tirrp42cl7mk1imkPlqswbLC9/F2JzZ2+el4yEC3IChInwwzp62QdMpPsqXlBBDKEoQdSEtR+++5
Kgpx4DcJl+lcnUXQsnUYpUpYnBWNdy8YTJmeI6z/D2jbkMAr7W5LsMd+AceVY6WM0NMpb9MJGom4
DC5J59QXjmk9G6/wAWPpCz4+H6iZ2twEeRYVtAoaSVajw0VxNI33u2u9aLrCrpR/bxfKKDTvo1HC
54QbOnDR7RMoOHBVykjS7k87af4AWX7opzYW59rAS/3GUGsMKrKk+QvJRTrjx0YLzWHrC6YH9HzE
rEDFdpOre0NICqVuhPL3/4AgTeIezS5Rfo7SdXcPpubqscUpTfpVswANjJ5rsPReCwx1AeRINTIL
Q4ldr1HH5PKHqjLoINKQrzxDQ4tcJY35ZSjLa33TU5u/xpiiw9ZU
`protect end_protected

