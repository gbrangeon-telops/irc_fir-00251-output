

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rLWvNa4xmaUmUmTsHaZZpmf+vdo1ZTZAwtQ7nnw7ufjv5GWZXhLdNQy5Q06lrQkoXFZkjYTdRiP3
F6m6R2KGJg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hpohmRSyxraB2TfGOSuLyUSGGabJEMublC4fhU+HZ7LC068YGUgk2aE7EHkl1WtDE9Bb6v5v3Qg9
2I0FD8nMKFfSIsem6wrqx6FPpal5aJB28sq90dkao5/Iru4xYelKhv5oyEvq5w9fsErMuciA6N4Y
mVn0CtqFHil9PLQizOk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e2qQeTSxab1fevbjz90nhYXx0vSvMvWBAXsx6NPtcQGmGbeJ/S+FZG17TXPSmNs8pJl+7MKHcPRl
s4fPkRF2q+UUqzkqGrUfIOlc9iDcSV3G1jvuqC/KwL75+As0dV2zHDw3g6spyRgrF/QyMSev2EDX
wNjTOD0D7tDHqk1b7PsRTM/m5LabqbFbAoaZk3OIm0Vx4hjx1H+Kj+5LKlzym1OWRKYofd9Pxrcb
EMUCk84oHB+E99UNC1xkjUMB3ggxmGGz+tj2pQbz0ixGcWE5awa9i3czC6zJ21Sph72Xl+p+aRC5
JcGtcY8i/+JbJchaWispPX8x4NW4FjK9r8JxKw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vltTKSM8a/zRJ1QJ/9B9ijVL2/YbgBrtsRTG74WarkSfaW1TYFA90LAMjfijw4Dh6V3t9bzMVLiX
18WW94nb3vnRj+WAyEjiDaLRKxJmoyxgwsVe3baoS8c9YLsCvI4C+2FRQmKh6kD8j1o6xfJUhYAE
QHwYAw6Gh1Fc1rWYuMM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jeozeC2hZr+0l/LK5n/W7u82KI9P5tCxn4L5QInLhVBS1ZXkJv19EUcHMrHeYhgivoQ0MQ86TEXP
Iah9T/vQMV+h0mk/ZiG6XOYby7qUUR5Ipu6A3NdkCDCZw1M+w2At4X13RPUlLeERzh2uCLeznee9
UbtfGUHB0e0CGrBNEj1LzA1bbcGeOcLXMz/DrWLUmi+Iv7nTaL15UXhNNoh+XY7m46jwFf+dQiLA
SkppMG/4vt/EhyL+TyDlc4FcuyPEIIJCq1gQ6KO1U+4QL61Qp9FOEA7sAw8XZEnuD8uyPmi6wlXt
gqJWUq4qR9zExL8yZmy88nYYAn2YB3+3OVd4ug==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 123472)
`protect data_block
b6OUu8e0RU/76XqU3Ct2Dz9ydMuNkvGk2bUIOyjZdtMd73LHDaEJaVlNfkEO4ANBq0Ri4mBnKCmf
aVf9D0F4uocDTxJjsCUutJFkaYfJS9Y8en403AWSqcl0aKLDjI+/GBuCDc/CKGIZ9odT5Ta6Jm9f
B4EVn63zFp++FLxktj1SCzoFqAULUsXOuKrUZjaym0q5T/yE7K2SILnzXbmpQjG9rxEC5wdxUsIJ
+C5nQgZgiRjzhoYN/SePifoyu08V3YjMACfeoU2LvRVZvTV3IJpXZq+8aaYFwrcvsAb7/YA6iBig
Ngi3y30uNvjUVCkpnCYQJjZE9vmgCclVHSji8uEhppXn/FgdxeY+qX68YnmLmli/xUEf6M6TjuBR
uDvsAeYWEbLugwiOQ11PX776QhCoSvadkcTD20nAedDaJPMAbM6ECtKNR6rEAeR4WuFZ2kCIUOiV
dwWLQJ9rTbQviRIR7W+Gab+yqwFwPPlcIUJvSaXSnDd/bz0rPjuAtN2uZ/ijs3FTDdYDRj2jfROF
66FT6BP7fxhYlkMoqAlHq2FZIhAlGdWRg7MtO/yrWeDDvg5e1+GsaEYs1SCYMyWum6EAU3ZvCppX
0UiGUy9cNo/SZbHA5t7ZkORY/8shm73k2fTdrZJIc+sxi7l5AiovOUvAYIXchTLI/3ZZpJbhpVVj
LSuPUyBb4tJw3WY8/3iYiDEewabQez43yd9OxqrWAgs+PWJzUXQSH6le9bk1nXZIVIprvlbP+UxP
ISpb2oJOnmVoKjBKgTzPPKnnOowYTkf4UKM1twTNeDkqQ6vP0oJNH3+IhZnNOYFjCFI+goPW1W17
w/QUyOo4OO1frLSQ/X2p2ZUWytGSm6HrVYifCreihww5A5LU2eV4GPxtrUcQ+4G+MeLcHzpI7ePY
nE0inmdNYH8sDQNvp0tCJP+sqm5OHEwH+zitBsjljeHDYPz0Uy1N/s0oeDN+lwSiCri6jhMNgrX6
MCLt0LCB0ucOVZuNL/Z2ANniCgcnrNfbvtpHqazSEOmbIFG/S19PVRKNF2AmPk9LJWCWFA7PmEDM
DQyVQMsJmZ5HnssZTe03wP7/02RTL5BW/KpLgV6XSSBtpssRJhvqi6M2sZHDC1wcAM98+UBGDDy/
qrVjGv6WtRmzHUVv8G4lpaXxo+fkSNuN0c8Zg1Wj2tdqSzzLKkZIzgh+XbrMJAxRr4dpLfEsb1+1
+Ak6i0HAzQkk1i3dOE1L1AS1MgLLG+DMr+M7KKer0HgefI8SBScEDapYoYk5UP4S6KKbxZNXO8DR
djHpaCUo+DIK9YcDpz2AmKbXa3HzENK9RWWJouXppV9KUyOj71zdbS/DccVqz2n5V191OmayRDtt
TWOv05CfvWbq2U4TwBidk4p5XevtOuB5ovu2zU9OoQJe8QOzy+bJpCyo1gwOtFXkw/Z1r3Oo3WzB
fNxKjULfHnXHieBde+eiJORy90kKPHpAKLpoztAMO6H9Bh29LBjdg8xb+m6igJZugapM7Wz+XEU2
A9ApeYARWIBEKeFU/1PJKoqgdZ3nGCFY/qdssrcpYag/npHnS0ykrcFQONfO9eEFggmdqHuZue/R
iPJ1MF16gAlrobaNBwgNJr9E0IjBqzEvuMdnNWv5fNvCTKfeUKXFq1flXNp5iW8XhL1QT7ABJynB
kTzM/EC2o/BdBrk2Hwu6qkUpU87bYH6LFWtOvcY8+quN2n6JtV7dU6WJw0Emq19lDkaCc+yolZxj
IQZY0+Aa7jdQvKia/Cy35Pd8rvHfhYF7XmB9+EYqCjVZbzjZxUAxibEGGS//NEXAlBk2A8QvCA/A
R1fBqi/Xw1H6JJfgdoNCrmG+awRLh1E395ymylI4+irOptL5yL7NQAy4jcEFW1GQTgMG0aNx4Man
P6zSGzGFiA8utuBFGckr4gdGnOMYp3TD0iSXfPl059Thlh+8Aa+axHgyhAo/mJIzW43rS+f5BVQa
mkaTjVOkONkMXzr1SLNUE5Pz3c1Dvo3qO5Abj8jUlxnm+GCd7Tx8FBpVbGFEDG5yqTHy/PvnubmE
mZHYNDrXBHcd9KpEuQL0YbYC7p7PCAB/OtVwKXYUYk90KddI13gTi2rx0xI7GKhvqCbTf71mcNE8
cP9rcat8VEpNtAS0g9hhgg5VfYY3wnVH+qIRi2eOu3JKMkecXx6UuIlsQIi8n5/Z22Jemzx/Hv7c
OSZX7cuYCnugzhGzN+0xX5Sh7esICbwS7hMy70efL9+i7YogHBvKtOZbHX0yOvEqEBNtUk6Kkxdm
MWsqgMPjen0XrC8pqdYGHQXH9hEqcb7bRxgndWVrYqKlc6lFbLJYOEx+vH9JYWERVEHZsjrJg08a
NodhRA3IGapSPplQHXKWZHudUAO5ShfywreMgYLo+6MM0A/oz8NQQH5jGzf/5Jx9Y7z8gOdgxci0
SMfpcKLYRebPx/REjsjGRkpFBCYRrqclVwZn0I9J9PKJZDpXSzw0XVQsNrQzjsvkK5bKZY8Zxo3T
tqAMr7fW1h2POINQAWiupnpz1DCcUWrTAi4YJ6c1qFR/wCdHJY4DejC1xhwI0sjrYV8xDoubhe15
zezfRhv8B8qaELJrbKgPg1mi23F8HxATgfaQplb0Ov9GulOWwT/FOwZYk6pXlfLLfzLl5u6J2DF8
9jXKiSqfyT61stUAUKH+T7w/NJ0z/hCIxt+GM5Q94DKkgyfUMSpxJfT4smSj9MkCh6I3JOxe2lQm
tugaMIXUU8WNOCyzNYqvC/Rllh/fNJ9P97xYznpgbNx1HB82BI6MlGFT9WXPrdJS1m22dZDsQHwb
YXZJdYSUsNYvZBbpe4QutoZQfsPgJyt/2u0zB2rBsemB1o1s44CmOTWGe0Kwaxb/HVdZWamtmZ34
GRnkLDkNHuFNgqSZlDtQ2sRPk0yBsyd20z0u4ayAAB25Oxd7iYcCC0vPoggqDWToVlasTsTGRRLM
oj3EWXWMirLmQbD9ppDzWVgxam5a4PZv7PQo2/YtVj8oAHKaqxLaGYeRc/9XHO4/Nzcs0lNV91G8
FAKnkJ/KreRHspuzbpC1S/geMxmzjr7sTlZivZsGltBOjjKyOgIUlmwsvAfM0cyJXe+OHEVUOOir
oGvrWDnvv1C5+wnbCNvqJjanehiXw7l0sc8kF45AaqlQpliesA/AUdgKFIp7+9PMhyfCMuwPwEp/
UdhKmB5GLjBJW3/Kuxx3e+r8flcSp1GTJoefUQqUu6X51aJZL9/8Cgmm6Ud4ZjXWUc1onLWKz3MW
MXoac7Yrz6tF5kKqG5+8LOE2D3nzDzBR9W0jxi0ALlP3qHdaHCX9S+vk26eV72sHw8MeEc/1WuUC
PQ2x6MxLM8G/SNBVkex++/CwQ8/Az8t+sudIauHzsle3+tVwibCa/qpeA9+9wT41+Du9cBM+WoFP
t121lCeJV/EgfRj4z72HQWyDnnrVLUB2IWHVQicu3l5q15jzFdnw/YrZ9k0dwFJOe+haJyYy0MRB
4XLnoZs2IlD37iymGfOkYpRS1ppYXiuoDyUF5iHGIrCQ3a73fhTBbFJb5d2Xw5uYMKEbiVhAG9of
w9kGGGeq7VhLGPehvlu8yN9qCoEfm8h1LGK/aYa8/90kqdnMuO92rs1RYaC/GbQScp68uP+1A2Tg
lCeOa1oxfyD7lI4C62ReiUVmKS0XbX49YcDjqPeGfJzf7lNWSCYylKcxMg0CZVjpkhEyGdrwt5qs
thnVhXvIiITvg3ARyfYBFFjgC+uIucL0fe4UcT6UGjoVycAi2E45i6of6kHTAg7B1GIvoEtQpOEa
T03YOinmz5EKBKTVgIl8fKKtUNFWyt67QFTlD3+lqylAcgirXdGLYJ439NEoFjprgbRva3FEhmMV
MgmtVV9Kb/lPrP2VV6UIJg+vORfyNNrAf2aJTm+WDJaXI/N0zZoczqzkvhHSBv2MW8BdMCLWQbth
Gw8+c4R0YPQuHfNflRuxx+E817hjZf2RPIRUhAktwhGAx/ZjYARKZxCMHoUYlaG+itvcUxSE1rWZ
hJULXgbq+vvB1qhzEfEmawz+DptjHNB4+JM4NbT2e4WEWlmTh18eM6N1lPh5Vl8xNto5SdoPqVs2
YbpDENfYGgRKeWUyxtdya1+1n9g+V5/qkMO0JO2p8K9N9AQyMiT9WF6WjMABxHkQO+ycs87yG7/b
qK+hOeExsvKJiVVjyX3A/4cvDO89yDT29lIAZrtX8eVH56j1PB3q/9RbvFmb7B4lMzmBNUatBDkq
unltT8KhDhcyjMinHbuIIuWQ9tk8o26Ch0KKYoark1gLM6i/mqAlE1dBrj0pF4QAHyTuyaDqkYxE
Pb5xmwJ+5pKfj7gfVl+wZXabFrRNtSw3ijqRXwip6oGvqpKZt1iR666DhvR5yXle2BX21oNIGe7G
nGRAONiDUYAeEWW5VWYkARmDN2ZcJ6egmpzt/jeqwdxxdEf6IGgJTkcR3x5xhCaN4cJKPk/ZScQL
aFg0eM81ZR7Ly3nb7gvyjj5inFQbeS8Tipn44qTUvILitfyP/k3UiwtchFgpNWJ3Hy7ui36nYTdF
I1Wbq7BA5phuCWTRmy/tSca5hgchQ9sJ0kmqK+Nm1y8CVemTaKGmxcguQBLY1gULaMR1MWzK39T+
b10opVl9GX61rkJRAxId/fUchOMjIxH9by9471krTrjdwzcV8os5PXUVpAj7YoLgzar4uv6FMlYB
1ITLRdcrmcIhgJKybMuL1yIbWkHwxcPv03cU46DMH5xScN76Un5zUbegvj11o7gN5rz3wn9J6nc4
JpfKr5mA0MUfBuIVfywSlwKJFCtbkIUF3MOhKaDhq5dpnMd+POCpxXdC+o1RW1bNgjkO/XO+hOQk
G7LhHIXthVvf1z0lVoS2GwF0/yor53X9loqMPrzjEkcjInUoAPYCgzLpQFDK7GkHQK2Nma5t2r6o
PDDj6hKv7ISEzVP5UFrMA6B2BJujoAsc+ZOdNwNGhdFDaQ3Tj7qTd3Lo48gK1lnX/xy2VSArAwGm
P3YDa6XQtsqsju/HG/BtXhVV7W7veB09VWPovUUdOpmTyRBXGols6J4aAKcQ42+Lqg7BKaCI1IJe
4vxrotkAWnPijhzN2TsFvCY4zCNJRV05VK4V4AALYTBcjiDijqyLcjNsRNsqla+WdS4NaC0c63Sl
fPh9e6n6X4cd8VBfcxxq0mJfihayUMFx1K4lKHBvV8GY1lEhLihdGox2QtSLWDypE5sKoNx09rlx
JW8ZISGlzP/DUsiTJPEAl9k30ac1tCQ2GD+IJTwLrxKZ1USi1zRj1k6VxJ61E9W0Kii2TDmiGjds
9OnzEyHO489Ivecuky5TRPpbbwaxFPA9aXZmyk5b/pZ+EVVDDdXsSQ6Cji4SGh0BIOZaqQMwcgoj
3BW5/V/9ia/hXEJrd4EbNw6pgjje8ujRuPT6SQfw/X3fPFp2i4hs+rxY2ZWl7/lvmFhaK+1mQ4KQ
XCDqK/2KLno8Qqcy4BSdExqDn397Kq8JbG1Cj/CUkH6Fd5JTYatGV8cEZFznnvL94mtP4la07BFP
XJgcKg+2Cm8ekl6QY5qf8AsXNrv8CFevo9S0ZYi1YnX0cGelsw1KNSVm0QbSJEQ1/aQC40gJzPQL
WWSn3ZVzhVbVrvGLhRMt0h/vVAYywxAQifiXlZN0Z5LiOJH1cbxuwuqtZuYfSX1+fww7//+mIG0P
4OYMHSRQ4/A6ZECIREeGMHuhaCk7fCGDnDZfWYfaCTufWtVmMHK2SbRTlaGfgQkEBzskpjWeb2yX
Yeoa2Q87Aq6h+tmsZMgbWZaoXVTXEtB7KdmxcZnGsc2Bk5FbhX1smW55T9lSydBBKsJ+41MStGFr
QeX4P+wKzKs/5cHzn7Oux5koHMfEIM7YGQLLAHCZ/NOrR6kP6P2B+drbrWX3K2jcQMEt2DHm2qPr
eL6G2mbUvBquwl/b2RsWfsAjJ2yXqY1zAJSOcXOqw1b0jy256qbJqnmjwtoEtVUWvZihghTfNR8r
ctlz3kBuG3xJ3XxyQYOusclBjfYWNgMLc+GFvm0NL3LCnVru68F1LlD69C4D+Ca2r6yMljdALV8T
BhQ1gBgykYRTr+il6TE5omcT5C7NBw2NYsTj2P7yIS9wThnMe4EDS66QrTru5lgTGUt7g5e02KUj
Mfmm+Iw1VhfNUwTqIMaX56uGF0Gttgu8QFy/BTWWjxPNtOPKJfeoWmRyZHDktm137FcuYFj3TD7I
mmajrN6yivL8MV3Y+QRLK3+AWZDeqQFA6DggDlnzKMwZ/wM2d4TeuutIsXR/8EWcRbNM4sXVBvbN
to/IxUFvM3M2jncNnNVkPljBd7IaL2mtyu9m7kGM4DTdV+gB6JHl8iZemHiIjnHyt3B7ezXUvkWf
wdHLQd7CPWeBdGcEWnkeLN80dH3Quw5nYON/l3wnhzRWqhMLjyBBNR6muB/hAC/LieAhtTsUlZCC
3W4tNnugVKu0xmNRKHiAteEg9BHK0PL31Spe5ceBELW0AFk0ZFzhTVVbktKkjU3IJ5TYoKFcVLYP
Nql+tWwbuvGVETnWIIOE6szSyePjTZ51PR21cUcB4EfYlyQRUiSFXRaRFSTR9IVSJX+e0YCAx6Fk
fPbXkEpnz9QYwgRtYI4xHmLnK172x8gHTTVsAxVOBa2Qzi8EHfbhkR1vgjYkRhvsxeM0wmpykIFz
6iFawt23YBs5SUDPdTD8qzswghntOt9ZFIYvQa3FvhqLakbLP6mABNhCzlSc7UUcg3bQ9WjXvygp
uQvIMwx2aQMaT4yQe+8k89Pg/nzWZTazsohJGZ/QHXUtBZB5mGAYGoNiDLhZPUeG/niV0KQtvhfL
PI6eWxmpFeTgU66b3qN57ChcAFqZF9MIIywOC4CF/1uFSL/TH5t46t6dfeX14ZcVKvvnjeZ7c+RH
n2l7omoNrx6VtsvK0oDIOQiEGiUuP3zXkcF+4cNbg7OdQbMmWv6DdqfRwQuzVwj0mLFhvvCacDVh
Mrzxk0lwqRJLBGJQ8qmRFCr+ii1iOlO3f9oprBoWtV9IWuY8WRPP8M/O4xJWlCLfi6ci3aOJ5stf
BT9BXP5YOnGYbl+hf6VLFPI8Qr5iIRAUsjqKJDH84O3s1OmPMnWhivuztFsLrtb9sLwBFvHm9pGe
QKqB3cmtgSreKi63ntxjWhuQx7a5w4YYik4l4nv3xGBtaJpIdPMCGl3glf00BBiq4tKoHlXFBYjg
grhc97oXR+kfe+KH4ZtoMKJ9wVXElHJViY4Igw0y43HN5yhXmfs1eFJLFyvfy9QSWemdv1Q+Rxhx
PsCaiGZ3r281ZkfLaqmSPdHfSNa0zMmpnjyZ5nxC3BZ2VQMu7vPjSo7Vd15r/vU0s6qlCf1cM06+
a2URsktXWk2NJYBLY7b/Itd8sT2XRa/0c9r1Swz15NJXDojVJaXL1JDCAc/1y41wuArfyI+pAeMF
RndzLBVlC6c+0THDdziK4E0DQ4oVVfcZgf/3mSpD0L46d9fukaaoGOryNdKHJj9PLkHRET2nfcmp
v74ameFbh6tur0+fY7G6+MQUeyEebMOYeOBZD7zMD5eoHL9p6cPCSBTH/SZvi8mfse7DvqSvYoHK
YAC+FvrLixft47P1M/voi07Ls7K4Ea9QazobK8chW6N6X/xxaVDDOEcpFhwtKHKBMuV45e/EnmoO
vGspKzXe/0uREJ8GMi3Qfo5dkwXw0YD/nGnX7lTDmzkJHhAilUpKHEl1UVdQcrvSXtP/UTQt1MWr
ns0qckCZCFZU8gnAkjNPPIhV/f0dVF/0dFPyywyWkRDclxBoeVbQVdVpQBUcqrstMAUf0WRZq7JY
YS4CDovU4YT4n9tZn56RhkJzN15Ga59HLeOvYudEGwKnCTnaBbsA+TM874/UyheLQiBwZTnmFcD6
pohgsvy/TiLj50sok5oF0CbUogsiwDr75IYk8g7Afqt3vo5eSytVtMxbXYCfN8sfLOmKPO2niGvK
1ljiR2bnMLWsuPpBqeLuFNk9ObsBquHPHmjho79JyDtGbPRFXQYnr4ntHRh9Sz1sPLv9ib9IW8hn
v3da355654E4fFzIStVB0SIizBjx9l+kVXmqab6J46ahkpykWOxT2MV5XTe5eP5uaDB1oLLy85pO
3gz339WExSLF3EhlFo2G3+eDAkIdutmJx2TrSC11ZunjZqf7s5SdPN5lcV+tHVT6to/DcZcQmOyb
u4M73QnkwuGIzOXd3D0bwspmQyKusL1owbOAh/WGZOrJ929ih1ayQesZRhEGSW/hagyuttAcqhIZ
pW4uTcxNrhu33BhSgNNd9eIivtJhDBJeneqcWIEWiZn+w0+XO7ciM2kAz9ydyQ3OEObq0/aXH3NL
zMHxkJS/EPvLZl8AliNV489sOIaL+ptXcCw97m7qZt1SnNFtKdcZWdRUzd2gzAkL/HMmAG4hgzoh
ARH4qxVplxfA3QVMBl4QH8/hmkuCoKHNLmQkK008ksxauN9Oq6z7R5bkI5fzMFPOHXJXeJsHAsSB
z2CSiCqR9Pg7KFzIoFEYU/0vVXUcJxWXRR1DsE0dh+B1atZA+1P+8GOsO1KOMGGWR9TcoZhQaJTx
ooJ1FaNngUbT+PL4QqL4apKWRga7uF+jDmNJ3lPyCkcesClxDTLlsFWylk9T7mErDOG9sdozkgm7
eMviVy2Y+x9LW/+GedvujAWo5+5kB15RgV13lKX35NAeUHZ+jW1oF9ngNhlgepHgi+q+f4MIzxno
AYuvzX4iQNRQXHp2h7V/48sM4rUr36ITZitWyT4mzuwuHT5IfiqH4zT6sHGAt8yDk4ILsKzlnyk5
CohGlDseEBANjnu8KBzl09w6yXp+x5wytgwi2onJeATFekI3rsGtOPxFWaZ6BuVykJ1RE2OQCtlO
TNKSNiBihwfU02Dw4XCMAQTYiYdOPFdWy1Fuw/TYHZgk2o2DEWzBq2oWPNBSPhl+CiPnhLH8FnCj
4RmJD/P85TQ0pyeoK6Mim0v9L8x0W752/0nGrcCpJHSmVFdhuLXMiBvhE9XaK5ECjhpwmx0HNIL6
q2kq/OoLFumn5ZVYggnzVmUAxWWz1fxVjBDLqGFSSObasRoMSBAGxm6NQcbyh/p5ncpUQol8xUgA
c+MTDlF2txYYRGz2f+bTMlSBUG+9rgIoPFNfybjwS6GUFeGKY1D9J7IeuUnp8vhrzUGi1zDfDBY+
DT7P1NZS/emNG6lImjaB1AmhsFnG3JDetNexsv/Zp47ThX8qvp5FnkWDzLx3/JJpKz/yZ9fpi31u
0B58QSk3FFpGZAX6aIg+RUextzsYpPO1c1aH9q5RKh0SjTCTvyVUol7aRzg9W4CofhljbL9HFWnW
JF9ll9wVME5VQ7oYIYybTh17gonAKioqNZkt0JkCIUMAJOHkM0pTFOp/UlHJYnZf4XAKev01O6m3
xdc8L/pmnlTsg3KhiJ0UTfjaYzooIdeBBnoNWSpoFMSNAFBMbhVMCtYrq9WEKayA35t1RXWQh1wb
HycBJyDCmwh+/QOp1LBlJ0QlqX0r3rU1p+9VoC1LJzdf+LM/v14WEbAqP+oco+tV97igOdEHfHMq
9KGIHwDddg0CSvINjCGtdExP8f7eyNcT+KeWDr8a0JxMzeVgkgwrYYRI/VCmnbpfbpMnYmsq2cZy
xd6AMEyW3J9++ic/Z7AE0p8b45fAg31nAMkPUg+uvTcL09i2HqYBqyTQDrS24Cwr4Z1YdB7sEeg5
5ocaT8sJStJLoaB9/FXu6+D34MKsd17IBWAHamvyh6TiHzfbwfDbvkFyQtEr36ZP/utWwVtwmQAF
4HV7E4FnfbTvlyp3/cSiJaiazFEwI6sFi7xDQGFPc3MnPUsS1DJFa3FmT1WgAfAzIgei4wXJiKej
VvS229MczOHBRIvI+r8eQfdmHEP1SrqkX/u/tJwd5wgj1o7VRpMobyACKN65P5P+fmOJo/REH1uC
qqcoFojAlkt+5X+TlafpNRObbeLUnPwg+E3mLAqWAXpDbbl9ZRrLp52mofZBboj58KujZlpK78Ha
+V9uE3Q6Q3xLaG6jQWTUhnebEp6L5TzSNxkttxcvRTa3KQr3qVO1q8w/O5hP4qREclIsqB/NDDtv
nTzYA2nS43FdNScZqPoobKMhP5evOXT1/fIuWBSXOQIoCI7jI/uMR0jji0fwZnQ/LFtmayAIzOxQ
E6f81u9kzJlLLhGYhiWiMnQ8GBGxgOCAVCITthOaViZvYFARyPvkaY1oOGiqlLzZTRt09dxaRvE6
tD8VcRqfrVWAJWUtw/Y2WsWQsRTK0NLzpnrK/yschIsNMlVpWgshV81VFHyKN0slh22Pee0iossg
Tt9Qclu+dsi0o5GKFKlhDwdF1hdX6o8ecaW9tXoGOsCvP0Zo2FZ8ffuvf/PXENqZKHPPmD5c585J
mnmlFZGOohFpd2bhzBpF7LJeBBbyScI0styMs8LWW+eW6dDYVooy8xFzJCr8bPqBxDzxkII5R6By
VGEZ6kKYoTSgs1bCWeVPC/QfJtUSt7uAUW1yhvEZ4LG1WhtUbtDd1OYma39+ctGUIh0Wybzn6htV
yFKEfMarouPmVQXYCBXLAjeSHqTaOJqQCqBZJcanlwPiHWQwC69vwSaB+ERT9cwFvi+DMw3CjmUO
XOFx6S436ynCC0GUd1lraQ8xLFKg3TklqghvLLEY20/p/92jof+yQvTW2D5UpOoOtkTNrugpod4X
Evr1fC8uxTc8mRkDZmfZ51P2Xdn+OrMfuZsgvayWOyjj+Iup5hkyHTbUQvBwXDS4lTgSJuApQEp9
3tRhotmEzWloGijHRpGhrLRhK5YIcXm0wFNNuqoVHUjOLgeza8CpPR6Zj9bFtepArEFDkOCbh/8n
DQbEWxB7nBjP/ISKnTRA+bQ5jbSxKkFoelNTrBqWthgo31X7sRPaB8WFEZG9YiIsh17S+7BQuwpY
T2T6nu33aMGPyM7ShmcMOyl2BQdwW8pXnSVGBcGsXAkqiVbmb3872rAOFwIlEVPhKv6XqjwzT51b
5ePiVX0mDniFm0+p2gCV9e23fiKIpPuD+Age4t4u6Phc71uv72Uj9OUWMIvQeyMF3WIA157sjPLZ
elb/E1UX/7Lag7wMIA+k+2DNqOyqgzzCfgy4D/g2/8mSTVcOrpMUvBiOjcvwlA42fZMZSXRx58J2
IYttxcGWIA1QY0Vu7JIl4QLlFWCXtCKL1RZ2um0BpOwQsvlmYgAE89EHGQtGg/MeQPLLDwjn0Ist
LBvgTQSYnfyTLhF2H7dSF8EA+kUOV+bG065sTIGCD3N7hGP3vosiiKGdfPKRB4lh/CJu7Jv4afMO
D2ug1oXtytlz5awY80c+WRYvDO6k8OYh+xShcpqIS/zuqK8m0CL1h0ZLevl3S0MYXQtphADaEjNr
3c51E821qTX8GRMD6wfrgb3z5NNOVKwNLw03jT3Q7Rm8l54LguDiTYFF6tA9iUtWuVyMUiDKn9TE
2BR4ZLZlrrtAVFG92L1tXnVdXbr10+/og4PJjY0zpqQaNX8qQMdasQNSao93+vCu7LwE8UOUejbE
wSf16mOVmce/q7TMsS4AFsO4XWxqWKtD4W5KTn+wW18YLSqfPN5r5LmgJfm2pfCZ+jB6HcULr5Oo
AxOW6DDAkjCwoS3yFhalOHeqOmRXorTD0+zo5exilO+gOgF+KekYVPw6Q/Q5Q3Ia4Xp6mURea0ZX
o/OBx2gHZI8Z8UcnIaThXExSzWpZRoFLtCkN8qKZUNoqLf0rd/zhkUcUD5iDIaPZlFwfhDP6ADaD
t0qO+ujzuGLLs9habgqYKu2S99Gr4vA1rDnjKfOAu26y2CdSSapjutjjqze7kdMMAsyLNlQeZx2X
qJn0lbF6L/MDA4Gvx2WgF8vG/bzgGpFe4A5X+e8THoBobyCNkDcWIWGTSLraXe+2yfRK0ZOzg1Er
zcAGzC4KhMKZmFS4R2vBqrE/IwEfledd0/J8D5RkG4gIPRe9YCivLiCkEjUD3HPbZZ3ja6gXC28q
yHo/lLDvhh8QKS3oqZur7ylvKu8vd8dMrdFdPJShDeJ0EUPbzTOv2zDWTjsngIZbxrQ0pEcqmdJc
QcZy12kiLniUp2+MAjNBBPCvgYntTA6UAtaMuk3IyoGMTSXLgQurMNSTeebUlAYUGu/r6o3UMZWw
pFYQZec/eXEfCuPVOdFOkl6LqVD/1FSkqW3kVFDM0n7Zly98kXJxmh2G7I+KQrwwmoGpPAwzlYWD
4vDDyNu5AroI+uB8VgS2Uc/cQx7K9DxYf5leGoIOfRO8TxEDUdLXhK3cB2q4Qo4BDIEOVRePB398
flXb4KLTTNzMFqgXVQo2znTcUev7A6+VoRnd6LBlqwCuxH+pr9a+7M02gktAOToEgC+/YQ2mkvLa
AG//EiW7f8F0GD8oZxuUPPUVTgdafnofoSrrsZE21mbAAkE/VQoFOmHLxJE+kynvDE13RdhGCUds
dMcghc62ckt/2Nc5j0vtk/tq3mvJvaGn/czobH9nrTMhMj1l2sLyNZNeki6xbzFHxmo/tJ1c7X9w
v6+mefZkj/9EX2c0nJ6zoPmFjHHrPN1Hw78lb4MK342Ejx06rDfVSpwT9Ba8q9KDpXtauDC5Z+XD
Hma82YC3irlqhN1ySFHODeVzds7TlEOp1MWp4eHLOgEe85edJpJ1TA8BzQVMIbH7lL4/IZD9rlIQ
64ZlyHdmLGFZ5pjdfuoRW8yDAxkQfpf4qvDVn2oC/6frdqY6HMmUBHfIqRSBnuVTP2tS62LSfsVj
q7kpTifIhQzPJBKRf2dmS5dxTI9MlYypYRfkMKnvLu9B5Sixv8D0xyj3fZVlc2fG0FWQRznQmAOz
IgVu/KeuYuivHeGNrT/DYyoa7JWF+yVCNXCb5pkiNPy6In9ljnAOAUjns/jMCft716U3nvuT5Gim
8nmCYNTyU/c124wk2ZVrfDDqDr5dGEr7xbnwuuzOulqLiBqgQbx/ljT8VaVNkGdVPsW212AYJvxm
8TolJh14NbNHrwREHJmZIsjebmgxDq0YSDFfztya7L6/PiOGxInUWFq/jVeXZbqiDMuxpnyAlxyH
p65huLodi20RPIVTw+6ymjP+oULjTU8RDbgFOqF6KP6+LSqweOyjwZ5oXfIzA18ipEQIyqSSitV6
gZgbRcsVNE6gm/+SYwsnrPjEKVloJxAZZR16IAuglPJvZjiURLYqwtVn5AUTne4vo2Ia/4uIUp6H
ROdrZtZMo6SJHixq+vT0apOsDFN5iVPsI5g9VX3O+ZQWoEAJBP8vWpELAkmHhdnBIgV68cTIeu6Y
jDjkJMRCvntaj8YEiukCxuu2IDA8hguDSrHHtlgCwS7lZnI6ChN+AaMFav9AJtwOpeK+EbKh9Ni7
AO7OoVp2gV+IaPU2DVo+xzSHatIZDrXlxrTMGJeEBHFl6lfHWy18FgT4QuTRxwC1O/BYSqCWclD2
7JEwLX5P2h/xxjbtotKglw3ukT4H0QuU4HxpYZvnhrvpbs0Ib5oeil1lyY89ppC32PEeIA8l2aSx
JhtYLC/6yYjyFQAC2KZK2nn/svl6FxVLDrbvb87TyS+zK2OIlyNsHKMYtjKhjejUQgQK1riBVYG+
5XyodDlPuqYhDgRaTaJdvMpe9ySs6pkLuHf/JUO7NjZRtz840vch2QVnlRHE6yn2MpGYRxKMrS/o
/OKymO15x2DNf2QaD+5IrccVhi6Sq40sasto46B/lrB0Svd5M6Y8AG5AKMgWjiNpeMd48Mkb0PHz
Z5nTCb35n/KPT1CI2NLQLqrYhg71PTSgqKoc3aeP1WFX/jNvFCP3FgfKZ3y7HO/WLYt0qHebya3w
Fc7qtHMIEYqLYnGioTwmz5h36DSOXtk77ZmkUbGRNDkvuTRPrX9+omdcELRAVX5a9JknLCw8SJNs
i13d/ZAGFJMaNep2CViNkGfOajeHfRGjJoNqKhKj8uRPMEWD5pO9e39j4MG9ArqXr5AvaBzg5l+l
ROlroe5OHhsoFFTQo96ILMhM6DNvJ8fP0HQX7muqfPJnmtZP4Uza74bub1/+snndVWgiyeuLelH6
zcx6w5UrX4iidvyLiS1sBTqpe+UQ68GxjdYtNjrEarGymJtB1BMPlsO6ay3d6d+z2T0qihtUD0HI
2zxb0sXjT7hj1gcvLccDrlnaszt92QDsECo4YHkIGBpCthawiM70vbrUa4BBi1+807w5Z1l42Bw8
N4F2vcNL3WsnTsu2LN87CNJ8NJZ4BSRQ8FzjrZ5lLlaWgubeL9E3eX4lkcvRe1aQFvdJd91Pk9ql
V9PocbRUHiR1hZ73NcObUjopCKFKA7Jeyu/U4wnLwct3+u/DD3tbh5riLkr1vIkVl2zQkK8yqq3g
a6DGxoTcAxe/6fpM8xpNzkxg5FcmoXKVr1+j8QCYFhfeoYIXMM2t0VfxwNFuqiUqibim0slX9Cw9
a1q6n642y1aoqqaqUSumMvtUEkmcL245wXPRs4aXlIOThwImUKYI87oGQpRlBMrD6uyLtRHfozVh
QIWtTxlnlTRrvhHSvEdNufJkfadauzF2xn22p64okDT05BYKuASLtUUK+DBHM8EQqP6VdkuRLTJz
edb8nvfukS1c7Yv3ZD6MQPKWFK18WyqW/8bKwjUTr+YL89nZaVmnq0cDIWggfo+giwUNuApRFjUO
THsWH+oXu5BrvbD2fQDwYkutRcrCgKcYbSx1DMnWC8BheoxoPMkYAo4EC+knPHU0bjUbbQAs0nnp
Q7UFO9vFucknM/XnDreETKaCsQrjLqtGkm43Xq4+fR2I+Ng3GQImKBr1CahQtoXiG86BqlgaiCWr
JYQ+JJT24mTHMbYRTK6HQM2UAQHs1XYk/6iTok8SpJyc9mYlZwpi0TPVlNcQS+WBS5ZkMjIZjZd8
GNKIcBmqxlGDkpTUJe/04cljQluO1fumeCVxfUZNXm8sg6qjSQr9Cz0W25b3VdA7gADtjx4+gxSG
XmHWXQ67PHzaGAOymYFJqqHcGTuISCo4SVbaV9kR3Ar20ONxr1Zh1m2SsBf0VQVsGK7uqh7ElipT
J0DV1bkAGo2ibrz97vZ3i5r9+xEi/v3wSbJSVl2PEIHOjOD5FFI+HNV6GWudr7SVtkOROuVLqyVx
Z8ldYnskvSwz2BRQqqaQiRtgPqOg6Mjjg4a5uHaVSJh9b39MHPrsbepbLOxlN23gL251vB1W8ZT9
iE7XPNV7qsi0MnpDqEkcxrVSMnveLo65k+714uQhhIE6f5vUtD8VIbpD2CjrdcsUOv4iDDXfNA45
WDloWvFJ3kaw+ORPFA/owVRtG1p5TF9Y7t39p2RjEPp/SWU6X+94HBPJmiP+Lu+M4aIbYNGsFa3D
R+uDjNcFD7pH3UkH0euQgWK8LcWX3RT3BJCbMXqTk7bPeUsqWCQBSYhfm3Mi+mlGxhcBLSRElyKs
M/opbmbivLDQqbcDGcGzFoWxfVDCdFAGucj+QId6aL4w2GGqRDjZFrouZ6C0pT8vBAgsIQzhcFj7
m3tlIcqgSR5ciKjL0gj7AZ6CCT9F5/hjWqfO45zcZlBKJeBsqYcY2u4IiR6FEWLSglxTlzO5DVcj
XOjxTVcjPcVbBXAiyMOKUYD9BHS6F8MFXxUdLUxJwhC7kyBoiC6a16747ieUkJjud9SzI55y2D7r
aye2tBkf7QAfBmwmA1FDSxfcaSqKszXFor6CF7VyOk0+hjytg2YzXjEi59sZAZOexK64Mb4o2pcB
P5mBvpvIn/Mqxkr9/DSGeb41bANCzxJHPu97Cfr0WOkq98Or0atjUw8Li+ROj3csR3+jIzULzCb8
Xae2mCihnAlhio87yr+9h83J47Hnotet9fBBS3drulDcUCH0awgWLpXKcnJujDBHDo3Q4hIbJCxy
8cJ/J7zlx23K57vKDhi66PYDT7ffFfJM5+mRkVcJPi68p9SK1Y9XrSipwQ31RG6ngakYetWX+Ec7
gdM8vT4uMcpnYzhBOXjqNiFmhzGcqSXTaE7yxqMEM40q/rpDCNFalVKMpQvR3pQ0yP9fepGBa82H
mnIBz+l89/YkKoDdc9OpCnysMijqxo8AQlkPPVHqGlLu0QhdFffRdMa297RXzjlqq+tPBn5aApo+
VboeeG7J8gUBHnYc6hlfenpYihfMsOjP9lnGp22MVvHXMXs8dSGl6N5EkUQM3F90aZk2RIgQ5ZLL
IZIBY2AaxI9J98xLdeQ6Dn+WdeXsXTgToY5/1u8sMSbkE/W5Eq5E7XeWfbRrU+4qgxwdo/PEPJWF
ns5EhdpC34a8egT5/m18ik5zCN0XeKnO31tn9PM4+qrHT3Py8L+ibcVumUDHcLAEGcimzdiYl2ss
0+RmD9t4VJUSMZ//tUO2VWGRQ3rv4dV4OQKBH/Ced2gQepSSO4LCj+8zsKwhQG8XZH3xbNWLiTiE
cG0s1Xwfj1pHVPMhehN0TTssBtubZK6zHg4ZxZhMDaGH8fgNLurIqBbf6WImSC7K3tcXCSxwUIY8
0gS/yV/SGAywJjHa8YhrN2qn5wzHfFi8KRXT0bEMQFPr6EtJ6/07UqwAn9MyuuwA9QoiVOPh6KR3
qAYNNUKpWw5Tua5etpKym/JzWXkEOcykuHwhqgYUXv8YHEzclMfqK2oxWv/SqLKukc2F9GyFknGB
kM6Q3Etb8Q2OGe570NZYJip/8QBY8EAZqiGqU3itsRYbKFdbGWeVM/OLHJPkDjq86Nf2IvG/umtC
gWKxx9uIMBNw/DQh787CncLbKqJbZvqmLsDyXAU2Rh1AK0u1LLYkqBnPUfNbctXVv5RwQrhmhKdb
jchcrAhuf5mZCimQpzb7MX1gHYFR4vuvV4yQpnoxDA+dKA5q7hogwrWHMA6gMaS4qkP3gEi0rk6d
32uF9t38rQFMxbrRuvQX6BIo3Hk4lrUXh7oIY/2JeDMlB7Tdw4Oj66yU/W+ac/GsSjh0a7+sBoAG
yKTmaL3AbuA+mlcjqHooRy+X2cERxsTqM/psxdo5ZTj1B67fGOvx0vKdFuaD3F20bif6UYrRPW0f
DlapTzzp/OyzjEHDhJ6o7EpKI6jZ7US7nOcupflzuLvZ8LpdXOgl1Aeov/ZeKURDwjzEggRv2ttW
uZVzaWrWD1ndEZ5LlNnACuQCkzEd8v9tCd3mDHbtUR4QfpoJl6qiMjuTmh1qsvNj+vHlGhlq2BGa
y9/Lw8VbxcC7E/9vven8EW551rqP0mUpcBBSa0QWjVF2U9HOJMA6RfszsHf/pwfoDEyI+W4/G7Pz
dIAgNQB5zbkWCiNkDnKQx+M4J0fQeYcLdb6XHa2Q8Jbyu0Asc+mB23GLacdEEKAK/ciCwNe0kQXX
mpvr88G8wBnF9D8ou3eSDvmvE4+1cFrflGWJT6KkhSRLSZ7Z6sjeDfH+/DtJamYRp7votoEViReH
59wWY+n7pITVFpgIkn3d6seOH7+hTSEk+8CAWm8a7cxP8FtlVmIO+0O9rWkG+J2NyIKvEdYqTu8a
fv7ridruY1Wh8lFzrEoouk3StUvX0C12tB5BT3RGTLEaWqU7xxHSSEOys8ZDQ354K0XVAxrKifF0
qqWC/Kj3OMYvCj3dt6Z7mUOJHJJwtSQKy3CtLgCKK3ti201EmzetfxiW+WySd9bqsJMItfuKyvtT
noB405QCBJb9XsSJf4HiP5Df58kxHZNJbAZU+vXuIEf0jz0UAFIT0TX4NsrB1jtEzSe2OhAx4uPb
mRe2a80N3VBSwIluFza8tuaLtyZR5r2IJcBhHghzS/Yd0gZoSz9kmpEYtOmLhAuYLLsJwt/XcQRW
H/iM+9i4oXMfD2m/tQReAaQdHkpmJbEmXtjh7F0eh6vOA6QNQUKztR87bPWIUA6xErhu9ASRQURv
l0Kb1exBXNTMYiXcpLayNTPNGqkBNhZjSR8jH9QWhOTi8Oz4qKWlV97ajO33hXIQGWScAWi9Hy7s
GqJ5s/J+9wDr+FOZNIJTpzUXQ+rv9iEE9yndbOLMfmRjlBJNM53q89fYCgvarnMwec3FiCwckuQ+
4JqWL+dJrZoeQJnNGr79AVvXH8CygtBSMy9CM0WXtoj3VOe3Cfbo84v1RDwCZfAf48XJjnMNQ9dS
356OsNrnxc2cfzJ/Ewrcfw5YzjKuZmAqnv+UwQfPO9OGpLljn7RV5YZ681WuC8fMuL4roSp0NJ05
MQDWE56wC8ZuRHMuI0Xeok9pAA912ACyKFyP/qQHuvETRedt/04zI2eSN9DnFmHYKPb7EwdU3QRD
NhbstOqKDm7mGhE2BVZATo4Jr5FkbFuy8MSRks3/XwEYJL4nyZPqe3FmIkNiEvD9yaUJu2CE+jdt
3URbVkDgZsB/x95Xrm9dFQZ6uq0zCWlbumSJP9Szd9Knfz3ioI1Kx9yebhlOhacXh2CJ0NNFm6+z
cMxcr2mrd2bTUc32ZR6nEMglIpjBDV4ERojOdT/rStH6T98CVZ6q63r/1bS/8G3F1wnHCNcsEZQG
sH3EGMFo8NsWLb64JBpyiU0oZS8OyrotyaqUENPssXKZ7zhdCUtfI2aMhRunIEpFoMwTyTgQNPvQ
eeOmG5DHHcz4Y5QCaymsoxOiaU1gF4xI2l6kJVZHra3T0bhAckAmJvlfVDWswaqNd4L3c+BJsa1k
/nmmA18Pd+LIVFBoX4hLOqfaowqt3LHP4YpTLkbYO/EK6fRFgtPvlEWQL3Z0RK0HYOZDA48Ll3Sb
fvbL6LW6M9MNHgz4h0S3EHuBe3sF7rsFRzGOc3DBkPA1qWw/eSDntfpK4N/aprUX9Mb8awPQi52V
AiUdvX5yYYIyPMGG6lTqUNPBpxEaVqM67vE/gW5xvrY1P0z8+coIHgsKTFPr6C1T51LEio+MBhPu
UabCYjxcnx42XK5K4BwNgGBEubfduyarQwwklwD011vB60gIhxHxdUqDG9dRgfqboXK31F/TigkY
9ZingorP9Ktpbsqr6S09kmmQQ2+8/ziKhpoyZUmrlIKR40/La8844d2qw0qgDgpB27DIlilv142+
CgM2onxDlJNiLuuF5j+HkxAYAmm0IUlfbvkDRU6CN9pqOxrODzyyulKAUQKg0KPf9r3YztaErB56
r7KIl/dI23iiSm7sRQi5ji4oNF11md0cgMSi5Zs2no4FZMr4dkVmhVZoVRJKzW/kN2rJBXAk+ScR
ESBw8O/4Cjlf5m5gUboGYmbHrcxGi0PEOyFTvXvmK/JCz3TtuXR8YdwuLcL0KOvMbHofVYbxvMd0
gcg45NIBud7Kqd2u5fbSbjOFwPfJFsIPC0ZA3muCrEDrz9MeeJTW0+5Vk0Oy24HyGhknFuGsyGYO
fjToAO12YfjHUvqNBNSA5WX65hngpxY2Yjt733FjmUYN8fGXNqHai3ucBFbpOw/IRx+QHznLgsGb
45nvvuPNTl2UFkUOJhr0u3piteBXlNPWAMYQb9uUnE1vfGbIfg4HJpayivhOWYiSx4JYvKToxLiO
lLLmPBt+A5lO2uQkI1kdjh/sag0DKARen/Act9ADItuztL3yalYHE6NdP+vdh6l2CIbi52VxYIS/
ERyKj3EQnnNOBaCAIurchAAPqRaWg+uFiNtfoOxo7QaAVn0YbLF8SLsPZOr9XaEdiTGCP1eGMED4
b66Pee0QUsOiOOdErUAEUuK06Iy0k2tFokpTEDJGiBDB4UcW2Az4yfpK9qyPGlTnHU/rA+PukP8J
+BKNpCB0we7+nHJh+Ulq4UdKwv9ZNv75/I3X1FrmjikNvKcUsMmPzm9p1a9Lpcqh/5tAZXw58VZ7
egjNFySlUgX5YwFmFITFsZEh6W9r+smDKzQesO5FIOrFSkM42OHhkcyA1636qtVVDRUh9HPBJN3t
9xBcCePyhLPK5FITwGR0jM3P7ThIHv3OHY7ErfgcYryWb/VVlMYOrMsextVC2sHSW78ytlxmAKjZ
93zG8LRqFvE0FUrmhHOp1UOgOxyeBFfe2XFFFN1DEiRfkuHyEPzpOgZtq5CmWvPQlbhCO9o4w4Xx
Qv4jU6xRjcZbQJhS6uhk+/FMrTeXGDlfiSusPqUCY4J+hWbxyn2Q7EZ7KuaOUJ1vOj727Wnflszx
KPyaXJd9hlqmAxexQwHPNzQIrembEjAnYjFRfaEcOvP1w3aziXeyWNDvmZPzcKyy+hYVoBnwzlmd
/v/GUznWK1gYj0DILLKZwOlyV6HQCs461iplOHTk6n9DxICNSjW3eGsxZ5i+zESBxpfwmC2m0XMJ
vrl2ll8wWVIcOHCdhs3qHrgpPW4RsqFfx+kKL9eoG7ceLxUjVWotrNMUPlgfwI0p3+EBMXSa21QX
hMFsormnjdajf+Wp3e9JcMEh3DJYuPuhrj3QXFrKbeuw3ExLLHQnRqdnWSGjUniW0WJKJOIsgCBg
ws29PUJ69JPr6a8Nq6yZc22fvKE356eWNKPMnjhryeUCfpLHVdBT7KSSyzbryK3jgr0eHhkPKEdk
BFtDiRUTn0b5Re31R56e+ife9xUSd1hPLKE1SJTlIXpbO4/DMxJ1u5eUJZcA3QUDReieCBhaIuwZ
eCWZwlRHrxQyNvqFViEM0UcoVhsO6duobRhkqp6SJOtQJAZmuOMTdx54DXtodgA225cyfHGmtDSw
RGHoG3RJ3mVPxtS1s4jgB0zw6a8RCWXnpnufn8I1V+f+2y2fU3Wh3dZnccRbw5tX764fztl8A1Yz
3Fb4OEoYOWMGRj+W3/CtujbRFkoMbbXpIMh9htaqqDjZvybjmCfKbS5s9dsXnTStZspskPL25D4O
BOlFi4STYOu1hlMbAs1BcbiLDslHFqAAEhXC8oGVPVH2j1qkXlx9M5HkvkqDyldU9G96bkX/UTZW
muq/qyaAgP0+MtXaiK6JH74XmiqdT5i4Luw3UIiH4RzGQKDATnGavJb7knIUyDJ93hCF4rCHT66K
sQMgtfhxadQI2vC340yXOaKsL4YlgTbwKr8peaQGU4b3PyVxY5v5UEAAC6rBkxqQlG1GO4n3Qj0G
25p12ZxVUGoLw9LYuAD46In9hdyXXGYq6nQ4C4JoRJgpR9wurIFUb2XokmYlHlMCiDQx7eCjcOc6
ykj6F7qzrdgJtk7jo9xvlrgWlDektFW6ICDMstyGwphoaX4d2vXY2qFfjbfVUwIkwVZ4n5w8Zsno
iGGlgynj5e31cOwd9Xsdxs6NiY1xpcbusKioiZtBGtv/Sg9SglR77d6vbgCODJoBwIdyv7YIavbw
hlluB6sprKv/I93HRMsXCciafWpEFt8UlqPapXABqLmA33WZZdE2esv7pUpu7DZBpFMsActAIX7F
MxJW2/gp3IYN9ZfNHHjZrVmaMXCHKdthm2x2l3/yGWQQlwz9MkAeBkXhuzsehmBqGU8w9OdfskH9
L8IISrmYu9nF3Sja6u2nkUh/fnnSZ5JBob/c9jKph0/1In0SLbh1erc/nBhBVNO4Tmp9VXJ79i+U
wHD8rRpMP35sR1Cui2zpu1S0wkvKJ7GntqTWaApICs6X5Bin5k4vNX7Xuy3zRnaqFUFmKq9o7+AA
3XPldDAxHVaVbDQU520tELlWPa9dixSN0WCzwtNSLNeGwmDyn3fbn7nHyGJUmYVSjAdFRDUSEi3Z
aeEWJwDCHp0Qu5uSBmvOKUKcXI9hZntdTU7ajqyJlaMZpcKIYAZwBzHBlyike/iY9i1cxT0AQYuq
YY/cnKRIEII+LsF/qsR4lc5V/rPPN5aStoIE6V4iBTkk0OjtqDiGVVt42OHo/tjlHRNUQtIsBx08
JVg1JnosbnjZl4WO975tNREdc6KqqPY46OeJEEaWez86faP2ovpVIw2Naf9oYkMt7nxDb0P8oZ16
0D8pkSYLu88qo2S3ikAYiHimo7eMnQh2TQNHBuP81bW2ZD7bHpV+5Sn09x8ET6Ph2OPnL6dJG33q
Wlm8yEZZXEYA1a+6NjfoQXc+7RlA8yLq43KfpAN96xL7gDxpjK0bkc89pRgDmH4oUSB5cJyhSpcH
wuYMEtLQKOvS/u54AzpPB405qUyfzAgI1+ypSZTdT7yduC8ZEtaCEgyXwvaj5Nq4SiIwgtYg6+Ra
R5fdSs3tsT3HJ3W5ZU4hQqkMiv3pmJ7y+dYegjK2MXvhPyN5WGeCt8uyVPd02FinPkhZcnDb32Ja
mi3RlNGE8oGlOY0Plvh48/imwiNA8zkXlL5CEC/EqQHZ1GNUSUwN2Gh0RYXRRuUgYhI8ubMc8b2p
FylGZewdzNiSbni+Ngbw8Iak1v3v+VlygB0VmlnM8MC+B6dPyptKtXTZPxfxwm22kT+zX9kReUfD
4r9cs8gOjT9L7qEXiz9BR2R+cEJh0CCgN7TpGEwfqteh4His0S/GVX3gZD7w61QX5KM48oKf/nth
OAoSkaD/Ru6t2UDhciSgKbtowrmKMSmk0/Gv1+zhXD+PAj6akNnnnDNpo0s2mUZQHC62/SHwX3sB
vWsZNDPNp+0wlFQKGsaCfOGMKEpcF79Vl7wP0upyKFQjU9jQ9mOoqwHZnaQPx3Mf1b1EhyzOS7xk
sxKgX1Wtq0IauKlghoiZdtwz5TEh3jvceZyJ4Zt1tTW9PvUktI55wa7LqUooZ+nw4Z8EsQarPRH1
8JWDKeFva02qzpXgucR2RjzAZq0uaNXf8qDJuxdVwTDPTlLt4gZsSlJpRdVnX8iLkziTcc+xo8I3
ebRd8jmJ83MDe8vDfg6KNYULExNVtEhF8jb47+Oj8/J0IPeLY1iydsryzXNYwfr94t8wIju0LJJx
+7x41/HIXLzQtjkqnvyPoi2iHMU9db77YbkMYZj5FNEEJ63m1y7l8m2AaoFj8N2XvuYx2y72cZoH
8OQoj0a6RxiTuHfVCjOnxaosSHqAfGncuNmYPzt3N2DIAmHH7416GbewZHkkIcLW7TD6h9A2ZNxF
nnUcS+j8tvsf4tDJZIEPyT+Y4YwAdRtmNOinLdaNtM4JxPnSvzS14y73hxhZQagbZN9oM0l/hPN7
4xrYzgckQ5YvXta28OmkB8cAPBzIgn6VgXIX/XZoZIFjpp2ldVeWF9VCw19zF2+Scw4JhuASQygY
dx6M5+/iRTo3Hj3rHy22FuhBRNiFBOukLUwKsQkCoXFQJ4LDy4qrwZtjkzsjAvMdyTZ0PacLOBFd
juuUDce+wNABmxx65uZeTMeAgLh885BIzJO7wKavpI2vKvkovHnYFHzejEymbaxz2pAMYiM+UKKG
rCTmLtaDPtaDhox1CIpSKIJgpXctpARlLt34aFKpZKClM8uBfdoktdRemVlSZXDL/ilgesNNHErn
L47yhUqGOHddgV6opHX6cd/FCB4CNdw1a3qNhFvqOoif3sYdt5x8jJgeTrS6LpqeuoV98uNbYj4A
RH5szxSD2Ih8+c0UkmkzOxglOk8DXE1pS0HtEgUdZ7HvrC8ICgrx3zTVBBAu1zerfzjapsqi9bzD
XnVefwGtNOQepiCBGqyOY7FruIguxQkRVGb0UNZcSrP7JXW9zUBa3ADYXU2h4sMPA9HU4D1Z03Yk
aOGx0OlLLtsRz2HSbEil8io+u2yaIMPBR5OOg7rD6nfCmlJHhDT94xB20rIaGjHbVwEuAgP8s3G8
8t3MB57esJBjvyM3s+x7NRRHOLpmmbAIa7Aty6fh6GA8D+ycYaZCQpAVLdLnAWj7F0ssXnupgMvd
RY0OHcTcdThj6QSpbEZTkkXwuIa58r/l9imMf0lcMMQO8qAq6O4GN40Roek1TsQ25IVV1upVeQfz
nSVx+7pQNGRMg0vKEE0dKo6rS397Rf0b//PdR9fkWqIQBz+3PkYaIsT7iJXrftMedbt3VEzL1/Lm
YUAHmb+4b9Z+GtGvgxbdQG8paHGcr3Ni53hJAoL6OjlKqde8wiA9C5+yk0SjnMIxk5c7c7GVnilg
snTwEY/+95QhvqhtRfMjRL5PZiyNdhmmga/B+O9HMJwM2dvbZ45PwcVtlsLG9LsMvFnXXQZIgiX5
Ysiy3zWa/oEwmIRY/483slXBeHdnAtwjga6/WAmPxHPm+MvWB1UyT9jLbRS6OtV1kwHgkAA1vD99
kj5yXazb5zlkW9fRHs9SG5gnDw9A/vCaVkMm+OxWaJn/MxXn175cnFhVRuoundXBI4btTdW4VpPd
BBhmg2hgPI5yDBguBG+l9Xdzyu/4DzxBFHpANqtxgRM70eBhWKOhst+HNkRtI5k1VIVJ4eQoYLM3
PV2ZV7LNIENfmAWGgLRHsiIawNrdPw/QdzZ4cCqDfHvTUzbquZGa26YOi+qGihdwOIlrXEO2lxJB
fuN+/4EmE9k9UFFMwM9489hPL1DKE5sMH68cp02MTxqghvbOQyCAudkkwZXyJNoHMcyxel8uE0LR
JKQvc9iUKJEex4qh/skY0CSTy8CwTclSPlqjTE/wy2QHKdGzy0TcZyQrU+ajdF86IxZtBoFklEiL
gFTAAr5wDxBogQs7QLMDoKq369MXMWI3l8rQkW4q9mhtQPnfs6auRk7KM9UEr9/VkDT+IRXtosZu
nvJjUwbGKBA6ub6VecBjkFW5vupnQ50KIAPAA57GAuFdSq3OiMzglSjTlUlbgF0AZzqnEmbrEW2F
HyrkyEE1WqD1e8w+wISyR7px4bLim4bfB1CIVCnU/glM/A5+4PQLvBea04uow7In9GcKFgHWlKUp
vnwFy5cLbcPBih1ehUnNVGdgpkvkwtUEg33SF3TYBOtXpiIP8d/QKLKzANyz5Qna9t92aupgoW8p
7X3NZqhCO/lFqkDg//9VtGZwiDZipeVzYyzodAZQMOiRi+o8w845FTtpd9JebN6+cFOtbbrkpLCS
cCyypLX4w77CJoOUHlvX/5HngN2OhuX/1ePdKRzVUl7SfLlUQSJLdLG3bSeK1Vb3ZCJQYr82Q1Qs
3z3MW4dBsN1dv8ZFq+NA+m4U7d2wmcGjsEyr70AqIVAy4XtLWtsoXdHbDFXR60aSyVY354RXzyMF
Itzawzclkee/Ztl1+DfeufV8D/onR/qWeZ1fK+nyT273afctTyya/mdlGMoEpS3wWPzNyi9przwh
MStPLiB2vti/QRa1DfnZEvMAaOM9HldWCAKx74tTSksNjl+tLPfI8pYgacsJF5Ssnb2dYElQ9ONl
3Cmg92roIIsLll4XN2g4zZgZtwDq4UyAgKc9y9JjuzPR/W2J3S6JAjYq1gF3DzezAKFv9pTWEFRE
09wM6PxUhIQGX9mvcc1304uKfUYrB43sZwO3RLqFtbIIppXVlbo7jTbN1CO3xmuiLVUiUI6chXwQ
2BtNR2JfXiXKC71G/fAOFT1G9J6l4yDjR/uNzhEyMEULnYQnFAt4vBoUg31PuFuPLfLDZkMgXRd6
oBYSHvCjDUyHkCD2cITa9xznUe61UwmSFR6IQV714qI4qEgeKrbobxSi5M+nO2wf7D383Uc94M+0
AUlB/x9cQEWI1oKS8SJRE5tTC8GKHpC4UF3smHP2Y3MS01rLhUSEm3pgfZaP1OpgFB6+/OOu9Mp/
Hc85cQK4/VH0NxjgaIYjB5G7tDK0sQqLJLjNgaGwOK2+qrtpguHln5Xq+tN6BPMDmOse8+tUjHnn
M1NgV9DSUdk1wLdwDnjbPyUy0W/ys1RPtyy2s4luLHMeTW+6oxnncxUSrjfsUZOAmILeHRDUIf7Q
+qM0t8MapHOer5Y2Ir4vcFUlMqEDWCTQIx9gjQVu/0X+Rug3/z7Phe0wUHSUIVa5uCaN53gesLlO
e71uQ8vGST3vVRGp80BBwhbFbmWzBh5TLHeFPivq53rs2zwuUzSVkK7q51EeHIz3MUuHaEsDJKzy
QbKQNCJl8yMI1t6TKODLBwJRBmno4pqTGamOWTrt0N2VPljuYu7B+MvF4HIj4cwZpC9tbG43VcRx
VBzAyA17kvjJvG2G8+gTQ6qKRCqUYP5U9K8nBKoUZM3H7ndR+sPGX/La9GPMSY161yLtADulX6xP
bHhNKt9+p+Ir/nAKWUyrPstufhbzW80ustVENhyhxDY6iZB66tE0P+wKNBFE12BdrhTjHg+Nfmha
qNgTorgO0SW/UqPVUpCRYM75jqyTsQpWwPfVZERVPpjKlZYKp0A1GbelgCDvqID6J9JzLNT9iNbX
WyuywWebOBwyl5Q/YtYw2X+H5FljqT7/qXmdWszB7uTLr0e7db1kMQFDIOOW5K3foX+2qRmwCYSI
A75yh5lPiJUBJCgzo1aA8L0jWLWuSei+Z6gXyI/vR3H4dTFh+4b+9TtbmMc47anYE5QBn2UMg9NZ
9axyEn/UVOpMOLjOQnDKP4N8wzBuNX3lKLWi644Af7grAjwwQkTFMMMg4wBcHC4SdqpJRpIeV2xK
jCFCicA0w1MpSGno1E3ALO73ngqWxamtLL45fHMa1ipZNugFg7W2lO5IWvHlURbpjxZ3YtHTNeN9
qq9Q7sA26F0yUEyXP8adBUDNNqHI9dOcQvR2xyAYsfDDopKmgMWs+ycPdHQghTiEz7m26slGChJG
lLDRstMXgY61eE3cET9s3XMmSo7GO/JNc3rEQuKrGg6Rcm5junveyngArNKQYZXe2jbdB+PVBS10
/WhK8FwuGKLqTC6uJraSdIz4OHopF33zsL/UZOvn9p/7vznE8rJeuYKyW3gf0gPJRgyhhDh020Nz
72nX3QVRgLcXavfvVR8LXJrmQnCfIsdBv1LuKRpvrDzfEVkaPRI20XfZCztqEHUNUCP5aDw0G7Bv
gSUfLcw7GgGbnmQCesXPJ5e3ZMOB42wFf/tW0CXy1nLxRfh5fvDHpV+he3JzqI21jgS0BLNapqW1
QRhQTuWiylzozRxdO8utEsP25UaMJ0oMchEcrh/bwBhpwAPuSbxwwNHRBKIWoBxBQBzbjUbg2XL2
6t4N1qmRRAjP+O4G+8V8MIneI5bKYzpHix8aOYbw6sQRchrkm/MGBwsd3Gipg3c5glDvaMNQ5Pbb
Z5GKjUmJN+RDzaPOdN3cgz7WFqQOSHLH17xbBos+RC6M/+Iv2cqoOJDDRWT/giUmwUVxup6WP1lA
H+N88rmlw9y0dYuHKuvKsYO9dEw0IlBUkVcqIIYNyrv35cpPqJBjzIe84qeKlxT6FmjvReX5GBFI
NQjDNSLLZc1YHkX1aqUEG9BTIaO5ikmdsfVsx68nqVblPDMhEtvpFeZkbP6YpGmAPI1ZBiYxxmrU
S70Pl0Ig5gju3HgXmhQpDZRP1DULnlQQXLZuFXAl3bYEu6BHOgmTQWCkzDnzw1vLE9NHNAu7Ce8C
QZiFmyx41yNDG4m3arwARI0LyN+Dhq/txEIHghO3cic5daV7cYD/PVfsZzaEybyYcXZDxqeOC715
UdTWWQnLVBwvJWTTBRsv8XU+mznLDYc6N1FdZxfq3m0Pc4JCsFFF+/76YmcEy0lbgP4quoR6i1BB
JvCcjN7jLVZU98hEBHactEXTWrZb6T7qB++KWVp4Faza3hhcT7JLw6Id7FGYOD5F4mXQARLaqJIG
O0NESMhyIIf8HzlWIHSocz2TTSiEorwSWykIWn/xLSjsXoX0ZC1GWgYYjt08U61n86UX8S9rqHmr
1mQvSbtxITXk0g82vC10iDTXFQc/Jof7ejnOHZvmn3VfB50iCbWG29cNcxatx6aw1zfsy6O20xUK
1epkhU4YsbfOUSb1/V6X3RE6dDvz0DW6p39E9YYxPmmOtY/BNIVKNrc//MlSfIUBIie6dtpzhP6Q
m/ila5umJQ7d2JEzNsGoLGjoiHZfSnBTuTS3aL9APYzZe3FSQ6H0WBDi4AKjc8XjjGGsm7yAix6z
Vj/WGPHH/tWqjAIWWRw/d54Yugu95E3+OYW7UYQTLrXE67FGygA3bTGzodAoidri442VOrncLWxj
39E3aQnofoDydtiCrpRZ1lAXrrfvDgYdJk9A+t8QmiFn0nGjNlvDzNwV+0QtvP7ccyHoIV7GOLAx
qR8xGY+3L4IudkU5PBhQ599G8NPeRUIGE2qFWGPllo59l/KkUhy6YwT0o1PJF3abfTmVgvNXurjK
51dSvEnVDEZsvS0GSfAb/uSNY3wpJz3iN4ql7Qgky0pGYcyEERmEiMwyd6ACpbpcrW7zOHX5pmU+
RZjN5yxsrUhhbv9JaDmzJMG1+Oljkee+ItmseHRzuIsyr8u0tQWVjF7lbzYSHGw2dpo/ayocXNwV
AZl0RubI978OZIOcF3KkshU0uoY2EjFGfjl3SStG3lWKL38WIqr1THgUO1Q9BCjYL4zTQKhVv/6F
IQjXwPhG+t74+R2FvidhvphU41d+I8G9+UklM+/9BJzCr1tAX6qVTDhvTBtpB/CfYZuQ0TkcKpVd
lnP7f+yi6OFA3DBtYTu88UyUw6aqZY0uFveDNcUtCnjiI2QN6fuF6Lf/vz0VSTxYPLZB2df2RpNn
Q5HS9Ykip0vKQTGXbjm0pAnPAhE8Ix8/SqZGrIA5MXUyS1J9h4EWw9aQXfduEb7mwsW6351KaCMj
kEqvq5QlTk2S6QmYN3oYHPFSyIKztqUuje9LcowF0w1pc0KNh03kay1dKX2Gn9heosKf8Xl1idHN
tMl4VTqJ1fT9eN/LCyaDqoIjYzxjWJbLUnBov2XrtU/iT3/hP0bS0oaVCS5muYFv/Bvtyqf/qR6O
yaHVN4ZF9ada3yIQOH9aT/U38I1+e+kxDWMmFPmISAjDVPDBfOsHDpM/qG4l1uEGRyrKSX7p6gOS
MwudX4nVx/jtLsMWTjfA0OjCtF7hzw2fa60O9tnRPmQv2Ca69FFZ+M0mqFDLuKZ3iNxjpAGrRuuR
+FXqn5WITYY5m59bWmhNJrdmzZXltly7P0m3YM/Gx0m8RLgObKId28kSLk1tHlGRcoVIEUDFBFro
LJVUTeMqAdSyZJQhWGJQUiBBITBXUJStRNEoIsYsK4RPWFu8A9M+bHwY2DcVDi9UXLp3KYfScVd8
GboovOadOuiKvm0jfudHKa0Uu2CE5oFkF+cXPtMxITF0Qqaz3VegAaTLLYklqpaIeHRJqkPKrk10
VAizo5BxwgmGC9z8ut0257z2yyvJ05JWCiGWc7R5+Ib0gmgTnn0gO/+Xhf/34p+dKqXl66/JL/A4
p3ayz7NDbEkJRvz3Pxdci8EotRmaz+iNIIjKp3ScpE/y0Enmq2pUEW3k/2y2jpstjdPDONVtsAYs
HPjXbOubgk1Fw7XmsASIJWgL8x5UjIZNOldTDalpAH3IlBok1jhOkYzzxl6xxeYWQSI89i5NeS0C
zZkZjdxgf7XvkrtsSpDOZrEUv5XzrNkgVhKptDknni5F8VV8OS/qPr6PM/t1N9ZZmMEk8ovsSPpR
0t5qtOk87lNo+F55+gdDSriHB5aH6aHarKUnwnszt2zObQkFw0/04wO0Nii7WmpuZnLPLrP4xCVa
PsFxqt+4yOg130P4U9b6iFTO4WpxFdmLSAGA7qmnCjLesx445HrkdEMf+05zM5DEZ5vaonuyx84D
Lu30nqLN4lIzgaVfkvvqA2Mk9prihK3zCMm+PY33+GKL67pxDShAlhs+oYJAexUgWViEK0jpmowc
0nXkW9avjNkWvLarakXPeKX37KzRiGk2UDV6Pj+2K852Hp5yCUR+EG0RFnOWYZc74AVSkwCbsSSt
oUbhTD7sv5VejZweIvTJZCoiKtzyGfPpyN1p0uM/G0sTvrowL9aqTWKfLILFe5s9iJJQG2xHuksh
VKTuWWj3ycIq1j24JXQUSmSsGJzYE67Y3wUP4E4PWl6c1OnLnvpJcSfPRsUTxW/xbOE/y2l03Wfz
EOLdVLd+NrvWpOgaMBT0t4yHCpj8Pyu/kwfyfLL2y+7Kt1JCQhnYGLDvV/Xj0RPeobl4aX5zn8cS
fXT3BMfRVJhYVvxeKmmUF39o/V4vVPNm2ogEzahL7mQ+e+GWwWFHEaGUzNikt/vzRWra358JhoQD
mrRTSE34yUUV5xkQX2OSx06caqsjL8EKxd7NVqiSGFfhMXLDHh6WLHQr6e+jWznFIToMKdENqjSn
pVybkfMDr61jdboWjqW7FD6WPpk9NKOxRKvVocdX37cmv52Wpkpyldp6STNsdOCl/BS5Y9wCEPMt
S3UMNW0raCNutXY6EiBxuv6bm7j72ST+SV2dGAN3K+cD+pkvRU4xbmNqBymJrn/STl7IqebaEoyw
+Kn1uffmBTkcjHjEAf4Bqq8c+nOUtZRITU92PeQZIdcbL4cJRkhYsoF9tzSea0b4LuzdzYlXdrF8
utGDXwYDRzB32Xnq5fXxeQZ4FDJHmmd98XY8MW7Hc37C3ELDsZRw6byTUjX4Aj6R4zZD3ugmGevm
L9pyIj5c1C3IPfMC+fQcaIaeIF8SUyUkkr76eR/mU2F4YwOisyyJ5VhWD8Zj3auZvQjdc3vXzWXc
r7hsMjxt8KhO9kmIGgBwR3jsHmKmCj05dJMSUDtRc0sa3JubJgSI+mCXM2ovC8AH6QWHt9JHQcP1
2IGRJXwjLuVgEdaEhLSrTCyzNUKrPyDDcANZOwbI1++grqnxidcmdu5Tf8ahXe3OUskDMLHOiw/B
LtxxgEPJP7FzV8NCnCYWNVDgPhfoUWoPlHRNQ5XYaP/1wtra4KTJRV8GwIMD6Ml3TClRqT9KQHCq
HpbZFougOtM7GAiQAUhWb8SdJoMZNztBviK6Poup+RsD0pw0Z1vgIjrW/fqJog6lDdfuorSgiQms
y4YZiuVjKwDljvfho627801iLpR2h2Syzg1PJ3dsc9TDFv8VVxxnupp1o0aZbTYjdWrNCPNzse4x
HxM7dQr8PfVDAFCAgZr0mCVBS96Qv59PzhRor5qcLrZO1tkmj/gIOe611A94hv61tRMXws9w+Cps
JmSG3kJb15SnyafpfsyXC9C44zwgooXqAIIqbAbYXMZdmPxcYF/RB/uXL5otSuFiyiFcIZvNKGoC
I1wS2kfUzRTwSP4P7wgR7SuM6/p/YXNgnmn/Apx3uAtYgFtMtSD1byUchbeTEpVbO2XSpfrrP/qS
PftQNO91JMIk9WWH+PL1L3BhmmZ5/uyPdWptD75XhL8xNaG+UnbhRmGDsyC0kZs6SVRq/x7ytHKf
V+yZekmETvW+nMr3lIdh62e61eJnbDYUvtA5q7/bOCNz06c2hh6hPpTF9plRGAuGW+WGMn7MMPxw
2bFCUqxQWnH3darpezTHrSmUDASpbgdsio775DK1FXwQwBedO9BhOOReKDxnlLICUEfVzX7qs8g6
rmUr2sTXBVrWfn2ENa3PorlRyrpFW9JzHZSQDtZUJb+ElCLyFYwNVHPlaITQnL6Rngo11W2CJCnG
95dDZc7em5DWbgvEIuhbjxmNNinatWoKdeBHpEqQtB6yHiF6yPUweTyHmiVTIRqv3uYWLHlR6B/W
h75Z5mcYTfVfQkT+l6OP1pVgR5ZaCeeFfAE8YHshPExBZUXD376+R9DF8MgAG5905OyMdZQ/xICb
NudgzxS9HuW39WYTMBSWOQFKoyGpg/CcDeKxJKuFqqf1EtnKhjcLLWWQNuNmuArHiSkvjWofZ88j
CSpggXDxnlyZZ2X9iT9g2kjxoIgv4t5bm6ofU5D3PxFBtbM3H8a7Eg5VhsCsmCxqd8g64FBVsZ7j
i9LpZlmaTy8eM1wGc5OgV4DTNh/BDziGKVZM02T8eCfG6EXVt4gqbe7FIGrK9wpAf1pRqEW9Z3qb
sLuWp446JLnPZizkklnwIF3EEL6wrPZYC5GPwgZltrjXVLPVOL+YJ3b3F1zLyGFQf5TryM9LdIYG
WAsRrPjIkHfySi3NVroP5T1itUyocrp0jy4KbULwqM9SdtCC4nRm2hMY3rZOt5qQKYtN2rWsnsXe
wZ7DeNi6HWSuW9803Q5tLpg1HZIwLjFopKTvNJMJ5mGhypFA25HUZvVUYUCysFKBYvEPKhQb/K/O
ENOA8xH0m1HAcM5DTeaVmYkBmHy/lwD8kXelYNXmL2nUod54OgKJvzzkYyd6H2E/qYQHJEDhdzJM
3VSG8NzTMYyNkpXDfm2P3mNVdtgybAKEKHXhhB9CN7MDWa8SkxOg3LIoYTJNnsmS0XURjDT7CmUM
iqVK/btSApli1rrbd+T5V8jTH9Dcqp+7TBK4yD8WKhHKs7/Hfa7DPJqgT6vI7pgd/gPd/laRxx2B
jKq4Xrublu5m2I17b7WlJWQuIJgPgqSY9R/y/bBKIyt9c6WL040RcuqoLguasUcMlfBKth/Z9lwi
N3vGt4ICgPfCR8TABD5OUpOyaambtgtTTyRZC2lAFqfkEDTZ30Tbwosevw1i12CUGxI15+7eBwpa
ArkkBdFi707wxDkMqAQ81EvTI+MAhvDMbSdmfw1KMpqiF0Cw0dMVc0BYkMQvhp7E7+VB/BsEIEuM
95KmZtpqG1/KIhI0z7r8d6CN/4CDNiGVUGJwwjoqquwNhSejE/ZBaoIuUHsgUW6cbbM0QJ1JpsA0
Qqx4dDtuc/INzq3wpxVkNYuUlpjgrzybczHaa2lSgnaBZvedAODxCwzuHYPAoiBqco/RBV/8WgIo
iMbJuLFV0eHTK3cG5UKG8px8i+bkhnK5LXQkCaTWJx1wvG35bP4+C/1IXmLCNt70nkniqksJ7+eI
9miVy5UimCEoUPY8OhDWgTEC1ay3ahRLk53UPWTrRAAXQYYLmc4tS09G9RHjDK6oa5ae/SDUaM5X
O//X0Um4d9YcBRB3d7hhS27wynx6dRtsbX15112rK3c8ltpNg/2S9yGRsJO/nwd0yK8+/r6ptK3O
/ViDC2heTKDeAHY2SaIBcAYVUHelrE/YoaxpuH+G6GneiBguFeoA69LRWjGHLR3uVNOREOaaLiSj
djl64HoiPfDCMHgv2Men/9rHi1Xts42cMW4Rj/kGKUw6ZJGVs+oO4nZfjTAMDuETTwuMS36lCV5C
hdJlxvNRcSmDX+Vu77MS5L7hgJtNf5wCqKy21RjD1PVQG5SYFyex0C20+2QJ4tFuyd56QNNu+glH
zk5IC/eclCF7plfRMoy504j82jmyt8b4wyrK+RyF+o8ZmtLxaZKVR/CLQN3XD6MtZzBiHwTGd86D
07vOq5j4IP5Vy9o70KmLbSyLbrPQglqeWRjnfcouM2cyBXmAuwQ++GgsMANKDoIWNo1qJKOQYZQs
nemwD/X2uLiynerrB/xejGDhl4kCudP7y96dLboJnl1i3CJo0HTVDgQXXaXvnAnTq3aTOmdQHbZq
/cQb06hs08xNWkC8MqwxPp8pIPOfavzuLCgLYvFT6Z4MuytCIRqbzbvAd85SKtuBEsyRnUrRWR5Z
3kP45fl39mlPl3alJFRVP1j/AbRi127BotcFXCSbEMXjA5Wf9Ze/iWdz7GUcCiRvtlMs04kh7f0r
5PQXFdWx4TMSQ3Q4Bp6Xggwl4CfGQMzhYA0fxx91cvvpCApk3tRflCdWYbiNDJDcmf5X+4sMHe2k
rXb5+RGqqr27elfQmnjFMBbLqGsdrARB+96248EFGYs4LAwmcid9IvcVpzZ8vjJgYQYGh5qd5ypV
Wv1irAkjIGqxJpAkYDKYRHeNCei/thFQFZric9Q12d2X+/aQuZhwroyTo4aLTiouKfuewtxeZ09U
ygS4O9NB1XXc3pZiT1YWMYhTTUBz0UobYVQMr6ls0xNgN5FNuoCaM6l+JhpZUJ8M5LTD06Jrre1P
nU/78STMVpPb9x4tCUIqyhR8rAylnsbRYyLyPbpJ4x5B1b1EcTc+drG36miSmVORUsTUq1KhenHU
ZR4SwI2jSl3t92eQP6JEjPTYClnFWqDe6UZKdcHXGpwGqzWvzLWbiPTGrKr9nksjwplSNK9DBEX4
CN99jTNAa+pMIBRrW9Es7Ri6R+g+M+JmvzZsbV/q7IzyTh4AxtRRH4eYeaJPGFgxIpV6BfDgk2pZ
WywnrJ1kk94FF5x+U7FZ82TvcktMWu+0wu7mEhD+bnz8f9USYVKcKikJ/xAQGOSXISKtNYWF1bI4
/MkK2nYBZFEQiWfswY9Hxdt6Xo2eFGFOWCE76U95BpSyBZDIhG0Q85Ycl+KchGoLpjLPsERWMUYW
Kan9X6kplKFz3wVXSsFkiG3EJgxyx+kLBOtBeVDcO6HpHaz3adbbOJHc187FLzTdtj1m8qofXZIg
8uYy1t8wyAjy8VRW+4XDPPy7OHIAfdb6T8FcPnHHpi4O7txnjggEvrKjBVOK53dzqbAgYlyO81kJ
xx8QjvNsgPne2lW0QMG1OD+SWEp2XtVRsGeBn/Qn5m/OeahbK2vlJ+AdOsLj2lVgVoBDeQnmcYzp
0Yo6gJ21npj0QXqxt/TSSJ4L3XUQg0jbb48G6iJJE3czn/AS/RG5QsldcN+QEYtLWG4eHEBQvUsB
0w3xKI9xQ4Wga+nIfifsjc0bbXrF98jW4GM/1FzCUrKBOBv3ge74Q67jzy3UYyKage9sbKRu5sfZ
81h0Xp602LJjPl0uECCYBvH+1g19rEym2tr4CX154hXspaEHNNldkzpsw0GMWkh9nTtpz3+e/9XD
FgO/rA1eVrwxSub+FmBDYCNrHQh/2e3BgNGsmEIz1AKDghDViaDxTWMb/uYpvJmbsku51IxQJAks
A8UfneYTAiI1CsPdnr14bqqOTXHzFG7qGZEM9FYMsyOiD163IezcPsB4Zjrut4M3ahIiOPB9rxLz
i7KCueud1HaCmMti1B3aVOMvY1R6VqpKbFBrDNGYs4P8Y5fvIx4/3AQd+ESnKfcImak956hHbOzK
3xlQDwoHi5VKFeLTbZ07z+b5bAAXquU+bm1ZaVLFPoe6z+BlaJXT7rgi79Fs0Jl+539pZRcvYkCn
jat6Ir1YW5WEjKk9JbrSLu1vkrrp8lPT0HUyaYLjswFBn9cYqLDlqmllqi6VydmGMX/n7Olj9wwK
fEZVxirJKiGWyVu6uaIN+DUxmzXF1w0b41L+ZZZhjnz9Z8ZQKXjtXh6d57zx40+eY1DBbstmb3UE
MK5L+gcJJ4nw+IOfoTFiDNJRn6aqmfR08mnZkOFkCjd0opaswIbZ8jm5jTC15KQhvEfsiVZvLu/C
fwko6hV0L4tcvQyQO19+7WCCJsje4kpQsxofv11ndyHzZ1ANqe1J6rBH5W4U71j4iGDJxTfQyc4B
TXH1WnUXajUp6/I3LVna7vhzhtqmh5n/NIwQIwE4esZNLlYSSeLqFIb9v28f/qjHBUUgKMwMR84p
lL2z6VXmuqXHVEtCuiSoRDiHy2A6OxFQhDZzWiC84ygTKk/rKROdlLd/cmSBVs0dbySigX5eLK5L
myxY3+44ERr+Bt4kU36pfNQKo3gVZBHQP/WG/nyKe6VWOIsxQqN+ViBt3ZTz37CtZu0ueer8kBBV
PVbXb69m6B0hwvsgOLLt30AsgCEwtTws64Z95fPhEG9BIuvv/402RgUvUsgh6EhapgmoS+4zLrTT
w0DI52kPsOqalEpI9E2xjuL7KvF5Lu9I3XSFEvpXbx91N6kJ1rjuy1cobSNDCmlpfX9JSa+usrbz
LTrvAnES6Qk6Z2qi6Q2wSul6xAZrISc+gwnRBdFkcGFOs3g6kvyxdkx3vi6UwEJdI/uimtuZdNpE
ZRDJWOFs1wp1R6hloKa0QLPQu9ybdqI92oq5IpjwasvkcNJmXfaOadGEaAtkh8X7m6wbpg+wh9Qu
6r525TWjW0k/omQRnfdv+56iF3ZAaeAwBUYq8GIH6etS5KkTXQE0euwLyOuQhFJP/lhsClXqKJTJ
jEqBcwmTN7Q/y/AM3lAsvzv3ifFuaVDA+g+B6XxqtiKaxSAJmwQtRbSb76AMFuCRIXIogdMgtyda
mrLkGgldKJAOeFZxGsrBFFgifFfiZU69Iv5RlsFOd0YTCEV7tB7WwpenV+tmqsGq2aeiUoavJx4T
Qj0+50xv0MXb6X3djB+nZeNW7oN7JSF5EXrLuYCDM0Tybm6QHxYV2K9QBlO1yaqNUyNiLRPxh0TV
h04zvh843j4TBdwmlFuC5yUztcu9dR9aPL6Uxnl0yCQgIjaSl2ZJ3isylLeKxMApJUujcXjBYZxm
/eY1eoo93Ng1HIyQWsM5+F/qREqqw3T0gMtW1Ps5mwApj7vxy4RkR1Fz1eW8kmEY+vaaf8fsQHZL
xbwF7yeQdiH+RhWqDgEvPCkAbOUq7mpw5Cp5g+vKwYoY30Lp/Xt6MYBwKbLb/JiYPkEAWyMwxO7A
h/TmQFaSa0rvwGiM/sHgG5grEE5X3RBeMazNh9RuDudwjXPRjevc2bTGxBuHRLZsUcRYzxCqzQ4T
7LdOXCw5QAbFqyVtB0d49dJ9yEo5962XkRtLL6NVTAUt6uOHwoMjMEdyyhvqFYBxrorMIsjFPIcB
iaMnmG9+FG8RWIUGLX7ZlTIm07GdoFCkcvNf3YgI5IoF+yu0tAUveuTcAaMVjqLInzfCR6zeZgW2
TgnzyqtNUO2OkyFTJA2N2RnTDIFyU68xXKYKxDJixXFZt2/bsgIODQJEDbHcOKCVfaL8utM83yY9
lZtrDtZ7evDGBvhodMm80RYc03JHccoOQErP0d9NFiy7sTnlK0NQdDWWQv+z7TUgMxOSrgMxQ00X
R5L1MuVvtoiNcEGW0oGDIrnFv1H6IUOctrONztw6jLiOj4JAM7ERwKZeioRyRPbT6L0hMq3goq1k
Ga2KbvCA9pr9lsImCservxa39upJuhC0ZiZNBdXqZlY8GcQjVY00fLhjrqkd8XX3tJcUWLZUMxje
pj3BGlfhmfQz+vKxTkWdrzphGQdU7qsJca0iUZ7pVYj20tgjmh+yPPQMosy76wgoV2lAAYwbtPAt
dGSEjsXrgHLeVj6+u0q3PyVprMo5JihONAfZ6ThvfeAq1dcL/uxObJ15NkiPP9jQLBH1Q0I2PROS
r7w/vhN3X/bB6WRyqeOGV5dm4X8oR1NcaUJ7t3kn1o2Uf9xYUhr3apnlGXViNYNYZQoROP/n7gNN
F9n04pN96B/AU7jJAyTGIOm+M87TVkdoMwtnNgqgNHpNymDhqWH3nQA8fOy7lJ6fDevPuGBtWQ1h
GHQknK4FEbK2KV4Nbn4ZYrJG4ieINFrbmUTwKlaIFZvJLtN0hTtFgxg7XCSp9aY9F0/um3uLQrpL
nGMDE6ZaSFQxc23969K+grHHFPQs+UQvuEh0JJ16mORdxav2kmWgy3lWjjOuyFD1tonNJilpq8Ne
qI+pO5olpIpJdY/18qXfkaxBn9H3NK4KDNq3fBGHtvxIG4zWc1uey5z1wl+JvsLxNT5bAeWdwWT7
tf9Wt9CSLea+V1rmY8sibjac+o341TxQX0j+REtRkAmRoyiG7EAtQOShKtT1NYyl7ge41HnqcC2l
MCBN85E6wdMSevlt4YUM53K/QK26QCJyx+ZPtVtLbPktoDLZky+BCR5/GhNwpgjFiW1X+/h92ncQ
mhXDQ7FdoKvlY4rEwu+ngTfJa7SujoeulBHlkXC45Y409v/beswf2WdM/YNCYflJeXZcxE3A5NZI
OuqJ45gY93ZEgmxnU9OLCcEYJYQlpwY4jtXFV64e9Vu5YUCPpo+tLGvuKxF8atrM95ED3VQfZCuA
HV43xaKWPnZDFwwJ4aKyLddELi9BXH1vXvAr9AFaP4d0zpGKnzWnajIO/n2BcscCtovxHruwtYki
eog+6VWzFHDZELWiPn4tKEGqednwZpuU4O6NpNY89DGAtqjV+NEMVfy3P532kg0TS6sK/SaP+vQ7
eT+3wgEQ7rKdEcZg04ZsDkOtHCV6olESEFaCffRYxrdf2ZuR/c7l1BQggITuecMYw0qemtn5agFS
7og9G7HYD8E8NKld3zlkxs/mKc1q6Lm0SHuOEZKy9TE4g/nVUF514PJYhW4/mK2em3xMQoT+KU8b
lLv9DQi9PUt2s4zqxR3nGXri1obe12LuEHGfUnrK5dXi1nB2JCbdjPC2BSmx4wjLt0S7R019JSVs
+VguLD7n/dZEXZHB4LHWm4TWFk77AG+Nf9O1HzX96IrwSIUVRoMbFqjGa8HmeunzSFOBjFbHMWBD
onIMMTMaxjI3B9mOdqVCDqI8iYCOK9KooBESghxE9OqzY2GnbuVeEoc9409JHOih9OCZ0p3N0hyS
GMjToKGZQ5rygASXpFl1SqEbw5MzaUUMivc1ILC96uY9mGN3fTQp/B7O3itOOpbGaCRXRnBjUrub
tCzJFzAi12429jkV/St+hL3S7mRnc/1gqsQZCn4TkBuEYGsHTghQlPFTNQxbglyMR1gHoviyLTJN
buGX4+31AiBoXqmg3hc02W5PcASdsedIPo8ewbVdIhT6m01/N32U+hP48YBQJ1UOkzuSP2Rdlc9R
ksWOLTJzR0AGwT8zk368ZZjn5zNSfWD4IDGSDSi+DVwz/njbsAf3tyWKMS4dfZCZIoyJw3Va7MnW
HO0sqiS8wqF0CxDev8graWS+kXMIXHVd9bMrngOWIgnAj8tYGwMdkVceqctTWygAh3ymxvqLyjvF
33KVyszh/iiUx1+OqkZXUCbGD1tkmA1UI5enazPHj7IguAtuFMxMwq2PPhqtFIX2QbHmsojRbnDt
QijpYwCdHYElsG2CjdKmNYdF3Stf/Usv3hCx7PzkeL7y3gFM2WGybwl8rVc/C+vcfkA42WsA3V/J
6bWS7siw4tVI+5OoKsDNqWQ5HVtE8mc/Z8PgLDP2WFmSGg9xq7VyLUe3eDD5XttatOdpkkZmL62f
dB7gaY4rR+wBSYhvhjyjpZUnZhMD7n3NgfZKbbIVm6Pa3mNh9iz1LEyUkBQx0xEbAwABlcqsh+03
/JmFQDvvkUxC3bpSYWkwZSEQcBEgHImaGOsP4fNbUUYlwhAqsJzyQSN3kJNsEKuklcUV1YB8ukOv
DEGFUFLtB278SaanxyQO9LHEUGKwSYmIWE89u5r37x7Bh9RyBBTylq9JKngL9zEeqk+z0MKK4Qkn
Y09hb4a0ulYxX/8Rs2QdI+Q1Y4oB9TzNZBkkX0BtbBOhuDSmRM8k1KXTmifbczx6h4DcZHE4Q50m
Q+KqAjdBK0ofqNXvaM3fAVYCAyt6p7WbZVrUDf1qhgX0BHzlBVm0ckrDB+eSg1n3UmzSJ7/Jd3MZ
7S7xghsbxOGpL/kC/0RW0YTTX5Rhy3D5KGBJLcN080dpgwLgs0jKtxism2yhvUBS/wxNrP7aJ/UR
IrhI7T6fvQA3HS97NYjLeb861ucjtueG/5Q4tgqVaokhwl0bpCRDPdffVz907eHKEVKwehFqXUee
NeIkAVix57+jvxpwEjDC1JJ2JheN720/5Enuz5oTi/ZnuCDYh/DQSUulX3YxHGyQY+rVn9Lebnfd
+7wJVNaKdlA17NKzNmXLvVPkPfNcIntZiHFNlsqa9vQSJv1rWFqGVjfUQ12VkWMg14y5OXdUFQld
bv5vPAYLQ/e5zGcDqKGsfEe56x+4MkQneiByWPCeFoH71gXQEluVYfwtXZj1t5xLdDmG1Qxnj+3V
gQ11xEzrYmeZcSPhSIij3tWShAahZo3s1PqvA/S1lXAy0xPKzrAwC2D2t/AzkB8TEOs4XB08Gy7N
d/WVK8pxkFgSCMgIoIfK5snCy+lbeBiWUIA8dTlyvKGCPd5YrPonGAEISUG7BZQgonkDS6zzswlm
I1KEB0++QGGqufEK5rNiW9UhNNPUpERVwngdxZwxKAHhrvlLWb5BaKdKWPXgxckBsHIOGNErEKDG
7HPMN9Du7yXY4U9ZyFRiBd9ZHJMiKOTF2hjD2BzqrMO2OeQr9ief1GIJSevMhYiw2hwFBgNerBBS
+sknDZtnOwf0MMLdgjxmHOEaAg0B2y1luQmG+2lI0JSToXIdE15sIACmmFhalWjmjLEI0w7yMNT1
MU1yEIg6ZBg0+bctm4DzPbXcjtA4doNGuLs3GtvjFm29hP/n/7x3N69/QhQ01v6X//fnyrCQmG93
qqIeKI6pDJ1UR/rQZE23RjRAulxjtyHF030yNo8aXWODCisy4BoBf/nB5JxUdo0EKxvmft0kMPVv
C4iGmNhzB8B70YQmlkq52sTaJq/Q2dIJ9Rp0sq6OtYmLJ+9t0dflSiE781YsNUL8F8D8LpmoXH/Z
pQzlJa8/pXp3L1HdgNRigWsswTk05+iyVSo0oUdQPDBBcDThEs3U3UTzdLd4GeoWfoC5rXLMvpTh
uUo8XGEu5OkNuJ1vvKR6PEZtQbL0+ph1PTTGEeNE/QmubLCXoabfIPc1jXarAAte5NzDKEcuNR4e
YPF8Q8/5vM+Th1uZgqJG/sHFt29N3EDu4D0AAYDq5I0/PipRVCWKc6PpEluW34JBYe9PGJump8jr
HTMoB8Nt65AigKm5/+al3LX9GbSJo93s1r8XcLVbv0oqloaVdYWiR4Jba4CL5FvRAbebCWPmc6hu
Q11RZRJBAO3m8M+xXmnCjXAspMayHoVuyfKKkx9S9QY+5KZo77UxgneD27u+S4to7C8Sb9Ckek8/
zSpERmEvBxABP2HsTw75UGDuFldrztsbN8yPn2JAsI81CaEOPCD2mz6WtoVsmaNCmFTpXsOMG15b
WTkrJuIhHC2KKf2GmwIMfPL7PfykwRAK06ohHjQn5gkr+JY8aLZyMRFAKHLLecLtI7tvVWGNK0/D
hYr1f/+u0lrZnCPDaPvol+dMg3vy7efabvegipNjEyhF3gB+DQ4qJh5lNCqtNs+YYUUFCnTrMI2/
Oc9APkAy4nbWO36B2YPxBvWowJGzRRIeBhwT8LUiKD+kKSQYa/qFYySB5TTBCdwVZEBQcxDa3raS
TTmjeBWajtgWUZM3vyUgpCadidamuBq+A6hdkIr7WDEZ2gF4STgQ30O784C+lmxR4b1wwKAPh2d5
32NiVA9sVPsgvskHzX4V7ybvK4gO8QfgkiQU9mhBP+rQTuQGvXfq46IjoZUbKNg1+5HOFUgUEEYe
ie/dL7d8IWgddo2tR+MU6OmCf60YksYAMYc/GFujtby86kLAqxQ4/Ryt5y48o1tp5Q57TXU9gYur
Sv9KpicW1f1wz0Iy5HC/vuipmZqffvliAC7O+3Y9rREu1xorwDraoQuOq21n/EqiKAObz8gmm2wo
QsRJWUyvo8P3avQgeD9mAFHoHU+cAETB6NrARHpL3JBPEn66kiA/jlvbtdw/IX8JbDHiqAvQbPl5
tbistQ6MBN6WbTc4Xpnv5zKrwsWR08wIq7UKdYxdNHOg/aVUJRpn9q62T2A5eg/x7cRPgrA+0SUe
bWJljT97JJGr9Ycy/q2f86iO0W6y+LdBi9gx15PcdnQp19ruAwBLAY+62QL2FhzygM41YvjNN+Uu
Iv/ixKphvDeqNp4VZPGZ22Exzt1ZPn4zIZyT92F/6OBFR0w9s5Xq0b165cpMIyuWChWU/3qv4V4r
737xCd7YkQstcdjEZk5Izn7d4pfx480JTNKHlKyzHAaz+AH5dkci/31AjRSdcgzHpIYcJ3S4fF8J
MrdWqzW3xhsRifQHNR+J/9Oq2Ic2uTsJ6aBSj5MjHQquuzds2sfu0c8C+l685Qf3PKqb8j1Ahn9w
2UM5FhZVHd4UwJaKvIQR1YqxUrr20Yk83qQGLp4ccaEN4UDKYH80EQv4vwNe31e49MQZ2FcN4pF2
ZaBTi8wwt/xxlWtRa4NBmB+m9yNrsnSfBP6HbAQcyu52IXx4mNoRjIKM6h3w5VKAJZP8HjourdAW
zH/HtoDZ6Ua+8X7Pg9eFsnU8udUDaNtokbBh8rDY95m6aF2FnQHqYY5j8jXsDsunbON0VTDW5oDt
/olionTzeZ9mmKXXCPxdproaNB/k0yE1MdlrPCXXOOv0g5UPyjslou98cDqpFJPgcnwdMBHgR9fu
qH7zLy3N8nh552I2ODmH6w5Ls0eNATxJPSGNK6yMSUNSDts3QeEsnB1lHdXFX+7igWFE0IrJxFkK
lf96Y9f6RwAJdC/q563bM55lmWrwEmoh9iC1Reoh36SjL8t544C25Wgo6jszc5YyiLdLcWi13O7O
eU0s6xVdH4RFUZD5M5/QHTgOsCi1jhC2J4lK9uF2oplMjqZybAo2JKmsl9ZmIgcxkI5tJLm1nELh
SUGGUi5Cu9fzVA983MVGG+TRmD0pNUo/Ls6oIFiOXHifI1pt+ugbLDxJEYVj0x0IHnxLUX3uECfS
WvcgVQ0Y4l5vxiHD/MvoKwero0iHGKAjwpSAZ22qFFfa35HdixXUa4xL8xKoHftJIJV0Da0BZk++
kKpeqg11UkldneCNbjYw1n0P/1dbwGcGSt7Za7irDeHqqYv/RWyMxHDeEyUMchUoDFw8hV79LSDU
1u6sknDzBioEYU9pRVCQTDykd2IyqafPtko4R3cK4C7V8+UhG3iE0olqlBiXHyzSQQr5MlQpYG2r
UJUATAEEST9XIZPU/V1oJ+R5aB3H9AHjUNT1n0yQZJF3k9Uxz8Xgk9FTzsc8y4XW2UHeXYPHU/fa
ZSzlK27Vx4qGAWrSVkD1+FpJTSdD7ypcIJk5ZjSimloidsz+ewoABFmyFG/+YmoXLe0YkSPLZigc
JipNxvq5bm4EohP8TBCJdoLDaWviu003msis7v1H3rSvdYXOgdU/zy+UmE7sv2Q+VzeTz3VMt1YT
xPKHs4jo6wYB6DPRHnwuoQIm9+aiAhgBg/+3JTYVfEg6LODXKSJgJ2IlGWlXmIKbYtavSgL0HeZB
pucdUG0TlmjEpBzAq3pvzMaqHKSUyGYkMQOqNxyAJADxfUsrqvXDsooOZMN5td2nXXCW2LA7820j
KkrQVgxZoNN2ENQ4LESMiuXFiXnMeGfh8Ut1l3EOXBOeCC/dl50Hxc9SNBYenKrwS8+A6u6zGoE1
Jxn9rHg9pa6Pv1SNBvZCvkn7heFp0uRx521zjqNhmOayMDziDdZoNv9uW7m8wMQuODArSpkjPzBM
1107KOYUf11kmvV4yQbn58HVxc55pekXsPnT1e8CMGZFIVhAOeKGoAggN2ORPFIpUpZYiHyyUg4u
JWEL28y8FUVwaKLwcXnNp4asVY/a3N294UPJIvYlLBb3Dy3c6GgcVENeZScRSeX7AeFzW9cLeUCU
BEYFDOZ061loflBcDNbfZSY4FwqgKUZ/hjejmcT0YSdhgcw7NuVtdlYLHya904BCkFY4Gmg+196D
Dvxlz9yPJ6dw0o5BB/LXlGLum/BiW+7uONDFCEwaZ+9qpIbLgeRqMfWvVGV+QiB7ew98LHKXKH+A
vHQ8Vo4Elx9ovnArCfVqALsZFb7R9S5jzYjtUONPz5YnhLEJL8iM4hlfB4ry6lt4PmnO5LlZ3zoY
zpkXy1AcOyozuperSFhA9vgfnwX8CPu4jnYVvtNXWypD7HpLf3Izvqceh2bvXZdjSQjpyEsaH7fX
3297IPP2XQwezyRi/kMNbxGmzeOAlJtUR3s99ODI38kRLyPhbSMecvknfOXS226chTYbRodfhI7D
FJ3PYi/KF4zf2kGM/L/09LBa1Rp7OfdFmt6Qs4UQ1TBPaPQ3FYcSqMYfddahN/fK1vCiihLO4R85
dSNQk6ziKupr7TrVO0qWIxqXPb6mJwq0yENDdW8pSgJN9EG/OLvVHmQJjzOOiPMZAcfm0s2GOX/s
c3RfwEwC7R+GdxFSlt/Z0DJp6+z6niq5Tvu/j90pg+758B/jL9PLdSNFHnMlHoF8ak/4wHe4ojec
6tcW6UtMrmZicQKH14bv9dSM4SoSwsZqxWg88AdSqNW3w+e6rFXVzGpUUGG4BFnHcwrNuBA3suqa
MqtdKHS57Ic6EbDGb6hYyhuQ5hYuTLllx8+IE9AF7r/XbIvn5K9cFQU97XAkQEF4/7YKPnE4AXhX
iSrBcGzeGRTNulySPAOhEjhA/ypt7FK56gi0MZ+Tbwv2EKFnUKrryLQFpXiPwKV+k8snoQFPuwuI
r4xQ1UoC2iWXhZBun/ANHeknu5dwkVoVraaD/nemmymDK44An6phPRw/mbBeaZdfqTZi68oVPBud
u37S3q7Ik5BZ4iFTuR3HWP6YqbCSyGE9CgKvNFytLf6Rwb33v1gVUJyPEobgo7i4HyD9L8AB4OFj
ujugKn2rMOoZl+ei6LZCYPuEOOa4EBfmM1/sdi5nivqoc0iQBTHhswj2n4GCqxPN5J8hQbYiYFHG
Y/6qJQFAp0+Xc1ridsCb8QihPSoaFt2r6eTrYLpu0dU/NUtQ+Q69YeLrA44V+BTFdx0Kk7C5grIp
OYUtucnWBHMvM+VKTnlwhHCYrcVnQI+JUKw8wVLkHy51v1kqpXwQEj/Ed/EI3OYu4bA/+QmjWT3B
/nd+tmys6eWXZMMQBr9Tdfo9PFk2rnXMg508GcXw4FY6DF4VSeGkm3GVUKXWJwEsb38JSvHUpn3h
wRsrQcHCxhQo9qlUzH6tVdT8cEJ8KQp8r0RfwTXLXKq2wjbtwW6+jdvrEkmEFgqgdPluFFXzS9e3
cuQIBRl2GngMfZNYkCLRFHcdS2AGRQBqJrbbTtZ9T554WSePagyQSmwos9dV0ZFZ19U0QfS0J2VU
J8/UmsK8FjlHTPLXcYuwAvrt0mt5Iy04nPUAgiZGHR0Z60mvtZInd4Ze/9Ued+ggOCc7gvl1Bggh
JA2PP3jQBzPPlkgLc7BuIKxMYN16AH7sOG5uGFOfrpWP2msGi5Vr8puHhS/rPJEw5hilt3ojvQha
1eX1hWxUIfDzdHn6djczQclej58Y6eunllWyHepaPlD4UeJLl+/tqTiWFGbEvfje+pEtnd+c9r3t
9p5ExlTx2cr6dI9ksgxJw9ucBuVhHtAhiLujLfy6Q8wNobpkGhEqa/dsZ5PcNkG57XtHx0M3xTyB
ugy07gA35wtb60jhDlF0LhsHfUw6GPvd7nUg5IDp1mwUE/QgOZ/uV5JSU/+Q9L4YTywzU2/4Y4G7
mwx1w9nwpLYacBIhG3ubcDL5YzYVa27+OmKQ0Vl4OB4uMtExbzjNw3qWDzYMGutnjrftbevtM8rS
8hGHz/akN2maD4wCRF/YkALn5SgyzGrKSSlhxPsSJTdBPjZhAq0+4zEKqsHoHr6hqtsgDh1dniv5
6regEz5K52UvLkO9N2YauEmR2jmsLCERHcAzr7x+FJrI+Xz4ggRzmPQOExFnpS62Z849HK3QTdPv
/2snAfsm1TEcK6ZpAxgziOKz6iZihj4+4thXK8cNNzugwwKtN+kMN7CDbIkL4cWnLw8HA/KE9gF1
mzRqQMmAjb7uc+2VjSw+JyO2DAHrp8gsWeQhFqxR7XeygPoYv3ed0w3BvWSdIvn7PKqLGdr7hxQY
XU8p1byZH7D1GuoEniYIfulHuxUWdGdgH8P994S5rTBdUBCD3u8G0MtCoZahUa0DKJM9RJaTydyb
ENqXqontFlMK9O/6/hMbPnH5FWCFIzsTcv9MrHQFYex5rbGV9WE6Et8Qjrq6Rgrj+4SEkwaiiE9Z
BjK23iYmXDttvMoxIxem+bQtKK/7h4Mj0rcRYEiC8GTbwV/WpCiz5t0aeDclyOmfa87z1NX/9U1C
uXgiwKZD0spgf5X9+bWLC5YaLnQ8kj2+N0/lBX2G+gZsUTT6P5oR+UQCpiOw7C/oXyDeTj2SXGGt
AXtjT9ijupl4hB89sydmPO21UvXS7E8/F9DriHEqLqRqzeCVqIdLrad7JkpoHOK0W7/CIN3PPcvW
VL1Nex99aLCXedjm2MwlDMjsof13vGX03ATIeZUiD8XKY5Qb1+awt3K2pZMU2Fm/kZMgDdRf5q0O
jWjp+KURAlif5oe8gy0HHcFUojoNvt6aRjwUzsBnSxkLfpV1RSXSXRi29ToIYS1+MgnZ/xlQOy7k
VlcPHjQDVaIN/GU+3S+14rjm/Oxvu+TQKriAYhgx1sSBpTq7+2ctd0/wTNIaNUaHdFObO9g6qlmy
B8KDIjcxRMnFRXYBifsa29EurSec2nG5JvJdlYC0Xwnwko4GeZYvjRZXP8ekTw5f+cWN2zml1MoQ
7qx+yV+njS2ZMKaexfd8bkowhUWdQmyzoK2S37FXo6WzcX3DWc8ja6j+3v11pM2xSyg+tp2HG5Vf
iKYr8vFCUDwh09elsuX5NFljid5jdR2XJI6yKT5QEcq4Xmh/y+Wo731zgiQJN+VYExqkkN8etnNI
JrT+aVrrWzcEbR4A5K76h8e/pyf/jovPFmaGK0RM94MtYk3waCLv2t28P7j2nH4v25C7quwdcNS1
9jPryIHUKK6BUwifXUzHbz2Fs4abXGYtJXhdy3YOAmh1WBeCBuIRSrUPGvlW/hJK3odXDmr+ZifN
9JAS42BA1sWEuq0GoO95PfbfOau4xRDnjBCKv5AR45ymHlIltWT0DIdbHOoJrWLYLsD3CV3eHwC5
Vo+6PZBqchQ6Kjyod+HX/Ig3B3ip+J/Su2+cCzjrhyDgcVMlmq6mtaJ4tKLdO8RNbNl6V10iMpZ3
PwOLwROvbig22LJy2bVEkt1E+W4PPWeeTQ3eJ73R9zPCCqOVzhoHAU8J91+xi7f0OMWYiY2mAzB2
ZR8GUbZrsFYCVRA99e2oReh21ijWGTC+hIDppegEmfo6114HIaSWijtwun+RpRrHrPpN465Y+wRv
iSux7oHEFZKLuz2TfrF3ro1HOOEBnuhc5QLL+VRDd+7n4IPXiU9d65b47IvmrMJ2e1IfoJtqa1wh
pCXIWRCvZNquVn2tMZ3Ocd3ExYmi0dAHIFkAZ7CYBBO0B9Sp19HoF+NjWN52Rk2wLUlZd1CKuvZ3
aP8wcDehiNPzvHBkPjIPgBd8RtWLbWHTi4j6gc1di2cAvUNS1i/pUhBDv9H7IpK2yyJO4USYtkqo
r70JU003dwQz5YdGgpVF6BUlpurHBr+0Rtb/Sb++h9fE81xo4pRvmLKKilb+mxpYcQiRjFwznqiR
C1KvyzmKrKTUDynz42q4ITA9X87+B/uUrsTTudNt9qxmzQdlBv4M+RNSxm1sVmyCpnY2PLQcLlgQ
jsweDIcEyIpDM7NB+EB4C4jI5o6S0a5DTgj5ifCmEz3KpatiHyI2ePY3/2CuqsLmXHlRjQ1Ya5ms
nLbTjryzpD1onfRAlN1DDpB7U/JucJ/saX0RD8+HSd2GOEOd4qcEh3oxlivncABe+PynPqdR/HR9
o6wvNTrU7SaWH3/1kjpQLl8KicAxjopkF4hkQqlrv1cnMzMVX2/Fhljta63FZsR9rQtNmF/+FL8u
C/OXuhJGsRoRq+xbvkzom6NMGQ3tjLI2HvdNJ9N6dyZg5DFdoFslsjwotOilBu2S2FbQLkctHHDS
6gdGm6Qf18j7BxmUznFEisI19Sar7+4kFxhhAlStS8KCG1xkVNeeNsne9Am9L8bZevElU497E9/q
DDGDslEiu4GEyKTvzbteNtGJfgUSFYHR4fI5izuNraxhEMn7OS/GekRqSlp/rr1sqh28Rt2EzYJg
f2xseg1LWM1VoOPvas+wFLYLBUKyHH5hYWbPV6aeISwQp2Q87uWSe7e1zLtik5LUMtlFRUub0AX8
gC0aAlWl9MDLLGDLa7hA7oMElgOoPc99O4CX2KYzSxryGhuZRWBpG5OhgbPpX2iscjJ12tKy4Hdc
bejn2ZT/mxHfCXVJ4SkpFZR7VvWqSWPomFRrDCHWiUhWiqDWkEocWpKyYTKiBMDZBil51g0KbIqE
8LuA0A0kzJSmdvNCaAjbt3lgRsrOAX4nfve4UoE/lNXmuZKqwDVbgNyDODzob+Jyq+DE5vWLWI84
P90wI0bJrph7u989vP4QpSXZ6MY/U1lBNNLozIsGm1WP2/DiDaE6LaFWBucsLzcZzOdbqy/dNwYx
zoWA/8yUt4SWFgD8B7YICfqZYvzBupXQSo4thBc2ytZTNl0luOQBNlGmRqdO1/wEsXC3XMs9vxD3
jnJrtEnpER2e3QnoNpPzEihAViN3OcadY9gR4cIYlTTNvMv+esEjg/gGuzF5YUUEDIke0oxtN5dV
EzJUGVNQvi05ItAcbKtUFAay9UESaLhC6qMwHxJGsyUxcbW0zJY40P0z56fBoBt9kFTvX11PpXNb
/C6DzY11VrCzazzQAr5nZnesa7ap0sUzX+/HrY9M2GlTgEtEnHsyUqR/KIE/Mmqps13kSlWgithZ
wsnsljEP26AKvxFAkR7kRgfikEZrMINYRNm5hn3oQO1LhsEbnODYCkxhUw/X11OMjsxJGMXmabHw
U4RgrapwaYD7VY8EBxX3xrwdp4HCJW+2Ea+O5sb26hmLuF3n4Ho06duXZ0S+9ZH/BwUwAqfJ/70G
3L7N7ZAiazPLnjT5sMC8n1NVRpGbASGzzR0RkLAyTCtnQYc3mNrpaaoE66MfwMRQNc/61AFJGVMm
SjlDcF3KbQphz/bgapndBJWPOJ/cQ7HeFQL68g9WRxRGBIXzxM7xnDx1Xw157AtA8S6FQkByJ9J6
8EfDWZz4QVmV3nWCC4GY+L9XMleRefaeK7fICG9Pvco9jWFC+t8GXlEepeyJ2QvPRywtvkniV5kV
rBe4drE2E6OuhMPOuCTiWVD9Lp9JIL5M8zD0SpJuFvbJpC68JGOUCdcgUZEkdVNA/v6nFl0KgbRz
TDozCdaj3M6+QjIVbjNzzaRfVOBugb3pu78bTM7JkjOixklhEpezE143GIY75cJRlo9gwrVAR9h+
C5qVS8kUGJNWenzqvyOO1aTblzcQes5lr+E7365Ks5f95R6WblKOz7GHyjjjHZyxQxRoUhK+0/vQ
Zm53jHfszn7HgdN4YNjgc8dAnsHyW/WPKds8u6T9BB9WzMLyf8FhIgWaPZZc6NqoMz62l13btS9U
uWkmq9DOM4qRaxJnYhkEkuh3puUaaBvzPM1KKyUVOsFZvDWIaGoqwjLB2yyb3IlgJrdK1Lt7uUHw
9xXRCeVnuPbImojrZf/nIKqdWg3/PEaYCjPXhhdGsrt40cqxMQHGhoOFthpEMCJgA2988UEiJk5s
a0ivEw+nS3J5K65X5iYlFFEiugo3bwr7LBTdktGW/oFfDdhAkzxfVOr3qtMR64SDJk2YyI7GLMUS
qtlRwQ+cOKgZvFIntW2PXeWy+qBd81g29c/SCS8+BrAwIFaTntbJfSHWcNKeYFuXlE9UXqLuBX5O
kqiXOanm1KhPQ0xkUgtYu4SIXbJiL6l4PcAY8rVEAt1WNYy7G42Vbz6HONM+DWWBAGvCz12PaReJ
p+DItuFZlhdBJ1HckFll8S5I4nYwK3LMq0LQw6D3m8YGrf6dSkLiOPksfsD75Qe3kl6+t2Y7YLqU
n1pZdTtUxYFgeHkigF3LBBYjGYgIo96Oin1QYdbmoBeChPu6Hz1XsPCgDG88rvxaw6HV8P+asPe0
tEoWEU830BhSsTdZoheCWKpaZCWaMdvBPz05oNlaQstVii1tWO/JCk7KenM/9WIiw6tS+Ix1pbiG
XoU7XLxffP1MlYrDxeRmYhXua+0qN+/1UXIzIqMcsmfV4fWMvN3ZOmKfMZsVbx0H0aWPmp9NPVGy
HzlvpadwZ2puiwVQIq1F3mALvA+LKkxi7McjPBHEBHR5a3rwpGkYTxYfqRC0lcW+3qEl87R+subI
xNBmo/P5YhiPHTWNQt/1xyHwtFyKr3c0IPCjX3P5c9E2FNaZzvN4IApgwrCXYyg6eaAAhPvX71cw
A6QD8PKt14Nm3RGub0it55DRZE4Y8gh2O8Rw6ME3Yvuq6SueiqIYTdEDWnKoiDgD6K3YJYMqsWXa
oJdTBDSMKIimfOBHg0LLCXON2W+CAWlhvvlpbfD9XsVNxPYroqGxy4riIk5I88r2tCUsZy9et5f5
VD0WtVvK91d2uu3A8gvI8wBhkgQU7yik2pOv5oIEOuifIXfHGXZN+73AfCqxEIoPzmZy2IUXMuWQ
ep6PJSsdPkhc5z1zcZt1Ps/4OciytvYyTTv4r2+CsxHXi/IrVGh0m0SJcN5Y+AXMgFH6qNwyuOBg
NWt1/4xZ8zKYBoEZNS1kjxtkHtyld5ciAKpP/EEdnlfKz1j3Txvs5zjXLu07wVuQt7piVB/w1Yk5
w4J2yhi4MJnEP2ATBGWkDO9SMVJbjrx1+V0Ll2xbkbozCzjtf6bCfEaG+VCqEQQeUJu+MSdZ4Upx
t6EsGu8s+e1lohb6DXUZP0td+61AHzmB4St7FkRu0eCS3fZ25S6ZIk/K7zh5Vg4paT7C86v4HJIs
AJyovBhZ7NDy1QQqDcG9DbtQIRaqw4GMHRExwqM5kchJ2SCEYbY8e3R5Em+tnTSA3DSacI9JQJzL
VLxaoLrBUKPv82nTv+YDs2sK5htf7jEO3c+1fv2nQ7M5h+P5F1xt9L9B1Wef1crAC91t00BwmWLX
3Z2iQk8V6Z9k2w/Hdi0+EP5cNiUE+uEdkB1SQ52CdJSTwSM9eINpxHQfHNB7NuRRgZ8ZzNw3J2bK
L3RqALdDCpHLDRC7/NjWy80T3Z/uvf6O0bN3QmC1TzLQlcMPBKqIvDG5W5Fv7VN5gAxBCkNGfPok
lArXZUuy9lR8+It+J1MyR+i47/uFpcHSnCYnIvMPwG0GFIbZ2kIkuH5KdlOVi7te+5xmHpfgMWgr
fLA6XZ5G87PiZ8AQiqxlQWIWxIZOPEujDkNpqHOq860B3WFRx3Ipm0KOvhHjG41uAT3pn8IUh4vj
cfoI2VoAzhij+Lhy3HauLyUFZTJRQb0GtI0XJ6TOCVNdmZca0aYWjK1LHKnqXmRIKsYb2qcvbRBR
YRoZodUMa7ByvdXh1Dr8HOsAhuEnt7SaJgRum1hnOlRcXCVBCTCdIRcPqWdXz3mDyLlqeu5zhTR0
fVLm/0KCHP56u+ycMvEUVgEa/UOpE32cBTBne3kO9K6GYFRhDshYN7RghLM3aCvQNuCg8sBofxvI
nwQW8q5+p/1xBijaO+VEsqIm+wZqcdP/5sTRSS7FUNijS+ybMg7y8wATpPzr6Fq7xAxcfIAYAJ0A
pI5HBEQKI1K41Pl+FgcXVpWviFvvBcfRJQLG0yHwGqD2j9d97AbQNNai9Mes1R2dWGPQXJlhst1D
Ol+z3HV8TcWSD/czPdIrCWT2K3jEcZOwydFHn9s2f+wiDbtQuCAB9BNhoj8eN29IbiPA75VIGccQ
SSHAU9JM7LAwERds6xEn9Pzrb29YW8AfWsRwHx4mffmiCyGuH6IAkfIs3GlFyq4C4/qzXjeDohw0
zmAe15gsj1/Jy8KMBfX7WqfH6UtpcLL5/jKhMAB+Bvl3CVt9utq05MR/Mx1mBwNFMeFsUQhfH6tJ
FywEa7AQZlMy61VKQIPvmaUcxam/JiNONUsnlxgboDng9xE8yWydDrA9jxqagfuQ0Ev+e0V+jhKX
2TSOUFSPxnYfwkc86zbDT/l9T/t6Wj2ftx+3gyj1enfnhqyRh78O9XBIiXTA5VEvxVCDoJ41/osq
AN2DVoS5QSW/3hInfKEZzWjKoWf8nYKp6aDi6lHHwYNCn+gxH3nwOFDBPxfzeZA4Ayk6ypxk/ME2
HrzpigJ2bYJp8i8vKVBmWPTxMr5/gLHSV3omz1qVHIyjE4FoHus1pcZz3p2bYE6MBPLJXD28v3Js
Puwe+KfvIj0wrvZHKCKvQy4STYsdIMEuUvVJZXBmaS/Q9ALgInAswldj69LIT0ksf7LGRrJQ/GGJ
ez+/oAoxBeiqZ42GiQdNobNuwHrZkxSNrs7GcS2E/HKLfYzkRnXGm9Q/6DUKXs42LO9aCBdDSrA5
HKodr2MXs1UNmAT/KkzYqYYAlVRTiL3ReziHqUW+xcprbS3pGrzQICMqsTY5SOToxCIrArIMiQhp
kgqPybIa0DB9PIgv8XHjWPdJhJ+oh5lHjOdY9toFxI1Jetw7mb+LM5/YOEB6/twFHurkpd9fYk2T
XCZant7KhYhEJD+rvo6fUfWm+D2hhBINS8SCFCSzRiengmpHuLSIbzmUaGOj7jmGT4uPRdIb87qE
2qixwfnT4ImgJWRZLWVMRSUBCsj2MNUWpjgTiBHF4UIOjWN1NyEvxY0niwAwvZEWW+ILwe19FKKQ
7Jay/8UNp7YmpzUa7uM4hpLe1DbENhjdDZ67CeqH3mc6qH0mCMri6VFWs6S/FgzhOrBaMFNf0hNi
Jc4942z1LqXBdLWXkjgFTAjknsQr7PUrn59F2cu8z+0nvAq9BPdQyUf5zv/pPgNrAJG0JxVTUYDo
nLmx5Ysfx2E85m+zEGWD92EsLamTAAlEaZiqwcmGBC8JhQEV0lSNGjayBEliypG5ZCqfYPYzUQJo
w7sOw4fzQ77Sf7WUANYj2DEK0KXtQhQx3hFbYkLEJy9onR67SUVFlzEl6HX1uOYm/R9myiSivbwT
Ds64pdQzSCMlZJBOM5GuaZ+TWTqsjS/HLiFGWe6BoS/2CCDaZKaHeVF9QZxMTXE28xQWUVDPzXUP
UjUGtPxK9k/jhkkMIIveiJ/lbuJ4QVzzP9IYSBO+UNK/FURb2+WjNhWxv/EDS+tHnVvkDx5zfw96
9D9U3QRYPPElMTa7ZsqrSPowlOo6LGCh5v/sP582U+IgURxda3Pmc8V0vVOb4uNL8zYxvQ5+zr0s
jPq4c9pyMKWEu/mcSrbKFXeit2wktDytmcSLz6mMK5bD8W3Zqz0jh3elADjJRmffkE/pIaq2BQui
KcCLoDJpkGzL0rpNJYufQxJ9Rz6kV5aTnpGSewTDyANVTnhjsyaytW72wgyk22Db2UG3DWYAMQSf
M7JXXAskKPlrHiPXragyl2S7c020FFNd6U9OLRxaY0tqjmqz35XcE+fQgV/k/g6QmQ72qoXSwe+D
j/Z9tIvOrNaFXvn9sz3olQhSN41XizpjQj2Mii358NUYnPqK4BhR1f7WDOty/P1IEP6jsexM1E2g
6rs5vSEfq53LNgan7aCm43ic4Q0asUO76fMZ2gNZNWtNrDWMmwRUXbIL1Fj3i3SokqssLfYroMXr
SvR8jKmMnmlQq6d8RbQi0JQk2KH99B/vTMtoRXuzHwEgHJNFVT9nFnRTJKYLVG+OI0FVy1G0XtCK
BQsHYHwtFF6m4BsE+YWQC7h2BFZpKKEO3DSCOZ7osTAu8/2JQRYPHDA8iL/Is3QCqBn4wptXUZ6C
vLjUZxhsUoO0C3JXthTQqguKltfCa6GRZaUETstTX4TLDq9WMrteNdq7oaxWHMxn7UG43V7rQ76e
pIfQWSCssqyIIzh27fJm0SJIDJqrCcOLCtAVXHE4eM10bMfYBRo9fkkRMB5R/666Xr7vUO44s2EH
csIS1eyfU49O0UNpROknUN36yWqH1rBx4HQz7zwR6j2HKyAHX/+KTXCeHPmHqsHhnu7XilBDlAGC
R5aQoz053txGncDRowgCOWaXRCGYEqSxDUeKRpHWde2fYr206IJYhekP+91DtD5Dn3pslbizXv1K
IIRfVsssSZBe3vz340iD5GCUwPRr7MvDcaU5NhQ9bBT2bdJ92pAoK4JW3CBTMlB6N3cMyivtZXUv
13cRw5KMOCIMzuOmL3Mw1/o+iLR5a4TSdqt8IMejKK7DIAl2J1lZ1qo4A0EB+QorykR7xp5mfdWK
d/mCq8DD2N9rQs5qsBvQiT07zPPrU0iH52p38okzgnMeQfRAO2l0wnl+GhwE3Anp5aU1m0X3UZjU
nItgd8uLBZ7fs90jEvxEmTZXegaVpECu1eKqbY96b6yae/UDDf1GaqsSpv88ZtpBmrorawRHS9v2
/rq6UHtpMxTUg624w3K/307l4elIMc/xdnmdUN7Iex9s7QIerla+7c8MjkZ7KEVJGnqMZXixbauP
mgMPM7ldbYwtckd5V3q9mjcRLHxuA65nmlS68YEce74JHKXoVZKd7Guu4KtjpTzp/9wGFdA+0nEb
LYm/xmczz3nm5yMkRLnh4fPaAJYv1Xfx/ZJ84PDPBVy2DrauMTHM3H1HrZU+UdLs/eSo21aipAZk
ZBkylcqy5nj/HPqIEbIbzFe0YOi4v0d+yLcDDhXc+EvekIvCXX3E8sPni0ui0J/jXnMb59EdEESa
SPsPef12yWo3HthZKpyq+XVLOZfK7S05MfoH1s9SRvTCphSUQe3QIuW9eaPpX/sJCzzFwl/x7ilt
grfInKTIYyHcK0lYr0oaBtELC1dE6xwmOLY/LLlPasjeeczenH/2laXjuKB/ybCO9lq2mqbab7YH
sc6joitB/LqiiheMvG1CzpJ/Yf8/79gIvIWGMWVqu/vH53+V93GcBaEiVGNBOsqhuMy9bVZGLh7j
U55GvJkVwUrKWPaP/F4vNbC0M8t6n/O37U2raCeCQ3JntWy+nj/RyRg3TfMywysG6QsSqXudlBL0
ds3MXwNlIZ6Q3qLyqeGHl/lbkT88vv1zLQDUoCgQf1/JK39grRCHvCCj33gHq+znuLHmLper79GL
JB0mUwwknCx3tH8j/MILGk2jTRsC955XFP1CMjlLGJanjxRmJFtMyNcdIfj5+c5U1vVF/iqFSZU1
WjrVrTEIb5RrBh/jjRo0PPnhWlHvTdLW65fRCRWKxXWjRkC7kO13UKksxjnmQIpYK/WVE9bzlC6O
srXk3vWVxt7+MAzmwUAUBK3WGCr+cvOhVFoUpqpvt53XLsHQf5HNq7XXST9OzGi/6zO+ucHfHrfi
M/rrRRzJrZoOY3LINMLKnpczVcZpCKhi8TLtoJvXZs9CQhDQIwYvEPE8cD4bA6Cv4Hjj2wUIaNJg
KWy3wKEcXr7ZSrnAuuX6WYBOK5R8yKYnrS9daPAaeVtwNOF1544o0rFc30NxrG7/P3OZ9dtk/DJ7
A0hWRlPaTVuqEuZ9qlq2a2eE9BxinfjfNTGOFpvefptV9dwGS9JUopzV+BpCkStRL3xuASQcG1uP
XI9cKv9o939PfnY2/mR/CU/AqHk9qw5AMuvIT55HqFfbx3nYy9AXoaQ8+Hm2gyMUQUN+k5NWIF+H
vjkdooA0U1cFRq9i1HznCLcB1BF3ZFc6KMxWGUoXIP/fMI3RVzfsqMPTBCfJL5qpTvUjtrlZ6AoM
ALqxKBSXNDC1SkpFqpd3IcL6Ob7nq+cQ44MYuexnIpgzxDS1+6LXp9HeKDSKzJ/oR/ANVHM3wJWi
8KAehBms8PqdoES4nqurqGenUw7j11z363XFVNz9GoezEvsTo1lqKPdXoEiosHtNw4cl2BkkClqB
bjVhor8zpEkcaGAhCsDNEeqRRmQfPDVHlKwI4aXOO8VNFDygpgXF4G0dwUP2jMdAx9LVWxJ9+Wfq
ErOfm2szVN1n9pyJgYF6jsBe2CpD9WpP2mHTK+/x1m7wN2DQyZO7gNU8D9ShUkVl+eH3ivaIZ0wN
2pC5YDKxWN4hzI/cfrya/L2DA34XTe1aF828PXL5+LfmhFrNL5uQfjk81Mb1jkUT0cuUPEeclxk0
TFnwNVnVsicHX51rL2bCN9Mgp0mrDipNUrIE+cFDozOZgjpsLRP3HPnD6PsQ5SDHKFtNg206gzvA
umu7jk1rKNvNqrZdNRytIwUm+SOoDhxIy6lBWJk0LXZiKwGZ9ZHqPsxUtzAJDVjgKYA2e84+TixB
cgQRMNb01jYAOu21Ja6utBmE/Hl4PaJ1dOqaVutoogysjpUCA1A37u3SVwHfX7sLDO70eS65chJU
8BDhUdGFf8tuM+R+2MbVSN1zCR26rnNeZr9kJMS3z2/1pcjT7eI7GvFhlCtIfPi/y5GDkjxCMKWc
rA3gWSfWoCYa2hQBMRm/4N5BTLw3aPD40SIoeHzSEmp0up46GvNji3Zt/ubwuTMTKqEEl9fRmOPr
pajphPiWfilbI4/p8ZfKNXKJq9Vq7fy06QXcys7X3AzLlAXLpUBqysZlOGoya8UTyIrvJI3Gq4ug
uCF8bX9ompgGnPN1UmohrN/Zj7vV/w0p7QrWhPCApEA2lTNKsF9KBbMZDuKx9Xg3wqnEMoEChPIp
3KEyK/AmCU/uAPuLEoPfqs/R16RKZHJjd7MqcWSkvvVH41WpNafxnqJ9wUtbV5LR4oV49eek6KHk
cLTlVK7+AwLiEAOtvgBycJ4AXqS6N2czwcBPdkgt5vXBaQF18lNXDsX7/P+IK4f7viIyFLRTxHr2
N/4KXDj2gJrTSOO0nLtccgPatihBvZ+G3wBkBeOj9Vi+chEFEDvkUmrDPJ/zPljP5O4YBK3ZrNCr
g9zbT6aG+sv8RQAYAU/9gkxtnkaAltaWn44HkC4ZDyr+TpNeBfPOU4mzDN2E4rhPHz+TFoLvF9g1
Sk2A6OcfyHVhlFws33K+bIQ9XwuvYQNG9Cwq01KfGhtRUZVqvLp1E7t7MJxqijw3A1ZJ2UjI/1ro
mzIjcXk6vzP1xaR5U8HbWOzKSSSGWjkyHuN8qy8IQ9E+1bu2a3sVkgE3/Dl3rwqIpCqOUeCmkfSd
y0n3RLj1Bb09Tmhu+P7cXxVuTOpiNOuWC3ag7n+kxz/kWTeECQyPEQ6JZYKrc3in66uSVjdDhoFC
Ar+b312RNovrvGgOngYE1aj061Nvv2c41rXkl9sTwPRsqPkQF96RT6yPvZyoJjSfAyqCz+ilxHvW
JR8LOOacSqISkD/NvHMls5p9qAUlYE5aAZfo3G3PjOStbEhs0S7C91zBCXcIWK9KiDbrBHwPHxvJ
HE3TiNTx/XrWlqaCCza5qCCuQUmVXGwbQeBgZ6bPuOaONBa7xezs6DGoaGSpu4FCLXaO8w90kwth
BJAM/givkqUoNzRR4LpJaZvZW8r2HbvIrIGx9y2Nbqeqvir4PnRGAwV5zzpnqADjj1Dw3adG/7i/
zSV9OrTwY1mP7SjXm658tZdUViF/aN/BxSFz8YUdbyQnomPtcA/CUYNDHsHUl4LyS7fnv8VvOD6G
RS6mlPTkR9me36oAs4uW/uMYNxmlirUsx50+2f4U67sFLdMV1wiGNOwN+k9Q4vuVW2XjUPlYpLfF
qrdjUKFURXre7L8U2QGn/FS9vDO74vUnGLfowQEyXOtqzjJ7D/BW9xo5YGgSOet1yNs9IV4DbPE0
n2/3lTBB8pz+wwZ7QCC0DRg8XnQxOVu05sBRHj1E3aVHh2gUAsmuLSKLyRD0CHPLdyx4quBlBTu1
sOMZ/WJGwXkF35qlzpoj+rLIxCxO6vzBkInelpG6IQtP0H7meIokzjnlUat2acfzJreeD4F2RP+y
/A0bG9uTBLhsCf49puQPSqZF7U0mJGOORs0XsfMHoOOWDakO0IplHTyDud/s77Sb5w8Xz/Yol9eH
J9ZHMilV+giu+QvvgICw5//rQMwQqKl7XN176fcIZBRDmsXQKW/unK3DNX29QuevxZ6MwbLhG1EN
S0x4xM/cUJr96XJGBaleGBO3tklpussfo1Ofyqrj51LbvOVzvGboOTSG4AwwIS/24YnLDwaI4yid
M54Y+/92P+PUdxYEGkwz2jvgtjZBMJC4kQBEefzw2FzqSxkAMVo/Nj0x5jlyQ3kboxI19hY2vMjD
/GC4Jn1Bk4Bz43sua2E+U2ebuwV1d8bdGTmDEK0tOv+5wUpM/1txCuOkednUGjECnVdMj27m7K8g
bGf0QOJq7CYP9rpxj960mBELKI60bzTs6oPd1HbnZk0PAO3RKHaVeoOcvYZSA8hpGQw11rDEbroQ
rMvYRTg1xaIDWzqqmzZIHq5jj37K72si3UQH1R+cLCMtr8a14L2vBUkdGk2sYygBs0sPwdkxUFTa
xKIz//mpgg2Zd4ayUhv5Z/6TE3Fly3ZodCNp/P33hQBA/xh9+1v16Slmn1756qYyJWmezjZERHTv
BBl6xbcP5KN321rsJLn4uFq9gvzBB9NAubyc1FWp1DjSDUO0uoY4qwH3Kubv0yUH7foquTvT5fj2
Ke1esXB/y8mc5NPzoNI2Xo5r75UypmBtLsZCwrzlNYXZxLMrjKMGJcgCFJNx6gScjwAORJk5mH8U
kjftXZ+76rcJFT+lB23CGn42SNA9DkMA0omsFRfdRvBIA1g4/px2WA7+SrgAn+e7YDAunB/uNbGv
6P7cg3ePpIhwfLILughdzOrP/RNeOSOBN1GVy+OKDBRi4/HAE3sGNC8Dte1/aFcIVJbwyAxapnhO
7Dft3GiPBCS65SFjK40iP6IP2PP+VHruV/kk4H8DDAuYdNsTrHku0K/U2e7hQ9kUkjW+C3Z6hf5p
mVO5D4B02nPsi/QtHEUQGizAP8joBviPpUGf49RMcwKiTbSKwGEn60FwcqK8avaOH8AxiTsT+XlA
p2nBMSd3xuG9eM7Wshm/nW9bddQNJd1u/LbGUptXhaIV0mMnfgWJLIeWefW9re6ePenH0Nyn5vkk
Wx2tL0L7sRK/1AGpGsuqDA7SbqAPgiqleoENCeW7JNQrFTf9BpHH/kXwSdTP6H/0R82I5KZyQ93T
oRwkMV7EG3Su+EdlY1CrIYa3HTqO+DzfrU0RS5EpEptNQgWY4sNDPjDnx33eTiiHWP55bD0WRS5f
jRDBCY8OGyErlzU9i7jloHNcq+TAry6lSCEq3IT7/zAsK75rYNLJooV9yiVaytLJOrgk2BXjMzzB
Ko8jLMIr6A0BQySB42VPm44pMGsioLCujcvrdoLxLLbx2Mya0KenwIbvfB9xIZdKUhfS/7jMVdu5
NVvjM9sccn5vIjYtJngENOVWEvV662V+nxuThM2NHtDsmFRUq0uqLKWZViEatGHk8pwLTDtjrZoK
88LlL98XBPcYYGmiVOrrceSqc3tBO0QErHbsMqpYB0Geyt2MGqCVuF+SJXDmO7JwaqXQEecxu8/O
jmsEY1gWF/SlLfyW+u9I+SFqf0XfCeZuVYt55mz4CGfc3MuOwuDb+ufN7FaGMe2bflGhJvWroixW
NG0aY5RDoZJJV8DC6GMx5E34/fN6K2FgJB4sTw66DIYghO9/ZAi9PO6gY+Sv5FimJVfHVtZkskjS
QZaGqCC+v9s2JXdhG7O3WjQazV5F4sxoNQS8U9TVBdWhyoDomRGGjeawp3ZJhMwePcDsfbaI105Y
Q6o2ySxYjL7iaUmo3M/D59wSynkhzG4US0R7p8qL5QEU7UyFvEM9ENpEInx/B5d+vwNFeXzvcRQl
HfKRL4Qztqlf0SYb/G0LaonjMNIfMQxXLFB2Y+OsNjj9w2VQZGu7PfKLDBFTfKlWvL1gohq8jePS
GV4kAYNQ1eTPpWfdQ2FA3YgSHu+SUZPV3hU4abQQMkF3HU3IhhJ3x+pYihupJaPFnUuP1qtumxT+
6yxfk2h6JJOMBgTl01UVmkDgzan7hGED10cd0eYVO+087sNY2rWAsXHHiFUL+JYhgmElZMVni5oi
O7ytNd/Leg5u01CyOtpI3kpt2UX069JjQS2Noxzxq7A8Cg59S54+zuRXuVol6zQdBvPYZ3cCttjD
nz01wO+dBR1Z3kGUUJxP3XIdmIV05ZUdxmP0sFigXPHL/dSFXATiLP9uti9V8NYctB6Q6HdIm/3a
drDBjuZR0+Bz4nMGi9aJIw+6GwHPN/aT96UA21LZs4Ok79/frB68mU9VXHHAImBT6D/yFBxD3IqA
8VHIKZgZ0CUNp0oBNkC3473hn2XlWulq28MVk6VHcBOwh5oOpLhCl+B2X06iWAfVKf5LH0RZzX6A
AIU7UpLUaaNUURVu93x/E0DmmdTMdSFmmq0+9Jl1UOHXR5aWNpYVMgw+dOi6RFoD1TApwEPd0GGC
w1eW+bRk401+Av+ILHuGZnvrGbOHW4Owkfv5oUEGWFAPMwoQW+5Fw7Cp5oEiU365PKCdm5525rIE
XOHj7jlbjsvQdPPPVn58VZnaTz8R1JZZi/AMSTKh55cQO50Stul5OOqZWV424qcum+ladcs63dYR
6QlegauM03fkqLxGXPjS1l8qrrtEltg7cJ6um1yRXdnvHMMgTAWu4HXHbEoG5f3MkBdEubD3TLXg
FdDlyMc1pB9bGUV31pQSzqNYCe6le1X9OwcwjflMGPacrKQNTId/A89tVMalYvDXANcglEqCxxUU
9QJr6NsybrdWw5gep1eFBgoppDz70bLJb+rvddYQ6hxIsn19VNH2T/DhabcfvpBl1nBKxXKm31lG
L2V0oXV2/3Gvj93o8IseLtaeEGiE2NWS4KhStOwL7silHTj+YVLoKhWOpBEIpST7ZLyE6nTDdVtV
z63wB4368DskuQJWZHup+NdwX2lLq0Tofuuoiox5igSt6P4RSvOIbdHf3j6L2ROPts5sAy8y1zuw
l8DT9LcPs2ce4H7+YXKGR1eV9BKQSnpxSwk4mNc3UJWWsHcvSDNK3yrQOQzL36xJT10nkYk2Ipus
lxKq1tkdmqSh50IXOKGV7fJSjxnc6DNbBHPUPpGP9PgygcDWsgVEAK8QPdEyJyLKGm+Pksv+wQuE
t0FY0UZ0l2vhFgYIIoWnnivpNmuobr4A0vaIeBgmzOSy0qCUO3MO4oWaZ2zAFjJh3oAjtOrYL8g0
UnbfXS1iriwVjgZ7ayX6YGvIO/iPbxBamkw9NC2L0sTqgME026AlJGVyugg3LjQDO7wBkePILwrp
L+mmlVCIIyzYThlKfPq6Bq4PPHlsoPVrIgRCPvH5kMvQTMzHFnzjyLCpPcPYaNUzTS6NZBO745yj
Cs0+Wjb6s+bIUkvbVAhSGm+6mj0baO7W/yQmykWvqPzYX3o7zGenEDT3jNrNQ+uxpYmWbNMTSS99
41a/YvVHy+9Pf2DXmzVgDMckx+Qv+TvcANf+6j636njN2d5srEiZWD1BhWs2aYj+7xXGwcjfqMCT
LRjWfLm10h75U78pm9VNNLxORJkOmHdil8WBDri0DlvbcrJpjasj2jlyuEJEM3zYHzG6dUnvBids
mT1DJElY677+YJXiwj9uyQxE/8W33aqNHQISIUHouB0PoeDJ3qFoToU52l8fxCLv2sJ1wzsBZKkb
OoslJu+/R+qbU+EBgExUav97WE83BurdQHtTGi3hmvZcZzrUm6OU8A8aYL8LbqO6wnlHQ0GsdJ7u
D85USN895CX8diuH4XfsLhcBQu15j8avqJvS2m+7VyZFEw9CsVj8v8HeP/CsRb6dYfySRtudQ52e
mfGQcn1xfO+wuElVJ2KvPOe/aoaZmxlOrB0qi4/4b+ZJ4rJF5NBGsAecu6NVZfaU2qM3fiiIWg4A
5e8tRfpTR9AT8yM4/j/PawqqXYHGkphrzLTYbH0dpehEVynvg+70yqsJHwHbK2kMKLL/LWf6D4kh
aPnCq2+Lz2NgMHZcTj05QV0XD6jzsgl+nohl/mJbpTmqqalKnS5qXAeRsyiW6fNo1Wfip6pkXBxx
h5A8xZS1jNj0Eu23G3SD6EsmMNIV62PsTwP74Sz2jd6nowSrnk8LSUxanPy8bHRqOYNftiInCvf2
LEZLtv5t9eaTy9GWmaTmaHFIBvw4xpZPRahStmr5zfs/l/QaIhVNOT8NkaqVwL9lM/VbNwxXzBvF
7ZJyp8xbXN78jhVFJ7GVTO1uky0tTEOD9lYXHqA0G1LgwbgyL4NsMqOkETNzj7byVb4z94u6IcxY
7re0z9sZoNz1Vc+cW4DMtu8gUTtgKCX5ayyLKmoRpjxt/Fp9A4OVNAJO5urTjNg7mQQhQ6YIk51p
uXxL+Aik++8Tc1qNV7q2t32LZ1E8hoZhduYTX5QGyINnmbdGdIzv5CDRLn7/nXDkrgKGn85Lpx/L
j16ielruGXvlO2qAqnDo/bPxQyHtiDMP0aZ85oN9RpLXQW3hpT4oS/FWZE18hg6SMIVc8WzRwQyD
6pwDAEBMvXogT0H3KPPnAq1kFXL+sGc7VjcwCPM6BHnUUy/00D3wBAZoRyWQAUU3CCcbd9NDP8q0
HLxU9slh/G977OR4+dkBEROKq2O2FpqGXFO7Vvptcg6gOWEnYmdFkmWW4UAK/e8i1u1OFoTpOFzQ
H/ede2AbjUePIjMmeeH9C4yECt2zIzzX31flh4GokCJRy5lkDFVDUhqesw61uFL2B0DioEqAxDjF
za0t9ZikQuhOeW558EUFaAI0Q0zjwheuVI9mXTySY5/L0CgVxKOR5DERLsjTU+fZfPWucyh8W00Y
2JXKbk5pWSMtZfYiA5hkInmr5h2ZREqImWr3uQUA7KNillq+l3k/N6kOSBUOeRZbMlaZQVT1jZZG
biRuvW4/NJsvOjP+COgoRVDNJgO6gZrMGERfw4DBlKsL/zkYxm8tpaY9Mpl1BPIAt+PL5Ie5eBF4
4nr2kWY/+8RIJMp0rVtVvxjdnxW55IdJA+65R1pA0i9kM74Pd+pEwdARC/Zcs3YJN7MsDqq9ptZZ
hJD1IMW92V7I8qt3IrgqIXwjrDrlqDzRZx0M14boz6cAaZwYF061cEH4YzOYmbvIaePldl/0sLpk
czyQpUcek9UgpKQA+19yL2udZOCPC73OvFjgBj8/N55w7oxZE79zqaE19RoL/aGiWUmPh2z163w3
BiP2iwZghdzrcLyWAhrKULPDe8kRK7oubw3iFuywluUPjh/kxitjUW7hC5HnnuOmQHhCmJVf5dsD
H5dGTsWiY/KMAv8vM1wk3IB40RwQ3xX69pQmzcK9ovj9u5fsUZE72hXvn31EYT5D4aoGuWvuDKMV
4kIBn9hts8DGPA59xxCDkTE84Ef5J0pFLvLNKTiVUqVber2brFKdOAHyEIQa4MHoxdlwBFBZCtgc
K6SOxeKE9s0OJmscpB8l7ECNrJ7yaTVYIhmEaTpIAehRWBQ0rfRQ83/tZIK829zEld8542m0XJVc
nkFlW4rDdKAV6S+kxlOVLlzdBxXdBy/5/Qkkk8Xaal1qpYLZQri8hxGoW3cfifH7ilJ91ktsUYOG
7+9fAnvcxpPu/dvZsO7ndqUdDLPEfeaBP6WnFszUBROoChp7yegA9E6K2OFZDlONnkdNuLZsTQEa
3cjnu1jE0TPZG2Lxyltn8lAugObj02Q+k3WJTuyvqXfAZEz5FFT+5Gw96Qt7xuxawNtU0wKb8xVm
dBNxxouV7ZJ7SuJCJfC1s7NWTrYGPktO8ooiyTkx+r1bDqMvzmSSDAiKONV5dpk3gxTNXJsKyvP/
HGhpjedsOKtpvdOIWO8dA/N4uc1b+ZInH51hp1vCijrmNSz1EB2DII6a3YkKSTCrsDb5iNLbCYQR
EEfd/0b4YYPolkqqj6a7unxabhpGdAuXHOXx0BSPsYH7cLkvhAJC/1k7xWS8M2SYlgXUl0DurYcA
qL5AwpGl7sCoMDD2cX1Mgugf85c35/1gN3J7yqP0p6A/y1A7oPhma5yP10fszeyVi/UWtQtxLcxm
3P/fin/jExqjDGWacWxnFtNqc77UmVSvZ5BN73SOfzT6yUiqQ8FDpriuPgJu4vsjAOvUvcCj2llo
2wiRYwIpTpq3xglQb1qCdjccqrAstW0w5CVR0O1o13dYCmIAIgDbfB6IxmMU0MXLgiA0oDGFaVHM
Zha2l+2BZLZotyoQdv4M2wRPHplrTgoAqwSRcFUUpAfrzFsiReiS86eTcLG+R2osJN77FKYrnjBQ
2E5BO0GJHUZwQy+hrye/dECdqRWSA/qYF0VIx9r98p5+gDXQitKywRqdK2cZtvDYD58kws3h0bxH
M0XMh4RHgTUVHjhPLUkCQGCmnvjsTlzj1jXrIwwQMfyffD3n013/Ecnu2ItrHqzydohGoWrfNIJc
RMkc9oShufjR23s3FbXXNj71AxT7Z0o1dgiE06ApwyJ9TGxcJsUU1V7fZkKZu6z9SWj9euuhzmok
l9TnUBZBMuoRW+ScYnk9yFoC1mkDJRuh5LLn/8JoCLG/IA5WqMBhRDjUbX+hnXoYPvFpUI7LTqXh
0oYFgs3tBb/B5KLqi8tLhO2rqVX0Ax6m39O6xzOjCErjnThSdoeXsu5y4YAE9xspILDlWpGS+usE
QbPRo2pLcpqqKlmZWRRUeOxIykgroEm/otJyETeQ1G29Um7DpsJcPbTplqWsLEtl7YFDvqmpEI9g
W7++dMYbWV8k76m4oB5/R4UKTrA0PcICviAFtPXwq27VKlCcZJoFA0uCOMiAo/g8UgrTT0ErlWSd
eW9sLHeSXCHJwezHe5ozttbAZ/PVaghdpiX6Fh6gE8ug6sIgi4lV2VycO8zKZ1ow9bjnzSSvbA/W
RQ+KdX+77kzL3FiLvGsjvLrgdpdYSTrlf1d3L+EqUpMeU4wG5tktBbhhTManN7gYQaTzK/i4QWRo
t34VI7VXa9fLVxwWe9+tiEmmX0vTsdpEG6S9iq2msydRp/sRJVNo7BAIteoudYaz/D8eqPVb31Ts
oOV7tfJSdSDb0bZVZ64GPoZOP62MbR2Ge3QkruCjmlPqYfqC2hT3pDGhviy97fLeHxcoVugihYod
7CU9VvLkVom9JSkiXIsewkEgVNcbV4EGk/KKM+D11Ej8T9clJqpY6F8vbMs4r+vxrVNENHAIXQag
1wBp0lDAxhzBKNV1A7f84vpb5z09fWMkE5m5rGnl0m3F6WWZatqWhhRlkIxBKB+9tEEaiNQljCNT
Digf6SW2eIVaxyR+O3ivbstwwQrWaBcOB6Q1FbNENbmJtRX9ReyUP9vV2MFLezurBqyod/b/aW3n
MvwJXQ4HAQLt8YZZl10xwcMmHnvWjd6auRm5sivBSkwNl0rAMNo5u9g+HCHfDAazhE5JRGjGEQ2j
tyMXFQPB/zH73WFDqwUtibg3UBS2zto2zFg027ZWOWLksHqODBQAW7mqrKAIxb8Mlq5rerGHxgYX
blQw3ZKt7HNwS2Z2dlVEfww4x1TttXxjl5mmpoBXZ8XormIk7Jsd5lNIrXPU48pQxeMbu/iqGEgg
oS/dzA9ovqH4qIvvIFNYuiQwDMg3+1S/DKjBERN/tFPXKQJ31wlx7/qZk3kwkty+nzT5ASc6DyIz
rxGZOMGRw/G+sOI6TRDDSLQJS01fusUABFD8ZMcE+qChU+tBK/tCl9XnpMS3MpCWYcWxK4X/YhQW
RE5Z72Qbb6mA9JSlESVE3k4+qpHLg5ll2K5YlXiYl3V6qLSYkii58w5B6rtYwMzIgH0IklvU7eCK
UQQ6/rxpL7qnPxgXj7Mb3S4SDVkW3ehb8SszQwbjt73NmLN8hguwoUNjVQrxOWgGDw3CoErlhmny
oCeM7GYuthRDnWcDVILjJf0BIaL1P0HTIyrpldSnj5/fCc1ALxp9jbclBvgmhJL1pj+hLZ0ibdv6
SbRXb5GfOTQwUGhdKRpOPPCtu/CAlFk0/3qFHNkMezvPRIHzFTSAsdJrVsMbnr2s6L54gptZeT/o
9is0r1XGBmU1FiP0ussQEqKU38k7aMikAG4Qj/inpS2J87eELd1dREwRm/czJY+EafnFY4xMcMLU
qza893qSpf06vOLu/mpUo4GKqKZPtlmcArhutG/0v5DhNY6o+s0ykSe8NszQYitdXJkDZ3vKAmxj
oPGlNCscCkHBvLJ8M9MxX5kJJBjRk5BP+p9xphR29BvYLK58H0lBowahKUAGTwTu/GecZ5ybCkVZ
Ym3XoGAQKYG/LKxNljOaNp0lPrURkMcZV+OX/FrOzp85/jaYHTcuNiOnC3KsTRN/p1gYnSpn5n8Q
T70C3ghbCWDzEgsbS1mWW5RnSeUza7dTBd59geL0sxlHsfn3KpW2lLQxxHE9uuQnr4nJ9OMR7k5w
mVTyWcJqIjciVcckMi2cCv68zX9APYhBxTsz5ZfTXMsyl+iPKlGsMIbmdbHCuIPpFHNn5uH8apMC
SqQBmKiB/z/RFVoLOlyDtunO1lQncaCAdn6phDzIH3UyZsWK41DB80EqgYkXfD1/2lqXRq5hTKDj
tAWyKlZEqsoZlCAvFp1N47o2KSEx/NRx5oOI+gQZWNk4WrpOx8a9J8xehR77G28SOVeyc0K5naHt
681W0sKGFRK5LpyuS4JlZE9dCrBoHrTc3UWHk9sJAd2NgzL/sMSf5iK+zYWIanTXayeBynn+BcJP
arzdcP7LFf9INM46FoX018Zk4VTtvlcXPDwYZEZy61mI+nbwK9qignLsaFKvcFdL4dv7wdiTeyEL
eZ5gg206yIUAGuLAt7EtFmknMUvWVcIhXTsrf1UPww+pZYZQYVhjPLfH32+rWHtlac+TL6Iish4v
oQXOgYWQF4t7GvzsbXwbo2jW7o/CbI0DDFAFU5cmRF4D4KCVQ+jd71kCTWrUGVy9IsQORma2hDl/
KGlvsZBM+kIW8i0p4QR2J/R+Eg8eYE3Q3S4elmacHVEHXngl7W8XXd3tnki0O5Y4FSZq2uL+lYjS
34E59e1q3Ktyxzpw22aW9Y7VUpIG6ijYD9C9r0bGu6Xf4doJpbBpZQYaHeIDfnlyT+OUtIV6GLXt
LLICJL4IeKCtm6wLnoOb5smAp3733EDMPWH2gdmrlbXa1APPUyXF3SOfGb5FR033Vdf/LkuPePlE
DrKswmbm0E6sspm4aTUbIvdOO0l7/I+LrAPGf9ZRRcW6LJeB050qyyzG2jmyaD3qYZDn1LT6Sv2D
anyf/aYMNvdEK/jcA8m1Wvk7kQKpiFsNhyr9ym7xViGpgFda8JQJC9oigbgWsTZ53XeSkGcf/huw
IXUlh9tZp7IlQ0bqQ/uR7krGOGlMsHN0i+K+vLpQ4zrhFuS+JCn/88YS6rpDAl/xabv7HxRB7WU0
wZ1VXnyVIwSL5uLFGnSOIYB+OS8ia/LNgq4UH4kP7FwMJ4VsrSMVgIk/9mt9ECm9V7ns8JyplJJ2
AyRhKz43z5fzocBrQpmcFto/eTMejNCc1WwM+KgveQKbrZD5VoELUafNWnOlIQDHjgndYDeWtyQ4
fPoP5y2MotO6bTznMInq10YCQwrInCbMjKNBJwFUpWKPFrmCssk1vajMfpxgjK7iAoF8DDu8wrz+
YrXUu8kk9eYVVxEGfhXx3gvz9rl13CSHK3iNsj14rt2zQND0A+yB835QMm+rel1MDJ8EcBPxWhLd
HaCAQobm3LPOYYnFCIvKOaLT4UsygzndIpC1I4boW7vjdq9GQJ7ZCXKCMTxJo4XGAVddXxFlWOiu
xYQdO0QzLLexdSL0JJmUlvxNllH6W7WvjOg4kKPIeTY6pbM7hjMECRyQwqDBWraw0jeQHqAi2gbY
EDMKFfE8XfLwQYx+zSe9xKXlkaTrBASfHikCvEAXHx5mJcA8M0jIolIVnMyt8d1x8TmVtB7cJfCh
cbhlTDZUnjXHN6TXBLggiDouGJDbIFyl5RDo+FL/38a8G/R8PZNRjQ9OCu9bGBnvfFSsMDX5Fqv8
WoL8yRsP0gRkXRW1+qHecfRkW3AueulQYWa7+bhKCZwOfFJGGneBWZMwFZPQExe7PsrkjVQae/Sf
E5bS4jPPzB+Ro4JeXS5j5DuCebZvYH2xviM65lhGUT6AF064/8j2fJUEMpD8b7C96ZVHvbsi024Q
cXjxgY5ds+fxa6doXPTXcuAyGfHWVxxMIcngD2v8APVO23GrSWJaLnYckCqwF4vOAskwdjMxye6k
5ATF6lLSJbJbhoX1287CX/PujlGlAOlVOpXw9TpetsMSp9VOyZG9VOQU9ESdQvpTCzbn9VdyEech
gAmXM5PXpyyK86diJNAZRIGqN3K2oJye9ZK3I8F9p1VRFHx6ant/IS3DTPO8Wb51s29RwK9p/TEo
j38SFuzWh+8YobMwme4JMRbemnL0FpOq5ZI91k7CDy3GYN7h76KYK4Dx0t2sbdfHXqf1mukUZzHt
9a5S+0fWtRNaI3UIb9szpUjUzkv6T5KF2tQBcErCx9GaplV5ovSs1cv/lij4IwpS5i5OfEIrKDiL
3j/qduvZj+TS8zaOr0NHApSjqKq4n65LZ5HIo2/WNSxzQb7oDq69eZPlZIuSZwe2ObCf/PE4LY+G
g+8Q5qKn5yEYGyZNV8kFOPOlsuYt4KTy1XJydChLwC35QWrKIEJaHdVpB8jbSWhwOBFJqJoPRb3E
z8fwoBlpn+j0xT3ObfOv4MI0R7bAmvoa6MrFwbKpor4b7rt/pRLGMqo7N9f+tKzFxluq0CzXzaha
F4VIeVC14d9Guk4ZIBbxiGC54HDwNT0dZCiQfeSuWoaIFUeKhy1b76F+bEINLSrCeZipszYMFiQR
X/y7kbBUu0M+Qsjdc7OVpOdpDrModpQaNEn0eNk9YQXyM012x3SlQLak8bSiFypJ+68L8jv6NGHH
HnTYpykVLLXcyEvpWcTD2en5sx7C2b07BGAIYAdJGqMOh6T+Fnk9WO8gcQhvFuaoZYwt8HWR588C
hdtxzwjaFzy2gs5q6m26RBnzDgtObl54DcJnW2a8vl4LHzgKOC2jxCltGQ5G2Z4GP5z5H216obgK
T2VHwPQBC8G2w0VtiTLJtbCoWU4nEkfmRT/Rnjv/15fcFMA3H4t8xsDLvVtgAv37M0EcZTzxGE3m
IKzSn+QFEP0hoXM2ik+zc9hUbmEdPexUIZEesC/mnycyRA8Bv/lW3gqd/5sNmZzBCcHWpb7uZeHB
6+7bRin//iYOv4ZmHQZ90N8gOxm7aGlVZBH14nUfSoz5CM01GwocAD2AGj7TKWPy8fdW3xyabwu6
wdXKmTfoc1M/w9kSYji7m+3vNQ/ylf/1R8EBSVVurCZtibr83gSoybSySSIN57gWh36Suwauh7ym
UUY/tAC0fgA2RYRKsv3/IshAiqQPlYVgMIAIa1053PbYkW16XoewbRJnduoDMJJNzmTWtjjYFuhC
8vzd8zvvxxDqoHRqt58tJtBKOzE1DY+DEYHV/Fa2Dk/Eho7ncTJHclv2q0x4dLdHFkWYdsPhYtv9
NhNbaGGCVzcZ0gpQA3KuemZpymrTBvQbm6++4Sa9LiIwBBUFSNvqn0S5+BWrCxpjzYjWUqLbP1ND
cVns5ycDEXLcD0uw11u739UCV2ycrF3NnHuLAtYwXsFohTYAd739Rr+OYohO9viSxwqqDBmp3FbN
DJMYH1HmBTWMT4pajqA148RQhnEpLNNuwnn7ubsy+IilnWmW/zFZB3WryzfAC3gOB7FX57ygAzWx
PnbJhOWK8E+59ngbGWek14hgMPVv1u9/4/3uT0cZWdfcrQKbfeVCa+FktaWdymYcHL5N0RoE/nmn
70rKRYw+PbVOCZbmqVu5GbunITeWgOONF6doUWloDPJ8Bk8fzFzKpnB8vCTP+sYRAPiLiN67NDJ3
CFL1/3/PUJa99TxdgmQMrL4N4mn6XVo6dmWVDgehPCeBBEq3CAX2nvYEIbf5rWTOEZJ4r+oMZQhL
SURcvyWWJWYEy09p/rZ9pg+YCx0TqrX+oQROKecrsDtAsb9TzDPjH4AdM9XbZYtu+OrCsTrLJGv/
q0BZGREBSaxRLkAA1Uxf/C9PrKMXWkxd/N5TUQq2EkfirdkG1/T+n7yNPL+/b0b+quwDIRbc3GvK
kDimGMPuZwuBxthb1BO9GQCDxe1QVaw66M70efwAVm0M+5kBYTN8+aaSUUNRmapTX1VYEuhTGO6p
tpUSs8scgQYzKQKiPkMuRvoA2ysilwcmPkH2gsAl98f8wBtdodSDTK4FDSuU8CcGfbs//KskVZ1n
Oy1qLnbsmjdLlkvdCWPyfLrHflXXzTn9IC+yK8H6WSI0ddwJmKtIOazlSr4U7487aaFOSftzYyua
IXVPNlehppWM2VUevsF16+nqoeRWYGZbUB5A4Krawx0oUMEOZJv6ZoWy7ZmSuBYv0kFowgyQ8NhZ
z9xQPdj42ECwWi5i8NvbYnjFAsRF3erShXp6H8qHqqiee4AdRiZNbiOCr3OMFZSLwszgEHzG94rl
9+bcWfSMPyiAOUHgtBybumY85U7weuUAUUjBFbKSTz8syHNVwmeKjrOTbzWpxtU62Wdl7Sv0sJ+8
NTLywWEpYON67axParAoiShlRW9/49hfN8wBBnM4+PbV756uHaSdSavAo/YxAQUomYxYYuIaqPHq
nKvWlUQtkYtKYSnisbby93yYBbMZ3JqgF5Ohud0ea/4GGQTdcoAlWLz0myi9MKnXLdCSoDbz3H9T
x53lTvjDCEntIU2Fu+ebt8HvJ/sASMiLiUnvTNfSR0k+EtoNGmHggws72R0AKC0gJpp9oflhKekZ
2lp42ehHq+pXi3Y1NnWd+KWmV/AlM6+HX3xSQFbBNQWsmHDUOpPlZxHT/FiIF9Y3ecWGPARToIhH
qmLceL0hSHUbzFbfBO59cdEnDzksg1Kh/32amsXRQI6+2+yaLkREYjYDV1jLj9Z5Q1xx6FQcGY2S
DJAW/wPZjlHAnjLbmmEXPKnX3WAJeH6fBpWSjP6Ipn9gmJKXU9Y4c1qzN+31MX+0zfEdgYXf69Qw
0f4aWy7jZHClr3i82ol2MlcoGg2f36LwSGRgruVNtHM2RNTrJzvP8mvPtddtJ+9GDspFHOuUSb/a
xk2GatEGOSJNEU+21Riy7TIsj5175vrtMKAxy7XUsOB8rpIETiOxhLuMDk2auPl+5oP1tylXmq0b
tV3iAEXHQIUrOhBYa+gsK1FcH5sQmEEQjqXS/lhcMX0XBo8XSopBJ+WDQkzYXN8zLghBCw7cDiXf
556Uoik4CKMEri8IqwbVhqVVvCkGL5ROvVV5znrV/nQpwmaNZ+QDArg2mV6oGpXlEeaIWrrb0j5B
CVqQSaVExK83ly0/b82wqS3g4WNgnfi+Nfvg1DJ3U4Nj3Jxav5vtekNcYsTJqRN2MWsfvAN0WkEB
HjAJdG6/vhVJZu4kiswkXXD9L1oWtGmg739t8Sd3NsslJGdDSvfSHqsl0P+UPJyVR/0IWNbBujEO
UQvSLdcNB71fD7RtSknCbCZw3VGvagKZfKHFQDE71hMoxjHvyOcPVmicBStHofat/0TC3GwdDbin
NP6uYifP3qLyrjudMtOjJQqr00scbjVJ2hIy1QPQ6AWGuuiCgvf7xANS/7WCouNSyN1J12eDlFwY
qBEBZpjKQYFx9wla85waS/CHRRujFECuT3p9MEK6aA8EvQEA7bYMVxa50xEG3G30rpl6GpeWaFX9
sg45NXTYNwEQmg/f9kuIsbB9deIuX3IytaDR1qY/TCv3xZSsn8UE7R9tfHNpctn8FP2+AyyDypBo
9zyXUpoKwfD/3y0g3q4Hbx1+8PTLlDQuEHG8zFxf60XQ4EWngUJkfOxDiFhDxL/NbSDpvO8NTGJD
qRXWaLTHBvhkW9kHV9WBQRH/QdsNV7lyxCVPReyb0wK9vw3epFw1mBW4UIdD9FKwCWPdqTXTir5G
CjSmkE0wcrqOp7t43Ty1wEalfEJ+65bY/binZrXdWsg8XfeMlwbJHUEla5xKMNRYAmjUnZXM+OV3
DbYDxITy3FCjC94UcJOwcE5ujtfFXwGBHyz29v9xJV5rQtTU9Nh+0AiLBEdridsJnui2mLP6QR2U
64IVWCHlsW8yfMmpDblB7/BGkw+AGpNGd9atcWg8MmW5vBbpkSGAdvBAnz4D3AS9lVDQs27e4VU/
8Ol94dMXubkqrY3bMlFg2KHBy3P0YgZfPWO1hqFQRQJVTuGPAPKBo202+wgUayabZkDLoN7hmdgb
T5on8DGSk6dtplH8xfduNw0EkA3uOZot5/uVjLNIC+i5GguCGdCISagHJWeaZx++VuKKQf1la0oy
lIjYc86vYsrWZ72rYKzrfntZm3fKBfKhc2a2q+Py7HRYK0KdAC1O3UzsQG3TGiIXQ5/jTIHz5n5b
0vBsXgcBeOIPKBU0bXse4QALge6DLd265DPdXIiLGaSuTe9vqnlOp6W11whtL83U8Qn32azd2tcd
LZPI4cTqMW55eNhFbRqKxshEVFOpNiZY31n0XGK86DS3ttC52LaCe7E5STRkw6/2B3BVDP9HvhWr
rYQBmzLZJwRC6D2wXln4aBKn4aFMuUvs5yOguJktrOFe5TP/kJX3vwcjuf/YiVeB1c+uZsW4m0kg
W6JDTe1kMdTiGhPhQC5s374/P2V4IP0sJkK4X6E0GVh1WSmfoWPfNi/xI6Zi5WI2lmrBE2boJqF3
T+yKfnU0wehcyaBL47TNNeQOZYxJHhMu1jmm9iSavciqqkvesmU5euli7vqR35qVZvpqm8+Y+TL4
LaPDn71GMqPfLIw4vpYmtyeqCriGEQ8ooZWz9w/d7u3GWOL+NOPDhcccUcsTmtRsF7SmQMZUJ8GK
YsXskb1Rta+qrvX1USUUr1TMXkRHm2HSFL0VQGpr4etChpBgwLpM6ChL3e4OLZJUu/h0x1/FN2Mh
f0BxlfAsiOeN+iAECTu8+o43ApGcQXtgqlyM7ztsm6lX5TW1WmB+DKzIawYrIALk/iqjfz4HQHuJ
bJYK38h044Y8OQ62M8MlP4zFgDgUSWNmD15x34ZTFGFc5yQX1gMKeyx4oGaq4Ao6sk7o6XVoRk/2
sQj0MZNXtyYRcEJh6XeQxtFXzJGDbaow0J4V6/6GtcFvR8MI9m7mNkMgOaDIURkJ9Zt7lArVDtWC
zCbBCiCFS09JjOhCbAnRKjcG+lzbzWcVcyGtlRx/4GxI9a4nL1dk/MLBogKwkF9lv5q4qtN61DId
Jj9iESVCYlcHatv/2o9Pwhwom9e8yM8+dSoEylarzXZlNMNueX4mB81IGBpecA8F6wKyJQ1zzstF
4VTxTf39OErRD3G0xFrQ8b49gypbTK/umyrGIrPGbvepy3M2QFrofTZBes/viJxFYqSAK/vMASWu
FzNR7alWZjgfcIVhyDupAGubP4KQKCN3DManzTBaOkNnFRwvHUdYEXCJNNUvvWi6bjhVaA8lgzua
gh52f8C4YvQukA5b/ECYI4ss4eiyi+eoI/UnNxNnTBpLaUuoBO4R1GEqaMbzzZNSTYgGoUuVNooB
SxG1XIO5EgVMoB0MJx9J8DcLWjU7Ocse2Dc496o6XOCcvHgc4Sr+RzTs863nnM+wMPLBUEnEd/WQ
x+xUKRC+8bQQyKlaRuM3vsKD1WQYX2J7ahE4Uk4v/rotHQ1VcqqXhflz4xzJvY1jLB16EkAK7dFz
wT35wJpMEwLHWFBIJAsgSJtK0feUElmtK+Dt6jjliMF9QXBckeHwr2tE1vc0kP3ukqa4lhXidXtC
Qndioa/zRlJ/Xuh80QJ3zYaMJbVVtr7dE/O+cl0o9AWBD/KDDC+x/6/F9OedNXXuRvx6utVg1QEI
qnPsnMd/SMMqq5Xon1UGFXdlEz6gDfdbHiPd52aP8RB4Fd59e4Z0exEbzmwQEpo0phgxuLxcYeeJ
QfTQRzPwa7A5+q1x/nxwvK3jOhOgL75qhKTD8OLIsAufbsdxRr/MF1r/F1lt2lWiBtTrTuNaq8me
7VdkmmCQy4R+mEWqsxf8B0y+rRjtXdzma7c1DoAwYSVke5b9kbnep8Wr/L54S/Io3x/BRL3QvC55
paC5rbIZ6OY+WcZmrh9eTeXeqATqeEJo7PmSh68AdeIZ8OYt6j2ygL3aqB4XhyRHFKm3f5SvDJRW
qlbqI5aKpp2xezFZ8zWIRnxG/Mr6w3pokBoxHXGonpm5ycwOcmXM8T7TNVeK+V6IZn4375QT8SMt
iWmIVsvIlKSYwaHEHTItk+PKLoFOxNiE3z4+nQ5Y9098YRrl8yoVDvIqSdDqRoygfX9XY9cuL5Ov
qXoMHyP7CJWrIAK0g1M9KZJ02KEyjs1sEyye6xgUvPgj868bK72PC+ymIkkfo9aXywLlUCccxkTG
fKfmRF1fQegjMbWdEHcudxA0pVxsgCoqt4CaZwNe4/9QVNr+BD5zZYeu64v7c+ArYL4DF4TveyTl
164Y2BxatePhBuHdvm5P19TE7hFskwSBvKCjG52+6ypoFGPxpWSuiELIEKnXzVEupzWOPGRKLq92
hgKvgynK2Lk+oUAPDnN3shfVETLL9XhagcOIsY9n/nbvuJhEg14QBDp+isF0RCg+mmoVBZV14UOA
BnMUdHbF9S0vD2583mQevGC7ef7LtUoA1pP2W88rqcP1o58n5ZnZGtzZXGcSFO4fk/+kuhXuzIx3
EFJinOo4ONiAwQ4ssRJWMgQmwqqTsDFIA80Ax5lhxkszGnpPQJ7soORLZccfM2/9tOJDv8V1pJtN
h7xmg0MlBPmJpxA6LD365AYX/7hOYWTzpA0+uQUZZLIzsXD2H0vV7vJw07LbrAiQTZsoICojC/ZU
gjDWKqxsewyjCVIEb2w9hF43A8eiAtj0pOQX9vmM1i93PxJzh4MqW5wnHt7Igh+dOrX8hPLVJ/4V
AO/3+507EyDiobcaNVXxCB+e4pfxFzNyjiBcTzfXIUhAGcLikPK8yFP3nwhAqpH7lvEKkf0vmGcK
9NrzEugPJxyQR7nJw6CdpYBgC0Hx5qH8zjgm8Dqf2iXbW7CSqfDiYCYvtFZzDEiBBT3CxFLdJpMF
65jQEPQl4QAGMPSRZ1vBb4xa4QA1NchoRIfr/gbXOLFapLXGPGWnuabUdEX2swpRj/9fkfYysiNF
oa1IQx53jzgTtMaPEiBa9mnewPjGemHfmbzjyaCoMsDyNyoAahIaxHFIPwKHnx0lPDB4JoyouEw9
Pmr1hU3yn6hTMV0gSdqLk7a4FgeoHix73c4BH1jyjNtaPaWbhVWI97a4NJsdRJm9TfLSbmviswS/
YZH7NjVyAQJisFys/PpLTqrJ8Qb4khzoP96WczTVmGAwlf75OWzHZ3vbi1wIlbnjC5G9Nen4uopI
4AhJqhOAC97WSZWx+R2mSZFxeE7oBRG0FCW92GXra+F5WYWYlQ7JrPvmLKIgv+E61syzAiHYgHWS
EsgDB8+h+UfFyGAmjqxLjSM3CJRAGI19uJxVQPcSxaWBBU0ONeKHSRkb7bacbO5Mr1HWafObKjHr
KFSOVLuNCrBvfZnZMKOuwkJTYv3SAW93MjqF9KV3rqz4qlmUpt5II3Y6xqomIBFkNuMley3YZiOT
b1kIRRiRBsOcfcpdTguDX5OHMK9jO6KR1Uv5VJIa+5lBTm+BDz3WdXasoKEGyRKUorxof9OfjjWv
ZbkdHYHGca9oGXNnrJa2kJKFdiMtWQwLBTiVaLQwYU8XjGAuKNsZIepHtWg+KFrShqvYEPTR1/th
kT6NClsE3aHxKW8PbQI0VpsFm562D/ai7COlW6VqL4zOZpcZtQ7fah+yh20pXt/kCrluWIJr6acI
4K5pu5t7/yAAM5ARKZoduABFaS1po48n8owBLuS+r90aUMnKibDNtH2zTr/DvCFeW2hTsSayuseg
z8jOO5Y265aIIvwfRj2p8vD9p/+adpiQw8lNdB7KcBZQZYuNj4tYYvQM2M3da8/3RsplcYlB6ak7
8D4iywZzpHgfg1wGnTgmqIJXeCYvrOh7HhQpdtPqjP0B+NqdbimTY967JUWiSz3wxZMkEkyLuVDE
+HlNc/9A6+DcFzziwVF9mRFtqa5BfSM5kSedBdR/NB1QEx8kaD7KdzrN/PQPE9yUgWCrwALL0CjC
IuAPBlkbK5zYpM1cmn7+p1KMY4RgNo687ldUyOqDhkfrmo6PdE5E9OjxjQRClPUojWF++FJgku/R
ls/RPI3zGskY/U2guj+1DHKWyNoXLfBA6/7lnmuSWcw+g8OZN8PLlaVqJEflsKlkWMslxrOfeUhS
O87YsjSALfWQUa4k0aXCLAoVqODGRNYqLGiuum+XzoYTC4bRcPWLI+1AL7xZDeBQYhku2ujSt0OZ
ktFJIdCV1QQuOeSj36nrI+MXs/3LMq6PBHBkwPL9t/5AZmzXwVNixyOYJAQX8DnW9xtAUps+5Heu
WoW6U/LBvjsUoe6+McEYWJ07WZKZv6CVVa9Ixmg3hRhKA6XUZXeU1Ada3kJ4W8gsQhbtClabBl/V
scy2R8vsxzqnYypptMoXctL/ucsmgRqXBST6WjTXzCqkYT/RHtct0DZYYwH1VGgvPdNbbk7PsBJI
w4WNOzCYV60mXXL37RDJt3HeTrsX0+DQDr6DHnflMHyy5NwYC13pRKs7FAXJJGkfOP5VZ6OHI75c
GPCrenjDNpPD2C6h2XyHWHdRZakFmfuc6pyIuGfqeAjT2RrQLgNb73mZrI7wk9O/jjChGygiMidG
LQE2PI9YB3smMXA1DP5zApXdKDfEGqjQ8YkHpEvrOEG4fx+kKG9XxRm43P4JhRftiyb6l4mTgflz
Ih69HVa1cWWfNfRMeLI/MMAIdN7p72yvUT5Gt7gW2VfALqbsKmvkqXSuMFFzz9hEaneeK2GnWfkS
z1BrCU8XRoxcxwgqWff+1pD0xGJIrNgwVgF4uV4v827PI8wF+PrENwDX6Ot72TFFrPkVrbqw5nMf
ZDE+rpaIyVSpDZ4hoXnFoFnIDa95bj9XH/jwApvptyD/1KPUi84zfDAiqYuLJYA0JMYE9/7EapdV
a3jU0eigmSH+s3cooHBw+IDmKrjZp/ZUAKZm6zZWSC/utON01G04IPy66JhWoVrx6z3iiXediqas
Kd0JPdyNLs22IOrE+M0vAPE/vwuo3413aQgL3JjtKRO1dzBC88j2Aqf/ew77WcY9kuGwqE0QxLd/
8EO7/OhE7gwteDo/y+YS41lIzhgzLUbV4gb1MaoVyL01V/Ar5mB7+JG8agyK04dt3pOSG064akI8
RfeF9uGVjyhWLx+4VnqFn25k9xQ/13Hb0/kuDF97G3Q2i1nXOISkeE40GJ+lcoVz9215ruA+3c0p
4RnpvWWhA4BVqiHd0rAstnCWRHngKvEKB9UJkCWpN25MBg9iI7tBte/f2PiAypZIv2MBF5yjX0Sp
NcbyKVNApCQiZaqbk2flDWZMGTIdGaChOTX5iQ/UihA5L1dFTVoWCaOITrU0aYxF9KVLxD/I1s5K
WoZm6d1Oad+djQtoIJqrTsozdDR60TzXokZsP7Ode+QWNegpFhrnTN2lMmPjR4nfwHZVzQD2iKv5
r5Ab4GKIRn1Rcv+e4LWt3izTU/lZly7LAZ2WjEU8gA9YwYeCG1XYHP+6WeH+ZB62aC9u+YS2vaMg
QESNrM4qzDwd7Sexp1HwLUNq4qaDdQJWFiC+U7WX3b63vgi1NowRACU4q2iAKSg+iAZcNagOYuhs
gI14ef5kT1WDGAzNqqUptbudc8GPlK2kUV24ybTgnBOHnfOwmS2NCuOcTmjkXLbXKaN0d5AVIpgZ
ilmL1f8+SH6ZRIgE2pcGezS+67aK+NWuphbE0Gbdy0pmv3rMuuKBwPlkxj2LDB7l6QmZe73OrluM
AUFuftMkJYP+lTJjzA5ahi1Tk6fxaCleXZNusB0RXcVplA3toiGyM6sygbzwP944aDSqm8Zslt4e
prShmXreHZoIJqtxqeIQlgtu8m53In3Rjj6ScASWtILsEGMEBxyG725efoje+fo5c57PvLaC15JH
A9+SSj4x4q/VYayIGbnxwTSYalJVFdfQLgqPhe6n3oVjPNuzZW1XU0U2m0yCl84s96sQ00RYi3cM
4AyyYNNjbcHHd9Tw/YpX8OE7hMShkJdnfeM7jKCPO1KsxQOQ9JIO4TonQqYChVmTyga+Me9sqcTj
W8GqquJv4Y7p7EtmSp1/4zdYFMLfTzQiwcEapeF7rcYeH6uyNdkFNwf3o+j4JPsJDX7Opj4vBZ6d
P+UEdfGqpc5nH32+iK+jnBCUpnfCPzE1HCxhnfeiJTY3tNrKYv0ssPiGbLRExtKKthZHDVtpaiFP
CnILF1Y5v0Mp85IbuWY+j+/lSG2bJoqIwX+xdb6xqxNp/yFn/R/bPNxnIzhYPX28tYJKU5a4R1zn
J1YZnwhXR104Y+b9A5wWmeDrwdfM+o7jFzvo3pF9yd+QcV9sR0dCffkNiRLxSXL64ID4EhL9cX8e
3fILXQEpwciXcaCR36R72P80KW8DgGlhTK4TgawwrJV5WRWSE9bFMF9UhdWyC48mJNnfNeZQ/Lq8
DLwdd9ewMb9uhamzFw5xogd3jK1Yzxg4CThGNIov0kL7a2S8Ch3m/ciIq9COi47eewI4KfTPcn4m
6P+kmA7ZNK8vpMqE8dWUyviuc2zOn3YjC8mYjb67mx+5xPYsyXut7Bw14r5xMlG/sNmCEFAPAq2n
uPdo5/8iCE0yIvkjZSZZcRmmQbkUYbz6CFxB0Ybh7fFQjrp4wSyfvxPZkchZeRzc3FXN8CbXWB0e
mtL8yEQqKadQ32JCyznGv9kVazynWehqAk8tlHKTkC5/Hk8gn08mgpg5FGQ+9HXl5ZjckQ2KsR3f
Po7cQMqEmTWLWgCfacz6FVNHrXI/sxDyDhpM3yqw66AlfnLaDW0pE1A/B5tUcU2mgVZkSruFKfY6
zmRUiuexJg+jkyjO0HEmOU9DztyLDYduLx+5ZlE7gcOX4lo+JdeUg6FVVyMke5qRXS9TgtsGBjpR
iaSB89jFR2+M7JIXLa5LHaYW2fvxHjE8JXRMfmaZyj6g+7B9ZPOSBEvNr0LAGOtfZNW7o7IHsryu
HJuEaLz9kxVL5Nxv3q/q442KNyRyCrVHXg62Dpz065vXmWIHoYllrNH+h/m5K+83zGiLXvNxmgNF
N9IcvNh8+bfIk2PMfHefkCnx0/chMdWakTVh+Eqvhn2gCyK3085Y2Y/gUGVsyuh2tmKlgvWrWwPT
l0TgGEjnkUgSa/z4NiND821rXn440jfF5OQlSib+s0YSSg7jS2BPEJzOufeXrUPbQxllbLqCKRK1
ji6EOXIcLFfCEV6hiCI+WkMArDVtmyjR1wihpMA+WaiIZQXRZ2RfiEvrO+qHGU0vmGInGNuY7x9a
YMsPSkXBRMCRBvsIlH8Y/oebx2yo51QlK5/1JYiIxRgP4yneDFUcPzxw9ocI8LOGP+loYYMN97U+
NQGYvPPcAyAWs2mwqwOMOjbkXa1ryMgvH7SqzmDLV2AiOpx/5vOr6ZcmZP+Wk4Ke9WTwmLD8wAsV
JqM6QwqYW1aFiEGK5yfZ+Ex2ijmeTOGJaQ8U/RMnDSsS3eNhyEoCl+3Kpa7/OzxBoPwRCz64Ns4s
x0jlwZkQu9EyA+ba/btMrlEHFyfw6pkjF1HPuONmp0dhlNbCWswid94Ba0hnS3dysIzEgdZUw2FR
YYtRA5eJV1sE8RnmtHmN5T5kW47Jt7hLCmX4MxPh4BBMUIXieA95B9AwPwjeDVN8b3GUn2PcZFq1
6rZHYjOkIgXwn+3gB1mcBic+COm8wOG25JtP32yiWq9qKVSg1xEXC0UiXaixiHl/E1D7Jz3uudVu
xXx1g+RECyT3zSsgAZuTSYumOniJn8wLh/w7f2YCp1TGbaZdpFxEsTvh9F8ZWbXrcdJ9O4RcV0gv
fT0iLsWcjpellieE+W9y/A5SSObTAhpLR3Yoz5bAeqVJPz1Ex3jZEI7rLOMbFe+8LWVuz5v8CVZ3
iu64UcSw8WUbCMkzGy7B4+QW8SWUM2feLwmvYxwqTSSDnKqUYyxpA3ymwjALQxzxVS4vT+BODGxZ
7JE6aJAcFnpMFVVTdtYGTVA+0cC7+hEcjGFL5P+n9V58H11Fz2Pko9A1rOfII9M4X6+oHBh3CyoW
KLoC3F1T548IRv0R8Vf0QEmBMJvgDJ9TW+7XeBR4WkM0sRuVe2KEBG1uaQ09o8HXmbeII8vBhzyG
Ptd/rExMxytyQ+eqNp2C2rzMorG2zGUd1JCPuCZw0itbekxurXFW7NEdHvRe7JUY+B8ihVRZ2jHP
U1pVXxEclWXjm1+ndyKsF7FCgVgobSGRBeoEdywHZfYQMGj9CDPNCDunD0johYuO0KOION+/wBDp
mswOmx/imsfp93u9DNIgB2obmAitGpqpf50j7CME2KIbkFAsIPdT7CT+veCgWw4iw8LD3ZNQ/mpp
sBK6sI2zeFkYIAWC9PWJ40hCNsnibMpjxk7UfEyfiGur/RGG8rRBK/ZMHYHmKBjlGQzapxiwXsqn
VPHWjf5hRx+5ap8Na4jLD/62xnTKxDlQsK6RbiFW6q/2uKQq6aIYh3Y1F9mg9CnhoTI3+o4RSvcw
ZKXZhIAy0LG/DTSsX+75S/WCPyGR2N5KysP6mbW4Erw6IPfoMvLaS/lGrqRiyj2Hs3oMbnfgl/nz
jI+7+2Y7MmkgS5W0wNXD5ItfkJ9ZzD6iB5N7OxjmAqIc/Xu67aznRYitGIKN+N7DG/SANo54UXoz
44upbgFYYLbEXb4U0ii7S58iC5DE8fXvmgvqeq0zPv01QTQBs7lIsoz2FJqzYZkB6jESHLP1ga0+
4PJ9oPGiQFUxF1IFAbLdVV/68X9PBGFBj2qll9tl6YUrh5jq+Vl9qIO/F7BzFnwAymWzwu5umwIA
OS+XDrsmAx3uxd9DslkqWexdN7WOahImeWSGBBRDUkKvA7xSvavy54GguteaNzbpx+CBJgDB7yMl
PDTf6ABnpPHZkpem3u1wouhGN2lvwMv7P9teCa0EpcKiMFtJNkBmGvwXr4bYUGynSuUyVzhL6aHO
jvkroQIj27m408JhoDIVWixZA4W1wn/JCyxgCwupN26e3hkjxxEmje+Q2b13zsyP9RvdhiAcZS+4
kRomdUyHtMrNEWG0zkvGo9XiixZPQ60ZeH+hqsIo0Fs5fkBkz4Zfx7sVb4RUsEvflPIiJHI3DCAL
cuEpZ3hlZ9luZ1pfGLSyiRSDF0gCB+hKBF/BvHGcQx1qErKDs1L6dSypEbFISU9OzCeyr5kO5SDu
riLxMdHbbM7iQxuBdrzhgeJve9UmcrBJAzbKrSdjvf20ZbWxIpdtIoGF5h+e1FzhepW9ou/kpxTw
kxHzSoR66VLSJV8C8+70y1ng4D8Da3BzP76M2/SIYj8633ladK7Cgatbx60GmLp4443uvOHfWgMD
yEdjQ7ksUjW22u0VZfuBIHZDURb10lBiqHtMofpIfjpKWUpoQfUl1baV2AfizGt857i2YkLFCn1/
q3YVCnOI9xr176j3kENx+V+s07kkcDs59RycE/19pN0A2K3lFXV3kCfedrLEjSabqK6UAU0vrTGK
8UurQAWcZTydCPIeiowQuhd7Y2lDlK2zv9IjFyitcnzgYxMygM4PNSQ3Q9VlfQKhFpiM7FoRoW6g
XQL46Il3NXpt5sx/EejGHX8e2Pt14X768F5agnlA7QjIayFCzua2tDG8gkjxa/rfLkRjB4Tpx4i3
wfvXSDZ/D6KgK+n2kafVZp8AttEjwmg0hWY2SEBhPSpjB3cNrzQXnxPV1qNZ+FD0kfD3hQIEFcq/
DFH0H++oaTxuXF3mygB14SHUv9Q7suhzOh6XvR6r3CLsUNHLhlrf3uxUlqEduwVZXmExOsWwRGIE
V0jwIhsR2ugLaWrrWI75lP7sGAjVy5tjBsr+xEBJuMdyE5uJfHoGcc2xARUKkwRLNNWSXHS8z9yE
GmD2l13QOZTwFbG0Ln3RfVmjBY1TDt896XddCBz2wqREgdKoLnBuMcdcN/+gfGmM6xwj+pSJOb8D
xHAwTFNGskaM2F1Mu+3idCO+F1HBq0GuI5IWtp8Fcq2MmQoobImG6ICG4MMhPZ94tsWZkSobJCWa
7gxmhLB0iZ6S43MMhy+joOo5k4Yid1NXLBSGeKarLZWLfGpIZM3dA6G9IPHMjxkkzyMjUATHMkv7
hRBFk+s6skRVKkTZ55uPlkKXbMqwuxkn5P9FZTZMalqoeeCYhYneUSAlqvMEe0gbEG1PNs17Let0
saeL/nJOEtYOxUVQ46QDjA1kBGcbaHJ/ymrT6wwF8RPX4TFE0EVUNNrdGTnlQcRrI2qo8D/+Tkhg
cyFIswUZ2MzgQkFhk/WyjLOBHKnm/fzEsmEUnfBW6iCffhz5TyOzDeHHPSkEWkMuKRaNI11/ikZ+
dLnDYBfhYWnC7CY5Q0CZxTIZDGaewFf8Hr0EMgpSvzaJ5nXeVcGnUtPv6EA/EgjBYTKnI/GTkZUO
58H28DOJQbsROJ/8jlWw8vADiJJ4uKVt0CaWlSYM/pHG/XsLlSdWXi2LfOnZD8QfkxBWrpyQ3TJX
aiHgNHYFdalsk3LEGpn8tbP1BBs/7XQPrG81XXapFHDDyeCJj4Enex6gC6tTblxIGdgEaN4aeySt
0ikRuMtBXu+yqblF3rRQb2XsuneSswvVfsTjWX/JhyOrjvBvvzx0tPfrCjVl9uxJq3v17CjViILS
8yXh0BbTZ83rbJTkdX0G3docrHyCRy4TXP88tlyo04A12zkGIlHeR6/fIBucEWjO8kGwzw97lNtA
mwnsihFDtEVTv4/WkYStI66sTDJOKIonJ7WqNbrXYw6rEiqvCoQJGOHKN3RLPIuy1csL1AEXEyV/
9hrOEz+IgibCWd5Wmigp7koLkZQATcJWQBfZCOGbHdpWedktfepZjnuW9TYI7QC143OF8JqhzZdD
BkjV2vJZx9zQiwhm+RfSwOSt4pTV6xdbDymgnFIVpXq5qu6CBz1vNrD+OaeD46MNRTY+EILy73mM
W5uaTG/YZf+vPC18+snbptbMYawNNmeJEl0q4AsmsEJJQebdBzQhBiI1wXZXCTeWyp+4vuUaRRAz
IxlD9DxXxJmvceVpwVUMo6defIsUbmth8ppinZNno60EqM1qAFUzWZpj4DSs+uKz/wmfQCL2zzTY
9VDQ7PtZP8O2TGumcur5emIOwAMIVPcdHUYDO79momJSQ21zprrZ19SaRkwnpYvnsqXytuOEvQ90
KuE86QiFLOe9K3wx3TMMVEl92UkLX/VFHbfjZKXsvrRBvz0fRzDyvU3qA2FaYcsMqEgsbRJK9V9P
enNh36ZZub2J5FsbD6gHR3fmCUNYrlx96XfgD0+qgG2aWg5FESsVI3x5uaBABCSj2OVkTBd9aaXV
uNuhr7DNETDcd1LshCNHZhT4OLjyFWBhXQFvq0rGi9RXH5a5bkH/S7LuAR/OaRFqQWTKnXoqmvy0
Nl7ETJ1sOnwTzKVtoys/RZTIJ96yrQOcB/LTcwlavJmVTA6KDGTNDXrvnXdImBRWWnHdpD/Qzfqw
l9chuDJlHxQkqBJgbdQ/PYXq2FCw92sz9RIJ4KL07ewANRNhaW4fZO4ayymdv1i+hkGbpg+eH3QL
O9TrjNuVAssn7jq6uIvlYL3k357Rc2xDHgm/vZu7rFANKyxzeMNj9ZIrjmFvUH6KDnVSAZA/Z27q
xFn2VePjyHSl7I+3/wATvYNHgC629/+zw2WuMGRdv6MR0YEff24AG8/HROey4XG0agRoAH9Gc3Ph
rQNq7UkhtDaRJpGmEUoALsZKx2lupF4NCab6kvv1JcGFHtiaoHOapXM15v6cU690f+DK0KnvSzZG
mhlHYb1TdexOT3q51IzJxZVKIvEV7EasIAzzn0rrkN6K5a0qixuveJDSInKBGkugH61DX11HyIo9
RCXAE0tnWkA4snKK3TEszbIY14wZJwLbDjs1ZIrwLwAsaFey4eVz+gZVxQ71yL94LRECRbQ5PTUD
Pm7hCzHPH4rgPOsFG0XtimYMpzrcaL6R5uUqvVvUne1JhvI0sU03uSI+dPaOERlZX1hq7zmAb+SA
QZBuQCZw/395wtHR2xETmXD3OlQ9lipSZ3qf7cQOymymi/KSHmMbErad9aYLztkc5aMvPSvpUT3A
yEmOvrKoNMBbOpDgozR3Jbvw0FgnlWMzeJZ04Hs5gg+R8NhWQoJFunBnA0yJ4mGc2XrYXwYx+GlU
W2dwAYQjJnVaj9se0SMZqBEA0ZhxOCPuoJt3uOEo6Mul+WqdVZKGKyk5+CxkI/HsFdb1gHpjes/3
vJvdJi3aU1NEpqrNoq9N7WmAJDhHbHI4mEs8hiprecHZrM4sxePGURd4ix3KWs0yzd1TfgXVpPjv
/J891RpQSmkKVyvNUvBTDqhq1+QdaOpGbP0yxqi4okIoFhvc5SD7v7xEdHGkkS8GeIp2UYbBWm9i
pAqWK/PHbrx/2eGSOSvqS39A2ufmvPS93H+S1CA/YELuCsO97bTquSJmtUWdlzSHGAkA1Clh02pD
n7xAqF5YVf6ZPCxdO2Hpx8q0IhM8NIobS5xfl1ONd0gB2za5N9JiUt0zrlXmxT+Xsc2RlbgOO8uS
b3I8r4e9wgVNfxHsOdydUX06EWvPqid/uC7FT/NIDtX4NT+NZ4u5BAa74flY4Ouc+MoPrrOt0Z2G
MwGJ4ygCH/YwD2TVc8DeUXeorjrlhCQQmEPfiu5VbTuz/SHH9xsitUUqfIKJvrU6iXwGG5B/TbQy
fB3T6BGFDP48u/x+7BoVXb9twPfdcoWMPZQfhadiS4H/f6+5W9Z2pboU9LNYlXx4xA/1Oi5j6OHM
p97tHPm5WsoVQJzW0nrNdnxyWDCbVkaANuXoFSZE+ykfjohoMuohKVp8lcyvWle6GfuDr7qPFkR7
UK0CcxSKJB8g1jkgreXZCKXl4rCicgW4aqO3RuuOX6Uouttsw3hkwR1J89HaCBffN5ixFbW4u/lI
1NQr6MegTYkR/lZJErVVpbRkAvADsF9L0rdMAau6KRGP+0aX0s3ukUTSFKpfFDtTYlmkp/Urey77
aj4eYKTRXo1fMmP9FQyhQn44VQMHwhWGBkzq3B4vRieSZTwBrDsNvX4SaFvzV8Oql7Uy2x4/+fK2
tao/8zLvrPJ6iPtDPKM0zCOR7rDifJHqv9jV99p0upUbxG3ALAhk7LY8DEBRwTHZ0G2CcxeR1+Wm
3Xr2Tmyj/QpznlDKk1C4pVAmAtS1NJARkoCQJEaRgodT/SX7+xrOxOhrECHvMus3Gol4ABZo+z4s
zjDuni6hxhmRLwqS6Yg6Zd3Nkeri4pRSZjUhoeBwZHQDfEYwMyLulXE7x8V7I11mT0YPUqBLl3Y0
k+TlOwYpiwRGSmvoDu6OyTtIS1J2CbKIyo4y4xip40y/HmJGhOj2WLvfEyFBUOoJTYKdZkrBXmwU
IBigrYQF2PtWqrtlaImhqQHWA4PlJaeuWdU24Sg+zilQvoVHnzgtamJG4YIXX6lgYciN5zIYTHan
uGgLDKFXBkjgYE0MwIGYEscC1C9uZRdsK99vMHdu55wZRMAwAbxvWDcmdbD8bllwTPvfm0ScXHKJ
fxPivtdqF0ywHYv2LSF+HN1LKm/m/iHqvuGl1unoPlZY/Bbn3sYfhKBxk5OTVpkrc1Dc+SG1pYHI
2Ny4shQBbUceJ2BqZihjTqcFLvMf29jqnwx1vi4GRzZ26GRwQoP+pbxvllVN20qCRVhbPnC0E8hp
56xOoi5oIHe9Y0ZYNEGo3coBnGcar5KKiFrNMPh37emeVBFi7ZylwCkgMrEk0HLTC/wuwmfDj9wr
Rk/zs96ee+YpaGVeRjDsmeJHA6uIJh/y568EsNymz4Rmypb6uiUdDn5RuFSv91Cs7CAC+TGFVJB6
VYfq+4f50aLzd+P8GE+A5NID6uxMGytVUOfKp9lrYVLBHxnDNt9iCsB1PF9bCu8kCCnAVuCMhDRZ
xgRqfIwp7npZ+glpZ6xeDKJt/Y7GTyrdquPFWmTLcIt2mO9n5uYTTWeBhMvdB4wYHw94qTuKqolh
W53G9ldgyu+PthyvbkuxzgmM1MzjAl5OPruiCuj/TC3P4g9zBBcuefly/Aa6BgufuBCkOvE1Qb8r
qWbaFciof/yBR1DQXTdlzy5O7Kliljytsk/nxg5E5k60tZRqVHj40LZdB7/oRPmNIIA5caei8Xkq
LWL7RjAWknCOuGZfEtm6CJ9i3BssMnE/ye3ird93g/OAAZ0WaByBejXUSbkC8IhAJ5gWWuGT2dAg
ouyZBwggatTJezgHvZh+2u2kYtVLalmXR4iFlOYLmF0hr71uLM4vDJUTZ6RibCMWFoi50AIEDvCH
sViUpQSvla4tz0EeGdll7SuOTYEV2unDsircVQsYOBV6MF0EBUQIwNUGsT2ibQOzmTie8JGNn99D
WvDe0FMLvhBYqCV42yCDDUBlZvHOOAjqA4N2ERE1REbiEfJtRt/3v/j1iM9a9oVvDjnurRwm2SID
ntPF7ilJNJJKkY7pFInt+l9FvfKg6ipVB0uscnU730wg1LkCs+35EWKJP4cXwQV1+d1ZtyrtQZbE
C//DpGnsRkABW/5SfQIVeffmWYHaHOfMUIo6BXo4ziWf9I35C19Cb0RIyx7P7DHvrJfa3hkOadZJ
Sprg75cHmbuKWoonIV3QUdxxeJ+wpcvZvi2f3dNVKwOYI19puk/2C0UoN9miokWR2ik/MNs4/2UP
USUXLAH1WHJs9/5jieye1HG0hZx/QujVc71SFmSV814Le0wOVEck+ldpZdniW15MvHX2Aetrxc+R
h5pAlOT2kwBZqfRFYDlmcM54GYo3HV9haQjE/Jhera8quBgvASgvXhQvjy9LgtuuRxzN/SBilTwP
JGAPfT0+oDBCn2zqXekBBRTmX4PRslz5wKUuS0YU2BGV4HF178SpgCKNQy/b2xCbAoff1JWcByhH
+HQ/tvuRy3Y61xp/wgGx09vEPG0WTxGhy+pPXw226fE0M+mZgxhoP7flm8OscZIPbYZ4pptb1SfZ
u6BihwGp0NudmLehjV0FZjZXjiCEVQToyu2FVXVzSCrOmgwb+b9wO98YbJhO2PZZz8B/vrvLrUEK
IVyYevk1lWKxlhvN8mMblZ2zBW2JQfzIDwz+bRiWhGDUmMa4z5UK5N7vm0fYaI5kTl9iOQExDsCG
jDpzOrVEj+uXeNVA8qUrpGV49IWOsa9iWqXUEyLGReUdmNmtomee3KWPwZV4mZta8aKF9UI8sLrr
q1vR4pcvZIn6VQNGYiIQU7w6ODPXn1alzFO+v9LaQxwAg/HIaoM5CRKM28j/+Htuudg3t9KZi/hZ
cSN9fNuT1ty/aITElIPpGn2+186q1JtWVWqdXwXDgvnm1mkrkBY+yHFNU4AFan/hv2Lqr6Vea9sG
b9680ww/m5iS3Vu2gd1IYPXDno/rLtz4TdA+ALJ4QLRDbM+noqhJulJeLDrab8j70KErphjLf2wr
bg4vK9saFb2FZstobjxWnyRVdmYql2RNw+vCEHNa00DAXgIkgstiZCkAatXKjwpEhm9TF0XZEmM+
dBncuOOcb+lVKgXHVjf7dtFlD7QnC+2RB2VZuR1lm375ZKPrzvNkAQh0y68pQjIEeYJiw2q1pq1x
PzR1A9nldCJzVdVLyrHVCxdzwJbjxrtU2xmSjSFmyI5M1S/Fz2/2hexRVmqnAEsBCehZpCou5Y5l
N9cHQv6fLA9g7yiYSgp6Nu7rP02vJ45ld/vojtmqsSs3oqdc2HQkGPet3sLH1OIUlwT08tIUVvey
4wOD0KyqhAWQjfaGcPHkohHoOKnbZbLUw2haen9/4EmUNhHNP2Ni8pru4l1H9f4vkzsBkc2hGiB8
KGnYvtIylO8HOJZ5KUPdkLwUZPVPZlFdnEl+sYX3jZnKDyxpNXNvo4QHRcrneKs912GGpT7RoSrL
7zwdvQTX4JCbSabsYJcT/R1Tv51hWuo8AvUAehGqDKVMlzGYkBSjv62ByiQkS5cUDEx3jRgVtSHC
dQD6p0PhdI7jI5eA4afxAN4FTecEfvtjVqf/XsszdL4DcR+YV5mhAVBIqOLx+nUyeFyhpV++Vftc
f0sPCMIn5dXIHwHZ8ra2AHV2n6y+QwCSVwE6mrRjC2P7DRYfC0f3Sd+SSFi55ic+ju+zRC0xzEX0
kPOHK/NYDbAZwwDe0bO/IY7Yo4lJ77gw8v3u9M3GUD//1AqpMNxBqeMYT75dGHr9dqDhAcSdVr8q
5qIM5eit+1V0Q7XwpZPv8li4nww1p5xSABlKTuZD1ymJZ2IK9cypdG2v8sXWeNveD1OjilqsIVhr
uZ39Dr2W/ly+DexBIiCeO7EMv69NVKZTI83mPdh2kg1P7CV8RbKl0THgFTit3iGkVLbEakacFgJ/
JZ0qLHVAlB2REahNAZ2KlJAn7+3/Kh3NROS6Gx8LAPOd1+8u4IBH1auMwPMMYSfqmyP7TnTBcaCP
OydOWfELmqhlSTUdGLcA3tMTIQFrVU1JCsakHkyGmfWeTyiPr4ICyq26QaLNFYjaFg8diyfFrAet
ge12MUPFFvx6wbS/vZrTSu+kqHBJzzvsk05uDV4jwg0UFgMtm2vSSG7bQW3gVIvRVswRWcRWanTQ
Jco/R0bl2y2C/96DO7krBgbcoCLax26Q17eisXMnnxJ4LzjfgzQTMEmByXi3DBsw7bmSs3Cq6Noy
GGqNTcr/4mt+/IeiQs1hATzPrJGlkOmsuupnXO5kHfTK+t6OsV1QxQ5TUHIfXC+j/QUk3Gr2EgRC
UWuJOaMcZmqLIzTEl7YEVDs0Kqbd6y2oukvdu2MPTrBI30JlJzFDf3MZps+S3Y+ENXGx62JLI0/j
1moF/D8Mi7XOl2oaJkNZACCniIabhMQXMAUgBwGLwz0T+Cw0Xchdb3mchgYbqpyCXWifE0ROze+g
CYpBHeHxj9TWGqrSroLoTX5idGsqGK/zYVrLUTxZyRjbosOCySpafRzFnloT3Xz8twLGe8pjJ+Cv
wK+uFcuUPZaMezZvf6/PZi8sVoxeAgKdnP469abL6r4VIB8j1zLmKmYrCP6ceR5buBzzsU+SLzoh
TZa1XCDFKSt2qtGTZEmX3qHVMa1zxkwTEAtUTEhA0yZFiji9n0mSIHVvqJSc8XN2Z5ziY0A2Becc
zhXn1EpsE+t3US44WZIYtl8GyK+1hFCNnrswFMzY1r9YZHWzHXOEp2P4CxCxV6Nws2VI/WFf1S3A
gyGfU5yldh1A3gvMpA0Ock4Wc/BDSL1cMvg2OwwgsPPuaQANBa/ZfnX+TCegdIvbATzHiBvHdrz7
pFyd/6I4/5RX/iaRWgmYQgqbPWRPvYA2fcV0wNCAlGs+MZ4lXiydP3QpmaVPCvlNPaOQk1ZhGS83
/qNol+Et9OKPyzjcc9R9VxujwtPe+O+Ro1D82E0jWpuK/OZCvhqbZVGFqC4Yw9SOFxjYtShM57he
3i66n4FApO+URqzsN5Li2Hex1XFZPsKnLFN4Fb+p37ne8I0JefU/yyewoovvoWOQ5u714Qy6CCRr
Jg0p+T8TpogcnQDrYMcEsGF0oOeJWtdbpZX3pAVNnPzHvBtgOzt7AZoblNNKj1GAkUjd8Nn58p0M
O9asC88EiphpyIT2mOMJhBbg4m0mKQasQZLVstosfK0ZdJOYSMPy+2NONP79p/PmMJSsNDVhsTnA
2DNYzrinkNSabZAJa/lVTw6lkyRQmnkIqHpoL8EwPTZbnbKQDnjJrD5FDw14VQyUpI95WlnJx0Ib
czMIzdBieWjwuKYVCjQuieVfIzCjUId/sD2sDAJvQYiqA1XuE3CVZBQJfGZdnBw2XGJyZyD9mhLy
2uac5nJbP3AIZbURHQpZTe4pXhuBR9QFS5SAZXjf5TYvwYsyN74cUudj1oG08ghnZJgaHOGJyTWc
Ox1OJcCjvu+UGS1hFpMhECwStvf4UPJRb5QrgNlXW2EZnKmuAC409A7iUADffvJvouUVf223H0iJ
NNV8FhBJihH+ttz71DAFqNdo+w3TaGMfvYj5/rPzV4/+GsmhwYcMW4nPjNlQ4APYjD00SFIVg0wb
XLLDPP32ZEZeY3m2kNf1b5PL7TN5hpsczDYfoulB18Gtji2lWYaQdaFop2IRv8cXLKyGivN39NOX
PZsXIqdP0miZQjmSdAmJ3ZC3d530A7fVFsIPeP3cMWjcE50ut0HP2C+cT0jiCVPUTvsEDOVtkUkA
y57qYebXG7BK+nNkAdBbVj5p7NXS77rh7DH8WC7nMp6abYD2+ZoXcA/lOzHvVXLOa9lBTadT6/2o
fayffdrpNv4EimGxvrTgyGufmZhgXFAuluk86M1/DdOeV3fZ4lifMbFh/lOF7Z+ocFDKjeR4hLZ2
xHR3n46InksLCYRHs1VgTgl0CvgugmPwqBnzxraxGZz5EPJzgfrjziX1775pJVjQAh6r/isJTcGF
tisUEXi+0tNu8lrh4wVu9Q1v/aFSSRR4sobY+/Bn0ZTgzMP5RGmUhzyodzYq/p85MdZ+mViRAtgS
93kRigcKvXvkpFiOnfdVlNjOVgCF9F0JT16kXesfXlbpZhkOwztJZH/bfW9uF8lMdaMqdFd2TejC
D3pl5bP8izYaW1S+d0GxFy/1uSp8pslEJ94SzgOud6vK38J6+44sgP49H2asXkrHWK+G3lN6uFJ1
exyOFxJeThGW0wll3EserFnShrSODlPbor2h9A1USqN3RxIoGI6y4YFZAE7SVg5n+UYN2fLymn1A
KxutxXG8FttC0cTwJOgnu0Des96tn24l4jHjq8addk/HAKXqaX/0K+ENGZxrN0ghTV3DGPeCyAUm
573OYslTznVSuSp4Joo3mX6uYtPOv+qXVHcEWzFA/E+lTO0OGS6Eq9Qf+LVu8f1DRzCugtqRiiPP
2R4Xqtg3olHDpUgRD67mCSJKf5PHdmScKyIVvu15gzWHAI1vCQsdXkAHjtapwsdak0ijdQ9axf4z
m19Abxry7n7rEVoegBY3drjEsV/D3qVrjXyd2tJ+MQYzlsKW5d66/aNmSOYcVssAAXzXw54vFnJI
E+M59HjWvaeGbHh0k+uwJS8km1sbAIgkJDS+y4W5QtIymsIWFDEylqkKuukAkutpeF4wiCo+ndoQ
cVTT0yGvnxkcb9nV56zxwz6GeOIdtn8tOHCLdA+G+LZ0bBgm+WPftmtcABqIAHIyBYuidupGVVxE
adO7OnSR6TGTIEcfad8rQtMkdc4Es6RjDVgmNiIY3slMHWpYSYQCs2OS4J6VMe6FFsdJ8kf5WRdT
SEP1lPLwk8hBsvfyasRnVaCiws6x5GBvJ0OacoAb5Uy/LFJrCrCq/oWJvTmyHIAq5vvLReWwsYjL
6qO9v986vsNNID/9Al3/40fBj7sr76P0P6IetVFpkGGL+CGG0iNjdNfdmAf9lrtOeu8NCGcuH+rP
o0zN25D2w/Fzj2H1F3ouldfoA1V7WbGj93p8tePYFD0GGy4B/VSk8dUJKDTDSYdgvK9Uwb5zuDdy
nN5ls3Ij0k8rQVx/j+NRry2ORuQZKkNbz8DjjWAuJ9sYJ0Zr++wGlQI0IaVB8wsavlgE+54DrwPW
G23/2i51PzsuMaF/m4T9DIdv6loJ2VCPlx3ujUUsRZyHjUvjG+0ox+ydI+F/4xqqUQwJMKmnyR/a
nOw8+Ir2ArdGBO/hKtuo8/JHnvtPESykwu5uVHuP+UFc52REMe//v4tpIrbp433BiTc0knprbGWC
YCGvFRZXSijzxAGner+2dyi0AwOD3bzixZV5eTCgk5OnPVreXFY2jpx4NHe9jeWEgWqFeEEhCsp/
tQNSWjU3UZUtpeGYES3zicI5x/kNhIdeb4HY0N9ON65Q+AWWaiIIpSiXkrI33oHOVhMqynsks4XO
GvykEaKLnu70BwZocfCNq1YWM6E+cyNHE71qQIvbmdmhPydBSvNah8KqEYpAfo44dA2IPB5gzU8G
9B+RdCnfj3dreSeYU4hCVO9EZ6mzlq26ri3ZZO4YNBtGsHl85WKEJjvpSEAO4rXdjntkvU9Ge8IB
UQ3tloIABOsiHy4Uah+agIWYkJZqVyP03v7CcLfohHPUvTZgOSlf6dIZTHez1Eh8GNsKauVaI1W3
87RR7nHfxqt7LtpxgSzYpee99nIag/zY3lQTGkYzJ38YTxiE5ACb9/ixOT281EOgiGzu6b8Bjp2F
e/KN0BGiszUxK5zdZrD0/t/0uFv/JQQtD8TrTyoOozP1CNPexEz+ae3eTI45FwnRCFeuV1tff4Mq
HXY2YqbXFi7yE9yABWLKG2EPXA0Bw00TpLhA6porhaSSJ/qnh/fegRhtlrCT/PWgQa7XQk94u3yL
uSt5fugcV4cnJSRmnHZ7d73AiTc8DKL5AcSwbhld/eS8f0i5W9t8kVm5Q5vrhZHAAj69x6/p+ozw
DTwwLveJBSf0/5AIowQZxztTjPtkICBfYV5XUEF7yQNhO4+s17tNplQ1mC8ebhlND1kZugxC9Utk
WdVZy7z+PQ6Jdw/xRqwFCmC2eX2gZIPpmyPDTOr/jqUCDaxEIitz+AAccrNkhY6tZ2XgBwY+Vu6T
hYsIZ31A+kVlEYlmMb9vYZCzyM3ffCAThRQvcGH4/hVvC2/OnQRhLWirZIXfsxKEkEV5Dfifi5bm
5/2M+pymkR3SYKYDZ/M5ip3JIvq48and3bqwMRhWhpIipSyi4I4fT03IXWL8dCB4IX32zbQW653e
ahxnQaiqjYsFGh52y5+bGiq7SzY0+hPI4MaoxuILgfiq91rx7geeJ+f93ycXOeDs9oxAINN+UbA4
YUssWG2Qqk8Uj9IT+jy6ndkum4CGb8g2oRNzHWS7Z+irpb2LpJO7oSdIxOPQIX82cd/aTybvMUQQ
ddY+gFSVI30UsyYH5stMcYwqsU001rksdHM8piyKF683f+AfyecnuoOtw1kD+TE3P43HSDjiSjuQ
GXyWmgT8rEbKPjcC2WhD5k/c3gDeIBBtCJ7+EvghnOR/wPVqng8UDzwfqFJ6lJal+RWyUZ/bK1kF
FRffTYGesoz5503hfaz8Bh+M1mzNv8ZMJ0G/f+4GV5MN+zr+oWrbo2PWlj61dXAxIckJnlXlo/a7
TVq7fQXz1YvFAF5H0C0tLljsj5EfrgqzgIlbM5kCXyNmTVgBhB/FdbTisT+6aRifRR/8KoC7pmxK
mKHaLAh0XAE+fRLuNncp8cPZsEZoqOnAmJu7w402sprxD0TE1zB2QynZ7EdmLNmz2Zc392BuEIf6
eGGWd/fRxLiTQZvVKMs9xLEFQB/FS3KXq3HtkBMz6jV8SkLy+GX85qOsSnpzKNwlMsaq6bv8vzQu
hSATGTXt1Tp0tC4P/hBG0rcweroOVoIaBh0c1lIe4bH+EjwdtUnM/NX/LIlMquLir2J9A1pSFPKd
Vpy6zS8hrCL0N59twltVQ/m2HuOW7nsS68JcqHwN4+ysj0uyGoZLVz0N9ZeZnNZNXCKbF9u469Am
mnaLZ2lO5N5m5fT7kC8Fh60CBoYC4ViFDjw0St/OJWAOukPu1josoLNFv3NC6pblzB3SpOHFq0HZ
EDme06TG1vCX/FNgyvyonOYGpypUoOxyCTiiNf4pcf3WreaytIa134Kspfi9p3XVX+qrzFWfMBGs
/JFZA7lc2dgmNkohxXgdGggDqytU/P5FSfFp34fJsEiQ586RXeG6ZLkjIQWklPgOk0AEzM50lwHo
M2tG3hZZ+uuZq7mxcMH4agi8a6Ckj6PZMwdqzKrUf7/ezw3unoNMRjzjfHkFHrfv7QHGC8goW6sB
tnME/iLRkxPkicf1oTkDR4GpdisJa44lOTWAwRVTAgwHYY2ODVLmIwh9Ki5WbAbF8l2k34Hi/wxZ
kz/ohPa0bKE+yaHc2I5oZMyGp11sSImCjBHKApbnGDawvSdO3ObhoBEVAxG5DvVBI4E4vvbOVsru
YsqQOs99+ao2kPnmJFpy0GjRqnyEGk5G1zIxQNbeGetPG7U/0ctWnPlBNIYgt4sajzD+p9ZnF74M
vXZ2YZKoHfWF6yysG5BgfJ+aaJOKgknGa3Dnh4aGOwpQTvkCM/E2jWsuQoXcEmAjGQhZkhbwPmJU
1DxCE0jT1DxeP4vxp9FOJKSjVTfQDLvTlJe/JxTHg4+AQQPs8+ldB3CiAI5HeYXUtTT/Qse+l+18
MJSFIUY8lGsW6FawC9bgrEwyiGiB9ZdaIqS9Ki1edBwTrP0/uhc93M5NXsmVJnKDg9LnXCqfuHW4
X5mfzY0zy/3noSPRB6LAZulp3ScvJzsaUZ6OgwE48Js4VkOqVUdUY+mX1qPGGGJfSEHB3JPg18+n
z6dfuAdxXiwn0cNsEnkJLNuF9kHA+F2eTIDooO+60zBfEyuNihvvtKQ8v+NTP5A/YUniV5WPIjtn
VQaPlzdigEvzbwBAzoQ3YCPySQ2R8bCc5AK+XNIPg6Q/snG1YfhJtExI+JBJ3d3L1P7mZS7+e4bM
EVJNjySp81xsQp+zQUhyUny5JfcpbZ/EIG6019NOWPDPXPEMdmIZ9gkfr9eBf2PzoncVFAXwRnK9
/u/X029+gXWdoTZSjY47SUPOC7M9OV/6D+N9A8WEdlf9eKfoj3wjxD50WeEyG/e1N2nTYul2yly0
AfA3O2H655CSWVZpdjY9iK9piv2BZtkpIOJm6hs+lFvMiiClXavnjjXwToBGaax0hS/Oj4JlnEKW
n3M2O8BHqfhQqJt2CJuS8NT7u+jDQShOjy1O+btpE1SEU2NFdlbtgq2faGyUUsLg9TuvedRwyPZG
uuq4kql7LFLbxfq0qPqEyP1nF8cTVGytrK74qycflq+JzeFPrOhCbBted3guO+9lgufwJvkahOVE
y6NJlIqaR1zwU0hr54aJ1GstQIvmPU1NPz/RL6Q88ev2rH6FyE5PO7FYjhKEx9QrHopMR3bV91CQ
d5TBUhkrmxS5YfqxB20w9pq40bDo0CLAUt68zsIH2eA5HAyJzQhV61aCFqnqJm3wQuKenSdRPhed
a9o4evau1DZPePwlyQauwelND5FaWbcTpgwoZneEdim3sgurYL6XZQllxJVIXnlkxFS5TUjueBtl
eVCQwPY8yFx4rhynTCJ3lkmia5u+Ea0aWbtsOwMz7qNHpyVox5Yr/OVTV6E6gEbqC2cz3kHJMuFO
eHGdGinJlKw9md4UsUI6h6XHCtjI6N9BxfMWElV43buyOogrQmXHB9HMH7rbcFFaBCvUeliDqsKw
G/NFoLvPP+nGrsRSbiz5V6KUaN3xiAd49cYpB5/j9GpbR5rPSYsPgOjXC1RrJ5LA6Ra9hiLNcboy
TY+ySnpMfa6h+hI7+8rvXF9CQyK7VMCISPOjTOWLbzswgUo/CAxGzj4xy7y6H2osxeRDCX6dc1hH
nHL4FIjgHshUDP2J9yajiZbQ6xEZNyrSEFOnxjnsKWO2M4qQ05Gkfq4WEe0t6Kw7Y8PZmxC4r+/1
hoOu/pki1GG5M3ACBi9RU/vityfMELsoqkaoQdM15Y0hO0IEIiSdW0vDV+zvTBpVfO+jsdjOhnaP
mSRir8UbQfzutoY00phF2mUggq40eF4AzcwSQNe5RzLbuRK0KHDbHg9zNM5cCcCjju9lbcr7S0e6
7hkv59bAvSezpvaw+A2k8Bi51A1K257vynrvMFfB6KKR3dLaEhyGlkHntd5oqhwhp0hxwj3dfUsa
dnhs+qD3RaGFEc6xw0WBH/+hB9eI9h5kTiSO+NmTFaIF/JM2HwuPHX0JvZkUwsFDaXaqcrkNxnOX
74kpuHkFQk9T7ErZXAekrsHB7vaLcPok2b5oLxJlA9ohiq8bdIWWRJWLAoZHWvmjNBTkxuTj7WnZ
UaCpIEaJQaRhGAhgaygkKBF9A44vDKGTGpKLlu44Ky4bAtlIaBbzy6mtTsGy0cpIkoju4B49mwX6
hLK6ezDjwiVnmhvNypfzMfGNfWUjifKWqmn/fhnj0bLTEYjQsLHiV9E3J899AOPBSur5oN/Llzr6
J9IITNg+wxhfyLE9r4pN7naGs931MqUry+K8ZdOmWtnbAI+3CCmnSeYTgMOC5+y4cisnDhyGgc2p
cgqChhCU76MN5X1iTkqthH6XuietquCV/33yN4B1aPjef8MKBBXoqQwaAXPHTripXOG0q6x+BOIW
liYD8j9V5PvgH/fsmf44KyNUSMgDbrKBTWM0lXB1/554nKyEpcQHGtfYxBz04G6puqcgCfc3sv6U
h2RNpTp7Q5k6n39cnoZFQiut990wI0AJHEjFlTnJM+VwMVWoMYFqhZXccV3epnc44qVCy4yQjaUx
AR4CqnlnMJdflXLfe9jl9hFDbdRMaoXG0O8MElTOA7w9ooVp/jFaDGEIPahg7XGvusWGx/Hws/2S
gWB0WF0yLsdpchSFOtj6TOe6PVYCL9gsNymBJ83UNKy9+XRLDU2docfhfd8k/TTEUEFxkCbT6+X9
txrbqI9bGJ4+q8JaZfYImyYX699CjUCR78V3/BiSdOvMY24E3U92Px0pcPe9x6u791uhH03Goavn
N6nU2vtKRPXbOrRw9Y/UFqOR3U5DA+nhfWOVooicT6HTqifsdjlaMTtdodm6sAKS2SlCJAglZnyB
Z4vpxGIRclsx+8Zvnd6xnc5gSsPvqZ8ynaoX7P+vaL/mZCoTxwqL0hgb0/QChIyDaOkTntbeAbUe
axBN2IB53aQwNkecK4BStDyYzTF2qTh5PjCT9OrgTm4APVZez4zNepkywWuy6qbs6OIDIFC1hKV7
9nUQV0iCryXA1aaCtVX5xE1A7dzNc/MoBiJC5ZlKjzGH0mioT4gnFcBYYl+twsAy/lqUI1inkzcd
qcW0ocJguBRE3FqqGQaUWzPXBzLm0H43ahqsy/exPSkdYGromss+zqZwliBSHaKfIdzlBp2h7O7q
IvtSrJmkrNF3WzZjdMALwWlChAM40Fxn5tH6wYhh+gpm1QeGe7Xxcw741K0mw6eKuyIv2CN1RgOk
Y5uXobCXRWoCrc+PTCJEkbzp7RG+aZZdqBWysqbhz8/jfKCEFrto7FI+z5bslATNCsaonLjkYn/7
WQ9Zw/SC/o55kcGNySM3fQsrxWNMXu6L6mAOAIPLC6QgLYSiP7JlWV6mcD6YBkeHQLMXVa9WpY9G
wgETP1WYGcXdT4XSgFo8U6CT8oWFyb2kcB/1GRQVaobDjqeLwLWrMMuGcFmTnjE07FRBMSf/H/uX
Guw74hpFbYU+a6IldlqYdDoK2An58uL6mEllLc/JZfo5GL5nfc0DcQimweDcTvOgPPb9mI2zNLLc
0uPvYoNoPzrB/Lui6L/j5st2WtXjuUqYIB/JF8OYE5+wwkHt3CcjHFU21Opu6qwgU9H6/tzzu0eG
AFgUXZfjwJucsbZeLIj7UafU8/MVxl6dhZctGcdTU9Clpm5hwyEh6iZGodijX5qL3kGWf33B3zUK
9mT1U8s36YmxWDs87nQN5ZJlkQB1o9pTTgsSLcNxgmoBHTsXDbc+cE1aCag0a3LMMBz3O47VOBjS
A7KXGc0z8QDDuE4xQeMC3DAUryUobtjjn35khzYV+5jTs/lx6C5QLUGIJfoftJsNFlBMTmMRN03A
wQVt7Ys4oBmJ4mpya8kkDKxkOo8x/gAYd5KQJBSEBhiCAAFpF6KHQn8yBpr2qCpHMlaYtrnhzpNg
2FkUX52FopDD/2DDh2sjBkquIgHr1K/lGTbTM3OL+F6Z0BPc6oQAYbyyyTk2QPlVRVJ5jxMWnNTd
Bt1TidjDmauCiOSFKTwYuessdi4EEn8Fqlgq9mVo21ie+eHSKiEFRMKrZO6vENpRwc+1+Svuvk/l
M91zj7Peo+Kb1DVM0MLjSzg7NAI2SQCXmMjVTOt3uYzB895ammrVSMdgqTFUawCSMfJu5NefnoWe
Y5nrFjaWnJLzdKxKTz4AfPO5TnSdHINsZJbA0phfHxOCHtYNQ2FMYBN9gcVIBzuHW1HO877Iv1MQ
7PC2I+KnwD0zKJ69ontm335IDQoCcjGIPw1IA0EAeOGGCf83I2YcpJtDaNR0ygMp/AKS4ZBCCG9z
XllnR6L5rXRVtk4Wks8qUeFWu5x/5pq0KG590lf799tP4t5P/PpS7W0kupX55wZXUjrlD12vUHhi
Z8/s96wk6sZHRbGhDwRPWRA2/YEyU4mkMgYKrDG02XsCdKLV11EnD33vnHTO7NQCASuQMuc7Yw3s
ywLQDIZmEQlCZPhq47e578vLVJxcqL2udFxe4VgN7/Ypa98HHiQvTCFIE4rSgmCaDoM6BMuRnu9E
jAVjSlGvL6b+NpxK5N9FLFmVP6MHWEnFcyRX4gkd6dnBAHzBi+0vjVcUAJl6ZKyHNvaKFHHRl2lE
vZDHbF3GDiHQGX8GTbqelMcgcvD0YbqmhaJeJy/9yKg7HLZDQKC4K6SlcRbNmM7WHiKXmaXkGWkt
BwnHfCB7du+hM7wtDVD+whozuCfxz0FSXmyEbThpGMDIgqpLZqMvC9qJ+m6w7XxP2ugOAaxIFqQp
XgT43xU68FZ7gJpxIwHht05W2KF20Ri7QA6KnPxXcKUFahqPlEgxNrBZKVebdiqbSoAduJD0tAal
OJc8+eINl6ryaQ+sQVrK9PO5g027jBIoMm9jER1xvQP4iQ1Eteq7Wcq2vOnCcmMRVxl7fCCh0EHn
cmLiO4WjbS2E0fk1R+SiIvdDPEXVMPfY9js/Nc8tlK2vYVYLkQ73f/5ebYch2pV8TOf2KGK6Xmtw
wSHSTgHodjY5Pwu0/Hby+uIEgV0I9G6zBMJyE2u0hmaYvUJXVKzdzWkZFycUbzeBLPC3E1ziC8pb
95gF6IchSa36wsdXtuZbv8jE6mh+pZ5EAWkizQSSG1zGPGrMl8rAXs3429vWU011WlIURxnUZnz9
iHIEsK54Giai3+Kgq9oTLN9h7x2wLOZRb/p4JqE0gAuGUti/v9HFDt2nhQAo6f46ljHeFkN5AZAd
19nXTI7f6X8Kme251LF+E0gpUSoGx+8JgTOCv6sRWiOpbEafHfHbBjtvDdX0iGHCZmWNJEODMK/A
7+psrEs0UIiHA1Kr3Te5ea4vtEX/lPtgYiSVB97vxEaiMWv+ytYZeA+tz285jlVok1QKBtGVIGlS
tdWhs7ixJ+iVK/es++ci41kvHKRdyskThKwDlPbBC2IqlJkHFBgNsrrY/zL0LTHAV3srLIP7+I6d
wJsRcbZBUUN0K0JIt228P7pZD544GHXwHERb79jrOpFtzRRTdKibAb63WPv4soZLZEU5uXdkPOXd
v/KY3oQsJW9H6+iad19psyQ8u69T8TJ61crzNavOMJHhidOOhEZHQVRWHVPpcpwPma9nsJ54zns2
g3bpvHNtEfRs2j8DwAic1tm660DOTMFEs6VIAtRmGwzAsd3lXkY0R0YzLTDXj31m6yc2k5TZJjys
UBxEgH88gZZeTcpBHf55egwQaMnCb673dV5PLf5AB7WQEl6B94CvCZthJIcvfXcLksSGix61T0J3
9mwfYUBafxEtZWherb37wtfzXotf41nla9J42EI1xp4MaI8sY/Y+1gRWURIZSx0xMKF2e3Mk6fSh
4SZrtUMLxMnQW3pNcuch9RbRff4MGGadyCmx1VXOCbNgADo48l8k4koEK+BV+RR2ZIsFL4EflypZ
s0fMlQODTSJP5WwFxGrbbbNPVV1wl0qx3DGqdzKhKRCWd4SD+rYUgK8kJgY7uBBGPTcjN+rhzL17
5jfgu3MSMQ/kXR5ByE5+WuxBC0m9PB4SahiMD93Esmj30uQLCcOF7jQxFAPd31qU54MEogNTvEy4
fMZZ3eA8qQUSWAxsUjkZVxgMq3Le/0xfW+3ditqXj0Q3qelYH/aXcuJ0aU7R+4iYFk625pHuDWgM
IXEsLoNf6NSI6Gf26KbcbNLj50j8WDh+wF31KKidB/TpizFe8Vp1+G8bYxJXsBUMzSPlbESw7BGE
LFn6DVQDeYLFj5arjI0vZHVeuOZOct6d3vEt8xSph80x1XNQbLa0AKYZvzN6YT6N1JM+uUkFNBAd
gKJbohQMjymLdvbzT3QNJblmGrskSqoKl/i5J3CfQhD77Fqy6unDRgcn30FSbL7nDiZLMbaQSvGi
P4M6MZ6Ky2jzqpGs56b6ZNYJq5sx5RCnVz9VQNlaBEQBlcqAk9ujKSt0JoXpF4ZfmepnGXuQKuM9
VGMRGQeP+WhsucT55hmD425k2VnZwWajdZKTaR0K0gtoXWsyV6G9RP6Vm/jLgK9kRkw7VXuWx6WV
FHkuKG5gpRrVU2yH7NBIFdj1KiyP3UxFCTyOeZc5kOkynUx8hX0CkX1tyMsiV0wZB88kOB9UFOn6
rlKofYkhYrTYdTJi3Mwd81jrmSkaGKvKC+BUGhy+OkiGU00fGe52pfU0jz0gbWY16IlCCTgxvkuA
yXNQqOY8bDbdGVELoCv01LHg6suHwSdfIPJulEWT0YunJuTvt0k1oS2NJw8vC0ECw53+oPgexB1g
7eXxVZBxKO7eJ4C1iEn4ouDvlO/ZGQvTRM81uqzdWMhcQCZWxp2fVMLm3rd1ipEYuPkfPymqnaid
qaIWrkcUx6fVBNbxo065gZU6lPEiJEwdqBGLiLw7Empj6x/A6heDIVRg1MW+IGXKX3d/RFjZdERF
EnQVyyjdT0hhWGHRVkWLavxeqEhdcNvLxuBwZiSsVRQNcl9jOILItNt7BCfMDiCZXmvqdHPgQ0dc
I9/x37wvM5cTJbLXjPgQYSE7hX1UAQIPfDp33jQol2YwC3IUrNZOdXfpvO8ZKxZUFOEir2TLcQdH
ysmEh4U9IpIUd8uWzIRskuA7y1UogpankUJm1IFqph3PfdwHJkxEqGFrTkDc1LvDl7AKZw3Ab8LO
ljUU9WC9yhLr+2Em1IZHhj6sXZ1UDDx04yTvi5NHDzhXJQg2S68mWkEyjdUFChNCgxNSRGDZ6x1h
7/5LxdXfMDJIBL6Od7MgKX1koG8Q1nihmohwwBnHGCz7A0nOmDL7KjOGSMyjEmQDS5KE+SAxb+Wg
WC5xX4N9cqyW1s/Fb0xCbVfBmBnn5W9K0/Qzjwzfx4Yu6WJIDkCm5T8ExgZVYpekVzEpNcy9pAdn
JkEkn91UV/rqordJ5NIxKL1BrWg5lYVeE1qIaI/MTB1uEitnSfnGoSHYI5awpxIIEeQAaINZEB+9
2ZRQpNNWkELtT12AMNz6a0VZZrlRjo7fwVBHRzEzn0kJitTWmbLE/ybvgFc+H0BN1fdc/Z4NGiVN
vdsZA9oy85Cr3FMtnZ/+2F/HXL0VWqQvsUIq/NBUHMZcPT3cdsHCLOwNBr9AYfGAEnZ61IAM2sCQ
EEskA9GS/tue4niwgkhOxuHEtDgQMi7YF2nFiexrndjNDRCjSQ51HidS1Khjoy0ClBG0n0cmZCvj
wuYyFaJBUSzrSuWpxSWKpty2mMB5MNtT/dcbUD2ad/8aDQiT+ka6664CEIzG6P+BXlhkS2ZjfuFb
KrWcSyb/mA1GNjR4C11WB5cFdAvnSY8Vqy2oCrHuctD9PVR6f88OFQ4GzcF+1xGa0VrO4rafQU5P
GwR5ApKmalqhuYU5F0B6W+gtIZEOX6QbfpWCImrYbR4njSQnVR0GAkWtG//pcB4CFlSkcRoROVj8
5TdTPrYLZo69aiDqsTIWha/dmQHdQ7wEzMZyzf/YIczJLkMApWHlHPI8eW3Bw1ajeyUhxTVulq5l
RcMg4936u/z5JwRdRaEGPPZZMJffNQi2EI3BVST41ugXa3qeTEdY+m/5Hk5cPZzzN+CvMSbkeuvT
ykqUYJLGEyUcVvNGt5iy6nDb3uL0dbkA/Z50vklNlCSoqToPkyHD0Sme9nJ8cpY2viTmKNMPgl0f
/ehSbjB4BJU2aR5RgcHSJit8EvjSEsbxaF06I6XjWIJfil9q1B6djJBoXRXTN6pgYj78SjYo1+kQ
2Nxs8fBYi6a5lGf5Undn6Q7KQKJd7KD4qrHc4JbT+xF3Y19Yfj7gH1qAUmHzq2NEc3wRLGnymE3U
ZxhiGOvEWsMlf7T/9mVVYqr6LyyxEtRr+6/2qLaYw3ZFak2uGPBaKK9jp3D3TcIyWzjbcpSy0UyM
S0OUTH5j+3Fp0z7dQH/4GtVomCLJQnMOsOwJW8yZpVMe4STcttH8M0MMpdPANXI+rvvL3L8gMx7u
tGQGeSePjE7cDz+esfh9aLlx0Uf/wyeETNLoz7F8z/s5HjRDbV8IiDC9zxmRk5lQGIcz8zt8Yz/S
4x2Q7qFwR9NAaRkQWsgZQcdCzMDqwkCqMqdfu6WOifWqdaTPkhzNrxwuYF3Xsli0QJSEPfXb+U7y
scZ7vKdrhi5/w2ibdt4QsDuPcU/pG5Eky5TN3YDoCLlkFFSrMovx+geDFVEfF+yubCn8JSmkB/7o
ATp8YSnzBdHzXA5eeX+Zpe+9x6E39D9iGHn6MrREswgZD99SMeHXwXsU8bj/EaBGw526DrnUjdrr
lg3b4CT88S6mPYBuHbFka55hJSeoyZZgL2GSXz7zBeFK/+Xfel2jyZtE+DR2c0TBQQt84JVDWygM
1766GAPzUZyUXhzOyV9+jH5wHmgd3E2Qv96fo1MvTwYqRfYS82sMiwlChj2F7R7Ol5KSLpC8eELV
HX5lCwKV1BZIlbe9+dWTy8YziukuNNkBQ3bytgfbV/9Nf9M3sFplBGHJIJXyhHRgSDUc/ssgWPQS
Pdoz046TGtvrYmDrQg7RCvEjXNHmjKBaSN3lDthd5hvOYEtkFjJZ2oemRB1t/eAOQ997bdvIYwVT
nsyvPpesBYJ7+7TtsWGdGZnIMKa+xX/ekiTk+GsTRpmWs2Rzr9O6KHYDzhwufFRR6SVPuB/FN1cl
8JJDvDRw7Qoi+WDCzWhyzu6SDxmqgVstPd+Z3WIJqUe1sE96GO88692RAXtlEDt9YNaTKRhEXpnZ
VnNqJ141vkoS9+URkCXC7S4Bh/2gSGuyRQYX2z26T1d8Bcg+2KUx0hwhKeXsnMotMhFEj7zEyCzu
tYwGZJgBTeUV90ZdAJtw4sN0f72AoMlFrdBEiC26LvhpjgxjCKgkKesnIDOHX5y9gxSAG8DsSF6h
ebuuNqK054AYmUa0iBTk6CYFWoRdL3wuC8bCQnR5+wnUT1SkntnWW7Nzp4mWEWKQWdPygpVPoegq
FbwxQpYHP7UumfciD1hL9baYsqk/it5VPfBwymn/lVZN8nG0UVwqktc93u4NNkXed1Cf/9TpP60J
dDKRgolqhjCF3dwGG+AMGO0zhd3ymzfv/FCdYTiECFYOT8QRfVk1t4faeyaMCowRA6Y+cji+pdZ+
DHV/Yj3JHhIsF0if+xU6jUKrlzvn/n52TN/8qsotRhKlLT9t8f/FED/DqKQM+Jbaj6I9ekEWTZLR
BFxjivVlaLvGLlXn1TWAFkSCyOzpTX859JZNy2YlV3NGlAEPQpG4+Lr/Aqr7VhtPYBQGSJdvwYWs
Wsjl94j+xg32cRwthh73qxDMcKw2/T2B6zbpOwK46y0dBg9+rD4LVMyY9N1HPYYTv/IORiqxHN+H
vFcpEz8xJWa9Auk8DNrfV8oJeRrwgLLrvKADc5zjAGvS5Y/B3axe5tNTqIdDV48dNZHhv0jSFGq8
IQLQqkUGC5rHbdzEGf3qA5PwJYrgzOwd+IJpyk7AhOaXDxAZdJ91Be/Y2gS+pNDMgJVIgDYn+rFu
sypMH374Vwce6rwoGIAWSqrWVX7Ul6P7fvoNwN+I/LMEhBTZaGooefhYWxZ9eaJH+vTUjuP5zlWC
RYSMTKIHUsZlFhd1aJtvo/GSyS6ZPdrPTKPcRPxBkvpEt//OrtTF3kwNETHUYrVrmhHqN/YHdYf4
Bnc9jnLFycufxo6dHUlsIf9FY/sHUmnL8wzYsCmps38HuCWXrtDTo025KDE+2za7eTbxb96KCh2N
o6UGGqGueXq4cCPrYFn+her31JzjLHY3Kz3vGV0yFti12Axzfeb+6tvG0XkOTdQavtkqZyK/8Sy3
bV6OIAxvIgNSN2CUfptOHoBYDh/5MS/aCdcliDDx2D+PkgGJCiB8iV6abJJBIMpQsxxsnF2PlUvu
y6a6ZN15xgqHi5Tgw7nK1XRAHABXkB+BmXG0FW2SYR5V4UEtRQ4Ybze3JFivDHPaSOOVHxviQTE5
s5MNrpJObFQqxf+jGFdsx0r6M1WDFCLl9GCo3dqrZ/PmQKQat/JsbZNfHnLPPis4/wWwE2+P1eMy
rQR5XJnl21jpELQZmfuI4IQGhbbq77kWndO02x2mXp8/WUyJzs6glemwiqllldsEh0W6lVoubFjW
bi2qEtp3yZERl4dVzWoOZd0nUhNbliQ6uQrnWMXeKBjaSkPQi5fK6niFkbBzFXD9w7X1JCigeVfq
JehBtkdNMux/F3yDlUcuG8k0e9WIVBfv4wMdQhESWVmPlDrt9RqR0boxBH6R4419m9GXaCsdCRy5
nIuAPMcfzMbM4I2Y/5vCb+85931q+IPGZDKXZDuMRty2VVUk/B5ilKGONdzFsysBmLHtGkiDSII8
NN4GZGtyl8hcsDFnOjasCEKoynte6gBqhPjoGIeXw0PhoqTHxNt75LZ6OTBBcG6gCt9x0wsKf8ux
kELDh5PFbQ3Gi8T70ozvM3mNC/olFzKrmbvWCgoPdsQjBICt9hCfSog34yMD3PLO7eVLB4TztOTG
OmV3SnbdjA3TsNjdU5gQPH31wrubWtk56N15bYvOxmIrKtMRJKN1KwoEf3GbDZjXmoryoMNJp79z
7kQcrpkkIgLkEtPhm7SsGriifE3/TrRl3MnoaqAa+ozGrKCZFTa1s3XbUgQN3B/Nvl6mOBzKY7WP
kig8lX07nOxH36D+hdEc8jQFCqkfpR+qkbc8xs/2xLBjFQ9/2cZta7X+bgZ0NeFdAp9ZLVg2bmoS
n3CvZ8ifZBYlY9fdaISo+NxvulkKbQ7eEJeMQGUWcVe0NMeR0I2LxYjLKmNSz6+UafuZSRtDvXNg
N3tSP6ODuR7C2vYvNBDFPC+dSyP2YNB7u2MjktC9l3pF6MrI3BJAgI5N/yuH75AcInqoBwW9pTA/
SUNGodAAgAEvvursPG2ol1r8azXxjxgOgETy0+7TR/1xOMu11JticzBEYxVf+hj2Un+vOJjVsX6B
Ro5ZhbAkqA8+d7+xmd4yPXJapbZ9kJ2tjSIhSmmkNLrKHhNFHb1kiWfOGSTh3vgpoN4wxwqFiA+V
Ns77HbTFRWOxmv+I0qWwd90Z7dIJY8v1xmcj5icectKrJb6gA/GoUFydkEUy7F5/0GOIbbMv4Oz5
WPVmIYTj6wVgu81KGK8/iFR89cUTrh4XZl2qACUP5ZF6aYoxKAiOV/oQ+yald9u5Z7Qc2G5EJ1s/
pqxVUfvONuHRaZlS/bU0WJDK+5ZynXCpZQ4prQiqfHLOJWEc6nMbBrvR9FRy6zDkgOQ7Db9CHtSf
jvTwF15pIXCOx/5qr59H+q21mpfwI0IL1RowQcD0YHQ/PBQISfGlWSMCIsV6tG26SKLN271WGv2r
6ifQlXOBS1pKSyqa5BvYjk9xVz+MV4tBV+gxtTJ32vRnbBZ11el1Mz9MJkHjJYV911cciF2Ux+ra
ycrs/sL8Qo3EcVvpV7rhrN/RN9/KuDpNg6bNOU+P30InIX/mU4D80TT8y9NNJoD839dZ0FlOns+s
3G7iHPsClYGA7Jn7DtcP6Yx1/kiauGXFIEksK2OryX0xAQeAQrXnJMSy2VoU1d2o/ClUSO0mKK16
H2wy7g7lZ3lybqTv3Ryyt24LlRDO3jy8JUiRMOWU2KGbEef04qZUTFS13XtfGfbb5e392ZCc8VIf
Qr4qiIMSeItcN0RxwPlTYdzX3VDUOVRghRt+ARe3KcvK9q83QklZ6PdiuJt+3JKxVHcsM4l0Yj+t
TESmMgtFwY+VhpBYLMtCjU8Paq0bgKMjDgAE7e9YgrxIpA6igY+PdiXSXEQkFEwwA4gBsd/qOuzZ
Dc4nNwHtaDxWQ6DQRgwAPxkQHCYBEUF08SrDGhmHmWGKqD8G1okpHT6PnFhODvrdazihZVwSCElo
U0jnKX3bjZeqWPHS5gttsBbRPASozO9RyU3nVe3yor9mMux64+SxEvPpHVRvuTRneiD1QKClVHwf
hYiJGCgPb5pLJc6Mn0+Slx1yj7MSHMuutMkYDvH5jwpiztLnZXLohBPdyXR77JITwU5XNaynTC01
pE+n2LdNy8xFkyqGj13aOU7WQhkX8Bk1vINRmNPlwmXJRmNeyhVgoZcfeRpB3ynzVd1ZSDfaCSMu
qsRCU9e3h9u22R2fFunWvHYrCjvPST58zo+nOq5DTgNe8/hx2pfEP59KARlOSsLrP2oK1b3+6ABC
GxI/S1nRSDl3pw0Q0wLqEXIcwCN1bG9XXdyHX7cWn0oCDDkZQLrWPcePhItEX1VdWnuXzNRO0FQj
cCrWNDWScGQY+g5T0MXc6AIb/dqcgXwCIuBZXZ0Ecj9lQwFKDPuP5RDKi/sgR8nC/hRj53VAhJTQ
UvctUzgM3roj3MugDd59uN28eC0XzbFuNe71F80u1RFHs6ollcLmStGqpb6oqgAn1rxo5dTQPbhx
yTO5s9PUL/3ACJf0RqNaC35rMDe5UsnTYm+4HI5l+WZ5O5uzCw1rT+JQ5UIwn/kafgqYY7yYHSnb
Jb7OIvKykfaS4wEYP2ykkxUeJNC9hsN5PfXGOUbDwgKEccUdJTVljM6sMA9PShSxhLujbXxqNc5o
1uY8lrm6ryQGWytz4K9kjJG/EdQcgTB6TWgqjjtRJYztSllVNc2XOZjSra7M/+xwhGxaLsxxsTPy
gjTxcLlw1wIWsbATUwEM8Bs5KnGZ1UvmU17jusDQgIQlxv70BWo69K5TuVc8JMbflbDV3NrUohen
Lj5ra/xdUTmGrAQFmgVLf352c7/5WFWt7CEhwQhU8oo2fTjH6eRAb3Gd+xSe6rYfndHYSoN3URyH
9FeT6Gjq3SA0R4c7YzlN5HOXyGp5hdXQXuen7j0eUMCRSPXPYQpxL4rM+sMO9H5Qw2roJ+DbTFGX
TtiMu7VWQHSWzS5ORzq0uK23wYhWSFsZUS7+xX8/OpTU1GXbafO8qjv9SYmBfcKUZBbck4TMvCrz
8eGX1QVbFI8NGmG1CByNDh/166+QfLQ4lLrCqEJ7UP6TMVGixw72JT+P8Y03wGy+aU39ymL8NAj2
1LWxHp4IvlXd4iHWlxkZ5nqf421THMriMpfcVebKrntk+hwIfNQ2X0nZ8/N/Nxni8MZ1B409FPP3
h/2sO76rANX5xcUFS0m8hPo3TK139L7rsul2FWGPptCkpIvBUVensh7CTnURih2GjX6jPHDXJu9r
AZxshTsp9MoAAHDi0pRN+R3pFssguPkxBcyxEDkgQnBEY2DA5yVfIauwbhSFK/Ro7Bi5qFjjM4XX
A62x43EqHvTWhAfeTepC384H0a1OAbN4Z4R6NqIIcuqGFOEDZfmVsUb7nzVdGrSAXE55dy7D/7sF
SnxYRiU+5uopE+VSpACMx5EkDujeOwD6GBTf6zy/qAuegGgxKflHBEWH8xD1lAkgrDTm0DsyU+qY
jr10shjUVom6Ob7qFyaY5taeSiPTxknvaf1lYxdX9hYxfUYGBF8J6Lim5v4a18TDFT4s6WpWakp1
OZZ/dv6jJlor4x09Dl5BuSY0q947rcjYC2qFNWRRXsBYH0sHWmYBx2YH4aDpbIKHHZKE+5ThAPGe
aih8wf+V+t387HAj+n14OU3wxoLkb63IhRaPHl5DP0GwzZRcLxEwlKnZy45PnqZp5Nzeor4nPNFR
+stUGnppZnAiZ1Km9bXGUNYnkOglhLHREp4wUQyzMkoD5Zas7dtLE5EsluyPo3b2I+GGmWqdiW7T
QafUSnVQTFphzCfKccEmPizGOS5YA+HuP23Lg/jDv3XkV2uZhqizACHR9/YSqG+dy/94rQzpoE8X
bwRoMczJDJav+TXomCQ6DWLKjxVR/y2wza3WO4+THDES2oVRvLST9+v8WX4QIZGWsO3U+E4WiMiu
xIykIObLIJVm484pdxmQDVsKMvJAPK+YQL5rzrVz/Mk34x5otpQUThy0u6YpF/YBtjBrVSzb5/zr
VkcaXMPuWYGEtX2ACI6kTMQ8uQ/tQ5MOX2UaugybDj14FEdlJdkmFKrOMMOJOhr5/5iNlqZT55h7
nHeljmkEHbspHOaQheMAOkeArQMDi4qfD9DnaeAP1Yx1TUlI3x0tdLL4LnOaE2FCe/1eafcMDLAG
m/oremvp2y98QglhOsqJx1xdXfiSoNtjW2x7X0fDUb3ohe0AQcOs+nRi7hYP7hlL68eAKbaySC3e
yseX6JIq8MhYBxqzxuOozukKv46DtxmrKPHVWfLpk+wvqWyWJUP/jCBvFY4m/CAMiJfV7CpDC+wh
gvDNq2N133PmKCvzVEmX9lpKCOnQZL4M+qfcSU++sVXzyk/C1vZW2H1G5oR5LiDJKqIJhTkBcuDP
TxOCOTo26Uo5gOxpzJIb43ewnedaderTvqH+MURPUFIa8KH8/D+TaA0QcpJl0EtLCu9IF6vQ3xnv
zWHQNH/PQoIUfY5Nh7WAtrz+MGA8wTuAEJgz8Tk/RkelcJ9ueWWOs3udSh7g9Hp01QYxy4lvaK31
Gd+vza2Obtpeq/6Kt6NleN/KqltCaABLaGKpxbBCIwd38QlHtzUQB7uUP+wDh4mJJqb4AvcI8242
eSeKtd8GVLM8bqagt056+LXvokAyEO4Kdfxzf0QNSk3t/7zRvSQJr0ma5FRBnvmfUawWOhBYJpyp
qOVDoQCihrbZTQp7xw3g7QxMsqWu0V1+FFIeBJ9d945PJNiNCsR30kLPVt+L1oLyKI751MfnVVyV
mVnZxUY5Cz5HT66G5nXwQsSiXRb9qsJwVrNi1mqkjOj9kVLEvUydLBGumhKlyZMnUimDFK42Bn2S
xxgVTJAIfaf2HIinhK+xloFnhsguMW2QlKhaD1AonfFpoHtXnjlEBtusosVHxy9lvhUVcUZPON+t
LwVuQmkOx7WfMA8Xq+ruUa1pjxw4VRmpzaOHznaOnjll6aEbP5GdfXLqKTWZC5YE7Rry+LESygOn
KcVLr98FG36DkKbuDZiQbjEQEvl9U/1Zs+FJwmjrRL0muMWY9ikuCIxPrjnA6a+sAbIQ0itRTHpk
pWT3iezig+Ig53Zs1DrSF/sX3NbXbrD1k2+nQ41Xq8lGzDH+eu3EhuZg6nD+PAB7sO6s+cz6x7Uu
ClJWgH5gyvP9pwd0nl6krwiuZzB+RtYWwD0klsGfQryPsWbmyx105l5ub34wOpRczX9rNC+ydqS+
zrwiK9Rf86BPZ5VbVqD8/3jLGZa5RQHokut2a6vb1mgLuVJtRIjp76BiTsqwyIWpZ5UGO+tC43cX
ku185ZyLtAhafW/R5asFp/jURTtdODZNgoM4Mtzmf2NlL1CL8TjLx3LBcFkpaYsiHskS70VXSeu0
LEhVi+qoY/FEop1KxWRiqZJz/FOg3YAaEhbA/klg6fjxrgE1BUdDVBBcjSiEQU3wL1tlRajlYJW2
6n5fzCE3x6T67c90bGGezYUe+w0kwlfdTs8uWt1tlCbfsc75ra90d1ZVHGJ1+kuZNGP8uiExtyRV
KDw/uL7mnZi51mNerChoYYTnFe90eDYLqCP8+CFGolZX7W/pqrCjyWjFAjxWus2D9te8UxftmZ5m
hrQDSt1LiJtzj/guqVOSFMW6XHayM+JDTHaqploLE+CXnsFKk/n9kHTiTEMVrzPlPQAtwKsfWgGa
08iH0kEQ3bEKS58p/1bKMkIGZAq/thkTJGjRo2lirBeo6o7XovlZs/2wPa1r0wQ6f9moNXUaOaAE
Lg1ePcJ7rmnkpqdOhiz8CGX+jJ/4YYW3Njx2VTtQXvPr3dswwYHc9M8h0SF149Owgna5W/M5OHcE
WyuvDWJN4cbBcVVgwmFQmk6vsUbLuSqiUzZlQdS5LKFgRq4MV8A1LRunS5YaGSox7LhjWbZsfFmN
kNJnpmMPtMavYrGla0x/ybiiyXiXkum+w/w9OAgZ3jPR6WHJauhoAOYxuy5Y3RBJ4CddiIW83jxA
+hOo0fwZm0tri3lh1LHD2TZxihG56bn8mXG0mniFF9JYSrqGGAFh1G7ghsXSeE025pg3QOeCC9Do
KDxiWzsCl+xGJAt7h6W5wZwZjbTTljDmGRdGv7IqVs1KYFLct3K70hsaxmDVkEaot6BAm70Ae/PC
yw2vp5H7r5f3WL36Pw+KKiJjQFVWbOU+1Abgnho+Tiy7udyA68NcLEd8DgTfP610MEZ5HXKhusP0
Ed8z0fZ4YUdlENOwV3aTO+2rMEcwZwE5+lvSfdqDLITIw8CGkg1ikD93BgLP4nNuDvH91im8CecX
aA7uEM7o6f3kk84+eVw7WfI+XcZ/h++hUzxozmnlLbIdVSmcxkrzjc6pVsk0PMq+oM4c+R+xmE8A
fISzE8fkkTuZHiMFskK4UNnhDMVQ0GEf2Pd54i6s7h7XO7EPe0ClY6hh4bEvu6ZqRZ/pZ50Be8pH
hnJq76ZaMV+uBYyeazxQVxXO4HUZNYPPHDU87AtBhRedi5SMenknAWTVmL28sepqdRUlJQu15MMn
lsaCLrv+rJNOqFNkAaLO6AnyHcMe2w/p8Q+FcYzIXq8XHqxb/67yp/Nrt0kJC4ZYbE8ChBOnGd42
RbVPi/P61hHEFGM6dqAluF+H8G+6Ym2XwPjpph+TDmZuhKPTqxso5iYtP3iPRKkygUzhI1ID/S6w
8xAtt+tbcUlx3WaHacVUUQJGE/C9exGfvpQoH27EQGAFndnWJRIpSyqafOozVQoFCMfvl4PK6g3x
6c559NBPaE8kBNrPzaEG06kxiWVT9yBvApROIGxER2vXdHJvE7t7sky9Rt4VNEuBsIXnkOpGDV8P
QA6oyrWJePtckg/GUNeuZvo+N4lTyf5RB//2Ol0tE/JhhMGMPI+idpa2K++PGCQfsfjUOLXVqKr5
SLmosr7nJvhXybM7KHZ6BI3Wbkk7hpjzXkMEQTGiOEx0dG/rdajsqF9PzjGHmu+3MpVdFMPotL7l
fhKpgpUQjXZG2CikzMLq86rxcL+9r+GeYgDRwTC0O4YwSM8rnyimK9OXrgHWdLBJS8hlMTCUorrA
aShd4sQRqRciGNDqTOcBcMwxTbzqtx8S1XXro4k1InI/UkeFbrFW+tAuc2d1vY+RwPAq+YxEcyIg
GWfzqHehiXY5vuz0OVN95+jF+m59xy2OEjtMnLEEG+VGElBrgLPQQVwdif+dz9F1QPKmXkVO0WLJ
2c44Of2p0WH8ZbJwhQIezhzuZzdCAsGD41bFXelfUsi75RQtDBr7PMMc4npBE+oPk4WPar9EGhZa
PAom9eOlv92jwl/j9UpBHnsrgzl/tdGXUpf/9dJklImRLloibH7ovbS0Rm7w8oYOFicZB0P0BB20
isCHin1lSDPlHnRyS/whqTFXTpD0Fo7yUMds44w5T8n9vE8mX4OY2wkn8qtkekgqBQWr31YxdvrT
3Cwvtf2RStiaf3I1BAVF1SS48wM1IcKill9WLOgiOd7wZ/n3LHqdkJLZW0zWSXu9jFAfKz7F10kI
4lCmNQ6pbAQpygTGq05IMwPEDyG3sKLgkcyz6ayAwAbFeaVVcjRr/Cs73QHrMgDVYzLAy1qVWkeu
+ej/Cdk4IvuxhmU1vmBr9F2f/PQRPSCZ7fSDkfe5bfHFV6HG3hpmY1+nrC2bdaH7+yNfIgR/TrIK
P6zH8m304JHJoqX/n0utOI3ASVXzdY+FZioZVaeax1UNjyBC+szhy0UHUBYmtiPKXDb9yBJx8Pal
mQ7E55rRQwQoiltHgd+Ks5TR86TO6V4r9R6MJhgvcPUaqlznJ1nIDGFJzaKvPaMfcRnz6QgZFq63
2lHU+JiWA7XxCYA24mYgB+HJe9ZEsOkHORC2Y2sFKE91iuWDiQW+8y+RemFbBoDuA7BPx/c0u+A+
gZ5nVlfguZd5Y/TcxftCx9RFgoPBJjcmICLK721TYYunEUR2Yg2RTguX8U/1SNzoMzdPvsVMPjDh
0MwBrZQ0JNq/FTrbSOMiBIZHZQ2M91/ZPhLrxsyN0mnghyn+zpEjQePIRTIPf/F52TNkn5Lr1Y/l
Y+2eNIkm5M05zt1uIATZwT+eHmyAPkKq4hBC7am+uKk7HCQbmLOEjH6h5Sljqvn/b+V10XtQhL69
PE2cKgZJistjBPi21tRLUd47k4b3mSKEDN8J2R6d7xrQC9v7DDRpdwgmEQ0TbzfreBuDmOIedOCm
B/qm0KRRLEqIuGqT882IDHa3ScU6kH4XdfguVkynpQzwz6o5ayD0X5N4sc6oAeNeVoYElaYijvcG
FlCZMgo2Z+NMSE+aN63gQ0nDa77vSUbKMhIgHAwUJbpnId1pwsSMig3V85OwaKoymzRpwlj9eXId
K7po6vUwPt25IDd2cjgvrD2hrQ0Jq/lVEpuz8yIOdofLOJxS+YkcEeE0CU4TvXwG5FkInylqXf7k
nYGs5u7rOjp4JtWG6AoikPphYQ8fApByTioEUo811r4GHEwHKd4jjKu6fEl1V2AJKCpsxCxbCNF8
ciGHaHthkKHqz25S6Yj/w643+Ol+wFL0U8agafIOe5wk0DxozxVWIM2qxDeXaFHODS+1zV/e0/ax
RJ8Sbp100NUN+mrmaNYBtkBNiKjgPKuVEsQW8pHgHCpU0BJ9uS70bfciQxn1HQ0GLwjpWf8z6pOz
Zz5gPabTnkQkb9451xjMluq45++AygI1Z2m2kkY3dHEdVoFPKl0M7jj7fBv3P3qMt1CZ4OAa9Fib
Ls/ntAFYRHDyb/PzLzXargBw5i6YtwBQnsWkxRYv8765Qy7f3yFKSUXB2/+kS/UXpmfd2XbDve70
BPVZK5iOXMA3nSUO1CCjvm3UjFAXAG8Pw92q+tclcjqlkcZrEaXYpgy4r7WzXfR1T1KvcNd4wudC
9dV1SP+puzc+vFkRqOkiXzzOtQvehM0Mrhft8cCQlQCpyHN47soa590FUeMF59poygpxlnlcOUcO
GPhWNaB4RonolzcTTZkQt+i6FEY6jaUffmK6k2d4zDxNl0pDGxZPDU8ogZ9jQbQ6P4bsLF7ENI9g
J+WdsOdokdpfr2Sv0hq7p50ItiMolUYZ+r0Bgt975nhlyKJb3nx6r14HgrZEKmfF+U5wwggXLozY
ouR+pqSrAyey4ZK+l8ScxxVAFvX/H0jNBUFa7ukazEuv2+WMAComSN2iawtcAxNHMmUUUNgrjrx+
K/6nJAckFHgSo8FINjyGw4e/mzAL8vNDeSyD3YpWIkXnSCS38b8zJaXrGdItlDxpvQFILvrFW9RE
nMgWHWMyoty0S8t5YKuXIvVvsYl4qrTnsExoVPWkN5Ux7S48UYyWRI37i2e40a1rwLwBuh75sfoI
q4ZOvK+cusXfytfJ2qwCL+R8PUU8uuPq0bQOp5myuy2ThNqM+cTiJ7PnAk3GyUZtnzriPZDFgZaY
8dPgAYD23Je8NoFRXBLDqMsOtTQ//ixpEtxE/FZ4ctBXWDKhAuV193NbO/1Tn1nnSBgoRSghJAJV
20MtixYCZiAvBB2JapIKrylW11+1Y96PbwUW7HNp5+cTqO2Fr3nPzJj7ldvOO8ZozzU3WLNWNxVT
8guUyKDFY3hWiCsn844xV1t4keXC7ZPoS3sTnf7O2IzSlUkqH9dnlxmznv2fEoZYpD3JIdCOp2RX
eiLakvw23213atcEYFy5uEGEHFfufIZDfhdy8SiIh8wMQXlmhENGjpSsruw3twd3SyqUVbrbeQcM
4eIub1ckftCO/zgLohJLjzlojYNzTtf0CjRhL4lmZ6WgK7aqYALnahvhHXczJCgPNhdxytt3xW4i
6Mx0DfyMVzvCIRLEgx4kPWBREtL1fC1nfRwrfzoiIm/T2c+rLOMOlAeu1cFrBla9pUi20pSnbp/m
Cc/O0UIA335RK7E2ZhW4lo29X7W6oslCoFeYNbdifu9Mi6epDiD3unR0dyJddmkp3v+RvNcVFKEu
+xQ7X2+d1YzWLEF3sqbeHbbu2aHASizj2+pwimSWZn8V0bQIL2k79OwH1QxLvm72Hg05D/01HkWc
SscuRbO75bBe/KDMG4qXr06tuw/e2+OHuhqMzQfMZy0FDGfhrMInn+lPz1Z8V08hhx1o1gw7ScDT
m+z/AhqXTFQrNMtyaSAf7D5YsJOxQ+ei7dH6vtCaREBvSeKJWk3Gl971jFNe7K1YUDdfPo8hE4Pz
DW2m6q05MXUS36HR47JiUsNuVjYazp9ohCCszLrmNRmZTTuuG9v4gsYT/WfPWVwzzUlYGSKe66gh
0h9T3jhKfGy+fmQZHCMesibJ0RsQOmbdzml6RL0dLJyEYmuiReIatOowk0CGxrVEGcN4Gv22c2Bg
LZ4Y0eHcPNBNM1ocQ+/kRd/GP61N7xJqrchP8ewWyhWof/aGAKmMXmAT8Bj9KbHDByu+9Nyrs+nJ
3jO6iRLXlGIzw6wEPgJc7WQujOAjHOTfq90BVYHOoTt7qRvD2eA06HxaJWtKIhCGAMjpPGJNxauE
+zuI/TGYHoZrHLW27TZnpaWyfRf9NzZ72JOty2TCDHcUNguAi2RTWUQIVyuTxhIESLoTUPajdnz0
VAekDX9qq8fNSnVL5LrVgq0ex/rOI1mnHf3c8w+i7Qiwqh5cGaD74+jA2DG2i7PJT4b3K3FXKwm3
h9WU6PZHdE+mZ5vNI1BYR86FkMMGWEHwfBYQe1ws4M+Ak4pGJvoPUnCK6uOC8D+gDGlvwkWL7W+x
9FDptnR/FvkAnJl0/PqieT7Rw/KgVt9gUfNAH8pj4ylQRO1mfWwKDpaV7ZRh/+EsoD3dZkq7Opo4
fc+8yCS4f3UTZtNRKPy9ocBcgGCVHMYUFQyqTi6o4Fg/lGASzP/VtcXkYqXX+zZyD2Nc66NTOH1v
8mg4x7Mze7PujDtl4cQh3DHhs12jZH6jn/8a96z8yEfJrZ3FJandACsgDy4Nfd39xkIlPoDm/Ikb
KzP99I+RFfcAExAkIMhuZfhdbN4493Hwrk73p1ToueH4HB48kk6zQkFNTfTSfw5GrGMRkrbNQ3Y7
dCLOhQxPsyX3GE0Una+uJFi7FsI0InNrkZfBC1Qp1raKv6ZXdv7h/egFCXh0dGfZCuuPa6Sceg7N
N3hkXt6p9/4HTRNhfY8YoJNsD6csYfUzRJNWNESl+aG0a5KVTgPghuh677e5wg3tUeyiEOfIWD/2
meFy5ADa//EQrlBcvc8h8DaU/x43bEAZL6peAracv5HuznMJtfoBPb2sYzK6uqI5jBilflwQFbFe
ZVifaK82b03Y2d60MRbKyxEgrippuqppjrYmo8s1nbGFVmM21QrhOx70d0oR10DOs42NAf3XTCJe
h72+FEBsAu4hCWFLXxIp8KLYgtck0nOZsNKGQgaX8GTbDDibhm3xJ7r1HEzdOuROE6Ie+2zxCdtV
toDlIlwPzkSGpA8WHmHGvFYj1ZmBwmwHGcqwd9dfMg3jPPVE2G49SqsQ8SBw9/DmGuRkHvIOOQF+
qa6zcYoEaWTnLxN1b2G3oTT+MabWbw/fhBQS7OK3EUz214Vbrb8HKzbB4QRVvRDQwt7l7xAmlPbH
0G3qk5LkUePkOGvuxQ4frxfufU3e7ZHIgRu2dsImx9cmZGTofStVRp5HqyLE8IRz53HkCIt5aTjA
pHGM4DLEEEU7QCA0CWw3TV0YJFVwlYN/NQhrS7N9rp7cA6KBO9SCYQH+LqIe3CdZRhbJY6dqWYVg
GjilimvIq9+lQXesaqljoSWPDfurqcf0/ThObh4c5slNywKOII2/84VmmnLWcrjvxa7KRO52A8FL
QGKf9hgFkMSxMkkPx2k4TxvAmW4/WYKRnzEhif369lRNMJjzwWsHSBvBfXfsuXuaadj1yGArd6jc
EY1O2quDokh12GhC29MfA64i683Maun6jXkoo3R2N0nqwsFydTKXu48Id2sdeEQo+RcKfeaSA68o
hb4lBDUxOZzn4lNCDo8yzTZqAKNezsoo1M+FCieGDZYRkzOTk+bRQFJh5ug7JOJ3ratg15vkxetd
b2W7gQNYMxrzRT2GbyNNsaAcaru4RNTqO8XXZmDRLdBqO7Dz6Lhe8ms1BGI/qtOnWQ4+03KRPxFY
64976HvSgEf0Vg78m28oQ+/wW0GhvHI1yptFD0kNWTqGean7CGF6C8pLZwTrUHo+FX89XzsTqsn5
DJLfy3a3Bq4GbXC4/SqUeOa+t9UcU47ZIyCw0bNmcVAVox+fuvdcJAW7wluoF5XiYLZIEW5uLmNs
xh5dXCYnxqg2ecM6VXHDiVdD30o/yJwidhAy9SN7m/j4NXisr67QkCucqItPsWS/lSNLUZkWkwkK
WMcYlrFD882i51PgQHprQA/HnCMQJI/R+xrcK7Pc74dtqIeW/kT7eiF7rUEfbhx0KlT3wRPBxyZ7
UaQjJIA+9kgc9WgP1SbLzgehyshwFIXz2X3BQ/zz/OkOBobNZZ0EjdR3J/7AvqfX4u0I5l69Or7R
RbctzVHE6x8yY+p29eK1ZXL0nMpRN4qE0q8KQm+GCfgt/AqhDJ0R/m+npVtCqtECP4CzF7PNVsEr
xGRJQ/KVZkEiCQufdAyPAA8vdl61CB3FWzh94XTJXvBDx5urM4RtWby2RD+7ESZsgL5pCaBybV55
fje4NdWW+HzHLORdM8Gd9PXwy+7yy9SMY2QjMT2k3awji8fAu+SqcfYMqh78Q2HEbHornOsn+o69
lDPOkvtHKZiOrFfMIw3s3mEs761EVdNpYB8aIwPWL7IK5d7hHoOQX78Q1rFvc19O/yobUex2BgIX
05XQCesq/tMvhJDCDmnxLbfrelzdlyQIYoyNOD9YdjvFBbq0W5XDJGnKSm0Wp6Pdpc0HzWES6qYe
Pd+Hg4aDIdF7X+ED7//E+88Rmq4M3wGqwz+xzlUyxYAZTcfiUF+GGr7p3kNGMNXRkxfS5Qcz9KdC
bjSFaH/4676tjEkAfO9WgD1pcDeZPUYWxF2/YRSQHh5KypJXVzhWiD1gZziWgKRT7FOOfGlzWKdI
I/0+TQNKoXc3sLhu2dGr1W8OXSqa4k0j8ZhcfufF0U7V2l6trav8qjXHwjVil8r4PQfJjd7WnjEC
WPfLjJ1k8Y1fT4vdLiRtjZaOo8hK8fSTM9hQ7sRKwDIZXY6TYJni8/ZMBI3qm6m8WYub2DIMbRVV
rMs0ptOoeKgZlMKv59PveDmBRhYTb6j4+bhi7/BX4g64YV1emVpqoElTRR4ydt6gf0j4oMj+IeF9
Cmk7Dxbfi90MGuUt0t3pAcGpoHZkp8060KieoU884UGbKcOgMVBD7Ql7gT2tnSBgHfIAMDrfpsVn
GDB7bTtrRYe04RzfQii5gysHYLX3H8I94y/bB2hXAtmY575HKeif9BKizrYrzYsj9u3meLYF71z4
HvlWpB+LOVmZC4cCQTzXot5ClHbWUGVOcEl0Im47cJj2Cm4mwxEIroIRtbrOTM9W/qIdtdxkranF
0TPXDqAZ/wkXQbIqgpN/bdsrg2XMY4x5sVugaXOW8CcW0UAyLktMcr45g/nM7rzqhyxTpVL/Nn3H
grdtT0UYPfcbzl5dWnCdHdI2bd7y8rzu9zcLR3acPrILGmKmksutrMBpa60KZPNCgribkK7tVmUW
KuR4YPR98EGGzH1WJeYVo1Uk5FMyMy9pTpU0HjDr10WxUZC4sRF0LL0Vc3sXT2yNIXH5BFoE6x7z
R7E7XkkkxTVGOEsf+REL5QCS1dwuhfs3uxcPswFso8iODfa7FLdNns2+oIHqowactCmZYTT0JlEp
IOvJKFIkXEZRyqG4zT7qX4J+TMMx/by1eVFnVSSykzTfIa08VucmUkGXi+OTFaMuvj33A4xORSe3
zEtEtrHw6DYaof96L7FqhhzcBmPuqceUBFSQILCRjBvjCWi7902WP1HyHcr0DHbZinyWn/M2+Jl5
sSK+wKPnmQCq4i9TxCQ1fCGUx+z/bvisk+ScLsmAm8LlZ1jn8vtEIQ87GZRFrPGluqkiKDHJApUb
XJk1YuGHWLkc/SEOWGj0w1WsjA3qAVh/G5lk77LXvcIlMKL0WX2CRYH3Ak85kd3bJTeIurwyzzYb
WitG1sGn0ZU7NO0oW2XOcZQ+OQcQu6z8N0lkY6OpbiL6wDxV79wJtD1izKR6Ul0iJgeZKp6TDFNg
L2+7WUOvYiOEK3s9JflZIMvHFSIGnbVXTRV87RotfpcpSiOqppshMQOW9qldcmIhn0kH749ZksTp
1w/SnlEgPf9zrC8QwDPawspVFIEN0Yz746wAqNe4voBCVFFWVaQgZL20xu2YZ37aVqtb4WZphDqA
cKUo26mUg/NxoBSmYWrT5p0icEOL9RTYfLPJobZ2EOrw7vBtesbsteURVEJBWpqQLOQAU82/aMCC
N3cPCNZcrahcKKj2GVzKPiTRnmPbgMXih20hwzUB1QhodMof6Rl/uPhzZeKTWKYaIGtqXIwVXNPl
mFziq7HQt2pB3Bej3393jG8hlyQeEIKS1FdTaOiuygZ45lLIZaQDUAjUAIquSn6Mz9VOcD35Ko0j
s1Inur7AHlE3sqKeifFcruuBmdHeUkoS5qfiiecyCVRoU3OLq1pYsr5oaVbjsbR7soz5LlnXOFw7
2ljZT67SOK0TLqmPtloNFAeeQ1H7l+w4V9b+KHgA1Jt4pepzNmXtmAc8P81PpYvNhCz6tq/7+AGp
+hS34wBcf732COcNXIt89ad9vfVZ1wxwJ5QtfB1XPMNjt1qD9Iwn2XR02N9eBbyF3j814aQMlXmL
FzzygAKU8u6XqmHIMTFN26DWWhWO4Qh1JVM1Y0HYMAFAS6CE9pqyhaZ2wUZHpgsGDLjV54TIK+Mr
YFmn933fSbuHCLNXJIeDGsDaMaPMcT0YPEBvpy1ItoDte798y0uSuLMRjTitloWJ670zTE4Qj6Tn
OEqKNqUhbUHc3yNkVjCNfRDHpUblnqZ+Y6z4d+FodwY9ZWZCKyS5laJe2d2xf1E4MNTxg34KqrV0
nzWQgJk93DrJFs4j6oEZU2rFQZE9pIw1ptBCd/eo9LqvcmEIT9Lghv4gICPV0yFmfQw6WrCd8Ss8
JnkiNeqhJBQoZVdjamZ1oOJuaT6j0FL1DfxK14/mv18q9hdHJKtahgGENEfuJmQp4TVwvdkNdwCG
TSoXSpiYqTORtj/08sfJBxb1hKggs+wCMqL8mq3VAHuz5rMZ6+KlJeb1sTX8R+x2GMyLCblGEHGo
3r0FDD1Czk49RBdMtcwwhe4tqNojM4Q0w/e8gu96hX2Mi7IyUNBhX+Ymm8Can+r7TWeaRpiZ+3zW
j+QBceJ6wyxk6gNrPhPm7INXEQ535fvD84E0aV+KhnPe5/O+8E131IHIz8SvCuPh7+iJ7NGSrU42
4Leb2a4XXN0dVLs9X45Utc7PKDnBfkV67SfXzwsuaBsfJa9Za9vo5CYzuMnLxnvlULUqopOBWjjY
oUl/u9RR76TIfzysbcbu9BLtmwZI7MRugihCcCI3xFo5kSbonSSZQINdrJM5H03BPDHPHQxGoQCd
UbvzezSbnarnOBNMFfOxgqksD5vPnmxIJd083FnziJoXOX4rsmgVMMtSwIV/fpZYjj6B6w1p8txp
pq/53s8Tej9yk6H2xVSawpuJ1nxVSVyHxMSDYim3p246uD0yqETTsor/BR6ENtvYnF8YA6ua3PHt
3j+NW1H1s1xFfFfNBbzd8+nNMSjYZwdj06oK62cawO0i26SE2b2aONTZRkhrtCNMY9/ixV1K0Jhc
bBg1ehWkP65UsiwDw1UEmOdvvMVi1eI/aAv7FFR/UzsmhhuPeKS2tdky39J5SdpsvqaVkP4JXNNW
k62FLjRqgWWmq81CtEYrdWF+9oS4W8In29skPwbHvOJOHjdWqoUlo+3p5A7fF4SCaqJUWl5JDWms
D6bl2C6J8kY+MlA2RrE3/ZGyb/3nDZqb2iRwSpMkSFNGDFjQBrs0tq+FJDDLYbQ1NSOiYqTI5O2A
f3iNlKGgO7HW3Y49keT++hHdIY6GPI9DFxygMDzrmrPPNBJuHk3tYe1ZBKid+Be3XY+xtHrn9T+1
KNdUI/NCgmNCSzlvrAeFOcDUnlYEH2vAnKdU2MnS2kCyth4MOWVkbXY+5v/quxfUxIUukJOo21Ja
r5IcBuAhT+p1fTJ1QrUfEJ6nXD/RzO5lsHSwg+AyNJgXU9eIAGTTyxD73+bjXaxzrYrapvZwVXkD
PWKwZaPNBRUyK6ufUnAr92VVUoo60aoSfr/V805YNCfArWV0LyfELY5YcfrdfkyH1rxNvfqGCeVQ
om3QK95pzCpNCcIUKi6tLix2UnknulAstGhaXB9Bj7JHpis7uzQABZYPI6obN1ZwAsVG8kHkSJTe
2Zyg5ta3V9pieA4D2DBXzoxuZldgfsCQWdeXGn8GiKW72rr+zVW1cUvpbnyXCAtYnwat3rcY7IwA
06VNumIhh5i5ezCs/nL4hC6a+cx0krymSODTkUDFMhL7HI7fu72jx2bCRsQrAGG4il4eoI+mCqtO
1Ie/qncYtmVmnIw6ihLzCx2TIygLQrZQvpTmGN3nfhZ0Pj0WOXVrawEBzFDo6Z6oPtI7FeSJEEYq
RQrDKcArnj8Pve/tMUTVnE8DrIaKbEe1XSy0DPGLI6/A/Jm6Ri6FMdpacylOi3iMen+vwdtR9gFd
EXLr6c/K2L5x8g77kPbdLt6V4FgPIlt6gnIqHZnkmW7Fcf4r1mW/RbYsm/qh6yuzeJtA+kqPDG1a
ocDhlMcSGElEwZ7gINLdILxq028v0ZonZ3LstGsgzidXswhCuouvXRxCmGlLnnKx1suNvbGLfiW3
QrxTS1XyEpydA4sVQ2JSC0NvKaLm/ySKjz3qXjJgMVC7R4z9vzgm86PvqtQkLjYGRPuE/p7wkAmO
oiSAeKh04R6XgPsSWdjNEiqa2oj5Jo0HTYSRuD8Bg6YammzVn+Nk60QqZLS1AOd7qL0h0wqAi4U9
EBDFqW/oshMP6hLJ33sp9U3em9w3rE5UX/ICWg+Sxl42rLI7VVgNpLRPTFwQKRO9kJ3bFJFtguPN
QhHl9XJJeA4+5ZK5eCYjNkQDYUtnBXYCOuoymR/i+liFeLbju5ttW+mQwbVh2WAQn1ANUSBDz1eE
ShMpyvHJ4VN1/5HFlCFJUdzL/q4MV+vZICbpRVGQONqdnr72TGkLdW8sxssF5hHWWJ2cowngI3cn
z4fEPoxsNZ6ZjzhDp88D0MnPnG4PuRJPadtllnlhHR011TSlgnwxFvqNFOFMHkmASNAUACOJQ7Vl
71FcKN+VrBQmk2Hocee5qb4BWwSm8UF2JvcYDse5q1Aq+LzvmgfeFe1cxM92iXOUAHwVmdFZnujp
PERjjKb0ybCdXZ3Hd5yIuUQivV4jrsofdV6akvlW+bsIQ7Yc7ltK3+aCcpTnKkEhbIEOx7G1mxFJ
aBTswBvupKcq42dFmJHDeJUCKxJBODG/9h1qWkKOL0eJUZPuF+3FNKTEAzvYJW4eA7qqJLl99xKp
MwgwnGVfE3VebeCAS/ensb8yz3EvQL1HVdAibNjYsVysbYbXDpaMZI4GIWcVwHDRdCqzig/m6MmY
6ki6qCeghibO4IQKUPmsQzc1VTD9IcsiiHrx9lmfF8a9uuWaCZTXes8XggD02XXOY6qCoxuvBLCh
Nw12LS14z7Am59YWqRPDx3Fp+MOb6/dygWHHwx5qaqBEAN6M3d+C470WeyWAuYkZ9yss0L6Ja6X7
jtuISJIU46NvBce7O90gXDZv6aj8fLvqbph77fVepzEf8RzTfz8imy3hupW48Tmh0E1s+W04zgJb
wo4vPXXEAI/M56S6riTF8HderXT70qImuedzOU3xB/zfLwHGixEEylfu8ySBKg4FGJefNp4m/5XL
Vy61TbtSpQV3yyQ6OoxueoLQub1q9jj6xSv/OYQH8GwwPo54HdazkxyDy4yKU3lxaaMxVd6wopT7
gE7kK20ep+WGArROq1m2qWBahrWy5hV0Az/LKbUcjPyXg3VUupS6hY4xsVrX89N0J23XqfKByXC7
690dP7jvXQJxAPwlbzNXTY069LiR0jMEfProksHd7Od2x7A976a0G+XRGxzxTPKxkJkUxIRDpZBM
nmxqORpmArStpLSElZb+GKOxcL9VNot/9fBSebSt61RAiPLYGq5GMGE3vrdLLXNzzbLBRRGVOdgt
sItv84oKfw6ihR53H+qu/xXHDaot9RQwReoe+RENnXS4tfCz7Q9KANTrksiCsF6v6GnxQk/tls6J
opdBpwcjvpnoB7gXn8799oMRj682+jegY/PbGt45SvV3ViVdGO25n5qBNIyXRAdnOaTm8fsKPgCw
nVfGaakhGz0rRwFd/UuHNtbZcK1FtzZc5KGcXBcHfJHAdgizBWTqExRvZnOZhUYew2Dc6TqBfjhr
Ow6QeITv1mrSMWG3T6vrsr6tiFIe+xHRqvuJ5wZynjpI0ECqTg8owsIakgY0S6jWkmE5JnoTN1Nm
x6zTH0aATgKSyN20LIxA8jFpPuGdKSvrmaqkMthvUnCvx1g3u0xb4hybiTyG5R6l0+J0pQwv9gLR
H1oTMD55s7A73Z9eQbqvSuhyrrakO8feS49B3AhR0ALWY88SZXql+IOg/hQI79/K18gQ/aOoqeRR
Ca5ZUA/pZQW+dfg9dZBqr6o7wiwIX61+j0vvRhZIPyu2rHTFLxj/yTTqyz6k1x1XgtH1nw2tz/yl
vxjn4dUqPpq828iKYBfMTYS/CDLK6MY+6YBZNaMLq7RcVXt7HGysHtQS2YITvPfc8mkyrAmnQ440
BmaCpHFEZdMR9/GMoEqDQYPq3qdG4MjrvnorAAYULfQtQm8SFwRw7Tp0cEiDALLRxr+8l8IvM4Ca
0PSYXOaaLGMPL+p50u97XNBNjdVLHyKpRVY37mHsKjUhD3tt5k+K+kT/Pv95MzB4EIj0YhggZBzs
RahMXhUsO1LlXEf2DY467ShZO7zhR9hwLqtaF+0FOL7cHL7ycsPr4LOBCEZKNYesVEYq24KJWMCW
DXHND4Z5e5LFeSJFvXYZzTFNEWUHQ3eYcg1E3Ja9SjxK27v1/lsoS66X2XiEZPUtKG4KNez2etyr
/za6W5ypwnZxXwVq6MWhi7Z8UYitDD2TZnoRQ8XbRI47RkABZSVCVVeNoHz58YJdb7jfIzI/BbB2
ZPTCYBxUisIPLl+XEBCe7lenSGCeGGMcuo/29fNZibRmK2iiu6/YqvfCJpnC5xb3c0XQKgZzdc1u
jnVlI+s+wFGiE5VcHNC2BXliWh2IZLD+PC2v8JwxS192n7pLPLXpiGmhUF2qyFqL8ZD0M8P7wCQO
bRo4F7Diu1dQMqRzshmwGcJeGLuCa+29SKoClBTM5m8w5OZX/aCepPbj5M4RjucXXWDg4v6BBqSp
LUBiTLT8ICzLUgxlp9+314dhG3OumF62CC+mjbd1eu2vhF8GlpxuimqTnBRn+BFH3HMtaMSpg5+T
BhalkijkMn/qxWSA63fYLDamNnsLRArlF80e6Tx41jPFAKip1gep/ggcT+a/foFGXaP4UHTDPeD5
2t/8b00mkPPDBHWvhp7nurDgk95RhdIm/OPJsI1G8uiBkicJeBGNvhsW2uNuJpOiBt+L91+7FvDo
jYSV4glBBqy2+o+IGOkopOCsVKxL+iOYGnRH5xo12sRrRuzCgFWKTExfMAaacnT1koZkKfOz6Esw
zW2dyKCtrN5FWLds8oqlxJvqXhNhNBAYLW8rXE6LSzyYxBkrGXMrsceRSaA0Y808jjDUcK3o13hW
52ESz99IvYxIN562xWJGX1okQA78EBI+bO14Px+N6ibl2pBuVvASQhDKsUf5mzbRLaBCNWCFslAs
Bj+aw6Za5VBLeAU/St7Ifn9L+GFbXYzbSExXi4A8NYfJU2F+PlOGUIzh20PJ2rrghBDoyXsJboI/
3X4neT4oOAOUZ7ryEA0x5QxbXiqszEwxvwlIcEmzIFKEloxqzSRCb8nWVEyYuQXeV9eO5CSJlYZa
/MmyQoOPueM18SCRsepX1EQiLDty1LUw+bLe374uKdGApCFMG25Ew0dGLgDEDYXuneJb+Q5l+92g
7k2T4De9169fBaZSzj/Fh8PoQYIaQVH0YHQqmFXVL5Yi82622n3DNUUTBKsC5MWwtafgbHDeTcqo
Z7GGYfLPq7R7fMp1B7t0oj6PtdH6k0c+4W+utWobeMmdcjI4WqaJqRqNaktCu1y/P4Gs0/LLK22O
N2grkXGmUIKgNfaUzvK+jASmZa9ZErkpDXj00r4QcbcjFTlb/3WjTcGy0NpaL2sadGygUOc6HwsC
EEddfFTzGFC6D+YKnz3C6DGdZCgXgQIIfwUMwiy+Et3kbUjJBPkKPCGn0vjY7TLS6ZMSTgaLc6NW
fdq18VQtQXPGywJ7pvnCsQGwkPu36wmP0muy1toKn3kiQsUVSONFi8rMiyPab1KIUXda0t38HrjQ
NsMV/bX7JbG4dyH5Xwu0iltCTj44DbFYGVbLcWQGQMoS04AKbzM+gWH0iQk6FH2C3jLfeyiNb/mM
vWsARXtFPXgjpVy5k2bK3Xirt7wosZHDw+ttNX4u5z/5l335Dr5dTB348ebUj8ZaiKdv+wfWthVS
QkrKUuGIzLbc+Iwo5uvZVOApJWs3zVHkKfgHb5XdBGRM8QWYpUPhAfzNmaxnTegnR2OJzaIPFlia
T1TewkUHWPEPMnFH/pFmuZ22/TNoMZr6hSaDiNHzZ1XdtsP4jFjihxXFnstbk1mAUWEAQQeMmYVd
Zigpc8YAxopf4FK+ycL/ncUOq8BlXtpQklWNd76gEubl/KxlSPw7sHvuKzX1p60+ui/6433LL8A6
a/jIYGfFzfJdXRDtGtL/sX+E2I4qR4zDaT062KmUYqpTczqJhfqJO/fj39+eIao+2GTrvR2do3FP
dJTtOcQNRyoAUyUCe5EqTfF3NNlXDUZ8p2vxmqd39YHlneJXS7BDl0lAsvmHhy1p5htucy9BtNlm
jkKO+9m0W6suhh3Q+vVtof3QlgJ5eEYB7dgUbnmYpjiVEouXaVTrdo4dtlYJqD7kLXBsybyVAmmq
sXaVqtdri1rUogKhWoTuxnPd+7gwv90IJcmcO8TWIGJy1OZKD6ANx3y0r3Pgv1l41H/NmV+j47aL
dO4F0zoFGqmUKOxwoeSnMldB8Gr4/O6FCBHBjsMAITJeSUZhHWDqZeNMWW9Zhf8Y4jYcmaokvCzF
o0irSby+LNFe8JfhPZNRqp70jVx+1ry30TnhYl6LZq8tUep2DAoIAo0LdACFghwWC7TZ0n1ENV6+
SsbBh0gmvoWPMu+VYuhyrIDGp1708UjGRuRbHoyCBHw4GeMY5oZw9XZatfhAb4Rpav1t4JhNo3Jx
mJiLNfrKWGQ+ulE6rlKPKcjnvjrG8sbSYEioVrc3kXmqPmNKGLXMMK7Qen4fW2E1IxDKzfRPj3wM
yFcSypsF+S5VKEmRnZHW4xprxkp14YQZMCkjXq7LbSEPphJBxd+rD1T4QMzVsWes7GkX7t5unbT6
SHjMZvokNKc/qBc0hZ+gUVWjq4TCvhayvDkckjiRQSDIhoT87Gih7T7S7Xcxu5pSpnONDhmC8zPW
BLtPw7xW0Y9r6i1o54wEq0bjXpmsPM3O8GojkxvZzfieEF91moig2J4MI6KGGipKhdtliwofuBzl
pU57h9NaqzGM5Hd74DWdNwPTSeey0g1HxHPQsCEk5b8gBA2rjxguRZD2jYuRQFrGKhzC2LghuXTb
NxJ5466kyXSpaChhWtNOKU3sfqiR4SQHJRs81jrnV0DYnOipSB36o6qdkyCqDC4SUWjtb5mkdTGq
NyobnEdLzrSJHJ6rhuNeVPEjfL0UlTL5ruR3HhD3dmTZvO4OwygpfIWM3Jcrjnw49eBODsy1BODG
xq6i4JdHHAtMw16JzvYU74+yRE4iRMgv517fkQhO0MsYyfcHK+0H5Y/oRhrQr9aGhHvwBBJHrasJ
mec2cyDNZIPXgfzkZylk2uV2mZcfYxVh1ulmnoPd7BHwvm6/JlXGAUD9A3SlXubBU/ksUF1IyaAm
yjLoYI1hEGCD/qV3BxEaySLDLoIOTrw00lGvHVhk/GyRDEF5U1jLZjLFB2uuGmlcKRsAUVdt2tqL
3D65pqI26osaLHxd+nd67l4+sHUdcpl1yfoUgwZhFj0T//0yWBB/vj6ZKKkKCgvKjxKTTW6lCQW/
5YZXOHagR1VKb9D5RwmNQXkC/9PxTQ64nhCsQSf1viKDyPH8p8cjoQ2ZfgWq7aQdU07dk/QJRYnB
KI+RsQmw1wtdEh7WJ76PHizAeNHdbXV/6u7XkgPI1fSJotf9ogUYd7ErJRPIC3HyAAdcS6+95zNh
nvnHOClmzNCmhWvofyLMhHORhB9XUgZLKpuA116MdrB0jIB1SEIvXee+4CDWkbNKcClLAqCbNev4
/n2wOfEbh65r9FRZghFgjlJRwSlyWPPLsTfAzqG2Kvsp0F8fPx7NOyEOf2BmhK4HqIxxrS10Fjg7
ppgvcIMS18ddCor1bvgxRbh6xApj9+Rl/wY/3NxJRxQV4QLJoyOCrnwiCKmdAWuI9LBYH0uhf70a
ZBjosssHilwmSouW+1gpAbIJDKCRjtr/Ne/MmxR77RLcZdGBZWVoRIdTCYZpqKj9haBI1odxwQmJ
JNWtzVxKiAKsEmgcmAmHwsfhk1lFMTmfrNaZNxptYTOT892jQKNQFaAdyx9IpnUpruB0/Xnx4q5r
CfecQj0dw1QOYwTltN76i9wJgDmsvWJ062c5LNQ7XSUfhw5hoGO84QKss+puU6ab3VJxoqQkPi8I
873ZlM99cmMUNw9ai/Yf5gADJqXV6PY03ctN6Ec/PrYlKqpwHOydOz+XnlmQdm2gmdIAcX3NTGN/
+8W35nvFH3f8r57YMmKNwBGUHM4Z6ZD/hujNz+0lFm7EMaPD/n0SOC2yIgPecVSzucwH3JPYVZ0x
qgRRIS5CfTeFzse5n3IZ+6qQ/+qdA1BaonrfCNDPcYAapn7Uy320S8roHt0RSa+bfnRmT27HTwkL
t+NX84D++M3CqiGc7CnVaQs/RCizD2JqGgX7mFyloEBF9wFCHNyS5PQ/OboNPt5EhEfTyNLuEjM3
1KZMYVrQozOP3vkVl6HIFslRmimUksVqfhdqvgbj1ItA5kuZ4/i3KNPfxtcOR5/XL0UI1GkxvfAq
WP/yOb62sRPrizxKo14ewoi0mwiPAzVYFdD/lupQSftlL+x9O41GBhDjWQy29Uc9KdSZTtEEmDbj
8HNLqgaOQCgAr27ChpIhSx3GKu1tR0vIZbO/fc0+/awPAook4O86eZbOfH3ph9QCmTJh/Dc626yG
7bJM80cu0Mqd6eyPlKDkWpHD24brpBpSs/uN8Yp5CIKeBJwVX1Emj5XIn3RVY7SRJNlLAnr1GTgF
joGrDD7EdcwZJPNE9bMkYlmt+Uz+yoTAigJe2PhpC6Mvrwf8gYHwpQi5jShApXlKKKB6H/EO4K6F
fVqFzU1lD8RcERMuK/ebcdH4iMFrG9BNesHYnUx26wf7iFBEEdpSsqRjYPsMzIx2JJNb/fZT3nnd
ug3tU6bnbFy3sHXH0tjos5yhZVbCGDQ0OEVJ6AzJ2jILljw27H3K3UrWMi75TEfbq0LzaqysD3CH
J7oThQjZwzjSqy3KKplSttd4G0+gQy6FYkrwsxnNxH2pdzIDxw3LkNsXzpT9bPfL51JkTLclTGbO
u/rQ0w67+m+hpN3s/GZcPbz7BIB85zhWdhDgiv2SXbFzp/yEUBBfnCco2Y6SpGHXAxESlHGsgEcr
NYqnqPfTNdOooDbMNW7ccQeudadkDfpnqelgjWkT2pFvKwJT15HqnyiC4QDJA7TayXPwVjHofFIR
VbsI3Ya1tKo6fXxyY67mtp3KbpQEz5FJwUgPLahvGZ8GzpzEOCv6UvpylAifwNpgBP/p5naWlN3U
2Ep6y5oelLkKMC66dn25XhUp7JRCQtxoXWawYiuRxxpQRLp9RHpNApRIvrKS02KsHLsK/y9nzmQg
vNFCGa7NrQU4AYkhUcXb3ZlxuCHpxvGR8SVnVHcPfKfAHQXGaYWwyEgTOGjzvNm+2prbvc0ceJnV
nBI6N9NuvzX3KiSynsveIsoRshvZE5SVHwo7+8BrvjzSsd+sm0kp1RqUe131snvf03pL+Z8IwfEx
S0hUiYb737PjClpY9cVwydsI61JlTe8Hhb3Hd+h2UV11fykfTidlR48mjRjHEUieoGnTsy+DO5mx
qigkCWbZBR2u7SzVXELWvtrVnhwHyjcwOfqN+IfbjZPdNi/ckG4oxy81I/bN3BU34/s222XORd5H
cibRPw0oSrU8q7KZZQKKN6ZtR0B5NS/KUvUKXVM9v+CDA7+B1+SZVegXx7NGf7SsOZRm2N3cVqta
g7Aly7AWpe043xJBHNQ7ddn3O8Ud1XEO5x3+oyp4rzx9CmK1l6jepvtrHn6FAwrJ89f/Rf1GVxsC
u2aCRyUTgzcENlzcAQKfHWPbGE/UIElPssW+2MkWMbUhBcS1G5pr01p3lgxnbhsCl4xTviFHT8Si
nBjdyg/j43ZsrCkEQM1gnxkgvnjx/4b4VvOUqkPupEzwxZnkYclmKnHcQoABAJONHY1nTLzPIExa
CvmLelCzGv6FAzkBFD2BD7v2tUDo7IMui4Y0gKrAiy1pBUSuIgIyos1vtNvNeWWiEiHsEktIFGHC
Ltv353AcpG/DPVnekd1kxAsyAkjVV3I1wqVHlKLOy9Vnl0eBcWB6RJmggCWPQMatHAi7lDUPYOgq
zebH+8CVOg31ypQ34EBlCAJhsbMEX3Ki7BZTNTVhXnpjl4gNzETm8XLoyKbJCffoZ983fhPkr1D0
UiGw83MsFnerIe5xCGW1nkz7+Fy8iTWw5zD61IPEL9P1Wg27nYwibNO4Rkv9cAQX9TFadQHNwiqn
S1bADOwRiX1+MD9tn/hpp0NCxCFmfdZ9nJ+MugmGWZlXhsWh6VEHCbNwJf+vOc9a8ugF66+C/Uuy
73JzrOeZAAr5xiB8Zv5xP7oyhEj7TYgNUsAGtlJA2ZYISVT5JKBtVOVRFoNDYBeY+v5l2HzSm9BR
FA43wzNKkKwFrIouwspNDRoqA0QQnJ0+LhNan9IxUYIrip6EaE8Dj4EBDjxYaVysLAei6zIg1vj2
a4kAyF7MSCBpz+VtGRbQ1c50mSvgVd0PGhiFlwx2n52Abr2JYfgNJv5nFOqhCZCLKzw+tQqGKCL4
GWMlZLs8NUOyqX32S2/lRcW1KSI+m6LA2Ie5MAJYootTvbzzccy2ieYwj4qScYT/u0AnjFTxPeTv
sZEWxTx8OWEjc9JwPdSUqVuFbLFlAxdDAaFx4usJGZd9SpFXsFw8H+ywU3G3RTYfLiO0AUgj1c7J
Te5MPhiBhXNszxDMAqtOr4w3HBuF+/9gdPoUdX8V9Q3HvcE4zVIqlOgXBWGmw5PbWXB5T2raehj8
vzQdQKTrVsh9M8tSASuJo1rWnU3KPrcHUsd7rWP5FdYGPugXB7w/J78cHBXEfpvqOTqWVlU04ZfU
p+Li5na1+vkQQNCktLTqtH4bRr/mO0klCV7+l8sbl7mouXn1RkssklOQ8Yh/D+xDwaKKk8RvLyWw
k1pGXem1ERwzMPy046iylATLCv9t3RV4eynGUitV4IX28nUA7RFAQPjXcaH60fvx0+j8xsZxKDri
iMPvp5MgBthBBNyvAbLGlkZ6acWFDXmbIM7egGtvuLgla4080SBXqIccNdTSwqnJDq5uI2Z43biD
O4ZU6xtAAieeV7/6D1pCdVXYHmT+r2ikRh+/oz8KuE3az8Y3i5yPRYu3tL7EBZbNqaDZezLObynq
0YVKDbPMmBK2IakPlQ3WDO+9LeB4kLT+cKHgB75Ah/9Y3xE2lGYncU98AdCSqKlE1qhZZ5r9Fwok
IUAEn5EbSTVpt87VPYm9FmgvCOQspFsrKHmT5ypenxopMVavvsGkCSwavVH5ebWgnAz3wMG/Yw6f
OYBOurfhysd/FMcpVmEBTc0dRCxPMBOlTX2DEk3lNCZ4CkqM6UA8uTjRHM4JASuv5Z2WmHuU1Ovq
D/fXWhAEqSpAD7oNBt2jPzLuOzlg/leFLXsG3WGc/gtsao17tgZcLJcW5vtpdZSPqUR1lD2Z9rUu
Jn7nw1X0KHlSllRoEWItBakHLuxmgtzbPF0ltxirufkmd2Bn0vjXnCOBQ6T2tDQZZUwxRXMWTdKH
End42v33+/RtVUM8M3Ru7tmThTEigV0qVwuEjP7d/ra/d7zU8VF8jO2LVKmc8dq/B5KNaXWCsn0O
nmHD2YP4DOmlE3vsvT0tgl3uDY/v0OxrPA2Cmm2N1qCS65QLZP8QqwQ+aOcsDuYD+d4b67F7WRw2
+ZWneB7t+1FOAygIFYFosPDPJvlIatwB2I1z3aownduQF2Tna1ZUlU8buDKlFLOTes9T6jiAM/2X
JKPEzY991ovy3SlmMfsTngTk/n8CQuFxQVqFTkiWlWdTFAvqv7HDAE6JX1UhwXzmjGSHO9/l7+R4
i6MYhpnVQnGXJYxyQjemXCpuEcNvDh8EWVDk0jFUVCMU68Xop9nDwCO1BwFWltwc2tquYAHo7qGg
gz/2fDVTeIoARPz8IFh1g1wXzaKLxVqYk9ESMi4p02/jzn/exAY+tqqlB43YrxHvDX0it3IUv2hr
LR5D0wSPB/sgS4mcpZHACIyyEcRnuaHcdn/YHzjqz68CopnplDt6q3Gh1pNAISK8vx7YV++YTYjh
5glQY2g/jOr238AagUEYb38T9VItJvAtQxypaYrSC5PD/4QVCVnjyvH6Ma0VRjdBLkVQzvFBCuFh
aJbtl9LRzgJPChdLuZqynVOAHS9dFoU+uvFIvCrPnoKGz2xlcGjKQz00e3ncKkRNPHYRhx0nFIz6
uUix9LUpHeD1QHYmzBz6LHntfl6n+jrkY2mKALMh37lgpkLwUEuo4rL7sQjH9tB6JwkD9Xp87Nzs
PRQdD0UZ3LM2/s61vFua3V0kBQQAyQUi9M2NlJQQPN++ft6qUpXnYIJ8dDBrEW1nAs4PdfACl3jW
UvjuEeQm60tbbDDFMvvNOhc89HbMANiFmE99A4t6P7p/m7mF85aLQkBzJMPFxBaTpEUWOp4HFN5w
uJSnoTSifUpJ2XVofKATTG67AJYBeVGqlI55m92OOZuEIeQ0103cJ9ig0ZfGbkEywl9Q61p7kWFb
xtw7XVUqqoJ7m4h+380PnsKPGOymx0LM18ge8FcovQ9JLZFDxQci77zghv8Zea18l4NUQYlGykGC
Pf0cSu5ku8lfT8PK0nhuISJ88TppQRvxdVDCVUfGTmJwPpMhu+s4iY0rjUlE/VxuY5C5AgmPJpT/
OsQwE4TzeEDerkPnh8rkIBlkUO7FocyJW9yrRo8heIDHOXQLvovkgPnaIJJBfvW7uXLRO88RCy84
1SLb5PXAKEuQnlX2NABvrR+lEABXW0VC1qZePfeHNFr/f9RIrGjrd6kylTJLTb8cDcAY+JS0Xp+9
2fs6o2dAtXTtzbT31MJqUXLRANoRS2KNUWyoaHrZk98RbbSW4cdN+Jj2ZoMu4w3bpqd2vqQCkGYs
67sIpwSV5vxROW+hpI7So5uIoTLwHqbnyRfsURSfl33OOVjNjDeS+KNq6iY5LKIYA2oyuDjmXkVm
wrelh56pBsxACzRkTdI4YVT7jprCx2VddJoTyH4asUBli9xu86MFxDMHbHXmEPB0/Ka0SYPr5GnG
kjfsZjrodp8LjafAUkoeq1hQzDWbLTVXkOY+laEo5Jh4GfLx93vxNxXc9RuNcCSBgc95k9oseaXI
GBW+Gt2uwEQ8yXCPqKyAp9PXDRLWHdhwweIMnGjAgb3TfGYhSt/1/u9+3AwLa7YjgC9PrRPiyvZy
zx5mgPJu8X+C7dVxg4b2f/in1yK7NDNecICt+jSTnhtXDoWlM0wgxYDcDaN9N1epwesMBZvWHUUB
bPzZjuXsHn/JNzRETufrlXYHqGBmYHvPs5dTwWipG8pFix/pJpS6+4sSVPFvO7nAIIzN9KDdCGEK
wqKmRq6eGhAOrF9Dzs9f9LFT4GMc/07JhQfpGOWDfaetrcgw9/ICDTBq/7wmjeCdOh7QoHMgKFdi
O4ANfY5bmYUmO2WMGAv2Sfi9b8SOmuzfAFVmnfIxaXq88FGoz1AHGwN7tJSkHi8MKna3vFzvZ6GD
/zbgdQB8qjpL7wLfEpYZHz8f5wdXasumFGgwpP3RJM0Ql5MasW2qn/+WlrK2ww1vMIlTWo//IpS4
lMJgKQheNj0NLelAPdwZQUfxqBm1rLE0t3gc6mPXsMGA7OgZ4CyRw8dVbgo5WJ+cZtRj4q1tC+m9
efaG1GPUlLYWgOWanQmmP/JkCHDfSdANHIoPWS1AEZvQmhJjKskfErMnG7rfWuf0694Z2VGoa+Cc
du93++AvMoKdVk4tDOabfQAOA3MtPsiuCHJw9EvtmvQz2AqbOoyvGqkvk6JT3y+/A9egDpCeqkfY
K2t7YgXrNS3cHmtDN/paKyXQ+ucy3LuTX49C/CYppBj8fUO7h5EO4sOwzbAKGPYtbn/1oPy9FNOM
bkZylMMBweZOP49YbGAoYTlrGSM7W0dyfPQxA2Mll3iZX69gGTnDBSJqmcHjq31R2QuSD0lIVCQ/
VEeMyzXTOVw0GhoKygFHw06tzwix7KSWQ3zfZqhdO9o4tx5Tpp/sJBDyzufqUVgbObPw5y+kGysq
Ta4kXifxs1B4H+KqUqoW8OfalGW3rWSILXDu0R5sOFhbSeR499XHzLYEfqHHUYUYeicxgoKJZCH/
lnDfvdgXrkJOTAQFRdwzuorPphYqLi48yVDWMsg8kzPBOR1/0FWLSFCDf8DEKJhntLOGSvSMOvYt
BYerwMaOwipFJJsW8ZWzasp2ODHiMbd0IvsAXniYk7QXsKFGZuOxNFvDfAw4OhjVjw8K280xsQwa
RFVBjGfyS2lxIPtuUPPPBXEv/leGzlodxtYOjHCtL/t2ZYadUH7UDf+/ZeO5jAoWMEehtPdcc2h0
/HBInILtVUk8O9SCyUe4x1JBn+r3LHNr1hipYmm3+/jCBWejc9PXxURzVq3jctY9u2YsHJbYu90U
14r3omGl9wOUsYFrJW0NCaYFEEG3a7N0J65+Rf2vlRwf4empWCJCIR9B7Nzm0ihxXbT3j6rtCUOZ
9K/piyRGnurwv/2FGMfMIvaTRS6lhrIkkmquVpnBH9gAz03qXXpPDvcQuk1yc6lr3ls/aF7gR61g
y+ZWjzRBxKtKeTz6hB8qscGsOH4WtUo9EjfDS5dRZc6BPqH9WLUyJ1tDO9dP3uGKHu8+IyCypnvP
dYpEfYse80cc3LykWwZ5zJio4mLf9K5QZi2N9j2ue1+GpSy+NP34DMLP3LemY+Ss9SgkflwfYjpO
N/JR51ShyN/6KqCTgFOqKWPKhiOSoBRv9mpgsGxRfb4MS8zNnBnRdjyMd0T/8gpoVDcGWQeAS+QW
2nTdEji1iZGGGXS8TxY6oJJBWwbelTbAwcEVbYV0+Auut5/lrbO4wUTMDe8jKlPXL8YoZ2Cdmivs
T+lvkGI86i4VpyRbZNUkymMer4728yJynUM+jXB5GE356kQQGZTsjtqjZ5v0iCGtEqODfyZ6uO52
9ffT3kkay2Ic1/xMUe5kj3dGUJSycPP0RpDEYCYSEKp5S1Nvesnt62Wc0mBfp1Zh0EGuQlyhPGW7
TLwCMI8WrBBafaICPfgQ5874eEHOARsf4UVmdZU+2UaitvUieQwSYf0hT/8C9WHua1+6/vSKemN+
7ngvoptzi1plJToogR+HsFsUCEN7N4o0pW8HTDGby84m80Fdf6NqMfNHWvbpcLSZWKG0sJU+4frd
J5kL4l6o8C3Fpj0ba75jGdNvCFAWDQ3YaWH5sI2TQg8EwSRX4DNxCw8bgchbOTA97GjzdMiWZ4RL
6++QQHZs2vbOMA1Eb+VRzh/hXbiT0vdZYFnyNff2Z2gHuJh+c14hB9PiVEIN43MBkUN/to3E8RG3
14NjVpTVSkYhetGusNAfAwEjl6t74UPbo0yZUaXdCG4aTOqnzKYIEWyEHevKPk9DqCwMqKLsbl5y
USHc/i4od9bR6XxHMM4f7gwNP7wk+n9wAH5yU7L6JHbcvQj5KYOiaUqXWchAKsaJs7g5xpXJDAyD
PHidwefQBRcwPATFwInX4YZUimw91o0ZEUkuTqCg9/fWo3CQnaTd9pYtLohxcXdu1hFI5RPOR1kR
dCDI/hZH67To1LHHnP7LfWvUUWKXXr12FJEUbhwd+6w0wcwXmRHqKIfrlVo96CkxYhZ2qQqFXjOZ
dp+rESpezLDo5+pSiXtZPB5lTl7SosXGxuY3f2OjY1T9DShZIg35ggqirs/hqOrsBPtaZjOo5D+M
45ri4FDC2Evz/awWEvelaTtEXssd5blQQE0VQCrr9EP4cWAETa2o9d3ffR0413wPkLCjbSlrTGMK
XMhJlptzwayQXPhiMfLamwYYjI+CNbQAm1jM3vgRPpJkLfMfC3EQSP/8DEmpIN2KRSzYlWcMIGHa
6ctnBcYNK8lD+WUzNzud+saxqxMuA0N1/iv/r0/4M7BWpnhybC9zvBNAfgN5jtLtyAmexr/hq1V6
iLSrYVVigl3GMXKuwpVsPMiNiSL5LHQt9b4RDB6guk/0CjTEr9/xHFRrFyhNTwQOxU5Xi2a1UthT
crKT9nLQMcXrmAm7NqTuRE6OshJ7Zi6j7mdn74P7RQH+xppDK6Uk5Oo771aM6LwAaV2tAKN3evn2
znmnv3cbKt/zgsDoKa76/fe4kMwaZW2boKNMgk6wx5WHBj0Fu3Mqms73dGHoYtB2ySv2kp5TBFxP
q6zKg7U5UUyP15ekq8ZrYe8jE6Rb54zVRnVLvBKwF9RAYM638SLrJcQi/FHcvMpx+SQcc5n57qOP
yZuIXCOZ+nmERVR0PultrFrQpcKxCFvrLPgJzG/EhFuoSImVTSAeyHSbG5rgsMDPXOSjTUhK6KGp
xylvTlZsE0+9Pk6ntcfLf9AKChM8oc8Z1mVtPlAEkr6aPiIbax/fJ/WTwjMLk4Uwg3tA7T9X8NSu
gYOhTBKv61pyow8FbsmmyumPM1AqER/w1YQ3l4MF7yDQciryl5AccL415Tz5RW7qtD6ByFFVAYWg
4qvDylR41/C7N3t9fGFtGzj4P9YXi7ZFyPW1kdtFRymSedoUcNFwu3nNHDjpcgPBCjAWIFtlDudb
K3R4JaDaLiAAay/oskpeJeRrVeJv16+YltcMR6HaKFFYv8XQKVuaNwSJ1r2jvx8gTdyw4cRmpvx0
Cs5psTzeVndSt8CjuLrdhMENTKQA2iIchXXK4n6hmpgMvYApXMhDvSUpE66epBoKN7vxa2/c+Hj/
uKDL1DeoBlika4zsfXdu4IWoFkfb8kQognYdIxXdbi3NVDdBKBXB7Jyhl6IsALq68IuErLVChTvA
26tZYZSNArypce0C+JSSYeR3c2I+ZBIypboX57vzngNCQ9Psty+KJxHczbjbRVPQZRjMnDxxE1HD
+Y04reGKsnA1qgHyIgMtec95B0T/tZdinWg3iHfEmxP/HxGAl1MkdunIgrWy2Cii6MKnuCYqEMLH
f/w8u7zBFINl1WMx1L4xzN23O/3KDXEoi2IwbPIbx3Fx2fuB2aCwgjTUjcyhdDyyUu1MXy18ZZ/i
iAZIshLOrDjD8uC33MP2OS9uOOoH9Lk0906tVWUah+Kg+jcpG39ufZHzmaYRuOrOGIRFiiDZMuQs
uFigjBQCNe/uiEK2C364mwhqvSFVwTcHIX3cAswqNFPxr9iA3XjA6ygiQ3TpHL6NDIIDXt2Dnvko
C7wbWD5tWPr7ynHEMcv/6mIY/McCuEFMOtRMoGxRMDFC04AP86MfPG8xlBB+8615MiOrzICZMvkP
mphm35W69wwyZx5uLb/4tsyoUpANLQw6gSPCUw0NS4DwruA6o+hRFWix7qIHhShs5mPMciVvgHPZ
1httsAfwDk/4gxorO1azoBvSq3rJZ/15QNGsgIBPKRVSGVO3HopmbYjc2oSXpGhzJaBAakP2ihGR
XyJ6YqUmztivKpHyValnDqltnK218HFr4W23jDLxqQdwWmIdyNCLt/k0TUsoEyY6HP5bPwHFCkPH
I+TRIwUbcoskPcyXAYhhfYKWcMrIrTtGldBMndKN2jA3RgWqFk5h01a3s0VDYZIb+yCjE4e6/xhc
6Dke9NZpdHwHY2cGDbJs5dFn1v0wmyyyaYB6qiTPbVdg9lckGQO9jdRMsr/Vy5p7oIcESP5MvLLE
KnNh3XjTdUX2rPVjbfI61tcRNUCRL6pGIjBZwgjOA7QQoOMRT3AkFTztk1NV9hAUcvo6OoOOsms/
dj4AF8tzumBcxJ7smdmsYMviOkv8FVBt15Z+Uhqoo9JeZdgrdU7ahrJ52XOkAx1rpD+4s/xvY9wT
VD3zBnn+Khs6AYwMyv/cYjLjQCmGb9LM8ABFG2mkDPTyoCcE9hZQZMjdAFjZ4zY6eSVk8DTlOKQz
9FaOJmyu7zgRCguRWfqBRQ5PRk+oHDuf6R4j89zM5qX+pXmEyauw+n6jQgcfCFAHtAxtlHGCA0s2
Cc90U8NsvSEmUpgoD9KoYT8EFhBHwTg8zen1Eo6ekx9VnM82gKVImqt+vUpt8AX3Ec7/R9pXlkdE
MWdBrpLYKr+6R0D/OA4+2dZ0X7lmSVFMkotYboZy7EjUkAc+PnbLlqU8nooy2od+Jz7JYKaLH/SR
Owdi7Capr853/9y7+20xl0vryZ1WBMxAHPc69LtD5eZf7hhGjV6lbsZSrQTYXS/vg8/DVY9C5Nxo
ejD7aopa5fQRcwtNhNen7kMnyw2l5Cp6RJ9KNAgkoKUZi5GzxV1qJV8HpkpGZf/1fT0LWiyido1I
Tq/dOkZntKpj/+4+pUiEu0NN4UcidocQ9BtGhvQyXbrtmMcu+lRsk1k+UhgGwH3SAXQnPuhzDKyt
MkewnD/zV0WFJojGQ9GPODFsMxRbQ0WGdiqhzRoT0QJAnyAPhr5xLMG9+bbQqXQhomBnInzY5OgZ
9mAboZ06PzLjqU9JyxL5JVzqYpUM7lQsSWKQwcWmnkr+TOxxjmx/C+Gs+wWeKc7boeM+Q+pDLtax
rMGoE3+E/RRjT61y2r9zklJZpN/8qKRESYlLwXyd03c7ZP/3ChA5BThcNDLhLBl81HJIMZflwUcZ
HIQlkDI7Gp2I+lwCvRXWIWvvdTeZ1B2JIfOLvIY8i4GJ0hkTC3n7ws67UIc2OYJJ0MFaMPbbabsq
4TfRykTXU8HwB5TT3Z0nfddtzglVHUTZOZVm+UUNmN2uSWgBhfzS1nliHiHUjnfBnxwiBGsDVL/Z
BRc/OrT2ZosUThD1NnNfZ+8TSJ9/wJy1jwfVbuAZvg3l9hKJtgxOTXe+QH0S7CZh8iF5j+/0Y9rX
ON+GxzgYuSI3FY5vk57/z7bwS9DpwAMsYu5lFlfdj5KmxhlsKbuDQLNkaIY0/U9+p2ioCP0u2Fcm
1d+2FfPxvl8a0lqfgo7qq5lGQ8TvyRTDivtpt4+F8MHgRAahGRAjTRw93huB3QpEliCTKyYHor9W
kD/SlhR8S4ABZsDNc0asSXF9Aj77VG0Fd+lEuqG8UTw5/eSqI7IeufhJIOX7me21at2XdLm7NCUY
5lVQO2/z+edG6gIF8Ud8C1X9462vB5PJLsQjYYvQluUc/3pqPtD3HApLSrnBwuLCgNFMOmqLo/0w
Bq8dByZv9ijSEhDPRqBW2+vsk8K6+3cdg1g7jeNBFU68nNV3lI3G146PobhiPFheLgsgHY8YbIVm
eAIg9epP2sT8rxH3UQr0Oy1Wn8ccyPSsQiUPRvBrXb5VuxaWQusOAY2O6ZnYbEOqNawVFIVRj+ih
YFUmBEcnamew4Qu1CIqP1e7n6ysQR2CPaHzEtrd8qtnDl6oTU3/aNu4QyBGhJk9/rSNYOzHGpt2s
vxQ4EKRXoU9EtC93Um6yIPk6FS7aFlUwxMJ4zdX5EzkUEs15yGyxYhlG5b1FpSeR+sYhFIWM2XEh
eS+HMtx/F/h6sC9QlpGp0m7RP7irKsiZeaLczCBEauwXWrefs2m632soB3XKI+/cJWs1AOTRJd/y
qHEvCLuS+iRkIPz4zxzJDSSNZhL4p5GIVk7lWsclZtLQceWTe6iyFTFcGrM8cwov8iPd4coJZ1M+
4xQSgsVKIDa4kikuzk6d+9RugHuwK++FcURjY3WoFV4Q+QxRhLBqt7EmroPmoNBb2j2yOZOuHkzz
9ZtRxHtMjEjDjtGNWCdsKxnrCDY1095zY3Ohr1eGGVAN1cv+1ZUtFjgrYzfQaFbVWYvbVh1Cvtkn
kzLx3UiB0E6/sK9ga3qt8JWFnTEuGaNC0yV1Qzq4RcsJ0oDMKwE6aDjmnF8q+WcckurZdeClFcor
CTIIKqQ6EtovPhG1RJz3a7fIpGje2vFZKlLM+DO9ypKo2HAK+L4hqShF6geBFhYxiQPufoSAPvXb
U7pScjyIdQPm01ft28Vsg9+Le1e3iyzr8UCSyFHhKf16A4i+mtapFIF3eXUaDDOTjtv1yS1U3JfT
31rA7cx79kaUbKVutQJLFW02zRkBIeJoqhZtQBiTW7tF/JoIqC/geLq1l6HjHiW9Er//VCOeiWZ1
TJ2ft3uL+gEmK9voFBRU6TBr4y7zSJ1V65KCByeAjFyKHpn9rSomkrW6hi/EEoX14GBKWVtRzJ0S
/wlA1DP0JzVG68URMukR+YLu2TCXL7Q3UQraaSZWhamfPM/QfiF8cGWBhK/kVoW/31DDmqPMMaLD
OFsd58GQDBOqI7r9D7bTrPjuMPwWc0Mnv0yi3s2FlnvBUaCr+kbJibv25RAVkFDV7Ytp5IpoYxRO
J06nrppnxgu3+/CKs7R/I1hfa3n19HHP8U965nkfDop1Agx9PWDhhWQnSoMpVQjMSAjcI2iiapzG
JNtF6voLlEbhoB1CtxP6L6sCV3zC0OVi0eNhmGDVGWJ5LCPVonY6+F9xFZTvhg04rHs8PzbRxiSp
ONtZ5HCG0SJ0DYHIpY/m3IgzMewVJmBaYxbs3xbFnxCxMsgC0olOvXG4cbAh24NDUFWgzaxQLpbq
LN6T6AAKCIu1BeOv34wwT6iIw5obFDSPjF2HXeQYrtj7pm48/PPgUTxoQ0OpAkPXZ0bqsykQJg2N
eiyrxBGhLL5E07GAraf+c1fENBLrhOHJEnAkZXyRM3k4tj6BfaXF2s0DNhYHT/ERhXBe7jd7Jhhl
wUXAYKs9dSyJUuZhUZNMmttSd77167DLBJz6KBgNshcLODxsCnvfR8mYw8hwOCDzv8jCt640Wwb0
8nnEducta3eKdbhXwsL+Fq9zQV+av62DG5nA+y6d71hDQnHRPehRXPFFEK6HI4kggO60sdYc5frw
Y3VBv3qofekXBfXP3rWjiVHDTqsF4a9wxwQ13qKweYNbIeQPSxfwX6stJqeomzEO2pRo+EB6IrOI
7G0/C19y2GdjRv8vzdKzPLeT408P4jrWQY5AbBGW2UXSt1HMgK2twglVR9FW6Mm24/uirCWtuMOK
bPzPWl3Gnsks+bGC2VO2DSGHlHUO3BDsW/DE2LBLq3Nffeu/WGfzLOz5YtbUtt7djuyS1kn5Q6L9
LMwNI/VTUBRnI4ZYFSJQhzvk4Hy3hjDL7j7rcLK7M0im60n0tjUIhbvqjvdXep28ekNQEuyFrV5O
NdQeSO80gITdDb0qPA6KukA0WmpEJIM8MfDj9Ze6gLUaTPrbWQA8+90gxT+5uAYnqhOeU705Qd2r
ADNV0lGFg8g1MWwzT93S52ScEjS6/R9wwDgvoiGicQJ5K1VQb/4I7hcNXjEKUbuoODx4ObxdEJPV
FNCO2gwkV4p5LSG1k/Y9YSwCsMXVip8tYmm33CSHN0HIy7DkPz42veNACaU/mI5Fpye0N+OoBtrr
s1ShOLpobGRYQc92B8lneLdsERog+832bqHxlN0QK/ubNQQsYNYAqbyWiE4u1JFrVbctnrq5ggtW
dDtK7ML1eJequ+Bn8mmEyIoBkb5Cm59UaGFtgfVJa/df+fBUoBMJsiTNW1HwMXNuNCOr71mSR8je
4VDYyfKaZOeffdkY4TpEvdtYwv+SappYPtMkQKUo9fBDwfxdh+r1tiYh54HfT5aznt4ZBt3RcLLj
0Lf/yfSPrh+vqX7bGGfXlHtR5CwDhpPYyxyIptJw5+3gQWxmu/94iHT2MosJJei9bNkm1sVaX5K3
0yr4gw8wnfPJsFe5GEJ6lS53SvdB2LzWTIqdO4QbcOKWLA86eAwK7iMnYcJ+s/VRaxLmVCHy1IXq
smLDzqZ2qdAYgRIdnEidlGkydDSyqoVX2MPKOIjOQuJaiLNGpcHNHMJ7Vj2dsKU3bSLJmyH8TTB6
m5O4jM23cLnyc8pGqcnhaMFk70qBQ2zZeYsLCy4kGAbnES6hlaZGRpGfH64NLlqB088xlShazR8K
MOVILc0YVvmED9ycI/QYzjIl38uuj7r81rPXrqA3FTHvkbBcGd/0qt4SsmB5GFf0Tjp5Sm6KVE/+
HELegpbzM1hFjQ/U+On6SwAvBEz6x1sohToxbbvtlRQcbNsNv2xGAXBoAw6ofI6BvlzVUIq9eljG
1Anie06MSIA+52mw3Ye8mDM/1fdfPM/qQDh+fNofukuCIUF60dOdzWUmy+9Ngn3lqpOOxCbXkr6Z
vPaaLArkSYx98hWvHBqMCIa74rd3C3uPpr09B6Ms5stn1NzWNPiJp3uVJMK3pLkO0oJm36JBRU2J
F4gWVRbzNXA0nKChrRzGq+YXw7u6cdTuOe+U8E8uZMrseILfELQq/mxfq3IBYWsr7vRJ7ORBP7CI
hRniEZLq/8lLPg6J5n8ZZ/3mOLj9+2SeSLqtP9Y6ugaX089lIfmHdURSbTHHTlYWfzPz69eWRVbE
pd7z7XAV/7Qn7xPnGguH0BFSLWRLPm9Xl3RoVeIP4I7xlh4zFDy7o0jkT/TSSy7zyIYM37i6UgHL
qG4yQHRwF4hfmQqr+NoZP4VCwqtQUyCmZnp45C1g4Ls7tKCKQV/GrX8yJqEAs27VmRGg7257LAoS
AfXn4FXRRKdkTaVUonWT3dMwNOg+Hak+Smq9scEyWlsgg8kPaOcURNhI/+c2zCa8ZusXTPrfF5Yc
4rje4kSoClkcI3i1PDjXSCYn3IC7U64pUCuZuhYxyCBDR1gV+k4R8BW5J5P0s+ylqN0dDSyISA4W
9amj1TJCUy2BepvyvHueDuyMJIWmQd3Wo9mBMhNKLT+9x49Gxs9MQSzo9990Fh9Mgaz4tpjytHeB
aZelcs8u33TWojwLHu/s4CIFmCks5ethxjW6s24TzRzFdcwPWPPA8vS9I1n4L/CljxzQYmamt/S/
0C7DoXNCNelJslEioirK5Q/z6QBX/Zn+AoOp/vEQ9GFw4Yj1w8Xe7ve1mjYsnwZ3ycBGlYam7tgK
G3tQqtVgZKOqZATaDS3sNnAdzpezMHU58/l2dzdrPU0C5ngqCQaC0fYUr9HkGhaHcDw/Z2KOahYx
OM3qG2caX+Y335jNsmcHoP/928gYvzSmKM/ElgsVdbh3vEq9tgZMO4OfGQiHc1vjP7z1LS8Cz7td
t5VZLjtGJVzwn1yY6itSLZfKZIUFpSUGcpVBC3sh7Codtry79n6UVB/JzjCvnxR3mKwEMTC8d5vf
PhQgZ964fMy4M+rsEXS3nJ31ydgI6Gq525zzREsUqlpOGd5eXCONplk/R6WmwMcuZGHbQ6H9eSJe
UDTjrV7Y4yy1v9JOVqWasvzFBEb7l86VJFjPmPTnI84Zfr/NLKMoIDiPw2450iUW98BlZoyhX/gU
40puzkJ49l7LqcGxf4GkNWggoj2/cPkhux3Qw9xjrIF8PnBJ8G53cvLKcKHKIpnMCtBVSICmO6rw
u41gdLvKLHKM3D2A8srhf4+FRHWszjJb3Hs1xdKZCTz2bWoDM2h4+OEyTa9AyRH3s8o7Hxr/KMuD
qqKz4duhd/8pCeipxe9o220wMq5fY/olZTS3mxQTXuZE37vSfIbGexsxS2OgFLR21eNpZdmbdVlx
E+SCQcwsBXEu00xg04MlKONnxkJZJNdSjXYrNw8nPVlU2u1tIkYMcev/CDtsqn7TiYwFd86+21VU
qn/L4EVpMhD35eHBssHVtqHeTr6rPx0BIcfMtfdy/jEZcSK0B7GvRztnUbcXIwUfgYiPpASzDhye
pJaZpMe5vo5ylMLS8vfy2vJyRMbHzIZRupI7PLxRO7tCnuA8Eaj7dKGGGTYBBZmF7sQILhCRotD5
CwWFrz8VNBn/y3E7j9j1WtQq+v3YEzO9M/8elbRJ5VWEBuXOmTpsMZPeNeZwgTso0kdBOLKi4Aaf
FGThZWxfyqOCcmi1SKV0+/DALe0ZgjmFYxr6bf3TUTM5jDkTIRDIN/QjhBog8/HKaDLznrHFZSkp
XV16Aqqtw+Nmg8qHeY0ORaJf/g7u6J8FyvMx3CJfcABV1MS+Z+XFyhsDgwYJqW6LZ2tJOhGamyHe
XjUeB4KPBZj2nC5x2T6bwR5Ehpk3SS4SswROpokPgaZxy58H5xn4I/BQOUOZMWwp4keI/TfP2Psc
5neenFXkCKHbL3iYv6smK5P2io/n5rM7P5jea4Lf3Atnfac83Asu0tl+Mfqfw6pBmoQO+3uQSknL
hvPxLg7taxFkpvsHQJvYA1Cs+G2C+9Nv+kXwidse7oJN12KHo2af1fLhn2bNpEvdBAhmzoiZeI7q
iovQnlplwZ3w3aDtxk6/08Z6poAbBfybMkY0l/mC/HkRW2c4zKbko8bZHnWbcOyP8EE35lVmzcMM
HdKWnxY3wm7XYClp9KSQ2HY7iCMCvt/zqGIQcsjpRaIAXHWQjcBoDLbwhk/iOkk1/rqD50AXJcYo
kvBNVRS/tcPn0L/UfVwzng3TooLiIhSrcDXnjnaLYfWtxbBZ8+1ndRttM2ndGKooBPYLyUQfYfFU
5TpYespX0etkycUUqswfpG1vxWLehU/AjlX5K+DZDWPF6m2hzV/CScymggY2ffcBbY5zxm0iTuSl
Eyv6Q/JMzcxIOdi83mMb7T9ZI7oF8gpNr25DCXTmbx0Ej0lYT27t1rwDPFoURuOLJdkaFk6VhgDT
J8rdf6KUagfvDGoASzoeT4gmd06ZlIDWt+Z4/OQMOUr/4eEpvAn1mSfhQX8wsldR3w8ZRzBdQkGL
bG+HT+1uT6zNfobD8j77Pu/LZl9nLnZBneblcLDDOuKPP77NTyrlnqbnNoswF5Nh4BT00J95eg1v
ZW/Px9f0o+nhjVhKPChhY1JB2WpVeTLur8hielb8qJ0GSzV1dnFkMDPW8Vnrg/+kSZrUAN1v90db
P9eH12u7dt4wbKatHMHp/t2UW79sls6vrknpLUCkcUQoeH3TH4h0dS60mftwv94R9UzhaRROfW0E
IEj2Av9nFpWpXV0mjvUbTzTFkb7qh5Q2S/qq+OVJWeYSR4uhYG68z0IRYvVlY52HnMjZVCJeLXxe
64zZHjrEExy4fqH8Z8TtS81l2dUX7zCip8A+gK1Qtny6FUM2pZzXNn4bvw5ykMLd3kIybtnvIOfz
Zsa+uWEiQXTGwEPwWZcTsFLIc7ODNGYWb/OZhV2VsREB4D4CqzuN7FpFomLOrLvHJUBePlNwEdWG
h09EDymJwunjN6L1+QNedglhtRW2VrginZGk9XnkH/TAGWNMWt5hf2rX6LUSzMjg2TkdOuw/KAhL
dF7lGK3ySDgweutvhfpcDJup6DpvKvhMWZ56GmneXSl2cZ7hJTd43Zs+7u8+uf07N9xsrXr/dSQ3
aIrNnmiyfNVbqhaf+pBGiDTg3VLwsysiq9SvR+1f7RlsgKUrbjG6c2fB1SvT2EK0CyKEDkOTDFJs
dKZfZ1jNRyxL+Hy63kX511dlAV1/24ses6rlEhPeGZLRscVOYky/b7aZ5VeW6+hB2Li1lRGHamGw
0S60uPa5T+54VHWtburRzfL+5mRAWsmpZQO/TIThY76Quj2faBcGi+imfYmLdW1kMLQI7DyZ/yt7
HQ6Zfd0dX2Qa/BEvlpk41SaoTFPAQw+o1dHprr60ZF9dlTQIrWPAU3MektHt0JvR/cNtJPof6/e8
yvWQ+7zuRKYXXje39RYYKwXpsTN4saZHwE3rFMeNxfQeMV8ESuYBFrysFk0bVwf+sJ3dQOLXA5eX
tfxZH9VTFlkgbk5GZkGAt0RNli2VIkJZcWB8ZL6JbZJLtke2PFCVGmp7k5hL99wT8j6kMehedpoM
Fv99CGMPf+VmCoG+4NofelYA8wGvxfBDj4hh30f5ase3m7xW9OJUcGWn64pBF9/d5nmTzfhhLDTA
472OOZEm6JvC9S0rtqtemd7TrKtTzH8z0RVXPUm76DvdcJ5y3MvomX4l0QmpovuwG6MHIaZ6t/Cw
Y4XZcFseNA1M6H2Eypsmf8Rr463gAmn0Vy2ioyo4lmQy+iJz4cqhboE+jNStJtDEkIEq6lqlGLmV
LB9kaWaOlbnXsXEBdc4m8RK1OVfVipDkII/M+FXn2QXrkt2w44Ld50DymklbbLn/2EwxgThquxjh
G6No23VQn/o+wO+fpHP9Lk9DYeikti25u5D97W1ixcrFvU/r61YS73pihj2lTxJYf8rkJ7qZ8xu5
VLTw2hZzUbrc21E67RzmYO2EcvOlrtChfKdfH97aDEYsGBh8itVr9FGwjwA6BaI3gXIzgiJI2vnH
QBrFraaDFVVjFMqrAxSg6aW+XDeH4oVqwiiLOaaS9KJm53nXzepUsYsPENvZQBGmqkGEVW7HrkPw
Z86H9oyfKmqGpW25S+OlcwBY0YUGEKXyHQXRsn6ITA8Ca6p3C+C1c1EQ75DVz7EFAJaws1RGc8E6
QUf8bfALfM6wsbg/L5QinmZOUGWZ0v1ZuKz4s+xHSkvMwpxlFUH+AGpqMARxxeoTjZPkZBDpnPER
2UfKoyDOwA7ZNfR08Cc1YjGDV23I0vk516QFTBiGnJQ/t5kU3d4uWIMWmPMslBFVQNgKizcL3eCA
zKaHXMb1HAvUcG/cdeHgGeMfp9uhuIlbFoxUaM9UYH0v3Ju+wTmqPW1GxFxi21l72T1fXqHDtZah
dLFLyST1l2k2kdj++sbFY+fg3KRWjCy4S8HBwXW2pwSV1m6kGTYy+5+M0H19sgtCffBL1TTiJ5P5
7pDfTICxZlYyClZ+ZAu4stRdmKbfACVrFkH5AT4gCrt4XZnJlgirya+OHRkQKvZcs4IxCMGkCmWy
/iFtt483+rM7kn0g22QB1c6aZoP17YzzfJurp5Kbg8rkHlRgUN5caAQRokKwttxZ6QqwY1nQOczi
Sg1SeaPrMkVshuke4KPidPP7o88VCC16EW1n1Sx+Z4liWlw3dGYg+lZYoM747gNZ06NPHeZ+B0A4
2ykJIJ3Ni7xIPUsf5ZwlT47umjBOj5pX+aag9D9gPH2sNZGpY46wgH8SaOFtPNOJGHjicgxKphvw
xnmiOKEuXRU+90LSlV93AIrOZFKsURFxLy8384JbrwbmFMhz5ZCpAGvCsOjFBNG4xMbsn2hmjzt+
Es9VfPoftWGoh+iJbF7L5EaPhrCiGoxax2sqCajbKaN1cjrpff5Ne7K2zkS10vj0RrLkTfEybwVC
Q8vNapUflSRMk1lrp3iYvYtT6lbZV8lNl2rFt2Dhxe6EuSZ+lE+F0abtLzp5+h0iUEe+EAJHYN00
YSm39/Y6gVh0Xs3U3W0dV7rMYnHctEyIE22VAKIrtVoXlABHgGOtEdnrv2E2//B/Etg3g1LVjcD/
nx5gBYF4qLwqSF5nTIJ62jYTwYC2wmlkbQ5thBpBw15U0XjFFY26Q3cPRdIzF+vz/LoWMLNnmx5T
5Iry6kdKx9UHOnF3xD23zjSofqSsLAGt2JPESXLYge6uocm6Vx59tZBDU1sptw4B9vChFori6VE8
F9qLZ/78zNyVtpZLWCffh/b0GqhFB86yIOUMk7l2s5MM79sZXm3jlFLnLXQNddlBDTAxkCKwmAwe
Dqm71l4Wa2FlC6wab1yTB8AcDYCsFwhW6v5XEiMDj+tkv3pFeMLoKnSjsxXsySpsP0Oek5U2aW78
pbHvGWuIveCSw3/H81HbUzHqulh2MLB89iUdp/qgdpAkqzONKcBbd1P3Tasd8PXeMLdhNchwlYBB
0piZNjCtNQqDZ5qCUF5uxpxEKALbToaQNmJFM4NDZDOH4HQU7kP9C3Cet/YJc8Ad2KPZalXgOstJ
UT7obYEcay+9dUkZesqqB6bibZ1MkRAFG6JAOAwxxiAxPKsi3uvqWKVwNdgeCh150SX46nXEwQc3
AZIq1+aI1EPmWg4bKJ9sEl9TXtfuwZsGoHtNHY1eJ67/t1Yvev9VDz+RYbgRF2oJswEh3Y1EoKj3
1HNH42HVJ8yaFJaNLE1d/xUIgONIpKEvs/dVg037PCgzhKmLdDnwec+tFbFNNPo7QNyrcit9nlOk
4ZFafEAvijwGVmwwo7C4ng6IR9O5lfF82iaH1bAxkfFGgt54AUymSaIzuke387Zozev0oClnlEIy
uZGmfMzQ6AVVRXb9Rdms1BJVVJuOAfStntLLi01Wl3JjwOPvfK6rpLOTW4hfpzL74BHCaoi7K2o4
82uyNa3kF37SkGUa1mb5jt3t6shFaMX7qsrTI+Ul6sqd9mlnNnU8k2t5hXca97ghlBg88p52tmlD
43jOMU1fVwc0mWmfZbsdwfs2YGRcCBMZKm7Tz7aBGa6GTw+yah33Af09EquMO+ssev01Bt3sqhDW
0WHjkSLBo4JZBdBOpO8Xs4m6OSUYbJM1AJqglNpTBo9uh4YYAQi5U6OG0VvAjmgR0Ogva1B4bbG/
M1QvEXBahOGX5ylTs0oaamAwE0TFmWICzX/ibM14T3F+1iIkbsfDyGSIbofzNiStDA8QCSQ7HHGu
FbGKM1LtaOnKqwyTTRzP+sVb9DTGokOki15tcSvQqED+a+juFacivzJ3NIPQZwuP8zooUPLSgr9F
wx5CA+mWgl4LsEG2Icg07zFVAB75H5Nlh01b2fFL2D/WUIzJh6ludML62thKWl+1D/js7UVLoj19
Xi/GZt7EJtHfxAPsCEb8OpDhuTuZoFz9eS2MoBkcZH0Q0uxdM5Zw7Ny8SIMSscFpy5ECnvKg6jjh
Tyg9So0CgjhQJi+qoU6XDfY1pRbkmynVF1978+029mAmyabcRicUaOfnfQl8/ELcKYqhsQQkzII2
1Gm6WQRgVNf4oXL5Xw7hNSPulvsfMMaAM0I8hr63v7cFKPoJ8QmNeNywMqLeqsXLjGn64qm1gay3
GVR2hX7m8teVYQy4+8KvW//GfRrQ0p+G/4cnGmKw5+7MOQtSIxXXQUifxHB5pInF0GpE8kYAwNF4
ue4ZCQpQoDjfBOVt9e1vNFF0WxfwpmYIKa8ZmlmHKaF6f1jsrkpzQVUJ8X71GKHau0I7thxZ+6fx
9xNLVi5nX570jpbewj6gA1bUlf8ix0QSBNqYnhjwFZpewWKhVwDr/HH3IZLUNN/3sbdDqZoRvvFI
rg2YXv8efBOFKZfqeKs7kEFjIfD8tlNh2tMhopP4EsbVQIFk40ZNja6Efld752ucbg1khkvqxE+S
LuZtjxeq1WtEt2nUxJpyFA3KeMHfbSS/RsNETFRivqc5O352shUowDE31Go1DHj73YBa5W8ZwWhb
kXRXEqfS0Of0EZf7Ues8Z6NqqqUUUjmTSiOahZEOKVMTipnrerFXSOg58y6boaZXzD/OfPpyHwgq
5wL6vdq0RLstqF4LxvxvBUF8OmKxzWWJivqq7C8MzYfCmFpjFetvMQ9I0Vh6OgWpgOEYvX53q+Kf
Ppe2Mw3nNwHvBjoBnTzylNJvTha49T2PjJKFBRxIg+OwKKkXG9BtPycRrzN/H8dUR5Vv1e1cKmgE
b8cb9/lO2wo2DpT9h3qRtc6ddVrUBWzi2CB9fmXYUhjLK4dHuF+Sq9R26l0q1DxbgEs9espav+mZ
ZLvnhsz21oHJRY0iDqFlRDA8D579LPsCcztsnzOtUoIXWbU1kud6ZbWNq2OcOKaEWL0zHFQ4f4nG
KqucUg0zxCJYoelcxtDm1+/cbhEUIdIEYzoLIeWF4wuMfbbaqwSjUW97fSh+N1RJyjjysyjx3tYK
S4gKrhjz8nL9iFJRiphcUwZ9v6wSetZF/M3qSr8lJIFMQkC0il7xN2DIZC76PvXEBwzQX/9aZ8U1
DthKPJ54OdDls1vGMixXqP1JFF8miBjgtO+Jun4MnLonltP3iDZjwZh6ehi8SeacfjgEfHCwEcLG
QX1kfgYIGjQHxlUsZoKgduxsmW+0ysRF/v8HjLyTgGWQvpTncGvtkOSsJ9ZWsjhYzabnbGdi7eAp
VU8hLZ//i2cysDWtRdoMyHv3TnlYudFAbc5ZR7xMhkzdhFOeUE6rsy2XPxJaPQjsPFnQ4ILhmxBH
fKUy2ZL5ICEJJ66F0EN4kbcSWQDUtGP3dNdKb05TV6wXL9wO7ON6SqHWzkNkw62A4PI1tfRL1uj6
vRSk7puWxdSzMUdt22R+/cq1NFTrFF6B2PbzNLJwer/rLg7pCt1IcVx8UugvskE1x+8bW5CrA90i
vOwqM7PKyy4bLBTXv9ABeHXCZMYROpHIgaYx6inHt1z/WlRx52hGhZd+cwoY2t72sCr86CP+9wl2
T0dQFOZLHgZ6Sf7HZXGGuAU+yJwi8+Z2BW8gAqJffH20+nrcbNSBv+vYJVPnMjiEGGLtyT1fke+8
jXFLELbLeJSNPQL2thYLF9WJshVZGB2L6PH23IuKJfdD6BfftUgZ6Y42STcaniflGnZZA1HGQohQ
PoF8OPdQZ7nk1utOlcDNKkkw7y1qgjeyFWdjwcg7z4b9fq7GarnRqhTWGDsh0EaOE0h3NEsFOmth
tfRjAGwTsgT8n2/boCuPnUbyaGreIoxyOIoU8oedO6KqqC9av+dHRkXRPW7v6496vWthesrGcskZ
T9cT/dJFtgrQG1eBSqLXAxDhnrhFjrIZK7wpXp4nGdA7A3XZPzUTmOTNLyYzTEzq6xVPL+XfyTcl
BGDvevenvYIioM7W1t7E66bqWnx+IL62XdEbsKoSZEfNLvhCqfohhtLfcNvpz71M7N3qvzlCg8KC
/PMYGyzK40VvGuZez4scr44OYHydmc1srqXUK3M78Yahpvi1FuBPOL/T2dHt5dvnhaBI5SUUJwqh
ksVZ2B83yBG4SXJU0/c18b2Fbt7ppqpaNDiC7U5yC5Xc1J6Vb9fkiJN5ihlu9MJpO3eWXJT98RH/
wNbSAa7cY7gPlFaRGmYP70xzFxV5TLLPY+f++TilWPDeCzDXXbI+lvuCX8WEV4aM3SNCpgBzTux9
YfxcBanBhzB5FcVE5vMN8H8B/rhKXOqsUds5l+7ItINpcGrgtDYSKuBcM3uc7ud2LZ7jyX8+PAmp
moQkMF0FCxDqK4SsGsTXHWLtfSbho+m+ObpWwfuv60cFK17hLES7q3Qt+TR20Y4bGQRyjvJfyXFE
QWbb6l/1NIhd+D1W8fLGYQ7bJqalONBv3kavFnp47hiyoKNDRHkZe+rA6EDZuuyJVTOmMMsoZlTg
ZGWSmPFpUeOVoOQYU5mxVpt5v5Tx4y06PXsKfQcn98UMfQZaYqhnheQlGF7Zcn79+8HWn1LknpGc
GoaLBYBne6RljVI3vKHc3f7tdtWXSDBN6FySdfm6SiKFrHK/QntnEh6SdVh149Hsc6KXslxt+Mc7
OJOiAm6FQYZpLJNmjrh6h5K2qLFTmGUWB5AdprAzJ+JTVkwcxnm3fmCgM3/L+nXWgH4jZAfZ7voM
QMeWt/77yeXRl149ywAgwhtbsrnZyc+EyK+W+NKKAB4Npa5Fkls5tIAzgrUA7pS6j/KySad5M+5z
ta07PF7hCbpSOI82bafJ6+Rh52y0KXkchhqTFZe195xQHar+DmyS1czbrplHXq7WR1Kr5EuBn6zM
JHufeUUfSwhF18tWunokPKFbFOxPwXd6LNMMB+ZZioBkQnyExgkNMuOgsDBMNzhyFyF0P7bG6hmL
wtw+HMrn9zY25dA9TZNTqfMnWabOXCoRt08ctzInEruq1J0jzeHy2PZaF516a59y0KQmMSWR94tY
N5M57Kr9rUXDcbmBkmE1KIzKZTrqPs+O/baUZPvIJ1HmH0TxBgUq7SfP5fPqvk+GfMligAmhnO/M
Saf/31PdmhmhdyK1QqaihAt30Xe7yt9DWluLFQlGl98CwiudIQBiqyAz4L/pJLwuYdYV9ayLntBm
ybxxT3BpNBwy6a9+C8zRX15GX7jzNfJJ2CgHGtWaDRoJfckUFyNc+HGdGLeo/exGDL9Y0rL2qqUs
Nfui49zGa6F0mkQYCKbMPuL3HChkMpn4nBpAMTfhvWHVBIPBqaq84wBrJV+Umtdiwuc4OnnbmrVK
4ilIdqNxG/3JXfXV/hU1xzNBtdonL9fkfIKi7bEwZVaBup5txQBWHlYf1V+gWOzH8EHbZdoofE68
qBi741t8MRJIy/E0CbQI/e89N5/Qwj/6fA5X57V/4eDn+P8oeHT6TCyJCAeCMX5VgcWkRUTVVH3E
Q5Upz4XPCaFz6dFavyo6CJHTGClW32wR5dIoWBAY6JS4kf04ySu9ac2QvDt0u4J9fCwT2eg3kZrG
7UuHw4ziWSW6/XZ8Q0c/rJqAidZGlvoykPEbpPIopQxFlfjvk9sXA5mcJIrf8MZJaHPxppBav2p8
7QMJbTD/36Brk84n+iGImLYq8IFj8Qny6AePPTyV28Cotj5C4SDH9QeUiiO8MlgFtL84p1MWVHby
moKYw5mPKbyClAhYpv3euq+qjAPKxmq8oL9y0rGnIy9+7wyn4rccuX3cofH+uVHkUSIRliF7G7sR
M278yA54xOg41VMBDQlK8R7TODfkjy/xfemel4MsItcgGFj/Y9y0xFHEbWsfH3gZc7Pl+miJ1L22
9hcSBkgPEkeeBkd27nfcvoR/Aqual19yTFd0tau4/KP7t40zPMGLl48yY5UqVtg1UC6B3+umwoHe
AcPVwgTKgC+xih9LeRdktN9Bty5SdKPW9rB4BcVK1jrNXo9pFFBHt9ng0ZOxJxwXik9hhwVkK+Ta
n/vY29Zz+5LCyhQvi17lWvWFIyTsiAb97wGQ94M6Q3e7NtGoqMQx38FwHALMvVqYSBDnN49Znqm7
TeLaw9/LUcoKlhQGr8PDrYGXzRGoFEmkedsCPLNE1HXW2rKo6Tf4WtxbjWVXF4RZ9CuGzwG+K5T8
m618Y1ez/USLzQldzl/wA6rLjzfhS8brgQMktEXMYC+aCkXpUsWc3ShVVyRwnMEcCSXFdayO1msC
tLGMnkmR5phP4WFP6w3xEch07sDzUHnc1WvHgDXmibd/oH52HG+eb/47z2PLsYVmHvH/071bTrrs
uM6ruLCDnYPOhVtkNS7PUB3TuFAIndQUx0PRdS8pb+zzvFLriH9tiMfK8nXsDTo68fJePHoSsJKE
V3Me7YR1c877+QR6SKOjfPa2OR3q+ltpWLxuemyPpmMY9vRWYoBV1Cgku/wXFHlswTb+bDsjHRyn
MYHwjf/q6VXQK/+Mo+50jJ6AnK1PhaZJFh9H5GBK72e6opKkT6wAvX8QD3ER2N/JJUc19uP4mlzL
TyByKMt14QUm7AwW+Pc0pMJxk+7JD8sr3UMDVm00Qmhq8WwxAHF5eynRVqhy3IIy+mk8GY/hmJXv
9bH9JFCfhQEuSZxq/dMamYcY+BeeS3Olq2YfxGAD60PCD5oA6MtUGa++eQgB09qgpwSWVR6R0lZm
pWfIrzEOqo+o5IRxxfa0NjaXCqbbPxAbon53kOEx50vp5qpPnSlE2J26/EpjBmtBsh8vK6a1+hbJ
lqQgrxvFFr5TizhgCYDWJTOb67q1n6PDZec/NkHNxtWunZlLuBXQuwy5EJQFBHqLjp8QF6JVPyMY
ltaM5JmgSCVZ8wibtYG2TNK0lJPJojk2wsSlxRM7Q1bHKkp+aXUakXdUNo9YTeLapIM5tOIMhXwP
cLfaepOn2sTzVRoL9HIWOdMRZr3fr8RnDG+T3LnSwFTboivH6uBfBWtIenhM5C8Mj0Iud++IfiUI
yENzXVucQIev4ZBabcFqha9MVY4gFVI3V5JPL0VtB7ND2sWGMuOWTcEvYev0x6pnS86Q8w+CdSwt
Tr/Tm4rabuWubDdv68MOvLPCD2ApcrDzcdHTAeI4gElLsC0XyfqGtL3H/Z0PQzFn90DEr1PWt+50
1cVCzjs66e+jYVauIAKcGvI/ud7cPxBaanfrRkY/CYjlZkyCfsKNls8wmEvPEVW+l5DnQDlEda8r
xA6Plfa6uvkuF1OmgVLpvjs5AOL2x0koFWTSj+2O+vjcDoPfujiwxhK4iXR1Mxlj5fRWmU7nqG+f
5mFlIecG2AvCRNXFKUeHJz1xtDC2rI4PUtbhbJvrfb2Xsf5HUE7Iv/TUvI8xG0i098thzhQ81b6O
1ereK6kCUNflXX+soDSWLlCx1go1nQkD7+7DaHaLwHj7LkqvmDm2a0JLA8WoaB7iUIuec/w5lTdV
Vs/Ki6nvNqPxY1YoHxage3byToIr5g5AU6oeN6dY+1hJpwYkTpJ2oUgu1oGuKga+zqA4VYmlxBp/
NjgRANl5A36ZZZjO1S+/j6swuXz+sRL+KYuc31o40U6EHo/IkzIWjhKZ9Y3fhpFtceYGHBsLAEqn
edRmkcb5Xq28N7dZGH+3wT0AkYm8UTVmggHt+NO9HKdTv5IM3xoTPKdlSNUz4bZhROcdYfC0s8Rs
owQGLy/LKJNNvhDDqYBqupaJJ8/hxvkn8xoezfEPwLpAzf0Z8w/twcoI3bYdITzffDaui7MAT3zb
n3LBsFYoUNMeEgrP/MOOW1njsTjMsoGUyh6MOjXs6YPhGDsemaOYxYLPEUJgTQaf2Nzt1mfx5I9y
HJ0ZO1V6LLlao+TVz5hynlDZQ446zXtN+oR50M3yQ8V/zsmLA3qzGMeiHZurjHNq019selYlfdVd
mBZO5YKyzJb4HV973ThI+jy127BFkkF3EMpKJxB9wBdvEuFS071X0Vq3rE0CZ6N1Utqh7a5SYMqw
KP19w7Cn9b53oxwVLF+E2DJkLmqQCQOIYpINfmQApuJZYg7sSVtYAyj4SAn7tVVbn4HupgazMRCx
WBUCWkw9g8aLMJ6dDHbmcfY5QS4lq90tvwDabpivUhT5H7Czcl2q3OCFlRH4oHZq8W2TISoCLpx3
PdhmUnGnXzHO0eKYkytbbtmb0WIuqp6pWeGn2gq4Q3pAiNhbM/7mcxtzWtQRtw6h6jAXSUmulU0V
4g1nPJEmmXnRim1lnWG/iBEm8CM86wYjOLNMg91s1+Ti8U0U28eIgNJlN+4Lo1hTaEMRj1SDzQTa
nops5INO1nKr++Ue/+/AmkcSAGcVyPAoRBtGxZmcaJQzkjiYytpXDY7wJ4W1GmLxmTff4juqIADy
nnoFdVIHJtgCEoTSYAHeKv6TynGhTs5qyGRtBX/K7Z5pykmkVO/cIJ2di52ybBQJxdqOSvPLEZra
avIjVQb3u9VwUyQ+Np85pGPMtawAfOSQTS0Myzb7KgQB5FFgwUbTEAwxNP9c1d0WDBqG/Am9rI+O
v2X6lhpPqX4etyPV5oc/ldByuFT9eSNuokBh1tjKpUqy+HrYeSr44btegbQ3mlE8dPV2/PWmh2TJ
FOR/gP8PR28ZomRs/LFk8/mVpoKN03zsEqa7LHkVzoojbppLAHTctabPlvVl1ASFIjmMopayPHy3
n9qq8OThqgy32kV9MN6CgPtJ5jEyWP0Y5MDVnk+ZtxCo2pCcnTD5PAquJTLogO1O/WvYlvanwW+f
mORRsupZ28X2LtyGsjPC/uKP2ZtnIIHb7hMBq2JRAZfsywPVvIaPapwEf54bsbkEj+Mz/YgJbiWU
Mk1vgHq98J50ZyEA3mw5/D/2zKFWh2Cp1CX27iap7EqZf8kLBaCqwl2rFJDjtsEPZNfgFlFl9qXx
NWzMHx44HbYhs3X48jEBl6wjEfoKoHIa3Cq7K7mh95X7gYk94GV8G4k0PKHbjTFlSzpCgml1e3Wv
lsdDqtBbsA+Cra7Z7YlEk72rpWwzD/9/44PJjGOQuPVM4FsOWQraYOm52c+YwQuKQvr0FskCqmRX
AybI2hXoV4Ruv+Dr9PpgGG04m+OhxfyvK6m9sSkt1CA31Qx2pyegcRwFpTrmu5xPywEqka41zv+Q
nCFv+j61lvgSNdzH4fTSTIZZrGf+1ff436HBY5z7QJHbkMju2LbzLSyr8d6pHGVBXvRDd6rNvcDm
s/NIxHvBQeTYKfHlrtMM0Eh5YoSrFmQGKd/X2ImckJ9svr3vA65jftlvC9kR24gx57r/ZbO9nxAq
Gd2HaQ9NiXzp5+FByidIvj9pPH3ha1Glw6GiXf+uoc3mdJfj2vAaryI5oh6rC0e53wQSzg0PmxcM
ykY3wsTNBRYKyeVBujPRvXJoawDKDAP2TflcAKIKIlHIp0yb+jPvaEFniQpmbtsEOem6gm/GpFVG
ChIgg87xBrUOVAJySEpBg2scZwGLUfWaNofMppEgFodFiKvcoCpVpfAsSmvSoowUD+LSHTXWHEUm
UnYE0ifu7KWZ9pS6tuSlwHnQplgPht75wub31Kc613k/VVGiJQboosVKkoNrMmLMIUY/z5M8SGLH
yWzzRF2p0bhsgz0IR6Nnx/oUCVd95yVndoXqcB7Ky2+3GeOBwCdkU/82jjFzelDqNYLPwVhyL6QE
dg5RDVlooYErLC3YOh1w+TyP0GBrVdm0ABy0PqRcNmNl4Inqhz358O3OAzK+SffmCOrmusxfDWEG
idQFOSHfez51Jc5RIql875uHyBeqpSb2FGQg5pozffkBn/OcC3DDjp6PYpcxGiaIx+I4V+0P0M9H
UAM6ZseI4KG8sKKB9pIDQzwpa+RIDEsyhFQlamlC0rh04aeopLUnfbDsUyGWSt8/B0BV+IRmXf57
s493fos/+cDaKihXrpiN4KKooG8zO+X9uceCuCcs8mW4G1nrXXU0pSZx+ybgyxH63EIaItiTzJU8
E46H9PpA+ap0y2y7WU9SwRfm1fsy73Stt+YJMtPrNcdfYXaHIs6OvsE8n4AYvsYbYVZ5YIeSAZel
zoXiHkpB3ya/G0uMKe9MySeBh4yQP0db+TjGwXiKyxv9IJuGak7gBiNjcjqwryg7iGaiUJguFR8X
krBW1Cp9qFy75c5vXTmpHcrNh/n1PtBxw9Nvoy5WvqIA2MuTss5ehO0PAQS1OgWQF1G9sX+Kf7S6
DWuvYXv0PcDMajo8rY7W5EoWohmofRVFUyek6EEOIcHwgFxC1ewYdhCAh+gLlpSDjMJBzYtJhD1G
YO6UITN+XwlPOKAnxQHHx+PCU1s+OttzHilUP4MdBP9CkvBEI9B9WbKAEIj44zDt1rXlRHWBzo4F
EUb4c+21GsGi8Xhoa+ANs/iTrMYBrzQGuQB7VzM7KkVuOI2ba1V9KRM6rWYd6GsBydV7ck6bDJRm
SVVaB0iQFLtr1TJ1oB1zrfr9VvhQQ91nz/vTSFvtbNQA8S9nynlVonoMG4J8lVGYABQPjF+2Tl1n
5yUI/X30QF5YOPkNkIHuSIPUWupIewZ/854jA+7kVpIPJ17kU3TkWbk6bC+mEBl/K9k/Mg6bpEMQ
yMX8wuiJsQL5Varw9+xNK0GqTAhxWtsfH2QYjPAQUWND25zu/Q/AYDn8xPgrrDAHUEstcqaBg/5S
5qFZNoQ+bNPj5PZGmKqp0JRRf9cXcXAQ0mtJkzDCgp3Ulwh30JuCNdClVpuTIQmRLT2tXf3e2bfb
Xqy4FRBQQaa1XXT6SbYYlC8T+5iXPbug/pgMee4mRqsR+ttv0+gO+JYEOaPCq6GCAr4E0144Pn6a
bz/BFSZKqnkVyI1K6ccidFBcfkN9eXFNTgWSv8nggQQVrllS+bxUnwavmuKlOTtSgmtqNZbzkx/y
hDymtPMeaAmNp/XDGy2TcghnAvhFtIcK40nLNMVDHLTLV5zsuZBgy5eVM++jVpqEmFgnoprjFfyM
ZPU0xind6Zq6dOhW2DALevQsbTothLGL598JhWbTVJpFybrqh06wE8mQkErw6citmSPaOWoJDT01
0Q/nV6wwvLSfOJrTNMc8BbVdDpOYKS/YcUkRM588l2Jiddihy1WuHqjV0ouIuP21/g+9yeN9rPh5
dVgfFHTEUdkJfPTWZGeLKHMKV2skV4ImFG2x+yNpceRXsDX4mU6iYhjkI9rpirQfh2aYVVB3GzZ8
oEOaaurbQXvU1pELXmuM1VKKwVBIq8kRqmKzTiHBblwuLLB8laTH79oEVLhd5efWpnFg0RjQ+6o4
dXhqg3j3AZyyxdM0ThomNkm0NCXq58B5PyRigQ7IvWryCilzYAnX/ieG3HJLuINmETAMCK84OO+0
twQxbDumqy7dToF5kayOd7ba8LDUcguUuAF6b1bnXVYEbXS9CjtM8for33yFf3duH0Cgye8FUx7I
FXFpjQeG1nVmZ80x6Si1dDXI878atsZMGUjlwOKFjW85uk+5SVSmwYTzLnMZSwU5u0qtYq53pZIL
FVODKuBU7is/CvvUxvJfHD/1TXDEXCuB1wOzaZ2VFTjazOa/eDLbe3VL9cZFE59UVSTjCv6fkIF7
+jF7Xh3wIswyE28kEgstqCIsUPCcoZyOajYtrAp8jfqjOwR/c8jqh8gLvr/Ywqo2LwJM7t66uOGN
CE1k9Ycn6mT2dLd/zQMTt2kckhHG5RiGsH9H0Aq1nXknFRanZGneN4O7kyXDIcRn51+BjVnbLDmn
9K1s6KwX5C/107NJKzIyY2Y05wyNcmztONonKMRuOZ+Y/QWtih00LTSmlgma8IVySUdQOEy0+nWg
YX6kRi3W/T5TmJlq4w5m3k9f8Kqf0GTlGcoT6gtc7V1om0WaAOaO4BfhjhTHGdWbCDtiXpmQPI4V
9hDeTQ3QAtiRAtzPY3GVXQvbTOFrLykGL8UbgfLsyjphhyG5iad/xCNhHIKDd5VYZok7xm4vJa3p
2kjRa6ol+bkdcknrWVA00nm3AnAAhrG2gdONgjugbuV5vNHx37uxMAixTvAdidhjVmkMVOZsCmBd
KHxbp/x6BHoJKCh9lRBJiVid1P2cZbb3ycj7U0rgzqzN+OGiOip0n8jH9TVvgUmnhvnsL2J00smW
K0TJAUAgctN0qK3fVODbXjkyhvV1d10HvrJE32gUcqkCxAmzl6Lk5/g+LKEFGQlbIbhgF1P3utLF
eBNcbpYEr7W5TWF45LTKDPchBmLQpt2WUKGEpMHTBc2U6drctbX2Nx+IdPmSHCPAs+k7dT1PGRY6
SBQbl3eZ+zMr0MP1qNoiiTzCum6NlhOkEz7tLIKsWYYkP9YP380dHRi8dl/0uPH6RlEvaaW25txN
U7zzlaOKK3lW/NB7zaqqWU/iOyrSQ4tOobXtkkTDOf1K2EVrbCaa86r+WdnLRzCaF8rp+0PR9pZ7
oGFWhq8sYsFAknrA8K55RQl5hE1uSs3y+DGqtYq77gpkAhghA7RcrZAZZgJuKg2s465DwQTClikN
9TA8f79gno5zqOFoYrErBfLHolPRisXBDzqWVdfKYRoBC03w+bCFsrH2KyQN5KU3dg1v8cdD31+q
7NVNNOFUa/u120x9y/8TSY100RT4nz41WqecsrPTeJDLvEOyFqAX0xLgc/Te0IkMenrLnNLN+Y8i
ibH65G/5g0H3JqHVEbq9Vt6adbYlSKHTf7hK0XO1fS+Yg8Cjni6i6360wmkqWYTijeedgCP5OWr4
AlmpC/AjrcvmZ8MqQ0ukkJ8fBgmjn5X/e99X+t9Ouy92zwUKozORI4QW1QL9sKHUr/YBwvA9BcrH
FzphKeCdFThw/uCio7g9rS+79yAyXgMu5RuRmkJdesCMfqRvM6+kkLn5HHpIL2LZO5ND3RE7aZX3
HjKAKjS7fmyImu0GXCINGaKbI39iLJXxXceu4UhQ2i4YNoNJQ3UcSMKlU+G0Wf0vI2b0HNE8Yn6l
KfszWCek1UD0bmvInEvYfXGAWkhxN0MXhaoyXg8+FmrV4lLYvB1Ur+azktZ2nFjM8qzg3r5YoxuL
mISLzRKgJn5jNlQ+6FQxeh0h6E36sR2l9alLdkrdexDT2Ho1okSze7U9gSWq4/xjhU0EoNfA5vXV
p3dqB3wSd87KdVDuVYF/0uAEFQU7LobluLrhuEMCrDSeEl3aNcK/9yULTb8krP3iUq9mz4S3CBG7
nozT/yIVqizFe99xiNW1D1pZLf9VtlaM/5ZkEgj/fScZqqsm/muaKlOPJIvi7lPvS31X0DmjD7co
lm7mu8Gi1+kYEUO+cRBB1AcWTqXBUkUlYWPRYOPkpsuzhxK+ztiVlK+LN7f/26jFEcfHgBbCIr6q
Up5oZ20xXk/UKE4jr07sJqDzuSp1h8IaM9byGs1SL5FdtRsLzo1f4KYc95/0JTsyVWCjBmVJHTH3
3kDS1lYHwOSkTkDrgJDZf5N5bW+15P06TFXb9BQuFd2L4USo7Fea+8UfkS7+TpRMiGnBNxLtswed
9mELdG6HDMuv0Fi5oibHjPiKdjWEEhelMoSd5XHc7vdH75bWsAF4KgWEJR1zRxDO6IeADYd1gZgM
SFeRSDOdvUS07Y7y6d162xSAXyEBpcPLuGP5zF9TZxMl0qTKa5Rw4DFv7vg3fpoNfsPyCJw+VpGl
26w0lCP/VFryTdCcWorRSdUE+Z12IHLw6u9xBFQJ4tAqzubizx/ZuNoFmS+Tc+nbMVfOhemJFNQV
FiihD6mCXOrOFMnx8yWBiI8/GVchA+GMGA4RE39DmuLOwxYj7v7LF0jMG3GtxeJ7w9gQU9pxwawx
33gmzFo5N/biJ89qfcJcf+GsSSg5kjPqbBpN5I7xVYnsrC7+wiCLK4TTvwYUbR8RU04nx9kFP9sa
U9RSOzckS1e17f6gAgz/eYkU4VUVJmBuGmn9M8wksFQEbf8dILIxm8u6AYyp1AFFuRMNa2yHrqCZ
AHoF1JO/oNNX0t8+S9xLL24BJ/Vq51VX0RQOYcLefbZAmhMLVu4vpTG0xMibGqACIrn1+2BefTtb
/gcA/xGpbPLTeI3Jczz1jOUXM8KqLPwVfSuREJ5eBBm9M9+coaBX2HW0+5u5KU1m93Xu1PT/XZK8
ibBt0RJNAXOAciXUb01cEQ+zLOYyg9Tr+PZB8/mTJextz62OcP2Q2zYmWNdnXWzj3RG7W01EMlCm
An3QEBAvwP/WaxpxPNRkeTKxtDVBW5M/LAAl5xbXtO5yhizwjjEGTsHlCEdYoxwu/VAeUO/8et9y
74awGzOEfhn/N7HZnIrO+/Osl+SBYdz/5z7smeRschxVJ62cVooEHyg73Dx9t+a7B8txzLd+uo2D
q3pd9di58iERZzyjRDiYYL1qyXaxGmLRCtxqwDTqGwmQZL7BFteTMdYDmELSPxw4dueHiE+NzI+i
ktT4+mu8Uv/lPmRpthBnWkrGtPNbfsgofIxyViHnpAq64edKd2YbYdEIyywzfJ3cksSmg4mzcJyy
McOTyiM3QlpjY3RfpBF3laqgQgdVK5x8i+WVNIgoFA5GBmKBp7w3wqgqrVlhoaCuNqjqc7HV7XKp
WxhrioEc5QKAcgnTdAaf6FYqOgkOx0nZLYxXdAkGbzS46ryQf3R+oObcE3VgI+SS8x2FHyDcOkh7
7MJEWi2pOEf/naUFv3gPgjIWEgzHJY64qRdf88tuLd86L5yDfk/OZko+XGczdn/hOcxEv6tM3al6
WNHB2iIAXlGbIJ9hdFDzwzDdEzvuxNNwPfUN1GCv3SkWyeNIKRM7QIoOY1FEyKOvRqJDB+WCegFL
J0kCqOMf+O8AbM18OFcVntnkiBx3FNE4K5qwX1wfdIICVowYs6xOHDX7l17Q/nliwbVIdpUBJS8O
eWu/XHVBJzgsvc/YCja0Ui7gJD2zN5pzSy4SNwsmjo8ulqJZyzSJagqYOZcOmmf1/Mafb4VkNyj5
o56iQ4r4L1RrzFeV/FBTzIzF14u9hIdsjm0o1q+QjyPC9wgx/dkO7P0tn1zUzxGvzWWLVKZdZIir
Rszn7GlZICeUcnh/K2ZaTVqlSX8pX/ibGBrDnhxlDX6jaxeYqxGK33SiIKqGDQwGk320BBqTfJkc
0XP3BaAfX50N5WYNgalfoMCbXqSsGThLxIlYdJAMFPv88WhYERoN7h6J+8FX0pjab5zfXk0bFwXm
oo9NHgGsD9wDd1cbXIjVnWnlWDzVAeXoIjMz8FwKvCOmiahtE37+0TKSoyalykRVDQ8v6MEh+GcE
FpW5qf7lOo2Js5k24SkHeSeiqsPXWYbhtH766/8XTc9d9K5LDHqscxQ2/oZAN4MWfI057HTZOKgO
zprdmjCAWVGVz+Ismzc5HsBdoeYWswWAIxrHKaXPGK7XRTWdh/UDH5SRKuDUZmC+pAi0xQLqRQtL
9GEe3rneeE5jQeVQwtytPi2cooKkAxQkmqrXg5hZ/rnqOkYr22biu2NbeVqiY9Oaxf4XPbkz+Dw+
I6nrvxLySKEmFsrEWmu3szaZ2VGVjWIxDhs20ZaxpFgHwG35V6WebW2fboWzyy3OYT9N/gl6DICt
FwBmfZv+Ja3YrFU7vAnEGlKlOl6sacagO2pOUfZisU++HZrMR0zCv/RtEDqNOgIKjdKjsfLgnkIy
cq93oHuH6YN1dxtXALTJrXDShqExrWo04EoxAeu5S4b5JDoUKVTJr9vm2SvM/BCT/w4qN9YpETSb
XNg2quqUe6za+FdqHi/kLJ8x5zbCortDL721kf1znOsuJH5ygA9IpeJDfE8AHy9zlFGM5o33NM9m
FEb/3lt5ydY0bJ4O90zp6SKYjTCjMDpY3gCqz0yKy+CO6inSIEiFE4+S+NHnNZQv7Jsz1ov6WCWt
hraIsMYQYLfrAl86xOv49E+cAfFEeepSdDgSUC+jJbsNgZrfip3riVetIb0wQHeqUns8JReS3KCC
UUpKN+3qqhbuUx7duujRNypFhDE3ujhiLXbmg2xQZKN+hEuoYlAdw0QVCeynLHyWWKP5Un9e6Dpw
VqOHwGNnH5GX9TC52l+3J/v7xrfAugp8Wx1mLJ6taJ7HyqLDVDFAyRIw9YgT/5a7CuV/YjD/ts6L
SyE6JaXR23SCNjfk+G8NYmQD60S7kO5mGXq1Ncm+GV2SuSunDbc5galqcuN/tR0dcSCOr21H7uOG
3lGKrBdpWMKDw8y7alTolFdV7Cv0vyfVwYtY/jo86Q7z8dapj5Dx/4aRK6I+G5SpJK9UBGl+xCD5
e7s6MaokpZy9pebqgn58SsFcmGEls4DIE0YL5SsrM2qEFdTbKHVGd3EvJveAwsOa2LBJ6x7wyhFZ
ATDXmzNOqdApZW+kkoy9Zv08omkcxNR82dIc5Zy9c7dlr/wWR9Dm/Z/XmuwWQq+Z2r9IqWNCNr99
QpaDF5nXMn9vE/tZ02v/e2jVGsLWQexx6Mx7i3crvhF9YhV2FTrdGmLjHzTyiLnDjvpqqKR4edvZ
jSWdfw4R18yxRXlJOS3XNGQh4LZo4k1y6NFDtw5P2JDY+YBWkSKikA8TvjRKbWewTSg4bMCb/nEd
v+8k/hyjUe+EdWxaO2deGirzBE/IfslBwkZzQqeeAXVhAFdcey59kVT83symNZQPQGm1ImPtOHgm
nzhcsMfFYH7jcInq+pWE6KAc3xqqWFRggDVwMvy6e7d1jI/zipOzv5t6G7YfbcZYuUUH3YGb9vxZ
IY/aeWGQU6veJZQXlwxmJC5KiLicAOMegJfhi1G7AUc2L5yjB1KZ13nMe5SKdjikJfrxeqwSXVKG
urE+fEW8TgVJyLX/WbaB+OsNB+v25Ue30wfxpNzDH4sRptTmUlT0lUAjpJh8ZnoZ2QdHD4AELHUX
0+JNrjzfUiEPzC/iME3H1uv7L5sbwGU2QHaQzFgSl8kpl/QFbC9bUO7yKtPIwKmYnrhCjAQIUpIH
ydlcuLJEL+89IXlLcoPfmPXQXtlFWSPMgEKeEx77mBq7ldvhVm0i0aJ69J2mhgJmOmwPYCCjHZiN
Rj/iQIl4HKs7pzKgifHFLFra7iLi/m3GKo++rvzgCUWu4Y7MFkqc/tmMMDuQ16SFnZ+Wle7W3Omj
tD6j05Gbgv4gJKcBIIh4sw71BXbLlkMbu4++HJKP95V9uB3NStbir3iQZoE6HUcx8B+qyXGeMelS
Mqp9E+ADsKz3RyHTF2u4sX+/o+5uRyWRwQAOiYX7ptRDbGsjmy+Ca3luPgEFwrxgAnpnu+NrNptp
dw/8bwKqBW9zR+7CsttuVXl1LRDdB6fBrmCxhGOd0aPfCfOrNe00PhstEygPOtzFrTvTOga3k99z
G5oO+KwfzKJ/15OuBr/T+zbZNfQ25lOyivH72OxotMS3Ul/+HOhmnEtSME+2/VLwl/fEyOmy9W+1
lE/mySXFb/8ev2Iltht1KuBSyz6rZj+7VPCEJ2Ik+eRcQciYBkQmBHpdkYzyljGmGUUaqDh2ZZJR
goro4+xFBIX6zwXylCjIk2qQOAPPqX++pggZWvifpAil//yz+ZdqJOa2yAqJi+2ASkINiSgftBue
YYRlSzRvbhIn6/BqSFB+5YQLN9L2Q0DyzgasOpVNxOyN4TD3101nWsbluEAL0VzlmMGXEmqLgecV
TmDJNC/GGJeL9cMhRCRjQgutaD525wam2w1hCb9FjebBU2QFLqdBl4QmXsQfIs2U0fwR/c0l2/NF
YDFPy4VmWIrHnOApLqjWA9tXJWng1gCjsULPxNgApLVcTK0FAFI1WYV47MWVEnv21IQKAqUTWoTr
WE8iN+J3dQOavGYWUveRchdoVuxi0e3wz8wzw/HSEeSE0V+L/TXfSPR079GEjp0lPbeiXEeXUgyt
t3jYUatS/BRUbcOMXKmJJoCw6DW9+Ge+N+YiYrt68VNVYdrQQyj3PsD8UZ21MazKAohqerzFj+4t
wfR4sO0AyVFzP8BJFTji79tKQ8Jl2ubVnfw7Xf8vNbe0oFbRkr9jaAVVuWe1ZCTFVcc91JHp526e
bTe/WiIYtF+mMDEUFb5Sn37M/IgRybgzkQkeFubglC6q407TFFI7AbjZuGfhD8TVfQXD3BfUbhs3
6fgF8CLQ+uM3PibIIjICcwCp+b4IWg5R/lk9M4CtBlvJsDbNoMsxh6tl0ZQZ4svKtFBwziM5ONNT
M5j7WPl8yb4Xj+rrhgfWjlIbFL22Noz07H5CaAZ9j6i3uo34G76dR5zzcfXhwJu9CT5HpIUVwx57
OcUoycs/u0TmCh2miqJNBcGOVhSvtlUmbpuR8FcG3ja71hXoY9L9P+0vSEAvCnNNX0fo28ScLueB
F53de/3+jzuETNSfIm9ftLiyY/pRa+tvq1oOQ+gYRa5NseDcySW2X9YAWGAfluX4iSOnpS3G9FNN
k9dUoGqJaNETWCIt0UIMDfPjdIfKgTnTr6unmjkr17q/JfR8VZmMmVqTJ60Jf3auiQifVJwKRXT5
hxgMZOmsoJZDbzG+ewcXpDTjMC5pHBIRXA8zTKAKK3bMH68eFO1N77Y+K/tCHV+oxRNr+tE90G/x
Ze1LU0lpLbeFAIm+T5T3vGpeP4pfgy+RP1o8LRzv0GnKvHaOSIi7C8YSgWRgzPEJRhKlkZ2sTBxF
fGmCn4130hpLtUqcG+cCSVrnC+D3aQrtBsrQ31W2xBS3BiogEe28LeD5FyLXg7NPRFipyZY4lOR4
eWw7zVoRB1WssVQq7Poy/iAjTcJB+WoCZ41YsH9XM/LPy4mwZBW/fpMnJwiHKEDZ8eXyFSxd5Zch
NUCAzwObo7CXt+QkpXuk1v7+orBRqfocd9LexkyAYNv60vOXQjIW+CPne7uoZkPpMKrgM3ULMhhN
sKwPgArOuyk3487AgzkWlL9I8akGOL88Dmx1z9ej5JfOvFb2cEpTskVGYL/jofBw1/l8dg9chOCc
fxfNq/d1oDZjr2hLINVXM4M06IBKwNAqxG0php03WauARcP0Ry4NVCG/uIVpRB7yhzndX2WOAGtg
bn/MQAVjuK8JFXg6CrxvzFW+hyk55mDuNnoilu1txB/RXGfgfxbbY/aIlPlztx5wCt2T8b5NCOW4
2dYFJterx5anMX5LcekWcvP3M/iiKofr2bKdkMAtpgYUvcTGazUPCDEuww+E1nt2Rr8OUXM5RnqM
h2gROxmj4kpkakhZIMDeiTFMN1zfNO7kCz5yW6guRuMJIC/6XLIFgK1EXcPXURYppnuajoycLUgH
qYCOQUF8wqpw7+paHGuHyTPMaK0hUAH8jlDUwgJFtIh20GhfwMWYm0HpOklZnqDjFASHKRS2t7uG
Gwai5x2N2UiBeC0IPP1Kx5nVD4wxCy35DRd+yuCAqAhu/9Rt86lXrkxisZmsQsWcYc7b97/hTaWU
SKLoa4vAdDdukBRyLAm4QqKCJAX0mk+pknI1YeiHkU0wLl0qarvzM8Kj9wcu1JNBodUDg/YPGwo6
uiRDZ8WdIzF5oPZWdBDDTSJfi0zdTd39MHksr/028MijtHdz4B7cG8/47leEazu+Y8wamh/kvj8R
qlLI86O7mEJagxinNNl4oyiUdcBYi3LchX8ffxcyQXTUpP34QWBha/B3WXlWPesnJviu1bUmxqiX
c/n3hGtfwXHByquB0xkDdcD1QeJf+IbpYiC8fUp94sViCD3SzyEwceuIb0Qyi217jy2Mv9hHcXV7
gIaRAcAY7SUxGT5xOIarKVSi1IR89hebkn1PJY+zqnZ8banWsPq1f+vvdeqoSkF7+qyJ14NQbjZT
TCESZYzynYgyfckH2HMDa7BJdBScEZLRIH4yHp9o8kW45mRDo4MbvncMjm2iuA7sb8j+sqEBk7yw
1dxtxKVoAs4USzPafGn7J9UGcnjF/RngtgudTCTS8vQRcj3ePRxPWbBMOUwIkRi8Z7SHa+ky4jT1
9mGVHMk1p74NkI2JCuu7HE4GnYqZlc3Tb6uV1naarM9EFbxqInBB0t+vDeeoS8gGjhJ66bgixrJu
G9p0IbMMw7fBw0BphJt/BQeRuaAzSTQ2hMoglsG7X8Kdr9pDXbXaOib2WjWKDAbz8TMvD2okGqRv
zWl4qRGuLSIe3sDN/VoV7tSmuHFAxLNuQr9kqhk9rjiqACahWo4q3oVP7TlG0vbdodo6BY2ranvy
CdpQdnDEeHXDlRtoVXhcaKWCFAuR24m9r7rz8iyBvsvbwFb4lNZrPGg+pKz2irw/82z7I05ITbNr
fk7u4sxYvIwmfKgnqDpxI/VNhM1VD7fmOoYuKCha7AHtv8vbLKHfVPrXZioH74gNMpVZ+ciK4AIv
1tzeFNcjkoE/EBocZoDazX2zw0R9xEfrknlCCJGp9IG3QZ0ag+56SRB9+J67AKeh5EJGlRbVoFBU
7IAjnXVyQiTcK1T9wmnrc7YQ8yx80lRmfTwTMF/fMRkkmFVgc4bXrvbVCgUWjUOaNe8U3vbvgd9Y
O9tT4yJ83Tut3i1/aLHfbokWwW7O/QP31CrVD3fEqqlQC8GRiwtabb8FQXIDTJOBAGGzugeRpnLR
iYGRzQ8Ltj2Kyw==
`protect end_protected

