

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
H5lQJsJvaeLLGFRhK1oe708p9zTtXNXItx2KAtknEaAF2yq8IXwKFiVPbPTO8aJ4G1wQZMrKgMvb
6zlyKbmneg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RUvUfs9jruf9OSb6utxk79ymugfgdQ2mgDnw22tbcF4+w9YY12PtlphQ3EwSjE1BR+YNcfcg2ppx
nVp8oQrlHaYHLiZdJQiFcET810isTDBwI9+sjn4Ry8+ftUrGRDkzGQghSG1UFCnSyA55dNVCduAa
//ZGtYPCXRggO0BwEzM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GRoj0md2TTeeyD4XkfgAjr1JI8z1r2plHgATS4H88EONpa3oaJwG10L5TE6c5MDXVxHb/m1WeMVh
VBt3w5S8h9pf8c485G3a+NVnNsA2vHPB4cEC1yhvDIpNkeqj7HvAUARW4zUkp2MDiimsNN00ZMVQ
inLzBlDW8A6T3Y2b3GmoYzUXaMQElMyS/PaVNF6Se8+PIRjTB8Dv5G+A8K7PF3j0h0gW5LdMZrCx
isigyN5NiqJ/3ZZGLkd5XiuLlr0DetrgHdwfifFeF2dmLtMjIx4kUkMG45tToYmkQS3jwm191cux
eXIUgmzmvPZHik85i0iZegdiOZ1LzY1yO5OyEQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UnEKB1f1t5V+eYV1nijBv/smbMsJH58WebxNSKYwmtj2m6R5AlGEZE0haiR3VYCxPRjmiopDDdr6
uBQOF41DIKvZSm6YCypTeVt9WvkLpXTJIiHnLWz3IV+uvKXohhIry2Pg30NMC2EWPfi43aTNvtNH
ROJrUVVcDZeGvVPmgRI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U8EV7GGC48XxGZ3G4wShg05dze1bZdqSUw7dITFWVJl+2U1VEqYTGCRl5zpa3cGdqM2+nFugC+BK
YIux1TwcaF2Ng1I+Bp1k4H3BhUPfmkZlNiGri0KnFOiDYzBROYyyiUUX4IECNCLZnG/OtNfakQoI
AjU6WqtEEQ5JSpZpL5mpGWt7jGfdl9gqPeY88IdcWnasDywKSPqo47azQ0KIzwP9UejnEHChmHgr
3Gpvmrmywo7/+/EQRujU1oGF+ysfAmqchOGtHLtDFJ1h2OjLVkv+puXArlpXpB9wZah1XCGw2FON
8d2jAO5M9wEJ2bQpFyxmedBeZ1Qj0cJQKZW3Gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51344)
`protect data_block
54IuO9LEGZP68pKxkluM2vKNfpGxZiKaMoMpPwH28fJ2nD9q5OH+p6NmnRTqt5v4vT0qRHgaBBbW
pD4QFknXjQEVyPLEKYAL/j8FOAUNxJLaSnonXjK8hkIwTQJEt6M7Co6isKgM1xzNqGc+6YlFKRjl
2JJdKQi+W+iNxyVPzwUryevTRhChlrBf8DhGc/KyzDGwmAlxQKi26Mqs4JpdeyckaajU2iZet2xG
pODv14Qs82bJEQNZiJBNn+ak1YQGwIar7hHW+wY3yQcj+oXMiQgH4uMO8aTciEFnBv8x7wk2/BY2
FYMTGxoEHpGUGS5MJbbIhnF2gic1yC3pzdZG+k/r2h20q41pbOD5DkKUpSMcNWfQWOP0aUMlLC6+
TgW+MEXD1Zw26VPZFv+snJxYmA2zcTQUp2tZJthiAiT3mOtAQZJROo/eLt/rPFE6kgrw6iZ3/tqh
jleH59MoAOyHVnQizqh4a/XY7Mw9FU8zm3flS4ptRJLDj0CjnZQ3udFt9x8UuLYmrN7gZ6xTpyRa
GfBPrVwXYj4OTJFIu9fNYBNndqU83G5K3FHi1PdBVRAGn8SqbVcUjnBbT5al3TTEE7oxBSvnplTS
DlHVrV24vQzDuufNHuhNpQOZqgVQS/RpURTleJTyDskgkq+aFGH5G+ADEtY6fWjDaONb5eaoZL9s
Z5pRTKelrbu9Yh1tjJ5bzLheT4xQFlmBCirAKUZdF/PelIQmiAE4Hp23swnWMeqBO4SrIocNK0pC
sD+vO0UvRIk7FheO7xzoRID7EMPMcOOI3FNEifmxOjWUJcsbCVZqWueP6r8YDfXiv79BbvsFXFiU
EDVJseycyBbOZ6owykIWYYV2vcaK43orkOOsAy7NP8gUb+dNjIJCChV0ETp6ssOZlo/6tO3+4R61
y5LKrV9CPl6mofgAAWI7hvDW7/ym8z8b/hWgiOcTNDrdTxYY8UsmJEDTvGDeinyTVnK8EJQEoR+e
UBnfM70o0vPAFPfYAQ8EgFU14JrLAgUK0BVVVeKMmrElitsgQ6mFMeTjchvsBERwQdS7pcy56UIM
DUbrZkp9q6BY7V4OV25yaKNqedK/Wfsn7syl7OXHwQcNTBzDAgp1kKDbn/QW7rZLXagGbp4Fa9oG
hlZm6e+bbvPt7OUd+fFnyQuWrZs/DglG5OK2BuRcu0v3dcYXpq8cUHT/RuDPTKm5wHXklEaj9YkC
dZEzqE4sASDy5S0ohTZSz3lN0k+7YFx5hW4HxP7pD2AFmM2Ach48ilFC6e47K9zlfi7fxef0pVLK
H5tPs5Sg4Zt00dGPNHX8FKlT1cFPAkxlq7sNQwVnKbswDHUnpDP4JZuCRK1nZy1urJu1a2jMwYDR
tZzbRdZqOwUVIfMthvcsotXsgbnz0WGLkBdFjDWiJVjnONAs9R3iB6SxKvXBjiBn9MQexEzCY8o+
sYWEZBj2UI/BCfVuRkrH5obNv5bYf1oD4Hfm7tEQvdHpOPODynnQbVkKwEIYbeQuqYQHLFZBMTKt
Vc1sd2tBjNzuM8vLYhaafuFzh0Ysk4SZJtPjF7kFs9kuCPLW0EYp2p4eQD+tYHj1cJKeO0HOZNlA
Z78hFf1CntzaxxBKQafY74l1Fuvx1GH/BPIEHz6kAdvkeXZughfoPDAwzHeuzmtTQLUY6+o0G3aT
FL/5uudNBmg68sayhlRxvU1a2cBK65eHKRrJIizvVDyeIGLt9OeJxB4MF1gXe4DhodJ7qiSX88LF
9GHhKq/jJISAdtMiren2hpli7gy/zb56071C38M4Zb31O75Phk31P0tisZD0A0tfUakrhzQraWdn
91suPedZxg1XSf/rOJbWTLxaO4yOJWFmCFeYNou+ZO9j0yR/PYu2zP03ugH2ESbFL7jr0heXhKev
gbuMo5l61rLZ2N3Bdt+FTbZBYFgDL8HqTEzlDRTA7k+W+86zMVWrQEBqkxJuHxEzsPDDHc832Gp7
Vj/bpnjOcWOLL752qRJe1zRn3wtDwkSI8RswChuQ6J7dkweVpha9ZJA9B3VPGsgRBUyXaXAFbiQ1
atbE/Q715iUHEpN3mVSLlfRzzoXlwcMffTGULcBN/snQhqjGpF3h7gF7zWCbYCxf3K0e6/XmnlK7
atiXr7MngmN3XfxkNwIlRhO62FAzf8KCBNIiH4YxyMEBauZ78Y1+YdhXiK5Q0T5u/i4liM7WpMTQ
15BznFY3nlSloZpT9SQaKP72D+SVksR1LcHwaNA8Ody12h8iWtUycNzKsPhpnBhz0VRVK5KYXZdP
JvOv4xqkfqU4w6ObD6DZE6H7qOW14oMNfo0XKtBC9YtZoZqPotQLLGmLHxjbneOw4QKOK/UFhdGZ
vF+3TtkH9cwX1jyrubgeqGQxXmUNiHfosUx9vHrOcTtDHdGqQC/4tOmwutmc0uwqmjArqSot6HbE
JE6B3xr/DFvEZY4p7q0EF7Mv6j8wVifaLo8mF+FUSKqyLW5Qh1DszzImDsSeDXBjbIt3KeTuXnOt
Dz1lQYrDA82bcth0oo7MmZXRtKZ0F35CvIngp2WigB2qcKd096AVNxbksQDCoSm+7xGyyrX+4MLS
+wE7Lyboso99ELgYZOTmeZe+HpcVVKGCmnUUbT1aO1po/HwLG4GS1+JCguS2AK+j6BPR83y0+xKF
IAnOEOzOdAoS9u5dC+sq4DQ/5PUqIvjigSvYzjBVKQ0U+lCSoyUF+A5PuwxQ4CP7hp51EbbldoAG
J4LWrHj7WiEQ+UiZi3NxkvTiv4EgEchPsF80d8v8cgHu/tHvIBtKSL8h+6Y+RV47ZQflcWdmXuLx
3nCPOmcLtpCsbrEJUAWC42eJQlMFC3cgfNgGlj41GtMl0Q51EBg3yxR3/ot1pXp3DFNzRjFkVswq
JBiAztiS9D8M6TMv6Corz/PvlcZXNpV9BigNbPaWJanLLSZo9TVrF0L8RsvgzbCTA5ea2A6aP9Um
b8Y9R4UZ5cLC7ygx1hXcrj/zeHWtwK6EG/CKehVReSUCxTkFXVqAZoquIPAg1n+z7mZDo0J/aztA
Vs0seXgQp6qNroQ4E8O2zRYGf4IHGlK+5LxyHw0jKsTgeltPrR4v0QMilwN0mo877RIZrggIpLgw
mgvOMbdaudiVqEgTWmlFgx6uTi2kNqNs0kg/HgoPwB8DPvztUUjcNJA6GAbGsd/wsYJJ1VWEQi+L
SfiHTMfpz+YAq2MqVvDcO+hXz7552HNDlMeiyYKAvh/kOZPFgVFjUYbtCIikbadKH6joy6R4MGoS
cXCKfoDPSfdwwCwZkLhNjh6mbcNGsnrz5D8VjBn3z1e3UoHa9BpEnevGHqelx4rLAcDo+sFY6l2q
VhHUBnGL/B0taDxH26YmdIQMlFHZHHpT/vFXa29HnHkDY3UAowh52Ha2+1a5Md+HGPU1MHhN2/O2
45SYJlgcEID/TZvrsMabO5KKrGrWCMYS+aKlqC8CpAYyDeVdaaoN0hr0DF6yvrncCwYGicObt16h
zz7/Z1Wc9qNv+3OyNHIxyYZ9TbMRy+8gw+y1f5Pa7ZfDgjB7cJm1NEqYPdo0wQhIDF/ApfemUxqn
u0DDnhEXpSqIoT0M1p90WHAv29+6XBer7fLpOG9dCSAkRV9nY1yiI5etFbmmAfd6VZqAFjs733eT
06ab/OPfiU52RuVQAWXMA68hYTxpp783oJrOI2YKs5PL3yzJgrjaaiyXVyMeKqSusUJ/mICumoW7
DJlrkQK5yXxZT6iSpbWzvf+RICA7lp6GPLcEjbSiLKtkkxn1Z9dsKd4rq+glM/LZrxiN2kTlLYKR
SiIFDkB7jTLtJQbKiPJ+mS0+yHhSzVKU8du2E/mEVqIxSj3hQ3OLLxKuD07LHjtHdWHfaPo58ZJO
e58bvnIiqgkmHq+/EzwyQSMPZtyodzSRnZ4KiHg3UmZFTmJJ3X5Ao1kPZ9GTkwIMBZB7Pk2CK7Ze
AEtwsSRXpyHKrOX+pTCPY1tDlqGo2aLmcYtG4sWq70XD3r9zp42j1/vWkL+akqivb9/cWxBuyV0W
aw8uA3Xdn7caMkaPeYJbD892FPUigS/jM4yhB3H+dCUMBQppQmcrufbvpMQF+E/4fBi5xDxtGjee
73m5LaMTcvboCxArLFpVykDcwWrGCxpr3d8iBSxpi/6RZ72nGt01nE3mnu6BMXoUi9yUi84BLV2S
sJ69rDaLLs26tFVX9xUZeF0pv6j3fxqlZTRcXP7frCnSFIYIUoft2CC2qbW9tZLvjrXNdz3EiAhY
fJASrv8ijNBLkEQWkp/yVgbLM7jx9xTjb4FNiAST8pjyYhLKm/zu8QOAltdjAArx2qFw+PzM3p7H
fdJ4UMdJ/7WlbTeZ8rVS/45AuX69j6LecShVoDxYZfUO45C5pYFvLlH58w1/FANX4USxKI+DB+D/
gddRYhuBTC3oIDjowNO8byXPpFDWcODGWANiFJVgZYN8yzSpg6n4mexKfVAoLUHvNN10sPpFsSm1
ar433rFkOpaJSIfN/S+EqW9MzK0uVY8/8zkprSvy1CcKO+tHLSkOUMUu5H1JwIr9cr+GDM8bMJPA
37zHAmBVoT3A7slW7f+j67YJFt+ui7grVvGMdtK4wgv8N12Cnslf/l12k8dRft/chsUni/0jL4gy
9+5D2cYTw9XmSKEybrG74GSeDEeiiRNacAoRbUNG6ef3b55Si9ftkDv3ftwF5qZU1/mkdgWud6dz
rdyXUf5JLoYuOYJvmO6m05QxdEyd53jUJeaobKeBoebeAPdIuuSJYtkRhruP/wTzEutk5/NqXCAO
K9A7OWfbKFgLatcySmGLLmOuypwdWaENhtuOyfgoTbOofly1b64Z4VteY8cZEYYbuZmmCi7yhyYu
7OyxFnfgg3onyPAkR7ms3HHRu8jeSmYlJq3/zOFmY+9zgWyLo5bhER5j0lbmkEdTC+SVQaiWuFDH
hKWUJUPxQaS1uLToCxWM1ZRhMfEDeHRVMHr1RS177apHyNqHwJtmJQVVs8ko4NHdWGWkq0/bYfML
VgfW2F7Z2bI+ZvLKL5O/FlOY/lRqsWenM12FkDoViGrE40a6TnvgsKE8I5aQdAZTjWe8g6fnqHE9
gUvVZq7UlRvKAMeGCCfGSlocCFMoVjD6JLCrMm0h8CrR2cHBRXwYq1YJpKCk6dw8dB3DDJPvAi/u
lpIeFXlckfDZK2h4WKDi0EfO2CHOeOT5k6blTEjD0iu0XisGzC7qZIJS6zNq8qLW5OW43E71r8+x
XP4/mwTn99RmMSnRCf/bcdY4f5m+n4xBZNOZ/X38DTmtJb4Cxx97oRMreyVvdYl9jpgWPYkwbWcS
rJDr4xKCEsbJGOsOG6UA8x5R6vXfKvG3Xn0cw6P0UeqhdAnR4MTXHmT2l573h1D/eaXGSiLJRKzf
ubhlRtT+Nr1InRkqah/oSpgh22ZvlozQXrrgscan+thtWrYmIklnQ+B8HxAJukbZ9W+b2+o52BRb
QDJOasfAQogutHRBbLivfBnjRvuFBfnxZPvFtH4xzkXIxyYcgQZ4rHvtq7aLTSGeoCeBPa1tUmRm
+30zVsDzpZrs3lBEdGZTe6t/A97x0wyAg04fwy9oo1iIYWOZEeN832Q8qCD6RGoDBsZlGqWc/3Tp
JtSPKZustNAXwSNRLZebsRFosqKfjmbyHbjbUR0AP0kVFwx2Mg1HskfCmm3CgpqoaEXh9IObj5fr
SGDOuiHvqdgj/HQpMlT3nHEplBolXJEOuwP/TFOgr7vYNcsne7W88np/HWSUp6oWSd+EUPK6HLRX
7Fnrjsm951cWCWTEUNalG0E9wy/uUE9uMhpF7MHnZqyF54CcaTCXuLWJSWOsIotiAl9DWaXUFEAK
yQ8NEj9AwPz7zx3DoB/fxT6LFXV1w/mBqfKDL9+maVHumAD45XnplVYDTKbQ677dkY2A/76NL2vw
4XBVW1YpnT5c5CyWhtn+JYz0Qf2JwOYLwnmO+3C4RoKtKZDDUf8sJx9SDf8h/pJ5E8N9911b5bmQ
SWj5EYenOMTseShSy/5Jn3LEmkQycKGrAhtGdcJeVYfUAuBsxBDxP3qP355SWhbtOeAVlJR9XeRg
54voEEyFI9LnIPr1du7iAm7WMcKAxtTpHyQO7TY2OokqkC7K6h6XOqxu1iUFnHJQ5PHlec478QmW
YUM/DBYORycUIz/rNvK6RExJNK4G0pmPBSg4uYVh7bwqObo6KLchZ2/aJevGYL+tZmonEN+MR5MU
CTpqTDfrtfTKaz1laMnjoq+XVo/J3eGfuVcU1I4vioVPRM97O92D0kQMYErzpMFf8jMfWSXQ48Rr
7nQkGxr812kHnDg5j7W95uX+lSVPmgTDiMg1i2LE3v+bgJMQJQmxaExOz63CAEweS6js1pTbYlP3
AzOfStXkidxo1ADnbgJOk4dlKBLQZNJcQdMpEihc8Do/9b0iSlu4WcQL1qkI/MyhhCxVz3Lkn8S5
yUxCAcpOGHYEekl8WC33KfjWCRPZSrsBrZaGAfbp1aeVBLKF65jzeeMBht8Lhsedvm/vNIJwKwyE
O8hOHpC1Fry0Wh9s21/IDR1hshk647R+d+0FpQ15sC9bmO/gZBfFXopt8cqDt7FynVe4R4jq7maN
oF0G2xuMeyhMDEOjn94m2WIVEtS4aR+XAKB0TfyLST0youboVP0VGYyawFfLDTCkjabcXotZBoE9
u/7ZYGlMpfC07CwkEAeeHGgRJbs0ce0eLjP70opJLqx9/xdfE/42yw1U8exdpYnuhnN6M6gDYsIV
0b4E7K1XwXavQVLkt6OCIolgG17NxGwpXNIecaRHfbTeseqC+hhhEjoA8wvTMoI3tBElE5dd4jV3
DS2AKa/RBvkPPVgdvQG8OrCU6eUO6+6TuC8TI/HAeluMk4RxLHI7OOBORvViE5ryDfDLL+pLu+Gb
8eUNOLqyX1j4CF5HQ08ypbg3491Vl6YUykjddi/p9S+GAHKkEaLwtKEyD1tLmMMf/709EwEEWA4b
HCXjrxf/D7mkzkmWCY/vEeFPJBTnhPAvcOJUJwWETEwQW096ahg6D2/Sq3gwwyvaiV0sD4hgmqor
w8XHO7giaN3oxBwlTTf6+ELz0Xn80st9BPHpg3uVSH2PRnTculwnVb8RoXIonw1U6UBVQKxugEhV
etag2Y/57EOJDeXA3zX5G+GlJilRAWe1KMHnzdCDciDLKhe8gEBFMre39xd/JozWZzLVhnHE6tIM
a4KCZa9yP5ufcqDc81HR3Ed9X63cvDuouWctuSzlgB0WNrHsxJ0F+Pqll8hAV5jYJwCWlzgNIDDA
kmUJ8kdRVCmC9PJeCVoEPKKz64oFsTN6Kd5KTpzqKKj7I2A/mTrs+suuo0AAAhsQerfvLbS//8nj
FiX76HGKD8Ku/iMHNyzK//rmkfbSuik90baZKVI6X4N9hJCRcS6S31GMujgJ+XJNBm/F6n20m+3Y
IhnBPgIocfQ6rZVwNmYHTw4Y19Fcqr6GFU1H0U+3lQtq1p7uTr0YbOtyYGCjoWgwahdAwBA+j6Om
qFyxOE4W+/TIGH1YtkX0fsQFF5/LK4/OVAfa5iLIFjCIGOpPvV9y16kLb0y7XyVh1mBDiQjL1UxD
aD9YcXQ8HJ4c735iACN70HyHm4cIHmLOHxfoJmUG6iJy8rRy7l9C9YGjDs2JjregDgSPdUthO8pK
v+BzPW7T3DeZUcQHGrefTvZpu4NkScxIpY1F23vvEbyNUKWhtaFnE7n5BZaKidOfrKZ63UnvCJdm
FIidcj0nTdN8D9/IDXbXSb57zJ8tGX3xxv3wz03zDEsEgSxW3/UQBkbm5CmEsQ3qzQHJngTvio7S
55zDjmlpGqCMzDSEYGDmRp3ksT4BI9GGQUlo9NaILvp9+XggXJf4PD97lFsHFsLrAq8YureM+kJH
uFQVkx7wlUi9pHCDf485cFXgXou+kQpDOv96GK9t6CCIWfOi998tSULcuMvmftY5Llo58C6Z+jOm
G+9c0ZVg26G78fDuOw/Nvl8dLA4EITUoaf39UewNMUjInDjuOAxc+U3CuBeh8gCZndtcyVHcA5tk
o3zOj6f5zszliQBOoncl4soJZalIJWRTG73fU5lA8vHXgQHmyzvqZSza0bfzj3DSVEcnFKceke+9
GdUOl2hY/XbVLsBygKXx89aM52XVilN+oQV+NeR+7ctjGJI9tbLUTYR3A48UXmOOKL9MEAi/YEs0
vZxldtwf0tqma0rf4U6fVu8FzHL6slHv9Xm+HFP3nbg7/wGejbg7CvxPJvPW0FIDS3oWsa6rKWmB
qx5o9MGbS0LPgeUt/BO6X0b0EvZt3m/78zLo764WlXstYkemD+P6mJALUdt6uMt4OC2Jm7sRV7Ot
xzQcOEtR1ffKgV6R5FcnHKx6gAshHevMtGqgfzh6yIQ9XaLhFFLxAhnKjbj/NUIBvZ22XbNV7vNr
lmkap9j+abp56c26zaA0yWDfIb/3vQAquuHnQpBwMGiibOZdLBmV0qHrcrbxC/E/9Re1KqN1SWAN
5nrdydvyEQSwUwuR1ti4Ifj8YGiUbI9QUF7jwkfI++gbAcABIWO1Wg/8qVZ/LXsv3jJdl2Jywnpj
DVirmf4ZXBpqvBwGU47/G/5Xd10lT2lEstEjCi14K0HHAQqhFYbKVk7NFGYQqfnO9SyahpRGxBtU
lJHTfbElBCwZBOWQVl2ffEO9vnN688bWD5TVyAjs6bb3MmsB/+pNMBT/RoKGt/z2098zsLf2H0S4
h8e2AO99SPBWOt/Ej70XDHJT/7F3elBUKUwHmkzj72jUVr5Fbf2UQe2nyHGF4MBqcFG+2Fv+AM0M
XyTy/P/MF1gQbc8t5ndFYoDAh84g82bprGbgDpyNNd/TtuKP7i6NiaM4H289OeY1bGgQjJP8kvoB
k/eASv2qZemzBVq9zcQK4y/qubUzN7qUUMDTVeisoq8czPrIJ7LtiCBV3IQe4KJlFzhBS8f1UywF
H4tVmY/rUQtzdcF0ijgQzAeOyRotkVCP5EBy125u867W/8nMqeN+yRWu8D2S1M8d2qxeunzTVvdF
MJqM6kXCeymWBTgVFMHFqgmW2jCgpgd7IRNA16bAhSztyR7oEKMuM+xMwC4IHDJynp8M47hAWu97
JD6Bi3LiYp/p6K+KZaa4+/frGXBSSbgR7/5hlGJEl833BM+14i43n1b20gTmY9rxbqCLNdxOvmp5
D6axfMRO423d5Ab65K66umg0KRQGjWBps3a7jW7XjmQh1gtru6VNpKQHL8/mr46IdIh5gG4/rxin
UAlAbXAJfNM2Xg8RHvHOouGicI6xO7PkyHX+6EgFBFaY0cNK5iiVLrWEz2VxKePP/rEP8GUlpma8
VKxXYZd457VSIEYgZWs5xryr/KaHdKDh5TkwJP9/kDkDT5TMhy/PQW0Lr559cwfj9xwa9idfrspi
7+cxO5PicQr9SA2L50CtRokKmXjespwO5SGNzpdUEuGH10KQQXEXZJOgbl3CgWnD0Ixfzh+Ks/+5
mKh+4oJzHwl/pKWdqITytj/y2IW7/21EZwLbNgjHdCPBE79qOBfFmpq9E2Cn68i5aD1DTTBex0Pm
f/CzhTcc84DKY4VRT6CM8WDDH5PEgJQwwwOlz9BjJ6r7VkftwN/kFXBCEyusDsT25pzp0eX71nL6
xw9PxydG9KgQUav/iEO5CqHKNtwM9YAv/EFEyFJKwK9D9Yo2TL+0pwlmovVWUAhlQ8FsstYOaUJD
dcLjjh7rvX6fATBXOwAO1ItiZcnJj+PIj2WiDRUqLXY9uXrR9JOrQOYeO9812ckQtopdCckmxBFs
5v2J0Wv23oVEFELuFLnYDNRvmIpIdkNuyID4H1Kb1hLIouSqwlScFpco1TU7ysIlsPFPEwTFLx9i
waJDX5D08ahkqriJeNpQD7C+Tko05q4iqA8g8rGrxm48J7FnNUmAXdpdCdA9fewQPZ6hKw3KGwYY
wNfOhwvcMeDyjhWVQsdfHBa9Rj7pkleY0iswZZraZnIVqJrpllEs6iv9t8R7ZJ6Xx99LpHt6wYSY
pv7m7ngeURyLuQTfGQFvsjML68KoUFbmuc4TVxTeeGlzYyRxNX0io93IG5IVdBVzof+M1XT1LLXl
RGXI8YTD079SjcQUmB4cPnuKj4K3pbtfAlQJE4JoNVdL3l9OMNW6Z/WRajxVEsqMBcInqphwDpuL
sdoZlWpKg2d+1vKjU5Q2Pof4ra32l8yJABKGrcVqvEWt48Y7BEB1LjouepyK/pZhMlMcNjyB/Yiv
3k4YRBXp07hbu0cgXZn0NgPq1k8SovAwz+tfVFDFPx2HO6WqSy7F/GGOA+YD0yBRMAt06wwm7GBF
otQLMBAvrDza0ja0J1UbnYKXZnory2B41/MB4NwgHhyvomhrKeF/WUwXsCMCBWY7SvVCjgYHbMmE
RQ/TaPpzR6hfMKTVRhLFqblWAbCRO733vEdOA5b5zUmEnRBfss+Zsx3CXoh41xcl+ZTGNja0fpHA
XjL9LTLoxgAAelZA+Ni5xCnQzvqzOHMIGOGWTt/Bj9QtM0VT6GZdj7yLE76yBtjYg22Oc4zyJcfs
DiNY/XIDpBRSsYbaxx7Q+ORRAZe8/jXjZNoPHeLLBcKglfI1iJYDZDUhGHtq43Wmh7A4o1zpXm8C
q4RxmZBT6jloJ8dozh8U42G83E+rrZAm1umq+ZMxyiVn/u5fcYbWqZNNrCQVNGX14N4cZissZaBC
v+s9vcKbfXlzTM7VOu0nSSfODKuJLAXj/ERALHBAY2PRJYHGGsNX6LB/2Yl17dxhNmFh+hT78zF0
XjGw44v2KUIgeI5EfPXvQAsaOpYHW3eSIfmNVDdyiIqsxCFZsQct0qLVbjG7BEkTUn4I66oluKeO
js4PTEHtPcZ9nh9Tplq838aRvmB9tGf5zpaIJx1d4Y/xMWAX3kFbAprT6EZnT6rjRlwHRNTyrMf9
8Icfw5UBYmd4u8lnwCfW7myJbYdrfwvjxMlJgIHyzzvZLDhubF2eA687E0GAE0i+SAmGkocEv6+V
COT5nllQXdwq6vbP0Sf9nSjO/6Cd4SN7qEh6zofitqex6ht22vssZczQHn3ttehG2BCSC+wYsUqt
LxIuLulWMNlAbfFBZXPb8B6IvES8XRDCH24AqWCphKDWNWSrSXMYWtWA1dbWa8HwJlslZUU75wto
G6wEs6hdWNE9QggjxGhI3wOmCWIXZ9gLoI36aTUQsITg7nS2iZDQXaSjwwi/bkroP2jAEgkfNbin
lXP7QeV3heKbMtYCdarmSyDE+8hYOA5rAUYXH2olmsfYu16r4q28KPxqq6S4EqBdW0jR1a+5CvSc
b+MayH25ZNqmcZ0L5OkWU76n7Av/eCH1OdvZeibogU1+gsu67ustAsQz4POCc1gKy8IxA0/CyEfL
pvvNfeUQu4m0fwhs9KymjFAm4r1IfY9mgxjQpr8s7VBKHqhHJs4Eayz7BU3H9MbPgfLKfEbZRBeu
Yx8zXkr+8j/CMQFaQN2TMlpOWmAktbRPUHAPSIc00Dh6JwRCPR2YixGcZi5nEK+fkZdsgYoiroqr
A9N6yblJXmTWN5bJsW0DAuyWJ7ci4c3VO5BxdF4iLWR5+MNkC8+m3TPYkRtBolWhwEGo16iEFPS/
SvgpzdcdyUjArBWkbKtvYfKKbB2TTj4TyJ4wRtNpumTjmKyUSp+Bo9svjSDurTIgKheaNXJXtgwf
f7/4olR/7msW+Rm21WN7Btk+QqK2lbjVKlg8tlMQwhPzX70mufD+Oe+6kbVG50ZpootKzNLeij3/
ayp6x1n/YE+4HW08vK0fMnL36ZOP+50/ymUF+KV74JktsGC4JEegKy9xO3qnwXrqc+DIV7/lWwZN
8HqLUk3NYyQDAOFWbFt2ltT5NYjYtG3kLzFC/6ApjmqtO4gKLE6MU+UW717qKnDbzKHTr5sbKb99
G51BZlIpC/6ws1GZw8OLeZDDjUjk/q3tYgr9hdjW4Xbw4m3iUzmlKDwI571qzCsBcqKwqNaMrFoO
2BmgIOA4zUC8yWI4IgCA22PQd4KucldDEEylZs/elijxhoibXZSuZBp4JOBCq67JGC0VRS8irhWa
1R8kxzuDpc9J7poixq8NgPOpRKP61pX5cAy1e0YhCEw1IUSV+TCmx3s27qjlt/kLvOPD8t0szS6Y
PXE3TwqjqhgCeajPMnzfAlK4pHri9dKY2E3qX0fSc9FvUOj9CaxrGJKUesWNosZML47sCGVKCFYX
naPS/s14jVBVR0Rl6sRDQpQlzBMaClOV/jz3cap2GrBr+v3B2KO1Vww65DGmuJMsuyoPgVvTjnQe
yvarqql7YuNWgRbIpZWl+jbSiukMMC1KPaJsEFbfAg3aqPmjxSKClPiZDJZaalfxugyR355x1/5c
uCfXFXbxg14cip4xyKKM2hmCI69f0aPVJAr/S6n+dIZTkzWjZWm76xjxpLxqx3jM769CkzZfSCOb
9OXV1ya2PO4StPUxmrZu0i8YA7AuYcGuYhWuCR5WOvq/Z2Bwqn8sES25+FBH2WbZTxz/hBpxBztW
FN5TuppCMOYZk0gG2Dw55W0r+tTlDeDa4rCwEoptUQ8637J8sJlM0rgX9hEsSX7L+P1FNWBprmDd
MFjrbVP4gCi3GoIxWOKk8O7WLcy32q6w5ZRPDlZauiEx9aPGN1n7Ip8WMNcvRdlAhSynqGGwfOUz
S8efaTfnyJr6XloOICVAH3YQtXS1mzqBxUomkir/sM6Ky1s/xf+B8dvsVYBbKUQzpthtjCaG40xR
ggSEjEmpkDWBkyCB/zD7L0hNHsfTY64yp5EOkbzkMB/7pUfPCjXfMaEzrq+cQMKQM2F7Ypqy+TIb
nquBj/JrbvrntQtam6nxHc7sZNeQh9AB5p3SQXZZuvocUQQ/G1jG6QBMpV7kEm/M8v17RGmJsf78
rS1SHnV/eSLWb0wsJRPlQ1O8TKFPkpZ9RNybOCLneKtAobgpBZiORZlaR1gbr8rEI5bmCumK3Kte
9C7jYJvJMWE/aPD/q+/TBE7sXsU5HwuDXSJxyEEQq+XiCx0xAKFSt0ApzW6i/OGbA9wwxguX86W0
kiUjiCSHKhcudcQOuIG98Qcw52GzkEAWHvmgsQVqzk/MjzLgkdwChWvXFYw4SvHsGcxt9YpINMfy
Un54mbRwj2SQeeCQoCJtDhuoc14vOfQwgp/xU/02jQcKiSh16Qg7dCxOKuiFE9Dd/osLI8cTfmZe
oTlVg6Q1Fo+tPueQU49u4Ic9xM/++c1hCbXl9WY7LQ8acDS7qoB9YQ3hhL5u40c7icQx6HY+OXhx
iRlFcnRd4BCepb+0K4s7lcwdnDe34Oeg+cJaMnfvt1O6vi4tRaPZLuEzo4N0lp4S6R7jRfercacq
ZH7yftL4oKHosKijW2flnWNtY919oebSc0+xM2e9pcCgsLsjp91A3V51Iqh6BeB+Aar9HWAb9jmG
zww/YDycVeFDvuupJ3zD6Oosyy2hGRXquaWWYo0Fi08XM7yROfah8i9evCOmW01Jm+6NAhUDXi2A
6e9+1JS3Z79924vBmTvEymU0AOR3mUsoXFsJoZoA5fiKOoGba55FDDetpEXGyglaSgLni4jL9oNt
Xvx+74d91YvAPRFfjvkp3SZxBmqShAREjhw+iPd+gNw2Yi0ex0EdgaWQi+LN37Fa/m8wVw6mSFMA
VRZoHbjRmQvdaS4uhlvyKnVPZpeEwkpn240v4nRvcq+s4KDT2ygKrqOZzjb0rUmCOLPEO8fk+c57
4PL9eZQLnpAtCaafc3pZw43lKCUKBo5KABiiywjWESg4fJmQCkjwVRssqrhwG8/lM8jjZC3Sqftg
T9rMeByg9rjUvbobbtQCOIneQgHajPI/bfINtLWjgqd3O18VqdSK+/VXfhpvgsxXiDj1DmNaDYfn
4smChUEfQPeZNiojH13Lc6iKN/8NbcHmwOJ9hdMiA6pTFep5zVMDRM4i2LoE/3nDfBAs3Mj9vxiv
1Jz1c20WS2W9ZTivfvW2PwRP2k6ZuEWgbkRSGLgmFvnWLnxUqKlM8luBcKzeNOtNoaHeQdHMuA9G
wcNU4+0yXyjuFh9SZpjjjGjTwYKD6lWE+qBE5v3LhA4RvDmqgN91TIQKKt+NdQEvye8clNoIMkVH
qBbr6m63p9fP0vnuYKmFxhmvBME9D9+ezFKsHA/fBqZ13abjq9Yz3nwD5Bft15IUfKUBnv/vVZTR
+uDo4QherUjImHXcVee50JFAIgf9+T1d4OnwHwshhPNxeShNxy8J8aK+b2OvgTy680Nkox9NLxGU
zJjJ32T8h7yGWa9bVywqSCkneK/YTUzO0xfhhYi3yFnxUz8xJefow3xkQxXSMiz0bxU1uQDcNovu
LrR8YK4HZPfUmHZTOs4oPM5FR9YcbY9dFw/LwcYNhOgEeOBXa7LpO5FQFf3hccTzPV+XeQmj2pQK
BbGtNUq/+nv6bKQ5mua4oevTDvqE5xpBvRsNNIqHbwU39bNNgdzBR70QkBCp0V093jDI+xALiFFV
kuF6mxeAPQP+n5iAY0CV3/Ebxo8WnRO0iYiPIF/A9oPB9pm2gi91FgFyn3UkZl+2TvJnVHMgdY9T
6pgEBFfzH4yi+CImB6c1bej5kNVJ9mw6/4PhnGW5A/C9vdAdOpvyiAkzsyU2srVu+r0XQ7o2M5JH
8SMdJJYswY5GmiNVF9PaGepsr6HiDi1uPRB30kv9IP9UDIqXnyQ/Am4tUBls3sS07QzqhR+REewU
H7y33PqttaqFNP2jIX7S6w3PkNiMjQjWLBdzV8EczlQaqJauOY6PwIdf3Ae/0d71YX/B1bGwZgPg
/Vx+M37Bc8r+eyvqejIKb7gi5bKog7FVnEfvGy49pT499Wmxf4sSfSi1rYbqC5hAWAn41VYLrw6f
ZX4dtgLLa4/tGZhFcEAZ+9crOZajAnvcLjk3e41MmqjNYf8ttZDntpMHt75ggFDNfj/7IGiIP9gH
ShOsv4q0b/y09Slq1nAZui68TJpxWVdYtQoRrtLZ7F+peKa12hBt3e8acKj4VM+T6EddEy/m8vlm
i8m2d0GLUv8jZ9gynjO71HRfsWYzMIoNomhEKJVHANpuKhNlXsIdUDlPNqbwYQV2EwW6Cy7bfiT+
xs4shiqLx95E/LGg02Pbn/Rce0YLtuQr2Hkf4l7mAvAY2Cm9mfIww4EbFPNGs3L8G+PG9WYMNkmO
W7OMwxstAeu7ge0RS85I/QsmV9QJcMYOWM5zHabonTeDdKtaw5ftd63CxmWGbU9/xR8nIqg9iEQL
hjsQ47Kf+7WtoFad9KljnsL41oySFpjBrgmVO22rEkkXVbDjTCsjMP+x72ghqmZbjDW0TkekxDwN
cgN/tOH6Ua8GbGrfxPpLCK4ovA6N7GGq5k8Rjp9ujADTTr0kLdaxKbDPdbix/0BXJILWEJGWnqEX
0KIlAePLbhkLmYZ5pgEZi9lS9o0PETeOiDpMlGJsj29aTTgspjBNIBtlJA8VvVmxRhbLatatNTWx
+JytgWE8rE27yNHAybrJsx2TvpNZ900h6OsqOvaa4BXpDbWgSLYIllr050LKW0+cxznGbbogPI7g
9DZ7jL0JDf8usYSYcYGcnMmh16RDpBj/04ArxJbX+r0Pd+MeYttSwTeqZZpHdS1l3ujAjo8qWJ7C
XVA8RZQdUgZqmrdTX522Y8XIYUGtN4Iz1aXVld8VvwtHknYXP6iIS3Oe0i2WQoHi1Eg44gfnRolK
Nh2DjRBWIBZw+PL7Mcx9IIfAyk72UzI3Aoce5INXz+HoAPN7Vi6qjIhHoXTVlOpcUUKcT2VLHtI/
pkcII6Fa9iO0IzPshOQJH6kxAPougrv6F75h2aeKWNcnYfBMZ16/6HRGe8bin5syElO5Kiz4RA1R
sJYtORt3fLrVH68s6nvboT/UkYIiK7P+I/5/TOVOH/ldf1ydfwmEGizJKcmaaMEcoG1v4c6gjhkD
EjvYFtoaCkeTjdvZwxW08e5Ln48T2BSpsSrbhW3BM4R/Z3PQGzBGRNIFIDlkt913P/qbXOIPGiVe
pQSeKlZjX2aadr7ObZ2S0R0jvdcAO7nA8Fb4GGunlYEODfo7Rc+MubW/6ediF9M99M362zIoRwG3
eAiHe3d9ARQ/gonEHil/qVhaJa4KD++mONNa0p7hJTRf0SCv7ZnEXNizIzvy+4DiF0wH6xLE7Q2u
NNH12GX/us/5+stK99XBLXtbFoxCUneG+jcG7q5GXJ+7b8rztsaTvU/zI3/04uvGQEglPLpZ23Vh
75Wj3VqVIROlc/9xLoLS+oswf01TUdcdBKF8sA0ZahTJPz/pI0DNcpWJc/s7w3NnNVWQ/YjY9uVC
7qHpis53BRcS9D4pB4j1NyoyFU2GniuNMgZ+rp5kg8e60f6X7no1lUWc1kyk6AF5NyqLdCrNMgP7
LO8pxqKy/KX9q9tUOTEo9THesc8EbO6mub/lF4Ix62q5dTCoGTCR6rWvNP0hy68Ri2VKQ/LvCa60
okCT0Mg/GTPv1pQIM21Kecr264bvvY2A0X8sCjysbN0OPvCUg0e6BxVMNSQ1UU+vkEs/VdikCqh9
QRRGDUlwC/cDkeqTGFYskyUDrnM8wQLjkrIJnLvBEI2e89mNmss3ovc12elx8ncT5oKCoKqlK8qW
12yCztSyqlW3J+RwEsxh30oEeD0BAhBiD2mJF4AtKBOj5NR0DjkvSI0UImEJ8lxNQGJuLIfixScY
opq9fhN58bIwE0YGAYHW5Kg0wQySln3pc1dDdgb2w7GpogkziLWUxEx0WRCik1xGHVIPH5KKl4vX
suLv082kp2snxlmfXT9cK6kOo5aVaV0a0SkT+iPAqSxxFCmRqhY0jB8nsjYxw1cgA2OuJUCl8g/5
uQariOiuT0srnRpm6T9GvNccXQuSjmK6Qnyt2lDaM7BBzevR5sgjsp2d8Ex9579/7HnMsw9wmmdu
slP468BxKIj3k4wImj5fPcyaYrcQslKJk34ivvRqq1ewJlcDFLRhYPIm0vXIv+Nqjs17H/U57vJV
pJa9tUL8/SgQFLeqROslmHo8Hv9GmoD8d7oVo7Nyx7Eo6lLJDd22mEb8X4egfRr9cdNq8AthIKsZ
rggxIBmRp2T3dXrrvpXGDF9NDBLtCFh9Z2ZVxDzfhARK74VAIK7aylmfckQHQPh6Q23RzsgRapQP
XGT6+qvPZrqGfSuDPuSjZKHf8nl3i+GbV9rVsftJRKJxgPt15tO4QvSheiKq9UUOycF5ocnMPXyA
r7nUkIFBs7Xc//3r7XCVoksKI9CC4xD+faN4gCUpE2cgj3EwKj4jri/pnl1hOkAcLA69aN4EZSY9
PHL8P9rGs8SLM7EB0LOJb+iw+mkuMVxcBKVBf1OGxOCYCVtas52iNupSOWnVJwi/wsl9/yxJP+vk
j/rkAfeUTfldYBjoJ3kPR6XapIBf9fo/CpjCistYpFAS37TOTwx+0SC5TYrB/1YiYJyVBmd2DPrf
I3QU45SylfhjnTHr3GODUgVgzDr3YIMQYDTR82/x06CNjiFVMVgfH/PSuzCkXMkACce+t+qrhnla
VeW3ZbAUCBumyuB8fGpJ4mw6pbirLWoAXaE3CGtKYiLZh/aRzCjJGYwzbMnq+LihOVBKu1eL2GaP
69HgM6+/i+RpKn1advHl54SLao1tOdK1pWodNnVhQM9u/P8yc+T4Ua4t6+kYDEzlxo9nTHvYLkRP
kQNFyhM8GeiNF/2EKXyPbnvmF2rlrTTNdhWNfq7PZvQl87w5Nm1k+UxBB/37DH1GVbl9Ijsz+LPs
H6f4WM0aycZSYFJq2i9aX0/GiYbMJ3tQlTu64391fY7+lKnukWqAog498YrNhu1AxgGPslk0TxOE
4JbWLJpWTTcsj2NU+FEU2rlV3kehxkGZL7gijatipQlJJt65/eX3GnF6o1sTsvueMHSqILoQ68Ul
XvP33rnXuiMx4FagMyRr8e1jdmBxQHv3p6ntsZ4eimTQ/48wEX3ACK/S0cNyzBK+RCLs+TAJKJud
VXP9BZIgZRbg/gBGpsMDIo2VHk07NZ6kK35MGYZoSjH98JS9WpswNZSWQHZPYBJzCFMWwNBscy1x
M+dnvC9O0oA+0RXAkptSn8q6JazZd/emBU3uSUTX0sOOW1WWIEC730k4IAoXNryrDPgg0RLwq+4r
OvFbgjAxEHv2SQ9PZf0oaxcGHbqC1lINj41bA8C8MMELFp+rVrBw+ZWCMQGPLBaSK+elRnrbN0h2
8CJ2JvYs8jzgrdBRZlvQDV6f6VS+Mnc65JYZgCgJekY68y1E24Hlr2e9iEL0qJe5Kbw6lDjAytiI
m8vBYLPlrTgsLX78lNqS9JWwI8xmMbmmqt1RlAnl2vf/c2ErDx7syZIJLhO7eT7uSRMfL9abyRQ5
r7SDa3wAnW6m7L0LeEcRBEuMuMb3gTGlETZamVjz6lCLpEMaIWMD1Y6uM4GUFOkQ4EpRSX99epA6
eVHj11WeSeq0/a+ub7cUjE0454xZSHnOU59SQYA2oh1GGqXRSsP7YvGS2EoELP0wmLxLMhPNq8P+
ZvmlqTWsenpSBKD34yay+yNIgQYikvTcbEGGQ182QHE7csXIA2MLTARQZQoK6bGn/AQKNK3efyD+
kY8t+krIJt0I4Sg12P3oelP3NVjAfkMhDcQymilJEBxF9NAk9eqmxegdbWwvt8pkMSxuLm83FRlZ
oQnI/479cUBSG619Dog6R2H9URcG/38UJY8W4WSalCuzsKkF7y5UhsbshwD1CJ+vFsr3dw6uAt62
3UQCjj32tN1r2G4UpqWpaZdtxV805+T0GHkEMNSpCW5ROGUlMaUEAeLmNG0lmEFbLaxtqtOSwrb+
957ZNmjprXHOjeYyN+y013eGJIpRW2wfxBZNIrWW80Xvxne9KGEJll/8MqnCCR0aJDLplHCLBHjQ
3pmiCSjsd18vX5jAcodK/qvHS9kZnDWMM2E5jeKz/t63ZQ1cJEm9JaUuZ5Ob7upY4vnF24MOxI4Z
L3UA1TgfJjclJ2uNEwnRyxtbU9Aysp4XgYGSG1xn34nqtExLztmmTiFRAjCfDRw882krSEW8plcn
nBLwwGcgN9hsKOQJXs7r7tohsh7NSlR12X6wCUBmdxqT5x7wL7x/FRt63rtKXXwD1rgC05pm3XF7
SQE5wf4WllKoaWWqCgz3wIOTn9kDNKlSrhpNkuHRpFa4OqOZkaIT+HDtBjqVPXDDVZLUHDDO28Y5
bh1QJF13k2dLBk5MXzEskHK3OXde/zVdNT7XLKCzckEyiiZ0qnHKlvkBlCatGMFv+3aQbh9NLX2m
DtSOUZbE+/FfUhhkanhyxG3wH44qoMDa0APrl9JF5HzdpVRR4XAq1jgCxcU8EmmvQhJqKH7Aig4v
VD/bW7VfZWdfwrqu11epboZGAQTM138Nfq7+oBwFO5QDh8p0x+BXLZ1QZSeSAobx+kJTS9D5hpbL
tFeKmfddDYQNUObCZASRg3/Spuu1pUCLBPvuBnRFA6vW5egBru5szeTMgDuoM5/8XbfWyFBaBlS5
Kw7KCKz2eM6W+/5k7CeCwGpjzEw72gpJQ/Zxp0gALXUFHhLPrj2C1X6TBveQs6ntgW7ixVfk6k3O
q1AzD3I915T24QwNBAAdOkYHeXPzES1hrj0uHoNoVDtEjErKcsF4bhvU0JIFb8fUo10FO/apcqHU
1AYuWcL8znAP1zyxBD9BRKJniNqeeDT9/5TEvXTMKHxyyv9E9gH7UKkUQR2+mKMHl+fVt2NtPHdk
Yl+8MqzkCc6qd0pBnGlu6GNoR0t0IUifQyRRhzejAdhAanG4mvg66FiB63CaSUWtT7eXAB5YYEcc
TwsaA37jwtXXYYe44wa1QSNEKrZPAz5ZYAFx1GyOjkYd7Z70dbrAMdcHqhhi5jsf+5DYSvp+7gge
ypxWg+epQiMMdwKuh6WiUTabmtMM2Er9u8TDifctzAQW3c1KCy1dEWHExIRSjzSKblAYM3LjNd7B
FJ7Lx/TBaXK0aQnDKG+LYWHA2W46za4rRKPSs4i+W9EjgCeu1+vWWwWNlhRaHnjVhCT0GPCMitVE
SxnQaS3KWmKCmTkXWgpHEwCWiwBtcbWX5XoMZ3J7zqiIsIRObflIXn0EHXY0bIfW4kNWyk1rP2nk
oDJluF74Ieme3WWTyLu5Kpd46Q37mkeQQCf2o8d0QrdywDI0jk2Y2j7PWHoLpB+ovLVbVyJri58A
7MlthEXQvh+UFavBkapDagu71RBhhGgTd963V1O6E018mfHcqbLwPAygMiyh98d02+F4jiBvVUA6
7Y5dRsUbmF2hiL9QYKxMO2w92H1jFS/vWnNmanHa4OxGflu4YZsBCdfcb5ZTZaf3Mbaw3vu8ZP4x
+PjyX0nafvR93zICpznImNtOf0Tp1zphWAj3g0uNSMKVNnEubTTzmrmtVPa8myL52+iS5Wg0jKbQ
ZCuCIVhGkVpZQ5K5wdN5xYd0CY7w5yTBh1jBqBD6ro81EGJSpF2eJ4jhNaOCvDeQCsl0A3cYwCh1
bgV6YoHUpQQzBPFl+2s0/TaaWbK6M54ZF7o+rvpo6EJNBkrLvkXOLiePT+rgSG4IgZvSQH76x6Eu
mSyXTjw7czi+5BFk2GWQjJ6UVIxrWS4Tby20UByHqnSPUiZvrnch17/OOZLObg+FMnUkb29eqLFm
lXLNhXviEZGii7t+DXSlgl4Tfg0oFcuj6gUJy4+V+asCKnBwZ5TdaDNVlx65pjGma1YzhJwnPpaZ
fEnbTAP/VbPHk6M9awn4WEDjz/5mpKmTOP+ByXAxRKHl18KMfFAHIvEQ5pbkGsJLU4w47NryLhLJ
PBDmBNCfoGZOBBc/KiMQQnSBnyaeW3tf/RMt2Naw6ftIvh/G2D0dJ3kzza9KLJ5plSK+N/mdnrHd
YJXEaCllCat0jrvTHUgWVlyX+JmLYUB9/3Z+toSD6rgIXygv271DmVHaQuy2KloEsfbkY0kU8uMN
OL+px2ysyeMdnvqXFrSJKaGBK40lvX6T4D7Ru6T2+8d8jDIf/WsJaBNk7LV10BNx07yVaTrjWxVR
To0+kbymeHsW15MMHhzDdF/4ge9XvScHIbNhw4KZMTzJ+d9CcurFwR0Un+pCmRFushQoKxmtwnvr
lcH+MC4l7BEowyh69VQwAr6FVa+ADyWPSZ13QLo7Yq0cB/ZOUrXzKeQQGF8ZRmC4gra9kNjiHSPk
CU+Ulmo3SNyWgdmJDosn3ArM9LKXPG+a7XQ2V4sSWlZywd19kFKgQeyt9rkttnGiPSN/H7FFPAvG
n29JVjNePOdeI/Ek5FIvHl5yS4JhNzMhADdgygWh47gLhKrZc46hd6eETqZlXid8MetyNdxMZ9c1
966wcqNSkEug2XdDPrtje3/S6w4k3v3YEZv939wwcqVjwhkHTaHZ93u6vzE/EnusR3/x+DpYBLMm
L324NtrmZY7WeUZnigMX7f0AYHyfhU88fgZa1Xiw5AST5HwS/KlVPYbS/l7LEbDbRS89aNo9muaE
IheHrMaItc/1WPokShNg3SNR8r++L7Epym2gf3p4ob93ieAmh4uoDX6uLUAZ6wvrCEr2If5Lxj3u
7mWOdECqcw+g2VKYScsAYGajgBX2oSaVCcQz8Xi7n6tOvVSh/6iwD1txtzi+YNOMU5vaFftgBqmv
XIs9J//4+yj1J7cdMN9aKWzUIH0yiN+zbDQ5Dp67scWm8+tEyFlpxcFBgGAwaId13WKlVu4CxqD/
KHQk0eHlDn3/ScMcr3aT80FMHTEXquXg02QBxXg9mg114KOCh81vKdD+h+uyxtoL0HfKrTK0mxKz
WWtwGzDxa0nZ51hGPKJxUYU+r2KcBwCYhgVNGlkbPo7dIMsEJE67ZO1K5CUSrOLQ+9rYGrB6Vonj
z+IPo1KXOcsogf1Gz111j/QZLVoZ7TkDcwC0I+uv0RSlohm6APCNyOMOgy40t2EuvgfTJrARWVSv
MvI4VpI5yqLKb4I+H6dllhrm6M/pJ3680we4AfNdkpMRRC/DRcmmDzfv4fJN6VFEn5wy3coGjo05
3F5wNpx2la2yFBOQNnQPyrsgdnR/3SiyFQS5gy4qHXBbze1W/QV6JVxhZb/2FcJGoEStNGWUogJP
Q0uigyK4voNbF7oc59l3wIOeA8qEPC2en3oExy+2oc+FBD6hYjHSr5oQrXV88hG3h2f+GEl+Mp9I
dOyQf+pr7KQZFr7m0bp6ZXamb+nxlRiWTR6qoklZujzzS7HT83QJsY82/L1fQW91jC7g7LQKu7M/
k7CfX+fWtrvPC2tBkWguNW06W44QEXTbIq9QA6ZTI2DLRULQRSRNgDCJQUFgZZPqKKXhLB7/Qejj
aro3Xa7u7fqQavOW72CdQ0nb+17CseaLbCe8Zhz/uq5CClT8ZNNgHS9V/JtVZ8bbctqhDThcnlKw
x/+DrtVscev3+qXOwVHBuwFbRIM0p1cgyBZJRZXalvIme5b0IRzdnHMI3Oa1AkRZPqBydw9PCCUS
WN6H7AkmV8jdFZAaUu5Arwnexri5B4yrp5uGFs01+5fcFm7x5BKnmurTHeeZlAIe/Mi8PEOVE8wN
wLxOyzr0tC/RJSV5+dgw0MW5IVySEQ98pTz7lHO/3Uf9UyYWwgP6qMvQdmbSggdI7Iz32/NsBMWy
OJR2dOAOtGLweQd8oI+/htmD6J/gk6SvPVqs9etEB9zb/fNfxvS5DFHyHCxsmIV3sJgtdMUyig5s
EXKlW4Ol8O/W29r0d4CB4p94+Nl5yL855EZNalak8fXgKg5N/7IwIDbxmXCbFL6a9FPv58SUQKJx
LORhuIPJNFhXqE5hkQtJTejHty0fyHolI8hOAa1shIhrKIOijLlEIMJdpTNY6fpvCGzj6emHAJBv
8+38ZlQ1wm2AOP9oB3rC2gB6KtrzZoGredJifyMD+tAYYeigEabrY5WPv4Xhf6D74ArlGCEe/5a6
93PLLYkRWr/NcPbW6xTEkWsvVAVLkprjy/+7em3eDziJCgPWIe5wjKrAju76UaqRP0NfQmV4ReGZ
68kH8oke28OH/OXQ38qMB+r0QKWuAChBr8jqBsLUOXO1hKrSCe1I9C7X6BebC98d7ci5z+aedZ4j
G4cb2jxGAZifyI8/gp4Cx3lFm5GEkQPJNYJ0iEl9+BD2OhaI9JTFY5jjnSCy1Jp/+DPMioMCda/Z
Qw2JWIIiZ6L11txTeA7ZrV0YMBLSxBwO12ZUH+ReCsMWuluAoS6sEoyVSgk4JXSoCHDF7fTzv9eC
Ptrdr5KWRP7mBvkV9vRbgfxEI9QyIWdYZ20xqoKaX4h2Kz7Ji9CxCv8z0n+HygvumsaOPKFdMF6G
ywBxrf8C9o5Hf+hWPDFN+oUy4RgbmtITl+e3h7A5fTAE6Sq/XCD6XHUrPq4VYPaPVilvwMShJBPs
Co0Dxqi3VoTfNx9IM4mwdtzQWILYrQSrNNee9kGLg49CyrWUYtS6zPffSLTpIAxcwl1hIUfdz90O
6dO8IXjUSRV0pF6GBHaXCQm0arnj6UBwLmWgz1aqfHBMMOX7SRmnuOvB3qX+oiGkerkLOSSGIlHG
sSQx1cHfzQKeU+FG5jr3Bpw9h11N8ja9jxw/BlCCmk6m/pvZzDzE7fEQQ4cSQrF65QgHtCNOZGfF
juMnSi+yIPjR2M4LCsISwegu8t8lwNTLTI11DHs6Jjd7iJjgFUyJUreTTdtGLKuP1NdJPDxn64GP
6jsli2/llQCoRKCg31xv6hq+GCJhfdpUb4O/9dFT/kHj749+wAnfTsc5VeKkdrwh1lSEqptlamLI
B7NcS6yqfXkI1KSKXDBu5lK7yjEaAIQukFZZ4MQDbS+SkUNXRow8Xj63NvOdrG2QA2KFaY9pWd92
kT2R8DiDLOFnnYfN72G/UtAOlg6JBXfxrU/p+pgRpxbWctx5XAPqhQusYqcyAP/Ae14wEXmMV2mS
ALgxUZ/s5U1eKhUkJgAl45sbJ3+qUHpCqIn7kkc57/aAsJ27HaBCKQHVKWoE10VIdieSV+tcZnMQ
OMIXSq+NYzfck2d8051CG2OouShYvBPAV0PO+CWIBirUkqfSls3+zjWVdSDZCTQp5/iSq2c+MoGv
iMncPETIeu2pNjSC73nPh4hyIsftMWoA6fzkePM48sKeGsUyfM8oEnnbuACwb0X1vZTa3JA0MHvJ
MsBkgK+iN0npZwckt8m64pxtPN8Vz7UOCsL2AwynPinhbwsWyxk0xFLRuxPKe0Z2GzmYtb++jANf
CP3+KOIOQ3ZhqM+ove2RsJQZaFTMpgTGDngQPA7WSrLCRrzHSJAZp9z+sR9WbsJvsCSCVmG1zEKc
Wku/IdSM8pqqIJCoaKW9WoAsF2PqX0t1EsswkdI4yyZUqq5IcyIc4Yj3oVz7+PYJN95tlEYnGRF1
50+bHWMF5I+5yBjrg8DNeAjHYZzlqUoFnupU+ncoJbizql9o0W30B4UuWNEPxk/qKMmAeEdqgqst
CnS26U69vwqUb6T+YjtKaRB0DZQGZ1+O7puT1MbRtZWrsn6QmI1wsYC83wGOYNRaXmxPfj+qZAeR
fiuC1fRbFqVuaY9J3lm/8awr3/IBm1s2z3WtBKk3XHUqLtiIG3xycZbX3XB9v0rEZ0Xo/HLGnaas
IIoP+Nhm8cmkEh69PNgNTcu46lZmnzkdB1XnnpddqzQSxiqhnVhOPUx/kWc1OdTEMxMaWmKEMWh0
tzqiYoFNqNnfP4m9AYEsUklyqKXEPJI52D/wEuYY+GVmUVGv7n9L2O3mELnTY5WPJNoesDmFHpmE
oj/XbeTc7sH+tzKnjmGXJb8JIFnBAXJym/hqaS9xvBRIBfx1mVPlT83norVa3i3SbBtWbio1lYhW
C7/0uEA7L2LA7EQR9kPU6A4gfuGp+o7zK9Ti3v38e57i0y9jjXSGpuIV9KSiRV6JnFDYxijkXQ6R
8ECklcnCs8EuagHQl9iXV5+so6pQ4/U7mYfeCVDRtmNxBBbjcImLvURCMF/Rb4sbOxDRqFsGdjuD
TB+XYroIQu+FnejEgjiW8dMcSyMM24QdH5U7EBKh6Jiat93dXyHXVPCCMAc5WOUZ5RIplUh/L4fC
kE1fgdLMv4RKd8NCjgIK9DSsY6lWBzuIGv3Z6QPQWTWXzuAYBcqLPdHIO1WluVvfonxk/q5U56A2
IMU79VSwMQLjpBFB5IBrlsViwHIoNwUMTQQNnT0ZFM/LUOqirDL5GWVsp4FEGip+wzmL9Caz+Ukg
HyYK9PjDWE8aYSJUm49dLkuCxpo2nIxaED2Q5T6/7e1QKl3bEFJUTRtCAUaQ/nc7vQWkQ7A6fxO+
Q+W+VlOzpRpyhIr03So3kCMLwuaCyWhLYHuGYHmJrUZgo/fqM5DlSeSSaxzlvxiy5Qc84AnA5TYm
fLiqVNQyg0W69/fFugxRDpsny3HpL3kfsCeQ/0JWh4oPdYhWU5H/vjLu33pClm6M1tE+LW2vQY9g
72J1jXri6hGT7LLli7bI0QSAm4NuEoKhcdCZAg1qy37/c6FPJXU1NQaNClufOqwtNhOHfE7mISZw
U3LC4hIQ83B5EVTuHgQmTmmsfxOIrMlD4bxPd1oZrbALuDpYKNXlAp1RNFk3erAy3XkawBB7aoGL
XwEkUH806b8+dVUCn2yaG/P+p9t2g9cmP+DKLWJluskY22tzyGPtKreG39GDOj4AgBUcOWJl2jY/
ntz33gGjHYD6heFgWZfTDS64OwfkQn6tECgo6nRKH0KrsCKKB9N6vz2Nw29pR//LT8dKH40lmn7s
JTaQfePwxZbgQ6E55/Vrb37dnH/KLoh1QIQxGlvJIYYbPZ29ikVjJUzhNsTBkZi0evg1FOQAccyK
Au9sVxQVHiINcHYmM/pBqsNRgmDtTsp3he9eBlzZhXRktwEJRDHqCMQqXb1DywbTaXhDMWVfKpPH
LTdxkVw75yzB9wfDxXvLhk2OeNVUrLvZ/8r6csRnoz5B59JEi81aEbpjoirp0eOnW+PUukPvslrn
lHM99fNMXPHPgN0EIlWNy1BJPicOCgcWSsZ4m+qFM2/hZ8E3+VPDIbniWjCd0yEYtbeuvWGu4Wlj
JW4NjuCXGQguZJRG6VpwsqJfBv/guV4DD2YW+ljiHWcd3CuBAWxcQzsCLAjHp1cxP47dkqgBWQ/R
EhP5VGSbJvbQJV1/++eiaKxqTXEKSqjqSOQWLagHEvpRSpZCyTQH2g0dFkvLVlLAc0PDYZPa0pTJ
Hn7s6Hxor4sxiozpY8i8/rMNUpZllGBINnn14Jw5E5SRFSJz8XFHpLPpHM1agPNSHAa7v3rCIeRw
9UEwl9NjsLIx77EgyyRWFZNfgFF+ux/1Y5BcypQcHJLxeJwwkR0v6rhTqSzc6OQzM514GikUGxF6
lzDnn+68qncT0jkj6vkU6eW8lDz5qazuK8vMMKASgYXpo0nhxjWrClHBKOjIJyEMGsQ4UeppcasM
p5A3WwfuYs7cHikmih8AiTxuBjU33uN0rAUgmBEqCswqWT8oV+gwOPf6DPjjSQ+/VqzqGNv9c3GF
w90HkXnP1Pusaqge3EcEdpQ+ZbxaCnPUptWR8gapYvHz350xmYgggP1V7/Bv0uztxJBnV5gxtPfG
ejQyN+nNAxlv2taadq3yq6OQtzEXDRNvFo6COfiZzG6Ms6cUy+VTx1XI8IEMyixsWvdtwLZsmR/J
EfwTZt4+Mty2engQDeiwfFKjF5MFdK8BfWCQcZrIc5mx/Gnd+puNMKz31f4Ilv1CYCAsJEoV6Z0g
o6We2MprAxYcELSKpNWtmslJbCEU7R9U0lQcxSH7rlZNDd4KvjxsyuMpnxbbhRYROgHOGcKFG7nC
id2JH1lDTdDs1ZWYydy8jBlE2f3/bpypox3ku0xlgaT9TckXkBiNXpQdQeIsQAizQamm1xfu1ivM
wTfz6pVX5Nw5P7z3707Tk7I9MXYGY294E8A25MZQ6hRXa1geSQ13WsXVfykTSDCCOajJfBjzbeXI
+j1M5i3JLdiQ/RRLqnr8VKfNKFj136rkGq436uJi2Bs9eUY6j3NW6KMu8btnZ9zxrT8u3P9BX7vR
wJ1i3LC7OSYFpkTZ7Q6RSUY0c6KLb1vF+bi9CopjEmQVo1v1vRcZrWHXjZ8ITt0zAHFfAirLKVYS
H/Kjw+82cNWXecoVAlk95cMQBXdSn6kOhSY0Pgq2t1XQGe63BB9PxtuT41sVQ7VxAea68JHupAtc
pe5PDZ7xPafSE9y69+LtPBgUmov+wjefmazio7KHDQcMaDz+5FiNstdLLmWISmGeubseXZfMLssl
Ok9GRj9sFL+6uOFJJnzz8bum0ESdxHJp+Lspb8zHhdz6WwZHscx6Jlg8sLfd/KK8ECfMc8EmBfox
LJzlxplgUkzP/pmwL4NGUUgPGAsL7MhMHYda4br9c5/Chd6btjpSMfhLRhMFTrBxQmeOb8u7wIcu
061fWXV6d5MiBX4XvtYBhNVZx61vB8GR/QYJ0lLMsEB+0nnUWayE59EAWqAMd3A8N24lxhTu/MEn
ghEXHCBo02LWUN+NvME0J0D7t5aIibkBl7jOCXBrgtm06LxbD5Ow8Bw+XsDmj7HQFDbzfSgK4hIU
oA/ECvTUm5m6WMfEReUKyKybk3+17Xpbx0U6HMawInWMDcIPpBYxUtmg/RdZhL9MjizERJTbUYUd
vb/PrOgCYEMnaa7zjMuRXEXIupMqyCK2MIfFn2O75w/xd/Glo9X4D5x3/v0jBUsjUd6w8ZQSteZl
eAObMiELnYW7pqRg5QM/n2XtfQ7KY8qg+hUXrf14QQJTS1cMRxyTaVCfQXTXNBPjH5oyUVYPCQ61
2lSpdGtJ//HNdz/442+B1MVQ4BV3Y88D43KUgoa1MFrPeNi+Ms7HNsdk3gzuHCgyy0cw559F9Ue/
BCS2F8cY6TJeLOgOuugabDVyik2p3cURnLIRlpctWfgmTLsHozQDsw5lbIjDn00VFkWGntK/aNFZ
z44C7KdItOPj/SlhmqZdFCTddQriu1kt1q1i4ASY9UNdXiQjiqy2HZuWrici6/oT9SyT5U2bBlwx
9WdUei6DIXaeWm9a1DQlFW0+K4Uvo2aNwxPTSuupf+iME74EKen4AV3vehcTW5kYu2XSoGB++WsC
nPgYBf5OsHtWqegOerxEwjGlcmQinWK1RH6i9+Ls9CizVEmm8XJ+ebH1ekK390yylshQ+3OtozNL
RiUBlnAmHFr2pePjvI0C7c2KKxo6Hwkn+xMbRIrCXdPbBZZrz6KXJ/8tKV3LJu4Wp4rRWJxSnBcS
boCr9124nCfKyIfWlkdSphQKfeqG2mmBU/MRMhoyUB3LtzrtymzD342AFg5iz2nzVyn5FGt5qqFb
5QIj04Ug857yQPYvJrUFRkIQlny5LMWRDt8YeDzhzg81D2ANVu+4xx2xKQZVY+tN4K8sl8/+/m/9
ZuITIolskpa9aLgIGVnpIMseevGVa/2LmbP9szlE7Wdsv+f+rWTmOH2TcjYADojjv6ZKk2iT8MJ1
bIdukZD62nPC3dWTfjxjTABonk0WkNq2rtvz1bWGzR2KAr83pe9Mwi/ete6VxIeLd/ZuejUwF0Jo
Ha5ab1hoIsq080n03tvDySFtQ2Ch5CUFVIG388R8ztbfpshgj3//Xj3e6Azu5NXbOXQYK+VL6RAR
TsT/MJcJHC4IF2AK/u+uM9DF59gKpjMk6Mti9S3VPiR+A5SwKSpFu3mccdYVSAHnsF/mMsFBsQoT
o1J0H9upUqJZvXPeJ9pmJtcSbvbjcaKH2/eAI8tYZSkwnGPnAOUMMiKRelp4ijqpd7eCpzjeUBhO
Lffd5Z3H7FNOQHbUxOff0leyic7Czw+sc2/Lv/qN0MQhyahEan/XRV8J1b/YY1stS8q/juC2gh35
hGk4e8s3OODFDnxMzkdlWNcmjkIIaUiUWItxaLYoHtm4v8TlX0CADhJfxQ4Dlr/yLTmkYhBN/O+f
hLa476FUV63dWew9dBh3PYw9GE/jRlW136hE4NnAkl8wmkBrx53sPT/zgVPrlVujMSlldrG7POzv
IKe2boC6+ql1ZzD0X2y+xL1Y/qYt9SVbuv3cFWY2WAQuXNrGr5w8eML2GCYUkE9lYfkyDokCxK+f
PO7FdLOhtdM5lvjyapPrSfPCR/D/9Oa0IYOqTTztk59hyRn7AdqJ+jl7X+Jg8u4D5nuS/FBBDHdG
pQ9PMKpSTh02C7Cr+payZPy9c5OEDc6mWcnxeNM1g/QNr+bgBdmSdC0eXUrvSUIIyzBcozHOkUKC
Uxf6NiS/Ql+5Bv2WKKLct57j0W5AAlKukAge7dAt2D+0928uuGtmGd310t/onQV5i9D3MZW6vjJz
8d2B0Sjh/TJyZxhlN/+yYkfKJV4zla9vrPI3MAeexM4Pm2RFQ49hidDK3kzv5nyL1tiemxi4hW3L
wmEyVCNKvs+S+ez6JsX6WJ9ih0QJu2VRCiKgeDICWCuXTRZqTJ4ktLDkNDu5FURoQQzr/Vm2gTmZ
qJl5xX8hicL+Pcb9OAJQuFb9aqjmuwEDYlg+qfZjNQ/KdpgcqlUvlqGXpcVpAeMDMyVJhRO7K65w
QRqhfvbWzqGHNIOALPJuVO3/Y8nd7vOIk3ow9Czz+K00kUVHy+6CIMDcZc0LHoUN822bTL5F6rmb
ZUDtN42p5XScUF6qFOAQPH0PPCL/JpajlwHXMRIF6hDNKh3R/V5+OlAqWigpq4ue9LoyNGtcoh4R
O3snL+1Ysxy38CRSw62ZgS2/iYY9YqCoPimXf3y1oWypR1rQT7p9lqG0xdoHpTb5KxsFv8MnM/TR
tskJDP3OOVdAFf+j3hM+d9xFMbKGjvuNHg7SuV7FbsCpjFXeiZNcWehFcnq8tAiqrzsQxY2070me
Ms4w8quq9kgQqur8BBaMts8hcr1Ogv6k/w3pXRMzGaPCidkWdTG23ZWVrxdmOda8fFcHokfuQc+z
2AIngTj6AtBn7f525MiXQ4k9ung1e4Ibp9IWACqrK69LQPVWkasTY3v/pAk7LdBaZoZxaxx2xe4V
CafKoZzDhRnMKnl/oQbEUTuesCnDV+q9O2HnUGf2OG+kyigi60rGhI+IobGuA/v30lDxZdzapaMQ
J+AcuaKE0+0da69G1vhi8G9tLUb69wlZFdZrAIUKvxS7qs4qrB7CbreyyCi+FQkq5Wdqersdo9Ba
FtUuu8RsLozWxUlREt9EbzFRM70bxAlhxvrE4qdy96BtRMtxF0ZsiVw4hCZLcHdEsn+MxQ4DZ2qK
tqx1gSVPRp2EpwvIRVWWUWxFpXJfj00i+xJ+VdDxXZEO1kG7ALTqJZEoVShaKYlermZeLFHQPbE4
urxvrR4pioRc8dYewywiRVp8Ph1KyF4Iqb4BAILloxU6FZRWoR04jTudtgx4p/+OSZen0rCIeA2S
cIVLiMX7ZXDECuaj3VWoNm+LK8FRbiPpEPKbK/ok546PO1Koh9ZkiXNeH25J1h0mdoUonFGZwAGf
SXVu0UiQihU/F1+v4dVyQXo0J2zWU8dXwQ8gU+lsmzRxkW1tldoPwhLD/U44+XITrLNBqsUO/ULw
GMTS0anzlTY491/fxZbSaShA1WlLy+nbpkt1P2jSMjnzF82B6XRIuO0gI4mzqcGb5eJbuNLpfGmR
Wquv2QYi3tVvEBNPvr6vYnDOL2Nllh4a/OZFsroNJCg53+Rthn9acWktjrZrfvay7eU+796Kgi6d
mFFLx/SVkjYFDOk3xRcAXhmb8RaX+ZlHX7gcogrUeBDXeQ1YSD8bviXlGVj48onL/X4fjCuWZagG
fK9vXSDGh3oKqO4knhsUyr0E4ZkuIAfnHw2rFFdmtdEu0Wbm7f5fnYZ1NabM0sPK0crIBr523iq+
kt4NFjOL9r6vgkoCjHqiptuk90FmbuQemEI0TTkwzphcUPL/1gFrgoa6Ie563JmqkMHTHY2Cqtp6
0SbfAwnYaF+NIYMBEEkdM9VO6Zq319bBqSnjUF5rNRb9iAnqdRCQTuxPklQ5FwpCSJtWqOnLOLhc
1QcQYeKy4OLwKM+2k4gjSot+ZGxCTomBY9WoT4pAJugz/IIGSK/CjTpN2K5V0OUR1BLdmOLOJlad
ij/CqnUG26w39MlF7RJNcQVcPoVlhoey502ra/lDHX219ZSJTyBbnTjLuFFObozEQpvMxqXrXOnP
my3xNNtCCMmszfCRl0hieUaSTuSrzK4QdGnjYwCaBkI2dWm+kXB9w4OwCdoeM//2ceSDJ6ywYIeX
wXtsmQ4Uhllev3/J1YRw6SmyT7heHBDWKeT2b5RAARCCQSVOObh5CLThi6sgx7mG84OerwcGYCKe
F0/WJECfEoYBJxkScvvBZcCdhuiHWCb8SjukamYnp3pIZ9SRRi2NCC/DjIPj+bF/tE29GfZFgKqp
2643qg5OYZBBusNyVt2EWkxObUBpWuEA4mrF59WHFWO2q3w6orcmvb+sEcYDCivM7h1WMz7LL8KR
YR20GQFqakq2ThLO9m78APAu5owR7F7eOnzhROVnHXpd1dJemx+NlKYzJ3XC2uwIYsJeT3oEIiWT
iNpBaGMTPrD+DcPA9C+T3rxBksxsEGYBPI9BUPNVfafQBrVu6B5fnBkKbTHciwqMRI/Bsroh5T6C
eAamvQUi/8HPq3np2ZWLdBHkJxts5xwMXBiP4ZdVKuSxNHmSMKZGd/XkryZTU0myKxyc4sInq7vA
wxBUqHG4XNrC/Ynp0uVgL6DAWpFJvAx0RH0NgFbwlEiSQctBc+S6vod9E/ea8sWSoVcRKZo1cBxD
cY/YPMb4KimLQGrVLrRCL8mflkFgb4fhyuPy/ocfFFSAsUc/IHw3oCrDwWtihLXoWqhGJ/6sDrbh
+igmhwocTqlFg6ye/17Zpnvwb1ZD092JgIT9G3HGUGvMPW2Lnh4sgeFcXCHaJucqVu+bZ1n00GTw
f8BXW2bXCBIgAMVOw2hdNswFdq/b56jXZimQU83P04W9483GVeQZM873pZ7C36DIwkaR63US+Jpf
+ubsaBs1DIxLlfvQKJQll9WyOjHxFcgmTCRTJggb/YVdZZ6Pj+YCmlxcsX96UB++8RZjwotIML7f
HQcgp7TYmZqTkqSWmiIAgtrfwEdgpi/pKXJiw89WNYLZpYcWTuv6fxiBdkjOFqVbwXxCXri7chUy
cJaZLGEaj6kR8HkJi7g43BeJ3zqrkrF9np7KF2NeydKYdj3kjNpVUvKrpIQ61UJH07wAgjqubZ/u
bPYnR5eFdlbuOQ9v6DWOKjdhyFLHRBZvG2Uv8ZUwEzD1SjuaWb7EmQ9qwzTQ9ZI/zaAB84+RZ5Pi
CDjn/nyLjsjmye711FoHFxYvJwudbVHi+H88rhnoe9DzezBGm2kTkQJIBff4quV6FAUBhPIgY4vZ
N7xOfQLRNT7jZX1U5HUo2+SeaYrvqEKE9s+/t2MFvKUgtp5IaoczGomt+HN3iPL+qMAsIXNPePEM
39c/P+pv0ga0icC9lt6XLfsXYfyfVG4Pf7plpu5Fcbmbt6etL4duABEJUzV0MZDbhIEHzUWXFJNu
vKkvon85NUE1CjyiA+Py+4K/O4Mb3m9TXKQH4XddLqrtZYo1Wulf9kIQIRnikNcFymYgwcUyZd0Y
2qiMtpL8HSinzDcqB3/5klAB+1J8FchZV+eWXcFZDGUlrVbeSfdQA6o0u1aoO5GT+qyvour+sHFP
rHjATlpjwM+E0skl3nDTTd2JdT6W/z88uUxah0ol8fL9g96jzFRvR2KdA15CnLVMkx1IrKjuAsrq
7mJFnEpBiHIDwxBXAX5yD8NN6tisBpW7bq+mIc8qaDNtYNBEmgsiPDEvPq3xkIGsIJhvGDc2L/hC
jLz1+uMpNFkG4JsfsyInUg0CKF9d0U1v+dgxP+HinfL3VEt9E7vlX1m08IojS3ivQzQmuKfoLqd9
H72Y7vOpD3NA8xQbRu6BrJzUowT0FTyxD/f/fCnSjo0KuD4v9LIx6GSOK1f3JNSuouhGPU6aUE6p
4qPdNoejd8SWrfsJcvB16pKuoQJpC7KI8VlrTvLwtTaJm8RMjo82JO5UnQ1HuNfg5MD0+3gZEvjv
mEaOTW+XtxWXCpzvBYQYC6Ayi7v2y3UPjKPjGWPhjqjsgtTcgzatyzNbsijSSEoqpH/LjSD4fEU0
TAzNcBMFiToJVPvYRrS5DGvTUAing/nAlmucnfDBwK8QnE4vXzMRhM9cBJvYohYKoYXYwXc9Vg2f
UL7tNJgF+wpeJNjWl1oAoBKwePD312HX7a34oDmaBVzTVSmkNdCAcLb8fXqANS1hIpjgWtdrBCOP
gygyL7FIvsqkdzYwsDQYcsN4Hr1bKSX7rl4pbWsipH5jD85YcEGKneeBtjFKc/3g7rMfQObgl1wB
YVtbXzLno6L+mE5RD76wtGCwIsgOd2vQ0Lx6GlQK6O7af2suQflhgwPfu/nHMU+rtP8cTkAHWfEr
/Kq1mM21Brc516bbU/aaQ4Vvk0hHMoq8AcgaSyhlOAo7DpeHTgbfu5tOploE6oL27E9ZPT2NgAxV
4L6m2ENTAqavR0D2ALRBlp3OyV99V6U21dfxJxk0mkyhvjGmqdChdp4JlFfkFE0K6sDR0WIOdKdU
mdRFvhWgUdRsNJVDA9ZfHp9NXjGPiHre3bfXzjIZrr8FdRqOofWpL9meYrkF1FIrt9PHNrrIx05d
g2HUw7/DmDczZ5DPCJVOhHO4JixF7mZCIJ4P9SEQnBVEx1H8HZu2DlZW6iDNk+ylzXVIJO04iXrV
vIIt0HzP47qg75bt8YsQaEzc4fGx98dqnmutr6Wa4elCagNkOgPVGB7y8ymoEIQwfi4qFwtdA/pz
9xItDK3TBDdcaSmdpDsPsY8x2BZlS/RdFJ3KkjeBr0R01u2Ok5mbGBDzbfANl4ljfdZHJIOfUrXc
efTIJmpKWHS3bTK+n/w5D8pCE1OTJ2r7Ez85fJjR2zRWqgNrDYX5QyHHwcKkeecJHljldtqk4BVu
cg/jjuN00GgIMmQPenv+m+PcwkofZqXQq5Jlhi9KVSmLeCg4i/hQ2r/6pZ4pJEX86O3u8a3+oJSo
wzeBwImR9ViSODDj3rO5cHvy0j7iVUM4PsfZWZy/QzyVqYBk7Dc4vyNlNAsp5SdF4n2oihYKrYM0
LhEpgJWXyeJI2EC6SBn/wrjPCaybhvj/HxbC0ZoKiiHO39dGxEzpAnnEfTmar7cVP/O9hOySZBJG
yzS452kARLa/P8PYMOJaySrIscj2cLAhyWCLDUrN6WS2aJuPrf9fQr7RKgDO5qeJNfqu0TQK1to1
otONADEobbsa+uwzGFTPicDB64f/2lPf0HxmIfVu163leqg/onfKUriyOfd83NaefyHKh+2DaZkP
d6AoLa9JpSyflSZ2ckf/KleZHnaX8fGnDuoFiysYApqo/ghg3rno0P6ePyRpP7D8Ne5FsTyiXfQ1
/B9mmRqQbvySDg3ggh1f849q/x0wqiKM6hEMIHh2w8Plb4p0wjws3w6Z19u+/uFRf/difcBgQZH7
PMtOGp54xqrd3V0azw5GPSZvk5/9qw0reEsSUCBD0W/3Qqt8H1M/GO7uIPLe8xObUAuqf2TpRhpp
qWmGfcnCYP0PNjEaR8610a3BpvQB6zo2v3D2UrbC+dULNJzG71PCXD/dnnl6stQp2jAS+YYo6GE6
mM2rVx2mhEL5pij/hSpejieQqtbTfozl5TPudi6nfAtR3zyurnG5b4v4zG1mKCCLYp/6P+DYsx1w
a56YooRMxN2DdUm0GYbveTcgZIJ92Um8dkDJ4sYdjHIy9Oswwzp4bdIE7pWSDB6w65aXNOjHCpvT
ZK9plxAUbXiBZQLZwAi6Ku31J792WfJcINCLxkjJ2eCm1bForCCgKEWWl9KqIu/3CfXJLjwEVe+3
RRO3pcDcy0ck42Hst8TVTGE7K59cGmk0GFnAB7AD++HKdmFE8jMrdDSyLBgy59jmOhsWk8alDVGE
x97bdaBtGzE5ccZ0X4iEXOoQ7JL+CuOBMwyXLIVAGMcbXYBhQxo7843lwN7zyiYBEMoWbD3WxAJ8
2t0uEPRyl87nHcF64+cxKC1tk36hJa+e+t6Uvz7219VrH1ROzhYbzP9BO88vAfE7o3e9J0ptlf1+
OBkQjXxNfSEF3EsdqLnFqzfEqauf0mM7YFDfxsM+MYfB197WuuRfvjj/IK2Exz28pzhTRskqX/lt
0eKFh+03ZHa9xHtL/SFBMgGnmLuZruUuI3cTF1J1uVi4VpkzUEdey4TNQiDykDr68zFoFm+stfd8
OB/A7Ibm0XS1laE99r/jNO9WeYyAp+dU1sTfkQ+y0hNIMO7FEYP4hjKRPFCndh+u5jVF1M//5Qsc
vrYk5MgiLV6tU+b5IuvbZPRE1cUB27FXSAdQGQWdbMXTXsgdJkzkPJYz+XTSSiDS7xHFWd9vRoiO
5LlA1PGnrCE0OGxHjzuZYSMkEDQkgtY5+YulJxFdh0hV6OoNv0uI3K8cXELIVRMEsjltaYlGJ3s2
fXOsAAg8TALNpWKA6hLIa+yobYEQ2GS5w+QXT3hNiEdSyxL5o42XmZDOy1M2WY4RJuWjrB3/ZzDH
eCPhzXM7BjGyIe4M7ubrOHjRMUSg+aQj7SPm4Kv60EzBSYyKayBzoNQimBtHzFUg++i8gAXHRVAY
CPNZPlD5DFpX6EICYveUKLdpkdDG2wdRz8ay1Q0C7hR5G7f0NywSwHj4KiPmYY7U+a5IbrO+QcYj
Aqm5x+6obrBSFhgyxPCWg3fh/LXbmnnecS79kX2VxI9SHdQFu1+nq0plQqVhArp84QGCa7Hc69Uy
NM+Kx/AunFlvCKTqj8zPLssHruSf6vi5nJMSZssWGl2UmMCwY6Yl5OnzKP1FtFWiBCrg0kiY/nXi
HAVLZbEh/ibmyQS/ws9DUdI3E6CDlgYhEIrTkyEfDpsnsWWpdGeCkwEEuPnWZHZsOyDCktLuXlrK
+K9re31k6BlfG8eqsG7Lbqkfg270y93NEx23rBAkKu9NIXejvw25ea7S4BbbnStG9DEvIINFk/Y6
GC95gjJxx9jjigD23UeirzT+k+qfdCulPZwJmD727XXGJnHZ88BVdwfk4QEGihgyTmrFUVaA5YJt
SLP0NB+CkRIaAFHLdw4OV9watQOWFA6Jqzs6wuWecpHdtdk8ZRROSfJ9aF2MNDEoCSXHcyxIVoLR
SBg9sEOrNHlGbkXhYxxXJSu9xAurz6AHDP1Bp89kyXjgGp7ltOAuNopCwMawd00kaXWjg+Os0z9u
6w/bJqFD2vPHHlk2VLd3Fda1THtXBsqZirS0UZBaR+LacAZerVfXOsT+Xuf61Z5mffWIQi0vKPWL
LJpubhacRhzte6jMljNzmnfOapEfataAOCRiyd471C0gNkHYR3qYMgu4E2E3zi40LRKkginvrQR+
IxYAx5HsY9QlNkdY6cXoi7F9JFOZvLcxDlZFdbJoegrNN9Gc5ep6QFSrvWTCNOYk6I52AuK6BRo0
LwRUs7qDrsHEI+wMeLCt0ArX7shCn+aarnd7f9qUd66Pm918vzajewXRqRtAGCK0Jez/F1dG9k/O
eIF71NJ0qbMO4+PxXEUfJKzlzxZUUxHAcyxgPjCKLe6KlaSLEeDNUHIAl9Ex4dmIX7yWdD3Pj6At
JBziWlNfnETH7WwjPct/dzEShnwgC+bKD0wjUkFIqMHCRQkBXL9d/+w80axZwe+VWao0UpyIVAh7
6Q5uSGKwm08cm/TIZsg0XUPSYL5xS1s0copoUzRMVu3pHs+f3tKaLTeWDLQCGJof1XY8LwtWq688
r80M4TL0ObH6VIeYsLFk+CKCI11kbFNuNcva8YoDCB5f20FCeTVsBzRCI3Vhgchkw9t7lH6gCXT0
+dj/g4lgVewf3xblINRBxw6WH9UkpmwMOxjZRlG79L/XiRs7UU3Fp2RrlZxJ2y5jCZ15M2Ehv5Wl
mzURrtfYcp7Lf/E1YiSm63Er8QQCgBSDyDf5FQdQt8Y5ZhrAOlvhaW0RnNWCzm+YYwNmS1aoI69V
Z+Hc+mOC7RoHxJS306W3Bd3BZdDfoA1fMbzyngpACNIYBBoUWkUvjxnBbYx7yC5ZtQk7FP029nsI
VOQfQBDrC7OoguWFs95OtAu15IjzCfzKe1q3SNTczDhDgKGxfaWdIvuGje3f3nFmJPzMPiEH9OEs
sw/Q/hKF5TRDr0rTEy5GS1tr7sZ05SJtneWBF/p9feidvqtJ3k36optO7lcXmXkGgj462R0nGJxy
f8Z8OgIgPJWCrMhZXqx40Qpk9FkHZG1k+jdLjIAT6328sQR7Vx81MvOC7ZnlpizP5GYH3mphXv8V
+5pJeQkK6Pi6aFC78ECKQy6+CpaI41S3gv/Yddad0UdJUxyRtl0JkXVET2aeb54xuP7/qU11Ruzg
skbf2ojJ/BTzYCeV+cieUZgZmCioa55nJrzlDLU0367u60X0lO+qEUpYPadTBoSYtolO5lBPf8yO
kAa4m6JQTrdqRNkh/CWy8qKPNMJnTcpFFWZe2LF5iKkY2DzMzqe5Inpr8zYIE2+fBaYh1gLiU9tS
IEDLKJGV4xpUvJGVEn8o8a6wiDTPn9KaAF1/zYjpTsRl9nNKoCwaA2GuzT8SV1+wbRj4QOtrQIoH
NrKjz3WAPEe1hyhjHYJ3nWQNmkjFPdPSM5u6aQlgTcLXkM6cbPeynccHFLilLgt9MpwpiGAfp32q
Hop/qzes0fd0Joclj5vDgjGq9p9kQBx3hV3vMPEHy7JD5+8WSHC++HDNxmb/4ptc+WwLOIvV0lKo
Fwsoej0UxxkoeytxnESpZ6sLRHx/0GtOLnQx4OKDMA5IeyKxZ7SKxp13yqHdVMgujx4TZhH6UVfi
EqsoZpZbdl3ZE7zON4DMsXcJagoyYvK+tDnqfgCaqeZqE2tLGmqdiCgj9MAS/8iUy2jfVWpbp//S
syoJl3RSWtXqnF0ShI+CKyIlLVben37/5tofDsvJ4JRKMlOOflXB0SMtwnzW7gMRPvNWTsKLK+iP
ZU+V7kZU+Cg5+D8NfIJVfuE4oc9WrG2xXPu3kTeTY8m3gspBKkmi2lU90AxYNjROUkWp2YY9Ny2S
fzjmexFjGvWA30yexB/sy5SrVHHSCf64xn56+pwmWXoX9MYLz3ogACL/yYeSmieir0NrZ6NHSjl+
Vqr1Lj9rOs3JkEw0x0o07sOYsQspBbRVeosrio8F21h/tFPjBCwWqyXJA8zP8TP8rkCK+Z3IiT7O
LDRsMfGUunK41XgH2eKFJ/wppTgnaMJozR3H8maOj1Xtq5Nvz43p/oTonvM+/lIy5iZqH5sdnQVs
DFU/j/e+aQ78ZhwNtLIA34E7dmiPAdsA77gtN9js5WZj9iCacWZjwxDuJdXlOTiYBZQt0b6Qb/VJ
+qZg8fe3LX+ztf2L7N6XzMuJQpkGst0Q3gEgvHThHkB5VOeeGVbOY/FjZ+KXpxAIQz9dvhdxTO7J
XrqBNdc5w3aL6v/fYDFCF1+bUIztiazJMWjaxvkmtnW2KpimxWdLHnF6kN9QFCVfgnGgXEdYs6I6
Pcddwj0DIC44kBsQMdyxDouH2X4q9eyLrZCn51kft25o25cDInuWFwEYYBXleomEd8ECzvn+mIao
XPlfxk01YzgoYOuh8GhAx8xbYJyTO06AoxCPcSvlLWXkeiHG+DaEobwM/cGDBk2uuTQSqVj477sG
SdmInjOOaR+jZC2vVI2iB4tkGTynjXhBH0lJlp3N2uCVxvDuNbP8xmlHP3PlmxeYFHEt0zDqfGKw
BjHXTbwBbsQtLgDlIVuG7gwfQs0mJnk3D7UQrq9460OlukODkua02kmsBVkGAQyYa4nKJK3lwPdN
FLKV0MkiyU6Gn3iPqqlDeIiP12lR7B1wnoYsKsIuHSg78YzLurdsyWEXkuQlaynyB6+d2RRq+G18
yET26wb1hSWniXG5R6OzGLBobDvSKDxX1KPhkD4sDYPrtjZK8kGq4OVF9HQqP23FXqPFjYSUAVMB
7owb+j0pK4DyXoZiKBhJhmS6IQHDdyIZ/HMweUjDPq1LteTXUuhWfN1ZFUMmqs29W6/3LHEEApuV
z+jHNX/RcW67eZxWVsjntnwqLYBMONpm7MoY9nxwrvQ7+qE5UKgC8a37VPbGS4ivdg9MFRT6ujTh
k6u7fQpz9qLgSzjJGlKUnTwLKhuG2ha6JyZWK1KZbfWSbyNNqbn2lcgux0HsmW9Op+z+G5G+8w8Z
SMYcWFVDgydi8YAxntIpHqXobAsUK9WXcXur05l1QhhxSyABMiAk+sjKSmoKdJISCN5ywYP+EeXt
R6hA8yAPxLJZ/ap0Rc2Plrp9ZwpagYhNlTsaxXRq7OJTFjtHaPivwVDvW2l+xOzhCbupGK61eOlg
4A7e77fNPpsbxnGNVMeNcCfmPe8YVObDRviymRfaWO+ya5bKMrMuqm/J3Lswce8jStOlv7kVHBUa
fCtPcbPjJJR1K7z8Pu/sXLLeE0BaUoo4VjRD+s8OTOeb0gTG8FhKEkR2XPLxb63c95Wp/2ZTqB+1
gJswUMvMbFf+BppV4YXk1bBZn3KkZ814laQV104nXngZm6kYFILkh4IkBHtlUkAvH9CAKxOxtZOE
7nOW/N74XBmY3sbXflelljTg39STL36GcDFsV+MPu0yuiiMlR3iNSw7QFdYNWO0zO+WPywat5+RC
7UQGM2IFRIIYSKjPIxzltHSW9RyCBM188ePUgsr+gRB/L3JIk7wKCEyl8gpDb7WS4giyCm/RwvR5
oUPmkiJDTY7KRAW3NO2vNUUN22YdOpQb0g4RNcyhpglZz08vAh5NbskucfV1ReA73Zv/wycAqzxy
8Qhec93yOwXq7dnIy8LWC/2cflqhJIoXM98tKRKYBnsbn/TV8uuCCVbngWh1FWfGzKtrwB00HD3R
luSQU+RngKTiWjIkeoHQRZ4R8Mvf9d/aYBMkExmI1+uR3IdeFReYeYBbompKHWwUWnDDhrdjIg+S
pZx8MqQj1YPcT4eT0I16ifS3dKJrjpyVJ46OQA3HLsIVtfk0FN+UW26JbeWkihcIVo41qN19LjgB
NBM1d+eQSkm9XA+BWypoaMPcV2ZghIX7v0F0LOARO0v/iCvkCyW/a9zaO1LTPDo3QSMHo0hYKj6B
yP1i7OoCPY1lcW22+yINs/NeQYFj04B6T7CKezX6AplSExUIeLv2Issms65TOcUxI+opMKeSzZf2
Iv/dAe/yBq9Milb9arDTH/nDqyT7SRwKvUcb87+fzkOcsNMB0GHq/w+AZFIUISy2VnBbZGbfq+NO
0I+2t3CT6CGSpmomHgo5ezS/yF9fdd5TPUQ8AvGpa+pBBpuw8THjlmtpT/MjA/MuiEeYX52etfiM
67zaPXCiGspqqUqXCUPLBB9XQ1wOrmiUSvvg5yoUfCqYBpTBxlKZWrr8h6TubsFfEjHM52XDds69
5lNBrSHVNUMsZ1/LBI8vDeLRtWmGh+LFkXEIUB+2SfHlduALJIt4sAWDbjqVBqwFOjbqLq15rQdO
AFbfUxucxWu/cT2WxBaY/g/NUo8AnXKYDX0YalgUQ1yP/bdjZkS++hE4Ny0Cq6lgy6gGJlmVdziy
/gtk6d/+fj/sY9U6oWC2TyICudkEHeyEUZ4lUOg35z37qXjFthrPKBhpFq7KI6mAYcwtq/OMQFoZ
ntgrp81qeSZFbPAHIEGNOeqUUXy07Xz8htQ5O54fSXlNiR/dMXzTr0BYE9wNdTllQfjnVZEJMgrx
Ok94Ertc8wGxH9SRX/syigbHgYyVhD8Xe92b0LqKtMwwyeTzBtBJLtUGxOiR8Pwuo0aYLznVgqbv
Uqoid5yH2b97pTom8B9fEkGbFFDdDkgrG+WJKsUfWx4JTsEdChS0CM4u2viaoISz9LgyPbTUzrJm
SQe628rJCqYn2CquTJ3CDc4hp5HFWrhdmafYku2oFYCJRzSPSAXqsDTmtC72kb1qjDZlWO3ZhJUo
HETmv1LPSaW17scHIcHm4jouDngJqJErDJSqC5UvCDqlzXJkTW7XuigUKsQefXCqk56ox8Ket3Gs
CH2sKGIgoLC/qL6pB9Y6YxqUHb6RryMseBBbdq4Da2YzG5aVfdNpfcPh1hrjyFBhmyQ0xb1Xkirr
rg6FbOpPMUqXmpUHeyk8Q6mnngCteANHqQ7OZZRwquggA/MxnV8WrYQygnKRwGIDJYIBjAkaiaWc
Xotyset5dlQExF+z0XitkdO/YMtI+tU8k09B4XCnBhhlLtCHi0ocrwmQbbhC7THdTM9jLqq0Japf
Oale/YIEeSCcxGCYyK4WZYAD1Oxpj1xncKPD3XNnd3Ox0NvE7fmiT7TCZKwqIFmNyWfqPaU5GviZ
XhO4q85x31symG4nkw0vLOhjQTTC+I4DkggVIai+BWpO7gZDFA0lWYHmpB1pPRY7Vd8Mxqe7IOWk
PityLkxxQyn/DvUB2e+bJXuj6JFxmfR+DGF6EQm+Dj7W2EM/6s3IEeqCnwpmDHKsHQcee2hJH4Ri
8Ibn7pu5V/4xntZWv5AtwvlnJDCXmy01BWC1ez0gMhzc82uCtYrJgQh1jKYnM4dAnhiu+b6TSgMR
BA4q+WR3lXOvY3/55ye10M/VJGEmV5vWa6JwoDfDcZe8uVuB044EsJQyBWWxXZkLaP0sSLdFMGrz
wSDZIHa7wv3rLEjFoAICjqu5kbTVRpl9hDSQuDkHZxmO+0WPN0F2GEpKmsuEVld8mFLHmvKdNzj5
COH6NtoUE3r+dYaAvhC8WCnx+w/eHwAofh0R+JBZaIcPcw8PLHWQsGdsFITRtY+qNM+H4FeYzI2j
fmFqyKeiohEPGCSm3Rx9xINFZrmragh96sqLr6fxWC2vQ5IDbTMiB86KXNR57ic7JoUyqQLLu7CG
Sf3LqseoDOiPv2jQ7uEkNAaprKFGbd19Gu07B+UYF81jMDl5oKfRMqTYGCxqi8JFNPHuXlXDmSc2
S78GIU93QUCYgolNEeioZB/uXBW8TquYt2QkTjxzp2xr0P0VjGFMeP2UW2zcn6SwU5PMwFxJTiL2
UbkCUriSoj1ugN6r3NYDHOuEN573/NFlcOSd3BkJgM3HS2VpXlHFNym+it8xeP0HQa0zazWDp4dt
hGeyQANCO8FAnVuWODw6S7PmFQQyjE+JKYhO4Y65PwUVvYo/MWYZgKCaJLXRXjT6BgLHqNY1QsEH
bnrksCrIa8FdBogWCAXKX3SyYMJucgmeB7ZZdDWyj4vXxoHUjDqsT8bzwfIDr2sHEpgOp86Y/mZg
MxLtNFmQVhnH/AXlbpfiis5OXBa8fNxQReqLoqMdRzzc/HLNLDNEvJyGYW5z/K+yzIarTJlYz/7n
9AAQq7sW0FzCxNydZU6+CBxFh37UhlJCWRbzBQzhiYqnR/VM1PwqCqdnz5q9/SWGoDq1YY/umeP8
PjJ2M56RU5EwEbGoQls6orwkb/6Z5MIH6bU19vKOAQxfbP1HcwOMJUFkSEW7bGEE4XlrhwMrZmsW
goC3pGrhWaM4zKdByyZazIrVPmR0MkRQWUOJC4eHIt3/sWeGr0wCEXvWstbvigEn7acb4AFquOon
izDagTMKrQ8WiynY43dzS6r+NPCbZxSS00+l/yEdmVI/IMiQCXaqJQON1xvs8MzONVKR4ahyGsIR
WstLRolmdykA7JW1U3TccHHo+WawqZbDmjoHXW3Lo/gE4Y4KM4BqKc3R/pTrf3+s1VvnfcCEwjG8
cvE29aj1NiedaX8Xuj3sTi2BPvdR0lItsi9oPzdFUKsUDDPf2PiiywJBQgvD4V00okWNDzpNcsi5
v+PgcqIWupjfPRqNieiR8OR5pM3JWTgpuH37FfJPkKFvLolzBpGn/wuwnwvwwbcg2c+xkSLywJNA
nJ/iKZTV3h7vk8ZhrulFffZeL7dhNbr8cr9snop12ng/AM6IOLUj+u3ioXEnntU2A2Y8m3P6ujU+
b6nJdYWU64EI0LWXSpeeApoBGVoMLw8j7IPkG/uRGp3ZuPl1F3KJ3rcxnITTQuf2qc0J7Wv3ULtv
6egwsv05Z7/q1SruXK6HHyNSEDvl/kOZ00sb2fd96El0qlZSGQzqfkxvV2mIOXjNrtt+qfqFbPwR
QSVU/cXts/fvC25OrA9ZTAddYH87RIirWo39NZcDl81K/61CThxE0s//3/p7mE/W1eKxkwAovzT4
/zpXUfipxP4bJV+2PKB2rajn4i0Wf6KJQpJSGQknZ3lUeXineK1ng2VJuOQ2ULQGmyiPDTy7qD22
Rve55G//Upbl69eoNEylG3UIfCoLqaU7UqthvP/mNx6f+79jzxIzxmJx/bNFIIbYdIp2Knt65v3h
wun53YrGtneS6WFIdeMDWZxi+YAhFXuBOlG2uguILPxJgehUM8lB4P26mQXqg/8orCilYSTEvb8L
UGcJIKqHTsIFphkXAXnRgNrLLzYrECZEfTNKgUgcw8v+Dj/lxdb+6XN3epdDJYnCACtoS0nsyNLM
Vb1jqsNtaSLf3AzSd/zyJBxCGCSSrgJnTZzGLPnfKBf4HQb/L6WDCiMewg81xrdin8RhSpzwVjHN
V6BbGlfm+icqORYWRz2tu+MuyQp8Rw1vO9c7GwyZmlnVYiF873QQC3Bd7+4gR/lzKfqDhFTm0i8Z
AJpw4RCb855os7i5AAGx25aSGiXr7Inm6d16Qtno46uSAvdXSu/21AfwnROpZWc7jEnN47FlQ2rI
RmcpYWYCrBbLitrjvo7WsKrHs1nI3QHrDuXfauXJj+3/nNdmCpdhTU9E40zj5bGduAWb5sJAPlrN
cOkaew42dg/a7A4ZliRQ0ZWniVHMVoa1GvBw/+kLxlJt6hQPXLImRhT4idqS4hltkIIg/IshCw0T
a5xrwE6nkSup7R3YHsd/qPy70dfrVVAwK5vYJO73xFovw/aOCxjFWmbpDGaTAk0BXEn1OlyFXzZM
wddqZFCTPRuHE+b4MhPjEK+SAzg268ypcWCEoZafNSdSUQY1hKe7OOGl44dDWZ60aLxpZgw5jNde
z3X/HJ1MypOjfQ2yrs8NGYRyKW2kIFoQm75VABBUG4ul2ippMvLvTBeLZtGPjmQ0hu6wV6cM3gfw
8XdqIT/sJibCG3571Mz3Bt3KqV9v9ZrRXu33aAj7cW3vcx+2a+q4FF/qPUy0xFoplL5lZbKReO5o
brcIKYzNV8PliZMbc/0t2NmxAGEEveCqOHWbVoh6vKRi7HGIddUDD4NYEi5mbLWs2QMGZ1rElC2E
XRBOeK9WTSkmLpG4tMQWkM+x2nnOQFLNgU88bb3H98nmipFkVw/Y9fx/AqQNlAEB6sGaN59gXAXL
8yjajfQaVgMC2OVnBcdQzuDiR7XuVRB4aPwUfVIInCETgBHerx52Vpz1zUXuCm75VTGyvYoTj8DO
30K2KWIaCdBo6EAv42MIU6PKjux5P7UlvK/LxG6FmDFdZqcczy4vrpkhtkh7m8ENlaLaxzIaSil0
qgvsz8+C/XdajIbW+vvc6RRbIzDHoN4hvPEmCae6TwK0TtQzzwOUmVQcSrxBbvG5Ey9jcbaGcy5/
juw9uQtSnyw/0LhWTFJ9ZDoWYNd289uh8mDdy7HXdHxGm/59h1varpcxi0//Qzthpm3UjuFooAId
a0hahTGxTaRl2L6ZPiWb49fM9xhJzSXmzhg7TnT4XQCiy1x1VFW3n61a23Up6D0Y3oVg7b0aKBf6
GgtjytpCIYOT0u4DPHeAamyxJS2MIWDmyh/OB/a/m02DC4ihN1zhTETKf/SXlApTnsph6OPpLgTQ
NLI/Fr6HsAdFx79afo5jfwfzvBZGbABO+ehQAcygtmfimz9m39qUFG+md8ifbS7ic2mqMCiqVt9R
bddq4tunZkZMN4w1uysPQUK+r+BtVki3fhls3a9YF6oLo/0TKKyUcWSemaXr8zAZcpgPJEkuagfS
qAuiwzB3zYo8w0v7FGeHIfCmZfgpiFeolv2CdfFlZk2EfsbVIf3ZIhlnPwLEi7HUPABiPqw1ZRiG
5y6u0si1Gda6RfWmCbwux9FzX9CYL7JVL/IMuqAosFH5Q3gqEpop0FnMhWIP4ae+76boN0FRc01c
RH+Gl5lhcKX5tlSWoLDvL6C1UGGo7M1UTNrCmuis/RBC01LzPNrGFNvywVTNMqNLGkqmR5pEF+nf
Z+9A8iuDgJ5eV+egy8FANkHBJXuaDPYOxgDPovBQihnisCZ60QLvXg7WViWQ9uN/Dcv7JvDCEPTu
FPaDJio7qMvVrIy8RgdIbtiWQjGAT9WguUVHvwsMihxdpru07/21C8M4mXPdwOKd6rKYfDEOG3on
Q76bXWtZ2pYNwyYyqYKUPE/3Q9Vl7fARnbehXnZyxwE8bioC3Ulg6JhWTUuZq5V8B3/fD2DsqEze
HyoldY6uoSWGrbs1kL7dFLhhmR2MjZtpjfVTHPsUi1aDCyRE2UqfCopyQL2K/NuR9gDDlQ/mf2vF
dDTQj04/KL7PTmvk8dfJJReoLZNF5dkXZyfGjdHV69cHBq8vtNzMyb5UEJpo3D66fVyP4XAtf6IO
86tmGKl81nXPjysSdWRRi5Qj4rgeeq+PvJFqvyNLWZ7SwiOKT/j97eEbjka+g0APp8yuAYKzb1bG
PIFZnIeSKh7Snk8LeIBhW5mODbXa4DS5nV8+HzWt9VVG/2DG2lbJJKmoaC0JhD0A4UppYpoqOA42
Z8vuqyEoNKwV4xSrLpAPBIEhIcDvB2MYPreoeNqQ7WIyGyIm6x0XFU2G4xlLKfbPL+ZNs8RUp8re
dh/bPU4hYoMjl2Ks8CJ+DeoJcTJeKP3kg/URghkxcwxLZ0SLpGmbzRC5CpocDp2Speg/EWPfTxSb
jdI+6CE3NE62MjYS1l327tIhQjlSpKCC5EbgSHC0byoUZfQBTN1Gvn/K4UmwAnv2lU406r2iKrrr
JS7XUFpx0ripziODbG40p1Kmn7Ve/4SgvS4JtEXiQxuXvJf3DNXiVF7aRWPgCxVZayTkM+f0lLNK
FIxjjEA4/iOxPsyVvyx4urjpPVrCwxJFOWZ1YLQ01vfJquRtHQ5SrRNmj37SYcOpot7DAFLpc5fm
CRKu9C1qgteTplR/diBL9TMEBdszMwDXo8a+CsT3xpv9AbBnZxA9WqR9+R+aqjJLTpytc0AleZ1N
11fmpDiMIVQI+Ul5zaAKYpsBCo4LHckf7FPUtjHPEpW3DE/sJTVYpIz3e9to2KOjCgIlakGG+p7h
jqYXtc4HqaUGbJowE688HR+vs8B+ydXyHmk9j31P5wpTFp4z6GIwBB55debP52jo2m5SfRDsH0wk
8vLyslzwUeAs2UwpJiu1GUhjvA80dI5ESYz8enVJXs+o9/aC5F2veLPiehYyo6I8/jDiaqDw7ub1
j7XhN7ZsA22rXEGfrVRrtVmrBjUcC0hbe0Fzok74kPEG/ijYZ2eyxjqbXiVpBiq3PIwohFxeLsqZ
+cDL36ujqqneigQii1myALqK070ns2/BccAsx8g9EjGxFX3C5zGVXaZAZ04jRHwKTkKZHuEgv2rM
7vDXb2xgCfvhM8lmqtWvLus/Y1L8uicjG8jH3edHXAnyEdvYK7t6a0TdfNlcgrr1tcqGDvo7ITpG
n07lXlOn2o9XdiAeDolXaDp6RGHhNDO8KSbZysK9nSlFiJq9RkQ2u+Apquf9H/062SS14SwqqcRY
MwxTnOULDZ1OMJOYv0qxcGdESOqzid8IJf//x8yBW7Ua1gD2kzopba3JmQlJjNSZq0eZJsUl97rw
/c0ehxKrA+v3v1iitL/1Pb8CURLNYfPcqRYc6/FUBJz3CBiIPiogkSDKi9OaPugVK10rU9pGdDCY
lJFss75hd5SMU3OY2OuOnftL1IUpyEMbZV6Qap7uFLuEPm5BPtoqm+EKLnXjt55c9qiNW/7ZhiBM
0rTOXExzBpx7csAAqpbHC273AIkW5JNYteEOKx9tmn5GOBcvJ/FRAW08huqo3Yl5Y+ekI+vLPRbI
U2Bo2ZBavYgAgtcGalEI0bfVoeUn/uJh3nuWZ/HmsCFtYOQ9fWzk/gxipLoVis/T4KzQi2MsUrJp
aRAaB2JdefqoCpofC1VgyBWfSzUCbBO2TVfFdZh7ie9YIHTRIbFgufa1Yf44IS7JzhbEpKW38/HX
JHbMal/R0tKiPVgczfTDjSdy28jNH/ToiBKnAsOa21fzMg2P/jC63OiuPCr3hhRBi2nt2bgMk8FR
YoRYnhZxQE//iSm/PneInY0QLhJ0/1x0e5gscch4mnAx3mPKnIMv6T6aAE4/akqf5J/Xbx5qHMeV
k3ef0tkGb53tLNr/losX6LMNPinkhmxjBXKqGfkEtETK/mYaFueLlMdRUUyFx6ElHYBYkW8Z7iAx
gGpVjF3saBHVm1bOYDEysECQl9F0PMMFdq+EvqMwHUYWD4gqjxIMHcL8YRLHx8qgYwro1BEuB6BG
8bM2rWzAza/lZWtN1OvNlzPTA8DrhL3sHQJ3mUP2rkQvjRzWq2yIUUmlxXNUJ8f5V6iOQOZr2JVk
YCLpv2QaaonXeQfURlJmSLfbMFUp9HXPhnHIOyGRQsMxHyhW575yNwVUOMxDRzEzDEBWX5uanUOE
YftOOhj5zJbSMqbphYsuU/Tu4e7qK0QD8E1F/YB0knEm29HSzdiCnBPdHf16tm2cDcv/VysUDb9G
OnCtTIvy2K6iUPsDtrIPFdbo8AXqT5DMVj+zh8o35D5pFNJ9ngF3Z5yUdF6ehucqdeykKrf4lPnH
b06TzieoMb7JY3rVjC7Si8tQ1DHHpfpetQh4UCJiuj0NcrFjrvJnyaqk9xaQkiJG+iHl3IjftWl6
oWGA+jPI73N/EtZGdSqVSBcqOlon2XAqi/tiCMZhEm65jIX8mgBeKyIgrC1rkq32gcbVLWGe2awM
8kvb8qTxBBcMOQQ78uujXJjtjQCFPsM4MbnEuH4FnMaoQo25z4/CACL7J4H3EGoTLEdDnFvrBY4c
yecbEiSawrmAyg7SYrGVx+p7Yju5FxtCp78YlAlIDt72iZiwW57m2RszeV/tHQu47CIUAT3XPt7N
zx6J6qfMmqUFLtbhGj1m4cFTGaKL8m2ijAQ60+hvUTdJohhdDYukL+U9/1bO6IzBG24HOyve6w9b
n9InKcHOZRO342+42/WFqdWioLRSe1fUtz2ifdi31SLg3VmvYIY4QeXcZWe+yeZuzKtSATQedFGH
D8ZVsfS/bRIUQToJLmCWgBCI5XQp2mvIXm76r/b6dVPXXAlOYmh0l5v02YbVsRMT4fyUShPpKTCT
oP10NhKUilNGuK9KdAqAmxV9ey54FNarU/HNGkFjB5IiuHr9D9SjjVNgsIhkYfrKFbVEyF2dJDoc
Gt94qE51K09b2/4fSYlTgw98yjyQQMhknx8mku71SgIFTRgyUXDS/LqN4XX+x+B2bBrEfmxetfDc
orawEjdBg00D4wLZ/n5cKM2RyUV4EtDRQqh/0o+a4F3RcVaM7ORwSyy06+ModPmwwFblFzgFCH4A
/PEcaD3xUWKeT3Ss5Q/G5TtwnxBt7PQ1TWOrplkswwnh1uuS/2/rQtKK/vdR5aQE8V4lDPuTTgmn
KIxJoA4MHgoAvXqFvp7Tyv3xq7PNLz1+5SXaTMIStpsL30lWdexfFqmGXoOhU3LzOl4utwkumpWG
8VHGIgwCQFKah6e0UlrcazDzAdTm4YW44DB+nSYGmiHsbdd7USJYKYp9dAA0wFfGDxEd/gq5JCN2
pU7GsYvHwMrlqLXTb609drMFXMjqoiKl+Vd2zAzVUX2Mm+NQhqlrodZC2FYkRJao6bn2dQ7KZCmq
m4816o6PEvsE/Mz9WWOlzfpxUvNffFltxVz1ll+JH/Us0Hz5ibn+37pMGs3sG9yVMG9H18pnotZ+
CUcMjz9EOTbyYwDFY+QIfmmUI9FhTGKbvn5I8wwKmRgktoQb3gDeRnktVemgmbV2iQve9VkpXQzl
VwKNzwcMHrPibEc70JLC2mcWkLlw04afq5Ek5eTwjo8h+sx/ot421QoqdbDX4+FQ615mpQvWVrtv
r1+B9aeuIAvjvTt41njGZTtPlJRD1U2EG+YJhu21+zgBCF0IO+uVtUd3cN8BUxj9mn8+Z4Z8cznH
/b6uWZElPYSjaUP5o2oxe7G6gh9itOVrQmOXQkTF2fCXgRTv9e4h8/Il+JX6RuA71vJWecBGdXHX
LTvS5KZVWeN9P7eNW3p2pnq1i7lGrPRG2+g7F/WLK3nKKkw7RW7JcENsApE3mMbjuf7NocQxZr1X
/HuTVTg8w5dFaBF2yzr0cUJ5kCdk7SSQ5t2j6QI+xhos+w9J7AdYJKIRRbQkg+Eo+OwJvOXqZSp5
N1ufxQHV9oDbs7Ud+bWvuyOjPuQ0KGsTHHIe44Qy46SZQE4wnRcav0+MkTmDSTMEOi5dIDd3pJjK
0BBqi/wU94v8hAfbaVotNlsTuk54II7u2YQoS13MKgEQd5ns8AS1uIhYAAGoUowT3YMjIM5O1md6
DnN/e4ci3noKlWt4HceizTvwwlGShv5d8pYxiyH9sBA6RjQDIYXDmXiSQYHDAueISfhF7KHqCVc/
zz6EXYnhhcVzgRTTjMQdc51jhcGmtMYbmorR3OtfLzGvN2oajz8pxXYr0Qn9Y2DRWK4CyCTMKba8
nlDgwSUuG2AWezMKy7R0NWzkMho8rcuyiOxbi8pfOkh6qoADVbBPbOynC9g8NbCcvX6VGPyioWZr
LoUyBiduiH5ol3fonG3no9xENEXIUBsrAXheTT/AAIfKiktTyOmZo9W4wScE8AfkCQ+28ZS+1Z3y
FqeYty6cbRKBVDXthWOvnx0gbhi7OamDL6GaheiCc8M+Xz7DMp6St3BDoqh6TBtzkBrR8s82yt6K
mIpFG/N9xN2X0UKi0TR10Z7bw4CH/WXxGG76/Pj0pqoLaEccxunkN0si3BmLHO5tYuIwQhSVtl3q
HNV9ic5Ij6v10P8DKjhPLmpaE7PXyuwVaZU8+rPUXUyGw8TculZOy2GZcn46l+p920QRDerryUra
SNwRROCb/5SNSvThqkEkUblDrWMlcHxe0N28M98khGSROtfzX6+XnBWVsxYCXCRSPiYFp7I8tcbk
/z/ieUY6PiRd5+gCWyqBwJGX2j3oGhQ6QPRrFDnK5RwN+PdxLZ3wKmxkZiX4eF2EH9q9vCabMP4A
meowt5nZOihN7b0F57QrjHKdEZin6wZluDs101KwIxQIwLdg34mBnoM0uemeYfmohBLLeI1c6WVP
biAuulAeK/yTEw3IpssgpFhwNmGNEQWfz9eqXgXIRM1xCcX0gtL/vZ8OwV3xuG+z08221X6xxbxD
ptbIP3j2Qgv2azOI3WA4BMtt4B5GVrvrBMT2quuMxKsN/lVCoE4eawXO00SGlbPzPyDaAkhgvRGk
dtCYMWLK2SfUf8oNcshScuh+rmDIZ+zk7iUT3UoNRRUJjXbnzjWI+9Ltoxz947kznehlri06t7En
aVWc5rZjT/ax082GAwrrJld0Sx1Lm6Dr//HebuPW0XJnuUnI8cxy54mmL2O4Py4sXTUYzqjYfwxU
NDRCLkUGnOo0MSszWWTh8VQ1kUUZfB6yhfV2chhcimU04cW6Nu38xhoFBdaJWEgKgfxwOfBmc/Vj
CJEryDddPylpP0YMzXjEzUUdkkA8N7nvb+bQ6xdc/diIKQNtNLGi2r0U/0lsgqkpgTHxGYe5u2or
w4FXgRviVDA49/WnlyJBshIGAxjWJwXeryYISH2LebVTHG0JAKmw7mrBPJOq+Slwd71KB+av6pTf
U2KkfazGChhGLmZ9uHchD/6z/T+Ta5K3Nu7bQbcRrcfjcC2MFuY9by0talkiTMJEwNMt72x7de8c
4tTz3uZ+t+hiAMqtfKiUasilhblFQAc3jtWEhrSmMMdeZCzP5VdILtb6Z7U09OIeNSvNWLcdvpka
IeO5g8SORKtToMYkPBLLg97GACxQeqLtBH+UmhLUC4hf31olkgo5KP0Jtpg9Ca86FcFkE/5ksaCr
OteEMO1JlvYPuTziGfroVK+ljMIHkUkw7M83mEK2dy3f4B7nTDHsz9i2DIge4qJrAFz3uyfFjvRV
VIrQnOHd46gRO0UUGpoHo5EMH0nvdx+bLZyD3o2kOG3IGeLaQzrabubPduQAtB0EosOwo+P0XJYY
nZQl2VbWKayNqHbCAP+oLbgaSnERu/Wr8x04Z15IkVC++0a005FNZd+kRWmQ1SWEJHb1wslUgE5N
3XgMHHDENUWDI3TCw5jJ+qHtCqf6XkznCKLk6i43PFA5NHvgiGvkwAmpE0bzmFNcxH0cc1fxxBXl
g9+XCELcsI2YqKDGOyFfQLxrh59AzQlzGTLHAKBflqhK5cD9PntoI5V/I/xgL4Bn/HUbWjYgsKmd
6bQeUSZZp2cwLQYyawYeZ7jHIjrUoxNKUk70+mYuhql7x0RxIvsmf3H7lOrot/sLZL7XPaW7yNCa
v2P94KAmiNqBInl+ZB5KXJS2kzo+C2W7HOhOCtt5eQSjMc3PlYLgPomzCWac821J6uWPZbVi3L38
EXiDLYGx+kWiHVpbs8a08McfQwasL4At1S9UbnJsEHH5/uSyWBsLxTxGyI0SYbqYxXdZ/yZfX79m
4qpKStw374l0h7lJZy/GCKTzFkt811gVpqCF6G4qO+uTWRIsGRoM3Sxif98EgGBhhNwEMLdFUV1q
FRwtl0Z3vzmrkmvDaxHlCb0YrYJPjNWtTBqlDO+HI9F0KqeX8CKdkdKWrBS3LI9t+hplA6trNidj
1zFLF9pdo9XlNaZd9mL1IQDXY6Ds21Y2Wi8VuFikD1m0Ed1mJ5g+o5YakTIkQ0Tm798j/bQnD3rT
16A9Xga8OX8mloM0lcXNHCNcmn4cAdSBDQuiA357guzMmfSmdbnvRcWRfEgvLy7Q9Jyuj0cVY528
ZNsoIcsMpija8CQAniUhfzotsasxbpNukrEOrc7uciFKYc6YL7JfNwn0DOAy2JCP0aY4479GmOpX
UiBgAQI+92+qGC9vaeZFiuSfp6fKuuCY+gVLeaPuWMuqQ/ZoAlnSPpgH4rKW56mvtS3pWxgDdTIP
NI6VScKMJ2vF3Vze1uVefkQJ4KbADpLzARExkcH+MiVeU9c+P8x2rNIxb2gesb61LgLSj3j/tCLI
BldxZ+x3phoMbffJ05bQ2V8kEvqUOCfxOynRVtrlFhNqHShh970tibVqejpdZtb5y8v95ZEBV2ZC
H4bgFTyaoFz4LIlNvdHfaV4DZeCKj9cuXfqxeuzMNRpzpLnpZlZBa5iJKki3f6vsdxSBJXaLQ8qK
W3+5QoNGhFv9vAMQZNvFe0zPksgTFyYItonJPBjn63V2bpoKbU5I2tAJBcOMHnzgleu1pkdEyxBP
VTaudLRCxjHLef8QHnhCvKX1PKM4wpVyz69zZI0Go2AtYRc66emfKkISLUcghXdxGqzxVG62K+Xp
rzJNw5FIRTeBc00AQ2EZ+MTnU8Eei1wV9fpityrSu1q4GrSpeQCvh0q+4HlJ8HEkcnNYdmKxh7QL
ZyJQYFB1WpIdmfL5Vw21yByZyub6QPlLMexUepuouJ+JMGB8yjUPkMq3m20x43hLHpK46grkapK5
psY7IbNN1EhveP97V7zz59+T1QEm8Fw4p3DBROWKz+4AGQ4fpY53z7fgYaU+G7RaMGJx/JiJFl1P
w//LeOVPPd97serBAr2nOBeU/ggcibFhiEvXI/UanT6ET479ZHgGSjBXlFS0K5nTvioGvsLusG+N
UumIbB6mAe0NvattA2Gs3RE7df+12TJlaZ0VhhOaL/+DQwtoD5kLQctTwVH6DCwx+r80w/xBKKK+
LjoYcMktR58WHBvUbWF+f2fkiNnhSxl4ZzEQurDEWI/VPmva4BvDp0dEI6MK0gk9Hb+nNFyqW3nT
VbkvjZEalI7ZgQTCJ9lorvzvbKNIjauvt56Exrpt3BwEck1F8kDXU3B9J0UAuWdWGQ2E0ekM0gci
CutwGNxq3lPmpmVOB5ErRhOEqntMX5MF6j2hRqtVP6KO4QkunHuNudskpLw6CTSelcHxbYb4kqqN
NgW/rjEvWLCVu7FmW9S3kKM0GhjU6YUDiicCWivxsyKvbswS9n2Csl+pK9IHLXhuvO10RxMY4umB
RHyXgrNzj3x7l4/XicEhdyLPqrDXLNSvf8kpMrjLctb9tLrxsOFZNq1wo3s/y3XI+2sl4llgfrHF
ZnWcRnr9N4gtSmblg19JuyijRSo6sgEz3GbvUPh5yqmV+mqAkmVMG9KVi5wilVMYOSPZVN/zNBb7
U3V3g8TV2HFKm/qS0mhedy9VcGrAb8HJ9WNujRULxU8GAVBCAb4Kq2jygLJ+wU1UDeure9I6O3qK
ZttdH/Duqe2+CHlkTqX5DHmzGaEctxS6kI8v5bW//8tnY/jUPFS/rH4wj0+CjEViToolGifZenC0
ReXomijnOZU5fPZhW9edIYl5QH1Ccr9QsECyD6oQ09DxjzBNBcV1AY+pSKRQYrNZZOZ6dazt/YSh
6PfX+CAYQO9ds6WzhW3ff6J2pqcIGjUuycuEuY1BYCaQV2svQnG5w2rYN/RV6mN9J81tR/ih1J/a
SkehyfnZ98/uHh1/5FcKQy174Tfvt6HU0DqvxWpaaFlnS9xzNfwxTyWS3BK2A1ymCtF9lVWrlYUX
/zkhryMD17NaZUihHi2y0H7A6U9o9PeNUHuNy/8Deoms9/0YejyyTBhhQ5kLk1H88ndbaX2dFywm
mMLLYEVhmnsmL8Qm9p9bACw4BZEwOTYBeEKqI/oc1TMZ0eYqRfJoTmeNqpJ34mHSor5Bgf/G8MWq
ytCIQ98pKj9SQn2SrcNw2Bh45Y9ULhcGlySvduVH1JemvCEwxeaChT1uoOJERjJ1jfJ9uHoffflB
zQNv4o3x8HGgnzv24LB44CdhurpCFFqs5M33nHzdST1UxgZOWhscJLin5rK2hnPXGNuoiS/tPfoh
QERz5Mk1CKAzSza7Zmj3PQha/+/EjdL4OblHgZcFQE7dt2tGYpELy9y4lRpghvDFB137neTCyPhQ
1+xoc+VggM6l3sjouSU8l3sZEgCSMmDDyYMX6hjbYjTpVhiOtB7mZ4dESlUhe0NXCsvdPGVEZh1c
T/AhncNUFQyP2+PgUWe5OA/HB29a3QZGRebGnsnpgh6sLzIBp5VHXSABHYMzZ2f82yjl/GhYbMPH
Gyw6NWa4pSNxRQbNAdWQoooLvrv6uUo5ws0BNMWCwzADOTkapTCCvVycOr9KsL8JX8lBqS5196XR
1BvlOFI2y5Y41Si3SRnsXDZDoEYFJRoLIkr71LeMmhB6K1rMcUIO26ERP4Di1lzjDa3M9fFr8TNA
LKt0FKt7x5kUoNPO0npas23uurryNNwbF2/wYkyw3JgOAryZNCjUrwQKISnliLPPJ7BfgIRxgRDb
5HMGJnkRs2alwapC+Dq85TGB/JMkQxwQ4z63zHzvODLovuP4baPS5a0ii5JuC2qS9I0qAXtar24G
sBK4gnQbubZOVjlRkntKC+Anw03yVIR5tcpwzcpHfEiIUazPw2IfoKyiqqOM+nLOQbi6WqqMmLmU
Pcr1b0SXBHP05OY1LXr7Rv57UXxzq7Mgm+1wcPTk+7iqaDVwWiN3osWplvr8idHPO+CokE6Kx4qf
gnZXO1MA6tvqKgF6rRRIsz/RJgzixrAZRQ4jJqSjLK6WKKQLGeWoPPVmUcty4Up1fEzC4vjt+3rY
FOD+/80jmay8TC3WImJfgLq/luCI85R9g1srxd4MuQpmSmKKroF2xbAGD2a6aQ4OgEJZJjfLx1ha
VxREAwxfJoJDE+YQQk7eN5ZXNACY/OBlecO3WcsyWTajGz/EudPHsIiodYKDpYi0WZCPnGs/Lfie
AfPVE/VB5iNFnELtmVo4MJ2IEoMtU/bYud2QojO8RUG47WTDtmdbT9ZB7SDgr7MdmH4dZFXDp0Hy
0zli/Sukd5K6Ds62j7FWzv5y/osjpCd1KrW732HBAOL4eMP6A6acLGJC/VSGTWjG6gWcTfnhTsDN
jIHpqqh6anTHM+QP05e2fZ4eImKg9XriMJKalYoi2bmJpcP4UJBTaEO7USIikHmVQZ95REXaVW4f
Xfdtj9zoKdMx6IueO3sKBsCxtckmT/iEQBlXOEBBU0A4cXTsZ5SQ0c+ytvqCC7rRRnFe7uLMOveb
nziZ7w78kUuM5LKNVovgXhsCWD0dL4rdvNqhR+Far7mQQ9VQFYjefZLR21De8lQ4shhDSlQ6f8lZ
zAAIHqovIlIFKdluM/lzskrwuvZx6FaTG6sQZ9+WDHlwHVttOLKzLitIxVFqHiWz64bdQvc/nYlI
ewGjgaQxCF0KMJvpdGHzWb7KtXU9lvePd1Bm9vUQhWJ7OslGOlx6Eoaw1jBRdggMId4VeT+gF4CA
T/KxBsU2pTJK9hB1v8Uk58uGH2MT7az1wSwzJj2lYPKER0qyLMWw1vjnct+qZwgyslK/gztatrKH
h7V8dukzOB0m1gIEe037+SgCcCeo0RRnBDILshsDPVBDLpVfnAbw9z5NjzLgLl7RitqIqfvx9Rfk
rxwxCs3wVF1eGIJYhtY1aroRy1Bt/HFMpq36jVuQxu3WoNAbiuuEd17gwADcZT56oJNBFXVUfr+N
eCecLDqBMAAUvGtNA9XqaT9+kSg0DngZpvZlNRo4AkCWJ/mgOdChu6DacHFGyGMwiTdVKZdbPKlZ
t5IoxgwFlQc0GCU4Zl1ZhJ2wsdckTL68ho8eRzA6paJhymbFuRjSJfjp/Z5nPdCCpe++yKAcEcCv
03/34lFIM0Lp955qQPASwEKKNg3YU+VGCtnVnEygEon46Ev9yoW9j/1R94UQ+0WtSSBAe8pmUTZP
NKESHCG3g70oLbwa+cib9QsXeNeV/+7Ot+NLsOJ0OvF+oq0nchFX4I7ecTKxjniHIqdqqMb6gCSI
sT63I7JRq05glkc9GrRqmiPCHXXFQSoK9CVODeX7S6oHMfHk7/keAhtTKaZ7FwOHoUdcDfTNrsE3
7DCqEqtDPUPyy/WS4ScCI/aFuvbMRmKsahskKkJSN6DveOu/5jCl8C3kCOF+WvWns0bDDO+NTc6d
DNS5rqMFGvW8X4szlWCoN1XVSRcqP+TQKf7O1Q3akNUjuvQEA/MvtKcoOV8VSYSssY19M6dzns+H
EoJG7OaOWEoJPsYjzxOqUtmII9rHy7WKmjNJdgAtoIFS9PZlMvKu8ziyRmdk74Txqx0UzRr6Pxgn
5wKkwtA9LZl0dTnnY3EnCK0xuWV0BB3Rosee6vB3FMZgkKLqc8/uIqrvsjgDxxGkHQEgWls9/7mX
XmPLv0yAiN24Jlmd0/ES69GbuCDuqYH9n/LF0y5L4fKRoCaEIsuFiGgAktjuupbCFlyh3IIih3UJ
NgYJcj/MvDQBjEJYFLTeVfRPHu4/qvuV+eyhBfkQXDZaWA9i3kuSWnqq01cK9i7CgeNplp6Jf8nZ
SU396BmpAZmXpKlnHN7cCLe6QKy7NhGrZkm1FbYY+G3TY0lMExTyAEOZFuai3Iuy32owMusdip1I
VClCZxMC4yxC4q3761CidhcHvym2vUsUG0fUTl0A5DnvwahCpfsDTU6K24Y3ujVpiv8cLcoWvge/
jEsorxIqR8gHerbokO6k5mRc80SAq75ZWCOFEgc0vOlxxRZoWtqIU/OoJnXs96PSiaGHN0xyhh0H
uTyBiu15KUay/ao5fb4pr6kMshyJwpI2VM1docc1dHvxwJBelvPgcml4QK7/0fW6NLcedp3jKwpL
TQY2GeNcGEYJQwGOk0VO0TaBSVCMuQDq2GJ9pXgtgsK+fM4S0r2YbmcIyW43fJjSAKEVBnNebxHi
A+t8ltJLPXdUrTpjdPGmFi2R9g9Lq3zr7X5cc8OGfqGdcM69XpnXO6/p32LdkzO/q6zkXh1hJ4AU
K5EUJTHnht8Rl8apnzTCcsvjR6nyh2+ehQJFvYIgcusdDgatHLFPMv81w+mNe7RdN4lcreQtiJlU
hH8RlRkauZD6MV+nSW9neEOB47eH+sqP2/7Gbnxe9Eb3DD1Wunwxb/UANjYfh/znym7PVOq7FqBB
VbGZixnPkX+qZhNE6HWzBIdSsWQKopr7WGgAB9qhT6B1FIA/6whBIAiXdi6UnXviTI38iCIKrP8E
QkWqN18Vo+s4jMGkB6fEbgLyrWq69arcPURyXqXqBFLNLHUGPVEZZYWly5lELAcHrFNhXPo9xIe6
cCClSZjyLacRnj7xoum23xgMX3IfQyWvIBjhlzyxwORfNiszX6rJbf+nXkDpEwRo2PE4a6Qg96M1
xlVd8Nrpmkd2AVxhYR42KOinq6agLnwwuu/JxZq/nx2F5ZrkiIwRDxiJVC+Hj7s2w27HhetBSy69
pcQzPUn3rnQ+PcFzzKjgeVxbsyRUwiAFvrWkZIEoWOpT+iBnA2tgnuaaKdNbH4vHAX7buvCPL/jx
R2uSOEyY98QLGRxmkO7C3kzYQbeMlY6x2JlStZr+2jmA2mVyPeFNKLh1fM5+XCRrZo5dY/b0PvNC
dssd5bUD3aOBBzchgnYO6QXxazJygu1vuSdyLfpleYt1wcZ1jmh++6ygnhJhHTz0YM+yhZJJeO9h
2njlFetN1RzVLThKXENn1ZegIacTUZ96BNFWJjjhZ4Q6glRgse7LjxNTU/W8iXZvdoAxbIrL1fki
17x3sVTQoASadz5Vkopn3QccEWriSGCn9O7b2W684fAg5ILCYaxOmv5XryVL8W67R658XOa4kJhr
qXTvewPyw9yhLFEHphmrFUJ1Isd2gSLuYNXD6am1QkmNWTutGgOvCF4yjRz6FdK4ukTh+4WlsqGn
Yi7FwXTpxOk17TQ3J+jQgAgT+JfXwwWCiEDoxpyQtPTjBtXMR7b21js7r4+rVIYjAS/SKZr+Jq3e
OQaqqJ+QSZnXtoQr+cGhAhgnBZnFEuBuF1xQHzAxFom3JKVARRqzFk4FaXqBGJp6Vte1pXEhZkJF
nG60Ssi49xohdBaVUBjNqhzv0He0DdYrxuyou+mNUodgifQDXeBwBu0NM4w+7fSPM3J/pvVwYLym
iN1HNFO8KfsZgKy8BdNPj+440K3QDniWWtT2CVVNfwZb7FmBAF02Jwr7UBY2bZSxtSTsbUyBXYfz
qp0X/6nBi8XUfThzn9hpYTqeGXv1QtvpXUuo29eK5Rm16U7wVnoeFyQiO6pqvqunBMaGz+s1G4g4
juPTN62+uF/VU0/LI9/gUC9oLKycKuiZAQqmUngAbvU4q7YCiCtIhTu5A942HwPROGa+rLJfL/H2
12H+By4SZI0faevqCIc3oer2tzbvLSx4KawNdZAfmy4Wp5ORGcM9rn02SBhmzAyN6tdZMrb7cql8
WxmroTSrfJeoKZ3OIGYENDqdoDcpB4CGDIA7gJB06yU+Oey6wDfNikEER63+BnFjKoatrH5ulmU8
3LxhS8XiDO6xYBLQiTZIM0aaaf8v5a4KyhWYQgoQ06HkTq7ubAWRWbnkWv6daBBMBaj43/F0vkR/
+fgdND5d35P7gUekvUzPfvzXYqWCcZ88J2nuztsbNjH3Pw7q0fZAPkU7oPCL5Xsfq/5OJBqIQboi
S4GIOlBOy6yCBHLDersgSLIVNsJGpAMwBKzdeAZ/oHtz+Xv5Q7Mlv2aZYQfSjzOlSx87PmyEp8Wf
EgNG8snC/fLLO4DWB8o9Hv2CF9V8VpEACPx6casu0u6LAtGpTowI/rkAqJgyWLOrSPRrMaA/6ZSr
z8cnR0QVvFJqL4PRt7x2kCIvqbfKh4M8Rx/GOpyCMzQOJDB9hmwK/QiwpU5G+zYz5WMpClZATF2M
rYM5ccU4Tk98ds8wZXiskBSAVZoSgRHSYKcVBH64FpdRhGmUiRitJ8a+1kvuLSKsEkOi+LKiHT4x
ulqlpEU30970enfmrdpapYD1Kkf/mVhzJiGifvLUfE6reG+pYn69LziUeKCqbG+66imDviXBsbtg
Af0h/a8G3vYADZgxeWrpAGs5RmMasdPg2to7VcrtHVUH37ENnfciroDCv2JCj66h+Jov71LZ1p5U
KWjoJJXASW+8F9slTtN2h4y5I05P5ziGUon/jgr4Wf1pawxGVkU0sP2T2rwwHrFyf094AgsQmKhD
8rad8P8N3ujsVCZpvbY98/UO84d9pO+iV01lbJyim/G36FwKH648ZeKeO7027XOHG1poQzUVgBPq
XAE+jC5F9eLAWqIG0K5yYWLvX16pXLlkiSPWzu8CWfLWjl5UVn/5jOzeZgjd8sb/JmlfI0SSEYko
giTl8VXv/H25cBmsVN6fqo0yxOwwKjL6GJQOaCXz6esi/ANLd2WHgabqkVFmziUKpKzxTPmpblvV
zTSYYeZVrVbdWQDP4X/ejM9D+U91idv9dHy+mbATHO7PHwt05IL7+5jDJoZQqY9/DgavHWGLbKJp
RJttXjA6d6UtinTEg9kN5MC/2lC9c1Xdrx4gXXRvYSBJ0LfiuYpj5zSEqFT4W7wyIhuZGqntDkN5
L2g98gsAtT6ecU3YGtw7kiV0N0+gKoUrhiSF33gWJeHXSnQ4c78kkVM/67SyM9f3BEX7uSmkr2U7
JFLU4DHJer2Gtwj89tSJIBRi4TL+SAJz/Y+tEQhNg2Ur51xhx1Grqa1cY3Ds/PzqOe3YWrJznU6e
Q3+O76wAVpLZkmnc1nY5aQ70oOfU323vg5tLjYgj42WPw8cAKl/CKypGXz45RpNKwjWzYMu+WQ//
77I+7v1JDzOZpaTKU7tYFJVxhkaILEwY7ngG5QUOCkqUseJnbCmjoti8dL0ZBCjBcTQnnc1qc9EQ
r+vMVsEefThULC+XCh/M/CeIHrsOq/GzDlmswfYuwgP73wOUXUuD4sDYqmk/MvyWn6ytYRUG57yG
lU4tNyG/7kKqHsrDKt5FPYzqN1DRfYEmUuo9CiqHzO6h94pMkgJ8xd7OfDh9JoU4geqP7E9dLpmL
/dLr6mGEV8ukt97ZgtUVUIEioz4J/hZw1gOrIp8haTlXwiIkoHJPf3gtmLuh2Fl5nZ7+US4kBaba
smY6Sa4qxru/fH3/+HyLH1HVkosboUMYOk8hod2BwkaRseaWHUcvSJ37P9viuzfvcJs/oSrECWWL
wbIlf20WfNT1zUEp6sm7FueSTtyTeIX/fUnsnFojBpK9nrtDtKOlwshR6PDQjIiY9jFoGfr3P8bR
9PKz3mwCA40ZfoahZCwSwDTyDnCmb3rQFqPv1rB4dD12zBast63BSin1aTFsq1U6+Zss/eLubzpB
McnSwC+yrWwrg2K5/mNTwU2vE4S+NLa0uDCagn+otywVZgWSTb0gG31g2yK+GxOIOtRR+7fO7pvo
7jK/TbsPHVLjpm8zEppEagc1z5qwftZd08EJA+BPh5t4p/PLwoT9o81kS2xEM5KPgo0iW9A/y5E/
nwGZcN/qL0CoD/Df9m0onf1i525xkwTae6uww7c6NxPsTanshmTK9C3PlgMkKGvZm3EDjB3eFEwd
jh8snKLW6YSsBBaavseLUMvcPiwMoq80ezYcfL1CARy2cUMmALi52h5l1MzhWwR0fVSviHBN4TDh
rwT9vTFgW7lyDmFQ/qnPAGQAu+oAPymLgTn6rSOsGURrXcR9Nk2xuMHAMdGmYsLQ8Kos4b59nBKs
QPqCWXBi69EOcr3zBoskJbJLwanpXWUOEhFQOrYKk202DWIZDNMELJOuuF+xW019Hwc74SpmMKkG
3TcMUVXkRPenAArq2El+wAy8ccEk2Ity+QzHQ2sstwBmChOROnXj/O1PlykQBuD8sSI09Bf63W4L
r9qQaC6Be/IMcrbjzgYyyLpy4syKtIX1PGzuxTaiU7OwhAaL73AXZ4wXqRELqLwXIb5NwQCOC+Ll
8C2qfJLGbS7bdKpRYrMn7dDgoZG5XhtCCAb9M6RFYU/OgsSvPxbmwBaGLwQlvuCCNWc1797VeSWO
hsohW8Yp5nFKpD8qC3OOLdIYFucLOCrPNjdGHgmNGeljdM9BKfIYUXP19rfbYlWeicqK7bUDI6a8
Z6OC+pu6tRn+mOBC2C1tDkKL2CiL5bDj8wq8HTu5Ws5ES8QF7P7e+O+UPF7lFIz6M/i08xgOd4Ne
7VXwaHXbTt12jqL2hxkb9tYmfeZtfo894Mnkfo3VG7LVxUPxOY8JoVGRxyEaeTKwTlHd67U5N7ik
dttTLGo8lQV0HqeBh+Uw1l05+4comZUqPAC/jao3J5ZZXj83kHnf3RVIttGKLsI+CSnBinpOSsE7
h2zq/cfCkduPL3eVPP4EnL2bvLBEwqzvdlEevAof95P6fQU3cwCmqhk1iAlWGi+CCjNZEbnYNrBQ
flZhNNCsu/6+BiXt/kCI+uThH10F23+pBvp7TN8M7IjLl7bfdgXOR0U7t6SNS0bU5IogwxBnFXWk
la/y6PM5e/eXXXwhJvs8M8MwDygpYdMHHM/nfTZZLqt+gdCdFgo2Wsc2KAg2SCXQhoqd2gxGcUu7
Oi9kYbnZC6taVG995YzBnj4K2WvTdRQXMH0Jye6Wos0bGc7gX1RWYCTQxo/ajiJW1c/llCILKDTy
vwR65xfVtJXwJmbX84RU9XZsdKDYgjXVmOC+YPzjf0fjWowFLgq9Oza8KNLsNqPec6vRizWAr8lH
aR6cp1yoIRF/ByFuCYM5/X50RtRSVzJzkeMZN96O1ZAU+kqxWrwiFAyJZkQzSDuKQUhPPXgV8SGO
X9CeFGBLngpxYqrP/4b9J6F3OpdkUFcQ8CGVrMain7oGctlpUyqNiCihSBoA/aL/XrBv2OUgPJoA
G3iZY6URfx+K+qTqoufu5jL+0bEA+0Grxmdcv9zfJXJ5P9AbF+ZDgKq15qFPxYYLtfjyxY7Q2COL
4zU3Q/kWClG4OGYB3GABW/m0yWPlV1gEoR0x9kdEFWSEapXpDEL2IpsfFdMiLPBD4pr9qXk84j4L
yMomFeCs5kVid3Kkv4oU1ZquOXO9GdtEq0bm/5nqfNkTC0+nk+NUgFcLQbtn3rmYRIgezsDIzpkv
SsM6RBCE++CunISptBMZE8Q3EFUK2xL2Q+TdV0U3P8y2rJWhjnxPYNeap3Q5o+FSd/SQLY2R3I2t
cQZOJpNXfMSpM1p6PA66j7hLrpQTPJB1wduvRmEhvA3+U5BipLGwspF0ywncx+aDG/ATSpWcnu+z
ZzI8dS/qXVznGw0PAuWVe4AWzdcDvFnE1kyY/WcpNnkxt2D/P9mr7CSHnXWNoV95ETRyVK/fWUj9
cL+mDLWwbZoLW6pQ3vdJvNVufTFVpETk0H2gpgNKrhUPt23hH1CAMbpP3vk4iLhnPf6QHPxWoYS9
8naUZpMog8d9wV6S/b2kFiLWCWfHhYE0NEek3cJhwj2zuABto0+XvtVQ6mT6IX17QuJpwMMrLIAi
/3eXIOHpRPMqfJBw7fPiMuScfpE+yUHQdcoQ5tg/7m3Bo+4LpHXfSrx3ij7fUaV6OC0lC9f9AmoX
IYoFKbfiNnLvf3GdpbhkFFOp+e6+BWE78WZHJnrwKyNcRr0egwNv0xvadkJyf2HGIUiYDAeMk+vU
6TIgGX7K/rnNbEO63I7dgtkY7g1UqzLIICsKpfMYQtGe/rkL3YkNUV3oRAP3PWo+6cTnDwgcrUm9
xh8VhuDwdiC5H44lvETivpz83afQaWn8ujl8YIon1oWzgY55A6YMqs6f+w55AfeLzUiMpelQPgG8
7iMEFW1sLFlwo9Sm0rVTIBUE/OLPXFxdaBnSFzQMokG/GqnK3+LmmQOBbiT7s7sQ1bm80JkMUvZK
Pkf6vXXt1cY4AclFKu4HNs5aIhHIPV59TW1Td93nIHH68rCQ+3jT+NFoxQsGqu70P5fqgmTEWYTv
eYAveUHSrnnv0ZukOVETNVN3j43QpCiAafmg2opywLixiq0GjkC/VxW7IfK/cpa+NAvUTeIDJWXX
1Roy1IJiJGO9r/dNOXIzBk8HdHv6bjGZz1SPTo8KZ2S9Q49q9K/dnSog6rYBnLglyGgz8xOxzJ3z
F2aKEnvPmZatRJLYx9JyUX6RRzYF5BZd6XinsvyaG1EvA0Rizehp0nz7lkSQVlWxOKtqpMePfvqY
wt3p4ASIL1ItXZ5ijBKCReCbQp6/k+KPOulYsrKbShT5offQdnIdEtrQj9SOzMny+SaZFgMtxBWf
clrERQoNZiopyAPhP9Xshs217kHRkxmifJGpK2hN4L4xQu8jbrDnFZhiM6315rh7PUW66Bw9o/AK
0/3DX2ueBvT0jJkRani7k0wDDAig+Hw+2YKGCGkENMSmw4qmXwsqyjbjn4E/QDGuffR8C9JZJ5R6
BM6J25ZEx2eLQKtUwnZ2EsBdbjqIHf1U64wku81HHCfsldY1E9PzuGEkfhxtS+epWgFH77ERG4um
zquAo211H7bSCKIuh6+VLCtgMXXHdNwgN0lAVeJaeBdCQIDiAsieMH/WHe89/numyHpz7M01L0KF
k8FRJ8nJFPH+09bBILv+thRud8ZI3+vvPbcYdkvn7XG3ARjHG/PvhVMe0t99uQ/YAJck/8RZ69QW
+q+MlKIEPTGrqXZDd0bi+qISCOp8IxKaJ+HyzVtQrTkG4Khsex2CohQZB9XnQ6vqj3Fox+slp6r0
LWukqexKfzl6PE9iC8s9Sj5Er0S3ZTT//4h/ydUphvjPwSyaKu9Yb8hHHtCoU9XII2dEdOLy6jRD
hfptWXv6druM1vD4qGrtiJQ3yrJ83Cvdt0TzTTrjePjedeba7yLkOeGwQmf8VKyY40CF+MygBzaW
AEvCqoWhgYr1QsAiAM5woKJmceNVbTha2BAvcMRLjcB4DLcbwdmK1w2TESL+T9YOWLYDxf5pUWUZ
zowb51sT4NM485giPq3mFyH7eihout5GXOPRvHUiGZPJBrSU+zTtCjJnL9knzTHnftBZrStibP0I
NsuAFLISP9MFDMw8NvPRxR3p4JPK+HV6mS9LIU9HktUFK8/gwtFeFQH61dA6q3O5kxC1tWaJI5kR
PJfMb+AnW8sKDB0naHbpzL8tdxO62Yf97KBTndKeY1cS7tGsfmtZSMe9GNPiV9SzXFtTa5q7HuiH
jDBBQG1Q3pFx74RlJDPEt2wRoO4nN65yh80CZOS/N5I/tfGTyJEJPEQvrikqPldVi3djES7R2aPx
Yh5oRTcb9QPaHtaCJuE2GVMYMp9EOCQk2przXtjWA8vuz0YymnxNDKKGOWcvVwq9spbC0lX+Nrgo
ZJloyAyIlaxBPe4igWNqI3DthGKbBd/mmnBuXAz9TY11q35garX3RyG6jc1LHknvo4da5sn32gz8
oMHRJkNQSsHjyDz5GaMNcMU9iXyqkocS5xP+VzbT7sivYj8q024ZE2P1El4Jm/HI55CSP6WQZs6B
KMIl3LAGzmRO+9sh2OwHI8XIiz6L+SIjb4Cp8+VLvzTiwVACJznffFgnr7thvfZNGKXPRdG2+G5H
XfE4EMcXyKFP62bxMCmDJRY+o/Ap7IOHxpohy+ckuxS2MNTaTiNlsv9W8jj+N1D5wIHuf84MXWs6
2f/mUMOTyiNtC4aqYt3TdZ/gTpu8MOHmzT9I3B2cZ5zg6+jEypEC9xQ1hjyRgLCGe80Urjm0ZWEQ
O9M2bECfxPF0VRD/5c5QojD8uE0fg2sfB7LkQx91a8Hc6NYPJEgd+t6LXuDsLhHOGwe3AJqdTbTk
fgUucVP6CEaxt0Emd3UuuTkXkyuXHm2Y/tz+C7CV2XcvoqYDWS0K03RzNbX0+xCQRDh1UrCB8W/v
lc3swXz/e1UtyIMV+UzLaycgxh5J02AboGnX6AJx3KQTT3OyJTSkuCHHHtLv1T+W5IdHCYBf+6eG
1YcxtOOD8FvlZ7pI3XXwz+75+uD8uZGe0V1lyExHiAFcmZjqGV4uHpaYGdsODWQq/8NiaPohmA/3
JkSDo1/6D6fvp2iPnLMG4lxpHtAmx9L2RUeEvSojS65g5tffHpnmMwzpowNgBlfQLUHdgwpGN2Bj
0Go7Zt1z+JSYi68qrKy2i+cUvFxC9QqQsHQDPT5Lfc2q9ZFmEgETLAy4pYg0Ex2OoZoStYTx+f1T
1vvGddHZBW2MPNY8IDghmVmpc/qpTRzCsBhMfURyF9ifH9vkuxAq0WJc55lSFzgGGXG6fb2z5Vb9
ZSyYhS482SnBpiGslQtGC1bjAjaBkT8gEtWka5bS8JaRTQYb0LvjmyV2nk8aZNLsRyERLbk+54hu
774pYhYb8ugmbNPF0TNc0zOt6isRYMMePv0tr+q0EeqoFKlvrKbB8mc9Bcj1+4lrNC1MOYpE3LVb
up3lTYjieHOfankh68R3M3Tz0RSzEYheO/TAJ5qdmuMkDOalKxYbN6wIUFjBn5CtU2kPUhvhitaT
5kQTmk4+4Gdex1itdg5z7/cIq02qLimVu1PHcIT59kHipGLOnCsP+0EGT1OoACIadSXAR6FP2O3a
ijUVz6TJnjJnqIXeuMNqT/Ep90Wqd2u/U5x/OimMJQ1PS0jW/IBxg98I0M+FFIEDIo2c60tz6ZTU
gyIXq3dFjBwmyJdnZ9VqtzbsT4iS+xX2/l7DqEa0KzuXVtZomtl7ekBm5AvFGslcnj96TYdGBFY1
gOEVVAF56rrLwcONWEGPSNGfYa73cui8mspYs3KGpSkU8KSq1FvMXKl0rS9/Z9l5RSf5P9p967w7
xB4UhmrWKnXTUmQEALO911CEmZXedIqYyMcyX0594Ze+7daTXKlzSYdtl9LoOc8OXqqWJgOAyCQg
Zodsy7RaVzY6SUQFEj1HCoh4uG6b0OgfQN3gFiS33nfOpKgIF9mnn31Mi9PRciJogkMh+K371e15
z6L74nmjY76IsIMgmzGLP0bJo/fohcxV7EqLvw3UlBQKcCwck1vtBiMNVpzaHmU8Z/Xt3v4Vhc81
zWDz2iph7viAjP4l8qbV1P5C56Uq9wSYB3oAPznPVyfUGtLncxGTwWCeCEuvUk/HhMh8hiqZvZIH
kNsJoTK2FG745piSZNZIS8t0Gu3W49QzB/12f0+HimjgJACWcl+pNvyKLwIC4wXFoCHZ6sMGNVuk
yK2Ki+WRSzVyAsfvdy92SCEccMBY5fwufUWMdtip6iq2BpblEnnPeOAi2PYxj283S5pKaLUD6/Sv
pLs3nAU7sx3sS5EmFrqDu9ZqiMsOR0DkFi0np/QZYK3WJxC9GWeq387SRwMjGCxvpIN+Chrfpx0R
K+DtdRLUdm2FpRfF0y4HY/69QID5QtC09zWfU7OgfCZ74nRdAKgjBwODbulkG+9WeNzDD+OHRQ6z
X3z7wWZ1CCtIEH969GLv4Rk2iWynVLxbwLF+c4GzmMsLf45IwTOcwjRok+/wZHU+hfC/F2P5y12A
UFL6Mjgogigeqnhg9BKw/s9xs/ZOT49HOUr2JnjTIIewwM7ARdrG9h0Tk1ovU63tL/UDOME14Qz2
sPIF9ax5FsPcTY1cAG8ib2P6M8WQx78w7hp1q68QoLVPA3pemY/wnfKv75uckmGEwR4C1MH2LxLM
rnqBT1xGxDNhZ/xjDya/VDYg+DJjSTmKt4R23fQ0OBjGPaAxhwol72hqxqNiBy24JCRzyk6CYfjM
LgQkg/WZC9pY/N0B1rK7E7sWyrMr9RaxQ8ryZMd+FgQtfkDQ/UwkzDNZEJXGUKxXrSfsVXKoqTw6
lqsALQpalc7MAXrmgUxu0bLh0RryGyCtf7Tjyx7UO+eq/YSvcU+RiYvocWRsq9OL7ESrP1HoNKoz
XNwP+vUtY1PUcXfnR8tC0TxQ7bX+DbkAFndtTG9V3/VKdSrscQHySy8MOFYV4+/xtxHiDR+SiqU6
xFiq0TZiMqfpxDyI14y1V2aSgwzPDlFRBHTIJ5WrS7xf7B5QPLxnrz0fKxMbS49IWRIkXf3jN5oe
DhNVAxFt+LSd+gU7eXO5uftozxwSgCogo1W1D+y9o8paQlx7rDCyfOs0HcswokYdTSxvn7VK52Zc
CKjujq1REcB9wCDZI+l9mlegUc79W2tmFEp41MndGacWatZMq1c6QuP/ehsdIW/BXUSD6evjCk13
xDCmwtjO8k8ypJkc2mNo38JD/sT71ah+uhuUDOmR8GAZhqjCYJOo30JfAw0WUCFCQExZa7q+FWac
dvnTZNO98wKeXHDzk/k9JTYmg7G+C//8Pymd6u0dG5Ff5BPPGnWfxxMQCyW6/txgXzs6rAB5pCEZ
g4iZ6i/OhEPiHQ5srE43KSbWUNzqR8RuthwBVzYXd0UmT9JrZ8R8fZsMtho4+4C63XRbGuB7U92s
NtNKWthqTWdzqDwz2oqbVLyRnySMH3WubLcUkpWd+DPyptmTejqglwA09dxCWiipXJEbuiz9lgDo
gNylhY96LTAwTaxH3+k76CG2p7IjQSWfEw2cZJseUXrmWTkMTDaPQHVmxlR4LHfcbkSCU6RYRnPc
11j4cgIaq8Kn02RzeCUfpV7VngEDLFjDCJNpJtHvQfZFOADeIyOwT6n6AV5LZjCHHatI7M5pnqqj
nN4G5VoX72aIr9VdFrg39HMMOW6dtdTAUW8A74pTqp8AGnmVk8UeEozhlJHQskuKol1SIxQr3cPh
O0HRSaVQE0jc/jKQR6wjhLFJVdF7iBo0j+mBXzcyCW+WhiCPXbcMgWmkbWEsLnnjw3GN1k1DURh7
2RECCPcP1bev+HH3+kcl0vZ6zL5XmuEzAPcpbFsBtA/QZgd0fNP+4Jxo3zV6veySxlcuCtxfRdya
oLw6ed64JHA75PalLbWWYGFmKCTHuMMo/5WSDM4cDvydWShrLyQplssl2jjz1dS76t6HH44fcE/N
w8YmR8fvW+yPXnl71lm1efddsjYYOqkTKzsEyEBLuR8HapohZOu2SrHgQu6B08vtQZUozeTcsaJ7
JPYBk1i+gP6O/G54M9W1Z711C2fxsL/OT+1eOKyb+lOKahA39OZLQGCc8DYrYQGG0trpp1Kf08lL
i704kN+HAZNFKb2eChaaO5sB0OlxiKwnXAfQjkGQAYuxwR+VXRsujOGGFi9hZGnFQveMJJ3KpMyd
N0ZLnkxyKYtwtGMyo9HMlHNWPvNOoFmhBaZKfQoI/DnDQg/3miJAv7jhGkSMASwdWKnyN8y7U8cm
cnPO3ggqwyh1GRFMUz3A8KpbOCQ8QZTeednB4HrOuqGXsrshmaSxOpC0yO3vm+R0EASQ1uOevWMU
5hvhhqE24T5PQivZ6oy5qR+wEC9MWPVOQbpSlnSWGReEqCQ+5+CkaXdMAsjDW4XIqghvlA8/aMCe
eT802FWx65IwTiI5N71KZJfb1W+qeQCax/FDojV5X8sYOVQx/QAsu5bN8iR6GHqNgU/q5tGgb24m
ZPRxsVmX6pCGJwsoXXUQwP7a7ZFmNCkXu/WZ5oztQkOmNFggHW6vIN4pV5lfZErD2rw9SZEjk3uj
+dmFmuYjbfKiBMP5nD4VG9r4L3sQZMLbl9QQ6BVtOtHm/JnDwiqDSKux8JE=
`protect end_protected

