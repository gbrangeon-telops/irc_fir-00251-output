

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ksr82/EJdyTi/ZnocplaChIHl5gVfg/QywOs6WHQUUTVobYB9S2t7HfNHkvfksORtftr4wgSGG59
dqflxrTk9g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qqej7lC/8l20xFx7bklclhPhbKpE2SoVMnU8o5jHyjJozBFHGWWzSqcy2OHoxuRC4svtWcuXPZER
AveySsBsquyvS3CpwUhQC4HU879mrvq1rktu6YiGUKekxqqq8XWVjGU2RErpRUag/ydvNbNrFWxX
vuxu46YvGNDVpOq465c=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
439mpd6b2KugK1Dxw8VAcq35Q01RTqPVrzIbAJdjxQbya32eEZ7i4WNiFuVZ/MAk52bZBtBQiNHc
mNfbIfQciIHmnAXJEN9w/4VODhRIcUMrMjQwAjn4teKfB1tg762rR2jvGQ50Ai1Ml+OYADsAGJtF
URFceTs0yqpLMxJ8Ov/lGmeNw5dXmLiwn/XRqtS/K35VTjZyDUeHpQAr9q51KY6k59LrSFC7lxxB
mXX0In+fzXXlrh0dFFwLWzscDXHiKjrU4bwWBuzmrkKr3uCoEG0OADwjka6wlXo/Z2cEkTpiK1Qy
MmZH9UXQxrxTgtpOMmK0pjs+MfXf5/7XzeJsOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
porEUqarzWQ+a43o1KcgcLOOq13cwiYUyYcVmnYhbdWCiVlWWfN80U7oRzW3NODV8vTOFdEeX0/T
HiPsKQYOSEqQjf71FVXt5Qu85a7gangJ+zMjyuk8+m1c85rFqWapoLbPUbexfLeiEmybpwcybBzj
rIVwXl1qRv1R4JNRI44=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s6/C7NZuQyYs48nVSWrZBvdUw/cGGwVNCnxc6+Wr+hB+GSdh07xJnxht3+mpM71wbe2jyi3JRq7M
A8Qq9KlqvpjZ87ZnAxTvr8P4OZV0DRnim60u79JqHUDowRtwBKuWK+fhBBqVkg+I/GuK0CQAje2N
3H5CzXagxYQGmhNBvdIDYAmWiG6ymENT9OP+fdf/JngSq3sbaQDhuOCrSGCgAWuZWv28vEMvXd4d
VKm66HgH4TXtJpDsYN5kTW6gEWdi7cV3KJRDsY6jA9RzwyOOBsMl8Gl/UvSGBWbIshxBeydyVUyg
0jabYqp6ODPXSowz5ZkW1y4reTS+cozycJAuMQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11008)
`protect data_block
J8tIxxVhzfnTuE6Zdfx1q7GetP2y07WsjkPvwbzT/XmKDLJFjrIyIU6cZWL/ljE2/oxjfsTeeGek
kQYuCwe7gG/wIAnh0x/dUSn/k73AtUaDs5CmGBlNpgM3XLluDWcDCXfshn1pprI7ly6AWn6Q4bTI
pcR/L8CTEiss6F1UNAkPF+b2JJkVQUvgu3wfWeuHD0IiKBL8/STmmNlIXQS9OKGbOhvogeLN+fVP
BdfLr672sdLFpOfmWp3jgV8OlJVOJObmW787vQJydfQhed7Gq9KI8KHileBgXX3BkdTElgajiy+I
aAhhhkV7ngMix/2AvMJG0iJASloGEG6zh7X9o6gJHwLtIt8qatvFjOJzn4i63cPp1tOIn6KQ0nTo
PZ2kFUWUm2h3XQTQaQTbpROpLeyZs7QhXZH7KqlU3H7Xs1LoKgAsrYJe5hmMo8Ycm6EZQUnwZC2p
NyBJTXo8oSUFRE8gVrCXMb7gBGyg+jnztLRPGEqazGBCrykXWirqtW3a+t5AZxVaLVaALCgZTI6c
6n1xFKWy0wbrzQsaFue3D+MjYyi57Lu1rjboBwoeDhFfoc7Ct0RQdKECyYHRxBiulcT8CJxKJxsY
gqnEq1sKjZWpPIjt4rwZf//bqNS5FdMYoaO8doTkf7uBYRysvBWUdZgSZZRIIL73pIvuiR7q2Rqy
U8mnFKCRglv5Oi+NoYLMocksLBMWIRjbnMh9CvAVhrQQB1efWxfkjpGDZ1O0W27j4mcM4xl1FgtW
QJbIGf3jZ2+QrqeVzOcWXkMMoWGpKUIcRwb9ep8t60oZgvTpcT7AkMOfnNgozhVvrwtzxxRLiyhC
uoI5VkX0eyY48qZMWBDCejpj/Q4XPt0qJ60bcobCPrlhkti5YBS+XzjmCfCdxUpIgt8+b6Z5x4VY
DuA6enmXNw+KGZpokrPgHktxkEtvBSggJB8hSLd7e95H85OjyZ+IKlZmW5fC6tGTcuyyvIWvt4yE
uK1+Dezhzoxr63xfqyVvw5nWrq2hsNiwR97P+rLDI12IrBmQ0dJdvofkUsXbEbf22iFDCxAVNwtt
PMQiwKjLeYrXNy5urA691fZNlj8+vR1tOp5TxtYPIRtwKF2SykeXP7BkGvaIAXH0ONckNL/dh6yS
+xbPC978TSzh9G1obqq6fZN2VcbMVgtZdhAXNLuUue/OqP96leYs3nNfO6Tg3aa1gPg6TQnYa+Y/
q2bjFRrW7mkvEBTVocfgS4iSEqS7f8CJqQJDbkk8Zd7GQhacMbkfheFpnLGJG8D/NwCKUbVkrJOM
Sj6SNr86yI2FKgpH/QMUnHNf+ivkL/SELwkjXBCeJ9asYuDZF7POqyMoQ7D1O+k9NWgfQ7rxeo3u
+lKAzet2coi/LLZRN4IYtBO5UR9tcKdNrqSsklmpp7LNjdZBbGIlDqkVpGz0I7saTMzKBT0Z+ERz
koCdyZCtc8UfXNFo08m79O/XkK+1hIe9uJ7u98z+X5fkZiWlbIFzUKOQtC4xrOYsfZos/spgBmrp
xWRaenJgpS7ARdAACCYmzluYETpLBwoxlb+T/ICIv99aUrcLNGyWQ0ES3VEaT9DzbWFnSyZJmEOl
5PkjXbq37Hof3O83gQ6+L5dqu509Eqe7mLqpJIfN1KxWzoWxbyx1igo6Kzm7U24zP97oq0N520sp
OoVWyHtCGqKJaYYawDpz1LhobwqGUxsa8lJxeIr6f06pSDALuq5ouSGCL2iA19ZVqpUJy6qh0vb8
w86JJTi9MevaSBsT1gT0AyJfwZhN5vB5vHDYMFpxL/r9foZhjTmrZvodvw6XC2JHEGv8wYo+74B6
10h2HGJ2iQJHVVE470EwnazqFFkr1+ILWQyvNWLr6txMyC1EeRJ9UgrDiLi/wh2D1FbKvKaegIWm
Q4ng9YEP9mlymaYhYa5N12Zpo5gmIs7pQeQngUHWCc7EuXVmbeW6/44j6qnew1uqSN1k/9V2Whh7
TlKzO+Y6usHy1+ueIdfSlVNkjZR1uFE9di/5tRipRkQM4b1UMc39EK70xCjskSltKw5yoSIYQidG
bwv8OzR3/HZto3vtqpqbUaNNm/QaSKQEL0anuY8eQGcHXXavZL2IAR1L09KQsIyfcu6UBh6D1qcU
8qZCoJCDn9kbMsIm2Ic/UPU3MBlmN92rdebpi9Dcnwns10sNzRkzcWiGS5aak61t8UPsd5ZqIFm8
73PAje5zCjvuyhMK8wDwYWvL+9x0lRguSy6vhgTj3dmmL5q08sPTh/7u67t7wzVHNoQ/LaemN6oL
gD47215V1HDlSnRp/qBOvP1ODNOqx78AchiAkTuq1bbxgV8t6EdzdWiB7KHws2oGqKrTkqNNnlEL
2S+NdhNb7bGIFVskQdfsGKCpK8DF+LKZnsz6gtxchH7RQdixT7GzaxFxsJGOjlX5ln90nWOBE7xw
49MukXgeKVII3N6RVREHxiHlRqjc4g1wgpjPkMJLw4TwpXzDihmNmG07b9/yRxlhqYKD0LiXMQoy
mx+WjCTGftUOCsBmXmz3bq8byAvWwOcCDPPpDi2d4W0LRPs5Uq5VZ6Pm6WIecJWDL0lFZ4glPlY5
gF3bZ3G2vmkG7k7O2Vpd4GwfbvU313AGVme9UNxMM6QbE8MT4KlDNIcIUrD00YUWP3HUPTsiYRbc
nDU7SJUjRhqjkpogiU+URPy6YuIRluWSmYduUehZGxhMyMCQ9oBj7ajbLAzCtOffDf0uSfG2GLOo
VdQISihSivRpoQxZR1Ohi/5ZTfGuqi7jXyG/tUJ8YSiD5fUys/qvUc/lgeDexD9ztfY1zWYXjroX
i7LP7seTI3wGgmJWrf/zxBCA8qIA4kHyAWrBZJ7lkk6uPHel1TpjdJrPoupWVrrw989zzqHf8WBY
hGhd3LjegymC0Hcm2WwuB4yJtxTN/C8Kh7yKLcY0mshqFnWQUuZvqYfhnRg8WzMx2oZW+pkVIZr9
RBMNYYnrkjRVAX5VinRJA+ISNjlgc6MWweCaGzxGpv/ZTUBjd0KZx14CZ3hrZCckAW/bhztFZp1N
GhSW1S1ZzNDRaJDDlzBnRA2KRCe/5BEuxI7sZ7jK82RIPdV+wX7BwnCCXhDY6+uHPjaHoA16Th80
9+64L/riRWb5swzrZcHcr5VLOLuoBBlg6osrw8H+NWP4brwSC34J1Ot33KOuoxdRmWGvI9XWq960
5X71/Z1YJdzWI1iuI66wgScGffuUCWDPeaW1A8p6+2I8SeNGHDVyZlXwgNojhzu4Cis+mn/L6CUL
TIjDPA0AZuDzjwJETA9TLRxazAK94oRTR526ju6hfReD8J6xBCqlFLFuaA7uaL92rWiYZOaJ9QLl
Uw9VXA3M2q6MFAMy7s79nJwRUXQy2KU0RjK9dbKpIl5BvVRI2giYhvGENsnzTZKVDFDVQWFg4Shq
6N/HhEri9NMGx36LMpf0pe5T37OAwM4iY36/ibLNTVoMnBDabQveTKYipRo4cUkyttHYWXIbJRvU
yUTnjJTXnu1pttSKNvnRqQekiGVDoYMzZMw6peiMdosn6KRYyLypJBdiYcukDQM2YGkpXE38bYq8
Ucj7JBkGU4zF0UD0QfOJoGUx6dQ26/7Lur9e3O0wQhvwFKl8h6kfevXVeNj/9tuds4fWVCAkCmW1
23qBRUh4hWfmJ6mbrRn4tdwurQayyW6OoxmcYgX8O+P64ufvigTGo8fRlthrbfWhq3Ex3DLxKdfm
U6FY+FAuKvb7im+TAVx7rhQ9j/9EThaKJLqM/AY0cJnpvdYqoIwekAVnFvdpShj6rfu+FRX/ceTL
Kdy2J8EQYmJsj7aaLMf33yWJ8HsEXYH8kDFVZKyjnThl6LuvW2yM6DOsQ3cX8T5EwMb2ABy8hoPI
WFyIfavBRt3my5Dvdr4TjcZ9TLYAO4C6ApNpsTJPbPf9RmZd8tVVaiM3RKLH6eHHXUzNz/3Llisb
Vqk9vWVk6i3a93CTZt75CeR3p7jkFiBn4gkkVXvxziinv5RD1w4VOSQKULxQHc1OQEUVC73aRLVT
Da6UjNP/HeTE4cLP/A4v8QcSEV1vDfsOQKXyaVqTHR74lLa2SPIb5Eiocx9Iv45XUjOnn7+mFADO
O99a7rXapGlLWBKMJa+dcp5nYrAyo0CkQ6WWvKizEIECOi/TkFxs3JoRtb16uVNFlrD/Ru8Eo9Uf
PrUQlVejL1Rv8qDHpPI3Fpk7gcesxwY96y6YIPDCdijEyRNdeSvIr/n1etjHkJ1U7XezP3Wgb2fC
f+DhEB72KSEKwAYjYafyfnUkcwoIORInWWe8uCauyJrbiNZjRe0ozVVcfW18GVzg9ahlLtYqDTN4
Jpsi2jyEs/JWRZURCzUZqx69dUOkRPNMBupuHc+cmz47824jUgNhxwdgvUj5U3NmGHjhzQr5Dwxd
tV+uZiVEtUj5PbfWDArzwj3bAzr+RtXILGiIC0KcFmYmlhCmXCk4szO/375e8d0PeBjytEgolDHj
maxKD7Gh5YLpk+gGlTllIWfMT3CwrRfURPf3baPhdgfZ1C0C5mGVHxOZwKVoQ1aDFIZbGlNhkABN
EugHyo4dWIpaIOQOPQexJXUv8uyNCpyuZRWNr5DcoJPVQllZIqZFPaDmbrtNad9hmYNQ8tZE9T5v
htSl9jb0LiNTrl4C4lApv6a2R2IJ0KDtvloCEZvMVpqnK4NrtppCJbBf/tutteDUbjm8CNi0f0RR
CkSg4MemjS2UEvXK3G8TsB2fsEAp+bbyXZAcWXRcF9HM6kK4BoAXCuOTS8URwsUSBnmr3bvMmzCp
TXbnwKPnGryo1l0+41fUgdcSDp16BtlVRomXYSDUPcP2SfP1+qeubd0oug2H/sDAKSVnBn9wNPE4
qQtbINbGoIcFDp9nzOoGqOafv8oqte8MXXo9gaUb3a9GnN438lyPUMFPLSaDnZ2kFdK25OzU/x17
/MerM4tMsCr+lHjjuqfaU6yHTFEZRhlzvMq8fGKEoXYtfW3+gUoPgaSIs/2VdLhESU+5pC5nyffU
lv3h2kwJABj3tVrfpt0qULxvx9zs3h9sF5abYEB6CSA9biXuBQF75GJqIdtDJQb1UzDhKOrtJPLX
xisibsiX/qlhsGa3q/27QAbF0TWYz+FO3Tciddwg2chw5u+cO/psCxCIaT4Uaynzj2UrMvPi/wYz
X2PbWK8o4qquvfgG0cL3fbo4dsObWwMJyq8Dk+xWk3vapZPz2EXNTf4SoAIqsxZnLOmSkXN6N/DQ
NIrHNRT0AsuOSNsuvI3f6919axh16UStnsxxNZF36dKgEmi1GLOlOcY78x08svGJc4De6iyJuwWd
XVRCowcKM+mK9OX6C+bEusNnZUR3876ofsF1fRsRK0SbmjkcJk5JO5+YAUY5wmfNeof3GOXUT0jq
zD+Io2hY7JsnIQPYHsVufTpNojptDHjAjCp5BCIyHvdAwemW2Laj6hsamoB1XOBX41kB0AjZnAVW
FWvBuJL1sjvJrYvu7iDGmHpR0kNPqiDv9YLyqJQeZ1F2WJo5jOibJ4m42vzWF74PMYb9Tv6gY8UG
EDlUrxdkdq71zP7b/WQXjdWc3I6gYsw2Jo5CwDOPNyCYU6aEn2YHjkY/88P+cKWRF3JKUci6J3Z4
XovZKxm7iBTuWypT1Xc3afnTZUtRcr3nE4sYfCm27kgrq61uaZN12GlwlbhqOCkDaNhTSch8uqlZ
zsxKq2ZM4BymnY4sQ0uOO5giypmxEQcq3SSz96x0q6NGo9tSzPSVMedDdKtZBeCBAcZ5ZAtm6Rhv
BlvBTzmStZ0Ah506K2Dh1ifpH19OPJNoDTzaUs00Nq93DomrjUScNtzZjCOYa2gU2GqNFJwdD4dE
aaoVESTr8nN83+kw8Th52GcN0FNsJwAAzjRCjrR9sZTFP+vHyWvtYFrulv7Xf7mjD9b3ssRwTpP4
geXRFDrlkbcIIpIqTOeK9+o5CtibbYhhpQS1aArTcwUyJuzZtVjj7YbrGlwEKuXapG196gfFRV/S
y+hq56mOxgiGZ92bMlexgK3IUZCIisyanr0d1YIdFzpveDd5S1hB8ijj8PR4UQ4lbXkSJfUPFVtg
EDFYvQcrZhNRT9mciRyXvbkP+rAtivuoLkP93nMUYJvjGkrT4US1WTgVIR029ysZyML5E7wvqdVN
ZScByJBXFDDRpdRebkuNsYQ8T/2Rs8/9Cvf7n+SLCLbWtgZpcu5Ei9YjOM9ddwsBO68mnRHJCgoW
PVpdTCvuivcL6phlBzoaVwItj+6VfQa0zADnWchwnAxd/rrWgcDHkMvxyGIhT9YbvBzjoSJyGJi/
KGnJh9Rb8eqJkrIxwYX4+n0I5PL38Hj3bRVnHSGorOKwG67YXKH5OOox0gcebnZq1Tj78yu+Dtk2
rtp8Bna4dr7zERebvbHvTI79CjsjtOW0NBEXkM7Il8TKrysmMlrzSA1CfO3R7Sr7YdnHoKhdTtpU
jqr3R1KMpAfaxU7c2QKDrNUlLmgcXUAf5IafMaNowZ+lEtXcZigjXBfnndnv/gFDwPbCxv9ZGPCr
TkCVAJ0YIO4jvPkDwTPygjtXd6RYVhJZjtx4Zsj/EYrfQBZeJYi2jrZoAmqKLH6zR01G9KLN6R52
Tiw+nkyuEv4KJKW1e2Q7Bc3jpMjkkIsKDvz3FK5ovEa/0uukSIeFIgek8QAsziSBBN+WfEHIIZ0E
+5OJGpiFSLw7VYu9XAsDW9I+jkywPyv6WvM1IWU+6JhlvNBawkD/70uyGWpRvqasFv8/QQsp+hfA
ad5E0eeTTr+zR5z0zIh1PG7IjgJDcMsFSd0EDkcR3EtrKv8HM/HxH0xr7LC0VIm8R92wFH6RtdRt
wNz4RC7CnyI6kO9OloeJmb7/ar8wVhZXQzQG/VMMWIeqJ4Wr9PPlrR6XMJYE8xLSeVE9rr9Fb8F0
z87N5nHowazCYNnN0VTiojB2Ih+pmtMMFTBNu3a/27ZuPz2+WjrOHvrTMFwWiKkYXQOcT7iUXU2+
ELi2Z70JVtVBQwTS/g7T0zOv34ElD2qh1MNHQY76qgGnkqfmN1N7l+51DLwrSVWtMzCfX5lKC8F8
eJ3eEoob5WvcwkerjRbiPd7RPRGX5UZ+e6uzPKRZExUDGszIff495wG8ctNdzxrsP9cBGWZPpe7u
qSiuvmgj3BVil5camcyGeskCrykDrEAXqjRwx1l5c4VMIJ0bi3wRYF41ihpnejtI5MmyZcHXfBmJ
W/yOzFU77EZgsbbnuyNpHQrqakM9XovSYHpYjQT4HKDQHWssoTtgjPCuql7U1WRhwnEfCSyR6Lmu
JSVa0xHM6EglbVyPtRpk1H6sE2TrqoEdfB1pvmXvd7r7wJ9TLYPi97HsNChdUmgTMjbPx/R2tBBL
xS7bOw29pKgMNESNpqLZs7Jpap9ZlPRVZzl/0tQt4EvG3tdG7MiTfe0eKcj5EW2qjVLqqSpkGBqo
kcoqT0s7oQwFjAumhPTX7T43nSbVc1mFwurs9qUK/H0lNmgeAktMKTmhR6NwyhMcXxHsHvO7j/0A
u7aY9BqKWtdrub2jVyKYbh2OWIT5opRw4rWJ0xTPLTQjsOTMGlyqOrhMG9hkm+0VeitACG+x9zyM
7qSsTXj6mV7lC/XbC7H0FDPzUUSlJ6+KFT37d50AoOFjbA9g04cDpCoAwF+/fDRT8lTFqyz3ejRY
i0TIqu80oBDDXtDoqLi/EVfjWIGrXqe54ajfjxZoF9mOYNkvfvvc9u6MM1Z8iQvNOCg93haiOIN2
bPMkY0Fv10lZwnIGebD49zg26w7rRdzwDcBoTU8G508DtTJQaqTCcgtSghM3K/p0ZWXXMV28/iu2
92n3HjJ/sWnvOVJcX0lwrQdrxSCuiU3r9pOTBMC2CpiUA/3IQg/uFYsH1+lJzJUvJveUkOoPc8FZ
hZ08VBQmohcfIJCmS19ClEDaK/TdVBQq+Ja1xSwH20Na77U8ejNLhSMZSSruLAwUuT0+yAyMkJJS
11s2/11Utm4ftn2aIuzwPXxElha77gOpUFCkV0t8MdUrXRTpOlhKXpj1Ukdlo33OgRis1xv+wtFE
zw7Q0tjvroPYrLJwj+FWDG3DoSO0DaoPHEWq4X492yrzHp8sQsGccJ+1OEpKp55fExRpu/eGn0MM
gyyhPdO1QZ8OUoeJBCZ7t8/a6zrYEMv41c/bd6f2rfxhMpM7uC7Jw8iuotAT5yDFAzttyuj4SZFy
jfFIK/421PvvlNylq0OYZvWT5VnsBIixVsH2WLGYdZwLLPBLK32ulStR/xM+FpFUakK600uoJpeL
nsbi6f3resfuOs2tOuQ+9Z9UyVnNLoDNyJujDlUXyo3t7IUmF4r4C31/+ckIel9NJGWaWvMrF11C
TWZ8OUItL9YcXNuPoIL+uR0WG7vlqeR9fBLIfTFfYJnF6hqqkRx8OZmHanrEgfIUITPI5BSz36Gg
Sq23OwYzRsY5RnKWbYU6RGodAzYDvwdQKR/gVBm7OAnqyzfdmr+v9o9cvqH9Xb3wkKwrbSa7dIgb
LdbDhLbf8e4ILttwZpO6+Lb3enrPIjMjJgw5Mk9rO33CAhIz7szpebip5bCUt1g6soE7XIjyKN2w
6qAzpwMh64tkEwzTjbAwAPiHmujCcHi8/K+kkQD2+p7Mvm1yObpwtesFeiqpJyw/n3elsR7Fg+qd
D0IqWTnMDerJsi7thGSUEEDuMaKV5uHs8VxoLl1vy1o7OOImihUgthoDW3+vYWvpW2hjALmvfxAC
N5iMUKL1+qnTC4dg0rM7AkicrUkudUQGnEeVkxeY+31vmRRW1rFa763HOjeMiZoxJ0AYTrFR3d1c
nME/WY25/qfS/c1J5P7huxbc68v1lMz9M73BH0YIYy6tQW8kXYpW8n1FTSOF4IpQ+oVX9ryghUNm
ejTubbRVWiAhb7HXJ4B8rlOVCosyoI3xSvw/yT6GNUm36uL0aLlCp87OZWiQEJuztcrs0HjDrzo9
srCs/1vgs3VYFRCeBHsBFaIqExKqrGRv8tOSpgu/9XSfAMYKsj89NvAmlyZzaCbF4j/931hOv1wG
4Z2IOJvkrn3liStbJWPcYLFNA2b/8BDiCoTsdsUel7NTOXANH7H7Evw1uYXAafwKIOJaXgVh4OPp
u+6/L/uCKeGxqzP8r3D9uApL5qL1VikqeN30hrD0imGF/cqfb0kgIo9L+blMFdL39ogbq8lN47Fk
aXTXVxaQFa8Wl9lOclvb8N/kamuHFzkT7RC+/Mk3+E6jq/2Z340ZLT/g5cPpxtFSp/TdD3yUcOXg
vWHt+1K5l9G1zEfILVWMr9P9vr42pw5zNBafNI3of9deJVALgKsYpv3Yl1luZUM6pf1OB/V0JjI/
RX8LCOPG/OK41FQ/osE3RktN0L9b0DMi+RMkwWlXtZRvzRORSaF0GWJqpt698Z364IlTrxwxNip7
0oUo7wThALvyVgZ30Nn1bAlbxUCjVudnAaa4GYAUsRDV3CO85SpueD08QrADXRuPPSkBFvQvUjYV
bymFgZC5w6QPRta2ZX14M/7T5Rf4kJAmYVo3lA4wzpobOgHcBuwHqQndg1xPzhn1rJ/Y72jmatGB
590rAG7EuXgnYrbvvRW2HKdrEujGhIjlWSq5dIMbNU1c71eu+81euTJA7JO98F14ugcNNIZUG1ak
9S+AEECTD0FaczFbUUquy74ZcVrl3gwI/01UdZDsQpP9lO7HlOf3ZbBO1bQyzgylOnPF/B7C9xWb
IsK/vAiecfkkH8yMpjnK/9osn5N7lR2a0H+Bau4B5e6b1cvXVEC8oL4gCtsEk65XXzRcOiu/UeQw
1DRgIX+P33356jhBeCcjLu7ZPgSlhCI46NDW9ytZXcjw9K44nimsFSCQppTakxS4rGzzsSDuzCAf
6P2XipdNLFPDanIIKlWKEsXtzjRt9Gzleq5I0oj6LuYvk+SwOJbJsIhXNNbV/UrWXEld/EgevWkI
pZrc4fifYFGQO4mQalFAF27aWKrO634v2S9Tn8AeM3p8f6yip/TiwYS59Xr2H+4xjDwknMekLBFr
dV62BqDHaSP1NBdMxZS9RQM9nvktwTjXTiiKtvAJPPeXLW9Z172bWkQJaTCwanZ5v7UMaFdnPozV
jx7i6KFLt09iTxo9iuLuvVO0h2u270QEYJXwC40FlqSZwSNgOn6jPsdYpgLsAzL6cggDzPbwbBLU
Nq+PqyrCcL9BA0CmuVoogAtN0FThA8UmBEhVZdgACIlnwxq5NlVPEyoF4VPlS5MANHTY87U+SFLY
gq4nF4JHXM/gxetGy7uuNegELQHw5KK5lZuleYwTvnxyR3Mudp7v4XEGiUCKRSUx9X/qhs71KsTB
5SdQlYVU4FHt3Y4Iy+mFmbGO+b4/3HuQ78uNmz7iUJiGZpN4sus4EOXZxxuuLUAfTqbWyq0DdyJy
e2FL3lQs+5o+sU6Df6gBOxXBhVDLH/77TnX+8vFH9nltBSw91794Zg51ODFntrCmbTzpZNhEqOnm
EUX6UFvDlb/kqdd1oz+fDnM/71owNMiIetbd+XFS0N8CZ50kZPtT+cHBEiCg1S+i/ZPWlYqzrwvF
oQLV0aQqaCLIo6YOulTkKwOOS33em8hxc3UkKtT+bU/cejZNhPQJY7G+wC73nIU8nkADAxEA6uF1
qirCp1V0JYl7pjvbFO3FuJZ981Y/yRRaU9teNvap2awutifh3/fxe8roM0rxBBBFQKZXV8zWk409
sPi3eWpYtlABAl+dInY9stJGvWOsuHKYnJGPiXJlUWlmdBpSeeGRuU9I/sldnvqlA5fbV4a6Of8Y
eIPUCNFx7QobvQU2IVVNKwMHZMRzPf6SXEeCgJxcELhlJ+gQh3XMnDNqVLzQfLfRIYAKylC5Rk/H
rJdQRQorOmL0C3Hw0ynFwc58xfmyn/l4Wi7sKVZVw4SDemCzZZbc+5R4JgONVuKsqJ2pZJ6JfMBf
YvaiRPuUVRPSQpyRN2ZPuRyi6UA7OjnP8cM9srNQYR/Qi5nbUOV1jmtqy0fESyfpAHH44zZGOfdh
zEzY1oGfkOsfPMA2/781NybJZ8/6hSbY5TK3jdvJV4PEJbnZgP71u0xBGiOz4hwQ/3oJnBTQefY+
K7wmtFIP1pE3QHf2kMDIpFr7goPROctCe9GD3lhYcGVu6Z62R0yqP0pGlfbks3pMSSXLsEtiQner
u7M9TxpFE8S4R8HQcH4isXvkCOrC3CFpo+AqwXCtldUo8mlO2Qbb0MFcuaTCN8n1f9qQgQ7bE+Oi
MwEA0X+8I/WnIG3QVDgwwBZOTeIQB4BwQBP/+Jp4kaxbJgB2EeuOpq32wDBFzKQjFh5S+qA6/4lQ
bt1yt+noRVChjTK/znzbopBJfyvNVWrUTmJEqN0W2ryViBBL1iUMRVX2EpWSa2jN2ZAXn8jzFosZ
zzFGZV9+wkR2eOoHKy7yAKH0n3i0FFDyBManABwbjO4Xoytrq3Mhw2EeH8atra4apngrkx0Lhcex
5UyFkyBkn2JV+/ygZW0jVrHLk1SazvG/j18CqogFarpS/U5z5e1J1it9TCAwj8jbjAQAIF7NgfNk
z7da1hnYjM0VbbaRjUYZAXTTbOCWfTpCom9AvjYY7a2OqpGyDzWlwzgi8fNLs9tMj9XVRsB4G8jf
xqFNhTrQSk2YWIFqAj2uY2t+NEc7I02hLpbpIB8fV50sKqOePX3bgilxlaN/wb33hCZ+X+G8WuN8
pIWo0VtCtdvOTRTzO1JmWsRJMf4GNutpkTc8ESNphr0IGVUf+yuEyAQV42aMrCQtXJksAz05r7vE
qrpKzL/K//PNi+RSpck3e2SvXRiv/7CKSvk/WuVxaj6KBVMeW7Bk8X8IY561jOzITIFc70n8bqK6
i2Pu7q2+Qn09vnIR2JdkG4MqhEBZyDFqwu5be16pQ62YxoA93Mg/98HWdY8LjXNOR2TkWKHvbYHR
zp7jTSHHk6SoLjunnMpDOFZ+7isdtn2gniPuiB+/WYPqkIuCUdtmaKWmZArCEr7I+KxogsEAxeEz
eNfN0hgwIw38VEe/TX2IBQ9PTVef0jf/AoionfbCY9ArivcN4z0fazT9ljy343Ss5Wu4/8kMRSFF
69XVgk7KnuV7Q7asd9/0+sK7FtRvCW/P+GL7gLFVCoHVrLnpCZXDlmCk/e1ci5H1Db+CHBbZ6KgF
QUz669A29vZpmXJL0cRerWupmm2kgJYdozBgjGKrjz8oWABaNl4/XD1df4BccgHp5dJtGUb7jgub
S+Rtfofuc5aFinBRxYvDAeLiAqw35fkY/NW4VPoKf8h0VbcbDgQdoBW58nTntdPsiDJvfYCDnryp
DR9TdgXOtpZOzyJA65z+VHFMlbWPgRDwHJqGgvH/k9pEytixVbxsJAV4mL8bQ9l1nXB2SUfZdj8O
sbTsdvOFjlbdxBgM5hBnRSuiJfBNyIYutQyKMr3sYcdVL7Xu8ZaN9LBUaYwTuw8UDUbjzlzMbDqi
czguB6K+ZKQAuANZEnggo4oOYFcRFjJPxSTXMKpdslbeB0JVBt7uBEVOVRfL2mnkDMd4mNX/BMBu
hi6vzAoUEhqXut6e/TyrbaSiZr5S7wKTRX8wjjLEjVIEbX1FaI8BDZG3bUYJcCyumn3sZwMnX6pG
J4ncGknZkEFGfZem4EpB/tVFMzUJHxUVixj01tPevDZlcYTsJDXe8M6fbiXmGLjtWScknxLqW4Px
1L2wRCCeKL+KtBIRBCuiTPrwrj4goZHFux/70nWtWUK1JtsV8remJoPBfZoTGVft4ABOuM2wh6k8
6YobOtEW4IGvBZZYNAmV1d6yg/jqt6RvGK2ll/5K+wg78sRTSGmgCir0huTbIuRYHHHe2fhiHn3u
lMb9/QpwyGd1lvkxG50v2PEmUxq8ROEd1HOFlDP5BcG9UKKc/nXVzW4X7QYhufyG1QkDnedqbGWy
fXX8U/tzMFTNn859/QuYGviOtgZiezT54MdIjYej17xdDOyLqfRGy8tvyf79k9Pkp1gx/WtrdCKm
8F9pdGTqK3Fdqrpqd/cGIO8yJibRTVq7f3Vtnza64MS9Vj71O0o2WvxK9/YilH+CHl+clOIssRO6
upyjuykxWjFBX+cA1KGziRGtJ1/pSiD9+LOriYTPZCGl9Iah0D4M9Io+2HX2Kw0/brL9k0UaO+RB
HoxGIZXWr7tJD5203Fb3SzIRYzyLNcinVKqT0S6H7iLsyC6InU9q24wW1+ZLbBWNDZrAqABt0DDb
KsxjZMDoHdTkNWpUlqVt1tFZK8I0a9uxMWs8e3uGcqZkBUxix4S8OUKisnqdAy4Al2RCLiF/clZC
9ZQ2FtPXb196DhaSsZ4lduJF9u4fD3kGQTUuP2EgHfl1w/eJsKzEmKRdNKtzATqN7FvuSO/n8GjX
QkZ3Apq5sEHWptQaS3bSEebOXPZ2cK6abeXju7j/UEAKSTbz2W5JOX/VWMPdrSbINY0S1vnW76gm
cSftMMSUKJOehVb3tJ626u11NV494yDanMpM5BHtJBXmWzdoRHah0WiWm+rFcIv1o7kfcJO0CkV5
cQtEGPGq8ORvbGJF0LWzb7RxuXMgx+ladcA+toFZ81wGSmgxoyPGY52DbBlY8uW5ttZ2heN7rK3R
HQwjP6rqAReA1vlhxUpwtGeN0aTAx8cGS3HFYvJorlVcZywetbIBwmhefo9rT92jFPxZ5lZYU2gK
lUUCXS6aUs2VFbppDjiN0M2tub5V6ND+BRNmZxl8xHmYywBE9npMVkPnx5JyL6UXZch71gs1ENtb
X/DfyGWDi3cxFD3hae1DS/Xx6GW/PEB4l3iGNl1QkCU5XfBOBu1vjEYhz4a+Gj33eJxnlthulgju
YAWAwJy0bslCIVJtOsCILMhsquPkMPfMfArGOCopusw2boooHSesXa5GO1W1ZR8NREHl9NoEvqDj
oWge6vFdkhmHy1W8O7ChCOGCbQm6qp9AP+t9B4J63lv/1oBWLXkCIq/D3Qb3oYvlg1OsdZjqTFTl
WkLwBxKKAUPR7vELkpBLVgcz6RPbRfP7Gx95SCywLywlwdCY0x8FKwf3YzyAnur4V3oeJssm/oz1
C3UDfwJMlG9T5sLte2oJTXCl6Vjjq28mMsbKfwJo3tcWF3gDTcCNueUBowkNSDdu1LC6QBcO+Xre
xwsKGAWY/fdgMfmCTOvbM7Y+i3VY9UErCLBcOLLAsY3dCUc5SKnx/9iFWpDPocHUgxGehnotfoHW
d5qrROmNiLoIYRyE+6cHtnzrmGKgkv5jDbT1KXsHxMFXkJd/R5UlspbM95sJDfKnUgth+uq62Bwm
XDYcuFakC3Je/xrBL3x56Uqd2g45LIbcDDfbjzzjRcsThKi7iadAy52fqPFZBo1APg18FImHLE5Z
hT4E5rdn/E6g0VlOwIOjHn3A1oaGEHoNNEl7r4M3wPxwFGB7FeeZCDEW6MgGo5iNNqthQfqVCz7N
cCW/nOnSYW1say5K0iGSA1XygVB2F1OwV4AQ7MXlz4VPlQblypUYQnGPyrKvKNBw9FQLiaxulDPO
6l64LtJoiebha448DiUSIiSyAI+F9XROl/rdouvjkwMoMjZufRrEQgLmUe+7ID/bt/lkq9mWtXIB
SlKc+mb2ug//Rdc077y9DZardykjvWXcY7i3eYJFlu0TuHnAJKuwQx/R5H1/Ivqd18mt9FNZbwNC
6QQr5YvInw==
`protect end_protected

