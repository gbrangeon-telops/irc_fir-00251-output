

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DYkUg37UnVRJ+X5v5iFDmCWObMw/mUCrJuxa/Cr9wGl4FgcJi6OQesLI1M+aH7+emQJssoNWrh+N
iL9trwbpEg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Vb74X6mc2H0e6MLiEAhBKZ84QSTgHhg3aAfwLeb5H8AGScZ7UqNDKDmI5IhuJ/LPpdHQCtOent5+
I1p5tELHTH0LzN6BILTKGZBdaGJ2AKKoofyljqaR51srCF/ZJLUOrn1XUZMkdlutYXGikghh+zK5
6+/HFEYyz6zhpfFGpAE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DUY8u9eRLqeXCDG4E2/8OtDIacK06AysbSio1XfMMKnofNQFNkb8eAjngrn4u/YZ6G16ZNMG7YoY
jk2Rx2Q3M5GrNkHLNcW1r1FM93KBIPYna3s3UsOdPXI8u/gdrTwtTwv/xpFT5pO5KUummozg1ol2
CfVK4phP0ptL6RF00qSF6IA3NotRdVSf39i8Abyti2fNqAeVQtQbe8y1/1WV9RrHHqEjarv5sqIY
6GslwJ8wdJjPL0QS11gBEh6rDpndqUhWIIFTUrFMd1tEU2WzUCNSxtbBPYlWfpU8e4/l9e5xSsF6
weW3wzZvwjgR473vdWcupdpbpXFjQjfOA39+/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
p0GGQgjzPW+6PIUsMdZXTQnjW6BUopNyvt7ApHmGMwjrt0lKkYFdeq6NnHPNeKi9xrrloGAO2Tha
FhPoK1WSUQvFoRR4uKVUk0OywXYhciTgYL90XL5T7z6pvP+T2xdoDnAiUPoqzH/Ubhhi84EoGyo2
+zIDCCcTvvnznOBjfpk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m1/kaqW4ETEcDTOeEJMS5yQHRelnhe+7sXgpcKiP6lTf8NZHj87LtgfMx1Oh7TGMtL3OsgLwXKl5
B/MVSSTPV7z0P/OvFd/MWYJqIMAVI0yV4hJ8dwWC7KK/kawdL1h0Q4iS0dxjn9/392LJCmqkJJmj
TEThXH1uoH4tMKV7xRRg0/MNNOk8hPErcV0Sx7ZxMFsvJk/PuOEi0wzy6daa+A+gop4M475HPjAb
iPZ63o2focv37v9R+NETZc+LyDzZAZPFDxIiHCnZlRMpU+rYc4lLu+Wj7afASerzvuIcVvlJO0R8
MuDtSunchT2Nxfc8io8WUTVsWpkmP/zQb3BvSQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18992)
`protect data_block
XOuycijkPjxcOI6dX3Vjh55f7z+uMKYhQEOo17cA/rGLqWI62eIsCc+KNPoxNqRfjwO62dj9xv4A
xgKwF/KVURDJXuXLfxUFJvh774NTS1xb+brCSXcv9+ZsYdRba1lhSXz737Gs3RbhZUsIOQ6ebYPa
oHWYmCrm3VdoKDk0dG5PRCygSqzQiT5Xu1b2Z3C9umrz3pq97T9JRjTbJ5Eas5K2xLfVH2w4rlE6
/TZ/La2EMXQg8Lu6+OwBLuQiRKNbpQvAm00VILOsxJm/yr/JHLWR9dKd7PD802+Nhl3KVg3X3jPZ
z7P3ymcuuvxTWiaoPTuj3lVOdAK2UU98/QvVxvlRvoOtBxW/oiZUAHrMiUSPs6a9T9raFd0/oN1T
mvxfal8CJkfrxrSvhSjfC2Av6b4CFnwQ1+EcAkBsCA1rlTNUW1OMBDq+YX1IlCiUaJGCN12yX2nc
9vNLA5T1BJ4497a4iiE7HO7YkAVcUMSbv0N5bzu0ECxdB/RWKoy/11N3nlFjZPrkXpBUMRtgESzz
siv8vkwly1gNgZoZV9CV5fZRasX/xsLqBmXDBepjl0SY53n5r+i+DCUuOS4Bv97dIxWX0qETEd+q
GnNSCgzkgu8nHtEmwhYNphAV4O6CHHggIuBry2l4tHQk/Sw94+CFdTnYO0LHaoSFMRs5G+j7m/bJ
jav793M9XVIT71Iqyo3tPCf/G3xi+en6/NWdOYTENdIucPUcOU4GqjbJNGE88OcHH8oFme96xHZk
J1O6zQFT4H1VrEaj+eeQnhyXX07jLtWPoVDZeKhsUBanE0WulOkGdDumIanVzjJ32denyWshU2mU
3V93RRcsJQgFiXvfRGtMml6REf7+7xJqqN8fYQftxB4bDlkECCPLxDPCg2hxc1RRBGHjcry7/xHM
WILrJQ0ApYZU/8MeRsrXNherA9eytVTWd4FT1zGsQUFNLnnEFxeaMpv/yZiZ2CXOxiNVjpV3rgc/
bqV3i7Kwxai1ocVfE8hR1esYUKKcHh2RuZE8kJwCDvM5NpbgaDUuZ5YAQ+dEeIA3ZVcvNtsNIQjL
IuC/llIII3qs7KZoLnNFXbYxvcTEbLe2g/4cO5101t1hXPuCCRWty7QDn5jJZU2asrUK4ukAfq2F
/CLK+7mpEirCuu8+YxMdarFfZDvQU9UVWhNDvG/vyjrsCp5xHVr+ORH/2thG1J0B4tRdwFhYAROg
tEPT7L6uroEiKSYfoXlze6iifenhS0t0mEXY3gjL3KV14fzHOpnWQDxrC57wYtHR1HC46S3UqX7C
QL8TCyRt1KWqp4X0qsG7SHlejcG0Uem7VCtFR/Ggc9+YrMIC3wkkf/OciwO/UnqsYTDOfMj7vFpl
05e8iDavL0N9+UalU46lRwP5dxynxZakKwKe11G951ubrdd7qdKFIaJhfZDlR2FHOCEK1FsIjaBm
NLJxgwljWwUmSIYcpUoyZ/cwzTM/0vIkgqVMmBzByDdlJITpvldRMRJ+B103PEh8Az6rI9XRawpt
xHdh+YH/0CSD5M08eeomt6uKBloV3G9178BNfFgJQHs3VwpzGhhaBU/WAcnoGKTDsojfVxARFqC5
ZG49uX+A9XAIotADFCUXTNaWhKIl3UihzkdaCZg8Mzt9ZmfipNdyT3fFyOWMgmmxG+PrVvYPLBfm
0gByetIDpFFZ+GAW3uQ+spT3AHsIbdleBQhdZO7GGHn8jKpI7SLoWsVe6kN4fyQ6Qblp4daMaV5E
JvFIrMu0QPfywTvY2gEgxwW//mwyQLhnUpbVoxucVYKgEV48swvo8T1tNWjjczsAN3k7q+qKlJhi
swGQ1jqUsN0S0GcZsbtVznk9plQpKzKoJFsrqo8f4mQ6viwC0cQGm+5ZuG6fvsmTI6wfZl/MV4a6
gYbVnXfipTzzxnbixCOeDW+lmKf8NTZOXtIK73fhuUR8s2TMHRFYodumHYU7fF3aIRyM5333mQK+
CFzxPVfD6KqnsIYpO6K8vWuugscVhNFfPSpHlzqyyw4hRyCntpmeHzu6p4TM3CbjLmch0wNuwb12
a++3YlSpwcbpwY6IcVw2k1eRF2nMTko0DnvXJDcbn1edgng7rnwxsRF6z3uSSGY2TQRNoQJTK9/l
4gu5wckvslLrA/1QGWtY+46TDcAfkp52N2KNJ5h2reNN/MvxH3+ChEJt9vFSlioa0Fk6WwTCNOVL
5AhgAT+lQM6rfqlBNOJtE5g3WKUV5/LELGfpTmGwmBpVVxGyIDKZLDqK4/KHfx8e+jY3t3/5Z+kp
ZQEixLTwOiTvCGyy3tJxK1fWmD60OZnArAg/7CzFSruyNHe2/zl1wqvH1qqsQXuJcKSb/VT+1Piu
DPJMvxa97hB0+ktGgxmYVkoVLsgg9y5MwrOiXOGkawGt1zXW2ka3CbrkNjc0ukCygtC8Ca9dcic4
tHFb4YGtNL/FJ8UgwrQql6Jn4cpidilLBB5D15JRQhnFf4NyxaE0AulR+U2hSxl/+tRLUzCBmkFu
bRf53reMdr/zwr8aWyUMWREhDGFNFtmtUrxx7dsfnOLMJXy8twESgb+EqiqxtIMGVg0NG3jloTlV
5sfsOybUqVxu9JhOWCJpcLUQLysOgBs4d6OCQslRW+C2SZj25va+BjHqMDtmshbpLMWgFSLTLM/g
LOoDZjkQ1smn9nmX48dudsNGIQM4vp32GJjOCE28KQ5COWaa7mlq5ydByqyQhftIej8tYufZOylw
Ht6hjjeKlAVQ3/ETTToOyZOxQKpZ4KD0Oe4tyFO49Sztl7lO0dRqgxfFDAAhHiNxZQbx246mkc3I
17rVXzX2LMhP8AgysWyx4KNkoxyb1W9WyhUqXcHMhKKNO9jg2KsP1FELJHHMvdvTs6J8p687KJES
Bv3fbsu0EbmcXHsJmNGATGH4s/knA1817yTCxYCP1VB4pStuPcxBUhjNjhHfscJPOzeMcMpv7K4K
VSdl0XrFWjywdovgxtBk3983qfPAfuP6W1Qvy69bisuWpc+lynbqMbYG0wzBxcq5PJ6c1dUECkL0
jTwbIM5wt3ixHZiHSLeioosEP41CbBlueg9A0DtNG6r8jgv0Azx20JIpX/SnUioxgWgeSfr4b+s6
gof6kUvjtqsTG7vftbI9TQsaq7ZTYUYPCfPLqPeLE3JKS+cMgW8Uo9PsSO3Jz2hX8jvTA44kKunJ
M8a4THMUkGjwWzjT4c2UBZ2JgdjHNymZUAxPn5Vh9F/7AMn614pWixd8DVbDwd6LzGWO86BBGGWs
4xogUOofIMsu33flE0yHfOslgvDjPrNkdjWgZPBhLv5U5L4NjsdkvaE7jdV6NiU2pKcmAJQMmFbb
C5lvlCdgyPxh0iWtmDwpD/wqk4kkgEJIzD4eKUd6tVVjOioyFzKUpeg921F7wAUjOD4QZOqUeT+9
Steb9cZKYmaICQSC+gWELqxuK0t3LKFgj2ywpw/rwVudmC7I6BFtd5PLAODY3E7St9+cBh/34ljC
7baGbB6WdhuaxUyCsiQcH4I4q93oRlswdOP5z20Pd9axQKdEAgtgDODE1PtlUbQGqjPB6qRIdpo+
/p1RfM4Zmczk1xXlgDOTFgqjWB1uGKeRxGw9o52OpRpVms2CUDqPVj6fMBzcESkwXDJxNw0sNp7p
9JRDy55YFkXkPvnKt6fFGScQPKcD6xTjxHc6LXzMk8AewITYV437QUfjmXLXwuy+KZoM4KAjAnNA
7gB6iPlnSz7R1MMPvah3OWJUNOEpyIy4RXI1Y4i4YrRy0Rq8ugFDpsHuk4h1m1w1GitI1exuoWh2
WLuEO6lsjk7/36jPpLUGy4rAUDS2QDVLe7FHJNKcWvVAAGJrtjv0GINvCDOLtKgqYBAl5n/ZahW+
os9R9oxMHFW99oEs07ZPiEatW+4Pdzgz5r5aD2L3ym2et+Iru4feBU6ENr8niVQ2oAgASUrFLHxd
SQqBwh057h5fpBHDhbBxYdDf6Xmg+egp1wA8nYwBRscgmSb5ClzC8ZcKmucYcDKU0hNQLw8J44rH
5yEKnRX6rxD2O6ugY/QQbI7XOjlZnqXdYLfysvu7/SH2/RmSdL3A7KJXSZD6DhZMag7/o5RT1A4i
gDwYrrjbG+sFwQgIyeuaSdhiOv/KmYkIC+ugJ9BlTYqYLtxYfoOXb3d0ZpALKxDpoLOCKICWF1CZ
7Hojg0J19iP+LFvH78wy8es95OJePFsbElpAwiHgNVi45pnzCNmQZdTs+RX9oT9RQBdQgqVqDxEA
yenH0RT2gHtaKdArgqFIpfZpqLtqWN+v5O6epcVJm959Nhga1cEEQhbCqFrxjufEKDo5s5m9Eig9
axvCqaXgscpX8Dwgst43aJfNaPNSKWI9ZNcYQjwfAz7NnjWgZT9B6rCNDbx6KumALILIAeozYBD6
vaUVjZOf5gdNHozwli/HAz1jO93cNbKRQx0GUSVxYG5T3DhJ3/6/Hj/bVCFpuSiLr7FhU2JMOrQ+
zfMLlPNAl49el/fbwmLM74sl5/PYDdXsMXNXC5oS10crSWA3r/M0u29eqlafF2OTw7+ccdu2+Y3C
1PNIX0BOj9ojadr/1Rxc5pKlJah1tBXoKoJCv6TrD6Zj+jiVG/0eh6wqvX8KvK1hT04fncD56sxm
yzB9JsNyphilBfSszxsbe7SdxgO6O5IO2t2fzjWgmN1QDJ3HhK5d9vZrQ3w+qom2Kzrg2QSl4yM5
W1sthNaQO0CMvmF89P5OGV51Z1biExv1kcetD9YRd6bCVVusn8aROp3lY+cg5+BBEpE1qYG+ihLe
P2GoAh7s46NcC8E+FqX2TrfJP5P1c3LB1cD5sknKxtahutGKSoWdNcQI58k2sX8fU9Y1uDKC8cBs
InKsQ8MBAT3eJp9ZZ2+L/cRwvsWPmOUb49/Xn3M+bXjrzzf8BDgAZXI9r1oml4tN63K7E2GleKbL
OK6zR/Rq/7eB3vuCMJGcjwK+AB5yYu/oqgTo8f9q5NyC2N2wndOUAd3cIcc8ljuAiuqbJ0rm0z3p
HnwgVt46psFTGULoixZJtTGExtMKLLALmAubrukzNLo2L5jHaHLgggKY09PfETlzaPlYyBct3V07
RfVhcj6a2pS/Bd7g/ualqqOjb/UXSAJNotBrnkJd48BVVmU3T/ocPg8eeNDxT7OaaJIUH8/8DCqJ
PgTtKu840ZY5YMfHPW0UIhek4NtRXOs5WQiVswWpS/dA3giNyIpguvSC8AOAlIrxTtKcgsi12/9u
J+YXA6hvpVZtMcS+S26OImzpsxOjMZN8uhJGVG6vfRg8LwlYNBwQpk9JXEkqwedv4wOYaDUOx/ji
zkBuJdfMdW34+OU9PIdBOg+BgYqQlgStjmDX6wBumobTtQQ+05X3CWvtZJJgowBQOgvH/AJ+nMI/
PNOTYCdh3Q2sg3K32G7WYXVsriAwSAs1/ySR3mCenz2BqUiUzeytSylwxLZYHApkbilCIUWcbCFw
vhKi4/anWY92W2AHGo42MZUmSVVysAb24tKyFIqWaQYZwpfBW2uG8JVyMFuJ7g0ipLltPamS8txF
yswkoZSE32QBi8zi62+jSDdWSAI8ehkorKCRoI8SRr1te5kyIk5oiSPxDvWFZ66yamHFhWTI50I8
2CVkjYHd/9Xzr+hbr9y92sgxeCN9PtNV3dS/vVeDvZDh5PAQ68J2JgS+0LBRWP3PebjCWWcwJNoo
hDAET0zP7ljIq8OrerlFz6nWOsAkQC07ggj22o8xvN06UA1s1knR8rJKhm36CkU8cCl1KDLezpby
/fJ1gcB8glLylnEizRJEYFKVFoboOFh+DG4Iajld1xQuDYiK9t8n47GPNCHYqXOXjvRJNjmcKcLB
C1VkaaNlnADugqCY/qikQUAL26TI58Ql56iVhxpq6wVxmgmpBJ4vsw/8kAEmK49qWTgMI7wlcmsc
WXSMUWWUxpiQvc2geN0kRvWUozmvErlvST90SEWkY7hf1wpM+p0AgKwbBqHXV0qXNMOVK/k+0Uot
/wMbj16LLvqEgqexeaxlNPqWVQ9BSx43SJtJs1K33lmEHzxgwWpjU4zuJRJbQhOn3vyGzZLHZzbq
8D35odeh9GaKiwKXmXcih4ibqTcdJQCgHLLfI289qhSjl/G9uBcVxLEu6wvVUyegf7lZwGqK6K03
5hY8R7M7mk1EYW/TLBtn2YCdfpbug9sK23kOqNAGotcHg0FRySKoyIWJTRcgXGlZHeZwESYIW8ZA
TYKuK4L+Z9q4kK2ZNtYdIZYPeonfGgk4Xq55nwBlfCNffiCxE5amJPuFQvHxfKLeeK3YCd9IthNT
vb4KVSpU6LVhDN3b7nb7YM3ECXyNbm/N8uAWz8X7Mw0qcs5YFFpSlTpb5t4BITYhpWnf+9BtQ5EA
i6au4Wpw2QyHwfqzuWrO9B0K7vpHQlmd37mTdAyyh7QhzraWPoG06sj7zFFWto8SHQXVaqnSi4D4
uklWO0V36ilmC+AkASNIavg3qOzHvH1P058SigpluzPSjeRKEcoV6jVZkM+d8JTnZ7mwmgDyrJ9+
4YOA15DQ7rBbr2fIXYXu08tX2ZVKTY7kUuIIj4RnPWYGG3GooHKHetIh+N/BDJE+T75ANFprsBU8
j81lQ3GUX27ZR7Fzh5N5vodS7EELlqMjQdGeixB1x4zahxDtROUuHVcmhSpf6+eaDij/oqyB/iwS
r3hfJtvGRHKLgLNRbhVHTPfqwIed1i4Mq9KN6r9iRR0X3sRQVRk7WFyTJuXvIlohxOfgg/35dRti
GZ6pFQjYZR0OvI0w/wT3+MM1gf1mYteflmNjtRlR6VBjg8xAGtswckpbB1OAIMrEZ3fwXJ3+lniJ
1FLT69jB6QriL6NG/vvcLmZUZs2ieh4rTWkqT4Te7jnEZPVaYqTHvOSSGQq7sSdGgLIUKcUKLG2s
kVMs52l1b6EYiFgLfNdWcHvTl+k2y0ZpOogNRpxGB5+dSGu+z27n5lM2YTNpQH5Rlmy4cGyKjfac
ICIa3eI+PnIx+2FZAc2b+OgSD+5EaHCeejDvVdAr5YiEVxBE+ZPAaAjq0L+ExL6dAqqgy/YsnPZR
QIL+9BttyZRIl03iyJbYKXuKkbqQunTnOMmDmGpBuIQwde9yEb1eLRZdIT/MqWT4waiaZR4jcQZX
OgVN9qqDAwSBWML38P8Yzxrf4Uh5NWk/xRE2Yk6eZBZmN29mBuFFjcwDC8qCfhnoks2V7v63l/ST
AsUdjaehbnwf6edr5ti/Ly1Z2JXocpS8CfNb9i1Vh2O0nUvu6bafGwU29AUV0wsWLYGcu7l2OtHZ
lK/OUDPZfQNgAfCxyt79zTcwYoPduPB21CyxUDtQWcchmulrMYqemplUZoFWK85gHG7e6l4OcJOZ
svlEXGWx7LAyzrV9Spt5g0zyf4W3rPkx2VRMdH3ysGDlIKN5kadjP3yzikUBsvF80GWrv5AcDdm0
5Pe7EtT+k+4S6FAcqVPAMtmyCZRIaujF/HJa12Ya+sYXeL/Sh9BlsmK1cNGl3hYRblafjlraZnRT
XTAd7Jw6EXP2TFyDPDfr+nob+RDRS8jtq1sBv0DaUg2Z3w22prc+sJoTt5rwpLXnaDUbp2uOVkO7
ksgt7l5SAidykVx7Z/6NXRVZSDIA5OcZ2YUsHjH+GD72gX6/AH49GIJu7OALUBsEjkW857rk40e3
7y+mCxEP3UF1EDriValhC5z4DdrbwovFw4TWznA96xApnYZqvqNaVQ0X9tcdT68/4167o+YLxydt
qPwJGIrS4CH41KhF4z99cU2dX7ZSAywW/dNN/KVsYdJPdquJ0cDM5GAyOF9IMJ/LA+YOw5M5lytR
rW5uVIl5m4828JIhFtsBYANshltfT80SMIpNH94wWOXmG3Nsx65LTAaWJU0ezpdzy444u8Sx/FmQ
OM9RFMx+GtiogX+hv24JPo6pWaZQFYW3aynipV0sh8eIj/5hqVc/I7BToVWld4h8jhnSXy0RmTVd
fshnaf5HBQSkny6Frp5iI2fRy+G+IXB05VPVfqSIXxGlmdbFJamdSXp0rvTIphtSvV4Iw5vb6OwN
q0H+PsPLdKrRH1lrjSyVdQFRL30wXLGUoT2LT7Z6g10AXcfjRdlJOIKmxfqDNzy2bWFwt6fa7/Es
IPnCtgw6KndLDxTw98FRDxdSMfJfi2ZUma+flSkEfj4EZzvZ52BD7rO1SapqPrioT0yt3RlMmEAK
Db2Q14UUuPzXA6JwPAl0dlq2iuD2z29hTXi6DfcxNO4DmM+roTCpJY1gY/xZVYMpxUaWd7ShzO3y
z6Ct6mzbT89Tzi2MT66GejCdBhI+iP8h1DCERqJTkvoChnpTOnaS0TKBicovhYe7VaiFYXIjEWkS
LNYbW1AqRRgN/0I/E8umz42s2o1M09UVirJtCGstiSLh/MFi1wR6QjrktRtwKDkCavZDOz53UTPr
sgUcJIqXxSH7bzEzscnlQT7Vgei2Oyfgxp922PDRvy212VsPgu+qtWirQsU5usVbPenHceJ98waF
PojBSbn9952aaUJFpPvQxVrXox+lHGCcUPS6Ue6LhikRNJL5Dox8gIpYlxzabVxCVx+mm20cwP5i
o//kp6OO2n2zCO2memnaBYk7jAR8y5bj3yuNfkqtGVhhh8Izhg3whl5Nv3FFNyhTjvxnltOuTB5v
6oclZ8oP56usGunKdq1GDryVtc/GG37dvR23tFHjT4DYS6oA+tUmg30InThki6WCnWeigewEXxJX
aK/JTn1vLD5XFdyAPDkmFw8+O6wwHFGkhaujnc7g3LYU4YOLnnlMRQvJNIX2MvJqNoU576mXgA4q
YnTpZ5X1VNP7wyns5ei5sULk23LdG5zF7HjByf0NSo83NLlMtQhRjjSZwlLcmKzRJGmFBgZUmWJD
kAeRaiEvPEdzCnbgaTfCUvYhe9CZk954RowO6FyKoxX9iKRDBTXmSQ6xB0nKMk/m98i2qwEo0CLE
OzgY3wpLaZmYBt8tc/h6JD/hCmyLZIhR7H4NRdODJuy/yNPYSfbBGPB4mnzN6CvQsaDHBAs4MI1C
IcoXJXSehN0jQfyjyoq3fFfV7gbkhAuF2wrp1VdUJN9WX6CMy5m6mIFGEtW5ty1r/+m8VYfIHcrh
lC7hVU7j3ZPCNiNZhKj8lx1F9pqgo622SdlrAgmKxm0FGu+vRXoTBw+U09LhfmOM8krxvNTUCn5+
akNHJBJugG8QI8U5HrD4nJJ0Ct78mOMLY6AHXp6CdozmaTlBqIJrMRVcEVukXb6LvWsE1wTysxol
6Vl/7n2mQ1zonO7FC8Hsv2AdPvMn5XHEEyMZs1ccTpTXFyoaELnlv7u+QaNluccLOR2T2ixkdxAX
o0ORmAXr76BilQky/mR2M4Gz8inzFNVsX0pQ9ifxMmkbpA+GijgueC9HhCa1PJd0pehJbPDgNNBx
pPnlYEz+PDEScLr0leuTBIjo8IVuNO+qULbe0CKz6M/9xiwFZK9l+eiYC32RRxCm7booxsNFNKe+
1sXkzSi0z7owTfQ2Q2xSJRMyXbPUFfoRmz03E0X1u3edqSTbsPJQArgEt15MoyPaZBpW/NHzN3h8
h+zpr+A2oC6xT9tehkYw1qx4/f+SRPUDUtlE6V8EYe4iQHVlP5ZgYPlHx262fnmzA6FHWubILhPs
bQeBmc68hSkRE8b8CuUg5zmbxb+p7YOffA/9i1vkNhQXH3Nf5oNIfDyWO/t4vM8LGs9uyYq13wVe
tHFM9mdAcVr3Kqqgz4coOtxxJO+Sz2TE5lh4CYIz8Y/dPjZ78FGHH8I+gRvaExcRkvqRrdmldv+o
3ENJNdE817H3g4Y1rqT58ayLFGptGpG+vCsa+EoY7sTUkXpHeOgixiP/sA9M2GzbSSzTyqjYxCO/
H0NqRRw4GS9XKyHuxFxUYuckGipiTon0zDpKBjJAS1sNa3pCtUSf0jtda8nFl08lUKnYarZKt8wT
rDNjZXbhDBnERs0mlG6A2C79ZsvePyUYCntCDVDW/vXY0V2ST4P2i2Kg97DVtdwM4rdqPmNHRcGk
nJUCKtekkt04O1sOoWiYkvbZFNQXuSswABKuk20Qkd2tnhHWOdZ2w834D99WGrwO7Fnij/zWjWvd
HAOWiNgpB44JzJ1fuR8PYKEluobIcoATZXSMH2fFsbOyrKM+nRSA55KH9OhGNvQuUiAzMwctdkO/
k+4fcdnao/5VSgiCxVGMgxTa/ZLeFmPDr2b0hZKpH54XmOuAqnDnYvIkGUbSD8XMTnG3+y3XehD9
1IOV80/C74FgXAk+pg8lG8VoRZ2NJ7QeRIz68WUnkXzDFd40UjiwM3tdQ/zbyjmsoi2NSuYMtM8D
21nkuORZ4LYJECgE8/b8HIaS9ExAdl1hSQuz1NQ8FgKRKSOvbKSgnxTuxm+WVGYPLdQX0pyxh1Xb
Gnk8PBDppnPIzjAdObX9gO32YVnMozeec9G9QT8S6m1WpPWHEtoy56Wv/5MWHKqG/OiKP1xjzJmK
tQcwP4KXGRm727BqYnlBGGeVPNhdmYqADsogVenBEnSc17XmwuzaOj1OdgSjosyZp4YCd5U9phGS
81vy042B5uA5/EebYl4ilns40DHm3Crql2HzViKor+gwS1MnwPbMfrNZojJT8BkIQiO+Ss4a7hZi
QiIZqnHxfU2Ytx/IS3iWaoPHK+DEZJJB4K/tlEnWeiXzx25tUKv0Jo/2jPPIC3smYV5HfUIVtsiO
C8hZGZjBfNswdC6SCdSLDTl6ovvVJFEiuybCpTqb0mZLqh6Sib0Cg047QAS2ypcybWLfrbbdi2sB
djmGYK3y1TjsOU6eU+oEbcaXtqisQTJvsk7ZhL9IiICjKgocv/uikN0rBV2Pz/uFpB0+bOsSGCmi
bzv4Iyh3Kre0RQ1AvBjtqXzMcDTPgCxxQeUPLtU1mZBoPMI+kmIomgt5qKYhvV73CEGpGSyw/lHx
ttanIaEhJnWVPcUxZnd0qHO4mDiwtKAGaZi2F37hlyHUqVyDwalvw1fdlMnXPLd+Mr9zHE+eJhz6
Mr5Kj3iFnVKRIX+VdWfbWY27DwEuk3OhI64S5u8rSDklUf/WK8Eo3ay+YkL5JoWVgZB9PGiSx3qV
eef7+c4P2BAlok9jZamYiJj6t+eNDc/yIXjKgOEB65h3Wz2adCbdjetGUwr8X2APBKxQeS6/Tc6m
7ljszW7LRzYWLduUj9T3cfWqtymVTS5LuDOpeCIAFwJGopSIsfoPHvDTIv/YvFmpeheUBRKiMss0
BATCXfJRH82MdtKT9Q2/hC3biRyGMlpjzIAHFBRNRIsD451eeBHOGLI+IR7HSv9p/stvPbt7Et58
aGiy8jPYOekUJ/vwrzz1m/SNwuhdiFxgcsWt7FaOuVKerPsu+OpjFDUpJOTfiGG/azpIEajK1sVU
i+erc6fxFcdTtq6MLzjY8MnJl7uSIRicsnCQ6x4dQlOnbb025WvzfA90NbXMhVqhfIP63pWX4n8j
JvKHDnXG2rOY8t0c8J/eNtpr58zXJz+8FN8a64wX3ARZhYFOGa8pqJHR0QaOS8a70E0Azmt9h/ly
M3gdID+7flXBT2MUeX60QZA7pGaHxq5ODXiTBi3mZarFp8xDp5rjxnrm023f89k8jHqb/o0q2zrE
ARJw4NaE4CKFwCoMW9ruCfZXbK+E9FgqoU89tuZY9l6jW1nv3cmsGdJ4x4o1qNBT2ADPJPqNpKOM
D7oeKrMxcBvkDlKdrDOSNsxsaPAoQKvN4UJCBpZu6/3z4CeBR3uGb/J9qinV4AP8weYxZhimR5Gm
ud7MvgkmFWN+Q42mJb2c7KmC86Qs31DxImHEDd8kXVuKcW2WTpWhedOxcYCv3jwUpNBKLznG9jyx
T4k7/9l/F+uKi5ookTxINPYKiPeSziUMaPlb/Q38JdGEOLKGbvYOHUFg0ajGdxTItG3u0u4OyosX
EBa0KIuf7/C4BVvJSURArWyeO1MpYteeb8yAS+VzVNDBwZJnrakZRuGngN8+0srnpGtWSdlm0CDx
KbApAt0WJYwAw4V05tKPVPY5Uwxm9XosF7d2ckjA8YbTWSA3mxVRjgrJAs1WYQSr9TEaK/q6RMta
Wk8Ioyqv+VNxN3vAImq5f+/4LaI58s69Dbb3wqMBea8Fau1wIirlCdT62lCkkSEC7356PDzmDAwh
tq2q9MAc548K8AHaUo8TBHm2CBJlA7rKJujB6D5w0aMNGDBxL7a+G26bnAyI07Jhrr2LObAltgBr
9kUUaqnJz/0tVkzQLWxuEEGTIdivePp6NyO6v0lju7GFiui7DNfM6GT3DKAKVBL0/0B7qEqjKvpI
nLoWZdglyHZX7b+Zv2iridAK7SNUncQ9t6f2QTG080CMLsI5NypqaFP7ReCAL2n91+86oBITGGGA
IfAwfnBmJbVPW41JuktpN4AIVG/AZLqLRSN8iviBqNstuB4Bz5EduLqO5cEd8fMg3Tl0O1aiQEI2
XtqU0kl/jw0GDintjs6LKkb4eRBgEo41L5SiLyz//4fh0W8eziQinHXf5fS8eZ17ZrQqWqFKNQsW
BIsfJMkZkakDVwDgM56WcJwhknC3d4dFGZ59dPMfadMwukH8eDw94ryQl/xllMtFf1/rxhbet3Ug
RocYzSFSkkI4T0GK2Gb7ZiCItJNYssy2eMx8B7+2nkrwushfdICl2gBx9yf8euoNVF7MsEIPmIwI
S95WGah7He+qCwGKTXthTTXK6G9zstErJ0bJmUSkjtUO+ZcGrRHK82Rr+ZxYbleHg0UdbFS9EoK2
GjzBwIBLuOthUtvOJ1zNNJLEUCR2Rwe7U09ECogu22LRGYDOvNiHyir/UNylqI1CFgTFS2vyIHVe
lDHjtDoWCVgG2n4V/46bY/X91le8PWA+7l436PMTN+M2l9aHpgcwJnsVqclKBk/zNFNRQNV5Rm6M
oKuZCm/tvkbEB5ITb+ZjpD2j9okCD7ygPWcTTCVWAUbCXsJMy18LM97oNFA6Os/IP5SNmfdtr0jM
lb2blsucwcPhn2mH3iv4F43HEqpiuqbvq49R47elHQ37nUCJzSA0Z5kGuSxl5GJirduC7wKRwoJc
tTskNuSSTRxnAHQ8FgDz9R3iarvN9rsiubaBooc1TAbtbRKO8Gz3nysrzErHikhXUh4IedfaL1Dg
NDJlLm8sgCJIr4oNXbiS+/zHwBMlBJ9yinAU64tYKx/S40be6LKwq/4QKONnYTLzl/K+wQALFdpv
rD7z6CvVXdpql+9/Pfl0dfrgL+OqnyfCppwZe2QlGV/sMyo89YE1VG3Cnwe2fh8ChNMyiAF5eXXm
8XcoqcEXQT5OFKYHnDahziTBseKw6RiF6nM/32YusNtikDgocgchyycPYgvZUWUClHAh1JDNiTVE
6lDNjwTc9fupZg0SW2VFsLx61YpSrm0dlWD1FDhH3EwWWcOflj4QIEFPIX2Dg7mToo42HaqlRlYA
6JhEUaZVlW3zbmeoMOvKT44YpZyULcXFy8GHJwUth5dwP9J20nLE1TdUc33qLPZn9kHa1EDGetaI
bkzeruQ7nNFX4cNUvmFLBgI3y0XM+dLGbuwbIiNye20PxNkkVxvuxXvvTNNtZdGmX20N7AUG80zX
5KmTHkKrzDETSk38Z0WyK1wlW5916lcsrfrUlQNSdf8QW0uUChhz+9lZmoGtl0hziQWjbrrU2AHK
dS6AxbBN9kSFtA7bw9bigm68DI82/3LSPWdAmwUoVFZGnyFH1FWZhyP1Yr8thh2uDYu+2ilBLV/c
DAygHDYLfLxD1sZutb+C1WgrpNpAa951uDRTF5uSaxVNxiCjny2bezRMahr4kmuzPD8TOjucxeV0
OY+RW0xbCfFfib23FbALqBiME5n6ch3xdX6SaW8sXnZ/fhABHi/lOMI0+NsoCC7EKnA4e7t8UKYC
FxPIgEbWEcxN9s2ZY6QAlLsSlUm7MKzjirhT4CP4smrGkVfx4XmnZ6INbTDP+b8iuMU+rfH+j2S1
22ePAZD2tA61swH/spvbL6wrYaICLuv8CzhSIQlGn676LD1kUV9frC9129V0Ptrqp8qjIiA3lfHQ
I8ee10PW9u/qYK8DZmHndSDfy1JMtG4Rwtjj67Q0Qx0mPEMxZD4iMjamtxQXvI+pcg0tN/k73Suz
8q5Ppx9M4k/8sHQrkjHwQu4f8aQAaxpZoQcCTV5tE39e5kJfZ6t1yuAkeQxfwHYpRpxE+kl4MJzO
Xn/LC0CMId9ugtp/KUZ0NlgJi9Uorwy/okaa/IKuBG23hJL5A9oatGCKxrjo4DYkkeeLw0hKSajv
9tKqnMG2/C+f83WZHkjk5rXiCfjnVq6C3n62rG6BOiweStxSPWzfdX6f+nSv3Xl6lktZMZUdHlv2
ZO5Ijyw0lM61CDRw1PePBnn0KttoWVkUzTVS+VvaY24SvDfl47znm0O04k3lLHay/ueNP7DKLdQY
2VkldnRfAhG+gMdAlryP51hiCiUFSbO8Ilg1qeQduVAKnjQHQ+1O33DlVv5MMR7/fvBfIJYiv6Yn
YmJA5vPy6Iy9aWS97j3YCvjuhyMLoePdbeYKK9+Cb759Oj8oZvoY7VzxPSSGUeunAx1icgckt2/r
nA6cDTk0KLNba784qo82Ux2koxIAV3QEvIFbReDEzUCravxrnrH3EIK6TQdRky6ZvvD6bXJ7rOHT
WV7dL9VeGp9UGFHGaDhgeLJIW0suPEtfItJTQtXwIbZEjPCUfI8vm+denNYHfp78V5ulQR0P3DZ2
v9gHvOZiakq4R8BDbW1f8/FntVB+L7+WTPVrWY0wJwHxJd7H5nAnkKY43OyACd4ERIScZebzRzJB
nFTUdKlh0yywBWSWTWD9eXHy57h7lME9srpijQBDzmryJ67Pm33ThhD4qJyaLVMhI9lIdqcBnZsn
bvm9qs2OZyTO9qUrPYar79zqGchKdgQZ6p26q8+10iashk/uLaRZf3Tu4rIImMABUO9glbnIXy8x
E5CIqfdQyQixwxn1GSTcZBpV/CnYqcu8PoxsNlE6KFTiZVX8ykf+wWLbhmnoSgXQcYO8gX6A6lKT
XhmbR62sH5q4OTUnLETKrS7dPCJD1mz4B7mtImmbRUy5eB+LllDJLCINAwTbhqVGAXFA1CbGc1zh
ZcRQGFM/HAKhJPWixRr/45ValA14ZBQKYcfWOx1WzHSjVSebrbGdqTUZ8t+v7R1HchcD7rzH4k9Z
TWBda2m5DAJR1XWoAGYLdgIm9yhhiRjagVHU5+LnyPBI9LziLuHZHesiVpdpEbfVC+lYc8QEJ0Eg
JOZn6qoG/SNNdsSeyJ2a5ceaXJqK1UFy2j6OEu663/vagBm+53Z/muoU19+Yt/pWfouJ4pQukvsX
W6g7AX9hLSMFzlOAHFSPEjUqXDfA6y0oQi235CeWjhHAhCD0EUW6vnXq9twuUT+0tGKCe17JL8bX
/auRZCVmEjQfjP62W+Jqkz8o4Hq8PbcTfiqJVlSRWB4HBVNqHCkKtkeIs7Hq7D6HwwvofUga8c9e
uPRNtKJ0wavezF7uvG8mM4Rstj7E0cfIfGneaX2HoyHYZbX6WE9UOM7nXheOk27JUASXyM63IeJO
gBDYk3bO9w0HaFWPxwoMVa4wCvxrjG3u75oOyHkbzOdUFP77u7rfO5nrYh9MA/SEWSlEvKtO3HbZ
BUiBFActd5VmaDFCLwNMAYNe3taYs56dPQmfV3u7GjBqVcRriiM21rLUaknBG5QPtca+KRWktj7a
8rS/Fx3KBuNWfIPSmfnCAzpUz0raipCtO5Juh//e0956Lmr9xOHR5ea4fnG5GIyBDBIiHIuSpyW5
IA7N8mdFj5w3NfAEkDUCfU/Zd5WBrgaaEYy6dJtA705HU+zKb7BCQn9/MrnUFAh82w+n2hm0WL23
9ilApjeKBBx+jRfJj3DjquELZAaWoBFjnKfVMOmO5DcoHV9hni/Lk9P89vWT9jg19gXtEJoJdnEB
IOwmwuoRqthmVu03h2x8mIXi2RFKfbjHY/Q/a5/z804PCL5pwyA7NWTfA+2OdixZ9P0hqT6ebWDA
QW3n1AvNfvZDfrZHAkN6QOXYDiLfphmxUZP7v2kwyJWsz7IZieAtqO3j0r4IW9KJ8myBStnBToHd
lp/Zf04FrkyEjQp1akXhu5RV8TyLhcjOIMeIenQt6YmJxZR/bmg0/bvDUjAq7Jpru4bz5lTvmtz1
e5vZ4vNyJX0UQC0eiddBsYDh1+Vr/hG/4OI3IlAqjV+pwTDJzdqfSpg/ToD9mckWVvu3lAXiLOW8
oOxsfAFHuCrO3hyv3qC0mVW3jpMAKd9INcvcaT5z8NIyOaMHaW9bEqs66Wp0JOToh/Mx+lkb6y/M
q6oFISYY2rJr8wGebZ6OtmwR80bINGIycQUh6+mEEtlV0fch0coWYQ5ZXmYhPlThj2B/R5GkxlfR
3gFPHldHdvyDM8Anro1N2HNSjAOBHTczmpKXvIij1gFdnGICeSagliCYgH/HO9QTU4CBKABAmGI1
XAj8mAWRRVW8XbrP89Xyzn52TEazw9j8NtDIIi3MYrWeHY00Jdkb2x3xNy+llCi1R+asNf32cKTB
TJktDaSpd6RN3rG8Hp6wwwfghEHFZez3UuoNmuRBLQMWb5qZLQRxhM5fY6J2YeakeJQ7pZNGLEKX
xwqiRVh1XqFzn7oKFza0FcA6P62keNfA/2kfUPyiGTqRJMUcms3X5mFUmXSDykW4snd8TyrTXg9k
Jnb+nLgedDXMHCfe8WgCtPiyu/CckA877cb2uZ0+HbAk/psReW/KeYktLl0SHm/7WCgZJ2wZeshE
E8CW8ExtOQIXHc+wxYD/3e6uksnvmSoGpdnvqdgLbvH72ps+6XC5LUR46hL++WsVsOtBwQLPAmK+
D5Bch5iCBIs/LvMMb12pvsEuLxCMHziMQMoxRFhWQD4R7KWpD8IFjshySMcEgQCqUu8K/26lgPPW
ux6p4c7tq64okj/G2gMkkleF6uwTwra6kA0p+scb8pYDFuI+v4YkyrPShzaWhDk3eJH0FHPgouw0
ww3K22Ho3vntLLeEohy4UnQfBUzu8/HgbvC4j4Kb5oY5Hjrj9x5Hm2hSixynXl2vAUQdND90Wtlk
YOPjtTysxxbQVga8xv8s8jRhP6HTax9N/Wnwv76WVS1WMVHLNGHYYBn/MzQO9Dg4VIp95THcqdE4
1z1biRVZxJRvnS9ZDtRZe8qtPtQ2paONeZjHrZtdgpLSXG2gxIyEYeFSkFeR1DS2dg9u1mY+c7AO
OiaQ65vl0bPjo4YPmW8ec9sPO2NdWlT8daSxcOuNmfm3KGrR34EWxlmbzPNtwQH3HU2Ko2XXiZZK
fs6L6gk/cJqWRoElMIRUAdzDkV3Uz/N+AlGjyoACDg6mIs05+GrCF/nUBq9wixLSz/fBm8O3+14b
m435PT0A5Zo/Ox/hGyQMesKMxJcWLzhrUS+YCT4bXdXAPFzbkTXrf4KypvHO3JK8MkITg8Eav8QE
xZndmTue6hrwR4dB+EqjuT/2O+PME+LslriWTJm7tpl65EKK/X+35L6iYxwV9ld483XSXEAk8CUN
F6lTNt56x/J3wBEvOChCg05t64cROf6hg/hTBQV9Z8KuVy5WvJNfrzny/Voec6Q5sdQQOeCAfrKQ
n722IbNks8qyylZ8TVLexXDfWPemTxaohNxomDFioITigUTAsLABQ6G//K3CUZmuzJ580KWw7IaN
pHShjumz5A2lXoT00HBu5KikymFq6x/TharNDbE6aATV4gZ+IylQIZ7lm4Qxh7MY1UR23T/uZ/TS
dCfBWHOnT+M0M7j8yiLvF9hCMCxB975UEw7xM9JU6EE+SihvMoUm12s8p0BvZbtRj/cmW/0A8WBl
wdb8gMnhRNAoojSqDFwQQl+fvkR808Ws9kzGW2oB+m4huA51OHR004VnRNa/Su8SQizSxmg+/DVI
o6QpJU+N09Ny1fOvu/GcthtAgELFofBe9WVN8LrvNjRAeWwFSN9BdKh4RhoENZb0DGDjfaGGqT8b
Z+sewGMbkFet2sD9WL4IIFaF5ufjh1Lg6BGJYX5bF5zOKQEoo/2mauXoWxSv1YFadE68AYqlrN7w
nYwKGRSKPmzCFoPHmUYK4+MYowXT5B1R/uelvxNR42u4eCG9eUSYWIJAL8G7Kk7QzcIOn9lCFrly
UMeFrgzQdPE94pFjFQDCaFrYFh1amMiOK3vJHz0HJH0TBWigGIrG0FxMj5wtQA5+jLB9HPSue48V
5gHvQo73yBvKo3UULG54cwfyq4x/U2JgcrzofpgjZ94hxYLSbBFqzS8tlud/PGMCRXC3VDVYlTqu
MmE8ZZ5MP4kiWCASIO0WEzEWfnQT39+dTR9c/ElwU1GwJ9DrEwY1LtQvX8nv5PfntI9EmlD4EXtK
NWzVaZ/MazjXiU/EeuqPSecH6UoOHNfAcbvCzNc1xW9qMDC2YiMIXm3DVWzWDpELItERveYBdIrA
M4HuSCBLKwsnU5l3H86MkhDwuL+1VD9tLl2h/1J1da4bwi/Agb9U19JI1qv8cw7GQygHgySOfz42
j2OtwDyWfOv80b26EgduT9a9/IUjIhPU5i7wJY7T4bCgDzRBKt2uIb02QtyUurTbi54UqIMwQBs5
9ZI6TY5Lg0GRCDUijjneLTdg5nkdmot2f8QKUkYwes9/zeEYzeIJvLP/TkiBBFORW/62obpccW51
mjX5b0nQufFxqqppWvdBWDlv5Wbos1+pYm74q9iMCkvZTIUxzNKIeEOvPhBPrbpEv8jNb9X5HwRE
zYdMBguD82LS9lyyoBHre8d9FV8SaaWpfD+FVXOaLxp4ORYIuPlQ9BhtOn67/48HF9ciEztRyZrE
2SP4Axt+wY6spqR0UDu1tCe3bfRu+R6fx1IiFhBaRYaW4uYoKjFIk3f2OyfRvpbQq0cRntvqUvNf
KsLCBWFaPlVYHV+TcgBCpXkQeGmSDeOb7+CEgV+JrJRACp/+HTeKJl/idOhzlim1Wp3iOXyDah6C
Pz783+BnqkIWCjF7YW0rPVatmjZcwsrlyZss7LieU6CDDdpwwGaBUl402x4Rh7BbahERhUIXckkt
vIWFWpmycCk7Y0dR+K9z6A/BoHwNbMdTU4UiqLihv3YCbXPH5JVnSbyoFap4lCAgssyNTSrP61fn
Ho+3pX6jW6XRQgcYW6U4yu3GYtzCuI1ObYirp5pUwZWA6sVrtt1HfzmYfLvS1k2LJ8TyzOcFVOn6
HgZLP1HaK3dNa4UmDrbk4MUutYP98/PUfzpYWm96iWMgL0T8iufWtaAE1l/42dsYhOPEB3tdl1tW
BYnmzujyB6lmDXiE8KJxPPdIOjd15Fpz4hdB+GcFx19aQEXy4vZo/sWOmXpUp//XPi0AKJGsJR1M
KrZLtSIA7lIEWb3abQJC95JyoDruqSswiRh2PfBFbIv7N5ggx46o0bI/aWSjIQU1yOUdpddTUAa4
gdFdzGepRIWmGoX/9nFlfp8PjAsdT9enrvi0YXWVbT9vmU6yhrYW3fTasJ97vhvQZbrGxD7n8tQy
hdm2PbBKckEGdlUPBELj3x4jOLO/PyY74sCjQpJqY/DeNQJVjTLXxXan++bP4aFtHcoTnFKFsOAB
e4ev+EyN7rg8WAEYyoQjhJr0kK+IqpPMV3LUTUY5EFQnoU+PjKgRyMHQfu3aPG1tkbBfYyxfIIfJ
jujVN1Whpybs9RWGQro+5w4P95+6KgMwnZh5NivJj0z+4a5zGBSCbnaaOKKfIEtHYd1ca13HN+Xi
3sh/uE1d1w6yGrMXvRH7uwlvTI5AlQV5okeqIMo7HZ7upe7PEoMS0++Azlb4kmcdTCcp+uwVDpVR
bFZt58ztCCFV+5PL980v/FJ8RPX1vPtHtQn5CFs80sTQNSaQdbYIKLmeOB7HT/oId3EkugvGpHMl
K15D4M7BwKSZxM50CEhMy/+NLz7iG/x+/bD2fYRcAERw+q1NhYYTCNrvU4mFu+5To1Dg0VvLXEKb
bvULEU5vEmlQV8tnZuP9vVk43EVjUez+n5UQQfX0nQPL0fngdxClRvWVl0qYUD9jsDfXx+QdO2ia
qElDuLKPrRYReRhT+G32xjn/XxcxdGZj9HBMHZp0uWQOK6rPfgzkIlV9v0jiFL7HGhdJR5cEd5lS
/Zcm1b/na0F9VdQkNrRtYRpD+EwOxQNV/L+apt3MHX6Tr41F4z9HhOCJYddo+PiDZWm2T0C1Wy2m
bykr1sz4x9/dCjN367vbfMg8+IjldsHb4i+HeOftBpcQWIRHiWJtYjS7eb5KrmXgCtnmT/uuqqE8
YYEG5ZbYyIJqmdVHQdwrlqt3C7R+e9Cp+kvbXwrwY7zhcgWdAMiuYMmqjgMMqUn8BZwUrPgknuos
kQxworXjFWck9biUNNPVSNCfoBu2ojVFF3xBX7uUkXdKOZvnswG2uigyJoWhnLNRwNpOY1OazOm7
wDJncjUhSLOeoWtQhxLEdDQPnKUzwh7/z146sivlJxhMXaNuHfMbBTdmtpC9gh0rd1dQ1ee47wBD
px1A7Dfc1/VYKFpluQflxYTe/5xTd6uyyT4tlodiK5rhpUAN+GNj7v1qRyXeVAsT4npCgSP+T/lz
Ra9o908bDCN/a5d17Dx3ROH/JEzp8wI0o0cRAjUQYvm2VQHses6Ch2SzW5aELgUlw4IlzZKAZyOj
iM6C/noUqdlK2m1yFCF2eE4PGNEhWD0XlCzwAW1obiKz2EVZ9nIBSbGQPQHAFIfZ1im+CfjAnV2J
Ou0tHBuTF7PlPKmqeMPfh+l3VafwI7iao2qvEoyLnZ8FSibad+qJ4IiqcrhdYaV5D0PA5ox+e5ml
i3IIR7pGo4jXWSkbhIMSbHp/4KqhCN5SCogAxy3WhCoQ7K89UTwxjEBU8ikRavZZJdu/iqnpg3RE
qTXIXwBVAksHLqIgtRHhHKEPo5WF6CtZ3nYZQV0+kLzQLHgIohhkZfDHXETL8CpdzdkghZT1ffFM
cwEE+4GWuhdSb+23hYHCWYdN3Qw++LdEj6w+vSSpO2AL+RiUaGcIMNNu44iYeoDhJK8d73mXvSs/
ecYYeiV3j68Gjvotk3vWpSNVjokkN+n80+84lKU2gx20U9ur3Hq6NLgivZmzAnyjUwP6qzhcqFTm
rAk+wuZBvIf5roQ6YBHk33/1Y/MOwKY1K5l6qxwev3+lR4yxpQrYBfKvOIKyUBfdDr+WcChu4Hws
DiYrPF3gVhcTouAY9a3vfLL1eIxjNGpQznRvONl47UfqPcY4YQZep1QhlRgmDIYB/7yFVAviPIRW
pTpWQPBPckHd5wbRQjGGcdvxWolzIQ1ewdqRDjwB+u2ghLX498WBH/i4cVxUVg1xsZCCdDgHD0E+
al2zb+zZqqu8sNdNGXHwAiCTGAvzKUFo9PcXcXx/dqxF3/K/ecpvcvPMB214ZyaxRUUsp9aqhd16
1nwtff/KJoqDS1deX9D/Y6uLcYlEoWdeF6WeEogqnRp+JclZsmWj9j9bxZYMHSYIQJaNI2DMBGpu
R3eFBWKxt46GWVfhvL8RgbSDNKdfxAAke4Vu+ms242u4MeGdnq4+ytTL0fNBoiuXbyKALA+ve4an
0RvtN0c1iMIFRa9cYwnxd6D08Jqk3Q5HUtrNiiRR9Zyg/lEhqWhM+Zs5Rykurp2IigX7NTVkyYpH
0i36d8dlt7EthIBL+BmUhNz8jDFT988uI8uRarGGY4RYcsnch43YYh9EqyIfoS8eQTFaBEoIDX8j
fWiO2lpyTaNDI1WSICkr3VxAxB5Pl8Y5uX1RBB2dL+fqv0r26nueL2bOG+4VTd15Ewc4DWwYTOcf
XXJg5wNUry+7E8xG64aJXVgtauEBSnBERSDwp6LAVAHvt/9D0gk1b1RkqMdqBFYqqEGBtjyUoOKR
NATi7jEbnpvP7AoWigMmNlQF2Dq8bG4VsgdkNWdbv2pCuMKQyPwkIX9nqCSnT7C5e0MAdLduOAQS
a2Bpzdm6Hafza/yH9Z18sDeaGVTRj2qX5UdKZEqRWzhEJsWwEZEh1E4qJJY1nMW1RzrpKOGzCNjv
+PWl69ikzIkC71ET8C+0sikW05YgJ5UQrs223w7DjmyyTbi8pzI1/7EbP0fCUcXblX0hvi3RrhuJ
zq1213PEuKclMbRd1uBYKW9RnfvPtlTn77ksvU5yujZCLHj22d9tkh6561a+3kLR3oRcuvd8J8OR
JZg7XsHGGnyARsQdM2VN9QtJmpAU986bw+eZm1Vo1vZqjkxMM+PuurNbQAyVZpy5VXgE7Pj+YDMZ
R7XBY/bN7QdjSyDsuc+cmrybEgrYnPHeFr7CrJFdxWbZHvgKDcsxmJzDCpNvTmEECUEZ5o5c707V
jxHyMzz2mQ04DRasaUrpKaMnIjYcjTEsiWaMKXpQ99g29gHDFbMl2gDy9tPTp30lkc9sTptkuy6w
JXoeKQlS2VKj42p0cXr1aJkACz96z+I4+f8d9fanZtuf5SQkPsc42xiqxQea+6l+5MK8JhNqT1Qx
dfgLVqBoL4TyFYDMhHDNJXnfOqD6FGtGXmFh37ZEsAa8fbtOBcYricG5HZtQpKZ6D5DWHeQa/Zx7
yILvsnilNb9PhjUoSXGmeiXaV/ofiMt/Ev8c52MYpm9E8Hn3QgLvb27zfzFGk0f+D7l49UnMLdHv
j5xrwK+7NpP6PieYga9AJ78Fz4GrnULwKe2wTCxrD6sdVqUDltux5y/oYLNEB9lWN6tGVzIGj61U
JiXFgVeLpdbNi+TQyD/yIMuOxwDKgVsfELuAmrnt1SDeIsGkI4L153/MxC8uavczFMIsu36eAZjC
7C7QeAqNEoJCT9uUVcOe4h0D0F2X48ttoBoWijoSQJy1lDZWIPE+XRZoPHFceapH2mdSXqylbjWA
qm+XDIvCUDVcTJaMMHl4bPI/qBO1raE6mp1aoIqUbckZCRbxaYB3gPognt/N0bl8J+gBmNn2gfaO
74cqXaV2cAVUJq7QSpZNSS0O/hAjCLtJssoHjDU8sWUC1zNoVJ13W1s5TnJl+uXWpRMqYOnMA4Do
4MJmV0EpjZWnWp4mqGopezk1bGN/AeLr8Y2gCryl+WHuipRqsRMCVrPyCnYUeQVQwwLYptikqdiM
d2ZZJewv/vqQGp3XM75a2XXkGs9vlCkWngNLW4tLyB04lSM5oVvJ/Ku5J3iqnKDSzgnEk8lVMRUw
fSl6XHaHOgJt0uiXRcnJmhvjnWe5Rru4AsNBwWN77Qy5BrmAWV8TMPypPJwVUSVL1Fuz1sUlVzHl
egdOGlLnF0ExqNY69iT0hjZ2lP6fncMQ7Wsnjy61XgG07WxFiiyULvtht+u9pwZRtK/YA/Whq0ZH
2/tKkjA1cbFZKPAg8k9GOSo7kR1dr62zmxMdMvoeemT5B5pnCUuGVy3mneZINT9QpgVYMTv3Y93U
lZzE1yb3L2k7rf7czf3hHRZhXZLxbDaoIfIbJX1J1Zl9Dk6oKaf5pn5oFLMXZ+7gezUrwUwLozrW
kvzWt5U5e8HP2szwREeLABAMZ9z7DUHAcnV/WrbAplPkAkgxmYzNd1iDraY3PeETmtLJGIaHjUxe
tP4vSAwWzKebqmEU+8IfZHfa28W+FNoILtTtPoC+PssZw2h+OztQBAPtH318VezHWGJp9KxXfQgX
DgCSRCmrO37fXsEM7HRr9rCVhw1owKHKfPpY6C5eiGtrS1kdvpjW3Oy/qQjBhnjA7QV69fuA/fJu
FfS7s7eeJC2kmhDOAWAyd4boIAYWbnP9cG+sWOm542HGMA5XleVQY24dsc1BbkX3DYPXDGl3IayP
J/lxCj1tKYYeABzpKJcwhEbK2aA4XtoXihLdav5sxh892iWwA/4Ms13bQWbXwvKD61QjwoZZG9nk
w/hfDBz9eO3xj39keI+0r8NnNob60KgQPLTtygowDYGN+pMQiZw4+OhS0ifUpBT53UKO6fGpPD/k
F/WOs51XE314yCh46wvyn6xZkTPsjma9j8TcHqRYWSyP0GXMMEttA7PPcAuY9TRNBD7ATqjMvFSV
hyeFStkP0/24PNSh3ef15fWng9jnHFfzEFftuUWYqkbQe8mCnNg9jhdmANTGkLDCzUZwzA7z/exC
ae7TDjds5CSBMLDxQXKNhOv2eSRbYbPDJsAHhDtWtAvRju3cGKGKddSzUxgvvp0MIzecFz7+HKbD
WiRdHsnQpD8ADbb3643pWxmk2lJudrPgDyAeajyGTLkXPDLUVkiY1MmPRR3y/IcqLJczyxsPWNLf
I/nM0Z3aM3w/vLNCAJ6dFJ20nYBIZQ0gay+v33moQkGo54YjOX7XOTpeiYL7WADOpgdHH4ORnzxQ
x+QS1b9scr5sZvOk/nokrKO0bZD0MG5lndONiAquJK7pZw/UiiFbHqyPJL9RiP1wupz3Ci8SrOuM
2MPGDDRQd8qRU5m7UT/y2Wt7BH9WZxJCzWwTDRx6YZtjED3MSLJSLg6/H03RLfSYaJzD4v2WnDTf
68+ZpzQKjdY964tLM2e3ckZylFkrcoWejzP3vBYYtivAA0gErBIW4MKUA7COLZOFLMNdmpmUUYjW
lmGDHQPxrA/TWjaolOsKQmwToZEpQdHA+O1kVuNEiBhdeHqNG/Ub0VmS8kO2JowAd8j095t+gIPO
SfbCoSWA1maHktn47JwLaimxeiUmKWdXhGPci5MODji0CZiubENFWHk6x/xqgB6VyeUQt77Qy6Pz
xQRuAEt3QRbW7IQ+KpH+IMk9Dnu3kNtYdxKSVrBZDWNkp1cMoY+P0GwxVLQp8JYEzlcREK0bNfH1
mrmPScoLx/dYaByBGQ2gGxlcSQl0jq3Ha2fq4pHtA/wEP7BYbpAVab0W+pCNesmJPUp7AnQ0oSQN
QaGaqd4vDNytPhDp3w7pd8qFgOATgH+ta3g03Zc3quWN4zqYM8jGZVoMlxXrBkHyjZFoWHUi0yBx
AJjhq4FxlwixE6uU6Y7H/HK5tStYyQ6fLRIW0Uzo724Dj2EbmKBo9udH9yRMxj8qVFZisosvPFwW
x2IHQWklg2rtofGdsGQ0uXBD/0CDC/WkyMeCaxsErYf3SKmKwh7pOAkBjIfadZa3+OqabRZHNfN+
g0WcMIReOGOQtXffhApaJ8btgO0gncz4Ghyxct5cih8oJRyY6V5g9e3XmHAhWYW79ZCHui0kt2QJ
JeF2bDR9VeoGw4jbKT3u3fFQnUpbk0lKMvqoPPuXyLoEb+3oCQGRVB/xsZ4wecldd1W/nj2XdRk8
CQfV+yHNzQPCSELtRj8ASh5rPUr8A0NDDMT0AeOBA3leKO9+l0hvr3BOVDOGiFF6i/ZpJzo9tO9K
fNiI0HmQWxvIcZU=
`protect end_protected

