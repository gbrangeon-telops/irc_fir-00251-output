

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nnA1LvIFtXuhnEgnrDveU5DQhO4oCdS4/TzHWVjuSWRiJTWamPLe1zKRcIJ3OgsD949QJsbaygaN
jpuk7BYNZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cfy8I58fHjYLB4BFaw/VxzidETwabyuF6c2nxAde+hbLnyzOfkymKdOr4Pk5oDTY4htTgTDRWzMe
dytGdfmZXjp6SJIGysindi/Logxabu2rWzFmbsNC3Q0gro5se9+3qoriCL3M82gnhvX/joJNLiXg
rsFmmSylhS6v32W24xg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gu3bZVKL/oo3WMbeK5OSi9dLiGmyQy2yONRw6Nst9yei3DenlP6wnhfHYdkStFXi/uvWUBEeZ7hN
0Bmqlib8vQ0eJP09mki40prhGAwrKuqYt+2JunlvLYMjlmKGJOXPgQJfoYTNzbZDTWMAPlUaZkK1
oZkHNa3Wtk5m49sk7N6rE0lY6V2L8UfgTL/MmCwu7DKHNfTBd2W2KricGJ6ICGb/eh21T7mo+KTw
su5JPh2xN6VOnDqK2JFdz2Fe2UsNNdpq35qIZsc5dRna+xfhp64zhbzGUq3oNeTCYYFL7/rkWyjk
xMfq+Y7aGpW1qrNdKLCLUa3C0oRubzA+yEUHPg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CjIoJO7bPG0vgefcLg3HndCtGBfDCnGBCSVZItM/kv6K6ZpvJnvEpEF/v7GEKszxgiutC8bTrPRk
/jMI//klbN/ln/AMlW7lDqpJ5wXp83c77tloVq04bnPwc3DaApr08oK3Bf1H6JgBuFfaRFUfxoRB
6anIIq6YC6xrV65+910=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D/ZhWxzQ+2vaiYn3/fV/u9o/WEb/ogG/V9KccsPCOCWeaD6JXzbX1wTvk2mHL3gwIIjopxpeK8ct
Dd/kho1WYC462ZEZ1ijvlrdcQ6jRucbVeVK20vWFMC1CO9YW54zFCdUIFDYoBjMQnJ6IU90guAMg
K2P3LVnqKNh7XA5585Xm34QBVEtkbFVGa/nBjX2k27AaOcjv8CeFc7ihUp4B6D6YzM34GhHkOxNj
NyMvVJlZ5HBA7JHakPw8PSgdpMIr12xEOrEcLpR4AR6H6hPW9blh2XXVPneGey+XXrhV6WAB7P2G
TGbniILS+ojY57htkmkMwgWfAakIRm5HfiYkdw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4720)
`protect data_block
WRLw1DZLNLSLNXWWIegxO7YqYHIvv0t5LJvYw7psrtf5nuf1ixiqorvt3eosf2PLnmWL2OkBHqBa
FhWZ/pUfUX64jc12OHy58XOWBKIXsO1W6jzpydrfxUd00bN+vZhZDm9SEsKjv7Xs3JqqP8LEH8/o
ievr99lfvQph+FDNo95Wb9gm2uBc4QxaWJtTky6SssG2FLB3rzy+cpxWRFCs6WDsdW5QqgedWDAb
DecEM9p2F9HRPwQc8r0Xgg+8qtonZvsRLOZ20t74tBJ2dgshsfQczjT2rBgdOqD+6gZdrDTKHgaa
OlaF1bnsd7qTKP4PNrd+51bAdrvR88S0yCTYfrMJliUiQ855NONRIRbD7NYJsGduVylDpAcFGkAn
GgcOXUopPhubZvkuBHezlQzlA1q+Q+HxJgg5j1XM5XRfAK9Q5NmX6cJ9B2H6jOmKG1HyKt5jCNNK
arIpCRy2/4Pe7jk4Y8T6osbVEyr/+DcjH7aRe5IEiey4/sTOdtWraaBQPAq71Cv7kp5vgM6zGuRy
Akk0/FnxkOVljki5tbUALD8V/t+7ptTT5WCS8H2gqS8Lm/Jm+qQdbCQeHEg4mZ49gaOlSD1Wxygb
pi5AwtKgGWdnP1HnBTpwVJpx0zD1ZYq2VQeH++mY4jsIsN2RTQpIGP14tB98B2Bw6NKFMBSs3Som
ZCngfRoi7RBmyHWUkZoq1m8GUjIY/EjmsFwgcNaEv/w57/GNMj5j4Bar0tp/8vHXQB1zjuKL7ttP
PRzCebL2H2SbhYiYYu9oMjXXGCPnBUa7+S92YpA3S27NyqRsK45ZSdrbvO8hRLNTb0LbGtjZ+5MZ
z24Xn9Pcol9qZf0xpsQCRbnuSf3Tb0Rt0/NsATIOl3jnq6KkLirirAqC35TjVNsDWKiVbUL8hWU6
95QXglci8lc6b2qahAiZ+R9q+3uDlbSf29/VhsH0cVOo/vWLTWWjiLxkb+58y/EX3LCN3O61tPEp
N0Aqd2aUB1f9oD1/WbFsGfTewN4RzaqHOUIW722fU6nYaBrYUMJOpPT9Tw0V2tkFL2pS/CY5CBSJ
gXPQpxpZNBfKznWcAXU3z64SZnIbQ7rMFE+JUkdyhoxCh2P3WCZD4EF1c1XtYkggQhoQcoDr08rx
uxWAfoc70k9i9IW/CGwjAfB9ETHiA8fE6FpirguVw+7+6LXusiCiPOH0rB8+foeZvhpcKsdA8AWG
Mm+B+L75WwLidcXD2lS30SWUKoQShRzC+KQmoJEg5c/Z8Xbedpx5yeqm7C0I+iDdwnVWn1rZn8rH
DUK9Y6NiFjn+COlQx2Xklg1KgCzpOUHEa36dVisTraeHKICE2uMYsxNkhR+R3REPx/Zw01rRMiH3
iXBHta7yQsjqO3CzmQopFyBNi9cEmt1Pt8xxLryX39OAQQX6UlTFDUavlkrQKU1ucSPjzexbd+L/
QbsQXEng+Mbd8Om9U421NDbwIDv53iwJ/Vhxsoly7RtHIUOQLCJh56lnYrHmFvBwFVVeGQYmwECj
yTZ0POoMSU9lAIAY5+7QeYiWl4ZJRwEGBfq2oJCzItXXmo60jWr1G546uN7OI8C/mCjv0ZOWwxO4
wX/fEok3V4IG6uM6oZFNECZAUD9En90CoAK/HDsb73XCYTdBoghMRYj+5z7Z/uVEdxuiLLEcBgsx
rKa4ALkJBcqays4QZ/rb6tSqsEgM6kSfgiod+kJYu+mWa9wRyTHIO+x8qudhevX194U5vVhr9OZ/
4Kh+bTPoI3h+0+ckRD/Sh7h253eTFQOXl51EDXfReHFwbZtGwdlvGwsOEm0WkRqbsFhH/Fn+7n1J
vfadogiU4GOkOMm5JB5+ZT8V9P/o80CeZZdMZC+o1Kd9x4jRGOwMCTgbLxm/7idL/gQqYHLuqfGM
nPyiwTrDMHW7lDn2Ed9UNYuNBPCYHndsowQmEF7Y9PNGinv8MxpnuONcvKXKQcrj+AyTlY8FTW0Z
z/WivktzTBJ+DnVv8KuefxakCc7gAGI/Li5pfSIq5HQ8mu91nGWt3zjphwLoM3vLYdc64my9fmiy
A/b5NxeJSq6dMKoXe+NrpWVOoiTAO+jwXPAv9WfF8Y+fYhEi635SnCRPsd59P5S09+mJdgNs7bZl
+pwF8qPkul7X6i/E+kX2nJLiU8hnTRY+0EEKyEyyNxzTU4IwaCxZMrNhyrJBsC0bJZZD1aQ7EPqy
FUI5g9kBbl4euAlXO6feIY5QwX1b1d/hjsleesAnALJOgQ/Uw7ORaCUophMz3ydjuDOwI+4+aQP7
nDDH7+ZgIpa2zUHOy/eUmVZFleey6TFdOTYomf/0c2woKyiUZGkNKLqawzHtysbi46Hr0igD+1mM
gYITMIIKXQhz/0ayFtAz2xrhQcBfQ5Ti/00c+JHoJXnz9PgKn7PGfUIkbyiiH0IJ+FdVmRNlTINk
mR8J+TLxyNU1vMa3Me6CXRJC6gwEt1/zH1FROU/FTdGOjJfRz9JX6RquGvZCiWmqNr6yUI26/5DZ
SArjzoaDe4xaY9h54F2z4XmfmUPTOOKUOvFSp9N8sCc3hCPlRQmcMjvRCJ+FERAp16p2etaLp7EG
pbsWjJU4NyGULDk6z3NwZOsbNGe31PVJUyoBiEuqPTFiqdfSJ7DyP7/KgC3KEneELcrweFmVQHNA
QtvgHK/i5Qay6ktUJiWUKKMlRR/mtKC+6pZ4XhjS8zGYaC/gWKNRoCkx/FOITRau0uic+1eWmU5Y
XCN/2DbQlalB3jzPAAPEqK6bJhTF4fc9RAQVESn8zXTnf2C0+8O8MHrREorLlVEDG533M5FcD4dl
R+fzcBXKwXC6UHcXYD1kZeXDpojqqMDkH2TAsSs5CIOp2fUqupFoBEZV/U9n9byBaQO14S6DNzBt
lJLCKjsMAXGVDuvZXQDi+OvtHUAiTlYYYCEFTqs0IWUm5PMSKv+xZmjPArZw+hPJxu7m4LXB5LHq
wcygKRPyiWJNyLz0bHfWayx4vWZrlWZDXAnEFOJPhSnKEd6rDNs9PcH18FZC610olSN3ev+MAYga
OfXwIbsU3rQuEPsf+WY/WdtJwXdl9evEYEmjtT+H04jUsAhuNyFha6DRlcWB06hUCRfjsPmC6pLu
ulEMXtaECP+1u6Ww6TwZS51G9mH9jIQ4fMRrZbMqLnpaMk6Mpl64Y/1adQodmquIuxhj9I6zasuA
uJJ/0oMRqK96UWekgxLU3ljV6/+HoiDCFq6mtunDUN1155eQCDLMr4x1tgeOpLERQaloGkpS8jkj
H/FzFdRs0ONVsxIkuLvwCYuuiufoucP9jn/mV3kasuWyCR50QT8sVxynzBjk8GzkgPEFb7LJDdGb
LOcBMKdlXvauO7ONvj76MeSRzmJHdzWhCqZ4rVBqQUI3JPZag5fiK0VAB8utvWUgL7IDkDxlHyoM
6lN3w6msX96beEO04+VBi95pMJYEvfKpkI/6TvEjMwlx/03j+OIThK9DKa7FyFwtGbxt94XRyonn
gpBM4pC2nxwu76WnSVUVl4T6O7wseb/qqa+IvidZMv53Pmt1FBKckgWBPGnqzvQ+OrPC3FDZFe9S
DvTBAmfEapwO94T3mxDovIhd7YaGhva84DSE0/SJIdtzX98YneKPMMp/0Sc8vgItN2pdlJQsaoWE
3gH3paUoEciFRvUYrf8bsjV2edT+dhejhS3faJRDLHdI/AR4LSN8sNL2FbdiVHb00j5rj/3b2aU9
FYB50DNMtwAEKsmzmIlWPgdqLJmz4yRIhfNFF8gvrL+zcFET3dOXbWYTqOVz1P+YdOMWyMi0OHYk
c2LMBgsEnGhYn4o763bLsULwcRqbDioibdJlc2wCn/hX1ZKaUA6GIL8PUr10Tk60aV+k2NMd2ZJE
o2p8LmDmuucqRhtDREFy5nO41jFG+6TS3uP2VFkbQwT6QTqtTeB3XhxeJoKqZZNpQrV1RJfN3Iab
NhcrcHrIC3mbf0ozFea4HR7sqPtJVrfJTj87cp2A1jJCVhgY2sAMI+E1BWSpT+XD2CvfYcnyOOoF
Iyvm0O7KiYxTRMHIGfseKN0JP2VfB+Yn1U7C4SzhzzsRtVyQUN9gIGDE4FLFnB0lFGxojYxivMwI
mlGMQE8zvkUbhINgHBZEE1G6Rk1fDTt6GXdsi4uwr90hbTvo/yRU7y+QZavmd4sq0cNjzuMRfbas
fZNxu1Pne1HS04i+Xsq9nUi+vnEuAqr+2oltH1wAa5AlX/Crg5Gjw3MewjoPBLOBTPWhngLxvLTS
k501iqLYSzV/Zz5AyEQpHwkiTPS5MzQQurtiph9WcKGGrtH7sTVwWnTi/piVdIKSe83DUzj5hh0G
HShepKRNT90UlhmGZGArmQJivQQ+8mSDzg5FRXtYvIP/DFxhZrVhM1am9yJ0dBLEw3fm5XcnnA88
lyi1+JYXaVjhgPAr1aE/NzeRq8vC3MJmNbwE8nUeyfdkaTtRzHPtBq2bbwsUyot8BPVE5H4DdNJm
MC6RHWAUV9CgU051NKXQWnSBrRj9I+yi2D66i9oHpe926q5YfwSvYefT04JpKUBZFLB1dsqaw7WB
aXVhYs9xqqab/y6VyXfYMEpssfVrdOiYNAH02Ir8udaeEPk0uBass0Fyz2/vFfuNHrGh22yWCf7H
aj4bkgOd8j6nA5kjUx7T7Msav0rd2plavwFfiuaFJUda7An8eEalV+pKxEALVM7PPf89kuhc4ttX
I0tRE2QQRIQ0fS+VEdraFqhpChZWSrfII3JV+tzh8beEBpJAymcCcK8WdJ2OqAMcpzI5vz9PJGB8
IOeFH1WgEYEtQgYVa9rkAid2hJWZ+e0ZzATjYrr0yqB2DLoDNW3U2QW56fWJYGxFE7curwSmtwio
veoXhZ5Erli0LDBdqYdY3gNJXuk3jzX5Qt3lFgL7U1uE8U2ZeeB5FiU3lZg5dj7qZgoqmaaVCUqZ
tBZyrpVg4UK81auAWF9mzoDLcdaQW6lmJlRlCenP3VAgCKj2ChtwGLCDGkyOZIvH4cTDXJuRClN+
VIr2L+HuM50pOvpVN8+32m7AA6HIwV7lcd3vSl5AX29e1la3KRr/acG+vmDw/Wpjen25V9qnn/mi
/2ZS0QXmdTGN/8ONAO/h1NHoI5/sYuPCYpGrpnQybEeSoHijMhk1qo5rQHY/AX04DtpYfLsGXht/
ui925Z+tQTsckfFUv4300LrJDDZbkepVnX0dObppTYlZZSWv84c7b+4Iispho1k747/T0iPCOKbC
7lnKI88+wajrh+nszTr8FAnWAukEbK6EH3eE+AoQuUfdxPrYm9nmViYtp1KqY/PIR0iF7F4lO7ga
ZxC+TRwqMAxBtsdSIuCGpnmRq8TamRlx8Nje3EWx7yQy4np9OzGDBQdkbDfGAcsNi05jkaxBx5uc
C+YAWndJdMLI0ChscGoi8e/RqMYFBJgDvKPfr/gvRsSmdqRLsab8B2uCNcyD4ll5O8ysNhlOPoSo
mu5/LsQn1wuL5P0qsg6q8KEio5a/Vqsq0akVZC+fbJvSXeGJpOwhoeo9oCZ3P9/D7ECXh/x/p8ah
y0RnT0Ncq+KW8wwPo3V3z6+0s2e3sLO8j0+uc0HtGeuOFMGV9Ss4qZ3NtZZdXhJjiKg/+OXsC8n/
24cHnHHTTaRq+qPjoh4wGtyT8TplL5VfG+8kkyl/xR0d1hYdkzWfwH21QPP/lp+FxG3C2Du4kLhe
E1KZXOhk8xn0Ta/9D7rkhpH5VbL6maD8PtTj4oyGKkHMBOQ6zY5d36CQoYrO/yCOo7qY7naPlHxg
Hs/fAu53cowRKiO6Sy23PinRVXCDsrFcR9ORmXOAOVMs0yMsa5Uo2nUD9oh6U9Fx0bX7BAZl19EP
U/SBWJK8uj9XPy9Y5C3BBgqxKpydHwgS78Liirz8L1EsITFH78yYIcukGDjd2FPBJu2MrdX4QiMV
gJZmj+cnRiNYVhIaq2RNHaWvv2VShnmTtjJ4F3+/x9LwlSvcWeBbpVOAxwREp2wA5M3Yg0KufuIy
j3wERfXW4f+gJf+BZlTjedr3eABV9o+7nuxtLOel5Mb+kl5Q3V26DHRa13ueDrjKHMBfLkekK0EB
4+qNaBsTYgPlDppv/pcLlso7fhTekYLPVNYIFC8wwBYsbjJMEIciE5e/aLjNgp/3aGcnS3ApxG4n
SSVfiSDEbDqjmM6WMqO2lXrWFUZUZo6olzeah9FNNX8Hul10/WOiHKt2+yorfB6ylhxCctUOdzcl
sdh82oAXUdR/T3N9FmEQyr6vLogsiZrECRJWjvs9EABxgAt0ZWaYSGy0MCldTg==
`protect end_protected

