

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CJc8rmbxQK7PiD9FE9h/V8z28Q2yjtwOLUGOHj92X0D4bGhAiTKxH6Gs6WbTk3x8dF6WKWHXW0Xd
imaqryWs/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KUGgnJN/sGLwh1pfD6BBRkJkdz3qYXsMmFAG0D8TIT3kvn1DM/WYFdJfNjuI3TZJ+GjJhgQt/TQj
vszszvccproNtKL+iK2kDAI+dODbmK/3dk8pZpjNIY8iqG+SZd4LOHkCbGnDn8J5L1SCb1FbgOpc
lYLzGKyKMfpMp2H5zrU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QPilQnlZ7SkqHJ+uQKxasOWlKPf9SmSQp0r8PPqOPGeQK2aUl+9gzicjiy17/DdQAM7rwf++nyUV
Yi5HrcGStcw9bK+k96zmiNT/NPvXPX5xeKvpNagObga/il62MarkWpibvt8B7D5IQi80Rp8/xMyy
QM6+TtOf7NVahw7dZAUwr3krfROulZTDfEY3oalO/PlnwAGr4Z3udXzac9NTOUWxkjpW4cmTbWcJ
unHhHJbyMO341XtwkTUgKReezgKFOpi+gREeBT80YOKcPQyjGyGuc28HYVmxKisVh5P7BYL5neLX
P5GVK+HA7MCB8DsbsorDqal6rxwDeaIF/kJcyg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZE3LPHWjt8FXIcLXD6pONgldgtzqHVcVbUx4Qj9ztf/3D9DwoYFB/m8dT7Cv2OabvKVMu13QC5lB
rxR5Jhd+fouVouDNKYwIESeS4DEkgnwfSJpsmeVaPW2tqCd21tzGTVfcw3Igam9PcTjnI1q1568h
X1Tcmu9paLkGRwvQeII=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EV5YorhH0risCTPPpyQGO+wsA9egdTVjrRAwQuEDG89jVsb2NsTih5Y+XoLrashGMO3AtQzajDhF
KB2YGM3JfNSzKu3jU5R247s9Goe6ZA8J4KFFzdwq4blriCHlPX0eNqXwJaOF7SeF++njAnDs0TkW
tSOb3VJRRI43LgFv/CHX80X62oIhRm2LIRAjPrPj7KevSjFw7diU9sSURAffWyrhgq3XZsUY6ovy
nAWzeDeWY3xrRDkxjxQAN8xOlyfUxlNsf7am6Prp3DCG9ANkw/MCyfCVBJXBbghP4T6GS/pNjySW
+j4cMtiThQqIcJCHVcAXQA0FAf6PbH456gYJfg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4624)
`protect data_block
pXbYHvxJQCyCOEYzIbdeR49xruAuu5v3VsNBtp/nXdoC23YI7YyffZjCw8sbmNNqko1YIV+sl0E1
4szBcKZh6N7mrDbDtukjpxYyk67x0PC5wjysvQrFGKT9c1C+ikhBsnjxX2tyUoGo9b6yoN549JHf
NoaqrHl9FXx4aJYq7xW9ivVCPXo840z5ZpOqER8oWmyGs0H+zKgbWkdVp7XnrHyZBp8e8ngkH0QD
GV2WSB3iPhmuI2Gxd6y5gihOhLGVK7Q/NvHoo69PWkHn1uXRturkcIazVvQWOj2w+HA6152tpw1m
wpcl7nB5jrgQ4poFVv+I4v20KNbv/jA09wfL2Wp/2qNy+wnXut+kk17Zfl6T4yHo22coWY2Jhhtd
tK3LbplFY2SpFTUnPuVM+YRdvDomkj1D45Whmaio2Ftd7IoErTtjDAGN7VKmaDkJeo45FcFD8jfn
Hck48HYry+uzQUgwfC8vEFvMQmlEzvfzTVP8dZ/oXBItmwmy6CGv6NJBJM1iQYUviBg02fk1rp6s
CTqU42S3ZzZ+jMYy+DR7WImkIZ5IdxEWn2SVZRNCo47Q4TlHnbYkujR/uYoG1heV6wwOks7pTRb4
FgoNWJTV9V2pPt2HsFCZgTvlck2sYsLN8aH8Ha2t2M6X2baPkjO93j+9Dx+tO9h34WOM04Wig/x9
9YQxd/dwSJYYgZEcBB1JRjQkn+aUxeL3cvS4giu1PkdsMbaccVstkzVnDwnFaYtRTWF+JmssnHBi
9m1Vht0oP1Wo8S704kt8pkI97iyPKIlH3ntcu0LzIr031ypTrp/XePJKvveiQBcnFDnLl5I8ETVy
p1JzZZu+JmCoWCFfH8rWBJ/PpIJXfXY4f7s0he2xXNNV9UULEV53RS5S7X8b3pYeL/9LzfNqvrlp
pQnWfYK82+4+xkJGJOZ7QEc1Eep4UseVAhrSPqrQmkTB0cvniQCSELV8bsUN1zqN8xjeorDlEYkr
d3icVAgfwQ1juCi76xQk9684jBZl7Vvbf9++uFFdFyimW4434VNyf7wMKjgc9rhogxtDztYAULnl
g3YISGV/n4csLILwRggOQINu8iNozeo2t/DtzBkaxNkB9VSIbUxCseRkzRUnbfptXsnyL7zWJfBQ
ztXc6B+TldexoPPUsQtV0/ej+QnJwO0LPGzVuSTqIig0veMjx3RxzeLw1YsJ9tQQdjPOdqKLZu76
kHAcd3UNW/tx6mG5CtRzzipck615S3KZftD0+6sCsVxKX8icPwsT5sZQwDIocpxyg1zxkb+Fxqon
B3cUjHlmPYnjJJ0UpjAJknjNnMVL2UspErRO8gPB9ZYjgEvse66oUSSRiehhk8EayeWB8MYgSdEF
7/KC5TPh5yqvD67zSi7Zd/ubiS9/OdkZQ3Z1R4YVtHlqQJJQvE+umvZ1hVAMv/8w3M0ijj4OC7M6
C8zA0eArfqw9KDoGjj03n7FmxnPj641ljuDgeZxsDypiCMhk4qFQqljXntHXZXSPWjYdPE6YsOYo
ffLSSN3rMjkiDDKoViyyO7XEX8Ef11nzPCIyFHrMSl9dpY/+C+9GNVJfN9fh8wghmwWaD9bUsnO6
dD7x30vdn6SW5qZxa6GXWCyQbSo2xFoW+nz3zIYiPJxgoAXSvAvgnIIJOJGfGdUowrF2mvB67MH6
WTx2L0OmGHW+GT5O5bf9VMK2yEcx9eV8ethyaD/CoQyHVv6K/dv+xQ90Vs1+NBpfHPztYwE+2mdo
J98Q0u8TDAIDQAWnwnPh8126JY1WGHGc8iv7w9pEdXPqgrF/4gPoAv/WbqEB3AhR9+79sZEbCC4G
xyqSuulKprclvljzLNq5m2sQnwbgwYX794NLoNxxm1TDmKZeQQB4ETMZr5P7fI/UC35DNcpo4V4E
wQD9JWlpqDihaFnxwA/KpXx6Mgm8w24PAUHRPTFPv+sdeLdzAgMtCdPqelUxgb8L2G9bPtXZIrJl
/WOYdsax3H0uMWHFzeGz5rSZb3yzG2FL4P4Q4JvSRO3n/bAHDklb+ZYqWYQ5wbHhDixZfPcFf/W9
wrVXuU6pNbHsy29KceV61e4ft6QfoQ9pkr2xOBPNzd9eQ9lbzk55rxb3O4thI59MER0yQLCvYxjt
gTd6Re68IrUwLHSCGzQMZutpyfdHaYLBsXJ5PTog8Xs/34BkOXVoAKERqeShBQUdcgFV9d1KyBBZ
yIORD/2zbbcfeLNW8RF6MWHQknCGIpFm1bKkV+qGbgP3W8P5pjLeJFf1nPuZMGaSomeB8ec35wfX
xESqcIMmGCbP28r41A9wUzfWa//yC/OvjXtG7Igypn8/04djbCRTEVTWLKGWL/DjlGPEGoWSK/zb
SeOPs1KrkDia0eX+GesQ18TrIuOLVly2YjS5RUCkCCiEUIQz6oj8JCZuOrFDtuHX56NM2NoifOOo
QgamOAjM2Q/cPXiwVPvgF80C3dCl6O3N4k6C9dPSsHtW1U/JKMtzKbKxkxQUfSW9+iBRaltmiMYj
Fs8r/O4WYQL6HbdnR9wWTfaSiT8MGfxPbWKgEKKIonfQip7f/NUZxPT0bfMrvpHf5xYiuXgFlZ5c
yayfubDUFou/EZXza+ACpKH8FIEuAW1e7vUvJ7tOg0RjonD2SWlbMf5GzpomwrhdJ1jaz1YC8egn
ceOEC6G8dCJiSHkRL8sJX6kQ2rktufMStwioamlNA/1kXpnUCkVdabfR6oFq/aRaZV0xc7uWJikO
h6kigv04EkvsoB2ktPcfNqxT9c7NMteGWJo925gsVsxQH0S6zqB402NUFUI9n74voCQ2Jymnny0T
aUfai2SLe9HtiqDRd/oGGlJglUcYV2zF7uHuB5DcfRD3M552fuuCFGcYo5un/7lV1k7U7JMkf0DL
myswXSa/PFSUyn0PwNsoChlXkAf12/UAko5sQtEfgFvnMwR509kmHghINJee49HJ34CzvMw/plBh
Rhj20l3nSQ94q1SxErQtZTsy84tDM5toRX4pTR3/KRV4be7PXaovusTXcBkhBBozGRoq6bBPUlsz
r80Weg0eC1zIOH2/imlJdfFVR4Hc9qrxp0tenH+ZXH04qERVNr4/1zKzzyttrEKae53wtnml6rYw
95yXymig27d77d+137YEuCBOiZUKcUHzr0Z3shFzNHpGWXQ+xnWG7WBKFhKC3lYL2DqPBbf6ekHY
DZHiGfSDn4u2dlpIs41saxZLOEgzz1SB8CnT4wtLtfI4k0Rp+QuK6/jF0yInJMNl3H1DQHVlwf05
+WRB5t6xCpTnpeIIAgTdSVpo1fE35QFxgha4cZy+OG2gM3PHr/U4nxDwEb8ZF2Y3C9QhR6txW43u
mQtUxzzb2tUyYehbgspxwoCkl+PsfZMbTCmgQ7BYlp1wsoQThlmmfPxdIvtksK6iYounNQaAlVkD
0VQYY5DlD12vv0zLfRItbg7F8GbNpLSQqSdlat5YyFa/zERTrb3P0JIxW+yX/cKQ08yhrbLBirR+
hjPFWFcr63jqOwfDwFXFuTtK6Q0Hlh6U8SLw7EhhiggAzGZoTqDuyGkmtoVL7iSkwHNrifEAotT0
OSsaKqpVxmvAwyUSlghPNk7x5lsSVW83Gsk6j4gdqb7BQfwbKRGsYnWQ2Zj79YaecouMaa4YyQtz
CHrn/CWs6U0ualKiLOCGUrAVQ2TKvvBFeUkZjhVqBPyzNicXWkGGaCunbpklesEN+Y4t9qEi6ch3
8JfBNXwSZKEKZbCdRKozM9lIauJjP2ek2MLV+cNH/dQnGUKvZ8o9gNHEvWcjNjynRtZD5Kh4UhLw
mrbhgiV7FvXV9l+Qb8uqZlgrWHhnk2JILpJvRAKhz8nQw5LKN2vpQE5L+b90yEWhng5oSvukjkoP
0u7gPIqpm4E2pPxNxFh2C22RfUqVkRSnEN/owAkCfscQ6hSjMtB83VgdpkSdspTYJ3rohNoK0gNd
rnCqhLdpQceSb1+R7B+8O45EJ7sGh8cnrPjy4xFDyjdENtahZUx/HyjBVbhECKc/1+OcJfjMAU2F
jTQt8O/7XHYfg1MWCW3V7Vl2FQVl6QZcaP7C8uOyEyoqxdEkIiP8g3NPiC+yYhaiBgBSKVtJ11Lw
G0dJpGbN+xSlZWfKwonqIWHLKnp2kHktfrazYQLipDC2Z1rC44qjcHxFbDTBybssChsKk2/8Kd0B
3yxITfeG6arTE55Oifdy56qRd1yh48c6t2BPGL94oBh0FYks6hg+lhiQ7mF0WUNaxeOoat5YmIUt
6RdD4/jnyHg7uW53dklaWEmGHTzXEcoiITNNJ9LH+rtZgMnwt7MDUNtWqN6B7ScHdSt05rC8aLnT
679qx36Ye/qrWFDzTqhlztVFks3P2H8Bs7qgXmejkgV4GBezQKyCAqmQ0Woq9pIkF0RM+zP2RCM9
UpSj6M5KoQfXi8YkuIWnufsMMCMyM2Q1/7iO7BAW+MqI70zTI2WLznvFmnuWqn/9XdQXCPqleX9i
zsI3LDhFhyx3W4jPSmaU4vJhXl1dahLa3MhfCe8GJ5L8tZkZMfWlXK5t8bnd0FQKomtshf0PvzuC
mXUzFgd9Hj0YtuWlrMFAubiCF+er3BZOotjwGuziA6ZmL+Cok+V3F+mT14F5IMdahuOr8+VoIcqi
Ch+Sck4EHssovlb9RXLvZWuGLlnZGMfx3s8RNdCjUw9EF97FyxHgsXYjKNDUYQJSMb3akS7TsbI/
X7iH1x6xP97S9G8+5YzHUp0JhZnohMGLoLAB1BCPjS4HJOivzL8Vm/yYoqObg2uWZhzWRJ8gy1Oi
ZiYLgXTgdnbemXMnYp70J28v97BVm7srIHJ0ibLI/8uEJkC6AUWYXp4o/rWVVVWMwoVUwnSWKCeE
Z5jmzEIhEP0ctYACDljkrdE7HN/z/PuM6WwtyYTWrEkTNMAb/9cZ4T1RS4ZMB/zA/ym+N58Ma7IN
HRdjJWipgDIJA8ftJOe2cQgr/P4WPmhtzFfGSFWr/yowvkmycm4joQXLmIOxy4t659Foa57c/zc2
/7tjDkP8//t72SXSS5j9T88IQbj3Oz46kvKNdTET0s5cCNIRayiXvRbpp7KR8exv2NTKnt1pQD45
MjSEy+10jXarOAOmdU4NZHw+h/RNNwDp3XDaMG1I1wJqpeC/p37M2ZnNTLgXcXjx4jaytvkOKnMV
QywhlKqQXrZO09WANiaujRP2beuZlEc9EQ+5eMaJiCzmznlN/HuB7wtFZU18mbpOiXzTol+ft5yO
/oZWtRol/SSaasUBnrdik4hy1Ndm6rBu31e0SB8fEm4LgUldlYNCtsDkmIgtZm/XZNkoARtlVhcG
GayLGXM3H489sJFMzh0xIFA+RcKhxcnw9pm1YfF6aANys9ETeNTkWKXF4ebZi096K7HzHBYA0btg
gHxRw1BSxod8AlXSQsT+WSf60bwga/i0eA6oOuwjGyTov+j/1ukxG9gq5y9a/nvo6HzDZybWjGVh
LyfyuvitdkHQtBpxN+voQa/w+6WeZvdls3vJ8ILnEYoD1kaQlr1dnZG8Vtq6z41S5vr1ahUDr/Oi
idMWs+kVLgV5StmK8DX3dVBp4auGIJKKsRSI08EFttZRnKvCMilSGnY/SVlJ3TgNpKB6VQLVm9X+
4+QdHJlZQ9i5ATmxFWkExV3N44HG0ClhexdhE1yw91XWZQXnsFbugrtLUhpVABCiFY0mvqFHQTBm
aR47l9M6MeeuItpaoHsFaMp7YDkDHGq++9hPBy/vqs6NiLbzdHqwKaGWnEICgMWiXig+H5chKqgw
KCx7/9OL6lfGGc6Ebp3rqAkKnK0zzoe/T2y4domfCTa0EITX7s6hkUJiYfJNYEtoZgRw1ctjaiUR
M78eAw1HQj15v51SlAuBU5nGkgeInzu9O+oH4bfIWY+S0bY4EgEJgQFjhMiE33V9f6RjacuuIEQE
B8vGbfMFIdUvS3ceXDpDmw/PHI8F5nP7EHgEwzKxzuypuN6FoGU6NQM1FGY3WKeBJpibkGWgnALy
jXqdIlF7Hz43Bp+lAibeyvgSgLEbHtfpzxnwpZ5cYxxE+u352RqxZsiILNY7qMkQqntUaZdh/8uP
E69EMzzFf/8jIhIwBKzxiFrfHdLL9V2Yt++KbxJ0t1ydJCIBieaBmQYsaWWloz9KojIHX+gJHkY8
5OCPiISYug==
`protect end_protected

