

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Qn7IteVsnZ/mdHCLR8tB/KgmTn8ijcYuBtDLGh2oUVKuF3qoFWhv7eC1IOCXLirwb60qousghfg7
0xqsSbRyrA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VgzxfdCZunpPyUwqbYGeC3ulpMsK7w2LNEgFOrFKGlFGTp9v30dyUA7MsiKFgCrzzKT+VrIPwMvw
QxU3GQIE0b38WJ5xx5bDenrFuj9fMfRnJLJFcG2V0iBV/hYdVoEecQkZyqCPVfkUdjfKW2nQQ9vE
YSgHM9qDx8fLqyQ6zAA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1ig4g7vOmzvtScDRtVb+tZEnSyg+feSk/Z8usEB/u9AljT40pDkFhR2JxLDYn3XXgfKo9dhNCFm0
whMJYjKNylxxgSFkNtQwR2XIg0BWg/XJdnzmvhE+MtmxAUvbHjuEhgVFiobIjRufLvFlBirtf174
Rb6IlMY8DFzGP8TNtNYlVuQtzXS4NvjPSDwmxdLLBUryIvh8XgTaS4XKcRx4c9SU8usSs2eZmKp1
PQzsFR6KYhbJsoU+KNdgC0qr7WxKSf9E11HFfNp3O241b9T36xgfVJMNzGcu/ZHXpRemcPttjJFK
GMln0o/DwR0gidlS+JLK6pgrPDgP5/6nmLlP6Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yE7rDdP/qWpLchJqOpJirpc1zOl8T978Yfk6G9kBcFGYD0r+ZC5agvccz99iMwduJEgIxwFmjnzG
7g7dI8mK6Rjj6eLbQ31Mhsmq+p5Y7KQTNM1pfCzFCw+oJzuBbgsBggo35NClB7Hfb8DM7OriNRWJ
U8K86UkzA2Prba4TIBs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BN9F+vWJYtgfrzbWbiAE08ecWOdWyzeeA+i0U6sGshkhExwtl0R/3hfy5ttqQZECat07SJZlP3jh
V4CCuSQw513kvIfiNR1n8KZK1ODiyg59gOwmz19wCVgWfDfnfDXmgYxf+0derYmc4F2n9+pXRhDQ
enznNCCvV1TM+SbAXbMWWC77ZJDkWposT7aeuix0KzNLkoMsiFOvzPJVJxWsxkGPtD/xLXraVjuo
/R9zbJjLpYz0T/O/R4G6FwuMiIZFlEBmhA8YI04Xnb8Of0h/udsHa/BIz80Zs9KgMYw1jOPT6P6u
7aYcNrAi7eu92a51ZSDtMllbDqQBzVGgrUZg9A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15376)
`protect data_block
N4sRPZrUknmQ26EKj7eGpBtVgblVuIT+Xc2o4UWvaO18T0chUcez8oZOEaetJPfQArioBg2cG8k+
7Oq4SxnT+H9cspqBlpZf7YvUxhlivGwBPIy9CI9jk3GKyFBikm5KiZHyi6AdIaheqhWZhXnSlWaq
UXppTURLCKo309Pon7DG6k/woI68OBs1iG1cmzv7vKWnMNeAAJ3jWGIN9qFoCSNPAh121IAGlq1g
ZWwwpM0QnWYR/c6bxI/VLqP6bLwIbuskchXSqUz3TRq1+QHDRW5hbEOOae2Yph+4eGox+5yxy7S0
88i7sjQXp+0YNfwCXVI9e4vrGdhlQywEHtXEyDXd6q3y4r1HJ6MvziHQ/3brlxwQVy6Lh9Pj2R2W
FEyfPmqLP4U1qP5RkELGn0pghQbRcH98sp3j/T5wWFOnGAvw+9SfPW/TtrzL4SPCx0HLm8aXWZcT
v45G6zfvbpBMJgfxhSFabxU35YAqh0ccPSx5Uqk4Np1M4JVSJHA/gCh/AiL+6/ZNUlLxVvo9mHAq
BYZ9nkRr2VOvIluQIk34TQEN4Ed5EALq5c1e5peTRMC9XwdnqiZsA79xbuA2PduOsHyB2mI5JXmO
rfqLQIA9iebOjpIK32pfx7YhKN8+EShJe9fPgbnK6dfgL2wprDu4NXQHKvzr7xrG7IrLcklLdcgc
T133SmhXzA7vx/HOJCo1cGIzwkvLgBf4NSAhSIXZcerUA7fxY9QReLclORuaAO84Y6lAdizjRRpI
tWoDqr9Ik9zancufZAGD9XDIkb46vRW3RvUsB08ArKyHlcsZblucmW5OXR0Q/x8VdkzRkQm4P1uF
7iDVo8/50PnaHABOZDsSD37vUl4dnJKA5BmjXkf1yFmRESImGfB5FIollWszdBl26udyOWwZX0zS
xTUwbrDDQm3qSJf8AItx9mRJbow/XkabZ5SuqnW3trqM0LHUaoBQZK/xje7JE5Y/az9FZ0OQEN7i
IxpQh0U9DAxKFz6SuTG1qJHWWx/PQwicIZ8FyoXJy5EOCSjTt6RCy7KS+gn2hkSy+6CgHlQJ6IAY
1dXejoOV85OpV1DJUTsk2CDRQiLG3TgknnAIoV+15TrmW9dAovLRWHs+H3jGx6886HqH1NwpX9h+
mFfnAWz9rXXrzhaj4oa+cOR0vRftC4+sSRXO6ntRWoH4ZTb1uLdfH2VTWJyzHiyc7tvr16hXAtgA
cE6vI0jCfOeDiZd6+FHD/2X+FiI8h5S6KnhfduvfKo4P8EP89mkvyn627RNTkrN2rcLCAeX+9+q0
HK5+iSFUFhyOHDOWM1scyq0G6AG2AMBDqvAaIFV1igD7exSb6bHEBLWp+bZBUPPzxZkMsmx8dfMY
S3E9k+uv7uyZ54P61PjyG52BO7CzthHIfHWxYVJJ7ShzL/OfWVpJAZhs0PN2NS6ujvciVbJkaWko
U2ZaYF5eBJ6uEKyeJAdKhe+scKoo9bAwsnL+eGWHPfyH/9P3BVqmLaXTP379towsyZ0zzS+h7guw
8dfNdE6GEeZ6HRwssSzPqNflGNpBJIAozetRP7F1TzsiX6MII6wfHl7SilLGcjGbiewp3rR0mdhy
ljqoHKB21Z85gN0aLMKvkUpjn7dwtWRMV9n2oEN4LgQZHryQqQaCnTiX2nzs5CKOS+Co2XSEAgKW
FpGTagZsstNBLK8/5AeH0R5uT+K/93Rw11XTOAHPrnrJony3i4f9JIEt3jMVGN5vlHYV+vI86vDG
qNBg195LWDM3ZV7OEzHQ9YSTnafgHSFubUEJbdA/StkV1FcPpSlfTTGJK8nouVV/Omm0Hh56fTPk
ArdXvHHWX1CVq0ZfIDyKgT8owHoWGteMEOL5WYCzWfMifAOX9IkFi7ZGARhVK5+HMjzxceVUNT8d
rjxTi1hVK7qSXS4PcJ9cvbgiLmBIJQnd+BzUSaCtmy4oFSoMmEafG0ltm6jAIGW09qq9ePISB8hT
vTPLDHtoxDI1vlR3rbvCig46q2deNQbZalmLKULioBut9FP/6cBc5oh65bRAtd6IaNmYwV08YsCD
rfksaTNKr+d7H0aRr/zQXInxOiIgqJneD1aUHOFQNtR1t8ovSAdfZei0eGGnOiXC3kNwRIoak/TO
Ggc0I7hnjrZObLAHDNuWmQTVvwmItVE0Y+xtx5yGDvhPrB99jrIHDF7BZtFhJBMe7epo2YgdTVmR
G2OdH/bdMdh/J2ShNjjZqQiV+lAEiFilPRYDXi9a66qvG3Khuaqn+q+jkXUW5fE0x+p9GUWRjMkO
fzXXhctN1CHDuaO6l0j97QlXqfOgPegsFAP3JOarU/s37S/VRZk3IC3tAR67M1AmEnXC4Bp/LfCP
QvTPKoqaxaOzaCKQk82U7JN8qP+pexGKNvmZy82wkCF3O/+TGTgNO9qJikGA1Iac4/toupeVFMwn
BBzAa/c9UR8pTmS22YYySgzF8sQcho1l8qaRu2Hnh0BUQ26EOsmL0jCJkOAbeUodV5hARvE76Vum
Gwx2JioGw6xVOn7pZh0PfJxAd+HWBIxExPd8Oi3eiRjQTFa+h9ManmhzHDTNg8iCPoYN99tPHErU
QebueJuMnQFz2v7ViCNuwwQ/BxeVxZTM5LppgESEtFMa3fJDyk4ulGf57kX2dX/zPmw984ylq7zS
Mfvi9VMXjd8IHY43itiidqALZ/1c3I5emtX/O5pfxNhrGDyKbptEugCEpCoLsCW/DFdh8zGYfwMs
xvV99OjlqyZq1jRlRQhWQURzu0l4qE/7OP8khg8iQE1neq4QMHkv7KqbnLYKBUvGvaok+lAUrdBO
BNRBbowRq+IS69x4aTM9zOJxdonaIJS3tkHn6bZL5p5pcXI1nEOlgqH3irFwMbK8A1FAw/BsSdTj
+e+FD2dzmTsigdQeqXjbOHOARFd12Y3bprKWqvUV89E5qMhdyY5HnA2TbLSbpWvKz5InrPNpbUlo
y8RNDx0FGIT9xsWMngoWljIW8CRIb5X5NeIYo5JnHSnLJ5J8+u7BV5fn5bBT8Z0OcihCDtvKIJDe
iMjZLNMKJxUgiX7kZ4rfY/CZoyJDOlv4etMzkSXxp9NO/VTeq8w7f5hEUuhxCiWwgy7qf8eB570R
oHeA+D31ROA3N9SFybZBRkXOEpmQUjWdHwe744e7BtrPBWWyanHdlVZpIWFIu0BMNVhi6jZrhRVW
9smZuEIFbRLYlsnDcaSLk+0R16d5MDdFVmH8RbVP6+aetsLjxlz00ZokMVyuGUTRXT85c5+DjAm0
jX288EVh9cnz+cFzMc7ycJDerQZMvS9EgunCAri53aWmjPhZD0exlRvZyZOAc0DE+uRMKUKQPHHW
k141v4PGeQCP+jit7Nl2q/vLm9b+H56JV4BgWVu7r9cur17v70fLDfFDlVDNRT+ADONyOtNoLkTG
M07m0WprnqkLGeDgWKHnmHJp7yzs5RdO4aPv0PUNqvFIyZw6VJcVqZQ5Vxi13YFLFLVraG/fvswN
jpYY5JzP+RVen7/ZGjZ9ZSK1j7o03s7e3CLTgH3KdvLHD0p2oDK8yqJCYWZKrnzfOkuwaihWEr5J
SY2oG7WMvbEqTVUtcoUtbC4rwQrBHp6mju6wfvwczsBFo+cT2QTqm81mEX+bnYqUt9VKCVu5ODv6
lPcyjdyV5uD1E2Q+ODvKFO4Zups+GGzVTp9ZivM+lTaZdXgB+JWrstqmKv9pggR8D3i99+nm6Roe
+SDMaJsXyXQPwZH/o8ZT/rZ8kDFo3DJ1sF9rREFGkvw3fummrwfdTLr26A1Rh0goBHpDaqbqH/Qo
jAcl55FNnicKIwzTajd++C7YgBNJp7P1RN8bDCz/YfuO5DaVL2Ccv0gqrpdwGT7hQp6cR5eALeNQ
RedsLIutUAsvU7ij3coAQnii7nzcdqbinvbBzzy8d6JwdSqqCG9N8jgPO4+cnWJeHpP6eZn/CFQC
AzOsXZXc6uKb5o0zQaVAEVNzeCttEaHgdi24gQVaEPPYL1/FoTIciTJ+F52jTNU4eUdjjSL3ZcN5
UGKut8HcG8puWl8Tq2v35pB4f2xD0TBWTtMkkQAV5q4TKe5AvmGjgTgABxeb2nsXJX8oix/4/9Df
Mekw9mtcaKQAtPq7iGzKIO/XK1uB/0Gd460U79epWBdEzLzRG5DnM65+J5qhW6BeIdWg1Zu4KhXv
2h5vB5lajVaFvrdA32fyOKLtKczNl6q+WAvrnK5agYOpyUqa0/mi57BYjOZDPqs2w8K0VSOVgaYG
l4fb6uIjF7DffZXG6wGLBYuj0jXgvZFZrx+/FclFPLJlJtW92es37XQCXWLnk5MsxvxhFeDTQ1+H
4fDbIFTouDqOdvXiDnTXCyl0aYSSQIlQ/SF2ZV5tAy/XI5D84Saq+NcoHZQDbfApiCV6DhNrmP0E
/e8BUcc/t3vXVsn0+5xnO41p4Y8ARP/4zuIttNsddAvc8x0FNEtEXPPGIoB7Qx68YdN5vctf6S/Y
94ZHwg37qljN3C8RgyLLx1rKY+zYPKv9itpcEwdZRgwm0rvM+d61sDnfxvez7uQgCthfX4zknkDU
0/ryF2Y5oIK336J2DLeESUbQscInGSXPYWoNslxfiqFpzGJpqUW9zxAIO09v9f+Uqyy/1J618iu9
gJ1Ug+zsb0VJghjTZnYX1ctqrsGBMNulaaoqMOywREDT1G5Qb1wzEYqhtdx/GkSHWZP2lnEXxioP
KcRyfo7Yv15Q1ymK5zLoz9AQZBLdOE0yF9VkHpxZjDnjvGonIOw14lphndpQIQAdC1h0/XJaTPua
g3aqbCigtPjp8Iz8qJs1jfM45JluLaiHJ+GrDh6fBLphTP2blMWyl1baODYbDpUC55zf48k65+nZ
EeA8x3c+Rs8XeMSeMm7XMFdMJKp2D8IWzEH6mnNeCQq9PE11re14lPPEyG44XdQc4dbHW+pFmgPt
KdKkAvor+jKScQfpIhBUOaZQ8QnCKskgcU1HUePfzs8elDlSrotb88mqjaacF2juKmw6amvqy92n
5t7iFkUKowWLggJYfTvA44sPhGlW6onEfVXb13k83vyLPVjkWQ9+FLNW3se2iOWPB7kSvfmVmvco
AcO0v/RL2LxlrYf8ogSM3qA9+18quVitXZ+FFlLrS5CMnjhHAtM751V6pX4n2D1nrg36yzEfc6A8
j0FxQ1Abj5O7TnhEh7wfb7E8xleDjPW+/x5VavEC6Okpi3ifbWlGDzdi2JY5kDUIlfVrakARa/rd
kSfwQAkRixN1vpLgVOjESeikTFQAXCbia3XOLOUzjPrumb7w7ZTzixc8WxzmlfGXZqcWjjkP37Cq
N/uM8HaxeNscAvO3d0V5hwIfTqD2Kh5CiTVnb6ESA5FuVIpagwSonhg74edoDC08RoKEpNwhEGaF
8w8RTIFL2nrrqp2xZhMKFc0U7XSNpFkP2guPV0a5ijs3/5TEkfqvVV7LSBkEm5A2e4UrAeniAT6S
nrNSack1gfWly1bIOQOy5IMvIlWUvxWJYB67zKzMcUkCbThUfziXb3uldMTkuITEkGzfLHguQeo7
6BsQzK8wjxkna+qwfdzkVZIHZ9cAm7IJ5dvp+/+fKxDUkQW+vY6wTloTMUHfPX7WMKVo685x6lIa
HnDBW3R7bAIIzfHH2gB1AiYKx38ntJtqCUpscfnQCX4fKfl2q5XskWg3zJBQMnI6li0KxmAJN7TV
Cy69VTjJcjKi55eTD8OAkG7qVbdFyXSqhp8dhok+thzhiBenomlC9+ErlF0b+Vxn2d25jhkPz5vR
MdXzsdC254J8Sg/pLpImkx7jof906o7qEbmH8pg64RFqJ9C6bSCE/5x33lZp2GTsVKrR0A0+UTU9
322hhCjRaA437gyKawP5FkitkG/N8p/k4cj3phfeLhHlVHPBIw/gb4BH+XJ643GLsHtNMZV4HRHc
8jik3O/d3lo1xdctPl6srDOuYtDw1jAPrDt9vefsqEjo0BHvlhk7OQnn7yocSorN44KZsvyZPP8A
iDzavemXkEowlYzZO/yOcuzqTXSi9hACF4iE159Ud56v7DedF7jH5IKhVkX8JJcUtnRcQE+WCACe
URSDtvsMYRYnLUYaAIgS2s55FeivaEMeNVLGeV1cd/+/MId2JRFVY2FYJMrXtvDAew07EMtNszLW
+1S8jt99PW5B3zkZyu5vPdv9owL5xkVb+c6UvNMRbZXfWJgIkJLiBnHI6xHEG52uscRyfd/0hx/k
W5e9Qr8c/Yli66YBDPJZPDQHd47ByFTCiFZzj22LNXs8TQamb0zj2CvDIC8AHrQXaG7ovN2fk3Wf
DfYf7vuCGPq2ybnNffFBKKIAfzMahhisfk8H6u0GHksVPof0/k8VNxk7m7fn4DdNj92HDo3oNV10
UYLnNqcIOrDbMF+7Y9vji3XA1nLxaH42MonD2zlBEbS0BMk/0V8qzG5eu8fENqgfvOFhihKQ7xaF
K6HZmr8KJiEjWzbYSrT+NNnSG1SpVqVJqjiKguuoJBTRNBN43geFYYsWPoVXBRs2ZBZwOMHhWuN5
vUOpIJkmUE+hwIHgc6vq8pZ5OzdkkbGcDyUnETW6lqqLx4GASmaQJGTTtRzILOe6lAAfCxMj09Bl
k1lqcI/zqf4tKSNS2kjUMXGWA1sCm2Kru8vAIqRQpuSSxWKnGb0eASAhS+sQKJHtU2+SMuDhNXPe
iiHCuokkfSTN0qees/pDnQf4poJqO7Np7Odd2BOExo1VMxo3ZFm2MwZiOpIAoeVzt6SOQYzCgB6c
RFNAMGfXtHh7DJ9cLFODywyQiMpsXXSB17KCyg59fdCINDp3FRPUHN+rJY5hYUXqycwLPJYRYoGL
hlRfqloYsNUk50ENeiFoWn2XdkfW9rhc9HvDZuPMTzErR7alV1T8RXdwVHNgbhpafQis3Acnn6he
bBCbCHhWKOYF0v3HfQn+46JAVVcTOt8ccy0QH+1Ow9a3i50/bqlUj10j0mxEYPFlYjsJMfua2a34
0Y4lP8V0g6G1HG1IdsVzSAI55K6eOYwUZZhTkV9rewP9+3lAUtok2pzLvkdJdSDM9Qs3JfX9fanP
IpymvQf4eXPPB48ylidoIJ/dpeqTSQZblEN9UgAi55TTBhbNf13liQrTjJKDMvHe1jC8h0/klNdm
D1HyTaoeKNBzrqHtUKi0bmgOVcw8ESMvAmPNNoIrxTeZ5zboHEZ6HO/2NYPB9LAk94mzlG1jVUsl
/cBEAfEvZ5GFNZqY5buI0arNGE90pYLmqQYcp/NxBA3dqmC08UN5VTGHg9j4zOtqFpUfOMKHyLDd
buaJ/oFcZW6uJC6hGH72yNNTjB75wPPqchpV3rtWiHkHCBOEoGSQuW9cGFl6J9YJ9tqWL0AF1Bl7
7PzlbeNdZRPt2fYrX86MRax99iDVD2CqpD3V6TvM+7YGeBnAlqoSnT9N0bFm1OHjWv1LDCx6w2G3
t08aCznxMtdWaBib9QMvejL6bobWpn8n8HE4Aro7Haz6ETE9K6eQNbkngbxzbR2OOahh570G7CIS
PziBGUzroOKG6f0/u0/WVoSgExpCvR3RYX7zZGIfCGsESTAk5NhtoaS+2ij0tBHvB50tscCo6sOp
o/+6gUzvPf2FGMK/oP/2c3WkWEOkJpGShXgNwZL/6DxjJP9U6wqimOezvm9+WV3Av/i8rgdAz/Nk
6s1oYuwpabt/iqg7BZaEUxYTS9J7ey2cTXDJUz1wAnZQlEv0zqYU3127OBagtHu01BOebg3lXAGd
67ehH3l8Mc5Q4emuWb8NkHQfDUqav7P2+dskhHNA0VTvJfVWCm73gJmr1IXbKXdx25k2oN4mXggg
7WFjQt+pHMFa33LKkhznDlmh4WBJtGyXN4H41DcUfhNhS7Qs2r2ECI/aN6dqAsY8wvPZj1w8X0xJ
4tpbaHrOIWfzFD4V8HqjVu8/yR7PTN1rsgsRldYAHKTVxz8xWGgixBWkW3tFAouKqhbZRVvGTFB7
GBxHzwoXSBOGy02AWUnBevvpShqjpJjlBN+MSIKi+JjL7cCsT5RePztfpbg2UljswU/RpKql6dSC
Uh2L2DFlpd9V1B0HJVFEftoprVWfAiyUhUDlshhWvgLUSlMXB2b9gbvnl1MyLq40OIMfp2xAYqgs
XNDE55cMCda4EJBEKNfCmgThUnOl+jME6WBw13u6R6YtkGx/Gdw5SY5Pu+l2chE4/Q2zwT/i0gun
tEVmWGCj1RA4oo8hvchzBMfkOe7fCqPxMGX6+rsmhH2jmlKRCJTIAjAGKFZX0rrT6nLIEWWqLlv2
T7pP4iYb0Z26hdeuT7lgwfBoBXBdz0iF1MN5UtqHZEjtwAq9Sl0mDHOErtHl4+nRFCr9ySof0sW6
x5ndGuipto4qrtKjSQdnmeN/2Joncd3dd7StWOjWlOukVUZ55rp1GzOd/3W1BBtBt3y4fLJQzFdN
AWXcJM8HGdCKa9qmYMrHh0rMusDtMFyYEu8ByQQtkuZkKQ7NBDeJ+9h2I9p52op2dI79vyGtSb8A
lFjFXaBLltzK8OR+/wsZY4567tPQAGfqeB5tXA4KS+Kjd/uDAqyxIL+IZRVphL+A2ShZ5KAALyZI
6Q3o23+nrPTdTFCRFDQvytstXfwg4JXRaqN5WPj7BSd1461fmm1wWMLu8d63LHDHlzDSFEiuSg0m
cdo8MrfQzwEr0ZHSPFScNZQhgOdTtuqvBBUfTfzMwQLge2dcSBqTtI0UrYfmUII/b8WXd9PqSJ2F
Yti9ixaOBdlyi1NSQ8qZ1tXKgWD270j8Mlij0Y8X8TlilHqRnH0hCUIg+Rqp840q+ILz9keOX9XU
fC8w76mKsvZkplM7Y0H+MYFjG0VN8XtnCJzxf0C0Evxlozs1gt37be9rQ89ZTkGdxcj1gnm7yAIE
lwqvvmTQ89dkOOIiJL5hEjHjMN6nvdsDatRLxAe+kioYNJTcqGcGNQXX/CsRvmUWTHhcZxgpHycZ
bVVv90jVvuSW18xQoqRwvxuCQtCxOVI2j5ZFF4yf5YAh+Mk0wq0Q0VxTKrWkG+WMX90E7u8xwiWq
VjAksvxvv06Y9Vfp1H3pHqUSVblU6wnK20c5vGg4Q54jJ9M5bb4oRjLDamFBl+oZOx1b8QR2Qx1E
Xy9jOhMcWtJ0PTlh1KWmM+qUFcu/8nPrHmMKKpM1mwZCxDdPLxHVdQgSpUoWKNuV4sGkCKhNFeWn
NU99UoFgADAo55mELIQiKmyM0R+i4UQWlG0WLuekJad2V9WHbFAZaWTXU/AKtHdsb8zcpO40revk
0x3fpa6gNT+Ys+R/QkKNoprfIh9j355sXuOekjOGK6u4txVWNyWNTIUnP913FEu3rtOVU44hGwMw
F4SaI58sVZId///8soyR1Sq51lOqHBFC5jx1L5vYMPltnGC9DaLibpwM1xxk4AWreSLwHDo2ToLG
rCoLmklhjiSxUdxab6nxjGKI1uiH79UX/ApRDgt3+ufkxQqCd7ObYb2UnBUGXTgkqkfkJDK1tGnZ
CN+YpqNPFyEEtTz27I5vExTqrQQnXgbfWZBWDx1Je50J7BWsiIIZZ9PfYPZC77Y/6ufSbBB1/zb7
ec9EXFZk+V6RbV4cFy3XCfcwbr9S/qWl/C/E1rKDPd3gvoPNzHcJN/GOVBA749duRvrqAbgG3hRU
nxLkIP/caj0EIG5als6pIptlvE3cN0lIzZ73CnB3dr+NiGBaVFjYyMX08S+Rs/fxew0rjdWlem4+
m+w4eZtSvf1bGoNyGnb2Ib2cgZgKldZQYaemECj4yRdYofrT3dJ+I6PDdsAPCRXNM49qojPzmjUk
UdcC7E4nsvTouf//mzw1xp83ppq2Xt2+/5eLQkVJEa6Z/mUkR85ITLzh/jDKxQjBwXMiS5iFxfoT
tPHXMaxI2KIh8pBrUCqpDvxHcK16G1Gys5FmFqrlG0WChPlegTczgRwkPSKwuRzjPHgv+/5ZIZ0H
1A+jTHNMfOYvma3djF68T15ZIbHxN6wdtiVHYXzH079q4MfUqfiI1WTZNU7bPoY2OWRWp0W2bhum
Aop6WT6eJKKpxTsSObB6HmZ8CJdau8q8NlNQeOHbdWYDPbJ870KuyQZ4RajfVBfVzsnn+Q+3l3hU
H2iNiOLkTag1XzsNV+9lIyOTuAV1n87SyNmCqfPYxtTlm/jlAjKMlhVP+riK4/eYUSHCDiPdyoGx
HpcSXSRfeNbPt2DB/6efQYDWzttTYmn0bGFgM7jpzrDTkxycOlC8nCA9ihhEYY5A32ZH3b+uUm2+
Ue6f8qHiFwlYHyy98bzJeicFw+M5qBmac3tkiB42P0rp5ibom/4WuY6jKtCCmRYRp0Lr/ctiZ7NI
28q3LIwVnwIOOw3/KUz96cIrq5/lQrcCM0B8iG/4/wqeIb8FR/Oxr5f2FFhSoTn1kjNIAyhoWmq9
hTAh6jzgXco4aZ6CD3HtFTSSMG/PpHuA92oEXHHVU8ofSwaNawbtI0XmckKPDLquNUt+lcNpyfyz
rCwZ31m7HQsSOlWiEojSJWCBiPKgey6eRX9KxlDRW1y2k+g8ul3TLM93RypN3DOmf/Z/9dbQHfgU
pb+kfYWs17FB5zGh1eAb227jeYXCLdHK0ddqrPLMbSB6kuHgg7TSlWESX2PW/QMCbQVpnjBV2OYg
oCr+mrsH3+AIzlN6vRgC16w3wzvGS0U/WKgTvDlqC50p2LMdAO28HLHhHILgUZgtEQ+cha6fM3Jj
0r+C0Xdrxic8gth2MhFP2dC7HpWizZFNb/CDH3h8fGB6eW/7x7b9+1IrKw/MJi19qFkOotdpoXvK
KIlXX5JwKEaq+deY3qWq0wBDWdUSPBdiCOz0D+7euntI24/64DIiUNIo9AGQuJfUHYJtZRfDBa63
3NO3Y+9YhFcx4K0ly2o8HT48EE2q4f5jpglDRzyMqvHB3QMMQFtyfZRga2AdoGACLFX68ThEwS+P
/nIrtn15rIs44dWYoTqPPTAO4AW34RjgJedIslpND7ihho+lSzg6O023AHSBhOhwcJa1jx/xuCiQ
7dF48joAtNx4IxYyhmPQxE7Up5++4fQBRY237YtJCvioPBQB4LiCq6+8Hc8THk397EfBgpA7mkce
7d02Wk9ZtrkAhYURdrYyKhANcHGASaKGCfMtrwb+y8eDL+veMNWmreetcDuLPlKiWLHZBDYm6Izx
j2Q9cgBgQX1JESw5lAq8vClk2VN1EdEwiK9N04Z1wqd0K71pKfTRjoF+uP+YE9YjE3ADakxfKmZM
C7mTV0ccxW3o4WS7P/Ufsc28VE5uJacQU21EfF6Z9RsTVTOI54GihJMOOoHOacTcbYZZuAsVeV07
AISBsVJnZM6iYPhmuGD7YsofkcebFeg3S8zVuARuq2tHsmrbyFiB6UiH+Q8NIHha8a2NlwUX6t7E
5KBr/h9iqm9h3fOFo0iC8g/ukxCzVN3S5QN7JSGQeKSnxzlU57qj0P1ulLWEzq4X91tezhNtjkHx
0U6LzxnHTuK75wZ0n24PX9iQhoaaT47c4F10psQ6jzaAkLt4Tgp6v6mUBIV6BYFwb9/gVQgRas29
hK/htVYlJNK/npprLn/R2kLdGigFLcrAlWfym1XxhwdvifX6AdvxkJBkqWJwZCYF60yhcEuLhIzg
QdJ/k0pEGpliYeIRGJ63PaNe9Ak55ug0bNTMeIpl0+NRS5oS4mZjjATgRaQCLjtCa0DJj8QZepq/
uvCZO7dSKespq7GcpIySbzTCdnAeTlbti59Q9ox/TrhBsD9Fftz02LNN8DHPYip8hphVnt8DwGRF
IcpYCOoZU93fuXKo3zWcYTK4XVtwG9Ihau2tYGNaY0d1ztULf4SmRcUXVqOm8/p7qm5bGa6i6RDK
gImkT7xBDj9L+YqNALCOggZOsJmHkbVJlKAMGl7uShXIuN/b+chbjPrRJ5Wk54K2JuAq29G90RNO
Rsi/ctOF+T4YV41hRInjtgMU1S7ZK/qMk0snFAZNdxzTVnUpLuCUxrDAboI14+bhjcg8A+zPaweX
bPz0tJBn/WKwQlytw71u2+D9PWlZTKXIc4PJOK/+F9g3UX6IQ2zejbTOrSCDIxProHgjWfXzDq8q
cFU2+eS9xN7lJFjs7pI7nIhyvjaY6tDiOOpKs1IBN7kFmd2orLtphh4aEnHkFLtmNe1P6MgJZqs2
lUIhOgNR8HZmQWep+RsnwlCITHSWpkJRsGs/DWgdmnuxQ18mxRaKMvbbVtcLbGNwB1PdXFgSagna
HwpIyMf9PYhYr5dNdwV0AYjGS5l3OsnDlzF0OIOQ3R43NhW8tmHiKFYMLQpdWhCNM+jCYVNo6yBv
w8DibtCuzN0j3J2/pfsoM6PcwsLkTCR1pkrE2vLO7sbgtFsNo/2LaqkS0WeyrVu8+aoO+wXW/TzR
9jcMDORo1fJ+8GIOAm350paRG+6RPROb/d64nZt9Xb9IosgnbXEBGGLdJ0lDvnnNbXmXOWy+A5lP
n2UGkrDj+fJadIsxti1KfABEYIQczt+8FCgPSbZbAzJYwpXKwnBbibd02bM0SP9s7VlsZ4uddx7z
BJYnnIG1RQ5T8nYGLfU/w4yZxtwOcwFrr4ZqC2XWqk277018pTw+wFMIkX3YL4p5A86zCPuE4YM5
9G9VnzR2E+7QseEr587e2/7QLX5IVsBciWVtg4ew7Hv46Ro6UNXuK6JLoXw70C6Pb//j0KfGKj1b
C4jAs289XZsscDYmFPtUhj9Ns+oM2NWJVFC6rpB31p6jXqWo8A2AC0peXO+ImoxDRsoPrUi06iAe
frJ91BpMsBaN3JYuCF3LMI3nHiUnWdQ4ZGGgVh9jiFrIUWhkiIVTy1zYyrDoFezDqx+E9RSh7/8W
1Q1Xj+xmuJMA0QJAEodaancR0fKRSx+43GMDd5aMvefh4BpAA68GNRKlAKCYKcufA/UQEPYnzk9h
3gSWkCCfQl0CC4XQ2672OsP6uISu1m/7PiUMwnLradtOeYr5C8k/SVI0+BqKapBgZBankFajbZnQ
nGBUvhcmUUuZ/j829ieRRF+gv8KR5uXj3+kCy81ZQrKEUutYZP3UDyiVj33ypUsEkDHPzg1ghYsS
Fm2FrwWrfQhE+XuSLC5+PwjGleEu4cxvOsFb39BLkg1iXjtRF2T5xNFXApJ5rtEib769qYDcE7WS
W//gRgYae3M/wiI6Ru797Z6s8kGKmcaVS8mcce625mai+lIhgIoDZ3JHS18zuu9IfikDARnKOUo3
cilnTX8m5dJXm/eCRzbUVSFyWsiydGOljH/gVYBtZVvnC0ROaSE/ExUASp4rq/3SZfRbT5WxQuQN
N/6ZID0p/wYwRf/R3d1ceLgnfxxYu6mVwn0T3Erxdjc9FTlFgmt7+LA9fhYYB0GvdUzfSo2usvTa
YsWc3ivU5AQ1GE/7IFRLY0qIXeb8UPEUD1NytJMMIJvM96iEbEXOL2u850XJ3NNdKa6hjK7bjRtH
OELE7bstQOAlCroPnscTIeaUSqSgyp3hC4zsBcHW1cZqwivn5k6h/jKFzekj9LEJT3nO7MgRvHXP
fjE5HSy2a0DlQeadXhoHExVvaUUB5PkuY/J9q0wZSVzxPz+piKHeWINM5ymPt38Js2a/SzssvuXl
emgYy7q52X0JLovFE8Nbnc06JTuHEVMdhwxQeFMmprKOE+3IF5h2ly/JSJTvFtn2zxmlsZoy7Mp+
nCDN57b7A2FTwOpy63D8xrLhvpjGpVHzPQw1TJnnoGxYcWaOm6BLEQnHz0UestPGy6dYDPMU+S67
u8qbfDubmo+FoAJcSMn4Z5BiprxRpPUcEOkR8J/L22+bvrbJyL4JjzASQK4wDpU9uk/vFAbdel6a
44knJQmfLgii90HL53EEWxzTtKFOwnUxcEnsfAgX5CsmT3vI+w4HDZYQ1hMv4mEAKoFzBmyA7/rr
SRJaWnw920TPdmrTiwivWzMCrfa/Md5VIeRAQ+6Ngvz7dpQn72UKfQFgTi+jiSo9kVflAjbWwNXa
VMRdzxjIiXgbeZxf+4niZvWYg3miOPCc6dgsnvM92to2UOlZArfGqc82zjAvv6LcEj5x1iG1SIVq
uRZPI/yK7ASqCIof9qapikf9XpOWWv4Hxm+tcn/gJlGyy7uMj2cDjfk4GYj7NsiUR3Kf1H5Y6o/z
3zQB1JOXTDqSMEHP7j8kACV7+OHnsVWAtvUtGt6s3QX9G8UyszEFbDjeJYs3JS9WlK5JBSokuL82
AYKzO3kyZ32n6lL2sArFg4HdUVONypOMa4jml2YcbnLfdBuDMbWmxMEPW/Du4s/gAQGToT7JC+vl
mqtCZPVwNrpOfyNSRPIy4yy5bVVUrB5FfwN90MJLSkNHJ4Whs1jmBZonQIW3u0rTaApY1+KwZJ+B
hSIPcxubInZo1yTZrsuVcX7wsq8WA7pSuri6Ypz1nIwFiUtblsxaHGeXOl7dJzOOn5OR71JZm5Np
U2kG6q4oyq1eWzSM207G6P+ZONMUJccImOMOZarUvKBdL1ryppuWGF9zsBzuEZRyd6B7L9UTkqA/
w7ryRDfzpGi95lyQS34HBV/PRRPvXgvnSKxPqU+MX4mtB88zraj7T0e8ak47PYvRFR1GlpXBGVin
KrbiRefTG9uFxleEmCfyRDYWlk+C+iJBuVyW/h6aco7oP9urLDi93zR39m95VKF/NxgSA1HyrR/z
hZUyBZ9nbzaYQlqRE69ItOiV22se+pK48ccCq1i2ggiN8xKEb1EEBwsT5bvijahQkZ4pwxwdQbbP
UyNR1zluRdiOI31Q/iioDHNqkR7lg4JnErWUkJQQ8hOo5PqbRP+u47+Ihw2r3M7vEP0t3VU/hJEw
gtR0LcnCrIEkLMODN48NRHMw35gb/m93tdxGEtAfY3NWKMH24QYEdmWX+g1YvtMCSUVTPH+7RJKY
IvjhVyrlYNGIpAuOEXQ20V6JfGLC4tcnbHs33Ya/RhvJ1Tx2tj7UH6DqY2tpaHYK2cPvd+0P2273
mG1AUcVSTpYF+AErF48gg+ZVmg3MX2n/A7NQplN57Ee2zDo/ZB2c8do3UftRazFMirXd261pA63/
1bcQjMG4PEzzHrHnAxJbCOt33Cis/vXyNfEysYJQUJ+bLNUqUjOUQRgwnB1xfuYDK4Wa8dwB+uJn
+5AOGkTFhDNcWPz2n1mo+wxu31aeGCONZr++jZXWDV8TjvBLdIETwL/z3n03Qxml4St46ZIDe1Wr
YXVR143eAbvYWIaOzwpKSxKGRj24fHDRShd2GaUwkBCzOaKUWA4GDWS5k00yzZFh4N5m8wdRJCdS
rYEegiIXDvSavpSQkTKBYJJRvlN1I03UgRUyHcX8pEoAZlIgAjqNLJA1GkUYEhjL1KOCT4CVUA+n
a9u5/OyrJyhJw9+MlLGwaZNFopJIkT3ckIewiQA0mOTQpHGAM2olsGu7dVFFzmL8cIldwlJOcg/q
8a7Vv1Cj41uUoztw8DSgyf0GU9mBPNNoLULCbKyxETU3JkRdqQeixC6L+hWyrDlPDPcdjvl/Kkfn
IfOKf9B0zUH0d2otn1laQ2uNOjoXrDk31bOLwM/RP2TQSzkCrJAUsf1vfqvccok7W/SUGQAPf13p
Cv8ecyHi3jADXRCASoMzFuX7OBp5J9dMG+SvX7B5Kw9GNGFtGz0bxHsNbBs6FC2P4j3f4z/nueta
WHkuWiSlUHHqf0RUVtyGja5O5fwx7S240qaR7UGvhz4+XROmcDzOCJIfbgr4tL2uiyB9/R3kBONR
a6JqpvILv26LSl7wuemTRgl5p2IYxQ66HBSHNJo1nf7rKcGlrAclN228zfMX8So3XAVyJUoBUka3
ldYd/8lpGu6nAHw4793zDLHWL3gvxUGDLtacGMbKRGdJUVSC+aWPNwNz9CotUUldD1E8sK9Z5FeU
HyZV6KtXGIAtbnVnzpDbmja6UTGCMU2ccBtgDrkGQBW4PE6V7C0v1iWNmE9+MWXqb9iwOk97HJqZ
BafX98hmNoCcV7a6TyzNgphs5GlisLto25W2Eo+SYUOJ3sF5Hk/EN/y/QxFJ/CCDDteVn5PB9+UF
/6OHa4N5mbmrYj8xev6cfSzBRBNSmNTEdpJDTFDp9NvdfBZmLSXrJ0nas2GBwSx6RRAmpRxpxjXJ
CT0pH8G0WCI7fgu9N2UH04qJ/+A8kUwJNjlxdZbpqd7jf9lLr6ltcOfVHjmanIwJzUgmNEF6hKff
mwDZUYyjgoDcmakrV4//XeDoBlFVuw9h4qIPFrrnQ4wriOKrKlgQ4tsGeJA+s9ivkBSR7+NVRTrC
nv729QUrEyxylSbsCdC68PIBmHwzYTzLad4K6flJJTX9yc+yjxfrcKkyuMam4jmbiWlRoOOQ9Dzt
HUs9FddAJeEA/2ECIaSPFMnYSr/nnJ7jo6HlTIfHFuvcOquKTFbt/CoaQS6l/Q6DvOZh/Al8SkpZ
TBmppRTlSOcm0qxjexCz6sQGTC0ogihEqZtPCKc7ZOPR/GTFbz6bu3ndIdnWCTOsasdloyjdmPs1
fHydzoIgmSvTVHz6jT6Be9lKZsyMbxRCCF90Qyrn3MWWSHObfDoZM47PMrDhDfaKlQfCbVRw4a/v
V3pqlL3xgzE5KAvAor1pGe3vYzY2aDe7zZDCFr85RLzbg+YcKKYhGqvmFTIA7kiiwHfxsAdCCUzC
hQxPUUBtchKBZTXI7/GxpSV0YoNqgZVtppLfuPCSHbM/lJ5OkOLNRQLgKsRfw6+UekV7psnaiJAA
6MZYwsMhaLZmN/W6JkAm+FWanqVTMYD00quGIBxIBgoyLl6eU9OZSLW8iZ7dOE5cG1dxgOrNfWFG
9Eva/kgX2fY3kIeMBRCp25fkrKKEGcJkwOY/Cqb4x37Eq+HHm7HUVViY1TO8p78VIWtPF04lXZyx
JsZ76KblOboNN3y8hplOJ9B8/PTNP0knXjccOI+IyioCc6RUArD42V/hQo7UEvmz7QcFSadaj6Fu
VZcvy8tTdYMbT/Te0qH5fl3mcbzxgs9IQVNhxKzgJ7VeU+BRnA8u0l4nXN1ma0Hze44g5M7lqTVu
+m2CDQZE5Vmk+QbEFQnMvcE+gnw3ECPWK9yL/UdR9keVevIJ8pjM2OXgcixl9vS6SMkLBU/pROqC
xbZY3x936pALEZnHj4HtCGHA/e+uYnvcHKpOzH0GCeAEx1ucvaYk5CObIZD21ujIFzTOdyoBbbnJ
tCVv1qHdfu3Sdi8pup0K6gk2OQLacX14J9sfg8hmjEPF4oJp+DqpTDg+BB0a1Jcy+owY4gboJgGI
WhrFSqRseUIWueXgNY5LIHPvlfoebw1lj9xZDDlA2qY3XXyKYY25kU7OF1IGeoMj9wkq4QnW0AAu
E72ibhVB68HAHlAXxyhywNw0lswXEP8rVWk0lbEJNYL+43sWKYN0eSIiZ8GQQkNwEv+5KYoQqkZR
jTBXO/LvTul0eFqWLqUquOsJo4hDOoSDYK/xhALruxir+XXhZZPtweX8SuMMCLFM0varE78BvL2M
ebCinpjhd1DETl7g5pmnkKNUlSM6HtGSfQ0x2PkfT1GQyVS7DR9DiXkg77j+hiRX/8h35RO3KxJi
KuuCAb8LQdMUT/FAmcmorvdCWJKtpIx4Ck3jEJeMQmAHSsUeif0JdUzUda3LFjG5DJ3QTACwlwFh
ciNe7vifZJuig3SCQ2spM/jzep+9i6s2xqyl8fR4ChMAKw4ZkKwsF5xnDrojLQE215HSGtmxbhqM
eCwQMk0dfQ+sriLy0LSeUnxLWVCvMKLPG97KIk6oC2cjqt3eQuKfHglMqUuDmSWkd6ojwRfHwPz0
nF6ra1rXO/fRXx0ZAQ/mJ/VQjPPstHABsW3rktGG/17HuMWvIA+Za259Pwa2aPM7C+eeyMvGC2Qe
74lGtWrW9CDIOXaZcgAyf8JSPhuPvmNqKXTBi75M91FKosQ2mlrDtfvPfN3002jw9z8yIwpAvDFr
iuJ65qNCdnzMTjbw0FpZm2I/CJrq8E8R5NP/9aMnCnP5d/T/P4qggixwjh38yXfIW0uq0tb4lB6x
7wESBnf125xqd/7+smLp4Bm6yALFqHlS+CADiuGb7q2Oii9q2jwHHRdrBxgcXlje+PsT6ffruUyg
zP7b7a8w4R8OG2M38Af/Zkk+sYZIJJjLxhirmitmWrOoqb1qD8ACSSQim5tk9sS3XpqqcwuOktwu
qBsMU/cOOzWB18b2M7YGQK5znaf+IHfbPvg2t4k7rU1w1mgaw1kBEyKq7EK7SwD0aZFkhQsJ7ay8
YsqLTz50ErnfV9KMxAEHDamWakCerWt11a5jxoePXY5ZVAnzpP/yFFTAFqxHeWZhEuY40FRw5OHr
LdnFIila1wcx/j7Yyre++1IFXACjHJ0OpQ92cdyU8HOHVOItDiwU9R6JDVgoys3GIrXKjSRsbZH8
EVD1AAHJ5ff49a6xiCiW0LJNlAMFqXOiYibqna4ORSa5NtWxApLi2yVDBZd8FX+4vb8kjUn7UVQH
Rz7HUD4DXzVf3a/rYgQZWlqDdteXXvCkansOWFwYS9Yop/cbIXR2YzmqTZ5hl3ESf0a68sEmwNiD
YKG1EF4Wf9/oO7bnLOg5y4N94rnNSdjej4m8xZZ1n+HofC+RC1epEU51zQrrxp5mcQncePP1VIyV
aUZMmFrMRbAY+yoWdHJvF6CXDe/wIjOZPwrMfiRh57d3sK6El60dhpMYBd3VCLv1NCoeIbHmCWJt
hqNToOHRN6Y7Gl0elMO6Q+t9LuCN21/OAtGYv+2hySx0nBTIYmFIrxWPV+0PbCkvjui50RjOawAY
3r2vtOcsZ2Yd9LO+k41SRu3beGyKCewOtFQjO3AmlYjj39qMcgsvDQ1GJ0l/V6fl2WVu3LXGizGZ
WQiOdenjayx42INj0ZiINRldLhPOgH3muMwLXAGkFWWu5SExF+m2AZI6GJCoF8SCKgHo6VV39knE
mc1h50gpshK2IjrNr434yUqPi4p60iUQkD/z0QAXgYjOYQP77aJYg5hv/Nm8wFn6At5UFMCCvjyG
206xp/LFiPzvhHMVphyYhs1ZrMD77So3If6w4IDal3D74TiQo/C8mJdQzSNqyRel/6wPFTbDx0eF
uoqMwhfyqeHSjLN0i5Sta5G32XVgh2RuMXIQ46/iYFdmjKMoJjbVJvZmSnzIyXpnjC0O45RSwxeE
ldqPfZBNd2wnDoJaqIm6qq8N0zkI5Je6advTEZk4UPTRVPB/HvEA6lv/ZFCZstpZXmkv99Zm5R9d
Hunm+Mxfg51unTyZPoCWE3oqLfE6J/sszuUQ/5PuG0N5dsQcjY4/ec9+AEcylVsCk4panoIfOvla
Hj2cek7dRcmZoDQYfvmH08MHcb4LRQYlr57UNAmtNph6CfgqMiwnKOVGJmTInNi6cstvD/DoQ18f
8kNuSpPgsWKom/pcvlm7hpwjFzi464vKiIgJ5Lgoush2AJD+oYjTDIqYSDa5z9Hri4yLN+V9fiAp
gAIpuiapVmn8wC9FnidUA4Z0Waz5YNomPv6xlOpLabrC0G9+MYxzWLZJy3Lj8BnmDe7TrHCNDDoQ
y0fShF6ZlKITFYQWncli7YGOt8W95+4EHNO3XI9ykE/2Etoor9nheZGU3tfVF/KlMAdpNBXTuauA
31v1LWHaw7u6Eg0AOVj7jcumeWXFH1IaszS5w3IbZnXsUeY7QrHStoI+kkVPUyKNEZAcn+fQLdHP
vcoHNsWOIXm4CgmTULJrBXc+ZWXWQYNigtJ1HoyDvoCYgiHEQHALu5YDFPlFI92TgdB/pIwPNdZ7
MFwoo2W6Ww/81FqXIY8369u8YGKx51oRDGRn3f+4UV/WZtBiWel/u/Mg2tDWKqc49hRKrj5yG/ds
yx1KmzdMlw5/Iqo3YxTN4uxNMCuoLacBrNNSCO5EyE9ecvkkbZ4tychO7b9mrsQ3izyP0h7ih++e
3l+ZIummEX++IFRF4t7JjwAhJ/p6OG/7N9Cj9z4IwoawQloZYxPSYHDZO6l0i0LqPriZO6MilKlH
5eWGQC2CumNPD1QC9Ed4QKHm0K1pUgY7p4OKTIWFCJcxspJ1FFY4I5iyYjv/f+7xBsrdPl9DgV1m
2WflUZIi446OoJwUuNFtQllwL+8MPP/RZT0uQLa3CtEiJpiVPMkJJzBxHkAQRZk3vJinNoOdyi3T
ovXj61mIqpclfm+bDlN9cnQRQOu2rEoOAra5sU8qHlmKtlQ8+cgrRd9RCxqPg5jfZVSqoZCk7GJe
O2H2BCO6NEduiG6AkvrhysvEKfYehptLRKq93bDDpliBJjreAHRjHByvRKtOEmAdx4NKOLkZQMdE
pj3BxD1IpUGDLq3umhBSoM2MjeFLS7/9o6tBH9geqKKXbYNI9XGl1QFjpqVL8YjJqL6edzzwd1ke
sugIdJOHUiO1suP9POz+8nJCCJ0sQnHKnoNdOUG94qwbxqSMJZMxQP3eV29EgAMllKa2NKGcTjio
cuj8QftuaXB1V5u4HvHM/kiF3Lsm8j8SlM9uQMjO1dB12UnVczLYhojJZQ==
`protect end_protected

