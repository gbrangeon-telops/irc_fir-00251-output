

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EHhlU67zSXzve/de+KpY85nXXvMNuZL7tYgf9fn2xs2MMX6KZ+NkxxVYV7RC95SlNzgUt4DfQ4/9
3ul1mLnDjQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UlAZFSxNoqgvPPKliBxVt5c0coSpd2sh9B8mE9L64FOLOsIE10QbDZBGLO1c2gEWIwuQ23M7QvQA
5NLCK/AU93Cer6u3Y5Kw85Zu7Q3cTJ6gtsPScNo+F/wtG37D/TBvZy9QIxLBvCRLOZx77GL+Y61M
X3HQ3kaL5tpBN9LRA7Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BhywTGDm5IJZmP+63CSoL/TDCpGJVG3VkCIbV3f5gGTJ6iLDPwvtFhhY8681GBR+EoOyUSMbP3AZ
DMFHBgscpLa8vafzBYp5kDkIAp6zpVke5p8WT0T374mfT86d/rJV4lUvVArJtTXZ7Qb2BRu+oMwW
4NXsxCdhgqbldJw6uUCqk28aEPgcbivrgwKY8foWfBnTw+EKHyn/oWDvwghTokcxfEnmhIMsR0T3
yD/98FKNKviERlHfn1BhQ/aqkW51Vp/q5U9qrKs/+lZwoRMsy8lRZRggDQnNmQrFO+0t1Oq/DlpL
Pzgpskdyam5KjVkaaUDiD9LunE1mnunv1fkvkQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M0G+I4o5qs/wY3cBNkJHuC5SdvD7yJrXn6vr03zDaDrjCzuSM2xSWnhAroxnc+rs8YiB5XG+kxRS
nfrpZghhDmt8SYAMsT5eb/ToWHwFcmxPkOwf0TCRf7UHox/rcVr0f6gppZYuBp8i/HMdTy7/9hVi
Jazk/jJ0qiENaXH3lhU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
II8O6ksX/NQP2v4t19inJMyzBruYXofFp7EnZduWuRh3lmwU4/uZj2tsoMzEFI9GURJGr6OGMrIR
LHPoTtEBaHFBnPNcL2m+mOF2hh90g7CmgF4J8nr08oNvCPZORB5fd/Cj4ujbrC4saBHdapCX/nOt
W3mratI2AGAl+T3t7Q0k1PLokEpC1hOrn+eLqLqV9hKaNBlW7DfM0Swj9M60AbHp0kL8sQjj6PfO
zKNcq6Xvq1JnJLzZ115Py+hhtw8g3az1/vAI3s/sf20/ggZ0t1s4m7+wPif6Tf6IZJCySXPmKW47
LjAxEb+MGgXZe5eFDZ4nbVPt5Q03mtQWzOAzTQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6240)
`protect data_block
TOhwkcSATxN61hzSKN1SWQLaCvi4pD4YqQvH4Y0LlXGkKYUNHBnQi3itozmWpIj8YdWn6h6mvpgK
3RwbmbTjBiredzZUY1wP2SGRqxsXzSn1kmIgCjyr7natlcgZkJEG4tFmZLQq0q4Y+yZQhskXU8Jn
uHzDR10PzeWduJ1pbyMpR7cT4bCEkftOADU7sZUJ5CQ5pW4C1rNrm/9fYoOoLbtlfJJNrvACvR6q
uHDZlA1gT8BifSZuhGcPEIkKcXDdLND9tBSbpVX6pAYXUDYK6kPK9Z/4FobVQIIRg5fUV7sTYqn/
k271hv9tDKUOwNw8p4PfZhPKurdrMdRr44Ly7l8tM/8AxJ2RDD0euaIAIPhz4KgWfwejrAX4f23O
4OBVu1TROhXcjdvGLJC3KC7LuzotyaWKe40S7gXwV3ndq8S3LzWPPlQAlVa3BVeowfu+QbQfbgsn
+l6UbmHulKsMw5o0WVVmvVbY+As0x8Q2V8/sSjouTgQKf898CgndYRnoL6tIFU56z6aLKrxERfwm
1FAl9RS4behtNwe+Hc6c5w3gnQ6PTOV0WPK1+N+ggKdbe4s2wK8J9bu56LWHs8Xgb1X80QIbw+1G
Pik0oHZaMzu8U7b+4ORnUleeqMHI2E4qqFP/vLrwtuB2kICIAu122q5hNzd/CFsN3475OQ++lq4l
Aqr1rfn0y2YZg/Den9BJy6wUHh4QZf7E6sgVn1+2oHKEcpiYeR2MCEOWCwA2H6BVeUpIm3z9lHEU
0yVsaAT9FZEtnmYujieBvm8qxhsgG4WO+E8wS2kdXklB6SuCLgyFmdc/nxk/0eIh2xP/a9Ib/JB2
pIqfaDyQMntyIDMSiabOyEQHM9kKA/Vh+4ulyx0veOpI4LWd/rP7ZReRL0X4EhHh5ccTbC5STfGo
gL3OvJtu2vC9ZOIG6Khx8sA6ydHotizj870+5YlhG52V8HwQHD1JLegeEKQT1gP+tf4ouEmQ+uqt
kqckBEazp7DemBw2HSfxHDxhmbr/C8/qo8rLENja9oxzLiX3/wDQ7996jcC+LWQnE2iUyEHsN1Ja
Yqlt8fJC8MLzCpGS2G2kABdk0GSprpYE0mEODp0yAuXNiRubN4liUHvNwBglLUg4uiEBWip1jnF9
HRYe54EQsTHX3y/S8F8rTVYYGvYbQSmMGW+WXvGK1UPEbZh+pOkSb9wvlN92GXx2X3qkZ3Wwgauk
k8/3Qj5uLBLb1ZiMHamNXO+cgyo+ZQv6+6RcHj5D+x0gmMw9QQeUuB7QsNF1SiOuT3JtkJo4Bxou
G1L0z2YwWuc85CeaiiFpksYoBP/uTyJ7BAyW+UCTbjN/9P2ReD0F2LQmtcmR3eKJKCXAPTyU1ObE
ijuctAghK6Qkt5ehBLD/AldCrhqLJoAqdOatkNxfGWr/1cTso9NP1hMR9APqT/OhYh5oEZZbkXmN
flwDYGXcYgBqpaOySmVtyeBMLc7tU8u9QUEcL9BLoep98zFPJilSvgVgaZCT5zc0C3q73ClMNuzl
YY23abviPphveXY4sdlqloCB1ZEnAB9gezy6hvpE6W8pUCSKAKUs2wgPwu/q4ckKLTVbDGXHQe7w
+4KXUT+bVWwmp53DEDCzditLVhzIo0+u/47IxDuX8sEpA0W8re+l4icb4OQjlQt1rlf2W4zsa6th
ZTjeKDYKG4jigVMyU2i8qXd7J7kCKGEaCXXfJipMVMABs7fxUam8BGt4847Ml84yd0nrTzdCui6O
Sq7PANQVnx8SdmBOz2v2+lMtpMAgkVLZN8wOUNe5hHVJsxFm1Xwr3MU+1xS8v4Qqh+zRV7C1Jkkx
rhU3oPtJAXmUlY2NEYmsAeDTm9lIyO5/uedjuZE3Fr0I9PNbRfM+xeLMD7DoNdGR6N86Nc9hM1rH
2ecOkAQBrfk5dBrNL1pupJjJ2F9s9RvPTVW7nu3H7UiHr1giLPMQIXWiTA/C//xESNHaOxA3dzZa
x97l00AhXhkdgWdS7sa+4Uhqao62JqlcKPXxX+SqJ3z6+ev080w7fIgUL4dX3+pCB4mWigMoQz94
jBp6gDQc31a5WskuS4Ew/dMAFBegSrlc/5n0oY2irobJ5TUQsEo4oJ3a41D5TxVHg/dJHHYKqbIp
8RSh5wuHzfPc5OHKeJRmnz92rNti0yDsCOVq0bVzZiu12NUBhz0G2CW2peu6FjJy69W4vEau6Sh6
4Y7GGhZ/EeIQzlxGR0kWstAZPfoTO4JMK7u4fLVCMUycdXypS64z9B538GmaCsQUiEZsRjHEcrdE
1GLB9tp6u4VF83dGIf7V8HZqdeO0PoVDF/hgBbu7T0G7o9Gzriy4klJSVP/z8G6twIvMeo5+Bt8k
ncfzKea1AxBjjrSg42ZL9n2iNXMbynqh6P0bcBv5HUqBYciKsqe63Hu08dxzZjLB6fkQKQ3rjhlY
AmamZWOePhK8IDyvCRrEia/PcOMrD7/PQGzJFxbcG5UIDCeCw55P5oQv99wLh2ednPp84JgY0kEu
CAenFoLMfI+O5xfiaoyrXwC9fIO/cuLTruSqwbVl/chU699rPYSPOuSAqkgjCsQp9M9ebHFxojHu
fvrJmvfGDcQxfmsSH5gjUXzg0YgvnzXaxdTVbFeVPSS7NIorBjctKCt9aIKJzYXISlq4y+DyZMqz
vd/iKWpOHrSkVrs42htvhIn4BLzvFriZLTABvGelhrdJlLBrtN3bzXTR47z5yMm3XebHdzfi4NcA
+AVwTGxLu6Bs5+B3hKSA0gxxuM1JZ39DgMejqOqID3eDctYC5i+sAFp8gz+B87c6Eum/0tTGKzaz
Ocd1lmO2sF2shyvzZJz2f0nYQYMC1IrwEPLcyMLh3lB+d39KtPTAUxy8hd+QoIEdWXBkSHlU1/Cg
t7Q16+FrP06OpDUtYjF/j7UxevY45qrj9RZ3khYTCDOpzgp5CN2c2zcMxV2ytRFrUNvZohjYD/ML
FQkuXPDmv18r+6c8G6QGjkAeyb1+934KssrM4JsKeWRrdLcTIVQEwex3ja9ma4TWTdNCBJ06Aukt
NrPQ+HfaTrvWKfXHH65ihRBNLe+OjToi10aWhdIdL1wUzocdUAYNtTti30c2aQgHASBDnf0Gnq5B
+TJMBFKLgoDFH25VBORIivenNRtT7d2nHssjZ2SCA4AQeiKFsgAP11A9WNM5AMSkBPReASYCKi9b
klgpGxK9zLu54kVPa3L0wje1f8721u27tcTwgWqcpOXdeADQsT66Ecv+zRRB+zelVrYvCWiTFJRz
EHD/KWio+URtuqD4QRAqxm9NVlw/27Sl/W3WTKnAT28K+mF+/c4djzUl6ZXxhEmixeQo08ZJk+M3
RjI86/yA7xH2mZ+JlEcjBmRH4cIc9bkvctLGulPMvXk6fru9r1nycO7KUTTA6Og+NxtHKcka9xou
mixiNmMp9tKG+ITGhuSs1FdNwApT/rIRDyV8uFIgww8Ni2CAzrvk8E0Soa9iwqm5ezdsfGLnM6Gu
Iw+CmyIvA+KE3wy9J9PqI9NDsGsY6Z/EUckp56gAC1c1zr816Xfud6UkAoKBhF029o3Yo9BVJH83
r4QLTtmiTDm3gPZMwtnFod/JvMMtzYQ1aspslA2O+Pi7WFPyXq6Pr/IS4XKhe/HYXY9ePISebpC2
cQeHOwk7FKY3pOsqEPoBp0qPr97CFRR0TlXlASBXrq6wKRCK6cNyLP91ffSrsx///cQj3643Jv0B
UyrmDqTIGqLDhTJVlJYGNuIn9VqXh8K4tuXv+WNedXN63yX/lmIeGzWgCl2vEqJ8hjAbtQvNoXH+
5hPxCiCd5YNSzrC90j8pye7vl/LMhfc3Ig+FekJkljhqJ/EiaJXR/yIx7VUjDOhg5eUYw7D1iqvd
nHhIqkLbXEH2keDnKzyyYHZESO0hYcEuXrFYOk2hCUUiNxqZakkRwFrD8atbPU+2ult65S1XwNmK
pbwBFVUmUGNlZP5OA1Zp7g8m3HwSzwMFMeXPo20QXYXZz+Xbsp+TrPKiJ5o/fwDOhj/Mn0ZoIVCa
ccmxXcKNQA4+mklhWsR0upRCZzYtW7UwTou4ONG/Qc3KFsozX1zOETlGNEvAu7nV7FtCfLZf4vQp
Ct7knWIx8Q8Gvy7tOQchDryUcAGYy1UyjgqptkTSm5eklQynzagFBWnQ8VOtoI7QqrWBfs7VRa3V
9nWqn73xwwR5w/bUKx5QtzhxY5FVIyjGeDaGQatIAYW4QAr+0Tj75lbf9MVfRKdP2ifnvbssJSWt
LzfG5JUvZAdTfBJDefC+5S51AD/IwlU3E9GjqdcVPJIcdseEj0ivDKrlEo1H4apZJlZYDXXv2chp
8IFffqZYoqMGPbsJVfalHJT52zFPbb6zaEo8asNfbSkFYa0/Bubwghf0ONEpCnw8qXRU9QsE08sS
F20NUOZpM/HJ59CSZYcdELjELahylPXuJVgQbTmnfGpz0LW4iv2P9ZLoQ9SQI0wiIuSiF9Gi6AcV
92oaSkoFAuU5h1EkxWWtcSh2A2CLW/XIAxLALgCS7Hcm1/n1MUB6eKtBoH0ytAvQP4WRTFke0Z2p
C1n5UcB4Otok8zXZkG9/EA92oj5qraux3UAFi6RLOfA1pdfA2sgHOCEYIHagPW9CQUwpAwpRUvLq
3FI4yXir38XWv8sheNSmYgDtUnOjTEUte/sAp6dITeTr7Yg/xX8TcWVrs3xJ6PUmnOc3Ln+GmY/U
MntC+TU6YlmCFI64VSQ7bNIll9JD4R8gjjlvo4fb5rtK7nYJ8td1LRGrzYoodML6QFOUPkrv1xB+
OR9KJd+fBGorB1yPw7uJ7r7raCE/eucDPVSjT50+H4Y4U/oTsUo99WKfNZZJpJSC7zUWpKhLG/Ri
KHXQBn+fqc/zH+pnnBwiaEnDbzvpLgj5lVc1/hFxTKBufOVtAprl7txZEpuQ+iTy/Bvbjmg2cBiJ
YBKN9Y4V1yOTlPv7LoeyzbNuFxWqYysIl10LwKy1DAncHO7daeONEyU4ySocolTxRbLB/KAuKhs2
TV35EylRjaz0Kv5AHZBhR939ZOeP9BwEXbkESyK/mep5VuFQnGG5Jhgkqz1AsrkI8oIo6uiLe9lb
/OgDsTKyG+BnK+MGhayvaWOtqBqeBOBV7GKuF1qx0krFTiqHJFnhL+Tu05uhdAT3c1VbGOfJmbQ1
MwXJfGfRmtLnT/FsuHFb5b/083okFlXDDt9BCwmht2AaFMl+gCupW686rtpVcnHiCimUdLDswRgk
0IZ1Z88vi+q2L0uCE88zs5sZjx14mfpO6NuIJDBb3HkhIV5gyrTUQuKQPRL+gkUa1ct0damuK19z
EWiOoiruOIF74q3x6UTxfvEbJX8eFk/8kQg7FGyC7G6hrj00MZYcPq77z1nd0b2MpL37H+j1p7I8
jM33LX8r62HqxZHvfQf4J+zu8LiZASsjn9bPZqm8FOMKR4nUsC0AlpeWBmZM35PCXliY3WGsStVf
Wnwc3J7g5b0ehzedqdCck4Zp3OZiu132Md7gfePkkWv1bTqxyoLhMGAJeYlmvyQzTJEJw0ERKvk8
OFXW4bKMCJGxQQsga46JLi4W454zhBFDT8+bLZZHu9nKH3VJtngf4uRd7suXNsZAfQ0DCZr2iCHv
Y7t+Ym3cWDGnP3P/5TElIFVg5bNBV2BGGiYGTBhBESKVBeDIhaYDenlsgupu0o1Ae2XDIckNsev3
U372k1DtP0EZIT0GyOqZjLCH/AdKordW9vgF3zFC3rjGcIGfTyLiMoI0REQiSGa0MmXqSOiACE5G
WBjCgEjwcyW/q+Xlw5uBdfUm40ePGV/3nMR+j+JDctuYgNIKKPtLRCuEICo+52YkcIXyLMReSJaN
775/LM73EDXw2AgoufPuJQwyAOKDa8LsasLX32cpHUcRg/sg1tsY+87CvRz879UZ+dl23QTTczs3
6/+5lZBbkBDCAiPHdIYuw575iOMY+ZxuMykf841MSiiurmnXxL6pUGtU8Dn+FFbzjSBLCm1L9aRk
3//99zxzvedyPBL1Bo3WkTp/XpL0gKVVm8dxD5LVrOBhXn7jUad3R9hENBhJ7FPV3rOMH3wGDNtm
4fn7a0/KvwMvN9fykPxcG62E7Q308nT9ARLtRHGo0Ic+5nn0MdlmlQYiWmRXJMH4cHsBp8msVCfG
V89kQODOQrCoiSMsA9CozPp+RrTCmkd8mxqWemO25q3IgSuU4kuOpBDqrRivtH1MWU6dAnAoSzTU
d9B29E/+ZgWDPxu1ZwoGQ5IfEo/ZY4oJE9qmr28maP3TDF++OTbghB6IAh9nqpVNNuDtopwMfVu4
UfhxCdotqRL8tTVTWR2EXU8H5FOQOTR0Cr64bC4gXy84oRb3oIOlbNuzu9n3QH6/EdO4s7UtCqp8
kvEQz28LrhtIE4nzx0Ca1J5+qn47myt1N+jvcq23WnhDIFc/CzNsGz8J2DURBTS/d54oUfH3KiIb
bcIAKsPU//SDEGWp6rTQ3SCXQ1zIPfiDa49tVHg4V5oMCce1Hms3j4gocVoMaShZzITWE50PWkSW
isL+olZk0kxlLOwn79AGTMCcgQQ3vl4q+9azoQcMoFpAEznMDHZLZJIPGBNkDCGN/D0drTvLebjZ
5TdzStFCECbJRDisKz8PMT2vJO/N3SibgUNo0wNJDMav7UZNY+huSI8b2cB9UHXd3cTP1OvNY5TQ
zOz3MF/ujz7NSIGF8J3xa9B2imOWNKYpCeRSRuatw/QZOXH6G5+b8xyjUAPEQnLMJ0RIFYtb02zO
LiAeoX8HW3fwkTdxQD/5akrog5oAJrKfQ8Ih+fcCbDA09LIdbJHjS7N+EaCcYFtPJriM/17uQM68
5WXq8UyE0xlxwrdsPhG85vvxHZ6biNvKf0K8AvIohEeDkMH5EnJY+LLXH/Oq3lH31zuXKKjR/xVW
pQ0eh2eacGfCr6zgiSIPqsFSuj5D595OJt/9v6zm+NP7QWCL68/73SVFN1qOgct3VruAy8M/F5k2
xEnKFUHRww7xowgSVbw4ab36VHhEz71ySh4DNp2Z7PaPa4g6l1WXWzo7zCs+J/nOxrCk+8KFJaCm
RPgKeQp7rOeRu9hGMf4TtcaXLW8LT6I1ihgDSTKlgpERVZtOXg2eWPJGTn7xPBgT7xFBd7AjAIuD
VsrDb1L0U9mnf5xDFRhpzJoiiRQFg+hs53XRdTiW6TN2lItyLUNg4ulunM88ud+w91s9baR5YM+I
m7LPB9sIMspknEE0NQmQizc/jnAOJ6UgHt5UeFbhKKY9Xvb7QTsPF6MBlSSLwWdKN4p6siwjuHE3
l52xC0rjVICKisV55hr2DSm/9YIIY/YkRM1eC/Cp5I5nQFTXzJRCnExUmG+jLUk/ro4mHQ8gPhYQ
Z0UBTUgKXbL6huBK26AfBckLr9gaYcWCa4tiFWBIynd5NFuMUkGKvVMcgSkaeQCoKepgD9fQYs3t
Y6h3Fgi9xpVAtUdnaC9/713JyVgY/uX0pjbOzNfxalu/ZGHiTUkV1We/3ElULkdyPCNYpRMx1f9r
Inw+Eutiayx/52B5B9KbqcKAWJpwnagjGXxtJDI6eW45+tlcFp1Moh43WxpxSvJiycTbwII6Ke0B
FSWeg2vRF76LEcB2xaeqo499umIhGdktU8DymLfjQEujijWGInItz2lYFiJdiLDlv0CMOmBB8BEl
zl4rsZLtyww0twDj/90kc6ZkQa+DrjxGfiqOkntP2FCeaHNhJb7BI7tqmz0eNGRpqfuJ7Gfl3K7b
tN8hvg3ld3qmxmBNWYtU/tFsd/Db6RKZZ6XnsBvh5VebJCz4lt7XN57JjFjapfEfwEW+vYTEBI6k
dzW41AWZKwYEEl31Xma9Aqwe/skqXaNa0EaCDI1PJiX64uKjGgYE4JLeSuZhU9EnDvSUirweqYB9
f2VX3jN9HWDgBjSxmKEu6QXiRBQjZ2RSHgcy3Yfydx7sylrW0cgIse+W1jjMmwBBL0vh6+fOqbqM
9L0VZSoC/7GhpmNQV4uEhKngCC32xGwNkwVce30JJw8oZFQsU4XLled6koW9WI0R3EQx1nJDjkAg
B2c4qEx0juvRx7ydkpsChYNwG7XLwSoGtf/9O6JEPtNIj9tNlkfXRmpl6FEYoRozPIJmoHKr77NU
xby9RwtV1BxUDA0XV3DXQPyikZvtUcre6qCgV6EaTpszU2Li4kh4puRNVbzlIXG2Hup4Zc/SKLF/
DZisO4tEdkNGdF3YUtLKc1v5ttsTtbvq7V6C/KKi5nO4KyJjZ3DouU+bGU35/AQ+ij5CpkjBVDCy
yIcRxN2FuEwIo9JNGvoVa2MJrDawOuNJAvtS
`protect end_protected

