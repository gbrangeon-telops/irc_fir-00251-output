

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UXXDHK9d3YtwspCksVg3cn1OQkWFk3QQ1bnN8kcpv130B5dMgVD8+qx+9EwjTR0JFb8FYrcL/7dg
lIwdmlKGHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lGlirTrah5ntgtsTqcFN8kWYeCxRHbehSLZqyiEvescJE+ORKShYIOu42/ExCc8hSawNVl9qCirT
UlThiM+Fc1evKMQYzaFIzbKiio/Xw8rjRfhTJKjaxdK3T87LnrHcsuSrci+tl+anpBCM3X47tPxD
oNmgZzATBY/NVtZsbvA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UAOAU0ylQuQrszr15mLZsCg4shnqFlxQBAKcqwUoJfM+lTESkAcOosPqKsRH4IbbLlaKiP2HCFU1
aKEFZccPWIgd9WlvneNU3oFbpPCOyV9eZTCX4e5jNTf/7OwRRATKc0mjpd4lxBL9xFrSwNaUKgs1
3vjH77tdesEDAIn5GZ1C/7l3wjwnB4tAiaRNqLY90lB834tlc4mPcP6x8L3rhv5EXfqU4jyJC8B1
4zsO/vH5+VVa1595cRZ3xWXEGVMvmWhY+6TDUJCMhztjp+p4kbQ87UqJz9ddvZWB4hRfjo99Os6I
PqyD9P7zikHIa7jafFMtZu0Vj7u4HDelVYnPyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qRFhWXCy25iIpt8SG9Mt+xW3HRp/MFye1jJpn72azeuP+g/A4uHCFxvcKVhzcuE8lYDqFZ9IBM4P
ZjcyPOhURivBaWk0KosUyfzbkORd8yS5XcayTSj5/d+90PPk5PXVCLjTrcMbg0+NO3tiyKtPpLQJ
f+Ih38e2az80fHBgiqo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tjh0p4bhQQ++Enuq/zxHJnIk+bY5nNzFWlWKnTVXUtnLIlVGko6ShpeQRaCrGzeMC58aHThmj0Rv
eUmPmT2uqc307TRbbuUeFDYMANj1kcC6Ygs+bdXnSkWnOQFu5reSEq5SE7OMIvzdCIaR/FDvSj26
cuj56WGV7WVTg7EZvTcQQsjBPGe7MBQPj6gVbjkHGUTFOQ09cS9h1BaC9UWWfJNQjyJE48PH9w0J
tqmbE8H5AkyiSVZzE1dyYA/E3WjYX0ib/4FRIxCW96Qs02ypuSbfnvJpIyeRwyQL7ko2qezd2p0h
VgIw3omrmALcnzzjpdcOgkkF7sgouCeIApSqBQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51440)
`protect data_block
IaMMjR9s3mjamk7TEDGM9+EkXo3GrJv2F3YqB6fJ0yNEaBUlVDC5gg23nsp4drck6658zjQMmBx4
Bx/Tu/xiWHj6uiBYoqinFzH+sM/7jQZvZh/AjI6XF9d4lcFpc0+S5fusKrQRfROltvx+pkL66uM1
u/QwH//agFbzy9KY/zAZV5PVzHCwmZ4kiIfpY+CVAPLaYPmjEl8XMI+FG3UXlCcHuM1eU2QzTPYM
JXTuJ38uU7wftssIiNO75a7mDl/Fme/vnyTYU+RzCE+bndGhlv7silhP+on07Pe49zmNV/JfzuzQ
zucxZ7yfzpz9bj3NKJhexKOpIlodB37CSj7Iybck1AYEud92wRrqVuFCuV514tFGxbh1nVc6DDBL
2TboJlR15gErb1vNxdukzG5AtRfnRXNc3TiSMrTZxnIqSJCRUAGA6bjqKpZcTak0J1j5buxiMfkZ
vD16MpyIAVc8FxTYdBDcPD0xAiUEVgv4vdoIyt7MZ+2swyodrN31z8Wec+LZnlztrdTF2OhgpHJh
sb1uD63C7PB3Q1iwuEjfrjbLDGMS1qW1VEgqEkaOAYxInga+F+QF6rgM5KbpojflYdQ/mEJVkE2I
2TS52UsUBX7X+T8GLe9n/+mXk7EUkSFcCVHZN0X3SyafIyGviZDSXZf3eRxPrLmbQjjWM6lKShQH
6u3ze4F7/BS+sX4uUx8fMHkb7r2E2SOgp8srA7fu6/7a7qiwqCHhYpyKvx6ahAsSRAk7XW4JLalg
YfA+md3BzEXLMlMIDa5u8RmWLAAWrMOJJS6VTqgyjNJjkGAOs8ezFmRtKQfAaxOzN855sGvfq1Qa
XOb1tk5oRSQ9hYjKbIeU1iGhEJigkcYxRryI7/cxpTD8Wsu81FA+/yf1vs5z7gIrWnULzgBR50m7
XUOn17oBQNOB88HhLq4gPpHq6SvukC8yYJH3GjjdL7EfJ7cRLAsLR3dXsqbuOZnMcRlXHSkeuz2v
VdmLfE9aUxJyc8drazZVycJpHXu7A9OpVEHEy6zaC9wSRCfEEvfMbShBJDCx3vmnfq9YEAHOnB2N
FWU7VBWDdZtcNY+xtgTEXtP/xYwRtKGCt8Y3RnywJhT4N5OUo2rIa1/6PTie6oYxbKrL971kbDeW
mZ1YcVZpe9jYA7Wr/3JfmtcloeFMChXm61XJ/vPnddXr2rDKv6MMU9+6YxRYpGKFMVwwrPRE3ZPS
+B6u5xxF0gPYUgma+Drm1yQQW71t1jFoF9wi9aoQN1HEH7LKYGwSF1/3J+upMW3obbjrkuZej0hQ
LGV1AhoLdRPYkz24eEd0kFmuh9BSeJktz5l5eQid0+SmwVqP1xIMvmrUcaf01cGxAI1ZilKJHZ/X
taAR/La5mJKuXSKWp4htLRs4bz5NXhk820vSvh6dspJV3BuvB99OHw+EhnqUnycZzVZDobkPHolD
x+PajKvY70Dgv00VnuPlJ0Eo9oaZ1gKKppxbEqHWR8m3lFYAJh9oxTRbIvZ8CVYwSRagh6gVwbT/
hhz8hqjbz5cOIV9oQSpEKonCIDmywAgTpCyCpORW/f3vTbwCeFOfkE3mOE4zAVnMMqGXYivNPnw7
kSNge0aOj/yXJhD+ZyiKC0+gUSvmXtMk3AT91PsvAQYMlish+REAMpq0Cs1VJWXM4JEye+SPDYtw
qmh9ehMrzvKzUApFeLIoNoWbEvjFU57GzqA/rzx4HTJgTJZI4sCsd08OGHYVt3gqaCoDXDx0HeX5
pqikrJx7TdUFO23WKnit9FfDvfApO2NfZE9KNquaEzM8dQS8Y9elQ8wfAS7L+mPKwMeBGMRIAirm
70EZhXtMmusXxUZlN4b5lGFCs+lh9DU7/gXPDV3tgVIiravhjlPDq7o9/ifu0t8kp+7MxxA9fCEj
98IFAXn6HsHToZuJHZDZsaFqXZUVeGI696XzDmBRwOZ+Uhy1DppNqd5BXflbEUhBUqtZg3nHpyky
8NUxp/Aqnh9PD8JW+yH3oxBqz3VH58+y82WRlwo5KAzBBNBYjSc+bNFJnZExO0Xk+9BSoGFqlcNr
0c4L9OoQyGnJt6akFPGbBLp9xZgoF8l+KThIKkOS/9obR5uM3fjKOGiaJRrGECKiThqoOe6ymhNR
V15MyDTmVjAa0UdEgMoLX5/W7N/03NQ2wB2PA54AjayxryAkGym37RQ2zZu26iyn8henD9x7VG2v
kjPjYe2lBLlRLDlH6dIWetZ7VC1QsO8IIbw33BB4Mdyy68GBep3W1D+SnNoly6JFFOUMbwaZpqBQ
mkT/oGwGCUd3s7aXV5LAufmj3100K+rCqLvp+1POjC++UcYeYVf03VhyS3wlpSHY5DWMpgjxmH+t
hrrTRa7/Pf24nR/t+zs9E6sunk3lV8RCDoI2yoT67GO6InZ5ie9n9tCyP1LqMBmDUjGWpyzj4txe
WLGSCvLnenzRew4CHCSJnDx2xObB5ipODScG9/aFXQdn1qFJlcuESUdlbege8f/Gi5slYy0dTMuR
pAaJwQ3S0OlvoGF3mFP12AI2IxdzzOPW/BpNAaHRk/kQm6VAAYXxc74JhETubbwWF9GmfahNVnNs
UV0N6Anys8lU01wN/bn11XYs9c7T3Ui9XRE0EiCPALg6TYm+uzxUvi5mrwl5OuDBUQUAs1UCtjuH
Y3s0YtmLrb1pdMf0qjhHfvF4Am9+AL48TgmBKD+QXpFWYGvqs8U+UyRedTrhMb6tE7DIl3xzdt/6
HBwF9yK0DWqNG+mEMqaB93shuTyrFUS7Rg02I1lqerQ0Hn4Ivnu3gTohvsOUzqBu7j7Vp9NYGXAA
La2H+3m6L4KzEnIhmnICqvmDQm2LAy/+rk78HnenYxa2dP1q64vs6Qggy5JPBKOFdpSsHpM9Mzt9
+pkTa6VUDHo+HsliSBm+UlyAMp+NvIy7Fs5FpvbT5H+z/hcbdDQ3qh/Rt2cUekNsU7gFyXWwuok1
s/6EHF37rOctxu36MZUvr/ES70IsJOq/yN/dtlFtVWqtE8gmZNHTkZr85+WW3jAsVIE1sEnztOLu
/MMfVquMtidRBJ7AbCuU0AxiWawsNeSGDkd+i8nFsz+Q4sfXT8merGGvbLlamKiufCPbXQViARkk
9vuxc6ZIRD3ZnDtiFjumqDathgzJdZOiOa1Mc1BBk4DbwrIhrFBmHtNQ2tUSv5LhMSS8cCaQO255
GrxK1OrPWTGAAJV9Fll2wbtPVWXfRxmX5yKX8PoMVwTSCQm6w5Il4tgZKRpGfilGC3W4Kv4mc4Gk
MRRMymVGLSI2Ixbs3JncUkz7yz7FFuN1c91n0ogaMRywk9cJCajK+I837sa3BgzsuqTvNfqmQDsp
YLd8uwJpfZaSufv4LAA+FxCNMrxALSFjfdvH/q4m0tvixnqri88xXj9xIGKOzusbed2C+1cMODtf
H1LzGWYfdzUgiPYqAZns3GOIDkWLMvQ/PeyE/gNdOD3DgElZ9WIACE75AVRhNhOicK8qZJni1YsQ
hSdMBtvYHl2fxKyH/NdA/A7MXRNhx+DjlShZp44NlOQ+9oiUrfk4fMlMRMxB81h5gdAWgIEMbWEG
BZcloCPbsM6uVj4vYRU2YI+As6C7Kl4y7/0X2eJ0Yom1xPcHCfNN+Fn0aZA/lXMrqDuNGN4G2xUv
PuqIC0jvSIwkoOZb7dfsf5qO372c/FX/EMCK6Ugb1OJ+OxW/ihGFuQdhXFfqN4Z37K9hQKLzqdPB
ZnAf8xdrDKsdwX6HXguh8kvqWVkDtSh8CPj6ymKjOdqgX3QNhk7+o27RoGjtqnTBffl82tmHWqQb
kQQs0sBEe2y/shs6i/w7YFYvtyDVPeGvtRODG1bTJIoMaC08OnruhLWN/RSHjoekqXAF7uJqH45p
ojVpSWZPnl+U9fa3H9ck0pRlYrfBzcALE/XdA2ZvVicZef9zsJt27hGEwgf7PQmLVvS91r65HXJb
tbh8WbSfPZJWUCDdyUdnz/U9Vq0fxZhzzHr9B8WiFqs08pFysIsAyqYRreLNpxYKbl0W1kTAXWOf
snllpoOPRZxMrh2uOZbWbaIi0frrW3naJF8Evskj7g5txXlORx5Frjf0nzNK3szS6MN0QINsnSAL
i/0bRkpMCEgK1kMOh9Y3aQ2Ic1bLo95l3GSISdsqK5Sjrl1YefLjMBjlccJZHoXBTgFOM5swTSyt
rLB3zl0XdPxRuF3jnHr9e+LlQN8QIHWQSIw7kFNc2aUmwrR3WtWsfnb2IqfOouaF7mQSaTawGVyF
/qaM6/Q4TSjinMhEKv4Xx7XVbZk3M7REUJFmCWtTxCYVvmHX/SsUkBH0RGvb2rsSVB4ovaTYfvfX
LI1iWRiChHCfgTeJ3FQpNWLfniLF+uQIxsSd9U9m2JVoxJcXXbzz/vZHJzCCOt2TgjdCCtGUHnE/
bnlcezaAszauQj+mNVfteeyvn29x4edW59fQWUG2jCJabGIQVM/i5HfLfEiRwPI/fYsONILZ8kJI
q0mhdcTAvxmgPdg695wfw2dFacRyKSlAxXKktR6a3moI2Ovt169VQ/pEC4dlxlVJLmt/TpleGaBD
uNob1dm4IpOznm3aFb1ip78mS85qVkAhSy1FAUKz0TOdqaw3X8EpqU2R41D6FypWuXASjbCB5hDI
w6SCvbK1WNBo7LNDXyqFv2IGYmHcBaSl2jLCL3mW4SlP2bTO7FNuOsWi0pBir46pJM3Qu+Y7LLo+
3V59aWkrx0JVC14L/0JvOp34SFeY9J8HqqSYUSlT8eyVIcAUg/vbtcRHrXrT1p2K6uGxb/HNFIJQ
zSS7wQ9aIv+GaSZMSuDHfnaD0HTvYiUTB5d/tlBqYzqWzjhJyee/lb78h6UeNPJeT2+fBfre126o
5tXD8oVrqKXmWdsbktAlnikQlqRbtM4HbHd2TecTbVvwO1xNlfrfVf7844G32y2KYGW1FBTCG+bX
p1yE4eiLEPtFL4qY8gCUtDiCKdC3VUXzn9YTvSLcEj6xiow6jWo/ZNkQyll8IR8jKqzvUvPsXIlg
NTY+EdLB9iuoxtjrs4Ho/KleW5l/Ziit4E1ndBNvrDpXkyS+RgnNZ7P+Rf1lQBmGCndxQfvmWuS9
G2ZSAUe55PvB9m486vl0toeqyhg1MkaRAOFieyzUL7FzxwfGK0fUSGc8QB9F9c/sV5hmqUaI0/+B
qlbP/EAFMh1GmaZEi3ffskbu0K05ijeNwZhTFWsylb+l7gkRo7hTXjckKfLkhDTHVNOj5G6DkBrY
32HuIEM+rYyeFrjY+5IisEUcE2frPQiNp2oMFyuO+cUh8mUIKmB322niZawvJw1CkB+jLMay6tfb
13wRDfMtinJIXltpQuvSqdboO7+HxGv/AQkeAOHxMm9IWEigJxanSAd8kO8GXNZxRIamvOZCscby
ViWYNQw4ULS2EYpze793/x9YPDL+Wif4FaOkpicBVEKUp8rOSJIYCDuSvF+LJPfXLHcmZQvTUbNC
3S240anpPYJOUCP2CCyRm/rkUgcYOrWrNILfDMqq9F6mK/eeyOcHggoabXkQ/y5BtantMLmIX6kI
NNahSJeUNzEYZctHi+/K0NiRmGDqvxiSKiDqS5BcZ0ShUc2lEx7V+zidsfwGqWp9AcqiJvVwv6gV
a0Fy9G9eaU3XHqZx/ynzjmkoUrrolwH5rl5GLKu2/WO0rHGIIjdaTvVHY80L1MlgZXHjizHMgrSr
b59pdI2C0XlCBdzLH5a3lss95BUZBMU5ZdRe9eLaNk7nOiPxRmjbKSrogAO10MlMhpcrEIaCNgQ6
V1SmsBo6TNyEnZ/G14B4U/8/LBKBfn/K0i41DrC4zmj5eyc49O9sZZgLjd4eLzCo1NQMNMJnkEeH
Ua/rtj8lSjrrtoBtOcDCrtZorgvqJ3v8WYPPN6fzzP4jy+qHDD+NUnQVUQvm9afxoZ5YeFQGBmVY
A7/OP14Hz5O0LzZJJg4wXe78islW9jeNhJ6ifdpXHgEmtzR56vbAECoEkPxBRQffzkDbrdJkj/OO
BxeaQdOCWi0Qx9C7uJi1F91OCTC/E+EBOWTZlY3iANMbxSgFKvmNdsd/kbD2hcTFo08AfVnm+VOd
tcvOXYUKWM3LdocpGjmaBSsf2Fr79EvYghxGOfuiIoBB1HYPBv7BUFNri4vuN97r59PYIEByTN8Q
6mFpf1eu7i3zvSrfPLHq/9gC74lLhpCRD0V9o9UQ1Dkb6Izl/5iIxnkgUv7I1rbLi4LS4cMKh2PQ
qpT/4mERtOXCDwXCHZNZKPMHRxAMXdU+TZhN6q4euA5/jlcUPXSQFB4wfrRBSLFMgDgu5uD0vvqO
ZF0p1pPe67pKSQb2N66J2r2O56rIRk2fLhbE8b73jCIxoHYs9fJgCY6xbC8tQUXz84tNslEqSLGt
7bCdX1Ncs8LDK3j2UvPUsqdMP+difRsmilGjajUvfWvYs26S6x9mbNyLrwjR4T86wIGG9sPXE9aK
jqnneeJX9aq6oiSpBLyGCV8kTjwbYTXn28E1gU+Ep+1jzxWdiX0CFZKcMyECWSGHY4QaHweskCHg
JcPGUul5pHM0F+UjGkLoPj35aJYhB4xTwiaBd66AaWH5W0uH3bUYgf8spssi2JcMq87kjifQZb4t
VRUbtnfHyDVTFaRm2CWiE1lMFKUPDPDCtcy9oEfEPTawyimuK5nKqKWHqS+OAVPG2M82zvz+wT1Z
ttCcvlkgCPc9d8383LUYZfQedK4x5dU7TilIhXoupDkuUmszYNcMAvYWIC50rKc2KTnQB9X4AU+E
aU2p4untwJxohpp9XKNA1nZvXxfCunfpVJvepWc5vZc7nv9klGcejjbBAMmx2MVzzYuDrI1GNPQF
GR/JhZTOzuW8MI30rVE0c7m5NhY1i5Op5mNOLZ6RhkeHxSzLTcfoUPUBLPLrTgmmJ3eisWw5Q6+U
mHNMCQ9XUVexr6SrqNGYqSy7iSd/9T/AZTwoPN2aP99WNH2kwlkRekQgDlHd0PKCfW6BSLLZ0clb
cAIpHzLgPLAq6+sQN95G5eLN8nki4oWFz9ouazSvc1ZAKOHMw55F3/9xma3OyMX13ywyKMkvrQGP
B0LiFZ01hmA7oKVirUnif1XSz5DEvi43QGYPlVDa/gJjpx/awcN2V7uqdyvetYrvkO97otW2phKp
QWBXWzai7IQj3VxOzdLb4klujUpEVefgq2rmIxVQuCTtOtfxU4IzFZIXU7qfVnQmfVZl80OU+0mQ
cfFzaemAje93XtKFgLu2Wgul3FFmks3zsxnhoR6YS9rVx+7JprejQjpehBr8pf14vyEF66JxI8yK
PBTTyHxV1mbJrVjbUzYsKKgLkOVdoh/2E92Q/inivdu5eQ63qBllsLEOt7U/bpnw/irCSPff9bdR
Y7HLKL5XLt6GSzAd59Q9LVnqn4MQLgfKOy7muWFYG4g3ZCNNz1/i1CNkHKtzITwFz4axd5oPHjIh
EM/gKKJ/uShV53YzcmIxmg4tVEdKug9+DOpjxUhl9CFYw6asPlF092oC5gEExD1q1hfB72xsrRN7
1IOfnhAxQZEvlddha7LFMZE8Aa+Zpz9xXOM9aNv9Y+10zsTgMloGRZW8RHO5OhGDTLzCvMRvFVBs
Z5ek/bHvdT+0KFBEizwF90x79xAzbMr25ehPpwIWs51/xPDhoa1dxY6qSVVsU4RpMnF7ao8OPWBP
HF7g4M/Gcy9qnuw9dtHjf1GNekNwbpV6RI6+kkT/NOsW7xfkh5rMBVfvWRJAt6xqvU746dwzzPo+
KclXnszZ0V9CMJdG1VOlSkt1sOEcSFexofJZdmH38qN0yIPpt/hrW1NRTUKu8IkZrJlzoBvpsdgl
BpRoLUhmpktptEG1NfOahJInrjjR+utUoaYrNWSHxJaX7BFKhQDyozBiv47+agzA90RpR7ifTa+N
xi3BoYWfkOoEBCYDB7re6lj39vZL8GBCvZd6MYLZifxOuCSbMc9ZUYaWmRwNRbqVyL6QRT+azrfZ
fLagvWjPcd7QvON+gxorFWETPIQs0X0tCp4qiq/3vFiZYAtgrTd9xQ6ZoB2TlnzjD8ZVArHeVHMt
aMQLpprKn80CKGOf1g8yCcXiUMrLr4MBola/kMei8FyEqJ6E/NHjN0OtvX9sBkmo+QhEoVjiiX8I
3BQrfj1NaN2L+qbYf0RdTvIfGZhYtzNGmT3mnK/r0eBACaYeaCelAOWqbovdBrhAPBYXEQmFrpMK
04EAR8wLe7zaM0oWwGyR5fahJcxjgbap8eG0RbmgLPIwCpXd7yuEFtfGpSFvLvvKLCm1gt925zaz
gaaeFZipcjWP3NwVtxU36LKUoJH1ASBRvVDMH+PERs241dSDJoa2klkAbVo9soFRmW9lRIYBMcjb
3IIT5myGzpci94UfXdEAzcxJ2QzLlTO9Vgw6dgZsh7lwvDdwtaM//z8ZqzIsC6a44QkrOnZ7lts1
dgNqX7riivdCi72O/Q5XRR00UVPl3SWlJkphZum/QvzI9ZGTUiW9fsbb6bCpH6kTO3fbP9F+8dBi
3zG0eWFGz8kg1CDISQO7YXIyLBPw9pwj2Fvixi11Nm4U99xhaGrUdI64DQMgQdfv6cJTdevxiJXt
LSyxBqWNYAA60e3kGfxk6g3dlUybQKIOV6TW06b2HI6TVeZqW51JT6Jm/MJshH5a4WJba+nY/I9F
NokLKMh/ZITS+El1Af2IxylGq8DCj2uCYhJWuXWrvsIrwz7boQvoMQSzFctGUsBD2hFR5Bnv5VwT
eAT63BHfdj0Hs8zy1nTEOz8OcAyZuUh452VPt9TpxiDwItIzhtUKHhxGXhSyYG+u12FqLz3eCENZ
y5IUjvDAuhW66sTu5UhqBqbgwQIxnNvik2agFlyzh/1FH7ieV+587L0P83NYbJLpwG1W9ZGJsuoy
QIEw4Xo0Q+nhS2XppRNS4h/NCEIoIPI+ireHsSFRdR0n9s/M0IM/qNlC3fBDhD6Hi0F5V+ZI6Joy
IABmOoWZCTDjhYZHatzTxXgZsoxSHe9l0+6h4y2ijnwa7T+vz5fLR3X0RvgGaoH7UF8WOWPbESmo
ARt9lp+JF0f1rBV8QyNzyzgN2k2ts7cI0i+5tofGYjrMiSNgT/1vo2/C5r6opmzfVUsgglrRfCcJ
949eNapdLF38WbNUKjNFEU2MRNPkP9ugzPYUZZXaEGUulIQspUZthvHT8Cvpq9XNlVr/yueqcdwu
lIc/81Gmcriiij6OPTSrdGtQWdBgxoeb9/iWbrpUCaUTdKxKDCBauop03FJVHSRLi/VKuP4Kezyf
ZaEVVAf5wemz3LzfmHlQ0+sOMRl0HQ6N2AWRrFiw+P9jEWlejD6JoXi/5j/Y3RbXryMmJYosydYK
xnnuaQ33sNp9e2hbuiZpFUMMePxynnLJypCVWF2t96rbwAyYz/AFeUTpjB72bt7uc8/wlnaSguhw
ooOzBW9cuh2dUDd8IjuZB0Fsq5hE4c7YCfo/b2ZBj58Gst5eDr6gH9/S3yA7xubNg3GoyhdS2CPf
d5Kh5ndXedO3LKw2JKqgsqhNl0aATeUd3sqv/oYoa9RbVUy0NXmXA0rc8wu8ATraVjXma16FZq1L
uWaUFKsXdI/RclmOfH23Ed8+tZGCGB7VGTfI2LI//02LnXMr+h+cNeM+29o61vgRG1vVMKIvn2cH
WkkX8yAq7BGzL7gveIVSdmSmPNkCybdnH3xtJ4srON6tbe8WZ5AcIiu7vHyp2KZ9RDhmUh0lhYA+
pmK1vgjrbEy8twZI135SukQI3cYhd1YnBZh3Tk5gXsjuT6tWmRhQM25AgRFFoXV14mIOag6F8kOK
hOtCxupQIZbtKXZQr8pJycWuyN9yZYt3313WM7XkgNSvBOTTwbblWR0o+1S+HKIVL3aUqxjAhQdo
rdgQxgAVhOz9OfZoqqu347cOGOvtk4BlGaukEQl2zbgQWs/w1AOdzA6Ay6K8NcFRgDToJpSl0EvV
PDD4yFYTdoRVlVF75rq/RdWGctVUvYreq4ivmlBKmr1PzJdIRt3fAZgYtfTWzxqOzce6KRB0sfly
aZ4LnbBu9aGp9FF3xBBiPMLDuqujdLKjfdPeqpzWQO68v2xctlm5O/T01hJ96IXmPc4Ebv0zjiIZ
+LndpJKijTnFU1yavtYPm+Id2CYwp2Y0/g9lecyf9I6rrA6pWUnC2238SymIVEpCrqzKds4NauZH
TnQ4jTN6dAJ5oaz3ShOY4uFc6qBxUUtzHTvAa9yq0mbW0bdyAW7L7OZe+YVqudXm9um4yiFLgtp1
/s+ERLQEMW7a0IGX6Q5k0ql0kjgkZPoQtLAdz5KHGKyNLEkMZbGnr/aZMrW1Q1zgyhnFx5BAx7RD
dVauR/yt2m2vK4eTdNKR+hAkDybo1ZXHKOekirE9WkQuBrkHeu1TP21shX3UqmIVNb5E1kmXJYzK
I/L3RiMZsv9bF+mdHALT9w1iC2z6SBuXPnsPSMX6vhV14Vwt8TDUVds3JC+CscYoFIsZpq8v9Bj1
etGx+ojMiHO0VYs5gK0NTUOXhm4oumQqLCvo0Xi4gse5GeMMD4vQI185BV/hEVXqAzNQhd2kkvVE
vZFaIeTi6dPgLAVPHkS09FlmqyPsaWlMZLdKZE2rtFmFXgddZz5DvpVYTRLz23yt4JpcDQrUbKe2
yeXU49X6eepx+aUlfAQw0U4gFC17ef8X6bX2zdBr9RijfZ0B8r0M4BaUJEyfBoM+A9oO4t2FvZ/2
fqlnuBYNVhUnS3xYD4UDywa2Pxts/5RProLO/+p0MhICI9KDcnpNY0SFXL1+ljOfpel6VDgsGUfV
jS2s/Eg0ULD7pJAF/IndvrcsQqe0znSuBlWKtxceMYXQK9gaRDtb31NRK5SUWI/uqyH4s2ACvMpS
auk5q3rkRmkydBBTeXZ7uXyKXSCeZ6PyefsMdnPlp4fU14yIH/1BS7DeLfuWKs57xxOlfNscOI39
zL3ga3KxqD7D/ArSJs8fT4gd0v4sXTfxRfkuELjjD1TaTTc1CTgCKZ6PbpQf0lmn6NEtwZkOog6i
tjYKCTvKlnriO1fOpaEMQUQm+lphmqujQm6dFiKB/Yv9rHkIXgIj2vyYAOt6yFT7t1KXu/Lb/nbC
yOgKfuhWBZPHxYqht03KCOuILoqOYrk0oyojNT83YUGVBuDwJEEuUAl1gBNsaX/GnCWhmBjmj1ef
d9sAqyX8/8Sio35vioVEl+qb91qDApnQ7h8OhHTZBQEO7SyicKyFNojCjM8KGErwipaVgefRg/iZ
mho2gU1B84H37awBEiNkdjec8Zh0pCtxX62lXe6ABnkPrcGIuKSKd6mpPP3DRt8lXDiVU0TGAgyc
NwaLTUbIxy298cGf7i2JV2XKzykoXgM530lBWTmFtWYuA3txDk5ayDyMs3c9M+OVKCYnKXnnzoNk
KJeciS81sXSsGxkiM0T0Xoc3DRFiZ+kpzgiLmSzxzkIfxw+u1x9el5I4t1l4mEH9gDR4mRscBtdY
DSf/WHYeNm+YIHBXUBpBDNkhFsYCE4K16mLTOYfmxs5Zj2g8lN57S0y9pGmEOj/4UfQ3Ig1KddPM
ecmdtwksE1L4+HGB0pRDG4eW2Pa9Ig9qjekQ+dsdcNuw99OplJiJSyn7i+81AgR7t/D6UpX/VFWh
LBAU+uRK56ED5edUz676mGWPnvWdHq8nge4T55KbsB1zD5LDgmCQ5bxCMwUOFdyD9XltQc361f2Z
F/XzAPYtrJWcICBqMrECgA6+om77WnOpfGjCnady5n1aqhw9Le73CwqGLbQUuL8qbcMooAbls/C6
3VzU/qh8EEeKtd5wRZA8FtZinepc+FyoQPb1u1VpVTg6uxDYwQ6FFCy/CHhTAIlSvyUU4Ld4U+eU
Rqa+3JcnDEj1VBXI6ZsYvdCrvVv7rBdCSUnzY7BfVXNpU0kFaoNOXeUuRNYqwVDQs3w/INt5i8FL
UDrlNnoAJul77jjzxMIOa+osqgCWlRRH7saplcIopN57mInb5fov+BIYlqbDSX/v/ixRZNbAv7ra
UF359cBv2/1XtWWWkKqz6frXHZkWlBFSwCKHGJGCQJsv1cV/rBvNCpd3AWGTdY3Dq05W+41NOaq8
npGmgm+YXyD1HdMM8XU0rHcPwG/wvwg+Nn8Qpxok5YsU4KodZg9IOy4Q6UtwHNEMn6MgP8YACVig
z85SK9H1q1AihyLKA3HVuRR7B9yTYWBU/LK2K5A7aJ8t95GjovSSd0deO9swB6nFNcun0RAGBL+7
6+UvHK6ZV/9pJRQg3rUtcZso8bJNXptoa1a+ZRUhx5a/U8jDa0cJARUHR9ejV0Sk95V1aTwUV2L/
g/V72HwGSFkz6AM7AGxQOKXCqqvDNqQj/oKDuegTY2MbPLn2sXJRuKwYHuQa9LkSjAMHts4t4ODg
paGYq6rjXcPughG02Nik4pDGOFH4UHNlaySie5oqLC+ZDYWCZBkNCGPWsriRD0DNBgo31taYJJtO
iv7HhMn/rAGGSb1pM9Jvwumn1UH8EbLjB0zun2zDwm4q8ZKj2bbHFSDzPQ+V1y9SmIcxj9GKp0kq
MImEtu1x7zL/OeaPRm0EcRyWO7FU7jwmuJmSUuY1/bWwG5GQh9EeOEm91GY3d9i0AA/kIu/kI9fW
siEX2e0+8uUhiOJuuFqTk/00tRGJmSZTPdqEsA1w3W2FguPxbkUdvd4rDQZrduPuOxkrdgLEOhej
ec34z2GkH9Ba14v3/ReF1CmQDNXqg2CN+nD07lonUIOkY4HJTq+T8swqQLNE7rq9AfgwLVYumbOe
yGgz27WJzNpFIEanHRrjoERX9bS3Kb70Sj1Tbj9aXiDp9MKxArVGrDZkf54fEtYhAvXM4/0+WM7a
c+VKRW5cfG9DgCu++Wyb4hYl6E6cJQtMyLLXuoVkKJp7sIzrO415xVJw6x8e9jyTr9EwA5xG0+6v
a6sWTddmoGO6H4mPymKYhJpDdTuTI9JWSh9wb3YmBSPWugbIxRWoR4fOZGC2yaT+Q+bVMA9mjh5T
9ZwjQMkbFTZIKGWivRvtylL3n3AIPTMhOHqovNdUIp6g845q8mLF6tCiFCpdIbZC1fEU909OfKZv
V6BAVh7bHNqLBnEwAmrEQAmQRa2mUfuMn6eB2z+8xAsjEcJ3E6jE0OcxsAAcAuCXpx6GVf5hixoc
myaPiatYMuDjlt5/9vRU/u64tqMA5/nN2R+12L1L20UhZPW5LjM5Ba3t4ZOUXrSFghxKyTr9nL96
aqHcscjHZI948sbO6IM9BuXbS4Th75HX9OecYecfgG29BSWbhSbMiVz8GfASgSvcwXVEgx4s/ZCI
ht8+3yIjXnidMM+z8oAKsKPDGrvib5kohLDdhoNsHaHXN2OMAntMoLQ8XSBbUBkWQZ8QTAUEpxsn
MS35smevgoZ1yescMtA/xpCVgWN3bzgeHSLJtS67SIPuz1nRBH6aS4/8wwX521x2natcT1EvkAwJ
9I94rvGKSd1oxw5MBb9a+Si7U0hiPhIyGHuENVBjrn7gJ3OGLbkbFgmxk+je+gRu8zJcJYonPTTh
iKimi+c7uNHWz9rLDB/4qhEv2uY9rkD5fcfb/HY0eV4jUYSb4OtF/qk/ucXTt5yaVn1gBlfgdYVW
doeGmp+YrOtcZu8y4EDbL7plEaEZNixJKNRYOZiHTcjQ0f//jnR+VrKrehT8LnNY5CKTexKDC6E5
aq29JolqcF3kRMnHMVkLaAXBF/BLKcNFjtCIDaFho91efdmHuYhwABOtSd4/uR+M72w0NOTgMacb
Gxb7NP5I23nY91nDZAA/XqBhMqnAuLjDRRhTNo+4N4LVoJadSNqjrMAr8IEkhwzvizkgYHMzCv3L
t9GevuJef7IYclS0Z2247Sma4u993hQlaWFPfOlxWyiK8yketQVOA2K2FWtWI+JCqVFRI970x7Rq
rF8qqBDO7qnY3i8HBC8oW6/LkqfVDUUFnJQj6mPaSg5o0Xat26sxuRHNtN3a6MXx4lSsmnOSAlSJ
Tm+IFPbHBJhw3bJsiZio+54DjdBOnI7MFtwJLsRiqBPuERKsYP1fZD1GK4SB4DUpi1mJzajnbhzD
RF3AygwCMZTGxh5JNJsE2U/XpZY2PzdVgvStfcIdNhhwZNEP+PCDHx/AXEhMhi776cXVfChVyUbd
6uv2CfVckkUEa8eooWB+HnIgcC3hg75qpYPw0vrescFRk6/OaWuIzWhvROswIeBFKRkcub7KtzeL
DZUDRrdgm2rmPr5GvptG9+Lxk7zXcyy/JkZy+QscoYnh+6+Xx6aihz0Zes3bprRSJ7GjURWyn58g
GQuE32bNcbtMtHClVHLdVZJzzAA22LEKBP5/mb3V+3FYcaMAFnTJcdXsKDI3u418LWJkhMz0JofP
SITqTui7QYH+jKtyojAmGDlxbTEQEcYjOdssiS52JP6NEcVyKken0Ho9REa2UK1dbj0QXckhtexq
fzUtfWBrxFMHVupKzSWLfFvsqb0ELjxWn8hmXtsouabso4jS816Aa4ot9RK9KkY2rzmW5xqLTmFW
ONg/hTDoKGcTblV7xwPMUvFBZyDWS4FJqiFzJaXj1KWc9mXIJtNjJQtCevGQTcE+T54zwfihTel9
8pjqWOg4lxJg2b6H94pvs3yyMLNciSxPQQ8a15b2Rv1Q0uYD+sh/N1EcqaDCEjcQahc1hoPKrA+d
5+55PP/z3lyiJIMqAC/jaD5QDkU7BGyEJIryS4uFib20Dcf0BC0Trsnc7P4M2/dIYmrKm8+otakl
C8MjPk402Rwo43kJ3xqG+2Yt40eTIJt9lAtYIkBfkqPXUG9ZUNy7RKO1IxDQKosNPAVIefrrfvVL
jYReYUphNbbJ5JOyAss7oJSrgZG930panZPVdJ+XG+gVTK9K2GF/aLvdkpjdmfQPnZkyQHJvfdLP
NZhICuYIDM6X3fd1EpimTe042yzCJwXN9PMLhFRyckK4uwuEZR5D1GqHUpKANYKGwEWx3fWctkEm
AiPBXTYjbnZc47Zqp3fcM3qUZA4z4U7qRCJl8etHV3h6po3PBPTAJJRSVpoVbJTDlN+G+1XG1Cgm
rw1WypoGdRKx0d/3GDmtIy5RQy5qRJ/nS7/0nNcYBgxuuPTtmERS32vcfLI9P8UnNjjfPMKSMI94
Fvt6k3o3lO573Qpo7OQdcJjHHFP5ozYkpVHTugXOiquJ1uC3DhUJmkL1UoSeOA7zIh347feu/43h
zWPComk3cL+9o6PZ4L/aO0TE6tAn39SyIA7MdivdktB1OOcOsJTiTQUdeuM11BGWknbKSmGdL2KM
ex4WdNZwIEcFkkmDAw4HaDGOIhqKaTb2r8c1dV5Y+GKOb5LKJ7rtuUKTIlG2CZ90CzFM9pZncuSY
KK5N4OUXAOk2utr38fQ67X8YSr0ofSC6XhQpku1fq0rvISE28Xthuns7pz3tUicmupAoh+9B74AL
3yg/eeoyg/QKAn13joybiUYxCbvPF7/+Ah3M1kqvamvAxFgbCogUlK26Dhc+NsDUdkSrMVa2i+H0
5l8AWkzCxN+kKJINeiIepPfL99WTHFlJxt+Kj4aUx+dSj4bwjyhgkKIiCm9xZy3hdZyMdvJiN+q2
ISKTRo0nspmdtL3bQK4CXaUAUZAnwp4eXuHjp3BzCN7ijNqHbMhHEy5UC+YaXXgAQk32A9u6DsHK
kZhcXdRNpg/5Sk4lSqJqBROa172vjc6CYklndLj0Q3U+T/BDSZJrRaZZTF0lWW1tGlRlcvWpKmTe
vgxGLj0+S/powQNGvFi1+8QSCNbbn7AV+BLw0SQOrEA6X4eADcqY5Seu8sgUIhTqavDBGrq2ujtB
oNlkMh3uqRcjUX0JQjyrBNqI+0VDNbJ5d5fqO172QD2XokOpDsjVXXbDHjLzR+gWoKvjaFRczJUG
epQ0OsLoZNo+C52TpOr675gYKyoZq9R8mWx74o735Zmm4svxBo/rur/gKukdhk3fLHdLE5Pydxhf
7pY0JhNvPh0eAU96WpFAwH9l1KeVIqaYJcTIrYflDYjC1jJMhBSZfxM9DtMorVSR4y955ylpFwwp
GKaxsFbvCiQu4ddqfIjYKw27SoxAdExUdLEZhcN6a2UxROisfi4cb9hhMDkFoaewph/Z4LjNRMjr
oEw943pzZkIKB4z/29ZshFEtGxlmuLmN6QneuD/MLA/ZyigqNvqNuhZot6LtYRkW85RVAeEQWDYe
b0B/f2Uo/5xT0rqe5eTg2pvjLVQxWj5gbAnjcJhbJ1Kmg5V4ScP/ur2TkWmnXbNDh2qaJ9U6R7lg
SiHm1mJ92JkMD+GFo+e2d7v32Vt074TmOLMBH2VFtY6vxloPXaanUaZ6NCErdWiecRqOAtm6QKX7
f4F65dx0ObPhIgWdFeIJJh8rHEgT8Nxk+/QWYXA62vuMiivsus8HW680HKRwgQ1wuPgj/wymUSzQ
szq9IE5TuG6b+kWdD9Mtf90DXmX6RfmCVRIAHa+uuwxsFx8Gbsi9Iyf7yu0PFn2ZaseEIbiAhYVM
82wzh8rlLOq3vt6wpNMFDNltSvdCOD71SSrgceYFmAKbGGwl5uwTGNTY4R3g+yp8RpAZr4rZa681
CTPw2ygESTfjydor07e3Ni39u/Lyj6I5c+LKZxjaYpFuTA22ytd7YQUpXNYYfguv6g8Z8LSc6Gn5
LjKWLhyisrlgu8BPr3np94HAb26pSF859Y5ovECbTxEZZdnovf4qufulJV9QgbJfqy0SZ7BtDoAz
irMVH0fJiIeiwd9Zq3SWKltxHWoANRYbz4yHBFdvQfQQOOtgZgzOshuN2kARnAp10V0EO/Ef6Kre
5GHH5xjDr74j68TKD/7ZR+xVDTnvaFdAv4iJ1/RjbykZjbJ/ezt2TI5TQPbIB/l+5dF4gt72wmmE
ZgUPYLoIYiAx/fKkNsTCxOyMgLVME4dVIaIX0VRsdZgV0FenWVuM49X+ERg9uvoLrK6Iemnpr8S6
CEBhH26WZfrnbs7L5Ek5ZsKAvwM/ed+RwyQ+EWQ2TR5mhHeKc3RQa2ihdv+Oh5EmgkNirSgbiupN
10sbQy79qlUCbgR8e7lHorDNMS4RK5VtYoRagmMU7CWck5N3dXGp4vYQyN6TiVYLuNWa2/USGIbR
/T96PzNTe3R3mohydws++0K2rKuhcLS1lgNWyA7kuVRXV699lJ1SF3npTMqUvkhnBVI7IP+utU9J
GbwZniSbhMODTQpBIEwE3K4ZSbULBRaml/RfUVIKJJI8Sc9hTHp0Fsn5lBb6GUk5iDyI3aKI8y8B
4nv2JwbHAgo+Vrva462jAbI6h9uDIi/RtJDtL97swwOmou0aDHWJbvIucpQOHvsKOE4gZH1NBDb6
wg1pkV6Gm+Shjiu9JSHVJRmkD8vDyp+N8e0tQEtztfUG+0Jw/LbTGywwaBiYwgkDk+acvIUs+OQe
t0PncYHtHRK3S9953pah9JJ9BwyQG74eCws1ocWay6FL6CPgSW7jmPNLHtLzcxWCD0SMhX3GOGpb
fSZVRZKSz7NaKFHh2QeDmPChzBWcbsXVxQ0sHPzaYb4rPDGvi00rH0u1o733r1+UKMtLwZEB5YMt
p8ke/vgpFN+1On7+Bg//UFw/acdqSC+oWLTF6M+6hP095ZdXQ5mOsGV+bLPUTN2RSfp67FbpZ48m
3evYARqUIgkD3uDSa4UHVHV6YEhkgdz+SYSazx2mZN61sO3Kw1+EMPN88MLPS2xT/xp0pON+ShuZ
D8jJYZOvj2YStIyF+b2Rvtvxh+W05jP8Joflvxqy0PUMdbQIAwgP4Ol1l2c9l5yBQvI/rU4IU5BG
grnoYNeX8htMpyCyZgmivnSFEXTLVvQKo/DeSax73J4LhdwT5k+m+I8WkMaaXG2mMt0sUxqVLarT
8EKDIBaSYR/AxWE7Ihow3GWitHXr7JW1bNWs4zvawEvGrddyppgJ0gTMU31fMTEkNRoxKmwTzgL9
gcLHs+9bWncjKQAVaBPLTEa7rb4Po2/H9ezTNpY6gd2rCBPq8YpvdY13HsBCTDhMhWuAN3j8fPF6
CIK3MNpOck0Pm06QWTWcJdGDsVU0lnWqmS3cIlycy7guUwQmihcla8vb0yLUIrYUGISpkDojpDvn
+jZrl8azje9qwhAAebKbn1ioShe1FrHaPETjalydW61xjc2zv/v6x9jUIwl0eVNoU53ogaU36RAg
nqDYi0PlsHuNTR1/zqKmhLgoB85i1BU5mcXn7kQNOXEs7jy+2bIyUcPWSlZ/q6zs0CJ5JjUa0yG9
+qCjz4bLvAyenwc80vjTWIGWeJButpTPG1LLUSNOsHVIvIc4nOJjwHjZWNyr/I2I2y7kVht9rBIP
y5MI2yYW7H85/oYD2B3Jroohwey76KXQ5poIOjIWIRXFOMdrfk0b5GSzHkswg4sL0J5xFNVWD5Dr
q8NKuLj/Dq9Wxt/FXmVJ9xaicb474ESHI/sdrsdjz7IDwlJbpCUngPQ0OZwNh9qegVoHbfwscK2Q
FuWOV3hzthKIv77+/f0tfZQDzf6RL//q50p64ZLc0dIzJHqxkZNfWK+tGvMKB+sFhGO+WvygGATr
c3HbI2cc53XvnasipNykwnyGnsOgjcPW1hCuWM5S7t2nkorQkAKnEJWL7N6lpxiam+WF9ebmMYjP
jcYffhigg/OsBNlnspZeys2kTeBxlmGffw3I3CouynwRDLA/OqJkl9GKF30oLpukseutYWs5m8/Q
nDLnDVUCyD2ZVi4N8Xmf/fkPuCnRcP+Er+P77pSmVWplkhtnwK9xDd2672BKm3jgNKjktMIn2RiS
knxVDaUI2srBMwrFH+iplY6QrJV0WkVq/unHweaHMbLgKee9zv8qYqTnm706JuIjY8yWoi1jq5vL
rFw1w17gUITRj8NZCyOwG9/UBR1ZbAqipfEPpX+XmW2f9YlFZInpKni7cAsdok9NIBXfvrbAFyzr
B767Zr7z9Yxio+VmjgKfD/XRKqI0MZZ9XgdASMNFowWO13qKO7p5+KbqAIaRr/hRwO5bDdswnn9d
GlwDBTJlK3ZoHe3ZIRCQ40V15i8Apw0aFGAAWN+BsOelXai2j91LqFtdQ6t/4zWzL6CqbiFBVZtF
jFBxuCGMl/jGBXDhHoz6Nd3MTjO9w2AF8tS6T8xDQ2iiWfdIh+TgwwsxYVlUxZ2lO/x9IcU5rGfO
a50OqVTKnesbnZDCkKOXy580AcAIBM2jj/qQj2MTwoxn2JfZeJG/qZ8cVL1LHuMxVL42+wWOxYvw
x6biPCJR9itdZLPe9O7lj4AOteLB5We3jtpv1Ad/rStGLMu+JQnMbM4BdWqiJOSlbbsdHHc2RK0X
c+9y99PjD3DLae4qwzRM9m17rwv7UPXFuwpOujFJ1sN9VEbnxf0nVtisBA5xyOz6s7ptlEYmBQMN
esuLfTM0CTfFHsEbRILziG945jLWdW2QsUgnQad9wL8A8xb1apjenrRFwOIn1lYB32uY2LGgqrfV
ezhGdS3Y0hoKMgFAY/KxjA+EIAs7lfE5pVa9L2Cr481vu1xdzc0X6Aw0kyWSAgKAIiy30lyVBMto
pj4enarKbpWbxws7pRLY3cvfqZXg2Ni5ZKmPdE/IA2W9hfc6CDiudK7ObJK+1PNqlIldr0PwNY47
4vL2eFNUHI+cBBD7UBbyW4LNs+nb/lco2F2tPzcH0W++24b9D//gctpRTiJWmAVnP2KWNlNy1MmI
M01d79nOD8FtW5S/Ay1dqxpi21NR7v+ySz2705zdFsjIc3UR6VRnyDpPVwQ/cZnjaszC/oCXkAI6
FaA4KJt0aM2nxqU/gHzGABesPozo7hKk2u8+zw5BMvYXEQVjUG/aZZoHJgjp0ji5SdyyRM1d25e2
eoBbR98ye5tc+QwfvhY41xP6IUnT56jgwMwrasi0z1nz4i+yw2Yen2YAj30ydJcH5xrBnesuN3I9
Z+M6SGIminlF2CHV/NUn+CpDEIfmtlECgvnXqCy3+GElLrQggWNrWJRWqJyQr/Iuk2kHkfuRqySA
C+YSq7ElIsn2ialMsGxT5dNR5QShnvqFjFMWOVL2wBcaZLzfo+/XgJcFncoG9CZyZplfIY250SjE
FmaEzE3Bwfgcv/oroQdZaUB5TwOfkbEnTX/ufow7AGdNpiUu28gYscZcCaJ9pJgF6raHuqIARbEf
hRqKw5awcohJfFr6Lmq+z9TPtf3HToFo2B3vNuST5MJsddA20dbYlIBecJZcCoeQoeY3ZjzFo9ti
cwHfQ2WuYhRg2E51O8SomrAEzekZCLWwYlUx8/RlSZ4BNYaL/4SlMxIbchJb6kTzOxhuER/ci8/3
Yh5UTDTmRNglR4xqNgNtFpUv7db+rh4TIEV54Reed/xWM3fLNxB5P+eozSbNf0YW0bDYu4Yt59cA
jOm4Jug44nuwlLiT8sWfp71T2GVgx1x4vlskJjSzUuPkiPY+3/ISby2qmjj6idm7xY0jcg7uXLrn
m1e9yNTD9rVEES8sY36Si189ojACz28sT6QleRTXh3QXcLvdDSa53YACJ0G9b25igPyDamL4qZoe
3aKiBOiXhw1UlAjmI/qaD1UOycHtZytm2b1Dtb9yQP4zClSHtLhSRHyUAuuvoVZfs/juSY2aEMdV
cSaw7iSLvIyFuA3IVwG+rfnjGdiO12xCY+3sad2RqQTuWhT+1giBxno+dDwgN/sx2dOP092i3HXd
qNBws/11vu1II2tfYXn5FrRBh6GVlQXhoNeuzQf2bXDYEmeVQgfzRSMecXOBrGfAHTuOUIX+ACIW
5metIZaiM85h51V3xmFcYU7ATZ8nNFI08MW2D72DAPTakxTpjeGnSVkOWaXEdk4LdRPskyRrDHG3
zm2dLU4Wg/9VZ1SjVKzV90T7ouWIPTqAkKxWrHBV6F/Xx5a/Og9PplMXIqo6YpwvwYVw9welxlB8
bjaH7E/CcM+p/euO0n89DTAeFtFGdW9fWZhx4XLrueWY5L0ClrySHkrnEl98Jt4rPmNgbGO43xBH
gywQinARF7F6vMqG0g/tqSYog1lINcuhHJbVz7Qq7Xzzlz8ARBsovZ1zs/iX/G13pcIBPziQ/OEK
xudZMcG0q2oBwjUGNONrW8CHQkktenBkoH/A8cG3RaJg9xXZegm+itKdS0ho/FTydONe8kfxEnw+
8dSSJvW3wo8RXYehmpxbBA4sjydA1dKB91/0DbIgmZfEpTCTKFCka6Mi7xn6XTVzaUVSTqzCWUzw
mlFx963RALi+uRRf9RGouRk95NbfyfLRNcb0Dgx43RXRCaBHjexHy4Y98Wu+7WfLp1ALYmj8cD1k
AiVMQPcMhATsOD6meINdR5INcCtxPXgwC3wxzEK2wLpuSZQuiq8g5IuyYhFQWodvpgdNMT/AWt7g
Q4uQzxOJLson4YFn/Q2xvpt3C19ooyosRc1Kz/q8h2l2IB18qnCZ3ILx1y7pGW7lYfjaXmnnRLF5
6KHygz6KxTajnYZ/W6/vF8Vrgyi/JQFPAc3HWX0Ygb1LV5fgUByMaFXOKmbqVVi04o1SciqlF2kl
WtUsp6yACT0mp+0+ADTcxA09+hRcNbfMq6Q3EiPzZWg7nEO/5G7nrcuZdc4gtze4W1L60kBDShEQ
2ki0WrTJQZ1F5gTYL2LEjpRX5VA0rMSu9uV4RGLVVVrKmsHYnb9MzbfPEdf6TGxIBU99cgxSh5Ok
knId0/OO3g7ILTu9LHMcvhvb6F919Q3fVOGYZWjCOAo20LYwDtqdsMqUTtbA8KCr96P/py2w2Vg/
b9Uji02CdJyH0RCrnpquEdEc4J67hG7DaLkpGElQsOUueCBeuG52C+hcFNpk6MQWB6c1EtyV/gDQ
7pDu1DXu/nT5VN1VDLt/wQ1bCiUhCP0Lv9ngiN4cgllzwZdOMTacRwO7YlD8qnDJO3mIwvbMuE/4
a0qJfM/Y+5HFotvBKoPNiF8cP1CS+0xaq2Ply+6JExl936BRvWJeDmpH+iaORneVFMlHBHxZado1
whxPJjbe0VLZjIN6IKIoCVErnMP+aehkMDHVvz1G1h6M0GnMELDFhWWvnbo635ZPyMgR/eIWhWgt
2E/ALjXw67IzwQ6Yt1I/cyvqykuDqiZdF37vlVmae/5yjgVrzDAAm3mBJX6Ss9WPRipkwVB5wXuh
0rrB5VsnoWdQTBgeGZKz1ffGrieNVlFIOxWUIsTOe3o/y/0XcFXHuG7D5cW0SGiC1IYMie/YE3vl
gqSpjG0QvVn7FcKATt2rOpU5qUmg4ZtsXDqqDnPF5zxSJ96I7A3Byv5QYjICmMiv70rTXvzW50Xk
vUvnb6OlTt0Vf0iE3Vt8LcWJJjYOefWi7qQGXYaHMOvP+K3lxY6EJhlJRB9dBXKerbnzeOWOyWPT
VkUaNXDzguuHgemBy1GQNw9uBOp0lNRkh54kjJUB/1iMk+8oVNkW8PFtThHhUba70KbRTc5jLdTB
c0djlrYOfPfDvzKTy+vehW6C/jSl5VMtXUbBOPcfBrm6AfDtr5ONF14Ta7dMHJTS9laDVzD3IBSH
PZJDBxA8KGMLD3AY12DuhdrtWDSFwIsQm+RDHTnMk94l7nSFXY3LDQ+7oArIfj3eYPrxcGQKMITH
U5haj44K953ONkc461u0qMkeG72V5n4PU3vHTNiYOt2kr6Qau7eo+oh3N4w/TpEehN95zHJNNqA9
domfUqPhBFHklhmTJb5fJI+yIN8weVKG1kuEEKe85ckPyfQtPQc20FFMZbKv8V/vdzNZ1y0W2QwL
aqQW14/iLx9Kf6zOFLsA78dnlsjsR1LKrQEcCdLJAHJ83esPLF/g9JwSSMVHpZFKSZa6GIXMm8rw
V5xMXvqRpunBNRm5EFTloByGfam++KxE7n8AIXAshC68CWRdl5MxA5V9edskTljSpZLdjRyReugY
sYsoFwO+8GPLVOkmd4t0wCYYgyNAnuAeQAnlz78ktnooBoqEUZBL8nJJgq1OzMmnaAaziUvOg5cq
LdsHx3qywOxOiO9m74Lm3DTY2YzrIiFj4GTOAPfpmbIGzj/YRq10iBIisej9f7Rl1EKPWGQIXexX
AiiXJssBBfh/whWYjvGrx+RXqgIZkT5j3bpWVy50ORMEsZ5RPUqSK6nEC5/kgkjteP138+wc0SFY
bvjxB+0/49XS7aiD7np9eof9HU6L62xMOi32xDfRSmbQ3zuMnefB57j1guiUkTW6UdVqJrCta0u0
D0K5sdQKoCPTznqQtUzdvNfB1q217YSNX3bZaAE5WWfiW3svg0CpQMRfzaTZfZIb574ahTNCAKVY
hcX+UHM1IoGRBJ+xwMZjpTwsfIcLI5aFgLBWNlZPacx0foJfHzOqOg4OA8WqD79yYO9EooPaFvtO
/NQcuMFTyJ+x8I+NTT8j3im9mLvCHN8PocbIOzPNj9CR23nqefE+ScpsxVHf6Rk0mRA2NROW+atb
si+HcZiwy3KksAwGySF5dCyR6xwK8ghojeB4upgZvrXqgYM6CaYHrAv5jfk2OPvhJyEdjIUn0z9i
+n4lgOc8IeDwrTOw/6NCxAXw4KnvBiPjRdUWwYLYl8mLrCYkF4XXcE91VsmsexSRLG9BXIpKfbP0
S6+zuyV51tN5OZjWuBUVz7xeajmOAxHGzwFWm/BeCgwxp5fxT8QVlK4y2U/N2XfzsNL4oCZ/1U0Q
3+sMAECZN3UiYIc/0nvoRTcKR939nVn73z95YbrcxruvFR3rMCj7oMkpl3TWJp+EwY614rH4ciBb
fZqGSv36Mg7Dwli8TDWmhyfzb6zR4OKS6bjfLxZPswmQGiHlpHkzRpTA2zJcoF2ZxQsHLRi6wajP
yhIxZ5SWthaM7gtmYxO6NQhO7RlmFEx0lAAgo7pfjTwnlkUee+t3wejkUfDyS17FbfYutB4l3AAi
QFDV0G+bU8ZU+sRbCVmibusBF9T1COS2Q5FhSeeqITP4k7cXPSM1Cr3knTg2TU00NrulufBiDPrK
Fsq4ipCPusNb1on4Wv1dljcwn4kb8YzEZnoX/lcNOPR97DTwuHmfVE1BNbUiCIea2XlBgjg9wWtY
kBLHuDAj3xpdPC/bULp9qwCuTcvwsw7yGu28Zpmful5j2h3ShnpQwju5DdNw53UBak8FoIlAegcC
fTmtG0sCnItmExPWwUFIaM27W4aYRiYsFReYyYuhYOwxMgMoUsQ5cTUPAZZ9uMn6SNzDPsNZyXAy
rBpNX7jb1lmXWVydP0zWgVw0hlir0E4Z7BOP1+VnX8/tq6GI/y31ZWsMLRtLGVMmeayvgGERnXxs
q5HRUV4aZ+sJ4D/CFqRebJy1T0E87/UYTeS7ZLrBojXlj8/nk4o0b5FqJ/gp58+GkVaqISmgWmRF
WExx/edJlphWcu5Krj6qpT/wzxDhdUUYtl21OZaqTimfSgjjusLVmtGhPFgcj4ojGC1sbTaE+BDh
ul4BhWQffkc8fQq7lRN3lQoU5in8XhhM7tRCQqYc+GUIp3LElEjXyMjU3CmN2Jocpb7iP4x7ZCl/
D8vuznIHBi0HXMnv+GOcH8L2CGEpxttsNZTcQl5Yvlx/Fz0+xixJn3YZLq4PJxfyCNKxEjwFKidv
AWfts3jtgmZrNjhXLph+p/zLQiU4fvKgXFc9+ZdMtXL3wrI6GKlvX38IuYSI65xbQQSoc2EfzvCC
IG+c9eSrJxKkK8h3zJQPTsg48/RNaX+RrIWjmhKvbCoBV3xy0Fv5w4CWRajlWuLJeXBOdycrD0Ec
i708dn8Pnx2Yjf5uFTKh8kVQ4xkbcyiL4X6nM2FW2zvm8oII95TlqZ/r4Je1ZR5AQCIMfQr9K6h8
f1pF82nTs8qRRzrfGYMYGQKqzigocmScwut/Pmz4DSD66CLSkejXStNVYpdspuKt03lC3rX7LEzI
miM1xCv6lJfKruB2MK/mVWPIm/+fQfvHtNoo8ZVOhdj5Yqk43X67HtIU7nX9vA5rf9TeJ39y0Q1M
xhSTBM7gOVodCqryBYmxY3KdCJFKNuNjX87QUgakTeXLKRRknLT12c3EIxrBiYkUU3kTf4gpi92U
6+V3pa/gwSroPlaAB3sP6/Xaw0MtXLIVCiXbs8lEfuFWQ/1GCrz0ffV7TDHfeho/rB0Y95NWLFNB
WjrvBClo2zVLbRpqcQPJtOcdpGjeXknLgkox9BtCo5HGCRfE540SG/mN9NH30xbl9N0JIZeXr3lA
79eWXebKecW4xz1qhTBeplOSRaxRy9Puw8fBSSRSxD3EKCGQPQ5Wm7kFAm8h+rFLU9KqEhxMjt1Y
lgQOAf247edj7UfT2Tn4J5gJRogoWioYm8EHeSwkQRMeWS5I4laR7pS+99w5NSy5Z0Qerln8tK+k
ajGUjEnw1Ptf/TCxizajkMo6HAsEHyyACMPbZskgyfBq3ILEda31Gf2OTo0yUSpoiQ8yBcynOhkO
KvH6yy7d1JEl8qqXCWVp9iOCyvvAcZzwY5PtA9d//20hELNFV56ad9x0xGp083kyYRgatYDE2czv
jS5Rt7GpMIS8jEjp70l2BJyMnYDxqaMSuFoEJwMb57rlITepv0qIjUvudr+T1MtK9rnQrvZP63BU
ozUo2s0A97Uon5X0+QiDJ/mj7t9u8SPjyL4ryz3M4H2YovO4nmEIcQRfMwRgi7u1CMo3Uv7s2J9/
fXx7pgUGwc+kB4WOYZOmmjjJMPne9j77eEzPC7vnz96LB0Qip5DCzDXVOImj3cdCVd2mxCYdEROj
S93tAiB3THvwehop/5Z1YiuiQ39keB6gjw0Ikl3xR9nxAZIwW/j5f7kQOKpybR/78TK8oUdKBvU8
AnMXdDg8GZ2HF9tmBOumU8Dgk8JUkMbQhlqMX0ntjkGqt03QobDGkYJsO3Cws6IKz/RgPqTRk8yP
8SXCiHAFQv+I8h+wUOqbuUALvko7xFW/jjww/bZp1gXtT/+pCuIzvgsxPsdf26oIchlPfKBBTuM9
L0GHkFkuH6zh6KSw3KTacN4QA4mUh28uys/LNcGy9W3UCQtMrQEH45BqmCrBoE4SXU5/RsEdBa4w
gz5XucA9FvQL/PCeE/MIINXhikfmRihdUP5uBljGCig59S4U9OOsVLUQd5X6lHWz0NakpurCB8n8
mAZEkIMP7AJvZ9sUvXHb+RNC4Ih4wlq0NIDJVq/BpvBTF0AUGxhe3Z3F2OcmV683Zr/g3OUEiyKN
AYT/KyfcgQ2sdv0k0Y/RDUMS6GKZ+q5LonOwXjvgyhHA1FemtZ+Qwx7GZ/Z305/gKPEefAdVS5ca
KXTilom6aYnIUi4exjDL2zkr40Hm58aRZhP7oaZh/EssbiiJWQyoCkqC5kqiFraTyOTfEt+qYQwS
M7XDwtPhuzk9Joztl/m4ZOjxZAbLNj7F4zQCzhty1REwh3BmAFy0AVOLP/9QfvSakb4fblB19yd7
pewn+WYPfbk60czqY3a1AuxKkgiz+7lQJB48ME7k3D+6NF3oASxxwqt3p/yoc/dESBMTLd3b5ZME
R8oyxX9Og3/FkqeJXLCHsO1rqTwK0si1j77lHwZ4caX+4oWw0feO39HBHtb1T6c41tmw6cHQjwvd
DUgLsm9FWSh1p1AjEwlDg2wbCowRaAr5r/BkiX2fe+FEkxizbhXEPQhroMjZiHJBRtL2KwVn6m72
DmytTLX0CSHFY9wThC3dH/DkfnLHsouOTI1SpoWW57BhUKvv0UguFKcStw3LjinQvHyyoCP820mt
FpMtFtbwXkj2tDjq0jDdDYmlekx1gFpkIMbb2sN15XWiHfEGKQiLTqy/5qQC8EGe5hgqAQ5/XJ6U
ZSfu2DAQg8xWjFQx/lCXfgvo3yYk726G4UXyZxuGHorl8VKlgBD2MpVgS/JS+aVJcznOrsmWe8YY
2Bw4F35+RgpuOBmcJbCx3PtnmVvRPXH7HRLMEpm+EAYP/X3YMsLiklvE7IbqewaCA4GugrXVm4H4
aNJEUIEM2gKqEuX/thqxpo1H47W7DR8VoDMxVBRTJUExD6ry0ivIQuclNqg0za7jOQenagQHMJ6F
mL53Tdd3ss96cnAdhFLQExFe9plDsUlDdt5ayjRLA+eFQhKZIqojmLPRyllnI9IWetNN0ycYu4E1
AVm9pEfLGa9gXYeaUfRygHMNKpinvRwkLHanKJ0bQe+QOnazRv1iokjKKLhOC15wCSB8jhRxYohI
kxnHChzVWjW+0iFKnKR02phEFMz7htH/Sf2ZYHiYUmq88CG9edUzPEb5z9XwNSzcvrSz7R8uvf6p
zu3f09zGPxTdiDOZQYNNJ4Td3evVUzoeOxGvd0imHG0nC5W0RsSN9mf/KEp8oKeokUgvImjCtHaO
RglQRcUiQoB0PtkMrq++czv87WsoHBBHcKumBPivUWao3zTNTqJIxahVWl3nGmSnuS50J0aFjDbZ
7j06KU91D6OZSSxq7oaMr51C2vNmr2lU3sYOIjVfxuyPgr9tiXcFjMtYWoVxMDw7dPuv1EfkQw/O
XHMeSuS9ZlnaCrxj9cCsC7kRgOXXL06RFzdCnoCCSPMJnTYODNXkVajTpOs6RE2+JERn46h3wsuM
7tgJCj8iFt47od+VpGmHjwwHlo0eawcnC/SS46qnC/vocbfu3P3bEVLlE7+eJYRvBAB8P7TjtWbR
moY1uyslx8262vbuy9uXG16n/mpbt3serhh3vUPh63391wZCNmMdU10sFJWHa+Oekkcdib3rhIei
nrlupthJV0yF39eYMBYNRCujKoUTArM9er9Uzo6vb+998CM2YWQCpplUYuu7h1No98VRfftgcx3v
jn0/TFdHq2ttR/z3oRxFlFZVp9G2gPTOAng7kPZnG+XUzQEiCcnUzWxpaiWgAO0xGgB8jUz3rRdK
5mEaOvDU36yhwFmFA3KDjm6pH7shP7aG+v9SijKHRF5/zaevhuXJZJOh5OT7yh1xbscwIBZTdFuZ
Dq8cUhEoIlU7Y0rgaCXbJzqnvKPVATq2jT2mR8mXvS+u5M1/S+JCbAn8r/JXa81dgz/3Sv+o7t18
z0yfJKNowcEMxKEU3qRUfOx1Vs1rBTNggbNpa7y5p0whgSuXFOokqqDnnpJRKySZCpT7UGb8CEtN
DhVzsey91mjbPDXGhVtoYYWkGx1fRxyeLESqnJZFgLRpGl8LgqCu3rY4+U3IPXASqw0zNGMYVC3R
yFh2KHGBNEp1mFie+n5IoOM2pnvOhL4axub8QrQs41w2gprYsjX9LseRSUmHSvhrTkAlMHiNZf3a
mCjwE1CXNTvibb4Jl2GpBycQ7VyecGBMidN2sKvz31670g+3uKCP2rYsHTQlgKqTmf105tJwNURt
6wIGQ6CZnNiul+jqR+A2GAbRlXvhM9m77Oa0ob9YwhTvXnK+jNRO9Jo5wj8T4CMSxi1DJ0Y+u90X
sMbug5Cab9EABHqr9LccP8Yiw2EZMl0Zz7hHV9hK6vJhbx+8kGUUD3Li0WECSslpLRoMfHm8ntxM
BZHgF38/Ygcl29uNUdudSg/0s0CVrYbd+eCn/rfjnP+GwFlA1EhYRTtLVk6Ff7lwO0enEQCHjp9R
x6ju/6ZzL+5Y963cAlPAZOPUS+qsN3y4wgSOKrFpaKn69VUmBqVBC/JWSS5LCx66PLpBR9Z9GliC
YZLBwCfcHK2zc9q45kaEU7QBnwPArL4r2yaK646CoZlCmHko/JCYG3vyHZiINju7nNy5xcT5d8fm
tEUwyteU920wZeh6mXdlwwEzONcljtup4xXekBOynBpmeYkoKpx/DAc/yD2gdds9MQThzhXH2+1b
dX4FJIunXWDlL8t5gKaWn2sDQM2bMv49SfgOFR2okN6vZeMiKV9T3PcPnrUWfFHTeZcvhwsLlDEJ
Ih1iSkeT0nfXNh6sDGPgjieSvPQ7ZRr8+ut9HlFO8sf0hD8j6uaxEKR01FPwB12pFKJU2uC5UbFi
oJqbeJJKbHfx3rcgCAvBDeXswffxm61cGVB4PjCCVju7VsBi8nzlzjWznD4pqapJYlbCxQtEdDty
zOtQVO4EfSbnAHct6Gnd44SmJsLWCQU7oAVj9aAGKwIxvwt5GXRW6gz0NFzExlHH0k+riH9NK+H9
lch0yqHd5haEaAjMdOm9i2WMb3hojMfttFh4/jGVMkkjlpjEHt1dxV3GqWzOxIHUgqOXb1u/N21C
1HxD+KUbzQqKp7LQNPjYCk3aIN4LchD3DYxwjI+HMPxvX3tb+pw8eg2gGJ2YFSUlNcNCpDGbGOJl
jH62Fi2YWR0A/WnFOrT5xDl1WbRrNilr+jwxZbJ3uwmm/MrfIGarQ2noO9NHW34QE9IGQQ9VtSm4
DJcUbLur6TOq/s2SCm58N+M9unhgn3lF8WJWUiCkxZR1nwC8aacOQmX2w5che9MKVFfIbKW92ioC
idCzDFAFWpWo1lO+XVcgSaGHLeIg5gYM/3HVR+cZC4wzmfrtTV/70ibco2ubwOo3ZMy6IUNRKt6J
52qBopthQ+3T7pGqhOGw7EfyfUqP/BFyoiDp1xeaAmpzTtqjoJwl0DNQ5ofgmhp5/8Xov6UyVH+e
+R2SQ0EjlhxzGv9Cq9iFBblXp5ULb2Q4koOVEiKKWW0dY2EI6xrkRQoDc1tG//CBo8rPIcTNzWzI
0hoOXKM/o3O85rjf2saAZAweYhwHLSkkVQJ5Ql9obgGXKf0UCfbUkjsthVyKaDxhQWlRVwd2Z3cd
wcGQGm+Oxiiq2/A8z1LuwSho1mb/p6r6h9tc4QNgHOd58nlE2VkwxKKb/5JkPn+HzmNkj07e/H8Z
buft8P2n5AKiln6bij6FDi+M12I7KNdteM6IgbDpk4MtFdxTDTcV+1k5iL9R9em5LG7PZ9RmqkCX
vPNOeurhj3co4Vnmwjv6l7YehzdQ9m3sZRsVT1wPMkYigWTWkvOVygF39oZUMhb0i86RbUhgRgkc
Hs1Zrx5Orq+2yfnybeAbATzpHanl8AOd6+KtGwN6MNOsyNcHi8HZwGI0t1FTNgB1gU/m2ENi3ZQ3
WfxACIYtOmj8tbnsc0oMBs81Bwt5PH+TR2vIvpCrVnRoG180gI1LiaOa+A9EDILlYaBnMVdDmkrO
UBCHylM0Ma+zv6XGcRgnYSKss1toYK/yh5tKsPMim7JhRUmFyvXB9mCtAgvrvOmPVJI1U5ekxeao
J7cmad6ZnD61bYyZ5HHnsKyyP0Y4rnE5BifAdpYHbW50ShBvFl+zzs14tQU6CmZnKbVpMt70ku4U
EDg5TD7xmo0aLPFlj/pb7znF3W6LaOv70N1x4wr+q37wQV54n20Q4JeW5D1Zb2GhR7h3K1Lv1reP
/M3UOCjrq8qh+Q0EtqH1bnwtfFEGr4hB7m8r3r2SSsD7mkSOhVZ/B1Nb01QWuUr2615K6wkXtoNk
pXaK1TQOxMtJiODUcJ01iwblF7oXqXSTUVoeno8xI0946dy4JtbB3il2nR2aG4cUuUPDj1/qfZr7
YMCsviqdL6QqX2ILCzwWTqXgC9Xk3l2HtsrLTbPe09Hekt567M1+A9LC8rBDJLckfq4/9wuXW1av
Ej7tJLqiMPdFB9okxIOesz7JGJlFU+28RspKqM+EI1xN/CrqUuxtvUwO8hVn2KF1+9S95rrlvsp0
dv3deWeb/bvDCTrVRq1bDTN0te267KL9wfDvMZO4V8Gp5T10582wjCHdbGB+dI1xSy+9HT1FG2uY
pV88M+RCVW/coE+fBJb7FdZsODN9DroCJ0D1ivoBIoNiwDIbo4yJdUPSfB7KCu0lIehQBH7JWVbw
AIOcMK7T8cbey0IjZAweAQp0+hE0MPghL3sowTTWh36QYMpPMFsjF8gudsrz8RWJUEJYCp6Cdv1V
idyivy5Q8M2Nq3eBNFsAvvlHFD1Ybrq6Ow7LhzP5eFhoxeYB/PYTzzfiyLTnwfmqzx5ZNqPGXGp8
BMsHTwXa0XXVwB0f+NaiyyzS8g3VOXscAa+PwzUhOaIRSmkdo2/D6VJYA6YyrYVhwrkNZn71foWh
1/SON1AEzjR7jxiSwIWDVrCnzCsaMa84AXJahgVUjVJs/vo49yoHqqYodT2yF/Xf9hBBPOuJoplB
SHYlJeSBjzxyrAegC3dI+UB1x1P9zexewhobR5apUXWMQDkQHifwGV0wKyxVhbz6THb1fN6Q47AT
90eRQVplpTL1Mq1Zfy9zWRQssyZVvdj/E59IkeUWQBec2vYYIR9m897M2XPHwwNY4WlDiESUdXRh
6J0J0aBlYADV16VEhQV8P5sqpMi8+8mdx0GRmZX1NR24Y2Weat7MQ6ZkpuTkl6doffVEz+zEx0eN
Gv4dM0ENQFTkLSar517Fj4gJEJYdjiTYq4Lw5vnKkHGGJVA6VddM5REaJJUSPGWvk5AdPGxMnS99
VmFWQ8AMIVlKLjXFIE8SV4tduzvQuiBFIqPjfS4niZ7SUJnh4Gj7AthD8jMqmcayM5nmDFyfIMnH
SdB4KFuS1gjuJPH7sm/joHreXc+Jf/bLgRX9YkY7xkQ9nb7jTrJCTJq//nnZbG0DsJLbqY/5394t
lfR6napL7BOLKmalBry45sl2VY7OPSHdUrdf7Uih+2gwuLZiw4LRRv7LxqotCzirdWx/26O+/rXF
ogZSZ99WyXUxuRXt3exYmyQXmtV0Y7hHX4F+eECYGZy3LCiwJa90ppDZ/Otyo+O+h1iTyuCBP0pc
WcoBGTgboKyV5UHFST54l/+MevqNVIbyW72TPnqY+wgvf+1ZTxioTvvydke/GbKBZLFpXjy7LeUR
alP9GDVhT8bNFbx4CCKS1TlUWMF2Jbkc39osVup9QRvTJBhM+KONJ1cv3dQX5bdQ4GVvF657qkAI
dcXFDFwokk9bn1NxDvbCscDNKFpmluFwMQ/6/tYKzBOsgbE0MUfHCFB9ZFPiYZkJ/O6vZj30gpt3
LVoVeN/rXOEBAw6hSt2yYYZOBYGahkUZlxXO5MlnMRyUMKYXBHxTKzWbyPBF3RxMddjQ28LCS5Qj
rop/DfujHlcc5KK/X0t3Xku9p5x2pxDAVMOxSvtsJ0SCZnYaA3G9kMIC39xhQQoeGy55b9WUJ9lz
5DDj0dPOPSe9hy1McnQLMniLH/PQ3yg9KOvMEr4w7UxuDxYVv+7PI/AX4EgMHKQdiO6J45wy0HiP
XQR1BSblexSAXN2pWwy+S3+h+IdWgIUFH7rSf6Y7CrEqm7PZaw9/KnDgbqoNnHi4Iqd/TaychHkL
/681PZyDVhXKXrd5mlsxZ7yHkbAonVnPaDKGNB4eyV60BUCc7jvRpCu/aAHhasH1vd1X8jkcFsHf
/kp5MnwBpaZiMkhrruXs0GkMZWe1M7v4W2XPYE5/uyJ6mCK5QCmJBcbCVb/JKp2EMsWhekwQ+9qf
hMF0SSqWH6xIbj8bO16S2Xtr1DE9ofHhWSQl3tDc9wstRKu+zHhepnWsoNxT1HesV/yFGvRrQow9
ui2wUOz7GpIUhJk8J972W+5U90yCnej5bgEDHU7CoZY9T937xMPSDcEVcNmxsN75ysxw64P6CA/A
iQYWl5xPEsR7Nt3SjMhZD+fp/Zwg/lzBcMb6t7SK29qDz4C3MFzwlWivccNIBd3NRamdHf22uad2
H7lQ7GnC+0zp7PydvmO4aVQ/ZSek7otH5ROlZ41QvJTn/fcxyJZW7/WV4g7hXHfEMi6cXA8IyKaj
mOlcXla2XOWnZqjJB3TqW0ofCWqx65BKVkldkI2k2KOSxrLqGYqzH5jLyl7RuumIr9gK91fVANuG
SoJxjYU2rOSY7sin0wUOprh4g3wGk3oOkxXrtiQsGh76+e4SPo1m4m5BpBVKOL4UOlCL8Kt95oOD
oLG4xn7wC3ysuqNBcWJCIk/tQV4VgZXfa6/QJanoOnMvqZyjGzXpSTbEKJw2zHy88G8ltcsdF7Es
B5o1AjEQxZu09PrG07ybiJxJ1hPO15VhxWFdLChGdDv5wODeKrGe73qTj1Not1WOYQ3R6vyC31wl
pjK7TVt7rbZLddi8H+dvPLTl81wr1NFcpVD5uJ8vAZXC4bgtQ6lZASnmVKJj1kI4yYczS5aTr/HL
obi5xagnxEEdn1kCF1HCnGf5FhTZ3Oo7mZWCIy42koo0IVIeqytUAP4h+SIPkafKht6EZvUXLPBJ
mhZN6J3aGIF9o2AleUbUfzFB55PS7okaEPhPNWECzxAvuDlx76nPto7EikdmXjEWyiaLJle0p/A7
JuTsRWYji7DQGaAd5KurUKnbv1PxntLbQGFf0d3+KHRSU4R7ommh8eXIKPyMPYuhcOsbEgT/FVnS
7+eomTP3ljsHgSt8MyotKURgUoKCb7IKqmRzYiyragzTc67hHSiyX6cY0tYZ78F3Yk93iCzZPxzc
XVd1cnNhyWftlJlg7OklwIR7hPFMLfD604fZyn1fsisHZF8LvcpK9PqLXo1XOgPOAqvUyINA3mkw
IvHDk0cvDkvzIyW6GvWDjZzeiJcg980xbGJTT/TledyPaNbOhNwreiS7JUAgSD+MUBxxEF3xH+zw
UJ71srUNv2Xi/qRxdKyaiUpO34JanmlqRSUFo/x+7h3FUZL1iLuUA1sH6EaAqpqe+zNK/xkBdCPO
A2BZkPRySO/cat5SCCRB+WcUOtCPDwtMgmD449/UEuMrcwqmzTwV21BG1tl8BgTVhYdBWE145+Fv
HxSaVH/nnMONXf4QZ8yOVDaJ/xq+7JB19Cf0PzG9nQ5/2irqMDeoJj5lFWJa2W7bmZIO9IuOmnBw
CyaLltqJT2gWRY7UNCkX8j3M4z5KVpEKxwz5mxOUYRtQ/mU/74G9Rb2DjL7YH7irSdkRCDi0zfdt
W6IERuyldQ9aRz/P8Gyypl1CrvHy+9YkZU6jZm4cydjqJUYQ4n9PKAPtQR9hVS3JY8iGKsYLTY6g
202KDUBPz95xN3kTFZwfcazfsaAB4x1VXKbsuJ5wem7SG77S5q6UGNVdLdgCP595MKtkXpdCMOps
5GRoY03NLDEX3iUUFC63w3ynjFg+39TLO2VuMJvvy/CZPYtyBbg273mBpVTbW6Fyc7TcF7XaWD1L
ISzWp/ag8sxsoaOafMeAHGfEjf4200w9TC9uKmJ+gHJ69y67/UiIn3JoX601GmWJF6B4ePgqGfHj
xa4MNOcRX4+AA/A7mPNbmePyMsbgR9JBKz+Uw2ilw43Rk2SGQpDfr/lo5i4JSpmKmda1mGn2hg84
kL3BP+s8r2RVtcQn3sOuZpg8kl1RWrO0DgNptNCbMd1bxtoa9YtcF5wEG987Ge1n69TKAFj+dNgq
Cr0iJqSmNxjoyO0kwtO101IWRIqTIQQg19YL4go85/+lZGPjJOB+Uen0m82XlpJZOC1TIqRoUJ++
NgA02/EjDk687Brnm23qxbX7GgJH2OQM6L/W4BI2xFsnPH35V2P8hOWy7EHqBibmNMWvSPEAD1wb
PdxdUuoUxXpPrkz1/gQH63RquEeWzeLlAt39pjj4xBBNTY9C6Mt7peT2jOxO6kGBVEDYSMt6t73w
uE4owuGOnozqM18/onAMAKOelVEqmcM1H39ve03k6uuTQINjh280EcHflWF3cTNw8LlrCml48A+t
BFXgoyfIgPeUV+aS01/WhTllCbXqOEUWumzt0ZD6hZNM6ESWDG+kPaME7Rf2tUPLvSzM6kFjTEjt
gaVA65qCmj3aq2sWz19Nwo/+zoXmMhaHwI1Ng4J4Gy+isr7hwrTwB0SGfXWwCfK2t3MAE39GUU/W
apCLPpGKHWVabHEu54zuRZrG6qpB94DKB/nRqpTttN64wnjq8dgBeGVW/B3cl2rzH0/STW1699Zt
pBPdvPyobBmkWIv2k2QXSxOhIv445jpb2KwjGc/mSndOip15ZwCxc1A2PpG4mVBNVyP6lUY/PoAH
SzxINHXtouqJUVmU3oRXeVTPru+Pk6D8EiP11BsEMX+l0IGUy0XwLkva56aEnzYl1vyBfO0OgarF
Phk9XViq92mq9JJ+EivekVFBF4aoWqorLsAaTLxLUcESAw4agrsIJeqIDB9DKenjPCcjEj4ul0wU
fNpbvQbNwefQfC8MwQrdEunT4ZWscy1GGYkQCglRxGnkvXNFJsqKduIFAWa9WMXufeSntoTFUPQH
jhKiuQ053PVVl6n5G+5r+mQ3AFYWfqNueg6+cW7roeTgxwWPjfps9g3TbXc+OFlE1MRICW30h44B
G+jzv4Nr1K1n5t+c2f6yx+YbxAXP8AbgNaKpW7QlvbIktf+ooOhGJUeKIAIoPy6aKghMA/FVpTPQ
/YcptrXOt6ygomWEyyqFx93wccrVnjmYFunSZiC1+IqFiBY09HJ92ENquF8VsmtkjTKXEDMSOT5T
sNBQa+5HgJNjcuz/TG8VllPd4W22Q+dycH+6xnMhvQqmjXeagGSJQjz4/T9RdO/CaavvW/WBxstW
e4ezsraaV0TxuJieJI0mnqThXUVfn3r+TaOe9LD9qCD3H+C4KlaUkkMJVnaYPQO2td8BdDwMGT56
kZXAe0l2rfrM9g52GFFZe11BdFWWlDmxQO/b1wANdJZjbBMT4UCg2M6T16rGuXGyTvVVqmhSm990
oCTESG1mwNqbouXDghIFl9LQJnbMn1cMlP4yscjaHSj0V2rMlf6YlLT5kfUNRAhGqKC53VrYC4lS
oIwRjfs56TiTygB/cm6meRFgcaLhl2BPXAXIEYjU5n8Xm1E1iTOw4q8Lx0iPj3OU9UEDVda9NxDR
3qmhzgu2/XrFxqhYmeKn/eGwAtXTz6sbQnzHdklcpKtls9ABP84+hJwLA2c5jnHYfEYxs1Cb4Aeh
Y0aqFc6zbWjvxjWSDUTMWK6tby4mHNvSli0PnAaomd0LCCq1uAp9gPDlFyU7yYSmAjHH0ERkrs1m
t4GCbT8C6CwfKcSgv2JMLjpOk8q/0EYDKNjDNS4gE2WcWLUkjnfExf+51OoAV2NWdciEmVBjToVV
v2xpfkgFGqjgiWNaFqAu7R93kgZbZTJbxv23bbUkOy7WBfmumj39LKd6XA4D2C/4qAHrBa5CoJYL
Y6zqPnfdWxps+tsTWXqDfWhcGVor6fcb8pDnbafm7DHUW/L975CowS0uBQc/3GA9T2dZYtHfKYCz
73xUT29GSDwBZdKso3WPjKGnoAJH83fLonMQx2uBqzx4nnOuu9Icc0+TEgs4znAuWZQB+m1T/vX9
qdoKZNHvfLq5dkcIdp3EBtlAkalOHMkBN9BPRm31yWscrc53jqYrPTnrJI1bfMr8Y1X1p7befXwv
0fQ6xOHx0W4uqLB5aEBhDjzVtMOKAQqRFJRm5niV1evadPyO8CiOnftXoTZ7kcF7fpZbEWJrxwd3
RcTRYPrTVKAMgQdzZwUnBgM4zZxNGSjDJPFOPylLL15I0/q7IC2WshFevbgQFyrp54dJ77ZWe+MF
3voR7uftAmtYZyb/kJYI6t25jutjW801j5lAYpXUonjObTNOdeNCCFMEzZgjlelLKiu8AomYAlYL
TQeUBL93gf2RIymJUb95C+xmhie/7/K19GhH90KVmRkm/3K+iRCx16zpNLHLCAWb2hYM3O2oLp9Z
grL2jS6RwKYnJGgD8aCZ+Xx5SX0mA7xcIKwOh/DdHcSs7Z8PEE/7bH2i/CoedsBB9qBwS6+xW528
cvpLdfgV7Jno+8+yHPzcQe/HUdbV5SeunBExjXWYzBu19AEv7lGc+1OEhxvAxoCXJ5+crHWf4osF
yCsehhQwAZJZup/QNDTKg2KNSg6DjOOj74QYRIH6RlNEHnQFDnzYPClJHIw05KYG/dtIc1QNG6b6
j9mL45e298zga1kXyTPA+kS0FePstzHhCI4aJKXEf+KhhRlJB+WkL/jKj6dqba6z2zSEhYoYfOgi
4OifCLXitQJt0J9u96ba2K1l5bk2jOsQ9BDouq4x+8DO7jPJLwyOelljPyRBPJRBtpd798COHpGV
qCN7/JkxQX4c0ZwXVfHtb3bSPq5EC8/pokWuPvghEDslArFP/VWxhU/OYxwlGfx0vv+y04eZf2K9
ZufQEaWE9KeWwiB8iE0lSJncAeUGmVdtUZr6LghAlj/YbnibOECjnf4J2pYohRB+4X/xMJnt0qgU
QTKN6kLxTCUpcR+o+FJ1cwWFtnERntRZOj+DkyXYYH5Bh/nCzG8Pwgsmj4uWgzDm+F9t7klih4TP
GKSw3kpKQV4n+X9VschLfFvSMq5DZXNw4lir/TYES3vg8p6Uqw4OyU9n4Hv1rmo5K8taqbFDEttv
coqB8hg7SOdBFfWTIqRj9vWNFfJYTbUrrg05xNhclqBCzi5GdXuPI1Hx2angVUC9qm9LhrkUZIhD
SGmuKs5WlkyykxBKlUXhg0RMsw4oePTkkERFfzrCF6mTlszOcqOQowds1MEULIztK+1FBG0ZSqtr
mkV8ROcgzX1yaeehA0M+hQT6bKI+0mngfQ50VyO6nlG/2taIahaGm2KsSJO89FYKKBRiThNYc+6u
1/fpTmWRX0HZrWeSZ6A3h+riMzohtqAqpCXFfBXI9bmgUUtYVfiuzynI3/JnH9kh/Hnd3v2BimKS
bxb2wH/vZ0gXFjbt325c9+dSuAFaqMZJm3W9wNpVX45f3aGCzKzH43V7GmLaoAW8HzDzXvnrOpIB
4VlM+GunqZE0jpu5Vz+VU5XtWxCQKXUeTH1JwOZauKIoplxBNgMp4VdMsnhQNuZ8gbU7nNPEDQdi
2L1plFN+6iwQEyhvtjmakQM/IfdYPyBAchHFPU0Xw5GT+R/jyLZJS8S6h9q2vr4C7jSF7QL4a1J7
zzO/9tcVRtvughQekRPfAdqeJbbYiLwnX+ZpUJwkSyyzpQ/4Ed40m+4hOSFE5YlUNWokJMufUY7K
kdkMMbZHbbCROWEg4dUIyYYvI5lXYrfBbmJA3kE+YVsoVeWnIUu1gxp6C6Ke9uzE7R+182QkRqDR
7CTHc9lEwppA1joOT9HY0m/RohXfT1FKEVJ5QiY5n68FP+BLQzo7bDV1YWwa/BgZLtHd7ELJ4lEd
6QnMSYE/fuNBPmFkwiRftiAU7c11XiyMB7bbtGJabLKOgzLUbvSGXKFe0RWVxyphC0AoTtZjjiUB
yWNDlbqjrFl86P30PpYlHPw5f0NlSBSphekOf/1g7lomAyzCz9mIYoEFP+noS72FOkQT1I6JbQfF
3nf2w785IydK1LI/bscHwsBMeFCCnvt61ZuiQ3lif9hyNBppfptUusEvDrQ4kfsF7PnxWpYNjMsu
wD3dgsi38BNIMaQUz7r4mWB7pdmuBKRvLMM8oBRhWaoby/0MJ5VhTltsLaZ/LpxONrV4/Y1jLWkH
yXuL95U9Rh5rgjL8GHXhOL7/Ft03m8vBjkQgxuJTcbtQoJCH5i0HdAELLvH11JqHAv1LdefF9nws
5Afds8QLtZPOg64GtFtquixGHtkdWK2AW5csnq+eazleusIKPbBahji+15D/JfVH9Uf6pTvOmZ5h
4xWEN/zaN9ruKj82JbRnwoF1vON/FruwJ0fHT3EZwrrtwZ4s/tEDUVh7lXgqHILCgfc+WCGIKWG6
Uy1HKIk74E825ehpcdK3wrfJAFGHsuejMc0dJYLWctn6NcK1wnJJQfWi5fk3cgTi0JhKX6IOtgiT
8jrUfo0yX6Pfd7l8YvTiwp9Y8qhKx/fHQDIIesOA4sp9H4moojGNlzTdt3eY7TMbVRTg0KrRoJvQ
5wxGh8WP/6XFVUbR3XLgPf9ue0vISJenulgtKfKig9sJxnqlXUXXtVwUEifpx9tMwcK+w40Tqk5m
2a7W+ngtKrpC6a19xyrg9l6LuX81M7GZxtNPrkglgVf9Taw6opr2oSePgsi5DY4BhrrPU2ioB2mG
nr9df/CxwmLYyZEfWP8k2wcksSS1X7lzjiHB2XcQp8XRoI6xBX634fBCpDXe0KHOLFukWkT0WPJG
FybQTI5A+mfEdTw2V3kl+91l7cZoRFdhGTU5S1M7siqEtNyJmUkzHtF9K4qE/4wgSQOyMhCjl+5j
g9GPnWA7tIXburThfYizrS6GHVrQO0/79s/9cgQl1PMtuPqihALO5yqeNeodIhzAS0V9pYfp9bXJ
3mCJiylUGQ0CGbXBPVDLppCmE7ZbIxg33uBojtB0NjbxA2HWJOM+LjQqmSQxXFu4VUl2SGQv4yHi
k/Clqf86Iyh6xXYSqkQu/Tpu8qmgMkLesqFZ+lA5rMHbKqXTsFR8ER2Tu0jbtjoHwMjiL9jtr1nB
1a5vnzOmmAtszbNx30LN3g1XihiwGiOZnVs9SCxg9sIOwKbIhL5m4EY1KrqGiUJxqUJMfl3TCFju
z0WqYNi+HLmp+5y9ShsSzWJw90O9DYKkISEUyk25ya/G30t/28em1uWuuVKiz69FW7jdH02aeoHT
iU1y5nLxDSYZ2pRlNf7U7WCuZvB93wI1P4uP9yFJXRykIHuv+APG5Fc3oh/45zG2XBarWF+T/pvY
/XbF3fTB8T9ewj4PK42C07lheQXL1M6IisqZ2AbT/darrBy8YAyAOC946d5qvOndH07ZWmvw3UKw
dwYyf7fGozAdaFMbU4zgUB+ruGFhmBABuJXcJQn5cpfS438bSbSBkT4uyfq98Kef1cNDmqvP9BUL
yRz2MzKPcQUp4kwKX4PkfIGPbbGrsdGwNDonXPMc3yGGKzHZY/p9mcCABbX9ljtmQvt386EER5Z0
lDxbVmgg7zn2MPiss+adPdrwDZyoNP5AMOxbviimcieyzzWPJAO2X6fTBpOIz768yly1yZ+jOKSS
2w4dJoYiiLpBdduRz62YwTAHQvgzF2p42ALNDQA8UaUIVRjxuOJDSRM65PH8wD0b1PWkgm+R5ZSL
JOwzwaapRbIyvPxCt/WdgdXrnfAqzc6IlxOkTCx+Re6OpelTDre6ULsFMIuC6WOIJsvjbk/Mck7Z
5O2KHCpMx+Pv1lROWWx9X+jgwv+5dk12I33AR2INjkQVgCq+KaAJUJGKSmJz8FNRE2SzY2yZZvXw
g/Llh8farx8Eei0eKPzXJ2sCnPUV+ra98Z2bCfsZ7Qp9ZcXofKc6dAvF/V9YHTBbNvJjnLMzKGDm
fq2uIKWqS9pUtt026VS++9JfdwHJURsfG4AhfFw5AILpnJ5mskixD+PzsdflCcBoqumZ6KjjxMJD
CmnfHB9MD7cZHJYtvd+RSIe2Rp13TKrCS080DLWwqVLP3EAKPLi3zCj+nS3QD+cHF7F/s8BY9EXd
haam1eL7AA+nJDs3gyF/2tQyqo7ryIjOGsVoMs5OK8GVNe2GoO0472T7MXPHAtU2DMzThvtQjQuJ
WaeZhOC+HGBXDluUYSrWmGtTxhsPHXhhYqIM4UCzpN+MOZjbR/eP8xTbM2lPkM1rN3gY9TWcJeJA
TiC2KpBHwvK897RVsOaj51X7YEbd5vjUe65lTBezCs/oh+1B9nxc7kuuW9KQ64juCfODWc1rIt2S
TNxnjqVVQjQfmawQGXfISxVI0hQdskt4htCZQrDgqOxl6qsKMWiWavJLxQ7rtKcerYnkbVSdsVPf
sP1lNoIc0U8N9m4O+yT1nsMrza3g1tBpKAz48YtWwkmKGGEhmhp/na6C4jujtjQG9mJpDlRegk0V
ZfTdVyMMa9jr5ZpliRbMTbR+esWO4geZCJmKBF6141pLPTbcFZNB1VNWKmUU5xZ9Uq0c7xZDyibW
VIXnZJ4QagODzLXbTPY8GAqQhWC1IF+CkIVHNr/e0mcG4vFsNEx/GctBIDGM8TyKdXHc7grQSfaP
SQtk81+OZOaqWNH7K0FQ2Qf5bmz3SDKVsjHk1FxEFVFsqF6VKxU3YRmGO2IFyLFqI2zpIuaSve63
dN8n2X2bmgrgtAH8tZFHCnnICRH6YyZ5ij+iDdfCVbh3hjMhBmFIq2zFJhYV+CwSptZI3oEVz9+F
rw+uhtUWU6VVyVnNwB4IFFdczMSFwvpauxbgWnM6VWtVz3T1aMYVGvLBCAkt8lehwsJlqd641RW1
EjTvTAR6fYGxm+VxU3uG88y6zC6kApCYDEgKRMeuX2F4I4s0oCxiMgGrcA4h0NcQ5ayr2Vy/F2y0
rPH5n6B5GKPt9aQcFvTjtv9la380GibI8yG80BBcOf66QRJQC4gmnSRdMoN6Ah7SamgvdRmXKucP
U+7+B/TAMHQBRSzWOw1Q368g9R7VkKaiUPKxTCyu3vbEGYS36k4rWWv2NHUr4IDWYr5K2tZugRxs
GmM7D/3MeNo1Q7uqnJ0wtloeshBSDMHG4XYEVwGq+PlKub5teSPMG+IrNrkXj8JQ5CZTXywKvZwd
UhmSP3SuuXSJz7FN61e15eA9kVArwFsA9lHD1lgvtV9Iym7y2jSiXwmdC0Wql/K9fANx320jC2OE
yzA71d86qP9hvEsvQY6Mo4oa3Z1IAuTMydSKHrT0IXaHvMWha8faoyAyP2bMMKEXwJJW1BnN0anf
GgUaZcFkW8Uuh+yXZLpA6NoGI5GJbhxXxk3cubwrWqs8FcK9n7g1JZELPTfPs1dKef9KpAedf5UO
e8uEXn0zy8oT5G3Re/vsI96Mtliy6Z/yKKUkoFsuTuMq5oCXqEbbGr93tclhZ+Q8bpdfiJWFo++h
W0AgVu1T03PJQ8BZQjT0NnLMnWdrCCzATD+CBY7sDdO5HeA6eGaVBE5zuwz6CIqOFk7FF18c3sNO
RAXZ3Rnx0CwSc/AO+TiBkv7DAY5YmMENUvp/QLUqwQ2QntKZuHLrqB3q9lKfMecWgWbXeEYfpjKy
ojBKjU5x6y6/V6l63I2j3biqke+JgfvrLnCIDLCV7Fte3GNFwjFY3UsL21FlambLsUMKOGelY4Rs
vi+HyLnfBDx4shnHVlyxrxf05W88y+BEic1JVfxx+2VtRHyealByPOgN8CFwD3rphsCEozDnFB/Z
XLTCsVp2BA+XmhitGRE6/cuoeQ/izAwNFLx6xMTOJnjPU6BvsHX9EiFEaeSjQ+AmAAsDEVFNtPAG
g8PXmwR/AGkw6o10pI+kOixioGpv1YONepKl5NTIoON2+dYi4WhwU9XXpqZMx0+lSdeGh/ULkJxk
64Bd8+EfXNwYbbLZtYoVa7g7UO74C2RKX0H9Bk3d7Km8RmG8O461RTeWMwwvTzCkdCFQ09mastO3
jnbEedpddlh6i5zFOHtylgcqhsWW12TtM6S54MtKYUHyFv32MDcGoleSi/hVuOW+moxRaxo9YslB
XLv10au1MyUPfWK1RhFWXA/gZoBiEw1nATeUTLDGflgxe+C+as6+0yl/WtHuO7lDiurPND39Xsbe
9g6LJvjJN9le1FP8BzxCWpMTxrqWAqYFX6GZKmUKIfI2g0/x3OaAdqf1KHSDmTi7CA/kbo5CTmn2
jDIeD5Gx5yl/KjdJ5KZUtSN9Lzw5l0kwTw3SSiZeqv0v60flimzXbLGkxGBKNFmzm2YetvOQbvQG
zZgRVlaQDvd6Cq8/TxYQCUKc+B60c6HPWCNfKyRWqlSzc1w/B9GEJuHqk+3FgwUfc9VJahIkO7HA
kDjBm24zXplhyTJLbr+5L+k06arPY1Grlej/QDq9GGbSkx/E16LKZDl3/gO0b7sJRn8E6pkdNqVG
GTEKwHY7h6PQad3+ki/QeEIpsQ6ZphnDUypy0nD6RxpfGl/MIBTh/ZWkftY4AjMKeGGj/ufLgfkK
AnPdNIDmRjVLTttnlTMvi7MX20lR2+Y2rM90mrzgUpPBLaDBkZiDJXIEcK3+uWA3vsMTBSOwuTeS
5vxOojR5i8LLEm6ToLt7Te1wpVrfcFkEMDPC1ocKt+h2a1UsJDYnl46toHkzl2/fdDqK8G2+jZ3Q
PxO4pZP/ad9VDc8E78Q9WDYxSHLgLjxEfiewgPY1SA6E9uufC0RmrkI/7mi098+lZ5gHg2O8//W2
ImcP/+Ym+p4714tAeifRGcBhYOnNa5OOoop+XH/KlWoJel+Fo8krTvpcmqpDWgFwr6mxsJO1sdpH
HTSg72z2P4f8YS0afwsw10KwIMQ+KznLDyYQ4S6XNdWrvU3x8nWxiSjfdYL0UvAEv6bnH8I5SfoA
3Q4PkiUHPHS1qpK8LLPWYzLGQByvaZ2AHtfPRRhhDBWeWH5B9bAdwvcVYwFWaiigngfUjH/zER/O
G2smL7pPUr0bzzgUY7cknDnMyyCiU6b3X6cNA/L7H3l7oxm3mcvb7UdSIerqiLsJWv4m5pIP4gMj
jSFqZRy6rFx6dc7MYnK+BZMTIWInTBNtEvJhhBykLQ6hgw4zZXgyad1PVcQtNsk6u1b5CKTRHgk9
1MvoFUJUKp1vSaWazpKvTcX0sTSEY9bQoYeNjhb7cOE5PGV5exDbN6tKl1D+0zuU1ZQdh3QX23AR
r/sLoQ/EQfjIGk3HLXfnQFGjBBRgJHsi6daiTbg7jZ5sfO3Buw83NHZlv7Y/xuPsIqC/AQFUq7ZO
vGiC7RzpSeavCOkzfe8+/92WX1JyoEQkuZ6Bxq3703dsmzQwqEqS9Tk9rkM5mjyB0vLzi2k9eeUW
5q46+92NHX2Dp3asTOz8LJPyLAHxfIjlECLO/Q9rZxCiuobN4QIWGGHcXXcvGtMjIXioKI8eeDNE
vIOotvoe7ceouYe8cE584RGsA+uau7TQUYU2LPiPUdWBSzKwycjjkfL6gckuU1eaMG/yW1mYSK2L
HdVej7PqyMgSd5LLHODeekXYRxCcu1ES5YtDhIqPN7cybO/ciiK1fYVipRd/dFF/zYTvW3xsrzut
/EGUbEACdKJHhz7eRnPYa2xtyu6hBAV9neEu/1KZmOBVgPG9xIxIcxbgfwOgodG/M964PZTcN2kO
mO0lKtOK1YTxZcyOV1vTP+Uz0/QcDujOmIJnw0Cj6jw2wdzxsqiNvsXWnIGYC+zB9HlheKsD03qf
AY9S9Ko5XD9TN0fYRfwx6ggDoadrFY3U91R4c8J/0n4/YZGvwFn+0vmkxAinY1ShO8KDemYIl+ao
eAF/+vv2FZreDQCOh5pjwiiuRS1TCFjUk3p7kssYdvwXBvhtirD6CseUR+2tbGumVMrxwHUx8k+4
Q7CwevF20XBhPXweKncUAi6qrkA4Gw/XMfFOZi//3K/EaEoDsZZ2ZsfNE4SnuIJGcItwBsmG2OnZ
JtRiX3ulcy2sZMkmoHQf6dty+/sUr9hqqpWKr8d3F9oYazF3P6VRDC6bdwEkpwEGykza5s48mfM1
sYLYoLN30qZJ6r2iD47438L7cRktVH8vnmyi6IoFtmNdKzjRv+sL2nJyr/bMW1cu4NTfdyU91sYo
8ZaTIKNE39EukuDFbhupE1xrL+kBhL9Xk6AxxPGd8/njK+M1G8XjY1WlUtrM/Qc9CCRbesBQD0iL
xNtnTKMpRMDdsxIHolV0TQcNZcyyfYksCgEsfGElK4yTgtaGLfVl9m1pSgCGj7rsWIG+tBvLhizg
s0T9Smewtp+6Wunesnt3rnoBiArAp0XafAzZFF8gKgTde7MBMrkDES5M4YPykRMZxmkxqNY4Q+iK
iR2BQNBhb9cfzaVuvs23DJaUqh5w3IibE6uRahtAbT5uZJi6jUe1Wk/5GRExujHCkHNSpZTv2krR
YYHmXpLBG6sXcQ69axyYzbYE9RdfaGUXdNAmkiB+kwcnWa+C4YxMdTB2X8sufg7Az6bQU2QAEp7q
H1FaJ6TVxoLH8vxutGd27Mev7/+vlnaQ56GbkhIHX9nL3rAs1XkqN2tCNEwUqLj1f44uBX4Xjr1x
NhZcYh9P3pEwZ47ngBD8ofsYUUcYKmXhVJke09P3qgHn3vMpR3R4bpdBJVcEaIEK73f4R1XC8dJ5
+LaKWJwvPH/012QSmrOjW35Cm6wQ1ur3VkhIPhzjQMH0gou0az7X9LRFuI+TfcGqEU6AhdlQM7ry
ZXfHzoP5HQOYiZe1zhTaVClH/FYJmcPGAJ7YFU7AT9W/FBlZ1ONw6ziAoqBpUkqdeQ46tJDCJXcM
qHgDYpqHbdgvMPBubIs0sTN+BdTugc2Gx/oqqrImPYNXMUJOPnPyiHZlBxl3AS84oPV3RoClwTAO
NY8VppNMS1PcAa8KjXb8B5cULFw4uKX9kz+vknpYFGKafZaMfzF2Q3xEWZti22nduLtRhtGLqZ05
DEiLuayacV7cvanb6JbEZrxrCuYGoartzS6aOciBCL+rio6k+De+fc7gQ3dejMDuYOfiN22BkYAB
dnN+RhKCfhkZZcSNbU9+54ufDFB7mV3cGusYEj/FQtH5lJLmxJ2vRoyasuZCgU7uy2M/R3BEmMbz
AzAxwU+jFhl924Y0dhpFedou+sMvAHO5TqJwLdXWbVoe3zbA8Mfigm8ypZZsKX2tf2fiVo34x08t
wPjMGBfnxVGXrTls4stkfSAF8OUIjgSR6tZJoVizNrgJ5RbrsuM3eUsaOgCN2v9ohYKhjVk3WK02
UDJloEIlkZzxyiHjXzZ4eRgMMngTUdTE9+hARZ0LAUA8j7b0Y1RKx+al5rII3DyHI26onh9oivbT
odnOBuKW/mgbipjzs+Moqjf3E9oL/0vfEax0LfiNXvm4xAwGnxx6KlhGvSVkOtD4ZGEAQXyXVwnS
fq7zMlXXeIDQcns/2TH+C/PdZ0PpmFg1yWm+gmvl4fY+R7JoOHCpdyoaf8A/1LYp7MroNPKFGqeB
XggAOXArGg8ttodqcryhn9M75cuVa6Pk7TNP/5mvsdlUPerzbLSlwufg6o+fQBMZkd3+cobyVRpd
hmJ6eHRRiiCHUcUL3O9Rf9xyvSbakW/msqQdpcPyXNN9OowX9cOuw1/fdGUWamYSkIKo19w3VvrC
gqaCXW4eMOAxQ+q5YDR7NoJLtunDz63efGd45Bjyzs8rkCOtir7D5kHFv14JKHZ56h5Q/uSNE+oO
Kux3WNZpOI4BaEeL5dik+6rZ4KTaLBasoNIwSt1Wl9ide8Dr+bzc2QfotW393Ro2FKuo3XWoLmqM
9oKXzCeKtLWe4hjetAXDXTXmR5si/JugaT9RFcZtPxMzf1AAgwru7yqGAlHmHd4HvAu1bUkuMHJe
IgCh9IPQ/aVj9I/Hz8K+XILpR2weq2ETFSO0dMVRcYoUtnHv6jHZKGlSb0UhcmURDW7HExagSoNQ
wxKx3ThYgtlrCYnQ4dq1ummYMSIi84jVBRiCYNtCtBkAzL10d9HxL7c3rtJWu70t7bfgFhnOrPI7
7k9OIdEsa/1yCfnf1WCbLScRneSmxg6MOE2RE3R5HNOn53mK0vB0wTxMbhp45mZQY0mkrhF9AlFg
gHEqs/I59wzz88ZV0hfAjD/13UJdpktkP5f06IahtvUQ7Wku5LFQbrUL4v9dd649qJOR+bms5yTN
LyMCFFE2McZOfHIDuUdZ5eg2FdJcrnh1rRo2I4nmZFtBF09XuJQaZypwGU07j4o2MgL3/v35Cyfg
Iltos+1/AchkrjjrJYBMUXdEJmvmYMHRYxJWCcQMmj9Pu9kUTmeG7pGUIOLTvHn2709h+Uhabava
sI+RaF5YUonGukaNAc8L8O3RH8f3hck9MsAHlW5qG8Vz/mIT7AAL9Nk7SlZmr+fs/bUK2/nAhq0E
ZQYWHnjHpkTCQbDMQshJjLzpF4DLeQVkgWdk/ac6iO4Ov5rCD2xeTVjicuQ6jMfSiNoJwNKef7DR
EiJ7FCRrwGxew5wxzyT7iel5rGrDTmtzg4MkeMHPpsGiPGHspnPeRuu3KusXJbwef4ZxDa1A04zF
lAQiLHtFvj5mcJ+SeLiKqUzzQd33tfo/I8OHuI09YB7HpE/uLDYcQj/xLWm/hgL5MFFSaE7hkgy0
I4uZ/lLWW6Zi2Em7GlbsjdJD7Zg3PNPnOz7X/S2hSykerbC5jWL4Xr87Cyt8BT55OpRFO4kAyxiG
UdXVimCwJ5LUHwx/xtB+Ds7BbhHJeq17xv3a/Pxwz5fWosUlnKh6sjYTd1NGrEyFtmgk1CUvWB4g
2DyV48YKcnPGcmHHDPUwG47LgQLDXEf4ancKOJ4+v5zRYPqkVfwEORCSLu1SOMLJfWDaqEGBOtt3
VxPj542z/MNs5QGo5+N3GncMDYEHJVT+kj8jfLF43zGrqFMS2lXs7icCaqnRIGY1RR1l+YHAp3wx
P1CpNMkWGtDxkoVoDWFEyjhxYUVPpEY0hZwA9r76Fjo1mWABPJDnUlVwyX3sdjMu05I3Ng/ZTbFm
HlSZua5PaNEss4ptSvI9o9MQVjw/aLr+GRORo5b9Yxgzs81y5+rxhAcTuxQQRwOREJLuP/80zELu
SsfX6AEt/gj8+Y5aDwMuJEuiZsGPUzamrEyU945rXa/0UKzEd4Tz45dH0tJ0n6cBYNoKJyg62n/p
9bpm/qo2HT7B7BAfULAEa1Bldzjl2oaGE8Z83iYIF9sStxe+IMFIokipKcfuVBI9B4adS8MH9bq/
X2bqIKWt1NbwoAOeJyYQpePKL0M/H9OCL8GRayCEjo0HT1WvnkNz3sNC1GcfjzW3Vrhpi5nNXxrC
hOaoQZsysFmbvyRlvpghfpde/qr4ZcrIPVUCl+rRs6pKx6xDT85ZXKjv0yfTUCveYdcOWpqzKMUV
DRMmDMteQua8hiqHCzc+KIF5k86bgmRCciwpXlcdf1sMQ5CvYT3wMvFyUvUJkmWjepSks8m2spRh
ijwvLQSAHwPXkePg7bGAVcIECaezValukmzMEYvGYe51jvggIeA6TPG/p+vF/R2h6oHhGvO18hrB
+NU6104U/MDfTLFnBcN/3mWcl1NjnVvyRU4IxBLFkrpqY0Ig0DxD1LI1a6zxNkNfhrFulwcO4pTj
VBIgbCSAqrnwQ4CzrcR9gpRmc50GoDxw0iNZbUHvus8Q+zX4/9Q/QfUhrpfJbTkLVzuzIUAcQctu
M4qj66OwpqoowR27U4JuvYP07FXMn8V7Htd7SOhC76PP09cyAWtZPnHURMdFKJTanD7Svp2pxTuC
zof8OOhmAUZeTXqw6XS7eN7JfmAmK9vASSqBFfmVMvFjguZ5LH1+RRlTzW3eg7tPgewSXJaiAgUZ
vXOBzHhcoRreRi8u9+JbzV1PZPF3kQ4gEFXfCLzYu9wi4pj9BDolMkjGQ3nhyWhC2ZhWrhvTazMt
n4elrj7HCFZLv3W51WQfuivPE8/8dkWJkcdjCU2T7Zv5XshkeitTjT+s+P0KcR5FVB1rMSogvHfU
1Z1WYCjf37GHjKw4BR8pPO4RkwxDSW79w4C66DfF0Yt8KKeipK9gmzATbZU3/duRLS+YCsAa6b0l
Rs0F4ADVZq5BDbBOaXr+3Jref0PcoT5T6lR1qszQa9j3afNzx/XH8FTKPx2cIWHgwrmIkVe3mrA9
Vgo5wco5OznNHYBpQ3Xy/CdrgM5hSXhoQzllWsW+zP9QpUZEa+0A3a8iS8qeNuP5CkBBdPk4j5W7
NolCtxnyojkPemm97TWxr4l4yGe06dG7xHNfPTc4r9AfCK/Sbhn8RCHRhQdKRwNACG8tpUyMy9as
DPuvhoUl2brQ9t9xguQby9v7fWcG0l4GpluWZVJ0XCVVq27xrDEDxFERBpO00loN8pSgNOyZ/pyg
pRpFIQ5ARMqtxkisbStT4mh+9pjDt5xkHqoQhtjU75P59p6DwhlXEnp2AYV4q/RLxUVQNeWizved
Ql6sESsiT/pHZXYIxRQ+c5BX0/Ppl2hgl7TOTNI9uWMqUbtDrWtRDc9/FuzPQtZB6DrovBcvS2cV
0EdNnfcwYjNrRItzlRzkX55DRrbSIRvAsM8d2LF0u4Zy4IuJkjdavhExQY6igmEMfWrV1ntmldrv
2H4y1+CLkBCA8LSTzrby0IkEJlq8lJXcZUcFvEIKQ7r7SPu6sOh1t81a0+mC8Lg9NoRBCz7U6Tcv
L3v3feTIExCPykzNFVGncYhLqEzA5GLD9MzwabrjGPfw46Eb+/6UF3m1kpvPm3Od6YVr2DzrTZqi
nEeO5mCLUM3vcs09B+UlZeQC+KA+nRbWh3+3BQQddxzE0ibBMk1XKJTGN7JDk/UuG6vePfieh+QQ
l+dyEL1TwLfEOcO+StNhv2MZewyapmFre1OJ/8Rod8rRgQXv3Rj800PJvOEMfV1UcKfb7VWHDruI
l2PaAtQEdYHSFKfG4LmlZ7gHPr8ReqrvHLMn4ZOq3AtoLfd29RAbqG8rxC4K3jrAo/QI8pVPeBRd
qtrfR6xBoMvYK3lK4a6SUHbrCgzvCpN+vHUvW1OJdiRPYSwGmLnhEI5Nh5pc/775CA8+YlSOMmrv
t+sC9IIgkXacrcpYeYCYtcEcw00DlQcolKmNdNvD62Jt8H1QHk58xgShJ78W85TDA/LuuaojAGiO
soafhQuYkq0chR4f3GXovPPXs/Q/PugWXtxW/LqVg2DFFsl5WX51sqy8sdSIr8hurXH5ZMQgw/l1
zcLnM0V4eQH/iX4Oy1UOwG+yNiQQTTmBh8GF/bD9GYon9J4pW8AUwqkqYgMHE+Y02v4qLT7waq67
xk2q8p1PDovdQqHkMFribvoBPodCSKXTVqMkgV20RE7DCW9z9+fYkHrnslWq57r9nG3mbo1WE94Y
4rpM046IPvjAUVkV1TcKQJQDBBzP3L7IulkS1b54bYaA90OzAvyaj8pZ/egX3AEtEObTRjhngxSG
f2z1HddvbiBT85yui87+ZJzBKWDzH3UbCcaBPRB4TFOChM4dSX/EC1Hib3YSCZZWgZMWd+FV+P+a
iq4ZDU6s2GO2tnvAiRsm//R/8xzO023S31qsqxswDL1uiRpTmi48ufPT919qAK+zLbayN4Qi+U3p
R/3R2bIohXnvPTUVgcNgUoHRaa8ThR8AW4TbhGXKEezM3FcQJyHB3n8ryeU7QLd1OZwEwB2Ip0cD
TO3fRwsRUP5QtB92AjrM3ldRedz/xfVaHFQS3qj7r9IsRGrH//AqcMUGxPlRoG9G6nQbDTFSAHMi
8JRqT9UTOWMfYaBZ+ABX/SXV9aRh8AQI1DhhsldZR2TyqNm+uA2WMy9/WI1Ta28lNlsrhCtFZUPw
xpf5rJtWbQxHyyYN5iAlWKpQYuXp7oMnL2yvM0S2cAV+Rax+/ACaspAEoFUG3cVXvVQbKsp88GLj
eHiFsVqvy57b5PXXHlMR/SrY1HnUxEbaM8SOhzSAUoPjN0vO9Of8+wB+t8C2Eococ/LdqlRnEjnb
iF6uqo5Z0up+idoXTh5CcVfqToihAnsyKwudo9WTwlNUf3/x41tCpTG4VjAhuTwL7SjV+YJ7CRWG
AVUl8JxrsatXNrCIyQV3OaG7MCDHMrA64MqLaYyYvev5SHWKHvuN5QPI1wKlq32R/8QKKlsF+P1w
usIY+TmugwY9RN3OZMedrhQtViUXlFjRjlQan57q1eEHIGlWQ6yS8DHGt/3M6DVjpsnYmVkLNz8m
aq9UE5c6tJd7ZXFhG2GFr0zlVhg6ngz4Dq070zs7b0O2UWWneW0S0f4eFN1tjgJQcLyOHfLEmxSk
wBV9+X5QneYRN3F1sNwW8QEFSdjJhREN13oU1c5iYG1inU8yUTLWURfQ9a7psLWTs7smgqt/XhaO
SGa1sXeibwceOOmIXthggRI8z/PpIdjD5L+AK2cO96XK1ObvcoQ5CPqMw6kEvu2XBhiq1wQH++ba
LhTRvY6HmgHv3OaeDvJTdQTyHVV/YJwbJrk8m6+4DpefIFk4Y/nuVFXCTpGhPKbvUSGiQta0Jzcw
q5Gm4ElcfykupnT5yb77bSc1VCIn8QX/U7vTu1K5k9M755VdBVB9RuyJCVyl/9nrTvRC4OmdX+Vn
FbHRfoJOn1ZE4AdhnfZmkG6y6PfI8owD7RGWsE0JE7bFJ+bqOoLiRTaWoon5nl+J5XwRlrtriGSr
AEbmfbk0RUo6oh8xdIKjecdJIrMRQ6QfRQfKEgKvv+aZyTLM38Ibf5LO2T8JbvzxI5eJCPfHUuJ3
5I6fdZP5PDasiyvEscBLqyxVOAqIoBXUtjPy+o1ZT5ZWdXgiSs34jByeJlUQgCJofM0t7OO4RL0f
WR5ZM/kctgy44aCaupt7zuxLGVaVnhVLkaniqjrj3gsVzdtpW5kuP0r97aisRQIoi5vkKpc3t3dk
HN8agXyRg7CA759xebP3955mHeiIBL0unVTSVhJFVwxuc5V0s9wS0XjTicFANqb9vC+w6RZ6Dzmi
Uc4AQ2SDLhkO8qncfDYq4ap3COb2pZ5CYC81NIOFgy50esnYL7xKBsySoxA+3VM7yb/H9sY+YBJh
tqEx/UPwpndWQiPwy2+DTOqNHHW6ujiuI8cwHT3bWpKo+G5RoVPcbzwlVQPE6HV+D1YexX/JeqkF
WUeVFsx6bklXSxVBSm4cMx/AiDVq3E+5n0QiKbBOTw/fw0vNlH3B+XvHFZc6QEpH4ALGIqXsZ91z
27G0TEWdjFU9fNqDN7Q9JFPZGt5e7aLVlgIoQkpNLCX/yfPkLzsuOTrWDtwIRGl3ryIvlzFMVAnk
1rZEk9/d6zfmN46A1YiSGtlTFyGsYXg4nXQaG5Tan6RZdXT9H0bh/YBhNOp2a1vdfyghgh/kbvQj
XqwKjT5ZJ80rDUXambq7J9d7QPIIJvZyaWXTOcRqx90QS2A6y8Rh4QTX/VEHZqY3yNCsOheCevjs
8MuucUIKoZ6LhvqXUsBZGsyJCYyXACTb9ZSIuUTvb5ztnrbRzjatnfeeLl+MG+MyUgrfCu2dXNMT
ULCrmgmBVNhHMNcxdfWJH+CoudDgLHKMeNtOKP+o/vbq7HM4v7hwB1lsi+6PnVLmM8yUTNfkvQCG
RvdittbnqZXpz365DAIf+hn0F5E0NAvjW82yNgKNDwbgEIKttlsyg+5alPhLcMyZA1moTMskD7k6
21dfgC0we7Y1mMomyRaYK9IFLGMsEjnQokgWGhNs29FIUytTgZ12W9uaW6IhnKJecQjqfktKzs5g
V3MheaU11oWUhub3SDkAeqZu6GHc3ebffplr/9fUugn02zSL+qy5tdSsIP3iHDrJoZYR4WJgOi9B
Dmi+tLxpllaOg1jQwTSW3Xl73xgbFGP+8u932Qol8BRjtqHgaO9XrA0V8IANdkZjJHLrj7a3bRVk
A9hPz0WGYLXdqLNwKNlmjKdaVqLvNAZIpFHnZzqX3IUZPkThIMCE/Wz1HnLI68I45WGdPbuya/rx
3XN1lDMQgZmLY2Kj1ujgRD+0+B6e/boLW5nQIEUSaBiBxn0DZ2TPMSklR4sOrWLiOYRUdCU015VX
Au3vV829roXtHe+sDbhxJbK0BmBXOk8h3Ts/ftdg0MyvFuUbeNH/khEE/PJYLinwUVHpbZP8huFt
V7t/OAQhE+QlYmvI/agZdxkrEht/oNOFoq6yVxgxVFKKC9GIgPQjjyfFbDyi36zQp/gc1kgTPxFM
FbZ4mQqkEsyfj+fSSiUfxAc1ovVBqyU3L6NeFE4dpkTOAVLHF1U2KpbxJ7aRbZFOJDks0IILR5Zb
GARvZ0xJGpI8mDvWFlOsUwHUe8/qGnwRx2UdTHcin+M3eUfgNmCsNLOGolbMz1KbfNlYwxq2yqKd
J9YMZxTuuQCr3/Nwu7iWgvQYifNhPxwSp1YCSMmEm1JVeI0B9uhhgim3z2qqNyev6g0QH+sCn5sP
fqm4Jw0SwL/l7hA2Thmxp1mMoe9l6ff1lKyBnqtWZJ2g5XyefoEefmDtgdqYP5s0xe/cM9TDcJuX
7VQzJ84DE8RLKksme0FLn7WYA2EwYS1lOll2Vnrm5PPYd+HgJF1upNy5Ar/zwf70wWUGWap4oMEO
WIBEVXZ5IekBnhZc4XW3/bsxqX9z/WYsjSp0YbbpaoOXMzBt4r0BFzoyCNGYo+VGz2ug7+F3ERCr
L/rgmpn17ucsG0iXS3lGeVmwQ+0qequj84VRLbG3mqAoAKkdPCj81yN5nWdpUDhdJVcssAwXbHw9
TPbRmtXk3f4OCPWijaB+OLnui6Yw86ZOHEgXgG4wjb10QVmF3M0zsnrOFnP8WwoK3CgvHlu3dQMu
SxzSmDyHL1CvHopotTKfXbknm3D/AhsDcTVJik9szDX6/cVhmXKBu7CL/Ktf3SaNE65y/NIUKGbY
ldVpQyzRO/u8EudH/T+TaPoOa5nPedW4eCaEvQr1GCglwYD7QSt8Kl/KbsMkh+7MzD0f50Amjrsh
PVWDoNVROOr0gIVQDH/mrikLx4NC3UzbKUnwRL7i30ITTJxiFMwXLqwKjBa7jEU+gCNvZ5bZuk/j
nsfzW9QqZ75AvkhA6AjAfGY+J0+qidUZPV4YUAWnZt2BP9SfJfmCocTvCWDNdUB75KzI75xYspKC
rHPA5pwlKWyG8tpYk3P5hI5IRw7f6vkwBICtxuZkPcOYPkMBmINjvYt+1Jh/UUfIcS/qcRFqjMkW
2Mne9H13S0hdmnyl7OFiUtQPs92v2yjYyVm+dY/Fys9os24X7XG4sfbI4P7wgooC5uQg96BWdAuz
YpiRJhmRaJ06G5DGjyG0DMu6t2nsv7r1f9WSTLgR9hBDXJFncDHpKJRlH9NL3orN5X+EgKdJktu+
SVLEAvD0f0MaQUEGYBQsWhedBV3XzjUx9Bg0GRazDPIgvO6o3KmBwbssV8Z4ilBxKZB3nHaZjP67
p8E4bKttwzRLxVMOnyDqmRsKE41CVYADRVPE707Mt+CqLs/afLq5fwJsoCZNP5NSyDFrOmhk2DrP
IHG2RFqK3CbqBP3rbD4bTXORoYH/Lqtc9Uf30SGSLuJxVCOt6zNdUSB7DiYX/jBF253UIXEzjYkE
9ryCgftSe35pjtbhwUjs7tx5WANnBXbGPuvpPg5RhNvjrCyqsIPSf/oE5XvN7ok16HnhwMXrMBXh
wp6bqdRgmAOGkTk3jBfMLy8Ti3Y/yn/SFR5+xzLbT7jqE4hFBb9ipzdLDfi8gUfdE6TkmZ7TYnJL
1JDq9kRRtPDKLDRWBXwhs9glse4YArcMlBGGOBgwolUzEHmeu8Et2zYNAzTdDZeCdCAgnbMk1uR9
z7MSWgotO5uPRlkbi2ZqruKGLLRDWO1fYncYSClDXLf5j9IvIdtAqZdY0AVoS3e0zeQbIRGt2Ygs
LBzhI//sGcFQfmBhU8lupPEsl7wPPOr7YoLZaSQ1Ooy7QcfFo52NOsylpGuIxfBeAwPhSSedsTMU
ASJ+uhaBpiVbsPLISBklw359lzFlxG+CY86fsTieL+z9y8TZYvDAZ1/XtkIERYcZqvl84ELA7lDY
IlnpXU2Ffu2zhMPo1/pnrg/eHB9YKlBelzfub+9exCwPdnUufSpZNlBXutvKoODwaiHqwJg6UP9j
tRS9UgofUAkJEaeUFokrTkTzP7dYTP3DUNYDU/6KDBXiUtoVHzd/WArHcxUvHyAyFJmTt7Nigj7c
v0DTsCtzzVx2ynNLkXmGKsjJyp7Sw/uB8HdcUyh4JoNj/YnajFuq1ux73jDDMeQ1s12Ag0fhBmqG
+QQAC7Kgfas9GC+t/aZj5ur+6Z29Bw4ggv7I6LrCF/hY9tdYcHnJht/GQmb9p+rFFY0Z6ttu2ReA
H+3+cblT63WtkfK3UsScuRFn6MciG6qVGG9vLZ3ntwqtRUIUUVnJ0ZkiCAJVPVX9p5F+noYmdX/E
LoXkOuLb8bA1qCUcpQ4GDC/0hAN1TSQ90ybAuyvJWeboZZRae0ZVoxm+aNIgJm37QUr9k9xGZ3Kz
pPk4LAIWWyRkVorwn5l5puu974fjat5DyoaDostZCFRGA21ZxiyZ3sA8bIrv1frcRQ294+KCYoKF
P2WrMu8UXkm2+JIEfom2dF23mrxFyLyyrD43D02hibu1WrVUjTHOYuy+kt764DqwJHQgqfqlwqJd
m1+/QF7rBCY802GnoMMpFT+pTEyvQpxMeeG/gtM30eiyjySqfFHItz/mc+Tayyi/J6V3bq6N3Rdk
5xqvaf7ld7N2czOo4f1ggQhRO5rBQabRJUG21TmXZGJlh5KGXEUJArQMuqT8jEa8LtdGYFu2aEM/
VOJrkjbn6arPK8G0nW8VTFu3/BnNY61AvM4OII/1uZtRA7wOTgMACImTLqsIQz0fGO8wo397tEAB
aI2twOBDkoNYouvusvZOLQYGZV5oOAxNr9mvQwjQ3pExK3uEIatGTb1jgofuNEfPdC9c17a329g2
JRSuJUB3K2z0989XknvMJXG9f/9OB3w0sZB8M6fZMELzFqcXrWhkc5SxP0XX7y3CQGyh5zjZkhvd
oeRFNR+JpKYhemGzDmicuclSV3wnJkgofpN8SKDrTS9BJO69VghHY3ygv88h2qydBbbRt6lOc5Vl
rLvaaGFlwfKWrGucKNfWKAnE2ZDcH6lqi/YC/7fueNYBKlGYvQbPKqcnkE8uu4CNlwQhYEjYHhoz
BlVbLTCYqJVEwNBYGMr8cpZuRnwmOYykuSrKnGRrs415JHQlvQXGO7Gh589mnWTk4dVe+byYBZKm
YjvmCMydvlahcnbPYAUHiAlI8Im5tDMXsXm8k16RNuNztSmh+E6E3TmBTfvBFAtN0AByVqqXX2St
H+nTPN/YmecvDYbXFenEWLkV9WQQzTSUYq57GlboylMQiSrHq5SGeH0920ALcHftwt76V+hPQRbO
fJ6C2h5z35vc/ILCBQ2LkqI8J5EVUUDOmq+ZVr2k6KMG6K0gFC0Q6QUeWPWukoPULa4XWAOrwyMf
CIok8YD4rLJkHMl/zY1iCmvA4p+zhc0NHeEdktEoY02A5MZ9aURZNKyme4xakFaD3TPL2N62bDJw
GBcp9gDFDU0ZlLu3XTZX8b/ly5ziuSGTyQPTQplW1/M5MiXMKf53ALRsBHFhaMl8wHlMySHPhxEA
yTyXa9lhpiet62JIgTQqCJH29lurIKPEMlPwdHX4EOQ5yKY0S4SekjrsldmR1pTrHa+CjZ9KUF1r
jRevTB5Zcg6Z5XnpFeVYjZLaPj3Gi+pQDL7e97RU1U831WEX1XX1evQwVGp2nq/DcPF2zsL2/Y4R
QlrwNylRdHfvOBBS/URxGZ0qknbvgJ3T41ZCVh1qROoexr9cPO8aoKZ/GLJduzq/9rd8Q5kFxJc/
1kOK55rMI8SR5W2Vm4q8472xsNbA+QBBPUJ+/5+XEw1/21h8OmJdPjIKerSNS2ISAQDHJngYSH4t
ngYs6IEvchWemxePj3x6zBpy8fj0/oo0AMaNSUrBycf/B5jWDR/qNmpCi7FQqH3Qmtovyj69iOZP
vXfAVcO+t/4w56ylGFZN+x/AleeCU71APdtSPdPsOMg0zp5xREwvR4Uik9om+cc7ry74vpiOR9kH
OLE/TDb/vBy/7hf/tnKglZqNYDI04QXd51lxNeFn7aYGQbm+1k0EYGbRFzNRdxRg/f9p1YPEnumI
H08SzDaBJ82cJogjFwJV8fPYd2+2fZiOMFeL3IERHb10h/HSrx0PzpDgwv8uVW/9ahwdkPHWizvV
Od+Mlk5hSYeatDQg+jy2b7C9lfNC7nlAFua6hP34r+bEbDejIMmPdP3AJ9VIynaUXp6YVk8OBeNZ
MovjdzcRa3GRht6CKgdR37OHIAzywZqeRZZe6XZMTxmWrnjKAo10dm5KGbYkmSfLsYauZAxy3lX2
wCbbkDni3/Jee5Mvin072taaKzDmWkty3HaZgQltKz1tm17Hlceev/l+lqfC1uaT3tUfbbYNwVG0
r4/rMmruWBwBem8Gw4oOTQghW3tiUtlIsD2J+9oohYHVQD5P5/+1Mr1WUva71yf82lXszTZB98Ju
JVYXQb+d79EHHFZMTOV4dBl/VyW9yPKk0VwN5BWxpf8nYfaB8k8Nrq4DKaiZ8qkegRFJ1yIwTiOi
2o9+q3a3ArvUeT1dsbR219fPE4ae4VvDJxUv9T1+qNhB09NRjhn0Gu7pbijtQT+IlLMw2DkZyog0
0w9FmSXC3di/3cGfsNHW2La78YG/DEhv9gkfW38j1t5EKA/QOirEwp1BhFGHI22Wa5JGC95y9U5D
H1AsG2ZeuVPTyGnlUZQIJt/3IVyqTVF7mjRy0ZtxjZe6EI+rtZevitA7Zvwi41rMIOUwk1BwIzi9
S4ytfOPL1f+RjBSCG7zerVtBUwRUkyCQbfND46bh1fuBj03yZ3zK/qseCJ7oMjWnhWgYMjvzs7Oi
i5FiBqrfKDpOlQAyRlxtgDCwBav2R7BO+FJphvN25GverwqjgNSBw6EGRlMGuh741pA0pTixnEL0
29mcsXjOn3VKpS1uno8YD7I28zWKeBidr3x0VW05ashJP41/41a5zgj0SC83eAZlDVi69/c2Eqnh
DjLl3ulMquHRM4qpcoQEqNzYj+AseuP52AhwPJwQPdNr2wFE12rSDizyf8E0lE5QpauRemVq6itE
dPSo75rSF0iinPtISJ0n7/su5r0CzkJOXLfdksCE6z/dacy6kzZn9LNRryr9J8q56ZaLGCnWb9Q8
MpvWmSdIgrfvF6eDncoZd+FHPCTGO6Zcu1647lW5QVoNxNir6mTPMh+YVDCluv77+vT0VFdj3sV2
hir8O/NXesJoZ1Be3i+96o4s4GhgSIkJ29MN+SHootbA4I8I3ICd3yjdZH66lIY1GLsH5mUiPYN0
msjAwIs5QVlqWWEo0nGjqBvFDZJ0DPT9Hjd1O2xm60DWCDrfsMf+uRdCSMbctvGekSQxstDWF45g
UmffQPxhrBzpshumWam9mV2nQ3YG93mrp+hMQM/6d3sjO174/J4H+Z2qUPIZUGl8sFYJ3IJgikHy
v2UQWUR0HXE1j00i7muEhm8M+35HxTFqxggZWrhI0NWjm/26vb7tF+fUcCDqOFZ2+ALJOw81tWWk
RnA6yftubpGn3G9ulcOv4M5/ArIXloWQsdeZk+5qcq9NYvWKQ+6z2X5aOuMb+8hbW1b8rPDhNvdT
7bhruSvfk2loVqyLoZQPLALV16cVZFqMaFi94BpWT7oyGlI8nWu5IdKRDlGe/DZBdRrChoYjprxo
Y2yQl73h0c/zfJcgxI7Pzm/sUkarv1kK2IDIV0xhZArui+sNL/n5Bp7LpjReoAepTYvHyoOcAk3z
otgwd+fwT2grbe/+8FIIAH56Pb/+GsgsaYo2hFxz8TlhsDMrmrhZwQop+LNzRZ29vrLBlsE0g1ex
9ylGIVkD15bAeos9QmRFQEPAzw8jGhLtEcpIaesKKWpuj01NUkgbNSxnVE0dh8ZcoY6XhuHeW0te
tqDPmPIfK4IOIDSzjR4aTYKLhBMl9F0Qc6zkZ9F2Gf6NJcNJdRUBEanx3T8J+OSW+l4y9TSYh57/
K2L37rkkpzXKxvZirouTpO81hvX+duO44CfgRfLIRJon21BOPmg59Gj7fI/9G+jLX9v28GaLM8x9
gizFmw6jK0JoM7tKIOY3VLEd3bvS2dsoY7VL3pKmo5UgYvNTZqSjKzsEFCCAlwNQ3tdshM6TwAhn
EpT6kOFtt7jCDVXtbXc1hoBzpXQocqXwSoUahdnTag6bG3r6V6guF7zJWzYyd6WoJfC59nZaeNz5
4bOsLLGztY1EiII5OluhhyPClPL5E/RpOy/JqL4/o+AfMvBpVn6a/M81/thJKcPOlCZD8WgajoJE
WfhhO/NsRAd+bmD4nmKog45Y1BkYUCELeFCzN+VM6bNfq/edS3erjOR74ylCwcIDQepLh2mjvGpC
rYiUt2nnl/K0RYJIYrgmdpsOGsA6XbE3GysNd/z7yoetfI16jQd2/PxB3U5YLGB0QpPaoezzCKXC
c6KDLuU2hwlii2wsj55THcKH/cuv3T4U0918UNUdvGmKCmq/n9ZG8JDDKIGNpraFEIxw0+Jwqrxv
tb3gg+1pKh0tBXMWd8ad1tPq7+qJsCD9otp9mUD5ChdiiEiCFYPDZB4yaWU0fYCat3GqQogfOu8n
uZZXBzHuuMsxrHgy4OhftAMHEeV6UK7rW6jY7RdLktgPHdSRmVx1l1KYJmKhVNzK80DuJ1qEUAAr
cFnc+Nb84CYv4mopLuz50Yr4HU8rRjRxMLm9ZYPxpUox8/nqdAiiHFMnyNOaKLOA+kiFtGk2dTwZ
ab0yJnLApIOpgxmPfTxHZckEGKi1wXim10GIp3m05BLPhJQi8ariZlUDeYzOWi2nRVJM1tBnkU9X
4oin6wkZkcNVcun7EBkByCk77qmUhaYc/xa2h7DHKNSgJd3HzShLx0fA72OfUP8nhiHuITKtKJtl
rc4iuIazOupzajF6Qw64b7ArALX/qvnGkfNZO7UOJNE8/hiLWPwEoE+BwVTrnoAEj+tb8d9wzfEQ
/WfAwGY/junIJ+qANSONgxs7+wpN8l2B/2UOayf9aQmpfhAGhmKj4UqTfdkGfRyaS6wmpadjpra0
tagnfGQ8FOBVZaHcEW/1nhLDgV1kY5JtrfUnwZx9uCw99g7wCAQQiOeMHv5P7q9CVcO4qcSr/s4d
4vjAiLdo0r64SQ7I8H0p1m8jHbSGVudOwPbr3BQczvKta6cebDVJgClWacWKk+StPJYtlbIyrLKJ
bQd35SHPUQI0ocgEVcDmm60/Q03t7H6YEclBIQCjkveqQgUQUsliFQ8/Eu7FjcmAZ7GHrdSYDb7J
Wo85eBn3vhLst5c9JuPcgjMmEO9JIoBUGuZK0jaQdW98uaH9Ss/l0PKpx6YMdhO0RFCxpdK1d4nP
0Tzc7HpoPpEl70uolkKFE1vWN4EnnyEX+kMfccP+3Q4SX7xfNCew8hC0WUTPalTc4Y0+HLNe03aY
aB3s441mYp8WXb/o+5O3//eSbDC7j3gZRkz5Fwo1yEljPe+bTVVg9IjsfmVW+C4a88J1NVa1c6HP
ndPGqmkid/GX9IMlrfd/WXDlvjcv4esyMv5HniY/Om2BmnRP9/qZxdITC7G5B7d1v+On3WUWmdHv
XbN+7N9aK3xcNem6O6X5bger+GMYcRG26uoDO73wl3vKNlAx1XGJCLQi6mthSRhvJJWJTcOdapWl
xGA669CXAF8IhVWLWArUz7HWQEnW5mqCcmmLIHahEzVBgru3Obtr2viAZSwl6hYPu0T382VDkwN5
IE6caB2sv6AVq4sBZUD3bq7ITdDEcpcHKOp73QY5mpUyeRWHsjSnEr4IElsYteJIuhBnumq6tazl
ahcpOKps/ZlPWFOyRY5URLTC1UyIg8Vhk1ZuMpfU8L9fVSvu+kt3cLpHh8/0Lgu9n5oeawz+TeNx
o/di42ZN3SW3TtRSS/WnsSqBYOMbRntslFMuSYtBh82HGaTGLNRqajl8lbjyHO2eM5e9hPqGx+pD
jn91AgrR7w3nfKoOXw1MlXJjyWQ5h6oxnejEYhPRU115DIl4mUeZxcM4osErtHvIbvYZaZaS5GTL
oG6xTbxye/pnSf56fa6jRB024FiF07xwzxJUhOBnU9KutupE2GmXKs1T5aSqh03n52/hrnsW63Lf
SCjecupHMtYbvaezw+n4lfdHdNphuAJ2h+NlTwMEApai/HhGGcT1el0AN48Z37J4DL+I1CMHOGdB
Ht/jgzFWB3sjgOwCm+AemtKB5atpwwO7Dd86kxOrBd2xkx+oMeQbXXCpEtPYSPMd1sy/E7y6hlGu
P4Gl+Zr6Q1cMcXYAPcuvPTa5twHIwQ+y3XoinDdPp5WGFY2B6ra8V9F6pLTTOfPXaju0fXz7MulK
Xw1ajvSOKJLwralCgrjtldCXiGan0G3gl1A6dLL1GPCncjFHo5r5Imfxy5ImfH+AuX/Jk5/LPol1
Zp3Urm+TVjQ1NviHwWH6GROqskXwY8CNjKrpXqfDO9e3BRBKkdey61sDUSXUt40OvVGl4S5y4rf7
oeN7herl/8cTiX2nEY6AuuqtMEZuuI5HgYXInMqUGAGqFDIEQ6D9+pp3r56hfghbU1o3P8fN+q40
EDWs+ft5edgPxQf1S5nIAyeBLjSAyRVsfSMMujbNTnZ5YZOBJuCen9wuduvW+Ew8LqqQO6hIwnSm
QdwMp2vcLTC0OC0Kiz8ZyNIzfaf70Itjk1k972lodDxsRvK9JmeKxeQ4klFd+PW6arBrbBSMF/6g
+J5CYoGe4ZAlvoU1stzfJq6uG0Z5J35l/cWCxvQL+vyfwTQk9O+GnXlu/pEMOekI6VjWvyUdTGjm
da3tlsqm9AtaKps6gNnWYpRfeILgTvI4or4yffgiFIlT9g69YdLdC04EyO5HyJ1WjqmE+liMt9w1
Gv+2cohUi+EYSzguJ7+iaA6uY6LkAQmpIFSSWNhv7o/xOVZVu6yzJaHqrAfV7Ez3DpxOzq4Wm7p3
QCqBQmE2jMTlSXi1ik3PJ38lD7/NkhNDj+lXyqVZRQKXdsFwku3UN+jyGxdlV7e7/pvbcqLkRG4L
pnoUmISJaHEleVvXSRLo/ozpy5w1PNK5lfShGaJD4HdBb6S66WQdLeXaKykQMmCcyPIQNWb0gWeJ
MSI/XxdRgBIZNL28lwDdmEQ1LTC+Vuyr6fuWdGT57ij+xSW71JwuHGMm6nWorYuZQsy5RsiJ1Opt
QK6YlI2QeT1UBsGmYWE3O2QvZPyGaf4W/cHifbj+b7CXUtVeBxMlh7T4yXCZlFijNAp9IxLIO2ev
ZRcKJDs2R/GPOL5yCpo057MuNc2KUuQqg6GILTYHuojCmAVvySIQga/z6JF+rKZvXBoA73yOm1j2
eVv7m4kC4dzizhdT1HQBooPbfOQ4MCPOBuLdEjtKrE6qJVZVAuaXycoeqpTPG42thEU+3U3d0GR0
+A1Q4HO4XlaVs5ojoOKutJLxoINy8DSQVpYuS3paNHGsBkM0ueV+7mCPpq66/fKeC9Tzh5I4U7Fd
aHdHYV15sncVsQeWjz6Qd9R1HSK+al7b0AiuHbrs9g1rn6GX81rdvc2TBwDVxskOQT3xiNtinlAR
9d25GSIofohSI0lx9oLzXlDMMkKv7bg8iS+/ee4bJWuvQqo0mG5zTbiy7Rr8dBH/luthdRZcXO2e
+ncnsAugM3S2wrXQmWGeCSOTwswRSUZYUW3EYf+vAl18qX4bs72vRlfRrS42VIhaOPM53cw1XnXx
zJuUY/W3hT/ItAi+VAB5Diy+H8zYbHTXMbAGIfFDfFuaPDZYuBWJXsQE7+PuISHOAD/f4wRypOcF
7wibNCtP/qGD1phb8ez3wx67k2/4p4c5zVc3s5W3TdTI/lTYm/nByQTx+c14O5sTbf2/FK1LoFZ9
0JRjGLhVBoOkJ4a6fq5r+FUv9O8RBrXHW7fccoS+bDqoimnnmUe7ApIU253+DXcc/vpa3QqdVtv0
XvmFHNZV53f+eqjmtDyeIKUkBk/rHPlLF8AH6q9YpMgbLoJcpQYJveJ+xgPrR55G64sEYWXs8AXz
WUAh8aHfEpUHGZGt63UxWgqm76ROa1bWQ5PgoNAfd8jN/uv0j3X60gLRIwGe2f5sWYVSFhK8W+sN
YL06x/gGsS9tIC/vr+ppJwrDypsR6LzzUv8/U02gVVHBLEtdQgLIlyjQeyt9DskWaEH+sUrpeSPD
h44cv8/5fNXEYiOlqXNO2jYyFihwWXDpefUV9SdAp3K/xJFfMe21VeKvab97TRZwoTrQ9FXTlTnM
Sxlxs1K/fd6txEbLsvTyU+MaYqc82QXWlFtGQwGcTHoAR5Vq0gSrspj3Lnc2Bakg2aACtONQcCXe
qdEL+3hkC37O6/RiN1UtMAtxhCgDj5ydYkto7f6ljFKJP14RWqi3DuYQLHhseK1w0vIs4odzyanG
3RIaK3VgBdvvgTtiP5LRsqYpfbnsA27qd8HBkSiYhZgyz2Ya+MMHGeVd9YtunnZESKQn9HMF12FO
h72w3udWH4Se3kK1DZ4pxBC6x6Zzy/0ehvxwDabrHYurm09EYAfhvLUI+a731nXEovs5KcStQxrA
a0gtoSeCYvYxIzmN+1k0ADYpQCq+TglRvfl5M7OUkkbo/RWhMRBHqZ3gyt179/DqKGRMpJSc/Tkc
SX+zstzJT4Ef2k4fYGMSyezKeWM/9Nl1sxDhe77zjjDJAL+CaKAyA79hEtQNvr2kv02R2YYrlcPH
Hi1luFkrnVL1dl31hf6ZuRthosebr4w4ZgcGgXuZRXv9AGO3/xI2x3g1mIRDE6Feb6ot2zqmYKYh
6qEKp0b+HhzBNwkxYcIlXOe3/dlr1Iw3fkqjfS6iubJ0vYYqGVdz4DuqN06EKDM9wbuH+1H4h3By
BjstqHkZQkKLNPc29q+SH9ehMvyb9bQOAlMDNA1ejw9oOQEMxh4nWz12fPP4YLvlEF/vAmpagn8P
lhH+ILpqul8+Rj8Krni/VJjATu9LuBEVto358lJ8jWB1QgB5R3Ad7YklWsNhkzaZzEkRN+WG30eM
Kio4++ITIBRVpkfLtJhIUvKvhmRi2Ws76a3LAy3RibIL+a+L93FdOsUfz9bEkiRyVA6U8JjcwUJU
NnSl406AeD3f2bxWzZiDWVFd6jYbWROmlABynDb2nqmRx4etyw0BHCLImN28ZIimnUQi1F0NEO7L
WgrW7/UYrS+SDWYjnJKSny0LQ0E7BfYta3C0Q7tSmU+XjxeNsv7GrJFpSdMa9LEb0qqfm81QdtDb
V61cYVTAomJo2m1XIrYFnTInQM16gr/IzkVOW330et6j4f1sC39CRugauR5uQoARwzqChmkOvIK7
FCRXJAOoiK/Ng0BqdrTrG/pgRQ6jIZdKsVQPeK2hmqLQl88thudczBZpg4YOz2wX1fOYtYrBzr9I
6uVwJgSMgc2kRy93uDqZNppUw1nOrFU0U7JckVkIuESOV2CF63937xPBfN0xM2SxLoLUAGmb+DXn
VAtmbOHf2ZSKG/UdRcsjwk4uJb1BauoQiPJWoyjSPhHVkf3UNaV8kGWFH+qkO6T0c71sA7fLhAIb
UxMxi3oFaXyyxpZale8Hqp9X4JdH5Tx3IlxBJt8FR2sycj3Ar9YzFJOYp+Ytu5gpgn1z3CK7LCD9
R5/JN53N2JEs9qI54ueVJRXuFytx9+V6kKKhqzc5wpt/zqmEJzuO+9K1UUR76UXM1crfkU6qsVmu
VC9QcQ2KMzzton8f5Iv5zhmTG0elSo5pPn5DkZZqkqUPLtsv1rE8idZHR0icrlueOq05rhj7eQtM
Y0soIjsweIiBlcRiDtJfHBtHYCGfLwEyE7w6PGvVxAUwDAQ8AIdGD/7W/WKXtcXwrPWQR74wuofg
hCiRiXx5MrPeEi1vgwBNbasWdUi1zAycqZnUgnSr8WxLOnbMLbLE7DSJMDslGnb9avNR0dsojSkE
8Z67Dbl17Az040k4AWMP+hMVuMFDmSFAb7DM8b6Khrs11tQslobIi4Os/dVQe36n4swcWx9O3vMq
83FD3czrl7lctjmjPIYacE6Rgzd/rsuyJrPhFLIIi/0K7mVpoBgUoudt0pUZqSUna0MXrN17f+hi
9YUj6a2itrUgctkKMgv/fP2eIT+cx43oYMCTkRgSlUmYhIGm4ZZmqNcc1R/y0W9R3KaYIBX9QX/o
O0+eIRjM16Om6Cl8PonrYVnNPT8ppZG9qIosvT0K++n+JPTiGC4vrfJReR9ob4uY/2v1Jm1SpLm+
/3C6nMs1go3SOMTAUJCraAw9OwL61RnwLbgvHeRHozz4Pg0fsmeiifAk79UvN4Qow1pkK65IqAh5
3ujlA5ml2pZr0ENnVzuzplOf1dfa2FI9L3ZL6tPgjfSkRuMFp9jcvpAlJ8Um/9dOadLcZ+omGPa3
v+DRRuxAyJAgw0/nwZ1MaYwmTH82XrYhgsC8rp2H5Ai8VHDgMsSu7nuPbna20tN282OkETD2zmeC
OjoEmF80FaanRvCekovFaboSusDSoI7lfyTPEu09PAbRcmEatgzj9onYab672qm4/sgV7wlY82DR
UAeUjxRDEq8vrtr/6PMhERD1RKT5znk3a3FtobwKEqysAIqltaKeOgNU5J6UkUFcloBQbDVPcaVm
qQW5cuL19+ltrYYNsqdQl3RjXhoitHLNmLMycj9rFjPm1GnUKtPoIOwHezpzvrXOlUeE18GlPG9J
haDb04/lj5aL235Kr/qZxPotwhjfKNwoR8V0keP728J2qBeFyxltpxUOFBaQdV5pQkV9irGth8nk
Hiahxwvwxj98wzKvN8LQSod0hc3z8fxQZZbEoBvWPzDPcmDURKJocYdnLo/Qe1rfhwaRWIFLMKBP
b2Hkls6yWHnQT8QWJIMpNRnPNQvwMxETyvF7QFR+s6M8VxFITFtFR7wVIRW0hM2quHVC1gG04/6J
b8wo2NoKjQFZd0czC5CWCnWd1idoG1eMfVezlRL8JN9X5hXcppd8OGDmsOlQKWkNbwdOwLXexJtq
Kenp6BpmXEDDu5iFqwRRPmnYgeZhiI5vIJB+cEWvSoNUJ+hlrOsRl3r3ydEDyFTWUgsulkKPOUqz
NJuxBLgNq5kZdEhOT51yJvhLlhBXyD9z6jLFWopwR4ug4+s6EhFt40hmlYD24u0BEYCJhHblMx0K
HLWnQ79d3KJnSvTCzs8OEJv/B8QeuO6rjQASS7TsA+mIuLiftUhSJZ7l9LZzuTDYUwGlySnVZ8rG
oCIfkJTjWuFOX1eG/SVE0w9nfIpRqEKyN2rL48bm+IrAYRHTBrmS0oBmnV+2wwIM2TweEkEWU97y
3loswWSPC4A9bqYqDWOa/n8y3wUua5ChEtKskxIJPAWqZndq/00trEDPjVyPLY8+g6CKqbGA1H3l
J4g2dojDty+5jMDg2G1zxg19rgGlJ7KshV4d0MjIaxwK2/+YmHcEn8nel0J6zDkcwp7I5arH0AXi
ogr1rE2DnSOGjgVd22BDAbo7VfcHmbgVjuE46ivWu3GtqUbnWwZOJZ/aBbYX+6YQ/1QYjARR+Ati
5G6YHB5KOl6L3BoL4ly+gxk8TU/7bM9OBl9Y/aXwRnRbE/ACrIaucdpGIu75axbDv2QTDnAOnItN
UsZtSy4cFyiCVi8iIQaVTyEJEv65IUsVtLFfkxj8Xr/PJRvW1TMTV+R6xzCtfMzwDepwr5CcQRof
sR1/LTBL+fxNrIsHwe5CXH2NFrXwJaLiY3FUNw1TQin+FDQPtzt8/BXgiYSoD2wAccdCK9xyLr9J
hs+JWY0BwwqQCfZOrKZU5h6Dur2r1x7qbc1e/uKcxDJv2eVKTzgL7G8YvfW9ETJVUOmzTEZBBlGS
QR1dGdAxUCS/tZbQajvQnzzJdwghsXbOeCXw69+6fLOiQiTcudd7E6k7isYJ1KM4k721QduSngJt
xuF6Mny6WMzCIVGFe3Iesx+3zSuldZ4soFUGcUaLs0dtX7EgLXW0LsP/Hf25mrZPsbJu65FdGWQV
hdDTWV03Cv/h6O4r/8xYaXmf/stkM3VU/d3p9w2LD9aiPNqyGyfOSWw6q6F7GLTpnKu0fg4mFo+O
ASKtTwiDU6M+kEu/muezJEyTmSno5cnYWyeGVPe25s4teFsUH9QxWvR1vikIbKagXkw8kLe5o71D
cCTNqjNhEYupVGBbQeijWpdvoNv/luIxCHJos2TpAmdAKnbrx8KyTMtw9WlnauXH7mb8wJvtzcx8
xjiiVTVpU9IZH7xQ+5E9d8YIj53gJjiVu7KIMAuyeikQZDeuBzTk9QKJf3QkoloV7bbZqoJelVc6
MsqQmL7rqi9Xf3N1S/csAkvrqpgMCAYgO6Bkr5e6L/XISk2qzWgZB9G+33qvxNHdhaMBckmspJxX
K53yONhW0L5VR7sBqrW3FLFbTpPvmAiRMBpb7QTExbNfl8kZ1zYVq2wahhZlKNDMpNnk0r6gw3Wv
/NPsA2edXA5GEogP/+WBS1Pq/WxnoYZp+FjjziKIb9KAh6VNzK1Q4BII0vyciS1DqSzRP34PugbE
TKJT3yZ4sIXN0oF6UrrgkgGX3WzR0kBeMIw8B7vsK7RKpTY+0mSAEZr6WDC2VkxoVXqqLEliqvkh
xnbTz3iVmkXMl8npoROJTXZ9DLHxQibTplbjmAU3Wlz7Z+E6FCYNln/aORhjRvCqKuHoXZRlXYOb
cemp5iZUF02gy/usQFcpGzJyl83ufPUBerZ/4PGwEC3ExyDDwl0Qe3ibBW3sKNIyGnSkG59OEVf1
5pUu+US/grCbEE7dNSR3qRhQQxlUFaAucrnIjVS6UXH5sSDTOJrzskjqfj8NsryYTw1JPeAGM3mC
TG93DSemcJ+RfVNAyaBjimCTuX2jjisKnGVHj5SW3IGA5DApahJ0aX2v/APqxDz//PM8FxsPpvbj
Vpf+FOKOG3edLOsNNgQku6Drr+j/i1fwFciq9hV/6LXmSzIKvENR6OBhe9dzFeu78wqRSlZ7FRa+
57YXi8SlLAZXE1M/nV/FfcJZ+eDa4dGzM5YTwBgcVxmH41Ifio9/EXaFuuoLG6J1S+eof+nBMd9U
UInqaW/Q3v04D2ej0S5T4opT6qVrDxJeBBQLt79Bw0JeLjmgjNy//4F4+0bsaMZhgaKoo+InXKtv
L1hKh0oZY7OVaZrQZ/v8qatO/CFU1ZEIr5+C+VElDiq4bWDJ8EO2F2use5f62B9ODhQ0DIpWcslc
LovJTOwFkvtoyFd9/uokDeiY+1x1am7aQNO85ovez52Mj8SEypzw+GxHDJeKlZjlQNHH2Tx33kCA
LwbE/tzltFELJ3u/iLSlU4oNyLKNCatPT6KXELk+CszjCJUqelM0j50qMweRtw+39PXgA1gfs/+Q
TKoSsQbSvKPayz0EtK8cEubg7tEVMmv3WOiiOKM994EIzcnUJN9z+VDZupuCl29JP7ZtazMVwI56
uhDiH5NP/BgAre3h0TWwtgGUOLA8VK66ZBGR49IgJMr3r24ns5ehnXI0k1gZgfQytvcA1PG0obxR
d0jCo7Rnbn83So1CxXN0LayqMrwTJ1VEfj2iYKKkT+Xkth/ZCEpmFP7VNSTzIkdxoDH23X54rcrb
LaQcJvwShP2gnNH25yJETubPrwa4x21MNUqwHV3+2HBXndk5HUs9iWb0bid7aij/z7KqzprOskMM
1zDeeXmGevABkNpPq6MdGgAQzM7PbXdYFWmdKKkuxQECHR00FrTgmjqHY4gO2rzC1F51fEdVzywd
3P8TWJEvjS2+FgGdklPCa79VVrT2miefItlwHU8R1FG4muoRdbHzezsowGWXUlahpq6dozwaGT1B
B4Kp0ZpTD7xVpVZj6PYuhLyv4jHmsotpBolc1xpa8SznrBqb1bADl9Jns2kC/XxC28zV1gJrcnb/
GULOMtuf6DZrKZ0J9perWIHd5WTyPhN/Fmk2zgdtM6Ks1vE3d9jngmwWMhJytfrdKl0ASg2TcxCv
b7dsNkSu15ccsAdMDWPp4kvew4Ai+y2M/O311bI4qeruIOiicQeXh+ZLLEuEc4jaZVevmyjkZsNO
KzT53iIbsKg8CMzdi8S1eATHoV5fd72dP2jZRSTsztFxPar+qmaupyO019zkhr+MXEM0LRzZohbg
lgSUyXRYVinhe8BzX+CWTfa7jJqePyA5NX8nPm4m2TVwotBrhG8GipR/Q0EBlun6TjQJVZBwexyC
McRynl5ezCTcEJGzKaLsNabNZxvDIqIXZEEd3nSma2FkhEEnA13kvCDu/fr6O+RUA+lyESmTECRu
6z0KIfsSUmvhLM3HHOYINkctWgxK8XxTQXI/edY3XhUpwCadijhakBr9uysESbKo64EqpTX+SxR4
EXIXpSdVCuGfy5VQl80U7iO/78hcVT8Y7vzXHSvirbb2QvNOpksqyORmOCbpwNN+wOaIiWUtvc4r
rYqLHHADQya3XJUCgd4B/wTIJnZvtuscN0NF1Ob3E5w7DN7QPimAIGX0geBZMO8FxCa07uIzCBpM
QNs9SSfjeC2/WkSiPBvFN8M/X+zI1Xr3tBs=
`protect end_protected

