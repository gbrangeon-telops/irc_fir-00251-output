

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IVTcVKz+qqR6KelbIxn6hKss0fyLwIejVgwej+TN1ST/vU6syUW6hxZyGugx/VRu65UT+0QU+88C
5SDN434/fA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W0uuDuJZlgdtFvYMz+doOP0vwnGc2SXfLiGH2a5FulZQF1GjNx3fjKnarWbbCm92Rksm2FFSGof4
SgtGKAeCq4Yz/Vqm5xuP6QHmdBwou49vkKDs52HUud9c3EaEYtdNlkb4+DCcueqZu76yWN8rf2DJ
ekmu+LGiL1dmyzv30tE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Da9hmR0COgf/nsNRjZU5mrjIzRjN0/ufJQ7crbPh82WrNgInUm192216ks1D/Quh1gQ5TieAOChY
26CHNdLfPPmjLAo5/cOIRsIuy2JD7JAEIDFhFO2BcC4GrUAhSArSC4/9FyqXrVJUKuDybwv0tWSf
qpHjmJw18CiVw84ne90mESBOJ0fW1ujayfbI70yaGaFjJM/DPm4Lq+TC+TFlaimxpTFNrAUzQNVF
VSkf44Zb11D7if2jaL6ua4hPGgYpPcisaJtcEYpURXS8Lw+NjmMExnMpUW39NqnMiTEPom3YBwag
JMKm6/EZOnBvVc8SljH7y69fXiGUXgw6Z6POkg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1/llP5a+sEX6Ky1I5ak8Fr3e35uMro1bXNqkrntPBRVTqUhQPFl7wfr/6Abnu74l73YggylsZJi1
1Erm6sC9oDhL9IE4pENErrDQRZHuFnl4+DlguLd11swTlNfBwauGoCBXbTtZ8+O70UI/sRzXqbZc
NDH1RywyQLhMRmSOjCU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OI4vyCtRzSCtjYNsCqL7rYkcvPw30aumOHoxNPQx0NU0Kc5/zvGo5pjE7sDqPsv0b00mAjKXUE8e
pVllo+uquegdt9Smrq3DaiQC/9hKGiZzOG1rJH9JbLcfPMXDGpwm1inP51BNgkQwocfUEAVndeWo
GE1Y28I9gt/5q5Fs/OUAX9cAh1VoS1OcnYX2wbgJSlzuLqnGWRIxOHl4+NkNkBq5Q3Xm589bPnnz
m+d2tBEPyqaCTvb13xXW7hqIf0ahuv0AQTuiClY+KmF0GjLdJTWJjDWPuRd9WYhybCp/lrgDnhAK
cnRXJnAOwP1Vgr7EPuoyVc3UkNsZTxEr3wrouw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11680)
`protect data_block
2viakGP8XHFgRDd6v02pyn+r285gaBNH31qA/G5g8z9Lwg8qM57V8M4pG/e23/7x2GHHtmi72aoE
u0DW4dy1yr8/UO4MBxi0aTwAicFPHSLgd5xr8P79rF5afpUtNk0sBSeKmpT3SXwCx8x4wH8+cx43
djcNOTVByN4Zx1Nupx/Az+BBL4K7A0oUqtulcBWyuo7s6o65p+ABGEM5t6akFiqtKwPx6qLR2p0V
nWbFT6TfTJmHoxSII4ZRUe6BXQXKkgbo/oQUhRvwGh9Q9/tB94g+WibCMUpUjrhpmdrRZ+Ytbmok
+SdJJ+Nbtvzwp0mXHm0ZbrUOTRO6jBiHwfhmmVkvqFfSKpfJ3iKWYAveHPtg2B7R/B1z0JeSgPgp
dyWLic7DcASxMR78oXMyOqQZ1GROufwfP3hGgFC5TvG4EetC4gOyez1biDSaVF8ZZ4HkoDrAzD3i
92DdmqpClxEoMwgl00HVRO0ap9CGyoCFthveqHF1P1VZQSERurtQeuKGZnorus3EoML3lBLTuVUz
IF4aO4nhxyc0N6RcrhUPr5eoiQcrMJN/53FoyjYahAsrHKAt6saBzkAhGXeimcp3Hau/DQAmIYIP
Ujqe9dY0B35uEfo6nAQN4fWmmIn4lDgUuqmkoWxZ1iIL9G9ABs43lpTtN42Atu3kq4iWa04OiGaV
anXg3wxEt5+29aAtKIDkbd1fS1RxqaKvFre3IN3Fy56GQJwSMpqp+7IgF1U/QD5yp8tbTNAs8qsP
bTojdak7b7XiV0Ft09L4hhDYtnSljhGloPqB9lP4jHFm8fX1YobZ9J2MLFFJpjb2mSIArscNJeQC
EsIfo46/Bh/iXESXi8pcwtqcxQqjT3lI0aB7YPTYJpRdVHBZ3PXEduxavSLGO3Vy9H0ALbGOzO8T
r4nmnaxhCbdh6H+JqYtCY4POoEQa/rjogJoHheWE94LjQTTtD2Y9PUHp2Jaxn1TJOHYQhJLMkfiA
MueqnxF5eFP1TvEPQdufLLdtLOhdx/nmM/hu8HgNyd9dLzwAthBs7LdMc2eoI2Ya5iCz86e4l46J
4ctBGMBiOHVmEKiE1mpatPiwHHR7yTu8NjT8t1IYNweXEwRcFXW+qQgC8bDJEIN+y+oanTULVyqL
ldRfYPoG/IpL+BCkGEjP4sQOjW2kWwoVcyHz6x3RjIPhD1anpK77uV4CnUo4MzsqzUuEvN6X9Hbi
QBa9uGHneQxHFKOBdscPc7+IvIQaOzuks7XgSUf7Qu5wNbz/zRKE8ie2FIzh9wu8y2aUAoi2fKcm
jTuWVnQmL5c+hzKrF/+aMJ8CUCZ/sAmlZYrX8wlqut/h1RE2U9FHtW4aO9ZKxRE3Eu53ginUlQBP
ANNwc6cRJBbXk/v1o5Ti726ijAIZBmRHhiFV9O7yMjwVpzAIDgTwV2DnKMC+Gz5WYhfTpwwKU0pv
k2+MLtNorWO7XBNWfOl469p+KNoii4H57Lk5JEpjBerJRtHWsdzm2y6DuWN+QnGpQAXA3x+rEVkh
6EylNBNdIQKaTBMMW2EssI6/6e9Ckw/rTZI4Zp8xqkTwteTEglIY7nnYoBN769FkqcvLUNaMiA6w
FPgDX09oDFdYuNna8s7CO0AxB2gZt9bcl6MevLd2jr7abHJWCPekx11sNnv0ugS0PAVgfxE+nUhT
pwMr5XAX8LePQ6Ao6BglS0ZH6uPoLD8xfK+QpjDnEUxmn/ceTHKVF8l/JEMwc+IDTHwAA/9Ddi+K
d1ussiUfUSIVRlEdgECkKAODyU4TGPp7nql+4Fx3LOpSu6tkWK4E8bgotAA9V5PAkPpi+kPP/HQB
1Ku7fALVB+V+j/MfxreJH4UJPgHwqG+s3OmO1pt4PDCHaqY0ObB66t8vnMcABjI1TLOwBwre9a8d
9jd30HuBcfCsCQippj0wbLMRxYw6Q+eu2OpA9ktx2/DtvwJthFwNulCiOI8jC+gTkm1PByZs/NQK
Lzl6lkIZGhJlQhfz1/t1PIuK2KDHLWPZdLGIrdBILDC2F7yBdFrI72Oj8kdCmN8knG7IaDoc2sbZ
Ui22TjXXPxGIc0raW30eegUD1iKiCvJQ1CcbSimaUMyqnUxJF4KeLpy7i8qS1K/V4zx8oBxfcVEo
IAo00gU3fT6J1KDB9TSif9Z1vQqR8XY391IRAGnEXn1/C4Jkp7TMph1cxlPgVe7SgtWOhHAZQfkv
bGV59LfgC7T0WPPB3cmfVkh8ww48x2DI2ZgJnlw0UGvkkUOWhnp99P8ZNRp/m93VKRCwz8zhz7id
HF0QbXepAl7h5L4CX2votvZZljeuK6JVO2LRLFG+LAsHz+XjEEgywBllpHBzdC9+9o66Lq/qzqK5
dtpzcwSnU/fWpEDFsd8I/New3ZHL9mxTeW+uDWstx4scbC+W/K0EGUoLpmwY1q6rdmQQWi0S3Q0c
6MBYUd7Ljw4LxmOyh2RfqZ0JwYD7c2TkB6ejV1HXi47Q46ptgY2ZTCYf9q/9Dx0l3DNaPD7oDpJ5
jc8qrtLMuASQWuOZXWzEcypdYqR177IqtN3Q0LyNyZRmwF+KBworxFVYNPEOxcmdlxZywMYhFNb9
mpGCRACZBVxKFa5hr9OwrRXQEn2c/dOjWQaLtkTMuHW+aBVdAWNY1GAs5mT9iYT8u/l4obW5wk/Q
oBV1zYjEZXtLpV820LgxFO3oV0qKSb1Zgdx8IdxqHVbVxNB9FFUj/Ptms+oLdpTKa064B30K5jOr
AwV/AylD+l1WhchvY0lF6MIJYrTXtYZ9c1M+vZq9wPJ3Jp+1Da7uK4KlOWTffVIj5qAS2Oe7GE7W
rEQlIVpzC4/rhLVKsWiXl+jasGZkQLz764qevXOdXVBr+If5sRNvozGsirJaLpxi9TWbNMl2oM5m
C6otLQUdCd/GQTCEZUvUajoVK45Cxt8GNKIcniEBH35cJpQzEseEYE1xFhdxKjNnUwzpSG9kMaA+
jB1LVkwm/HybdxC5ZM4y3UANE2kdihQWYUWHbPQyzu15vbiz7A9YmLzpNKn1ADLtF8oCLtUg9ckA
eQDnDoLoJaBpopPwJ4TAkZNHsD3P5etFYcrtZSGoDp5E0eVpqA4hF0CgbfNr42wUvRQloz038u/K
9buPLeqyzsMasmc9TZkmcsIiSYQssC6sEqXi67YNI14Lh8wv1G6Am175YAqxfLMMOPzHb4DIho4N
yw0xn/ikHnuv4YtLF05SM549ZW2lJCjAPjE68AbNVq8STLNl7b317G3Of1H+2tQbwl9WoVvwe+oe
czvZeV2fLv7UpZUHxhT+vtdP0lWhXckG7/4I8DAafNmekD/GwhaY9zFEnGKEnK20NxmWBeyqQ2G1
HTja7okMF6K7QQ2eZmzbJDXa9OcSqsB9o3OpRApy5cTnmJUUQIzqoxtMrxleuEgWPnZVtjcweK9V
P2QXJ4xP232KvpcSBzHnyhri4kOYwFllw9EC3pXzN9QfBUYwF/wLWJJlbytHQZc+eOjoPYWnCiA1
8VDTZoKKigqsWTWnS53mB3X4rYtuPK4HXJ1ObzGc9e7OLHV6DpYi9+4OPwRZzUbi/KkJpox2sm7n
EYUUxBLq+TpagrmCgw4GNL+MC1/yLkECL8CUiflCjwMR/CTsCsQ+F+13HX+TdmALPRXlIFTHJSeU
rJ5Ua88MECIoMs6Gm8m2+2XHqyrtEud9QTVojhtjKLTaYxstiloeRI7xx+N6Uh1tuCA4qtEjOTgp
Mon86b9wfURAsjPWP2eM21svgQu8aS4R8qBjsfjZc1jPIYXRYRpdcf7g8y4mY3mG1EdvWbLwcspc
SMuw0TOGCDw2SqokkBBYdbXsBK03SVGcA5nK/ofBrWRTuX0ufTIAgBWBZgl9XwQzL6oG7vdRTTSV
1bBsHmVKQGclTERTKU0wBj1yx3kQWpeE/QOXNwY39V27l4ePli/3A++w4GjKhSE7Z3OXsK5qP5Bz
jN2lVDLcE2d60/D+/X6gVN3zffAW/uwCfpZucoI50ImB1cAvF0Z9YU0c4szxHLq3L5KdmCUQVcr1
fDOm+FuAaMWoXkl7djI3HHiE5FGs61fz2VRcVyXlfLkBFNwNSsccIQwlYpZVdRY0Es65smVlOV7E
MsIKMBc6UF7bSD+VZb5PFGmmXp7/ax4WtoxmtD1A8AFxv/FReVwGa5d7nzg5Jbn/BQFEk92XJ0lZ
5gamv6/UYLjOKJl7M6Xs9obOw3DCoo218aHeC4vav86O9Y5rtpunfWWJ7x13NwDqzfTnaqpGDVA8
R3gBLF1e1bvaeKL4wpctdMH5ULBvoy1xpsDOIMXBJIeJ0GF5MApakrgOLGqT2FjKUhZZmL6/IlJT
NMG/0a+42b3bMfq/XrUvRz1NHhp7I4dgOWsca2idXU6tJiulhKiuPtBQfMnrE3vzE5UAwhONzjLE
QLzVRbzV9g2NGwfXgFO6daoO9oVetSrEgMqlMjlE7q8D5ZfLhJKf6n+O3U/oOK7zWawp1ap0vhmp
/wRhLUv2w/ZbWQOCGm5xZcz/YbmM5dojubV7lZLgsSK1qhFzYVEQDoM6s4+bnNhBHkinFxwuejx8
Bk0I9SGByeuEKrktXrZm0FeoXHdYUWmt6Xdu51mQAbYda+MR8/GGxe2GjXzh7iNdErXPIdD4VaFs
SMZDobiK1wPkumzPFn7XYDO/IhuvegISvb+MB8zdDdY1JJX+o3oSqBoKbt2DX6YMIlUN+ehjqL83
tnPmPraxcBFEUnrdGXcYVb3RYyVwEhy/K1gNBdzK1hxSzhzCqNCt2F8ryZJfo63Un0Hxw5PeYdvq
VZB7ddTyu342ZYfb2VuwQeK7pZ7DMJ1qpbiXWojaa/41IFrSNvZiVxP0PVv8ir1krOQF1BpT5oyi
gwJIfQDHOnGg6uNZ06B1tGv6hYWkrIhYHQq7gmSSjae/VZ2G8YfBXDlDpupMLFMfmkl0QWhmotfP
uDUXX1+x48oIGV7I5bCCsJuIdUGoPTURDd7nY51Tzc1YbRLhuNjxjOj8ZkQOgqoG54Iyfrouv9kF
VYAhliGYNVOSFZHaghIjRkGifGFKXf/8yh2/hJVjHmlA9tZ5Zudufkh5e7USBAO1zUNvb9loYUfD
rl7j9jBbOcH/p4lyPfdJ7b/RqFAqItM1tfvdG8jRFXjjr27gIYID+W85ifQ9p/+z8OzNNT2z8oNR
suOG+j9xAlQcxTHBiD4NewkgXvl9KMfvl6p1kmVKyn7npXptziGiK/YM1OZWheN9j3i0zNAwl+Ec
vYfRc8wT7DSWDpJ2CPZBeaIPI21QiFKr1FcTkzSbsaR9FiAiCwdU/6yHFGBFsmUhNx9UE0A74nwp
a9NpRhZfDjTpeyocQc1+bIl4a8TzXGDDZEpCjEuD9kYBcf+MTs6feFsdEmNy5MiU8yoMDOWzp13t
8HBOmUTqX6T5h22cNwAdpTPsRmEMH5bJJm5gsqRmaI+qAveah0I704EIYrcMeirS4YBqiHkLncjq
lPy8uoTRwJoaB1JIXsmF3e7c6DUa3kJoEoQkobtnuOqpmFwohhZHj1hoYhZ01VMaVi52jNwL2iop
7S+FnRaDrzVOH1VHHwglD0hZvDxIo+nB0Pr1P5dl5ZrAtA9pDxOshtsBduKnE5DcmIsYcIaVCDNg
x/iEzUtreeqTkphuT6h0CbulvFN/SLv647u9xMoDUCbypsOLUVoCuHd87+Cp7CDYoxZoA8t7gtqC
q/1Iffo7wWKX45Zhc8AVavMz2rFLcrnHde2uiElkytAZfq0FtomiPXRWDCg9TyJfiBFQTdSCTzWu
FJntU0shuPkKinBntc2vKMwWQSQjNF3HA6+G7yNHY3e7LSGSAivlXjuv7pMZFm4SRMjp2hX9WmfX
3S49VNRj/OSeCfjbkgtg0kXDNbeTwXid8DDXAjsrNV11JQyzXHNIPUJFCm/GVHmp1tmgLJY9vrmo
DahoG3OPX458heNCMHGSesfXiVt0xd5pmch/cQ2kOuxBb5jLysel83kEjjt4Sl0CNwWdzFUV8ijz
NQWgdGJnf/qw6pU9w1ttPOrrsc94A7V9t5mA2PMSoRI5ttlMcJua0VdKOUeaem0o0Otl656aGynr
RVH7juuLhIEygLwGa1nv7BYTxRcqDRyReOLjCRO6+1K7evAtbNE/C5yj49WnO5un3nTv3Qa1Ify1
cmZJy/PoOson/EG/V3ugEb2xryBE47CI041144Wcxd40D3Yk4bzEp34mPsjKrdzSM1p8RDQefT0H
tRrP4AVJLSQFnW/O24i7L7lrhR5VCNTJVd+iZmUIgEvtQrqxNyfFz0+rmaYnLvvlKtQUbrfSn19N
qdVn89oVU6fGodOgOrf7wdglPofWMsgrEEe+LCqQPMDdVl2Vy7Nzs0hUBzOxEACnpVFqMAdC9vFV
KJo9dVUkfmWqspETwKwLBA5bkAivflWYRzHk98ML3OkMt9qcTNVFzH6FtSwx1JPf16gt1dRhisLd
yzB1B+p1q6P/94Jo4eAky+dHp3+cTwFgBoFT2mdAPtSIZ6FP7S7ZL1Rb/z6hZeNCOqCHF4CE0vwK
J0e/ACmNosDaWef8QADP7mrKqlr0DV2XDX89jpfuNyT7f0Qsxf9eg08K0qHQeWCntL0HPAQuWe7Z
cr68Phfj028ArcLdvaO2rQ0rLs1ElSqMUx6kwVbWdXGuJf0khDxbJWgAgXM+WHgzwB9/9vhZqXzE
E1bE+hqgqwTHJVG99RVVrd4MDR/tR+40RSMJaX/OSEGillurr4VUHrpqoWM5vaSNoWqdx7HhD5Ql
+jjxpEa9DD8acA/2ckX54V8+A3ASIfdwu0D6CyVLeu77Kq1PS9RYTrFv+xBG/9z3L79HLhQ1e4vx
ONGFziFpwnh4UL3R2eYnd6y8TrWEqvyXYyQSNti+QSTyZsZRuuaTdrW542VAenVPFQ5MxeK5z2ph
yWktzCoRbZ1ZxeIUORmCr4QtYcCULAPgjNv0K6pNWVEaQjByvaWqiTbM29UIJnkJaZXQy0jC35Qr
ubVL+mWIkgnsiT/llN2dbhCCgBI7/rOOnbCzGEBDnhN5iMfsuo+ljDhmnBLqt+DocOHcFrL/DOF2
bxhB9UZStPU8dGoNSk7emhENlUA8ME/I6TnuhTiH+Gdm19bNLPqj59NPM3XoLSN98lTLg2Fvlr0s
746G4AhbZ7jiMZQlfVNNRcGbxHXe0DSPBTIctDpggPWVlT+iiU4c3a1YP3sstFOX/UoEgrtD+wW4
AA+97CZie+Mr5IxCjpbdE+jxPHa+KyBHAy9saY0sQFNXg3KOHVsBZchtM2l58jXgY3nTF9EOQztx
TDyeOVUUHb8z0mqPOQ8EeoZjzA6H3rFlxwOrqC4W5tBDEeW+ktHBIXPDyeUcwH2RYFq+gZpFXFCZ
u7Hw63h2vxnMGxqi3vWYcWeXN4LExMol/bSNsQv0en3Ssd5HFeE7u4XzCg/hFLaTgeUZ8nyCMgv8
bCadL7rODc7ms5nomITnLsLSq/9tIpuh+wRrILrvUnF8/oM10jlZmPCElaMi6Oh/tOrZQ1MXcw1g
O9lxX7iJ7DRGvf1WgaLOgocb58jyRKFozSMCQQoF2CY17myMDCkDMiUYMEWJ3NrNYAyNf8jr325n
7D1XMZPEXPr/2FG6C4k2NIOEBVKxBveBz8n2MWqG1ftKHaRQlUl+Mlxn6G1fQiaWvOLmZQpk6y4f
ZbL+VX1JCYBt4LE5WPt9IxxbwqNC1sYkEp+Z0BPHu43FKDk7CaYjAAueo52r+zvZJ3Xfvefz0v6m
5B+6fkLaWKJltLz77+CpswMy4aS+3i/x9RPPcBqXg2UL0N2Twd+wE0J3O5urlDaBWZ7YCjGGJX4f
N56k5nYIDLRsu+JGHXMFa1NztphVk6NJdrmoSElEthRaDv0F24JgvA5OA0BYlJoHB77nyASLhUdm
bOY/oFs7ieYG1FjSm1yfHtWiDuuGejMvMRWfP2rZXLTjjBhWsmE4eBJVMLmtKCwtzBAxqi5w383p
ZngSLHp3QV8B2+kVFdvK+IfqPE6FBTqyKDY8FfrcvNZHSVDsaUNuJuieKH+2E1PtCCJ/KNgzFzny
uTu9CjLuvfQmAbugdSUwG1MmKG4y6kYHJpnVGZsyA03gY7Bect9x0o4YqJLwrwY4kNgvFQm1COQG
3IJLroXwf2Zfio2LuzBBNN/R6h0ygYIwzvzw+ELbfxsP+8IgzNGPf4cLXGK1Uq/ji0oMIYg7+UvN
ydtt1/LT+8dQySkgq/sctIKREhtOEbY+8DzZTMADvtNrZKcGBF2DSEMZpyZr5l4wa0IX+K6lOwM8
5rvZbJ1nEkSHrusD0gVCDMbZYvx+9/8227tRT41tfteUNOanblaYVbL1V0BgCyWalH0OvKJ2UmOR
SoIfCvF8mk656EK3T344xX1F5KZnpVfhsZySzBYjDmEHLOo4lTu8lsnH0t7na+zr1g2SNpGgYYx+
k6HnojWTKch3IULKKQLt33iR91q/QuP2UeDHCTOKdh6QRYv+AZo8pe0cLhjGOj1yOkY0+lIYG3KQ
5hc5HHEqVF0zKvJLFKhW8P8H+FaCC34Fu7s4a2Km/Mz7fSR9HAUJsF0iBtQe/+vWOOwup1oTfhIz
u6hPR5LRGnDJ73yMAQWb0w+njGoWo0fmaw9sLS4XknmqUOesIukxc/YJ2CD5ZnYPk0kadnOyTBuc
ugRx6/uA289Ee1Qcxi+rh8CWIy+aVbLGWrmng7Is75M7giSvADZYCUUIGpL9lgsizHH98r2mnAS4
Jw+F9CR9aJZmldtr4FwLbIS9KM9GA433Jgt2QsMyejvO9eaiK9lsNTI4NJSNdpGYZolhUn1wocA/
y3BlG004AOSv6yRW7VqEEheL1DyfSj7ghhCXZmHaMRvBdORyGlUCFbx/YhFuAUVCzfWVfPZ8Gtan
pYsSUKoqZ+zaKfH0OyVGVtRY6gLNoB9ez+wR/fkWUJOa9WSaq6jtxGy9oMvbpgYY0KC5ZdrjOONQ
NwlvTAjeuHbeDgG6lCtqZRFvRibd8n6/apMa0DcU9/Gdq6+0zXOh2XIi5gz8YZy3LT4ihIVHkvX1
tiRRkL4DhXHDJ6U0CADmAL3mmyemt+IFntYBF+ptN7xcI2vGhpXSzpLWrvpIsB9SzVlvOSjlOwLY
eLB8p9y8Hwfd99FgwUZI0kGeXRHRlMoFiNStZbFOilAu4lPNBeDh9lNUKxBu+1uJq6PI0RI3Nidn
0vd5Iuf23Wxbgzl/IBC0+cSdmF2N3mSYe+S0eHGT8ZdNT33F0XEFtjrcbzOqpl2CqXzE7k52TPVi
AIHFxrFdeUG8PCxpVfQEpw0DBtCzVoThC4HBCiMbB/cns4RinMC3tNR1zNRP5g5xgzQfS5rRu4tN
ys45xs49Oid5JrU6iUO5wfaeGFCGF3K+eAWdjgu3cj/39Oc9QtCXsAtlS0hlZh/q5k8++q3n7yJl
XeK2CF0IZ9gWhBgByoWgqz69oZMFPg7VamgwOnz1FkqvplHvlkhx82Jw1UNe2AJqbBF5JwB6KVVh
zd9lMzd0uWHxVuxHL/Ef4/Yp8/OJCIReKU5NhaPKfue2gW4VhkVrPeXQro2dsaZTikkr4BhntORo
/pW9c5bOFGpLCDlmNmoqgBX92VcE21fJIDz1IAhgvpKpnzutIFMDXYITtwZudoJw/q9dtu7A3GQZ
e52B/e2mPJXYY1kzq5EuhqaJR9sxLUAMDjNSo/8MswnoK+X7xPRd2nFKVHtarGfhqrchqIhM6u2n
3OGhuKLpL+tvp3pP/J3DlVfNTTXo4ZT2mSuXwCVTYadcSu/9zOLHOr98KpNDZFwBzCIt0E1/htOR
WIdHdcBnjWNFxIcFaVggMhBv8vDiufFwrs5wq9jDkF9iMCfd0Vs2DUo4vJnvMAGDb8xr7GQJ52h6
q7vEQQflvIKfaAwkDdw5Lyi4+UTanvkquttBHRJiW1uOMRwnQu4N2L0fdd6RQJyQovgZPIMX26tb
G65xqNizpalbR3urKBcYviKlsiirNWOjzdcYvbicghWHDMUFyKMlP0yczhen+rGamomNZ/om+UhD
AwxuPUFUr01j+I/qSNYOylkX+HzFW6XAO5cidlEhgkUU5bxDdZUk5FWdM94CZtkeEUAnV7HvXGPW
JdkAqi7AYbw4/R+1YzAJnXGTzWgbia7hmVcTDzZrjiD1WGvWSnSo7xksV+Smfi+OD/bQLc5eYVCC
I4pF3XkhB2vH3keEYh0vqkxZwUysCVhi4lT/N20wqyX7YeTOk0PN84rsArBimVOEAEvQ/CTAZ3CW
ap0PKgqqjKuWeoUYgbiqPp30HCdr3UvinyZlgilR22x3pTgdFDlR4FfxSa3szghA94lcJ2vPuEPL
npqMJdiu2a5s2DH44ZA9UWSoBIwShszJD0AlqR3VbaUxm9hEitH/3BK35+69hxngcnsSxTJJjyu0
isBFrA1d0m3l4+UVZotbrgWh3z8sti+8irHzr+M9EOc1dXXmFDFwYjGwYM1mZ/6tQwZHNaXtYSVX
1Y+DjMaWmALHVVsNi0cXQ2qFOHJ+bFaGOoZxs7DYPmZDdjVKcf5LZKPTKPc4yQQLc3xtiXWH8t3V
uYESYMlFMcwAXvfW9AUt416S3WKHNg/LmgNO6E2r5I2fiY1h7JJ/vOckZiZVF+fYONjiALkKRIRH
WXm9wIRUTuS7PnAnvfWRkM5BNPwtyu/GFjH1F2eXLLK/9Pa91YDSRJGe3iuoo3FHNaWLfu9aG/lb
7Gx0sH9COCywFmgagdQFNrDAmdU+2dOLfeUIFGZbNp/gnMHD+EnJmeO4OTDU5JYXv+2wuCDTrdqb
ro0EjEos31YubbwHYfLkebqofrFD4xVamm3cEW8IHEgEHwGKtzBCBiHzs3m77U+p3lA0pBKxog4H
LYtCllMSpZx4fu5m+hOJsqxzb6TAD8P2y+FKWCAufTj057cAtISH2Q/3onBq+3ucDpLqoYi6pesf
HTTEKBc829MnsWYQo1n4xpUGB80sHs2gEb5GSCgGQFBwLDBeZ8G+YgQlCfRvlLUufkUxvKPbu353
t4/fxj2pbrIGwjheSOjsZkQfsrxi8UwRNomHFoTQUNFCKAjT6FsnbzKE1E1XCvWtLCXL1fNBOBii
1zoETLan8f1yJfl4oKmgnr79nAZ+B8PdsSGdHeLbt1kSZQScleYf8XWJKnRvzZonXm4/gzKngOyd
J6+jbwkJAd4wEAGMCwMLHcbiZvn9Xjj6nOvsZllqaDYfv/K/3dkSAa4I9C2aMGTUNNNWdN9mKUOM
OgD5c6UahEdgT+XJrfPZdFmK7nCCLpzy0ara7mNb25vhT9/6KyALxJiAZPuy3KAtUiroXCcmV/dR
htH4tk8KeUXVrdrgYv8tL3gVI4VqMOZ739jWPThYQ56eC7hHcL4MTUZnfRJ0ftkFK+koCWz3hV+L
xyL1/vBXjzQ4QrkUTmoYMasSkZeP1WM+o73qNYlvBFHlihRpgfsRn3FdIxTSxtTy/nqSG6pphtqY
prfhXd57/7UlYgrp1RdDzyFa4I8aHf25X5Hg5alLr3TTxN2VQg7kBfmFXW+5wCk4PJn4bazQhgVM
jflAZiXBPaz5r3ASLgE6xqon24wQdc0ea1qRTcZ5tS07/MGnBIZO4psRHJ8GOUhV5YH69bqH0Pv2
02X4/mDRTyLdo10F5qRTe2YL5aX2mPivNFOsvidVsoGQRPPm6HwZTuIje/Um6uuK/zwTNsJPl7Tk
sAyV0esFn2zjbMlBuV7EBaqEZToxkr1WFG9OVDjO5CBvMJcTjsQl7TxyUgJvrSJ0DS5+bHWMyMmO
QZb2j97spwrDYbySOzn/xfZ8wKh/1RmgsjV8ooc9mrzaub7wPrKlr2Z1f8b0rP0s4I8+CuNa2qdH
t9Ts0tRHkuEY/XfhlwWmbvWpIreeCfYiOM4LJAK7LGiQt9ojLKCFPst+zICridKt4Vxaihmwirq1
CMG3iow3t7rZIdTf1ne5U9vOhSzyIo/jpwMcROBhAYBP8vCIDXLYMjEyUNa3mOLBxuDy8NLbk10I
lls87vWy0DawUChmmQJOuPeATEpCHbUAkPhW07ZoGDIHxDT/DNgqwFwewcGjaDvR+vFrToJj0mD+
1D4yd4N+0sR1UVZ4ztHm7fqFMq8oOUuJ88miF/55sqfp/1jU0gxUkjGNdC1en/2T4BIP7FKw3J7/
AXKlyWIL1lN6ILrJbFqz2mmoeGPhJykyRw1KaFZ88XzH5z2m8EAHP37++3uAhmVRFb5VABDq5Z/R
l2/cpMPaMLu4AyW2MKMF7P142nRRSOjQnWtDgbScBceGDv9WT/idF29kMyRwJKiwdUAW5MJtiIay
5niunbIsQ+Oun7Ya6q2wmFKmo15iwi0I44V0oQdjNeTK90FiyAqUzTVLRMCaMYdHrdJ6tMmN7/II
GaHIIOOpVm0oBpfeo7EVWT1ogbBQzkiqDRDEg21V/v2mOuP5VpBm0t698f8b8aUx/INu4TK+ESC4
UnG3myC8xFxw4hMndD8egLAFDPabp/BqFvqK7ex78mfGBUMGsYCdvVP9UJ6S05Gk81kgH6lA3vZ/
XeuWM0yfe3tkyZLJH5JdqL7oIVQAt1zloHhbT0BsCCwJ21BVOVm3gxLFKBwup4J64EJSOZ1hT3JJ
2w6S9M3s4eSmQAwOEWkpzDj9Px3vXn835BIm7SFU5Wg9l5thCneKWDtQQAsWdP1MFifGHsPZUVi2
FKbUAE5Aav/Heb1BEfYvpwZMABXiamc3ciJC2BxsiUXcvewClDrummBWmyS/vRwuJ/7VeOJO9ALR
FMTae+cNrRsXRhyaRtOPwgbSc2NWvcLSaQCTvv0O+PoN2E9jFOwP4OjFWsMfkBrvQZ2BxcZLZdjf
W5dAh8JckjAlpl8YduM9nMEbW1L5LTNNfUIySe2xcY6YDCV9omGppfkTzn62kWAzrGFOhCj12fgv
zIv5B8/IBseiDhL9Y8Z14XWgV32GkXZ2Mzmha/VNeAkVT2UE3bgabllKvsKIeZhtJWhodMJkElqO
v8+4VBsRnqF2UBAAWUv4RaQkM5/tgKrhOe+uWcKOydJt54QdDQMKy+5z0tkmrW1Jpk9qCcLw51Pu
LvyjAHDdnMHES/J+5ue35AK3j6KbY5E+BVeDw7FFtWOSNlfP0fMcv2L9zviXwH/xptTtpxPh5+IN
VcaYK766v/MEZ/sh+VUiKWMQijD/gt7jB/h6rwQKTY0xmA0LkffRyVJBBwxQwYrlTtYb5hVuoysd
dTtx350IsG8CvLsj+rQt28REFU38jniIGdsbF+iEmIFrFSz1q5rK24P/ZNv8PG+viBd10chregRM
rQQZkJX4PFyEROs5ZwiU1ZqRDCc27MNEritFZwvWeoFEhqo8jg3BNxhtI2SQfzMeK6iNfu22WXfG
+i9958/8KuAkUxAsCiZxBAc5vK7H64Rf6AmIpiWYLNDcS87xU+ifHy4YOM1J1Gug690DxwUqE9v0
o3g2YgvfWqdUkcvnx80/ADZ5UHnCtOzj4DvQF+4ZWtMZp/M0IAZCzUKfpg+ppS8h4Pjy+SKuATr8
r+Jm3BsrqRolj2SQxuqRhWiMg+RDp86dnjSffoAgKP1UmsXCp9LtDTluR6H4BCTB4GrUiBQI3hEA
Ig9tSv3QoYwnBrqozVinpBIEga0Kb5G5JBTKEAt165TYYqYHlZg5SriO18UwKAwC0ivnlqz5SITV
epzBJ/kNroPBiJtV1J3iykhassp/7j9NSXoARR9l4bMHQjDwlgLqlUfeEYtsWJ8ZtxcMUAkwHV4m
4GYriFlDrD65M8yhCVrudcOh+zx3NhsGKOo3fhja3VCFQXsJi2pprdjsO9pTTNwaWAqVn0w+qzrl
/d83lRMJ9RUepGypIVvXkDAU/ELZVlp76L/uekvJrZ7mnWH8dGbVYMttqqQYRSYuPOZTAtocVYUN
xaLX/OQ6o3fGJbX/5Xv/KWFtvAOg7/XQW0JmwA8dsUhEnbDbEvfHlEsthefbF2f3c5y9YtAGhqHD
8BvKOxx1+kQ8cxSYRFJjtTFKNla20ARWnqe01HD/7Cq3iZZtv2A+oDpq7/WJ7QmmZfJzU71TeXPS
bjQEIzbRalEoNFU5JndeY6umOPfWU4XAyxAywUjsGqTzAGSlb1TC7yZB3uWrJD9SwiEdG/x5S214
fHIuC1nXsdsC2IJUXXQE3pJZDaRLqrNvPN1UDDGYS/eSbOD2JxoEbst3+Zy7ONDiTEwBzLHZeCB7
xADXSi8EGwAzqW842fB3pT4VYnJsB8CmyO1gLUXJSsXM6Q4j1L2zXSKj/TOzZ/4xeJc+zJ/bbYdg
8JRxghhAJqcKfCXsnETGKSHnI3LnODyvGFkSK4uG73/yr2+Re3OkBJrG8ExUx/B+srkORthYMrt/
2nq7Xzw6ST10LFMMHbGbxfL5vfJ4GzO/gNWk1M8rd5zqhY7ALQWToXW4iOj/06OsAeZVYrJor27l
A/DDG8AeezZNr2T0jDYbEJh3eFFsw+bGizaGsId/nk1sVjDvnjoCkpbrcaxvL65HTYq7CjP+537a
AGQVFhyCxNjKQHvmesg2AH1Wg9sT/NI1by159TwMu42Wty++UPoFRJuJJG7uzjfoa0E4DA0tgOs+
Q2CxX4kFfU9rT7++OWcrXOLekmANpgst/GnG9Z8KGyYqqNNSmEbuNc7aSb6LY/WADvtiXqCiH5r8
4zla//SjFlnfxsrCQPLzdjIY4A/35oZKMwhju8dWuqEs4rfbjvjZVKY1nPmUUwzbUGScsg/+3pns
ftNMn6k9NjHblO4VqI3vkpSgUcoKIQ36IiCr7e2V7mf2W9M2XMYrVRhyvOTBNvYnq+nbVVPVlA3T
TMzXQUbXU0nPAGVkS/LcFoBK3Ybcsa8wOTFmmeC6xVjFeJ2uiOyvyt1Z4wsmtZ4KeAqQeu/m7ZFj
qSZszT6c51w0y6HN8LBaESZXLNCPm1ERp3y+gTBCFDO5xcfKnsuHyeFOoWIYCi+alAqWJ2+S5Tb2
2E8XGQbqLmb80ExvHVdc1uRIK/7X4ffRBnfEpcjblXI1qKaHGRgkD1G9TbunBOb5gah/ximdt+GM
qJag915FmyG1ShTur4EfxNJjcLjcikApGzJdSZZyBjJh0Lc3ckM9WcsRTVM0NXCEctmRBxUpvAsj
KfeQmJJDhWu7vu+MqT1ZHUcDvI5ZUYvF0NysJCg6DQW67itrJG5PwLqhdlegMxXH7WuqPZr2gaLh
tUOvAJ8ApCD2WBS7/ImCnmxMK2B8jOAI2HGd3Nxm0Sv2lBqXhWnFE3Iond4bpei788lvOdDiK067
F2ajG45ecPHTfxHo+pfwoOX6u+JHxoMDBeUru3926fDXD6ryLm6Z+DkzuRRnMwCuXYNLVI2HXc13
npCkqsoTRSTRLHKPRT7IULwSuIsGmkl9yc3WLv9i1a8pa+k792ulQX2lbfrS0/9x91ppU5X95P5L
Vw0Vv560mG0ZkSyZ2G7dbjWTZP1IfX6E/ByWh9S3DpBUzplOeoSogSO3wLEpgXj/s3WN2TqhEo7G
CzVn6tBuVLJ5R+V2kKeAzt6PtRZ79WpaIgxAgjkmFgMIjmXjvqJZS5uJ96i4gIeyW8bq8w==
`protect end_protected

