

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gqDFw5NFAM6CTSTQpb6ewV0dkTDze+wC3QoGAxwxbjcNW9/DsOht+2F009+7g6jE2OnhGLtqTq+c
HspFg2GBAA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OROCzcjj1wgCYlIqlabkGZopoXwccuhDPoDiFwbBlsbzl7flKX8tC5m+07o0XejIs9tQT70vCTz8
eor9UB573WqZyEwu6nS7RfReZTn9rXIEfFTmb5LNQYR53WQufFJWXVGGzbi12Azu0TUMNBykYjra
GCJvYkOLjulS+N02/QU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y306+4wGPVAAsHa7Tcr0Z+Y/dNy6G34dYeGbx7ATqkdiT3xoZwFMriTbyxCB/BNDpEEpWtR2x6B5
1geIXl7xRsYW2a/OzYZ1VgC14cIMMrlyvjd+Q0oeBhNwIf7zzOU0YeLe10Ln0VhNNlM9hG1yxJpm
PklN0o7dbe4z3qSMhzdrqG9CNO1AfE0zEYRDe4xK7ci9EcGBPeIBnjhSSGUwaUeKV6BzeVeTBH5k
pFfAdDfvgi3P1VwvurSSAL/VyrhWR7M2OhP7fekXRqEU99K00pFciI0NAEcJPUl8pbYtjc86ccu3
OmuQ0fZKcUeaRlPX6glqeiiehMLm/EPWzCdMgg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gSn/ibMO73s4UyV+DQBAOvPjnov0A3ONpbzDn5S1gDHbJc8laliw/uAOvABs0KKAN8Q7GKr5UYxh
qWYO6FhJPBG8V6RCU+sAaoeSnleJb/buC83HgJws4chUKE1EbA08UnkA2E57wCSfAlSkdEQl5xrl
E4NsCY7zrBmnjMH1Xu4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lI1FhNfWvnI088CMtuEIyHMeXPGNhtlppeaUXaQvRzrpC6F1bRvO696fznybaYq7K8VPJB0YyXVb
8oCJzTtV2jMI6KoF+McAzbvubpz0ru0XOCjjvcTsZJ3kGxHGUlKh6xdlB0Gez6kASJJe4GeTuEaI
VZNg+Q6ea8OLPKgQf7VICmBv1vM4svyVLDI/pSGiGOmfSMrfWDP60zo6tHpkaDS7uHEj2WN7lXT+
Q8c1SGnQvLeKyHV/kGG66fpNSvILAslBR0l5Xt1/csaBtahK2IV70dxaZkLZ2c3pylf+SxXTt7v2
CzVvxEgWwmwKjiuhBgmVM6qeL7+tokO6P+FlQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 41056)
`protect data_block
qz0aGLCwb9OfDd6oMobdXUo9F2VRX/hyg2LYvLNPjuA9vxsm2uEuyLWX9rMobYjC5VvjzJ8+FDMw
pjAAUWuf41U2vz1t/LHkeV5C0eTIg2zp2gvNl+9gM1yWcxvj3Ays4ZnJEWgY6DKqh+hxeBAvH80N
u+fsHjuhVOGm7rFv3ukQzNA4x1ymuMtCaT+FZoT50+69ZeeunBhBug4HrSCxrnYupM2eAvoDm7Cs
a9zf9EqEGJz/223draf3hf2Tfnn0NApUEDu/GNosBXfeEdBKh0HSCOH0fQmcutf5Tj/Ao0MxJvre
atyySgEd4SStS2IHgU8rHfPogxaf9rDLtGFbeWUX7amD54XLRnjUcE5U5VN1M0TX2bLdOCVUiKzy
YqkJTO8dre9b9H+wKNihwvpMnz1TMRnTmHoRkrEiFkWzh738NaB5YLLoomN43q8k4SAFYowDCTDh
yONR0uz5Y4NIIX3qfE+vusD8mtwa5XFl/k01xkRO4pEmVkitpo5eOB9tyUgsgRySctwnzLpo5Mpz
6jhPkExYei3CFQMu4hxHUzMVzLAnIIYBvRpNw26hFLMJDqUKexc2xwyA3uFaAZ0udRXGpLnRaSRh
+3D55HszPtadjmLb2bxngSTQgIJbxgUFcuKXIHAFA+nYOrHk2SLsNs/V/k5jExK1tCObqnjoE6YR
6p0MoEMdLPC9r5SP3HebQNSGK1rgHpIYedYQjN7sJoX+ytHWJePCJ4g6uaOu2/fbf1Fn05vIn9bG
uHFhOvRaFONjmyyCKlpNkpFf6DKxZgQCp1OhiC4CsKXSaih+YH5yTUJ3eWd/0LrNxTeia2wj3qg4
ncSJ0d/NViZRjF9wCBxpr9uUEnIbk0kXPBKKu97HOq3vXV7VB7sHxZWAjW03FMqsaCz9ZJTD+yL+
LMohQ4+xPVBqZm4FrNwynTpt0OfB0KKaA52Z/5DwgHoHqltth0H4yX9P7FivJYN486KMTo27gQXX
vqNadQbRucazjK7FpOPFEnIVsJZzW8FjsfJL74AzYrZRxalIIMVVI+uGJaKxgnoty6New5m//hoO
f0RK8Xu9kwDgKBvvf4xy6yDKnPMnB2MZWOxadWT057vBeUXWclBoU2CoNpL7JSFUvgGKiHY2gnzD
uBzlHTRMTvyWbfGpz6Du7etSY0kLqzgZrcMPlalapS2kQeQ3dtsDnlBBnglgF1LzfJS3D4LjB6Hf
5s2e0vqZJ6iADEon03UTzHk8E0ibK1F0n6qblLEha/cNb9alnI/p0y+r026PoxZegbidK/RTu28L
oniDouyRF/iq72zR/dumxoLMTlceVIGbl1RYO/CnXJn5hFgaPS1QaxQ1FoMGmlthGVy1CxA548ro
CGkC8chKxuWWbSke00gsRRHhPABamQJjXV3p1Rq6fBFhH94SboKK1f+BF1K+eHg2QGRFfzcOU692
md8A3/zsJdVftwDEqT7Ut16awOfjHZk0oAc7wPB7BXwLnZ3UdYhfNof+0fyO0FjjxH0RPclT3U4V
b6KH2ALCMsKIcLIwKP1Fn6zVZhEQ6GZB1n0RSx37OBE/NGa+7u5UjRTD+cLi53go1IAS4GlXKW3b
dTFILKcDB8J5UTYx1XLSjCL5T3466nxFnCU+OY3ByvL52Dl1miLutwosAxMLBcGX5WMJcHlwgQJr
iqOK666fGwKFvrkPeznMRPsnWVuwmLKWC5QvW219CoaCRJfh1OLRKg0YrsjKAatE0jzfXHX1iixb
W+ufUw7zzbeQErUPp6Ny0A7kQ7c8mTYJdIfuIl8uSlzXn14agRtxgt4x0POQHZwe1QllLiCwoAx3
O9eynlwg/WBC1R3UUGbpP4stvq22Ry24pBoGurQK2h77xSE0Hb5Zlqjp1IkCron4/CHfaymXSF93
Wk/sjGIwmAseTugEgnZVpb4Nt1Ev/JHUhrohX2glPvbSiGV4qHcgQcMejPUfVu4o2PFu2k5mOJqW
9AnSGuhh0CwLWv9LxiC4yhXz05TWp8I8bfPRiVgSOvEkdpmAP0GkaiSl/vswQpCIEG0Fbrbupcq4
AoEmqEAUdrbdjO4lnF8QjhGTHne1sazGpC/bc3cY8Wo7Z+cKR2PxlqPYuZOk54ukyg/MclLd4ADc
4GKi+mfTal5SZA6IaIzZYA8c7bTJzqGjTCK/tN59q4bb0EeTHfkx8+xG+4jJ89YQtNr+EEbWbOYt
0VHFtdVkqS9CPY+gw7X3TbhpcCt5v8MR/50rCh/tA3HkOafH+7YQqHTmhtAhd+PJ0dRgUJV2WoXo
w3zeFZ0OuvN8k1uKTzFe+w4vqkwiTAVPsVyr0rt3ZcMdrLWx53Siha8dih4JDjEDPAP+oAXLrsIx
7uG51C5gTvgStPg7Nbm4EeYX1SRoRnMGlVlacNTPG/YmYVMIWXt0oTpScJaIkLvEJ5yXfpReROXc
GR1haHJDbcGGQls89ln97QD6JUvCBuBlh+7U1hHgJgF89/s3gRRT5MQgzvZgiVq4Cymsy2dNO80r
zsvUqMnuI6Wus3/Bja2R4XBN3n6pDsYM0FLFrIjPDSwhO/CXUw5BwGwxXdpc8/wsK8Sn/GL2NGzW
ZgLe8K7HkISLT6IMOEWnDSLGUOLnC7KulpXWub64a+ByiVU77eMX0lYlRWuU+Y4D9BGTI5HuErLI
MrtdxKLySyxXH4djpYppHhazvxtuIa82yeU+QKfNhzuTpE37/8rGAmWQiJStdyi4Asqnn2GfxHWK
UBhHxcYnmVMnMJqNzbendkMSIlztfxC6JnmDKmryb5IeJtkoCkoTnlBXntMTtcU+fYe8lmnso71H
RBcMR8d7v5syR2k28u0ftVYE7DG2BfgUY1IcmM7vECdD9QouuASHwHOEL9Lf3JxJmGiIdXBllxvR
6vxzL/tu4kuHyy45CklkC+B1QizHTOdrqCDMPCD32vOBWeNNAIMaCmPOiIuYvp88Yziy8+noW2OU
IWou6eU/BrNrC+ElHDQC8eeEbzWVZVWGRuJn4meDxIpHwf9Luz9Im1Nj0Ol/E3suZ2HfhRWw1Vmf
uaFHgEjxx6n031WkxudQR/DZmEpM+VDBj2B3L/7R+Hw4dYGzW8ywh3HLfmpxGcs1KNwaJJhQM2/l
qHsp1C9vSxs3DW6DLU83yLJc8JuWu66IgC5PqToYh4ar3/VamGjdDZkz2pnhS8G/Fim3ozcFoGJi
y2pOdtYwXRgI0GNj1/seNb14EX0SBJGD9s81tqtddcF6a+1F5bevHhttCjAjViuz4EG66QKORPNO
UOMoXMjnFgA2HFtSrGIg20IwOR8ddnjE32V6vxZzU7955IT/fek+UHWVQWAjx/s9TvSby0eq8Vwu
bqjXOrj8CRB+GA47lE6wLh4h4VcjLtSTyQcPZg2xRtO0hGPTC49RDm/eCS2DGe5lJJo9RyWcM3Ng
L4S/6yTdaCi7iM6wakaziWsfta6xtBRqJfsE1nRVJT+wH6AP69N8V/YEYNUTziMF5RpO4+dJ/OvI
FP8Cj6oqnMpZnOHjdjZFHMWd8V+OoLIailtqR1MDbTglJCIxaRrVpo2CvKI4AlvOQ7lTMfaCzs8A
+8MQXmilXKbGr88EOpg9QzZoM+EI0D765v3x+yzrt0OkseYIVBIqycFsHkNShTFu3PdOxNeSJL8R
0PlGJR1C443k92dhmicVUGi3UO2FtHnHSPVaTNL09eZtT1GvUvOcgRUyc+DP1UIymv+5TM1hCvJC
5GMZjvr2ua7Q5SZKxvSsBiajjoSo7Nb2/iwgSd8JhO9P05SnTzyKGfbzoP+aiXMUPtgHjl0cGCuq
9+R7fLWavip/qcUPhpQH8HvcBoa8g/kSXJ7UO9JHleKYNFr0na/p2AiVhUVtEYSmZ98vQJAmuTI2
nQui/HTEe7TuQH2ADLhaa/xqmNOJ3m5qvMw4s04npemFTM7OiIIaQXxr2xSQpOXm7XwHPRb8oCqf
YG5WtUTfbiwksAJykdGbdT0F5JsIydz9ChNh9P876Y9/1UfEivHZ/aOYAj3VitBXH3qQwPSq71BW
ZzQyC4UASGHfL2JdHWjYEj+AKDIgag5CDvPLN+YhwB7MQlNlHMQ6u/P5jnT7sdX2KLXK/RCrHzJr
iazv2nL4WIOXhSrmqHbPhz16dRhwoGEol8R6eiveWw4nW0tFUlHTasfZvLxHb08ri1WBucgkAofZ
TLUyEJB1KheZoiVhpafQqaCrPxFsal/86Ephr4E5NDl3grSBeU9bCZYUoJyqz3qsx4Rpt+FIIyVK
dZiDahela7sjwBavMZUZomy1fIY+bMk+8V+UYi40Mra8qUWmDDlGl+xfaFR+mZR67NKzywkJaqct
ifd97KbJ3UUbtBIOGA6gdcbAYXplMIB7OBnis5UMa21Dz6aD+cquKWbcTjRRYH6Kd7ULTxtD/hm4
Ws7f/KLVv2uxEdymORSWpomp1s7+OOnDupncd2wpWad4NRQ7YTv1WEfAN0TqKZj2t/C5CxuIP2Qu
d2ovAZRcjDsY9olQZ9pfxr+gfLCAzrTI6/lGZddAVU3BL0kno6N2sT+q+7FwDjKkl0w+TBcVySyr
t9KHLHxIZgFMInHeFDR3sKvpaGZgCQ7vwCg3ofyhPYXoSJ2/qQ78PwX4avLr5EO7tKIcD1SDCTz/
W8bgJCWT/NE2kU33hP1zXUKmgVkMBPpK3omOS8EMl3BztSKv57OLWj5fRUwOo1Anf5S+E8uHss0s
JX0d17fRAUaLcafQYxVtmlmGfqh5JosIK4PGZry5Jb0H4AV2ylplVjSZ2QUE1NPDXccvI1B7Tr+q
SOQpIQ3fcr/b/wl/EyvB+dfjzcTTNt+g19k4uupZNvw/AQBwHz//EkaNtXBWQEijNsbB+t+SB9s+
tq5dg79A+AFqpzQlaJbz6I205sBOJXH3cZq5lty8KZKMIGmVXuOTRvvr9n2+Jpu6HKA05oF5Bpzd
JvoMgzQJnaqaznC996L1zMWP9wYJeY+dbVcAhpOPqQn+MlVrPz40JqNeY98jOC7ZrjWAp/xv0hEX
EsJN427S6lIKKEY4vmR5NOPEphyomp8KyUSjGyj1ViGDsml6bgb7uDWC4V5WvrxXJPMUmBr7NxH0
E6W/dlZWQuGvhuZzgkBKOGzVpK4i9tbOVUdM28itJJvGOKfwfto4uWcxlrm+ZwVTCIb+g64Ztjwa
bkcAPwT1lD9QrniRPRcixe3Mpdc77Xatc9+vbDa9zNZtxBFE3tmLK7NT7B8OKTOFlY4PY2cCr90G
dcUW2q6RWgu7bwvyeUPM1Vkj+J+xY4oeEa5Z5WZAcdIBZGiS8Ud+/nDl+6ygZxY7JTU6ZS7T7R1l
1zfCdMos4srMdU0TKq9c7Z2C1AhhEVVaChPcKJpuw0OOfAMjzyKEQZShKyEqpybJoduO7+GPIwEU
y36m5ZcfZuJSw4EvrY5u+JPYlvKf9qQTDbD4xU9Vh+ZIf5z7l+2bqshSha3X9nIY1v8keYYFmPMa
i0hGbnwmzhi9lDf7W+Pvu8TDfy6BYFU8PlhSBRg7AbIo5Jx8H3iN16n3J2jQdFYViAnsZrCJf2JT
Bcw1UWyXuL5pBef4kDsDSHKPpd7CuIr7SOY9eRkrI9i4aup/Xoms5vL41LO/gJSjz5E/IIkXbayH
fx880UBCHUk0id9usL7PjgUiettC5mEOr8ZOx28RwpDXc72Ax03/yXhtpw368HBcZVljfL3uTHKL
oA69h4ohteglWK54U5RI0dNDWOc2Gufv+5thiiqPGRhFx4ILoqwK63MBAQO8Jmix7bJHFkpY4SiP
jSph5Jkf74qr2KKFPMJTKujUK/Gtx47AIDWDudvIWPBuQi02BxYO6ko3NOy1s4oyRfGZWm9l/z6R
BRFykYE8Zvmm0Ggx+amQUohtS6KMHjOEX31ZR3SeuV/WZ1FdaBr4qIYT3gnVumj8z1C3WUomhWc4
ZrkuTWLS7qf1CAHSsOtFdswL6/labyOZ5aolNl6VWcaW80HjPAPt2Dx0pGqhzDFKp87vHTw9IgSf
CSUXxgTEpt+dOJiA9mxr5uXrqa2QUN9gF3s3mwHzo9mDH1Iw+IubZ0R6mSQwcQ8uil5j4AI+aKcO
btvve8wruvtjMTcZUfFRdkOHtOS6soPfyejtEH0wrEsXKAeSB61ckS7Yoki4lDYu3WMeqHUC2MVs
+IIOd/R3XX1zKF9bIu/J+xAI7WUtLMa/yvpdzerKhHxpJ8L6b2F4gSCn9SpCb4OwT0KrxZ3YA9By
22XmaebfaAfFnOqEJ3NWUtB/DW9vHU6JnhZt3zGvC9YglS3DDH9iY0+7rXfIHOpIcWeKHtYan8Va
9jT5dpuN7hEd4JpHFs5NFFxbpF+av0uv1d20Jkn4cqhSMu1Y3v0oehBX1NpE3OtD8wF9cPegiNIK
EFTz1wqyWXNuhyLUmBykIBj2VU6xGl8DuE58x/GkKR5jDBiBmoh/jDtflKj0a3w0Vlkl2qlGn7Dr
7y7WMcqpgdocafRs4/8z101WHqdHdFlli+x7JzY79ouiw78lnvOM3ywHiEWh3T68yCmQNx0ra02z
2iH6MmfCHJlBzbcbvJtCvNQGElyTXovCbpGZWKq6d49XqMXhrFcCuu0jpN7Uj8Ddj8zMCaIPLh22
4jebHYV03BKeJVwJQh01zCzlB3xiY26F9d2cUQ6+0lWyJcpAPfR2SEyLZFJOQXDJPjP58Yag6shY
eOXGarZ4LC+Ssfe1fLci9vWyxCiQbmH1lx2aBF56tHmJQkuzLYg0Vm0wdGf0QCNEK8dQ2e7fTvaK
nf8cEUF3TecsUhTtiYzrl/kjB9f+0yqxoCm/9w5i2dQgw9Vn9zkrVzp69sjznDqMV2PIV0YNdp8s
7ZHCVfVsBAN2Uo8MuSg0HkmE0mNjs132W177UghXcfuXIS/fOrkBn5pLwtwb1PrO2Hgx3Cvdgkau
eaWs7zCS6RFbXVAm3ZlEqGPoiIrYa4R1C3Saaogpbl969e8Y4Al25VaZaSp5RXy39+HXtxTHj3LN
aRu3PI7yXnzFBMFJ5f2LgQuT8BiJWU9YjeawovD+9E9p1GhfGu4N376hP51bMl8x6qF84xJXU7d5
Aovc53M00yHM6omiQ1cJTMR8yKMoSfocD6U6Ho1lRpRq8v+2fkSCNgPiLFEPpOeljqLMx/hjvd8o
6KLByxLTI6SwZwZKWDXq4+zBNhveyf1/ID5C3t03SokTRCKrHuZlF5Wj9V8hMZQvvs5se3/Ssxa7
zDbjxAL4bzjfaYLojvGZMzZ/VVcRW5kpOLG9XjZHWi42twth+2jCZG2HdTMYWyqhPuSiBK2cHdB4
UMG/cdGY2YOJLpno8PYBxhRNsrGUT2hy8ku4frmT78cAG3eD5fkZofJ8/adHlH91ASb9W6xRjbsx
HXapXtmhipYDxBqLN6v75O9alNhUnuPjb9ZN9pYf2X3YRJ2dfeL6gvam1UsvBI4rgmue/IWe6ISV
XXr96jriocyG9RBswDOFeMNNSl5MqUcg7SDCYJORvrqhjn4UqMn9S4WRnwyomHyP50SreQszuK5A
smL81ELZWhwLCblWPBiYBSaPt13wwVemXwg8n5zJspp0d9e3M4AqXp0i4v1QDOPvQkGxdLsRGEtz
uQXhUTTReCEsEDAbOBKNV57e8+uzi7flBFYxt/6o88pin6e0Jbu5U75LvCjHji6XwqYavbJGfvOa
w1iPtQG76PLDjwvg7Y/p4lJX0sqjdKE+aheNHXpzyxHU9GLp+Szdybi6aGlb16DjeyMVgNn7bRAa
BKS/zwPosTE0UKnRPBFq1tHP62NkQyl++3oQIdN1lRlmkibOcjH0qobCrlFaiDDW10YHVZguOrxL
tTuaMlFB9vfGy4anM13EJCvQADyfo3Av/BJ7XIfnEIDs6z+W335bJrSfsxywA3I4F0pG4x1/OE3+
rJMuQhjqcmQyr0RDIQw045UiSkuO5wvuDLM3KnRNjXz+3wEQZZrTxUT4N1L8UdUYM77Pt4471Kc1
6aU3Qgj6Tg56VLEx6KxMU8RgS5+BSkaAlMYj/uxoQsUQW3ymvPHerZv4uHv22E5Za9rl535tS3E8
6QEc5oypGBL+FvoMMQnsVZbk51Zr3G1/RXjz/hOhSIjysx6jKSDF31T92Yn5ewhK/c47rjrzWubQ
Pv7sgF0yE8IPPdUzLxVnJqu9RfQUmLaMNRpLU7jgaSBgE6toJRrI2iJXLQcqFzP/zohzQ0sIITnH
Vb5+aY9XP6LsY1PDQ/TlEbuoFeDDYbQm/krF9vfGK9Sw3RsgVLD96OiRcAU3PuFAFVoz2xnef2G8
RzmKsfrHB3WVPBwkDxYxrKfhYtbH4plGh0NFwLrYetSqkEvOubwMswzkHoN1qgrN5aHsI/UzNd/k
N98roXWmppXtFSg3hr2YiuYdXUpshE/q/VdSVfXMHHkafd4OUWuQ1sRA9hW3DWg1PoUhkMF2LtUM
U4kI2t60ahyQNUNT3EQoY3LV3NGRk1DxhGidJHOT8qHL1H+Ajg4rKONn+o/IdrQF1z7CaCDfhv+7
4+I31s7kOz1zpTaqDHGbAW/2mIcXntA8JyvB1Lcjxln/HVCa6PBLsEOCleNcd45bGikkY9LlZqcD
eAZX3mMnT4kQYFANFBtVKDvX3jv3ly0MX48iDqOPlpRPjavY4VI+pVMFcu/MCfNkRwjH7jAeQw+P
1+9Xta7jlxmIXb6skjPKIT0yRJed7sA0xn/g7pwHo8ihRbe/S7YGBIal1F4FGqq4cwJg4WGAJPdT
A+PsCNpmPRmOfk8Vtgz4Twn18trcFqKhTWL1oKKZKl7Ub/MXrxlGNpRTG349OXDApLeu6b3KqV31
pbFRgYAo8YvzmSr4g+aW0HN3Tq/usGTVnnbUFEuMwEwnjsZngk9Pw2KV8SEqeBh0R4PZg+kWmBH+
HYf9ShYwxLXkRpJExfglk/CY26mzVgG6mJ/lNCR8mT9ERdfzOBmTcHjOKidFtSsot6Klk52ziWrL
KmTVNSNcYW1GOuJY35O4ZtJqppgj5hf/uNh4l+Zr44nj/z11DJ8G+x8E/GssFk4E8vdnkNK6rkrY
KxCz+kYE/Myokg7Nd8I2RsSJyduP7qAwxLQVZspsjJgEX9D6TnIyZ0R+HXEh2B8+SGDzoAxOE/Kr
49DPW6oBQ1+xLPpUkN+JRao5AMjhQNIx0NDs8x0J5/8EwK/rnepNb6l17cq7cRcEB0wJdMV9jtZV
eWkEzI0nKWqd0W2oNmW8cThJFrgSneBswSStNhOyoaLAGUHh0zBq+s7DOpViOUHPWPLXJEERSpJq
ir3BaUu4Fjhiq5atBGtwDWosC0iViAReSUBvrDW9QE+tnJa7LusvPM/GNHiCKig/qNmYF10l9asC
yV1UjT4R14+zZA1183NlmEM8xwqYW4IVkbewHSqk1TO9f0xMv3o//vR5b6wZZONdNJygvMS7Gwbs
7J2USuZLWJhlViBshw2ELI+ogUTYVV/psMKOk6n5A5SrP6RxZ9uXCd2iVSxkeXOKLNalWXJUN9ct
e0wjyMx6Odh7nQ86OPezW7G+tAbRQC4AiWUIdv1NH9coUKiOYURk3SFuk5+mF9NlYSj1ssVOt1ci
f4xINe2tyMWxn1VCS8a08m49nNwh/7B5+wDZ3kqwR4u+Ebyn+m5LjHFE68lVOeBZzIT9wWilNozy
XemVjDfqyOorMAZI7NidUyHB5N3ceBwz4WJKDM8Zm7ttGtHswS1K9mvufPa5J0TcI3+vuwkoIrfy
tg1v2LAo/hghBhHbeen+8Y3pOj8BOoiX+X+3auN1+OAmT02Kb3ezMghGz55p9Q0PUHfXoqWmQAgN
dxkASW2dZLxfwhogoMqxqu4rk14sjsCudDUfBdk4BKXsn+6QmApK06HP+xAvYq0lMN3jsangjDoX
lcTOHTpmUfxqH79+6HFMp3S7QO7p3Vz/VlzxwyKgqeWX9nXlTfY5HtAdmWNO36FitcnOt20xOx8v
Q1qnZPap0k+vzn7TMHuVf6Fwq4XKaLXKR7BZahuuSQdD02JyXb6UKYjAm+X7B9k68VNxrtd1rxVK
g1bIFPJR/qD49tdyWD5NRSLHsTkbnXl3RhrlspO3QeHIc1hBi41e/J2kGWYFd750+PcjKdOaCiRg
FvzsIZGVtsClcrY3coTGwDC/2poeQ1hf9twlDR2iyJ7M4Dkwo0NbGCL7iOLaumJD2uVSVk2nsWyK
VgFPtIlzMhg9jA/HO5jhpI7cxiNmhu0yRBJlqdyJuKidRJizOmZ3ULiacE8wvne3sz/cf2YG+q76
B3j76YNQp05japnQNu/4C+FHAtN/XJi/LzSQ3WgF7Rgz7VrpNdiKOYkaXs72kQriGNwQTvsaRR4g
HeRC/XY6o9HNaA2NpAWCjmnHSi9IA9DISrdasWAE2mUL3BDEvln1vr3RSvG+u/9EekXUKSqrJkMA
0+dG8DojQw2mUmaZoNEOdqd34qXNHrhWU1DXYKEGscrEwMkGQV4C1MCC884D4nYES0b61jZozxZV
bx9PKAP5XvfXaZqtxvfWv9nm4wiEpyLYdyHdAynXBNXDdakPvki3iU6t8yJjJ4fxANqJgqnxkyQ9
sKk4rMcLWUEe+W9ebWhlYLK3nWcNlH2VUbCE95aRKxYYr/iH1tKafirhmiI3Qw7D45T4a/Xsv2MN
zL0hAOlLe81pIAITSE3FD3qEFoMvDAkNyNPW88L6mlRIZ+B54qa8Z/nNNqF4RRFMD2PqAvSwvN5F
0/XOPbkgMSVDufFkjd6ZuOPMcwx9TTIOZ5gd4ljN3hLGl5iDTp4PI8YH6+Y+rFg6LE3hiunIYVSz
rJuy+WUPArZuH26XUctgV/Sb5HzqOH+ncP82YuaoeUy7AzLm9fAqbCMrqdgGEk/h7wbnP5vhnK2h
hXyiqdYoYaG/ITm+/LshlOwXeKbc/YcsMwaLPI0hEmY5gYCVYtBhQ9v4CA9rQ/7Rw5X/Y5wcuriI
pr5GuSGj4jvNhAf8Wh6rA0FQOk0zj4AE+w6nT2/+6r3IH/Kk80z+Z1W9FmeXhVLQ40a+CPbpKJpn
qBWMFCmeB2TvZHMBG58UHVe//X5Z2RjwqKuKzOLA54d8a5WfZfV8LrCo7y6gEHuHWpOPyskonszP
B49bIInmyDkTiaSlDkoKKxu0zngyENw8OJ/JZG3rHFOTxb0mvTZztKSdLniQG3A9ob0LMDMO0YPs
dPpUsNx6kgCokw9QKN/oAW/xD/EFlPMJ8O6pYT5/kK6EW/3aTBSTw5JCJzT1H+LbuaKnaQVP3lig
6+UmwoX9WytNfiWJlg/ch3x7wEk2NhmzZHTIwtTjRN2RMPHRykSu0Pr/OIjDsMGanijwiH0Mqe+a
gBbJxKAOGg72Q3/ZoilM+WmVtPbLibA+NmbYTwrxbc301whHIs9oorQJcE0AHOatF2GVi9CkoPBi
AoTEhpd5o0GU73tVyzxQyjX8GBvPv3Zesk+HCq7o7rpuekYoTK/NAo/0dkhEcHoWPxoeMfcRfaLI
wUYESuD5jBAeAxxhMht1ncE6hqwI4Yu7kFMKIyEnKoNv13u6CQPLs7Mew9GvrEQmRQQpDrnyaRNL
d74TCLi6bQAKqKCS5ZsjCFyj3q2cR/mDsfePpsJ3vPW2CsHBfJmEcZ/I9hdRt3MWj6Um0YXtZp0i
SBexrViWFX/1kWpIBBaS22iPfCH90vH1CiG7q/2Yi9KcWGfItG6795dqTsS9AND+c+bVz+eHan7m
b9Q0fcP7xSOryY7rzFk15IW6IOWcyuXVwm34Lq5C2ZQVgOKnDp/K/8Y61hf3Y9h8r6+ajHMQy/YM
i272utMI/BdpFJUd56V1A34ErMCjb6xWJ6x4NbZIQEkLTCxDHImEiAZrOVYvobIMjTrx7wASUau/
ekKhJ7d/ZbEcU2zN9H6fSrN0QXnXXic/KNbHS5+dh4iglfQazGLeHtypApfa+5WUghYtTHVmLJ4T
+Bn4fX2ktPqSyep1cO9W+GsIeKYrwQkF28uX89SnQu0tg9Lxum/FN7gBaGXmp+gOq/xALBbow92x
lBqATIw0GksRu75JU8EIazEbFEq9Xu8Ip6pGYBlAqzMrqz8qL6gd9pzGL34nc2NAGakLtrmPr5ke
Jc9nmq85BpJkFpak29j+LrapGZZf/UidJzHUJBxAVavNQL3GxiEL0C2OG8Ptopl78pjKy7D8LojH
d63JyER6YaTReJfAKcdhdFeOnlTaLGHQRMr6rer7rdoIJGEQ8lD+9QB5BQ4WtUxXUmExxw7nyQtK
WYCOh8q8QbN68BYHpqNxU7V4hWfwX9hOaDc7g/UW3mtZrNgxCFY8KYz2KfDk9eBLfIyziJ+Kc2zC
S9miwSl0rE39Y4ZTFo5qK3ibWC5Vn9U9udYPEQ9cT1w8v2es7JQRU6Kd24xHoIuW+xYymJyWV/Up
J3MmThY1ufi3cDUfytbAnxnk2tnMCJM9+iIvTFrvBarRw7hPJ1MkrB1MD0aL7gTiHd8tUixWH6oT
j4yE3MeLY6C6AmMPMrtQ5IlbIGXH7Dfnw8H7DQKLxUOusG7JDJ3qsZlbT/qlKkdbgAjq4c1qlB9O
4CSn1b0ASBVuuFcLE3PBx4VuDYg7lpnXGvUduecYgS8+5o9mx/HpQ9XEma/Q12rzm2wkmQRUOZtm
fvyM6q+tGJcZzkIT8nMo9nyk0+vHTRrrabd+GxLKYA/nLxgmuXsRRQPcMS2g0dRuKUcMuA9NF3T+
taVShu/0bVr+a/sI63b1JOKsr55uAX122+VoZKtx6xzBUsUyLSvLOiaphJVjWrC7W4Ya4SJYHVki
YgT9DwfBPQqOHYy2BhaGYIlIMJ0WoV0TUvSuwSmeYqd2pNSC1Mkkk0MIKAOsEfto8gFlBFik3pQD
qL8hH2tOgUNBH/YBhGc1FOUuHAbaAhNB0vC7zSE+icQDIUGbUVAvkW4y1p2nsUzxq9FvJYgumGi8
E9xCTVRmHntHrB9NCFclZqA5PILu9hT6/FUi/+/Dk4/T3hHHntrlwjhtzomVN2OK3cWQd0vR3HcG
F1CB34w2MC+dm0O7Doz916ln2cyipTE7R6byoHQpUJTPcgb80HyWsqxSB5VRu8DK1HkJnv9Vy07E
mZiVmbmuXudJbr3nql3Ct+5zL6xby8eZ0c+9B2xZseXgvZlbG6s7nccYKyEtXtU+/8XiRdhkbYbw
8nxwJXsjL6pVk8ZRFe+26zt0T25tW+CgiG67AVFFZaMhpkQaVVNGt9cY7QSHNZj0eVAfxe38KRxK
dOq7FT2N3OCwyZDYkqUUNVw+MykDrN3mtLSSUTYhTNgu4lydj1xn7Vls2v9Nuf9qkZLzf1JG3gNO
9qJu+BzyElRXbAMK+A8D7UJgwJgYxoWXxeo53NbhKG2QTpDuQuh2WZvS25/riW9O43a5SubBn7MC
rCAs83C8KV8bGNrXSKJhc4lbM+rCx9qFnJWMMiAIXWgsjJu5m3QyvEijCKicgmOUwkaIIL5pYW8q
q7Od5PwC6lhq4C2iJ0idmDKBCnS8sRKwFn8nR+cQgPYMnZh3DTuA8w/Nri5iJue6WVMobw2ao60k
yQPpugYBI05kLv+u60BwjKtwb1CDtwW3Ad1AXRQMbAEEHpGCHItfD307Su0HiAhjPTeIDhuZUpiU
6+wtEP8j3ur4E95+4eE7/ZWNu7EDrQhq/R/cM27V1sMCLqndQfK4dgeTh/GZCzSiivXH6uR5pK1o
uGyUD4UGKtQltUIeRXnjJhGlLhnqbR9Ux+qAR8b5kTZ+nbfn5fyesiSQc4zFhSRebpRTBfwSIXks
mB2MpUAoFVyy1J7o0KuTUHaNPFEvQsoNA+bdJoj4Mp5nxX8ZL55R8yo8JIFwZgF37qCi61MV1xJU
05BCTqYgvnvvhJ6WXTZhBd5eXGMdEipkuyd6hzHqL9DKk1uEGaKLlS6JgOEJr0P954mLdDcX/3QU
sXv7Qh7rXiPohwSJuV5d4cstNd1qAta4puONuhq1fUKgzyEksQp9KLLHmGfodP9Kj58QKavqGCFj
Ah3WUvqHmiN+28sOs8EeFyoSE9ZykU0peR+LdW9c+1siEI9lByOHr6LtzUeZybwSfHB6VVULpUjT
vOuKP1ekgmwCf3JoW2d98mpYekAPxvbILeBUOpyNVX5NC4D2Xymz3w5jsaTUJyooXbBxL6ELvhQ3
x7Yxj8td1jXYIQF7/LS1DrnB69oyYNh8Jd58WsYYywVekYM+iCpTVhszbYSVJPi1ElCs+v5S9VTi
F4gnhvalQ7l/G3tsSdR7so1Hx01JcnTAkeG1rcRHewEXp0GgRvCBV9L0K4br8wJj73SJO6JSG6pP
lQwTRNHXW8+Rc7vXr7KAv1NhxF1jUxojgsrI4Dl13akDCrkIh37GV3G5VPhwQC25TyDTDgTdk59d
OeB7i/yC7g0akVSrjl3552QhIRsmYWSO5TUkuUHTiyHWH5Ld4Y9J3M7UYSXjW0LaU2PqldR8LK7e
Izio4rUw/BZUWzLWB95o5/q9F1LHl1IfqSuEzYkbBmD503N9/PkTS+fmCpkIs0ou/F5tTb/7Cfbu
7t7yGsUzn+ozfVzOpTtpTPIr9yWCSN3qRUfV842sPgSry9P2l/VL7wKC4oPcD65xz6zz9Qv04E6r
+GCMJ8ONxgjenjB6pHKWh1iq8ROATExsyXbNEk6l4cs15I3t7z36+4CTotnJn/kaIzGzOksLExhq
JKoLbAZEV0xd7uQ6nKfdqixUhoJl779wjbtY3+4WRcF1LcCePL3qpinKEUoyMjZA4ba0BjtDI4QS
+kidKd5GgRBbhKU5IGTt7CFYTSKItrPndmhev2nulO2oRzfJJra1UVnCoimOmR+eXpsSx3KU/yvI
M7FDElw8+elTsZo0mCG1b+5OO0dOaQEZ9JpP+qheZe+Z1hKms2C9UbHyTZqdGKJ57ScPa875odD6
JM1x0/xUuQA8l1bO6DegMly48W5xFCOOzXHXDMztIdrkUxPjGWue0qw+/wrrpRwtbaT9Qbb+HtsS
W81YgxpQSzAldgUOAq2g0NOU4FzkVzXTqXejK0s+F+QIlusaobqd0FGUG7K93ljI98JX079yL8b3
G+/xQmtp7ekW+92+O7ZCCw8y5ew2wezZURh78RcV1iKmmsMB1hhfyR0S6o++MoP9Hg+qZINQiGXJ
mcWA16uuIL7q9RVNjwG0IbFO6JNasphl8k4lQk/gQg19bXI6uUUDHomr60Jl8wMRGBc1g//2l8QH
13rl7A2GZdhK80IZ5kXcHjFp4YhmKAMmEwOtNGworQ/RONN5mcpU4fHX68/1iX8TCyiRRdKiWaHW
HPOjuvFcLpakf8WUbolgjRZC4xxUoyO6k10xFqgOQJf8aAY2AYHbMtiow/l7LHRNLPRnKewHx8DI
z/JrhbIg+ujTiNcnPsy4wJA+Qq/k3Ay8eoJ5VZ63z7pF8dDPnn/FPFsOfdoA4ZF2fUFvrwIzxfTa
QobHcZFQLl/mQ9ULzCTYbNK0QhHNAN6M5hY0cJqoIkFj662z7ev1Kq05Xp31zwgoX/MalzulVlhn
xyT+20qoArT0d3qDlu/qyGZMunx2KrkBULbbMToPFWraRDOcXhxNxEZ0KMkVD4ukYBSVmCuFNU8/
4jD1Mfs0UNBX6fR0/8xEjNMN8IgvjLCZE8ZJkrKf0nWE+iQALwnQnMznyTOpIiecL59+dXWow9Dq
NwNTvR1bDFVUrGnIhUkjXWK3EPwVY0gIyBahfhngKItBxI0LF+De1m4dXM8fPRAV9e0/EvnBdUnh
5GvwwuaszQ/qByBCmNL4BIbmqJNWSDT1hXJrqIPHdesFInuDgjQ00/kxV/MTvehLXtVsXnDd29Zt
cSbRj6g5KR6I3+jE2L47kJAAplmSRXdKflZN0oMXs51QpD+0iEaEHeYs8yjxOFPZmk0ZHr/uKhJa
HAR3tuiaM6uWkdL5vm1oEwVJ9XrvRUUxQzl4OLfaF5i1onLaVobDMvbd4+B9Y6lq1Xh5UZv94xj4
S2OEU2L4A0oEHcm2m/zAlNrbFCarQWMQQaJtXz8VjcvosyKsFqeibl1yUvCIhfIrSJADPksl2i74
o53RlNavR8J+d9BIyfV2UpQ0IEY258Za7YIEE1mfKYJYltXJVi54OcNvpe0Jr4S+Ya8X46HuIxvt
rCROvO15jpz5SUs2DgY8hhTxTrd9bt81iTq6FR3lO5eOwjgHrwqPLONwT54LS3euq6jgbXmwy2NV
cPAjM6osyaa1uArIVQ68AfGaXbFVoWo0mVS92anhDjfbafkv4zqhztsTkC57jFgTzW/4pTWI7g8k
aMAvev36Jl4MO8mp1W7HM02a1tu2IfP/IQFf/Z6QhC24PxixENuchiegJTC45oVpbpP5slKmbECi
hhDDEPhwCTrWDd+VB2FwL6MAFphme9SDnZW8B3XnLXERlySC2Pjm1E0Tcu9pOVnaFRtPj1Bgirld
2sL7PvZ+0HoRo6VJHbzlJpXDMfemKkcY38IDd0F6cGgGCPlmdOdGz1vEBkWleEatmvf4gZxrv81F
A89rUFMTNNlQ5YXW+rS2S5g23vs+xD72Rkuv6hVtc1rHV30B2SimJi6zizaf0C78PfD0YaA5mW8H
UEvOwtZmoku5kB/77PIIbfLpyOJoGg5+30pf9ijxiyvLlLrbagl4KE8v8wBchfnKRRpBS6Opx1++
pu2CQahZ/LNR369Cc+plLAEe/Ep7Wq9JORniLCIXVnPq1nbzSrgjrBsFSNJGqMmvXR2EpYcyPTHZ
lyRy7Tt739aVNLaTLsDScM2ZqiIVPizaoYGyQHqnve5YVDK26/C2/Kn39Be1shZ0a3EgAF/Bt+QP
O9wMeHGClQCxxSg9gGzEoyh33cRmr45wy17+PfpvY7qBSxuim4cE3bsF3poZC2wDzdNyQ1H9Fi87
e0wt1k1ihGdjvVwxnUtn5Of9xhfQyampeqxi62sN2KW+g3mqX1a66D2tN9N6YaHjSE6BFV+iRx5u
Zhfjl8wqkoITPgjxRNsdmRW6vutBObWPTBELpecTeCxmabFNhG/3qm6Kzh9PRZPEwC3jtB2P6HnM
RHmPVSghh6RWmAds83dEpZmkXRTPsstH/QirtLrDAnUjUCpqj1nI0FZjtyKsUFjWgV/XZXEcfvjX
62CEqH/+BHbEUvOD4U3549xitZL7ReF0kzeNvxVya32kkwFDrF562nwjukNWqyIFHPbzKT80YNrx
RLIqDL+cUhnMyGmNEWrNc5o0zxvrAcxaXOwVvFUSBF2XOPmub58yaebFpcmUxMCtlvJveMu1uY1r
aN0NAEZfScacYLcgZAOIAzQjn/00RCbXXtcmmM9WtUrndbV+EPI0wjefU2pbx1niB/cZ8nQx++T5
JS05qtCQ+T7w2StwIQfaWQ6n3DuS4UXkfjbN1AOY//+xDrMPBWXWIgRCmpG6O+l7qM72uweSGxfQ
yQwQfOE8kFqxM6Tc0lle6/y4GcGATwqsDwV3CnQFxzXH5SvltLzBAW9YiISe2Xe7fx4QkQ0lYBoa
ELVZimTGEitG9O6fJDfYOmha5VcQ8z4bL+CKJSV1wMIiIRwIHnzDZ868EFsN0V1nGgjZ1gcidxAI
6ercCiiXhqZwE2/yq6GHLGy3Xg+NT+qemRvqjYUHHeawXMpkJchrud/slHIV6qFPEPHCkPVOdYTR
4DGXXuzCihRuk5WBhJMHe3JBMtNm2LA9GD2xh/baANpEXfEtIwOaVMZ/IAj8KundJsML3UTe+IYE
/Ql2CBAroD6KawLuux6w+DcDAn7QoVpvMnm6OJ9Thwow/Ed7rAqX2R+/reVe897pdscVNickBE74
kokuKmcwfp65EqGbDs+1v0RcJX5XHFV9J1FqQSDL7JlEs9KABlE3sOt/gr0qRQrbC7kzTvTnJErp
Aa+bx5ARbTOv/92c3jj+bUXrEt3LYngNXHXx2kExTjibHwIEdW2Rvadbo5n0LcnYvqgK1OXK7oB0
k0Qj8sJNOlj+HhPMSpDKR93b1PezlJ3595Zywz9FLdhIaw7fivmNPEHWSGHj/vkbZUCDpaVuoULh
LU9uAXMoSK9yoLzKjtHiAt6iPmbTn/tFmIYLSnm0QLbv8z/ZTH3VFT8STmkom0ik7STT1gkvtg66
2hTomHmyC6Vg9JSQzJIOvClHZT4LF988QtvoJeBbYcYQ4IjpDdpZdX3pxIPO/JgW1aAX5IdZUoUu
YLwiKFvpy+hM5VvziFEMsk/fbm08VM1ZG1cf63a23lsji/fhC7RQ8lUaC+OWYbutoJMiKkLPq9e8
XchHJlAIWDnbdsEJe01uT7o+Gq4o1XqLFqIwcALhhYFVCofhPFuzxHpuePWJ0dr/S5ITK7BbcfED
GieHyWqObIMZwqUa2oYpAKkbltCg7+NxFENm+XhPRiay1eIzE8bJzfRyzve36tymdL1J5Sai0rtH
ygQu9me3tDD52HdcX9gcWSPlnctul74GV4X4vQvjuVx4X4K5puv0RaTeD8eo/+fmRHS9stfDNydv
hwQxFnQZWIhgIiJnZtw9p8y8jYSVFQH94t/6kZdbY06pbjLy6EuU6ruMW+J8PLT5RCP7mqJ5vNlv
8FOIDHq1epST25uhY/m8aOsHIz30Acupw/sjZ3/3buugoLomnRFZoEEC/SlTDgsuTsGwg69BvsZp
W03wlUgS7yuRtPf4qcgMFsGVIapvahWp8+Li0yECDtFr70C44fUAHzprL33QXaUe0aJPl3Z4WRWN
sMhXKdFV77PncqCeiM+6us2AsnsWQKqSJzqWCrsLaEE+sNJuat++DZO+j1jesafZfecGbybn5dq1
IFm6Y7tRDj/am4Cznt7uuiOy01At4mAHKm4Hg4lfKuXCABtQPyuF9Y0w/bXM+uN6tZIwZaX5i6+I
1+4KjsdLdzT4S7uypdcMVaraDIrtsKE1FNkmzaru+qbHRXWXJ891RNqfScYSY941TlG0ZUUNe6AJ
2efN4iz8V3WLpERPLG66jKzwb77MwM5B28xRthZNQo5Iay8CJFyrIivz+ESu6D58kKWnK3Uv4UGT
hmJP+YoLiJwwNobKZ44CWLe51SRiktZpBmmhLX9thSLxFEMdzB8QdT8OANtzSbJD7gCGpNoKnmiW
OlXtO1FDfldbPvdSd36wnyfduy0CJetmXANQXpygMds34ezcLRSzEEfVOeLNOFDZRzl6AHzVwuoP
LPLxNrsotPMcZnPtbBVkCjWb1sdxK0VfiYFkt/Vm95TVG0U/OCPx6pdUOy616Sp5T9HMJcml6RqL
wNMovobVXsKmXjtbssldSZjjnbEmipxLW8bwcEQhrnU6l8dhY55abSPzvEbIpHnv332xzsKMxrRn
97RjkdYHwlkYhT00QkBj4UIAhOR/w33BY7ZmCnoGd7hMbxjiXPL4nR9nLnMdfwDRtDc4ZJkDGARL
wNoAPGItpSxR1BCWQ6YxkonjWXE8y6rUAzZY1UaK6sC4TmWKGkoIdOoxM9+InxEsepW+mhVxmqFJ
7nbElB/LSFsL9LjhOMs8yPgtPpY0OYtz6WAUWgUDzcGIPTGTRrD/mSphIQX7jyi4jCSHQEmnJvyR
k5vUU37cXv3t0BkpP+BG0BSzzvb3F2S8qx27H3tRmz1efmNL7e6gSxzGUW0b0tRaPzCaBbBGYEMJ
+8Z+6I7uk0JwydMsY88s5Tj6YdtaeW5IyDIcx05PhZOXbO8I2hvdDmG4MswugAEXeYJrv85GlEo1
O6Q50bIIxVS1U/O+42CZLMAOUJ1Wrp2MYpUL7cjaUqZlVP4z6bYAChTis6BOYqwTmnwHfQRrKgKE
aW5XgyrxAaYimkGOPgz8yl+a8OBFVtiiih/AXQCog9sqsEh0das639yd/Nodvkfic92l1+0xsgF8
ctGe+wBI67XEZgmPm45BXrVlyy49qlozTBvCofixOd8OznO3tifzd1Rj0seUIrd9vFOC9XJ0CrRA
ScEz6x+o37gc8uNw2yH0uyfpIKMZ9eKpG8vlt/bP19LGp+U2bZ1y/Lel/zKRTvjFAw4sWpt73l5a
d90HikZPcVT1gzxImc6suONN7cRa9GMbY5Kb6h7i7r9cjQ16dRfTnmB5toKlvoTey3tpNsuq4pEy
aSECezsACVMOlOwxKgHADRGsKtkPrcqJL3bw/L6GI25QWrbV/8oRkKsnTvo7HGxa6sitUOOKMQup
pvD85JgtEQWeuQydpkugJBJus2e/0N9NfMAUJ7OrI/5PkJbN9aDgnblwqhRa0OQYnTdWnkL9mTM+
m4ifcvyBW9JqJcKDbH8lUNSYctSIbo/GKmQpOJvWX5PA/MUnQ/I9i+moMoti4HLv7HYeFjsD0iIC
NMW8ros9L59h7AQUYd2sPT/1q0BH78es+Pm204mdBmyM/BaraVCtyN78TIuxj4PF6LCs0rNBSBef
lm5gIuQ7iGWq7vmcyeMYOOeWWtpzHrOtsKTSQjhOeixawnz40R0d0tlUp5zpmrkncx4iACQfCPsC
IDy8/atRDHOEQq2x4EMXEcX1rHvR5zbXNE0n92rwlnrTDvCgnS5Gi/rKDfKNwGjbhITUaCuanhNd
u4PrU/vSzRh6DAr8nYgl9lIlknRaOpH32BVJyvFl6A0aYod8eYIB3ytcWVArxGULtJbJEo5OHVO1
GUCbMrIHBiMdLY0vxcyFIu8Kqaqisc2VjrsasEDFHrikmEXIR/7hska8NnubTIKJyWxG0MFf2XqU
FohhbLYr3OJyBC70igPS3JQPVMSD5veHfRdXnNU3lF9VBLVVq8Tio9eoFFLyqmPYDoVb0Cmq7TBP
usLvSBkIHRoPV9Ub19I8dOPJTrEzRxevYdwvt1jKsIxgTT4EpNUoLYfcAl79kUgbh7W3aQdhjDcZ
99Wk/RNIU4QaE8boVt9OaOd8qbQsACnfJzugFGVu38wcitjg8MO6TaeXQ3UmmznA3b1HnhsqkiPJ
w1StM9TZD1heTUsG26XR85ZnYEAH50iYxuYMFBdX5Zo5LiRfjaxB1RjQfO+OvbYc5k0fB0Iya9DZ
qLTDAECWrNGS7t/KhF0UFfturccFjgYSBLQyKuzsxmWOBCdCNB0Ac/hxd6NQTMUPpjeawGgVB2nb
KqbFjx8vhGtkBgfOPRZXMNUWE0miMZ3X6hNxhtMzvVpyi6VoSdicoLBwo1HheXP3UfBsie23biEs
GAI0WSOfOO9BhTgfBmPOrA+6XFcWZx/RomSTA8f97xQPHjyBqMVEJpJdVTyMJpSHVH2l81zAWkqU
bdv/Tlj4qdAotUUqNw7+axYTidWUJRQAmlFyEQY3Rru/0PgFPAEf0HV3HyuCW1aJ4I7N3spkRjM/
/STA/0A7Ms25vHRl0VuKPCmrT1dB0cNbirgeAdfn3rln7ktvzfU1+kkrjextB7dJ7bYWKep7dB0U
c84IuK15v/9YjnrmIvLyZ4pU6cuDcHjW7MB/7qWJIMZe7pv3daaG8fFFucHQ/T+CwvtMgstpM4AA
35Mbskme5DBHAJo+/98lcL9PlYXBHEbHz4o837BOrCtvAtJv48kbVw/2IVCqO9LAIP24Lw24itG1
SAtuf3UuToKh5kOTBdCIeml+P+kfwwG0m4SB+mZLfRmYfQbEavlAlNQZbxO7rZCnpDU1rzK+2MOr
Anxh4CU2VO7sWBvuwpo0p6KnvAU1ovlyl8i5JaSk9vXqKkT7j9eIXvbqw7MwHOWkrWUcL99aJe2c
9QV5vlSoR+ZsiXupWZXJ5AYfjUhx8ZbEXDUVWSUNtFHb07aFsYjY6sM1L7OD4/vDRJBFd0AOJSVS
PD6KZ0wxPyA8jdOPYJqkpkIDnj6dYop2ItIFWYfPjQfov+HGLHm9pL269Frlp3DiGGee1QIAq6W+
WVACneUMwq5XeyhDBunDqK0ZcGtEQdfMWPIKBmHDMwHYiqYclaOMrVyFIBSEBGBiNkqdKxtaTfBO
Mh82xWSt6vZ5lkErDrqP0EDvt1u2IbmJcToMzJEqvtS3TrQ7rVb7rAZ6vHv/vEVlmwOxFraLu0GB
JG3SykaAaDx/03s8FbQC+1MLzuJMv0hAOUPBX6YqeCheSNpJukU6rjvd8RcmXzPVjVY/AR66Z2Sv
PJ3ExqoXCrmsBFKaz5maR7dLomq244WpehDLhu2QnPvl/w7RP5DGLDywnh50dDxMBSn/XIomxCcJ
2QkILSKbitVVwo4u4V+LZmQ3szikv/cxqdx1T5OrVpAzsbj9jOydOsg4Z4sw5f64xvOaj8kDIHBh
vZnm2ShKkRGb63tE+tP2ek6WTGUsy76syIjSzf+knD9LLEpD2k9HkodaI6iIVvmD2krIyQrYkbru
LKIa8I7unOY9cstg4VnweRkqmxvkQdjiM5lIrkOiqjWgllm4zAWvabzKYd3uriibDq4Psnr81YO/
TyLyQ0LIs5+QpU1+RwgywF9lBO4PZ9a6EXEJXaGjSh3D0L7m7KWv+uytSU6eG6Eiwt6leRjzNRQe
8UG5zkFITtdz9BvgLaDldPcVPmaTF4U4MN8yzVJktomLaDDbUCmyncxozTYqWhFC7YXixeDGFFm8
4t/0iIiWJQnOMFQnYLDKa9bLOXGKNQGNUUULoCBSg595+FEeD+Z1zSHfHsBo0C/TKs+4Bm/fhJ+Z
v5IHgsreGgTV5g9fn6ehVUu73E1lT4vTcbUge/1PC9KpPWK/mrEzes4NghUgZ7fgEUM5ac+1ch+4
rJGyNkRGG7kopB64F9KgKqWGst/knI2A2elR0KMRJxGLpG5QQAm+oMMz+SHF37/qYuLwWmFsSCSq
j/7ra/3NwiSVNcVjudRRtJ802UZ+fO6wMnJ8QDelJ4iqVzQAJDcBlmcwVsT7iBsdzJMOqMGR00Fu
Pd1SovIyx2AJTWcEtPF/arATHLuOnEDUMYfgGCNzCIXnCydDz0u7AS4+ZP/kM29+zzkfPTgtwwgC
SsQK8FtGkqexPDH+hB6wxtCmDrg/YoEUY413o/Xl7jOJq3dyQlDAVLlmNQaXbW8dOa9aWmxjjeCi
jZQct0jLzeo1lcK/tEUyR6k/EjKx66+JDlGCFlXx4wn/X3ZN7bBz/+RAfM0VKXN9mWSHob4OSx9f
UYNjpA3oKIQQthvuHDygJz2d+lS23Y8Z8r2d3l6QATPPVPIg0pLOtnpT1aCS1HJrqutyGniVg0bk
OMT7sNAQ7IpWyqguiI48WJIljUvOV+37dl0pftMi2qlXhuHtV5NSeLJa+pcBuc89Poivl4hH+pwb
Jt2gR0cw8c5kq81LLWZ4lV6AjBGunuEtuQazVqlAsXtYKu3uVX6y50xiNXXRRuYQ9SNDJknhX26C
sWyX9t/cWlyVB9kz0hbUXx4sFDmDBXZ0OsiSs7c3ByWHQRyDRsapZG5aC5nAn8q+5xDFBFFLkQ7r
0/7+HFKR6dqzmkBu3e/aU7xrF4pNl97Rs8wafs8cFYjGM9L/dw+vs4D8Snjuzoc0JR+Ak7TNkkkV
4RSyh34qK9qhhHRehOE7qvrkkMPPLEmRtJT673YqxX6EGn2I3Q9Rktj7TQUGkHzVseoYg6KIXWTe
jAA+c+n7oC2dG2J2BTMKhEXZg/BlxOwRctdn7AWA4ixoN2cCKD0P8OA2fnGyoDArZYxl/rhuGP1e
higMpx0LgsQKT6SiqQ+8uOEIZvkX7zVvMqW5QTbfUhGYyklMUw/ybESMoSU/0tsMrQEs2uBQgTI7
SOgrNoLthidqeAlmD64P7EwAzybUsmy3/epNnG/1eStXgvJFBTafrKQf0z4+zESgQ7cbNlMGu92v
Lq5KWhz8OfaVwadl+irbfJjG1mhWCo78Zi98yg3ARoOjNuCXRvJl//vdl34MUg8iZZ0ewEfeWGLN
TvW2wccz7AAz0WsfiRUJXf+RAh57U+KzpY3HOH6pMm/MkLpLIlujuQpOu68UlUuxp1ukcWp3mFUc
AVLIBIP/I1J7q+Sh3YMYD7LXjjncCsikuWnGFxagyqaV24F15d9omUd8BlN5hGJiKqPcWREGfFmr
GrX1zbp9sHITOEgtK8WZLI/WIVjhV6RIhqdYTsxDl47Xp4W/v9WUdZLvGQZT4AlT2sg3yfXY/JMW
TohmAwFtoY6vvSWpqGmwaE3wy5xE+Ngs8Xi8Q8eR3MeKLYcGy39PtwlO7Wr6bSWezcsu/PC9b4N+
xHHhOcxBWOcf/luW9yojCRTHtJGHnIYDhzmh3DPEZ88zOsNr803nPs+7C0JzWca02DLhw8IhcggN
NBeG3LmGhHi2J4lCmI7RfcCHlMwk1iDHTV7BPG2o76xcae2OUdcK5uRD+6dyJ32FpVfQiGhsXb7t
3f9cJPO1VhTB7zPX/BUQGPTTqKLiifkUqiWDbBT8dG4cvQJzPofZTXiEGwREhV9O29zVTQULFr+f
9+w8iks61h6CG0HG1o/0BQa/zLQrsU1FE6vwOzfnaV8kCTBl7dU8cnXT829J1qXDs9chEbh34Y+g
4IAORkSEFJp9axuAQeISypisdG9Wb5zJAiu4YAjoifmG3MYt660LKzMrmCRI44HbMUQ1WU709FiV
1lFoMw5+JcPmtmev8XUs4+B3slIBX2O7pJ9OXKYbtQWTgVNFmAeHfUpShLTaVO7qD1f1VVccRVEs
r90+ocpHCjsbwXOgkkfnV6HacLtnP/qDgwKzJvXfXrseY5fBKXHjaPHjziAD+rsOtj3Vf5FinTgE
xaZhE4ty7JKxxK66BDlBUy6zMaas3fCcQTCnUoDqqp3w6XXjwwCv1+8KcveN3joXbMhGwPKk8A1C
o6kWeQS5QpoJHVh9PWo8vDBSqVPguDJdxDZHoip44adRwcHP82ppeBBg4+DmhF1vhomJcqNH9bOb
Qo2KcT0nZaH9S4S3BTyopBgllKad43t/sJEMtTscFgWD5TxCjqFg/3fw7O1sPkpLJ7WbovY4VxYg
29LViPc4Sgcmg3ShceIIL8LNxtMynW0Oceht+xJPzN2163g17Bvhu6fVuzgAw6Oox+h5z7OZO1DS
9izYwMqv0hwIGd1x+RV3aqtj6qKHLDmCMgjtw0FsLCgWAiGpJbEN3qi0zrKksNQPKD1x6XorFoZS
BcYuq7xh2Vb6AIayn8Wo/AWS4P9QwTCmiKha8uW/J0RdHbRksnPbc069xapgPBTxJ1Ye3xHoZjsq
V00+KQp4SlSBXEW4EJL2TfvooNT7c4kJqzNkd8tGhWaWuQU3L8/hYiUOb6JpNlfm3lu5oO13EfOc
XmO7tt0FxhC2PpRdnwMtDLuNvBQnEvuCxeh0tGQwLazaLo04twQFvsuPQaBNzyJWrGpBazGnVyz8
vuhEZp0Vrc6fsj+HY5mlUPXYIwfNfWZzEh9wNEa34WOExqBrpA7PwOfEaSqu7rRfJTfsgvODSY4I
32FxaBinnMx0vQZQk1SDfOJ5W8bDHfmVORZ04ymafttTiP9zlI5JvLxjA0yFYZ4m3DdzYiQbrIc7
aZmJKnqO7f6+uazQyJ9Xh44/AUfbm2QKeqlwfbmczp2T9Ig8DtFncsQBDqR2unSR+wkiskRPnJlF
FNNgjIu65zlV4s7M/i9/+WaZVbyN/X4eoJXcLTRaKiinHHmJUzPOmola8OXF6ktzsZuYme1/mwd6
AZNNEXR8Te28PPrmmUC+EeE9egf0jgOH0IgMPywDQCVq2cS+YOY9iPWn19BJZpcM6W+kDQOYYXmi
S2YDiQttypJjJzZ3pU93kBZpr1ldHO1GYXw2etx3OYGHk9Q6ncgV3HVufhV32rJ37atBtI8uhV9K
ReGWwG7WzVsh+x9V81Ao4pDZuxJsBekufRifeQFvI42I31bHK99aJqZZtTKdhUdtA4lVB7IfsklS
QtAAsjEgODnVQXTLfe1zfARQUOZTcWQpNyBmmVjykR7mwKLWy+c0UFjAr0o8El01kS67MC/2RWhK
Xyx7Eb+QVKyd1YNXSWGFk5V1Ag2LCNebQJ+N0zMteiq8l10aIj7ZSbaR4ANsdcA2d/+8oRMnuS9l
RYkZ1JLgHp7Bbf9Y0moI7Fx8CxGjm8CTsVVnI7wfbqxLoPBWpOqslW411EUzO6ouhQ8Njbgim7bw
12Mexo3mZ72lMF1HCvjT5k1kOVjhkP7nvHJnyMBySIiiekvhqVupWCGIOI2BFia0HQCu4Xoh3+dH
X8IXeXVHgLDGLSv/jaT6jauAG23dQH/4qBiZ8u5MfSi3aL4eCSA/pS5AH4JIg/lCy+zJLWDrXHFd
mRuqnluqvOeAWoTxfqxK9qwWkB7s/I69hkSx68hLWyjJOY/TU7jjeZemkVKypAFtSM62jO2UxyS0
TS6PGEHPPQOIKqZJf/iGtIBzinnALENUDzomX5g8fQpvW7rfRPsECYZhfx/ZyRdXbhGsjnSPp3qk
Ld0WPMd/bPWU6kqGWDo9THoXZgpFEim6FOofZW95y5qW9QEldpPA0vowSY7nE3eOiL/Ml+rVoybD
IUHQc88n1pi46CGgZ+5j6FNpEzjKieTZ+57m5PXu+zDWs/cZ/6F0qudLEucCjYN3+zNxjVDcJaA1
IGb2i9gJcgJ5HsiAnIdvnuKWQ2Zy55ynEGlBtgJRXy66W4FIBkZREWJwTiox31HClOUwRECHV9As
h7OFTlJ5SJGxZCqbTA2kbgsqB9/7ajQWx8oUl+x8gm9IhZq2WGAqpFIl4qodBoVM05qJEaBkjwTU
ewX5+uZh9sRZtvUND0mcZre0W5ILNfLFQLVEHfhnrzGJoIH3/yJoylmgj4ahhafm+1hKoF0FTwwI
GSVTc8jL1caJOmK2LnMdfbuq6m750sW6cUn61cmLkuJSmdv7d/ZKMtA8f3i5tWdLZ5X4fPp3wPDX
5IB8s52c9T7FLR8IEWDHuQeyvycmQL/pQFnt8S5YecXGs5tVNUfuI1x56tPY8bgV88jgBZAn+Jxr
T5i8eDWxoMTn6bPihGulZJfGly0C2MVF4gQ3tfoz3Peh3IhxhVsRt8+CHIyDIm1ROTUDfIWHm8Mo
YJnUWxp9ZSsbinwPUBK9tZiOHQ+S1Pwyzt/F7wzhQNrL4sJC+UOKLm3RQkmhpheIEsXEN6IBCpv6
J2FEaCQqEcVxgSUFjdkxaPi6iwr6Ykr8pKyQLRRfSjVfB2zorJqH1BvXKXOOYfmPu21dq2qAogbq
TStvbnraiUpG42PFZlkxclXL7Fe7EtYj9VtL3rm9Kukk5iSswvtBClxq341PnV3hEtLf946lL1KS
UzuX0aJLCZAJoMC7hRnDAXld/4SPDJuSHEpKNZdydZGd16ATlv4AW/gPAgHqSDLzXnTzSp1dYuCK
cSGWmhQlfZpF2kEZAe8ZxH/a0450apwPxOMScdFKFqVmf+50hSlT3BKJptQ4GYfuCKGb/ptd9gPp
+9VuXtWZAQIc0o0tKSKbY9b2kr0JMXy0/KK8d5N8r3NmfVdFku4+eeEt3haggyqliibqAyhKivrD
7TP45qfJb9aWe21SuLlcodCEgOq9ScrguuBxqNLRHVV8CVqfyRJBx6MeiSVITsXkcivmFvW+++Vm
IWYTxkuxs48tC5EXyY4z82Ss16XnPon4uvGoKhv9TlQNttBm3bv29bptKl/Ros712BYYDQIoUnNc
mVoSy/IwvOelydvN9NPOso64gtfZXhTfl02QpWY14+eLRBLNbOJY+n7CQ7VImF/vomR9tIO3NCat
SKfPZKdZKfAzGAeeDhKtLUPlXONZEYpaLXEPo1kNrfDWYad8KkUMMvGc+wwEDqy0x1sw1szDkBXp
c6P+Z5BMA+uO6LN8DLhXGyRKcbjTOR6ny1VXmw0HJVvieNoUxh8goo323xRHKOgcCfolHFw/2hUF
j8+vcqtV6OCLtf0mh3tVuKJ/j5oxHU1NRvPVnbSHDcgPVKq3hakVELlAQUD9LvORU5xS/rsrTm4Q
r6e7+6bR42t0xEvoJaxVIuSYalYGSS+bxawsEx/H1Y0h5TO0ayACldhtxhRBnwxfxhj4PvOMER95
1/wy0VHuUYu1d+f3O1wOAmETzowK0XXmFeygTCiPD/iqD1bOVhQnKFfHKhfsB8UpLXAo/X+pcXxx
bgheS2j+bHN09XsQgMuwPRCQ+LbXhZ15/IOLpnG6eXRTs6dtdUnGoWY4L6fBwn1I6SbLaMbypnzI
odkoYiEjJa+w7FgRTLA6Dioewmu83UgT1+Cdp9g7Y2gK8iQMR+j3CVKVeAz4QBBpdM1UDdBVbEhr
0h/TH2Dbktg/pkA5Xu7M1byaJbx/Sn+C4SRokxnN6m23UjHTUerL5VpM1Bsn5uVfXUNxfP3eEdKQ
mAbcoTCIlppDsjua0NYGRGzxU9dj/b0ESzbL8hR1fFWx+sRM9qbruMGRxTOzrrGbWuyS/xuCgWdj
Nk6JcgMQ/EMD/aqPl9tYMSUh7SH/VaEJZyW2YKzS6RiSscABXV4lwhN2o8C6NZljvbftrcpysh3J
pf1i7vBc2jQbw0ryl6GEnZa1ewfWNmACovk8KNwCm75LLciBCMRC4S6zNCgAAK9bUuPMCeIXoDVz
08hhC5QpwQa+zOa6T2dvzyjfl14kTWod3cORPEj+2QYL06ccBz39tQPBBbBGOf6evvg7ihFxF1O4
PNQFEYeNzslw6giiAFHumCDvpIyLjKRL5uG+Iu6RCS/3gRQnHgwP/5ly6Iq+Igwk6CUB2sm6ROPG
CwB8D3R3+jK4bGwwejZWrp+QamSEqEmORuhaUXyBFY8n0619IfIR8T+mjRTbr2KGkvhJsKVcXf7I
GiyD51iDW0ij8Qy/cmpWGqbWuaY9OJ8pDr5cguN4B7CJS7SAgQ47zmCq9dAmjpbOUTLG6OXZPfcT
TUOBWO2bBAboGp6U3H9W5BrzOckDMR39I3V6SPib6DaaFh5ux6sSkiZPcRARUMGe6FHToc/gwpiQ
QIXN+lyC47QHQQyQ0fLizvdB2m0b4FV7WJAxC6RvRdEE0fISOAtNrlXelnySdXUp3CH9vlRBQNPY
5Lv6TA62pxmLFYFTUltNcumDWJsEqB3ntGo3F95FA4gsRyS5vrea7y0a5xsIxV/HIiIlhY7N39OR
/P8PYkgFf0euhoEJAFDitm6wPLlGx0HXSrZIVWl/lfohEqTLb02zJw5dzM3731TLqFhS2VUT2HUt
vIUtzXiyl118fU7yss/Ui3SMcEmTR4rNPUwWg7CnYIrBOBtvFuRpj8glHgU+0kO4dkgKZ7Iqk/FZ
3NWdoCjoSU/dYuice2rRnaivlBlS6oU2IIvYfkuc/eJbJWJn4+wz7YAD3UT/hwFG1AyH66JLkamv
9gdVro0B6vUZZb2InsSHP94RLy4HFE3F3WqchonmupuCjrsl6q5mNXeC6gn6CtuQ+4QDIVJ1a+um
+x+KZlsdRkgs3l7OY24btihPGTaW2U/giou4jqWN2Bv8CNlM5DxrgqoZ+eTHQqmzspgs6G79z7xQ
NeOqbQ0ieV6n9WvHrZXZqvslj9y30WaOHYJaAe7yuE0PQ2UE9M43YNMim9JXKAI+7PS0/rpM+gj3
1fxu0hu2KIgdHqJtlLS7lJ94vr4opDJWb9Mmd9ud3F/t+yUWkovRD296wbSEAv9rWlOvILfV6cwa
sM9T6r6xnO14x1e+XYcc5EYAcbAgHVaNhPg053Z6eX9q9YnaC5O1GNwkVUseDpcQiw4/EvEbc8JC
S6qPeIm3PEVuQcfbQ42DAyoHTQYLDQQyptd8/zPgbEl0Mp6MYmL/vQ7SMGVKDTcTrsDWVE7/Biec
8ko6/c/EcFyIEzXyIXj2LMuCwznXE7biwHxCk3zFplq9w5sI8MuF9nNtwRFuWV0sQQ/SQRVejtbc
ya7exnV9H1JU8CNdZVYih2M+hCbO0Z6rwmyd2rBV9vl0YIik1LXKg24rHPhhKAmvSwsFoo8rsSb1
xx+P3mAL97DoCNfjXV1lli4XjPIDzon3kBy9kba+UaAfcumTaebL0Ytlvk/2+0Qv0seZWEjpJ5YD
eTu3E8QUpFvNQx4BW7wJGZD6M4+Cuj5h+EPo3S8rW+NycsRXnYNuJdqD8YAC7GQq9OgcIpiOi3HG
58/2f4w/DLYfruWYreUMiZ5V6pnQ0UNsWJf23CmqSeDrrM9ranHgUJHHmX4jPOPfiu/T29LRIFpi
cXBFZg4wPScHf1ki6Kk6gdiNOoF/Gk45qMfcsateBj3VxAAF1f8f+ZtoV1CfPb6Uoi/KLtXmMivb
IBMxd7uw35Dpz9mY1csTWBT9T+axZeY9iQ/1MYFXPoa6xtHOwHFA9P2G652Dcb2awVOQhEWTOIZd
mMhrJo3CGe/N+y7K1ok3B2KsnokwEOdFg0w6dj3JzZHm7+Oj0XeDvWBYJuiZhhNw146ptR3EeRlk
JIIzuWGvvZ6vdVtiMrbPhPia34MqHkf88bLczdrKgkPzxfp7XV9p1br8mVsv/jCsstuwSWPiE0Rx
4ZIuN8cbI7WggCEM5WBpkzVKvdegI7OUAgPjEF7HU8n/Hs0jRz1N1ERJ4u/IiPgTcixvOqKu3U8K
AKtOG+skX25jABJPJStEM4WmPJPAsSrybVqPdlRilqHr8rx7SEKcGGXUCEdTNRM05BdkvhN2Nebq
8/8sQm0K5gBRCq7Pku9Hu8dlvr1NzjDJv+z4BerrPF2G3sZgw9DSGMhReW+mK59s2iIm0scEL9u3
q4twuXLwjIo1UEJL575mLJ62Ij1WFLJVcd6hos4gkxEGZYIs9lOgxfk8TSKc6Fh5QU3vtZaNZiMh
yVWh26dFOP1Ys5u+dZ0Zu1rV8uEcdASSTqQEgWMhUFZIs7CHli6tkAB7aSUIOb4H2TU4v2D8uMrg
KXOat7SvAphrB5hdGbuIk69GMqeDz3qfMWiIcH9risDsjcc7D7Aq2RdBYFio+e9NUFApwLoUsmkE
bbpsCKtqj8q4sWermyPIrK6sciSJfAJMfNTSW/Rl70vNBdASSjZX2GQn4vpi/qSWvpQNeBEFBDms
PBWWLfTPm01GVQY4n7ncfMeqFRUmG4EDlFwjgcqVS1jJn7pY9Jb17sNSK7uHa3BM7WT1Ev1pfqGo
5e7dQ1/m5yVgTodekFFd5Y9RtIzs2M5E0CM38ecEV1Fcfm5Ic/bdQWuDHo8sQDSmxhvxV3yne6k6
u5BgIPdaCiw+mxHuhU9d1kdL67uqNcM5eTLMaKeLgfrU5fc8bhJZr8sgiZHeoZwR1c/LoyKzyTv6
Q0i8+achnYd+ZcB1s6M8twcmjCYtFLoezUzyetL0Jc+5MY2bC4M1L9p4hAQNBinGCp3frWZ5Bqfj
V6fkX7+2bIQ41s5jzgQYZDmMufVGhqexc31B+YLrJOBrYUkjCP/4vWGW82wN0khlL8LkCKJH7zoh
oLrpsOb1jwsr8CyVvsdhLZDFojtfGQbly6uheEoGYmpjWXuJL02iXEZVSlpUgLlih2Cjy8UO8lUU
LNrug8hy9O4R/+h1TEjCGwxQDEbfdqg4M5cm6SV5kyU8E4HA3K3Jyuy9ee/bPQwIfvxEhD9YjkyP
T9ciVUofG8hBrV6zPmSO8eybImVDV0TQjeH2+XZql8JNPP/6VnbOBr0FmZv7M/NPQ5RnII7O6CtZ
1Jwt+2LgcWSSbojtxwEi9Uw0hqR9GJyXCCnP2oDjEpv2b4iU8qkxbwYm6GBr4ReX6iI2Okf7NQKS
pGJZjVZXbChiqcDbLy0E5bXQ9t/Fg9NTsBquBg/ZmkN1kj1/kSsjyuea37qV7XYzaobTqIcWt0+S
BSSWjHuYxF4btfbxK9MY8diSNonk6VGUu/WbdKFahyw0n+QL29f2cKiNXn4HYAyUBNyWy2dI1DB0
x0ypaQEkaHeVcXZU0YE+3edVZBwdfByj3rt3v1Hy0silR60NKoY+i9SrDSaauRSXaF06P0meAInO
Rz1EcrIMM5+KXbu1kwlmzErHYDXj/hQc/x8qnOoqPSBjRZD1kZXuH2BkQ8pgjmMfcmvjJjk7fzQN
YgP+v7znq/YP1YbsJHywO5/VjH79Xqaio1brjAWmu+Ou0VW1bl4yDx9GOdNU5el5A3wWwPL2IYOf
ef76egl9qucI78opspdZTSraagMxmdqe9u+AgaiVA3i170E9RCI0YWHlSipx4Qih9tXVFwk9yTtE
YHhDVzw0Ma0EDeQY4a8yJY8LXPoOUxYJdnaSUY9V5I2cZ+QkotNNk3yYSWqRqxMqqa7NkNmSczdw
6KxOpRqRp9vPLKkXS0j7biqxJKdAuB3nk+ZrUSd8zZ7+cCmk5xUxJIsrB2OTkbFn7Y0BN8PHkUNf
xZcoXwIBa0Pr4otLMuMMMAMozASuSBnWusq/rMUOUlyfFKKvDxtapDOMby38t1jLV1P5l/UgaLZS
S1OFDhr8WnQNBNG1rprJfdJ89XxxDuxSSHQRx0Ba1kx7ZAmd87+774G6vqYRitx1k1n3ltbpGHdL
m9BqtztgTKSUmruC4txDDIw2LbeOd45QaF74m/ilKJIycRUzGQZfJnZjmSQaF0E2BHJuq+vzIG1v
8U9Zh5wyFpQlpRubEI3dfxnDoGOe2pIrjQf6iHkwFw/RV5O2+Eb3aNjMNMUIaWi9qSBuLP1Vn9CS
1rd6a5JLiuNhEtJC1scE6OsQpujg9qC8AdVUPymQ9rlPdz7a3K9mIc+CouaLtq2DH/SxafOpOPOu
T2W269hsmQbZgkRp4DotNYod/K5t66Y442m3LI5Ujg5fL1W4RMkbbF6P3Cg0Fw96UsDnDj3mrkEj
xFYvIooDlUh52t85bSOfecCJUlS5Riq6QXcwM2QZXqRuqbVFQ1mIVbfyJq/wV76VyeYlX2yQ0nb2
yzhOcN5ZDrwgb93MuI6luCaa6IFdfkwTptcDjYhLgPTJRCxYu/3Lb5CpMD6y3xcNzS3YMKV4n9r/
fVS5OG6851rKQPpQV8GY8hxQrC19/a5tCuzZ6gIdVdmRocfV7c125PlEVIMN+wFIQs1vdp3Ynt9i
LVwWTnZtwu9Bq8n35MDfOdDCaO2/mUnOG5PovPt2aqPUcrgHucBo9QwiheOgczjJ78vfej2lahWd
JKGSXG1Weqy31mHTTvFC/I4oY8SmUrnYCv0/R9HlpJZAwaJI0HxWHEQqbWJj4LQnU3cG1bgCFl4o
jchhOm2VezYL/PG1cfuy3I30Sx0vc2P9aoAhqxMiHRMbmOL9l9jf7QFhTbHyMgls5S+oNntw6moL
5iAAxQR3JoEVgcsS/WajpjZgblIXJOsdUuCCR/CAYt4K7gsSQT2EXJXsUAkJA8mauLFAWPespqVZ
TtNo+M8QhdWGg2Fh5aE/U0fUCA6b/4HMOUPQnnEPHNA8RsnCQRBG34J0A2wsynXXmpI0FJm5pUh8
SmUJBCPOpFUFamP01PT+Fzo4GClpIPqm7CNuS/V+kGU60z44Vzj7QUQVtiJghbfc5q8BWuybkxc1
vsY1piZAiM6D3ttytJigc3taoIU0WyxI4KLFa+JK243e1SsMmT3MQDYoPhza6lmRyiERAPS51fQU
kP+jity0gNbzRJGoksI0x5kc2xmlKytxQ8XpCZ1YW9OdOlNO+CGApZHHHF47qQeYeL64SbHrQjhx
Ud6GD2bJtP5TOQLtHt0saFjXO9Z8fBWarY6rJK8dKoi7hSh+DeWrrCV8eBe0CAd+gJz/HkPoT0AZ
W5aVecygCXsIwDbuUneX88r1DhsTjXNMOROyU6cjyyAmSn/U4KMF8jmH7i4CMaED5OTUePSpb9Ia
kfH2hyDvaowTOwCHdgaTDV2ppxRgz2QMNS1F8qazxyMxcHOS0/FxyJkc9XKOhfPozegTPrGrFfrN
DvLd8bjx17axFCNP+gq4YJPPGo33Rl0LItFH8zpGZMbVZGHbeFXkAJoTlhECUj6OkUWZIHIiv1Dq
mEO5hnRVGmtP199jLmVOCv4AeiMThto6xpmrx3zgjJENhogvTsiUNJi1g4uCm4hMD/X9BO7mhQ1M
QxX3v0iUklqO6vYmdX+g9VGA9CbQ/ssrP0RScnpdrrhl1+eUHjGkzta+n1rmaXcM6YWRpou5Vckr
za6+LZWv00RdXTd19jfoBUoh5vXJMT0W8JGyk67tazN1/15JRedAyXsYjLcNZT7mIhQ1nH0uMJLt
ipE4SQo2zZ0/qGU9zkrIP+ZRpbAw+TiM/TQS5BuWR5nyscohS+oQGrKt6GJKtroJ/2SgmYdzUTGD
yrySHkN4Lgu/NCHfdv2mqoerVeu1eSZPk+HR3JEj0VOiGpEIs81KG1f2d6oxpx6rrWnIOezV98im
yuetAZkL2osSS3XkRwhGfnFKVuYHpKs3wZX2dQHlk7Sqq8xd7GX54Xz5h2uprJimvopKc1lfTIyj
ALEcwVYMfSfWHA8mkF/lkKxDacjM2SSwfzhle5ZBIv/Bsu6ofsf79N7mon3rqeOBqB0PKhGBGGUn
1sJfGzI7+Xmq+JAj6jZUtxVwlcH4ioideiqwnA0KMJFS7biPU39Sycf319tFFh7RpT5phC5ajnAM
0uCnxy6tOKzegaMe2g+t4RJHn4yye7LgndZdC2+1Cv5FPr5LIKYTRo75y1jnWH7Pz66U+B7rBovd
8hmpOmIeZx8hbpwnoYgnrYrrSwJc05qymGAmEnqHiat31+JVKgldKLtJnV1We9fsRDNPXcked2XX
zFneZRkLzDcjsrA2iU25uWU1bu0eOnnn6hww1aHBZScBx5+XsCMlUWLQP/3LhQCp8PgswVrkegt2
RKy70EpNskVe3gWAgebp0xZHzmy7QeJU8GatYHWkpE04bSB5IkJooWqR2SuKgImN8xfqtKQ9Li5V
MJvvXRHyB/goVCuR+AQ8BXLWm8eNOPfkSrPpSYpAemgVlMyA2qt+nF0ZI7qZEEiHS0mspOUsYs2Q
WuH6T/R5UOtxfmQ/l8rm4ptKM7C4pbzlZYUJ0rNp/yCjklhpQb9VyfUfyjebmBCh27+fqUU0aLny
JPgJLkICQ29VpTp0QhKJrgC1acucZ0ISHE+EjHynFmbJy6o9ghIbBvAj+w5RlpcaL1UmV8Qjf1Vu
kc46+JVJg/YegF8tFeYnPzNd6yFOPFhcf5Uw9RcxQNIZLZ6QO/nKdhuiKjDedDoUag17l38/pZQ/
R/nemDMIDelGRi1PPgekRYNC8j5vC0zBi3FpoR62pIDGBzTNLIRU8IXHfx8kav3Gq0eB+AwZPAkY
NMoPRPhBACnrmT+jLEP6mM/dDUAfwhPjrgxeqa7AmegScawZRXhuYtxYsVdE6AjM0c7fnRWlsRl0
nQuW4mP5/h3/67+MRT1vik1INsrBKlqrSoXclAsQ6SEuFGblf73eLa4QUNzq+rAYomxcAIWIHCrH
q1eWEhLZI388GVbfq/RgrEnnLCsFerP9zhINNtZ1p1CXIzxlLCm9Sj08Agyn+6tB2JCdEXLYdnuH
zLiSHsroyuuiYchkQfeB57LT87hLpiQoTan3nZ2eufCPFA1YJVV96G7NPHS2ef9uB1Zn9C5qKTfx
P5wLQ3Svi6Rd0wrxrDgF7YkwsxT4m80gD/SGkElEB1Vn3e4E/4ESjK3yo/obBXHJCEx5GqsWbEj6
CBYZnXDjoP/HwitCNX5yy24c42Ui56WCgHc4C7pn0ip0ycMkiHS0HcgAmozLI810clWgAQiXvl78
cPc85jHPWN53VG/GQskWDp9xVAe/+JXqOJPTeTNcFI6uFGFaydJ875OOGHbBWsuAu219Fw/TKfgX
/qRGBP/7KVuymhBqmuqX+gkZHSIPtgLZ2Z5zx77xnqYCB57adhVMSuEoMdrFLsNE78m7crSXiOJU
tB5z9i3KW0DUPdMjX8PJIr7meu/mndxAEP7XrOt5SyJsCX+57Z/yOVZ2sSZGZ0n1QzwsBX77lqGS
3seNPYHVP8gDfjg8b3Z2X4raWk/yoSwq8ULOD0ZWCaFJoQhz23eF/BeSNaIJdtyUYKTw/V+0ailp
KB+Ixlu+URr+/k+V/tDHyD+DCRsG+53LeBupPjsdgSXgMPvdoiKhNvIHacBnqjUqxg1gWNxINK0m
dQhJWcdNVDHJZj7/AkVIA4gHfy+m+4gm5xEKW2XpJLov+TFS533iWDPe390+b8Iswowc6Y6W3MpF
RvcJZehaz9kVKzDxPHuEqClO5mXWNp9RZAMiNOth6GVoasg4oylySNNxeglnHUAcroS/LflyOuxd
by/O3+1XdGnUAIQ1ntt7m3vWlqUFuTpGVHsMcntOuUYg5jRHMsp2UiGewFd2Qyc8wgrhvqpQ0b61
XhcK0sfPlg10RVu6OZJGzqNNtjeuKWwsqKGS68peBZeomkpSH3BIqahmRXdgM8IuqZmGg5KH7mmT
2gEXd/AD1ikgkZj1pZqUrOyR1Oxcji0TrMFiknCOLndHpEDFInH470+AnYvjXicxaIRS8BwJfvYo
FztRpY6vUrLD+sPLwNz4hkSQXPw2nUUtbhX4dWLuYTtqzZyDb7zAlSCxzY+laeK0GBOl5tRFqy81
rr989qm+RN2KHYeuNd6HGs/hks4sAed4nDdhbxmCYGkppvXZZCFpNssNhIUGpV9PHKYsRJkPlzTI
BQodrq3i9rej5Iwe2kq6QUWBu1RQv/iY3ulzXfSP3Fu/Y/UHgRrSqRVma9yciayg8CBXiil78G55
BLm7KuvvGjRN3TRJbrNWxr8LtbaKpWWGNoilyygjrxv4K09svcimDVVZNCF28NcfkIzjbn5sWvMt
AicFowlIliVh+4PpNtr/VAVwTrE2nLVKopIPxgOtDUzROJ9Un/6y6SpLpMxO1lpDoGvZmaUDTYO4
lJ06kaj8FrshoGS55SP/RUY15yYEyM2J1ZjKlJrRJuTiM2PF/3UJ5F4JhIco9oPUdq4YN8bfwGaf
l1sYUc1ny6Pez321XeXT7MG+eCRn1I8FpGDp4RH1mc/vKk9ozb/y7W2dPgQNC/0+VvFog1p7O/3O
exX61ipwLPl+KkmW3TRsqEbEeRdnLviv7NPAIomuEKkcDXNIKcARvt8Iq6VaGcK8sGgVl25iE9qM
k1n8P80MFQLs1KpsDt4Us5/CMv9KJB2sVSACpjGEQexR5mdd6roaZJC5wwXB2cbRn6gX5GIWTbSl
WfkAh3VyRKc9IyRI5GakWe49mp5UugwqZOeI7rFYfXFs3twzGpalT58yisDEXb/mxDNCjURBHOfC
o0y2HeiDwbabOY2uZhP+tkhLXAXHxsLR7SQVPDav4PwfANUB8YgLPgAj6D5eB1/8cMGf0YyQzdAd
kk2Ez/ks++B7f37BlW4Kl94wYfrIGLCjMXOjVSgcnj87MBJj1rD2FwoZaqdN/VTgN/GlIULI+1rT
2BGfhwjgMmFehos1cFbwMJG9w9m7hfgbqozsBCZuOgT3NXEJ6m9nHe3YJmD6EHfKQoeQUOJhFZtk
20bb6E2Z9AhnqX7wph5hBT4YW/NSQto5B0Di2tsYyuRo3wGR/Sd4woLukeKI3H9G/fcsQj/8IonC
fwqjJs6u/6J3AdNoh27H0+HJyodqhFr/k8MouEDZy4J0wZhe4mn9jF7SILTq+0Mfq7fjHibcHeSr
R5tp2D9qFS3bcq5EpES1LHzdtQSVLzPIT0NrN8IFdzOTmgz0zjY16AP1TdHTjKAMw6YDxYlvMSI0
UQJa0IHNRppAzNrR6wYi2IpGCgr03OFJauASUVtvxgxucdUSsqGopc0y+eptUrvHkt8v0OjLmV2i
peHmW/1eHEPclrPkwMiCCs8fywK8yZM4cNYyWipA0KgERcYmoVJu42toBlzKs711eQvP2ZbxeT+5
Hmo9m2qvpevBgMSO/1IkTS1Kpptwf00AMQzgbjhi2NgU7TRsO2AgRNLoFxLSB7kEQj4vcb4v0QXv
KuiSpVeYve0kN2eHvUN6EVeaexvwLlGcZ8m4lO3wdzlU+8H/1NnDd7ceoVHdc4x+oLv2EUQQM5kO
IHRSEiSq8n6sIoCAK9b4vTq/3JVV9kcl3dU5dSZxluAsyMoIkyeTgFq6lfTOOMhax8KD+Lh27VoU
OkXTmahb94Q0UR0Zwl0JiExIYyo7UVsrH6E/Kkrc97/0nurXzQuNQ93MXC0z2hUs7+Wq3lLUWL98
bvVjeL1e3sCFIi3D74j87J/Eq09tDk7RWAMoq8c6hPgFZ7+frJ1RsJQFONK4kIVOODJ/V8syMEoH
VZVujV6yFMb7jQly+RIquOU7VJH/nDaJ7nvaCr9Tc/8u2B+1i6wj7+o6C2KLunH8tew4tQ9Ln2nn
04PwjXOeNjwDTyZt47e1CYajybuVK2assdBG1YyfJkmCeaZprTUwI9vCJrX/arCyzClbr+D+z8PD
7oQg5m1t02eRIV/lpCGbCP5oeP97Ag6A4fKFJdnTB1GS5fF+v+qIIxLgC6HzeESFUgD8Y2YEGRMG
5biRj5p+bbo2eJYX9fxx+b9zL50BI8z5i2p3lC9rdEt1vkK77tD5J/OgLWz+HVeiE78knUG8d86K
mxVqhrHQEK8dIyzF/265bwEnsJC8HCzpAQkOkbcAL42rWSMqA0q73GwQPnQ6D60x0/MWXSauzu3D
IRhNzNU1JQwFF1fHJNDcRCAWHVRJA9+ZHMn+et5MH1ddMbbLBIQXrNi2bN2JRbi4PWzLxLeweSok
HAQsRXnktWyMgSVNJpVDcY9gB58qBNqehQb3JJ2H+vCiE15mEMU0KtTWNCdfwfHthvhuf9VHdoWE
4brOJNWJsNX1WKOgj3vCYIc/dZhsPVvq1L+hR3E8Vt+1DQUb9L76j0KjdX0ZHVUv5w+TlOevTVYf
jtleWP6tmiwiCsvYlL1Rz+XFoxZ+KWV9wLW1U0DBY9bQ2vDmhaG+eocRS7Ax7Vq2U+rxYqueG3rW
mpMndP4W+rEz0gyCmMKdf3JQY8Jdx6czdtVWtQBMoKPwEyeAFTjEUi2gJikJI+38COv+5z20zbWC
kT9vK7XSF0/fJ7KD6jxH1RqpF7f142fM5aLNyBErPEozYmK1WFnTgvro15ybH1Wmcw/AKiJwecqg
oK3jYAhTXfhoxQkDzh6i1I0gy7gQ62cdCFQ2Fp0NZdgGwwMFLt+jcdeiLCvJDnrgZU48Khamoa1z
IIjkg4tftHJoJIyarsDB1Z4+y9Fsf4Hbwg6Z4ygdXLZ5xh8Ch7jkphTnoEZUBnfySRWFJczQRljy
qE9S3TMoQtWJxGOP4gqkHm3C3slsZebac6GpJrh5N3sAs8o25i4o6kVNdTkRC5v4wZKmXM8G9zr7
5LzttAzBrbxR95Xiw09DI8tpcGa4XWIrH5mos+K6fHohciheklYCokLoFCXNxqmiRhSCYQf4pdis
zZaCabCq5njd0BLS8Bqj1lAUC7idvR350lfAY1IpfAezbRLKz92yPx01YQ0a4shiO6CXhb03ly3/
xVsKOhnYB2CHK3Pa4YTCKGFppqvKHqSngY4Gbv8og1ArSik4wTLNmSIS3pu3H6DLPuhIam4F8vma
QsCkiOW2HIwydsSb9O5CnhFkklePScTC09FOy1G0AS1cAu2XFVHyUfMlKfWhKCwlAo4xTlkw+Ojd
63wbPFZM0UB/wspqzFSYs7DgGbSalJEZZ+rMPiGtJnl6YR2ywwP3qMMnAo+dS5kRukHhXSELdqlb
vAoh++MrI4ANuBo2x0lRCSDphbnHiDH3Xq+vax+2asZWPD7HxXMOvM/XWxaLHygSkNacxsVy5qVL
Llz7p+DNdqT48+jeIamkj8YjEDQ0yaFvmol5J5MOX77MjHNmcxjuEG5G86N6LaphSYDbA+qub5G9
Ty+eZ/mDEknIyHFzQDbFdtlsGGEtNOJtQY/Xc/Xk5Oj+yMT2NzNFmvKBmiqGZ+KOPmrq8qUWytjP
flYPILPJUje3dONFZwKMtzdk3veOWn1Ly7h3XFT5tSHJyzMWF/6ixPsk3kTvlUGO5EfNR0OkPewL
WdcNDahxh/vmD1GGnnMMgGd1MxtK+kCc0aRiSFRd1YIYI3ruViVWXAjQur7PpH1IyPGlfzvEEWV0
7CPb/IzdSsUrrG9Xa23fQSRxyDR0osOGL+jx1/VLqAd7LMnAiyxpGhPGum4/hcHeqLRChrpK8WfR
toHaXBqUfQRc7NRx7/CLAanPuNB99raQ0id5EqBuorG92eWmJ487xmtZiETwHP3BEHus3uNSjwXA
/SSwff9rABDrSTQf4588ZDYvF8B1uGERkN5ISLayZWG98zUBW1lqbsgW2cWoUCAyzHixA3h4BJvh
NmufjA/7hFywwFNbZTSmd+UOGvEnXSAOweSquroGqKifwpUtGIsygY4Kdo0sYCuW38BrauPCDJmG
vgIDzbIIc4HIbmpLQR3j5UWHeSUGy8w5gWdloeczBbjHWKim2ZsI8g+1Ga3GLoyy0Tez2qJiHcSx
KYm9/L/Ca5ST7DPWMdiL6dKiGjRls601qpwK8RK73zL83tU4YKoZxeQc0VzBEvwQ7ZGcADLhoJRX
zrzqTx2oigVdeGP/mz6fs90bFepHTypVmhaJahLs2DeLYtA8avHHzqZtwFlGTVno3MV+WHGggifl
NV1f/175nsCqXK56pZvgtoWjtjesxq3IFoHUJZaWYGHyiIZuLZRkBfSaRRVbUAx3mlpkASizz9DE
7pkjbmWoyBfol0yAh944Sr2iuTgh/NiCN+bJjwoHqE1gp9vJPQ+Vxh1sgNwisuhDZp23N2pOShuc
z4HgQzvXhu2tXcuHc4T+cJtvvGfIN53sk9Zgg526xK2XaZsGTSdoNakmsJYxkEwpGg16pzUoFQXB
TTcWdiSg1GMmVfXy6NlzPMYQ+H+CKCFrYxctAsmg3oYv1RSvuoM7F9C3k8nNUSbHzim7DXjR70lI
bQ9uYlDl4MP24nW8rpw2XUQnAcj7ONEQWoLCxkW25sOIg6TTNETEu3BA8R9KQpGJbuY/n7Zqib1z
R3oxzjPbAS1O46Zaq1bWLrzlNvkkRMbovZ/6U/0pvzTWo8FSKGAjq5VkJp5t2ekUSa7nxARSidLd
PSKe4qcYBVspYuM5m6aKWE0hl2f+8rpY6o5LxRB9D7dujW/RV4YxUzsllr/SjcigY8kh2NUd1A9X
kMElKzdIxtS4NzUmlGCrft656kL1x6nhXYlkGzFxjlY8MvC6TLnmc8a7vYCu9yEw2DXRDf+4z1f8
0BEyfr79PKV0D6X1DbEtEir6j0emenADn09lGD3JAWZxjhfIFEs6udupN4SHp5ly5nPkyKnLZidC
wGblDNvRxa93u4SJ4gazVWYP4lwEktEKhivFOJtSHtFJWoDoAgTjxbhHSLNc89OdsWIfT4k40JKQ
iTEpu6YeV1wY4jzTWDdLZS5MTICrXHOv7EaUynmoEZFqLADTX+rtSoOUcZFf6B71YWAc4S4ppohS
sgvcTUmRETkwd+IZRPQT3BcDuFXPQLivTyoIRde1EKq6bfNUjS/mmt1f/l1EVI0zrlBI/OP0dzCk
CaZPKsJOFOVbsZXsss5BjI1P/4dykH61PINRjviQWrtFzn1q/HTojO+R0a8wWjJjnL/WpBEZwpxM
dqRbqv9uhG0yXRu3Ss6bFiYk+XqturQCdfMT5FufuLbJtufD9eRybiXmESdxUBtsR3RVJO0axJwe
6OKr3Wh2L/Q+ZVm6Wm0xlecMWbb4eZYBelxacpo7H9O8BTgnzp4nM35ru9qTBgkglmNrPWrL47MV
PqLCjJ4ZvO/INZNCNutfSOpaAjT/STuLvfmBaz5cWaI5+O85WVYxKdMRENb/vz+CCZ2Bn5bPqtqR
EFYfWfov6reg7oBonI/F9TVzi6ReCwotWCmnAghdj4hyAzmU5cpgDm/whZ2r4zSBo6+6LhuIcGGf
6Xra9Des7tQuSoXWBt2YVe7K2pw87BWsSIrPaKj7rvlaOaUmQVF00N0q48Wq+UfqGtA+n7gHE7GY
SsWm7jWl/HjWY2Or2v/J7+ddlSvg6pDaFN1MZQVVRrs+zycmzQJDwWFgGUMZdDhFwgZjir8tvzuD
/IvW9cU372U4dOMgV+mMPZOXIfj+0kJoRWMR+ByxTrAekhdS+i6PY4sIeXqADYNU7JnsLLWoEX3u
oHr+qyihgtmcBoSbKWyOyJHik5XHj/jwsplR7E7D7+W7T7apKPDWCJehztlNBy+4kPdGGaZ6Zvqv
GMptqxcLur4SdTUOriPy4sYaEq+F7lDvcjmLayrz1osA/Gd98elgcGc7lBTdmb8mrAAyBYfYG+f5
6XQg4ZOJRCjA3Cvs5R9TDgmhCUbq/ual2GZNj4n50bdeHAQcshklMRuynNOIeJrh4iHQQzNibg6b
ifV34SvYA2YKul9Qco50H9BtS730MpJMIX5rUtVWpqPSBEEH78Sofqmm9U5J2Px87p4hdZw04ye1
ltVD6Lof7xHMDhzeu5rHb/2gq3q+HoThN6W/o6dcHp7gQQbqE2OT4Tas1LuTHG3SYySWl37ZL0I1
gqJF1BYvyKx8CWCoHWOe0wV4wTcnDgzbyYx8sBS8DPSIjdTIYDLM3kKHS/KPJAl+tjJ5bt+6XQom
dAoxX53c79+STtG6kX+RXPVBVVt7Uw5VmIjhBw92gN+BWuNi42jEifuSO/L/c8PAYLR8C5VfRi/y
42+mCVWEJ6NpqCUV0ybOTn/7eCFfdzrotTnclJIPKW01eolRZE21Sk3kbWM1UsyKul0FwGMQffPL
T31vtW6ZK71vOyoEwNCY+no/Z9+muLNEYKo3+488kuWVawTYtDmNw24uq68c02RkJwKxb+2TY68k
/fhcz96tgL5kWyu5n7xTjQwyVfO75Wd9TZe1Ru4Kfbaho9sTsyM7/qV7jj9rwdB6UaRMgufqbkM2
OfMJAtwcA3EOkE8DykEF5+tE87Ru8xbbfTroZbp9/evODHHKLt3NA+bbP+yJ4/xx0/ygNrZFKM3G
XApDGse7+ZZiOPv9eMSHrRtuXnYOBdfWEgKUMezPzm6qlv7dA95FPwGjMoAaq93LBNTQAEQYjvKS
UWVRlE+lhD/38fLCe/ueyZU7h8A3pW5JCnGZmsz9nafhyRFo1jSOcyap8HMzKFBsuQoRCEo7wycj
7TyPKlEz/Rl6CGtrSYQR1Vmg0UliLd8QARjlB4r2kENbdNlNuSArcdYbC26ard0naIJ2EQXDrNL4
uumXxK9C3nP6JsxgM5RMm4ig1Xq+GD/+WO8twvxmdv9NhOUHHtv+D/mKQPDjju/2hccXVheu4dPI
sxb1l8wpQ0xd3WC4nEBq+d0TTVacTO3p4i8ninBWkKGjOcFGWs4qjlc4vUdE+kWAYayRiUR9/sxa
82owqSz+LvJzOJTfzp0wT0CRwVXemCxKNJ+vhol+d5Pw6GOcylDmlvhDn3Uz6xXTsIarE15ASCvg
5UsdUpLXbr30vtR38SG+8vY8vw1u9MzU9pN+xNo6Y8Uzk0Z+auNhaEeUfyCnDnoIqCK/PIecdbpG
zyjymQnwsve667ab7SGKyAB7yKNyajeldWElAADHVskfgYnVUZkIN7Ami7yB7lOpIs28Sd60BN90
hvxk6+HqIKKvLaEne5+XpNXIUz1QKVvYbGCN8u8zPzm4IpltqkzZfaETpw2C+84+WifOVnvn5hn8
X5PJlICw2bxox+tjxHwuwYE5XAGAJtwojGCjimS/4zOX7fzwrHpOcbKNUagyZnO5WEqtsjUZsDAa
FgALEKPmna0z2bePkdmAj66mgpZRlmdvV2mPhs9YgQSs8d6sAxMi+VVQzwH1OigN2H2qDl58S8On
fl4g+fUex9k5Rr+sotNFMIgB20m5JXFF4Kp8v6HQa6y83HIiI1XQp+5px6fkB0A9s0g9EHCCPai9
AtE6WDa7DHJ8UN6Y05p71NmqZecyEOULAObALOHkIynF8cIScWEeaZZ5W2blvLNxpZMeODSUhC27
D9FWtTYmqj1dlJIwJYy5d6W7N7vndMk9j1bwNU/aYEgamdtYNOuBLUUT+3hxlfqiH3sOVbMd9jw6
uLeM3a2BQAiEd+y+vseCKKxHyeWV+VVVQAwcYl746+hrnEjUl3TCJFgzsij+560d+TFCUam3JEIp
FPhCxWuXbUvYfAJWVmFGUf1gOioNa6i5IVGQRHiBn6xIqneq3Et/4DrQx7bXAbr8wPA5H9HZ+zEV
KOQbenB8/Rf1Dz0Kk+fbluPgTw8pfsrKETXvbMDOBwQbl5anfTdHLRAu7U10Ov4VW5Oqtssd+NTc
nb+ZhG09dTClXC8zJ+0s1Sz2hhxajbFCyVoB4LXrlS19HRZju5vN5/njp/d+KB7n15Bv8dA/kERm
Yz8FJ696pVspg835wZ3sV79PXXThCZRDsKzLqidA9CNl66ywj50SwFNp4y18T3kV3NEsVGpHSRhz
gTmVieeZq5XtguLW6P0ncZeB1PkKFmlFVQuhYfqS6qxXc9ElThbLP63LKwkyGUTzAayneUF/otFd
U9wSINBjNDboJGAmCzVCXBnIUu2R+X3CdvM2kiRLyNxKbRqPHHkZGfZCjPjiQrM+WM1DcPPHzVu7
+u+Gll8qJVHQAVFhdwy3eqrSzgOwgXLwVdz/Aj65g73AUHiLxHzyu1b6zuE2wtNxsnUOGc55gFqd
ZWKUmHdIw+07QlPyzHrjo7qsvcKVW7YWsd3cNx+qD5nJszTx1DHYFyiW1S9JZpUuMVX4sRzMyemn
HQY9faLc1544QyK51L6e1aicoeQgfpsjG1jy49Xub03hFL8WriJK8EYvJX3WHcN7NRlN2MO/Qjjm
K+JgK8lzhpl7TFEmVbo0y4+OiIRBqpgIXer4uEavFNyxO3MmyZieTJdGZb7eDjRGAq/O0L5nxvby
V530nLm4z2OSu5eo6Udn61gfYblw01M+4wEUo3BS0+Yf0xN24zUgorb3h+pKGvBpaYzYjiZweUpE
q5FL7vgKtYFH3J5gPzn1WxVhKTM+Zm5tIg/OENDawYE4A8LYsSL3YQlp2gi8okWJPhKwwf81xtUS
6lcu4T4FdpgTPBvjHRBqU7b/yraYFJ8dGjEs8xkCDo86otbkoJHgO2lrn+82CrUV3GZe2GGhXBtq
l5EChorAr1paLFH1XETaAkupSYCIJPY/sD0HKGTCogmwbRiBuS0JteoAgh8T/qX6vw/eFJtT0gra
QRRi5IesTmHlTTUlFMQaEJ5VbFDuNevTcrig5nYsdb4HgWmvd05WmA9ZfxrmegiBTZG9aEatT1X+
HRCx3CKBXFRZ44xeA/iBWEBeitncgZExFhXD7AvSd5hkgh1vZO6Wu+Hi1fvtR7gUKd7Dsld4BugZ
mCFSnD8F8X0DxBsp+kVSlB0UoNMegy5Gn0RJNPGOKpA3ekQ7uhVNRtXF6gM62Msh628Ja8TP4BRV
EVkPiXgJ8rEhWivkj9H2eMXWoFl6YnU3oSDSP04LtK+SCnFZFJEVc0ZDE4ulTBK3rJNex0TE4ybN
7fQr3Fqr0/HDAkypr2DCkZu5UGLjKS8iISBDEQ66tbMv6cpp4lJErUk5dgGdrrdAqLIS8qDcYnnI
KncbTBIzTlx6DoB4wAyB5j5hhMkw7wIlSueGa1pFezePrOiuLma2Uu4tNPdrVAwUnim2Prbl0N+7
XXD+OUnEDzZbhK7MN834kFMdHAHzIogL6pQvvl6lHatA69oGzr36zDJk2iiqvm6G02+swE5pyfWr
WvUDwxcvKSRNnEpL6M0DWjxHvvSrN+HftO6e28/q5dmGs88PjrtNvCW/ZwZDhuH26PNKLFt1wK+y
8GofI50o5/U9lnBr6IbG7iLhE68L5iudbPhNStI/bRQHf5vqPzeDET34ZdSBTjy2uNpTJJOM4Z08
9s+wQHRzwfqEVXhGF68ILciwm5+he1aXXa4xHs7H6258ZLUxF2ZNO4Ll4QChCNoOBI2cdmlv6AAA
LhgBkJc+lp2U0zi8uGmRvjoX71tkNGjVVuqsTJxRm6FlBR7FzS9S6ZdRS86EQu9albZ/g/bUzgo2
4fmNvtrFiqUC+zrl0Ek8UJxzCBRSpQxy7UrBBJj/YWlPBYB7xsaDCwiiWXasx28SBz+AIzLn0f9a
3yiQz4x8wvwCxjOwUqN0fx0ei+Y7PI6DVMWvnUSlAT5L1u4G6SV6llEGOSZI8JZS4FzXOS0BNnQp
JpMG5T25nXnQJ1vLAJlOoVmcg5E21V/d00uLagiPhjclZ+cUvw8soSW7l8Lb3t2/cJHrYRXRKxBY
OyfOkjnbWj4Zna3mZQEDKkfpkbyJjYT02U755tv/4M67276DvGLJz9yiV8elycQtOFkl8P/V5z4o
TGQ18hfxwuuIa8SC9tI6QYkMtx3X55DGShKVJtiTrByR8hRpIXPufSmfZSW1CmOVni7Iv+dWwMxX
9Np5IWk8Q69Ek3Xf6NiXdu9bmg+CgClxOZz9SJ/TD2oZSOlGkWvcQWTe9b7Wy/RXvTfNsmbSOU5h
J17dqpGTqNF8kh4388DHzdgTJZvy7bM10fJ90VSn8uy5AP+FKggmJwbzbcaOJ3/AvypnhgYyiLe4
hxm4nCvi4iNdDmLzH03lmhO8quF13yzOZxzDE/rd3p0LyK0ujjvM1ktr7uXyfhs1Z9TLLO05ouyo
tW1NHehJuOaXB1ikroH1kqMuFZm4k3CaaQ8W+jyITkEflRhlrosRfA/t1zOVTmAzBKdRoJTPMLJm
nQ/s6ugzJAYoEbqRp5bGFIjmbTnFKRh4sGpdIXwuLErIwNtjuQF0WHPI3ErjYfvLM4bYnDE6kprW
NAOKOw0IIdcoSIG5BbZl/7p0CkCEOjDzZcdkL6LaqYBUT68b1ISNnyuA7pLHTrRCsHLubxUyyAms
PIZHiunPezJ/MK3nf6hcUC3ltFiBgeLNespoe1NpsM21psDJGBMJkesrPDDwfJ8DikHWgNGSiv1J
HP8uJJQ8C4LJu9swWCTTo/bC/AjuN/iUUf2UtrXzuQNoSiRNyJZsanERAOrJkHf6gOpJ5PTUSnUO
ASdlL3+Sx7bbncmdx9rH0UuS0RplzVSWONFYoE7J8RvFoJSYDVU1At/uQkXVcIMUZ5kn5RGu8eD9
LsSwRxeRKOe+Zw6damhpL7Vn6KxXiV+w56xPl9AQjldYChRXGsCIjK5tKYkO71exzrSkaSbHI2DS
GYeAhfJbYSk5RCKYyNl2J+oT5z75OUyE3iKLpCKPIWCQZUmOdmM8W0LBJc/+2V3SWE1xau2EMBo2
fZFb3dbaVWQY/n/3nLbgOaCruBCG1O402tZpZofM0EnqoHDS0wYznotCi3hwm/3yxpx2y78NKpC1
UTXPBsZAa1GdaSXYBTv60Rtoek9IVMogD/2IOIU+bEZ01xZ5/aySzXEk9txbzJNvPy58L7o9+sup
a2ede4s+WLrbfRTJlYHA7O0BlKMRsqVIzaIWnY7aOrfBju097/IgYAEiAIvxWJRmc59MLzd4MAYR
4Fj27XoZ6l2fEs01OFHeSDARxO/pxIFwIhb22CGxbmwRz8lefaFkTAkNzSdg/wxMTCobd1CL/pLD
5q8O2rLYQJQtmxKuQWTCoL82nDJY4oi2qdxY5IH6haGLeWNBdDUsOWXp7n6fY54813I3/RqMET+f
7hE/7Ge8GFZtOEf3ihieBA/qzRynXn238sb0ECm3j+yyFzIrLPAonNVUukGtgBx2Wkij7/8CY3IF
ABEvtGgrkug20BT1FgL2XMBYuOFhofW3a3cYbBnCvgO1O2HBRLtEvDbphlh3TxqvBSmNAvTOsJ2k
xIdH309Okv6bNhrZNKg4AFPYdgwj6jTneeD/YxKkrQFoG+TAShg8wbMfb6sqXLyeWj3V+HfrjEo1
RNWn1faTLjNq5QM4wXb6tazVizYKhaRHFM2ecdughR+fNwQd1Bp3cq83lts7U/rCqHVpbtgfMv94
8fmu6SIRW68dtaCB0EzVGxk8KY4AECxzbvuKrTUDbgePLsCqg4K8REsnIt8CQ198LdrxjLCeGu0a
bSDoazJKXX1LL3kHHoNHRSf3nNpiVzCz+uD6Ax2qS5eD8bzIPJdp17VprPqquVOnPMkuahvBp1ni
kcj9/b4CMp4nOvry+uHVttkgK86lz36yMOdCaq/jauUWq3K7WrocHDXTFr9hSdo6HlsOEcJt+yI7
3a6Tvs0/4U2FPmz2D0wlvLAxa8qeX9W57y3sgj6nf0cNI8/mCDKYV66LSoPlt/m9audPM1cQPGzt
s6XY4jQuiQLvhSd7S3v+ULIk6aFxi/Bx5HIhQFxsUBMYRe7YR0oROjG41a36B9KSp/OrpbecTPqj
nkrrIzbpvK7bC9o6vXoaIuLPFQ0k+adDBc3cxsnjtTr0RLB8GgA/SjHM7R7aJ7J2y+bFjfVPfGZX
fBnLeR5LmqGSNU0MsOyY70ossN9hvXZ1+5tPWttVgHlEWi/YfUkUAeDg+uICg9Nay+D+mto7tgzx
q7LxW4qO2kA0msF0pHtjEr6FlaFIt1Wn0gmqYojgh7RQrB948qYJ5jzAeb9wXfxc+QKg+Gzgs+vF
550RmpPGYfDRxATN15+oiEpQreCi9JDizCKJL37ThiQ6MIOmhNexzTiQaaYzcz4Q2GB0pchJC769
2JkFMls8eluZbs3LnpWm57HLM8WBzFhkpLy0ohyJgjEwQpxRpHG2Gyp5+cjBadRWDgqfkZ2VldRj
k1BBZMq9q20CQIF1ss5xrQq20amGQn8eWTL7NMIAD13zNMUN/pdjY/W/3UT/h4YTjn6uxkKBW3gd
P4eIBszuxvppzkatt/RmWwChxhSkgItiAIuHjO+qUPt7fqbfxvWpm6dcrl984C8m49fSHQNzrxHv
zrUDLbKUQp6Ypihjh0Wkq5RIgK2TxLRakSEmN4RjbhrselnSVHZdt/fXpYxp5ji57fwuhpKdSlMY
as2kDB8AnsPik5u1Tntrnj86fGgJ8IMPoNzyI1px9QAD/lQ/7UaxqmV8LsWD5cTecLxdwxZY8SW6
WsrV+xTqR7+gVGoszjl2ndPOsyq+ZoQ7gvMXfU5ByrUQoMY8gnO2ZcB3NMrulcFejjg0wmHNWE3J
gbUxdRRAA6FoOxlfZuv6Yz7AL+1bR05ZPwI7SLTOIjyvsHOSMWlU9JDi742BvpH7VqLNQVz0yuxh
zfxDJZEUClHVE0g3SkdkyF7gDEwnI8HwS6G5CX0tQu+dL8XdopZQ0AEQK2K8UoRbSeg3gHz2lYxC
BLmGpjv8vicOVsISmU2iuxZtVK7/1OBcNJlXTzpShTKrEF9/2w51JbICWD+ljF1lSn0XPCRherfn
KqiaAjzank+hnSXl/jY43fShq327eBn7fA0mfQGMBfcYxrwmnX4s0Dl4ZNAb1hqXNXsKL4tUcDpy
j2KCkGBJdX3T7QWV5J+YAJKYZW8QEh2LNRmFJAJi9AuRxH7I1ECs6lrlVPdl44bTxml8YhwabpPW
f90KGdFvrOXSbi3GeKsEV/JacyyE7+CCpk9mdF+XlbqSsy4Vv0Fgn2y6JMNTYQfyV+t3npaCSv8p
9P38BMpxJgU0HCar9hw9X7lFCCSS/RR7eXmRIuKvnz1DILdKvTtJSC5i2saM3Oql6wC37cEBeify
NRYNRQ4gRth9UefrRSBt8IM3vhJ62PqIpLBOSIhX6sfUD/EarlaIhRPiyNZO3qkX6m23J2fCHSP2
G2hOoUsvyywo/9iP3uMhnrHPaM3WDbvi/CnnayFYEX0qNVF/l3owiX4hAnBW70XYRusevAOWf2ul
fuSeyr04N5j8o6nphz6MEewB8+plgVLXxlkWDoRxiMLDchUDQgKme4obyjLY80xPOLs5WcUNKy5I
hx9Fp88Gue2zF9T0YbHgShgV9PGJEkNW2ewvWGRhe9sLvleEusRk89EbQJrJ1IJT3qOb+fOSl8C1
8RrLH/+CLcfX9t7YeOMpisykqQdv7LJdRWXQlRLrfhJ/KaPO96TU308FFGSVyiN6HkwqhHzUvZMA
sR+63PqY8NrKlSbwSNrwQWH18JFsUvvfja1TAhyzguN88HB8QRZK1KaxnIWRrJRh2dyXEskR3UIL
9wZz16lGRRe9FViwakMsqKcAJZb3TEdxUPKZhPlhs6CLwZhV+KCQHLokuUQiJCq3tQfUXYUvVwZq
30wAt1HnSzvz1xTfh0jT4t+zx5jc2pVNtYHgdah9k2eQmrSvdDZ8TkoDg5vuTf9IdamBrW72qgXr
8KmFu6In5tcedEs7pbxAE58dMcs9ynMeWl0eb8hozdOdYEGQF/J1pERPL7kRGA/H0JT4BhIYspFb
K/lhDzp5eu4f/jACzvHSC0kwFCytkKcjItteKEDhu/jHL39gzHi+EUzJ8xjCEoMmfvSZxn8yD7or
qrVrpQ946Ok7UwZUCXoDIwyqdDjs88essyMjgtT/fTBTEdg11IjNUUlFpHQkIJ4xhKYsNG2kpwc4
zKnYfwyIjwbhjz+FqEjLzrkAi1IoPi7bLs3UzBWeOHhGf2fYbDrjJdreN8yF0bIBmdQ/iVO4abKK
aqJjWSAJz9jxOJ/imTtpDsSjm84xZeJpxIBp/+HDRCBeFsniaHRh9FOqTsNg5aIIDeHW00dvRhUg
LRTrW1wQV9gPLzrvMhqV0q9/gi5ROGXoKsF9XlRFw//NvKB6WXy3nmYP6gxpSuydsP0geIwqb3gM
XuBZM5iBlZJlz8aJ6pNKc7Yodw+dTcCiwR/Edkt7lto2OM1aaX3LMxxvqZTYpmx33/vMRxGU1k9u
RWs13RL0nRRj7nWFc5FcGNnd3yTb0M6dQd9oewOE+kfuYYdT1+WIRouD27JkD9byVUQewex/0bcH
TP5gCLLZhGqrycmbB3P9t2r89968PxJVyWU2JLUCUGNRTFQ5Bkjplo9OdV8NU1HkR4hBWnZzSYrH
RE6bUcWxZ6JnpyyV19kAEy8cTIhS3JsNcEHP3lM/gPHPHcjDl4mCENWcOco6FxJph4VoJVfENHiO
/+I6UxPmkk62Ha6O3iKOUs9lfzW2blEDXWKQMErQzwBFHjoffr+JQIW8NonDzfC1uCDTeDow1BZ9
0l9ZtUrImrUYfihgsnweN/i2ADisUciPwYrbn0w3gnO+r6L6NJVLT4qAHbM6gkZyMEdQW4ewIkGH
k8JTMS3gnMeKt7yoRYjfLDU0XFC/sJlcjDPwhrefPXATeohDfkUVMhl7u3ChOvmC9VWXbRShdqiN
gUsuMCYX8x0ceBNR4cwt8TotUo9qyZdwYhavdLHDWM5E7GbrnZAcfXdz8aWwwOB5rpGOEZHZGeFz
SmkIfLbRWfdAHINtSguHAhWV6hZv48BmJLRq43wmaVzTIoLQ9T8p+Nt/pm5KvQj6XluNpK3V6zTG
qOL25nfrLzMI7A1pRAt5V8sNW2WGitcZfDjMQVTZP4JN0FO79TeYMVAKQ/OhybFQuZuSpTONNqD5
ni2ZEqR/tUOqNE10j2ZyBRKwXU7ItGrHFdeXjkcFvr8/KhHT54WisFEe0SIgF4t0BZVHBr7C/HpF
lWStHpyRUHL6QT4Ql8xJcvVp56fPFkZUaP2NoiP3QrzBI2bQpC2yXS9XN0Sy1oXBkir2gbGdXqJX
v5E2o7Sl6Dcl1QYpWPhyYmtOrZDCQWaWY0dn91oQJ/uBRPPtg/1iJfAxGWyt6SI6FW2F0HbbfE9H
3vmBQZwszDeqZ07PMlUv4B+oUoyfZTOo3MIomMr1QRJIP6/Ay97npmrLh+bAhEoO7DmYokL4t1OY
rdXwOgbER2SHEfP1Y/FpSn2upUFZfDuXvQlJxhp+ltSklz63j7j8oMveBRy8djX9N15Uo6Hgj5W5
ons77yBJOQIAc5MISi/A5Zq0MN5CBcyOoptqbG8rQS4umj5Y5nsJQcgpi9+wZaZa3Xk7IY83k47e
BFNJriA5faIJ5aemVw2nR7K+FkLnaUK39XHR3js/TqA/JvajUiTLPZQiW7gsT4YH11rqcpRBx+uI
GkbH1uNWqF8/aUBm738LFlmG3WbXhhCRuwVpLEBnSHGo0XDaqBrJsBCYvXktKLK6flULN1DPZgTb
0KqDKlgPcfsn8nix2xG55YP5f1TYHt2egKNACTJoYvBIcgo3lM0c3MMRkyeRKONc7e/i3s0XHZ31
0VQwdICelgtRCYb6GsKVpgTMRs8F+IiRhbRg2FjdOWGFQ4jgLCO0kS+ZH3ntY7B2+J+dhBSgFpa/
4NdBlsaH25V+vn9M35og7+197kAZozyDKZxqYDzoa1/RqkpSQVeKINV6T5NUICMapNBOnxLivvmZ
5uN5tVogXtP9lvg1kwsxrOffYzsay3yAVWRH+0v+cpzRlpsaaSDpCxtZ1j6LWfdj+AScQdzc6thB
WupdE/3uk9xuzlvg5wCbdziW2iysU1UI72KEBq8ji9MuaP9CmREayjVvGCy1/zG594bZ12lgwzda
QwmVaMtv9Z0kHZf5iZC/V0vp3pYSi4kX+0kdeqF39AI9zSFsDxW2aZAGVw/FiAuvcL3NQow99fl8
4l2mNEkOlg/2Iuoutdc+n05MpBwp3zSuz6Ib6oB5a1Pb27gOj8Zb6e86ynCj2UUFGDNfs0eIhGWD
wu8HSe4+4KTdZ+z4DzGf/xotxEGVujkIAFgleBthjaSy5XTfMFILBa8aoO93i85AuQ7P2Aystf7G
+xuNtUXOUH0pwrDQEBpMRUUAKiYBrcwJ8f86E7B4dhvXeK9q4iZYXInYftRRbmSaBWZ6KP1OFA1Q
tae82itzplHfQ0COpoTrGiCt04mQB71HviE1gZf7cJKv9uIeaaQFK/BXOHOFy0EQNz7b1wr+nmAf
4Y2/vyf2D8jbIEuy9wnxvzARqH0dJY5RQSNFgI3kScgxYc+OHHgrMdR310BYrTtzmHvby9i7avIm
DOLPHkfzUL96Jet3K0dQ/D+fvPZjl13ez6sPc+gjO8KFn3cxA4i2hmHN7Ujwg4PGJ1sS2aDAuTgD
TvWHNephxrhvz6Fz52iYApretA9pHE5fs0NQvcD2ca36bX5cxKKETlNyE2t+gd797atY7xpmWExt
5drMJKVTgmyl6fgRQp/pO3TneC4EdbrY+VdSgyX/R6pjCXzTUZlrDZX68S4Q7ZrVUlRONXMfOhmv
ZNJodFaa/AD/67u00AG9RvpM6uruaM1q4yjWfRp34gF6dPPUDcsVNXCiSYk/x0pMPYXb1OYUjj7A
1bkbyYFPejbGF8xxtTFLTzBw2LwTTbNxIF+IBPETthejuWVqhE7nTQigqVbpZsRWGzvTzxHhJQmg
Oz3mOh8Up71/O4sBspshp1C7pZS/kGoLu8WH4fRnzFQta7ixNkTp7zznbrd9one3FG1FqIUEcxRj
pmz/GmA2L04BuOk2T7SB2VSxak/DjoqOIOIMQ2sSbwOAf4zu7+cxgspjr2vozjNWNb/E9LTGf8nd
yA3JnPz8ncWG+FoPoGghBVHApIxsiKnQVd1ceQnwXsLggeFDtObKraptGqQSL6BNOM7Ke11Tixi1
JCmHFjsYte4F6VdYVB0EMJz4zJ85GtRwQLIag/eezevx1RChT8b19UrAwI26tRj6ryO5WLvIL2+t
r7RdX7eYndduZcpqa4ha4rqmFEO0F4fGnGTfFGLXunMztdmHaormyDGLFTo9p6aSlyL32TYREfJJ
E8yHzhTiyYrvvr5H4SN7XPF1YyPH0CacYW9w+Vyu+KmMeeKGyUqpnH+qQEejqW7VJdL/yOyB9rHs
QrsmFFvE/ejgx5N+ZcuncxwTVQcbTKUhOHNOJuTJ7UoWbXgN+9xKgN2naECHnndfyaA5IuezG3sU
2x0W+cK9UBQlKahG+AsX59mQFy/uuuodTA+jUWEGO6NvvPpaRMEFPu5ZB1HaKf5jUtrXbCBnac4p
KwEU+eJprufhwaMaOIyPVA2XzEr4w8MFTreLuQx2pB69z2PZ+73KC/bjTXRKwNE39eZxhzJZUaWX
eeih6UTZcebT7FjPj5p89Dg+UshDmfLsXiI4mHaQ3Y4PSy5KwUwFV+/f2oatbj6NzMvCR0uofe2p
ulVOpBp8FuX36lqTHquHIkxe4EeEhQAFir4+M7p5UkeWH9l8xKGCx7Ro6RSf5OK1q+OG/sufesXq
ye/u071MzhcEU3WrAxYI+RDiVpDs8HuexDk504zfmmmakaVxwrrTcmFw3kOJ6kvKJ9tWRziPQCmN
kLp1XbV46/TY6BGKaCIhLaVmgFIy3O7vHTTL2EmtYpd4lJf94fi/C5Xwff29dJk7rFH7Y26WS1MG
LIiuIwKARiM9V98sH18P5ihscmXq17PASeGdkT2KrsClfV238EiJC+GZHkL761e6nzlGyxFYD0cw
FUXTi856VqbR1EmAKabcMWE3RrkEB7iqQoQrsXUQ0fpdH/2lkpUi+SDP9mSgAssFTZfv3Ea/ZcZl
5dMg0fblGlXZqOQS25jXrKTtT1AS+4Yok+E8dINYKKkslH/gSgrgR2SlI62svLnKM8iihCG0L/7D
LNYH/oCY+NpDECyldzSDj5DF9zmD4ZGmWpW8Yth/wTcyG7kJM3dGqXSipghYj1iXVxIjgh0Hhpdi
rZjTawU5KmcBV9FlRXkc3AuJ/u68GCKRBnS0LXXlHQIML7FA5eQ32X6l6ENa80n+7ZUNGxQDEeyj
jBWOhTZT7p2/5weCr37t+nCdgazRagYTBvT4FwI1OTtYuvktB6BWEVdBDaa2OYzUxqaNrJgyOEq/
hwiyY2wuBeGLx5iWJZOqtpGVjCtlqam9lnotbopDGz7UjlQ6rB3gIBADK3i+ukpugGRxCV8V9sAt
VyCG8QU4XIktBLR+QIuJkV7DugH1hK2ty31qPPcV8luyAr0nxRvGC4vtrE7pS+gNEMOOo0200XvS
mw1EiA0WMCbnkD3Jq+Z3c4XdQJp/yYj/kXj5bcF17yBD/N8HBe0p5Jy2i2+7YzEUXcjLFuQAwhoh
FrEXY1SMoll/tJz1zaqfyNHx67eLuMnLjyP5xRqZSA70jdoNUavOnbFRWmVO7nL76TNn++NIHPgL
9GXk7W96suOUp+60lzEubw==
`protect end_protected

