

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hB1MkDF7gDUjtp9+r0pYANUYTDYvtQO1sWNXspOA3ppM8SYB929/qlOMzanhENZQcOQ3aiyEm3Wb
ozapXP+k8w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nob9JCRq6vcsk9H9VmyBE86hdNvS8BGq2p8Ka7dLN2J7EaHNc5IAaDkHipJixlCbGOjVeeUZyKme
HUzNgZTvjzVoRv6O00gQMvGJEhPJ3XxSJAOF+OM+ukp/m/tTtC3aiC1VdkFrdu6+fpapkZIb8cKo
kmCmWqIF3vlM9zcrSOg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qx+ritZx2pDvnekLOZeaFDvpDAtmg/hs096HU3U8xSeFyrj9v1CUwvI97hgO9fhp5hx7CLb4dRhp
iabDmveFs8T2afhIu9MmAO0ZqxUS0SV94sOYT5DwWoTjy8BTwRuP8Xrs/EEWKwKuWJp/Wjv7M9k+
wpkev7gSf92vj7uOWX6J6ECKwgIRjUGLc/NIrHrXqaq0yVd8j9fP6cvhVKR06OMq6U/6hMqO3Mwi
SQI1xdCXs2NXbTiCZKqVDbSBBvTJTo2cH6JXLB+E/g9NyF0e+z7oxCuyReCUVFJ21DVUfLxU3OhZ
gXG23tcqWGm/l3ZWHVqrETjEni8mwIO1yFoO4g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IXrSnaP8yioZkxR461AE2w19esRr4/fF4dA2RHFQL4fY5TpvMbkL+7RQBJ9eOLT5OFH1DsXcS+My
6KW+sTOsl2ndsfe3ttRCDI7Oeo8joeNZ8xJuwUGdOxtV0ae9PUAaVjkgDttLOomzNLph4uCXW202
bI3eFzZlGpn1iGIKiFQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iqW10+NxHcU1vbwMjaJKEOrgcrSi68eS0/IgZB3xPrIkkojO6+T2kz9ISwjr3CN6PcPo+hXCdZn3
Q3TnU/fMPFYF96Bkmhtr7AtYZE8GinVZHXJyKmm5x7dcsR8FyNv3nSOE/XYU/dyZhfnBj9H8LA1H
EJZm8T3/SQk6AB6tpXwh7kVAfE+bMsPCp98Fijzd/ynv1FX6O6GWv4CZpIVUKm7Fr8lIGCex7lCq
foNktfSIPTqF27RC3UxvVuy2VPf0Ck+rGl7pVu7l375TxqfmSlC5QxbXyTQ1NByeHr2LVJZwC+Xp
5uMCktl5vyr3uh4gEJyZSJlJ7E+uSrhstePVYg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37424)
`protect data_block
9dz6tYy7bVT5uVdoXw62hw788opPvi8IMhu68AEJ76AhxNkN7oWluO4RTfkwUL9R2kentxfpQflF
On4Bv1FrJWbiR3ZWpACmaZzwn+5YMVcZWRDdadBk38z4mK5XY1i06yoHsIavTFFEgIhqKZKyG5xq
vrX+htaBDSktA3xZ+aPzl0kkP8S3R3iAOHSv/pPAlGkfFmluzXEIlXu7mcnect3I2nJcSgfTOqVD
OT511ug/AFSVHAzx6yNIsGjVocVUmTC7da4mOvc1Q91YyWXNbXhh+vpg4De6Dr5esMp2Rk93z9zQ
3YSgc1f7G3fVXpLcEmWsgxXOOd+h+IpEcoQCn7Xw2gx6llBhLVuiZUxt6r4zt/MdlaGGycO3UHwf
NuiVmEvc42ARgvjnRcLKmSc4i+h8iS51Zf+jXXCBoNIjNwZdej1IvK0CmQ9x8I6eWtpXNYKix76S
iAAzgm3D/64J8u56BkrVSkzrm4cE+ss3XI8CyQkOJVHHnYQVsWI65u4N5LqwZ76pOW9rpvftD9Ut
+Ob/KBdESWcq7yTtRtWVsnu/KwAMTI6mJQv79o1JynYjpVotiOa+Gtkuvu1AIn92Rl128ci9jnQj
0WtEjs62a3GCMqrgqjLA9amaJXSqUZEGY1ByVy8BM95lhDt5E1sEihgbSDwpAbunIT4yHQdpe58I
vHZNDZvrCMo5BLHYegS8t6+hE0LfECIapzI9KHViv31wWdpg3oibvMR856PSOxe05EAp7bYFtePS
Q+uxzvxh6uuybmwD1ZGJfknHhBpOuJuAbI7GpGbOIBr+29/RrseBkEqgqYB8mBejuZu617ziVOuO
Bp80AA0WBI+RuBCWk4EC+6cOEYn1VL956oN9pnxHrdeI0/7U6uQurKXrY98Wjmo6EUCQ1HpOmoHp
ihc+EF1rWmSnYYdl61TasawGa5GUySTQmek1xiL6bdNV+H2D5cao4IqMfbUfrrVgNOc5oskhgm57
XTExoZMdf8kqzsBA6ih3ptolEi11nH4p+dheIyFjRTEKBYZIdv9wQNZztQGzgu41rru3IUkYkg1y
0DzDdMVTlw/4k2Zft76Qsx6GRwEw8HAsxQmBg/GBV80/Sk1CP6Y1Le8fuTciVUBvCvBtJXg4alTq
KC5fB1k5kVErtxNlWHlTwWP4FKzgujfjBWSlfEwrNZXJIi40kWD8KXQ2cPCBQQSrKAKTMafpMAmv
5TOwQwh/0SQNmvMFVDBiTp//E0nJMnKb6MkEFavvSAijNmW1m8eGOA3JIQcp56YZz3LaVTo6lMRP
DCXQbUGpHAfX01CYoPaKbRwtAYtC9H5Mp4ZPBclHZd3zOjdXNCjUeeBS03l6A8AFerLaK5eQCNe3
qdJTi62Pz0t7+wLH0HM4QRCPbTF9Cs2HhykZjy8pDaVCOWDcLrbOv2XquoZPZaLu5zyFU1OYAzGu
bNPEU2Oj7jQtwIuS5qT9L09owGq4SUt5qamR4Lb16DKqw9cR/olz3wVEUIxRk9JbSGpi3dgn6H1E
3osVX6Xqik9LMNe42emKKF2yL9KCmoEV/ko8oTdQUBNALSUXsBDD/SKZx090lWtj2msMuL+uXhjG
a29sMIqpS2YPDN1izNhlcBtBkQpRXan/7SX0G/tqa5Wj2HrsBuWS0WbGtvNQW2gyZz0CDNis9XBt
QIT8hsgjXsFoj8cpYpV/ZJeCYRY+MYSysOf682/wbgcK2bEd0hqLBm0IUiJ122OT9f5pnlfoeDGM
rp2wxDPAGneeSHpe3Sg8dskLmyxkSSeum0sSvVQbD04YFht+hIhF5cimKXiii1GOoyxXa6uc9+3C
rLrQMEWmKLoCCSp2ZyEasb5lTCEV+ZBGNasKqEmqnwDBwZs96U5WgOpy0itM5pMPr2x0+Lu24qK/
3Q+ofLFx1NSVLb7SqT0hJ9TkqHKejdbHyf4KStitWFcPa+5YaCt6QRdiuC8yEXKoWlBdmoy0yp/r
KAOMFgREDvD1KKCYJDTGhWA2Z22gprertQ/0X1W8YIEVmFIK2JUFfQKNlYpuT2sK9i9OD50rppdD
gVQYMG7XG0wu2Y52JX1cI64wFRK5cGawo+7AgrHPwaml4nDOw+X3Zmmw1PEtZV1QZ6mZKoWe+qNf
ccgKmbVHOhFlzNP/rWiep8ZhIbwK1vPDd8GgsQ3iub0wFVGu8YsGTkJMOwxIS5SLoziNhyvhDpRc
0vtU1vUKTMd5oX27a96Kq5WZhLfkFHdivCqN3FRRrGJEcDMoBojp6fwEiEvLikOqeXzB1eB7DM06
b09hKmOEvpUlU8zFatPeYmNVGDsRPR1yZDwWGhCNndpuQLNgGcwN6toIKavxW95l2UTuKy4mPNWq
ra3u9Gq7QhrSsQqxRqD3kLuKTpB5Pg/hgx04AfIkDl+8JcTxAxKvsFvHNuSU4CHFVBVFCMIwIHdH
1bpie4j8pYa4ABlDRs9Ar56lYr82IZGHVNcwO8hm87+cxVlizMeptqr8Zu3BRp02TNU801ebEEJX
5FunJEsWpoxjy6Oy5p0TL/CEuFhMFZyZqurigIieZ/2ek8tWRH4IpOdo9q4bR9a+IYdWV0c4oNee
mC6r+DnPBqzSI2M6Y7TpKIqe92P2WwtwqVMqNMCVMazvzpf512IA0D10waTyzo1+1TaolrQMwnCn
Dc/xoQu+/dfcKUopJkkJ0t2sbfQVSpxVPer2nMIrDjWYBW9cAW6hOKa7PX51EDOTdFQyt5+1QVHW
qvkEVfrqxoCQU+0NbC0taf74EIFqll784dqgdRP1y8OX1tj3t2ktXXbcFYzgpGWMh1DUl91AEXCD
/EEPpFeya3ilmvkggng71bFc1CappBqm5j9M9U0jAFx/tA2SODHLKv3K4sQeM+hCLPsYCtQfe1vo
SzFXhmRKcIXDKttz7zcyD9Am9NSH8+Hd7nQInglz8bosc2oCZfoMLYj88N4XsHDtk88XVRE3yF+f
GvuxkKNDFCQswFdJp6h75B9AUrWtqqcoCFr+TOJoayECK7IucfhyqnnlZMRXfW0pAx9sqihygVdS
RNdQiJhF245C0qdZYFqo48+JHWCJQkc965zkVCrloHCasBGUqBFc7ZHFVy9iIciiiVnDJZE+UKWF
Bj+ozGABejDbQsj+9EvRAYVclD7pUOK5aQGT9mK5fg6OV8EFndl5HMKxNn4yHWzLr39z53p5Ye/v
FRWRkupS5qXX68BILGqxvI8CEMPz1u3Z31KB9ly9eNzQcFVFx9KUHtMDpA+E7ryycKUvg+4nNhex
nMotMTxlnkkefu+xlTxArb7kLtdyXae7/1HEB/qdFU40v9lw3t5PO1RNG3HYszGSZcTOMV1gdRBn
haSgzDqccJugezOaMJRGYd4wSMh7SGcmMXwrUH1BcMCD1SyJnAarJb7KBjbMTWeQcYW+FJR7S30d
ejXflod6t7CuJgmzOilWyT6J7tKb8w5+fsTkc7HbiWlCi0VHGB7rqD7ZuTD4fIqiQsEWHrjMK5XT
xTcZtHKBmOs5FR4bTgHnSy5OO3lgszVXMRFQgwfXbu1e2TGW/6ErTVK3b4aFa+iDbrifnF6W/CCT
17pS81IXK+f3nLnCIN5fVm4FKVeervvFb5Sq2rsteobOb3g/0IWcW82iK+0zLIB8pH1nyhMY4Hyk
gSvJOT/gFxJ0loCWz3UsHHiGiQVne5zldgC7c6VZrADhytRAjTzfRV2oOdxEc/n0SgshONcbogZ2
tyTD+Mva9S2V786nOIct2JMXDa9jkh02U3Ho6IfBPOQsK+JFCswcO1XSCo2S4BodtdlloZkZgGQW
JLeheLQDODmhrXZxifkeFcM6VBMKqxXnh7GiPsFUz1ErkvaRdHS062UV5tUchtvpvvU9aLmihBXN
oHG/bospuZEjp0aAn01v5zaLNjAtm667zUro21oPn2b8DDF6Qmkm4iJu7L2HlIiT8kc+9YSFDWgv
MJ95nil+DGn7m+RR7x2JHzsCeWwscqwFHhC7/JnXuLW0OSUg/JB7M6A44jgwuJBIhT/hboUuIMuN
Yyl1JPCKTBAyMle7lccZ3rc/hOJpTewh/hSQHFGjpTq9QjAwRCaZE9/vTAQXb9QdzaNkql143GEf
HwvNEf3F3aR2O1S38gfrdhyYXEyw3QDl8acq3Bscg+fcH1+W1oSoarsgSTM3EovJJ0qCMRgNFeHV
WtV5Mu4Quk/8980usZx7LQLNF5XvgSOO3SOO7JxBS3FJqyRIbAcJDt9ySJBZ6o00OdSxpxVwmMII
wYvgp+qzNVNNlE8yKGSIQR4jWuXtf9M5xDrWGMGTPWQAfcph0hXDw365oi3FJSPqcp9eH/S8/GLn
r+tMTPTEJkDLzw0hzJ30TBWM7uEFwWe5EYeDLZ9P/vsbO4c7imckmbaMihFhb15usmII1Z07iW/N
4HhLiSsTxCT8+wgsN0q2wu6bX0DzXAHK0dp9lJTTmkKBX5RA1VJXUpAPDbpfsLxQaF8MIVPQfRVX
pjGnNCF8whobvCCTPeY8lSgumM8ZXLuGm3IySeIw8v4hqbq9wCdNX6ZPk/N3gaAl1IyR9k2rsDMo
3xg9/xOmpDIxrkW9U6DEH0fJgPr44Lw2SIXgd4iQHkQd0VZlF5rpEZ5xdNXnbRkpRftA6YX9BmDV
j+wHZFyFC0tGJyCT2r0iYkGB/XZK/66GZtNpkyNvgyQBVZmniV0zE3VWilFIqtFuiyaLNJTZGDc7
+uvro750z5TDsygfpMm2se1ggnmPBqxwVkeVGyAAAOMFabmXO4+0+tmFkFyZ/Qr36mHKVHXWKKyH
iFjx9OvRbmEuJygQPak4xM2VFalGu3XQtpDmTz2pOK2kE/ssAKbZvJRXn8wUbxEf9XATkrZ/aQgB
bJy/qpR4rtgF2z8cx+mbcOTliBZJX9KhnpUYlrg0vFK3E+YVd5Hc/nnUSDNMga9su4D+KBD9Zz30
hu+r82arEDkGDMoOgT70J7oHDeoyWeWzudRl3eaA4O2cMeCNow7DKJ666n9x/wHaxjGRYhx4lhaW
hm2ocxsYJOI3KxuEs4dYbPEeEjq1lVHn3tbMm952zC/Q3MmQtjlkxhxph7DVt21KnBzq7CzIsHzC
FuH5hXrMyYuZw/NPBZa1sNNkxXtV2P5KpW+x4f9ZlLLa9WBFj9g1IKQY8ZcMSITaSknM+JBn+cqs
0IMAcfFBan+Xix65+kMoAt20uTgwUP+QlyryzzbxOf/izrK0tR3N7WB1ABVIYwdxaL9SxJ0U5R8D
9Uer50Il+bzRYTb7ZVnZTCnQFk4jarKGu+n7akdXzDWVZ8wwAYqyYamMWZKxMYfrEYM4YI30GYIr
Iu4vXf360XHO9Dc2GIKjJ94EkhSw8waUU5izjF9Tqb65ztRmilWUHy2Xbt/6kgEBo27+qAy1hP7x
k44p7tgBSmtelDt1DDRQrUUGgay9ZbPnzE41N1LxqorEUh65WmZ9+AyIBevBpfnHtzWr7n3i5/6m
AFjFUKejDytAZRdyt+4wEgvTTP4H0CU2gRwQGyinx/E3gHYDITpfFrX9RU1gYy3O2lGLrL00Bozr
6fLEL/xatAxYrGzyHLLhW99r49/662Gwuf63k0F/eBd2P4wkoOvu8LMSNyoM03Y1Ndr10h8SuRLv
Hb08/VgfALGLqYnvrvM6FSEvNvi3oH9mDoZALrweP4ias7euO0VSvADdt7ZhdeoTZCQe7uPcoyoW
Ekg1Olbt4rx5muX6OhxMrIytdvHvGFQQ3tqwE4QXmY1M6icYc3Eo4ivwD44aijSMnMQhTFJIEKsk
tBZ4S7C3p1UnXVr+QhN7q9BGEYLzlwjcQfGw2mQmRWcYoy8pMQ7ykUjLKHdCBNq1i21quZlDxjR1
egCG6/5LziGF1HEn8OOF8Pgwi2PA0vnzPlZfZm60L6uyl3QrV0YT+l5EUuWRbowT89BVPrXwLKQV
JBJLo8VuigpaCZMXWbkTqZP8j2GR2Q02+hsWrYXILoE/h5krVbcbiAzWedZgOROkLN5DhheKF/OF
6y8Jqm8FXIrJiWUNHTJuccjQwXuNCntwMyIjWesJzmJ3dQG3VkG2MhfI6idzXdNd1adqKd/nbvPO
NKSyfnfsEH7YAaMFCDgnLUL6ZNlyFqrll7EmirRBZql8cyebwA+D5Vh0gff5msRRBiZRhU0NoE1T
AIwPEuuyQuxJPsrDEaNlCi+jD8meKJshcUpsnQ5PCHuA0OPL/8kcmGCLvZsgyjFwSGI5aEDO3AKG
RTKpDlQf4nboT3vPxvzXlMQfuKfiqGPAAZskQ32AqDwzYook53VCWsMako24qfWt81BUY8aZ3FDm
+rZxrNBXT5gHMmmz2iKeaWUR71Ok5ygFKgyc59AvNskPFpU0P8XdQ2YAp2WPXMuAWlAQ2sywiSNd
hvmYHOcj6FpNX4mkcu4d8LkA7deeGkV9/0AG733mtHpiASneiGwFmybw+R6ZYUnr7GNQIkcvFxkE
pZsKyrWHaStYgy20NIhJayUx++4Vz8owPAkpN3+ALf1SREgRoKDXYhsv1fwQovSCFgsE2I3m+zUi
uphjMTQ1mQMwndHbbW3PiGAHVDJLHp0UKVhzm/UJwVYJdVrCsA7FE6ViA1CXK2ZGifs0h8xJCWeh
d6BfD7xqFYYNBifcy8gXM73QIznklFSn5cf0T77KJKPCkneZszJWT9/Cfx63Mci82iKOrZUJ+YLM
0YaFRuSVAV0ISq17IXSYuHih2qjbLc5b6ZuktFxD/XsOSCovb93PxnC65EVtfCK+dgX6p0IB03dL
cEJL/s7oNfsSZ9XAuO10xL4P+kdC9yX+n5hA+q1NFGhLD8LETysu8FiLX+Kztk6/dMJGY0On9dEc
t6ymK9ewycdT8uL33HpXRA69YIFS25vEs4+2zTVpDYOLeijzhWz2kGBblinM15KM3ljgiledhjip
FlG0coLk5CPxWgKhCg/IxIL0pFxkYg1LBvPDkdE4vvf7kkj82ZCD8LKoD7Z0OtI7hxGb81QDYLqJ
JK/MzzOP6wRH0qcANiF6oMvdme/KdLiWOkuBa3pgP4hWayGwEYYB9SpgvUwJ2kn70Q2hm/pRLNW3
zNZshOokfUT5lTwXAOpnh0AUMWpDST5BOdGSA0QrbDeKafmBX7Fh0TlaeTJvEJkfDAZOVeLSajlU
Q0egjcradvgiIrxz/Yqyhjde3FpOtl7Jred4BQawpaseGya7ZVkex+R724iR4oHdwInawdMXp1qm
NZ/2T8aG+MB1s5SFblTbscJ4WGoJbJ5CXXnIaw+tZPyCI180fp9SQfRjIsGe0aZpmIj1Owei1pEp
N5G/F9J9pWP5ueq00NWbFhyN1Jj9jgiG1y7rZH6c7ALLHEMb6g7k8RnAgVoH7gOFujOH2v/taAZy
LqVi1Vs5XUUi76jegO5D37JAxVYOb/FD/rWqG4FEtpAkd/KgbQTy4nGtJ4E+q8/EfzLUCQEH+tl5
wRGkANGl9yljyxi8ZjZ3S3XWgx/qPkLK4gewddu2qZeUeveD67kd+NL5MHqhxPsNeYI/uuFWOf0q
6+v4H1fMBLI8p5xMDWXB0OOCH4sAN6eYfP3INGo+qvAneMSxDXNOy22RiGt3jdcOPxgN1ZoGj9xz
SlwZ5uWt+bwaD5AJimR9ek2nwkpPQi13aRMzcqsjT/qGvy53wExA7Wr7mxZHbe4geF1lkeUtPVkS
IgTUFmKXjlrUSqEXPdZsgpSnOAzKo5NZXz1SIXG7RdZR4C39KtLUGJky+qUjU4c+z/pLAyqajANY
8TuSNC2KWaIiYdSvKo7Cc3bUO9QRx5LuYX5jsv341Bh2cQ9iEDgpkeNz56eUFXIRv7+TgFf98nZs
gDkH6en2FWAzdP820rP13K4tS9KyA0k0xxY3yN0WNFZBoOe/TuI/nOjJkoDbsyBcUbIErJimPo2z
CVZjWVtndctAEAre9ByMV09beoLXnaeOKUqls05OeiXk4phlsg+lkEpF/6V3ZcQ7xDmzJUA9m7Ee
fltysHyItRn+IPI4rzVy781yKlX9FUEC2R8xTxiGj9LerWWnv56qKh0HMCm0sgJeAphzr20Jyxq3
PNgcfEvg/vTq6LJzd/Eu3FP301Qgs8MEHxiqeJNcKGDnY0xQp7AZpZKZEg3Bxz4V1ENfRMMqo9Bd
EmKIUBsg89Kw3atRffmInaEvhRb2yr9qY80+rIAIqTJg2bxQWxnvWOxFdnUiV+fzOjxr9T1XqQ2B
419OwC9z2FApeGzuWUcrMiSYy9Xt9xQ51fcKkfTQ0UPy2YOYhhN4zM+qx0z/LI2PEG1YpmzDgASC
MnFfpGVPwYUUJJhAigfjUNy89W2TlDynA0dW1KvooCgKISyrttBJoM5zRXTyZMJHEngg9B1FPrg6
3lEgIgyNLOT3wGkRfJh457jacdME2Q4DiEw417maFx2XHCBLiUgSaofNVnU+0oabGi1keyLv3nXj
rni0b1iovKBNGqnIIMhx/Y8mLj9uVTzhHqgKq0fPFTEpBhlASPspGejncp3XUug7jmiNg2YDQY6I
s1r0GHPcE7FI16fK1Cb0xjfL+8N7HlUFrGjRctWvAVj61YD9ALyoXuarKxuCVLr2QtZhjrPqMQOd
8YrGg68eU21MnSPUbyFe04tQR9hBquIG+Xsq7VCrFx328w2C+Qu0br81BlTKqU1duJT0aVbFP1ES
yGt80tRJvGhhqWSxU2qMaxKtDv026o5bGPlaWZGv8apC/2ttNdEkaC2hHSA2fqC4nwKR+XElkKOH
J/Az9wZT/yUF6L8onB7t9acm1a0/MjYgae7JnPfok5COqNWiBoUszQE5XwjtQoqqd0l5BW376iRy
GT28g9qlYoTh2Awx4T4bg6fNzLXYzwJ8k3D1080N54aQZONvhpU6uzC3WTi7nIMbudarRqRucLv/
UpIEh+ZrBioVCg2/F/EUOsexCdzBL1satmO3MksstXCipDbYUkArJrJeaUy7efhbPAMYQyBMRYHv
dKPFgJZPchcNfCr/nvxQpkg1bM63GfjQpUUb+GsqrD17BJrqeujk3gHm4ryR2wRwoAP0RH8EKD7F
mgFt+ztjt6tQ5CvK36DCgvwUXtKG62ZR1g2Qolh+Y9Zjgi3gx4bn+y7WGLUSJjZpto6eHzDHnGjB
TZyPNrBSIxXCbdO1Z0e6LhO1qV5QsAaLxNLz9TnooUtgf3WGwCkKx2E+s89K3MLAwdkURQc3hbUi
1/H3m6d1mHeFJNl3Vf+om47C1E9w6Vk38+mJ2mRSywutN5L1G+z1nWWsRJvApvnnRtfEW9MAnUvE
bZf9FoWFwrBO4FXhSIrIJ9XZ6EgNAF8lfzdDfVKLaKRXLG8g4zP9B2XqAgGm5LkibWqB0B4MLWvT
DtTVJlfjZIzhEUo9EqFjPrrPj/3S8ePdFhxMO674PasKH4VS5UG2ugmewpuCZOAo561yaDqkKAgO
eN0musvuwutIi/lAvR8uEwZ4E3KaeFJA3mVP8lt1Pjy8OPoRKtmgXlIVcbOUq573pcdrs8AIjSy8
IatsrXyZkdhSgapii1zPsljsgJbyFTXgsph9utumsCwEqKx8haY9sx8FYef61PIvSI14M5g0WzUK
hhXCFYVzluGNHkjJ+epza29bbiK6NBoEbfMEC2tSMZ3fOYLh0Ebx3jeLjQ1So+GdgyxOD66NdFwr
+aXqbW/JvbzukhTw83u/lhsWVSFnMQgWz8ngi/avSmA74MnM5JIB3TIkEYCsF1ZstHCRRAH4Z+Xk
J8OJZv5nBp3wVP1QIbTbYFw1ZTcHYx+gANtgGJTscPORP6wnaohSBLEyqDT38/YURFaVT7S71xCR
vcw1SIaEoLbE9wbBBMamM2rZBdQ+Md7OaItoSClKSwGuYrbJA8rrj1H54vZVv2+aQVNaq1Dn4Lmi
MMlSKxlRBYfrLLo+itvHMXnuajDrpyDFEVaJ1f5ZkmlcRw2TGf85Kw7hdKoDtPBgbZLqOcBoE/pb
TaAtDHMJBR3OeBpYI4xeDtoVpV2CHCkrb2+fBIcjmPcTu/rTKEaACa09p+6fxzSO0eN6wC9jJLe3
vfpZd83TB2Al/2z7BWHWCT/15c9vtChhS6FDS4Lmat9fn4LZPfcth+gvmHA7fQAzGxpF4+aKZlzq
HUNxvYyd846/IQB5VJ+kL6ENMGCkeENmyyUIM4n7Eg9FUsQrH5/MK4725ek0IoOPqmB/WfN4H+pc
vPjjSltYpsAqJcDELP61kLZ6sB8jVwFxfyppB6bNP6pvopnXYDp6lmkkpslo9CcqVzkdIAny+NLI
z8RVRAzdIb1kIdaKspQ8eQvL9QNOP1+JW0WIU2xxqASIYTreGrp8i2XUNqvUa2YByBZyp1qLdz0V
DJ5Wms52TjTe5FUyEuL/WaePyBSOE0jo1tQD5YD49AaYRZN1AFEqGN0538UJcC3F01lxhYOJoFiC
Rjg0YOI8ridd6StY0YS+E67a7+A4KmbNkumwdY4KL2TcRmcJ6HGFLCFqIAc+GymQ1KVVAgDQ+L2F
gNQRlQJ13/uRs35KmJtcZSKz8K+GGWrLBHRWXGyZpcjHEb7tOxHFg+mRuXAko9VBBitouyl8+atG
zgNroAVMBh8+HaHbGPuql8NBCMfhcgHoXkO/EWp1+xRUV4i3vvD+dN+HoJdKsrv1bs7Ld+MdaD0O
cFcF9Bxsrc9i5FErz0c5drn5UqV4OYrRrOWkiAP9KL9M8PoGiorjqA+BExHdBqQMLV+AmZ58CcZb
mv1MtyIhlGRbBLjeg9QYuu7myj5nT3ZG/3FhSsDyPgobaxaUNH/Cv+swQzVdoeX4ka7kGgcbPoW5
vZD+gIqgq4B2LfQTv/HNmmdR+31celxFxZUIVFJFMlKLXCEvDOKtA3mPtVDKfcI1Tj8VsefMPJoe
79SesuRvlUskJvkCwoJ9dMFLJxV8G2WmuVxNRJaVwPQXbBK3uVsX408xlYamxRtxvUqZTTm21Z2N
2ZyGNGkt9t+kJd/LJejwSrBTUuTX37wqtZetM+9PvnR1e/PhzByALfLxeitcnzVA9ruD3sMHlq9h
V8OVLHEWtWok/VUwa8n5IIzmTBb4DYEJ/2zeGA/he/eBEzs5dM6Jhvl5DJsMULIm4NzNzVpnV8TZ
2WCVncJQ7ZkaRQFCDIDGeTZcyc8W+CBzyCTvn+fVfiv6RMwxQeN+ZJ1HTXXjybInYFwfuZu6WsSu
N4q5pMcY8Wo3OATZpc+S02ZbGx6skJKiINNpUvy4CumsQ3R8BO0Koxqxs8iuK1Pjnu9OyPyjhH46
4rpyE7CIIJNniN75qudZBLRor4CtTo1RkAWSEO9xSg8BQjE36fml6jB9vR3jaBPskva4N65NDTf5
qNgWXs1KxYHaKq8O6i6RMAjkCpR2XefdCS/aRe3jJbS1rAnswedmqUMYDIVocGfjnS+lCGB88og9
2hT1KXHQunSs/NClWFZAZdiO9Lo/0x2FGHuS3mVM5hte28PN8nbu7TG82ivvb20Y4MUek7k7roZA
+YtvMJYuSqrXm2//Cm6MfaWOO+Jz99MKwnPQlxcURKCwKRR4gAg1pA+NMj1pdejlhvlcrVUvyrz1
CA0iXZuo4bbBKElUJrGiX3xKQz0aHSuLgnvOEEK+ci+gvFP1dt2gDoum5q4K3NeQaTNEpRNJQXXi
EgvPen9YFloREXwtkjiYoWSaVzysBHipDoXUvDgZKd4wtE2QcTjagKzQfGuSNAcobeun6cjAKwoX
cb6oG4itu6jP0EIITxbjZkQhnjLvkq+hqzg12RvogJDVTJ1pYIPtuzczGWJESAMvgjwRpqDeiKWs
OE96wmyxTFHn10tT/i7yUAfw9e7Et1tjc8+K6fav5TJvB7D/JKEV3251rz1sBGysEZtU31TDxCuj
JSaF8XXJe5KwiYzn4v4k44sYKMlJUwx4sdKUdS3Zt1bt2v3umRpCsGw3NgyiPZ2Fp6SHG7NKvXL0
E5fTDsrR2rhIciiwEFTgrJAtrFKvfkO/SQOb3MfxVKlbqOF8nisJKxNcoYd32esqiJpgTy4I8mbo
yG0M1wSPfML3yt4soDxZ+fkW8W07GoAcQK3AXiLdtGDEgILRlcMPu9iJ/egNVdt6pBUStujCS+jx
3e38GcbR5TnHBrRs2jLctm4Vh37xRv3kfTlIskzlpZg38RSe4wZjRv74cqSDuUFqNHzARbN/5gKZ
0z32SBnLu1rbUtkXc+Al6UhMG0SMFoniH1zfT5F53p9H7Qxfn/JN8a7hF+co2+VSWlrCCXfuSs/w
ExVUAAU1KJ0kbMMJiVrrMUF5bxZSxnUjBsYm8g+C483ykdDpDWLWPZxEFwMLOdaa/HLs/4YVADlo
Jt/TO3dw7UKtExvUmnY7ZHzDCFc3NZXgSZbOUL57hncPAoYEE/E0IDvh5LhmYX82TVa/JMKURDeV
Vkw1X0lx97SwrUCL5RyR5/d1ywYXH8auUA+HnNqoGQMVVFLDE5YiSyJvIhzbKG3sEafUyfhuu91B
7Asf99hhRXJ0UvNWpZ+xxv5pnWUxo6y9mlpQUI65TiP1rlcPcwTR0PacAvnBn0Cngnk1sWqnPNKK
a3tTphNVSTBINUAe/PwO6QtOC8il4IKw3DijSk4Ec7sIoNIsZq8uwB+1UcL4TXwuj8y95BAg0Ycc
mQRPnUKaAbrD0cTlo2JmdLp+cfEe5/kIx8Fr5XssgSWvxwpcpIi7I+1pYNg/A8w27E8TOqSuy99U
Qw0EIekxGLV2K9yRE8Xf99krSDioYgNtQHFhWoEHWZR/h8Eeq2kq539Z9nCaJrKeuxFfwCRw9XVB
gbHkOY5GymfZDwn8D5k8pi37t0QuBe8cllP85RRJbSSMOOJxmqsJ5UsC8LX6o9wsFdX63HB0JEw0
0r/zv3N5pcIEHBYuYtUSD2XiYAfkfqmjfJhMS70DR/aMpSwbEhgI2vu4xI6S/oyNM+URw3mj8f7G
dlp4e7EomuKsxij7/n4ixpCri2ajtfm3DHibiUxVBIfmdIRb2q+B4EQAGg5stD+hmSgLoySPcXhh
l87YjBreNc1B3iSTrGFbKr4I47W6tWkt9EnTZsq70jyko/WTFNCQyVXvScm28lcCQNvbEBXhy5HP
pVDrd9toGBoS37VXsrPSWFp2MV4+39L6ca/lTf1Qqbbvj+W0KdR/NzG2lrOJ+AtlxuW4CdJATQ5a
Ah/9Fq8pE3eCck7m5xUvr7UZHQLq9OEUqyLcfcf0k8Sj5M5Nue7uJ6/6FMLEKBkG171QssSnRLU2
rf282lDeq4g7ofYpi+qtmsDzsOjVs7Om/WEESds1gFYDM1afpn63J+zXgGgRMgqNgJy/gX8TsMSh
6sS1r+9OlhcYlo0rpp8jQbnk/5rh8jrcyQN2EYOILrFKMBB91JnF98HoVSFk17LOXqnsAy/SM4hh
FkhKGbnniHLj7/4sDXLGHQGghlYPK4cNrFshc6UVui+FFVJzFZ1iE/KDVyiK8TGOowYJius8OjXj
Zb6Wzp5+8doQ5YA0E3B33ScuJbZPq5XoUMMM4xbrNpVXp4YTVVrEpJaJtg6w3hmgoxqpu+7ek8xz
1T7zCNgd/gAOpljm+bdIXPWDc68Mpkbt+0Fb2J/MMy0atHJk2xLamM5kBt56VfIIbqeQ0H4YFN4i
OQyu4jT+CtHI/d/qT11/jDoql5p0dnnXKCTDuYlDLWs2WEaM/Y/ZuLwuhfZlK4fr4x8MaAxONp0Q
CEGJdAnLkUoQ7/HUsb7mtD6Ykpzbiiyihep2x2KHyRAsmX7Tgs0oxlXkQzbHv0h4FbVDmXAFYUBl
zDKRB4nZciLJVlNTW26GDfFL8hbYNI2FeXjShP5ENmbZTdT1BbiC3xh9RiT1Fc8+QsjiXV4eSzzG
xDIy4Fhr64Elljo9oOEEzf0qrvb2LWVGhcLnzBD6GsUO0HBWhrAvm5o5Wimy9SN7eEdnT9VM3bqp
UC0EVx4sER/EYBRTS01wOnr11/OWoY3EAgre2I0eEBZiOLHnr3B2mL6TASUYe0bLSutNzQDoMCuG
CSFw6syjzanmCB+D5DyBWOVOXgfPbXezz+B94602W5vKONU8gzmbKsD7OwEZSbyZswOZEz6csHUT
E9YLJqwu0Z018n43t8XlRv0YJlXAXB34pYUYhQQnMbfHZOX9kDlNOxamQjlwB+nIIQh/DmQy7GAv
kEwmrLwaOzmOX+7YsuKVb5jK3gL4Jzsy58G2ST+sz/bBPesXqDGJp9DRc7EbNnAYcD0h8NYNjVHL
N96bap53ZuHLTWhoIn1xFbl9ntv6iZL4QK3Qp9v3dOBOAGwxRSt3ewl8L9YH2tOtmLoK4qMMOPeL
ePxbHeIkb52NkvUxx+XbAzsXhmT/9KS2mJcL72TFX/WyAfgzf3s6fe/PU3MrFZ1Y6DvU+BHSwvB1
Fd0fhyE0Ei4cfYrI84xoFZ8bjBt90zuFX6GfiF1C0iUGc0tCcF251Z4uiWPD2vnOHEbupgeWqxSm
ihJTlInhwqSBc4IWksPinrd9jL7mTNAuOwqq1Z6TZWpKTNgrGwWTFi3+CSyWQt1CV8JbCbeK5Bd+
gCKG6Wv0ctaJqFmN4bTQmMXwRTUn6/igRk8qPVxEDAdE8n1WIzeOMJedDdwdg/21WacurvBy8p0h
SuHg5sXWW0J29Rw+yKqV2POJdr9VUtfAS7DK2f9WpkOzop69K1L8OqfpGFwZdE0UG8vcx0tflURc
BOTMMEYx7WZESv2iv27lHMLvnQaniGB4OcEYqp6d2Bc6kBgERAbOsXIpk6gfvwM1Iy8+LB4fK28h
jJDqzJyYsEbDpdLtQToGdIufBvQ0Cdp9GBITMl1xBAGuqgGkZHbuyWdmK4NX8uVWF7fG49h63z2X
1azGaUglMLsbvZzti8nP0olunwfmhQ28IYHCHjs4obxo8GqFaW6yDZRrr52jcMFgdPBWBewR2HPI
fOqy3BrnfwVYcqIwZS3oFhRff56dyU1RoSIWORJykCB7yHNFWfDjXyhjSTIBiYKnxj5GWXGfxu2o
khLRe2GoZhciksVlbZOaSzlVmRyTTDHlRvBngpOa2dnSVCJjB34M1eVCFA8ZT0wELTji3B5rKX+Y
IziPym67wV4HSVrybzx0WTzK2NJVRTM4lZ05srdkGmG4HieGcDNdYVAHn0tSZJ5RYQIVd0nzUOxG
AI85WBihnesTyD/zLWYfmNf6SyI9WQgNW/Fow7xlu3CWbK7n8+oYmjboA3dcgIg+M05xT2vzXui4
SyhK4bCnHtiu/EooZS1g1ehu3PdiDclpJaQekb37XvO5OMW4hTsCdc9twz1cpmG2NhkxPD1MQnlz
WNyH70wxVUpSZMH2E6k7ZF7mG2duKQjC49ia/Zbj6/OZF3djnWZkL+ePbQ0SC3GoEd4nkNVsj8z0
iZ1F91dJ7k+Ffo9McCwF2oyDz+zTrfUuS33OQnjEiYgm95mda0+YxJBMJQiIewJMDbwuPjQa444B
Rr1q4FIq38lHHG9EI66y9qArl6Y3DG8H7hGv/OR5x+PqvDoXDrNoo2VgLhaL0FiZ4HRbAoNwqng5
Ex+LwxLyrdIu7TCc69lbgBUxhQuKNmMT9Xp9kEMtqlRn1/KWFuVlUqDUxiWxhLdZ7kWuF+ZWklXP
+FoNF/2dbgg46SP4BeDURXP9wjsnJX44cHE1p+gx1wtnpMeEqR7BQ5xx1KR/7vPMshLVaoflCq8/
yoVlDLiLUGh58EZ//XJ2XpF0quF+ZPu5gNWngWPXn2ItleUSzTMZCfbHXPepwGH+XrA3A9GxSsrV
hAqMviu0hgXTvfTRtWdzzjsdIM5Fx2uyI7tvaNTZ31alnil8MJJ6uJLDbtMXHg5kPCXLReMCs3b9
7HiFqaGZuX1STGfRjAcuUQuCID5Lk9wjfJ4DzexLX81eKTWH0ISpMLsBLAPY7wX94jIjarN/sky1
xXVUVWKsYncQktM4Gi7GTPJOVQ5aOyZUHuz1HHb7OUKPO7YJIAkgAQCEt9/SDmzBOemrfuj2Ssz/
+zrCGZNLHJfWzqmmor32yK4TM/VVC3TS4MANFKp8lDHiT98aI9v4HgPK/HcEWTAw3YbG/arPE0UQ
YD8lCVdo+3byWHrEpM8zZXyhnnytSzpuUeHIiKfPZQqsAOgug+byZ5hTAP1XEdIIYQTSiAC24m0M
HIkWiURNzq5CdT0elM8s4xtuXC6BAzTXSY7f6g4Zr0bkf2fHi3nz+b63rEfP3UAPrQXVCz/oMZVT
5pwpdTef4IqwMg1ahBj7YomU13XB8QMrEmpdRjDEid+O+/S6HKsMwu6421Y3qFH+2V+Nrfy4TXXB
SBm+Bi1Lp6ZEiuHb+t4sJOqulER2b3HK2aFJhonhvtmmXHOifW2pbvcEbrkRkAYbm3KtMq6Zmpav
EzN9NM7EMbWDaMQlqeDALtS+FqhzoH/9uKRNWnsby4Ps7g/zdVQ6Yh48H/GWpcMyAlfClIwBEmlz
mLikBsFFqw2Ws+mHQukjMOzjEdO43DZhifiJ6rmOBGQuLqh7j/FBZ8aoz2CIOHJ3XcTxeWfOLyrm
COG1UHtg6y3tCIFzdXeKrav1kKW0cw5q2u2wUgOJ4+iMeuLszSlkzNZG9OCN7hZESiAXW2jON8Uk
MxM8hMb0a6hBThHCmWK6zNRFuFw9QPnk7J7RpLZkAKnsgXsu/QCdMAor/AMQU3q4AV02KqGIEqT+
VjLTplhra/h3i08uy97XOKPSMwI/6nguTOJJcNtVjcXa2QVngmKBfChDMfLtucX4UN1hjXLAfvHE
5EGP3mtubHjX0ISCxdN3XB2ytwFMuaxTb2REUSSipPD3D3mdzznWoe0heXAtywAi6Ytr0yODNp02
XHbTyhUay0sNIfZ+BxY14kaIfgwtKlPzX7xHMqIKAvhYpjNcc4SIyMXbeiqg8rfwk1rffvSHw9L7
U2HzQlUj+wmH8OE8YfYEcQ9R1Dp9urSZ/rlN5hbFWOZ99QYMAEDpO5o75ampiuf1sh6CBCpoVH1J
87LAQr967vUluwo9eAauvlJtQOZ1ZL/Lk5UEP3KamvaVmrHr0cOr2A2J0msXA+DnDvimXqaaeoDB
e1cwF2FlV/p3FrP7VnBIJ8F2M49qTGlt4qPPb/Si5Ldu17RNborGNqHU0WQovh8c6orNwR8MUp6R
mKISoNLu/FfucxvA+aSj+Gd4/L7X+VuXXjb5cgKcuzgPLl/ZbttoI3pS9THs9SHgBppbkdUFBRKE
yIqKkWAAKGP2NczveRoF7sw3cjzQ/UkxWmD6yHG7TV2gi3/eEfOKHdaXxCtFGwal7wxJQzZ8CbH/
oa5p+2kYdj+GbGDDDzk3G4qzh9CueCDtnk1biRoWm9DR2r1vhBj8MFYxvBj7evSO/2krdUowNrZk
K5ZUPxMR6LR8M26ocQwu9yPziV5SEc086xn99fE5loPQ0Ja14PHd7Y6QRAPj6Cb+pokTgK7RKuKl
DL2pIe1nsDHhs3MtBahs7bmJbZOh/QPHF7bv+4Hu5DK8Dk7Dr3VShafPONSfySyswh6qVs9zN2iH
7fdBASWR9mC8npsoqxXFDATTvqCQwH5NQCN+sPX/BPQfErZjoyO84ptcTzqQ5ku63a4LZTVM7wBj
P8gr+KA6CTVyWg0sXdB8xpNpjX6Tyv0lMWnsf2IMaFuYhrB2FxXs8f3HOcuvbAbEqz1CbDFgFDNK
HORNOUsLzeNus9Sicd7GE+9JxXnTnI4tRDVrkufGY9qTFKmvU3XkgimRgCgfDPjDS3D6EnXCb6Gu
bhNb10tqPO+/31wq4ESKz5lC3cUtCOk/VNwWO7X/s4BqUB+tS+9Qsi7MKZxLPhf6WJWdQR75caXM
SaXuqB16lMgTWZbv+GNn6Y/8vmwYr+NrAv02FyMTN8FZxGNVkm3NNXMIByU2Q6jYSZ1+legyFjMN
iniDZdztqT4Xex04ACo4NKZ7ebj/nlRpfyEUA7pzhprO7L3hCNRoSLjCnjA/Ed0Z0cO3F9QjKrZM
9+Bl0Gb1OAqtvzlJWQxyW5lnSg9RbGFvTppiDqSaVFOGPEiBk+bwXZt+Ei+PjVJNdan78QXLc9KL
v3eoQrodhnA3+rc3BDn7SuqNdrpeZkJl7RJqmq14YwltR1USK5rghzVrA2jMEqwdAM0PZBpSlug9
MrzyF1b/YgzIbPKe2IlrvLUEfnO5iRCEPoSQZTbofZbGK/I7VcsVvg6LVBEVCpkQgmauLHaJv7eE
9QKgwyrcTaCZstIQspITvO/5dsA9LcWXP10hrMUnNywk6BYzRtsYbduuhghIroSM7jMuJSmgKL3u
JxtgZSghJdrOr0bYgjVMKs5ulSJJcBOjIWMHD0xXA+WLB6Fc5CwpwtPcJMwwTKHEifTuuhshxDpc
FAZ51oR1CUH0eYSMi8Us57zgp9wSuJYU/7Lr1R6TiPzI8/d14W+xJHJ6np666jgWZq2MbvK0/1wE
D30g4jyPHCscOa04OoE3uaa0YgEQxFlO/Q2EdqoQ9ETe6XXpZ99x7eoE9lPPzSCqBR/9lV5qvVwd
FHYdFJDM34dM1W6vQ8/XyWde0og6HY8p+2OOWR45fD1MOPFpFrxcHGdEtneRngNe3OdHkGVWvyEh
LkzI+KuYytVOzLdI1nm2EZl7VLlGL2R1/iT7jysS9JV9RbxSlNFcQNfeKRACcRXQmrRuAYvK323j
R/l7tsjSyiRyg56/gPRBPCmGHzCTrOxdDXPBZt2c21a7JgGUbRiP5dRE3JT6Tg7rymPLCrTbc5O3
lriOZzwPOQUlyqCdPbAlsPXAOOAihZcC1TVMG41TBWWJS7EF7cHcxnabykycIimHpPv2To1t7G0Z
9fchSVVZFC2U1V+bmHMR/xOv++1NMGWiG8VRhSfUXg6dxQHg0/qAYEQPfWheTxKwuwqmiao/3T9k
gm2LJitPfN5tKZcoqNLFpUHnKJa35AfIMvmDiDu0DHhaLe5weU/cPP5b9wDKwYg2tuY5xroU9ZT7
A27b7yop3U5DMoZLA7uVvwiRb59lp2ghN2USl6FPbOOozZIW5qWnez/6giMAoT+RHcFF8o2QBHJx
abn+AGC4oz/8Es34FITquYYgnHKwZA+N/4Wh0z69yXm3J7xkgPtjt7I0LJZmEIj0RlrMJjRLuQD1
qmHNl78NhvQSd5vgW0MKdbgGDl/Gugxnn+8rxdNcaNDyE2Q+iIPFR3dVv6WrxZikWpb1FsFIjO02
1Cyshf/m1rZcF/tzh310NKJjORozWHKPMQEsY9Z1w+BeckazGSl8Pflrycll6X4rQrqdvauo0tT6
AruNaxIx2BuxbdXdKBjm2xJnNJ9Pu/G+zyjv2RWR8lUkGWV/d+pDDNkrNRgJEUjuTGojERhx+dnC
+NPtnk3G4P9c+Vyy+B7nhTt9axHUanUkCzZT4M69blpmtnKr3VgYdQRNgvQlsEHS16BgktIHaPyA
87VeqkI62nTisDzSOezeKt0/VwaK8jpbHsbo9ZQag+O+uY6HWmAN1Fonf74kfaaX3BU7llyxASzq
4I8lCVj+ap5Wa6oF10WJgmOzaIy8p0PYFHM5GdHRA7sTf9nnegJF7mQu8TcylVYB8th/fNt5mhDn
Qbp2qTWdiMTwlNfuUJdd7UBkWnUwM/cadWeC5yQDgSx5M3Ji3ofc8mT5eXeB9xo/SI8olvo/JbQC
H/AkL4fg/zlkXu54dpQGRKnzF5jUMjrvjor3/DFwFNFI49EHbVhx1npRXutK5OzPhSOPEWQJiuZK
OZzt5ulUO3fAXTpH7TldCc8f+35pZe8B9Gw5Os/Kf1SiyzqIJchG0T0MdEWjxWP/RBUIC47hlXyE
MedVlfFDB3JEvMeyvV6JzGRBEx4HBz0pVxyiBOvO6Axg4Cfiy3x6MN28OJxpgSrW9yQx9IHDxh6m
azHeb9ohOy6No6C/AnEs9dEz4eXpvfZG3CvChtO7lZcuZK1bSdAVHgUplXOjA4relZxH+pnczcXO
QunNb6MIdtDub1hul2mFKMqQUeKBOK6oFzFkF4wROSRquf7KDNFBKaKbFK5PncD8PyoLocXywnxR
A+ikTTfwdDG7srHC7IK1DIrL7QmShPG0EUtV3v6+GweP21PVYkIKYtf442rl4gu0HiBDK19RDJ0m
709fMbTin5IEe00riiMQ6q/+1SKzUmmE35CgOjWit+QlC7AWwrFdgmJdbcqF4nX138HZuNNMuopa
vXi4N4vNIeazpxdrGsKh7tHh2qhTgbA7GOGtwEXIfr/fOdX4MI1pnbTp5fTHrqo/1kNburdvexN7
8FLcSe8FO7Ef0wuqsIu1sGntioJRVX6YzpxOeha8fj+Xt2s8ma7euW/82b1UqnJVDxd25KuYZGSj
bo13XZszjbkI64DMWSBQ4he1jcv/t+1498Vp6rtqv9EexxxmRULgcK5Qs5C5zDGGBuuKl0CGXfq1
ERTBaXznEsHL7ggp29mI7heQRRk4yW5U1S6ewVRP+8xOGkK8jDCvKvIIZdzgAE749wRVKIOXLiob
ICwNH3vwvhv+gAcoQiFASdMWSVzzZFPS0okbGojCgwCeTluKCMgAtVJRERMSs11QZgwwsyhJlaPR
yenV1I+MAHQ6BdgZXZIX0IHJhBKKAU/pPd2x0/Gy47jVykMf2U+m56cJPYYlna8a+sqtAtf2Ny6U
1csOm7ZBBg/7hS02s8fCnu/fLmq5rfTIglLx5fPn/Wx08Si/rCAR8OL7qSjkVJy0H/7I2JhsEfv7
vsmHpiodZWSbQC129H3GFOvyT81EU77+HFdOAuLBVkflUk+HvoWmz/JNG+SwhG2Ddn5jCXHJwNmZ
c8ove+//8uMseJnEM4iOtCme2/7TCO1caQ6HFX/LXL0mE5UvDzya4PNHIhgCQl+SjE4w0EEXqOQq
9P1J5KJ25eNgWYK7cIUc2AuTQXe7LN00N+5d4n1064f1QAAi7EUvexI/Z/uSjKhRdBx3N6Tc7va2
Okdkss/9fUMMh84yhdrWanhAmVimfP/KOg2a7N5qwtcnDGllEZHT4acNOVrsOycA0cJu/itNKGTD
HNFcseJVD7SQ0tU0SwrU9wqc+U38g5G+qnsZPPpSznNnEev4g0ac8YK0anXPGxQHYrJj+/Ynoj2s
2PGkOZ/XmHsZ13QJU+sKNB4p7HRAx4t1S57OmoUesPC2fsuPGjwwuU32ptWRTYqICJ7Ji5Bj68/N
+6kCj6CzKPSgs9V9HB3m7qzPuaGeglPJEQoHEJItcvt+4u56iJyLC4MUGlqMinejqeUdiADRxAmo
fs7UdjCfzyRg3zUPaTvjerpbdy34qtJjj/uCuhZ3uKKn96m7OIygaXGv2c4q4IT8/7dyBaEdee/q
otRMHtfq4flkZ6njHGOB839HHa6v7GDGQTOIkJNyO+h1q28eSgmgNY6tj0IMRhiFUBA0kw1nNBGI
Zjgtjgc3bOLzvGfCx3HJICDzakpaViMY6gC1PljWR6V98Lg7bfd1cS5Z/6AzOtATSSY2mnVEhnOs
uuNSKUbjonex8j9GhAuwAzjWbQTZ8zmBHVKDwFlmGEqUaQk2tw1AcUMDkD6yXlqygsvxq2f1P9rG
aA+2dlAe7PXdH7nXzDzAejOVuipDim/RXrC+/s3V+NBbFO4GMTojPNHyy2ufPxNHL3CTIeAZyYYV
35zmIKUV5uWaY5banhLpEX1edNp7zPCUBMpwz0NIk6qv5YDe8ImpxSIgwuXz4EHd4WkHSe3BicEt
qd7I2wU/LCu8uUfenb8athYqknmoyczGe8zaGmADCappBmXcV/Iq/LVTvV8x8qD7G7VxfeaQt5RF
NWRfYzQ4SPVrLUIDl3iU0vmBMM3CUHUKjQn8uol1txdzXQ/x8HPrBLsVTnD5aVnH6p+K2vh361aY
QbTjTycpRixHJi5LYVK4p++YFijXPn1tUMXUStIXf9WyfU/TV5OLvnHQntEp2beGLeJO7lEwWWMH
539OoDbGsjmX6lKfBuisxBOmdK1R4VDCnMzUTBMiV8Y+9xtcPGlBDkXw+JuuS1C6IbLT3KarjvtA
xBbknZWJLPzWRc2RbEsydQZpZlA+iY7TVHrmN+adlK6XJgoztbyrjFGoUXw3X1rZlUQUROXhyJOO
24oqh1UxU8W4daX7ekh0tT9irAwpdDdCkiwlJhcxbIrpsbG/CeFKexBhmXh2oXtdSOwiAKqyVVNu
BmCEvSEyXoeT7byZb67kPA2Yz0pcGWojg4UYX2ifj2soXKXN6G8BiEfpXmHosWtS8S0Vy43+MDer
teoWsu13iv/nOvS6WhzD9YIh0lNQzOwzm32/h9VQxDkIpK/Cj3jEmfwBLLpgkqYjvlSLhpLSM27V
dQaKyIYUmpQwL+bYnkv/CughbOYUeA5ks81swfNkN2drSL4cuFQz+quNKChmLNUI1Gn5d+fbq4ni
DDs1qV8KJtkfcRSZlJDpBo7dauBqk/A+za434q60ZG0HlSq4Y0wmF8U/NsaRqfK6AWMq2xw6jnxh
QqN9uYTzcNeIOua4L2JY0skL321QETP51A4cBv88TRUnYNYjdeZ6w7rzsCghvr8TW3XxR7l7ttOw
x9W6gehvpkv4PrrCpb0HSWZhhUcuKp5AvrUtopkDEV0m19fM8Duu91XUXYJ9VOPg18rDXaA8Li80
RYbYlju0N/OsQ/Tj+eSMcq8tPhpiE5Qb2zHTRLGt1i0u/ulrVNGZ/sW9mYCUAPohlXnawY9YStMY
qyVscOC2BE43jk1XwEfjEEcQN8h1XvpBhCDueWsg7Hd8x2+301IyALNDQWObVCQqQo97GhMgEqWx
Udxdejm4cBHUaIahXE/hwqwx1dGWQkcMQ/x/tXge8as1IWWDINEYZptxDtRZ/wkql5CCZOjeGRPl
5uE9cP3KZgKQaTuyuaYI86jyyYIJJRazr72fJ8l2iI6XAvQf6eB8NauUyaEjRfzoQH49rJjN5c73
RoFdaAtHJGttPYoKw6NjMfNbLbETJQNU4hIMI/tMGyT5O2dy6y27jwFN40iEfhyYEEHxBO0iOKBQ
dMEPPOUTdwPAiHdLDIIrZPcQCwEhiYo7JF1mAgMPfui+uIVq3RBJEMujxYClKaolezYrC84BapCc
ux+q/nNdEgXx5NfsfK0neFfAGpZBj4AvLDFVnffeBTAcshBIyZL3N9cKoMwMv3X5sq5CkoDdOEIK
czHiu13rQN5TbUUOyIqyhaBC58eycmY1xQvLHgilE3Fxj+aVZrGKxQY/Yr+1xOS1Sg85kBSPcuCO
oH9VVKVRB5lxBLqrcYdLpFsNUWJO7AoDRe4Cxp0czh3xqy10hCAfg6gMi5xWKpuTJUSjbKr0QbxV
BhlQ9WgGCTsS71LRlMm6iTTgB01qBfVM28UikXfXoNK4OafTiRnji+UcxGltraIEWKvq5OpJUjTv
H3rq9VpTzmIgrrV9dXZgB+d1zii/ni39sFcPKTX0DE8SGLtlBlpWbK3Ede7UL2/FWfvCmPqAE16p
cNvPhkG6EuF+M8xFX+dlUjtzpx33A0FiUT0ycdsan+e2kyqA9ldtjLUMn6Ho9o8yMZOCxaTg2zhu
ckk2RFO9ciOUIz3L6pCWtJNsI5tJwgwdRvoRGSemUiktK2quK6TEJrfT3dp2+JFURXRc9oHmFSIT
IUv3ya/a5OGvy5jVwf8RPVwFZ9intUqVU0QqI8p1vddQYyMFNY5FpbCM81TIqIBTet+Ap/I5JO90
2wdI1aGYwtkwGrudfzQQvpLrNPG/cWwIUSxSjpTsW0ShIElbMaUpa3rsLwKTvYeW+jinV9lPdlWB
8K6ZAxS7UTupiBEq3PLTsfNPm3h7dEwd+jy907zpaB8nJkndq5G+Cf2RQG0mxKTsuPFw1y4pYtF7
4dXf88+HMU4yr3/DR8gGWdcjzMNSA2qFoCeq61vLWuHnhnA4fLe7yRYNsWMMrVIXk0ZbyL8lmUiG
rlyiMVFS8b4xbuaQNzY0/8pzGBA1C3/LvR13SO95N55TydnE9wR76G+ZezRJludkzxSwY1vYRCPb
nwlFgFzVRyUhpU0xC2eAHwC3SmWYmY0H9+Q+GKaEACOoc951JdfGs1S/jS5SkS2zWGLqpqCwmwZx
SqpoEKBvN1FG9emWu8uYQ67FvOh9TjQjCKkEAZsQmPSbJfuKa0YTExDgF9cBw9SLggmCi800uIzw
7y80tzi+23twGMilHUyqLXgBPY63hZ6qULdYR3AJVJvtJXi93mzsmNrzYdZK2UrZacuSOBDu1pJN
MAX4TAAeRQc21p636SW/mMmcnYV5FxIMyyjiAccOsGgz9hRs/5w1kQyFVd2ZYa9juYY+NEWKknFa
pdxw5RQyqGjFQwpkOD9NgzGpjOPf3vizJCZPA6DHKjeyQ0ZmRgVlufO7nWST3nGi2NIcynbCqayb
UVORDwriK7QMNMaCKdAlHe1wLDqjLACf+Nm+kSi3EPtoE1gwjW36Pd2sxZdp5a7jkEgSg3ZdvVY+
HYbmc4tUbH6r8MoSUfpUNbUluu2Jd1EOAZ/w7dshJj0FkXE3UMgU0Hq+TMgYwRpPPb/3ZmMTxShU
nQ/b+Xc19WXRsNpIldMMauEP04iVMGW7sz3bU1zT0SkC3NLgwwfA8yy8DfPpZa/o+Whg0KC9KV0W
1g6JeZLtJ++dOKllrFijHIpkTKWflkOyViwjnWj8aGTaGmMyJrUSs80ugA4t1Q40wOs/Wjlb5Ixq
3zjA0LGbfW/2GLYJAOmo33ycCZbtjonGdoDQmdJLXikLW18ONLK5d7W2DYzWEWEhrYyJ7a0pWhKq
20cqgfDNbkvLIOch66zpjH9GvgG3pEqA+h3WxAq5Jz1oE2hhp/dFCiqOVxpyCKsgllkRvaDVoUj8
q7fLo5FNxccVvm8aFRSP3heqkwffMKhcS4lMBKKMPdXJX3CNAH1sJH0TkEXw0ZxuNjZi54kzUHDp
ZQII4xRkXqb77RCxVR3+M+MJMmm/E8jL83w7TWo6gsNfMJbIYzDAOMvQssZh8y8fiBQ4Vk7VkuXW
dN9CXet3T7ps7Va8RMDb88O7y3Iu9E7cEuqebGWsHkcHm+rcUMvZ0zibaCqi7RgCH2WDwQtOqER/
1ypMqkZrypxsKLT039atPlZiY8mJP/jrgw7LZyJhwoR7Hr5JWDy84AmQg5KTmAltjb876r2G7r7L
v89tZFB5AD9AYI2goLCEjn6EBfS8MEQDEWCC8PMEz6G8Ldw3SuQsLe9wt59zx00zJWfg0e4dK2Ep
pXjDqHChDLvPCckYpBWNZQGP8HfwSU57RhQ3K//RzXYateVfZ4kQZGjl//433zLbPZTFRORFVbeQ
SbYQH99rG07+1dQRoxNqsQQhwighdsIQm6iLZLr3oddPr6LGsBbirD+WwOm1qt7Y6a8TLFLKqbUE
RKubwg5aI3yX0Ss5YCY/ePSx7QNBOLe0uIKLOYj4nfRwy+8kNnu6HqEN+G8Ci7OIhVznBK1ljEh8
CLKPvWCyId316dswdoxn1TsJzuAzHtsqDjkeMQtR1JvFeUFd7fZf4cXQu44w+OxJAcVbxYkJBxyO
fIso9I5l+WBA61lb+BlPEsyNq3yoKT7WnSHc6O2gwTo4+RY1eVxqTDkN+2JirAtuuS3c+uAF2A6b
+lEIElNDl4Z6PCzgbQvr3GjP67ZcvkWDIZOcMNy1IEKH1075wTsg1BEZiuxyeb1tkt3a+5r5Dmog
8qxoKSm0EJVXJdd2WGa0i2e074QCQc4XfkfoVHruX7vROPZ2lCi4cXyj3XnIPXhsVVYlcxnOVY4D
fkM9qn2r5Ztdke3uI2JYWQ7bbgFCoJMVa3VGNFGga/8sChOQ6/s99zm6SbFQVmkH3+4LLFwF/G71
LP4LBp0Jp8DdLafkWMK2BdhURjeWeKoEVBsu/G4QHb4G3Ej1KyCeafTzEqxnwX5+rrFwxK+j7lyB
5sLTmDLJFhEYOwrC5aGyLoIUfcv2DMhKbSXxLPP+pFuUndG4yakcU4YGLSPHu3g5u9ZyMlm6RFQt
nWuzwCxIAw1B/cuvki0/QoYQOAcenBvbhlPSYMCVfAzCRluNciJfbVow3kBlsi3I/882iXZxh4kk
ubqe5K+rRy66EiX7Heve79wdeQkGnIcvANvU2LP9oYIogbLe9C0ukaLu6VoHWtfzl8FVc/UFDmr8
fohoARnMiBbW66yvIEpyjPcAwJsnA5mgTidt+EMdOEo7U75JmkREy92L0rhfXOEXeGP8hKBUYd+f
e6jhIkY2StD5NDAY6s1WBlkMUniTKGfxeFLyX3r9vHNS/Q5ujThjMIP/UysOoDnddXadZPLEBcrt
cIdeGEE2Ga9ZSoVKOCbj4melGYyNMOcqhf/WDXIrmx7n6gJHG8Qn2iJecIRK1+4O7wYQtPf2DA6Z
wlfBgU+s3QKiBrHRxhX7UGZYo8+3++6fhPs67UaKS8NxDnlK31+s1Q726LdkJUFbCMy/DsjMtDxK
VZwApP2nP2DJVRkElqGOWam+8nnn87WPVjAsgpndy3oc9ts24b2mMO3kQoe3KCOEZBdkUVAB89YH
U3sNARKcgGWDnKGRhE34KVctYgyWPV79rne9Sc69oK4htffBoda4TJAH0P/rsa9PZSfuOP2+NMEI
aU/g9VvRcPlDoFzrhlN7/ijeZwTuw07Mww6qvS5MMZC32hleX4n31JlD90TvDZYHqxIJK79O8Ppk
Uoq8hReSvqxtaAZU0DZRo6s9Adf2KqPtQ/c64U+ou7is4PjSuJoCkq+eHuRSpc6nJeyIGiw2Lfj5
+nMnLwXqIT0KrtA7CHCBNpUAzlNI56kHCrJ27N4DyG/6t8DVQDcZgAiD+TMgfl9pD71a2Q3A+zou
A/7bKU0RHnjB3EdLwm/KIpQYcFQlm+J0GfT+mGCnLL6hawKofaI1gU1jKIJeXvS5si5jTktt3onN
uGxu5iFu6Wxz3fFUvR/+Ycnf6wV8yyFINqAhDaxr4wnIC+A5nWyTchBVQ6FAGMlIp8XGgiTZ74D6
VLUpnQrj/8dAc82ks3CGfgR7cPDReX68L7O/eU9IQZsdQL1dfyDQZ2oXFNV9yqN0JwZ8lCWlNXp4
fX3FRgaDZVa5cmt3GHn2loKv12o37bqFXViU5ck78OvbExu8CEKO7JN4OgoTWBr+M90gqn1uiHv0
6NUJQ/Su+022P+zM2xEmsO/TFNkYOSNCxKr/XCCdAcdbem1rOIatCl8CebafoOJ9nKem793sXMkY
Mmscrye7MTdnirXTX/L8BU6wsvTmzJN5BF+Y+FCLHlmttri/q4Xeb7N3/+sgTs2Y99jUoSlWQNMJ
ZAaKjQ3nnWt/3T1XNzX2FmvzATPKbuR5vbEftOxSQkcapLezHXb3rNDaitukkbkY0m10oCwEOXVr
62RdeZ+d0I+ubDbroam+CXyZ5M80yGykpMJ0Utpih6SaI08miFW1rVyb/IpanJcEGHmISKj05/Hv
mKut91xFrDXT/nMIhijozLigv1WjM6CN4rvvjBVG87pAFWf60XYnNyKbhjnydOvqLmezUfj89V/Y
G+AdtLLUNvzUqFez+AO2fj64RIVDLg0CvdXofzzqQ4hS+c4bjWh7suyXJM7UpiNea3oO4PClgZ8a
cNXQNOjVz++iwX5UEhB4m2yHu48vhNgjruYqjv3KWuPT9tqWOWiO16hkx4kHIZ29BjsU2cWwje6P
lW5azW41lJKhep2wLG9QKuYxdvkHhBrkonzxL9j0CAukkLHc3gQFA0YQPRxdjOOV/NJO/f4+AiGu
iUTqL9nlz6/lsZGRzQNhaNKt+339DgI6KCTmJmy+E58HZZRP+6c483p1jrtQLJxkKMrQ5/HQhv0C
IQAVE6qlezt1s6Z5/0rNeuFQPAscAexQAvB3tPKYy/8PsB1sGNJSLbS8zrK1JPkl2XeXUxaQM3yK
V/C8DShyICabq/saVq98Lh3NLSJzAjVhBJe6anRH9GCAlL3k6i/VtQL4lNTiAYRclbLru+Gdjoti
Du5Fxh2Q0uKgRHihVyUSjwGMkoiCrQi0f5Vz8WuHhkU03C7a9/rGw4XB70PT5NAwtv6GYV+jjSiu
GrEPKXerLhBv/hv4U/r6BZvzw5YWGgp+c/c3jHmWtKAfkV/ai/3wduWbNkK3/WtgnSLd62fwJTXy
AOUg35JjEKAm2r793ZayVC2hoEIEm+Fqock8OpOnb3/YJ7WEA7RBDAzytQkVNU1L8fz8XF1/A/Hn
HWxnAbCh0uy9exvaiESb8zOVi8FE7kvUqAhFvf6x8RZXrXj4L4fzZ8lalcVVG3alaZdZsrRJXb3s
9BOrFhoh0VohAADoGVsjo1h/o9dGoCEfVqfI+SlGrXjDNxwq0T7Ihtivd5HhFclAG1PDVRCBSNcq
XPKSzpFIgrnLQkE1PYOIkokApBMKZnyxdEs3IEdpY8ZZELGvWNBDOt82pq8wOhlkAaZU8dw79kIr
Y95EZR+dcVkNyOiyscQf6dT1LGD9/TFn1tI/rtF69wxBxZElkwo8MkTYBW+3S33SLmmTjizRl2Ro
/kRORNJ9GLKB8GZ7LSWgTHA2efz7bN8jev7t3Bhr4hqDuw2NGtM7SJpDB9qRfzgf9nYxBK/puBxj
PqDorJEzTM9EUNzqUe16WqaDcv1aHew68N2zwyHroyyw3EoYxuKltBEETwinqD2+3ZeyPZPL3tKx
Z/geRnw1qpVOxmslxAmKcwQ1kcWjbPjNn66rQ/Eh33EIWjin1VTWn2tjfdCIutCu8E2lbxMBMTly
cwF8npSv5RDo/F2x3MUzYQ8qHbt/DiOg1VTloRUvEiyrIn2WwPYrSVReBmrGBHpJiPbfZV+egOpv
0rC49KqAPJ1B69Dh8BK7vpGIPXDUFYiOAltIviQuCKjEkbgLGbHK+KTvWlAgjmeENXtWu5r69oXZ
MyXkZ8cGct+WBABhxgxtMCcjwLGaqXr5ees53I4/f1eJDQkJReVgSrC47REK7VKX7aDzLSkAVIa+
A/Hkwi2o365UtSVOXI2eeJuNXnskuWfhgKOYy5UNUb+LGmWdLBS7cTRVgNr4GOHypoZ6vMiBX4R0
fWv3Sou844GLLeieSWWPwD7jYNR8RF/K2SqOMYiVeB2+ysE3d+LRvNog57z29mKKeabqTD0lRA2G
KaQm1QNxmhawksSPV66wqzT1DHQdrjYo9ZARsDyxqb3GYUXZucCTZsMOqARA1miF3+CXDmQfQGIN
KNIfTd62yruQIdUFrU0dJ+LILhXkccvRwroZC4Fg8+Hm2ee9vv0PT+1YFYd+G0iCmeNxrCeDNJkU
hWUnYP8ZvvHkW4ozjdwH6VV4z0+zV3G7B0fTpWVtvRwYWHez+EtOcQlxaUIJ3GOe+lxjArDUWsXf
Owbbona48PtdAfnnSMGXQCfaoTu8wSH6d+NI3g4lzYUvzLb1tk7VX2c3w0L6WDjUwRf0O63g+OSL
h/g/uqZrkDQHBk0BTnTzlOwPyrMJdbSfILDGWgbjdYZqtj/pJoYHfnO0ey5wTXyZrM/KZYyDyXAZ
zm11GJeKLsw4SUIjlmXgA8nkcajSptf+RFjQ0Op+/VOPDROPlAUiie7yYp7R0aS4DN6/Z1XgPngI
maf2OF/Mg/MJaOX4dWViNQLskglIfnts72/MbAd2MqEmNjcq9t9hKkLxA9b8fgpCP0SZN+v5hgnE
KuyZupDAGAy1RMeF59z3i2JPfByTTI95TfbGkd51xIianT+vsr5+wjFjXtpN2FIgnebLJEPIe5+c
20SZ/q0/RSh7kDTRdsey8/HGHURDyutU8C+yeF13HRb3ts0fi4wyIRvbyb1b+ZvugMqpsv+g8jit
4+BOpnJbnGwFH8dggosVkF6b45QanQilAvf+O3uLYJJidrKIBxn7MAdd0I6pkPha5M+ff3oE9cxY
JjE1nygJEN8j47kYuxTQkkDcsOgUFTJc1JAtW3pFUfblqm4oQYVUAA98bWKTt/N0iMoNljp/EEd3
OvU2W6kbkKO71bMbdAqrDdLI+4z5qVSUufyaz8j5uWyA9mUAKcY/5TBZEOTLOJxN4EgpJKQKIaUG
WX7tLwsAmHQzvfEc3nPH8iRQSkmULGNaBvcjmH21gcxmUPCjyoUEgz34L+MaiRV57YLGAzJVARCv
Izx1yC8/ni53RRHqb+UAbG9kSnFIyuBnXC6bWmJrlFYOczg4SqvVMQzG6aHMwC7DLLlgGME78AR4
WdTNHVuh0/djKxyTJhSRm9vRRUDOmlW/K3ByvqucBICxMS5JJ4Ti2EbHpcYbYGaTRJG+NS/847Ne
1oKhhwbp+wY53lgkhHKLeEqMsWPCcJIFfkkKf/xS/hyN5c/KTQ/6cc8KQEQk1DZzGcIGtw6LiR06
ZA+53aMr4ZUgo/Ye6786F6y2Sv1xb8v+VZ1jBatsWYTxPmttSCRQbgnE9YM4Z9tBFPt9Kq6PIzYu
rPYlX2uIT5qBvIWLzZrkTwupBxWcMxUxii2nm14sOPNiMdCXeEwcKS4Do5W0Qdzke4yChhT7kNHQ
1a+sZY0tTaMbfhXbXy+IVmyLcaFO0/PYpKHukSP+WcFA2e/RINy/3+BV+slr+jfqEHRAE6BuW+27
fdVFZ7ZjMH57HxQA5+QwF4BZ7AHgwyyWhBS8jAFYQ7OH/rHS/6d36RbvQ5sO/N2rs/Uojii9wX1b
xlm29RmgMATsSPVD4cXwDXE9r2NbI046Ea/wZsCasm21QvWuoz93TvKkV1+JonK3V13uoMGwzm6K
ZcqebrSR7msIjU/Cp5hELjdnwIQ9a0o49ywj5F4tPE0TRor4iwFoSxD6lUrIfGYKYqJIz7dTAyRV
sdaTRG6QWG4uS4k+mVHGsV5cc8G1fMe8vgoSE5gmhk/ezcvd0/FaAxE0H2uGn8LlOQIvrwmUw0RR
bkq4aUrItlZPfWRliuS9MpVu++gDv4WZyQ8tOynfNCLQfMLuLvrsmplAjhH3Z7JSSWL9XS1zwbyN
RKRr7UnbrBQzaV8tXj83WpNl/vVctNq05Ohy5z1qvwlJ7nqO28WJ3gh4RNF19Abu0acn0Fxpz3ae
xejtBd+fhInOelxrrCZuZ5GDEJ6tRZXQfPA7kH8OUjLAvnjnNVLoQNA7JEnSv33ptIP/zYAnCh0Y
G5LG5CtjsR4aIS6AxqxFJiE5zCfrgvodXG4K7RLITR0JyLLs4dGK3nAotExUxMmtwNdrqJ9eJfBE
aIV1au2Z+EjRQX5xp42ErmPxJkqkvfQbwidhPqxHihYX3jZXwjUSm4XxJhI/krlBZeZnk6pED5RS
DMNqlRtSypmGudyD3TUQjFe9HEMYH7ck4LtaEw5mGCXFeOIgjE8WXa3NxZzBWIlw70IKeq6DCm3i
EMdZjlZUpuIfNg+DaoUGMUvGipfCKsHYd2Y5mNt/h6OCmZZ/vfMqXcb7ahNJ6MGTAN5jeONWRUxC
e41GJ3aYVcLn/ktDb9h3dEDgTLmhz+qzpawbkcX1aeewjBqaCAAITutyi7vpswWzan4nLoCrqXZW
VqrP1Sqs0kyYWiCLGr/TaUmMgW+cCsMdNUIo7tybVvV2Mja1gGSjBZJPdvxpSpMWFX/N01vVu4WX
u5sBQWPGUmv/flxFMvmWtdBQX+pJCeu8t30QQMZesrulGpwO/dF1s9wvcs+swd2hXe5XPYEmb/PO
szZ5VqZsYV4Hke/p7UpfXV22jfyGEftEC2wYWyp5tMdKOFKagobLZj1puxgWIt+bsW98KapDSDO2
D1W9r5np0dwHnU0Jvc4kktZtlBNVwSvRfTVtsAFGDzihH+4Chtdb2gXl2jdDo3n4nnUrAKOI3YUB
ij9njbGbOK5ghhNhdmy8Cu4z06alkMiigdfog6O2cdFNk0usOEnRPf7l1wxTMnmOdWaJi3TjaFtu
iPTZc0VxskS1v+7cse+4Q23DI9wYcGCsi/dC+9FGVepioKChwEBYzdHRGTfPS1HCTrz6JyVsKLuf
aJweOBwdIpEGDh+GzIeSfEQbrmIVUupIVXNxYDvB5g5NIXgvXSiXljniSe3SKRikHsEf3Hit9gGF
Z23wgdtJxa84VY6AJl06co5kQzE3ioKaQx6DfW3vqLtLyHoxjt2BXEpIecS3JKIRe+u6WfhnaOqt
ta9fRa6LsDosJAS+Lyfe4LJwULzKsDqt7OAfs0DdFvQxGfXOkfZRQ5cehgaLEaTuIZ9vW4w1/N72
aI5pfj+G7TNnefxVqUJfKKcs1c8XEw+YsyNh5HpLS4ziG4pe2k1WIpmglIcfzBRT28oUjGQ6NGmG
jARwH94qAIGjH5cN6L+H/zvalJW7fmWPTCA0Nw/NlT4dTBczPNWqpx46wtOa4qxTWy6SdLGNXdB/
DZn5o3WWGPeepAuyNbzKVjre8r05A36Gu0O0JzYyk/Y5/l6q45RGZ9uAXvEq3zniRbwbkYsPZfBr
DGC30afhm4yE78bIiR7R0Y/Wpb5f+am2T2s4m7cvlv8OFpW4XGZAMQhnRKcy5h9eIdJvjTWr7vji
CdzXcJwtBzxNNPv7VfqQ/HAmUYEnQDo4XafyGil/MGH3cM01Eox95ctJa4jQF7QgyTdyke8W1BRQ
CJcCf6uC8iDqJwSrZRGt3aWWTKsUCCg+smskqNYz5RSrHFsQjWv+NsC+CCvpQqyeKNBwoqfYwoge
LZN4XZy/cLEWeyzrx9lvbErhHvMUL+iAXAe7Zyrq5YMJvppgcl0J37RwC8mofg5l6OLcG0Ao0eux
nzA9q5/G/jmIuVev7bCRv+cNLyUKT/QNK8TT5eZldJyuxp8EdLLqP9OGloql+LRbjCzedDaZD+DZ
kfxIbhqfZvdsU7hV4pbU6rvubyAG5YI0NEeWYRNlBkrsNkGEKkk8AufvF96GWKlT0Ng3JnRF4u8/
rofvekB2cpZEkZKPJFFvciZ8WHkuyM85Tcg88xdCVneJQn5nFPJ1Pcm9Mr67sq0dpVonXEp6Ntkb
k5j+sdNeWBqQuxvygrJt5T5HIodtH9PPvl/lpnZJwJNX02e4KCuuMLkkZlvLFHLcbhA/4MXWWoUq
ThGFc2QZ+SbORwZ2J6hLnIPhLmN5swq7JDdwcEkwWKmjlOHx3G3nbdltj/uPWN41/2F5iD/9J0Ly
LSLVdrseHK0oTFbxGqGQn2TGB22HlygTQoIu9FOn3HupctOvMTtyUnNslTCD6MX7fm41X83RkbkR
dyy3cXleGz4AsXKtgH8xkrKu8A7O3qjTam/gNCPyQVVX+S0SMwIuDlPkcjFMI4IY3fp4j1Nd/FB6
6UrQvaOgMYLkcJbn4fIT2oUn5lDsvFjFMkwzeKjPj5Wga/C5R6NzGecQ+np03cKHYE6i4zmeoQsK
ZXDmt0eV4ZTj4m9Yqo/O67d4GSZddHQRvuhWfA2gFBwofu1RgDYdF8yh0sff0wisQVJU5xnCRjuN
pmzP9vQCvg+XcEkfZ1aQy94nb9f9pjsrwc2sTc5B46kAaE9TLAgRgr5saaary85GbBGiyQpHG4iI
tr0ao/wHc/qQuYeJ3zV3Uc/iQOpwDxh01N0h9IE2djkny71t9MpF07Cbz2FXpGZr2PN89PxE4JTQ
00/Sk5hnNFSSDzhyKsqXIQYd/hm6AZ8KImfQUJT2TuozJdOeNJBEyNyZ1lJXR3wMroh5TYu3pYX9
s12trVR/EwRkRQNHrbaN/uXzYUnDW5hrDURvq+HOyFKp2rndLbGa2U9a0D/wGo3TotlnVbz/KyIQ
Yo3HWy7EEpFtisVPO25Maey1rgXsBZb51/MWWUgFhAbPv4b8z4z1nZOI/dOLzufXxQcNlQtC7cX+
RcRS3mrr882RZA/KFU0yiTRl+ZDWoWaYt2sbVVAhKasnxYgxfYwvmwGKcATWvdaVO77LC4vT125/
7IDwq7bRAQJKuh1OoIUBn2dc11u7CMrIsU+wMyj2IWOAtJy/sRnCgsIyB2eOcb8RNBgnVGPCR3GL
Mp9hhA3QiacOAigcQs/Y6AkZF4/aNrcGaZXjs1ChnBkcGM/5h83pZXvpwRoHjYqQGv0CAwIilRHU
WvSNU5l/7Ib2HLWGTlTNXHobZ8LhiYqpjHQZWyWoi8udczHdjDHrfKnR55Q2w6tOLRzTjPt1IFAK
1KX9EHd2owamtHFHEE9ZCEeC18IPXLbLG/r5Pfb51e7UXcf+o9k72+7YYpoiG8j0H+Or9Wel9JoL
sfMD53JyNiLF+Oxd7OxoMVSLPzDWFkIsq9Io3CugTYXmlV+wc9g1hP8OA5E2ExjQPW2TqxmtRU1S
U2Fi54bPkDIdtGBjPNSTE3BCVzyRIoL0efh26+jVbRdg+c0wB72b36A6aaBeB8Lk5Q8n2c4yzi/Q
yqX23vgmJ9vj4tEeDfxG0LkdQSddYbxAkH/trjydI/D96nWJrDWCjWnmN3i4UCCcm5mKaR6mSFH5
xFwwMGPrq4HYD49QrUyj09Tq5kNbEpMEjRuQuWM6GlD/73PedRCm35jMF20MWCcSlrEiqrCGjTmd
vkGkj4o4n3hnYD0G760jMlo6hA1+bMt17b0h1fUAwqpUPpoLZ0JiqZx7Y1sZsK5Uhl51+RQJCsZx
48HPDzMwMikXvngpXn63vGKe6dASm4Z+r5NwDpei9zZQ0oT3NJqRSqQYQDbF+OWyt9Fg0EB4z53N
TA/wn0mEka/vobVzN6t5PTeIL/qkjP7PELLwotEd4SH7ou4mqfdaOKpRFXhAunuWEJe9UPripogH
cZGw6CtnEx3K9jL3HnCSZOHJxF2hc+ZHIuejdecSRV9ABNgzaeUt73ESerYkjvEMGK6Ha9yhVYPJ
LjsoEH7+OnYb9SuIN++Y7HGWn9OAgto7FMBM9lmSf0mrs7f3wbFbYQk32CWvd+fb0KLYKgCPEn/H
mWTV2LEUUtmzk3NFnDNTasJuph+OtBIWxzzJwtLBLIm9mz+y9FWv2EnBIpYdA4//P6ZsY7fo7vlT
AqYK9pu5wrJiaLDUJJJdsUaL7mo4Iq7DxODzlnfMIt7S94u/ZtBSsoR3+ItZYPqDHnf+nUoOPi1o
jOBC66pZzPa2e4Ro8RlT4njo5XKJQ1i9FgJh/sqechhlJyOnBKi5n2wrIA5c3UWtyTX3YCm0kiPN
RFVH0x/WyJuf+gAuYtJcHIhSr2WEdY5ZQApwbgPLAHWBDpCEkzcF17xg9Gf6wF884E992uRy7+e2
1BDbp8yVi53thF6JfSK1QpwQ1k5TwS1AVtOYZR56gdkcKuBMpnuAX4j8rEk04GTxePsWvEwhHpue
uOEVBF/hVUt8E0dywxZLeF76lULDzaoXhy6LN/VZ0jlXfaSbfidRUvh6DIprkm4Zn6m1uS9LnfIe
+JUdgsba1ecNDBXgR49OUcgJjKDIdkYMBEIzbRGuU3nc6vjRO+9kGq5Alv4zX8RNc2X2Kj2qdcW7
Rz7zSa0Y+CmwaDiCBM+9v8PTT4sbFBqqThZ8gzRYmlY2EqJJYgqGNo74oBi4KIbG7jaNEY4sMmUt
GIo7FzCGSaRBwcLPWP6JRk4B4+m/rQVBji8pZ3mDcG+7MOcYT2BeM7QqvTFZy3xrsdICevY6FDEf
ukJ56lxwTunVAp2KVKHnMdLiKcYox4arzCX2dHpjPoE82ITVrSnuuXQUXIcKnhad3M8euK03pBXv
pfWWeqv2O+3We/QUNMY9CcHd/k4nWJEYbS4cmOvkXdyjWZkA2bvUuBg777N3TQIdVXuG51+qv6W9
Kvk5cTpfevrW4TynOhOpGDjeCez9hOOVs6uvcb1tiw0J6h43bftPL4cQZtoaDHcVpESuO2ps7RYi
YdXfAZhDWjtgEQG8KFjITIGzbByX5cerJwBvkNVBL5DvwWrZlbPZaecqUZUmWLwv/JGFiERDENpV
0qUoy9OC/9LxUYXbMbPOQEyZrpMTY1hnyo3zn5XxvmlecS7NmPBi4EcmxTSNp3S+lnoLqrRoX3R+
7EWCmr8Gm/22cq1N+SE4nf+MkzP9voxeSkNPCNkrlvKsM329bIyIh192iRhPXeIDbLhARE0Doy4Z
IMzyaSeuz/X+zDvxO3C9s4n8bFUomeQ4QOieGnzC+R0Lw43GLTSoSM0p5ffD5slbv3rbprM+bL1E
8UkuDZtchm++XTAbXZfjtFgNqSzF8bsaNs3jV0mjqlRr8654LG93wZg3UkgKyneqmhb7rvWTkysF
NsDzcSJJ9Oxh1xmchzmyu8VQHvqDuU00GrXNDAjUBWQkeVOP0oEheuM2zubjcwTgMkE+kTgV8WyR
Gc9AaFuvqUVxXG3wxBzRxMNCW5uw1zn2LmgB9wQXsnzt0atnpUpeIztCwVUHsqirifLr8Bm5/qIy
EfBZ9l5XQiC/13Ll9git59slOSNyzIXaLYbS1oCWrRmacbcluW86d3gWExUJYa58Hm73pybAbTD2
fgY5Y1NTkMWl+epDgPsdE84actJbAybzXwo4XB19xo3B+5koW4CSgnze8Cd5+iUDi67GiOLlhUrC
JSIBdn/L6q0z9C9WIasjpbm9AR9F6pMKvaPLP7z6yLwqvdiGFvPdrWStjvjptDHHP+emvCHzWKCc
tUnyIZ1N28dRNBwAc6QVYSRDGNSw6Im+blAWIulgBB8Lj6YPjGZ1/v05BM0n3Ti7Vz6Ip+jLYWBs
Zc81iadSIChKl4DhaARdHYZiq70SsX7jfJGCyOEkLHjukJ16K6pY3VHKBqO/PJoXoNlnDIZ/NOTl
ZJxFwONfYcMcBjudavWTJpLrvWr+yxDBOTomX84Ut81pU33NzSMiAMRK1WT4jP4keiYWh+IpniWp
0ne40kW6Ewfjzc7woaR3qNRF945f0hAV+ciu+6yznR9VGFTdZEQUUfLlDfJRfkv27IZWgfrakfdz
QqolEYCHFkiDmSWI0gsPKpRftEYGb0tfpeclyZQeEBVzIHhrTXCCrHtBkNU8s0JZWAwTlNgcLvMr
xuChb+fZGT17G6xdMvXxLmCejVTDcY+AHpKFMmP1qs2OsXQavWp0WxZagd4fWs62mjDUWEeDb8Qk
F8bxm2npm6oft2eTVww9PIEcnMrni7rVcJDZ8hKxXJZFBwKNae9Qm15V2jWjPyNks6zLJy1WhFN0
0l0agnh7PnzXnJz65P0DfT3/D111HWali/n+BLgdLBw8bZxs1W801s5yOFjHcSciEiV+o7iMSNV9
7ZGAlfaPtVfwgITp3cIv8OKAC//OYbqtZtmF1iZA1fAIs9g64/R41RJiG3EaEF8IkcSf6AkE3tC9
9n9rvBMKLUOf3jR3/StYP1v2IjZyxnKsg1HkXbQpzLlrOSrpMzdplzqdC43kbAb/GTL6siVcNkGS
rEPH8Ad15Pl626ZpejSmo8ZfmKyc1QSsjgL0l772hRUWTqWP8vfYjojnsq1wUCXsH2sGuCptyYCL
3vk0Ax8+AxwMOKfc+hH8wVxJqIwiUIp5sIda16nYU4L9GyD5BtzRFyFd8Oedarnct4om5pvpDc9K
H0fuh6C2bI4fzOuMnejFzGmpnCJzOH9lbgk2o0Mc2T9A9mmAeEdhkuHQA5Z3nQ3MYQ07tfL9gfKU
ktVfSErWfBXq//S6ASkx8pMPrGY9PY12pNyHYyHjj9uJrNg+vHupZDm+bv5WJs7t71znMI8nffRR
i9+SAnEg8JKa5yMUdIQK8rGImmIe1YsqrRX7dCP7dAchYOLh6Q8U13ld/HSbDh6o3p/0IwqvFqj5
Y8QZ/Bly2QSkM8OatAyAjHqc2aZGBAiwe/asdVpdSpEIb8Es4oauScnC1lIc0MHAEBkipEPwM0WP
QQNXzFq6iDi+YMppAPXLEXeUBvvfhZFS3x3O3HPZOYFHwRwGA/x2zHcPH2u5BcsgvJs9JZlZZUb6
Uq+IRK+VlXivp+jcoQp1ayNS4CDwMeTZJTPYq90mo4Roz8f67lan+yVG/rElGLqJjRJtAORD9z0M
5A0QCo62o0DjetKZf53IuT2/GK3PYWdmg71BBOsVtbt5Nc7IgfrZfqGUdRLQScGWVfVgC6aT8YiS
804G1jz2c+7Vlibiy9gCTyKak2rlkmtyOgu2zO2dXrcIBaC/tlG1Nix3abwFK4bRV1uyNJkEHkE4
unlE0IU9h7NVFwI/E6dHxJ9C/huGVkPwlV030iop6AmTcebOzGcXmx7MgTHOxAbG6u4MInaGBMpc
hTy6Xy31W7i+i0QOC0hDgG3B/vcu7gNLbkRDgDGgTOQOKENUoZOGckaGxaAbeUDTMxVH17H+eE+I
3SPza0EHbdKtxfjO8cfyTpg4rNG3rX0FhSguCoRICfLYS8JEfG81AMmItwFTOQ9R/spFxqZ4M5tO
XLJeWq1lGQeaQ3BdxxTNQ/iYgLvA6KmoUCSMPKk7SW4DtKAcsJQDjWm9ksqzfDiKezQecGPM8JA9
l+FzHn2XIzsj1VYlrXowUEu5CTtZMLllnI7ozFhV4MhtbYkHOl2qr99zaz5WPW6r7wNbY4CWball
bbwU0gga+X7RGvZhYEBMkvQIYQa2C1gwCRm02DzUoJ8rgcCCQWrayno6mF/qyW9FXfIVeCtYcVF6
+YU0KCkC+gT03+ihP3AOTfmzBsuaAq0wbJCzEgdTQ1hswWNSZEDP/TAag07DLDVmiG+TZx2eQnxJ
qjHmbZjk+h8AM0dKBh5CwCkqFPxeYSmTGYfENRJg2n/DcFb/ZIhZadSV271CNpCPftHfeWFLMU88
RLnF9m+izDh5lUKMe0rLwGQGmsl8fh5BBTjAFtG58saKyN4bYgNwadTqhTuvil9JnX0uo84AJGkK
hQYvEfUvEwMd3t562vZlTa4dYD6MWcxHjIjr3LOG6PHt9zwFXM1eoIVgD6LLYq34zSjFVt4v8JrH
Rc58ogVZMaA9lmcz4n8ntIiSyIFdnY1alwHO+r7Q6RhegHgH4lU1h3fgBMzm8zFxkzboopt9/JQi
wYO3jaAUFEHxjcxoWJ3yxcU8xnexhBFupDObu6JPd4xkZIwZGKxwrPhl7acVBzKqz0bsEZluymXK
sc20Sp8OhvfL0eb0f9ZpEE+qx0Fd+wmnQbjMEQRkuGsmDNKe1RmWqU1HRVJOcM/AMtT3PiqUkGxT
YQgF4IS1Hropcawshp2RFTJsOA+myUeJHmsrG8yhi2bwHqH4avV4UJxpFkJCEQ3dSMnI8yTCEBsf
pZKVOLcG3i84jCEHs3AtrqczuobQJcTme4zN4zB8D5dfRTigd9W3a2Vg6aGgYUIzHfrN4A74Pyzn
A32OyCTOHfPTWXKY4FvaSO30WPvZRTF4qMVG0IN8S/Us2A3FblbtgzRnpxznM2dVCa6uvsAH1L73
zP1Okv0PPRntSQIJEHR6GmFIqdl9dzgHlxVwbfxISRlia+mdCQiiC7vpFPJ2idd0BORK8gyjtrvi
r589r7XoX2xBn3pbfTtMwXyBNdtBjIUUeyXm9E2Xz88qQhnvPWVz39vBd4u1cS+Q5uJy4CfL9wwu
46maKN4HIlHEC07lh7Z0Mv9+DnBG4DeKYYopj2RbiKtjzvEyGsq5UVYQnrBPLRBDKgpoXNB1bKPK
KrBd+xCNgSBnasOVotKXneF4gJ7CTyaYF387UNjC8T2jjys6T4UF+9pUdAVnZ20EFCYhc3NJUTAo
UTtrjG30qhEd0WXVizoO20YTXBGSXShNXiWuHj/wvxGsTnrKwIvoCBBbSGh5gOH7O3JMVtI8/u//
J69TIO8zyrCAqtCwdfdgwE01DstIJn8bdzGekCHTLBcDiyqoqarxtVdDMAli8vc3/Fux2eC+iggH
W2E5PMOmtSrM5S//h8d5l4ijulAlL5gvF+DTPZxg7p8Dd5mtWI56OKW7jZSCKPDS7NokbZMwR3zd
HVK8djVx14+NLu3tGZVvkND7ieiRWzkqIxlhCdI7OQqfLGPSLQfgJLQPAMViQurBYTKPfVwe+zC+
naYDzE59rcIERGPWZJys1Q8AwN3zxQiV7j3KmU/snGBubrnExWBmdvY7hLWDF7MPNv5JGjPg/Foh
H5wosN8R5J0/8XRUoDBEMVkyBqjhpLO2AvW+vmTassOY8OpKtHe46Gq8TKlcFV0Y/4/PNPHjDe5S
myil4xLuIkNpfZLWsnJm94dTIBP0eoV+9fjQTBLg95pVGWQBzqqSnWrcOh18wiiY16oDWNvQz8iG
QJNUenkVk2Z3DUjiijuwRunWComgWH3Gs/ZN4iBXtL7we46bMF0lasPZUWmGhAIGC4+elbF1uVxH
bJiiJUr+k48/zFGXd88b1oNZqp2rj3D3mpUA6RfwRNCBlPZmWLRqhdxIUAc5uQL2PnXh5cKmCFIj
YD88q7s3pHkKkQSXDbYD2T2I0uhQ1CQg4A/ZdYiG7d1xucWQSooxF9VIIrchRe/Ed0vNE0rMBEVF
E5YP2Z6eUS7n42OQevQncGnYS8BqEZOk0YS0Go/XGF1sp7O1eyuPyuZtdij6hrxjpGi3Ptc46VBA
G2v8L06yRVlUfTcGSq7UD4I2nGLZ9VlrnsN03ZTr5MtLQinmzoOC0qLNXhh91z8mIwegrq0p+vy5
I/9VcOpZhSZVY2plFwiws+SKsSensugaxJPSN/OFpi4eCsA3gHu7GwTnfrrlRo2XoOkhfil1Hcit
Ed1k1zMMeY6AMQeajgHlVeAHMLrVvV1hy8o2A+NeW8VOvO375s5mLeBFbIjwOA37+pOzu/yJayjb
jIKET2PgZuUC9QOu1yvzRTsws9ZLxBVlI/Rb+TIFcswJjly8/h7DRFLkdS4A4qQ5CoLuJdW8CCvh
onlXW4C0AXPMLLDOWvs9ZHev36iNJ3wixZ8dcXfl/L7mq8Bfd2YgwoUDqbC+iKcROiKUI3S/dsUr
zezZfeJELifB4V9B8PnHLx3i5wgIR9BIpGE1aDfd4cX7PmvuI4nhmPHBDb7GjAVPafmI34ZyeQSI
ApMnQmPqtYkMFBv8mYu56yCdlg0v1IXOeeKr2j0vG5YK+jImthgU9E1NMeaTTd85vQ3P23tzPerb
CSPOBXwdY/f1JAsBT59bx8ZQPDvGbPnuEj1c7k6kHKRSQ6tA7Z5yJ22U3hHZeRkhTFSOSeM4LSAq
/slIUbsAcGiq5niMOqMmhiFAjpgKn7+pB9zz1gj3LMPaajxpRCQXLZ1tnJDatXbwPC7I44i2Lm1V
xuodVIPxvTZWkVB4oFNWXgBgf2J4EDeHDTB+1TOvHccbs4nsQinAfUJmB6tAwTfApq1dddmb2gYm
7J+QL5va2XYqkH752OunRmXUdTd7hXj25zw78QV2pJOct8vdO5ef3VZKWFc6A+XjFXrW78qk8INb
CN+KR5GJw4wjN090b9OZrtwecquVpSOHg3J4QnRm3ZNyGyzYhUK3KpzhgbA2T3qE+OXlAkj8sslK
Vom5DifQfZNPT9H2x4m2R5VP5Np8GRBKtvFIDPlXyYIOKqVK8i5zOK7zYS1oTBYnEEJi4lThmiQI
bz//b7wDSDZBhtD6Qu+tOeWF7hczA3wJn1XBwBbYzKkQzkM2lh/X9CzQJLPZo+h05+T1DPuOsQ05
uIeUPkPH0hLNKELlYknhFxjyV31IqqronAoyWoMugbDj5/iixNjp4FaGFvp/6D+vN0PJgortBOIF
F10aEP+H28SlFiJLZJQ+0orXOHAEpwvD8Iy8AA+JxCWO0DFGxdm4tSOH3lfraG0o+LbZkml4QbYr
JlEbBIINGcx+ZXRxl5CYM4skVBcZmXHto+jnVWPJfFfZ9tiawS7QZu7m/bnfbYcWEy0TRvVflB3y
g7n397aCpXPf7vglDfKzv7ld0Z6ZUBU8mvVMV5E54cHC8uQwDvD0rzZM2TAH1VyvZsjZLlATNaZR
VF1fED06RBjdMQFd0rSf5+nFT9zBTPTkugw/CZ83N2seCXDlSuqcBTGdjwmAqbMl0EzvCASCiZAZ
07WqkN8ZHbcVHUGD7SXEkIh0XoyG8uI6YO6IficBNgH0GRIpOghNLboqadkYqsz1yxaty712W4Uu
sl5iFpQl3sD5f+DhH5+AHvpTBXkSZEQXcGhXMI03CU3YWr4F9Z6U45r7QNwBSwIUnblNuZBU86Jz
kIrz9lUvCwC1+uksbwo9xl9mh8u/LFXTZ23MKWUrs2DoTI6YDfu5AkEO+F759W2wbUFGQtSQ69+m
23c8giV7eCwRqskMt6Rw632diA0sf1pouN04YHPB9Vlz+26S6m9L3uA0ElaE2JO9XRdf26Bz0rGZ
7piYThOtnTQuJ67/sMlWnk5WxPsN9U8wcoeGZEYdoY1Si8BNhlZKEgSoCSdktP18SW4i3kA+B4Tl
Nj+6+NlhUOkBw9g0RTwxcKGCni5auynndwT9SdHfl8D7rzhyZ+NR53aQoyXfp3u6YEldcCZEgHkk
z+62mT2OOx5aSmYdaQ9yRVkyNrmfkr6CsxHuGDQrAGLG0GdHsogDTSXTiw2JfNys3cKQjpD46PRx
zXvhtbidCZ3S+TbAsq457UccaXWyznBEE3P2SLShz5PiH9DJwzSRqlWpWXW/6M+b2qBc6x31KKYG
p6PAe5oNC77IaGk8h+YUcLPjtWXBCw/7Swp8euDjkTUazCyOB7sNcrcTJqxpYUW44i2Im52IEQAY
NRoNoljNFswXKzUX8Qd2bLpGMEeyixIDzekG9wmJWpyO9gsifDEobmtaK9FqJoWQUN+YI2LdNqiS
op9yMLm5JxU9+iWA+93Z9ai0UUNIklgCYY/qOUWboKeguciJrJ55250C8VdMAEkILzy2T/QQRHtQ
rtLgmuk21aGt+ev/Zj9FSclt0MKkT26UxsTPamyFYmlkUtyEKdc1mjn9NP8VzwRRWI9orgxoHPIG
RlfvbnVPq4j1Ne1VoXZzuIy1FU3e3g+mFZvC90j8sBwo7IiHzrG9/qL3VIJeuKYVAlA8WFyvpmjz
2JdfmT8xsE26YyjvcClJcYsVtv7h7uN9evxNPo1LHyTH5Yi6fxHCnf3IQ8FrQaHf3pi+bioJxbsF
Ujr1yccifb7n6erR+vZ4ifxA+P0gYLjngLEq43HBVFys/XKlCyoAib6fo3CaFlcIVdX7pMl/Sx8T
A7So1MJpd3TrW4vXl6eM4H/h4djnwPnSb/EPkM4CGkR8Y8jSFMVrwcjZlbrNIG4Ep0uJJT47npgA
Sn9uRozFW36149ZeBzYfgmx4YB0XGHIzfP4MJJ9hWlobuTFMkwfDiDXmCzHyyihBFfaiwdZWYmfP
MDeI81H/Pid0Et8G1rdUzRoGjQcAuhrEravmAUCVcQcGjpKzG1IFAmGsM1NYF4JqnbPZoLDpjxo2
JeAeQ/875vQV5js7jWB50xua2siVQQlkUQkkFPi3cdII1xIg6DP+SKWFbtP7UJQh5i9K4hH3FyGc
YjkFxPtaCKnlbq9WMS7xghEIzwW3ReolHgh9f6XGto8Nf0M8qk+Ai0/GgTjik4PRj7PRFY+fMJ8S
aZSuEPvxmc92vnE/6CbOdMdVZBLkW+dapMu7NYGuS1Bq7updk+o47q6yB0tBCgbTfzayGkxO1z2H
DDy3TuB18C/Sj1czEt9Bs1Xcj/SxXnpoIhEawIoEQmJ+pVzEL5Id3pF9vtP55Qbpj/Ddd/AH5fNI
P/R9H97EDIBxYqjxUB8nL7ZtmmBJHrh0reawzmCcczyi/TdUtq901uBqjkp+Mkyt4Xi0JB5CuhP3
LzCo9h90OzMcoKcN/UU9P/fI/yGmHTFb1xWPuv09cAfo3jUNu4BgUtEIcXPS5pBYjYomvgoblOuH
VkKWGdfQ1vfFe6Xcbak9IIl0q/xHYjqOEUH7rip7MmleGmWIs4HgTJvW3tW1HoG5uMxPk9FUgHcg
BGo5kdCOL29TaYbnyq2Azi+ly0budy5r/LwViy1AsIuO/p4Zcngvbhhk126i9E2eJ8sCjNxclpag
IWvFY6ov44TaENg8gnoDqhE6IWNoKg5JHRe7cAfXxkbXjp+bCN8zDHHXoKA+cTlev4gIc2qIF1uJ
TEOO6hk3wP7y5VFAS0wNjZHfCGF4odHAp0AUZ6gt3mz8tGQT1zeo3ub3IfGLQ9ZE7rnn6RxKZiV8
sFaQqUDZM85Lr4Jg3vx3jHgk1E5sA3fQ70N+wNmr5oMJ6kJLeJuRn1pVh7J68OY+ngPvtLj9rQZY
iby2+ApBnr2JPiEOm+GZKiUwLtS8yqc/ZYApHkvBsdYgHu4OOU6UzzKtRjEYkRbQRxuR1ir/iObm
iMfr/OYsCJjhYL8ZyTU9gRlYJ59PgbQp/+ZwOvqL5nXxoVou2zUpEmtTxui93/4TWYGGhKjlxVXA
Bz3S5VEW9EYPs/wcP5FOui8ustU7UdrfXeP6E3uUQwC07p8gFVfRdLWWQ8VJbUp5pGxITuTsHeYb
anXzAah7rtuQ8tVkKvLar1dTPuWKjq46xEamBBmG+RfDyXR+Q0omMbge6GkK2isrKwNWmip1iK5I
ai9bi7swUIumXn7lGya0y3pyUGnB36EFdp2zMCfVHsQtd3ksMj6OCiCaCgekSmNdNd58Q9Gwbqib
6an/MI8tSBNfhErRN11w/41QMmaowjRi/9VQVywUNDcRaCsfLCmXTKEuWX4h0wrnbIhPgKDO4SEX
dptRPb6Af6H67NSs0mWZuH1wHPyMS9Fx/kIiwQ3CmOa/L6OwmCi0fEBG8J+XcKj4hbzN8n+sdP1c
SGH/GXxU5ri13p9eWSZGMOXIQ7MWJIDYO40TxTUsoQJ9azI7l6+nvruNdgcfjTT9dxcVAg9XSKTn
Pb/hMdPwJoBtr+/tjBq0Qemv8R1uJKuhM/CQeLZjqKCX8x1t4WbsidyS050Oq6NAz+lGJ9j+Sg9H
S8Ge441mAld2s2/l3g/hgW4VBT/MfaJ0T2Knh/HdgHmS1XX26q8qS2pHK80JZiNZohEZxrcNy/TV
Q6y7G3p+lfb4ECMWKdFu+YDT4Y8+sXI0sXITNZ0qn1t85uB9hfqESWk4jSj7ZXdxm/Mx2HRttgkZ
sxUWP7qk5SMA1RVFLPplmov6JEdORJLIgKTGE5iFdqDb1QUZJE8MmvKJoQcyU3GOV/gYbJw8yvBs
nATl1QQTnj5hOPoAtoJGxzyIIQa276W74zjW+P7MtHldhaEFUDh7GKLJ6fQQloMwus1x8erprPxL
MOJxtp7UcvjX4c7jIp9tdSQV9XyGP98r65Zr8lvLalYGfdvGMGocjANe/3TZlKBhbOsHDzMWBFrT
qYFS+Sq/SpIr7T0juKeJbLZkTHf72a3q5gZFLsP1KGGbnBVyqZB3851nYJojMIwdUsTP4/U7n6FX
B16JzozSpRL/SXwTMJOLO9AkxvSsr+mjU4sfjdRFSikQWJJF4PTOtMR5WEzwPrzAiERXnkyKigRO
8GgFxYilH41ST+68XiiTGQ8NhL2726Ha3DKDhPI5mYIrxUpwihcn3uWeoCd6iNB1AyKbXsL+/Jdf
9yjTdV0CJjpUl7ubpS9Qv8YU7ZEE2XGiljtTbBKxPxjJmYWbjekyL7GZkgE+3LhiFssKkEH8eltI
hZtD8LVQxdEAi/yTaUij+/2pknjOpPnalgRoJiXipPvlvSe78oJFm2dYf7a4h+Kj1B3vw7xtw8a/
ZcxpgNy6F2yQThjcYFUGWhVgTu4zfVn7NtHUq0vSeR0AkZaHgpogNCvtYgz3KX5I3Kk8yRhORFDu
QagRrSEoG8Pm8tqYddIXJDSYJ4hP2f7GqgZZp+7q4AMJjLa7iqHo2k3vBIJ/xxl/ZGVD+wwrNOFG
nqXaRtrBWKA7I+WdoWmJYLsVJKyRjzsAsobpAeY6GEfnJqBfiOG0Vct6rIN9PcuZ74kdaRY9Q7qb
IIGH4eDuvU8O7ee87w3W1n2oHhBaHjxzpbCthxD4hoMPQ1hAqI+1/uuA3C7RTy1rdrW3aRE5vj/Q
uY8X/PMBhDT2AetA/aUoli02esPEqD7/4tF+niW+ijHnqgoBFL+UrVzNGTGFTz8QeeIeojuGAdCK
dDZT2AfG/IkGFHW+rls+JX6bR65l0HcyBRsqIR+cE/qOj+N8DlnKwqz0yJODT+O9hB0YmKWIhB4b
JCKuOVetScbBRljhF7+I3rhGsN7Ip6Pw6cLvaBnag+OmQcmf3dV3sAhEFZIUxJ0E79uKK2dp8PUr
Pk2qbUVjGda2xomRDAcHph6tQlrxOQJ9gjkdnOQ5LzzcO6CswKkZ4OEMVytkoaVl6uty30RowYeA
uF1Y4jP1D5al460t+Q+XYMTDHo0Kai0ugbLkQURXkwL88SwrsPT3mDMIyZ1FCEUDkMsj6YvY6bLX
w4t3dhJNhkA5a5LKBUvygYjkeUjku1wGgAu3Bxio1dfDWfA0Uo3q0T03Q+cRdTazoiKcRk1OH2oI
rilMKUeyXeFokXyrstmZ+005aOkRqOp43UUjCzrSkSBzaP67tHZVisZE+r05qDlNoPLdHCUAOgNK
PcMmu3rKgoXVearl+6Y94THUux1OSc7OMIDP/V7Ie1yqgtOlDUBHu5h3MRZzd+hEQUB20/MnDT+x
lSWuQGz3Ctq78IjGZ6l2XjD0Efc0hXQi/qaNsLAGHPDqZTVlxn08+tN/fFCM7mcKYTedfw3XD1Yl
p+iM6a08Yn+3h889Jz6RHKCwWy+lSmJLNmX6vAGCY28jQ6teBUDvu//aXzLYH8DtcJ3tNqZbODA+
+u9DAkt4jBVHomwqeG7ImFCXQWYo048+4u8GdLOwuaCmp2vT0XkD+RT09U6Fbrv1LA8WHS5/xopm
7O/h0A4XhGw2U82c4ebBek4bL0Hu/T294ufMEZ3RZZhNMSB7DhFubjzXu+moIsRGi6AU6sRvJp8P
YBvY4V6VAX4PdroboVDZ/9AzE4UB9lq1G/IQPR5MVd/ST4a5os0PLcnwJKeVEyS91GdOTGC4yvGv
C+H6tWVB9kdRsttKayPU9OcS4Vk54GezoY6QH+Rv7sbkSTNVkp6vayAxwj2ZytFF9tw4xk9C06Cq
5dU/fNkC0L7SKtEDlGA6x8uW2jqEsNh0uyviuKIMsrpaqyFAh4d+/Qh37dfVPh72yr3qYv+4jE2l
8fzJp2ILB22zXx1V1ew91Rea3q5JO+Xzf30oHCdyxxCaQPwklsJ7h6yrarUb+AdlPVWhelsSUDmA
owti8AlA1Oi/FlvmUjAlpi5agYB5vAz5jBx3zJ62cVWiR4rNUlpocrkhRXeWxqCCObI0KRQpIxGN
tNTIrM9poBtPeQPXjMkcOxrxt8UAWSrF20sUKzeI1+dOtUo7jHT6JRkyc/g87SEBw4j+QTk+FtRq
8z88dU3qk4FcrYAA3lAPNdmYTKNBiTYm1hS8Z9KMUzq0wMVgEbXI/FrKHZdJwZ5L/m718OtK2lRD
arnI2tCPrO8DCVi5GYJUPImoWkb7acXcjrd6plJ1ZyPVCnMMs13mKBoaBSqwoZmoshpIP7Xinh6p
deQeUYVdgoOoIY8gV1ER3d+VZjQvP7hpDea8B6XvS1Rf+J4aBz4sxd6trK+//xVicftRCoFHqwzE
3mrUgO5F8Fo3YIloDGSnAhAAiqeY+xw2VrzGuvuXIXFmSmLgEClZKfxXPMyh3Q1OcztaPgFZDjVy
jveE7pkI3J2QV3jxj1G/63ei7/algyDgPrgpGQl2rAy4kPle4DuEZSvOojESRnnkUwXhMm9Qjyc/
FHaJjOooL/zYO375aZVZyld9tUUCxnomoLyCKIO1OGtbUMemxmeXlEUS6uOulo8ed+R+imSvEwwj
mn/MEK/a/DkYTsAnVTF5Pu4eZ/kxlVSFpmkdAhgN+i3HTL0m/U7aGc+NpK2nKk8r+QfsVx0sAlJM
6ibtWxCnxNaAW3xISnFRpsCDkfpvckMd6mjEfMbDhxRmioA3LIOPmtqf4RrXZqHFN1na/5d6jkJo
p1h/jSrh6Ra9DZ7r6aoIkZJOygr1M7cJ9jLslpsVOiqtM3C3HmdRxKZUnG14dupsswuj6GOll2zC
XqLPKL39i09PRCHM3AvUrlFSm3PhSpqhuKmzX6PXRx0e54prMRK5y0XotJgHpxP/gNpOUD4mluXl
pUx6bYvHjFyq/VWQSNh1dYB3ojppePzC5flBOBnFSJU3dlOYQ9DiHJmB6L/5LX/K7dn1KfBHSebk
58sBixjTeNBF17Vo9YIRPbKAzQ8yEc0nD0Q7cS8SrVU7SGCCydDeK7o1F70JH0YFjX+gnqk6umks
N23kYCQSj4FeaogXcq9B3nyQle7/WWHhEqTydxAsWyEHzwhzxawRWPkHCCbYTr4Pt4u22sjgdYrf
dJiuqUHpEWh/x67lWBewNBEBbOvEhHg78BlKlHIw3X6ZUpP/5XjCh1lkwj/roZqND3VGGO2uBV46
kxjYjW3f3a217HI7ePF0gES40lvU/lfF2vyL3xTL0K1aA87ATVOa8hWkUrC8VEE/42tHsVCm+T4t
SRRIwHq5M7xjgKANKkVJYcYZtBLDPWXsX8lTGUAnukzbVAr6lWTjHw38FYhl7z6sCjAZlXH6H9qO
58dWVAJO6/6cCq8guK36aIcD9V0YwFqTVi3PbTdBRYfGDmGOowIhUSPfln1OCpucGOcVsxA6fnBM
tTT8yOBEz7qODtyDX28r4JHcptGodCE51MY218XclNwF0zTtCRMKvMWgPGOuwMD/+iWrzX99e3iJ
OvsnsgA/v9MPNATlu7wGO+TXWSTDdcqSGoRd0oQyRirSuG7L+SGdNJ11q0J2L79KA65HyTzLiwX5
kSJUV+7I8SYfGknj75HnfGKddhiCKClXKO9a//mcVl0SOJIrL+FvR+Kgt022uVnpUpzL1k57A5UU
w2gvmMNMcxi/KkwxON4jmFBn6fxPIyedsa4kevkTHMZ0EzPSvr5c8bLFL+WjfUHJK+KlMJAAjIt+
6QA3lMCoI8QDT4FnHb66ticbWdusdeCUwPtoirAISFlSP+cCXerTSGQE7TA9oMBKCDLsZ48iz+RV
5XFe0RIZf2JIb0cESMWzzHfnJj55UrIOsp3qxQowawJ4r7Zg8ZDD4SRq5/cLPitt5KALzwkA5ZQu
4sR3qg2Ute7AKBc6/uotNKy8lvmiAGx/bl1hN98vO4xkOsRlRwKf0z932X4dwCfavNVrlEk5e5rD
QsHpSZg7Sv+xS6wsOlkEytlbhoR3U0QHcViWVJUxEqXmACaZBGOmkUBZEZKrEKeYdEuvXNtaIcFM
df9WLqOrjODwrrR/5VlYOtyKWGEDFW0hmH/pfZrdWlnmOEHuW1ygdtf+7fScxB5zCLwUdv+3CelV
mfsSqucy3h+znyUVYTRafwdWgaR1oQsMRe5/zSrG0jt3v0Uni+EaClYyENKzs7leMc11sprn27Vb
OIaO6ld7odZrqboIletDJeCPABseMdYfeibqPtp99l2pS6lK6gVlZT9Ens1fdPjgx935FgLLPO+g
BzVZXswW/ceOxbp/syIHaelsAhKS3AQvO5amcaLvQrPIOFME5/qSNDLuJpTJt3G9jh3XJprcAuaB
U8noZs3UBO3H9B0xEq448c9l+DzkNZqzirtSfvOQlzcOyosdRJ9xdqzkfcGo0xvisCJ8iQt80Zz9
IR2bZqylkpDHw/5LT2Psb6TBMPCJCHCvPs6wWLB/Aazh5rLvf+yx1GmWjbb6kknaekXM2rpdVTH3
j3/eLd5mtJhim7twjCFdt0eCrcTZ6GM3mj0dODYXxrzVBHRGIM/Kx+bhkcozaP3Bf7shcXy0WtaC
Ft6mAHIWiDKdDpr1df/Cqd5wgXBVmx6IVIDVvpXjdSfe7mVpvgri4g9qq3JKXJRp8BYORGpyBdUf
dDBotyg09rT/rC131Vg58qLpR1ckI4Ee3mPNCAdv0pG7TcZLrEE9gNYTVRGUdC+jeGnJEm4yUaV4
5QFk3N8f33vOBtjXqSicE66qjzoqWGB96ovJ/My+0HhAg53XW0N98x0QV1qzyQFzffsKCaBAMnTK
5E/jwCeI6OmkYb4tgttwzEuNk2pO/0+gup7zXzrwuEAvtUPMHLflYA2eGi/4Qg4ChOJQK2z7Qmv7
Dv0CmCx8kvkZQpRLnfAG2tUJeC9VN//h0kE3PGY2BkyO4NZtTtpmiMeYfJHwB5sLuH7wMfAIc6wq
iN8+IqXM8+sMKr5+nRM+R6ad9bnC8zOsz+kFVfOSnRg=
`protect end_protected

