

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Zt+Kvzwu2Ua/vrjhNueC6ZHFBDEZvqw7CYHtLwQCcRpSvR8qcFedNcWPERpPju3eJt3nf1a3JFkv
PrBPNZe2dg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BgYona2Iv/0k72I3J2JPeYuzuEtaXjhj+ZWCoU9nVssKXxrxRKdrDHt5tFvberHeN9tDv53k+E0+
zSJEc8s7HUTXqNlaEROAMDRbOb7ChasXXdVxfl3WOvXTlUGfsx+NSKJ4/HfkR4Zaiz3A3zH3MCLl
LSzFeWSNT1Mt1+XG8HU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FzDw40mQxR9kpm1uxLfUoItwH6249dxMvWlSzzE19zJKjsyLJvf8oLgoShFkGPrtSiP79qKNxcUe
hzH0hyrZBcM+hC6bI6Mi60dC4BhdqclOgz1qMMvUNpZqrzZ5JB+kSMGHVFW8GUXvnFCCxYuu5mP/
ywkJGUeSDVEZY2th7ObJJlKEA7icdJ5tzO8g4W6w2f+MHJPOeHFy+SupHzB+1djuSlirLlm4nhaI
hraNZ0zRKoeVe6z0EIEqhB9JNsFNiC91BziwCnpzBdkOsKtsrb3RxMWbRRWbmc0XLssKg5Ki5yKr
zZaZTZk48RIng0NJRYTCGlINVIuaWueM3WuBUQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gVm/uXv2qQX1H4bUmXuUswxUb0GUskWeA1MPfdTQVCi9Xt+VdX6mOhlgO6EFKXSas+dhLpimNzTK
aBHFEULIiJVFga1QEdJchUQ/rBMO2ShyfVm62wP8vvP25+deZ0Ac63uVlMRNhE68fori8KTc3x2X
Z6Nr7gpu2y0w16PhA7E=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UyIHMrvI7wZyM6hLJ4gE4jKiSWW2iEuHADz2BcA+kHWTu+vXmBlODWfGdNNdgy52INFMV1nxlqnJ
XDvv73yssq80S34n064XoTXJBVIQ+OApIu1S7Z1OlLjdyiOtUW3Rq9q1U3A+hwbuiZ1x4LA5dZoj
5xr1PfS7YeIFNi86pALVL/xngSOmrya7h0pb27Yqn1ZWp+ZFU4zxAnMBdh6smb7IVFLN7MVgfSOU
BFsRwVHyMW6sC4c5q5LyBHJsVE7Cty+4Vqow0WWDEITa8OtbnNcM2JZrP1+VHJVzH4AYNHP/h5/v
rWvTg/dH3ZrlceYDFRqzQnHfQLNZHJkGerETEw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 42448)
`protect data_block
DhwJFVEv7I5AMXt7Vr9cFA1nWzXzGdcPJCl+OWeZNPNsJe0ny2H5x/ohb4VK8Rto9QITp02yM8Ym
DSiCIshndWlHGqUyVFQJr5DHXteiP3Oj1b1OPfyo2kDIC8tbNMMvkttgM+50eFs4K3CfBRShk3Sn
AI79G2N9v2441GXTeHT+jl1iP546GLPaAKmVoDCrqxcuGHZD5K4bL9fzZFiAXEyS6oHDVdkFxMKy
lqHm7AjvZ1w7eEpHUXS2wFJAX8xPICRIJS8wQtjrAuXde7VjpSlOmVA7rfi77XWozMRz8XesD4cv
oMemQAgBgIzkv2MZihds3u+I9iU02npBKvaXQApTkbvrOCMy8oCSjea0fTXPMGReRFdnD3Xh6lEY
6VnhPh0l3GSfNcd7M08cXbWVaj58KaQTzduTCYwUrzxNfvIAFOU/kKnRLmNLuWl2QupDr6JjUfrg
mMK8/VZrb2CdFF/U7SuuRuvREi4MuVSEBObDTOdeODg2CffJpaPUACdX4rWAXyMtPoQa+Ryljxmm
R2aHYSVMDWofyN7UJFH9WTuESY1wO2j31hPk1NB8BpzuB5dSCZBa0L52nJbzZPB3NNqcrk9vbVjm
ZdpVuiOCGn3kEWCfFxs/ndjX1io5C0opA26oVDSdR8aABQnDGb8++E4apFTZUFI2+iAE5Y8rDsbX
mZ95T+Oa8S/7a5Ola0L60j3gLof2EZq5ReP6A6uroeVEUzmGrDntB34c+utTwhLrHKP7DR0hl7H0
hWOh1KDRxQ553KPPy93jlSvvbEUWSl3o/aD6cZPROjn6My1Fw8oHejD/jYXZg02Tr2qfP1V09ZkS
wp0YE+Y0bIowhurZSM7tBdZ0j32GdnJK2+xZduWtjLFhgndZs5D/CrFS2ge6Dwdg167MNsfUAJsu
H2zDtoUUBL0KQZ6RhlF33LOpiU7+JjZhKc/JB98EG3w/SkdHrTtl1kVeecSaP4RdVRZ6K5i0+9ED
oqFlZdEiXhVyGZvaIVUG8fQ6UgBgP7E36MLA8vSxKWTH4hDG88ei/kKuJ9EhyouCL5ggPZVj3646
VHmQBMs/wV5j75OvvZrbC4zLhDFTVPlnYGplGO/q4Y1FhjuvscDRx1s6HSewqacBaSfHEFpVSVzd
a3pem4Sa6RqFIur+dWjmEEA2ZUUA6vOF2QN3Nbfr1RXWhJd65gqpWFnlTPXDpamhdSVbmHtF5mtH
xKGv17IaMEFZqob3J+3E6fEBrj5OFT4XoRoDXLoEzdraJfVn09kOkz4nNc3vs11q9zgGX3bfQPpy
uI0SRs1O9o+KeeveFe32zAgLDjDw4E6ZIWZDkbsirmqmkBHtxUawYgeqQPzj4iW34i1TcgTxt4+d
JTwl7G1k1JVDAc0YIsM+M0YP6YTJHGDxbVvuXjed22GfL+tYRM1LmsePBSO520zXUcEn9GEMhfya
0rdam5eOmVXhDNr/s9fOkAPoeLfaKcvwkyy3DCD7AeDXinKYSCIZQAVfdpYon7O71tzhN473uGS0
TFrYXcZpR3VyZ/o7tSf8mZpkeaSmkLElCiBIGXOkXcnoaCpJxj0p3JwOVU1kDlOwxuvetzDVU+pV
CSPTtUOpR9Q2dLUBcIo1XP4B5m7sSN+zDuYVTQ5bkSLBh3cpqAcmutmQHBMih12opooz5zTzMDkr
LYDHaY7EAfQp4/GqgfhHWb01yeJoBtu6vfueio5zSrKXygq6zlT5xQbEzuKQiaPzw3wBjGfMNlSz
n56RMoOTQruuav1QK9Cat10fTnZvMS2EThI7jnqN2ifw0YkYb9FtYIY9Z2TmB+X0B2MRberQjy0G
krBev+K59gB6MmEGOE7LfTc6GZS7fAP14gGwlw1/9xSttCHp0Pu/APdyxvkwzMnBsQPZDZVQ9KpM
FQ6H8HtZxYs/TL+TQ8PepPi3WN5wcdeGgnS6Sf0grXXl+esvnnKNnnI8VamPlfPyqoVK6hXPlLXZ
iRNISa2Y9Kb5zROtq8DA0olYONYc49efwtip2nuUMn7ntJH+GdIP5aoVxukM/4zxFbcdaRg3QfcS
uaANJOifFyutSHQZCAUvvGauntHkAqyVJije6uZ73B0ImZI6D4pDe2Klzyqlz05T92JPMk8jPHf/
iNUCK1BzjPs3VqCQJ31UGW6nrgj9FgFZjlcEqvGz4afVuc2kUVxTDc/JYStRoWmssX37/+xcPIFU
qOpSOoDuCoZ/DYOXbwTO5uJy32i8P3gRbtR+Tx4sk/5JMzWs5ARwhMyMhK2S1kjbkFo/kBKH1PLk
q5sZAw1x8MzY6TrUcrMaf/NL5XJGEWaOKBzDb/IfPpvmmNP7aeOCqWdZVLg0T3W91I1ERsT3Amhp
nJ0+nVvVcnpnHiahHLcTzgKyDmn1kmi8De8ObcFv5yep6x3EkUK+vtrhwfK6UDpnJUkc3trYHo6L
86RR0oXeqVqy/RfX2UqV6YYHclxXG8OyVDdiy6saDCwxahfeUbSR0bF4PiKGZhsPS4SFf/jDeufL
JN/9V+5W1KlRnctNZ9R2nx7P3WqZ2NhSwM4LOquD5q2cLX5wfPlM2LXQDHwXOGUPwIu8RrjD5Zn2
a48fJLipQl9KCqu8Rfp5hDEjvs9K14Nigd55p4Dc3l5Zx308dmvQ0RRB0WJAQwV/SE9FvcmXMDV/
tMGEnxACE6QQ8IWaCz7s635M+jc2A0X88WrMiJVO91CpnUDDElhrBcldHoQq91994rjMkT++U1DB
OY36wALgal5ZtJhFLpncjRG33cLryadcP/rVjZWCPC+kjiWxBrlYp0vEdJjjV4sFxyGAJanYI7zV
pd5/eUFRrbmIysFFf1w8kG6rZyjr+e0e+yTRjR1naom/OXEyIJxR/Dt3ka44GS810YXGVZ/b2+mT
9RKHK7h+G6bzBzjj43S5PmR2GBmH3p+YgSAGoFF7o0M/DNfrvsH0C99WwA1BF1QGO0iBo6Pp4OW2
XIE5/wuziWnfkO+f15f14nsuwfoxCip9fDTFFEJlU7qOG5eo072/q453Jt3P0HYCvpyWHm+t7xZT
cZq2xo4kyQI3aBy/KAeoUfc8GusWOiEYn19p8np8wb2tqBSYNtfQBLOgMJ2wp8fyY/1E92ZMIDYm
b4j14koHtSTy5KAw3VZEz8wJjaPamdZHOMK3hAutedm5NIhnh4u1aA145Mc3LjMhVy/fP5w9oDXT
W7KSlxN1+FfJ25p8OVC+E634PEai78BXt9erQSdgZsWEs/mTP8uvjJbl5UVnkn/atlGDZfSxL2lx
TzGGRMFscJiF4UY/BCsJgZugQm6eW0j+nrFrLJLe7xHhfs1RY4TDG3+MecaDtodid1xLFosG2ZEp
ve1z0B93Lkcq0XIfBo71rOIHGKwIcqjR+i0e4bhYdh8HQewtIPLakNA5Dgx/eBaFfklB5UpyPzHJ
5V/0g6bQiiZO0X/WWw2Ho1NNU9JYXuzkYRYdYubUZ5z2fRPDe9yblqflwzvdOyezPbpP3zFlpf/x
1PDYNUoVQslYb1sn3W+0p2uZ0Esgjb2NEKAzkosHGzk01O8Qj1bhANyLJlViC1+72vczE+c7nJXf
QCU009fF5Gb2PQ8QnNsAW+gKvSPdJZbMh8leel97ajNyegYyr4z1ibZmssW2x57DctjVT3DBMIeM
4QQTelmkyT3c4qyprxCzNivD1C1/0xDccLcTYxrWcJixMTjwoH4yDafNA1C4GinZEfu3M+2qFO0O
+ane/sVSjek7/gzYn8KSi5Du9xVLETxmV278O60tnqcGrmsPj2iZI59zb6iYjU/VSXBqbEmqHDp2
JOMWKcA+sm0dv75h32OAVz7tDOd31zFHSUwZPRZ5iDqn/IluRKVGf++eK+8Sy3lARG0WyLjirGqZ
7LdkiuDiDes5qD20oeECEr0UEZu3IPa9dxQfwQ2IfRbozmkXsQMsp3qnab9E9P8QV+j3Jcjepo2V
9osNiHRjHw+DZw02nC2mzOIUqWClXmqwVtE/nWLwgoJCAOOqA1EOdWIrODO3YuwXm+w97rrGyHj1
jKIxkwJQA5QRoAXuWC0d9NyccIoJzEcP1SyFVQW0bTsfno/jjQZvaVtZ+OywveZBOSYlqbTrVsNI
QP8g4sG2o6H60mS7dCTKZIat8ffMT9WoR/BUqrzRDYsK4aM5WyjpYDXzVNhGOrRGWBLbJRV71d7v
N91RWvzFLSPKLsmS4eGdG+H1xRNrh4lFfv7FCXMoHlX0zElenz6gTdSCuBfPWI3rGOjDnhtQQljh
AiSJqrsqIAZi/lP6O0idGPJjCKgAVybsTvg5I61Aeo3nNKQVVjxN5a+PRtcpLaeI+LWUozlKujHg
gOJmk8NacWovuvv2oepnZozB0De1Yo9nOEy8nfefkkHsnaZh7kNkdnATgBaE0aEBtESiAbTjc7R1
rbbZzMtxxGe+OPAHA036TOX3/u2Hxjbq+YZlWwOphA4TUYbczckCBGaKPL2RkOZi3jJas/jAJ9MW
U9LlhcKMxyKsrq5rHTMVTRXARk9mmatw33lSL39V0QujXkD2KlM1zR++a+2kxvDzNE1Hlq0C3ugJ
nlODzKe+Jf+0zzw9esM4b8UuiYqtf8RiOi19ANmeYrGFT2Y5oqf/+e5mP6oMczVm+Efn7nN8Gku4
U7z5N6bLkP/EN+hVYrxa6/mUL0mN9UdDBd+cBZLEtz5dBgL4Zhm4DmXCdTnl0ncYzyHrqhi40drR
Y88mZchPlNL5Vv/md15d0XhHVrpzFNU9mB5R5rykBjWc7r9wmSiVmSqIAho6g94qUj7UpBt1YCDj
5QxIKpJ4JQbDQ902JnVUWtgfb+0xex2uzE7M6REJHtRp9yGzMkl/gK0eHtx14vZLNKY2N2yEU8bl
x7G4blN7NGAiTM716e3N9oxWt7j8dnPlyCOvxj5lywvux1oNxL4BhFcpgxM7CThr2Xee7unY1p03
PE7+6vdPn6Of8O0Z7XYq9s85udhrUQlajoSvOayfqNpAYrs+VxOqoqr8BZ+yqu70cF8aRFrDVNlK
YOF/+Cbx2O7YOi8qP4pIP9NyD6q2axoX3siYdfeGFS7tg/dGqgzCDP5xEet5teMk+YPFiZvVUyGv
8m5ppZBDCh1XqSNOTjlYhz9wjI9ilLz6/6AqP0C1xZ9zoO21l+IzSSapSl5xROmPXHMIqi00rabf
f9a5FxJmDAqmUhkqAS/U/gTeNwOz71nXV6RqI5rd3i/bMhMSM48IyrI66RTmS3eJJoIfQIBFqCS1
WM3Z/zM3lMWhD8wQxqCQeuEVyY5GUe+wd4qQvD3KDY6gVednEBD+y6zcPUDVDzh6dIvTBmieyvP4
C3jgFuimnVWoyMCBXgqPQVGuICARRSnoESDm9QM/kbuDeEDY/uEMnDTtFWl3QgarfGBc4uJCiRos
wt87ih8jrA5H63hqJJxv5qyBxTs8086vLgCLRE7+xImELBWhy7oDnzDtAwbD3saUEI+NTKrYVURx
Sc/U9DxkYLIZVthW70i37fXpPYYmKWQlLW1LS6wOp8VfpwKIHKkL0SekDLs/U6OWj6WvG/LVrirU
hUW+ei5v42pEJlN54evR0AKjl/8S84w2WPwSsuQMrp9VtWIHTlqiXY6gMFQBEdXSGM4KZYElBDiN
vUp9JtwrgH4cEyoLTZe8N+HwVPpBOuxjSCUw+O4idxRhPQjvt4QzK1aA6gqimPSjBHhOozCEb2Eq
Q1ZxSqvp4yejKOL+3pXavL0coPTCN67H9s/GqUsgwxvcleTFpKX9V7xNpZbNCgZQYR0CqYPKPuNm
GinN5pxg6cSuZZHYNFaCoq/f59c1mIaRv8IbXmGC2s9uJZk7DlO+x9wh3Q8JbFtTCzS9t20txDIy
FLjGr1UF3IoA5I8K3O6mTvwhBZRDZB1Q8Nm3yTMo/cBOWZRhRPULQUqVdmPVkaTzPr5odxtbOzxR
PgunMOqVwJu3NZGkyi/vAQbCEYvqr2kMdTmWFD6cz5UBLaZN2ngnhRtpsOmZjHiansP0HGT0jwnn
iZwIoadZXO93yvILx4dRg1crH8YwFzwNBviY3MEANyvT5Psc36JlhwKrPmrVguaYsL3uvFqjuwP2
6caTEEsf9VRaQ66NmkGMU6MQEJA0wExPU5zsWYRZzeWXSA8DwMu+LVFpTVZOygelzxzPHychSu5U
IzP2CvWcJucWIQNyOPUNl//aSPS4/8qMdqF8bdjuzehEmfgkepuaZ3HI2yBD+eKyU2HoG0+DLE9P
FMbhx6i9ye/txFE01+Bh0/l+2Q5biGFfT7bv1nDSsPDCW5uLxw5oE+U/pnNf2+HeK4DaGx4XINcX
YXCvIt27yVkiP/zYqaZ6QwuAZtU1eTRa1Cp0mavAH8xtZezHbA8d1uywJkjjDVYO+tLQlfqRFqOi
9OgOSQKSIgMsGq6t0/2hr7Ls+aug43zJZH4+mntxNxygA+VgpYuOiozr6HrUDw/P35IISXoiX0Jw
y+/f5oSKY9fQnXcrEIJemvwfJjW40KV2r/9jOuTQJxavb2+F21WVi/qvR97STBkgfWxNOucA+3h5
RXgzukHxjzCN4jBwn4Kh828J+EzC0a3HW70YWvH/01RAc26yP4T/feq73+HIYSOEy6/wKygsxOAh
ynW9Adyv/F4MgX6G+FYt9SDnpfudumqk+Icy/JDwQ0r297BhLu221wnZLFBPXkzkxfv0GDPf4n44
8zuzFdB98wyFbEO2XAvWv+Mv/i8FJ9DiAnjLPFBB+j4RjqPW5eLzJLH27rXp1EqFbjElx3uvDy5M
apDymuCMhco9c0HD26TP+Uip8TJFP/lXQMPeZzFR6lBsmFaXs6S/jJTSy1kR5i/Jro0kbMBaQx5G
MJlVo1Hhw4ZadxlJcgUIl/LtstAmARylVwripx9o8Ltw0fiLylYWBiVRCOwonWLpw2bpvD4DOyzh
SUYESZjBRHUBrZ04wTDMKWWjyNmGiG6qwadajRCkieaTkdpd4mB4npKV9KXOe15A22zLrPnbriGj
yzre7riqiwP61+gQBAhqPB9oLwXvXbV9F4YARSJph0Zfive18n9xIF5cDRbrhkPMqiiBJ9yBgK7e
Ab5dRCWP8e42E6cso3Dw9GZxR2ZhHvfrI6l0BYVcKy0FjD/1OXnKa0RFbu/PBIFFGwn/QhjnirIG
Zk+0bkxE3Yebxaf/4C3proxzpoQKPLnvQSBe8LGJ+mwoZDJTB4UocEBNdcpFhHIfpTmi5sF7Bubs
+0mVD91FGskDSAzCUoCmmgUEGQF6sovvSZdqBjUvRfs0E/7t3+CDSnWH5YLcypCXvXrlPSx7JfPC
HVwgHPB/9jk+Rsl47lgXtPTiY89jputks29DCWTi4e0gALtEuT1B3+1QZwJB4axrY89NgNHzaPLh
zXCQBGm1EWNYlVaQudQOnkRPgoDXF+5rwA/4TBglM5d7f00s8zGgaQ4myv4nDuCmUmVWIa+S9hmK
FIwgcmCqYPj7AmeIyQ9AW0xFo9sl3W3SLoKQeDrIvKHS61sCPnrrx8nY9zcbyvYinUSK5gh3b0jj
iG3iCsnDAIOB7RJyqHKpFvzvxzsHGapBTZ5gYY9M7z6A6W9ST4aPe0to5N4doMXzI5WrcFKCUWgW
5y2SgAd6HMug587MMLnH1S6MrFVg34RB/5lrVJ6o5kpYFwIOmyCKWY9QjnCF/EJu4qs2KkRO+3nB
dcs8+x8bnU21f7QwTGO7F0zR5RPn7nzvavjasGcY+PQOKpW7ICyowQo+RMk9bfEV44Bnk1OIIwZs
kz6J+nyeFHKqSQOj+fgKqmsqneu80xrG22mBH7DWoQGv9JtDiaxpohugtDf1WAjut4aFuq3iWdYC
0Rn8sfwumW5gqY5abecOew15kEESkKsFgcC0nOiWjslkpZ+BMxwkYWiJV2MDALR/TLZM2swYytU9
foDSbkoBp2hjX1aUTmy1+YYJmDSBSOaQTR3kEo4QZoEeCsXRjefilZmWM5M+gRMO6fgOywsUFeUr
YvaA+AJigW80nZjh2oik1zwXkW8zlN2KWT/NXt4iLo2JtVy0Vgt7GUPg+t5AmqZ1fFWb85ZxfB+9
aVC3tgRUxRhxoWT+qEz3K8YaHSCJDSIbJ76Gjf6GJw0xeRJS+oxoSzyOUJuKGOxr6Dg/Vd5K1xbS
YOo0tApGCZNVImNWA18vWUYAjroqIJgKXluE69rhK5bWbDClvl8ikZmDgpPyO/KGuaUr/fwDQznN
yJCHxOY55V/lARHwbJqRTuxTu866IEus1FYRHP4cVHJqfMylk+L0MxDDQF1eZyZN5mW37JFlNHkJ
R7PSUF4dpnXIY+dXoHs142/mtNHEEjYYJUwMF4hCPMWUGVZJE+yHNoQzup5cRtqzsVqc/EMxyjWd
XkxPJeZNu06igTOTzw5MliL7hbZqBVp0ilqVuA46tMzdTyGvLeHG1KScwcbZDQXuw1LLYTxdSajh
9xYTRzxGs2rw8TlRJ+/plkql99i91tw4AoieHQRo1pH6iOe5VyYlRbTHbfIeDlaOfPjsIreiBTeW
tAHBnoyQlg7cuYalAkaBi+lMExQg70kCy7SSIrk5xgiVU2Hz7e4FJyfpV26ksZw4KKlarp30sVKU
1MdJV7tSx+S442DDlix3LA921RySSkyLoRVZPXLHEfen0zULPips9ntaJ63DaBo9P67pvl0vEmxS
yflMAPAV9nKS9peq3FxyaGtzA9SFXoMczlJs0KkIyi/bfaX+7OvKYrf76JQ+ffGCuGdR2GPfvQZe
ds9z0zFrgzpgRVAXl0bqagJhkFDmzirNxG4Y4MD3TMDbAPUtpmnIpYGHo4W7VvaYBD1fiBdtLXDY
mtWDR1+VJucppFxacmUbPiZg3URPakiYKYclWUH3tKkxkSoBRmb0B3RGbvxqk7uyTmi+Zx2S/7XR
k8toJQfC8LLSphCCUqgRb2170i/0/URto6Znp5ulI5ATjeZV5E+G8W+SHESBwNa2mG6zxpFaKeKg
Z9WcWb6HCHqtHV1hKEubQq2/A8se6ZeIfmiAPiNG2R9IszLKXDEdvKmUNANznZigrjXvjjTIBh8d
PHyXESFkcdl+sO5EKr9bKQFitjddM44gBwr/EkxH1XR+ETYbF6swi+yLOvPzljDM347zAyORl3az
2htDbcHAPi4iZqoo9ZVKm55OSMg+Mrf9Fwr5yhVNhbnZTj47W4MHw579MRgY00HYfXjcShrvdYQr
88FYSTMQunp6dfGGkMkz8/+CPU0N3FczUwmPnp3zyxfXdbvctVF7YrVdbcK4imyp2SGXueqvkId7
RanIEkAswW33yz2nt8iK8oKceRgv6aocZha42BR+emONMzQ+LhrnrwcWap+ssIEU/FnVxVJopo3i
CqCgl7ZrOxw3mpO446X8T/uLtkhqqM0M4FIFFoOWo4GM820ddu+h8ZS02OKsM6wdzbvNoMafr/2s
Nt8Nj7NbHas+s5bG3q3Hp2wLGNu9rwyHgdTmdYFfTF3igA5FW4RY9Gsj7oN0kpCWftpimPpeIA2/
qCwbz29kv8Y1NMwfOQXc8IJW/wKvWZgW4xd40eyjEb4TFQaoutl9Wu5z+QGMpAjpRcNLpb3w6UpI
Hsugk513RdXD8wYAx1v77rmfN3nNKMbgMroyk29Fs697zO9GDbXKA2a/EXVD0L03lR9AbZPcGo3D
4qTJct02T7o15riBRrBO1cEhG+aRNdvVOrXpCZuOlJKZOkTqYvp//1WhtI0j29eD+3du1oWZa/yN
Jvpu1huJVhoEWK/XvpT6wZcOxyXBsKAkqNqCb45Z0KpWcmZu8ejEFBQkjoY9Pgkp9SQLLsFxxN4D
JdjltGm51JfvXCSFlyA7i1F5e2Rynx8W+O5i6LnGA0lFForkX7aqU6rsOs8ZfHtr1YtBk1ep7t0Y
igYGdETVkI0Hh1MTl+E2RjjhnKax9oH88qBrS7FbR4B0Il72Asqvpig+ZR/9TrimzmNscH8Irvs2
aM1QHGhrhQgBxbT5F7m44VXAFmdr4Om5Z6lP6nzF6RLrFMeRGi1TI8Q5m0+4l4SEt7olptDT2+Ez
PFMgT62T82gjwm05Z4+7xXKJxSVmgaS6v1R8Pg+78fzjJQj3t8Bd9h1hBASIxVAkUCLUJZf7HmWZ
XAxdH103V9ccQ48UBpj6/1DcXkYGzDTtvSt++BXPjINJGx17CexfTKHAhT49QgQeznWFOLgrIhSl
ZcnO1V9QB62CgMJeYSCjRhgwiLcdYNJhB8seArpN/EH6uMpRA4I9bdrpRKfasmuh3/bJUxg3cPv7
6Wn80XSsR088yi/wfOSizO+VWa1KfshgQojPTjImrY/jDYj9++WDiakvrvT3q/7f8H2bS2HbyPNg
kT/xxN8VB/BTCn1MqLA/T4Cg4fMlHdycGEDiCIbWHHxLrrAgIgdbu6dBLDdCsMNUDM2DUSGwBAnS
7z/eXcjkYnHGqdumot1bYR+Xw2ot6FNlTap1e3vO6QWRy5F3kIwUArKhdtgfZwPFv++wkJyy6dtq
k/FYh1MAJ+Zpqy9iIeAn42/U45Hw94WmfzWeW9D1pA/LQcQUbtLzFhcOU7RLsaCitFSf+vklppTj
wMZYaaN2reN45sjKvjPMHr3ggujQy23W0CazJqi6L7OlyWIpGWTX4c48+0dNzBSLe4ievsP66Faq
GpSoSOj4AssDEXenzW19YHBlGiB9naRNsGr8qbOV55csM5fkOSSCEo29zfivPon86HTq+5MFRKeZ
vARTgVKK3iU5NNdF0fuTeHC7KI4u+2lSjNZnM1LBeOp4GTrBMM+j0lBoQTxLeu6tgt+kaVA08uci
tw5hRjlqP6+BvOLQUuBXTe2c0EAS0EosqIl4gAg1Sd4aSgOXNFU0+BDNs3Rv35dCy/WuB8xVhTi3
IhR5gse3q8/RXCx273U7DDYVf7R4kQlMZ3wSv8AILYGnKodB9sktILK6TNQ3k3q1pN2AI5s0ms7U
cBTEQQixvhRNX4+/3pWeTu0IfFOl70yGBptK2lYDrvOqXGoJjI2dlbw3qY8UUbMzaNHIG3grkBfK
4a5ckhr5nVBbQycIam94UNBCAW6LjcjeUskzVoXf0Zqwsbf2G2tswC+Px9SrE+Z1VSnoViR4TE0c
6DLdT5iEy+XkSNiXgaTbFi+PgQjedX9VkbK/TxkzqPDw1hoG8k1DVvgV86DcxTff3LSdBAy4HR+x
KHIXbHlOffHecK/m+3ZZ8YENZX6QkVEoy243NtKDEk1YVuot7hqhJdQHjcX1sLagqDSCg49n8giQ
tYZKn6rpLUzxCnoFW6DAIMvMnjTGxS14vfK3zuF1GQ8vDKirPYSeZA+uAi2IPTD/1xIGmhfCCUYY
5epuNzvWxVUTh0dJgTBQLqcJOd1ymApHegk3Pq64bpTUEUMCNRhLzmUmfXCjF1sfPEBzDqAXf3G1
UZSg89oq0sAxLBXJRMOoX/VH8l63UEKw0zqsgenNmnxT2keR6yP+qH9lCWgBHpiuQxOnUAi+qQPS
/wwODATh1Eyco3hlIQy9BH2ZQomYVT+A6NFblrzEdibeyuWTyd+EyF51ExIUEZnaMcYyqIsCjKb6
bI9VtJRLYHdToDkbI94aWsk12JLOio8ZfGlDLfMsL4n1nPxRxF3Rlvue8V4avSKjryoCAQWlhiK2
1LK65yUxFBGtVNkxDut7Ke3BGnrQ7CmMZrY0MLSOTfsU6nNay3bWEM6LRwzkOj2Qw3hH0ogQwfrQ
3I0G2D77Z/mO7MGsPEyVFriPM1Xf+omjTi1W7q7iNNt3G0RYtyote30rNhcUvaVDWhOzxoDWTd03
6KPAoJEV4Iygnmr5uV0ATEZqkzgYLYQTJZ4wTdK51l/RHBDILwQrrJRIB50hh96XXWxA0jkJb4oZ
52WUQOMMa/W5WAElbvlNtS1iAX/31eYjEf88IogD16RL5+WvXbMBAjbd6X+FCmVK4faCRtVyKgSd
hCoYBhc7vbU5rvIcVd3MVpW3qBgcGWPzHPRVu34FfD1dFrw02mtq08tjF+YXh/i0eU+CxRh7QOQP
9Qar/LoNWunbgK4LLVT9HF8VAwFIJfxwAK/8WryRJK6esok4StJE5MX7R/+E4xnEwlrp8MvYH0pP
xAZpHiilSuTspz5uYyQN+aqaAo5as51sKGVcnoMGmAggqFgBOEQ7hJ2D/f+oC644oQtmeTNRfKbI
XMbb97f5hwjnb20WIWE8yaiR9X6+eETTORjlYJygR+ikRcsHD+b92ZNMNQgNscqFKaST89Jd9DUt
taTmVYU0PM8Tz/J5Um/3tHMM8S1fcguffZjHZVk4JQ3krg46gnJumO8wLCzHip7hU8c1Fz5M8p4t
JaSEuKMz8L/dTbRqdCoor/bJbGQnx7IPl60DEB3YvFzTwvXoX+kI+G0iCB16Hpjrbuikz7MAr2ue
EGLOSm9q28tW1mar7QPJ4whfAmblhdm+4URLFsT9tSJGrJUe6P3w1h5HFk3ko/Bk/lp93sX/s1Qk
/7AwfMKpCs3g3/7zmcj1gUxf7BB0Htd6lcwH55ETxmMbVoKyyZ7wnfCM2dGF2gkjZfqj1kpAkkms
XzQgKMHl8gUUIetZw+/2FpU9uVMxBhzVn90eGxlKC2Rc+KrWmglQkaDbif1Aolc0OjlIbw8sQeFV
3bm0nqycUNPaa226rr/AwO0kvO87mkq+wtj6xp2lYNTly3Qtz7oA2BL9XxKRKuBg2sQ6Hjg5MFei
kIPLpkMSMsGmeI2Zlyp0M+1qsUJFrJE3xg0UDVDwU4T/EZEefayc8UUQ0beeolsbPQvI+ebNQUqY
aofUN5ctksWQq8HlYGIVOBWXUShivITbiD+WXYHMlcnK37L73q88FHJG4PHtWzMccYvMZ4Nn/lGj
pKSh1cBTcOLVBz0ZOUGK11+ft+OQDnquhrkyfPAoUvTJzJHOqHxqug0As6rZgFf1LpOpxScT2kOH
uAZ98GS+v5cHngvbH1gVkz/bwODLs5+0T9ke06H2/5ZyS4UpYk1pbApR3xl9gUCSG5IpHDtLbabt
QjvArmsZRtzjXwpt8Rc3jnR2EClTgPB6aMXyzINckXdK3Ja9kQhw7PoH8/PO5uUg9wG1SFGWd/VD
t11FJl9iJTGbuCZjnFgj9WsD7LAj6gvD91pHYVVJEj4ums/DnM6N0Ik45OnrmSH0bfAWY0HURv+c
li67ldRuYVuzWOi/NRLZAT7xGmx5Osh/IqJ7BAphFSsxJ/AIfN4NQxGwXbtdxDTDAf8/tasJXELe
ba11mZYC6oAThZWyMoOTlMtCnAmSML14ylouyWx+RHAi0OY41BvCVHC2p+ZPl3Yp4KfCX/3JCnvr
NbJZzhARhqIiN28Vw1Ln7Gdh5ejExUdNbXFCxY72k0oZNdMJDTaBJ9CDFZ/GP3uIDhLbfFH3iEg6
hbEDJIugBTfPR1RsjPDeCnBNjwmvRmEc/oisfrDGxca97pKByNbKQ6R7PJK4VtjoBOJrqRR6BYHi
13t4csTfZEDoJyvLeOSRNU9UVF9wJ9FchtvRmrV9SsrEF1RvZUV4+XjgdM2QoihFMFnJnO+GtyEN
r6fcTi/WZyGyZ9zf/tJ00x2P6n8U2XR32bboCJt9Rono/l3gX5f5Tz8+xsi2FUGbCar5cSvIqIVJ
6u7t6//qYps6pUxO/7wbw/X15ztItTUDAcJEtNn+KIgxp4vPhKxQovAnNGcorP6fyDQOCaJmzK0d
B2RvsN1BVEzHwvWD8vv5uZqtzBRDI7a00dNCtZqRQ8TKe4rdqqbThX+irMl0GX514S+zR38oSFzk
+qDf32oWEB72sLtSs2UHqMtb+rHfEHtO27GoJPvUJIvxOqh9szQ4TIphx3JgPbEDAx2fgj1q9+IE
eHNqFSseSBfEYr/GpbMFSJwGNjuJT/TAot/1zVIqXhRlX6FIfViCVVzQr/NLUVZhbpZgAB3RLNFe
Gkp8GukgdpRxqcPCb8fnmX0Deg909CN9ZYNgjhVeZEnFmQn5O4j95U81Vj4VAMfixGSYMEWk09Bs
XD8XOZV62mHVxbGcC+AX4kGDuVZQ1wUFqO27A0m3jKycu3WiwrPHnZOneWN3abIjPmEklfmj5wfM
c7pxcsfH03+s8ugFMJG3qKXe+mHSUiq+Ff3kiL+mV968SyKPFPIRdh1ncIn7/E8rzzTVvwJQhxO5
AEWDrHpw/H4/RbFIhXzzHyxAdWm9axpDliBCl9N34N9VR6YjLCDTB8IVnF/yYPvfVq2v3RxO3r4G
tXqB0ODYR50gq8aDG0g5OqwdRJ7GrkEh12c7xbiVubtrNMm0L65PN7XaTAEglE3X1g1lSOF3ACbv
WSmbjAhH03CEuN3b77C5ecy6LRph40aUPc6zqDXbbTUsoi93co0HfdkGGVZz5GveaHIN0rzQr0Wq
mCtKfZVVCXVyrJdSimF4sUOSQ8e0ty2S7SGQvGjgFEOGXxWekpNERClhkObMH0GIqtR19olkFx7S
7WCWwpy1P3ELv4d7t/R9lGF5LDsw4jXBszlmSvjJHzfKFjlYocWDyWPagK2clA3mYo3e14OyDMLo
9ag2aXL+UmQJsExwMvaHo3qEybNGW/khFySAgKHfLRJMeuWSwT+wqObDr2B1MdJpi+DGpfwz8zFr
L0Vf59idfMqPpQ0PysewEn3LibCpwDI0XPjraG6V9kl0DZbsUrGkWWkuQna14+VZpuN6+X7dHYTn
Mg8uZ5TXhcTC0KsiJuErWj4P1rTKhhT0Hca8Nm3mC7vV8IXGDDZ8p3IBS6mgNvMUHPZVt1VZSCAH
eQ8iICKM8MrAMwXcQPi/4gMBuJtLnhI+PCFeOHQ1EXfM2yaC9TRZU5OLzOjjEAjHoTeDKAs743rb
eBHSBUZq9oVtpmVgQSaHOWk2CUievzW5nX+fqpduAOc1mD/1ypj6EKwGhJuvsvkVC118/1KlY9du
4/V9/I8JzlDOa9G5InyyY4N3rHhH9FMHbFfJ5HM//aqGfOTz2wbMFSbDcHDgINM/UMh5H6iXhDUg
6GKHR+Lt4yKGNYMlD75NB7qJBycSZ1riQ2kCuAz39YRAzheoGrDIXWposercSrrDraDMItHhH6cM
LVybbAG6HoUbeJh5npH5TvONV8gsVktrcWNsMTpD2/oXjwe6403xwJWbJ4+pPr30TadM0dKW7i+c
QXdQDn9gyNV6wFkcBjJnxhIz0T3CWAKCIhiPgtfypqG9ym8ZtDaJM6pGg/RRfJX9vb/3pwYnUk78
y8z/5SHzAMIVWfyQ1TrURF6HQ6rI6IJiUREcwgs13YCjebSfTknuGNOpxfj15DCbSAJdU/wPQfl8
utlfKA2j6jIfbd/k9Ml2KnhkIGlgWz7hyg6Gf3BTDTZVYv93ZKeNcEOkSWUzjpsJ1jvT0MaBhwk+
bUeXGr7QGdH7IplDfknfq5ovz4m9dVAfRmJxadZjAULKM8SvNSJb7tFkNQ3tyHBlzCwLnH4pZZNK
zJzuneHUTg8zF9Kxvx1Zyzps8TYrW80RVIFCOqIaoXqiZypIddLpE7EZwuZpPflw2wZaUkpwZNYK
LGog41ptOIC+pXK3lYKa6IrWjtNFx0oqirnKXew/Zrcz3gn0F9tgDxQ1ryotcqgR/5bCv14v03zs
n/E4YWMdDaYNe2rGuCpc7eIg8yyrQ+WCVyLWmCxVTxi3nV3Nn3a4wIts7Vhl91V7uN5Y9rGQVo5L
EfAIwDm16HpDVSL7cc8b/fsgzCDwPshVBHqnCwhO4H/UMaW/s5E9+EsWkW1tzOAI5DxpCmi7fdPb
LtPY6dAzXNrG5TibpHv9S3RdmzHTtSHq2nkhVo9ugZHhuAAYZJmH9vtuGNi9qubuuUEy1dxSidSG
K5A70fF3gXyTd+gC+LdmwtY41tr9B5vUZbHE0TMqlq/SE9P+dRcERKPV78TSgvjS5cZ9YcA/yoQm
HnzrkvKtNU6Z4zcl/2VrgvgQRWm6DUlR15DKCifNM6+bKQnQT6BvsN0T4dTYMb7Pk5Mk8QZfgPcx
eHb1tUX4eORbcAvgBmqsJdqKHsoGXoXBqJbnxNE22V423Sod6LLiN/e3AoRMMDAMCBWMCqs59TFf
7RtEvVV+3WiQ4yNvWI51I+TbmQHBrry3hh7elz8Wovoq/Kfusis1uvRcgwyp2xU+PTShbrTRlHhK
bK7igGr/Tu46KQ/BquHO6y78t8pKTRmAZsKW8aJ+UXb5r4pR4wRdBgjYT8ai63d+JpcZt1fMMQUw
kHrtNO5NlZPTB03tuw4Y+yL1ly/Ae0iIaLkRAUPCydXPIJ0H9c3xeNutFcJHabdgkh0kYag2AbDW
umoApV5gOBqTvAieonbYHBv4dNNOagVUm8ql7yWaH7ZiEfGfd8zlMzE9fXm4l36/BdFpeGVkOPyx
ak+SwLfzSS3m501nvMoui8J80PxTQkxRNZV4G2DS+Xg5q+fTYPBGZJVfoRuhLPdYN/oqpd3gCKaW
1qoiL77tt+A3HeCemZLybqeMqwPJw/D15ziCzR4MkWMP29CiNVuBA0zd63LhTPw4Mcish89i6ARk
6o4myttNCuS2QyTt351yl84/Gp1qLyYwujbfWlN2hCVbZtyGf2vwVFnaGxgGkdIYUld5rSpSbzjW
pTYwYOxdtB3x/WYfrsQ0Hm9RP00YBu73GTc5Fws5Wu6QcM0sEKoKIYZSWQhzyKq9c/MQrNfn5aPd
s0yYOG4PaQWR8Vhjpb55d6Pd7i3bTmJOJOWadZA3oPOgl23CW+aYkZeiscpwJBqcgtzI7WrFa18M
hwoIdonAdLkW7gtLNxMzQI9l3g5Z9nedbSCPHzpNnctWTB1JmDuq9MTf/9LXaCGQP58B3h93DxEv
065U6XairPm+JD/vxSNyWeHwlgaPfohqora7FLKgfJ7qPB7hgQXPsYMl6t06ODAUktSY6rRuU45L
+2w2Bw/MzIy6IfLWc3mj0jeIFO+27yJIfD11t4x4E+68l9HQpKuLhmy+DxPFw1Rovs6Yr7Hwz4AC
JguyxiG3grbOjPMoxZlEO6oUlf1GmXWhA7wz0wwYDscFYJmytfGw2vYrkoqFLFTwNQiBQwsFHo5F
qSNJu84f6fIlYMmAJjIimKOYXoZlizXrLsNnHXu4nsLLLhjRt4R7KV4BxBfd1w6W47S2MYChMnYk
658AIEA901kTNn0phNT4Ow0JKUNR+jOT8DFnJxE1AWrQTQt68twZUZmphtr+qxW265KqlV4w/1hL
sFlijZcNjC9dkl3qGHydU54QOkuLAPu4Y/RoliXhxSJ7RMaa0P9yb8NBf4zUYtWyQcrJhKQ+eWu0
vulH4mQa74Lr29Or3VOycJcsQ07BHI1xp6g2YcfURPoj+kerPxQITxcZXcSWPz9nzFIXWvhxTlB3
H6ih5Yo8OmkBGNxFXfUD2xmeH3QaQH4DjD3bl6QYQAkZNYQmW/ldF1+hJxnwYQ4lZ7PD0HYCxERT
z67SjwbOEWb+/7oUZc5a8DBWLZ9fmGBq9ebg9HhWKXetUrtDSofdPbsXHk5ggnxfdmfq6J/TdE76
UZhoQGbLqq0dqsMrHMta+cMoKAJJjEof8BEFG5mc4aX0h82GYeCJQvJoH+B67zcYwZGDsIg1cft8
Z3wwYzb5muA609h7PGS0+rce617GXepQdm3DOvVXmRCcR7oABP/zdOPUCq9KWqX0gAxjgCuSE7Jx
Rxz8JN69iBUs7PGWQXwYOFodkAS5xC5qQuQGkrBDeQbLzyfVEqY1z16CciPNhixAH6Av5byK/5cy
5vgNKEeZUvhjgaPGTivhwfJsP5CZzK/edujd6dAXjhcVTYyaKpZAHpwPHyJ4GQLJCif1UGYHS8Ba
ZdfHWuHUyCvSQyQxa8a2WTwNuimCTiAXXp23eLt/qXDRQvpiysmf2gOySuwQe9xFX83DJtQQXTZd
0xmBKmp1q6/s4JAfZe3xrPz0GKZA7ai4sQHRKr/M7ln+iT9zfJdTzQRe8b7kjXLHkz7TJ/H+n19y
le6HpQgXIrgI2SeIv7mCAEjDbq3O6G+tqmpCqzq11tL7QyBzaC9VtXf2c1vbqDz1/koOgWvyoJN3
Qqqz+l0j8nkg9LEWUUZy+qzNI0eZAmpAEbJGrBdGFj59lpwx+utgl0yjEZXYS+QzL5pIUzkNA/ol
e7IEZPkmC2g7tVzPt9+ILKEDtX7VXI73ProIZc9OSzJxZd+j34yI+YqiuGlYn/vcOB3ndNWUPDaI
u5L8xuHMKSSQsTri2DcDMTBsNdVdwOs2mRMTugRQ+dc2jjY3TjNPQZYigZ+6Kc4uc+UkGd/WfbLg
UydcvSd+8FXzilPaiMNztJDMJh3Ii3p628qT6CkzphQvYOKNb7fYV0I72JxtwbUkPoy3c/ROYU6/
5HpWIkRYVAIq47c7YcXsDyLnsb771xl/48k7f7vmSF9ZZwcvQKslin7WCNKyq/bBV6CE4824HbLQ
rC4UbJY1QgX7zOAfRn+3a0ZnwtnIyhl5PpQMc/Z9Vp0/aiuEM6VZJyzfG5l8aAa3+YMtvwVV/jK7
cL/cvigYsOJeOed3e0x2OL5Wd32UdFjvYyxq9QCLrJpTJxICfMkLh+jhcOrA/jdWDeH7d37daHl4
vD3PJmvDX/3xd9z/forFEvOHbT+qXuP5l2x+QKBzBJ5aAw366uG9/8SOvAymL6VKXL2b46Pz+I7j
d5tz9S5vFM9bGoJ/btxkqELSfM5TReeo5byhQDWBJNTc7gSNDMA6cbLDoehbZSkeMLlPs6XqOn8P
sawAScNkTL5SMvMvNsXIlYsQwaJCRAradLuj1Ziq61t/VJmUcigO2yENt7wlQb7ucW6PgGYbS01X
EkLDLMfS+QDb8YQ0fGZGKktWDsh1I9Mh08+yFBkyahAASIclDj6ImijgE4BRYf229XDB8mvBZxeh
28OI5fORQcpSdViwB5wuF8yu2Kf+HIOsw2C34sOligRzp+4SDsO1OPd0DkhyLzmoQfQxBtBettbI
X5NQHUMRPnsXVbHt2vQ0kwj8O9PtQDoPVDDYgmC9fkpdQvHP7eSfg6K/PTppoK3je9i0B5oGjcvL
3vWgU1mtJ2YGyJ69cE5iDmMV/jyuTHUfxtF2xhOtNV8KKwdn3bKjt50lTegR7r2AevEz7pNaQKWz
+QuvN1OJXYeYEe7VsTLvN4qB+EFWwVEoBKViJ8CIoOqcw1GvsaIa4IRzEWGBsi+R5WegwSyVFt4F
E+nhoSzq+MURhU5GOQWP6OyRVIupzdgnEb1Z+sOXHXdVWZ8qrmhh6zMYIkRadClfE1Mc1/RiQqf/
BDFxS2zGkazltJfcLpyBbP8xj8rXvYcjR+RTt8zd2i3hUCONkyJiRP8tIGOCxFjk6Sf38h8AfeGX
PUzwkbJ85Rg6FE5nv1m4/OAIkLr3wsLEO+WL5JzCMGwArX1JBANQokOuYWt5rzKSE+m+f+RBJ+7F
1/mD/vwExXWilIP8Wtsu7289rQQU67YrYZC/Syfoa7peV22Yq7mWf0s53UgXCxLISGgTtPHRSd0k
pqrCavC5NMo9o2YD493s681wUIS+D8TJKWhiMdNltokaEOzlKuUWE2WvnefK9lZAMeuVdgIfEbwF
N0nm9VmAgGPRTzFy8Zfh6JGnC9RG1MjXaUr22/bbc20tCNcgH5lRHYbnAlQo0/Zze1HGEMr6HdyV
PQja10hBWhG5uXLzmnNirtopHwSTCXfZp8g9M8ttUArT/qU200LZiIS4sDvM6eoe4cK0TV3SRnwz
xtdgofcINh0KzR2/yFy0CuAULaxxYTkczx78auksbsOaqphMLYw5PYPjx5nEv/Oep+I1tN4xt9/6
VZxsTs1O2z1wZr5TRBvsZFwfU1lIVAlxR+oSOHASomt5ZnpvcCZRMHhKjJ7vg6ss2X2bNdZ8AV+8
b/hAnCiszKsF+YZTT7Fip91fCl1tr5C68TrzFRYoaH9uhMHjXh2lXaHVXJryQ+IZys9ozWoC4Vrn
d+M7IDobYSMCRSigTbBQOsJkSB0i7S+p654+Ifp+PTwm4M5k+2OMEEiCR77ThQ/klcKGMXjtr4rv
ibzWvYKD3/SSwJrDbIxQo3kkvmd02zZlqKvdkfWRx3FaaZ89mLyXZwkRhMbcaKNYJUTPB1CSuJMC
luQB6qqhZeYj4gW1x33QrfL5txT9gAel7yl2ae2T5wBbX8JCE6UvYB6KttmpQdqXyu9qLVGIrKc9
1SXvr8QvqdoHNwdGBBaTJuus7KqDZcTyc/E3Hd3NZ36hyst9+tivW1hblNFMqvRGBcDghySOdfPf
Gws+0XpWZ7LtpyJG6HE/E99bAKh+wtCePhr8RHm5enxDCt0TXA1iinLmoeC6ITRJoYeb07NWuZtG
KYZO+r1LCSDKscKuoLi6MTsF5yqc3YZBx9zcWJzo3DrdI1sleXo5vpuNaV5hjt7ycfy8NTjQit/T
qA1oi0azH90+GqxXNwyVhXlPyfH3E9jtXO83HY/2OG2n2g6LVqn1zLMjx1il7bTKbxDfNi4oA2AV
3XSUgtnP8bEplY3icy53p+rNWfZEEKp+EIAx2wJyn2OfgMeL0opkTDO59aCy5MbTnF7E2Un2NHVG
zafLIX+0//gkfzDyDvnvCzbc0X/XKLcS2uX40Prdh68yFZKUcn1moBEkaXjcm/nWtay+3seicddX
De32hGy2iJbQ8lpO+bbYfZBK77DF4rqGBz48UgogzvhOM5ExqMmJlOrfQE6Zb0GHKVX0OiiBmmC0
/jwAoczS9x0QDBSTyy+1iyZ9wMqp4CICwHSfA6sw2N4zf4kcYQX2lJZyeib5rjmgsaX/3toNN/ue
tJ9Kkw4zn7daUVrMMABquoyOaYLr/wjyIQV/KUi8aO2Cdn0PG27Y4Br0O4butBXbfox5FlrRT293
JAdbYmI1g74DiG+5VfqXsT3S2OK+EiEcfvrEvL8jxb70JEobwCxkJV593uIyUYQr93NMkk1pBzSX
DMXDSsZKZVZ7ORKbISJQsDozw6QHvNWuC2JikMacBSWc/yCjEy6AQJTzQoMQWCgqbzNSqnsZzAJh
i4dxuJfwEsebdEbeLIZg2v4EMOGLc0D6jHexfN9bgEFV+WY8pFG1FM4HZWdrcT+y4i4z4LvoWNDd
VVb2Mm9g3BPrtlXP3aVq4eeFGiwHu0oqV17BGqXIv9uW6hP0ZGCfoiRqxnKxJK9wMGFWW7ppNIDE
ITuOj7nq7GViD3IinIbuqdY0czGWgZQRwp/DLvYR95Ekz9yeMN3Sbst//lht0GbiQiNwgJoBvGpb
ZljsuUeEAW84gyAifsAGLRo5LuPfT2lviMA3nx68xIiAFH0dkCjyeBWa/wxrL96MrrLZxDkNInyg
ttVFKdNkM4+OOg8AjWUNXGbaK8tcO3VH8R/YGUVIC5QWImOHrp+xMbfDmkEu5LwNUsm+AW6rjP9h
76FZxb5W5LPLbWJuI4TUpxLWbIvs56+O4vL72maNExuv1S5jIMCrDnvXFfQXrZJFRYgdtpOeiS29
LSVoblooUjKLi9TktAkRwJwDtK/CPaK6XS87JXAlQvVGS5eS+JKNlx0v9yuBKBvy4Hz2jMUeGMVM
JtQoWlTnsxrGCvlfFJXwRawLsewnzwr8mjJb+3m8EV8X3FNXnWFCM1mck0Lu1KcWFYbNOLWfoaGm
/HPeBd5f4ztGCVMZ6TQn2MYyfuWa3YHhvcPrfDaYrj/2M1Bs5h4/Pus6fL3FQhSXz+EnB18VMcXx
5Nd1nfP5Z6jgENuijbXzzZHEl8Bnb8XSmgKmI52gdgBLI3XSVeM+01GuYdIEkss8r2NkLuefoPYD
emuBEsMDLmQgyiC9KyYfPwwM+Onrt8GFEzrKkFb+K41zkuSK2oRW4A4r3jr4Wl6hcD9QS7Awei3J
OeqwvYQ6rzQska6zA6VN3zDonsnr1tSp+Bog1BSZirFIyrXJY+/YR74S+8oscT9+Aw6VoLzbuTr+
cjLKIweb3MFmzazqPBwSvpjccq97o2+9mjv22VWZNdc9ocYLZNOZYmLtgLdX73PHD151pezuElpL
MvX5gMe7DywFKU4atPU2b7+Gp6xgfOtgu4+BIo2oQ7FKrLmcztbENcKTI1x9L4n7DOVLdqrEqwzo
MTjPeBx7Y9/yDTrpCf9vE5vMf52roM06QJDZymYQcyZF55tDy8xf+bcKNeruUNrOPSmb/VUqnTSM
iEphnvx6RxFcKHWXav5m3Smp6u/fuzUo5eHJG7sKt6GceM25DsHTfI/C7HAkS6hbaM9tU1+/MetV
sD1LMq+A6pRNePhwX7RbA8vgpvg01GaAm4cgXBLQ1ABIbqLikyUFZ9lFS+WJLr5SONXtQnAo+rS4
A3z2rZdHxFIdnVYnrYTFwGDLUJ2+9jcMA/Wh32aYmobVjKDnyAu6aYHB+WTkYEPg4Xx+iv5+P84q
bIOZj61O8DTcgrJwKmLfbprQl0aut+cRtz/ILpwbhJaUpUQrXnyL5byXRnOxPqfcVslbC/SORaI1
3iyKF9g5Gbg6tB3EyYWCfy0v6DIeHBZLmCoIiVasxy4e3VWEt+/I51+pNQX93BWZoqLnITitSP7y
lfBxo6ghIJ5IY+V17NVCbdUHMcUbTi1KudNys/6mHCpigSqs/rIk4famQ70/sELvpcRBoFcnl7Yc
21JOvDO1tqXw991R52QtR9bM65W3MtnZ9xBsBFHSS3b+m3v2kOY9RDH80jaS6CFFXEAIUWqURij5
vYLrn9qh1zqgrJZiF3wFnLUSuII2xbIXlrtm4ksmV/4zBGDHfWJ/a2/msg6jNwiqVLJQkAEKYdbq
fdi+Th9/Om+R6EyIV4St8EyzsJUk2qUtgEJXDVtZOzlvyE0SR0pveeoZNaSOZFJ+vFViiVG2kZXr
U1fSQWmRZlt76WtVwxGtt8gBnFLMiFLZe8NSNF5Ov02bonC1/Xx2U+DWDTnj+6QjnHOsBesytnuQ
F4w/vI8oJj/8dWP+vU6wdVFvYdLGVW/Wllhh6yKGBey1SBgmlxEhv06VgCWPeH7YkOSF1PXaenEg
VsL9Y6gMuCo/rWw3R5H9sj/hOH3x5ji9PxYpfuFfVFy13n+sojzRM0lhEGQAdesQVFTX4rIUWfHC
neYKxw8b4ywcJHpqVY+GxYCPrBODAQLjK5tld+m518XUgwlZh8UnZLnk0qfPmHkmnyvMvSOq9EAE
uq5VVJsbjPq6rpwrN9D4UVax02He0BRnCJ7bxEv2LiXbtvc6TTzacH6eyCXx+7xD5i0BlS6ori5j
FKx8a8LADu7Jaa2EQa2cK5etNsYfp+4oU67ELUtAzstIelUonVDFlQAcvZA81EDEnp92Uof4xU1r
B310lVNMCGnUnhCHlw+oZd77Un/I12YKx2ihESh0V+Uykq+rrUlkctRAaGRcvLHJCcZ0Zxsy0FXt
wrIGsJ8lDRbYXexBWMbKurNVKyOzimgRwEX9WJ0AnyNKaUCELX5apdYAZF5919wgkWzTXzSWWCb8
4g6Drf8JQZVYgp/BYlcqpeZiOCp9rh19gjHK3CUHQGG5JNfW3Huu9CjrDr7wqumTYmaPEe3nNlnR
Vv2mHZM6GUXcjEftfHP1uYVq+dt4vsWuIl9ElP8q/AqtfCFk5yJwLZjekhgShUoScI+dRPzNZgCJ
3p4KPFpZTNaAIUmH9amLLvCPGBil/KAfrMGdVv+gdjNgfZBRXiNsc915h+DfyMyyNdRfYJW9BtoS
u+d2gHeQUxOQd2xsZyK53oUiMKJj/yhj0+8ngf5/fe6LVLslRoVa7kpDOIOTCoSphTH7gVyEFK6s
GmjjSD8R3MLuml2OK8dqKAWogFQA8YWi1cJENuivS17ljOQYgxDbX+ufCNZrMiy9FRqOeHGx3anQ
iUawIK8wrpCEmpFqwTkqrGHaGFZgx565kiUkkcJXXGEbb2oeJDMTVCRDvP2SBfZ7KSOS2CbHOKK8
Yh60+brTX8fxEJK5jKbTvRnV/Z8kO5UvlT4sa7cIPc5wH4HTARaDvfZBPUhrumWQVun/bAmNb9lI
CTqEGYWC+h1+7mI+0sl1KgnDcfRxQaXA6bSkpFA+Q9u6T/9UjAtHaMizYEjNfRncTa+MazTGUCBh
UjO1eXEN697wQ80v5U4+XtRJwoo2bu0l6Z3C/Zmt7J210sINB5JVGQgx1G1qGb9Wp8Bpw9iCV7ce
TSgTqYRGGrEjO/141G9xeYf+RBahWbnknlKoIiZSiuh781lx/lJTJzWp+SkOrqlnhBRvZj1C3MEO
bTbEcCy+FgLkiJzfGJvIFfyvehfQYtU/dJn/2tMgw/eu5JEPYGssipJr66MjySHpW+bv3nssHmli
2blmP/8dpCqV3Wf7WUXCACEMDGlJtUy/OHJOCe2SIQ/QEof6EWdajWunwMBS3KaiAVjiqNo7gCa9
9NCORkAupQLSjpDjJCqdRQ0lwiHAF0YR6oEDQlV8gnk0lK8Ke1vq+jaq2g9fWNsTBYJ8DodLOfPp
5I4ki+OsIOggl2fzvrE4f9jj6F1ZQ+S47dNvaoNDvXw5HWXUorwPPTbB8XpVapcW9+kp0vGnRjRI
0JDx7p0HeV4dyyjVZbk7S66IGo8mmVLanHmXOQOpTF6Ar9FSlMHZmFJZ8zto3NykAYr02UV7jfMh
eWqbROH9IrZ+m0V5/Mbs6zm3xokmSjtgtP5a2xijQejBrcDCS6CRiNkqaGv5Icu+cY9hJQMaxllo
zWiaFTbDxNtHxOOoib3wK9HwphpR5vduU3e3pryUfUPtwhHvW3Jhjk3KVRJueYNnI5OcjPnbOW/6
61vanykwEVvb0UVkiyHFE0VvzYbCoj24ySrXu9+NZdhfaZZUseV51OZPczqQCGn7SNYUeeYMZ5UQ
6mf0fXLReNN5R7KtpVnZrT3IbDibXjaOHUs4ACLjNLje9mjkaIVMvKso9CeypmKI6P8QBW8r2hI5
Lxr36+nvtFeXhXb9Oz+1YRG4UCqA5kcGNTorAHYYb/cTpvpK6a+nb2qRu7Qlke/zbnX+7UcUkoxC
hQdGI6AdoGjgS15MUxMxmbOPbBhdETXk70mZrMVuUxKZH94MIDIOlO4OgXl4p5ZVQM6u+2CDvIXC
UNUxjM0BeokbkNXgmYC3tVPRajdvMjAYSe+3ePf3VgqGDQH2j5WPSVI1OuAnCjBh1Eh8mwCu8hYE
ZvsClbcuWbbLsRt7oZH1JrXLxoM6m0BsWEzcW3FLpXNy6rybbmgGEdekE3ZBs7KtRHsy02LrIeSb
LpE6V9wMkluxhJn+9owV4Zq+fH9OEuGqwYCqmzoprv2UdgiUDtRhUEfwwetrcVnFrwDBlZA+qTza
6AI9VSv29t3mtY+2H/mDPyDKEFAqgbYKJ4xsBVYbzWwkf8lkvEIUQ+/YRIwa4tO4iUh4L9OXioXy
BDlPn4LVkGxKar5ZoPKcX9LbbM6rtD05j+/ijl3X8pYKWpuoQA5YmWs/HHHbrW3fI9bdzwaXlq7D
F4I3ovGuUMJFW8caR22rLr73Beb20I4xiZfafHfV1ChgDhBZCumEfSISCsJ956zTt9/TIKRSNPVl
BJsu1OugDi36yAIX9OHusdc/RLo6ILZqH8JsORZyrouqqBNvRnvXz4vwRe5OVX7uFuCeaW+KhL8+
6HpejLin/gPmzmJ4Ts5s2lyr5MbF/olZ9sExVkYdPHRtGQ8D1iYnKGtK3Xi89z+mfmk5iQ3XKB1q
gf5QSUHF5O2SFMVdOVDTNkLdT9p/Zg1QWrXVEAjLlpHUQT40fIu22O6dtEH5NBwuvn2pCiRl3LOi
tk3Lak0wOLAoCYpjydBD1g3QIofGLr+QLt+7t6pfs/Co4SsFRFztbfc8CuDkblzk5zNdzdGjOdN/
NjpIDjGbggXt7Zn+coxaoKBEYpyVBjuksGe1DpKhQFF9uY1MqziHtfwPBMNoed9b1+CreBDmxo1t
f8os5JGmrcrK8eXAE8ZYeAiJUqFMt7oa4PXkU5/IHS76UzWwZeh9C2pkx93vtA5cpQxbOqEhLltj
OHCEA7aNCT0wt8Cyei9i2f7FRvN9pN6x1fYrLEDkksIAqgoOr3LQrTg56TatsV5iSt6D/I23BbSv
R4NPQZ86PKgOsSPpT/GXbcd357CSaUUaR8/UrUOgwcKUytBhZnB5DEDiLpv37UQJM2a6QrLQLfuQ
nkUxGjCyM6Rfe+Bm5RWLT2LyfoYAu8os0X6pPoCKXNiEiAo27R/qufDQBR4Hr2TL/52K4eUTvmUN
7tCA3fO43VW+InWRfPC00+5KT5lVqv9uRO/BJ1jm3iITi8kj+/2c5rPtB0SAeY2nTcpw6281LOsz
znkxHl5G6QCpN+gBfpgzq5ZBs/6gnZXsqN2CYDHRnfChN+OIz/9cEngWYK+rvkV35V2jAgUggstP
xkIOXgEKyi4e13ekkwk5jxBFeWuOk+KoviHsMIfAtKsgjgBkhoVknUPOt8ECcOOj7SOvYfvS0z4F
OfdQ2x38f4RdvWY03cUi+Hk3H06LVIUIE1kyjsPvVOtKhgo5wJhCkTwrF80mWq+I5X9qG+bizR7u
9qgb5BOI5R1sZBGR0cpcjL27kTSU1zmTfXz9i0a5cnF/Jo57u4dKJYMjfeOzLA0czHHeE76wfovM
3MW/iNzSP7wpn3+7SMd+PmEwE0zpFrINOgR3JhkYsgw7cOBhgPEa5WY+53Jw3eTXFWuJfk9DBEm7
2hb/zOwbNoj7kxt6nJ3mglTGKogLPL1CUZTAzMd/L0PxsjF0m1S58ixMQ6VTwYJJxAx6XYr3aH1n
CT4448ZQmUBPc/lGmkSOStqptQzeCbd6NgDLUyFRjA0lpFO4WyV8rJSXDI0zwxMnjuHXHtira8FQ
zcgTu8F5qU4rpvLTf3g22sXMeXAoTN9zVyAOqkEa5DU73UvAvtj0DLzwSD2s17LGxzt/fqMhAC0J
ELfABfz/J+XB874rz+uEk1aeg5L5WgJbcy3q3WuZvyF2dCDV91Rm45lGYpc/4lc2ucBnE63MCw8X
B8E9dYg7cgVuQjqQVOUlPUbWMsOd79adbtPsK83EAXxlKHAbuz/2FkRXah1C57UuxjTxy8FZYhRh
kPBgh2k1js6/0YWoWlPhLGbHKxVTfn9deKhs11lwaF92ecld0fcuW4n6TxPlQjrBgPC1Rq2mM0AM
cwz6PFGzYF+q1rLKNe0fmLm9NnvwG4OGgnpkeOFzizkylMU0l3RMHKgPvojYRow6g4PLm0ugIe6m
ncywWmpFKgPQIpzE8CfkVkMngN+XYOKjek8oIYWo17GSoXHKiO+0qPMiOdRaHvLM68fLplVsJ3kH
/B5roPuHq9fXKKAurvd0lvvx1hhwaMcHUq/Ot5B6824/A4KJM5NzVEZZk6xmsKMfBytEWTwIZXE3
AEQZ6UeIfxmslyRRKJ5mQZ0fNb6h5aapZHCJH3D0sdaQ6aHAGPuEuz+gj6RPpbgK0dvBWQjzIFq7
AiNdDZDBqN5jBEUFblCwCWnsgxHmKX4SGE2f04yisrZ4pIghZkdWqzzqqKClSPSAL/EIZ3VpuOAB
drA1TQt4cmnD6hRpoCFoJbxzDhLUg4PuLyW/Qo5h4ynSPlnPjuB2X3t2D2/+ZbiJWpAvvhZpVHDw
fbjvGufnOIUr8mHnCyBKXuHOO3wqVcfsjPfvdDFJ3DsVZW7tiT2OwB9U0fNwCDYQTRGY5DTiRuSB
okYJ1Q1IjMpgRIBGOudkVN2R7/+RmaIYEdgYIc3kBtJQA9OsTsyai4WkQeS1KPTv/IdWq4RXN6KK
LWZjWA8eSuUM8TrOddmg4dr42pbWBLkN3E5x3nwv+N89WkoCGPQ1jnafTECcDM69SOFoi3rRxZfH
3xp5sFSo7hyVePSil+7VmrUzerL0VRqc8Rr8aujitJpy9G6luWWjDaI5Z8ZQft9BZ5eQZpD+TRzl
oz5CUqbEzwzcqyuvnkrJPk9woEH1yFSOHvUGCoOEEH2biHnM8IvRIQkwLZdO7mjEuNqX2PX8LaYS
lCrxwkxQbASDLXxW9CjSPerHo7IjwWkHxCk5j8uBrP48aAUXeQR66DoFOVyVco9Q2mL5d7Lz43dR
2B28jJ7X8H2JNVGq8Y3mdmYhUM1gPcvGFFlLkZSb37tZnTcEKyedJWyCb5+DWR2MkKhjfMWGMzrf
UM5IrUqDfrIGrvVbe5+11CQRBfO9Pz/2J1RMJsXMPx/grdzpQ+ToJTi+P5A9sqDO71BmHCUizw6i
0or2LeKgkYPv8rGYzeK10wN9Rs4fR3dB5DnoFU1Eex6gqA7lxrCFXrRbw4pvPN2kIe+CXC6KwOpA
jgE26wGNb0at+Nl7VwTXaTpkjb92DELVj03H/ITDd4d2ZkHMmI90CLICp6WnFGoeWA2pak2Tbz1a
AnvAvJvlqBL63pMa19bUvDF4Z1ECqAYW4w2qM09km37V/BijodpGx5ORF/tdyL+49KQRO59W4Dsp
kdzGd0DORJdi7HG4dxsh1w+NoKzGsg9C4vrPc4jKwxrQsOgm7RkAUBPn1QCWAqQZGdeuH7meHiWt
+ExEWyQyAi82wH1k8kmClO/AXhWg87gT886R9RnOFwHQq7Q/g3jyRmWSCmQcYiV7Y7moy9WyDFCC
38LZx0H5+AhwKR0pBRin2YuTadhG69IcXxgqHox3/0O90BGI14u1picraQrjZxzK6WM5HqtsQOtR
1g/is5XDQqk8984eG0OEL0Loof4gXKnfHewCFwQYhdvheSlhH53XYS6vdPL4STMh/GDKFXslO079
ETPWMzrVnqgbdWZ5Pi0ZW6divX4T6rDwIK6IQ3U/Isljfo0pwV9idKCYwiigNduUJO8l08inkAsL
5EgTAomxeonVcZdI9DROAesvEH6NTrPkJSYIoWWzOS/R1hT/jiBfilmbXpi842uYUSEOdlrp3dhO
z/DPXab/o5VR/NDLFX+z8SXQHX9+Yw9vieVLCctv9YTnaPG2ZUl0FVxymI0tqdPp18fVvMi/fmpR
trmr2V1EiQiRMUtE0t5ejvKukAy2BGuoeZu038V3hFEkJosjnX7Y3QS0IdfLEez4XRbExTRkZ6bt
i9FbCM/Q201HIkGVTjiJvFqM/ZYRhlwSTg56Wx26EVQhmoSGfd7kBcfGK0m8jhMYH/OxNMOOFObr
3St6kcpvlBKnfYIc5Dgy7hmgxD7dhCuoNJbuXz2FXnqrZU059CD9EvABvCjuH0nAksmNGB1LF/S4
CEi9Dv6sx7VnnTKnqjGjwvVZLXRjkZZ5UHAY+tr3Xk7VBZKgMo6rJ2FRAdTIsVadbZup+JGuKMyL
sl+yI3w15RrJCbRpVzExtGxr/SMGxaHbHwL1KS8cWk4eY2RyXFX/MQqhyJ5sfm2WgugvJRMB8Jyl
h/PJKBgo0qRyOTrU+kipZxX/TNxIr8JPK98V0JLbQpTUYQPLXgjIVC6fJX/FewYmJxb6ffGeh+1e
PsS924e/pnTAlUzIy1fmW2N1lAtaJEFx8u2lKhHDI7nmfsyGDcHgMLSps+7Lnp0MQXNetaqKM37N
3DalguAQaG99ZWr6upZVc7hlXG6iW2mSPn1oeGcTuVmPLnX5vn9j8W1vT1J+zmqUYehQUwLbny/9
bWWz9DPIg9+CD6HrWUN3HKM1gmcuJqmyL4e4q9HYvCpHrZgr9loQO0zR8lYqlE+5iWQXbG/wnh5c
jomvT9yE7eKqN1LGk20/zoHMY77J7nQzEKq7sx/GUjogGef1IYCCwMaSHnQ6hvu18y+NDurEBWi4
vdu56QxebHIEJ1qoQ3iYk8Hf5iHntjR7mUVq+/4RJpUScLzhzPXnMOWW17n6PY6zGUwlS09eZFZd
5ruJ/0eFx9QpcZMhhgP+L004ohrK/3NDOJ/RcM2JJuu2yU8geLZ7d4wz9mNT2fvZdDB8XSUCwVar
xG3BTU62UIEAHAMdeffnszx9fjtOOiXIbbyMVgm7SA0s6cuz2VYx8UmxL+URSPFM+eDNlyg0OFBb
kYtPilYJ41qJQqicQ1qTCjkjhRufyR9KT2XYbeelBAjopyJVTXO4HBp4WCzG0l+iold+ilklMk5R
YrpZIZ/A87Q0hf6mIHVdcYOqhdFiG7WMlO/kJwS2EzFrIOZOMmLxW3K2xLvCdUcDbaR0wVm2ngWu
QU6+cGq9f79sVEiRiNTOSJPtbTFh+k6ykMIKcbUvYeR7hFQLbcHi2pO+ryEYf6Q6+ZbmQwKAqzwf
mmumJhUfVtNmcGrpW/GR57YYHj+Wbln761XhgjYyyQ/II7ce7sYp/yl4JGSF+JZXgwibM9qqwr8z
47q+Egp+P4laT55O9Aj6LqLbt5ym4bG7f8t3pf2vHdeU1ho4/qXEfmRzW/OPnSL8UY/vF5bym00h
+wa6kcUfax1z55FQBjr/lRTAtt6WKAMic+BczePzJoftfVR07Oem1yNCo6kTqjuocRsgx5psSV8R
yRP24axX7V88163s+lPfHUbhV8eOd9HskL14VnV/jiYjnvaNN8U7Fvy0LsMt3tSQynp5qUapzMc+
ZgAal4iEChEIkPcCjxjMC67pYxexxHW2VDnYmfxca3Wbz9ILCdPT3TRctqFN3/9SEtmYNSccZogk
mPE0hB/aZHJF1i2xECoj+b8hqtBpCYPxkHbQ8b8vzw/COdxRK/8U5K0EOaXc2ZcP55HeruU7wJuK
LOwGn5xhPdm+5rwvMNRORpFk7mF3YaWijYtjw2g0v+5tXr9i9x0iz+m0Xe2Wy01ZHw/RgvbC8sOm
m1JKc6iJVh9RxH2lJiuVXE/vqdvxqIzMeE/cENnd9yL+m8ami+j+/W6Q/H6xMRxjKwh+vAzPjZGf
Pd9LsbnytnUZnr6o/VXGw8ITJ52sVKSAvLdJjdnoPN8YGL0n28p0/Zy1OzH51Eom9dnkMzMPYSud
/2ajWIYlhSzCo/SdNYa6llfacIhO1xDy4EDmEB2M2B5zuweAHZSz8/Nrd3H9uEym8Kb8YaqiLW0o
FIGxrjBowISoXGRRTjPIyYACBiBecKmNMdZSCx5rG5rMZYlIBP21/JveS5JxH5NR8mfpnoIE1hij
hor7o7CBO7EMxtRduFi62+3IgvU2lsa8k08awp3ygz2PtOZkfAvZj1ZCmXxXuprPt6jG4HFhP0VD
2ODZysi8i4h7ctbinSI2weaJuGnpd7wKNjbi1Yd19ru6cnKly1MPxrr/xpuFuBFTMDZWvLtmDAis
1BIWYrAZAbBv99dIp9BZTro3dzNT5du7KTw7yidtJ0RLXj8NK4BBtlRsPWT15DFh4Z1u+sUXntXa
6usuxV3398m7THt8A3C897xP37W6hIUV0JOJ/03tSxra8qWYHJDyMOKYycfSygDuF0xCZDwtlVkS
6QzsmjfQ8zt+D64PtPpAAWU5lZhGtWzCKc5VzSZznmLz7C905utAXpCisf2I7/O+mL5kdPGaNPhp
Y0M/GbSbfw9Ev75rER7T9/Yl/Ci41ej3vj2p0QnusakCK80yC0KEEvw+LXlq2QP81U+r7e5A8elW
EokMgvqfiQf/JM3k5WhzrZ9kixE9tK91qIElXkRucL4A9WeWpbOAAAJeludXRMsFU3PPDBsViGzi
M8otEeWrN3/33w75qrlH81UxxA1+cueJu15ntO3RYd2jxSLMHFsg6ixeGysu4vNeHJWKSRtOrOlZ
rv5XPEFgr6rFGECXnFdin+1uK22esajyjae/i+GeXV9tnVianQ89fOWYdVdkSO3u8hWQRQ6yeDIE
H/wFoZ/FCiET4NdaCVp1yuUfzR52JnbikJsCCMHx0HeeEIwMWs/4/tADfGxjkfad5P054TKdS6iV
iTEp9xsJswijgI+OcTljBl7yyZUd30C15zuBa8VKzthNQLGOq6LHfiijq6hpRIiEOoTOwV7bQC6d
GZhORZLgbVFP4GcKpgaW2SVqaupc5/djvB0H30of0+4jRGrJcobCmc5RklzO0mwGmuzulrkPQp+r
nWLJfKw3J/fygOLGpYl7srAYXx1Bb1hDmjubdKNa9gYCgutCW1uSXVWLbDNB13nQDajJNamVIi/5
nAsACAqH7dxShe4zYkClMIYbego9v5HCjoOHkZVSNAOfBlLv3SlFle+azOqARwkg89LPPLh10jp1
pr8DkXU8ZBb+a0yWE5MDU6xalGELra4fXQLURSehR+l7swRS5M2tvcHrc8lIZ1iyQaNy3buJiPDz
f/Hn8cLhB2v7KnTE71/oXdxARwXIdR2BZwB4He+61q7YE31/R1YdLHeNDhUsGf4jIUcGOwqXy3mK
JNr+HLxQQIVtRLyWtnz+cQEdMBYFQUAVf1O5mfzXqg15rPFCDxZFrrVRJWmdqMyEBxw3CDGZY5Ks
nErJMfntKnQ0CjsnPwToJjN4V/ZqR0lnC5CH6VYSMv86gBCc3q/hRvPVXePN03N/tkoTOQ4y7Iu/
nBPfJyyfnGetBp/+sMRTihWnU58+iTPB54YL4g7IIQuzwL6ANyhg9tXXolsxzAUf5q6XOlg/ZUEE
HVnaz6E4d3KlHfEyJyUkkmaQ1PhumkiJWzSgfd/4tBb/pNXHvT3BhykRru/FUdca8v1o/LRUoWeu
VRZvLZpLclPtDMstetmrJ1UaRB/blXhyeqsP0ahMFog0GOVCs4cwsBoVzmFIPBpdCC9RhBuYi9go
X6ZhcN2El43Eu2LJN4+6jXQSfdGzLFYhIb6ePkB8iHCi6cSo6nr6KEsAuwn6Nyy9m8iT+gWEqpjy
uol3yNg+kTzIDVvzEVDDK7LwjG2i6JbGunGM69Fu8/W4ty94REwAE0+4iGFQ9y4AXnorYRGPjmO8
qQCJpjBCqS2tkiQB+yHGjIAKlAxTJyShWKbdIFLE5CNNiROV6pSgqO7u95862Mba7LOE5wRHSGYO
0ZPXsNr+ZGKsyUOdYUwRDKtHP+MPBlE8rkLbtdz+jP3qZadF6M03GfBxYhhX3RXXlbE+vdRlVGLH
nmsS0E04nx8pBJ+Tvdr3F8q+s0CBTnFxwSe1WU9CBYb97aCeKrBT3Eef8i+Uz9OWxxK0KurANIin
AjYOyxF9XXlTXEVN7Vp7oDMaSVm7VGcic9ybJpbTd4n2ernlPi8mP2eGdxWvR93k1Iw/yR8WaP3F
yzRMrYuz3aC2R7HdSpm85Wugn0tqUzp2IYxg76aZ1NfAueuwf5t7jhwfoOGJb84gRUlkJyzF+M71
ez4gt02gx8/wiSQfDA8s2RzMG6mdxyWBSkpaEdy0Jbrkz4LQtb7lwece0ulZj8OdHBvA8cu9qKFd
gcjI1vVkjBcU6q53pqtfqeZFMUS00K8+gMyZkLXVtorBqh03Z13QYYeu1lh7wp/2V8n9GZWTrLFG
SzfIeuohrqs5NkBGw0fMILdM3LNZU1RNUulpmA/WOFrO2AtX5n+Kf8k7vFXI/0QFvYYGS7JxgNgM
a6YiVJgan92XmAXKEiGbYxR3JvXAgVdGk/oHIlnirrCJE4NpyQWCqykc1GUvGgqpPw577WxGxo/7
YhS0OS6IPPUmOOdNOOauzJXgGfbJlfKl32neuaHvVO0MCDxWbwPSzQ8i08lEXXGwDpW4uzW4ESum
G0xWRhgYzAX1ySNlncDobjXep6vGwIg7NGAQWJvzJd4/CUlEIpWU4kF2RF8eB/bsobktdw7raq8a
q+a+/QILbX3kkhYePPUe5XILbsaoaE2DLHv6inXFmo4ruiGp8y4s5/96iG0WNmyYAtOLvCGBk7r3
oppR38hsvrqfbQMf2JN5sQbbuJIEBX8iYljbhZYLnoS5BcZqD5/h42PeKpdQZAnsR3N4giPHjD0i
ZVyYmZhkR1ygW4lCJmJbxV8K41TZRAaB05U6l1NnO8iufkfzw1aZKI7GhsQgj2fXlpKZEwe8j2AZ
KBPfZhCqn8Izc+lsgh5FJNC6djafdnLxlIbheNuE/LQQawtva1kMDOq3h/NKZc6fTx1cyL0mcqYI
/qAT3ZSospbGzCDGeAw12NpLqMH8SxQ87846lupymaExn3UxHeR/Aur8pC0BWMzgWjlrwjubAuTc
aICY0HVwddByuIXL+IUsVqzUQyJAN7aT1LsGIOt1uoQst27CQnc2DIon4GE3mhi/jKJD5ZUA94fy
bP70adJ+l5A9PjyYtqJl8qpcvDf5Y1ye7f7UetvkEXTPQcLUGSU/nlMhCzGwyM0H1BMVabcHGjJD
HcyGcpKPNjtX64ecs3pf7zSGW7PhqkLGWYF8uzpe9vyYIjYAVHFiOq/2+VVa+BJ3rACrD+VJk5UZ
lw5vtRHadR+FF0F5QYWY7oTaIqOO9nAvxY+7kMGFs9N6cFYHJF0dLE3OXUWYgaNC4VQe9I7D/iJN
UUhP1dCNwt4ZfFGJLmJyRX4JqzAh5g39xJ9kCaDUOcaS+gPbjvDDh8RodfnvL3/08JKt367qVFlh
iBQ/ahiSrBw+4E0xIAdLvyc80osccaDn9SOvM1xFivKjlFwoPK4y6X11rFrKpXW/3UpCzIPaJVmK
1eTApGRGnalqLKjOxJXm/f4a1fEV8PHQpwP0l78cfhL7U9Mo2JrHMiiyd2ECaYHbe8q29WL0XJhd
/tRWAIsGU/gdz+bGdwX1Y/N36Kth2uW9BcmlPpjZSdv2RBrf1m/TIzLYRHQrUmDH06XBUB+NOt1Y
9JK2MICRTp2tLgu6uVl+OA8ZEmoDEeDQsPJpwiM6/KYivMWs9UTVPzWM6pOvN/ucKLXEhgkdOV6J
+EHpNAtJ7EC/hB1xoZIW54hg72nh39HH0vLKFw5STULTtYPpIT18QkXVqxk9pu0tedFjtDDnMBv5
xLOP9+93m1ybcmskGVyDq8+iciPQN0ISSAe0E+Nigra1gghZ2HGu5Dekb4+qCMaacsfoOE49Euy4
P/B72mKlEvVIAcoj50yUplz8nGXU5TvhmzZI7dgxvrb4e0dup9X0nz40T1KCkRqtZtBfaDhmbqUa
72uzlkONNnacK/SvzbPwJXINCpRuDFEnenksGb9NpH5R3xgJJsV9+2XHJArEFyNEGlQbXqmSPgeg
L0gxoOv4OtrjmBbZF6YhN0/S3htt131MU3fi7ggR/LuunU0Z3+cR32lqxwR23faWne0f0Za9R+83
8FOcSnfWImoCWXJa+9BNGPCykYsDZ68Tc28RAfdy+WZp+EyblgAnoZUzIVi/E9nIhDiPqem2g/G8
gF25J4U22a0PjfI+hkJ7O7B2jTjjiXCln3MRH5GLIR9BAg1aedoJXRvjeTINlaJzRl5nEqAOmnh0
4TzV/TzkDXyH54Zyj7cOkEbGySks3n+0RCq0FhSxqVhV+U0LvSwzHF8tlxrL+PvqC/WA9Fygx5xr
lF8dx6/8I2j3IrSkRF5T7FZhInK8aMVRl2cXbzwONJx1YiJ6YXF+CYgjG/3PveqH1ksgum//oFek
xnpNNm5bWBbXxDOQLIpxOKeMIm0jZr+5esXiavUtnl3qOMSVSUrl90kP4Z57fYkyRGvNyv9/Ue9B
6aHbKvpm2jXBKS5R5xeDrj/UdW8L3DG1awesUgSoNodN8QbZ9C+hyNdC/gy2G/xbjZydi8veXAHj
qiwNjg17eSpfpbebmN60T571VDueGiNh122R1/DOowLrvUJSu7sFgrST8hwgJ1l5NwDiQqxed/8G
5D1wBqLxfL/A2vnS4qsbx5BuDKojhfKQRPmfTAPKnvz/shawivASyjmsnzzDoENmYA9IrGSDtM1v
uU+iZKIMyXiy20Qs+UhYwVCFoIe1c8QURwMylmfPedaAnyb/cldceQ4ICUfTDlag57YNKj6KS5qD
5GkuKivA6WTSL6LSxwbI+TQTcH6KdaGJzTW8tkHbD2U+AfW4MERVpxEyUmsV385m1BsJNT/aiupS
GEbeknOoRSRj4cFOxC/CWVyDsXne+m/IRQAI1AMXie7JC8xkGNAf5xK3rK2efrXEPM1/20K9OR8s
mcfaE1xcVXop0HbW7YVqbcCrpLYn7Npm6/TUTBnM/dHQiuiYLl/uEjHC4L9bNXaNbsPl2qNzCJEU
D3Xy3dNTuyThycSTcCsHMkL/zgyt2Z/ORSUrbhcS2cDi7OU9+k0/UFx39/r2ABNRfmp2xVhAmGLR
IkpQxugsu3v65xHzWEMrIkAZ+Mc2UA3M/hsot0YcRDYq/oYkl1Dk1R059LDW151p6O4RGogN2YqX
jHTL8WIyGWVl5F4rLsf9TXZP09Wk8eji/qFzPVjrb+OI4SkOw7KM1Oqe2Jj2yWSN5fAP2FIDyfFv
MMUXalsu7pxofF1wTBCM8KHxXzDj6OwBFdZGzDEYvdBhmRELMM+LUkCWfd1r7Qcu9w660R+pHZXL
LC3MMXpQEez6AT3JDWXmUhc/9+6uQ09c8x1s2UVxhPTeKbhAf4HN4u92IHnJzjSs6Cs6POoxiAkr
JH/LhMPQGQGqWPb0XXdM84E27T3h3FJagUAlBagM6Eg3srbc3BjhgE5qFqRvmebAqj9/7L8n9NLH
q+6v0tN1zgi9H+MEg4ndB+jYxbVL3AxVP8QQjV4b82ITqnaWBqnyF650f+w57U7DswKadTrnWaga
LZqTANdfwnG3PuIB+64nVDSsFxyAatZ00DaXo8O+1pSB6EfRwfPdbaNXaDSr4Q0+rrbrMlphktRL
hUrYrYTPFfCFbkiGbbQUhjIG4AMAFHN5zM63c33F1ClCJU+jqFy51zHIAi4D1QZdqljB0kpHQWTL
KYE8QHZIhSLs+12uWCPVx8bGbxKGhUUIgayHZnfeY0FY3d7cgNN429kg69EUn2yFbrcfQf+SWdrf
9ob10JV3S//2xXm/tD0AGNl9Ie+bI7F26dlf5V/WWn5Le0YvYgFAzwOTttuaIsY6HNRWCAPJzGTh
lAFM/cPIgXzCHR2S4W0cN1WSFeoUDoY69wtGZEZGxPVEkugUOE0lro9DbVQOyTwkVtpbtzKqx5u3
pq9M3tJCs8dZOLXIyNEJzD9Pk7sPkxowTbECHRVYssJBanNWA1MLD6Rg8gWlJoFTa8PD2T5p42fJ
89Ojm/okNJpJ9DkmvAJin1OHODWhqvSWyo3Iz0rh0FH/qBZW39KbzMPbtHo/BrgyhUy/agwBN8Qh
kQefmCrGUbTTiNaD1tN2LoaulwE/AhQTWcupTtrg9v+41DZ2Cmssa93n4jUbe/xosqkA3tbSNq4/
AOOD6Hz/elZYHPyGfmZAHZbbIToTzX0DP9KwfS5RdB5LPUTXd1NEmwUnWV/7yfPQxZa0De3kouJU
jDExuDkTo/AQIR85YbVlWKqvApj2+9Ylsq4Z7xjuUo4M4JCVixVe6AbQ5Co7g53F+7guOtoxHcES
A2KtjMMyI+KuzDNpdiUG1izEqLGMnQKs1EyB8DW5q01tSmeo44BnWaWc4K9bo4t2OG8VZXbsU0RP
g5FhDGLjzypyu3nyNhlAlbNg38c9oc9j9rXCDOYmMnnED5C7o+D89eCsP/W6vB1ukDg+aXf3/XCU
9e3yq35JBuzHGuuF1ODHG5wbj59cj8ojTPy7CGXd6Q2cx7A1aUdNI0+/AUuZ5b6znU27bn381+U0
04kphNY3XQLyecghUo6XW86EexegJSfF+2uznYfmiIl/gtKy3OGvT5BNnUt3stIJh8qqG7Ro1Din
CP1SdqqR+Dnr9dL4EtDFExO+ciOuDZ7m2RPj83zSy+5SMH0wUczJPWKxJDKcaEw6coyMQGn1oh5h
T//QRna94e0R13yoUJfTYO43jxgnnV1KFvMzj1vbLuSC5M3FqW3hPk6TVSYu2JOW72ZBDurLIApm
0FJI4kdpR3N79OeW5K06CXnc2Po6OJzt9Qz5TIHMHOS+kvf/6EVsSJumfLgcqZrDCBbRVtn9Eyye
TrewF7Oamj2Z5PxyAnXtuQK0kBDFTOhhjFXOD0aHsSvKy25hgJ716O2tXawKtZ0dPgl2Wflp36T0
kIc2E6P7xynXHTERyLvT8qhqjXD1dDZrv3WsIWCP2IghGs+xM+DrbmUa5AkvzlqMlL8B2K+pBdEa
cFx7/6Gv1bLlG6vaxmQUbTOfarrKiKryh/h3R/GIZuuBsdCv3kxfqYOVjisXr8ZRCVQy6zthrw1s
gDdo/YF8EcoLUIlMnZUH625hTREa+yYb3irBBBSVyjgxnhMFu8+ByJbY1EPMWp2zch2+RArLpJcO
4J1O8cpFusgLgvLjmsGAuFwCIjDADu5H8G9ZeVCUZ3uqSy8aZ6jxbSToYh6xsuWzIpNyiT9Uvxsh
LwJQ3xGu0EQYFpSuQi/jet2QE96q9/V/m7tmtjOv7zPpPOg+47h3JvccF7qSjWqbkGJqBuvL3jhn
6HyLkCaC0L9SO7OZ1cl5SBtnnrKxx6lo8V5CY+1Lq8xJFZjhusoJK6mAUnYGBnE8Irez8DU9VN7n
6B8HsRzwZ1trcCNHm+p2qVTAnHqZpqh4V95JEXMOmgYLuXhB6Nihv1izXBtQ1rU1hpiFFi2rY5OG
N+7dbJEDOBCqcDmXRKtsZZkuVn1aL8smvM8IE5vlObEHB/q4evKbhsRwrAganlUoYmKXhxcNTgc5
8xaDGIfN6isHLWqQgCg8wI4gs5dqKuQVqPApIOB13yErHF5Alus7nLb1W3iMVi4PRMCNOdI2jMN5
NkXck1a9JV57c6JfIRVChYnuw70BXK8sEKR0dBWrAvzlN+GYt+aanBUyp0NFBs9bTSwcCh9cvMT5
ejYmZVbXCHhbABQHDpA6fflQ9axiYfP0epnZsUJ5wlSN3NZqedS65VBNXsIKWADV00ElwRiFIJzE
TEuTWpGzCK3Y25Zp41zPMRqO3zBoAE1Jbq6Zt9LDYuv1cUZvTLXcMOlkMpBKmAru1HwqnhHjkPF7
Wv96VJtcIRnD7MmxOVDj0j9TOY9Bh5/v2exAdQnaZt2dlaoKFTUHJSxb0NWjpyN8TPTvuCz9/C7J
kdZ/kTH70SofI2T4PUM7RoIgRKZvuehXb8sEx+kyS40jAQBpaKlYDuI6qDiutuOGDHYZENn+f5NN
q39tRhSOATdijLWD+RQqHxmjv8hdw5zyQ7v7X9q+7+qNTcyuFooCCkREbRVo+1BNGf8SSPrp115v
IohEuljIJ8qGfOe4m8mYTv5VZM00eWd1K/xnAR9T+oLyCp6teUAa+CkCyS48I7KXXbZzIFG5sluf
rFJiBeMKgupF3UYJzudglHBZY1QMpzxcvHtIWvHYYgB9c4MO1P3UBPsrPNh1cUeg2GRsXfDLC4Go
Z7DAPqb0UdW0loAtEBP1wLkELmf7YvNJamj4kncoOoZ5AHvKtSeFV5jlC9GzSLnyYPi+aw+uqLMo
gFsXinZxi5jTnkUNKNOmNNSUftcM0brXgTAFNrE7t7EFrWH9G0V2/tTKf409RKr0l9CIK9YAFa+f
ZPlg2EEGyEddiRz4ztRZjIhFVLJvdsK4GWxZ4Kszl7/VD47u0A0DrMWoERYUO6pEwcKRLlFJRgp+
D7qj/INKfZEirN6ictPeEJybITimu51FjxoZqVDEE9qpELHDvDsKJQWExtXxGOg2yniGAd8I6Wm8
t8GK4kdvnG5ZMqjHo9SijZa2T3zoGItPEy9fq65tjL0xR+Anl8cXTCqLXzrvzplAVFPqVajYCKaQ
W4ES7uX7kUApgCK9WlVUfgO4EPf1yaw9aEP1aA6PFz80p7YUqDiWAjA/LNL0GH0p91QWDAySgGgM
YBYdLght9m1KvdMO0KJJ+2qlfIBhFTlWAw1tuENsjIsO97DCXry2K1fD6QCoVM6FYdnjSHh/DeEt
Y/1wYDcH0iT/dL4oOaG0dhzSp4WxJ8/3A9lXs1ps+k8cAC6D4mvBEY+M1CeRGmA1xkp+qoi8I/xJ
7BLjeUJKM444OkigRAAWWRc/YOnpL+TvI+YHwKQTWCnKYPRsZlynmAa6Q11Ed1NgwpzIuEmkBMym
0QYqQr4/6zNt1MOQizk7TmymB/t5ic7n/4OG4JTKrZILclgemxUw8GoRsOEfThvvwI3OBA9TroZr
hp2r6XEu+E38fOGs3z3PAmIU8Yvh1+HLvatF32z/OcEGUYitUIXB1+zt4I3SJ9q6G67P8ky0LJzv
AChCyR4fBhwocHIRdRbc8/H/PnR/6MJLarmWh0j/ejXjQIRnS5gG5evKUMNhZ5OHOpFgt7/CDIeg
yJYmcbCqe4gU+WTyzpjY3eLDCBcmIiH9H6PhKSdVbnkjYNWX/NVnyQHiJCwRfkKoGax5ouIZpzZA
PWo292O+57vpSTarVyqtUzpyfLoVCpC5xsDovdEy5zV4VyiNjXVG1FdXjS6fiSZVHR6FK790Uc3R
FYtmouBdDkIYsevqv95hT6IlnQOfPuxu12imvU9C/b0Udc+t9Y0XRbp5LfKD8XTuCG8pCCL49a/E
hu/sO0yMdKhXBng8t76rxWMq04CAqmWjlWNQDgMvaTJvxIBjnmhlprcz2JBOCqfnJ0LBAQmyt5zA
ycAYXi4QxPTFGiVcXYayk/vtXMpdlJU7yw1TB79G9Mk4pQisC69/uCSQ81UwRTrNxd7u+OBlK5Fn
a/IROcO4pIVjuLVUym6+yQYZeGZbpYPvctL4z5xXoJjcDAHe4CXpVOrshhlj8uVZu16+kvWdMfaF
h3vZ5vEbzg5l0qtl31ajMDULzq5ABfFrDDwN1LfnWQEcjU5wy+4j3Jt6gLqg9FuJoIDOPZ3Z9W+j
oq4ha7OJcRhofwD3s5UcZ2cFqxJpkjoN6bOvX+GJjTO0VEwavdWqIpiVUgsjVjmmyP1qp2As5QzX
CPvSMohmKj1ur8uSWKZp8g2vdFcsX1rokPlOeT/h5kj7UxtIzMRcH29WlyVCV57GfzWDc77/MvDH
4DUfb2A2nk2ZMAp524gBy3r3fw07SAmmUEn2rLJdIs7sbpDORju43VdQA8GCxRqVgFnONKoI2XlS
9pe7PXRhxcpHA9c+SiMn5Jyxrk0+46DXJgRPGSR6YLwEAd6znat3n2V7RGeF5opGU8Uuo4VHGCFJ
xeMJ3vm4rqV+3XrsitZFFl3E3UXWPaCDygUzXzM+/KB5ElaT+uSVKanHY+kXIys5Q+o7RV5oCrCw
av08+tQv2JKnctnji7j9uLKDjLvJ9mc6/k46EliJwzhHsjIfjACNhUVv2zjx8vD4sOUGjYSFnLw6
pi8lMs1g4CxzqpV3ifPZ3AVkqlyEJDgIprkkuo1eoqtNMVCRJtsL5B39kJBbpj2EbReSFW5vdet7
hRQhbUjZje4CwQGGoqhfXaeh37axQcV1T2SUD768QP4A9tBDBCr1+HL0N/T51/Vwca2Ki/pXgiPZ
L59YrmRP0Era6VrkEwD03gmrOgYWqIPTtPaqmvaez6IzubxJ3zSsWT5PvP4PeMfwcjpeEk9+03cv
k3/5g5gkKd7cug4G/7CUQUXgv8zRV40QXrNhWVVMQMHCUzz06q7Mm75eYvK1QwIPBEfPc0uScJb4
Qcz73oJ4WRBHqJ+LaeHJoJJ9av14/zU10C/mv1UxzZf5d5Ymt0+oQQdmRgaZ/y/2vnn89G2Fjx7n
jrJso2K2Z+makBUBfbnWOKyXGMruyDbq8wxxd+aITeNZF9j6Vpva3jTk/RgtbRj4gxbt8k/zdECp
7zP6X0LS8LJLyxuy+GETS9xzjrm3DEKCgNV4geRB4KpABT7STZAWfGh2I0tE48KXXMv3PoENP2LT
yJSlGfdphtdRsvSpxQ2bk9Ygk6K+D3rj6rLOkiI9OfgxMN7h7ujq4klmf1Ir/C5fcpuCOvtbVwku
DShsvoxFnMfk22k7E1WMHehX6LyIfxIHI9DJULrPaRLtcXdr3+zlj9Mibc7fZkiWDRQaYRVn6qk7
SGtm/lKgvIm9HtsHPHzo7mPiZJceC8Hh2u9OUNS8k58DMde7Tgd8ox6ewQq6QkTPIevJJNatl9cB
s2iPsIFQDd0HLQJjkERFi22DkUT+/KNQkFBd7/ziKx/F66C8IohxBrEXUo/Reg0/iQlvf5E5gMtL
8BGLfgtDhuKS3Z22T8x1Xb+6OVLj4JdayhH/gPtD6G2M91cgGaR2SUaUK8l+EoscBuefLnDXwube
2uFB6jENldbljUVtmyomNfPZOufAFnqADP1YgJI60lu87fUbx80+g+ESfuvdpKkzH+6KC52yhTHH
Y9Y8Zqf3iprPjtRD227OBBVXKN/s8oW7YymzArxNpWQlRznlqxRYBaEonvmEUmvmTY0iw+jp5FYf
YcPFg60PmRbAyNh9OUmFuR/50rLQXQL7422mIqBTxIQEQMmpdb6LftptPt/cDHm4l6UzGdmQaZwm
lUGwA9pBeHPJYFFu2G3lKkcx6BECnlvNbU3NO4eOu3kGOg+soi+Y4w16u00ZA+H0vlIHXFrvjuEG
gtZpAVCSUx2oeDYTO4B5xhcakHk2kHQF5xQv6ajJ109CiX0aQGofI9kAOFkDAlmZI2MqAyfblM7S
Vc13yMYeMSmI7ny3kD+G94/7Z8m/A3Q5HI58XfNX+T0l8MFeERh+6mB4SbuTiidtY8grnr9T6txZ
as12Br3Pm94AKu65UL4CY9X35GRtMaacNKXCI4Nmlb8VbaE3V8HHBBqZTMPurULApivikRYOmARr
2Lim9NsGftJBhNabOcgsbSdJ7FIo0ez7pfW96wtXgpiJp5eYzrU4jsLkiuc3IIP7OyDxxE3mZln/
BUpwGCvs7b4sskqDXOWqne6GEmYFectI1M07ti+BPSkTyse48OsPJD59mIIAyX6X11yBHfQTrndZ
SHZdk5nJWAfwB3vt9eFRBi5rnfibf7aHTl4/pN9GnDv8T9OxkKiqzGT/RPbe/flUx5weca8L8QHg
xzIp1t08mGj5dKvRnD3Nam/dBgx7MhopcpCUWs8YhupIHNzGelMi/xGDDJeGD5XWiQbHAIB+qdBk
hADGTwybMTEllTwWB8jWFl+HcPU7YiyX6ByPVq4jBFg80A+hcaoPYh6UCI7yTgd8fmf/x+oytaZN
BicuPhgX5Q4+0mn2PInr7J7msVBBuRFh7KH+kE8MGWrfpm+larJ2a3Ea2lH9b1bwqSYGjYx2+HdJ
7Z9Cd6kgWbIBFxm3RR5/YRtkYfadhyDn672W7uGMSeMldWUHudv2b3+JYxG36T/YpGJkvR1EdsgA
ivn3DKJfm0O9eUjp56Uq2+1AVKEtkLR+NC1EerkEvz6/KfqSIyIxriVQR6h/f9O9xPq5NfpbBYKa
9EH+0rdngfZrpyaIgkxpAkEyypJXVpBcbxit+MEBDHSmAxUlwds0xevixzooNvYP52WZxqgAhnse
RMEutDTThcf9cbBJ5Kb6dW2kcSNLt+Hs4roGBLDmahJTmkQogOskerT283iIx81UATGzKdHVNWaF
lKBEc7zA8aLilphhRjEOII/g8FlLgz6c4E2wV2HpuuCsqrIVGJN5Glsc6JRRNCib3M4pPyFYw/Mc
7eekQHKK4fDVMdrYj3aY8gNR1DRXWNFSrpToqKzQ3BDU8uVRwUvYbPSOfltWyoUJF99VLuxnxPRq
HQY6u/FYKsAA0fBJ6Z5ksZuLyOSpL/3dMfa0LIrISYyy2Ki1kMN8Jnqs4AqyhyzsumK1Htkz9vJB
XzqGpC8RoE8QPnUfRfzAy7LCTYqlvMDrkj4j3QFWYr9AKcsGVxLnwOKkvdrn7/itsS2W0GKJv2Yo
M0fil7RK+vTUxjW5H1AaTm8C5M3zN5GXTks5v9lLD2kdY5rCm6yHy4I6zwXbau/SibNYLJJsAFRL
rk+X96pgSzWsn2+2FynNHjkoLbsQ5MCg/FEEx7EsXOBNswCYKC3axcOo5Ag8ppaIPXLU1yVYJCpd
Ssezt+T97ED0Hv6K6o7V39yP9oO9vu/+3VApon1Ts/mj1iDbUS5CLvoUrxy3eKGhJB7WHcIOQBYL
UMJvcsS0dvW5uThE4T+KWCcac/OqCe+9mhC7jvAaatjDrDfzLT0A/HuZhTv4DsQ0y31BfMq2K9+C
iTZfaVXO1zFULv/TR3ABjJRk5u/LZDquFlDh2TonffvEANUs6YfsF0WMX/wH9QdgMg6F5/DREdaS
YJddryRN9HBvVlaAYN/saXh9/RtF6aiOWg/Bf0mKd4GdL8+wzeb/FDZw3j50gjUPPlYy8amEvl0q
+eK2JMOD0HQ1TfpZGOIBZHKGW+bQ10ilXqIY7nHf79WDA0d6DzXErmbT5wKvOUeoqflMWyPRnDMH
aX0xNY0CZYf69u9QPOAE+n/lhvHSrlycJyHqGmglbKYLHLb8HUapQvOiT2NZqShF6brc9Ihb9oI4
cCmFMQOaaDjMkj/mFlkkC6YyFG+CrOHL5NIP9IGtqAN80i+KnOdnFn+JAtokWSFChDW0Nc9mJ8Rw
RpYtk2slLnMiOpa32mFbhDddSUonjDHxHMbieqGsE/azKCuEidvAPZFN85+ocg+BOeQWW2ZvqMTM
9d+NAPtk21rY7qyV9KLzxuEOYzEzv0ub1mEQ/U52MelP5nbVJmxYbNzW9OVzj9OLckkBMwNiBRmI
8tEgyF893judMPuKB30w/L2wacwyf/oH3E4DqM+4zTRZEnL2m/vwoY6xXMvx0xHNX5beRMjHnBhq
tnSkbDCd2uYWNglBXuj10RPkC7RX2Cvtq2y1Hexnu8KN2rjv/fj7ATP80BF5AqMOe8rwbgvvd9dz
z2f4xjlDDOPZE+vyyJnJWsa81bh46vzrzuMk6nBiwiiSa5votfLDZPiHI/7EKCCjbAIc+ejx+mSZ
AW+QgdQS64YMy+oKS0zBTmTabQZjz+PZo3khAG8bn/4rvOSLCEkJLanWFJ6b6+9xLYdNQvHPIR/I
vLBKDEjyJA1Jpkxo2ahYqD5K/KPjCsy9DuPPbe2Rxu3yNpoE7rDW4+TMomzrU9GX0txCpYgUHnk7
oQP3bAENH/0d6cRQxRRmPqOhZ3U5auqWHEmVuvjiHb5pzFqP1AuTm75RO5m31vv+WiASvKyHqb2Y
Pfvm70kaeBhActjZtrEvfiVle1H3+5CsdnZKsgoqgkK46N9Nj6HHKauYAbwx1Dkzp+ytd+tviDUI
sx9NyUxotnpAc6wA5LCmnbJl0K64pEn0OT1AtBWMCmB+1kXK73fEHHfft6hm5IazgCsrhE5Yvnxu
xH+RFRP1BqT8h3yZYweNTQBvJvBtaqWMz3Y1Y3R681Njsj37WbQCdBHEt6SMjCT7h+kO2lSmRxYK
7MR/7gF6dvBLOfJdwv96HbjwQbyJv4MRhbLKvgCdqVWN7htdWU839ghIgn9rSVubfbbicmm0Ny4Q
Etmtn4qT5IDhaEyNk7LKl+o+9spKg5/4SNq1yQa8XVdm3zDY5bZpGyrWy7uthfiKtwAbLTc0urtT
GADjyZCRzxDZXQDQWcBXkOgeY66rr7GZLbj38e9ph6Kk9lea/L7XUkbMFUS5c7BxgP0P8bLHrZ7G
l8EWsWfkIcgMwAv+2/yeh7CHsHGRnzyyQR3edjxddZQU3r+z5jm33IHmVlBMe3qigxj2xN8XzUjP
V2M81F0nxVXEnpEibBxlL2SyQPchQCSUHUe0dPTR6qN0mXxNPMsK7GUTyiVGJrdmwK/kR/LCB51h
23ortYwOwnFreT2zTUtNzJakmNJ9ZkBLU8GoXQ7G6WyBw8C7+qKQW6EsxKGBmRk0TvE4k2grWx/r
2hYLwaFsfnNkVPUXmpIXDwzrP6Y0ZE3g0+umummMbBduapoxELh9xpL6xY2n0TkseXGmHNysZDJJ
xCbQNXccs3G/NABQzcH6QyfmaiDoeHUAVDx90ONodA0BzBAMIiGnAah7VK5rUMiNWbbplVdKdcU6
aNiMYkOKa8ZmF5YIwnMkyCjCbo1CXDtcHnzzP2GmfG832YhobHCP9bRlFOQhzkode9wRMHtmpXTj
O2nw6oxiAKC3b/xDzE2gXDTNdhJx230wWgiuCWzBaOzy2Xr8sG40FBeU3mU180GXNHUJyqAV8wXK
kwMQ8pRBk99xg54TUK5+sWJrz3/sB1wQJbJMFv22A3rWlxR5zO/NUcFGyfuIy2toxIcswQQcoGtb
OWNBA5pRXHUgcvfzkWhnFzcbn1yEpaOLN4D0cwXk1jEf2ipzsPxVMiGrkjY2/1ZRGZ7tSnBM9Bv2
5nypTSBYe5GKRR9ne4zavxWJsGydV8zGGli5k3ThHT1N4+9SUXXV6kG3ZTavNdxvo7P381NfRF8k
T8r1thi/JbchWIlZAMzslts4PMQJAsMMjyqyYVOJMslyqYwQ8tg1xiO4yRuLCRqWb1rxcJ5VZIjY
i31kDdoucOAisjDfrqh4Tjns5p7A6pWCsQV3H5WFkj1oZavYrlIFllunAMtKAxL+SGhu9L/tSf2A
pllUcmpPBP+YtvpUejO3P7/CfLdcQR75sKUWy4mnFyBf5A5zB8UHkE0ppZ8+ziuLZaw1m8AWdtwi
L4I2U9nHvlY/H5J+cbwog63GXxGtRfoTnsuDXlk+xVRC8QflFUdRhUeW3gomeG8hpc2BVlUNQx4n
eg5B30N5F3ez3sZ62grqo3vK6RIaaCLwd+ChY+BCj3+ep1mKLdpBs9xOMe7ZnHfbNfDe/xc6UaMZ
IDE3k/9AKYiBgGusvJc60OwTMIXWABlROGDeMH1okClWbBo1IHkb4J5sRFtLFhpIjU+QUOeyPk8V
vJJftdGKOO9VI3LOVNs+v2PtB89VuQUlg216BpnOerxjXjyafG6Gr9bPc96n4xMLxhpfPnqMImqL
XTCcV98qJPBMOwx5j8s4JyzetfuNmK2viLB+170C1ghiSElkzjjq8nF1gumM1BA9FuGpEDHyGuIL
8ptIc1TwkjOZ5SCjUIHWvbPkrkh59wO+BMPl/lYyaVkzQksd535ydee4IC5PunJ5QvYfQzP58L7T
8hH419HP3kD4LlpsLbNyD2eRg/ZpScFusVchfWbAyFDopTrAcKRJnh07PeCEStlqjslbatLcSuRC
1PLfTHGER9tnv7abQVIsJ+Xb6A/maSch6QdpPB+t7QfaVRuAEoljhu+sTWhppbIHQXXEVM8qLIwf
cdqEZL1/Z0n9zORV2X2umbEsWq1ulgLaXlBA6SoD7BPb9VLYwVTM/MqYphinaL0KDKLy1AOy1Wk4
GEufIMpm9m8vUeICoIQ0We4MnSLXGu9fY75eo6OrKLnut6JJhffvEoxk/aQUh4x0ixYDTj2Bek3P
i2HP8l5LBfNpf1IR9VAvErYgGHvrf4U7FI/1YrjQKI9hxZ7U0NM5i+pTCwwDaQYInMn9hF8Pi1Qw
ISdMLQ40Uf2v8UzPtEl7+qmI3E3jatHVaeh6F9tDaSdprmeMuqrFP2Qd4LhHz6JZEb79MyaTMylx
HImFaPX+kmRMFwz74iXhroIkQtgTwAEPkNHhTVQ8a4NgiZruRJnkizI8Z6P8ubro45tjywvz/LMn
Z+YIWxu4Ei7vChacXuvYBglggwS8ybqpf1OK3SmcCcwNjdsU+KklOhYE6i1BCZukRY6seOwKuDOp
o72dsA7UuoJ+7Fmxs8BKiEPiM/z1lm6s6rTk3RgP0vtSO2kUZIbRIthrG5NEYJ+bXsxsq/Oyk/20
/gwrTVUBGJPTImZkKm662wIjvA7ig6USt/b7DBF0qGnihCSuU1Y3ReaHh78I3So6qBHsDw2i/eUj
leV56pAexOlN/Trj7FAxEYSC2ZqCPpH2x2hepa8kSVklG6C/u302F2j8qae/dFd+pO/R+dA2dBSB
1+Md2dlPJbG7CNq0ILaeyJInWLdpRYbsr8zZT2hI/oZp3ifPkZCqY8oWkfBCi+yKUxl6AVxBKCw3
sHXjdVPPJoqZk0JqfUv0K/nuWibMZk+ZQklsiCnGXmLt9g8K9HY/wD63ptnuGXp0Ut6WuI+1QcTO
E4iYY4wSjvWoo7XhBwD3cC06S5FuryNHdEbQiJYFWIN6l+97B0KZckiV7cjP9ZR7VTeASz1kky9o
mcCPdBXNTD+C+EMQ41p/VvI4ZbNeD/sXBTW+PP6K9sssIHhR3wDzgz2cdLrcDB4RZmt24xK8fwry
92BDjROD8DOPxcxByP+Zn4pXdo7muwDsBnoH45sN9YHzhTnMpWDRvkXdEzAKFKBD6jhAESCI2XEH
tzOAjrrotx25XW48D6hAni5gJ9xq3hk1/MCBexfdhB8eMsAVPdJgQhE6by3ktcaxAZ6GF7o31Uwd
+2ONoxZZW7pMT4Lp4bJS3ZDNcBfcGDJwPDhqs7Wr/QVzcjSNU162StqdLuwpwxm7URHMSBqIBJNb
Mkd5vCudzEEGdEDnpdZcIQfUgCsEweFottonWlXXu74sowpJXrg/9459xC7vq6fenbOjKNpa28sa
nUx9IjILvwlpvu5CiFTY6GuhYoDlbgH2JDsAOoAikjTMD94guYWfx78uQ//KbN7uMkUPHBgFZ/Ne
cVqjrwho/mx5vF3/8QOthmWlMB9uHjKfrnTUGqZxcAH5p1Redm8FuBpunUqy5Tq8da7sDLX4zIf0
yywQCMwbgodrLUPvv1Hph8O6/DW8WHeS/K98KrewzjkrHR7JeEj8izT3vfHikfLzqULXYVl6aW2p
dxBoqS1535y7dNPzNxlz0Mpw2/GzXZ3f+dwEYCpyJv88GPYz7oudMbbHRg195HdCggm4rFUyywCL
6AteNuZJ+cpy7nlShoz914EGiV8FbEVgljxeXm+O82yc8pPiBhtotgWl/Jtb5oMDf6aQEaIhhJH5
V7O1/N+AyqCx1Sm7b9XSNBE4XH/hI20rLk+qkrHiXIN+nn5r/uIUT2f4k+/bMQZvQ5ZApkP8YSUv
oARkwnY86hqFkmhoMUzJR50M5IQ+X9KD7ERR1T/QMRI24m+BHG1T8Sbfv7ZvaXzkVKdyc8ThCmDx
7b95dCmBicPeq1aGdGz7dHNM7/RCaMWvRIeKinLF0Cz6vOS117rYKIHoaapd2peZ1wW+SL5CfZ8F
X7Aw2oakKRKyKoc4DP8UUzVqnZ4nQEZGwwrc2RtvnDUctuJp4Zr0Y1DW+rIz7mN7RTdoxI3iDSvs
ZOvNn6fZeDLJ/xF0Ee08m0GmO5Qs3H4VW2Tj+bAP/wp8Ytgic1mVJcyb22qv+IaSfj1FbAp5qG0n
Z7jPw82xnksjqx8yEjtdr+9nSYHQBdDDuz5hIN7cOhrMe+8RqEgdXEQFGXpt3mHgb3Jp13CQfKCD
HegPyy6dCcO2qI9VvMcgQ8EE8z3pzK+Rb8A6UuREqITGO3GbijVd7tmkK9ro8f+63x11Th3vxIdN
f9ibP+y7952sc+7g8MVX1GcYsbQnNakjvsCzUCozOLgwZNP/eQz7CIIYHgCsPLZhiGuripM2w0u4
IfAxO9gsYadrD5Yh3ZejubLlkjJTD+zU3qaAIYtZiCWFtjDuuk9YyYBHDOMlpVdtDuFSfgrfMYGq
vAuYUmLeuBTp57Ag83Etb3IsMNqjGZDjpXJ7Zu93K79B39saqwq71LSgVNaNAlZiqrfG7p1CA1Vw
GSgeY91iaL9V7YaxGu7gcbVjK0YhKOcxGtUqYL/hQd5LcCnNkJ/5ozvx/XHohrjAZt+Uzrs9KlVi
omDD0Gkq2aJC19F4eyFMe+0iSs83fuVp7M1EpiRck9ZNL4TOfHLa6JHrxFYspYuFDh5rHc08eKf6
0yGKl/C8TQyjboBTo2dLDh3TsXlIiMqE9Or2Rr9ow7ZU8xdZq+KGAa9T3ls51jVdDmBC31YqxhbJ
P2RyImTGisitqzq/pxiGAT2/F0U56d+W184AKsoV/VNbCdEu3lXehI6u61oqs9+1rbaxcMP5dBYK
WyPXIpEuLiS+m7MlzEJsiTrFi3u4T27Gwqxjo165CBuFdydwbRhKbvQ+qWbsbC+uYfVJUOYAcwPw
TuVCSFcyqDdNJK42zOtL0hBnkzE4E/e5WIC31qnJphxyRnjWwwIveNMLu7b36h8LtGUMQL9wZ4Qu
2sdN9+XYyiX0t3e/z/WXctW5G+Z+hGzUqHBOXCwaQcWE62ECjdm2uKjKiG2RLH83WTq+8LdwRcmD
12dAF2RKpwNkik2JGFBYm7epKKtoRCeB0czhsdaGqUNyVvgWcLTZaJDap1C3A7SZn8BfJvOa0WtE
JAnzXeGcBhsqF91YAPxpDWnyEVZCO3ZLBzz6hSLiQ6+zX/90snFQntelFjwN8SeRHSB2WcWRTeP8
noDoAQX+ZeBLDDHQCMBApNNsqY99d6RBGrvCNaRjuNgoHuB8Guit50xL5Avkpe0uhjB4oMq3udRn
SlQOYtkcAM68JC+u4oJVN/qsPmf0eV99b1K/QgkVUt+HNLULRCjzN/0U2V6uqAW50hIlZTl4V1Sw
ueoRVWsjKaxYWBMJc1fsngrKwtRJC18EQ1aCmFmkssyebuMUj+zrhi+m5TM0eBfK1AOsZ11vyjec
b3pJ+cuOa8Lo8j4lxfmyiFWRyJ8G1WaGi46M5xJdKsVG6DKCngmIwcT/STvx8ALBwQL3tNQPNGiR
wOfwWSBe5dbnP2oEBVrojc1r5NqJ4ympTrvkbAI/B2vxj13G9OxPDJnqzIjgMauPRKpEg9UEKUBl
9SoOZggyOvuYywVsMHRR/ekJ3jjbPMoVTuG0NWZBzGjRfOTmCwgmZF0HC+kM9v3rftaLI3DlbNe6
Gao3AkmBj3zEYhCdlwzcFPPy3MPZ6YjLYn4Ih9deQHBsTf/6I5CvZZiJgtMAhCx9NEpgS3ZoJS9K
zsoM1IF3Xzy+RWLf1w241fNwzcMLwtBFgi5rVyprfns54jChkS0GhS/1vNneF2MrrqYU+RKdlakh
zVcqUMM+apNSKaYxPfpmB5egNbVYwy/Uumd6IYyodInP3WuaTBgGS3TA8IC4WGx4+jEPjcmGz9wJ
QF0nWDd4A1R1HXGZG8tiNq0xbH4C5fYarZAE1F+gPSe3BXu8rdrNe3fkqwo1JbZTfK6stIHHruke
mKNYlkbpa3h47NwklXYviktzt4cjMo6omTPbymBu1wkadX1BYCBu8v3FyK1FQs6LJptIJdHXLEG3
VYCS5//bcuJ4ZZXmLCM+DTaxQNnmk55c5JTHo8bFtt/Cp6KiEIt6Daap4EtKRV4AkKE/Ks7K3pK+
D2kuAcKz6ZSQ1DUHgUvXBVlL09mCW+2eauTBUzlalqs5RrNw+yO9tt4Q/+gR2TLN+l/czNqHd5Dm
MLdhVqcynlcxgOibzyEs9ufGD9KZ1sFy/C6mZIxMnuaTHEoW6rdSYrI+B7CuV6lmMBWX1Im5aazJ
zO2Csdj+vNDHdUcR4hPWvIBbxNFAGIiMJyfHqKwi55F5aHhq1E8o9porZh0BPIVLvi0BRdOPyhrC
kuR5tS8nyM9M0dnZwb49q2tP3mZmdcnh/v/64gzsB+B/DMqk6YZCg+T2/D2vEyR/EcZeIQoYHEeU
S2TBUkExSTCYvibbALDZs6dRYCyA5gLg7K0uKWrh1KjCfyJpQV5U+rqIzFzbJEP1/5BFaayCuE0Z
/tCLmvA8RCXWJdqsD9K+zl3LCMomSUyVhgA9YnK95yrJ1dGjvtzcFeULbLnCC+idEM/5edgc+k9N
JhW2dxvH5DL9CwJET0moJa7OA7uE73dmeSihB7x/BXSqO3sP7iApp34KczLyGmqg5Ed/JVs0ekbx
KjS2zxghpx92Ceh+My1GT85VMF/JWVcMOP6QK64rBsZfYXIX9OJ9JzMlGT3kEiMdC8vYAAsJSBFY
XZcioi64mmABUw/8hGKO8JeRD68iGzdJHvkqZl6mx+qqwab907wolcwAAzsvlhBL9OGEzDr6McL8
EY5zvEDhBATq87YR+a4QTd0Q8FParwAfG8E2KVDF0o7LCDn/6U58eQ//8BHm8Iawgag9KAAa+Stt
SKtIo2BNHofSwTeKD17qu3InWD0ZvTKO+AyFf+w/I5S3UWRBaRwjXl6Dqe9bYJECU1K7k8O58hzG
aG++l3RdjmW5LlHmuWxsytuI8jAPL7CuY+IlKyMjsFxFoDoWHKC2SPW8M7wF16bBzoCx4WQ3w7NA
0gdphJHohdOhM9XSt0XBE7b/YS3vtKWeNnjvNV/44NKfTvNrjM2QLzKvVGjWe6aP6J2xCf1K3upd
TpmRFQM2BXJD7HM3o5Zh/eYuK/V9j5wMjdUzmTXVgI+ZQyMLFXQvgy70SItNwC64o5TqtNAEXIBd
p58lqWlEmhKupqyIPjIflB7v8HfBjF4n0XT+xDTTqUu+X7X+fUunLeFOTNrEKekojFTKo/4xCr88
mmzfWSXJ8LzeDOMrRnsznzcKw+8HmNN8VeHedctZZnso4ydzkS94IdQZOyzMaSJT9Xeg7EfgL0am
yPBgfydpWRqLoWe4wEskwcYTHGda4drqA1dRc18SnLOpOt/7U9pn0zh/B3tGi9nXA4iJUctbAXN6
dZcWdarFHI6qATZ445HYPLpvk2PqO32JvkQGhlkGnTWCY4dGziOSucClP+VJdU0D3sH/9o6Tov3M
1sjM+ys5kBOZTlczk5qAiz/LCwdQlu9XwYVQTvF/adiajqnApJXTuHOIh6eEXPC98jP8fEczjexs
NwLZULRt8TN9t06N2MIyYQFKvQO7V0RRx2QvhxRVW51DW9PgR5WuLq6VPMw2rfPyJAWuWyutCAla
8p40/O9VhtBkdW07h52i+xpwZzMlUWz8LJT6epxLeTso6nTed7N0UrjfZkkrCqoVlkxgqzbsSN0X
wcjDr21IPocJuFYnO8E+JDX02w7trXPVE220ukXTceFVMxK2mNJyouV7FrfZ+VMZdVscLUAjyw3i
rvbo8R61IbYPeKKZsFFNsYkteKSpiEd0S+fam7P16sVq+M1glDmIRYVMxnwoDJRkMLbcpkrB4jxc
Gc5FC1wp2jNuY1sGBLi/JsgPk6ekh76dhgy0U26l3CnFE4DiHX1D0XS8QtA/rx0QPwdCGNJvaEK9
3AkmFhT7MACdgVkx5HphwIsJqgopQYSJC9ri60PHW94r50kbTqBJo9AsZ/Bh6Ii5kaVTrp+WssIi
v7oxtE7ONFvxPtX++O439lM57WGXyqHyUNQdEDMPvExzP0nrJVco+WK1t2Y6EOqTtBIDW2Dr8Tbl
BID8Xtr5xupVA/xytVTdM1MHUFy9OgJlHp0IPJZ05I84vAk9BkKTjC4vMciMJUe90Kc1xKRJUTyK
sqIVVcTxYscvySnWck82jOhzopJWopY9LFtor1KZDMLHk6eCfgCFe8NxFmRHBK5mvecReSnupQSO
9veoNogmFVJiuFOkIpEZgh7OnX3POargO4zJRNndmLz3IaeRo1Z8jkcymN21xR/vr2YdimuqXA1S
JRWikLjw2AtbvEqaklCkzy9oIZvPa7KjFmu3iVg3a48TNC5Nm4/H/aD0PSLGb/67gEclEKvwxUTQ
aAI+d2h0xVk3OxZ7Thst07wrTRrcNneMx0vaM2Ba+VxROQb5ZBoiYPTSQu7V05UZROh82TX1J1Lq
+h11YWLfxb1xCy4ymEyzXflnzHo+6+Rx+lQihRzt/FG0lVMVIK5Veh8HcBRXqxp6S8vsGTbD9uEh
IkLLH18wmGDvJjWnHWSs95+Ujmgi7e26YnTsBF+E4E4pWYaLU1k26kToJWziX2jJ4F97lvaRJ03I
a0WrCrHGFc/HwDLyVKHPo1h9EAFs6mmMDtsXC/2nuqNrnVo5MlGT63/95LV8i9tBo3bLMWYdODlW
+fjGNFhk63Lp3716wfapz22ZsZS/HAxLhW3w1adn29FIoPuVK8hiax9zqN3DulqYv2cy7v7NACSq
0CGBLFlyPWcSxbBLDZV/ua/upM8/17Ag15ly295VU9PAoEHeDLIrU8lDzRouA2DiJExHjzXCCuRT
76XoGkBRmX2jkT2c1ymMdRtP6UvImT3dJovf8pVpnx5TF7GhIBhiuGBRtYdIMDgARK4gsYtDodLG
0X4QKoNUWlUKgC2G/PmUsxfgEXqN0eDnxZfmM4tcmftkBJxWH/eennPCZEF8egqnFSPIrscRKRUM
UPUqwzbZEJL4jn2Nrx8lx+ooJeYQ273jSyDL0hcZefNzLpnVhaGRnyYPKjQjLLNeDgiWc5Dm0mfH
BO5faj9mQyJbon8WVDpWagH5f9NdgiPmRd0CPAFeO5xfLCqFuaCLXsD/oOibLnzawxeNF6BIoCWS
yO2JykjPtBTFoAisGShQoWJqp6hSdnWKqWelCzG6Ir2DNEBxaf1vNKHJlyLcIU4j6CajuphBKH1C
uPfuF6SrmHo+ceZyei1HXU/AjrJ+V0F/UNFY9LXkHDkvfLgwBED7sHyDHqhewxipGOHFNzOJ29P9
YFBbDiA96gsIzcwmXiSvbop4X1421yPXv1Dd2lV8JP/lM3bP8ydOTZDg1d+eLg6Um9Hu/uHvyG7E
7MKruGRYjnFwpQ554PGPDTKaz+r1EqXcYiSKaUqn4dbFYkhFQxcYCqngkMwPO/KuFABZQoZTv9SB
W+tsR6C6v04bxi6uHq17FjwGePcd2CNN+234nztRYvkEqJOlmDd7yNhI4+uwc486pNFHF0dn/np9
wNei1RKnVjfS4ukxRgDWSUNioxgv5AVPHua3MSKiS+Vwbd74iLWfkhhFNa3pXkEY6o24KTsqbiD6
jwVvCuEobWKr0aknL6vtR9mx867Jbl8BgDd4m9Kj0LXE8t/qfZ73pkKp8yEJ7A5UzWUFkwcb47ZH
C57LVevhyeWqkGukVFGi8vW9I0X74dOkYwB60z/ZArUZM00n8yVfYLi8En491sFvNHWvm0g7FwTG
iEA1dCb1S0sWyAc1as/s1mykr9alqDJeTGpkIj0aRaKykwMC9N02wGwtp17np376O4O1vJpD1izZ
pXjzaLdKc2MXao1rHw/K/VeB+785vX+uYbua+DTks23Htuwtk6XB7CBgiBM8nzVq8lOBClsmO1kD
M5o2XGHqZPZBYDfAElTmVw7iUWCjrK8BgTWWapv1aZFPpZWBv0sKQ4zige9MTkK2ESAFnxim4uk9
JH5tMOeD6YtuHODV9BjG4Z09lk0gkqKW2I+uHbIryAnwVaKMuhR0vufssWGy3MA5U7AkxDHIgu7B
IN7IMRO/hli52Jn8eYESA8UK2WjBtk2XwaY9d6T+TAInl3hd1ZD9XLN4C4Wdf1+lVXpMzEnqJsy2
p1Mqph4LoXlTp2AtsTFjRUg7gTjMod6DE51To47i5OuAkd/3oORyrwWfJXPvMGgqDkGO+sUHlyZU
CTG3/67yJFekU4WQGu6zgh5v3rR2/w3+J/IwGmOAkegbXONsvJLixS4A3+93iA3Y133di8+QErI7
Q0Y2pDHTRRyzfXje5EIs/t0N1TZ2F8+KE03kOiSMm8XeM85nIBbjsfGsQmBHMCZEm/zL3zDLWOSz
sU1DcpxlOqAT7EUu4OfBbwD8SRcXgX6T2YF/UXr//8r0SLdpjgDhLOAeLVEWV2gifOoo3o5ajKld
VEr2xyDjsftN52pxqA0Kb1rCekbZUbAwIdQEdZuV+HqOUNtsbN+bBjxt43HXU/W7pRZNtMUfkTQI
S2QI0DMBhWt97YmEnRR6Uan1dRUG39E8cvZXwQEyiGoKt4rryV+a9yiChpHeBdo6B6kAoWPXmGLi
2PLSVE01p8wMPEB/hQZAEIB+bdDjhsADwd8g1gFsNYJh+rDeHxTD0QjmHyHTVDfegYu0sURPEOg5
fyrwFjFrH1YD69p2XKJQw7HZl7eeYeJwkIZQreqE5pG60c/8nOI8QaWf4IQTmpknN8DPHllUizwg
zgR9t4e2FBHVe8xtuBtSp2dHSOvu2IsVcYFvN6TvarY89ThKYTCn13pjzzml4iZQQSp4rVswJXU2
F4ZOmeK1fe4lCck/hNQV5tBlNICcdbELSMXtLiw8Z0lZNVzFNPi6aGi5OvLs9bDHKslIMA1lriRs
Zn17uEzyYLvBOfua1eRUETjCxzWi9tvMnmKPYLszidwWvmlwOcBllzA6NiaZ+tR7wzIAL7Xh1PO5
jx5T+gmOdnEuoh9cKiR9IXkQAnVEpVx9TvVdsRHoyNgtwczKrbazS+3+5XAL8m048GmpuuBYbMaa
joS2xh8xTjKs8R0sjtO4xWXc4b+6BSToKY0PxVbPXutPwO8bzDQlZyZhuWrqJstGRC3xbxHYs8/F
GP8zveBmi7KF8jt68KmggsyXKUYSRhR9wIE+JPwtOjBRWOKeHm1bWnnQwz4YdlZQHSk2Cy2En0+k
1fz3CqNe3sL+02UJjxAq0hm49yzr8qMNnLDDIPIJf/IvnQz3KPrLcPv1GV/zo8ipda6vUtY6OVq5
yI68VspOBvP1ySJh1If7x5oU8N/x2JPgTyBhSlXg4F9S+x5b+fy32sQabD1rni51FCVz2GYIrP3T
sQYU7zgtNa7YxR27Db7kEnC9KqWVdG017heSFrqkQsO8uuSXaI0FJxUufWvrk0PJUgPtKcRi7l2S
3b/X5wKNjUyYSyLGkU/vCFm473U593NO6KGTJNll1ERnFIVW6U0DpOJSpHr+og0NhiNsAT6a6qGE
QrCD0BCFE1zXoFA85Irp90mX9kqphIbud3PQw2Sch3HMp+dNmGduwy8YdO3RlSlWPt60tzf77Fid
5reGRqN6vzARsJJQNFjjvNSoiGu+KBzS4X14bRBk44bTQy+gL0f43CeSp+QYaGEmqhv70C4lh5kT
Bxe9sFlWr7b5mLtBP2rATU0Jqngq67lwSpohV8xElye9vDXHiSqKfJ3ZiNjv1oleJA7SR9KzGe1t
qtMwk3Q5N/kcoHZPLSUI2g0SC/P73Pl5PGKTefZk/PIiGRnOKeR1OuesHLiF7egNV6IgR60jMTkl
6JE+5OCrIGeUuHvn2xejzCuc/06zSScpsq9Y7B61RnQSxG186sw2mw==
`protect end_protected

