

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YeJs3h9nPnCnr3aRxIBZUXmhDS7WeTgKjgxxU15evXAwgLO5UoYuCJb2fGld8H5MyDQGWc8UFp3Q
QS1bcwQeLw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QMDnsLueMbfhPqb347LcBnHgrgkl6fbZ0QORe+igLd+Fn4pMYglXhNwzAsr45PWnZnHEuCtMe3Am
9p5sJ/ms8icpsPjNhMihj0/+LhkVUeJEYGJR6AGOi4DauCIoKWFsirWy53ZScEPa2MEe+a32HUq7
sCpglfzmrbsWEab4EEg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F3FpAl1oCeVkGEm2PKCJ71S6Z3CGasBF9SuzLFWQnXwmvUuKd7HyekhOce1QfyX+pLQcgfmP3XmZ
qpZIDWOrbZbtPCk3pZcRYdM0rjk3gWPTq89GN09GyodyzYH5nERal74RXFzqDSlXYzgzDvsSzAku
WQ8fc8R6wi9d8ZzaPtv7Mn3RMOg32FvlzTpy40zwgHFS17RZjspNh23gqb62COtY3bIw5wgzOnnc
pwYSu+4rxmNM105eSJdh2TJiSEN9+pTEYMITQ2PUZ0OLL5Qstj3GHFD8/78u9ynXfzh4PnzFHX+c
DtImYoh20HOPJeCFpBeWPHfekXHEPhbC52n0dQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lq9ua7Pc8cPhzNKkRvioUx2DGTzaswIzLnIP4rJJ3cLZM5wsk5kiUTKl9rdBpb7G3yE/zCnmkGDT
ZEvIhQ4CGdpOb9ZjoYg0BIc1GhYnGIexWpvkFarqP15NwctZCibdBpj579M1D8fvQ9Xw1j6ILLQ5
gUYJd4OzxaJCHTNx0vw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qzr81pSyvLThhRepJmzjPLJdFa8x8hA7KFKfUSPL+CaCFf8sC6XyXYts+1DRzPvdthUp8ISKrFAv
jy1EBIdnZB3D8J/YmjzA1s/E0S3V/3tyfjjyCDrQgRkpjqKN1zwlXCzBMyGSBWpl8ENwa6XmbY6s
fYy2IxFIrKpit7mWPaxU1OjywKhHRwk63dw93KzE2hJmtDZhJmXSPJNkgusdN/mkZzbIYUj8bMZ1
mRTDgqzRIp9L2zyHSB7GfUn9cIiKtJb71ztIZtRMoFGfKpLMWPUiRhyoCIz55vgxKfE+F3ghCh2A
ig+nnH/YWVIR6bKztafV39mEL7utiMvwk79iag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8592)
`protect data_block
SLfECvTHuK6E2Qj0XrUW8eM5gCCnJ1YjAUn/mgWetDLiwxYbZryTiU5045KD+iJ1npOEh1kO1wg8
98NUWtNUyPglMz0Yqh6z+9cs3fxPzJA2zddHr4lNVZ0PC9FpPQA+833GtTVy5VNuzcfPmpCYQnRh
80UyDtbB5KAiLiFm+K9RzG3XV5GSfZ7EkLBwYz/moJuZLXro7LQ4e+rU/XivebYMGbwGvcxF9Rpa
zZx+ShgC5qjppj35Ilc08qbkFFmpnfdy3xHtHPRIyfFdPUPYIiQpySoZPgEK8jvCacTyGS57vXoe
jCKplqiBhdoPlpjEBdjESR9uq57led0CuRmGnwa3lliaIVkUp5UE/B8oHEYqvVinW86Vaayr66iH
st2/7onL+z+4d5ctpfa4HqAtsSBxdpvHj1hJAAOJY6bhl74ca+9NPNTRZjTVty5Ul2fJlpVX4ns3
uJRcdt/rjxkJi373PDF6EokvRW5oZg4qNJrZTWZOw02/68BItuJuVOB7UDiO/knG5cBebPJwd3cY
emQNaNsaE1SAwYU2fBJUSzTfOyqAUWjDoms62Vhci8DKVMSiik9P8uhToY3BF12hA2eg7UEMKmcy
Se1M7Bc4++NdIFibgSIlq8OUUYdQR50J7Mr+Z9MpbmEiIGcuukT3E7QAxpM+Vy+m1DlwmQwb5k6N
LbcyhPnq5cMZsAN35/yiX80gLAM9KGzLr6QjiAdeoIETCq9LdViuxnas4tS/7DSpx4aTPZAohydY
zFfnwksm+PJqio37e6Pp/rvjZ8l/Pq5oc1nVKdP5vf2PVEid/IMa1a6WhUwE2GjrfLp0zo0UabVq
CvEEdScVdWJkyqGQPrMawTMZYyREXjKFHweY+d4Kj2e3HNUzkjgP9HkRxxrMX+VXw0mFq11KEEJj
m8K7CLV7tjbocAYoge5S7yPLbjop8hFbQj/Ua8gZDjf98BccgkXNMN+uQMC6bf95pHNlB6vs3Rti
pCTFzZr4UksNZJzYdwmzyuOCt+z2VbDhdwu/hUBoZJvZx46kfaWmPnIvtK6L6ppw1vviT1fMRg5R
uIDPk2ekZUSsU47eWksXGfwHcnQollx+q2vamHzuIP5u8e84doWfMTQyfZfVGcZU9GsP9MpsYldH
itIqTmpMQt5UMMSQOSAhmapChOz3ZG4R/tuveh54k4geyCF3qC1IGIFMprTpS2uCCFaa5DJ2E/4c
4wBUkqU+A57SRFF0AI3QuO9ZXdCNqJuYCg4zs86DGHNJK0ufOJooS66uKrrSmoU0ZNyMSGmnJiZy
zWoDYAjXwj6PGgrZT+HftSEAkezEdCXSlrquxXQgRzmGOufwg24nLR0ugVkl00jeUueqmOJWwUB7
DpXD2Ww/W9Ce3BxKNSN8yBz9A1Uc4VhVtuEeOSBRpE9UhREq+CVtybmV7hfGrdKr8G9jla6Iyipt
sUbov0Sli4UFzSI8sSXi8rmpVWaIoQUePhdjRzML45TICSleBT1vc3PwScU2lJsei6TUCZULRus1
P96BOsdP/qWXQsfZ3EYjqelzsoOA3pbuVY2PO3/t5irGZgS4rr7qs2UYCFE0BhQOy/0eNan4+kIa
8aDGG6Ols1o3LBzwh3xJYQzMofF/+BrE4zhenv5FI+ozQ0TUENqRYp3X43jv8wCC2dFzYrnGbpH7
0hRsgTWN4J2QmMU1tyZo0gfYKMDeywbhzzGgnjIHGuEDjf5QxfjFc82Db6SLmzGzPKTkvUpeFyIK
kWPmNCqlzU3Jn2kqF3/HFN7zlx4koqnzjEkLzwkY07oUmOptXgOOLox6iWyH/p4GkNw/7y7aEcGg
sw/trrTpJ+8HO/9t23X1vxNkVdQ+CCCuklC5Uzqjibo/5w0F6hM8AuOw/Lm+KYIrjxR5bSRd/rlr
uV63Ht+Gt3V1PqKt2n8uTd3VTfiw8z2RqY+u5V9NjIIHb9aYJkPWjkZm6tLoH7jo1O2pQYI/mLMv
aKi2ozUZj0Y97xRAqWlqGS4VZbnWsQgkJ7KRtF44NokCl/lZBH4vHT4JixM7M77kpeXMnFtNbP3K
vTWfkOonMmqGnJHak6jb0XbcYyqZZS1n3Ouycag521OaKuQqRO6SE71V2zTDkuwmAM8kWNOR3HSN
Pu/BGZxn6iH5Dh3cuT0/ZIDgeiPfErFXWPqDo4DOpWhe4Jn2uTjucINbrbExOILi+sqCr/Ho8VvI
oqwvsN1IZ/V5D+Bwe8xFtKyWH8CQiJ9uRIfsRhwYgHXE0pBKOXvEgaJvgDLFOIui6Z3ZGoLnZp4C
eXYuUf6zBLwmBQ3EFLLti/VHX0SaM6BkdzZfxSleKoWY6ESH6Aztmsw18EokMBVjcWGknJTYhoMH
5FSceUL95soB27wCSENPunXIhBPPDTx5yTuvK1aJ5ro12+sVJ7dixbTrGx4fwovxvMI40g1IpbUu
DzZMdPztX3S47bGgV7yAgZZvJQUa2xfMwtDlLILO1gQ73+NLNg1ZmhX8VFWQRpbHKbjAVcGZrRVN
ux6gz5Baom0NEXIh1OStQq6WyH9oM4szZExkXeTi8+lXKsSOY/C8x/6X+WVCDWwO+w15QortjBNU
cgsPDnJGrxOOLytre02BVBMawyw6Lo03m7mebdjkZKDrMtsV/UA8k5Y1zfvpeiWVVYxBl3xACITb
MNUWWapj/qdN0Jcvj0SHhB/u+U7vKgtWANX8FO2WjopM/ZG0FsgTPnIunKvBG76thNbrFdYTSZt2
/Zj1kFFnUCN3VaK0F2FCLSstJEXNk7DzeZe8On/hDjhndqDqt7M770ewaqsf7Mx4AV19okryagru
pcNL4LXHF5YswsiqnYMynf2g1wz0tVaDHL76FtDAmZJp+WEnAPEb3JrcDiHIGGDRL6MIbnVCV0ux
K0ulZcVmXRnLl0N5mW25Ajpi9LgzbZXrnWIxghFe4bdslAbqvdxNOokLue4apiL2P6SSXZOU8z27
4GtKZknR0r8rtzHg29qT76HvX+spT059yo5VcpVLOEpiqTcB7JBUMcI2XFJBI4WT54KU1byWGAWB
fezOsPVAu0MjnGLBTZU8wMPQi4X8q9MaSpEJABreNN6Up5sLTBSzx2tiVrDt9CgoSovikGWvB7V4
VHgOFdA0TJDzTA315ImOeu0YOIA4YNtvS3nclJavqeq2BdWLBGISnHOqfFUAbCN0KUPnFe7JZI/n
OqfkQ1On4mxz7OXMI/0rVuMIaTRMRmHar23pfMIip2C8oxrkeMwVUrUla2C0YWi5d2J1pIxO5xkO
u2HHRIZc5BBRJimNQ0oQrJXDAxdx2oe2AqMVmEnqqzCumOmVVoMtl981H1DVP5Sw8bzcJaGpB6G3
4SWNFJnKv0C0DkeuN38qOuHcyBA0sQJ1asthKu85KOtwskpOqhKpL6xewlShJY2tJD5GEu052KEv
9blLvuWQf4XUu6kcPAn31NiwIQfzAcw3jGLWDLTkmZT5f2Mh0jmoeFZQRbVgJyLBVl8wLtdzo2rX
wtfUGl3CsZWlUOtOzU8S5Jtv1woP+nWr2mnXuvM8hgjRDx3KedWeaLMsDoUHolZ0+OsWe+ZjaTa0
XkYANE2uQ9fkAB4FPy7os/oHAOhHctgTZovWgwrn57ScJl+NEimHugA39drGUXl9Q83BzoUP5Qbx
sIjb3weXNSJN6hzizQ4y8LuyY/sP7tmVJDTEZ93lsAJdSRm1vXLeYJMXtwEAHJujv7DF+XxjT+vB
99AQ/G7tYzICGa8hHAEV2rRAIQGJfcfle2FbDZM5pOn9YeHF5W+hYGuXfnwaW7VT29svDho4CauD
jyJIIQsUiCGRzYTY3LeyBYCoEb91FRUmudLxurNCyWoISM8KE/R8EaKJckCIbmKODqJYM/mrVZsv
EBD2nVVKhuha5dUceYPUYXlt7lBiZTFZywL4PWpoVUvhFyzCvXmwPvV9Fm/YDNuvvI9RDC0VdenJ
yoPyj2vcW4kR0yzmQ0/7q6c05ZN1a7Aytc3AOkMH+4L87/rn8CL3d7rVGlCU/5qlGmMDLro+v6md
20V+cKrbAFV0bANzWGbMzTyN/MYM6gh9PrH6CNihOSfBbyDzdO7cs4D5IeVXiN0lxtsI5hh1cPm9
V/Q1YzJGlwgG/YGT8x9o9PJdhRuwEPCgm31+fQYcYqGldQWBHg5RvH4lux6RYqQb5qxSPIlCXHsM
2RRv3Fbqg1xcI12n3n03mpwXXavPilGz3iP4RLIaqYUCaXGxhD7qtRi7gyX5jzzd59MNU4azTZhz
6gxNgumhRvM8eMoKnd5WW+Cm8C4Jf+KanAefKYpbiy1Cn2PDuDGbS4BKgwS4z5xpLzyrWCrHdC8k
J3rRcTKKpu4HzJIV42syouI+LvUen9LGEzHBHnxL5MMGrciaC+F8/fjkJw1LU9fUsH7+jyc1mBUv
3YB22HN+PV4H1UMGXWJQo7hksK0+3gULQdMOJ7FgAcIL368Flg/K6reBAvJw6poiYsmnPjqdcUoP
fYII0DTvmJHJAX5R6WEvRKs+8zITESjjfBpw3easTLlU4Q3j+ShN7AEDEiXbAMXu6p5s3hqXZb7Z
bB/M/wQ6WYaqQk8I+iTlewYBhX0R2uKfdIGnjUH9Sabt3WlazvWcmggyzc5tuec/YBMxLezYrSgy
EIF6yTE43cAY71IyukUOA6yTBFYXD1uhhXLJOPvbhv15CKryBnl1gnUXyeBDYPRWyyI6OOTkegh5
djsrGsNLmx8O2xxxfQfxrKth0ScJLgiNNEcgAoBMeSWDgD0PBjtF6rMvFB3UaZqOEfwUsfNgMlfG
LP1BPTzEmiMGa7ZjzlSUG/DXnvj3r8bcdXPTT5e2FQetHoKZmqOhZCuwWuWz8mC8S1bzw5/6/Sbx
MtJjVVcgsDm89QejhwtFgKkRzn82/wDsNCBK+UwgqP+2xRDcUH7nUpbezuho4IsJTIIIVQImdwnb
YxoJR3Iq1QQoA4ud8yezyhc5CnWKKXDjqpGykq5oisQAz/z5g3edl1uvALXod2fFR6AthxP7JglN
dZGH5sWjvq1kr3PbnK3dj6o8zjkWwt6oCATR7cwLt6g7pnqbIVBn/N81cunQsw1IkrVNJTRGgG41
hVZLqC/oLgVrgtOsLnpg7LsTwqqau3i8y1jm25vMaoax6Tj71+7vsHATG5DKQRCm9JVyK86ohhpx
1wD1wiOG3Hxv4GQaSypWqHPjCwd03arP6kegG5KM/gHrPhzx3xCdzOJVyVsa17W+I6dXt28T/IVH
rnpPZ+0P52F5Pa6YjfdYT106L9/1dvcRQltIa5WkgTvXYL1moL0aiezNOKhJJHnTX5r3yKov7pbi
PspoplOrQdkx9nOVbA9iWTzu/867sKQoLtSFU/bZo+Wcy2KUCYz4jNZWpjB2W8OjOiVEXOrq4vqr
8dy1jQD65J1kyG17/qIu5GcFAiyME5s1Me699RntbxiTq4vWhF20RkdcGainT7NVcY6l3p2AQTu2
+2IpQLug9jBJ4eKk0H92qOdmyLUBQjIHeSlZ2Sx+zWiO0V3yy96q4XnobCdHRR9ZCrixF4yGBSs8
eBd/IwSb0f+iohUXo8/C1FlzdhJiPLHs2coa5U93TgRxGXuTucnJv4UBEFikCcNjLaj3btx86mC0
AJqBe/wVnSiZmH5qfElQBztYcj/YwYBbmEJsRtdR5RhHEcnM5ZFJyYDz6ccMh/0NbqwtXQgI7MIs
eDqFswaZeepKhV1oc5SGcHSErnk/V5TEfc2nd2nmFAn16XM4skRrLJXSKlveuPdy34eWxBIqVkgo
RJsnBcj1OuwN1EaZ69eW5f4icfIawjvQDTB2GJl29vBo0OyUuUKGKyYn1x7kn+drXHsb5+HZgQcR
R+2B3T9hpEhP2y42K+vGOS69UXW5NCfsWv4Do7BXJBp2+4O5zPYCbeVlHLfuQvUkCd9BMY2TpI3h
Y5qg259sX9CY1UZui1yX2JRmRuJJeAdOxRof7vyYPMUE/caG5wPqwHyjHAmkIvyfUHABEMwazQuF
j6PY6ycDzspTafbFKsx2mkAM+hVPigy4AXsgeAk5XBGFFe5QXdINJnzdEpRCOakIMCt9ImUZhnxu
97jstSc3A2rTXehnntasO2iES0L1BMcUJF8/ZXpG7JkryNdNw2G1l901OBhW+005srQdotlET4Sq
V4CmjdMIBR8wHSdoNJ21L6e/9QVagDEgbQgsOvxmjAScwFuH3rFauWcZ4P1fz/ZVyE9ZLXbCHOmV
OQ8cMiPng+Z04xnIwePoD1tFuR2jY6OhgADQQhaRhlcMTAE8gZJiszouOAz6AX1ms7t6m3AnOeh1
G8YV7XySOTcBAUDmUhueHh8CraerWVkS7NdHPh0N7qn+gQVRtt3irinG71sFlchuHJQ+jiHVlcI5
2HjhF3KLQh++VWSkVqWGR+fGJnJDcAZzYovmCobcLuitHD/hqa7GiiX8N2DqW1tpqO5j7J4JJIGe
C5tpIgznJ6dVJoDp8o70lP0qJX24/Tydk6qsIdaIHNEhE6MgL00U8pj2c+CE9kQjqCkWLc9k8BZY
MLxmC3LlaaYqL4VFR3GvuIrS/5RHZDneBmE2Wn1CGNdepdV9j8ouOBxJcd+OrdIhYf7HtR8Ec3WD
fLU0QMSoK43yo00OHhBoWM8qbt/pCTDcpkt3QIIjuu9cqjj71/EgpEYDNpxFJWHRiG59/R5BmuL5
FUWva/OJLcVv0iGmh7d0hCqhaphO0N3ujXUKDEJldDhNuvn8STVL4izEkt6ubc0sbUeaHP1H+7lM
Zxop8zoYRZhZ3v0JMjBE/L5fdfSTzhbylXIdJ6mTb5OE8ykRg9vpju30XMwKFuRk5L49p6J6h4ME
bQXagcBq1u/YBBdhsYUqPSBfV08hj9bFJUf0M/BeQhJ7EsvlAnpPp7RkbZAzbjpUGG6sbPUgF9wZ
SRib+4FtCjjZreNzoTorIivMf2RKnwepHV1XgdZZdwW3eaFdtrqsDmyD5tBmV0SLv3e9hmttOXg8
w2+Cj2d35nJgrJPXZYS2QEIZMl1uNy1E592gu920UDeM8qmK0DjpVmiS1ES0q7MiDYG9s80ANOG4
smjtS1OjoUXmv2JREuc3l7MrB/G4fHK40IkbdmNb7M3RleoFKUYOPTX82mOsErY/d/GkK9Q/29K+
14rXN/AVWZ7Yhz+/SlzWu+rZ5JIAa51HHF4VKEO32r7T+bP+w0myfnjK1h2oWSyHyeSaloEMSVI4
9shm8rheOgaTs2ay8OxuGfKvKRlwXKXQFTFmnE0AUayh7Q5AemtIclWKEIr7yLfZivogJVRaYdMD
4Kyr7FMSbVBst4tBYHSpP8Z3ep8kxKZ4zVB+akG4Up5tU7BLq/vwncJrAodft0x1Gy4oN2YWY9Vh
DB2ZH63g9/sHz9A/oKfzlrXhB4sKIkGSg6TyldJ1gc31YYSHNjWW6VMAgi3FgcUc0YoSMRSCr/yX
ASgE7Gn/IkyWldcAVlytQ72VQVs0FhrEQLWLJHEa9I09ibzz4L68g3R5EoaGVyvnPLNsUoGcDvyQ
zuDqeTOthI4hvnOPuzXHtmkVpsUyZKpuycQP3aWMzbS++CGa1KO+gZXLX1o6It4eJaAcqmcujw0X
gdgS+CJHjfavIGhZNgAflDhoLjYtNArXPWLKaCVDBejgFDA8PY1jl6ixBEFZW6Eb2UDPFrPNZg4I
X+tapt/1QwlmzT46gU+fgDUvi7AVxGuAZRV36gAc6l45+Cq4umyy3Eqa5KFX80qKDUcoSiZei2RB
+Pd6F2M4dEK9vWQsWhDTE4zjBUSZ1GAnrNvt4AwJgRpE9amIRyydl343IBJryXlWcRz09PxW5vvu
AihnTTeKcaHa8UVN/Wmmu5KUn/52aLrcYEf9buxsxisz41CCHvsZyWgazZrrt5cckljb5/Aa0/iD
7CRnUfnfjy9mutBY8yQFq1HAtsuTmxYOXWrCw656PxKUxEg/s9jy3V7Zl+yMjgUFcMo8kLeh3MCb
NRjsnOtgRecFFskdjJaLD7Hw7xvlExDnkAfSP+WT2J6jOINje23RSpXDbXoFmutIVAIg7s9PtPHc
4FVRDWmBuNDkYqMpTPlLe1CZuHFe2U3F8PiRjRMr82NcbOypvzmmdi5G1/ig917BKkLerDpXIypl
tTzZ1/fXMEZARxhXKRDdAvXVHrl6bCt7G7YySUAVz9jKVH1zHHQgCg1DUxzgw9qBM7FssACjpRdy
t3Yocb5LilyhXEFQHhFLzuw0CDueo3PXo5/HPdGj9PEYGlro04jmPQqblku7w+LB1b/Ma4j1Mc1v
CmLPSZ+qwB1atnoqjdST2WU7t981OzdGFBkkDxOI6Lp87Z8c4Anx9Td5a3GKoEhtYxZRH8f4j7VH
GzP9ChaxHLeBB9BxOir6QLXyJO9iQnJFacMUsDqFEhX3nupVTxi0O5SFn6KoeN788TW3q7+ab3/r
7zdejEsJ4geZlSq+16cL1aYFBQ+ebsN8PiRdV9jh3LRWjF2MfG3PyShPHzgLe6MTtUFFRqc8JhtQ
IaEdLU3FVPnoTa7/0iBKInzjSADY/GzWdb0PYNEXEwsyLI1yJ+NgC8k1BG4GIVHXC+t0XUNmBaT7
wqGCryPwbZ09ilID+7DbdGn7FY8IgycoqHXre24XNlyT46gqoeDyMmq6fMLz+36C6MJsn0BNT16f
eIaIKOiZ04lp6kDU84IGQI24cTef8m9ddOdYX5Cd6k1kZW2W6ZUWXhi32Q5rbwegjkrDWiwcAsxQ
1VjaDG6odNMl5nfMf2qXYZBojU8jEQdwPSbynZH1cV0xdNxQtiZ8yb86jF6AbJRbhitrZ7jLHy2b
Hi1OE97QyLfJOIUyCIEw+W1jDg15rKsLoB7AUL6+BklhNgPo/zuxYrN5h6vTrMO9gRxz7isdu5cu
n7m21FedWQGdOKab3f7mvkMYlW/c03rkFpmjr7CPe8x/f6J1M1gkuj9qIXdnNn6N5VoiX0AmWYjI
VXuIYMDTYq78NvAeOFh1zfKB24iVm+9b4RZWLkeqy5K2IFrqKIrqcQNB/heU8JgUbxoYewUWK61q
KU5JHE/0YiAwVkP0pW7+l0ct6zXFrxKg/plrKMVx9cbs2Cw+OPhpJsCBKJ1b3ioyxQShvC+3Vo5H
mKUXWTk3YpAqZWGB8eZ8Y5S3/t7DeqC8MwRlorOkrcLG0a+pQ1K5GyRyhePWXLnWGViXObcCkyzl
eOCvYF62hEoQDbmqIrVeLqMSVskPQZD8kvAuy2ncU3Noc7W6uOcT4gWEivC8yyEuwWII+/J4X9E4
kBEP+etXYZfNwahwARi0HmGQmJqlqH2sIaXMqQGyK+bJ1y6B70hG97dDJA3qY33V1Jd1WwGT9Mdq
GsO6HmdXbAHwXlDv/Ckz6up0raB8pxFved5DRbzQ7v/Rmveas5jik3LKrVqrysNqW1XeroytEqB2
EK4oqQg61mqklPXlTI2pT2HbdjaALnpxQVobEclPzqTHn8/ocSNrM+UelGZlbB8euMOPgvbiKirk
IMV+8DvpcquTMjuHW3DymgihQeKzr6FJz8jp/sNA05ugyAhp0rGXxbFTNTz9KHJi5mBcf3u7pcQl
sWlYcYktfrSTL7I63/T4NyJx2eQ/+QMJHiupRXvZdoGDVDJqQaC68GHQMG2TEEooNH6moWzwjTE6
0K95111OIYfVRtLNLAc+WrnyL5ZbreMsq87/8O+jUMivuEvx05gmF9NcqmlgWOIpHYDHbAznXdaB
me81L3Mm+9Ji4ukWdJZz2OqmIxJLrNZc4GetfRxDUuyPkPN8fmhHQD47y3thTzApQZTkQQkOApVD
N0fzueVh4QL6WVPW2PCVNFUn8+Abhqnmi62jcBsgsPoE7z4vA4dULStKYPKtiCL8lcJYBSySsdl+
eluzxlblK335ye/RtReNmV443Yz+rR0T6CApuspvoHvcZ7kci4/AvXkkJB0kOGNUIwgMw+BS2N/K
cKenZjSPGfAxtfc1BE7V3T8ePEHv3DbXw0/ttXSP02tf1hdsB8h7yQZfOysW4z42DyHLF7sYtEa8
/YR0bNhkEwK3vPtM/zc233w/PfB9TIV+QChIu/S35kIGM34WmjC8QUMZIDtkNtnCOp9YU5XK64dn
CAT4hG62P0Q2LXLyEbsIHMItQ4c+t16i2tWnrakp37Ad5B3q7pJSnLutdSY3Zw0UgNfQWatfD0wY
yyjF++gw6DztyKXq+KDcB6e50msnGivi65KB1GuA08dJ7OIydfCPOb+rV8tYzLezZUGNVLUj7AvL
cGatvqWzP3HXluZxlKYj9GQYLsQ2j7qlbXvEuVOSIFwsJRf8BF8ThSsgBaJwBWOm5/toM5zj7Nes
8ByylsXBaaayZ2jzeIwpWcLgz8jebOaIFCaXpLyA3mt8YcVbcbfUsyGBO0p6mf0jS1QUI293Zt5c
2V813wA2hKMPua4L5wnQnDTyG8+hcjHKdRkTcLmp2n0jXjpdjUJxh3qKFpXLAR1/8ZJLZXRYcS8O
Dcya30YbBpKY736L5ft0rzE9mBNl+7P8W/+EGLuGxrsuq3/BZ9hW6ZeZd2hS1RzzXrXZuaVO6LF5
Ovz341FllBLb/eG/qLCXItTVsJaK1uQbyVHau79VdCl+BN0EEt0CEgCGdfmiQnJ00dVz95gyidWQ
vNUfeZPNy2hI5ux+MTmrfEnV/H+oJg73E5FEJC9kwDN9ewF0rl12PX+RKwJVnYVCGPDrwSYX+9rG
wTW+n+PjtMe7UBiiGuim8ziXGU4Kk1dh25OUuCOZIkBNgsgrr67mzedwOePCPFSAUnPrMNCsB+uG
uOwnYSj28yUHvVdJhe2LRSPifwd9HJZ7swnlNQjYzvPuRPPJT8k1hCg/vORoXsryOGHZkuu/Tjbx
E44HQY4KP9hvAmtW7bzd+Ybf80a9RJvdltuBg+Ra5SYDzYfp6HWjof+lyshXB33w4yz8vh4fD4YK
f7z84rXOtj3ukG8cvL9VUrPJbBU11226Uom+aNGkWdi7WbTKWD7TduQaACsr+kDxL5FiAqTcLuGr
1vc8v58naOAbPKhmudfeLDDOltgeA546P4hdoHcJEkFjcmMFb9CyTVNi/5eV7pX94NIteKeprexe
8vnsuRni7R80ZAHa12mSfQ1VIdEY8a3jjXWHF/n8a48Re/u4yk9HKJaVKbLq4+U+F0bhnsewopiO
j3/MTs/VTWb1AEX2TTTWFoJbLKfy88xejOEbUMk3jEnG1K9bvkJG9tAVN39hUKBpHpk3Ya9Eny9t
Rorpj2laGYuIAto2U/U8qNpiah3Sj1bjKiAdT1ZQColENYT2DoB7HjkOjalrVC+rmmu7BGdE1MYa
2pGqH4U/94eMLsToAnuDlkREzzKGao0t5Ont8iuglECHcOj8HQphzoZNJ4ipfJJQORZwLrRvVYqA
chafLxN2mK4rE69kI9OIdgYXGvFRAgMjwCeHuQQHX0vjj4j1JLLOhNhb
`protect end_protected

