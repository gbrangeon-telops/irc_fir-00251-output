

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LQ2vJKYKktoZrCpK4juRqJANqbtQy3/ocOY3ZqWcaeltVJ85vibXAMA5tlVvS0pp5GAf58wutyGk
pEVV5Zv68g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oMuoQxHU8xamO4YIRqVhC5y86VVKXTIB4hGEIvLUCrdkutaN+fgAx1w1DFW4AV5UF4/dcrqjOzkY
K71n5sVp1APv9EcDNy4SK12rfM6JNEmec1W0js2v54algVfB410d4rZG0ryxf2jOEEtG3y1R1uZT
docKTvmf8ciwTam2vyk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RwKTb0xAeUUC/Zlh40ZbRUmoUjB02ejSjmyrw31uw3LFcwmpLfrEGeQFx9W8nBY5yWIBOz4idUaq
fc3pMxhJHFC7jCdnh3Y8hC14pp9rspO1hZLfCOxHKu7GOhZZlRDfFJE9YTYvNMQlQ719mBEfy5DV
yB6StZ3JnfaWR9muuKfjZivHmkGfCe6IBabrX2L7+LYnKKp4Bj89EkuYxLdjSsxwwHL5yBSzQWsD
f3NymUlojWqzg7COUuAovEX4Cr2S0yo+Zr9C4jJ43pknI50nQ+b7CaiUKqbCSj+K5CzuK/dZ/FYE
aO9kMeHqHP3vuIYIBhuz7gnYm8SB2OlUmalvFg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yN6ERKfUqtxcEaZPhTWcKmh6+v/ubkhs44a1yogYIxw8eK2NURIBs5ApjPyj6y69SFt7ufKFYnlE
zs+yxTyZOIDjE0iu1eOyuLmYVN1yfs8OFxlynJLngPXQyLVxs9254patixjWMGwWk4PkkE6mKJuY
ZOkdptcpF67u2/mYpXY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t5IcFW6UoqOUfYz1GOxoQECi+9Dv8vBS33YPIONcGWTXCbnB+Rky6dyYF4Y8M27ZqAdkRtAsKEP1
XbHsYeeN9tcVjnhsAEW+ZxZyVmGkxa8lAjUHEo6bSWwd4akFKgw3xIpbktgKgaV0fLwj4wfHvTcJ
XEKHWYqSYc/CYMdUUlUPXn3ng5DzustWIyUHmy7pVesXYKHPGiFba8n7HX/7Kf+2y3k3y0XUfQRM
e1vWugHsLB14SmtA740nmVJ5TRRb/gYA8FobWc86Rp4qtvRHvVvYBe1XopHUWeY1WEaPGutqYtgU
FjBA3NC9aJ03W8dZxVcVFZhyW8E1aSZwJp996w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1517888)
`protect data_block
JWQqrOUMotH7YZt7gtKmIp1FQZE4ix7pnWT8X0pk0wBKFNjrOKyRqqDT6PbNvWNEyA1j/n0dChdK
zwLumMkF9p/vBOlt/1iP3q8YDx53OP1mcHgIq8LQlQl8XVEkqOGKEhdvnXuJp8P+7Cqrxn48jrav
ur60OlgReGkQrXaBPqc8jI0NlGrbMEUTJ7WFiEceh+FqZtbjBjSfjKkYP8pUqq9IrPVb5+IbFgxa
0FNip8ipAuWustBnIvTHnDgOr6COJ53ju9QYHdMPbS5GsXx31mEjUJAEE8WsGH4lWNEI4wh1Sof3
s4oDHZ6vAL2u4yJamNNtO/8lPQJMmvwl6t/ND9wrmsY5tMl+AkocNYH59jcsbxwjen9Z0S1Womh2
hYGbMgcQOzhBicbseY3HipSPvKgkou6R0jUloSuUorWcKgdEhaiywyCgcGq+61Yg6l4k3hs0pQ0g
lbpNywSaE4HwLxoU5bWf3aw0NuxBDRWeTcI/+LnZRZKQl2YON8uWswcCRjVGO2ZLOzjF+pbVyyDZ
d4TkbPJlkNDjAn0wHjCrnUQ3n/FTs7SR8BvE0WaQtj1ZbdbE/V79bmiWUSk5ChEYK1v3cWtHulC3
ZZQkw6AXwz2nVo4Uz1VmU0Mg5msG10xsiDOZ97vcqVKRTctWZYs4T3RQeZuANMM9/54H66jYjwqf
AUGwqHxd8EDErB13frnOQ27pb6wy1sWEFS6TjtMYpDtuGQE+psFSbzOPKG3+jVaSsXxOuHqw1f61
rGCKDeMUow8c5fgWwofKXs5az3wgeBB//aNd11tGQU6TWu1yO0X1c6EBwQDvqDfYh8s+cYQ3HCaR
Cf6E+Z5SW5VvrolY3fwoh7S9uj2y5gTzgrugXpkPc2YrSALX9K13J9KCw78iZE/d2UcKOQ34qxX0
PSYhuWJmDAW6tvUDMHKiz5KsR5oTR0jg1jUi9k1icv3qf4yUytRSfJ0FiIeyUrfVYdlFvloaqwp1
E7Y6Rtapk/ZKI/i7hCCcKznCErFW2Es3XLfCDMd8rrjssAEamU4KI90ymklpLm+PalEmizLFbPud
2l4c9bCcU+pGkO+aI0IjDRxMZ5edIYS4nTNj4QwrHXn6cyz39DFbiQhVNghi35Xw5K5w26TPAp8T
sQSbeazpTgYWi8FMVqALiB3lJTiu5dhubt/4lBjdWt3Rotf3HzzyrUvr0Tes3KZQ++2t7jx2sn/Y
r4SwlZDamMWL7MGa5HkQgcB/VnVcT7aErWnyEEQImf2fGhuZckfRxQVsPOpgDZsm5UtfxEFvuAQW
B0LrykfErVi3Q259iKEuHluqmpsgskgqKiMwtAn5IELFQZ8QHFA3k9a6V+fw5chT2yGQEnbAzCPc
4tP0p1xnsS9xPTRy3xv6FAK7zQv3/av7IcGcKRWPK0OnB6DNAoTFFUbaJxHjtcFLni2lisTFGut4
GGKsxEsAtd1xLXPdf0JsilKN5VijCJgl31eI2x81NIlLZAWpBQImDjq7TMa9FVF4SxmWFlwN31sr
JoggW1YbUqUalX+jheFw9FMt6+nKQmw2XJCJwLwPjoD+P2df9oNDD9P3lrw5P71Bcc9TqKpbk38+
D9rUknJZiaZeBa2yg1kGGCC4+/pVIFnco+rGU633KwucetkJ6QpNtBctQmZ+XUnF41bd78tdabmh
bP5APTRf/Cs5+d6Comz7pooyaR/FXaF7rm5djbMD25BXJJ4mlx36Er+MUsWt8Vg6SHKgcSsx38nT
IWJ6Z4xXpNEwDbHvTAzywQcmLyv+rdFvOEUgJBANnTV2oRQamz92OHRxxWWjUMjwEJHqAt2kGjPl
5J3v0B4DKy2JC9+mnC10yIAJVeFLo2FcoUKI/tQfeUfkF4u5yl+0IoAC+ijBqp5/QLIrF1FCf0HX
JU3BIRCWt0h9jWSBskS7ZvHEuTUa7pIfGOfwFs87X6FtcufROtRuJJ8lSjbaJ/haHE7Dakf+ZX/i
fIhCDNhvAoV1xHlne5jjJwSU7zwHVVAPFmdvsCYDPyn2hxmMKU3+nuFYlSQJKh++yGgjaV51BIru
STjsNcynpeL4mnDIT56QTxyXYgAPFmMO19wRWtSqdSJA+iTSK8+Z8SC5jz/4cu8mW1we4HWTHGus
uoCWPhrcDVmdP3tDhVGOVvsHY1flXN/3/0kINLtTYqAJY6sqatjoUj7S0wJ5yGRnnn4Hlex3/FUU
Qr4RSFx8eYw/yXUqL5kt+pooPDb7RasHhaxTHvKM9AjUb55aw98gKuB2BtEurUBj17PrM/XvvH01
9W4lhdy/UCeO2qNYDQbNA1tFn4q6ciQsjHJwjOuKcjAQReia+GCK/EWn8kvj5cI+OuTveDIhJm+d
rtE1v9fjCaHDw4ATB6d/Zs4RqyXD30IF7BzCoed5+QWXQg7ouRqQDZI5IWNxLEyOZ3RhlORGUCgq
iz56JHwej0eTtWyfnIldoZwz83MNO9qxTdEXZ5BmuPwAT/vqyrZej3ssaYYVuGwRBy9G0WtOWql8
G9VzjnaYpGUxmjmJggnsZYwaXQy++Rw9c5EnjrliFpruGAShaXMCMW+SMOgAHtN87n0oio29E7oJ
auZrtj2MkRG3K4Qwy4CpZomK9DjjCc/YnvusGOLbGTfgEPWIiHO0uswK0QKvY0YJjnHc+mp0Whgc
D4ZdfBgkfg+UbLnrNyow+5Fzpn64qm04V/j+Fv8F0Bx43OGChgO5PytDwd4iq0bugCeRAckw0Zkr
jk2ahlLDzQTE+ZBqwFzGdFe6CJlKGAJ4ghzG54n1EuTnSnNkjA3rDUdIqExE+sO39/sQgmvrpfRa
V8GQ5NqtoeBYjzRARN9T43i+IxOzhmInOpZ7w3pfNpMNG25YA7vpApylzcBHZD3Yit9a9OmMXIui
nj3mS6aRHURUVreiR9pD/APIXCQuKFkAkSRqLwxI0ixgKkv8HJTH5Aupk4s6HCealIUYC9tNE/91
XNTd9Jtzsh1YaR+JhMF0x+IRCQWc897h1BRmTnzjI2LjKDML2RXqEVWSf7/VQs47LyFMDCIfGNgi
owjUcT25GwEs25jUbxfHwt3xy5HV+fLLRZEXxsV0SKLoyr5DUtxAyICx8C402GcvcJSGIOKM6o9s
kKEQ03n1Su3vBte8tFaljzOojX0W6SQgROVyJCTl4sE8pwJtEO+fngZx3naexYpfQr4NeaIE1yu4
g8LWObrerG0MsNSs0GNVaurg8xSXgXSNsVXaiKjt8064VQrXQoHB1plqRgNzbku/0mUXIHzrSwPb
iBZzQem8c+G+FteJEsL+0soMlM3qQDCNk1MVOVxYr+i/dp6D7VKqTcLncUM5Gsbboxgcj5O3osY3
SO0vtIi2WCsWeLzguX4KzVWRSIn6UWWXPzw4RxqyQhZlrBDQkGt888YaGrL5vODPkyBTK3V4Iecq
/HiCyQKLDxbmUBAVCcs9iprHkC4tw7poKU0JBJWEQH4gbyDrm6d6wKgp058WSLGQ5ifR7hG5DMns
tw8Mgdtok//9CclXFoMwpgbnQ5588ADdD3A5PEMJ7MDngPkrY0Jolz4LbRwalF/Rt9CD2V82Daxv
xFrcK2dO76SFEsGpuGHt0G70/xLPZW84IVDdy0cwTvHq7dboLXI1o3ecBtrG/emr2pah03eeltPg
Ud+mVMb1b/Z38bHYMwyFrHQIwGv9xuCAwaF6k5Y4PlarYjM89dn2PcZGHYK5EEeu+6FNV75mt6VF
zwtKDd+BtKO/bvAm2dp3Jstcz9iuvEmpOZM78giXMbjias/DwZk/j32C7BaD36uMisKIE+2WSln+
gvL22RRod1SM+XkDdSM31wksaQT9Oy+zyCDwpcIQNiUZ2BxSkLeKVK5rPuLqeX6G/UpGR/nUyS70
V0I0/qVD8x92bkvO9Qt4myxEOaF491d1nONnZcGf6HE/RC63cWKEAFfXW7Y+2Go7fgkihqmi8FrL
dQoNL4Csu21vTga0PvYtdvq8F5yQ2hjOFjTHbtuC8a+71VJG7YFeSCwb4BihqM8Fsgmtl33a/ymE
8+T1GHLSOSm14crpGNuzG0b3i09I/eWxx82Qj6AkVBJvl4VYMWoCB/X5ASorQh0WzY3vW9ECiKi9
iqVrDukm338N9tTZCLzdIsu132bk5nUE8G3K5nsJ6FRDxkNvfPuE6Bo8fbyflTVvZ0NBUOWtjeow
1Yk2koaiaqbP41ZAK7K1Azvmd9u768hZMZMOJx33M9D8VIYCTbxRsRM/oxi7fB2T2qfs8EbG5FIm
T+Ldp0n82AixJIwv5rZkyXc+KL13RtYZBsLy8+mDM3YgRgCBngwwBajD7beyG3A/6YQY0zYRmW1q
+BCS9KFGEJCzKAQA44qHclYujHtTbixxjQA6vbWVfIGk+2XpJggkplkjPXbpDpIB08HYWdj/51cn
syeDuGs9f1gVFrEtG36nQPyU4OF8OHbUS8C3vUkff30ZUhcA72NhgLKH/JGeyXCG3UpvcdV9SmC4
1a3cQfBJ4pwlvCmrw65sYjK5o9fI6ejpgBI7c+KUH7F6fyNbAmewkD3OOE8fLb6qDKBzM6vek14Y
uUiLC3F9HnhIPQ8Bfi8wUMrmr0yB/iiNtqlFgkhdjXt6apPsJlQxeu69DyBmduaY38k+oJSrEV7h
qTeThbCtdtwoSfHxwl2uNylZDYw2BWux5To/Ibl0/eoHMqB8nSAh/BTXj+/HMpz5SG9EiYEkSPPF
+NZqoeCLHN/Aui0zhpNX8BnLD9YApE89z5rGAOpBFEVJEAvkozjN9GzDmSzszK0D25B3Z/DquzW7
sFtEvE0OrXe0Iq4rRQIUppsXbuszsJq25FLqcDO9RvLu7JJzEbfrfDSGfDZfmRCBi0pDhx7yGYsu
2ifdm7KHX6YOM0mNWJ0tEM0nv2jft2QLbIyzXWSqxeqoS5j6aShSVQVSWwJvNL5/GvOKvZtgFVNs
25zWjW46khM71tPgIwaZVlVxtE664nTZvPzjWdEEX1dWnfJSvgMcEOh5ZKEZvaITisgJdr06z5U3
fEtI/mWrbxx8bgwlanmB5DDixnvY6UzPVBavnBmahA3tAIhCHfypL+BRTNXyQRvofqUEutBaPhsh
Fp2AQck2bQYfkiV5WfLfdHf3Fy7HEr+N/NM+siJgV6W7fG5Mz4tyFfKM6ViGTXpzV/9QnLVftl5u
Cn9AMfir2xU15dqwg/SHzvNf+7RK84cfvtTpWT0zX3CSUVwPW56xDj/v91BtfF0Pj3aC+tAdwS4k
G5JsUSKbxNOHDraFsJBpZKd8TxYdtfYymPTRlU9IAK6dg2Opwx26QhfoxiBjtvUjAsafdbWYieyZ
+xYuMHwP0Rwp2V2Xbgu5MI76/iycJ4oGZfpwaQKN7Xm3UL05rf6+Rm9H3qU5WeQj9RcMDC5q98Gu
Donnhdw8I+mkPYbmlwa2Dim6fjpKkMV4/I1APsy9P2CP9rUCoro32ihcUiECgxlrHPtdGHu7GLPf
4Bs0lKZzrcFsSuYKpTRkyJWBcAgI23j6ZXmv+g2qdP7IMOmBP0JWm7Qqze91KKl57ckb2eOR+5k1
GynOq3dDuRO3LJiOjllH2O9PT4DCKoic7u55aojMvXS50hYHAPZbSGo1oSpjbfAwXLLGPempDarf
SUFOyza0mzODYVntzPIgua6ONAOQFPPtENKr8Rix8MAdKOl2UOEipGwLS78EVy9ntB2WXxzZUGqR
q7x6d8c0+s30j7oop88/bBPPrTZ3YXUCv3eYbd+fITXMQZ5L0QUETjG8+2oPz14hBdzk3wwtJdog
O9yMBGxyGC9u2n/sYD5QIs0Xv1MeTjKimZwgVrpmNeHNeSTNuPo5xANYGxVbUr8BHxANeGkNuqsO
G9DMqxiDC9HG1ZQvXgHIdUOKRpns/GEMyxjyMMK1kmSGFNkKZkOV6leliAJplZxnEj7KJXZsTis/
w1haxv4jIG60YWCBb+Luz0+R5TJ6ECnc1YuOlMKen75UnEzMWVwhTRLaJzduIpWwTwGvDXlxvJR2
1RnLl8uGW4/X0IIFdKrWpGWnInejo8SZdDPaPmGW2sXET0bV0cmjNSErbuWSfv/X/yrtGu8ZTK0N
2LK0ROtsSq+Yhtc0vRWSLD0cZTI9s7c504NwGhmkfef0z/vH3dHd2x2/hmbrYUq2Te58B6ZeeFvr
A9nHJA4b8E9u3viUk6l3C8ddR1n6S6UaQh2S6ADZUbrKYL6F/2jawyLRxSHjLL1P5W5LoxzXuCFp
nf2ix9AOeyBtGHzq64eo8CKUYNWmOXf7WXbUGGGJznku3fxckFa6SToEzsChf88UFAbrhkQSq0hN
+NETHb5R/8O9jFHbVOxKVrTv9Yog+vglVEknA36UaOh1LpKfzY+O+vJG6cobtt0a2nbmQla8XoN+
XRT53MlQkeUlQq9OCLeQz5GXDLilHfdzyIyoRNQAnu6Mtotwx0/rXon8eT14jpwMYX9JmAEJZ4el
L1GRxl6kPE5FqGeOhnmQbqPqszb7knU/59Rdj1b97xMsUHY2iGfpdbayOvtopQa+gbgN9qZr9vDf
zF570w2NvebKJUOljaYJhBPieWfgteYLD2KBX/WL2j0R+Io0TUbs1BYl4SXzKZy0C/jf4lIJtlL+
uHFRmqH+J/DI5jBinftaL15mt/rel+otWsRdkLluS+ksGQ4CGgamuGJUJS+rRfnwPiiggziA8oQj
zlCcAiNkW6kiP+wyCDR3AF7psDc9ZaQFm2llqQuD15SU8ab1U9lB6ergecV4SrTh0XTnwR3EhxGU
csfSaJ7UEgdAI8HIAHZoIMo+9wYRJozCa4uJbJqh7bj7RMhd+lkmwAp9Spy82uMe1TVn3HMQ13Sq
uu7YBSDeCSd+35O+07KgtF2WTSR4rUCYdtMwNTmGo7fcZUfRwmAzWzwGaSILmC/L2O9A/PDZViU9
XGdENXJyk/c8JtBAzVSzgnjzM27icHuYJ0Y7K3o0Ug8CZqo2ytm+PQd6K76YquIeZWLTRsv18bcm
6HKXb9UD7IBhdKq8eSijRtmFegjlWd1aosKT6K3XysUveC4JpWlqLVGckgDCwwuHfx015ARSznE1
4s7c8a+GYjkF9Y/bimPpv+HxOYEUu+7/ph2sPvhWWOXDKyQ9WpHNeTxjx81NAGaAvXpfFL1ANVHW
+JD/Wh4mDvXmJiSWK6+NtDKPhaAt15WbwCOUlv8b3XBm2nSIg1jt/fB5S5i1fMP4g/ELFkwk82mb
1zP+G1AFiU3jYlBGk0bVkaOjojZ1IozfLrOw0V1otR+XM3r/7kcKxop+zIZYlIPE5ZwotczsSA0F
FyCq1pclzUGQtFdRTdTUpR9O9R2MAUyfiwKwyRYIyqg+1Vk7DNlkvOTE+Ubctm6Q8sJTTazVrvCW
BjklXrhwcEQTxREnS6zyjrfT3X/KrzW4/PIZve1+O0hvn9vztV+AY5NJ+PfgGEh72cifx5G1SJlZ
ofd/bckkFd0HCGIU074gbe9hVJWraSctoOAiwZ3wt/rH/gz6PTpBQ6Yt0bdZXzARH+q9lTlaSoxT
SmanF6ZgPvl81DElXKdGp6pwDOTlFMV4dA9OGuDc1x+1gzijWqxsoYyG47BoNx9Ely/k2tJH4miJ
3pc8mufRc9OqUA1rpaiyzg7qrfxVXbEeLOwixkzyP0zYaREoR0ZvZE/7/9C+kaq0sHGTfzH6k+Tj
WkffdCZS6UI0YhpM9kZ1kN4RKTR3Zj2n9Bg5q/W1236kKMUYnhvEtrHjG5dopLvFyB7vcPGRKfOf
nsB09kNM4O5PLYrDrL4jNYZqNmbSybP0tZ5RjnDtC2jkWdM4c5WMfb7eBp/CP9iUrTw6R3+7Vcol
NNmtggtEXEUwwxONlBE3NfrcXQ9R79ZEQPd+O8gNjlyZ2tvsuMmTkkABX8vmKN2/e7T0VInjIYNn
QZwjOigUuJeETM9Y/qGK3uyRL8u2ILymjnGs3LP2OkmEbFxUfwr8iyqMTJRt03X7n3tQFh01PPGz
Zcf3QKN2v4loZ/2a1y2f01qjWalaRketeYSmDQCKPF+rXweYCKM2xZZhyLkNrQW3FMOvePTZRh+I
PZzwAcL+yqJk79D1YmzGcX+cpqfSw80krPKqtvqRQy8V0c8q+lZ7QFdmQvVyyz6YoToRkTfifVJp
ZOXQKBZEC8tL9ScHfqpzZUefdH2aSCa7jk03UgRr3AabVfFPr4UGKvIeVtzQDfTU1YNfT7Wp15xx
NIRch9eP9sljMIkKxNt/DXVsYqw5tsOsJ6UqIV3Cik79yrSyqjQOnV54A/D0HMgNDYcGAxuc6H2J
dJQ0+fO3jTB4rNGJcuKBKj3LkiKCsMdjhroG9xBhT69H0pIy/RCw8dL4Gnc79+I33zMJ5nf6anRT
Y5OswH180Grsmd06ZvxC0G1DiQWKacoAQp/cOoRIu7y7mwx695sjiWf2c1tj+xbSDdiezcQr7kua
AjG7Z7ulWXP61lE62ilQKrPGvQhV/zYFHi3VWbeJYamFI1p0WcOA0k2AatyTOGHP2lq7aMm6gYcW
bDOlgYp2uxpvRzCP7djYjnz9VQSVpG5IWadcO5XiB61SRf5cJibnBYyXR1qSnma6F/jGAJxR4LLI
nZMM6KO8UAANIDYApQHc3Osneumm0Lo+z9Ay0V+za+SLmP5B+pIp8u1TIwE3QYJHkFEgGOS7+I/l
eiIBK21P/u/hlcQgk4yYAK45svuycZL/hSBFn7gZYC9qUKVgkLpcY+LXgcYdroiNeOXA7KI3PaSi
ko7cWFyhDQ/sc4EFi1mzyspug5hDSfsKyxV6GdNVAS3s3T1uZ3cnuuD5h9Ux2HSNFCGIn42Jkkjx
COzRchKVbhYhaFrzpJ3jBtm1i3kVBUzHJQ7lgekhYBDxbTDJ/UBiuvl5ZcNYTYb0sWu0PhkO30R9
HMAyteLSCzNQHnAtZ+GtQeA0/FPZdghdQCZ9zv2P6+R8ZI8DQCf4rTRgozAtYstNggp9mm8D2Ex9
cDSLT8/vdCe7n+Dl1kZwr+MSMsJhQexqNky0w5CNpVlD/0HHK2SA67QnHztfl2SfMj4vi24yaeJC
ztazd6YqkXMpnT7uHxtjyo9D/djwKtoEjywfmInqfQd9ZK1ByzaY9CxW3oB/4qhAwD+sZkXMg+qO
qlX1sOJlRI0Ffm1Cm+lRr9CJe/X0vRQae/MWe2HbDZ8w7+N/eOzaR8B6d8fxoWJKf8JH4oAbR0t7
4+XP4p0OIYhJ6HCX6QtLpFPAbsibk7D7nvN/Vv0wFdV2Lp1Ier6IhrjtbS8m+Iu6SvDWQtR66UYp
pYqYOf+YrVFwDpj0FiexLiB7e+9j66FPuwxrj+QAqKv6zJ/To1Bp/a4RIPJUYd76sH9Mu3zE3SH/
E2SxVPWAuU6aEmF0jU/U2whtncbGeHY29J+C6STuTAmz17XOMUySYj4j0L5ihUYoRcn/0bj882Ou
V1wQ5yP+dD5uJ1V3YOpHgvMHCY8ZQEOlBsngFZ/QfQj6ZuG2c2iHDKR8klCRrmoJ4VGyMI0rDCdS
RRQH6y3HIIwSn/WO4yKpl/E052ml4XmvQPxVtYqAw0jpGNXtIMbAkyvMFHUqZSpGxh3zhacz4grX
F9IkPPUzhY31JZr8/iMDdKKigmC+ctbh4ee10ETR3QpnoojMhBVb5MRm62jY8HV1Rdb4TLCCjgYf
8K7ZQ0SPJ5/FVwRW00cnWu1r3qOXEOJeVxYeIbAe9LAG4PCiWd2Rr+bV2dZIRUj5CVmEMUpnVN1L
e7CVpfFduXoB0fNdiORI6FoZk/pBxXR16e/3UV6Rjpog5QyfD3fA9AhK2lVpqxpu8rqSZecymtvq
R+BZxG2CqxHhYcKEy1OSdEYBC5H0DoaMehqfEffUhAKRqxkdNUGhSzcGI1AsowNeMrzr110VjLth
m4ZtFE2GChZyk/NPGV5HNyWiLTkfdArktd9FjQc5DJL8JlBlH/9wRkMN6DQZ50FsytJcQgDAKQBP
dNEAyq0le5swFLAvW7zRGi1/bTgKMp48607XpIsNoTHZOmdIQKMkC5mV1HpZCIP4HkyeNtObCTEt
vevmEudgn/Q0pYP0XqRTHCmy3uE4kAslYdTAr4wsIL/qP69FrTJJJpo+4kmKiAb2ezRC9wybZ9tn
ugmyeRJiUC5dC/Yf7K9Egn6MScdfPFZeY/XLGLtc87wDpn7rHXrudp6iFqPhOh9Q8SfrWRvH6+Lm
+GE5ID+HgLZ/0rWdYqyZBee6291ClQd5D21TJsP9z0MKqKe2ocRKiqudjZr+B/hRKr59+alVGpjE
19czgcnFHN1kz5pwmhruBpeiz4pNMXl4a7EIWIk2xTG+ma/EnlXQtZ17mpm7+HEFxvbUrxRH9cK5
K6RBemU2GDzHieKrZUXOFDZLSGQobPV2LZPTuh18JVWDyOITrTq+OfEiB5lbTkXtYcBgUdWOmXQg
HAvBNKamTVtAPNDPV80kx2D/ObuBsvY1eXaYoV7k2JdbXzSRhPxWWBwxo/OQc7Po91Iu+GCIAO3x
HTwatDLCtjlueg+AFHY8pnfAH7eepv+3wPRvR2VZh1TTC5g14bZdJATPpxtvNy3Df4PpHiyBYXWD
6ZjhNKo6xwIlx8ncMuhdtDYK/d/t2YhXU5rIE8lbfyDEzrQrH8Ffbmzu6+kic5MOSSLokJdd+0Qk
V6co//wVTxW4TiMrnYkGIw4s3zHnhViyXsYrvfDhliQiSrsKocS3+B4XSRM76qr/EHwQNjbfbnY9
7DgXEO+TkUfrwkwyNzHEKdVz88U7ni3Gi4pEM/lhYWHIbLsxP7v5tPt8DczXkJL22GbdHkYHSwPN
HpZ3uy8Phrlq4OuYIbMLOeIzZcz/TCLQuz/C8lphvgo3NoqsdOhK6H8vu1zydphVxF3MNoXG2eLD
jOupcQiPJP8D6iBRjolhio8BMcqMnTCbyqWXgbk8zYCV+HFBHpy9lfBYjITwowLzPveMmKzZZfLe
JYXv2A0CCX0XZLlYIL63z5Y4lBh9kzsWTtPXpjFRi8rL/kYIu6H+jmOnsDRFz8fdTDE1brjIY2md
9D6I/trgH2CPCxlqgT0erlyEqo9o1n8K8jpeLgJpUVckzNislY0kbMHjc2px7nXwzyNluRb9Mxpt
Xyq1q9HrYEUKZ6KwUG5dcq/XpldyKOdTr8p0N/T9QewLToBDwJqyA/bQMxPWQGMHDFz870v6T78Z
WkUUKW3teJtracwlfGRYI1cekx9sTYzb7m0wyX7FnbDS6dZ3vxwL3ofNIyshUjzaAxOsjzemlzlK
F5BuAMTcu/xBZxf8G4wXmI2PQA/Bx0Unt0tdU7CUFjysd4cLNgSRBe00CBX+N6J0950aYtXtfLXN
7r9VRyQqYEQuxXBpiXYYk8ZbbGzMLNESiq+ZUMJKgsb5JBBUiOg1og+ynv6ZQlZmmjmU5455AbEn
bzFV7yZKgmJ7+yivP7+DsH+XDSpOw2bUCmzKHBZJltqkdX//8jloAQLDFvdyWo3hXbqF48Nye5dc
mJ8vpelNc8jSkDM50Xk4qvEx0euDeSTJFPHB4AAzPDReyUqJ9POQa5I2Uz6VAmT1afVHtBsDb8Ip
e3Ra8BgRrNAb8FEJeQktFa9wSKl4hSEYX9CVGEB6cf9wdmVnpednxCHpi7E9/MPeDqS9Jp9vfoBj
Nks5/Flvcrc+LDCnaToCwLSo3z/zJQGwsYPDz6TqOjoqGyRtWWScbseNtA9cIcqL4AKoKL9A6kPz
bb2CQFkMGYENkPQ84ngOuJ0csQJs3Aw7AlW15lJBNgB3eyytycijFTsL6MiwCEQwECdsENctw82R
dtXVMjzNNWihzYiBK2Opx959Ur5qCU3COG2OYuNbYj0ddwiByHGxoej3hlIn6PdUS/LhnBcg6wnB
dj2RzGYHJZZ1/PDLd29OERp+mwl1dXoGFeZJ2tPjZUnb+Vh7gUvI0zRQJlB2MVXxOHFFM1xlBtZV
drX3pQO6eag2Rthhs3OBcp3QxRYokenYcjK6hd4XZyGcBcHBJIwwzoLF3KYtRldU7XT460scceN3
kF5NLoCbXICUZvpCYZxalCYF5GfgNURUnpCEXVxsy1NUYFHVztKhWeTIPGokCZuVEqnh47AEQu2I
SWh7Jzs+GGLFN3P9xI+giA1KgqNpuQet2ZTpvvBl8vzMZsf0KmDvoJTErpOB6KigtALMs18PBU7w
kujW8kvNVo+ZKZq1QEEcCAo6O8wqCfv7/xqOk2I+5eNtaMV0Ti7F0X4rK3DwjCkdLG+EtPcy2Kp+
CDJOkVCFRnLyoeUV5WdM6QexoHvCSXvIhp5MR6u0EnueTeGtu6UTcEbR06VsI+HswAPbeZ2/XcbX
Gl5G76ODKU0S33wMiKS3tlz7dZueUsgRfT/WbgCIIWA+fDZVnFCNIlTuoGVFdVfYtBvqNQjlezuG
Tqhf53qVwHVP7eyBLboxxPm7MgHk/faSplC733Jf8upSFnzF/kdaamer5Sumhq1sYfBcMEdocGjg
LoyqfYPksvcVO9sL7qYY+YRic+JVeFHor5V/BxdVq9g+JPuGsEkSTgDZuZbX+g2dZgYvNDhcyCYE
7uITihIpQUo3MU3lTdwImAdOZ1I/16FlLUo9W33QIQ7qhERbYVwUWtZdwfdLz9Akx1J8yq83crVJ
WMiAZb4tTet1KBItLtPRoI2J8zgPTlSM7DsB2R5UTEIcyDCiL2jVzaJhODNt5Xl7w97EEQ4WmYMW
E5RvX4j3qeRpfw6i+UbIzNZ1MuU6tdMzf7KPNwJ0Zq4Sz6aqCnpqPcmRJeSSy5xTYgwVsXEcmzm0
bwvG2dhTNnwJUonYCmq1/aE/uYul+cPCSLuDzvPNwrz8CqB1B71//c6w+ZARr8BcMqzU4bgOhQw9
Vy2GT2MvGOWlV3oBgTRTWC20w0kdZwbntZ/1pKHrn4+31vkbsYQis56WBahK0GsShWFOIBVFI9LE
UxFeYkhOA4i0whNIxsdKPqDElqy+Yy1i8M/X/l9+v7hZO8sGMFtxzJWK04zl9SBDdaZ+geRa3HLC
RjXSnKR/jO9Zu2MuMbmjl3FzGFeSWZaSZBBUSnoxi2pZD/8RwrLpjTsw2GtD73Z/BlBWRx9oNUPU
Kf62BmfBiTqsySP9lWK3CFtVfd8Xm0ms+mOWsjy5jFkEmtxsgoSZcUcwxUKnhUg5bbqh15vqTVP/
lUJnWrGIv+mXjzt3KM+RZs51BLgnPA1u2vFYM7qbZ0bZFawtd/Wgoeg7rgG0scq9EfInfvu2NaaU
ZKr3K2+3N3wy2nxEuTd4BMdTO4Neqpq0nxSbOS2Rz+2x++fa8JDq/EvN4qL2MJkW0cc1tBBIpWM+
4Tz+60wLb0BrtnHy3FcD2cGgXHd/Hyttra3Oz1aqL4aNhN7HE5AMvXL9Rl9lomPEL7UZ8OcWGe4k
6GYDHjKFjep8ZVmBKDVNOSPRMZdAPSGnmJcPuLjxg+c1nRtCBlV4cSVGQh+Eku89RNfMtcyxeG2D
QaxNsBot11eLfUZztoWHrcyTgUgKPqOZOdwjtltsoB6qCVI5TvqI/66iy97o6OiRH8obYpykCMsc
XQqdppsVQgoNB8eA2Xvgl3Ic/dvtU3aK9jBugRf5U/F40PjtWmNoVQpK52nbmLq8ESvjXPDLuG+6
ZuMWqb3aPH2flziDnWg5hJzSB0lH+X9SD03y0es3PtPcOkxCT3mkERmXU1PD5wUgO4dArWmvgOPa
Dmoz9bYVdeG6XpvGT0K+2BeDUw5ynVcuke9Bje4tZf8Qwcj8R4v+RQzCKjnMagnGmfFuz5BM/U1q
HxCyEWqPSmzBSIZn+C9HZqjgldS1VMpC2BnC7KbxcEZ6YTiTEuXuicJjEXD1PHJaJJGym5ySb0F1
1iU6xent8P6+yE8mmG4lIaGqyl+YuQYSs9SNlu3AhCBhdCn6hVSmjKOxzsCdk9cCMftEnBlYWu9z
dasgTlVyQDz1Ve9+aYvhwl6gpKSX6Vc/0sw48tbqTant4/CiszDc1Bu5Hqk8p9vD9rjAHm5iCP7p
8uZ0aXzQ4RlbBUM09X5wkiNqXTMSwc3yCKRwzGFStOmjyCg5RRixqJqC07Wg5Nh4+3YWZayVVUpz
3f5fmBqDPG0CGV87xuFOeGP2rXlVk/1z4XYb6zvZFPTXYz9oOHJc3I3XkiFlCEWu+prwfJwfUGqK
0POJsxuBQg3H/dMh2ugCpptfC3w7pTHJHN+58O/FyKLHj5dPtoZT/NCUb2s/Xnum1oXNmq91Z4kt
Fp05QL2XZH6Ka4tPQdAFFDSbkUQsLmq/qw1nLFsjXRSl0Vp7zCn/9NcMGMRskDQmKGuPEjX9nkWG
ge/azNUR5EcKWoFZIXhQl3f6hULq0QfFXYqpNlrOdrlvq/+W1Kzx/q7YClagEZlPFZ14MQBuurqZ
vav4reYkFKaXkCYvp52HKMLdtY8SakseA/WeguCidieXyy1dvq9Kqwow8xtmCCVfJf0SRXLlRHmK
SWrzpZY5cQOPtlx9KIFHJKJ4Gq7PkofeDWthZhQoZGLONhy1i/hr2vtpj9sjO4ZyERbdkyBSxN4L
IbB2WcMhxkY+Ba44+syflXNjdKqwiPcKebmQevbnmr+iq4Y4H/BYIfbUDiRtxya1KYgsj4HGZm/a
/N0n2Ov7+mqurFrG7LH4HkCAH8wDOV7Zl/Zh8ZnsmUBBqJARRhdV648QbfRHjU+mSczJvytp9+h+
tldvMjkSojBOHNnqy45cYBDw51eVyGXLd4DmtkrcsbVoKe36PW5xVnaJDfqJDEY2OeCLskQWZbIf
4JMzUrJd+IMA4BZrTP5JoVkbDcmgGBnsSNurl4R2sL9KsvPIURAleqMj3G/ojb6FkxLNvBJTtERO
eQrxBtgHkOaUqKDh+fH2cOdPYRenxyRDAh6ISGmyNeP4ClmR+p5IiCKt6bA/4Vs5BEfb03Hsr+Qp
7jpuDoQD5gwg6B+Og9mdvLPnSj0VG9KZBAk9ey54RGtHW39AYoKfdF34QjJRuwMVC328mP8C5qOS
Uj/9XLzHnPz0Wsy/NHYCu/bE0sixtFvyN4U0mjIC5kosbyeX3XmIL4zBKxvE01oHVlPqGkwUn9Ms
U6gPoyot++77dj9vE1Dvq2Lb7IdcfNBBpKcFaDywSrY97pTuF3Yucf3sXNtCljMDj98Iy7qjmNJP
7xV3nd+qxoSCX3MT72milokIc0Gcj4wodjug4pHpTF5B67e/zrsIIUn/+P3ei262CFTRW17a0gcJ
q2IOIDeW1IjN1AR0+QfIFKMqcY/HCETuvUc2BfAz+zSQxVaHvBs6U05NdPkjv0FxanduCahnz8XR
RbYi9WsWpvkk+5LwO8G9ipiiNPbyl4VvtKsjQ2JmmI/hso2Bo22wRHjiA2PVswVkcutl6PEEN+jU
9g8fUMocyTK46MkVWt6Ui/aDbFwKUA4yV4KsPjtSJooxjp22csglChYQ2WGUPHiKNo3mn+ztHFCW
b1Y2J2ki++YadtSioN1nGvb9fJGQvRUWk/qTdRVs+1p7mToa5qp0MagXgxF6SP+711eA7h3f+Bpq
GnHePSTTX31DsICL2M8ikYHGzDTYgTpa9IODWPdzf19Q2S3f20cM9gNMxu0KRhZuDBfUllK7DQsi
9WStd3LdrnHjEatLKrSRT+wlWCDTHhu0cqfSYbEqyDgUc7S+u9WvpqcLkiDLFR9QQO2hHMXZvH0K
WBtIJ7PH1ZmUyRUYKvHXZW9O6rrLl842VhxyqlpIP5QddAAIPnMxukY15owS19r1Agepk8iBF4pJ
QHgGiDoSesoZAHwZJvSC2PQAKweFSkowNIMl18D1fWiGI+CGhOBiRqnUsjDef0VcF1E98kw73W7k
4tnl14wubuE/ZyXWqWVzU8zzWVUcqmr4RCrDSQpWrmTgzR9y9bVYHmDW8Hsl2eDkV62fEJj9T0F4
lE3osPVAgjqL5wYL8ibNBjQfutsMV+Afwx1xI5qeJYTjWSvdjmEFWLI2XntrcOdhWjX5XhP3olQm
D31ZdwaTViJRBZ7u0dnG/53hnTYVPkqG2Gdb9cAeoqYpbAyWhPH/Xt9uTS6EK9Vb6D7+kzi9rIe0
ZeQdoLSE7+UzRsikloLG952rpGUqTN0gVLBfPjjs2DTe0P+4sST+hs077WSDMpVVOV99fssuBJND
rqeS/37H8ef4GM/gSHYW5Rmdf7PUnFGcrDfIQ6GCwpyx4ciYaQioLvUHR1ePuwVE4IMH9AQNCKwx
UpG6PispFCbpkN2euPVLwQKnYV+xUrs9A92gtnYyr0fzQUHOl/Ez14+Bl3S/mz3d3iBuH/yrlJtg
Q/r6yIqCgyJjqKsDcvsbkAO4qEmxGrOXM+xty0VVoXODeI99Nw4DqUk0TdYveP3GZSaOUb3CDlsm
985p2C3uhFIf0mxzjVrUy984zGnYaUZ/3RX2DFONcTeBbsyzSjQsd4Kr/sd8UrNHWM58mCh6PEKy
JCk7xo1o0VG4s8DPTcFxnFPf/616irU21wWaCW551eRblOJCDiLOQhWeUpDt9xAPX8S8arhYHekq
OHdmZMN8bZlH7ao2FEb+d5ZhDtEP7/7FA3iXzPc3pPxxv8jxcEyJ5zeoIhbnpo4wjUX0oC4SSTPV
Bb26C6v/bp1MWnZXnBoT6dRTL1Wbcjyl/FWuiZESmvqo9T6AFapLJHHpVXa8hE38vwz5EJQRwI94
L2coH8K1hTjr7WitOr3tKP43kX2cIvF4u/TWZbBHgfe+6zoxB+GHRN9PjeRgDWaAkOQHxyyjFKcB
SAavtBzAYQ/yYDcGDkMXJqfytELp5IeFNSh61FKQC82dJKs7IwiWVWea436QI/J0t2/fQS7AONb+
s/O+0m7BNPGr/POwhtu3Gz+K2RaT9b85GORZeTmYtqMWKwI/SrtAmIkeKBN5O5ODomW9QKRUS/Il
iAq537tiww2lvxhVkt3f7PbEmq0z1fGIR4mD3ajt5G8jm/dWeEIkJ9jkj1ZXsTAB5T9iXWsDJM/5
65uQ8CbNbuUmwdpDEjrNSr3RmJRfwOHo8pcg2NRRcO6nhu58VkSEOcNsTrHE7fk4tvLDzKzA/uKq
08PClufE7fwdAfQut4vtjIIL+7MIoc1jvI6HVj/sglChEwsrTaPpiTnAvvU08X+6RiodzHHL+xMb
39FC7owXeguHpmLDcn1eNAm8UNNaL/eKwCBsxqQNW1BBjCRaRWpS33scPUZiXXGj3uLKbK7X8Owa
W0RmFRwLB+xDv9y0T6GtO3eItg6PjjV/zb54/Ibf2aNUq3mOjcgUcRG3YKe17pcO5uhsX3uq3Rle
or1f18lpj7FFOgpTFAFyEGvs2y/FU4QCVgGSSA0IlkFYw2TkeziGSGAsDpZtND8BfZmvvqsxr/L6
9Ej2D6T+fbAoUR2tNBuH90LHfOIfIovFjdJ5U5Fnjx4csHWNnybQytqPwcSrEgzL8aLw94QCExKn
J18VGWEUtGZ92jJ+FsXnYJs+d4K8l0MwjNl+RIc7DhqzOsUGWacj156KF480kXIIDrAD7UG0YhD7
d8TK0uiARmS0fZoxFsc/lD27HSg4SdYxtjDjunidELSC1uH63ODhj/7A8SJpb58AoI1IvF99RbeN
zoD/zA3aBxjYmReu/AkNoAOAAkZgAwgIJePulB4E+DcB9bGAOqUPab8hcv5KZamDleG2ZFy5lNfo
oMLhMBbJ6d6K8bh1v64QzS6toQZ/xnLOEPLmTPDEu6rlsg12uH1joZQJVKQ6QhpTxfKUOzkpr3YU
tuhvVCCysgxluyU72nX8QfjVjEy1m3LIgKjH/uKhZzabeoiS7hA+eCzNqdngTaQ6AslGA38Lzsg0
skWuN/f2DoR6HNUUPLM3xQTs0ZT2/DdZaeqyIl8RjEF1eXAqdIwh9waDx7oluqotqLC0RrrYoHAb
bpmk3fYi0gAdXMehllgMeS9k+O0LKgucbpvtLyW4Jk21NpeyGvfVox+ngDNkhGWpdy+z3v8MyHxx
i6KEIBzda0fiHegeyiWjPyKNVt/OPAJeK+xk/W7J42fQaiSCa1GcBDNBZpH8ilxuXcJMnFdE53c3
hjkWbqsXFYfXCDjksdVKVM0OPPWCe2aY5G6qslxQiC3gOeunSAXuvcUthVIhSmtcL3ad9YPUBvti
vDXwWRJD34Zo2rZClDw6tQ6ku4La4Gb9w99clrH/64oki2EEdhUHI5LHKg1fqshpaUENAZB5k5wW
XUfpaQM1jd2F8sJQBYRZQLqVazFLmwY/EQ/moLyJHL26PLqtTd0yS9repmmSq4McvRnieXi1HgoU
XtUHTfYGwvUToxORZTbu9ODNuAaeXfkjCNeQZBLWvXMdv+wbDnC4nm2ekq8K7+eDypUKdpdWCfTD
2aglTfFA4XDitWueaLwT+f+GxcCfO8NFDjilW1tA3P8E5pOkcLJP4rT0Em8vCJAsRk83ouFFgFtF
NIyukEj34428AHSO9BKNez3QJ8iuIaC1p2qiizFuUeiakkmC1DRfbL0PBay8oJHv207SVl6FBc24
JG/ojYs5c9sepog6eGHMh/uiKw02NRGJe/DuTyJeHiHg004ajAoLB3cuDutlfGq/MbHcaM6JZ3Rj
hUZ4/QIxApwcxJfLW3TbuWkc0C6Pjqtu6jNuqc4ZTfBWcLcSGrOLGs/eummCnO6C6LPcLspjmGDx
UaC1Q0SC8ccGvSxJKBtVkP/WbzZC3f4bYdr7WgCz5mfaWAE0K0+4FggbJsFanjG2dizlSgn61cua
YOY0ievmH12vWIckHUhL+BUFUl7VWoXp0G+Om8ELz1WuxDlaaTNb6iuWkdVnSxXIC490+Jst6pyQ
ig20pM165b/Cg7KIbply+6wdemW4Z2NJ2125KachTV5eLkP2WlYEslINpbqv16XjvxzMOjDjlma/
pk8IjxvbhN+kVUstv9dZluY5LcKz2uH2wQ8ZPLQzFUzOSXJLBfXb0bhfB+d9zs7g4KjO5EJx6oF1
ParLzzKINcEGf1TGvrpHyao2hAOEBalAiciwL0NZvW+qZ4fxwpQn0X8b6RP4Rc5QLg6jO4JztXgU
1GrOHtjlUfMrmmgq3Xm98X7dzGh5Z77oFmaaHQL45sUHDryy1LTLVN2yVgf/hIWvj4yyPGuw/x6g
2pKvJMHGoNsnD9jtRFlycZ3U1L3zKzr/bv9kdEwe1dpc2g7CcJUhp/OwNowdK0HWwZK/qxeCX07p
HQeYj8AC+VEk9FAhKy48PZ28EYKR8hvnFfxZC3Bgi5HN+M3WyOHgBzYyshW4BgIhvMRjq8CpkfoL
P9JSxOYxAWUH7c5dprZjawt4akOHOGUW1MdTuq3t9UbrjZGNZ+z7twLslSo2LTC2Ue2LWJkhwcv1
EUT+vffUQpYfkDpmeAhmHgH6desxO9jA8PJCkLN6qt1KkoN6I/NeLectyPmhQath5Gk3+jdkgLqv
7bU7ay8upDloczGMQDFF8MjoXJzxoHaSDNK9iBaKvVBp7GFpaYPEjzsxAPn7hhHYL24zseQ4SDEG
Zlnpw0loz9KXZi40KsJp2qbbDb+xuuxcASxYsgKOmdj0zMAtjEBn7z1bNzGpK/Yy/n4hMP2sGNVW
R3w5FvKmlXhFcsDe5r8Up2bEVvigdvOhg1U+5bTi/P94jrpsN8vzPsHpZCPF51gF7tMO5YP0yQyH
UTyi4PmO+5M7eru1zu71zaxEZkuRXQuiOIZUzbdq8NtVjpYKfRNGhFOVtVg8oVsPadVwv/CrryY7
a2nUZy1nfShf93PJPT3R5gmxzJWj5nnV/VxkKy6S+uD7awN5d+4cyDUmbrhhLfeSNWf374jrMUTY
TAh32CLGkaXTTwbsi/kfcdNM8NJHRykCQN3dphfml/xkEdKIdajInyCstBN5MxakuWP1MCcXzgcN
tRGTH0/SMDx8n4SkBS7tzGMijroDXQKE3+GIM+wFDFx1Y3ZKy3TgfBQi1E32vMW2TOmBLN7Dpip5
tnIAMHDBGEJ0TzHrL0bKHrW5MzDdmOXz2FuEH8a45EVHQ+iyGmF6aHHKi9NVjPNKVsCukUcmFYAU
L7PRHxwSsOOPqaeCkFnVa3oOfzRRYZwu+kEh9PEoENwwuXqqkz0P/38lncmnCyDih294NjmrcUlm
ofJWseEud2evfizmfm+a1rUQZ8tlWhW92znS7gJ8MP5dHG/aEQfx8vVaXNWNBEbjNzvkqmuFXjLN
TZWcCUNYRYBnHZTGDJyfE9+2UW8X15MKG82BmN+fq80fSqv//obBYd/fyI6/vTjConRtg5YAX6GU
E7QnQPK4ez3ripFgNI9RujoTnKOm5w5CQf5wxYWr7BCJTLjg48N+9MrmZxapR+iZ/UADTLo4+dYa
gvqA0rO9wddDcq5rqjCDs1uD4uWnetWDw41Vpamy4pIOULNGueAJT+aK+89KnzEZP0CXF7HFsWz3
82qfiMDPbI128XQIheC2e8iFR1MvKV935LQdYnbrqsLBwinDBUrYMzVK3SkanDJ/Sr22SjYDg+A0
n2WfsaXwvDp0/T5hwRLRjHTvdzTRw5h33GkQn0OyOvNh5ptcilp854v7BUuhN82bx68nVcENp7IK
q+ZXTHvqZjFnQZUmxowbCManlj/dC8W/CoJmjmfIMnSeC5zO+Hllz5wXdK5Bn/d2fiS169Yem8ae
2/5yenDHBfY7b8cJ/bOGWBzcD94sG2faqNp+s2kuugtTArbvKlU9CfgljzvIInDdJ/Bxb9ZTetBj
iD7+1TVHQxCLYUhPSSHzqX7pLgqUSFjJtpY9wANcwyKlGUjz9ZKOkWvJdht/jgcrUVDB91MjrTzp
0DQGoQnbV24o+oM08P+XgRhO5I4TVE+ebs7Xo2C/rzCY0PUiFNzchr3FRCAEqo5X+TgqBSpTtTer
+f46TEhigO4gq7Fo4MiKVFeoVFlDqI7UmFRP7hnXzOMxPTZ0+3CmsA74XiG9+PoufDh2P1q/INW3
2fkQJuOjosJ7VS5VUbETU7Tqz0qqIysWGp8XxXZ0814oyqIX3eN5ux6QiyRVp7guoSjQ9MuZu6dI
A8MDGAniOzYIx0vK/ck+4DVBLNp3lG/KBk+iO0RBkPsRje68tkK1ReW73c8vEJKOo301coeft+31
3yvVueDPVBQZXNfJ4qxynn0QEqZIZ7HozMgnhdNSKV5J+LoXXLb3spbDKJHQK+atKIRYB1ON2CL3
zx/BQwJxj3589NM1EOVbL3mxtslzOTdwKFt72p2xqYWrSkWPg8w8InS3bGSbkvPMHRbu/3H3YUew
klLLdwnkbJnY1gN4QUoeidSbTGAyLXTOhVEkGPd3DFnZ21PwsjjhVBl91sv/9l4x6CAHXYvXKi+b
gHIaQMhnsgJ1v4qVpASJAvfydv+JflP7E66sSlffhKPD/rSNZMgfe1Qw8u5YBN6zWPUu8OWAaZOF
ZMFdOazNFo+O5wdcEIBduH0PlusI0lLnJx97GYlbeolqcFEiFqrZAsFE/BEv1KhlRUpJjAqFQw70
WNxTWRCdFu1XFO8nHxZuzfj4CpTfcSgUrUY21R+bADslJ6gjGiRb/Fku1SygZaR4NFRmkkJYWBxb
uJFfQ9MWrokZvIHjmSUaC8olORK0Saz7pRwhjJSbaL5OhhTbXfZdt5V9YruXnd1vABbQ2kU0Vt1q
6XIQrk0OIHTEaDiFg8bJ48pj7ZF1W2gMYO251Hp7/YCW7Hp5coB0dIT/xES7WbdXAmGa7g2ihYek
zMMzAwpN1UT+GEXmO5pkNcEShDDMnT7Smm4YF7px5Z37KLv33PbBYxYLl2ocstzCW24ktlA2ckCQ
OcWCxEhQUdi11l1pNu7HlV8TXpeyvFyw/Sv+cuhactlu7FM/rqGi2V/fXAOGX0cQ3av3INdZsrnx
E7gPQsnqE3es8Nc9agPBCoob/ib8sEx7BLhsQ9vS1IDs9yZ2faBktPt9m5xT8cTy/Mw814BhvHqF
LRcehQLyphbYlvSNIdtkoqeUljJqTqF2jnQ8mXvB5oyJXkzg3qRI54x/2gL9LwvlyqGmu59rp7Xe
8LMvV80jv/TCPTQ+KGusgd+ABiccRbg73WxHBu/LJWRmLeX8QJ/RTSrP8ohHN5yV6LhoAu2vsDCA
px47x29rpB7IudvxRzV6w0wB3FHzME5DezQrkEcKzIf2KYYUi6WhgwxqjTzKev+7rhwTWWqzrMhk
zapG2TTOdHOJSM/xa4WnpdMNCZULiFGA/7y+FI/1YF+zIYLQWS914JiAsiMkHi6nIriRDAhFSrSj
JITCe12KQ7Yt0IVrCnLwD028Vz/4FSst37wc7uMTokOMo+j7ewzRCGlM7VF0P1EXRyJ9aVo1qBMJ
uzPteMymfREzxsUPMW9h/7FY2cpae9hYVcWTGf6l4VWdlKUSEVu1aQxWLRzLzhRtu9yHWMAFLXKV
DbnuLIWh2bKCihEujzdyopxENJ9aQYXYV7WHiIg08K/gz3iazICl335hflPde0hpJ0RFM6XZRGUe
mdGPyDmLxYBtl5IT++Or3wyKdpCBQaiIgtDobOoY9ZbshQ42i2/ZjraBpLLpcr8JJseCmveVxEvu
0Q/9XWi2yUpG0VCmU2saUzDCV0vMP6MRAEbU7nWr6oBN9rK7jFzOXK8MjCSWV3pUmXwwSk5LHOwY
j3vDfHnFchX4/pLa7mQiEfkGlS6xIzuu0I472fu2+Tx0m2RMNVLVQhmgyUpnQL4c7XB0UKiPhOCQ
3Vp6MiP58Po/lTcwu3sF3njjzxYq8P0165rgw8zB4VNSbzu8KGUC5WaI7ma4vdw7qag7fXaEwZ8w
iOUtzDMEHcmpolt+S9jGKqX4aKsDWt9iM14VscX/gyDY2Ww7RPVhUldseArKGEFMBeCpHzRmwqxq
jOtQthMgnaJqPoEH+yeWKcLq38EXqGJXWHhTZJ7ox2IzBwsv2y1tsyPuJEB6VLO63DDQGvWa0Nqq
u5ahpnLIsv2vF+YPGkpghGDRAO56ZOxjB2GiUBZaeKPC7YxUdxv+uQfPHqP7Zp0fccFZx7E4S222
VqG++Jni8UT/5TuKbGxaC7/TY7+COfsKvZqiQFC4e7kXyZ4d+iBeXeopW1JcadkenaQ/cgPLwSSj
RXp2osNC7yHOjrXPChK8agY7cRGhVMJZCk7zX8XAQGzJEUGhDmhQryX/2+gWa3eXv+wFYkFMEoTw
f/p/3xjH6CLHaVI5QlP2W7Y9vGOsrZekm8ih4b67Hp0XrDm87k27IKtReUre2LCfDY9OBoDMfC3T
5ypkJhZ09uCxQGdu1hNPU2RVcgw/oQlTog6Fecg+5FAd0H96Bqylep2ifLsDHh+q1n6af+8c7kKx
t3kaK35RJSE0u+2Jf6hGZrFzloBPnMS0SOMOo+zT1pWmoyUV6rm394SioFhci0R0NzfEOIPPM81y
gt8o5tXOAxm4StT5b42cXUxXRpgEPcPUJY2GB65W/FMUctRv2kuKMYr08hzkVW141Jn5SvkB0pn3
4X3jfA0gx3ngEcDvgdIEqo/2k6R+NH+REJmYvOiMpZcKFk+bckNbywQOtxhtMJP823L26YOwPi6i
+qkIDYZWLifTwtvFrCM5tZ7T7lK1NKVpxdYf9qdjWvixQFXxc65I5VEW1UDYEB6A7UlHdjeFIo7H
XDJhsfZbA5B3haGuYVHDRfJ82nXUr32yx60qXuj/4/Tw1kkdByqMqynkB5BskiTUJH8Uzknprc8K
umtWrEoDmGxMviTn9rpRRxok5fkjL0Yis21zzjgVnGeGt6AoXB1I9o14IPFmFF1vlhuDpap4QU/h
tbZcSUyKbRYbOXo3oqRrYawcyNo/iZliv17sS9Cy/5sYo8eBmiJBxyJD8v/h1zqlHEVGBz4UXx0E
oIAatxMJdKxbMsBN5U8P8v0T53hLgys7YpnRXmHLOzeHE+EE3np+T0/RMaTJsQ9O6DG0VXcoHgYR
V8QHDIDAtSuiMcQVIqj29ELhxoI827ux/Xud0MIRkP9UKippE6gp/shpInNngW+dzapmHKZ/DtV9
2WeL1vPH4SuI5VVsdHOVqCvhdqxNpV+E8dWEZPT2x6qncbR7NDuo/CcLGV0knCbjk7q+DReYwR9C
Q/1trmg3CzRdUZwP3skO+6CRctwXQjND+3ovv32bvfdGqXCI7tK5q4+5L+SKOZv0U6UrAwhylqTv
AFvGQG16judzcKS9hka4TLiYAr1iFntwJVGm2RIIC940uTjV3jI0Hf0/+nxSM92j42Kp37olgHkM
1aJNF8ISiz2RfePLKXXQ77Mz/QxjmxLIUBF7TAmkHjAbeheJlfX1EWfoOi5ls4jHgWho9H9cxJfq
Rc/5v84zk5aU533fVHZJ+uIPZwi0V4HGiDMyyeN9MHzCfzMnYIsNaK0WIbuZNNkJTVnNZEe8LpfX
VseNagbw7JVhxmlh+NQPNVg05VovMPHv+JWXGA1KF/uWDZvijGm+PNi6PmQ6MdlRbDF8SSU7oqJ9
I+XL/J3Oa/9+d0WdD08DWjAbfWGHv2kMLu0s9ScGiVz+lcOYl2J6Enkg5kKofG+Hk+GoOcPTAnnQ
MwDdliUlDccJetp++qQridgqOhA7w4FE1SOrHGc/WPhKHzEShN8ko3w0w2sIKEx6Uo4EMjssMlsc
pFdP16Lr6mg4NL1W3cU17rfry+3RdZDBVIPRw1+KstDt3vp4lt8CDsy46S4ZJ+bCA1tiYb6bIb0A
Go6QiPv7Cqzf3q1VzAt8FAvyTPeNDa+f6Epviw2gMHOehPy3lTPmgVW2TKrfEh5XnR2Nl76fvA9f
sRPVGzFeCGvBtUGJ0zATADtbQ27sWw0lQ83iQtWzPNgT0vf6K6IDq9w/PrTRiL/tpE7vNC+8xxvj
KT4f19a2bLt4zZO+eyXrUx4Odnu5hBaxESedhC6pINzgIJnR0YuoJRjgYMf/if4i64y23mhPFArc
jjmiChnhEtJbYI6NzAYU4t0b8uZYrm6W4uKbPhXGkQOQyHTHMjYBUNRQw2lrouCQn7yld69RBv2u
+1UKACGKiGnj9CzZa6jK1y40OzGGvttUXE1YUMta55xJKWEZJXG0fxwrDsg0IFrKvNZnWM9qzwO+
kckE5QsntQ+mAs13Mp4aqbQFCayOonSLwawV6Vwzsav6UhPzpeM+LPwdZ9AQloLpUML69YURKw1w
oA9iqZ5QrnYGADQtUTqWcOhMoH7zpqUVuE4KsEm6vQJI/f24bRWeB8itJynKlyfPtBcJHb8RIbm8
6PKY2RP0OHsO08jdfx66PJRST1a62D6yMbJCoWJDn7pw9Ska+FgNrCoQCdw+/FhMJoLFDSPZiytg
pu6oa6Oohcqyz5n3ChDdh5F757R1Kmu6VEDcy9rpmImnFo4qf0RZSZ7UcIdbmW6NGv4OFbrhHB1R
Xh3QyXL6f7jvYfYeKVumiNxmXsyOmDPHkJPqYtpkjm9UHwhilI0cSKJEcpLrQ73G4jirltS2czfZ
czsrEcC8oLe+FhKMVBojkZ2mEohM68GHby6WOZJzrTKI22w5Zi7EyvBuvxXDWOjri5UzNaHDWbVw
+hNhmL6pQy3uuuzUHBasxodmYf2Una10k+lyryTbfcPsIVIkId2D2yLg8dX/nfovexj1HlA44wQM
lTPmHrVEBm8qreLhlyaDKbzVl/m9Ei3Jks5780a0PRWU8oEtKheT4c2lxTdU/ub4sJ8R61yEQWGH
aOY1iwpL07GskdvcytKpwdPBQTRtP6Myj/VSnW8uIYm13oBSw5y6oRDzTwlMbJ7RSOt1LuV2RxfY
UQGGAmhj2ZTskRFq3kcGMUPWXxjPRhL+PW72unWCPzYSX2H7SHUFM/yRfCu7C5A42ZfTTlNyjD8T
D3Sf1AHZlD2DfwynGZ9hNiDSvlmUqFT6uUtmTfFRgjNXGzga6KV1/7zzkjs1ZCG6F5Psw44jHHj5
cQIfQZ3KklBfhzLO9kZt2UgIZOOROowBakWwsCaa0XObo8VH1fouW/C+crTlyzUuXfjTMvTqsr/p
uhTGIEEsh8c7dtmp6W2ORSUyUrxWkfcaicXkxttPnOX14crE6ca1esItE+teRDjiGZaG7gzBN1x2
usFmhYJ4yvPqkJyNPDDXUxsw2Urd8OeXEZM/xhNQO90qEmog7O/aT5PNVaphXcvbkpkgt6L5xhFg
P9veL9DhcHB7f1/yKdomMibI3P1zPlInACqMGDTYzlufqzOKw+ySPhORBfitwUXAUj7RXZEXdFCm
RyKe61puMcX68qNLvFbz2aZwraumnM41NlJhW0AobVNSh8cxoCvkonglLXBisFJLe4KYI9Z/mgIn
UdMJ76mCmxS42KPREZ7D1ErJ/ocDoZNDERWIvG0vSRGnG9YEj7upCUOjJ2/sO8sVvrw+QASFpIwL
eh9tyZgiBHY0cwtzZI1occ1q67MPMgGHWOV0U8vInFkCvjF0frEcydd6yWz+/jNTf8bKNiCBGERc
pt7aaefUCAZwZ9dhXFWP+ej/c7jpVhPpmvIkRKGsilZPKj9TFM0R7ih+/7Ob3/EaO0aLhfqpAZcd
IsOzb0BM+2RJL+APaMsMH6L/DbNo6JfbVp7RTHdlsGzQoa3IrtJkAyawcEgCD4hepDVtfs3lNAPk
WgDMAE5DsRt6JHUxOA2SSdTm0GfKJCgiaWSeXxLM7aFSXTzRby5z2IVEImVpcB2UY2tMpwbOHtZG
IcsHkxSf3CdoU3DkPQCwGMoZj6eXP10Z2lJADk8RoEtZdCkKNaRx7DYMIBAWlQV+sfYVYyaEczwX
IosnShqDc7Mcc01xv/XlLLzRj3FKxOyoQnry8NFwQNlbk0IWiUlTnkURuEPuUDwXK6hPBiE5Oret
gxZozjmUiZUYisOQ1hQMDPHhAPaabQES/J7mRHwk6B7RGqxu7vGVwB0+IhvL3U2PYHKqNcIwCBMv
+8qP2wrgyeMwqpCU6L4HgMjt+VEy3cBVUVUghPDwCQnUynTP31MecJ3Sp6Pg5ndp1Rz/CyVYaZ9Z
hEPA4U0FGOg1wAIuc4QaFTf4PN2yn3rLc5ao9MGjL1s0j2Cm+sQhb2Y+2SEbosdpFZ01L2SbNhh7
JcIT2Hyz9ZuEKmUtn8GS3/sp2kFnJNWkRYpT4fJdIAS3pau+tVAPtwpCV2y/bR25gYECTUt/j3Hb
OMxxqGTT5R96NJSITvJezJps4NUzq8UOOXvIrIPrbVECetdhSm8g6j5XmgLy9Jssm87Jg9Tu1seL
GTTjWp9v3i43wU21c/hxBLJ95c0CFuoDbxSwXtm5FuMYPjUFdDpV4uesUo2gRLQnzUjtnOd1WCKd
ftW+7UPDIk2NxzcpCGeHS29w2+l4zVLAuDTzp1sODo2AmFC22zM2izq6FU0DkHSWSh/YbZXZ2x8x
gMUPYy1Y7gwQt734Im9Vf52Hs0kqlIb3PPIXLvYmDSADRlxIHWWXylDD4L0GX3n4VTI4KCmkqtDU
RI3F8RpN7y7nOwNNG5ngaIN9BrpX7V/K9GjkirTUFWRsbf2mV1S4vfIQKLYbg1mgSk4f0D757sGT
h6koQup2Jy8av5m0sfLrGDQbpr5XNevKDXLvNLxJWwmLplki9IAhycKVzx0LT6whdmutDHamGy1E
Rt0SAgbVvbC8IcwiMg89/HDuM48VQpd2X2meMO3prFOsQOUezHXP/eXoWFc6zxZ02Wjq952hY4Aj
v1G5OpV7c20bcjTcKQpB/ARux2iEvNg5ymNTcSrkZ4apc2+prW6McDrZ+qvAj6UdjqYr/m+fsjyA
hySScnB9iJzUXEtdjqSl2rpTLFD9TEn1k4dQhOpaX58mF6j2IB1Cjeqm5TveUU+8hnamVTL4q69L
DJwdqkMnryCywXzKu4FDkIkZKcZTEU3NSKB0Rfo2mvRxIpWs4lu0YsxPHV1HubGp/MF9ozaQDBZL
XLlTjVSc1rMqGow/h2P1C49M5QRRhf5IQUzOm7AjmOTO1PwkoH6A/o5mX4kDpGxHDU5KG+CXLehC
Mfus9gqqSA40JfkTPkobkbg3elFpAztCup0dUBPWk0f8hqxlyHWSNdSGTGWBcbvSz1VHIJYeng78
XiyoeKhArZuOnkdYXlCF+KApFcI5xc8QefTpYxcClT/4mj6VPpGnvKND3OXGdLdymhK70z1Hfvuk
hh9JrJak3+m12omHDFwS4ZGVUIETDptAolKOrvGgdLGDfTnV9pUFsmXH5YHDQB+J5RcGfiEKEA7M
dbn5D/mf4yuJOdFoJWZdw4ztN6OpedYBE2jJIYnUdw9QxkLkXMBbxUILKYK+Y7Op4CyxwXSmxzoi
7Beh6QZ1kAedsuROO/MRiwcUmeFjuJRoQt6SGA6r+I0nT2Nnyi4InrKe+feXspzXzcb8sQaj7s29
HYF569SK/m5J6BMygUtciWhDAJ9zv3cxsAxAawHpLpq6gXDlWZXhHqQX5ityGQQgythfj2nrFIx/
+n2zg9Cw0eaVZD598RiyaJRPPWpq7ygyz6ZLhEL2tROpmSV5elG9grPO0o77bFxa3DH7zlQaAwyU
cpzJ1NvSUtcJFurWI/7rwomkF3aYyVZSgnUeXcVVAkVLqDJYZEgYWJ5tORqDQVJXXjsSJV06QIBs
3wsHlqZIUkeRZcJ7fBsEczcx+CsUE3VykkWqXdlRnrkj6Bl96x89RhZJ6ml16dxgx0dBqHKSxR/k
YSPYKfRgTe7coqAgRKkazSXlLggM9I+rrPKs65dvCM3i+fIq5CrAwIbn5pglH6imTtONzugctkP8
8bvxe+2Ekoofvp+9TqbumAR72qXehhPS5J0cNGoq6AXn7tggdLys3O320WI2wKeXFxHAMzCPL+wj
dO/ibTKiq7rsRJur2SgqTcqA67Ueg6s+9Jafm3dmT4ZArRI6oaifazZqZuoVfi0maLxj1mx4ydgX
fCDPeNxsQfZF7gj9zDDLJ4mLuCQGr/UMVJp7izRLWnVHkDpaZlPi+hap1v1NXutpNF7WJHuZQigG
+FAR4pT+KXThUkVHsCPJxqTOh7aVJAtDCKVJ6RSwbGsOjFisyAxNCkX3YnPj37cupbnqlGSwB+OY
8SKqGyLZ/UIG9ODqGhZQCDDXEkfU7Gu7bs0zjw7p3H+o5YXSfGZcqoVnc8b4pigdfQHBVpYWDsSM
AH/HbAJI5D7/rbMc5FfR7el25aFLOSZyraGjhRTcwy0MwDJWU1DoFOt3UI3RCK782QJsOMYRO663
qIWdm65bQQyKExHoaSvx/VtNPOaxBZTuzEXQy9e1qlubEHNqx2faxkdXoh7FhWzQRottPS+0Kb80
AP8ZXikTAVFFRk9Loc0b5On67F+ANSjdFrDkuWN5rKSIGw7FtiIUvPPJA9hiZptUmTDPNqIwWzEQ
yzhaL23ExckXx82yQLQJvb3jpSmOjemrUjQ/BayGlIe2hAYUnx8OJpYIBR/+u+0M2uU882Q2Yxj2
Ni/zXrro2j9hKT7DR8DxcJc+5sgsA9z5At9vKY6fqoMJcCTsAE6mYAHiZJpaSItHQ5cEdvjQhcJF
0Zv23nyBy/IvxZGx491vf9MAbtvKd0HhIjF6OOelPNZC0MPFBG0FjgD/YrvWaCLffKlDMV86YbGt
/MRPOQB226LuFMEPCwBcdwQG+GIw+dhOKRRYMy1iqc+xjz3M+kpQVOMjYCWUaGgroGZJFMEEcTSr
hcbS5f/ynRwDYRkWAhT6Y5/OQF1Mc93yMWAQkcbGJfBwd7oiHd5yVn+lshM+2UQ8wW18CJ8727R5
eDjkrEWzON3Jie0ku8GMkN52Q20K6blTtF6Oy8Q6KaJN5TJjLQp/q4Ek8M+XbsbW1Smcdsb1PLBs
hfmpd0tgHj2grTbTaGvjUi9P2Uypb6zjegmA0DFMTFmL6vwCisAt7F2dNYXm6dW6MWod9SN6Pjaq
Kblv3qKzCHxv7eeV+nCoNQ0kicyw0QrXg0xMw4QjvaYz7l8Idl/Nh45VJTAGOC6pum8mWFdreqij
c6AfHPYbUYWY6YoNnubBJXlq1vI+Dt8gItKxo4x3uJVrxtoFH9wUdaiyue3iyS0LopIzG5sym6UC
4GBadj4d6myIsp28xdHiVrMbx4eet1DBvP69ykdj0GYKIGewg4Jsgt6MGyZ8tA9fwlJs0bgQskz+
KCmbGb+ie7ENV4anyPRA8LGYeh2SxJTzPilo3eADWqLC4drydRyP2vOlMKnUKGHB4CWaIxd8+MPg
M5de3+QhwfG++mP+TZHoa6XK/VfjWJc21utha8FEMrWbAqBRhVwz1xTBMxgTmdD1VRxTsbXN2UVJ
8sIYnp8Q4FMVHx5cubYO3KeOqaLcV3+vGoFF7T6l7ScCGAVpVrZ2ty47oU0eWG43lUYVdXNscaq2
LHcsCOyy3+ks7aH0pgh1h00+e+DpecOLGwVBoo9A4E/NTbWDjXZWHPqeJmKVhSFqJ7BGYyw9B7qi
VPIWZZYlNhVua93pefeTTshSo/Mh+Z5GUWG22qbwHEAxijGCi8xhCergL0Yxg8FzRpc3S+omKX0V
uqcfKy9E6wOFx1R6aANG5ntqMvSBzj9zwDZSYKyCJpcDGdsMmhX7LGc60a4v+tG1jMNeqs3cDXqJ
mDdxMuBLbf4rMXWImrn2I0wD1BZOGtCdwwo3n5npNj+iVjpkWTYJBxDYzvyg7ykZ9teylLaE1Pbw
vl5ab3q27NqP8B6SQdFIuoMRHQ0PicK84QPPUfW21GbLavMYiGY5UYcQ2m9EvmVB+3FnNpJ8QFuz
oUnElKPjHZdi/54dt5J51ZQ+FMvUqviXWhx2yEyPgbNRPWs2IaezAcZhNX4K2Bn27J24I6jkC44g
Xkm2q6FR+xSd5JgFBRhhXBLWD8A/iW0x23gwr7Z+DoSeqOBI7xRfGhez/pKSKUh+o0lP0cmPgj8v
1QITA1efOBIDMQlSgh6O2EHkaWAI3fYNUjXTDpwgDY4PUBkpgaNnIPliooSoo2MH/LQiSpr/CnUL
TIGsEkePxA3w+ORy+FzO6oh4Oals7u3u9tftGickyDYoDvtn8l5XlfQmKz1J3TsQklyvYP54ZzLe
aC8dTui8VOo4HlSooPMP2WJsCej5FA0/zBC/TROh6epGtyUyR2b4i/v0dM+nguu/UusuUzzhhSL1
uMI8Unhaem/Dn8mk6KGJxu6GIRVu/2ts2Dz9kBLUifnOJC7FlZXZis+XL3OyjnlUQHOMqYbU7gcr
+BxH68Hz/SqhfWY9D60wKo4bYtzgOFg8uT3NnnPf2IdMoncrbjx3/beZy1WG57IEduE4KwTchBSB
GaJhOqwcohQk2r7tIQMm9RoVnIDCinku+6sZyJhE8SGpxwtmibcZHTiErIzu4btNQFfWCdjW406F
W1W3zUNchdA3NAG3k6uYFjndoe4h0hxmWCeraiXI810Ldq+EG6f8J+tH3SuRnu9ZdasXYBPWfA7a
q5u5SN1jWOU5fDN8CP1FG+NMVyiq6TLqrncqu/StjVT2ljXG7YeWBKU0omrbUN0AzmkCPoYZeTLA
zugr81lAunX25z0kH/rObhOlps1aXSNE27mN56fEvKpuv+1F9UC8itgsBgG2WHxPJdEixZcWec7T
0bpkCYUD+094NJfY4UqGmpzWgHcrwJuLHVb15mt7nkQTuXKVf0X/5i9umdTT43rg/qug88oWkRNh
vnRz8GP4KRo5PMA0KCTz6OgruE1UY/k54205MVNt3l6q700YNJ6CNtuVionUIDcQ51Ao1XEB/Zgg
D95nQJ3U4sj7RZiA4/ZBqDZgoQkuRC+/sxG94QMl1oxziehraDCvx/PtHUxB7mbtjVf3Omlb9422
Zngmle+JdRyIHz85ki4G1F50bt3EqjriBoBMEOLlAtFyxx0TFD6QR60CDEigVKlncEtjime3YSoz
nj9tGM0jcmY6a1VaxVT0XvA2EZNVgChlrl47K4cl8E6zgTQbjXizJikJQS7kOzuy04DUKagiFxOt
mR/rs+Sut4bsuCla+AcvzgLL/oJUNj2e53pNx63sAfViz8WdUnMk87te1OI1wO5KjX3dnMp1GpPi
Kh9WhkM0f7wB+RvcyWObcJLL/geXi45qICHRztlqNNAm/xRBY/dDc6NDUkAESjg2ESz669ssicO3
CGOcqpW9HLSPXTwlzbIcj/ihBT3iTbcCOEq2sivVMtlzrYMxxG3JdfYE1ejmWEea4ZQz2YYH7K9P
cFb/Kn3wYWGRElJQpuXi1vDE3pPncjTnEKKTM7gIHkOGTchQ/JY9BcRmJFS534HMgA22znX/xuYR
Oebh1Ow0UawvMj/H45O86L0i9CkiuLf97mUld4XOl2S7yuNTTeLDbn5wqId7XSYMw0oq9HDBeWN5
aq3m4gdbrcuXacLzvlAXw8HFqUOFxVigotbUQa5wbSDaK+2ZjxBtH5f+hGpUd4A2WV7pKCV8pmd+
xUF9eIDErbhrcE/FQIWgOA1E3F6EGX9tffXfXf9ZfasBOaNwsPFjzGyiJreMUxFVjHp4YauW0Uzw
aR+UPvcELX2VdMqaDN05HBX16WKD4ThLv4Xd+7GtI9FH7IZHVu9Pj7ajA9Yoh+QIhCF9/Tns3qwd
uyYxSrRCclo09yUzylTUkQb59ENZbIeLXrUvfo5QLML5xR36LQjwY7LJ/HzH3cRAv8kZOUm0qhlf
I40yVIw1Pgkj+BOAJ5C9IGlzUrDf0l0mo/oWlFwLacDjVjFjUFATzT8MLY3F1P38XIEgly8eL7z/
wlYfBg226i1mdFePj83PMNPS1lpzWk26GCdJuARIB+YtxsQBzp5MhbmoemjhefXwe4ctgflNqBHe
t1LL5mOvlVvuiRbmSZMw/6RsQjsKO41GY48Bh/qzdUBi7s/jBu1B5vqwUhONk3N+DlnEXZ4Rg0G3
X+YblLduo3GgXI7KY5T4wGxFLFRxkxLUYiHwbA6wU6BFsq8apBFhehjOSJCTOtGNRHYdLKx1pRxl
m6vA5VU/23H+HC6AVOzKfx85ttQaAZzbntlDdZtMqEelTjgL1UUCcytEilP/pWZux2NEhVmG4c5v
rfZOaoeZXLTE9h5us0ekhFyGSyTG62ivS4l6MHkDUveZJbVoy0ioxagNm/MIbMmYnGI2Wzh2jII0
fOIUN8VomkVCyl2l93UtD68Z5iC6VonRpZYULP1T+KL1n18e/GLtcISaV46WVKrRM1J+EuO2ifAp
Dn0qCHD09oP6nnQ3zGWbrN/4E0qYrKgVrfqjZcKyXFuyL9d6F86a8Gdd/75uBKIwvQwc2O521t+z
c8qov9/AhPK9Y+PI/iTWO0QX8WxCHSKXOQeDD24Rxrg8+vKJwRUakQeuidQzsTkn1wtjndaNU16U
+ktWRD+ImEHKcc4A7sKLx0BT5eBNQke4TfhAHZXg9/56RZzfLdoHjzpl6P4VDx28nrLDiCGjRu+y
+v/U8c60kLXTK40f/4XNLCNOP3b7N78LRhGVKKGm4dJgdtn9jnzvh7zr/Cq0TIW8I37wrM4d+pUq
Bs6FQFh5Y0RLyh2ceqwM1xPypwh1PDv7YVDZh38u7HvBg5FEBzvmrrEaU7NNhg1mZRt7FLzF/lNf
b8lQBqam4drmvbdR8Q+2U14houT2kBvJ0PO6/PTBuyXpLVEaXo+VBrdvZ20bOT3XCKXZ3xZYGEmS
3zYegIUG20J/TT41aEdhvKkSTsEA/OsjYlGDlaR9bvdoDhICldFhTHHSNrf6SQD//GLilFhOSmMZ
aPF8q6yuy7P1wV+DFIzvpizzflMSU2fQyRKH/vu+aRMjFId9T74LvwpRCX/B8s8vcvLIuS3wZaMw
PF6I4ZaCyZbR8jsZRN/yr0n093Xb/MKDh17OrLPyTFW96MUleoo8PIG9WddkMZZQoHqlBKwYjLju
H398BC4k/LeMmyOnAFZpkA+0mtJlt0GiI9NUzClB3C/vLmvdHtrx+SyYMrUnAvj5ssNDG9nLi0Sf
VydbgHCT2Dx8D/MLHjJAaVeHoDRBd4Ax7TFFUNQ8yPNPfbi4mGs9SMu8fzryEXC4/CcbJMjjNg16
bFMeoNrknlfWAhdNB+ylRqzwnTjBBNRHQaImVc1+AtXEw8hQPdV57PVxKvFnhibtzWmNWkfyK+OW
WAfM6uYkxYD1O96fRG6ChXinIaStEg9nmS0kDr4ao4cZnAdq0/wj1n0bn8Z6YWh+v6UEEmwmzu6Z
w4fkXvQMlF2HN3P5wqWyXAWwtEEuVzkmzQmRvXMZTUCdj6+3GT2Ssivay67dYW8JjzteQ8mn5pms
W40HtNaft54+T2RDhVA1pMOlqI35YV/9gYd8PVPC3NdE+e7f/T5X7w+6pTznC+yfWLcmE2LuEOli
4jSXWTGM8Tw70Jwig4ZwQNbUE/g5Z2APnMWvhzWEpo7eRGMxFlkec+tfzAsqs1GySExgFtvh96U0
BllhwGooLxejcXRP25Q3M38ohTY+M9XCtP9xzNHeGViDp116WmDDBtBRSYUp3rAF0xv6C4KY4J9c
/MnCNjCEG8cy0N7KCKfhAt7evWXY8BYu7ctSZyl7Hpg/qZMnos9BcnU81DafIO7sRxIcAYD5VgWJ
YHyYmzad5S4y8lY3ye/7BDV9kdNufW2U9JAhAC5/zQwOKpDsKuwBmbrUBCqIESuy/yxki1uJPT00
dlDMBrGK3v5nAdw2hnFIis54pwnIpXvMtyfDYOsuFmELdYDMnz28AZhmMSvjFD0D2FEKL72X6vrP
0pB462KJIoZQykNyd7cE6XKrnF07ChylOr5fIFVAueEoijY4kS2SZBff1WVvfyKYBK12dbGDP441
AicpPwqSDAvgyHUe/q9zEbNZprKxScQZqufwIoNeZn4S8wWrB99/4YuTVAXBqqWb1xzfdfP/3DvN
dAiyBlsmIgM86V84j51SZmn+hAc6s1Mvd2iwNENLb0Se9tyM4sVi4tK3PZ415yZiTpKurjiGsnV1
cCGwXe1vTi1VDUq32e35u4wQCIVGWcgwpqGUcTcLuSwr8d+zApK53/hY9oJtkCSzyHlGVAYwqbBt
onb1a7MrVZPBMHk10Af1p5rg1UyXwfXipikp2YJ3ivFYug70SLg6Y4DV10k+Gcs9X9DLsU6RAIqi
n65RhL5uOozky3vfsnKD8Ag1uhn7attFeT5JOmUL0fcn0Dy6vcr7ioKcpJgI7E4LkWZ4ubOrBlAz
Hh8GeeILvxE5zKq2gnoEZmmqlMc3jBUBSAV2QprJeZq9PkF0m1D+VOdgP4ULw3DUSKeENAfrOWPJ
R7ej/oQ5LunDlDYJPemPbsIQiQvSK9Q45CCCCbPCaT/lTfwSpWM27HGQtjUUtcmqLsrtaa+KV1Cw
9JISerlVi38pvvSNWcPX37mNcpRQ24avbvkFqwH5n1qpsgw9ecHjCoFc1bMANNz8BhOPy1omqCls
UlR6yEpuurgF8v2jdFLWdIjuaTHSdLq0/QxXiVWrBR06XqEb4hixe0tCXqd+TnBypkUdVtFXBsyf
cDDtN5O0kVjigJnExPgLVUnx2baoa8euJ68nNqRN1ZeLEeZN6Zqm39zSBLqyhBJsb9c0WaMAZPcN
v/N3zZfjkSh9c6ksuNZgasVyJehDPgDqHt823eCyzMg9/NOEC2vWB9vICjsOCPG3HRWSIvJl5qiL
l8+M7gSdSblkliH+tuaGzcB3bTlYWaSISmO+xlIcjYrBAxMtPhWJFxkDJiwWENNyFSI3/zOmh0pf
B7s8N3u6oFk5T+vVPr/VrKWilXSZm5+P7wmocAixH4D2371lK5VuNEEErhLOx0bcHTJPg6MXTpyt
dpitFku0wV6BbyOtBo3/jTmzTOwmNFMXEycIXh6S8Tz8KKWq3rH5FPkprhl8L9er6zcL/EGk9kBZ
Wb2z5zbiWBdZIY4qUDaDsJTg7Es7CDNQr+Bkv8TbvvQeQlrZoowof0BEBVNwullNVBNQ9cmijE2W
7bJfXggkCEg0Fsrrz/ePZ0fbzJm87wUCCYkAKtdUhdTZL8yfsSjsWri7a5iUlwfl5N7ILH6JYmq/
gODimfbXbLyDkSzxY/NJt4eqkAPpzwQyGjgma2U/5YfjefjKk/kYS17gxRY7i2CqRcUFxmQzx8mg
jEC+5W1RPHSxHHO95VZ8UzeG1PeMP7Zg0NV03qOGBckovCFA+goXsRVyQFZ0GQO+52/0VGy5i6YX
hSDG/8jRbtu8i79tcXDuy950FxLhEyhrlGHceYrnLF9tnB3iNUt3tWZQd4ciAblz/SfCQGHPmxGc
D9LfeHejRcVABKIrY1jSUzqx6lJztxDEJOquhfLn5d+76iFdlkid9y/UtJWY4MosgTDhqJbghPtV
ZT8CaMjH0p/9YzDQ0eupZBv/43P9gDz6Eh87yehvXreyNqE4KVmwMrtMoYkBogXA8l8IPOGfQa8v
xAHh6hoCS/XrUlQBUKUM537NnGvd9j2hmotniBJzjF31HovhkYz7+ypO4XtWGDBqgMwjDC7Nf+Ve
3ogw7Ytg6A0ylex+X2Rn9XK4ysghxTVKMGFJ2Eb3hSuvdd4HCGemX9DqjpKRdb1fjI8M4ML4Z4cb
52Dt6+010dPgzXO7LBNCl6BiwAgOA45DFxEx8GLXiwstKEnMPMlgIAQs1gv3MQPb99870dX4fZYO
DhZyvySFS349+gmE5uXWUHvlV6I3EvFSyoteu5sFKnH2syopatR/d6pPklypmyGAIFsyHTspuJTL
g3skcfscDmP5P7Vm4x1eAdBJvm1bdZQsEhMsyFABTRhTHa+cHXDnVXuBQ2VqxFgblInaooQSEmN0
NWpuZeobgRmdo6BF/41WjQp0XMUIhGZwdo3gNjatpScDG5TPxcAunEzRVREUIwKfI2BaEvCt1p/V
hxgbv9jKcfi0twBsYZmlJ/iICpYabXjO318NfR0VI6y0K3MfLYMGEJkiUYEDaYZG66UJGGH22Zld
C5eAgo8BemdwsRbTuaira34sJE89OCHrsl3tmipwJ/3V10aIhAQfJOQSHkLrCJdq1fmL4GLf1Dqw
/N2eBJ4dWhqJMnL8+BMAgQA4w+dTlGa9O4zxHsRFfjrD68DNG8l5kXC5OSrMT3FV5RhzDgpJ80am
nLHcQw4X5PViI4IiGyOz0DVN7HWbQQ/j1qGIOHlSfXVCH3zMcB/bmkxzDPf2rJU50tAZkzTxt+ht
kgLpwXRo3wBOW9HNhecOIFdodfV7OIDG4bm/8P/xmWMIGykj25lMuCTcq4HBkYQeAq1mVpj/d3pa
tWO49Dw+16G8aoZESA4SNBFj4hA1sM1bODaniGZwbwUsoEv49Xp+LJjhO2fSJVWHY4vb1RLCIvZW
rTCezAa07uZSdhF68gp/nB1s+xlJeplAqLcMspRvD24wYL/ZA0c2erV6c0AitAJa67TVtSz2lC/R
Kf037kpDOokS8XsjrqIJlKEfZKgd/uS51Gp3Z1x2sQI85VY/aIw4gCYoKzgS5Psrlze1276byX0/
k/Jvcl1uztFklImO/auh8yDl5z8G07IKaaenCzCk//hYtuc41lRtoc0GiZNFkHqxjw8m4f/PYnpo
kNRkFWcHOQuM+xRK84rJMP9Us21hGf6zlrV76Dh6z9DZf455+ynMbsr6eScey9Gw2nNHms3LnOAN
y7z98LzVUU1vfVARqnJ9y61fDQop4dr5xf9DdehxHtXrDKzG6J8oqdNBcdgNkierjBIIhtJ2bT/D
UCbZ32GDs1wiVxCBEiOI6YHfX1OWLpY1tRDDvdSH/iKR6Gu3G39Rcijx9YmGddgHqe1upvU/2XXd
HUlxoIxLinYF/gSD2Cxwrs89nF7deEKrwErDo6cYuykE5XSsu6kxyze0IoRUyG7ga55ynVx5c8TN
BLAkHE+Tf0tWERuOx54XXoFfKbsh7xmRHzfG/r2vIfTTezYRuPCrRyOMGJOV90iT+sLKg1FptmFZ
6Ga86n6lZVFQByhaMv55wPQCU71hEipclvFeuQUOp8heRO2QEIUY0r/Qqztud6QSqH+e9P+MPrt+
GcET0EtC8la0sVZt4+UDLnlS/RkBSVAif+Oi9jFDFGxZDWM8BMaRPOK2MYVSezk9tF1AaQGJ+5WD
Hd5fpWKIgjDNDJeeA26WVA1ByDGPWdcL2XouqbPCPzE3XA/BXmXeIbafdU/xQxWLzSbsPt8tKLO+
aevrU4OZq86FFTPse76I2WnWEF1S/ViAwqs7Lk3I6wZbT34IUGSaK0C94TswV09ycn6aa9+g4LGK
c3gVW2HHDzn63CEI6EImwJS7k/hTbOhZTO1pU0O9kMRrzlfAAwEOXNyqn7c5a6gj5JT5kG0DR8ln
OsTWYsHbP4TrzJL/PuIEidMRK47tycfboDcm5zRHFZvG1oKXM6ljh4FSAcCwXQL6t6MS9RotHNMx
KW9iDtIACNzvbGKRZbjEoCnlRJX+dF/dzCbVXpYRsptLvE6DbwMnS25kQuf0FZcQGUgPGHRmXM9Y
LEkb9fNqdhAKUXN0YTuBGWO//2TkMyh2h+DZTqZFJAJAb2gNtvA/wiePgTw2wgifUkctd8iPehaL
ZnptKrk3OVz7V+NqjQ0Y1kS/qmw8L6rta5fmsaUxQ7BqII76+wJRyC5s9H1VSpvejJMi32VLY78D
4uVQgzVsBFnD9Y3Y+89CFaMs5RpOOZKUn3z6sKfqyCyMEffuhOKo4TiKGzQRG3Qja/507G6eSFdg
iC22JaCau6qF88mQeLNQ2yPWKKY79a6bEb0F7J5nyHYJMNcSBvcRIk0y/z7uEWrlrbJMz9EmyowC
KhKoi428P3Yu9+OyCaajyOhG/tF4mMKl4ddxIqW67boVxAIvxWFwoZuz9V/KAdmArhMxEEk9x4/C
VKnBn9P2FfXQWZNrcA4RywlG0DE0fYUo4a4sC4DKI33ikNCNArXVmBevTnxROgwqWb7Jw003Vtyf
ospCcT4YV+x6RGbS5hmNQYa2/vPVSrPoTY6dyZAG0jP1lKqqknU9CzhxC5EQEya0eO2KvxaQz9Zm
J4VVfwLuPe6yPEgqlw2CnkCcqRt5SW83dSumtWuNVTYL8bVyaZzr/VCd9atjIRz0HNXDo2MfDX1R
EHRKT02UdfcM3w239AnfaT1uPQvICBtQK0m36iOaTSjnZMTxcyaFkYxskx2x2XJZpXlnkRgnnmx5
khoQdl3xPDQEF7siOU/3km6htJcQL53muoeriPamiqhXgmCmIGTa88aD6lTbxBN/xKAdaADkOSgI
Wk24gRwX2i/PrL5kUUWFOwVi49kHo8z0dWVIAJo467tbqrdgawxwW+27ZjOqGYOI09h2Wi9Q+h7l
2YC6hfM5KcDLPv/geXExto3jKNB2kAUwY1Di8iFX/gP5HAvQXi5IpKUNZQbFpFjciWc20qh6EAW5
1KlRgNeiggky81NkDjsBxwYW2NoA9aVvTYtzVGWeQe3KjsXK8nR8yRZZMLOkNZY2VqzHAIg253L/
OIl2dvmeKKiZj4YmQsmcapAMDKjO5zIpWEiHxQc60sv8OpupDj9+iTS7S6kfk25wlEvCLSh07d6c
WHLNJ0GawIAiLUXjM8+wT1uBKZL+tpIgQMW7tZl8t5/9G0ZuJ1CLI1cmAJvH5bRBYK/JmX2DbCt2
sOCskZFnPT7T2MjBxtVsI3QVhO1bYZuLth4vVL1+qeWotBPcH1HcNGZE2Qrum39DwEcONlH3SFJ+
QI+Ubsr4aXIfQQ/HYuZYpesSHkRKYCCkwlA99c91c74N8GiSOnqJqL9e3HneqWtqS9i4f8xP8cap
A4LF/Aku+vRgqouzHZGfuhp2LecZcHbQAPwzxVkmJxSi4+otpOfzD6VVxE0wPD0lCvY5/80edF2t
Yo8RAKmqvXooXY5VOMZVjR6g6/Tv1b/Z9wfVsomtbCpsTMbjZnhSOLH1QaOqMBhpRwBFW9h91UDu
F7WIgY4yoS63+e8Hl3d8EZdGR3iMuZBMWkEkQla+2XfcSHJa1Kn2ulVmRSyzHYv2Nuv0IXzwddRv
R/6lZzavhnY5TcfZZOmZN6kUhMg2T3lcLZfah7+LTkDJMAY8uemKQ1tG5j0rheeWZLCR7XRRytHV
3KNveZFDGPGSMFICchx1smk7sqTBJqbu0gODJHpU+yzgArNtPJpsNpw560L9AVW6QTd2bN5wC8e4
GYz4tI5wYpxIevOBduKT9nXKzMoBEKnPr3mPVotpq/20jl/Vi4KI5GpKPAvF48wHLszi9TlkNe0/
UkjCbOEkagptf9baLct911dzZsQtJjoXB2jWjzH5qdDUv5zGdDkf50AZlFuz7zsm12ZrU2tyM68m
cPzrNr3J9N7QerLzG6GpjaeOs+KNSjaw2+VuP/tn+gYPiHNf0V24C6+mkM5Za+a/5maFDvkAlk8i
xUqKkBwzULjWajCeUhXC9LVZvJPXX7T7C7IQJAkXvTrchjxoX3Uug6LB/wMIgjq6BefIPDhDH+N3
sA+9te/xBi5QNkccg5PqYKBRmhD+O+oX5J2aUsHJAXIWhurm7rGRPvDymc8lMHhsJWvvFgwTLL+d
yF6eriiqehjTXzv08jWahjrE/VSUW2qD1pbbn9FREd4jAtL7Z/3wtyLOtXF10JCT3yoL6XOGQkln
1qwg2AdJriv/McuOXcm/uN/+GDDpYxWd9FSqheHnLCv8M7vjlOXCGbFY0EfrXUadkhkcdrocvCB1
JixYL1/2A+Gb6WQqCRbO8KHwvgLFIhMfms50tZyxlBKmnzc6UguIljZcr2n/ek76hxsRHKqHtO2r
adWWH+ALALE88kq0Q7AKStfKT7QNfLXLhROf0RtPYHOCyJIuXc+14eXRZklXPy+uoMt/HWBkV6Uf
+Kc7qYPrbE7GYGkdbqv2Z2F28WxTdPx0JrUXESWmBxUB+mrtIB/8hLT94KfpWAStXmen/VOQcDyX
sTdnlGmog26uW2RQMj46koTOPDQpNDxB/dOqpDz+FHBoaTzEZv/o0QjqkBm5B16Cvs5era+t32Tl
CrtkI+mNVcx7Q8U8+YVy0oEgXnGHNIeMiuf2qjHvVwT4/xmZoqtKtfsJ1OKdu3kv2l0gWanpFoS7
JUprYpR0tonSmBUSbxyfg6BvUeG8xQzpHMGZ17i5mz084P21vwdYD1xjWLaJbtt7JPtB5D/qDJn4
uQ8GTexAice346ViiMYycxkllkocgG/6bh687Kk0mL2htzXF+O+wSHl9Vkk2cogjNgGTVjBakqOs
DYIpi3IbIsHBN4PnhKCAOhbGIYwM4J+yP0TUeMXkHybDhIUt4Dv8qyMUDlfv03SMWKNzOxYMc9w6
MHW71rW9ib4QCM8l4cKM9nt/aw9UXufHJpqSkqlM59dphJduZ4GxvVDIddjIGEC1Sk4HFA1T33hS
tM50k+o99LpULvKy0Tfdr69DA4DMbNwPYlCqmW46QXsepTdsFjv8d+b/AyoZdShdJKvLUZBEz6ng
oZsgdb61jPkmYIdjJRVGLSg+Q+AdnYKIlqWcCub4ViPhew1UaCnRyECuch78o3KsQaR8t3oMiZ9q
GXZvGRYsWiU6DUurkNGGkj1SYiWHtAw9HdR3I3qu9sFv6CdKcG22gqvy+c9shWvbLwMhPz9wKBHp
InNvAgrjsUiQP2n7r2WJnvf0kSoq5BeV5njgP2ViDGjF5yXipX0ydaVvgGsqZBTC1gBWzFoi9Kl6
k6v/cB+ElnCCYCWlTluRTbTQddti5RRSLhDUXOKmLfiSwOlinLoBGhxMEyxxM0J9foaaZFh5Cj6Y
YjLktBotoPdGGXEWIKv0ZUWdLkOIC5uEBPHguusDoGUDGLDFLA8MZLVTiplhZExmtBWVQvXBtxKX
QiA4wQoxPnuc0LxH+L0THLYqmm0L5f6oCpJhhzmjRjtW8SjOX+pmYwwiJrh9aSICTW4bYly7OPjz
mFjSw2dIMS4/UACFAn2lD1u0iGysLtAxkZBsq4ajcmVQJLCxGiz9CfjdXLMJx2e7inl272GuSusR
AS5C8IZ2n/oMThHza7znuNLunh9raxZ6LpHMLqAC6Yg70ogva9I5lJUIdyzlDPKu34ddFWd4ifoB
VHI3pv5/FGVxNT+zMUmjtRtYt5vOk8O6A/w4jaYJR3Au6nIiLHCFPbez72Wx3jlD3Y703K3bcyso
MHaG0RUZs1o2phe7/UqUJu2jJB4R7QdM9ovHLJ3MAtA+jJGMZ/mTwAF1buZW4i41RA3T1HwBr17G
zvb5KoB1vttMbKd/p2U1iAVH/Eeo2yHjSozdjmlyuAyzb1Im20EYOZGwG9tHR9uKI7Y9wyISBTq3
XCuMuLPwyTNBUuYBgRzQh+zd2Mj+UADFaH+8sOv/5ZpOvaaop/GoLdwiexsji2fBV3dQiDeJcatZ
etXtLAhDheOrrw3zaD1LWleah5p+1elWrBxPWSkE6BYpGpYklzIdE/Axd3Ro4SjBbKYSxpyBe8Tg
1w82ATEk1A6QZvgWae9XLezwPMDqsJy4Qj9vcVuvkpSxAJaahc+ESjYSzj6IoC00C0QQiivNJecm
6NjLq8QKVUMXVAIVcoaqI8/SjPDqArl0D/Ne8OjINC64lgk23ykZ4hVa2TdzkBBmP5ym/Q/dTD4A
2S2HDu/pYxK1BPtaDBhi8GsLA0LMG1TaAtfin+c1zEhaSDi8YzUWDsQrvkNau1gVhASwHn/YEwzg
eOPi+LOsSdYjkVIQObghPKE9cie7f+YeXON/lHhRQdyu2HGt/q0VVE5ME/WDG0vhSIwkMdkAoqhe
+3+eW8bEhTt9AhHfsz9e+1ueoABMi5bQyYDkOh3x4FKX9Fd1M1KEMqSUl8Cm9Jt7HDm2cJcCIFUR
RSCQRjKRGkCuCoho0CA24SQBOe4R8ucb1M4rKy+T458i1P83fnP2v+xKvSEd8/gjLmID14lfoVt9
EdwIEGu679I1EhVl+wikfs16PIU4ql4xq/RGXmgzRM8CYgHLLs4UaYmPOn1cn7GPw8M0AI3b4AhW
GYhlQSiuo+HjnImjRYRGyV7R1PkGmn1XsoAuCc0yG8dFwys6alNmGkp5S+Ea9UQcbrR2fXBxZuAa
11yEj/ziWGrzWLs7ambhBV2dx0Hhzg197nAtMTDvu/3jWJBYM0LhhpqCDR3anQ0Q5WwKLO/w10Nu
uHldllr02ljBJEH6eNwmzBCSc+8iON1KjnYONj9rgZ5RI13j1+xpMgjxP8GnratQfPz9HwQF/sDV
c7amYthc/L9jst0U5l7vyeFdTJ9iPtywqZxk2eVm7DTCJH44wLPUnIImU5N9rKfmZgTdiN9bbTBl
j+eBBp0rG04YDek4FcTvZffNibbdx8Ea+5M06AX3sKsaeqe8IQCO4CFxWgxbGUllkgQu8/SoqkMK
mwvClPowlZiTMk0rGPDuREIRFVTATIZIxzvyQ12TcCUurd3NOATerMy7r/n/Yg9FudSvAetLODsF
ijt/pxmu9eLxJX9zmALNCnulnJ/hBLWPVFo4WyMwP8ybgHOFfTbo3fSOkl/3S/Am8XnOVLVejL8K
aShgp4HVw06YtYJOM5MMWX3BlLwGH4MolfV2jOvUFZ8L37hnYUYbUqy7ooYSiFxVmC3xiKI5m855
2hd3+xRaf8w7B/DXnNdfH7hEVhnkw+lweaCfwaLBxQ+7pdCveuu+E3FrHR28pdqpv95AGBVHtdIa
vWZyq0JJFWt58n4D++jEI/DbyMbdC7tntlv6d+dJ9T76d9JF5oTfveKOnjwVzZl7IDsJYjhH3v9Q
Sad6T7Z0ho6O96eli3IHoUAjoDqJ+1WiNVjexSYbjLSXwSWyUqpZkbhmzypdcFf3bvaDbVq1M9Zo
VdnTCX3z0lOgUSTL/WqlL0GOVj9ZhtWA1iJQ7iXCmIccboDB3gGQmljLObxvlpAnqLilbb+kLzNR
e2ovioMiGoG2N1/EB0z62/MZdr3RjhCPOCLUkKTvMd7A2khjus9czKNGype2TZ5f3lsrh9T/9rbi
Hz9QYYf3N/b3PsN7cByxM4U80M2efBP0j1kIlq4QOLXiadLEvZ1Z0uU/4pcKH8lBF9PAYwvM43Tn
/x+ZqHUBBDGm7LwUY7ZGLcCphevnNANB/lBbq0NveUyb8FtU+bFO5epgGM4lS1T+D/2smlmmUNAv
E5iOw3zJuSIU5WKZOpeXWXBSza7WTdg81c7gxK7Ivbt5lVClU174brUZRZDoE4vDeEV7dwuqqZNp
OiRWQaglzJoN7w2ryNOp2iKRhYkMxwHptmsgCLZckgAkS0OkBGpj58R4vKQSEWnADagH4ggPlXvl
roQV8ztTYa+ZQohgYOOBLwBtjhHEQtXM+ytZbWUc9pZ8aY5mr2aotIj8uTq13EyH3paAcsICXE+w
Nf2X7hTpboyhb57rZnWJsORmoEbrDyBDj7bXi7FLYzWM+v2qNGX2aL29/5dzjsFiEpbIiey5LHav
cWzWBjjnz953YwZvRx77j/yTjs1pQqhi62Mt1vLbQtDCeYdl2BGTQtXBNJxSKhaIbzlZ72Kvr5Br
WN6kusPIxB3/rfCxR9BMDebwItJMzJ5/q33pX+iFSKwmJ+0FSnlGZcGzmw+Rx+IJTFxoMIgmoebe
p7I9HyYzOeeZCZotCNTP1IT1YjSWLdPxyH4xMOYrWPk8rVnU1ovkjLUqb7o4wwPcoQ2NBhPUISz/
QqBbl8qqAdS9xV3Yeu9g4v7g1+Bg1rkaessxLuPYGiYW4wSJMHKLDvtd7QPrsbE45Id9/pNEshx6
+zLxW/HXhNtt8980Z5tbaqZIw40GP+jbzXjqQGaJ0WSJVRa4SKjHG6Ctl4TFDhYv07uziTOjbQnU
8OSkXvD+rrka1dt9qgwKvJC3j7KS0yAuE/7c21VEkErlIo8VpZogVJNriM2Ot3C1c+x+IRbzQi2N
9G03LNwCbrKFVTu6ACFNOvp5y4dGMIvnJ5kGA/tJgeEZOGFxX38QoIMY6bnOFQeYenoiZLiY8hhs
SBjQ8ddmvRvyG3J51EWm35xjPbY7DuPQCptw5eBbEOlU3JS/KHGbxgb/sdxI41vCLhuAp9n7Gfh3
HuwNG/M8Pt2KRz5+sZwC2YIw2fem2bbOEvH4RPxSAFHRB821G2XvwP49GFpmJkMwXt6biewSRUTY
KAld2MyHI4vP0lHoWhGUK3qoA+eUm2xLrPfMY/F2FJutk7OhxZKX6rVZxnUtGCkanzpLYCn6aoA1
Sj6WREVSABT9PRjOPBXmQ1El5P4oRZYtWPozf+baGP0pqwJDvsSJRF4vgvviLAOk/g4M7dmJRTbe
h4uKV3z9G4i77qkkjfblTTEzmeT/MjbgwhYZgm/oEJ4TKCHLX04IrsUZxe1dazhH4MzLcKd2Aiev
ZO+Azk0Xz0vzHiU4SaUsQiOHpa3OVaqq5pkZqOhmGLKR0lXiwn92c47fyxNza4PiYgy2eKz7Lgi6
+Ddg7knlfPk4tfo2qLCFtHJ6CS7hROrNs8uYIufMocy1HwfX63IFJw4imZN6P1bNHlFfq2+6kXqe
2iKdaaHH/IKYX3VJeYsGjj1Y4UbZFpHqm+t8oQQ5IscbQNwx7rIN3i8RCz5/nt/N0xvCy+970/P/
jJumzURyGve5vL05t6M5IQ8ZOwWD8+N1u9+DTbM5FsnL99RFb2sxWdmXVlA2MIo5ETgelmFP+Til
JpxfkG7m7BkcARdhkKLQicmzO4NdliKojEVjoryNIj1VEx2NtrGhFSKbN5KJxFEhGvCqxfA3dU+Z
z1y+2UgSYXeB5t5KdH40lm0ve0hoa/q4u12VS8EzQYsRHMsZ0J47ehYUCEFY/rINE/sbSZ3lJ7Uw
2moa9if3SZwD6Dl2humTudV0V5ObEub1Zy4I+jFzEuTKXYg63nstDmmbWV1pJfEvOy7vF5c8ZYiD
OcE00kvGIQfZXVqp6bx5sGCOUzmMRFJe9eNvu3UOnsVHAsOmvL8D0cRivjuFnIxu/7h/xqCluCRB
R/afgQt1zDNYLN8mNhIp+wJTz3i2Qg3u80Hmae/dyJV4cShEpRAmrP1cDJBUAMamZq2vka41UJ19
Fvfl9zb9Zfa6is5weVs9DahINWoP2lkeNGD/hc6gysO6SfjbjaFVqJmi62IrxRj15hp5ZZzhxtCt
7oS+LJ9GAvfVLSn0kDSSe99gsIH9ir9jS9L+niVGWRExJu/2Qb/Xf0otHUa7IQSGL5jD/kX4zg+Q
Rp8uTvB8qvVtBG+nqqA9sSCngEwauyMuvKN7zo4obiC7gaM4II4bzPFqevZulpw4hRkYlxvpdI3W
0CB/Ncjh9CyQVqwn0FfFgEvzKVCLYMm6K0sV/oJjC4vwWDMycUL5yzOAesk8UY/JUtW4icgIjosW
wo6X4qP967W5AzTVV880JAQP55wIl1A2X5G90ZNqawMuZdwK7ZdvdvDpKIi49EEutqB7Eo7u0ucK
tboFzYdPjAgMx7qWmfZCrmh5gN0SdqndhGqdWjUuFFuCKUxUMWD5/FRblG2munZwa1QOhEBu5/OM
LbMNvwypqX++iSUaO1KCUpsfTBPZvIl40q91WpU4irQMut3v5+DZFy+TdFlD2w5hCA+4ch4sACnA
HAqZhZ8bPb+1NRTXJurisy9fkpSr+/ku1d5IVF/cWEz1FSHLB+l/evgfqUgEFOg5Jd2urPOHL8UV
S0glB/8JF1Bqiadc+zOXGn+ct5mbNKhhm9CGiosREWyPvtW/fToaP2l1NWyh5qO9Lagdr81A5juv
+qi5/vTwPYRJUJbRYhm1jxAOrIinmZMMq/rvlAUkoaGxb3It4Th3wCy8zh98C+pCIgU7KPRwI1fJ
g5hod5c8nLLthVNfeiT0Hhi46bMUBui5nZl8kdRP4Sio58h4Xb4lBDp++fXV/clW0SD6nvrbzO0+
XRnvODuQV7crH9wviQwRoPnqPRXGUo6BpROhEhHpuJYiZXeZCNyvigJ++weL5UkJdRnr2CmARQFy
HhDhTEwk+G1XCg4GChKalruQ7ujmWWi4179wLMA8MP8KZcJ7u05XEvxTOAULEYqt/z+nD/KXH6qp
vqUUGrOBM2oE4cjoshInrvJQALXgayGYDkRcS0Fhe3oL/uD+oHW/QqAwaBys82EixpMLaFiK+XIQ
7SWn64iyCd+Q+6OeSaMHqTHiX7xGvQkWHzL6a+7SkbU0+AIWhzP+9MzYvpjVU2CQ18xj8vpdXDnJ
1Q6p/pZIxZJN0wdSTEMU6D5xqqDvpNAz/eytdkjQoab7f+dYYWm4PVgiVD93YbPj3sjW7k9lwLVs
wlNi6u6nTvx8fFxE+fu74uN7NtRES3traxAx2Q81ywXxfmY6TgZDpfjACZvUdM7V9yp3vtpKb+Nm
8xn+RDQg+SwugDOJruMq83y5G8diAVxYkdl3zmXmqfhWzl+T39DP/72+sLvGDnab7iyIvOLpBdN0
8CGFyxEqDCBYIt8gxxNvlGzChcEkHauWvHyxkSfWVHEfrNxDoCuoPWH61sysyN4ODOf73deET4c9
8HwrDDJL7VrpK8vWFXx6P5Gn8thku7Ch3qKDelnugH4hdaJPJsnq0GFar8dR+BkEKHd4X1wM4JIx
9tp/IGpNr9nJMPkFA52/rBenG5vi9GRiPrGZID2nLCnNbqFdYUARoMaFbim2fX6PQz4SkOmB4+Jv
xTMaETl17oLTpDKhk/S+qt/TFgTBiafrjxJ+nd6R5cL7Y46/ngpIGInGDfddhZMK3iP+j/SlJGb4
3traXwKuVOxgjZimB9Ss5qe9/lHpi50C/jwd4QagxXsT6WeiusipA91RUhws2pqGD4VsChd0Fkz1
MmnnJ4VKK3h0GXL4iZoWVQCE2ayvmF7VswPhSh03xd8fBFZ0A66r+CdJ7S9b5CNF+3V7FG0uYbeT
siX0/CHwJd6GYh4rZKqYTEXk6m/3IZoRJyAI+9yZF2yZucMHKu2IzMyLMIy+ds9nABf3EqR+8hpx
TqirbpXHI3DcsW3V/C0obQ0sVqx46cBMB3fq6W5p5rGK3zz2fgRXFphgsPCY2+yjZEzYTieARW/a
pTdCECjSpXku96BJxwLGntos5oW7WoBCM/0aLYzccYI4LAsqG4PNm+TcaOlHybkRg8Ucd9No+NgW
SqPv6lk1jpt6v+5KNEPr49iMfBmUj2OSD3E4rSUVu94IRMHnla9HHBndIHKhuoKRlONxP4Yepajj
0chWJ8Mu2IJow8dC181NtUi/kFlbay6VukS9xrtQmkNtICE02RHvx8j+PLdIm56hVBd3BiqqtuMh
ELg5cC7ApKaEzMeyX8J5cPZ7f4XLmYIaqd2L0QZp1ZSdWKggcgMcYpnggdINEKWuqnncTLKj+65j
nCUywYj6lKFGvzP+1PAb2LmuR8H1f4G+AWbH6tVvVf7byo0j/UTSsfdlBm7knvzIkSjJ30hp7N9c
840Ruxow38zIj8uAFmxebwfz6vkB4D85rnivsJweM+Cg0T1zqw8m/lLAZUs6xm3dGu5TSFHt8iIX
3UMjev/kApj0Qi7zaj1+KX4t16itwpVaylnp7nYHz5VmUFEhTsYWAQGI22hiLwRcgXrfaKiC0fpB
YQG9bK3pYIzVi3nuzo/IJxKN117kpX6WAFGotvZQ8r+SbUR0TTxIR5BTpEWtdTLxtJncPimK3yaY
SM94QF7xv5lUXMR+x19kXuejh8pIfdC3kTPk/bukfuUZUvwwgMaib0yZ85qN8pHZ2qEY3YN1gKpd
sGs7CpXk2io7Ay3z7TVvdwStfdivVHpJCrcrwEeTqEA397kBz/aqF+1DHOf+DPCkSo/9bIl74gbL
6oJcPaiNRvMAUBHgWUbo8hk7NY7vG05DFoAfufhZY1TYO682VH07+wWETwtl/kqN4mvpFUv9xA+3
FoGRJOzL0i8Op/p2epRR8zBAfEWZOP0DBJ8SaAjvs5df4I3jhKU+5aRMjoRbdURBT6clmKMlaxFW
QeWUVaZoLV5RZ7IYvp+0tbZexorTqOKEzS3158l4aqR9uJvN9V00+XROtu+OlnHtUOUmKO0rs9U6
BlJvniatMfsHT/WzAIkGUsxd3CPTYGt+SdcRZen0cep+ibl6BQatAoax6FByWKx+QMjHIEp+77ja
2eXSh2YFl8rS3LN5KnLJXI3GTcsAi5NYCCI4rd7N6uOZ2D1SRS0InSN++0RSzHTfFBBWRukp4eTw
u11Tttr+ZHnzbWV604Zff4Gf1k7tiuUFgkGgj+TRX/lPN5qk10tIbfP3poBIl8L8nHSK6hpPPUcR
ejeIYP18ZlhzPSx8gLihfgz2PW5pBnvw7AgUceRw7wC3iG9hst2Hod7dEwsQtT1u2a17+E0JimBO
wo/BdvtpFigLYy29VLFpqFUuKBAFDIMLJDwt1+So4jMK5D/8SQjcB2QeEWnrWPLz+b4MsE+uRqsJ
ZEQzR/CMd1BLoYKSnXkIIQAxsm3b6und4cTewlLfyUQH0XZ3K6BMMohw7aUfb/Jz3sJhZPNfaVMX
Dfsg2eFq02ifhEepxc0mU0uL7rM4PYP4jrtGayZkNYS+sD+Yrd1oQtAqHH0RJMU1oH1bc7wyQ5v6
ML38i9po4Y5N2BPgsDw8atPRxE61YqVa81ZlukqRb+vgPsguD0As2QSD5yXv1Xh7HFs5vlpktNKq
SOzz/dNvaFBs5bVIMFaMdaNoq/LXBmQ7woeIHnmfT/I+BBrwaGMSLiIE8ipFTi39dcn3wWyUFC+q
BH9E1ErsDLfkS3da6jmMto5Iav4vL6Uk5Bvm9KzjHSEjK8vEns5NqXIVuIctV3wz4ZS0/sABKhPL
vU2qJCVoDBGMbYf1iZleh+k5E5uvM0kwGm3pCfsYOWJp2DNoqOi83o+5lBBu/mVh/F0b9sFyjR9K
DWywthnjpTun+UGtMc2FMx4H/xriGwMAxw6M017gLUTG14i4L/3Yf5mLLq+leF3CPBGqhrOujKLl
eh/a9sISypGJ5fQShJnHoFQzq+LTUhNoA36078LVSKMyjxsudl6yNW7JgOm7a92R2cqAHSbWLCn2
pJKZ/NVutgNZg1Lq2MQquAUv7v9DKwa/6scUeknOUgKJpjSRVOd7TYt6CchDj7zegQN9z2qcYBfe
Uj1LnibW2Pd80tNRVpIxWU//G99ex8RTn5D5P9uMfK2XqTJUpPuifVNdbxLfy9ts5XEpqxnauVs7
ZT44NHwFhF50Y71UWIO5dswXidAXRjnDfAUwgCSnPkXxcGwDFjGefbWEGfpy122mUhQVQ5bkWQoR
ugng2i77PMlJSkjnmNJ7TJRt3PIF2v25UC0Do3zc5kopflLMu6JK+Nn/imgQfhmjWI07HZa+yN/p
EnEkGYqxd+FbMcXQzEokY32ASeUATBDOo0BQhGtrN1UIBPv4o36yPzW5azgdDpjq9DfCKxP0k0q9
MvtJUG3QOyUHKkESDfoY3AfyVUH6SXr6+XD6teCGJfbSSs0sJPP0waZ5eSxzSI50yK/mI4IkUC/p
oBOUnfttrqv0r+vj4OkAjmbF+utKjUqOUqYvN0YVpk3vcwq3EUpMmfpRm3hz+UkqwpWgO22CG6xR
mAmbA/WmmiR8+Hc+J7Bz5oiVENYa+spgMKJT+3MIF2wBs9VKUroxf7nTn8g5762dcdyL5gUwFdjg
/H2sK8aUL6LcDCDJuSqku2c7E5CJTGoCtZISaIBNxIokJk6HRFdbLDVUzA6Z44MOd6HqmLTQv4xf
9UqHLM2uzmUkKFmB2y70qlr82v4PMLsKaDxWM9AfqX3EOQuqFxOc8l07tZYPEuM2sqfP9o2fNlOC
OpHgmdbePVvy8djhCq0pCXfwBi2JQA99oqnjS7KJZKhCqMGbM+BgxaJTSMetpoJMdLuzPl7iTMCa
8CtBSUtw82OER2CFarCfYElv6NMM9xPICUlf5+J7A60q4by+UYV+TpETpQH04SfFGGfbSP8hBf9a
svfqcz2NB25/19TMKhctw+kmQfoZHgPiRQ89I8mp2lJ6DfcqFaCM1I4sLCUqNxLsHaasudT6Dqt2
iOozF9jTBSbvjEDOXmwnQXd3OpOR/jyWLDXvUufEBD2rmeXQ/FIhAkFUnDr3QsKwvgG9BEHarHOR
MzBimksdDAjKfh8Mv7/j82Ppz4iibK1KezsHG3RtB38kcQU2SS9CSDOzvT98HjMlqoFEqY9NjMQX
vOA8vc5fb05OqqFSTTOITnid8n+HX/CnIw86pE+GJjqqPpIBH3pd0POPeo6lVXWabURVAbrjHXmc
Tf/3Lg17AXaDCb+GZwkNUMJpk1jp/iYKROLyV+wEP72YArIa9byPmkDiSivhoUD5ggZYHQM7IuJJ
KflKq22GmOyQMgNdQuZPddyDxwYw3MPo2JysurIQWBR2UptpMaHUtapAtiQ8V+DXJGUZP7aSjwPM
Y7KvODQa2t8Q7hLDTVXaLNIX49vORJQxe7CsZlkrYtn+kNS/MWX65iL7f8nAGCf97ZYi+NeWPvT9
BVh33rSOytS/0H4zDJyVGSZlaTgwGucAftW0cPLjCaA843IVu5ifla+Ijs/6uNzBmkjtcQyFKq1T
Cm6BA5/nrGwvmgGuEaTlhy2aX73SoVCKS0eL69egA/9ymtc++gFStLWS2tjyYnLtTKNQZFJoA8Vx
d6uj2QJEzc3Hm9Ab5oDWfHryBLp+jwjUPcSQRz1Uu8aiAXhKeFLnZEWznL4LG/rbJA4EWxCn54qB
mZov6vgCAZ9db3OTR++/7bRzF+U+Uhh/TGbuxSw1K18x7EyT80flicffVw8S8deICw0m38OoiW6l
GxvrUjhHH39W/2IiEQNpZZq5jRbwvldUdImoXPlGX3m8E0m+haKES3OfaCTQB4btdUB06oIg34+j
hGIaYcWNiD7yah1klqtorsMDoT9uVEn8GTk6jo1kupceb7QZP6SL7dXyWxUT6lM35EEzFJ1Xtw4G
3rAGfCAN4Bkad9yl7s2xpqUv390JPXEngM+DCZrzN9QC5rRA6f9aWigYrJK5S8G4qwJSE8s98zSI
K3GimFyaepePTJuMaVGGb2350viKmWIDdalvJ8Hb6WuV4Lm/9Elb1Z5OrSvCg7GR1VhLlPlWnx2D
1Zc+ikF88FqhNEBLI/lVtfME5Kf1jNkIeesv9I0PGlxOf4FzCg2ZuU9x2uURJ+638WR4Yr17XTp3
TBeGy5MKsTUaur7+fZ+ZRTXoGwbKUrOk7Z1PFZoFSQiB3qwmKehf7KB/HSeFHo97vm6rEgcZCdmN
4yGhxINtY134TSfoOILx5nmp5W3+I64Z12iDdAUF3RfmwyV+JRhKF0Ttn+dIMt9zwoRaB9qbWAG1
sI1UbszKnLNYkcAptXy7KrX0IE9W2HG+N4BAvUmcrQTtU8ahmUkxXRmS96CALNoIRtuchrMZiVn8
KxNYD9T/hKSNkAxaXjfqfQoygrvdSnfhzYjkGjU5FbUPkv5SqmhvwxHXzFF9kyetyAjyLmtAPof6
0XS2zpNOpcDEihulwcrm1zHHX0c/TyvKWOgI/Td6k57Y9nmBbjH49sVf4JiJWoKqhWiOod7n8Ypg
ugnJI8kKZRl6oRMpChGxNYiIeZUvb8zG0QYnBNqhDSoHTJ2rF5xhRbExEG6fDPqijdxVFizcKWsN
+v0FHMW2tDOIPqYAdoGyRn+YPfBCtZ3fcci4KKK8Dyzz2SgYrc0zv1CXgk0XGowqnLiuXt0UHHAt
LRkQVPbxNKbgQ4xN0lokkA99utG/OYA+oG6tCEk+pYAh5BkVDpoTmCrMtd9jvXI0dMhKJYmAlUiy
FP/4UVhDdVV/h8wqviycjzyFCWxqQPE+Yd9seUPXSbPQzg/zur2epsHPDG6A78zeqw7M+L8LSSyX
ajKz4Td3Ip1rsblty8Leqz4TpRamnLkK6+OOc0wfOAFt6laZ6n+JyMQ22LfQcyidgK+8KKDGWD5t
yLlubfk6qnQoqyDvNHMggMgY/tPGc46lN4S4C0Rf/xg/NU9ila20eZIGlfFaSt8XP1M19bF1Nffq
SyzVO73RYEG97ZBo9djDx4gYIzY4p0SlqvmGXv+KR7VLMYcfzK1/8DKeUp70NftLmqHPkNGuzWQq
BD99qMEwxZgbED6eaMZ4vOujT86/Jyw+vFNCwkUawKr93LtzYcJP8dSBXoD/JvZxK+4n3uRHML+0
kCBJwVT5ZZcWbaGKlqoOtwKalTLGyclOevv0n02U5N3muqWfIrLCnwexTrtdxcAIft0m3ehx+pUo
QTvJjnc+sEhCjO5+lEF0zl6mFUg46koaP6ES9v2U2q+KuqkcZNrRXIQOkZ35gvw5p/SeGFdvyNff
vtwYU6KYb3rRfI9K9QZl7lDXc3wyLGoEeB+ECoThcHUBj08rNfSu1ZGVrs+kXbipjQnUsP2/8SM3
ixuAt0ko27WrhG7BwSRWTdRYRdURmj0IluMkt90Yr4gs98EcqPo3iUZetnHmrkkY8FcxviSR3Dhr
wKdkvyYkn//sZc2P1F0rbSQLyNUqdh2JWtQRr8/bN3C5epN38jb7xfyo6VD+c/z22RNJhUQY18pW
on8J2QMhlT5AOmX+8uXfxqRNjqcyP/046bVLwvn2DkqT+sNM0iDaoqZwb0n2K9NLYOQvQ7Wvr6Ur
7YH7J9aMTUR1o1mh5HzQ9tw3icHx/T86ULd263DsuCrbPNSGpvzrHcmFVkJbP9UrDugkHwUWr61/
nMNAp76DsXqtXWLrkBnot6iGTHDvtaxkDYfVaFuHqG3R1HqabpvGyFtWr9KghvJQcW8Pl/xzhigV
MHV2vQ5ccFpcaporJ5DK220DXZNrDi4I5owzDVOXFW0blrMgSqjQH/GbhwownYbwtYgkOibOu/vM
QDIn2TWGlB0Oa97/jVEFWz9/zwlo4LAZTy+UeAikO2m2OiGB+7QafKPvQniwk6rWzyMBjpnJ4Wxj
HXgXZ/hXx5xh01CxZpnmN5bh+Kf2pfEh7Bq4yxl5/R516b4LG5/EsBVZt9t29ayBuVistNIGCfYd
NSXToYjlVMh1cRxgqcl+4Q6Zm8dYUwqDuYn0fy/frCZ7IYlsEBmisdXB5yHeDxbc/yuFHsYXHirO
L9/Fijp6IvQQh7qdpX7WZ+evIisaCqhYq8wGOoTGwsDikCS5BOyKyjtjDwy3iu6aBMTW6Z/s8/Gk
UoS9f9xsf/YpEYL3Xlg2UV4ezTP36N694JgE+dbHgpoGhTFVwldL51di46yne/pCXW9SVMUcYF0e
Ueb9/0niYJvjdHvmAP+CIW/RnCZMbWrHxmLZ906rCjDRS9vP1NJRGJzZvzXhO7apxsFUYLI8GcZm
L24TjGewQQQJvfwLv3EMjwKXpQose1DQLBtFz5MI09ssqezvkkJ8kueoWM8TWqABcC3JkwBUTm1E
I3tcOjKu5h3o5NN0E2QiGxztlYDb52OKicZqP8HmsM1xdZhqGDGSq7a8P4bUEJ5nrjRp9rLhx3fl
Id8ya4pS4avqMWOuTniP3EBHRSKNB3XwUPLt/hVKiKhVEtnrQFhRcuvHn3V2nf+KuYDT1fkBElgA
If/z8n4E4z8Wc3BHN/bXnXBkYGoGI18m8ljlIZ+HeBLs8ad4v/bzlC9qTGwkB1RINcNNC1qs5BKL
/PS88N/g+IZUf3+uyFpTr+KzhziW1+QGmPfAYK5052IidqHVrN02zH3Rz+SQdPzxpYKQ1g3PCyJ+
ocmAwmaOfadknvjOOy/e3Bm5HGtAN+/0IJfmpzTtfCoVXgTWUfinxeZhQ9cGuoh1zN/6K9b/A6jK
h1CB4H3WemHCjxxSOe0GGhAbGPI9AOQCv+odAGCH91ZqsnJ6ebEY+jmMavXtjxPALO2kLM3ynUy/
ZntrHp0JiEcunzc+XLdoaOWUZIAyplpKyv2YRqfgs8rKq36YOIHn8OVJB6tE2C+Zf3xUD9Fri+Nm
MbR8ejGJ4jATr4igd7eO9HzwbKTc/mgIH+3iwU4ttzmnAMR4NcF4PfbH9Prz05pA4gso/9NCQHGv
QzKTXzlmL6LkDlE1bK/HgQmEDX127mTMkVVixDIYoAXiRlI5mto+SgEg9BPjTp456PvpB6ub1xAU
dbFqfgFWG0NNZbIxAsX9BhUI3ZwfvCxj6utXmj//fJ+0MaC7BLwYpZQbAsysA1+SQev4zglWzBCh
j/cKT0h1kNvajcxal1grwE+kHaxGfTxOidSxgpI8bdQGhGJbsMKYmVyk7gjWIPHalIUOL8H1Uf3W
DKtJYwcGA/xdT7G1Cf2AlA79B2CmIYW5rfsKPZ7ebj/9w6eAix5xfRTwzrcZAn7iB9k7zsw+7Qsg
D7uPYTNSMQe8VdudwlfkfnApbDXJHMhrDBzRN7491a7IkWZxr/ELMYetaFmyPcKNTqHVWJVivvV4
kPlIYsDBHWAF7WR5S9DDifIHnPgsjDySvYPN0TenoCYbodnNUwYjowP/28Ae4KRLlEwyroVpov/3
5XrlWUYm36F4zNEAh5LI78kVuhC65YP/WaWoX0qSUGvlDJXmgXqJWCcU+1+DDUlvd9LNw78Gwb7n
NwtshHSTUWT+qaFxKQKObcN+ybRPwMgl365nqHurzNcjmpQYsg/VM5Ztq3i9sHxxKkGWiQNdf91Q
mTjSehGct/ay9w6VZ2dBItXjMhMIWDptgscaPalaXQ1jL4V2F7u2Y/OHDmfVLMZWgXnfjvMssQZu
aflkaUOVrInA7LbYyT/2bcrH+wljmVD6tE4n6zu1voJvNhNgdeEPwetr7e5ke1mMSdD7hWA9LKnk
T/LXNjaLiirEiM5DfyglKClVVadl+maXu5qWVK2V976Z5sCzWLHM2OX675Jbs8k5LovwKW05QjgJ
1bRBNFvNLsqUegG32EnZ6fJB1yWzYy/+ZZlMQTpROeMMPDKpTlyoPMp8oRCffUh4iC9eELjzXKvs
hDXpKWCy/iB9uXspI1AJvXVmxdaZ/ekkm3KxiLQ7gXdBYiFy9hX4a8NQmTiCzop80TBPl2yj+6/F
XImNSSYuM33ciP1RuaXYEplmFZhkJBedKABBGEPsbWLfQnC8JIijQQlZyAJGvhiVztQDNQdKtXWK
sokAFc1dGDDp0HygstOIljfpVWKrRSmais0MxUwUt6DjHNA5Cwrz4IXXw2vaEOtysSF6IPg5rFMI
0lfkiP7Cf8UAgKzRccZ8YYYdDNi0QH0RfdayuX4GEgEtb4gwGpIykCO0nJJIAVkOVYNOogkV2PfY
4CAC0u/YdGd2R2+O7c4Nro5x6/MVRvjAExYtCkTsSF+8feVwrmskA2PoX1fV96gTDeJrIAr8JRLt
pahDiLA0Q+SIMQwPtdum4KjoFZMPxNO+Er6xjiOTGLKuN8vsEcxQKSmLJXH6NCbpeg3o1bvX/xU0
VhrjqLV/MN2MO/EiMY+ZcA2S/s1neRA0KF1bwYrXrXDnW04DbIhKER5jimE7k/ZYTYi0pVy+l5NY
OEIPppROQFCiMDvhb4HhFSOlBoTGG+RpOzY+ucwH2j44VyxygW77AMH7ehTWb/7vgr11R5bxyXKY
2Eco8NCB7tjgWedw4Ro56XuSRwTP+q8WpuPTHVvmB2sRo2G9nHav33jOUrmH+gHkh0YdtsJiZXbc
FSY/yp5dR8KNs4rJwLhXF1WxjtmTvrEndr8SVu1ZJjlAmtYjRTjtFJxPgD7YxRTquIbZ6Fa5do4L
ezkWi9uWCkvd3mZ5JsG2QkHwudDL4Cj9l+6jG/7QuQcmgoE5c7MdZ6VSxjLxQwPixpzkRb6OmqTc
fTNV2OuzZemVn4dbV0l+u9G3Ek1xfNK+xPhIYw4ih3022BmOwhW1thvGiSHfdCbyKVz9hibg2hiI
iCLH6ktmpDEIjywAxYf9Y1KY+ojG8jKKHwMDv7iCfC+ek2AlRvX1IfOFBjIR/GT3uRnLZ31Aelhe
GzuZRIOHZymXvrKkDNb2YhvAllQR1uibwJ2dl+YBYrBvkgLiVuyUlC3aH1yEb5MhctwvFrpPWknK
KQHI1Rgn7rW1+iodFWPajQcFihxHu8kmp91hUwZhvuEgkHSJ/fDie7RJnl7QFkAnIQ05cdxZ/yT/
6+68fY5mMgHlEw2GlMp3THThepIVQSBOZtILlZnBVeidb3NlbWJd4JC3/e0h4Hxz26D2JLSqiuGb
2Hd/C8fyiwP9WL5oYO95owlPFuT9oYj84/cJwhSEHeDs5PT3uAFaL4VAkexI/7shy3e7Hiptsdmr
OxqwYlMPhR5uXiYAWNGGBSk9QCzxwXZE2Ka9b4j86gaJhNWSdgNDXdcCjaUd/8xvgtswp1Qut05z
LtzfXcyimskd43/PyN1cYhK/gzAetoiZYIkMvwkgCcGB2Um4BhF5HrZE6p2kbAdyog/+pgFWvCWN
Fpcm6UM/T2I4Y/1FV+eInnhc9TRjaZI6TpAAR8HL8A8CEdxyYrys6SK5BI5+NYtsu5LhNL+fmNHX
Jpm3bPh140KWuU+RUs+f6SzbHKlc/U4onjAv5hXbt5+oOtIb3S9MfBJGVpntgNUF6EZUQKbxtuG4
6NOJTe0cRm3OOtMemUSWrZlVASIgy1Ct5cdXAE0FYxvcVF+UkUFmZZwsVzJgv57fkUmRWHnZ7OFQ
sKtBiK4+mBgZxT1uGj+xZ4mJcFduS/BoYf3G0pp4M5p4Nb0Z88Vb8ia6RgLDUyTDL3rsoLIfTiiA
uP5lRz45bv7U5NNRLwfF6NmNigCnKy6aPgwlprf+ji77XpA0fUZpAlWOgylPE8hCfsNZa3oin81W
0699A4dxs9vUfQdr7NVSlgZNyGIdLaOfAHr1vrGfHAErytUU2FDpTd5XR9DR5vkVweslh+4NJeCf
vBs3ePxsSQyU987MKlxxtkTdc/h/Nt3K38VH6NLziwUQ8VS8Lb2nyz5bkIAABlcSP8LkLuxHOJXA
7m0Och9eBbzZdtUEVx+vo7sYyAG07zVwdNcdAuxWFvyu4N0vZprIiPICL4huXh2QK9Cw4qSp0tLL
zIuaoDp+PSak1aTbnfTH5dXZgDMn/P9aLLWXUP0CX/LIbvut1KQwa5gzKe3Jwn0Hm2FgAlw++dEM
J7U6K67JXMnsXRkvoKnr2jUOZyemW2xB8WKjqeJzvfYpyrjPcMlgRGLtRLlYmNNWda7eFey6w6u7
AiI2WxYhLDYTBJAq2mO+i4RjSwGB/6tLBWa5BxX+8xrdS1P7EtrcCCYqrrnWJbH7hQojLze7kwEe
AdplB/nOheFr3DkJmPrnDWOYZWM8xqtJY5UBn9YKO2vmeE7sofRQKaiwNRmTZTm6gyWh1fS2H/IR
wtVZDjbzmKzwJebWJP/pyiLca03d+VCUIABASPf0V/EbvYytDfCw+5DcGVi8kuAj40D7lDdtcJgW
hrtmFOtwALRxWzWhD0Z8mZW1W6JKw89PA4K5faed7+wuhJKHZ4o96ZyD5/PsXEz6fDfudDhuKptA
cqzGm9fquYJCPphBVk6C3zr8sO+s0+7jzlg4z+/UBRtF5MQJM0CEmBT1qSQ42dhLHOA/JLjmpWHR
J+bsZjM6gY06UGq5BiRStJ/7z4hvtnH9M+YowEm3VxqBmXLN6dxbayJz9Dj+npsxcio8rfSA48Vg
fNYUeCPO3yZ9YRhGHYRzifJlaygY/gskAfEtW+O8o3tf+cOOWWbZ0b3VOLfvoUm5mdj4AGhjtoco
vBL/6FacLy7KA/4tNLXfQFqbyUu40qE5gB+dKAPQd+UBBz4yj6ZImvKN/nVv4lE74bEo/bv/fsO5
1pCcn70KN7G0ZPctmxs+11hNhpllR+v19GEgTMFLG0ecWb/piV2Pf5C+4qfwvnld3A+VAPVoDG6l
h0BvFKhqisYSl4fEWuTbbYOMIV+Ya+Bco5PjK5yvK9pUz+taoFcjltlwSQt7RVkOXyzzj/tc07SF
dtRmGupTZSnCpeqfPipq00Oefkavz4H2uWcxcnwKvNGSuOyt6DgcqCyYYC0gzi3ucUqDO3Q1Rkm5
J111ctQi6pEggFBAMaZ+EzmSqa4Ed/S5KdKqV45nR6oXJxF2NlKIUs5YFCjDVb2uAc+15WtYHll1
w+HLmnjtLIEgUie5B9KnfgGkXSIWlWRhz2CWYyzRItdOXDdFTHiFa+MCFHyCTpqLmWRwmIJt2eGj
m3qLsaA3eUtxk1qKqU+eOXN7AFFJXWX53Agb+koA1X3ER/8k0fzcv854sw2dOPjNJqLx6wj/aaTw
/xaqm217Fvo/EMzJZ/NqrRd+L8nmDLtoNS/iheOnp0AUFHNQ0jeLC9MhImr9YVlgBLdJtgz/j7CD
2PI2rKIiKrW3qySNNgCK6YCRvmP8WOIgaRLhqnrZdoBXUtgGabrNpYbxkTjeuj2HQ0wWefc2X1Ty
Xpoh/HuUacDpvTNPS0cduukM935mnLDa5gyksOq+U9A66skHW5ZcEPNd9C8X9j7KFy5f1oTYuC74
73y4Euir0bXdinVWDMFXcVnjSiPYX1GlUdQtqab2TKkPirf6kUhps9btujOYoT4Z+mCrLu3UbD/w
e/rliDEd8ZxtVi3f0XelNbzZgBGHS7Us+1ymZqUUuvIkN+7tZO0lCSkCJY3WeF18w121u7AJ42Pn
QiVt0oKL0SrqQ6P3SFExpGtSirhjPZRCvWLeJ1WLaxlyHxmgaTrtxnZDU9lrSGK7WnIiXo8UyyyB
yD1iCOBDbDKZIyEazkifE9Qzxqh/WFo1TOvm/Kg+2O0xc4A9W18xwSiDEgUHYH1ImufnHqrGu6Of
Nv/6d7Z1tn46aV7m6k3gpWbcWFJjcJbmqervXyc9acJESe558FCWBhQ+k7eoDwRPXg4s2qIK4IMy
DBzEjOPpuqDlmdpxRaZ99HdPj8jqJ2QvYP/wEVglzfrK+kiRJJJGCgKACj8WnH8zz5egeIf3oS44
+BbB63ES70PrWYBbGsxpBwdaEp/ORrhzm+38hSCH+yOPtmp9TLyd1AA7ovtoh8MUP5YRuoNqFrgK
weZwHdnjRGbGauLTQ7YhhR0s4OuZxuijMlWcanSNMi+Ro2Cmadweo5kGOtGgMaYyH3z95kzLpx6L
n0Ap12PRyB8qWDRkbWuQK6lbhVFuCewseqce4mXOwZprv9xq6g0UAeShBfpXEcrLExruKfvdtmx8
NdOvtlUlNZjqwmYaiBSZZT1NwjMy3MQYl65UkyAbsT/ytrm9hYf5D6xh+6st3vgNaY624tP9nC9Q
fKEGCMnksf7TOblWm14BbkRWr9QhF3zPfogM0hVj3AZzinWWrK0jhKoUN9OyigxtCjZ/kRxdh0Nn
i4hnDDhGTB1aftWAiNPa35fQUyCnqZSW8U8F8PQluovA66DbSb2gilTVFdVYzyf8qCW10Q5bpR5i
qrJFO3k+MzazWo5uTzcMC9MuQEheR1DYjgEoWkba0bl7uMkxdWpxtZsmR40fdvWpPvJH1zyMHCYN
ifSuIVnGY9DeIZINWjRlmdiF4xqMJI2PVD4rQHDaG5XSHCxr8h94T+g/RPFOxrpxuzWZRwmDXW5J
+mgllG3wIUhwUtwUknRQyb9PVqxaD5NoxeuRZrlbRTZMmqaKT5QsVISUMW4NK0ADGe3801VzNk6O
Hee4JaG7lCi0njf79jyZdq9bHRA6FxjxHqZ8cU5PxuhRhDtDeqgXc+KELF5F5C9ouc+bo8jBg6Ig
L4uXhiTLg3ilewwKjGGFdUqI6SmvfGp20W3wteJds05aUhmirpuGj2dInOkKUzhrDFdA19/fuAsF
7Ml9LaejWKgzMupyF/2XbiM/5By6rh5RyyVqStp8ozA1WHA7L2bO1qWKAEhjgP/RGskGKHsqQ+eS
1MwJJCydWJr+AR4u57h3kA12XZaVKOjXMKgC9zsrz/nSs1XaibhXEgkeTsJ1A5hH+ODhNGvJC4xC
jsWn8mr22ttSZ1yMe885b4XRDCr9h1ZIAFryXMyAfIAan3S87cDrckLcvoJEV7v9GIf8Llemw/kc
g0iovC5RQ7T802ol8OClXRhupjXfWf3tzlDV3hMogVbf1HCKCD+nskTEBefVaYecgapQrUDo0jLG
lGF1p7qc9HaCgpF9MfkEo0cSgoJBpBZR6tmwk4OkdmESeLVbxfRfo5IH3NApWyeahj1YjrLwGL+f
WkIKNvcZ01HDplrbecUPu1829q9foJk8HfNmHsyCfjasxccXPO1F/95D8VYTcFQS3mwY06bMzmId
4agGjAlTiDxXHbZ3Q8zBq1zH70gIDXu4TnLwGOhQpODKAK8Bu0naSqin4bdVsh7+JZfmFRqEnHEA
hKcwo48QroH4np3o37FMUj3Yfd7fbJmWYuP3o1i8A4eqdSrXKcvVJYkWT9U3r2F/8D1u1+Mukjvf
AbikUsgXM5dvMnj9lHaBO8CeSlTeRXtGHX1NObs35rgju6iqqS4rRSVppdQtGPoT6arcADkmNh0Z
vAZZl7oHfDWE592xBZTNVdECv6fwEBMnKbc6i+19WN4LdyjQtliCOjPzcaYI4fbk/fDjmvP5N3Jq
i16bqdGmurwO2GkxKCyAsmI83s3oYebg3aQL5g5imkHHgkw9yDGL53NY6ry95XC2hHXHOj+JVJr/
keR7YdackZq0XttR7Wn5ukNB15LW2WyLklF8F1zaO9Gzk8BE75AdRyxv3kqq22whibLBAhyy7zwn
SXdY00KRBeX18c1KbcPaEmP8DOgMjddgrSKFszudR/otsurKxc4wBTWENMqvCkXxJnrKZpq7PYLg
miyimfyCsoag0U+Zz6lCjljlKPDysmIHmMzFFxmfy5eigv3+e0hL/RddVnJk6Kkc0RQjCxSYnMVj
d4azf2F4omc7ma4wHL5/DFDvHBCPMHtBLIOoA1omB0zmBfCvPp31lrk+C19haL03eixEeXeXp4+D
nElTw1n1050h9AAodMwhYsFYlTnEH2FQ7ESBJX8nTR5TT/3OsEcMQLl2/1M1QjQXtWCsvo+M7CFw
1mbZ9WUomivexUpp70TWIEpEIuX3jtnXXQmTZ0byNcE6gII6F4Ka4mRFG8i/88EiNPuAM5p8Iy8J
BqTbYpWHeYV0c71XKlPsgkFE2Z1SpOG3XfTzVowxRGFUawQ6LuY8aq76t5dKM0uROD97GwkssMeB
y75RFRSO7dZiPnEO0reuDy56mlqqTcG9cu0MTH2nMNVkd3NmXOz7a42ysm7LGr0FcootVE+rpP36
8d/Fbck4ji98Jn8+rfj4sPrQpi/FuZz0AnugIaEhiD7UlV2bUereVFgAnZpmhYSNmMtPsXZugahi
c2qJZ9ppuGk9oJt2ZhlFf2PhTP8Irb0DRc84S3IgSzkic/WibjskIFZyTI5dJkAXKVABgXhXxjqN
Q1q2lPTYn2ah5UDdqktfEYnx7U8dsri1Iz2mlQkQPBs/Hm0/whClehLmmff85zvGytkn8Ru9DLp7
8Ghj12nLGWT2jNSclifgCRHBF5/SAzNByfbukVeGPpakmNWwi9J2C36s6HkJvVEqFKj40cuNwYNi
xJlWdT0joX/yMHxFhniFSKrman7CP3vCrshZc1Y2CtIQvMr54IkEXyHfCFXCB9U1QE8A6t7TT6T/
ns81AIuL77zElHpwv1HWlFsXBPnZe7qYo/7lGqZe21LW1KwvRqIopbKdaH8hPQdlrb5dE5+fkKtx
Oyfw0M3ky2myZgl5hsIAesnVlQNge3yIBvXQgEPCROLo/YnTZzxRCNdT04bn9fvEpprylg4Jhgqh
/JMUnwURC6MGf/SHn7nGksNJRGBF7iY3BClqzpPyA3ioZZhPchVYYevo1c2cAry+0b24V5TPKhB9
5mSkH5wfNv5IobtaJySV6B1Yl+EwQYmPpZJwLzSqm6wItvSBE0GiR3yXqY8+2reshBxy38AyF9X6
9pOBmQ2sKB8IwZBOuhH6KjgcmhREvDlQU4kPn6fJ/z6q6DDSd6RKMihxGXYL3M8fW4WVUrSQd0XQ
rWdELK2icpV8ID1xge9i7GmT2Z+1QJHRYFXSFlbhduYc4Ryd0OghDc+4cbSjMgozcQcf9posQR37
+QrhewIylC1JJ/D84tZPNBIYLD0vvV3pitSZ1FpQ8pQ4+XAmmL84ceoDnZjrQVgIBSLAV++5jGZ4
gnJTqMZLFofM3C9pIT05rBsV26jYtNB+Da6paGEzBfHAu2urUDBGWIa/1Nt0eqFG6Pnd7IgnPt8R
sboNokYXWgKeG/lfiIdIF7nIXD+GZdXkt+M6BdZ98VnIWQbzlZinngoLGUsHneTVOPmT8fVz1/HD
2o/bXxlIZSgFmMr9MU2lLY1jSOqFp6a1jwJ9hyHQG62CpOaWDTLPRbwmEk5cSzX+vmBzTtCLmksN
TvJV8QpuLR+BDUliPrcTiJFcLgxQAUQikggXvN+59x/VhqNi9ChxhkB80VR7b5EJ/ViRKdSOmKWT
6YPzVmhj33X2G/K7lJsXGrBUxcT2MfmVV15ktLTfaS0rBu4kATabTfpdyCmY65Cnh5897Ap2D7/N
WftnWzxyGh4UWmQOJecA22XD0NA05tkbigriJvK/dHhnGY++xeT4hkJRtDTUB5tB9XWu/5U/5mPO
feRDNTXgEqM6aqh5sXi1eZbxnQf1yl2H3Szs+RQ9VNwhnniz9twYMrYIVEjaa0G0nZOuTR86JVTz
H/YvnDEDhBj9HZqLq9aOsd0uqVqcpq1Hu2PipjmqsyTePDzTYvHOgurvxt6y6xXj19rTd+b1c1dv
LKWCqnouSi17W1kzykH4Z6LXDf/+WisGEbD6KCmCE909VUKvQW/7tdBLsWJOzObyH1wpRigLQw7T
oWlbVugqowVB/Lr/qgXEBfK9JlsTBwyc3Lx5+u1OItOIOY3aznC1aHjiOLZNn5RGPybR2Y2GeIcb
k4rnlh6zoDONU4gRt830IQRxApPIg6/Ifhcg0nH7AvG3biZv+K+sgzCG6v85UaGxOZT5M1wtcno2
MKPeYBt+mFKto1/Kd3eTLx98eImm29GbTV/2NwW8SJtgbh1ElUjm5C+hUb14w/1wKNbZU6SGkUZA
E4sfmoc9HCkyHT20cvXvb8BkX5UiRMxEUPwlI45US1MQQ/hTYCC2OOXHwYh4uZ4WlzX+4NdFji6Q
nnUONYGdJKd8m6W4J6Kn3HNCD5jBvkXD+67UQQuwoHcQo7K0+8V7ogM+SN4wxMkMGRUk+fRgimkx
OPfyOi4lOl5hcfikPrekv27j5gQbepJpBXi02vcb9ZzSGXUMgYjUjNmhj7UbQXbxTF2alQTJK015
mmSNsrujrJJoUb/V6as9O/MkkR7VbA1PPR1UwPcUKEi61XjZeRc2Hmd2X6emkpmGyTwDbAm2mk7c
827z8CAgg/khhTKnFQMKjM+hXMd2dD2iqosySMLNwa7BnJn6+CDF2afsMKvvDFUBelR/6TqmF3cK
xRi/rxkPzc/wFxN1Nb2TWuNwKlOTc8J9ZlUbmkqrRGIIZHfgTV+cvoWcRrdzXlJK+jqf9cjI1/Sm
WA/92K1oZ7kofDe+T5zRDMm0/hUtG/rRaFJCJdgTv4xRXGLIIl3hzOR+lXf7wsrVXB5SjUSGSLJc
oEZp5bUFDFHBFJpmApbbvrrAzscoPuyYbCVf3X/inAwaiLF+ERRLP8jSEznCqKNjpWjV9Q/BMLP9
EgTLu8m0MsVCnthI4aWb5ocFsqon7cCa3so1NQzGKQdkUqSodizk2+8n7m5T+5s7o8z/yhugIEv8
iPPvAhTAfZkvC+LG40gWajeKVKk4j+cr0uL9LcdQLv9z+mJtwhXQR2WnJVqYeHD9ZGmik1AM1Ngt
VGGCABL5vwN6mZL7VX/g7fmW1Xvn/WQeY4kfnQfTOHTwioncAnFTS13ELPrupnUIG+6A5h2dRV4p
vh5llvJnLKZ1fzOuOa3RD7+9EBqDPrlvGR1sijuJgzu+uqZEX5QL5Cb8oRm6/FGMTx+BLStMTcHB
bSvBoox5AS4VDixBfbsIvDDujq0Y2mSRd+9HNkgfBEBZY/W+Q3uQFoLb9d7weI05KBFoSLe5kKXU
ry+1vbqzgl6tAXfwSkZi+jjV57usCxq9A6ja363PeayOzNuzl1E0inNnpWoeL4d+BOGqJFCkUyp8
NpSRc6mcPsUcuRXaNPr58bBOj43JKzDuwGzV/+ymkOMNGw1srljypNN6znXCLNohAoDEzgYpr9Rq
AOxKqOzhTEZ05vGibD35jylZ7eADHMfdZ3yrlyuxwLAmz6ZHet4cWmBB0wbUSpRyE/eF6614FwgR
4ARqZPAh4AtD8bQC3Adpnw867xNAETshkFUObMHqDvOqyVRvI0VxzYs26X/qVJu2pXFzyfKJM3pJ
vYYuxrCyvsxU05H1QTAaFTe3KaVnd9eeHBMe10gkT5HC2ZzGHiepROl/f/ltib/MSd8br7WSb7AB
2nvocSBmxr1VLdSsIKqEmY6edRU384zu/5it9B/wMg67wIm8RIKSV5MDsLsChtYnmguArg3zORuJ
zbIpME12QhpcahqU7SjsN1Gx9jBOuBhVJntTn3t779y1xalYSPDDAWx24gqJw+0rRGGU1vGoPr0B
27IM+rau74ofZ9kYhq0zCkXqjJier6E4tK5yh37hMvy1egKs63zuJ7WGFaKxGSFI1XxBjUB2Eeij
34cK2PfmhuXw3RiHpP6alOnpyadQI1uWnLTST+pyrGInNksNsNiikirkKYeG4weDNp0Raw4M+/Tf
04Ezs5msfVElhcOAT0kh+Ms28LhdVvtMrhmqeMGq3jlYfrfKoVyMvG/1EgHFbEC03IcMV7JAsvP7
u/zc05AoLpfg84JtPvl3ipgjYbxsuzRxxmtTeltwa8AVMcQilXhF+y10ZonvhSAdjHz7N+X/qjVk
6qYJy5j1qVi+zgN9JVRzeEKn7P7H1Z6Ub4STc7SLMZto+a5bA86zH4i/vdkztS5a1GPXgMIHY8Eb
9i/hF5ObG3hJiuhIOAOz9IaqxOlXmAwGdsfARQHVfqIykT0kwtHErJUiJ5b7guXC7bWzhOaFXUBh
Phk7jycJGHiI2vTzj7Tf8ZzzO2vWb7XCDr5SYqzvRV4wNPOHz+8At32Ee4r7rIwkQZhs79DBnu5e
M8dQ6G7r0ZqiI6RN5JXkE36rqEXfej/GXPYgxXVk/hZqPR01pPTD0rR8FPhL44ZrgoGrxN7bIEwS
rDipi9zxHp6cgqLtnBVRaIcTXO6B7xSv6z+5fIFmgPDueWOBmT85KURtKN8M1YCO0qh1mZq1RADO
5zAgWZv1nqtZ3yi0VJ1iudOo8PdBN3qvvBr4FAFzvUZ3GXR8ozXrx2DM/BwDwnERpaVk/fpcbqdJ
7T1h5wbyejYu8ejbV1h//YcBHHzhDwuYIsc4D00hpiQSQ+083VR+i8N3HkOld/g3KY/Ev5XfBuyA
URJ6X5dyhMCsJJR2ZuXMR7+eOZkuVgJFm9WTlT2thP4SCgGLX3sV51zOQzYy0QWn3zygNMP4JN3+
q0/Jk2eSzV/88TJXL4oHw+/QVzFVKXd0Dj6hHjGfRC8AdQtgVIUyeRnCHNBcccjfYOJI4TmpWrv5
1CVHrS83Bins8gmR7IICF6wBmrn0UpIiJjD8r/vCOvGeDW5S9ZJYw8x7XhJXHuP6qJPSvsJr7x1p
I0oGIw7DHlDJujq+etxp+MkXSmV57iFMucQla+s5Hb0vgrAvB3jVH6TAw6k+0wpz5Y/CZNjErxrb
pt4dtcfADpqJU0E3+LZMsttKdyn6qA6QzWW/bb1iSN1bSoUWAaeTD180jPDkqSxiQNZVRMGAShPT
QeEi71L0OSz346Bvrn+Jsp2xtm2J21wj/cbDJkmlM+0hSZ44lE51FmC1b6lZeOpXwuAAvXyHQt+j
FntBq+wu2/H48zDF3LFjK9Yk+7dZZuvQ4o/FcCaS+TMDSEr0WCncrAtXoR3Oqna0TDFnIM7ReEUB
W64ABIluSMPtwLoWvsyqJyCv6tbQZf+eBKlburX8CWWIUFY6Df7ecshAx+UdFyd8UJuLt7Ngvz/L
eWLCiIHfqvX6TgW4HlpM7/SCJ2LSsAFKGgG+/tQ6CjZES+a0xf+LFJXreSgaWLiPQ1lmehzn6+9P
wdgbXC5jMHbv+VHXfGCK8BoMDk0ibWKpsN6lpNAYlSRCeIMqK/Noxe3P6txnXUCgC/eBfhDsL5pJ
jfi2SjIVoJflfrUDEF165ayIiWsSAPHeTPzUUvx9l61qsPdCyVb46kd1dMR8tYH6NeN0+7GuVKjj
jOmudUt1VIsSA78M+99IAilScG4g+8lnmOrUyGqybqWHaNGbExo8jsNXkYmN1VXUYakAFWw0DWmT
zlwRFlJnh/uEjMuE6msGglFeNeXBxMGKPgzmgaLQsjB226Mh4stT8ackFv4pXsgYxiewipr2J+3z
2PhACkp6/Kk0izUapIru4G3IhAmypyQZiKECDpEKtJWNKCBNqyDizRHLRtUs74sq/9GMC/HgERXu
ZyzOLIu26aKY0UjYCgKwn4HXToQL6QI8Ondjx98BMBj81Yhu9M7fJ6aE9E1fHtjZ2cxMwfHgi/4C
0pFXoZ8TqXFExjy6H0MjnA10Dw4iNNRoltgxBWHgDCmo5E6dk/zz9bUrYKZ2D1pZK2mY2Y5Txoe1
sC1bPazTWT1wcDKHgdhCIuwKhd1k55+sAOfxKaZDvP69pYcFCDouVNifJ8vRpt0VIBVOs2at+XER
IQplMeEK59fMayZsRqDepaHgUo4t8Cz4r8xPdxinD24aUx8SkPY1PIF8nrlj+VaJ2HbAhQtbqsAu
AEytOn7rJ3FfanNAXZL3k71bd1xN3SOUi3IPKv8XvgvdIY1UeOgk1gvZy0Y4TPybC5jslnWVeI10
cSEL20sMYoH3aeEcXTTgmn4QniwbI39qx970sJWYarXoNBht8u0UVhxaapoJjSLGPNHJjuIMhi/9
CkYbJbG4Gv4S/9huCqkPssObCt5seqbtp3bymw7NBNwtVQlhx/TsH+KB+WHUBN6QT1oAHii3bcgj
1DJRl9avKzLnd9jq+DxnYk8T9MzSmg0shT0EpKdCyzYXL+uEp2WrsTfmw46XpzW2wkscZDAsF3mn
5gpNOPxJincDTeDuVZjB3KjZPD/LV7xf0ihsdjEgEVOcPT1o1NUBkFddjOcbAyLkbFdUgysSg62a
TtMi2Au/NdNuOsQa4wb1iWrSttVjFDZky2homyiTcXReYbl3Pt6KxlcvBDYKEQSZnK7ssB9hNglc
/oC9rbpsDfR0/zORBvTXBcg79pLe29zZE4sUlNLf2iG3mn3/dhxMC1tHp7wpOMCC9De5mT7KeNJz
B9HRvBPQPp3S/pgQUBpaU1gBFd5LeofUajaKnn2HnYJVxP6JZ9eptO7nEiFeQIexT+5WK199as4R
cAU7xUnuf9c9pYhrUVTyrqnoHdthD5UPAcvYPnV6yi+59p/DjDvL1GuTMNHpTEOTRNkFi7oX4kQT
mswKFFiDa08/6ZVTFSKtdZswOhJMuKy3e0uDwoeGfMTQxezCW6Y+xRVVYWbZxTNTADsNPRx6X/lj
tylIgbjBPAEegGTdJ9mjXzF/X25pqmjGHtPi0lta3ZWMxVCP6cFLNBVAFD5hs/6YT8ilSTzW2DiB
1DSYka7ZiCBr5QPUHw9uU66Pbj7ElmxRp2WWtjEGz0x71LeSe1CXTz43DFd6eZ1pZyv4URBGZ5KF
juC69wRYh7U0ft+eGRsEaa0zv5WXtRe0xW1DN2PMqcGVL28OHc5YJ/j3vHVAizr2SqMWpvq5G3dY
8D2F7Rjcf5a9MI5YLTwJjebGewT070ZXDHCO8UVbFYYMa89Ka8ztKaohkmqJMQZO5puQlaW4iGtR
b+ClhFbyO1y3QHJwctJ32nDm/TGiU/OXONuzGMez/JvkT0hbDTRgblbhwDaAK5rK7/7gYIRD9M6l
DmR6Q8CKppd4VQJt6OSKljikoJv5ASNnQNJqSuYP33yU+gJxR2Wu0dYR7pYvQYxf9y1CQDdM4AwC
XX9CNEBHzrufuqWLmTI8mQzPPu+VjCKkAausdjpF60jgLrb5Okw5bSzuDjhKc7OWmblCWQUxDXl7
/rw8A5Hqs7shcExNAjDdM4L6Ba26bJJsJ8UdvrWUnuDOJqUPy7Xv3JY9AZFz++7UQgbtn9aKm/K3
Ryk+UpmdzZNDfew0foacj+uH0XY+28i0S1AEyKnzNGy7zczC0ciz2KeGFLHDlIGVM7/ZayYUE+ml
9bfI2s19XBbXmpGSsoqYpKundkjQY3gc7VWLMwxxbpTy28Q0swS3PcbgIALZEuAQ8CJaw9h1YtGm
L4VCFcaTjzn6O7Z8m+rZK8Pt0+isRgYFLR+G9/55FVU4gMXszlryPjVDCJDj7finevQJDGqU2+Kl
t7mdjQqLQuF0O3Oup5Uo3cdorHwpSK0rLNK5lfoAtuUvueGl+KYx9nBjUo8VBnuD/4szw1mLcor7
EhwVXwVVEA2ufYYUXPNIoNyJlZ8Txgaxfa4AgGswXTNLUglWhxqocKjbTjJEMUPl3htwf1OAJw4J
oF9KwlCPYJb/LL91CICiJF1onYsI1oX24dFuXgzicf9c82IDs+l//h6Zzkac+hYnLxXAd9GqL9t6
ko05ocy3PUY/Mln3b47BfZ4Jyre16fJWh7wR8uq0ShMyTiK2FyPzQvlZE9XBJ5FOuHjK7aLdLTyg
0nQL6LDtxk0VxP3MrvyhGxZIjLCAXwMSzrtUvs9ZozBVvGCfFiAzsRvbSTu8G9CpMTcruLKzwGbV
7D/6COzhI6oeRPyxX6xVO3ivmuNyT/P1eWF33s3vC5kBMwqr2kUkGJM4Yq/TgEY4Up+tURcgGlQG
G2fUfdTl1+jHIVjT/y7S6WZkRti9VdwLqNEz+EFen59E9iXsH8yO41kCsXpNvfR7STMRxzdPlKv2
4nvwHnXnu0dMGD/QAq1e5cLfkQ21laOowrPaytssZghOyKhvFWNV+l1QuNl2yikXaxAtdU25edOw
n1EVWoNnG/ewQCRrt7v8TbyHCf+NaSBkcno8CfEOxjcnoofVaJyRNFLNjKb8WmiT3BFZrpfCF0za
ZDHM2E1hh5lfHPU2Rt4jQ+YrIAC4v+3gr99LTXyJWoIWK0grPuETGQSmITWyKdpdp+Fe6fhNe5nj
IJjsYXYpRgqzhQ41d1pARx7fC/7omyKW9Cz0ZN2p27AjS4H38PROe3CsQsG33DXYwrjGC/fG0Evq
kfqrrmv+5kNQOewZ/EoTsgOMqftwUF4yEG7eDxzaIrtmWlB/vORFzf75oUs+DdCx+uqXh0Kblqv4
ndC+pYmAFRZlmsfM2ALFPqsQ2X0/xcC4v6FQ7GYcpwt49h0I64YKp7LhTrrizE7GDma7CNAVe+7n
jCGE5utyTh0g2hFmHQWBCStt22dGqaUtYrO+Yb/L/aFSp1iQzeFjgSnl+At2oF8COi2A2SEwcHoY
RHS/DWvGcNfpDFdUJVf/78OsPoxgkqD0LCUKr9AK3RBois9mg31rF/KN4Mc3vm9k0rcTiPpg/1JC
eZsB1U83chzWVAy3PaF2Z8/seGSNw+TvWgCcW2HWGK0RrbzLmRZtJmgy/4ntHRlJpY+KgaULYV+k
37fJgut+gc3RVWPAbU9/5UIVzd+nMbB+m1T8H2SRRJ3wkZ6p4wah7uwdHxAx576r/QwT5j1bw4kZ
Q9S85qqnhFZDCbm7QLhNwoblYcHRBgF+MHmWyszAJLX5A6+NSG1YWTPcay6WvwToJurl+wdJR7Ql
A9aMrzcsc4MvmojyJMs2fDkcjuA2m0KtvaCMCCSDugjfm8NahzxPJIt+8ol4BeUXyzJlG2ncaGLB
oaZuR7nhKl7ENS4Fw/cOZuRiEX/OXbdAGmY8ZxuHXadlqZ1coIc/tkD3e6BNQ1g8yACWOP9/t4p+
ZZkJAqvK+3dAnB8ebEPr6rBDpyBp9BaMH9zBWdl6EXdNXZW08gjwxbdl6ClUTIIk3bFuyrInwTop
7B/n/B3mr1vc1fn5n2RbiCrdWYoOo80w5+zu4ye/Pcx0IET4/2rcLtv1Rh4gam1kUbd8Eqpgy7XG
Yve6nPWclNr9N6f7qprkAAe4P3h/zq38SP0Vh79/1nKcw5sYJx9FFRWYvN2Jof+EkGhZNfgZUcxd
k0l8OKFrVr31+PZoIZF6beP8F86mJamwmSsKHAeNU9J5z6BXtGqdHuoQ0RO/iLpzVMwmedwMODxF
b4Q/+t25VI6bMsJMFiLcQfVLQw0Gb8ay2jriX87dcAjO5e0duf0ENmsToin+6NiK3T572sJmiyus
Eg4bSBQgBUyL7NPU0T/S2RgsiHzWBEKcN0NYGyeS4uNnZ8NmT4SgVQ6lGHJhTLCk/JDqbS1SIYx0
Ku5FePN3IeAeIuWVpan6S1wDxvwlyzQ8glI+RChhKSga5S6HP2LGfUMjd4dd1BZdD7H3EY2elkai
Mc/OYrh18sl3gr2po7pYcJbWG1Hgeu1N5xslBTADkMYKu19EFj0xzyCMaDPbwhRZwU6mCJOtkGsv
FWVGtGHtLNCWwcUPMm/1eBSK76nCrX/7/mdcpF++qG/PKqgdWeYTjIZ3Z2XDQ2Ha+Mm/ozacek7l
mb2wKIWnrQ55kszHsfqY1J2k2dKFfzpJO37owpdhtkPrJVmp+SCOq8V/iNkjESVUV5SAVlqea2tR
OJg6kaHXQyc5m9ZD7yR2T1sDbzr+8ho09hNcI5EnrDAlIy3OsvuKNKHniBbJAy/adBPg6t+s5GNE
EeVlTzoymX9vWDYdl7p1XzBoq5KSJl47lCeksTK0RiqTPEuhh/YEP/7pJ5DXih99bzjDcf9y0ucp
s4upLTRprnySXWcPwL2UrAcpui2+DJ9lz/gpmZmRPs0eN+tYXeINxnWDKdBV0hUuoIcnDaonPAdw
Je6y3KwHxm3FZ3eioEw/TtSBsfvdmnZh0oPNk3sOb4eWQ2GTmxVgu2nraTIPmweusfOSKPZH4dwt
OIyFeSJ12l9Ty+qVlocre4+tOuT+GJXFwEjPtEv2/26cxFe4yIUAIdep3Ej4b+Zn8RdtGEXHx1Mp
dP14JaeHzoqMgcF/kIPAJTvUQxSD9ONvnbDuYYj8K4HiHQ+/oPEtlY2kN1EiAUZXXwZEzAhQDPss
Djq+UFxKtWpVp+xB+i5FSvywukZNgqRfiz39V5kFaYjPnzp/QolbsD7DglaN7nZ1KJQLjcbnlt4E
L0Y35C7bI85LhRt35fflYH90bINbfMjqTV/+YTuXwMlZq2IggBD3dRn4IDoBIUidvDVrX+6IvKcU
MCp3ajPH8eFrhQHC/kvyD4VctoGRGll/EPRSUNMRZWUvLMAjXifzBfTG3vHSWqcD1DqHb3vP6aWN
gb3H4sbldV6MGpBzl6RBjXkQ/+s6J5ZrUaA8Mt9pmPUV7bhygRGVrM3WhDkdyEIrimULB7Lp3pd0
b6pXKeBRTh2PO4bNRTASjycO35r9EPNvmGe9FCQMLy4lNDna+Aknh98kBTfsRxvuawIa05/0x+3v
9k8EweniKnG4/QgHA8GDs5xjE6IJaEczxOqVLcVtT3Tyf/9k+fHMD/yll7Oebm84yUNuF0oafkES
8KTH6xPzrSjgTDFXypWat3poS3kYyl5fRnGKVZmLPvr/01RyeJeTUxTVmaGi87VyF75Q+AE75jnC
jFnduXgXG8w6PSzkSL+/4Boq4jjKPvMJUAHRM/ptCDT8qlOHDfLAQrrC1GLs8hM9khNcyrjej1W/
pHOoTvtm/yfeGpNRfS3Qwi3PLFALrs/xZjmbVZhKAxhN6jMPCBLSognNDu8aMm677oXugjK02rYl
+U17oTJn36LroTbdp2rsDfLV2n0XMlZTX1pWARTwWfSK3gatI1/H6lLLr+zAbypIzKLbkE1ZfBL0
RreePSOWNRmPo/8sUXhr33bcfZMgadCVaD7Ih4R+EzQkGw0PUXNvbEIJjkOf5scziOvQyhiyTO9G
9LKUNqGA4BLRET55tgZPBRyaVd+gVc/RKhxQjzxdIo9/8ar1HqklgMFpEpUpVznsOVo3WmQZ5Fes
nZsrkcrpuuUY1iA0+hLbXMhURi8fYoIWyevEGnOsEgh8n9J1ME93eApiFhUNA5WFqs5RctUzmx5Y
9H8lMnscPOX3lsXB3ew5QxvP4xhu8dmcK+QXz7e+trkJNx0CXMgwsovVPFGUeqbA/8pJkV5n2A45
atLgyMbHSLv6VFfhRhzTKUv6OXrTShFtXU/kacnMY9oQ/0aswq9SOGl9l6Hl0wR96KN6sH+MA0+p
f2CKJlbp90maKzfEZJ9+CrLY+c4mq23z1lszp057tqQfCpnlMEFbORdYYzmSqID5lpsq6XOEkgFa
B4btBfmhMfmI5p/8FFRPMqtZObTeZLVuq8QOYXb58xiz9UIZrzpGzHf74/Wk7ri0WVjnSwFgUS5J
brk15eL85TKvMgczkTDhVMONE0UwmSJIo06AsLb5/eSUxTjliGNaBjgwrrqjNRXKP794+V3OWvzV
9WtGoRCyGi8p1pU4EC/tcYNxw9w45H6YElL5+2GG6LR2QQ8YLVRxri5O/fsUVhm4FcZ2eBr8xf6v
qWmBYdK6Qzdo53NjUmnVXyUWIhsiSuEiQXLpU9Xfd0rfSbgCoC7sfXiPVJoBw1ppt0zZFCCeOvgf
jqaT7Pmm2O34ko+lbJcOIX1GkmiZwPNw/VYMxo7b+p0P5eOah4ZOjxn++pHYxRuUrrFhHMVCz8sV
3K5c3B01HyA/Aq3p1D5bKWNAJ5e1X4JWQvf9em10OgFz7nFC4r1v7TGMD2FPVZebUtu6/Ro7o5aa
b+Pm1HnOBL2b540DFdf/wZHei1rA/hDe/Gb6crbWkXOXHnEvDilEl8mr/NK2CIRA0h7106+RI+GU
Du8cxM3Pl76gkWXQub3YfZLmRa2Pcs/cB7WZPuqN5pjt4HWjpwVuektiMCIyGhsceP+kSvFQXwGZ
OhDJ3D6CXk0lgn/oSuA3xk0/MCWLitSHLY3X7aOMOc97U+yYx6uYw98SuoZZNyMZ5oB1jdoQgVxn
T5t/ToEg1Skh0+a1ag6Q7hbHtUJ/E8RKarq1CAviovTed/FkJ16OMv1HOzA2UZHegFExkcr3W3hM
gkNc7kmh73slLLCiC4NSlqcgoD3eXQcPncmUDtTTSo4XmNPzRbOSOCKDef8eAfVdy60yhSkjDjip
9Go0YdcJTHqg8XBm4yu+HIk12EmkfgD11JKhHWMZjz9zwWNcNAih5+dslFaGPi3j4zOj0UA5z+4l
DTev/aKEd0znerT7DG5EGlMjN3psWZqSla2D2fMjy6Bp3ofzsFUUTbYH0cMGiA4LcDz7iQE7lfBl
jBx/lR43JlPm9rajNOtIIMZ9Xsy8xoEDJZvx9yetOZEyffeCxKuFsNO6saobE8s25mON95hh40F4
rcmeRHkdwDBLt/IQF62rUuu3qZE27dUV27pgdj5xPebCsqFOMa27zg0cEsuCp457z0vhMq7umBL8
gs3b6A8XsOpoXhZkGOyR9LUKtZUn2TqLlLPK8ODu6EOjXx4mcN8VI3O/CGn3XRbUY5sik8Rb1BwX
3gP9rOywaT3txSjrXhIQkmHE7aeHVWrtHJx44z7g1miv2p3UFdrpfKiPt0QoQL5mlL1CIBu5y/nW
dWTntN15q3poZYiNUt3yQOBSrdbzjOGASIBWAOhwbNwXbFlwI4FhyIjVM6W/8J6ED0xDQPBcnUKS
ISw7PupiDKeqYxeEZlqy2bl0A6B0k6f+hRKi28SoAefK5RvKkOqoJx6xcoIY9id/e6j6xL4ztjfv
4DXDlCsf8S9ZSDPFhL2AJTD2XS0mhfxZ+XM8B6a1CH5o9hYvIUjK0AvHshOtnR0VOaQfG2JGrh5p
CvJw1ja4ErNyYyj+sFsVASAoj1KQRnKNmhDEmQyWoPdme8EF1/nQHk0dWHQIFwc00pcjkLd36VVS
6uyYYUQmf0xd+9L42C6NhI3UW1ckkxumU6OfFUcUHhDut0tf7niOvzJn93oEx1hsmE2FsFw+weP1
TQ8DksKgBLKe7FSn+558TizN/LrQfibujobtY3feUwk/4eZzFuAApPV0XS287xqKdPA4uNu+xilJ
Js9CRBWC7to7aER/l82cnvxOGYoEtVNlyzyG7BSU41gPEFVOuXpTnhg/0eH/QF+mBMw4iUzlJ5J8
d3s4K3dGbpXg6pIpKqAsUIC70uubsgcwxVAFfZK6UxtwhL92uZ9E48uTiCxhapvVL94gImophma8
Huykjhex27AVg10U8wduCTmeVMS3ZyjjXPqdRjCtEDz3DKGeGgV3KcJU0nkJHioO3A6pUR9Oc9dh
CYGsYR4reFWXhxLdDdwsAgoxhYwFMsSd7YjqjK2H4VIPTnYyEWWme7+CXCT/wPxVbhwfrOEoDFU1
g4tl9psNZwrCnAJoUmR6rF75iDC/bYCFsqsumNjK2kfBPp72LgzCDvHNZh5eotGAcKkB75rn1OI2
+bbayknfP0hcauy6shb1KhTuS3PXr3DkL7EXx2H2cBNdXGg0YmaUGhNGFeKqlgxk0UJYZy9KVq4K
LO3mL4B0W34UjoGsSVXhS7IRL97ebSChTi4gRkFuIDlyMp9C7qMV7SfkEC6oGZ9ckJrWX5NUeEsD
k/3qyC3Tx6xvJWDWQompqRsvcQqnwJaeHad2OyBj4Sw2L+azvc/PIzHVkKyLYJr/sQy/l45eyVnF
vKqX/QbYXCE4cNw4+T0geNd01SlqN7x5UpwjRES86uvmynSfPgDZLCBh7pZ9MBYCsxtmfSr2BkOk
1n0tbYwwCm3nPPizAnKihhBF8eUBEUsit0sOTCbhQwUHePiwXiovSaOwbePT3ELA1wUWgneEryIS
HUKXQ4Qq+MAzwsTM5HdJJeUk8Doyji2gOrDS2F1ZINKUNJHP96otfEIk56GaIm9f2IATUYudk9q/
6+iFhz/CESLiNuFISidotUvLLJSkTOVKVp1HpRaKmqXpBh9Evo10I3oDGXJG6bki8elaoyXz+qAl
rFLIlmVfmB9ihOmTnqSqmUg7DEQNKAueDBHOzHtYYghigcb+uZDTW2RuXWWZfL03qF4LwxS3TVUL
JM+s6mqc7eNP06aGdKIBemfAeTo08qgp2UfyyozmfBMKbenV84Fq8jUBnuazZUislv/VwqP+fSsS
cQHyYhun84dlmchDyRJzkpFJAuFAh6u8VRsJ9Xyl7KD4FeEHvv2YCfCwlMdy0Yb1C5evFqs7U6cS
9e6X+GocVZI7dM07sra+Tli1pWuyYcuiFfKP5QLFEkml6pccaUAAEfq2i0Z6Cg/7j17RdzN1Q64t
6C7jbJnJdvXFKbYwsenpIY2ntzXcKUFxSdvo3FiLyUgtRuySL3x6xJ33eq9YXn24OPTDf75dozQ/
aHjd9HzJ5C9fllW9prvchEYT8VvowFVSrYihiE/+o0jpLnDv+1b1g3vkEEYyMUQAoq55BgZO/8tH
NuLD2rBTFOn0GRlueTzQohs59mvq2hr9C9hztrp5RYTDwBxb09SNxpQVzq1gwEmO0YL5zNqH/Nn3
05flPc/MPSDqS2+AYg2RY/RcIjroEcnuRa69PHckicQstfFm0JyWnubpkQgGP1KhADh9BPP1BqDh
Ny+8zOpx6RlFYzi5mHkNmKrAhmi0RNctBCFJsDN9Jgio7rZtTI/A1xhK924WgUo1UMBH17eH5ORO
VvE6KRdA+hIoJExGH+pxNirwz60+Ub4Z+NmIs/oe3rqp2qKcwvmFDc42LDsMqzdUfQZbRfplqFa6
U2cK7WPdUi3CzFihc4HSg8HfgVZ79Qa9Zy1mtoQ20EoUidfkifEt6G1chwH+5CZPtKBnFT8q3FWZ
0Ti+oDzv8A8tZXBWerqZqoSj17U2QP0BaO/iO0XToHkchKjqWSAFZT5+ny6pj/P9Wspnti4Xugwv
JxvkrSTFLNXwXx0sNlmuhdcXOquq1NO4y4o1kgsKP244rtS2wRkRKMhligJiKLwUP81tLLeZ78To
sxZ0j3fr3l3gMuClr4MSVNZjjaawI9tLv/1j4xmwOc8DzKDWTBN2liXX5YecBV8BoUsB5cTAYY1Y
OMkN2UaDx7jvIxEOTS3v1K0w9DtROjSG7325nyi57oiqZvYVO8gktxbWTHbTJzy07d5gfwgF7XrZ
a1s7Fain0fkiGDSKj6aU/ACmzIyWY0El0JT8/JTENEYf2vTxCbPIjOwpNbLv/h6+XNxGWLq0k79j
Xi9pVe0pN7ixbCBf7ZrQBGRGQm0SGWG3dtCcCPUpVkTbmUci/gDiEbDNnxHZTaiCb896Ugj5FrJo
nc9xZtlBnkRw9mglrzQ2P3EeNi2COtn07wSMNIFjpvCXXDpD8xWGfGOJ79FwHLLi/WA/oQDDflan
uu0Ir3s0SXXaRRakVGqSWyXVU8B+hsTsVe7QvmXyFcv7dmssEP2o4q64zjGZYvqHiP9G+WlWN1s8
M8LHqjh/A1xeNVAAmeMutuyUMR/+sZerzNX599B+eBO2eiP66CDEzdB6wq3z4TXSV1A3eK2BfxnB
6PIfobd3x0qlT+fy+pUKBWGD8C63dCD6VW4JrbFQCMyE4OJMZ4O93WnqYAt0Y66FOVpX9Woy6KeV
TMDCoy/igdNGUQIAc77R/oJF6aFThbHAwnXGMVZwaPIHynz5Whs4RtTE+e05KIqd+W7/HaVr5cdi
MXoMvSlXOCVYQOKhm9irhQ9cfq5akuFB/dhaEYElWMKjLzRZ4q/PE/qkJMuV9uNsslM4xda4VjWJ
qhHLHWVlqPNldnYNTDDJBoBTeiKINvvScKUom1oklw9CYhabBEOHlCN8HEEojOZhLm8GO6cSkOMc
vOuCE0jhSwfgGc7DWKKwhp89UB3TyCvX59rLrBDnYehjx90LHnFdlSRnfLFQKMvPrwgYchhdW/X0
205W+IrBZ9i7rskZpuduz6CAriwzhHOXUR/m3Y0iCJrnCCUkXg/dw6ijVWzIcYPiolapNzn1AHfp
ya0qJyxlUyWdWxPfujmNEfTxrRaawkdAeJkCNv7m6kvGBAeOsCMZXpFOjl2W7d2JcBL9fBhhyNxy
BCh0Nuvmzpv8GVDsDKAmuTyS6IKHgSAhVVB9iNb2e5LbhZ0V/cuu0VpPImlFOUkYzr/B3Ek4mDY9
+xcRxlb9FdITe3lbKxAkZJTwYW5soIEkZt9qZXt5Bi/wOVWJkk7aMiq+E2xNKxkYOY/cwzQ0L2wP
R0cp9L3Udo7vnv0bIe5xGWLrq/Y7ZBQFmMCRRRe/ricS9oVoAdG0UvNwtEA3tQbAOyF2Z3Kvfxk9
KgTSno6J43CmndvkxO9Yc5Cd4DrUDvKgxuVSiux9HgAlmNq+KRB3TdJ0RSZkLeWC0l5maFGsr5s4
gy1d3sfubPdpF3Cf50nJZe43cEj2VErTUVZ0DDpYgqtdUmh6WJ5qSrekux1ymwR8YtLQUEomzoYu
W+JyoAjX4Z/3uqwkEREDcJV69hacFK7Y19RI/cu5QDW3wAqcwB7AcZCPFhmu0F+eVOfsXWyRpVoR
gP7Ul1yUl9sqZUFOMH462ZO8O/G5MQpR71lqrUrcdyFk/M1/AvzT14mNe7YkFaUCr/tWQO8792BU
2xGXOV/3TesHDBREywB0MblyeobCiANu6NwDuNl8pn4qMPIkd13GIJppGnfeThtdsJhtVB/QWh/t
61Cw540VCfVYODGnDIZuOXwf4vx8dywQVj5gaGnZshCj1F87iTReUf1eveCuxTl0PyHibq+VXBuQ
f/JJvMDjsgbspUcwwnEwsjkVglM4C4tz/pR7ZZjwVa9cPtCNx3RNOoYVrdwqB/O+ZzcgMpzJtgvC
kpifbUDOAxJJ+qnpvh5oGRjc5ZroTZaeVHkZTv0fiMaGXa7JUDBfsr14oXl8jeSc+hm44xlN57BW
LzTzTgcMP6tK4p092SEpviPALuk9L5tjRmn4whOhzHoKM4IjOqfx1EWsiijIWaxlGrksZ9nEaolb
NF3teyO1eCCS7SS9oXi04QH8WAMm9TCReMrUnwMLZ1suoHP9zbdsMr7i9YV5jO/l3hGctAEOL2hn
JWDNTHx2nM40cSln5Osp2cv5fbFfciNYqK3+fqSgHL6WVH8rN0gyQAnIcX17qV46lpMyoaN4OjKQ
2Mx3mh73zWfPfsQIDB+j5uDgnzYex9pMHUClDAnU9JuBlpYSSrYHDp+MtbdWs21AXTMyxKeFiKXj
mVqUMABko/PGFzvyq4kFkfAneFZ2QFAM4ciE7HnWqoq+4bucehduEDI3ckBZXHVVQonNEaZWokzA
8ehNFCrMDUHpPs/thy/C6ZX6LLA4xhmCErtzQ++16jeTwmsOKjxBY1torobJkvzHDieNDpe0r7zI
+lyTCYNdnzV8NybSwQqBfjuqi4jlRR9fAht602a2CJBJg4bflCfNjpYvhmxcX0ry/6gYvbxOFJ6p
2zVxQylwVRZVRu0TODPuCbXMLbUD/D4sKuh2tvA285bRHC1+/Tg2jYo+dPiCZUom3f6DhR6rjFjA
VCbLO3RfwEFDBHkUzZG4Ikls/eypeLUDCQTWuqMUSUd2UY2/nhCsJyVdkrTSDovqQNon8WIdFJtN
9JC4XPRIjfwh6mVtSsJy61o6emawhRrmwBJ649uPlUogFIv7gtbSpFCcj9l+fS37/LT0knUMQyCu
1zXk8yFDzVq8cGR6flrmnJ/bFguTkFmG3VMdiuR9OvTvo1SA/ik8b0GsmhFsUZu5mbNID0Y1AWsV
QV7K4xtbvMa24/vlIfGRI59SwQVBO2qL1ez0+PcKWoSY/Ob00+Ho6tJYBFcYKRclaTySn6uAF9qO
UFV55X0yFLwnlVqXySDzyDk5YJrI3u9C2VgeHFemoBLkUgjVlqoAlVwZQRui0c+oKjcSx4J1V++4
kDr7fSJjnOHn9BFa9frE8B5LbX2+fuCDXNi5U6T4TwijoaweqEVvQsROvV5nV6Cl+IbvVVlmHxSs
VxgLap7sZNqtx6ztOeykAxuFm3HkRfdNq+pp+pfJA/0RhuDZnP4lbCl3q0kbJdD01ByS0oxJufH/
mhhbAvAhdnTvOdczz0Kxy5EAOPXiy124xIvqthqbjRXPQdEdXEXOo2yl31vP+9cYysaWHWCPlnps
7X+F3Ilahxa/6+BTHzFv0R7i8qycu7FojiI5GVjf2bOcVT/Y90iWkTnMAjztd9S5ZTDzj7lXmzVb
jW6jQniF20o113tyVRczGnyS8bk27/0IdWrQLlvsR4NIj1HUx6DsUapF2Xj+eMd7btujIZErlc5P
uPFDc2yaueLhDGcTbWAYgoDFEM2oPHSYVRrSA83imVQkWZm4+2Wd4JkMUXR7c0aJDqRwVHzUjkCf
RNbzFaV66ONzPEHPcvxWHsG2OrEXIWSBCdVKakPi1cY4PsReJpZ0H3IhjfRAkcKbihpYU9dRWWWW
z1n1s9t6OT06TG1G8otUR1vjZROXMR8R2XFFSYOYkXUdwAzsKWXGeR56xhMXlbyEjE7WL+RfI0ix
70w/sBW9AnSX6IPyaiwuh2ve05jgmDaTtGpY1pEiEkkHpi6nIPG0P3DQMsXuaKE9gEd5JJfyzkdy
eOPRw647NUR0XLUhtoO9epJLgZb0ywQ/cAUZxspbNVAl6pY+HcbZqQHbcU0SamaZeLAE31Q5R5wk
WqD6RF68Lfq354Bm+wqJuokf7Cy+uqSn5QSDoGaP354R1oEczU42z/rfjeo9iylTNMTLivOi55U1
wXCB46jWkELZRFHTKwMGizZCma5pFMKwN31Hpi9dvvlXEMSy4aOM1NpS3FSctYTwQgqtvmlrXT65
60uYmlEY/S1MHJbeSyP+mVZkGzxIXUSmVp0PlPGQLt6WO33KY9IUlmloYOerJMmPcncNKHqDjZ9X
DFOG6UnoWBKkV6CdsLpGIVUSMP4pM+mQM88EFJR7J4lknhIcwQKzqpg5B85np3xLVLHIhGUpg5Z6
xViJS/xlbhPE7fq31KU0y6LsNWEAC5OlaM2o5A12u2XPQrI9EHNgqpj19BtPMLZ+mdAREfHrrIBv
hC4lYHZ6FDELah53SKeER3jm1xQfy43W2P9tQtQa9tztrHlHFF26DJ8LG04rHK6MpidemxV8BKd/
0ndCXvry086JoyzVftBQ5MQgO9wNcqg542kbvFSMbTPeHEC0z4NidAbfVFMPPB7qaXJ+la5ICqFS
ponwZqoOW9e7aLXE/XP3ga6o9vVu1npwyTRva5tSnBHWrmbZAhDC+L6wljlACQK3bAb4BnHVP0e4
LNZBjV+wr/3pAgAe8BgB03npfTbLzr/HNMS4A1Ot/+qtByAcu64qyLdYYar71aeP5gcYYWnxeqmD
Ny89gdhca/I2LaJkgsx9CD5kmomT43aFbWaNnT1X7iB6ftW6Fxt4FIpsTEmqI3Z71pIaAFALKGtK
SUhvEwDq2VHStuH9I8rESXks6jbNzKj46Z8xFuShQp4wesPz7cKT+J4SRdGflOeqx85a+h6tnXW9
zCNZpFCXk6AX1jScHoBXBVh7WScTEgarbmY4ZlETfhc+gy/Z2+rcMgQhNqnTZWP1aaHKQh0Cbu1y
FE+njPIdhZIsOQAq3dAr6Znua2lOsQOlmecxtqRZAGy5PeopT1GA8103fjaiLgT9kJ2f/ya2AXyz
JnjKl6O8TJXE5mkQtn0vSCJ322keFqW8jtX7Wc96T3XtyBDEk2zRTNJJPICtY5osWVN5umqkswF4
GJ5J3j70SuEw3DpOEzvOBS9Fqw89fTSZ8LXwb63VcQTxAFhiz7U+v9M32+qse7iXCv/0A1pM2XOk
W4e6a32feEoamS8KpHXiV7Y8c3rkgAlYffiszoszuUbEwKYy16F7QrFbRDBaBZ4FUx7Bwu8KNy2J
fikUhEbhywL1MHXhyVZmkB9OTJ+VyHDIEyHvTH+m8OsiwPU7JlLd3rGxq43oQhXa1QrjtWmQCCPw
jiTFZwDCIKLi/FAHeLbQL1KQdwnQyQSLN+7AW52kUWIxJcoIzs/OVIWMfSoPanV/CMOSlEhQWXB+
9RNdMgX0EqytGbp21ErgDue1/ekhKIXL4QCuR5FRzfbFTGKb42IMuRFxmZU8LO1RTWN04xbvdF9h
l9vMI/CVC8e5At0i3pWFn1Z8HhBARZKNnGo/Bz7fbJ19T0w+hE6/U8b7E5craR2m/R7wOZm8f7oq
IwZoah4Ph2w4GNgfD9N4S6pJi+RtO1L99fvjRkQLNF2NRsg3QmFVh6egfrVGgdHZj9CVg/gX5BnQ
64VHVwiel/nSH4phttNOHUE9MhEdEld9ZnEsLMzmfIkog07RgHbBGPTG/7YIHEmMQgFOWh+hUSsv
HA/LDWVKcbOlL1/anHSUWZLPuTzU0uZ4f27MMSMcxVaxPWIkuYhATcnzbPKjaZBSG9i7TG/B/zrJ
DyToXbRJGnm8Pk6XyXFktQBz8VQR+lbW/iSsJNZ5zZZXQapcniEtO4mguooRWailEOp535VDLKXs
GbTRDx4Wc8nWzIxs6ZjBOqBM3SGd0MHl/3mnuhFDvTtBPqHzc79rs/YeTXJPvyxIULZACB3eMoAs
ahz8yTSGwfU40rfs9pBiDhDlHXmtprkM0jtHjPRNDvA52AvsZOW22+WHiHz6ngInG4LozdtO0Pd+
LtIusWzzmEg32lgQ/Uxg0GsziedFtRC134IfL7NeaTvJ7nYEuHM7VLGk9cbDbLZ12ZjA/v9WFC+Z
r62QcyBx9qncjsMHVTYG1LdlL4N1d/baREmzyxH868kA49/lEESEMjmwlPJgQYysK5+UvsyI4lHR
5q7brojqozsW+TtQThHH5ItqB2ykW6LKr8NZgB1hvPfP5xG2C+NwTy96gVV3cLePfhe/axZXbHBG
fpuInRCg84Gti7ioTvSQw1MPUUdiWdY8LRsaRHoL6wcmG1DQwHOKtCVqxN5E4Kbr3b/mXm9bccoH
3DKWCcZn+gYxLG5riyHlildnmilRJ7eBXLgIG7RlGaamm2vrDQ87ZrQCoTCUrrHiPqNPI4O026Qk
HEEJYoOAo60IlUxXyZvtenwJnKEnvlI5MIsHGY75inIz9/4btlQne3Raaa4sPSOZdlCkQpgPoiJ+
BYkgyCct7Tgq6IxGKjTn1TvLKv20bHcNDuuZ44Qy7O/jeap9Gkl/UfibS+gQlA2kQivnROtQQXM2
6MqLXaDtURfWop0Vyp4OXdLeP+kkJGth4NeDbm8pp3sNgW207Avjytr7tZHvraIbYJuAIRLqNp4N
bWraC7hW+56MrDKvqsM3fKutJUb4siDsl9j7g59W0D4WiWoq8v2DnLPB+OQ0vSxUATmEwib/nLkr
Q/2V6TDvsJS9o7lfhVDR6S3sLwoxYeJ5PBZpmEtWTCFLhzUlw8ZZZrANV47NZ6hbpEYoT0m3tNOl
nsnyabKAd99I+wxhFp/EpWRViLqaEr1yHIl95iS67pfcuvI3uqCrXpwG9msaSqUpv8uDMmY3xo/2
3DEwqAHq44P0s/SP3fkqAb6ZeQgFOPc5Go/7mbjJEUzEWyk4EBKP5o580sAG/J26maPU93TSximj
uoGejLZkbvszTN/YY5HJCC1LTxu6t0/oo0Fny6SVyZ6nq7XDinggc/wjytXbC+bQZuUQiVVopgDh
Lyy5/xZt0FgCS6NcNnnIJpX7VP5wvAwXEcz+iuZuCklUcFgnJOftjkefI6lePiEo8yuU4nQY4y5s
omH+cHO2k7ZbZH+Ig5LabEAsZe7Tyxxd9BIaVZiTjSzep77YrkftcaHkQ9g7BbeXszQAoglCezQY
IPonEYzmeFA3nBV7fQ2qlLzgPw+va9u+YV5Fiv2ChibjQcL5m/G44n6LXuSqCP63nPnKDqydMk8d
lvSqDd/JA6Uw69wiLdXQin06Kq/ZPLhfK9tpNLnBz7ivuuhNOi21OBs+Voo2H36ddzAfrC1KPDGV
zYg8KqW85kVZToYy0D5Q7rGrYQ2RNR672NXXdpSQ6+wGFMGajyzProPBXUzL99DS73P8tlR3QLCM
zGcq2OAAxT4bo9OL+Wd1VHjsulZr+3COTrL3l55cdPlDhAc8jgEFwqfzV8b0WpHrFvInp0yOxAkH
7+FpPcfhspMBIetOaDw3WQ+ZTihTnlWZjF6FLYwdIZdD3rcN+wSz9lXE1jk5T0UjE8B247QDhiRG
PMPeAXzgW645kQUeqMXJiils6T0QDOLEjoJNrUVo3UXX3LNXb3g328G1gUfrWfjX2rzVvN095gh5
YewWcM7qmE8Kqh52HavnN8wFFO/7y7N/6gDqiPAnz6neoRBucDtBp6Zr+1T6OsSjzZ4SKDYcJ0xe
nzowcc+cpfYUkc9dc/n9C6Or+NJXVHgxuBTk/XPinr1dZtUjvIolTgLQ5pGY9DA1AoXTcJKAeE6f
F/+wcO2ivQHacayA0lBIXJexuYb1RB6jROgYsQcjDS7EWOIJU+6kL3iY2q4bHOgSWWFAkDgIp8we
H3j9POIlfTMHtVTb6P2909mwsEB8xwU9x/rtTKk8s26zt7TwKMYEwLKyKqcvQjLYEaceeMnSm09l
V2aTMjI60cwK0FOVOEO89fqUxfVSIK+X+hJ+OdtyXUT9bqnBllTJtkqsrnuXkvDfEOfn+MFvGpMj
k5o1ogGsCXcqEBUWS8eT7v1cAeZOdsWwy9Rqu8RbVhPo6FQW4vY085rOr9eT9NLQ4ZlnU36OVe3V
EBAXck8IqXL0Y2dkR6gnwzIwjmxDYNGGZQIZy7QHcA22hvxqu6/Ofm791k4bjxrpCNAVNSPhpckh
1EaLYDQBST2IhH5jJ9gINhM4rD+GCIofhWkYb3tM70VQ41vwquZXPdyX6AgamfGReo6joSCS8ce2
It3B5qaKzM9H63HQ5ilRPQbJdhbGPDVqCXLdwSVYYwvn9lIs4y5NDNrxNv4GmfFyn+kPNJNEx0SF
1+yhtKUHIXli7YZGn74ORrAMgnhdVQibp1Tyw5s/5n2dNCfq0CxbiDtEOAt8kVHLH4dBdlQr9FOs
ujhQVj/hymXtzQitbKfRpNemhCvMdUQcFBnbDt6qHTvhzZFDq+IPVMgbZEJmzDCQI9CDs9cnO2PG
5s4jqnkmIsGy+THK18dICJN5vISzw5Tcnjl/d/apge8yCIrHmi2aVDZuCjGdJl8qWaxS9TuGIMIy
crCKoAvhEbxWoqxkiYFjd4a8/oAo3A8aTUJ1wrzv21S/6ti1tbJKK76DSmSwBKVMvjUQeT7tUXp0
dqjOmrxhvxEPqZH32l8ry7BQU0BZnrScNM0ZcCJkOmvjHax+tt/erkNM8osaFfrGWqDw49N6keOs
SmmU4W2LnjoRLnsHeZW0IfYk8xDaHTCho6/7mgvedYtw0TjakDa4ST8Fy+s0RFCxFOxzUcti9A0J
5Zn/d/+7GwxryqRBo9KZ7V6YOSuH9DjGy08VK5NFX1Z/da+Q/kJSo8U6ADw87MNUMjUommM0vOKW
cooW7MJkues9pl69Q+dXuERguvV9v6BwPtZbEUr1dxkxM/CJc4KS5TrIQq3Z8/Xlzbae+hSzo7Bq
85JKccDxmHBhFpW1xM88zgxu8JfGsdUAEqT1TtnREBppw2SSMhsQwnDrH87CxqUwz5/WjXOJKPZ5
uwDVEQFSqfDXPVqlKJp6oBo++i2aveMVvK8DOqBpknVfqlpHJCcCPgW0QbdhPXpO88qW6dCRYD1P
bvwGmwIgWjTwLTiYuFT68qV+LRDFF3LJ99AdcVtpF+UrR61s1n75+L6MZvzoksaVZFOyJVj0vobL
KoE4iWNGr+jYKiVZMDieHSju6KyEJe/OcuykQVQarn9P97YN/0Nd7/6Q3QTJubaf6lFACyUtzLgJ
o0r6oBlKYUkjd2ETIFjDO9rwZHJ01EelMooAQbr8DdW4/S75UKeJWHjEnv60vC4a17PdWVkLxiCj
hlbW425ERWW5m7LtQS4CFgh5H1tLhnKoICBy0h9rNTZ5XPvYxnqVNK141azYc+dC9JHSgDtuceUV
0RmPaMzTKikHE+E099iagaaH2+Oi3j0uKy9jGp3I2h6+jMvl7mCjiA7wdyUxKJl6o+6sFtJ6yvxb
e3QhlrIwQdMRdEwHJSPeTcPr4UHGMnQ9/M9PxSmSdAw061mORvMNUALZWubMe9vUX1+q/4NooZ0F
pm1h236K6Re1hfVDof6cS3dZVGoOX013JI5f0hj0jV5GnQmmobewOkvt+a6AoTDkpPgNwXNw4jKy
yn1/KIgfWGlsNWMIklJ1Iouyjp35usEzAcJL88dpyQ7riy+8Vei0FlhhuJWtZqiZatijHd2ilyOZ
Z0rLvFiwHzZ5lqYrGvgLf8gD/MckRF8joca4yAaltdqP5+8Y27j4NbxiM9WbmGdHhHF2UnNAdNwL
t768KCkgWoSGULPycW4DlzPb27jmbgLQc0FLYMtpNqGa3DEt7nQ8bXhN3HxiFlYTkLxGov38ZVzx
nkVAkpVKC5eF0srTHns7mE2JqfG76BcDD1V5odwCuj2TwcqUhyn8u27yf7fB5iciEmi7kC4RCxL4
RvwVbEKYUJjihS/RoHiqyiWYsyFvphJ4KnXmGmrqIYeuBdsRslhWaMKOHpYw8FNm3JhMDaJ36sq5
wleaXQkzlH8Yp7jOMU47JOtCnX4qyV7pYwlQDyi1bIoffr6RzrIV19yCi3eDqgtkzEmxsVtWpBMw
IztGuA1vyegSRM+vdBhhozc+v7VL69+hoPDFRUEO78vBwZ9/3p3JBBoRG3d9VsIAu8HNooN3zYao
mZlAx41qcVZuz0EvTZZBpRPTd3A5/RlOEUkVRtIf9K6kI6GYIiRij7HlBk/N5uWGpQa2faekLI88
eWlPveoeenLp8CB8ewDMfWfTb9kFzK5ah+NTd0f816wylVO9nX02y65M8pOPQwSZVb6Vxw1fCyRw
krMCTgciGOPfqbW1LQ0re51OY1eBUjVlyVu4DbZ5ErhoQNGgLSdSYweXhzFX+7cXtt/J9DbtOvcA
SfgLlsUM0HTKtHVhwGBu0nkppanuSufJFSseTg5h3+78EpgZl2OUBqNGKPGUXMdLMK+VCtPi/tfM
zFAoyO8pk3r7CwUr+y5oBL6EquejHVyhqkRjT5O87IsyHv+ep7G0XsbZiUlMXldTaUOEm1IQceFv
qSUYCNOIo80K8O2XowbwlKh396gdwROp3MimW3/7ADg0fZf+1gf8z66LDIbT6HyTcuVkbHB7yfpG
JYqakY4zYhdPISW241uCXmrAUlmJOe5NeMAM74BN70iP3XLpjhUa8JmJkA3pwWmeVxRPBRSZmCdg
oHiPPIcI3Bm3Uuz8637Zr1Q6gDqFjtgEC/vcdN4pe9f9ZecgggsjRYXhoSt/F3ZKSvLlwPmPMfHz
D1wMCKbVpGF5Cj+ZigWN84es2f1+YTqZDo4GUvyYPTvYdS11wJK4ocoXGGg0hiYVE2D1m8OhxWHa
jIj/w7uOFApabHBkrpkWPgbjJqIXc38apA3dlAdinptD4nl0wFL/8HktH9vdQSfB8Oy6suAM+NG7
U9zcFQPbs4cAAfhoiSUjkoCYhp8I1EpcrV8rpcqFjIvlkZlFjbHtoIwojNYgHKiMM+7b5RHJOa69
urNgCABj7e8KBQXart0H2KGxwpjU4VmXLJ9voOILBsBnC4auTL9x7tnQ7iE63jrZB6HVUxHclqvP
pi+aQzxa6RdTK8BBR49W1f0TvN21jO4efaJxi5ctff+SWAs4bPZGehVvCvZFkxqGhm0kYkaVUp2j
0QfmdG/GS175XAUfhM8qVC7CyBltr4/xzbHaIp1/jmDe0BlQ/xlU0+UOAoaIeo22pwvtin04ICV3
d1ruo78sjP0W2O9W0eLr7YTraAW+dilC7yxQ/EN8NeNpPK5Mj7Kp2lGos9IWNaSdgg5DgNhDOazu
OmPlfFcjc03hhGMl2JhCSNTPixTdjk4ORrF/V6xa51g2Cmeb3ttPUlNNO/mHN0W8KKArlWMjzODK
fJ884WR8PmCEBWKO3cm/9SHeXUnqm7v89rNHBMRSRpSCBvtbFgeHL0oYwNMkop0XVeyhoHL1k3Xc
6OLGJ/uTcHdu8UJ9V2C/3OiUnjNy7DbvsAmdSvDGRt9fwyL1vXqSt3Gg5mV6b/6vSxNWvxd5OKvN
W4SB0Hol6NzaXpd9b28sMYijXCUUVAXd30vKCGhee6uX0FIRyVQXpDNGkNMBJ4Y2sbkrTyCbxXBL
mesZh51zNwxSDWvRNNxNPfYQ3XxKQenLI/m2js/4X2C/FAmccg34hw/0undatGSdjrLL+piJUvn4
KXUyj58WisfXaBpYfdCeLa2Ax5RvpoM8/LK04lBi8w0LLUSwCtGkqIa7H5bodQg1vjrtdlW4xHWQ
yRP0iqCP6LbA3+Ht8N7LUG2ORij1xvwk6oKrLN8SsaJxJp95+VsklStCM+pCmpTnkOjWhU6enaYo
cG8USYUP7PvN6ShVWfqWEDsIuyd6jsqSYbOQbnXgdqAueto0mCy4Wo/pwI28jLFizICvE/ku3pwK
x8NaF0G2P5V6M+AmXg3gZFIfH0RWnUoz8SRMsQSpB4c9nV0L2eVWvQsDGy46UENR2xoH8pfwftot
SIIZL9wmq0y9/v+fZgBREwy48JzZXVYCfiypTWTQ2ZmQSFZ2MILjYLbsOaqd2O8g1kXlPYEfvUMV
6qhX2jHj9uQKO2Bmbj0gdZ+JHD2yJfojkrdKR0MUy33swCvkNoTYk4T8CIHhITAjGxFeVyvqOeqR
4iSXjZLJkqEhyyu513EFY6dO2OjXkqKQHovaYFeHWqZIc6QgCLn0BUsGxoCxgZUTwBu2Eyw4voAU
0m+Qi3gctouvo92Evh5t507J4mKQITtO9ZRR1Wu/Mzn8wgl16pC8f0aIPGlXOVqg5hzQ+/6pQSGO
7Q1yf/bFCBvhAQ00hJC02V5XC9/JeUGV/oT9n1aDATcZWCQLCFZOU+mLpHsI2et3cdSXEWd9ALFF
ISd7QDrGQb5N1htcYSiIGCZ7+xDxqmFzxRwylgd7HVjUfLgN8b2Q/t5NR8rcYyOAmovUJYAJEUFX
EDVsNbKb9fNVgL8iPkQqX2bj1V20AI+uaFgpPck9S9BmMtytG7ADkEK347/uZzShPysEaDJD7eIU
YeqEcQxkPsz5kK+wLlFg5N1f8rJkZML8mJKOVQqgLcXvHAaD4IfidLsl+UFQRM634can5zaO11X2
poLfyoUPlApN9oG5ovtiqjanRNiLzbre01x1BYukjN6oPtLfptqc2zNEgDzjc82XZTEaZzNlkUfR
dAq+sFarceSzlBbXMMGLX2mmQippKWYKij5voy9ILYB9WtAumf0qKd1Y4U+xUZcxK7H/akuKYLbu
4IwPd/QVJYMNdcxlxoONbKEV+I+cxHrNunGx+GsQegn4N+GdPqWs7XDAprre0J7KvK+kIqRrnjoP
+uMihYi89/2TzmTMyuLql8MWpEz8E1eikIM1xhtMKPR8GD7k0icnNgsCygxya1f+XnkxXMwF8h/3
yu7uvfcw8lUmd5uGoOhUq6vpoNHJ/3frBQ88My5LW+aqQbqRaAtNsJwk5JWYFys16Wi1jI97CxNa
NeI9EZ3BHerl/1QFrzungR9W9ZsiJsFOMlAB4z25n26CU55M4ENcJfROxEwup1uUxvMjX3bCQ1ox
tUBEWonZayEfKXYxGW7fBvqZVrWpEy5BNWY5sHGfvt4r1EK5AXVa4a/017CwLg9dkT0ZLEh9kEmd
1sS8nb/m4RbDwexzBqO0li/5B3f0ChWkGhrDbs6igp35AHk1Bik17g0ReqHXPN16NkqEtYmX1qg0
zqUBq66Kt1BRm0wFQe+vVlV5IPuDHpPwxb7ymd+9WZMJxF8c1HTDOtYyMssgk5ICb3r5r0t60LVM
zy9y/ziZ0m5G4pCKwMkHnbwQ521hWkq6gz05+QK33M9dVmutyRUlb91efHB53ypcS08HqELAZWu9
E2APK5OLtnWSCVLC8BBQy85QCqHdJjYBIOBgipxxUhi39qgJ4aOVBrNu4VwRnSnTbO7uGYSKsR82
W+wwfex2tXwxKFp2ZjTqdrnX8bMkh+beIzdW1wOlAh+jkgPcBSbyc2jJ1KaXMPJXmb4PmeqLaRni
dwZvsE14kueEWDrzO9xBz/cQTw3oPYUx9H0Bx28Lqu7Ebt/WgcOcBlOmwEgYvP6NtMvuQllq4yLN
bvVhnFYzv5qyjkISzDowIYKsrL+MDAruGhVkVVR6mm3HLer9P5ptGPgZKieeOkhJuUEDEgawXQ5J
6hgJz7tMhrmfLjDnRejfYPIWxFlMPGI4/llcYS74YQdqMMzD9gmkE3RPWgznXzbxf38Xf7/BzR6t
v5vvVsV5tAE+3KSGOYWFdFDy7vLxUSKBptZpJzqqCPzzFf3VQFOu0/dyGEhVeeJa0QlBY0EAay1d
C0sn1ik4hsVIj6pKWba5qARdDnUGNZHd1SGnB/fIUx+vtAYYSCVqKooyFI6Qf74Oz0mXwaalSoQn
ipTWAqsFqHVtikoDBb28EDq5b1rtU5yLMCyuKgocn2mNuBMKUzW2Ykar5oyBMOc4wehn0PUUBjPx
xhN/w8nkT997WVtbfFQQm93MYYmhdxIUy7zKE/5uFNLmuWxSsTsQuDZIEuqUuHKJKufUUBjeV8vS
5sKRswC6KAvafuwF86SV49WhS9kfGb0jrvvgjAj0qNiGz2yprpAocvNL5n8oFvML0L1Kq1AawGxn
XMXgVUZPBqM5aZAjFhe1fozKrp8zaHZp1ZuCI7ZFjwrDPxGy2XDCUfpqvZG7JJH3wRIYz4vz2MfT
Gc82YmhO/nvEqNhE1R3zDBRxeJvnNEP84sMeS1aHoF9D9ImOQcmZL6dX3jrQuYH+40q5AGGQ4Mkq
Q/X+dMI6y0hU8W7+VfFaYXZX5g+UL2+nuDRLX/K6YULsXshT5ymW7YQ6LxcnZvLIqSZG+KMZsfzn
PrVWYhACoQJARoWd3805FpHHyrxHLf2N1CFxnguAb/m28WpXZ6oXga+vcALk130Yr0DAYqQwmI6o
k1AFrjPoSZTmTWOxNHJYNGMiK//0CSUZjjvwHgu2iG1xOFKZyHWfJnOm3pfYtpNHkVysfW9v8G/m
GWRY/+aNkZ47rp5sLVb/z0AYOPMekxpGOZ5sTw5/xEC9MbP2QatBA0bVySGcP5ZRLgSq90YxDm7P
hPTYkQG28Y1JAohUDVCZ5GLZpEygSIDGgSdynsFbmfBZSY7/tzsNtOM+xc5uWjaPZQRrGkMHdR+p
jydJ2ZDHozB+XBdSGQ/YH1E4O4CdXFFdCgthMH2pmu546EoJdfjj1S6XGWStJeRznGpSIc53Sic0
xhFDWqIcz+DeFvVro2Fakrnilu4YGBP9QJdy58Rrl39pRQskgLOPz27DzdKcZwEu/8j3RfCaSaGa
X2h5byACXdQJzI7qh0Oj8FR0u/XHwDN3U7WlrhSGkg1VqxLJ5RmSATdktUylsxI6uMMlUBQelO6s
GFTLlJ3HpNLuEG12SnBBmZL5obv4D2nqDg4YGJc4sOoSCKYb1cc2plBDBvHd6hSvp1R/acJoiEEq
/VZrgUMR19eREAmfNi146q4PbL9CdtOEU+CKv+cjJHsMiwDZjVcCU1xuEuZ10BrZFsiDEf56b53u
nit01q9yrjl5AgjUIAqaRfbi8TQqt53SnnmJK4YfkjivHvsKHNYii5d9a3ufUnPDovyMP3ftUfHT
H2KtQgdYwUu13r1Q7Kv0Mtst9VRbSYQ4TpwBTwU35hA9b+ORo3cqY1T25FG7fR/OwKn8A5abZhy3
9GXFFLg63ehottyGD7N7OHGW6iwsgB19jmHwNN4ut/fHZKSE67g/whPZ97vq1QGSyxjf574LhiPr
giygwqXiBHFpyOZuzFFq12124HaXHpo+ZdAIQsI6D8bfyRDztwWwt1ZSK/oBqAntwp50V5uwdRNo
/K7tozFQvMwVTWuF1CeATr6rLuDe+SFTNd35PQNvW7cbDzFSEb5oWp6wklW9rDbALx/tPngfQlqs
5hKZ0hn3Wnntb2ZgLgzIraXKW64xwkS7kUYXYpzn3zhYQhNQyEktmiE88ka0Zc/AxufCMAmtAE+5
CkqzN3TdF0ONedZULlyLkpio4lnBppbAvCAB3i7UfWb069PjLoNY4g1e0iSXkNSAizsJ7LbtDufG
vTQyee5GULkz1Ok3T1y1qWdUb+SxCOZ0o0UFVbtMczhaTTRy/uAgdNuuLiVc+zxlPZT5U/075bPv
zRfIym/oLU7sSuOsqaNSLHMtFtgolHmHhcDjyBU2xpqk1Am0Rsc6T1puPmLsSA5oGPguGOkMDu0p
uCA1qmmliOUXdwGVC160/OwziHAew4nsnw34VY9vx4kfbOePoJlDWtsXOMy7D0vqU2iePwZ58PNh
QjtLv/vz/WHG5Ks0qkhiDI6rd1IlbqKoLDqrz7q4uqwUpNwneo9+upCK+Xzsf2CVs/SvhKe4fcSj
ozC+G97T9gP28ZfQH/87zOVyyJSdwjgreKY1XiXFP8z/hsLL62FDEpABcrXX7QXZtgC802/By4Lw
IZeftKSSRzSCdHuIe368S1IFW9IcTBZx6h/L+YY1JNbWMaJHLIN/MgYcHM4RxjjCrzimIY1vrbsc
V1j4Lmc6YL8H+7/QUAnz0r9B5IvErGDRIaRHPUkwoVW+Zjq3dmWbN5se2ghvjNtj/BkTVNioHWrR
7yp5M5j++44mTkgtZVNuMqR+zPqKne1XX07E4lqfKBoq4KF9beuXY5f4krao/lUilrcsUZiiNvHk
e1/cBh1RGwBZwfuTu7c/WvbLFHiSltdj4Sl003OK7RAKXVqLsRwAtcEZHOmneHAmTriVLupb1XkB
nmqqIYF0XjATDJklFWbLhvlxI31JPO7nhGtfe800Sca86OOcVAGOt19sTmiLxs1bfnoqG1+qqL3u
d0cgRXyGu10QV76BMegFgKAywYKfuYPI6qpXU7/nkBzFYpfUUAoQOmpODbjQoEI5/Vy+nCVL0wmy
IiS4eoITGpmkpgSAJHOC0eCuzPUSmow2uqtn7tYQoRN4QQcbKdunIBxOiVBpZyEtCk4csDDgDG8r
rDoULXKADPoCbmlLn7ks7NU3CIPyxSOByPmGUFuasrZKfDyRDRIcHGPR3jncUjFiTeFsA77nPcXu
XykIIWUdWiJK944wfMGYBWN+km96qk86+qdocaI8Vdiuiz1oWhzVmv47Ps1mDNRvJh2MjiXmAo0L
YPTDSC5dJNsafxLSmAwQu4bJlYX0vrp/dd5+ImEVTRjORnbmhdZyD/WhSxoYKenECtFVJuPyw++h
KD3TYZ7yCiDglMAmGo6G+fXEZ3dIxWw6fjs/5p/3qDlJ5qpDxn9tkzOBQzsJsBgs2muWdUsKaBWL
s4awAPLNDar+fokm6ZNS8hm0DLtKUI8qpYlHiEfy7ck4Fi6NIg9v5Uuy2T8Ypnj8Nl2i9FmYX9bY
KbbrSGACKSxYRJ2pzmH3Vd3GLlQbdszlSNpshoNSo8wBpjhLZ2ignccOB8mulo2u9gEQQWOSyYmJ
6hMqqZS+SyR4fv+/Qh686PmWnpmxSUMZtGR/d0tEd88C9YGkQvrd2MvKbV87/yAF3SfVX6CVBnFi
IyN1TANmNxfEzzTreRjbgqAyuPlqv4fGKRR0H+PilxKrKgrKgM+1Zn2pFjMdSh+6qEfqiw9xMiub
+sWwAGWnlFfNLupjuOE1bHQaC0IYkdMfHwo0zB2oajP8y3Gx6RzXLJvBm6boKLn7UFzh3HP3NbmY
6dgmP6q7oD0DtWTaAqFgm3Dtf/v8tewkzaMaL1g56fwPvLoyUWyO9Xck1bXZiHTXxp2y9yTR0XfX
U6ohf0LhSNISdAeTMHLZDKe9AnKyORoIL8hXrpkmjzOWc5T+tj5ugMgDeRITH4TzIdTIKI0lIy3s
DSORgrNyCZwZRpTVT3pQ5Zu1++NXSLysXIz7Od/jFR4y33lqFYDOVB4rwDi+0I+JJsGQDmlKm76w
rWVMuGtbZDAmYQF5212Kcl91unEc5jtBBvE/imdRBpm1WA96BNFpaRE6d7DlXQ1xOHvDEqchnCFB
riiadtmZXioE4fMKUP1vGlwL4JEdxBbeHiL92QxtaG0cBOoFe1lO/AR9lKSNzUqLE4bpU1H/uePO
5XGyNfjSMcb04HxKsBK54Z0ooqaN7oL9zOBFBg+5akoPFMHllnM9dFgDI9Zb5KdFfKkmOl8F/Dro
3K198iuKwAAaJYWAyjbRyqM/sJie/fxg1UIRRJktoVsBQfPN7CcEAHflRkYmi6HnUx/NsNvDaEie
kvtTLr32lhPsja7ofJJxckgCKl4Bjv+uqKfjcuMlrty3UNDSnNNgEZ2RD9ZWOYix/Yr5PN36d9UP
NCWGdzaWzmiyghAGGvrcDbzseJ216n8JrsWcMk/EGxBKIZmzxxwepaPFaRjbPg5QFZkHzOuM9cj3
1ElSaP8dnBEnvNKq0ZC3/FlQCq5MciHjLPoQ8WC86mFrjn0S5B0Lrqhz8X3qhD8qLqMWLbXENatO
84xumP7/aLr2a4Qabn0F8Cn69mX7q4WOcUUsHUShfWWODlFXbzZOEJ5GTUvYRFeEhs0tZSnzCMcx
qE/ri2qEvbERzZ31WmXztM98YI+snC7qJjBELnaJUsQvEMGw45lVvV6mshXaT99SW513FE3QEK/S
2AVZndmZu23yUAzIsUrtcW+IiXgcszKxlILnXJ1IUFzScfkdeShVzO5GT00I3bo0UVcf2E0Rcoqe
HoDIXFBazN757gIdYEy/43USWci4FtkS69DY7Pl4ThGen2QankRFtLNSCnDwMnxD+VWB8oStGxGS
0xazhYU4Zq9WACH6CTFXAF2jGO7CcH9dhlSczeY4DFeHZHUt1yOgBGtrXeOShY/bmre40pWkl8Hy
RhaHZVj/n/pDkWl7mcJUyqlkI4387PbRfZO/+RNvSr+koWMvgWe8y2HL7+FrAsUNN3wJg0CJXUU3
Cb8qhQm6ay7X8VORvWBh5MWVUkxc8ah3ItWgS+ehQnAEEHeFicUufsQL02RAo9I95OgK5efWzX9T
aHs2pJUweUaMTquCnp56FLDkdZtZPej9pnaehkX/rmd1uOu01+opVVUX7OQm//zfXQOTGAEwxhNG
zK2s+W2Hwl0bUQRloL74VN8WeX5BAzFyg9fH1nF3AjXiUqAha+YU2j6g/m+xx9iFehS+U22tSgyP
ocddTggmWMVVQoaepOQXmq1q8A33olgEeDcLF8eF/fiW+tzPvnTT7L3tD9gjtc+OpQkZ+3nOuv7r
aKEzWJYSAuMhVSayKvjkPxJ1Ar+0DnWqjgV7SYTlDK/5vytRObd0MOrpAgNon79akEWGA7xYwscS
GPm5Eh9yPo0544bOkL1X8Sw80OA1jYyhAkAYVyjtU4kg8TGG3Aa8zTiQ+AThNduMDE2CdRC/2rd5
O6VdooBoLz8CE3L/RqTQnujm8leDLQmnBGRNrs8RU2M2r3sdM4/VMVEi4L4LWUrmYjc8FH2t3Aoy
+Xmd4iLxQXukUdl7EGS7nG0GGwlpq96ZUW2d9G6qVa/Rxpu4fYfCOVa0FcY6Ww0MzWsbMa6bllOQ
s3PeL80CsejmohdHEfUDBCS2E5GjzNLM1dTCTzv/b+2K9xLZD6rdLhiB18cTi6YIHey3a4ofHd3I
2DCHGXe2RT1xwcS4QVEfbOJirGRiS/B/6w5AyyNV+T+8ceaySQR4kjqibKvff6USfU5CmNhNDzx3
jvL6sRkpQTAYBaPZbLQbMJ8vZtcM4TF5Y+t1emxtEPoDfVMd17XY76UJlRZafzwXVoaJam2f0Zyn
VuYPg/ZOMJDDnFuOXdMMKfi0Sdmk+JIB+xiEE+nuZE4UVNYnVJ+tn0FhDD0wvTsazXIHt5qXmchz
cTSy0ozicnBD7I+fW8iMjttVEQxzNt9upqzgJi6bxzoFVe0biYkTUEPVEnYHpSythNyAvCT8ohl9
zN5VWTwxfTsjCgYhC3NSP52+/hw7UfJkwWsStdS/vKQOoz16FDIvW5nbOrZRzO2hEZw0Mq4co6V1
bJ7oCm3y4rl713xkhQOcWlX+g4rzPAifumKVktjFguSEv55m2CoLNaWasdvCTjJiBCDZ4KZIZj+r
usA4eriX+t450pp+kkBZxdmASEiYCkxJEDlEci2EmuZtYdv/l05C8KIERUYXP3Z3uhEDWRCznwfX
ap4pVF1yM0jGuaZE1QWb/W9so6ECyAGBWIOkI4/judF/SGfxV8Qm1Vp3EPsOLXtNEU2jpLvXomfa
F+7eNEXP8ILd/2fCXXxN7wdqQXaG5ZzP4Ic5eRDzXrYaygqLFkHi87RdhPLYLHPAe+Fc9S7rIpcJ
WutVJmYI8dM/FGaS6erG+xMpRheZnDCXo3rPeErq8R/cyD8HBRYKCe7wfOzJqqPCvYmR65mneyte
gXryWlZjQT2pxFPWUoYh5rJ1w0jYno0SfeH5v5zSzRzDrLvdLa/LM84ntzEp/a5DkJcCUijM3Tru
lvPgpEMT0awWoD+XwGuyf/rV3+PayFVFIW51WMG+KTSs8khwqD8vOsvzoTCy6xVnxFhJ3XJO2xUb
vfa/cOmx+4gmY+9tEVHUpPiB9krPwaW7IoGZVWxgBo8p9F2cQ6AJwz05DXIl9t7y6w7Hj51L6EVL
CGe/YxRaYUBVfsjsm2GoAN5kC2fhZIDQTFxFDyryEuXJEwemMcaWppXdkzt4cDuTDAaJm2QE/7eI
NJAnPbDve3PMYhmldAZMV3J16bmlRXk9aeZvgOPIxBFTKWVe+N/LqXwDGT4BpLDmGcmUOTAme3ZK
H/B5W1DV/ljs8mQ7JZHFsuGjNhmd3WFkSu9RiOIvsJVJoJ8S3H7tUsqBDo6lCR9cKaYNwkmA3A/8
JHcs7zGQ/wD3HTDrKXE4ibtJ4hxSXFfXRGOUUYClaotAPoVNaymYz2q8ytxGfdPymdGVqOoIYNZq
OABklLdQBvt1VwO+y6qugj3UX0F2BqTcKWKBnSfD0Q4ateK907FIpST1TCbwu93rXi1/ymQnLg+t
CoCQ6YudfPO1B+YjZGoi+itd5He51k1jkT93hhHlkhZB5atyJl5U6/VQIScU2T2Mj8iNPOLTR9tE
iaHFMhjQYD0wg2IaAiCyGDhN7zM1iz7uLh3HmoJz/FDhgchvvDh9N0qn+Lp2U/+sVx+22G3cq47r
UC/Cf2kXirnMRXDerv9uEQgziKqE/Va1cj9hLJ9TMGehQSTXkdzcbvnP713PO7x5DbEXmSVYVv2K
5mOGpDyZon9si924maTDKBCY33tsbjnBAeok9GIQY00I8bxq01w8t2anuU2mOp6nHGEs35bp/fTc
6hhG3BxbZixp4ZV40ySTG5uUDhQ5VbRQ7K0ySt3s60ACdmyATRqTQMGYiOmp6hGPFizlWdY+Djwk
VTqfaW1gEQJ0fy8lFKBAnlhi0SN4b2RqSAVZfXagwmDtckXcLieQZnaORkjF+5av7vcNZ8qOe6Cx
LFwQ4+tBFf8cG9HNd75ZLNgaVqw018w702gxw/GSr4wwVUZ6lR0wgQBcLBZdGVt2wAy5FL6iFln1
QPst1nzIT46LbpSmA5cnLURoXH9wf/zRf8oH6yd27fPnXz5L6M9AFJTRYy+Zgi+awMYocFvDM+RS
JyjZPZPgduxsWOQocOw7TmxE565FF0gQ7FR0lW1A6IgC75vYzHGMLBUqJFNDs2ix05DON8N7pvDn
6dl+ww8xPqQNcsWGVTPBlgzLxGYpl5vw2h/Z95HO1Ob2ymKSbSpnb0Rn2IGXTVedp2ciWJ+Fj1Z6
ufmefojGBrBaTmBzGHZIS2kmD9X5Bmr7NZHcdiPaTDQCCDF4wGwDc8SGaX1PKV2qTMRXO2Xvq38D
YVdxbRfc5ZLsgrd34VOVXdd5INOoM6NYUeY+IwbaDkP3zzCOHFMvAEEdnsN+3vmEl+TaFZKOtOUa
2eoB7G+K8z4gagpL233em80J4+Db36y+28ewDXNcmMMOjnzJE62JSeLN49o6wyqpGG9IO7u8OPIF
NjEQOK/PjqmGYl8i9bnlnGFfCve9Ewek4nwAbfPd96fxhjnDKLZoJ9Kf0y2ETVzAujEK1UZAHuI4
5ggqmoJcbe5clAxjidAlJtnpWpNo7gR8ls7HpndovlSe/eJrAUD5Io/DVhzPOSbAwtFWCcqLkMZa
zz/hhenU4B/LmrmyJcP9gvtHxeReRIj20pvY/N/NEaX7tfnP4LQtW6gmtRflFw+wBhWmhMm1fk2Z
KxbEKAAd7vRVpHSgb00mpXetdLjtlE6spafBRkSPMAo0TkfVCiqbDPWiGvOLt3nZz7NYeci4J1HF
yg2u5s9Ar0ywabt/P9m40aAAqTLPkjbYORc5dH7g8WSwxQHbNPj2reZY8uOQiEW1MGtMFAjdDQ28
WVnrKmnQGjxkN3F+j+x20ugS4+L72HNxceMDre77IvPPXIAVjn5+C8Xn1BSoLC0U/fqR0fMKfMl+
ACHWyKAnR1RLggWlf7HKccBs7TfrrSe6luilo/LgjISO8S1PZrDNZH+/o49xaxjLZcnaeE3K83MV
v75o3SMc3O2Jar7ZFJoK35m7ji1OUVjQLA+Mj+hj9xq6V4u9WjqXwbv/dmm4zprjfnnrsVYuXZ8q
Hsl9SAJDXVcdGvxKe38KfiTGj9KvkUM9oTeEVuBbsMfUvDv83KarsS3mnaxk5npGoBilfPLx71NY
N5nNZQDb5Lg/Z7AAWCuvLq8OYxfMdOoEVOTuvM1FAA0ZPE/mPl4mugfeKZSdCrKQ3yexJkIeIrJb
08kHDnLcw3MO8Ozm5pdZnvO13IV3sJFhQky8lC6xJSmve96oasnWj+fmG/ZG71bdZ3oY4fDkZ+bB
wxckBsHG3VR+yRZ/bWJL6/siuRC7x093FYDYKpMd7v9vOp6ZvDVgjIaqWCnfqxS/QlH5zt6E4L94
56YN1p063Vhued2eqHqcsTd9DND9CWin+J+WtnAMT0T+Jh/XX7CXMQLLITEJ3JWFP1bW4NEwNkNc
BjiuG6gR3Kr4tOZ/E7uD3qXAFg5E37ZSzmdz/l3L+80VVvpXEJfz/YdxYn2kBUSCwTDwrvCggyfs
1qgvP5ImDMyL82OYz9SzvfBxtvJWQIy69TP+NeGgnID78FlQ7ayFTK5hj0cdkOqEbbOtRvDVm+Gt
GQPCos/PKNCNY+4Ld3FeganCuNoAppiwseZ3uOHOO17LeQSd2wxh5wBBk0A2209t9FhRShj1yR29
F+PJWW6LQi8YOliehgsmuYajzrwMXzjMn+UL5x0ic9a7sni3rTu1MzrcACUv2eCiT4TkyBtfp8eu
DReVFqWU33yzpncoL0ZukDnc8rI0uFak9ZULCALZqy9bqhIeB0u3kggD6FfwkVXElTc6VxYFrBZ6
2wCCrxbcvC09z2RF+JQ3r4pUzZOaqZ+cxFxLdLcGpKiucKalVFsrmPvMiyJVGujyw+ylMvDuuMId
+LJrUMA3UEfgX6SXKgN4EeZKaRR65JeTbefxmTfJgRHx6l122xctrUdFVU3S9gfpoMjjmZ91aVfi
EV61wS0sDvQm1eT+9imleS0y45HuukEooGTyifRSo2oFrqC9CChQ2GlW5kHFufRAes7Y5N5IoNFW
GWpcl/eXklP/Nn0Kvtx3wSqdEebup7MbihvhwePulMG9/z0OdNcnRcfTJZp1X/+53bchYPz5zWCy
7lnp7FHs0w5u7yGDAOrPkHnDdS9DjDAZ2qR+6/KUs3vkuWeZFGXhcRDLGOnXWN54SN4YVNmJZfj8
er2SvTvIZJjoiZToAry7ZuIpMFf9tvoR62yXDzyWigTkckLkHwiOh2kLf774RY5WNJjvSZExbWos
EY51JkNmgR2UJynRdsAtDsyK/O02qaC9ZRfNWHYJIc4xvzLoGGiebMW3npeRjIMNTeMMQCLPh21u
At04ByFO27pEn9TQVOtZp+X9bGS49TbSSrunyLuhmSkPTYAkvzhPo2+7NoprVBUvZTHzfu5iAyND
opq1Lo95kck1oCeaQKk/SQxVcUycYniL9fQ+h9d/nkDg4hgbYUBzt9Z3RajCkiyPS98zrAa2c5gr
K1yPHmW+SEUsT+b+WfrSBmX8yxXgud9fYDmXPPxLEvMTJhS6lzIgrkg8QsLUu1fI/rsWGVVEPaQe
AAQfLk/9me1aOXcq33zYb1OgazefwQHJg3Qxx0WfE2sFNtaAa3v6gVSvAUSQ2b+WmXK0Bq+sIMuj
FC2N0pHE1EIhpU8Myx5lIXSV0BhG9iEakHaRPZR1HAe56sP8/t6apmFVWBXMdFhbJr+19BD8au5Q
63PA+yxsZeMBD+dxkK4nDiFM9+7jTcCLOurYg1l13e08hUAlE7qdup3SkJzamjiklYYQVAG7pWef
3bTuAC3bw+B1gFeAsK2/Pf7r5v/LnU2DpAGJm23oBxi7QqVa8p2NqXO8Lsfw4SGZyqE9xs31uu+L
ehrhTPg6pWqJiG2MnMnwOGHhgVV2fT8wXk16bYUoUM8UPmOJhdDaq6TxiigLCLQ/6n6+yT1W145U
Y5rrsWe/k323PAAZvJKrtF4H7qveBByErWUoqGC82SpvXXgjuJrY3Fdvy/iNnVUOSL05tI3d+uHQ
ysEYLQAJyRJ/Kmwp60vXuC6eYt6EI8QCqRuXcaahtxOXJGTnB2hJLFm7q7f92m1jdXLF9KLRitGC
xyZeetJbxH2/U3rC5ZBLTKTPVM3G2vj4puIEdCSU7VI4MDqWKcQsI2kLVIc0kqE3H9XirISJgVzi
Liyg/YY5t293UfoxMgW4SQ7+yq3cz+oG0kJ5unthHGVmWH1cLoIgkFwxrnXCOwGLd6uyNm/NQ4e/
tTwDK3SAl4BXG6WX9zYmTc+AWr5bUH+Rvz0VN0xWXsEwGQ6LyOesdzu8rZyyYXg935IPt//2g5Wu
A7pLeH0tg5PcZxtzsla0jtvmTyiehpN2s3msc4uUaA+NcjJci9neo3eqVdXp0joLn6C51OZn7j9V
s7E9TAjatDL56Cej4bz5chQJbeegAW2v2040HXj0A/Dlad5UKaooHIfvNbTKCMXvS18DnMEQx+EQ
LSYpIzX3/EUL2NHcUUIe/1kUl7W6zFzR+EihfiJVa9W20kQT+xgIlO0tXcagG663fX/Ru3pfih0B
FWX7qu1LgMZKY8TEP0kZHGi3glfofC55u0V9N4Tz5C41BY9D3kynOC/8q+37/B43Y1/aUXM4Lcsi
T8PYuo4sIUBwO3Fgi43sc80pyLv3hIOeICLu7Cfw+ZXeVSNtEXUveFXTLByQfB8laNVp7DWNAWpx
qnd3V52im/CVZZHMXytHK7YOFAlCxjxmi93w38YQlqL2Fy/ctn/rMe51fbseVX8cYw4D5HVNdTYH
FAIB//OjOsfgFFt3pRTz9c8Moz6nm4SrUe8UH4FmUGN36oXdYWgbRdIc2OIMPpdZzLfemKV9jJRi
HaG/N+i7XG48sShYKp7zD+bu2Vw/S+CFcT/fOmCA7ioqPlv3FPSg/Xkg66QT8YT6znA6FuDDrSpv
UUqVblE3l/rTsmCtpzTQ07mBtpngDO1eg9ZOiynDc99fvghBBEK4mtlDGMMvApNlqzqv6MONPRBe
XVA6c8bPX+feKnMxUTYIQz7WlSrLeq0Z/1UOuidlylKKmrVhJIwebGJHHI1W4xUJCoTpD1y1qWWc
NplAOHWzu4WquMbPv6toFILv58iWAtrhe6On8FX0CbBAsPauLO7tmRiqt3NByym3n9E1jHMOUeZp
rEpVf1CsMBaBiPnqZve+5wfhpjnSN+dyKHc57d42Na5417WPDF2lk4wo+YotQ9AAJPCeQ4L9wVH9
y1RelMqL5XHiF2OpuvGux+juQpwXHWzFyEx3LhLYZfUdCfqAOQA+Lej9XXPcDYsnVONtdyt4QBWm
TW0jGu6QclrEE82Vd9U8DWFM9j5qTEZaX/GG1E3lNDUFMf9rbjqYDvQ0OMwmJimvJmOGm3OxTNTd
B2j8gOLeDVKmyMdz9auKdod0f+hrykmn2SG3RIVB39LtKKtOjF9JlukMme8f2RW3RRVKW/af0aNs
Rdo528eS0uickd4HCOiJ0mebusLqzHK2lNpd+uWlY01x0j0MVkt290Cy81hx429hcHSJRXjh2e8o
SDJsiSfN3j18wOhcqa7nrUVeIe2SFRzovA+l6T7OKbyeNpoO0yJtloP12pYT4Hu4BEjia9EXh+3v
gv8l3NGw7zxI4I3NcPXnI9o2vl2Mz2elEfFizHde30rdyKNKD9GBkm/xpoeBdWNA9+ZNBNWPBF2u
V7oyUDyZrKbA5q/BqKbCEmdGhO0T8y+w+Gtfxc1SDnGhpSqGHOB7ibhLJ/zz1TPAyucjmwT6GqCi
/lhDluRDa2PZohlr7dx33kEg9EAZXyBIQ8iF3+gAkuBek6hRkQoiG3l4Asak4LhZzgPVXkxeK/JJ
7LteqQTRd+F+p4MqSOFuuWtm30rxuaqJHtQ6evt0cgLNy89Pgd29r8l6EiUvfDZ2SZlQ+McBQKsF
5RL9xmdKxXPvuJIkxE67V77oMxi9+oI0vBup+vuiLAmOO822vll9hn6km1xVpFB17ta9gSGApAri
Zw+fr8BcevtVVzxHo6DZmeIwe2y/R4Ly02G653x40p/CixSt+iu6oIrPLM1hl0Yo2IClIg5h0by0
xSAV/0FXlb1YmIinCbj2V8wxldUnXPZUfMnzSVXr2R0kLCUQShMRvfPrp7ecqF62M+I7CjC5VT5N
Ubt1/WEOTfHrZ+j1aFiBE4kPRerqoFSZ9DZC08fJQg4da396FIqGjW6/Y6zmIAIy0/c/AQVLd1kf
H3OB8GaMq3s0eSUgdAqn8xsiuO6rNIkWRuv+NPa2FlCXqjP0f56cOUKCT6lVLkLW+5rXsuGTT0c7
HNFT2e2LzeihxT0CaAqYrk9S+EdDOop5Rc2FvddMMO4y6Ijp7n+OrAIya2pCr2iXXmHD6qJ0dV7j
xyKr3kKb/C7NivelUdDaGwLnzTs07KvNV31JfBUmpkVCOueLmejviKxWttfIZ79NkaEn3eaXUopg
dqA0jD2oEkNasrPSGIzHzFufVA24UYBP1Xzk+/WD/buUpGu8gKTftXlyJ7y5XaUob3ueHZdEdjgj
RvHME8N5ZjDGGRu3FW14fOIyUH0aUxBKXJnnieC7Flbv+biKr7jUmsbetMdt+b0hjzPdDz4qBMYT
svrWPkb07mV2CvCYcIxKhd9fKuuFo1P+QpsZ/QoYigJBRwJN7iuPLcy6Uj3Yz2+Hg6VPC/rxInXH
p5uryS7lD2CLsiQs6CuyV3U3kRh4/7xmJpOPU/36YOorOwrkd+g/+cBph1d90jmxEpchx4PtcuBy
rJrT0W+2swgFD7n+bRo+lTkKh0uNx/ZfKWRCe5IJl2H7Tlp4xg7+RNZbgkgYcI68tbpm7sLv6pJm
mZQGUbCRSqFHDVaWQO30mcc3vosZseWSfzgenqhSQwIh7O/gZd7Rf2sig3so1EmxsqQS9R8nFKZf
VIF9QMLexsoZUtii9ANpBFsfkJTIW7/eId5mjyP5irO3jEW+0PO1qp7eigwWRxdeMoD2cJes5b97
iBWXu1WaebrXQhkTIMU1VVjdb6veyOmujiPkoSwfJfssa3wbb3CdnrDtEZzXzFW1XHTmsxV0YmFY
Zig7XXRchOrzXZiggALCdyMNdj1mtp6Ks1iQ5Wrx7zlqDBIn3Tp3zDfj4yVpV+XGoRIV8DGSvUTs
J9S/4bx0LASnZtV0bSrlaQyGFEnH4IlIrrzqG0fF4/A5PMDNPSKYd08EA9UPlLwFsJ6qloZP/8de
9RBXF3lQcKs3AROkX+3OluB7m9qufvW7ZMo21ScHKCudIlYU79lSV5q5cVIjSLUj8wO5YNa6gaQN
THlPyOH7f0e4Fq+aQUPEn6J11Kx5FznuVZRPIvIg21EPfqq12mAzJgUa1aOHTTvVJ9rpr3sHqN1O
UQXm/PFAdldkN0dlTkCnpNyuUoGAuYtPWSapP4Jxv16I+eu5VFQjfQidHXiO46sgZEuxuWi9BMN0
ji26ioyoF3+VxipStDxSxEaR58oilIAO7/5oYKPP26TMI3phI1hq9jc0ikLjli94qzmlyuaMcRXD
rzqF89S/3jwDoKX6q+SyK0vRlymEtgxfXySU2Bd484+zN+Jci+LGXM8dPzoxAkGeVCSaEnJSGKY7
Ud4NcQU3yw8JXwcDqf9Tsptt5N6P/OIqy9rEX0MzqYMJoVMLsFL+8uZWdzgmuYawZ5YUfbs0IbAY
qEmypE8xTnoeFdm3ha6U8baTUS6JL+gPSi6QbnxTeZNjmkfd4wz7vBDa8jP2ps+dZ0kVmsFsNdGm
rnIOjGteAKJ7r997lsPi+KGwVtfTOUGB/Bg6pNGkB6vkyJ9IzAVWYg59h709rp5n4HvOICUkMfwg
AtpkV8ZczWdI8lIl2XTDO0JRTxyWPYmeLwnyDrGjGdHLz3tD4z2sUFcaxQ+AYRh70QekwRdO5E6o
vdBEp2vPFJndnF9rYEMnRgNtHmn2AcOx+EJW4tI2F3v2+p6hQ1iVzrmfn0KlaiZOFIXoN/CPNS+L
bd9OPcoGEyqzM37K702e3LD1o2UCayPpdNGlI5aTA4YKvOPcr3NpZvQecFAER6xaP9OQsSQe629g
JhriLAMKsaIAfWXPrC280jza/6lAE9SU5ycGF2RzfNLOZe+7fMbbCRlzYppnfqoE/kjKjLgC3baY
UvwLfDrOkvwarxmQzH413NYD5KReAH47XwIK2Wkdtl39j5wxizboZ1qnYGrmJ7UmCu+aEhGl39Mo
EkR6sBgNScRJUYhzQ2EIPlkJG7aE7reNec03m1On/n/Iq7Dan1iWaQ/p9bF9hf80+wAqv5Mx2/73
82qzIjNltnbYez28qmpQ6SxQYwSxqjsGAlO2huDxEh3pRhqHumQ4wlhAd7NhtZ4zp1yizXjVbDSo
R8cWj31OuAVz4tHnh/hLD8C7LmY/MOHnmwza+9+RLR6YJUbpd+XMq5mGtUUMYW2JrvLp6RfHyqjv
X5LkWAsiXVDGOUbkAB6fXNoTMF2EItG5JmswpeaShMjn3LucbF0oRsXS6VcANYUS8yA3jrbkWqIn
vjDPWXkReNNkdZlZ87GPPtD7cyL++6hXHEWwLPG1NrO0YL+BvQiSbe+mbpUTZQoUp3skUv9CuiFM
Le5jOdEse6dAVxqhDPd9HMRTnTrV65+djF5N8Is0k4i2OKpqZ+lclOqQ5YI2wUQvB/3ddJWE9H/E
IZqLvHX82V/9mf8xR1BmjOmiXvN3olRV+pLdg5iCAVXtxKNWXR652yJM3IgyYdDFEZ7lI+h+rjVV
YQvOXME/jiH+4iDHe/74zjV78sLlkotxBpDY3NztILxHrUckYzPQCC7cufF45rGuThl4NyWfm62y
anvWCj/a7UOdXAjN/QcJ5q/gptVh5VWAPe8AldHEZqOGOVhP+oVEmk+UvK+DWqCx3HNNnT4X9fBJ
wzsKZ1J5yLvEqqYjAot7iZvGrpAy3p1gtJBPeFybxF8dT7wNh9w0ZGczjbLSF9b06IQKhaULHI1L
qUCzQ0JPGt+DCuT1heEk1G4qFNM3ZwuH/BcQIcbanSpiLVoxw7nDUoxKpM8hTYDI9b+OxA4EAoGj
WB1N4i/SC5A6np+9icsQvhE9GDJeyuohwgtlSIdo4bmx0959K/kJZdvrJYuRpKsom6P3DBnKS8xu
lIFFuuuchqW3gDlzbNsUV5Wr7fGpEmHk6PX6VnyY5Tq0v8uuCCKoOxGq1JEADbejyAqV1guLMVKj
g4zZuBlWR2+Jo1jI5lB+xI40KtHMwFelb7BoYfjzmq1Qq24+jrtif2UrKcYSO3s+ogre69IlrbbH
bizIBmpCmOOKAO2CsIvDelDgllRCyH7n9gMuMki2gewifiGhHeaZMniiPL9PJOOTpJ/tXOo5ONho
xufixmHP8SRRLj8nMfxkndhKHeFNGIK4+vvE0Bmd5+WFhfwS450a/SWDISgAAzBUpbEkZ0hM1UoX
ScOYgyQcTMJn1BQCzXSjflsPdO7fbjV91thAbl/uC1IaW+anA10Ly5rKQ9j4eNV/w7PK4yuGmFJL
26/uLbDgXZUnjywSiA37GJenCV4w0KOC7RA4xJdjHG1cxu3jlK+nXXDOY1Acp4Smr5zP0eiX9k08
7k+vL5GhlpUZY3OEkXGzFv9mlT7vEYvCTw22fRoN4GzCn88japDhAAVJEdFxWhKXYcB/kpgJAVZb
MERao501qIzqMd5S3qO1yF8ycYjyH/FXKq6Oxj81Uc8/9s7u5sBraT08mcLO9UMh58LdsgPuWDdn
KI1xCarrmGNT2YyKnD728bpEYl4yTqQytgb5b98qGuA6p0M3wpd15jTgFxgf5rZDuRezxm5/3k+h
UAOxvYI5kRVkVDhr29MLQLffEPa+dOmG7i7663XqXBAiHHiaA2I7Rlh+i68bXXCjKDs/W9mBal4c
NjB2ucXXhe10ykRgYo87vj1rn5ji202PvIsgJblK3jvxkGgblRnEctNaS2WHQx+mtt29jbbLMJ9+
6kviNGtQlMqttluf/4nErha0PWSPOFSUdVUIuMyN5EvZSOHpxHTFlypid7fVzKk8cdgfFeb2Kqty
XKXIsn45AwAipidaUe/Vc+Z4zQgiNqKM9hGE4OqBX5g/5R28keOEFX024Af8YcsWzEyUqMN/sFbh
94Latx5eUQPuYWZZtzbdqh46fBBtO+HkZOp4Z/Ko4oU19VEcfPg2Z3Qb2ogkzHIU3+BWZ8RgMP6o
kT/1kdODNHVHC+MNdUC7f4te6jSopEw1J4xHBrraRHoh+MlGvbTLVQqnh78O34KkZUxDtShHvo5O
LETSiUktIIIahMBUgH3Vi6XTnjZ3FlhUTkD9bZSj2yd2pEArrQyK2w84OLxrrfIrSNmlcdoMRz33
geNZhuS0nOruCInl7eiiAnysmcw6i+tj/U7sO5rFLNSc88Eouc5SAbOhqKurnqM7hHUB6px10fk0
fOqawxrgvqx6P99RiEXnabc9oWMBQ0W6lbAt6Jbc6iDx9OOc4FSNBSqDpnMwNERSzs4YFNJqMRmq
Cttv7oNM72BvHeNXUjMZRcllcORjpcjkMAB1kl2X5RRgbpFwI62SaE35HOyFKP+LLxqtdVdnPoDu
JylSE38Wk1fFiC3Kax46V6RQM9LdV8m5XSJf/7Dm8yLkhvVO/WHHKDoPzEiuyshlGmcdih6XcBF7
EBAUTDG11fCwxd+BCuDU4x1rmymIGR8Nm2i1tOQRnH0gNd4xT7fEzXVi9mWpNGi04jES/aKWNVzb
tI4yf6FPaFiI+5xPh0wxFV723sO3XhkO0ip/yK6aRqKeG++a7FOVtfh80xkvp/ujLObOn/sUTkBr
E59Qwe8MRqeruxYOCBsGQIaeb2MYWqSpC0g6IBxVAbTuasQxVIbdBb8k+HZjU9ATkU5bupVdHa4Q
sxT4lVMyocdzLurDdZQutryq+Fudk5/w6yktWHimkt6oYqfgpvXru9EdYFTb1m/Gws5SqZX/BtLp
v7CtlnHhRs9FNwGHwBCFPepzbBEllPq1r7EwmjxEJbeTZgpBa6zMqHbdSwgrLN4Y1MwLiKDdvafA
ps/HMIMIVmx1SZGKGaffT0bEfs4YBpnHsmFcwVhYQ/7kV2qbSnSwqMT2w/njpGrBQ/VGe8Q0nIf1
L6IJWgf0ORC+NnKyfCPbHeq9AReTsvobUdnDxv5L5BeoP22RjZqVGm4BOY8ObC0PwWvCMUUDNZRq
Ljex3RooiWfk3eXHvpvhcbnqCytCo+4SBieoYCl9mVuOX8lMjx0q2uncRNvoY5bRHROJRlLtcRlw
62WxH11+nROHqQENL1JJq4j/M8cz3b8lFX14WQb88nl83KZ5eBLEPeuUy89SpiXdIHktz0gE6lpA
XiAyGevpc+gdNEYLMN+usO1SxSUgymhTuJN/+XDqrdHKWQQDvWURzIoyiN7cSfOhBwDiVAM9AkRC
WyvTE33fGXTPwOIKF5AkT22YfbbJ8CtG6SN06QdQdGmGqm9/q/cc7/OFnJ9vmufoypwiYMDjMDZp
pgQz/8xxTRWYt8zpSQFn5BcygBtZhq/aFWmAzMKiasZL+ASrxHNjZAfCMSVuUU8IPMpGVfMno4JI
c7fHKWFT0QTkuxYHzqE4NYjJsZrNOFiVoOIyhku0cExiuUNeLyi4kFklEzIuiArE8lhqOd+VjPh7
YX4UgX+4mk9i7jmOve5d2hvI3jsadJX1KALygxF1zWfJgLEKqEoLbJxjBuTJtzwzLMihLknW5TeD
O/XVeq/kfaVLIb8oaAgT/5BPN4w/SiF0uTNRdNrFnB/zLe6cU5s7bNVFvnIcxOj+c5726/+4NZKQ
8ze3QGyB4RzaKFzm3Y9RB33OJ9isrmnNiqKoYVeEa7RFrT2Tkr9omMrwX2HPlQTPoKxBHUjrkfXf
vLhMrzrTIT4AxSHy1T4s2hYMFgEIDjKhT7yuDWk8yIJshJEDpdSvTdMQoVYK4QRVXsfxpPuEjRbd
jXERzJ9xgs2aVK5Uw2lR8dxKMLgkX4WSYmIW+TcKxTX6P40q9mgIlrcMM3KYQ13sRRBZI9rKv+1i
74Xhwh7BptDAnp9yHGP0zszVB883UtiD7Ss6kXt3PyVciJNHmLBbbOeHrdX7WXz9cX1lILGgn/bT
5DeNUSDN5v11f1lQFmnDih4FCch3wkxN0SQ7eqXgXWuQUbXUzQp9wCD54at+rcYkWX+ziEAE9kS1
zOcNp7oZzY8mpceKY1KS/cjfjNvC2GCU6DxHvS16Zp0SDWAG8fo8ZW40ih2sfY/2D55N9BY1dKaa
jqdg6869ybvfmYPsUFkspAvbUD4nBbOZ5wVGrnDW+TpxRZRicEtvBtW+8PlSe8BYUTxJVySBHBbr
bvZp2JrJC92A1EYzt5TUAsNMjjV3VY51uSzMXA33rgUs4Yajny8eL9MHoLpx7HDBmspEwr/9RWof
99+xiusVFSyx22obRkeUm5ZHIKXI8zg70MUwpLh00aRK9NVdzUD3dh7hRvWRuL+0nRP7VMp9rAKt
0mUvRbWg5zAkaiejX54T685Q6N5mp27nwSLOrEimerIk//ItwmpRiQ9ndo4C949exMTDc3lKe5R/
qioSJvl4f+pYbniEEo/zV/QjhdT/+H6qmsn7LHX7/IDT1C2bMGyI+dUBXmSav8iFpiOp1IveAYnr
VAsKgOVts4FyRDoImQY0VZe2Z72GtG46UgCpmulll0dwWXor1TNmhmyteAio20fLe9RGwRRSugWn
JnUUb5WpV8FleVX6kGl61oOOLGxAIw5Gu6NJfezBtqcqSszgt89/4GRvKMtVjlJeDqjVk1IyaGoW
x5NIosXqAUjdAg9CuPs3eLob09wex1vBTj2Fpkm+arkM2gSdAWno9Sep4MEyVwBPzQFilVxqvxdx
FLqB7omX3odZ7UmhjVEFkK8ru9NuzOvMi9Opcks99gQRLazVLtjgGFcnnoJVtYBkxeBNfNl1G0y+
HjcYNup88oEbd37iBlnZQCy9ZIbp9pw3NAn775uFhSafeETmvC1d1xfaBB0aFoafi8gRr21llbTU
YkoHV2XraamDoKSOGEZ8vIMupVpWZYP4RfEUfaqEVTSLfcYLwjvGhPjo9qHmDGAZgbeYpsgs0tgZ
JAuNpt0GmjIuSmqtZRxFPPBxTOKsC650o9F/sfn/irIYsmhE+e8lEt6Iv2VJ7okqmHZMVKOPd0LP
RId6ssG8o2DjZ3H+SJ/ypzAkD9N8TI0SCs93MawAG/cYhXRvZ+b1+G8UfgqHYzta2iyncNZuySYD
/f4amAoU48CbzBS5htxd9GHNwlpv3SjMid6kJswHU0Xx0lIX6JnnBhuptjYOUx44aJVdFup3BeHD
f8cyPaAgpOpLk3K7dFKyOXxTF/qiOOKri1RvHyYr6bedtlrEWcMnQRjCODqoi8Fa7EM784OlM4+e
mR1IGlPMenqiWQra/68s70yel3frDnQwKANvrUbbqkLvOfV9uY9P3taM3IuLu3QI+47VgaLUYET5
HwDRaMHGVrR8ZA1JNW6K6//YpLEd41WFj5gnDLnROm9UtsYzfUcj9vNtiEj4ksr7b086bsZ94n1l
fvvM7d6sLPajGaeJSOJofQatkECi6d7TBre3tbcTCJ3NiIDtcSZwvmQ81nSqDAVDDVcdSQKyAqKQ
5OxIn9+66g4Dw76ryRtEiVJpj+gU7WrZ93Uu9HTMVn1T+eD/9dgrftuYEEldlhIkYdyf6B++yx0x
vR+krNULBp74h/eSuvlWgUk/Mp2dTdo3GpR7ATh71lbeuIlqk1WzLZDDhTn+YZYVf7GCys5SxFn2
XjaaN7z8Q4/9oHCV1Cau+k4k51AFK/8PoSBsJomvTQTJYZMa8OijHRiPntubtCPVo/PIBnRGE9vM
+VULz4CPUT5E2WQLb1ou8ZQusB/r+BJZnhfKbySWjiGgd7LbMOho4ewxUf/qqrqKzroeVAiq7Bli
ux48vlQE71s9dUNBGKRFw1a/hcd1xI4E9MqGpw7wIdVCoD7hgHKZX0TdNLqMBQsjbCtYkX6aPpEI
q1Stn6sCnH+SOOPsDx5df5DmfEAeo6lgzRabudCfQ7U4YC4vjuhJT7nT/+//JtTgm2TihR/VxfIV
svXSQdgzZvi2sA/qANJQrrmFefxVs4OlC9dK7kGarEio8Uc/QSeqgnvtUftzCNJlZlLGhZTZM/EN
AjBYR0RL2vQzYPsuZbORwu0PFffM7dz+LECV7DEd4adotaaSrGGzp9gZXY+L6vzSDwM+/D6z4Bwy
gJt3gmx3PRm8vLvVsH4qJrKNz/OiYjEoVSW+LEUJYpEclX64sF/G9kXhdNfv40UoiOj3WV4TzARY
WVlGNR0lyQtYlScb4xUlcV6AXZUutigmZSGOa+0fvj6xiCdAtd266lvrdoh63N2egtzZSg+AmTqc
U+z1nJYh8FS51HpbViVmbdsKLffhs3tfy6ZVHh5Xadtac88PMBAhRfL/xUn38BBeGc44QTic8SLO
apMYHPY074Rv1H4DOP/219kNuOYz8EHX/dTNSa4epDGrv+Fgp2rWTCs06KxW7+JqR9aSQ6FHUvL5
eJq1bhuMMUNj2fSXIaEwLtG2hYKWF0dIU3YlKAyEKh6RIhGqF56cS7HgMZugIF8afYWPt9Ez+A/S
MUcI0FqzvD3aOmpDOgip+alrwVMChr6qcs9j24gQgR9uCnxQ8OztFZ0VxMtFcRz3d7cvNGYGOhgn
aqr1wqAaqxfd7hXV9P5bm3AKq6TcQ85sgLPZaiquY9XuOOQNHyb4vOJRnkiGyXstOxIVdSaeWIfU
KibMwU5lAibyPVB2dUWw1LYtxCswSGk8rLPShqTs5xwywZ6OfBSONHOOtj33iNLrCJv1pxFtTr0e
gaYo7cLiKutpVl9qVTgWxICslHOyd3o8XIQiZAQI4UOrZni2YNfF+tN3mIdirxv3Mr5suK9QlU5c
DElGphyC1llR92BFH84/Qpm8WzGFH/iCf+yW514euVutKOO+rp5Ba957KXugNDGbDc7WBkFi5g9P
AlyHSCJ0UqbK+1sGxqEhkzCAIKHIrdJf4JXD7oM+KGLei7h0JojQyW+MZ1vG3QCN5eg9gh0x7SqX
ocKk50+6GcarhKFhhsYkLOgRkqcrrzxDczDzdGfqXfYeCZuU0ue791mQ15fzLn8l8UL+k33rcMER
orvRGaLidy7gSNZFxzkBVcxaz/0DWk3meciEFT3bge3XYz9/o7y7etvJAV/99wmS7bECZ2+Ku3Ct
UHF/AyEIA2orCvZ5YTXRK6y2yhjrq2j8DOEs60jLOJfhPIMLutEMVw6dGJ0Ows3EM4DiGFkKZH+S
kQ2m2y79s+IClEBw0qW2VpxKeMGWstCU2O5p3SKU8uUDHh32LWJYjknAUOxmakpnBm8J9dAEQw8b
mZ4DoIIOv2w9KpuumdT7oKeeFvtsxr66nkJaC6Cp1r6n+y5ud24l3OEXOebgGQhqxshxeYd9GO3s
fXi8HkeReTE73F7QMG5Zjk+UGWCg2woQ0PM5eJp3IoPefA2DJVz2RtgX6Q680E8m/NiDoxWRGILB
02/pRh0CZOQ4+S2enaExvY+ZHXEzbvaeCBnu6YN4xMhtaTUqD9G38aZafyrW98sxrXjM4twvS8j+
NA/DMK5RftG6txOWKqXZBWKeHcoYQmGAWuSdPokKYooOi64YDaOOe8WCp4/p7CTFR81vA6iDtHa9
uLxeBFCFdsjLXYIZjIlsSCv9bccYEvyhwd5ld0EhNkM8ftjqithnXqxBffdayP3kOWUja38d4huJ
MQbvcY5asu1w90VW+Bpk8GUnBCI/5+CDf+yZOU0yPJorvkLWu5pDNPgf4Ma5PvyjCmLPMZqLvXfc
BfWfDI0DMHY1cuGokktSjbwKD/Ur+kB8ZkwCSjcX8vKGy4VN4UfubpFL7QnAUNFEsKQyMIL+4NCJ
Y0tbfUkQEiYelVSJybelDp4tJFDIw267E78QfTvRsXJgOY6eKd4DTQ5JZN8tL489uPLk16gFRNIH
hw3NR5QklQTPauVitkS6BKExvx+oFk2iN0VO1lPTyDLlSFiC9ZTLxdxmntEe/U/UJ2BYdx5t/VwH
bhOIb1ipz7uj3liSGeyE9ISlPBEXLK0F0A53owPIgeCVPw9PA5kTk4d1Bb3FOt604U36DOTOjmGs
e5VyiidiXb1V0fMxr0oSxxbaw7KvaZ/R0S32io1r14dZJU8vz3pNAbya9OlfccwwT0VwECqsvrP4
BPeJN9Rkj5bKhXp5DAAFTTsmrIqlMJ/CfDYSXEB0ozwV49LVmMXS1bR5P2YoGUoHZ6+z5Lf9g84O
Pzv4B+RgIbBbyONo9Ax7zbNlcHGpI6dUBAisrWpqBpQ6Z0TqImy6dbwwzFFx4CDy2P+oH9A1QyDI
znKEoKY5N/q5HztDeq1G+c4MbU9V+7HZrup70364GAw0FY86CyyoSpolUic/ALbKbRvzB3/eTJvl
zWv+a1YtCMLQptCeY2+Dts+Bgn3TvPgiBMAV92bg55HHnbYjJ/yhwf9gCk6bHD9slZ06ObrE+RKn
uupiyY/hRe+BYDLHEIkHtfE50s0SCYjtuhQhDEjm+Ya2ex1QaTo5lcRx6qrrd3k9g5BBpL1RzR+E
CZsV4Xz352w9EsXPdcd/vCAmU61f8YfKetpdE6umaY+dNqpraKCzyRaj9Scdjbe547Q4A1/K8GKo
e6UHMtNsjWDsH60xL/9oGvFZ97ar9iBqwoXZCyCsMeqXM/dZjxmOFXkrib/0nBoSGmprYDShatAT
152n+qebIfOamUqrwxPt51JAqNzQ3qC114Gt1Z9yO8T1KcNMCrzgvXiE2xk/AV/WrmI6wvxgeZfJ
VdLu8X5KOgWBL7tYPIQqiDjdLsH859FUxXNLoH2yDXILFUqsMubVrOnCoB01Yj6dxOj4yi1gZnCj
KSY3BZFEO2gliG1264/eKwCx+9busLfMGHCuSS5FVBL6gmOpH+a4SCoJoDpY9P9uEzmyl8h8sN2t
AdvLQzJ0DCVwQZH6S8tG/CDdFJSUdtTZGzsaq/sMR0SFIC/Ye1XrlXsqIE6sF5PcEENBQOW52Wp7
BAcG+xg/S2zFAa5EI5VJ3EnBjGwmUi2bi7hBdXZ0jbkyrKCdCkckeZYD03T4CNVo+LWf1gkiupuP
iMXwg+cXJ3lOxJ95n22BJOeKIw3gscHGnjLbMsjZagQUIL+QcpYUgxs34OFwlf+zKVkr2RiuMZeq
5NcyqS11VsLog+q1X9A3+3ZV790652fFCTThV5/AfO7yvzIKsMT6TONPIgRgNm+/YZ2gWs83NpmI
MMNP3a0A6p/dA0kV73LTm7bAKKo1qrK/AzoGN3a+gET+yeHmgT3YU/9ABbYX1zICb9bSfEwPtkJc
x8Z6GZrcxqR7xdSf74+TqwaUsVUYaLP0LPUlFbvmpUROTxukyOfGRiireTbVoJB0s9NpC4idtslz
B8UFtLukgE9o5yeDT1KDkCNHDpqQ4EiFUWp1q5v9eFbTC3hAuWAhqfxb2ooRQxEnGAZdm6o7M7JC
V8R75KQssnJ5re6+JWS2PyD13E+s7GNK3Pbdn7m6yizEAtx3/VwiKDS2IHjSa+9LLX0tr7ImcpvY
R0Rh8Bb+4NrIYsePHmtEJLBSoncec2vveG1lSGnQUSxi/eMnj3ePuy5CVWlDr0Q51ngnEbcaghoH
uh+883O1e8aKSJ+BzofHuAvxdEdNcoMWEPW0Wmqs5152oDNQ2vhaiG/bQRnq4VB2aBMMzNctEEyn
cU9GtQU6wQrfRGd3fGryFcoCgWcH/rKXYlPg74nOi6ZWnOihhxubgECrhN1rLUrdbBDJwUFIaX4X
YfaS1EAVJ2UjNLllqEzpGLgLRdzw8A9PYvHOUc/6nwnC9HT/0GUTsTwtJOAgLN0VlMe9BvNeC2Hm
LzX2DyNs2mS+PtrPmHYa4owXJFQo2vEwpcSGJAcmJta4bUN//2IeXLCG5MLwZtMnOvgqsy/A4YeL
Yvwgn0bOq7Rk3KJK2yDgnQcl3dsdYAWaiaBrHlTwkwOGgKAiDtowUect6UxNnJnh/2iyaVoTc+I/
uqUygb1S71JfOJ06SA5wi6UPbU17UFOFNMVUjUqNrqSL4qfb1yaVFrxcMtNyLnT8nug5PLtrJ9a8
yqIyj/sjdh5qpI5GqT6n3Hh5hFT4kmE8bmGzFIGWIOXbNsH0p2p/jUydrjIraciUzIcNKy0HBZR5
8GIkLSYU0HoT26K3My6xwkCLN0fy5hWUIBBGAXjd6NSuBL/blvxmdWxkDVlRCfGcfQ3Mt5i5lT0L
vb2un8jH8wdx+mn+ibXMwtIP9C7pb4LGNzZB745rcadzaJKk6PrtgyI52RwkOUn+CVCbsHp/sUlH
jh7VIs7VCs1fieYjCOGNP5sFk1RSGPi9lh8gki+nCv7ovRcHZndvW4fRkutjGDShOYK1z1O5pvM6
ZqPy5b0ejfZxq8X5C+M53w/nHoadxwhgEF5MM7GONnU66+62A4l7pu3daBaijZ9qb2Y7Q8gelQYF
36hU5oUD26MWGIJhfYhMBBPUavyUrkhOT4SSmykhoAZKqUGmyLNYl/YSuQCwhQ24K5lxvgme0IEu
QvVJY3RFmsO76k/FmurT54DobrBdjmYJA029o3DMP4K6QlLiHhJ2r+O6FtLFtQp13EbMKiIWzDxB
qIX6rWeZED9PJCV3bkbEXvk/zd6g0XpavjP1EpqCU8iJBaQ64E8UC7sT9/3q9z5ZMCqygS1UhbYW
eOJd/2tmvWxIoWpMoGNyw5Q5x8sGaibYGErEzTyZb+3ZEgf8QSz8NNVnR5xUj0Ipz/fqZocFHFhw
PxU2rHci929MW8JFMw3Tc7IxRRHyKnDYMMwfW1+k3wegKoeX6RmB5fnd5NxY1I2cDthVjZW7xcvY
ozl7IzTuGfzQ2a+j1biMpyv8oL3GKdO3gxifxvxTkFP+AXEk/MJvUHUg9E/xjFUzWh/FEAeWUPhJ
wh7OTwBFfHEyZ6bg8/9hi93DuKZI09pgbhdGcRjREBPUkW+6QfNPMEZ5pjuq3qs6vx66rB71rbYl
VhRHd4zIrKwlmpucsXsUaPAb2mAmKF0speku/oNq6TNYuuzQ+Vgspo6M57lVZv6jz2Lc/+vM1Jv8
V45Ew+xNtf4lcD957jz/PbPn69HdQv8xCT0/EhXGDIRsWVeRHJeP3MwDPXSvzX1judOXzdXN1Uz1
Xa4D8yOkDav7tbJxjKPUSEGuTuUXJZj/LSDPj+/5N1bLePV8tewCrWh+LOZwOFMV7kQ6suu0bI3n
tcoiOsH/Qp1+FK+alj+xeBvM5aYhQc1WpV/M/95DZmWOBVA6usjHWvWb7GuIRDV/BHcZb/gKSofm
Lk2D4Y9Z0o2TeTgfysoknHEW1fN5GPHAEhBZ/cuFI3d9a/7/ntqItl1RIEAL45MtJCaAbC09dCbN
SgsrzcwGsdm4KmPEoq0oinghKvfcLwvFLIf9YGZ3ORI3UND0We8aJPH+9hOajOntMJBnQz21ezD7
7JLH9QWeP5TzKgBS17Kzkam0PvcVKohOU5bT5En1OqPPYhRZ5QuN4+Gp4dpExYJ8fP9hwboe7SVq
SuA7nrwmS1w2V05iPvLm+IL/0JHFhAd9/bpKXuknDIeRtXIY7IIwVH2QVh2ZVDhx57SKLDeQM708
NPaKH7DEuvgMYp4+ey3j5X0WSE8U5Icjl9QmQC0kZtpx6u2xTlkmW5Gh4c9R6CkEdLLl40RjcYc7
gzp7mGDYMxIqlMOlQVCAeuGK40WxbeXstM+IQzEpn1/km+fcBb0KPt3TPJcQsa0WmXSiEZ4j7Uzi
tLbqOeD2dKdgtjdKpc+ffXpPBeawdy7BzpxS80kG0kqDbNlWURxtA8OdT20XlO7R8iod6Ql+p8PM
iN5rUAntE0of5XcsG/g+P0H74csAA1bXjid1Ktweh+mitfL+C3YFVyYTmAkUfuidPAz8/452W2BW
9pTuB+k+BJqyi1e+9PzEDHfJVBjNy8Q1avDX5Ux+BpJgQS8thaaHin4aS3MHCrMcr42a3veECKUy
MlW5W+zFBNd9gjxzPCEAAV1SySgpg4cUtybnugrKudrcJf1HvQZVCqBheOTG3cKjggj4tBkAeT4y
Jn5jXGvXyUXyeEi8WXZN79TH9tjSThSYT8EaDghg09076OqSw7qnZlN/XXGf2YSFQwORMCyDlr+H
Py+g81n0D/LHlYUi5Q0bNNOAOZL899ZgRg1MLRCYxxof5CHzksSA7caxJPlZ1znfl4/MA9JzP20C
RUbn/2ko+ABvtoVJAb3uHbEVdEHP1E5wKrYtnstkORDxrjKYsLE4pAm+kI6XS2I3Mv80qvJt3RDY
rRXc7tG9qa2XtGo4Spd/Bg3Qd/4zk9GGUDyRlhdqmhfpLS222Rzj/oLd4cS26fypHOArw03dF+ID
USqBZWB9pCjF3/UwsatQes+gGX6sTl/mUYbaG46Y0gDag9NKOZ9hDyhVMDuTFYuBURrQpGSlXXCV
4Sew0P+jtPtt+kpFujDiRMBrS8k0xBiSF4DFihbPWAdeif7u/igYUu9/z5TyaOFM3zrHjEObcZzD
8JeLs2BolV3NtPF9hqXHImaIfmIrmhI1XHSvUJ7G7JDjAOGCCQdalmEbv2nmXXYng4aLY7Cc+Ukp
urRATrbn4fC37GgWupHvhsi2PaXWFVTBF9aN+eaMrj4z1+lMWGHVMBWDoimLO0DF5F2c0hYXi98n
mdwpc1wkRVMXDn0ndc9HPiAw2THltY9zPbVZrF7h24yBAcGQXqDCANnSODXJqoK63DYe1spQEWGp
M6pCdajedGsXSBDuO3F9TsOT1zInmaL/hq62SsivWM0bwZ5iQJxwlLyCnXc9chLq8sT7TEeeqW4x
L/74VNdKvwUDrWgErwHlA7dMPL3ewZd3pdwiRb0g3pNndW7Z5E/kLFup6TxiZyZOuPzGu+XGy6Jq
ym+AmNxTRicaRQOzpGeCeNn7+TuwAwCaqX5n7NSsvoQ8EmXMZ/92AUYGSu110ZuXFFrMJGuP0oIS
ZkbNj2Ym3E0f7SAaFnKcBouh0ZgjPfGFzxLQkONSheHLM7PYLjNsc0Iddb2aWipf0/drcqhku7VS
d2+n8UJH3Kvg3ZDvr5W16CaS27sTxv8Kjw+PE5XaOo/49RfssjsyRUgOPj6YCYA6YtMAYPN1zlwG
aw6H1Otxc6kFeHthswzA4F6xE2sQfeQtdBvRF1SgnaTpWVUaYSRD+xuOm2m2hvU1E+ja22kNdsaJ
w3ws0i0mRBKAqzW9ojM5KzWk9awBLUM72wtafm7/FNXRCv+TCdIG1crotsGHpHfr3gSQVbjCm8Kb
ysilwcyyzsKfojqryHtvGqScgGXss2FN4jTVyUqW46pyf6tBURz9SwFvdTfooNIlSCKnD8no7Y8Q
UZuk745u0W0bUIq8fFCZXkIzspc5nJrk3iyDosoPXMbYdH/XihSZPGAVF5qh/M+yRKsmzyOfLs3o
xfGZ+DMApZeTxKIuqbb2NmroRoU/Jy2Syzt12ZFza0KjxOD4kryBUd8mmkJtlQn5UWhPUse/4WJK
110Tus8vEC+qWIfsF3InS4jkDXTcDjzYvS13lB9PYVa5OlA7KYxH/Z1YJZEKdHRgyEOn9uPLvDIX
dIxwvbh5/VW3nd2cPkfT6tBAyrtBP5nxzPFq3QsgBdgjYTCyo6o/1P1WsEJFTnv9PYDNnlbkJzQk
In+LxCa6Nb02zR+jIE2JmUu2hnlYO1VgNc7BSmE246qufzVZnggCi6gkHzKqKHYsfofp5BLulrzJ
BcPE6QPTHrzBoIbrs4CwCG96cZMGmKCTubC5LmF1SINE1YOQ+r4Gu133437BrRnT7tBQ+k71lc6j
A+AH5zsXvtaIXUpFXQdrp70pSZNaElfqSgpD/GBy0VeDx4atr9nzCgP+0Da7GFDda5wF1uhBklzZ
Fwt7ASYDrRYRKJxuLLDFB5oF+yib+8Ts2bIxqJ/PYVE/xNGb49mFzoxMbbuA0CAkDwP1b+nvIwe9
hkNhfaDgHBE+3zaSXWIgjDDLast3IvwdCAtyL2VsCSGX1WvjIezCBfBfxVC+fiYnDqPF2TwYGUBM
RWElPzcrY9JgLoIe6DIh+rAXrU9uItS8ZvWn2waRZTHeo8lDCtYhkwnAGKT1WSmaDSVOQ928UyeL
x/GqEKerK/WI0lcqK/qt08GExjOEoabahMxESTOCN0GvUvrc3uotaVwFWaXjjX1uLWf/OjdetlkM
514/dQgNdZC1RH9JDEOMLkurYGgVCdoYSlzzc+e565zDF8XrlrimZ1RdfefeRm4HgtB3E6upMNAP
qUfB5PYRvWmxJBZfsVZBhv6FhTMC8F/xLTF52B0NTYHa6gwZ6sClJcZFPH2Rj9AcYAQUntjbZHd6
E0u6a/laTGhwRX0zNt60OrOIFmpNNWxWj+Pl45TEHn7W9/PQe/EC0AbDlbsPyHc01NNywFoPKe2t
jc4E8GUCI6HCVTvajl5XpGYeQi3TrExEX4YLy7VZdSF1/eusftmJ5mJGLsatlLGStsLseF2Yuy99
hnKocKGnC09fYbPcG+Jh/y3ltB/O8fr/U0ls8cH4JWMW2vEPfX7Me7d618/7YmW28HSJYzegWTcJ
OeTrzh9+/6rDKIVxt81b/MYHb+IA/ebpKU8Ea1df8jZG2bknSxX53DHlu3/AK+lnSNvqxfVA7qKx
9tDSafgAYdRaBtZV+DJwLwCNpgh50HQ9ryASyW4sQk0LFx8hKYRebYLcvN/CsamMQ30vBHaqrm1Y
2ro7MwGZfTbUPJJBNxcTPLxUsrZau09pPqlefT7JOqOF4O102qTcCt9gq1izCU/XL4oVX3w51geo
tbHUXULqBNf+E72CtfHQOODgF61q63NtDeXydCY/PZccGNsfo1cHIfCXSNhdoKJfy8/W7M2Kf2lS
dJ4XVSlwozDXSUEdzO3lx0CthJzXQ/vKR/SaeOhbQVfRy5qZsfHyrVeFwRe4mLiI+mTMFURmYNJq
0SmG2+1bwVkrwERDIXQygYK4EcyNKMDSP1PyCnZbJDdS6GVsijnTCpwQCqUBEkPg1k+2qhR5sZXz
MSPQADG3tFFUAjd+AcgfsmJFEiiTi1fChvdvzSV3RU4Advs1XWRQp7yedCLNs5dSuRsJsK9cpGU9
MHiT1Elc2anGasSqbAksSkemhxcMiFCpUpGCtggqmSeqKxVJlbUUitr+VEGFoRIFLHTB8JGD9Pz2
9oJz4nzaUKKaVtenbon1jsBHReJKZyj7CZJBvfN3xKtZbasdTaITMbWaoRr6k074OB5mgK7HXFtI
cDgvaQPdUZ9b8yr52SjUkwiODMUyLVkXgV3W0kxNpQO2IghDmxjgpZqC/Gb2UscEEAY45TauVr8+
HtxEccpxmxZBuAC/6Ksm5V+RFXQcA1qdzN/6a8N/NbONQWONdEluUbmoHnudTsYTPYJpfQ6pyQf+
rOhGzOT64XeUI+csD4631fyO/X7oumfinmZEjZtDD79CoqbGaBAbiUoo/r7SBW2f70+1Hx87ZfQd
Ghm+nkZRvxz8JsRM/ET43OpBWND2g/qc6hkcC78MOHCuxzYpTcG5XNOzgLoRI+7WyppzHNK0vU/w
TbqHuoZHpI4THfDZ4Z4WNmlzuzN4XgENqJspb2dyqLJKEEyK5+YqSy61GZbtFvbklXWnfvYFhl47
a+OpEAx6Kud01BUio8B3UPfJ+7lShxYtHcT0alHPtYpQAmVBVKLwaXXbAe85cOaMhrizgFqUD8Fl
ui+cI+FNyCGcob8+2eSFKU6M4/OeuqY2cuTM09fV0QI8EW71iSZMs45+A+wuLXipAl0QmhmDVcWQ
SF/hCctSkpXQD2mfdBxlhJ+/2l9aAJo5ByOaTaPlp1xJgMy/cf7V9052W1qJIc7e8q2jQZ6xv58t
0e/63N0BAKu/SzNQp+kZu0fUTexVLcQhxsYv+xVCYHv3qhJ9TR008vc9Wz2OScpV6NH3UVi1DREn
80T1pr1Nlt7+Z74JeYI6RqBxWb1iQgUpR75zk+JUHlDGECOoUcIYvtKE2F6IaGGI3LgY+1RcXJhr
37bYSNzviSlDQTn/TcX+W56Hfj7acWUkUOCOqAwJz3qifGPcPtUB4cs8cmY8+EtRPU4QPIaTsL5x
L6OJVrT1Vz26ha/DaaeMvnj1fTGIk/p5F7AHkB84PlWLD10j8s9R6zRXmhb0IRuJV8rE/VRpJBV/
8yW9Z5BWY25NundTyRJble0iUX5ecTi/IbvnoU+7viL3FgiArMB2tAF4OHhLlpbXK7+zaI8RNzko
tYrtDEJbUBcLwcMbeIy+YRe0I/Zr0ArGfHfvcZXU8f7mrh/QYyFzD4mz4SWbTWnhSE7O0bwaP4PL
3bgBGFKUJc5VrUkHR39cnehZQyQXXQolAzgyTeLJGshCv1zuL/J07TwJ8KdNQPTE4AXnW9VhSC0C
rsz0XjSaO6oqUF2mNr42sxMZWnS2KYYutpgyIL3ecfR3HnlsMKx6IEJbTP41t41A6OWbaA6+9D9L
D3B8qme3H+5sbEgQWCxzzdoqlJPbbPlWyLMIKW9R6Qg3GdUeJB5vzL4j7rBEptu0bhWq4nQqHdMf
ZBkW+PLEmbLNrX3P1hDODOU43kDugmNoSeDWlsSxcC8vu8rH8rDNjyG0t5HEeVfJf1StyXXLyQ0N
ZcbLjGGHuqCFXkIbha8+Hk7bJrcqNZmihYNL+LAQyyeRVwq5WIH4lxk3bUjKvCZ/nDWOwMxO+Ipx
NcHcnAPJGiTBjWZN6pEF9ydOYh031NdCkum0l/TCkSZFfx5XZVfAq5zq1k3GZy/Wr6A5xa1ESzN3
tcmfuPSrYVziitSVkdwRsAqG1qQBZW23gixOjFDKhEdy93ILTwHBAxMvkl5cxI3QFW0C/QdHHmgq
hb4WSicF4oQrmOhAYYQD2UqBl3hBIO1nSI1EptSgs1SIWkSQbzk8mUGUZCEYlOOuJhNI/F6X52Sz
8tA2ifDEx9XtwwXD4EDVs5nHaXBnjfyZlDOnytZYQSSNs4Ei24Qz6IhH6Hgj7TMT5CZtAD/q3mxK
ExNrwvg/HpN1gXM3+RB6ZAN4X031Lw5ja1sB9cDgwoIvDUbKxeXkAzotjF18aCPmRL5NkpQO5Avc
MveMie2iozhY9m4ykUqEL41P/cU3oBQYQ2wTLETyjSb1iR5SIV27F0xFI8Ih/2tyYSEfEHQMTVlS
6adFV9vOuuFXNx2Kt/PbUAM5B6Cp08ewXfkZW/01k85MVIcKNN5vwBPjrd2YiZETPeG0FZhJSr4m
7KP/fvBcKqJZ6gECfibOjMkuhDhAzbOECKdkXBCQPhpbNb1qFvtPjcrvs2JBHbL00gbAwfEwvXVD
VBCQLhONqFFwkdAt35+se6vF6hlqcSs/a8y53SeJKmsNPLB9EelwZCvWvA7ZgQvgTR30nBtHCMI9
/eRSNrzRjN+4TDrIxw4QoGchA28QHMN5QGoCm7bi6kZklJfTN/5Wk5+AOTVQQxOhN/XmiukAttuj
6UoCIygNVRA+RhqmPpABeGErGsNLrz4DII3rbstvasLOPPnzWgmupchog0HWmNsXAf6JzjhNZpC5
jzhOhZIIlZwORDVLT9h5aFsfL0ucVnof5pI9no2Sp+7gwLKsLx2y2xDoco90KZWETgy+Gkd7m/SV
JWfgq1OgW56mnad7/61QfbpKuWoBeULtY+kQ+KXNHZwcSeK9tyNJ6CwkCMyOaebYy7c5uZGl0hAA
G6SdlEVGtGlL7HB9nSb2dGnGzNwrWyc/7/DFDr+XE/tCXXKDSWeoRqBfZsGuKZnEfs2f6jJbkz+3
j1m3wUgUEi2LCNSDCwNHNi/CSrgukLtIo9Oyy6id4q/iQ/6pfeBhfhnWcgKFjDmFl4JswMqrqeE8
HtQ8nElUaKlaXD6so8EuSFzAZ4LKTf2KbgdXiMi3koXmbGZSY2ZFc2uTwHRAMLTAu/HEhqWg1kV0
J7ajj/CzI9QNw2byvFxam1G7ntA0s4ELV4I+LGCnf+jHfJxg+osOu9ZO1zGIb8fzZIQdf6jcMZJ4
0zXOGEUrrKezj1xiz2zFQLF67z2BDVkhL0HHesbWXd6e7nAa46x2sr2cnIWXB0bd7vcCf+Zi7nYA
uvyQrLzO7/Y5YSbJaKLHo8qdTuedOHPQyxdroJQUd4ygpOQwI9R9Ny6QNOoYEgT1W0bb6vHWBUwV
gOpSVLH/qXsrPYIMoMxceyN+FXYMb9lwSbuboddAbzV5BHkbdwAzREavJeVD33FPef4DEqzTlSi0
R8JlyRLMUsrCPAmFPxjRAk5PySJs4rKxSweh35X0jTgyVqUBnRY4e86ZAEWCWS8VYhK0gNxF6pAq
FOckQZE82oo/Or6trmA7gGZTiO10T8n1+CZFkGi5VmtbM5HRTzilSW4vOMHCJbjDlfy9ew/eRPVE
fYqPRm1R2+TvOaydQ8FXk+xluyQM+vBwE9A/MbQ+W5XgFYwE145iEFUixZMys8Z4hGMDhqaJFDpO
NXs5H+7LyKlKOocU5ZxpztoSuslK2+n/uPATlwUwO7rQBxQyQuh8WI+1shJsHthJxFU+KCSrP99j
7NRvT57yVyb8gFWeO4Qvf2OZ5aQ+9o1aVDDlyF8UsWhliu/QLwaEq/nIP2WG49N49HfCRWE/g6TK
WSAgdiRKdwrYNRssTc6RPWDJIhKA1t+eNRwQb+VBtjqZFtTnX/tjVJ4cS3ZW5w0sSGb3s+UgtRlN
Nx4Tr3LdmBRhExxG/m8c/esXSoI2dSX3z41j+qRxn5u+5ec6JcDOfgKK8ruKE0/5gilO5pkeVw+l
kbB80z95B5p25BEX9rcqanmnu5UBGPqkfol3PrX7Z4VYiVdeIJeNFP0rKegHSeBcQWLkaMveAwhZ
7caY5sRokKjaJkytyslS6RzxkTxJeAsOviRVgC2amRw08XLrkf81MuVy4gv+mfkwltskhwv3wryp
R3Edz9KotHAI07h/h4sWnotAkUgeU4eRETGRHS3YBIhcE3ZyU6U00zQIEP4eFHbL4+hqnvb9iJVS
B3i3S7goFJCtpzFhzOSzUdwFlScLMjIMHTP/6YxSpssjPXadXD19nntV8Ia/C1/OPnTMivLC05sL
3CgnJstSWlBGMEixKbyCJ91Mr+2wWbZ6pFvi/G7Olzriw8qvmzUZ0MsawcygnptHB66cpRrSBjSy
sxMIqIwQCJ+aC3OMmHgBVSreVDsUT1vJhB8HTWO/8RkFDApLiPg/cxUijHA2CtLaDDFc3qjdy8cn
LVpsFrS3FZZBWO+eIBm9hgo+bD62mZgGUf3a8t0fijvPyfxteZI2DJ9uZ/Sn8777TFHNahRxVt6X
QzSEvsCSLxFMIVxodVMCmOtWbsXF3IOGU/bwH+g2XksmrDwezoYpa7cgKZGtovBZUEyxBUhkQaz8
l5CHwj7h1Xagu4M9WDAX1HUo5WM8wbficj3Tk+zNWu2sqdxyq1oIHDL7k6Q75Fcrzj5bqkeV+6aw
j5hnXCV+b1RFmli1475GmJcs0NHK6svHsmo0SdXB0ICQCt2fYLFOsjYnEgmdkoG+QcHRZ+ZIrY9l
lNYA6B35sSoLA71O4+clQ9wSYwdSM944ngKHdTu0Z92lcpUqo8xtGj7bxaKv+vFKA9yH/Z/N3LBC
veE01QXKWapXvNSvfm6gedbnISiC+wXbLaNL2eTHwD40rieQ06ZPJt3EaPqP+gKt+QyHxW9OCUxT
/2bCyX1Ho8LTeEFwhxTgfaIDeFuojcaB+2qUsdHMX+QQhfQIO+2TXbGrgLCzYEai1bVhHvKYRxaf
+3+zK72eUohQ60t2gmxoDeXyfFOQ9287kfCUibtiHe+grQfSoe0vjLeP6Jo+K1hZvhrrfn8JJq/6
S5ulTmJ++9XFVRoySwGZkbsBpPTWreznHiIc3zgWMwct0wOM4wL+j1qzgGWQwhhRQgV0KuncgX46
IoZ5ex4jOpLyNFkB7LrvmhexrPAHvKTFw39Gj2OjKhYO9zgrr+hpL/j8IylmRjh90gvrvrnkUfjl
h35Y6k8Ens22ikukwOhugtMSDkLfi1hd1MguwwU85Oy6b79gMMns4zL/PYJCF8wzON3eUxMQFLtP
NgoWlx+lHhr3DBITMhUC2BCd8lgnTDV8lxAPMiwVOqj8PsYiXSxftQAB7vpZXXa8BnEoled03acd
fN0gqGVkvkQ28/SHMbPxVxywkXOAWg99+rODo3YEnHveWW+yV8yMHxacvTN7OLivUWfUBsf/Tkhb
pxZMAHQ0wSIQMnfA1hB9oXmufKe/qMmbcfUgepYhvssW97/U1XaAAU3C/ny4M/t1HnsrLwQgtIys
hagLXWZE/F+EsbrncANnGXPlPpxKR4YAlGGnK2+aooXNsFPnZhAXv/wPYAcR8c8dkmPLTPrkfE5e
3B6Ciu6AP9qlGfgjXJXu6ueiV+EkbqsqEOy9+rgtwYdoYC2V8plgRGZ78sp00VCVH6wdRPPy8kcG
P5tpu0WnLfWLXXysx7A/o2mPESXjoY6kqclxnYNic4+LgIn5czrO4mCeqCIZADJ1IzpwIsw0nNaU
Q08KK/JFeyeKqqRbgRlGjfW3kjvrSLmCRNAuH1XAxGjQMI6kDqZHxDTHOI0Gg+z2aYIIAIqUGOBw
DBuodfst5vgisgfN8YolA/8BVdj9yQCfkxtpZnHOiorLQA+hGzrX5uaxsygg24DUKBPToDWPwzph
41LTEvBew0ltnbvsjBCqrCYLN5POndQdVAuiwbyAQlCm9vJ1GdfZ99+/sowIVfS6N7GHMtL/XCdj
vjijXyHb1aK7ptC0Il00WUKNxD0wq+8yF5sTwD1jPh1tNBoDuUEa+xTGEGbt5FmbGJLwMxEG6+pt
pEVGerMPmKcEh8KJgKu+ZjqN7cKGsMcsYiKTFxiWonHwnklRHU30+JhS00xfkFIueq2uH7rEmMRv
AVLsIKSE40/YC3JWicANmm+ML7grB4knaO03/1xSyK5QVQ7x6ZlUtG23eftsq0gtdFj6NPDbqmi/
1QftJnkVQGS42zo8hYIjQgtOD7R8lQInkyzkIy1oVzIfot4tdhw/LlwHf0aWnJA/1as35P3ENLjr
K9NojhPCrLLvvp8DxattP8YPAJy6RdrtZHngvuQyqYX58VwIPYwI9Je7Jg7WKEk6ue2UbZ3dh8VP
vkalTYaw0GdVUEyZSdQ3VRaHiPiLwjsywHgdNWpHIxbrqboTb+iMrk8vNSI7e1n0kjo3QI0Dlghv
AyQa7oBcGLrULEj9oPH2qALJwYTqR8suwOXT6FIBWur/+7r3afmfF9s5NrmadEVNHOrOYjSI/LID
9xLJpdr29nRhzMT9nOQjpT2zvjX5Lf0DougtDw0jJIcDdAJP3DhtAgXd5ba3Ko0US0pLONt/aCWm
aYisXcdvxfXs7ZBwA4R59nXkEcnk+3wUkRbFp1IDROhZmVMB0H/v/PE56hpdTGo3AJ7LRkSrvcXK
7lVD6lh/lM0uz6QbSUagKD3NRNxzl32SnWROzrTx7Y0x3hwW72euIagB/rDFSaVx9vvQ/OJCrB3/
NuDa45VL27M8hzJ8+lnlbsO/tLMkeZwRAQRkhvSCxAmsuj2lPhvvIv+3qhoFbnB+zqyH8InSfJzt
ZTO8qUvpuLaE6aTfrKg8qqBSkHW0UCHMRJ6PzkePLUq5s7byU1iflphwgAcLVsiJh7+zAaUQIP0i
ZZQCrmPv2ZhZ3LjYtiITySHyuLxAEnCAnwgIbzCaIDHo3hxvJnEepNCwyWQAz7UO+G98qW7Nxas8
15FMyvywLJvGeNF5I4QA4UFgaV+hyXKKPaiuXKuDuqZowfFT7KZzrgWRToZ24Zsbuhs1zyGDUE/z
XG1ACr/Kz+LbcI0wxy6lDt1SwiatCs7ZTypmxC3DJy4qH07tiyg/RQxhfwSvC5/hVNYWHQje8sL6
xqR+xhipL9MAXsQkPwAabL7+ClKFEpwhfpCQBEiGuGZEbdPaUC6XhXzJPzeekP+dspnoZBYFMkgY
jnqlOkjQr9r7bHfNlmfjSZJ/rmZLtTIJDikaK60CQFsAhUb2kZBTGwlbaWug5ik21TVB48X3LKb2
KF6wbfDd9TZ+yXNF5pLuXiprG4Sf25tm6BvC+C8eK+nx3a3hr77ZRQL9c9Lic52OU04EI8CrHAJM
+KS8A7/ipJwPxJiy0YpCwOTV9FKaNwuiTb27SxrJTjyofK0l7HQvTB5oXljrKMFd52yqSwX33UI8
DR6KsAxLsaGNfAYw9/6vCw9dcP6SlA//qHM9/0SMMi8TV3Jx8LaMeRCrHgbAkuuX+G0H+dru6TYa
sv1H6DOsJ026vRNXbAMfptj5mnNVavzBsKb8svHWkeC6v84BUYYbUj6i/oFfsPj2typ3FJUARaax
5e5DAyyau4YxUwPOBfuX5umAU7KsXKaI1RJcW4+pXToq87W1+hira+QB2EgGlVFW3kIrddCaiiCQ
QXa8QuKmV+tHJX/u6a05K3v5zd+6xcRdhtxupZXmzceKXet1RMHDVzngbwLwLCPkD1LZSdmShNYY
rmdfISJO0JziEG3lHquo2SP4PUacm7xSxBZRnB8F/sbihAKchtf4wi43Xwezms1ZIhSDo5Hh2njb
KE34BxGCPcDwEvgqzP6nLlI3Z0lcmqdN7LpmMlOFr4TQa8953ieXagUfNSRrWbpo7koqK1yaOZgu
22s2CU4pQL+tqAP8/YNKxYQbEeYqrSFGWx5idihJT25OD4FIXwbpqOAlzvqno9ysrRqWr633rhgH
kn9F/rOXJ7RDFUcc9PV+gD7Uni0HKVEDH3C11Z0nWubO7ZdFekXuPx9VF+EQouw6PFvKeyBnari+
P27x4NrLYhAK9sctdBc4X8Mjj/4m/MjyPWUsGRKO7d8JFpZ2/fQcQ5BpHxX3yMlhShehxe9vMuvV
mZLOjgxtPP8NOyAXIOCS/jlabqKvLnAYRFr6dzCUrQMI7jko3btcFzPQRUIwSgj7AML0ECK7rC0n
udcZRf5GztuN/sFshyqxuXwtRMjxuE+gjotIRVCMoAUMO+RRa6VxTbS/yHizNsWb3ug/I1aEjT+U
mnwey7PyHyGmQS8v6heEEqLTNrraglCh64HV+iepJvHxRtOl0Mw8ncsDv7gkE40fEdYDOVVA3XgR
ahCsRebQHMgaH+E+/6g8lh1xVQJjaVcb8KETlRTmAObfQffPTlTPTso5EJtQhGPe2BBPKI3Uj2GY
8QmNICmazlWcZkHW3e5jafpmGNDjyXYef3G1QQ1R4p4CftC72h/rAjxHb60BV6dBZ/YBIQL3/6Gm
kZQe0B5L4MsDb9Tz5XMh2iWU6akpJZQ77yk5b9cphRrMpTy3iSvyQoAGdrXVeyi8CXtQs5Ijbfuq
RTwRyYFxxddx6Rpz71H+CBPLt9njjTK8ruNzUyBaCAy/X/2FlU/dLRbo5mQRG9Y+zIF0a3mnK4sp
ko7LtVAs9qodU2NGNi7xCdgQ9QBPbRDPw5MPHMs2OmtlV3AqOa8IdMka/PfRxVHxZQlgC6yLOPM4
o22iOXkY9Ww/8q05g2/6kylypPRumUTvSK6THkRsPFotXPAInaOHcvh2XUiyeDfZbxfy7u8u2V7X
6AQmaYBvc9zpZ1Pw22FlERfSPCFv9n3p8GzoFaf9hJRdcW5E9h4lbyzSXxHBdncwZcud71xxk4iV
/rascVqPHa018Rcr3NB6aBB5YX4eMoDJ0QFUBR8Hh0oWyxt7Q67RdTvJUlHek+LTdejnufyYjq8y
5vlvcYXBJ4lVwcMaOKubq8Brvf01zQwntx/Jy/fX/SKgjBuqIWC9/KWElXoUh4Q4zLYX5kJ3IWcP
tXCTegwCWalvrmsGVTzL4V8OyLCkOaLvMje9YbdBdCwG1Z8/suoXUU3R4Et1RSMVpqQ/dNXesjm/
sqLn+08ofUAa5iwlH31PSgoGq5HBN40fiXjae8qAXMs+7vOGVlxa94v3o36fsnZIb4d3ufrNBP4H
TcTSL8rUfnOtGNMdQcri6hAR70yUw05X2EtgXVxtIrUG2DbATeWr0L9F2KCJPa7vzO57UMhNyvKP
TXNFjS2XkBDamYYEY8t0dStb1QQmQD+L9Robi56OODqU7gcsfCOnxXrDt4gcPCyXEaCi197DhbzL
f/UAp+WYgf8AvAEFbxt/vsTLVO/WLFj87MFx02eYXwBpmSwrj3/CDF+uH32X1HI9eBkLHfmkSsNt
UlgwDfXiWvu1EVKL2EvMwI3mnpMIunOpO9eSYpGfiHxGutZn1HTk02orxq9Jz/eBmPMmnu0OoWH8
kX7SthtsD6a5SrqiXEDi+s8UWFjYXyvy1KfOvzbdNryr9FSz8TT0+Gtd8MyXz91aBmVzunlgNn7X
uPNRHahUBqBOIAz5OBoMgmC0ytCyu1AuwD3K4hQW3DuDfnqfifTamTPmdQlkvf+PK9+yfD8PjMiv
IvrSw+FaE3d/8frvI3crXXzbrkweH/Mme64Mep3dA5c2cWvRJ+qkUzYGFunGhwBJRJ2Y879ClJeA
rzz5QwXST4Q0aT1OtISK4bW48gq0hBGX7n6TLm2an/J4Rnp31VdMO8dsFKkHONJrBo3vGKNwlj+V
ccuUSNDPQi9UEqz4DDMn89N7dVgyoxZVxqJzrRqww9Iwsbe4OauMECx6SE42Rs51+DexNo3JGPUL
Za/DBNncwH7U/VYhHQ7HRJ20mQK6e8XDwuz353nPVue2yeo3tEjSuY+roD4Z8hgR4+bcB16OEmrF
BSOnHKwAikLD5jd+o58AI8zQ8nO97x62dcrU/swQTqZC15T+Uryk3o8qC/Zn16v52YP8B98U0AIo
AjZVdoAKRuWJDPvztVeh9WG7hNFg3na35bIYaZwXNQxRacQoEj13UXtRJsrEnKvXBRNntWzClu6c
BN2/cG90trqZDNCNPeXpFFqe6Sbh2+0pcG9h9YuY5MSj72ucOg2FvcsF261r2J58Y86mLD9p8//1
iIJpeM28UMRqN17CYPBomV6wzTDhCqoL06M695uX7Q/Fp6eFnrk+2DV0wvmG63nCvJ97CPxZP2Fq
RfRGUCPZ/pfw7BGy/Yst2vVLfAhLCVizFLfqYFL9IDikKlBbmGJKaM4KdjAemOGqaFleSo6GCUjF
M5gYJbjFbb7sSSFZbHy5eqaKZNunjdO0y4U4TH6WAaPq3twL5C8bp8YdiEWKxJAZQ1kxeb/IgmL4
3kvyvWxrhsVmnEQhCbyh44gG5BS4qCFg2EpqHhdsRqKiPbT9Sh9KFsVO2q9CW3WHV1jqCby45Y2l
ZC90ycrQaQ7CLilHLWP45u+kpWoJhXY9vMT2Ee1Polj5yJqJAYRoAAkE7qFujmeYsy+F68X0Va50
qBZPNVKg4djc4j6oKTHZHB8sw0tKGBewFyXIxgwphQux4ZLZik2s2zpteI80vXY7IvsHOySwMgng
fuRAzSP3kHNpebanPVbmtISAYezIIU+qGTWSkUHNCi/rmitHS2QJivRddWDQFzQAwhWL0rxVnAqY
mWBrgHnVHZOe66R5NPDzK9nvniTn+u1N4ItE+DGzza3/uWqdkoQMrPhcSMDnsViaPhsIYwpeFGQ3
WEqddlCMtshfnO+TH2B7cFNwDZWPSN6IHyOfJJ0kdn9jWyd+jrFsEBmYENMKMF1NBiDW0hjORzsu
Zgcj4jZMnUEJ3nP1KY+1hHtIj0LaPnqbfUltL5fiVtaD4B4XVf8o4hmvc8VNGFzFqBJvIlUMvPXH
4eTLl0hd048ApMTCyOkIITg8GjD7WgcMJgrPJUFc/kHurKH9lM7HtHy8P75zDJg6iENMSAmIrMOa
c1ovShChqqCjkQMMvRZ0Jx213OSzoEcr6CWGzJyiK6hoTCrl2AjgmUHXerkau0E//tlGLBSFjku7
ccCaIKswwEC0LxRWOspik0ogc1HGgOOur291CrboHD0E7MWlvBlPl0ImaAIPEeBwFM5+DQ8avUZA
+Xr5qjdRzOSNSzpsdewNosdkAjEOc22EeN14fn15gttAFWaCOLKjGdkLx74hId/RwJUkIcWyJDD7
ZiPFZjeHXN3dUF7LimrkCzthBBfiyi8SZo2bw8A22BfyASuxuNR6Fgi7Gk9Tzd+PMSdgyW2lML9K
O7THvDJujZkx7ZWm8LrBsurSKo3Q9LrOaXspWqRDQ8KRl2wRYYT/luuAK3Po7r20A2fk/oYlrOd5
rXKWrsIyCD+iTloo+TKxEZubrpC1qyVxyBrmLliTU0v+kKWrpdYWyFi3vik9C/j4MHFMB6OThvSg
pruKaaC6GBQiTXgQaTl2ytuSgGruT4jMCR0fG4m+XP05XZe7bJ/dNZoW+0G5sRWLPcuLSpIgXWZA
hmefgm3V4wYGhaJpuWLV4p598wNF6LFw1GPAzR3MucL3J5IdEQK5xH4oe3cimeJDG5bIXl3YuV/j
jlv/Eqg/XyKVEUQ2/iWh1U9yzBJ7DuUt+4AePvCZg7iiV+kscmm5KzWoBJpLKOubTTnxEgC+fNIe
9PNeMx0RFHpXizNzALuwEaqSsM/mfguVTJtp47MH7//C6OcTq7UrVjqakBL7nthmfCKvhB0AYTYQ
GR056d0/Wk+11ZMvu6zEdvGf+lIEAT2yXiPSPvV0sHv4GjbnjB6fploURHRpPchTvUl2EsxazB/R
jeRqVaAour/y6smfPYkXMCP3LBoSGAo9kjyYjmSBEArlQaf1Pu8+y9NaBpsaAxodFM3F3YRdC81w
Wu2fFfWVHc2828YB9tYEZHPJQv1duMYbHKKZ0X52tO+6g0ISQ5mSB4KHN+lyeLUXxu1WXB/gXO+i
QSLb5WV0oJ5UNZYEfgxKts/NSKw3rMS/9R66RpXiOER4omaKPiz1YT/XwqOt1J8YUE1W2jS25rVl
83N7UncaTcO20P/3Ohkpd2gtvGj9G47ArFu4WmXgpMkgjGsaQAfxqpH/UVxoiytfJ8w+vxxx3vFy
g2dgg/G/Y5piSHjMfKODGeP7qZVD+f+Kw6gMFGzM2aFKC6x+e3B2wyE/O6bSj61WjnKH2MbJCLge
Zl23mKn5iBT7MduAFvLi3QBKG3JAjFYeE56cZdBLoiko0cSXLughvgVr0ZPLxhVCu8wKTRLCoIzi
wKB6Komnq21nJogQWx5LPkmWkdVc0YB9CsueWO2YiTEMdytRREmtGtpxGYkdB5FKwj0e8nn7pT7R
jUYfL/LM5r2s4w2w0oThZjuCu10uV1zFUGfJZi29C9jhV0VW1E43OF8q7ZuruZYf7A3TKOB6hNYe
NGZlt5/xVf/Z4b10qMRsk0osPuq186nVeK1SqfZTZnI6u7rjbV83JLFYk+UsiAUKlZcDlRB3L8Tj
NVSS+zN2zNFLEa3/WVgKSjPp1l4S9IgmR5/RrR1hC0WxAKV2VTmxgshd+2jEhCVVCQTg2PHKAyMj
eceVHZtKPDZVlq1OQ+0gVy0TuIt0OLTcakPogenPb9Eg5DivM9/ck5RqsYG+ckyV9rW36UJZgDI8
1WgynYK3QiW6E6Dh2ThBkex+P9JXmu3mUIJiLyBGAiS4R+k7NFlvyXq2lJy2cCXOBR97sp/zGX0N
+ZPJwFJjKHoGVpCrLxxfAss9OinIvFx6wl1uh5EbgKPUgvwIjxjU1OTCfQ0IG8yfWUh7RcYfrSDv
7x4mGlcrgFg60P7YBq887TsFjaIXuXI+DyeiS+tiY0vuxqlQFoh+63qJo3198rEMeNcLv2pJYmCw
Jk8EMU9sJKuF/XT9Hunh8//j4/VxPJeb6tgILaGfjAGTtoCTT1kVPOr5mTgrs4ZSBSjZM20EvERV
y6izW4Hr1bJC5n0y7B/YAJnj9N6015oVAIlxw09bpYVYeBQpHmj0Wj27YIazuZZ79850nci0v0Ce
q3eV+N3/KEsytPt8gM0J9ZvvoUkG4kX92VYhbDRy4YVPkemUAzjU8mqTrm7Tt3etZYEChjX6Ej6g
mXCJC2iyK935PehvuEU6qybppflfz8vGZ2+snHJ301l7r3YtuuwFIpfNUCVNUmgyk+4JMUcdW6x3
xCAJmzABmQEk8q0I0iGL7m4vHChDPrFh44HWpP5jmgeZlnX1DjnuIX07mSv9s3ultsI6JNv0C38P
TDZ/AY4UfXNOOjHKiyVayGGIPoA5hXBhTa9G5Hd0KGie+LZSQPaSi/ZBF0gPHImm2a1/aeP/KwcY
sp8mxJdb1g6EsFHPfGsBQepaU5E6tXO+RtKMtYJzJqiqrMyTiYVZS8PwgSAIO1Vd37C2iCJ4uUIj
fDuEYleDEraZF87EHHA4ILMlnc422GeXyDcYBoOkc9l2oeNYjyqOndhvoSAakFYzGWPbOGF94qSO
8ClyVRHgYwUeZZSD/c4XCnzTjfJNtFQz3VYUpw2+eq3FPnnsdsCbhWgg3+xqZI8k3GaOb35XGZSE
pIipPd0kRd6Qpv/+WGf9IFT/2lIEUeE18WcwwjEi+0ynfhuTrWltLf7KD3dG+VlmXxHSJcyZq4F5
CGJX4SSk2gaQsFnlfleD2dpbIXGU66DrLF2dagzZ1hT5i9OrjPUoMvSN057k/6A/PGJOSTGOe1yS
SkIUJRrgkUiR42Dvg7LiqphlNilSNYlap1OCtZLllpC7FrywGWLwCIxNM6LwxQhVaeNVkkSbHTsJ
F3NoS1M3bKpE3T3/aHV2tNuIlwebaZpO/Ou2fHw8teyFKU9g1y9FJEBsjx9dc1IGyiJd6zood98i
Jq4tnuY90ZfpEXb2gGyydSOsRZLq7E0hm5XrnU4RbQ3l/KG5lj+l3oHhPYHOYNeD3g52IPTHNoQn
nIgmk4luIAoHDigY76Jx10biCpuaxWLwKce81SDpSxMrManbJ0eBdzrUx0ibPBjszDl7pJOmrsB0
CgJR0IpxtTQiLcvMHH9kdIRKKNkJEQchejTEU6Vu+Dvl7SBlyJIVWlUSn70LbRvzyH05JRG1OPAQ
qSIA62DhrYnFJpoVzzkeZJNtntcoFeiZP5Hwwp8kr8lk72AyVvGB+ijp2YVoOD9M+akkfPKATGjx
0juPx7VOKhUNyinD/LsfEmFr0ZNzqcyN0Q5dvHWV0ejXyhpC6uOncbk6yBCK/EYVtQQaQi+xn9Cc
pYpBnXLvaUehwYxoIRnVx3szYUmy+a4wtgC5N7WkSh6R4trPRCj3OhOU9UmUuJ8w3/dtsh9dB30R
eXtkvOcNtjKDkLxuhhjoSk+lxy0EEereuCJSKbFADnD84W8QDDPfCyyN48yMtuX8JwFu7Cou4Wmv
sMdR1e47YkT8pSReP7D7KFnxnK8ni5a74FLvDHXa11jcbdBaCClDIytJHU97GjUqt3CzLutI6+N2
fpjNkmkl8Qryba42APcBDC1jNMOzIz+3BnzHZpBDNhfoqI/V2V+aaf3iDhCQ2NG7Lg5sGiLZ7U9Z
NyC7Fp3UKK+/sH9dDlfFaua7cbOVa1LFoo73R0J9hRwHtRpVVOLFHpDdJKJGoQdTF4MOzlMv5ygl
yk2GqUmUH413y/lZ5FKDTzA49cgzYv8WSsVb2kHZRXQ+EdJ9Rc6UsNbLYhMU018/q2ekYt4kOZnk
3zWG6ESw8PxDpc59HXKXftW1udfkX50v9lDw6vT2ZeFk0COnKNQ35mX5gQ5/oFJhayEKBsa2slIs
kLxIZPd0p9v3Q9siplPCGgbKVzwtpyvZ7ZSFoOmapN0jArs4UyS+x1zK1Vx1HFrmTMnFXNZDAsOu
u4/d/I5Q4ZntP8uGk01XTr71R+Mkl+QTN2fD/65cUHOUhiy56RyrfZZ7nZXe3ufxhu3TZictJQnG
tdxk9fYPSqgt5if5kJG/RQA/WIXCNo+y58OkI6jilWA3/P19Yk8gFLzMBwP951NAGHOJPvD5HGqw
Q4SKKjYW7w9sxtq0u/C5aR0v7YOUf5NMrJOYE1/bSkaw0bPm7iPSa6S4+sRckT0yKmlSyZik4uE6
CD/RXYxYpBaa93A9UKosQbAyT1sYbUguGf1TYaM7YwpNnkqZ6snyrLLQHKg4OmGV9ig7QpvKZUt9
z4jgwCd1VVYZ8QAyjqcjF9bBAzzR5LkJzzAEwMK/iv4+CUOr9TCpzFyllBgleBrhVS5wfmSuy6HB
D3EHrXVyTENSSHK7mHk2Itj1a+21B5uKYk4uqIG4YRGjGJhRBayJtq2jFfSBmRSK5zOjWlnEjnCz
yuaSRuV81Di3eaKUWrjkVGuThzSBWHjKlxa5dgnWvF7tIER5tSgV/UnF7V1N+jxXtfWHIUOsoG7X
8B477QNGkuPzT0SxUSzuJyY1V+FjNGxDZpW86e2QTho+mzhz+TXNAexUodrWa4JHxgv0ChVK4Tvc
yoU6ABsQf6GsLO3zWUNsUldNch8FHEuDbxieHWAI+0i1stwn+sJkmHUB21mdBx1Zh+y8uuwpUOEX
ELiuK9n3kJy2PQ830GO0oNhDpwqe6nTH+pdfzSeH95z7YIKJQ0f7b3Ffa25+fqovJ/eDm88SNyKQ
QVuEFPPndXlwfanLcnCEOiynKE+WIVIN/74oT3zv4mr9BSoKiiwSTEjxit9hABuhL3VHWoGIjd9i
9Xf9/8aFj7PXFAXMTVrt4F/NqRptRyc/g3coR61NsSNBUaDKwlHelczXNiN0sh8lf9lEgyFEsy06
Opij+Zxzz0+1Qil/I+z2wK4hy6MPMzBxWUPB5xG4BeG6pv9wZuofcFqynYjlWC43Wd7DzOX/2WzV
By/z4LYelp6i1H8cuzJgUu27ueDhPiGJLHRj32X31j0JE6gTenPSGCkzDQ5KPmRWRaXOcNE7KcX6
uDOs7AewO0nKfQ+/F2C+yV8b+JKtHo0ZqwokEZ/NE8ybBGGOOMSjJLUVj1hka04/LFdk/8uV61Pl
r1YXTpxF0cGf/rTExvE4dDcTGmwFHaJarHiy9ZJ7GN5ef/JjF6P5P+jC9uo85xp5lmx6+CiHhpdp
9JfLYbD+wlb+/Af8jI5kU/nbUN4Yrir1goFfuOlwWwQ5199d86QU+IByrQlv6XqXxzQe22mptE0U
Z2Izmze48J2WIOtTKOq6rJYQprbx6rU5YbvBuLhdo6A7pUhaoFyrG2wH/AwBSeY9+SDtfozI5/Rh
HIPssGo1S0X6hzJYVuK3kDYXcv6xKETGcIQ3Q28khR5suvYU92OX14ck7s7dfmJUvbQpvKASPiHA
wEz6rnbdOVhg6uR7Cq0x38XbZpUyZTR3s4SMDIzXLukNrqpswY3vf8mR9zc52ndGDM1SzgsCwwKZ
VxfHrFlKde5gZZZf075xbIlsfQT6OPwk9xACkMqCZqpUNyBfveQUi/yr4rIb1SBhno6WOOBRnP9X
ExzInwO/el05AaWp4ow5+BjETWc0r0PB7CVp8uPEwWXE1ulLZuP4ZVL2MCQxOEHethliI4j2VeR+
okSP4t0VpYPsGmv/DGA1rcI2vW4I0DMPlT/cq8t/gVGbMufO5s4pInBS3dZTRGdSuamWdBmWlqzt
coA52jdvNlxePKusX8wd0j4lKqrNobfYQ9eAIJ9x76n/lwhiP5hlCpSYJElhhDLWyVal+hbEQvaq
+e2Ii4lQzrF934QgBV1EQ/gVdUrjlN16zcxUX7tizukC+XN1mtlmxgQRzErRCTaYku2AzKYBftFP
5Y/w4glKRXJ8xkkjOFL1JskYSBETrWCI3Aa8A8dzxoLa6/fmNIQTSMU7xVcU8fyIVX+HcmwsPN3l
SX064IWJc8SXtrJEFtdwcy51w1Xr3+vrW8Q7yzvgi0iXeaw7gwuCy+gyaxEO80+CBIpUuj/5ubzH
IlvzE7xmTlD2/+cCVFFN5QCNv2oBJdhaW0Z4a/uFoGnvHq9gDEm0K8gq4A6CMEaz7j+3J+35I6AL
PMtteW0unADejeSoB4mD2d+DgBDUZHGVi+HIMC/W4vP9ld3sjdlvufLVNumda2VyRtsE2fOTJ/e6
7ZR2IDZ36AR1rmKCaoZ5mIuvgZaWnofH6INTdiGaqMpMCihN3UBWHmF9lPweAUhDARD9nq1np23J
a0SoDv+7+CACPIdi7TbXAq2AchqSNCIXYGaNNvJgTgvp7bqsu9JakMmke/wpLR+u3/l9HzavMRMr
wPqHHhYWE5ahf5qB3QRaknrEHztSBYn0IxUDwYXCZuUcxdf5EeuWvrqSg6oI1MM5urvI1llF8p4w
euhnVqM/WqT+V9Uz+q4WUHFF6BlwuoFA/1oeg4crlf0V2Ki/g/Y/0zikWUOQaHbB9f0VUAjO/p/X
d1nVtfFHqZIiR27fIC3OGgi97tcd8pATK36zsuZhy89X9K4rUfKU80MM8NzQtlDtU0T30i4w9wyz
Iu/NRnd4emlMO9MQ3kOfNsLTc2iwrnuphucDrfBCp1NS+wDoUxMvOlzCgNaKelxNsuTlnPC90oO3
DI24MMx2S3hRIn5NStGd7ByeYACV1HfJFzLu+duTGKALiAAv8rJTX52J54NVLYc0j5ydXV519iDN
xza3W/arkl9OMWVHMVTTmryZRV7c0/wDKUh+BKYX5htgbg1c0S+3mGnQPlNPdU7HT3vFp55SyB8+
F5iuZCQmCMVakte444oEIOhjos9XgB4eOidx2p2aGlvo2ufizZ2cIsgFmvezpaBPV5Q+PATkqcvl
d4+WSMwJ+s/SLl7FP+HwWQddfItGdq/2o0CCE5ycOUdyv33R6nJpWuutT0hq8EicWL0qwFsCumQh
6KFck5C4+Jb7ahZW2hFJ46pisDuwEC23QHChf51+v41v/HJh/ZOZeU2qv9FpPUoy3i4MzWtb6oZq
TXlLxoLj73UB/iGtH+alz+I+VQ1/vUcxFJJ7+ev33S2VNps6uVqGL7xslzGDPfEBN5DMkVb1XxTi
6p9UA7WvhaEM4E3rr/3+2arNLKu9IXzKPHtlb53bMVkzZhouuzGRVpuWRFHq6Ps9RKTwYwo2FO8O
Kx3xvW4T+koo4uQLilSzkeGrnMiDn0o67t4b1kPJBrrAXQNvrSPOUHtr40VnN4/U69aJzlHQy48O
PR/HTZR7K90csSotpvf6TMb4LivaQSDQ/nhbTPXBBowx8u4qR218qiUUkEPngMcOw4PPKPwpl9OK
iStBiYkHbW96uSKQ6fZ5eeIOXTkNa/33sWQYzV7BZpCC4/4WMsyUSYlXhrcAoU+9ahymKrbbuscL
rVgMft25vIgFbrr0ViLGqcJUeEd7P1rPy2xjx+qjqGvCWRqcZR6zD385hGdbQ4TMOCzK3XJKMAua
e8mvFkYqQwzaE+zuMO9VUi3ujOidrEFANc2jGctaiaYeb9iqCuYRPnygw4gFxsNvYF+Sfl5aG9L9
WYESEbNRVOjKePKo6QhKp5ZkWripcAY1S118IZC15Nk4pkVax7PwWoFsAs6LlmWc3RHf3P0Y9yJu
LbvmhupYcR8ojti7rJ6K1ehmvVDq0MBEhl4y1mc9pNmccpg0f/lJuRuro1l/H8rzCq1vHEeX/RYM
dkrjcU3W7Ssc0J6MOXv1Upub8bUNK+KK+82KFSDAK4a/v01Aiz4cGLa9J6v9QNS2bzWQ6M1slJ+2
I4izM7CBwyImNTMOHIlWS76WVwJnPe1itnAKAq7fPJnW8JxTfua53CpfpEMKSPdBTnWWGF/nZOwS
MsniV9IjIDIP3SR4GF3YEYBdoT2Coy1LyVyuAepsH70H2jif7VBmxwNF3rhKOgatUjaTi98Xo5ck
RCXDneukHLn62x3asKSmREttJafEI2sIlhH06+BVSZGYO1bHU0WY+QnqFiDnucLmVEU9THbpRHsT
hgUTX1a78riNXabncQKq06o9RKZsDypoGM0uyWH+FVt7skRyC3+KJJ+CV7wgFhXNLnyGc9dwgvr1
IdagM1RYxOe3D+/M3ZvMB5QGUTlovA85SaIlp6ZEoCzAvg4WhCwHYszSFGSFrw0VE0vLdWAvYP2M
MyT3DVdqCnb0ohofj7ztMpkonu82AsV9z2PbAuXI7tWLePOTYaTWD+yce+vq/VNot+bHUT5kCkbx
7JCgUcatiL4LsBS6wn1L3IPf3iJiC8JVcdtWxZHSB1h/oCyPJ5B/Pzl9Lk5CNsaQzu09XNxoh87Z
C8A2pflnKz9/ADi+FlV4WDx9tY+V/U8CQ9GQ83kxt1tMr6zqCfS+kaN3twP69YPz/TCzN8ckJVOR
/pynB/u3CjEwHwOxkTZcglCybpEsvmEJmeszahEdtd2Coo7bhvDytOyeEnDG/r3pNzmZFg6b+tCe
dqjeF6ot/TMSoTElBueavdnuAHQGZxTlZYmQM32mjlVC2t+VW7s+bh0Mjd4ieQrAgm5MlcfUdncw
lDiMhFj4KPkcHJ+OZJjv4eG6FZJ5BYqV2GoP0BPjU/eYrXf/wvzQKEJzuqG8ZjYVADQIfSQNhs+c
QoJ6mx0he24bHTXdn9xkH34erFE9Y8dD8yAruo27UIkz7FHvTCq4C54H/u0mHL4x+2RTTy3+KcKv
C5j5rGhKQAonVBeHo9S9b197T7lFuh2D3eKFInFeuIUNHy1X4t0xU2fXQDhv0gPOfkHqChDz0hdc
RqzMdOmYo4oaHq/igw/MoC8rilnndtBrVjBnG/UQ+Z4Ke2FBfjfJAyQ7Slbwdk7Cq161R4bhrEDQ
xs8D/raOTCC7ddpotn5Tb+da9PFhz6Y2Y9ZaHRdRn0RhxTDSYI8Q5+FMjPmNp0CE+91PTN60IBUI
31PUDh71kLeO9bzIbVz82/JQolG707X/wxfciLGuyOtwSMXMW/etphwh98uHk0asTf4QFx/z/8bC
UpMb4Jk3PBMrHKzi4YMT/DogggoLVpiWiKYJDJCcM0ldPVpSs0CaBBSfCThvZ/LWgQqN9uHcfDBL
K/2AMQWR8VrdbPuy/BlwTb40yAlcGgoxXRQ1ZJPqHhDDfwojZs3kd1lc5xXhWcKTvBf5JCXLcyXZ
3cKJAMpzR3rJ04455/cWrEkyvOj0BhCWr2ChW1e3aEiaD/o+kVRDeg49KX6o7CSRr06RkGr9Ved2
bWDNWAIX8LY2zZZN5xGy8CSNRaeqwlU9EnMQdsa+b7hbZ4q7DMxnVtkumXaoRQhO0zCc8o8EuM4z
BgMKJ1yEt/cfwMdRi1tLI/82Xd/3MLrS1eSMJjAh5w2Ck5WIErad9gModBOEEkCEm6wyHhIqBGRO
Gwapofp6Wg1ghlgfjqYTH/Zf61z2DG4yx1+64T4tjfrMfX4Ml49Ra7tbrjR0mf1aRgaCwSLEVI2Z
QuTcK3dMrMdurfc8dF5Bi99CkSkHhBPC6aQ117lLveHXqWYt8AZu1iiUsGptVAguHALeioVg6tPd
/Rrs8IUF7hJIZSSvdS0y+2uO6r0PHKG4H+twD1/u6MrCmjpNFBC02jsUEP4dyfpVlVQ6KnW4oLtU
eyhgXrF5IeG7FdGDWHWwg3NMXdx1C5k3o0Y7qv/xbTvPuBC3O2i6/wgybrY9JSZkL+QBHfOkBQKO
/dA/+TroVhiC/G5I4WE9oZjEOwSm2R0H8e0yBO9Ih7aD+OL6Tx8I02iblRUQvZaeoFMZPMmCUdfb
xL0pcg+wtqoUqqOdFAYLsxg7yJ4FMrl1TWhNFicBWEHjWN87Z/8uCc+E3bUFCNE2cVGTuqiUg66+
kh7bD62elx58lT/kufNK9XXQGbMROLkA1xi/IF+LgvV2lSt4jFORvcmAyCck3yicIbIj5LLe7VaB
ZTxhx0eOpaRsyXuqcExiVnT2ukpZFGNp1UX6Qu38zWkAhtJEvPtRnEsks6wkOXDROU0LjZpSihCN
Dh1gxAA/I5yqYkXMU+VZUXJfxNnmfAey0vW7oSWKsoUXqm+rSMksa4vefGmwhNt/x4tdvbBp9yGE
rFaZFo4mdS5Uzld4kCegBGoIo8WfmEWnbbYblk6kJW3sWc50p/QFm9usuWIVtCe4HHoLbXqZvuog
MKMLtA97/25GIIk10MtJb+DUqogmCpk2mN5K0I0sgChXFtkG2DK+kEGfB7XUlcqUuPzPV6loW78S
eOVbxwHlSaNF1s2OQXkkIpZThZyaWvaJ5IAssX+w/CdlIG9pk/KT/A4sdblKppXsoq9/xSjDD+E0
kEsTT/lNcSOGHXEFtHWE7EZ0Bp3cItTiGdNYAF0r2QoQaNvCYv6777KK3DdjDWBn3wFgKkQhXYRB
Ddsvn1bn/8qmHHEmmND+huyuvDMkDfN3bVxhbLdgZ12xDY6ZxMkZ4ZJCmd8pGXygAAGtkkmLkNMC
uwfTGZmOGHBZPFLBKo9E0bfmDNprMQHsTp2yQAtf8O4/QkXbK+yXVVQ8ap9xmjSPHdzYAgBIMOyI
BhfZzbVcmcJXWnwTWC1uVtCsoN/rOlGtqR2yKDgAb1/iaFKuu0WKiSA6FJAMstT4BuLRYv6mgaq3
OukVrj04Uhs3Zsp2O/d2340gSdiSMUfGHW9DY4iWvwy59Rog06yV4sFE60ap7KVAPjs0KiB+r7P8
egQTMWAO3v71XJbieGwGgVTYmRyuGFevLGI1Ng0BX7nl7zcIJNRmrRuwZt68uzzzjItwr6yC52BJ
0pAGxk4sxMwtO7zllqy+jWsNGV/2eON4BgdCVHvQ2sAD8fNL0EZidAvaBoaxA5TVDxZky8cQF/2x
RnTp523dfPxiO98D/By+SFyrp7UL0KSnfTvDCTtSrqJXr0OQmBXF0cxzw4BnyuPbrMEaYc2RBlXf
lV+VQIMoMmbswvelzcWROyVWx7EryQvTPkXuNSt21qHS3fWOpDlfmXWSf3JWxZyhzXSl/RgQOP1l
PqAZQRgOUN5mdwNmQUvxffELWLRVueKQtR3sk23Mom2ODPiNShrQIsdDLmj65s75EM6bgybWctKg
kcOXcDQ324TlUu0DovgiY4jpnqYUtk+OQVWdubeqItNBURTaLOvT+7DvurgMC4l2FN9pDJ0Q+8rq
nR1+A/t+Cevfmyuph91LOn0xWOw46K/LSKMt79K6rK14uZeIM4FHy5ABGTGCJyv6xUCrIpafSy4k
xp07Zr/tet3QmJi7FAbiSPOFe/wW6YRtoORYaAKVvgHVBMlLBfPFSfKpxcsUvp5S0Df5b5W63dGH
FWqrkIiG0GMD9rrsEr/e0OzbvV+CPR1DHwHYsnauxaGQroBy2NHT6zVEYAwXOB+tDBfLrNTbB4q8
kf+SNvD2qnxJWP7Qj+WvXVR+q60GzfhCQmBtD6wXqAMEamJX2Dlm9+TUmPr8Bk9xrSH2y58SqU8o
0LDVNox8qbtDQjmSeYTauY9CyQWkYQArU4KYu08wxOPLxe2WpNjEQ27ZRR1ARE0tEKpcWtHuwYPi
3QjEYuKYv48LbUFUNm99F+o49sfPOqILjYgkjS7zJ8zZbMQMLY8YCilkybwObi6W8Rq4wLMwD6Sm
1UCtgavdm6n3qUfynWdMl+KiY8RjiI0+rdusf0gCh27vXNOjitFJ98awKVwXhewfIHGA8i5i+jcV
ubYzZLi2tymPok5tT41Ah/huq2OuXEMMEvYBh5IKyQ+BxORh3R1m0nr78pmGlFBR59bwONiTsOXj
6xkSi0FFetwZHp9uQZotZmF1eHs848ifsBPdDECqZhU6DuMUad2Hwj6kv9tdWLKEm3ZRC0tmjO96
ApMXAyiyRDou1TDGFyCo6A867gDeEXd31KCNk67FGuK4VKoO8TE6kVFNJxIhVi+iOYoGrqd8YvCY
li9BuWDJRC4RE5yhHFBkPaqzM8QfcmPe3QbPbnPUe1HCGIY4PvJOktPmXuBLwjiT09uU8N2C9u8T
Zv62kjhNS2Va1mlOIUjRhUR4Znjud/UGzMx2BQ+PSCBJuHrthyIQ0iH0A6R9Y4VwhZc7okp4H6HX
vKpOfg76YEXoiVlUWbI0D0ZL7RI2o750wmyrY/0W28BPq8yGGERaLjM2X1D4ft75cb9cEFfBlu1h
RRmMRr9CJNB7ou3apCx5a8bHSuMv9HKeZZlb97YyyisygFPwAmmgY/l3e7dVUisqEr8tBmyhIG3y
SaMOyE917/txzyRYF7oLkHlL83anQk9ZQMSM9NaL+Sx8751DPh3BbbdX8uQjUwU1A+t4vZhENghC
f/rfNhDJgio5msDWTIimiU+17DhV3yijJvbuNcVtxRc4FfPQ5lnis12o8r7AnIxmlNW2aamMPdpJ
MOS55Fuxx52qjHashW2j3cQXRSj2/fscAn4JK62HoNsLxLdwjAvANE+zKfJQ95ltomro6ebMFGx9
mT9QThkrSoR6A+8bd+y+T89k33S4a7cJyy1SabVt5pht9bhXRCAGX458FHUmVIB8LaIgeOxqtSnP
CDBFc7wAfukVylBmv0gmH2PSVYvYV2Kz2vMyO17AHhGW4QUg82ZNum42LT4ajST07kaM6iAdi3d2
R8p0MqZYN0YMK1x/oJJ8i/ToWDGHJrpwMRNxIqeAYNt78HRKFL6NCiAhhG/fpocokVpotoX3nXgf
6RlPtwVNiMbUQ5IJBscZruIYZqtHm0udcNcV8UPrMwPajepVlMCEjB6d0VFubLQzTvW9KhyJzxZk
kuGOvNz04vQx9RW8bZONufLgWxZXU6dpG0Pu5FhfmWZYbMHBa1ThOenuJ6jyXYhc1wRIV+jLHF7n
BG9Vsu6X8vDFGpKagAzhABmGMYkoP+shyvYrDSIbDdagt4zU+w07OCl1/mh4d3mwzWk2fSnuLx7B
q/IMnXgRaCW78FFG8+IAT8uHkK9OKEpn9kgn899ZiVMTN9JZXOrJ3fHBehhAQ+5ZmGcDxeYUZNKr
TlXCogLmK0E1PDt/jCyTljVP67Z7Xf66GVNwV5d3HQ5P5WgLzwlZs7EjFM8hKofPN8vQ6iKaepHZ
eKH5PbBtDwTAmtHLEptbL/JDD92d48dRfPL1+VTla1yIz/UAJJ5vTwBBXWUDZeJYvKadY7JPR3wD
1BNszXbVFaAjQnW9A5ptvxtYVHMWHeH/CwutJpeL7CJzZCFe81mTMr87JKWKtGELp8amvKovnTY1
X728bblZ1Gd0Zm9qlPIY7kiV7YSdsBHq905vdQ88k0bhNOFrasjj+aDEFHmWwDhnSLilOkc0z/4f
Q6ZTmvpCwwDSBj3T9jrR4QYTBRN3Kh9ctYvpvHskFUpsI14U1tlYcb8Oys2q45vHVD4wHoFV5yLb
1HK72ZuQ4IB4lzmk3P4FSFD4ogL3hYRVt5FX0y8xbqrZ+Ib/2OWDgJIlx4NgkvY9Ajtb+qPwYfN7
x7UjqzRI91QxF2z/i79DslSbXUwsyXyG2KmxvDo4Du0FsbH+okzWqBMwxIf0ja4UJGWqHrLW6uBY
fzUx2IdbapwWkt3bYQtPIcazy4Xzq0S0oF6+9vAghuYFtvyRIjzYtr0FJNXh4dgNPkvtr5s+Rr+Z
XErSR3qB/4Orq/8hKWEGjY5Nwf2K99kN9wv+/fcRL3yYOhnS/tNQrkmMafkMC9x1+bbzpWEfspGS
guGt53CX1ey03Ujdjs1CTOK7rA/bODt+XuhR1pTT3pquRdOYvkjiTmdVFv8OkhQfPZD+UkDQ+r4P
NoXHyegRHPEqcknTbcNjJmLX595tTxwwuc0iq9CMbmJXjR57T85u8Q38ksYgkej+os54A7TB54FU
IW84S/BPgQaGYZNCGQ2a2L3lrLqlZcnR9q6FZmqXhYlATai/KGoUiKxRR3rcdSj7AqnDs1LdpHxU
GaJYyqL6vIXa6wIJTHsWDqsTV+oxKQ7Fa4J4/w/B9LaXMVHQESmY/Pypfv+/1iAVRrKJM83N+XS/
K9X5KLk357bPlTui4SEQxI9zc2wubStGWiys0QgH02uith/oYVkzwRxmvWnr2oke6g0G9ruevYcR
1fmabZswQHmbsEps9/91QcXDGd33wlFcLFJh2cK9S0xAtYhH1MbL+oKFBJfXON9Ho7u7FYMJiwrK
95eTlFOE5dkw9JpMiEeShHSo6Udh9diggEzJWLYpNBbeu6+hmAvWDm4klh9xh7pczed5URdw6Zql
dgxxhExZxEuwgZysP6J35TctTprgYsj3qmtED+aPaf1m7nNshgl58b2n9C++aj1A5DRTqrjBE7Nk
U0ap5LNk+TWXp4galtS7Gmkshu8+gWBTgBGUwTjUDYopjlKK+3Sl3WMpwdePmbskDDt+SZDUH62F
dJF6LZMDQ8RaoviuK2w4GaV1jzUHBaxsuLQg5znONcQdb6H46mcnY9uUZZqVR9YDy5dxmGwst5Za
McL83N6AwEA767o+kTOBZjai1sBbOIz+uE2ACFv+0xOu2ia85FfneVssMImdQmSzo153nkAiUfS/
fC7UA1lSLWLLnZgClLx0UyWSLyDpSAUglte9dL6YUHmCGlytfg/PnpsQtMiwO8WNLdjl9jwSRCeb
yicaZ7zBK2Z3pej4gx16EeLNtWAFO03Osd3EuSWIWyIOSOaPcnMM01uNh8hvRFb/SzqNQYlWlwQ8
zYf643M33KNXcGEySlVoRut7Jsd5EHvc6wWmB69ODWW8Edq6wqHrR8MStdOo7oSwrP9/qXqVVdPc
o4nvYcIpaK2dwPcnPOdLZBn7xvLdbWg9HUsmWqoJgphw8MqMrJJDiESWgwMI7+LCB+r2quXH1aYo
TmSaM8qdtj+ljOIBvar3QsyO78yD0y0nIuHyIZyOXXU8qrtUvJpYQOGvprwHMtZEvt7NfJap19B4
RA8KWPemd7Z4/qMXE5rPF6klH6fNgoAN41TcVoUmUl6MkadMeGphaLCqCuK90KznYi+JCx9kQi/y
dupVPHassMbYHTNXe1MV5QwPntmvt5XW4Chdf+7tcs0ov6LRlKemdBEnCKFpTI9RNYiafGNbTmeb
dIhvAR8w7GZV1x1yIjYxWhaZi1cS6PkOHo+h1bcFXEZl25qBJVrli5VIzOdtfFxJgmzQY9vybn6m
qsvVV/FIbSfEMTcUiYifFrKaMWhfXy+URIK0xD3sWYU+ePq30B7Zc/iLceaYdehAtn3Ki33fC0HI
iYxag0R2I3wb8kiuPswwwVLpIfMbtoXxgbYIbEZQ4DGjt+adK0+mg61GszpGJwm7tWA3GEXU3kMU
dbrBnIKdDOzb+qQ6RnGpWRBErMsbCIWZKDjl9kEa0c/m9WK8W8Keaz2r+z1k8o2AyrQOCw2unnWf
YYmuJlmcPWzhf6O/lYl9BUJC6LKYOV+W0NQiWj0DzcEYai5JHuCfIdEBqaaThc0wgBtktFmy4eyc
oAIKUEayD4NjmUOLe2wbZ54rYhCfFhp03Y27E5w51mRKOr1xVLbJH42lgd9vO83B8TgbsL/WE1X3
BMd8u2X93RAbB/GCJmaYYw6obK3hdDtQMSLfCXjeI2ZxwncMEIbKx37YrDf0T+yyt2EX1K/48pMe
Ub2S9SMxbboEYoiWlH/iGgzc19tOptlxME+zsCQZHmlmRHQQcyc3emTIzn515oZt/T/ayj66WytB
rZnyz/usOoW7aKONJd970VOvJ5OAd+BFh2dZvAx1NCP6oflE/j0n7F4KXvrTtFl3K7SEN5zpjXtL
6CwEiHvzUrfb9FCc5Ljf0CwWHk9txLDImzu17eKIls2Yba3GZJ9H+PlX5uOymvHBX2128ZP7Ctli
CPIEUSZEpuICGaPzeISITHAZNhdehO/vgcf6c9gSi0G3aQ2zYB3Vulu2fOoVueKKb10QOYN8oLXd
yXdVnxJcclpVrwGqLQgKZLkJ7J7itzsU6jkhIe8V3sYVvcn7lF6WxqA0D9gDR7oj9AtYAec5xr1X
d1QMLJA+YwkQcIevrM+bBy3sr/pk0MEBltNDkK9sM4t2rfM4q+xDVw4MMNUH15ZdtCoHMvBxFUKI
ftZ0wQTGVV7Tyx77zXcGXrJSArG2CXs1DB7Df/CaUT9a+SXka9A74bBtE4h//7DubynBYdpPx+wP
t4k/BySiKxgz184EjW2QZ7pif/Do4niKZQBYM8GBzVnceLv1evopQ0CEWRg6ObqIcjz+0kqA6Y10
Jpv9VNYT0oee2kdgS+6d6liIb58ihowOb+2qq+WDek+Pmp98PsMKZayJ3h/XUxyYYaWZvNOUggPG
oLVcnNUngLY/Zev1GvTVaxW9rV8KTwCZCuebR7NwY4k5k3W25PZFrnAccs5ot6ifwUCXdmfLY0Y/
TbZ5jaKHbxO2GDOsnlV2cjGHpeh9kUpR5u8ljZ7nmBS6IjcRnER8zU/IWcfB1SbCfTTLn9dUVZdU
eFy1hpR0ET1H6Af5b79tEYFysF+ckF1ivKjLHEcPMKNsdGKQRqvqTHU6f0y4V7+gtXsibmz6yZyI
BF41OuFYVkDBDohIYn5XrFmCVRILTIFHBike2opAR32O4xVpAXb+gxLrxFawehUeqfGwPMp+eOoI
KD61v6UDQl9b3JF2gVij/agd1CMNIex6hBP7IKNFwE2lV8xeW/KktuVOopb+3uRHDR6L8vr2wjwK
ct7H4HKZjISq8I8RDfKbS8DQRzUMLLaMdokUem+b8OWGJnOZ2XVqVLDjrR6ceI9+i9Lx+gN2wnXh
iyMJ9RP8aNezrT4RZulcKfEBki0zftoeFwwtO5+z1+FPsZ7HOR98iw8052uLUwmvznzPnelHPvjP
2akcpySz/pK1TP9b5BRYbkYhWqpK9mifZ/aLT9L+SpDpfmu8Uze0kvgWBmCKH3WaRTnejiaa9ZQX
pSV3kQ/kaq0iChzSRD//XP+W5JuFkNCifKdVsD+lmTugG7HQBkA/AoIcmVPqCy5MQt+m7KaVwJZt
ZnGiQj9tcm6WMykDSP0Nl72dyJeuq26aFSDIcb7WyMGEieOPhAZc1KW7MQzjrwMVtyLY3Dp9xdxP
e6crzK5gF9H58ZES/JzDwZBQs32+BfqM7o2rfQ3Ir9G5C18ZWn/FoHmIyosfIFihMc0S3KHcm4Io
5U4GhR/Xz/IOPkS4ZxZ9BTtO35iZtSy9J0bXj9RqMSSC++UOz8awVQ0chSv5vrZ5kdxxuA/nwv1e
OMCXyGWUTRhSDsnJMeQGxKyx5sGhgqR8sjSyy/CWAm4eUCA+XqRRau/jIEfHNebOQtYgqMIfGj++
Sd3wIWZIjJCx5+CM+Ht9JGgj93gsTa+vDx8vBIsiO4Fki7757qasZGTC2m9W4Ycbj05KyF6ukbQO
HTquM4Fe6RHkrcUSFXoqRsPKw/rjaedknqqyFHHVvW/Pd5RQ9rGXF5a6xYIvwkveQ//KbQld+1dF
hb97iteFo5blDAYoLP9sU7nTKBMKHNZczMjkYzP567fsqDnth7jkKfc7fT+DQxHXP6ZN7mVXy/+i
9AFsGqLV8mpZIqH4Xs0DgvFr3EUBjl8pCiBIF8crT5ggfNeuI6GbRSoKqCWGGRwaBsPQSiGk0qtj
mqAkf1h1rxusFGZ7sBD8EUCGlt8s2wiEdkrUCjmCrLiAjDW86PHtjtXRLNFQNHa9JIpBda211yfo
QXLadDKxxQpqG/QdrE5ZILu7ZHWVp24+Br+bMHu1mwpKYVKd+9ZdcT2F+5Cq4s4BUUW9u7AJZnT8
G3j3hfkj3Ihitk7A4AflWhFacc5L3QqWbfJhdhlSdkBj9B5CAiG/9i2mfSbl0DUghnxsoxfhExfz
tTtFOYz0Alb2p0/yyafLXwp9o/i879Kt9MVsT3tE8zk5HDxWpKnxS4g32azBUar7IT5st88Yhf8Q
n5cxG25aF7LlcNCMQWLBzYZ8MMw4Bi/P+NJ1CEp3Wo27sqpM04YIWRRsGIGblDQVhng4ZEUf/ItE
EIYreYPnlvJ56nx8iXFdwmwJFlZ1xqXqENfpU7jOCyvtdjYt5SqopwARBi9IObgrqDGPF1HAk1iq
9vss7MF9Qc2OQZs39k/quOJPn6tnQcpuV3F0jXO1ytlsV42EKang+/tzBZ+8acIXNi58naDJ4Sew
znjCaDImvmlVK5ZhqTpCGsMc3lqFmnl31WVuLA7mmcxDpM285Xv4W9vcWSx3Gr9qpezVebZ2tLcJ
BtAmeiUxP3hs1dW4GLpAp3f7sjVrZppHc9NfPD6UMjWy5igQvHCVDQZEpSTANPlDRpiM1AD5vjd3
6grczcpeiGeuD9eETmid441G0TQWz+ZQVh4GhwroHWqvKsT+40ZSJtz/g9gllApGHDh2Gm+vTOFP
75iAZKwKlPzfpYL2433SzAU0iyqtlR5u85zcbfrJEU/dYWp6QrkLOFTUPjTL5tGftZCM0rIwHt/U
2YYRVvXnjQEyIJqDbMgvvlHd6z6ENJsE1KlQujHUPr7uGXkCINJ1nLquxJ2D4/1ElCqnzXx/p2Nt
2dXZc4Vy7pElMYqF31t+Jkk8EplOMIVSEI4fysw6jjYyqT8fs8AJzcEEYlDhLn++FUE2CQcfG2xn
wjAxhWPXpYRaV9ooebMN4ekt22YpDunE2xbYW/s6y7LWb5cScs6DgPL3s3GKyxB0xUjQcsvBe2a/
f0VviyDX3LBeDBQAiMuIkV/3rZuxQE9HqxWnbnxtQtzDiYAgNxa1euJpY1Az/ij+eJQaRliV8MOp
9yqjyNq8Ybh/uIXpGs+VFX9TV39P8X/6a/zsTn167SBRmlwA28TRBTLXFdMchdbNlDsB5clkM+JV
BRWvAUkscnxI1UOGgbYHJ3bWEAfuJH3vkeVB1UDyCl7Xd26JXLxiGk1qTy0DqmEH2yy6dSFeuvcb
JGNhtiuwV34vX3kWMiMIReQhtSp+TgaI/aTSyA62YmYvzUyxcsOi92vvWtaTZBmeidXxMGoU6cI9
KXC3nWzWy3HBP1ZnbROQqfsrK/pLWSAc37rfhciA6VTKqEjmy+E2g93JuYHYYiY6qZ3omcee8f6r
77mcwS7un6VPJCIyMIw8CuO/+Qm+xQlAutx/V6eU9dz7QC4uOSM3iamjGJJFr6JElCs1tfcdlefO
2wOhRay15wEB0XA4j6rpbHYlI112LGHcY+pPabfxCVUk/JyFTH2f1j39uxrUl8GzofFyWukD3mWA
nCRwuXbw5JXXz2R3tjQeJT5du/j97c8gXIDw4eShspyQyn7sEr1D2PZT5SIj20c4Cp8Y45uFOckD
xP4hBlwiDUqgImpwNTYF06K+WSUoR7RYUCmLZkk4hiOqtPuKsokcfMSBicJRSvn1Ka2R/IBC0K/b
RhdsL4FAhmtVkW2e4jnjXNpNqqcLOpFiP3AYTueq1ghLYNUW0DOjU9brdzwGh4UoY6jsauPnPvcy
uWTg4bFeVph4AovCCRaCy3nuXDQcK/x23S6WbqoKVaHndmY9nsBXmT1347C46wRS7vEMpaMvCXyg
j5wMCOo7rIzyXF1/AObZ6KkHVxGHwryk9p/NThn0lQ1Qj0/dD7oEu4KbV6+3ndYTPwJBerWKxXGD
TSaVvT0H9ohbJns1gf94UNAyLOi0BxLUphVYskccN2hbOkbJdvxqvYZ9taDk8pyBYEP8MK6S5Kfh
nIVyZbufj9XKSpPTwU0Vl8sB/me4wiyDbIl7QBGfSqVGqU1eDiinY4MQHKNG9K6WobnjZ3YI99F6
ze87D8OQldvgU51q/CFgCQIsas0bsMR1QnmPDiUy2Ns6mddVSaP36tFES9zClRV4TE0YJtCzQvJy
NJtyAYCpU3tXXcirvan4keKUAefSWrewLx6flmlUcPvG7HB0erboONFg0F/wBRb3+dJ9CDn2rxJR
TTCGGC3he34jeQNgGN1UpZmCxmwwLidMFqPkjiTwkI+OUGw/rOT5R9889rOVM2sk8ykzYsImvzT/
YCRgpnJTFWhlNCUgeS8mPfWtMxWTk3IOVdyDyLl4zW3ICAqpHMqa88UIbZD+DTO61qt7TpYoDDTN
5SsxbIi7kmp95dsVnLpYlYC4WPAF+QT2HMD2A0FXwaSVPA4R36/AmbpG4+SSYkUQmrbUX71yGktZ
+Ety7Kupd+EzBWboO/oAyot3ZXkYnbBF8Uo8rHEsm0DnPuUc8pZEquzfX7H6GQrm7J1380PxPBW8
SYnFJg8L6Nn9gGv6sPlNEnj2Ov9phic6vSmlmIsSSaE8XgrqDSd1+m/D1ENM0sguU4L9WqDJBYBU
hpkyA0wxD+ctTwC4318JTlhKL0JXS45D9ABtjJAvSqPuf4aVpF1xWzY4sDIl/pUp5sdh+nP6n2Oz
KoUQmu9jKEof3q9EUyoVNtbkQSLwJXZGenLI00r4o0qLL7AwwMCfFZZhWyTtZIJgARJdAaGZgn2M
hxaUfyEjzVFlq/pYibaHObhNiy8iLBQbwqmFSTqic2eu2Eo6cMdWHREccrPL4desfSn8E8beBMuF
iWdCtzOe6znj7wip/RcrOIEFq9yoT6/6MQ0Y185Wm4MHZw1mXYmFcSlsu7wEOzIgfoW9g4zuHcF+
g/EpL1Cwz6KBEEFDLNQ0+eyEEgqmeY7zqwX8AxwKP8d4VJYoCgEuOh1owlJye9udWTwErudu1Qs6
bgukBrXSxIV+koWeWsb/0Dd9Sk7swnn6wnBBHliWZGiM86S9X3yL9vq5Di8IW4PHh0t+Tc59DFYY
KJ99EX2hawlG8hNj+UmyDXI7NW2g//IZ2HLfYYA+MP/PoL5QJwDRAXewH4opEshdQgvrUcZ55crj
9Jq+3thsIN5i5/DvXEYFbPp3wUkoY3lZcOzmEBuKVM8YQTZsgynV4yt4Ct5rwCwuVDR+5Yj9Tu7N
KGj5JTqUZ2zKy0wasW5YhkpziD7m1CBOnt0+xIZvAjFPWOCL2v8vhZ4Wo5h9SHoLn45n3zUFCsP/
VTLKEkOw6CunTu+GQsC42P7wuFlT+rpBzkB+OcZKPfwhGVOdvk//U2ePZ1BfzhqVNoVhuLeeqsTH
T4QnUe0a4bz2RTDlwUSwd6XOuAHs2+ihvLErjsY1GrryWKI7tt9j56WzMvVdy3i8tE6J71AtmkuA
mnJS+urIQ7d1ul4YCKBhErtsI9UN5k/c9p046DGa21LKFi5Qf3F480TRSJ7u2Ln3I5CCvkfD6Y3D
oJlueYvBWyZ5VjRsaAi5SFvEDQTMnczIk6I7OhfYPRoKDPFK1fbY86c7k8y0HKzcpDLhet+xi+P8
RUBmQNb76QEFG93akwmGfJBx9o16riWwCHv4g1ttUR3c/p8U7QLO3GdStTpiRj0hvZROcQRAZbLJ
rlxUKpMrjpQHQC9HMdu1h/kZS38vTWa9Gk0E4GrnKtUzSXu9pLwS7DiKox8bL0PJH2wj5R1XsleJ
eQwz8E0PHD+Q9mwsAK2AECUxO4194QeAeu5jm/NZk84TK2MW/v+XxjUN3q63eP8UaQyZuIA/ffX8
pENidkqhK7B6YAUOrk7gtvdpv+LryV3Dd1qV1jgJOXGvBOvKAcC744gY1MgmJmg1Wq7XiDItN8LT
GAOUBZI/UX8X3m+aItlNl/nL0sRZn3QPwBGPk7VlHkG56e9OgioqqQkEFqI84gK9B/8bWsBTCYRU
IyaAy+Se+5R3cndJhraYJi9nD6rHJJirl+1r1fc6YOpJ9S0mp4Ep/ZriFY3AlVM1rGrHUUUV2KRb
8F8PfoX0zPbgfkkk31tnV0I0CY81+e7SXOJIGEwNL7i9d9aGQVwt9mXbLHUqi/j8SdvPIf90+fR/
OlHf5Dfihp5RCvNuRUhsuEoY5gl1dFyTR0F7USuvIxkBqvSPN11jdTHKzIS9ZofsWkE4NS0ssdbD
JA4Qkg4a+NRyWOrZqQTbgBtyhQxdeiAH5ZqYt4ZzhRn8KoQyDM4eb9elXupObYOj7hn4s0V48NRH
DI5upXJzubPfGBhDCdqHHUzcZA0mEjvxM1hIEGWB75vf7z7Vl5gvz9eH//7opKdxXJ2i0g+SNq5J
r9XLwLsLBUIaP5x1HnKE0fSNxjOLlQTgIgjuUoRkWmg+r/hDgzO5vNVUagMAP8DYbeeRNuXLxWHk
tBapAGe15DuDCzbsBCwCl4n3HpCoApulQy1i8oXLdaRDiQbzpvBK3oI5PDb9GPIhSme5L3bao5NO
WaJJAzZGPTBeaskKOg/L4KeDSznbvm6C1jLtanyG4HG1PKd4tMTXclLQ7mEOpW6jFALzECDH6vpp
jEaIkci7TvKWh9QNA1bzNBamdW8CnCfLsju+9jKr4pzql1FhEM7+XSWiKAaSvONWcLAStTldw0rz
MGPenREBqf28yFdOyJmoCI2OZ9e+9KxAwhxCjoPzB7ctRLjSXcmywkFcLGz+nWs4xZVUcLOFz3rl
L2MX/eJJ7icvQYhIojDoXJzY1IhsgtN0Rg+VCUvRRDD/e7hTp6zCusCzOQ//HPXXhFgXhoGskyRW
PiNP51o1SIvQMDmR2yrKSj6VgEX265cjXf6TLKDzsx9Xd9CJniFRIL3+nvqIRYY9nAXsKoA5FJ4M
wm8gd2jM8TXYmw8ufOwvplArn8K+xDQwUUbwR41jfd1w+1PHos3QR6VcQnfbCBL9TZ1h+vhOS/Ti
FX0NQYwlRmJEcSWN2sgQX7kF9FTq91P7nhjtyONPBLXjuS19WUQcd92/V0p+nkWtqfSER3X0Qw/w
1va9d3ZIreltl+LEO7m6wj5cPQ32P4YquRuJnve7tZJNqONXjJU5YdPi0Ru2pJW3cvaJYGrTHGI0
0bA5KgOpbchA2gu6xkhGOB7EMx6nJSAhxvPZVDt1YWUuLZLLdSmpKWcsabCDjigmkfRDj4pzDLhm
GlQ59WpE/W65Yf+I8UVjPabEsT5ueUZYPtzY8eiNSRHp0l6Bklaig3QTL9zcbBt11AUmDQ61B3iu
71xcaBKrqQzvwewiVuzSyVx9pdmcRlYQFxRShFF6jU/58dt6zEXbxBFmaPLf+Rj9MN9PZeL3IxWT
2e82bK+Oh5/lrO66E17mazRwlj34m+ukPDVWbxvjlMCDP2T7bRQXryy7FGfpzsMSvVyVk7azvG3Y
zXHAb4Fsew03aBjItokHzBKlZnA53FpiLFrFqxXbNT669Lg9eOAPyfl8oB1mRLWuoR+gz+Bf0VL6
YUqy/RgRnoBVm60UdivGhgpRtqwCv6BHKK/3mYqBI42sGg73ZvhNpUw2bXTlrTLJGMv87mT/IkpK
MFcmNuvPxIpI53XK0LAEKK71AH7zoPbqz7A4Rn6LQq7IUv4/JjWQqGlVcF65rEMtqwJen5j8MFql
RftqRLaI9BiXZ9jJKXeD6+uEDlUvv+TkNU0iKc2e5i0j019BtxhZpCxk3bp41RCoxF0MjDhcDO/c
5oCsAWATgx84u0JZdwF5+XAa/1N/KHgr5RQxaD/sNURK1Yyg9dESZla6kQis2lrvBWBOeLdxw/9E
nI4iM6chRIfOVBZLxpUj1e2kjqob4YUwvyA8SD/hp4MoS2/12OAs1JTub0nuhyPISEzFDAjqyDwT
drZDjDpXRWU/1JZ+lyLInU+NUNxgorsCPVK1UHSLitUUgQh3xuM6bp2jkWHNNU0hM02em/FGO4lC
SMzc5CkgC4DGRn73I+VuChBKXOSwaUpKbI7DK0pvaN6++Ngh3ZyaS3/hk2A2A70aByZiwTB6NAFU
35EojZPRelysDuFY074Q+jO9w9E6zrW9kX6lTcCe+x2fiUsQajF3SGAImN4C8y8OXf0D+JCtLBzu
e2+PvY/LR9HdRVopKtgDpXgUhbclevs+JR4XIpTqYFWlnyDatiPkP+gleIan2PrGc1QgH1je9lxQ
14uPU2tt0/KdnpnVF7qOfT06OUIMPKvLrJ3vHmy219PqUrjL58x0WnpoPPK8xTInVuYq/LaK/ymu
lo3++vscAjLiD71LwoNUwPrDFW+DPJklNd2CNgeNc7XTyUBokayCmiKsF5/5EJpjCjtaQR/zs9Mx
3GlPwgC/OQ7K1UyoYfcWfMcilwwA8mJSOE8tRDIRvGAysdIJU6fIBSwCgOuJ3M6MOyX07khn/peT
u4Ipl/xZaca1LQadT22SKduY3uN7szxDi1EFeWO/lmATDQ5PYWILtavgVqL8gNvrl1du/mVAM6/+
sJTrtz6EYARx77fzcNT/vLflwb9mkflvmftkLYGCKC28occMNCty2Imhpqh31f/SiFTfy4hbOkSZ
O2o8zy3x5doGxq3fBPpXA/jYVWP+iUUHsdycWHHTMlJn7YMKHYGcJtEmf9pX9F4SHv7OEykHUV6W
Zjg1tpFwamFLUGV9eqNh0VZcUyOBvNcpOB8bP4r4RKJf9YunZJik2Gfkq34iPWsDdifz8P2T2gX7
o8FBUslW38F1b8qMr19/UlzGIXT/UR1kZBCQGq28MqxBTOvkPRQd96nv5qFd4nV+TQH2lerb1FRm
d4pTH15SYN0DMQBjbTnWMHRtigIWH4zIbCJGfOlg/5FRNj9mkwEdJnmLToiASMuLskUA8tnX4Kfx
dlBaozV2wUxuMgBMbDz+B4aTdepXhypDIEolCYPaFsR3Dxi8WMFtNK1oi6kBntLWsNCfLm/vYxXg
t7fQirf6KcvyRE01Sprlk5GzNsqG3ZWFSN/KCsDsYs2syuizsv3Fmq1wyMkaO5X/CgBPIeBTefl0
ust0pmNU2mTWYbgEp+MCfyDwMciEumSspmqhDFm8uWOvqP/2ZjyyTh/Bgq2Y+e8PONQHXha6gScK
oO6x1Bv4qN6p+MXkTbawzN/8XZbU47LfPRDNtm2fBLRCPxVDZQ+D4NotKCAFkkyKfsW/w0IYqy3f
7pp1HmmfBNbnV7F8ZnN6Z9NkW7fn2d2DnM+qH9HAp1KqFRz/vBycN5PgTKlCXYc2cYm+jUVE76va
hk1VY9GbGijMrNvYdQM4lO/VR0/Th1QgQ663BVF+cTMAlHJyiz5oe8uSWminbk8xoMKDRuDKZLng
CqT5eM2ZzKnUEPE408s8ou00WXGZXqwJLymJ6jXzpKx0s1cWDnNmBO9AdI52BbU+5uDdUAjVgu0X
7U5XdWsJd1EIKsld0qR1khZICefqfp7eBcmTDonNCgsHwGunC55sPImYmWyzXmYApTqomB8ktFpu
nT72zdAH3tvhpc1g/YMIfU0ZpH2HEIjojYobdFYLFbF7s6YObkYXf8gHuNekzUWptDsT/ekMxljs
T1L+Qvki/I9Az+nSElzBmh3bipo7udt5PEFoXCIls+xScMoMm9opOzGpoYDHYDEA6KQnbG+AbWzr
80flPzt0u/8X57ABG70zlDwcpz4Wv5v4kDH7gxihuGb/LRQbjo8CzAmOofmB9POm9Vj3F0VwEAWW
u8UAUR3duH75OwgmuNJ0OWO7hgkmwQjH53vrh5y9VeFKHJOro7aXGa7Bm2eWetypkaIN0gavsR1O
q8k7A9xXW+PwCczcTiTsJ+oFO8qIeoMw0sj3gGNpdiDzF+TZCVnQaIoth5p35JvPhT6v3BpI0T6Y
dUhUAX8asJsLOVj9P68Ad4wQkr8ET7GL4Z3ClJ08SNry2AXMRm2d4HBnuVzDxnoRBEDzwsFaiAYK
XyISNRZaAdxt6Pjp0llcR2AEl2OYpFhd2C1Zg6jmgFvnaAl5ktmGqCQ60LYCY5urAx+aFK1kmoRs
DC4fOXOGOQX1RBBIycIC8buPwWFRSz2JM2Tk8lzH75yHFGIYfj9Jfz0EI8BvQHmGlz7BiePLKvaW
a0nVZ2CqVOeBNDwKcaAbs47GrzEB1KOAUvdjsAldXRIQ2i2QbeXq7WIuel5poUBX6nftjFyxolrr
HWPvkQU1I/1eBG88BiiXeCUzy0hedBJJA+i5z9DbcKQAQdM3gpN8AyuDvQEEXp9T1sFGCIkdBSOU
mVGMWvzysM6Ayyi0UH2x7qCooZ2EU+5ELgeuSLErbYl1BngCdVFCdyR0ZEVT8kPRj73rr+DXbGFg
zmNdCuMQ9LLA1v/rOqDQSm74iE1JagF+na474EJxv5pE1/5J7xHQAD2ME0NiApKRXrx7M2mRCdzl
GTj8li0j4dHW2PmZRNY3W+DRrFFKSS6oPIAauErxEITcJnG6NJKIMV2kYEsYqr+isS0YgDVEISUQ
eQT3Sz3GMOorvanvSAydpy+g/VvejZNFWOKoLpzlkH/TqMMeyAdMPVBjlZTGzVPzV0eGSiCZIHET
rhCxs2idNAWMxPpNP5fyoVU4sXQAMX7QD+6CJ+CyVzZSHvxXE2tmS4uX7NmCvc2nwlum+n6hC6SQ
lifR6xsV0ztuFipMnciiJ8ksoGpAbe4Yfm2d4Jb+riKlFMRVOWDyZV1fEY8RLlBJpkaAQV7Pp041
cGk6l1yRaupKSx8Fik+Mvz40i9U1YykBRuxiRtgDukGkNIJwk+zVasYnitYPyURALVbXAIXGj3yk
jg6fmawOYI5W3dNAPFk6Akxi6Eth5lD7P25IajjePnsE5cER4yuLHzG/c91GIeI+SOtth+lg1KGm
CJu/g8lIc2WfdLta9lnsOdRNH5o9AAgVzT3Ki0uuYGZ5Gun3304+9f/q6lf9rnFGDEDE3k+Xow44
lzKBnO157X1/D21rJvwIPUdyJL2snIJCWpGaks8nFzyhHBioeiVr7zw0nozinNHsa3fI4IyJ6RYv
k1gSHlMfMqD8Fr9CkItRSlr3ZxmvBYZJfRhSmdoM0Lyb0OXYBh5C5dtahjqTUJfo4aq+DoO0SrIN
Wq1/UMdyTw2k3aqiJHNjnq8ZGpr2A8lux5/RNwPARGuSOAsnfa1ddGQ1kgI3L+k4sj1yTC1vH1GP
zLBPpgOpUxvgH0pLcGruzv8rMBgCerXrRsgKxM33j54KMhluztn8uzL3pqyTsL4sTxCwt8tIx2Ow
MUEohr8tZxOwZN5ZhA0l50Ribnyq1fbbNQHHWDEhuJEyjzmsK/n+KeiY4dfyEWQpe8+z79jXxd88
5gzM104ek16JGfzDemUrwEJPlLqB2e3Py+9rYAA8QtNfjfJ5gm0ZdB4aaYGJ8Wy3jtaj2rsDHtcY
jy+GRSNPz6njo5Eb4VVkIxCBbVZU+xzR4po2kG3w0IiA6vzYUviEMpn5EVEL99su3yiAoYZVW6Y7
w1pg7lrwTbUwMPWgxeyNUu8pLYE1A76KpQUrdGvd2jBGr/DaT09FeZ5oRpBIezrg8AefYhVbf0B/
KKqaKdDDzNo08SXrKueDozBbgaahziJ69AAv3AErB3KS/GcBV5TVEl6h13Wllv8zGqkbdYjFqyPm
ej6f3UU3q9ho9sPzBRwFRZ0LA48R+is8lKcLGpWJRx6wEipDQakv0y2t3/b1WLpkUJ/zz6Bx5tJ/
Kj/0Gpr0uTAO6frTk2K5fGZSRFeWiKpZycsOunPBi2CEzhK44F3P0590YcF7Pwk7/Mg9eRFi9ukt
CT+EaKVHC+dWcK1YhqGIJfvBFYtQ/X36TWc+LHyDLH4ocO5qeXis5ayH+ydS9uxBCuQ2IgJlf600
As8oQSIRqA9h1V3nDIWQF/t3VJ8l2m0TZ3eKR7le49aOmXut6Sc5Kne0gqvBUSkYWenmMJuzIWSI
OI4H5jvS7so0BtYxOICd/Lx1xeYhqm2Ap+dlRkLNZ7fpPaSs9mksRF6sE/xzDnK4qSZlNrUSLM1f
Zf/EEInoL8ojTG1t5iB7Gg4WLMBBkhimqJcBdggjO/Mc5U/I4ZAcn8rxY52VC0+r8Z05ziSuccb9
VX72Fkv0kRMSy8Pa4sWe9kaIw2QqUjN4PMtB6yM8att/9AFOB8oytSgbDiKxX8ob73G2X32A6FqF
AhgvOrGFL7zaKinbleNHj5EPBwgJAeZRgyP8OuleUh+U2NEVs8afli3/2jqWtT0YdJmcduKBpoUf
pQJyDNH4IlKOvwYZDRN7kKgy4r+ngFQZ9TNRv69iq3frm6lOjz7FqDvBSX5rDJnBZGSkrOXDlyrZ
P+wCmEwUBCFB9IHWuZDpbjSD7pdSIILuQKohUGhHKRwOkPzEh2cTtZfFiIxJahxJl6BAM7y22h64
8+NjEinxcAnBARKjySsH9HsLGTw2Pn+GEUcc4xK7RdcbXAftJ7wRBwdy1pr84BmdnpAfWAlr+bQz
gngzzUfMiZz9HGV6o5UhWLThlewWX0/q4PH5oezurn+KUItFMcEx2M3B3wC8+7I4dncfQOeEQ+rr
V5v6bC5dG7pvIfPEvYuTXb7EpLooyXM9GQG89bVwSxf8FOHK2XDBlOT5Tc65FnEhR2KRlzMW0T95
ZYZSvRd4gYKGQGET8amJVtWZdRNyvlCaMNsC9FbLvQcB4dIHlbDb3aFUl0Ny/Qc030OSupmn1eYH
VMYwmxOtN97OLSp07W7WY7lCAAc8NwPpM1nb77cPoPONq09pg90sYvZ/WilPDeMHwlB6LpSeWopA
kFDVEmFJxtKeniPaJFDcelXnh9VNsZeCFh6phhcNvGxEZXftsklVeGRiIe52+MwJXFiPNYPH8mz3
gLf6pUF8hOoBEz1hfNbkntfDzJTBFagJ89JSR0C6TiiJYNWmJNjLlJZLcsoraSkpWnVio/7z8eWP
9QZcsxSFt4icCYs53Jv4UNnBVd6/S3SxD6cw6bLNar+nodT5m91ttdAWUP3KkTcglH8cKKPz4IRu
7aIw/D9yeeDc9VjPaw5lonfRAxQcHn+aVF2XdV6ZVCjSRNezUnecX7AXvTxUnp1GgHbMWa+leMfz
0b97pot+PhcWs8mSXISGajYoR3a9islIm0iMgdjFQP2sITYzNRBLA40kiPKGE8BOmtjw9qcrG6Eh
IUhznozeoLoUuZiMzrr9BqG3g0TIQuUh3V1v8yUgeSeHLkHQAFmQyfU8YE8IldL7UPUDremymkll
GFPGSSjBdKymRaWtxL5J2orVsRqzyXKDnZ7HxdOmNSPs75NOqAlMIogqTxSm1UmtvRi3ctA790Tw
5xLR16qlR095X81d7s6mhtFmXeLX3kF2+QDEtAB/ZhNCZgKR1EPUWJ9+04UOnSJRpb4skLEB/TtL
OmiaYfLcH1TV8FWjzdQJzXJ9fGXCDaFP3z8lzT0qLakxLEe+OiHWnZz6nTvn0Yz/U9DatrUO+/Y6
ZnWjgWMamPsgBiKhskFKef0Aj7LhgOUvboJ0epf/cAcjQ6ixyDWV4yfCL1dJwOKUpuluCp3tpXKg
cBTa0SxMF7a4s0Lb6zg8QzUacIZnKoHwTvX55Z4Db0DPOkXkSL6ESeZr62TvwgTCZdJykI37TZxM
O1hmlNw3Heeluj9jcGxjpiVBsy0eGGou8rP2GWhQucVy85JZ56VrHHNUKWOM7+/Auy/BbClkBMLM
xLSPMrMfe/VEcze6BSW5ZnX7OqhOfy2MgAb0TIRoo8L0eYgEo/wNidjHEEWu7PaOL1hT5kvEQuxt
p4I64zpoyZJDjtJjsov5uC1kD4ygopLDDeaMsO7eKEVAWgCYvVNaegfACxu4uwPFaVDUm/pOjmiX
G4zdtZX/KEkYxgSf2JuvUFrBGRo++fpsQpydFICQTO5/lJ0/rQ8IccTjSlRazO1/C5NlVsU9/xOX
09qMHYhCRQyxvnnKE/aGm+ZGvxBkEKbcTJC2O4W2OPTifMfLmfpw7FnGUKGCcg4v+5QaMFh+f2zp
/DOQVeFnVkhUVqX1DGVtLzFNzaR/yY159AS/ZHo4HbzzyLSbGAYvgbOf+CMUV60igIg7AWJ0BkRM
i5yrjpTyzsKELsR8gKz0BTY2hMKIU8v4tvSt02L9NceGd9Lernc3bYQBfhaPU0DcPgJtCfUlRRW3
WuIiNwS7fmYklo2nXRIrSZ12zYxuo1NstLSbqCJYihc7FKTu8AohXNlTXHUz0ZbGXPl1ahAoj9uO
98Bjx8sW3cHZmQZxB7IBObTRTpaPWGlQyG7AZEV5tkzZvYSb6UmjG6EJUt175sh1OK19JjN2cel5
6RxBpJHGALp2w+Foe8tbaT/k+ubLUxevt2lqvcpRQKpfRfsJi84nzpdfuaTtoEcWJ3oFkeG5NmGH
EH9LxF40Bil57JRD+9YhkoCHJLXd+R5xwSexHZSf9OV2s1rLoZo+nY36PPGQG5ONA4pdk4nP/By2
COU5pWTEODaXKu7tDOVf0Uvx3zi0vQhUy8vHrA6CWtm5swMQ6FeBV5LhVcbEqRAiMyI4yVDxjyDe
VIVfn6JTOTIX25M8bycEmZy7F1nqi7+R8AY4SIXh6tNYgh0RjODtUoKflN1jajXSL1oJE46s1eHV
x1SnRZn1R9voBeuS4s6tqRsOBNL9F0kfI73YABBe4zK5gYI8eZ4nWwLReb08YU+Gn56tTxMl9BzV
XDa0hU/Qh7aqpPCj6/udvJCq5lSzWeK2m0g082tMCjfLt3sp4L0rSrapBSGbLF3gp+pWWVqtoZ+z
FUkXzryrIt9ndz7CFuWtClRZTcAtOgWcz+Nw+oJeJd8qr7zlioSOuHnkJfT+s4p5Cm/CZd5RkUqh
8J6snryY/f75vuGZsEt3sWLYSv7XTXg53lqNaqqOLkT7VCWUEEEy3Yq/jxWF5PGbHeh89Ez3jS7K
3PFxibnVDViDFmW7vz+SxnGn5G26mD4S4fLTTnlPubvIaUwMchsMyAb0tQyPZXqVofTdgtwPQ/YG
3IuD5Q0ovyVDXAOUkSWNXmaizXlBbjWT55L+VQyXP2Hz/by6Fyug5oEnKYc1psiBp4jpWdppXVuH
Crw5Z2RpKqpUAd0QxLPAJv2c5rEsp9en4165geBxoeIEH7pdF8LEph5TKAmpc/MNXZCWpFpije/N
vvZLYSZYekyhvgxGA7KiCi/TwGF3RtntxJHKmvt80Pp7yKbkVGktbFqJT2bZdK9drOhgaEAJuZaj
uT1Kdwh/hw6x9oIYGe4OwJNr9TTPTSBSmCJn4aX2jVTtxLJBxFz9OuaS9FjOtX62r9k18kT0OFJ+
jH2NoiASB5LZ+vHkIi9Ftw4YMgkyEK1MvNCdAErH3YtIoN+hP28kf2sOFouSBydgkhHCQUIcpGBa
8i02EWHRkNfC49z+MSfkESMEA1wC9iAkpz6US0WbITLuOCE4xyEqB2IJ5zAZNFNqEgmhgfz5LTov
Pd8Ibxym7QSwtQZ0Ppqq1NbZlc9tOJgnJ/KhFnoQsST/Gk7FDSqSgg7wqiJx5svqdXbTXZzdGAL8
zbj60sVjoEghHDQjR6+5eiDq2J8XqU7vaPxDpk1cwi0u3J0fdtVrmBS2rnNDykdP6x48Ykenx6ez
uGXGhMvQAIpsxgDO4c8P94lL1i9STRFGcPrjCZoGPLadeE4vun2Ao6v9SD1+VBkbyvKPxaFjn83q
4Naimg0amkCp9xpj25a3T42s5C9zouqHzpspKbYl5dTuf7qG/40lbHi1H35CGZOib/z92W1HiVYR
vctnZTAFSeX/g7kXzu/+qIiH8s343JHIuOZJdriko62TI2jgbVIBTdKtQRLWsdGUAhbn7ZokUjTa
OO3kAJ+Sa5nadwcHJ36M4mH/95rZ0ZyNkY8spZ8X99hpEkDZ5a5oFYQAcJHP2PYFXy2bvpDrdbLx
IkmXa69u8n1Fc6l0kEomLYZXgBsiTfLbFyHpOlWlE085me4T3n7/r0ATxgw9gEtk/AHCCMmu2389
WIa67SApn+MiIMvEXbmS+hO88YVZ/e7AYDrMpJf+S3KWMfG7uh0LV5Scc3CwyxFURPHDOxTlp9e1
WuMj5t4u327sI4yKmutj30wwX15mOnlVWZes3rtVniUlrjIfXvC4LocZhnGkiuQObGsjYa/RQISi
BERanflT5tfb3ViNKA59RzbgdD43meUViFk7RIPqCbFu6uj5UpQ3D1tgwmklw9lutJMAL3ZesfAE
saYf0ph+OoD/3HgSv69Ne/sX95BrAerGfH0glyZ5puVMQE4xnFbi7DKYaYGa/kfHDtlLaDdeowRV
i3fcKWtq4VAyWO/5TdokNMSLIJfEqiEZJGeeUr37rg6lubHK0gWWORaRMsr6ZxuzJK/l69+h5eLN
B8iArRezXS5owIxhQ0UplTfyeY0JxEhWV/+MNtm7EusfjvccceaS4hXa3Gd5niRLLvhM7zdbYIyN
1Co3ibj2w+EWr7Wa+bBfgfW6ERBQIcRGv8bFaC7oRAUm9ZK+9C83oarBxqxJ8X+KbH0hS8pn3r+t
sDvMFQ2oLnyJTHcH+qDPCP4ZmF78NTr98g+IM7ERzYBaZFUc7N4QmtO0eNxo+VN3IRjx9/a6E6H9
TRDF5bEydanQq4VU9nICmD0d76m5+4Ty0QieebmRLs2GkzIpj25HCwbzM1YyUkWPJNl2RbhoNzka
w7SG8POQzuaW9CUkFakgSlpTgwAY450H6J3+siNpG3rtYVEJXbN6YmNTBhVinQnP+20zdz0pbx8S
zo89EENsn5oJGrm58JOB4gaU5lwYYs5jGgNkm4DtamOAqsEc6Sh3ONSGt7eKkRNKPeldisScygeo
FWYX24+b1Mt3icbFI3MuikDgfro+WbOb+NKw7rQaXcJrz7cSCiX+3GiTIiRSXyfECw9unoKVp8Qo
W7m3QOQ7mSJyq8Hx67eBv0Qu4+r51FApfM2sYjW8tGqsF0ciJRtdqDE8n4v4j5ubLzk0Hsb1cy1u
Ax0RiX+O3NsA0NvtunWHvHvSgiiPWrs/u4SvaGNcYVjvkO10YRnnx9Z/1KBQ5GT0Og5po0KRJp/a
8s1AT8u6u71EDSgH5xcMohIrpDDVh8IvdwZdBXSnILOW9M+NTJveeDwBqhnJlpGtKXfS1kGHzIzi
xZuG87lTmn833yes34yBcut8IfDSvO8HuXx5Ip83PNYu0p1T4Tn93w1mDojpWC+9VcYQAnbIRId9
q3BEp+FvsHydr/fUzrXNpeYQacOtKvfLePAeqHb/BmfoiCsp6DlGsya6NyP3IwidCghMuZrKykC5
1mrTvBmUV+NxtGdI17mL491TGBGbV4zJ7e9RmLx6/yQbMXgEQ0et6bb3dztVh6Co58HpcWSdNspO
g1W8CtAhRRxE69P3VSEa7nS51hBtG5xxIkcu9CQ54PurlbsvvTTmy42C5ZiZiheVYmqiDt4qSy5s
nQCMcrCdvJ7ToT4rMHODZ/7R5CNhAQrnFvMZspllL99zhMl9/j1BXJHrPIw+HrX2Mgq6lGrJSMBx
5YgpLbr4o8Q82r+s8E1IS83AzRNb/9QCTtFgrC5EgP8sWZsT3O3jiXfUPNx3JNl+hDYFnx8hU9AP
cvniLG6q36XISwqi7nfKh11+27i8bh9XyKTEwIX+krkQmCuFOWGsNpxirZNke695VyoY/MHZb4dX
0f//s/I1wfcQlUWwn9uPDSsAQdNniapl+fe++IMfe+ECwwKgWzvMXhxPREyYCEw2MVCQgEouHA7j
/Q9Y72V6oyl5qMrtnS5jW/Z49vUkjA6S0UB/egPNsthMTGUfyLT6I3sYWhBCS2zeAel7fO8jkli7
48hFsgKJVqwSlRwrjkMxrb6Odfcd8qXUcKPQx3NfviWrwswJTpKKoJ8dEotGuAmaEOqf2pKWMb1j
1IEx2sKDfChTKrvt0e1ZLe+t5x0QHDoFGiiPK9/fsOyt3mNQnLP1gQIeVNlo3Bp9DVoFkltcOKAT
h3l7D1+gv7Se91/HpwIpQppvsnZ+j/JOVuMvDfTZmiZMELgJyJkDdRSCMTYPJG0X/SNchHizOc79
053ElzlWHtpxiT5TfQp7GZi1/v67mkLE9MSA3gSmrXg6ssSJkMZWK9ImbKDZ+JFMoltxa5qmKziB
hjJF8oi/5hXCsyV47CC5d3Wvgfzp0y7C+bFe1p+Gz0VmRZDcnD2CgOCWQzSSd3NTr+TcSPZRio1G
CwXNjuFLBPy0CuTJuD7YPTz9talfkKh4h/R9KSQG46EA9Qr4ytKZcrysZvaWeddYZxI8i2iDreq6
enGff2JHS+oGQTBcu2LRzdq1VMeautuqTNTze/7qpzFCplALhYK8mwoZQw0LuMuOM3pVok/+uKvL
O3mgLjocmd7l3OkNxIjhPi4sKRCvCDaQqgcxY+KDGFlXc38aclRYFwyGNcrGyM1+Sle61TlpPUfW
bkx98FqV251lSgW0Rm9XKXZlau5061yytT4i0/ZJPFcUoseMo2QM1PzDeBYG6zpuq5GWawxV260L
pnrtALNkAyLYjJ8YV+b5pJFjNZBao/sRExrjc2rPPUcOUhuRDM+8owmWF/bhvSEYbmfTsGYRin6S
E49BO8MNhLEePvKXWMvpSYH4dZ2vc5FhOx+fvZp2bWc0Pe98twpJPoHa2F6J40+OzKkD9qDKnw88
N5LvUcssECHOqsw9tTPVW8Jsex4cdAx8Af5C1rs2P471JecfZUI31lbOGwgBX7zP0A9/7fzQdyYb
XbbKQI2JtYMA9EfqRIPnVY9tvCzPiuaIkPYW0+KHcwwf7IIapnbUZ6gY5YhNsfcO4+CVfgTCXzbz
PTBX8wZ2iT4T1JCu4wVO1o7d2IbqdrvB1um8UuYC75kWGWyjAEClrIbGwdbSFipoSK89xOhJoxGG
ZB15vB6YWGCXJEDl+S/bVvik7BK0XeOlqWZpRvm1wYZTgxhvGleqsyLDmrVfBA7hdiH2Zu3ikFgC
7yj8T2LH+8FNvMQXt8RryW3EeJhm0vMghk2Vou1L3D6e4ojvWcrCEx2G+Z3M4L+2rPwCI+kPpDQ7
Wx+k5XM6BDeZiYQ0izja3dUkrC3AgMtOKqgs5l350mSVI2oAcNZ8nkP1gA1w9VIGF0LyFGgDQeGx
4vSg7+jIcNthsQ7NKjxmv6d8SxXG0+jIER6ZsL3D4sJua+zzBba+xPtL+9WFEJLS/i5aq5ONR+1l
TFdcl5DDGscOiaR/Q01/qX0n6A1w06ZtGu1DgXFoDCWoQVAq5Adja0wSZcPi8Xfr5VNKGrXgc2jB
w8iHpYkb3OgvaPtX4r/aQMyDxPwmqOAzJeiI3ojwQ9jBqH0E7y0pBYAUljj6q+SMXNulgfM5hE4p
Mj1Fr8mhghIULswCbVDsPfrU/G3ns+CRY5uFLthIqnmQPkek+I8mzxd+eK1UG29MA+o0bTbYp5c2
frP9m+olEEcrztosu7RGfmdbw2/5wQqv91nUWqRjIjzn9+e9Vi2mr0eCyH3ONXJXqjfYeSYLi7ON
hnXALmG86uYMx4ox93nP7qNckaSQtcriIw6z7dlJYfkylricSzpLSxIge5hubY/eJz72/lh4wFvh
kwo912d+47lLXJLBBNh1YClRW4aG02QOYljWfyqqjtQw2DSAKDIaUKgsP1Ws2mCRFAT/7101jO//
i1aS1t7CUeo8+C+MwomkrCzxoJUmPgHs2y+zqOqBqgUTriKdzdKt5+gvCE3/4rWw+ekI56JQPOmZ
HOcMa2UgMbEqEoS3tGAL4cXA645BojcE9n2B25v3gBH+TOqs8MB/iJw0T41eX4OU9qVtChcWrgNc
MDenIECdIi00NA0Yu7DiCLUFLyozIckmVV57zGkAhdpWREs79Pn+hmi1EEuOnL8S2jTUu4JTP4rY
qBShRfi1Hvj+t6sL8vsKLIB7/0oaQjBb3ZgIkOM9KU0JhwC7ESa5oFxb3cCwRYjce6mwq9dXf5PF
7NdcxGUOLp8Ytod7A02v9aa+QrO9wjiGZUq7dx0Dzzs8xneFfv72S+k3haxK4dAFf3nNNjnnJPEY
69Sd6z5STAfkkIewVjvJnimReZKUNscuN1nmGupFF1Wt9sM6TOF/Y1hybljbW1ztibUsoSRwKAtQ
jrUeCKWJ18+JSIMDx/mx6Sx94Xvz7FlToTKBIL5ZONFafoA6641gU6ptqBHpFysqwkU8HlBtak8G
zpkW1HP/wZGK49nKdEKT4lgIViVyLtFMxWYru6BgNm0eu0nUXTz0XoHLTbZA1rR3PvWUgZOOriGK
jG98KuMDS7rryxuxWDhrnFCl5/z8Hgshb3FwvwW6DGC+4VtbSYdrTd0j6ZsrEbLDrbU0Jej55aXT
uy+ACKwB+3ceuCry+dCf9eoBiBsosMYN0WLQ5qu2oCC12F1rxwkbmFQLHkQpCCs0qLlP8+0KSnaO
Bmqchxv3CWH7unAaYtNJqZueEHb6Zwn4qGQQRVkg7y5RCqTCZqSK8pjj4pCPk193vxJwt7B8FXmk
NyjdR0VtwjaTE/EcawbFcDo6Qah7lXNW/1s/54s3TfE6NI2ZaRBwsssdRgrW3CGjHHQVYnz1Qwwb
LXFkgL0e2HmLASQEtZGJnGfm/6phvGmRsIiRUxypo71ObcdovIpRn4UZac8zW8CR8NLVE8kU7rZK
ZY0u6ZoARFnohwcNoLwcqnfkV4eWIBnw/P3CoUCmkMoCa1dffa5NY28eSmqccMRGX3KcTxOTPFKO
o+bzdzqyiYDNfMnK6RofUjoseLBNRIn7wL9P8T3tiwZvEampFoUVYhHEU5EWoEislMH1fSFnK7/k
AAmMrE+pogCU48IBDnShWq89EgrBAdNioq7/OFiw0Wjj30C5eDN6tu8okHnPSq2kQiyZ+a+2Ro1a
tOzvyxE28eoRAzTc0/ijxJLI6mM+rebOD9LnZsCTNa/4Z4NxYEL2qpX8jt120HZ50ZaJHVZavIWJ
K0trAdhht4gj41dmsHEM7Ct1JFfntzJm4Jos6niezBEa+/MYpQessXPR29JdMzP0lEZrlYrKlVxt
Az7EL7JNaEPwVW3RfemqQL+buCTzU6bsQtBs6V+5LT7bQ09AHSiTsOmIWKI4OnaeIcpLWR174cCl
HwAW1NZe6z+YqraZgzYYV00FLG0HSXr7yCZiValaQcmKoqAPTyF0pyuyQsA+/8f5DxVjM+SOxx4/
GPrOWCR6PTWNDHD+iJ8m8Dn/PAbcalUVpPsYdxytXSDFp2UlU9G0qdddZ2rMun+UR93laOdwdSHR
FPKhhyq4eso5gEsip25ABBZRrcs2HwyC/EzySahY1+6tL6VCXziRRM4JtBlSL6nHcY6CpQ8SWoq8
t9Yc3AjXKgdvXISHjZWrtdLoZgL87xU+LXC11inDNgOjlyAHv2WUfC2esc54YPa3vV2/+RdKBQtK
eU9Bzm/I6G3j8WVU1wRLieirxrCI1794eF5lzSKDpTmE+3HW9WosARYvNkrMB6q2NnKkUaU2GQMg
LbxMKsyHOX6k2WvJ2wAuogSnFUeKhExIriOadFtQVZBWsFgVrgvGusWB9q+qU6YfeSNRp823lY51
uLxsYyb+D4lV+JLXyNuvZn8UGxczWGk4hyVyUS26nL9LgwoqNmhbq2mMnEUPr4WaxqhRnS6m32L9
EHDp1R9ZHeSuQiV3+m2kEEClASz3E3c4Hd+k7xZoGXKIdf6DFdmZ0Lp5224DN9lovS4KPzK6gIQG
OHc3vo3jAFt9ZgncFUX5JnN+0FTtz0oeAxaRUMNEgm7RF5K325XpMVNhohn+J8TyZXwvmhcwICkO
WMwlOwnRMpXl/ZMsZws4PK0bRHdT3wYX6GzZvAhDoemHi7gEc4wd2Thuceq8oyEiY1jzzS+zYmh1
X7mTjnOasT0TxFsEEQ4VSL1jIEAKbGx8MpDXGd8gbtYfLW0lguJ3ltd+TM5KHSpziZAC9EbKKpNc
DPiCjXJNGW/15uJzTDfzw1zjDcp1gg0yYvvHIqw+mxGu4DYm33J/AFFafwfXmNR1IzVG5vvohWfV
996jqpJgQVorVyifR0RmXNXA+333kThzdCwCH8WU92YoVmoJ3Ikn2ivWtit1o/2Is1iIVDfGNW7t
UZe+pxVclDykmYXas6uLsS4QB5snUZKoF1QLzXQB46511LS5BmBE5IETLB2PfYPtR29WY2emH0oK
qc2bzIfJSBVWG+rdA4fUXZyeFNWJvsjby1gwNd+5xFn75SEpunvs4SxDO9DduDMjAcHcRpRlJ39Y
w141mVFMVNCIRYJncnekKnih0ainZYHFhYCcAPuxp1zBLnQcwCJYECrH7fhoKqODh0YzTcr0JJxF
rjc6QINxHclhckxS+s54HrtKZP8kcVXXUhKdvuyYtRBtbPto1DVsPcGi7MmCYntX6iSlVE2CerN8
bZcM7yh4PTr1M9ahtUBqDNOSMsAxRV6Dk5/yDz27GM7f56AQDjk/2WZJt/+EetqkPoDLorYBDKEo
HCBWWRxarKqh84jdnyHffTfK3KYwDu+sxwZAHFJM+76gN3xIkVRsqg52M0UzWJ6PBIdeUsPkig5x
D3BQb0sDUGBMnDkYPFY/Ekc2tTwmqgPySfm6OVJGiE3X/msWt1Fh7l/mNI25rS3tOcJIYEBhV1tr
HGnZVFGH2TDR1SUl7vGjPEQyZjFMPI2UVII8FKvJbvWP2QyNZFfPk2QDzDfecnkkIa7+tMehb73k
m8Zl2ekceuieFr2uMwa896ef4F+DFxjIPEu7S/2gl2WTY6NtqgrC79v0R0jw/vdzhERTRcD6q+fc
Qg09C3M7OaYXrXYD6MtX6+FLHHuAq9oABTLPYTFpWLdUFsE6ZA8ygzvfeQ/+CHSKCz+xgL0olfsP
GSRagyfcNi41j7u+UjGbdUqw7ppxP8BMTOlx68v8CGwDOaKkbHaThcaCXUm/Dwgx11pqTxn0eeh9
ZDtJO67NvJEGpgxIKYO0tEQoiFmjWjvhc1frGIKQdRbmOOzFR8Q/a9qzdnqBAarZigmUsvODkZbI
8Qagh4oZFxBF7oO1kKSOfXqd0KHochkmUwtIgrjB6EPTDW8v8c9fpwbBNn/aCmXRqmlDhvQNnzUC
yUnuRSRaM9nM6hVB42EtkEQRVQ5bRsL9SqygYnqFT9YyqiW7vGq4Jsz6fKSClTBuX9GDtOFzPmXO
Dvp88fCzj39MHRV0WLeXRG63YsUnZkHotH8aluViyXH+vqtxeAUN/fWVFoie3gWJUgRNPG24YmYx
H8ahqel1GUTtZjng4uoKwx5uwS2SdWJnHzKdPa1UENC+n8+DbdY/UY9D6eCAqGoLhfQqcAv7nYQH
wVITrzwZizaPF2nPVZm3zd5WUK8lvFKFRt7kpJN40WJcNW/OMLED2/Mny7g4i8bKRzljYjF4CcPk
jYb6bgLUOkwlEI5OyGVzDaT5nCqax6QGzcALhnOsahW8YJ3W8fGKNGmQFCbwqS115zd6ONZ2gkMi
ODG+nFJGActtswLRhDT+P5mCBkGHS+/VnCNBbRLMTqBonRSGYrgJ0Agr53doQP273Nf0hwYAOXg+
TQZwqEXtxUIUkFs4/baO63shZxbyG8FFrBntM8bfJVWwm2Y4zZnWb8mP9HnW23WwYOVDLROqprju
1EeqN/NLD7NCDX+qLGS8CL3BDPIMg9l1OnqyZbpyDEWRpUDDiNxGGLxxirYrYwuydkiGIf90EkE4
zwp8lZp3icnTB1Wn0x+abjq7B4XM9pRC+LzmnRDQ0S/0le6wTlN3T0L2pNokq2RHQBc1wAVcnD7/
WbCBtMV+Wi4BZQ2RV1/4e+VAI1TEBZgmBkzC+FQRRMvHbGgXroF4OjslPPPmOGnU6UMLBTGnTXhL
APWO6Z1cvOqq6dXO358KbFFEI8w72WZoB7ZdFq5I9xzUO3qavs9KBCgb51uf7I0QrjilLSZK1meN
3L11DFhvZjVGGzVFBfwukNLNjD90HhJOr03AnNOk9lcLSp6N6S7jcGepTzbatbAO+9FIY3mAPJqM
RGQvdXQm02sSfyNPiTPtE9gq9N5jt6OP/mKcrMB1gUw+u5ZWiDlFsim5UlFlkTLAlC9IVGsn7bqL
sZ0IvVkpz9jfzLaE8llqr2Q0gbH6h0hMOiayMwyUe7d9oh5puPDH/H055RPpXyAcH5g5wZMvNuQH
mq0xQNPDrYLpqpExWb+NVR/MrfDs8KwcDItjhf5eD06BgZGo8iWsOv3UL5NR4TPHpnf8sMbn8ZY3
bxfUDRoPwO19vYBiSRrR9P98pNJHO73e8D6CZ1wOnee+fXODMshg7LvbK1USK9cmRoJMS4Uzgtmi
kCKLjcPkGgtGRZEyXpmvE+LorwAjJQZdWKW2BXOOqd43hLl+jPQYsvAt7xI0UT4j9SID+0zFL1Ew
Nf5x6C4TmEViR8EcQS7QzyUKXyRERw7wTr7SlEmW+sN9sgCIZQAXzwRfJvkht9VCjAZXY2oo1CJi
DgPFda9UuKZQ2QePNznGPU9a0g3ysawvXAzNUq2qsCiVvXeUuxudsrIfPRW0Pcew/kddoFmFXlZF
MwvoglSaC6d8Ldvp+00V4ZEYbYDVhNCacZ0P2ye9pgeqpAIWzYmOcbuzVljUTOvZxE3/3EUOvhiF
ur6RU2pVz+iZGeA0sdI48XLGTR1wl5q+3WKja6uWK5MjnhZOxRqPsRt56llKdmmym1mys+dhUw97
31O0xLHSevUTx/n8dVVVcYrcHurb7+OSheB79spuJLDe+lYxd8lKEBbt4P516LsfMeop+Y8A4l8M
hofL6zkoS+3DX5LfxJ4rkBOxoN015V5m94JGy9XgstAj3CIEGzTpnBLjTaSX6F4cveUxrVK4nc1Q
R6FPhTrOBRw/dOcRQYR9RRduyBUM/knHxBfFPgBjaYic+I3QqWJCR2RbOrywMykyfbsXFmfnFdvt
aib3Rubq8Tv8XNegg2fRk5owgXH8cMwcjVH274AuziTbA31kG6Td03nzD6I/Ln8VBeSKSs1bgJ8D
TPR958SzvwYEqy3TwOBtajgzSXv71GCCQ02MaIlbIH69y0XhI09I39fL9nm5NDGFT3p5Z4gpQh8v
ZM7XJNFMUA+23bkWeafPC/+1wH1qqrkcXk8/g1AAsZgzXABbFeQzbuK1OGcbsrtHWACJqBYP1yxT
btKX72mWwGC2WYcHzKhQLDcudZC6nH8i/uLv1Nwvdwjn3U/YYY6m9aDt1LR53P0Adz8Y8QtgFuge
ycHxMZLaap+g9rJlwk3hFPfMnMY04DMmp6SntTa3hXCWiFf+4yGpHfz8DSbROomXsMdqaeeQHfFX
X39gUJ3oqTSzAQOmxH/jDKnriZ8XXaYryabWURGH578X+5wdI//dVDLaDN0M8JnAQOlNcOGxmm8m
DXL6xFbV8B66XRAu9hT7W0vEyHRRJncQPv4ryPCRrFUgl7+Q6FuVEm1QKVPSXruDJEnIDo5E+hth
im10sszvNuuOTihQwUA2ZvNPyQ44L/H9NyNEHv4lkG37c/QeYdbqD0q56Oy1L1xnk4iKOb6tdXE+
HDtoX0ddHalxe4eroq5kTUF00mygo1brnffN83v8dTxsK5GSfQe7+DgFrQ9iSvCCziz0e5jpAS3Z
fBWgKU0ZM+wji62XvWc2LsVJGk0a8Pa6f3lOeZRNWizj4KEGAb/bsniitUUAVn4qJCKKM/UW07WZ
lUk4+Ex0Q/L/Y3D6ldJHPzXmObLu7TsNWhHASZSX0wnCJ3gKF+Dr2OBYykqqEyMQ9pzgQloc/bQi
+rcCuyLOZalNYwjBWVi/x05uEiAyhiO+xvrHvoV/dWfIPy2wpV/rFOmJX7muZjHaOM23ANPMfjKj
n2mnddrf2MwjNTg/7Gqom7kU8V3og6MViwz6+IpUVlgOKC1i5ZZMKH07L5ZfsLExFD8A163T75V7
o4ull5lUPADwG1JSjnrJ0fQ7UVnUb+0PK94rtXZtSF2yt6ycT4bigCpUbRm3dnSbs9jGVPT+5AI0
sHAx5+ODM+FGZa/+hjhI6mKS5O6pws7yc4YGayJeOk3KIPA2fiBCsbZOBVHDmL50Xl1ToZGUPHwT
UJz3f3VL9qeUNaWnhi4b0IQvIRUaAhXZ9jNn23xSoOyfDO+YExpXuE8V7wG82kaQITwwTtdmMBqE
dqX9OXJ17aZQgBh/8fMic14ZEtvBplxCtnxdyfVc2aiLsVD4ePqIXyOt8DjxeMryWaG94HGJB5FP
nfBiYNz0iweDfXGWMZtldUYiFQghGBFSg0znkvhvT36s1NTeQETHtVHbPvjQ6mJzDgTqSp3tNUt9
SrLe0MQ+Il+KrwoD1U2P+LRTBurStAUmXSAvPD+EvcoHRu+dz4+wDM2IgI355uZ4q+RdO+i6qDp/
yvTI7h3aINSDUmrENqDX4azTR2S+eZfdv7kfe1PzxOqE6FmCeX0Fw6udT8JnZ4ZMaspkX62w1/+m
KQJtKc4TkN7OAi7ove9ih/m+GAfKXI9BSK65bPRBGaCwRF+yBFKceFnuKVHcSKEvC7wx32Vi/iEg
9gpepO9d2EQfuXy2ypn08L08zwl4Sh6C4zvN+cH/KntDzk8CqwmWN2NdyV1d8eZHs2AyzGQF8Qhs
42m4WVI5MKys7x7KFqzjSMjYgtZ/fuZ7xIJfTXgHdKdybxzFKZ8bGkm0Z15VLq9XBg+7LPIxXyC0
s0/OKX4DVxTOaSKn7PFV+STN075XYRAAZuvtQV/qz6tWYiccEeNNtp9GZE6PwcZWnTCgAxkNzA6K
akx9D08kd+aXVmqPt0l9SktTUAshxO3/xZcNJVtFclOIB/4MdkVTxzskVHlplmvUNpoXLM/EVPGp
4ppsWH1AmYVDjBvyM+SZtMP44bzpPZcmtjWIt8AQfEtI6bIdnYViLqWuLSISmrLI9LtL2ilGH0s1
5Ye9Ld9FJehvW6iiMyUJQFLT6kq2uLwnLOEwS8i5tjzQXeKbYUw/9KtaZNzvNUYrz+Oswf9XwgI0
EN/ifRUkUSF9bzegxiJQpqt3LrmeL+V57byiCzd4Mt7Qt8h+3f5wXcCsaOjNmpXEntMqX6fL4zaF
MXj8xauiRbcY3S/zX+vgj0BNu/2HcJmk/fAKnoDxqWAeATbC3v+wpJXQM9GKmDYwsoXf4qEm/w2h
sJsXAW5xJ9lzPHAzByD35MKDM0/+vvqwXnSbvDNQ8HDC2Fm9zj3RdhyKrYpHWqlm3Ue3jDfe4bNv
ayJZIO0E+XK1ODLBnh37acDehSSleyo+NpNO8LD0LVLHi1AQpffvamKoZdtcubAnq96oh9EDRMKW
rHtn9DXQEtGY4Jgx412JN+40mnejVOIISOJwasLwP0WZH2TB/0yfQSc1eI5A06rrRLbwXcAVmXIG
VQbCVBo6reVw+k+KuC3t9hUbRK+cZ/ZrwhjPLJgUZ1jLFkoavs8K7r7kcnobXt5TN8Tdpb1TBgMi
P7EfPlerd71Lzx1184wn3uiI3t7IhRr7SGL1SJMN2LVYlttCna01vR/Txb5ki/FDw/SJh7mhYb16
H+RFvbdGD0fywrxaqAXcwGXkbNv5sf8msF5QesHQD9F/qY6o8mA+8oXpfsT1WnXbI5laTPh5gl/Y
t8d6ZF8WsYd5WMnqrs0T+jPXl+mkLlbEo77t210aANBkmp/H3hE2okKwp3sfU88D2YNTHLrpIRW3
3oWTJ0HPM9rxL+kzzPtlxWDbd/Job3bUfTjUlBkMcJ0zpysOS5m543CIBoRp+V/b9bpVGlVSvmP/
gjEjAmodb+6fpfuESsv3pdhs/v3w8eRp9U+8NAQ8oxBWmpf6vTIyDoq/ViVD0peeFhLGURXbGxBM
H1ILWAaxZ4I2AqR2enp4HJD68iUPNOvdRUYYQ6YJAiWy3vRwIbtXMGf/piX6lztS/kl9cKNCNCCc
7qIysFWea0h9ZtEJxaLpTjgx+HHiXT9DhxvTgATMN6+z2YD4mMndUtqDO2MzZNRZIj4pv5eUe5Dt
YAKNWmcEygf93OWh8IPoLJJGBkNpiMwoYfoJe3IAj4fENgmBULJIWeEydm1pLtCwaGHS+VcKbr1k
inQJdAc8AXJrrRQbEHFxEQOIXZH2ctKk2aBaTOP5gobZIge1+mxxLIYc5LPMzECT7WvAmJlhGP4j
H2YqQ2y1T7IzzHyiOSGLxe9vE7F7StKpvX00BQJSgwGGMYtQ7AEPIl5HY8WuY87Yo0q+sLj29tsD
7CJxQ731s/GV4Ku+V/6MaqADjIulhutcmh93iW0Vwf2+RXuxvzAsk+Isp64P1njoG7uyLPHhAOaB
3CwhbzX+b6gZGrFMGfKg9t6DRJgr/VfeflsDkAeeQtms97x9xtxo2NgLNrZSi3YRojIK+kxhxKcn
5iZlWXMfo5bzyPGa3NIspR38b3Mzc+KuM1gB7qZj26Hq2+x7nqe+MugD7l0ToHUsLG7+THEYdrux
8qsQvenGeQNQqePPv4Ia5IF9FkEk18+mJ2CZ0ZgAG6lPc8DFtF8sQOQlIku70JCy0AwIItrqVAaX
B7jH1bSbNyw+DpAx3m/akLxsIW1Ni1WFbi7F9XIn1SqXMBT5hkGHFFFuDcBE1inC3zgg/5GMVtfJ
mmc88FG5yDFUzxf1ZGJrlj44ZEsg4hpR1ZxUI7fah1eBc7p9X9PnGjCRqUJSB0p/JVuAyjLDjUwL
MiRiNv5mec7+iOlYb+zBXAVGt4qxNMedTER+H0ATLrHTHDjtvOs0sQWbwrQsNRqb6P6w6RXgY89Q
hMu8L0lU9a85wzUGuOqV6gOjo/KTxmMQet7vnY51hES7WfvPoAj0etgb/doF7Wv9n3pD/gJ/n5tr
hRWyiv3dw6DLEroys7BVsfESYr8hascp7lZN+fbC9PsnFWLoKwDz/M+sTgjkxos5nmHwam5kvEGh
L+TBGXUUNsGi/wDIeiZOUuGR6PXydIvZ9HVnUQvRTb3swIWZ5pIx2zrKywiLwNaiO3KBAzEHyTrA
IOiKgi9SkeMVYSMNoI1USvxoYzfN5c49BXeQMjXZP+UfJ6/6ahtcAP7hSuDvWPW9UY9HoB+NbrDb
hvwViJEo+AIuWhe0zb2Sr71L2egMorIHizEHhjuzWJIKPXHdyY/2TYKUrNHmwSQ7spzQ/mdin9Fd
Ln8RiaLWQf8o0li0gehUrNysdXCvXcryjXrdrvWmGlcoJE0PGT0OddXtxW1uOwV69YEfXOzlperL
fkmb72E+hGt8CkAKrdzj3uJ3TBQ05E2ezIbjleEAJp6xtbX6JRoEk1Ue0cI2i2kz2UL/Gi52gqzl
JpZLnmOhngA1GXWz/6GWq4lBuyzjtGAWLYte3x2qmt/8geD5SdvzGyu1Z+fLAqJkdEBfu11U3Hbt
4wBqid2wI12WQ+ky0MHnqYVREtZysGnH4LuCmGrXt0zioQgvO8hPvlBMOiGW0sMUkQFF6S5U6xdl
U3GIH7LFVXMtrSta7uw2Sukb/FAzXrTqaRRPwr7IIgRC4BuQ6eimeLCEW/1JFwpcuSOA8CVBrPM6
HYuISR15C+xjouxX7othRmxhB2X8bvkWT3WOkAZhfqaCKu3oOnY7mVrirf1W7by4G3HIz1rjZrDw
lrWSskIEbEsOXFwezCt4kW0+i1dbM2ZKAyxMbDzhvcQxSI97kRVX7YLyd57vn5lEpJ6WEONmUR72
H/ddRyNbMStA7NK78RrOho/ZpJR2YAHa2rt8l+3Ma4CobrA45/Fm2OcBZynG71TtxbEA1vf9TxpE
mZyOxwTO3GwNpbykdtn3LlLEQJ77Aaf4Pq3qJUNS9bRfyHCY2TsNAswR/Gh8EAdwvFDtVYMrqhJ5
ii7QyQ22HZ8AX3M1bkdbmtpsmk1cngMztC87i1wExh1Qi27+AL5kWFtNEUVXUBUZnjtmBLzvC26i
4oNpcrcClqru2ftSSZADYM/2KZUzLH1+KD67PVUJW0iTSAk+ZqcXd6CcAW+7afwD+tkEeh72GUFX
NqvK9n0CMwpxl7/vK54NX6dy8L1luhAJN12oVXRrp111RHFlMLDrERViMKskRWsV18erVHB/d88i
23s6rrPTm+nCiYFG88NQNnLOhIqQdn9ocfosHsqdl4OPJLhpJIOjrxz3M63ADEcSiGauTB3DaUvH
lX3gYJwx5Mb6pnpw3RVmIp6npXObGoUh4xouneKW3eCoaHz14XXqj5GjSdkrsO7HpvyymjzZv/RH
HeanBk2kjN87MkSC/lVHAYOuEZjbCihMmEZBU5BEw40+XKstIDYXvmHhKvLrfyz9IBBt9VFUvpCI
D61UNgtyK6x0iBp2q2rRwQ/CY3cWvDQevZJWYVPlepPASxB2gHfS1ZwjBOB3GqDhdQawOI3cnUON
Zn/uJ8O3ZzJUe/v1uEPIzjas3ALrCZEqGou+2VrU58rLUAm/I0+Cd6Ct9f5ZWRL9mE9FDZvFtXIz
lH2PUkpqrr+AvCc279FBLCImikKsEb7YkVRAaIJBxDTpR12zWXh53uAhA94k2U5OAGJH6Mw7Y+F8
KlxrTKv5V5E+SfAFuYQ9uo72vZUEY6NepWHiaLTmYHN+y5IXACBM4wFY04hFAj3G0TMwtwzVTuMh
3NJkfLGXgoxQymxUmOuDnjwNDQVEoy5tTRXLTD7+OZWskFBYWTYvX6caWhgAhcDo1WPFauDINB11
UFCPpswM/Oj7THoH97C4yBWuRWRU6vUZ4O28FnKKSNl6nulnThNp7pD1dm9GWttMWtfq/nc2yxON
pf50FHl0+p2gDxoXOynNsXuzAsieMBbwfEDffLjwiT2KoJZqcrsGY5f9wJgmhmDA/2ZFBu9ZMi9W
1CWryg6yUjo6d+RUDrZlBw+9Jv5JA5SgGzNlIkuSKNOrTNgSpXSL6UgrcGUQbBLG9JQlA8JIIDax
n87ckziMM6TmQx00qfg+OXPxay7e07Ail3i/hsx4CU+s5e59YWQZPP5hXZDHs23ITUdRaNazgXUL
6pbRdPOybtqw0N115nwrzbdZekUTGbiMUMPhxQqy9F0tLO+BFHa1kX+hSnEhZRsNzMlr6zw7JYOB
xN/+5gYNUZdQlORqniD+ziq4zf4nsSTjj1vE6V/7CZFWmQidsTnS4JEMWOb0MX8iLW3CHFTw5YeW
3QteOABQdcJwySu77EYEoNk9QhtSI4bcaGL2j76FySoJmTuM4QNvEEXAGJjIWiTwVu4XiGnjMb/C
97jceAEBF7OJh97GGM7b3JL1Cs+jyowEv5cnVmkMY5NbNm2ymOsSdoyIiR/aJLzGOPCCf+J3yL3e
kok4vt3MKCzySml0pdT0OSL/+lzgfEDNPgr0udds4iZE6f1orPTnYc2GhVuQ0EK9EP89YuPZcX/i
y/ltymn8/dVMc9mfp0Ot5K11IwqGGybldwgc/CRb0dI4XCcxmZRRQILE0edcFGkARW4r+BD7EoJQ
n944uq59v+UZ2vSYaoBwPUq1sxBZHzMmXDQi+eqOYJd2IVZTgZqx3rVmjyAZVEYJUGySZPW89rBh
CNtDrbiiYW3tOrryKMpcsFNCVnBkTM80SysoI1Y/O0MYkJ487rY8hv6PahThn5Q+cwXdaEKsmiqA
Y7mFxM5zQD1y0glMfOx+gkvUUO6DqZEFNGi8AVQx95Z6oDfsDF1Zw1y5MZBIwMvtsCLaoNTAD+fz
xpMREHFKGjr5rtWxgBQtbK+ULu5uTr1crJ1j7uHUsd7CCYDNtZg7+/G9303GIwRK2U/7kRUDudtq
TUPDc+3Y9NVW1fdJq3h70ZjVdQjzMFlPAAGg2RHRlvSsxHNVDa4WJxazdMVrZrb3WlA+h5VU98tg
KDMZQpTgixvfQ5xoTfdctY0sxpXzxMxcZtPLbufE9ew4CLj7ssJS9B2ym9MeafwWWAej5jh3MBwL
CATLzZVWBU2GoXAikw0iuzkV5Ohf8XykP94Q7jaQx6Dy/xRLZzYWfOqs0NEgIXNmT2TOADTXDAEH
azzyesRIcRzrTn3hvRCiIgFd6u32wbLFqt/eKswJ22IICyotSvR+RH1J4aUDL9xGvamOw/HN4vJJ
m3+/3ZMnzPyhPq1QXUad4xbTjatU8UWuf/NwvfN4EwQvBhscyneswOaNFD6zmiPpaRkplvRyAxk2
3kcEp3AEVHK5y0eEpsppuUflEe4Mtn9xc9GDsqhF7rOqRTHAiYy4CLO4ic8PArXTLKEk6AIE+FiT
oLfIA8/lRu+biO6/o7DAwmCjvYuPKn56J6y4FdZev5urcH+o2qn1MkfNhEQWsn2i5qojoPrTnbAl
NxRYkzgY7+4B6EhP/ekDBnEvcgjSit8Ql2tK5zue0AwLfe+y9z9V2yTqAXWKYseiFmq6OQvWBlgw
JvLfafBYwKU2seh2bGOc12nUQ/i+zfug3XGVlmMtOmsm6rTMDTbYPvI71nGgwAeFo2t32rV2voVY
LLPtsXBLsHhGWGqHQnk/fmRc9WLYx4q+auAdxLt34qHHRoGrbstDMFiYIkvM+IxloP3lg/+Dqb/r
4FLRIt1o59osEiXfZei24ne331HJwbj3rf8ZYiajY6JuYraVt1mR5x611+jR9gczSiW0fNq7pfnE
d3JlPDL35+00DmnXKt8h7uiGPQgJNxX1GsGmJTYqpRvfvr1bEy1j1NrJKU7fZzLQ2hx7RgZ6YmMJ
lRvTXAC/SRs+htchFY8gcv2WuPfliuTFY281pqzcSXi8kDb9mJ34OB7miNT8jcAT6VBaMFKdbGgD
0k7e1i0WZkUmzJotnajk2tB/73dbFxkNyTUFC26KbQ2saF2tTHFtLgm+kzYE3GUzGLW1Da7kbN2f
BG/iqG1rKA9smoIupwQfwTPPBy6xBdE4lx5FOuLhNlRYA5s5O59eWwZ+LpITN3RbOiZUlaaew9tg
r8Lcy2sSeSYzPjVvNzJKTw73bqVfV5JrTXuPASP56JO7jhX4coSM7bVi4iExZF+omn8VZ0pe4Qfk
9+3hVgs6wnl7VrhfgBKMH9OANzmHci4iD6Rsb0Yma3umfaCf3badTNN1a/ugFmgK8Lg+9BZ2SreB
t52UDKrr+vhJnccMSExQ3GqlmRT6AQ5uz5teS5vNjs+KLLz3cHfha8A9b8VD99ByOWFICb7rLQIm
et4d8mcXqnAP+aFieLWUBIb3Laq2Qs8MM43pZvWccx4/vja2KQl3w4J4N4g8sRUxD/C1RtcWgn5+
i4XQM/fUGd8pcSXLtamxZBT/pNX5YP5QyRhkkKJHydXTBpLOfBg7yYkw+VGuIOTlBa9eyRuUEXCR
TURqIWTdHlh0etFP0BZK0viojAA46e2Sj5ZSUF6ae6IM+792NEikvFw4JCs2316D8apoZCmjndXh
N0vjhxU5qth+/gXjT21eVr63GIgUrvr0fzbrLn/dVj2YyuV1szn3QoIe3fsidXZbaNaxQ98Ffx2V
b8M3r2d8+jqL7aORyfToLVHon+cZo6905M46JM84mWyw3g8uC75Q6kSmedoyLqnxjA1m//5gPBOk
8P/9tC59LtGyoLFOsC6SdgNjQ2FXm34BgGh0hBD/hkGbiWCUV1hFNESAC72MKauWypzyKaLWBVZf
IlfPYgTW07RjgLvyxdAHr6ArrfiEpCq8NKkwk8lpgcnEyB070f97/Ug+zLtjzRwCB+zZ5d65IEqk
VmMfTSPJTa6xR6UmeeZ8706XXERIkNVPr7qHyv0Tk2Ufwv4VxpOwtU62QCrWIunleuPDsCH/MGaj
vSku9l6qoj2G0MD2Yo5knopXhOFpRRiouMCVFw6C1a/BwE8zFxSZqzUP3740NlzWHB7K8r674YzQ
/9i8ob6E6Z7jRyZXd/3tu+scwG8r4ZyWMJZO7mZS/MwjTmMKOpgCYEgqGSNRLMSpAcN/0p9oD9TO
bTyeHoH5DQkkNgJmXgz/Yyj/jJqWOMj9XnsYDiNLoKZW2HPqW3Fq5dzb0x2mgVBwFInkyer8O8Ac
4eEsy4IKT/xxpVmYo4FJ/IelNBprnVdhJyWbZr5FAjB2Qy4fQOIR6mXNynvfptqpr3JcFpQQGxBU
yaoqbnwU0QDtmqQ/uZr10cqyMiJVfwPYDZity3YUx75Cm8Yi1MFAds5TplkS4ANOAPXUW0cCh+PB
x+gOTgbXQ5jYF1U3rUTL6hnaAXZ5ytvI9I8CX38ZCj00s6MHeZewDmJXwBGAX/KabQ3sNpeYdCMU
tpzg9FcRtRGqdd84nl3qTxmlqGN1TbjfuLrKMDAGlEz3q3pmqAn6X3Wco9MhafJWsAQIS0b2GVgC
7pH1kjDI9Kiyv1rq7XawU7DRyoJK8Y0pllTRL2UhZ7LFT1fvD9WGawGCJOupgofTXVEV0D/J1IqV
YSQQf5dgH1HsVOk0j8h8F3sFlRS1YzK0gc7aPI9hRyDxnfvdpP5JJhoKjkOYIYJpugLITcf9mc/4
0pHOtWjc/Fq0hJG3izq2L1WZbJSHeQzzzXKpeVMEBb4jv5DBv2GK2dPN2iBF9QkAi2yyu6GxQJ00
bF0KnPHmj6w1wxm2N/8hBf2K2a3dXhvQvn6ca/1EUprpBCBS5nbHRUiEUqOKJFYRbVwT0wKF+qDp
5zfWZSal4d4HWVWSt/eX0DxO95VgP3moXZbvumusc0rPUrtX62SLSItcaHQqAyM4MX7IoYkS7XYG
445BjqE2/Al1wjRpfCIquSbQ69AUGW20n8+lYytt8MwuFJayU8Thb82DjOCEsRBU7XVUuT7PMbVr
SFkoUQ3OMGebgJRY7p+yvKlmijGLhIL1igxMvrPvZk9vl276OxZZir1AvuF1opFG0EprL7tCmHBs
/IG7NwqqYqxWzQ1pQqFo/vg9xaQqB8Bt6S7o1RhcyfXJMreOsP62s6LxZF6XhFwKx8GpA9UPj9wW
yo9IDjC0/3Unlzn0whxclW/eMqF46436sYhDRYXGDhek6OGvjk9taP2Mk7Oi5socH2OYVrK6hAc1
s7bcFn6NqU7JZpvP4+Y70UeZZj0XL0SThaeUiHZbcrirNG01/BMrrjM59nKsXbHS1fWkSQRrhmMq
AFNdg7eKGbZfn0QjnxNP+U1QdJpkHpUGTEDZjiinWW8kkwQSMbcpwf1HCAro1CAS/3euzW7TXqhO
DTMwBXZlbVhnaCe9I6NWQMtDuSBOKFfXu+xSuHrWDYjcrMcnDhCQe65mG4bk08J4SqmbXx9gEZLY
5lH280bWs28h1Hka3qbIkGWtU0S2X1pCov1zTTf5U2MCOuKBYPjs5fGCHy0m+mpG3r7PRCj8l+VZ
euKMHabX4bvFrIuddi0KRsH5TUOpDbQM1p75PpZbAxbVGj+uuswytsHaeSrsjwhYRVD6WpPiAfWT
O0NiQS+QDkcXrICdgjFq9/vKs7GjP6IeMcHmWqU+ZPNtRIShDJQURNeii3HXj8RjrOfvI0wPdj3m
BysI9EE5fvxqaBqebc8Kb7Ezqqz4CikwMMAB3PlkmzWu7mlSB1SvVMFwtIAmjLj+dhMx5xW1Oz+F
lWeInWlP2xSK93JpbiEWNsz3PmpDtke4VB5abK5ATzZh4m7rxoza/DhaIInkn2RzBHnSXXlZt4Va
rcUGkr7JjbSpnbvOo2YvJYmsL9GXFPoibqsszXZFbb75KphYtFHDKmPBx7oUUTkO8Xmv4MQo7tmK
l7LfucF6/n/jpT2Q+vV1bBkcMVfD7u+5eJEX7BOhNcKQnjjLxp8Y3JSwOhwwiouoIkEigbUiJJU7
lNwtoe5uy7OY0YViZd1h0ykfn7vGez3zodWQaGPeml0PiJyrz1QLYJ4dwUKAG94yRjNzQNtKRlud
sSXgkhUNR8lmD1bZqU4kUJ9PvZj3A/kNvX9IMAVssjn8qhMVYQe/6ias+8VYukeWMMLnVZAq4VSo
jCxu0bSH5gvm658Yg2OFYII+eBe4MZgi92S9+jfSbYcmhS0A3Tr2tZbo9CNH0mryjcEgdgzPveVV
r6CWgn3EGTZl6w+0m0/R3s+uRszdP3SWN6WkSDqtiuoZIrYgI9fmFZLpOAkjxUM/YWpg8O/if5uV
d/9NaSBfalh6lszKqCbX6TKmUduDW+fJlUrCxg6IzdPrq4a/T6jIpyhL5nsM0thLuphbQwlgg9ij
hpX9IAeg6VzvRMFdcTeKmMN8jPdbKV+SIPiQKINuKnss9KrKggk4vw6gsSB76lz/B8PPQCYOchH6
0afU8TnlmjkZdXO8qDhwr2/bzYq79G4zJBK283ay9VtoiNRC01zLfVThukNkDQzkHf0H0txJme+G
Ci0Z+L3HAQt3AsZjuOSJCVPNx0Pa8EQufauJ79BFm4sHUKAtRpyGbK+VGP1YsYculxQMweW7tepq
FECe0+1lLEuPu1s1KsGhD3eLtnHX2n+7GveGLYVNrNIW0yH9Yh2oKImufolNEu3Ml9qZMNQF1eLh
rhJC8sCPlFtPod8QhWszxd7x1c5fooiWEt7nCOAETRLffspvAVmPBdFxhNn5J9mFWhyTMehTOncu
uI3RQ4jLB2OpEv1tru2uMBocPrViXR1Z3nk9/Bkamf+MKcXNVhzox8Yc0Yt94wQwyheB42+aKChU
Ks3Ouq1RmG96Bx2KMZQAw2n8D6ZXGB5beRW6z76dziVbGY5l335CpruEitcrpvzoqIaj8oPUy4BV
m/+IXEDZ8Lx8Mq0eFO9WsCvJm1KtrQTQ3drlxtsCKk+T7XD+BYA8u36YZBKFWq6GVBSsbDUMbEuR
yj6SAhoqehdIGeAKMfVmBRWMUUeVCL7NhChdvmQEVrhmVMn96tcIJERyWt7jx3szOPVR2XQ0hL1o
lQv4iPK0jXN4GG3aVx3Cd3lEXfbgcvyuFN3yhn0sTZ68swDd2siN2Q3z5bzp87Yy2rfCbb3cxsyF
768XyKr7DjmS+qAF3rhJZHnWiy1Qdc5MCpOlFEKgiPoU5RBN3NLjhCPfJChZxyqS0uRdJunmItFL
ZBhzCs5iCpEIFq46XqOYw8OlttOd+VGAMu948APXs+NlNK2O0f0XG/1MmXz6GFUwtFb6PmEoNOkt
hF0ErcG2C8dZXtZDI9GFjz6a/kDsbbf08K7Ie98LPnuUFb1aRa4wxrE2c7iGtsbmEjXkW8Lj2Hcv
VSU8+1iJAnAhbLWrVu7kIgZHD/q8n53+vtsm/k77OwSC7Z40fYWsY54ISUWTWxud2XNxXHOKjo8O
EYGcQyKm++HNEYGFDXrqTGQ4+P61RXwqDEWrqgV/gGT6It2zZ8v6pjgz2aMqsSTVM6TfqCxPDwU8
aPTJZWlBjwh32cYJJTViy8w9rF352e95grDblB5c1yJNnLGE644Rvj+CnuMHjKudUcCdBUJ5hvpY
O6XGcu/pyliGliY4qJh1RfTFgkPI7TmjJPiXDgbckEDKm/oNLI5saD14/TCUpyVEaq8mH0BYqP93
6n9cvqnk0nAGNJ8EW13pQXXn+CPfPyzpuKFAlb8Xz++t7SJ2OIR02D3HwYQ30YI37pUZ5S+cSTAW
SOMrbkqRLGkxZ0rZ/hzEc9MhJgr6JBeENktHeRBaVXNFB43G467f45MhNCaGWRXEVI/Gw5jcuGu1
STiMDln+JZCio9M7nXEfBfyMI8MdH8OynEcinSKpoNV7f+IKD5siBcKEFl1Qil8n7tlfXmqMMDuN
vv+wW/aNLJYb3jyHcqZnnArdd+GJ52FZpVm2TW2S3HBNbWCtmGga/uiSZ0yRTK38R4N3Cc9pqtgj
8byl11faKZhoJEcLViypz40cgvf+wP6mpyyq7ITGclR6Nr92A8pwPmAX3n1KXThdtXaFoWstCj4C
D710Xyb60HXAMSnGUtdRh0rtgNH5FyNJr3iC0EKyoBP3wnPScznmEQA+ASOWEh+1moK1XH1ypi+g
HRYEme+7diLv3cJxVsg48IX5KCEsA7W9w7WFgP6lCrJLv2cYpI+AFe/8x46bJDm4kBRz4zE+W1dX
1Mqz2//+EgM8R4l9GivrUfzF8SHmZ2OigsAikmzF0oTD4y88vQjUMK+mGNdxNuOZjwxsMrbnMNGi
LQxatVvVB1NjplZ702/GijzLpypt5TOOpntfBOtvYFDxZhIPMSeYwyFsEN6rAhGwbEblTbQ8WByy
xcJFf6dvEEbQf1jiiKCinW16mWIrVKD49Ywafkn1XQqWGR3zsBhyeg6GUypPqSpHOD3ThLSxglfK
MsZ3kk65V+Q2u485OazCfbQjZD8AQkzVYHrL9YSZjHaXblNqci+qif1McUhudytbaOOliUOWG4Ea
4oQBDeOcVWqtTZfevyx+L44CHz7bmLqz6yrYoxq+Qd4OnsdiqepHjHB0RwJ7wDkfkhA6MDp2UxwK
Q5D46rkShNiMbdLsYMctsCEoscVEotf4IITsWoJZU/uIaSF3v6zsGbqZCtI3ihpXlJODeC3oUP4o
3jt2LDkVWUgTVucpNsAAlovC5g3Gcbgg+8Hjpa6phla83Cb01Zf4b+/+tTaXKA6YdsLgLAXpIMIb
SUQGdcwwRM8Jby7QK6JGnZzA8Nn3VbN6G/WriUixvqYuQQJ9CywB2PLsxctTbC7vB1wPmepSMfm/
cLJJsqSS3wKaFY83yYeHRdpHfioRFzPLM+aAzM/FxUhXbwhuMlUfxjqDLyPP+32ZHqwL2qH3VVSg
f03z0ovGMzW1/PN1jrA/NSp3hBA8Y0ToQ/jAJDR8MzrIuFV5x+0ivgtnCHpQXbo01mVeuQj9i6Za
i+5xryvetv5VomYmsgyyQJ8UkBCHK4cIJvD/p36wZwk/CXW2YzECt+vqmOBG9QKOtIg6EB+QFJq1
SFLXxBF5Kbe0Z3/I9rkHXPOropN+I0RSnfue8usx4a04tJ0xI0DB6FpO0NO4xp5ei7kFSnqryoFE
lv2SytzqVDeGfJtMzieSxrnV9nB9efCNSZ3PPdKvoxEjYi3FF7GFFDUjiE/dEQzrgxwQoj5BWa4/
lEKn+2oG6Sh7fok3E5mTTn6exr6svbRCjOPcwcQX81Atkxq3U1/ixpwPZadoeC5XtrlLkMJm4bNL
3/fg0IBzq5BTy3H7eQpUo4VFgPs4jmEKIbkxA8SyNsbUPysJlHwOnlOlWhM0xsPuOTEF2KG6uaya
8yMRBQRCkMqMnrCPbpjUVvX4W0+oJ8ZUcxENBAGlQa40tjwz3T7f+PmjBNBpeiFuIgn1IocKUSUu
7uhZI5ILPL2pxJj7o24KBbjBYGwkareEmHU6oe4STZjrDbfiBM6L0gNqYBmTOgAidkQez0B3Y4vN
7ol1JMi5K46XElzywiUxM6BmAXluVxiV1CjQ5OhNPntHM7UKkG6ObOLrJhL01sLnBUn/ePsJCAWe
mzppf5hRwHzia117PkoAvq5BaBEYV2dIhwRrB6nxMi/qoNpwdqw/g4Br6B+bOEVLUMcttlvXjlnT
rWLQR8VyhrTgvCvaIgJWKfwL7xGAncesE+YoUkn/cpH++ylsVOgw5HAm46LsIMB4Ae6yejSdIMx/
6NjIL5IOtlRyASkZAAifOdzQnDDN3bNh8QH6IBKsi7brJnWwdH46AKIgStB1HjY/J4AwITn+h3up
ZMLwJs/HCc6yv+u1lNz8ZRol0uvp7QZcltcxvdCIy/RdFAAUs7XigbsAXTAdGbncsftbiDTMXSwK
gl602gWGaEaA4xNbhk32lhKJm6mtdlGEX26IXgaBP72lv+yO0XS1F1Pqm4otHl8LPse7vr9gAQrn
vreYDpUEJZYBBh/PcSO+zOVhJsbh5h+K/U4MJJ55TMGabqbmBNSucTueWkX9rpr4kpH/ONqZvejg
2w/RorHQG3x4kCZNaTr3NZmqBz4DQtcAHzspvv9N1zpAaFU/H6YyRvZwHUP5Ck9N88U7IhR1iWvs
rzFsbrz6s/JebI+uLsaz6fEACS+fLEZ+8fzi7KaTWWHvA6Ow+mrNKfEQaE7fzyaCD5BMGNO9bSEI
869J0iA2jo/n/VSnNjgzsQAUVFgEOLoOGrtlhUfcqtXxeYGAjQVcoziRpOWIJJB4xqjMAXUhjXB3
t3j/v4bDMdfXKnffO3PHzU/KC0FQ5LI+v53FmOiNq09lB39972ZV/FKaKwUG1WmsdUf/gCafk6+h
XPToqUBccDZMQNBKHtGAA/O0S5kwIrhG3ZUyAg39HgZZ4LG45DoWcMRjL6HWD8KwyusIkA739YBM
6CZDNw/rLOcGNI0MC/bwDdcwz/sz9kC50vAkGvxxU2DPz9RPQEmgPhW1khYzRsZQrIJepgXWaHvg
bOyl08Rh/TU0kBETc48uNf/a8QPhXycFryoRJ5cPG6dc5PFwrNOXz63qFD3jDYJCgejulJlzUXzI
P3UvUnyFFH7ti/hGtVNhYsJA4cmSEXhG4hTZ+uVSqE1Wq7mvlnOjhmro/pthQ1nvXWTk6sV1etT2
DCNCzf599kEBSm2Mvq/KC4CrlQmqC9WgDJVRKQq2EbDc0lxgS9RIn+yV+TGZWsQr19J2zfnlTr73
XfpRh5iuJAejiAQ34E0TnqTqjx6QujkL+G5foA0iLceV2v81W8X7OEpL5UAviWIZnxBiPXPzJ+Ru
+ZPCvk8nzZ2yZtvqunudeAeIYV3m1FPSoeAVdBGeAQXkHbT5nMCa2C5WmLZS2hwd8wANqXib5rlb
cfz+m9Cgr7q3lFApLZTS6Dify+7PkOawJZ9TXqeh5hOTOXIntH6J/hMiP9XNSbhPU3KFvdrlpTaZ
2bAdc6jv17ICV/Z0pyzwgfKVdIFkJWll/4y2jEjzVfjTMVsTtX+B35a9GvC/pq+GoHLqUA+p0DU0
2a56E/uiyWiUU8iNtNMpUhHjUi4GwpEtEZwOH1rqLDnePiHYYg4tpoN9hvVKc1rhpppAjbS0Meb1
rI5sRwnOaJH50SpQsytKu7GvhFsP1caPgXSb2Jz31Nosx2oAuodfo7iYBWILP7bOCE7JtD0BdHXq
xkk0saYEv7hTLgkzZumSHg2Udpd2hjmLOOfie2e68pzHhIUx9Ws9DXXnief2wH+H9k4x6n795Dvp
YxQlZ2KM7jO20XHT2zqDmQsNUp9QDKQnPTdPdEqEslFxWk4AwWRJSV0vCDl3hrA4gVWQfv11u0KH
zyRa+ZqRlpcS4H7aQCjNW4j+qoOGd2Ejfi+Cc8onwFqqWo+A+o6FDldVYXZVzCMl9etbl0PSd6si
NBe551yKFIFnwEOfixbFaeavvFaFGVWHEBIS3dHZ3OGsDHWX86D/KMkV85G0tMyx7HnGyuDBn2+y
M0CyM3ZjEPZr1i5+uXQ1xg2twuyhEWJGKj5Kq2tQMFSL+59A635UmtUS5ELkF2gaarRRbDFo47/a
Ja94pPcnkuqq1CeWmACoSdGvXi4TOGI/GFPb0RgZj8okKBPynJwKL0nkyubCXOvlez0DV9ahGDpS
VNRWNNI1zRYe7s+tVBx3/nJPxreZrlBSwh44HvJfdYZi6bvIG28z9xqitvYGHycGD6km26azd0Fa
ehbLeSw2C4rn1nFGuEPWtwYXcRZo69xcS7VeSZhbPB5WCTEyuhTzA/f5Uk4MIXzAHr+y7MEJ1ARW
3P202tcHek/8qdQbIgoPj9w9/aP4gtAVvFfzl6xRWtYUXDfD9DwPKblybhezW1CH/Xel6Qka/At1
f8OkLW6hY9p9wjk81/QdhmIC4RCeRZi20aIg2EexKwq8vyOJv5Hy2bFzvBwtoZSZsboOodLe85Hb
yX6SJOtnGN4YFkiSmxxVpgsDSzxZ7O6DxKU5TLCFnf/614VYIQE7ir0Xi5BYafPw0Oh4sKcOqBax
il9LVCiUZOFx/+jgNoBhSHc7AH2zUP8mZpOnuS8rw48vzq82nuRE9K3kMjthp1NLwPvPI9TNGim9
DfKSR5y6Mt2y5U/sq+GwgF98xOnr3gWyXS6nCm/z2txGWyvwsC9pivRHbtiTxSvMoel6xE/0l2v0
h6CkJ19tMbploIjG6opy5DVqn6XVmJp/vyhfMW2A6ymMaB0mbIUL/EHrTQg0nhK9ACLUPId2h22h
8alw9fk0IkPZpaNcRutplZrJHki8FaqnuvDvUvPqL51mDJywdUTz12zOMmVkXer/7sKAdaBk2ZPJ
vlNxQgqdr+VzrDwrg0fYib0bSRD8vPUwjpI/TnBxFp2z2hstAOeQKKN/Y0nqU5lLKfRfIENc9BNI
dj5gj/6Ghoe4vRPXm62mNuy8lrnqX7XBmpYh3P9f4oJ/c16jy8H5WpE03y3dbRkmjMnqEca6MYtJ
XRPakhqCDB6dTuqI2ZChZ2HhoD+RwVoYwTPR+FtjtJg21CecHEd3N3SU2ktDdtut6YVBjl7yncYv
g2Nm0G+DF3DfBrqXNjZdnRdbz2+2FOLundLZ+Vz+BEr0ciNpHrrLnMpwJhILw13shhfeGTYS7Dvt
kLxWHNE1xo4WHCvrtFiSPSPxU35jpwVD9RsGwiKg5vBLHb7SzzLJRjBV4g4AmkzqIhqh+dl6E9H1
rzzoqqfDB/AtqrT+VRuWjH5Fw8/knx62UjR98q/+tz6xmZF37+plneHOwIoliBXrz41TgRwKARAV
2++EZBzQIx5kwlQ26CYCSFbrhC1ata2en/3c862Hhvnx9e6vuifdSdiTlc2/9bMk3+qdzya9tFDC
R5ESVi1e3khE177fvceLsewga6hk+LdOWUkMHmxVKpwTfMplfB5oR5QR0YnqDnpGJNnt49rtJLVb
6QyZrLCpC+ipR1E0nn6m/SbzN9OUKM/Zo4p6hdsqQYxsYX5B33L9urPWqVuKaPVPV46XHzbty8ZS
o1y0h/fd6gKIKRtsuD2yowkQwyGJmQFWZrtsNusSiNdqMPZLMdcJAd/FVcwPdzBWj/jzgXJXS25K
ZwMDl5TllLlZ2ttOVPP4f8xMnRW+/XG9n9FUHJPN4SCD9O1WlBEeMtByy6iACGIvFzWw08UygJBp
GgzohBTGkY1qghH+6TKRml65nflnDEbUdq8GKgkOmYsddQIJ+fjaLnA3/uIPzHBIEv7KovHK3L0H
jPVeXOz9MlKPWuN0XdPHA2dgVnt9uOYdPrsA0IzPAn+/zrMKR35ZyPJKOoQu4P76gkgDLJAcWCQ4
OViKk+TBJX7jsiDH3WwlTUrH5J30IlTD8X5tSwQr+yD+PevvA3CAWEo9gqgQRv52XLUN4vTpxNe0
tLOZSy8dFNXhciAuk0Rl0cyTRB90ZBRllxUXncDful9etogYCqN18KUZHUEJaTqf0nSgK31lnrFT
juEcjBzGVtrGKchsUln43QXSM6+95zaM8Nm3SUGyY37h/p49mCFySem4IX3iJ7LRieCy1qeUXT+m
ZCNA8L6gX9xCDzZQc53QZtwMh7SmXqviFDWKNpFosXflpndUEKJw/w2x94sRAOCNyg9t+zq8m0W6
7htGXe5iKd3dPIk+Uj0J8JX1gCpGuSU+erOMQTDfduzK1niK8iJg99KkyNKyFE/nANync0TKNa5/
b47iyHMiNaEMQ1bm8gUMf/qJdXcrE1RjBURGVS/7fVhq5cDvfspX1dRkNOTeiLB4I2AgwBQCUgd7
hP74HTscor2R/VKnWzMwdHrkQ/G3AZ7bDjq9uG11LgMQmfHv+XwuZPSQS7VZxOUsgC+bTonBdAgK
At/AkDJ/B00ij6MilImCh5MftF22MYhKNHw/e+JKWHTSszh7WXs47idPRo/+jfD3SE89wNZ2FaHp
H5T8/s023VDsiHVn3jlOL7lI0ww6LZ1v6+wWh4BM6ZQmIE4hcODbtONt+WU5ObQFj7E0RkSQ7mFE
kMoWbH3cn3ZpsdCU1Val28Pd2eo1WsXc/C/b2f4hOGjqrFBbu7NNJXKzl7JdRJq1mS3lKo3QoHp6
NnLvNfLkZMkPzOc5I930R7BEUepffciuqg/CD/ev6aRLrp60llKSierY3lCqUpkSGWYZihNLGyfn
gFv1Q1Dh2rqRWDja7ZphFYNGH7YMw/Lko9skNtIbC1WfGiIieX6QmlmPPksOUT5qWf+odbepuV8P
zgvWE4LGcDGkWDAvUPIlpjEInQZC0SkUDCgX3mW7BfUPwHfahnJKeR1aGX4SKLCIvZbvIAlBC0Vs
G7O8EX1ebt9XWypKGdqOOScFLecM86QtWHZk3Rprqvvy6ROqZfJoKzJtOlvg08zQo6sypv5PGBJw
Pe6RmG74hIlIxj0fWxdK92tmCd3OJSJOGa81wlCZo4+iiUwsLUU6hwDNwLdko7HgrRtf9esa2o4s
JDSIGuqYlfSOU6zKz3oSxJmIGJyqQP4gVDX6FvpXndNNg/mth5Xcm9Mo1qfaNadk1aCYo3rXkjBW
1XIq1GBiR0Js9HbYdDCU3MpTd6ZF/ueiuzMiSUyiThT5yX4f9EcMQFgO0tz0iTXnSzELNgrwSYBh
tFQMYs+YASX+QGeopN557hMy8LJDvHr1Bk1+whwpVX3YUAvWBouyUdwvcHH3yLs6OoLFbiYNufIn
y/mbFKht8GctXOZv9yC4SXH7R4jQzx/DAjUttUO3FnxrYKQy75ju7lZrg7QrAMRMggUkCMqbe0wp
ST75wizrUZDkfPLe3ALAVrmH2KEAx10rhoa7hwjCboPTn4LCu3OvdOrw7zTlshoCPBwI/VcDbC4t
4YeBs2Ss5jsWrfZeWNhWWn8Eq30CKLCEU/L8wKXinfVcokjLE5+LayGDsZce38j8njd/Ai8OQxcI
z8hVRjKrqujYPgZ0jjQAI2fiDZibI1+ZNsLAO88/PDQuH1wHhegLoKajpwnbQ9MHZzudE0m6ytfu
XlAPP8KDf+mOm5FMCa14XkeHTPSHPDK+eY8MPDEwcHGk88ijEYoQdQqstNxMebI5Zqj6crvAdEH2
SI1b7hDRRUR9/5keCpbGA8LZw0scaJXzbNE6i/8kzC3SY2blYZW9pqu//WP5gOn8B6KNxMdkF3eO
enuoUmcW1Es4iFZyQJxay3aLMatd/jP/EilBW3ShuQ2VMBRqt3l0Cjhk1iJ2GyU3l53VrZeuuDWv
EWnRbIwMe8PcM5JogoWoH7dVnOmW2E8DSoD9Ga9N3iHnd393z4WJbmQnOnw/2vwvX4FCzIoEJEpd
qz6LOLSYdMtHM3eFk2H07uv6c3iqZyTNQrtzwlh1jYTZH3WVffY4d3VM1CDUbN0T3HIEPVejlw4Z
3wlmsY58wo36jZVGATSsiArNmD7Cyt9mc2X4d7smdIOPvNcGcSuqaTp55r6ZWEScTOD4c8Sq6P8r
J/0R0idEKoabP6IAEyy0pMF6UXbgHztZ74vCp9caUvADhkMUsqKTi1Ch5iESwDzZeOvjW5uwPDKF
VjLu3nOIJy3nS1GIWe+i76wuo/ztyZGNyEmwVT/oFzuwbyyLSZfkvn4XE5ROev448173/xKBxoSZ
pngbBKnmib87J+g70iZ2B/VM1vklziEJRYabX0U+AlZXSWFzuQBGQeUi/FjXe7ELCQpBo88VOVKH
Mp8a5WT7RL8H8FlP3wi9dCvwNxTnrL+5DIGLTwv7v0UFII4dyeaR3eLf+nqqV2AXjT51qIsouuTE
YYbqpZsBqE1QulR1X8ThKZFWYZfuaKjc3cCVZFA9VIbifEWrbsrlwwoLlSdqeYxhjIPQGB5ukN75
08EFVCrgFtIN/pA/oPTQLN25XmHuwP9fKOgQilItuPuwWgf6BLfwCPxL3PBqDhZtaTp+sqdNW+Fq
sXpdVnW/7Ig7cvA/i1cCTl5bDIdbKEsp9yoWTiu7lqBG5B71lF9rFTiaacfwygIONjehkLRLe0Cx
h34hwxJFl9XaT6Ay0FiZr2QEpj3UyqcWKlu7Ln4J4QHWo39FS4yMhLoyn0vQZPVgsQ8JqRjVBV4D
tlTRifjW0ssv3G10A5P5gHD6MaK3wJeQ7R/VIc+gMxFdOQmHtirhRKYOyfJpU0kCmD/nlq6iudg3
JFEODBbIgfLPQF7/bpVQSgG7Yf3UaQ0rCucpuWxXhCFSzQZC2WqGGc2HyUblPwzRZO4xXSmGBCCw
hChTgHHha5W8zwlMq6LIBOQeU7QshmroJRwq46youB0CLCE1HvYJCJdQy4DYquRKsH4tz1P20X1b
lRAcFZZtKaqkbp7CG/BaXMJEN3kOePUbEvwNMrG0CYG6P6q1bG4Ewae1pOW56209hPqifFe8tVWx
L3W4Ybf3tJaPeMlMGJ1Jdj55/9mUiLhyYHJxmqy8wXdEljKlmMwRLtXR4cAh4m/5yTdwJsU2NHqy
gQ7GG97gFvSZr9jdZ3prRX7Ab2JyTar+8ErusLltVTGf/0k66gSyLBaEfwAu3si/2SIkOgOUgPde
3ryXY4e2V4qOQLhM098iLjSanAI/qrDBUMfWfVtZjDjy3r49khOdz3xrSJPl3kvKEjhoRVFfcgRz
sVzf60iMxPs0WNAGyDw6Nx6RBr2fKgZ7fHurP8SLJr60Y8J5fZAem83mTnkaDKWmHQWRWD3ER3BC
vpGiQhcoHj7Eg6UxY7NIt06KHq9FVjLT8E3sBQpfVvazHWq2MhwWnG0qB99/6Lj3cL/4L7hqPUHr
iDhvdQm8bK7mlM4HHP4KCrrsB3AUpmyl6Ron00huw48ljPDoaffbvaJKuWuS4LWcs+QNjraRTZ2U
WMn4uiJWhkVkNfp+um+qQ5uLvNPDm6hqikrWMoCA1HaSlGjpPDdXlZj5UQq16O4GAvzbVb2467cM
CSRQ1NZTQ79jGXUWic19j5fpuqZ2vYVkC4sO6hR/uHxUh+k9FNFVnrGeS3e1uTOiH3o1nm1hk+We
ljSUklpl6IFpaeI94gkG/k5Pyxl0rPHYkKnYY+Yx7O75ADtKwDXwjK2e7otuwGB+9bcUFxNbCbRe
FDvvhmp7WPN+IcWav1j4hdZBu2cz477eT+u0PXzM08p2ceu721m7ENnDG9dsw7VN8qV4Mj30WhmL
aiBvPCA783++U8RoZn2pcBoBxl89Kz1AgfN6DTIsZQ/vsuZhym/MWwx1+p/bkH6QGuv6TGPd5PCz
U4GyqitRxcHcHOC0lzPQpY3Bz2K2kf2W6PH/j+sGx67uYN5IEXeZdX+MThTHrx1ILTjNj4Jr2pIq
+vK6MKyhWuhVtQSD++qJ4d25jcJCM5Q5p0BoauK3u2K7iiKCAx4veHY4yC2wAKDc/3BikCJweBTT
khVIynjSw1fHE46JJCtVPFrz8K2d0+j3ZVuL6j1ka77XHj6J5lre6lIYt+zGZ77uOEpLrVK2s+j2
KI95SbdxE7dsBZgYseeSY6C5zh6n5JcUkszZW88Nwcx7LkSTlmAIyALTeWpvT1zAn573F7q8vJ8d
RF3Iw8IeS7W1JLfe0do23wJB/j8tYhFrgkvuhZjCcQpk2cDq5rNRZ0xm99B0alXB0ov6t5h2RlSk
t7xzsP4RXXwaMzz0HUHh9cB79HcIQMpG/P9VbzqXVdv/FJmUtv5ULFHA2YVclJZH5YBfUoZ0aQ0h
m8SwitJB9fmw0v43SGF0yx3J3r42fuSUj4qjyO7qh+NoR261iLSzNkd5p71iql2EApT9MO4VnNtv
LwiycdwC7IQT4v2y+QF/wPUe2ZFfPkioZK0of/8xaF0n9rfMLqZtJWmw0zEGro9CjyWuTTokGf0H
PQavBk1xDPUcxSdjQRZTsNE7jfEvpK9SbEqgkIQUzqbQGGI7KnSq6mmS/E1bPPE5+/da5wup+sEc
5XtPioxxCv+qAy6bReckv3hoWZ/egEeYr+/xPdMc6wmvD8SXNRT1aqF9lnzYnklWV/ML0sFMMNDY
a63H++oEnQreW1ix2ZeC8xC9RHaX09T/ZUgd7Jrtm+7X+YjLIzmpVsFq3WBL+oNeQreyLc4gltYH
FnoEd/2p+aw9kK9MBK+V5A6XlduBJo3F/TnPwghT+zs0SlGF/848MFSfQiU+XvzxnmvupOf0U4KK
KByLP+rdNjNFJKQAGkKgu/9F2Psk74VI61kzCG7aN+Y76haUWtDz7hKWoHe0rHcdo6KguHi2aTpH
g1fD/O6Y1gF7B7ID1JzxqcV089j7RjW3Ljd5RV0Ni8Sf40lpoCjSqJE/YZJniRj9bFnZmmEsdijd
hAw7cPk3Amb76Vl50OxMi6PlItMAB9Jx7bbHT5fKWM3Jb2FE8AGP0NLNqw1pKXGAHjIK4KNQRA/o
eVG+hw4QKb/oFw3UgSpOvqYiYUtWSSEmiVAWM7xtn1xj1ZPkQ3EyDPffmD2VK/Ih+fWrQCSHULYl
e42pKz4YEknQLIMZ6J5+xhVDR65b0AC1tSsyorvqZ18RQvl7UXYgBLFq+RdK2aICaJdEgdU4Gpc6
UJcQ1aX9k/8Bs6bZk2a1ZSDbT2jA9ham1Z5Yks/DtE6EKPDAuKGQ958PVxsGVDqNZMgCCFp+6PoG
ikwJHISleIzOzlz3vJyyqg2cmxRwsa/6GIGCralnFcg6Ww+vkM2xMbh21MMmCGHB0UYiGiPD1KtD
MTm6cC/TlKjGCN172hSEiqZ5KVgkhAjwdOZ5eGIInEQswpg2w0Z+/J/Duo8BsRNC97kuoQdrUd++
J8Qe4nY8kDtAxXpFKEyddcHjXTxNs2zYr4+4YukRzaeHLDy8+/BWhCNm4fyYkTwRDfzl7HYOxg0h
bbUUX7drHkfWDX8Mh2yyq5ywlNLAsfW3THw+vVL+LsXkgG+aXAXp4EDUupqQAV5qWYPNannuWdm/
EUDRLUyJF7vlVBgl3e3obx97h9Q2pbkkYl28dD9ZkJ1udqTt9sWFCnFson2Zz2xP7gEIcKNAn5D+
ZpWk8DN7xYKyxsKP8Oc07yz1mRzskK9taPD2uBJms0v1Tig45MUUDp04hCs6BX5yfu3s0Q3v0MAx
0EcvAuT2NhWEIRNE42bw7RZIFBmvXSZ/RrRCz2ywQrUbsc+22vO8C5dO1Whu9uo/PKzMF8YW5NV/
WEOPX1qkSpB/R8Gvw2UkO7IGdErl/MppDV8gGG/VEkk0lN8AXBDuwK6ap4rIfGkjtY1hRi2sPowo
aL3n+uAc5AKpGG9Gkyf5QNAKPPN1/Ea8evupkUmnZer0+YzrfHvGmcnwJsqm84NwrHkSUPT/0Ftu
enONyMN9kXcDyNk/S4AQ8a14EyDKkKKu4nOzHQPcR0pmwmLQvFyzusd5HbYkLrLFvr2FVYOLSQAm
avpNJeqeRDfoQJMKct54isW5xA6sXydXBEiiaplX6iNTL7Twm7U3TmkMI5inp+/p51UscBgejHVF
bmJmM0/MKcu7sDTWm08hGYtrZJUoF0rQMz1KldIGBlFGX3Vj6i2mwMTMenVxWGqe9+7xPmyytpOB
5XEmHhlxLcpmKkEX02iO9TWhtlLxzzniS5lmUh+PHq/dCR4LLTR8lWZyNZLu8iyExmerV9F0yPx8
Y5oRFRN2XxO1JAyooivKOhqP2EpYtNuGONkNiqgxc7hyFKQoX5m4vCtLpmaq5z4RZj4vbvNm4hV9
kIP3Enitdw2lgDeDXLb5V172a2kcolwsF+cD8mjx7rBvkfByKRc74qN5RSBJE2u7S6s+yxCJmyVw
E2l0fzZIo5smNUiI2GZPcxvHPg0wlXNpjHvlVBPAYH1x8K4l5VDyZsazuJh1EQIkgZd6n46mHdBX
RRuqS4321BG32wHbB8l6aEH7JLBVk1t78ZSJ+yPgLUlGYOFO4fkP29FdfYPnzdrN2k6+TN01aDO0
EJHiQxJj3qVuySTLOhCItX73ISDUs7TJsDse8mgtY/+8WKczI8laK4CEdqZ//tY/hzw2y66ORd9K
7SXbufjD9WcNeeG0/m+dYYecqhXlYe3AvifKfhsd+i333dOkAEVNL+FZ9Dhi3KaXYIe1OQ8FbqOZ
jyf3E19goZw3JDLTBDOLgPEgR1uW4IERT5Cpf/JFXh7DOnZG0Xw1Y/Kx5zuaPcDpirVdSe/4gGtk
3xaCIN3ZS8KJF8TQ1vRmMg/Waa/VpAmlAqei0yeDsaHAZ9B4BYb0sAZrhol96+EBa/TyTQvBv6uU
VT99j59ewR+eoJGq0ql5xieNNn25tlJ6rfFTl25CTTZO0vmgKzFmNbCDx5XGy4b5S3jvXb8ZumDQ
NhJSK84T/rXAcH6k2+ApOSy3lhWBwgVk/b4GwhuBp+XxgNpn4TdpdtD3zYUSTsvspLwN6LFpiKZG
Feb1XWbrpLF54KzjmvUu9y0eO8yD0/36w7N1sKej5eP5LcmRGlqNyI8mIvHsw7oBcyCk8eAAwEjG
qR9bBTl8ru36HihB9577lSjiaea6fA9l2TDsoLxpn0G2WqMhc5eD1bKktBGwsbM6yQzGEpeNNjcC
NOenrxz4GJqvxgvZWxyrZ28cOdOBlTZ9Mzuu/11FogFpl+Vdmyk5J4lUzs6g4Xqg251e4f4215ad
qvrCn24rtIZFd8C6q8g5ElZOWPU3pXEe5y6apWj6r7COTjP4ULJVpxzEHg6wrSXc0AZgscsbE/j9
hNqr5sgih5tiWw7vF15H1c1l7MfqyMYwVY/VRHx2JYovnr1MmCD4+Bk78qGKsZyoceD0055+zFAK
31N4UA9qrh+gyKqspO/orQNs7FO855ZB73lZz8d5E0p/FanmfhO1KJTzb4xKljfQkH0BH4xqsnqI
HusrZ5irb52Pr3wskmZh3QdrXx9MQGZftlwel/dYGHFOnR54wCRcZfOt6AsjctXrjynhJKmautia
Q+RFgyaP8MNJ94tioNafbVoT2O80lxesWue6/Id/iqdHNLTGTGzg+54qnsxbmgz3vWzPL6lhouoo
WVzcuL+pPQo0AfrtgAJOHMcaGHH34ZFBvRxAusvZMJ9kwvNdH5oXDnAK59sI4103Y2hBUXLh999i
2BzT37DG/kdmxeOQQVSAPD++jSE/M0w5gFuVRFGyzcEATmf2d74GtOsVQrzGROJq1mMGaymD4knS
8rN/A3pbUguH6Gijo9omQ3FxQeKzFtDGyPqG8JMS9bIAUwl3xRsNFafOemNMwQ56PfceEFgnGK+3
GuCwy4eWh/+Et+AgDfj2CaRueR5PU4pr4/c43ZGtMgfgvHAPz7MiURQEZ8hWGxNE9yRG43UoNAPE
o3Ojhr+GJfjEB69qm2ZapOXK10mSR/kQiFHA01VeCzyIIyNGFgJsnPNeCvT8vCkq/KRuhAdI/7iL
WgJ4XHbwIqwUsCW42Btz7QBze5lFCH/EQg/egl9MzTBlnjauLUgGguMfknW5yMSeKQaQ1zGVhYHs
fPMDSWvnxoEf/4hZZC8ONZVPcIWTgnRzYoHPhSqTeKxUvd/hQmm7xRifaFo+o/IIEn7BsPNa3iQj
L2t0trHp+PpfALx7SplpOlpHMY13ce65CL1O/5vmQJYLhpJozyV6eBgDOtRjh/nJuN32ctsNW/97
sQCPNMmAdUunKkOuvTaAUpiuUTSw+i3H4qapZj6u+HtomrA2kHuuz/X/ScqljwqCN2Fq2CRc2wfH
cfvs/e5GRg5/Nf11wWpBoleju9VXuQKHZ3TBdqKjOsQUCorTClBNsbWkoNME6/RdjaKdPMXHxdcq
qp2OHSuxE833M7vMIvQW8GeoaiQ/3qpnrJsWj1zPVegGhRzESDUmOlI/qSrRfUafqGxImPc1Q5F8
q0+YRGVYhTNjtMcZ4hoeWHP43hR/I3kYZ2txlZo+4PKWgJjIGhDjCKJIjG8j4na/pnLe44ohODZ0
fb9XDre9PBaK2pnQTTLcR4BM2ppdPufYyDdP2hERqIKsxbh9bWfNV3ZNV4c1fI00S0i/pA+w2M0q
jA2ScQycXsAEjqy6c8NknADYHsW2zTgUVTW+TBCPvF7X4yEzuf0hWa0gymEbj22Qzjj2PGDYjwCn
JTf2/ZzOvzto6Sv9nYRS7hQDBMO7cPvYcZrYgPunGtGQzHJ/HstGGXuyHVICQ9wjvvKfYm4INV7B
GI51rpGbKi66SpckhszkrfPeK6A6OPsdcLL1LRn0goEoQy2wZ5qJR5SGMIYJl+AUUYWnXxspT0ev
+p3HccS9oBh2owdvcXrk/m2UnfWkpP4tRh+ETFbxIt46+MeYBtgsvZT7n3YiVB7/HvfJDvMgw5i5
5H2szx22oZ1yLXLFSt4thwP11mDwchHbhh7RTZKaRC+XHMrPZ/Wu7t4F18t6CmfjSSlGx0Uh3ubB
r7aYkQDyjnP1SUnNfeghxUwbBwp0+8QH8n11AS1yAMNlfRpNjZKeaiDyMONAhFIQnG8rHNAZAanH
Bf+E8wDSy4cJlomN/waCPlh+NpdwrxGhcnhxFTa3YYG3pXU1JUPeo4vSve+9aSPfI6aFz34iTQfi
JXRM20zKRim2Zls7OCbmSGISiGQmk1AsUFibX2TT3yNBVbjaUKxn5l7dG8UbjeD2Ksk3oX+SSmaj
xM70eAeza56G971L2WfeJYD0RNnZEnnKaoBZ0U8/fMFP7ljG0K+VVBOR7pWg0CUDryTjGC4amNMc
Zpjwjn6gAaXiYqdf80WxvkPQcWINFwx7j8eCylJFBerQKTTPRSX/ldofW5dBk4YdC0MJxhE4dH08
0UQiWxUDhe2Qium3IROLutnAOZr4NZvtxrTvJMG2dA4EoqObD9Ikb//3bJKZBxmVxym0v46T+lkf
kL94KGf34Wxa1jmsqu5cASCdc6jnnjtIZA1n0RJrA62MZpVsdjPvgjv+0rq3NXlK7GaML8dc4oxg
CXZkGtBuv0/a4sw2Fq/5FFTXkrvQbNh558MtEN1aTFMPjZLHDUOMRjBHTNXEWpiqC2/KIJUggRk1
wJcJGjORelUZT1E3YVGRhdSgyx+RwE/0XtVntFJRaEBHPOpd3cur3XUjuv0o9eHVvaXjorPtwQLA
VGP3+7zqleraT+JNynC/sylMXeSejoZOdrjEWsMm0eloJvc8m9vGegrpeqbOqPfamDT207WHSYtb
4Jjfhb5N8IUjOlLNUCO+YW5fbQlt/vmn9G+HLF3FPi3OYJjIFcauOVpCoFmVTA1fJmgLJ0bMid88
DXQd5fjTJT2Sqs6nurs9gihZ5RDGyHa0GhlRWZBQ6Yb0GJnO4CBpSGZGZ0JHQaQWSwIt9UJnMsRU
jsarOcXkeEuwAlY8l2nykUFszQJ74VAz9Ecj3euHNmJu0XCjuXv27W60gNgI/zcq4UXudwvuQpBC
Kct2q4sdVYrenOtsJlGO5YyhjbKiifZpQm7UCDgvgcuBcdU1JHU5kV5Hsi/AAIBDHE/dcXD/HcY1
YJ03AgZWMG8o5+t9it84zuApjGiDh+FerJYZd0G5m1aQmb7eZLc415P7HLP34HcEruvGByx/01yA
O6elKElDbDhl+xbwhwM4rGv5pqhLiAc6LSbTjO/YCyt17wMTishET6VKQAGuc64B/ZgWlrIfbJPB
Vp/gY2EUan/4YcXFnzIFPC+ZLCiOeuu8vJobEaNpnR6AEYn2LsQPR6ReFvnbR1J91t4jsu4vcO/b
HO2k9UtGmRJX9qHaTK6l6dnmWA0FmVYpQ9yb6hbn6HrSd6ab5b112bOwMB0Ohe5UjL0Nt/dXrBo6
1LceJ9iYgxSzAx0FSAyAaV35dQvzqb69UWwPGNWcq55WRZ65LftRjMevI1YNqZt1MlFcHzspS6DE
HvrhmFXZmYIm4mmnqugDTC8SihoorDez1UKql0YL1TG7LVZWOOUdjps+/O2JtqASGpS4BQhk98Br
0OhsQrQkolX1Ai97XqbSUNaU20r+Dv0brYr1TQzfDNQvbotUT2b9F/X0RdOIyxOT5xA4G0NNBJC+
3TWtipTP3scALEYBp8LLSPMzMVsYrUJsr2MuLZC7s5ujqCPeIjseSUrK7snbvS6VfmIPrD+XWQ3+
IM41TEVzoU/bZzwsiG1fdBC5ALbZpOKpzYNhBINJYujilgykrK/Jml3C7XmJBVdYaHePb7V7dLaz
O6s8R/xNjJJ/txpPZWgUd6/Sa2moKOoHsWjO07F/c9f+pPBVIoTDw+TSXG+4qt47Xf872YPNk4tK
jOvrDIoicQosCBSJj3PI4jQztNN9ysnzmd+C3MUuPtsKQyJdEw3PaERCsAAzUwYRFuXBCgOI7LSo
kKbcb9O0xTdZtWGTSNfUdCmnlqK85VXKhJrikKIJ3xe45WvOwVipY3jTqW1eiYlixuKXI++4udLP
UUsn989FLXpGH8I6D9GGcZgpTu0nc7s2AoEsgznZjO/H3CvaFjT5PuhZ1Oj1UP5JjVM3NdBwTEIk
wCHLQ9QWe0vTUXdAF7abQC4kScry5cpV7ZBOSPsDvIXuJ3pkssCp9Ue8UPo+meBsVBDv7YbWAKoV
0ZvXguODO6W4/x4EazclQKZQFkBri5I0aB+N3va0aNlXDeKbec8U163Nbj+kYgjL3N9WvQhlOJzf
nF/ceaKgNsM0aLfcgZsr4io18CUxXBMkQsCmmSKs91ETCKGB4NvMPsSXwwlb/chaR6dhcogctnsA
1gngA9wFz9Z6Eb23oUBvEgezGSn0qqO2tdzUDIWhgQM9NNiibGV010gIPUSu7FXKO5Xk3xmB+bpx
2UvdLa+x7d2hqaQG/965X364yhZBWfHNV7tI9DZovY55qUQ+HMGxdDd5z5kqIP8Fa9qTtq96fxs6
eByEafimo25pe9F4/qpQzTBAQI4NoYi6KQ4t2IhfWtVe7q+KzidjzU5zfbgOBwnQ58vES6iJuukw
FzTcV++f8/Lic5nPaYYqmmIn5fzu7pWC+NJiSuDLrmwAHLpelceCeVMNyg+G9pdqXqrAE7Qnwxpa
Fo0DnIgeGI4n/JyEXUcqowSPiQD7vooihkFrPk1tA/ihGQtg2JYx96yCMgf6wyJHH6JJkiT7L7Nl
SLjCR2PNwPp0Z9QbXQVafsus2XUcRURlDY8Ahtx+2XRDkxMhS0UisWe7Vg3muymNOCf+QPfYWx/F
SswraT/wafcEBmuV4hLAcfxwRBUZ/Ve+COUz7QVOuH96x4w5YSlQ9pwiVSmEv/kFr9eSEY9obN+j
kyDye+CAoLs+ItweDQHfVaFJ5m0/lSPCtq4cl9dKO1iB/N/WvFJTAe1NUZtIpuMyT8ubVHwtHktQ
Y8jBS9gMpMEMDzQqjNW+AIaXD4CKhm4QXXEH99m3AHkcMgaZu/k4v01hq9BM80Uk0SgmG6tCUOrM
PF6qVrJv+lCxXMc1emVIekdmQjL307tLgqiuLUrjKvpG5Vf62tICK6kfOT8xraNbZIsjKmfonFBh
MVbezsP5bP/G0HioCnOEs07B/PLDHPSoUdSoCWeFzC+nGPwZWIs+I/rXFhwADs13Xib6vt1XwoGH
YMAtx4m0luHBeHhnfFZ5zMRBcaw1hyrwk3ELR/eiAwEVkD3oyiuX1Trztm8TsnjJNHE1dc7B2d9w
OCOca3Wp67uXPHrf9Ve2Iv60pnnGYUHaubvbzcOrSFrYU2OpEB0N1Zlzx+zFqR4DUtpvx8MO3cgc
ziSEoQZwPqLe+eDawB7O+Tm/VaYLweEQcOPcxyAM4rXAFtwpHH83RpEZykz5bb5F+855jucX4Sra
R4klZDYldvdI5GPOsSFfa4jJ26V+O6t6GGc2EZp8y+YQ2p6SPaLW8WfIERgQ3SQzRQT/iUFVL/hT
GxZ2XRGhBDLzY/YtMW9uXKIsNjwlMsEkLlTJLxl6UCrSRS15Xc9M+iPReXkCbWS1A+ICLAx0kcyV
n2ejzGtZz3nAiC3dg5MEiZDY4slOtzGPbaxld0OpbwrFzqL8P7mqTs8SRxoA5bunqVvrpNJ1uEAp
EduntjibnpnIsZ4lgfWNgq3DO01ZdLxDNK3300LzjvfvVD46lbaVVe7AvcT86YxAQc3uJ/BDl4RK
ooGFnNy0TWS05M6ec1lf/cWCfyhGsXYho68jTt3RdDuSqYs4p5PdLtxkVfj67RhlBhQ2O+Uj/cLp
ODG9I58hN3Pl7uwRdkgZSdJJakPmgdLY0Q0y6gDcmQ/I8uEpI2zXDoGazXm5bPNSmU5Qa3y/uu+o
CqiI3rr4FISYMJVo2oUuEwUABsJQAnywBQd8UiQoIEjrqxS3wW1grSCslVECrhfFx77VmJmbzV/B
IMwU2QACmaSGtUBBatsMjHjcotK1rqwsZHRgLM50VauU/lu9pEqfCG1J48EFFY5TYiqCERce4lFR
MtSVwIpd9mtJKce/NzByu/D/dEgM9axYb3gnX1yfsCgTj0E+q9PDRKOeacFZ399N2sCukjAVPR9b
wpuFBMFvLXAMazXPIp4kKbnJ8PdMUKjz+HztKP6GkWpH+7pRi//kLe3yxI1qNBztws5dVdRa1TYf
4rD5tnwCeyMeM4W1+szTRLP49VhPq1JIKj/aAimVJQ6JE7SyLz8HqLL2YodI3pgTKxtkouoGepPb
Lvx5DzFHTEgyoAg8myFQBMHTeqAjp0pn9AassdzFBuEVGSqQ8o8CaEKXYKKe7DEBs7eYYndMqOd8
EHOPTrsy7b53ou2o0q/+z7+kijY7e+0rQqa+XX/JRlKw0l00CEkiDCS8eD/wCJleKdJ0a6fG5qPO
7ODWaF5+VlxK6R6Cd1nZw5HP8MtRs5JcL0YdrEdCnWqe05UMw1kAzbBxXL2hRcPaze4q0zp61ImP
yyLkO7D8fCJCTrPaS/EgTgcUn8LQSgT0eqshP564PqdPsXNBYW7mopL4faTgAvriDUQkmF6lbRSE
GmBjSgK++MR7zDbGsDKBUXY7VTLtJXSa71//crgx7IJqo8GHmAiVqsuhmHa+gqA8bLtE5sVbOUYK
2W7DWLxNbJYQUIfjJxwPNMeMSGpSCwv5c16CYjuzmG3VK7nqkzVAFoMCBEqXtx9naHOnGBHej3C6
X2f8LbO01Ald7kaEmtWBv+IUM+F8l5vRznxwxxy6JDiuGfJAgqVI1z4c87lQ42orqJrhI+XaBqR7
RVtV5ooRJyvb4L+u+lurSLpzcgtD3M3woIfbwi50DXm9ZSrNAXn5WFyIgOqjqCf3GDdJZJXI79N8
QabRyZ20jIIC8ryaDeq+ESmb14HNulsOFT9g+koOFlm6TIiaoJS+ZwblWyf5i+V8+HXq1V4CNNte
fPdggv3pSK6mnEhbk5hHICG2bJ0t1mo0jIM7ZEIjPi3jQ2cKYLjpEpT92xC7mpd6alnPxUNXBlao
enjke9rGYpdC5QUjZIaaP1UXzf2Yf8uwxm0YoTJvP5KiZkAtx9DK6VpSc/ujv52ARg5zsAL3aCGq
Ww4uNzh7iwUq/cmFcFdATs23JRboXkkjjTXUXsesjQmkG92jXynm4ep247/UbJ8ZIpduiA5R8RI8
R8EbPkDZ8uWYAAi7Ak6mtbvOnd2SHN8VVftU5Nq5p+KMItVRfytpyzYENo0S7AOohKjjMEcO/7DR
WIOn0OsIryVqZAEVB+y10a72QDYOKO4MVWC3Xwhpzba5feJUwQrle8IFz22EKDazPelxYXJeULzw
JCxY6lHxnh3nNd+Ojqn3lTou+8GutnhdrTovRubpofHHKTcimK55hjOVvx0InVzJVcJ09Gkdq9rZ
h172bKBs3yatm8+/Pq/hPJDQV7OPyckblIQnGrHnEQ5hNNZdsRfKs91uOziaqFxCRf5Aidq/RyGp
VPWx6s1zPDx1LcD3SAerFBCmjGY9mAV/r0x3lmTxs7hreTJiLNA5SjD8TqsdT8CP+4RHgTqiAbGI
9IUHL07HvW2hV+gqZv2Ed/7IRt5rQInMsJ/BwPjzImW5MzJVtiu89+oasZIVN719EHoBVZT+3fxf
iaetdxUqFOoMap1s/l8LuDn5N/UsbDHHs6ebFd2h9okait5ambLIg5JhRSYX4IM0EhIO/dT5aL3D
rbpR6eUVwKGX6mDRSCgrGm4gnGTpXeUQjY44fbzEH6dKmwHYGzXstOdKa+9lxxD9CP6PF5yMGOY6
5VKS/6UlrOFPjB5/OGIxMAkEEH8GGChturhitSOGU+f/GyzsJz9PXpUl9l8BdaFfNFMPo5B3hRFa
0G8EhP9p0EdwSwNge1QZXugD3k6m9E18tBpUhIzr+TO39+sItpRf8YqbVAPFUmjTQZFCdLeEWL2S
V1OtKt8k5oloWuUgtaxpaXP8BTxZOY3OKSH3pzYXJpkEDi/upXCa3b/q1udV5YXhUTxJDb+QcMRP
fa1yJ972Fmgd6oYE5x8sBvBWJsb0MOiTCUrAp3U5y3VAUfc9WD8F9ZZWUdOjFb8pIP4NBa1Uiuum
zhJako1HdMgXRKSq96BWYqBzoIA8y5Cg0QoZsZzknMmTNARqNSuYWJH23K+ptql7b0EnYvCEnXh2
rdDCIEFbCM4rcUnkcXOs6zVViWbEvMuXsLKpt0E+hCPvcv5v2zA9twV6dqpgFFTY96bCOIE7xeqt
jhtvW0HF6twx6O4btNSl+K92h6V4reot4K0a9olyWJGJZDi/3+yggItK9h4Pv01PinoWYjImsYCZ
wyamJ13KG8TW0GVNbPHpbnewnYdND29w/pVgTuYtrHN3g8pyZxD3+MthxmWXI14LhHYsxCUo7hlX
C7ujY1Yw9tIOSfML8n4d72jWF+VIGhPw7k+CFatT5Bjx6Hn6HjWgby9wbABMok/GvV5OPxkPWQjG
HmhBqWrdj0uIsgHtlWIqu3qGajAV0vO+fuK0sdiY8jDpD00IaFr/y8qTDzToL9XE4vS+Ln5bR1Om
iH60QBtv3C9Pg3+B0MK10CtgESwpjrm/7jUnAi40S9qd+I/5Ts/aTwkHv6TJOy+2K5M+ZZ6cH1Fl
lniIhCC3U2opdYt5f3OPzpdId26lzHKTamTaCefscRYzEM5wLqu8jQ9rjBw1Shqj4TSxsh6u+4Sf
t+ENAgP8lMn0UwUnkbS632DiRTYMIN1T6MQZXFzEQQswSpCf6buLjhyylTqcDxFeMi7ZHYZrSGJg
kuXjC3CToh7EVmXtG9iodX9n6LbJlQaBtZKZb47tfDNEq/PqxYmPmSq0EIded6ZRFR/i51oMdQsM
9NrDjIpEidaMkkvZdKUi40py8WjwHbMsIsgT0MpPgRaB90+5dQjFcrYk2J7QdTBx0qxu+foyxkpu
8tOTZKDjkBWT3QWgSJPgHYznu6VNS+Ie5cHnYX+SH25g0UwrLUEijg0NhROf1AXkxPBK/8DoCXHx
wcRDgRGdW1mDf1mT73Nh0StmJUCn/aTSoKBaptijg+8U/2DVwW9YK/riXJPHnO/tnFX4K/X/iMg9
T40ifKdG6F9/jcwS9HnxBQJL2xXNmxWf+kT1ejCzPfG07W2hYE5zQlAw83dsAs1ITqBHT5DkaVii
LPOF0ScDA6Di93/nkcAo6th7JqCiELN2OEIwDpZe3+j7kIitvEkAHlAdIGkrP+cre3dwvSs2C+Rq
0vIqR4baDTZyPi3aHJYxdff6QHmTv+0Y2WiatOhRfezMh96IRKgnFHp4R37QPuH9mEiYHLhyuJrq
t7sJPC4sQg5/InxIOCBb5zgE+154fPFc4vEt0lIc4NjqCijneB2tMigh+wctIafcec/sIYa9jMvs
2/D4IxGRR5pIugJtDg3+UimQi1zhioOgNiFE6CEA0nxR7xtiyl1rWGRTg3gVh4qmb9jby1nZr2gE
6ZpobQv9RBCgxjoZFznRacuGLfQTBpBezsD8BGOoUwY4UXAtUBewAJJ4BBj14bsd5/rEW1tXntuT
7thO2xVyFQ0DXgG+4HY4v5rtWZY14bXkVEBYkk7o4Knmb8pp1PW0sMHcH/YECewMgEx2sKW8UiRS
zQEMVaDqhBGToUGK7bUsJyVeWTOXRuiZmy6vRJtnFKZdRpqJIpOLxLAGqHy3Kdnu8hyPEN+x8Ht3
8lcmMtP/5Dhkkap51gFYYb6pbo/EJzvEnfDSdH6w1jc6Tc/+2Na9GsBhwRMsQSnww62USsxlaWHJ
zEH5PyHaKfiDrbS/93YX3knnUh4a4RRegro5IJ65AYGq9Ujpb8nRMdvNxc3dhTUeadYUC5AMDlha
Hji+gsjzMcObL8ZsT7yudWDq5gGn3SZl/hUkYPNR81K0B9sotleaWJBFNVe4YsFrCu/72ApdGhOQ
EXSeRU7TXHaOnkMj3FuCPio5J1bDGTR/nx6358wbK0/rCkhhUGHd/xadQbvvzCtiWD0lDo3kJdm+
5z08/vM9+R8NiHgegYigHKRFcA8fsaQEevdu9jqNiZZG9oV5gAGdGCuHzk4lcW1/h5C+8ANNEKQy
DGvSKWKEjOA9wEbbOJd4yTB58EwSW6jWwJRn6P+4Bxd95VEqnqE89IOGyPACaJDLLSnhGAwsj3XG
iaJl4Ju2eFEHxLVfiLMJXSqsXHRfYhn1e60ofpBaBV1IxgknpGgd3Z+NkDkZKb19xcKp0iBGfLL+
dTevQWFYB7VOdvvrekQmLHKY9QbmpoMm9VXv7yEJ/K3hVA+YlFfqG35od0I/bZSjVYubogh/e5Un
exTaIkajrxYGECPkyltp/z3ktsW7XkqTlguwLyptP/jhwvCfFS7BeyUx7jEFKVlZuYJUPUd67Aua
ffG5Ean8lrWBQ8/c5AFJQp/GKxm2H+tLurx5W2rv/L4MdEX6qbZZ1udHNsbbL8rnb5VKpYFMWE5Z
7cFhOC5i/Ugc7VJU0kT1NhDNBB3cCUYR0Rkz6XDMlC3BWO2agyrQqK36tTSsaZZWN5hASabFSTwR
eQFuboENPTrDrMOgR1Vl7jBceW55ImIvrZpviHGqYWTXF4rToXkLJOfa5JAVaar0Ijy2M8i+s/s6
P92NBbuL3QfAWHAPbL/zseUcu0vYkOBn7Eqv+XPk06nRgAoEu+ZTR63wDCslmcpKL7g+rz9uGMNt
FF5GEo8IlwmYaONlMb8dEv/95OSFxxwo/dPfyz6rSyqHS4LphqtcrUA2EZ2noAvWzjXVTlWC519L
3qNu/fzgdkantijSnOq9+rlsUFfD/OUt6F06QC0TReR8bVZ4u44gHTsRT30u6kPj/0NG2it91g9C
I142RaR4qOhJTTYpOg1BpfVKwLbkIvf0q0t0PML5Ew2cDWrjcA1CVh2kna7fcc1b57GQocN+vuTG
yfBfDN2MpMXSLCYF0fyGIAEEaE9qBsSVXNvL3Zf+YgneeXgdvpjnpDD2BrjW/3BP9pft62W5GKo/
JEBWLCxLtXm4Zk3F3Di91XzjUxMkdQ+JFtsixZZNJ6ApCjSmtBjWMpjVPT/6XWqX7lYpZNt3i9AX
q8zAOcS7+Y4o6wbaNb48RJ3CHExFuFmE+EBK/B30737LW+Kg6ebMaIrCI99XcgOdTHQy2fiOWhj1
EsZgFmtIn0Yglw7r3y5bkMh8kWzkrTOG9MtZCKWeYBofuQL8VCI1Vx7ht8ltqSVDuka8LlGELWIE
lbSFOCzkZatZvq/TEBVaGs4IhzKBFhrhvPK61F3npyX6iPzbXB5gtJwEmwCFli9trCLoAZLbQV7Q
jh6f+Sfn/vcnPFShuTv8ZrUV+efF3qX3oAdRUcK3wuZu9O4v4ufYJyVpm/YXlHlyYf8/agjmiW0l
WvCsj0Xj3ZApDCmZDubnshIcXMjhd4tkYexPG/10LCtxdUEY+5b3aY0DRkc8ZuIE9qXxaA86Bk2J
Vzn3kwxM5AYUchqxyDuRUhAb+PcGKiMutPJAmcDLnPqGJcGIt8moIWJYM3CtAKz2UT7ri1dO/LMt
s0sf0I32V6+Tz50GZiAsbtqAazqkgJlVDbeRM4p1PykfiGL+Gddc/MxMe/0++wkb7jglVxB5rzzJ
3vZnEysHMcjq0AYfQoedPk5fUtOQna2JWIeTajkwBoyq+V493jApRxa95AVqzXwOuiJKbZ2HhCGf
+F9ZXXNQuW/b53ERkNqkfuAD8RMFS/mAwEs+kJV7mo4NObwovbp3D50aPxuU7s+VxtuMhvJxNt2D
9Q76vMqB35DgtlcHU/0tnWUXuJE7ixz8kOe7xe4fkoDacg1lTBA3VWB0NKSo8K9rs3FoC6szoR+B
fV2x/e5vHsQF6ePDXtjAWDBdes9UB/35HddH22CKQyX1MKxsKozIVN6rOZuu659PtzMsB+4X0NLd
0ItYXO65JYScOwIK/mkw7o51fJ/JULZ6PGcvqXijsw3GLNh3FGDbRKX4x6jNLb1eAzDQ3g9TC8JX
g/PruoyWBaq1HauXcOo2qBF94zDSz1Now44dYUsGohxi8HtAMnUC9oLNLu3OyQtFmykd3juJM280
69mDzJo9Nbb3Sf24mhcrTD4V9rTUXqh8V5qJfyDQrn1Vwo8C7G+kNJFhhv7JFgXU67zYqQYU5SDW
fFEu57WvKWD1X2sIP7nluNv0aeJqIf5OgmQ383kl9+ts1JvArUpBxCA7avQzvyiUDj5hAuEfcJzn
mOPpU/NXocVcCOk8fpWptWgFYSNgU2VYHT+oSIZ+tvUJEurj5j6aoBQw2nS/UiDC7tPFaCMeQxtG
1oEWC6M02/TWtnjNjd2zqfP4jai9vEILlNf8k2qV9gwyulqz7W2n9KoAWXEl7zCEzyuaMV8JG7AB
Tbx+WmL/1xOXZ0fIjLQvZer1KOshgKkd6WTE5b19p0AadiZ4YoLm3KLtb83IhR8MxrBkq5/U9OJu
XZo7XHnTXoxdNyXp3rLJrZJ/VLsGqxqNagqfW3OUEds3Wui+d/AhKUkbDCjFQArG7PZ/iLdLt9YM
fADOYusWf2PXUX1SrSw1xMN4AHklYwIbLRoAEodJaRXYWejNQpJYcf6YHe64nVnOhTaQQB7wo5/F
sh+ir4qWzWSxsAHIucvlRLtvdXTT+61p3vG6YXjXlZPglMZFfoIL8bAiFVWFnSMqhNhOhB29tC6b
WrMDPd8zVO2RDM0EiMTH29+XFhTdTOEh62I+2XoycsvBqO1c68/d2rDLSnHLs/rgGaD16a7qRPeB
7pPke6NHM9r7dIojXryp+21CNW7UogjBWqsaGBhxmpQyFFK8RA97Enc1mZl/dmzn8rECfKQlBXCh
a+aL8QQGyHYOEcedWP4YBu4Nl7zxX14fTWvNWMEUEcPKBjBCf6ZrTzQLJPT0UXD4hEQQlls4bfsW
JMhQN7XMdoSnILckmWBt8kvq7S/A757nj5FH1FSoILdjIH4DhDoc39/pYwpXdQEcUZAnpJ/2v8O3
n6U/AqeRUYxVQU+a+83j4+SGgj0OkEwpXs13rwOxXxVc22j18P4+169Pvba+wV0m6J01+KNBUUxS
5UW7VSxcSTlIziaGtvxnrFuD+u0lolZoN3ush3xdxSrc49xvbhutsLRgYWxYJ2vucQkz0heWyHgC
k9mtL0DvmcnCb3Dcg2JRQ0IS3zGLLuQ8F369A1Bj/A4eWkvrfsHgU0rnKQOWBYikof7PVOeTzTGJ
uTOQzdx7FlVIg6soOWpyv1C0W8Om3av5+NFZesk/mibHhBES390alL8r1LtdAm4+VXfgE8eJ8EEC
FI9AcxM/Elz2vryHXpFlCg3nB0fweE08I4VG2SUD+UzcLaKwyAQBbjUhFhxJ9UHl4ijmX5lXozEW
WWRRxnBJiDNj5e0wjSc8UObf1xKQEP2HNAUitfqSloCVvUyaobKSkfqVYtNeVLqwj6ewhonK1gnE
IUd89KvOlUj9hxWXROAdrTWCx9hKhfyiXMXUnmPWALITxqMBKIUpJAqKrtXzxBubszQXatVOiBNL
/ErXFRsPIg+dtxADw3hRNQ2ByuoXGk/t4HNLeRxhkEcDKYFFU+WaOoOxcqR9cTp45GMiwjWkU+GT
hdo23Bzivu0HtAGWZMO8a8v0X62LaYXZB1fqYIOzD9N0xEna7LLj2jXl7/NgeC0LVM1fdwhBAQHg
6dRrIRmmXwbrWbtjv4ynHysABZPrTgKB4PBzZY1TKLgDB1DkvmtnQM4IX+SmV9eqkLo0lM9h77N1
uIGwUni1zH3+sg0o8vf3lrY/+um6nXD0zIu2z8KqK9jtHNFdH37uSTQQXZNKJf3e2EAkmdM1ION0
xk+MlXmDRmsE7kh/c2/f/Zlc4p11IxF5gSZhh4e34BA2FIXS0XQA20pAuH/4423jgX3bJQrhRSly
/346993UU2NZ00o2kVv4H4HpQJWbwUzFLar8MS25UKbNqT1aLwIpemMNl3OIUzmBWtdA8RAWqYuI
1xP4mVGSEki+gbqI7TENOo1TMXrP8RriYDWJiFoDw2u3EtbAnfpTpjA54dbp58MpLLa7KLaKuYrF
xXQUCJaC5w8D/llgt16m/jkR5/VI+68nEnnM5nEQJKcYZE8ML1aMCqjbSSFnP5OWN5ngcwfw80Wv
6ZaP3gjS+LkUwo3Zja7/SNlpUVDzeGnfx8sUy5ZA2ySR/Hfw16yWCRH8tqIdB6l2qbj9NEGX5BLI
dhn49gTXc6WGsCmzbGzWTYtuS0OXhOAxCbYSht8bjZKcMq87gDjWbPIZRTNXCwXgPhMaIxdvOMak
s4f+b1WjhCUCqCU4c9dhArM0WGliXGHOD/VnIlPC0xrgLw0pydJYNkWVeFT+cwNTHtlmpZFc1sBf
HF54uf45QN/UVR0jnMom6mYDIeGJVCqF9xqQb23XxDgV2jyUaj/EDZ4HwMFK8GMJqGgmv6I7868N
BZ1y9UVLsmTgx6ikxIXfgAAwMW5I1TBWnzw+DUyzrpOrqTcOJ78+PNdeCvOs8vUUdVvojlCZRsmo
cxZABp6eneQ7Vgf0t5rw3rSEKinxriKqML9YK68G6ibsHJZ6DssADj05r7NMopzbEG35uQKcYwP1
oCSce+Fj6mtH8VSaNkjwblOl9s1vD+f1LaVZ0umwIgTxdVkEOzaJbGlRIXA/5OidL8ab89WsLS+8
QETRoZ9OdTzkbLZa4uInUBOYAT+NMmt7je/GnwyPJsTbLCsi3mQemZ+akDodLFBZmgiCWVdCRDot
6rLogNSFy6IQwuDOch9YEDqolJdc7yB7gRa+9MSeApmkiak2z12YNMRd/hEmw2UQ8VWeXfsCExqP
X10+90xV5Mx9y+cbcL3QXoj8smXNWYpp7AThmiDGgviaKRN47K5Fiyz/dGPsIP6LyuvGn3Ak46si
VicpraJ2YMULOHh3ed9ouocsnmVSyCaPkwfeJU3zR86/QxVxDoh6WVGuMNzykoP1Z9qEF5rejDZV
U13FQL/gji8ivJCDGAD9lf4I+Yd2Rr233a+/jWk0/HPAcMRaKs7vC6xijhUchrbccP5RS/dwNo6D
E9Xxs2iXrF3r29HckY8abgy131dTzz/q7bNt7v9oJbEq5Ir1M+ymw6yF5Uh3scr4cKoPnEUfVDkZ
G5dvV96EjqeafBfLdaTH27S8UQXUSbdSKc0Z7bwJcEkqoccUa/mlqq/vxsUoKJ/epm6tsPcs0AHy
C6jF0N3U0IOPHU0PGczCKzQD6BG8UGNNIjci8yMYthGlpOiw5KWTUWl8DTaBhWSAHLZvC2j4iWpx
gnRJs31SgD/QUC2+uO15UQ/DGtX2tmLHj7umG0s1CDisnrZE1DJd9biH4McuuwGciHVJknRmegLy
9LKLzQPTIH/6YPJjOH18C91nBoKmomNLhKk3ld4YU8l2w4pUnjIGeWFksD16yC7gBtEqYVy3rpYE
CmNVR8/3+YYY61DxRuXiNzPnUuCWU9c4C9Bc9eOZsEDn0ETA8eJyaEMrzct9qEZ7oVONKV94TfxU
rNjKgepruMHOjv+vZDK7VPgtiXVd0g5oIvTT0AQm6ZpRRehsq2LT/zqcXbTu1oQSgSZrHz4O+pRx
gbMjOWUxk53kvdWbYlb0n1PfgHFqQHPSOtWgnk8O+JU1CCiKH/NupX7pB6BI8vQXFqLVn4xin4hj
hB/0g5F3hABQ+3q/96PMoZ2qx6jxzTzt2zulqV4WB2fihW+0MtGqsLCnidU9vbrbCP+KsjsP8tTM
da2E1jwh8Nj51YwdRcVQRFkeK9odZHdm/ju7mdBLl8CVLCyZeWOCH/B95cHR5TM7/s9kEkInxv2c
LHI+lACf/yPbBzLjWauHmL4hTdlbl3VevEKP4qkDoSShAKHPAJZscFZNsPttmjR5RzHgSj48zSWo
32TaU7CBBYaIw1wjo8EX4AoXqhu6mMzjxg15YB+/U3v90BAzEJaPF+gPQY7ETgaV5tQXEiNpnILo
KQFxX09wYf+6okJZOIifRby66/hHgEwcEs6Ckqw1kFKengydqi/hUIojzdNH7tZvkYhZ4OIiWcPf
xfdUvymEwshfnPniP50Q5cre3Zwgf57lCgXDV893GyVYjREIbpECMAbXbjXzx4O6meT5/UHJP/fB
7usq9/w0TpkgESbGSUafFi7xYKHvxrSstehjr6CsLv/ik4mbRXonY9bGDh8UNTtV2hqVQWesR4uJ
ztvjOE5prYnIXbWTaz9KYAamA3i0OnB25YJWYep9Tlfi70r9lmYlWUm/Ulvr3hZysjKOVGCxBkBI
BijJfqVvZRLAoXM2uPmRqeSxMMkO5jnsZliXYavlEcsbGQLGSLwpSgEPskNTsI+Fmv7l7/sz9WHG
+nj5B2XsR59c4eiK8W7/yZ5ej55SPltZ5+3jC9zQc35AzePVsr69AapgAAerOE8tEVKxUtHbdWLH
dKXFgRHZU2FBa7HTEoZz/sKSRVGUzLZSLSWXosSkk6Qhs7jwUJkd1O5FrUd8/eL98TYy49E0UlXh
AA6DAH3eU8Rp7J31XLYMzV0DZl3pXeSI1Li6w/E4nprXlEfuLsKnGfM1lK3M0uVN4/AE7/9PsM53
3uYsCxIVRCRmHsi+kDoPf8yUlG+uLewRZu9e08GCRwVlBzQ9RDEr87AicGHHUacBVOD+81Cb+H1d
0d4U3SZ1pf4jQ9leAfImsqJWObrPuBkW0+a7WUlEABmEJ5ICdS+qUnkzmXhIZ/PiRKqnwIGHnBFi
a2DlZBHcmS+xw4nGdKKyjlO6CTPX17kq/EKbvGBZogXm/5SutuMd910xRRLoVtrcvHJvavHKV24B
ilvRwa82R4ud49WqvUWu74WgUeeWR5nCnCyP/YFSJc/79Bmc99hYQkGyQ/vXn7kMb6+qtohHeTSN
2CYt5it3WguB7J1fRQwQjbwY4osR8hoi457hVu74c3llj6A1CwieZWCpe8iLrOX3wn/WEQ6Ddy7T
PbztVdAIwDtvnPvZD3c5hWkaZWWddU91HZF8FZh/v3+lz7iOiq1t9MOl7KqQ1v5YUgqq2gLGNsyD
JIUSiz/QVcz4mpf/ZzRqSsLiAEgcuoJOfaqeRHblQmOCocSE5o5c44zPEd9uLLHQ5T/694qqY3SE
nJuvId9BQ4c4lM3APqnEGtCn9fxr6b0XCnX/kyo95/KHZgRIfrUo1F+mwz1DVPmbcxINpwKOkjxk
5ADxeenOe5s2ljDnkRUpW+crqAn7aRBTLx/KUFz5zGopNZ0T3zIvCVpdJKi9ccbOxblthO2hKfv5
rLW8xMcvtxxPJLSvY0XSZIRP3NeNCN9HDJI8pjAaWKdlV4V5E5PoVAnhdJyBaCBkHuvjxWsB9WoA
zS0u/3r8Aq8YaBpFSd2AQDwH9+VUJHDZIlQg+vPoGvWhyEjU0luIFtWkGmkwf/EGecsOMCv4A6jJ
egUqZ0w8zYAh1ziKqbt3NNSyuO9QVFTpcUKTUEtNOK0508ONUUWhUs92tNaF/Z8yx/0hx1b3CBLr
xpyFp9vdOhBsqJEFBriZDr5WP0gPUu1oKLkr4cu9Vb2LH9jnopVF8hC0c+GhxNKFTXCq/2T2Sa2N
5Hy0UVGjIv3hgPKTKhxGXzGfO54jpbN/e0JGClfvYr8cHhA1/9TyBWBhxJZbcBT4jXP7NnNuDe62
LudmTtylRbRN223tX1KBjn/WiuhnyJEzImXM/6XyVspwq0BBS8xGwArUhsG1zuyGXHssRQvbq8LY
v5mg+SsuG+IoAnVV0BjeU05C8pUF5rzKrdpNReXNVtlBq5HZJ6jQrCvYRkgq+4+0UZC5JLCZH214
d18dkJXnkq/AWv1wZV2jX09B1axJXpOeQ/v6qSosPEye8jvMvlFK2XNP/XxmuvzX3kZTi467wVBv
RBn8/3sS61X9vjc4D8qLbDkdAA7zXkn0NkgBHwWZUgORaEmFGJPtgF1o0rsxnxGegkyZpmeGgUtm
ZSbktgH8j3y5BJHTqBlLnHBU+lEYdZWyyYtSWa8pKHFQ8db34McPNLUV5trQ21ns+/fbaGCdoGkg
EgUGFCD9kE3CBdgARC9JKJsioWaouYlXojCPOnBFRntC1nZX33VNs+kToSrcMdMsdzvcA6GF4rOj
g3w8kgGDoX4/3Te3/BD5v9wJZ6BUoAJFK6NoqO5f7mkZjz2Kk8hcNxfgLPHOFh7DXRv7Ab0ps0fP
1/BunqtTGiougXPrdWJqdo8xfANnMx3e/XP3Z+448qRMFLIXCFnzXZ4ATeGDPZnBG5aBVW2r28+J
SYvvDmtP+1wRakuaxpIC5aVRddpQgW4WBxEzzta3T0T3w+T0TIq32Gh9Wme0rYNtfkUy6+P0z1sc
Hfz47aBNaN6srHprtACHwiMnbFxDBqCZL5w4/ZiFeO4qpeKP4j4JDZ241YBCWIBW+cIfSTAtGBXp
mizz1m9LoTWBR3rDbUsfteY2eRi1VEZWUhtk/cCVHAalAFPZAP2Fjs9SK/gffn8jOnrSTRP1qfhM
oF0PzeLX7VBGgbeI3BUvbMCQPRkafjZ+0vd6C7PDxrqcCo5rCqAQlf/LLY2NTpWuub40sQkv0HKK
94fP0T/4DZI4MA+5d4WhHvSame79H3nGFliZwR4jf8zAdwVy0zNIQ4/ezlm9Hr/TXtnANzpD0byZ
CQ/Qgy4fnb3yJuvnMW5dHb7/8x2DGvlvYTvlBVLRo8JL80Ptas4DXateJZoZcj8QFNbl3PTyjZXE
U1BVpIod4+ikgn4ZBnB+kzsCvAcLOZFioWG2BiiU55Rm2OptYVFeT78zyzkcdHFd8vp9b1IpoujV
p8amlZq0vhAoAxTzif4wKbRvKDR0vkoyu05CJ0CVzl7vaJsURUmf0Ekb5CyCi29hywiqMEBa85rW
/fktEib/dWFIrmQ/pCOOg59NZZ9B02yH1ILu1MNSkWNDDWQLobMgk5WucYb/7hUpS/5u3NuofBpP
y0TNHa9H3XA7nHJp8jjfDJTCGC7TfMCwl/9KtU8AX7YW1vUl1bSFIO/OiXcazd4XYPxPtThiZ9RD
ltJqSN5DVj8JsajdfgJUaLzlBQCyULh+idlAP8CxulcVs9ESxMqdplzB3dfp3o5h5UT3dAcYsbtd
eaLe+wyIWolenKLKNNdyZS1CYzcSZ5T4awmJuxwyQALsznoE+EFuDk3NTVv3ZD1ExZwVqwSs+HcV
gjq7CYWwWBjLEN3orv/swbIxcFyqrT79cCnyK5iUOxQVzWsuBMXDzwcEZ6WzpPZ2pcjOfMz35qCd
nusPzLiaKgp7qURpD7aU9C2vaXon5q5LhWQkjL8bmmSImvOXZFgOlR15OSFQVAk8jolVbIUeh/Zd
6Xmqq7m4cA9hvZKfyVivWkAYwXOe1IONmITjV6GQoAp9WGV5/iY/yHrIenN9og8twOsQLPfbcJmV
LecWBAgIpGypwUo1PiluAcbq06CYO1fGVhZaEeKNfugWwx+sfLtQKl/IGw1DjXdrT0rpqBqEHh64
c/Rt1YGfk4f9jxwK10M0qJNrZbPad/59gi2mX5wOI6cMjEzPhSBmjy1wwN87AWQnhIY070XEfp7V
9iC5pIqAZGSMFsNaOtRV4Fl48MgI0P27qELrul3HwCoUm+XrFglcxxqlhUSe5oCDJJvNrEthzING
slEdfNizUV102OguYUhtAA1hYNdRUIbrD74hCZqU5yCYJf/UGf0Sh+zL4TSsmdWCqnIbh5rHNzTT
x6T15fH1QGcmuaiT6jPmM3AjYXArK5sqJ2mZ0zGX8WMkjg41NWUFcdRd0d3IjHRSStGlzyWeL5H7
zlCNCrPFcmDSvUB4R5BRt7/7VJj92/QHPn9kxw5BpxzDPCS6Hh3tTpYGM6Ff0V3iUoq/yIWzUrdU
POwSTaf+ihW3QS3IAMeGqvlQAQEa72unMlvMdhyhGcgqATbRzs2e/+swezM2fw5FAqMgug2GvPFl
6Vb+A1Hfh/hEdOhLvdC5Ng9SZBZ2sL95tvuWpHV81Tajd9JFCCnlemFf6xzcU8n0Y1Jn5qq650FK
2nqK/MCG1DM//m1n3s7DwGyxuXjlKymQ5l1G+F1Rei+s4GDeUyC1ArUAN2Q4y5ycq1HOaZdJVQuq
5kKI9y63KHkCOh9WRgCwPL4MiVFZ7umPANGm6XPz5OG6/ZcI17Db3F+FVcZRxO1BHBKoWaUfwSYa
0WMGHB1vnsoIhijWqGPkUlcXvcCfhzozl+uN6We7cKWRSVPrTi28rWCLu+W9/BubfdDKpB2NTkWs
Hjohzraz1OzYA22NgAZngLJ/x3Udwv4pHcDcHBUjT7F6Y2k2TOgD57Xt3IEQZRBM/LYuCPnIY13k
OrYhM5v3A7g7IZjxvVi8BD8hF4z0i8WrOknTYJmyRp+UxhWwthCye45DbCJA2X2k6oUOCUSqt8vh
9tUf/xNzrJ2s7R1EWf+m6H6CaHM2BsyDbMU9kNu4S8qqikEjQjMqjKkZyosdyemO4VVh8XcYVlhv
zIf0WtBdWIKtGFDzQF3IRLMV6dNpbU+/f+RF/pjC4hD4V7RhjC+JIisEp88Y40HpGZpwX59hgtXf
ag4S2kou/oqHq8KblzARhEbm54qbyPChPk5b6g0i+aA1Ao+arSYFygaKWRH5a87rDubIy2bzIL7K
1M8RBgBIDqZDQyNJMrc2+jdrVnUY/H0FMSJ21ijwTaMeXk7jSzNoXaYAlpbKzv1Lz5bBAGwLPtsM
bYRn1kQT4JDjDcMVoLN8Kk0YnQwUegIMDCAOfC1SRL0nz4KBZvyU/+lsw9U1AvE8xf/KDTON75mJ
8p2UxvUoayeBpmDPvrxaHGVlVaJ050L1THBzJUca9aQzJDdkQHXmH15OSab7OumRFGA6rJ4iIGqV
hKWJDuYUKofDqC42V9PRpMUXbFbi/pCYYmcJxwzfyZEZ2zyp1x3EQUO4E+6w4lKwjJw7NolYUEG/
iKRBiB8vL+Pm81A+ElRE4nkBtKpfDXG2s6MfXaWJ3nCYcWlTQ+mbcJhiiCOku2VcgIhVQwicoD35
+j10cTMtKmObtYqOjRcNgPhrcRmNUL6c6ZXdl9+pw29D4QU2B0ny0sgnJhqsJfrRFM57NC50tMo+
2JOopaEJtAeYnWe/kqPGA9cuT/spoHCwxzpYtVSiVVrsgCpx8vEPOOOALjNVotOAfqFdu0Mhol1P
tiAeC0O106eT1T+8Y2ngBDbFhafb8V/J4wh9mzumZWj+97D9+cL13EmmIUwX4UaeFxP2d3T6QxLk
WMZbY8zHnHslizQF51zc8ZA61D+91zLEplC6PwcT4tb4+o5UkR102aDb536XV97RbOtCk7LUFDeI
Iy1jnkmkpAuH1JaU9QZEzSgsu/cFkJ5v6TEYk604OsFxsHR7EC+pNQDnWeAv54+OXyIENTN9gGLI
I+nc340fQqxAf8C06UFfRcQLNlCNhRHmsMCIjuJCyEZsV+fkCS9acO8EpExcYTohSln+te2Y3gRb
YfidW++OjoZFWsk/gFCQ6ICrF0Gva7PQSW1N5AnP6UGmR2WVb0JRF76m+JLiah7E2rq7rPdq2Ggi
HDrOC7GhXuG8+LkponErJttsaCCZ5FTPJwqixUwoPpKr5X8TQ2RQ8lkKwn7J0P7G0TiMQrxymBPW
p9vZFVLhjallqfMdLOrwqucb2+HGMWfu7FIX2Kk5b7MStcOfDdmi4TSE5GIZ+ksQMOchg5aX/+Ea
e7RzejrJasw6y9ctwqK1cmYVEdS23u692/nD0MeYfQ5iTFEOeGArhBkhmAeHy4PsRoycSY/feEqz
GKTGk5lYZFOQ3YXdHZGkyBSiVMngBO9AB+Wa+wLlwq4OwljhI4/AyfejVmxoJjWlo78sFHWpSmjc
WcYG2xIFsWDcb94izFEsVBJ2DGfg9SQQ61xDvSqag/FFNDjMw3s6wk7PFEeQDj4aj6mEdPPfLyYi
V12v6Z6VaV2NNZ03AFirOhvmN9+bRz3okkZyn9qAgLUpQd6ZHMqJQo1LPjqPazK97FFKRWPIRq/a
qTeACGgiT/Rq8W2+85m/4K5eEzXcAVQ7SI6gPQbj/2CaMmahyorfJuOB7cwVT2/sscIit/2zC+ei
oK2JfG3RSU6nSk8CQRKqzdovQlSQyy0S4MQ3I4ck8zq1uyOcNr46YtdXPtuKVUveS8esn7DT1H/A
IxEW+bdusL6JuvjGPDHQjYQy7hqZvaCdR957bLm2jefauIy2vHOy0wOqbuIOEEKCIOZXSFyl1ZM+
ghRfaUTk+IpkcyGZNrWQWYEuRqob4UV7uh5sZd0qc0z+yr9CpBsW5P3ntXXcKXj0ParyvGtuG+EM
c/5oY8BLnR0W6nzHx6HzGIxSXD30i3I3m30TcRwf3RUbd6iWu9pZtATJL3hdVdPbfl62hsO2LUkp
K/H5cL066YOXbC0cmx3u7NSkUOXmw5CHVF6JbSf9w86863lbr1RtC+556ZlZ35oJJdZQtz4+GvLj
6qaQyoj2SSJr10Wywn0caK6SNuniNK5cB+J4IlR/pRe8a0fe1xXsQTZ4PFkxiPTqeeuZAEErDiuz
CffUihjBpWK0rUHO491aQoSlDHN7lVHa4ztf8Rv4FMp5yBPj6X8jXNdXqFhgVa8XUhpFRDyZ5Wo8
oifJ9E1Xq94LPRAcM/ZrpQCv+iKRLGUWn4sECIf23+TSRq9bT6oaqqyKGTcLqB6vx49OIRHkPKsK
AUaLIsDHc8x8PaVzkSvqinh+ZeB99nvv7Y67faQxB+3P3nytehw1rnwKQU1Czz2gOeWJkb7NnTKX
WYK0hIruKCZNy5zz9UTjAWSPHIv4i6SHzwBtw6WiNcXNRhkp6khsVplvj+nvouPZu6bYIon3kYdg
BD9FDFWZO+Gx1+ivFFEV/Vhugen1YgvZnXNMAyi0ftKMb/TbH50YDPcZ7SaRtaMesevycPggZfUc
eavG7mPIoLYf7WP4LAm95sjGw99zZSVi+6qgzeKVQGDSYjQ73OitY+iKm1/QCoZuKTvlqrWhvD39
qtK+FSwJQZZRoXVcK7WHxv8wsSb8lFd6kE7J6ajGar7OM2ioxlAZXg4EXNU8YrEg0lYf5DZIyhjO
hxjkSVHOaHoSELwV4u3s6BJgLWyrv1kWoHkipaH82FgHWPuGrXCB48nDGnhFCIhFPlHAU+J6+F4o
AYlj6w+GjmQE3+O/j5S2iBitumcXHDYmVPzL08o5VYakOYVHxr+CefnCydbYy6uUbaIHNkieNHSa
+XH59eLWD+PzTnKpWiMkCZHsOhXQ/74IJaPr8aEFJ4pn/yYyV3mp7NS/wJ0T39dM0DR9CfQoauUK
gunQ/5wSa2NHgNgcicDrrNXp74ucEb/24LtPPnbFm3jw2t8mrbn/Bq/38bC+ljJZ+/wf3n1Hyxoh
i7MZ12GCc1baSDkv+Edvol3SIe6fY1MYVDF/CaceggPUEWD3BtQ0CG3ImLonxM9g1+Y6dmdXSgnU
nt/Gpl7DVGxBI00qTNR2xmJ6foAwmsSCV1NXw9y8gCB/2qHVBpgsMRvZKmKz1TnptsEmXKf/ne/h
zlAitZVWD7LRVextgJ50g+8p0JR9V64rD0obl6zHXRCw7iA5JVxSVm2eBpYy4Z0BtjLsk//pG0Yr
nMKUnVLIXT9NPNlcJignZsOQyo5ItdoVt59mA8AxpHQYKQPXBO3jwsgkw+XstNcZ+pzNBaKjH4An
U6mgJHKYxiX0tBCR3R5nwNF474GN+2jw3Hu+tUtpiS6a3xs5IRdr05KS2dswbgDjp2GE67DcDOlf
wVGTf9oki7bLG2KZhZU3b8odj9JrcBo5lW2y4j91ceYqJ0ETtFUv8oNWWm/Q0RgvKgK21bOSa9ut
sw8DbPbE/jcNsOcj7FuZGsFSvvcT1o0QR1T+8lymQbPmY08T3Ng/tnEnVr+bvTh+mQ0Ar7ggRFT2
On9Iki1pw/QVOxyxnhJXzAvSPrRVp59D4RxvX0wFSjfYLWewUeMVGRNAw32DlUMd7ty/Txdo0JeD
NYAPVuhbfTt+m6/1EpKpvQZpGXOkIahxQ7d7L31CocjavoQWZ4Jl4gSVMycLOLkcNCXIF1vlhagF
nG+w2GhraFJfTH+1D57aMJaqvjSuu0ePT5KiIVk5xPeT+eWZHkwyg+EOPtK6xs3r2ALaWI4SoVU/
c7/0Fn12OduOL5tDc4dUtiDHPvkQU8RLYUuHTojKfjPQrErSI21bBErpevaXnKJOAlPfTDveNTbL
Ks8OdhOmgmXEWrSuSTeSIbo2HrrTBRGHbpbHEepYrO7Gp6bBlBypW5VmhwwjDeUGSLpcshZI+gpE
4uhPuvx9Y3qNhqEpA9hfAkQck9XG1v997XZLI7io3PVs//FIelKAI4NCff896NehLwNpDIG39awG
9cQAyuVAh4mVamltCEkyk7cZyjtzgqXqzjn1eh305TgKVwjayPmMfo1SHrYhpGVHiHR9CrAH+wvR
WaDfkx2iFuxTuGM3uSIYVWT3w4Gr5kDshQ+0o1DJCQekhnxiCCyfjDWzNUa9GRi7W25ZWzBfQkhM
wR1u/VolYznGF44Lu9H1p1xIE51sQn2tWltLLAZWFfED9Nucj9DTUhopFHvEn2v4Y+FQ4UbKdlj5
B0+c9wSv58yDkKoG3PyIVjGPncMcoy8jfB9ul8Hcn+i+YZ3cj3OalMVhi1bA9sei6p2+koyt6i6W
gNsaE837V+TANruy1gxd45uoadQrYbA+30jVKtzDN0CtWlQN/4iqeSSEoW5qDF12UuGCYy08Fkxe
KLuvHVz1sHSQmSTg0r8pmpfziROeMGpD+pAs3OKktwvHy12EW5Ca7GGLJ9XatYk8MsNofJ+86vjl
i2NgeSVr1Bai4aZMoHoHva6vCrpN6wgaZ3jdfLlSbF4xuRn6soGBQOP1YDvAvcNoGXcSDLqrvaGu
w/vLGiXlV0GhFzyKlTzcJtZVpbU+GFWmYWu4fgjG4+DQWn8NVFG1QhzI138w6tfcggybqntFtmwP
uWbFCs4lWfKVTyZhkONOwQWl/wJ6Unmx95K2w5drR9nczUUYZRzV8O/Hvzhokj5CgiPPN6mrqpJM
ug6xL8xPpAzYYUJTzx6g9rLvA9d6yCXufZOu4wnVaj+OnBe+bKVv+z2WVSPcR9eMNPpy4MJZLbnw
4J1kqGIug1a8cbRpdcgqlf5TorOqXR3z2onnQgMG62f5nkJC2nrcAHAyTfmEGfvKjdpJZdTmi+W0
P46zEw3LngAZyMwdJCQIIqP4syI8PmF2oHOojrV2iSr8rPmxBP+utWI3Xh0LQkfSLzekhpWhItj2
YLWiLPlI/fLZQpz4ibUItnf/8wtE5dY8FqbfyXxVFYCCl+lOP6WxD05fQlSxj8Nyq9pW+vmH26CS
En8RjGvZ18L25PHHdZ0EoPqIl1DlNmv7wCpCM04Al4X2NWT4JSm4+d9NDPdrcex4f0kTlBJeMSYI
9XdXmsAucLZLekFrJxa4MF5mJ80ofakCditKr37T0VYLxxN368pyaYb54DsEVeu0RGaO43KVdFRa
FU/aui9goEHU02lMg7Rz6DzXFIZ+jBkK5qLqOuZpy53Qz5YvVQBC/IN/OONbOhzI+YbIKofIj+uE
i7PMit5jKiiBVab1SARWH7ZWaqhj0s+a8YlVZJCCPzbvpy8AU9pCbladj4JYRdgS3DIzxJaDqnSY
lJHcKZZRM4yznjBsrAZ6p72m/rDA8iX3xPJyPCSyPZ+PMOzTEVQ+hRfitdczbh5RWvt+a7D8VsmE
faDvcZjemjK9R8S8h1MKWch9AG/WhPKmfa444jU26r3Fj1Ynz3CDrrZutH+Ar8g8/yr7lX4RqKAo
WqMAwVzJOcWtek9zFeDrirC/D9gTaatXiv+zT/owxAR6dcU+Od1KrIjUrcbxlBtQdgThkMuDGkLx
xlg+mv9j++BssSgXiZTz2IkQveeBH/7VQRKZ2vuh4IYnEhTY38A3apO5eAbLtquy++qRGqeDbncm
5XUym98KVqvyvT44TwXz3MdoOnFwetV/PGfbzMK1w32L+GpEkrUy3QdoCJebP3RsAArvHBWbGNCR
V8Z392U8E1G2HlU0xXgHKEToJcPj4uY+m7xGjpM1J0leRAqBHc7VITIL6nuuSw7Ll+nmwFORlHgn
ikn9OmoWSjlcZUTQQ5meF+Ur2H6Vi8WcPggacoUWOIEZGfpCxNN6kV0h7Z0cho8blWPPbsaFQw3x
3Sz+xVIsxkFgHLhZ+fSVBaI2SHjih0rOURxbUh6XXIwoFSY2NqhVEtlqvU4NYY7f4E8ATY5oBZJq
rUqayujDdNR9AyfjAXTht5XfxsVg7k2L+nJ1ApQ3BIr9dIuWVKYKl8CtXbgPX/1GujGmTH8yLNQZ
sKe5FyPSnOhbuxUjDobpJDAxuMg8FlxwBOhezDTTSlOAOIHjeb1EkS2ifjhAwBe8lrcFv1Op9W9K
ETgO0lmAAzLQXlLmaSTjnYvehaeZaSwrQ3bPWbXJ6hU5mRPoCxzEGV+jDpBkao5L6qrpc0xJ/yKt
KgHtm2PQyvQWnHt/MXpfaOREas63ziVr+iNUjK6WvUV/Ra7rYeDYIxVhrXlIqwJH3v1iLRuXKYdz
8vNps5TIqrpLlibiP3wQv6OSfp5Hld4oIjeKEUlm6J/I/7FWzJcqSd3kYD8qu/fzP7FkZ+NbJVm0
nYvdMuJxIVe3qWXF7ZlN/XBESchUYBxUhlloZjqXb+JywwBZkqX5EI2Hh+P8771gpijHjVH+FvGP
raSihuO2psf+IewUWzrhwPN5YOcei1ogspT/Z05Tx/Fgpdp2ZQbmBXtQXeQe1Lo7phfb4dYCVEjI
3YvGj6FU5d19miwbUc55rqs/SlEd0pMKbdUXrUBwFNDq8itnlDhAyOQp6JpO1poyd5QgRMzY/RR/
sauY7h6YqD/7/C+ysn7t3PhephEuwclZYPFgcdXRuZHs1B4wH+3y4RDz/MuAiCwSxfIYXBjbFDJK
oWxzOA/Wq9U14+8svQiWqIlRW5NStfR6zM7vcSxfOdfPwlXhIbTfOyS+YGL7kDCGXLqG0tdssN93
dOiadNr+n9DAlT2b6+9e54wqJF2jKvjZbZwz6SuvgzXbHMX4uOKrcAs9VO3Qwf7xfonHcS6O8FKi
rmzCGGsG1McDvR3iWgAboh07S+IaIABvhViow5VOsFQEmpQrRgTePXe22WhGFQSs43Hd+qLexXgP
753DSZRcAE0VmYPuF5FZbXIJ0bZXVIqfxR2ckW0O3FkdsixCBtYJbmCo9VbN2em9TFl0s7OovfFk
8uAio2LSZCmrdjnPs+JvnLdP9Mnj1AdzLnha1poQWWnDx7woAaDi1FRd3UZ6Q6k9012BmFa6KZ8j
3PZCXPu2sOzZgh//D5W3TbCbFC0UrpXLF3iLTlVwgllXlpNTRHyOr60DjzyinkjGfA57fUwYNw88
Wv3dG/Q46sgHtTvMVlE8mAzOiTa2BH7RP/+zi+iP04nZ58turKUxdPo1yLr4taa16QfR8QNHO7HH
OHbS9PkoXI/Ln4zg/5S9lax4sWC2B+TRZ1KpbtMf0zGuI8OlJY8QEQn5usoX7xJxbAWrnJzA9Wkf
wzWZvFscq2XNwcjWkzmebr2eXBxZTAEOVFBvLsXX/WI48QpJpMv3DUiU40vRcJ/kWuhvzzHqm1Z0
JX/x3x2avhyTiMJWo9lspEJM1MlhuHo5Hj73tNyDBF2tF0iscpAx9bDkHb2aOf7alMkZr8pb5s+H
PbAcv4jFex6rZnsX3oUiS9IQI4c6bGor67GSbOtP0xvA2/L8o3V5zFuump5ATMaD1M8ei//T9aZ1
o++sxKRG9k1KsrlWWWuXEp+rvrDJrt+/GFPexF+cyfbxjs1ZLeywMw/nhsSktj2qOywtOIE/p6EN
k9dAu6b7g667W6g6YuEwq5L1d9spyvDX1AhfbJQ+ynNJUzGdwIQnZy+w/K3Pn0GfSDQCxctOPqnB
PmolvghamzErqdcU8b5ehAYIgb7tIGEk/+omwdzyrnuA6ThEnw7vMLX6gQSfQdYDoXqmSG1gkKzX
ipAFxYRWaLr6uuivQ+pt30lOyPfXmQEYPGuPiOlLveK8rs/xyQndONCx43zFWmKcLf5pyPYuObP4
7Q2/RjSjnXh3ThpGCgROM6rlULAwXw9+tv2YdqB7rpvWoJPru3fDknYe4tZME04qC1DRmzXrASry
d0KOxSxxk2bhve6vsbKe+IHQziB30xogSNkKneLF/OIUOPUqszvQWpRArEh/O1EdgYCROvQUOffj
J9lqxL7qfQAFYvXBqDKosEdnJCQB0hJqJJhr4LdOvQTpueaFf/aMp7xyf7z4cvhLpS9peo2cGcIS
6ZlVm/9bjZ7VUMPt8UJUo69mngU9YrcfLFivoj9+Yn6UbTJ/fRZeFm7IUWI8cgT6Qct9Riz+rlK+
iVXFDoA29ZtgL0iSggtFTyPHVgAzbC1iNzTvXOlPG3WlmZdUlwyrsuJsfiLPxCnUfWLswbgiPuGo
CJTezKWE0EPBdLy3h3aw2kZ1h5XZjf2T01CNhSCpK9jUTjafz3wYiN/KBMOtj/muAC5M57pvToXS
2/Wq80GqX+07gGsFDLwXxzj6iJrPsR/gkAFirmJ8xUJO8M1oANLRG3bnaucfiyrN608AoiWcO8g6
yffrX6kHs/KyOjUBLE7dIJksqvcqQnTNPDgzkEZX5XtocItq6saWGxOT7i1mhxnJYfof22js9Uwc
uy1Q6q/ooALislMYe0s+pTyga7ePl2mywgIy/C82y6ka1pjAKkRf1dMdBP6T4giKh7bNzBwvcwaC
K/S/DdyAsA+Ty2ygwDy7CMBFuPU8laUEiQMrl8uH+umXZxnuBgfGkC9PYTyCAa40IaHi9wnysV8w
dL/U2u4bK56AaAQa8b0CGHuch7OoY7svRz9MRuXw2xiZRR52gQmh/VeC0wNrUL/l+YHwOCl0ed/5
BC0ByKm4amXXPKf72r8otUK60Q6Z00oSAILKjay9ZxYzC+jcoHbt57aUL0aX2G0M0OST5zwPjtsl
DRGtHFfftLfxlAXvIvWv/KA4Xp4oahctMYfGv6IBfhC40vGxQjUrYQHKQoNOSXwSc84AAbT9+GSM
bGwDnrjM6O5g+zy+UrXJB1GUa5GkK4mTeXUmQZQ2RKTPkQKnmm59PTYuSAEBfShopeUazyPDVdhr
l1ztAko1Uu446BpKTK12Y33VZIybk7aMg7jfQhb+c117vBEPRs6IThrSmJUPg6+aiuOecWuFJCBM
mOZ7lM3E0mk8zDXffFJDSuL+fJRcL94osMAhcFpF/7dwrzU2NRt50RQlxZhD6q5mVhxJcVWqNij6
0VBoMS4PF+nSs5uMVZB9GqHzpKvAEQ/0kiYdYE/Khvq4yfvnbfEIhEfx8ZIT7zvCXwYra0+Ka7UQ
tf9uQI7nOymjmPttATt8jaMkVYqZfoFdtfnpqfm+HmjQB8ATrpTn7yuhjZ0xXczpK+4Ke3bIg3gd
ph2gcM+w6ZPntzUUtFkQ9CcWFS8CBjSwDwiyrFnxS46nVCb7EvKB2O/aHqr70nO2QUsUzibBOlpe
cPpHr72gN7OijKRaIhqinX9fKNQDrvBRXheA0V1076ahip54LF5En613SozgZEM1XFdkz9oHDuBc
sqE+F2R7GsSa4l8dEGOVPF+rp4eHvnmniUYhTeM/NezKQ2FC9ZP2fEwJ9bAOz1W7bPWy/zX2gyAU
DBBrmoT+rgrFlffS3iBT1/ApAH1UtV5A4h1GO3doxq4UQpU04jE0F5dsKs8+VlXWP437MIYk2Dq1
YbUxUYvrIoMIh9UkB6wGckoHlJGOOARKoKouW4tEkjwLKYf6vRAxuhd2vxjeB8MzoFP0INAnAZY+
bKh+MlRgquVbTCLbsO4Gcd1/6PBTTQCSaypztMT3c/kn2Lnl+7giLvqoZlgadN8T9e4tdEKjc8Dd
tT+rTBax1FT584xGB18UTfzNDxgaquCs9IhXxKtRDO8MmmwagOIdcYVAkKm8Y8BswfkKMxvpPlvk
yXeih4FNme5p6A26yy8TIoIDFhMm4K8o9UY8b2ecR4DovDQ7xCEWltewlgpwAivDmeJbo97e7HF4
tXppvKQWZcPxsjg2gVxVEe9RL7rkCU7XcsgEQWFyB1QXBex7LriMZIo/E0KfWKKzvT4ycL6ozxMj
dhcj2l6lYuLIqvkAZV4Rzut+cFNXvNd+5rn3Yup+RRQcxlaKnhJlnJQUz8K7O38Jj/PC9oBrOMMH
P1mgL/zUeINYykW1cBFMHED+8fatLMALkyHajPOS9waauszzB7CGiEfHk2OM4INOEKeI/cGqrauN
XeXBKC4/0G5nyI5S638rCMzeSYoSCBGt50MsOdizafch4/E3RFa0Nz8oeZlqHUulj/mHfzkm4E+2
z/F6QCLQ/3dqir2F8xC82MF2IFc8WYfqoOYy9kXEYGYimRmF6P+bUka0YdkA1/cLulvvr2gc+bjY
GWfIKa3PDQV/00oloXs4w9+/CqLYLuWPvMdn6bh21dlq1pxGByur8q7Iq3i2BYpTX+Zx7nQ4cCgD
YMGWCaexA3CxiRUb0BGpJPdcQGQEiivW2PiVpI7/ICxGYSCekGQvoPRrCgg69emcF5GU5NSbr4IX
MBFCYZ9K9Lgl1a9fIfGzFcCLShikznabKJ+XqD+eOeONbyZVYoTrQS7AuVXrR4o77dvY10kGyoWU
06MytYcro9pKdAoi8iztPNiGdXRRmXSiYFLztsSOspmONum630ChXB9xdgeGrN0iOtetE+1hfe1u
Z/xFAdcggMGwzwP7tkcPgrrLAVRo4gjAJkAqY+3aFRn9ZgueU7e6joFzieP+vDJxOaowtPn8zOt0
aIJihjIp9weu5C8NZ0BACYAnSURtGVjlxbzss4B8iVheLjXa0X/Y1y1On4z0kuM86FGvexg3OvyP
G/BDJyrpro1MMxbu1ib6ng6/nINur4D8o5Ipiiv/a+85YtQBKU7yvmx1+QOvMZ+47N3JtNax+Oiq
bUm3yJyxbgYc/ZSfuoUkvryLWpPPmV97MqFZ6RlWgwETDxBM1Tx5z4FFX28yOSLdR2SrICg6U3PK
3eEOGlB+2vLGMnj6Jnc90oDisCJ4V55R+MZW4VtqYHpzJ39cIGErLTrW2JenFkANlME/WGJgVxZK
uEcYBZPJCsrH5ydgSeKrayt+zn/oWfnZQIhNNbd+I/GfbryHYu32wVj04MpSl+lKKFIXdKxu1kTF
xGFollVTF1sIm6Cz2818z5gyHVukUjKkia0O1Lw44R4SauhFypsUkQKWk8p1kP9TjfpEMIW5c0aO
YiIO5AE6pE8YG8LgW/NeNxJ20gTed5O4WApHLG8EeysxRZ9nQHCgoBcVgyI7lmF3Z8PNkj3UhE+l
uzoGJVUadWLhlg3SW1bHLZAKELo9upnRl2dDfo7ZaL70pmzZg1cFywo3xcd2G8td38KyVM17/JYr
ktZ2VURyVzIYys8cZN/gd++r04MSEsylN+7z5IqW3jvV+lXShbOOesuB3lhlvqLhdMKjdqj2gTZL
/kVKWjzjno+mjLKrIxyM87Mdxdtf9OuUmlpGflg+fYFtHDqD1fhjVUcIEkxzvfZiNF8wXzh5jSff
uxMDBoEG5pLAoGYGzd9SOi/AGTWALky/w/EuEozVtVhkyC9g9eP4Ikw3LAGEmHGAZnBYEWtihEoN
cvblEQS7i4YIAdIcxe2LLoJzrSvH39oj3ADz4jtRT6adbTEywVEIBQjqST/HkO9+tPypsLJdvm1M
x+qX/tKMUnSHTUe9jWNf+fmUcnegFYZl6crw5/15/n2GyAR7lIGtjp2FjUO9tnH3FJqn6KvX9iTM
3Slj4umT04bJGs2mdSodKKZePM2UbSbyxyMbxiL5vcyFyP/HF89p0syu5bahMTG1V+yj+HHyEI9g
c29fqefwoA7V9FyrqojtcVcGp3H558LglzH3MwtQyY1sGElO2W/UUtiDG3nuOMfZOay7q4kX3CN7
nUChfmbmFKX9c/tGDW0R3PQpl1iio9ttFcD68NgHoiKyhGewg7uI+UKLedjpC3Ds42bYrbEYT+ot
w/PODxf6ioJWMpjtyDRuEiLbbWOBGdceKb9JKRJbDhYeZ6eL3xbdiNxUKHl/PQxHGMDR3KYFF06H
L77O3POdZyX46LV4AznWxmmMwrU3INQwsN9AVkFhEhER1NMREx9kT2wL6Bt6qrIuti3armaKEawa
anGS5tykUHcXO6sCI30OubTIE8TJpg5cCigIaIozsaB49GLHY71mowJjqpAvjI/eNGOtVIg89pBn
vIMsrxARqjrkLPvB1VdFMDjNErsghH87qGaOgIt5M3/smFtG2DMw4j8Zyx1u+DlNecuMBFZhX2qR
ChMcXIUuyVS/92OawRYFVoRYMYeJDM2pPAAtpiLGyPhFkD0sJBeRvaaZI8kbtt1GiDwJ1ZmDJGFR
8MQ7ekvTMFnljckAgYw6DDfG03TQ3GYD7Jm77GWauCKO0SM+JODaz+sW2h/b3Mm1Ed9EP/zEakI0
hESR3yCh3sKgMlNORHOrUynP+4WcOxSFtXAtL4cQn3FD0ho1VFn98HjQU/gRHui6Xqg/OQLVeikX
p9gJc1VEs9rVWUhpll7RkICzLvK7roM7MBF2rFUpzdMJm9mUoknmg1SQPN6FeAJbSMnTmM1nowMW
aJQieoKBuPR7/fnIJlfs8xKY08Ow8C/mL9niIz4la3LF6lyG0snaOR96JPt1thqqCy2s22FDTGDU
rprejtd3KVhn7ea6U2gcoW+MZ9gVsXe5PGqjejmV0NSvlhO8KRRMAaJDyC1HDrXGt5cWDq5chbiq
3pwxCtyBCSeJcEo63zGq/TF1hV/gE7hto+cP9MLKpKXU0DCmAvA18oLka7qeM9Wd1ebeZyyAKVTE
/oTN36YHb7/BAht1g5dWw0qNTS0d7JtCnm//gxylhlGCOz1rmqQRd0IWlXGvn4exWQQk2T8Nr7mf
DwTUfNZ7XEeSuLML1I9dLsBdZKzIJu0FFPk6SAFYoEOPFu1AoxXxPep+ke85M3L30egsGV2CTmit
YNDVVzRikoVsFWR5+k6kyPKVBWi+5fCyy/pLpC8uPu9M3iRmGElosNRMxQlXwjGQp+0AMIl2mirf
Mj9xX05HX/X8i8mgyAm6H7rgznvq0GHrTmZ45APetpDXP7snjAj5AT4KzYPWrHZLnMDZwVg85Arg
Eot1w1g09GBrBIEUPtvKjdQ5dheKPllQVLojCg89xxVpvPHAX7+TMPrQTlbLcrmc6nBujXx7m9rZ
50S9lNoy43K+7yxqc2/9jC6KoW2zcDf2itaLCtMkxGEI9p0sJ6LmT/GKfyNIr31d+TIBSzg96cqR
t7bDTI0peyjNTZv8lfO5HV6G7JbctVZDNrl3gMCE669DzmAn65jcV/SPjyxx2OVwyjHy+DKQunI4
FVuDFgPhMOps4Wf1ZF56dQ9PMVqZflfYoFJ/JyUnD5mVaucyF7Ka+5p2WdfCvMccRnaZb/5UjuFu
BUqwlWuKvlINgFjrKwDkCicU5W9+hqh16iktZIax6jivMyEYU1yti0X0JSdndXtfZ4sSQh6pF3QZ
wUR8hv2BlnYyfIYjZcZxSyfVyLRgE2mwW/dR0rQK90vwyTFWLz3eWS/hpQtHzHDo65SSIY6f8adN
m0iQsMliblYbNTp9BdBt2SVEoJqZLELCfBMQ6WZvz7Tf9rGnStTyz7Cql0JNLqraqa7CzEcuMOl2
6Tpz5auQ75wQjHXe+5Y9XGyYhfAIuMGgBeOq725cZjaSB7Y3onFbBFO58TkPCcAUt2AO5AloBP3O
3gytwFd0Xu676RVX7sFBdX2ZMl66dsP9nepHpxd/lHSLsp+2GAaNc12mVmAstV0qwQZbuZTxBKyx
RF3PUsOwe3uL5Gtp8ZK6G5xwn52+v9/jvvk16ZN41mQOQ8OE+rQoijmV1pGJfUDIIYfoTOlh7wMO
F7c6qdRPneUCNlW8ZiOcass0QBenP7uuQOqZFBwEmr0yrzukO2/++3PFfs9o4+tV2tvgDD3pvLxH
XJX0/aIUBzvOneAbzQBkxn28i95Ssw+rDU6mEPtiqlYCIm5pzTjeqV5+qVX884GUbp8qEK2fCj+O
hrZ8O7t2guEHKkvNoDy3Y1cnNwwcHkzsflkyWdAvGf8RgUTpEnW2bctR4nksoLFTf40WiAX9ug15
bLDXqqafUNHu+Qas6QJbYm6eKahQCJbJA0FE41J1Iy4dmwdUX+isY9cRo3AEKwlOOHUt3k0wK2aQ
AkuLkrBzhCUAU0lxCwalJjMY7vvGTr/ys0ChPkWmuEy/ENzGu/x/S4Nc0m7PQqtTbnJEqv3O1Roh
LTo2ReYjyiZZ+4CLPU6ALQytfWUVHfGkev7ilHjmNl+zqW735OpTKE+s9lGgpAQVQi99auvfbczc
KLh2n7xW/AGixzE8m4S8tX4N1dIx5XXV9RpPne+HVdC54tfeSck0DTXnGMFfyu0Hzg2CVFGghHsE
TZksDTLy5jbMOoQl6x6hJXaahmuqaNJ1X6yQffnCKfks15BIr986YsnMtX57xg5ZZ6ffJERpw7Tp
1fdgTMY9L0XXOr/9UROjk9J6HU5TVaQLnjUFOgI1Wo/sQvCmAM/kzc2H7Efh/wPg50YXA2WKoByQ
Fj0PCbGiuVrqavJircSkWiCHENGD0l2wGI90Gjd7W3JAE/LrwioQhThAPBPFKzqlWO5Psk7dxOLh
jvcQoyNGDmwiLsxeUBBkWC4R5yJTML8L16Fnlv1khdphqWNah3djMIjaXjQbr3FUPbYDrDISESS/
paWKm6+zz2UEQGkcrTdui8+HirQoY04QFzHlf43IOHLsbf5s8tBt44flMZiqYYkXsx+pCA/mb+ku
eL7kAiC8oQqc7NyEcZGXzLN7/BP01fMSf5tu37Id97tENBOfEEe7vSw4Xzbzv+p+wAi/Sa+B/yj7
CP3Z5sVaAJybj4LwwRRHlgcjKEFK9AlUCO1zq8GRfcdTJvIW6tEZ+Lbob/rBJ0mS4oGM6F4l2RiI
8Dp2MKImdmQe0jkIbwIyRNEAguTaiO2H5PdThb/WxAtX8HHUylaEwFKpPJ+aGTUOgV0jW1o0QekP
cWvpo5PZ23KGBgWhOIMDZ2coecHn3guU66oFsoRL3DPaT8VPEzHPYDRv5CuzlLYhwrAqpY96okbG
Duckn28pEjqJXKKaSBrAxwkPRD4dhg/fB1DpOUSb+xPCbz2rdi6F02d/bDzqDgPywwBLwXSJduS/
US0vlatz+NIa1UzJIvGYAOJb09pG/foYwKvLfutxSt884vkp1Z4GEJlmgU8Jv4gddXpjvqKVL7pP
Wjb9d7hh5J2nIO1pI6vquqKByMB5DYriWAh4c+pQvp1GLx1XzS++I6Sqtum+F6YE7UAJ3q1/PntZ
E9JdcPiqzodjRw/fiywPAax0bAXlggb/WC4qbY1d6fqh1LnvqPlge6cUcVGLuKma7JHPLIuz/iJr
2n6w/lfMmnouXX16E5sYkKWCdGYuK2yjCogw4BZbVrzut1xGIpxNAuDLjLM+kDz3xi6blDsKNjnf
5oPnmFQwFW5poikCCERpdOlgHECCiWkyyxJkK8w0aeVI8jQY6FoT+8q/o8xQ7b2kRp83xQ/q8tMJ
b590yGyT11UWai2tWp+hsZr2gAdSegbyz2vtlcwrahEj0xKVIWyqrml33u7laXGObCsWdi1SkyXz
qHYzIQkOGbT4U4U2fzDwuVOp2nW+pOFll2AIXbIDC0aoeSDzsHEJkQYOXVCRrhQ031iYiauu4KJv
H9G8Q5PdEFFzzZyF5cZF4b8g1CCb/vFWvxVmC31nm553c5jNNj6dZAqCwpOzMOeOiwqtfAi4eL/3
H7+BMOgvFxA/OkZTj8E2+6gWJUdCx9KAbpRBr46qz3Bxoz0LTqR7g+2dD1iLZJ0FrBeEWvhHL4lG
0FlEq9lny8UxL13fRL2g7VmRA9147jKTg0bRCqv5zbuK2uZN3WQorzrUOYr7xxY3Tjsm4iPXOWz5
1acwq+fjkBDFmq4niDit8mu5PvM1hsLmuWnbNn1QmSirdAY2dl4cSuCdokHYvfZje1Yu2NVdLNcd
wLX8byYRSASqLk1XU5I+5MTnJnvb5utA1Bhuqbndg4ZNYzzRCM0k32aAkL/YoNBNsq1BG6rKGLkw
dSI8yy/P7ijLsNim5nkgDJSCAczjKUkcpMdzpt+gJFXN9UK7W7MaI7Aolbbbctgx0M8TjjaytmlT
Q/rZSEchzW5PmVTRn3NYCPeYqFq9Kvc7fuDsc1gyNzaOvkPyg3uCCsRoejpOG2JrgxuEfKApYsTJ
Wg2YRm4P4eWj5EkdRAfFpiFPCYYoxFkSnlFZCEkpRRtM1yuYtmeBnJU3pXxS3gJiRwY6XlWziNbG
tknqm0kOL6rl3iKPEUqo3J0KL7AQzYHPX9j4ypwbEXGZmj23JDOwpufAfvbI8bwni56oTCwO89xz
WjiGJtU92xhPtzbLYa+hzDNFXnILT7tUkQV3RHqSi21c7KJuuCPkW6c9THHf2/olbYDlpyzDVylD
InbgQGxbVYwGjGs51d3HcSqbtaBfOB3jWOZ+WlDr6+4BcOz42hB26vvjJtfIbS5k64beK2ROEls3
md3g1JJy82VDy0Dh5vKtOHpt6o8UHONqvZDWl8bwHAqDiTNMSABKKCJjJpZOBj4opcFOknoQsnmC
RnYbjqnkRXphEpaRj9DsGjnMAcf9iJq7N3e9NfAPmVWpBFhJv1L1mlJoLJmtM1zszBcarX+9cFbd
5kanNmKw5AduY/ReBCAKg6f5fWIuvPrToXEYoD+qiJrhij0RCwJU1P+lOADBvOxXuw13oM5qiMS2
zUfB6M1UJSYRf34d09cRw260uGQJMffHRtX+7EdbDdC1ciiAsv8OArUVh3++4Qkq4gHwjQIyFF0/
Y6hXDqLfPnIHRsUxLPV2nuNlO85hq8zOpCF/4vvfHXVhhC+kMf2mTWP/zh+cow2sh39Pdu9nlJ6m
jC+h9pFJmUPKozsIqq+WHAjzpAkjFdt/MExwGJSgFL5WbbzPKcbvKRsgKFelaR2aB4wSYabBYvmb
d8bDP3Y3/0QapHfLv3GM6FlbKIM1vyLT3S8zV48iAVFmPc2dxGkM3y+ytof3RVzmVw1X0zkHSl2v
lR/F8BsdzK3PHXVJQpfLbhb5342d/W774YtK6PU7gqNqhwNXVL27DU99jPkhitCiprt765SPI8yn
SD0jV2OC+WJizrGZL6eW+loWN7g3eftH8Mv5+zeo5zt5Ofmwu39U/dnvuM2fwWFxLT4KjFGsQ7u/
Vzu2VD12Gc+uKJcIHtstZ9tUICYmmybBwPJYUqmvroxemSxuF7X2FbrcDlgBZFHT9JQNCEBOqyHU
87TLeDs7PwEO0JmxQk9lhZxlngCH67MbVwo9XvLCl+EmC4DT+e34VMQ2R8iBQ1a8L5mmtBbWfkjc
cbU6B1gt+JAo1Izfohjslp7i8G+LN7hDZ++dcwjMgKmMSKMbDIYmotDuAGks2ZwDX00/X09RZTs/
3rjiHfy53t3hPTNr6NpY9GB96gPKIQ0EpTDJ5e3YItsywiQCHe6gnkRcKywOZCykQVNNUZthhpPc
i9zB+EY85bH7Eyfzo7HoafmR5hgaBBW5gH8ZnjLntvq7AcHosir46AEb2R/W3ezaBh2Le+QZ6dQb
X7xm9YT0V11T1yh5BqUUs/fKZUvOhEH3EsUsQ7w67R619Gj5O0iKCKXmftjPdospKCoomn+0WSvL
u+vDX/FobxslVuPoqjfhwcQ7P7gW8RZvnbVt+IG8HPg+cvATNbzLWh0WrhC0JUrE/ca+znlfKuiN
18Q8mzBQcNOy/TLCLdCV9eI3b023q1GXTZPMVfsnk5FGmUQUzhTAa9Q0bbBy0fKtPCvCAS75ZaF+
pmE2JwARe1DdQMhTdpIBjoVSc/9EFjn29RLu0M8qPcRLZMWkjJFzv4CLJYHujYZW+xXdcZgrsJcl
GBo2YDD6SYrOelmNyqURjY5nKhRaPbltFrACe9dCGugghvGKNOD2Gwv1e9kHdJZiigdEqtHZouQN
KVn9139hYDBwvXgpCpvKEs1pjD+g+t9PApp5zdpBWngcGilp27FVwqXupvGF/3v+vhpBvU9OLnTG
k7RsA54z/76pn0WGee3feslIMZgoM4Wn/qCVHds7yHo4Bj3h7c5fAsr6eQlWVyWOHs9WMn167RxW
ro1KRDToY4XIOCeb3bGE2gmWUyg5IUrdFF28R7QHnNYoyhid9imtWVBz6OBbv5phCiB4kdNzCsdb
DOvu3W8Wax8n3yw7tx8U3Ub/b94jXX52aR857BWcHU0uNNNr5a+I/p4YNiuh7+s4JXIjV0uhyszP
E8sGF9v86IkNd3sxNv37y5r4BYd1GRpxFt6OvuSb9ipV8xef79fRC1xW/EKk30K361Me0oGuQWZt
eIqrTsdjKgVJSzGltUO2ocCq6ZFkK5eQ1jkfzHcNpvG23DdLL7xQqag/1YcyMnTIyJ8FTv+XL0Y1
WAUzqu5iKEo0HqNSHLjSsnAmyhWwNzwLKg7nZronFD61n+306PRQH/ldSH4FXTSk+Xl8ygD9tDlq
+8pDxuHvYgMW6xqlSv0maga09c2jtkLSpSYBSbIxSRIy6xphh6VbdexLfucXzzQDKyr6oLGGPs6z
BHMtFjVpg3UrgUGQiwPEEyFb6xdlsmtSYP51Z4kyTpt1eWwn3JWs1wS78hMpXO2lpdgGCMPoYMtL
MTsy706GStHkXwhi3RmBMxlsgXGZbQccwhbtCa0z0juNjzJs1JDaxVgOPL5TRBj9MdmiVizpwN5g
I7PoqG5YgsWzr2iXo9Vfl87VnKrfOanQ7N7ue+Qi4o4fK357VgLvm5uoBajAPSk5qkscOcBCV8Jk
l2+8bk2juPMMxqgqjfKz7AenPlNBm54/IjdLn3wTgtYxnIoe8HH8QJuiodQQK1y2kCR8OudcaCp3
K0FqDDsZ5E2Qfc5hrx7fiUGkKTzwOyaelB24PblLm34JEcKMA7oN10yNTh6SJqlbBtM67hZMze0L
uoAhF/FJJGmDU00zvPoig6gw7tnr+0gy70I/73TVpBv6Sig3LOSOcgjklekbm7b9ii1SlExgacmD
toPsMMGXLhFFodVZJ6SpI7f21LAm7678pQxE3WiydV4eevjV27RoTIwQZ+yA0I2EF0auctE7Yup7
lqC/36cu1Hyl1p4EjsrE7SjoHne40qgw4Ggd/EpVbWeUyWRd5ohgb7cJe60MUs/+X+m6zil+Z6NS
CZCl7tjtT+/4zJNQ+F5oGeN7oewVP/mG2WC9PLjdWapYXwmlw5Wh2ljgfAjxGnxgVuUFiP+Kxa6s
UV2pmZL8iywhwJswDUTme5bRFJO9KBl2R9HoPaB1xmb6FvlxY5M9VX6GBBKPH+bN5zXgxEJgXIYD
Wpc106dFKG/gCAUXiUzSCYu6DRSk/6/U6/0+JwIIr+hH4ZzKxXjIPtD9ZbnIkTkdkskLVgaUGibF
OMcWgKd6+R2sAplavLrBr51oV+LKMj+MBJJALb86IzJFOuMTvRE8Ge+jNu+j3TYBQGqO/pVt7GcJ
+Z1M4QllA2IUlJE45z8gNJYm3PnOE3bHdXEXVg6QGIKudwl/rotnKFdhH7wMFZYi5rp7ywMVtBlL
KvrO743RfDU2b2uIYtbqXdLwevTluTE6xhuqBTlDb9p7uHUbVcfoR7sFAs3sndx2BHtvpWm+cFSo
pqO87QAZ+hYK+XeGAoFg5Ot+GnJwNDA80aI/6qxX0gy7BXa2vgcO4xN422mCkMa50ocFei6UUEJl
hZtNMoXGr2bSuRzdy1A4sm0Xpo/hTB75b05rXxiAxBk6wAaaFK94AW2PgpT4rIHmACQNe55qZl7Y
FzDTxa6Bsu/IACihj0CnEiwmcPc/OIs2HRXY3dbASzXbvTPJ1P88QMBx3FzHYwx0jOWYBTZQUWvw
zhP2K4URJnPYW4rXP1Wettm/jhpkwXetR+OmjvL55djn3Tv5+dYlqkVNHbBaNFp01DzhMRDS1goE
Iss6r/QwwdgJTDoUsp3wcUraMD9EWosOIp2LdqKTvswEZ2HtZY1egz4gZbnQHu3o3Nc7JlhC90jI
wageZXttG+z+cnXMGnDKoyhfPwl2klE9VVxGc2TCXN1mZRSPcdb+7duBwEC0bR5Ep2PUtWFM+Zfu
lDDPP0DhxGdY0lpQUQIPxATk7VuI5jhdJvKfk4mhEdZkIqpddGsHpOlSh2HcyR0IyTz7892qF0bI
aNGc3CVsz/gS4E6xLpVzToPjYhfQacGtStVWh3bt0u7tt6VQKCry2bN+0GPrkNZnWDQ0HJZovNU3
7WS2qHwQ4P2FNIcZaTR1WlsoWiU4f6T9wos7KYwQrcQBTkG/or3UjctOUWxTIfGyhvTZPlDw4bzb
KXOV968+My0BE6M11ltF9q4JlzRCP+jeQEzsWs+Mw9rKC58MUYal2wOKN8z4QZ9mcju+TfTOFpAB
B7HDifz4a7qfc3QjHS2thznL6BSgslFwoIOSkKMmMixQQTP905XmZPGU3QfBVI58EDGcVmYU4Jyj
so5cifQiAyaK6HG0+vqPmkcHaoNK9EBokkHkqs5L1LnmJGbC2Rhfm15mUfQ2ZOnN/OlDRIiM/eN3
aGhqZP6uYje9Vnry3BU8et/QCg+NhxuLa0glPk+gWSPcf8ijf17Efy721ZHTjilPCnZRI1aYgAf4
c39bLdDBlAlmyiWsWJ4+v+RJBnd31nmvM13Qs3u39iWpEjbSvnwdS4dfrklCjmyzEOFtMVpUUZXj
4p0CMdg4m9NgcP8V/xwt4yG0VDQy236zSMhSRz0XGLso9zq1rkJnEAEKmIaAJu/VyN2Jv/skOTML
NgqoPnebCt9rSv0q9qxRk2UOXS6dRr7bY5OYU0biwv2nSCgbJ7bi1htLn07a83QiQKvLcmyTVgRE
SAYO8IXDD9n959+PaRqa8BIdOwYQtqhwZ4Wi0JFzILJIUq/5ziC/KrWNWUtdlJZnocK8ZAoJvtNd
XoUEWjfu4exv/nz/+oAVTyyUSF9N+JbeQA5TmZlY04skTRTBUHSixNm+dSBu8LwAIck5kwNFIWIz
BqX+tUo5SJX1HFPyJLN98HW7LGmuRrRrapEi3zH8AzclxHM02BF2uBVtIepLDT6xeO7hvR3JdVJI
CkocW6SsSho+14yERgaF9FZJJtd7v5wXrpL5kZKK/0qX9Fd5hxVdoz0Umwk1NyQaNbN3ZwXJZ9YB
jEdiOtc19X9HFR0I8G/tHV2WW4NYKlRIA2LrTYpwRHAFEuCIeKTdCfAn9OeJEoZCd58cUzgeNElp
s2TQC/4VZkgLCHmZOOLnHkBwgmeK+6l1FAjX5ETWKGrNVeS2S0L/sCrNrMtzSfaSx+elanjXzmYo
sKhOzz3eSycp7TUpb/8IN50HrRusd3lRLtx5Xj1EY+58fhQKKGIZ3wwhT2204z+UvPLLR5s4qgTc
SYOXBuMMFRbSydoarZqYhbQbN+KaBNL3dv3CKSoXD+R/Am6KqgEuCpA6qfuKk/MCSD5JLa8orLXE
CefO4X6u8iuXBTSqxQtgnM6SOcthes0qZJzVaq14p94RF4Bp7NumHIl5cAN8jneDRG4L8WWvcCq1
5Lb0DZz69X30EBo8XkbSmN6Y2x+78lhTUL+NbJyEnfaMxWNbtBcoVGIjH/SYMHP2CVEDYz2OPtuL
c+CTI0pWKbRkExWq8O1ZIT/QtZ+VKQs8YEvPaPmVgZUaWIiOF+l4GtINbOxnPybgnGbNPcEjS6Lt
LQa9KPtLNBJRObvMF5ypkYP9Vu1LeZh2yMbYgoTeu3m0CAx3vOXJVwgQpxBWCDzXNS3fFG9vHJX0
QhXsWuUH7xP7YPjvhLUKHVgUP5WQA7MsJp1NP9IIDv6N5Iyn8p0uIEV5N0P5LNL51yNqIBbppmS3
2pRDHhNKMGHkmF1BxQZyOkmPmP4a/lUITLMC8Ku+GPveJAHaXTZ4gFnF2Z383CElDqeHRGsv/pZR
iTGW5LmdanxhMK+ricKrr2izoZEkiNADP8LiACfbcRIA6zsr1O/CNdJgUPxI7V7bICq7LP78bD7g
B9+MzbNVslV6bGsNUMb3vDvQy5Ebnr0pHk7aRhIhBWK6R1VNODOxQn22fp6SPj+MbUr0AzZFG2Pk
Nohdm589ANYKd95j4WIHUHfShv8q1qARCYEvu4/KM+BIPnujxRC/kj2fi8zOfDHjqZRgQlfIVPxn
IHg1pTP0Fz3xsFyXMFiE8rTrd9myOVNmN5PnztB/Og2u8luhXoEk3D5Mvv6/9iAEfxO6fLMMpuek
N5CUOHKLn9vKbFK1zL5sHvFkXhEwdrBL7zfYfUJ8gxojjFxGrDP2LL7cAjbwZqkw+coSuvEPGSpz
vcFkhuYksu5d9eULVg/v5aadoAt8DFTFsPRO0d30OMqjrWTAW3jXXZGFFNQOVCc8fsHMBUt64V0K
+O70TKTy6FKJ2ZClaTC84jwNboU7IEZJ1JyISRYL7x/Z8HFGG+KPln2gjqF/Wpxu3k+2yFwILrsq
oOkDk/QJqcU9ku3ADt9WPtYuDkHtw9YCqHNkHVz/Pcv9uhy3YywrfTTGufGwCDyM5fWPSCavFlf0
Hd88/Zl5gH1rrnQglXCEetRabqjl7HJA6tZl5UklFuUcvH9FZPhtwf+jlLDeS0ztm7Cyw9vI+9qh
9d0hI//9fWZihKFyyz5jlCIXThenkHmniba3+CM89hJlKU2N6PTCOcYxjzQ1gl30XTqAhJ9rrA9M
mZC2ebyZzmtB0FSpvYDW0uuhMKMwZs11cl77kDmpcfg8NdDjY7e31scANT4zVzdqan/c7Lp7WGPq
2OCVSDgGHkg9yN/b6LhhM49f3zcTeKo/y6bK3qBnfrFjUGgQpP3cEJolcgVERWcj9sonfHE5C9r8
ZQw+JhRzwf7v88MV+NyCEZXqQhvpLKZ5NB4UoeNfnlDONsy4vI7F5CvxvDQYKrpo5jFwS+IiOfmz
/cJfThMZChVcA6o/V8sdXlgpeypWjxaR3yw8BotUlGo49cy7n1vMfMZqiAMYp5voq+4kdwauJPTw
hDoptbSEqw0EXJnbqkibalGBYOf6OolJdB8Ag0yQrnqhW74rvLzJI+2UiKEZF/KJ8KTVXZn3vq3f
XBKMTfDUuLtRzTrAvo8EMkFk25dLKN5nabRBbinCKNzauvjMAZzCX/dLLWjn2jP9GfM7v7hkQmb/
U+QJCY8PxQtf0+4/8s074LO9r1bahbf7iv9Pw9RE8e0iVhPvgmpaTqzIpggDmi693d5uay0j6hPC
h+68F7aTSA6JO5oZfFL2S1Po1xRFiQrJQtq/vzaLfoNQw98WlYjC17y3bUxZH6WxQ48xBwuaFz9/
RsTyOFNONdGzlAN6bs3+kbKYmE/Tl3ccqn97x5InWdUYNc+W+HjxxwVGQM6tWEVbB+ygiqHCXvaf
94rXjNCVGIiy5uO48w3Z7snYd/yNJefcqAPOOS+JuaghkfJ3stOOxOTtdK25NHeKBAqNC/M7crx+
tOczYbRlOf7PXxnzLTRmzxDAGvQ9S5tlb5rFCykD+nRZmKIcP2wIQl3JKtpJ+3s4V3viNCFQy+sG
3ZpQJ/xeFqP5DSfJw/KqdREYjFqpAdA2OYa4irsw/WV1W772tFIHWf/nvTb9DxBQgDNOyw6x3T4i
IZ9by+sQnA1VCyDphfdvKuzypcfb39XjGDSRlX4vj0nGuduEmIPTHPLsR8Bk3PFk1F6jbuhgDhic
lSh0UCwPgQZsIKAlvZKOV3eYdp4krvCSxP5dE9H1tKV5YWFkW5UFSg91LxlbNsZVyIL3rJwh4vx5
hNTF/jYSeCrrpLzeNx9v68fIQVg+xgWFAfKy+fO+3hM+XFuk4vIhKctz8MkfmTFQolt53FMpdzHT
Gh4xGdRZoq+r7W+C1LhCHwFRk+ulVydDUhgRefRS4LD7ZQH+ZZkojKAXrtVk9+wf1oxWrhaTaEaY
Njae9crhWtIP4JsqbwiVQMdzYczyhsU928Bqo3FFnqH3qd04HZJEjEPWtOAGZ9/tAVlOHnot7Jm3
BtZyHbdmkHpgHEX0zYnwHB910h7zuBKqfgEKgjDi4cBa2WZU8V/eB95wnhofE6lmvp/9PxKlrHXQ
BfZO243nCXMaN3KT4DjUV6xtsWFsNDGb/zlPbF+3bhz2rx+z7kkPM5v/Qw94MAY1Lla3LyKBWEac
9ZHyR2tiyGRqxEAOj/sKk0j4VuiOyk0Zulj5C5OekT4PpPC9BYp2jJzElzsZGDdjuoBvJn72/ckQ
AVWWizdzkkhubv80tHry0omguczdRk5JxA7cBT6x9OJCcqnD6bRlY1D0tyo97dJdefAMCIK8vO9D
WxuGyQgIOI5/QWck8d/QMd63ACLmdPWvKud7Rml9F/I48GxeqroNgsMh35Z4vKeoAnIsnumiSUcO
XeLpOcTiyX+/eCJxu8z4Epj9i4/xvuaLlU7atU8QOni+CmSOaJzHCM9/BNv85raVIn43LrX5zxGk
gVSgGzTGRz9wo36f3Eod8QWyq9/f10hhwlonafJxkZ+Dx7YcO/NhKJAqF+L2KzIpXQsjZdmvH2HG
BZmcjBAAsnb9CtO/spiMhOiSmPT7pihMVa6ie8YEgeN/YO8C2ssbUdqo4nT/PE6GFoLX0KRgmqi7
gu35BJGztixom4VKTmlU+p1mqEr8VkBSyp09l65Ebr2BTV3PWDv2e8UMErh6exQGM18S6URaIOqY
fOZSZAbLN/izY4/Rv9YoQrcd5EmfiJoD9DssSlVjie7xXWvZRCQHpJMCrsrViLxIzvJcDougVYI8
+RyhddHtTaxybhEg9WysxANvU4c1H4mH6WV6uKZxts6m2jK80lJ+iR82Vy5+/6cf/mQEBKZDXc4h
p+iAe5Lda7V6QClIQ/I85kBD8ni4uJFvVW2BLDz5BE14Eaqxp9KsI5xhJh4Xflz+ob3j+9txLlbU
4Z1jZ7+/p5xj07wBPpl5YeC0F9pHR5uF22Ahue1LDUQzC4MOIiFPjbA7Tg9yXSVRXCUGO/KP1He5
vynVh5MNJhXWPF9Gxax0uXy3mbSY6t67VwAq9bhntXQhxxGkGcDrPdY24dj/02WII2dayTNW6JqQ
LddWtM7jyinH8AFTCuF2VQluxW4x8gUvEg5HOgI0HREGxh0aTSN+uBGoaS5J7VxPTKjm0/CrboO7
92tq/ofX8o6alH/64cMS1giqA8t1MCgOZZ1Lh190s0Q0Ou8X8mVUsQPfXS/5MHnhm+EYBBVB5UDt
jYIyqkUqZtvaqbV8auPdKb+2y1Dw8aMLDSb1eXRotaOxmNwL2GATmvfiZglqs1eI1cY+SqnY18y+
TgGlIhCONUHAW/NK+9jgOWCb3FLT1K2uc1CGXEl9XbZyfkSfy4a2sjN0k+3g275MNAxZjmz2Oxbn
s7LpoL5foMXY3Wsz4fVHnk4yW3ggbihbwTm/nq6kjXoJmRGFa2nQ8Ek1g4L9jjFpCtxt7aqXQG60
w8gpJwzRB/ImuKo4zd1wIuitxQJUSLohortXK6poPxYvhkcJj/k/Le3jN+ZbE0vYjmDHZQcFFEmv
Jpoxn9TI5ad3nuHto4mW4JTjRp9xSfcCLY1hH4zqaElkmdLjJU7NS0CDjD2Cp8vEe/yaaheyq0p5
LNdllv8p0tPeCDP0gCaHug/VhVHZDGgZ7I/U65WiN1tqIEsB1cRcSFvwp20iwdmRmBzX5bybE2KN
rs7zC4PkG08rih86x4m5NkGszb1x2WIudUm8O4dTvDAK7WCL14O6Uv+0XA9GkVDRf3bBz2/307Q+
PBJ5yDeCbN2LF3CkC2NFc4ioF803jj6E65rv4RTVSQoCz47NpYj8SEuEI+/Oz7IerFD4Z+uGfDSw
M+tGMy0oS9JcWve7AENBxDFf4CbTPYIyth4EfcMp+bWnsj3cy/3uFnWKT/wDS9CyEwAqdWWbBM6s
rRbFn9qBZLvSIjELp+WdoSZu592Lk9A3QEH9xwv2wtFrbwK5gJnG2xmylY9UdOu0rhkMX4oj+X4g
5H0nvy4fLcEMsQUTMTGlcLQYJospEVa1J1GTZFBUI+79Ljvxy6fqz3laRvydHCJBMv5mw8yt57ZH
6eUVNu+eXy0/i3hyuVHRt8GBz+KDT7QBaynHqQrL+/Y+Fu+lN21fVU0ffUvR10sXA7PHYu3nxgEW
zmbR2C9og/zG3DAfpd1H2zcrKQ8dihO+O6j3NfZ6VfZNtnonPbfYaaFAOueEmv/zloYW3dcMrI9q
RhpGMHkQgqLzwmawars/LNz2Q7KP+Ilw9OCCKToLNRwpUXj4SGMOXkoZAVcEWPSkD2MlnDcrpiGg
ATaj/xk/mDbS1ZvKk+BKQaOwqbhGbLaCtOXYLMNOQHv3F/PxT05qQWdAk6AXeQ5sobEwgamFIAGP
KD1XToMuzLa72LWN/qMvan1rKgpRWBmgd6xc6T3OFxnPgh+g7fPtr9cvRLa+rL72xh5cp4YVIVSu
kMqCss040M/A5Aej0VsE+V5wKHBFe6jnDSAFOrlLujT8EAEH+dIBYB/WU8kofrh5WLesPd4y7XtV
P5ol31JTclRGMzZ80rkN8sIgzJ9bJIuHayUq4CPKf320eMuGMTTg7zI+XmS7aczTfj3CE//eKRwB
ASLxIzC+NTLphr/CD7W+0UFDcnaDJhWkWRnVGLDIAl6PnnNqnmsUwEdPcAhs0+LLrWkAVJPB5b+T
RgTjAxgVl5pZnkMS/crJxlsS1RTnP5DcktB4y9JCTL3+I2e+eqzdMugzjyP0fJVZCeEHiePJ9emz
lqzNaMW2edMrUFEIVv0xKNA51cmqGBAH4j6aVnvilwYywCNnDdWr49MIxCdRk2G+uS5vIG4Cus0y
z5gtuUA83U2+deXTbZZcL5F1dW5hjUGLeRNGmOtWkEl5r7Rs/+hqNQzLCjnhuPsOd93tq0rFUfVs
ArQs1gc+Fl+h1uH0XCGWJQ7yzA8wpdWyHWAzhLOAQVAln8r1Co8yRVytVUC6/uozOpEtPKfe1Czj
1+vLFLpjTcI2T1x0KybE4Y6mCGTulDQWw5Fxa/MYiJE7QDXs4xnNaF21raQaFgODKNXRJ/WcR4I0
t+LC22IAfa8T16E585WUSNeZV074IyLyfPejsfQd9IdIWnoN4b0Vo9o4Xl3DDgcw6Dc/U9I3C6AZ
2xWdjZf8dYi5h6ASETSmPTFXthwXIB6h9ghR9nGmAvQwMhcnrIzsOm4a45fM82WoxC8jcj23ECu2
Qj2eVPoJlnBkRv1RbHst2Pyspmggj8JBmMxX8UIPwNwDNp7FxYPGZ192O8ps5wu8famXQ6BeqvTd
VDBxP14OWrLXNw8sZJ0A89L33XncwjNfWN6LY0SXkUZawX43z8zuklzbQL6wkVsOExfWaEwBsD12
6EGzSJbyToXK1NCR+ogtddr0TvusjTKosvm/nHKSigaKaR8P+4AJwy10AIdbznuUj+zmy+JeM9Ni
5u9ctTztouICTt+9O3PcWO077jID6RfvAd/CWJ4CqNeySwoKrC5sV5BoaomeeVwccmZQzHLuX3or
7fs5xWfXV+FZXCdfysCQg0G4uHKpk/D8sWFNQ3WPMa0mRUFv4mbY7Pysjpd8WVZkC6zCyW/RQZ4k
p/ltSFk1zI/Mlbjsqc5ILhAuuqfGnOB4CaEdGkuKpXzjr3rsuv/wgg+swLshBStTVkBaMQhSCYv2
GwNg9paqWHIBXK3/f7MZAKoy7yTyf/yRKWorUfWKghTmcCJ+4kXcMAbgSE3JgRqAlufsDotIm/zR
O2FkLSIiHaVDBquLqPvwVcH3mJLmB9Tu8oFQsxor0H10pScLkhljMhf1PI/adIYW7UQZrOizrOAl
0qw0nNfzB3Bl5YttBn2XySaHBRWd48Ll/rrO4uFP4eJcqONivsOU+0uJ5gJS1pUEVBAuTawdXhUN
dc+z894PjwerPiwFgNqmcJDi8UwsvwKyp7a6MlIbMlapvQIGRNeQYbdIY/0DBOMXWbwn0yiNormS
7hTQ9FOYkq4jRBsZOmH5ZjLDeV2578OS+vLZydWQbVUx2ABIJpT5qVnRksIYA+JvxU62bHCqoHMd
rkNwhsagX/n7p0aTgOZajKbdvzO6Yo9c/DDCKXcHx1SFMZDzN5bJM/2mnDirBGwY/PCtDqoXrUHE
8lmHpVdfvAsn3y3etO/EOHu0i3/xShBM8k91bWX3o0gwiBtBpjaGsHwmkokaVgeYN7De3wAaHucp
tzpMOP3g1DsOt8XJ9VO7keQc2ktAlAM2bgYEW3Xq/j9s0jlxENXrRTnl+pSYM0rzhz0jcJnq23zt
ltIAnf73dx7ynzjhHYPudE/lVCils5SlHpFz9jXaJu7paWdMX6/NhTngSe6xUwTgUJ/hxX5d5CEt
5umwk/TNbEuYtBoK5KlFdB3/HBUesgP9dvT7JoT0HSbsB7eDhrAhTCp8Zoz+MVWa4mJ3u2ptg97K
DRJm+1I/n0dkVoLNhLx8NHE3vqtSVm2wG9sQrwQIszRWXloR5IZoYchuyAhYiBMM4IwpEgFBK8o6
57LRYr+vJiyMHZJpmwQcY7C3i05CUiuxRkGEEpxKsNQxamPx1IY6vC/jDEbzgT8Qb/HAWwQ0v086
49ftsxNkvLUf7g11y42VdubwimftrjW7spAZz60qqn0owAvpn/+ePKH44EAC/bK5JMhQOIlASp49
SnCJV3ZICDs5271X2ihyWnT286W5sJhdmht6S71g6ncOGd/6GBDF51TmLGtE7JobsmfFlhwXwXuC
oWE0FX5iZLP/CGO7rJsvd1SILT3NCwJdF//ue7oBjkB1j85TN/Jorjrm6eR4XDQFTJH0RTztYNvQ
LF6RtleZHMDi2LnUaIsQrgvoFK567X6Hn4itiSjmFVInlbAtklUc4ApQ8h+RyqJ7b9esG0sQGpSr
F7xNV36CHVCfjir33Z/UHgvfzF2ueYf3YGa4HHJNvtGA2bkcECrCgzVlCuAwuC4LiukTaRqA51BA
m3giX4R/ahZfJNezeDhO52QCZqyfMQenFdSxrD/6B1ILoEbMM+QlAEg7++JN/k4yTpmyQFaJJ/ff
H+x2GAXYlzwzcxnslkz985IAXlp087x1kXVqnIJ4b2wS8X+1YQIjrrbb3TlJlUB4M5qRsKid22ym
iklsit/BXqP/kZXwe9Z5s7S9zicKF8dvsFwKmQ10TMQzV2KSxVVUtJNNv3wMFqmzWLab8QXGr8Zu
0JwBGFylBzrN7MEfhFwT7wAx1u1fhXGdco3ooL+gm1SF4YpeWgUAlTCN3IA+shVj89EXSzuNuaST
2pU7YZ3VfSgZqpcbEpicKXp76sHXN8s/wywv425+9yQ1vzCedap2DmdB09WikllwZjCoBK5Z+Cjh
2v0XNCKsa9kZ06eE+n3vc21uqZVMg24kxUE5+fVNLWZ+j76s8qb6HKZRj5VJj4ddVPBAg5DOrMR7
s0XwRFNv+60cf6hYRjkMiPccNxiayS61lpp9uRJDO/S80Mzr4gJpv1Z7+jvCGI495H3lCzsno7N5
IECQWyPCGR//mr9HsaD5ZbpbROlkyfIB/sbWYVFXDNdyqrZGsiqGm7d/FdxH96QkEsLc5rLRcazX
SMfNC45OOL3r6BmBQhHFv5WqlMa+sjP8ybpzyfaMo47EPsUDyn8KDyMB0Sm/WMckj0Dc28OAMvXu
9doXpPA00tppqYw8/peegHPISaqnElSqrX3Alzke+w/jgBG9T8vF4/LuIZoXQOqUgijwIxcHpGDk
FYg+3Myl1F+jxkxUg32jyGkw6bZm1O6T2gb8/0PhOI7fjw4ZJXjsgTQRU5gUt2AYmwCrolTMp5tA
DH6Ys75p5pGERGTO2mBN4LkZkF8rAGEZC2b94qqHv3UkflW0YqQUVRwmclwc6eqV1DG8LYbvVBXk
4j2W3UhzKUQLt6N0mcScg3e7FWtFXtfeD/0M+RNhgy7IVcGbUFTqBMqFVn/zjsTE+v8RVfXwRNb3
/+LX8HRuwgWvnr7ecSuef0RUiIXQh6oydMKtfFGDzF68rMuZjaaiuYemrDKvfzHOdxgCsdauSg0b
vSVsQ3MaMJM1XpOoTpJzba3mrFhXStYwaO1h3sn7ghBnTgKWdN7pdzQwTyrkv4ZGylZ125ccd2jY
22Uo4pL/Er2iNpkbYHDEvlDV+0i9KqvSUtP33RQ7MeR0whAhUYNnEHPisSC+du6aPPeKLgNOPK/o
MspaVguGRzhI1+Q/D2ELZkQ/xsPzdLGOGEQooWRrE/3QKjYWetZvVg7mBBIm+PqUL+q2EzJpdDwb
K/ORgK310dZPizSQRc4Ol+magYQFF2++qrJEn1l2Iy42AwjB0piKLFkukSPv0LQtisxFwfSSjfIA
QGyE+rOvZlWL3NAsc8anOIZyttgFk9RQQ90EWdBEiCPcp4M0eV3FPuolLFEttC3kyCX/nZlbo6GL
CGsvsUb9HyVWqPUMfAGgx0LWC1QDEQPnrmyUy62HH36VpQ1Y5uKGCWiEJZNn2vlhJyZi0ln0bd0o
ssHbCRA7g+8PDaincXqjJe6Nov/dR+94UFKtcWdf/xw6cSXefzlRxROqnFbBxYbPa7KpgcIo2cM6
dyn7ADO0fRNC5B5sDT2fiWrWOQbbqJ26r+FADW/oc1/km2oJclH6NMt2gpKWgxnarndKggZiJm1j
PEq1Ba+vzBbmHaN8vu9DQm0imdwo6it+JtWvI+EYFjuGrqCz4rkHnaewX+sKAqOphPGyQ5iVk1R7
LWgq7fHW9J6aQZ/+Eh7F2qTOGE5h5xAQZ+uNpkYIJpWJ1wtqetPdRED0gfQWY1ugFsiR10zAXxsK
RRNAAizZcXPiuzJyPeSQUV+ELDWg7OOMOxuy4c/BnrQNI84STQmMrDso+qU4voq7FN3LZeMvabYr
pZ6JgJonjO8+ATviYQX35q9rwRb8v5uaM8BOVEXUULLP+L3pUdqPOpZhawC4KeV7YMdyHsN7GPZS
nRfGqxhaJ+KMbKOz09ENmmQD10QPBEzO42VM/E8JUAwk0+2jHMjPYPqojyVoDMaG6bB3oHObSLUb
WR8viYoPMN4pohL4p+QKda1xN9j8TawgsaTWsi7ebIH1AWcQE/Se5aIHsUbwggTx/hq1Q02yzHJP
lvLwhiwd4CuDJfCaBKgiUE0ZlF2T+KRifByAoX0NWMKXZoh5jICUrArNA3qNzxbiLTOObTYwcw2x
D4McCCsfg1TPg0KnAJv9VQCAyfFndCFmZwzxjJrDsuxsFR0fS9ycc9UEwsMSdoUTphJZ64px8U7e
GZTA5wYNCeg/5Ry0gA5tOxmaMBh64TcTSbho2dfWGb9vjFuR6NeEIUZTpNky2c/3Gn8v9dsMuxts
uojySKW5nbz/DcEkaKz9vaZUKblbunjpBl8wgBX8ex88ggaliv2vKkg1+8zEyJm5uw6k17do5v2x
X1dP8wnyVYF9c1Iw6fll8Og2SI5c65YC1eUm8gZBbO65XfSoOzPolmkv+cFvnUciTzZEHuEzIOrd
Y9pGhQZvT/qp9m6u0kCv40WkUKR0wtYQP6Ak/bwzh/d1hqeSFvRUIx5KtJzOFB0yGqcz/aQ9fmEq
CeKDlyCJn9Unp1YnisP4Fa//Ou9efja2ajbs8oDCfmUfOS/1pXrVxX86eJQxeUjJ7syN1/zYQ3sM
ltRVxY8rX3WkdVxglCKIMJbBZCZWAUZG7exV7m91uH5+QPW9npM8oUUzn1nRaT5HKSTfM8edWh6m
umjCE6Y8Zo77sof3l9LUxwg0zWDKI9fsllZzZLaRYuk7f/g9PFRBnFxta4nCDxlJsizGWNoMUlml
eHKaANqvokCq48qfgi5yDEeJIMyjcfbZLSIWaFljEbtR9XIRXKnt122Pag9OBlc7/1sXBf7IMhyg
QYOwPCEEkv89mtWejKDamE314dynZ7/S12hSHHVvgARtOdMKKtyq9Fuv+SIHHuA7GluZTAPll7sT
cTyqKRL1CcL+kzuCOY1vnHyhDJlDxbRGcwDtiB2sz1qXF9gLC4eDwGOWuIH1l8aqJG2r+cRo2UkD
M6t3xnnrZzJL92C1kEiI5QJT+TFVXjoSO2h2gf81AbTK+f1wA8MP13gNT/aPwYXRRXpWjBZQYFBZ
HE8w5KNEGGI6UFuLHPd9xzEI7DNaWehr7cEdIqHeoECagGwCz7Zx+0QTmCQdS7gWDy/Nhy3TKmgT
1SXAaXvm5PiKML8+0dOAeEjMWsRjUcLaARPs/IJCKiNeUwdaeXBemu9oswDFwocI0gLfYWT07DqW
9zY4GZy/HdDwql7DmXRrZo7lI1v3WIo5RDxTnmf+9yu9LuUO9Faj5oq8hWHcJRBgkCcj5OizJBmU
xpDa1A+nH5V19s+af4QmtJ611dYDlT3BFiUcTuq+M7lBeb6m955y8nNmTbC6b0kuVEE4CCvSKXVs
5q0Tw6QbU+8Yju9FGkxScolABwkE4lhj3y9KXjL5XabZfTKDh+bQ4HqRsHq/EN9byzUzifmMctMZ
UKkf88SZhaK6zBHRLqnhsoCYnGH0nTY8sgIZAjDDngzP0RFk2KQpWP2Czh36hgjYiIVfy4NtYYMP
Zm0SBCTRZGHNGkHDdWXvnBI8Es3cYvvbILv8GP1kgEAI19YGvAm9HgTbJPXk3pLP4qN8x9lmaQk5
sdFIVjvg/Aj2KE5OHUz/7Alm29Oxrx1534mEVEC+kkyPILB3Mi/FYkDlVkhUM/YpH77yek+7Dk5r
IEf4S3RYFgGXLmmIolOKtb/tr5h40Q0I8UzMANWAG9gcQf0t+RDReSbf7FKKWC2yk8XfX9X7ID+T
sGbDswjwIVZAXBGG5cw1Iqfy1e8gS5FZajsKQxR9HgUZhr/qdAT4SGHDPjq0GONQWxuya19ateaO
VUBCuck3vSi0O11Hx8RdP9GAU+9QYUuHemDADRadcoA0hgxivIkoLvONj7DT06yFQDH8+Ysn17Av
22Nhjue0BLTaAn3lTH5TX3Din1RfOooWPsxfwjwz8s2e7Vf/S5OvxYfowWgVI/MV20DF7ePbIDMM
qumjEpUsr0JFeQ7kpKW8kxQcHF3K3enohsU08mXCABSfMnalK/JTe7ZMdsPA7/ZiZkL5Kc1J/Q8o
NCAHEc3nqhKyTMj26JPTf9CMyYwM60zn8o6xBggvASdJ00Q8nctXGMJHCv+9rVV8M/9n7/WpiBqY
pEVhaU2HmaS2GUEpvOhUq1OiuyxBNiMZ2rgbRGLRBsrImgDUDzM6SYvGDfSXwWn8RQTf/ssvvZ/6
5DhdCLDozcGX1rumm7jjPcuBKXUPuuazoXSWQbUW3LJFajy6ML1eyM0Mu/P0g0UOeWOoI469nXon
FjtUw9RWDaxkM6KLXmk3SybhWvcvWXKXcBZJssO1WMYLZPjB0Wr44QJlXyA5H+Xm7oSJJXTUIO7M
miaKNOY62IQVLhqz1xhSqOwtkfVl04EAwx7t1ZoBXi0JOg5Jh8aatbcrdZV2k5pfDFcFMGFE5yk8
UkvrVShFEvjzOdfLe96FIqQ0FkM0+czeyNE+QhP/TGMt3seL3xsxYqbe4HrpWsWOPvdVxjyPaftL
xp7rbRhUbGRljMzFDbDLI4M2Z787NgEBGmicx/0oF6tKQdzFpjuKi1yL7AsMLbExcJQHELYiWMOY
D9tbQt2Owik/6AKzIyVqlsmRQ+1ynTKkzIUxSRvq+TIEIHZ/4Vb2cIEPxcVY5SlT11T78GYnSPlN
JBh2cJMM4h8qAxtM6nb3ImREZJ3SZ7Q2ITveyhJmy4DXcgaPMp/8TYk/NIyvwUH7WWUziuYnaBUd
/Xn0flgHdr/bZwaSjTJOH6TfVYBBjWn956n/SFOk0Qu48pD7zFi6+shSquqZPzCIHXl1hywwaWbs
ziLt9abm7D8T0LpBypiJboQs/0J6+QGZrgqU2J+/A/BB4AlYbBFy6DgJaj/aHIsHsUViPxHPnZtq
NLEEF7gASynuBz2EMFu0eCrR6X+z0B5qywPTk6vJfuHzHM08KaFoip3etH1Y62FTrifwE45qgYxC
EmxZKRkXFQkJG1bbFEEG+efoytrkwPZhmqDvrj50OsQ8z1SaGtMvzjO6rLdaLCG9Y7Pzp/UzsKHu
MXNDGnY0Tyc/cXRGAYoF8JMffpqrDtd+TgDmH8CjsG+3cMIAwJR63jNkEMJ84f3Kh3mBcJpRou2Z
+GBeZDIcEBrW8TIqIM+foZG4nxZ2PNaXIa1vOn+fWCZWGwabDUhK0am8hapYEkjU+yJnB4DPBzWD
rcMj515jNJq1v0oY0nK/L1Im5mJL0HRVvcv3hBYM8NHkgVhM2ewLmFBh7Q9RcWRuyKrF9thHB2qI
SOn1BJNw9nxsknfmMwPLPKaYDSu4koaHM6jlqMAGvYwALUmUiPNgU/C4MPy9vLHPKiIBZC0g3n4D
5eyL4tv2kcBFH95BHM4vBK87Aob2R/S8VXt8wNbG0ZXA/JH1E4xXnlpXVTQU+F/RZWDW8jfrV51B
udnThM2eiMCcAKnThCYXdcotZA2WDY+HBoypylewrBSNJldEfKCCShlxos21rR5OOndguYrH8/DG
iB4HtLEqg/5xt8p8QnwBNio+WaH7VhdDDyO6uavLFuZyb1seTMliLFOJkVO7yzK7cMppuWKPNeZu
Ob698rU41iUp1Qf/BWi79Q9zbVs+YH8uWr/cnSBY27CmEk/8jL9btSTXER4kLdICzwpjJCSetYNT
wfWm0oTOYT7eydZjevqtwq6C+0sx/OSw7cWzv7ZZ05U5BppCQCcNddTi0zx1K8yFwWTw8xp5/WOG
0eW1r6syKSl0JruNtwzMO603PEedmXtBjGOafdNzlnc2m0HcuYkSLQUiut2kSPd8/jS8D/zsmxfx
aTlAskHo+odasDjzvEz5TB46K5h/MufGnksibm9kK8xzCQUtasNWrq61Yy9L3M+oPNAutJc+QDr4
bjhhBjl+Fj49fxEaO0O8G2pInPGu3MpWk2iotuxsBIcSwf6i6gHLWQgOMn6DHyksPQvQkgshyTni
JTJkHggwHc3a1M7tZdmJ4QllIqOVcKF+yA2idbSVbZMjpwT3DHPQJWZkAU6CQf3oOWxnF3lrV7m0
uHo64rbVBgKjb2sd78vPeMJjjaYQfaht1+Bk5ogTFVYjEXeAKCTd5kr6lUCMXn9wBQ1e/g0IOnA0
0+TxnBv9PoxUmpSJRr+Yr5QxU8KvVzTaUeSXzXvO3D5t1keDFIJd/HNid5FcPMaihAJkW2mKtLpZ
1euevRDaAS4rnjzl9MzRLA22Nsz6z330z/q7JX8KV24j8wqA1VxTDgK5NvzXRxsc7AV7E17WBN1M
+yqafPx1vv5s1w+AFtXTZYoxTNmnQsW3LjKNcdoT0jAiyXAGq1JjAdMUQOThckUS2X1jkVkUM04Q
3pSzIrSM81L977kGR1B2HBQZelUgH9O6rSOhE3BLuBst1NeiYIAmbZCbRglHNpbzaKY7B9yjkYOx
oTZNT4uQZeMWTTdMjpM+Vf0yy7yJhGlGhromLrFpfymq0pCVY9cShMPWWydrTHYYa5dFKbL9v0vh
qRKHNPnUlgcj/2N3AZQ3OnHnDfxofOLU8NMAbli5m3LwO1StMFi+GFE4y3nHWvlEI7kdo298pAav
rkeUx1fQrkUbbW7MJH27XynC64hO1am+XHPGLX2ejpIU5qZKW3hXdu26RgudcKZRPvaMS3c27bAT
GPx5H0WPD7/Y5DasS3nAsBVmoWeIyF0BX1PiZ1xtVgxDM68tCUAAZg0ijGEZfsC4Lte1JIC1mEs7
VgyJ26L392Yvj6J7b7IwtyKvaF5Ln4NEWzmVEInXnbIx0z2KKrmIWuufhOswYTXvPymp2IBGUE7x
z4fHo+zRTeS2GF7doakiz6IBmWITXxXekfZd6L+G+YbB4mHlw+JKkIQZvzvk3BjyO9zSLfTlsLh3
eQ5phhbI+Eaz4OtRDEPmTCB8Xm0SnAgOEPpHuQjZxIHaTA6geC+SEJLloKE/4Qk6mTjPn8gZ4B9w
BbmdCz32FX98ns5M9TdSIXqWRHmMbCwN1Oa/40w6NCjumIUs//YH/UpnULKHQWt6j5RFTmWtnF6F
ljgqALYwOjRfn7u9MgMaXAnoTCzlL25TLH1j1aVLm3H3bvDO1HoNL8BfPXViDdrqwEQ0IojRDItk
PbuYBZqDjgHNk3MrCr1/4IvglIKO0lcNECsphBgxHVEUNcMKubhyPpIGtWuJ8cFo3IrBZwEYsOpW
c+dqPYrbr+MqrGZKO6Lb+kvswg65ZWUWVsExIQnZCeJitZ2kpFsv4XLH/TSyz4JeCjGatNMUsjm8
mbhXRhxLvQxrad1mm9xZk5in+/lGkQ7ANc//od+pPunkMOwOA3v4WEoNczqmPTPOODVIJkJDk5LH
RdFJfs0xzUhBsaifhxXW1TsUT2kZa+CVjOLIi5ahabcopTrDYiLA8N/blxkNTlJRWLiQuVWHi3y8
sYr2cYHunebNS7QmM8giffmNOJ5GSVahe8aRjnkk+OGH4yp/7pjlFlpz8eNl3iaq5Q4D9aSNKKBA
Cjxqt1WUB5Rxs73YmLGCLAvEWBbEPV7TyRAoUUdLkE2cJkqR8kAgYmI57GtUgeq1pm4tT4I8qn0h
3SSIWtnV0tmKEwRnaWDPmLDzu7YnTsgqCrac9QaBmGbxg6dm7fGA8goH8Td6XXtntUUvNpIxBp++
kVGWrcNQvB2HZYxu2x7935WAOCNl9J4xGla7onhGP6v1NvcUnY/DDG6rV/ePVPxKI0P/SfkRdzNG
TcKQbxEOnM5MB6VjzPVZgn/PsFfFMRBxET5CF7on6RlRomzcYoNpZ39I65fZDZTJzp9HgdNf9Zck
Rc0k+/U52QeobzNtq7xDAka4dI02U1/lOHZDN1ANvLxkEMdC0UemR39CXcwkj+c1JH3lrSUVU+DH
IYdAc5rreXMzblqpMTDR3CJIfy86pPLaxdBRxv0p8bQDv3GqVudXZFDK/wivPfPA/8TFHPqwUjeB
3Pde84BkDfFYKHrSZS8s1VToCOIJy1cqmmhQeH4f+Mv3xD99bgtrGPO4INSzHZYZikl9/GoB2aBm
2ZcPi3/JebH4ZDVuHHwBgXSlCui+pFM7Uq0pis+b9MXDpf9uG2A2n4v8Sh8mMawkbzSjAqSnwRHA
1tdPkDQEdo0YXy4XtXWTzWnY2RbIhJWtKQCt+pOLA5PHsipcKu5mWv8QtvjP8fzgiZSd46qXQFk7
civJDo41vASLZBfJoNLXHEOR6A8MLhqO17gwO8nGjJlUclYPTGDmPOODB7l2TK9GeZUmF/nuUDnS
VZdTC754GLhwjjgWHFgVoD/fmNv6HrNn6i5BCBVRzui0C3g5HGiw1+TDuTI7pBzHwE2fmAWZtf2P
LuUZ+qXNdSPaMyyn/qTUY/8PDYQy9fSLYQHUvjCsRvpINZKSd5PBNabOoxFG6dpb4xFNEvCLL1Ro
wjq+UISpPC8vixNOYV1f0ul/nQmUIXChuPma90ibRdfMqmSbaJUq/XACvZZiDQIggzwjdn4Ymbit
efL0pA2lzee1yzZz35bhYen8zqmvip2fYdVtqebRsVgaLOC2gDtpZyBALK/AyhJ1E/BbzMCkD3TT
bVAfcqeyk+FzvEOJ6kZhEdASBaHPc9wFNOYOcJJwXeP4tKRU4AERAquvFywciiy2bmNctqYzlUe3
HZx5u25YVc50uAzgIlUDzLv1msj0jQg11whdfRzSIVGgYd+5ff1292opyZhk51qpHtMXbR/fxC9x
lrodrhSieNbT+TPKIpXBnTwHR1OVkpeAr25RhcCjp/aTQEvnEaRH1qRnSp7/nB8vRWOywWEDRo5G
nOx2/N5nJpEJeWTtGvpgdafXEjslF2Ffr+P+CRoFMBp3Whpa5RHmNOhCPu6/ZVIvL3XknMBUZgt0
UyHCCoO7Ya6dJ9taSloYeKQTfpeyJq8/E9QdGLxAqQC9cteaZiaHOyUQ6XwbikKHP38aC2w4MvUg
l/fkwHue1zWlw+LpdzPzZTcneDlqXqGyJ7f8bpTO95+pjh3gHI16I1qDNcOl021aHxWcTzAMsl7z
hmE0Ow2B09l9HxpnEenaOHsfy0iVBG8kMnXsRTQM8zPbSA/rLKZjU/iiTUGSBbxhUCoY6r9zOi7g
3AY1uXwPB25ECqI3MNEyqbUK0H8qgXwHOvLglF5YHPCVlDIsvlyliknVrlLrXOJ31INzJbz3MniI
Vwa2qt7JYxay+QFP1LPfqNLtk6kd3bdKLUYO/V7VhafhUDiDtLQBkx3NgrZhDB8kNrODqxOA1XeG
+LP7QnRjdaPu5sbemgnxrDRfp9aKwhR1pHOtDuT/ZZUQrlwbNCROvji1bRhgbFAGZYnLGMXzB+Qt
OOFk9sLSdmH9BPwtUgjvdllr6xp03hpg3HvFSyZdnoy4XZkJyyaZC+s+9inJP92V/0opNnEKSJn9
Mxm/JV92gRXcSpF9elBfOTnoA23xzMiE/kQxOTyiy8+7VZnbiYtd0Xp0oR3q0RITrdBUkA4Dg33W
ZFjKf3BysmuhbsrCZhsdLqYiPO1LrMuv/bxZzHzRZuI5V75A1r5QvfGoIeUQRAVBvi0gAC2+v2Of
LxPvubq1x4I23iq92HtUpKi8RVmsHVR6LFel689J7nQORPb5r4+QwgA3nzTZWUBh2CTd+1Tdxrp8
rhBH/1In3vAxqs3xzye/P2SmtQ+lBjkwzMZmvAT+NtEG+Rsj25vs1cx5hn7hqBOICTxFa+aVWHgz
jH36Wt73IYKAY2wZSNPYQlo2XiqDOOcYaqEZgHXjlFmg4PfbE1IGRQSwAxnKWOQtUTTsW12MAbh0
M2Je9IiMc33YeMTgnD6KAZK9jfqxcTfFsuZ8r0xc/UGkuEDZAOCBgMVM0zJ4b0mlN3tGVAHQZkF0
/Lgk6uxL73ON66shUkNoE3ZiFJp0KvykUZP47+9QDuoqub255mClYq5sWTRPbXC4erNEcoeGNTly
CzH0te2Yh0Ig9OB1tio63KTa/HPqJvQ4KUuW7mWOgfP38DOC8XZ96dYZx8b5ob9rcQ2eRKD1Tu4i
pfKp37qUTFPXrw3eqr1BfJMpKBjL5fpST1cLzzyWoaPO8ixzUY/9wmTYrn49u+FeuPvCHjtsdgyA
3P+85iHlOQTAWdJbd60BN7D/KJmAbmSkFgjxc7bNtIoAlcO59HHH1R+n9Zke919wkLyZfZauYwTU
IIt85HnuGmWW/qGIMgYzdH6YcLY4XND/OE3qcQyuDtitkhEOAtKYEdbDOthUsvKSFRPZYOs93DPV
mHQ65Osj+Yk/7vp4AQ++SmC7SCaNfRj9uyOpDzvRf8rs8bMfurXLByLBrBdRjR1C05fWXQsFaBSN
ymc1Z9kXDYmmC9whynTVfGslTKG+12fVyibw5AGGW6EqoSeaL0crYuTDxy8/pJXDBIdbqeLWZH72
8hSlGFuum+KTMkYRalab/IEjAuurCyTcS5hPSt7Be4VLngJ+rGxYaqpCui8hvABkNtu9gm1kTu+s
oR1FxgHczzmeh+iumeG3nRp4OOB1dzD9ffQBnci0X90hY0fCJG9DVBkG2WFaqsoavcKAPFZW6AN5
h01lGnfJBh9MNDAC+TzWRdjVXCzxaa22i5GSP50iWUj9b9aq3y+7exNlwqH3RqjnEqpxFHBkOxmb
oQBb4B4pTgmDoWP2XnF6V6B6LQnLjNpXWXFTmW/K9aOdwMNg7xYgo0TRO5dbeIO93jaf+YJY4tN2
QZI2q/2rQoEe2qCDV/k+d5VXzsdOPJExSo2F82kZRtgwDtb6tSd0JSWZ1yd0V/bVQeJEeF+aB9u6
uqY/juSd3C9xbMy8c03fYJ2sWkT47C4ZV+r13L709D5Kx1T+q2jlFT6nY51M7wvUDDp1BnWrThCD
95UgpLBqvf+ZkE4CgtC+/UT1j0dixhgKB6jwKuxSLAqGW2/OVIupmQpLg7QOsWzpQ9bb4bBD+sAM
CbppczhkXJQKcMI0GDVoM0YqHY0sqKNvenewB8UHHSXHlVGz7A9wgnsRmxMRZFJ5una1YLZOH28/
Wl49ABxs4euS/D8+0s5Lw+B8hVVflDW1H0v7s6H7vsLwh5YdjCSKfI4W254Mg2BXWGjyLbnB8r8l
LFArCnF+WqbwY+zJrphwgFtL8YObv1tuKoLuVkaihJdnr3YbPVCSSlNf6KDW7G/OMkoJ/3GhL1qM
KuEgnAMhIhkgjls65W25RsawmSTrTW7npw1N0aU8RSrbjTz+LnG3ta4FLmlboOr4w5ppgjObfnpl
C++NuMh12sLYJ1wGpVHde5lvXFEEqKs7JijyrMmKXTLgQfBZlAcr3CiBqsh6e49dsdbFjCk/Kvh7
sEPT7SXExZ44iFfkGBYR21uDLsnrx8ghByTIVXDwC8y9eEyk7r/kkI2k7pB3GNjcltOGo2aG5ODZ
4vfu/cdOUaupUbOhRfJF5dFWH5T9vy+exxrwe9GReh0tOwtN4rNuQIpBGZe6A+/O8qh1mE/lWcb/
dV5t//XuolYNh//C9HAM8f7ozsNItekavFEKpSOkZlBiwlw4z2+770VWUhTmaLxBdJXEikCeglbY
NxTeKysK1bqn0Nt3W3t0Rb0/OeQGKb00RPKy10luxRytBrjYwLXamWqLAK7rrciM+eEYpLQ7CWbt
s6w7KupGDOxFY5aY5fjJPW7HN0u9PSAtLHZ6ZqzSI4ZCXUovzFn3XJ9bxQg8Ah+IDL0V/zY0DLk5
g5Fi5xVs1Qvs6yqa9utBMrn49sqLP+O7UqB7MAgJ3w7KHYsZERWogWcAUtBxQzdMxGMhcYO+rDpx
Vb7h1ia5x7dAYNquYcakuDDqCs91F4DchE90QA7CdOlsKHY77aS2H0kbPJUmYRcRrkG2acEafYmE
Q5gg2us8fbP5M6XrkUall2T2gCG5jqbLDBvZE8qxWoRebMUvIm06FHqDzfr8ayRZL/prIu96CQDm
+IdoGVScjY9vNM2rDi23QHoaa4jn3XBAwkXsJpblYQtih3EgydnlY2eqKmWL3sT+/Ea0/Upp4z3E
VWhe4lFl6PkR9EAQIqKZZlmNm/Kd56puk7A+GyPLSu1OJ5mnkS5Et8247eyAD7GOkbI6uuBEABbY
222qyeZPThTFmE0NTDTgwsLlGcH5GLsdyC7e5DxFGh+D9/d+Wb7nK6zbR48w5rr8uOabSOd7MgkX
TJC8p4n08app5ZJJMUY/fC6wLuhd9xGFmwAphUYIrKCYziZpMwN3R5faDjUi5f/1fPm3/WbYEIk5
pMWUX7+iKRDzMDicMyVcgxkbfTukcOEShNXbafJwUsJJdPB+cyXys0p8/CEZ4Y5157nF8UjjbvLu
iNfSl2GP4X6mbxZKrtQCpYXlQIIyq8sdg37Si81YyZEXRwDK8pey+LKi6ftO+bBxsiLICu17iEDi
D/6SIjxEZvGwlXjnu2yZkTSLyTRnf8ilKq/l6nSNMOdZcUK+6WpYmWYjoYmOXCTE0hcPF+idc2/v
DTFk+aneVLNVCFYRUrhxGGURyfOMwiET7+q4wiZOJGRONwfEP8jwHRjqUTJY876Iu1PR2WWrAtlb
O0x4A3HSJLbpbgmCMAwvBxIO+A3UV+LIae93PTCi1G9CGG6sxguiNG9GRZfQvZg6hsTMN8lklYdQ
WpElxrDb8yNtT5eVqlPKJnouQYFmmoeOd6yiC1MqP5vL6DLFIxjlvNMeGVbrc9kdBXtM/6Yv9BRb
5h0W2DLWUbwuQ8VE8tgqgl+vm58u3okFVQoZOm13fTf4uSFthrq7tQbkZmppD/bzzFvuASv6zSCB
dHXNA/NGl2lMHfeeZNjHhLuV2utSpwPDtDZBkObzRnwIKfNrD9RkcEt/2K4jMWHmA16INnyMTvvX
ueED+cGQ48spvbN4bLoSmCYxvW9WomaKz9ioMBSLNupdIMnOghgMBAmCp2+slEbStTS6Q+UrPLFn
ZyxwKhLdRiF7a83KhVXBvwQ5w+CmyNy1QaWI3oQbirwHjPEWqTRft/CJaWduGp4ZsYw5E8sMdp19
jIDxodtd5t7b/vGZ4SuQC5SUcYguowQpBhj1QtFjHHzgOHSYvqOsN/Adif2FBMLK3KbagV1/vFxv
p6aGR+ZOdeHi6qEy8dF999xw9Qo1ub2rQfBE9ru8DVJ7PExzXghUbQI6zjlpstxmTDXQO40AZ8QN
kWJWkJwUELuEkdZXKLeQ2rGpC4R/bvIyJGvtxDIVQIBu2EeR2zS4ZczaKupyHzDF4Hfbxw39v4Ng
HRq+Gdb2a2ckEziLR2CIduJMoyWvUcCBiXqq1vHYLSMnco8shFktOMHFB66jc6b0BShrd698EguZ
o9E+uaK/fAF1vJdSWSo8ZjI4Og4NAXiqNg5qoieacPTxHw8pa39sq/LLjY7MVGZ9n22FPOQ5zDw7
85gGdAlWn4yrRmxGWmGq61AYioMs2l0bBIdapBhImGQ+GDTGyBZ3BF89oKcPnuu2lZKXL6sWTotB
O5hx2DRtqrUKcnK3vUq06rsYZIFyTvEGvbIeY+07cS4DfXtacERlVsJFGt9CW9w9oUoSp4jRRIDw
ViOfm4F/7l4TEt+cSCSVIy4QHmTQFJG68vegX0iToPof8SFePPsVUXQxKMAGV34HjUpfJtCigBWu
jggaC2zCBvYLHyL8Hs7oUZ+gjP10iTCMnkgtGwEpKZvHNlSK2O6Dz5lE6ag/PnqVR5VRLc2IlRT5
6ZMT/xh2iYv+P8+wEEw3iFSCqFMRa6aNIt5+boRVxgvlDMI5oflZ0copr1CasP0u1JqWtETpvMFm
wRz7sAX//VadVPPMdsjk0Ey+GW/LsODBP8PJLK134ww5GZApKHBeGaycML6vB7mEc8K9gDvm8TMS
Hb3QhH26+rnqRSKZrUmlupAGz4rELEz1AIeVX1WokhAD+i12dlUtSL9i6DXdZ57Ikb6fknSQzFHj
6xUVF24R6nQ5mgrd9QLQrObqyZzmCCyR5U0P3j+Au6Y6tXvOFy9M0gDCYMqd2xN0P4wX3hJwSbkk
Lb3wQTn0IGqEeYI8pkodIhtu9/YbqWQi2InRNNkwjRrfYiyJBX1NdE6kSco7DSigo4WTRD1KnN1S
UYgU6azD356uZs3WP4NUT4SC4Dlr9w2cL8wzIOw+JLNoqTuozHwE9dueav35rvHS/nyHzUo67vdR
zahAobFn5uTggua3JJTVdJyy1nZvOE8fRGu4Uc2lp4PquZzN+hFisvuCkZHwtqNcTqVKc25drvAi
HfZ4uHLX0d30U3duiy0FjeMzbwQX8I1/vlRGzI4W+vazdH/i8MpjIMXV/6sGEj99YfOtXxXPWLvG
AlQuwvarKFgFS2YaDcrrepYDMCA2P9IKPJ37Epp4v8MNF6TnmgQFxwKo2h3liujEfgbaJITxmizk
OVX4xLD/JtKv+F/ODsy3kesDJcIh2Mooupd3OKOc80qe+r+7Ok7xD7lxehlQLDZmzf1HX3aMX2V/
BFbHhmNhpeSlyqNHD7Bri7kPV+5r3Xi9SZFCLAZey+VleZcTqIeIUFFoKRviENWgWNhhLvIX2HM5
pJUzV0mVHcnIDuObPBtEOX/jJNQtpxv6j9EdZEaCyWNk7B5l1ArlOnN9ynv0UAJt+otyBIcfcmuO
AIb9KQPXyMPTq6c18iM1UfKY5tPucRTGT4IxXUMRfcrIZjNKbSjFFqqudZW87TFrW+bkocaD3sR5
gUePVy0jL9n6DIZ7LOusEP0WuacVGgm7bLtjIL+5IuYwWndXIw8dIDBI5+0UitSOfADewqifqh3T
b9P60pynkBfWOuoqsudwRUIxz1B5oSxE21+hnBBzi9Bzhje7ZpIKvIsAi0n90Lrx9DjILH0PKdSf
BkLpUf0rE2Kb5B9waZNN/4oqn53h904LwJevKbqeJzfMMWgl0Yz4/LIi2CN1UXUkp6uG5EwTaEa0
u1Nx44ssA0rUNhe9tJ8FBA970ZwZZF1dsEAgSxuMuJ1iIa46L1y86fwou7FKHZiAKGf13AKn6tb/
5x2kyHxnutzvBIxlZtaU7P+dKyNDHjWsGSGuIivxm6D6dfcYJuMKnWzo4CbnuVzZFKBaWwJt3ZQ3
vqOZyYi1hyA/Mli9anKIU8b8/OpT8+kkp2RLf72meaaDIFo/VrB32+OikGxC664VzIBCj9OKtzlG
qKnDY5Fu0ijt4q6hfxwnV5a04rMGCHw+We3v0kqCxDJX7Pey271BlRBjnQi7t/gXIyse+hx/yb+3
+XvurAQXNQZEE0pe2vlUJPaAPXugUutlHXhp4QjXZJU2M1fLHD/rDcuC9dNurCwy70N1VidiqcF+
9r9+adbugZI/8sp7BRSES5eWTm1VmWQOQktmcjbGnMwj29sNR8q7lSaCJi1zwMKRQAJM+gRJ9nfI
cW2AdVs/eQu9OfPDwmHYSFUH6gBC6NN4NRts/PeKZDPi9jpCB8MUld+A17mbpix0r481gsVPMgO3
QyJ1YbVz6+b+dnEvpo7UkNayojIycSzA85JQGVS5c3nuzPzCOF78O2V9tAuD2XvaFUjo5+ux5D12
+StNYuFCHt7m4Ltvak0GrwsaU8OewPUclLTpnbfaIz6n22hqtWTYorcuxdo3s1Mmim3xzYxUdjbs
sjCyoYhtFlxT+KT79u3QyMQVyYh8iTxeNgZe6dy2M6SrCxSz+SiQnnIhn4lRhUDkiHRA6z24rrZT
qeyayHIyiJHrzI77+Gn3R9YNseEt+eYjhgZibgUrtRYhNu0kRvEcUxH71EQahkVC8aHPbmw6ystT
RIk90vnBujlL96M0Azh/mopEcf/3Y+bPaNpdIryUhAMDl/uIO9X7zsDr1gHBGVLzgWsuJ+QUkNj7
XTYuIz1neXLZmFjroCX66P99B4gmNMMyvAUfaXgquDV5Kpvy7tyjz2BaVoTvfVndH16S7ZNE3tbk
opyKBL4/5RUkBfRs+bsxneW99jM+XxYbqqXnvAOKZuOXtCEjD6NngyyiYiMvVeO4GKda6eNLm8XL
ZZCvzVwO5JSq5P5IevYvzffEOGZ+vTEA8Gs2+Q3e7nZ9f09GrAfmHtgv/T5OPFcl+W8MqQJ0JskS
CQAlElINVdXB2zG150DPRgnDZ5P/lBZDYOzZn2ikLdTS34hhf5mx2mMb+jPutEMFQqkSiVtaRRoo
V1Ta/xZ6U5q5kFa3UGVzLnXoJrWppZlsJNH2+2SRm+4oDQhx8369g+/BDa1vG50lGAjH5V43V4g9
XmOp5O7+Qw5QnUUfBokA7gEwICG/Ag5U+/AcNaqAGPSp23JfFaUsYHbm65q2NUtSCCg5PKp7YQWG
00EG5yryb7RyLsUdl7mQvoTVTXRnmk+eSAhWSXymJ0R++ZRbk8t0UM+jEO9Ia51/VeWK9KZgydGY
5dXjwWqnzGV1DqYPSF5sXn3TJysqPSBHU4XO98G1ABDXLYzDKnrnR3plSPmWRJkZz4to4UfN8zlR
87aH2qT0eDDoqxDCwXaB8bhX9ERXyl6FqtbbZlSCEdxt4xU8u/kYoz/DsIRUh6Cr8Ra72OaU44Jj
K7nUhcUIRidVS3jp657Oz+atmpY8aLzLC8skwxGnuWJ39phrWcd4E5gPe0b3zqrHlkoezb2fh36i
yBeb6rok/f5gHxjvjNUDMIpi7Es6xHiPzzwBgtY6p2dtZpp/gXa2L6ABwo9138qeUezzsFlGJhuv
1zD167SVaC3NBXvlX0dIeiNZDLrQttlBPmL88fzgANub23vFucbxPv3b4SkhziI8n45CyJbavbuU
ZYvP/RdfDtv7e7FHn1JUATmkJtRCt/0EnBw29BCKpPwmKTeNyhIZoHl6jDddhaM1MRQbMSJzYFPn
oPVBuUBOq60s4TzK90muRxjzpmFu/6BjCiB2Ar4cXeg4rSiWD7LTeblPfz6K+Q3SULsM9i3R+eCL
vH/QZ8mSNxOxqP6o3CmzowFXtuUdqCIAMl4ef8GGuS1uyw9qE276bBJDghpt2KUzfjLugOyybXWE
TgyMLBCVPdgCnYTmq3G/ErhJ7iAAGNWz135oFAfF9Uy1zdzOOmxp2sUn3qTx6aizp99c5ByWw3z3
+xtsSaawshrsTDzaVDm5nLo2/XqNkimvtVrTiFgHrO3pskRcTS0lmeWvM004xwTKRNeYel12CLc/
Ms0V9x33i0Ls2myYNvlYpTlLOCA4pLfgUwoMhdHb0b/bhOudsRCFOuz0ocBC27vK2Na+FXISaJ/g
EZDK4VD0wCRdBSaOU9zkA0Uiokh6HpWZaXuyPfVkvT2Se8c1eI2si259H4nlrn4XOv0Jv8AYXPhR
eOshAOms+7Wr+tMZUEjAFrNfwmXlXDaRObd8bfnlAXnNF0QIOATdhEUXzvYiTpMJexcapZum/cJx
N/kIQb6X3r+fJulJsV6OzlV+PiTjxVeoOfyZzeEuiqe2O2l0xjNzTiAYBpFAz75gHZrYK0BA1FqP
xhoT/h6p1C5T+JjsTf3q9crtslcAQ7bilfNYwB4XLx5v5KekOrr306oCFRxsfE75opeIoGARe6MP
mf7qFnOHtSm6ItB6yBPc4NkYs2RQvCQxxYzM9Yu7J0VtO8MmuAJzuRCMw1SKAA8VS018eox9ru9u
sF8uYHc9TYc/jjsr48MVCfTLBYBKfygRmrg4GQmM/RU8YGuoFQZ8IO9aQCtB1qkLcBUrKauy91ci
xywxiYXkiI2JUkEWJg/s/ay14De+bdAhrddcN/wrCkAbn40olyt7Zy2J9P7QRdf56Sn2NRl0vX6I
L32j781e1mqyz4Xho+k2KVV4lGJH3gIr3hdsJgLK7ycAra/fZbCFV34zFaqVQpMoOcRgYYoiE7KK
Ts9eC4KHISOhsrOmznbcRQbbnxKG/W1awthEtQzfszOhFx3dw9HWYFSlhJ0cDtT4RDqd7N4rK4aM
A/OU/BHiyEo5JOyGRywgQ4J22Bb9NUF7uhWsRZYg9ieHWteu5Naialgb/nHdOfR0qgWOZiDLM/aw
WKDkmsHnskU7UFfFySrs1hsAEKqtW63fq+P8GUgfA8FaO0M4obHpRJP0bBOaJgR1zYlNS1TNcL2d
SHyR35SM03JNSFeDHSRkURjrMnSyvRUOBabMn6ypPjBvtZQuHYWxD7SuMmmSaMpCu96SpaaOkPhf
rDPCCuX/itzvAey0MhBl1Knrr995gEG5RB1+ABc+4uoazv7B3HGwXAL5eR1fX1QzNjdMMsTIn2OG
pmIjWJ8qfjBVigpMSqX2ADkP1OE2rH5iJD5TLuEmlPyMvm+H55/h5rKrOUavP0Jjj2JxA2qqwWBV
FUHPPQQxkSDhvoL2DWmU3+yP8qnk19V6uYL75nJx4Cu/wY9XPUPOPAYE00waD7mrWwQYXWMRDzPT
iyhcWuzgswQd/yDdjQE0g08Cy3NxiJvn/TGEBq2g8Qv+lcjwi7pj4AbWOW2LA0Zn2dfiCYxX7Qmq
rbnGwr2xalXb4tfb3BlJVZ0ifmQeSlNIJlwKPIr/Kpt0sO/XStKYi5ReRcTSBFdXZwo8e2rgD833
+FpBp6XG3dR0Ffa27d5aBkSgSUkaMnDaFoMaKzWBqlcIFfuzxEn0Zr/jOyflV0tz4Nc8aKzY5N0X
zdQjHx+bdP5ZhmS5xyKvo7ip+6x1Bk+EsBwJtDlGA2ovywfwfhVwS7w0Tdt0xQKulcqSmWY80I0T
NfDtWjsem+A9NuR+5vdMTiFL3G2hxMjDSKyhtlKwiYNQugs7hRv6NjQBHXTuxDjE9ugg8cSuluyy
F4vK4N59G5W2GR8+bwNGhR0vTPSWFEE8q183RvqgEp/t0R5GEGW6KiGIXEJ1aNPc+TSCEPG4e2UL
qnTpnF5lQLJOfuxNsUF1haGoXA6yogacx3CE3OUx/Wec8GtKjmOw4CGQUesbDIIOt6ap6u4qB5Ji
4Vlm7oaXPGKmfqDJgc+m05vgGqx4wkkSPJlc7bYK9+aEZcDzg3iabaYTkKodhmelRxGBC1z2Q9z0
UdaXIwAYURalvkluUymSIMWKMa/Jiako9hkgE9IURGddyj7i38hNEv4M4oh5c/wTJybF/5Eqr29s
nIgDcTUseeE71NzcvZrVCsb7ahrFt8xnP9i35S9oD6ml4Ji0wzcqZy2/c/8NdFItUGV87AlTQoO8
DtImJ/+6yuyTegr8jbJNv8v5FV2zT8SCx1zUvrVZ+SU2Y5r7swg3wotGjilsm5DBITgz6U70ixW1
KREuaqFof953QFncmjrvm/H/eVHL4AAfPvVJ5n6FGnlc6LxOegh6c7BUHTuB5z4OUAhK+kBkH41m
GGall55ZsR55bQMTysLIdvD9xGX6fwl47Acrn648HKYmUF4fSLFjyx4mlBQrqaEqRe462NfdgEXv
9ITSdpUnjkBnU0hSD4YenpjGyVW7SNteac/N0IcY3/VaIUKnhGpBPxTOUz+oX0FObYP3JhIbLCa4
EKKME53EPgL3j9N/wg+CHJsrB32MYqKUbVZ9h+8UVMmex7izvPBcB44mq9ZIvN6z7a3IrU/oYOzt
oCGkaBNgooTuWX/IJwRNRu/bLRt6WNl+WKqd6y/XxF/oZt5MIQF8uIPsRnwchIJC9IhpKH2kBvJq
ckL9e4hiCNvTsOqpxJUZXkiAxiLzNHX+GbRxrlD09EoMtzBsmtpX17FSiHWoGXVpYsZlke6aG+9V
fMXMZsHG9xaGaLORx4Aq2XyWX3oWYt5XDqv/tkY7deyb5bWhSXt9Jzh5bNSsfQWY/MtN8ePyHCp5
FK4th0TQWsN1UZ4pInMvIrogoSvPDKeyyA6RVaSCOtVABfcRyDVnCZokVZaI1OIhO57VaOz6UZIC
/WZ9eH7gCIVkNj7E3CsmPyaA8KXMbIKXmaKMDjsgcZ3szW6TzrsiZYIi7Ks75GLLi+cNmz74gigB
evakdzNa5cJgal3ujUCM82gXBimg2lCaS9gqShe9JqTIYXXnCiZjPTgtrDgPCxck+i/o00B17J8E
t3hm99O6xc714p39MY5xJX267zAfURRfHlIKqhYxli6JN4PVdKMhU59EuISRsAQ35eGDAR2fud8z
IAEKHzmrDA9cQVvlOaeCidCsZHWNMkyJQi/pVrvmcgUUc532it2cu0z++CuT6OdvF+13Y5RC1xHB
AJbkufE1urrtn9rH6WKtTnzGzzW/+UJtsWox1C5pElBp0HIFEN0jZ1C8l2w1NiLWFYy1yBOsgb2p
5UuXtqybe59+wTMFQRrVkbI0DzBTVBh0d43FavwrhEsn10iji2ZYKKupS/JGEn6V0ghkW9HGif9a
2fTbEv7WmSnz8gRXXWLngkLvAzbBW5hQ26joMbD+EcacX0sFQGkGZM052Cy2u3tGCOH8edNo1Jrv
PC+vyTG09FhoktFHcORhXfFs2miMXoIq7+Jxbt8TYOuyqzro0tJxxWoiyym24VB0fxxq4ConvbK5
59gmEh5tGqFiqB0SZ8WhqTF6JjprFlygny4+ptYzMVCsbQnl+3xKj3pencFT+PNc5u0/L4BoJLgy
e1um6XCUK4DGXABbhsUz40LLugCqOyRTADs6BSCytT9B13imzdQ+qXvANw4GGvY3bzprXSgWXEVm
b1Q9U3Lx3oD6Tqb5oEjYV6GtEfh7TpEg6swu6PyHVW7wCW7X29i1FzEs1UiNekDe/i6eCzPdCFDg
x5zb3w+Jbb4LdqIB7IS44G2xRqwjXFsTiuh0ye7WGb3fR8mZ+Ahwb9s6J8UX0wRh8qFWfBPLIvwc
o17e7o7NA6fyaSUIYGztNe1BDTdS/OzjV/LjAZnW46xsxRhNJvqXgHcoVOOs0Nkt/hvD+vCapA+L
PwEBgFYcq5XrQ3tWkPjjpNucsaXJ9rm5a1KKPQRfAUc9+0ckZ3BGPef0lQkY3ysI36RQiOjpNHwz
8ixe8Z325ufRjGrej5x502RQMC1jf8OYQCDa8PiLmM1KCwPDcIEq1sVgIBxyRM+oGnBU2DlZtwsH
CSI9LrK0kv9MJPa+HvETwUCfuYA3pyVAJt7swLCSH707cldy4RRu0BIvITjMjq5FYDcLuetRFcga
+vZOKM7BgJpjGH//ymUAHjHA7OttVkDfzT5MDmdxSZFVO1hOqBpc6sNGxQxXvKzfd4vtl4MBfwBZ
KLk25smFw9SmusqyGqe0E9GsaiFmo0rXmiYJAtbG5waMJQJ6piEu2ADkTDCPIssxRs0LkitYOv99
2q0NXm+A2GrC02NLV+o0qibgmXr657KCWQuQAuR1C7t6wH0Ca5u++VatTRJl4cVbPMEngxZsg4D9
LwcEQ9dC0MOZCsLhoIgkgTMUqprDPcanW0Lru2dTL1ClEzvyIrMs8HTf19MbuEPWnIhe180aDsBY
KDunpR/RALsQJa4Zj7zEUlwkL0CDMPzcV6ggX6KvlFLfh3CTfmHNqx+xRH8U3TZk8gGQuD03mYB5
XCxuD5AMA2Iut3P+5Ia7IZ2yFx0BNC1mZPnnPK95ZGqo4DU+S8ht4eZyQGYXA0S4CaNlGCbJGu5m
ITksjZ1wnv/ExZp+T4Gth7ddL81tvLvdrSTUt9fctl5/kKt7HdTOVcreasw76KallBTE0tfR2Yfs
I6fZkQgn2wPtiZHafM6aosYgQBTUD4KveG8oCMjWWC85VZFBvnidFPJaCX1T/Aug4im0GJO+xtQL
OQPEu/Eu8nkFX1hTuwZiV6Bg7evWkBA7XbMkJc3wcVojJYD5i/CBCLK3TgazJ8jeq8Fqi/zKPxpH
KeueF/UOb5ag8ETzd7jKRwc5Sgi6kJLWMUfsBzTof/Q89YzudkibACaWSLDs17W7DthrCE0IQ/K+
zmRklprTAx5LN58ORfEzd2QeC80ipQw+aV1r+uLXGZQ3nT6i22A/B1INor70NXZlAo1d6f3MEQB7
to/APXbFh3TXOEUTDeggBz5p5n2Hexm0qSdPXR/+qznCGdNG64JwLIsqb3IbwtjJ9ux6uIaAMxbv
WymowFR2JYWk/O3PLAcz6BFpWnPQiOtov/AhFIo8lIH9D1MRhLoR5X/Nu7AZBfXhM3A8u3xJHt/z
dn5ZMqCK+Ok9BKgPrC2cIBL1QyAZt+uNqyaAJtwsr+BgSrXK/sOq184TsqC3zePc/T/17wzQMY5/
+DMJgDaNwlamKBGBIXMKNgMquih+0LemVGGeqgVNpRI2/gMzFIAcY5AMjzcqiMrPdIgfkpYxSPMN
JoRaRNW3y/WD6qOtyc3ym25RSF8hAcRGvN0TP1xXB5+TtbfeVnvAySeB/qSIqx/3csxJy1eXI3c5
gtokgbY1Ukwv6GAQrPQCZkRMY9T9QqV2a9JUKzMVyAEKXIKEB3aWIFDrlUkstqDaGcx0xDzXl/Vj
ouMrfyNU7u31RNwSUACUM0S2Q+RoGFI1BuMN4MOiMmp9V8fPJz0swFf2i16Fq1CbxjuVsTJ/yLX5
+j3n7IEAOMxxfwU4P8YgsnMBHVPPrbEtoS3fzSfFiHpMlWaL5O4tAXWQEbbNZ0FDqc3+su7sDnD/
xIu0rSEFiyo8F+25J/yo4XJ8Ejt4Iv8C9rryNsyePyqPsu1utwlsWXWmSk7ni+3pIIvzvE1rQeKV
vg/X4IeAP+5YAsmZtXKtcZDaNQmZNsDMVaEgMmZInKZH/cWkLuhIrH0Jhgy178pqB5x1B1a3isQf
j8Jzje/g1F97YaNr4jR1eZ2xsK1wCDi1n5Kvw9Yl4GRCCAnQfG6m3Wb2UQqg237AGSWQTe4yCmIJ
sr9v73o5UPCD5a/1ogkhBGOVqlCeZg8DeqLsb88VOZFgRoK42nzKuaEPXyj417LWnS9qvxHMhhiM
DfE0Jl5ZqZ/XtXwfKNM2lDr8Jn3QHLnL8XWPtL2b0Lj4Jr6FmHlTMNFBFuYPtbNe1/6SzFFPiQTQ
yaSw3gdtk4CnA9uxETfFmBHg8zpqVqDJ3ZBwBLhS3f3Pk5LHvW5pVRoF1cUyJpuEVNB/NW2ZHGc6
KN61sCXET6L0dptL9iaonZ04+vmULBdHMdedSYiS0k3HenbW/UuKolh/npOHlktngjPTW1K0hC5y
zNX3r73f/BXJ2/+2GLFflKYjSA+du9TqGbMgPVwo09mLRjdhcv1lmF5wntDMyni0ESsu4mGDfltD
UYlMoS18Eo+l4mrMss0Va7zNlR7hqp81+pH4TE33MjJhov51FbeF6/yqfLy9mmdqX1SoRO+EcC6G
cGccAGLKdD9gc6EhO/Ku3kC/xur41PFBzZTjPI8CG9aQgTtXLc2QeLCiOYSQXb9J83F4y4q7yakS
OEzCjfN0fy7/wbhxYC6rJYwjrawkt1A6LfCQcTS6aJpU70MKplhJ0533Ixv3lccAqaJdsB3y538o
UY7XWrQYyu+9vFCwNnL/bi2Hh8G5NrPQXgPNTYU5tOzkmQmPUrJip6DG5lvIz+fGxkRsD23PXTRy
rAchmH7yIGntasUqvF35rJ3MnciK3sd6aOO/D43QRL6Fv2zBvN1TlmAEHz8Ex/dtlkyzaTJPHwak
Pseb3sN6ALVh0aoGLOzKVnyrMrTZFxJpFa0RbXcV8B9lbfkhOukbg6pxXyNNAdcnpD1DYTRZUXPs
lOxBWj6iIDhaEamW+eANlOguZE+vPC+tQ7LN3/a/Ahr+yJlJ0qslXhg0CVlfDXsQ/2z9kk6uoxNU
WaLBkXgNf+pvIWOwQiUaz8hTk8Mp7X56ogs13cHUF/CgMabMwXDmXff9j9N9P11SP7J3IRbObU2x
jCs40hki3gHAElVfLLxr6+L/6T4/ErbdGR4KX0WP0wN1lihyfT0P6wIE/qOYiAC2YE9+w7LEA4Vq
nuFqpHOJXv+u0p4qQpn0BlsKR9TXE0nMS03So7nz+/7prMQE1KYr76VE4ld2iHh236WFWsq58ks3
nOxQgNZz9idTreC80QiJsPxMbyKIM4H8sQvK+gc2MwMeSon73eztwPHM5qTGIA55wmdyqMDeBqkw
8cN1g+T7h21buZyQSO1vtUxFccqGvZCPWorN+vxVdrmLK44MT8ZCxHzXnA/m634f7TJiwGesFUDS
GSAYLGDtb8zDbsuI0TXaEvyPzqQtJO8+H7pvuZU+PiowQ/5Nln8RW8afqxx+yTKNPCqvWJgkqScH
uscXMpAmsZ2RNDjj4Aj/1Vkzed6xCa3HNwatV7PutFD93lkx7Iu2r/RcmQOcQTeibcz+ERqrPnPE
h/Nj8Lh6N6STsFdY6YSjwVgiEiST/eWZ8y2seZ9lUQ8/kOt5p0HlJuA34355R5JDEVRNjTpqIlSP
gqJOg347hxzZzlgJNTUwDqssgje7qQCjw5wRTUv1xMfdpefH04PurXKZ7jghby03AB8FM8Spg0w9
xhZ8Tq/Z0Vp4TBQMBrlvrvGIWQ4rcGr/ajRvmXv71dcmWT4doogEIA2MMnRHmbGkothmuzZDBZZn
uF30gfA7iAX6z1OUT97bE65yqRCYul/Ykzx7PD7D351fyc+r/s6dG/pwIAezM5A1/OXVI2FYvYCg
iCwYxOuFsmFjZs5FEBPvLNVHoB99FuK5KsB3yp2u43fMThHaN5/MLzGJ/IICGi/6kvpdvFMSC2md
Iio7sw6QmUUrXT3JfiuCXE9SjXy26s9VUtcUmWfO5ZniYULSOdyz4B10gPOuFZVu5cNDbTaMxHrw
sfpxuhyHnxp8AqQ068LrhU4ciJuqes+ion0QmqNtEx5yRGPY4wvecmAY8r+Gsw9GIAa5caQENv/0
x8+klu4s/W5kTVkpJtNkeuUkc/IS7N3OPgCHLgV+he2Z6NRKHvA/VolKVCvOLHPkQm/7st6245CQ
CPbp4veFchPbx+1bNUhX3xYjV2ToBH7FhIy7x0xXgSzuacT3T5yQZSuvBjA1geDOyCU/bt1OKre2
wnvuzg7Bg44AlKVLARX9NdgHuucgeeMpriUsj/EB8Pl8CWZ52XIEABPYJisZo58zYmXHHhrU9jId
7M1XPfSWgQnGuQcnndOnBzy61J+g57DynpOjVIaO+4BDeAm5ZmpIHsqViztarK2msweY6DyXzQsS
KqNGRnYNnY2RB2Sw6ebHxjCggICQF1SPDmIww28hYQ67hMedg9GrHt6q7s4em8lBIyRyeJjwQba+
tj9ZFr+/40DlXU/HWB8wWVPDDbw3PdKEeIf+E8PYw1T332SDENGhgJLv0DFIIl7TOwAYvSY7ulr0
z33o968Ly7F5TM0VSpAKSSPwCXYPbDl/JHem8uvEx1Tzw9fr8GDURj18vmQURh5jox63V/BUmg3k
VEdLx4shJZKpoYP4oyhGGV6gpIOfw/PjHqTBXagH6xET/FZRJtvb78Gh39fNbz07FlBJqHkehCfy
7aIC45JazO5QmcYv2e54ZckYjngAFm5O+bgkAZN94+ytZGroU+kGkUNlgxc5QGZ8KST/elsG/SyH
l4X4z2kQU1ESilk0Jluef727fxMHjZNRIJpRFORBG0GkhnDfSAfz63UW2Qaou+S1EGEaNfdDErZu
D96RexzBuVixLryZFr24glF3HfF0Brx8hBgmZYq1xjyVz/SiK9Nco5B1fDhjzjYJr88qFojifF3H
cnFjrHfuuYHdhOkMbAbUOZh83WjtFIrrugO97gJYQ+AAnzeXV+T0dXALw6C6khwh7KRcdskJPx/v
IA67ZSC84uuO+tKhV0Oi2QcLw05d7BBOKh9ps49uLrftkn0O+GrSxvHXejOXqmS60IJlvdWeORwr
Xcz3cXp0OY2hmcDqwp0LvReIQihIwK+/4QD6caxmzEB1qAfyK4RKHPOYl1zwz60HKFfBh6xFLq2S
FHl4MQdQJlDaWGd7DsHlPD1FRgdEu2Im7vt+JkbIXP/D3AcKmyqPSV6s6Unz8kBNbZVaMvZkM+nW
eRnLqzTrh+StB4QZ7/FYtvL9hrLWpZhVTxs0TQUwmQIWvCf6hLtqJL+NTcr4knxZ9YfORAirC3f7
H6VUEn98FdSEwEQmClMTOB5RNFxBQ/+xDCj+sN37iTsyVkYvrN7ILS4ibdMh7OSps5afIeVPSUAn
JdypJ1iUmbdqPvTHWiKNrQtOyw2ijP907vqP5FrAwvI3js/408Vh4eV7O9luMYuPPER4vPicI396
dzL5FcjexLUXIjL8DyISeeZZNUG82SgZXQPTcimkGANNS0K3d26uRJtGgMFG3X+TxqTJtCZ8MAnv
bC1QvCn+A4e+rF3FOv+fiJDzSqYUC9boEmQFBwOSBrtrPXbczf9DgWk90zW1vhzYfF/uJ51GTPHe
rQ9qFex5dkzHxe+ZXMmmUPm27PX9Wb+//c92HlDmgPwDzSj2RVhSkFIYsiX8A8HOyW59Zw8q7Qd6
aAYpuyCXTbr8h3jyVTZYgWduORBq69Ooi52x2KO6Ty99gctMJ/ofOz8vO7lR6of3uXg3+RYolpui
vamwc/h8lrtSDkUJ9+wwPJp7Mexyh3gOTrLeq+bst7wAKJVl9UmW1ZUZLb+nyjqXjT4DhJdOhb91
OeQpPDFSJ3IUYfghygKm0O93JSviBCPjh5lmvViQahNZr7JTCw2u3xidt6rebSf3VUFbGt5hwN4Q
nONJo+irwG88p1GPNudFYWZcmI7bOs9OCWE5gC/ldf3r08R+b9IWs7IZAwcuCSAas0EQ2AV2njaW
FBnZUl1m+zvatr/3u8q/e5kVcKXhlWsPZlZ93hKKmMHWg5aSjlOh+d8nID78NvzqVzxTns1pwyTg
CPGtL7q71j1GTLoELa4QHe+Bo02ftFXipoBTXeIeKr0VcWekrI2x5XScOtSqANhoMgXegwp739ON
Wk9MZNE+nzxKNNAtwSozuEnxHtZhf/iN7JCjgtZnS82AXIq0+v+ywQpyuaImhndhkOUJrSyu+xDs
Z0aew3lFtnnufDaFRN5TSsocAoiGADCESeSjA//W0IHKTNBz2iIilzHtQZLAL/s1nKFZ5n4llG2s
8vCqz2v/x81uv8oEm0MlKGSXsXtvtm4rpRbkenr/ceQe8MXiqx2Nad7seTj12tc8Z69oJlYkAmjX
nzgn6AN2H8ZYe8hEFBpAJ/2Xa6qM7mXHaiQRXgEGdSUZIZIJSs6eo38LcsqRVVx5UVyS5hg5+P3X
jd6nOIR02M8SI5f4z73ASIuzFjC7xMehkQHBAa/9bu2t3l9I9GX0KHZRSUMm4+4T3vtsE2KP90ml
bJQf/4oHgjtqzehQN9CVjT/W9NBALnOprh8Gm9493NMRRkbE0Z9SKjhzp+bFaKXiABIbVVmbzxXj
TP8Xo7Pbi8ZZxzRz5isiXQ/d/0y0K5bwyxL3fHSOWL6zvcQhpFP9YLrFSKVqMk1ygs3Cil9S8OuK
KLxLGJz1jNWMfK8ayPuPGIvnWQ624ujT3t5+gPum+vVvuAKqevCKu+io7x+c+XDbRjHcX4po0iKE
bm+kzqiLa8jK0OvIS/phyyntzzKaAnt2aRzkxmqqo/Wz9Q2AA0xJQRPoLOeLO4704AHI+C34x9mJ
t96efqZZwQGiQrd6eOHXSwUYpSIMr9Y7HgEIFQikIiFHRej5+nhsQxqM6laALahQScVoxzWtkgV3
wRt0MfqnmGGTZaNjovV2vYswReEZOl2av/vWp10pXWfvW5MynveniAebuEVufHR579cndH0nX6Zp
f4ZLGqBhl3vFvGt28LMpD6ZrQMcxk7XIfZGVOoq/wMgLhlWgbL5UlJxG4wVKXtpggEV813+9/npU
HL9DIOgCWWibWJV906b3HzqiIBVSMF9jucgt+t5tj/VwUfkQQTxD6DqnaO1t1tk2SfMmY125d/se
9q2lBxoUK1jx3HLnD6Q9VSUAIv9EUHKLCKNDktoIqXf25B4fn3tXm0lmpXTwuNu/WOfyPMTXzSS0
4FEI9fequ07LyY7nMOWN0bLju50oKVvsmuTFZkTCUB1joJo2aqZhNGC2oHJLgR8yNQZfn6/fjTzH
qaIwbMfcPMXavN39DLVLrMih0Qkoiqr8PZIXY3OkqIRdtpFIlwVxhzq3aYlw68mv+7gaNzgmX43f
YObbhAkhp5oFq+0unhkP367LmzHmF5e0caUZQMa5o467kM72zLMSEFzeI5KmLVoXdfIurwtE6m91
SbRbPvwDiYMnUn/Ds181PZjbb4BFRJUzPjiKagy4IEenyxgD0FzXDnI5iBHxT/NV38OuXPoeChVG
URe68AmxWqTgNWuRvX7hjxvX7jJJB9muiA8qQrMn1vw7l+fxBOCfbIbDYSGh+6YPgvBHVmkO1r1D
LQjCQsLmo9pCQw4ZOhGQEnKfaezWPrnzibkTgd+uulRf4QuJAYfeLfj9GaJglt4jS8lo3RC4JMGO
K4O4uGTXcRVfKYs9np8Xw/avYU41qVhqDKX1g1pBGcFga41cSkrXSaDvSnYqY7y1UsBCgu+d3Bg0
MPv0TKdOVdj5vg0NKGT736VpZEK4vlPDoJwLXeUe8YipmdIoeqJCosrc/XXqTLsEsqb7zRbsczY2
7J5ZGT/+G79tFF9DuysUHObbpNgMWrniU6Sw1tYEtW9exTP6BbohIs2Ky5FSugAmDvSH9L45yEEi
70e76vPOuUheyVcI5pSr9x28jUXoYiz3xebdpMOCqlWUbzYOY7MZqGwUAvMIrVLw2GDdPLYv01i4
oEYv0xdDhC7qE0f0TQ5BuZbV7pYgzjkf3sNy5TAE23cRN+A+2zGuauxu8Ox6njDxzdp2uwF+l7UN
uFMH+kTqX/X4JWf4H+7w9IRJVpT/KUUivt7zB+2g96xKoVzbaXQmRxv6YCDuAeT6SXi7ZP7zfBwX
FYib3SJxBk+HZJtB/E/QDxCYXemXSHTsi+TXm0ynaJetKb2M50amhNcbdOm3iPTZgbbTk/sXl4QW
FRDu/bNfB+le8+A/1SZumCbBEfIh1+FhoODTxSVwj3cI1yPyfM+Cv1kpb9ShfaC42VR+qSr83uFx
Y7xQ6HbYAkzRt6Tj4hLP4fcJc3FWi6fTWXc91vOY0yI70ckYfx08sz+nIf6JVTFfN+YNFWLyhO/z
/ZvWhbyYsHYVoBEpX9DLsXJvjVX9TDq6rLbU87824LlwzKm5IqrephPSqIuFLk0LCovVIFc9KfLT
O3mJBnU6t9NZ/YktTUg3rPLxLUgvixCptbDLBVz94wBWouwoI2ixN7yEWcpPsYmFA/YeLRM3lw9X
mQ9oFJ1ruDxnfsI2mO5FsXCkIkME48k2HoZbapVqGhU9BashomUg4GS31CoIDTEY4ofDd+t/nq+B
mwT6+tcnqACWGlXP7Awb7zi15YUad66GXtiRhijP0R68a9P75ycuvRsYhsa1/KUFKNvsFGiaXtOB
iKLc2EMEFMc3Y4M6xm9lQ/UzHpTfg+rLLpol7Z0VdfyViE8H4Z9YHcMeX4NSDHsEP6zwiQgMSb9U
N16UgNwLt02BeNPNlEnRHEBeUow/q63QQJftcWbJcooM+63jxOZVEj4ehFZ7qR9/9rcEqRdGISF+
a+TIDiV/S+n2dFMMGwTdWZ4Rcfuq+dKcEDKXXO6nKphM8Lspc+dLYWuWmiQIzz8C54IlGnq5Qjn8
/09mZ6+REidfyqrfr5vSSIxx3PObJ9uytEDl6yCzisx6ppEK54RI+Qux9PstgrRAMrmrJL/wdvVh
mjWpivIogaP3KrtS/BxeJ2vW+ShAOBeV0nqL0Q8U/P7t6WKP5GTYcTyF8nYE+0307J4ctDcJxEyU
YiwtIU+X3xB9mW2Ks8d9J2xUG7NQgLSc+1mdr0eetOCQGirqpwmxye9e5LmkHen+bKhpO8eKQRaY
p5DHvvlXl1R4bOPglwHrNM4vlDoQBh3Nc5wrV+skrWn5aC1+zYg9Elmg+hf4sAoTI0aXcwSf1b6M
cShdb5egOoujpynIWYEAitdlG6bocu3kJnsJywQaQLtf7OF94mdlechfJPwXDs7rOzBgjaBF3Qqi
kTZMGFU1yCkVe8vSX4U6PMBpypfGw6zUrZbzzXdj9qzeoVM8r6QS6qQCaHluMiNFFMhOm5G+cHht
QxhFYiIiir9gZT9aqt7Tcq0O9no011tMwdz2lA9zNYi9Gtbu6irc0bLug0iQPFRmxY+jBJNFbwGU
9F+fnFeHO+sga+jBH//0H3GSUZtekg4WN77xf9Ks3vIIfaF2n6l/9jvpMQsHgzVsIXbeqATf9zdt
SH2+0W3vL9d8BeZxZwGz9hPwUMnw/FMvkM0hE9g4W6793Z/3JJ+MLfcEwdmZDis6L6uY2Ti2EteZ
CaTVyRH68bilSSS4mwg3SMYHfBLb3369C4hhAhO91IbPdsu3EkHwRkGKzro4xg+mo5GCq7zHH2UF
YIHjbkSJrrGHsPV5DUpZogAArVNM1/7jmkW7VeqFIA1iryg85nGnSZOVqUmFDjBAKEHqgct9R+dU
CwghsTBZXYSJ727Ncu+r7uVjInLqODBduq/Ktwgk1rGVkbQ5EBcK5HhxdBy6MuTgl8R8lx02p8vE
2SWpOHKSaWQSUVEBU/4JBcunRKcssNAC5kcqoo7VP4DnTqImyA3LpnoOZoNcXFUP13Rba+OSKTGY
uKOMss1zqMSNdd6OzUkBMvZ2apDAb1pyFM2aQkoWk+/hTT+XQ6Nf0SwG/FJl+KdchOPVElsdEMaL
wwvr240c5o5f9SeqwT83UMnjYMRGCxw9zzwvWP7EiziKd1GDIS7ajCV8w5kqiSSSnmA27FPuBYuo
9Iuh/LrA2JNrOymGyKaoe8XZybf2BWjEZLRb5eeZOIyiK8cHPoYJOUjLb4PErs4ceQtbWd5zo4N8
JeoDZtRtpOWcz0omTh1dwMSLTPoYWi/y9gNHZFxfg910L9iHoqHrh+yTTLjO0s0LUsBhuU/qjILT
c+CTfUVoX0dleo1F7uhuK7ZvnUgeBErJqCx6W6qTYFf9Xeyv2pBFoXDjJNqtKA5I65abkrA0Fmze
HqDnjTNvF1eu7n2qmcfxHnRbOY18T7/7M7M3F05w+YB4oHvYZcyXB+8BLXlTamQdHFUk4a1UAPwE
GmxiGfITVQi8cOA686AasXk+QhgpYYRzBJ3r2jaGSc4UG/yKF33LawBnwcLRW1gEPPv20N7K+SSP
5H10goHqRsrwUY6MzYSKxB2oxPC4ZWfhfy2sbho1APXdFjYStppSiWOmhWJZpVCaiW43oeB1xIr6
8v+cglsCKD9a3xVgSrlGlpHw5VccxrYvN/+/hVP1VgtmTgftTMmkf22PDILbBy83LtVJmcHO9FpY
Hza4SKLHMsLvFAjnZpXNUP/GV3GHKwxMVt7Ck28QPMkwFV4wpbjSUlcsoT7wp/d3p0m06FXnjySK
6UgE8K5XXXdGPRzRcBJZ3Rh4XptMLiMlYPi2RiQEZyFw60m8IqU67yvcmm9+lRxK0yi8WYp2MmSM
yj/xKNo5U4Hi52v01029qrJF7kWBJhkb53ADXlhnNqC0PX6CwXsZngWpDzeYma1pId4f+bi4jzkp
jThHHAbbXLZ03bTAnpTZGWbUIiKKiI18IbslZUxGxFdbRGpflPI+1Yb/J8CrYJKHztSPRIaz9CYY
7ujsQo0RZFxhsw2udjm+NP+KUEsTVH6CEV0YT//fZOt7ZZk2AWB40WzWB5GdH6LVgbKBuZem6eoI
UesRhe9wZ/4IpO23IriNmmG5xNJ1VvU5W8MfUyEQNWVkVrdWs81nvQ6Tk366oIP/SkkRYz/Y/4lB
gZS2uZDCoqzFJdf3etrmKeAd7HhRlq/5LXRxyluorUby19/5Y9avc7gZMX+AU0HIOZ8+5c+3Q0OH
FWExol5+XBgwou5ZKOFeAns5Kt3rF1aw36l50SxE725FrmCsHblJnRhKHyIkCahbA/kU3t6eCu4h
CT/h78qnb8UkFcvUmjrsXh3YEFcivoJxBciZiGCBLa16+K5g1nfTfP2nEiB+PJxn2KOD/uq4KH7a
MJy/EBEsc36k6fU5NDfxatnzZ/NYM5H0ucj474ksKK91MZczgAnojvro45hgvYtK2LtdbGaJCzZE
5hm9qfb2N/XxS7Lm1wklmj661qlsnycXsBNtjgA50JuWSR8QZyO8NHyPb4XlzSFoe9P5UGKMe4Ro
NIpZyXISyTa8M9RrK07kmyWYhRAOO5HRw1wWE8VvlCy3kOt4FOPlFh9VXYGnwUL4qWKP1d6EDSCL
64703doPLotlcp2ODhtLX9hWkwdmJYFD/Gy9KKJe0/RV/A7GaNZlVqq8JzntvKyi1/uJceHVjgvB
0KZr8fDOVbvHErjsXEMVBegeInqXJQAMM7U0yrUF5sY93xifsRA2ZKCEIduYjyyZIpzSN+6qHxGY
xLb0E4szrLAtezdOa8fVwZd2tLrAUFYowVkG01wlMGL2ImYPkNCg7kF74phq22pCaUqhzhF45hwR
+t0sqML6rrkXaEDz+yCWHx/pLDQPTLtwrz4G4I+4qcKhzIWiV06rD/yZFi8MfcR6GCHnj7nfKCN5
d9q9/8oppiiKJqxm04UR04y4G4aTrvd9OVz1Ift8AA5/koIvgY4v8UsLVDVBlpWl01T9fdORADaP
8557qokM5V+5xLzoe30y9IIKPFZxUQ3lLNziGuP40/ykB30W/TyCZ5ND3+csLmjr0U2hF2Z/CeIy
KGWsaSM9gVFATFCyPdJMdqDmir4So6KJFkooKlgMYomCTzVymhuvR3YDVCCgZ7H1v3Nxfl5thTwh
01Hxl12eMx+c6OMXTKKnIL+wPU5LQxFIGWLulFCTCjsr9Uwxqvh30sB+en/UJk1HMvwYslmUMToR
N5d1TDMf0UAuV/GiCppgiM2Ltnx6oZSChbU0acxIL2sbq/3KAbBefyyjM8R6NMSZLNd2esX4QRZK
j7pOPGcx3524j7LEMAIILEjL0JCqUPHlSAIrda1jCpcp5qBYfC6OLdpNerTFHMO68bAImTsiAMWh
vvlJExAyvAehkfQXiUKdlmbTjJn85gJHzQM/L58IvzDusyG6029inx18ee7v6K1ClSCQIDMQYux5
iC7SSLs0LLXbAPmO4ZyzmDRZ3MXT3AlqXgFljpFvUIHlKE0tijrGCy+oYg8Xzv9YTp4SLaG9Eq8P
+8DCdxR20PSyNNoYAaWlGA0TsbfZEePwrPwlw8CAE0GCGSJLxs8odWFpSNO5HoGZBAbBwClOIE3A
jqOWrpQsP2WfCAeSdNRwoL3hM3uQpFAav3gnTROeYD07nGd21D2eX0SIRst0vRoSmbUQHHn+f2Tb
VACRQxUiD7V8LyisWO9Bj9zhiKWS+faCm+RS7X0z4pRJSQMrQw0FSzXeHThsBW8Cllol3yImRoSt
e6sYSFe1YgGkFRm4fxtYoivgcy7E8IGXKqihi32XIVYotiTl4Cl+GvMCPJPS34MoYA43EV53qYzt
81FGXAqQiYnn3SsneX1xNesKu0La6ZKSsh+XsFvDZGYrEUe0DwszG8L65CAV5uMU6gLpapfjeBUe
/63LZGelSrmuyMpa61gqp30JMFhzLTZb2ic84pY7C27YvzfxIfGDrKWmGebgm7jpyf/FwoW2s9qn
s+hyDC6Hw4Js5F759nd72AySHjcjtKTHjfYVXS8wXbsg+Enf0Au8iJphZTAiq7nhflJnbKgUZCdU
Fxm2+boi74wXnvahUipemYX9iYSJEzvpysY8Xf+K7B7ERC5jVGdADmGHjSIw3ERPnynvCFYCdD86
wl+nEF4adDXLhI0lVgicht0clSUki9wyMbvwaO3du9OuQOMFX5blP8IHKcenunpguZG2Rc020JZ7
XNQY8TMga6TODYt4YVprMV4iQ/DUceUFcGWfOrzw4eKqtrHMoBiYer9Z5xVZ/zHfOXIQAcWtM5re
c01k1rz46C7uyw38mUMGKA0pVjpf+T/LtFKXO1yXjemZjFjjx/dqL7u72hNqqiOZl+7O297XgbEm
8UZt1w1Am8nHwx6tI9VJym8bdNI5Ev6qyotaklJNMSN69E8W15bvCVZiJ6hVXIW3pRbAtmjezaKl
+oQp6I+nyXjaUNnL5Kiiog7Dv7z/74NrRyDxQutYmCXFuJB08fSyeDW5Dd94iubAXTJW00NkAMWB
DFeqNdgTbgO17UF/cozWoCGaPvvrREiTbVcYPWg+KymP6KkrXoQ7wqbcj4/+JuARJ3ay/6K+mn25
h/1dfWV1fKguB20P/SQM1ke71dUh3x/6KChyVTi+qHfzlDu5k/W8x0w/WSaCNQEwOmOkO+rk8la9
iVPwJcAG8eGOduPQGJFP8Ba+18inBccPJk9Z4cklm1hkjB8O3Brx27eUpQke5vEuJWcvUOzJ9uAf
tBVmCpkGlTX/ysOA622hXZo6AAoSQEuiioJ1Gku0/oghJ6h82IzkcUgA0ctgbHJjvPQJ1uzCmKpf
LuycxFz702jHTpZQTrmpAoXvBJBzHYo/O8PJnFNIinwMornNIFJ7cJgwpxYf/p5MqkXjNOUjV5Db
tSq/icgAve94uxD09tJUPecsWYmaKwZ2+B+GTKnA0eF5h4SuovxOCRSIVjAjMIGJZ2vchwQGvUdV
JsAn8lvAK2w0B2aOPg8kUvJPd8ZOZ2Bje0gUxdhDX1nUr3JH6MokQTgQY/CrsGZYoq1XXlS8hQ4V
YnKPzBa+nwRdsfyzko3ke/vm/PLcRQXkGOZMWXQrwfFAvi1YfkJ+alXg7gj5VeChryCwcTjYHgbi
J72NF50UG+rGhRnyI7IwMkD9Hix1Qy8xwtkCeKGnooHIpncp6etyQ2C40pk7k4MO1dMoHTyM08Em
2JzNFJqFqiSs/AWQhsqsu3328pNxrrMyLpQkdyM94GkNWQH6Uj/L1Kw8gaqkgvoK0PSpMgdCbwIf
ZksDg9+EjOLRzbqtfFmbkRVWijzUcln5mAG8v2JH4Y7S8TDNY2vejZhIZaA1/MKuvKHxZvwlEQD7
iotMP/cdefpoEvOQn8Oh5TdSMQ/AHCfN7Lh5D8NDH3Db8fK63luClVl7lEz2S/3SHW87J1Dg3TZS
qw2zQUMbHptRvddDmYPMT0sqWYhxcf/QfJgbvuiplQXeG8C7r6yim6oTy/S69KPCm8NF6UwYmg1R
kVHKtWtLV0iDbBB7b0yqQhlbiG9ZtdGJ2CdidN68WQWyg04LEbC4kOWzlL6q1zCMj7oxLfPbWa4p
uHG34SI1C8Z0DEOQMsdEFlnYWFPO7lNdN6Hne18XRgCZGmiJ0ymj4bu+kzaFKDb7n6A+4jae96jL
qicoLQuiHRHx2g4TNts1pFqBrxg/zPZIhhrDo4QROeGyMvliDd1L3BUlHhEgC7Rdd32la9h0oO4q
TvxvJ2/UcfNUT/OSeNMJXASGjt21YVvmqOUFxpg5b8vpffAxaRgUngBvDvLFI1KjhQ8qhAXge5fD
nyvYd7+IBaCLYK1SwmSisbi/7xbefstzBl3XUrbwcs5Ig8L7usSacXeR2YL/RXdKh9XqyfUjgC1h
HE+Bk+8ozDC+/B1wyRZVD9l/khqjLWRpweGT2wJXb/dbO2Um3nTHuuyLcqbBKROIUbyYdm4d5eGM
Wfdb9K3Ju970lQsOjCJAK66Z7+a6pNp3aY2IjJ++rs5w10wVY5ejqa2DuuCO2IWjrZazxj5fTU1S
qZXysU+pzATWFVRyzvmo7ybuRp81cZHHsqz5yIl9axL1uE8KAC2TIqnA0z70hf+Eask/NmBR44Ti
9FD9g8wxCa3rD6m9/kC7XhPfv/4hSHpIZklQ6ntpAcXZZ1AQL+/AkxyMDp3mloOiqgK6mFqwMNyV
yL2fPpLOPvtUHMGx5gw1DXOAU9oMPJoAcX6f3PIDIL7ZZmM0uyDEVix3iEDU/rzVma9874i6uWhh
ggoJSekFDgATz3RDuZ57VBXBrtpSQrh+MIuiLEzt9qjRKDC6GPpMO43e+HsKDBu4gAt/kp1L930D
oH7iPio4WdcXmFXOmerWIgNLr1pFXVwqqZpOfo7GNEKB6N6H8gvw6AmahmiOrsiy4ULFDTNPo9c1
O1DH5K3WG2P/1X6z6b2BqxmAZOtf/PdS5nsjWCFCrdAXId6NeG7fhZZ1Pz6G8py8uo1dGqrfedFv
jVwME/qjGg047TZ7xx8hVRIXDvIwDQHXW8doBt1VEPvhXGhDHThpOWtIZcr87IHWal88grl058mN
L31PKtGLHQ1XifFjLJp03eaQrm2HdsPxpOaLH2mfSw6F8i11NMgs9wmQk0U0h9gP9qjL8W/NlMZK
Y/1BDMJG2m0AFxHmTNCUVvWr5O2cZD3BFxvEJXI+z6kHQ67ch8uvaX5xgfCynk1M7rxBF9ED5RHv
oM+lyfY5H+rXDUftZvz6Kb5bV5Z7++3gZETyPSeu0btgHtZv6y63xf+EMN9APNHrAvaGVRUFIgOj
rmd/053NrP0MkBRpQCUoybdttlo2pxRhGXgFcvKu8QOsQNa1LYFAghqjmDIpUJS9qtGo25xMbhV5
pssBFx4wybLhKbiQFGYYCEiTsD2updWJuHju4IbaOBXvg2NPv7p49zq+2PnxE8JngHJyM5BqLfCg
8xc8b87Gpx195JgNIUCWPyNextHRMp6xBnFprwdwYgtHztLcg/rt3zdTqM+SP0j6Ub9PyYsTY9OJ
XmrpGlyqUfEmVIoHY4RQiCsvR5qREiSniK2N2CqggsjahNrNs+DQ7qiecJvK9GglyOOdA6DgULdp
eI4RbE6XBxP7RC4mmxhlHrNxVrrp62360dgc7D7KwE0sjCF3BW5SM2/TIfNsUoduxtwFVgHW3AsS
5FjVK+PK41SH3GiO452kF4kVYaqmTo5fspl6v76Zgxy8aSBbkWcXD6hnU46rk8ARPy02uYUrmha/
Hffu/UskX/SGIQ1pS/lfNk0DGtheLZQ+wH9EblZGWZ4UYNJVEjsg95Uo6s7eGG8fF0dpX/OA2HrI
Nob4qsBT2cD+ebiTIaSSwSgWT4fnnAtVHfpSQEzAYHjxU7Q3RcrSK2Wwffap4Z7zV/l/E7HIIigB
baX4/TRmyTiMTgiYmsM+bjGk/jwgjJrc/urbzPCGm3/XB8LOG743Yf6+/0kDA+vjJDrOlwLoLoir
n9yJh5ZcfpaqYqV1VLBccsJuG5a2jvm7vmY07hrVFSCcd+mH23JVszzi4sxLMKiQjxADlR+YllIg
ouBb2gGPEHDW70wzzz+r+w1Cdzg2osphhfO+OB4eD5npCwSNPX873iD0oOYQzoN5TA4BEADB1UGU
Us3HlF3EtRtL236WVJP9O/ROmv8usJTg2uJ8tfaSyTdOOokVk394aHZazuW0mTkAk1gdBwSAE7Zg
nR1+MrQjp+00R59hCDIlgg8HuaHp3y5PN9hNTnZKb6xsFD6k7lqiaU7Q76Pfk1D8Q/NO6psXVuQZ
qNvOv21ZXwn3wkfiaaNA/zpKvvj6VlbecdTcshs075ubuFbWuT1zN6ExzG3FsquJfUEZ0gQq34D7
oP8oHThd1FIE6fWM7qctppBKeRAyp9n5pLDj0QyOv0SBPkt3DzLR6dXsMItZ569Vj6TMeJQ9y6xe
7oFeB+fXoWxHwFzWAeNF7sMj0D7EXqzr0rh7KW9GJw/I8yGPm37nce2Hn3t3S/fbee5kkIxE/9iP
dNBkN62o2PovG7MR9sJIxE7s+73smA1rdNUTAg7XZCIGzAHlOqVOyVRdf9PhdAVziTXPERUjockS
vt+QSokanIdlCio/MhDttxUjOldRRK706Yj2GtEkIOHWYGYbDH2s+kaWQiBbxeXnde0t2SNE5nD8
XkbFwrEX/SPF8t2ncO8ZxQ4yQWH1y5Q+es/ecJlRXV5DT7BGgSzxc+1ufsfQqvJJaHKFOaqUwSKp
J3TAxlpM+dRp9p5jtIuMb2o9446KQyAptyZpqlnfgNRULpv2GCP2kcWFLF8+DFpxulLJEZbECPUz
8szIlQeNu2sZ7Zv5FZ8f9dK0Rd8Ec42Jd+TB1lVdtZJgsSPLARBPJZ+ukRQFekV11v9wwVUKkDvk
xWDQo4qhRRdGmuzshyy62N2E/B9V23kfUlDL+DlWyW9blOrcSY8YfDKh9+pSn+U6+Zz1ISLBL0mJ
0hw0fYuYvMdAxsWB6QcGpYPJfm9ykiVTewl70GAL+FQQF1+USzBOmajo2QyfTCaFgN+Gua8Tgfpl
xZckOBWAp8D6iv8/KMScHQ1Or9ES7Ayrl0CeUcH4+YOUTUHgA5CUDu9EyzHQJgfpDaPAJCTwooGU
0LWA4xRm4sDoTY1oQm3jqwY3NDce+aUmfs7rAZrOr7xLp9ZZLlYE5stU7dDHIYDdpsOSXpCcGS5N
azwNgj/RgFlApsj3X768fF+oC0QHB8vanuwp4xgw9OKBQRdkGn1anIYE/IRMR24YG7J0hb35ivLO
RDuwNRkIPQVLU4wAOy0D0MADJUri1uHHbIvo/xUhfU8VUqefgq9RFvGWbQSkhIE9Dan40uAC+aK/
gQLtIi96rmMUFQGhbkGwa/aYAvmeKYsLEgHwPshf6h8s2Zn7a44Qzw4s/rCwMmg3iQFVeMxLGyU3
Em4XQwNMxJykG14Z9sxxuA7flb9NDfzCvWuyGwyE0wBI3b0pEJYFKJAj0x1+ncewUtUAmjmUffko
II2GIkbhsEVAdhz7GNELyNXOJv/4NlLRP+A/BoLn3OtRSS40YLIVXHfaho6UtS+xDGs4GY9keZWF
2ZYXRm6pg7Hd9gChMvVTX2r5DN5NHTzosG5EqxtprRgZlYQepq5kdHco+9Ufk9v1k66An/R2dksd
YCA7/pFViXBSwKHhq8TE/r9BRmcMZa/H1EOYi7jR3aqbdhE9VSthZhLC4kd+fDwyX6Kv/acUILyO
m4p++OtD5Fvdzu/CKIwLt1f6QcEQ+dpBBYq1Xod0XtKhoP3gKudVQsF6n4KJaVx4uj4NIeOIidQW
FhWW2WIKrgGtBvAosE/peQaFLzw00wDK9A9bnYB/ofraLXIEfEWgL/SM/pTbsl1P4S2N1zCZSvQO
1iuEx9QL3epcW45Xhrabng8Dh3pPWuj4YdZDKvn9rOjsWz+VElt+NM2Z4+n4/T+TxaIOBLKiFS4n
TiDLsst8pd4SyfzJMtTAqH1heg3fSfUi2/YKNxtaebq9Mx847WIAjCujV/QEVlfQO8YeGNFN8PgP
yql3munRQiiSMKtNpfca0f1Zys7SYV24AdjWP+zvaVbHR3AQ50A+tmJBPTBroAqgO94LLCXcaZHh
i0RXN7Jz37tISlyhqzHBRVddDEE3wStWkzw4X2xAajcSskK101AasId3XhGzhq1SQicbvIPXW0mv
XC6J6iB9c8yLUdFMn4+645D9pkU8JEAWB5Hh6z9WsrgJTiwQ5AABbUANlLhCfebt8TpW1U1XwWz1
1gYqBEfhbS8V/gK0gjFgIf/QDKe4MqxbYWMQ9kzzbh85j8qDK5MwplLmNMby7nSWpiISGghrTcK4
wqV5aC1FZfsQHpqaXsxsV9dGYHGCq7Z6zJFn8uLlamikjn8+oBhvvy2GMNzLDUwSTzJMtXD9pWrv
8kEQhkNOV8Eczup+NtpsO4S1sLyQWie0WiJf4tu71WjeIN/fNvHWs3gJW/B7s2GTdOxbDrw/5Uu4
UBAYWuo+c6RYTKp6vbbOVHGbAYeI+8bYd9/zBIGBdOPvpn9zGrBYDv1OIaWboK2Ez0TkguN3W3df
hzQBF3XiD6RFFfUsamuxK2SP23RT9Cw+K/uzqr0rQp+IacetQ+IEIZ8TJpqq/uKXWPlMYAO8Y35Z
Rq45/bYE/gXreqxEd/2DtLOw7z8plHWQOhLqo9DCAa5UDRXk/iDcbDl0iL/x+LZcf8u9FOfUhA0n
PJZNhQ3pmxi0Wzmd61MNrw+CguFR4dl0leXbNWT0FRDl2TY5xe/L/pR5ztNUwaPiQA48ijahktbh
hQQdHDKcobyjj3YetDx3SvcgWteBlLLzOnhu/1PG6PE9dJcbkt2+3MztQushnilG+qIyeyWywAHq
qtm9Aj5ZoPe9BYk05hJvuxMVM5mK0VvU6sM1K3rx/iHp+JVS7ZGPzy2AS92PQP63DF5J2zulyntu
5txGwYdieU5e0IoerSVoNiNsjiYOuH/NHsu+a4B/TvHBQsKBIMhRTnIYAFPUxlrUFxDTzgfqqT5p
NAni5/sBC9hCJrBx9iTjcVnKVkIts8iNtOwGXpG4mmaaFTCVo2puFgsZtoRgYch00YIaQ/OFwEPH
GuWjgQewhkpASMLoXygNjRbVurmyYD7wFPWcq1ln8D5Dx9DHGo9oywNklko6+gUBP07rlQrE3lab
5iF9u/rVhA0zx9FTKnCifK2MXRtS+y7CwZ6yXn/aC+i+9vWinZlBM16tuPfX6EwAYsfvgiZZM55l
dApgZxqMCJJubT41SLaKLum7wWdqfLCcpGQQ1Da/CrCXZCCh/aCG02MuYGBknGsZNqGmuKz+And8
gEBvwrikRnFOPwaFIhEypDj2R2ilQEq1cz3LuI9k3NovEwFrZ2FuqRgnDUbZTX340SIOhyh9qMWn
Atzz25ibBe/IXjMDFWVNCfj1qR9DoG76azuHP2OCWQG5B6lVQ8xzOUoaY3OFVwteq1/+W5OUf6IA
CDIQ+TX8x1ZSmevgnIQbkxJ5zsqLpI81XeEuTHfQ7K6/LtzcPda37Pwt4CNKIv7ugwYJWu31YSoY
Vn+68WwUoJz1QUbBCTKy5fy11lmVY+Dn5Iulan8624/WrwD5W9MmXnFSCM2khA481pboDzimTcr8
go1fFS4SYkiLc8I+i8sBl1agxhws17tj+MCaloyGkM92QTNIdNfMQOA9rfwn8q9uW5T5XJk5RpXb
1y0E3odHj2NW/w6s5JhExv9bbzF9ZHfC1y/snhawYg981jU+b6s3T0/Z71B3mHb2z1LTU734tZAU
CoXpAlEIBvXiX15yKVhhHvkXEbIvp9eWZa2lG0X/0QIQZAxyyh4bsTuV35l+1mPxGZplV6A+279G
lnVCgbFpisv4N7TEstnfALyXnX6xEWfqil0dXk2zsq7gOEHsfHOp6wAflC0wBDRSFLvwatjugRgq
O0G4sQPzmj2a7+U61YoX2R8g6kXDqoI+iTyCtcKamRCRXCm+679OA8NXKF1/KHSxUovEJWKYV25P
Y8esTgEN0/O81w85pQmsBgc4kb9OUqEa5/9A4hEfOVsJVHRBcef1liBCNjoQ3tBx5wzUOlULv8L6
arJXTBoj/knZG5xI0gEUnAXjsSs0vtwD0SS9D7Hur3Fs4QNIiTPKDnwnMuyDeI6kvCx/+/vyVWKy
wWR6pkmHxTvzpUzj5CPzhKNeoe1DY1Pqj2Ji25o4Cf9D/FHHF5nIkX5HWgarP7f0uBNKZqXvMz1Y
wFatvoyyI1OCIfDjmeTD0MD3sgfG6s+OPsrCDj+t77GLKTUO5ekW1pt+qo+Ni47OdNYenF8cx7KQ
pKWnMg7wCW8XzNs8YTJgtscm/cMJR1YMV+dUOKTXTm6DzVuxqCq7bN0fWIu5QQtUFWAQnFBMFmOA
G0op3t70ao8nuAsMtJaxfL82UDJAiwhsAguLqaWaPgzHiBlAhM8pfdLhDEPa3jm4z+Ye17kSlCi5
zoKZNfS4ElyuIpfbIFH2xUUA8Z2zk1TokMMpdRqjNSAsLiFDMC/JaSQebq1K3WfmxSW4NdfFwhb7
0gYopXHlvERJsqHOgcUwxIaXOl2OTdn79aZrNjum/eTnIbeW1EeavrcZ4FXUFG10C8YuWbFjCIDq
Vhi+rm+ZCf+91X63vVkXT4IZM/wTf2XMHNfN75/sqEMT4CAm81nq9N3ovWCWXyIAtR9UCdg4j4Fw
k7nwIOW+TEW8b09OO/yGjR4ui0Y5cNWsIj13Mm4yQdbH4lpjpRmSZgNYpPWhdcqyLz2Hi7MTushU
cBXzl1tcgQOBPyGqbPRlNNkqIO3Cj4yixZ2zFzj+1BWYzSaGcCusp1j6NnE1A0xI1wg3L7iudGde
/8WU7XoxI3N4Zhe0HA5EmkdsyupGB5qMqzlyOYgCvPzIYM2H2lPxSfAEXED+idOXFtrsHGYIhp8k
e2Us3RRjOZ7wCOryesIykOnkgGUkehDLiZ6yumHTCu/snzvu/QYli/UnVsBJgCuQsF65N4G9yzMF
frElkGr8mLaKf7onFwXrOLOTEBojjckh9EUWpwJ8CzLtfrUZ+g6XdHziJCEzwHQw3wlDaPL77cEu
ehTaEPFRkpE14Ddf0wJE4P5Dqd1vK+GW3YNKZixrrzzENJw7Jmep7aUJ1DEH0PRSXrwRNI9ik7Ay
4EKZyPfG2ZTGBk0KcnD5NnpuzaO/QNuwosQk4LHQWfqCsvzjFbHP+T6RGoqOloekMIDFxstR0ei0
TuQIybv6e6YRoigf7GIxjzADfVF4WgXBuLOhb5iSRLzJLA8WnDQrJf/xbNBs6DtHJ1dkwBCqsr8f
ywB7CMcCTh/TjRMIfiY16Fa52B8vkW9abo1OmoW31YmFR92zdbWjka0Ag/SeNbQXTEtwA1EDvq3r
R6WEo9P2InvFQ9GsKsmv6Is9WPMj3Ydj0ntNGpRlO7mta+3K60nzGWJjtgD7nRm4SvFmkIIAULk3
hR+cAqgModYoiKzljEziHv0/sGnz9K28Lgh9ZNhhJQH7wAgw/m+6hCfDN+Fm6ofgMApvxQNrvV2B
9TiF7IjdEc9xz+MSZstnx3F5WxV4MM3mMdt27MBnnTwHD1MeNeVPdKS0PiOGCM6kFyKpoDaVKOJi
gICn7A6h2sb7x1381ShW5gjGJkZJPJtsJkz+T8PYuM3m7ifS/XiJBvlLKhaowTfXU6Pqin5FMLx5
qhchCtlITtAs0jQCvEGFOqi6MERviLcXGN0AlLftrmqfikE/l03yHEENzUIIjY/r1MZJB+itdTsp
sxA4kTQueAjWYXaCD6XdAoMit9E2QsincVekqdlkKBvQUBJYwJGXs7IqG9Cu3i75zwy198wLVSMU
J3nbBqpOvdot0/cutcC53vdUDSk/zw03qTwcWkCwnbKdRgWMiLZypXvw26d4wrxsEFd7sj58dOIH
5yjWgzd223orkoj33+pz4spw1xeUTx3InmkKbOK2VRudESqprINXh7Sx1Z8Nrgj5R5UhMA0rZTAk
fiqV9hKvc+vfaEO7AIXBoNrTF2IBVGgGZMVst6SyNXEuTAU5xhCAFlJuZUU2QZfZDcQJIdFPZAdw
omVJt/5j28EFgWT3ApgNGe55xHiW66/xWdzUbfdi3h88mSfCrddZ54QZKA/kdmojtlaR8gw9MoV9
imbHFsdTzuKj/tHF/dx9Tc6zLb0njsfUbiUVqcjci4ZdCYHIpGvrxlZImtcqZF0p0WrVHBJXcbG/
OOt0/lv/iU38YLmCn2M8IG1kjqdXBWAmkJokKLHovBarFbBGFJ1XxQ/s86Ye4/wt6s3gDBDyRDNq
0SYbFyM9aRICzI++Vz+FORuYmv5rVhX2JUX7a790fl9x/ncWFlyIBN4T4cePQakUJq20pbwGQUkG
vdHQGHQ6QAueM76ND+9hzw5wk28dqwT/VHfFOL1g60G6c5hu+eaCCWwNyDsH79q31PnidpK2OK7p
q/+L821Vl6ko1VGMzArIVKFen6sLyYUsfsTdPUWkeAjDUg9Jott1NRWGcYi3JfjZGd7H+u4FbNTs
wh+QEzm1gArdTROU9yefwfgcDSDf1yJdELWWtXT1F+r/VPPbQ7S7zopnRuCcwRXMtgWENXefopwF
xYqtm1Sugd6gLiksGyCRIbGgDdu1Q5HVERlq+J7hMLoIWt9kgCSIMBxTBt4eiYAgV/cs3zjayQ1d
YG7pclV7vFHtqSEc5GyYrVXIqXs+PupcBgv1RdLcyjrgae5M9z5lNck8SjeS6EGmwVyJ+92E5euN
Dczpe4BzU5amtwGGs9imWcDYxOcyZFOV3Nhb4QQT6qilm4veXgZvw86yMXbM7n4pOxdZTbhGz4Dd
vwZoKTiSEgs4D9g3CXRp/XMptlmpasl7GnAHRwIQLqGsIAuX5iIhHqzO4BLxekr6GWp40krGE5lb
aa4Mac2U1uNG1jNn8hpQtc5OmeXy6N7QyTFMC5hM4Dd2v2MwHF6L2XapsJP0wGfT/TDNKugWKRGv
xTM70QNcR5qmRcagKhtNjIdqQUIvgjETydyT/+sytVzyOK7gftZVjPIhD3UH8l1JWjDAu32jPRxN
rCzNU5GB8QfHMDgR3f0Kob/u6WzsicsvL6KWgNcz+U+conay7c/ysacVE/Mp/gAftWRWtY7nxzmd
+4xgB9W4YybxfgyeQ0UNCqPe+3Ma226B0t2fJWz+zwnvkKlYBf5vG/yuXyhVaDSdAmUf1RzJcYXB
NY5oqborcjwdLkYSrhx7swIWPiIRIaOpr2P/e72llwSVdYWe/L3fsWS77bF9nPXFMmBhPaO2X5x2
vHqI3thkK05skOMxoVYyyCzaZFTgOgBU0hgX8BFhKVfNqbNjC4NHPpiry+3ddAAjiiZ81WXSUFTC
4bEiFFssxuNBLBUcS5Vxy+dftB9Sga2YUhjy8P6+fcGTHQNV081e2pMVbS9RfnidUbas/6eWFsPX
N1RZkKjaM+xe1zlq5+OYLTND4KqQI7tEWVxYV421Y0NN63Sqo+kpNoNCeZp3xPkjM28muyvAqDDt
7qAF8qknndM0oWRIHqMcaucJgwKx3fwajWQh/sjsea+0PTIfu9CR3x8yYEWsT89sGLBEWO3OXFqo
w2OdKJYJNFPiX6oYPraZ3wxvTAvAVnIexwi7fBu+vU5JB83zTTm5khDYGo30jDdBUCLip3auGwBa
iv+iLODzWiSJt2opoVCKorxq+pr6zR2g4kzu/QjpnyExTdm0QwIDtQCLnuWP7b6Kc1B1f3/zLZPZ
e4PyKjj7JvTvxAWGNW1HSiFoH08uskMLz4WMRbva0U134NhfumB1RWKaRG5jjuAV2tAPH3Ayshrk
nZag0iWsVyAJitcMh8daC3Vgg8zZzY5y5nF21Uv3PQsHUnjktvVNLaTI5DzWg3z7boXCp5KcfqkE
AtiTYqCamwo868MJI2ZrBE+J6OC8El3tIxUg2bIGIy7q3VSo1SaP3vkcx/2BtcsK05PLQConVVE7
fb80RL/lNAhUe5lrz9xR02Be+SMpzoNaYFVNT0zTUnvc6eDtPMR1x8nR+meqogEcsnP+Z360Jaib
SLQjJuEMXABRceZNJhNITdWPYN/pbHpzy6ZUCQZII5+rgcLqHLts/ZXNIm/n154YYfMZnDrfcN3Y
4Pk1+1aAdkN+6DRm2khkZIszEnJllJiIbTg4cQRVVymOPeImmjveQrfvFpr3zfKx4Z1tLWvDNXep
It3hh45uhkZVHeR2kmIiCYAHAuqjNUfogkrq+N+osqSQpvGDGCUck1rUUnLkCQEb8KqV1YSm3R6/
qWH7y5V7agVK00HJMt63Kaao7PiLWMCQ1y1rUTA5kvb4V6IOZsQSaKgI+pFWLb1Dt8Xtcub43hdu
141pzdbmJn3lrcKVbRimdyfNRmSAYX9cUEOo4hUzVscj1nMxySXvl6lVU13cIVWzXWnz5CYJpvGB
G2/X+4imAMiKiypIpGircq7iPeIZI8X/rcNr3Hi1Pwy2RLtZDlybG8ZOrBF68ljq5a4Q5EoFFssQ
cJH4HHZHDoB9boKKKimJSO7fqLTTDG9QGp5Vn6nrh3CCh/bX+d5sdukhrk+RGMuGRsXXIrvxcRlR
8MLk0yllMsoLvC+2V0rxgzzK540EnXK1VtM1bcgcglgs9sVoQEaFSWhdtMC6A341xmtItCRcnWp1
W47pEzmpZbcNuS1gEZYQXwv8whK+o3axaG2pqVAifXZJdewnHw/1axO+DDmA1cpGnQFA02cJghIm
kKiZm0o99MWf8JgZeuiJxUGtOw8c6WWFo6++/2DF/7aECpfawVpwqofrPVKTR0U8TMCXHCX8oeRV
xIdb9A9tvxRCJETHTOuBApk2Om8n4flicveUPRAFCaJOjS7VMuiIGt4XVQOkjiyI6wGZa94Cy7e5
1pc5u622+uNK0IxJy2sQb/Ac7mLAF3bTf/7vplnS0jUAUaraXu8j+HS2CiJwBXTtKyc0CJaA3d2R
rLA7Ise8Ig2DQDHushPM6avAWNljfXUhjCp+UckF5FnwwhMRAzyJIIJI2alHmfh+bNLu+iUAekSv
pWggkaT9FbmecsjCiFZDbmVpgp8bVilwurSGORtLjaSahD5vUR+n52HnYGeEiVzbGdaWsbQyOpXr
CyXzWxByEc9ZJAedjGgRS/lUBIaZ/EPDUpJ3WO8F3/LEGc8Eg4ip0RIKSEIUhOS86I9cDsazIVOl
VcvhO2GksFXPGTC19BmWqgxsNG25pXbDxIce0xjIYGoP/hWeiEWisa+5oLWJF6Ru/lEcAQYtRq8E
puc7ycQIiDWNpSZO8EGy7Q/iIzjUQY8xJ9PcZhXDq/GWQoov8Cm2B6FOwEpP38wWGvysKxJPYkge
A20/vDlO6MzzTV9dA7mMiJxO/b2Z/NGoFPHNE3XXaVCnZ6cooIF9maDLY4DhqjtCV27EhbbPS05T
vPsocyGroH/IuoZZddV3Xs0qumyFkL9kW/zpEOtAnCf4cyn5Lk4G8E8SyuDG5BRdcdZabK80y28U
kjQvrwQOo0EzQNOSq2doaIhiRBbmc0rVXKvA0QzrUyY+46w1Mf9VpEcIViIZyJs6PbaTfCkYOpNZ
6mANsxOTrY5De5m+4YAH9Tr/5EWp9MVRB37wcakuGOhYawigEty8YLrSy2OdI5ir7b0ptNKxlN+g
LKi9rNO0tAtZNyWkTy2IDGyboU6qFTH7biV4j5ol6Fug3GVlyFRBXSPMUgfZNBXsHbbrYx+sXmtQ
ShY93f5dNMLzI1rTB1QWVIfV7yjRgptwC8iSyHIAjGrBy9uvoJ701spag11gQOi7PbFtqDo/pc9L
BC2E1v7T11JamrdS21O+GYNXkFa4s6A0RZ06jgZoRKhs0oc1wSwszU2Y2f5tE7mBQ9nH7923osPo
xcOao60WXBn55e38vpqrQC6y5qiE+GmN7SizRTSSlSm7tSMdPnpS/tI7ZeUKEBplJ3hENCttknlX
+GbgKKX35y6NHDsq9jDR523a1MNqQUrKcUhWsPJb8cH9QF0Dnl5/5hbHpBX64BbrfWe0rawqSbfl
avYlM+pgeE5dZH0NYIoGdc0klW47jJKRaeTOXpfbfy0Xa0JA6n9Ia/Q/dMrJw0mi33Wt+ZvD8ONb
5XLF+pZuJ22dGihwYpcap10pkglsvlHVSmOcmvKyKNqU+KdhFwEb/KUtVrZZmN05NR+XASIXg17/
vmgIfv4yY5txBuvstK2jX6KPB0LddU6Uc4QoVaRGKVmtKGe5uNEazwFEVoaiZReuFSACIuqBZxjN
JElxdtHqbOd4wamtjE0DdV7xkx36BNI6dbnHbWv87K9gwSV0Arg0ZaEy95VG7yPpaE4gx6lPG3u8
/aGcMSDxc9VnmlUVXdpb5eyaNR9IBhPd+5e+mboSvD8+KA+27cmW+YC+XeOfkd5IkXKYBHrN/nHC
jtvHaWp72lBk+ssOYgMn0HuYQlRtpcUxzSt32msfCDGQUudJVjrfB9bIR1OV7ro2y2O2pbIUme7k
LqhpC3b2k3stNkNFv9Yonc7jLzh+i9DhnbUPWCMH/OgBg7cIKLJAe0VVOfFP9tYet5PsEljLHkJB
oADPC3dkTnCpY6IT3pmLOh7PW7ZHg+Gpkq5w6zb00dWuqoFbiXTmsYq5aMfHHKQnAqgmDFdtd+SU
PgSoZqcqegx4R5cBJkYnRjFO+J434uPWpleZrvmJfpRXzxcRApI2sc4UfityGc0uOYYtBbTgOb40
Ruacjjw0yk2GDVYvuixq2Gx+G5YqAXId0B4vqr2/pi02FGINTckN6cEuTr7102NPbck0QS6a5u1f
4O7Oefnv+I9r7hJFTFGiVdTheZ5Cg1P39WOBLGGII0+WgX5yW7JwAV3ggh63BUkowWNtC7HsxDjF
296YMzCiuAtZbVfC4Xstdr/njCnfiX5rVv/A8P/5rWUoeF9l5e60Pgdqx7nSCNm26W+RuzUlsnEh
NZ6gRhW23t1p5s7jElvgjKE6NJgl4tR2hKMjZuFMu47KzRsUyfAqHODf3DUVgIJ7fBEm3W3KmpbW
o8lhy8woGsNrUKLccLLrw94kxO4E8x2qbqSHFlV1GPbndrc7jXSKXgsH6EtBJD3CBnAtTZS1CQo5
uJDpTXECom5JyP9YGL2uNaKQD7IME0nyx5RFG0cawKCbwJaP+kmvtqMnzSupgbXZHxFKFPE6Xesy
jouUxxL8lRBoWuOpf95t4xrAKhQ1PCTmG53EBW837/AmdgaICaJikSn8zAElpZZcw4VnveUyPADN
PjTEcRDSRTk0RZWAAl53lpCzoP+i6nUr0vsCru44ykBAxR7JteSK64Zp1i715o7CSOoNPgp1rBTr
kUqjPBN/oT5bH/zJ9d530js6RXN5YNEXQBuhmyaYgiC3nM7jR9CT7O/swnImNLleknTGvBlNgDou
pOHS1pTSocSt/Dq5n9wpJxZk02OP72kqvnw7sTeDYUkhIc5Ft5yDh2gfC4AgXUmi+3/rjUElI1+O
eFIO5poP2qW8FxsO9VTaX5GP8kvbmkUCpk93AXAH3prL2M4N5pMq/sWNpN/WGxtMsoH5noMfeQdk
5laeuer+f/3kBDkQ7n6UW9aw1+PEgCq/1vIFOyb7thre1USeU3lEzmeT3Ccp2mT298+mBXcJOBpj
wa6odeBYGnjtl55YuDvKhwoMrVSl+sUaUg9qUfjn4j1efvGuGVaJOJ8Tug84cTe7zmSklAiewh2h
0jjF8tRRnJgkd1T4kDLJetky1ZRDcRhjCK6V4iz1QYc5tfiGU8ff1pBek0rWgsC69p9wuvQxpIwn
CSDCWXQGmTVzV0Wq4wjUFjO8PKTHrv1EKvpYM8qUGfwOC6i3+YcWTl2PBG6lCPg2/BBBessQ78Ka
oPWC3Om6NtmMDfZ6Hh3GCSGSqdwT+NdgRqnrHadVpcHYZgtsd4zEyFDPiqyLCkpwRmoXzIr98kmd
nmhsQm+znpKyBQyxQj7AVIZOwNNcXISU4JRrCnzG+TkwzGbs2qg9oc+TIzII+USjtUqZrgwg6cKs
ssSBorelWKWTveZ6qUWoNv2IuSVZ7RDps4Ym2+3v9+Jbw9A1QRCH4QbJ6l9bxMBxx8yUivKS/MXa
zGoHfb3eunv2mJaKkSa7lFgWKMeIA3NgAcYpU43F4ZtT7RgheuTX9qd2AS+li+R3M/LFjdFX9V3D
2Pt/dSdS1BWba3e8wbJdhnisN4SD0m91usDYq/sQ8iY3eLy+AlJLJ/etYLkZ90yywaZh2HBggJlz
l7FCeE7ixDk0ysuq+yqOmHFhWPmSfQlBSeT1RJYygnaU1U3VvoTxa6eIyff3j0jPhnyXlUJalQdw
biOH82oyMlM5UjtOVXp9H52OVYw9kx8HRfCml9VUfetZZVwAYoWfHXreKiGerGd6a1NO8OKXIVDA
cOtiZ/JxX4uj8aPVv48CInmtLaoPQVgXoXJ23iPr5OSKjWxhrF1XKB7+5Q1pkxadLOXlmL7brVdN
eZdjrep/HKU/v54B79pujvtQv0C6JDEx7yI8MsbcsCPDnHxd5JHD4QQzKIhBZcyqTWNGD3AmdSE7
JJFoUsv3KkgvWHgUfMaYsMhSAxx/7YY2ozbivxcsX1RYx7Mka0mFRw9tXjEKhxuZmSRqQ4dNbiYq
33SlJgC8mCODL0u41IslRzlGOW6TuTrUIK54RTfBpqRRgrjhJaQ2Iqoa6UZjAKly1n+3n8z8qCLB
CbJCh6qfyHRMQj/YHF74od8LPOsIdgc0fEiEbUxDu3DBuB2E5ux2maaTCqB2Bhm0bU4CGT7/0jlB
UC4DgBQFEvhrQWlhrq+YW6XSebLsZeBMJbWP1/qRUIOBr/U5C1NxvVCc48sDv4Hu7K8YE4a9ZJ0H
+ThvtNdgiSHkWphgZbV+Yvujg005R6do/acqUSW3sizCO+rVPwtzMZouWFYJrjP3e22jFrZpSJzO
a087eVswowLVcB15/tqZKuUDWC1+XuX0/mvZeHw+o3GLV5DxpSV3Ai/Hb6RCUzyzQ76IubUeMljd
G2VZ5mn23DbGXK9MuCD4M/oCGJpnh+FjJTnepU+Sz9wabTJ84Gf89/ArWDeTahYUOglqsUp4yHlc
DLONICpOEEsO+8CPIQcjPDMozkH8jctXDRBnrYAI0RyoTQo2OzeKCEBO/dnRTqE9L+vvDigYF5Jg
dyokSIAE6uni1Al57t8oAIM3/mXDCAF06ZbCdkeYV2NUeG0EQLo+SmJfmOYMMmpYJVSdCE14aJFm
QbM6jiOf7RJAmlX5ebeVb34g9ir3l7/QmOw5V7ndp6LRsAeMlFvuR9W7+fmQJWCAiegBVLd/ps9y
pRDMwct7w8psD6JivOHXx6kGfQeb1bdEwAms77g6PBb1/fXO19M3hn6aDBRHihVI55kl+m6SBoLm
iDYuXCafStm5ieq8RVnOeGohDi83mGESss5fSzfAUKeGHlxSTp8pANIYjRXEiFulC5upjzOGpOdd
JHpXFuMw6eUNXAofdEMzsL/G1k545Vp/BHghq5w5wqR2sC11fyguXA3RFo5h5k86Q2H/OoUDEFt8
YsMMq/FVuB96ONCM4VwJag1MveZH2I8tR9idYPtxsuyOVmpvLGJj/D3Vlg45XKDbmXnCOy2w2NsO
jOisPDHdS3soAh2Va7ednuiUje/lblqobbrfpyqEMcSq8VG4iM5wApUKv8/l1X4XUqirnp7/SIeJ
mzHOH6h73wQn8dNGqTHX6rYR/anJ6FMKGp++Ld1xRFNhCIKH2eE9ItFiGvBXp8ZcY1KVwqw3zTjH
kkqrT41qAwbhF/2Rk9kBKGO5Aty2PEikceD4CXuETQVXQq8G02btR5ROpf8RxLbdVYlgYNvFin9a
D+JKESqKgBOINg8JW3WJpQLwAf5K9uZg8v1USSsPFPnaubwigdH0+Rh4Dt1/DicXerXa4gur1R+/
Ze3HqIVA6NDxVqeOLaWjkgaByak/FdhuYyyMpWPPbmQZV65iM64NIT7kTJTr16p4zlbjy1dh72ys
GUzjS0XGINGxERCvx4WrFuZGZyAPBhwSUeberBOLk/9BuRSYtn7FUvD6yFc+Ogv2aHjx6SoBCJh1
tvKnHbnWifzxNR7DqIRSF6N5wjjGFLA7unjvxk9K2OFNj1bzglPd0/aICJ4xOurt+m5v2tPJX6OY
pmIh4ZlMDKHoRV9OAFs2pWhPkgGfrOkarleFf+0Vn2TC0r+pxGr97xywkVHxI+z2q7dyCuEb8knX
V9gXzIMHz9qjoCqvh6NE0LWh273YeIL9Zlwy7N47LnAyV8Nno11b6BW+hcZ3umzFmS43RST336xR
HQf4WFeAd+jCxdYZg79ImIwdH43A2aCNUHAZ8Z7vRKJKV6BxvYPYNnFbGmmanJ2iRznbW2Wkr7ug
uE4sf3E1PyatBNM/fZoeLceZewMZMkMpgEzMs6rN/jWpoFuwzqnU1NydFyTcejWli74HdMBx50z1
7DNk9WFEQHLSKhP8+CsyeFyeABSAex/LIFwRVfuuCqlg2S9sWAP91dZl3w7Bq3uCD/YDk9ThDNZV
i2japxIe2DrgMouP85pct6Fg2Hr+2AyEzqKhvRVF5m+wy97Wy9jdo5pTnsaBXBydXR4n7nGQcEyC
QpdKMwKX/GSAN2cEUhRp63kMfu0qjcWD/1I7cLJrZAAZW4O1Mnbnhic3aqSc/uJ3jq1ZC4kTFj23
aFLS9e6ivuEd1q1mDlUh9Nt+/sLZKHGjbbYgTA1BtNDTlk1PWCprJD+8vTn8OLJwrnPnNK0MNEKV
K98c3xCqmadsKP4brlVxF51zLNhzFot+h1qCutb2Lzr83H29CwW5+KtdVDoDT+ajkgZ1qnqS8k8N
8uILAEJ1l4Xiu5jP0sKLiEnIoAhjnrWpsO46NzjJYq7S1XmLzUjZCikSzNTElm40BhQrAgcwfRjn
pHEqvud9P6YcTP6wJq/jnNQPLeiJ9y/gmSaAKpjoh8vRiqTHn7j3q8VL0vwiIN93UxYt2xeuRHhj
zn+FCn6UxSt7yAtEK2eYEx00ZrO7+07vYHZy29tPwNlWOzcLW0BinHRNprf10XiGicMP396O9gCN
KTQGCW1fSYZIlaCEp8rGDx1cBNL/7dOzijIAspsSDAome+WNWRTpgiO67snHc8BBSYEu+ahfD6Pn
V5d+vnA7fBT0Tfr+PvNnkOQf73yqs5Jn21niUxFIMZweN4qWvh3WH7La5qDu2BvYZFf8dfmpCOnL
6ImB0TySvY2TE4NINkKhSYm7oskBp/4bPTguScjADn1mI4OQ0MuHGf8/QcR1Une7gxXDYI1JMKQK
FruiSVgjTMqoraKf/0Eix0Dkcw8zVSBbDBxkiOCZv1FOwFShoHFpZPdqviJA4aib2OHMFytKQyg1
0mYQ0GHk9WMnWBm5R9WG7TZgtpJ2xxEID4dW9aJE3f9XM6t1nt3ILNtQE70jmBgSsfWcnja+tq1r
rDuPgHws41Qv1cqwNl7hNjl43sHU2SoE/nmLfyRlCVNqAUH2JK5GHyYFZSSNX6fJQV6UaB9Mnm15
EWXL965pAQQZnJOKypGZo+BTT+TTKfpWodGMFcBM7v4vvMQ5f3FYL8WNcW7C02RSXqO8/4COsyMp
pG6gA5doWA2TTw97bu4QY1aKhpa8i6URcSiK/yvHnrIxaVKyFotQy0j4pd2eE2aBQsDlpVGZCMui
olcLtExpXkrzqtNoVDYTEySqITXyp4hLGVI6u24hX45n/w26WF+2qegGouyD1pWoDc+jMnXScvH4
OBdqDz85nrxQJ1hMg6VuQhf7Wy6AUMwRx2ECtq+jl/uGgCjZpMYSgEjypwBvMg1r0UFiXBMOp00b
WukP5B7w+mtbqbkmH7Jpnm3aE2HGIAkPe1+RGrqZV+AstWZ4ufIs20EhG+KSdgYy85yOX1jm9h44
qvM1PqefiS5aDdUvqM9ygcBnEq5mNNn4xEcQ7raTy632IToIZboqOzYPEf1/KpvBwnYg51iSsus3
eaB8uuRG3Tjm05780foX4KWQ9GpwRj31yamZaclfFDxAnpcbE/ZoYieMMTRSHxgFoNeDS6UFUH2b
J4OoY6XxqSuhYKu0IKnciYaW4MYtiWHWiEbZp5oyCNoiM4gA8M435ypSGBQ3MSAwhKA3SK6nDKt6
DGicfVG2v1HqhUEqN7fQbj+XKpfKQJZuHYcjI8/zakvSbNrdR0tNvfxKw5wHEq9MT/kZXaLpaSpT
/U52DxI5riySqodB0q+NAXYZskOGspvEboOrc0KUcYjYg7uBdQHFw9bgVrVlMih8TRF1gFNdrd2V
I99ZrDmltMYN8LfUznj6wJ8gtErTuQsdZOlrmp2m7hNV1gYfew6fhhWYzMQrqFguNo7Cz6Qh3gUH
wIkOiS1r3TB781mU/7imQypWN8xlO8fVvkTgO96zYBYf+88mTWHgzxlrGYY2Z3TvIBhu0tlTvARE
/NINKEkcdy2D/AtvTi96hc1Ec6apOPg4u5QA9xdHu4bxtA2Ys+ft/glYSCu+a/eug0dS9YICANlE
4KiaL0zGrMfsJLYdIbg9QQzdaahVkrR2UQ8qLseylv8yb3rTKPehz1MHPEYf53pnutn6WOUtM242
p9XdUaG1u4C82gckunNe1bbyJiyUAW4p1JuUg0KUXAaWo4ExTe1kC6utf6Lle3ZRDmeEy3dKo8jr
mC9sxeumltl12Z0jTq6wQoEiu633XflmvM10xoRAd5lfHvITQ2/4hpXOY/63CCixaKiUmzr7K1oO
FF2qR1bBBJFp614+G3MTYxO6Q0aUukNZcneFjbJqp1EHwxzbLL7kN/jF2JrPYNriUAaEMk8cgKWa
lGWAO5pP5QPu1Ql1ZcA4tga2xIH5gk69gdjSiNEdvyQxYaVu51S4T0XoQTI8YKEUoR710JO6sUZo
0aP9RVDs95joxw8ZNIQ8YtCIPaDlJtz+LP4OKEe4Gp+k2xWyMq/w5ieIccQLdA9tPLNS5YWq7akz
TnfSKIj/cBKX/Xl0M0/vCRudlBDZobKFKXW4gFNZJQoMMNlzwk26nm0gKjQvdoAJe6+ATOduvwPR
eNBXJVjTl7mrvV2g8qEoJw4hxqcZTQjJyE3aOIswYk0/VS/t+HSrs45vkiVoytXJrzqJ74kQAJl/
4fFjXtjGnPYwqozUeCcVofWeIQ4UsIy20FRbuovOWZtvqgr4G3nGC/D10Pp2R92cOw592Ia87pM0
rUiWgI5JFN987A/M7bU24q5yge4+mmjO4yTEtegnqNfW1aX6L9VIPUj3UK+L3jcL12ZT6J/LBX0v
bmnVMbSIGfmYpFy+S809gIyqzd7g7z9yxaeD9Dgn3hVPAVigbx6X8MnINqdglDvuQJ0XhRQq3Nqa
olz174G+q9+bByIYdhAR3Y3D7yBZmtMNkjtafPGIeWmiSyhEx3/ESoFR+hyxahHO7f3RPetR3jBn
6m7Vuqzz6FGMggiQYLtOgVcEoqn+EHHbIDXoRwso2DuXzOJXgW7Wxd5OWoWYEok55CqBR4q5Rqs+
N8hXRPT2iGw/BAriXI2c1/8xK5B8+NoKigYVvDnvRbYbEtXxnrtsLfwZa++rc3NvUeNyDWyNoe8M
mXN3eDHz8ig55Jxwmzek413eFVO4YKcsjxpuB366RAqC7lbo5v8mh3pDS2lflR1TkU/GFt33vY+j
/JODIHZNw6qWruO8K7MdxlS5O/YUVu+8u0YM+pcjTQM2deJNcysrGpoUOM0w7OezLNCDTM0s77pc
jRXwCO+VY9A3DrlA6Yu7XZmaMUcbQD7NOaYJjBRZRkPxQ4DRwGAcbSxWP6bzCQQXsG98bsRql50B
CV/3qxYU1SS/1BdwctLKJbazw9fFqHllKDpUfKkoM/FQOQsczccZoaMQVueaJ779lGtX9OXU3y7D
YrKGHkAwsGZIDPilDpw/8HSjbwKu2XFIr2BftKG/I2idRsWi/jBY5O2K3B7nthIxEPQD2qSNCSIM
RmjxYQ6xvQnVUdCWk+4B8P8VnQS6CYmSLAXCM1Zrmzyz2uJnH2NbyvVqhZeVIdLVnAOoVhelRebp
q1ku0H85YQueZC7noYsbFFVPmAU9aKDKSkE2ZDzlXL5kRWW4BenWLxBptjtQLBoI/5l7F4XvOuFo
+wm4azHNwqhvRdgeNJi82zLIfZNXe5zFFYybbGluErg8y3peKV+TQ8/YQMgBjkqZjYrnowdoCWKt
UGN1tGSSgEZgPiTDW779+N/vTT1S1Bjr7fxkrSU9wcZEiKF+zLp0v/pLRqvizJbVPKObLAepr0C/
GvLdx7hLFTxE/qjaLajlKEXB1mCC3CYlvU1gP5KyhDVNrjYG5hXGnfSrLeJp7dNuS8ETv4TvMeBO
8dY8Vi32LSOyEHZiXQwGWfdouUOTppi5+hLHriV+azeZ/Iz21NvKtIe2u9aFVoE3lBTTCNFYVL80
3H5SRzc3LlMjYSCG5KnWWCRJxuFVYh8Vw685kWK3lk7gjrsL0an793vbwFdVzyhDgA0Nz7FBoSLF
hxIFdOTpz/rwwTYTK8ExErX/S1GOCkyBaBslEQY8MVx7ASwkBM1BIv4rf+T6os2rSkjokwTqjqRJ
zbiZvhei8PbvhbElO1Ic1Nk7F9mKaTpf7JXEYEQi7U1FCsQSrYTOrwC3Xw35FJlGakgxVOtJtEgS
xRLGhLAp7F7gOgi9x4x2JsHVD6Y1TlQhLYXZPzVTto22I/154MGRFEq3HWCCMx4+gNA89a/J+W3K
2PcWeAqchgHclM4MdVcSkeJKCgH5tSkLNHu8QJdVwQ4A4A/AxlmbU5KyrbskjGjcBQYj3Kj7Jrkh
Oy4ei8In51rcd5/N04l0eA+9qfVOIpBGq5UAIyUcdVs+J5VWw0Le9QgLEJK064oytlv4Ft6xPoUm
LdOieggL8uAhNPpquvkaI+XH5LXgg/dkz68XR8WjJZIldiWLeT7pp0U8XCYNLPKAo4EzWU28baLx
zGwgTfr/7WjGJSays4DraKzt7MjiXGDIbi908Eo1U8r8R9SMk14lJXGx9C44SS057vc04+bCAeG4
cLBwneUODt+8HxvJMt5EZ+uX8dv7Tc4k9/4wp0mcjWMz5cPS7aebLPpUDZlViEazdv+LMx+Qqwa6
MXsxKz/wrpDV1R5Pr7IrFg+XH6GNhHptSEw8e6VFmZ/X5I8izWs6izPyC7D9//nCAMTGggHxEaL3
1V0kr0fnk6p1uxPTRMsgNj4ZiRl55Pqnu85i3BpQE6fKRw/srmWt320p+K17wHTHaLQhQCknFB/t
CjZJcEEjJ9rmpdwoQBptG5MoCR0UUxk8z6HUz2IPJdZz6CAxyE36Uz7+B1updiiMLLA7mYwY9x+r
NlaAJGhKwZOkG5zXMnnOYYBTFKGPTrFkuUUDhHTQYMHJFND41Y5Q6GtT65JCfznaV5o+EZRvT9WF
d+aND5Ej7JsKDcTy67mxMnHxAlQoIHQdauPiDVC8XsGuvLh96wTyJEJf6oDjWH/zR5VUj2B0LaXO
xu/XNpcYy7UHSSnVW/EpFtb04ZdB4lqwy43SH7x8lnfo83KoHktkI29VDHIhKLMZSBGaRdbAHSTf
B1vxLJalNUfl77z68zEuGkSubPF4YVq4N0wWyKAyzRsQwQgSpIxyBrUVlxMwWMeXZtocQBDSPceH
9EnzioGIVhcMysSijTqUpZ7/vN3a0klalzSiV8bvcbTZC4ohJHSb41eSkAdTTVgVJNzRyfQ8dh0F
g1OPylOFPbSyv4Jmnylr1EVTScDu2L3ZRJcJPElV9OmwGUH3x4et86vsmcTNCmnt7EkpBCcSxsTe
wEH3AL0+/q1AF5LVhIxRyL8CuToCSWCEaw5JY7zuY6/izPGI91jjN4qRnP9KGDuKnUs8oAP4F76t
j71u1aNEM8AIe/lQo+0JEP0Ar5NJJ45F320rMnmxPyJoqoV0hgGjQp3WHwcXUryfsKyD3b7mHcu6
N8UJ+hhChXa+e8Oo2XaJfq44t0siT/ZKhrGquqNt04Co9CPnp1Sal/NI4OZ6v1BgbCQ5WLmL5leC
hbCicFHko7YSYRCuHlbf0JSdmfKatp17FKPaNgUFkzjLHEFLBoKd4oE1RnJEDBR7c2MhyW0YZtWo
2RgOtbGWvWOFozOf8tU876D59+j5h+AFuxLgfYQyb3Tn3oTtRCbnP4cV9WSSJ1LbNoxo1F+RLJ3E
ZgHKKkM7Krldomj8ohYYETJk3niZ4U4lfB9IQ36VfCdPWRzMf+L1po07Gk6LAoR5Wj3E9U+SSN8o
jLeckGVBKVsVyOuD8wf32RHZY7SbuI0E3ann0p7dhB44Sdvqj9uKDTdHNnDTqFd2kfBSWqvPkp6w
G9l16dNUMUgvuIHhkS2iQtrLsfPq6lSUGfgOE0cszvDWJRN8s9a2DaKqphGE/7qZOnSmJE9gkNpU
ttreax2952iN9/tX4AejsOLUSDCn7dC4OddTAQsxeOaZGpO9grlC73p0+fQsSx6KIVXwv61WOkdO
ulXGuZPsJDay9bf4+tfOtz7B6+zvv2Gcph1oU7p9Uq9z1TryglUaObCGlHjCBUZ020fCYxi/Duux
BmzL8nCwojgiduCJDAvODd9Psd73jBQDWWp/FI82/+kej+IIVQej92p0c6DRdJTjUQ+QObglrD1h
SejOONGbxLO1q78apywX9VqRRZcbTDC0awIQH++ONJ97Yy6G95qu0KojKj/lMpbeynBBlz99u67k
rLYiwrZoelXc8K2n9NFnuy/vFtvphx0M/QhfUsSj+LdQa8yBWLG1PZYtikl1patFtc5tIQaBbTcw
FwowAIDwcONxrL01G2AqcGCZpUAJHsvOGnPsDG0LtYbhGbosWq+ZaxWQAbagvjQe1hYRkmFjVK1+
GyWMkueUMYKCZn/8PNw89/5hZT0dOwTGPyJScnDFJ7KUVQzShW0LOCR2GQ/SajSWetSk3C1nWxpf
f9eD26X44mV2mD+/7X4569Qt1l55fCkpGGovL/W56SsoVQ5sDtcyf8rF9EWDygsf9MZmcik32Ph9
wNz7WvvMO18L3+rX4bGlDeh3m4vPCD1PvvUoU1WdzzAb6iJDEHUmLSI+tZkYNUkaRU23jFmsZt+O
0r3lwUeXyWvbry0tyEoY8sV5aqbUnlFfLwOpmP8MRG6fh5sQ7kotbyGznDJY7/6jiBprSO6dppmP
rCAoqraVc2U7IYeW8mfkvcaegGyU8vyYjeV3QIwo48BWXV3UqI2i3lZp/7S9w9HQF8gHiJeYNFCd
YZJEoYj88E6biiUWXmSs+uhZ8TKiMHzji25CK6tO2cp6PkZwA/cYloS0W8WuZpqPHOJ4bD3CZzY9
ytJ0u0hGz137i+pZSlAMHFalB6vzNfOeTcaQYwU/zNC6B9PR5nD9MVRkNiZDwhk5mcNC2yVmmRki
AQx0uVYuzx4tdS5jNLIlm2sOdbG1HaPZCW+k83S3gz9C+Dny3EP0IWvdC3zwhWB6HPEwt3WtCuFU
FbvDWE7mJ8kW0iLb2FNHyW3dXe/mZQvKjEm8pkjoDJD5b85POP8HBAL6vWka4pYbhdhPcKnhY4uO
o8fPSACuTlF5wKvR11dY2uNj9dvjNM1pBXGKA0dlbM1qAlD8bJksmLpaDZMJXzu822CDOh6eaV7G
Vk2pRuSeGxKCPWJik4jd4w0Rf0PhhFv2SxjvWAU2ca+DhROfCR/0lBYs4u1DAmb/GgEhp4tsoTs2
r84phu+hoj5qm5eEOQk2Zy06PwSymdhnsn0kkcCy8QYx3NsaxnGkLmbI1fFNufwcCA/b1J7fKIDp
yvm6/iz0kGgnwYZ96LI+TxCNqZPGUqh8OtUUB18pXUBL6urXt4pr/o48LpSInZP3E+Ky481h5Wb/
UOIgrQtyDPREV6xjLQK2VtCbKgBVuXqg12RDC4hTzHv+KLdDrH/xwbmikRGR189LRu9fwvVtnSB+
sZY0surQKjkezEjbjF408HqCE+lfORNYNAKuHTMtu9so3Lk+uPfi+Jww6H7LmU/pmn0/8zTHFKyS
9PcOHjt8cu+7+4AgO/sFs4u1v6EM6f6PBJElUq29lPY2saWKiMFpmi6KJSjCLLMQ1Pff4IJ3ndit
qIBb3CzirPBlHj72TpyZbe6p2Gifduzl3NXzZIocUr3IxLK47bApbskEfvI+jXnZ4WEP+GQs52SH
PXV/KooPgVhGlT66v7leD76XQCBHwsMwMhYouLg/uKylZvd8bvgx+GOYTNvjn/zHfVveBYcdUFK1
NRafouMf/9gnFzxBWxGMdJEdPE20T3CAfymtAgwAiZKyooq1oWfpw4c9q371JA392SlP3v5a9P+q
DqXio6fBAMD3p3AN2bgl6zXqHxTsHKu2ng7jSxXGIbuEOkWMiGOMhzVpcYGoodSntHujxvDawrbT
XWueJFhfFOxVBTup9wjRrut8+PDnGonRrERsCffDpL5HTgXsO2v/4g+xN5xm1R79zg8VT0R8WBqZ
371NJ4cZRdFx4/JwS9I3UkB/rvTEDi7MMESDTgY4tCyk1TNj9NX/N69GqDU2a8/F+aCuz82DB295
QjI/KRoZ7vsJkLkbLN3TN3gQMGb1LIiVEagkNyLi4iD7HhW7WlvVL5oKLbrR1J+NIZDQ0oGEMCIY
ocIxK4Esig/nJaeXf++0R2ldSOh2bxVjBLj3igyj20CMDSYuDkb4+RHI22TQQ+TyH06DdKoLDsxA
oPUq2OqWTiBaO1Cgd7sGxUpZGyBj5yWhcTmZ+tArny0ERZBR8NJrYdKjWGBtRdAJXoqvtjlzSZig
w4zXZJnEeWEC0W44YgI9IEsstpz5n1x/kYAYcZTdoFB4EYxtXYth85TqoZGJi2L64uIAxJ9TE9jH
eovO6bybbjtGKMGvKdk5h8zamUCpvg4QcyI8ayfABbMn/+MIYUubam754Z7ZmKCLU60eZPe+zV4n
3JjujKGpnYk0MNJLNNpIKv8egUbPpYtWLYCo6WY6fwjk6OLiTCOFt7h/qLtDvYygWdRVG8r6OZ0v
MGivV2oZJW2MLA8NWYdSnFUfFW1FuBO3Fc2wjYI6OKZ5W8vNl2JNRDYJ3lblZozEoAiL/L0xTosb
YgMAaiVgfCYBn4uKBz1JXmFanBcvTpdCre1nTOvLtU/4zmUr5dMDD/kw7vA16Lj4Acw+VMH4IAFK
9Lcds0orANXK6LulsF7sYRMPEnpxRD5QLIzdpODLXp4WqXX+upKh5ZapWLr1gNFLGHe/sD1IwSin
kjFGOZzJvrO/ruDdRhtcN7L6mIP2+zrsuW5WCgaf3FAz0xBYLAQthy55Okq0B/N5DTsJ03HxgbX2
9rXoKC1KcI85VS5avrdNph3ozJRpX9JrnaX2/C/tvZlBTdRbWiKEqBsjKslfPHKZ81CQh+7b2q20
kqVg2ctfJl2zsr1ZY/ClWAvCRYH8fEo/OZ5xF07CFIMr7AEkA1+OHdojAh2eeIMw44KbTWIOBsYH
CDmSmk6BgPJW76gShBflJY8EJP4SzOL0CsIyX90WjdH0HkIZO9e+v5MLS8hIbkKXLs1iaVlrqIaN
VJOzO7smP9HdSvbBnBypO2uOnN69f9Mi5y7hdvfPAAvKRfYJLNgh67hTKBtp5XAB9aIn7Y6Yx+3B
pIvVAE0IdnX6z1zZL4HRfFjxq9r2Uc8Hs7dIAqy192OmSEZUFQc6Oc8OgHJSF+zJpXKyJLRSyAhK
1MF1F9IfLEmFt6Ay9IJnosq5hdl/dAuNuMpkVoulifSqds3Cl1LDSBddgK3Vt3mzv6bMIIqVd6Jm
H2pGHnWvzPRfobji1RvxujhLhvRu5pKvyGmBea+631VVtocF+HBzNqAjyZDnviXVQVbGjZwg00fH
f1+vNw7tLtzeyCuNTPcawU745vX/0zkR6sx24rbzh7Q8hRFXiDBQSgXjAMmTTIZA5nY7j0EzODGh
Q5VAygYO3SeJT4Tnzop526Uw6JcqU/WOBqTxSGzo1ih20ou/EY9JiGXJt1Mn12UA/Q2TKVDa5Thh
+Q3y0Wi3zV3ihTCvYPoAVijoxrI4XgVSKCp32gDkf7qSCY8rdrxUHHOENvSwBZNUknI3iPAw1onv
LVTJYq2e/DEoTctgb75+oNFsY6HhXOM2TlqacCdDE+pRPGmCHenC3uhEgi6Xf2TuRP49SNlUc1bF
/pYtF+/Wr3XX64qOWFiU9+hYlHkBGZWkzpgsoW0JtVdP1UpbZxXotSF7Sszo4ymc77sSZJbmS4K+
6Wp6T7kPqXrBFs9LQJntmYYFYnQmHQjP3E9oxD4e/CHvPWW16Mhd1OnYsdGK8qcC3h9an+qVLm+q
14BQFBw2w5mWEoRDZuSJWRIyQ+qcVINqi5Wf8xr6PhqwoMJ3T1l5aeyv7/skLxUKDHP+1UbdvVuI
y+gZyzMmaSia/dod7opXEnujovKALa15Bzd+pOoelmbm/kMW1VsdGZr9Tw2Rs0OOWnoNwL7E/p9d
I/IZU0Y/LBknyfwx5tyXDgmnJahEEB/BdGybhGwRYTtNv7h+KA40h+KBJzBet67v+0tkPjuWego2
lXLOOALE+97e5iP2zUQTAa+MWRQud0cDzHDvjVzUzLL4J+D4lWvW8mCmK5HjJNZXhDGUhAsAs6ZF
c/b3uK/Swm81n7hf884PxXnmk42W26/fMw19claAYORyKMXb3Yh+4QtS9WBxyFoJZoV61IB1mNU7
honavmvF2fWb4d4tI054lj32lmd+qkMU6rg2h9saV4NZO8Uuxv6JZIqdvLpEYu+RAt+FRtIrqVA2
TGjJNpGCuMkbYZDFEktXhyDPO6u9HEEcjKqRpzgZ2D4+0GdMuFBOVx6BvwIhWKl4/PMrPkVwiWl5
J6y1EXjxsnC3ptY96ar09goQOh2BsWHG3jFOj49RaT9DY7x3NtoZkYhrUjrepbjDATIIKJZbmeoL
mJoHgdfHhZ3kaP81AEOa+pWSA/2NWLitJRe0kM95IyskMQNhWes3k85f5Yk2oiD+9FkFmHb8s7+T
NG0XwykERJO/3WG2ho2ZZceF3LHgWWtiUm0DgHvX+U6ItPcyuq2FydW/+z0Py/XXxMhmXkwFU+eM
i/m0ZleaC6iR6N8i5pk9aOPYXNRgD9aHDkNNU5CGQEahfqv9mOkxxlHIJQfDZWvTjmSAL5cy6fZR
sNXszLOYDMt6H/rknzi6QDRSq3A1z6j8vitGujoyf8Zup1vCPcMgxDGGtQIJITALDPLq1D8DJBmf
Am77/xr3y6UokmChHmvHkJmBAWak0rs8/9rmnDOiGwiHqvwq1/2QFI62Gh0ngpkzzIZ9MwjR/+1m
0ANak3J0b/vysnnM+v6yZ3hS+JUooYkW00u6fvf+ol/IeqbbAxkphkMsa9M0lNA4dBB6WqjBwFnA
vMwogwMVHUfgWAdwINxhTOnek57OOVKV8SYFLDO8rqfk6Gs6/bKAwbKYavbeqOoBX6kf6UnDYusS
TRP8mh2qqHJZA7eYB0VCNyTU6m5AYvhPS0DdnODEdHbG+wGdEmQbs2NOeAqZhj/mxD3gdFZqezzc
gT5q9EpQqlMd0E7C1s3uVj3REyHhD3lh4845lza+9j65BbZawwQZ/dYJiaL2zhpSHZiXC6xBasdN
G6hbZnReUQY5oslXfUBhaf0Y2fygGoiQ0+dju9WZtF7GTacYmLGmpt8YWNdSOI58s54GfVV9mAaW
Dls6al1W5xSFYLTvabitm3Nydtjg762z3KLVcV8Ae2p9/jdsvb6Iz+U86F5d56cMkFHaupS/HX4R
L3Z/vsbD1NrULe9T3k7mTf9+jR9ApQl0c6LBRm3jrTJtmzvxJVhaYNiPfL2eN7Hr5H9XHfxlFKR5
yWH7A7481ZOfiaZWNPUoor0qe1K8k6PGo3jpMW4g26Xurxwh29Wvu5IuRpu7GCT4LvZXKHYE4WJ2
BdKyXFdj9GoFhDJ7agT7tU2pXVBsvaGjbJHaxSWZGzSRKJ6de3KBaM1dK8JNWYPCzUuyAjtiBtkr
Nv2qLfyDhPG03PqlKqZ3/SVy7qJNVY2pny2I6t/0HbFUxckQZoNhYzA+5easEtUA22tuR13uEfKx
bk7oJD7KGiqDRKXeM/WPEJM2jLDVN5HsX3iXkCGsKWC3/dCs4/9KcKsSk7RPKimD71Fq4g7tk6+E
OBAH/Nfc2R8UGOO1b7FtIrMME1LerIBjcMNJhvuRUQMLysCU24lbd3Q+xBzRcsDeapJIkj3Jn0CO
hNl8ic/0F9nnHXF45glc7QfAImaypG94tM2twQC8x70r+QlZRJbqN2N3IaoQ+MwphbXpBb/XJt1N
55PMpRYqIiNzWiTGJ5/6WpjVRZoOi34gaPdqS50Mnx6BdCh2cZww2Ha6Ufurwx/5/Ze/nfbKIIhg
a+5gxVKCsEc+LzkGj8zESUQbZMEjsbAhliXBaI98biUzGTIsnOwKyspyRqDziFxPn0VaDc3z4tlp
MgmzYhANN7QRbfUBZ2jWLhlQlI6xZsBKyCBtnRddz+WqVT1bONB7oEv6IpweNHngb9tsu7QkFewz
Jt27DXgr5S4tFuCF6Vf5xMTOmKZDBzl4eAEl34B8jJjFEb4mKsauGHzxLIaCTjhxl5NKfxtNQ0YS
T4l3lzVVM0gwlzsjLgUHeFuW2/HSFo91NY2hGa913qvCGRszFQ1XtaZWWjqjVrfmrY1o5gflZVjx
xQvzt2Ds2K1SM8vj66axoao5zT6Jbdw6pBgtEx4abbTWIHFI8SPx0CIVAuN6gGyjNfSZv99co2uu
9RsYd0hNQaz4Yej0PgbgFoJcAC6uzsVHrYj7/fBGJ4ZveG9Q1l87S2cFflX0J4Ab+Ulcs25SVqUG
sMePRLfj+re4Wr/R+ojBR2W7pC/4yjzEP13sJs16Hd6ri/kRdROch91bpejoSxHrABDz5uRjUO9E
keKRrwlGZu81U8SqrUlBRkz/TUGiH5wg4i+4Q3HHeXIsw4KQPUVtqWhrTldrhfZ5EVSL80PMzBTr
RHz8+6syUm33b6Z51tkKc8U+3cZr51+lwWsYesZbNaoLuuPFD74uU6SBWNEXFzPOX4pPJVh7ukH2
7etzCZbWP1VH7FpWyQMha3QyDqO9W4cbOEASTz4YnB/x0X0bNRoySqL8lgICd7jQX2TvH8QbM6f9
otI4RbbaASryCkJ/Rz4chKunNECXiZ1PD3j84FHID3PCJTBnwkse5zenXYEKn0je4IofUNXwfFxU
9a41pO5OfzqF00SvOav/p4oao1sIOqgWyuisV10uGTyyjO6SlpnsmoWYiQ+lF336ZJ5ZIw4rLTOv
AyEtK1j9dPiP5qr5hB1f8VAgsHj60zeUsItt9Ysg52IZHra+BtNwLoY34SMo/C4GT/kV1bPjbe5n
aOLtwz5ilWlv7rIwmcurR4Ra2vh+DdOIM7knrP/4NIueJ4+P0GksR19GV1MzLCsi/n2Y+TvgQ1gc
fG+taZDIlT3dJlY4cLzqycvr7TUcnNwdFI8NxZWG5fF4a6Wh1cAqpQCYmPKAVn1gM6EKlMLI2Ged
I/OmAua8qt9lrdUXPkrgkSX0wwRDkhA48KW0RnpeKAd7TNgSfngJooIId32RPqruuEmBOemrJwoK
anEYc2Jki5tpv/5cgcCbWQ+u7LyJhnCNiDUUOYluzYe03ac0Pc8agniM0Uz/VYXORxqr+TFWGdT3
ZxqQnHpMMhja/MpBQMqBm0F20mbNZLJStzGhYcBn4sQEy64PBE1MIRr9YGGjKNeRqjXZhaBNWmJU
zDYYYngnQ7VWIMPjoEi3rlZrdtXvg6NHqNgifGXv1DSkeUswrJaQjdva031lyKAoGR498H/qASqy
JKUeXptyygrztdbwMOP5WsrfQTg5dM03UhKjjq2mnPP8Ij9BZUKu2MZPrj6NhN9hncu24jmAnXbY
jNFvnyMcZ+Bmpw0YLBLpkYJyPdZvC8r4VG0LQWKnUOB1hy0/Z2FwF0YSlzFRRPUdPxD7jBSkHhfF
jvXXGRVkpc+4XUtvnnjkDy/CZRv5CVf+9z1Q6fZpiz2/C7M9foMuelHt1W3K6hT/7RsgIoGxuwIt
S7XPvGqO4GVZN7bfJi9QqjOIJD6EXVREg/zJMb3fNL/MWg5lgtrfaeLmYRVEXwTDWrC39yYdIgSY
eaVZ1/g9b9pH13M2z0JqXA+8xPoDg4Qg3cy2mJ4n1Q4sgrL6Zc2gFVxozi17DsLhXxu1JMDtO+U0
NteISCSzxp9EuohJVPPRm0qBf8QK4ymuQQFlcurQCKaFNuzKgWel4tTuEBuYDpmHklyPdASUthYX
pr4vQ78leWkq3rTZQ0x8PaRAX2WqoQ1pc9KrQPgNjplY9UxeppHmamXpCZjj+h/soF8l0WMaoXZD
gPoiqpYS5ZxXcHLEm09a7RZoRY9wb7B+g9Dr2sXlHaZQHrD5vTK7cMPGDHbQQ/HNuEEeqDhr9uPt
EM8V1s7MLc3KLIts7WTrIK+wByZExUinC2lGeJz6OXOR/K/DGS/rR1XfuISnJzkf9nOfCg0N5E7t
94Uk7gqcSHu8CMFbehYU9r4qujvXBNnVSUoTSNeh4k7pAM8nuwQGE0LDq6QEcnTbsrA1dXoCVgFr
ShIdFOH5LOmG/YQXmSloqfuk2YXtAJhHMWlUX5Ae0pva9Mq8DrElnbma24nZYFU3WcSnlm6adtJi
bxW1hY4ynssAo3w3tRY2agJMED7hbdHDwitqnH9u3T18o1OpWQBGDDBRoJT5JxXnKyeBkIi1pCtw
jQDOiObKuNCjjDc5vUEGjoz1OJyNiWUYJChrUi3ej4Ncdayj+QfM53paNgOd39Sr1GUsMZF66yPZ
Isr4wLWH1AXK0SZcH3aw9KIXhn+8Q2pzMA9rQMnP5vFbkyoLsCbSpwfHBDtmXkNf3gO36WpggXqY
7oTzoX+R3Fdrlw3g4iDe+uPIDiU16xC+5oil1LGUzW6CI2BcRm25uHp6+6GUKZcAoOFZ6QpTKLLs
mkOmwRIzhOM/4GRVtyL/lmE8URpfN+lVqZsrCKecPkDVqHVUfHo+sao05YFScApLTavF9nhcUbCr
TqD7Bqee79Xg5QYviR9x/6mwTtz7JNhRafF71zf/tykU/gPq8ZMPLcU1Fn2cmZvE4Hckd1dFlcV4
Rnyvq7uPMg6TFjiP3XQ6+M7wC54taD/NIBP1y+urFrCBlQgCZzg+e91nJFYNHt8i4DWia7MBSqlq
KIeDUoZZaMq9PkmNh+eVFTjWppEhc5xayVi3yqe3dLa4Rrd7tXK3dT40KOkk5Ss2TLkujMbuLiqc
4IK4DCxVyQRDwJO7FrLnswVw/44YrktmlA9PGW+3Rmv4Co0N783bR47t1PPZhbI+hM3kLLqrtNux
Lisc/YQPr8qsJ+PyahP002tQaRc6nIGRoKlkz0utB5Hdkq8dzFGPbUe+4LDyFWWc/HWUyW8gEwpG
je/qUaIl5HsdvXAhIKcVPmCMT1Rt98l9P0TxUrwfrJeJiDm/S57NnJRG06v3zaMdhv3nxyf0H9yc
OovumPGp4hrqKCt245yk5ohjRNU/4GM6I2PkcOtjLCCnnpvqlu3t/XGpzSF+PtZ+UFOKCU3LieeD
BzV+nfxNpLNor8frmC8AyHTLezFDcY4TOv+AvtXisr48ZzXKSThfIBwo+O+0Iozw4bnVrkY3fcAY
dAMU5K676nGU1XNqRjMaP3NunMTer5B4CGAftEUtN/35pZi5LFNKEGDgHG7Cx/6ddF+eoG7xY7aU
IszkA3QcJrcORklzpb4DAJqGCZqeoR2Q4UNsZQefiBT29D0HVhAlHsFqXeCLelpiXBch5Gw3oCdI
mA+5bV1XSOGC9WICdHmkJcdHkFXOlmDwzUGRyBC78qFBFJ5z/TcrTReKawQl20uyQOe+q0mUZZRD
VLwNDqKffGZqG/YbDwnAFVrc1TgKNgkPGyXrEI8Xde/gA8IWZdmm584Hgvwi+k7Mc2s0XG9Cdk5X
+BtUyDxfpMuSoCrogBho0T2R447lMgcCI4T6GxSpa7SH3JB0MwNBr50KJJAK/jZS86xV71SuCDnv
RtP5kUFoM9cBWzQW29MgE8LT+qxKXn+6TgVc5Ve2mAlVrB5GkLoOcXzCaug54y2+3RA9Ql96dQcp
6/WPfVlvrCOo1BS28G1GrHsDc28VpYu9xf0sUK5a6s2ClkekCbPS3LndftR9BK5yWzt8jlx29/5E
jk8yla+B73AlV1wXdcvHaJTlHQGjzrzFvRGGY8VfriPm4BpBtIDuL/be+94HXzXv4Eh+4ooSzeop
AgvCea4dJA3SGRylPzvKz961yl5+JVAnKY1f8LgEAeTg3dYEI2W7pDm+dSxQ4fLUT180jpHJhIIP
tqUwzq3oafFZP6SejWYhwpJaM2ubtwU7kR0LteLTI36AnUWq6zy3OA23clzUHTPTTuevDN1tSP6K
EMfUZpxxTM9QZog99ni/f16XBk36v3in2caHSe+o3YT/5ZfN56rl17pjjrPaPVw0E4rud4Iqk4vF
sD2jBIZZpJk74XK3mC4qB5oXCPExwRANka1ApaRfg83+HCy1ww6MbyZLGdoTIKFXJ01ke2MslP1S
hGKHwnvXinQo+7buM5O9hrXzmgGsGsd6ck0CKhOT3Zp9avRe7/faI7Uyzni9WA5kFJlkhegRQymL
UyHE2QQTWg+cK1wnErTF5CCNy0FT4TDc0c3JnnXmYHnhMtim5olJP9XNv/ZYtGozLmVONPP2Bwen
vBy3uaIghgOzR9zCLGw1HXS1MJDpXuxFw1d0wD5JMPZui1Cup5iqWoqL7fOOTy8yY+8crHALhV0b
m85uVhlccZ3ZT27Gs7bRhNaWK+fEzyI7Bkaxe71gSndZDGvjlbSKP9fxs1fjtT+46I96yPwKW4GQ
ybTYMVgN/aL1a+K/nR2ftZnHtYOtIjjzLbcdrX8RpSwa7FlmcAcEKpxVm8bxqoII504QY4oU+iQV
v+nFYuK3HOGRl7ytHCmtUGwtYoNuArwy8LdYMQtcGQnbvTJgkbsibu4/X7Wxbcd6aDiB/0gluThK
PuHoXSTwK/n5p1kvaI+ozTxjRsTspdqTEJs5pJDAvUvK2Rw+Fp5oRZNQJHfuVthlf6hD+HWbvev3
FhlAOaMTCBmxm2+QL+zIeRqdBbyEjus5inOXMVCYyTD0En1TQr+nABjwH7Hz9OSizMVpa/r0v2KK
gQ9U13C/4SXIZP3+Mz4/M7Mf+KFFiR8GLdLSm32Bf8l+xhafa4moiftlBiIEo4KZuMV91cbzY/n8
bZ1WPaUOPtvs4Sjj2WmBbPsae7oqiRZzw3dLuNqfKiX5TYifGJEHsth9KS0z5+QtZ0YypEEzTY05
5KcoT2osq2Drdpjz1punCwy2OEkYxf/6viKdE3obzcXaj+Hg2jU+Sv/JJP09dXlZQ/DSB2OzcaRi
8cGtqf+hpHmvsF985KoZ/PvTDgjgY550ftJoXevlL4vJd91jLBkIIP7Lv0iQwHyvTl/ADFIsEYIg
yVbHQ6V7LIhtWd3owkdNKk6yisd7UvKRXxZFdm8tUXLgjzmRr60q08sX4eC7Yfx0fygQ2dUFVcHP
QHcMlmyUcZ4vt3lseu8mqrKQ0nHzd5u/tOaUm9lMyTWDWIzYjDJHsNkdhEr1dWnYNi/jHuvPJGr+
HI1RMbBMHRO7VqJzO00vrxdyRDOmtbUOxtZtuXXBnf/oiYWiHnKJ6qX+Q3yYtUG6FYpTebnsNN3D
0nmubD74V6H9jN9Vt+3I7VtCBn/++HHaX9WIZWaO65kNwE1Nyx57y0OW4oWGXyORtugl8Ulw1WUh
lt9bZRCiJvQrJB+v5rWDS3QqsvMSDyoiRfP8W708siO4pvI+FCoVfJi8xq9cD2BVQZMEhs38qwh+
kYx2bJYO9GC4a523MnRs7VepnO5H0czf0394pWKC/GPHXtzRxc+l6IbzwR/wCrCTaVyCA/5Celvu
qsQHttnLeYY+LkcHIR9+I3S+C8dnUhrAVxdr6LHzrdXoIYx7SUpp9S5O8OhWqBNNCaB5vuRxovSn
w0futAKYqktgJLWbW+QuHWledQOKWDGHn8JVL0zpGjCoPA2jo5o2qjPtdt0b8+aj/7SXiWAQqEIC
E7z07VOa7NTuGNjM7C5DzImQLw/p0oo4Yhfu2fuMtiEkI7anzXzWMBO8nhqBAoZxeOnMV/ZECeAr
G3H4l/qX2Zp7Ekl+b5TewNjZkUsodkQz3438xPG6EBIrZCLwc/3g31Rbzekm7Pxj7qaS+E1phFx6
NBHocGjIx8T6lcHXMlF7oEYpVEUoE5mhnzC9lm7p/xCtM31EnNnO/hYXgT1/2QajrmwdAWEdtPch
a1WtKQ4hMOp8qmA/JOiMgHKxGawqrZ4wmLIsJSFZzhbkWjI9so/OV5Z/fr8us9D6hVBjh0GY4oLG
ojj9LOgYA/kkaIDWibyIRaH3muCWN1FiIDCcrfmKszwXS4dIO1AZGVch7XfXwAlcqUk3sN18sB7L
bI+RdFxTwuiaksztg5Oanbv6HVZDQ+UnSgEZk21bA5hxJkZR9/TSni3NxZUw1bZd8rqCe5NbRH5c
6NiMkNlTBBXg+yay/hlsuq5VEuUDEyDsJvU66c+hsO1lXycRECxfjGvAYx0nDR3McbNYqH2Daton
LfCUTKv1sk0GwfAHyeM/F+czlgvSxz3LEZMx8eVdxxB/xhHvDiHZYBbyiJCb7wxSpmZXDycZoHRG
4CHwN+mIw/NHI9UaAdHejzH+9PnHJ/7jSctUsfwvRQ+UlKBmrLWvgt+B+OVwhveKI2wvygwJbkUp
IdCNo0g6S46UX0BEofKizto/wBvFwRF+6wkoLTw9Ic33YgNPGYU/tfliyvZgYxpUzAmxM5QJ59rx
hOcrKTJaYK5u/t04ns57x1byLPQYOqX/IXrVX/TbX9K3wXW0bD3q4Q/KMJ+pCG+mcogODDIoKhgY
3lJyOE1a9f317A3pEoG7jfRDDL6uuA28xIhro1iZo6Q5to3SNt3KP7mtTh9VVOIs7xOZSRHigfQj
PWu63eH2x/9ch0sS/9f95KH06/DbbEkEIdKlJ9sfpdU8O9QkVrV35U11LLl2Bd3p7ABipQyg/jQf
/kZgZWIc8bpYNKlbJC3+iiNasCBjxfsItztKl3nI0FsliXWn02MWRNhW1wvhIyRCIMEqpY3Jxn/n
WKO/spjxN5XVjz7LpZImhhjCLwgRg/Lkim2W23zQMz/oqdrFifR5qiafgPU5oW9q4yksAhGfzasB
X1KFqkIdiWadPk2tGEewLL3Txt0jjoeuFcqpvcKBAyUlJM/guIGcw2hOWW2OmdX7tu8YwlPx7LoR
BvovUxCtNLiQpv37jm2p8ko87vFEIHtna+cDMfW4lysUQLpbMNwUKUKJwvfkx+QLjYKvWmozjbqL
SkRUkpx+T3nZwI3ejzwkH7k2YKBvZV7SvJx6e0VYHXYZQl2ChLpwq4MfbmXWtJkl3SeExA92ItoZ
gnmqD82JLQRsIH/dBIF3xp8fy86QYz5j/D425pedMV3z35zkBb2XHVTyvugamKtnfz7ug4XS6eRX
NOLci7PcPk0glGrCr9r+dUnLt7s4NTMRMEkkeonB3MB5WBhCsUjqFtqm1XyPQbdxyWWhvVmIBfxH
GNtfXjGa9lQZzzpqRT4VHW4VHmq0l1oFAhw2scBvGZ0S2jdPMUb9mF6fYOzhjrZFR+0bxMHCt/J6
ITt5DZEWywKYb+Rc82veo4/k8tlSENtQaYM4nJIMTsGHE4ZmN9G11kMpGMJ1TDPObKCjXClUfWAF
Wfs7OIwT3uKq7eat7MNUcDiN+NpwtTcYMeCiP/id6sqWeWGpnRsh/B1EZCpmjwwbGco71G4dZgp1
aFJN+/59Nk0iN4YZ9UxcGpZuCXEI3OLYtkAC4+juPVEdm/27l5F24PsDsNCVksUymapEsPbwlgxR
04CM3jbv4L+xdNJ5dh6vqKJaAuEY7C/pHuXCAyU/vgkX9Yl03tMcrR/4D4lC0UM35XVPV8O0NK8+
Wcd06GGLSWGQs+I302DRyoFdMmU7Lfm7gIws6WfYgStg70umRnnW1hKKddy4BXixDksdfnc8Nkdv
NvB1vBEGQeRRlmERWgJ3t22dtOUh1VgVwKEs/dVL1kNM5nSB4O10v4E8NUX3wUkjkE7o6Yl2ort+
cEf8ucVrTL7i9hg0lz0bHHPswu+L40z1fKuJTFBX5S9EmNB+aCGejh5G2kYg3EhhdFzy2OPHrIjD
GS5j5G4AvXkwOnlJxm5RX8lxV6at1J2t+zy+Nd8SMXQRyd4fIVuwOfALlXY1eWbDZre8+Rl74lcf
OV0oWfpw7MPWuj/gPlRxWRVaZ7bEU7LIBSi42Wx1baDZQGFxnohBYhRdzVgZ2YbPbRZ8G/kszGxB
OtyNyHwcej91IvcLPCqTt0n0Mob2vaZTZ13Vd3yCyii0JZmQQMNdxukwdylIZiP2c656U65C4mBn
V3nUEBSvK5Qzmtfx87NGAC/r2G8ssWguJXhGyi00VWEuXWdh0pJkMtBCnsj0yn8/wcEsdoepedwV
gTfT1PKSOZVreLlRKC72+rJw3bqKooShOn0L1jN/VSp/jlFEaUzgU4hspNxvsGq1bBg6nKffXwX5
tUCQsAJRgbGOGlWDRo2KTXjtpJx3FclVk0YFGnU8pNvMcdVWFn7uEPYvuJpLN7Sd85IsZj3E6YW0
lk0Z1u3GnjRZ21xqjDgVcPKu86x3tfaA0GnWsKtIlLC5rv/TCwGr+YzEjZ7cK5aQnLVXHWQJaiyG
NY4rT1ND+djz6gvruDPwuLlohfYoyLqGdjrD3KHNrhLujHEu5MAzhDGTMS6ZKyf5NcNcZXwFG/dE
De0MfTlqRTo3Gkk58c50BjlSTNtkNZB9dyAzlpnjH3Kc7864CJeVuuBiTMA28AQOCit25gIGtqEt
xOGoaJdKsebSb+8PEko/Fg3cggZLjt3QjEfmRe6OT6h05F0viqi2eB4CQ2H2LgDLPj5cYeG6+845
xAevIooKUB1VThc+fekLyRlt34WFPqZ2abkUdh9lnqEB/gSUitrJf3pQdpr7MHxFUxKKS1htXeC/
ZQMqwB7siCVMKAIyGf6xhEr/6szFtJP9hPfZW1pBReXrcqzgu99ABcipgT2aBXoVeFp4yYFkPtIH
g3tjqZaNy7KcwEP2w3x1OgmlU1c4QEIn3cuTNGseDrRvnKna7mYtJjGTIntwYcG1+eq7tqWAhafW
aKQwR/kbDJrRx2jXO3fpTm0nR1qUq02doSe+/RTRlJuO8D6RtyJKPMILNCp5p5Oq0MWIV9wl8mNV
5ZHilkEPptp8sOsR7pK1Uiinq0bV+0tMASsMN3NnVUGfiQI+diNf6DDseIBaWFJ5cckezjzYYf2M
hrBgTsi0PDh7bUAO6V9+TkT6afEXrlmNquLgGo7iB11ctL30NlLAyb6LkUKko+e2YOI6vrZtRctk
FvnQZH7HlPB5akc8IYI2++960axDh3sok3Pm3pw1maVjYmXcjmPodcUDXIeCPnlWzSoSxc0Nh9yD
I5DZkqiVl9sTLdXjPWharUX+xzHMtSPzDWOR0Fqqa6yHO51RAhnDSYTblQ2dJcAWxOn+Z2I7pLOU
LJX61HRW6g3JYeFv/BbEjo+Wv5RoTiox6+8GAnXibFo+Xcdmo5pll3KXPRirX4NNKZFqx4T/Phma
4h6qp+y0UivjFMpOrTX9iQM4ex/RP26oRcuGMlml3lN5u1bwZUmYjz42hWIgqwEhjC6dINWto9b9
ios7WHgmzlrUSvQem3oKA7XHTW2jx9hoBDxeVvY2jxz7gzm/pE87xclSujS+eeCLgNw7sYxtXOBW
FnDI1zA+f9GXjLRh7peMlzvQJOANqXlKq48ghGT0Jqu4GvlncDZlkVXYbgGWjAevwg/EL60oYUTS
9/8wOW9B547za8mJg186qoq6rsIeOdnZPWHSgoxcEcRVC6rXc7MtD3SyzF/I6uzr5h8WnOVOGEo3
n+JCZmse0uxScCM0kFypSzFpNp2jBI8ptRoiKEmmfbF6jXkzhMyMLFjQfUNfZfjjgrYurahiAlV6
7QwsxpKlKya/ZAxIuKj3YjmiiBLJ3Jm75JxGpgEaks/inNbsOhLT80SdbI3ZSik/Bv6WOoz5q7mM
kVjaYHDN6eglbPJB1EsP0C5dRJLUe20izOkskk5mIGtPpfF+cRj4F1TGwGv2jN22sva3WATnS3eH
l/s3IWd1BIga0UGuIXAGXbLACxPfGsyFeR+X1yDWhkHHTcmAA+HKzp77v6OdqCp2PfN5nHLRm9LD
fyRW172bCfSfwTxshkytHCJ+FOYcmvGmMq4KflS9FLNCqr6y5kHaTetvrxFMaE8UdWUznmjLFfEn
FZSXLMy9jf0yQLo6xSwOF5+1UtjhNp8YtuIfbaiPvfyr8FvFuZXRQRlnwqiKnD0RgFefgR14F/J7
9DYGYo057kg4xffiJ4avNcJjaLt52Uvu8aB41KoDAkCiQAD/E7kzyrKp2Ybrx46+HDmKTl5hdrOK
HiIpeYu7jXgZTT7wEt+N2emYdhDkMctlzG8UQ2hQocW6oeuwzbYHihCRsuUI0vbn5WuMT1tOeHx6
DhHMZLK6ZYejnVJKGYGhj8Tj44tg/g1mWp9PYnQN7siKX3XpW5ZzMxPOm8YYAr9FNd4kXLYTU8Ag
RgtkdDo8vUeNT5ONR0GEIyePZHJaZjuM4qYhMne2MKOIORHw7456xxFUHR0VUGRCfa7l6Bngmtvv
PwvSFAHOUQW6x+3ofzaiE5RJXPk0uG5LIHL59aapXE8kYQCllFsirEGsR6kW4sww4qX2CJopjeET
mE8+aoUdrUHEWSQB+MFTmqTRXFyMZzqUk5gszTrIp5QhRPYUn6SKw53jt14mLIu1+I7WjpSzepDO
PkrbQQUzzhyCbNoUGVdQHL8zw90NHSgYXMIMEkZOk0aXyKsa7fGMkg3gwawPVAwnaCD2x/5sVsb7
jKuWg8nM/FRxA+EJlHNQ9IJovl4SNxg+oQaQgaV1pV0HKHGalZE5iLCmNiPZ+ku2r1IY+xhoqAIR
e65gakNgBlQ4GbeA9l/2KmQ8twrLX4DbjbWZ8bP1P76oXHeXTt15xrgoE9Qk0aj3FDCb5VeHqOov
kXSqvZy9a/R0Pz6+B4hjLUA3/RVQaUgx3q2wb7h1muFaAA23dkmgW1gAL5cx18gdQvNG4UDL4dG7
0qgCvgLq+ewduaEIDI4iylbQ2+X595Z9uz2XHwWSKDCX1hvui8K8hFvkbNvDLmFVyAwuBz387VRU
c8HcEW1LTCGUlEjxgDoQNZ3XxuoCAEbnbBroeARJhcyKHzsQ4GhdCFdevSij6KIwloA3KeF3jeRA
90T+GoyWPcwcVra72GTFRUv2PptyHBLaKFZ0oCYiuIQawpwYmdYQPT/iK5E9rXqMzoZS68rr9PNW
JoLmiPEknEDmID6LfQBcHK5thzn1y7QYxP/W0SS/SBzRGR7T2Ezu9h7xbiB3aQBdOdBt2dGWRK3o
qzs9NFVwJKx8WAV/Jiza2e1G0wWSonDTu1M6QQiO4PJIAF2W/t6D0H5vZdv09/dSWu1mD3AMRlBh
8X9GcwG6VjK4ijpRvDtU8bD1G89x5d4zzyIKLYRUR8Dk9UEFJm5fEFM7ZXqZ0hmT8MrUsrGGG+3Z
WSp+H0LcuOUQ1JhSViqJJ+yQzSLr1GJ8tdVqPgoSsftf4BElQ0fRZDPzkUbOxTa5qvey5eOIcYaU
XVxxXaEDZ3rbLmNe2/8fTgAawK51p6o81YRX29hgQAVWA4DSUXnS+F6lkkcKQoNn1v6z2Ega3mZL
Gosedq+MeEobTLn7pOC9VaIf/lxgCcJ9/fslv1n6o12laIeLqU+YsCfEczam9Qaug+YCS89fsAfG
zbOS4VJ9thIiUjhL5jok3vLHDokMRZpU0o95UAkmRG0/W7aKp2Lrj1rhm7aQ0pHDiKG2p29AUct7
dl9apfqnrs75biSN++Ug6vHVNvWKXs4Fm+7QoOrxqII79Lj2d18YyXOkAeQwXNQaBICJSlurYggH
AV9d1fHTdqcZ7M5h+TyM0hqd0I71/p9CY28CbvPHLfJkXgg6WvfIbYOY6+Anfh2rMqCJUWcMWWPx
NiQR3BLELWswO/hwr80ysVTRCP5F0ovJhaawKQ0CNEKkUwf/s3fRtIMBidk2wubViCsUUUIZiAij
aW6FlsDKxSpvBDVvrEagN1bLbc3k5D3uE9Jf+MBbErdITzSq3yfc7Hq+p2aX2n+94A2QYFI/XDNB
Iir8yJM98SwHJNWLgBWysk51/oQzhepBex0M1MQ6NH885JDiqDSMdxgKr/WkjKuZh+u3K1Dzipad
Zmu3Ud5xgqrkz0Rlg06GcR3b6gCaPUacyGIwr2/38k5Jr3d18ZX1vLsrZWq8iZpTjV1K4tys0s6a
xXtibzItNdV3D/TRHt+DXqSL+/58Qdh5ZuiAPiAKfDiLqL9sNJziEGZ4PaaXRhV1FhgpbD7SYGwP
t0E2ICcGFzLqaG/5ADt6jbUKfbfXoQVjTBImNfYE5tlN1XK/qjcOmVWLI2lhfd8ArIs5QGfudFzR
yKrsEaz35MKzG+0+p0l4ojk8d6j6wSoki6MUUhE0waNV5dsuSr5OTwr8bWDapODT6Hlqh/j5RgAk
azDgz7hDp9Ifg2YlX8/Nve+eRtj68wTo6ETjUM/P6Fum6Fku/LnmajAt88Vbh84VoED6f0pmn8Tt
r4aJyHPfqfexH0NkeMyx+SdW2D0s/AhpVQCq2noNIWjYy9HD7lhtchD9EGoY7ugSCBui2YQ21Sv2
1tzzQfQ+4H6imnh3bbGFFbT7gN4E7/ESljT0oVrVLppnLWm5xSXvQdP86HuL0+s0091Ftfme1tNl
B/yYG10jxoeRJI9FfpWwW9eqFoQhxkXMkjBGjrm60hbCVrlfEO3D7InNW8GPGgGKhnK5izZOlRYd
xyEW3SYnHVTBlgOHMG9oh35QBd69VGJz/FhY8YOfTypkCur9H0wlZhumKvnQV8zgXlLQbPPDGmve
21GW/4Bh8hof1tnc+NCy2+03683IFGXgao30jq3l268Nr6+tI6Mge9Uwz0lyCb2uJAZeakCkhKYp
lEGPrY7upwnSyXaA8TMjRTPeSWVJMbGMrdvSMW/3zK4AL5GIm36CggElhZxIgVEnmdnoJVVkmiOv
TcBmabdGUcyb6LEbtZ9sUIIwrgm/aix4txg0LN6TYVJ+TPv4C0f1JPjlrjvpK423NvzUysCfR6BQ
hTSktnaMEy+htIW1El5VPswchSbmymLE/6gLLrOvDt6sb2WkszJFVNLlHBfIUcxU5sIGuHfMMZDi
5AjJIUvXn30vGxcDswWLi/iG2WpGeLaoGH98fLaK1lmf//cc2mjp4LzYGdGPamcHRX4g76a0zZc1
cTYI2UBGe3vbuxqG8lDbVoqGIb2FvGDrl0yLUjEUMECZcoxXAo5pWqrJowPNfV0LXJOHi3mtSvYZ
n23cp7BdVoQfanNZBh0ss8sgm9pwUbQ6L4RHjn2r3iAL4yVbguzbcGW9Fhu9mY6RWKBsWzHDEijP
bnt7sT6xNnwtZW6ea5lP3ceYkx1ntJUJnN3f6fTvcXPXWfa/r0in/yH6LB6sjm+3zGRWILB8X6/B
0GNb84IuzE8AAPDfeIWhpxWuQw0mb5XzBYW1UxSkdxwoEEdUfY++iKsoFePLHTGIT0zyOyph0ORd
gOXhpssfGbfkg6uSXN12xmP73ttxN82QZHkpXY2mlQDhwuTdfyWqOjZmM2t8pprARX4NCyQ3GDsC
FyNdEMUZnCAkqu78tcrQ11KGXkaThgjiNAB76h8XOfhvUmMTsENjVBrKANJuO9xHOVe7Cqivs0fy
lPPbXedl1hdcDtixY9a07ZE0vd0d1ji7N6koFV7sJQ2EnPeUFxGOr+DNUDETwvPhJ0dk+E2cK8Uz
OOHD+XOTpWPfG+tPdvKrRf8Zvj8iBgMe1pANQ9lFQ74w/bIYTp5jkmFQVNHDyshLH+cDNjHHhcDR
mrIQNrx8sOW/a5bBxUWBHNgmDVzoesgss+oXzNpePTs4xUe3P6473zuzoQOztp3PGiIEIPRs8cxj
rf7oIefF76Io3u8Psfpnxmqvy6Xi/8plt1ef24wMbj6OcBtai6XWLDhsErEkGsZPahYdJxn1UlAB
UToVOmG0+aHiGNY4LhBmvwKwBt4r2t+642xXByospDJeAXKwPPPm2ndEMLb/fQZGFr6jngeevsgQ
P4hfdUlB0S/U1+/hWH/zPelQ2muzC84aJHiGVYHjLc9K+IlgzYsg12OjQ+L0UO1KCk3muP6uGpZu
aaoDBPOPyFwYmWDpqT/pqqvE1J73HE8R2gJEhqQWE74kPb0cupnCJdXJDiAAAhb79AA+R7yz8WoF
9rGHkKCK6q2ki5uQi7aOKoCvmufXFPnCqWIInTEmMtL1QXgHJdckZqWLZeT3Kl98VZs1pBL/3yc+
ZFWKF/nq0prNlPKZeLTCts2axMTcpnyBfNb6Xn7VyUz+U0wIa5AOAwsHdU737u+cEybQepq37c9m
UWdhmJU8kQaJ+EpZCdaVK+LObNUkT/uj+NNGH436R36SI/D/xyuStASM84xb/XALwX15fJySlclI
tNZFWL65rIO0ZYpOWmQc6fmNtae7yuhh4NzH2YszoRd7FywyWmmxGmcnpy8/Z3LQmZr48KLlsu3b
q7fTB3vt6ErBEi24IooS5DgfUkHZB4TmkHsIEt/yBPQTuS7DUaFooDBR5zBJxTpvltU0lpeJosqL
lPJKgxCdK3CRzJQlrYwMDbcrPYEKkL8yMgFu3TR+ho4hZ2pBOMoejB8EuVE8f5VZfkYItwZGiijL
qwZWnZb8y6TrDpPNgl5yf2E3384OmmVYXEHAJeQPV3EtxlVm3CbcsIsD7DRJULJKCY2LTlRCqOxT
l/FdIrEWqj0gaP+/G+Tn/h1fpvIFIZoEcLIZVI713Y1zCfxHb8Gfec7PjvikAtIiHC7WNeI2Vm/b
F7AF+Sy/o9nQr97Ri1dzBaL2+OeG8a5bKYX9MFTAol0/ZbBGY7tH8RNDj2XHma/bGbHkWLo0odjX
HYxzpxZkTu2WMyT9ZBjClmCtWOZzJ+mb/xPRN1wXOK9OMA7qQDg6LZ4kuuF3ihFam4Ac11S/P2lv
wDMmwZi7nhdmnxkVEeemvWg6G11b7rzzdGbUl5HglWSN0+giXx2uTbdNveSJF1dzhufkL5a4IYxb
L+YZ0B4wYthu/6MYEVy9T7uy30xNBqyNu418dp+E0NwHHMRthqWx2ezm9BF3kTlfO3D8IH61Mgvf
Ca7Z0zWmIecOLYWPfLYjv59k3SpGf/WIQ6cd5l3fXaZPe20X1rZ9/sjenSCsDP7dSeQnKq3/dIEj
u8fdzJEA+lUcqGHves5Fzilvb+jD0zXxZ/gDwj6llIUr0isfX+3VDa0xkU1Da15+cknky2+rMzOp
F1Qb6RwEucjzYq2bNfkGjsMXdahJQ2vpUvvxny3L2jX7JheqVJMxT6gBnt60RJ2kZwny7YzrTjVV
8H3uI9nZ/fTroJUvj5GMeAz6K4/S3+1VyOfgblRLvxabNxkDYJ83YFGBg4py71jjq7nciDEgCygl
G4dA33pGdoBsnb9gbRMMCdvtlST9DgjQLSUlkEg4nUAerQfro2H9OrVzSrzluI4MaxCWumjPLJWg
+iWU4VFF/mlq3/nUnPUjJ1YPJHhVV+7+KkTro1EVOpHgfzr064JwmTFT0F9gvO4x3CCQv/Ubg+m/
IbbB5X2Ua0hPODcM+rU9CF5uMtTkMvdZh1xE/KsDcSFfIxFIX5yEij+0rJ/U26uU6Zkh5i/WaPkU
XVsw2orFhMRq9hi6LZ+/GoIOOLjjaolYAIaYyPv7uGND6uV0slbFTI5cIZu6M39mQQ9fy1XJOh5t
XTJJF3ahm8pYHtAztsGWv8U/WENV2WdCMUS9o4nW7npyypBgRNGWGerQeN2NbDd7YX9uvmfxC9HM
St0aKFMH7gnL6KAp6a7sqzAKjqsR6y4FTFeNJXNHJRQ4sxo1FzysmtpDyD9v8SJRzEL1ld93tpj3
i6eFH4JI2+MKxiUO0xEM5TyGsqmF4S5f/6RnaFpG3BH4U0dBt7hqAAXstQTE5lCfCnr2M7DkgLlM
OV+5zdDbCb8Tj5jAZW2Okd6cZC0iWYuf8f+s9qA92zTH4Rk6/1JY2QM8rcurgsQ+0Tnf/qxlDrt/
z1FKBjnoWwIEKYbVblGM0OqP1dsMedgeCGDM2T5fu3rholOsOMTv8YA07HmwxIItIf/RJSkV7oLk
3BHFw9QQzdUvm3fHiNsj3iN1N5+0u4eRKyeTCyfG03NFxyDHsf63WbjNN1DSvbibACfFMkF8kFUZ
B6vzRwg/E9dMs6g6WNTJfH1PLrsFKDlKzMMkV3s2Um4+0RjP5JcUN6WGcIRGxdXXCI7M0zZYh0tU
tG9GgIItlfOqrQ/VR2cAKBjCXHI4kd2GxJcZJ5TC62flrDmFP85upq7yFqlqKCiZu98wjzLLGcNn
wxINuTCr0YzBvskifLlj3B71zDpI+VEyI65GWR+kLTHYgtF+ZWfMjU+NsI9JSfyNqAnyZGHMF1TV
V7bjq6DPGXZikr1zr9J54cFLCqlhDuXQTVCqfug8aM5EOwdieYXMIq+NHbXzm7McMvAfDWMVwgO6
yLwiacIzPWwHkWwlS07Xh/XPCwLhiEA41M69P1hdwmVZRyLawXtOkRGNmCl2L8yvlItb+lvr4nv0
QQEz33u0moeg+kX3bFwHfe5mVGi/ezcdsEjZ5Xo+Jv1TKC27m+g2kmef03YkRZIp4eRZc/NRJDhQ
6MM2j+VcvIH3rZ/IfIEi4bdRL7/VEvcdb6gFQYXhfa7hAidLuFuVfmwKmB+6MViSLnw280J4N7d8
968CLWAhqExljIowzQjYUsUgXtLaypDVWfAefq1E2Dkpy7k8w+Ze3R3lfDvSGc5597Ug3jqSRgi6
Jnk3eKU/BIFL//dnO1wK22GLsW0j8rBnBSfL3ok4vPLElNp1kZhrLQazUZK3/VAVj6mJpkmfTK+F
OqYc3M2NsjgO3NVMur3IhNYeF8JOpNqRrk5hhQxoqMZEJmRIsCWbmhydgLeD/Jfn+wK2asNJq741
kn+423+4jeqclg/aYKFaqP3ehx+XZY7SLZg5AybzDRKabTtzAyll9LEjKeuEP6a3YQHLfPVJB/n9
/EjTqYAXbNnfq1dGvsCMa9pCV6t/ZllElXEemBvJQJlbRymeGL/svoC9hLHs4lQ1UIOuIa55Ux+d
bNy7vQyQ3EleLT5dIsKLSoARQ3oXMJna0At5JNUyQ40yP1kZkKk+TdEI2lUElpjh81VAoUhurgnj
LU35SNbusUnTXVeMPdFSJvpKFPDt2HqMlAHMQDwWTPdQy531HvvIIe2J9MROk8XywOuqx4BqwTdv
HiELzwBp/VGUPTmhuX/DA5o+bwVY8Rp0B1nInIvp6vV1/FxHMA/SmRaEN9OwwcdLoNWyVBSATKQA
anTSsAkiSrARsd6E4yoPynXROYKOyK45XIjTVtBeu94AmmoFUnzPwvuroRp6aLYWN1VrboCgQTUq
me6FCA57yUIHC4bXR/eM86iy+elWnsel8hYoABXWqBYyxoLuMZCq+7y/Hk2Za4QRH/OXRQtmNqWT
or7cYF4FKvWD+DRPdt5wP1NJATl+iHyWe/v9n78PWYoP2IXT4g7DM152riqD/xbxlINOJz5bZGCX
dgUr9DZ9bvbAv0IxQihgeOpzRRd8sGvcmhe5PxtqVF0SPmPjBMn4G13X3srNhwJlhD5JJL83e8x6
s0WVIQJRFd9/PK/6zrW1bGktKs2ccu7tLpUn6UmxHdjcRpDZkJx4C7e+LRP335Tiks7gyQ5OhyA0
VA3kPo+dy40DXJEPgza4UI9tZDYih3+6EMTVPBFnDCLgFB9egbiBay1kXNEslyjDiq5JZFWLqfU/
bky+KNdydkyUF6Sba/sL4PJFY2th1SGME1vsHzPa4BZPrm++Iq2lX+pNKZQlmKNQl5xxZAszOKzI
upC4AeBzyvbW6rZIBdt+KBbinfgYgciCzTR0AtxjpRavLeDVRJXPYSiM2525VcB6TnbP9Vn+6DCf
LAwmdIEYAtU3A9jYihi3k27E+rXL0YjgHb/bm+W4vzhLtfHFqiB9nPXKKVn5GgR6k3l2qoIjLIWs
RGumQg2In6mm5pUgxAriuDXWlvPKxaokOQAdnqdyqGQ5oPA0GCQnLPOAEQduuoLGdJCdSlTqpFDs
G8eQsbfYJKcIkoPgzq9ukR+jP9B+YSiKltjNWJDzmLnE6Yde7zSUfrQ/L549Z9a90yM+CoFDTRL2
X0aeZOXlDjOiT/lAqRcpLv5iTxS6xTqYQYJtuyIaB48TWSgw/7+/W7BbbXL7iP/a3AZ7dnkQagQS
ozNlV822Voyly9FWR9kMiX1OJG2p4BU+RdlAFLWr4n41qFMR7t3ON93lG834laPVXdmu5NLbuJNr
iBDCEjyiHeWlXbwY7hy5bR/7aQPRbmi3dKcy49U9xIMJa9AgxyhA0L7uTTrMhjYM1JDX0OTYgRpu
iMzuzRPgHFD3ybRYmukvtLYMUIXUvyfYPSCdH93e/VJZ/QE5pHEJlEdyxy2N1k33/hJptfKIxTvC
Jc+cek/ZHEXlWBktwNGR/78ZbJa9JDJL3bQiafoLTnTnaHEjdjAzUrXe1ifgUOn/oQywtZKQqxmr
Id/xwNXfqw3U278XRQJ6fEIt0mtVwEkpZWTROlI7B16m3YLFf0z9/r91cxd6UNPjs1+7cgNTv/z+
tyxtaqqQYQgbatg5a/svue3BlG7IOlDzy9WuCPi7mAKY4NJzRWHxD15cV76eIA4Kl8gExxW6oybs
MGA2KPTlp2nP1XnsdG9NE23j7miFrjCyma5iRdqRB77fz5otjSDU5Q9IXI8795SWdYRX4EIzeq9I
ubfYQXsgH33luETAFH7MByTSPIRd7tB6pjlTmis21v4osDwcFqDlbJq4txvAXEXMZJHs720hQhkn
1EqeiqI0JHG5IdmxUx0K1p0tiymWsXUiFYkMVpSKaMar3HonWnlEYl297rERFIRhzP9En+4S4Q9B
HmypdfjTobBSjcUeGG6eEw8DrjYBQgmyIA3+W7icSL2i3ZHgY7X8NeNWBh8mn8bupuSOzDzkT9xV
MWenq10+nPO2FSm82v9LAnwjAa5H7pvROkyrqPNdS/zyuqZ2jwE7B42cdnPMfydVD//lsJ1Yf2v3
Y+Ol8kCEd7tqnEozIem5jdVcAvsB6iFqtNPFbQJ0mVgXC7sSj1Od6Wlsv0tl2b1J8bOKcHhUxfgr
dEYdclIqNELNLMvn/f6niWAgqllZse9VgfMxzm4se8RGkj42eOhWKJPsDgC9ApFVc0lZux6YByTD
6+t/3xOhtsF726u62b//WzQKgxIO5/kJTlnTUg6dzQwgDyxhhRmJwaXg5icdZc8OCAtqxlgevqX7
4dmEafMOQYz1iJLPBbd1VAziTRkodCJ/kQ+MS5XsgRVYErq/VzdPhunRtQwF2Udnc+81XkuNMHEB
Pb4yhXok/cOskE2tTiHm9DihsntayBMAkVdgAIv7AQF9SxgjXmjT8ANUjvQxjtaSL7tXCu++xn5/
kNREBEcOAPiUvT/fZhJQHRPUu8TlB7+qlDGw04/wQeJKXDuvzVle8qw6EnydAHZ5UuCiG0Mo5qkx
LYUKDoEQn4/I9Ni1mucinTCwKGY/TN+wO6UY8LYpGrqlMdKiPErKzQBx9nyoO/2IYq606mpAhrcp
gvliso+jbHjh2hm2iqfYhVDpstU3ajMdB/JOVDiO2049OvkRzp/nzElA+hX8YaDmUw5PismDMjOh
yyTCbR1bx9fN0mlOLiaqztxjBRLz0Lne4WUeI1S6eer52BGmhYib6WTxOKgcQFkYXYRB7ypBRrwz
iGb+By8Vz6dgIzpdWsdFCu7nCi02wLPhnDmKf9izUYBiKg6IFCxd8HenyNGNfJrkpVQuxLmps9KK
rVBcfG1m1JuJojvsScnJnpHit/M0g4MTH7IdNU4K3kFWJzbMkEsWYSF2eY+QCk9nqL4xXGzE1qP5
8lq/8sIlp9DV9ou+vC9bRH+AJMolBj3g6tDMqD2wa9MLDbWbSAO38Xm83E3cAbC4Qf6NcQM2Fm2D
D41bHLYIqpWMc+js1H1BwYmfufxcepfC95Q7Z/GhfflA6XDAeioR46aM/axwCcNt7xL9o6ibfuQY
lR8rP3blkEQ4q4G457uQJfbjx6LEzYA0UnJiYooixncHpJjbdnFWXiFNYurVrB+tfc99fuyik87J
5dYqDBjIuUOPPlMQ80csID63ebgi5xN9uDVtcdfed/ZF5aCFzR+aqx55IYoJ5gNpQSUXuEz4ixD6
xMWz+3ER4qhJJPxH4EB9Gmz0wg5sazj7VKNb6DROBD8wRGpOWSafJVQWsa9y3J41IWBA4AkWmTT1
p+N/4uz9MVfHGTGkzEGgQCi/ohEgzvF0etnR3IQqgRJ7lu3cs6EHrRbbh8D0/m9u7fGH+msCYQIa
ZZx/uiQMez/89ZErkdQH1YD4k5aIHRkMSwM6OUrockQ9Tj0yohHNuUfP7LCdYishUJl3QdfMC12R
LEReQKLaycELFjgvW21hAF76LSw6/knh8Se8f2g9jTnnP/4gGZIudEbcBagNysPB4vONtpkcFi3X
VkYduyMI70utWTTg5Hno/Ud2wDnjfqyGHP+VHNZ6IPI4z/RKrQ4D+KjVlVb7Gsk3RwzRXIZQp3wP
U7/Eug6mxLZRWeY7IqzgZ3UexgM566e2HmZuyRGeonTavWUHxIgkgUFdWaa7nO8hLVPELJeNopSV
E7kKnlKSsZezyf/TMSG/DG26cXwvC8A2cTFc3c3PvCatmXO+KreVWnFguxScetI9VevsEfzBDOQ7
t3U4r/ipdVfzgJ7FDSVG8HPL/x0QcqbucfoSr7ft5uIbXW6uj1aV57apVCggBHzmBQLf3/9YWBSf
AkSUCJJwqXlff6SGL1o86FV14ZPzZdBUyWbCbP3cwJqbQtWGtvz+9KBkXN+JSdl9ImU7IJZsiAgm
y0POUKxMvLP3gTpL3st4U19diNQUcNt3qLP6Kz6a62p26ATUO8/vHmco1ICuUSUueZojTN6ydEB8
AYX5Eqxd6eLICznvdgJ1coz8XGzBoAsGQZpZWbOdth1WBTb+fsKBWlQs6AM2x839atEX4kINoLbF
ILodZsHYGEhAvmUDjTv1Tr4uQXDITPLCFUli+dGqH8EVLxNjU0ec4XQ3YUsPTLb1YPLohu22MmM/
k434JnC00XAqI96ulpaVI1zkgPFKGCggd7u47Nlii4jkdK8qxku4Ys51uWRIJNQr2QFJgF7qtHYO
8yEU2bsYdjIz9oDjS1ZEqioJxcl0VvXH1XSxhztWRCve5Xgzfg+sgZmb4YooA/1HAFD9JSzva+aa
FY59AzJ1gMNCogoI1KPAgO7GMjn7DO0/wQxogSX22cnThQZ73Ukv3hIyuF53z3YQjDV8idru8pXe
qxF2tyF1BvWwS7AWmyR+RcWdSr6lxa3uIq1F+qmZeQ2lO1cIkjhGF2/DDGKcB7QtBCF7Er9MzjGC
1TVoKLKpoaX+odos8LYTy939OvtVW7Vioa24bUwIwSzjfdKc0I9BBfFCr3ZILgulkqDGT7wTJMwi
MyVOMSXz9iEtW8ieg0AsI78DdYADYa4eL+Cl7uj1VyD1kXp/6b58bufrkYeSQQEoytKfowydQtXv
GRGtyj/QvsnBv46HbTotj0uDSFkscv3FkT0ahSKSEPNAr3ntBq32EZXm6FbQ4EzEGyI/PJ4IT5J/
vsLHwObwSDe9P1bkuHlOeiF3WILOqv+AMUdgQVzLDTF4tAt9GJ2d01xQUHNzhvu0pdwU/Y1wInLH
89z2moW10px8g45SjJA5qWvAPUVtjsMr5No2HP9/176MZDYtlK2fGZV76755LB+/uN0jmdYmNFsy
SET9bZj6Aoe/PZY5CKvZ7NYAFmgIoM3admCW0Vb23JvElcLBcC20+A55eeGHrQSMgyZ2U/HkEVoA
slEjo3el4bL1kO/p6mR0kPOGFgHdl9FogvppwOXvLzlpgQ6MGXEv/VguyyyHWwNXn5wgnilVWCAd
IdeseIQW0FKfVN8Rxx6fr648WPdEPTku1ZN2/GxJebRoidoq2hL1roRSMtu3y0UlLp5SEKTroXqW
cTjSjjo/IrVcKoV9JUVpKA1kzzBQKrAjVksOtXwatb0Ed6RhkKmUdMtXZjTgQMaQ8bCaD4UtvK+K
ATV4zKOUIKaPMnpH+OWafd+ow5f+CLbph8VysBmkavYf/WHASUEIBrwQ6fGZjbcJ8pykUM9REOTu
fY7FRi5u6u9Ihq172wKsOaGgQB6XcFb7Su91zvv26D/I3/Kv4hx/39EzU5HAjOYrKXgcOdopv/3U
ZPpczXDYGc3cJ/PayPQlxgYTMbvarEZaJIUZQF+p7bMlH8rHrzaDz9NLjC8Zlqzf3rbostY3zwET
6eilydG9/9VBHWw8dzC0l4F24BAr1/ZqKcXqCRwAvpFbRrkbalWQkq6WN1xumgGUhwpZIk9Lg/IB
m/DbxLH1/nNrOaGBDOZgzNgzZs3wi2zHWkt45ap+CAKzOEQyYkNZLDQC2yPwUiQpawmPke+u+Msj
xbtRALM0Kdnbue7Xv45gX9CFA/290GABOHY9Wuehd6rxWw+OJP4xDhIobPAM8sm/LalRSXal60NZ
9WRX9kJskeBicJOynyb99ubLBcmdLMwlCFCHdqwvxJDi4V3L+sgqqrjnt54sl6k2Cx86YyMo3CKm
qVIC6BqBg8LjCgCcFuyviMaDep+Z0X9A708rfbAzKTmr5Cm/a7i9JIbRzZ0cAWWmOWcUM1qyChIZ
4elM6FW2wx4akWakwTLBEjeJqNUzr59fYVhMUFu0oPxpVeU6HQ2+0gbkeRI5/icU6ZijDWKVioTh
ir/mJ3gkY9/qsVqwfXFzmmR5EH6JS19U4a/UwULIILz2OOqcNlFgroEJBJFZkxIXRbawzW8iJbNB
DSDCCYAPFUBnyfYrHqF7v7riR0Ve9QtEMGCuM8GuDpPIi7Mc9DZSE4ykeRsuS8zNHAKUtt90CQ2P
SgBaUkaFeTsexLJ7mIa42rQZWdF4oLc9Xxjlw1WiwTLOZdC6wZ/lsKFlTglYg5rsERfKvC4M7UWY
IG/fVWGiyegtUQh8kkaJj41y3jgjLaCO3ns92+/bpnQVqTbUmhdXto0KaB2Mq4Xm24WqUw3/plik
F7bp2UpeG1v/fSZsDtm5ZsAHbACm0gztoAuMZRmCUDDlGEmU61zxBoWhpxyOoEUOQsrDAJ0cZECc
DEELJmMDMCe9Pup7lKkCM3eEMUgsX6a8nwmAlEbjK8c2EGOxYOaixjVjYsf3/Gx4p12yOK6HSAbU
06GU7VL+Rdl/gMZhOv6Z0a0qkLOPLKl2ZvmBu8uwHwDqE9f7sJvjCFwVX+UhZvKNmLmu80hbFDCI
vmE4gVkNEEwOQFdK9xDipM7/Yymw9ZYb8bzw/JSO12slSEWgeByv9ww4kcQQOxpIbbhyGlOKzrxn
Cul6wm3p4xZ4HInkiI7nLlmQdiC/lCbex43QEqInNQIqBkff+OBK6G5u3ZVvENJ5qxrlTxMuqKX4
Az/YoDk0KbwRvnEjZ0tINHxv2LNrs8iVCyqz3COyXQV1nsZ2PvrZEkItJbehNpnsnclwUEnjhnTK
ybpsDKPcp0RV5Xr1qsrEGzb8fFJuFVw6E5r+gBSqGwXKvhmkNs7VU9QNoYSPuU0fJ1o1aI5WBhGL
FLFo+WpEOnRNef4dvxmE5Duvls+b7iUtOU0lkgQgjai9nB1QbB9Y5DbkGU/1bBzL5TU/pLT/dabB
g9JXSIWpt+Cpc0ifPFFxKKQWub67nHYyB/Jshv4cCC/8mrks2xpqLvsu+g82ZVivvjI60eloOg7e
L6wrWuUQHOtjs+h0mkqjoQ6OZrBNv68xiQRIv7P977ImSWQR3cQTeR/r4U9xDZxemW7ul7BFOI5A
LXT38l72KOe9wu4S2XEyBuqve3e86sN/6D14oBbvrxz+A1YZUQe7E6sKsZp8/nn+WkqYA3vAk75V
2vIVnQNuIN9/c/JV5znvuRd1xKMuf3r6q/fpF2vU0D+pH1tb7Lmdk06GzMB7Vhpolje1yDnSitOZ
lGdI4h1Tpfm5cZ97S3kC9qOtGg4qLWJLXe94HhNLBJpuEBxE9mL/9CFwrxwf1IUuqdVrC7Juy+BW
qWRQiLeXlN6eBHpCQXyHn2CvLRJDhS/O0prhSPxZWdqvDAiSBD+B/+thAmm2W4zD2I7XJ37q2Hdn
DBoX0NGg0D2BP4gWz+EHXZ0HmG6KzL/QxxTpMKV63Tx+o0G265U4jt5EszCSvUgjFTfTqoJTXgH2
FLtG1diQEmUEALl75VujJzNCokCz44UNTAbDwIKwAG+8Z5SafnqzbNGCbnRzVvxIekFEcLU1bwzJ
OX4fuyfRE1KJYbJm7cQJDOrmXGPk6d01uKWTHvAzBzMn8h0udLMoKlAQlrzdFdl/0lPrbWLC5KqF
EVZDiaIBX1uIr+S1uR/4rT9nrehgirYRiUixuyOwHpkXhiyml+YFugxjuIQnhH8TiHU6OkSjNb3a
HrH3IKn81x8YR3Kh2sD0dcNQ/jCiQX53tCnK2wcY57hFLKEUKBDRX/dpOenstndEiyTx6A0yva2D
QtocImOIWRbECACAusKtMoWaOYNf52ih99vUKSnsdX7SJEKYX5xQ1yBq9X7Zmv1v5WMBkqbfTfFG
1C38uiW/Svs5CbARnDXFAIurDSBLTBvS4eGg6zJcrVRP7NDil2od6h3RUdIVm6tq/L70pUJ/ZpKk
fCQ/ynOQFAqsS7igsFySJrM0w5XEwPvjVrc7AuOSoYGQ/NdIhbA5G2LjwzCzEevjPRAaGzV92iPZ
606QY/GJrtgrmRJZt/C4dqolC1MASETSOP79bcEd/a3MWL50l4X/XFDIdUWcHqY0TATPWAMkvSiy
xlK29N7bCENoO573onvAQVDiaWzwECi3MyR4wj9UWjagmqIbe90Zgcqh8Is6kdXDHgsXuCDXSXaH
rKh7QU9GOfcv6fAdGytpd83d773WqYN6glfStY2QEM9yj/23534iCPctPrBlweohSyMIKjJSWY7a
VFVDz/f0zgc4hqyIfY93XP+0VJxoCy6Bqg0+9fx5IF0jt9J4+4ZdQ/AEgNZOL6ZWIOBMpd7xhkMa
Ja94FoRbH3F/YxAmqFEci2y9p4S1k86hvRHRvcDOhEEAQVLv/sfhP7Jdm5j7ruaOdAe1lVzRQbgh
EnwYML4LXj2DllCa6qEENNG00ouoFxdy4aoo0xDgBY9MRsXHi2fz2sv4LfXKAtGwFsynDZA7M5z+
fB96eX6DPlHTYwD3t8TW4s+iQJsmxiuRmjgPrKfXAo7MvupX29+0aadv3t5QHc0R2vnL2XFEiLGB
xh+qcS6bW6N9ZZ9Ve+e3rr2SQmaNblpHT17PhlfiaJOItvgA33PLqtW8anrZapS6+JlnMgokCZTs
DCfB/kMi5AxVGfIKwFPbLrpfBXyLFESncSxaDuriSqxEFmPDXi/FpmZWIyugyYJq4iuAipk6PltQ
uOGvYs2DfC5bqDq+U2DpxTCJVHVee4aRB71rWIOnxyPWC9bkzzA23g4LSeYKUUzE0lcuwLOTcxNr
7ueiuDdlFeVPrqiXeBpOAfW1SCM+yql0OhY04ucmPSRgAqNEZAaMM02up+BBkfMIeQxgxp6ePQeg
oiDIxe/y5JZxa9oC6OsXckvJElUKW5nvuL8ayVeIRve4HfmIXz9Gq+Cl7W92LlbI0Ar7i+LLdDfC
1bz0jaTHhUQM4twBv3j9+Wse5DKglOh72iIeEJJ8qtyYT2KgKPUA83jU4Ti1GhHi/kBFzmWqR1Ky
wSgzQlZ6kIrZUiMduClxKI08bKroSgaITrArap0VBen+FCTPw+CX2nScg0ENaVyfNuu1oPkeqEz4
JBOy5p4eO5W7IxigPdLsH9OUA4cnuz/7sZuF//qwaoxKEvntEQQJ1tZVgXvgdL0Tax0UmtTu1ebU
cvIzyNMms+N9Bc3T4c5aZRrqm/Cg3fROnveitCbUXSw6dwJvhjpvNCikgmHKqSYGMfxhcTpbJBQE
U2boPTOMWe0kmRn388rLh9rYxADL6kVGOFHa9xAs/1zOtDS+/epoQBBqt96I48HJJz1E/8/9h8+v
N3O1rSYg0VUvsc2yM6n8yzlKEfhaZuCdGe6wNQMgxnEsH85+3AcdsVKG84EH/H/c2sn7w5ZnSl/Q
qKkoDQty+UwMMFCIODk4ygEAwxQ3eWwst5wQBZAhlv7rlMcZEj2kCNK8NAD0b33VMhh120+4FFPI
OTMlI/lmP0e2W9XI2QOHMU23wRMyqJcJajyIppGgh4HMXdfvvX4CrGLaqZQq5pq2Q1JdJDJo7WO6
pqlDXY5/LVaN6laUKbPThbvo0unfYzNs2thlrePYCvS5Aoj0lBYbmaJERFB3dj86mnQbPy1HwxHl
0LW67++NHsFrMAPno6FlCAV9xyb/k0ze6JyH70YPAlg0Sy681x3ylO9XABlGyrrrgPlDND2IihpL
wqowIrUNi9AmqPX0Qz2fPxqggaRdTov9JklUuxfole5CvzPjqrP3NDulosknZDwcyxES/d3fPBLU
siCXI2SmcYAkoboF+vFSYVeHFPQPOOfou3qBL9dD1H1KnArqRPH0oPOM0QKh4ql5/9yAk9cI1zPL
0kISZ9IUltsS3/xRiNVmV+1LQRO6AitKRAU7AezGJQpTxyztKzndz0IWLx5wLNgzo9G22WFsUOxK
gT5G5mXEtkxOOBwWCxoTvkPXdjmHfDwuSN/awfouOY0Lmjaj5fewfUn65QHlpAbo/t0TMb9dVSC8
j0aZqpTBI0kBwVjq/0jQMCH6xawQPpgAFxwBgI62MyMjoJwJ2ES+gC30iAVPnsmAJ4itg2gPK4hR
YFxgmIIrwt4BEL0hCvSi9Y4nc2on9J6sj3kXP6hOTvPOFWvo9e5VTgdbj1wbcf7Ov/xQ2IokTqEe
nET/vXOTUpaU5qVbPYkOdGVYvGqhe5JY+7iQ/lXsrjUlLiwe5c5RXRrAwgg92L18yTNPRr2PlaSD
nvuislO6te/TqQL1XIaN0ya53bjPs2cxsmIqfQ2FiOXwGbISfQ66FCjJZ2PFUTW6TsPGNDHjnPT9
UzQnq5TBHQeT1bmV/fQaQN6EZplP7hjJHo+WIOycglB+yjL06Tz8heJ+pHa46rPV2GJPqGJ7oXB0
LrWKcXbhoikPhs2NQ66uQ2OBTHiMBm22nFIoJ2gkNvJcdBbkMR+P+Z6whusJ2YL9ENJYqXmjLaqi
oVS7Cr7REy1YdziLKOy1pF69OIYcZ1he6mLaqmS7ois3QG87Dy+l1A5fGgAAfUZw5rdhg2cHRaR+
VjadbHouFw2n+e9/dPZdgW2uHCEDWfIxXttXlsGCASvYecdesgF4yZd/N7yDr9LXuarBI4hYe42C
TOyTeGrMW+KEL2LrsBSbEZy2sRHjuKUhW4klLWvH+6fu7DAIkFi0gLZCE5Pw4butJ2YGr5HYzqd9
JTP42513AWN0gCjvfO/9BBLcHr8v3fA4T/10iZpnOPiH/P/ZyuGpOjLc8C0Q6ebNiR+vbTmc8vDH
NL8AWsnYzdCyjHTUzeRJCC65wbeHvjnIl4Hw33aFeYJSrgebzrpQk8ReYCkZBqXc1NRYMMTsS3lX
LpB3aR9NTm5WyYEqp/nWXfjn5Dlb6eH+Hvn9ICjPKD9SWYfwgVIYpsArEpJxrF3N6wdRNm0oS6jG
PiQhEjmRl3fkGHtWhT+c0/qWEQaaFC/j9E3kMrR/gi4xSll+uWXitA8FAhj3KV4eiJv/SmLLN24b
cXw3UYbd3oaOu9hgM+S2EQqFLkXdsktfh4xMSJVRrdjPSUvVZj5tQnpy3z+mUWryoupr/zD+Bqe+
rnIwliJa/IiCcREZHqIiJ7n1xpAZlqa+DW7ePgdNfiuhlfCxTFZpWUPWWOa54Mz2Ksi+HBeJ6b+M
9CmpFS+lhAx80+BN5OcfFKSDUWB9qn+DvkvTyyHMMAfzY7PM7tq0wgeopI4rdYUk6wsIIktf/yZE
4s6NaoKgo9IVvw7IUkl2+ymE7fUTqP89aormwef4O1cxfqbtIiFRBjdEc/EloW7rO2cuOXBmfJhl
aEE6KP8qakWnognh7B3+lIJ5jwRoab01Lia4UX1CILRL1cQjYasFQPEsYZ2/DNcBo8sXfP4enWcm
Nm2j1wHVTelIDfLPy9LzM/gEmSxeids7XLj0LhS66+zDHOr9kZ++eX6ynHX979E8ldLiiY7nBGCl
mJlmG9w/ZCUJrmABgAVBmrtFOATOGuWOLNc9mZx40Lejc0BiS4rM4L0TXpMlgy6l3LIt3C1scxtX
6BKs/7nvROc3EsxFxS6o+OU0ZIXKXBsm3UC7DVtUgM8sAlmjSSHTZjArjQkod6eEPrgpLX/1kk3d
0JLTiuKOhsjdt3H6AT7ioyYO3IxrqxLZ8GepCPCEG7tdcr1mHsTYNhMUHfSVbYEGz36xOlixQNsN
ywa//qW/RShpM6kKRHX+tqKPqhC5/VehVlTN7Tz1Rk+9XGO6kt7qYhAVuFYNR9dWjeXpUPEbzHdC
4ir/h1fdN0SseChpIrkHI3B66iq5rLnBGWwywNt8VVYFKc+l/8JGtnpaOhGEJb9lViJ1VcnxcEfE
CXbcZG+ZNgGRRcwv+iAUNryXso1fig+EU/dkTyrjz19/Fa2EtN6quocYtTPEermv9zvLa/0pNqXH
BRG+H1LX/58iD+Sl6AFL6ea2KkxtKEY5FwOA18sgtbV7V9/oYpzE2ijKPpc+BPWc/djTvbVnyNuN
Kv9tm5H1TtvRMWR5t08i6L9CMQamQxnbG+ScgfWYGmlL9pIQycU6Pm3Z3g8sVHKLowBprP1RhyVy
oUuaenQM2POTnVj9cPU8KoYUhLEwuztsiC9w0UeywUa3r2wir696uw6RxIRkcHb18WSfB9gk1yAA
lBkoYTyu/g32EO3zraU974qFRsEZ3UY+9jJBumiePIDu8SNoUlU/VXihw3NySt68JANEOB0plCOi
mq8dJKuSBZrRSvdhPiZS4v2CXLe5Z/SuyTNCN9MLbYerwK85dpNRx5yt37x3tErPPTAzqar2qtnK
Xw9XRjLmPpCv3Jy/JeCH42lX4xXRVjqvSLnetyFUiV05N48GmaZkPzwB9TwMRVR78icM5GYqUVax
XmSvGaoE/dVphWruJYP/kNHbfOAD79RtaLLMqlzqTbBhxb3JG+uH5ZfmWjCj5b3W8Y2nZlDajnd3
0o7yoer2pz8tfcTa4FoTyV8jmanlECXCx7xCQ7J+SD230FI+AHtorPvfo4/+ZBnGyoMQeYm5gmUu
eioF3o4iY12W44X1zwECNP63NZIv7MWrtv+Gm2KwN36Tbvs9M2wZml7Go4DOM6t+Enog989OeEmu
QPVM0cBoqti0cOjzhtCw/2ykyNTRJ7CnVB8aA4xv2WzxNU7yJY8cz4b+nrNO/4j4062FAwWhSjsP
LgMOKai5AbWGadTtRfLBQLKVeBFYT2UL451slVgThPOZl8SstRm0JlVegDRmUOz//F7mYi6y5bO0
EfLOxrouSEN6nJaRaLS+S4dj6BmlTjEoXESRU2XjzIiLLIRl4OPgVK0BBouW7badvVWYGCiTd7t7
YcCBHJv/w2i5/Ku55/iKJmqDoGDO0GOE9VjVmud8Qvfh7cAiToqIcDmswjI+9crEDJjWyVu0ppdk
xrG3fAQ4jcfpxXSPle7KVlp0OVZrXqTsSxqQmsyeBh18BlGKBWzc9m8UgDyH6PPU6DljJcymh2o0
XWtUjG0htcrGGqpdCAf8Gt4vwOqzyuokrevKlldFv3k58YF3ZkPThYjVLOPpmP4r3aNskSZmA6+5
REa6PYNFYZbnZFC0p5ze+1KQW/ho/WCwc82OMmO4tJ25vdBFvo/28LwUMslA+6vd6zjpuIE51mn0
yOPJC4EuxiL0w1ZvXky9/+JHLqLPdQeFiSR1JODxXCcnk9JSiOOEuiTiABKl/6tYL3pE9qu1+i5x
jhbeJqnNSz7eZivjvnKXqnOo7yuCpyt84sDKhesrmLQoLl9OWAXQ49nyM8mlY7erbsKyTsHckHUd
midcr2sQ+oIL8/UNLcV15P4z7XPtV03G6g6Lcatu3z12mOIA8Ydg3i0Ikzo6OBzBovhzCGdBav7K
bdlcBVN13z76Zts6lHFi68uVlnNKpManKBVkhtBHRi5LjgaNTA6wVum7VFpci0KZA0V8Lgri/RaM
H9J8CDI4fyfVHJ8renALVm3qRiYltv3oR29QH6Sk8ncdIWP3lTaPWokNRzt0AUbYzk9BlkqW0sPZ
1BznZc/wCK5YKjC1BKo0jqz1/edijcpeHtIiRZzR4Jdwj0Rx1S9T+9ZlNgx5bebxItyRpipTfR0k
MZlyB9w6tPPvq7wYuLF9edj5EG0ZSz+ykNCaSZHi4r3MqE2rAHxqRupJdYCjfWNqsKi04rMXWBuE
JQY7w2H+Ya4y0SYcYvUyngOd6agZ7i02rbpWC3GvPa+guyXVc7KsSBcf+soQTmDRLLx//BN/aoh5
pybdqtWgm+xRg6UdTBXX0UPkuHfqbpTro9feC86j1y2vzSNTbgc4mJCr2em/QIpPpT/on5Mbf2yj
oBbNIOmU45kUgInyzKj8zSUry862SIrV20JegPSxqUfXFBJg6b+cL46a0bgZiRYJ/DO6O1nE3zfL
+9+7edPrHJijZxunBBAveBP7Lh+TTGoqtsFGDPh8QAHFsRYBg2VkM9Lf6Fc0S73C4aom1PBNHjR9
MbiiYu7vHwaB8uMPkuBePSjC+jt5CqFvg/JkEEIIkWnR9P3zCThllq8eM1YOUrsHRpu87d0vZ1j9
lgGSZUoST7FLBw2Uuc0ufg8CgRwhBxZq1Wx2pPmDiSIWid3gg5kHqG/Zk5TQsoG/VBCI2dhJ8YcQ
45F1p76CKkNIUQQny+FhN6KjfwuQrpdIUb5jVgvZTd5X+Z78+gJfNwZQy4RIfzAnndQqgcWIbucJ
b71cngx5jY9CL21sJ5MQhWOdNorG+BH1g+7L/9j7RRsyJUL/FZaDAclzxC9lxafu91x76xQd+Eqd
UM7o+jxvQkA9ReQwk/8r98tYHGcu4CYkf+2JcYVfwXIj33Xlpdr5/7gjLDjbODzA8geMGuM9iHHe
S6wBV/YJQI9Nr8zPSMXJg7+qYWlAHJYQH1nZo2Y57l/wT4RWMna9UPtgShdJunyLxJOsx/19f4vK
jSRC2/ggADDKUSxPzqor/1Lq29V2bO612QO9lpBOvHfb9umVA961EA8RLeHVjyR9CBadw/ikjiy+
A9as9w+i+PEnXzKXpzDiR5RUK9gb4A/n8MFG2hBDplqyCDCDoYLBhzvyR6o7GOndVSY404DtNupx
VThKXcxXRdBwXfetXGVbAoFLWCJNwnO7GKi4V8fcBtt1+d4up7SDL2ivyhraJh9UvR+NdvyGEMKR
pbJnqwdDcPJyAGabxDT75UZRNFKJ0PX6nxHsWc2EazVz3M/08WRzNAsLsAR7n5zwkl0piidHrC8M
duhBgzSzHc2DS5BijZQmX1r++drfyBknsgra0mefV7xmC99m0ToDPpVCQv+ogu2KZJbYIPO8Zd7O
6FFkRUFbJaXLu1rpQRZFN0b+PeLS8Jfp0Vpfo6oHqOXO4Wmfctmm5afVfm/FwdIUJOy4aXt5GLKQ
uzmG8HE7lFfcrg6UQX7oZvpquS8wNd1k/eMV6/cIhhsmWJIW1Rc95UQXvbq91kdMIp8vnaXdPWhb
/2rWH/zYfNSdmBLJR354gOe041G67W0nbmKDZEsZ85DJWXJWI2hLKNry9U6Dy0zWxlWqIdT5U6hq
FwOEnhu48IAK9A2jNW0vpH6nNR3DufOYvgG3SMB1WI1K6imx092cWeAClKdudpNIQ6Pf9h9N1NXs
yYBHv1kVnE9w+6XMFI4Yh2a89vu5Z5fct4bw8/H4IFKTAX96R45tTWUJldoMF4VsF0hmwqCAgoi2
3RLJfLctfpgEJVN0sMFIwxyNhir4VlXne5V3lDKp7VuXKGS3BdY3fmHrDESOnvUBej/VU+WzWuj1
K7Dgv6Kzc4/xNGfdNOi/zSNq8Hf7fY4xPtHZ0Wcd6YlLEzJonU9bBAJxZ6n9HnjhN1YD+7YKs1HZ
kFIK/IA/S32C2+crwzZG/pVMk6xuE2AUmozWCPMF0t8CgKUq23eim0MZ47wreofyHYnFywTvLPmc
CKKaXXOaVCXoIv2QrBQhsDb1jwYGUXrttr6/sWsLgdK0q4+cWacYoudb3LYzlWWNuXwf/bEuh36Z
U7YnFA8FToYMt565YYDiFBLxbuWGfK0sr6K0yXYotVfjwg8O702Psas5JlqYRWg3TAiyLJ7lR60w
CnRpRO5kxQhraWTPspZS+KGJ0LJ+Lk3WFd1SdtcAb70jAf3rCzofVeuhZl8APNm2UZ1LmW8WMOEU
TBwIYPOPDz80qfbyuYXrPJleAl1jVrbmfji0yv93tmUiYcVDd/afz0hoHAdknl2CBFu1kzjvHD4x
GCYykEdmgmjSpKofvhc1T0rhYpPtJslXt5/lpvtOUOBbvKVH9pE8oZ7dTb7WR+G5OFEFJTAsedn5
xDwW9b+iOx79SUPe/csa5s8hmcVuAvFGDKvqZtOeqfIyS/JUuHyglyuuFyhFqhUEFIN49w3CgZne
2UIoo5FGi7iv+CiV/nIWgGsTWKQQs2nKKRU/soocVg3OL0ZW/JmdolQjlSaUKVyGrNCJAsfBmTCs
AP2BosRPqaskmRvElnbgIriOsKeDVmxqxd1tGDn7nfX+POCtfL28fjcDdDqLdVrqQVAI4HLUF/ga
mvymraNTs7OA8uA6GeyMbJMoZx/Rw71dE/Or/9s9xMr+ZWH0dFgTqzlYdkm0ji68RUiWOp6h4YsV
Q1xzxcHg9dGnf6kqw7xpgqZSOEJ88YkqWAX5F1c9aWI+4BCjzvExgv5CY64tCOAgCxjSTniskL8K
cuhe6ErgCvZoM5wZLvIhtrcVi2/NoCfIfT7yrB61hq9RPmvJI6mseQb6ow67Px5oSKJPBmO+osLY
aYZ3vBbEdsd0VfgcT0+eztYvw17GTy2g2oM5PVVovaimuXwmm9d02ZEf5hFCjgyZeLFb9//dMnun
AHbEcIjZs/qYkHzXdOVEMFsBgapw+f7+gLUyjM785r330tERxFKeVKbTU9BXdFJ8hqofOs+2yxum
6XzwhwYk+IFfzhmATLV3f/O0k02R7/VqZ4/5GrBfDwAV+7+c8RR4dMp/AJK29/NyjshI8PsWSGja
D+KGvgej+Dy7JqKDUxrWq3TWvvZystbVg9c0WAU/tRqJjerwxZs2jxyYf1JvvbQiZ6uPWV2YbUcG
pMpjG6sHyxQOn0rMr/l4WhgUcq298dS51FyFAu7BSauIpTLPsiNvIKH7/Y7pyswjExiT5ENvK//x
UgnmKglu6WKNGxQ89DLvHs5ih0q15l8TcfaAISPt7Q6C6uXZfE6e/OZ2E4ecsmwq5Dn/8dxXMLBt
4evP6uHViB7v+vhHHUM+at82yF62tcq720mtGwQYxISpCytU4fzA+AqmolY7sM3dVkEEZkFOjj9m
/dN1fpgTkChytU61GH+cne+ZuCxAwjTzYQpSfTWlsPNf1ANoz5BBvTczgWQ5dsCnmLGv3XLt+iV5
cZv1ugxmOhHhcB1Lj8iPPb5KuGdShGOi3UEKT7MczLXckHIsykhbVJm92TFG83MbzYstxjgcAJ2O
4QbU/Uqn/UA/yEkfY/W/F6FaHDS3GvFNo8j4BjMLyt9aow+uzEeui0/WMbG1TdI5vkW4r8OTSiyu
ypF71kj9xf5+9bO9tg0yneZawhIgfY3uBd7wmFsKwctTuKO/elExJ6UgTHIuDuqHv1IJQ4jzDbHf
DgwIsEtUcS3DAAGNtQJJMEJ5/bG/2kMg6szyqad9j20PHY6AhDrrU6EF1BdpS4ZtT4LMLQBaUIKV
TgliD0ch0S+eH7/QRWbYZ06WIiAWKz0PsH87MM+Hj/AWvdaKaC9dpg+QNq972Ec9srIkqmMcm8/U
C5DrboT700z+bafYxUxTwgxXboYOE4U9Mz84aLmxGm2RBwqHB9AFmoac4p1oSxzrN8EHy4CPMBrG
ATuHCer1WJl9rslgtDVkYzqr2CFF21t4GJhaqYepDrgiCP2z02ECSnKejYY+MDIDWXyTIZqE1I3w
8itGfzCqA6nZ5KjH7AcCiqO5Yd3seKPMnRd7IF5sIYstG2OtKTyEpbAeCltfXomEpYWYIhOrnYUv
NledbY9ww2Z7LRiVKB2Bd0f/S6iJ0fkYzc1DRVFArjcnnQSnBqpgJIgmubyKT4+o0Cn43v9E9rQb
e0AriY3UWWRc8RJ9Qg6iK1ruJV4uz5m8URbBiVVZ0FircJ689CCpZMzoDPxqQLUXVsXy5mjBw5aV
YzdHZYubM6HqeEpttmUHGBVU2KuCA44XAOnYPwhiTs/xfeH2HdtmXlVe3DiRPZd92sOGymBDrr5A
FBtr7BwB1bK97whgnQ7Wl9gETPKOqjruWI/rs3jCRIpxZmoyJX545anICpp/C8Quqkz1WkTZJc1b
mHlnW8Yu4L05ls+v+9o+br+cx4P0TApFtiCE9R6K3yok3VvwPYcUQfgGxh59oECLDmf4N5ioOjML
V/yC4tFE7/F/z4/D3hl+NfSkHOleo9OTJUZl85fmLb8x8w/RoJDXjYFwjqkOboh3cnwhAatBo/rh
0vClfwdJcyRf3KiXLsZLWl6esIHAIfTy+ZLvFFanB+cgOuiGSvJRggcQh66Nmb5HpSyGaXMj6jrB
EXBsrUusWnP23gnZGGckA01R4O+FU/lTX2FnkAfpwDZwF9h7z5Q13rNn3Pt6y9aEnT6uSneUJt50
iRk8VcSuF/v1PXZOFk5qEAT4nLJTTW5eCp8CGKK1sRk67w8dSrTjwieegN/QyYoPwXhmxHszkLkg
8Gpm8+wMP7CzoUHKnP52zkwpF13CLFiftOINXEQK6A/65XmGT3DI/i/a1dNvhru/y429V2ByR/IO
KTSJoIXTfd4c53ebNkjAQ8MuV23AyBreMxFbWKByXQKE6gqdPyF+khm02z7aln+NlcCQsgF18FxR
KForIUw31bSlgycijRXYcaHbjmqrYhOF7OFkj0vpmZU4tjQ5cD4hKerkl1/IAZ5uWr/lJpFUXrOS
PIOQQejELoCJhrTNZFqCIG8P47sXpkaMA6ci40sfASRCrryMPcjRGfpdoM2Fw+fQmocWnVINyXMF
P/je6Tuh5YRkmQVFvROyzDm+qD/N5OHfyJ9Wz5VpAwF2JKmeAllBzxfWua12lezVb3qqzIcXde6n
rD/gVVine+zpof59vL/YROdb6L2TeSP+K4MUzpVEsUezL73Yb0jEANAkuAOciXowDhfDYyMJB7GB
6XCYw5X+MfXDrcrZNOvOPqMYxVz29V/I6voANu31CoeG9sSnpABzYsTtjn9YH9Zvt6rgt5pwwRjD
7lpq0ZhNodU9Q3u+uZHZLAo4eOyNXFSgnjosrwGACibrAetItHdROXU5CuXbh4srG+9AIdXQgfJC
iHIoWMfpmO2tPpkAMm9UOED6FYakrwnyRpSd4MDP6yG0fNVMtOkDapq502XTv1EdQeakYvchVhXS
6buqzcKGQBWftwVQsrrbD9SNw+GsMp/lyhZA9lDAqXRepbUko0mpAhSTdHmBQ+p63wNuqEJ11hH4
AxWf2Uk2ELJOVXu+jNfyvscMWL13FH1wbrMM2jPXRTolfo4ngF4iQO2+FSLun6IzYqNw27kjS3IE
dCCeQPxIoDhj7lwWewuDq3nzXBmT0jRhaPikIbKrnDChykIbt1xNBphFC2S5yYbKj+Utjzlz9USl
pl2+DqaMpP8qIUC+E/DHybR6e1CxIWNmm6AFoaHLDkiOHKU+nHn50RKIap35coKulh0xEMM+XWF1
bL8rAwKWKp4mCxc1jWKWLt8vp8Nh6Ys4K75FWpufOzhj9AUxnhf9PpzHRtKD+kG1M1u5EXaep6jb
kQS833GJkserLqZYWvTyCWuhxROsNWt+e0/j3FQ6ibqtFllo2VP5wi179GCgq6liCpF8VUbdYTDa
VZUvlF+4NR4dpAzkTNvgz0pjU72zQhC45D+MPWFQa0TbzM0ymXPuTXyDTy390GWXzQyyqIEsyApq
3m7f85HETw6Lsxmc7bWNdU7T+bR7X74jtt3OsQolnwqDjwELi+bVXynb5S9etTh7aG9DqxXQ+SCB
g9gnFx9QO032QkVhL/ULB/9dK/6A2gIbU3ag/WpupLOeQahQQmDDg4nWbRKNIp+O7Xom4J+Vlz56
uAQUpL6O17VULBRBwfOaSPRoiTul5gROIm8IAZadwBRLbuf9Fmi4TMKOVcagGXAlGGuHfVz3Kfww
f0gjhhEXUInaj5Q36pgom73On7DHEyPBY/DVBqLuVhSfI3stSxQajCtWB2+lS2cn+u948iV6HKRg
ie7is3IN+aqurvcNJ8ywLhnisaSmUoCG3RukHqZIdKRBjw9FQMyOsG46mPkep2SgbrZSKJtQEGRU
UTgAfe26VEU6MJZL517sG6cMa7KSCl+eR0XfeSed5qY6Q6m/G97oA9/2MKhFCw24pE4jXveipIwE
OUnCW+6deAxCbe2LICdb2QTwv+AnuSSrS8cTmwqghH/U5ukaKif0gMGJq8lLzVeLKpXQZFBfyJOL
nXPSC+L5L5f9dfA2OPNP8QK/6kVXN4H1FUMucUW2A03Cy8Ii+OQzZP7m8UV45omjww1K+4hHIETX
q8vhN31rr+SdOqJk67N2WXmsW1ec+DVQsZJycvJXsD1kBpH524KLRsHLQnwtz4IUsUV1Pg4E8GjV
8EbmL6cHqkcIHyiMFs2lE7K3ANzhdWIDvdk0jNn7bjn7ZLDkN+B0c39sUfiwH1J1jqD3YAly8GAu
mBxLVtRxKZnGgySmIcEwTHjnPYOvdZHen/4HtJtlFJiS4nti9CCKwsPGmP8yLY1HxjSAjVTJgOb7
xGGBQGLS7CCN8EU9ZNhWMR5l8HhpemLu1nRikPRy9NNUIOl0+zT+tiOYMXm9LNJ1487g2COudPVA
qWqIJATRuoj60B71w1BKlT6ZQcFrHkKdHoq2q9OHuMkgu2dDSD9VmD8KuZ/G5miaIBkA1n8gYKtk
nozssyShtEm4+7SyPvdYqtrQFTDyin8gdKxKDkkHMUBQovcZvoIfM+Z94+KN9iM8UvKPEryrkUiQ
CrQUZZUgBSTBQ4AlfbFix9YPamDYDR1uWEzpoxPJQq8vUPVtE3fZNf7nHL10ri2O+y/GjAq3p6rx
tRfzEXnMXKeFY1gl6jYlmZQc1HBh/WxaoK0DUT02oDw4xjmzt1KwlYwVTiwAup41s8Jm0LGoEZiQ
bplYlSTa974WjarHKkVtjcmbSzZk4TYyTTf7ABaWw4+pkb1vVkkDX/tTySGXfeTOZ73uyZ1Yrubh
mi1s8dLuuytpdfxKUBV62h3RP6BsZEnTcyuo2eB5y3sE7CFdqMTfM+i8UxM5VAv9S1Io0i1Pmulb
ehqCdNvCivfA+4Ya9B+2hSZh6NTBmN+xMsXFcdDTcKbkWuRP+62xCSHxAFsLOzh6MImdb0rsbS+g
6gynXCk0eNmauTV3gaUyUOyhHWquXMziWM0ebRT2wzOiwKOKpzoD++mKJNL95G/a/Y4pFOhzZmmz
m0VaT2d4T9SGR1kQ0l+lieWKt7y8wyXd/ssP9M+P4uaMBg8+v9VOOukXRdtwR4aIqa72lsQ5GIi1
K/GuNsA3/yuiSveloWN1tKDaxEAWqtwZydBFXH5GD+6Jj+5G1UC6xAj5jlrRBzbV/JjlWfsx1Zb8
RJ188vzNB7c4AUIinUmx3+nRUI7Nb/JHABz+gJfDmcxSaO22GMNPiLTJkug1R8UVnNUBJnKyOx0J
8jqlCXS2cxC/s144pVLxbGbAvkofjRmUEJQifMI4DrjY56scG56XKMRUnb11rTLPQCGR68ar/TCv
exqi1Uc0BIepzvN6K5aknwaxzEFkvaowoAAtpfWrZ8mFrr+SO1z5aeh0+MxCizop230mCtDV+DqB
Bh5TGKbUPWw3qaM2nQo/Q+3csu+PlpcP1U8FTEtIf/KgGb5SN4hG3KiQ7Iiffj/2gSu+Ioql2Zzw
iCsGxhwOZTL5apLPowhtVz9jnvdrn7JGMLIs3XxRyhgf3wX92kiyS5lDAlz6nkYu3EcpL2refT0l
UkAnFS8KRGZmttKwz1+Qqkfokoe1Pnaly2yc7mxY8KD3hZ7nR1S6GwW5HpmWfiklzx3wxngYV/LM
edlUiHD9tmIjDlDwsFpmORwuCxIy7KKgjuCalf/kEhx9PPZ2Rc/qy3uqsjbKXeZ1m6EjAOq3WF0D
oDP060af8JsT12/8YGY6P9Xm0ymlKPPQEGrIWN864vCJVcMkBYgqJaJKJ9cyMdGDD5OcuxOrGXJC
64moQ8eeyuOuQ3MwhQm56uAiUCEJe3+0Vlo4Ktsm201DQiDperoudLgMispHVODxXI2HkepQGEkS
3LyAaNGXb4IeTJbtDNoTaR2f4ljcqWHyjk3j4gFgjgGZhfCzQsTdOVABIrsdGIqMSFedVyYIoE6r
SjMAfdJ1pKDjwZX7yvhv0j4biHVeYfpAWGMr+wf+GG6l0ZbIEJGDIZFBES35lOVho9Z0Gu1+8B5N
FwSm0ArV3v5AqXkNQ9wo2227BsUYNgOyTBY4knabKC9ZtkeLDtvgV+ML9rn+Djdb8EZB4/Kc5iDz
fR8eiTq6fsOclCt+9ETO8VidvsL5jOzJBGBelBnWbcYVbfJ/nTmy0fz1+y/2RTMYe/gY2B8EdpDQ
7Lul/E2p0Xed9Ra00GGzySvVMTt4PXIPj4aSMxRMF3i2fR/zpem1X9qkRx3/HK4xtGnvlyY/758f
7dgYOL5o/ziAs9Wwc44OVJIrsXUWkcaPYaSszJuoHT0NFelU1GWIXNQGdpsL8Swd9FRR3ECRvsDh
0GpwW6MfhfG+XnKEsZh7aT55BemTt0Jo0sA/Wpwk3Gi6FoVeekEvxUFuWPg5M6F/rcd5gtH1A1nK
0xrgCHlGVLHkjGqeQupGsWkHjWYADKfg1G1Ygfh+LArutSW6udwPN6rquzEkY4kJPilaIe6ymD5y
rzzYyqhtts2v47x7MLVTDCvJfzQ8FpwvkJtSZjJnblh3YPb62eJy8NF7juZKb0Vl4x1zQwt3frnR
dm7nVa4VswP/myfM68FDem+YwTiMHEgxeGjj3GpbcEsbA1RSvSlWp8JpcBhzbiVpTFuaJ719Obmm
as1BhNUK+cWLZHChqetIwINetJShskm276pdVBpPjenOT9WrqcKWfiv+Uc5FRQ0uzBRJsGcLxBXq
xO4qBgQaUn0Cduwy+dZthbkyP/N2iRQsTHvVNgL57FCzrdy3huEEAuVm8Nreln76az8/5MajbuTg
wXAWvIZFo8qCBOyjslKc+toGLpskwHAsRny4HyXmlX73I8OLIliLHer+ZNrU+BmFRdimFWlVfYhv
efsagU/1nt06QYCncl9O5PXFvc7x0Q7lLYU52ZAoBpDMruXGMGQZYRxe236CL9kdHlVVptiPZHWc
ePY5se/t2n9UcxXLOF3UDEL2k0hGK0U3gaLETVIxWgTYlvxJ4LvUUVgsCjwEKivxuei8xAarQdbU
7hV3xuqYekj3RFpUbHgO9TLJYBsiUavpV6vd2zUr9WdhMCUKiCgxP1b71aj0RB9UviBdcq0WH0BT
HdmGotWz4o+CPv3ybZ6CvcyBUx3A97kU4NXSl/MWPlA6KV5pXoklWD9nhZXyYXaCWwDeycHsiqhy
+UwY1CR+Mj3UbNFTmA0GSHMXwYiVdm7BuiOomELTu5b7fXl2BLXTX5HnqkStqUHyE+qrfGaS51lg
sdbPOluiuBtOlpTC8QWCw+hXWTK7cjBj5NnM1p4ze7uMZ2UFfwFXxsvdQK5LTSykoQcqI3ASH8/P
FyR1Jakuz1clRLf0/BDtkrGp+6FYwlprSWLeMIHmY29seoaLceHahn5vd56cFzzbJfxzPoJgX+2G
jUtM1WhQN12qy0yiwjbuGrKEkw9YPG09W0XI6NqRBzUtU0t1DdC+1Dacj4IVmZZ23cxhAT918PUV
BB5D8E+nP+OgVAeCB/2mLXnF+KowK2/sKJWKfJTTQ1iPCBUlZe+oEzEFJIBBj/232Z5dMa3FawUB
d8uMFjsUp2X57Q7S+Ya5gAjIH+4QGLgVe4LuGNwhwoClWGNUjcO9XpkNKdVXT2mG1Qc05tjnebRn
WdWGCDizoUJZ64JTvs3Mt5b5iRkdT4hVYN2wUAc3n1JIEPhjm35xlMN9Wj5gXLP7uBXbnZRhHK9q
QvUFMkLvuWDOyKlMxYpgc5lecYtGXOGKgQFQNBjLMrDYui4h4c/A5WOpDF8+zOIvZSufJJF0dETP
vFeoVuMdnx8vXczRT6X3kAxBqKqUfFgCGw/HjnrpZt3FcEzIsKqJbjBH9qwFifUI9Ci7y+eFTnA8
64dScUIYnRILnVL8/oNIPQp4M8aBpUjrUKcjxiVmgti9/GE4G3u/rhp5JyVbBJpqll0tjKZpJDPr
o8flwGTemgNR5VOlUO5OjcrWx970OVc6Zj8RSlZqzJQn2C2IH+xUayQWyM+8ydMyovOMzNzPCFdk
Ojn/shb+hqyQyNjhrwqx03s+aNqcHNtarkxbU/dcLDPbVbWi7fN0JJamTZ3JFXzuP1/C4N14UDI8
tLtJgG+gVZjbu38xeSJQ2pIEZ53cN7qK+PwBuSSS7sD50eaxS4YXqsqGREiX52DKPO/wFW8pZKpe
VZy0g+MD/Rbtxwj4iYYlgaqow7Ul/rhVlsCAVoO3OUBu1hK4BbownxQX69qf1Wx3B4nOvudgAw72
ZD1QlX2jZnPnbMvPkubIsqG3L+IfcOCQSoJcAY68KSJSRqp+jbdVH+5IfimldfoiEm2KKl7tBClf
PzWq0t5TNjK8p+cAvY8XfwGtb7u+Syr156JoDcEg35djIKlz7NljQyPGl5crQH7aYJfEIUIrxUaA
t21OvqDk1F26wqX2+sz6KWkat7Y6M3Krnkacb8Ob9h3I21R7B87y3tSbK1GONAg6fz2hUDYE8ctI
LKtlQ5BCoqjAlVqAb/isBw4mttTimISswQEB6rDeuvpGN/Z/IFLAOVontBRkd0F47b83oFtKJbHI
aFUrQZw7M0V8lARVWbS5A85PVOXi6J6kvRzZm7eYdd9kMXMmeGZmkwmp3v1kyKnBPIR3CvYkFwzZ
IzQXWUM0FKuQRpobQbgPmUBOv2ug+N2tvIaO6EfUfna6b11paGY+UAhZNOgC07l7c39yayxyy4OE
bXJCkWq5gJzlbVWwNt/MOeRlZxMQujd8s3g8to7qxaeolHiOzv1sXPgGRC27F3JWx3IrHr8x3SHB
MhVF52UxfblE+kVNHdhBKAdmjfS8CeL0XSnIkIT75OObdcZLAem254XXcLP2RNiji1kFMOUCkH4F
R9kvwf7HWZmD2PIkNcR+19qqJvIOPd6vBO3pszXbHIdHE/AYJ2QdL7+14FUrrN9m3TipKu4Ual6F
mclXxy2gwvPfn9G/cWDTq4M1L6woXXg9tj302fghcmkps4il6lxQGSgvyDRSuMP3ewjE+ePoOPwq
PYk9hvr5D3HPuJgHSHfNVrcNDAX8qQzTss51jv5iAz6dlqzNai94rRAC8TUh4kh/yBXp7GOrZQHx
A9CnMj0FE8MXj/DBMMDBqZJZzx/414E9RSblPdFqqCSp44igC65jYeVpjD8inkphKWd+pj2Ia3h2
HPrFyG3g+RKKF6TJ7TWeYyKif3+pggxit6bi78NOoiJ2P9YDYPMkd5zqD0qw90s8THisacRGSmhL
JyDDpljTa1Q1swHXLNBhfIs8XgaCAhONg5rA0i8mYJ5dx7DahE8XSIQP0FggKei6/GI88pIS6kXb
RjkKk7ucKbH24H3J/yYES/rNPvIKEsraIqNZXo8xk4A3UjeKeegt+ugfA8o7gCiEA57m76aEqjf0
8PwlLtlA+7kyMazwTRSG57zBDx7GgLCdMjq0c/aDDNkjLSP3xABMb6uWgDBpIgKtz3UbnKlNyQQ4
W28hjbpEPFv8PJMwClsS6KDutxPhmizgQwPDSg89Gau3wA421IO8Yiw4MjqYw33YK0gSRBFIOH/r
y6d+i0/gUtN7TK4PUEFJga+sVQ5U4ZIGWZJqOu7ZGtrrA2rfZZPKf1wLb5YirQQhUSHrNc1evImu
GRq2BbV74fExsZ6etv8zlwyOsPmPAnbtYrhh/TW01A4kaFiAiLfg7ie+QOGoErJcnjTnO3UvsjxP
aOo2ESgDFNjFw8QEkr6EDmhpWO7jDZCG7SdnJ8lZgEnm8RGCw26l5bfn30GIUE8BwA1QLy9ZXZAS
y4IMC7Twmduj8+A2T8A3p2ig75nfSLvwk06mhlZFYmLzi2CpuX9FhECqezBZ5CvxAXnz+VraOOri
ODwOhZLtK2A/8lhP4RD6xgVXpbXVOypkg1V5YngthPBGxc0yL4aIiz61gAIuzgoX7Pj422yEjeVH
4MBJHDVIb/OnuMyOPX5KwU2pKLhZv4HQ75vfcZ7OxvaDuVjEgOkVeWngSVE3sheDPkof8uzBOt6E
IJZRmu2S4op01IxgF+20H+HJyRzhU9YcAeccnGbpCgpgG+luQ4XLSzsvqwvNC2sFjsnKzqUwtEKo
KjZ6JenNSnpi520eIoWTY5vOdN7FWu+kT59687K8hJDD1fzSBuRe/5JDMofx+2A8lm4wqE6QagKq
4Cy8tHzVVclgGID2nMG5l3IIjQ0mQ/iTmmQE+CRF/8RxbEtmSWgytHDkm157OaM8qo1sEU+5XXtQ
9u9uPqXMfd0VhpEKawngbM1JvTcdUnN2945w3hmlAXOhsgJK9Y0JijIx3UDIsn5l5RaUTpMGaopw
dEgTTdNCMr5r8kQmaLdmMdbQH0y69JynDHXanagnqWexPaHSsy1vqdNLhbqLfg3+/GIuMZrazy9X
2GzBnfo9SZYaVoAeIoEHY4ntVaFP3etVoIPipCRvmWva/Za5RgXegOuw1wrU+qUyzVKnHuTwjcNq
Mggu3t8GQFJqdmwQNpY9+d/JF11aeiaH7Jd8euc54o9dJ2ZP0nf52T62zljfTBzM3epXOzC9fFs7
AWQ8AyPQ2G7VbYUjrfZp3TwEL0FJjnZsnrxnTG6+eyURha+uI4yVVVXGLRbiYTbT8mvcYhZ4jxQ9
gHAPJG380CQgTATEkREfPvW8SHEkoE8sThGmTUzDabc+UoDdNGcF6L6Zw5XmUJvSPGGJOKs26kN5
zYmBwiuAD0yO2GMcWak70/cnZSeeFIiwoZN9bFcsH+p5ltTYwGnB73PWtZ5s3Hyvl76KUvAd1nQd
9fJu91mHBhIeaW+bgT43H19VunjufRkZVsohCZIiqf9WmXdKRhmlgahKqQNJR/SPMpvPII6X5HkY
h2JBy8DLtKUKaN6J63VY/N/UpKM3HlpUcTdqYF+knfQ4sJ198AiWVN79OIi/Q3QUUad65oosnlyQ
LUV4PgOFnnNpmR4nqQw1OuyLhj3j2+LOuGtcYBUjiJ2nwLgfuckxN5Z9LAbgChN2s4/OiWCLlSeC
h34Zq0uDpsfYIZT2MOiDl/keLQM/T2BDUjL/z7wzppG8DdqoxCz46meJwsbPnCfnMW5GAFpDGhth
wSjNzSxSQd86ed5W5ok5EGplDiA3EvI4ezJncSs+FeJGBxzmIPCivvXCo8sw/AhJ7oJkU/LTKcFb
qiyjMLXra4+9NQtnhcU1QP1DK7xi5JKkucBmgFShdL6CP+3/CcbQG6USjTjmSXZu8Z8xN98CcXmr
zxF3Eroz/YUYkxjrx4D9OZ60dwgG/qqaCRrQ9DrnlfIO3Rs1KEtRYnO3p6nwDe+Aq/BsuQ0PRAHN
dSBXc9RT3a/hbEZ1S1CqcYgfageORYDuUosy1k+PGCMiWPrWqwlq5FSOMrzPJVpuOq4/FGUBMUUM
DyjuAc5xJgrg2yuVwW4KilzxAL1yBVw1yHMbVLQT4IEtCiHRuc93LISmehT8/Fx8Z5Dia9/3FboU
4rO7EaCUeuGa/kx/xVELCX2VmaYDLQT5L0iUMQlXnEvANecS39jVFPItTa9XBP4drbtb/acEp8Re
OKHo1ISuY7Te89goq3pB3c9gR5bvZtYEVgyQBXq4rG5bTbbFHVSeNWAo6p9aAg24kN4CIz6e3ICz
qa2h6pCME1epBWCWCGNwVAPivTdt49srtIrVmg6mFE8FgzhgXT+INFToeOsxPVYhIMGOUSUbDbvN
P3aK5pYupDATHLXW+8Ft0MTNKFDWCDPNy5M+fZo33vQf2J1+hnrM6cDmcnuHCpKONlvQkKehi723
x6HlPud6yy6D2zpdTwzdCSOW+OIKLSs2j2yjy9rXO7mGuT8Gx+Ek2Na0VBJvgOCrcjSm+KaO+rLc
9Xo8BfcTCxwlhobDSmHae+gQytzvBzf0DudPP+6sF/Jp3MgWZc/KeunWiWwgSwtXPeyvt4caeWO2
3exk2qesCeZLnUTteB6kr+y2SbdvcneW7BjerW1Id7Yr8Sfv9UIETiOwl6t1+38wu4GLyTr4QW0W
2aB0pZ+A40pRXwLkwgbOQ2pV6TMXAn5TpD+LMZ9cUcyjZgp00ABDcP2QNi7+QsCFhpivQTexzPh5
rIgKar17ZDDXc0YPS1ZWQHWhhtkNUom9r3PEfn6oK4oPUg6RltCakYCwBAB4DN4S6KbuqUAmVIaJ
CJZoIHDxWsfJnN2MJZrlghQPMzKXPjHRbvrdX7kTPhSRFQwNM0zRcQTMY69L9Tq60+GsRjzGtAz0
Sq3xVWr6OmbLbPbqHJ7g/f2URygnFZlbfjJbEW2OB89nX43qp5eiyXPKH81qMiWYMb7xxu0fv8Gn
FbHmFqAxRkp+s3tO+0xWViFp/PoMseZa+96mKwApX93bMtVz1Z9QiNXuPSttzrLcwcqsPW1G4Krd
lwGyJ1gp+R17lpOjyzKq/bLZwnCElq9g0j6j8lt6Yi0zfNNaqCAznjCbWHzi7k5iTo6dcSSmQYCk
rNui4d73db8A85sGfWlK8NSTdl/pv3Y0SKrxgyXhRZZkqNQ7bNMxu7CsrnjZtx/59KdN8rXFFH9R
f7tux19E3YmXoOj3eTAB3smHudYnDdUYuBkoC/0/98WVNIT2Qg+sBtFjgTE7nT2iKjJZA+G+055K
LIVRCj2NQdulKUBfxWb9AswG1pGoDB4oqcGYVCJ9ZQ9bEo4vAqBye2nqzm528jhU09aUajuvIVzK
Tq9nBwlowEiD0G9S2ykcmx5QnIW0JVfaj7andX0ApHUsCiygYLTt//La5EkNm/xsh0ty9g49L5nQ
KQAHeoqmj8aHFWzMHP8zNnH9jIG7/W3QCr4upLYio3HorTCSQdYIvujChLR+tWtMd40Q3AqGnTtS
CSIphK04OT0S/3zAtvEXraZETvbamNG3n4+kIJs95nZ0msEDwJ8NdSBu7yUwdJrlpq5QLQc1guMq
c/bunMYseaaONW3xS06oZVE+bzcv5l2Z4GeGFL1s5iWfa/2aCcLQJ+c8DEbT0Q2aOtbwED1ZYrWT
15kw1VSx50zoEhPvlwqL0Nah57mk2zN3J4y3afirDaiHqag3Jd1epBj7puv5kMvx7wEKIbYbaTFa
ftuWRq8LB9SnxuT4rtv4mnzNBOKDsFd6sNy2K3+VFCMgXTaORNm+FhpAD7GU/pS+ctkMSV+a9B0G
oMQDzt3mxbrqvYQEUQlOMbBlkqd/BmgXlsu+49s4EHPFH+29YT0YG3QBd8nBOeTtvZj7wLV5Sb8r
aX/cFG/YwSyQBpnEmINgJBpGh5xa4+npHZdlEdXWuzoUEBaj6Znq8IlfIvYqFPN4zRiPVpUBAqbk
7tOisN6A+41FrAX2SzmY9XOeNVeoUD2O2f3sy2ywXclPuTg9lZez7N+L6sMyy0jBjL52pYTuG4oy
zrtKgL/BqgTsMQo3grSWSMCNbS5CN56J0dC4qDjWLoSVww5Gkv9ScTzJDrna1eF4ynGpBYwnrD22
9X+IoiQc0pSMD4SP03Agae2cBkQSjHlr648jsstIYclZ5s9a84Su2uVh+MufFQGuZTSQn1GF3uZo
VPv9Tzw3bVLj80kZs+wL2yJz4UIGPZNMyZluWoZhTRxlz2R/8PGAN4XeUVH4GtMsD5R7ELYUIHdf
wq+AQrWu9SHYbo0hKbRZTUbNIlXb0qfAjq5mJuYjzDZTrj9qScbJasIt/6xn21ITuDScmB8wLedF
q6TEq9Fu7umPVJmvl5cPbr79FP+ek25yor8qUT9oDcca719LJFIoa4CF4dv1RG2ckvqP+485Jleb
+do7zy68iCsfcomhWGqgotDYrJVnvCXw621l0BL/m9L2qAOKBVAn27w9sN44aUioxqS5qM6gxH09
2K+9/biVPAVqBtbESY/RJKVkMN8mLCbpYqf3TKMl8BMzRctSBWhYPCQgq2g4uw2DBufc4mEZw3tM
YvXVggxH2VuIMiqNnqYrJSGuuHOqxU3QTnwqcWcaTWaDc1Ec/H/uxH1nYPcXRPStEHFHXEv716wN
l6dl4sXFi715UDLI3EQK7mwZnIBl8BUvU66Emc6iCTwCSQqGTCblOZFuQN8CRlaiA6+O8T8HsFrY
4DejO1qTpTJn51k3cQ+yzzKjnvtlryaDBfixnxidog1i3E7iryQ6VwZz5BsIOXpL0GwSCGcFTOjY
Xx+sd1s6pidcpDEie/GXui9MLNOcEoiS4zYI9JyTDZbehbjXFEAZ2OKTaKwURRdveRyClhN42MiO
udXi3QFBzcP04Ad5ZNYYdrEwPT+h22Dobi48NHFx5GuiISwxhampqPDpCAevQeoN9j2K8Ansln0p
3wgoz5Lkntk+9bU8udJDfQE1QFXVIA3qT3kf/7yGYJiOsfSZPriYaomtynY7kWZIjQ3sepckzpDx
N605x+cITquWyqAlZGV3OQwZu6+zqt0k9iJ/oSQBPeanyFpwoyErlwQS8OcTm26LG62eMJeDZElX
aOSuumX+m4AfGfrNPwZUNFQ6Cm6X+ZCMVa8vWUsoaZny7n+YSO47dQ6vtTo6NDP8QFYHpXjwO34K
ZSYL0YJZhXwcHA8cjUeQ3RwMMn0pDRitENHLpAwaqsii/1RJ/TV7c2U1SoirALxLhdlRQcG/ULeS
P1JkIp1DwYZLdIBtxw4g9mJbRwseEh7DasG9y2WbcCMT1+aTt4JUivAdSFW2JDNW4BQGqpLLtYDf
9daPT4GfdZkT8ACkDFG4j6VbtekCk7d7wuTfL/+ahWp4i4s/27w9QGrk2Dt54STNS/ThJOx+CztQ
0GnkSVaztuaMBYp7TwXJStNhFGvuOjqTNbHdgEV0orC7bPfWLnV3Bf7l6QzQmFxLiC8eCfCP8iVa
4TQGSZ+PrrVYgS9Zh1qkt+cbZFTW7diQ7dC0+8cThRbZrvL7D+Ryd6NY66X/iia4Et7Q/omZx928
oXFhnhLK1MzmI8I16FVsYr5Xg06Ng6sTOTL0obuATpLl0vHG9qLSb/mlbF0wY6hsgBk2tLAvsCAC
ez8MYlMot7qTVsCzLVmpeNbpCbQEA2hn3w7Fx53JPmiWrUoT/raoCYBAbDmIo//603GHcsvNgJdF
PZ3c/i/qd+BNc12VLYWNAEQVRg5wRCz6M4jTpnvA171MXfr0NwPEgGLztAE8MuWQw2PWDPch6lfi
zWp4xOdLNLmuhE698JkpatPawhUuvxBGf78Z1kh9eaG6xTFasNZ2ZmSXakB5Zf765nQUkm4Njidr
INdYr7aBihdje6fH/egxcmfEuo1MPZvhUTtB6PLMAVtZzB8In3bEtTg37tbLtsOSkRCvInVf9+x4
6B5oUpmzlvi/AEMBIQFTmct4WUHaRiTcYPJSFz2286Z7CxtVI9lgRzuI6Em4I5jGL5wsU3MPuIHx
pyT++u9PYxrFww6rPzIUyZo8L5eRnhcJSU0r/+kHtGX1xlpdeiz4+MJPFz/1+S2IDWn68s+3D+b4
8u+AGYon848YSeRTHctdEhlovavQlYeAmlphHvLxvt40AfURy5Yv0mQcXPRuZgPyMBVip63Ynaso
72ld9Fk96uRVwoPUl2/6tst5iE6TVKBr+cnIKW/bXmVZmegC7OfZcORaIv7t/11cdDWbr77fMN3F
CGYvcOUFG4qzkaRFc1ONLhr95rCXWF6HmagbqwIN0R4QhAH4SwDOiHq7tPx0gcYihmDQUfWq4aUg
UT9yuM0I5W59rDQIgbYCv3nt0CENqW37V6n+GzzccT5S75AOTX+fCRQw1+hrJpMIu/hXZD1qZHPE
ufUQ8vW9fchQzY7BfqVN74O6uJpQsJrnj6Oi428gdw9jzuc94Kaju9QpQQJqZFLEI6wHxdO0vWSi
nlqMGSdGDIQcwIB6QtNHpTynPF564ydJA57H1B3jA4tCmfOcPO08fE7QyB8ASuFHk3ao49M8vpCa
PMYgDneiYQ78lVT8QRVt6VrhFI5JAz/6MmLSYfRjWCLfgD70/9yNZznUGukt0Jv1temYZ815Hd5x
l90lPdjt1bJvdt75KKIo/lzIYsbG1puc+wRP30ajte5oCGRZXwzvxp8KW/jvuyeI3mfT/MPDyCc3
YbpR9Jz0LZWhlJ5rsIKFPkBw91UCqslqd37Z4j9ETmOxDg++db+5VcQrIBIsJmQeZb8Zndt1vcD4
VBKznM0L+JyyqQwuPDf/8b3/ystCd6Dt41aAhEl/aNsjdCdkKHBYxCymzwL3FN7IHXoCp7SAbHjE
G2STzN3UBMxQJ9lE7R5WgdO53iVpVbMKD4kDFvzieK+LftfV5FQQayXONTE7wFxJSeMFITJyvFRh
rgCs7drB2LfTjeGMZUBJfbEztWJPDv2QnVkxexUf6mJqzs3Uw4Qf9RlksQIrHj8epxtL5jtpn9DR
aQh7saAzQpINIZaVTanVHXd3t1Q5e4Ddo3niyB7Y163M4L8z4XT9dyDG5w4Eyq9+qc0yqK5voLF1
9opNIbpyB56CcVqqdVrVnfBoH6P9QLzcNeN96z7kra1XeI6qWbs5dLYyrY46QCzMWWDc/RdANxFA
pfWNZPonBn8llIHzWkDuIR6eXCO3S2TckaQKjOcfOBpl2sMHJtoedmNNHSX+uSxU0CroYzy2DMMz
HJbMsi9iMnWnNdpifUrVOv4ZiyCBbviZaobYyDbJTmVRPJc8Uj+3VpTVJY3K6g+IsVveiwiOuI2Z
l5PD9Oy9K+Mj4CIRXYwe1X2CPIK+n2wBoq6P8OSRBXeqq/EhQUdclBUIjUizywHAcy3KCuToeAwN
HlF8nlezWu2O93ljbZJryqbFExcGkmkEHD9r2u3LCCmd1KoKofEaUy88Rf3pJM35f2eZSMCwGmaX
SoTwlZDV7vPquHjHjt2HOdMA88aUGVZRW1AdknJvcillDmnny5s71vifBIW0kLkOnYzEEUZm47s2
/iL8i9A9sRKzTzg9VPPf9TiHhJSAB5ya/ksfiVG7qTJd8K6LMW0Ou2xc1YM4sgYNlZA6AZk18vKQ
S3mpPCEdnpMaRjR3yJZ7RL3coIKx8HxYxT4ILzPiLLXPePIQXRUvHMJE1nRcrzad3AbZ7DXS6/2X
Hn6fn3wiWlUGRUvQbTWYCVLs56WzZFW64x14GlE6Weolh56uF67mwj9OkHqYwwuA5y3026RgzDPq
e0xtsE7vzZ/jc/8S7Idb3yfUqKJJXlsuTbAd9eIIeDmfRXSdsfX2KG4EoR6CJTxxmQ0RB7r+o21H
wplo/UoXUPRG//7V4pou0JRRzVDk5j2S3nhk6UYPczIutvmM6fqRKJS0PCM00Lq4CEoGXxuiu+0Z
PwS7L3A74Wy86CK+3kKAm2o+CN5Di+3JweTdHPwvjrawFPGu7So55uiy3cyISAtVz2qBIePveZKy
MmkPGQK7Zj5MB8a+cMO+dnwHfogXslh9SjEoblAJGn7cqtUBOHoRDkYjF7GMqNOteTlrl2HYR/OW
ckIP4QYavJiwv1LLRRqO1FmN+2Y42Mpe5irMIu+oyyd6lBerPM6yisGJEJPMZdkyvX8n3p1KP4a0
BP+5LWg69nUHZouRklSOvNMUfLBf2G+zU+2vaNZi7KicTTI2DpdDOjJ//vV30rQ00clDE94sB5Ut
CA6+IyRwePhwhQ8aOt4BEpR7V0qus1F4t2XFzzA9V4tUTlfxyy5eOsWBnn5gra2VHEOVG+nrXEHJ
MaqFP6cwyUHWmIlMw5Fm7hGSmFhPfi4BPnPF24uivz22fnh8QfLU7TG0vQZvtOIFrl3SzY1YdL0R
4RKVx9nHXXHrDx6k2w5M5axEhkDK7DqqfyeJlDraWxx1eUIs/A3wF2BFnZdO91UaFM5k9PX3K8c3
z1fWiUwfqmI277kSyUMGIFocksN8WeMsCCZHOcKXLydvCuLivBzMQYhHdbPDMK+0Y7PYIyRxK+oc
AIoBQEJ4/kWmDIfkb8lMA6IYVrt/CpP7rtnwYs+S++iBWh/Lg5uXwpkuAkxj8wHRxfPn3QkZhTVg
SxgzrXjqwIRzHRBPL8sMEQ+GEa7D7xSEWIbjmRR5+qAFTNgOuTy88hDlY0fc5Q5zUWjAhJuSmYuB
1eWXzD1XoH6t5XZOlWnAWW6X2p/CRnHfF2mf1TCwMC9Ip8GJYUYTxpzrqKktXdwdQpsCCW76oKwz
n1nIunBVzEnpLHnmXpfPDaN9dQ5IGlWZM/xZDpF9GeOe0JZL85WdAdvIYd0w3POtm9p0Q0v6sdKC
fZXJGYeD3VX6yOziqz3EiTETOE6mG6AUrD2S4lhfFpehB0Y/JV5uPAZz69kYS2vA+oJC9LdsgrGF
68voI6ZLT0dEi5ffH7otH+hOA7/u1eC4oJ3iJkCwycZYEC5ue9qUkvtJP1ni5pe9q2MZBleObDe+
Zdg//Q7m3wxCjWnmNuy8ywYyqYYqWr6HV+EuQGqyG65RBQ4hXqGSPgd8AjyuyFl0qow/MqAkTYfq
8MXB9EYp4/5nvwzpJs2W75rBd0hB6/Z4J/GiACTOnAC3zSjj0ltfRxmlbjGH0EUnNa/gb50fiU3N
soK1yVaLRINuOa7bmD/QvvNU4UlMa25uR0sg2q439GtBRMIZWvrIIVXuaXHiVobb6BtEH/EWKufA
prZ9cVdnPjDgEOhDkEWr0rAVt3yTLhexd+ambkWeRSJZLrFA4Pmxyz2RPGqIx2Z0NWISk3+3US23
7jWlPXqXg42w2J9hzLPOwogp/WsbWyqoKvspI6BNuns2B3P54u6MBMse6IFs6gN04+udfg1v/rIp
gp/BxFvCBXS6IEvu0gjwf+g2BQrl3WODInyFnKcXK/wzXRKuTnhg+svOwwNms9r4mPpFh2YP9Aic
0K/9sZVc+FISy0sLVrqvfaikT+VrqFvbax8vympa2miTK9qQAVZq0ekruWM95Z6ljasCksAX455Y
hiy8IKtXBQ8EnS5ASWaFbgk3Hjm/Utv2Y/xi7RIfxZAZ3AjidzGl920Cz8pA0w24SNloDGYbtdjQ
B+TW0othWcfZbCszyTGcJVUf/PpVoKF13C1R73gS8bO3zRrFYfjRyw/A7kjAe8PjXGDGXlovFmuL
rnaiyPCwduhEtFvCmONB73kmxOZ7TXGWGMisefyoTz7bdu6rCKrfN/KbGS1f0nQkou6QhKdpOdvH
yaSWQZIGjxBme3h2rk2wjTQdriQzOOMkGb3YRYd9rsbf4vrzf1WPMXD6R4s4Y08LEcC3V/sdANiN
IWfaEC4XpLrDwQCHbvD0MckgPhZcarAfyCndws7AMHl8L8DR24MK53kQETOghM3lvk3K2YpRkDfT
8LbYBP092u+djUUi35fF4aig/b0aNMu/aBKwNEjRzpL4yGRYSBers1HSTo6YG0XgySpwhG3dcvsH
al4qEgwWWuTHxiAXv1LgreUS+GCOJwk7UXMTUSht0MWX5Mm7grpNhOs/W4POHeV7jAmYKd67scN+
EuSdTTeL20SaHPK5bOuJLQD9hgRwv2xIandd3Q3mzN9rEZUOWcQ8ukGpQ3PkvXFyHJM394aBeG2M
H/SrBxE7m0ZfnrH9yIhNrfeqz1kqbdaSKys5j0kzLujuKoP9henucBWBcjJ+0QZAryB5yKuc0kNR
pTIMEBunsdZLzK3cTL5iSJEou7FhRdCzKxXGTNJG9/3Ka+5EgYtX7nxXOkwZpasE4ouxCV0QJ6Wc
oKlL9InaB+Ihr2vLAhcL6kBHwP0/ayruZFVzNJyBgdeXJcV8YPUGiHmnz1eoIW9uW6mn6uT/+IWc
aDE3Vf/KgGEGCnY8+kXepyxI7aztKOBOn1DhyjiwG2GXgPtsZbu0rYbZ5pnpEHOHC/Up0UWl3WSv
GezNvcskqaXkfawX8hsf7QIKzso1cnSvFuym8dPdVGPs7zhzZMGqnxzq0balOL9068ehV2MGoef3
FRcwE6T4qtJ0WW8WxwULuMfr8dyZgDdI7mXQ2RMg/rV299doeVNHEcbvIgBd8cNI5jTqRgpFsnXW
NB/7Vr3YA+Mv0UGQqgSgpg6gkWaLzXMapOq7iwnXphMA9Ns5li041dTk6LvrxFnPjW+Z0WW2Bp44
YLRz9naFskgON+00hKxUro2by86ePNPHwI9guGynmav2X+7vgKo1tS1FvrO3T0yUJImHhk1knyMq
1km5kSsuDZBA6HVkARtCYB+QQU/oIe7fC6b+Xv+aKfW8bJyIFqmZwujww7NjWmLcfwayCsLBQb5Y
ADFfDzXM/9E0eW2bgB4gEsdVxOsD0oI6Y5deWrS22QuH/qRmT83ekD8cgsg2WjLgrSzjx5HFWKHa
knRMBBcNrkABG8qsNbgHjifSNH6C2iWeUJYOQYNkM0WyI9kyPzQzXe/aS7VEF6U7BVHmnCUWPqFp
eq1YRq7314Jyx5q49/GXcbTEdcJd5s0zGaCU1rfx+Xk+21sPFIV87hreeKOKPG8d62KJhdzBfc0+
SQ9zfGBr46d5uzMg2vbUeGkBV7BgsR+Ggxzrq4zeySwxJrTRn3opRzrv59DxwiVXfx58lAZeMmDq
RpOmr+m5LQGDOnUbTJuCtM5FULodhqPQUQoloIsunqMQyDl3vd+gI8GnULlqubwyls0CmsoAmV2V
MxdHGymgf3/vjHAS/0KvE9uh6zo1JB40cA1Cz4VGn9SVodNOB34tppkTC55IFv9D0Pdstd7P4orM
yKBWxgKRk4zrD8Pi1ZuV6denl3qqOEJ7h+WDaqZhQ36Cg9YAYWsiJELAOkq77Ygp3ExjiA14wtWO
tTAzV+CT5X+zQv3zuLJ12OZ23ICXm1TGcPT1yVjMoCIXbu6t8GCaCOpPUpnyk5Q74oqepyNAjej4
8sKIwO8QbfWmcYQ62DnYsc6kzhuzustvsyhKnmISGkFhOg19FG6dv6e1BMVm20uGLRyme0mzEFBi
31/MNq+EFyvX92o+r5aySHKpGb4fc+jnqNDJyHCIT5cxEa30ckP08VMprCpyni0+PIRML3yl4T8r
xFTgl65abSOjPLBZkGv2U38uBXIaBjytbLhSbnqXW0Ef/5l95Q+QKxIk0X0bvDomWk44GVK/G5YK
FXq4DLE3zIfqI21JrYlgLa2ZWkSENrePhEvj7KgWQ03EaxLq0gzKCm7m8yrkLu36Bzj/+5SpoK9w
b5lYPEWfi0TmuTSkHYRZgvOlYkZ+cIqS4JULnPJ92GnKzJ7FAO9r4kysjw3xi/UmvDHqaH9ujS7J
APt8B7oCnXSiNL17LsXtMoo8Irs/abpT6/60NJMEWlTTAsBzVUT+zjrvHF3mwPARf/l+DRSQ7qGV
gJJbm7Qd70bp3zAyutgvB3MeaUW1K4S5D4bFKoeAqvibbx3dU8G3Mi123bMtXV79vD6dtAVwW0rQ
Glk3SvF5y/0PNBHhSAxrjcE7R1wIzLRL+oBTzDMVugw/Hc5YG71lCZnackXxc2dBIKdHFiAaWqyt
siEZjSrzNSkJf+AB/dSzq8U4Ku3/BSzaC4+sE1DlLRqFU3YPkkZqaV16Sig/6nUctMl48U4GQq47
KbXWt7yW7NFatVUwmt5FUu+ol9oL1vfRo2Q1rpKrf6T/Kqjm+TMJISgp4fFD/fM27Q2NH/zWLvZk
mbg2y/vESvHD/SVQKxV2440xu+KCbmvaZX/pcqcpJbANUHYGDGWYj0WpRyV/tf5VAkCTOaBwTysU
iavNhBBZ1Q3ynzwpJocMbGmWIedb99xMiVMLQFn7RYQWH3jGkP0BP/CNyozHJaiASE5oev1cuyUv
/cr3yuD3SK7IZ1qz82W/8hFypfeYs48kLNEwNADDhyujjdkcI+3Q45P9J+J6n6GNzSBf1WRuNFyE
3P0oJg4fkUotAy8567L6eRYg6rq3MOkwa/UBl/P3dnqxIo/eUJrDKuWe392gmxz0eaBQNwugtLWf
19ncqfw/4zctNoeKmgV4cyiy/NmM+iP1DXNSZFNV9IEY0cGeiKiQ9j9gbI/nooJzmyQcb5St2sSi
S0w2m70RI68uA7k/k52HFXESj2A+XXyBfvbsFvyCKaxMspk0GyXtHUlBpeaDT7f/+KrvmbmfKE7k
D9uxOt6K5TrmixEwRUPxX1o41i8+azUtWxtcDb9bzBKfeMo0EKjsx4ZTngtiAn3qvcRH2/WimEgx
6r0/gtyCM3XnQTYgZkqN2TeVwXgM6e8v4uTVl2KSY8mCewfBYoUN4/D8kI1wkOxYQD50x0PCC5S2
po2K3JHtr6oP0OBxp6gpAVlK5l9AZcUUh/Jg8Vle3MUH2X0eI5a65+ysFn5ndxjOgUtrqAqgFcYN
ZzHJsYUuCsyAzonYjntFgPVohpDVhMetB0YwtvgRp25BPV7cTUsou24bUcjQd/5PvjAJ/9eNZ5aj
/n3ZWISfrckHjkxTh6d8XBovXa6eELnVe+8fnYK8noNIve3ITEc/hSyb8WCmePCBLpYxA4DKsIZE
n2Mcx2m0hlgAL4Ygbyj0rLHokVW5ohxshDg3tgl6lv5/T29B+5zlzCAgnrZh5knPdcLetKrtyAM2
rWNkXPROHvVNV+920/+lixrHL1JQ8S0BK5L7bOdDJt43Texfat8XI31885BfNkWHswZfrsjmvMZk
f1szW5Njp7Ox4EHltiTxFPDamggDZqzL0Pe/wtwDr64YR7WVcpOETbb4S52uSIB//006NKrF22zR
l3J/J9Ls2eOj6SjE/geNSUs9OvtU3OLR+1+qNbJruJsTp4oMaK7sJCe5RizpDJIJN0X0+nVqdwrx
FI6QAeserh4lKHFJ63nKjBBP5NGJ5xsCFF/CqKvXBHlt3QVL7dVZJP+vw8zs0+2y1bm8X4I7Hshh
C0MOs/terCnhOiD29rITpKlt373Zl+4Np109FT+ynem7mUa+MZ7UGWeUjgPSNmw1ZnEBIsF4glUw
b08TCjcT4Sesb8E2F5qrPBf+VLcPuYS3Abrclu1DZhz0c6eKd91p9+dRJJYRgWQCBtMr3Gzir/lr
b+kLDt+DslPtQDP2VVPXZnCDLJPfF29dUyp5kWpUoE8+mf+9v/LcuiyS/YpNZUNBoCJxrSSrVz5+
wfpxvzu1eGx71JfaKRf7EPmiA7Qn11/ADolGkGzdsVXqxx/zhznSN1DUWOBUDdCSNpvi9WGCINtW
Om0JOBROeSZfvsY55+c2hkkQbNJC+YJEvHNs3JX2BTagPuqyyCE6mfySGejmiGaSznr0lrx28NPP
5pe9E5jOKDf5ldyyKtjY8ZgGXcPnYQV2gQD7haX1+wLWRQZ0Y8yLZvZZ4WsZODoSnQMrkOb0cgN9
XnhCVWnX0JswcOj/cnjCTUjBlBxwhiIvSSgwTbnl8duKze/cGsMoesYLgRVChYgkc8DcLADpUZzY
e88R+tc7vAzOGPGdBqiQ46FoOiJ+mBkBZUFktmE9AsCBtUTiRlbauuUhlpkVsMw5l6fX5SXp9nJl
nmG2fXDYu2M+CL6TifAKwl15mS2WlAid0frpg7fYYgAkDjTn1eHZswqER8LcAhXP0NvsKOQ+EDzS
GKTQ5cuUxO9TaMZyFSHUtzN17/elznRz0RxFPv5KzVZ9ZNI1Pt34utd8BpZv41ehL9BbMcHF8fIa
ZQ2TpFaWC4wwErn3Du5TpW67x5GmvgMeBPE7snO1UORk4SeuoMdbRE+Z7pQvJgF7NxugVTDByDNk
noc5Ke3eTg93Ie9G09L22elD+y+ENTLpaF71AZCnCur7ynE0ruQDPBZho69L0k4Hr4wrQZjMLzK+
JX+S+uHnUZMmkJ+h8JD4YSa33IGrgB5IDShqWFD9EztwGAu8H5i6gdcS5DSE2tLebGV3S9twsyBo
U0kbr0eVbNxwq6S7pMIOLIcr3Ck6v5YrTI0FnoXtcrigMC+Q++OPCJUcwUdXwLLmB3QgNw//lp8y
35bWrL0jm4friqwpScc6vpI1k0rlDlRlbCIfe8NugxEn23Xx/b39iOafSOrAgQtcNaWUP9H63Z+a
gKLwMwOPRSbsqRBCqDWlE4CKPP5duXh45xSElpnEJMUBVqa9yy+6WtPFY58bmbQ16AmdPnFwsA5s
8sitaUggPZ5aqCoMBA3fDPKpPgvubPrtVcvSDjpECT+gOiflqcq+Rmd+PxMP6I/AG6lLYJqULUtR
shM2jamxNcYDH/0UjFTbMP8yOIHXtkDErgPvZB01pa1b4qS+Pvvbmo0y0wZUaZqIytfSP8K/vDOF
abMnjmaRvZxID3zS8wKuUMsuhCKw1S2GH/P6WGS1pdaMfX/UJIG4SwmLSuWc1HItNT329rsUxFhi
+UV6G4gQ/mo1C3BAgPK5y7tR9GY6YRSEwmc170X0yiTyx8gnH5ScL+5wLdDCKiKUdSvurqekLZuf
UBKVfVVCh9e43oy9rIoeb6l3G8N4z7MOmafW83AqNjgLeXqpW1/xwsNRcK5GRXDA+vclOhdaf/hV
JtYAfdD9UWnA1u5HL72qVW1FsoJz29XubTQ3Vv/CAkxn1811V3htqOMvHS84q0i41Sh4bJ6Ur1RQ
dqNDlw0NrgHToxaqXS5tjWSNssLwSnbBrzx+RZ/npleO5TvTsDRIZNqWmW5doYtebnlJ1j6enMl7
D3l4L6KTL+UJkFzu9CYIx9FoewhMlnYKNpl4ewvKQaoefop3JX1FgElgfbH2Rf4SefEC/joKBoEd
GIPhCjNQXlMjyucZf8JHgy1N1u5UDF8FtyhwnLOG2z0352BRIXBJdf9LXakN10AMZa2rou+Ab+dz
1oOQY+po+56ndUHThMqsDEtetSudxsuqiePMOiRQaP/M6yElGurzlVIDIfjXIj4A7buEdjKhmRkC
kC/JpZhsHcp868XrZm8oYvTiv8esh0Z8g/NWuBtNy1+UWdQSE3Qk/1kb0dR9nYQm88MAS+0Bwe0O
AE1ZfozFdffv0NZrJdY2ITWUKWVjQaNXhTnWWCSZDg9ePuMEOq286r7IKGrihN6ok40PWMkU00F0
6M1c8TwV417MBXcIw3hD9rYdMn6p7/kYydj1cy+lNpDdZRZ92/itS1rxULRaQmKAG0fttw5zHmew
VWxKknvmtj64EC3q3CyOyfpAW/sDYtrE9Oee/Mi11RI/UUSZTcWghY+f79btYsPZC0u+3vnDz/7T
9Aw+xn58aOndOTU2JO6vZg1WDi7YRmRoNGvIsR+zpUdvFDzZF+sW7m2ata0lqrci/NoyNa53d9HA
ImvBpG4Pm/r7ajnp868gDfiuZhskYQHG7qp/MNgH4r/drJ1maMCi/NL2VbdqFZ/y6HFH4hIWgyn5
IVJVWdS4jACj1FwBQZqSIb0FF3ghQubbXw4Z8+XEoqVKhyNiHgP9H6YuifQMj9vK2tI3muZKCQCg
KQLw4Y3mRTRsjlciZ0KfEpFF+1mMcddursMt7cUyvqswC/pPS/fctGd3LG5Sgq8BSVX/1+Gwa3kH
3HiX4EsD3UJK+kJqYeJIXtfn+/PrfrGI/t+JZqqZz2EJ+Xli/KL4EzK7sUE3s3uAIMzvT8e3IKJp
UqeNdSqjMdPumIu6wrWXTcH3SEk8c1LJzXx7F+OSLkO2pxOK5GU/cNfCu0XHU00KafWzX7/bUyC3
eY5qRNbk5Dlux/X8STeTMhLZ+Or5VRyJ68Ew9yXZPNnbCqpsmi5JZDiHPSS97yKxrvs7j9gQhnix
sZ00eWaAEtLlrUn2d02s/CP8qfqXECqV9xnWhJleCJp6QT7lWJCLVdVoVdC0+E42m8qb5fO4bYQW
1xwVey3nlkNyqSXVApjBZkL/Rh4kMyVHWVGUer7s8otC/riR06NpOznbx7KSsbRgraKO5GlZcCgz
nkSz6VMDpyTCjHD74h0CoiihSB/27RO5fbFZ+vYeZvSh3e/cQtd+u49leHWa3mE5+CDQwK763ibK
aJGm8kQSPhi1psLIBVE0hCKE4OPAylRZWWJxjXGFL4dzBPipJysC+fMCkxWJ0PdpG8ICiGx+nX69
RUwW2+FYmH75b4iZ642rgIJeTKp+MQUrN+yQQKoDKmaF2ax5s0f40KdaxLj0vvh2HwtRGrT9nvDZ
35iOs250Ts9zTbR+JsQ6XwQcUVSFbXJEl2ySHO3KCIKaZUyoC4cNtq/t/YikygE664J/Wq26aVja
YaNJlGmmE/p3OBRVsX3GAh0ltiQ3W0XTM29Hsep/IA14UN+Panwlts388u+hyJpwtZ4uy1Bx4Bri
gF/W6W0Hr9UwLtDtp0vtw46Tm68DUdO/Xxc9jAsXvnQvHzpJPOMLTNVc+6aqNJ7Bp5eE0msyVJE6
V20OcS7KkV2BBKvatxXBQLyP3edCvE0PjPwHR/YZtKYFp17oeUcjn8ROYk8wbMQMEqfmAY2rEHMD
0HcVfi/lAQrv8GQry2qU7TI2u5e47M6V+MPbQ0B+QvjWHWVsfwwm0zGtHigfk8WuQN/13Iwcczxx
x77SF3TF+o6JNqK5y0hdn7feJrka/G3DxxLTILNBHiyDS+wxol4bC/4u7ffHqKS1DyoXHVkpu8y4
ZssDaQwAvAu7eUaEzW8TS4GH4on9ig+BiVlilYHDFcKiKpvApP7blxvEyyEfeadDpLz0JeQWEG4+
tZZo2wUqts1+jxeQUCSO3xsF9cp+6L2GJMSXuFlcc+Rr5ivJX5zCpUfszJNqZc+nD1a7M0VyKbOm
rXYLz8VXSxen4IKnNjL7RnoTuTvQfnNySHxy2T5k7tDfi9/1aPihlYpdqmqa8FWYmAu9s6RoUIWU
JBo6tBLHYXbk8TY9LaSN+rm8z84Op50OFSzDC/Kcow4R4wJPbz8qWzfcBeUxtoy2eDOfO0arsR3K
RA3Y/HUYK+9jkvvv0GuyCufIQmM/QryqDKgVNAiOApTL9ZFCQa1w9U/ZgnGKiQbR2DidUU31QQwH
frVOF3biEv6vCVA7zVX6j21rSgxHilHg0O87ms3c4GiKyrFSRLLH5At7s1myPazho7ckyZbgNT3M
Vb47JsfWNnQKLGACjM2ajdZA6/m1btBK4v+Nr0acDsj2byeDrY3cD8/QEIgQCesqY3hRI4OMpfrM
ZyeCWhqViF8LbDInKesJ/EiLY5RiVjuxniNIbHp/EEoym9nZtW8l6OHmsYDNl61BrsCIrX0D5QnD
P+OSuH+n7M+8aeVK1RRyFAZNZQk55DwJoYBSKATEf+15qFqh633BDGdyScmOD8xPiMCiCTI8PJvH
vSkur178seJqBoa8q5DIIoGCF4YBSgCru37+Ire1en1nsJFE+/Ze9hZoCEHHZtCAM4JHLlSzw5oa
kFVTIIWvXXyIvkzns1+ZyExtJ20u7l+BSj8ed4OGLMVwo0s0CClkw50akfk04eUsp6q32ZVdctDB
WdXAnCmxGtfBUHBrROV89qNMkIgtj3MreRJsQb2FhQZTMvhH7MndlpWWdb4FFQ9+GyQSoLgxytCD
4Kr7obHGR9jr3q9lU0iJh9DRyN7ay+S2QtKDXQofybrzyYvcs8z0UPCs9zLwSBLDPR6FyLILwMGz
3DBIat25ebKtaDJYM62jOFyIp/GFGn26wW4SNKWMGIuDHk+OWZ8RuroBzOPjtadDnbXGOV01e/ia
vJuAbJc3UyYuKLu/84O5U/Ibf7uiDWiwfr09UZJxLypT2DH8pVBX4F6O82Uvhag3dL2dItTV6BQW
euUx2bAmpbmlCKp/W8TM1kI7bZ16GmtYLQx0QstePMroQKoNMcGeGNqY4Rdm+L432q2bfssYjkjz
PmNZxS6U0k72TmJLnDeadPgPrbKp+Sql7qi9fBRKY6d9rGy8YDHiFI0fMdrQu3s+tGWv4A1Dv7cg
+t1mGAzZlkLh+RiBLmM8SnF/3e5ZIxytAp8HGugDWBXafG4t4FF7V+yN7Vck7Upab0KgVdba7T/o
lKEF9CbUzQZOvOG9xqwwAVe9uOgScWM4j/3ruml8Gs01FsXIg9DumJ78ixqdG7At5PXMrU7E++zN
BGwYTHqLimKwjpU57Lnmg6X9tSBi72knJpo4kVzyUSX0HGSE2gA8pF61uWeRtTbUq21qs2qJnsnU
VvxbcrPDZNfpMKPwu140HwWGb2w7N1h22e/2yidMioWUm1mxCcqGDNNP4YWCJAokDAbrtkpt6CRq
yC+l76lXB+/ikW6sAz6ScqSEfqcU5wBzOI1t7ciQqCGwUxaFQunt2ZCcvmLNiFynKBoiBbuqHRHj
jqn6vXB8Ob1MjmwQ9ioo3VqF0UzmrZVl+P7MysAgQO9UsLU9mN8vx49CozeBk95K/fnrZzQHlrUp
4m9RFWU/VsxCevR/jIGghocdmMa2wFwzhrL65wi8f8LcBfDJQcFB8KVJrylIFIeNzs9DW6DWkIHT
h6xVJZYT5FNgvb6EwLc/ekLGgTaADdHTlj695WGYCmn4XpouwMp389E5NCcKss8ylNZnTGpc+yKc
lIwVbtuY0eJbW97kYmF7ncsCCb+kRTtzVO/+UAL6O2EYHqgBzFm2Ry+UpIbIizybXbuQcALBkuLC
q0yNrgE1OKr685bs7KbvrFkC7DfSxvZ7mAUHv6q8vyLgIJayrdx+jQwclr7DeXGxLcghEwB87MjG
/HzJl6/qlmy7V7JUuw5mrLqhWy0VLY0dOPPEFXWAUYL4S28iuPMlg2gv6FiStZ0+KWBhfwSrIUVg
fberHKZyXnvLSGh12f9s0SdWQTk/J4+9g1V8oFvWUqxD9LCeq72tgp1Lgjss0zEtXGlNrnlyIc74
TOcmbzx7Vzvf96DJmWdN98E1cdYKRL7dRl1DSj4Sccv9KXmbC2C6tLB+ivz7vd9jIA0PsCbo1iLI
kGVCTPLaxnc+8YaAwgwMU85nZJ03ITXqYOTFJkOZxX9CpbjJhvhy0flSBexUitndyEmt6UkJccLY
mo1d79MhefbxcTULiJsjuTXs3/rQ0YrkkCLhUmIrLzeBx7yYW8OTco05AzQI8/MiJuhYQ4/snPc2
JhDbIlDLXRD4WIP26ij8COU03/P4n5zcs72H+Id85DqB8e3S6dWBMc7duK6I4+IjD8SVbgMvEtk5
dreUJnUzfT96e+32O9WDYECKRJmkNDVt2EgTuFbTHoo2xUlv3Xf1Ge8EgXV5gaRBWwIFDeLXS/jN
++INoDoApA35fRrJknV2wjgCDivn9JO0+rJ8JetZwCoh3MVYRQAv0xFiLkNByhqsSQsCi77ebghR
Nr0e2tr2+IHfANVFYPzdsNKCbj2VCxEOiagAulOlVDHNVN5MOX1g/f1tFc+xFUs0igTh2VClcww/
RtW8G/kQTh8wiuhlE+y/N4NteVo8EtqmUB4mWZg1CwIqctofvmdnJujqOWRTz0N8ajm0YXSsOsPa
RDKfCfy1YalgR6ksEKGIXRr629PQSv8XqM1jNo6uD9tS8Yc5JVC+FeAw3IX8wdkb+wt0Yl6sLkox
GVDVnanrfUd4y5hWLbEOtmGc5upaW5OUsexNuCuEEGaEgK7HFdmfMFnnCId0Amxmy86waqjDs95r
NUYVvbPJuFe1aFogvAdnlpLAd5plCEpLfzPG5SQoSC6v41eFLuyqxKPruTT3Xq0t/9eiuphC/DDG
ZIUx+/atj7/zGfEsRRVVR1DCKI0aR6Y9PdUqG0pMpupn77ExPPSoIQHGTbxjlFytp8hAipcglV8G
lGOPSTuLfyS7UwKEOaPm6C9zxbpyXQDb9qU8dG79DbAcmaXACbIWKr1Fw9nvLoDxy8AK/1jrP2C0
LdWn/BTP4artjXhaIK7StwOxa/29cSHv4j2NYTkSffgHEoUX2tvjthQNw0WVXB/Co6PR9NDTxc+u
/U+B2wygm8BU8a+hMMvQd2THCsrs6ATW6maklOOjvSJ6kgMO0sAwZQK1r+PHvK1OlMTVSfjC4/z5
xtELv/d7kCs2isKNGJGM0nMTtNR/8wyfag7OOeAAk0NsSycBLCwH7FPgiCR1Ly2ELeEB88LruMZc
/MZhh6TDwvujBf7J1/uuyZCYfe4fClCM/EoQUlbgQyGeiTA7h9ESyaPWcD1YZONlEYLbvpV5bzXJ
LKi1sxrb+N78Dii6N9IEYIKA5rx4LoeGXQRSIQgqFSPIAEfyT843ujHd7I24IoIkPJF7P5qw3/tL
8FFLg/0E8s4WDpNOvyA8gZ2ZeGP0T3c8L+4I4GvC7usiB9Xegf+QNVDC4iXOpDrSjPazsmARpoQf
7k+AbasJLGs0ELlz482HnSzorMoU0c5cfHFkl+QXaHQmQBUcbZXa8SiFje6eBSVOV1s0Gc5LXQnZ
x2OwZ9OXlQceWUghneBq3DNSiXJ0jYvOxYX4ZkI0rAKwsb/0j/IP7zLpzQvColqdWDqhZGuTb6hx
i4JzjDGPLwusPA7AeWUGGuCWQhnIGCUwd87K1YX/oCMfXXqCO1zvp8jsNEjQxwoY1WfzHl4MYe0i
MA1mhnuoTIgNUEG4kHmeroHemNK7848nxzlQN4cmEofa4fFu63H3xpbYEpuQDqCOIeJH4UyyV7R9
q7AuyIV0xmOWx0ykfkaIv8d/eDc8Pxj8u+XsQiFA4KMT1rEDT83NG//d2aLQTrF9VW/COap6G1pr
i7X98GnxIV5+plEIdk3XOYa5ulLkbofiJaeXJqLbdFJxRLzS9rTg53HQfMEMC6KaTOjoxk42WOOQ
91x908kewIeBLFZdrnnmOhq8LWiuxLrKN5JoGbcQYSKFcubfltazB8Wtc8+TrJcmQzUKzxOqx00J
yr6g4TiZmzd69PFbkYZwL8zlq63VmP5PUKiwrik7KAPl7helVlvINZQx3qC4rQYWa41M01to7aTc
Ot5KgdeDMxHWFe8kruWC6JUzcwpNNDDg6l6dWhUlqcjx6SEuRsQlXmKYHxqW+1rEa/VEBwZFlH4N
zQjEiNV86/rnuVzxYMgrO+ZAAHulV4QNx7JavQvk7n1ikOj5hOPl5ys+cwLdTZ5ZgpmVvCbUoghC
vWYCWk1J4tnm1N4W78+2Fe3qNjg7zEQ2KXV6ncZnQAEqbyzK/jQ18w10N1CUqZTgriJKaSpvzyY1
eqyQIy8E/zuv46id7VKpVHKqLMBcMpMErN9vwA2kM+/nz5WP5mD6xMpT18TRRPHKiZXxeVWTNUhu
oACOQvjUnXCRny96AcW9qWfY0CEtIcdwQZMJFJnjGUk2YakSSjAkFwVJzCXpP3HetvxDCtEcsuYN
PQzAPf3YndnmfQWexMJUJspe7AHAKoJkyhxdlICqt4sxE9fm7/ccf1Ts4HF9tS7/xPG/HlurdAjz
qzJPFU88kKPc2yL3SyEqd7UsOFW6SQ1qQ84JaYFCa2xGjxEDKZh0nuTUiwOkTq2mw4pyqWKCO0g1
7lyzcy9ISc/31aLtqY68yw/VH1Nwd04L2nsddK8K5J59ZS3E9Gcl6OFADBWTLauzOzKXLZjC5daL
ePyEn6X9pDIuSQh8O6AvzJ3e2oNA91C+xVG4pVYenqfGt1qRYSI//okIYwsDFbDK2iTvJXF3EA95
2NSTYH88JNIyqzzhxzVMOIqSDajUJ4dGuCPjdUJpVGD4Uu9jcHvv4mDcid0GHZS3gQnhybdTvwF8
xCXVV7m9+dPygjEYb6hcUj6X+0EIbZ+OQpb7wd+Ss/ZHr06rqOoG3ruFaxobySKDtP2LyPPYIArk
rTUd9hoScIH6yDT5KaAOvGvwiCLf8ldKR7hrB+Dot2RBaVwVaIgcizqy7XfxLrHlgS4PvPO+a72I
WXNKkIZIl41pU2sacdnh87cspjHgMFmmERskq8pG5YcSxB++K4ZAJOFs4g1h886B7iWNi79RlCX/
9FvUnsObwFjurKWnQSI5Zs+CK1Bw4xL9sK/LKB1oP6PI8lXNzg+HywfgpexfRwsZLpoT9V4i+pSY
0Ve2j/Tzn1COGMRyAmDOtVtteAXRc6vtNNxPvf8JYzp0UJtCVRRRLIfn2au/R/XTzH/gXe1XwEOZ
WbcCQ5M7Cy3giJEbBfX2mPVsr6Ac8MBHF9JwoNK2Y/TQay0Rqex9OaNQqGtqNrITzFKasfqY4Cyb
/uYSYL0XI3dSKvNUwU+aDEWWmTeVmIdQDsT2Yn85ByI62DsIcnCHyqlI19gVtP0AvzO58Zh9Ou1A
NjuEpah58mhnY5qH0xjb4+IJ1kp3gtWFxsXxxfRNFO8mx7XmlkUjAb2MG9UJiNworBQ2kYh7Mtdi
ca+XXIj8JOl2QXurDEOo+y5tADDc7Cz2Kd0nwm3zwcgzcQ0GfYK8RNjvc/eqXXwzN3aeGJIQwxI0
Ujtvp592V0YgEZdwAiwiN5ITtmqSqPqhh6S9qpRm1mByT3VKfPpapL5AziHto6sWpcZYRfL1oLiS
04oMVGp3X4k6RIj81an9XKiCgYa0lJyo7aWufbj0k/gD8AYrR9G901s4TPiTGd0wBaIWizls1vzA
nVwS2Gc49rrxNLppiAn9k/EDMh8nnQRr8s7irCtJUpm5lA1t6hfcutLzGMwqU95ufA6tLIuF3rlB
SRKdfG9fScARwg/k3EtNZtbemPsWaBktjdC3Cs31jEuKd6w3yRY48TZ3Yt3rMaxKsAMxxzpTZVWJ
K953KNbvwz+3knR0+ITwXji2UoiDrUWkOTeRd8W49IVI+NthytH67ebOl1pqN4ShtEZlBW87JkFd
C2OzdcJuMBU63HTJuIHYtgKJcT4z3wc9L8hJ1uDUzbbs23GFtE8HQDMnIB1HtopfUatOOxmqGyRK
98qe9m8AQ+l/yaX28Sey43UZaqwcbVwNSWkIvlze9SdT/eN/Rdn/8cMPnd8PCx+gFD+ZOiHh3Qc3
UupLDQEsN4bMlxceaPNnZ5YHSXsERb0M+sdcJz4QJMELUi3Nb4tQRnxOKeUSdF9oYaE8Uw6waS6Z
1I5BWfHIa5iFZEuXqjTw+8reG3gEf988f6wEKHZU9gcXNNcxcRTieyUxGAY+eQolaclWObBa3lLZ
TAsqNTkW7abbHjvzDLXHfKV+qXGibUahMIxJstTHNtWfDgOg5proN6ic8rBoKAMcg+LtzUi97U8T
JIThZ7rnr+LsIy4otchLksFFL7VOmvJW8o13W20zINdeKbCn5ufKt/AzEDb1kUcx5uiOmoFYGqAt
gpb+Vsxq/WGOvI64wxRqgQky0Vn6sHxlqhnSkrOiiyLI5fuXg8hI1Uz2gxD83Q1g7HQr0Bt+Jp8w
jUmYZAEAuS0Nz/wncDNddGpMVS6fazNpVbRCvlC1qstbkjownir9Ot1n6leeU4RKzHa/VRCk5vKF
nAN39d6wxO+TzhwCjeV/zqZekPFh5kz744TiHV5uU03YgLd9cMyfb7oi5R5en6FqZ/MspbouQAB8
RxF1IqJVTYzKb75ckFHuPbw4yB5rjeyfxPfZx4zWZP4oLnFK2h69FJ9m5WnvAHWU1JA09eoO8X/l
59F4qQjoL4zw7o8QgGO8xrDrqOOBPEgiGDgpt5FaCzHyvxwW/d6f5YxEsZ61Rh1Ax5OzVqHWKYT1
nL9Gqx0JW0v7SmmacFiTxsRcompBEF2SiQL3rXsivWBQSYT8QEoQZArDfYTQp9aXlr+VbZ9+jGiV
PMxHQiYZsFa0kuEGHu3uaANMgzuyQEEU0cXJzA9QNqg0j99CH+KrIr0pWP/b0AbQmppFaAu9pzcP
E5CC1OTJkFg8Z2An3/tURVMC94Kb2gzZS9tAwLx/ScSVdJopE5QCe40s7Yl1AXMbfSsniPYBvA5/
GHVzkkm/pdR9SmP1NqT9K4w9cpWz34sTAeyTVUX5Artf1LLb3PjW5vHzzAThm78o8XMU7fmKxVIA
ZDHxydWc++wUUHvGme9cVrwYgueERcd7pjvuINyUPhjaYMmIa1SKbl0vgsHBZ8tZMU0GmOJPqMSj
YaJEwgbbVkjt3vSGVAJMQyqsSKK8T1Imz9+tAtQEcjYG30GIu+jY1djfY/ElebvlE3YpSxb6s92K
rNkbncLKy4xL3+/ZJz1we4QWh8n2e0aDK5e5gFlU2NIRlTbn4BHD/fHUEtOlmrnr5yrUu3FQb2K4
PDnTDOcUqtR+1M6HeZ7qcBVcIXSFGkRwsKKc7neZ9I3NC8o+NJjSyt/hm6Z5YaPpWOYhRqT9Nt6C
vzes6MQfTg5FeE56gveUmpVLqlRZeIjannn1m5sLWRz/A+OlmhEoeR68lfCplQY2oc9t2EoXgZ33
vcDNTMwmp/G0FoQucaZTaGEW4rB69UdJI9Q50d3KBrJh8C94oobABPy9Mnk/QUXBPvq57sDrc4Co
+FeAM8LDvANRfYrkGlTvSa3ku7t7H6RxKwlfcbkS7rZKfBjFgvX36qZNQ2agaG/NNt00/WHCWVe8
eets4ljyd8H+Qpm5b1bPyiaRmJm0LEe6H/uB5dL7P1AeEBi0WRnC1Z6emWTRs23JIjQl9Djc2lz0
k/MrQ8ZfEvoJIaRzYxmtJoV/2PD97kf1fod4RfiWwP2EmkPIxjItym7aC6XF+sKzYJpcs77rdP1S
JJDByVSv6r/ErjiuM+XLi6g44rlQI1mY3q2znDoQKZsIOUWT+nd0dWk6qGlAs3sJqFAbUd4EyCsw
IOJ5Ymz0mGK7GJfjzuASS/iFIfidkV0w5bKJc9eewsSGUZ2E9+wLsLuJ6aICPl57KQ6JAeACTeG+
rHB5HYZIwZMWdXq1GWUTpvkqRMbnAL5L/R86YUYnPGXdnWBgHkwjDMGRNU+uExHEt6Zlv8yYT2qt
VgfZ4NTbbXRu3ZDgSihPDpsycK3QCs0dXF8qlk6xGkGW/TrO0IweEtG8R2pOa/VenhoYhf225gaO
NxXoWHcafFNRUg4O8OchX0SkGufdQtWt8m4bXTzMCRnt+gdGnY/nlIRzLyUAlnWUkUVGvNb/UwGS
fCQ6bvuE9dxpjVbYHSUQ1JijxvUggH8nd+tkFeXZo/BJZNDPA59uirlJp5IXQcOS9cdw1cr8vGu/
CPHJwTPWs7EpsLQMRm+MxYtq34echiadwDcDMvDBjypYbRCzOOVeV7a7pcE5JRz1dOiKyqZJ91Lr
69oU9jccs66A4T6o+dKMjEzcIqaQTuiF57FqUOY2OfNyo4gFApDsuXLgXWQFkEL5ki3JsAyqhZj1
Lm+WevGcaDw4dt5S/tIfxzdfZNQfKEsbpQtxokYk+elfJN+GnsrLYNTPYWMPUQwZwQ9GPQM32SIh
CLLU32Vr50jt9WrSVLF0uXKRPyaqpTWPg9iqjK3NyceTWTXXBO5+y79VPr8o1m0+hK8iNq3Y4r23
2JaLT0iD/08pIcD00RmwsVGr01wgiDxHUKDjiSkVo8qZYvyANjx5JcQLIKcJD+xMtWvdxi1ykwua
Zzn2+k4TUFIRAjSxheNkhPS29f0g7j0q1IJpR9RC6i63ue3ZtIMlgW44qJabPgguB+YFY4Yg0bJT
S9bjLj/ksgqnsSjvmQvQ+1/nOBmd9R9ZF3AhEw9zJz3JQsp3sGnHlVylLQck+A+QenkBINubbLZ1
ehUzD3drvWQcRq2omH0tXpBLswtosBl46zDkavDAyjpphKXFim9zC9pVyQnFx1yEe94GVauCxyw8
Pj0vc3iUfrTqTG6tnVdKgBCCkoinCeZHXh0thwpXJLEGdJksHXyuNH4pSn77UOk2ZtCnkTjnDcnl
eJ98cNInCxIBtI/Gxzlg6wjsk89ZBOTBnjGa1L6jZG6R4R0dYPoKmSq21VagocusmPkEZc93jX1l
CQybQLd4eecsNVHDt7L7YD3VWTVHeMTmW0vEaTKDIFIunaMKy9DI58Ri2lLqt2S7JOj9q6WfoTgp
ek28Me0Dy4qqalkz60sM9HPwr/TxDU093NDhXvXAN/OwEg1Varcl7lfnO2RoDxD4FRjHwEhN0LeE
ER7NLhgMs5A1fKJq8CEpolVRrFd5cONswdF0lHqLWSS54e2iT3vy45U0ZOgcpV/TE4XaTBiqxxAH
9IEBjWr7xwV4CEnQ3kXWOm793jid/nYMjNORdbNPbc6iV9PVYDp113SIuHNnFNsPpjOfZ69DxfZS
Djfil4e+2au32y9HNqXaWOBL0028K8ZGqNcS0ZGdkPt6YxNGv7tU+hYomMlHP5Jn1ETHf2UvJgB/
MqwFGYv5vHqRCbgsyWm0NBSHeonw+zt8bnAhtXkLssVTAch2PzPCa7Zgzg7B1GJT51MZNdg3A8Ai
TbwgDM9mom876FRXNDUCk2q3PatxU0AuVkVLtR6XZP/my/eT4kEcJyB5O3c0MBQ9a2XRLuiDGqDX
OODTuoGA2QOJuns94vNo6gEkbzge9bSWrxp0ITEFY0T2Z4/S+pWyrnI6StMaron+SO5zTPkpeVTR
ff9P/zHCyk/krSZCnMwz6uDIG7miVayYQ4JbIoO+YNGl0X4nRBs4bw4G8XhuARXyJBFoeGG96CoM
YWoMSMVA16sId/EqMEglVvgee1+ttk630JqUu4RoSOkY36xedlyLAUnioQWaBxkFTOVg8d97w1rj
bj+iRlinKangXYqYqf8nLnx9UMT7/nHrOndLwqNj/wnAJcBrK5KTy8nrilsr/rub6umQHmFq/BnW
DyN+koH8JqOXGlCAMA1Cd7oTrwLQ1dbbqouWerynDDAk8BCzHmq7+sExtvGsNVuf1gxjFsYorNS1
M4sE6iE4Eoy/i+7sxZeJDfWPxOWTsfdnINdv0lgpJwAlAWUF4egPpGyTVydkw4jdhJ5dG73mEYbF
Dv6nAPPerQAUYa24MPfiz6RBBwHssLLCnqs2ZSDXHZ/1OQ28hPKmmRjZNESCf5lgx0TWKn6bEw2m
kmG2MkD7HTe0agWItMoD08QHjpe8ycQjPOY7jds/Ase/2DeKkKMj3EmAAY7Zw747EGLUCOdfj5cM
dagtf+/zEgUIeUnDJC+tr7mD9ELx5ataZajvo4s6rq1H6O3j7X64VTphEcipVU0mfkVtqOCvZkiN
PXngOg/aNzUSdKKpIoIH7E15wZFbFMvl7so2IENoq7lgw1PKujrdC/umFFzi3jTsgR00rih2zt+J
qF2RYjplRIF4JqtiW9KGI7zgGe9UDgTDPyxdX35ekP+qR5vEi33J7WG5S5AWlI0CEO73kB3KSphX
H8b68hMTBaYNRxqC3fvKr0gpYgRIsAhbmqzQ8sPzVkM0ouEkYs4AuO2e5XsBU0ufUHAMsOnen8TO
j3f6z16BDxqO8J3xXZ3f/9Rz95GEu23KJVMdEmedb21pYXQhMUiSJtJq64dGR0uiDmSr43o2QxKv
fPsXrz9jXGhOd+ZV1IrMha/3BuNA7dfrNf5bRUTi4gkJcEqyvp7pl4pNKaBAzBQO9gCogJycSGOr
dvAomMVevO24wc+FoWhNpi9Ez6935XaStcmEYPZnEXMHCKVS0000HbFxavXb/V/IMi2i0r0IKg7g
amfoG6gC+DS8WLvH7nlGkU1a88S5TapSbmFmC3PCM5GXnCLyu7QmGlNjfAo+6MzlvjmYWVVIj923
38oCE8g2Y+I39aHUSGhJZaW86WE//u03YI86J7i6k6NZiSQgu+VDXixVybIZOtjl/kQF9G/hM4Lt
8G1dde9OEedKxKolLmWz0n0dlpIEXYn6MqQHuiY9L64kQZfrzqm7sNp/qZ79vlXVGoTH9RiTV+A7
L5qsSiGQG7K+PRSFqnuRXwW/4+UpOPZbyiPbc8wexVktMor0ZWxMuvoochQZK5jFD/Ds3Z/ggexC
Z7+csG7y3z9KPdd6NQDW6kOCMOjo5UnrraHGmCi+yHs6stpQEca7OV5lkPSfKeMFWoCnawQMijEi
QHRP2O+xvs2nIIj7sRQ1V9SjbMXahyAtiFtzxox8188yvQfozBaq+pf2a7p56WoZO1916/ZMoXLM
wWPT/+U+RxbZgc6uPKgUC6T7cNvM6gLPEOcls1Lg4RitXp4QDHZumCZEeliHy8GDTHOMxMRCWZbd
k5KEpQviO1W9fNjO187vKICMwp2iOffYypXGxuCrYvA4HLPoTq5V2GGignZNAPUyle/KiLUZDEK7
sIo0mPJoemgLhDAaZePbPtyGQR8lrzyZRgkZ44xReMXCkcVgc4a8pM0HwgusTv9NqUMe/veKdQZK
SJ+pS2ITwbZa8gyyr9d7Q++6tgDywIrd/9HhvsdhFD/vgyin7G3GIsLiIWjp/Zr67vm3SBMcwZVz
7evin/hES2GfADkSQ4hD/LNmgdzVI2h8gZT3OmVUBqNOwxt/YCHwlLlNoaOxrnr2+TtGgDm8c9yi
+xerV7gF3t+jdKviRjVDKwOBAy8NenvyXW0MPkILE+416Z/dGv7+8T0kkLqXCW3H/Ef+ACWDTuTW
4TWwMcBYUo6GcvpEFD/XsWtmlQ6KZsLxlVy3Jh8HHJiTTCJIKj2/K1Bn3v+xYVenqRqDoJIXOeCB
sCP/MXBdXHH648Ou2H+bGAMPCRoSgOxtDCmJ+bjCOmYarU1mARxYgl9a72T+jI6AbAVe0exL0GQh
y5O1433URsRZtwxu8zFa6Ab81ptVwoPsR+uC8TV8uX9GbW2t9rqcX82BjBJu8jya92PqaCv3lZ+H
zgXdWPOSFkPnUnGkqjz7+ixZrknsGUeARsgc+VvM0B3K4rzUaG42HxnATbss5GqgksWXRcMyM8r/
4YSXo1YahbC/E4ufc/7C6NU1Tbg68aaYE2gS4wIbXEOhB9p9VvP0Q90arNy4QHzBLFVlIedL8t6/
hsC0uksfvAInRr24cx7nnVcrcJc+WGIWq75392CkDl12FiWM1V0GcuzXtjq0rXsCKzUWnpLmjyqM
3zw/VZP3l2Sn+9zeuXZF5a+1bjSgH8huewfCCzA5GBcE4gsC5guDeoPDhgSJNwqX+IhTi2mMfAna
afXlwP9irt629ZzmRgXi/eybcsOZe0g9yKmJLwqIlCNyc2CrQsDecX2tOlVxmT/I4WkmEA3a6whR
kKjefkOKcNKrlpqJU8JF/orpcjJWB4RJzKzcMdb+HRVmij0u7fpEi6nSUB/jMohGLU//xcUvPc5N
GOfSgnNO0pDrScikpDve4rh2hYl0qO3HTo06Z9/L3tHZ2+c3B4NbaBK+dNrGAyXVD+dgGC6/n5KT
ymobvx7d3i0u/Q1Ha6PK2VLQmrxYfuqVrcVILdTGwSlfV+o+z2KgvyuguKkbRVNIPnSE8Bs5hshD
HdeN/2Pm376U/BUHGAEDQuAeNqhoP8ODerE9JSrI2NUpp+of7EUMtVocyRjKdswb3b/trwxv3hSM
yb+sTlKTlnqYXvKkWHUe3EUjKzcHMC6GCmwYfErhVuwnm8oWXToW4sE+lCX/n9bI6mQAAo1S+MaB
A+dLxIftYtkYZQXT4ofNxG4VmSekQmGFtqZ8n31GuhDeD7twoPApp4Sie7Z6MFehZe3XaoT9URny
/4Neo+HLwpIZxzzPMYVQfA9Fu/EmvoWUSkGMesysKf7yMPE3cRCdnOLfUgqgTWZb0qnAnZ7+z3oc
Mrbvxo4TgmMzsx3F/eCiFUjwb+/dCCn31Wop2knreow0xmni5+cN24HM1gG5IhIKwlwh7+Si9jx0
V4bnSJfKwICh5kBiKoHRd9kUgooz7BKB+NbTrIh0OFmF4tL4pr4faF+Ui4IjOaCMQBnx9G3Kebb7
5CyR5/S7EZRYumrdYsdlXvgJm2b39EZNNIS+aPsr72DVDle4xGwdymMegISW1pUbXzKAUbg6v1GT
fdtyIL+uMjZDoIL85Pka1s9q61kWo0ibtfLjvACEUdsOtQJxZtyrH6SvLhrR1wLaHewBdTWugMT0
OskCRGGwvG7VZZFJeNtJQxl792REPieejBlCZddMR7WPvisQRxgkDpRxgn4OdluDPYoEqB6x6YWw
91MrRkCuVnSNdLTZcKbO3ZB6/i0PLiHNWeVP9PqCdZIykzO6BXbb8Y5WUxCPqsL7P4eFGRYdTO/g
6+tuFYCzqY7uOx+NuSovhH8OOAQ2wlR+DlS1pd1SeE22AoNDwr+GQsIxnKirlRyfhI8v2M4ChMmD
IWCdh7EOX3CCVXoeXa+HsAhyHypfxVDLlc11uPXiFc0UMMJiO+XiuNFXIJvlWRL/gfz9DJ4nBbHZ
eiQ+0oQ8O7SBSVezknkN/2iljBb7ujHyQP28f3bjFZHhXIoRJ18ScWr2ne126Xp9I6qgDFOMxHqr
mtuPH3yOk2JuQLdhFpM0/4WNO2eRf5O1hJGCVQTK6/fQp4HS1pmmozsefMopklSjjigddDwj4yPc
Fcmgh4cTBexnX++V4JFKhsZgDeobtN8ErcKclo0/FBtNzNJajskktTQbIhiCaZBR7DgUX8v8p5FM
bvGe2o3SH/fYfrSsmYvwubCo9bIi0ackzA/oxiiTM5/t2ActhCW4mhUNGsCBQvBfCeKLK+bnlRUF
ujz7yjvw/YTh9JAs58jb37yz0xhL/MEZfOE/x7TJdTUgIi5Y4IaZkOavyZTuNARnuy3RxQmlq7lN
6c7hK0iKWB29l6JMt+w1tburOV/oA5NL83QZUbA4HJRsL21bH8qFh/T664WXTqymQwmieGIqPqA3
IrCOirB0fyKNYOI+7+cMx9Vq0BQvW5MnZglSx7RO/+YoLBc1rI8AhnZ3mpf/TjQ51LiN4BDnQNXs
JSz+FoDVfCrbPk009afDrm3vuLONG7vnEu8L0/82XfV5bfksg+2KdspCpnfi/HcBezoV2s6/2dNU
JqXbDMAzn8LWT/siP4YsEAF+k3OTF0kW2oIGA+LRCYL0EopMnSvJKA3oH6yYFeAlztYbiDtpsi6Z
EebFsfZqV52wZVHQ8MXVBqQDZKk3yYoUUvScAv1TjaGGI7zVUDAotTPXOn5mtVdygpwwNuqnWsRO
E2U50ubmqpMiVca6JuoE9ooUDMLnqxpwTmBK7014Y3QoK3Ozg4rBCmZaN5MPb6JykU6et425qsqa
BrNlW6yrTPFAQAF3LPVco0mAMwoqAHFB9xnRSfRjam4pk0da6G3g6tYkRCSkNHmBdZ+a/m3Hnnth
bmOTmTUVGXW3dAKwY/1wS1kY6GlV9AQrHz/rl2uUnPbq5jE2jH7XC2phtD/rh7xC5lbCBkSOo6dS
3OmBVgR7Vp2ylhDXRwdTyX5FR+DZdYTzZYTVJieVc4t2EDq7bSN4KVGmN7vlHnzVDObfE4pYd99R
7fZfPmL72G4G1XgNTjSuuV5FD2D7qBlfODQtUkynJS1Y/mellhJ8bO+olzna7Nj1h/wOA/DV5MEI
pJRF1JhlkuGEld9TDhtg1bc6UaUdTVck27UWCE0OgRJ5twc1YJ3Ih9YA7mVulzHGvz+ipjlk2WRO
DKzA+cOeom2hI3S1gZmJQ81H0iR7vNyOTcQdzdvKLtMIcemPIQc/wf4RU2Owxarta0WEYXap/SVd
AqW5EW4YQNn+DjE8gNs/kyt4AewV2Ew9lVuxivngPCZRHfhLriwgvYdH2lTHSD9rEUOj2ynr8bJd
k4zHZmDRAJb9iqKcfOlh31Xoh7e3nCjzzeVsBpy3o/nT3KlOc3L6kEWfbOWF1NJcJ5WtJnL/bGR+
1O6AuPF5Okdsc6cvMT7wog3vVBgBpdDbzHhZ3Qh1nhXokWevY6r2HZT65hX5CJep3e5K3zzcX7/R
mHdEEtgEZvSDnLkarOHgqI2BUYO/Ele7fLC+Pi+ulBmxPW92Xne4RiDOZ6xt1sgX0st/zf3l+sq2
Rs2U+ARnupyKREhk3hCd4j+bQ0aZhXc4saX0/cm8SWM3frzxddtdVi+GL//zA+2LtuvWVGcfX5a7
V7nCydkg1p92vXvLzvO1pJ/2dFyQfGAvgrgbY4fFV1PMP+tr/Gucg+Yd47QwbX2NTy8VebRJnrlo
ohFJ+aYFYH501oSBCgtmm2rZBYcr1ILD5UIFyfveO1+V5Zdr0aU37OQv7LAYAPalJuv3QSFrT1tD
6Fpcsga2J/rklmvkKiP1FKTkYr0zV/bv3nOrQ/34h2pMDGiKMNHzQbwEk6uJZU1x7s1/fBzgdZ7l
JzFK1CrIDdCw8tHmGshYxx0BJIxy85pLrdXeMQ9H3eZW3xGekQJQloXJR7sg+4QuItYbMWYkVWAz
euEWsVKPF2agdkho0BNJRTM8C6hWRY5u04R9mCPm+F/5ZMLkaBeX7W53KH3pEtVFGN30D1qNOqtU
WVu5OIgCBlPTD7PMLNuwez4VzSqozfii6R8Fq0+higB/yrul/igsDLe/BPzsQHmTZbd4cKjfjl1Z
WZ16GGinURVpmRAY9XTFNF5XF/sYSPPs10J7ltF/UQiM0Y7lQRxj7g7RUv+Kdl5JBW5jhWib8CXY
u3Gy/Z8uy+SFvtgLwY0gnCnPetFWViXyoNQ2WnsIp2oZH69gRu0W3p1HE2Lac7eU5DxQ+7Da8KUR
JttSVZ7UyDkh0nbDTeo9h+XO0pVZPvnV3hv2X+BPN/DfVt7UkFE3LM9j9hz5UfYRhshihNqi/KoO
QJEiFCiUwjcFvyvlwLUElYzNJnZ7tDra6CoLGj9Ht9G01CaGe8ANKjP0OY+y1iDpiUlzyLElKoTH
NiJbtIZ+g/NQvMexJDjVjuS099SMXey4JWIlml1RHZ06yOWdN4aAq08iG2rOmZb5XGy4dINc2V+C
Zf3bMO6+ESWSw7n2VlU+sm/T8lmRqYkQ5xRwesfoYnMvxWLH/I5VZNdiJ1LswCwr8wL9DaWmbCJn
MgvAhIZ91NTb9vK2fwUicZe35+waRUYSnpvqJTl2e+2qe2Gki3lMH73oiElGLOWuxRCSdP3++SnU
QomVMXaBT/SET3Wbs8MhafmwSneC/dhAhFCCqHhGVK9uT4A+LeCxA0zPXkgT9JDkIx4Cm2+yMvJL
7WGZwDLzT72/eWuGbjsrjkFO++HHLStVywP/tL8D+HNgbPwk9rCS3dcljdgy6pFLaPx6A0nljbVt
OQPcnRntO3AS1OAm6Qdt3UB3cdZL1ILyl/TkabuipI+iRm1SxZWBLoPDBuvp7ci9PUgBg+qCISAu
i5DS7dSqNdNYO9CmjJkfYd25HOIWYY94qvRZHw60Lz6XJOx0h0Q0rpIp9p8QogcaNdJXz3c4K16F
o51SDWuyYcdOtRxyhMhDCIEFIrOqbdSusxqRZ4CPr+2fbnZvI/+0+EbK9L41s3RHcU7uysrYvuRT
EAYOfWJRAeBrMlehFlcuGKLjgFN/qzJikbLgRB2tfGCEizeyKraXgEvX/m+IMGlc9SCyO60IJW0h
H/VcBSQZWnpm6Y8HtuY07PZKtQN1iWQNkXbNkp+a2ESkt2eNyDQrJkW9n9Zj/RQZc72xrMbmLl8e
s+BYcoFVMoirGpt0KujbREDQdiTDfJBb15kRhW0Z+4rTGnFeLEbMNONg0YUKpQ+TFQzw8PwwwYxP
fOG31q5gAED9uT9rz5eP2jl0EoC2xk/mT9Fgzyp+HtKPxEV/CdOtlZoQqLAM4cWnPyj501uTirTl
zA3bJ7U3/KkDj7nVur5eTFmjv0LSBUHHEkY8ZXjnVmYHJg3MAd98hHfcKCH3QYO1BmJEtSqgIHLn
t8ZLeu1IquwSNfwLGROuOV9pgt8XuTz/4X5tauUsvasGVLCo3lqXZPTbFjTiJvOFSq0HtDVodMf5
q/xDkrP+v5fkDbCyaJ5USfXLd8jMLDix334iOOhSpQiw4SpUeMQ+5YkHEzEGUvWwcHNRbwlCL58w
W7VWTfsi/DbMHXqfYmIhYF9VMJFxf0F0n2UaH2aShb/4ys723+HwIDuSHYgauoYGW67iF5wBIY+R
xazFlsnOmQnmE20UoYln+MRaU74vxA70q/Mpz0wkcCmXCv1XhbkC7gWX5dtUfnBuzBR72rEM9u22
WQLZASbTPY2oQTM2+9vxuCevu6LK4mAq3tYXCfbJFtJcHheT50Y9IMYqMoxDbC/Ebe1yKbkK0cS+
DOMByXs+MEbbUb4ulJAiHaSqWuE6Kdo1UsLPMBfYFeLbeuTqlugBRgYl1IAa1xg5oEY2kFnrVJCB
gKuwbLvCNcSOdhcTs66H78jleqc5n2iZD3fnzqG63wpjmCOQ9fLk5PkLRLraiyUJv/JS3CPC4of1
DrgHZ6o/6m5CuroEUupKwMsnsIInG3Jlu2MWvYnSZZc0sZweGHepVhbtvlNo90Gx0OknGeUaRc2F
z6BvfBDMX8mqW5Hk6MZ70DE/6jl7FoLq8BfCaQnKjJBA5HNROJO5u5XAJ2sFA2znksClGrcdA7RZ
keYzkysrRgCIm6UOZvtOjqX8lF7Jgfo/53tDzf4gVWnT2M5eVrCbGCGXrgRBc9w5nwsPEf9LhqNU
AylLrrm0/ermL5e/se5Zzbpjh5i87f0IQa+0cC7nJcrplJTAuLhrnOzBzsaLO/ckrbkDcV0cWZ1r
k1VOyWn+1YMeRh6vxzuWftZmEzD6HHYK6PMT1uPC3A0X/2RQKmwWAQPfoKk472wXUxS35ou2u51+
CsoDKNv9gpTp62ATCp1SqAO31BX4FIf42vk2NMWj3G4ZCIR5EE/3Fs3HLdTrTDZjUOWON9bn5FpF
/0o5JA2z1dy7ntWcFckjYVmRd3DtSHnVPS6+5YuxP3sAaaSTawffzhaz7y9szWmnB0DjXqdyExCa
o8piFRQ6JGizEsuYb0UQ3cRZ1HYRWrFCvyu4i8SyDnptwoTzPW46O9yWmFGXLbrO2OPaTYeEM7Pv
E61LSdUNwx74pO21NY2z0i1glmllxGjSBjLzEQQAB7uakLzchJibz5yJQ2qJSBA0ANdbIi07RS70
026UU91Lom7xq/LBegODN92CoMnUJu+UjWhmFoa8YSeNSyv91PeB4z9I9c8fBnRHIhAr2Rq22d8e
l1F94Ff6+vVdlgVsI+xIjpbZr9KPGoXx8eiZUtEKlkRMIBls++Oz8RWVhsnr0HOrwbwL4N/rIxRx
oXQml52/0vF/9WY0Cs+XMNPJp4VgZM3KokM6LcrpNZjF0B8PWGWc4BTA+XFe35FF+b4oLVZBX+Ou
RCcuKF3onICFQAZcAcsAbi/Z0q/zAWsGGuaGxjlfwdyigcbo6c3ZNEuQjWPhRnBreMbn/8sZaHZl
BZO4xgpS3kEBFS3dhkbQfnGIIO61KExNZeS/mflHJaszA0DFemErcXfavmWGBsXJYd00yjti3w/m
kNNAg1h6Whp7n17ucHSPyB3T+rgS0IjudPa9x+r1KXzF0NGxWuqgliQofjYrIgjw2TqFRDnaFZtw
7WeHF3mJNA6QMmyfIQNECHwfJYp1MfrKm72s+MeWURjX+avfvF/UMTBV+rrxQB8EhPOFJUpavsZA
SXJL8SD66I0PYV2gygh2W9/LWwfNHhfbCVVElBa8ykgkZYHbaiVI72S5szX3IyUgCyXZ0VUio8wU
enriix2dMzMASiluQFWew2Z3bxaPgDtM8xJN+EkY+911XbFG8q+FOY4GDQNIMdnETaDf9FFenTPq
zlcVRcZiZFFQmgpMzZ6u6nIY7C6KfL7W6vv155LzaqeZj6Z+t/T+EPdyto2AU8A8vZderu833s6k
TFqts4N000tbUd1IwDy1Fey8tKVSvyjsj60uaTTghhC39p2kRMOA6XtPVxnd9p31IpBAN+2/pgCP
4ZoAs3uKcyPK6hymvVCJ1x3IliT+rJZkQf2WNsS3xnTrg9s0WrY5S2GyP/m9rrUkoiuO5e8YgUUD
C6wsv4NadY7TrrExIhqIGUNYXIqKcOLaIAD9YkvIgcG3rDHL2X4pL5FtlTl4zn2tRhrSkIg5l7Ay
S2zTN9oACEabs2KokaUTXzkMKdb+0cuXjcyadplWdEYxi7YlG7rvhpigFvmn7R0g9WV2pY9zQBYL
Ooad8+RVZxWM+HwYqVc7GwKS57qDZLcJI/OUgaALYxlDp8vXENT03mg84qMtt48UtzqNadsYykO2
+IM3Rl2qEaNk4IqtdfNy1Gfw3yvZA/xUj08Cg6JFUygmulGNSV80MvJHuQ81M0B0VEurUP7HPchO
y6GtyvbieDyQCffQ6wEWLalTP050onWpqzSetMIh6ptvlYI03nPk1+5qxYxN8zsPl4mOq+qJ5KWZ
AApoNOvwP54+F01cTJqys2T49e/rHPMs/Mlf/qgtOWeGljONz0OWpSXtKcdd3w5GUigPIIx/ibQY
+nHu7ZRha3dnngZlSZhDKAEYzFV2C5xFTVNr1dVpcMnTLUNkhQTn8i91B2E2LA/1N05oEUVnoOwf
uEQXASnw2D1VGnrxk+WfSy9iDN8HaZ9H504H9Sv/W1Pm9QHGHqD5YO7OE39UvjM/bn/2/gXEp5HY
BUKPv/cwnbvlEnNQkSxBkEgLTOl7/OrmW96jeIFr1qpppVgDf0pZJwt0U4KF4HDkB0vqJKB+kEz0
wFxXQivrnREukUtMOMO2oIo8Ue+OjmWfiTWS3Joq2v5MarSRMYOfGl1vW5f3VCz5VWewQhLK6A7K
+h3lCb+aLoEVCbF0b0hK6iVPVpEfbe1fK6Mf4WHXhfu/pxP1D1k+FyOQxKwTFQceh1tQBjafg6U5
MzJ6zuZCSQ+pETNl+LdUd3UsBjyBV/1IOsdMyQtsKfNV5JyfFh+6uySSQ/Bbl2Ft6yh/YpLXmpxd
PRcsI+7eG5kVlZim6MxHH9tTLYnWxvQolvzGmVnjwJcdjU6RHUNQAcW5rgaAwtPnc6vdjeURYyRB
Vfv5v/n1EhC/m+cSNk1DO9vrktAdTFkCdnHh1Ldtku/O3pFisEGJT/6VGvjb6UO9aXwbdyQEa4KE
vl6FKcZeTeZI7Ilpw0yihHMWnT9Abm6duj9UldQ50myRpXFYU53+WigbRRoSolhHVRnT1L7tOjs2
vfi9n9oBGmvlXftqK7fRAolgf9tOM43Qmrvuf1rfCUjmPhm4kBO81grnn1fUqaxL1tBqGsarFGnQ
t4zOBjI1e8Czf2gaBJ5L6K4D+5x2TeTF+kZTDNrMnvPOyvpD7O27+b/4ii4v7vD0t74oCof69FK0
3JpYTzl3nMsKMyWDIpdxWOuA33ZYAWPyahVwEEsguUCpwpxrpRho1Ru9C8xWk4olF0j0cQMxZQcp
WSlFwQNwGw5Gj2icws/BS5yvyVBOoa5mx2GXrYnHLdTVtCtwegLyscNIFa+tCwPqhxM6EYP6ytc5
9LygT0VsevHc4EDAMXdVUDoHBljXXd3J7OntzRNFKDkkEn8p9dtq4/yQXKIvHlujhMRVlhONPa6r
Y53sCnxOE5Okj2+OppB066A6YTKHb12+75ZZw0JVnQzh4bSSoXaw3fLOaImkuMYulIJthOQlsjvE
gYD/t5TEawnWSSqzcjUPmGoueiF5ovLWMMfMa3Ue2neIigqxZWxkWYkjjWHbzdiWrVVYymfSnPbR
n99qi+3OnRmP4Dl1O/ttxHg1YfFxQfCsU0rpy7FdZA4KWhc59M/gjdcqYUSQAHmltS6BvR0K4MAr
jgRK7N7+ZfhjsRXy+RC0llRQX+1pXGbRLQyl3nQnTU9X5eCVolu5vqpWp4XaqhWUoGvqgDW06o+2
RM6Q92BwGF3tUgCeha/HW1y0ukNVDBaTGNOTIfmIUwMX3ViSurInuN5XSPTG22qxtgDusYsxRv00
4U5ZHZoRTpA0YR16Vs6fLq0BoJAEfD8k3z8bmYYL3xnLERXETxT68KYDsRahodjr9oxDSz5lJ7XA
GvrNqTwgCr5SxNK1DJX+rkuQSOaQGVKoNPNMp8MBuyz/lbrfSEVBTLekAschxPWdY+18Y/efDlDf
wJ12OwbRa+DZ+51RAS7A3meZLXTNesZX+XsJVmFUbIlhcL4fqyGquOmry+FmNCbfCu6F0ewlX42q
8Dw8RYFYqVBcLsU4V5u/qe++c7ftKV50opznifStgLzdFhcC9kjtT55m8Od5LmB8Cu8ZrxVBzEiF
pOBr3WkRNGWlhyokdqUvd6zTZyhFTlusUNJsQFoB7R8GebobEvvhGlfMhe4Py27FE9c4bjE8DoYx
QcMvgs3QNlSo/1O0BUjW1+W+N0P9k7O7OcGMlsmrE7DUfdacF+HLJV9VBANDkeFPtvV995Y+SMut
Zc+7Iem9bx6K1cvJJIr8RXRFS90rrjLUA094X2jBrx8JbTnrmteDVaTLB20fZ1nUqijySzkj6i2w
DLDIIApUHYiOGha5lsKBF5JqogRiu9cBPOp6BRQ47Yk5FbyiKh1nJtDDJrlRW/uKqEFrlq6kUyXT
DHpicFlImlDnYQVoJ4xciFWYgArwoYNoE4/ISfBJtuq0fk+2g3D7nioIirR/o6lz3TWWs73JqXFH
040sAhnANOdDxtoU7+oHnqJ7LyzDlDPSi6JAWjcWpQHqBz3Ww8UjXWQSmQrkN8QsTEZiT9MXVv1n
JixjyUpenxmfih77tkotrejwlvYVODceHRjWL90Om08Leasp0P6MG0ywiyBItx0No93N3Fcx9yq0
A99i7XJWxZilIFYf43EtQ1Y+fZrZd1ZNtHML1HQ47BiUuOQcOUNNr7HFFS94G/EIGFIPpBBEc2W2
wz2kmdRbvK3C/gbHJPrG+os09AfFQd4mgbTYq8QcUV4vQoiiVPDeV4ocfOX01EkRN7eCMENFKtiJ
JmP5NMLO18LQnbylS76YcHId//nCw44hbtRHRIslevYRoxF9wGttIre/PIaG7UcYjSa9NF9yDos9
gGaKNHSUueslqvMZsmAxobMzCd2ebMJNCHY7OxyWpUulkbAZH5Q/5DaxnTJ/oFxZPF7Sbs1AJgR0
dFHUa9mSePsNi+v+ONDzVQO/YeY9nfCNXbZDvMIcXv7OtXvIUh6u5YY6KnqoFeBfu3TzQaVLltdd
od6KtmJz+4mWPQjoAAeJURv6i8xXXCPYDlZZXNUIlLg+LFKKa0VJm83UE91loXYmt+hwZlfi/oND
aI+sfqqht+/AC7AmKkyoIxtw7P216V+4VjsA8CGEZD0Hh0StiwpPhXB30Phjqznm6PMTCVd8DTuo
jLvB1HaaG8B9krqZUycRPGGf9zHDqA8upcLKmZzmW7jGL5QUBGZcF5nRb+vMMkUWNerUwYrjxu6a
22YsLrJP40W9MLR82hFhKV/LezZWQEX1or0rBW96B3W2DUrj02jackbwakvH9LMTA4i6KeqxUoD6
e5hGo03+vmk755xazRGvhCxbKYwI43/ytieVSv4sWgvCXBXgkOjqmrVo5atYWImMRCxeEAC74haj
aVyLAv+7SU23dQa4EbzetT2WdLKVvyQ+PjW6QbnzJytdYKbjovLP/CO6Qa4a8lUYUUD5dNiAfRpa
wRXNA6U0NG5GH4BiRHAvtR0ohYuRm7pveT7bUOxNKyoz88V4iawOlJ+1JiYqmdCi7u6L/hBNBqy9
4JvjgcZLdD0U1di4abwGham6SdQbgeMOC045UqV0u4rjbivLS+CulloY54/RkleIH+KNMjyzbi7C
KGnTaM/9ZHqbX95lC4R4lGf6ZtDojonB7y+MKEVBNirgkiafWlaHmpyiZOnH3/t6FwrF/l22mzNw
rf6kb5317KyzlHcOxTZqZclAFQn+d6ruUot6VI0pgPZCiDSE0OgG9gogcsViqlHSa22LLTwkuEZg
n8U0wU3Ii9MNQIOuK3B3FRpAhxvnQD/mgmE219DNXNGMhh40X+GCf+TBHnrfz2CqPS+acml7FsxP
J4jiLSxp9j2vgfhKqlVk5rRs4J0upxl5TzBtQ/FKZvM459ePWYGl6tBXWJMC9/Fu6pNg2DkbbvG8
NH/LDEOIE1HIN3to6j+fQZFmAWXuEFKvBd2hh/yhGmk2bCwEKSfiUb3iwde6gdbGfPJke8DNTnEk
YggjdUAqFhVMToqR5xLspvandFRK3CoiP1W4rufI7dEf8dKU9OWT6dj3OnlcuY2HW+3RiC2aNrpL
Y6bMXKR/u8uGynL457LPSlhPs4iMWdV2m1UXgblWLArFqcKU/TmbjMQzN15JUml3LiO3aDzfXVDw
ur4BumBXtf3ORZFs9dIHN0slhq06cxqXVMAwTEc36+xiIW88uxf9so2YClvLorcZo6/iNmILzX+f
E06sCQaH9WOzN7m3nNHvi8jxsQ0BTJE94xTS7DLMyG4FVYf1QNA5FySftuYtUDRkB7Tq/kQ75/0o
sBXDGt//uSHTdy/uyVvOWLDrTeAsijxrjdTL9/1uw16A7KNyCC10hpn149O96+nop+zpmi+/hUZh
lfLoLT/7NIKuIHqrouTRSVBnLdOI8+XlISE+7/9GxqWR1BvwbjfMd21eqy7EzYvDqbMp+rD1G1BC
8EgMSif52jslXzfLPM6bSZEUtObec+/9R9i7FtOk/IDMMvsL9mjv8fh50viEZ/2AHXQHnBmSMBJ9
lQib/4QDvH1egmX7PgYH3F+mJ9ZzF5K/LPAivSDb0prp9hWfBqoFxp7dgMGQvdywBUqHpnwFsQ9M
BtiZ/TQgl+vAo4I+7fTC/mHm+O0eZHSDA8pNo8RzzEUJDpDLI/WSgXn+EGCG7dbj+VdZL9ziTi3I
/VvnhbZ9wM0Wl4cDdTiQIzwIKsHhJUDBG4DN2+JQZKsmC6bjDKv08ezOVcOb1Eono6ExxsV+h2Ln
ADVetq8MIqz/Amc4q4h/hYY/cbbvxT6dhp5FttsgudBRgXfVw81bjpuP8Hm8ayp/y4TL9PPkXmZT
ZLQ4aCrAqpXb/c/V/fBYo4H5QXXIE+XWkrmrLqQj+pSHUpquWNxyLusc8jdZzADkxhimgv+wMq+s
0dhnK2pEAv1q8+PPnLvJxMoA4/qXFcicjYd7v9g5izi4fqTudbNCxs/ZngiLYWz6Yrs0ybLU5ARx
wGihsKx46asdjftG5us5aj5C4d0LIzmMOPeRwRzyYHequlfQ7DMv3uRbbNg5N7eHxKvwlgjE4E2t
VLdmqNxa5KnginsNQIdR0GmVeJzQ3vGn9qvFChbG2tnpKBFPZGArfr6KfYDQyxiXxIhxAZ9yMCtw
QTRGE21eVOVeRJ00SbN/YvRU59asi/QpDuXgr0kW3QoOASHJWYU/x8om+vkkaGC17OP1Ir/aBa2Z
OMDkaatsMHiY7svA1w8WMNlOWiZIKgdrkABk67r+LyoJssFPYj9ANiVBWyMt6xxBecAtyHnCtHXI
cnCmLkI9urpXI7CO++01D9g/yQfpkGU8H0WXj1MOVIX7XuhXr+PgovzTJcXfmYD4jvFeSucAczKx
YXUYMre5oKu4bHruYWVvGHK9DoRkd+2A0LCLHqbjsSk0SawOJ0QbOeBLo9WEID/3S36Lb/ywq5yW
1QoEfhvdW36QtMCpJLEebi+/ePbxVLTC1HX5jPli8HxL6Lb1h8PKfxkuFvDSGmLwod6sJtmwIZrK
7xtqVlCOHnU1hzlZEZwoIrOKCqN7u8X3bi9CMXfVMzxEaWTSy/ItTc7PbjzUEi6qJd1RQcrfE4u1
Um8EoOu8Cv9wDR/ZkhoNKw0JH3MiRpbn6NSEgcsFgPlJtwtn9z04lCKOsvkyhVtTprO+YpcaKCyO
i15MMHXDKk1/FQUYWW1UiLnp4rQLE4M6qhSHXW91LjHJJwqPV6ETgnJfj9AErNF2Is2iuHn4u3yL
HylvRqL+fg1iyPJX904zmQj0PuF5SjGVUUT8KfPJIfZHQwTjZKWIIUHTAxuC8qxTBCFxE3KlJjaM
2pCBCcAOSybe65eKvQxWsvR99pGPSRhV+IcK/DDKB9KERqM7Q93n+AOYDh2ZhfMrhzp21b8pTECN
f1/ysR3O5xI2/94Hyi15nYBHu8PU92+9vK6s7w83eHxo6JYE6jjq6nrYjqEp4zDrLcSNFNEOMUhZ
AU0IVdiMKJUmmK5HnEiP0rSwYT/iIAwBbixgZJtKodnDtEDb7bGALbH2rMTU8o/+LsKRFpB3VTkN
K32/exQl8VXzpMVFRp+zUQNlGVfGsD9bgcslUcTNR1+0U/EwcBpFrIswfrP7fr3euJKz2cxNp5o7
w0ruVWFnWJqLOWTNkbhuQNHcV9uQrdPAkqbmIq70/461n11tpWTG6lN/NrVXSastAy71VtMDXvf4
zD8eHWb64F06ibUN5xZMnk3OqTRk3Egs1GiHd8GktTJG09XxcFzZZbnOlLdRlW7NrM92211hXJC6
ow0DsuUoaRsOq9iSh8tPeswUzoQ6+ZbT8gYgTlt6ZLNB8jRgfNtJNhdKI0IRRhZdOu3d6Tvrsfp0
7Hk88efRvgiALEgRojDBGaveB3jXN8WiiO4UNQTc7uFibaJtWqa4qc1mSJtX6ZpPaeeR+87PyaiU
T5my54V6g0NyA4erxMKfapuSrJCieXVaGFga8hl3opiu6i0sAplHvWgiZj5cyUDGlrXgLnkzclaa
aV4YcsbiJL2tp/9hRCcHS/CdrVV7Q5MvmZLy7L0UMs+XnOc0megNO0X0RBg8ogBV787Nsr1GixVy
cz+2RsWwUHBnQ/z6IczGr/tqcbrYTm4KW1oPwwsL3/W6FYSs+abfwgQR5S20jrNs5GVC8hR1Kvaa
jlEbEmQw9KMCg0MVC4S32OVS40ZyQV1oQRcusFFwV2qOwv9rvq0alLCCPMyE8mQzVkmTWyNbMuHG
1B6yXfnP9K41co85Ci7pkHd20hdKhzPCwBq+3nnFkugQsRvC6CXvh6JyW3XA0J2oFAEXBRE9KnHA
16nFzrb2//ZXbkOeiBxtQ8Y3jCskgnmsmO3/eFNYAT4B89ZDb9Fs1DdhTaMF7UYDOdGefuriRunw
ZYBpjP7D3GVDQ6t/p+6d515nszcAU1eg6mUQY33dRpD1xqmw0tVp8g5arOCEhzZ10rnF7/lIGZXU
oH10tC5DOvZzQeJUU+22X/oPjNL7+tUKqCuSlwBRqb+za5bKk2XNEgPNurjmKGiMTXGbztllXYV1
8tpHXtahHPRD8zV/J5544apsMaPfeOGkonlYKuVq64CNcv7tTaF/itbyEARUMakugGKMOPMTnFqC
Jvt8bO7/3o0/vC6gNMGKUnFFz5op46a5IZ7dNqH/8zDeCQ0eLtUd8zun/py/Qym0afmHZDkqJN3I
WuBNcmSUTUhyaUPhal5w7PKy6+sIbIllRcKX2eU9GLTCbJ6ao3rQRlda8PBa82s0th1TFhqw0guZ
ATHNT0oGZFWoSqpRcAdUI6+iGLbZ3MTkteSQ1jC9ClOF9E2g/TgDKkPTFEWJJgIFiWetvIenuqkz
ILyRGZuIRf8/qsDynjemxsSny98YeMBgsUeVwcgQ6YaBjv02DO6+Ktq7ErcQS4Fr5OYLK6y4h57d
QO6p3vMNlhd7cW1jw8PwsCcW/nDixriv93oqNLT0rTs2K3280CVRYAmzgIii+uYzT7GN1UBafMzh
Os8PvZBOiLKanZ67TffGhSNU3PIwm0OTTmhrGNLkmkIxvMVCMR7qf6piUISmbHpbxNUdMzUBnXy8
6RN6IvGrshpQf/2wYRz7BsABQFOx6s9HWdINjcoUwFzyBqjqtmnRynMUO5wH98fCRiJ20zkfGI4b
ez7OflXYPb02J8+1Q7YQHA8KmP3MTQ5eMS/fO6AifljYkCMuUlHInr4QtvzTIqdHcb7qoJOI42Wq
onMpHHN6hLi1tcYJAAWDLiVWErQTt4A2BYzxT25wjwx6LRtfFYnRpzW+rAXL4awk4PK8Q53/msn0
YbOc1qUcbVmUaRGHHURTBrAnbOEF60H0N62O1hsoCG25CJnx7BFCxSSC9GVnBqFdUWjFmfH7fsgH
jLERZ/sFZNAunYC1qzNLOcUcse40I3eYq8Z1RWGGJlnlsUUnxvdc4zkEyi4AA2IidoONrGKtuVOO
gGBk+JgnMbcIcgVQ+J7T8JFeY8uMUEGit8CXa/DBeM/EbskOHys5j/RZ9hCBscMdljrcZ7sUxLc8
Mr7cz750+wQMmsURSFsqtMDnXlZ+1H8Zq1FeqT7Xhi9Yx4aNGYWAARmnhEMUfYSDDvfNG2tkaV6V
D13lKJ68iQ3iltzbZ1YYDnEM3EtYq4sw/tiCDxDlZvSwy+XzqFt9BfHXUugsNOBFFZYIIu4dNSNG
fOeDijPg1u3YeLFDcSLTcq3AftNTCkdrwRcy/fY3wwkCebLoc0DAYvfHGqd/9n2+YJBOOz1eRz69
WvD3sJ9p4PuFj0cr1TXoDxic0Y5f6PgCh47CV62XlRI7+ElO1bTdcAXH/qcWZGEtxyCE9NnEINn9
TUf9SXaf+NfDoEsV5UlGjbA6d/j09C9O8zN1/BCn0fUQFznfSyjDuKH7xAPhqnsZlqaTKjx5DNMr
1XPBxPmaRNYfcHlrb8ZTV7sYTdPBwblaj/TZPW3XeRTJkLKc0TxciymTd9kXXgo5RVuFxGK9fVzu
K2nxKpIDPyaaBSYp5VEXdzkfTMtOXM4waXGJUesjvcFMG5nI5BODMtoT5EJeJgfdF5rFHbfY9WeE
L+AiDdPXXXnohj2IlHjdWbZ9kqIeazFJCtHm3gHYICY1HKBjB2wxwTuas+V1pw7yd9VPm8Rd1ljv
sEGZvQo+UDzwnnjDE1eGI8y6z53SSyopUtS4XWKyfRMmgntXbpyoa7gJEqvEnkkA2rpi2TYOOeDb
ApgWGRFmQrh44Cc+nXPymFiCVT4LfExX3F4+xcY+ipUd8XDxQukeA9k+FgrWGxMn5/mfNlpjZjy/
/RuLtS0YuMV2XfTVM4ZG8tF4q3GP6A00E1k0DnKn/n/N/5T5J3S1ko02PLL9qtmM0TuHNJ/ZIW6/
YF8348ZUyYb6PchtH98/F3kyssPgxZROV31etp6tSasfvUK/E9kaATt01/2EldJ4qZXiqBBGdRVa
0quiYlOAf40UPNHc5io5mTNip6vdc3OaZz7vOfebNJ6hSLraqanJlO6J+BWHeJ07mXl2vYTRfxCh
P3ZlmVcfdDeD/si6t/hoKzUH5GrVzGWh8uLdvZnul1DP5HA/DrzBHbzTztB1KLIDvb24vPyKs0+9
knzkhRspLMU7NREI8auBmmhyUC2L1M9DWnMDxNLHLVFSjFPf9BFe70+JnX4FW+OOEtbwL55H+5Vu
al8xxLxnGwxrKoBowkmE0yh4O7IVGb2UmKCJwE3oIE++lD+C01MoYjgfac9ut7AZ6NCKOBjNhi9M
FH5RMWWqO1Pq3YmwZ3wqniXIIb5tsUnXdCS9XAs5DixCTuQOwJ54qqdct76walIUTHSRN0n3eEyH
cOAuqdTmJwiB6cpNuiM/oii0sz4qD1FYlu2Fv6wmr88iZap4cJndu0uUl7xpFnHh4sdKfN2kfDCU
RB4LwbU8W1O66ja+TDKdQ88aQJU5ImlUS0Slbs8WDUkMsA4MNI7/JdJ/AZCYd+fVnLVbfSdTNRmx
3KPC/qApgGkGW5pFuaE8Rltg9GdqM4z/i3yEoif328fJ5ovQbt3+pfuUElFMgBqMZMDkiAkbD4ke
LUQplZqfYrJt/x+Besk3z68Ykp+C1rUulfGi6PcdEu62qDZetQXNiqbX0zIYKcKiiO0PhvCnsydz
zXus4BF8rq9wiRkErRhonv9HE90rCe5tc59RRMYoTRR52tc1d4oyeSGv/zD/fK98xLql9uWBtbyk
55WPvApG7m8MxmFu6xHrgyji3dqR5JB1iBWFBEuEF/RfdJN88+WfFx/rOztKj06aRjJdyDevIi32
gjflLCBfXHwkNfrfKR2kIbnl2bCtlyrakTNaz8BX4LuxdGaoJQuC7/Qh60y4plsuc4e7/2fJUCih
n3lKCAg8D1u9IWrY2+AFdaMN0kocibKU55LhpRAK3o0Au110Os26z0vtklBROaZGIpsADVylCqql
9N2Y7mIJ9qDwK7pF8mrnrCVWjHdfD8HPm0eTdPw+nlPvRM3IbAhAAjAnHvMl4oLCjjDFp3pqPBWM
4WIoxfK5rehKxip4do54MYY3CNhCUmmF2h3PcP7LKnCZTuqvDP47L457QSnOGSMDhLEkc1EOuEuJ
SGAnycA2pwfY+0e1tga45BaL3v68WgA/+Cd2baqOy9xhvFjVjQsjtADW46n5i+fJnX/zdApJd+yM
zo1XUGibiIYvvN4CpmSlTI8h6YH17M2gaXjHtZ5X25sQQk79XBwVh56Cv5EbRQheH2fHOnDqDZsy
G+2HMZenRELnuCrAg1tiU86+8us6Q7mgbs9qfG5vIVEyO5w80dNzxKo+k+fiKqdcX1Lx1bU7IUW5
6WOJX1259gO0m1Z1Le/pUJeka5LPCBBH30u9kUACJYSs91Q9WD3oxaC1oRSdj9vnRBS+7OZ7tamM
inHbQyl3Zcq6U2Jy4AfjhTM7wGEOpAIeLXyzL+9D1BLqyFcX566XduVWw3rB0Vhl9PhRb5dGicIy
esUJwXhhiodby7oP0Tu4uUlvH6BjTsp/jh+KO4q1/XCtOMxoyv4ybgLEE0TYYFKGt9jH/1ESEOaw
HQ8eIh6ZYnAS3+Us7/QXR5/cLdSCdnxb3aZcqTfBSckCxct8YmB+H0gKNiHuPAGozI8GSoj7k53J
mUudWIBGMIl9S1ylcbUA48UwngeHb0DAFPmC89MlFa5ADY2Mtu9AKWjZ//Q1HwNrGevc8KFhsIYB
QNi+yZTpP9Lmb9+rL1wWZ24RL7SufGlSpKUYJJlMmrZncPy+tEAkxZ76DSZK4gpObBaTMXqe11l5
Mtu9e7WBEc7tW6q2JXaZKcGrdAXcbNXScnN5JXOUX46Pqc8nPmfHvA76UtcFwurATBUCxbfxCJd7
5cPXmz9KkGAB0Vq78dyxuU6CYxgj1G6sveQ3M11YTwjFkxzfg3Bq8ifcf2074RxhHGWLKsyEw3ro
AoAnOmLN88XdDXY29cclUMAt12HTvwzdgmXSiSztAE2ae5d+QLi6kNqymB6+fcn3/RU8fN9/YUvv
3y//y4scMisaMC8KilycZqnA3n9XNrTEupspwjcpZlHRCbfxVTPnknLDMVtcJl9O/uJs0XT7D+kT
8CM8vbd711CiY+pdAzx0R8ZzcKyrDYYOzDBnCPQJl1lngpumDCLETH8yxacfGHz9jPfDHfFc9XUE
7W70tV+3v55YGE5VziwqYaaVzdTmWVX2b1dIV4DE0iff9Co2yERrTIRsMzNXcIXN15b5/Q1NkNPW
3jI+wSM4+lPtMrSCWYDTwum6Khd2mw9HZaJ4eug3UYpMpka+et8RM2xcx38uufG509gRo5L/HB7e
oUM5Vq/xLnwaTdOkQkhMtnrMe4mSW9emzZEmXEreHYpplqnXa6g8iP3j8ezP5liFRKRRPQJdygch
Q6ZfO/Fd0IQ75Qqaj/HIcCQ2bvNlsymKKSbKQNID7fotaQQ3gpwqBl1cOlV9/JSMfsBL7NHtU8o+
YEx5RZ7BYpJ7TKp8PF5aNZOyXBQJBAIdiD2rCtjscaTtML6cCf7uw5+fF5BftD9CPL7ovBAplJKA
oNndu8zFLmKmR1U3LssgAQDPrcm8AJ+7iB4pqQjOGMjie3QRIz+Il032+xXLAvYY42lIO/2LYzu1
RQu0kzBnCSDtv9u0jfMupSSPyY18f0nWasiCeXAE7Sca7/ZV0sL0XUcCVWtlRU0Hj5gk8OcUPfNf
7OrQItK7Ot1yVXtchk4q/kJTZ7vnWHoI78fn1wjZJ8ZIQJaBkQKCQlzXUN79UAQ7EjFnEIIfyFvB
DN4snXL6814q9Vw9FNWPqZZvUHRV9qmDntlNtT+hLb4i2L8K08tCBQoNIVDEWF5uMj3rAEGT7t7Z
lc216iiAdc/RgPTfL20GgsN1u0Lz96bGWW6Uu0rAZjw+1ZQ0S5uz8TpzpjMrvEYp/3WGqcspAs9+
8/sQqxvdtI8xdR85MHcmdxH5Z9VA3VafYWkS6t0yT9WvCjPPHixzT6Dyn9cqlAmfu0TpcPB6pHHF
BWdxaBpeQ5BcrxaWZPtkWz5+gtx10m0aqIGm9jf+t9Zg6NRiMrWxsvuJbO0yM0O1jlyptjuZ3k70
gGKFR1CQ/qboWVSlIrWeWzY8Dmvt1Mkmyq294InZ5S7iV00ALsm/nhMZwTbBXkDBQAkuEApyJ5jF
VGjg50tOzScDHzKuEzSc3o9wl5ObgR5OhdJeHtqyAppOTb7CNlvZid39Lw4/GKAJkof0k82QePAZ
6BE5BXv6IoEsnWmkQRH3KGvi8n2Bn4/gQRM79N61kflcBLsEnrTmFak4gdRzlyktRju5xs7Da/fc
lg6gWjWPZ0qDSKORrvsDUGmIKJn07Royb/RBXpMiqHZGfLDmNXUEp6uaA3ur8up0RRn9kQD7J2kK
iBMLN6UcmXIm2UvasyV+3QO/dKjYeK45y6/nLow428Uf0csUwUgLCMGqP3IciJ0VMnx8X7BXiEnE
YvsY8uKq6ShE1ZIzTEF+OHy0ECQwcrNn+gtFXlicbleSCSdZ2y9S6Xujgjq9tyz6qg8HhPygPePL
AZg1LzX5Jk13PZo43KDqHqKr0AY44+7TG+0cyocdr/AcMmwnvUxqCcHaF97mHUTLqRL9n6NHXGQN
MFKFKiXcELCV52aYq+mR8/EOGIqx+OeYBDnYe1Kp8PFndVppZ2xUA9B68LFup5CTFU1j7blDIyqg
2jC37cHKlkzzOOaoEjoKoA9AxmcqHumfHLEt1tbzAHXP9Z4SwLyHAwi2tc6MEDh5qfemshk0zh6S
3NfNhxUCjENYnP7z93sWXz2B7fOi93CSoSyVfQZaNt5T8VcSW7rbfTgAwtWnKlApvPprqae9irAq
gF6hVrjmOmTizrqcU92tHuQwi7i2j1fVSc7phkUdoOXazDnx01CQUxU5p4BD3K6aMfruc8aApJx7
PZsYkgOi+PtQNbN4d/R1LHxOanV4P/mzr9TprFQosK+EKxWTMuD4poIA3+OPBgDKpzi7OwttAHSj
mAbTHs4v/pno0RLd51HE8kq8nW+y9xEYaMB95SkKjcNP4SFBaQIw3sl407onA5vq+/qFLjiCmuX2
Qgy2A/ogbD4TO86jRGS+uyaklfwFAHOwX9C1DZ/kTRJsLS0uy6fRXr+AP6oHXTedOG4zh1S03sb2
8oszluX0qL4MKG0+SKf9fgtGnTWOME7F4PsHBb/GXP6+sKRzn5UpiemouMdvTeSJcRZYF4PeQVeX
9o0IGdrfpLIXaf7thp8cAekfjRqsyrWzqIAimKmCpsc1HJ6kpHNLQc/khM0SlkrbPv+iEt7XFSlW
K++q/kSH5GX/XsE34i1FzokHNA/2d0JJT+AmWCkpOUnXR8m+nYvKrC/eD1Czw9kqm3r9SJqaZwHU
/V3z+ZDTqJBv+Fn30ZVw+soYfISEuTBnqVQV3fc/uYOEQHi9nGagSSwPdkvsiD879JzSnthm4vBJ
dVqv4LpWLNE1PaMYqEy4ckZmD5F424xS/Rob7xFhh2Fh2LBSkPtSMf7iE/9P1EaOIhzKF01R4h93
yijAlJIZjn5FKfs5ot6Brseh+6Ko22o4284mvccvNKd9IRD2o0c0bBjiU+RRkgb5uxGLizF/5mpH
AF9aMUQLvY/YSh08gApmgRvGGl4YxOK+UJjE4evoK42el+z7HuBNiQi4oQXWRMm4uJHSk91ouELy
mvy1uZVtYXbaef38oh9axXkLhWkiXrGRiXSv3ci1MpYwMRR9t57GoysPv/w8e9IF9H/a9yp3Rb3E
Q94oBZc6LcFMjBbAl6snvO1AqyT4Kyy+YKK0vLvhOqymWUw6bNHQZTmQsOYdTojV6eREG7BY2KVu
Cqdo4goD+zfM7feyiwTO1gw0muaucqOnMb/sSKHQRobX1/E6kT9+4c0BesCOXatB9RJjk5B9yr0e
oBlnWZMWZzlRCZT2nHP9xRPCUMned2PpLGDoKGQe2sJS1bajW9e7ZnDFTDd/KbAVq98gWXnEDXqc
aVspTtjS9FkID4sAcQeTHGAaGpNY5AQA4mHkbH370nJkmF7UtdUeq8nhYG+qSt6l6Kf4N+3/tjI9
JvPLlGiZTpH5A8jCYwNps4WJvSFhNzTNr40LasoNoeNf9sbAskeIcynHoXFwBdTsHOPeKTt4QfMB
2Pudu7oj8NgUyxCRBGD/hLVZQol5Q+iFuSz8mCbE33V/efuuojArbKZSX4fNfh2dZa2iKsHIOcLp
JTKeDnLT60z+HohJn1OqtJ3rRvtEuoh9Qj0SRvg0TZWweySayg1WBSFjwACP87b0lQM6iZiBkq8G
6KNzi/sErVqsEq8sYsk2AH6c6gErNvGXS/EOT2W6zs3lmFmpwVs3DxFaXcYJbYj2c8FC8R8/Gypq
ZHOMDy+9fxTnFOPE71Ci+9jc3tsX4ZhQftIrJTmR3JkgXcS5pP3L5EgWVXaaQemqhLeXBaP64Bqp
yBrkiGftXIaltNRfK0BLm3l+iKs2dJxsG0aNVJqq0x8RTdMdK8sseH9sMznFkPTARQDCItSajpHj
nK+ysNhgkuNSMkkbkAFVW0RUhY7Hl3JHBPxb8pqRgViJ0kO97Yl4G0LWPTvB4whbrB8g60urk3m+
tvn7ecap8Ot8hUzIo6+uQ8DIra+jaGmTDxoSrNHs6pM8CnGBLsLtOGmCRvH69qwPojuYRjydw1ku
8fB4EN1Q8Bc8H8LlGHQIn+Q6geOTXmOjmlz0krfVe3twowdLLPA/h4veEYLA9aOIv1RrIf3SNfa2
mmG1mx3sTCalPLrPnaOMUPOv/7RJFR0EhM4k+ivGtyTST1DMz9YHCGNhXwh1jqAwizr/DkJlBG2/
tVF3sXPhJIu+gJ2duQYO/MLpvHaLWAxeXgLafjNuebbZbtoV+hzFrEWH01YUNb50M3kgvhCXz25b
tgv5LR1IkDr9VSqFIC0/QOFjOFSDxqB1m8LzOACCO5RklhNpa2Fveu9N9AD5lslPFd2WKDBk6XN7
U0x9ZU0sQklyJyqpMbF4bVJ38iklsQ1ZmkwbJNl5iDUkEpbLZ143WYFbdm3/hwWZzs+0QVaaJLc/
iIVAyv5BSiLt37RdK/QJTkI6P95MSJNFtPbyhWzH01Ab9LwOc6fGO/cYlAkiZhOpejwoVD/XvEQO
VoLwkgN8+oz2LAMZcjejnDkpHogSGANKRjrOJb98Rhst/rSd/h4OFEbMrQh7b4KxzJ8YZTjYYErb
tdDzwUJSJ8raBYJ8UyIqQNsbT18uJ4dBvb+Q6eL60lsJ1/myJnxClDOcMnv7JNM03IvSCRrpLTV3
Ylq5T+uP+hvV1VrsjR1qNubJlu3v8hkLyR4w6f3OQMPF41mP18+tb9JgDONmCu1aNVvAupmxA8U6
U1I9hKZXTQiDkQljLcID6jFdeT+BcTTm733Lw3va56LPNsBNIwjQw923owyA/PdbtRqwfVgG0R5D
WSS17J9AX8V9BDFDFQqAJW8vQ6kWfpMxHQtJLFuke2AaiCCF9YiwHipVSHUpV0sdTVnb3lDiZtwi
YVSVIxb6drYJ6NU28tLt/GNkG7lpUoPcJ3vUWA7lNrkbGzCHTkWYev2UYrmf7keRa/BUYGmYwzTd
HwVI25gHJj7jLPGMIqfm6geZq4alzDACgL83X6kZE7H1Y8j4WePh8kWiOJGVnmalbrSsOPgW6A2H
pVOkMmJo3qH+zvZbqeobETD++GhI58VjFX1x871KcFLmQsD+ch9DrLrpA7ZxawAW2npMxRf0xqr1
7glaOB7LbzYBXagy5SkR1oYdQsOIS5wRcfWyT9fZJgD28cuwUwlTrhgM4DlmRKFywNq6hwqvQNTY
O6RO+P/183/wAQ6Klc+LRkJcIDIP6heI/YNaSuI9ZgRz5PgpJjj5K3w2i7TUb0w0F8gFPpnARSca
CE7gNxINHxnJNP4F2sk7B7wcOgIN7YLSvMlK6qxii0W+FcvmiMlKHPfRubLxSi+fvmG7dcLdqDFB
ulC7ntsFAxDbYxxYiifx9mj/JQwetMegPwO9d03AKENiFM0QkOtVYgqFuCJ0f+ZnFcNIWjsnGnjx
vgRFh65wKHaURNye9k/Zl+61hAH/+Dyl6uAvZL78DJIuCMFSsgQ1hqnge7wxCdePD2TcTYokRJy1
LEmapO/w61uE6iaLY7lGsR3VISAI460mcrPwugl6IenhReeZdF36+gCrqRi8OcEJyAT4/aCEtvCJ
qgyfqCR/TlvjsgfhUToyFDM7bJ5DACpGSitTntNHP6pXMwHWg4TyEpJqmc6NrQC9RziKirA07gFL
Pk5jWJMj5WRun3vVuryFirVC64Yzr6kv5lXGLBe9j4H4iMeqdB1imoeYBixhdaCxkjX97YzYsG9U
x5QTqzGQCkY8LC53Cxy9px+C+bcIadp7hUo1bpEMcS8bn/4bOU1BR9cc6VnUTkkwXUbDt7byoGhE
Ar6rAEfIfCrBiNLhem1Vopjn7ogLrd9gqUBhvOl/Y8jRp3h3bBWbjc1/hnUZGf4fVgMSf/tm5CYB
IjvECOXbP8/0tyPat52g9QqCNoMtvtTRLiA+/dP78vPcbxPBydzW4dpdZlCUqXl+L/pf14U1/gPs
bjNfAmPf9f7TlWZ8oQeOnvSagZAE6eFz9Ly/Hkp8hBwmObCV1S7b1/iXIH3M+jfEH6WaFCInWiKy
j+AiqJygxeST+HtpAuoYoi/VPPvRRCh1AVG9MUhiKhicXr25A35IuLIfiz2r8ussTajmMrNn/nBq
+yqBSuQMjNAmUR4cvs8LHGi6h94WWQ/dd5EMtX6iVO4roDqNhxC8PP2q/nhh1tgpEkQJ+GKkZjZ6
8Ut/iZ9mdI0qm2Dkaxqxp7VDcew7wJsM/zC0yJwgE+J3ukTWymtBrriZyQw6jzr21ZtnaCM8ruaG
koYDxTlecgszfDaxgOpc1HE8TCuVvM31Ulw0ToqZUchsXpJRM+ycTDBldfPeiuMvEk4y3dI5STzF
hmyZUO0jWf1LbdAfVo5zSwLz7aoUd9ClqPmpvEvd028gamUSqLVBD60udIzj2HxpRdolz1qBLZSL
W4Fp+NChw7fyRxbHux9hmYtvAEl01VaGbsGhZHYA8DE4XFeIPYIWHIwAsuADsNjXdH+8QNTIaqeI
/79OVjrfLwYP0/5gCTrazHm/y4QhFxmAjtYWtTI38tJM8/YbbAs86Lx/0mw3/+P8UOYNO95r+cZF
yptjEIInGh7KpWwysz5P8VY4LfIDe93G2PicokT3LNElYv3it4o7XJ2fs7LLZ7cFB1o66v10stAq
zct7sbDeus3HweqMoFTt9DHd26UMWO/PngTEwg6Y83l6PvKUz/iz8+YJb6Ebc4zz9d8OMiKqlarM
xn8hzlJ9BSpY8CyPcpxg1jb7F1SAZ2Zh2hlfx1/gqt0pvbwc4z1/F7tLmL6OksQW5nj9G9z+z4Ug
lxsjRt2gAs0C8ZoeD3yK9o2PI54vOHWMIPjNSO12GqKnHD3BrbdRPA+hC+edOC2i7B3HqVrqwsS+
x7/zTYZik//qzPVQLw3/2fJKPkztQ9bymMtz8AOxYLtI4HtcK7q7SIKw660BBTN2l/nvZMrlAhKa
pyRx8N2H8J+XuTYpSbCY8pbFj3nvfvt0VEw+zkIGqWeXITJ1Lp1zd7WkeFbF6pOPx/CCwFtZaXjJ
XFM1eNrsMB0CK9/mFqyPp0mwCA4DTA/4DewRV2+DelMZSiK7HB+6RGBibj1HoaUORliqS2V1ZnFD
oGATtYc9svxwq+TzrWUPFHvM7DiAwroDcrK5+80QyPp1D1S2+fNVbOKS397yGL8GPUr4d5DcbAia
8fxZuzaBWfmhRZ75RNYl3Qud7BePsUhTtrZDlmTwVGKd1I44HhZjl3IxOV1l6Q0GlkNHNiNHvmJR
2XovkkJAvnDM+bBaihJm4m7TvbzUgjQL+jR230jcBle97eHhERBCbDkT/gFrWfR4SbfZDk4Cpm9z
e7uL+R0vr7vOGNlzhaJnViSwU46g/JwfnT/oQYQsBRxx1mk8IprOqtRsWmNB3mdF4mC2asfbsFYk
+8plxWQvCPKv+CmjP03y3SBCWEOp7VvcU0FMKdUQSNYVJ0BzUD2EkAQvCpVKzo6FVuF7ttG1Vkqe
4lEWsuCq1foFSjey2HNEVrg9FcRJgZlCttfyuc/vdAcN/HWFJhm39Io2ZkC18VlIZWdAR4H7Il/F
Ux2uA/N75RjQH50vtDWFu7fib87ttAfXi1FcBCkK5L/0knXzcgG94JS5id5Ncup0L9e12131ocjZ
ObT2hp0crpNUY0X1JSQxDV9VOCF3tHGT/AKEFt48oqvqQ0LNLeDbMKly3cF3ER3ujPnAxHAVjNND
ZNtvA8tSlpp8gJmFotWDa6d0FvBy6UYPLadJQ6jfIDNU8sjTom8ZWFN96v5SV1qZoJImhn/36mJj
sjEaSMisiRjKa0/PKUP9kfGyRcjYKs5hNDyUZbI3ZSWYrMm0iUrhiW3asjn+O3vVsNprGFlH8Lgv
5pA+z7ofqfpQIWoe1dvPKVcNFYuDaHfMbdSA53StV/+PPDm8CH8fsJjmKR+i2NVIH15+okWbRsrH
+nZKN7uFs4u9nh0n3bR53S63Y/JeZnNXnXD1NKxjzIVk+/9IkvOdLTuG9JuXqsQoAkKfKYOch3fd
DCL9n2tgccbIRGzns741btgO3Lm/dEjPNnDGTSzwP0jOJUSITeXvg67Dh7g784dGIJL4ysxbHgEI
XbrfZNeiOBbVHFmlqECyAJztU+cLDWoAqjt1OD+nsj/cdEJ/2534rIMpBfb1RB/R4KlMpXOdLqfr
3nT+k45fEI8w98fDrRbMYB03M7mu2axixBUwJ/BA/ScPkGjLaJ115JyUfVfYVjtmi31GoPZA/Dsa
+586CRHCVXlviNAxIPta8UHKI2lVgM6QIW1LIaOrPFNgJ0x8oMbf11sLExSOADsa1GDVfMRTnimJ
OuugmzGFZcNpCvGfC0EkacrqrEAfUGLdDnsH3Dp7aIWPG/q/RE0anRts9xPIXS8eTWiOCAzmHB3l
250gWcbSW/pKGiu0+oM8pRqBO2WH++sDA8SBJxD8mOsk/aCAM1mqL2Xf4TY1yUUmluc3nn8hO+na
gYVq8KdvsNDn2PdBb2TEMm+87mV9vLgfDRLWs/4zZHq4EHyGQKJ1x5yLaPs4VKnHTDY2khrWYsAo
ST85hWXuIdF9qttbRThB0oYJWcHrxi9hX3jCD/nct3icUSs3FFMPgrUlouLyu+NPj+TtM5z9Dv7X
sbqXSU/xzFux+E+FY/6AN1SRaLUKfmLldwIkNl1D6/mqBUnOTCAfzWotS4cfytJNoQfpmslCeQXs
HsCbeqz3xHHHvH5KfVNX1sSkAbq0K0URqIqt2znKSEIM2qxVa/WB+CbuN8RHi98psd/e6Q8kpxWT
Cqh66oWJ2yWjH+6/vYKvCPmsKHYXLcYwWpVURv9mjNkegEjEmzmsUfX8LCiEsIJ59GmSXKAjSWDS
rs/EXDkO16iRrLS/928pUuRf0PQjbEAQLZz4vB+RX1pq6U/+HYZVXGV+hsrL/NqmG4MtnJFo8b1s
HJAatn6k2MtT6RKQP946dm9gwB24BOjSqoGmxmGjHk/WbNyS1xrvlDbiJM/cGq/LCXuXlg+LObrV
ZXLTCdttDlu0LArgoMBUgetnlS46Y4Uq0NXfCQf1HN+B+T2JTDLySBJByUrM/IjU9t2L0UH+K92R
iVWaRgzYVQHJVq+m+eXSh2t03l3U/HFna0CP8V67Pg3nhvMMp9lhA4oxgauC6WvZfde+XF/sBBOT
+coGNHNlw/UNU+Im9OMH6TGixsuSreVfkbyhKJxEoO/tx1XpIRsgQeYXykTjrgO4DNZcGR3CMSPF
kzOxZ4ob62KUObj8ghMyoSOsu+mHIrLChXtWWB8uevPS9O4G87ZDYA18iW2HCYl3xhBmzz4HJtqF
rSPV93cP7WZYfF6m/QhJDoPtKBcl1PCGtr3AALd3hgQ++W/SkLItbDUYtoIvyrvz3uANH/COkEL1
KITzywFY2svRapTKeOTM+qJeWXhOjyC8OV5OBSe+I5lqXo5TlrnRuDrJU8sIk5vHS15mnNL3q8YS
Ci82WcQ/rd0CXrC/+8Vry0ZQcrakuglqjCVZnbeDuXLQdfyNLwhdMsxFf9n4zpvvTs3jxueGQYlq
zGzyzicGiXxD7MRRAdhniUYA9QA0dKX/uuHBxoj7Fr4lzfLfNTBIjxewjMIH40/iBlWhi6Ja2Q0t
P4U0PfU2XXPEqdXF4RS4KmnNsFmvbVRrG6XbwHMHeF9IJLYoHcBmS9MWU8IuEG7OCqDqZt0Ba0dA
a0k05U1llVGV+zpVBRMpMD7PLBp4NP+Dpe1DPbdM6DH6ImrHbyMxBJNmnZ5c6p6ybB+EJjII2USP
2CmUl4BBfIrP91miwAl+1B79O4SDylLiFcPPD5bDBf1Pj11CnRCUm+2LQHJel+Ua3JCMrXjMw/Fk
7WgCl/F0iFgyJvY4J+FYAxojkEcZwtR/xjlKcBG/cQRFSQVqFQdxiEakMzQP+hv+NoSROjqywFRd
hPaO0gN0B6OB9xIKBmfClTXBKpf+b7ZTs4uGPJV+5Cv0oVNhViE6gYi5GKkQR+zSpJsrkLp9rfVY
4c7tm+x3OvGLOLtPdr7KNsFDziDdyZ1zeLVYCD43uat5BlPaYih0xAbFsgWUHK75/PjhpdpEFn64
pb+6MFN08DyzxNYwNzqiO633P5HygzbHxF5a9R0YSIogiSVvz5koQJe2flmz/EdZ05nc1QIs7ob8
2MYosRHBgYx+xp2kdnfs+NkJKQwkZ8aezYLlp9ItWp3kIxXn2jMA9zQuizL1lWriqEDRE5ACjYaC
ZjDxMvkIFtpq8tQASw27inKT4TEB+lnPs931HH7th2BxG63n7fR5VsrlERxQvPtxFn5vPfsiviL8
L4iLsIK9kiLuErYC9XIqwH7VCoLgbMyN9lL7IMb5Vqpl3JdmjQzybk3jO5DEM/7cLxtgvPZLLoTi
msNVvzcpgkfhZ0CsyDtjQVWAhljyvxiYO69xkrjB+I3D0NmD1ePxivr+kL29MOQnY6yRxAacVvKN
YO/x40cfV0FJOlJrcNNkVpbfP8Kmmpf+5Ufvpa8smkzTYPa3HlnEoNFbExL6YpsPeNJPWynvplYw
MOg9rnVR/pVqJxluuAJ3I7pZy0yjfndo3ZW+/odJjX/er9KpGMrndVEz7IUcUZ2SHLhEh1ktLng4
EwHQGLyg4z32r551lKjzkLDib/pa8EbvyNpghCa2Nqbher1anZstOuDCgQwOZzfn8xDdvrzZZi1S
/4s9FAoR+H/zM2xXukKhcwzqIeygy1hQRxs/K2kFrmJnZLEWDQH5F0s+pU/ZlC4wYHKP4CNgWNbX
+OkoT8rQNoVM5S4baHUAYIf4WI6UtaiYV0389qIizksjJT7FobW31KUAJxQkJUV9O0BS+pH4ysqu
THwsFwb4GnEQrOPxvu1TLUFFrsH+gAsOH+jQkEt6LQaucsdrlfTT9DrRJIIWPItqqPXzslJCLpur
+LpoMTrimkZe8iMjkFshhfCDxkv9PNB7mmHYzfAvCKxZ1kxI+rH3xNOv5AvDLo8hThIhGaElbKTS
mq/tJWATAsQZd9FLZoEdSUFARUOsVPdmTjAhA/g6tEsKNGBLLLMBFpvx8CINTskNZoN+lqV1mPyU
AOu+Q/FGXd+8Q36S1IGF2lQ0+jWQNJQBi6CvRIJPlFLJteH4ddKGcA1WwFosCHVU3xFLcWV9DSvF
hfmKXaEWJ4QkP8ahwPOtK758WfzqAxDnFd7zBBLX0tiMuAG0kq3JmEm1HbE0GPqy6S8VLnMhg/XK
XSYIT9XcYbWORKaXrlZOBSHnK6ZIDdJfpapp6e+qrOm1swrVzOy27TYMHEwPdTa59V+ZQ/6jXXKY
PSEJhznIIkYJrX0IiS1tHPZA6X3C/dBoiChlbnA9n+cvbLLARajAfpDkEsaKvRHhMWBLg+5VWIAf
Ig3C3swEzdmImX7V1HYwXdqMrTl1zMdx65OebbMbN0c+HzpbPrdkExBOGnhSiPwrUVDH0LHLrmLt
lwZbJng1WM+RtUE5XolSYFBHsXM8FnfYU6wTHF/y0iphMrEev1SbcZzS1f7urflXr4sEYHWOgS2b
k2g6sgyhaxpVelrNDt2w19/qkr6UD6SjgeuAQDyj2tCS7ZWauy7bVKmyVVT+1owgpYxq2+ObDwMh
x1hiP6wdNWMbBvM40FQs+EeypcR1wp2g26bFuZPOXBVVIT/X7jEgM0L3I+S8H607mL6jS5APFkwR
j4JgHjHIBGZHfw9sbR62xbv0cn3PGF9wz56VMfCZW7LTANGDKntRrQMtWG+rN8LnHB0n/RBL6JaJ
Lm6WLs4oQtsgxaCnn8aujJA47AR7kf6/06qhpM45OBTQTG8s2Zw8CyBh+CFGZlY3eiV1JYJUAhce
BQEjAmsDzBHi3g9wDq4mc3ylpwneo9XxCt9XDV/nzVyMELRGSfvYCBkCBRkhUXA67vlS91V5FOfQ
Lk2oVR8gSs+r1dK9IW4TbvO2KJsXMquSkBopM0q30gynTS/CCialihIOlttRqHuv8tM6oNrau+Os
ARzGNraZdtUPPFabYdtS/B5nCerNx0lgnA4UwHhvgS4ce8QGJzYj0KCbJNqaG3DhJTFJdqrqdrIE
vdXfZwT8G8ZxxZVe/irHg+2lLCVPhnjiGDJIXjMAlkAXZ4/mw94zvIGwDA+MAf5Gkr/GCRNEZUl7
iXlHyRMJt+0VAcHQqcjkGuK2/XTjSCSjy3DPIVqqr86//S0/yI/lFnxOXWcv3glVWWeo9bLpVVEA
m9gGq+DJH4p/gaPnN3LM/E2c+P0yRzak9R7RzEO/GIGRZPZ864N4zNgFWuGKccav3CtumS6DRYU9
QnBDF0FISvUoR3Yn3rWdCpRF0eRegkMqDS7FkwYp6v2X6aisjcf62QL4kNGzQvtXzYypeV9Q4gHT
NpH9acWNG9V3bIgtbejs7MtPUaJ9XPNZu+Kai4DDUM1xIPsSCpSIQAEOpZNAykqY0bqUvckTvCLn
TBPaZtc8Ef+zVqqI9heLEVS3euxihc50/IDCgslVQMy+I1BUvVG/g3ABTxL8UVRtuaTYN2r53mq2
YR3zlkbSqtMEucdzhOzDS3zHoLvMmKa0AZJ26YTiHS9QkJNvqIbqDjp01E0w9/y9GuBIWSbCFUk9
wuMSykbIwMUJCXpaODVISgsuuUXn4L+55x6l1votBFGZcDSRLxY0ZSgi0Knq5edFC93kWzhR8jJg
NLLw0QFVdb0ahd62G7wJwYJptGssgIjPzec+/SqO2xKsoprulMUvEagVTYefwDUh+tPM/dNytBRn
TIdAhQ6XIiGAI7kHQ8WdDUvYDcsohTPrOKBzOBis5V4/6eiPQcm5MkGcJOL5qulkUNnAKHe8KkuP
b1nYvr72QtmwViEH67pBULHM64HBEBSE1gZtz3u0+tIO+hnujNS360u+5cUHR6dzFAby2h+EK/ZY
1TDBiP4DQdJXq9buY29gd3ZolYcdycfyk1ijs2hdkEA95loOaZ2pMdo0H76rL3bWo2sL8TqvSVFy
SGZU8SIzRSDPoCjJv+dOF4NAUgbPd/1fbQUTyWFRQXKuirV2ENFzbHG+OOF0ee5jfdt4tGYno7k/
E+LV+lu43fyfhh1DP+YXg5kQo2sgxklhURGHOT9655CZIsm0B9Lwi1nqhTjyHag1LFwzw7GHzN+W
WOD3mNLTQcbBWJbgqzXIGM6eUvhi/TXU31hL0Ah6BznSASbo5/yWEN3jQJfSQNwPGxRcCYWKGSJM
l2NKpnYDOs8cGLs6LzGXt5feqxpT8XY82pOU4oKRlXrqMYGl3JN5iilnAC/Nfc8IQbgUTM3Z6hWb
egDi1QX+zcmd1GRq5X4CXAZiY2Ib87jUVYYrZ5VqhTFZGQBhj3jUMr8OJ6f7fxtadTjWexhUgF/x
+WjwtGhpJ+wHBkqNLa1F1/no7Nakk+5k94ZAKDh8e4Wk9X+pHZDRoK5eCpaM04sbkvLkqciGP8m2
en0n+GyHoYCEcueVHNbd3Urd8Q15dYWymj9s6y4+0Et45FyuNdcLg7gf4WXefCGsSxRtQbYCpH6F
vLnMu6W6MHRdyEEK9hL0kbAyIci2aPmJJDb1J5RKldUojNqn2h/9RI3s8dGqiRitup4XBNtJjO7F
YtSm1eHJzlkS1JC2ey2B9Dpkjh36zl0jmfbyNsskH9Nqg+gx/ScKHlW5gd0cHTWnn/Q4uqB3YRCZ
oHjrbZPKtiooBB4aaqK9LmoqOot6vSPmRjvmMOjxGkD8DN+1qrfu7rp78w8q7w6fPswuCYVzPUsI
UAJ3zwBM7pcwn2i38jT8rnuSTrVB69lleOb++BX+CPuiswIpkUtviQtYbHf7IZqfH5lpTLIlzyHM
NDyE1UGeYGKRFGkGiS57L+RcwtozqVQ0SBDGRpnNmqnyL+Q5yyHy4R3Y0wh0xteC3DGK0W0/HtcI
FmIf/F8vKpLQp5updsboyFU17l0blp0UaWetsER2Rc4S4fgScNdhLATvwwX72YPASp1KBQZ/J5+B
PWpleRxBuTFIfVZDCWizqL1ygPkJzXEeoYdvIF8D5zFqO1s6cO9382FyaqEbFQJ89Stu8wUVQcvv
SdRDxpzbB63TCWbLTAQhCKnIJ9LHb/x06S1KsPRG/lwgCHVnJkLuqgKveMNOU0SeIJzujt4KVO2l
aHMVSRluZbuWzvWlEK+o08/7Cw5fmAhsKMj7xrzQxyBvNXuFnUkrEJ5XZN7pHkRqSJnrywcTJWV8
PrPIFQBljFR76F0Gc+WUTLGMJ28MhtuIB+h5C1B/00B7GTG+nKoAOInUjuhu2utPdg9EUcbYDBJP
h/ofzIUWJWuJCtUmExpVE+pDQ9HBy0l0/dDh5kP0BaTjkMFuL2Ofn9+B/WNURAIeSligin8uTqSk
ULq/u5NA2PKhsThASLP/pdfOyair+lcPCupct7BpG0dYUi5a+HOJ5Q63t9/WHzk2yRJA9OJIxj4J
zkXqZycvHYz/xhZgjrve/xDn//YsfK4jlj6AsVrTNXuNzI1odYl4KHw0QgcoFMzovapwoAs+LC8Z
7axPjvKjL11UaO63z6Un5Nxd4Qi3+FVzqd1542KpGHSeoDAdwOPKOF5hx/QAHXCm8FbySJQM9nq0
ZUuXqp845axYH77v82McQbCoN5LFfZiqNQylOYRYm2rlgyuxbc9AA6SlYd0AXrHfpR04qQr3QxvW
v8ouabFOpBBzoTRxoMIuZY9frI9hkQwgXzKDEXVOer341Mu4xxf8/28Vb+8ecBrTH0Xhisx3NSLd
M5DjggeLq1020mKsGTNTqDW7A84sxFjWDXmmWmXYtVrVHGC/j56zg4Ku7HKBeSZ4RYwsZw6oxhs6
QG4gZU/ECNMKnfEbcTWIo0Zf9sajRiAIiwrd5ZsYoBn4CRR0akS+8qcvYOKbhqtB1X2Ywj42jOPs
zIIWni6LdujdoG/d0TATB7yABX0WecMoorjE3Ur6nAx17s6oIK0plZzAYYXBH6UYHTzKSriPrOpv
j6guVRNfbxPHn181mRId5pV7X+QzSrD4v1h15vlC03rFcuGD8aVVO6+ZkaCp18VDV1TMt5kt9gd3
FGvrJ6np95a4FlNNcyKV58l5g6GKKceXrBfhjRgCHusDWv6CiCoiBnTxGMghtDdvv2bWasS2ZWCT
fnrNxjfRFN1Wzv53xfJRf+Hg7jJ2n+gqEMZ68VoVZ00AfCeD1ndUeEhBi875QbAyTN4jOW6W7PoH
yKiuuAjcVpo7g9OEJbdbCqhty95/KW6/aUA7aCK1mf5DGI4kjqMr/HWMW60t8E+y+SKcjuIUpOt/
s6G7ey28+oUvpPB6CvP5MYxo0FJW7085iDwnkgaQjDElqAIrXKwZ5SknMnPTFOFVykcMb1WWviBP
Fs0NHZn/j3C5reWioBjF7x23w4DVHeR7NNIAJO3Av5STShZP4c6PjEEBSrAJSZhNbYeBW83l53up
KYcYthv6XGI6IobRLH7wZ0Kv3LOce4QApEge5fPNZVNCm1ULWyb9XdDdD4Fhq+bv6nzdeW5GY2iB
R9UgktKcsP5SO5MMhwt5oS97CnTA6aU+mM715BN3WLNVltK0FUX+bO/O90oGyDVFi+hYZqm7Fj5O
4xLcmLQEoG7KM5FQEUYEgcpaBqv8FrhLmjvX3RMBFefKxQLHCOBah63TQ5ppn8s+vc3a7EDjPisw
gAPcaVv2OelWP756Tyok224fqXxpVMyq1Rv3axB0nB4I46oPT5m35kh5ZMDhrLyHJVhKdRiHuB9Q
u0dHXJmHiaPA5N/Y+W5ZC3m8cZojhnr+fcI/obv9VdRjSkv/R3OtUvP6pQqlTqSEQ+ncaiGs84su
vEICPwXsbvDX0F4rTSpkU609VsKuPRMc5ZlqQ6GG4pPfDIaekmQJRVeCv7Ak29AmAsilJ6JLwvEA
TyDGP6lNh99ltT7sbjbW1onN6i8fFhB3g6U1+19c2xi4HylUBAxZwS/eIXVJUniXpnH26IwkqtWH
cRa6GNytKJQqYYf3IsKAHochpGJRy/i5N2J3VLF7ser7/hrLbGhvJDIWPPaxt164UGYP8q91/1Kg
ed19icsC1GkQUUhubQEaCTaYkHW9lA3jF8u28TMkEQBFYAJyE4qREDRyBLFakXz5UGHH5UJ8/EDR
PenCTHQ6Vt2E3Ewxu43R6ScWVDrSR0aSTO4xjEdp1cAtoC9NEtFC1nDrXFha4bSFupwTgN6UwTGV
5biRV4v07uAyA7joxv5yuwb2WVX+XxS53qpSqaC0ACeBmUezzXNI7BZBv0tzMPLO+VxCcSJs7DW0
XlOofPgIovrNq40pwgVbJH0iK0Cm0QiR91/yWLEKMza96aAAJH3LL/chVSnvPn7ktFQqQcoX+A/J
GA/fCfHxiIMR8QlmtPO6jXyftDBv7iIYs10S9T4wibhjTkyPT+W7sR3HK06yKg1WMEsrkpKG2/9S
Lrx2Dt/OzhyUv3HBoLPg+RCXUAuBTix+MNQm5lfy6j2Qkjv83Zlr4OuxBIr6v52+sDJGvegeEmet
cFq6MJXFc3KXykX6RvSSmY2r4FRiECFamjkxz553IBitrwqF9OSxetWWqIYTdpVHFx6FE2rOnhRn
LWZIV3YClIptiMTdacdXngRAoFtJz5ht+OAh0xibWorc3sDadqsZDFhscA8fO6wa3SB9ZivWD7P2
sRXnRTf77FDFaaPSpkkPJg2GToPlA2GJlG8KdnYETi34ZUIwGTBLE42O7LD+KjYcgJI6Hte2PFxm
2GdCdMPd3lHdFMW7nwKJe2iCP1UQ2PaXpAbQUsBpzJkRr9EZt7WbWanH/FYc884msuEAiPFQHtp9
/iOsHhw+ijHiDeSh3dGtQA6whhBwHUAdonXnRFvblfGgC2atXoPJ/8VnD1hgm2UD3paBLV1/xuIO
Gk/WuWsplu86xDr4uivZoGs+0m4gIQo9b4VhlQbdBLTo83mSt0M1LP0q0+1L5OZFcTToLyAqX893
kyuvy1m4qy15MStaD1Xbao+vS28RaVFOUbjWtZAh0Woijx75ivnUBytlrjM4UxkAU4KV7g8Y3gCD
L6oFVX7oDYUNwIBurQRZ2gFd+mnmeQdVsJvdH8aHWmtegPfUDokqCx5gWB0ulW9kyUsA0WlVgIhn
C2OoZOU7k4TqsUm1FkDAex5CUVb1oJDUuS5uwgYGkotuyZI8axzw9bnwS/BWho0GNMRwJMdbfCed
EVZrAz0PDgkTf3HcH23DefdzKrltB04oyufF1fZKEIOTFmcCCfTENIKmS+hfVO8X5yqOLlW/WdpU
oZGXVACL7ElNH9y4ytByKnXLnghV1ph0kZg4GmuRhzIS17JPRV/dKXsZvSkZ3Km5I3CEp7v4ZyuB
5sMvStS9m76j8JYTB2balxypmsgXmcS/jFJkC/wbr4VvW1oePvCtVm8Zgh6u2oZp/DoVJdGz0QXt
k0/eWlE2VZObYkSEVhp4dQ1UCeFFXwnAeLwZXOrZmO24kCISckt4j01IxYBO4yi5hMK3MXsnb9ea
vdMNdTaneMunC+RRp1FPd3dPnQ4AkH/83yPs3E4JKnEwHy/h2B0kynncoS8SFjQa5dUSZXzDu6gh
DML+6w+T5nonu8xUuaO5k0pAzxJjF6FI6ls7e2XYJbOiWHRTMfvfL7xtYj63PGP7l5XyKWo+QuaO
BzvDTIgtgR5Em192sv/O2xADS24viTnJpXNt+AUMmNcX1QNYOVmwa0j+H+DPlNHv7UtTh2m3yIfJ
606VC2kA6CIslMZ4hpc9C+0TFqa2HZS9SxUOn3VzJRwtERzzYjZdWudaH/bo+RkPdOGZJAtB3CQX
Wy7/EqnkgMpJuymeJTCgskiTUO1PDtBjBlgTOieM0kX2fCY5srzUTVAYXESzOvCLYYAXq5IFViZx
8MZwno1PTsfnJL3QD9JT1WFOtV7O0+tm044tRrfyahbKmd5t3zCrqwLdqgNmTrXof45I6nWqaujm
X0WD0YAzgsOV70FbI6bJeVihRbowfcvkE3esvw4eI9u2de0G/kEixCvDwFjJr3qUq7vYEUSCrrID
ar612tmWrg0uxhSEV5+ypaMjMsAAG4kcbXj5n1FJ0/2Ck+efByQKKrFPeOMsHLWu81cT3AoNbjoW
e1zjOiTENL2EN7h9Z9gIX+fgTQ6duWBbaNqpC6NZDorXu2Wa4zcm29Xak14qCmB2bHMcVWTjZo8X
Z9bCvG2VmKPipBF59+yBxseSkuCySZJv/JU+JiJSs+kkqKfpcRKQD/zzrNyGneovLr7Slcdz3Rmr
7Us0nHGCV0d0ck2T+5GL/MB5LkKPPsXn/lsI6/odLr9ILf8ALEspjNgJ56eOjNobzrzbih0PrKK8
56/RhQLuSDqoccCe/HqzDZv14Z+IYEQig26GnWsgDNR+twH+GC5TXfdhWjs4ri21rFGt/ofoHUav
6oqOOtK+wKEmaBzdlawA4cn2kzNi8ghJvCOSf67YM570T8BfxvK2jHyi9C97X/l5Z75K2o2JGVeq
n8MiWJXuH4JHRth2NytXizatZ9RrP+c7ip3mAhBqHLOA40/F/0hcwhrTA29B8qHwFULHkmW6ZHZ8
hl4BAyS4KaAGSj23Tp0i2M1cguc5skaI7kqUGI4gLT46ZPFgs4Cj8jmKJNEEcf9W8lmjaVCSHgvm
sVFX3tWXzSbj2Y9ZY/9j+pgHTzv00Qhe9OeWOkZoMiUi7DZOYv+1jOFpLac3tgspLNtd81BIAknp
Qf0m3fKZAQXnAyXQkAad9yaQks8vvpim208Q+Kr8Cju1HVHe0YIojU5DPLw1tCAesvCBcNDcnSMq
U4gRZq8vt2Fxppjr1yG4rldtT95KXWCBqgKD2rnhslQ6zwAt4V815T0lBSWNHTQMN0Uwo+j73ybh
FdzbwPMCvRr5Ptygoywa6KTlPcjHx6aj+mMNe4wUQc/0k6voo1lMBOhn+gg05NswYCREngUWuwUl
LakFpyXnrLmSFebaxtDY2PDWRV8wnFwSISr2wh2L1GeFH+9vNtZ4r6B5c+e3FyrvzNZSi+r4GKzW
XrAnOpZj6n54uzfGsoMmme0j4Mw+vgd1ZRXZhEbJGGonG5wvytCuWHONrHhaCGA/nd68H96sBh9H
RMo5Z9KpZllLWKpx3NhMkWQ8lkuP62lRagwIsTNasJhFmTX7SNuUe2/2h65fzc3vy5JueC4LFYMF
dgfNz2x9DK9GaVxWQh5f2MgcBoTr5AlRaXpemQXwYWLOtBJ6EsZbGC7Yq30BoA5M/r+OawBrUql4
w5d5Cb5nu+5mWgfyFpzOFdf6IkAtqral1eA2W9Ygepp5RYE48xTLsvERBjrEVQulFvXC1LqQnguN
6pUfMRtPwJ+EXMFfFZls9WhDdxLHwW+pWyDvkzMU7eNlWWxQHwqhcCNFjR5YUJu32KCgSLmr2r7+
HtBytKBfznolrCPeULBkFQx4kSR7LXAThupkg0Um1obtUOTBpfuv69N13zTmyR9X/im3weGHHYB8
EX6bvWqcVaLltTtKVyzaM1LM4KiXx3Fu17s05SJj4Z0lyPNITYGFz3uPmsizDMSxna3CIcXesAhn
NFpn07WcJ0gq6fnTF6/gRG5C07d6LaMxHfTs7SMvgFTK2TodEQZWqrINZIZEsYRBvSaXs+TgHZWW
5VHXSwo7Zd2mZAQWIUcwAvzXAOgLGUcoFHiX1IXrzwc191RltiTuU72KpXX5z89vyYfICW83kH71
UWhknzxrgl0mWS4cz/3OYu6PulbHE6XxkvXOyhQG2mHT3mndGWQAY5Fb8MmbmMezXtby98mR0yFj
yOK1ylmwTpGa+4gBHTdpyCiAGk4gjKQbznbDF8dNButwEfKcftN+5oL3QKQBGXPNxebh/KsszzG+
YAyWsOLYSZy8mKH9/Ow6abrm3morqNOb1w4uRqEAMJdS4AUnnXbBuzqY6pmrvCHEfn4P//i+vwFF
30IiNfSRhKG54s3KTQmKK1tRHFyObK5JQaj/giFlupGHQt8jyVZe/HxAcWj3rGfEFPoeKEJwtmUy
fm4stX5pDaQLrmJh67oXWBEAsjSrHWWGB8lbXe/ns7trwoWb2/Hv0sdbEfXRTBKRPGIxquYwNVb3
Rtf7YDpGQ5B/k/I7ofCQftzv83j4yK+Svo1mPd4rO6LC60dejnZUVvmbWou7/E/0Brvd3jsO/zlr
CruphpuKN0/pyEREoKVNqeG3KZNIQ6gAS00hn23Hg4xHaO4N2VcEWbBZKcm9HbRInq9WZXmaTY/Z
qQs9Zrk8ungMuDI1j3l+9fU5r2HJgdfpieyhnuhrhOvZxKjQqZOFzIlJP73jwJhxRtAk5Xeu0pXg
2Oyvx4VbA2rTwZwCCwpMS6CK8RS99ydlsCFT2U44QhtGovX9CknJsyqrV/WYsAVFMEm0oWlSuFWL
bkBOxgMVXiSkZ6uNOJSpIa+bzx4FcPUM+dHFThmnoZPNuS3FpjrBEC8O9UwE8u4gYOKv5rl5XKH9
5+WlQ0R9jbbyFDjr3znTdLbohPxZXL4pZtuqbTLU93zO/qoZW/NsH6t/8zMV+Vy34KTgkhcVJD1m
NQa6sRFIMTWHkDDsU9U9B6/SrwRpedcqiLT+u5jY0+q2typ/be2deQlwgXTqRuDfBamWvPpo9CiF
vFCd5WUqx25xr23+Y7viT9iHRI3zm4Yk7hxJDlMAjlDheqw5bYDPLbCY8y35Tscdk72vIuS2DKHg
XWF8+ulbo3/xrSuLH8+uk0eL+byorsLrpXEEqiRFj7+66lgBCdK2kM7+lRVa0oBYrUyiZrasc8Ol
lzv/mHIHd3LaD2XotjZbuSKRvJt3yZTxzBx86gWQ3w4YNUWaWTCEQeNESeZiu6lW0iUqMjEr7TB9
iXGcRjPVdrn7H/aQTtAFb2leH5SiBxWLSAd2MAkuhWHkzG7c6F7FPOwhPo2xRrg5h8j+LpwaJw7r
zbCGBG1KvyIAUNAnIO2a+0gKVdcGOAhjhOeacqESEjyRxr3JyoZbKmqTkcgVKVUbSA0iO5w6k5IR
yzopoqmur6nAG3j9oYd0W0zh0XGpXL83+tLUQlDnMGdw2/ztuLRg247XSWT/thXyqU24nPDYyMJW
uAPEvhNysiHBdkCrfI/d7cFXmXH2mqtqVOIGeh6h2sM0cq44puYazUHwFUYYeXF5eNsnU46icI+S
0S3QzALHmfcOau3Xs0okEKwZ973SD9SwRkceq/+5lfpfYfG3Dlu+SkpafFRYApkaNGIdTVbihM3Q
b8Dci1v00ZRQWH2DBMEB2RvtAXwzZkCKJ0aANMXK2Ikl049EyVzk0gXjRYBIfj0BHrW6xE0nyH2l
z+UGnMHrQVqlFlXEZw9JN87h1YZXcYPuDJwkZQBq7+s7t1maLR2Rkqin/DSW+Pxb9flys6rkjGeq
BY0u8ytyxo8sbnQE19z3OXiW3HAK4FtueW40/ldZJoI3JeAWMG+H+80/4LhysSCZqrdwRzGTNg7K
AYLcvj7RtIW9fUPloW9cTaUoI+oaC+iawvgX3zJssmpUW9CA9P+qe6IZ5A6A9kW5Syo0nI2ZXii5
EBxP6A1zeFzuW5wVymxqiZisj+qptlSgxxvrw4ypNMqYLjiUpHiKLlhDydMwldjXEMKosFFXaKpg
+6klsRvlfUTpiPTUGABX1kyxdOu8351E36fSuzIgl9rb4vBSv4l3a9L/DeGRYkv5Ef0aBtTJqP7Y
gWUCwPW+zAHfvP8w8MijEx1eq1oE+CQy4y1WQtylKXUpBzRuM+3C769UPWdx7bmLa/Uv6Yvrf5sR
YAYMeajaTcBZK97Ljdk3V3mCabhpE0HdtvcO/HI7uBEsyjftzmFKTGHOQjoFdBM0SDzRmCOfAroD
cgkcA/fBvjRSh3/5RoZCE+TqjkTssQD+mNXd7IoJReHCvIHNTGEdjHnwK3Jltg7VIr1stGWud9GC
7/WWFOCwhdnjPJOmJQ0YK6SNDqu4H6E1EmJm9mag1jck7jWtoiy4Zi2U1zNlzuvN/2kGLn50Af/l
MP+kbFd2fn+Sw9PgGcReQCBR/7FKzSEYAtHIOPD762gPVgf5hu1KTjqtkaKZzbYVPZDB6wEzV7Kw
QZz9A/Yw+idLeS3SW4MYyP0lkirIDjPbuWPuKLrM5Ml8W5iqDdsjuM+h/zzxHtMvm5RqQgK+fxUf
tdf3DqIY2jpW9iVYVoWYJ8NwNmbFAfLI8xjoHlL0sE1a0cbGjBXEesac3bYUrmq9ZvKLIyNe8niL
3qhXA+v8qGG4WwZNlZmd5FjML6bo4p0rEXO4nujRWWT3FbQxeN4THUGk1orVfDTIUUt0VEqD8yeb
s5IWJAJMTly153j17JL9pjbCrhPpUUTxdQMovQ4/7BCI2TQs7k1JvtvtfVrC83ilMarDPXCxrxE8
cX8YydP5kyONYuOKVBjr9kNRyTpls0+Fhu+koEglL2jVqfZkZFz4Ttgfx2UTZW0TlzQPXNthrevQ
hp/LAvL5awVU5j4h27/MpVqheTUfnwXWA7hGhBhuy2FgQucpI/zmyyyxLxm4zU/YoOqeCZrZHMxh
MIQrYNc2QrhAmXBJcNnyK1YCba+6udLSXI8MMx/qr+9al1BjxlHfAuzn1JiKITej60L7ekdR5g5b
8b4OsFs6apOfZq9v34PBd5/Z64PEw+T2JMeaGwhIm6mBbGR6u8b4fdAO+CibjnS/kehkgwC/9ghq
NCrUxN/4WxlVG5D5YjELpP+MBMSaL64qsWWwna1RiRSksPM5L1XJcjdO5T++9Ewa34K+KTzLkrTF
wQ3ZvFPoOLjigi2/6tGt7iubbIas+RXmulv4h0vizVbIL7Vs/STRy2LFAdzoXbiAvghEgPo/sk/d
knpJcB4k8sZADN2yUQqpEHKnEa79EDz6wzl0D6IVZu/gm3ooD2QXvZ88SoXDLbw3M/Or+XpMfXzg
IneIgeb2Viaa3qqg4HDN2ZklmwL3YHR5gjcXcRyYkj3LaHAZyGwSmP29KWq+PSB85ghauYME9oa1
wpFGTl75Z3eFpaKye5sRxx8jVyT1nzGykaxr+OvPP7temY8oQWNgSdCFjm0gmfCWdWsqnBRGLOfY
/urzSp7RHmr6n9V32ZoQAHbreZleyGzA0ciUe/r/kRsZ15AXIiwysBXlkmzLxfnUuijnZhhPl+ts
fV2w+PpgVY2aHY3l4MrcCB2nbSzlyPI7Tj0zqwnuFpLpwsHQ/EgHmzUbLdIjSU6Js+TG2EcGlS/T
q6UDbfN2f1MQWwULxoQLEy3CXvNVdrewvxxLtsgJZ5SjREuKqqXQrzYc4yhN9RVpNZZdK1GlReDz
OogDsrzvgWgwkQou60t+GV9nIOWEnSasmEiuRNEZtOMg5g0MCqA85fq3/UvWf3034pRzD6+MPkAZ
+79vTkds9sJUYdAex6VabfhcvGJIvd/nk1tH4HnUicT5cU7iCel2mGo/Ss/g3aNajvRRhP0DrfFj
1jpijl5La2UajQDdMnlfEb279s+yglC9EIMjhL5SyAnkVq/hoRvOJVRSCEUkVOvpxsrfPU4p7ilw
MzE3OOg7Njap1OgkSCGJA1ThmlZtkFKXoyNStVyytz7q9NlvsBNcONqtGi0ldb++EAGzmWdTJUqL
UyjBcl6iiLWIiln+NfhG0gSekR9gN25t0u6uykqtUt2olt58afQFgrmGkNF0PoDsSluq1Rs47vyt
VnFVKKmEoWHZLVLSbcHetEhLIDdBJsUO/+2q2xldLkywORE7KiLFpeVp4Hgt3VsSS4dynrOhIfmJ
QwNW4dtV51nx8w5OSRY5tFVtM8ielM/1wLYZPOdA45uyeuWHsDwuWYHFBEyHt1D08QtWCKy48HtB
3IlRPnoCyQ8ZUXj7kzGbkBZ9MekjcnGmllt1n+vwLI938b4LbGso+6ES8SDYHo0QvuhmAdlmqpnW
SxI0iGQrveuM6cCBWPRgDnH/EiwFpy42jUvn3aXnGNJieetjdrCERYvHf2rINzAcGRwoytcYsmF7
MAcCHCH+72r2alFpT1A4VqR7RUMVYu0mfLceYi1aHYScdR4sv0H1CjGLDjVGdFdQ6+LzGU36O/Ol
GqGvOoX6rNYdwXRp3CX2bPIHMLXzDwVi9HklPreSWHY3Ag88G4rN/peUQzwNgrYBufC8+JcpDG6N
IfKcAiS0eMoi+qp1Y68wjmsZcpO/xfmJ9F1AGnss8xCVms6zjAEjPRlaPyGxiuQBNN2RdLYmkjRe
AUQ/DstjSe9ymuBiSHBnlW5cbiwjCLptz+xpwEmwedUhkBlRWg7zmFRLL+OVKQPW0Yusl+0m1l10
/dfT7rhFaD6S5Xo9EjnjnpS8skqnSi82qML6GmtutoM2QIRYO5k6a9J3ehZez0pSrBciX1rBaBra
G185AAuLzeJ4W5u9geCIoERnBIGv+x1cxWlEwweEU95biYc9MOjnkdEVpGc/dpN2bSAT5OmBwxUQ
Lw+KWTFXSIs5G9rFTCpn9fMKXHTjLqWlLBJwPz7WN3a7g7sKPonKYXmWjgHXqAHVNK6v5Gkw+Obu
7uJHyaL7HtwnGkp4rNaQNB41D6Dpevc3V96hvalYMS4sN5ATQChAwP6Z4ef/jTaAXFukNn3E9lf0
EJkU9787tCiCKtuP44yWM5R3aQs9KDEOo/x7tjZ53lPQS/u6mrz2jTelknsKAK74spGOPleSv5YN
YlEB1/5Kp3jkfTrP2ySMq6d3VmoKUqnONMGq34KaSjovR70r3mb7nZniRfeH3D4XZsstfcYAsJhJ
QKdV77A3GQJXEFAqcbBsrEcurwauilVkshaGZ4rHOG6JmVFGUBm+8QPYEKz0ue+Wc30ji7lPEFeN
nXWV9PZ4gKuulw3RhcNSfQY99bRF7Rkp/QZ/ByWrRY1hkFEpNwO1D+Hk+TKRL/QbZlNqwNYbjrqK
413/z4g9WW8PPfbRbhvpGnj2tMJt7NeAmgQRmC0P3TC4Dmzgxbk9Hpe1NvmK0EYFLYgjFUpEwx/G
l804yctxgM83Z5+xcljIxmEl9gLStEyE6PUNPnaHMrhtqHZ8kbspdBbfgeKoQEFESDIoH22kX2pz
XQctctwIC+pNAoTU8JQFI/CxckiGkAbD2JLoxPPr14MKTU7hq0uNWFQauxLBYJb5WJTzrcKjKkKj
T7X43woWijXYZuk0fEzRnSdWncaHRjj6mpAXLyyd8ypcvXxErPmbmoR3XGhFD1n/kt4kjAVhXWUY
oYhtVHvbDjp4ukVCL2xHhenndePrXgygljtr7JGviiSfMn6I8+f28J4vWDnfNci6CIMy4nhFETOE
aiYSixQigHWoWf9l0qmNoPPI34qgGjMIrAD0O1/YIrwxrDDThOvItxj81NEkjqIMIZmWSNKmgNKN
suuxtiS9gR/D8sWpVJ+OyPSo6i+KJhWHsFCEhn1Jn6ryym4htDu3IfyAZC0LxbNJg/cNMbP0MFS4
fLTqT0EPaUB3HD/QPXYpV1empsvz1LH0Tn4zhZEOL7IW7t705C/tJIq7Mafa3a34MvLgVlUuvD6S
RPrvwnAq5HlAZtM6wIT7WtTzIwWSUC1cUkVQ8pMoI0ZY/ybsOAJlzWqKzPgu/2A1cXVZyQf4Ugky
+Z2dEQxaxiwtmXjVTyZtOS8Om/kIfNRsRZR0dflgHKwYGZCbCf47HzSCqc08bVQR2V+Qq3I4kDY8
JECsZ2+SQMKlk9X8gIkMlJQ5Pu+S9CTwLvc0ETqtBzEHNxdBc88kHI8IgdGJU7hrigy4uEavaQwF
llfJsMZRxVFPOGvM5LBFy10cV+0RwP2IP1D5zXw6X4YB4w81mcOdHVfVtGy32luIktJELoE2/rr5
+TvHVbAxusxH2sYlh2Ubg1/GxqexTUzSJQNhwToKNWNVrSrgk16dSqykDHWh0tIDjak+YPkHNjR6
YTdVda/wDNbAzctFYlpU7K/zcb1YdVVma22wK9rCuRgdnjG+HnD66FFk7PyWgaPGGg6U1fwze+YW
4F0DcWZv78Y+EpKmUrkfp3jzRwdMMicYhcVpAxXgvet9w2v5iY8uCgtb7fwfmt8YHvwR3nACflRg
aNIGl/lycGMr0TgkZLtJKd8KPXCauI6aFOIqbvvLVoavConW37Xemm/iw46GsUAdR5h86dkX8eFv
JJ9ZWfxzt7GHa58Esf3hO5wORNJP3bBhyUiLl2Z71Aw/arz2ncKEE4Ii2z3+rNvEf8+6aOfmJO4v
snevqjyf3C8Rv7tyIz/cvgb9H0Z4alEQd15RNk7ScR/xoBNOZnieHF30s1oRTtrMadEwNhSILi9a
r3Uqq7yRS2hziOiQ0874cPrjUk4O4Ufm8uUy8f2WgInJ9cVoPFgCB9AUHx40wsyP//1AAG9WXqdI
ox9YPyHK0DPOg/+CSJyc9P5rDj5ACuKeMaLrbi2yyhfT4YrsvvomN/FgVkWIOEMQfomhTWZ8RXEO
l6z57+N5VF9eQOsOwpdeZd5FOLGztvLGyuiYZZHmBFtpP5/c80JUJeckiFtLTFmXf9CzIgLBh7r9
nq2zszDrchLLSx7qBdGqjdogqlHMiSe32uw43dOoJ3fHVf12NxNlHLKIL7jOh2uCAdPKfa5zdGEM
6uvepEju6wz99WY2XNCRg9yw9czgD//uGeaqL56Jo5ckiar48L7BX0D2NMtY15pldMW3v3sbRmbR
a6fzsnOut+hN8xQHB2cdk/gCCoewc8kl9QyZfjSxTqaXT5+Xxfyf3puchcnFmcGhCIMMhbDtPsHM
DofAxjfe8Y1OIBy9EItz6HezsHDTBqZPqvzylkilni7z4hQixVpUcSoospBUkj8jytclwnk4qxj4
OPgMasP00MvDOoTuNtunjiFe/yfAuTehNEsZ1+gG8usjt5mJRLh4Q4QHnZdNXnM8ki2y7CV9cO9/
8ZFZrkoii7xtcj5pa4UAoUuUGxC7Q030P3M1Ia+gPkOe76e7RWvhJYzKpQHhPsJaRwQxjZytnLkF
E6kjRcmpXjI6cTrb43Op0JHz+7F8Z5MxcoPRS6+XWDWRv8XHwLogoMNXbqP5YJrMhkpcKC5UliTG
9k4li90AelR66hCQkQSOc17HhRWQR1ORjoX3yPEA15y2n1nVdukIqYvKF5OUlDL9KPxsuJgt3Suf
0cGMmasiK6ZB8uOV0FVbjFNsaB4TGRA55JS9mBYDvee1QnvOnOYbz8epuFy4b/w9GUJwNNFK3AMQ
U14CKCP8yFRbPOnwI+YIvR0VcvV5X2R6Qim0xvUS4374FtO8uEd2NidHricVA9oaaKv2HDAJ+KMv
HZGQmvn+W2afLd6PUw3bGm+pB1obwoTvn0MCmK6PmEpyWN1kfeMkaszHMg9rIYjPgnLXv6meCxy4
p3MghRip6cr8y2bNeUjcNbBDcSIITtuxNtAAfTYe5tghvlKPn4+sHIA5+mMV1wrAcfQlg5e722qr
pzXuBpeXyvol1TICeqTpE4zWIyimN9jliXPnTuRdYPp+n7fh6GMNDPkdc5DKme0YPEtzYfYkgAXp
I5auudrGSN/iO0GWmtBar7kn9D7NunxvXynMNtWrL426Mu7nc24NGwnJ4LnsZxECj+sdKWrG0dNN
JYRlF1mWY7zYuaa2TWcDYJgvX69XXQtxu9mOb3DCej4NUhrEVr6/BYu9R5/0ijhdnrhOJEP5cmQR
2GJAnadF7jIHkhaHw9SvXTwGvcg95Hbdh6y2y9cddH6nU/Gj63dwBL4Xd2r2jQWGXzPNUzs9YVa7
Sesps8N4hdNqi/s65+1dDRdOXkp/isapBhUOxXLaMC/raYxmnN1BHoEeW9xl1+IZbPlrT31AXLmH
DYA7uF3AJ2++Y8gNeQdNTSum781zspJ5tefAdioDsYeWva85Lnutb77S1ejPAFH48hgU3Nn1gHbR
WkVl/C7VgTmP0tfphBXxCFQfbIFrDbd31oXyo2+LRhYb2BCKg5Abne8U5EDKQRVkVPYtMb55Kfbq
utvvILM7MkdpYfPwvt+74rbgy4g1D6jMh2hhAsP5S2jxxPC+LPBKeKUXDNaKl+MoS/b5Zm/IBbeF
p4+FKqIWGrfvvnTdo+7zoYVvsSxtgWMlxwN5YpXN9ihowZD1zbaZLbOPnMpRlH6zjhx5roOWSewa
Fwrc4UKFrVz4S9FaCbqSubPhnEe2bHdixa0/r4gO+xuYxiSfIvoNX7yALdlbIbb1FGN0OhRLbwF1
3H3YlyjTg9qMDTeAyOJkf/+bl05nKOsVLTvo4RiBRl3aoyC85yW+/S9xZUgOOv61vs540SPSt03L
g8thEtlxROtzoX/y969WB32sXvzqzKG3XX9zsLyYOy6ovCrE+x+BUxA1NEoC6PIgfhF3zZW+0JBR
D3vuhLTu1rS2WXooFZyWNMyfcQJvT9JNi4vhgttNmS0pkocA59Y6xW1m4cV3qhaWTiBf0GrgtH6a
JQUNoX51t/xyAZ+mxkQLXJ0XBftJxxbBzDo9pilmOguobctHDlsqd+75KIP8B++7D1S3NZB+R8tY
XZk23fqyknXuCiaeTX49nIndXO6kqv7Zlwcx3MOujTbX2lJiVKvFDckr4wrYWaqIupV82qdJISt3
Zw8sifcBSGdwBw9omQi4Iq6pkciQLHqyFf2crcq7xbYkI/kTg4iNIBTjMug+Sjfyu4wHlTpkdm8Z
+SPF4Qplkyo4ppsNnB+UdFTDi1c3tJ+djYdVdbSJTr6TIZRaXMgKCy/VuWKFDcGKZ7LsoLfeZUSJ
RhVSAsSxMtBrgsD9POZY4ZtcbC4QDksjJOT/yQudPWH3TZkk1RlLJ3XwdasvpW68ZOR21YVEgJgO
qlHy4Fd3s5GqYQfG9umlRpnQBCQd91jcKipOJ2wRCiHO0/EZSNMPCoIc6USnsl/zgK1SGuBXO0nU
aaWntz8XZff6iLlqoFVUSQ9Mnvz7Nb/8e9VUjj/9pRnbKU3SgW4LO+3RTQjTnigbFi7MMenZ0aZc
N+j+EgEM//7xRVEu+IWfAGmKqU/pVy8yldi9jt3EHM+Y8XK2CpaO6nXb2kEmMexgRHHndv+WG39G
LyN3zxm3/J3V/6i8OPZM/gBVTwbJdDmJSKDr/IAJG4Bnkr92kcH25+p7/VFvcTwGIRQjpFHo15QW
33+g///KgqdXdBjAAXebwsc0imOVqo2rQL9gUyLrXnH657ybdLhqxnINJ7X640edc2jv4qpKb9Ye
D14eZ15UZaadBQTZW09ohWFzhTcjcS9XwZYBV4ZLU6Rpl3Z6Xew0NC/0xNP5rYrfZx/rsdFYTRYo
EEfFZTgMseGfoD0zqpc1ztzFt0AAWZ+C23woxxquMe2HMHHYqgbCAA5g9ky45EnVimHizsss3TSW
a/BMTun1uKTrOrJuQ6LS+/irvqsxbkfkzhunlQifPx4rCvx0fO4HbPaX/yx7mXIxXkXGxzTvUmuD
MHKj7xGe+3xPYPHeQBKHKXJSB3MU2YnjTY/WLzvm/B+FwnKafHzAM6whDcbBs0gvTtYpetSJhg26
InN5QBUeymLvgwEsRTIV/fgA3wbXmsOs100ewRTAFhtf9scl1Y1AQWnGJrtI/lVrQ338sfn0ST5L
AHcYjmtP5hXLxPu28g6wEq2iBlmfVfx7ZAv0hmQ8mGR+LF9MNG5qkPb8LAJ82Hm40qnOGDfI8yhD
g/kc3HpkG8UPKhG5jEgf4YRyXmXgl+0QDqs5z6Ms1japIdLvAOLPZ2vWGEiweFka0AHiHxwdWNuU
V2neDAEfQY/eMSm53NIznTuO1LukjqJzlbP9H5K4nRTAeecHOZUj4YW0gPCGMzzTBroafdHAnbSP
9FFmRlG5+64Vxk354eABTFohpYfLwaVWWVXLcUdAcEFj1HkLvg4OWucjlI8ENNpEHWo6z+fs1qoh
sUCSTycB/lON1jvNFolEN8PXN+8x/aHOn87nVAB0o/OdGBAyKJpJPVbOT0tnHSNClAH9ZkLOWOtU
Smq1+UuWLRYDeqbEuE/Wg53Jj97C6xChRpAoyEX1kz5fiYu8T8kbSLoKnS8EMQboxvYYgQKFwrtx
yju2ZcRUtlsVaPnzplTdrou1F9a+g6qAoqrbZVRFQaIIdR9NHkOWF90CdwseziUsGaAYwcjUMQ5s
5xW/W5n2JPHFl2XC62YD2Zh/qw5XdmjKpiOcoMFZdzrWWl7vaFauzSBaBRldWCb+3sibeJbGEo/S
f8O+N+zlimHohss8T5IWZPx1PSvf6be0defuNhQp9l+yJtBVbdOm9GgFSsGmuTsZ+Itb+OyfGz4U
8uduXEorx58sONe/5Y68N1dzgYcmvm4IBg7f39xMWZbkcb24VTVuPSoUA8kSp6g89TJ9cl1L1vN7
YjLFFdS230iLlHA91KbyBbb63ekfh0yjmEne4acEf0+j931UQbsRJ3sSNYFs0fKAxEdeTRinVx6T
TuVnWVoQerET89pcwQzDFlGoaFvQRvwOQF5WT9AdI0M4iytd+3TqUfaL8UhL+PbTDRui2JjlpCFt
yZLf4xOXD2u4hXjP9Hva26pu95nmiT45/33UF/MVJHmSAW23mHs3jBrsZ2AYtMwoiYhRQax/xugI
SZmp830/gdDDuK9SIvJ/IRf8facZyhuICbbjSsbyB07g8GY45IDBRdtHSMeJa67Y8zZl58h5Hu/L
nLCmHzsFvtXflW4AjHgXH2wi3KmQEyNPGUjc8jsj+P4pIDdrm8aZEe1iO72sY3GY706ayNW737ST
i1ZGkVZzpkMZhVaccq3cEkDv4gCv9YL9dFrs8SUKbINqOmvAXRC3QKyg1JfxOtVgZOWB/pKVxUu8
0KIREDIitDD6V8crjBNg3sofFwCDQHX9EQXWMEEJn00hLyd2vnLr0QEB1qV/nsx1hSOs5CxmezGU
ZM9vwOgVpWjk/57lBjR7/AxHKu3fEZJQCF73CL6DFWNG84CUyogB1akkwZg8WiZ1ggujbUjuFEYk
1Ol4KPdF8GKhG5GEFnMw0zMLD93qWcsFbsmsCdxzzV5q8H6G8y2s4F7CKf4w71XG+kt/AM9T3LGK
DWotUAL9PGB01Oqly+OkHHaMkH3qgH5eGBSmT6aT7C/BWARXcs//evxiTGejhhd9yf2fFnlIm87Y
mUsDB3K15pzthuZiVTSQwKrObRLoenXSmyVCvsun7XLfN8DCBMx0StJZ6uR6DlSG1J0EMOdGZnWX
m2RNr77oM+DduNWsPcDKYmKkOw7vfHDtDuR+PtiY/Us7Ai7bjpAh89HcqmEra5xoUJXxvMTSQe+y
gKMTmeblM6eDh8T/oxzfFtVe1LktNieYFunEUz72SVrdl200AAINgO6EOkHAEIl/O1VBPUIuOrEv
BjdQ5JDIhO5Yz4+bomwKRrqtg+DWLZ9aXWSrqO0HA7SwM4JSo1BN9h0Qk3oXFd6ZnV+7XorXc1uR
Se5wl0W5fUIrhJGv/bhjegOmHyaxcwIVSvtBTeAtbvOMikMoKzKnwLoZynnqLBwy16KlvICFn9eH
bcrMP2p4BRXybsS6vZE8GTWQJHmRzYIlXNtRGLPnfJt36QpC4ex5Qoet9M7MQmJz/aeyIPgFNhdx
4FuRYEZZ9DCJFjQoxj9ONtL460TA+sX5Y6ax/eKtP4Pw0Mqx4wmRsjl65obn8BhFRxZ/zGWheei3
iwHrmGpBCHxZmfelclxmDQMo9E2DiSChoLQe87/6y6cIbUSVu72oGoY6veQ3ghkjw5nZJRo0bpUp
3on/6Je54toBU6Pn33BmFJssRjn51ZiQth8IM3t3ALPPSUSaGLPHMmhuypZm8vTReYoyUmbyokYu
aE3XLIiayy5tuwFuGLf98x1cpRG6XdMJ8H+cBa4TBZ1p7fDQXqL+xNjZHzcxnkVdr98Z2ROedQNJ
5lSRj/N0bzNmt5woPPaQDRIpBAMS162AXeyCAc6IG3oz370UwQB3UrgMmsmBqORfkuuMtfDlRbG+
jVX7dfXA8XJp6kF1v1kuaEf+lcBBY018Hlv0nfuxdECtc51YraKxV7K4/0gQu70qbfRdmc1ZAAUn
8GderR5xc0q1cO5qc800M8SP5A4Gcn9qLZv7F/Og9hs9wczCrNVqZ7AENG6FdNIW/RnyYCQqbhsE
63IhwK/sdkTN015/yThdg08H7PNRI4wlQIorjIEIw133ZNh+9OjSpRfyzGqqqw5heh/aOp3PK0Y1
IroK1t23hfR7SvL893VySB6Qjy/A9I7asJNbFlaQIqRfkM39uHzRcg+PoGhH1U4j+NI4TSdoy2i8
z0kr9AII+60s2z9jusp3FBealNOz1BesKohKPTkrqHfyyZP5daHZhHV5OcNTquOl5JHd08vBdMGr
YLjVOZOgtWGFXJSIl/Mas41Xv/sb0eukbn5S7XmNFruTo6wUDoHiweDGBldIkvbEKaUASiY9ngFy
cLNb5+67VJbgRuxQ+gCZJuaXFtgb2dKchAu9gcGnsN3/kdyTILq1CYhMLurUoRq6YWzTR+oEUI2i
M8XC3bUO//f9ssoAKWHGZMwWMxWxRhAbq5F4T+VisWj3lViPMmpjrYSXs0U0gBHpzzLhSVK0KHM/
d8JaeeL24MRxAL0UeYXN9XnRjdGlQUciGaQYO3zy6MUc4uowkP3ZESJ4Kn4xa7r0tz4lf/1kMITU
Od5SN2tuH9nQSL/E1jN3rY2JvUYPpH4WJsLTG2XKkYL5RK2V4c4CHFEM/PzhgElSqb4Xrp8pkyGK
yLlSLcX6iAROEhbkJPN1X0L1z+FYVoKVJBKZkEgJdjAtm7kvGotde2DlqBsLsab5kHdzxuD+Mg27
CSxhyrEM6hmuCqwqCbwLQ4ZJiQAw5LquB0DwSuf+x97QdrTG8kDLjWhxM7GLV66vDKrwtuJ9M5wR
X5LiJhMRoiOOXh9Xzfust2ch8tCtZEcDMVwtr6vh8mJT+4Et4oEQCqUS8A0hfoSU87Sl1RB4MngO
eOIWtgzl+Z4OSh+7mWydZzF2yyFMzFlkKQeO+Ag1+pbnpF1jXk7MTgyxjlSc3kl8xpEPG/K+cyGX
iIwv9g5fjcYCR7amL/EmIgMHU13jmQFam3iINyMbpeoK2h3RbRfj0eL6zFlkd8BT1UKRx5iaEoRb
/+yJ3O02J1edLj9cCj1/QX8rDXJCHGU0G0S3rdBUWvpuaCJy5HpcuFiIL+3iGFEamGQa8G0+xDu0
h6p5LeiycR1/TQkcgt4z2+xL33HRiey3IHkg/WVfzmZCPPq4nL6yz1+Sh+ViMW4knCjUer9MxMm/
2BUNo5pLYzlythcVUFHyo6WDv4PcFG7FnjBmae2bQkgtn7V1MbXlfXZob+dPPwGRgKDTv3ZvcTDI
Ec1PX1SowEoVuXvXQwbUqjRe35acPtkSTHuH5qnNBKAvF67mYXnYopLd4o9Vi+A4mIjCUcTWS+k+
hGVZRXprRS/HU2bUs60ToGegxf9seE9yVCNiw5j3EdZPh1mUkQ1NizqloXPq3rZ5bLK3NePfcres
cK0aHwLb2450Tjc1LCgzUvTZuliciDdK54foLHTXoWHm47781CsMSN875WT9c0Qea3bNseUnAXTV
tpFfxLjdK/3PjPHCo4LaNPJwWDQP28kRzcwrLVFaQ/wYYHbzdQsxnr4Ex4mBQjyazGmDCAeypwZe
tw2gE2Qjkd0Y5JHIhn5McRNSuIH9c1A8yXtOVWbGrnQYkLkS1bcsR5GE+HCoBqaUOnVXe77reSqg
xahgYr391aEPS27JxpG3o3rBRBCnIXUW6GqrpRggkJXeJ2IDxxrDnBQ5euZKsHdlZLZlR8MZ6g51
FNFj1t4lhB86kiIKqsyH6pg6LkorNvk7jU6uuV9dBXh5XvKeVAmsxvpi7TzdFxJn75qQAmi3JyqM
W58b85DtTYiJvcSx1OiQuNS9i0BCfAhorCaexRUbPo5/5IQl2R1UpgqZ1n8qi07YjmrU52/4S4em
GZ0Ehy0Rahe4lpTpjjDRY1k1OeQpDX6O/+wnvBJx68fQobDPkTfAPEf2Po45ibqkJwraVDZN5oh1
+30eah+6A+HkzaeDRJsIZj02T4Gbzh2u7kOJ8Y9JxYEQzxiYtl3SRGXjaYn6ZTyf33lzuxT4omXo
c2bG8ON6gls+OY1apxSGFsj/iatVad4R9QoHsfaOH2hs1tQcf0vUu4JTEaC/JqZgrX/3eON072b0
Y+DV0noLUZYh4zitkQjyy1rap/jrGh99r9Rx7pudMAK9Z6+aPlWX2veGFCksyauF7jmGH5g79OTN
YLt/zFcEpOL/6BqGXho0ifrOv7w1g6I2R29oEE9OimaQe8WmEr0fqkMQwrp80ctVumhn6dNJD39q
TQyP3HLlWUXynjyJVx1OS1sqfJic+kCFsOBXeVcPdZONC/IK1+P2NJOH6vyEQPaqkD2luP21ucFp
VPnFTr1kZwZxF7xhGj2g+vIY3t9qg1NXxqh80Emeq49LQu+T3ZSozTwq44I2CWpxYBmKUOXPElzZ
Y+T7Ehc4zeSC64JQMJi1WZQ7iW8hz4tg347VFvc+BQLzgWqzUmIXgn6FQJKOpYk/d56ad0KArq6+
cR0vLcYRR4yTDOpJwEjR3dj3z3Ey3Wh3aOaw5QBc/cKHDqOUhJ2oTdAjU5BQfPFuXer9DMBC67Ad
J7E0oj4rqOziWy/HCtL04c5dMerP0sVhuzyHLD83GMs2j2hMm4CDrroMXtcWwn/hN64e2hJJl+1s
lq+KNHdhOizrwfCkfCkkSwovIgCHJhMJqv6LFftG5a6PL4OHhuoyD+bbP5Nj8/Oci6XYoWcOCt9Q
00vEyTgunDryEAMYbDGKQT+eGtlM892TLahPMS0XYPJ74xVoQo4PTuF2SQHB487IO6n3nYBF6wAU
wb9ugxuoPhef8kSpVkOXBR56aQlsXr09NtMoeZWtn4XFfrf/5AjjrpCLnlkMb86UOJc7Qp+WKhuu
lzu75xXs+MQI2v9pMmL8n5HC2g7xNNqfx3WsacLq8a1wqv+Vrg6X+atEPjBY13GAbVSCY7Yt2XlQ
/p44ZqvDoWvjDKPBQboVdnhhc7BfkRtf60pzdlh1IWB/GPeqsDhgDMj9aTLqr03R3HxRika0JZYi
YlypHXdhXiphJjEefHsEmo3X10+lao3Laf8Rx0fl3LFJ8Cva4/b/Cqtp1IDWTDNoJdfdCPBftuKZ
z4A1cjqTSWiqxzC3fGkx28qlUgfUXz68pjLJdhTISGSWw62tFKtfIVuZvtqB5ChMn3FYboExOxqB
/XRvTFDovRKgrx68nR6VuScO3vbBpAuSpiHOlnFRu0z0EhJ9Ida4ApgTWMHrqEgWSlEO9b5pbcGR
rVB6bD/UVwIrb4kZ3bwPMV/o3OlzTanEa+moruOGU4W9kxOoTJaHxr5Zou0D4vdaUFjvN+ICWbkp
P8RuSYItKHqrhU184iBiu/G+ortSVufNM+/q+bZ1lUnOvkH0fNl6L8nlRH9Uf3fLwOKKPF+BKo7K
UTHlSnZhwH4hWn8TjJPr1XYrX7WJ3gDH4Tv0XxBY5hOuwE8x1ybHlJZFdyYXvNjFHbhzBbB1Ny1f
KgauQ/Wz2aorDwERwALInEy5KaB+Tml7j9t6ECJHCgmoY+xCGCoKoYIVo4LcXnSWLVpYwuRHFu8f
yYGI+S7n5xRwpPPofdOMfVfTdAQ0vs89BsnbI9/iuHJCNcz/m3eKFz5eRl2+Hg9mQcx1CYAKZLVi
/RmyTKR8jkx8k3/7nrGOEbC384620u5UlMxtlslJX/cnT0rY5PCBRBICrAMRRcfM1geVT3zg4ElT
l993bGwg2CYnwb/017B7s9tgmH/kzaaRyfnq9bhd77OZfxXBUPOAwtKCeU/MCzM8o+tg0Yy4zrnR
OXfpowRw7tbFMSOtK36ImjloiCwt1/ZaTnyBm9JQW5MrHdXLFolDao3bRvQAumnC4GJ0d88542fJ
tK/P1h838+Qx1Mf4Kkjjy5zBWDztO65Bu5zX+XFZaH1OZKNahKCaeZ5OJr7bQLDKbwPk0hI//aB3
kHcx14qqXBlLH5ppoav3T/HLnbVJ/SvIg0f2i3rxR5yGIaATBKOXxOaWVspmOXaXiXStLYUknSbY
s4C3D7n4E+cRtb0Ssob18YLHVIzfCNjJLGkkaaav/qun5tTXUQCm1mPhqLQEOdRuEFPjNfeUL6Xb
WbBnWx00Po8Td+9zL2Ae9xrqyZQlFoVSLU+gu3Sg3bn6V0byCLPcwxdnBaajYBEAEC9KBXqz79uI
UPbPZrlgnkeu9hS4nhkCd5WL9zp7hrgOmBdS+9vHnbYzUg4Bb260/41tz1MNuXsRX8scy2ili0t7
f4o4E7VZFL13yP/ONRrqfl+03GU2zUFHZtqcmexgtbZ/V5FAr+ebu6JwmFpeJvFIixIhwN59hYTf
tEkMFwZsexk2g3JWRwuAU7ab/35rMVoDs+pQp7bHheXy9wtcidqr+bbF+z5hPcRuwH3hCnCHfMwU
3VBqLm2LqXZNqRrk+3IV7ih8kfXnwz1BHJx/zm3OQ2tYhT1yXAlnDGCnL1OHQ2HYjoTjCBTtF3VY
e3O3b+/96X2kQyE6VUe0+56ravFBGUsMmZ7ARcLa6544kgMEhhlxLvuwP3o7GskhG701Rg/cxNnA
gAakl3y3T4OFixL26SBU+7ZCpWaWhmQSyamXnPUTfXwdz0pOX/fM49Dh37h7wV2jltspIgGAFafT
SuXreP4u2W0M7mno59NFhf3a004+IZBmZIp0oTNPr8evZ74A9p61aEzoe1jCtctI5erCYYKKWDIQ
2s4gPt6JCZchrldCFldcFZ23CuxrJ6MLoF9up/bMuH3myQvDe+G9pa+/VmdXg72tO765rsZIm3ra
Ug9J4ii13o1AAGPSjAceCHa+1fQXdoTZv7Yi0wNPvCIbYRXfQfL6wnjZwmnh6DSwzqRenK4E+X1g
8KwhHV1l5hMe8CSgAZrsby5BY/P0QLrzlXKt6mTWWRHFHIWMRaRSvv2ZjrMkIxltU2zD1KVqKLHC
ONniKbWmmDeP8YI77GHhkax7wfg71Wvok19tK8GMFcixcPXnflWxgySni0BiMId7XRP77LqyJI6g
9Zfs6ZpnMyWQxxAKMnjpfnZNxlj1VPufg8UAI9V6s//LcNkabHc16Ku5DnNw4Dfm2b/xhOg+HS55
kGvydFxELDIa8cVrOjOpxwTjZMCPsR79eXlVSnP6Wr8v1LAP5aeGv8px0VVa9otKcytHj/4a3Sf0
vqf+yFtpTcmi8qwDzqLAA2d4F21UxeZutwx0t8Vbkbea+Lq6hvDu9HKxJApSzf+4LrabHZHmw3i2
rDOjwimQ0+lS+OYg7qu8RzM/BZ7E1uJyADsmkxgOiK3z217P3udZugX7WohvnOsvjv7a0Gf8JqB3
1xTQOk5DQAft0ISdPJkE9Roq+YNPjpFRN/YIsNcjELr5dtEVk4epizeUAnO0tVg5P3bvhjgVjAEE
3Jng8pQgjoGEzVRZyYvvGZjXj4U6BVjT0gemI4MHQWSq1uxZBaTdK8aw7C3xWaXWTEGAabQVUxdE
1Jw31V+vjGF6XcrYuPQn+BK5O7kGdbWC198/JDqVolPEr7v55VmhojfEJfqNdsAiTqjPDi1x46F7
yjPNbp5r+4XMw8PghgU+vllzWlhcaP3sXdCbN4/M9nRW7SdWFrHEB08YILA+CeyYszS8pas1wbrS
WtS32AVBRh+DsD+vLLikz+Cyc0+bHl3MXbN0uBkalDc9aPpUvo7VkKlNdul2VSZTwc/zNWqEHNZX
0vO3Qv9KZkatPJb0GxKqxT8At6H69DD6uRRgt9iNIx8PCFiujndIyx8kITwAvEOc3DbPLl0PXX1n
qxvtqip+qAwDUrCGkmHhYqwTz+8JdGI/+QmWt6mWi5U/j8NilyQ6AFm9T0VcmfCXtlOz1tSi/Udv
jrsiQqEV/TB2R0sf7RcEsf/u47VA1iFNqD3KDn9Z7tE3LFIsTGmWlf2UwgkEH4UIyWXrHrdDoxM6
s1ZDO3jWR3njyiMKyjF6PSVDkDZojeXlGEhif7skpsOMDboDXWNAQCVKo6OQZ9k7niZj8cTEfW/Z
g9Z+OZtJcnep8Tpc3S+2dquOt7y/0POvzRw1X/0qAekKyDmVX/Uz/IpJ4cXflVd8nduOg12NpnEc
qSNItW1IgzWLwHRbjap5fU5PoBNoDjELWETuLV1wpNy9qShBSifzCYJiESDl5ofNT3S4v6g+ktOn
+K+O8SE9gysRNvmfr2AfrCbeAJSdzsnZHqTtf004SPP2rekoLBHjL0jSeFxDpX18w8l18Vcr2hlB
CwbuFt4htm4jVhiYr5NwYrXfciYVzghg4+QWpKX03K8vVbpmtgStRihnxHv+dVk+UQtH26JLrild
6GpVuUBdvr1Ev9Ir6fT41OVmVmBczgVVnNjqrd4RgdayOjdGV09Yy6xdMhZvx4Bb+AwojaSQXole
FzXiY57Hk8jbIibXWUWUq4krCnAkA8fpikwunGP7PC10nGiy+b4ql6hKroZQSx7IkDbTdwfh97Hr
se51IMjX4F7tDlDrbtGSehEyKFHE9AYsi9Hj+6PcysvRHuSI9ON/PH3BeyDhItbvkP09gvldoLBV
hHUUiT/tsieAbxa2RTpDapGh5P7VwxykVp/a08MYGvvnhVR3l7GGVKv8rpU1nf1QUjmZUV5F7xdZ
WOQ07GdSZ26DjSVWaaJXUc8N2yHC281K+ASW3MDJt4zhSWXu8qp2OlGGAy/cHdBZP4Ye9ZEUdKek
1eoc0WRLb/VPu4tVGnbrnVfz3bWZhj3KMtr5RiZG7QaKT0VOsIKgvS9HQ6O0z0VONYiCJ+vQgcaT
MGKDIer/nbjMZE8IJ2vjs8HJ9a7pGV8rg+nPm5QxMV6TxAo1VlyA/eSvYFwrxv3JZzDaqqtw7DpB
Gz6UgPuttfe7nHEsQee0t9nf5lxFRwrBva83U0qAXY6DI1HOODOcgVR6d+FwAPP/OT83wlXopZzR
vbo4ZumJ5W4SDG77rUdxqhhI4xdd5gqshFE7pQxVgG1ZPg4t8qUiaUKQWRwFA0OsvIXI/XucSsjR
UThCFEjrIiHJiElBKXdk99+9p/19IG5MhEwSTjTOZ1itq/+VCc4CGCpDxu3XFbOjgDTtgZcBtWBF
xOUZEXPYgXeCkF6NKzVNp9KlgnPt4HrlbCLP4WG5YghwDqVNsA95i1aKABaQ1o0MLP0szuk7UoZC
LvlB72xSwA9NcHeEMPJ0PwlPicKQvYhszHuhTcRibpxXSMU0fvFCdKz/qMxA3tWBbYmjnyeI2zhE
09z0emHmt/ZcfnxzeDwqhTMg80hbc2pkT3D+IlxX3cmjoiEsCojP/a1pkG87C+n5m0ZaevIOSqQm
wPspMv+LvRAAg0RmY0OR+DgBN4eM4DAlTk7FfItssK0AX+bcp4v9qJujhhcwQZJmrObQEToBKSqq
PynCG5E8wn8SFsny0gVHusK71XRPMscNO4h1SZSYyH5vUYiUQIuewR99BcywobsT+wbyHGl2wLba
hkwhOZroKzn+gC7P7NOmArih6c2gusoVU22d6N3PbFdrowAEuF5FfQPQs2ikj/BLdOnUjkbKs1eP
O/eqjNEKdpowrgd1HVs+GN3iSSlUNdwHsFrpkWNbzOmps8hmAs+XKBz6Zf7mRVsX9sRuAdd6jLgM
XRrH8wTE05VsoqhdUGEsxm4qvIzv+opP2lCg/K9Pul0y27Ll/Q65nGZNxYMZpvpugLctdSoyoP00
hJQcRcScZkxrGQ5Apuw0apAUQT3kJratxBsGqxX/Gi8V6UgC3rgGCszsJXUC4E871NXaMYyHOjdV
VCrTfyPcHjWU4QPYIQQOwwBJzacLek7ayLuR+jVAtVguSdR9MNK8mRkAMQM8x9iSPohVQRaw8MNm
Uqqtxi0Aub7os6jLx9d1cQOyCzwyFG9XaK5WC5Rguug4e5Dgmd8q3LIL33s5vJaIElRhu4xFJ9OH
ZxupafpPoibccnlIH3rZ7sNVP45R/zwR6TUI2RKNdjamCoN1Yspk+efrf0d5ELu+zdbB4LF3+OY0
JymfHTI6iqui/KTxAWSSUpGmDkjji4tvvYUanI2ZwBp58/soqTi6X09QYo+MWkG1H01d9rW5+zug
LG1RNbndvQmiifWVhzXE9DvyphPdvRz5uCtlpQDibV+TABN08In9a/nB+PmZLAM0rTqKs5DNQt0e
mrezI+UmgdZAvOPZDlgc8mnFmpvumU8GbjBjRWMHmGRytBs90eOhSPSfmj7yrF4vUOUmEHOVtqSi
LpwiaeHa+feBSyxOmdVpwGReNyRV1oMDmwJ5c95LYZuc72bkFCmXU4pOXuL6jiuIoNdpjf/eFWaG
GbsgoQ7l+rLH6DB/URI0elhBmPcSI7C7wA84kd6hPcMHb8gJlGo2REzazcyQB/kNXXuV/c/jUC+d
k7IJLPzFoZc3OJNo3bRv1Tx1qudFt/Lzc/YgEIkAx59Vxuja0h/7Ncj6xfWnCyKtAoUhabXvisou
Til0rlA0RWAICJn+fV2u0uDHaY0n6VYChnq3Sni1iSRyGGCBSlfnxqd233TOt+mZie9h2hhpxGKD
7v18GwnrB1FANrgBe+tqbDMPybKR3YWACrA6Fi6Cq9wKlfUGyg9UMl0wW2RaJyvBIHuMX42U8LBS
ANy9SWQxg1dj+a5CCB0sjGItpsXkJ5Z4h5lDB+IdWG/Yb4tE+szpIRQwuxsfBzoaQ7DyBM0+uHSx
Vgx4fCoIAFBGg/kmWrv5r284e5aM0743kfTtgPqDMiJv0kh0UyyqEj8q9DN0SCcn5aa4BU9tEkew
7xTniDNEjKnsFDwpY7DH/aNPkmRNTmNCSiA9nNeDJsta8Zpzfy+OWKVgMDDNoYkPO3fUIu58ugLk
82z9BPky+YIts8wGm7pAZC9P2oQ8nZeABX2fQGriTjmXbD6kph23sLDIoW2d9cHoDoMCPcX9soHH
nO0zRbNCWUXNgwOQTnfD53sFm2MdFsC/dvYz7cGMBCMMl9fIqMu2VAI/JGJE8G9NbKyxHhVVtItK
zQOekUgkcptbkYeeAr91XwCsPAg7aGwlP60F2g+1/1byidpvgcADnNHYHb1HIlOaAz2BGU2XOmR2
qldbp7naukxlx8QJeApkJqnYYXLf0+gC43St5uim3kL+z+/bTHOIhL5dvMyQhjelwH4g+gnOSMcw
geN982ChCHOELeXtrVP/cKp4Ok3D43OybdMucSdTEuUvA1wyzhirdgwj0b/oQdgd+U59s3+irbuI
MCTLEeiPs14U5bBeWfMSJPKkDxaDL4SvmlMkjqQq6xBJprlVZt130sjfJ1L6wdi8KY21OicxVRoP
QptKLiuqLs9/qIZzjTu8I6sGdt/HJJxk1SAa4IunEezEcRso/VvENoOKN9rL37D6SRoFOx/MR3yJ
ySNVdt6Q8BpCtb69r4WvKWDwnfMmcPh4xd7bKT3oLtvyQneE9md6i6lJsxfJdxT73yOydIffixU/
Gj631amAndE+D5gN2e/OACi60k70/Pkz6zqgpixQg3fXBuwm+XK0FilhkynwZzvz+STkidn/Z4N2
E4E1tUWeJRkG6y45habiRAEB0YecATScyamoEin9KYRDj2mINCaI9jbMmxUcn6m0pzEHrnQtMFBy
/QMWSNqX9nAHdMLslMgBOh6Q1S83IaBumns//tYY5xWUaDwHFhFs3Pd7E3+TYKnCtelFjJGMjUjU
vYUXUFtekXIhn/T3q/yetOpD9H8nrAhA0jxk1pGd0EiI6ZNrWRvSkACNbEfuCRNbBZdbEhjk9Eg5
5Hc+D/HXuCCwjl+s9OXi7CZMaX++KsSxcOLyYLBOtW+RwGlVsYma/M1VnT0RTEyxaNue84fBdnt2
vVDHBx1f9tdE7B2TiuD/vPwNsd8IDbth93thi8r8l9qJ9qDoPggiJhwX03kn6sWTho9HPgWrpayv
t91KscEUbFIv/da5HyrZDSUFtZK6vwjxee1TvzjY28tWGWlcggpy4lCdkE4g2r/bbkj6RWnRUnqf
R3BkP7ILq5ajvt6JcyStOD8tK5aBY7/CQom2Lh6S8fhP+fzsUEO9KoJTwRM2YCCzAo6Ryb6Tx0nT
aJjwS3CK7kjw2z1hGaB22YuYe0x3a8ILDL3acqIMV610q7P4NMeu3sL4R0U30edbtYRsRDgsRat/
rwhZbzPlGposAAZfUohO07GhoPpm+1emcJUXUBRnc0t9LLMkO3wxdcPwiOxsB/fofRlyrPG7sMDR
MhP5jXKGEb1IjGl+k65t/YwCTNKM32zGMi+UcpDOZ6f93w2n5DA5UL3oDKr42oAp6EAbKL8x1RKU
+CFRsQ6SvBLYk2qaPLeHmYJxxgm6Lw25nHOu4cR5wAXHZWivoBaQbjToak9FzNzqR2goYXzhs1M3
Oo5GeL/BNMUQvXNbMHd9Fn9wrt7rRVlSB2eCQW+H7aLA2oEiPx5KT5PUInTrwumtIKvsidQMPSnS
b65S+e7bCJ+5AIXa6jDcIow/iZMUgeUAEpoS1aoVBVYWGS24azSENaW2SSoXD5UJYLYOUfudyERn
hljlY/aHmswFF5KDLTtPyHg6aeU8yfOWdT1cPfQjkKbYmn5RXomVB9PqzsnkxHGKrvwMCfN7ivPl
jzgzoO8ppA01fdo5jqoMgzbUmiRa6LYuzddFW0Wro/sABJ2oQnSQ3QbPTmvKeRx5zHFHfwnOW8rn
Nk3Vd5b6Nz3K8iLDjZMgjbDMxj0TvrZDhoo4j3VsP/cJz2G4dPT+IX2oBQDYnhNLzCxvpL4o3gNC
xw0VOqT7H9Lj81jVG2bpmj7osZ/RFGv5tgi2fTn8Ihg8iiydTwxn2WECxVbfJUwvPipT++y+t2+c
rvVh1PV+Vp/75yx1WhUL0DLY7ppnzm6xccvEUX+IV81hiu/C9oB2iHwBK/eeShSbYvxLOZFFjbfe
d/Qv73AHR4E9/4Q9Iit42uEwv75l4VkzXP/FRuvSMPMwh2/YsyMW8jeU5lqRFkhhXypU/Mo1S8dv
AEMFIN59id56RT8J8XjM2cU4+Z0qXdHeY01yjchvS3u6uWp+WWnfITq98EotDD/COYg6uK02XuAn
m+MruIDHERLRfYqAppiMB8cgN8hNtBoeJvDvqCZIfiphXs8LRsYL8dhaSMoZXutg1OsDrNpPZRLl
njnZTdmbiT4SOmXzpKks8Jy2U+T2907HGbW/0dAd9dUNVX1VrshmwEKPiUAQQKw/0Ks8g3uvszUY
eOJdF3i5W/0lt1c5waBYfmfZS46ZiCgmzr23GQVDwXP1ZfsfNl+S/TDNnRuhRPHFSqg3GVmiewI9
RwyGgYkGb/aT4ddF4C+oblmdbAVg/iCmXFh1Uek3sEGnAAHwBElFb+b7qyX0/GGkjOloT3xruXIN
YvxgeLdtUmp8MT5Qto+brCET6xFmdXCGsPymTkOKVGCvTodutThUGBJYyvaN3opKj1ACyoPQfApt
0c9ZoJLPn/OjvR4RaUALBwhI6Jy6EVib4QUaxJAnbaTfuT4x9Ee6HStx59p6QLDqa8h8NDpv5Xao
uq8pHeUui1Z7rAmYbQEi+3Tn6HkRFYSxc0y4YyoPL/VMTEo8wmYIKldsAKXk6BuyOzfZYVLUZsDL
Ei5F3oEHndk5AYXP3vVko2/tlkYYemQjk3DQ+hI/2jNpwrIZZMwkqduexv/87YaJ29ACtV04rfXB
GC9wKeaa/1BZjdiLQBAxHDC2YcY2hgX8qXVKJ7sMVEP7n51FoR21UhqmklEF7sYzkdur3APTBGoT
rgI7Q0IvDRtjbs/0+Cv2yqzJO9NO/wMBn9Ln7+zbC7rSaef28a9+cFC9yapulOpwDqLQzxIdr4aW
oEj4VtsmFogSi8ZU1bQL/1EpmbT5+sx0w4hZz5HNlJATUgr0t3rJMTDqgzIf0iqhnkwHqfdddl6/
9emKvl0Stk1Ft3vmaVzzE9APSZoUeXsSj2mRVmJMEyNwvfC/BMfsiO9feIDof3YP97wGudQvz1CP
CvA/eKNTrPkpgH81dlpv5pZWr4k9CAwG4LBIMFbnNpGJ4dfGB4AtCLnrvYdzQ6f16YnJd9OB92AB
ls4SdwL4S0eNAF5HBZlhMtNixPLuy0SRfnAXGM8Djq+SbkH+aSlO3+LMLtBbQHiF0h5N6mN+c+lD
0yvZxld2VsMtYtgtN7eMIRVPFA6FB3U9gMfbml/0hO/ho1+GaWxOqZUa57E/PQuo+vBePXN9qykj
DRy9FcKPCpIHCGVq0eb0q1aJfKRQOEDpFxL8c6bDe4sf02WSecQ4mDO3dj2TzyKkGmmJA0Up9c6R
VFabE+nGS2YeoBjK1dd0kpk7DAVn8DhsyGjeRiFjdKPy1/mb4qbQUrpfl6uEiFOBhwUrJ38cpzly
A/E7EQ0ZHUMHMg5m74njBDgLwlUZQbje9mlnUaerCjBPBY8Jw8jDCTk/bba+0wS3AR0YJfZHbVk0
s9/AVwmTmKe2WuY/cM1R1gKhOKZZLBpQlP7/MSkVihjBQeWm5z1qlsqukk8q1boi4sG4cU9T+UbZ
EQvue6ZrMOjnKHThuc/ZBja9rgAwuezUbUP6SJbAMJvIMWCw+uRBHasCD9gycm0Se97QQNZObG75
4/qQIwMLC5M6/49I32GqjFYmNB7VsbMznCQ6CuTXKGJpZkChEHMWRONmzRHBxW/vY5mrvdhjebPB
xnTu6o5yMbSK7nVLOI7pwb4ONVjW31nnLo8YJ3Ql3OQ/WQ6U6blCmUPIqt6AGpWKaITnzy/c9+XV
xg+96/XmAgOk4N4fAWphzdSNP+kfpZoKPRSOgLwCXg3s0mgcNVxSYHji9V8EeJRoIJfueRuMwmq5
dwJtwd/CmndJ8Ykmza3LdQxfn/4e6ESTaPJc4ksLwp13NRfku1DVJEQi5vofKn7LFFl9SLdrbICE
qRjljNHD2p3E14ds8W2wzn62DJyVGgGZbV6qyoAjqzydpv8mYCpbqzROaKDJ4GYX5lJmDbvx27rV
tjDayY7L8EpQRdudsN0Jy0LmWAf1rNUjL7EBxVghQMy95ZvrwHqo2zp3TOR/f4die4AwOslYYYfj
ZzTstl6NLlZJvJP9V6NVMdAXs8okWljs1F5GhHtwUCxU+Pog9s8c0ndmwOtQ9GBiaDIftxpJNLaT
VD3Fn+aOnLqiRjf5tgvXBso2BTCY/NBGUBz14HF9pfg4R8eetrOpPE0XgSx6yEhyq9P5iLdTkBGt
Q6Jt1eJb2mw5QTrQ3MWwY781tClJw32skSX3G17meUAOA0J8O8ypgo7+bmhZ7ieEtIJRvLaAd4Fq
ci83SdAQIhuGj8+MVYEBGeleZVa1ix39rjLTPqVcdvRAxYJHNZ792V0eN68sBWz/1L3ty0ivASrq
nftpP3emf+OO7wXNfC7zsgidVsbUkEdO3nPM+Xmkbd1QYAml1ATk9jYLZRtqY2Z5fmizwQOzXM9i
tStWwSUpgfGGmEMt3ehWbyHBIK4diMj6Eh907g2gnQAxenWA0osY8SZWErYcWf9k0/tZZQpi7sRh
JX8lXCUwRRqfbTdt4Vuwsv6/UbjYZjzDxJiFcskP36pMjWvtmtIZ+fKeClkD8mGd7JjMZ4Slm1jk
Ou5SqT3p69eyyTvbPosJkv4aGI+RsOvMi2T2XL0FHd4Qe+kKAax6+dCYAlK1YDYmWEdpmYezOQbf
pqv7iJjh+7HNk9BKxNECo2kKsVC3w0u7Sedvoe/hyuyzKECQT0vtVAlBijA9XukXorUf+mY/AQf1
WVVl3P1gK+ykjMUQPsxtgEoV45sirUFTydN9pe71Kp6t4mVU5Xx4q/ZYhD66bqegjX4YLda+MRiE
goMIvvq4eX5qdJkYD8BRT1ZZfZ4ORlde2duKrTDynJovbchkwHZyb+bHDkdYwqU0i3BEe0RF3HQF
ojjZHOTFEXjEuvvAZO0lsXIahkv9VNXuuNxBG3ticb8xC523Yuk9Jz7f7Zd731YZKX/lpBTC0FSK
gI9RdVt4gfWSb7ogDoZRGLcSpPKx3uEWN2YkerugRGTa6S4VB94lUKUuDEK479N7JQRpUw6tb0m5
a7+p4EvexVu5u7hmTGN048cFtrBkYlSqAg4GCL7SxDHPbXMyXFUdSC/MbfMxMMt0TZ1tMJbxlZ4c
3gIQdx7BIfVyFn+eVHo83IxNUpGHLnfRARPv1JT86Ir/hOHz0NAX+DAyLm4N5QOFGt55j6vmtRKL
FkbPExvuNzUPw/VANuPdLgL0OBN6b5qEVCBhQ1J5YrMGTbk9Cp5Y6kS1vXK1DjSudAoQtkBDRFuG
fTc36fau79+JrXEMWQ1khDXglPMfk6MyOA02YIAr6gjmqetMfQ4JFv6OTEkU47w3bwQvIcGkIocR
HKYpswRqsQ2IeKlhzFHqaYHDOiWrE+1psnWbKDm2P7KSsZgPHEnvQAys1X6yKImV3WS7RyNPAzt8
eLvZDSX7kLG0eXA4cUPnUVkjDTv1OTYhxplr76X+/zEqsxAF+H5ZCB1AaBtgwuOynY17DDWz8yZj
1oj43LX4dyfh3Hs+z/eQZ2QHm7t8WN4eDDc3aYgtgoBvXEBoJOZMx32okYgiYK+Tqq5P8Qx7MAsJ
vm2q3v1btBizl2m2t8XRYaLO20IcqVWIe+wvjJsrlNs1Hd+6o3AajPxmqYhiieVYpZMemfEBVqk/
3P4MuhRKtEP554qehxJm1q3i9uIvxI6ErRYI3sB9gmSSgmpAjwRM1HavYUTouEhOOmiVwUbVkxkN
QIplcCSBAetdX4fNRPobXLAc1htmFXRne3FX8zSe1ypfsCjNNPRG/KvdZZqQ5iXQzB+3baBNQPPj
Fmpr0kfCxYJPmGS1pzDj1cPGNYlFs4DttcGH2Ga98wV+aD2582VL/7xHQ2QsAZZLIzPcwqqr7uCl
MHoCcoYo4lhq3eovOiL6hkfYCrc/FuVCUm3TuTUZBy5lWWamvmk12nhMgYjgKp55OOyvf/2PKp40
HerQX88zgj6SU8+HOd+uwaZFhPOq0beUoZkesh7FpQ9yMri6ttsf/HJ6b6WyCkkdnBU5Nju9Xb6q
XtatLPQCkADCbzx2pmUqsUCZyvyjWPSlVjwyGRNYPyBBPdAYuxQJ1BCzkYeEiypyKH/PNzPhCIAp
4Al/m9khXfF22BNafOqQjvDDdhQj/TLrf72HAOGxp2uNuKG2joshw7yVJ0LzU6Usr4/EDsK4RNR3
EKhqjB+dJ6gqDoGC0asWkkzJgTRKXEsmTV1Y37RIh1YznEy+Unc6eIMB2mNACuGEXoHwM4gc3vAR
X9cnUwL0OB8JfkJ0J0w16PHJRav4Qln84gBTv5k/JpxXusE1hjNpJ4SOpFpJfMCL6H71Kg3jkEYl
OR0eJos5Z4icyjsx3GT6TFiZ35uDiF00vwVh5ZdlnUxsrDeJva1CKBZqIRapVhukvOnfXjj+V7Af
xynrEjmPvVljkL2dBca8g+OSUttaKRkQusSalUByTWEp22JJLgH03RN/CpM1FsRYq0S677hxZgf4
cD3WddDncyOtM8vm74/9Q/W8V51/7X4M0E7uCoxACcYTS3VsRTXqe87LlGJO3NDMg8XNhtBbJ6SU
SqmgZOkDJ2V+b9tHrTxNyE17DrEFtj9d/W6wxr753159qnlV0uLM+E96Z4uq/NoMXwm0MB/ynizS
Jm0OrnxPcVjjcUY1BAASnpbnhhzjJG+sNgDyZHE/dE1Mh52iopfm/ZwriqAgRIj1pgd6APx3lJG8
GgSIU2YKR8OzwNTuV/oWtkPa9c130LxkpMydjA30YVnFj470MSHli9urb7geqvF1f7T+ntlB5VSx
Wqjpikaaua4qFyRkZ0QY5CX8JRvN8cPhMbbbSW26BNfIZsBEYPhwMDrz9Bz5AEe2qwHjRTh79BnC
IT8KtC5W3u5X7Os4WHYQqGhEIOFlK1l89kWKhKTOyxtKldqj3ZywpgtAXgbabVEgmmiMuehwS6Mt
S35v5WdYnXU20hWgOqlNp29Ch+BOyu+JAtL2lScMUTxb1I1fYf22sdr+trXGw6fYl/vckaQRkGy6
M9qpj7f2iF6vg+JlvyAytFuiJnNL/sCa6t7Alnn7I1cO+CeT+K2OpPp+iuWPZAMvj5vnWPt74F/C
smsUAoOvi2pbVJ8WW2mhYBQy0oSHl2iVV2UHq7hTPzBKI84PTc6JtPUdEEHtj8BKc84vMPYREa23
pzqXHkPrrGNjqwSVH4Ii+o6qjvQdgdEY9Cdd7+AU+CYlc/7EIBnYfIQP0UlkWfZ/hmlBOkNixBet
fEMgzlIcWPUfx2MQ/kOZpJ+zY4Gde3usbgJXlElXuWlZmRS/GVqKeuZX73BXj2H2d/euS9Ip+8fo
/DaOLHS8RviitdWg/Ipiwt+sZFDAgNL03BH+G4WKMpKA/5lXaiDrkT+bsL+regfiGnCDQHDuFfP8
BDV5iQzftV+Q82lpWUfvZM4d2b/bkMPXfcPGFCjOk2l8Zc/iClZSHANsSQSQ4ZC2iOtknhMtdpNo
ifj9QEgiqw+E3drv8HfUmvuuFXm/52YM0BIdpceJ2IxczSP2AueAgCSBg3SfxkpanGyov1x84664
pYQLOWgyR3W8U/0QbWvtqXV9NoS2edBjIv2deT4NxNhGUNaxd4+iB/qtnCrrT8SZzXwStLTbCyM4
lct2DwshpGnbb/S70hb+2OxhDmCIOWqIo5A4soc75VDYfKvJmfbdECIwOSOQiPQkpZvj2zUZqoAO
QhCMg86LLUHe5W1MlPb+EAez+D0F3P+fV0cqx46neE4YP21dnCN2maYTQ7Ydvr7VUf0XFuwdTrjS
US7veZmlY/WaQR2oCPX1MCh6O4Rgnt6VcZ35mKMxcVQ2va7fmLy8sB4G72YfZCxoOycqeZghMVWQ
ftEcwklT0OGPhCcQdMdv4orwNaB/K9ZWmNy/s75kCYnQBU8D+SrC/oGJThjWzoImv8eOxVh4LqRD
DIE3elAeSNfwEP0oxGvxEbRyscpO5TNHqSYM/wuW6oAAuu91TyZNhGzxizSEGAf1oVFh6F1JG6pk
PaWm1HZRSBKh5pyuQGUnXFYg5/KyCdyhhOB8ahKM6HgvfAsKX+e+A4dRVXEZ9hJHc8A0GSgS06gi
fug8mDSgN1KXcHDnwgrk3RLEk5F8iRdJBx9PlKyKz5nvV6uRztnwyHcpaJ7JndgLBM0THLWG+Z0r
/oqTnM49sAwMRFpc0U3BwtL1hsfu4IDrUFnliT6cUN8Epjxmvt/gTtkM0xJXYRY3ECWN+bWKw1sh
ev5YpEjbNAT2JaH/4q6dtoOt0LGvkAvWLAENYQOxF8u0rB9DCUxzbM7qC0Kf/XVVD/7FWGLEE7gz
lzrCnmBEy8NfkJPVKAtbG8HN+foJHcNqZHqLz7CdhYKqm+p7vl3y6f4rDpSHLR78wslvH8rCaoX/
1MtzFmI4ME0TAN+J9LMECmVzjBBlcwNAfc9R6n+pWUvU/dmGP9WuvmW0t6gOZYFy6QhPX41ikIy6
K8uVdAE/mY+3p7noAW/8kHRoDK4PogPpjYNj5u52gtxJYhUgqVjCcCNUTdC3xx43DUs0/QpdkmAT
j+/WCDihN4Or5V78qsWtbfo0poC79rlkieTsUCMEN8sVMHWT99I+Rr3gzL3/EIKVVjtqgSXa4D6+
RG7yXW+d6VZ838rpy2x1VWtRoZz2o59OTb11AhAbEw5SU44ArKyrsIOwF7l0798qyyflHCffIH+5
hRJ8Low2gLVr3BtBfuWZDLtN1HoyA4IDLOnG7C84/PERXhHb4Ia4QR3C/4RCQ399EkSF2bbfUm7R
izp2GVDETke/0agsYE37FzZeKEuuwx64VMaHGpF6VdZuNNu+bvFxOEKq0g8Ncc3X70BEzqSLSPjw
Cl5cx0NyzRjL2Q62Hgkug4+D3rYyqppOg3Ly0lHqMoTqIo1YBIjM2XiaUO2zm+68vCybrMhOXgi5
9ZRr2PF6lpumGqwie+/AzCYQ0h1RYzqjeLFTGXKWqDv9vpqm4orjMpfbIqq3k1I+VXJT4nE+g2/0
MMlPo34qKppUOURzVSx2cZ8bk+atGTPK51SEgvXMSMGTXVqG+tWscs2Y50uvIrJYpdBl3GhaR7yV
ZWOw6CwDlWHpOchqbRFrpAc299hvUFmpX8Gindm7qzg9Z2rcFE//f5UB6a7iauIVEFZPX0HmqDnw
cEateb6RT6HXueGVI6LeP9I/2yemFH+LIIbmLmblYe6oQq/7D/Lke2qLMZ5QUYKEurZenS4Bagp3
JlfguGYv3kbmq/N7MiyafIjgi2ZZqW3s24tAa8QPsQUuZIO8qv8Es4jP+xyQh+uRCAEpVcud71g8
6HkcyCo/OjXMNCKSbOQmA/DHUi45ejgpcgaqTZwzFqB/Yciq5e8ecbPETTojNenE2hYXMbvhoKwI
WL+bPF7jdNQrzrDzTqr6UFwzu7hreox1BCtensujhlHAs9HmB9kkuaydKwlNohcX+1XyAUEfSlcX
yxPiD1sEBv5+M3hzdqK6z8eli+ZhvqtoDJbX5ASXZuqjgcQgNBhru9emQVejJ5bnlx+mjQYNs1xM
uKhEWbZE24nYInNqJ5ROB4YrJe6EIDcH1ciSIEl++2mr+R96aP0S/OzjG3JTtZKJF7IaeoPbehxz
0NfYSEbK6fwKo8SjnnD1r0CLInsIdbGQWX+UUG2nE8TDb5JnHI388uIC29fynwQabSj2sUqpeh2F
qOKvgyTr4stxiz8B62qlC1YjRLh9V4cuNGb6+cANJs+4X0gyCpKtozSfxug+MQyT3gDdk1NzvZPM
uthX8Xqns2xnMhcx9nIWut6gWOstqa9GS/7WCvE0gcYrBNBM6I3IIILKOX+YgbT+hCVthyNT3Wbc
rtpaeoJTjEF/9IIxLnsda0HZbPcRxfLUDZBA6z4ZzlPFXU4RQ1OA8TVbPg0nvD9fxfETCZ1Ctd58
KLVquaLHJUYiFa5DcuxT2xdyZjmc//o8PEdfbXVaPap6j3Ed3ig3UZBrItvWA4UJuvBPj9uD16zI
fOsNtgp+G9nHwNXHGwmp0BZUJ8wIRnpzXptfKe/ErEL06WBcfPv5ScqbviwPDlKxC/uYqCvm73fe
8EnkS3JS2/RX0JDsD5YwmLV+iYchfE5JQkSBsVBgoDvbXaUxkVWms2Kt7J1L9Te0Y9TiqkyvZ1CD
u1WT7gSBEeCQ5zTGUGKTHGug3yOGo1CLvMW8qB6h8+A76dOjhOi4uUkIq2L5BsT02SMnF/OorsNr
gYV1Z+TP/MYDJgplwF1UwZ/IphmXgl+VYsmLNJ0CTnz/+VXmGSQpJ+PG8dwpC6/4FhFh0Mh4a8LQ
SPnPCq+oyo3ui/FgpCl7QcX9W4A/APITNBkB1KpooHir3RQezSaTtLvfkkN+9uSccU/SAzCRXR5h
HsjDJpYE/yB8LZGG3YYDfSMYzQpLxxFt7TmL5oiFvIDzGAg58Z0KZCRGmwFl8SfYhvK6Ax+rdYJI
W1NajX3ugPq6UA2oERPy4tQlEnF4Yuyy/XRwR6XoKUFx4y8xbAh9YBMJhmfSj/m0+lDVsylvJbuP
EqL45+hbK/K6sIIMKa3J/03OGWp4QobNJrU1r5mvC7GnA8XUBuuBu/DMFBHkTcYJ4r81jy9WmwYt
oJ/qfgb55Wp24nUb+HuWWovIqF0nmvFS9xdwzHK6JaaF3WplZIL+k2fRYu10xevJFsOA5+heZoW/
wPNaKzS8Amgw8CMrbf2jVFrpoEgKQpix4qKWSr4mV+ujpdJOhunQucLZELEvfS1ItPkdmJA65Ozf
A9S01W5UfXS6JIj97d8PCvQZXtwb1QWjN1vp06fPifQo5aYJncP1r01VewBHUC65FS0YuhOj33x8
TH58jXCubNZ4bxohEyHKzBW16aDWXGqMnje3sd3oz+7eXz+OfrtlLGSEq6BHksLFpKY8yl3oli5N
9Da/uXskfYOGpR/b5EbpWt0kMj1vRnmtyDFAsjoxQhm9Jgu6/eNVxnnfccbGQ11tTllH12o9Ikj6
qmMZy2WnIhVvx/MTN8kF4/daELKYKgb44kAXO/DkjJbJizSs6VOlBG2a6MQcwGAYyuCeDMtgz6K6
PGZZYVsxhJMvtxmhHVWJhhfPe7362IdJ+yWFTqAi9CHb96iSCTro2WdKAWdjpltlfviyaF95kxzv
zM6cyWCRTIi3Tw0miNkLvUsFq0kSRPqJwsfF7Olfb9D0+VtwkLzYzFWrmwLCEyfGxkBqVvvCW7Dg
jQ7zDmo1SICQZzul3ZxYThMGjXcxCmb0DBWk8cE0d2mjwjf+RSzFNdBgmAfYbn7AStTCpD69KnRx
8Kf1kV7zVF29MyFHxEpNqljupyAQWZGCWDB3MgSg3xHXgunrhZGO6qWkLq6REHlipZK1W/4Fyn63
UmEV/HNLmvVFzniwcSpkmT2JwXHg/BiHraXXvXCW9D0uGVuVPGQI+gAlFksA7ogWzQKN9bAPove6
uwRd7ytBe6gYGU4r+ySryvg4r3/2vnF7RTm7YQXRFpkgv9MHVzCpz7EBbsWvde6opW03k9B/AU6s
gGTH0moU7nmpE1i1CM4RwpHB2Y0mwL5KRTFtKihJK5cSV0sLHR33aOZgK6CDJZTW+cqJToeVbSy5
G5jI839UOynKmZ5sqr7HErOBzJ3gzJtk2q9+aghyTwb2PZlcOCtSEFhsFblWLVxvNbpN3fJv0SA5
zdMht2j6gHWG7W1xCpW8jy74DArVfn6DFRwN/dN8JNoxzRTfJ/FoVWz6CCEfwTOXneGd6s8L3XYS
IlVS780+jxq8KrpyQAAP9I0D8st6OrJ6NIxlpoBsNwAYxhnxFv/WL1SCHEXD7/c5HcWVXSPtc1qu
TwkdXWzocWjGlmi/YbCsn0Y0y0n27Wywnmot99iFUtLcK4W71JNG3tyqOkutzymwnhUz8LKKnDgg
Q8rhc6SEbB/r4s5ZcZqqrm6kzTXZJTNbWBh0Mw80REI+rkCYpVSsU7KXxkfebeiOBhltcEQWAR7U
w6/yAiwdCtDylqa74yKMLeRlubC5xp+nWhaD7mdF71pbkIlG21RBQdjUfX05J346iw+uvWeEKZz6
3j5uyTThO2+uDtntJpGDE27iRvlQi405RiZFt4X434NyLrUJnZIIeQGtY7Iv6P54ecOdeKQdRD5z
OLCUuratwbtTvOMOnjMI/tTk+9YmXbqBjZDP3FaKQuCbt3qGonuelDmvlS2WbllHOqVnMtusORDz
OzMwOJsN6G13jafplsmnc1VwDYD1tMWVBUKLwvTOQBLgjz6FR4row+GPp9+6j0qm45mTDUnDaPuh
M0HbYoybc86miz2qyBo6WbBWrx4F4/M4wrh4/BBL6Lkka2BFpE7xPqfSzjACYlJweGyK8QVu4mAR
l1Fq7Q1YGX+48INScKGZ4xH2zLuWOpiZ34ULq5oMYLWFkUmQeIwlajXxch9BRS7xsyY+V0ts2xzU
sF56DG19vSj5SBlETEQZEECqqQOVOufhakt4MGK9suWDnFOZm98CenD2wL2Hl6F75flLnOZQj4Nj
xwhmd5AQOd72VlysqFWp41KWEW7ZJtf4i+l/VyLRoOTfoOcsoECb0ip4FIpIl4hmS5rfGubVJuTK
HtPw49rxxD6Cr5fLDhCMmzL3zJnCwxBhebD42uDNrFNWSjoym2f5gLIQ/t75+8lPK24gC5vhJJR9
3oLZWWric54tRuOr/4uo0Nj8vxGaEoJCPC8lbDOszi1SFRDYeyQASywGVtYsFqlJnX/MtoRuD/Wt
H2g3C+U6BJFyk9S5OYlm5uavMKSQyn75/O4by8KdUldNoMJU8+AMu7P+RxlEJZVeO9ow61LHqj32
WI8EA4NYNvLMgp+n1VWnBRFx54ukhj3V6dZM5/MRk6AyKcApTEOldFop/uZ2Y6u96Onye5NEukmu
C2E1qSoWnab7W/LNmI/56RZBfI+rstv7lhfdwYXxWiJTYLj482f3TdUEKDrx7S+JjZrE8ZCw3hsK
Vjo5AprWsN9QFbmBrj3Tjo8ExYWUu7p4VYSundTGrfBjyblpL1gneHh+Nc7+Sd11JtolTr2/AkH3
xO2vBnuc7x2B0LvD9z3WkWeWCzmbBHodLgn0ua+B/Ok5mOymomGMxLV+KFqOARGAMkamzXQWzL3J
f0SawxOnqQ1oXOqxuAxhAeETFMiUhjOK//DeQ6d/t139wLHDD7Wm82aP/Qs++2EXZRef54AXYVmT
jGSw2u2Rxq09BG2Wu1+IUiXFHQzKma0AHoBJnRRSKREH18L1rrandCbJrPih312b8LH6vL6b5Pbg
Qgh0L4eU1kjOQH+msyiB8Rqu+ZSnj+0BzUTCoIESFhG99aV9gwJs+oeoalKtmvirc77Ao8eiVvM9
U4gmIqMoUGv9fHifyKFFcvOyHAQqBcwO4/UM53ouUTC3dgn9pw0AKveZv9FG4mYT9BLX1Lr6HnW7
ydav4ongs9j1yU1hh6OnX++aiUn2XeB7JUPXLiQpA9a52qo+4Wo640bZ1J6+NSyvZ78nxh4+60YS
mFdXsVz3dGSYInHeB2Mw8QRrxFn0CRihOk6EBWH21suH2Bk7AT+1haMGy4lHyuXEnFT+lFnjCFr7
gyzYytNCHubjwtDKzfV2zNHC8OyRmLbia0zNiapK76yRH1bnynQS3JTiP3EnHP8nlNz8cy7o/WMl
gqs3XB8B/USatNC6sIAEfyR9ddQF/YClM60dTL5LQoeeLu6AZ0yp4cjHr9eUcoB3YYDL+6FlNbia
CIZLQ55Rz/Zx3IBMP8Qqecmm6vAV+1vDsFLH/QfVBsy/htJJ8z5OplN3g3t+v1ogClUTc+kfaZd2
13nqC/C3SxjIic4NuNrNe4wF6nozO6RXvp1Od+8H6b83wsLK2Lx4fnwbrsN+Ok5lB1uaRrSN0RWI
Zd/M/VVsXRVCo+7E0FS50MrlmdRSUpt6fBgE2OaQLkpcEvhm2FdLb34piqv+ZWR9jO5ZLU2Eby+3
AZS++qD2PA9/kJjB7AFUVBA5jBJmoV/LhDU+zi+U2T71Hry6UQMZEO7G/+qmjDqQFz3oDH7qDY42
uBm9RwESOOKlH53vs9Tbi9lNi+cv9Dv2YP+i41Rhrf4EeotaGPwTlXYCXZbrnx2anUxnOi4TaLkV
t9s4T511J52pr9DLTjSsTj9z6Jf1SdD7vXaJwg/sl8cumnrK7DXE0M4MB5EcbDZvuzlTT/5sns51
OyKesC7HhLFgsdNQX4JOmfi6e1kkQ93B7ukV1StX9UDJhT7J4nrKJd31yO+fKmmJQ2zhgZpCrQKT
eRWR8+o/rj+ZVp93bu3PkEcVfLNUSCN/NAgZmw2L9j4dqGrIT12ZF5yvcMdrFyQimxTZ3qWqmHCQ
p/8mZlZHU5rGOcHyQPJBjp1DU6nRYD76B25gTU2GetpAtDyAAs9h7SV5PYRV+asoLpu2CgsTiYmD
4mPx+4DWfJSPJ0gfNWP0M1tKMoLwMkU+xqWBH7lm704xC/Rt2F903s4PipZY0Bq8Y0t3OUJmsjL/
20YqJLN9Uw/rphZb+Wt/5HbVzOTkM4u60KF+s1ab065fpRxJHAtokyyQhd+H3oagyLrrYq5sfPso
25tePvdu88lcmlNc3YTVhPPi5HCOCSkMKZJUUyqukQCwmBNDw3jaeXHFhMS+0vNck0jRH+kkd33y
xLskD+v3tuF+qwzyFBBm6o4JWZgxhLrXlIjq1t6dQIO/ogOcV8jEpJ5O26PyZV8SRHgJ4pgKSNYL
osN1+MXvMTD3NxTM8cbaBWZGLJQeLwoJCCOrChwASZPSy4020c27j7/VAqxPW1/gStJZNS9dT/jL
tCFLSP6doeshTI6yXtAz4HQ1h5DAmLHTVK3eqPID4/EFfKgFt9YCMqkeTN30/GWC3aTmJuQK+c02
18gdX/YdC5V981jv8DCb27EPbbsaYbW+Izh3iaWShauQG1hPI6HSxbWbBDY1IqKrU5zE78az2Fa4
weXteaKN6335VxP4D52BWkLDeI/8GesIM6MK/YULF6KnvbsJKkZxrMes8VAS7cnA942N57u+DR28
VPOupQEvz62kqkkqxaUAEoiDZaywwT5EkvNE2yBJCmc3kX/iTKz9sajwz6KIqkBdRJZ6zgfCURjS
fOPq5qmfFjnEzL8KF/BY5qDdP9kLLUP0WUVx5jB0jYzoHgatmdNjTXyKnxuJ4Dn3w/gnZKnnI3qT
vJYapzhFdGd/Gef8aAqScJCAaQZWveTp02cZA2V8jqjBa81gNpH+LvNbmaSekQu3mgjjMRPPdxTX
C7034c73qpD3eTohpYFRGu8S4BrvEOIBAT5WFj8nMqMghAqZMRqxLaOMPFiu/sn8RJSPCSiEv9Kh
+7FsdS+UIYXcISI687dILrZlfELgGGEJaA3PYnPDMvfRTyL3sakZh5WrZ0Thj/JnG/UBpOSCWxE/
nVE3XZsfkqOw2y/xN5NWMJ0AWRMVRSZtGKsVDW9q3P5j4+dBpXIvIbtQ5Qyfw1YZBB3CZMUwiPjZ
T1Ag5i1VUzYIuwaEmZr8Fc9p+G4H+B0M2VIBcuDETlC8dDj5L7fDD9tg7M+nDeVxunT/q2IeVMK0
833kwEfqVWI3sLr6CBFYIAKZSzKiSM+FxuAhT6nabq2ug5d5Pt42auYxWPMuj70bEBBjjaSJUM2P
zHaxmq78V/BPSUAmsp6faEs33gnason3Hfa0568dFu17VZ9nwhlC2LzMw4EboqUc6ZnBzRFVw44o
B5ihmCUC8uk6AKHyTvegwo8y9KUPtxw7RSxSJq532nkjSRplFg7lGXx3efa8n2Tyckn9TaitciJz
h+krq3GJ3kDgfpd13vhuFfVF0pqVo96SFshnz8C1CaHhb6tD8sr7PPdcdAAw8z5Sy785DUWIazH8
87WJNZcbyELqlTlGmzG/0OePERPGOryMCpqN3J480M+pSnkQpw8+bavMjs0AMmhTsAJCPau910cG
8pIfZdnXLO90NAEWJun5e44HsjMfMNsd2RO4tazN8m0s3gDHs7Do2ZfTXbtzwSLDAzCXOMJubkWE
leRtZ01C+6d4tLL4iKrpe/ZaD7vRxJi6vE4r3/D1O8TpGJc4b6dRWhF29vFJGlYfAUN2zUNKT5Q0
oOHpKH3tnK2TQjiZc7b+9aajwRGmpkFrb7hc/0LDwda+IdJrkwOxD+qCtkYUmKEd77IOwV9fEPql
efdgRrtyWq0HZlo24C3M378LS/NXRKhhhGTxa/dG0hpzU7nEZO0MWJUfXIgPed0eZi5wl73Ztf+F
L0lM4I2d3+877rcEXL77udWWu3strasnVrccFmL+xQYyJAKmojNKgGVg567kDbPIUP/eRUMkg8RL
V6fwvOtYuojzEU25aWxvTvz3jDMYRWiERCfp2Z789c6bcfJffqz3pG9AHZnnarC/HsBCGQmHM3Qh
e8phV0Pjxb9Bky6xE8pJtrgUJT5IoKtwHE7fL0sQQQrWWy4yEz+HbX/ADMCSZi5UEpYBDXT0v6oE
OkphtgJVp1V7dyD/FTIh1S8vd+4fs5ugvgckwlOT/t/tMaFHhxpfyjrVlnK9Ffj/qBJHSUzooX+3
JWc/dX8LurLfzYUoYM/NPMYUplE7P+5rRx3P551UExLH+03TuTnigcwtHokbd9R9XIb+6t1rz/YS
luWYbjNVD0b33GI2UJDVV/GiUQ4ouUXZeeKvE1SoIuRsLVZSBYRfV+o63ZZj82j18TwKQA09VUZD
9wDXDqnFHdmY8pRWBDgl52R0oSbw+wu5JNs1kv89yThX4lXwpTFQ74hzuRjnW5wulu35rqP23Myq
Uq6XDtsToXOkinqe9Wlh4ueaoU/sWYKCdev8+r+PhL1JayPHNYhH6hDzrmJDgfzLUZtwpu+ufVUl
1e/hvmANS0beu61XacaWlWL1kM5ppUuEUkpzJRsF7DdDfxluCvuAQiqj3KBwuYCQZLf15fyplyJy
SfifcOJTQp+mZ3dbH9kZRXANdj1nsy521ECVOM1Qcl0wd4rhu4xQpWFzQk6CJIf+qGRUbFJ4o8Y2
DPo5lrDQdzaK2mNibbtdZGby+j6sNBomMp8eSBF/AQCJI895vEXIAXBiGT+MA1oLrqvmid2FIHNa
6lZW9TVPg9k7lW1XmeZEKLlMer2LoGkhfUfYZ4ZFgP9iF9RjLN3af0VABpFHJYxIyuzEj6Ocsg9g
atVnOvIdx2MMrBsTcFXpoMh5VTq1YfyvIi0SHSXD5oKOj1TW/ZYQmwNzyNcH8TKp4cW0fsUgjOSm
9O9qDgy/7uDt/GZ4T/UXIGPRfGvZ+9e3JX9pnLGqJTbROnEpj0Gs0gVQdx8eR4W84z8RFS9Yl3Rf
tr9EGUdZtAeyojV7SSaf6bshO3OUUlzrgL0S5JkZehomzjqarDTdLTHKrvN+IGgOASBnZLw2lG8l
892c3MO3XGshw13ti+D0oFEVwCqzkiWcx9oEcMj1qlyf3lBs8bYkX8FWtmLeDk4Dvw55ND0XgWAJ
oYncmorj12flsIv65Miyv8iNogLSESLm82uxJ0SoPkbdNN9o7VJLPFOOtxVOb9STcokEMw0apfLn
byBkz+HRVC6hnisfFZ3OGbjs5E94KjHItBBReyg6yol7uc2ohwtnueAF9h3VXtmhoW7ascoxdval
WIMTiD3jvJkpHsHNyRzxVqyc25X7KIYielTB9WA7HhFN6eI8FjwLbkTryah+gn4Hmw0P4TJ3KLGj
W2UmdRiiEXpVNikgsdeeJHjLqn79Bh8hgkSrUbK8Iyz4z30P4Oxq/xcnE/CfatzkHKYEEyAeQo9w
ScbXeDW/gBK/UX0/eHBcmyeQ834SzsBaTbwoVHl6s6DmCEXN+dzOTKdKDSdZ1SxYnPTI3nwjSiYR
Zcf4V+im8wd9EhEEJcWDQLpoDvmSOOB8bPmOO3+ihLXvKp1Q39c2XGSM7jB1SAxriVvxUsQdzJ1G
B0dn1L+Uugs4+g+7tdGJhDrMqMCNAEYoOhkJMTSMZdexCPE3TBeItpG/TLa7SkKUHVzRiC4LYy4G
9FlHnVWk9vYhpoV7vAWgjwRirfMHLQv7DviTK8RawNRrDgWzIDa5UZcmSV81ax6UL13FSEnfVIM9
V25XkQyTPp2rWCQKSKIS9OnNLq6vuYzIwRlDUcAevTspxRrZxGy3ht7UbPY91mLTpcNKLYggu89l
FBRFWP6SVlmcCWCVvB9aUYGSv8QLrNIPtegdPjHGd/8mREiLHEP86IVacNtAgyBhkjU+2BwHh20C
AeMKSbiAvdem47/wQSGxODgmCZGbh4KTUpGRGwIlGOK73pXz3qzuQmba2RhGh56XO5y0YRfOfFX8
EmQ70hrtPCTXrot/nxcxUZmKurjo9waJGXADImUBmuOG/mbS29Ioa9sP1jyEqZwxW5NC0EKDGS0C
RDP+hCIkszLCR0xosOrevUhf6fGW0Qvwlsvh/oSv87N9kp4vbWwBTyIuBCXik2shC0a4o1B3gOBr
FIX0pOe+KBqJtA5xx4TG6WQhl/yUxUZdcbAi2+Aog31ECMPX7+mXYAcd6ZAgojSwusnXNQkdw2+6
lfpiuWTgsdS9rH4JYvNwJ5EyyjhYkD2RvXAy/nqyXJm/ggxWQi5UUUQEXKZrFg6S+URWkN73i/22
nSgN3VDU4ryVOuUlULWLT3PqfoVppYtm8hT3I+6q7+8OUDvOXx7mO4FTBmmKoP/9x0Y0v1nPGL+d
UdUwL4iGlKi1cOe7AWixuo9uoEtvGB+QVwB4WlhYngkUjhImP1JbGpHIrzcAffuB+Y36RuLTaD9b
XYwm1yCeWs50t/wXU+J2x1kTLKF6MVEebgqH9dm13hG4/HTz94HsbWw+RfSn1352gK7Om6oGPa2W
Bpte08NHT89xNJyZUseBVlaZGdbyqx6aWTEKb3pkKnCHB/26DBvpKD/XiyYF5GtkOVbqECfHKMuS
rn0ITt1Kqu5dTv66UqV5vtDR1NqJpY32cGDjJIaIYetgiShHG62zkUjx0krH68n5lLicK9s2NNAl
kAbcZgpXFOAxsz8sWyrxpf9OSE5E5zHcMFDDsR23Vg9yCmSYkLCaca3VbX8kZRQS0rTjeX5h4fyS
uVwNJdYYzVBK+TecGkyEEkzoz0T6AqqkQ1/KcsQL5GElWbBeqwb++UCBTEXq/oXpM6S2zWgpn+MS
BzTzWubxUo85OIII68gCGXt1u+rs9Y5/y1V+En+qC+E9GwAhjrzhyiDbNIxLV4uAG//9K7HPqVs9
xG6V4gBhC+bRc9r8WgGuW3oSWntkD9X1N3rdHlewBdKOVsRz/gVhMmncTx7hygx/uNh70b4weS9h
05aMtrIhpQ9CJbGcwCYpSgO/Tb/cGqx+F5gP/Dj4o22S/tOtscEGOSLMjB1CNuiEhIweReSLJz80
iFpqiQaqM0gbFZRcVoJC0+BWYXDF0xUN5LWpJjlHQdEerfAFIEDmaJ3js0gAptK4AZvoVPHtksC6
q1IWMVYyVQjUFZRhT6YgI9vinJ1NHJ6OdmlLKyJ0pINkY5YmFaNmCdbedTqgbRqT6wXbKW59DFvn
JGJEP9EFL8oNPmztgPLjKJA+MJpULthyNB+4FexZlpZnDhjVk2Q4aQZcw7ZQlXG4oL7+RISA7LAp
w4yrz2HFO0oamo1ki5mAPv5zo+LJUjCdGwBFzuaiwHsPAOkv5gcfhxZG/Z8LId1fEV31QrDmt1fG
PxYY2sjd+WbVB0DviwFf8WiSQc+F/OR7nhZGM5dNT326dqFB7Ean0IKB135+e0FuZEG5l3OlUXo+
iBcKgKZHaORyYzkY6Wbx3je/DwLiPLU7SdQ4s1zoDKobvwTsU4vPDBqsZ8X+96wiBDRUGzOnkdoc
CpnH1dBkh18j51VWHEl7qmWVmSuZIUmNAJROFcPdZaVN6GvA312I3LTPuEDMjUr6z2agTl/3iZ6h
FzG2cCSwFqpp4oGnP66FvabNudhDrQzLs8ZxnJOecWGX8Typ2KNCuYVy/EDKktx8xCUZQDQg1zYn
glYG3U7Upz+NWlh0e3ILgf8w/HPEzS02+uuRbmeTrnBe/qtC7fFuQoYoPVUDYs1FrfHPZowT6Ncx
8eW74/Hkc8qqRweGSU9Rqn65gK0Y2yZ/Dw/0L1LpBGOOmmUesi2UQuGBI0CXM9Rc9aB9cDz2w1qe
omUGzQ+vj0KrVQzGkiXD+4pK0IK9faYWtu6EvfOyiEOqzgD98qVgbVlS59QNDefFs0iLrra2wyp4
RAyadlLqJOeobjeUqRsRbHjQhJ1r+R3oXUnGqluQoESSZKUTsPkBDkL1Y/YJDHXq3B7wGP7rnW4c
toX02sbYGosr474+BjMvIUOHzdr2+Wsd1EI5lRFLSBkmmzJmS6BXiJJCOjS7JkMRitK18bowtokX
9F5yAR8pdGrOZdYxhbJQ2jVEeR0RWZ9XF77aTYWwIKiW4ZGClhtxWEZNZ71YlDRtasNnxt5XN3DA
Lhf4w0qmuURdGrUtqDBIhk8AqbIdNwHiPG04F6ZdXsjJw8o0F2gW0oshD2o7/NlFJwAZV4Z90dVI
MuPbkNAa+tO2q2mUBeHtWxRXvSspJpzbNG/nsSPRA1igXfMMB0q+exiKdUbeKi8iwdIqBMvQeU9b
17PkDU1D8fIr6lpV77EMuz7v99HrPozLVUMv1/L4JRSvJ+DZbyQCHb24aQkNDjqhWzHb1vkpX883
OdZn+3xS9j3ZX/WQopsOLaptIVzULodpog1lBnespLEqav7aMf7bHu0qBEqx6s4OPacpjRh3VErQ
osk161BPLFtfAVdZlstLVfcOgJztBPSm0pEPWoVbQbNvWzd2vb3yEM62HE1Oq+bcZxrcon+aTjwl
JwJBw1vTKm/jrYbb4rAMy33BJlUfcEichQXD5R+8TrPQ1dtkfWr7d1bB8mPMHOe7sfc5d9Vh9pz5
QPf7XQIXL0i78Eby9iT8sqfQd4g8HCeNYGR6lBpkJLu2ByiIkqs7BSOG7cL/jLtc3eSSGTjn5EjE
7G8Zcdg/0kROnFPHsHfiAt+n/Icywio1QfjMVVohfknBe7ayJamMOVYMUgG+AdVsy0iapcvEyG87
kW7s3GAcXXtiXoH1bEM1LJ8qG+onBidjIceGwk6N4SUGguStye7J767clTMwDLfO0uZaep/pWjxZ
H+V3hPE04pDDmW7fPuh5zdhUyUMX2vJUXzDVS9j/74qe0qkLTcPYqyEhLfv2QWhUDrN7h5RpSSck
IYDivA3B3iA23XfnHme/so6iMOUm60HuqxSZuglZL79ZlfiQ85FwZP7lEWM5/VJDjytbk2o1Kqz9
Jfc4Nl6ALpaIw2fVSpzBA0qEgXP2z9J/0QXxn+ZeGYdC0RPQTSgKbKtZ5M0wOQpTIg+SDb/5hcGh
+6xDdf9MddW81xbCvV8kZFv/cMcChmjBENRs/RFRWzvLuvy4vbtQ0w6d0WuKE5Hb4srnrqQMyg7Y
ozi6g9htUkqA7/T7EZ6pUAMd5orO/unqYTlfYxDeEhvA1Z3t+slJa7++djowybrZtwOX6hGzU1uG
IvrwRadfzAH3UDHjj8Ta4sF7nNRCwOMDOVM6c+Qu4K26eJzQnwwrvgG8sa3ySSWwdRaDRvjSXU9I
t73dyz9q6aWcHBokezExSopiLPozOV+zNoCoU3HdIP50Yat7GSoxKZvL0QKdBcE+k0qHmnYivdqj
vPLEyfKWWGP97qjKh0YMnmRu0vcoHvlTQly6ljfmfvGlQg+RXWNgDa0jvMUvZAt7H75BHHpI4V5c
3tLQvkCoiEaUC5LqHqGVFpy81nbxA87S5kMc3pvImMJKFM1Ha5IBGqdUgYPfzlUXdW8PJ8+q8RJ1
Dqrf4Xl3ByWmoxCg/Qyxto1LYoQ7f+1gWTrfLOHdrtsWe8GLvncYynk0qNTOyK7rSWZvBk5JPCUM
maRwvaMZkmuqZh/N+H7BvIsXraOWAnlb72KiAy9ipS20XFif+Wm1sxhbaZqhVCqH0yaD7SM3++9J
NXebOvnz79QnM5HXknYaSInBJs1CQ9GaXHsL9SoXV3SLhd4F5uRVT7BuYyAdSAku1xtFOBhL38Hy
TXeZz6LgznA9zX6jnJO+5MeIo1LtqlBm0ZidW2IyZdD4CelzYArl6FaILMjl6jCjlgRLWptAI3pz
C5nxTy92DWq2BSMvGycz1haO7PGWLAn6thEBrMIQrSqQLFGShnyPv5FcVi+IrdM+676jV8xE9uPc
7hZRqgKqpvO7SnMdcU9vBNKcQrYj3ufveqDs1ReJFBZj8q7jXVGGPRjFNoPS+cLNBOq6dbSpkrez
CLCqmkG77hoHVu1Er6UIarcaeKAq1/3uBAO27Di8DJWgKocwRbaybhVmzK0xlj/P14ITEnEWdUOs
ap+gUWZ7JIodhp5GBAzOROJhgDV0dNvxsoQ+cnPYyfYLYdj2dz83IQM8L8DC7F09EF+R01LMr+Ly
Nn+90gw+u2oXw9mhouLF1/+kx9DUCBgAVlCTgbnI+19wDL8oLY1R6bW4wRXOqRj43qtXYVWhsp62
35OksMkpr/AwEqn5FMOxxT9vOBvpsGTLCFOJ78n2JhS4lvAfATh0mOlEbiIV/nMJFWrpzD4z9iAO
F61iNCu4BHQdRGUtNkiLZX+7EoHNRYWeIx1Vz+5kWxPCC0dS3y32WfMjhijBQ+75lL/aP3pleO5w
Xl/NdUJByMmMQQUqRELs3+wfMjvD1RwI9ayR40YYeucQsOi93yvJgk5ou25Ubu/5WSyuwQlj0aD2
nLM1um8hWTZNv4tjYcS2pTIFG5ROI2suKQDBwne848C6HF43iL4VaKYWE21AFiR0dwLDif3bWGxX
AoDRLzD+MOivhd8vU2lsg6qseymt1WUokiSvSuI+J1qbYBFYwyWefmwZHlCtqjItj3L9G4NSQ6QZ
tx9LZQfDf6ncPukESmxFkpiFNYJa1xJP/auDfWAR1bkiRugltZVb40LRJ/HGW+UchGCeHuDN5SIK
PkxwFAvCNyIHtpnzOrtsuCTdqxcg5SQfq0X9J2Gll/RgIR1tMM3fcb7/tSuh9J0LOOlPHr/wxJEe
BaRAA/Hev/0bTpuEFSyOJf/363GaIOezOe1ZbVLukrM9+Qo0WtBH5d27IDDD3tw9Y/g8n8Nn6JSv
ECqDf79mo49GGIPJBkKLNhPHvHc/7WrBn1vvpcgDs2t9Zx2E3C3fB6xs4/TgQ26vLz4s7CbT9dJY
jg0JGxcWV029LwPfIX4x4IttZ8j8QXH2kBn+/lKrCUsoxNHJEym/5bZAHLRE6XPmfeAktBVYKeap
pdiUgOkQi8yig7LJvg42ioP9ZjkxUsO+s//Be1uvAGcUOVzkRwtkRJtsbRxP6jMSt7n+kcYJYFZV
+HB4Qd2mqnLiCA8R890FUB6koLHEj9VhVbSz8YaZHA/uH6p9orA96YviR8GklgaEGxP2spAssr2B
wGgDfgBK7+f4JRI16MZycHMnUfAfwd1FtYyiefaiCuX+X/vbps4D2K2WI4VUvxCHgoGNoHjTEwMO
GcxpPv82BbebuET9Xu41xupaz1RzOUnWzGLin68B8cdmaAq801XsIGDXRdfz+61zQqreeQjpp0kE
hXK8TBSgRyQ29Cl2TPNTgWImteAjS2GoLUEfR9paki6GmBDRLyvAbhCHiZA10FC85i3MlCAj9u3p
C2hoCPDKJQGuYf4MhibVOSkEm1/nlVVKBIKYxP5+Ma9/vpw5w82U25SCnkdyqfPtqL7eciyOppe1
i65DthFtajdXmRV7WlUUAb2MPzxqYqne4XQCrT8DRnOpqrcC+2yG/YCLxy7Zm8XJkbUOee13Pj7Z
JC2/SdRGzacdMxctp98hEILkQwns4zmYZpu71G2m3WzQz923wAQeo71XVOqLNp5V32ii9Iq6b0ow
Slwrk9Bkdi4Up0cv76NcwOy7YT5M9HHn3sHH9NWzzSdNxdEJaF499ruWh5ZF/K8h8iEvAjlJRDI6
Dwl/IxAxR2fgcjrEHxX/hthKqnrnP7gKz7p55YgM1vgsb0ourIcVMhKiGNsCYNQbTeECpNr6cM0o
xyy+YH31vpSqoPduF98TEHqC4vk57sLw+ZBgbnsBS0lwSy/5khBbtcbtMMA3J7oUh6VsiR2VVfPi
AOrBq4+0WVnAQdV2dytkNNiws/ggj8Ycs4d1TVWSKnzarxUdZeNsNgemYuoWOS+XhNTSlDvToXTA
T0RP/+Nps/SFWKeEoBW7zbuqxI+v16iItSscIflSgitmmARlZtBI23w6TqkaZUoihU27/jCs6drn
tSly/rXIuuk8ESsLKRcQDDryfFDWyPi5lzTiqcUxde0INEhtpFZCqS/QZbsiG2PZz0ctLK52G6Yv
KCF6uhAUmX7+265jt14a5uFARFjai1BWk5Vf5MoDtH7e5jQIXeOn4DX5VSFIRRpb4YMCIMzsgEt2
74G4War4y5Z9ETSeeyWdCCtvbou92LLx8oWSMIciSkyjYLFm4tP09hQrK552EeFDzG6uQcHk9J1k
mdbGzL2KsijYeEGeClK+vogfPPBKzCAejcgmEZDtB7QhMZBsd7HMS+5qttCajjE0qHctee88Z9KY
FfIJp71gCvGEyuuTc6YIhmnLJWNK6uBdp5YP8o6z/5hFye81N7Pmby+z4aBowMtPqoN02KzxQd79
D22/aXwwQvX3fbgml9q2/pTPitApGUyMuuGWQMMM5O7mwlOsjU2zZ0yJM8Ii2I0y2tR2Mhu7IE7B
R/2kOJIItIrqz1cStlG+mbnJJYGUL96LLQtEm40eRkvmohYr/kfnJH1Xr4eMMNb/MURgQo/DWR0d
UnfTmjfS/kxMvupfsysEr4Ai3rfI8SWV9K/V9u7SvL8yX6Nc6GbJiYO+YnsiDEyIechLaFo2reG7
OGzA1rnitE+6IVYehE3CKttwY22fnVTKC1LGJqvoNA/Ync9Z2M6YFVYtAM68B4p+/hPKMQgyyvF/
hMwU4e0ViCnBH74CzA0MSDkKZzvJHz3cwsuqX4DlPMOy+Gpa6t7OEr7JUD0LselnitPrD0R0WP/c
JwrZcvYG2JUKyyxMI4AgSmII3SOZlRVVfYPhLlWcJReSlhHQfsh2TXTqMmg58a10nOjcEQfU1yoJ
ZSaZbj2ghM+aXZhwdSSjQJQxGkFvSaDF6ZFRnLID/x09rwKEjKRfAQyInKPBFJ7QLrPM6e2SBCpC
R8xWRQWIDbP7UudIbWaIOM2VEVI4pV5FZUaORLDPxFgA0pLHc7InNyr31AoFDuOOkUiLLOIljme5
PCfWMNnXuPBl5cOTOWfe9NFPl0U8Q7QqcrWD5gphFbx7mGuCTo1S77e3f+3KxXdKMg5YkT/+1BrZ
ESS4dy38Vc3uotV6vQb1U4giRfSG6lRdpltrPLU0I0UfQTbMEFp6paPwkRyYXVDTmixT/Rbvfjvm
eTfEedT0JSGlBiI6+XCTebRSsm7rloHP1ecRtRKbUehMquEtA90gWpLTPsWcHawc5OB2l4FqXILS
Z1j2N5whUCH2A1VMpGitZY/aCZannZaRIXyH3Gd4C7Kk69pEhq1LWftmJJYGxqWT7U9aAynHhKM2
n2h9Q/RLVebo+MBpwoAgSUk6NmtRF/ur2e4V4XxQJj0fdc+z1eGrZxXVZlLZGLamqYKc/50WsUMN
lpb26d/glHGEOQREZTJzAaDmIG+26wQ4HSMMLneNI/i7o5wLZm2RCJG0Lze6m1us7OUigZbww//B
C8Uswp/fiynKbXYoMT8NH9TZj8x6cYnILgAvI6h3Wmm2JJn9m96Vou/2m39Za8Qs5bj7MaEz2lIt
OnooXXFiD+c/we4kbWy5Lc0pacH+JfsnMQGgfIIxhhxxHncm7+VQcnMANgj5/8OfPhEEAFm6iKs3
7ynPgS3HWSd74Qio6yBb+6fO/38lnElXbHPsttfBte8tF9r52nxcoterC2V7s1yIphoo1Q90U0RN
5moTzc6q4S9iFKjBjQJLFrCPaaa05tjJtImrNP4KbTsCEs7zjDTcjAxctFJYfWKGmeieryv83+Re
lg7yqneOc0q+gL/3VL/0sBtnH5JpwjQZC77IZccws68QvsCiAch3Tm8GhbRn5BqMLwDcd52mLOTH
14Xvlaehctz8okWx9FY+t4dv8KOGuCYIxKqYd23i28RYJSxnI/CzHMpI/IlFc064rNh3WDPnvWYO
8gsYWCO59B30MmzHOzt5SRpQ5QViZaUbZOXZoH23p8kMlDMJaLfBf9ysph81ftwHSjJGgscojCyo
ovQqPdZad6qIf13xt6Yf24FPFMuBgmrEagcygMGtDU4fusY9uchjaBDH8Fvu9ZdUJXRu/UyL4GRj
sqcketw7Fv9xDUg0Due0b65PMgdqeJal/cc7Oj0+3Z49PHlwhj2kiWMv1zeA5PzLRTpdhB9Xv3X9
2XdQyacvcaEssboEUZkLYX/MHJVh0T9VYQ7IW60qOwjhRPGqGg/oYawvUgvfj+y6fH+5qsrjBi6U
FP+qCIA1cTBDsSjzMR4Al/V4gho32BOPgFRAODIX8RgILzgS4pgRtWg89qsFKcC6om8DAe3p5dev
w+pXWPrUa4XjpQBA8vG13gUbuvfZ6Q0JepHhNUKNT3P4z9iKp8vS+Rv1A0IMitrke7vwS2yfCMz2
cZSAlDJyt4AWZYCEYw+T4cFigtyxF40lnmlIImV2sGyiErrrK/xuHb8vTsnVMKl1Z8BOk44DPiiw
mvHDVn6fN/jcJ762ObehcRJIQsfBn8BcVEfWKSgfZxoed32h1ZVw71hnbRy0lUUaGBt93dnBNh42
p4vWK/y/HMuUjyYs7O9enVOmrMsPtalKPuwFSxN7MRkhNBOZeveGOtBZK5AWCGZMEHVnJxDFJTE7
+j0vqGzm1vy3fYxXHlb3YEK7X62k5KIUrSSDGFJ2Kgjr1AlaRpViR8pk//fNxRnmG0hU+5fgpVtn
+jWSxmanDnEM5SWgcPOLETlxFaye0VpO0sUChkZTXJK9UK7su6J8AZu8UKhJ+bQpEqsQ4kcg3Cfb
0qj0QuHtGiu6+sx2ky3VBZWLiBZNasREKzT8kb+8A2wsoWXPvMVB1aIrUwIMQD3UCTkqWP+pAjzC
U1lagc0wCWyOonMKjZbHFSKeQQKMVGowPQQKG3VQLd/WzR8z0npRVnQb0J0Q6UlajFP5qVN4FUl2
ljiOCXhor40/IldLtI5hRSerkeFCzY1eJG+hCmGV9n/Wa5iHHORqGm5umPJJTDDtDwfkGlvgTXlO
3pkDtDy8+pHcebjs3IaMqrrqyH6BnfcBLfeueXGwSlQbyPTz3vZc/G3yHHNlZjajMYy4Bm7KjCI0
Qnwy3ZH0B+LpLrl4wEjb4wSUEoSLXv1QRKEOpA8olYkGhVbBZb+a6LXJT8AlMOmTVhU+E5SfStP+
T86iIBmlD9m0PnT0PgNLG2uE9g79SrsR3atrl3E2+Je0h4cHYA/AAxaRGOVHdWjG4FwNWtgzMNvI
j99pYJ3gLzx0t80EG7a3hH3uhcmhlIUdPA6drUBfhkKn6LkC2sY+lXwRMuweErVt8AQHuQRfTE6k
xYg4NETZxyejryHg+9Pl65Mk4lWLDraLLjYj0vlsNk5D2hCW5WqxsKoEqd2HQNCx/0WLOjiTXuYJ
l2YaX3b7OgtFI0lFvkpp43sRkrXYDBl07lCd61m+jy9CI7b9SnMUA5TDxutTyNBCJKIomdgLLovZ
9JlAO/hJWxRt3IpHz2mGcUcS/Sy6h0UlpqdxZ9PwJrxtcanYgku86de21Tcrf5YV1Dik9VHk+qKE
M4nRzJm0DgaO5P5Ziwh+ydATKvPeMuM/DQ4qwCeqaTQtz5i+dr9XDC6TpQlXs6Ao8JMCz9yYzt9Z
H8v3SRHOyl9lvboZ9cuJTUXvztcgp4aHP6oqCDIXFpOghu/C9iBC0ClSVi7mO9XKAR+v47HpYRO1
aMzWB2Mh6fl++xsuLPAVe8AYiGL3uHjbVbT+0YQYa0e+WJ1nykw6sUjHAJEobnr+7RmVT/+SCg2X
UXVVyp+wF25E9y1+LOpb7HAW5JelbkMDn35uV/hwLh+vgIsxxg0WkpRAzyQ6l8aSiTUNQNbhZJBV
A0uN+giHJ7JcliByBUX2byquiuuxgXQkDqy7gbLo/YPWO7AiDpG+2iwrEns1OM9AXqGhjN+i6Xbi
ne+z9QBaaLEDlwutJBX8mx0m/cech4oLvJBBGDHf0nl738fDt09LTYKoQAG5HC38c5exd5B4Mava
795hKvK4zHBDZZph/X5WXmiq8vDad7LOTarWk//szvyirkVhYsgjb6kby9escYWwNGqJd7fVSOsm
OjQ5neNpFqTyVIyfodPSaX65JNDDdsK/EWxF54YgSJ5ml1hIT7fzKE7jOi1tQYYamyXve7AO30yt
08USWKAGsOiUfNKpueQScSglmrGpm2M/c5h19DLfM/2HyJlGDFLINdYRW06wJbqxZ7BSouRaBhB0
rC6qI4+/oTMrY913TEzvCqvlPrRLq8RTlxl6W3tnOMhcsGpOvYsSA3uOi/Tabt/obWw82xuzPAV1
DX0Jxj/+DUs65RFBAwJUnW9tWt/WrAnaAc9nJh2T6DNkqcjRkurMlPYmKWssjnpEol/oHHnV1LqS
Wyxmnp7GxluMVCQf+Mwo4sfAXkvyGEAkF1wtNJemFXiAkIXZSNjOKP87ob+MKFkorvO+dYprqExs
7UK9QdeK1/TQZV0i3aZcIyCDCb/ukre0i70XYAyQ5yPQFu6qTmEKCcmAxcpIyYp6dnp91aAoYMvp
X+aF+CN8S2ejLwAQROVa+BorVR+cQyxlYv+kEeVLM0tlkxuf9xTyYIfCMA/1Bz46JR/2GRslwtPR
KEpY2v7+JOyy9bawnJBQ+W2ecsqf0vI1dS1Yx0ik3RNNfKKvfI/VTY+pXlsu8ZdbNmO2+amOjsB2
1QORIqjMZF/9jRYgDSod8PsrUZj/SjKW8iKzDpwcxkB5V+reamYqhQ+CrNHuDJ6bGGtAv8DHz/qR
eCgHtu/6W+U0qVrBkYVT9k+JqYT75uScoHKwXCSxQiihIlKskEQ5hEnNsVcnVrFqjVROi36WRH7C
y3HAhbGdnFr0rEgVfNEN//Gy1mJqiIQ3x1A5B65xqwaHY2ZaaHFEY3AEQlxT4SEBf/CvfqnZFj5+
6sXb6GZ91Fy+CLvOqK12D34qQYbm+EklTSEhBRrdl4JsMjXsYpZBC+hYDuIjhJrO+9WXms5LGB0/
r8jDrtdrS0NauaF01VGlRjA5tHlkhS+toB6l5mLLq5VH0ZXqvetKvvP7E5YQ8F3Ey7xJA6Z1RGfX
ZwXHiQrzo6YIpq58QceDBWELysub6D1WvqXhQWrtcE1bhghvVfdqoQJd+PjN8zlEtBUZ6epPUeVS
yF/lZHWWTAEDaTOpjFbntZ0VLLgvStj2Sz1Gi7W2e4eBecDY7JVfQ7UUOZhaIPU5BasuCVKbdjEX
ua2sZrXDqZ8fdvY7ovT2KGTOtXhyC+fFWA4j8uPGzK2PXswPvOc9faoPMZCf6PjKbuhdH6r+KLyM
dfSorNds6nCb8O49hxOAxOa+mIGdEeSq/5Zbv1X57zEbel4/Nbr1FSmEp0u9X/4L+/qCC353H89Z
Qi+STGu5pocrqNT5vHw5DAEsprlis09sj8VFJ4Bk3ZkaOQyKZvJ1tVOjYvLNO289T4v9AjHzK4dD
e1jaWBKHNB0EqLY1RIO4gUnp4wGSbqRi4UiICjNGUV9he7Uy8gWQzqNExSt9kOWDDjmZnBzJfFn5
HYJ6OEAlv3ZI3hBrO33gPqd10UzMmTqPEaS2Mi1ERbfOTlIa8zlpKE+zdxJ5tYfC9/0EjmqcCq5l
FTfJjE79Hyi5wF4QZVFNwN+/rjWahDBhtAGS2IrkZmFVcVxGu4dtF3AZg/d2Y0eyPcHpYafL5dV/
RiFDWfYxNHin2dWs42amX0J8/xxrfMifhzOlX6O83wjMPdzKCtBw/9JGCUZuEZZPuZPMd1Fn+Syw
S+iKzCdCA24IIYOrbYLIQYtgbvi412s7+DLyLRT6yk6nhLsSwXFAKuDYp2wgHTM1xSVnkF+BQxxC
h7PiMiu3F9BzY+4Qlmbaj8PG3AlFKJUdx7G8SFqwWYIkmx4g3GHTkT50XcrjhdCZn4pMEr6guARV
4a4piideP18zJwp7WIW5xuNiwNT1HbuzimvqAAeuH4ViZLbh395Uhbo/3qiuaZpwT7WYWO1uEBF2
3YtJ3sj65gtyLrZx6KmiEyUpbiKtN/nhZ+dAqXPUzXXhV7hZP3/s7bYvu8SkLYN69MOVOdzeihfV
QNjbxyKjhlX7YTGrhuUss3P2hMLFcVsCjBR1prkmxfyc5u6+OmpfdJmktpGWcJjgM2I6dcQxhTzP
8Jw5YXkzJpRBAeXIuztAcfkJ0Cx5sgDvqe9J1QB5YYkOaK0RrMbKfP5VCLqt6spnac7IWJYF7Tbf
kMrrJ7x3tHL7bIfj1/V5XxJmzEc93Hmg+YyQUZnc04+NX+gtlhb0toxgs73QgP3PJHXp9JRMs4M/
EPvJaevGe3A5JwviLp12Mm/eMWtRkcS25cCPOkFCo3KuSQkWL/Ht/jJZA6eUhumswW7XOjutQ+xe
5hQd1d3UkwuDeIrFiEYsvcyIBmjSgtktDFSXPCGpDoo43vtM1wyqRiXw2r71qpH1d5QkfE3uoZe2
mCZ7BUd3m9vX90i89BxEiJRrvvRP9DhAfirIycuoWyIaW+7ryetJwIX+jnvIEOAUNZ29TgOcPL+h
lWlQtXRDqUzJbz+6aCVd+a++kZZ4t/mYKEK9lKYbO0oVWuM3ECxrxmr7KyX9x3wWZ5iCx2/+YPPm
2OZEWwqoAdiKe7t/cRTQjKBGtgjWSQvqj3p28byKq27asP0ISAuqOPGN9UmTDNcWE71DC9YDxe88
LbpX5us/quOkA1htKmZTzG4hoVduFD7FZUKCO+2jfyxh5NEtqRN4YgDAEYwWHdnO9UCVBSGm6ZEO
gilvzBqX5Mb9Iz4J9TP0DYY5FrJ5F5aIRb+Z44+MrxooGpVyvrgVJOlOwkt242RtSfOt7Y5K5lSE
utlIUua8l7fTCgYBjJenRfqRRcSceQIH2KrQutZbFtbKmrnUl046mHP+cO4kDHWIkkIOJ5BIgc0x
VNaJHth95GSBXwAMi7Sfu3JJRRwPcF9UCX5HzU54Sr4kTU64hujMVVW4v6ZBeCn49GPl9bWil3Su
F43NZH1VCaLfX07+uki5IiKHGgg7NB7bQ62b7Ju2ThLFfow0Vimbmsc8C2FTt8Y6sHlI8MX2j9CO
8HJgOjB+g4uWnW4QCzZTMW9tyl6tmw9o15oR5jblp8PUG830yxEzjTOWydhQ/TDX5WLBkVCqI8H2
+NwK2xJudXpQ61mO6ZbNDUolicUoFtaKR4Wxh++1utj7JEJwBGniJiA+XVEse8lGWWuunDISWWQJ
BlXRHeGi+GCnPFrmNkKkagaX3KzF9JbsXoPUrLTpMkxCeXLfwtOjOOuN1MnhPiSLIqMItT2aTBIj
ytAqcnl4Iuy5+PSvfkS2LP3wRgCrhIWSrwuy1By8lS1jjnw6COrtd87iK5Goa5bOf9oJ/AcUBKoN
e2gAQQYoS3lik2+Qqky7HM6ay22ELhw+N4E6DkYmG8vpsNVc84Ga2mLJ6OWS062Bdv+QPVJtaPZL
idcEydhCZvPhROnvFsz3KySzrJPXHS2oR0Wvx7OT7VNCEGBUTC8oDbwHiMfvm3dAR7Jz3tesMICy
t+8grMrjSLhUyhxlbN4iGH9FNx7SUFrhNB/ZjdYzgeMQskhlW5Bs0gffxMwmJjQR1xzols+C43VW
Kq2b/hYiU2P0DXCoavTVVrE2IwPgLHO9iE1ro1lFRCiRti5JFOgD+Q+iCgTe5BPZ9IOQsDXlfIZQ
gfoWUz2XzWEDnzrWQN/mvvPii6lYWfb8d2bWeNIR/KUfB/FODs77u+ARdBqrmV+QQgyNvCBvlL2+
cMIJqXsbe13t57nQqxywowAqmI4U++Iu0QqtR5iHwie9PIS4ExI1rHJFjbCq6qHL5gllLwYAWgXo
3PL1gAq3b2DBIE637v0BgSTb8F2HGeKCt2Cu3G+OYPYGfz/MdgeJaeGXzD0Dpy46uG7/7zwMrkDw
xILIypljzRG88XiItBUYtIQUIXaZBtD9Bjqubmasz9gJ28W216Irn6JAXavXx5REjTxWQzrWyXyl
16YUHEhxVOXf3osZw3sbq6NfVK3/r8cdnNSUFyfhWfZWJvcnW/NP+mm0EnwvGvaY/eoeomNXfQTj
bG2LfKN126u18b6XH43J6EYc8U2yZEP+R62o4QcuxtFoB6DDYdYhIqUFnReCL/cKaFamTAac5PRv
W55c8YM7of0n7l9ELORs3EC8+3wapCU8PIt49qw6POR8bRL/OsRnTk1GabDw8xtEOdzpMGZjSRSn
LiBqkgFxEElpA6DvsvcwHISrorx8SDnghnkGdr3Lui1HS6XzEQBTu9uMYKHjCcFgPJxL498VhLRO
1AZv6zv6qP4O7Js3Nn/99QoZnuu5GUQJz+so77kS5ETLHQNDMfECV+RtoHznrgGKHsvSbfpw8jqZ
JqnO00+XIruZsTdp8aDUNXoewEBR68wY/RFtD77TyP4VJkLw5O4M4G6rDTsqvhdiYgOsywaKnaXZ
BrICvkfrZXYTe/l3aS9/T/zF+btRAS3PmkSDyZA4EoYzGNVfKOoKpSe1TqPpIMn/bFNJxnY7W5gE
j/VBv+ZTm0WERudNd1UxnloQ45vwLzanbKt8C44gTbwdTVFYyXc4sYq1Rh5I1TjLRNFmX51MKXoW
0AX3XyFmD1uN5EMu5cIuznlL/C0fYULxFj6qEixBMhXbuUW6N9Cj3AWoASZU/FombR57n1vOAbou
I1voZRWJw6BmiaBYjGqidKPeE8cJvT9qROibuEfD35x51WpnMIBFInq2cOIzl4Z+jUKhahRrtGUE
Ikq+CkBMj/FYKutJoQlhHFffIAw4WomVy54PGhuBJ31njE3xnHGo50DbWjpvdU6RFcxWU59HbUm2
yRUcG5z7toxDvstj1njC5G+xSs2aYskGdhO4z2FFPYSbMBiz0GMOCgEdVE7+ggAsORTE4xhLEfYW
veUfYTCMCcuLM5f37BDMyZ9WtmUKQYae3ahB4FPUomH0XNDPsKU9VyOFVrT4ZjuojYe5b+Bo7H7i
SZ6eGYtjVGBqdOPhJqlDKl15xjxElxRk849AqUCDR3OO5aPWk0PmlKai+L9wOV/jnyOR58ETlcGr
FBE88bomsz4qa6CcW7zla/TZWCtddvEcWvUKnDouIhkpNebIMSgInJ5FIsRHBHXk+ylZHi7Lq4J5
4RmZfAqLQnR/wtQXOEoIrAAbj5BniFOtjtx408ckMa6gq9VRBaPIJPmEEr9H7tbmS9kKZ4A8gcG/
qxTBnKoJ7MGKAm+/V+Jp24akv8aQ0KF2SXJ3AD+0J+laiXmPpZ5eaFujBzKomTZGSoCKdmE32NFf
baZv6HNRXULFu9ONNyOV+3DhzUsNzCnH8CII6ktVtKWCZbWYps5irBHY1aBv1aXr3/ek8Dd5oW4l
Tl3lfJKyEdu/O5wup3PbJmthSIfRE0rPnDP00Mqy7TjtEiddlNqX5wSHac/d27MJdpghC5tBkPwR
KrvMaeQyxyinD6OrDBaqPjmEtbL65mopZxnfCmE2mDID2seP6E3ojSYdIl8iW/PLyQuMV01Xrkfv
z5pE6dPgfO7xi7mj7AQJo1pteVOwYn6hXOXwrRz/FHjzrTfrQqZcuxW4ilMVJcNWFbQH1j05h9o5
9fiQ+t28V9iBnllTgGRtnYGjCkj49lboP7qRmWqCyCyPYP323iIvgrL355JQQlCDKSIisGEShKlp
YvQ0DpwkSVpIU13tP/hRY5DDN6i8hfmTyxqIJQU3rDgGVDRRAqUhyxxMzDmBA/oWAjPfAkSnkPOB
TmFf4QCfguQ/pj3XMS+ptn9k5P8TT8PSfVpLS89lNoKhi6Ge1uRis3Y6cC3pQ7kOQjd8u4Ka2fIl
opq+5b9QvCDIMbRy4tAXU+0WJelP/F3ktPuW0vY/GbnsceaBZ29IYLqUgFThC4On3UPtYYshx5cd
PByGPnaLW7b3mrkPm6PKKINeeh0SVL3IUZKFQADNKrFDF55j3oiEV6lNOHEmSO32tTqyBiwi3Mr+
xGSQ3wS44uDiFxfUXbupP+gj1Bq/VvX8xT+FUVTO9XEnjQns9AjRvA/7ofnnTck9Q8Uw2pm8O8DC
ndbxDMsK5sECjxmGaPQQPPKjMsg7Zd2NU/uHf4u7R2gi3XtVnVtLCU/iVw4cx7BXfkPo/MT3p/MX
xXN4OdC6d20qeVuOxlgXN90FWKKnv7fPWdScPg4UlyblVKvvx6W0HfSMNLG2xlLUFkYoknGGKabr
iA0K5ASIMSSlmewyitWm5nDWZCoYzKj0S+vez9iMP4DNhlQ1Wl32ev07DSjpd72Xb1sZXHr4xjyg
LrSLnsHzmlF/HXPe11GvZ874lcDJCSPhWacUsMe5OeRG5UNgYyXnqUxgEtevhkZHIFE5QAZaqRAp
znV2cBXwNm6+4Tc47lY5RQEGTQ4iGBKjb4JT1dDov8e1W+ngkLHGWD6EgiQuyJTR2oFhzoexIGG7
sN4LZ3cLE/vMz5/3k0aS+2M3T7LsHoO56A4FKEHRPkiLAiO6o86OQw38Xvu2Qv1ni5y0fFQ77lX/
NXcTGbhQ9d2G7ErP8B5Mx6hjSWB2kMOCOoUQv8vegd1phXggJKSlly35YfORJF2w5/WpYQfKH9Ml
XG/aEq0v3qIssODyO70e/0o5fXPqwI1vaQJ0uWp//Bro7HymAOIYCP2kOh9o2M7gk6t15PsivQzO
v1IWCm/jiQkir+coZkJMocvMYbDp1IWtPoX64i/i04JZpAno6WJ6xKTFSdFYMFW9A9jf8PFgjOll
NY5g50kt/0C47lLIfepeOM5QQtpDz/G8TamGM3v1uND2O7pjS1uI7U/FFBT8p/lzWeH36P1bL8T9
oNc9nk/qY34PuAFsNOgqhMzzJj67YFMjYy/6sVms3cORMztE4ifAmYZGjuwgkCnDPcRc7q0Qvrmk
3IvNxMWcntszyZXNdu8s3bFtW1wOey0zNiENuvwf2LYMwNf0tqh75oi97D9pQUJwC8/8JPHiChQn
4U2nzpfo1J0xp8HYrcO3KWg4pDpWIJggfm0usPn4iapJX68i9UBVge/AlenGbW0SZVYhQjIGuvPI
k31Q0dGAXJFE0Gi+WiyRxqubxvTnSsSB242SKxMx01S4ss0jLfelvb295lS5nT1+ZtTeYaUB57dQ
S3HkM+qcFLZbhkX/t7pZ1OwTF66hInNTL2li3oU/O5BRNfArsViZQWvYfyX2kaaPsu8sd9UIPgii
LhoKYrJRjj65PHy45IHdDzPYY2Qyxjgm+GR8uyef5lVAJk5s8oTVHXd2VgV3N7XV1gx3QLp5J0UG
Hqxa7syBsBwnRONjaulmc8q02+VTTYmoKdh9pn7GHktuQHtBoIsY4YWRMjMoRmf2R1JhiAUhMmEs
gClnkEgI2TXS5S00aD8gvnKMcT7u3bSKqToOriyi+DwpmSSoFj4fLF/k4GL7nmg9YPM0O0q4OzRr
JY70Y0mH971FFElvCtZkDsrRUMCR7TG8lVr6+6oP8BYyH6tEknMiQFmKQ2YfQVqyDJKHmy4eKrG5
nuay0orsdHgO/rEMmm+p71J/239KeGau8wq8ELgQcJ0irZRr5IRfum+urpdMl7IQy9/0laY2qzWe
8Modq0RitHNOkBrenyVycxtQUy9WNTV4Lg359Ivp6/CWvd70qkZEkTzcEqfl65U/3xLMNItTRCI+
qQ3k/TIBDiqVSGKKyKiYezP64frgXmHKgB/aoorxmgXvjJplENXq9pSoUQedGRtuWw+uYItOsmLC
og3p6n68xF0bg6ygchkgAYy79w64CJDAsyqD1jO+HBi6b4eSsm82wA42goLtnlwrH1tl1NekFHvl
ipoDqaK3rHdkI91Hj2YO4DjF6j+cKjkXiegK8o10XLm0bU9380d3gQ7yb55uNkT3X/kA/buWD+/s
+NmOYX/wnu4Zfz3LiRcl+cDbcWeUkDyu1ShH05nMravaTP6wVZTNLo3dNXp5cNfjwV7+PiK1LeZE
iptkenKgS3tD7tywDxWzMR1q7NSwbnRf6M1FsO3qxmk0mO/VbAc1zYcmChhjGndSlEWxWrf9PHbl
Mv9DSTv4+S7yQfMv3QphPn5Hg/RZ/i/JHdvwpmbBt9r4CCQHwS5G1seoFg+ExmWDTcywgyJWS5S9
Ms2Oj3mLPWhzUOgg/HPMONQf32Q0G5a1fg/B5smvYEXwO9hvUSXX2UuzJlto3IqnVutbPe4IVIlH
O+pQI6hUA4vyFsfy+1hMAatLB3kAPzASaQcVyy+WwP9jYAoOIi8MPpD6sO7MrAutSlnWrUtgdFzp
XUKMXV0pKZN3s/TpqfaA8EeBidm8IK0xfGSlmjWApo9Pst9tpKymdurw7nsIooMcoYxhZnnGbiU8
kSk2tCUAiP/GDxGitFgUjnvn6hH2JyTfGkzUcpJINALohnFXuT4yT2aHwbRiMLTLGlhAvgMn0VrU
rSSNBjdQhJReNPRn3Wjp7ITRiTkWp56B03mIQgeHYNkz7E+2RS2F0UduuRmcPuBYfq0sveJpZu9R
aKca3kv9/KmqLOhhDbcJYvl/aW9wcyNzN+d1YJM6MurDQPv33P+ZzX7sWabh1M5wNPhl1TJlUHHJ
qdXhnZ0UvEdLCtwzw4M2lukK8/hz6U1PH2bKRnToiEwf+oWS4OP9sKkEmNE+z9V9Z5HUxkzCx7wm
Fq6qq06CjsULu7TlhHpgi9Z3/oaAm8q/XDWLwF1s6tXKkNgLWtUBa2xc/Q7LfYNrYB+MCeqbxHBY
d7FD3+3uG7aLiHFUKgTiAxiqm6NgGvymVhUf6inV+6VC1OzeRHbv7TuIMgWcFpJLR5Wdj7retCr4
9uUP0+7OQrEO6XlHskAfJjBiFikXqgm2QZTxRheeYEjkZm5R5XJdyUYdjoFnqxATb1a9OMjAI00n
nV+8Gn2/gGY8AIU53G4o7RGEHw17CfQ0oYPsN4aLXm3GuNAGliU5d33IhJN+QHGKr9L8+YjSxLe1
td1BfUoWjs67MEQacmUsrvNq6NIc4mwKKGLT/ZswZYKZtQpnbpyXq4NktQuEKs5fqI1CE9yOEHv6
zpmd6GTXpklw7kV7zAHnqofMGO25VgzH1egyg/98Qw3VqeWI6wbVQWXQYJYu9ATFTaYzYSV0pP1F
3HRz9idhpR0gxHPUDxhUE5VXWWZ3yN/8rdy8CX13bllFMuw9O97ULPzBqaIn7MrXvrbBkst1LSeu
kzN6zaKP3E7x+/B1BEMUJEpaJ4y8XANeDFyjaCeBYBs+SJi+4UtPQpgfTT0mRuTyRaQUtlRMjOgO
EMSRvUyLsPNKJAPuTneLmQ3FZfbopgvLhUWjiEyoK4SFEFVEHqIfHE6wk399Ohlyf1VcMn/9f/zF
xAO5TVUkQQQ8ebTwujazpsH2gdJI1pOm4kGIrTlZxdyE3KtyvCzrCMq/bH9VcbIMSUcb0h/wr3g5
0GChLu75StkhFClFWQXES/KvuOhE6aSJCUqsA8TFoV72u6RkFDiqSw/Gdn38CtpoR+SUgrQl+5Xv
dZMCMl9AuyDx8kdhSVj5GR0543hJtwSqpb7HIx/VfeALfN54crpk8x15iIfD0HfbUPeh5NWq4tw0
nxUFTKEGPg0pIbg1sauwodYymPefnuBs4s2F3llyI4hXbUKbLgpoR+4+X7XxYQkQFA5sMt45336r
a/LP7lI1y+EOY431kEuudgYytQTACiwG0I85eUfgaj8tR+G5ugesene2AejOqJKRsAYe72Frj74m
s7SgyI4LgdRvJl5V0qBumA2DpcHVo9hGsnWzl56gcFyR7CMqDfGMSzMuH9i0Th949EEzXgkdq7jO
vW3S0VTXkpqR6QXPXkJeoTnmBDSzKQqwTxwKViOYlHEw3Jx1aC38ninTEQpYUDRX5Mcvskxaq5hP
xj1lKSnXnt6vIuXuBNdnHBHJw49iG41go1CH/L+VO+ltOO6ZeIyGXg/wiGBhFAxM7aZvKeNe9z6S
zDs2alSuwYZ4he0x0YDIFH298MHfO7d9cOy3EpPLH0ARs2He4yq7/TLLZKnwcRtgOy/QsC+UMM67
eiiQCYNGi1xPpNm+jZRUCenN15IW7BN9c/X3sty03OjN+YMMWkA1qECoeq3bUftEn96ByTzg8w9z
rTfBR4uK4jwcpn75pup2ogmIB6+cSPeByIyXoJXFVbk5pddxOgPPOysToJZONWKyE/ET0tZsgJLY
WbiilxjrM+UQYbWdjcXQ2lNnNhINtCWWVlcYfrsNbF/xzvvJHooFfjFZEigDITa0b05MC4HoOdPZ
qw9XRcjfvk0xY1tWPQ5PZatX7IMzBsbq44MZGOmQTyBeqLiWv8eNbSVgysRId9/5r7uMcb6nnkZ4
FiMyiBICBvLxPa9CW/+Px4rxs/iPFrYVqRTiKXAFLq2UP1VhXDuY1/eZrZAke97NVcY37/N5YNcS
kwaPxjgqlJKzttmui2/bbtyc1V4JBXgnzSTN+ebmof+SE1MQ45MlMmy4BBTeaT4wLI/QYb0Lg3dJ
J1HIQBN4Il2bEMaUXwCbTwRk1g381evwUUQjvZiW9WkXu3YKIUNTtVyaX0DooJK6a2ERM5SLk2ON
ov00yFBu7D/wsmEKswcXELl38VbVsqvT2Bl0igSspCQVkY0WXd9x/lf/KVidkkKA1HF1YFQWrz9o
+yvpXDF7OruAalgehZg0K/N3NpyGd//F8aiFvo0EsM+PJ4OeO4gW3wMSYVnlimSVPvC8w/8Iledp
uZXesLVC8j0+aOHOz3s+Tiue34f2jtlhTTW1lbkdZW7fnZ3+HF4EboBUzilctZ2qe23DqPngeIOj
91ILZqtSyadGjYq7pRHsi+hjvvrewjQdjzayC2viqhm9/HJqKqVko70gHSJGW5PcLSpPtlqwO60t
5AwdlZvgmPlOxWIUcOL7vcBnK+OvzRq4oejmXy0x6f43Dun7x5Wsj4gBGA7TYAvkFgvieZtLo/WB
x+9gMBsyaQkzDJ/0WfKk14pjHEijE0B1MnQyGF/CoAVuv6y/eY7rkyxQHNBPVYRePbth0RpM5IuV
fADOrWz/0aOLyY6XlUNyFhZ1DSDRDBVKwebWpHlsnl+drxqucS83whyuTidBRf9KMthNFSFb/Y5h
5eHM9g3nEZKDg8wVvpSFP/oFmo9TxfQjIvm3ebuyiFpw31WALodBH/lPAEX8pRhRULnUkCLKfddJ
vRJnX2AUWobAAPbcUNHFbZrql+JlFvywNbaWI44jNxf9X4fTzEQZt0gfviNCiMnF86XmaGrbVCcd
EH+BNLOwkbnsD0D58BWsgPKWSUZHZFIPu08lyo0/u/mUhIqjCpqZPDNnGCKtljnAsES0ks0KjN6T
MUyRvbTw6NW7YIXp3xAe5VnCQP9WAr3QD53ZnLxfmZddTk9XbHOMW6IqHX/YolbNmbp3uekWuHlW
HZ3Z6otMpTQwTm4O6DQeEAD6+36kf8HXyDOEa0baIaIDrmdwI4lNzYZ+UX2ZMXkJ+DJxlvHRLkyf
aOAnxMlE70nuzA/+nelVF9xd2pmhc8unqGCsouqjhLSdIL5i8oCLcghvMWKl2MhMVhcKQc8n/GKc
TqMGHfq0rL8+uSADMFpWJUzy21yPgfcOfBGfc42eXFI1Pi0NNl0oR1nQ2kGs+I+JyBm+onK6LWj0
hL6/xmTk6XSmiHN53kbr40VyeRt6AMrT8SNVg18Gb5bxB0AEJBxr1pPo8TjOVz0K8B/7FiTuDJC4
V7TCCjRN8L3BPkt3a1C74yPSTPcQ11C8liUmvc/wjo/7UovQrwSjvGgnSdlhrEgwoKvRXrA9SfLO
048JsCSzz32Ls+50M7ZFqeRwpCxpUphrOyxSJx26au61UzPFLNwCNHnP8vFsFfCFCB2uLnrj6oid
R+yHfUfkCOohr7z/iqWG3N9itCmokCwxJEzfA46NT7jZCCPwvSyJhmK3s2gMO6SOf81zXQkN3kC2
KLkzIlH1zti/qlRuX7XQvRj4u+qlOllAsSVVvHC+7rV9YJHAhL5HULj8bfzHxhA87KwHtK7B6FLv
KiO+Xog+06AhhYgKVTw3Vcnw98PnLzQlge9iqv93EkbQGVLRAj24L68vmTUWbCl3wQFyuZ/MEFtx
Ti0slOiEdsL+KZbCVWve2VktICiAw97BvB142MRIaIoMVOGD1WlnNPxCGuojX4tu0qI16rtLDtWC
cclpKkBYAqkoL+6VvNV/wrP0k3HY2hODWk2iJ8bqy/qW1Dgd4VlSAzEWzFEL8rwzDSOEKTfNMXSe
7lsmJ7sOpPhR7dBNRu8bXxLGri9BNjUhpkkKQWaI5BJh/XNPfWGUzrOjqVmo7MsCWb00burTm8pJ
Pd8WY0KDfEhLgFMZpjbqvv1H+SXrDAWNGAkr35RsV91GGTIy3HKIDqnyDyLIHKPBJkiks3KxttVe
8vZHai4LG0FSbV+ZKGo30UXTiY5YhgQ9F2k0iteqHN9P0OsLyxopZRWqJxdR5T2qufB1rCLYDfXg
C+BYFr/v4ZdRuaeCM/sINBZzVwMx9ZEOq+ZxLelkEPhhcvfgc5VrHhJA5Sq7QUxUFZHmHL5JRkIM
2OnQ4FlvHB2Cqu2mJOUkhfaqr9ahxwdapkzCC9b0UqRmmCfeZfVPoBDpSNKMeXMAdaLajmilFTzh
hjXqonEy1odqvElnxx13DIuLbrTyMJC60YF7/1WNQbtfxLWM48y/d7huPFTEVa7Jd3JWcXGErCHt
RN9aYr+Of6ZoU9xGW9WOY7LHM8ZZFJwjWWK+1RLWfAI24x5LPdFGME/9OUJr1F4yWbC3gKRKOGqE
1yju5K0/3qqvnHIuaJQssEuvNLoyGmKuGTMlqw2B2ECJ3pGT8X0t0Pi8R2NPM4Vi0fb9HnxQ/1KF
3kC7FZ506zDU21gQ0tWL6s4fCqzrZUS01jh8BBMDwYlEvGyIYeFq2Fk6i473IIarT18Kr+xi4GBJ
0Nt5rvAlj6U/I7OcllFrcditt890Jpirk6WMy0Ss8cZNJ2/rOTnSTMVyoor+q5VBgd1pieRD0/IT
VgryOAPWlOMkvJ2abdtzxZo7fQ6sWE4i9J8UtAWvH376a0++dzPFQUF+wjA7yPdc72tFAdFYEAcT
k0reQPaJFFC6PkYHLUM+dnUKni7vTUn4uSTN8u6FMH1Q4XUJ2nJZUMasdfs2534+3mZTi9AJGJZe
yr2aGw5+Z1+NqyH+oIfdNIyPRjNlsaih/GLS8tLdKJAqW4r93UspL0D9qB4HLYZb8VqeKOqx7zMw
t0W9UEspBouXkOWfb+uux9H9mo//a4Zx1wj9k/HJl35WNPowBSbNS3POYtE8p56QuhNmUKYZWoRd
rfiiQCJDG6Y1Ed2feaT0x1hJ7tiNu+p0peWlguBDmezjmDZ+BQdp71+4PBsN2EaTB0lEC3H3CyDT
aTAqbNSqhQ7ON55viy/uIEO34ssC4lzZVsrwGbGHxNLvT5Xn1GgnkYtk145StexWrah9WNQq2Y9d
pbeTv5ZGdf3cHW2jDD9Sg6tttCdkTbiUFZqtfMqLnaqnC3k3clnGOspCp9kWrErU8mYj7pVb7eC8
EBrUsEO5DbuAjF4+F8ixKSjCn2X/rbkQhW8Ee/9rzJqyHebSKQh/Behr5a7Ve0gKdsaPAtb6jXDX
XyVsuvS+Rjnb22GdIrunb0tdMqbHcPBtSha5pCjWqvZUTNhs2DxIE9H4MDUrMT3cmDYgma9xowRe
UdSLPmsvEOCiWVKjV9wZXQZHt9hA4jR+xVnWe0zphSKjGuI50fanoZ01xbls9Lz21lcHtDgiE3W0
e6lTww1yKUAEdZ83HkptI+l3asL48EHGe2+7C8l4Quj9gfp4/GnB3fn8Xt6dwErORtd1VRdhedmx
EbBjRvKVeSxKLnxfTi2iaamjrysPLMNZW2kmyvOMk5y3rzrlEqlrGkYyFJy17NMYIwSfo1QF8AIp
ivjv4nnSkV6QkzWbWKVi89XywJFySY8FknvM5VHlXIRRiPUFW9+tb5LfVfTb/vGfLmw1523RF+81
IEcMsyCTWYwSYtMqMuRAI7IFKI2HxzaI9oFTfsRM+vaWn2ZmyF2pYzvcYz7/tHvkiAEZGcJ4HGCA
qLvsKK1pg0gMfXBYdOwOJo6WrAlGYa8mi9pZ0jQpkv38qPInIW6xMRIZnl9GVgk/JEBxy+Oh1yqm
CMTrM7DT/vLbOy39v5oVgG7KNmV4GjIKxQ4DWtPaQ5M6RWMpDmbJyC4H0rG++QJlsOH4HtoEo3XE
bDq+vWZkXt4BiMb/MhANx6ucR8G8lcsA6im15OCF8Uekur0Poxc/4uay41zbs5g0lBqHo94SBCt2
/11p238q0PojuVDa8CNeUgd/aqDLzkMjAJ4/5bT3QIsGpaiiEwc5DmRwbhKweRHGVwssuGe6EEQT
3zetYro5T4z/S04MVOYmsVGxb+8k+u90Qbu4jVF3iHGm2SpiMOba8ZQmGZcWtHj1T93F2o3fgJay
JyDirbBaU+5YJXmjrhcJAjNVFolVpltNEApu+L02aqpvY0YLWsVBkDLQTSyEKL8EY3TGLNlTwhoi
W0llb776saALX+PUTKxXspEeQIobrMYosXxFr9SQr0ZAC//MCpm7WdHLd7SNa6fm92naGJyv3yZh
ShnOo4Bv2HxK4mjl0GCXK9mdKqt2kR2s8OCbgTI4+UELl3L35Hzc12gYcYFncHG4qBdnTdHoOg9s
yipj5dWyqJ2EjeJ6jgP3LzOxFAWWBVj+X6Eja/APQPvIaP1mKDdjy5wojeVBhETqC1JPBRBRrHuZ
fhw48zozDrfmAm7MKzepac1GVYzQxU/jefUsgeAiqg8MhKGorf+XXwPaFifTSP6nHnZi4VEfBB9P
GBHBDPUATRIwl9/ypRQD7aN9wAJxXFkwyjSxYvVjTpgBS8dlQmRJjgu6T1SbxUHwWBIvA1p/kBZa
qh23sx6bSWSvWbZNTiiPJKu63Wx2ax96+Eft4Qh91nBiffcSYGEgIjSTelHIW0LCYv3JFKDdRDmk
2pxpBonbpxu4Q7P6gN1Y1tyT1LscO1mSa8UP5uHmwmWd8XSoMyTsWfSriIeYN0z6pi8KAIsYlNiL
fH1bh8G1EM1P+qjHyy+egnZ/7MR+bpByNj3eWpi7pd7aXUg3jWuH+griM/TRT3+jONfv17rRdACj
52ywaRXi9uLvydUUpDE929gGbRWlcJnWC7XIv1oGtGm+pZfWwjy1nglBViYvH2ccFcFuMfr5jptO
EAHJ29308qv/ivkC3/ED3Es/nFEn45hEc3LzJf1WyL/ob4HWXBaZceLDucoeyUlRhksqUATD5Axj
55b73TQb1umLjpKESWRP8DMIfRGi+OqrHeYFSIzBCOYHnt8SVXdGVwXPUtJm7REHr37a/q/LiFY3
gn/+xmQYDSu6g6pZW2pIBTelinZQcjre2kw9LE1qT1F8QW1b3fZOdfnJP8F+BYmyhMW+kt6st/Wr
5jOA8XwFNGtoIrNk6FRbpMVDiizC2b5+h2iJ0Q6LWBLahcZZLmwdJKu4HoUzpjvx47cP71fpUxim
aEeJpBE6zHbN0qPc8U7JFPLG6c68klDazWwl6cqtA7Qtz4wHrB89thDttYOSMT7rMd2gD6zNzGSt
lPjj1nWJR1dH9Tn4bCQ8I0k2QM138aIZmk76M2esxDs/lPfoCy0ccqbQ3oyiDppz+HPT9csd7Bgm
QYehbX+Pwxl6W4X2NsjuVMhvXZWaQ1wTGAwHLM9l+UnxXd2EA9kVHh4R8zSw9lnMA27MvD8viuBL
TobQLfe3yjkHlve7559D2XmrrVhwoKOkYMskbn+IHduYNFxsTBsBykTruCmymDH+2nTXv+JVSPN0
9BO1yokN4Jq9xvB8dOeF+tGm+Xk5KeslFh/07LjT1p9u765XBPL+fpe+IpDOCME1BH6NtfykMWN+
fTnrRuV6oAzRgr7+VNZHQfUSBtzAlkY0TJ2N83mRoRh4ykcXWykso6o0TZbA+yrlodVPleetGx/N
HPCZ5WwWK7KpY5Hn2hkia4M4peQL+qY4fqvOX8fzt3oGh7z/0AnsoKJlwUhEWBv+P118obTz4C11
YuoAf8Wx9CGhxo1gZex91SN8h2ze5ZIvEaz385jgECXKfxfkpMooYMwuC4iMEGU70oTlYokds18A
Bh0BZ4lw/sJ7jBuK9FjcsNyhclfkhCbGPA2lrjNEYk3HGk65WVskxhpr6NroKxClgoxxoIgMq5Xp
oW0WeMwZaaZD2fK37H+MuP5tqblK3MQRT7lhvhyuZ4Nw4IYXnq+ZgnFLUesh19TwbjV3Ww6h4gdV
9Xk45kfctk03YwoQCCdEQE8HquI+jcZzIz5xzslm1p0oR1j6Up64RlLhwPxRtNyvRLcprEfwJnUU
ljG7HF4yIvYh3NCHqEAbu3IrUqU6DPqvsSrnWCWX82MrborooTDp2Jw61k1CBJo+V9lAO/6zEkhp
Sbgb9QaPg6xcU8aeTnw7j7CtaF0omVp/h6u5fliRMHxT67WavvkCJ4UJFtnEplMooHttsHCA7KaK
OuyjYGXYxcBFO5jN3tQS/hyKfNIVuRcm7Erk7sT95zfIMZHzxo13kkN1gr7bsw1GJOOZ2iJVEJIe
wX6SChuG3s/0fiqgkmbKFrP06U9iaZrLsMyFapWzUlcMU20VUgo9kfpop+bswM6cOSMRYY3HSsDv
OJ1x0rk9rc23+wIJ0EM6ONlzDFElC/+H96pz/Ju2lnGVMcdALj4bU4KxbogVvZtt7jZt/SUe+y0a
j2fN3kD97M29Xs/PnMdpmVOx7qmSwbFlgmrSAm5KAywla8/P1Uy5oyWO4Tk66zcSjJEMf2CCeEnp
YDX2E2Fh2HnRLTgxlBaqCujK14twyqRbnHWxTOaW5IHdzLAqKmsJR7KNHXeh4xpOSn7C49YKqZ7O
k/FUkMWaK5EMO1dzG3z88a1xHp6S4GzpiQGGYOFnzxWnbuefEDe39jN67VcGKy8+07X5qTtp8N6C
VVCzFfQf6J+wOXEge6Tgy3muk9v/ndnrsQEf7Q20NXgdtP0m/PoRbnnqtFhmQ/sQfENNmf4OuxFd
fMs6uCi1dlP2Inq0CroFNrKaSfcN+2258j8emAXp64tn74OrnbVN6VSb01nFW+lPNpO1yqOGTiF6
/o5gGd9+7HxIq5T4tqCqra6wNHWWGSPI/vzPNZ3JnJwZ5K1mRj7YJBDT6n1eWOdAxnKIjGdI9oWz
XlcJTWvaJGIgk51dNi4d23Jf2LTaOPzL0uue5CQlgSkDsOrnLnU87TSOmbcFVZXpZ8XV3X6PIfPm
SqAmhS951bWtJ/RgOB26iu8zut90QWoFdelzRGgK0nfrg0zg0JnNoVbxUWwnmbbbKqVqgv/9XzMr
lplI2kMjHjY9k1Ub3TKmn0nSufaUtNati9imTJubTpkLwBNEMaWOAYoVEcqGFNfAym2Ju3Foxa9g
eRI0j/HkMoYObnCROh/xXQRu2TeImKOpIkL90ZG9xyrMMosXEQBm/m1C20tq3tH6XPk77nZ3o4S8
VpOqEs17nH3I5r6TniecBVAyGWEsnghcS3PyqofH666lsvKhLqXABlf5kpwQtbyUxzBpAFKfa/Ia
9kMvfziRCrFuKxTwvqS3H4zu8juW1EE+D8VsOx0cQPNKgOAkTFkLneE7t2x/PHGjsQ7tFk8wNIh/
iAhbNF5umT07aSHWtN3MVJqgUpuOIFqVdot5In9+K0W/Kyb+tpocJ6dqo3PqIG7sIf+Z9h5a4BUc
KRkrMwrYrPPli5GVFBqn4KdXgayqN4wMo4Nr7cv/KTveDdriKQUx1NU5AGsvNd/rfHDuoR9OLl4U
QnIgQ+ArS4Iu92FTe3D76yIqbixZdfWo5vB7G9ODajaWZnoaXE59tVY4Jw5WLUwktpdfPRtXtGLK
Mbj/N65t8PnZweNPRJ7ChwDOkEyNHanlNAGeN0T5/hBtGlGaYUFnCrfljum9nXEbmeB/R5jKXNrL
diE472BhqyqW+N3qIkd8RWDf5uLd9rezxR8IQDSTFxg029PbwufroDxHprQecBdF9rZ3d1Cgn313
eJYbgN+wpPGmdSZwaMVBy8w2JOOhLYwIyVGahb8MLGjjXoR3UMYVy0kDVK6/6O+KUCAaxt4wx/PI
5henFl0JBGv1nFpllMnJvAp60+yfPEqpliQOulUY7FTaoJRbO6dXTuPj0+JY4cynZFlt3RNivKfY
f/teVPg7+R61VvYO50C8Blt3G0NR+vjFJdjw6gMWgNMXEsZbsQodzj+nqUS3IXnM8vV9RyWkubhG
/dy2i5QAED3tLEL2QRFyiNN0buddk3zvZ+lIIhWn5IQbU+Oyz5JBsMnbNTXKCRJBStPo6dBeIOOY
NYD52EHD81hRq5Qy5e5NGpbuLlQ3IoHEy5ziudSe204g/wp9pEUQvSWoaRdYG1WeJnWrKK3Iscj1
52Ye38Mfdw4QZpX+RYCuw2q3KSlAbE6zIjEDxZCUyxOffVudqMdmVRg1WWsCphOdS4WWK+Uv9n6v
pHnl+pr6s/4ZU0EMjwqwo13yBmqVKId+LB3bp7lB0FnZhrQJNTEyWXTfCUCkokuc5LeuCCPugY70
wsJTR007zGHD5yBH5MmdYUP+j82l/JxM4UJSPxhS/4ufLXhQO0+NMVA1P5/k25sypLmdd9ivg8km
+3wPNWZqwMal1RCFgZy5MDCgu4dhnjbf937mNg142Scte7S66ihR6RAFGoyVuaTErrST79tCoAx4
Z6bnXQ2+6e7QydYNRsLp7w2ziL3Wwv6UL0wiUGNCUAcyg+bQVFRZUFmeGqSo/dUgIpGUB0uIh0RN
iLsqL/x7KRIrphlKmBjiKmcZAdqcYn1yjhGviEmos2S9501yvXyIA35evW7Q1sywTkYFvYfbQaWb
akiD6g/TlL841rMsgnzpSV8mgBM1Xw7JJ7IToJSS64E92XI5HZYmAJHy4xgaun2y/3XNnzeA6ZVK
Kd+Vt/uMeeJKYuhMzxZZBCq4wSJI8DqIf12pTA8XCe+OLpjkuGUbW1N8Hhod4A/3UDNQoNIayMZy
8GnYq67nb/A+9R9Bpb0P5COMx428hIsZjZ8+11aLKNpe1AqybNkGeU0oUukuOKE5Ihhn17X4uqpG
4S/p4wyS5KRZtk4U7s4IAm728g9XlNnzALIs+SmSzijEaekUxiLU/3DRLYRwmGBgWchNUsQf768b
eZ1O74Eyj6C4Va+dy33PY3RPbS/Pb7dusq2WIliNih71J1EfNXvjvvd57zhH3SmC6b3YpA1+YZ+E
PiA+/C6oU020878Vk7iMHNFU3r/X33f6Go/1kC1Zz4vd5wE13flU5ad/LPoVGIwPN/C450+nZbO7
0Jtxpb86FY93EP4d+sQkrMiT7kSPvP0N8j3IT81Cv6nukhT32LayhGk3PPRQEPZomhLRNXe7TNMv
cxnQCe1qFrOC5HQVGTfzD3uDtiERdqw+LqR7Dkb7cF3Df2gt7FOvSZ2BusQuTNhf6mchLG5SpeH2
kQfj4P26icYnwKk4YJvefjBEsl+llrf7E8lsAB8Sc5rHrpBhAgnniF0aVW93kBF1+1CcnRBYwqA4
6tg1v2l1twwBhZzg6qt5UKYEPmnyGz4gSrI4ozfGuCVHjiCx87bXhhZhOjsLUFN+rc4ylShP8sUJ
x6h6zVQJ1KkkwG0EHiNWu3q6yY+H/01QAit5SGSL04jA1OMZ+jaHtdIyMW0dTETKDQRH81Nv6SAa
uW8WuzvEBTSnAjPgr4/d1o1icowQlGPJ9jACRv3RVOxONuo/fB6rlfCXYzQ2BF8bGlDTDcvTqgpb
SNGeVgLl9S91t8mp5Yf9BDfF4XTWbADj3WMeYuUNB4ehW1MAW5EtRdvgXoDHtSmTolBodAfkZkBs
RI09WWLVrsukGh24pywhZL3H8YeEXvZQgb9e3Kac0Vap05tO/2VbPKzLN3DRVDg845n3+zcswFpl
pmEINY5jcokB/6r46RrDrQXvNKwZNaWoe6b3N8CLga/l5L8bEs+NM3VyDsSFkmDhJBja2mrhSycY
ON8tkq4KA1djbmwJP05xJXfQhYDK8FFzTrVcsjZKuEbSJ6pu2MUUaDq6QsGny2k1sy9x4kGcr02r
gpdjqjzBztOjJ+n+O7DZKfznwNMGBPImrYweRwrFw1E7PwCdGPiwU1CHjzKh0Yiie1cNA2A8Oaz2
tXNd/vuY4MaLh6CgQWBshJO+xTb07l4ah3Q2V3QNWBufKuKdNZdJciYlBprixAcE/wDc6C2nG9K+
laOlWL5adUHWBgcKfvPWFYeJX/wXAast0OlEhdssx4BTeZDrv3KyjQ9PWOmqDhrHN4HXxQyKXVIC
JERJh+obd1Kge+hXgDZ38eVB++P4W7LBKKkBL0Es4vPX3yF2cnduSjM60e31ApEuBGBk3XYj1QU0
AfX6uMpMkkcqq9e5zV36PFm/f71IaeFPLdKYDAU+uyo+mUfBL4WYa9iawEYIPID/dpRqFlUWbgyO
sgpYTMSY8OqrELu0hims1aPC4VemhtPvD1n71sQS5+hloWhTIr/LGeRpFb48c1D6cuIhu/UAR9Dy
zNrT/9cUZbM0adw7eKG4Jz4MZrKBIARUa57LTd0r6+fBWFAGmIylsOp+VUoE4PhUJDGpFm2Sv96A
p1VTrNDfwFWnr/tGfZfwrLWy0XLDKWsJ30Sr0Md3c4BMUp6VrRbocj2NRsgQRBn7Wn2TX0zRW/3q
5wXonKmkMxhhItr8ralOdPyPWyNK/+DAnS1fxZl9Ma14q9vp4fnk6c5wHpMx4qDjKCkh6cQJHIr8
b7Rq+KnLV1ArR9IfPAzs5sDZwNc+HCgQK6fJoyZ1skGDdhE7x1lFBA0scVWVySYydXlwHaUFY6GE
lVZksOYSdmUrkXl43TFARilfNMsFuoUNxGjd7hvph5jfZ4klceKrnGzaPa/QCN87oIOFAT+Xduzo
LjqRKyeGcH0rKc/uARL4b1jFVCCKvFlypxIiwjJFDNlsIw1Be6ObYaNQtArjVX3O+NsCm+jUwjID
4pueLUoxVaufA3LN2RfGbqrjg3vURwZrJD+gw7laxmVUrJM7ZfD1Kchqp1iiJzXu3YrbNUPczMLc
fyBR/Zqb36cBNoeNikplYZSeLnC/2hVSL8Fqo0pH4I0k/UlIN089izaaUhnXp+NZCbDJtKSbcJvT
3MRr9IKY2k1/UGvPhWZjfHaRVdSgAcKE8zY0bVDuSFNpD2fesF0BbcihpHuPtuYR90wzYg2KgcXM
MHwtjpIhIiVnyuC1LAbbvmZoBsHO4fCKbR/fofsTikHexghwGgVqDeTXgFxLlMieW7k3caub9gnM
anwO2L1GVVzUGNR43ndfw+F65qW4sBnippAyG/1UGb772TEJfRpDC83/IzcS+0V9rVQj5mAy3llQ
9qU02cIIPE+hT4sjafHKxe03345HsVy0ajK096mOcHi3YeBq7teGbzZPjSq+qm36MJsmVmtIdAye
ntXXrlU/xNkDtgjkyBMtSE+Mx4BvQClJGUMr2oizy9sQ9Ocyd2BDDuPPfFVn88aZioNoeCpRxSH3
bOo8KvARTKqS6RyS7ionJlLEQV7F7gL9kUic8r8xjGtZ/IkkANWOh7cuHqlBsTKQbi9EyQNbuIef
4yZ8aJNdCfGg5Q9/Az6RDWLoQ1y6Y1Ko8y2lYywpUCgMczFsFfotzY7DZuMc3/R0RQh0ri7Qd/To
Yo+wMf7QtZfY96c3imUmTMiB4yYsMf5SiWxp30mPYfFwO+YlaLG2MCIHkTlBPE7yBMRuIpdv2JPN
ah4JcdGa2bRBasVN3+Ox6lLUaMWT8MzYWeBvRisup0iM2SO1N2jnDK3tZLcI5VvqPZ0VT/7EScUW
7kafyEA8YZte4Qa8ok+NXHY0mqt8ZbY/51qp0x3DJmS70ynGDlYF7BF0ROQChOQQFLkX5gZC2fyc
vlBwSm/ffNbtFloMRF+UMidJMXHqBdEsb458xhidM8Per+KJ0jyg+zFmKJHzyWbuGW0hH2hdxGWv
WmoU1FOvO0YMQnFMlbBwg8k/exTnz8dktutf1Oq1piNs5yu3ve/esORdS7Qr1OuGe4j3vFAgQ5OL
mAsvC7CijLdBmdXCrsOz6UvTZcu3+uw40O6AdQRGnD8FUb6Buw+ppObyZJ96S9DwabncUxaSyhWj
q8HVHv01G4xqDnsz8XJCpdsGyFD0wSeGoNqLAfzu91Zn2TjlHehQyTsZ8oOqO9GKjtzP3KWU1RMT
FlC2cAAyisp7+KFuDyK7TszSpTBn8OBn1YBRZ/KcFComiKJ11o1o6RCMpJmGsuZc+dH1zlukA3b2
CATB390tMAKp5Bgxs5ZLjmGQk60LUnf1BsTG4wr3pzJG+zZmUeVYRJ8XJ8H7oAtVVZlQsxNQn02c
iUHuczSy/dZfF0Xs5gQv6QWLpw0kHJMp4MrqymDNWap9wf12oR+D4cPqp/CnilwknlgsxoDYRPw1
rPXgj5de6BkUMw3CDzcGD7W4lk/+ApBlFU85LRqIqPVLh8gssKYfp/mj8zOsr0Rpe5vIm4SS1aLs
iSRE/+9wlM7hA6fgFYp+PYlYVyre5rUIOV6250peoIlou1gaaPauvujk07gK+N8w/MAaGUps8QYc
Sm5WFIJKQH56kt00hD/8kcmmD2mg0nw8JU10BgBw1Cy5SO6fwmpFPBHNv3ff/K4i6pC8L8fbwDJl
7TDT/2aCvP8+jRIOWuHHirOJAAVX1htx2F/Sl/yPPFjDNcghCioTAWt0piI8XZ+qmGZlN+MVqeZ2
9ijniz9xTnb2XiXpnAJQMSio9sC0jt0rGczg5MXrqWDdyrYqN826KRRW4ElGtDEXMYPkN4rMtQvV
r9aU9L0cDWonI4nQbGzpTPaD2PN8Y+ltJV6i3QgHhIimcIKiyBOqlUuDzp2l4E4vKknpyq4dhugl
CbahMAPtzFAo1JLkCBsxtFbcEVTpTfnhh1btLa3v0zOF6dEpbOmlihZdJ+aBH+pX4tV1Cpq5FByW
7WLKedB5asJoUIDpWIuyJEYQgcev97x1+amVfTdfj1eK9rdwmSEhNorvLyzlDknJkmBgCfKSshyz
xjqjyk/1oTHWLMhx9zo8JBY89JYE6JtMlzg32eVs8aVJRG/WY5ezaJ23PpYt1Qe1CgCa8NhNMiVk
bTQ1Uwsa/SMb356gj0XUrjh19SLLgKQ1lfUZb9qYVtfr2W1lo1WfGPghP52Qr3FUs1N986wJLmG4
ICMPaPcDrSVIDSpL9dXr2O/ntOz82+WOLcw7wfmdht7KsD9qRcRZboIMC4t4IW22wt9EqA+vLBfW
Di/2G470MyRdRCvmvqw4sbFuRRnWgC4pUdmw+eOnRBB34pG2OTL77I1VSDojYJHv1WEDqsS8O2KQ
YiOoQDIRc7tqEpB5qgEE9GXWJnB+h2bWK5X0fLR/c7X0mtg6H2NAJeE9PG1InQzdyXTupQnekEHB
+EivcmWi97V/WBFY7PRZbs+GMwZMJk3GVAnnqOhbdNm0mALA247cy1AH2Epwk021EamtGXdxOiZq
4WaTFNduza/LxquenXG+Ahsb7iowTAzBWaF5jTFWAtXb9Tbo/V0yZI8IcU5mM2vPo6ICkHYXRR2l
GHGYaC0p8M59ZWW1YLYhFxLzlu0WjJ2m3JGeZRdUM8bh7eiJ8ojbKyr8aPuHuk+Q8gwhQM+FGxIp
fygepKr5KWhaGCXpWhuiV6/CkSkTV+H8gHlwthP+TB4O7dH4OOkY9RxtfSGz5FmFUAJKKH0y265Y
Bn0k8Eh56+moAlrpddu5f3mQtJRcCNV2WGHrhAvXSaJ5ih87RLeFtLUfIlBPZfu87v+XMKam3WOM
WCboGD3ZE5DH9S5pOyPh1hoaRw8QaCMO/v5ei8AWZ0TmSXGWz/aeO7Kh9FPy0y/n+eFeT+k7UN5p
I37WJkmh3YWMvZ9yZlAjp5zx9lFbmBE/kIKYat2FsCObH1v6IYpQ21/ryIcKOMcEWY4MIQDtb6/M
+Ho5Ucd4GtSdAoQ1n3xQK71FEWFUJhf8tYb4uruDWYjpNGvx8OmlIFRIhrMBuuHM2bkqnhPg6xYE
z9K+0xUhYBXUHboAynFrBEB3xhZ/SgzLgV/QlzqvQlUQfagbsXfUo3sBXszFJwlTHBxhh1PRbYFy
vARgT6xkZgJoWvnmN/DnHldjJ7ja/MYRi0IpGj8kVSgfHBSjRLGWl0idFWEMRtTa/ERYg9+0i4yM
e88on8USk5j3+9W2P2yQhn/tyJF2Lk2kuby9DLSVDP3E7kKdpGh837xytJDA6KoCMcIv14K+jLuc
yA34IQT/hpa9s5gZzGPutRnj0vWCWJEFIvJnP1Ppt1V9fmlkQxM47BTUtlUMVPYYPQy5ROoKW802
sOKJkvHqfPt0+ImaXHe57zpCa9zETMIUTk4pFQ/B3ka102xBcx+b4qdCw1yoQucKJNkE8CcRd0I0
2lxDfx3R5cu31+O3bXZJSQ7idS2oopPFdUtWChjC/iwlkSCysH8ffhOg+P1XskreKH6dyhKYxlfv
C8Gfddlg5L7bm0NDwBBWXZrLjOnitD4RJFBMnzYtQ2shXlvU2TKrEVBrnWJNs7Oz1hnsSdd0pVnB
A20Le4WvSSTZeCEj0DQA4nrYpO/SCgcJ5G9fdqJJpHbkOH5p3nvxKxtWqwfM79CZXF2i634Yp6l/
eYqxmvc1TYancCODya5HMXkssaWlUuOOpCGLSaBtq5v9Uh+6hUg+Ez4mtc1HJRGh7tLv6QP8UT+i
ENhxqTfdgqfkT/XdQ/XM0i33++t7IdQLnr776tA6nBsFZJESZMT46iDsBWJ7UPP55f3WmWhG58Eh
kmKxphxt2lrws42GoW4w+rqFo930LZK5gBJGms6OQvCz73VXBD3fxHEf8MZ69uFhcHLj4BAnVonV
c7cQwFsEJXSmxn0/XtuJnmkXrcQxvcmxHa/mVT4AW+AyZnUeZPvGqu86/wRCtWENEkLo5drX0uL0
u6xoPaPw8F9eDzX2QnaVM8qmWwp4KN93Ha+EY++dU8S57ANR/NRyKcVJTHdQ2c1p2gf2iKqxgPhJ
V1o9+lEj/qJOOVl5w3SoXkVUB4GIwTsrxFjqZ0dSh59Cduiek34+oDxZ4HXZbZjbbOc1Z6WXXL17
bx9DQXLVwfIo+3gaaKDsEhbAWDY3sHTzhxSOPtUz7AECcmoUzKFuSmfxTcyQTTqtRJ4XpOu68uQz
Rx7Jz1soQW8euu9cVvcPx4tQvQJZ8GFiBuA2WWzikiNLz5eUWl5HucHHcROupUG+3Xf5+W2B2Jdo
BHIG5+QiEYwpzyxe7UY7K5s+hu6e+wJ/OKRWbSWHHKpuNAweRsEFGy0MtgyUXVRsGCtUwisgIBmA
HH/kvhJp8S8Ob8Fd+fyLKCxlxOxpd+WZM2pMf+WMeKsiKAG1Qnwt+vJsF/D7loxRW5D3fe2/4YCF
x0zhdSh9cpL1Sa7u8S3NNNKJ1O3n7YaWXoDgIWphI7vN6RLORX3t2OkHPZv2omHBHGV1lRaUToyh
UxjFy0pjOp6G7xhEjPMObJEPiKdWl/zmohzmrMBGsi3QC3KRPNv7EdQH4R2hj362sQOl4HJHlh3N
gNknTBYNHO65QVyQoRT4rAGSi0owHaxF9rVJGojnUNPNxGKMaHHaXXHg/9f0EZKuRbSo7K0iObro
8cbj+9Tqik+MABTHj5HjuZQt4ODMF+t9Kli5SE/Ne20nbyywffIK7eoK3JIY2EDcX9E0SqAE0rC/
zGG0TEwu8qHzL5ugi4NYu3soz61arkiXuVR247E5M0l1lUs5/z7UVNM7dbQpQF2vYXqaRRu9eoSK
KwKz/kVT7Q6v2k4ednmZbyWD+WKz+an5zV8XhlGfoCK+fmDpxxgrg1BxWy5NZXfeTPuYi86KaZYp
OKIQrFwDb4pwnrH7dCwKKMlCI7nhbEu+tnzblWn8yt9542SEkFWiJkvwy90eOvJ00LxEjC+40TLi
jtQ39o9M/0K9DTlmFGMzckQjSbUpy3m2OMckFSZEnNeVVkv6O1dLWQ52+LlTUTS5SVzVbPydYYYp
mgRMYWpBhsupXMzEua3I+YO8qLg/5ULPgPkWWOhao38HgJjJv6Z/rXKEVM2eKJJDoG++g5rkSkNY
xYbFKDpadt+3yXlsaO16yA/yhRPU0iE6BH68PSRHdf/LNky7Z/LPHkbOBIg2tr1iq3V4RH2bYlnZ
hOHI4YuJqsCL5S3P66V7iE6JZCSsw866ihVX14e06yIfYt+1l4x2qxA7/93t/nvTdA6Lnl3Nai25
FWT7dIaLQMc/sO0OCKFUC1U7amgBSXpwG/62tzPUbqH5/J6NXcCbApOkR/qab4wsx967QpzqT+14
gCxlyjwnMYpOB9zUZGL3gvFjeGIXYwEEBGlMxp0Jbx3szmU3CaEQa255I1l3DGzVCGgJsR8gKJmA
lNMlrK4iK3Awa82SK4/0M95UL0uUl5EIBOSrOKdklrkm4M7as1fpu3xrKu6Engnz6R4wF566u/d+
rdaKaEC+sti88Y6DqbQ85b5i3v2B88a0G7osqORTa5dvMall/BKjVJ6nNALH0cF6/ZPeZ3UhyBW0
KIAvog3S48HtGGmO1LeoNlDMOwqZzg73x7l/rGuQ2se6v1hIcG/Ul7tG9aZugn6+Sow1mLFc89c1
t7bH9iQhIGaW7fg7MCJFIm+EmMdk1ex1HTnMcJDsHvjSskHmq0d3NaD2UI60H1nR61e2q/JhvYc3
sslTQUSPWHvs456zGnJF/Ac7A4DoTVhbLYBDVEd7bE7XjTz8MC03U2BKVmsil4VohOOGALRSxVv+
hf6RPHKJrxo7VyI+ai78/rlrQRpViSRLhMpQdlDqvXrAmn+T4aFt9wScIdvGr4p9mhFNdVfUo/iT
d+YxCo4kAARFZoWoBoyg53WVecpZjUvPFqOhGbmjOdpTnC0UDoBEjHnkchGQQ46Irf/8DvSn17eW
aDswoyaFFNDdQON55htm4OsjTXWex7jun707q0wdaiZn9NMsXHwP4gcy1jPUHhBSclTCba8QpZhl
nh/xbc3uy363JUzuk48Pn92+hgDNPlZahm+lPRc1SEJHHVWjmvjq8LnoymStYoKlpRrJB048YIzp
oNZvmyLEBFWkZA7TO6SJbG3tg0/O+PkPh/bApLBAppnsVqpx2RF0zz7zthyt+DKnXYTfFpyeGDey
E/gIElrsdxurTMFL2imDhZoLYg6hgHXBj6rmHGcc9vqqfvrUt01TvYeT/l9iqX4X4ohICY/S7NBm
/sYXXCNihzqK0gYaPjonGFvDEsmEPZfCvPY+NYlvok+vTWe8kFNB4NPQn+AVtmcsZRdw3gsZXpBE
jUCK/T+x41JEwMySeLm2OvgCPHejK2o6QgSRiK2C1yACbvp+I54dnQyDZ7Fr5S1xBGmEnrmaD5Kf
tYO4mgeB3FKqMr/6s7T4f/2FdDANQlWF5W+tKwD/Sc+Wh/bG+ehWlZm2s8f/mIzhCdAdfCkz6Suu
sRDY3kjkCWm0DTYG3QdqmnxDvFTX2owsQ8kZmMHtFDalDnHvID0AtIbkETgyWPTXZx5GnR0Xnmln
hhoRRz2afR//BShfSCXk3QHxhsem6H/RaSdTuZuKkyKEK5SS0T8k7ZFPeEy4yrDW+L54+ilI+fVT
hZ8sTPi0rOT5cwuKmC2481WCKd6uyguZn1xbG34FuyYTedDVPPBBJyKgKsaz6JS1KgfNOrmoz96p
60tUWRzpcZf0/UMa/nai+dufiklAUu8eNjNIDJSEjnJww4VWIGSCON07jzN6LdYtXB+N7dJihEqw
iLK7e22K/tTQ5N4lo3MQXi8W4L5qKeuOzrfwCoszoZ1POLArvvgpOgkCpL5B4wuyWb13jKvFkgdE
s2yagoNhJUAkf72HrQ3QptMFO0FWXhjgjN84itLOE+H7UJ3u3oqw8iizXozvbjsEtr/8xsa1ZCOi
6NWwwhNawJ0Xedk6AgFquGK7a/VfD90t+CQSQoD1vybIH3LQ6jAtZxhXpQX5WWPFl1RsrvZsuuQn
D3Gt3zy2KpLkqzUFd+oYU54xJnnHF6bnef6QEtRHyl31UbSWzgH3GQ48o9ydtseu6+Z3hMaAdF9B
Kn9K4FSBkTYe8yhtE+zdE3Fv+8y9/RCy+jokeukbhRSmMuC8jDqrChMNMUSKml/8BQO0NT4Zh4F6
/rzsMrmsQaCg8Vo3Ck/HVbBSmMwsuxD42AC5azRgFit5P8UwfHI/uXcSP49wKgck6Jl0+Z8AiYEL
EhZhcwSHqMT5D2cBMy/CfBVikuc3mpjtkNgLT7zu5A1g1XXuTg8Kh2WCr2gRGsbcgQG3QheehYwN
3MXiG/q9MIQIZQRcppqmj7BtQ1Xl6VLTvSyJPFXmOS7b+NUs+M8p+iZrKRxa+rK3UQf0dvDdCg3j
MWBV1ZlPm6CQk4CSfCla9yOZe/nMhcDPNQQ++3Hy/f8eCi9YozsP3Jf+T51pFIAFR9Ycoe0vUHL7
P8lXXsfZ0wl8FCAVh9e08VruNW5vBhIEBkeGbXKw62hSab8sjcm2iJArpyHnqBu2x7E86AfZlakF
xJ+/mhsVLAJ5oYp8dzAaSW2luYMuG15UhD2dnX4v3bviDFr+CtsdFGg6BM1R6oXq3By7Vr670Pcf
tj5dNmZflPBIevucWQtwVNCm0au7gQ9ioykBsmA0GSwui4VDUi4v2R4iWIK2Eoi7PQZRuLreritr
go29hYlGudS+2pH2ivOw+7voT2YhrbhmZn8YWawmDeHtoAW8aoBPOgQ3oISF9HUC1goGmvrvx1kE
Lc3nLTmKhy+9SHs2Q9BLq6FvWtjprnJFA7EqQ8aGq1nj6vOYLf/GOzsosI7dlLSeubv25zpRw3DJ
BoeqAfSvc3irl43YWTCJmGJUPjhATWQEZpKPcsxIYv1cdtjyYnaMCGzTZtDikH4alXeBO30ulDye
mt5s3YTwTALWciFe8L69eIHr8ZPnUyssO4XdSqWBwSSJVzWXNRc36LyYqeNKqi+Q4mwd5zlSa/ZX
tatysxpl5nhwpg9RUKpge8pcrfRJqmsH5h9WcgbF9ipmM3Zzr1mI3x6zLkjD+pscPnAnnLFwnPHS
rdC6N/ANc3IEI5Tl+YNIkFoJWdKEIi5iu95D1jg4GenP7kPtin7bx/Ysc2SmECrc7oM5yq6rOmls
EDZGCPVbAI1ygzxKsZQ1j1Dnee2zafeKcN9eVqM3nh8D4hIM90ijDjWp4arx1055yJ/OrTM8Incu
1p5LfH3ncq1G0zXbMelBnWRfqHbcBGCL2kJ36PtjX5CRbuEKgtMLRkzh1ltDPXn31ysxKjes0b2U
LZmGWTqFC5YC6FXVgyYUqCBVmWBTkNWr5N0IKHf5I8VW+zQn7r8bByJ/Zidm3FOISHhRdum4c3ey
8idJT3uaKJpTfSEhQNlIyWlgrz1DlteVMS9pa7xKHo1qra+4BRVmpZHz8aDemhYzvGazG++Cg5ug
H9uSoEG5fLVvsw+eyLqbzQn0mtJza+ahtlV32Iem513iYSX6DK7XdLPAG96nf0/YiouSaIyQsC/Q
J9YulXdgqkRJ4q9rfcHDmTjcU1LnNExt0DpxJwf9RWKNh49jodlrtSCjlxDg7pmcWsCWy1dIr+se
1Ig3l9Kkr0NDxXoQM8chcSH30ul7yLbFjnwW6giQtS5Zj/Mcv8cgCqK+FjjUuIsSxiHJWx3vxKFI
PBM920Ld8w5u5vJOjuuo3DnyXAhImhBel7xCyF/HIFwoD0bFyxQrcx1ij/0Y7OXg/7YV5kms+HCe
hUXZ23Be0UGl4FkwHGJWn6wi1a39bzagTnBHitU6Elhg4jXyYqcC4OM6pMzns2x4LUunNAaZgohU
+JdE/zH0NtHATMtBmbBz2Us9nz2u/K83Zyx1SGuyTxvBjX4CbMJ3ylalTGZWU98Epn639jb/GCtm
9+77wbDq/DRWmnUkNI1tbyyMqx1VXl6ptB/01cFPQ98EPPqMeSGZvDodsMxfD2lcwcLBwHyKVU19
IWr37zSVs8tZs49gJntcfiC0jgfHMgIN8QcZ1ZL4Iqxljc0Gq596GuP6V0IDquI8nVMuHJZYFSIm
aZ559pdruSJ//y83O5yh0dQJmAgZj1jPV5RtByspwveaQj6FiBeHv+JkD1flFpW3PJWV88vjs+q1
SjBTCjVTQPMb7Jlqy6iLEdXE9iSgi9GygdURjVE0ZhHCwt9Gy9iR+mOHELWOiWtQXGeD7xzoZgF9
Mu/dKLnnpOsUH+OIPl1/gpvPbT1ogWBZtxC0Cbwc1Qs8B7Xqw4a/33UNNcghkko4Pe6CYB2yw869
Cvvj/8jorymcbJ+mvzgdgL/1fWman3eeAJFJlmjiwOeF3Sdfc94N0JmPPuAPAVHvvEggw047P1vi
7NfPRFo3NhgG5NsjGbnNsv5aeAlCFkTKjQ4YOK6gkvMdLTSS7rkzqtHg8Sgw1EeK6DS5MBNBMt0T
RwutuViz2j9WwgyOl1hcuHOesaxGSmK5bMF3PlplyKD5dkfUgVrpnnb3pSi8XWLY+z/jhMpPNT8p
kSQykrSppoqkifs/DKXcSBXpBLFrwDpv5CQY1EGbBEVTUSup70ZzW8SpvVU8E3h+bVwn75IggRlf
M5awAE11Ycd/xtIjkdclZlXp5w2zsj+1Ucq7qEFPrtrCZ/o/p0uZ65Tfs45QZ2pyOmxU15Mp2Hxi
nGkvXt5ams5UAm9aMLbFlF15BC7jM3NgNMHwVPVARAqpKDirSKnrsU/y0sQBTcWl4Edg4LrZmTVb
+1R4ioU4DQ2eImcX18e16gQua66o0okSBkNw7qDw2yjXz04FoM6V+u61wV81OVXPDSOdW9yEbWE4
ojzS+px/2tZmp/c4eFDqFKSsQJAxtkCUnyuNcnZydLBB+qokjh6nlaNPF9KRT9BX94QdfQUGdkCn
be9JK4N42DhfnltYAeJ78rjcPXq8mBVMfvDS8Yh1WxgcGjg00vfcETCZ3NPUBi3xh/m8/b33bEMH
WobENDM6hsAgR9UruePkuMc+I2q/ykhqwNUVlQja2iZOdjyDXp9Hl7dlPRApCpbtuqdPmHBxIFOG
duixc88U8FRa4pIx1+EJnBbkLgpBq3InT/tRCIO5nGnDUo64dfSSj7cSPUKFtAgR+oR2TkR+Wh+j
HmcX61ELXHKwvAf7krIA/sPF46ONuILnlW++Sk7MjYITY3oSlyD1iNh34ZLJYzMNDX24nHogbIUa
Cx5DRdi6Q73IBmRsGLtW2RBqLFa9KHnI5xCdJZbZPe4k74fZFc0xLUG5iZIs2SDXNvW1ekfmDcZ2
lRaXeaJoqCg+nNmYrcxG3qKCELswajIpnVkYRMDV7aLlYVFkGO8mLMkcNBmSn+Yh9qDyN2ok2K6E
77VNSxjj5KkzQXfKoZoJ05PVS4BvxY7BmzYkEQAHyTuI1kJ/76Evqz50LXY9lP2uYTvKuQ1N5+Et
IhTaUqRI6yFMYKAi6hr/HRdUJe4m8Ghp3+mTEX8yDIlrFTuEY6TpeAuu9E9h1OZz5iH+IIqFpi98
En0ryGf4TRNO8PUE7ZKdIGx7AFvbwZI8DK793B3HXMmE1Opsw2slLjUpPTGbJVle+uNRpnlLj3fH
rldSBX/PhV6unGdOK2SyWSsJkBNxM8gmJ7xk2wChDEodiMp5dgQgeNrOKAIdkJ3tJeaVSQ/voi9O
bv8NE0UbzBEjbcMt3SfRisG73BsWiWBsn7Mv8kF/im85EHigTYvEfauemWk5PVOO+WaN1SkD9kjD
nPTNjQBIWIzB3+eCL3+aoM5I048cElK3JBy3Nd4ISEs7PsqXDe2IEKDC9NfSgu12ufZsObT5r6q/
hOQsYEH2bINrrVcQfgl8A11vEv2enh2CVklpHreFBbimfEZKAtWLMIfzJtdxUzv1Mx+/mMZQAOKm
nr4M2f65Kd2ZB+/wcUO6nXf5KqSpDgg0A/C+cX+pS5eUDU4Dm8QxPC/dZmg5Ouzs3TCkHmWgl1V4
vR+YTOKY4/CkPy1LyrX4DLeeuvukt7ubYlEsuHGu/6JWivr0SowTJxpIjOuI+mCm+Hhg27kO+CLu
3w2po9IdKD5VHW8EqV9pfLGXWRYBq6s2JseaU6F3T2RSGicEfkj4HZM10Q6vg32VGpNH7x3s4ygi
I4JSsNECbbUGZd3SRvR1iQTh7EHbIgCDxzoQf0bB3R18hYS7NI4wZDWs0E9cH0hVrRToErswvh0y
1tpj/g+fH4PSMFV+HPtLu8ESgWvGTQHvQPxT764enwdfmLYOywLLtolQEtdFt0DQGzKmn1gUnH7s
Q8+YbosGcSV9rapOZonn/MUdZ1jPIwIEHEklw/gi4kb8VgAT/l2g/PTLYF8ci34V9UoccO7CWkYs
V+Y0WyNCP0MWVDyFG/bs+cDoCgk5JjP28n6UYjXaSzmu8M9thcyIua7AXWQ41kEN8DW3vNVlXf6X
pmB8UOuDuZVKZ20DvNnhioNwPHP1zvU6fPUBtwkij+hzcu0DVTgRi2H7VipUzEkpwRyjIsxIhqk4
3eqbjUrZV7tG8ZoRRr3ewaD0XLa+Q3B+ddO7qDNjry/GG9vqScCNYixsjfmJQZbACLIMYpXQmbph
NDWDSAYiPdO8eb/9OOpKuHq2gklatgIllHteliqENUasl762Dc61R1w6xeDejfViXHwxuVKfL8ED
dZ/sIARoNRu0xObNyKwWGSatO9qR7Cewtuk5nMrfeMm9K/ohO+XhdiwB2wUDOx6UmB5bDA/5l0nn
rjx7BM14vXpLEiKzUvr53oBRiRH3thNqnpVqGN9Jz7syzi7gFm6vOClaA+rgSGKpLMWNsOEQiEUe
g8T9tjcfNTvz4wiqDowNbkcpVY9gjtEbJOh0/l3VpLnxGwxtx5nTS7blEP40iYNP/AJKvH2xcP0u
icuqO1V18+5LBpK7SYrKLzAwFx2YG0tUZWdkZr8iu7Dzhjr+yG5zqDA3FcHjDkc+GQNib/iXKH3d
do0H4gQy8fGOCyn2mVR+P/zX8H7hTljGty3S2jP3DPPvB5/YycsHjlXNJyZJwUWXBOE4qVt5dfCT
07V/uAn5SBTA9kMQz8jFDFNl7/s1KDbhsbdX9w0GO2K71qQ1AcP9XDXADoH2t+ZJo4oYBzguB1Ad
91r5AIsf68eH56CO63aVf869IrYKaFXvSs2LbMYK2LKeTOx4rdG4Nu5Sy7+ACYG57RegnZBgR1N3
UYRiTY92EtC5dnJ9kEVs1RCpWNOcDfZLcHeX35SEGnZzBWon1mwzv5u8yQYlaVq5+qfO3DbMDMdi
DN/iJhNScdImZJ4/fw8c9dGPnBVBMCuFqn0767+45ZXKeRJgpCXgThXqSGF1yRBWx0rYixlqPNQV
uj+ZTFoEtgEkTp+8nI8B9fiUc1BHaUUL2YU6dXIvr+3cyxvXhMNIeNrTLoWynsohZofsXhwneJsD
HF12RaOqOyTdisyPwCbh4oshUvUdYcuTYuTDsKV7JMUME+k13nzElrQfOwzRTsUXGxoweljVyxUN
6+I+gdM2fw2ldEPk4dR0vJF+rFwMO2MwQMm2Aj67iuqKrj/2aHHBPgr2foNAYM5oVS2+ZRfg/KL6
hpgMl+gqdmV1PA/dvaUb2VCWVlodSjvKvbCaLwtHcjve7aLTJCSWXCxW9j7HZrr8zSWBVm06B+Ds
aPuQlNdbW5RODXfwe2otBOT9W2YcaepsAZ7zeSZM7M4S6UuoQyMUhvWLrd+zYXW+FYLCUYrxN471
6NETtl/z1fwYWDGCJRk89CqrvJbNNnwD52W4BUfU9UENaQUB/PER+svOGopLMx5Gf6wua2fjxZlH
3h/ordbQ6EGlPhGzCH97ECcpJyUBGrEeMoRpn3qaS96xwPMt8+jve4OWlQtrw49fLJ8Ix9Xvr2hq
6xeJorWwzoR/fu8qYxRhX47uL8PgHA9OeU1JNGHmDSIESTQqPMExR9F/z+YBEsDO35OlFuuZsQrZ
ufQXTmz8Kf+UbkTzEPZELE2AAQbGE9zRDoz4zTzh/In3k6NQgDCzuJmL8M1MwOfMKQTkWB+b9hqh
2MIP0mKm6wAKAN/5/94S+aI9dBFSY55wkJ7RRMYYG7lOvxpklzWfWdkeW0VCSwHyQw+EtnZ2Yv/D
ag//cgz7kB7HWPdw7u0KUfLv5qH0HZwCPSIo3answQGHfJYfSCIDMiEdIV32+tSn5Vc1YU9XxoQk
83DMz/oEZHnJa8khLx41eDJYGEhLu9ZQnzxlRgHtkSiLe5RMAMqxJp8rRMZeBtWlyI84A+B6hvyi
GXWx7j5TBX9tROLfFdvwW0VI0n3to1ES9FntwUgzmtcAgIqIAO8rXG2Rlxf/UzoUlVSdT+B/XIPf
V20h9L1W0uNnhMaim+31CgxuwwVOr2Ukbme84IkA0SF1mpqopH2zo4H5JXZzhf8hHrf6FWGmR6aa
qUdiee8pTbJcTwsORAJaeYbxe+WmMZzj4ORxXRQkODS5XZo1HYYYzykqlNF/TZuaTYk4zGQh1gXC
MHG5UlJuIALpDMJZJY+3UfBTCHLymp4p3eHGL7jtm6H3iy7PwCCdwdn6q3ifPpATkocR0JNa9KlB
HquXEkh8A3oC5Hz/u8SVfHuP3nhUMVCZWhEgORmPWEQki4K6t2JSdcQCrPIxY+DBiviSEEhu8g9F
XmJHvVBo3WAOD3QvdoKWgg7/hTjWcpBHDBI7KpfpIyiSEoZRzhziEW5Z2yQ7mArXto4fBxPDZsZE
QjjsBxxfDU9iHaA0heGoGzwf1Qp0uqv2iuQX5b/GUpqs82yqrsHaDEsolKkMzkdDS7RbrzCKqHD7
CYBZod7/0rZLB1xctVEBNviK5uopkU/dgfiCD6AGItevnBGczAFYzmZEFnLbMjwBN7Djn83W3dfq
Hkt9zLyrqgx5SWUPMJ66/d9vrCXB1Qvrt6qMl6xnj7O5wYnvtEvickUdsZSviclz3gAN4xaUn1/P
tDbTNa4sxalfiigyMRIYnJWmNCONgYJ35iHXhKlMEi7/DnjUk/n2MqD9EVw1D6ASxlKuhoXQWApC
216cK0M59faqiXC7VIf9a+WfEd2qWEy/E2fxUEuXuuooQMQupXqhIYg/D3lIIy7oJju10ikYtD9y
y9Ukqho42ikoJfDoYe//iE87tVq0MliWHP6vrGtpk4yHXkrQkIsYEZ6kxTAo1TKVMQssjjYZBFID
oZar8FAXyQdU6iBaCS/TDkAkNYvT3GHBQ6ZA2M/35cJyR8182b6eeO4FkwGkGhzKIcSfZ2VSaK+f
Z0lgTYfC5Lq/9Q9M24FpfO9LNUb3JaDCM+HgqQTqapY3P07qf/PC5GGbXjgTEenfB5ERF71VdMC3
qJswrstsZ/QNiNqCmj0Z+CL2nNYWAj2U+WtTLfLvo5edFjAYW/H/43VxMFNmE9zttMiK4rUxkiH8
H6C1HObJVonlk5pg5I3lSbPA19CwY/2GtxBq8j3jAOa5Kghpdit4FCo/B6wu0fd6IkQv5mF2rKHM
18+Agt9GOMrdu1V9ASGDkXFl0kNOmQGf+BjZZqIy2lAwncpQCGCeWGiqIW3dNqjghuhtGhyvT7Oo
NOfMrs4aWHgaYp9k1VOpg27utsddaebcjJPD6xUn+DBGis4aCY7b1pT9f+CJEdouAx6oZgcueidJ
kDQsiru3WhkGiWuPky2pFzCznHZkLS7OjPqyYcygpcEHLizywDkNgqD4koU9YqGp2gwWz0wGKqik
99Pwn+UPnaI195rc1zFzvI8BVQRGCHrQIKK8hasoW+gVQRWXypN960wIiRqWHD28N6L8isyzQbME
Aos3R01K7qCaKK2AfOCTZXWCiv0LtQS3dvokSzAjabVErCf1F9qBwHZfS/KbkIeIR480QPf+CmKN
lk0BKvaogr1v6pqwtVAzto+osLik4T0HndA8Kd3A3iVUSonCmCHIMcEMSnpqK4F/pPab/y1xptC7
PgZOJFZ3RCOHT9QflI1c88imaBUYNl6LLqPMG3i+JL33vs9uFTzoQSvyJ6ep14m65HAHWA6HkweI
hEu6cr7f99pWj7HYAGFjTGlUqf1qIKapB4FSO3hhAAni6h6hDh/LNXqqppy33NM4mlAOu/oGG0r/
6/GsD8lv1za+IydY1q9Quufk768JNgkKNL4C7wlHhn1qjXebroBXNZgCmQbPLkyfSY52OknMGg+D
x+QJj4x4rll4TdEFrH+EGxsnjbIfpSg5+/IanvIG7mHebY84KiDg2OaEArwImDYEpPGxgwNZb/oM
FStPu1WbwgO5gBbuxTF+KvNVcHnemP2dhMJ9VlpB1yauO+1bWoQqy1q/jd4nEexqh32XVubbIpTF
zEfPFe2UvAPme5Zm7BISaQE58rloQRZK0HvyO4zCY0Xm+M6fZvXChxZV3uNNi3fr1olZgDW2/88P
p/l74uyYM/fs6Xkv7d3vz6NFJKpjolw1UzwnZG2nRahkmyhCG4W41p3yVpW+xDnochDfo1Ertq3Z
Keb8n+yfnK2meZmsHRSKBxQwwOkeZiXl92VAabUYbG3i4jq3mKgyKK3V11xntexPNq6V1FdR8u2Y
1FI8wFxvjxEPqWJsHqmucvjFcBm4T8zW393oZtSOFlah6BumPvAXtTXnrUyxFWVcuAEsIOHLOuGA
Z/0Zj+qVM1GEaZUTxmkIUnLjqSKG1yCrMOsXQy2dNiuRsDUsEs8aLTtEF9VNL3Np++94kxOF74Tx
DKrjQKGdiMlEihxkTXPvQtCt7L2sd1mcN1RK/PjQAg71i8bAArfJWHAdekMDBm4Do+CXhE6Q1T3G
41FWIwa7mlc3aYzCGcGql8dxdzqyPFydTbsvLSZtg1bmpWPYHi+/cBcP2E8QTIyU4Casrk/kA0Lv
jOymDyqRkdk9yUPVxA3Wh37N0UlUQTSmGJgLC7UtXl/bKk1nUa4Arji36Ds6XOX9YndylHbbCTrU
ppNEkrnR7jgoF3bym2gpjB82AFoqZtiiR9ibcNZcdkn548tLQZRSdqjI4aZcidTY4yqGhXsXoAxL
73MAtoBXfzs7+G+UXIdd6TBSNMz9iF41UcaF9v45wgGHU6MDXSx/1aGGY4yw8AIbloo+mr0E9so9
GxpWNDNPMdoFIRN4XrvAp2TZOT7EU5McGMBuUR9/QGNfKAymintKr6B7suAy5OErw3WpaOzcL223
PBH77+PU/DFSNaf2TRP9hgZI4s5FSEsHoXGc/ve32PKZMX1jZoMaMG4V/VYs4iACznizhlLn0fX5
m4xCN2sPuiV45jMQG/VGjvetIQahLDPLEZz4JNeyPIhM/eMnSC75L08CyQdcMqjsE9KdN5MOsr9H
ii829UGYQ78iwnp1mbyQJlfi+rJJ0YWqaa66mVdJDnSrhitPQlaModVg2drpGtd0649+bYeA5G4f
lQc00++Nshdz3XbqxANRSw7Dc3sZzQhtifD+S+yZjO7z429BRRqwL5O5cFp80zs4NctS7d0aZ5Fo
5OreL8slcMdu0it7ubl2YOUvGj1eNk/Hx47iQWJBXhuoxy8218kC06PDfpcU/peawhrQjWN9WIdM
bv5VS3igRO473U+uqVAtDXVagIMnLcPnHcAI4soXNhChivvOJXfF/1po2Fe8ZXlj1qfzvvTxKp1D
RWV0iyO5kIAQ6pd+a4cXCGONP0VHLgwsHv+dEmiQytlIC4zU31YTVmGfaVBEp3pQ1Kdx3V8WaLTq
utFwSMWlflw6ub3yGlf47au8WCDGUHf3VC0ltDs68trNyqJT8YKtRtVc2lLV923Zt7AMclJB5Smc
XSfCu0qFg/bQDqP7oJnsd5oLArSb7S5Pb+KHd89FamHuYaZhSFuzX4/21niiZcnJsbnSEcjL06kO
PhKqN4QAWleZV5DR0jI2naLuX6/ocqbGDgW4qJ4kcmipHXK8xFQbbJ10LSi9jccxbIoFZfSReytg
Wu+OY51pTwORI7VqF4dhSvRafe1qNM6fw1TGkY1JKfhQH6Uji+Py4BSl5yReImHKtjNiyiW3LNKF
IsnXZ2QKC+OL0ndL24Pq0J4FMgbZBYlnRTs782CZUI8htQdICg1eXDsLrHsGCNk4WddCpgJywGJb
oR4FLp3/ico3EaTdoBLUR7yVCvxGQb3dHTFZtsTOoyw1CNv0SmrK6ju3RLMC6+7nkaG495FNYjT9
shoMP8GclDFpRwEB6BCCTrPxTlhW5acOca5H0ARGDfdEdCO0YJdZrrsOELwu+7qCmRLyC+mPnZ/Y
ncNv1hTnCPqtgyvRB0ZCvw53xv/xTtt2jE4zNueOCRynHOL0Os/ggZDfk7dc4ozYwWXOTxx1SCff
ZwIOQPmM12NjeUIQHUgbo/tdbOPfq7RXzrRTiFKXz9devbMAZEk9boq5RUwMS0R+5Pb37S1j4rqf
4PaG1FjfW297QAutxxw3iAonKXs4X5udqe8OrBYOuihJYy3q/ijemaVxe01oiOyRHemXEAx35wLG
XbnaCp5u+l6EVb+MqvCBZTQ9JOVBQxRa7I12Hlli8usBmBAupp6EwRfAp1d2CjeJwvlG9o8Q28a4
ZgLYQhciFbD/SDNOsLyj/RhnH4bQogr4BlSDTcYBXjPzQyBGh8zhf6WkvRde5dqKJdzD1uQqtD2T
9h6/gHIcnYUU0wsZpYIuofBHb5OQWGeHGAt9/uNF89FYWRbpEwnkiopI5dLt15787mOYMjNEflBz
Pnw2ZnL3TBoVB8rHYuGHEQDmsAEIK2nwnFmPZe1tdjBeck1jca4mQFs/JOhCTjn+hPZ5EElq1USc
t8UtAMzPjfrVGeZHyKk0AMQk4jp5e1QcnDk/wH5tAU2BRhvut9MIe6yd9u73So5vDWKYbC8LLHuT
SHpPe/Yhe00l9Ek0lBqsj0cdOVJM1hhzTMvZ3V8ol1zrTv9m7CW7MulhCdggzJ0b4Mvr21+GDCvb
rnbDbd8YK1Z8KM0RLC/o+yJyGpXzF/Pp5Fgb3TN49EoGUnCSM0ORFfVwMBlvqb39cVvNMC6FLogu
SO374N+pHXMmmo4VH9/Fq2ugYYlpKilsKpiA/SjhpRXTGpzpbuFA5FpjSNF8snsciu01euqjUUc5
neqpNu+hkTHq5ttOMY7RhyZQZDQ458tM0DXY7jwu26yJCdHspf4lsYrdBJWCYS9dfdvM+AHxC0iE
Zxl4aluBgloPQ9V8AgknuJA8fD4bpx/w2VUdiG716LnaigcG0gJLfRVe20CDnVp+3eAD4wMKEowG
ORtCt64kst0CCH43j47DTDBzx7DEujnC4NDumhaNY8HaXbxVZqvW4Z/8Dhm9kD+vcNvxN2OHT89U
S8r7bpO8+L7vDLYmVJT3X1C7g5zvbtU+z6fHe5qVSjohI+xDIdHcFKvdLEiMRJKf2y6yMouwwLn1
39NeHh03akiYtx7tbKuSsjImPTXgjRY1Ke8VN/4GyGnQ9nj97qiGraMotzbf89ydmUx4dK37ujyd
/jPgFr2NPRoYLHzrSGCxNghoc9yhEbH0/TBsYgiHRXhRoB1MemInE2fRok5uv8Qd0c7+QVYdzEeG
UYsOVUevvDleZT1T+8swrNfVHrsNrgbCtr5u9qBrbDBuMlcEdYN/DwHcT1Ssd+smHAHARvWKQqW1
I2QMGHJKX5B+nVvnEXEQYtoSjVK0tYBwigxxwqu/0nNHqbpLHtVLrkbhXIGb8r2AvFjAHltYE4XM
Td+XdqbeTh/CxIKbe4Tw8G2ckeJftMBvvKV5zqG4icPBL1vNhHyebgOaHTAaonzFEACjBjM8bqrv
qFg0uqH4D6SPEsPuI/lT2QqSZ7F4XHGa8nRonz/bEaovx1xxi3h3GOd64rYgVyuOF1jNiHQX9PJW
OCFzt2Zd/3IS4DZWDTysNmwUHn6Riip7Wt0loLogrrtoOu2KEs2qotgOPSUajVlCASiynfxUvcQa
x3fFf3ysXXxsJvHtHxt83D9T+zxfATq8EViqawSSG1D8I1p0yBmALFZPAHFwwpeVWjECPdlXnvEF
eXKESu/A2Ajy9aezbfPuS4KPYyVgGQkTlo6+hLC4TVknHlI5xjRSGfEfjH+7OQ7PbBvDmLK1FaZe
ueZuQn32Qx+hjHTXufgyfXDB2XUNC2zJaLPzcZ2hGEdQRC/xaj86weYhe3dghULaS7pgUo2ZJXG4
AdsSBxxiu7J/QrelOkoCLWsHF4Ihl8WtsOnc3mtJaxvjfHRlLlzJ3YoU7qjgaeNi2DJcSomplY7V
o/YYZDJIKghSrfLooIGXuJA43yutxS62p0R4aLz4Dl+PIVLJ5aYgmPiXGyQx0IN0q10Y+eiXEJOw
o3rJ4wMZz5YwmyBbGHIpMPsyHYKpIDXIkIqhseH1yfK5Cq9Nl5zGONu9rmAzo0GNq9ciFvjrPPuI
AFPUHqhK23EGXsg7aAUALEZjBDd8pt4uM8Ng76U55Ax4zF8CDe+qWdEnnREKmXv9w0Cqbf5LiWXl
n6BTxnm4rmg7S+RybC7wr4QDFjfCz08J5XonWWEWKvMUvenEr+ekSxCfEcWVTRHmsYgE9i3atxG5
v4HbzPUzMNciuw+OoBOMb50ht+7z5KFy1P/wqRMd0EjT+G1V8tbhggiwYAI2m2GPZfON2miMdRVN
MO6s/yWJve0g0IB0cO3/pWMQZFt6ZYMSE/D/nj4d5gmABOng5h6ts+dswJ57rw23ORlyv8pYMpof
6aO/VSAgDj1TDDoaCsg3UG+qOm7KSCRWBm5ZMyOlHfpNKQSvfQGJQ5hFYwLH1xATQaX8OochQ91o
auPYqG3A15W9rPOIHWGqje1ZuGTyJZDFj/IfLjiOKgv4DvmDv+Av7MxqQ7+6ZrpH3WijP79ieOtz
UMY0fJzdSpx+8EnxWG986FsAoL8z12g8hKT3XlcZoe4exW2wSWIrW58WnB+gG+RoX6RLkID67pOV
evJLIWpYvciZWKDbJayoJ5v/A7IgpUwomL1Dvz1uCfZVd8Hqna5bD4HhalCnggrQzqnYP/OoLuOg
YdGZ3o/38BgaypLHBSKIzWLCK92QAzMXC98u1YL74QlsbcmXu9g215MWk/pltNGenjmPWiLla86m
XrrLrbsgMcan2BWUUG8R76oP1aJu3BTEOlwEix/RzfOlGHN3/KLAlPQrPq3NDutcwLSIocl7v608
T5aVQT2SriqlW2nz0rrlM5tCOWiIcbBnUR6axXM0iHRXtw0Okp4S732anMWVuS5x211Ia+Z/utV3
DIwiuG5W5qPFHCTMNxWX3006RZADM15HIzF5DAKnRO94F6DWcLIKQKiVIQo0TM3F7UjSfgbwsDsB
F7fRlodWDx7dy+EsKiThjGY5W+Q0fzWX0d2pN32cAQevreHQYfPuH+jTI7lOGSCg3eargiZmhd6y
PizhmQBWnZ2vYpqNAR4r8YIxCDpMVc4AEuglg49Mu0Q1bHqyl83/1MsRnHqYTrQ4T86HSrxljqjd
PckqQT4Zr+7FiA8q1P13jJSsCIiLX9zcjIeoT6e2flE9yy2h71cLEocP4tLjapMg9CGTAnD/4rzf
LU9LeWAGCkdrsTexfPJNwX0M7v9smc31fxKMSCLiWA7mYpjVa1GdyodAZZSG3frP7rEIjifKF/x0
wnErnC8moTSHWAatYGbzzYZZxX/+ftk02RwzN+Z7rRu3+IjKNU6KUE419vw69sEZP2r//vG5yt+H
P+KlYxCeNbbDit6dKI6qSLza6p3StkN0iKPVOYAKv5RlUEa6fQAY6npHI/Jg9jGk0vPJiCFsklLz
L3CXvPhnFVr3JF2YnO8G2wBff53tnZsUpYlDys0oQZE6s944sBFUpHUPCvN02+IIoSH63L0glalf
/Ef/bx+4iR+dZyEu+KD+0EJxNvWHddvmQqeSNBHEWPWkol+nqS+7v1pqyUdQ9far1rvP6hYmIZvl
wPlIGLubZxkXK/uQHgWxNuGUM8caIB+fzK3fITXc2jZKhNGrRtRjmSiIYSzcg9UazP0kthr8QFyv
HkVoPxsvL487EucPNv9NZNXc6y30d7pPhNK2mYgtiDHn+H6TbWzb1kPtbIqw5Q0XguzJSmA9oQ0W
wowxOkabky7LE8OC24nT9yq92W/h2ZS4rCj5s/nwuiy0Zhzt6+fZw6TUCRv5ErbAbAy+GzWIDtnU
IUkCY9HhynsDiEJRkfR0hstUZxmTbAvz2xPYf8odYJHgG7KZjFQb119UPdSMsdgjBN9o6gHb8eNX
W20VqNDtDHujFSpV7yuW71VLPlP701aFPvHDJ46rMBFvaysYjUs73wsMGl4e5VlqJ17ur2OYW8wE
OsuFYqC8MwjTKf3bKcmRV6K4UUrd1gl2asJ5Ft73Uw8Qp1GeQp7AXNC2oiu9Q+7jy0vf3rgdYigE
0oONnyZqCFLMet5xSFeflAKSjv3304A3OVKswiUdUR1SsQd6MQ8PRZMDCL7yN3cmyObRxMsYBh/r
cvpPmm9uUk+p6p4b6HgdjuIFO5F9JRzVxRT91q655AlIj/yUoYH/hdlvkOysHCWUDQAPlmEucreD
Gl7C1X43n4V14XkH/Q/EQxQaI/DRSdndrHMsSstKms5H8Q43K1OSkoNL/RRmsQbIKJzOTgoAx6u5
Nylb/b0gHe609zHbfsJdXkcYxAjPWSlepGuB0271L2oTZ7SONkeFuuZKNB2A/W5y2yomcrtrYkoC
NF2ekv9iscQpvrP79jko/mCz3/o6Q+DkZxnlj98U2gCkWOPEmUep+KC+BqifJAtbzvg5HxaTf2VO
eA4fDCgQwdyzDhveKX0nIJOTf2mBbEgzfQ6Td3Zy4IXld9J6AFoqPT4dWd7yiSaCHbrNJry59OFA
w1HtWcWisvwNVE/ErMM7MetDAEyT/eGS/AnxqKYBUQNg46HfPvpsO0RCFeBG/NaCYLrcI5OmISlw
7xHwsZZhEwavGTyA3rQauky7zobGir+iLKqp6ezS7eYfxiJ4XqDBIXxdwafrIRuIi872d6fiH2iX
aWnqzVH8v5/KRveJuBYL9fqKL+vl+he7oPKqCJVKhK2hRtXrXtCKyGqAl5S/cibC6uMuWVxJJORY
6pCcMXyTTnht+6DReXkUT2WYTFd1OGKt68DaQwEWBJM3KkTRvEGDeGQv9BBIqsmLT3Lboik3YOrt
BnMq13NozwMlizrQWn/9/Wwrqq8iRDULzrxwh5X8JBtpDmfP2n+KVlL/Z4Gh2sYgLFTz2FdoIygq
1oS5ShiQCA2oSKLT0L7XisTHr9PFAsAasuHJwLyyf9Ady/YkA3HspxFVCTrd7dZhXjgZDk/vHTZj
m54QWunb/aSV5ib8oAuEiArFNgidBwyX1bLAej9EeQJI28tAQYkf1PCPLgMcQfWVswxJZP9cmsxO
4iZDU7Q4TROzcL8ZGqB9H/j2mB8WYfRN18zLJj8IHQBvrXmwcNr2eEZUQ4pPwIic8Fmm6UoLiM7l
A6Bu9u+JbsCkvsvWGuWgAet28slywYKMT8B99OP19uE5+MRNIjdBPX2piXzkQpbN9/bfPc1/fGTh
7mZgkqkM3bsIZSBz/nZ+I5RDaM1WFwu330XhIcqSi2/StfmqRsGHv+ATQ2KvE9vgeN/5/L7t8nBX
ijgbRylYI46Pjw64DYvE9r4wfkJ0fnrtYbcUBrM+vxs5M5TYWfUA7CeFbG9FKgWFknj1ftePd3t7
MRdL0KEKXqcBh2IBNoTj7E/nyIBSfiLriyNfyiGV5tQtk7AxviS0yqfw8fEY74FU3lu/ceAhzg8t
+e71mfbksgD3kqwa2+8BY2civRQWLXmWmyOd7Li9jJO7VVP8Y84lI7whY2lAGaQJ/sHaxfAKAPTu
THkLYePrP3ziRL1WwkaHfZzkZuYeF66LTgH/eeCYnTGGq8i3Oap7Wf2NOYTuxshKoIfjcFUUePIq
y71OaQJ6ipsa9ZVrQV3WRv/7kBi30kPqBoRZ9wuzAzGJc8whS5fZQ7JgyLhoRIWqC8++szfLigmD
4/CkkgFUrOD6oXw6FobHLSnKGiBjLKGvBeL6AP32YW6l6/1N1x3GrF+gIvzduX5TMbshMJ3xBtP+
SHlS6rCufcdKKJj4pg5cKfop2BffwaZrm3H1cMH5ZP30n00y0bKGF+DsTZUcQUHp1YlBq8VjQV+q
YHRVzfm9UxRhdkkyZvfl+dmunu8PeBQUCw33XHZXvofurrEPea3oTyZl/NEotzh6XMwGmIeFTs0/
fvZ98toZSCQFMDmwlU3FnWvjVzRkYCFjeZ0sx46m7oJ4VbLpsrSXYfUtkYbTE/3ObRxi90cLLcR2
ii+i9+TRf82ruqDgnqKFj0Ygf35AUxvwQBmQqAY+8qgNpoXqo9FNkbyyHq6S7a+k+HDmf3rkU32j
Dd4acAGEJ+2ZlUURtbDqgRRHLGsinKZpew80Dbj9pm8ErPjknenwzBXoGeJruzqIuvUtJc2jpLVe
+BANH7RkpBTcAqhsmmaXi8ZjbCzYt0CcI4VSpYI8N7EUFbVkfYtNHpu4I+qUNzCPgTSbxJFNr+sG
Onh7wpDAVcvjxRV/+d6bFe2T77DDu28fGW/HKQKzCWjcGr7IbrwubZG2XAJZSPtiJn1zTdMeDKSo
Z0NWTT6wpyUgaX0CsBxyTzWPpwVRPHl6uj3JrWtwPgRwdC6gy/e+BllX3jIEjtBugeSN88l8rnP/
rDkUsWHlbS0nUqUkoDt1LSN/RgCCCl1N4LjmQgGe97hvMg0nRvmBRH4uiFBXXtVhb+si6cDGn+q6
u3DkEEcOBf/gDf6FZ7DlWJfQecKWweQO9IP4eIEWkHKrjSzsB8HG7X688Eq8YI3lh+/d3QOae/q1
ESYIhEHpb+I48e/LD1obPrwd5n7F8Mf3OMj4YW+TgLeXGUJs6Ob0GFiWwRDmG6wA5ayDAOQRAcY6
sZtpoW1YTE14yMJOBJtAomQogxGGS+O+AVYT/mkVkHdu471wI9jGBvV4uarimkkx4NnEb/HlvFxG
FHRN4M1FcHS8Oyqd2RPr2NDbvUmbYa2l+IELTnz09yuO4GCK0/VcDMg7VcjuuamG5X2vwIyBBBJh
OQgjFhGOeDyu9HcWHOFuBUo0RH4lFYVTtP1rLDtNn8sxe36EiaSZgioNsMD9aLvTdh8sjRfw5xpd
uPSeZKpya+mnXuC9Y0HWs3d+tuWDV+sbduJc1QzBiej3qZWkNjwqYRI53UtnlxwZlw394b/CcXGK
EMjwX8GP9TJGGWl2KCWNKBTwjLYgp9DiUNX2vVeJ5TbBxS9T8UN582tCs6dHQtRuRS9XL6mJzhcc
vpYfYe9djFTatNddtt8suIPjnTPvzP05w0TJNQELfG0e5+5kS8I6vD8zAUOlOcEgnii1hIon6C9F
TZiffBgsBWzbwsM3PggFeG1H2xTKyjfPBdVQ9xCCu/CIzVred7w/YF9lC1/Ia4a9cWU80TcwIm2G
0wNKvNLSCsB8ZCa0ImSDyf9eQ0WodubZj+OPqtnCrW9++xUVI8u2tP683/2xUwmYiD+ufDBQAv89
UHXoY+2/BVHjVTPLq8iiHEAxYfqV3UCX1W/0tE1EIWfNIu8I2wxRk0NCtTnC5dMWTuL9TUrErA/S
XRsut5qh09Ga6ND5POk0uOiHkdNx4pd+aOGqZhXzfom4ZtueZSm41cyPL6yvdygWbztjJtDGBKNz
lLJrvfyeUErJz2HnVsSS9mQH876SI0vC8eRns1Q/sEnOaj0N8ibe4h3TYGIeESkYBnGY7Ts7RDJk
4a6wZuTS3DUzIEd4vjfUkJ3M/fCLw0JjAGFxhEoeZIsmbYZOdCDtQPE5mjn3ArmyuAmDsQRVQ5sP
ngnJOfTo7L5karDq/VG1RFcSjdBgkuJdP7u3uebDzCGPiXbEia2L2zmqUjmD3Ziw0lTwfUkrxL/E
EI+bDOimpNv1OJWFm9iA0jfvONoqQmjLrXhaEwMLgUAet12NtZpEfl8jWjbpN5kQ/8d3m3QbfWcf
6xtfs1oqF+iZPjIm5heQN1Y1wNFmpqFL11w0B5bvkjmQQ3Jo2cyEGmXFdaJYSQJNHOZuMWLlcgZd
Jqlo1Yt2CPGohUBq6azqFdfu3f9zImNOfdUky1rwKrQGNVJmkv797Py/QE0Iw9dEal8EQlyRNPHM
+QOlcU8SGYf5OKzPhEL5Uma/8DstdBRzrarLsLM7bQfTO7yKkc2HoPY6Hv0uxR+5eGrgPMR1CvyI
PsXtidLxXljumHXlny3skBA3/5jdFBhNM0abW/h5RuX6cqKK2TtCeTytTgbNa0Tvzo5UM+xm6ljv
bQ6rXHMCqF+ImZB/UT9mOM3z8XyZW/a1uA1JscjwpO9/0WVohJ1frLvbnwpzL9lKskRSlCWE9AXi
hbB8BE5Id9VjCQ7mHbjnYPDMmQHUzwH46IkBv+Ms+Fo1LYq1uOJkr08W2aEPUQR6JFQyyCI/Xpd6
bwdhXtUjRCqt68hIhNQgb+P3jOahicM8BhNTjAICHc/gQZt42Lc8TxbhNSek4Y6pyhfstMO3njzQ
iftpC2JNjcuTgG/j+ny8rQaNuo5crhJuyAQ21cisB9oiRSJb4s9XKt+KUi3UymTmbkN7GhHYqOqa
vXMr05jVv+Y2TQ+yJaD4QufcAd4uZ7cxZBZB84DLjKjoylW2ZLift8FZkn06mUzCc4Yr6WQv09kw
47a4DIT5auElAMmTZYpZABpPSCKWvpwnib/vDr2CEwMzQ5RkWsvIaam5uq5ktZbre8PsyTXcQuw2
XZkaq6MrscuhdIeFiGRwgAwqvCEMYl69MLfkoK24xa1+gxACvIOqHgyTRKfiPAKcIkLNM3Ca4Zyq
eO3MkyvXN2NIKJ89ek/UcWYZaA8H9/ijDJk4T17yAW4N1meqBq+0SkZrOlMsyywNMSkyoMM9GNyk
kSLFWPoXH2WmOx1qiqQW/EzBrXbnBRzK+R8DpIENi54YwWqJ3zfMgief0kiE8lmqJ/jkW0FRHOG0
hg+zrb9fLx/M0PbGyGWa+nnhA7GfvZuFUS+7GgHEvW2uy5d7GGXrHAKsdTkokEStW+HriwWw3lPi
OL1lz1Tn14jxFjsomVbyZn14miJpDMXMuVkiB20k1KyesoHnNIl4gj1kjbcCh9aSK10aOjoVRp35
T+4uO7ei/3fHGmGiTZEXPAFDOAo0m8puBpDJg2zGCXD4YX4QkhNlg+vKywc6M4Hx4dvTWlAhZGEU
QVxgXISndDp05ZRQadGzF3dY7I/Xca3fZr8rxAbhrZdvW6Veo+W89sNAJX2iET724KoQp5wcO9dh
7o+3u/6ywzrCPw9QELV+oxwQxiBajaqA/+PwA/Jce5KsNkRNWAL9eaadXv3LFiir7054VRVPLXi1
IwQtoUelvcCCI13F1nefXCokz4pqh/Icvd+KKOpaCzlLTKkldH/6gfcCxb794kpmiNJYuBTch9T9
usZ3/T/1h1KdSrVXETOOlj1UoKWdAaFev1dbGCH1WAfI4PvVt4SquCyR4moP2M6JSQLu3suQqjoO
SMkufNJiZc9ICIyR5t37b7IVYZPPF11SpQKt2WVN79JfNrl+rHnB/6nG6jhIzJhoylxtCyXIRaXM
MP5hcO/yrLhG/M5O1R5PvSgxMaV43SSBX4Z24hjrH9tonmXiAMRPCE3+PP6dHnAdlBrjEJjnPcW3
vHyDtLXGsDa3eWP2uf71vWFW7g67d3Sc+hPT72wvrUK3suMEQB2J408ZXuv30fJS90G3mLfjUxQO
SsXAeKB3OsVkoe/+UdvdjSlWmM6ZGmHR0TVVi0s7oP0RTdHqC3Gt9JdP0e/0bw781GS6yIBadk/4
VJ5Jk7+QI5Yh8INvYn6PXqG6E487HNX8klX8xEvbFlNEqr72ddtAeAQgCtM0Y37+xpczVy1mtEwR
WHmExoBuAs19ea4osN+rfJX23lv0Tk2FhfWSWQRiV4YC0Z/CbWmJ2fTKv7u+UkqDIeWYLQLMusu4
pEdglZKqGSvt5ZNI7htbp84xtJrU7WrhFYR+D2egzFsQy91Rb9F+uhVRP5gijkrroiEbujA8CbHW
JEdANthoFIgsfH5PD9I8QRokmvQ+sEf8+naH2PPO5eDbrlmZhVz7fSY/QNY2RLh2YuFkxRQ2OJY7
VaqOZPs5+PHXKiihc7vPItDdqzW3i7Z1nXbUKSPTsx9qLQ338o1Z8J8hINkVKZNYZJKUSC9rpck8
A/CV95iiU/HzkaOAhwLydDd0CFRK/jU0KRLVVZJ5B96ocW27T2p1QfHjGY4OuXAre8OXnNHdD58I
sLavoF8P52BQet+XkHKdd3txz/FDsJhT7XV/I3YpZMm0XE7rDYLnnL4LUjdYa8gYO/KsugNZZBKm
x49xCJMp5A69yxqgu/x1kMIwsDmt7TNQxGl50bKA/SJPKNk9Z2KFvf4MJPhYf6TdeNVg+rRU500j
TPnA8jMNtwCHAMTreNGhX6GMwzyV6GvKGzyz5fjcNDuYioYa9kfyvJv+E+DQIsp0DHbZNJ3yWmY4
VQet3yXSTdhvKpioMZo0HvkmwVV8GuYjiV5ezp+J+99ueoFZMWhPdfRZ0W4opcXqfkB8DB0K8Q/9
0FX7bgUlmfAAas2nBzDaObR5sDNLl4oqKXeHm8oKBKTnsLpHjkA5YEbq9WVUF34BZNV1Rdv5Awz2
hwSs1+XTQqbxLFkkMtc3KGE9aujaqSYzbumPRg28V9mIbA3fpHaZ8i7WWJT35l3L+Jzd+m70R7Fg
aP1f2su1qKF5rpOmUtAhXkw8KXkr6aUk6TclFv+xoWsJX1bCcCR1LZr0qqzTdAmwC17d5I35UACs
D4q2Mp3Zr+XjO4RMr2zai/2Ldfrf6QAV10pRHRwpGdVOCJFwbmaCbSj+l/0It3esHECwhI0/3xky
May+z/kYWEZUcH6Ru2kxaHPHbnCzzffd9nOb9vVJJ+S+vaeNzH9xb9Y2afGqUHo+HDZ10c66KF++
mKLX4/7944x4M8LmmcCDBXa1ljt6ZmYh1RgZiNU00BKJGeFtitutsPOyAgzrZrudO//oEMa/bvLQ
glW/GMq9jLSOBmhibM4C60tMWYTOc9Ff2wtRBO/RfdVUr1gJIYbFJlJ0SeUAunefj5qJQ11QqTr/
BMbwYOeErhRtsFsBikKPLdVlgDiIrhlALoyvx62yNskKYqV1ZU+gcGNFNsJCUsbF2WM2+7b+l36o
HqnwYWnYv6d0rWvIm8yznQA35yXQUaqfulbloEWHWbuM0jVs7tFRQNEj23Rg8sqPg4RRgNqbO1iW
pBlaGFJa2+6LQV6Eu917q4DTmqh+0d9/w2ez+NnZiou7bCx11r2+FVHxI4XVYIVL5w5BueUeSi7v
81ORYCkvn8vH3cC+1nCxm/UugNrDvaiMpoXbzG6h4ddLh3x+Q8i/wdi9IHnuWsJanY/0TAMZQOXG
/StGAbK6BsIzapTRCJnjnBGHIxwvH9TsC5uN4sJRiijuXF01CW2g2yEUIVgReQ509lo3WOjLrQXX
fRE8YX73YcQdGshX4ojZLUgytwBupQJ6hNglUOehe96MDbMbkSbWcPpep/eG22QBiMw935HBlLa4
W4wF8fKSN6U0Dr/valdxnRisrf7aRndRbVOEjH1G1Bg3MD+tEADFT8J3TDB1PdsEqs4Ip8muniHt
okLMZpwiL77jaeTbhVAMcY0eOX2zHSgtqgO+7RD+ni02jzQlHApVd0NLarls+eAC/FLRO4IgRjrs
KLGqT4Nk6CkyjebpI8Obx8AqQtbBdDE+CWqOy8tJF9EJ/sUe7O+dUNMdnSvG8kRRVeHV5OrVn14H
mmE7Vek/l0+48l4YhzuSZhah8pz78fGaijBq9uQX9mdEugFX8SDdF27PlDM+Y4o9usM0QbN+Lfmf
IW2pdfgaLzrqVt3Wu7nRAbvHSATeWNqgQ/moAP/MFgLEsLdyfhqRRX2JJnpVDxaesKPleCMPrMVp
NYxoONrmgqkDDg7HO7tZ0mBFNPFx/C71t5cWmNK2tEXGZKeAOTgTGhZivTVXMLZ6IcrDVRs4Q7NT
BiOUVxrEVWYpgSMAheBWriyb0kSQ9pJvStAp190B0Dv4IfBsTXnWODtKdW3NVCNPcf843cMd/w5d
duz4IWH42QP325Uz+nW/gx1uKDZjK9cEHE34STtXnrcoa6VerYVSZ3v38XQLfSKN8NgrStxmuvqK
jHxpJ9i9ECDphCsw/pyTw59V9xTYqxayDEbedMKqVwEh6JlXXlaW5BEjan7dqgT4nQ0ZLAYPWDFy
DmBWrM+lE+kjWihtJEbdcib/laGBrwoyzryaA5cUOXIYfOszLJsM74lRG0hrJ3pj8V9uGnNWRfWU
nor1CXH0IvwxdiT1/o7/tJqPG/JwBM3HgYiH8nERL8cfoU2sXH9nWPnchnb3kSzYS8PmwrkCrUaZ
bm5uArivYGjCXHKHTqBoEpxFCcbG0/3osv9vWEuCB8oWB7B2YTXr8ijAH8c/67Do41C2Bud4eYyo
QyR4HyaROaOdWCUCW3wDPJdMAisMq+9hih5U3rdRJ1AO9r6rHeU8fnUbfcEB7xP08eI19rT31o/W
kY8xOOKJuKTGamTPTiaRBO9L5eGhqx++S07eqSd9hjvMtvDR+5JKPrdXVCIo0tB2Y5uUGYpvVkqz
O1d44YJpFBf96ZjRJfe3f337y8IfdlZvfznUSakwB0RJGF7C70eV6ohH5h4g9kQEzsS90qaxFu2+
b0yaq9mLKolIv1cdDNyQJmxaaWn1nhuD7qY5JZgX4NB/jM7Ve58lcdpZ9fpr4+EejuaSA+ZK4mkb
5OxOCGyRrwKGrfrkq7nsZmNS/JaQdEdbqyJ4W0bHIAQsH4aJKW1gaMZ0wyVo6VSMdZYrvn7LRkzD
ThSiyqw7jjAQrnTtcCZnUNt4qHEjjaIPlzRQSuKntZhbfXAnSEn5/dia/GBrTC3qjwcqKrX9oHOQ
XtXqdjRXEm5M5Xe/DISMmfS85LcqxnL+xMpZOdZk0dLpAXVqgWqfgP9STUJdeGpibyQTrEmSVFQ8
+M3Sqm117ORfx2GuwACdDvyH7myCc9bQ/mK3Ic+dHsAnv237ZhBRtBq1RvsxSqu+W8FfT8xi5T0n
GGhTKfS+dirAq6gr3TjdOtQYUjzH2fKAN4O+X95nJZ7nxZf5JL/uNMnNVqukxdLJpu6gOlknPPRg
uMKi2mkcvzNG34ExSutfiviCTOHoBVXve+3htkrEGvXDuovu+hYoEPqw9SY/3fs6M3siHHWfZnkR
TAoQgbOtd8wSL2CIRvzSTjm5rmGCYbs/gueaoIjEeCdeS90Sml98Qt7+IbT04M5UtqQ+MQcJXztG
8PR58kFWXbOSEb1j1/e9QTHrb5mUDOaleDKgenT03MXLTwQaPSwf8V7vJwndF028mcQH8fJdpAEK
nGCjSPLLuhq3cF1WFXcrQcoJtdrzL1ry30OqmfF7MlCPgT46E4Dge10SmwRM+4hDAnxwbhwa1Tfr
ozf2FCwwP8v0Pdja5CPp46EBuXmLeYo+TGT95KK+AfLqVp3yXFXLVo2ro7RD4V+NkM8OQcAgnPWE
88tYmtQBZjELD6UqCynQxUp19Iel7XgwEzWEtaMZqWpC9scltL6YwpaFfxa1j+8+WT+B/GUvKRTL
OH7p40rSlMYGmVuWpYXN7GhbUU4QzQUnK6DIPKqSaA/sNtW6oFSkwwAfYn/7Axzqn9BYuX8L04qP
W+UaBl2DAD6byGAig5CYpsbPQ7EMqK6Y31A/1UxKWulws3MO8TnFkLEDrYttw2DVgS7CKvHksapZ
EuIof0dAa9aeXYZ0hpqWO69MdmziKnMTrhQWe839KCjhsqeasS/kJfFy1y8RHPq2Nze8V/hri8SI
5tVQKjWrV/X98CGjtoJs/+AJ2HCOXNfk+I/w4vLgZEoLcnStXYPdr7yXEiHgC66t8AhPrbqfsH2T
POaTKNpq9gYNf4/84OCU290ozZkKSy58PPQadVRW22KLjLm72Z5ggQEVh2af4Zz6vZJk244ZFUh2
3S6+EIfXrzQOb6hnttqe8SM/nANOcstdxVAItqfKeM4eEn+bwdJ0sVkOU3szOiT/106k3flrEWj/
xaZfNatZ1NDHHVvFKoFqVQfdr1SsQeem01HcHoyouOE8ir8nHPlFvv10pXxNl+l6fndbUCML4RxC
gL2u3f13+ZZ3uh1KpiqbumjmGH8R/VHAy/hckF5BKg7nWmycU2E0rtrwFEjDWjsAxhBuy95th4fA
GBPKjZfOgd5HwZATjSlhzF/tWH/Mpbao5wte/eTTzb4j0o90Le2vFCt3TZXbwJ5gAZ4338HkhRmJ
waArgaSPYSCpbSh2uR4ebG9k6PMIoOQ0da7QIjlXSA8I52W7luxfVDJAb8BCjYhJ0WDy6qMIPRPV
2Y3MOnBNMOlwAv+evxJKM96c/YUWPzJj5eUf/elDC1N9CoiZl51xBD8w4wNuWZA5b/apjzdDCk9a
HDwwLeObXOlfuONIPh0gUw2xBCgV91/j90H6dTc2izUimcCC52EFQTkUZx2lx7AM4x0/6YWcBJMA
w5f/XnCWqingCTF3vaPAzXtGQs1gMzNVX6PCypRpWOcYBls7HOYRJlkmI+tt8gK6nVLcHE6szWBh
zeJGN1Ro5vIM5+VNm8dIByBoPQZCWyP/MuVICwR1JNe9/EMHX/CBDtmEkX42wo7hS/dZ/Q/HUDGZ
6KwrAR724sj0pOrzJmSJXFdJwuyQc0RjwSYfSpApj1HXf8h7HfvMFMN7if4+bw1Zy7Dxs2nQoyEL
ZOlOkc2HpCqk4DV44/NsOsqWFuLSlpAupMOkiVECrAYhiCjxKJ2BNC/xPv51nM2EeYC6qV6COM+e
GGbPvyVrKQATcBKLv4XiCkhMX5Z33AIITWYKX/fuWvY7JY3V2S6TQLY9JXH5XjZ/2VZNF9Q4OVVL
HwQ0ZCr5Rv0c80jSJ3XU1UATU5U04cpYQciG9eIc4Ii2cGZDdH6DQtS2tPLuwT+ra99abw8OXGDR
Y1wnmGPyx0asvNfE9mpjGoMrr5ProjwmkAiBkeUY32XKhLKkL7jubtiJuKyPEJ78kx9ktMir9/kV
9CSKePyQIxgi9lsOnWgKvH7H3ICE5iIG0o/bAwDuvGZal3Trcdxd9k0WmMiH/wthI4PAqyHwveG5
SouxEiEtUGqXVGh+nb699bzRw/JTcfsbiTGLohp2IVTFMauOxPf1zh///OMQq3eL3DQAAs683pxp
/u0cdjJY+Og/pAtAb4cWVWO2DMbsW4g7/AUjHVhwdErF//nE3V+HfrrcT5uAUvIRy8P8DUO1r3vs
dJu3RsjTp4TK3OD5OzRKhv6/cnfGArfLVZ3EqmbNCOcH9I2mk/cdZXP1Pfh2295a1AfF5LR/jnY2
v9MemZQkC3aL6vQ+Lb0R5qZMhpbI2Yvu5Jl2HSp979cPR29GNeug7G5F989bylMfd9L3ng/r4+HC
ZRBb3FdNic7nqch3a2B5g1OG5cGKpwFwFWljxofi7pcV+R95erHohzDO6FpcCdGSKXSVaFQvh9Db
hrtzYrQ20U6/Hdz8WnVEg5ShA+q3LW1JhBpX7ySV0TMPmYuZNZVZGN/8Gsq9csNTIF/Z3iTSlArj
5EaUeWHtwOzZVRAHkQB8DP1sUtEQskdIQ74shmiX/WxbpynrMG9K8P3TrL6UiPTv7pC0NhLUv1qh
oq+cuhIbtDqA9+clCbE2R45dV/HcBfbK3HqCy9Eh8UiVi1EYh9Z2377oDa316qCUQG2vCkAnrF7v
urE15mO++yfJ9Fq603RmK9+TMj2T2U+3gXo7dy95zUhrJ0FJQqDaBFlvw0gyJvvPey/Grt1xMj6R
E742dQfkQOse/jpcPDwjPXCafCYiXO/+yyfsF86hojVYCKhE6mwoqIgofpgHN7b2wsNimpwYO96C
mLd2YKCV+lK/Bpz+bxCTfdCpGEf1lJPryoTA0hDKEyogQ23JdA34iR5gXpa7EeXv9Tgd6zXFD0iw
ovhjHSuu+LgRzoQgtaeSgT0VJGmgfyLJAXKJUaof+kcGSREeqtAQKOa/UTw9OyHfYpQ8Z3+x5iBE
8h3/GzaotFi7J9VC8UaV/og7YZfm/bOyJNjoTPg+ptkoDQ6NjpHpFn+oSTnEq+b71eZpyGRHp6m2
rIEPE/KH5QFykmy5O6hjnpNBTe7TAoQS5gZPSLwTGHg1H4GDIcBIdeGuAVmjIqwK04quis78dIdf
wZwhBE08bab5lf3GZX6YH/Cy2s+l9s9JjKodqbA0uT4cItX8K9T5BLs8FO7BkZ22mk2vKxvOtM20
61EIXDQAjarRtlTDpFVGb//B+bE0XZl0QSjKDukaCQKqOGxWRSPUnv82n+yrHdJIu+PBe/vm4xtH
tgh45gyI7YT7y7xZys2WKvGDZpwm5UR2UWgI6v/U/uC6RV931Mtyjl9QfoIP2osvKIQk8XOpXckz
8RpJg45XO68XFGqndhAfPxeYuinon+mD4GsJ3v3z7qjGfZ+4kZMKO1LH+UGyadZ4rQFEd8N/pf+k
lbWfUQVeCyjJ/uTWrk1T/tZFJjttsjZxWwpfmJqBuWshJHM818lB60Fu12bheI7vqwTzilrbY9LS
xDylKnBh7/fgK3hJpZ5ivEvJYSqF+7Irct3iL0ZZXt75OIs4OgualoDMNzie0Kh4LG40XNhoe5zg
EAce47NwOVIliVLEh1ZtKh61AfebKdnZaH3fyveXwIzGvc/O4ui6oDCJI7LVlTGciKm3XB1T/rBO
OEdlEWZ6d8AbUePx13uywW1WQUoa9csy5rGRu8rihYbvYIzth7r1EO1PwCI+NvMYFiOKDgqlULa9
HaWkOwFZkloNkJ15dE20JGSkcic0tUuP1TApJKd/+BkLbYg8p8/juprdM57XtR6heow+B/RC+c+m
g6tF27S63V347HALxS02SYP/nv4NDQy9QCqMCqhy59hlOAJRFqBbZxEKai+iUa4feNeqHqgjPsUj
q0mwRcrw2RSL6EeZF/tD6pZ62oMi4OsaarEH/cBjcxR+Ef5Tpm5AE11LYBm6wpiCQVM9a6MWhk5t
eon5warHEJkcRMhlRnnJgIThljv23wDdI+u3ltEiuolESLr22+PS3nxROS9fIaerdBh58Uv7tAAg
gPZLBoVNVTF7hML7i6txbTjlWQVpBHtQLyNXhYH5YS9kTYoJ0NX5uxwmM7mxbz+w3i0sYTaai7yS
ZV5MotRruIklmslgE3GJFSu/2VsW+aR75Dabf2zD59BP2l8IFGOP1Dt1s3SgUjV4NaYZ3olbSg85
p++UIOYHNmumT3ZR4I1hmAJAyecRe9ObxcKkQP/YC2/RA1g8CNs9A4M6noO3jareqHqzGTkfHuoh
3+O8vvkVfw11VvguZaV1MJOGRPw0oUI+04TDah2vDHwsD1QwxvbJjEBEtAjLSO73TugsnfshVy8O
bCss4tt9VDI8MDFWZStZrbMzMz7pANQWUI631NqdZcgfn8V95N4/Q6tdQw8oYpubvcmByeQEMol1
XUa5NAKS1guVYW4FycV/THxfC9IE9cfsY2m8KBD8Pcil7nMWSU0T1oOObJreimbC7ygWnOnkfe7j
TTTAICBpq0ZAZWPj1+3d7PdgYYkZCgjJcnpuywHpIm/JUBIkpU7m4nXYVtaYMd4pum7oZqI8bIYk
LH01tZQHwcApr7vbWxH6d3IGEVbVi3B7GxzxzEvccEC2GrTm3F/h8Y15Q5YESotXwrEDMbWcH56D
66i8YKYh0I8X2piymvc8ffdz1pM4kjcjHBt/yljDOp9VNWpycymPLHM3xnP+u+0Cijh+YiBY3jy4
yYAsCA06KJKKn14jqIZNyYe5SlKknOVKFLczAkaePVBwtLzQCsA8BlVN14BGqBKwVUfR4yplgqy6
CMkCv26He/iXqiOkEzkco80DMKqF7iA1IZi98eYwMPKhylBbWWWknS3Xbufjpk9k/XDCgRZnSQou
WjffWReSY6WOlYVPNIvmUrUB3xXDdUFHPzO03fv01QsQyllC5NNlRbFGN+8znoEtDyph0Ohgn5Ij
Tvc2h1Coa3eLvcjOvrxjYQfY0OouxDSaVv4+KVRHN1A1eJRKyFRQr+mcyF47yXpdeeEbX979ptfi
38KXl7YUyZo2Hq3/GcIqaw2FT/FMoQ40bKmGf0RLj7PP8lKqnQ6mUuL5DLIm8TSJkexl7utkpzc5
B1EaXhxIQzrWflA1J2EC/DQVGGepmDGhIx+h0JNOkmQvuQc7OTs/vXjhaAqLPp21VcsGqr5pY0E0
e+KkBVIqPYSFYh2G/UC2ITCU1iVximKstgJmojRdwgBkNmw0j6WE9n+aKQCDeGYBSsTawYKof6dl
fLl4eMcSzsUNvER6BL09YutU2E7lNHcyWC9n5uvbvjw80g5wXaCS50Gn+4w48KVS1IrYakRtPydX
xns83m5TtbZ48VaPlgox+r/EPqmRJtlR6bFUvu5pbPkRY5C4t8iDFfmW8on4XjrRY4oaMQRU3S93
kYdHZbyDDLx3V5YsXhcke3i5/ElHfjVgH+Ld8lYgDBkoXu+nJZ+gGr5aYis1eTJUaGEE89/zTLMZ
OOUWu6kEKhWZjaXQnM0A80PlKQybAfYq4z2EZkC4C4Xm5idBMi+cB8HfH7xwNgPi11AGJxQf5uiy
4xDk/kZpnKJ5DUEwhIPLhss8JcjudGTHUzeMvEAyacF0f7J48RWhZA49u+g2+6Wpsf9v9mai9+V4
ZtCzoLDJK4wbSjYsxfcz7coH82dkHnwL76iXcvdhkexE4Bs56XXOeHO7Q1hhABXcsqXI5C5EX3Nz
kL7dI8oyWAKK4H5lb0NZeoBls2IHCYhL0fwhcGQDomS/6MtcEY/VW0+I2ItgQKS23vCPQVTgbcwQ
YRmFH9zDE5L5aX25Ur1UaAYiVlt9hLBv4bbuHkh59liUrEBSSrW0tTBUQcxS/cRJEVwe3HM/6U+e
Q+W34XHjMUZJbM1Bio0hClwWe6pW3D4RNgkHgq39sJPUjA4krjdCOMVOKvqvaXIDUmzWSTrRUYFc
uXPZYtM/JJ7qgH8FSlpmn5fR6wASO/zUGNtN71jH7C3OJJ/XMFi+knYx/g1SKf8zkGYE8E+nabDf
Q0/xqIizKGI/xh/f2u+ZLGhGb+//qKVQ7Sl4viju2wZ8dta8RDmAEAE4KdEXCgCcdSi7vZcreOhT
5FPuhtfI0Os4HJ1NUP2yNj69Tn87/abzuwxA4xKNuAXmq5/zDnSjVOFD+pIuLRmKFLm/Vk+aE76h
JRwvEDu7BSBbwUVVZLFBmCuj2pH7VRWRTPybnf+9fW5vHnUdI9ffA9//PfyWTti6fgRd7zBjyt3T
LmaWV1RhHcttFZVEpZsUeqIeF2fVe9ZZVLRpwxw/Jn18AoRu5pSoF/2ivVCZa7mBrxj0ATYgCOva
acYZcQB+GP8NPK0DeVIw5PyuWw5RBAdR7UKB0NcAhN1erxV/UNhndyCqG7WMPpoRlww4rAIu5clp
6yhrpXwKgSgro9GxHRHUh1jcCFATqmpG3vfijWevUvaJrCk/xi3LoXY98UuuJ9qrH9TznT1NsCbU
d4/4PWftP4KZMe8tf8DPS2orw/P+O+NwNsEIOZXSpnJfzMC90TZJwUonjooVfHAI5pWyhAHpLMXa
kt/qvfHUvbE8riBCyArB1EDAcdkKnE1tPkrkyGuD3R2DYDljBkbf7qg6KUVE45V1AUFjdhe5LzHU
Lh07nwNrfuHQKu0BqePs8z7KPwdIGQt9qK2y8P7/PAnOjEYYdPQMxXSyq6z/6Zrncc+Uk0+gGkvp
xqxsLZKo0nL82Bh20Hq8y7e+wg6eeKb0LsmnByCeY4XHqvWaXzcgzKBJrMVNA4Xy0idvkMVpd8w4
sH29r866icYAaVTtuXxBs0QmhZazfPeevv07vQNUOnTkefS+idqkWFPKeRKIrkRIwTITMJUNMq06
291tbLZoSdPXElds69BaiPNhghbcFZS+3ipDgw3AAtn2h8idgQFWBPtsBbOeswxmTb9UOO01QuR6
vqb3uNL9Py5wfwQ1ASPNFwjW3yeKwRvBozPeIO82rzaR/WYIahW1xStg/7YNF7GvNywnoGEiMr4H
mRAIOSvx6dJra7vs4G747dR83Vy/JM5iDLVGN56HXo6wt9gBy4FgGnbej+7iCyG/brOBkJEQLBDq
d51KDoauIxiVO1Hh62ebqxlqdKDQ6lyGSJEGGvbajp0gOiUlZtoG+QDc90+a1cotRTrDNSKTKLZc
ROhGYMGgFkmeW61AN5kaUvL/WnVt+lcWsvyMCLacdr7rEtTAGhYFUa5HeT0EiwTVfzDbkGnE/TyB
9pgumK/4vURGy5HEMna4iZhFuWJ3Ay1qjRPuvoLkbWLTSc//TZY9v0MwAslBhaxUFVQ5P2jWc5Og
YqprPy0L7tB8ARXELirHOYtWuZN5dwc/ghGAEJ1Ky38DPDoGl02GlX2M2p/AZQegzT2R5CFv0lwI
FARqJg5zg8H8Nsn6TqYBLEjL3RVrPqNCe+jt5eD9IP1cYgY1+vlQlafaZ4EippwuaLPMPN2NE+5G
dAaftivoOOl3gM30+0xJVUPnLKNxB0DTiDpXa8Pwj2gG04J27uPe01T/w1lvYNE7J0aiGbbqC6MN
fciTe79TiDalfh4Y7tvLxFK7C7Hk4/q4gq9vANzh2CiTevn3ppbQFr9BQgnkb8Pb3+RFONHKrfLp
wxyuf6/tOjboSbtQ9lOhXomSrgxPNfU9hwaihmLb6XR0Qhn8k0qlMTTnsUEBGbXsRS2CkvMjwCQ1
bYhXszznnxio5L7Hti2oSHYtRbvUvwS2bHi5/ULIWs7qMP3rL6/GKU58Rk1gHAL9sRKM+Cl/js2d
0nH2MIdy466uaAvR3hSJ++Ko5HFcSFTrVJcROnpZUM+XpMdSVz2hTLT8FxRwga5SxEYx2Q1T069e
Izu6xeVhKTS7IfbFMSQOJdf4Ksj/qBpBF0PfK7ZTBxzKw608M6pRDE70NntVElqI5do8hnuyq/8X
doMjW+uAzsZsbaTcAJTuhFy92srTAG+tDP5is9FbFpaEIm6Phnp1m5jtawwvn1dSj/NjIgTF1s7+
oyiEP/nRppBnfwlaJQirIJoiIlowt7slF3OS6CUyAx0+i6QVvbxkzax9Dvu72y+HQH4AhnpITeKu
3nUDhGw+9Q6xJbdOYS60RXxZtJaQTWMpbP7oqC2c0Hngi9RKOftwHUgTrsdaZRABWorrrx4TwAfz
wLxhQPK4RhkdOgDYY5psSsdaysP1hqqgZ0PgzECpwYvOLVTGGuYFgxaXmoRd7AAlRfKsLVCbrpao
zUx2LAsv2qMKK6CapcRJ2hlpZkgW1LhKY/Zjly78KPBhCTyx2WRRjySEGp4tSdMhwqDs4s6FESuE
MRj/t3qm6MliHe3xYGFhpuhd7dT5Xsq9Lky3+VM1Hn5Ls8rMKcmy0Q2N/Jkz6xvZsRef4bwZgE2k
uVLdTXt+UZnsZvp2Uvteu1AumsK/XpE5uovwFSg89eRKcTTQhMDpeI2bfmZ7karsJYXbuQV44qqX
sWGW6jly1CZo14GK13nPGh+XL4cBo2MsOhQuK4U0d3GUQRb8gKjXTNyQBCvPa61DSzjlnCW5a5zQ
nPoVoNkvig+V05GM4Fo8m8h9Ygvzot9EHRWuFqMA6Oca2LqERUXsnb65Mw790H82Y3hcO/FS2qFJ
71c5lupvCAOV3oGceaFLg8Zp3tk9WPx3Dkd9gPPbxw8YhlYhv3nVx2VtDJ+bFkAM1dC87AHjgRxm
99cVklGIWDP44e4zoGUtq59AYnXHtGC5JRr4Bq+1uKa13oUqsN3EbOL7vBDMu4xzEG6ivImoUcJg
WhB6u22DDu9MXEKUFcgprI5nLRT8gxcJE7eXMoY+JQ5hETG2NK/DxzTlRIlEwQKIn/CJEqObYAtV
ptdFzHGZMg1C4OJonpW2OUUTGjuYYK2anh/ELs9lehHWK6G0sYS+/8OvggerVw20l9ixnjio/8QZ
D8GneGiEunCuUpijca9nFD3Tpp8FeXy98aDnUnjCcVjkEwTcnQeT7N5Qk7URrghxCu5VTxVwSIki
7PBzgWUT2LMnjtbW4jRNamZZx2cyquoRf8ES82sSOeCqtalUKvXxSmD1d6w8KOTY+9LuHsrr+szF
C6XEIkk6ns4ixCEjT+AqG4NGG9/W7Giinr1O3h8xq7UOf/45gR1Ur2wpjd+FVQ0k1OCUN78t17Zp
UEKYOdxRv0DLuB/uKq/AIwJrTM0acHibNAaKimn10NsJ6TsPLzemhVCiUxYmZ1qxhxdiievXKNEY
Opf1TBOgAMzkHyoyWqBKF5i4D2VXEEM4t9SmIH+1eoJgUdhUPm7WeGsWKp0kGkLIpWLx8tvBLU9N
X8+JiaXZDZ34m0nD4TVFXY5unb9IfRvxh9W9YiloTNdER0PfpDwPd2rZteTeIDdqekFFUZPLOzlN
KxRnsXAN1mSaa4/9P5co7T9LbVPwGkprzqgMMj4ZqPjYbMZcmjbGjZiqzCARnqa6sqKQa489fgpx
8/AfCGDd6f8h93lOfQeQUeFtgM0CsShYrOjZKuEDj2FrHustUk0eZSzeVAZoflA88bunM4Mmv+Cy
AbZxjYs1JmiBdFrSTT5dlu0s8ui1Z/oOZQVhYgkCSRZ9D9a2cPQ7XllvR8VLcTAfUpGxcQV62TDb
IoaEJqUjOAA3xGMNy0WMQyDZeYjZ8Fc/f1ffeWiAqbHbOqofP/Xeb/8Lv2ZCAe6opBsI9ZEbtTiM
/fp3ecxqLLFLtNr1Juz3/JMA3OT9YSWbrne5PmpESwAwDc5h6t+fU0YJs5eyyL8XCi0VW6c2KsQ8
rkgWBr9pZaEcoKQ7P9B/4Gh2EthUPs5mgVE3MckwdoDEGqGdLEdEOVsPcNmjMtVMysRf2ctICYid
WdJXGiwdhNkvZdP9LVJRRWzjSGzNvRf6NinXOtLD/RHKTY3TDCit2FC42H5KES4WXzueG0RdU9XP
eqhTbjJj9h9BB9m6VUb6w127Ih3anHEZiqTmqKAjttqq3teSa+nyi/myFQqsedlLTeS+PrZx5f9m
O65o8/yf5BYjCSpXaRoEkNX+sHJlOUFOjW+FswYYaVV9peY45n/V1WduadhNa3aHf50C90Zz3O/h
AoGlshu9GiuV/VgV+GbaTJkXB7XO9vGsi3FoMKNmS49opEZeM9+2pH/ROSBTfH1YhRRRo3t57pea
GuY+hsKekQY3644oEhkFAKZmVN2u34ZlMsf4uKGHVVBAb3OHIf9J53nvSzPGtrgIT1axZME2Azdz
/ckKrIXAuk+G4gQJifNhCp4chfaolcINi6TMBIScBQULJzgbNzvkAOjG3mFLO7fd/rwKEULsFJ16
A1uyJXIJwvGMmkzJ+0yl+Rh6j+Uttme5E9N1Olqr7OD9kgeSBLcOI0RKDAvu4IqtFV+EAlZDcIrr
QEOvKSShyqWGlkV2YkD9TMlgQYTArsV2KVogrRz+ZOJDZQwNgM6D5W8OGAY3l/eyup/m3Beasb62
atiPPNklOXbzh0wr7+N4a+bhoY745OZ3P3JuVnWxra64Vnob3Cq2tZo04uj9ECxenKE9hUjb9i/3
0/gc/9BD9TGPB0X9U6WqA4rOcpyKIZ3iOLEhNIVvZ6FvlgVXMPRZY+3cciTlvgAtGvCZqodmMsnj
hnwjo9YcMkwM4qIq7hHXpRT3B5VEfAA3dxCqNfr/a3AMjQ+3wlIUZqTn47GlysWilUmaVLLEMq6X
dKDMg71fg5DlLmVZoEpHUhIxdn0XGiyY2EUU2bib3z8n+dg2Fyx+mnLVsJoW1HCRokd3LBbeHMQD
wwUagHHeLqw4CLU4G9Fsp0evpwjnnvcO3zwj4O/Nnfi4KmfbJmqvsYw0yMYtlFrvgO7J2GYQqUcG
HczWVgFbw+dtcm00/vuDNpz33p48P5HU/1PYpPYNSuxIZPxzwh9LRmHIJwPyk2Qcx1NJoYUs2oyd
qU8GsA9EaQwoCs6cWk94YIttZaSgMNWeXsQ1ZfnBV0i6yfNqdf37CkzcLudXNRiAoI1NbuaNXOVE
5JcnDgSqIio15AijWCvcljleX/65N67neJKltzUo7B4dRJB4ki903KSxjnZU8eQeau/8Z0yi0qqE
mUBfG5QoZ0LShPoZLaK36wCT1Ao5Zk6HF7E2vRjXT12vXtStzYzjO1teqnPlF6zTzIxOz3D0z6p2
cAVaGtL1qRcGGQk+d6iJ93zKXzD6EnT5Gb9GHkCXWoFL/SfXTwL4CMiiP2vdn1j8vKunsKBWaa+e
nyqxvd11exMSw48Y9kegjhL737Un4rApgfELE2A/qzDOsbr5BMpTNMYxzxLmOnGzHGqcIuyGulxf
1yQzjtkQlCiGca80uMrdUWibG3G012A5xSfNv78CLgdWfIW6qCocv9kQFPUpp79BOHelZ+ZzTVm/
FhiSuYCvmP6yiOeLSC4PseTdXb9lwghhyukMO8EZg5thbhoUXvCVelWxRnCkf7i9lrh3pDCcW5BX
mvyagCipbhKzSxRky3A/MrJU7p+u6l/NERvLEBq4m492mOTb8Gf9SW66UB9o0PWbcfyEKs05DQ8Q
/X9RSHFF19VVkxi+JZ5D1T3G7I3cPgekC+D+n5UB9NfnBqJrAqMDv6QiKPD0CE8oRafMqENa+QQR
Hq9wplwruR0ScxDLW4CfnBukgfW/CYtJKi5eP4UZN6N3+1jtCCBQ+bigRTz2oB2KxGyWzSB/MLfi
DilHTkJOrVS9USd7G46ifLV99OCAMzKhc+rwH/Hecb5khB/u/qX1wgMIljZ4ri4iyKrBFGaIzm/G
wiPugRcyCWDbNl3hGKy4A/+SwXtP5kWhUh/9Zg6CTkofxXFSUtN21mpKErTH8kEL7DjslgB1eLQ2
+jE6XG+1YA7EEa+yGaL171XZMIQ8u0S88MMltLk/b9e7cnu+c2zrS2p8jj0JF2TKlq/yahrSrogj
zYkZZTVHYuVbuaT/whhZNE5Pi7XlnexnC35lux8v+sfKtoQkzceePiCXC6jY5F+S6N1YzuWZj9Uf
djs9ePXSPtPXfru6xSqHmmvFOLEBtRgk0tT6XIiy4aoZwY5x2I5tSkJ2BQUPwU2PmdFDsMKs8ufC
VOYBDvb1MIwyxZ8MlXDTFIiNn2kZ2s32jzHfS+uc+rvvUBXvFjGKQaH0kZn+ol44v8ziMsbJLIRT
0ViEFeE3UZ/mOTatmvKRunxPbZgo9qNwQ5Z/bSxyXWtyEGa1unX9YL5K7bUrXU8UKz0Zwd/ns6gy
1hlqORUDdTtfg9xMZ/iZl11iPiwxsuX/ptUbgjpeXPqmwta6GDc9cvxmCnzSOQGEyAC/ity+bZbu
hwp8mbMbdjKRfc3ckJjXmPjKgf/rl2Jlm+jGzi3JTklfxrgKgvchg4ewh4hezZgsQj4fNWPIysWD
Gp4WQKaYGn8hOHeRwrH/g5sr+8It0YsmxfiewcO9I2PJNlZC5cDqdIkXUG/g85yuiS01nN+7yyxt
GAk0PnaFAxiQlP640ZOhQmj/EPMwPKGzqK9qHoDMB6PBPpV3PFGyV6ngLVbRji8qWhzwZ8IUtw0k
RCHGGXMS3OjrW2nS9SF1SBgWz+Zh0Ty7yZLEFexLoJnDCH6Ej6YecxGL+nIBhhC7vxkTotn4XbZd
RwB7c+9JSD6NppTFloVe0Tnog6XpRPRkcyn1OddiQjt8CfgAqldJIAcVLIdG3xkfJD0ht0Nsrrgz
mthfkfe1UUt1SDDiYZGjdsUgrgFTWccPQTkruKDsS6o541/3ctqGL4axuqMDU6DTxpcQS5V6mwsd
BdU5DkT8E2CP3jlGUig/rGmpqLZ5j3BLlxf1ZKZeSASsdJ+ZeE4HPAnESzyTqtdS/oGCJFtrTMoq
/MMbZ/HPCiwLTex67JO990RTHYnw1zM5j8/hFMpzQIutPPRDkm5w57CzX8+fD6PxBKDWCK75s91J
KPAZVM08KaT2S4gP8H0P9dnwWQ1ujICQo8Rxty8crA6a12LRG9ThikLC35LUTKxI3DqKcM5z6USz
notOvrvXMzlO8jiOcyEV6vx6KuGJQMvkWx7NcQaGdWW3tyRB0fJbulTQc28BJVFyTU0T55CqkVE9
6lOSgen4Poq18jdVW+ulBlSSMbRCvwOS+2UscnnVwUkyP9yaWEx0bI5uNH9pQxnq0woCmZIb9l/x
rlzdKS60dg+/2aRvzT5ChRjhR8KWsGqPS5AXO2g2owDh5xmhb2rYV80Blh950JM58nEMMocAUfzy
hzY4sySewK1OQPEVnmkSCB5ZjM2Ja8GvocaB/6jniTRLRA9Bf89ydkDbbz49daM1LNFVh58GhDpg
nxidaNf2XYq/R+FXdjuyj1OSgQTmiIv2YJcMHvfhuW5MRoSeHhUlvTgJyqlTHpIk/AhJdouqQ/pZ
/5E8T7YNz+9+u6cAHkUvq4LkK01+MLSOBMePNL1zYCKQjrgS3FJoeJKwUK26cokHbYQZw2Tdtg8A
99O8NRytZXn9oCpIfXLCutb+NnzNZhfh4NlsWs4s31Msvbaj1gNVscdGliNac0v0WWC3K7+rbLkp
llM0hafxxsLo5xCbAHMCqbxJhUnEHEqODFyNKMpLUWSAOGx/3ZTDopA2ETRPmb1w3/6QerHBp1v/
COgpX5AYYyrCd5Jyhp5D5Ma0JkZsaCnN9ZnT2GGSpxCSOSvYDsGGGi1gnMOdWvHcF+4i1gijJmVY
mw8HmRoaRNA1aXwN0ePBkGnkvFWfJ+w90+nk/kkJ/JYLHZWDmZK7fJZK9m09rvoi7Vcl5VocRb1n
eLutbxtOIl4/Hjfknwuw+rJDVUhWzuBo5X72dAvuiFILUoCpKyX4eDF4XNpH0jkX+2s6dj+Qcgam
a3Iw2chYb076w6cimSjrHRd6HxwNPNKwi3/qsYPJBNIwHv8Ci/Kz4OjnBrGim9LBAHpRLExv8wPc
K1hDZTHgtSPi7ejd7agILpLsvIwUPQyVWKqv/mQMCS6JuEZ3D+JuNatykUDOr/tfqAMh7v0742Sy
8DwoTkkuEBJNcXp/69FRlBn4a3a6Se/ZY72i+1+KInXnnIgvJWIPh8gLNr73vliinXcEBulo+nkr
EA9OYgpOk+GFe11MMeKwBmuJWy/6y2A4PWv/N7YDOPFNaE9dqRETzC1p1kb9bdPsIX5VRY54Cxy3
IO+cqQlUrBNsfm5AAWJFHyfHkGf9xa3tjcD8cRQcuOiDzrQrhfOXc5W8A/MO6mCHjKW9ihg3epL6
wcjhEIu2CWqtb7jCyQqM9tWHzLwuvwb7tIBzL3IVRqfWaTplmaW0HHNX49A9VTpCkqK2LmOpRzVI
4r91wQr2tQBSqaux6Nsj1Yf9FLnJTK8AEkvn7SyNOyJYIofb70yb1SdtkSjKgSTbo3ftpIDGlTVp
4X5Gk1hN8QPssgVch/wshJhqn+HyYVFGaDdzYCMrBvsFL1NCX+Ba24ng4JNnFn313ezpo1JErilN
V1fRHJAlbCtxnVgk49Qd7hgpvcfioNHOOSM90CHbN5LBlUkl95ttoREbDttMOeaCA+2YxizUo8dh
MU//FYFBE3yi0+d4VHIKTHPjvvoUwVRZBSjUa4RprqiXoez8ORoW+reIumklQyc6Qd8eW+micTeM
Zh1gF8HD5vKzOKL5vVIPGd5cmnzVhWXJ0lVXhu6w/ARu8eFQp3Jzv6x8zLyhDqiEgvFZsL4IJe+M
A9Uft+zSlSeeW6O5JLIiEoGIJI/cAUAwi1OJiKQa77rhrOZz7RfXoTn6mq/dKJa10lwJiTI76Kjj
t6A99iZyqXpBfWUrxdxzOEfIDnZV6yRIydC8lJupn3D1QBLmeDpu1omIigvp7cP9jX9NgfG2W8uS
ryCuBt9AWBC4S4jUG5VQY/EJbie2wq/jhd2u/r1ShgCjB4vzLcB1UlRqXLVezuQH3dlErTeizDNn
hyUr64t1alVJZE74yjG/+XeXY90xc21sP3dEVuRX3y/zHc/USFdb7nD2aVIWaU3zoJjHa2uAZxWV
whkP6Sb8e/XXAvyp/1X/6UWXK0zpfHbTJMNiaxKwPA/DpDIz2VwMbBu6LQn3u2gJ4qTArYeOR2R+
DDw9Nie554RQp9zNvQtU5+PSFYOtmzjbhG8OjrFxetZFh1rYhaD/QBVumObbxjAuGEZcupJCZ/Fc
L2eA4LwaO+9UIQ/HlTZbb+AiBVj9/7/2tur/JNbgH8l+4YLmX53n+feoVJX9wTGu75bZ2lDMoBKY
iTK/3QvrTR2fvGsCB4DfByClvETVWDIwE7IBHTZd0g9fUMmC9omHTdRT7+BZixt+7AnwG/yj1iPC
yLp1jk4d8M2+TXf3daLVm4bQMiBXOWaR8MsZ4CUdiJG01sqYW91zq04TcUX4G3FsYw9ovCTULNh7
bXGuRVNU77XC23ZgVJSd/t8ZuT/hGLSqpyYi9bwX+xLauR6bbL+XWOIySg29TS7KSAjtUaAPUVXm
9i4gaAVsT2qsdqPR340cJm405g1lgxzqpCrXhAgk07r3lWGTcnnY5zZnDY402O9R7tdPXLlJPqau
kthFE8dPHDQK3hQNPehSW4iNonklDfaINh8pQDSdrC9FtQVPtCyJakdx0f4hB6R4iQBdBcnO2vLl
MIeKVDYyvqnJEu/WzEPJfDPr0TRv65TrbBc+wsROKilwI7oudZ8Zz3T7BsC7reywB1TFlVb87Akb
gVd9wiEMco1pY0ieMEFjj4ng3l0HK9AVfdSDPFftj3qvNZT8N9Cw8PNa5PX64BA+F38M1FCHPHm2
9sZQKRxlEOlKfe2i21Buhyxs18MiOBgYkAdCuWzW3jQkdnvin8WZazJD/TIM5orFwjmfB1zFBlMk
nknzVWaw+QAbo0C6H1U/xlGNzjbWkrcAccKtFySIUd9UgIFViVJGmT121Vi9kXOHjKf6xXJO/ekP
eTQ4zIYjtaFuPKFUVDZFFTHkJgvZ2C2s6jAl8ivtxXLcj1KLioyyHntqWOk/ST72M+ksPhk7/yrm
dYtzTh5k8MSapB/RbduaR6gztE7/meSomApcoJFoa9l6Q3t4tEemyhgx3TAfGIvgJ6KevBJHvEyL
3delynUgRpu+n1GgZGk4eKzryNmY0tI7Q6F88kFBG/GxipRio885gC0Cs6FHNpW4SZeaA6hi3Tqq
fZJs3wVzZ/4Kf84oO2i6TGILVvWFypWfGT/MCJW1FhVczWrZGNfHHZ/PkiCThNNWtQN+OT1OJu5F
udZLfh1fbJOctXsqu5ZwPOlpKPLxCm/ktGs47hqBPfx8UtEpg1O4JN87IVeRY2DkAsyMVASE4RFD
thFYi7/5b6vkXKusFiuws9RqRBBYMmhhM0sJs6eMoC5fSFYfI2f4tG3ZZudYoqmzR6+D9+kSSL8K
9Ylc70qlQPzEr/F/kB/ERIZ6KeWD9M6OPAcH3TDBhcS5cdQotL7zM3WtLA9aEyPRlFhcGfztRro+
FokihLPtTCDWEbgxjC6p0GQ3piukMaHn/ERCpIVRDqmpS6+J1YPSrGt2kxiGhXwL9SLWrBWaTURf
yN6W4D3ki7rIoF83XIYm2GFpuwIuz3KAIJ6/vXnqyzNp+M62QqRP9yy5FCOI0/kRz5jcKa5rFsB3
TN2tVlZihG/4MoLTpYDf76ToXyJv7w9vlUZfU4ep+L6Ph0xFMT+o+67iTdapO81evXJ85ZilKSVL
+KUxPa6kb8kzPTMMg0XMwoPMhgJaBRfNijWKOEdhdmdu41dSsl24eejlU47rbZm28o0B7lgU4WCj
o0JKpzStFs7uzwvu8CzHmxTonMgH2uSdZMMfy4Tm1J6kVTNfpqXz64EwhWGdXIvRS/EnDrBX3eNY
JVmgd60tpnaQNX3VftacLifBU9dvFNQYayb5o1+whQJo9VVOXYlAYRXkLw4H6tiJ34YuYg8YlYbZ
FK2+t3U1La8ti4156BUPo7ITCinxTKL6ti4lVVn4Rht8St0KzhPOIL/6a3V+8yywct71ip8kN4+i
XfTHE8+0Geg6yZAmQJDHzU/NzRg2l+7sy1DCJ+yxe71Lyv3vlnhIbhJuLCiAyg4mQTNP454JzWw8
rUVx3z8CjHXcnXN4IcDPQQ980rYlW+Zcs9weR9ET/0YBuYXlkQdMti6FNlDQmVqrgJY+SLphRKjK
5tlpb3lUMjsdB+HhyqCR73bKwX4nGz8DJKEFTcLhkh6GinawmKumt5awzBbA/H6Hq1FHWSZ3AXn1
anc8/4vfnfKaPytgJ0POpvlsIKYrQnw7zjjwasC58SLAmZ4/KB5ZqzrEPgTT5My2kpNO0DMsCYJP
jz5hrN/G8O7yB4zJ+RfkEKcvvdzxWJDBZRqZMXj1IOgoLlIPzOY+Dmw19vmKkxyEmvIsT/cVo7vI
fkAssVjqUoVI9g7mnDofjgJ4awG3LJEtT+N6PUN33Yk3lwYavrZ9lD4cm/KLzu+v3pobFf9hOTOH
KN3trzoRAOiCGZMUOTAepd0ADJQj7D4tGjJZChtHYigTf7Pyn+GLVolJLEeI5hxI6l1RllcVXdu/
bBPjBlIrPutZ7Rawoo+oumXaYHMaALSgZyEz31xMHrBNCNZmmmNg8g+WxXaRikjeY4axk5V0cjGX
LLdd3YiJGoh3HfUyUzQkJY9+pxtu8uFspBEg49GvMMfkA/iF1voiJVydi27NaMRAqbXTl4HWbn5A
RVxliSw0EYm0SlIBtHg1UG//vJCYCWM+vG3Yq8YXq/htwfEIJRo22DJLE0fRJXkgHDWUOGfUM2vw
j575WTVOiUTRlF6+gpXymp3VJpU7DTqnVQRwcHm24U+Wt0E6a4QV+mY3gvGhQ0WnH7w2DPyVUPS+
KqvL9sX9R+crrrvS6jbqHV7qMVnsdLF/8EQbstPwwqrZ0QIzUOKeqspGPaH3orSwQz9+IoVjWpIr
Gb2p6IyXBdj62/AI7isHiVD3xZzcO7bprpJ1CcgcI7xhV6INbdCt8KJRH1mqVrZFuowkf0XWrtcs
rb0N9IrXJIS1fnTtiRGqE3Pdl+vr+29tx+VbbsvvJoFoq4uSMieL4Q+fSpYwNxDFEG2BAz9OHSgm
CY+QPQ4y3Xhh1Sv6x0l1tPg6K9NvIJj0PqSVAq93neyamstttVgDcR8z0E7z3M5xn57PNw2ns7gu
82UmhJZ3Sp/YFnIk2cioAWY8ebPvL+gaMCFFHOj0p6e8jex0zhosy9b/cbrFSkd3RrI3KzFXp2dk
P4VfuDH7r48/8jOrpWrfrL7vBlOLWl2Q9MRkF0qLAHuQP8kPvQhcKIX46sd6od4put4ncLLWoBVh
VdHaIHVptn02KfWDeQi7okHKH806bM3IxuIFcEW/+DBP667CLVfF0XDxjGN+fktGxCpk4RsXIXpW
sWoAp4N7/xwgIeG89TdiTRCmR3kWIgrIsLII0KKNB76cHGWJh6w8Eg9kSv9YiPVnnZBjBavhaEdx
kA1IrRL6+OQr+Ztc12ZXGg9ihDbZMMEUiQ9MnkBNcmXapI0i4lXK3ad7aNzGbfcaV7QDrKvVWDqF
axoJmRyoK9L32hsdDOhmvIMQVvSh5lOGgjZzdmAsygEuQPUaUQKynqaaoYipN4rlQY0aTyj4X8ch
fQe6aIB+G7h5ts2xUX0ZDcEzM2RRxokW3jtainsdCJJAolH9NDa678ZYDq7Hm11Sz1iUPB6mK7qJ
Q50WjSQUgLeyz51hyMGfd1pLo+B5n2hDllNAeXJkDTVh9ZBv14qMKhh6P8vPrzPvA9R0sugvkbl0
iSRxmGoH9uOgpWylcEZh/RUoe6t9eNqrJQZGqEnXcWZzUKrtvAcSh6sphLduPBZNe3LdwIiGLia/
bxrYx65i9E0ZslxMvDXReJFF9aCH8ZCYWZw6H49oBXP5wb74Kxfb97e4Y23HrIJnZdzhwqjHpFff
y6RqcibKoQif6Y5YVQ1u+4P+N/KXLuq5IDZMLJ4Kk/PoXzgAqnat2WqxdwduJoAXDoAxvd8jdI+l
pB5SOX4YSB7z3X9dUK/70jjIJ9yOieQrysdZHCLjRi8IkXyZxZeroFPZLowMG+tmh3WBXCX8UZdQ
+J+ouYRthtyfwjnZivov6JiZr00uECbVeTRllhsDs3tSUVI0Wpl++pU3fzuhh9f3PG21cBQaFK6k
j382/lkTADhML1tfAa1C6U7Q1ko+Nns/LF5yEfTowpxEYhakdevtcAa+OMXJlZj0C9HUAesuTluT
EelMIyPfgSVXsgTykU4JkY/GeoPW28zCLVn1xMh94Ye0VZ36Fg01jCZBlXnvb7l15NUHWn3cnTl5
4tcYiraBb0miGUguJpxnI7K+4haUa+BaZhYzTaSuYwAQ9qxwaI4vnsruumGIwtsmoOdlTeoq+MOW
imDV184Cz2Q4U34fctL/3E0lD99zR8+N+nd+vt6OQ9WYnyJA/UCsIb0dba+NOTF1iJH9vRD5epin
ExXrpj0wpqZaNOv8NUdaGTM/6WaS2Ewg2oyvMJDi9dwxqkMwuMTZP5aA5IIJYrwuQGltkeOs3jgx
X//gzZGXJSi9p0BR60ysgZhIdnWAvTaxGOAXfnEo2dtyjanMBOYTwBXARCQ1lj7c+UR6Td8JtFpn
PcgBg3WOAoN13iec0e7FqhHiD7wTYD8REgWwV2MB/CPAMmX7Yo0YaWK9WW2M+da+Oz5BjSyC31pc
1AVc6FkqWUZ047Ng5vvsaoyUHqaY+AQb3/U3RD3GvpNcKwUAjDQqiVxADZYAtTEaYIReq358ifS6
1urjT+DCkuKHlzTG9i1d8mWYVB0trwkt3vaIKTtIAQvG5aFzzl3LHyc7asGuh9Cf6AEndpojhqVd
zgTA7qjMItAFbhmyCGqPMSHtCzo8Y8Z3qn7MXKW8CM+0BwCRpg89oBqn/2o7JYn9Tw54mRkNAoAd
7KV8UR7IQf8ZcnXz7NEuKitDT7MlIurG6H8C2m3ySYnBy3xCiXkeus9KUbWGWAjG/w7OaQ5BTWbQ
gi4b+rpLCqCU1J6YCS541qQrZfFR2nfdbxfDdltZHa/83yZe0GqM8X8aBDaU+MzQufLCw6D8Msgv
m6CMr7QW+A2rUYQ0TzDGPHTUPvIqIU12h105NcP9sEvaJcbQZVwjKJ/H2yp77BEZmpJEv6Srkk2L
ws4rTYR3+e85XGnQ5fbqTtRtFUsG+I91MqVs7S4ED5Pb9SK9TRGHHYVlh9rSEVqIkGPBzlKNMFaS
IuR657vsK5KBbvLEQFQmNlP5hKm0OmuuOhRtvBz8jMOHR8QksHBK1SS4SvGxOzh/v65N0rzf+6g7
2XkkPiLfCmXyZWd5F7qOT7pNOEr7SRRTgZN6cjrK4DdaQ7Mcd5/EHD4wftDPHsxWOfd/aWDABoSD
A0nCRsldvU1g3v07b/kuTUw+eEEswwjpLSfnYnBHoEbpQxxxRW51bajxScvOzcKuLC4uQ6QnC7bW
TCT/jdpWG+aA6iiwIdFCm7ggIxjcFKOkaJQ/76LADn1m9+vxPzdU/U0NE6Ch1jTRNixyON5mKxO9
94HdkspE/2vDGnU0zuQ9KiV8JZ0vR+k9cCs3gFh4REmOjQmm1PwSR5dNUCPDY/Ws9aLIrlTucWnu
VSkGGnCXA+GLd5ybmTYN1F/veFk+9jzhe1pvWiztTuCKDrSSwl6snyYDUqejROjtqmTy8qMvrppn
Nfl+tHNszhnptRnuUHhpP/tFzaz+KmmlRDtKCmfGuF/7+FWEYPc1klQOdpU2cgkGcPajrsyeI2nh
v1DuJiCFYqsc9Vk0Mw4bAgkZcqb+A+2ut3GDe/kGn89j9HqV2RAKArSQcOG1td7EbuutM6g6CiFm
1r4EMONoAEtaO2MxjSUrvFzd0cPLwNo4LvUsUSbLDmptjy/uN3tfAoRJyiQ59UxRPLMPxNNeJoH+
k+fbBRLDHIizWI6rSdhD7bWy1KolpF/wqdIzwyX9kJOK+ad/pTMIxRNuRQiN71D7LvxMXyCJftAV
b8gM97C0BRR3T3LtlCpRZltJF7jRdP+XtROgNprY7pAH/9PCzj6GQNLc73uOz6bwvS1Sg7efntOP
WlaH/11Q33FtfF6Rm37LEy5TQNxjjSgyiaKF09kPWddJkx8uTQb+BneCFJnJ2yiVJDwdKVtmuB/d
u/Hu74QugpFtFbuXtVrLKme0L2eKA+G8kDyWwAe9PthubGdyuMAM7IxLL0PYHq/GjMB2i31CETJ2
GrOjA6iii3UTrrMBYq5P/3qzk5C0eEZYU5ZUBwoXNZQJdXZKU3BJhiEDfbFIqryU9TxApluQ+avi
ml4wD0wT5GezbTOxS5ZpDO0JcFpJ2ssK6mwENApJOWI49tC1h7HpIfYBC0n013wNHb7CpkzKBuBq
8PJU4ClA4+m3mf8L7t/hrq6ZPrS5R6vn9He2ltx1keiH5KYlYkJIKw9arE8iCNFC5wPIXwXfJr5F
r+7UmkJAVc3NbOw3Lg7RDVFavxMDOirm3a3PBQwQjKNcuxlnAD0dMjDlVhcV6krDZI7o5eiVzmzT
vJgw/nd3uxSIRr2WMjjs6snQL8C4ppdKDlKlWFoCCNBZ0F6CcfgRbdUBGqo3AaiFwyvhQKvU/ltV
5r500oQlNp5SRnDak1gUwar13K5Fa7TriEQ9VliP96UTh9JiVr5XBrorEF4pXlgt14v4JGq4o9g3
3sB34Ajt6NQ75ZmirElH2ZVUjhHiVkOv5B4vf0T8dXv3nANBgaJICEDchbVShsKmC5mYS21tUu76
59Ya8YSQp9ZBEnkgO1S1xVrRWC1MFQBvXWDo4bevclLw6mWJzlpH0+9c+9jC7Xu/fpJS1czHCoVb
mjZklq89ZGMJE5mMXvz7tLw7e0+lrW/xjmo+laBHpBmhwHmezHTg2lO0G61ZqQ9H/gtZ88PN9jiv
YZy5F56fG4hdkF+d98wp1b/4spXwB4r+P2bxKHsDG3ae5lN6KPGe43W4iV1j2d9JHEBzYOiE6I4V
lzh7CescKUxzmmfqEz/Kdd865j53QoMfQR9b0IKsUqA0z+8cdLZ+nEYcNUxyElGHzVDl2tbmJvUa
YGCYs4zzPkYpsEmUQqouLJKK23FPXzExzFFrkr4Km5LuKJA1zgVerzVsIFQnsfHIOzVS8k5uCHxk
MXqJQo6BVy6d5lkQQ62+8vpRoIeAcxFY5Hh1QYqGLqc/tgA9B7chqxov4z1i7Q4O9rKeZIivC35q
U0Qr5BMVAT7QuvaW9sR3rIVLFT0ry94aMspWry/pfSB10+kHTVPTYKTCznwL57QGvix+EBQEb5HH
gXiM0hATvoTWb8LkzH1p8ws4rnLgc7PA4pD2XQ5o2lzgPsTWkJfjB8FA6eGJVo0z+f1J76c0ZBk7
PK+LHv3Hbp+bx1l8el9tH/Re0RsKQ7QzsfiVCzg36179DB2e2pfnI3te/CuJFN8SUEbluFM0kinE
41CvtGhiq+x0fLdHdWI2mB50h+fDLYkgQVS2eXU/GoOY0V0af7E3bXbcqpUZwpEcJhVNu0r0JpC9
WIE8QMkI/jMkfU+C/5gloX/nlB5XrToxOdAxzPGMbIM4pS/frBYgza3cPMk2fPso5fLmoVC5dEnq
yZfs7unWOllI2IssyUr7qLNRU2XB9+l5BXVR6LIX6+ey2If6r3aa4ziKnqRO/NXuJgevVzC6Ol6P
XFxt6i5GNvXhbZ9E7cFLpmGQHD1iGZGvnimXkQ43l1SJQaK5xGx7goU62+xDLNcGf7KeyXOXH2KQ
ms8MY3g8dZvYfvNR5GZo4kf4Y5zJhSABrpjqtjEVZG2j6wDwxH8It5CYZf/oRKTcF+zhvW6undBQ
VWvjzgvBSMSwG5UHvY0ymSILGx9ToNfmaxpMzD4+rAbGIUNe/CdrkVqeqmb6aPuoxqRzjahGAl7+
W22sbvMpniBUO1dfrHmIJd4fVzCC6GTWVLDK/sFYLV7A1VvKxklhb3lznwc4Fk8Q8DXI4NP/H03t
UnB5D9CmWzZO+n8m4Oyq65/tI3ry6y1qdGmd8T9BAF7cE9GC1HyL+s70BJRPRB8NCUx/pxjSxe4d
NMd6D1D5tfyWHw0UAyFlIGw5FByj3ebplaVatfwHxxbjtaeW0lFZTzXP8I4yN70PjyHSThIBMMC8
4ECMxksOC51VxtL1Lh5MetP9pn1CHowLa/TmPTUJ/DqX4lJpoPYhDFaXRp5SdKKAuX465K1nhZqn
UDdnqgO899uvAmeTyKsqSl1NmRvmskZjFYrMyzmhdyzfGptGP9wiEscIV+TwVMjEzGYH4kPooz+q
VhbhKS7Q0YSPokdI5qvQm1hNloLmZQ15E2Xs8z/d3WxYLOTH1Jek/9Zvhc6d5n4v1JapVM4dHZ3k
YvNhA6JwsV9p0Ji6yP0gr5tNjIgOoDOfv2wM6J8kJ2SPqAXwjVQXfd3pOao0xs0oFjRWiGFNfYT9
9j6BTTktBEfGuONHi2aCHR9cSum3FU/XeA71GX7u9QVklVmb/8ziqgaZJn+2ShyqYZGPERchmIiv
dLtlv1S5fTVEZq3i5n23/E4FjSDJ2lO4LQTjeZZrV2iJDJ3/5u4xh74SyDAXJG5oaBFqT+4cPKxa
Q1OV+mDl9V8wx+hyoh2Ee9l0XNdVqJbjfM+K+WuLz8ABstqzRqLQ28OGyjC2AshTn3Y1IY+sVCs4
o4GdUDmxTU/i7w8y25K7SoD1Juk0nmJmGvDBgqOHJaUKy/X2nRgGBFoy9rQFLymXuIGZZlv2CNAF
Qp1CYpFn/XltGInxirAnbdAHIM03I31NbSb+j/UD14STpqgnKO5mcwc2dGZmRnfROsBh2y4g7Qxz
7yFtwIf5UcU+XX4gI4jkj8S9QLrD6a2TJi7A6M+WKAYd321C+a5M56PuH2Goh4iy5BaKygOVeP8z
kNw166rxA7B+SPPaF94lBCbbi7HGQPuCghFGp+JMQw+W5SYXhZXAFQ0aF6M64AGhm7yPQiD3hJg0
eNxWFxJnMtpWMGx0WHi6s+fWUEPSDdBchleuRQlPM3To4flyh9ugoVBibFxucusjyTxvsheLd/Io
d1VcxbmBwRiDweHw733xg9eGzZkYE/1VhPeQofJzNYtEhV88goraMiBoTRy6z/WjoUsTvKjL6EOP
ZKGgQrFN1XERc2TvGHkEL7P+ofbRxLfnPK6p2zj+6LNvXR7Dyh8FfMnXvlCDLUKVjjZTgnS72X43
52mWpSRFpjzhtWFEQ7Pp/4FJlkNrkH3cnPcSICkEMiZvHaftJHGcopw3sWsrCAB3/Q0VaNFnTavd
ujPRzlOGyODPcUB0hRSvFx+CbpAomHLEj3upa7e60AtyWL6Gv4LKlMfs3SyzbqswPZCjpOevM5lC
NB4pnqrbEaPcYpqmIYNVf6aEdhTt8MG7NKyh/LRdPnQ8bQEAaOjplcGDg1OD9wKISmJbBaGbP9xN
Zl+9BIFRARsELNDGotCfOjCHQ4qWYq95YPvcy539p7Bs97byGCCFwlOC9NPGsZKHD7Nnp6/BHvIO
58dFRgw1WYvrQCKTz4waLFOD1+DEedmQSVScHvn1BIN7U81G1AEF15FITDJegADKNF0wLYncUnJq
ackxjBxb2617hsj1EywB0Z0hdOdWVlWNUwppSXmObFFzIkexJgGIS7r4Px7VcaARNXBAPbI3MF+J
B2+FhvPLx3enqw086qrIBjYhfbsqqY63QfLASWNbrtz92PBYYyCoyDLQHpRTC/GzYnW9HwrpzOVX
GrvjJYAYs2S6bgZXTY1WeE04LgzCzPkApvPGl/jPfzXh5RRrL8mNaD/CaD6xIh+qBeGh9AWLrVqY
nAVc+R7yEAD0b6dPNKB69maxiR3mC/+0wTppYTZvTl8dXfqblVMmagf8sfcL0InVPdIPgBf3jqek
Ak6ZTFRh61IxAeXKCdTsxXs0WOEKlGy5ttwKLdXBj0bve8OtFXlyXI2X4DRGREH39BwFAzvbSDXk
A2yMUAKCwJJWTRSjy0YrjN019gOfE/gA/JE2DM8SoFTQva5nU9s+ReG/Q4n1/ynmDvV9hzp3j3hR
6sefyhiUijP6ITVfhg1NYLv8VwCTDCxw6tvaq5p2qAhEwG/96jlIRaWCRazwgbNZ5TpIVccu8m84
Dkm+0GsgsLq056rLzO50ZJobM6OXLo1n1UK7RDGYHTFKAJohmFx4PEE19/GH6XFo7x2yk6mv+O18
FfkMocuInzq+/y3MTiK1yl3+OSUQwqSGXyB53Kk42TNsoJOQHBq7gwxU1z6f8ZUTQwHWUh35wLEI
omDB8lVqaa62MwqkSp7UVTt5Iw0eG8y7Xy3oc/C4PNthmtQfudmMO3nX4vNJjPV/7Xij+AjHd+9p
IjJhCu4UQ0rBN+U8RVyBWWJv7L6wK5pTc5yaJyfWOJ6ZJs2xqHuBCQKsdTqdr4YzJ1dXwXs3siCW
eS4JE+4eGjxZUuOcroPwI//Sr71HmIJ4j4Lw5i+QB6WcAQ9lwcPIQWoJxNbWEzVI5G7eR1miURqr
QFLoHlN88kmWeF975c8EblyG8KuHiX2ZY9xvvtGOAiG3L8n+y2w2uvKJC/amtnT81Cxh4oLHTIkv
OmL6BG2KNW1WZn/subUr81+3Bglgvos2cSHXyTJPyQK9FkpOFHQPnPpbKhGbIHir9Ny7We1UV6CQ
rSD3WekMSumtEZV4YbAVlpdvj7ow2Vhg1bR2zlDxjqhwcn3h/tBa21d4pdftKD7mRQZ1xdqhgKbO
xEMU4nkxRtVKMSqWFRPN+QSzt/IozaUwF7BzxlYZMFXa8v2wtW2GgQuOIvQjYvtSONL5q2sMWA2H
cH7naCsQWeDNpC0pqrY/YsPTSV19S1Ap8AF0j1j47XjZ9JBiWfnxHtF0O7nKSRXiRFwLQtKnRJ+k
4HmHXmnpsKdQ7c1ntEM2QCyD86QOOrFSeUAc/qrtZCkCuhRz+MtmeGN/NB9bkJNCHyqpTikVro3W
c4shPabn8PRxXzN3AwCRodVXJr1XZgqyDVb3d0vTPMOmYwhd8enSMusR1fUdr6wpKwuKGQcRZkpz
hy8hr4W9DcDmDM8rwKe1TbII/m2WL5Z8dGvCuIe4PEqMDqZcFCDVwNeLj6zlG80YLllXek24V/5L
Z3k0eeTJ49Y+MUAYsrOghQMNOszgY74DW+KsrOjdAqt5nnSRJmDXeOL3WGutaQv62r6OTMqLN9xO
QwqSyZoykUKNvvP+jRjJ37wjxYbeiF3msZTNnkwGxFVogiTjAHXscWCA7Lb7FMRavOkU83Ul0Qb0
PZeAFe5H86OWOa2VoIOPjIVHehH84NQ8R+04zB121nLowDm70rMmSxUl1w0O8X9iwxnABwieS/4u
5JDw7nQU0z16cJD3PtB5kg+u6neIXlB01MumgdGIrBDf1zSIybR1isoT3jEMlIo+gTXrIWPWnoZb
d+quvlt1iDzANFS8UDNUJGjxxxPdjdgDnXjqmNokn9toidWeEu4WIQzENjQXPwNkddefvBAbGo+p
rxSGzzkD5sZ5d0XcFE1Q85hyXvDP3NGhL5ewy5I8jkdByfwIPIwHXZVE/vRGi436P4u3Doc8Z0T+
1hpkf8IKnFB56WBpWlko0dC4hGZzhBem34e6dyA7IgEyF0krpvcqWUlQP1DHdXCQ1Ljc3XY6ZmFi
t8cuSpCWlMTlYc9QYHtIpEHbKWORk3gKKXLJuvXqjlROW8ktyaP2m7lzkL1NiInfGrwc/KB3AwfL
aB8dKGh8tu+7hHyU9wiQqN85zGMPhqpQEa4hjILtz0A9cYM1ygrm2BVKSAwir9AHcfoolxLlH1p2
dDNHOxeEQfzAzyHxWe8TTJc9ff/vIVFhT2FBUHFMliUC7nzI3WKkZoEyE3kwW9N7lLPi0zWHV6WK
uNvo4ZVwRKEiIE/rMRNYe7u8GIhJ7V1Twjt29JlxbrcPYMio+FDD3XAnJx+Y5GVL5brSFMWgXDzy
k+xtq1uz2qFU/Y6PZVNIgqQzbRhk2Xcz+HlG6Qgo9fwC3jkYAAKjBD1vCw2wVJsRq/wxOi7iTiTi
pF/bktZoVVg6mveNUi2ulV7953nmsEOCbf5nRCFrqDq7oxiZ4BSWL3+BKU3ipgBG4wSVkhAUi7LK
b7vXAt8CEbrMFaRGhcelPKhS6cKz7GJE1noFnRFe/dCw2QHBYgjueh6BJ6cezQpMSL0fRrChLZC7
q0OC5CJeTfX6kBDmyKWZ2RTd+T3V0RvmNFcadkMO0DgtBS2mLBMEhHmf5ZECAbFxbe/2IMODBg7J
fW5ywuqLLWwoSuCzgm0P4YFh7ey7N/Wz9SrdxfrbOumqwtYFKmKAn+O9QtqGXcD/ZiCjhM+xRlpQ
POICar0PL3nuIciRHs91O/vKzrM20TOdOCJH4tPl27rKef8zgeceLCY1OI/irAXDGI58xbYbyrT8
GWnNm8ebno/TdZYEL9i2Z85Xrfj3hRCpotjtNz7UfXIyEd0gopxI8DaGoY5O5Np/3x9HPZCqw3TC
uQcu1FfQvNC5dGLifsMKfcui/IuHbz0oU6EqvmhHKeR7Szo9gzrtPihwiZlyptMLkNVhXJMpwLrP
/9afnrpFb5GeggwGKn2bDddZ16E4jSaMph1BkjCODpW0TyoKrgfoISLgYzvOxWhMuHEns6UQ4MJH
4idXEX5umsJMhAtLPEvSbRfzkVmvJGXfKtZluu5B7XvDfT/mAniRSqxWFEH32pph0/Y40+PbhPQJ
zwKji46lQ7w7jbbR83jA2v+/bE+FIKPXddyX0o06VK0SRrCWlzh46RRvpCIFb2U+ie3j0LiEpbez
WZr/WN6e3Wgv+L0tWaaqSKPFrRGGOtlOFvLJVa3ROAOObk0h0fwZL2AUOXRwnGf601NySi+tmbMM
9ML/vXBH8A5OxSMiuW85nyZv1V8fv1Kr6f4CqGNG8Hp8DkGqiOwmb88O9n2lxGlIJuL+hLQ0UpRK
CRISljnTZQX3ED7P+D1WToDUKTwZ882AHRSN2Y0faY3YOOwPZ9k3zKCZYS62i4oT96da9rCbd8nC
ccw6wYFlJH+wSNZb2S3stRgw2YucuFqwDL53eoN+fl42U4imibDUej0sN2o6uSl0wyCr38IkC1kK
XlEXvWx7TsLVbIeP9CSBVCeUZviKgr55A1ScBUG4K9DxYNW6yCp9NFxRYcRwuiwblxkznxaUxdKj
srQthI52Sl0NHAeJVtNtopj7Er4yGvvcRQxiYHajxMRuyjFZh/MVoMvdhb8RqNbA5Vk7kLxLORwz
109XZIxMbxwiT07vatSMevkD+OZ4qnIrZMCbjtUPjXbeKDxcdRLTdidxW4i75tfQBmNG/6mk46q8
JCblAYD6/rZSqx71tVE0SXJ5NmQ/HrOE+q/zRxRnBBiC3uD+Nu5R+MUSJc1214N/mjz36S0PQ9g/
eaEavwpvlE1cZSw5UX/BKhO2alB/cWXlUNezQNYf3uURwVwHEd+egbdUq//z5Lb/8HvfYdE64em3
Cl8vr1JE4FfrbmCn8O0YYoBRW9WEhQYxlrW+QFmbGjBTSd4Bx0E6dflL8EDq/tznwXj1lUCyELHz
UOW/Cb4wd02NU0vJxyF9anyLpPCQATRzZOyXF7CaozocWDtVQ+qQXtE+HYIu4MdLsP9AkTPT7BBE
VeIz/GOtGGr7EWnriqvjPel1ZljP/XXzaGz3SNWJ6z3ua659qtJHWmtoyOsSqRBjLM9DrmszPdSA
/kKOtPybhYV4KGIJ13GczwskS/1fa75YyVpOkWxZAJ8mMwbvpVc/gTsNADE11/nRJ6EhFXji9mgJ
urMJC/HbhFHMnGRH6qW5T8v0A3hcQMsJe3eTpm+g4+ByxoDHmeb8S6l4isA65ir/XqjmkuTy3ksB
s5DbvW6mDksBLO0wggagwz0PfHaRW7Kh7+/R2vbb7IgL8g0C++le9wSp1KzlMphQa4trzd8bZdJ2
7eI+Yts+rcQyg9KaULz0p9DUzGzAGfiMbaW8lQt+KKNAtkDdsIZVcPiUsTmZLNppp+Gvb7noLuS3
UcaTfKzUzv7yyAf4UHsB8s4/9PCZBYhp8+SXokT/TGR/d9GPiox+aTp6o5//+6IBuCnc6r6hdiCj
jXnsPVZrAkjN7AHFRX+cWs7H0nf7L2giaCnOdkvGixylJkTmur1Ok6WKtUs/o971UHTPft9auopf
djU2K9cdqjqZ0rnijABId+QXmwwafmaInU3x0b3gt7xBVpqugE2XrkHOLsNWjok7+jiRPANcswoo
TdqsUZwvssKNHhL/f2r2bYpFxPX6mvNeM1UJvfk1jSqdiuANNOBzBa4f5mw7epzwe//xThSUcPGx
ZXoEQIL2V1w0NEHSqbcV4g1clvGyvST0dg6HtvfzAErbEM5R0Il+EFOyCJGsb3LtXXS6MusbjhWX
KWxwVVJuZor4YSZFibtb4lOLE6wcNFPWz3WotXOFiWuNHB4FXcKUccD0kmzby7G4Lw5pvlUERqZF
4SAl7FbOlw98+wxe3Y2CRZhxDH3cQ41yjOYI6rFYrH0sMKitEquJW5PHfZxHa2IXE9e0+3yro+gs
JOMewJJ43XRWV2SDsQU8OW/Te1rh8vzRvjxvrQnlHciQeCZAU8JXa0LGG6GVvzpeYYQui3b7KAgI
ds8iY78QB3mCwPawtG1j1tSzA3IBKYiLSSR93AWsNNiQprGZBw0z1md2hkMLhwtgMo7R8hQxYcEp
LKKEMmK3o808PjCVI3jM6M+j0wCINRYUnMgc9ogxqcUkpokC10x9EGPjXSryPwWdoGUvupKP+p19
uEcmckRJSynHKvPyUmdxxQ1OG40lv5xJUc9OC8n+HQbDw8OHmWduz22pEKXsLHBgKC9BJkP9T9R1
qLp4csLJ0XlTm5QAoDF88IWjdDcJ/vLW0bpIRyUwT3n2QoSahhagsdbBziZZ9Q1l8xg7Vo/cNuNv
kd+lT4h/2An4yojqwPEV0R52aJ5ToTEbydfO09nnKXf4dbpP66SJEcNNb3y4Jm+u4HRVLc36CLLi
ExMnfAJwzf8jUQcTjtx0nPVwuFEibUnVK1ygWA7ZnZgTQl8iAydnTnQUH5epXSX12uV9wLB/slyE
NB0Xtvnb8SvmTuJ0P30XkxNC/GnmzE/C/n30Q9N9CjmDBQZ6yZvSNYxKLNh87FoCMD/3hRxhQQDz
zMQMIJWr7DM70msCVIYkOG60EJ7gj0SKvKFepbhZ6HnNbVcaEId8cmkcuXpFiP+DGpymg3u817Jv
og6OPeTc16QM2D2gYYHA59Xskkkbs1EPS9xkV4x0NzreJBF4/A0VpMg8Ni6z2TzaGcIk2a6Sk9sE
KVC6Bs8Ffg06Pl/fQw6wf8PqQt00fNFxArKPHovE8QAfcsCmsXwJv9lDMeOiaXoBoYOhgx5BlIIV
AKcxNglIBmCIGbWV9mEChUIk89BCS4/rr/pumbLNKVtTM2lGIBQaaPYkUf0TDuyFQdUt6owSUikR
uHbk2ExI1qcUZ+og3Uek/5pZ9CUqNz2UeBVpSzaQyTLIjxFSaMsWNs72yZODCCcFWMLtrIxvbowc
IWIU5r2Ohs+cpDsi9pZLjqUZihcbd/kMrEZZN006q1AhGdgcYFvxqJha8jdiJ6hlbv0PY8xbuw03
tKzbHW5mTWddNs1TGLs0nQsTuMFVOyQwWfl1HUTM2w/rXiflrQ8zCdpvR2/2r6PcBtSsirni6if+
9K0b6zzFQY5xAsx6Jf//TfV+eYsvDe1P0YNIjbeIxhGzZud1EdY70CkuVv8mhp4beMwm8dl5D/Wu
1+OakMV5zUj5nJyFs8rzQ0cCp0vroX99Tnjkkk60WZiRXfYl4ro+yJkPWqmbt3AXhRHRBw+YQZVD
qiz2QW2FezL8anM9D+I9CRC0CHT6Mp5tVeJn6TWsgVszkiSekFRleTVAvEGERggwSBDqH408rbx9
sbvEfP0UJIU1TT7/0yB14nVsXdnWHjZU+I4SUsJvAP4TGmb3KlfDqTwd5wRFLHI1dD2JG2A0TUC/
q4uJiVr4cSV+igyyz9iJnMc5P35JJeeky3PSIn3vEWVtsjKvNmk8UZIdF/fCcQAxhuw32SkPFQwy
J1cxfu/klPX9pxdjNwuLdMpH7XG+Zy+47ncBTGNiH72xgl3HXzdKqg22Cr+StRp4YX2KsoIru598
C+2Hum1mWwGxFMJh6TWDvROBK/CJwjsB1T46utBVmMbNeZUzQtE02cjnO5zUUEoZEPa7KhJPUb6K
9ouH+FOC4SBApOdVRT4xfnCySBajCo/BkzqGP4B9Gl5jEn5QSJ6HzJnDWR7Iz+y1hhts8Z1OEKTq
Du3GBaPRWch8iMdmrwUVcCnPe93vrUBDb/S5e9v4reWMoTXLqqG1ifoDmsqdNiBiaVzn4cpVLZPv
4hF4ZO7YBLmgx9FdLpQUQenyNp1Mhnp8EQspXxLVwdXkBBBgjzw7J1uLJcAW7THXC4+mWzRUgs4l
dq2uGxtRDRBA11PoJniLiCqmw2OKLXDYTSGu3X2AzxdoQZJ80luYeGUQS/XKtEG8J36ftV5kv1tw
quLJiNuYlNB02rMWeTY36Sn3rqsG7tFbIdWB4W0cBWAAEBToSzYq0lx57m8GsXYRF2PfpT6vBfoY
KV1HQNcycPyfx1xWXe56U+Eg9OmzySGWEo4f8buSEdoTqo5pQVEg47EeVlwdm2LG/iEghwohOfTy
LOMQ/lxhwuba+oephm55QNq6drhkhdlFrnBsnrD6xuP+lOwzTUKhorArLeZDgUl02JEKjCO+6rQz
QiLnFx1CHSH+/mXQEw8588ua87ygH0PH8r+EpBkHUiWOd1Az2e2gzcg9JlHCJmwydgz3fH2CfX47
J9JlXQU/DHJL1u0s6VsIxIzC5jpdIZLrVzXFbeQkKxM8sgXaGm6x9dAwnHU9hBr4AdQffvnuCCKS
kDKsiqJK6Z8lufIuu8BIzeNkTs/hLGy0K8phiC8X/FQuq4xgDh7n4Ak84xGzyduuSShAk2Jqq/Gd
KSFefHenJ+pwRnRbzDGoE/z+d2DqOsEdUPvpgq3KPGl4KBZWYl93onT0jEDM5ni0lGTcKEIPTRJj
MyUcE/YTUjOevkFrdCp/5SctHQpeh47m7oiba26vtP3cvp8SXJKtFixbmI3FUvqvXxIZGWIsbZIq
JU8CEImVoit2CLX7DQ8rhZSy8Zn3f9yTklrRnAv80gTOCI7FEcB8OM7pltZ6gw+9/gDVv65pSukQ
R1v3romo41V1RujMWvENhu0Urj+ZfdmFqcAJAV7tfQhXVEAdUdR0fzKTEfcT10iXMt/7QTV7MUek
xOXUFH8k9ykrmEQ4nk1deTVg02kLguNfLZT/Jer6ey9eWOpQYvpeVWS4iEBjkSovtta4LZZyhGgG
yptdpPZqqOiIIUIzYEYu6xBPqVN2NxVxoYnZHVmV4dD7N6+e58LNv8im4k0WFn9VHyMli1mqsiib
T0UPUNTqyds3KVIX7JV2YGmJG/Ecc/TlTKnoZRZSiHsogRoLQVgjXfyGZ2EflcetKdhkv/4n912l
8mWHO8YmAHRsvvdS+fWsonnGOdi0yLU5FRr3lIWAdE+3IP5NdKHgXpZYr8Y+1mFeV6qyDy/lOrYH
UiHsxMsn0GcR9VigoDKXU8WQKYyK8fadazt/nIehTkeF28US0iskBKDqn4j09lJWcvNC8UY4Dxqs
knaichhI/b8QvJ3Kx2/LITy4nwQt9ZjweGiAglP3eb5dXKcAofSch+4uA9uUBAQQVXcbHzUtsmyL
Y58yiFBbNHAAR2tCbTJ8628JVAd4dcasQuNVW1ggrYfHRdX5UwD579EWW4oBQmVwBtskBlgx4/8J
z6zT35zxUZ6SiYlNDY0xdcsZDLm0vYB7MZFFg9H2qBrI01noGf8DsyecqFNVcoD1MR66pnr8gdfe
RSam/1K7o2LsXxTJ120jL5CMZxXjWVFPaBi+r+eDLlZzqQfBUvG906JEOlDqWQYOFOZO7KVTjc1X
jEEtIMd0jXKaZAp+lUMn9KGR18Fd3HhfIgcHT4t+HQQ4XSxj3JX8jb6fuG7uegnfSszYrASD2o41
LhQfAzyWf2xEt4Uyrc1SXF7XibKMCdcQn1f0xRsy5iIvnnsNOuObvouJFvppbEfIzxMbEO6Jr1zw
L8o2QgvYXhho+IpnGxpYI3r4vzj8XCC0P38b/PZQ+bY6VLi8DFWRSkWfL2KZ/CntTcaS1VazATf3
R6cSB7mpXgRCzTRriNSP/lUAFgxYuFHHQGNwOQu7Kw1Jq/+kCEIHs4KetOXBbgXJI6xJVQAgc/FO
nKSbTkWiv2v6tFEIdwbQARJI2RH60TV9gexP/KNLeycadjmB2BzwMPoBsnNRdmYvV7OICdQ9bD9K
oQZnvdvXquUZBh9R8aoTSubSglbULRsV/DV8M3klk+WP3xqjKBsJBQvFlapmkvLSbGaDlr4RoqZm
ogefrgq1fgVeuCTzjD02kOTQjDWq2SXjRVuY5ESzPPDbNi6nbM9XW1Mj9Sa8dp8bxJ0zDp9lV9Mb
II6TOyJeNoII+aBaAkqvtlpwgUr7hBJ8ujsiVKpAM2Jn+xFGCntPXsP65ubF46LuWl2xd1RdBLku
xzvkKDIzVFwXkoMXNtZ7NC3nmPxKAafYZFZTCxHKVQGshUwrJExgAXMrEKynhG96etFbkWQi1Fua
RSvigXzfoc/KXnxrMnzC1vObUL3c8K1zTQZ2tUA2OdSeS2C2YzSn97ojHQUq4s5tw6qGyQwyedRX
w4udZJKOpCnGByWbjZuI1oe4CV0dwt2paN3BJVS1EsI9ncwiG8w0f+6Tvx2o20dYfbd/74YkAzpO
+reIsrqMmxIoTo79so61qICTtysZkPdnyJR7oeFJuD+LgopZ7qQeVdR4x4jmO45rsF1GuERqAY4S
C3Tw130SwTt15Dfnt3/kOvVO0MoXLKIinPu8B7W0AuRoLAipf2j8AK0FwG7WKauRh91n9s66QEvl
DlkseEVugsmza48kX5NfgGZ6frZtqVTjSL/yPzg055p1ZqTxkw74sTJjAN+3+piRgZi3r5HYac1Z
Bg1//xGnlBSrDe3Qd/r7KoC3nM4DOEALsa5O54CUdfKgIfA1/6yCEeTi0Vv3lPsWh6PpF5JVZjWv
Sds/zLymbW4LWXg7BRH6/p4XJLTpqq49V2nExYh35TtXWlKGifwcP+d/VP8qMerc7ZERIjhHUNC1
scA2iwYHDg2Y4hnPeUtg9S8EVXYGyUAZu0PdAipyDXLu8QV3KFzUruhXtdbr/g9XtZcfAq46epSN
P/4OTT3jQfhdTgwGiyzUUJKS4LXbexEqsUVb3lXzeJ+sje27AJd5yTNUCmdxOLaZ2LJaC22uMN0j
ZxnY6aBo02BjKDZ158bg9Ns3qGhZkepJOzD9sTMMPbXdZc6TIbydsYUZDaVr+GGNjq5jDXXATLYy
h+b37vFwplf3rz/Sv+RB9iH62F9BFoZWVP9CEMqeFR0xaG9ffRlwMOIUCaXAMe6bI+TZiCR9gabQ
4nuj8xJ3n+4PnH7R92pR92EA1xI2yOFiownerkoe6OjsjNNOte0+dbda05x9Z+/u0xV240GvYYLz
bvT9HJzOgeH8tPsdEqn9todUrmpPFjzmELtbwxIZXCcDfLScahqZxBHS9VnyNkldJpvBLB/yYlPX
rHOlL79EIrREeRNZsWmUs6Lqf6L0LzLr+MIeUAkp56x0PxzqPuanZ5IjnKDfbtgTHP/xKe85M+RR
FZnedCvnOWrFZHBQ9HKc/WLfJNJV+L1SR94xaOK7Hbgl8eWmPh8i0Y08N4cdFDQot8sd1ihyuuoZ
1n/7tTFKW0anpZrIvoMjHgOp3Ut2Jr98p24XWsN6S+EXaEvyntr5Em9QGtPBk27uKnf3l2HoWW7U
Lj5cGpik84Hz+7L926FcB5l7IkOqhmqWyglQkjoh6FtBKcsCpjG25cD79mpaJUB5/gHeDGAvZd32
7RdbDTzZDEixs1g+AFsMAriX23PDtAGMEs/PW30dvpHiOTVmHnhpL9gE6BPV2EuSZtL822WDITdp
PWPPTrnFrn7Z7gXafJUzuiBxgWTCDqQr1zzKaFIV3j8GohuBQEszuMVjMDD86jSGWoud1c1lrucE
hwHLyTKJM0Z0uGbAjM0/Jo1dcuVRmDn29eS/dXINsaZhKGlT2Thbb9zkkqD7E6ufkx1pESEaOT8I
JDmXqIOVh6KvkT0kaeAMJW7sq1gGOpwcUZWC41+wxlYA/f4JIWXVlncDC24AM6H+yDCsNM21LWnN
BssnG6EjwpEz1ZwbtoD162aqZ7CqaJZSu1ZFMbGAS/NTd63TH5IJHV+h+PAKa95V9CRJUngP44dA
kFoaLUSX9ooHRo6BvD2axRaWhcYUlZCju9lKHPPDzyKoJI81pagShupOh+wpGcWFrxLnkhVYav4s
s6FmeJ3G/5vQp/x+kbRxmmCGiU9C5PyDI/M38K779Hj8s6MSgbNLqZ0TpEvGsBLCn/QaB+XftIvj
eygIr/nsPzca2VTryqKJ6SQUIy9MesI+XNsaEjRFFBeuGhAnWrminv61KibpKNpVryijj09WYISA
zhv2+R9UUKxL4A22Yx6ugxr4nKbKopT5dgv93R3qkmiG/QKTbtthc7iLXY84e/zIqnMTlTibWBaH
H08dVUH9Zr9NoYRQt8Nha0P6NWuWHKkjbXN4WC6sry8DVp9CxKMSUWpWnIo9gLgmxGNX0oEM0o8t
WLk+bAFDMoT+S0nXkYyEohLo0XR39VOIiX8o0Xdn8Jd5Zn26F4khzQjrzp4JBu7iFuytLBNeT61i
EzszaAY+RXquHlJ7cTRD4gbxfT9PSfSuQmw7hzhVlipz+9RMgmdfwbE+xJpEXaGgWFIojKe/wcC9
uPVNHw0+WWtXFiLd5tTve3ZEst0mrl3RItUVcAF0VSw/rxTlLszb5GKM+3QIs6Tth8jGcjjpoAM3
nDSdFQheJTzHJEdNhUcle5EPyJTm4knoI07v6PBUTtxXrn8z6AE0Dwr7hiD9N+MeAw+yo0C/TXzO
M08hUjbDg26VBLhZjkYPx8+5ZkephBK7yJIhP6NDtAz4numTfyL7xLqBSzpzpPtdVlASfu3w7EC+
HmFLjjlIwpos16R0QYJWobWyczc8n4XcENmIPxLZG1rPUymtJl4fENQcpRrzr6gsJeFBCshJt1DW
J2ix9tTQTJ3D2nYUNu+TONOj1lE0md9XO8Fx/X1469LygcgH/FcJ3RfAZ/2ElmjCZaEPtPK8GG8C
VGUPzxy/lMiZuMK5w2uvb4YNkurkAPmbhKYrInIk/d2bTlqz7j3cumhGs9nrx1z2eX9VA8r1VAfK
x/CzSsTc7REABhWDyvHtI+G09ArqTZVEZu9pNGBUaiyGfSaHG0EQKYU2UFOMswTThe6Q4g5nlz6J
bxa5OfJR4ENsX0FD+1lncbdOIbDvXB83N9mJTj+M3iCB6r6cb0PkvYRQxVbnp4baPSp+2ZvG7N4g
64xgjcuUaEahjVPF1fGzif/tJ2OtPuDiyAkVurYRxixP8ROGX+4Scq3mb3xBZXHPWfQgAihvJ3JQ
q8oU3Ro2GyRali9d3jEXa0Vk+seUdGr2FbssXZ1Luk24qTAJrNyOAAzhcuVO9ZgB9iuvHJCIf6oK
HYLuDGf8QvuHU99aKzc6tWt56N6fCrinQDycVS2ZLK0kXmxrUQqNyXB2bBNVGwLb9tZo/ySHdAZ0
H91QMABN4fwOk6WEbZq8c9xnoHbMbqMFmdcm0nb/1ShYSqMYLKBrGS74xy8omXk3xA4P5Q/KNN4g
A6Q4PU6Az4+tAjI8JoVT0bXUP5t0VL0+0kcBe4fUfeXknKlR6PE9n4OTubox9mlV08S8h/IgZxk+
kGFiZYqF5FzOme4vjjmEVa2WBAbEUPAqFeXPd5pGNmSEHp3aT8R1qKyP6Diq30ggLwxtQ6WPj2zq
kJY3aM1hVQ29VrXLdWYGg21L9lmCiqlrs+ISjuSUs6eS0stMbRQg+CYz8SVojWubp5APMsiITUxr
m2QMEvIlHQ/ZqEV5TBf6PrkjyBoJwSPaYdnZLbEk3XFVge7Dyv5yloSS97920dyhcH6HGu0Fb1aC
I7N/MPDN0CxJVgk4nKpus1FWOQ75arQ0b/4Wu6sKrGf4pjLx+CE6gzw4yMahw9HGJfAiFfK6JIth
/XmERPw8ya7gogjsFE9aDtmi4uuNGsswwgHVCRObwcEcAk6u0MdXcgkFx3YXbPvRkR6yKgmUnABD
94b7RY9h6/tqTNq1aKRJsnj590LVKVZslWd0EfMC/kZf0aUwbT1vxVKt9HVudfRlQUNATtvILlKh
Mdlzf/Cc6mLmDie1+XVZJ73g1SiumbponHsD1wt+0iqC7B59Jkd46wcaPS0bjqg0GwnGm3AFb2Ou
MuYvjp4LV3ShPc0eW9DBZXdCMMrUFHhAnALZo0voBqNPRgDr/p5Kj8VrYFQ7F6FFBZRKyInIA81P
aFG6JZW9AMKojoflt4XKHuErfRE9aonJhUlI8VjZ/8OB0Q6IVEKjUw25O5ZI6xkC67zDfE6Mt7+R
dXN6oAWuVugTtCceYNEjMokLO9V5VpIPKHeVNlnMxM34CY3WhG8/8my1U8WHgq3OeovUb6xRWpJ1
WiJcGg3ecOQNF5FfZT7Mi4DhCFBsPyXSifZ3c1+q7XsJ95VqQNUGbEhSANCTiq6Cab0b19Hz/Koz
zesPcRZ2Xf9dj7HBI71wvLX5mn+tXI3JJjC6DiJ8cWhgasYrQ3CIJhUj3+E/zmcANJvifcYE3FyZ
/MApmDfF3r7bddjMmAGzpu2862MnxhDz6gfu+EdbMLq2j4wWEQNb4gI2jPBBQoY9mR6vEuXEWV1T
yCXi7fE7tqm+fG/GVfayzSbJEv0fAlyStOVQ2wpyhps/1pZADW3pCIURDnfWV4RVmoxbz+jytNMa
qk5zLEFh03bS9tWsIpQzl8hFaK27eSV7xMfVLb7/VzscyTFACRj9CbB5Sto9m6/RQHAYA128msEE
x0TNupCFehro99CTNnq4dbl04nFqJs97I7HK37eJljsiX9cDEJxY+eapEJfgdf3NvrR6F7MnD5KP
h4dXigd4/MLhutM9kroprPxKLLf+ofHnqg1/Q0IJOnzMkIhANEssBBIFryRVtPrqJdI2EIxm/Ru1
ZU8oNue2xJt1MjrCzykZGcEolC4j6UoWBvGe0Q3FKru5Rc5dvRy6Q5A4OhswmsxdWx94ptKBVf6I
ELXAvnSY1ep+HiaJDzGmEmbSyZof9EEnMN7t7OVHWvGUFtb/aWSJSbQY2reVc4WKhQUJNal93+hm
3tw21Q+UQdfLR6BQmliui7CH5dkp1gqQeVW5adp1Yz33gs0UfzKPZIyhWPRGugQ4tvdLsaxSIVg7
mqg5yQ301NI1sToBDoi/MDa6r4Ay8MPv8JDhuIavjZqI9JOYhKdfb1w8OB8tO5vu6qEzRcVYAn4o
6rOyi3V6nKUaXON+auSyvmdDq4NKM97WH/7i72/VUAxLVG2+NOhPdi908llqPkRiKNVssk5xPUTe
gkGyCD9IIqeIf5o+gv5QHNm1LUdUli93y75TWS+/B49Ns5xi0owujbs960OVT6EiBkdcTrF8jTWC
JwD9s7tozo8L0jw98L45kAeJGbsCWrTl5HtLMy4nuiIX4GMfETl9Rg7QeHFucsbvYKgHkekZTS+L
Hzoz8gEKHSDSxdaicQ89kWkotTqlV6RjX/muIQL7b3tuPG1RqmDnpIelvfqQ1nsIci74qsF7xU6f
EwXIGmFi1++/JumsYlEDDvNAiPRZoCLd7TXlQNGuhcF4TSFMcm1Hpcs83undSGzUqGKEJb7fDQUn
ZBi1iYx8o35mXlC5z/UeMBfQJABBm8cVx75ucabgqMJdfL4o29/a/dH8I1qILxiqE/6tq2UK5RJi
bgV3mWJAPspb6NNL5uF/pl4WuQ53n3wAwTkZ2UVRhcO5mljFCzXdyZx/4sEPVYLcaLGK2/MLMktN
/9NsE8dd6WW3tkwpYsL3ijiU1/x6p3Hx7n80F9FoIrbSPoa4WxBbCjXHM44zEOe2KdMHnRHGOy4+
W5JebSKcAcjA2msl/FKTSwN88okmyqQRkfsDj7HFhy8Htg7D86P+TJztH6iw1XSq1upebLZkS3ra
95V0mbl9/fukTaV+E5/FeH0aJC5U4sGCAJOQ0aXhQ5jQ+EUl57RAebuQVCVCDbGORy1DTjgpe7Lj
pk7eSrHjqc5efRC1gzOnMyhqYQSWPTm1ujD+/pzuC4+jR8wV1uj5Y0k/b2CNd8Sm9VJ9OqUwMyY9
zTapecKzY4D2pZP/f+MrafbzHf/nlajcOonHVwRi0bf+L47Sp9Oy/2sW/4IBhX04t0741eM9J8rG
FvyybHiyEJ7lJV8hy9zewvRWUmFFsNvZ5jvo1Nj14UrDFvZS2jAhohA7uHUN/Aol62JlXtHbUeRJ
2jJWUfa7JZUnTYCsTQtpvN+ypJxXXI680sflPp2a9VP2r4Ra64KhTeGfhknAJNyZnsKPW4K18uoL
iODwem2jzRNGlo/V44uw7veDAgcRQw2nl5EGrb0CvJdhtLM+JZNOub37iU7MgCHUBKUHVB3URQOJ
Ku3hNlwgnHc1vfdV9MLzbpEIZfD8IVRPvZdS9Hh+SrYSGtYHNw8xir7a5NqyXxP0Zt75k7PR4mK/
Ol5IfjJm1BOdBxl6ZUgniAF7i1DadQBGrMLCBSuqk3ePVpWqweFt07kVPkykWcMbWBGcTlP6R6VS
VMBRUAUfpK5umfSzm82sJb3H7dhl8VtE0/NuU6pQgElcG2BkQS0vMObByY1fLbf2p0f6+1t48bcF
o+81DC7iKnu0V/h6Z4yUlUIN9yYfAiTbqRQoGthC6GEDpPOnRGkwh8fUiwZKl6rz4AUUrRM4Ff+3
BA8iqk9ZWQUrX3wshZhMeYXjTrQMuQuwAie6v5Y4NOJ2ZHFP0Iv85KCe5RJiY/PjUGHieumXcuEZ
/OAEuol0NBvxSILV4iSX5DOzc4Kc2yPsXrZty10KI8zxnSGzLFkk/Lt47/A9n56unGG0srKlFEWf
K2tYTw3R5nLG0VoFJDsvN2kGSGPyCpz3U32/yORvWJ6SUilyXo/NOCa/55OseFh7YQGmnY3cVuBH
UkhF6Kf0BVv8ha3L/pOTx07eJGCMCnCxHTt8d6AKlROABzpcNDjng+lJTaNrnmJWrAP6syF8/acN
g5UKIXAp9uKRn32YVPYnQrUwwUDH3VFad1BD+XSPKM2fpfUuLLvIy2HcE/rz/tWCuc+ntb5zRvRu
EQLethQTRr4RHHmWJu87nwGJkIMYWz1evCqiQlYzDusFKhSciq/vQgvWiOnZ0EtVgo9uSeptScoG
0NNFR8nfTEJoWg4FapuGoDerTce8CxcHAlJ2fG0tMhVKRtpvg4Vs7wTTro+gBD8zLE3orWOTWiQW
sXCFKlFXWaUEtaeH5szmg8DC2ebFQWEKSTcjYZL2bna1dR6vua+DYFUfmglnXKof418/n3w2+ObI
8sWPViWYv0THDne/wFVnkdLQ8mnNcbaVGXR7lLHFL5Sdt1LJ49vYpEL826rD1ZC7cYwCcXDhKkB1
GpxAQgL6C/UYM2T04MwaFSohSfzXt3l+liLrw5JdALPk8S8eVUXXrl6NZ5qZ+6QkA1NMQ2OFHXNW
E/hYBxRtGuQ1zZUwnlc0TTcaT0eYWf+k4tAZq7vuigAfC+ce/mQNnYpO9OsoBiupsTD22wV3Ii51
BswGOfhctSaOi++JzVDQsJA/yY+6peGyqHghk25C/k5XFFwLEMWoqPZRWktBTzJ8+YtMoidEKku4
g7aEA9hVMHF4sf/lQ/nMvFoRGucnXJt7ZBRunUaPeAEJeE6o9e8TdYjGzp2NCk3x5WnwwB+g6T6J
YumgNlYDCL2cfJkDUaUbRX79832guhFCszSssd3geUcyuO8YkAPwr2BdLA+uU/tIytN6cVvoNv/s
Y5v5zKdpKz6riQY7kwoCuvMyCI8l7dK7Eln9nmBotgHotTIfVVM0c4ZIzep3r2ojS3FDn5IrN/d8
4PHDMxrrr9hU7IT/mr7oocZRRA0cv82KsMEvBkA0BD/4orBLTB1xnHlu+S7F9cLbx1oSTNeOFcpz
9Cg1tcF3VKFSRFAUmBf5qlLCbxDMyj7gatPMWvoqiOK9t/Q0Q5CodkASLqzdJDMfX6tTa4loN0SS
59FCzDiLhON3cSIuf/w6f07aRysYEOlEeL0ir8xMRfTNxG4csL7QrOsEVlrnT/7e8YvSyVKsxaFs
lE017BTA3/oMDYsL2TgtFsSWp6cJ7MVBg9js8ZWG15FhJek5yzKAKqRHaYxXpmzUmMuX7yVcAbcH
/79fP2R74HY4oha45bhBGelLLJX308LU/AQEyjafFwz4g65q4rNgR+kaYvHdXRUzNs+3lGiVU16B
t5a3hPQI/gELrMFccj6mTLMDkLMVOaQ0yBIBrIc4ww0TnOB98FiI5YvniLNdvCc1hDXzo7SuFHjD
9IbfFGrq/FLmCXhuv+gBCBqGcz0vOlz12kp+Y+U1l5TmzIHt8msw3KNS+EC1fRDIc0g3tjH7lvrC
NqLu0MUV/GW/oEJFBPhCGJSquYT+gIlvQqbIScRlGZZFOd4Evsh+MzvZc1aOPdIujc5vx4CrKf7d
SXxS9jbqjocAY6sOSRVz4Je0R5RqKaBoJMihAQtZ2RJO8Fx0bGvKeGR6L8yWgWKlL52YezBHi1ri
11E/nuPXmFcUYNSlwyVRRHLrEbV1+CTT2blik3oTv7qshFi2RzxzAwW6P07Zy2OpdpedHdOnCe1P
2Gtl362J96GUAAHHv5xxFnexLzaP7KoOC+Z/EuFm38NXQ1E6qR9fNTA0I0b0+XYvGYKH/quzAY/u
jCEorPiGNKWOc2A5dSO5qFCXRBBJm7cbVQYfefuhooN+cYvXZT90VMVOgUnBbPjswePWPdPLYjkn
0ZLE10hhXKlLQ449SMl0m1kXtp9nIOcn9UDQ1yFIAfsZmbpymNsOme+IV4qkc3gxNrht32K1PQZM
Gez1pHP+g/oYmB3qM5gO4gMapFWbEPtdl6zqfXYB4fRQrI39xfM3M3QzXSGFOCiLfdlXYsvrCRW6
Y/QglW8uM/y994LN1SlK0XFj1sDO0X1vxsQH+7s8qCuo6FChETnWd4LdkGQGMCbcnbwqwkPVzX+Y
UgeJQjdsYkf2Haaz2LqK2e3pzPctYfZ04l3Kr3xyyOg0nbt1IhSPN+fKRF29PatF12hNT8Y7u4ia
gtYfhWECkyuY7dPcxAwHzOGpE70x7/LqUGvy7Ky+iTXds/kRYpdEWKGMxb0eTHgAz6+YN5QtK9oW
5yAFT6gZGR5eKsHXTIYDTUdCI1/SHnCS53H3g3+cBIVMPiqW6HPCLxVsT/UbJOCpUoSjBngbpdhx
OcURVRpl5Lv63DM8oY2u4NU0Qh9T6ExnGCz8dBNXxqURaF2oZJJhOK/0MOzoZ2MefXweoLV3RW/i
ZnzBAKM3ZCdV5i2Mif8sFWLOec8TfAaNdfcW5ab05KzDAU642ZozYPmf0Pt8VlVqPztPKgMTT2Dj
9RyOSdXxzcHd28RQqsWtJFmYJXFQWSwSxuy673CiP7/GOP5zgBMWtLCu8gaxLZFhYRbPQ7QSlsE7
KWXLQTvYVDF2TK5DTLJ+R081jy4pu+8ecoDL6i6IJHPGJzb5GAwRxrdTZLjUHNSeYXp1kI7YUjgN
rEgatGVbKl5wEgZkZfanwZNkoPDb2JB9ZWrGeVIFUBpt8ipdf8c/bPHGgT1YIdziftQHaNZ974pk
ZQnr9r8ug3eY0IsLoxqM+JNUJedR/lYJv+h4AEhQWiGKlY1fSdpk8TtYcYuRCh35EwW10ZREBvue
U0G2zM4T3YeIR4iUeAmaxfnQLoBqGhXq0wz6WuqcI/lCHD2mmbFt8h+N62oIv/eNdnxWJRQDAB/T
qbjDejjPO7Ny8HS1kojE8yrdNiRgF4IIPYy/4xQoUfp+DX03tJAR4UArmZHFizrYA1HLr+eSpKE1
mcsH26ZTttySvyA/MtUT69IzlYf1s+SmSXB88496lfA75mHTjjDoi2UKCxt12GVxKzCn5bcJnC0f
CViJB4FFcu2ACKEFpEa///bETKkm3faou2g5iXT1jiW3xz47stNH3ijN8U0OTviODDD3Bmmz67WG
QK2i/4PzC33vTlhtdxEJBjamUweuTfaBtLjWiTwg072PKNCBMW+jn5CFp0Wxn+KDgYRXFPmiiT7i
Y+qO14z9aBKFl036vcLW928Bzjs/eSSDeiadULV45j0IGqNkIeZBLqRPbE1mG4Xazf162NQgJJ1J
d9PbejkF68XyJjGgaNMsltrcHDNvQRqmaGriYXb0F3m5sOwow3rhP0H6Xk6HHuqyTftQCiwKAQRq
D8Q+c8i/7YfqWG+MqpVV1vMnTlbg1jt3Zq4HJ8t2MTpFPFba76jYfPGgiTvzT+b4Ej8y6ljarcc0
NgUjRNCCTZswY7I4AU5+F6ORxVO8KySX9FdPhGVEcIXIBeLna57XX/OqSVvsIi8fPu2JyoDyJnfn
5OYGhoTDOLgfYJbeBOh2BV0YE9Qqbfv+zo07qvTV+7IsvH0baGGhSFxN84thl8zgDcR4a9BpKVZt
6tWiL2Sjggxu49oOk24AEENQ4EE5twXw1zIP+TbSWCTeiu7KbzsJpANI1sc652qKKXlnFxHN1Hst
4OTZ/04DRJ2PkGLRQypKmk34TXhNFTERtn971Hp1lYAExHBEHcofT8Nttugyx3zw0w9D3Ku8Jx7F
Cl0A2GzX+BFes8rLQqibZohlESxxE+kSZTVxkG7KbfEGzffKnwseE/FxYSJlulRVijOXe5XWgZvf
7zePbSQACwPN3DnCCpPFfJ9RpuCge60gNRiWREUT4ukO1u433Qak/02JIijWTjFvEHoMhyKf0Imy
ZCkm/0utu0kxZxtlTc9bBJW/sPAEgEa1CIEpFj5Giie9yoW3W8LQ3w4yQDsBAgG0KuB6gMLYDmrS
La3DmqLUYtvsum22xqiq2cvOaDkWzUF1Ak54yI3gTs/wC3tR5Xoagv3s+hx8f4e5GtmLMMJvqQBo
sLF44nLDIH51LfyWC8yNPVbbrK5YL+wTq9h5+v/TI3zJ5ak9CiqIQbi0bjdnKUCGm3Aq6jJW+/rS
pj1uaB6QpqlpaJLc6BZj8iXr1xCFu43lZrUvK0f6Nosbpi/yxIMJRlhQKUrP9RibO5iBrfkKkP+J
Ju3p8hCW01EWApP6AwzX8NwAFLF9EX/T/O/XI2bwCPN58eNwdkHucgNA/pxEQWQb2gGafNpKAr9X
AW4LQnLBe+muiPO4GgfOU0p9KLXPMg0w8ZcKwyHWSh9gn/OMPH8o9pK09gLsbrUfFRQ904QQdNGp
g5F012TqMbvY1FI7DtaBnIG/j4cbhXh0ml1Ydv3PuBHqs9iBYPEEYx5aFMUx1R2LqEcYpmkU5iYv
5tYpgG3jHyc1yw2uIbTE3e6vITuwdlTpteEihux1v6B44W/6FhNv7LBS9Ku8XvCkGNMjDVvHUuiM
WaDRPxAl32j6w3IsjSpmFHRwcVLUDxHxWqMwqcUj6MU3TIObhVncd7q+mW2j0IXK0dxiNw7rHlOI
K8ZUwUnbapUuwdR7deF+2svVrSwOg1b6jonvu4n16ch5tiL8U3dPhydZSyO7kJTEMyMBmOKyfnTt
AHUMhC7lzNefc7o+iLeQRczuZka5Lr/IbfahklPEp8uOtbjIkz+S51VT7iiU06BdVBpsp+cG83/w
xYfEtVyKYh3CrJOLA66MP759HxXhvLRu77HPvqkG1JmVXJcSASnep59+PLxapgyI/tDbVq2bqplr
d9KPqYegg/XCfjacuCVyuz+Kja5v8qpxRymQ909aLfDPUIJHg2mBPxTa3gcwple84B78F5pXd0RK
0R27LLvYFesSNJM7chLZFUiJfKGLOhDd+/I7a/uvD38g2ca2Z3HTtsIS0CdjlKoSnEATNeVrgyhY
8W+djpkfq+HOVE9NZtY2PtM5WoauNS3pjtNOdQfLlK+z9vDpmKrQz7biWD9xQgJ6ZYplIV1GttBW
A14EbP+eNi/tXMsKH2FewQpne9xn8FvXOzGoCcO9Nt6NvmIjrBm7hbl2PGObLiwzOB+a/2yEGgZE
VH2WMtfP2de+kRj9RNSQaqxLIKExQVtqYTKb7EYSfGGrq2jpl3i2SqHYo5BRVNVj4cxKbFmE5U87
Q4OCM/bnGSnqbREg/RskudkzfTZLpq197/764qrIpWK/Ct5zO0kySBlN0Ot59UCjpi4W7go48jjO
ocV4pX8U03JDeLBEBSUZoRoTnMJjgeVnOQfzl5in+t5PyWhfPCmM63erbKk6Aa3vxt8u3eFwga18
7+UCLJcwWEpFUkki0FOdn65e1fEp7uHdwRisgaGRw0hG4/J84TjzAOEf1lkCSdmGpchQSTjbp8Q+
jIAzrAzU+4+vYs3qfCLHcioQGGWn5nsA63I7QQIzECtia9KbwKaMNcUr+mhldHEPooh9HtyDjJ5d
9gZHDqTE1Jiz5X0xS+RU61SVSGXTkFlQMsULVp4Rgm9kSpSSPphw9/UD8iKvcixO0K/QuetEYh2F
gtMgvoRNlLv/EKsng491gpkBcmsqLIL3W/JJZ2K+V3YVuDcDZaLFjnY6Ba7yBBBMZpj17ohOhd7C
O6GEjqxJoF/5gvMg5Ad3d2AgWE8NPLfFTTZziE4TtoOfvXlbgkGFEB2BjM37F0hhT2V8AwetpxAR
6DeKD9kk8N8eZkOtzYGhlqnIQTVFOlB6cKpVziE7iQ0Tc2BSqI9fcLE3YpTsI30ireLrYLDBH5lR
McH6OBRFcen5WPry0+/Dts0/owKWRgSvy0W6vbDzIErmVZTaSj9UeRfcFmxMdMlBo1UH8CFqVqiN
p57mY5bi4wi5n+BL3BPfrO0ShEufPpZ/qkIT9sCBH9zWo7JTZitWab6SJD0gIjES6wL0DW6eoqCf
UbYMrcJEhBffiofjqEbkcXdTmwZpXQ9DI2wk7MEHl2CzVh9oSBpXy2rsSZG9zBEyQ1cySkMi0EiR
wzxW/arCfGfr20TGupwZDislbwdtgvuma+EVBL1pTuhwW/2h9ZMNhyDvxQ/JgDtrT9xbVV4HfsDO
XJwJ5RhJA6v4B8oAH5V0klAmTInlZAlAX3Xj9ilCvppJ4PXJtkhPL+KzUOHtq+yc3e0kKq8UNJqM
aScIB3hgiVfFOyHSY/ip48iLECDR828qNirxgj9ZqWvQ33mEYAgzB17ZgEJZ/dqmd4DdoFNuPcfO
Pg2SADDfBnzKisllN1U511jes8A2ggpufUncicbByc5KIKogK8HEEnE8jSAX0vQbaAlGuV5wguyQ
c1/uyCenJrEeGsos7+93mPSKMBsIxLhCHeYev2sKJDrH/ZmdtVXwG+xNbCRIsXZxFgiHmBIupjzM
YMMY5Vba9x0chrSojksjEG8BTFhbAp5IcLMvD+8Ctxt6ba1BkslHw5Wghs0BGzMwn+agE1uo3tYt
pMlUfAMN/58XK9xvglp9Xu7D2TKlFDdefHvWc1R9+3+LP/F0CBaLZqF2PTVhqCfuv9/1XvVvx7x2
mNu+Z1wzI1KrezCWHp5tWGp/vtErhzusr3+xbRouO/yCdpYmaC6303+sWQ6nh3DdSnnMIJ07s/tz
NOaQkW9mv+nIFMhyfJq5w4WVroRtUokW+cCOpC/CZjn95nzM+boXI0PP5pXqYQOyaxd08wnei9ri
g7WgdupFLua84GbZA2r57ZGcrbS0LkEsIi5wtF2bR8lGTLjxUEzr2CI7Kvu5A0bkkI+4dPp9dJeC
mhvhJo+wPjccLpZbl354+1JzOOdrTPa3yfJyK32MXctWKAEPEyI2IY3DoqHa6uQfFyDto8mF2Wxh
w8yyk8wQNwdnQJEXaazSYlTpXHQ9c+WBL9q1oXFyWE6hxej/bADwXxU8O/+7EEqJfs2eRe82hpVT
10yWFIm24R2h2HW7CyGeSPLhtIdZ+Pn0CrOmUwLntCU+C7JNS1G6wjulU8x8q/iHkTYTMVZ29AJE
ahlOdCIkrHJto3gXTpWgl8Xo/MliEJ6E5HpEf7GQxfcrgl3R/T5RfvVWNfGm1dqK7RVRVIEqOpAd
Z00plZVqRlqhgHTYp/M11vU29Y7FsM9R6jiqgq+evXEk9pGKwC6Dps44AVEYCxei1oEZEOmRKklY
yE6zOCsZf65z1EGZXEj27MOoiFB/r9aWt/kj2MEmGoVldiqSkDizomNekppGL+CYU3gv3C8v9fN4
AKCWhTyktwK42dWpmOZcLSD0jGS2xEkgUkjwOZ3oIN/xFMAORtndCtAN7i8V50aLP9nzsLeZ6eVz
cTvufDLCc+eXgB24Sjc4RAEhM/SjnE+LbjbVqBA9pFSZP+vamLxJFRy1KBAHPzxr4AHO5rtvyRut
5yT9FJ2COGDfMht75lPgi54oxKS4SWsgxpOkMgOMOfn2GdpSPdk/0gOZmRxwDtzQnLSB0zLpWLCv
EuJrvGR5ffR2MDDPN+8scUkc8IkLS3p8jKTGuPP4lLJSAW6zftkVAEIneQmc9L5MyKDyoHyf05IC
46AKOdyFMhay8ccpGQ8keSG2nOHuApJzlNswy6P7AnzdTultEG6LuC1XnZUof+HpAWpDanBKmfvH
f9CmNtQwUp1K/Cb8CySwcHxZngTQFJPsqCVeTziFPFAIxu6MvlnfFCYhbPEyuIwzl1+CndT8fv4V
30ECCNiKEtGU9J/idvEOkhs0HdEdacRr15D/pp/Ppi8BuEPoFfv59Xi0YByjtAbjOy+cBtNQVTVv
VS4eHU077wOoYux8i7lpRp6V48yL9vCOlsp9aVD9oa3UgOLXAU8tXtP3NR29a7imDcoHy2V7U1QB
2v/TIzn7ZzQ15oA5xMuThynrp/AM9j126Iqgf11sMVwfgnawGoMrGa97kj+tqwv42Jh582rHZDfj
E7yYM5i0hSCTqU0Nu+/meRsmEY+nZc9wL3Djk7qkLmF+gRqxK6fof51MRK7tagXkjYk+wgKAua2p
PRm7lLmTfgNIu4NZdrhpvJbOFbBe3purqzGGdLe0DZVCNL9K/qhHjfPi0laUzfA1/3vs2Tg0R9QJ
5lxju1GYudSS8r9Wtmfpn8eZI3MM2n4hqzE2QcxvOJeKCUEtB3hCHsL93nYlJ+dqXzEKM33hIogH
r2oPWBFf0fG4b4jLPmLlLuikayV4wgoLzVEkqzO9dUMJMimL7yeWCB9OcCPTcehicjZbvyG9wl6t
R8anYwcAaW1IDjuhVejDFhE7KA04lG/YG9NpW8Y5PF7orYMS66j6PoRzOPpZKTH4H11G3Nv+ZatS
FArz6SqDQ6RJsWQEO/y6AxPXyBBid7yYh93dQ7M7rXQc1MYbb1wccwRYbCnNxgFmIxM0IBrTHD7j
+xoqtLhTeSHfGs8Jgclg+e4UtUnUeJyZ9xOse8CJGeeIQiUzqNxZOXhXVX+WQ7kf+P1BIH+0PAl0
uAmvzABQhGZAYPWeJl8ViQsRfbnHqmg5RBA9MOmqpGe8E5ssAT2mQGkIGy8VDGqrp+9tVyqu1nyY
FsDEWjZMvCpUpRTYVsYOp1jfAaF+rZVtS2R4z7CyYJLACgq+Y0VNO9FbVhec9SaDFEuM8P+fUfTl
eQCowqOkVTJXJ0LsD2rZS5XFXYxJbEzljkhlnDpWa6T7h7MUT1UnDCbRjU+M+kO6/50GpB4py/M4
paAYPn+3m1eFHCq+CQiQJ23Y9dm0kFlxrReVg+LfzcMDwEHwveWO/ZVgug29MhUKQyrIlYqkS8xP
4j6qyI1UmjaiAFzUtXEtOYDNifPCt4LuvKuBLIaBfoC+91pu88d3wrB9aZM25kPMnjXbTInwH2UR
lZDNNnfOhIDG+cncdGwyyvh3g4Fiy/eI8Uz33trIC4F/CyEpesoQAxg8K+9RvyI2OTDLfsYGxjHq
MC8VSboQbyVtEZir6ZM3RKXWagkrF0cBzQew2o2S3yxV/0hLhIdA5+IXJ7qFbaSPgc18fkgsLG/m
LT5JgBoVhxqZn7/GpvmUpWpzsQ/Zz1JF1zlBeYawjuxECmM5/kNYNZQpdR4JScKbjpOlCK/y/xTs
SK8H/h7nS6MfYiuJkLK9EZ+B6jl8/xZBTTUjrKh9ai1elg9IZHpv8m77Hf69hhCEy1jsJ8TMrpxD
abhhPWrsYKWaCdDQdK5dEifSm9R1iE7NqBuuxf+W0S1Hj++M6M/5PttxyyuuQKgaYZ7B3Ckm6/vi
Yt9EYJtDO9loZl2FU33nPCeC/7lQBYjytRcQ4On14c4Tv/weR9K0AN1IL1vmDsMFrnz4+AuH8ugZ
zHwY4lD1OhXkA92UkI/gyHPETs+LHVQkGpSjC6zIUuP1e2Sz2CPOguo81LI4Sg2nVG1ZwA3lGuEQ
aQM6Q5l1JNXE8X0ttXtEYi1jI4AIF1Q/ubrdKgkUWnMVjqQXHj/67lItY9AcEdxJ7Hd2NZ5tytSV
2d6sXrGy+EbxPxykk4V+XWkqRDEPvOapKjgKBcdx5lhTPBrNHu61HXmp73QLXNunsTGp5XjabtDH
JVIYLzS4KXNuONXXEBOtAn+x0HRXuDhNwaL8GAea0mYQFY4RMN4JKloBPh1Jan9JK73DmhOsXSDT
BMqbAj51Qpj7TSCnqcANYhW6xGsSVM2cRxlPLgtrpz+J/FfxWpczPXp3Vkq5md3YRLSqfHPAvTxU
EgfzeTTZww5lnYyJTUN2gkF4GQS3IdNhF67cjZ4srXfi62VEx7LoosQs90/i9HfZipOUxUMsZihZ
8Sie7Xv47Og1qmWI53RDEPrzG/KJFhdbjOyUvGF9XVYuKJi5UfLPuGx/V3yE+VMikLbLBd+T7F9B
ZkNdmX0xzUxeDWDpPw1GPUkxG+W2RCWSHw0MdY5eEyQ8aB2XQ8En6iDniirWviajjH79pmq2GnpO
b/49KHyB2y+YVCZamwbsGyiy5OWrcTycR7SUaZPcee2wxHGdp11apkt7V2BohCwOfYjwqw1HzI9C
QiDP+VrztBOMbx8nyRQlNxkFkuuYPOb1FTqlSsQFT0J0Th5CJtfb+zaGE5jvzUtKq3Gj7TYbsLZt
ZlGPW02u+z3DqcGqGWxb4ko77Yti96jSh2W42yaJPzcHvXwAy/vaYFiIvYS2gdvXbQYwR6FD022m
mJd+FyLtbRTBUeaI9J+goXLTGws1wgKeDdOiuN/slCnziReN8Zn8mOQOEDDZdeCsSJfAZpo2j6cv
KCBuHeWhtKYDDh2T0JYmM+XyH7IE3h9efR9Dc8+AXM40fpofjPKok/8tzamip6+BiXZXmYDEf36Y
aaRj/za3u8imvg/Th/2w7cqgt/zrIZh22r9hElrE3d22NojiQYSEt8COeYs/nbSo09p0BpK/7+VP
Qj40M1tV3vO4uMfoEe2hD35S5n8sU5a+p69wRE0RRfiTvFdodWiuQMiGJ5YNvRnUJRxfEc8ciPLl
AcRuR+j2mfTg54tqVFKoxj+C/9vrTmwjZ8CQ6FOfotst4wK2/lotpaddG278ex9Z/sUAdxgYomEr
+DiNqWHCQwowBz91RLCLZZDOdePthFf8CrHgtlWjEh9EdYekF4ZYKXE/cAJrPZR5H6A0OOIVIXrV
oddt/O11arrJ/yUlkZK4ma55IDp0sxU1hfUIo5wmHh3ncZbQNK1pXVwxKd9WeNmtm7NcfX/hmFiq
nVdWWScmieep9RXh1s4lTg6MRuvuMbXZ/1qyLDLJc+VgP36hN8hBOTD30hEhPUyxTh9z86uRtC17
dYcszFkxrBSDd7AH+mDa8wws1HfK864LihbTdwn00zEaVJGmeQ2w3twCZVzEvMK3c6BBnaCgp36h
h+LyFp+FFQ0k6twnbxxTJupDc2Fnvfom6d/eIsm4NBc1LkFDvU+DX0RWFuYEWmB3NsYLPxDotfN4
8poPeE7paw1RA6gKQKkYlWfQ6+Rr8F+9szyOEufOl1y6LaOYaoqfDApgsWPX6QmrcwN5WLJlcIuR
ZMH22JEPPjo7lpWVWsl2MAgl9gUsN0RdquRoBKH3cQgPfO6bjChP8ZpI8vP1otTz4+NfvESg7j7a
1b68/VUgNiJ7O0a28WNy1g/K0Y0m6U6pp5caupdppaLBJqQt7G30UZTFhNadmkb/z1ng6TCdUX5w
EXZc5Fd94z1VUGt4rMr94z/dVAEa4gOJZA7YmnhTuJB3BPSIbmyOFB9RviKnzj+NcC3pU6a8ipUa
hQmEPipAiq+29j4ZNWyGajavQRE+oUxnKVSBpDv6ZAt8PCmq1f5O2Jafofng9PvcJ/NBMRRUcND7
qLC0OlRdqZ5CUkwJ+z5VhSFzF3zAZN0rtPrPOOv9Ib9F9kGp3bcXGndx3jbws/PgfPkX+/2CdQiD
TwqwYoWoRD1q470z7Eud0fn4v7P8N5YWjkKnXXRiHYsxLbSmViLoqKXY8BdcVMcMo8/OgThcZuVL
ERPUy0ZeIZsOIWdGETtLb64pyCZbpjpGzW2UsStFREafH+zTR98pJeXZvBRcaOq4p0FTwYd1KEU/
X8L7bnHbB/1HPINpFGCAlrQkgD+Jku0diEU5crW6IxufIGUofvmUS04mqPuEUFQjSmqKl1Mw0Kmb
I5s7cZVITMhN9OROpHYFNRebU+gf61YAGSusV+hEvnqnA86ZhYakPiy0HuKJPvHk0l6w0H1C5L/7
wN/jlQ/5dVDd6zXUoyyAFNnTXEeZ1aRpkk8MLgm+G2p4HwZDWJRHLV2Dq0C7E3YVT6BC0Km/OdOj
vxqB6Ye2NoUZJ38RrEZHhfnwkpj9NMMB2d2X9M+JFMKYFpp5NqWaluLmNh14BXe0RIvRinqfNlw4
AGDoyop5WFhg/rvATLrABvn+5sOLzWp5GAAVNccTAzTzuw+tMSGs1ahSEIrxZzdfgRPrabwKt7eK
W1/RxnbtzLTuBcS0N7mFElx22Q473h1Iwm7NHwQh3FpC9XgBVe0q8HY4gN0qmEt9RxJAw+ZALaSD
gYWnWlfs4iwzR2nZZO9oXD1/HwOVddt4FHKKLGIXAyRXqeD7YTFU860y3NYNpWIxmd7VM+DiFY2n
ykzcbfLSrb4CEE3cBzVIvrOm+z1vggNKjNvu7yGq8TIBAb1OZgW7s2iF5wwpBc5sl7k4K6HgET+/
6vGKc+KADXt+ABSTV6VvjOZqBV/ekKDQNIMpF1/VvmjWDwlmxFdlOJWYrV3pO9Mi9kJKIo+rytCo
o77we1rBBUY2AALMkLoJtoc8Ud35wJjcG76yh7mQgO9FbeRFymw7EUoiETviBqIH8wYnTW28aGBc
iwJ4sj4TFIJx1x9+eZ85vbu7Ky79go4glapmzUoD5BCXOIokcA0LVRO1Se9IFk4wv+PlEgPDJJjG
mlXwCjxAqDe3JsRvOBolSEJ+/QwrEQsNcuaovjUH73PUWGqBSfCmZBsKcQ1s3f2Ho73YNXbk045I
dUSxQSIkrwdIgNbXX618SazDJEE7P26MBrwDq1rUYnI6jIRkdoNtfpsGjiaVMSsY7zJt57lPmx9k
qEiw+vq528WdDEq/LUqaFBNQ536LUgt9wniJsYr5Dc5R4bNOVDRpPJ1BMYaLsDtTMOueIb7uMOcy
jzPgz4leT1Hj0Z02JAWXo+U8ydFiyCoNet1Upt6QUzE3Y1uNt14HTl6jRoHOdpLOPxGHnyGn6jII
36XtynNtsnu8X1TrkEZ4p/+AzXtYZ76fL045XZgmL5+0/c+k/zDLytsqhoJy6f0kK5d4z3oRqec3
oJeokRdK0c23l1Ku5TrqvCqCu3BkS81SQykqub3S4rFaI0KX3VL0MgRrImhS8yyI3TLcqy8krhC+
FkU3vwWJhy7dHAyTQP2kVfiTIeUN/ngt7u7MaBm8N7zffWv2YfMOjcokEPkGJJaMloLvqFW8FYgd
Ig1GxdakmiNkDSbahUZKpKUg08nnXsQjGhcpk901z9bY8THHT1jX/9JPG0kxu/8Gesvz/eU0s9nH
m+7AfXpRyymDskD2En63yriH7exzt4u+D/WJKFkC0LUkTWMVmQ3oLFdf4nI7tLXaI6FRshXsW5Hn
M+vM/qUFagUry1cQZngYp+IpTzy9oVLSnx8Q1FOvh3uLFMhswL7xx/G0nlhe6f+KRBfp4yumYsIS
cwLormtOk7FEINplUJTo3eepSxrud8BRZQrwFmAZIa+xKBoaICMbzVD+bk3KHIdee9QL3Dpmq3Hi
gSg3yHlVOhgMvfo5atTnGCPtiIYDCm2C/GjbEdWYUsGPZ/vrMj9e3dRIRo0HBXqvfYnBdo+TdV/n
uVYsZ6SwyhAQiKyGEN2qO8haOYtvzO6HKHpDZlkcUCIcpuune6Q5M7rzXmKkWqKUTTXNEDPqw0Bb
CqXGlB8QlboPwSawph0kWQyw0yywPDAymk8FxtD2bRrb3U6WhardSDS1doh4RARvTKS043Tzuork
gD/ysNt3RM2rdwDNtv1piK4Lzj1HJ0xlX0b1krpNBuI1PqxndIIWbQEyjg2PcTYhWoVvxFJ2no4V
w1UXmSDUTYZApDL7R1owpgDHLb3wmoO7r87NKHPZ/FKsOoGQgA26n08v9/UkYTV1Ngcox36DMvT7
a3WdCnrbOCqx2FgtDEzhuisoygsKwmOlo8zXViLLUcNs5kDfdYuxBamkzO4P54xBVbPe/K11U02c
18UHRBVe1gqnCvIhm5nqlbYCOR3fv9aCwWXLOgfZAblnPh9Tn87GZB9wzhqCgE9TZO1Amz802kO9
FR75PonzwTCD/kzvXvqc0v5FLyWlS3e5sGryekigIj9sbsPjgpvAWYVvd8KlXu0oXqH+xZ2df2+X
wq4VA+ujA/uHJ27Mm8Epmn4FlEYO5WZ4fD7m1nTMIBp1CDWTgvRBP9Y0l1fQMu99QGzT4xF4hwa/
HhpBuvRLtrhMq/iYEip4Kvv4okzeZs4rJH1lcaqrKy+lHSugIrRPTnYEQKZ9khQqasAxvOEKqHUW
PDSaHBy2iOyDroZZnc4tJ5KmP1AJBgM0BgH833/PeCimIwS5+HpfBoFd714DgJxicEQ1h1oq/6Fa
FsqjQ7DB5YGqoY83lRDcqcnpcU06dxtKtQB1M25ZIDb3Ez/+KQqscxWHMTKqOIrB81lVT1F2SLIh
AdP+IMvq9i2+gFu06VrZm/wKhd5Ha689CKEFxu0UOe7Tnu7Ee5KI8d/cvLCQWPswqrSH83ddP2CE
uG4+Cqj9KVkFZNYUhBRqBiutTyIKFLVWdodYh+grIPcDZu1pJUPV1SDxsiJb33hRUcqjnLqjlVbJ
Tzv9l8cyEfqPVShNtdBFY272AhI4imF3l1K/G/XARlM/54QGHHIuzHoj40NDxgMxbw5cYgXJt//6
9k10hBShq9sAQcyrkctVIjL6AsRSXncuYwRdfALz7BqqGap79om7V2wp29gwLiUn6VeFXfdc7hok
i5BQplEsD2Oq4Np57xwgGwn5SoIgiT9RI2Eh6OhGbd2lJtsKduTxRhiR1ah/gSZ0YUg/rrBJRGMs
kT+L5dsAbMuzdV7sz45cCoDMrj15FOiD0ps1gJqQhsxv343UFpxLF9tD9CYER8nLCGwyI7DNVgaR
gMdKO77RnLfgSXD8ugGBqkaSRGzOh+haLx/3k2uLW/7Ha1HHQVJUP3eTkA6VL8HGbvLPXpMviNve
nIpZaOeupChUT56Lh/N42zOixZZAooLCsX2zEaJzHXs4Dd0n7oHlusbjIeUiob3gw4uK3zAYwEoc
PIjxS0klc2ND+og9gm6WKFWBxySKPV8jku6Qnyn+nwBRDaRbCzhkckPToHz4CRUlde3N5Ti7J5UU
IW0VFaHF95NkgyGP776IkOHRUWHY81zIKG5np4L2bLMgZpywCasf3QWWo/axfz5GLWJhCxvpKpsM
vHEX/0JPvqn7n3NdCKP3HlENSxa3nPgocpCuukdTGBt70rrzkbAPp2BwoU/AzFJa8rTOGS1O2e9r
Eplt92ClErcI5l53yaYV8o6mZjLlqu4vxhcIngT6CbGuN+iOhQj0VgIxHesLLBZ6XlLhoH+E6ork
Z3AXKzbmBGS7+RLi3hdFaShDBK61PVcJIA1Lb+9f+eGxXdV5I6v4+U7ahPp/ZqHLtHffV61W4+KU
k/kfAObkvJKgRffYPpatjYoK2qIziCfRlbOzs2luHEPO1fgVIOsCt8Wnqj+qkBPjwIhWjQzgolxN
hWNEX/yxFQyfXOq74xbPt5VgHaHLLQvhVMmK8p5+dTXKvmyN8p5ee2VJT591L+vO6jOrrr+y1qOx
Fq/oTNkB+t2CLAHE8tFo44eVgPpCXYaB4qydmVeat98NetblvGNXoh0Rg+OSNDaxSP0jeBZ9Y3Dj
uKo2/F4Z1PKSmjNP2bRjph0mFluwdZu4zRnOdt451DqQSGJTkTDCB8hfCWyi6sn9nQC/VcbPT7N8
MXVYWdkLM4QhUkIfdh7cUJBYxZMIFHDc2CY1FPURMQtRdl0Ll5I692LCwH2HD+js+s+JHMSDrtQs
X7HpZyum7BsNDbTGJv2lNe5i8WQe5qNq6KP3tFxomCgssaPm5lqxp+gBgmcs+anX8Nlg6EhlJhZq
flZfokwvXnPWXRjxJPOGRyaKAUrpoUr6HF7G1fTtQj1XKJarWZT1wGk5xFZJEFG9uMDYnZk57LqT
qJdQr2AV8PKKmk02WFVCnXC6GwmYbeULrPT+BqPIkVYldDbw4GUfuBrtFuWWmcOmJhnNg1v+aDP7
bgXaKjbORhDPh9uWkEzKQfAPA6o4viG99taqYmBzqnnjoNcKPtbpWVyKRfSXdT9+DgK5UzEXrQ5r
uqxRKzoh3CqeCVvTTTRqyAaDjLMbkAOdg3P5bNFfgXSRWhNPuz53Ub8G15+woW1zwccmUcFZJxi7
J7QS1CjXzJwSMgZYRE7Du1x5kUm9iG9XI3sYKrBzxTAtjYMZOYp7Xmh+e9zGc9K7doaleukerFAp
HO9qiwdKkf/2wojqg+6/hRs9KbMBq9RqUuqmc6X55cFRZQYzKsY4KssiYek+XqHrgZ3p6+uIkRpw
6AavTTgJWP+dYN4CPlXZKLDEdUvydStssMgLy64ZDIlCTDP/0lAre3awgZKMaExzOUddsHRtsfRC
lo+L2qlHp0iKHdvEsgTPAzz6Ham0JwnvMyBWXTu40/dXV+tWHl2JzL2Xypv86wwgCB+UAMZTtvt8
TwHHvgbNaPGCH9st7/wcstZMy8Fz4GtKeRMGGt+a6clAmA5l78JqMGvqrXcCp4XLA3H91wRDWK+8
T0dFZf8DoFlxklTcq/RJBzqjraAjjgnQz7D6PT1LA+sOXDHpGMTaZNotY2wAy4W6T89dLGIA9SPr
cwV94HLNHZOVyHM/Tx1z+CbhkqHxxseAxK/QbfXcca2wznEfIzRDaT+ZfzrenB/F9DUGH2OldCe4
VmSTqZ/NhokC56OHUhO/ug4dfnvWa9DHieQOn+ZZmbms852RJAspNalOAMZv0mK2dSluag5+SvBS
bscSoQujpVVNnQSsf7agWFL8y+eRaQ+BeTnzm0Vv7+VOWU58cCb9qAcsfJ7maXhQ4OP4mGqJxOCL
38kx1fRKdX81p/Oy0bjAXengzT0ELe91C8B8RKBDeYDmLSYvr+A0RSUdzoozDyuOKJ6yPBo4ycdJ
kblzrLgl6rjicdygIeUDshTii4VyiYk1QCuhjYUnvzFGLPGr6S/Oorxbr254g94Xxgm/KyXKrGVP
1wl+CRZ3JpumL65MXdwaiZERRoOVvNgwmc9cj2E9XwX0EzzhRQ7rnt+vGYjT5QxKoxmJbxZ5MNKg
NRFH2WbYvBvkTYwCrPBLRUUBIX7EcM3sYxQ+5QJBJfJraY5GDzSN8GkP+EvtqAqfyJZnG/YJIUE1
a9qLxshMsjFVOJ2Cvmhq8TfB8iNN40kCAfVvVlxzB49aOyk3L/q6HOMRU8wCaLDqScMJJvL3CdQs
PnymWAtl6w31Js1hCEb2rHV9HVNlco34SviiftnzwxtX4ZS3J0sSQBV8lliABR9lW25zAZQAuu9Q
+spIgrxvoRjOgBumePCnpYYFxH6NMriHp+vEFvpaoP1LF1HLJJapXjoA6tE0ZuGBO03sUFIS6S8x
VUEpCpGC/Q1ku9sxcixJASkvjhsgLD95mnPROEiYn425aJUQn84Op58pEfHTkg1Hoe12v/8B/4iF
ONN/Jm6QR167zUA5F6HnJVqG2SgZQ54JTbnALAeEusK74QgGAgCSYP9CaMysiOTa94m8FblZNRSc
yQtIxoRolSbPhVMUfQZrg+duUfEDqYOA+s0ZaS4YWsnyW71uBABdSu92VUaMAnyIh9R40SUPVMsd
B6Q8vG/pxsJUfpWVRHNJ7Xtvt0LWyDn3pebjVtYwlpOhgOKvrzHJV32G44JgiyUBU3aWP+7OiWFe
LQtXfywaSE7JqDRcmAQ6NPKP81RIqXlYMP6fIhWknGx6IpX3uAmioYmhqJc8gcuSZX1/9w3UJYJs
goilKcMsTDN0iaG7EB+rXhlv8wmShSi+ficLVL+BwyCX90JhGbcvH+Rmc4ZuQW41XKy/38FdJg1l
FMQAegNSiYKbRO0pGnBbR0U9rD6nZtvnxaRubKJpHVFEiWAfu+uImX/ygzVDvwDmhNM/B0VUTcYe
or5TsMHXJN3dmo8WQeEKHE8ng5ns8Hw1ydAeU2FwNVoXt1IHXC0O3oIAWcsh8Ytgxrgfn3m+8peG
mDMIxyinXjCZay/LzF1ALQwozxq3Be6BUMwHRXtKsUaHnKwZzBuX1S2HuJjCVV5EgNlHZbzJHqj+
Lt+Bg8aBQ8yyoOwp+INTVruVg2cX86EAgjKUNP+gsM88yhobT1f35lS1o6VClSPPT2F7nJzr1C36
Sip8yBya2P3PQEJqfi+ATooqB7vaC5Ydh6fhirRGOIZWHpRmPNa+bdNTGhmRACmJRFf613NAX68R
yOibUY/x8E37RsNbUI34hCSWSaw/UrPuAMlzuIbw8KJIBG+Cy0Q6cuwx3CJfRU5GVRleojh83uoa
svfi3RX+PsiadBwic7z9T5oYwgRjys24dEGkn9US/OUmFv5vsSdkm6DP2CKtKTRY+OGJDpGKICHh
KLImAC3YKyXbD3ZDjEYy7vo5jaeWMZFLizqXBTjEmhsu+hkCEWT7LwxCt4nQ3XWIRwp9eyW/tMuC
IKTmTLnB3rzK7ValTaNDKagtM15EUu5ZyqoWacCJesP9Uz2zKGwg3vKhxm+M20AGSoC6c/1oPt2x
O2v2UsCbX/DUUIhIzVpRRYx5XX6n/EXkHPSNvHVcACxjdM5zi5mT0Smj8Sfm87i0j/1ZbvJ7ew7e
b7EdLsHSeqY4UG9LW9N99JVFS+k3xMpm1qZrpiMhIYqMiQ4SUU6AAqmGUpLQhv6Iyah0/dEKuOPV
UxTfET6Nu/y+7YyVGJqjGTUDeCGeXDmmVgYFYUjfug0fK+2zQOzD1MmP66/sOLpd+oErL/zSsQoA
bPd62LkTiIBrAnMWbXgmc0eehum2gqDUb0fatOCTxs2EeK2X8dtF1SgXnkykO1Wh3ds8pa4Kh7Xx
eKfW+NdDsbUaOOCwoPfPgjTE1389Lmp+JPTYeqAUOx8mFRJq+8EV6hq5AtIvalRA9nDmTOGSUsfC
1ggQH7z6gFS6f1dK1DPq1F3mUj4ZiRLptk0rQvZl9yXMFrCC2yifkuWLb3tDi+Q9t0WqP5kWlFjp
FCt7Fn43k65Pa7g4ZJbzhXPXzeK7VpftuEuL9bI8Xr4daE342LEthIs830VgdDWY2zjzgTwHxVRL
XVKaeGLe5RlKnlNIspVuM+yvsCQQK8UnYIhlvj5sw93r2+6kAncCYP3ygJafuBrsEov7i/HQmNxn
gEOEXuBadqdGQkJNVi4MlrYaqoxOEd2VSMiKWSMUorQj90iXouxdhylk7IoQNNY0iA6RLDxMeJbY
lQI55w/R1Mp6Qeiya0gnERkbubFV9f9sFVXsx0GAQSWPXo9tJfrISp74D82WlLylnhI0LeBs9wCS
wXk3aWPwEHFn+U72P2p/ddAX6BHlKB7yYJTiOj0Uh9KjwO5bcdg9xIL/UNom8h+dyPTYB5c95Ivq
Do/YZgmHWrU5ISIwARP3/AWzc7FdaAYdYdGM7YnmSZZXifgu1GSgJY7WSWts/IZ+AH3B2a4ELT1O
XLqH1gRbHkF96uvHCIm0IZtRfWXoSUk13ev3wyOWkMDeQXfRUSQTy4J76RpwkjmIflhX1STuqdre
tv93Q68yithE6CXX/Ya/k+2e6f0XQpJ4v8Mg89LpvE0k4VUMJvjjhRbfUqvSy4nzCRIcnMVDrv5a
GygLN+wD4NhCXBfSV/CR3qlbRmzeH4+6HKKn3FTZY5eqUNQywxo/5cZAP59T6dlYYHxTDFIlJ5Ub
qDBx4kmYwzHc4jnHH0wXey7WLmdqvSruTSxfNPrL/umfULWaoElefJJpBFhufuqaKVYpzUjeUoPV
R1C+XN3I37JtPKHz9qze7MoOoE27ZM7lKuakLAcj9K6RQcqXsvWCAU0gdwfg9JwDWS7UZVyspCtb
n4NvLj9VI77NfYuBJRNUCv98OT2+EcpDBcpgKMlS2X0eWArJE4u8Ls4k6xMumQqP1nxhjpTqYKep
38njmcUk0gNcv9n1BcL8KHLcpjWZIJb7CVCnwW3N37ijfDCkHgIiypb1p0S2nLjzVgJJncWDb1Et
jV/FvTH0ULv5siPNm/1N4ttmCk45MvqWgHhty4XIaX4S+Jz4TnXEv760A9nLtNdyFm99RQkCYM84
rEKkgoF/KZcgWkwbZW/pdSuK+VWak1+B5sbV9u8M8p+47eQDbYcwfKXLqcIW0h0l36e9KDzT/UoU
qlNbjyZNYWKNNCarZc3H/V0T/CZ56qbEF+KOn1fozrmCOA/Fq7Y+SqJdr+HQc3MPCZ5KCRu55JhX
Xe/S3MtT6AhPYwEKEaeL26ofVCWojadbjNfzTla/Js4wrg+HD/wtjzNnmRRoezAn4555AXkuYPgZ
7k30ZX1FByt+ueDFBLmpb5mveXQ61hbFimO6AxENoKCxz/9fF+/cJUb4MC8w9rQiYl7gH36c4+59
qTk3XzZII5qXUekPPyh+hCmwkJ6Qzm4ePtpZiHFy3ZqlTv0uHBNVdOHxp3aoYrPO7B5rBEk/D8fm
u+1W0wHl/Es651+wp1XK9jxnIM+bH/o4V/smKYMGihjapAVT9U++IX/UtkYLXJkvvdZa7g6ZuQV3
YYGvYJdKcGMIcLHFTmgWQaVLYK4jW/Ungw8WwnsdM6y3F3lJL20Ff2u6/jY1xTOt4xlC0LfTd9k5
pEMWiqYTbpa0WkSKGVDFtajKBYqU7TAf6qbJWYqbJJgavvv14ZxNeiqKcDDzSnBiJIkG43YkyM2b
hLsXxMaoqwlELZUGqH2WHamFh7/mnuKeKqTViLeVx8iqhZDcOaLRgLMWhE466DDdZfhS9u5b1QOC
quEke3JnfK0s7h8khAjzMBjPreiB9rLjkKR6/XMd95DmGLAPP+BA28bVYVDg2r5kGjeXhNZyb/PW
Bofn3nUsuZUKXt3Va9RQTXzlulbYe34RubKgr2Q+LViw9l2aTz8xHLXkHMSjs5iX//iNuDsHxok/
PHnNyDNON4NWXarklYXFCWPpj0ORidf36RCHQhVKL47pYL31orILEFTs1FqRUoHx4TCq9xg2crDP
/RGOpNBCJWzQ2kC2EJb49kcu/QZjdBREeDlnngHJAwVqZ0CZYcPU1bUpkHGgGYbC8jtcfV/EnPjP
WZ1yWiSS+369xicPAR6Z5zJMQqG1oXM61cuI4K4YEkx45aUEd+kXoJo6DB1DLhnl+OINQcYmH4Jk
k5cIX+lBTG6VG7nUxOjsxTAOIuggbwdj3JL/hRy0HH6YCOeIlgzZiNLwbGBuAEjnkn/P1BS2cSnB
2aJvUNv7fv6XXjxjFLZcre0SRcaum8bMpggYv/U0lS3ZrN3xhdzhnTmTkBNsVNxZEAAJDe/pB7Fm
rKq+JoN9y2EFtZ4O6037QSXeMQYDCyo4TG3ct9mNbqnTFaLkHHxJkren4noL/XqfRk5TzbNSf/0x
2Gkxg9CrhttdUpR1DEvyyQkw2GYd4rlPI9fAMwToB+XwpoQnfawBFj53Lv7F0SUdeujOGu5jsnYd
hximJ9Zl42dQwq4Db7r8uNhOIZmB9KZNOaWiqhlZrgHh2E6YcMlrNaZimDzb41NtuTO/+G1XRdW0
tTtoxzm41+kLiGE41VUpQzEvUTeMSj9xpjx+UEkMFYv/rMQCSQ3K/7HeCHP3xbnemzFjbcS4TUCr
1wCf7MNiRts8LHtFrBx4Mq/HCaYjtpuYAE3NmgxfCQQInZkCodT7uxBv0s1LMXIwei8Il5gN3XUw
nKkwM086+E3TwUjcqA8WPNvGr+cnf+bMipXhNi0eu2j0SrxHE+cKoImwHHD1TqN18rAv7qBzJxrE
JGrs85cYB1jgoAykjV3LAjDc7lJf4F3oFTc1iz2Dz6jZkhF/TiHO5KwFbpJ7pB23IYWjXaSlHTQW
mH8/hrfaf53DKmWaw0lcgeBMl181aSswWS8PELDPCYFNosecYnEtDbG2RhHpXJcoS19RnQ+38EHk
A8xC6p7KzJonbEJqJrq06skrShZtLfZvHdnLB80WYs9rz6tN5TmW+j5//ZzDeD4a+HOXDfGGBva4
DxzFk2ugo0d5d5ye/OtzLFYbEZaoVULvkWzSTCcR2k3XB/PZowdZNLLuEFyKPzgZ4q8UG6m7yH0I
90tSmxJ1K7AzZXR4Ixt+CGhZHukpVC5/xnWx7VLnTyjnkfXIhnERoWm0iDeMhbbGzVSFAEQ6yV+N
O5RFzp6qEJn2VWjxuznti2pxFY08MHYWJG94DUgfk8TLdU6V6z/tukv3N4hKxCXl2i+JYGnnVNGc
hLGGwb1ETiFkn43zym6DZlWpXH1lBJZmeFfK/uMBXL//WF2qy55XZVRMV6g3v+QOGiO4XYTXx332
1LXqJFFWuXbUnKs+ymYu7FUnbZlsgnYi1LH90VuMOcr+6j7hQDe6cgbau1nlRn6dyQNjff6Q4SS8
Wp1eDZzS1DJ9bAhaSS75edbALb8LV+PNsJsLSmj+Q+Q93iHMk4c8b3GOMMQsUuMUQC845QP3+eX+
D5tJtiRM0BOCdEh6lDCTfqWwgSz3zUl7RTVtuGLH+V1z/uzUgBmxZIYOgJ/bF+pora5NWwT23UIl
m2tQvXTueD25tc4HWjHW9sRvgcCIIec7Fn+qacdPaYIQt/muuNSegmvXT8PXlST+zqKJyD6wpDYj
dPsRG6MeQKE1BnbpCu2hZxEFEL5rwK2SXIt56rjaZ3JDEq9KlY1kgWKRf0sQfDIgEGUWEf5e/nPk
j8UIwfMNN59ZR0xN6drR2lrlNmc3KQbFx8WT6KfiuRrcIN20wNca2l6Q5VApqTzHFwlho1SOvWrm
K81VyOUH/xHuDWgXSfIzraGw9w2ANEbH0x8+PhgfnQBZyig1S//VJ7QHjHY/7qV1oooXbjI0pukr
FIz6OKaOxljRoUhzwwQKLYoAhPQZAJzk/wtu7K2JLyyLCz11wamxTZ4iMnxK1QdUgWAvLOAJuZ9n
mgF42GIcSXnrbpoU86mb30PcsDTjwC0YgZJ7XKdrJfN65OHVWaboCVdjuy0EFfGVgcAlSN/8fUs/
l/Dpzcckghw3cFIdEGunf5uHUDjLMD6VbDTq7RjCXG1v9ScT4s6iRYHPLrDi/KboJGRrPU1ovbs0
kzY66zo0kE83/vFzOeARghUcS4/Lz1NdicyW51Nu4uheiiuXJsAQXKiaTES+nCUOIHnS/9txSMl7
dOufmhw+4dLj5CETDaWH8DTUOANW1r1NVuC2ac4GSElTfmfiXyy/Z1XO370S0xbH/qbgpqEfhg80
0KVCfwqYp2UhzKjKKjWD46BRiYp3YIKs1DUx+Fj5e8RFhSwHKI2KMJoo26V/FzN+FsmosuMVKGyr
A00CdVFGYeub/ZsoAT+51qTxr+63dkJtecXyCn6dPLD93O0RaxOXclEUh11EhF7F8KCuvysEg1Fj
+XACQ6A4lbxu2fSRq2u7mDYmsHEB34msa01y4dXBZyUYrHgnv6B/9KAY2hr4HnHFSV+lSObzDdJb
tA+wU5/cD3xCf7Bk3/4blseZBJah8ReOCAiZDVZ5JiK3nRI3ZFwQhpAnKEqP8RLkEcUab/8EZFqn
13AfvMEpsSB0SmO59uEvNpZcOznIJHGcH4jqKe4scMbcQlwtEuPCx6GnPVdbqkOHkpOr/9lkeQWB
Nr4qGyTYZiRLjmHZQoFdHrYPsynBDRf4SNgDenbTH6twPfhwYR8a+j+uspamBK1QwRuNkwkgafIe
WECi4vvUgI00f89TCGJaD6EGwiJ6kOK2GV8R1jcBvegdizhDhcMi5qAH5EaR/CzJRU8LO2DLaFCE
Y+kV7V/Jx1o8QRsPWGM/Stte4nUZy6PDWCVol48/qS1rQ2Xw0H92Vww6O19TNsH3O/z3Bm/1Mhin
hPz5NPDSQmLU6vYnx+cBfP4NkfWuirOkUllkJ8+VCaHmZ8p6jun6/RYPVUwLla3uMa4X7ZhIMO58
mIIMNpdU6j2VQjh8+SwYBJNK0sYh0SL4jKrag2weg9N8mGrTeLjd/SsFuH1/8QNtc/8blC3c+KAH
yCRjpJ4/8Sa4T88iqOy72NXB09SjzfIFb75G8iM7M9nlQD7T7HZkmrailMR8tIGVDfMZX/6Gkto8
kYTaKAvYK3ws9+whJFJfYdGum2ZGGuvwFutYN4Ek1qLOYqJiRLaKQuFHQHzD/uVU0mZ4hgpunWwU
iDC+FjcWrwMrSuK43vPRl9kTUjxAzIoyahqmDiNk+Edio55r50EhqNdRKCC2a/nUyDk5BqAIVGQy
g/ACeUCqYQWzBgz19sMXAEEijitT9PyNbNx5yQHgjYCOadR7zzsTHGoeSlnTgv7pWMRzY8fOqZgS
5MJJ4UJ7b6ZHFH87cCVq/0ssv9tibXj4J1T8HvD8ecg3iOjA3XHdv8lTk/bJ6QHhE36bG0cu0JLq
7B/ebDaQN6UV5Q+J1oEJYHjr1qej2i+hLJRdx9oW+PDY55GirDROC/klZaJ60f1UA5MG1deIMQF6
TP1WAOL5BjiSh6zsfzpM66H+/2BIykoExkToci9h+2p3Gz4+rWHI/N6ikHxl2Bx7LganVgo+3kCH
iUpeJex4oVJL/kKiKonqlH4uHApJ33Xo89VkLqzgwsc3/cgVNP1BigbPiIJTtPZGnAvbopuew948
VQuPcpYYWuQ/1Se+oecYvrtXDIk9br08kmmUPuJjD3uQrUmFjRd23DndIRl4x4RcVQg5ZhY4TrTH
SqeOL/AIkrC2py6v66I/Fl2D7siIIaUacHu8aPNR8o0Y7IE5eAKI4c41O/JhuQPFKGE1p99zZckt
mjAcxnyrSAJRjdpOohA4NO43ld5dv/iX/mhziqz5E8UvX42FzuSlMjcC8mPa+QbqIZgnfu+jsTEr
0F7q9NsHnT17C3Ck0OG6VBzx6TyT8qQTKXOzjwex1FHXrzHKykmXSNOG2bgPNtlzAXDldtTD0Yfc
z1Uwi+YgQzmynpGe+lXQ1zGUiexZY8aST3xCkwv9uL9yvcOWYYQERcZ4eve+sDYTvJeZ4uApPyWM
cJ6Mwug3qApgrZmh/FOglIr2hE9PSBWhZPAtv1fcHzcKUVTaEPDE0GfRKUeyw112d5U0XD3hDZ8u
JP93KR87UsFOCYydXiZdBAVYLaXFtajQiUr1dRPt2N5xAuZVC3nHULmdQJaYfAaodjE9FgiWnCMr
azooaJWMXcI8quP+xl5G1oOh6MLLlFIXEhnp4hnga+upqFsreYefqZrDnXw+2qFYOMg8rZiHEzS1
+3RrA2/qi7K7QaApvolXbCk2Zhchpu7iE506Zob+2Gy/5YV2gX6dYSibFJ7+UbrFgbmeattFTYLt
QgUKUqrh5Q48Q5T5lurOddx0KUf1l2UcjnQSVf4TiQT0FdrdT0Y3gq3tdcPlC4kOcyLCbw7Dk2Um
xh71yKKWcfDvIaYaOObb26Myvry+B75x/tyK6D4W8PikMR7BVPL4Mou9hYicssGjxxLktCbbsXVL
OaxONxC6szxo76PPrwqMoKgbMIVFRsAGVdUZUF+hJ+Z/17w7CspdToQYi/ZDhctJIwW5nzT9Vhw1
wmmeBqREltJB4/MQuRuJo7GyNgYz6eh7HID+lOhrM12PXv6LNlQGtbpEMd8Q9fR+1uKkVPVKfvDZ
brfu44+c+niMlCCOkpQNcN4llRURBnS3Wq/h8WW3EbwGHpm1brb45bsoKrn9VfR8Qd6UiVUmc+VZ
KyY3zUpagmpYE9tTLdysxnHFVni9ebxHJX7Twu6oceZQ9NELe0AJJEM8V8DC+jxms0dlDvLaw4Cs
TN2Oy2GdymHFbe5+REVfCRU049vwviOtn+2gD9ATB7px82IKHThUoBjsBH/1tCE6NVG6vhYVY2tB
dD46bXjY6v4Z9CpaPIP1AN290rScLxS+Fz+LQ4YqVXHhnzlF/tk1jwfGSRMrcpBR0GkFFMyfQuhA
HiAISImBxe85o874pEZPtLAQTsXSesUVhSrUvgYGZ/CbkL38L840gQfJt0hyY39Mb4F6dKoX1FLq
aRStfNvmhZWDC5CU0hFrk5mH4gZA079PyNV5LhwxQ0HY7mHK6iCA0curxozWw6AV9dt6gU/Ktkol
prjT+kDmjTR5s6gWw4AqUuMo2Im793Fp9h4rmUXwirD0EVI4R7HwM6Poc0e6+ebHSgbKZ8X4qSQi
qpfakF4zDHBjLI4o/exnJqi8tHMTnVNkphn4s2PzgmiV/Qc9wnSWMtQGPRFDeurITQGokF85ZaMd
4MAzfSetb7912fJOaDJCtSYgmzDJxF9UbrqbxaKGdSnKmTqJePiGG4opKTp33URH8r8vZGv4W0j+
i7aN1roeROaPPNqmVa8v/8AtUf5+Ew8UwS7+IE7YcEszxZYSh8c5nulT5qnDdckKACe8k0/plAgi
bj4KITqkBqZKYD6v/j6P6sqz/pftGuN99agh4FB+a8PqN+rAUeb7NEY03s/9eYhg3G2a4lfmyLyw
6wHhb9ld33qjkhY5LaYpNaZBMrLPqvJx/R0qqPAnUXOncX1kFnAH2eCz0gSyI6wwXLnE2T+WtnJM
4RVrLJtTYQP/p3UvdjTkzR1aTbVnAqPCvMxb9yeQkO3bjYbi0A9t5aZmUkMdWqj8XK3o/9lcL32k
57J7MzqlsUXhlVVbGUrSydd+Np6IAWJXJWnyEN1MzXGwaVu4E8pia+d3Zai8zc+9hbUQwxsVTYef
fPQsQQ2xiTZPHSBkyRYXMaR2d7fghTpSgSkNEqhfgunB72l00gwDUxjDqWNCOpInR8rXqk7d7/Jo
D0Mp/yQZzIsLboTMK/dHwcNDdGbSMzOkSvZsVFHmquqs6FeK4n9uZSDa/XSHB0mnzgdsHR4mV9jk
PwB87tgQ+J6MkiRDcG5b+akFIxc26/OzJtZyro9uZs2BwJgVr4G5jpybUyeQxHuGr2DFlEUjASde
lcHaPP9E3ubSrBhapnM8SgwWV+ruRHYv40ekYiYx/dEG536u5nhnPLIuG6YmM1WWSVuv7o/BtyKD
ZzhlEn0w4d4WnF1+7SXXr2nU3PM9tIl9NZ7T7MyIvWAIUKOli0/nTiiCv88sROaPGVf6JhmiNTsp
5UGju4HBm+42kh3UE/HN22J1PO9iwjq79ebyt0QUdXUZclEjYcXONOyIxcKsnyZ3Rb/rBzxtu8AU
9JV8KgjWm4xEo1/JCGY1u74/jYujry1h8QwmW9WWGiznGljkDJdGAA+FqEhro2HNJ0U2o/LUHzXW
LHjO0jHkHrwlrWMR9gm4gtrrnixai5wsvtdjKUQjG6CxKkiRlFYslF4qD1Lmsf8qg7ZNKchQBuoL
JITmvkNlyYI/RGTarlGkCuuR+DUuPf/bx95EnzkwDLF4PDk644qw/m/UGfVDoENeOZMIhLbLHJsj
kAr+47ST5W6y1ISKnhvArrQ+DN5ErhGvXQbjBGG2czxk/GY8YAWYXSdwqCzQY5YCHcqsBDgGg1Js
bo4oBDoy992BbuSEwMmgIijmSk2imj++3XHcp+eL70TIorCE81M/lB95JNc1iFvdtDjgQ35AF7ey
QunK2Ge4+ZrrxEMaiaHqBbvGtaFF0+FDzRtNKd9ksfzlmqH3ke8EiRO8hSabjkzu3oOqzkbfsuQX
+PAcyz790iF2DhWCgQVtAsxJ61DrcR/OtwuP0Dw6GcHk3bE6GTm4Mkmp4CrhbsnaOeE91sIVKWP4
AbMpBALkAP3FDQ99p5UgQDbYq8LGaeSXH0SOV30/L7RV2rekDYdjWNxj3eggcNSuUs1TplQVn/zb
2Wte0a/3efDwsFS/dA10Llu9Ftsz6nCtW7yMXFBzBZ64lRe7hbzi5bZ95NJqJ+6WopVmzgH/sj/z
+V6seXMKxJ1aOpjY4XmgiY57j3Q3ekl8ZuUl2YWp7d3IBzkAStpTDPDxO60I52S1LV1A7KzbZPVN
OThw4+wc8MdHw+X6xwaBFEQDbSmc/rLetdDz+5fXjNpBXi4fph18piZ4op6ANecR7M9DPJIpt9XE
cEqspNB1PMjh9sOMyd3SS1rv2F3iRxo0B9g7dCTZklZ85Kjkcg7uIEGABxtHXk/F/Nmyrrkom4Rw
u7o++gdpkRblKj50ExZSHB2ab2sk1hshner/xTlvibd/MpwXp02/6O7dfJAzZx2pGCM4XptcfDV/
WygiHZ0D+FHB8UH49ubiDJIC/vGDdnaPZsf3Ewq3eGIyZSsdufYl4v5K60RfXAcREn0ag++iRw00
n7KQ1XNxZDNaussPyy2Prxh/0swNRlGY3/6UPLeAVIqCsH5rFW57U7ie1qt7OROjIAtSOC5/eE8A
qeNd2sTuVhrLKqFRx5vuPQnmHmye+NgwreQNmNUM63pLiX2tNwOkA2hOo7PlDm2z8aH+QT2C4ALT
fmGpJZiXrvNG0aNgDt4OUh6oLuHkgJ6pJ5qU0fqDvutgZJJE9I3SVNYJPcP9PGanUL6JJuPxkxl1
0125Nl4ZEH+5HsA8mdgYqKOj/1r6vzw1gAOFhXa3WzZvfWgSRmMnrkgy8i0hLh2UzhR4a9+XdgOj
b6b9vjfPV3ekxgi7+qscSaC/wQQ57flNUWb/5vdFs1+2hiVMLocL4DXvuf7scqsenyEdrItrHr7H
Oa+cF6UGgjxNoobu2v2VwtSp4RY7KwlQnw6ODe9Z6+ges+QBL9zUdVTMXhdlOHcd7Ajtg/HM3CBi
e581WATHc9FoOvv5dzNfxFCs4p1EW5aqfD/2oq8EIiSf0xwIwtDGfmkUsl8ByH/9K7VoxCiTh3py
/OJjKbbZMR0AjEBiFPNrkpvVj0Hy2tJ9UZiLhMJ2afX8Lq0f38gQ07HHmqY1x1RJHAbarcjSKPB7
0kAGG2CfwU+6krZ3c4UXTUfUxDOh4UCTN8Jugv2VnNnRVPf6uay7qD8flHlfcUwSVtNo5GW3GpU1
ioiA9hBbIxQe8GWPoCzOoFwCQhhaSk6WMtwW6YbA6eSxLUdnUbhVCONeweCBqjH2CqAFTO/hgPba
ZHj+29zlZcRMv+nK8hDLuLVYjipkRAl9rMk6mi7t74SCG2kdzxJdmUK9OonzBNoUb6UrGgoCRQ6G
TbG+YNwHIpsglDS1XT3ow283LNMFPlBJSEseednXbLsLrykb5wRrEtFijqu4VRY/0VKXE21NCGxV
rRRLdmoMbBgIbcU0N4D/hunndOhJvVtCnWzSDJ5AJT5HHlrBLt90kCCEFZ3O1NjxT23ug5hWjh5G
gcmI2r0JIKXp2lq9/HD9KjhwetHFLFDuyOlvUXIr7G+sfVSIGFAw8ow7r5p5t61B+4QUhtMXV4+/
4M5fp5H4iUMmH8U4B6vofcgOtGtQ9t86M/LyHItCL0d/bAqC2/kiKCegHsmSHgOcqS1aKemVllb/
AF4NREeh3G/psW8vZbEMhA5w/cgRXrnx22Detf1lPiELFdKhXPsEMYr4c0pjmYgzaJrXPJPEfaod
105q+JGJ6592NTgdaMlpEW2HeNMH5igRUNKWuEhD4pDiPoxtjYYvBbg3b/eDN+0nhKFLCI/O1M/M
fGMF4x5N+Fay/MyJNm6G/kl/m06Lw11jEoiS3uMsDR2F5P4APZw5O+HAQP4NoLl/nlF1LwoMSujG
JCWcS3S0omzME/lwR9VuUFy2Vhz5K/yQC4pmU7GuEpzdsvcaxJoZ47cHE4laTg2TIhMBASbFdJDb
a1Zhx+XNF18o6aJkx35yq44bdsq69q2Ep6XLY9FelDD5JM87LMi5vjkS2H15By0rEGVwY71lMfU7
S+4IZO9Ke+d7++oDjTLGU1InaljghQ94t2WM4j36lRp6YTzC8SuZOiQb7C+J15Lu9D+fxThyMoWB
iEhGZMtbo3EeyaGkL2zKVA9lL3mvid0cRjZS5T30m3KH017S9jZe287qtpYmUGDJqVf6tAF/rylh
8UKjJe+HSTcsxhan6SL5torTG7xHnSgVKgGHE1kWvVifoumcSdcEwWR3PwJwgIh7tJGycpl5ZUJo
o/+2LbVdKru+BOAgciqdi89dWNEWCUFMOpI7GGT54gJO36bJBiQ/3JIWcB+8nzXvwX6qIw3Pw56a
sQYHVxco73vaH4oSM8JEsmza6JokZ6rMrklQDLJyOmnypFLZ9HSLTopNYAMCq0pgtx23H48SFXDm
LaAdA4Yf0DFIe/Up1GmZAEFZwSWlBRNa5wJ35cLxNf2t+WcpWYpMAESXR0QL8DVshVB1c3b6rCAC
Srf1YxTG3iA4BLLrYn2T+9+2g8Hx8v67p9UWVvwJjiXI9FOjMGCjRXctMdX9xse2BWK6lYOIEFxC
WQRDItI6mjNDxcySdx2lJ0DlfX3zQEbngjJMMAwgovB+dvj+62+Gx2ZsmS1HiuyTeI13J62bUKvA
HGyTGgDITpEbB8CD5tQZQt0NUBBcIJTTGzl6V74LabsEjGFDudXt0rI4HI0mszBN8ZVNYbOIXq8Z
N3twtUiMo4zxBv39vs0X3GN0W3TZBdufT5+LN5S0wYmnXxIhFnmhZ3NIazacVfa7aOb96eoiR3GH
aNXKcoyzpntqvkvuadGFq8UMqY1jYDKBJEUXfMDpk4VyQvGY1nEAe6KEaG3qH22REO3bx50Fs2IX
ts52KJryt51bYgrvyTwv9+BE1Ix5PzHdw9c4GWMnu8puOoQHDGtrUtQe5IdwaPSDvL/Cdh246qdh
hpqEfo+kPFL/+kHTNig1LWXx+UC/qwz9R+lTEYqi2h/4v6CiqabJNjv3cJ45deCEAPBJurohHfO0
0mToDVls75Q229b1IQQu8uuED9NX1K5t59FTD4mCsCeTfA1cxv7ejlcq4tAXuSdYse/S5X+OedL0
zO15rMK0CGV0pktsoq/U3bFU4DGhYITlElVUk0PxGuTXpyMVZJ7uZy1zGYzmkJ2polihEvw0NlTP
xJKZOsnu5EBrMZhOE7GV7kGGxwa+HuT/wT5NMo4LHcNWRSpM139z7cWi+B3rQd9SmBs3GDZpXfMZ
EJrV5AYp1yCqI8fDcHMZ0/aR+af2mw1oKvyCP9cdMoa7s5j7QY3nD7ByFrMYagJMgO2WXdyaDaNk
wY0KvTlTo6BZsOQvg+uLbq4V/d+Uo3ezFOXQ67XF8DDu0F3tV1wHmQ+c4XYZxec57gsccJQl154a
6fd9xv/EFx9kU//C/KtuY79yo2qMVyKOd8Ym6FNOA6ko/9OZRdZzwfHVkx5frfBtbnyjn+ErUuH9
8uCDNqCLm7/ujHwKk3H1ujegjYTzNZPggQDlDkowTVXeyCCgBRmOkkGfaMyWSiLlkpdHmQAzl55p
fpkZL5As/uVwEyoYbDJ80mH6fa+lkHxkewbYeeB3hhawI5yYpnSs3jIMHOM79TRRJkc6fCf/oUDP
dd3sHXHf2pxSI4S5BgiYMOKaAI4L62bxM3frO1gosiZNsXxcP/Xnt2Kz8c7rr9RvlQ5dsKRlIYsW
XVrw+6I8Ihc2r0FNV1GKCfK++opet+i54c2FICQvihYWZl2oVGTN08Pkn7RWyY1o3p4UNCpl5v9H
gli2cdtEEry+WT221pRmSnftuM+eEVV+m+SU8C1NY0yGc+s8I14+f6VkJ6eGAvTEJGibrizWlkH+
+gK13c7Y8eVI9cMz2eQbcTyq0Tykeb3nOMhH5YEsAAJYVxYrN5NPmTK17aIKSb/7X8rZ9Hyb+DKZ
9r/4t9jWnuo5kVsZpPc5f3dz+bNDHJBmBV96FaSeI5RmCCcWSWuYN9h7AMbizida3Qhs5lGmXZFI
PvXPIeyn8e5BDI9lKLl8cA8nd3P1BVGNUV8aIdKBiv+fRBOYfcPrPZVprY7W7H7x/drRyyc6oJ0B
TyrMNrEcluFyRNm+gyzPX5w8dcXJBJ9TK0fELX8WEA1ZHDc0xbAkfeD051nvk4kT8KAp8r4jGpvL
mOk8dQTypt90vXPFoS3nrpdmhQ5EbdFEIa6shW/r5p+mcRoKEZhbZdA5CZjybmAEsAZh/8OtTGGT
UuARrECaFmWvZpmJW5+zCL6IOuu49CB104BzZ4bcsUAvLKdaKHuc8KtHEWgk938hH2WYesJHrxoc
FEl6PICxkMDBia9n01wrzHxgpSI5tzepvKbGfP4dXJ37DAhfk3PyXU06ejc8VLrOsDh8o2DtNYCM
Ef8WJr2E3WhaR+cJllwFDPetBSx5rP8nD5rd+2QJgbYB4CMFQOG4wogVjhJhlfndRDwLqpZ4insD
gMih6GxM7Sx7S26lb+8C/Hblm3jdKMeI0aPFsOgyOoozlcFAxVDciODTZ9H+JTSq3isnmm9/Y2CN
12xDaY7HRJj+01a+zeE88pKkk8rd5SK7cvpZNWe097LLJS9/yVC3gUsBsG5lOZGEtUW+KDJZJ2L4
D52eRndE5NvO7vmA2o8OJVtXe/+ud/HzErYmJ4/e43AyCFj9EO+G6m6UbZzdE7Yl0t6T+eNk77cP
mnmvjDAkAYlQCm8kdvPsSNB1uYUPNPaH+TJasdm8vdsYJuX2Q+/aCOeduAoWIlv+uh+kWcP0fLO3
TOO0XwVTfEIOQijXuvvmGlDHCuzE4q0ZrDZ6EjBMhv1IeOuSfx4fJP5BneiGH8povy9WcQGca8OG
w1O7cRCqEHQzKuYMRio9rjg6NpvLhCRfGYnwZgbhaKGBo0mOH6phBCUWGNS4evqMEUwojgAJPRfb
qXW/DbXgq43xAZWiemsBU6Q9T38I6nLV5SbWw80KFHy2kmbpdOBJy85y/dNA94NpLqPhNAlZdZZv
GiLBnbZp6hNzw3He/weUEZxGCL1p+t6AKgt8oKSkVEMyaR0deCEfD4uCb2SGiehy79Q1wESTpcIY
pDo5uhowukCnCMpyVnWUxY99hKJPKKKTj2ZuDssb+7lzCQkVzvq0/psKLBQYidqORpir9RdEpIVx
N+04uHjFP64k3vlPcOACNiILTDBO/WtXqOZYMsbCtFYxr4Ig2M7pw7ixZWiSzsmLjZqX11H5FMqD
n75CNuoN14qRP6pKNZgqcVT6q8lCDVYNPX9+a00hbqMx0rts54dD7DaR3JRiOuQw02Vs8yn0+XXz
r5cKlwwjfQisk/XxNWScD7ObpsPTs50PEO+7kEqOXKkqFUH2qWk0+sU4LvzNxdHw27F7Jt1NrylH
KK99sAdNTVHzeOdEPduz0GQOWuo46+xRHrj2qwF8u0p57sFCmGkPKrzGU/GampqxQ+rKtjEHWwDV
TL7zkMtZzQwL7BenCExvhecC7ATEOPF4XfLP2KjRlsMIvo91jrF2fkn1OxTYqqi+g8lwF4euS/hP
J1bYIGmRYPANKsb3/bSKxfgHKOb5lbCFemEKqfgjlDsurousb4IcMkQ+/q9/imcn4ysHqJQpcJS6
J69ATIPhKZa+GD+otFazK59v3lLLCZAT/Z/pVPWgwLxlcRLd7rZIwNoJrmEH6iirMRHZIwYDKcII
FulBtpO/5/aet/ZtlXuNQ8qK6Wf0SA14frNlxIywRvUSc8btZEzcnVMSTw6cAySS7VtEzQhoe4Xa
AZB2yC0KA8O+2GuTt3u0oVVnCnPyzbw/v1qAnfYd6pGvc1yopdrLWjVgTZnmqmHzTJ3XQLI1Qn87
Nik44BIh4UNR639cW0dPK2Py89qLqCQVZFL2Ubuhkh9EK/n8QP7zwfFUs+3laZuEm95CU0FQyWrJ
Ei+Az2Tfgt/6iWbNQcJEWYAIJj73PqhnTc9Jxe2UhII63lyibkGib0lnh93NQaByxqxr55y0NQGw
WgVeEjaDedyTn/pQsLeGbKogazgepAL9YhZsCkR1QSsi9GEylXtdSCVes8Me/7aoJ05Ct56P7P06
yiVEEQAX9L148nzfb5G/lznEH+sPHx636+//WYi6iBuNHzHnqNGY0oQ3lRH+STaCMc9BoK9nw0jB
suvSt0PTKWmFC8lhGvOyM/HgeKelxN7oj10dODrySpOcjPVXmHsh+GbKTJiftQFl+zMUG8Uy4TWA
Mh0frjm/80/nuX96+5GKehBBdpDsDQGQTvq8XRQWUxb/DHH562YIKQxwl6tSf51XoRq0BZkiEpVg
60GFSB6CBGt96G7u9V7xDdesVmpM+bK+WUNXKg2mAjxm0anvjmeZnbJd6nlTNUKGnk6XEnbIBtbU
lan4JlgWLBb9l0iTFJduHVTu/Chks06jp0ad8ZU7eGusxiJejr6YLcBXCXHQPg4o52Lm20ToIlJg
0TYHb7BHyDmOEFmTtbAoXo/eg7YqaGt2TgkcD/imZHtmVsEH48r4abwjw70kHSzUPZSWAycg+3EX
17GXbMTSt0s4WPF0pp+LZ1aNkKGVl6RLy1g1AV9oz8LNE63ubJtqkFPdKhhVFv3a8e7BVJUHszB1
Le27gQZMdjx4T2nXxDhIy5rcMPmW4/kJTAIHbrcEHGzCW0KW/3cmYd8vNPnN4Y5acp+/UJx+RH43
wekqVBJV0ctYUD5hMWza2QU9eRQdokIhYU9U69Bka6JzH9+8+2sAcGk5jcSj0ObGOJQ8u0otkWMe
dZo/yLKNY/C1QD2tyhF7pqSHMsBqmL/MkF7QPDs9XQde58VLzerWeN94vHS3s8iFDa8V/A//UjZ4
HUCLPg6ZeuHeDJU3ccLCtH+/kdXlESO/ohWgy5MkSnp0usAiqeChAy/p6N5zAgj2hDtk/VJ32NrW
FHbL06ZeU6g5bbG+xbq5B39mhzJ+CSeXwPOhb65bd8sXZM1QNwhYMU/OkpUVMVU7UBbn10057rnK
hMhs9ud0XwwG/assTtRlSzdrZCmHj0WvmmjbDjZEsEN01HykFN6a6Av6p2QC8jbDYr1wmpnQlmxn
h+enVQxehZ42eDhKYEatHWQMiNsRrPAkHqhRyC76sB9DDIhRb+xbIIaJ0gt5/yoQO1yyxXvvkcmO
DDsAqVQR+z9T6tUT4Qz2nhCijlyvSgRjFqJdFCniMPKEsQzz/DgHU/XVOf0QGawe67XuYqOLefvK
SYvDdmZQC5DC4jgO4wmPV7jAYwM6JbYO/0LxObscEbBpnXYNde8OxR1bFRgLtGV1M7CUX5PfAI8l
B27z5MraAfhLxm832YRQErON/aOhFwlVXgmbO7MYou9csjtZPTCDlJ3Onpgd8GU2tBfOsK3OD3Nm
K/SGHqQ8TEG3gfCxeUSgQ8Qgp1eWR6pVlDJmWiD9IW9OfuPfoy+WzTUReEri0QLrMt0HwSgUS9n+
Mj2H7WmjR+ew5e8LZomtnQmv6TnZSb9Li8eq5P3tKtS8NNoO0YUMAfVY0JqEjtFH/UwIf0Anm4hW
bxUvu2Ynvx/bc9eRHt6YmmVm6emB3h4kujUDi/O0QQSuPtlbi+2fY7pogXg0jFCEME6GtqDUV1dr
TXTdIQRa6Jnc4Al6sylrd6iSHvL2tWCTq8pdlOiS8axz/6WsfmkVHSqxnVB7zHx62SKH64xAWDFT
uaeye4y/fQkSXR5UD+eV/vGajuZxiu9gg2oWbr9F6wqxQd24iIEBAOj96G0jMBldIwekZKDJkWQ9
GTgQepfjNyI4+e+u47i8U7txcs1WfzqwY76+BA7T5VnFX+1bsOkKiw9TvEVNgMjz3nUPWLAUsyQ+
/f8DRD6z1jmMemFAhtZrGJ0gAlB7p8b+64DhfVywDFC9cxDEaAJsnA2ppk9No9ep7cxVZfvRyEXf
g6ziBDnFydXa+YUkTWAq7gDdXqzGYlUOqj4DkegORI6Y/Io8kF/9DBObGoBxtRAa7sqp9Erz0MuS
hD1TWH92iIe3bWekp1srxHN5YK9eRx1Q1JpPPv5jSfExwE+8iPlE/kfNmxo0yEYgsViX6/aRbxwP
lyBj3YkVw1xkIY2lwFxP+Bwtb2Ko/RwArNFyhXkAJE+j7kgeE6mvdqoeda13knVs3fmJQqv3AzJL
fd6+2JdCcJjR6Nvv2iJZjntDOf0Z1wmiDeYCWQqvOIn9P0zaHuvQcXH4d7RTJ1gu6uEuZTJza2C0
Spm76lLLP1RcMyrgXENTWAms/jsX+sG3d+qxPRdtPEoDWZgs4mlkZX2aCPrKuFbVx78/KXF7j5Qk
MNpyilUDSsDJ/AsZshR1GP4lH9Pbf4e0R1t1fsOseiqykgH396nAdcmKrDuNjsGgHEF5IQasVrP1
57/xNdEOw3+BmDrgC7mong8ad6Uy4MZD/DuFyXBHV8ZWaERwytz2inP36+wQDKd6nREumfCwa0Nn
3DgZD2XVxTMdlrBKj8jpbkf6OP809DxViVILL5Aoju4CEg5M8lLnIrfjbIBG4uD/+taTOJ3f2HbC
G3rozhkIp4pbKWjuDSUaNEFDGj6PZE4hcMu3LSeSQj9e0nqO689j6AiGden+5SdzwQ34zRbrPRgH
go5lpIH8kX5189/ErZ4ZdE/mKngl8ksFYVpB9AzTEC83qoMh0ZRUZOz0tBVFb4OvPddj5N0+7Oz2
uiXMuzlMg/sm6YhhV1bXeAGHkohS3i3ywbqafA7QZH2RdJnF8K/kqBHadR+KdOpGWanhE5ySkRN9
mv0QoYe/h2oxvmUZSjH0YJvDyV0RrWX/6o1STyJ/LTmXInv8tDKR1tPS7Bo3Dzc0OW6RMmYBTsnZ
9ncmfyMLP8MPz9hUn6hEDKaYRDw4IYETMjx9C0sTb0+rk+4g0vz/0l5Gc6u2yCjF3IFFinAPlZ4z
rULQTv4YaLbVj6QT1P9+DOMft1GjE8IBtOposSl2L3fr+PI05aU595Hk17iTf9PI0C8tcCXLdFZH
dJQl8jVhz8ZVI8M7T/vhZgoSoj79+Cd+PQTpSEPXdA5BZGjHcChQiFDh1C/m7oJPN8Y+fjfzvY72
S8vUUJXAUtlyfVlWVF6Cc9Xf5tIOqTLX9/nyvdZnpglUF4LIsjrXKq1xiufUoAW8xunBgZ8nngKZ
KK9/kNCY65Nh70CfxEmtWoiVDtzpLGYmbgEmaDiw9SSlvnZLSwXVTg6cieF76MmoyL9J7ii47q1n
UtHmG47psO2o4g4uClekgPtFltBTAOR/Yfx+U6i1tHxiPvl8ggszTnn8ImByJoUEsm7gt9hvd8Xx
jBl7K95zxEXz2PL+1a+GrPXysp5H8I1a8aen0ITf1ay0ZrTewCZr+wM2/nvkTbgivZsZHllLKKcK
jWyKOwuT1r7ernpJqK4aG+b2rNHAKY8flyz6cLN4noOSg4MPvEiUswSPPUPQkms8GhCvEXMDmhud
TpBp6AjCN4sP63UjPOwp+Rd8gvwf3WDkq8SDIIRQ4nyi/pUPFPxxJcAg/VNZ2eiU/Lz1w/lhLMTe
TTW+Nkq5NY8xTmivmY+xH74q1BbL8iD2RoXDHfVDn2nZQpIB/6xm6lPOsAdkSSvXc5cRcw39xK9Q
AnKcMbejBpbmbT0k3MUlbGYQA+o18Bzjw5Io32unU+MOx21jr8PSRJoIrFPu5jq3zQMgJQyaEctm
MzmKDra2y2WOfVSoF7mW2bEuUw2Gbvv52hK1B6DQ+5JEWXsMf7QuvSjLkdAECqOe3R1rlvzM75+1
z2m4R/W/PUNKwxREseh/X133xzZ01hxKl7AcbrVTYSWvAo3nGnYLLgIbUqvEVc+i+HyWG6HkHZg5
9KaSMdeIlcGnD1mEVOohUuAV97ZEu5PY5f2jZ7R6QrTV5Dc/s68xBInMpp8uV/eCfiqgJHOxXpMp
EZBtpQ3xeurg6B9EIrAZNLVcMhBBdU+Gb0uZEgwnQ6ykTOZLv0BZVNZSpzR946eF3xHIJs7r2SKB
AnEBIDzGv6hS1wPLvbYmKvjXmDmfayy8pnnN9ygeVuQ+U9IT7SgQGYNY56K9F5XzU+DoX3Rt54/C
LWKQUZFz7LVcs2jlKf5Q0wW5isK4i5jK3snrhgX8z2+lB/NVl3hiOn9rKX6mtMJhbrXu+gyQOqq6
dg6iNW0Vewjh+0UpVlenfqxLtqeFHSWwaWFaK2LmPB5vXeMZH/sAgI+mrgr1hXqBcfOoeoVXLMCw
1WUtb2wD2GzQSz/vlJdYaNvPD+TQWl5cc7EAba4bGBtSetY/RE+cfe+MLl4uj1x0iM0nj21ewfs4
iWd5GFS58lgpHADYh2QiNhqwgr2F3UxO6W6jN2n2I4iEAgNGruuSEsdNW6cFxQBAm/rYI02MiMBg
DtOY/hBGWjhOHR01uqEiwCf4aCTeq5UdThuXlBHa6jU/hqkng1iJP4fBTHSq02urE/rTzYuuEB2w
T/e83y6l2lXbNHlCKVO2fMQwsqMeiIr5L27cqEt6DTk9jFtempXjf/Kj5cBxuNaYUZRGnD2PAsc5
PYfUsNDpxi/8FqO3+2pidEOV+cX506IcBItcBedVTysBjkymqyWZxiCZGlHFoHvXyy0Fi6ilmj00
mtldnWFI93QnrRC6Q8fOvwpADYHy38azAvI5WPf/97YmfDvgSyYiv6bGGzYrBMxk16GgjDBKscz7
4Z2F0z9mknEFk/nJIgwzlkBcAwU+oOlu/GNq9oGRte2hf0u2P4kvVNBJg8VMNMJ29TaOvWaUKOZO
6FVSdYTJNqcN1supLh6Cs/0rednJxtQ0ojT3Co+f1Ng9Y2QIPzfAPcRWnLZhA90Hvzld+bXuazlw
4ipPENlscRsWLdtyYKKszZLWcN6RME5+/5hRHhOw5b39Ge2DZqzrUVs7fx5GyXAmicnH6DYp9HHJ
NnoUDB3l7AxEz5+sRCwQRecQkEwackQfF5ljzeyuFXLNsTakvzxp/RLFWaHKNW4vmLqod7MzHndQ
t9j9F0Dn0sXEPZefvg5JBzFKfkF025OErGH2we31VRhnpFtvW/TpM+4ovD8BpY8eqI0aj5nYpUST
kWbb9u5pbe9e2Wwm6LlPhwCVbtNQARrs/ywN1h2YW+CzOeWB7XgtkASEENRYpt7QBxidjs5rV8UQ
amMqQp3bx92TCR41SzvsFRAXQ17RaSvLGLT6JwAqBPW6L3lwmFU+d9W/i8SoCfNb5xflwP4Eyq3P
6ou7xK4v/k4HW51YG7xipwmQoAzHOLkPbhVXce9ShPFnVEm+7vZsfMSSWI94RrxcFMh0qkLN0oc9
qM1Ja/t0X2Vcr3vrOFCtn5yPm3tqwp01Jsl+SrM8TLr5hVxTW69eVw20D3YGmsHCBa42CNhJd9Xc
SJsbJzid/NkYGA9ZCxWh3pUfopHIkPeIaqfHU7HhkQsS6vFRG9OsFhUarWI5ySiDBLR7wMAk0oRa
E6TYIfTHqFhSN08zStAuibJXhy3rtpyEcHGX755/H7pqH/zn8B3YZNkkXtancQiaLAxFG+v5d/AX
X8dJ/TKQfzRPESaFUxOy59+lhkVguRhGJFajOkk7/RxUy5FKJkPV4ONKRW9U48g3vpsZTiLRrHIG
avvJa/0/puF7Xc3ZwJFbB79YRxP64btP0IkoN2Y2K7DIrWnb3G4t95unKi4kkS3Jk6A/ZYP+YVp9
oNiDZEVTxAw8G+DRf0ofM7KhZiCVo5O5jzBSnzVoysI9Cg/UxnUd41YxGAE7sf/KdMtHTkFASnyC
mrw5DjclOwYy8F9lhBPgUWLCDqmc/k/Xy/Mt3ZTkq8FqK2At4ijE0s/Mj8EVolLrzrtJxlws14gn
P4YAMZTch/sL9yyTtZr84aJfjyWjw8h5Fq5ai/1M7qxRdQdWlprI6PWTGCz16PwKP3S7fBuifz+Q
ckwcPl5d99749904HQml1P8ho3u258Ox+DCBL67Ozjy9NUAa+AZdsTyQXKc+ZZz9YFD1DeV4yu9J
q1Cy7+akOl0NbfO8wwK9HTdUdgedUWOtllPxdx8xveGYx0xzVRe/X9cTfC7eJuH1Oy/PbXzfUxAj
nfbPtFaiorlfKxiAEv0B8Pfco2bANJo4WZO0w/Aaq28cLt5Gu0/kQOIn840tSuxlMCKLc/gEMl4w
tQTTF6zvqTegSpN+1B6s6nG9le15zJW42WDld4oHiVKsN5GxXqdbUdagVfXnkSM+xvhdzIAQlmAL
ECxcvDSe+Oe9s44cKYVnSwn06Y/wTCdFONdrGdJjPPWl3FUvZEHuvjNsJ8B+5g161j2FSeUAHBJj
WVxq5K1lOJlqja5LozheXvv0mI54n6fOFm/Ah3OPAX44+Wa4cIN4aQ02DpZxoz2x4wY2WGaObddn
1DxLSqHENj+GpKTg7dBJ1uvkonGSRy08JP2+uXp3zXGLVw8S83TkbcSvsGFGJyxvWohVApR3/wVZ
NyypkkcZKY4djQhDyljdBCoGv6Rj526IHQuvviqOUoEU+xbMUOfeL6wg6Hboq4aB5Emood8NeJ5o
omYxbyqTehyBhz//NrI3aZRRAmP1AGCp0ZFHKvMCLWl3I4+Ua3KcsKZGdUbjBAELE7DzMenEFozG
731Iyj7SJNChRRnXTASE7Fdw08xjO6sF5bKE+bsGukt3CcY6vjKcrx7gOZnvfMcTvokJiXBTfui8
GNMfOtntFiF/gkTe0r7KUcUlUKcXlHb17zUS5prEsxEUTqs7HcV3UrRIWAwl+O36VqHUsIAB3Erz
8tkDuG5FC2dtEtbEy4Pbijui3pGKEEv/5gEd5EIQ5+EjedShFatP/346KVRB/Fs21vbqtggRHKya
IAxvKrOr8WfW332gAe2VzCvnnQRUHVdLBkO9thZJlep9FVA32ho+F7C4bhqzGdSQ7VCU6d/Rnbb8
uStBILqnuiMvhEr/5emkDiplLS1zktY+MM5vXhbagBrF3WDqc7/JOZfUcchYr13MJQMz2WW3Q8ge
M7jsApERy0uVVZbhW7b3DTDl9Y5gDg2kMcCdTUzvbOLUp5TrOJSDrrXhkDTrCto6BMNvKBAo1r2t
liCp/mL41OnP4EV6Emr/0X3G7k4vPkASaLvGZOOgXvZXa9ObzOi7eIIaRSRCkCzHGqKBdroyxAcf
r6rAcIc2SbhBDSrcynk0dBD1R6sYYin3zp4CK/OlcgWNiLX1qoJvTOc2fhRSu6lTrVBLzjsPtVP3
Ezej35v+PzvNEfoEbZGRX41cgY+qaR5tfe53c/6I0Bzf+6bh3Tp6NVsHiICY3go5g3kX1+M7RlhS
A0VXyS/Zq9vlY8qOA1lnMT+nx0r67H6kXf66MemX6lBIAi05um7XTBTvHiG1XtcfHs9QSH8Efozn
WmPQe0pt2Cp1ZxSeLT2wFl+uIlVw18YHp//CZZhZJoEbYvZS/tIBhG5yYOwtNyy5n3xwYbScQfaN
cyUPxmV3K2aoXN4zPAUep8uV+hEpbm/mPJmKZQ8Ne8WSve4Bdh6IiJ7cUMA+MY3dI/gSbj38nFUI
7ObEr3KmXLlhx+Hg+5IOLpmj8B/Qb6Ki/5inpOT+6L+HDTy+/aif/GKBkbjCxEdgjdqYxpu5HvU3
Fog1qKup3t0HhCSRce82gTAuEIOO7CiOsLY7eQ2TIoAhiY8jDK3q/OVEAD1ECkUJ68Sh4E9brLgi
OtmPeHNY65Woi2bFO3JrkR+q58o+qTuqR+yKiMsuvT/sEMN1osqPVuFvf3FL9GiIkwU1WjwGfv+C
p/gVbppvGxNsb4ZsRAXYTDgy+FVW05QI6NZUsclMCkpT4et/tY4TMfLyAIepEo65l1EHMkNB922i
nJH9IdQJcLkylm2L5omslOpoO39ra3vBQ4wdvmrlNTJcf3Bm+19TuGuNueCfo1lBJ/rFX4YOV1oq
Y1hrySYhMCD229E2GVE3GE5ChUYVtmpipqAvBKaLZI2Oz3KqBAP+QuXfFOuDKuUiRdaEsXd53N4d
WaBO/DSH/LoyRt4FWuJEKgJ9P3T8Xq5xlNwB62qvGC026saL7RbyFpMvadgW1q32/yoyejfQ8qmy
CfZmGGg1rFNS7wZxt06vROyg/m3LnBQLz1bjlhJDwfUh1ExWxsLrBpJg+YRX6nH06V2rNNRtDYSH
JVBqVlXEHAVINdj1dmZ8Rh+239B0IqYGN+rI9ybzc3IQyAVjs+qUd65LIKkenXqOc2O/HIo7mT2N
FuTgWCr8KNMACB/1FPjJhgl7oqy5cyVf11VhOrLiZS8D2wYs8r+ieo21LBcwnzNUWU0DhBNyq+45
N3NUvN/2AM1mE/2fGOHjZQhNIqIthVc7A/5CqUqRhSEu5yCLfn02tb/1lGgSGhASyyGBrImBRC7z
Sq2qcsF+RtEzYtpKqmuroV2q7yc/ZOD/iwXjhrU2rXJMZ0PjjHhYVZWnROdlWq8pcrzhLQNDSGBL
79tABt4mf5WYDqzMHjcExWDFNGWERRAvT2eEFXDrWrFAHQf0ixzPW6LQnF6F4nxs3F6D+2nDnIo+
y/l3td30L0sL/eRKWEIipbVAS38Ax5i9/6JQPI7bHK8j/zCceiJv4fyOodgj+b4JlspaMy25m4Qb
/DDTM7NgLV1CcfdtCHk0gxm9nNKI8rmkamAjerkWabl/jxL4d1pcG6JY8/FDZK5UpRj1a+NHOH1R
TG131pgRojdzQ1qcIrUJFe2/Nq/25ys6wtrBkSMZlTqneSmYGew2pMJQHx5qMW89HJXvmaa/kNJi
TwgTPwu7epdtqt3VTI1uZSliBoxi7zmA1MPJhmV5636ttGCg0Nr59EzxF/TmwWGikeU5OSN9F4iI
LBeno+jVk3N4UR2ctk0Fz4Oay8ik/3fpEUFKvxsXS9LgzDnCXhoPA0jDzo8pLNEY3iRigunD0/hP
exp6V8ssNGKePcB/upNjwi8nqPt5SAZb6jmMJuKh7xIcdYZaMxuUcerCNf4h7MtMUqSGtZFmmot9
SKsmDAdVDeM4TR1dab8vwGyqE8bkkGDVMn91pqVbRILvrBDwebVR+AVtcWJ+Cxmu9MysvgI9KofP
OE4N/lT6xWZSaPGT6W33Q78G6C0rRW9hGXCUurj7qT3+vYVlp8tOELaGPr3lV2V9qc4jv9tVaGMC
d2FLb6+5TmOWX6VohYf6Hb7pVZFx+sSo6h/h1NUCppBIQ16GxEHLgFBOjeyUmpjhNqm3y8t6xnbL
RY1UsIFiTfen5K84rEH0+l5DA5DNtfsGSnrxu+tiPaEs2LEgwliesTApkTolYFo6/EMo06h5Ktz9
1dYDwa9A51Zvcav7eGFWDbfVdBeWEo1gwCGI2xrefZLNHJT+CSPw4gswwENCWGEaMNwsf+RPBx/k
9V4ETpjwYsXpmCvYsr42c2YpM9w9Qq9I5UjKj5ZowJl16Z2OGBWgn+nHAnO1vTQSYmnlAmk5s245
nX5wwsJEvJOVcignlL+EUvaUrc9/+D9WGlv372TpXlUBdp4jMB7WKQl2czlRl2d4MYVg1CUs7m23
R/gHQ0DV2vHW0Td3CzAiOcxW4AFqjsV5YRFLZfrkxhPgxmw8XIjqqFWqDAdMaOXPp7+VjadiBPIe
A5OyM0D5uYk481RmIN7vby9ZbSmqsm5QbcWlrg4z8oWD6QWULURXmHf7D9mSKSH0IUAgqrSUODYx
9Iu5sPpKOpwRisp2PZ8lQO9SYPwmKOq6fBymbJ8LNOBMu+EcwPNtUjWRsZ7iQATlRA47T6AO2MRg
Ba1iPUcI0Lp2U9zIjUPfNfLE8MD1I8c4gi7p8VwkynToHnn21qDa1fXFbxXjmZLR5g5TH1BGyBUa
X+1BBQwoqCYq1Vfl/ojJubcx4nH3wFCy9LybaZ2fJnhC8p448ygBSTZ/qVFFo3NbPDhOacbmV+Bt
Ag6qruzGuYuQ9+XbTuL7q7qjTi5HrCQUa7I+C+MbrNWZnsHMOw3ZTQ7rsKcAi0Ok/QF1Pn44mBEf
7059VmZvjD03T5/ArIu4OM1FvvP5+8z6IgXu4PEBTjOYRYibQ+oU13SoSnT1ZxHClyNiPz75bXBl
dSbx+C/e4qSgoV+avwzwjRNMuvKiwlTuQRgvIEPN1FC8BhDyXBp7ERhXyD7EM7BbNQPyx8ZmbdNX
MeGzPMmTYoZ9icuUaW/uhDvZXo+Nmz1kWZcz/ah1ooyHhYX1ZZeuRljS7RojLXdETH/OhSK53EUk
sSgl90c8tDkKh3tLpP4Tz64MGBfcwhibBllkzop7s9JX1KI2aZFYr/rqo23VF8tFHforQl41J7CO
miIe4IICw1bp3ldo/SiOA6trRsy9vIqwtu+KuMtqIcMellXTLlVYcJG8myxE/2/5bI6KouJ7H8Jo
XmFRoDaA1lvtQ/kXpxtCHhtEbolU+0fjDJHgbmcYYLr59hV9njt/q/ACmJQIkT5yCPM+lTfAJVa8
tNb/4tg66vEUAzkQRJ4e8jbr6cWuNYo5/j3OJqtVFz6Pzr4C6vkOTCCgBdpS/+VAUIkqbLQ3u9aN
kD3FmsetffWGLnuMIjjFw54+UASRQWnCThCdQ/LZZ0uVGZUJeqXcMcjp2qxgIuyfpxQPy4qbBxvE
Jq4kUtHDvNjSrm2xf776NPSAx6V7KbgD0vBSiRdl5JAurFDScqgtDrQbn1sZUPw89vF9cd6m238z
N/izVdnFuqQGg7XQywDt8xyLl+DbqK/2CAbnawhTwgHfudAa3DKIaWq/1TZmyYr+eHdc0ju3FWWR
3f8cras/atBj2xxhhByncLox9POrlAhv+okUBx0ZaKJ7wzZk1Tl+3WvEDY77DMsYBLZWwqFs6ju0
WJdfdz53mwFceM+pcRwXDqZKBrnkGqxPHcamz8+K/fgCZMeZX60jDtYozF7PAZUjBl4k5ngZ3C61
1nnKRYsNkFEiU+tsEjFmiAnBiNRGInkZtWYQppZ93hL7llS7DyF6v2vLMNHYRBd53c3Lq/g/yVTB
Qv5PDu5ums+ywLWZOedyTi/1PoQLKIj2O9Euos8/lo78i03zzbM8GW6jw1nxxb0p6fmMIjJlGJoa
gb7EOXPWMWJfCvRhbxuh/X215K/7SyaURISKt5I+v4cqGeIjZhb/WeBYKzB59og4W1NEdp6sC/oR
KIp79QP1neCXV1DFWhBa/Zu3J0+zYdKon2/Cfaokn9B2IdUAldLaXc9cg2QSb85Hoy5ABxpwS5nF
ff5xzE6mfErYrQeoI0+PbTkYylnwgHoQqi74VtiO7G0LYTBMoo4KthvdlC0X5T7OZCEHerbCKJ21
tNpjb4jjjorMDX38omtxxsY9M0KRS7ES6Wiz4zKuPXMwQyBLdn2RKj7RI2ouDoaAt7JRn4571VkE
ujQDOsuOORnnwToQZ0avmS/riTTwIuCVJ1tOCQhmZhJoY3TSN3IAoXiSXvdys4kJ2dNmq3PrJ18W
twmFP7AFUW93hXFu7p73dUT1LxfaxNYk/askT5oBZc5Ej6gyhe9j1HxY5GrDE5bIi3ddmaZiQTgu
87njtBiolfDnbXsJogtivNDdL61GZ3VBR7MFN1fnA8VJ64txcReCWBtHHVERwPdvVGQ4cL45GVTS
Q4esRKdhI/sLN8UPtaktn2lBuKdqBrCWgh2gZfMLxg9rp8hb5qqSt28TvUKkGBs7uq00JCE9Z5Ii
wryb+QMW2WQLRMwqZKmqC0a9p8Ykjc5UkYS3HNgqfCdnBELXrH5yhZ/owXRoJO2kPQETMJpRCz1k
u4Kll4qA61IfZ78flO/AmBYZpq31gqr+gFhKKorNHRBvelEZAhnqqzUGfzOWCAj37aM8w4hOZWXD
wi+bheIc7JyARnbrW8KVN8+CMf+/PvCnLIDjrrBWE/cX1jbqr+wFF0YGfCTDkI/SEoM7v8MhAElE
J+iromiqqBMhvad14Idx1oc58ZB0kmctHXHx3NBuZ1Ab4+iGz/7WPGe/a/GkedrDyKtYZkP7uxqq
jNmn16zJboF49C6QE7Y2bma1JAq9YbHa9OS7OuSDR5Z2bu+fGevWbG8JwNSCPeCI3/uqKngWcGBL
NVqQvtcj+R3GhwdQQ59BpIpQgTF7sIogrpdpUdl0p2+ebmjh5LZBZTUj/6Z+0KBgTW1kWOYm1snw
Lcpi3iqYQ8V5y9SBGNpol2uyWEoOifnZKBT9UEuOFchq0H0SlkyY7nVn3HMjYDIAY+hb/Pn+p4xJ
HPIZStp2pA1HzodyobsL+3nkImuGo4ir++7juMcbibruFAz0gvNyXkNoqUgrBH+EgKo0TY3U4YyS
TIdru/nEGBmRdTpMDeen8a/DYiV4rSp7u4SREgKMbwjy6VsTt0yFpyqPXKm0KAUYgDpcJkEU9Aol
A3sWtmBA1Hu4XB6tUm6g7urUoKa5WlDnkiy1dYIdMBU10n6nyQ/9HBMpmJRbu6kGdhBxUfX9tBFs
/SeeCXCAvnoWkVe63ZdvOWG3eBXZXA8bBH/qyuar0Ce8FdW+Dx5Zt9z95VJx2c97nf+90RZAV0Vr
o6N+4N71BvWk8BnNORjNulByCqavJQerdTrd2j5suN1u7XLRagbPKxhngeUBcZYfBMCcmdCIQKCc
p9/qPz8LetG5BRm0Wqly98rqyEZj3vgZvi13+8lRAJJJqdG5dbPwUGq1WHfYj/9eKi+Ihs+ZfEYA
7WmXpNuk4TIbhynRPZKqg+kwk3Or0gR6MbqyBDitt30ES+3WAJ1WanPqzsrvUFcuY30pcEIpQYZK
kSsjs+HaQf4S9iw42vylFgdHyrT7sGE3tZWw1iCV97kktWHDhUU+fA4pkNGCeDbxrI6cwSUlnZXa
j43J1Dng2LEMxdNl1On1V9I2ot6ON5cUWIOnO+3ZXvoIGS8lRxyCHS8Oa5Cz4lferfhxhucRg6y2
ZBglEhGIH9JUa33/SqTKWKDqOwtzAloMYBKKSfELhTJwU2XeOND3dZgSZbjRaZNBvLRLVAFE9T8W
QCV6ZUckSUsvF7x5pzqEEAHVbqKD2KsUUFpip4RJxC4ZfBy1SKITb06+A4e4jU88YI32ud2memAA
f8/3GvSQD5TwLEVhYMPKx3ksutvO46eG4VjHt1UMOgVBLjchWgbsPJPLJxMVYv+DYX9030X/XvMa
4BtXxunDt+lg253unqS19yOBuaiSq7qmakYjjjeJoRVC+QILOR24PUZaYb0ORttordzyvBTwxLpN
y8+hZGinxlO/VbssOjyGF+gQCghx9+qW4MQFrSmwMBwPOuygDoHhjpmFCBQa/HvjKTbZ1HQjW4wr
HpIEJDEtUp7xRHoYe9wjFe+G4ftU7LymQRJDiQifkUKOVo28u+SKB8UjmP69XjgyHyPDUyg2+wPd
Hp1W78080cZEILDjFTNY5aYb9HQB0wBwPuCMHTjxJ1NGTfXYWuqEB6eK09OpRfb9owlDEEGw20xE
M8WEqyWLOWieuIUSO4qpvabMMkL8ySbRy0U8DYcmWPuuhv5VKmKR7cvYcMyJn7lfpaYi6kCnIk8r
OP7oUrWQj7ADZSfY4Qdr/ABjfIb0kZ7SE4Lr/vWPS1NBml3RbK5O9DyEuiVet/DJKFFvn17QXV+O
iLiDAV+I2imyHD69uUb5nkAIrAauWIWiWFHtVGhfzODo2gx8egqNnL6QI30huEBQxbJgnXzQ88rT
0SfENWAmPIn7fyCa9xlLt6MnCfL+aBFKcv5GgTk2Lb95vY/uHWwUivBqi5ANo3f4KMrxZzq24h1r
j5OMEKL9WFIVI68XK7htvOnnxelQfNWk48TT19EDtd5kyFGWz5ETxCaJHR/aYQdWbi8OFZJ6FKRp
3iXQiqenziKIN4I1uMwo7/uZIDUvGXr9h4B4wcu0uMQyiucEPLFuwY7lSMkzXQPaGbl37sBryMf4
mNDqud4RL21hGGcIwlt6Ndfw3WaO6rP5MdUMhM7LgwQmtYVp7NBPz9gKt9okykVk9QiFFR76TlIc
xRNaLRaZZ4IqiHqPFHCvpOlDnK02/9i9VbUOuu2Nq+OvFcMd5ZcA53a/EJxD/zbfVXyXc5aZb+5g
wMZsHkChCrR+pj9Bw9xpuK8MfC2KE3UpJa/3r1jJgTJ0+7c1NiRj3taagExjAOj2jm6BPH4AEbqC
/FZ13EJkqdgZwTNv2TrjFzU/bbDq4d0cq+x2BnO+V5sCnRZlMhLVZ9rprOCNXHBhMQT5y68wzlvj
tfqXfBaJch4CqBA3T+WIE6Toy/87nmI3x2BgSGYJSFUM0yxKKBagWcIrU81BY4b+s5WeSUW38ULs
8bNnj12Sl9aR1/Z/x94Q3d9NUm3anyTZwvLhZsXiR39maLzGbnejtWeH9eUI7u6MJ2nReebvYnD+
D+X9E8c5nst7LU+KNPVCoOPGaDYkdlKnunNMj+M4LpH0/Yn0hRGyachEHj8orXFmgtsUyw8NlmEX
lRRCQgw6yTUJL6456/NJum+zMlUwgpVE6/53ecK6d5nC/MrHC/rNth+7MetSiBoTKV6bmPxxhf+e
XWhLUwWxGTzZUAFfoVCc7tglFHNxVrmgb8FgKzu5mKtiJzetLPMHukkWIftfDJGvkoKbEypNIbzZ
7O2XZJ617kQT/T0z4QsydbEDW1+FIAWemxeL6+0E8+bHpyoaD0XFhIWZ7gRHjgFy1+Oc7ezJGmR6
BgZ2tKnFIUojQocvP1tvFP3Yl2eThh9G9Ei+v7pkA6e0HpUQFfwLplYWvloKr8j+QqltOa6RbWuZ
p+NzSen7LVObYVYUoc318pjbM3z2Q8vB+5F9K7NFaES5209y9ANOW9vb1Zz7aPdfChH9CBkt7QZJ
9ZQ+MNKRHO3oyphEI18uLPZoXHg1vssNNXMzAjpYFiidSCQWEWwTG7m+ynkebt81hnzhJatSW3x5
ugPcs/PzjzAkWCXuZSZAUvyUDQRdLfQNXnkVBW24cTsF3xYBLjqpnyTjG187MI/MvyA9wpi83+Wv
r1lGkGP7ciwwvWl2/xSb/Xn3X8KlJDZXXCDMWZ8G2N+3UZU34kj7T6nhSvhMBoE54C31c1S9VpHU
jbEuSLD8iMylA7OtDSvGyoT+0UeqZSFOpmIDDqOZ85/wfFW2sKkFUheM28NGMpTiaJmzprGpg9VG
nFBiIC3pb076tr03sgLx0aX8oeW+zEwYXx7t2+YBBw8qeynevzojH97KjlSn9s/Zq8O7KfKNWRz1
XGdLRiitX5WlXi6MOnBBj4GkM1KP6QfHlraQhuVIo1kp6tVnP9pMljnKBieETcbb/3MDidch05eC
cb4bhbWtWF+322mZTyS98k+J22GWI2MI+K7bUQpf00TWJNsoG2PYR1MytneSIprNy5v63fZPUI3D
zvTbUsOPddAxlDXMSOMr+p2aysXLgRn/hCG2VF/OSf0whM8uqeTI4h/UvfPs0O1X/+7idcdXtYbn
jWubX/wKMh6e0NXups5tdO815t76/QrP6+6ZF4e5UtpTewcjRZe7I7H9vTKwlrUN04uIxQyPV25q
ZPZ7gNU0NoC64d/w+GqgqJb624V//hDI5i+bZ7zerBTAWQToEeMgtjw0di9dq87fEnq81/aili10
qaxOAvvqcaTp9jwDEqpLFrHlFAe0qZhIUmPkunw9CnV7BPOVnaT0WQiGcXDaK5jjJHg1h8pB5FST
2jFuPM8FGrsB/+Y2JgvY05uhM2Isaxtvyl0s26a3+prT1Xc4IMBvihNnvzS+gxqqezF4bhBChAaf
u3l47uzaQsTzBJgjc62rDYAq+v0crwJNj61VDOtojfT6eyhcTjKqi5ylH4vGW4Ooa/YiqYmokE34
k50FkJRx0iuhMkWVE/Uh6r8R3+ujRyHmdVkJdV7lIYG57pYaLdWW6KMUkO2fZNUUKsUSPjHFT0/4
bMynXbbBwQEr1lSuEZcXcJklct7S92nBEXwuncYwr4+DTthmFNDmAvPLJcu0lukrp2s1+m6lHyNB
Cvf3L68bNaCQYS3AVimuOvKWrNAhhjrej8KahvVN/syArqzp9S6U8bzqrgxQA3du9fbuFXggnvff
FtaA4CvDw9kfgqQUyDKip5z1EsPB8aE5BR9m/X+CNEDyXeMJCEsiVStBuP/eJtGCGvd47MqV8pQJ
i/9SgzTglYLKWiYsH64aRTQ1joL6yqh+TjYwvcAGbkDfTevC0niiHcxZRcYZ+PaFOa81Ah6taYrP
0c3Onu37UyaNDXQsMRxJ4TnoteGa8a+rJPz3SPXbCBu3cLXxsGzath9xPQqndogNLd5Z8DjovMm+
dfgxHbm0nSNxAhXC2RWGYLAcPiH8JwPPVST6WzPFjTWFuhlwSyi/5gH1Rquj0/8dbCSdd5Z6h4+J
Z41CdECJ1FrRUYfl9NYlr+vR38L+aeCu9Fgrdao8PxgPK33GyL4aDN8aqC/3oFuXvUbJu7wFewNd
EeMTKijOi7Lr41g+QW680n1/kdumljIFiF6CvsG+IzGFgSRn7DvezP5CypZ1Yb4rNTR+S+e1sLfW
uwg/qCkXrNis6w6+jm1JUW9JtqvPfdmpsz+fB1LyWUBJWABKYpfWWn5qN6xqsWIgYOoAmP7N8UAO
mHq9OvCs0HJZAghTxb7F8/2IiNk7PC0d26LY2CSHAm9ytVlR2DvOcdTpJcRfImN6raJ0aCD0AcBb
2xUmhl3pd4x2wtBf71TMO9DjP1KzFL+dMoJGV9BJJdnotcwU3HRLQV79G0B9bSNiFq/yKb9MfY1d
Ofhyyw5xU2TipW59oWDFuF1EsaAFWIe0ZsaMn57GtqMg/eIlD1hf5VDCKuVnKqXT4jMUT+fYxyOm
I6SKnxL7ki8pjD1MrFwqkB2MEnoZK2bKTR4w1jQWYKEKCrke0Ax4oN+onvTpuJIEA6YzJfcCTcFP
oU9NUvkY2Teee0O0ppkf3MYSx0LfbLhk7YmZ2cr3yWQfw8ffnr4sGAYfV+8xzG7mnSAeQm7BcHf1
v6VMtDrm+NH9p32DggoMMsZ2owutZ71QNGnwgU81EproQ+Eb3Tg2/NcRsp50RU1Hxot7HN1m/M7t
YWMB2ei974zLkRRPToi8yq7y3ztgCqZmGKk8UEWgIrt7w/v0vqpdOknNLjwFz31Y2vsdxjPFt1d2
VOL1zz++p6OQzjf1AwvvKKBvLOzfY/bRye0U+j5UYwwpwdMBpJ1KXJROgMArTvCYaBDNhp562TwH
N1qfFpK1238u+vAn+JK791YKRBRrGEJOig9HjbHekuMgwhSwCiODn/hSpykIhaqUoCnZQjodAUV6
HrLWRu9BG3gOPw5Asm9m2NeuEJC3sgjRbpIpBXdy/jtFI/xZM9zr9j7T11Sb8eNjCYFO9/8HHSu8
rU629uhXNW6KGpJHRWALxaS4Wgkag+aPUenW0J0xD4jItX6+KcrrXWPp8rr87TRVObeKEZ+8MamS
bvHlyYM3fG2LIUU+550KMYyR94sVDqcHl32ECw2fM6k/jK3jeptSmeFS+t+PzYsPNjLIjDdMLKTJ
pJihAG2+CNN3Wk7ppHDpys5uVXCMFbo0i5kSl5QlF9FtqlbWX0t6jPGqFxs5iMNj2BBzgNJtGnrU
D5fIREWBb0Abe89ITWWDaZqRS4peHvjDtqXSMGNhe7kOmU7oljk7sy+COBm/v4ASv6xG9yFZMFrp
uym/MD2ECEaGHIC6TWf1kYTjFkNVQOZjWWOQIMbjotGfV/kGeCOOm4H4epQaDuZOpTYGsOcd1qrR
sjpOdMFO6rn8seByfYPDDPr9c/llJAs5bKOaqbx8xrTjfseTIliFRezJR/IkIouJWagbIEdm21DP
MCe2NgpPR1mffkFb0WKgn4R58VWGmD8HjLHM5hEI4dbZ4aUMEm4BkZbVxab7Tpy/dYD5hJ5Wsu8x
pfbcdCCN+tA/oq6sQVn5mY1ywA7Y1d+SvoVXhBjowmbYYW2Q2/jD/uo7Lw1PKlr50ZerqumPKdgq
/VlQdcAaQL3awr5KDxqJFMbs+am64pJ1M6xZVPu4tD5SI4lnEPK7lSElyL3NgQTc6dwVeYWVsPGN
LZwupvWir9dLKTP7siQ1KXtLct2Mjt4yvv7DbpowikEl5Gw9fxwuhCuwIO6Z6BYttMZ7737IRGPN
AP8OdFlmKP5PpP5yPhJPYlPDdJpNzTCVgGM37wRW9S2bBXk9x/fNsBlZkU7OJZazARJwdax4zLus
rCxP9NDeKo/Y//PH9nQWIAD1FKYdO3FtXm28sHqLyfobsBYRovBdm2Nb1SuYC2BvfQAofjD0DH28
x6I/szhU3UPqJ58Yei3WeDS1qvdOQBleMONK2N+CygUj6QZ494S0sMmhkct31kp9uXnfyXwknhdf
eWakcxfkZeeKs9w/0ZneQPW1VxANhKgYuTdyZzw3S0w0VuFfIHv6n4xUQsJ7adk5O6b6RAitP+Ig
VymuIWWHCtq9/U/12FlaMAWqTXtQyPcAa6Vv+lZ/K7PHghgR9hN/Qe+oEENlNRER3FaBU89V6uTC
0Nkv4sK2N98gwXkPaHOzNHVASNRYJdn0Z0lObE05LWQHx/TKN2lv6nrXzSOivEExJK86J48Mb0yH
xCLsLJ/nM/K+Cg5q39BkqU9iRbG3HOkzyWqg0NMyo4tDs7vF+1p7SxJ679GMUh5ly8/VXVWijYAX
IktWL6u9E8QxWdvXNXsXZzRSsDxQd7PTw4lWHTM4E4QwFH7KwndJdugN6zANwnI4jtX54ZXnFZwA
vBn8mY3IUuGaucxZ3Jfq8Fq3MxRPXON5tAxRUsK3CQ/x3+gzBuDnL8KeLCfu5jxMR0OvZ5mookE7
OLboadsBsvVtnvfPWbkwWaKPiT6xPc6P5XRonuJbJgS03KaiHq821PZWpKIlBcVadpukLb50E6bM
hNdsMU6f31GS1ytCz6on+8Esd4u05qJUqcEJo7rYBu+OSbhQLDhcZXiHz3LC3kh4jNyZEqYSAF5v
TNKYTl3ZtBkMXnCRkS58tvALM16192bxjlFkz4/Xjyr3UmwbPLixPt3MXoKJGGrEwYdz+8kjHoEW
VVDyi4tlPMdjFx0LhxI3Q/V2j56wdIo1aPeFViAdGyuq83EybBaENFrENrGH3EwoX6aDRcsI9E6K
zfNbZO200Ji+j+Xodql4SESaCn4LQ0eMmMbhTlIPxQN2sj7AbqSQ+dvwloFg+Q5Mo++Deggzmq7X
JJT1tkQskyw3Abxsg74OUQsqA6ZcRJPFE2rrKRPrjrcxo9/Q5gyEW+5cUSuIqWO7GtBNQcZ6HD5u
1ucF8wh/ejLL7oMb7UU1lywf3IHvvdSkw8zNqza0sFlwkR5nNjpdc1fPbcvHaf6tBrb8rtQXClaq
1FcagwKr+L21pDASvYVMO/8y+dV1c3WiPo6QMBd7a8Q1I4Ie5cp8PpCoWB5i2DP58Ro+w+hdIBwy
mdZOC5MnCc6Mqz2/NYNohoCo3dMmYURJ6lKy24SQUJh2+FsJCA3/bAWuANpqQuDly/yNDPa/jr9H
LT5WjMxtTHSkvRLaz73IlR+2MLFKCEeDYLUmB4m829N9r3kZ+t1jXfr0KBh2B91CjxJ/UXIyZNl0
5d8kUZNQk14UOU429IEbn/qZIn2kY3NrlcdKuCQiYYOIVTuKqzXooKCkpLBDgAGCfMtIemd9EiFd
qPBnBc0rmnDFt8bMZh+m2SoFZZba5fr+FCw1BrO7Ps3e+u3BdEN3IhJA6oM+MiJCRuKTkVVzqD+5
W8yiO/z+0rMA8tCqqBnwdA+Ydp6eFAUODf/HiqXliDV48fOWnf5WTx1c5kTC51DaZMxwOXapVflL
80y5aPnOIyhX3GMRVtUhkHRM8TNR74XvDaps1I8WSVykG63d/64hotRIPy6dDOL2OT//G3jPe2lj
BL6ZEHeApujPl0HQuzT6wWXCHFXw+Yd3V1+GAXYKaHsNhWkfxnAShtM/o/iTH0nKBj89Cru5KQ+z
tX1s0676QxWdMPaXH8vDNc0chnwp3gOUztczKnPFPLnWmM18Kn0237Eq25VqggZ3ipNE1bHyeWaE
J3hSSwIgezlhVlnj4sFQMesQ590ahx9WplExHFYW37Z3Rp0hLoP5vFbZVUnQuJU/6Ip0/SK+XdEb
Rf3sIPZG/268ixBf3zuQg2MgabkWkBil4Ypl2zZvfDg++CWxtUiGgDO7WDKtgPRU1fDgygqQt0j9
Bqrm64GTJ/0vYCJRQUm8P9IGsba3w+pPDtWdwNoKDpjlj924uoFd0pxRSI+WuRL8QnUoZKFrVOkX
c5SyhJBsWfMiLWC6/HKYztZjc5DLA+OiLVyItpM7JoEPG01bD/zKLcVxDSjn8D+xnIcllNoSaHQB
1yRkSlJgKSdIJRMJPmzq9eeLKcI3HGDpTFtZ/oLA+03a/+V58s4dyY6odKvoufIPFwPbiSx0nW+e
1aeV4piqbg0eUfpCmzTspJk6Ze5JGLwEGCwK8C81M94T1KN/lksS18KgdVwzxX/Ho8mmsfAwqs7+
/FmX8BkcZbjiZ3iFqauaECSt5uCDXalgvp2ymXPruooJHHhvdh+B1jOoGi4Qi6k0o3MhtDPn3TdN
wmUxdKTI+oEoD8ssE8dimR7NS3aztR6FYIDvhC4fIVFpDEJJPdhC479IM2MUq2jyPt4Kjcmd2M+R
VsWN6h2FO6cCDox167qq1T2SfNt43+oVQwh5M0rA9eO7fZ28cTUSPC93IeWxGDMu7Jy00JsYMAtH
RSdbOiD/baxF4H6b1EzJGl+9bDzOpPZGYERNMOdkEJBKfQr+bn8uRpp6Mr3GJmpVSIow0Re/vzUF
UyXBcq8THqmRN8ANm2KWxyxPlc5S5+ubIGpEx2Q6ANpcyj5K6hANukN5StXKvU31uefUvko5DmO/
VJraXxMNy+IVi0JeeWoy4L0Z/sHOa3T36aei54N1RyEKlVbQwZrAR/EEh8It8TrT/0hZIYa5XwuG
ijEaJGwvs9kBVwVVH3TQrHcEOcNj0VT08WlnzNeU5M3xzIqBImv3ogvpeZoYtyuPuiGnvD8tQ0A4
1zCapp/PVsb6P5QJIKmLYCCe5B//UFkzKHaLkB0sMVqab8gVt+Y+4Iyio9+ZNksgXKcyWiWaz2Sx
37eQZ/0kGvpb+HIMyQd8/u3J0Q544l3FcD4e71UDE3VpzGxH9SesfMr9EmylexX02HITWD7lBL1c
eXWYis4GHSITYsB0haZtXxWgZKI0SDDKFKOYxklLg+ze/2nNmhB5i8x7EMeQStAQHN3d9Q1cOW2p
XaVg1U5msFlHJxjkB86Z5MyidqPdweUmg7jFcAK+G3v11oEwPBaaWWO0CT/Kwyt8admNf44mYfLZ
tEJI1gXwbd+NAIPM9vu/x74SDldj4/a06p/dxqKGLBHm18p2rmYDF/HXwIvKfXtlCOGWBO1H5kKf
aCUSMJ0oTTibyE2Dy+ipqEYvm6qMahtvUz3bNSU8BmeuG4VEibVz05qAPJd+iErx+WI6UpN+BugD
o8WW9+F1J/5zT6X7vrh5jqajqh2cO2juRs9gFrNs7pUA6w1YQZKmJYtUdFMp+B3imVCBsr6ir4sI
c4piJUhImKjRn5DiWvA6LUMKFDbDclMWQdxsz2kKW8qOTwqvFerCX6TY3KMnzKtTkRMGBiKwLHXU
TRhagqrXqbI+UDCzGXP+sRPdKjNek4GgSKBI4AIQSQhOprTgmATy8Cg5uGgFvn2hdsKVnx+y3n4h
xw9KTlLCwx+XFbBMDWf+mGvIH2/BJx4P1gyKWcZSIugU/biFn4Stvm3uwN4JyjTl1JxagcK5fEbD
sG0sJStiOqw/tqe+eZF8G+hcKBCLgWnAYYlwPKWUnOdvE6UByUOpaVLt2sV4ijoZERvKPqkWjJLh
o6H8x0aKAaFvAZD7QqssDYz2+O06aow5xmde7i876DLljqXB/9psfYAQOAXN+pXE1TzVU6dXMgVs
rl57O0DO8zANcv4d60jGYFFBjv4OdFLdeev0alt/QLTYMxaOFuwYihWKTlT5ApTdHH9BwQh3zryk
9JEMbkY7BtlSqOMJY42/MkP5fH6F6ySG7hPC+bbdzdTmIPznwMmuMPsRKs67XtCBmMwby0EDyDev
b6oiwJWTfgEYVCmSoBiBCD1RMqYW2qKvXOMpx1d2jOxyz0f5HT42AINk8QftO7ZzbJz2mvvnrmKH
FWomjE2QsM8q1fTEracqDrS7sxHKE8k2on1dsQ22wQCwOFMKFPHxU5SOR7N5vyMn/iUhc8lAoex3
GmcrPBna2JYl9AiLKz5NyLnI8f2IBqYj15EbMNn2ZkKObQ2xXUR72elIGHSEnqHSdB3rKGxb4+LB
3efJJRWGZTpCI/E/jezRLes6viavibglTyCnxWKUBQ1zIR7aymt6low9BwY88JmDEsCjsHqxhGwF
kBidsC0QNvkCZ3IR4K0P5BjcWTVZg9U5VCE85ROeVjnZXA+NCwU3y6VlU2OZ7yKxP2DzX+rqra1t
RFdaJecOg9Q+m2ixOmvGqzz+Otl6sbWlJIqDa/avlw2YdTnsFGGyVXPSWfUiwWnk1R7aPzmWEiqc
oUW/2xXv5likOUzdAODEWF+ijGGfHeqeRV2MxXMEQq4qKIt5mL4sPuH5jt58smgghCOFi/RuCJ1f
X026u0RITwBEjz+BGjPGUrzTvnLyID6Wa7oQf3svpkL/qGQqIyn+0EECn8vJ0H7jo2Br+boZnOEs
bTVin6ZFD8bNTtptdyPsC3914FGIXvgDRgLFgr7xT6V55iThZD9j5Ws+AJx8X4CBmg/bSZ82EZ6h
Ks8rGtRYdZkJIqTkwTFeAfZB8Y1w6jF43JRivDgWPEJXKXJltvYCI0OJU0JgCAdFaxRwsltzYsSB
0AFaIhoQkMqExDXzN0jkcoUCG6YgpbVfeHrdiBkP8a0tjdb6s/q8YddcdFAD01kwYjgv3Frt6Y+w
x/rAzaEbqlUdpurJdi/+GfpDUfqdaitzPX29INCk5pdpRlIZnzjrvXUEdSjw9YfZCug7YUkGNEwb
x+QhwGcxZZ5uvCGhtEuUUkIwSzxmfbkZfOjOm7S8mkRjImR9TqdHmFAHF36vi5jcWZ/hRYtQnCmo
YfGPM30JfWra/xbvipHnSvcr/eyb8QGunoUS818N+g++dbggIyuS8/X/zBfcdCw4dMNI5MHtXrxJ
6XIkjoMvXn7Npt1zNTPPYocERYxbjAKOJeVluBlEFaoxKVB/+LEbQLNjRiU8MAOhDhnE7djn1kZ/
qkPDcVn8JLxk31i9ob5AI0RxYiifPA0Sf0Oixv0iOq00cL9EKIekB2IzjUrQ7fYy+dzjJPL7ENzO
HnENJkjQLT7BuCdpXeISS6tEbUpd6r/8T3Dd35ZDH2lJTxp8ZURsv55YrLc9rBGUadktyIG2j4YT
3xCvYyk/PTDiqLtAIT9G+qGVrGH4f8Jpj3PVFJ/aR92oOW7X4M022Ujyd10qtFrbt05eZQyxQJjN
HKwkVFsPufHlfIj0MzH4ycwMojGfwQvwN1EFTdRdL2FYt5FRqjlCV2tGo+A8oLVXuYdVrINmZhPe
L68Hn1WdE3pIhVom1s9e2NgHDyK+cRn+YM+AJ8R8GyE/hKz8luLr4IC79pOs2IzmCB8LqbyxVm+e
ZSQA8vv8lSKfNjQSdfNsUomh5C+CIyNEmosH1YUR/lKpWOFdF6KwmQ4igA9VIWjv+yt47ksg1qZZ
NO+2786aaFr59pPweVirBFqS3hmOUtkHRlTJ/Wvrw21XsbHdazL4EPPh2eDH2AHuhs04+1Qr/P8N
HXwLFxL4UxmxQe76t5AFAvd3zFWpdY+3aTu8un3pTNEF9ht9ZQGDEkhVYSOOrWoiCnomt3iNGGok
r79qpM3DsPgOrlMUL2eLInBavFHuHB9KsPony/UQezDHePM5ERQt3WwwSZuM7n3LBISpS9158hQ4
dULcNbhCN4KT7vdV/sbmn6AK3IQ4k5rdh2UUIbpO8ggZjf3+1xiqN0+6apW2u8AUDFgh5jxPrrba
KXNZ30uS0bfc0Ky/lijoD2MDzwhW295c4reSJuFu55iaSNZxjn7scH3vL2x/UnsiZQBtp+yfnyzZ
xqWKNH6AFLE5s78+DDPG/UpD9MgsvdLywQqTE69zPbnzF5MycJg3HA/2RJGnAhXC4W8R268+TyOn
aVQ1mawNDjEPiQmeRNYcja3VB4Q+zwJedB825oyiDOnEE7zuv/sSoyYikVsy/U0LCYyhGrq5q/g/
lNP0RLDxtYmr2J4zk2APGN9oEsw3qVKzSB6lh7f+pCZ2xqqZr95u/7/xqIiOWzmUt/y7XKM2P9et
IB/EBlrH8fjNFSH+jQmGgnBWUjwlhablXs3hq67SXbSO4sQfB+RH69kkt4u3wFsjKbOpu83BvSJC
K257moVcFqGYGc1tswY3ZupBH9dE/KQ1AinmiYHJtopRFcv3akGKEyfAA3gGo9jx06A0gSVO8V+o
UTHYBh6UTfmFKE11lD9ab33MxczMcXRVUG7NawJOQz2NEu0JLcHv+yB+GcZ3rADuofu+b22795+C
3UMvEfP0xoYLXqOR/MwonoUIG5f4RQrXuiPpuyUfEMeOQt+f2sZi2F4igeYMzxP+tD1LkfSPSfIA
J0ID8lRkZHmlh12qyGLz0dEsEXOaQZzcz9nEisGzF37/NFTms6SxMq0Qn6Dhm3EPQLmFMGAw1LvJ
aJXqN3sK/qLoCPnX4vcYikBWXgsOhc7NhyOpcJOkX896cDitE2EX6j6DNPKix5Ziv8XYvVKl+mMT
5GITwK5miL7e8MyoKoiev8OD9WT2zdj2QUVM+XeyAC99YUuG9PRpajNlNZ1ozd+t5Y9lsYXgcmZh
N+apQ4oCZIia2PzSVdl1Jvig0Eeorng6HoU+qwJFATP8eM5l3vky3BBMLuLFPZQdTjnWYmW9/00y
pTVv0K13SJm2DFb/KXUbGsfMA2VKWLd++IZ4lClGsPNtipSMcvQ4nKuZ78wsc4ec57VbXHwrcJio
DiiTpTOuDjYGXAdVZueCYX1FElEG3k3KdRHDnR95icNBfKqjKpoDzyYXDKo/Jt6GGXMyxs9oliI1
d7AaHOyuCkAD/9POczCpJwVzasZbcpCima6Rztu2g3ELfYA/VlNi5XpqT0EMYapR0TJrAL1mQEoh
E8EUljl1yJVWcbVhxf6ODXVwdiL1hVglwviKu5DHrT47g35N4MU8LSb+jJL28hPqtdkvNKwBXVIo
uq3cnMcRcrPo7Mp9PDNry6yvErAIhn3SV1e2WJ19fW7PJHh7VGXuWWmCYsby7n/MZvI0D3RXta1B
2pRBx6AXOXcEtT4sx3WDJ0cKD8Oi18GdauqZYZGckRBKjAGrmjOQZnkXIAmad6IH8tDpskuWCNsO
EIrrWhseBYEpUBhYxtTH1VE5PX73veFXE2l/yo5/5v4/eh7Q1KSOtTmv4P/8/RlZE1poIcH6rXxt
XY7Et9zTvuSACv9RBKE9FQ8VW+KmjCci3Atom8l0oLNtdL+svp0Dn6Nea8EJkUaEuMZr13wfFEkK
DUMTooKWKW9vdd2W8YySLjenE/vMNrq1uPI4dVUgeLDG6oZL+klzmPE02/agah8CaAmjiqKXPOAK
RCnAX6RMaEarU6tYQ144cKlBflEfYORvuEwe+3dAPQA95zSWPOqQvcaVgOX3aKfeEtNt/O3YbtCh
+FRw1NVNz+GufG3PUJjTuPHsGT/sTH+TVyy6SpWjJz9EaN2lN8hml69fxCSfqYK/WmWRjo4khZnV
x2aKpzSN+smk3tuck4GD+dfQfsgXxfEbUDEAQxzeFIl7lrCDz/BszNpM9rHbCRBl4ru55XioRypk
hIbe4ukUF6U/ofiFgTAv/hG+x7rBeBdJQL490GT9/ErzgbSO8K7DQcFbODcB+Oy8mFaQafE6p6sF
GnesS1KFPDuVyDcv245qkYC4ozoG2+e6Cf4uYMTE19yVONxSmYJdzPiClmhdj0tk55vTnLyo4/Kv
bou8EKQ7DF+QkNPqunfO5b1ExpAB+Msmw+FwC6ydDcx7EkdpPpUcdgCD4vkf/ronB4fNXwX0AiOM
KHqns+yVb0mOQZ0rGTfcNqV4T6E2O+CPi6PWES3h3cGQml/Vu/kmzldOpWmrASLbAFDfg7CjyR3h
c3hfNu3udKz4t7A3ufhFeNMRQVosM7FapFq52r8ytsSbIjftJ2YCwAigMo2Dd/rGZsoFDq7cIxDK
OJUVoc7NlrptG1OC4DvZnujHQfVPKWrTx8qlVhkcqfSQLb87K0TnCgoaT2wT4ITiS8W5KVzNqS60
UVxoNUuraoNkhWxfNNIYqJDULQ1PgPBzuppvcaflA8r5yGg3s6W2GubD94bDcObV3NMuOVZxk6fx
DxaXRLQRBTrRydXsgQbJ9mIC9QxD8PT7usn73I9w1fYGUe8mPi7iv2Ew0kpxb7Cats9xAUXT4rJ6
LQ0hJLXcNxuPfe6pF9suXWGdXSvdv7pfnQCeRb8wdXxpaWraCpWOfp48t9of0d7JcNBIuwNzlGw6
DmCDejV6vZThgxZg/xCzz/lDdqHtlnWJKKtsVN5ecW0KJDz1GWjTit0gJAiElpAlHy+uGn9C04am
oXwEtAT4/COO35/0PEEOO1tJtjV9EPXHh9xLuRTWbAxXMOjvKAYbF/vAwVB6KM6otlhGLsWsuUVi
EHMOGvzcux7kaCVHatksQUfQ66GwyuvGHSr+q9JbMrLaBAhZ2OgZx/5Zgx/4d60OCNP3tlpIk048
AxB3fRB5SJTdZ1DQanSHsnkDhVHDXig6VAx4iivLokwYlO2QuVEwMDXNtL4FXh7WQHj9CRx2qqpW
2P4oljtdZvr+D74aGRZGeGXShYe0TQW+opRit+3W7Ei3IoA+o3Sj5nWy60ChoQwneoT/K0e1NSLw
zQYbZeIoHjOV+INbzcR1sTLj4PcIhO22xligJWasw0aAxC1M06A4VNw8MWYAjUbXMXOVV2gUHiCw
JBPIROjtY9YBm/wSsoyy0UTjklhra+XEkeufO+85Zyzz11/wx/nRlL1lCMhV4z/I2rTbnLGLcetN
hKcuxpEjPMxc5tJCspE9UubnVo1aEzSFReDoIWwH4nATxjSqYWK61lYnNsZPe1c7WZyKfK1CMxWD
PLtQdtUb6h3scif+MtTG3PF+Gk484KUMVtvYCeS7jqmw3ROQ4bVWMIJO/74zePBqyeZNyG5F8nzf
+OOGKe0s9PDBzyttYnF2sumaHlVlkqNEflMnArYCadmLDbyoI75Sr/vZPF3eh/YMl436i7KAe/uS
cc4AUGQJ+3zOww1jFcb0Bact4Zp9pbh0QUDuWgk0IALgmgAuzNttEWD7pDHKnIxtRW52tzJjNLKc
gDEP5blxUR2XeD+2SSPWzTOnM5p+g9AVs6B9QDBtZr8rq8p6xVTSGxFAdIouSQZEE98e8I83hsiq
IYW20DcgXXLBRJRvJe45wkWm4J3I7o2vqVVOfJSTt6qnbQnqLoUTsBXFNJZp4kVnOsI6Nw53KmpE
xyjRFDPtG57zyjmtDWSIfs8cIGP4Yy829BG0LlWkYQo76g49M1wIZOoT6oUANvmXHxgQVuMB5Hsb
fxu8u06dnJWYGSEUykt5qITuUuUgbxk4LK7ubwTqpPsWCnHfiTPBtT30+czGFyO9RKwdiB+aV4aR
nFZI271Tnhnf3BSQcWfjn44jw3+0f1QmpHScr7b0kFqic1CxTGHtlFyANhxuy7b2+s851h+Q2pUI
p0+iCwp5GILWW6T04ExhzjgkqogX411QAyTSNQqZGtKvKD/XM1rgvG/R4gqBv0pxX55b7rhRl9t8
h9c1cYr7An59crZ+Gb0F7g+P22JJZpbId5d+2ptm4V9GTROglLw3XphALagaZsrOQPRsCtovYDNF
0RTjxXf+eh1Bp0budR/VaaMFM04Wu0OgWZn6oFiNKmczXEB941vez9sMlwaNctvAgy2xnP1V8j/C
pr7ReTnzCPcBKVHLMpVir33U0kNymqYZciAr8g/aPlt/S9rwY4EYbOXLBOtiUvp6Su/z3rVcqUOq
CE7ojBwwq+Lm88OOtQC5IpOsfb5MciUqH8wWdMHHwe0Fuchx4efSPQUjCzAGOoe5E9HSzN/GV24T
dOCQZZj6s1u25226X+yTbexWqGLXobzUkiXYn5E9/dh9HDxMVNqTaEYEk1XPa5pQ4OMdkdXuxTFh
tMqXvF5kpptYKsW465Km93RJfRCs7CNeUz419csqVU9zPsjoyHGGaBTo7h7588YLH8n5ozUSKeFq
MDLv+zhv6xj9xtJvoGj6jQD1UnekUdoHemxCIz+ralT8+RenNgAatIwTU6ykuKCHtrtaTB7DPD/D
2syz4/sQnvUlR550ILVqVE0dqt3KXrWqNJINVDE2JRdHtcFv3xCib+mO1u4rFvSN/mJGz2ytRfpA
q3gXVQ4MrPlIMol5HnvVCyTch0PgfJhsPdFmgE5imIS+O2MhoNb3yWu1+hdSZ5pFy7AiZ7LZGPWF
waYhp+T2FOvYKGpsw2tKYGxB11O0L7xKPjmHhQgObQ1/Gsfnp3Yx2GReFh1oLVBjumuitQOt8BS/
2Vac91HFx26L3QpGn4fl40+gkbtn8S8EAdry2Wi0ur7geBokh8SVMM7jrBN1ankphMhCKFilrKlx
hhYjSih1oheXOeCtKE29QPxNg5fLBcr2W6RKk9bXEQVz8CQVmD8IIQo9WLwIMxmoGszAxUoCXFIx
cqVOd1B1QrpTwNxtkP2lYcLwsG/IMVGIpuC2Wyx+WFtCwusXwB0O6KyOu6eRzg3EowV5JDMmuvkT
z8jLP/S1MJ6OP7kqFQYY0IIwp793Jf5C0pLJOxikz2NQa4aldUtdeWZwHGW+zvjEEoWfijnH8Fe9
7mCKt6WLYbAm94KQbxEx5znT3+w/FTU/geyfxMhPO3czdvqa6Oap598ggk6RY40OSshbx9ARoMI/
68HS1JTqd/QG43ZCmw8CttGUbVomKyf8FwIVDJ+WC35kYOG9j6aXcLDgIrBsAooYhZk0dGcWOXVD
Vrkllu9mArCFmsjmPL+Ok7oflm7Pgm2WRKb9VU/C1rNu/m2dzMlI/+nAcLyKaxmLffdsVtveo/Nk
rU7roPTuJpx5uuWO9eb8JxbUNiizkQojMhhYCdmENihuLIlPzBgF0T3U/SwXT9vVesyzs4Kkl07P
bC4pHIb9yVG6Nzeei3FdhJ4iRiuLBDaiAGjMDkp+nJQfQDNmyf39qBRS0oc2zOLvxcdDaInlFqRh
vW3mO0XvqwK2YhnG4r8EOIioWXjywEELp/vTc+lSKPFQB4ZcHPLLRp0W3XR9l804ueOn7/4WGlZS
aJbv6zBZVIZq+E5aIrHTQPzDhd7J8l9uNBBXQKMU/r1uS3U+5i157WtaXSuRyWWhlFB3x1qPJJr5
7mOEg9oshZhgaBXngC2npnF6+gdm+QADUFAwEd0HSwnPRFbTuk9NwvWtrz/2ce3CGDvukzOPKdvq
j5XyftlRFoia6gKq2A1tLxVL6Q5JI7pmqaVeFHFdkl38IaUc+eW1LZvpH4VSe3nhycxHiTKSeVuX
0/sr1mUtXJV4tGgpK1qcTq1GuBjV15AuNvny3xt/wHZPuWpiEMQTIS/XjLPbD6/PuwTNnGezy98S
IFVbNsKfRhHe2XHIJWIe/x+hMXuxcAuCe/zrCl4vGLhdksPCYo6JihxbUD86q0mW76m5JM8TuSW0
5JceMf3660qLpfIRhaOWPvaGySRlPQPHAcpFiJGt9oTGgdXh0+qYGgAGL/aya5Q3GL3xsnNoi0ke
8Jklrg9CA+O/LwPO9tSYdCnAtzGVrIt1IULTqP1qt/hJd2gYu5/9Q7FP1ol/eBf9gWozImzL9VZY
3G/N6sA2obHhESDvl5yFRqycrQKDJX5W1hkbjbR8ZCaeRgxtyq20aGGpuPOPg1VYrqC4bE8t6L9f
D/x0zQxb1juo8khEVCbafNLoGq8C/P32WSNwsS0mLRmKjjh9+cYipxYyjdwUjpfw1jBpCZA/mq/Q
KjAgEFpfxOMeO8PaukZb0+eH9rlsORPlYAr0GpDu4cPp8VmhGMtCH7TepEJ4mHip4COlIA+5SMhI
DAwE06HOsvAYwVOxDXDWdSbBmhfcRr+2QcsaxllWSHimjl/5u84ytxHOHXDErT3Z4lTcgXIRnx2p
MIaiEBhWaRdlny+XQ8ZNB7+3I7+uTb2W98pXX0+mqu758fS3I7LihgQm0LSjRpHU7KP9/AWQ5Ic1
Oo3kGGmgUR+GHgGGOsbkWl4Vni0v2F86cTrYI/nHSv0cVYE/gwg+OSLdkGz716xGofoZcTcJCpPb
dNaLVQLRQ2JfwN4jfCkV51PENPJJT2x7QN88y984bqJtX2FmMe9UJu0G48ZeF6tuBVef7b4E/Pq/
9099gxcF9ggZ0ymflSkdyuB+ebdvVx9v8HSLqdQholAccnw8QKrZk9369+i1ma7EeQilm31iW13M
qEeFmcvenChFdJZ95GRIXj7hEOK1leGEaDqbZb1lNoxqJDfgPwvFzoGtxTLfusbVJ6Oj8CS24jdP
+m+OZKngQJpYDo0o/hOJ3BlJ+J84jb/yCqrlpV27TLIKOsxXAhauxuNK/onIhJI0YtmxaeolZuMf
2Q7Bnucm8SCW1MxKjfNc5y1eciJ57xiZxtkkUKOAUzh5jRRzQQmlNRRcKlNKHw+tEjW6nlNRO6oC
1QonSAV5HFmzqL+/gFdYcGxlPN4gHm9Ky8tnzfZAaznhg78IqVKGz+0SLcRPCuAkZ0nnqilcTDhl
x5UKuPEDbR5FFE2+vzbP/eJZvdHYGBdYdhOB/nHGHZJdyoc9KIGeb0RdnXC2cycD/bUJ+qK5LI1Z
7ETONS/N9r2ep4CVWHhbMjXdST7UTJf5mUdttmg9zFaOQ/LwVJsiYk9PR03q8YojR/cGnPTLBiEF
0Y4OVTHRMM2WvTAJMUS+rGYmU0L9AAkLyGRNwlvfJdq0BQzjcb5dlKL3p0BqUmQa6aGu9rBT6E6G
8PvbaKauBh/i2WBLAV5rpl8nNgeCL26Mz7sScAR2x/MArlBJK3LUm5Kph5qy7Nlw0m6zu6c2gxML
HNN0HQuCgsbj5C0JuU8g+qEj48FpdGto/9hJYfSjJ9I2zPlgXJ760Hjn4pHyH9kBSnzo7UsVtd63
4TkIU+XSsNmBCWDKx7aC5CKVj5g6QHjHEK510chfE90hDWf2Kmyr2irsDSObONYfRwgrOt5zdEmp
ihrG6n2qCq9l7WqEHh0hLuRhBbRqovuFOCtkzj4pCRiK9oezGB3wjLh+/BWR9TPZBqQ5eQYdqY6f
3UYFoykqC3uUGl0eHDnCcjvUJ1d3zuYXiHOYH25Rq8Gnvkrkwp1Un0zoOo2/iQd1K0xq8K+7M/Ch
1OkhbXeksCBvTEBHwbshBhWM26L0qh2xLoeZ+PuT1dzBb6nOBjHbFB9IiKi1DUMKWPm7428S+AuF
Vspk7jvVMGidcZ2dSxEPKNK8sJeL4m+wGz3flkVMQ9dmXJxbux4VDtIM0YS4NvdC85SuAEzqgjC6
0dNv83Rd9DkrwqlR8m1PoDwAuD64Ap7lnf17w0xZRhf8PgyG9gl3xBP2G78B+AbVhmmW4RxqllTZ
TDTg5wYxKc34QDzsD09xRqiQCazHAQyRta5a+Kl+0vt+xT88YBspGm55hkGetTFE/or2Cv5VUH23
ljttqI+JGz45tgYywMwNx3E4t85KwONdPS9xw7xGk+vKLxSexvHh8g59Diw3sAiLjHVbFTAOqnU1
szrSFkOe5M7cJHY6wqeLBiXnQqxGoCvBEjJxp20WB7D3qo+8yKUdsfDg4Ixnn46r28+qlABKxCFC
QWrR658NGIFikh4Yw2SVnb4fdn0Ka/+LvmLKb3BxUT8w12OqLRcXk9tJhs4FpArwU67IkaU2GXqG
f1Ugz3u9xH0ysQfPjinOKzbGD7NALYFu+4WKLbPI3JiMmc4q9ibvn8k47xnRbHjfy31+XNSI26+7
FfhMFC5hBC0MAaDd4S1CFhyhRdwM9sjh5wTL7p5WKM2aDvE93yn3W2oehqdN3ioSHECZ6Rv2lvDH
sjw192+vuDAwtps5kbh7OZnCD/bOYy3335G+IX03r+w5UqV8f98CRmXBSwUOGyiuGpWICHc4xdt/
vwqOAJrXEF9xMhS9GqP7VW7g16Rqs5ll8KiA45e46QLNDByrK50gVZb3MrNVutopzCiGO7WprTUC
5QlE2Q8zHUeGBna9r/8uNgDasLt1FCJEUQ02TGghceXLT9TH0RuJMH3D+W4oZCZbTW5u4xCmU8c7
SwKReqs9X5/5H5FX26bE5+dtNGZonbBDuqAQSpcbMWUR3+pstquHG3hcF21VZNaXkRjXis7OLJUi
tTNd1YKcPvC4tY9s0daJpupYjPP3nAgcp7cKIa7kiMgy1dhtBZeOgY4qnRMF6OiSoGzSxOnoA0Xt
5ikKxHYeZpnW0IA7vBfoxfQgKPUucQNYjWyYo0+SsJ2mIszufNmwGTSfMuxmJYPzKp6+KRSq7ghx
rAx3GMtr8te3DwflU7RtPUQM+kWrws25fC2G57ch3nYos3A0TWaeqNFKPwPNW/V7LCDstnMkDSDo
JqeNo7lRNY6057xcEOAWp3Y2dgxNlzd33y7L1ft7YPUYqQ29u7qtONfBYV1xPbaaJI7clNZLjcib
XAy8Qv7JN4iF1bwJQfrv/hgiFA86Ui6+yfANMoZ0lXWgzyDQRHtw/IdQipvq11HTrLOYrgiq+I55
PwJfFduHCVgSrG0rWMReKRTA7tlmkrbNZMDNhUe6fP6iJ1oRdsv8U+Yuw/wqgZ4bx/yR0+EeEyyZ
mkLr8e6XKKOWRjHLS8lpXTos6UtpkQXHCZDp4+4dZwiZJyHvUFyc4Yf9ntVpsNXKprmNSMoML+20
qfseEwTtdt1hSO2APgfficUP1KUHebtVqttXcedEP42pWCRylXHRwiayYR23+DnrjnvhA31/0NDj
ZptskVz7/EUU04VME2p14vkvV+CBItrvR8NVAItETQuj2HcOiVEjhLKS3ASnD7/yJZJpmdiHZ5LJ
OoPA6ZRwu9mtOxfQnHNee7tR7ZwpH9ZH7gQEp2wsslX7Weum5ThWCNR/KY0oIUbnNACJWYRWe3m5
oQq/63Q43HdSulrwWfjIVYYtZgTCRGK7TBtEGNGWc4MBhNmYRjP63cMzildAH+LYaT3kTlVKekIV
r4xezvrELGlW8zkp+l/6dkAutyzZRIyMXNkzdKZWw+Qjz8cj261xWE75eFKkhxWFiJSWbkPqEd0F
WuNf++lRIsWecuCxFpQj6Q2Se3BQ5YPIyBnxvq6Q9WdlC5xAWN4zMPvjDUDU/R1ehxbX1dzjWc5B
zBnLw46ViRMRdjc3+jxQq3tffDQ4DmAOm33d74JCtoXOUiHJtABvI4ls8v9JqqSOtyO3h5OP/4f7
oQWItpbkKr+6pvFZV9lJacPyQUfx+AFNINpCBuG/eEASXMkVuEZA2NoyCtl/O9opQd+TZMSxjLM8
KkpeGkixONrYPRowvNawjGY42JzreXGrQoB12C+Iu0N7Gw4DgT4U5Q/CbTZXsGKZm9SRuNe+095l
uUB/IUuCvyvQ4eVgbtCccLZtXat3+JB0yUmk7M861nevJC41XGjZbYqlg2KAanXu9tPQenie9HpF
2Ea49K+MTrEN9o/p7uUguHlXMPjGOUwjq2kzSk8CyxKhdUlNNXiILlfG5I20Z8fQ1pY6AiR7i4Iy
ri09GIsAtIFl0/VFF5gwAw7/GomxcNrLsL57T4t7oP20s1RxQt6kdCNudIySjTEkh+q42YWXMtvu
zTGZ1QJ6zlwnNUEqA1JfHCWgql/y1WnuMlVi4gZyfbH3Ed03VTdbs0Mn20CyPdzSmCzGYt3wVgWV
kbjFb88Sn4pZnkE+3zrKT4eQHr2juWwm7W4r7m99QHeaGDuIvfam9fE4u6aeqT48qI9Loa9TJpK9
w4Yv0hlPzoFu2lPOeu5cIFuRrd8xzIOYQPHLFn9xKJq96M3dkQZZKpik12kUheR528bOHAdXrxsa
jImhikEvCWsGP9MrTDcmm624iOu/i3fy98CKdnOOXgS4Igv8MeKxJzTeZcS3grtQmM82gSEfhEi5
CpQUg0OV9YnRO5vv3lvXy6kvEv6KVfpjQZ+GovIIu3XQ0GmjHkpggnJkqp1xtX4RtWyXFflOytW+
6D94ZMDmUUEO1BLAF6njhHyXbeqArE5TnK0sPgpOdFgapKnf5Vz9gDDfAJ5fEFX0SXr1X83cpfJn
ZvGEtSz2b+NU5vYWQlK8eElQbNMagRPf4D5D8Ba7sFut2PUCWfTKXD6BWA9BVhGIwBqbP2DrlVic
x8/tsTIfJ+ZuuYSo13CBSVrfjd3VPuspomSw30R0hfTR9pp/gSIvrffuViK+m4T8CuulVmy0CSXt
ckFTf2lA2+5RL5SFhw4awrrIS8oQID9A42RZ1W6Cybit0ctOOrw0EMyZZJNGuBwH4RM6JLMRI4TK
V3XidXX4hzbqr/e2umRrkvkKnx3jfFyuJrPbiEDGV8WB6RM7GXHZF2mvt7kCUvoeBR4pbOnsHDwu
pRTicctT05bzayQzSY0yg6LUPl5BIhNI3qkt3BBKF78L6z8NTGaoZNEPeRM0dDxKcZvt2xuz8eV7
+l+lWqmnAwmm9hcgru9/c16ofEF+iJO5SqQOlf5PUKUGkwWH6q1VWgIOqQ3NfdVJledTgCbDqsDX
dC983SUNozwr4DTVmF+DfOS7UeVo/izT0qjgT35yj9Yoifa2lnK6D8458/qzzpX1WO2nbiHCO83j
lOigv1P/lYzP7t7VaxLRQMPrtEKSzeX5AeV5u80Ouaqf8xJ4xaYuE3YQrcEWAXRBhYxv+0BGzyiQ
bXv8uC55Frey1ZgNA7KetmZ8JJCvNRnulxWTKy5UW6N45JmwG3EhL8oA+RDTrBuPAJZZZHJBBHxA
HvjCPUGst6x4yT9eCtNYhWjA85AuyDoAG+UBzmOFGVCl9soVF0UbXHyHuGk/g9OMyFdtQaez0Bxl
dbAc5M/1KCYyej91uIoCJfpJu2JPALmrAzSdo0Hta+tPr2z0ysEUmJMbrQlZJxx0SfK8ncv34xlU
6K1vC4OsdCM13KdOL5t3EqPS+g5qNDKuaH1sfAy8u3VviT+FN1w/et5v0DpKmj4PG90KqTRX2s+H
a4V83u6RNPJbWTNF6M1gJFQmGCYimJ3f4/UES/XSVXrv8OmGSG0qaZ2DgWb4kYGP0kccE1THiaif
25HkHpuI0u4qYWq2ERwd2UfPmByiNAkZ0HkJXhTDOF3KnQsypOaBkHqtwo+7dn1M34gkBen7ro2u
Vx4U0AvM+Wd1IreEsV4wwUQzR//hu+kRVHYBzEAzVwseZ03OIqvu1XFsQkuPaDyzrX4kluB1dK+Y
fiVMj2x88nBWTiu5sVf/PTh/vwFUkJG6aQ9/l8GuUgJTZEO2ckMQOKZTfCsmpWOfkTvv9n/JgBy/
8bLfg1gqzwIe8eDtE2PuRPOcp4kXc+WOU0srPavzMdPFTCmz/S2iov/hTRCmZ+FWC5hkgYooQjw8
am+c2067lcWP7GX7rPT7neKXvq/YxryYdLlaHObf0NLKy7KqdGh8cQ1XHK38JaWKv9T9q6HThZdA
1n9oDF3c8LrAFReI4DNvtJkwpg8lapPay7i5IVCf/1K295HHAcnYhkPmZr2Wk+M0jHhmA3vuQRrA
dzHHZidWCMZTy1oUbZ3aVdxlkCdSzpUO0ViT0Zzi/rmh3BkYQaCYjWDqP77Jb1FIN6tBkIT0aJHa
yfjbRw0wlzTJf3ngLmyh/06EZ7bFgN9Q26ha63H6MPnDNxX/AnihlGUeU11pZSbvq6l4dL96ySmI
TC95PREOJdfTeWMgfikJaIuqtsDjhz9f9l1Gsvjeyr07OH01iKbiy/ONx03RWpNb+QMtsaIiFURj
UJec4hCltX6/onu4U2jJmRYtViXnVzPb20d3zpaS4vMg6gzeqrpxXsqbtOK7kqLuI7kEubOrVQ17
Bu0oF5g9Ewr9d/EmZfN/TS+2dmOUONiGiLjTS6V0FuGc9DVSJ5/b7rPnE2W8lwr9C7WPPSN79UQP
NDduLZUZMO564jn7Ai5OJ+ds06aReXImkAx7HiaW1ukD5vkZTq2/SQNdbi7UPF6w4bWehBaTYAxi
mx9ar6wl6TpeZJLpDtQo/wrXvUSj0EQVyErhv2Ig1LRe5rpS8CtKBu+UzejrbH6XomYRyTX5xCPO
Kpqo3anCCkJC1USHR/V6kFDFuJ4wfuBQeVu1sH2bvY/Y+se+fqmQ0ZP/GGEbSoFm2YrpL4ZhpYe1
WczMI0/+6HHbXEfz62wZyXWxLYoljR8NyYwytIvlxPo978gxuhp6cjpBZFaVQ6E+3dTb3mWFstWL
sBRtnqr+flItPF4Plk1WLyQ9cmCKTSFY1QZK4qZ2IPOYlyVSDlgMvWT4hhaZQfDVe5HY1EXrUC+L
yHmr+5DJyqV6mhBm0B4c0r3sh3Jaz6LSMvbVVtifRUxjpYUL2MIzEgOAFCwRmjEIJjw6ZIe0ZroC
R/BtpukH0hZuj1voAZ9Esxjq/F1G277Uk7q2S0ofRye/G/CKeMB5+YY2RJCAzKUA3Wxe2NcwiSXC
qJnC57dFHJ5MmlRdI+3CXCJN88Dd0RJEUqDUW5+Qw0PpqdYtq/F66etpccgYfUAu68nDmduOqRsw
g/WGb8gVlacmGMpMnbV+wOTV7vNYGBTtl4CDfluPhTJZQob7RFvh/VBLOC3dAr7cKCeupSWnfQaS
kMSXYwlzLl2MoYA6INxgqHgMAzSuKHNoqikRYN4PiwKWSxqfApVjqsjkm26AddA/JJ5KVra+fX9s
xfGF8ZAkt8jgaucNnvRBESfXy271W1Dd9ioZeJ14bIUCc7JeK6jukqbUuwTJTYV9TZy1m6+ATUAj
p+Ivrr7OwBzhI/93SRuYTTjMYJWbsBsa9WhYEbfEl4wt/RjldIbAn9UawMBByM+wa+Jng8vap1/r
wnPR5lW7n5JEpJLjdIt/OfaZqWbCFkf5sl9roV9ktJsyIBmggMb8QVgvWQrJBNXe+nK4RrsCSM+J
EzRUsNyeqZ3GZB1qtCg7YX5suBmml3zwZ4fFSukTFVIWZ5ANRC4PEPAMwQL2bqR9PCEgrts311aC
CwtSoTT213WH0jhmXLtyAiV9gViEWLMmdaOpIxlOy00r3A25ad+V2jreN41yjcxQG4WW85wpvEJW
C2J+tr0Z527oj3Dplzmr4BYZQYCyEaCWHW4h3uzOTTg09KJMRYPYOP8QRDc+R7OTlDTbvmn9tYku
ldMBr3j+7yRP+SJPObcx7QcrmNLqeAcNu8uPxrUFxhF7GWrZ7ZjEyQrwljdY/iGDpeNiHwu67POv
LAT8fu7pVnD7EkpJLni1KqPJamG8WyJfbFbb+8f2Yi2vpu71eNvlExZL4fyVvMVaTp+j/rsTImx3
9bHCQPfE+wIzmEziNZoeDPd8LqLrHmuT2AY1oQtm4K5sgQ2v7BnaUb0evHoio3th+y1qd9rD1+Mu
Y9kBOTfaAZZFdwvCF8LtE4hSppptAnvQW7De2g2iFvB25wq2XI2ECcum2sMjpDwCpqEPX16x1btG
U7g5b5utKpm8moOLwCJJZKc0hKbjxuZXcS7QBvgibrwolrdXdORMH4Cmmp39NNcyjCzMnfTNF2iI
d/p+i7EV6FQgKx++8ljhg+an4rfR7zsZogoAIhczHrW1QSTY2RR/h+iTPu7BO95rmvKupVfX+JFk
ghNJdDK3Ozh2G9FsV8Q/mJIDPdUbevJfcMb6sIf6HoxtIOuSFay/pEAuDMoBCyQS7sdpiBgp8J8m
zWsjJzWko0+IPQuWlTMJtvnm4YMs4kKcajYeQ9GH6g0I3IjO8O/vcp8dqOeLCjrQSOohYpbG9Wtp
QND5IbmJLy6YFu4xVAcjEmdMYNLBvBLF/1o2QAl/5OLYRALGslkM7rNEcm3dEEMQE2CXpuhkmD1C
uDcGHNMpa/TwchL8+e7CzyYBTJiHs8cTkoVpQtSodTR9ZI1rxG4hiSpRdDDiVH6oV10gkkT+5VwT
hNoQklfGx93QTBimK4UkxZPccRrLlrEOpNraNWSnVXJ+6QwVCoP1KRnDEkUkwK7yleUlLArknr+u
bn/sNnH6vG3MOkhzIqhHfqoEd6K3Ik9s9lGh+SnX6GNlRs3LO2stjy2bPYI103Ry1Y2cA/XfCBmo
4KDOXqRLgXk0z8vGsFKHDv9VcF/W8pnAjWUDehzk0L2wyQ8oqdTv/W0KkM5Y/ZTPYYwLPVV806zF
GqbBzlP0ahELmMWiXw+FEVfa9y+K4xrbNnsSxWgtkwuiXXJVM9kLxppX3YTsA4nWjoxkOdZuDXdh
azcc70W7ONMMmUZAyIbWi4KSOZtwSQ16lnxx4M/hKx6rsy3UlA6ibOvCiyr5eHr+n1YBCBkW4YmE
jzLgHdwSwXVHihkVOKmk84S3ddM+pIW727P5nsBs33IGBxjGLTOEudZptjY5al0ryF6FEw10ZV3/
O01njE+VBS7t4AOxqsTbl9VXJW2VuXf/8d62ttk46pn5EsocCs3hioO7+FCY+wYkpZech2lZOt20
OoU+4OKC0IuCEhjhLoOpmZRPtxsKhiaKPGM5f8A4qucZT5qOySI7Azhye0eI+I55wDKMGczFl892
kIqA+u4xY9oeNujve5qzkgIkazYHRSe1TnXEfMSJ86/rf/pXwO0+0M/GV2R/PJ5hUf0uJfoloO90
LoKXME5HhsDEU+QepGb6E1qdUgzb1o+Mdz+EFDbMNBb/0iM8a0zTXhwz0YoLOpgb4pR32NRhtI5q
RCd/X2J74GTgkTxNyAyV9aXLZPGEg+6CmdxChNJN9J1HojOqIO4N5BPWMI53NzQ2jE5nV3BnVyPe
pkdnkk4a+VRIR26KDnqH02PLSDZRNApstfmWFdOIGht4DbLuUgb3D1dF35KrHCyvsJP5IVKfQQsb
BS6oTBmDrUjWbhndYDUHz+wffG2uk4gOZG3mdzJvzvoXF7Gg0CLQLDAdfjHruv1xGZTR09iP41Xn
fjg8AcwoJ87o9mGRkRLey73bOZADvIyPRp7Bq7k3vetu4Pwnqh0wvcNOHhK/pG/nMk7UfER4p81e
ZTqtJUKX0TngcJBB+mkb3jeAA+246NeuqgIqWQFHC+mvZAKgthdMOQ7FUq8iYvxQlq9SwZiGB02E
DisP9s5SIPMzG9QRRj58V59SQt5UUg6662mNEPEZQJapkuetTpCocwuP2WpjT10W1WY2v3yQk30m
CAf9A93HEQq0uc4z1IpShDongkgntlDSOcI5ab7RS1evGdn9IHYuX5MK1n8dEf36Vth1e/HBUUO6
GnW1WgrI/tQRpixrLhT//CTXhN3B3AfUlh9hp3Vpa85oiUnAW3if2AtyM34e9xgkQ5wcwWkNpJQX
jgus78TYIm0qaaebnGs67BSDVZEiZmh03amSyI3H7tnqXZva/OGnCZdtpOb9U4W3tWnplNuN5VFv
n60MDgsG8OX1krz6IbN3CafcRHpASoZqWge5Sy9euKF+HDsnwqqIpNBhQ40jSyR7CCFvA2a63j7f
A1IGxjIHvNg/qozG1U/b9UBT3SDSRzQ7AzN0WFAEabeL4OaBwJ3S5wQsuWVHfK669ZUGGHcZ0qh7
6u7nGvRXZDdIOJC1GXB6+s0eYh7wzvBzWALw1Blm9n2DsS6C7KkZsGkUkf0BOjcEwl+DEcISd0Ur
nsoE7OM41lgAV8v9BPyRCPB+XHpS7cZtLltl+9Fswq28VdJ3jqEO4fYrsA7qtJcN7eSVndHnV4LV
Mgopuk8DBTxPgsRd1yhFyZZnpTxKk7GqHlSiL2zxDVrmZYh/1EjmUmb6O9x3HAFX7lc85d+O6HjB
qV26cBgaClzjWvoiVENYK5UiwBg7IKzWjNqVOoWwzrMNW0YZhaAIzCqfEKBkPmBpryrAEpwhVjNE
B2m5SB12Ffr9b3nRRVIj6SMudjfZeIf2YrhERWp7sKcAhekg6A1+YE8hln30DNCvgm7V47Iil5WN
1XrPVbvueDuhAljuxkfUdLcdn67zrxekzYMpUeh7tOSGdgm98l+v6AwJH+iE5zTbYvmlxMIkg6Ng
8L9w3zJ17bhtTFQr6XxIa2LURNzVqMdKuzTbN7yI4XxzTB0qawQiX7tZOHhmsnydG/x8TfJE8dhs
8W7KnPwry7oXG3GmZETiOdWRWA5BmYmbJitiM/FeuBFmUp7qUQxDQmPx+7qnIQuMwqHVSXOuddJk
uSGk7+pGtCYStXSVA+Naua70wcdSGVAOpglilOGCv0D3Gk5hi5peqoDffAgSKHPJR8IylJWL4j0t
hjd2BtiJJpH8BGTCk2gHM+jDkHrM09lk/Q0Bff6FPts3s13CCui9HCtYZc8Nm6i3cuu6maYjsRdu
EZT4k2TybW7hHxM8aDHKsmcSdzMzhjapTRkOc/cBJt0AJJwdRbgKTrOt6iQsGLcHP62qjVipKBoS
8tGQtQ1bFvsjjQuORujLib8SIE3VIjtOW3BWLx+vlez3iVvAZGKokbA4xSDTyyKIrXpG8O04N0LK
HIy2KNN8Cj/95bqd9rwGTKVz8GtvGQQN4j7g19bxGZHCj0vnkDBJgeVMoIpcRfpzfVzsh0MLThhG
XH/8JdLzaCIqdGKa6cYELmoKN2y4zfLy6Ocqjf8zeLnDizJgScFESiFWlstKEtae/lcoTyiAeaZz
kCMuM1wLYDZueeoThl3Mxt6CebGLrUM12EPkF79BPdYVsbMHWAsbetP2jMm7hTRKet7BSQ0/FslT
TTvvuTDDSuTDZV1NKTcgKtJFASK1qhgdzGJy7bXs+C2LTGkQzvNQUp7AxQcB3qsT75oj+GO8VI+X
JceRAWT7DsDmXuifrdM4isFUYy0O2Mf+qMc4h94kB6hUnzE7DeTWSWudx+TEwhjJDpCZjbHE9b10
73X3imjsTkQ1V7zZHbtfqcBdu2J+j2B7mCgMWfFYtW+Q3PFBoHVlISttRIeFkf6NNxdP7QCEPiKU
+2Ek07N6LERBnNJQcUSxsxJXz4g3VQYn0FaD4KwknQoxbm5mj7Zm6N23pRAtpGS41NCdgeCmFKkE
RB3g8IlA/X4mK+V6aF/VE5rQwEq6BJzBgY6+91IzJjq586f2mMJucEPneDFEEPXwrdPcu5tWg3xT
xDfmHfqWHMtuYECa7Z6U8dTsFmcJvniqH1szHkN6wV5o5PIMAlvuceauMM8XwSBnRGQvLFuMg9S3
JkDfkn1WM6KNdlRAZSZNcVrFgUl8GXaE7YC/wx3AsaS5ECPhWOhLuq4cwpvdQY49jgW64QEdlCDK
Jl5SW7VuE+Fy0GdiMg15bNGhgafBSnlaGCrBW4JmlwhlA9qTdBwDlB2N2opJBnMTcbJTMBVfow0s
ORG/gacBIVwAnNww5mHqIKYFFGrMfEJ08O3NE6XenUCcIwnZ8cKEghMSi0luaTKB6KlQTwI1SUi9
F5FacP0HSL/DmAeSgEX3+mY36c1WQ+XV1CiABF/3s7K35+ixbUhVKuTbGKRqqIJO+F7ISo9E8dJv
dMFQ5RdhG4kwQgil73O27HznkHYpP1WvQ/6h2+O6E0tJRSYrV5aTYrOSUZ6lFhe4TsEbLBfZPjtZ
y+ytu3+/71tmkqbJuIR+JLEhoVDpv4O8oC+bl4D6bP2hM6RccsT85bSSCImDf0JV6exPq5wVdAiu
n9zJZcgpDMIW7eo/7v7benUOEvkcBbGvlAuJDuLSJwDS+o+xpssReyYUWlddqao31NzKRTxt45cG
yovYM8V+mRzxOdQEsKyknsBQwdeyHraiRMc1d+SRmuNBI/lav+PoDLko5jq3NPqIY96iWgeZLteu
PKntU3pd4YhndZ7OmuXWtP3ee28lRDs1aefCS2SeKIb1SzE3+HKPjPKMq7OO96h2aE/sAaI8jSPI
reXsoJVLv45rEakBlh5OKKDenTn1vG0Ns0yJLEJ7TiHznoYfVi8H4+zRa8cUYT5Xe3mOcZqlej07
AMTDJ6w5G/wvhJHTPcxyNnmk1wRuD3vDFvMnBe35ZLX4qY+hwTNP7oaGGw+3btQuDdrimVIBVPMn
OiAD6cc5Gkncb1SfRqe3f3W+16XpmmvKRu7s5rYlOH3jsX5dpUmZJAY3samxWetKnov/yMq31h6Z
3n0dm3l5AOfX467fCw+DVMXSOPvqn3mQRlJvj9at+NfB3UUkT2r83NRySKK/d1Dy+oHiKlJN+9HC
5f/xjcUrH3FWnXeACTfWMl7M4rx6mCcaxHvEdCF8t7jVa1Yj2/u9GIX2+OdoV7N/GUpeYkqygX3y
gswGicpgVm5CmzqU1PGKZFr+n65IACszzowIo0cpm1w66c4GPKxtmQ3Yu/IzjFH3Mt9SamDqQkc+
Dh5+BDrtYwrAfDvp7eQhYsWioKuLHGTPCaDFQr1wihT3swPa3F8nL9DjvFd69HtYOitPL3btWusb
WUxUUv5USCfhGcTINxMoOkKRflNEvpmAn5+zkEqbzThIFORfcdZp2fr55JUAZKatH2wQgH7iniI9
FJatdD7RnQO+xCNVx8lRRg1k2F9r9EFYponyIMy4v5kHuR0KUXCPncBk/Vnf/BOUBIl3u+eveSUL
GIxfjV/UmSGNjOIgNj0sDgvi7lGTmSaEWGM5uR8h6pcDSGacrEeCggOnQ8XJQz17t74bDWO83K3x
5R0ykBtRVM2KSmnr8APaqWKVWnBRADyXxqhPGDYa6yrC7fLSnyIdgZ+hSEfy2bdR4SN3F7YEJeJn
gSs5dvqlXX4znF+M76vUZ6JbixVLED0HI5beZSqNUZ/gVysPgT50kBoWNKrtHEwh3PAXM7WyuZhR
injX2U77j5KV7wMBTRdnRhFIhKEJ4jpzk1VVoE0QUSwg/Y/Du52Oj4lC23JHnVscWqQtQnujPcK/
GuegNHYtCp2rZpErcqco+NE99DuzV76gZkJsZo4+3iCbjrnE8AKD/uIlWpOCzqJDUS/l4fL1vIez
awQ/ThbPj01Hm1XbVL2LaMgnP6pVDcCzppxiuQBMSb3JmUXIKD18MiEfASHFsO9iM4bbIWwXtTAQ
TvgYRCaet5ocq1icoomscqlyTLfEqnl2+bXU+erUDLvIJFFcPlQ/+0WVTdvBvzMIPB4UJl1NLSxJ
lVkynq6V7LpHhcSHdVae1FEJrodRGVnLyIB9AJ5BVtax1qyitzgjq61G6Pj02ECasO1R1qqdSqA4
XYc1RGdtUpMLrKvoDyK0y7attUzCVWBXgO9zWXez4s1mvS/nSqTGmTme71SxrhgtOqXQWOusZnsE
pJCIs2qMVG6DTb9/VhFqp34PJnp/kiqMertaef/MCZJvvyOOEVFGLCCy16Da2/WCGx+mDGqucRSJ
3n0UQdXlYcwN+Ll0LohMKeFeS2hyBhm2NFleMLRh/kJTZtGlOXlE5ekfrGMSAsgaQZWfTn9ycbLB
3sBS2Ou4VpBd8fhZw94/JioJZO7ZXJuWtyU7hZSEmhKJONrbOPh6AB3iHCwMfQLzN+gGEGYKk92R
CAon4IEiKGP2WZX5t+b7NJcqOdd5YSvxEOXHzd7fq7j4emXHLxUTOmwJQrmCZ75wl5tND/Y380+Z
k1rLWINXsQjrwQjPOuSEEWM0JMGcPB5m8V1x95pKOYKWtoajm+5qOj+DjWHV5F3qn7pJf140Gv9Z
YyXnwtosbTXWvgDTrk5VtQ4FFP8MLYfgTDoAkdeTLzyosoRRl/ngha6rflpmiJfcO+UrG0bu5xgm
AeLK0iWh836qBNrqfekISrKx4rDv9pwd8Ejl4RAbgKcSImPgsZY1INP6JSnlG7CMncD19TS1Gdja
+JMyJJ7prCXBoVe6V3yXOROtC6XlAaid+46/ATTuVvBwVHlJw7fw2u3F9aC1WT1GrO+B5deL8X6d
yMuxcFfdKxo4ZoLqZYdancMuLguUiTa8xNiTfAGWmyKAHJgfT31ecDuRPzWCV5y+G0Ujwt+WuFKV
S0qnBvHJoS0Rwq4Nus02YAcBDQUZa2TZYIffDAhf5WjwthJdrQU0yOkRWuMQnyzTGhUk5hy0Vifj
ArPX5gQls8Pao76TMv8PcAN4lMQbZT0ClWp5gJtyjuHQ9PdDumA83rsQzC37ihpVyfXp/BqvwlXp
GRYBx/WKLy5pOUPzZdlQrwJ1PKdzo/e5dn8B8Yf7yJZA9UMwt5fCEKP1X0UbMsQtfSOpTQY5h4mq
vLGJ+6KOph6jvQHJcOZ3YxtQq+r859ICfZQRQydap125NKDYeyfqsIiy5ApEaebI9Oh4pQIryIN0
cgygpivwvNo94GXXy/QjXOKhGPNgyOcMfBvXtHT8KppsEEF+UQvBOsYrPsJKZODWX3M6T2eH8/BI
DNvGRro1Ikc9wGAMzAGoo/NuRZ80oAzBCRrKjdg4CaE9Ugn7NolFVYiSrnvj3RKXV07kvPvQHPCu
WlXyTXAZ3GUODvzn5CIMNL+Cy371wp2/i47TwknFWLoCZQXNBFBRTaFRiIrq0G24C0fbQBHQB0O4
jZSMK1cf8LWF//Das7w/qvp9OMTcJax+5liFhpR6vO6T+xclrPCjIUoA1P2W7cPctjRNAzmiiCV9
8yy1sn6+E95ru6TqJp34zihbzVJhdD3xcXy7cQSVK25tioi2o3KXPjg0SxrM4+GitULAK9uJy+YX
uPxiU8rQCYJWKGKvGI3FGYS9Sw25ORDUqxgpvDdizoI6d3cYIIYjI7swKk0ZVF2lZ+YeUx/gY81G
odAK14wInrNtodFwlOx+NnIH047Vgj4BxZadTUv1JbKqs8aEyT1hjFJi92pr/UGfDoz5Twx7Gemk
o2rDO1K79ATzKvTRDyPrMMvwNMGc6AfEtvnwIL33ER9ECCRhebcYJUNSP+lUzoeXNVVDvaO1u7zh
VzrYQOpsFq2s7UkA7GHuu0KF1rUEec55FPQ4QgAaNrADHpEB6MIvVqNs9VeYDhqQ0xqFX7VANAw1
PDVGTa6JOTjfaN75YdqSM4O0PG+GZA2gIK+694U0PY7flnAWXvftKzaiZXh0yoUVT09oNUnj/JC+
k/r9kY4MrdkKnSvq7JVVZmaOWlXcS46jkSGSqNkHcOIBYXd7aOnwNpwQQgcdStqiP8YtsdhuvVMI
Seotu4pMFCof7+tkF5MFO66o+fAmCakhLPgo9sxGn1XRR1GUQyU5XCKl81d7NFPzViKp6xcvfRNv
sBDiEzfiE9K3u9fyXwUQQbh4a3uFemIr9qV+f2f4hgsImU4/oN1faIS4YiIg/bVOR6Cav43D1TXm
Dcl97DvNkR3JeOhcDioBKbwL2VCMK7bCgdJsLfjaZKw4mvOURqQSu0nWl6IHaW6n+qzqZBDWnDRq
fzu6M4Z8P7l+nNJefSWB3ejMXD64r+Jz/w57cX3K7EsZI0We3tk9bRdeXfa6/JnEZ0p30OJZWPff
aFzNd+vusszIWvIxB4fkd83CgeqlgaQ3hIF9gGAFk4yWR8TDmWrAuo7rvW4Q0Cz4NaxYPfc1WmIv
t5FOCi0nmnpppOemYYoOUgZtdV42/s1l2XxaBG07OeFFRXJIRXurH+i8Y/CWBK8Zi7QX0pQNZ5ep
Xv8uAa3YsS8D+jNcBSs6TMw6UQea4jNmUUPd6NoQzop2bX7IQD154CnRpmfI+GwA/OjuZx8vXu4j
81XoneI8AtvtxFhrO/uWBWNZiWHdeRGgfVwgZX9IKM0HDm9LdHGU15vAo5XjTxqzVTfU4pdOZA9Z
j5yOtVHR5p+x3xyV/a2/k4r9kY66JJllOp2PRgZtYqM3N+kS1jD4YINUsuNFI3TUw9bQLt4g94V5
pasUpM2NB3WrbTikjcDXxfcW4EjofH4nOdcSO30WcYy05hxbcJonfjfux0gWgPdF/0AsVJx+cLrZ
NCrSG0r/88QQzMY3yclU0NZmu4fJWQSSyDcbDiGhb1FeJzAtG1crJI0bAUdYvdO2wtQATSpOCeSU
li2SSYnBHVt/pRKQCNV9tN/2hmN/anVpuD1GWXPnLNX20j2q2Gf41d67mRtysrG2V4yMJOwETU35
4GndwnOlpEpenNoouo2pKqN066pnP6Lmecg7ukH/8SBjjJ9CzhSa/Mm62+XkU3F0P8+N2QQ8TmJ3
8I2X9+4ntw7jSe9qcqhNUtgVzx0xq/KqFwjYhhRKJFzfERg8kHdSFpa+g5ycwgcuQkKMdVxFz+IB
9+UxMjzpmQsTpWAQ2fYjovupCd9cy7iJsrPgbmumWcSWbbPeYvsklSB+td4UNJ3VYm1gnq5icmzx
/PqHFI0THk817vHrK2Vwd5oQ6sVJxVB+SexJMEqDVptH31NE4HNTX6G/bEaDCaDk48rTmYTcmq04
WS+Deeus+FyYuDorNIDd7GIBg7avj9XYQEpu5pDenVXI1p16vGRMcjwi3o7yzLJSw0HSqSvY6PGC
ktkuttaHY0WVYv81stU40EVzM5eoimNMW5nyVhNYv12jCl+W0lxX1n2ABraT8I5PBwy1YxdL4edE
ccM6xC2dLxtammSUH6Hd+qsl0B7BDVTeSKRnValxm1+TQzx0g+XYDjYA/QioY82cvamZ0qJzQDuc
ShneGaPlZfSmXrjJGfydg3ghNKebNB4aV3iL0pMPEhqyS6TxjIK2EKIgW8Z0pftyIVEakkUURW4x
uRPIk0xb/5EzRym160obvLhXnntx/GpY5RjVXo6Cfz/gkl6W2oy8U5919kIJ88lSpN2/kQh135rY
bE7aAgm5/cM1pOR9o9d9rR9QhQCIvL3Ul55V5VM1Ax2V+roR6m7y2AYz9AFSMuUKyAJWhrAdz1U/
hkIz67A/7521BahtRl1OQQcP51Dfm8DQ63mhyTz6QaaPukzAclqG3dCO9eBZqqGkPJDbv50rOxXX
FoME9URlmfTmyblXx79hcV86mfkn+EUV12FkpvivYtGJIoFdY04FEQbEPoFdVeVGdm9NazCAdYzQ
/dalvnznAGMkmuZFnoT4l8FmRvyRCnGu2Op7xXMHJEMPSksvaXCKP3WKYYxkb0xZWRtFU3pEkYir
PNmZl6Uq/BU7TD1R1Lkm+etnd2LT33XS58x2RkZr4AmGU3iYO7CoUZPnpT0wv59Hrt9Ain78un7y
m92amouvDDad0CRQtIzw4zQ41IAm+0JSThGzu5T3GT3MGZ+dNSx3IVnfSdfZCzVbI6UvDeUmkEEJ
gwqaMPiikAvaMrcOfhczXzFaSsyH1sRSdcfz+pf53/55kzPF0fdaf5FuC1ulvS/TgK1BWK85Z649
YZoctYkEo2mX58J33eSe2CLQckJ9eC9nolqd0r2B7FjRlquGFGi0ulaE+7+FyidB2a/AIACgS3br
t8ttoY8iZFcriJ+W4JzSVLg5utHflddL7Z3jZjnVuQvmdhd1ABGfC+zsfaIonnFr7UqCLuUZTmlH
irKiODrXNB8rsRla+PftEP392gvHNKEW+3J6+k2arZULpY/65igpx1WiserWIV/FLDz5mjogfFph
rmPJ1QaUcmO/ovcXq4poF8B+L1/T5dGHZmv8CkGzXtHLqwKyIGivFXqJ9CQwhXeDikignqney1BA
a9HpiYHiX1jb42FR8xrQkN29jTnxXlQ9TfGhMLbh9iDMjSDUJ/T/hD3s6eokGSSgJvV6GVCB+kIl
60v7DHddXBiDbKyHKi5NKTHAavUhaNSlIZmY6Dx9+nGP1iedbC0GWq/7Jatzg8GGlBzieuhHfbf6
rbugpTpvGBkvRbD9SSPG/MZ9dHj88JtEJoj1TwVVnQfE1s6NX3KnhI0lV7Ot4ScYbJaDHrxGFze+
KZ9la71++si8ERmIH/9Pv2TepB4MaccNEID5oB90bI8oW+t2OQtNaC/2KtOfLw7HFGH5qMtPA5RJ
E6F8XrITaveU0OTbMiFf9Y9GQoa6gs2umNhBQpP16vSInT9FV+SVcZab/M5aMTfE9C4xx1gmzv31
wPcV0Zybmh3ufKsPpkZWzbrWMQeTalHvAuZ3ECGFTLfHeCUmVGM+TMH1LXoP3sxPtU/PIaPEuRU0
rI4520hR+ZNI+up0vKfTiqc7BEn2CvDXcdVn0Iuz7aPEHouFKjWVBpF2rYF7npJXi/NokiuQa3/6
MeJHI47P3Jkwf6P58rgsxibO4SuqDbF7osNgsttKHM216fDnAKQaF6wlpdUKp+7nemobyqptgCu7
jVHL3HE1F1sCJsLd0dq8ZG4SsJ2LxuduJH3caTYevNkMCCEcpuYMt5/ADRMUmCwnnW1YlrfLdBFW
S75i1gxp5oNcBobBHQ605HU2sm12YZtvtdiNv8hNV1i+9YCVOlrlY2DPLPb2khTyeF+/sJQSPX8v
z8UohNWAZ4gEPWi0KCu7nsmx5lPlfgBv97pOAHs1JnAJoSKstEBYB4Xrz4XAEw2zQ/70R5Puqu6V
7EYTL2wbEsQnZbvgb+3iauw1SbH5/3SGr+iH8j5M3jb8gmx9eELQIge/Jee3odYBOrPKJR3YPBL0
ucX70fUtwzepllDlZjnP9C6pTyjRukISJsjQLg9C2RwrJkysY7W1TrGQHxWemyjgdEJVVNHfjm0l
Zcaf9bSFdAInX3o2cgDGlSv8a0R2UQJPOo0Ekb/+FaBMDr/NaAmyqjsUfr5N2VOMeTKNPGRVvij0
GuelvV+/dADGl5a0FMPBde4SPK0ODR71mEuRhDxBE61YnFAKp/YECbZqMQQe9dlE05omCAhocyqS
tNLED4pR2vgCObrI4mxBc9OELaT6PXewZA6uJvVnjz2aMMb4lWgmoVTseL9BCII5fxcsLUkHS0oS
uRksh9BXrtNPC25AKYCfr4Gc8nPJd1EaXEFthzj9vXmshjLrdrND7mgMPhwnfi2pvE4FJujUd55W
IhhSQfCkIQDVGXRgDdjc0nB7LwFkgDQO/4imntGo/B4htJnEfG42Jxxg3budRavKaZdtc7DsWjJr
v5iFtx98oAVEUHl+1RoMPdDMRbi3JMqkaGSwhOW/YTKYWi/lR9hcy57WnElcMaf3Zv0Qo7jTT/0i
n2di/eIeeocuayZRQdnaOeEeLyn4OC8seiopXjVNr8pyr+Yu2lqFd0oFryw6ZWb8Izhgm3qnXq5R
GdzUSQ7Fa2WafvPSQWEzVHKNSCq4Bhn4rKINS+geUik312pTC5/SCwnNmfzBHUjR/VhRPDq92zB7
HKShcL4Mba7itSpGYRQInfRHgX6OwIoCQih/g4fLqrFhTjdQts6O6xnfaENMoR+5kK4YADt+kfPr
VnkBM+W+9WJ4ukEXthLxeDmqHwqR/qfAN18qkgWJzZWxw17ePBTEIPjXW5GVD1FeC5+Q0Z2pT0PK
Slja4aB1gDZT5ouNZFK3wTWfQVl6jtNTkRTSJZtuv6H1CkQbqXFejl9uBuTXwSHigU92aA4h92QI
RVa1o8thJy3Q6UpU3yebs+uHdMxqJzOBTTJ3r2i1TQzzdzyTNhwmJc2HeLaZXh07buRmOwO94/0M
0Ydq1BkqzpViRsuQfexg3VNOllcKL5nANvWZipQSKMR7R92L7YPKOVpXyzyAXTUflhKXVpxI1XGz
ANjWDe5ZjoOsP9K+3NZMzzNlxCXv/NkidfhrCbBQzVhfcvoL3wqPR2wc1R/uOuk+u+6HaaLhznk1
5Mof+hXAg/rxkCmxd+i2EIE5Wod3+3vW6tO09iksOS3+K5Xw6TbH9O1JHh6tlSvq55q8O9Adg/sL
5OOYZ8G7+hjrs0GCDab0zFevTa0vFE+wbOj5f8pxZs4uyJYpVGxO/lfBb+0XCJJWHnhaGEXApJRC
ZWrrJ3Qvsp/Ucia6SPuouGMibhSAF6cXDm4GMHNpdgA45JMskoWLAn2yh/yvttx8WUWhGl8Ucpv3
O9pl/b1YvD+orr5dzygSNHD+pxdJzAl9qJ3pQSM43obtdKaUmTHDn/z6VMUlUx4nU5xjzeSStHxS
NjHYV2zdtoD9TJqoTL6yHvJLf4ot+xxVR3A07G74eOqgjpnpOMs+VFBTERgOSDqzuwCWmDymuHGs
Xvbva8EOhUf2FZpK98P6dyhIT3duOHbJaw0dpHrxfF1D6CERk0PXnaansXopAS1yYevCLHwPi9O0
Jad7XaKrGM/eImFFWICKzz5TAwsS8wDBmPhU2yFx4SsQaFaLK1o7wKZ9BfuMuXW6oVs0iikNMF2a
pulgls3UICigAQCu1BtHwOKSj86opw+E2d+p1kGDZkRVUHGHGzrrqeULM+QcbIkQKD+t9L6BeIvp
pWyLVPx4yadT+lES6q9Ls0rVlizbdMZmxVJv0l0fThrW5EQ9cyjFHCCQkY0FbMDvfD1afarI1YTf
pQlMGjvRBLNE4fkwbJmNoQ5sNj6x1LBkPbz4IuvognUPFj1LDUTmNUQUUvgLEVg8TIWcb3IHrago
Zg9AFSdHu3j6bOIzSOeo8jSNHaDTxPKmtPeLhz5zon0+HSpDuRKK/qxm3X4FOZdxpYUyRO+S9f19
VaoXt4G3+bD+xi/nts24qq/S6WCs3jIBsx0EKMrKIyNJ3UJO87a+THuYSldaByhUbFozdPwGVg9A
Wmu7T60EL6gDUV7FzZ25dqvLkaKcDcrSzaoBQw50/qLlcSthoWJqHAJFQCfkc3e2Bg21rxjdBIi9
WxBktmC78tmxsi4pFhucTfLqV+ml7/Zxxh48EYmBjYlcVtD4XBt9L7JV2ilCka86lO/MWJEe2SrY
B4UDmGE2ZglsiAOo8V1xsBRO1W6EDHx04kbeTFl60PObp+gemHKmS5ffoyT4uPD3LllrP8s9Dbzw
DU76urzjSePFxdEuxbqgwvNSgfePgRJcheod2NmBrgV6F4wAyb+DFdC3rgM/z9JmACUhJ5IbmCho
sxYrc5l0kum5dITCFKkffWw7DvB0DfpCwmRb6Lr2M3Y8M6aapEfACBUkS9Z4F+f/6iKXB2MXz2G0
VKvWG38D90FSKvujmpmcBMDB2FskNphkVgku3cQkDToUKQZAzjqTsvirdY5vtTOR3KMC245CAZ9o
J4Za4cIZ6i7bXsopyYEND+ae2HBUJwB9+/WVI36TZgrvAKo/eW7b6cW+zIfB0yHQnlu9rUFgr9p4
VB4R67P+ox6GzS+3I+PBK+7GKpguW7qKzEs1LSWgkZ1rN1CeE4dv74tgyMpifWxebZF8Ufw3NYsi
NHGoOgE1oHPSztnziVrDFk121yTbkIU9ugJZBAJucz3QJ3oL/Gt03GA02PDirpbPFVAbhgh3pEuS
jBDkiVG4L/XKkrw2geD0bzmIppR/aDI8+FQDRDiXOmcDBWN4DRObc68hHvXa38ZC3ZhOUuvSN6Sz
xR8w0aDUigdxb9Wedx1+XgDlWwnFGLvcVWN/JAgRHOkM/GI7NJVloS2SjOx5JSVcmTTlyosgB8Pp
psl36IG3OZxF4LLxsC9TfLv5y7iMJfEg6y9LvAZr3pXs7SnnTRdn4fqbPyTTCGK2YRqcD5BtdSdn
/QZ30iwB532sDfBKOhmYLfj2Bied5/dZhXxNB+/IssGuD4Ghnv5kNEUQgHcA/6xtWADT7oHIwFro
iiYBPZh4s28S/dxky9butQ+qKlCrdfbxBYiGwNLxWGnnkx4p7m3AOt5ZS5wcwwmrr376uDOhEQLs
mrdBGuM6nWrskeiw9VgqMUAkeiXMS1ZYBT5MZeDRjdhFly2xwu4qqpcCUzHeys9Y/si6Wp9XkZrx
q0myNFjV2c7660H4hiWlcK9oEkjpxlPIPtKAlGWWoflz6oWQVeW1Z5ASU6EBkrp7YQHaYOetmcp2
kq+5Ekc9TCVN2++HxNcS5TonpVtsHnkE4WwfZiUH4xjQCOmuUTgLo6qMrxfgmN0C7B/Pq8taLj3h
K6RrXZMECRyLn7nugxwiY/ELOsXT8CHKHBWkLsIqHbPh+q+4T95YVYTkYHWXFWBKQNBy0mQjhN1K
5HyPA/u6VxTj3iUiXWgpDJwZ01lZWn8ZSDVAU3S0sLsuSdpXCK24mzK18vKsS07YB01sp8C2PcQo
NfyszcgbLxMCtFM/xs8+tSgKLhI0dM68Bx37dqSOliLEpfSyDvBv2OiNDuxavNvYV8+7xJIxBbNY
/ZxsJ0NUaZ46IYUeNDr7rvpqjT+zn7mMpSnRX6Le0sdsqxgwn9KSiI0RiuQzVtlnUzR8LBOeM/Qo
6ODcmAXxSVY+GUeozVbGje4Sm6TNriIWr0HttEzqiIsqAHPUhloq99ziEKv7KOs89byQn/YfInY7
eRBgqXV0ve58rH5aarLf+EyL/MwFiPgnMBdoDwf3mPl8v+x1gA2MeeUNr5ql1PHJuH2DtNlNYuRh
6nrZ3P08rB8ywwvLYEtarz8je/h37NctwTgFmiRPyKHkXuMxV1Q1/YIUxeT6Vm5XUEO8X+iiDPKf
7GN348vYRoVS8A+SvKUoEZ2cfiOAXV/qpshYidfbpGxvxK+8lq2FpzV3zYA+hSlJlSVQImqe5ZD0
fP/pOzdRKqyiN1VjNDk7NBB9TIcTMA/seHKPn55/HvVCuILUOmStk1Ns+7dl/WsSfkjUpMBRJ7JW
az1Dexj9nGmKZJDmtvpbQW+DMMSGCjJWeR14C6xj6PVKzNcFOLANnBBVE9dtvvvWv/y2kN69foSB
BBzY3Qz63tfi7gaMuI1Fs79Y/2h+lPvhj3Pc4YEtGOBSWYrW6ytr2KjnwfUGURoyHLF2ReghhkGU
iak/f7vs6aDB5O6Fr7ANr3tJfzD/5vf8fTdvph3/nBBIzm3tNoHiuZ+6tGeyX+IU/gsWAXhlorUR
AJFxpB1QHjWCrFS0dkAmOjLx8DNCOFEYXUZRuDQteMo+sT7GZjhNGaCQeDpOA5XF0JvhGbuI5a8V
LgLrFFYYHMoQbR8E+rNwdqYfuCwPzrYR2RhRSNl+BB4B2VHALHbeiojLO6L9Prko7yqOolpqli4P
0YzjQJwYa++tJH4Hu+n26+O9dEVlrg+IllQl0VcTlpQfcDDhODw9RPDvFQKOT5mqV0f4TwX50Wtu
PtC6Z5BX7AVnIi5oVKvBES/SHFKcllhBoLBeOog9YNhZ5Lw+tSCAcbNmRAGpb/6oG39tyyOcMj3T
gkfsmBDUFce26X0Q3WnQUpzer9iVSj1RyY+/bmhSapAfbrlB1euHgFroLbRgTs8k2IHmfaRUROc9
+MrBhVitB++2q06D4u9BIHrUmVcytbtiNopUidAy1SCnx6ZUiAJZx+WayU6CrruXktKAC9joS9pl
aUViB84ReJcVH1LqpcYoP/tgPfusmrIU6c9WHOEQlWDl2OJ1bsFi7Iij3i8gRiG+/DoxIsPdnuPi
xqBRbnKYdvh44J318rLS0MTzxTd+23VZe3m7gEj634Gsw9EQ1Gl9iAuIqSj1vtWw6dZ8TJlODOQv
rvT3sJCcTK3VOUiXI8sHi6igKT91kSvoGXgDZ2rzDbDoMdQiUgPkWqVC0R06yBx7NLCf6UUUPpSJ
zwvDN7CoNoWkOZ8tNo/lSFCuOgn2qsGbBwFovZnxexXeTePqIrnoYsQyGLUccKg+1VsDDioW/2EY
08SdeKxDOkZxCss/ETAxQ6iSC56YC3iCBrsM1lwozStPMxofCXVjLjc7MwqZjlxaqnObfiEwL0wW
/3PjP4sR2V1C9Il/4Tg8OSlv6iocFuPHkPB5nbkKIhjuS6HQrer0f+VmjqvyvA/nnv0LQUqRmpkq
Wp+1sHOv1SwjJ3FNZXGCjVh4kQtUtKDsxQ8+htLLk6bkUfOekL5g6FX+d4GbBEK8baCiKWff39bc
3OzVJuLOC9qtgjIP8+6MQwRBCVcJgZ/QA9A++oDbJtsvVuZEKE8EvLLzBidJ/UqCgwrZpdCVGM6H
ymRWObpo+EOkwFlwqhNT+JLZLfDqEjHE3CAkro1Z94uRB9ELrvzA9md9cdlZ727PMYpEq2lPzGvd
gAyT9xMbi889WS8vYhNPX74t5Mmw41G2EhVGK8aKA7nvzMrOgEcj8Ij412dWK1PXYfk2m4D8TsEO
s/pP/TSEyLTPlWuo9fq2Xnfo6IUi8J4YQVVoSDAQOqCzt3XYPkGzUgE749KPaLv4mAOP1qVO1hnl
SQd+6HwN8Yxb/FhFxelGnnFTPJxfm0Qp78u/4KqYGWiWvGIHXF7/Z0Oa1IaepvtbYnxe+xaOLhrI
NyX6snZYhwBKP9efNcPYfVP1gNCzK6FEqYl/F95Euc7NQI9TauSih1SFBiP4K3oYLinyweQQw5Dd
jL39M86wqMfU9vJCyqp7BqpJPCNaB78qrDTbRGXtMpdFKabgFCY/1zRMoORFP+FE/Lq971eoavTv
oTxCjf6zNeYAeVLZP70adFoep3r8WBGugKUEihmVN7Y4rWdbUCh0aM60XIt/AeBLWnauXAoagb9H
zKKbPEc90Ul7XmOvyT1OwyYLly1Svo9EGl2GmKP7aWMSFrG1LAz+jGMaRoz3TwbbrKM9LRSSLd0q
YBZOB98CmXCeeUZ5MdvEM8fYt3WP9dnm0BLI83k2vQEaOilw12gfLxQ1TtAUm6pI/MQnnfSIehYC
E6YO12Xr3tovHKHDpj6V8S+fpHA3VBnC+g83Jxv7ymLw1l2OxqTcgMNoR5Uyy/n7hn9qQVwvQnJC
iUzxrtiBT9kci/iatioIdt1EEwXIPE4LremmzMiCDJ0CwuYnEIjSoRZ8PlEg7iaJXj8gJJSlGfzf
HAdt0W5U+b6tbHHU/r+gfMZOcFHxPMCectVrwnDl7vwYe+VmdygWylz0wwJ+H6916UxdQIXwei6g
mqi6BRzdCE1AGLNt7isBeWhGKJI+AJeQNdwVVnyFVFSDTxx7LnGFwolVEOOF/uWiBgUx8Y7GRHVL
td8+n7bczwXp/rGui/4L8CIK1hQMW4mGgAWOooPv8gJ+B/ds6J4/1uESdYu9cRJGzxu2XMjA/WKa
t9y7U/u1Jm1uBZf0C49nik0243G+YijC14dJDuySqZqGF/5O/ZDozI4L1K9lomBAtuF1a1VpKXZW
XEMlHCkFyuHDEXxqRJMAHoq9D3zG2RCgUw7ZQkf5tNI3fniA8VXYx1os/wgh606yrUO3jBmHjUm+
T1AYXFKBzgbHjOk82nG4HpwXTmyHRX4RnkiLRkyf4Ye2WU0oFkT5oyAgpw1hPJgBLV4sfb324Urb
rT5wdkBxaG8rmGIvqASJ4nxUWlcQOHPjWA4+doun8ca473VN8hbZZx4pQMhGEjv278EaPk+kcWhc
IpvFclR611lm3Y9m30fmy0E+HNFiJeb2LwKSVtXLtdFXPhN+EZ1qSFKYyGG1uOyCZ1+Bpi0UczqX
hyEw9hl+NWTkNfH5fn6eLU0+B98vAr402oFPfyPum7id8+KJPvIPD8oPr2x2+KpOTD+QjvHE4AT+
z4Tk400JKpMrh9Bv/XAtW8JqchhdJVAuCDCeljTY4bfCR/7AgwBY+UdLJhqLlClhIygzH5H4ykjE
YK7KXmycHHD8A0nB+ItLuXWZxGefGmDVylXCa8Wwgl4HFwHh1Lw0wSJXUQv6EJNTrBKi0WSy54A/
LxGLiq5WsvKv1xvkOJR1EKieYMyI201Dh88qoxJk0bI+jIyqPTkkg1If/o3wJ4WDOdli7ubzfFIr
Vz0XU+xluTTH8BPxMaYwLjZdEHwklSvazuUCk7aZ0vNFOq8ZoYFDVJp0mSe2uXvtX93gZ2Tp+X2I
mGiNvSkJ1Cdthaz5IUteuxEuUlXAhZwn+ickencQAY/JIjxqezWQuDK12o/FujBE5g2PTIcBOqzJ
6sP9FIUcFG+tJ7taI4ZjPoaPBKgkaO6xw4KF1d/vazaM6VQpffFpxmFrfYdAZeeQm34Vf4KkgoL2
aQz/qD2nCRJI5mmFh0vyzLDBvF5FaaHWZpKa6WOcPTpFSyerEX/FrOaQosRFi4F26HhKX9mHJLss
8GS1a3aciCF1OsdeGsjqzpVO3nLjbHTZLa3XAgQT28d5Ws4TDKmK+cS0i1lsMg0SZ04ml0A1KPEw
TWfQsPxkb+pNOYAo4pQq8j4XynlkT6Bzj7CiYBjeSkMgStZh8MVN4J8yfcA5v0z5bSXl+nvI/P83
kzFzrbxRYWX1xhEVieNJTprRkanCIYKHH9iic9j76zhPFgZoQ49eaD6mdxsaCw/XcM7F16M4KQPJ
5iUoItBU39mCCEOGp/p+KqIG+xauShPJYRV7oTAqU734WywQyP1R9iQ7pEMenfv8PduQX4Q/7p+k
vMhny07Rg8T5YyzaLegFaaL8ML4Y/rmYaATdORlQX/1GM0Iw7/lpKqkcprIG4x+HozQQCAtkf75A
3uMtvmbC84UL+X1NRupTW8TtVc7L70E8eB9SzmvA8XDGYOC1oBDiDhiwY13mlCUQW8Cna+f6OYov
i3zUiGMwXz5QlMNj7tI7Z2ILzLfHSgDYKoxqzXXJm/cavfdsgxhb2IXg0f6zOpgIWHvp5EIJuuvC
UNQlGTL6mAW2jjq8akGNmuFk/wA/vRUAkx5NUXG9iDSbVCxmI/iSyz0D/KjRttEmO2MCoPXHR7PI
BaDMQerA0TJz4DUDEhhaPGnkDRZA8mXjUmrsnl8/nyHSft37RuFWmejytqItxekVkr7hYPl0IRsM
Ki1ArgENFB8+jvJeZa4254VL3vr7r71R+Qo5oAmZzwlcuY4GQI63T7z3J57Fw4fRt/iapwoF1/oH
KINyJri/NyvrrVw53cv2wjQdBg0M1R2q6kVWIIkO2xPqSgsZChA6+RkBvAl2oyFxsKPlpWkrHSW3
EpOSQ1SqJ0Ecp/f8EfwaK2HuZ8wm7gTvw+4KyFn30pDWyda+XnDqblRDAnuJIjR3Xng4+AxB6KON
eoepgk32cygCKwe6X/MPHNBIq5NsE0la/laNmhpL+rAofgFiY9CzjwR9ewr0And1xbR6w7IxyBfQ
BhlQ+YKM6/DkzZKtk7u2kyGa3G5QEj+pWoEy01xhfTrqtwKM4De7wos+5UI6/w0x0ClBP3Gknu7I
Bt/VfjAJC8NnW5GkUC28/5+F3VAa6Q6e2rKSIaycDEHs0dAcN4jfwgdvdvHiIX8mM4yf/2KR4one
i6qhtQ8BgrEvAwK7AxqT21Z0cpXCflWha4NOxjSLQVuklBLi9h0IC6H5R/p7ifKV4vdKZTrCKfTr
/jpqUWNwHY1uJP7JOQjRmCId5HLtzrgW2uLPu5y5Tw4zHEAPt6wQQcTgYjn0SNU9I69oXetcyZfp
v4vK2Vl9ybgpFCWTAJg2rx9wKOVeNVH1mSNjDuAK7TBKzm4nef+9K4sUP4PIO+N8nZHKyxVG+sOf
c9NmBTPo9zDb/HbvSawhHycEfJhi2nKLqCCNioCitA8eEJoQD2w8y9L/j+cvJZPLi+sd2CiycRq2
WJkns6VeFArwCBmk2VwQf3HE4JW23cZ7HTIubTwBAVBzZfplABDPxdsW1gZLg/VnPVWX9Gblct/T
0grRXAIdkgxbVwiqDt/Wyy0sjWRz477z0zIwkBcLqu3Jjfr/E7BKM1O4Ya4ZX/C1cXIWMSwESMcT
+fm6C+KukguxI3suGPAS4emHfLrUrwUeXTwxCye2FfDYYggXkDz96Q5wJPooGB1ZuHjsgxT/1nqu
IugpVODjzNEVVqn++2Njqm9CYJCMktYY3FC34tBEd0XO/FVmNCMTAc98uQDO/7mQqCPmoXMmZ6YL
Y1TLuxabng5ozNgqzdJ/tSerdjvdiap0x+oMuBxYyU23F8wwNEA+dBa/dkoqjy4Ih6wJSyWso8jl
2qzVQ5pT2oKD6MX0FyY6wspw5L3hd+HY8bSYrxOM2aiaPRGoNdUypz+uor0RSSVcPkW4GqXiWwl1
mjwD2XOUoADA7LFVS/cp6r2ZQPOGbOeJ4lwxpCoWPGSBM3+SbVVHshvoZl5eEj45I/9U4Nfr+P7n
/QsjePAwMTX9jrDsLj0xdligQYWxvnVj/rfCViGIH51BTmtcWRFZRcwPRWsyeBdOVN5DTtgPCYxb
8IM3xHyI6xkWM7AVobLPM5w1PooHbgu10ifvDNVP7xFYgdOmkTF2mi6MwH0gXzJnBeBVYiXOuZkz
A+obnWEdEJlN0t/HfStcTqnEd8dCp3X+Btv5eahWthxYxk6eDovoQb/xi3IBt1hBMT9+J82B5Tqo
hRTYWGDmd00iYAFVvH+EPdfurvy0gZQsI98Ubz7CQQxces25cxnwgyU7mr/AcvOHXksXdZu8dVyL
79SGz0HaRjKO4M5BL/IZ6vXgO1cm4g3DIlAln0NbIhJ7Zkn9sBcqSITPoV4gK+7dJAxNb1g6WDBs
JzglBMCoivo64/ebZBDAyrPNfahudvkn0E8h8xEzjuww32lH9EcCq5IplVKMFCvkGQxAE5wxoc3A
ksayK2DbU9tijWQCchkxOzC+xr//zayc0Q5Y5RQZ0ewqYGWbjx+sxngT3MFTX2CBAAbctWPdSykq
8hTUjpo8YdRTGPGYcZVPxry4+A59p+iUdEqzMguQ6WUH72S6PIzN3oFCWN97bxCHZaG+ogvFePL3
jrGHQN6MI6yz7jJHBYeeW18ClJR6qStcuiVFnWyyJj2HYkARouJgNWRDePQb91+01esPsEooMTpV
BsyVLptcYR0Fl8ZviSxs8h2guJJ9V35Z+lCrHmBzJ/J/qCt61aJF+qul20LNuURY9MfE2sKjRLrh
8j7tOktN9JzEDQkCJ4sj+t1GTcdFpGmILp8lsj16m2C87p5vVW+jcbEz9Hd/HV3W6pIZuulks7VC
3xr6hxFTi/kNXoLEMX9T33BgTn8GyXmb0gn0cs0P7de9skz49b1b4kBXcNMLl9hIegzTrfDmU/Nd
bwHAjRGGChizxWJx9SZvWel9PZkn2bDqw+Og5Seizbm2ElwIKKt3QZJFd7UfrONXRaziBfXMiL6O
8iEs1Z9aWVm9zrz3CWaMX3eb8TYYzYoZeJXAFYmRhAMSeOZ+RZjGo1PNZDdXeX8Wz7RnI5ONxnMd
deWQ8SwcTfMtkVPOkpGbbUoOvpnbkQ2u54gy3OGdEoqnlxQF4EKh1vJKJGnSSymYY0duhF6ZFYZ0
o30OvyhKDQiVyOmvh9669j1iTbQhB9pv3siWDkatXIsH5dZ+WetlTBg6nmzL5UKf3bGvjYtEX8L/
UL8mE9wET6xZxJG3nsLnIxYfq8d9aCufwdRUp0V2xGvsRMuIZ3Rr0uRg3zR2T1g6nEQr2V4DOphH
KGfHztmwmuczPyGqEfFx0BOt18QBHeY8TcgC4zR46zk1jDMvMGbQr3vnr3Hk2G1c1SFhYBh/aoSO
ViS+04xkn/UDPG4TO0FamdzSjHexN7A9kQLc+Y3rORaXNgUKG25Luys3JqqCURnxazswAY7TCtaZ
p5c6hTcUGQkDr/j/j90bHtuS2Yy5RZcGDa7Szfpij5E1kdf8cF9bbJifH58BuE3WZry+FPnLi1Xx
XXPbBiC7EZVe1OjAsSylLi7PUa7i9B+bzIWPm+Kr68eKVYY55UlQTKc/ghRu/gXLhP29L18fcFB2
XG3Iqp8NYh/ET5sjQm0YbJ9YTtZZeg8QQiw82WCnw4vCfRYL7fhlis+JXkOo4WfzobKuPdyKvbVO
8/MRM5dKQJUpXHRONkuOdd4db36XIQqKUzKaMMh7VkOJ9E/R46QtWas3qqKBzhfd25ACnoDhlmmL
qqhsiCrpdLYSPYCYQ5lJj6tM8vPjQt2V0SzOFQU6G/87ljQuRFB24K8JlBZU5AA/fsJzoLtAY5OU
TJWU9HLw7I1bQvsYTa03w1wxH5d0tgE2xeyoyqJgZqQZrmNqQwETJfq8xC2sm5ovi9zf60n8UGUH
T0SNW+j3SLxeQgxVI+9FCMFhr+oM8XQ6vyywBQYHic21zC27HhvutDYkF8zTwk5yQikj6Pq1BPeE
WOSbqH/BwTQ/Mucm/4I/UIzkv5UAsLIZsU3dTpyAYApYHQaDp3oIua8Qh4su2jMgAu3NioLOgNWb
5km4q572tUGYTuD02HVJNksGnfuvedVAe1Li+BlqG6mNxy2sEtaQZDaz2Mg9+9eWVFqc48Xp54/u
VhV20hhY/mZ5txUTWnf+/HAr7jbVwPum7IjpBSEBtUDcVFd/hazgGRGFujyO2ZjxvE4zKihVcEAm
1b9ldmBNxeUtmc0LOdvoKguivUuYldjXGqjbfcYQqd1WQwO5oGs+ERZoz64H85FVREugSQ5WLgbg
Uuj1pvU30BhekA1wY/dGbaX4muMTJLwR9oH3Rz/urEsaXQAiWLOAsLH7Vx4mw8HZagXezCDSb5d1
L0L9sd3H2iXWqM7GrS0bgaGNSPt6yjRuiF9KEDzFAHevxbCxHCMWko2Do7BV1fzj6watqFWwJW0n
H7EjeYtjVUG+sDhdNiJmVGZhxmoZ3Nk77/blDByXLs+VfOggB89jJ6e8kXRjRlc88oxvH8yURQea
bW+sChjPQ2cr6nSTWjgkVLvo0V+lXj0vDPWJo1DgWF2YuQZydCnmTRHg4ftLeUEwLuxrFueLrXSi
eQbiG5F/Hdy5K9LIYlkjs8efVTvOGGmgy7F4tNuvNuhG1ez5vuUR9/F1Y7JcgrU4Fajl9a54qxd5
VJ84yrZTbyzBcSiQE7GjvOJlfXmaaOCDYpJ6hCEOmQ1EZIqGgAd9bk0U7LTSpg/1ChS1G5eRCgbH
xORVV6/7DJk1eOFE4lr/L0Ls4y3H99IlxvfJCx71T/XBdmG9u/Q9Q2UANsO9HxX3Fg1duV+ei1/R
WXFxUU8pGz7cUQEUsCK0AWgout+2LVrbwIiwENOESTJqIG4UBl4cyzTBh49dVPYOM/emXhaelDmO
fT7wxomJb09yRFxu9q1kzXU3hhqLAWBlaVuV9TiQkpqCffx/32est69h+GcUjyLvpT7xVrGVwnH0
84rnhWudCn67y4QfIa24MKiR/QOEJykpAXImSzCsNtnfayKuon+RIJ8yg0JwxxBkOzkxJFEl0PKH
i/lRxpngqmpk+KrDF0LNf3pOpoDikrD0qNm9Q0q84Wg9OOK+9uZd9PplcuzQvUdhemM4eC7HN0r+
SIRk4HcyKm42C80nhdaGd8ArjVljeKwpSDJs8zuKpOiOr3Q8XLOnbDiG2+VTcIW0TfQF/yBhe+xU
Ca3/1UdscYp8bmShwe0EuA8aiSIjboIupitukoWFV/QftU6lteG6CpMxxoRMJNAnqHrZ7Weka0Vv
HYefC1AyfAV4kLJn7KBP601MtB+2qULyrM5KrpJJxm54qJSLVNoqJ2C485aS02aAoTjHyIKyLJc2
NmDwZSAl+1Uh5W6Vmvnz9eGfuwqFgTOnucGj86ESNvIuXoKdNZWLfOqA9DcjS0TPiQ6w9mp1zrnF
t4Ot5qtcJSHIRFw3Bhl0pQsqh8Fm5/E1RBYZhB+rKaYbLJ0eXXwQNv4AOSx8Ux0SlJYTtJ+vVici
99cThSn+TS5EoLuVY2OZ0iPtuGlmFE4EqYlSU+fnMWmXBkPRgg3p7htouSnannmCrTdjUju66GNj
cT3YDeV4I/ZuZuu8E12roWmXjv5Xzaj0gV2dpCwzzvvS08ApXxyg7b5t+yRFNUmLPd6mJz6Yz9F3
ZvlumhzFo6lurFuxTXya3SKo1eW6+JlndZtGjK2RGmIE5CTfSMt6fhTkbZ0pVA5m2uZTnCe6HRUN
Dq9EarCLU78o7CJafcwlAxdd0e6N2XJBEnUjnRZ0SelvZAl29+MBgogfKksfMxnjE5rbNoXAq4nn
PlPeeGHUZQL1qBa0Fmy0mXLHqQqtBWHqIhcLaUwNh3E4L3X1kkqSdzETjLMdwSblX0HeOVdv7Nc1
OQ7f5bNx9jN8qwmQYWvx17NSR/hwdR2nyhqMPqIMzuAOShRD1MXqxyg0+hlMTdFl5jikJpuYam6t
X2xsZKGkUWIbJ5KnFFjg2QCidFVlf1lX7xraFQqOA76Ib/c2xocLAYsMvfSa9kSPsLBJ8igmYRqO
HMPjO1dBAHvKrUn45thX91z5dMwBrl+V2v+ZT2Gr3lHK+gcxM/6F78Lsm+sT5Vi9g5YZ6UpnY90e
aE8tNTFkL40u/O4Q5SXTMrAPsiMRcRPrcOgWbqNCxkgPjxul5YA1ak2uRlg8YNmzQCC9kJMcCslP
qolGYArCNRiB79P9LLOtzVVEPwTnkCCKr8j0BZpnNih4LVHqdFqkWGGQZgWfPhWQrm59c4W8D29H
MF4xIu1nrXNq7A8ie+KYxor2uIF2mQrv/Y4xpC07tGVNUVNcY0RBTmPF6RbrXrCJvbvWntYHAXkK
XeuDC16CPHqRHhJTUZC1U99giO5v3Vg0o8ZIVHadPGNABjSklyQvem490CpxLq3cMOXztqWYpEco
5exjXzj+Rsg5T9xla90oYI30BqhWUaaoxfDyDBTclaGJ5o1sZp30koYKon7q4Mn0I+Oa5gRmTZwT
rGn94ucDqOGd44xhz2+iC6GLCC/90F7IxnanZuBtNMktedtBCyg7tyxzq4VsdBVBwLaBwjpgiAqn
aE0VRP0c+uXuAsA1b7MkKIosJ/KjMyW/ivl8yWQiS12QPIT+s/b6XBMAqhZlqDX6rhc2ai3G0KJP
e1vMFbC+xAxiCeqTzBxWVs4KEJwS/2SyyAqUhoOaeSWAqz1gFIej5GqPB4lY2vpaklTIHREqYruy
NslvfvPED3XynkgjWll146nHC1JP/3iCI+c6P1AWQgwLLmJAgXr1OZ4oawVHJouRu31nhfhwdQM4
MhquXoW7suHZkONRiEIfmYSPmf4IwmYWaKZ0mZ6a+U342VgFE0wpc01Q45axg/Vye1aLD/6RgCI+
C8SRPWjDeLNh4uF5delOcWsTzuIS19NkAWzCOAddMTo8NDSmW+7MPpdkKg/FLCKlSYIEHVuhcweQ
K8q2LaXUDG/Y1lG1JCeolhOOhKzQngJP1+svjaM20KmCV3RzJwoOoKEbrVtr8f6om1NA9kff+UA+
EGmA5/evOU7NDTVCzs1OW0STUOaMdNTQi85W3ieU6lVpzvpJGIC5mDhGym00EfWSANoFtpamS86r
6VDX1sWIyLYeRxYlloZEk8WkOUTnYm1j0/1RCngwV9Ez3i6P30Af0eCMEFEh6QDyI37GO4LCTPOj
2v3+SaqITnsbn9AhQzsSofi87CHFx0GXNluvZ0X2WolTQu48MS+BWLEY2/MhhFRh4xm0KLbIsoas
M6KuerpUKE3Pe3Xzpe3A7izlv0586IKE9mzhjd68wQnyU/icCrCQtXhvh9RhA7bEZ3uyg1tqTAVB
a3jO1NbtSx9u2k9OqFgpMYAE8e1gqN3ifm0tSZTwmDXvkVmBIco5RntAkLP9V0OEwFOK+sia1PUs
HVmSuKWuj3i3+76SBA1yUDEKSkWuxLwNpTirBqoXfCEmFF2lVw6Y45xXUDHvxKzqVQdL9IshXWy7
V0aOcUd4tCpR+RjZsUpcnd/OTs6ZhIhF70XWVY8wLByx+ny3GgcAA1SGbzyVH9MK+1eBY8VnZdc9
mDphbaMGb96nuxOEC95/YL6RHQeDJDsCzFvGdxo4X5AjpG2HhoUVPChT7oxzzeWjS412oY+aEpiq
o8saKe8OsjvKVSA/D81DRJ3p77DnC1mqMoJyXl4lBoMk7kUCzgE/tvTYQNZhXvtfsK6ROUW1XOCA
x5z2O2eiuF9O2bl2JoLoEAwM6YY38GD+UNiCzYab7Runoi/pAXLUyD0wiEls5wVh+Oc8z3M2/uyF
JWeda8nqt9IW1ZxLEapkVX0JOBedWelsJBh1vDkayaTgjpD0c2wwaGJ2vpptkqKtjxxvAPQ7/cSM
aojarQ/FOylurFaN4I0d7aoXnqb64dAL/yAX3k18BQMUQ8hOjXnXsvguHSWrZJ57NAD4KyIfTwYU
osjbSOJGet0p8wapM0MRFa6kjGJCHYWaPHRycdiQZT7hljnPom2IUd6om7GTcCwW2QCjNoLt0FHv
sOJbkcDdRNvlqWL6L99NPcx2OMjiWzxlKy1T3eHnIvvwo7zsNUgAfb+STqu+Bd3KMQHYrnJKBseO
WnPM6cFc2US/mVG70dtHmJTtUdUwAuBx0/Nzrv5lX9irTRe9bvKmt3jd0zfWO2wL0RTYR8IoyjxW
MgOGHVTFIYngjr4uBrbVgMx7GydBB8GljSlAemS76DUdQ02LfAVbgQiG068T3/Kb6PDqLIoPJgeX
UYdc7QHHhNSllJKT4ffqjCelEG/3KQbXRSh5DCuDPr1ckvqK0qRjFN18aG0y9K/IocKYqRa61pEg
x/YqTvRzUVqQ6V6rUsEuu/kP08ADeEpgckktYqoHKPOwIWFUY2t/r/svmPfxjRsEtXev6H+5HL9r
TPD2uL4nkI2LGAZ9yweLB6F+irWsCJXZrilAzEJ5hZgbqhCi49kJw4qzFtO1SMtyWb4L9+cBmxdx
laeZ/Rdo9lvY1jbK4G8B/Hm9Ye8Pqz87A7CIVuEZvTE0m4Rptp+dgBkvd5x7sq4PjxAj6Rh4HHfx
J+3FmMJXgNlaK8HuDqO8AdKjLq8RcuQ+S/6ajs8ePC8P3O298fP0QOxb9gOSwGExI7YjyIGTBrf5
tgPgfP+wwpTzKhQFo4uqgm+3zB3zh3Rxo1wSyStRrnXUzZIeGk2kYRk38W0AtYbwOAV9eqMktYI8
KtJ7cg/UIXzpkAodvH/JRB4ak558xvKNtbnEDlV9xEpA7LzdjySC3nW37E/n3QaNtbEPx7TWp4QD
pXX9SUjG5ywxmQkDwL2ZIXrnadABwxRAs6zWrQOWlUMmbpAskZ9iQgwBTnwr6zktu7X/PFk1dTZu
jjOM11XKZ2JNLJSxp6sINuF72hS+GYpF8iVTtmrGsoqsNjEaJuIHUvbxMpwEqasL5DZU8pULXOLa
8rmWP1X/KGZIBDhhU7wUoSGx7I64ctd8kBYhWjAQmErnt2RV0MYRVhtMNpc9Vljc72YgmGfrEp4G
G16QzXhfAWwsq4SUt4ZkuRRNymdIK+ZhnHz+8BiTubZY0GpGxiLoubs+fgUBMT7grf3ROGHxsxPP
gTdchxUZPELLyE2jnpplCc+Qgc1RYWX5cSXHdZPXdafI1y7UaAXVHx99Stk9B62EFnsTKZ0HvSF3
PtE67XTSk6V9Hh0XD+n2cgWuNs0lA+kueam8bI4r6PFVn53un0jm/+VaMQCqVs8O/xiKDVXF2tPj
popEaEtINYlJWhKVKyIsnKU4Z4T4iuitqPYMcx3ERHZ1T/cSsngT26Sc36znvH0Hkd1XKo1nMZZ4
HXTXjFBsPANrJGSDSu5AUGgVYl4UDFKySMBgYYlNJF5Xy3hXZHbADUivCyCvIfG2HPt0qXhZ0hZO
hzzGuj7haJq7c6+B8weyX74WUTNteHTX4Qx/VbGE2ISVTXvKK9t2xUeFg8WcHi02Abg89pGOa55O
MKKtH1wfHO2pEJVNfby1E00XaepVay+vFKvMsIEmkg/F6JmqpALsElM65TuY7dhFRwxuiFZvPYEW
hcxMQjgY6lF7VdPv009/58krm8RGF+5EVWj5IbSG/zvilnbBXLhnwrhYahntSyAm3oP7kHsGd86C
vO8zrHO015C+QI1mgW7FT35DIQ7fiybzKB2od9WXhV+4HU1b/Te/anfBs2NqxyTSeHKmvxkLLAKb
7GUUx94vuBZh1w2pZQiMAPDQXIJn7+yC3LlSpujKCJwTzh3p2jfkwNxO1/eMJz5qyHrmzzwwLqeJ
FS6nGRi2RglnoKayguxJeJy83R+031wMTb4ZBYHhNe1x+VI6z5u5L3OrmAtvJWjYzU9/taWLlPfN
/HRqJUrW5iA13o45TtQgXO9ZS+fVB7pTo4rXREI2F7zy5iXGO1Mp5PJDCmasnPXuZ4EvlHkEq6CK
YKqeZvd2ENSA/9BbrALMyvA/B0/6pf0X+fG9p9/eUhKm6CjpFucdLy0rcCzXrQe3gj1vOt5he4fm
pKbr308qj6G37bC6Hx1nekUhVcJxSVZM3ujKKwd61OmNvMr9ptruR99WOi4K2mwOD3i6Cpj6MrZK
EvoVlcIOcRcoyD9neUu34j6uklngLPY2glJMmq1QbWpuiQayxFC5EUKsYuApiBq1mwKbqLTXep5+
B++nn1dWfq4J5EKJOtcaFucfJ+Zd1LRmKJ9N82CTo5hXk+mJ5dHiAdjtqH/Te8xlllflTXZsApqk
DC/A9VaJgAdqrbNoHMRFUUEkpEqKWvgCQ+l0Ds5seofJvPGSzKIJ9NXzFhkB5RVoX1bQkQeIYC9z
jZg8vlqfZRfsrTgx9HYsAxypvVV2qKgnZ5lV1XWB7TS/A7x+jbnhGt4HeHqZ2mHHaUaVjo8rNhNE
z0vnMNiXz6XJDYoP2J1yLVci4eoOeB63vAOeZ4geVYhwTlTYrxzeCHFsN/pHi/CYL6JSe92U1mD2
vHcUm728VsyAPoECPzZiIJax2sbVn33pBmtbCJ20OhOUd08W9ZAveQ/p87zdUyEcOsJRoxHjhlOQ
UnBBmEDUqvOZVTsI/rybNE7DZ0I1W08TVkstH+I7S5VgYdIFBn0cqZrdkohp1R0zi+H0fKcWgI6Q
dKOYArPZW472MBfH1aprzP46OR0dgj4abINPJVlf8HVRHbhp/e5+iQZ6uzohAIdG0WXH1qMxQSQu
522cnonPwY+uNQaDVRlmUBC3PU4Bk+kw1dwFctdFTglh4BhYtlVT8ppOMYVruNtRBIy8c75rJ/Sl
sg9nS2AZvJXX+5nIp3EmABb84lmhTcaFxNp0ZwPz801ub6wjTv4Swqu4Udwv2bOLLvGhT/B3C8DL
nj+Erd60XrzSfSw3C5w6jMSRzElEnCOMS3F9QQTp1vwK1yphwdmQb3RS5L5Immh6y2j3di+gof1b
2NcylTd583dbqBYWKp7jABge0hxxw2xKqUTCtNWbMYJB80u3qFkn8LYpk7UiZdqgJrPXACGgfMNV
uzXYYwJJb3sd1FAao+IqWxXbJ5RwPHIkCWh6cEC/M062rR31AWkwAGD3ftWNPcb6NuSj2rgBF5/o
RBeHkEJEIirjJ18Mw7m24MPIbwAz3Pz+5GUGJAfyVb5GJ8lu0YJXlvdWOuJrvwLPbZuKeOn5FgIY
mMJvkzTvZ247IxG9xVA7EB+FrrSr4Idx+8FpF69PIEISgUoJSLHuQOfIPqH/u+AFWdVclH5RWIHM
0YQpCjmMXQdRj9J1bGpFXlj8s3fLE1VEnpDqal7gnCA1KFF+uU5vdJ7ApCxhhAYUMm0BsWEs3BJT
iTfcaHNsW45oU9Ibe2P16JdHHBUjA9tyQ8uuvW6YRuGRdLYmO+ObG6tvdTyu/BbycuSHEC2TIaZB
M3Wummsa+Ujj9mI4RCEiWVTIRUae9X+6oR7oSsqcTa2sX0nQaXdI7s2ZxNzhMw5VfKpj89m+5Lwd
mfe5+c6hEDr8BPAlKu3MF+92KIrXWQOyj/md37+cvRixiPtrZIO3NJyqWDfzMB5jwOzz44fiWUoi
YNm3g6GGgwQhc5jL9AfN0CHWbrCnq4t92gxDPOGBWs2HhGZTFy4xntoyxUK/Z0YjIwdYu8eJkh3E
nNGK8Otv5UiULCkiFPVoxOOsRHfQxT5D/m2XSi5BA8W2dCEwKkY15TCHE6eU4+ZSgHZLOBXPC/cP
7rPuDrpKCfzchranznvzuk3FNPNeaFoLV18jAVxEc+08IDmybqo51TdnVNNNY7yX4taB5V7I2qXl
sAPb4ct7sxCm2qZQM5wpVTghDi+MTjIfWIaks31zRf/uXoRs3NtkL1HdaDV7+T/BhhZaN6WS3Kqg
VqC+Szjr2YCKuu54wsO2IbXQnFaIeXw7n1Vv1DC8EGB1UnYGXNRzTaccf2eF104O1hpamUfiCDjQ
8ekEqD5OPA6lBnV5GJufCHDAilJyDY+BgS6UhRFuv/sPZiWoTwscWAd+18T6pEf2si1nKV6fcFvj
BhoLkLqdv1W2oGEFPw8QCWUns+MNWnR1GRhuysxU06+wwpPmkPrIDtlp8FvjGek18HQ+udlXNuZM
S8Jxg24sKu6Ee7dKTPO9TWyie0P3cuilOu69yAA5ytXgFrarwKpNL97MpVaqv6xpd6HYWSAbMHd9
WkelBwkxPJJQBGr96WkifqCkvBk6Am5YLyl7zWcjYQFat4OYuRIA87JYvNUKpFQvJ68f5MhWjAg9
oK690DFgszeqvXoIBY4oBNZTCrlS2koybLK5yjO65xpB95j1iYYkU7AeQv5C7Ck64RQWLC6JOuxY
Yz2AFh9Ic5+GS3cj0aMmJrib9aqfYJr6+9cfJ2/SrRXxV0BsdLEegNjwSic77gbmynHANq82a/7e
05Ib6hrvqZVSL9odyUfOkwM8BNp3kAl7N/WQ+nh48L5Cg8G91ymgTvIiJw12MP0cTP8tgbzwyBEz
WrRi5MJEW/FixBJr5J5aQQGA/qiWJ+kafKuKJA3iPeZdfSLDtBbjvx7lAlvbyNfNDUVwWb31W40E
+G6EwPhVgsJ3qSc30kAmBWO03yA8PCTnyNc1gq0lXZO7TlnX0zjQQKpGPGbBEHLywb4c1LcZ2oEK
w+wj7wUxHK7B/6JKR7WO9ANTwn3+G3jUQ9ccB5Bed70V63McFlJayS4FvqZvDdv54ye379B0qePT
3ju99P7uEpgwKjsS1CGnR3w8nykifQEN/Q8cHk0RhhzhVY0PHIRrGRAQkjP5hS5NpKOeiLCThAqM
9jIbUSgx1JqYENXL2x8hi88YQqdPq9cSswOlI5PljFJixc7bvXgyzWFg+tCzB4Dp/2vafL3rtfZK
lZBQHC/QJShEri9QRB/5zg48tYXxi2icjjkNoEliY5HSYlhrwBU1ynEGhykPw6EGUTTeCQurwNHk
i6K02Fj90HkKR3XA9G2D3Uf+/lWCEJItwCx5zboAX8/rau53i2yryFVQE5vIbaFxSWBA1Eowtqno
G5q0QwqONHaZ17WaMjHBa6JqA3KPYG2Jo3xqRWHEU/S+OBIC2uQTaKHz38w43gBR5KUyyKSziY5T
TAXGDOoMOfhigNm34XvGNhlm9eMF2cQkhV4pBc7lnfCNIMFni/m+5ks+52Jd/Si9bBYUu7r3QmpZ
1UgqV1MAcPOy1u2af6O7CYvdxlOWEN3odcQlVNTlboqzoFSw7laT5FGlWd/D07BQRCRwkDptbVm8
UFy9tH6PB86TANKSn+szBYye34t3bTccUFknQ1wEiKSym1TN5Bbb9bz+9L0mq7HmgKhMEEnN9Kxn
KwCZwzgK4QxKS33gIOmT/IvQilqiWERbfsv3981FmErOAXuPGvaHvWYoKdY7h1ev9547W0oJQbBy
kdZ8sUnK3PVmzbqkzfg1JzATF/BhWgcKlB0GF9s29ECskoYZahAbGYO1CuxGnbZxBL56B3ln5igk
O2G1lE5/OMPSNHd8uYylEVdOCFA1cPy2ogoMmMCguADDf6A1j+FYPg8y+AIBIIcqflMgD91jIbje
Q0TkRqhL2vySfBaq4FdORrZECPadEn0EJfwkzfqVKS+UKWoJCy7n2VVAZ1tj/Ah+TU0pAfuO6B4D
XgRjmq0q/bDTn5AFejp76NwRAjuFXky7Byc2xuWZHm+/qqo6bCeFA3xBO/2gKVWfl3wB2k5plw0H
6e81temS6PnhRTwP67SBbzLyISvXXs4RIpVGcAtkH79Mut8giXnzAy3aj5Q9cm/j16YPPK6EeFEO
oKO23yv1cvUScbM8VQButCCC4+P5n529t3yvKHWB3Vey7PyNF+SrHJX/G6CmUWMgGJSYp1vfO8Ht
twHe390Rzc6uUnxvkEfTkMHBKFH+HQijMFUdt99g6400VLZGw1G9NaKZIOgmuSfDTp/BwYGJYfMn
ROivUU6QTqbYVsYpVKbEScAsG6Eo+CaobI+2aDiBLj417iDMr9J6kCpdykNKRS7VlLkjiD5vIaMv
zuWI1HMphhjL5TsSh8CVnO+rT6RoHh/rS+oDx7i6oRgmNcRAAcN9jvYtefx7cg0mASasfc7evsEV
XXtsZFfpzZ497vz7nFtms1PzPRkYyduZvtM7tFdNjPj03JwpRCExsDiWgIyK6N7wPsAMhbucMlez
CYAVASPLmHL4Necn91TsgcTq5bZFRENZWdDy9/Ty/5tQ9bGDc2StMvBy9umtv26JJx3D1Nsuj/Rn
RoSTTgc/FeKDjm/xT3MBwmDDSoHJxUjgpe3/L/qFXZ0NSj5r9xFgSGdtEmOFwVCdxWTRQUyWLiEZ
7AEhfR4OO9USl609dxXWggKtL0GYQbbAsV/2T3b/r+mvnYkIm2HXXXNE1ecUlXVNwGrhQ0G5DVhv
8X0lMUBkBjVhS+1NAD9HQRfQWUt+S3yRZ8QCKuaCAnpJmnMbhZLZRlge80CaHKxsCFoep2PyOkJN
e0nDUVOAdZ6HfsHV0Tx8ckfFNoyRutQkYQSxO5w3X2Nux/3pg7QrlCNoGxAvg8GZcU+Z25yPIzUq
Xfy0BTX5GSirltgmDAedmuWFGLusAndGoifAg2+H1+4aCHmJv8wZA3IOiLCG5tzJ6v7QQFsuGkg3
Ux6BTAdLtcC1UM/XisQf1iEzUWTKWBwzuSSL5HTXkjDs1DYmaWc+FI5TokraHl23dLXLYpBljK5g
vTdT2rjEUmNURTKn31NcvMM7Hi09885LuCdZCakHftbXoK94aiPxlDAM+sPKkYsV8bQmZbpfv4An
s5mVnsFIuyUdx1xMv2h9dIdxuHBSGffEVSTrNa9w+jVLCIa3swGdeNDKo1zkgczrV+WLoC8C2kQ9
dosLsJ/XJTbp9fKnWAbFg2bYmVq+01lgFSlHPZ5spOeVegkz0f15XjABPuEi21dRDJngZnIErecm
NoMUVEMR1kp0gpe0KV6IwLQ6aXQPpXKzwZzdNKecLSXif4ci4PV9gmkPhFJWMc0egegi9dbmdYL0
Ghk1a8F4wwgeHemx34XQX8ja/2a92KiBuxy5rGo0QSgwpBvb5xp6ZdZ4KmODIvGJxZWM7nz0wJRY
5W4d8a5JHXxAGWNilhdr8UtaJ4jK3mNdmJrSUzmyxQZCytyVoXGmTDjAHbfGNhQ3wdVnHR/gcm4y
PUEX1ZV6gCXogHz6NXDfW7g/gORGZNGWvDcDhnsW7H6aunwUdnQKpybz4FrPC1gLSPMB59eqXg2c
XSS0E9H7jcZVRGMnyNaLmrt2AqIx/A6R6r1NA/NfiVzYI/m0r+Sqlo7a9g+EMbldRRaTDkcCPglS
B4n3WiH5xs8f1AI8zVHbJY3yiNNYsZY5MyvQ3hk2HE8NpyTv+bWN6fkBSqBbwM+fmcux1ryawF1y
F3xQeebScq/bHd/zpsF6FAy4PCRC8pI/1whf3//J9Bu0BBIq3ewROCGXl1MpEJ1Wu+T7t3psQYNK
/iVxrGeySkJyxpYwpk0KU6amzpgWYFGTUbGenVJkSRpQtKhN3anyQNuHWvV4jJBy544CYoLAjKi3
3vH7STFh2ruwcFvh8LZop5N6qDONAGOnK5m2qr8RvjvxefyluO9otlyEWPA/lXqgv8GJnc438qy6
VC1ffF60LIeew5m6fMlOFLZnEZr6atzI1EL0XXzEMXisUcDNOUK/BEwonFqTjEVJ5cWKHYqulWb5
XZU51PHieveXaadTB5Msz88SVXNrK1+F/Ziv7hzfVLNois7BuEXGwIm6/2endKkizOrQ5CKamFxu
Rc2JNQeb4++w2DYSH/sKjjCAevaWt3wdVpQovrlWnZ4VUgALjvTyTPeMBG9fug+nSFFLTvgtznfm
ctaa05VI+xOqKmH41ct8Wu7ZfEpHi/IPpjNqtvQWxqcnqOmCMKChXtaR91f9597C/igOsFV1vnBO
vGNHvpVEwkJp6lFaIv81B2ldYDngLgTAlH0azI5/ttgneY2u76XyOuzKxI1BJAumzevFvy1EJmB3
T9r+B4XcP38TAEkSH+VvkswT0P8UbB0nuUIrbdr5Umj5rlOF4tRR5GW8suR+o9hvvS7kTKZgOzrc
dmkixU/roZG1e17nAMvaNx9bQQDf/eMWFXiPlIAj2h7ehcS/rg/8JkpCJ09cXtI38+xkL1jd9Z7f
yLJ1MgEWZoOPtAy0VwVdJG4mJC2MnWHY1G5ZwtccyzzXZWJWgT/Jl24gE7S9IbIH2K9WWXxeKZ2z
3nWKbaNxzeWVjpjh5GnFs56+m10BqOMt+5x+1rZ26IRWSotp9rbcbjOxBRvd8cCXjMILdJd41/jR
7CHgID+wTgBzUKjC4iiJ8JNNmxdnS/EFxRwRtc0bveEEeVKMfd6Tr0TPe92NwAA7ZKl2UFxCF/sq
uTiv1QHljRV/MV/St0PZ3/oZKHezu2mlmZrJ31TYHb+VHiP2NJdbgPkrsfYXMrffRC2dDuyRw2PG
6lgStYvmatcTbv6kVm0Vr+c3CC+hoVYkTcMgUlUVlfMuMhJ+G30JVDObFCMir9RGg72tmE8Tvu5D
CsB8eZbgAv1gSkh9aq3VU78lNJ5RH+WzdNZGFGLT/I2WKYZP0mquKPhI0V0WL+1Rss2IpApGughj
53fr3j6m0j+6qTXCZlKMaE5UjWb43sbQhGjucTIU1AVkJzas2wVUTB8fBetQhd8xJxuAwK9UQEOJ
o3vGtMG//azaGlQP/2pAM5zR6H8PV6SvyhYhIcYKuWvmj1NowfC2gZM/aH4FxAIACjY0j3OW2TB1
yvixggaAs/OosjWqDOhwPO3I3/keSNPc2Mjr1dLO2UMRz1XFpB44gG6F8Cd/UcDI03bUWGOrU8Fz
0Nr+2IAVp5nhDhdYuW4CTsKJHr/O10Itv2/8+BQkvJ5Efy7HNMGqUZ40cTUAgwW30bsYJ9PAEcZE
CfscE0fA/KjMoKKOioO4lsvhO86B6p8Qcp++qNAdAxC+2qZ9PBhckdQYHFzZuPBAoUo/lBz1c084
wAuRpotB0NDJIHJnoRM5CfYRglYEbq0w37bZDCPQoJCJ0pHT1ABtjXgY5VDoiHRJrcKt0kM3Dydd
roGtxgjNKY4fUZTL1Dg8v+F/zc0Pvf6H8QuJLitBe2cwN+0Jn9W1K+1RG6+L4VROzdzPIGhSYNh2
ECfrhl6YcWR3hH1wvhsAeM2ncvw54zIi4xyt+MN9Days7qRNI/e7hZQbYCTf0K8wXpbi1QYoHmay
L4FH6kzY3Ts2MALfImAodsK6LTBExwL/LnOQ16FqyuoaaTH/I3AlDOtp3wHRymUC7hCopyf4UzNg
iCxo8IceEPda9mQ4b5/JBmsEY1trYcFcN77zDR0Ptz5DfWlsE3vG5vFQXzUSZRknyKc3qo4RB+Tc
rJI+ABp4AIfnEr5hEYIqLC5IiwwwL/dupQNYH0zIUJps4Qn8vmfrITKpWrrp16ppkq+mLrq50kRz
o5N3x8rgqwcwdIFdDiGakgGCLAq7qB1q33TKO0xhQKBo56V2gd5xvq1mKChQF336xs4VkQQ+Se0W
HWXHsuds+IsOJb55QdjPphtb4/8CmzWn59Z6CVJVyFuRxzq8ZWIS4wqzgl2TripFNgf0GEgRMS3y
tS3XCo4s1czE3tkj0/LRiWMGJTxC3mnBjZDcZ4xttfKZZ+f1xDOdDp6ajeXviL4ICrivbjL/GqOE
NqxYWNF9RC3C3nhIMtiuQKQJrp+ZGre+z5Kg2qNFy2pJ215o9x4ym67Xk7YKz3/Xqultg2wVb+xt
AqvtvzqmJJGDJ2YD8PHHs00Eny28+LSzcH1l7seV+LbZgiROoZHOLmu1e6r9qTdfjQaWM1pGh4Iq
z5WnWWy5avcZzcbrEmNpDrzohrWxPDf2ew8IbTEa7ZOa9fle+aYHxf/MkOW01rs/EKTWEO0NCOIE
9fWNW4hVb3Bg2uy6dTdoo7oMKor5ca6ctmwSM2y/qOwAfBudO6OXN1Xr9WurUyt1EF9FzIqTkM41
1+o3zuBS8HRmTlPR/QR8jWMdxVqfedeFi3qgEXbqBUOdmMM3KQjxs2V4CXDOGHR1KJUWQYOe7+OZ
b0M4mmw9mbpH8vKwK2hqd8lyH6Yx3eq16os29BRbWVVTNixk+QfOegvUhHQn52Fx2EITwpg0X5cl
7QbG7Uam5K+U0d4YOxW0ATANq2KbqvBlbbbhIkKIBF2Ns1BILgoQSI/xjuMT5wuq0sKZJuubF+22
ddP5XR/9EYFRSgDcOPW4vJ/0n+4HFyGkfzp+3Sj9gJ2vvlDXErz9w85psq9FIH0N4+Xy+vaSPIW1
c7wwfO/QQNYhuYCfnQcTYnh5EYThc6bvsbVA8/yLPDuVXIpvZwlfVC3GkCIdftRMOu0HJaterLFB
69NkZPFsYiIiMJJOkCR4Gg+5Eb5hW2vLQ8a3Rca0tGHDAyPorsYlQsae8xWWfxtfuwdG0mTgI4BL
tojLfW7ANgQo8lbz8mxnHW3B8f0lHuY9p1PNXaDYnEXBVrFTQJFeVl7QfBTIZdsKrjVtef9E/iZX
Xg9rzKmLdnxb0LLHeIaVW9hvKiH/oFgS45xQERo05DjJ4ZLYo1h+s8sS0iUSBudMWGlAYeDlLJM1
kJpFmgWngaSjzA+0ClpNOdIMTcx1jy5g3ieEYAN6rbmqQRMNem/VRR5gp1UXFSFVLBCHZpRaRdrn
/66Rh6MBkZ9FHo4rMBYG/1nUhvSMgs2AKV9Pim26xAXlAK9F4dJ6heU/skdKXpjbiFQPeY51XyWf
F6bQnBMtJBza8/IYngw6M/JxTeKZ1KkzAuSkLwGdMjCG/IyOr9u3LOQrKS4Q3CyhIiCStnocZGbJ
6NikEmsMXCjGxD/4guOr5WKOQCC6tpNv3dIMDRF2E16Yg9I2kpxxrmWE8mAcQ+EO3u7OTo9HnoC9
oIMWATvm89NbLirgncmYRLEhbnE2sk8ThDhGb6XXM3+3FtwhzLiShILV6FMSwKkaXwZyOg78/Xwr
T6dJrlXxEO0npOYMRT0dQXtZTullK8tBdJWkTj15FCdfdskTGgw43elGjn7SCzRmixjWk69kZ7s8
tdsnwQT2pmOcN60pnwq93vxfG0jjUqeJaqlyRqINif7EqNi/OjeUtkJOJJfVbqDCXiw/etUiP0b6
Cxm42NRAFCYuLSJ0fY0D42T9o0/plhJWlbrOrrU84z7e+VoWfbRFn3urhAGNNVtzEcBaXwnC3InE
ZuWo8PtlIuYZsAcp0tUshc6IA1P6eiQFyt4S0aAzxGuedamxgadvLFJYX4kxUOz7G5rM1NcmIYA8
NGDIwzu09/ycsDTkOhQ6Yv1allbdqLn0sbUA3SIU8Qp3zW4EOiAfAt2rHAXhbN4AcXhT+eQg74k3
RiudFdHrXZgErRJ29EZPJsYISSuVfvoAM6NQjhEixcxFlXUN6kEREnPaGtnuWUydVr+qRj2b+8Zq
a3UzksVhk9uS84hqEMseszHSuuhttcpIEh/SMNcIcFRvWLydNvOlos1581dD3XNa7aBdTYQkohVW
c16NdqhwvQP2LPvhs/UZNLS3bwV/FlrPCRpxdxVEEIAvbEh3jMfgbY9mHOl8KGgrfW8Kg/waMxbj
svCTHWa83WLxIfMuHL/JE212FO5cB4FQCPsoTQp7k1+Mc/269Efd8d4jXxbkQrZmgZZK7BH8UP2A
nhS5V0uPaP0puxFy4MnlHW2ZEwb6JkyJoH7qyF4VDM8WxD+hbHR4vPUfb/Bd66q0T5WSOney3tfg
iRpobNynJJWexJ1PQ+BmsPIKoWpjSsNiyIlXaegq6ElKmNp//d5GVKTxovEaznhZc6/3uXtNB5BK
hPv5fwzzb+MlBe1kxmx9vRmjHe07QBBnsro3DnsumcX1xzBwNJYpZ2lyxwJ3YQIcmZ16GRwGRsDg
o5n9Nuyf86yTruxAunaUCl8bLtiP/LsRqiqLgVrGIHh7+6g0nFs0G0PJvzZooYTngPWJI7Qlt83W
6/8c8wUCqc3H3nEc9l412VLre1hpIj3YyfuhsKaW3z0WMQRBt9S00oPY1MM37nw5yhtsR7s8Nsar
69lV5C0MQtk0uJXCIbOogq0PxZ8NZQnDmpir7pD/CGL08XJkMxaPMhXM5ENgS3b8SYDqZleYx+Q7
x/JYJS/w8AiPU3GSNhrGcmKkyT6+nG64OWg0Ds3k2ETKbR+6/MgyvbnLYByQvc6VJk1EP1IDHz2l
U25GR90RKecUX7MPdfTaIT2AvbnGzL9Ok3EanufLzK/4ww0bDGIEnsmgweZ8allKqFMlZNAqBo6Y
4qa8ytwRiDqDuViry85mBTe/vG53VviXAnW0f8BVSFnVkQ/prxkq7VTZVquHjfvJNLHd5saWfWTa
Wd5NuqUur3Qa0Vk8EFlwL9XFOvXFgfrbKEj4w2kf0ia3x7cMUrU1tOHMQs8Aj6ZLyDZX8RAembKn
DEeQ5OYhO0PuJ+oSfQou6LZPqKQPDkrX5kEebc62Nxwop+W1rKK/o21rWWFIQtlk3t6pVlr2JmRS
Du5ZJ4m78tYJvvkzSfoWzoMqIZ/Wb/dkdLyYAoNHktFj9aE1zz75ti1oCY4XtRcV9ur+PEz81OL+
y/Zk4aSB5MhBe4bKpvWyWIBeqo+TQOWYIyLghqUKofXYytuozQzj5HyOClcX3v8ycBp2e2kLYLIR
CIuKvtSLNpILYCfZfJcchXh38cSYvqk0cF8/CpAHzctW3w4QJhOvSSwZIJ70gJ6k2PW3Stqs8BNZ
uDqegrcMxZzkSblP3EJS6nrHffpAMQiK1cIe584HOoIqgWb/iaoTosATS6VGMVaB5wRGH5atX1BD
icoQRLN9INnbjtLQ7RL1vNC1TGKMKXukXCtff5MT8kG5zpZopxIDur5kQH3gVTzPj8v8za5OkhMP
DjDzP7izihgL8VdNWSxrla/Uae6WxCcErBqQXWB6+hWsj2waXB0sXqiQ4DquF/nb5mIIFcTbTqw5
ykofuusMNCVbjsvO6KMwsJyKqMAJVzHk78WV7gl1GUkUr45fd0+o0vl8uqZ0kVR4DpFIb5Ko1hJM
2yOLtLuLhtewQmc77CGiy0vRr22zZdbnFBV45/tsoGMjaFOU3YVhzrsfat1s8IFHOcwLpECe1PaK
CukUhisUEFbPlVWR6XQ4h3fPSp1og4fqPMykuiUAHgs4PvoSh2PR0wSzqwM52mtXy2fl1EuruQHH
jy9koWzO62Mq4IVWtsL8IrcpXAHhyGYcaASFaxRCjsfFhKElAl1lK12Z2iBdjeFdZHR6dOabBaGl
A/3S6aoAKsTCs28yM+CJF600h5Oop3fh65IKX6bdgYUEYlDT7sCVuGrgLkp7tYIA8IEzt1BpU69s
ttWDyiRfDx/YbLyu+iR+rtHpQUQdm0gb/9JBm4rxnmChgEoVzaPUn8iuS5ExEL157CiE6Ta+92v3
Y72lvgtwFg7LFbV8rRiWJq8fQgrHKIhERGfoiJrvp9gy1Zgew6ywooRS1eavohs6OZyLazU7Kxu0
mqeNk2YT842J2N0D7lG0ekiQOh9j/GeF5dSNRhY//lkEhTyT8kKYcKih5tVtTovsx4/ERhbteTKI
pg4K8EgePuVAZMEbjOu4yD4sQ/GaOmP5IpWkcqJjDikU96bqSalWQhW5x44nTpCGCn3n46q/yu3W
7eFyfeFgeAgFwwMsZJkAG5D+OCdExMed9xtA+ZTmGDVRkGGItWuYiaJpBKt/MlHtSlAdVKxV++bB
B9RTqMGmviGuoLPBe4s+2KhLbtmqT45uadyPGogvp+296bCKvC44XLvOotajGusSM5YSUMyJlUxu
uBFMlfYGfmjkguaOf7bxcqIuxO89JfOZfw4YgiuwA0aFgL77eVrcGSwxz0SeoweEz0Sl+d3yYlx0
s/sRTfpFci5mhrpVg4q+ZRKhSORYczHfEktCKT/aQJ2RKNliRZHi/2uX3lHQSOQRN+++Ek98JzeP
bXvA7BrNC4hS5kEZcucS4XKZmDJp5+aKW5u/PUYM2g8Rmz3uxAvmkahZiVf6G6dNTng7LOnZlgac
8fFnaFo/bWIzXPgQSDmeEQlF5iXfO9KoArT2mZV8M6FuRiKJLwO5tL12Pz8ye2CsphWFdh573Mkv
JhL0pkKWZTmZkiPlquadUWXHxzKSX+gotE5ii5tgJ1mg9NScsMnNLsEulT/1LfmsmL5Sq++PqUus
jyoFJvy+ypBiwWmkPd5age/ZYvp7laUP6F2U7HGKgE6ytze1fl0czF23FVl44vVyc0bsik4wZQ/i
rcZZwpxyn9m6PiGpxcd5UShZgySjcLslnAyM/K0PlxijFyQ8SrYGU5U/hdtlpK1eFshXpX4C/CJd
Dud28i3lp/DCFZIBqkFEqasSiPY0v0EjtlgnGIoVH5JY8iC+CPQZwT6MOjmqln/l9/Ry01cyf+Cp
zVOyW6ERxFA8Mj+XC7IJl+wIEp1KuzUZpho4fPOcuiYQkmwiKEr1EIgiQUIIqVJjnzq6DIA0nfjH
OqSB4coq3yRe6/e41szlp5sHFO6Xbr+40M2u8iHlXzCcNH9WevkwXQ6cyFzDK5FhOEy8QcDF2gQ5
aDcfUKHGgyfJLX6ec4Bj96kmzudsxhd+pptpDj9UNib1wqVDZPAb2NylbRL9Nyrc8kIt7tITsNMV
N3NNoYB9Y152zpIzsk5eRKOWWVq99jaxFSbY4P7T0nxoP6+lSxrPyy3XPjGUZ1O+3x29EDsAKaUL
Lwwi94laXITDatE8G+gv7A9hwMaw6qEGaUHFmP8Iarue+YcugOeT5O1DIbya9nksPtm7+d9RPc3C
67CHXBp0c6jRVuBe0h+xTN46nEvA8qMHW5DoLg63GS2ovbkVybKNzjK3FvmnXGnOSXVhJb48RMG/
Dpf3NJeVJ8k43PpQD65dK4rIzoSN528SYbYYb1mrJFXypDaiaX/6ektV4fU0BP2Pd47tJ3AcRBME
nHn1I88XyO9c5UU5JJYScKpZOfEVpENx41nXJEWz6TDWDoYA8EMf++8ddibPzEZVJNTtFyA4Dn2W
pqX9yEq6Zfbvt3dYXaFWEFx3um0g0qNz5uJf6oqKWFn4p1P3EYM1X/PlnXcW0bOripOsp+4w8sre
giRla99Qf6dyGegXr537d+MDGuauQppT9RSH5srjjGRSfKbgi2F6JHpNqjtzpmcNWl88pWClBwXW
r46Tlj4uqatfMbVM13YAzGw41SiPjIB2rNjRUnSj7LYMqGKPN/APxVlknogdLet8HyeAEMasA0K3
238PeXnJyvQpKAIeK5PRmcThIzNveEJj/FxAu3SNDE05fRlFHyZPZOoC+V6XyetT1VgrDvtl9Y0+
sJwiA7WAdWRv7Mtk57Al89jsDPmVdeoHYadNGLHv8Url/bgAGhySE7sqU9vg86c7E/rf9CSDO59W
gp8IoQ4TN8hlLODSGZoiRFCz0j6/rKY/qf61YFgvtQn2KPd9q3Is9Jncsd61WzVZzZAYWRh+A3P3
xdZyOmGFGwwJxPMH7c4ukMeDDCwKjNg3cMuQFAPyBBNR0VSvhIvK0NtALshGCMoXTTSuuPs1DPdN
PKAT/Nupqn5njjWKVeoFcmtWAEtOo/rL5vyq98/vIbcsXsbd9G7aaffftTGSN24RqRo8jYxAIRIs
XSu71QP4ZyWLgeUkl4BP/J9s1+QSqQCsjdTt479JV6gCxTOG6UIBGpr5JijCtExbWQmq1uu1gFIQ
PVSeTGfBUFvDy06W9HCe+/qMotKvCrapz8mtDRoKd8b4pHLE+32mM2bT61sKQ9uLxSF7rt2N8RHt
fA1LruVPa9V5qNYz1OeKuVgJf0620uLENorAhJ7LJ/pS+OJyeus8XOJO0wLLIA0uex/O5JUAlaAZ
z9KrupuugyS0c2IHWGLNfyfhKnE3yOutXzOsWP0kewpvbKjhstI+G2iz9L/LB98y230ExKAKmpZe
+KHs10G3LuxMEHpOnjxgsNpgMmgQU2hh2dbok8Nl3z5/ukT8oxKVbqcXNkA7aWpoIYKqZatzCWU0
97IDyO2buUqP/SaOuDIlZMBJmaaqq6VBgfk4UbhvhRMTEV79JPEFOQziXqwNbBbegNuNsbqzx8Gb
bz8r2TRL2MN+ned+7ZQlQOQvWBNdzxoT9R4yrCHDsOrXWo76s9n2evdO9YrFH1dHGAHPYp2aXd3P
WMN5L5nhPshruLarEwpTEW9mhnpvjiqLZ3sZa5PA8QNm0+9P+q20VxtSTY4w7jPles8o06lgwj0O
z/GDr1rPZa9PD9HXD56mJqRWquhbh4lhM7KzRLyP9u+7ycLP7a7JYU3HU9p9K88gfoDuwhKkHSLT
G6GIzYGCByXoAqvGT2a6B5E9mp7MHYSyM2vxAQL3fOamZSJf82etdCZtcNywIpJCWeNww29+y5mb
zrUMaoNyeu0OFJr5BdJp2Km0uowUuJ3snyt+A64IuE+KMPDhUNXV5/gizmOyoBD3LyF5dUpprcKc
f2vLYLLtyIiRAPaTjhNS+il9jFAcuNle4KpSjjPEB3RHdMWRgtPjYtTaxhHmwfliX8fVX/AVlKOd
1n39CvQc/PkeWGKH9oatj88qaWU5glrNgjPfvEr590Mvq3dtfPLUSvV462+Tijm2H6QGT5//ErVw
xAucY/KCZqqRLip2mqJIm/d1BzCKCA5gi3sy9dskV7ZmL53k2GA2vBWMrDEwue9pKoKJw/YfLKlv
S93s/usBT5lVCxEGOo+Ioj9R/Q2unke4HNTzPgKFVj7ZSXYTmndNlSB6VpYGCivX4LCv/1C6ezWU
1yateXpNpsIx5S3h6TBqYVsbwOAi+cXS+e6Ks00ULXN0JeGGntB6esgGxAeJzfnjRdijNyctq4wE
NbJYoff/Padva26eiad1oHUpYodT6S+/GP8utJVCJ92+sH6hGX+e7ZCGx8WdpQQhZHwFPSBsbE77
Gt8GClgvtIGBRwvNOYzN8Ukn9yhys/KnHldapkr6CMunocri++bGZM1ZtopYec9G62IghmJAU/c3
KRxZtuoEjjHzonXsUraHLWq/dVgj+01RWlUPhDtsUVajtLJfKaohyDd1cDw9qJuNk4Sw0yBCaMeV
XhgWLCALGgxUfuBjY/RbKIitm43zfTpnTzLhvE8DVsXE7XkMmIP6303prN4p2r9Aaztc32qdO6eH
aBfICaoiaciogt3gylg7PqMz6YTaufX6bMRK0VvXMUBBm5Nf+ymaT2g4GqWsReJKxbNd9nXpioyI
zHVyQyt+buUUk2fXoR5kdaUQKac6nAMo+fybBRmgbEzn0dyU+CsGpgpGxcKjVpNK1/HVIPbcbusg
yjXKUSQHnQ3+QSbQ+ADYPOS1tIlv7VADxZZb0dq3dw0sy29H+upPF7jRZfxjO0b2dBnGSO52xQps
t0PytDMp2xs1Bj1QjJFnauJx3EbvMeA/6NrNuUwvDgYsACJmz1A7BX/YtNCfrZnOe9thudzZW0C+
dK4SLBluF4K8GZOsYKHpOc7Y92+09kJbPzorJ8EG2pVAqGlrodXDfFE3w5RpzXZoYE+gD2BxiIWW
wH6t9s4hzh61gPCOwq/R6rqTj2YuoouWLeHf7DIvGfuB6Hs1urO1UKZA8P0Em0pGNAHahnxW94lc
vLJF92jgf9GR60jFdoVBhQtvr/PHcMzQQUDIuC+ZDlYecScAK2mieK7kCUdLL8eJ2ZBbnx6CIpmO
aupYxvGPOTOxf+gC++A9vaOj/sp6gAkklV+lfU69dL2wm9Yk1FZLONcKUB/3H1D+pE0u6F5bv3tu
XurE+/3Sut79KKDUA3NPmykFp4EZUJOBqpDHk9F6tOr175r6P0/71jjpM4zr/Hxic2OmdNco+vee
CGtyjlqU08CXc9A3klrZMcmUja5hxA6WcAEfLiAQSRo3eIi1IN3id/tbY5iOURZR47umnQiMWluk
AwnrtQILREZxjxXg072IAX64hIjMnHBaxJSsoILZlAnHtOLc0+R3hAcHq6JRL7jcbo7vAn/u4o1C
jCVx68UJO2W8xMnZ5ZwR2HtapjOReHdyiuKOv6z3L2C58wbm0+9QwCdV3dcAD1P05FCPUDtCb/Pu
k6MBuEPKdgXE/bVHkSEvVch64tj61kH96Q4i2jJay+EuSmpdK9IDvCr1GQ0zf1QevD1WLzIUqkbv
45kPFFUBKURj0I84MSzzTc5pePeZTm+JLCc9QBPp5f/KVfb5hkNWKbeguL5DT09m9IF2/wIg0W/s
b1cvRKKPH91cLalTRFdevu/spn0UNb8foymBeSbiiCMv0QMBvxs64cjWr/xm1+fPx7qKkYYP2h4B
vnP8p4BlYEBri4HSeJofjKEVY2DreXDWNU3Tp2V57EgxWUhNFlUfKDAZJhULiC2N/i12HUEnIBRK
eVvkgiIDQ6T2DKS4vnxUBhuy7oDRzfKSTe8WLPY6qEpNTO9Lljzl4YEU0B8jaR08CiUc84EgVQg2
K1AlvGpLHH7XT8JcMmEU68IeGHUJrXfxmElgkNarn3uJu33MQkGSXD767txlQGsfm4TpmhQ7n/+F
f6swoCajNjxc62e2EkhV0S/gBuwKKDRmssDCwx3g76dZi8cbcRXoIg3yepB0Vj1pDDw69PFE12GI
X1upgAnxygTrFNH8Vkxq5ZmCnKoh4U/At6Lfp323h1b+RcjNhtPx+0zkmAoVrDzIJitnEMjSnXs3
7f7E9kKGc92rX4j5UAvz9wPtHn4y8evS7I/3mlk0CXyToiTc8VsjYLLSOsaJLa6kz2K8lsmJAC5E
I7fVrmP7E8KVmNi3GqC5bXG059F+rNFBlq/SCBwwMMyZFDpzJmirpRELecIPa5ikG4FsWRjJAwKb
JVmnObzT9xpSjWYlzVZ2ihIFj2b6YCueRjiHR813Wa++KdO6jkTdLUgETgdRG9pqY3tFNRxzGaAg
SGW3yJ+kQrUWgxSDj98nrehDVUuIZwBB4flNo/WfREnge6ECo0LaeYkON41X4+0yXfmSRjbawpT/
t4jaKzVkuG7yAvwizliqBmst/Z5yQ1b4aRLZurhutTjMjYcMO93PH/rgLmJUOpuRnsWOkqKTZY9x
0EHm5myn5kGD4p4sGXNwKZdu7VXLxL3qykwu4eTugYKfaJh7f5Srb6PvRuCCvJLGDclLf2Okr9vC
bEOlEW+JKg3AkHGh+HFeQMOYq5fHm89dVWTdTJBui6KdlO9cmMqJKWaJ2iRH19GiPyTOMwP4nNJ8
Xk0qzilood6jGEVMLV6dPCEAewfHM/hysA1uOyc4aljfIpHg1bKXDAHTQz+Okh2iGFY3CCJxDLyA
qn4xUABUB9iw9uPM5uMXG++C6Bf18Uw6PQjTlW4PytFyVA5llPzWsQwhDoeWoEUzXeEwztXoVcye
e4Zc332A+idC6ZNNQrAllzotpgQzlRLIos1sva6XBdvZSyWBQsJAO/V7pDdi6PmfcyMm/kz8JfWu
yppfz9wnT9Ou46u1EdQkAOqfeGjxQ6g4Ic51jbe/C2NzONPHdGPIEjIBB0pddpx4kjsurLy5Pkc5
1TPB4/sFJv0oX+NvUC/+I+Ok/T+n6ogSbZfnnBZjHkv9pS4VKxdc9FYfD0y1J4Pbt27sQ84FJD1y
NMaAcdWxOC15onBF94DxQhdXUxgxsDoXus4pJcZF3G5Aip0NVHcI4XeH3PeTM0iov9fm3Urp1c4G
NFvRDyuj7amvQofqIVvmHVRaLDzlc6kvipT53XE/QCA5yg1T7+EoeOU455ogIC2ikGSOUOGxWfXu
EtcTMK66n76QaqQ79pR402SEH5zJR7RyRSnOWhIO7mrnkkMw0uAvG06DsEe62asxy5NDGenjiRD0
Brkaw+V3GygzAZwixF+qjiG1Ice83fLDC7hvnud1MGyp/frgeZJP5KiXWjufGz2Gy+zYIlzmp2pW
VzsgZO5KfUsqgE5/UW1gCcdhX4z65K43t0rqAp1cF6QjwO6Y66jhllsUisUQkc77FwC1xozNeylz
fw6erfwDPncmuCeqp916iJGiyzbi/jDRsxlTLLzgQ/vxjK0rr0M2H6+gR/sjTprZUqXB+tdZ1AdO
DucC7u+wXgjPivq5YONSS3saXwBlFQq2nfTg06surtBjkXIwy/dmZoGa/ryexoMkRtsGXk0R4U4W
YSnjLCnaYmFDSryEL9lbYbnlZaMnkZlauhxoc2m70J6oVvgXRJhxgZ2CpoXTbfFULV8arKfC16+X
BW7nscDq0UwzrPVGYSK+JnyGraGz0O6WVHk2G+Z0CWQKE5oGsQV8+h/dqaqOV7aHNZg/uy9FG3Ii
8oNeayBpDMbvgAF89zk4/VbNuJtA7HR6lomsW3mY81uayT5/AvTWgCuV27laR8MWmQZcgXnaw+8+
2+JPFXQO6Ao4ytb2su+d2W9p0nyptQSNZeVRrOLJ9gnguRnDWEU7rEulsQwttTdm7mxdbda0TKZf
yLJ2/vKV7SW8WS1xyNOg1CxJAzG5A5BIm8wceEgIjgQICqVUDFXVVKt3hawF5Jy92tKwKVcZF59V
rjf7IlHPGc95EfFzZV2QBNVd6RFUNYon4GQpXt+tZnaZH2rJwZKrqOL5SjGIWRBqQdScD6s+10t+
avGxC44izuhln9ZC4FhD1WINb0HVvahiGwCzMq4CbXSqs19orPC+SnxN7QChVX8Lw7QLMlC1GBJk
amnW6+M3aGrrJLRxW/jafxIegjSUWN+U3A8o3KzMYPRD/UIpAseg5N2lly8bbcoWNvceujI1AWFT
dtCUbRluxy8EJwSL/VfCurId86ZzEbV7XUj0dXc4LiOaFnV9B5s1QauKpAl+LaNyOI19l19S4T8Z
d8MVVMVgFKLRWoPNTNowbeLLDBaq08GBg+E1MQtwfXjzXmi2F+TRvjnqqROdO6PPdQdy5oqNDQTg
EMcDlFb8HUSNKA+OzLh++Mo0G+Fo+s/YvKIInaYqkwafALYhi40uS7djTcLh+nkPIy208A8MVZoU
/DPlmi9iqOZ2DBEZWx8Rdzy/GEWx8QQwd3utfDvVIkqJnELFn8MwUtaVwb735Fqsr8872dqmEpQp
buPnnJPuEjOCseOALe2QyRhUNsGBjjM2IKlZTiG3Taky8S/kCczHm5nLDkzszrOmhe3bHa/8hkf0
A/uBxfWNNq6SewNGgysLOA/hTibBbZbiwHM49RxmrDYVAo5BiIxOFnKTMS2RkoyeFHdE0TISiTl2
yAcrA76D0tHbHj5tP0ge7qseFwJ15WoTU848hpsKN8q6UbNUipoDVregXijD4JK4e8jee8l/B18B
2SlHYQnR4LdThP7o+ifOzovGfzU+NUdSSuz6tYwor+FLV2H+Bt4usDw2KWBK03gLhfB8xK1pWMpb
JQX5RxJxzLQ5EK2wc8sItPM6gH8jKCgD6M2fo4OToMCU4ez9IpbmP5eVj16E4480uYBT555Geam6
KJ5Y9foKvHrsT9vgUlJrhlOJSlYNkM8BaA7uzz0eFvvqcQawOZgK+gnLjaydvju+R0oUB94qbSPc
MGz2mqigjfovmuvf69RrM8rtiSmkTrRcapHC6tMxoJ6jPNrkLuQ8xMSYljPuNXkc1CRaauqMdqOY
v8kLkNdNHWXKrdOgMhdtF6DC7B2a7vjME2FIjAPqaQZNlmiMo4Ve+mQBIJiTRWfEwCqIxiyGpN7L
t8JrEyudSfFP/I9N0Wc7J5unMJOqTi/X42p0Xy/AxJONHfShwIty/zNOt5I4VMahGEbnM+/uOW7Z
xQr/cQ18D0mxL1ku5QJ9Eag7OqjnAKcPjEaFDH1DLcZq+yfocAVgeNURdo+IYQbqaExiwqjM/utc
tZASKoNxQCpLV8nZN4+o1ZW0gfHi+F4HYygux6C1J2C4Nr/rc2l10OzotKkZ6NlB6lDoOEzDWNp4
221e5IJwkrIYISRoQLN7GYfS6iAfFUWlFo86Vvbt+eWXWbBrIUWnnto2ey5gAtrWhjmYZIjK7yhX
r8n6NzqNnHKIxy6yHvu5Kg8rmlPsZhtcOPagJLC2nxvhcy3dkUPH1OqZux34sx4JPXvu1SC5YLyH
9345S4czBGOgVfMB7g2UXzXxm2nOErh3XXlaTvll5K5sow0p2M+ViE5xWgZP0fACYtE5O4X9oVRd
ssaVjkACQA/YLjyf3emyzkfoalFueAWA/nnAc92iGXcgoPG0UhK12W6o0IlplV/SF3Ynjh8ImLLZ
9xkz2aNN+5CJ7mjbZ8r+jljHyME2bvlIEcbOwLS1WIf1h3qhSJdx+Sp0eU1VdDRzK71fOcGz7Sar
H+3ffLse7I6w2DkqOXPB70kXgLmGPSmYJOiLPt/dTu19Hxeuom3T8x+8tBXonxpCYmb6Cw3pP7KF
Yi4jzeP8Va0G39D8wBC+TxD488ee8a+pni/m9/y0yqjopIROEQCiMmrWc4/UWvXY/i9oqfFZoYrA
nnQizdk68CBs9p07llCF1/GGYFSD2Z4TspIpDYIeajNqUPDxzMQ41EjKXqYgaXor3vgt6IjJZde3
yK+U1orUDCTlo6QTa00Bkv51xA+E1nhL3PqG6YVdYT4sqDUSR/cfeA5+C7pQHnpSbcr2CCQwItNk
vyK9tGVwOXqdqynWMPWtEOwNNMQ0nvCN56GIpcthBN5O/TCUkuwAIVke89fdqZhT+Rv4DG1R4q1f
d175iHX/0z5/4LOQ1AJUpCUIPqcQfThFnR+qITrNQxQbg9w97IzmhXVQF71QfsNaYORf8BJLyfse
+2kmp0xztPJZG/7Cuow2ASIGc9g4ikypIF83eoEZpVDI4FM+fMv61NAM/T5MT1LyIV5dusPg8pUD
JZsGv7j1uccWp/Khs1IQKC4TYS8wn3/Gud/QA8hoRG1rHmgnERMYqDseocu9Pkxv1IYefP0+QpzF
DUWL6tpKacucBwXxbT7a+cTd4SUTk9tUGfdOE8ftnVcBUESVvfTc8LirlF5RJdNoTc1jOmxXocPR
fTZQR2tymnh+0x2E07HGIo2EOFXyTPszSr0IZWOcXRvukKG0P8/PUtSeCQlBNyWTz+Om4Jgyw6KM
RBaIBKusYSdR7ZCWNbAHgBBeqO+qEVNqP4oN7uGJTVCddxtX3xtkWLlUdze5jxGFVBrFoIT/obFg
l9M6xNe5HyyqRLihJYlJieTP3Ipma7DX8Bet2LaCB2HuIT3GVLqJ2P/reePqV+m97mY6VT8yJgWo
U7WVO6a/AhQztRYkeRBYtWVHDCEGhgu3hhl719zJFGnL8MGC+oEH983FSC0gMomcZfffsbQWGkkf
KEisxEeePgf65SqWrCzGeMcQSTVCo+9WGKawg/HFMeFXhs5hnMO+qEAJ7i1iWBg+xif/2jNr+kh0
YWwWpQ1ywNo3ZwsBvvd3a/u+Eyjtn4YFatNqNWXdu2glEC1kRHPGE/9Zm6tQfGpY8xCbg0S9V6oU
+l1VG38o0+UnIFWleLVn7p9H2uu3iHBYKL6i4ETe0Lz3eARTNkT8q/dffBXoIjZ+/+DcFXkQd4yT
jDoAcq2YawAoMbNaLjrZ7nzEobfNGK70bMEaT0NAgIKt1aPHzz2/7dsdAV0XtO37i8F++uFRsohG
TslXYf/zyVPW87X/fsZJI71ZXlJG6gkyp7dkfcWbLdel3gikJsFZ2Pask6cdiv/AWY/hY23x+0AB
um7+AFS60YTEQVOdJUEe0KbqbggfkMNwrzgw5PyAwYqq/2flvtrf+yCtfK7iB1DR3hPKh15SXMMc
l2QSM+eP6k0U9GoAjAKe/r1l9a7Hpje/VnZVoSEHYXgXPlpAUywRhqr7eE//hUnJPr0g8isPKpE5
4zEAreFKDV5zuqp+Xv/cFJQ/l9RBUSd4/ba/0L+4Iw3O4rSCb5b7UNmECmdyKBLVNimB0i+wfKGP
t7m2rBHPPiQrZEtiOK1JFx+JVSu2e2QLvwApUeJ4yNJ0WqwszKXGE/gm+ryb7Ip9HDzJjaoRLJCm
SGzxzPGMrLFlLXwC/1bpYrVJgVXz7t/MODUgUO3NbNL9545AslQ5bD1UFlyQzNePw3EJrDrp6x4b
cCEOxiNSgo0O7juZ6l2Ys6AdsH63xKH9kyAdHwMgr792gcQ5EtTUaZEXBcjfDd3NWACfzBZS9g6i
jdKRqyav7qaTnStGS3BI2mOCITTOPbm9AUPjgjMjqND1su4MxWrdjdgx2JuD6m+29hP69H6VFn12
jyvCas3dYCx4Jop7gdf147rRkJBf4pFF/0gLoO9rRDosdcvIFwvWgmP0VvZNtE+QDcwl8hlEVKzf
KPkQN2rT9GHpAEDQ5UeyJGEcSBIRIvodTMwEoZmBdIRBweDXWSfV3c5YXMmHSZ80KLWHh3mS8ug7
/8bdW5ghBLYYaZA1BJaL7QE3gqhBhpRT+bMMtfLgIclZpGReNs0yK3oA9n4L/x0AP/pWBQiLKYAw
JN5jsKy/TGuqzYovS6VzUAz0sV2PcokAmPNM2ATdaJCSdPzlJVA4cCJVkAsf5p08UaKAlKIQqY2Y
4TPRAnKz3eJI+TRSMUSkCFXhx0dBrD/CvmbndeU22E9Ig2xsYaR614bigUT3lWNiPZXaYaArDrOW
1V5xzFwqiWLWInAazjY5ylAPuTFsOm/3qHzjwZN0+qh5ithJ3+gsNsTxuQDCQ+6hMjt0T3Su2zVM
yM4xoFKTHt75s6nn6i753Ke5ZtjIItKYwaaOMu0JpgCbiinFDDtTJIR4c6/Al0VBnm1BrD2IFlPd
/EH5yxO00IlurAa/AViZH22XNtBO8YLiCLFVBedgNSTqVsoYHXI4WzHKfaX2PqB4qHDoA52vmINR
Y8mKG+gzTfgDm7t/LkGA67dYnK1l5CMMynyJ4YrC4Gg2m1MHnHDAPiGqnWco5Kx5Iu8vVrClyMxt
7oPvgzRoi58C0x0l9voEIR9WK6p6LERW63QpmcdOKeKSAPXtGT7AXMq8+4TGmfH3rTH3NbzoO2ww
o13VzSv6M9cqDxkp9BbNx70aALbbnktYQrH1k/hqbhduIo8QiHkgXF2b8r/+KKxUIVYi93d7BXW2
J0F4gUiWFWX1LftqVys9P0qCuWnbwfuEKiHNMV//pDlRywzJFqSYMaZDOrfYU4hPANZ3rM9uYXbN
9n34KX9mD5NI/GxrvRGDCdMpxlYhDbgwpltmwya9dGsA/pQ76pvy1Xl+fGfaAStcK5QqKoew9YZN
4kLi+CSI6vFsVUmV3ZW9FTyaGIQVD+1IblX/XQR9aDpqsGfIDPC6T0kQ6oNrM7pHwesGC15BLkgF
CZh3nkKwUX7PzdHKyqsQnxHapZat1orWdTz5aY5gX8/AowEy9ujyyEPTGASoEk4XevQtrO9dtBSP
lWNZmnZt5GU0WlUWfpG1Fjn18doFR1STcYbSP0PwiEuuSPn73q1aCrFLrmx4l6K8URvi9NvF1+wi
u1o5inFPWp1HTeog7i6ISPeJCnb3a9OvlQ3BFzOgcsQe/AcMuUUQzCUgisW8eY+zF+YEKxKqvCNh
uryDf/k6TKn/qLoLpDKSjWT2zDLRJvFlH5WL8EDeI/dHULPPXXBwek8mXz4eTwN1vtyUWhiTfNr1
eaDcrjP02fYu2VM8is0ikFcLVouJOpuzrBiF1wzwIdjFOmR7sSnlz2YunXTuDWnTQBcutOsDtHoB
8K1XxFbS1zRAzDrHkfhoSis7nDtsBiRzvzrZ16ST5AJUpu16E2LimJQbQQV2tCdbZY7YdO9p8B/o
NrU8t5WZj2ymP4HklAr5VsSzuFwUAU4OoNPt1UR34QMqZxcwzeUUE3L+nPuSHqzi2s/+pvoThsWL
4lgohFAXLbzaA4HXmY3Zd0h1sVvjuy6W/kE1X9RT7YJjp9lINzE5ZJyrgCiu3m5MmGBWiiSBsM4+
VpXsKi9h3B/iK4LR3rHLKdb/ky7paBu2C4AxlcGXOhvBs0Hm1eZbM7dPJl6aowS0PCI9XnEDbgGI
Sl3d2XDx00JydGqeXj/QsYgI0rWRIHmkmsL0ic7v7BZ6lHdWdKFdfJ2SgXTS6OyDdH+WQnICpx4s
9FY7T0yJI0e9TSeJm5OkeYtEEvK3NTdfZq2NfDc83Sqy66idJb37creRMyWVgoyO1LJJyqtL1jp9
aq+qPC1k26RY/LzVDsn+0AFo2iOpnsT1GRIPthH6ILJwE0OVzZEEvrWo+FhcThkfUJOd/kbI+mpI
mZAdk77GOcAeckQQxijSUKaW+f9EAsyiHKB8yeVdZHPA4RaT9D+W0t4D2oxOPMwJj2syBmGkDIrg
ASxlDHO0XUC6NWI0B4IDCg2MU0nyBtQy9f5dHzdc6uzcJDqbzuEVRL1tfBnVdg33d9AkAoMmOfIA
b+S7QwRK0/+ewEJ49RpoDqM+HVO2OtICJoGTAL6TAOIW1fQzlxFDiUaGzx1sS7ufSwPWwaCZXoou
kC3Q05yYUFDlNKDlc9purlL37kJzsXBUVRe0kmHA7YXfE0SrVU2Hq+OBbreuYD1zur/Nni/l/BIh
fVjMMyNwZS4Ffqyjq30nnWp9MygMpEN5eF8xj0U3/0mo525aGMQAI2Dj7/L2a3zvIimCEVr2E1cY
YlLyv6tmqFHdfzVeTGWiZycJ+8hh6Q+dz5ClWrooNdJU4A01GllQYhS8vn9OKDeV1uiGinEuq5cT
haLMKpf9oq7S8KIrPKtfGArBeUsD0A5ah4Z6jQnLnC+MOojY8GR16QJeX2lphFxWZ7m2LhvxuttT
KHSumO8ShFhD/R6/q2GT7ovhb/8MjHNvUEcuf9Nv3BdQZdoMxDn2n2shpmvyt485Jlv2WGyr4y0e
6LbRqKA0blC35FQ5PfIa6tKwxUVBe5IfN5BZua9QB3j3l6OnFDZOiIETZ/c6P1JWgGsPB5qeIjs0
2yFgF2mKNHRCwTWWzuoLJwkNV3A/WxZMi0jE0hsQ9Z7WZN0NQugDbUBs5EO1oRt6fwdt553iNAIr
T3h5eFCwRT0bZc5bf4f08ab0LKzFiSk2QMRx/Elmr6FacusWEUBJUsdvowB34Kjk62Nb7+iLkdgr
OhLwdVp2VrODAUSyeh2/dkiEy7txoWEqpRz9k8xoGUsioN5MEHZg96eBKDxl/PnRH31Q5CTtqnMv
5OoJ5svTN/IAXmQCvhVQj5O3AF86ODJbbiH3E72JqFS9M0LlgGJexqsqmXU/qODdV/D+HUfPZA+r
CNBSyx0bZt7+60Gjd1bii3Cnr8viDQk096OlPzKMZmzKYrIYrYBjgPUhrKpAdmlWT8lhLUhwQJ8o
BQ7JFSyoE15vyp3X98oc8lpdl+l77uEg8sYKcWz/bta7P8+GQ5twXYNXCVUdODecyogR3411iChc
F3KGIPVJN3QAS0VGNL0r9g3wPmrhYPwSQOCVgOESXCPxr2IJvBuvO0iyT8b3V5Ax7pn/A9upcwLb
GOUXGvqoExbG99DQc16Et5iiXmeg9A/iPnuHRsUizpwCLYyQns3Qtcs1WVvw8y3x3uVEdxyHtnv2
wsfQraQbrhBkrDCxvljhkWu9gQV8RBNzL61Dc0AoYBJSqKB0Dn6uCIfuZn124dGJQ5cpLt0/nUV8
fCnXuI+Iw6Q2PUdZxpzne4/zzW5F1cVRPQp6QzBh5WGVYNNdw3swO7+7ojHLO/az9JB7RSsanDum
xKy2r+FUC3MAazQSGSpaEw87lIrStZbLJmknmYKBpxZg9y8FtSMI18ikN8m52aF8cWOWrfDWjSlF
LfoP8IaudFYS6UTEbDhyBcJehzQsf6W4exOAXcynu4ZyWrobsRtQQMXIP7auOAgZNxOzmeLVQMkK
SU1i+vWhrxJGHZjPpov8iAJfYeBdtCPA3Fb/j5hUNlP75sR25Lhdp2POXtE+DxhyVJytSNaqgVbM
UoiUPAjFjaezBF9iu7CEjxFlhvBV7YmIPidOoj9nPXTNDYZf3eWGayQObEAY0vuVwj0R00RvOk1n
OZ5SXieR3e8jv1yz+TL/Jlk8vMaody/2aOwUgSdfsRztu2oSkjN1l9a7D2gfDDQdHegsLNAXkgiJ
uamBUOM0hOhDQPwS/7n27oGl2thZZjeeZp5rHzmEMYPXwodh5jSXH3e/IedqNqZfE43ekQlAdkT0
MXXeoIVyDPA8radqudhoFGsLvf5NG6tqO0YdByfu1wWvcTyhtcoqZH68NthYOLxkj2HHNR9X2xb/
D2t4/Dn1/eHwAyvKIspNJfLwidVBG8vQKpN8icffVj1cw9WOHXN4TSucKI9wwYXOdXfy5Fnaoplf
MVgUIjZ9t2K8cqurxF9qmbCg8Zx0OAKR2dqnk8LiNmd2IcdeQpxI5obD0YS9a2CcH/wYV+pVEa2u
sSwgvWCQWz3wmtsjtEwDcAciN1qyb566CQtOiYaFxH7jz9NwMSSVVlfOY4kelfdLpx3P5JcDQETT
z3P60jm91y6dEgkU2IxXv8VetLnqrNAK8rquPtGYe9RKjBDqx0j8G+O9vMoborUm8xdsISZNga93
xPyVDgd1X7uyqp9VysLT5YnyDUfDJNLpitCuPby9nBcaJv+79bLRyd6EMgXQNLuhN8nNELkNsPrn
KFMzLBFUENLgXcxNGGDZPNMI2zGIDevJ6S51lAZgB0BAL+mex+BDxsfJ+WXBipuKFjVJaLavi6Hu
yeozrmonkudlD7H+/ucZRcJFXKGdBrwKxhYeav/yGx1cxIK8ag7T5M6UpMMTevcCA1cj1lTpWXZm
wWTnq0wDIRXyab3Q6iCkJqDu+LSpqLBTzawWoL+o6Bf+4p6jdOv9u6dcj+7O7PvUDQSJP9hysbmn
Tk1uL7ndP2Jfs0IYw1WoMyIXGHEN+DNWXSTma0ACZkbHweQQHlzUGaR37b7w+uz2Re3UAqbEho6L
VnQQRhjLkj1GkdhwGxZtb9KXzGq5IzyLr3rA6fA3HRCJP+xomrh43VmlhMAzZIgjbQ+4kUfc3LzZ
MM85hiz8bmvrnPdoNR13p0zc2zDmw8qEx21RKRhi0UjshuF2eFL69Yt7w67Qh+d+m2rXc2X8W3i3
kELhVtXVMLzeNFYd8ry9xZ6pKIxgyNdgWTeHOb1PrR35xNeuEN9W9WtEwyedQEjB1O4XMF1RifmH
mFUxBWc5+RG6vRNZbg+W11zmquyhC9vNOlsHsMK380Z8IY3Ofgm3F7ydHuK/635KDIQvmY/JwLmn
PygnndGbn9a/kYdd8oBFTapdSOQx+xHr8jnl/VJH2fGgTyRquqUafJFbp9Om4EwIoiBY/ygd9b9T
U5EIEtrX/R/SDTwXeAFsDWhMU5WBfSocVIyppS0XSIi7kxruUtGikNGhE6DxFHL/9UWwpWQeM1Yx
BMyFSsPvFvfxUYlKQPM7SImp3Ob5ySayTJtKJU7WN5jYF3pMzqJt3CHdW4SD9Yfhqe10Kdx3Q9a4
UjIEmSmrCw7Vv/Ls4WRly2Lfj476Dusyn40v9T2Y2T0sBhjqE++sBEeoWiBccFEnrNpX6CyfqdRc
cLpLiiVibvkJQ6UDi3cSWKfG4x6qolKm69bCjIPkoLljuf0XZdMCUI6E4ZTbb4iw2fjYF5MDIeXC
6MhvsvP6nq5HE/1uYxF/CoXqxMgLDT8XJ2p+fbfjFtw3R9HTCnpKZ7jY65KSMnjhr2Ynpo25gJGK
LfMTKF6DZsB98BaUE4ET042fJRbsLTTKXDmffCJxjaTiY7PNItzD4EzDe1QX9bjUkWmZ3RJJlBi6
5Wyz5BF83IjiIC0suPdUssra1OKw43BUNXK5zN+bkdAELFt3hz9N/XHgFl607jH8v1EQV5ry1sxT
WONEqWF31QjB2rHw1rKhoJJ6UThxf1HP3v5y2Rdj2Flh1ChrAJ3MkwHlucm2+tAvyFvAiD3daZ4A
2eKWvV2o2SyfYe9ea6w7Xxe1II79WMR3p2h8AS5Om6MBtZtEcCZvByG6JByU8LUDuwNEfh/KV65q
86wUaRa6bcLeT0EhIbJ5ZEU1452+SkcRwt65hQDMcd847ujlPD2MYOE6g9JvZU8oP8KC1US0JHjc
KgZoQF7MSBDj8R0i6DXjHmsLxaFQT5Nk4CfhgOoeGVEe+RWIqEorzNOxSLBtV5jnr+JSlDCrGvwB
s6ve/A8Ab740X1lcZ8xehoIpspwOC1CXbO/hO2SJg7LHrTpLJHQ8u+6x3NGl05XmIs8sp5hYlCk+
Ic1CG1isz1CvXuJQWm9RpQ6diqINDJR0YI5hr4C3LhaWtT71tAZoKHVZu7CtbuHGadcV0EfVYwPW
9mIQ7EOUfB/GzgDAYXX4qfGj3preq5b/0A33JBHMKNQLiDSmNwJAPbE6sc30xqd74JcJe9KSlmel
/3CN7jOcJ+ChiLfVP9usUfioZ7ZexYkSG0/ZQZvmXayMv5Pnx7eBQrsAebal/xeDO/NdsO+Ebl5O
2L7JTR15eL0gRkjvUQyRpbueGjzMNaJc4leMVe1wLIJ2OpKXTaz1QvPZ6FBNSWUn5qHBB/z9nJJ2
/gDo2mvif3XBGQpCqKVWONWrDQGfxNzMNhrdTtdQaz1ck4gOO8jiy5iBii5HJTqlFN7Hym1+Uqc/
y5MLAumHeItNVgK6eai3zTHn1JMVkSdcALxaa6eZhLHa1muDHNm+Owgc/wJCZ8ALhJ6LvnIl5Zxw
z7X0tOiNwvizWmaarsQ56p52LyuNrbMIpKUnP6Yud0jGP7qPFA+Z1hkxjSAij18ikFupqi+Q++gF
wqs5tpBQ0PfsWvlUVY7rLnBUTje4T5giy5p2CBaI4c46UUKenNLNR+N3XRDIS05I4MTC3LgQtn1a
yVi6PC86tMU85Ews/HwseZCTadONXv0xhQF3Q4dzt1yy8xBRrJri72xWNrcS/0hK7cooimgnak5P
mB2IYJcUu5b6mtjAeC7PA4hGV8R5j1fLO4AdJbtrbrPJK4gBXDocPGO3KnAlaBTroli3fa5CeMt7
IxbOLsRLkFiYvtjVYRAmb0KUP4T/Aghbb4h3hcb8Fr3SPov1sBKRhO+z6zDUo78U+8+myhllNLB9
g9dGWsaduB3VTncq8HIUlgBAi1gCbTRAMXnYWqISZMVTwTrNYSBWOlegbCNTesy9+VfoJmXlLHMx
LaJy0XDaizK9yDqNnc/pe+F2532AnjgWgVW61avacSW7518NYEY9COm1bWvaHINBuPFfWLANBxN3
XzsUgBVwgw+X0kxTB/hM2ENcyn0uEp/ORFw70a2AlwdTxTOcWz9NR0BdPnhEZaSd/feqNLoTFJ6Z
VQQnddVRdkGmd3SfoW7Y+YDP9/nhOa1W5uzFMyleRk8aQ+UrUyfHLAZcqFncWN5nZp6RWPHhDb8Z
uqiCeYNSqPUA/Pca8NDiubCAV1DXnamx1OPBCRvo0o383LNVdis1SCHQtAniuybKpc+DL0RCBVb2
9nf35yTvIV75ns6HB1Xwv0YbFupHPndsvhLhaVlRGhovyQwre5NhU5kCJF1IZleX440sxq6lubOq
uYEVF/FHIRvNgZftMadmsKXEABgcbeSyuZQ3iHldodxjFRXn+5R5Ej81xWvkfmHYZ0ZDjcw3ReNp
3YnWs+gwEtm/Pi4JOzqp68sWlvMAccETc6wFArEXNSA/YuzVnBc5HPBRJ5DS1nMUREItW1luHOsi
LumhrWMV/ps5SUg448J0wcXfjkhZ302nU2kH0OTMby1V820dCfTdxHDJdpQ4Fg0m3LLcZpSQN6VC
2Bg0isdhJ4aCbI0Bds6qS74ciL8NUBsYRTTJngPBskkaRn6CFv2uiCCVeQzu6ZLxoGftRYGe0bhv
REizErcCWKSVr4UgNWpY7qHCVLkPBtndIx3X0vCxa/zZffG6HOkMdTCLIVkM0xoYkZyIt3Q1WbwC
CtMRskjAJ9eO5jhAWfN8sxNEvnDGaBonwVQgf0hYr7QHy6hcP409Mf12UpJi5BULp4O5nkRP7UZu
v6u/rYzWqTI2OcK6JCr40yZoHTYYQRjj37aGi3UVJZIDmPzKLyai/vKAY4kK4G+BdSdBmEDE5jZ7
F5aGQzD/Tsk14Qv2L3oZwwoP4aAS81Kh+h8yZ7ClqjeD4nYxq0A0IyU3w5g7BZ5dh9pvIhBZ4VwB
pZEt6JW+1SmvEWx2DwWK6TDMlQnebd/O/gzvfU2RP8GS/K1vM7Gu1oJyLX4sXyEqLRN0KgLwBWkh
6xtucVQEA3R/VynChKsvsWrXVd2idXFvlyD6qFQFQDCGyBgrP0ccZUJCUgO035kR9cMR/I/j42D8
u5fOy9K17oiSyM4L7EuQiUz7UtXRW6K8NUEc9eYkMKnPNlZg93OoFf1SZ1iGa7NBuI3DXaLimx4C
RM1nMwM0q8lDjCv2b56QsXdpthaiVFQsq7rSa0AsYEV/CdEXnwl+XxbKsGTiUNMxBBY43r/HYwv7
kroWRWSGlD2pB8bbVTsWCJGz+dM9YrxCi/TInoSLoWvGut0gvaOnzPP7R5NNFnCg8z2ke7kqbfGa
IhSVrgopE99eHXEcrp8ytUgrLZIkq5omg8/iCWX4KeCFZ7PFgxuToecX1i9fM3P+L+k5F9LKH2nJ
YadHo6vUIofr4tonajbHkSLQ1URJeeFvHSpCBGr4aJSY1Av1K9skwokuqDBVp8o46w8K5IApTJjk
TVparKGYtn1jaof4pG48+/EGdP8u2XlMt1Aa8v3Lf9ji9lukqBmD+TmjlZ4wRhP02Z1085lnQXRw
WWG0ZhoefOucKrozPF3Eqk6oL3T6i2PUOL0dZKqftEhYmKF9+xS+teTT9o2fukCkPdW8Sd0HJV6A
FU6CFG664xY07EHimWSnNk8D38ntMbBvMh5x44c3SZ+67ORNq0ErJ9ZjcKOLPvgtALqfwxgCy6Mz
0ggpAG3jPINUKG5KPYw2+0MjAtzNXXSWmRaoKZjQCVmWjCcvsH+qJvEkYPJAZAR0MDzY7L/Taix3
2onlwrllgchJvZfjuGpri5odTuMND3Kt2ncnNk4c/ZExPXnY+VjI8MTig8qVxPAv1YrQSAmuYzMb
8x3HPSXr1dfgafjQN0Y6uMKz4d2731o1EDxHSZUXW77AKJ8H//tb1ucEQZHSM71uWbcu5Q8/D6xK
PmnSq/Z0jElKPNpdlMFmNd1b/rUjZxeEK/MTa5wTtMyL3acAnm/kEL5yobgnf/Ops+wOumHAo5Vo
RhDXD2jwAYzqSO11XJxAp+aQwsxzeOoPj3JEk2JH0rSzEvizAxir9WHdOe3aoGvr0f1OeX6vl6yu
PhLHjnAZ6FT5KGeBwiW+pLfdYjFFZrAj9ehMyE/z+IFMvDJLB5sRJ1SzZn3wv2ZKrBdrbslAadW0
nOOOZtDHfO3PhkDQhsc8cbc0YmRP+ZV1i/gbdeLe+HwuJTu6BpHDOexCOtc4QtLFWB0C8SIPkwA+
jCSKykYU6sHke4A0hnpbgI229PLNnmW8eMJuT+EpJ30fGbFAtZrfRO6rwyHgI0m+UQMrzZgNaUy2
/7hFGYRRM3G9bkmDDKSgLTHG/xNaKf3dtjzljxZ8HjzA3xm/OLJRd+9TRgL0NkmPtrOdZzigIv3S
DFNH+P8FpOgi3vOhE9LmWf42H1O1qIWYoNT22lcRKDC3eXvrnKgGSgvrRLFbuD0s9OmVmDvpHpOh
7Wy5QrhT9A3hH56+oMubR3rYxML4K29/TBX711mXkwY6bh3whVkfZvmlVCPQcxmClgxhoKaqEFuK
qv2h54uVqK5i+sukDW0fZB/89NBjHZkdgBZKr6i07DLHIZhWG0xcs8iQc8nHrwE/ZT5VLbmnC299
wT7eHQ3S804b5UyLKP+HoNK7z7NvKrERtzJ6hlAPL5UsULzrPWyXwX/9ZtZEdS+gVnk7jgso9FMo
haZCECs4Pu/uxYczCJuvXjSmT6BWs2rguVBqrF/eetUvLfjwJznJyC6MJicynB86AlpFejbQKK+q
7NzN03eAdZwVe5bYqgvUHxqDrGcdZOZJ2UgISJGyduXtn8bb1FPAx66Kpd2XfBUZs8STu/ACwsCi
lAo59FwJeEue2j4BGbY3MnlQiI2Qg+7FyWvfUkS8LbJITmwulqAlzi8mnH9k9MaSsBFv4/FWZujZ
hBeZo5Y3JuO7w2A0oHJv6mQvbvFqMQwKXG5osSDQcF4CmmgEr7C+1ZndntvaWeqg5HUukhGwelH5
TRhVaz8fpsioUB8TEhuIYGhDytdrPae2nFscpnLyvDlYKsxOXvY38tf8twswx4SQaskgoFUKMGnk
OqWWW7Be8dl2lWCwWWjAUS2UdwomwZX7BQxIVwRmTWhDjDBwFYXPIhLCu5qs3QmS4SuYQX4WZnoz
4z7M8S6VUQINZyKj/SEZQP74opW9xCLwa8VlMCNhwySe6XBlY1bq6eiEs+ABrvnh1xGgWYL0bLd/
Jtk9f0ST8I+KOxuY52gGPz1j37bG8v2vA3dvV7wrsm5zB3j4+NQDktADIB2f3V3RwCbfUCsvc27Q
DczJotZB4n45h+OCwBXpuvbYU9heBgPZLUgNSQ3j9eaBt1llVFN0RrKIZkulROxK7cpjMPiu5rPR
HI85HEn087zlLWwn/Y/Zu+/zEfPyLl0JDWziLpC61dBn0qfcR3zYsP5souuMYq+MaFPqdic2dS4H
qhBOPdXCJEM4GkEdRO3xB+xaCco3BeaN01wdtNg6yHo66e9QRl913D9nj2/FgBIVNPgiVEvEFSZQ
2M2vtya1RFVq7LWrT4UDZZeu/CycOsLwAge7lVbJcrb8Bbr+82d4mhYZ5x3utV/87GjfBP/0Gwqg
dz28xQVzG++H4a8GxdqD2m6l8qxAb9ZBAoGDrYKUxgprJhxfqXfLmiVXCAtpTehGDJf/F2O2hQq6
n585TekPN9N+udUk9fg2L6CYdB8Oo/SioUTL4HMnG1hkI4qHpoRUEnXJl4w+u6ZCGoDv2tLK/MVc
VJMJC1CrRoHZjseYNvAh95u4Nnnz7nHbbPvzg8KSiKfypFhSOu6TvrXzpAJ5CNubBCvI1lzxOd/B
A4ygPAu58NFJ+nYqiFK3e527EK37/0pHwhqzl74UoXRo8SRXa8Qr/E0HZUgubi9EbvSe4sAqcjLY
BxQ2SUlGmH3RVWh+BaqAxkX9LicSLMa5pON5AaSgtXqgzZLtTsBPeC++gENEvjwFPXG/DWqBbNJ+
LHNINKgGTg2svNUCX6fFkyOn8fBwAa1g16ISOWpO36GqATXTeCeOJ1PXFe3F6J4mAWslskiPsNA2
VcHzRl0JLzUN3/gPyktRS8aABafo4xGFTWQfCk0iBg33QTR6Axi4kOMxdscKn1aIGIqOFBY/ic/r
2xsP4vDwx2kR6HeuvFO72dxmOMk0mTgCECOM3JUegUGISwg8Emk7DDUnJAvgq5caczzAqaqk4P9A
sjuNvQZYjiN6V9dPFRaM6vGUvfXqDvsevOZagaSWsjXAekSQ5tJ33ur85Ly2gF2kQ8NCJBJmnqfH
TYbBBf05kMvF9Fbt+ESfD+aTi1vMI4jEpC+R4Ce3tF9WJ4SZLZiePR8KaPyVNel2JNG/2EqSDzcZ
bdXlSdM56QRf/RDuRpCkxIVTdmEyM0Aicvj4rJXTl1IEiqYUlXkdaUdHTGU8xZUbF4QbVF7DyiaI
MkQixGFSMSpwKwANGffbEoYZY+UYfkPlMr+RgYasRseW0d3U2XBzE9DOCyJXLRn0fMIPjq9YRaid
luRrQyneOXSqhuQDt8R6XyYt0iGr5uMSjTJGs2jCU1QB/j3o8De5ymTxDaC2j2Qe1grxNqw3e5Po
W+S+FKyTKCLVVIEG4PJa7fW2cShEBWO1kBgHEYNDiKt+5Y15EANZgXRC40uVw2v5SGplk8nvE0dq
ihQIq5n66yxbHNgtKON2yzVPS8H4GhldZleHPupsE4bo3y0HDUX7IkR1Moo4GN+ZVMH51rc5ufKE
AFHMMhjuUg62EzHz1H5SnMIoxZC8PviQIIGhZmREVG7NfVnrpIF/LoT31FGCvx4vh5pAp/Ih7Wlg
S1PEZPzaNaSAW6FHmWE8D+cZowOb0+qBlwDo9rT00anim0vHBxPz9ZMqG417NE//7Gs3w+kHK+TJ
fH0YRs9OV2DBtypz7cVi7XQdSGIAFgc74XKr0PDu4EIPElJ6wMUFZt3ncpItI8sbwWl+x+0B/MGb
CSWWOQ1IVCxsLDvLuTCyL4cB9fl3TBmAWn7DyRhk7SqPRZ2kNqrtiJFuDvPKVVsvb4uquD9KJN8b
cAmank3q2ibNhZWIKYo+2GEnekLzKWM8BMsxp/HbbPKfDC6vPr22BaPsnbng3bnFULsQMBRNGaoY
CmJSsp1SlIjxVwD6jhvzvyCLXhOFvgTOD3miTgXVCh7u6q+zfThTssczmnnrfxRmYJZKlfvhQS43
57HHKH0qVrj85Q3l6fjHWhd8DFnc8h2UAubmZNnNSNpWRhkP/DMISLd7fCSARaUQtBk4S63bqiYJ
fvoNo9KHXBjqRWJ/HNI+g0lOePQCLiEC/6s2Jctg2ELZP3jXsQTgxAWHLJp6DHAlVRev2+CNZad8
oqIjTYcam4I9arvVnXTdvKTzUFrwm5T/N/dwGrY87bNXYFISdr6NpwnTfpETxXt/4QWoZOEisQmE
uRy3VWkxjUijFyRxsvuI1yhBQeoFwcl2P4lIryi7pc1i13a+J4VmBeRtBSp7dY6j5LBE6ZOff6Ku
m1I+kL/O6FjaPn9Mv5klHt85tKEZTYpp67I8dk13D2uyzoTQUsVI9gSZtwGzy28gBP8sN+zA2b/g
uejTxBgTgirK2+x4zLGLdtETQb4jyVEHAg8EyjjK0EqYGDzGfw8ghl6e0mSxKIbyXHhJrndKOXFQ
WMMS6OMbL4yQr7q/+fEQT/NXB4sOM/YDyPATCtIjp2g2LINFrearFysfB9aYwpuD8gsg+zVO0VZU
outjPceTtAAXOklbx5Fmg/7jfQRgxK2+5Pwmb48lG+YsKWR5CjbMk8MyT6zvmjCFMTPj1sbS8YZ1
BVqp7WzPHuvUYsvmUe3GLmwkEGilX535v8tNd5xUA2LziLu6TLjTPUIpll+OS1/jCz8D3DMUR/hn
WMXF4vgTNGCzPYZ9hLtTQAhlSEA1hsOr+WzATs3vvf2LU6ojdNW5GTiMS4D6MQ4nJOLAt+FxdfUy
uKHTZe9wIUd9vfNUdvEIKDXdnVBMJhXr/Y6KSVhAnTBpOAjLuX83aSZYWcu4yZ/Ycm7KC3wnEUys
Bk54lWAFPDL7SnG6GKmvIxA8RikXp/31N2/FVktfAHkPlPaAAzz+4ZQDB7nirc+OjD8kvFUzK73d
Kd9mB11fn9Qr70e3a9Go5mEP8umCq6SFnH+HsOZPmhE/9WlchtrCfUAuzmKHfj/b3RdqhkTylng3
cGbyjSCjhzTwF85LNuiWxAUu6yJ3F9lc4JQWlaL1nFnmhMlBiQu3Hcr/kXab02HNasNkpvb2naTW
/bb/njD7t8+jGe9gLN2s9DcXIzN+9UM8dmZu58nQ4DrTm4pjVdEwvRjyVOfEEW0HC4U+jg0r2kHS
7xiicZVviD6dLkbMWlWSs4+LfwZbVIeXERoFIMTak+GSkhz372g/Q1O8fEurl4ZAgrEUIrR2Lgqu
SQBgsJCxLCl41WJYU/5Zi0kaWQyZf30+lxs76uUkjKHhOwPzrq7l0txUc46/mV3B6grCgF2+Nk7o
Plzi5Vf4KdS82a+3cSjwwTljrjriZAk/YTCh/CTcHNhh1V/FF7J1tHNN6Y88pUisUTcGxVNZjQ10
OjduG72L4v5pOhza9S0ky3J2VotUAyqL1gnhWmvJGjOakxkBotx2dhDfurigzOfxxlHMAExsB0M1
a4/QEFpNv4v/2k6Un5XYnFF9DhOHpt06n/cXbHNq2i1tVS/o805JojYSrBinHGW62iEQd/znuhKc
YGuKkzWAPHGYMI7N8tphJzeS0JOcvUQHApB6hbvOQH5XSJ6ye7oYUg96co1+QLwTP8x1c6WQksq2
QMGAQsDmiohScR2jQrjdY/EeHpQYuFin8GhkAEToH4l1GH9akP5zTcsmJkybPceq1PxYHW3jorpp
sAcpzmbaO56UklmsycQpDGHxpUffsttrmu+wqEuPeDRrxaQd+Epzjo7u/iYdf/kMCDYb2b3lFCNW
6UhSIUNTOH6InsCJUEWCe3Qy6klvDmHORk+et6ELbwM6Dy2y+PBEtvv/GtC/DEPYB7SGeAB4EqJD
lCx6PcEhiyebAjl8+yDJBRnGlzLVE2NK/pvzoySiuJwD+wNoGau20ow2xEetLyHEJMmH4oiQOW9X
uGFiZS/Jxe5eJ3mNxzWgi9OD5dQDNvqp60N3Uv7oz3WkchlyeDIRbKgOBf+iEB1dZ0FQfHmHQdOR
ZmMfdzd+5S5kQ0BZlYDQEEaA3/6+UxRHP9aVPL8/7CppM8W6gv2L/CGT0UPFx2Gv1zsFFxmOGoAQ
IjcabvdnIN5o7VXojC59kpoo+CPr1yjoWo4SV8aC3pTONZBkang9FhwoAW6srAURjWuKtNOS1lrD
D6yvrvlQDhReZ7j/39swdSNcjG0cJU6fYg/zVIktUfdhyOKYF/ic8M+/IXYM8C+3MI4eQSwgpUSE
AOn9HqB5WkjX225djjiZlgIwJrQSn5iK5UbfH44ameu2Y5gNZ/oly81Wp+WYVRrMQLU1ZUQ0OVXY
q1XhxUHHTfeHNR0nvCsIjAhYt3mOYn5yG0HYbkS9Aa0PmgVSPwH101Wt2KVIiHsiyHWAh3zPwG8s
n39ntEGW7nFnFVLV64/6mA2Gt3RjOozoQp78wlngEP9cfG4YYspItyYgtaiZWqfISM81YuVItpUx
VV0O0g6yZMKNlUTNo6P9tWhvwTwJMPmO6NiMTpsETc5PYID/n/sc+LSp92B7YTBihQqHGozslH+5
2F9tJkJ1TgccMYzWRxSPgwq2obQViyZmaMRR+iSze4kwE0Gp63+VEO0qYDgQAW5VFEsAe8fD1Uw/
hMP0tetUUcGQ/ehENfWi/PskjLId6rUgluafUEXWm4Ib8oPpDNR6SAzic9c7snzb/P3HHzeHksNn
zvP+QaU4xRT8dukD+6wXSwvdBPSpO2rDbas10BlFz+9AcvtoJfSWphoYOhgo20A8Wvq+vSGVjhGd
BmBMMQT1M54rIw2n41P9n4frvVuIbxyP8J52nVuq1GKh5ts4LpU66fYpriApUL1sRiihNb+nLVIC
/9mQh9qiVvE+gEZ4BlY2Mj615eoxK7efVEgBEAyeW/W1rxuat5dnlSQFYu/cGrlms0xMus9tRKiS
cmqNzr758lbWgS7dHop56AbZMOlyiIhK+IymxeRwcUjDPpKBJVt4vcVNttJSQVKOjV/4JuYTbcbB
fch4yL6WX22DnO2F+LfAm+ypfcLjSH/4GRwZqhUOJn4S8X0X6bSoXMGsrja286X/4vuCWugxNSkw
pcpFUnDKt0KSEN+YLN6qrDvCdSWrRB/NEc25PkD644df8DPFNCyweaelaphyaODw8eXCtZjbkJ3R
gG7nJpwPi9csb+MxjWyqq3NCYIm95MK73Q2IN2kENmQFd4OWhSwvh1efLmVv4Gtz/FZcXu61/yro
sngkOUDBadseCnpQMY3i6oB84/BSrk2XP0eEit30fs49W9OYGx914GWRqvXNO4wzIK552K5JlK5q
YLvQTaeGd8XEdD4FWSUfOuyVcyOHiCCnBmYTfEOj2+3j5AbEDms41sNP07iYQDfaLrJCIwHGwQos
TR0fOGzZBTazpatGtvDe/aGZbKowV2xHzZlCFSw+/U3fN+dX+g23P5SLGwVC8lqRR7D5zfMbYpVW
n8eQO01Kue17VNZjumtm7QuVmn/aEBfLDmfixRcGVY3/VY85Of6+QFPjH06TRFeK1KK/oDrSFYXm
Drp0nccGLj0pfFJcDiQ2mROwCSuCxdeUhRrUxqBwPotNn4CmwYZgeof7VDWFrTpPgGPBR7dmnCkR
EpJ4yAnh//FBMl63mh1ap7dfVGLZ8FTKumnzUftwwHB9oAMP9q36Y6reKLP8IWSwBHsynNQo5D0C
p5yEsyuD74tXnMvmFaTk369vB8n9nBovNWUvKfu4RDDQx0PggXl+aa+5J/nGVRsvm6/gLYzhdvl0
WappxOidpCTQVmxsY3WilHWEgSSqutM3R/l8Bom7z1WC1dqA8GrRVqwD4hqrIe9y0mTHtCKD4jc8
hCrXXOqI3dZZ6FgQK0in3AooubzeURZy8AwR9NSSV/2IvyJS/QdH+35NSJgUU2kSW2pdSQuq0GEq
ZvwmmhImE5pvEtosU4M8Z3ObPl35iSPLUHo/Lz3OtHUcOLNldRvWAlgkmdb9Czqxg7hlC+Bzk4Pr
hnjZihaKl8u9dYqTRoWOsiC2nQXOSOQ2FcuZKu9Nzg5CzdkSsKUarGZgu9VQwCrjwDU12tx990Fe
zT37ujgLl+hfr3phDMmVe0FWQhkc20XiRlpY+0MEPLQiYYw1q3/3lUoF0bbhGnQT9KmZ8RUyj0VD
yo90HlrVbeEk5rCqt/JaL2WawdBGoWKiJAz42vK1Q54vTw4WEFihUN+JUeOkdXeXlMX63QWwbnMU
tZLC4KGrbipX7txOEMXJWlo+Fii+oZL0wLVzj+jSS0bPTB5x4eSk24ndf84jGWPLGoX5EPP7eRw8
T0Po4L6kf7IKmWOlApDNLIYhSzStoKMAYP+LkGN2VBrBcMxHVY/lno9AepWv3eFnIOIl8IinPPYY
j82Pqz/sDw6dFKY1vHvQAFv7ZLigD2rxLTi+Uqr/ywMkLdxVZUknH8rRI9kXJjKbDHva0dKU780K
jAH6GxmTQ45PLaBtVTDtHWaKpN1FFN8FsGu3G1NgODP8oVAYahROgMz6NzTt9SlzAWcQgohTjjAG
RSd/ljSJci2pm//2c5H8Wis+dpo73Bwj1m4zr1ks3vjCNxhDonryX6JNOA7tZdAtWxtrdZyUTCw1
XKsbB4CR4VPlUB/a+0+zCS9GQK2qrb4AyEJzJDh0vkAGb226MqaXNhMNRT2VWO0uL8+E/+0V6WC3
EQaNM8i4KmHQIMynmYCz0NqsNEs27Y09781FUYHbIwC6APgvBMc5n6M/P8aBxiU3YQ32KuzldMhF
+MOr/kXVXybxm5CnkKhTuuhwcz14UUYzcpxToSTDUwScXGQnREe1f6ka0mcCEqn4LbF9rU2Ehm6A
3Ioq3VRl2blQ8pZ098yUkzhPddHcNKfm0qRm5jjM5rJzxTbUX++forq4K7zc7cljDGgBCvtMKb+0
Bpwyn/6209s6CDqlOJWbwcyywsV+MeHk9jB9dasBrdnJ0Nrpn7fFUxk1Rvm0RaInB+G71vSwlBVo
iO4CtdcOV3c4p2gimsm7zRlK9JMhUuFbUnCyVPqeyhce+fKuKGNt7JLdlqgHRaKm5Gn5st3TQ4Fq
FLi7kTDObYrreZtxm7ulJXUP0N17kOI0abrmoHxn+DBCDjvouQ6fQPweBgFP3YfRwQE+am0qwSD+
hP7lTt3obIRBwjkkY4idQbN6lDwUSL1GNXETb6/V7b4MDp1MlkjYVNUkQga+hlUtsVcUisH1lZ1m
aXwa2rxeLGyZv/y/5C0okX/XTJg7yZI0GfCxu478DB9tBKi7VHuFCv4g4VxpJ2O9A0KPxRlLIjcd
JLDb1hd5oNGB3MAjQbvtkj5eB+1gLUra4/ceM6S5c1LmAFw9p0M3tl+hysCGg8E6wNdQ4jShV+sd
yNZwC/bzaWh9T/gFtfeK7Wa0yCG1/3Mv5xNK9zIF6XbMp031OMu6RuzhOcq7Cg+wnOEcW0uavokf
W7tXDLohxKqHNVsJiFOQMmOPRevWYvPGPngYkZSFii71L6wTlld2BpypyiCBlrmly+Gpcd0fVnpE
10wL+p9IGvP/qz7+BriYzD8zZfqoy/mnMnQ/v1EDeEHnwwjQPwQHpk0+kejod8TnJzqtDiP2g49P
9cbcKxOfT0+Zrsa6V135hegg7j0WmDCl92Rn6G9NlMEfAiO/7KsTLmIfGg02pJ6Vce525i2dvl7v
iMB6DGMrTo3OGf6SG7dtRfBKhjFnUwhRcq3tenuKiH5zYPys79EefAMh1pKUam0Ou7BoDWeKvCLy
QQq3/D9AILrQKhibcBisK2ZeDcHVuNOWxrwYvN5QkhOdGPdcUWEv4mLSlqOOIgfilrcwEwtGJnUx
vz9znVwu/UdtJw0hGmFv5CVeGjxSqXiPkLUcx2/F+/sJ/F4UgUHnkKvJtivhPNdOSZe1URp/n33b
vFXmoovpgXPRiYw3yjr5qCTzLxOAesQLi99iq3PeTiqbRg5PzqfHrNNlOoCTUvXaZluZIfVdzHRF
qNqlgdWIUVubBc55ANDTyW5xGOyfns7eeKCtbhf4gPboMgoPW60ZlnupAGSz38Nq0WwS4LK7dw1C
ueTEq0TriFWG/h9kOSOCyb17VzvbMwjZNqLJSLbnGl7igdCU/8Smhogc3FuKIiJ9eOC0q3v1SUNa
MOUlymp46Y9q/lW/hdMhUzaEo9s1QXylhwMICvZV0qDiMFiQYStlNx16AtweFTV8Q92+1T+oJlrN
bAdOFlIO1nIG6uWVm0qGDnBFj91yFVvg7CXXtrcsD3ONfW9OR0+yIu/z6w2A05i3ZoaTZEAjPGG+
v3VlKJzAU+mAxKY+rzpuPKn6zGcdEPbM6pcMNux2d6LGAhrYXLIjLQVWXUeqG0oXBsIBDi3e8CFQ
MuKa8ougbTQRE5yNfYIldkJ2EeP9oKEM7zBICIt8Y44sBjWU9J+4zyBESuI//+vOM5K997zJjyKy
PPD7gXCFOsPEiVApNLp5FFZ7kBU5S0q07d4uuIVO8ubj+3eTWdaiddQWbNBwQQcCvoBBP2CMXZvO
pdI9ptU9FAvnAdcSPB9MQNcwaB0FFR/qFKuXEMZOoqAVpd6z6K2V0nGinE0r4QX1vxLrebm6biTT
6pwLLZv+w52M9PWy5FqO56Gcsrb4SM5fiS7xTw2Qqwjsk6jLCI2jMH16c4xni0ho8FrrFjX/B5/U
bhE0AVi6Lva2HMxJHQJtenXHuIk1cLHlixJSl3Y8WSthDHrNhHzxZVsmPDo2+IWx2ez8xni16n+n
laTT4AjTYKIC5IPiK7johm+wYs/BnkNEmtfRKX/iW4zOW+z+g1EyEK30vvccJQR+mBJlERKdmwIK
bDgz6jV1DlJPAI1sNup7NNDdBj2IEa0mTdrKKPwUIyuCflma/upQSVLPelt0zw5c1UOpqoUbS7KT
szjHgy0maiv75BCOuGemsKFnwm+Grmg2Ii1v5ujlBuURKq6ncgVDPybkvB4yfNu4f3e7io4tpH2O
CBUmU63cm3w6W8xBNpJIOLq0cDYOoUb3sqOutAm4ViFsW8dN1TF/sl/tzWxMAuAyrp7uVYBKiWye
IpZhrsJTpaip4sxiE3rkp89XiH/twP3Ga8FpQ+pA2t53Vn864Uv6WlT/Q4QdRxOIspEqDjF3C2jE
+ApomsmXgiM+1xLssidH33iWn7XEXD2BgGhYYChPG/mloP4CzeHJc2jxrWwX3eMqqtGmPZcI1z/4
8xHq+gxo3FqyESyACaNuvL2T1d1ZCf79A2+pFsZa2VkQFL5iuuCdYBig5MRUCDNKtxm4efDRBgrt
vkuF2+R1r7IehE/PBsRxf2haY8fkROI44qh6pyRZCR7x/vecNQHYhL95PVmTOw9aQNxH2w++GHcg
pvVllbMi4BFxvaKoKn97IJck/VtGVVfQJVFt1wCTtuM8EKjSa+u8lv58Bz279G26WdDGO7WM2vuf
VMrKpBeJxvS6VzIDd2rDrsC6I3rxi5cHHYue120z86aCA2j16cC9B4KD/fqVr53rd49o0AO4/B3s
GnifWrbtLidDu1oMdTwmmi1V6bRfGg5PGFEydfbmL65WEDZdh8Pi1nzENbu9PopGQGTo5hdegK7r
uxa6e30IgMFkE3FwSKDxGMFKbgEKxePG8kDQPQMNW25TXq+hYLLB7QDyEoh2TWxlqQLr3UEENeMM
noJkYU/y1oj/UqvBjL5Wo0x+zOnekadSPxxTvXhaWQqR7N/S+Z3tPO/W2t+6qf5KBnrhrBpezUoQ
58BGoEWCHN/iSVf4++CTPqVJayF6QepsX3luOs9pOPWpukeFuXi2yWaasIotP6+rT2G62/WmaFhd
L/BBjrCaFSd7z1MvEPghV/RiqwG2QfifW8S2FTEvdWxuFoel/+95UJd7r0H1z6B3O4/5uTt3SKXc
Ppv7Jhv1x0h/8FrGSnBayisqd6ZrUTpd348ZDX9ceQ624e4G9PXFcVyV+IFVpjx8EYv0KpyzhYxR
Vjj/c0NRPXpOd9Wcs2aAJsELzKA7Y0wQP1CJ31mERNrzqPDFKgzzTp2Pk/Fi45IajOHBAOwLF/3/
5XwNCoWFqDmhJXxdHmJ2b5ATofYwNvKyRTIbRueIgKRyHOFqfk/KFtCaW6PHyrFiBYRwuSD3cbgf
t+r9x9XY5AnRp63RHxTK1O0BzEOnWLgo5yvAp8EwC3miECzt/qb5hHakUEjNUSkPus9YVqU3Jhx3
2BZI+5A4xkXjaDCFwPbeE5i5GctkVtzKsI68XC4MPH1JqpfSEj3Ri7Jb1uwdIqNvrSmkrOWycWOv
A6ZZnV3BaORflNySumXcL5iwMj4r7prrwdRCBolt0jeKPumXgra7jtSZIrq4OAzMzCWH5dhLsii0
0gD/J9V/OQ4UrdiXUIrk6DDsd0moR/py7RXJm0ZyWtJlRjNdigVd04xEoUZUJAwajCodgJcBZ+zH
bSyZDYnk2OnI9vr0UfaxmUK4726HEW8A4pxVxUkD73fbavSj5Wy1v5gGdu6O+1pu+Og9HWicDd9S
gS4P/fa4LEsMW5Rl9g7HNA5NYM3MtytyXVd/4sW76RzV1WaJqh3X6wSAPG9mN5LuZAIIUBXs7NYt
XviMIZ8DFJeNqnGOppqK0re7bwPEoX/sceAhFMMHf8Fh7CvwsuNHgPSDiCnAqQgZA1nicTCvrZAy
8szUY9p1tBJMKjjA2MABAJaeUsMkX+CqZtEOkGtwjcNj9Wo7/3kyjaEHK62UP6oYMl8ONO+pcVPg
C45WEJV1rnYwen0yXK1m3CwLZ6nq19r6qq4DB82thIqZ6TV2aYIwz77/gozM/K0f1kGc4R1TFUFX
EFLVbooSueyMZavKG2swGiEXso4OS/ZUBajsrCT3ejk1MJKqQuYWhoSKsSgEiRCWjNZXVHLzL+2F
HK2XeawRQrePiTqTufBafqcZORwOAbtJ2hGtckKW08cTITHr4iQ6ZyjTWai1d9fgkRZz2+l2kZCk
docXOqYoQ3mxvOCSG3lbjop8WM2oKzHKcHmZACJjnzQ0sgBo88oYAo0jQCQazhqwQxHRSm55kNfJ
YwC/2nvItP7T5qbowt6BGEiva/kyIM6xUCJtc9dp+MDWhoZCQUYO4Q5suVIjZWJEoqVABYEtP4s/
MEwG4mUehbX8XytAGnktVMoIofNnsb58iyddgZyJMlKdn45wunU4z5Z4w0lnSFetyU3apCELsNfY
Aii3mp4ondRisTtmZfIXx+cjFUW18QLl9Ymx5i7VcfXs02MVQmYXhHqy7DeVmaxzNuT1sjp4bFmF
9kiPNyIBZTjg4cneFVBECsk+JkJtosCacDJLE0gmnipEs0u/MzPdnjW6UJMYZPSYvw60YvFfw55k
snlWGUy+2Y8R4SxmIRMSvVD+SgLv70wAPFt0V+/gMS0j5AL+ARZbQb15TLtIdoihv9CEmXmwyUOD
zHc4TJ+z8+jzyghqx1e69DpxsRQIb0C6Vsx/Iwq2K5M1D8fzYu7z9x9TZuzp3JNPgEhZ583TIA8W
Ks9fexAjm3qM0ZoPTBV/sAZVJBUO2wqemSOOKbYsuyq+e39naCwm+BDYHNcCP5SkkeVXgXLrZfmC
fi1g4ez2m6agnWljsrM8vjilQMOKz1iW7DiN2Zp4/D/0tjOZQpOoXbzcb1rbHXEq+mB5ESeIibqV
JhGrR+PEBqewu/CzKi3pWj06CZWVw84bwA/CtRCUsmSQrQva4u18dGyJThwEZ3LBPVjeqaxZzwc1
WU+aX8Gfa5rvhP5/8g79Y/5t8sb46LVdfh4DPpwD778jYdUCl+7TYTxIC/OeIuZ6yWDCCUBwlPGt
pS9VUtuWUtlavejibcq2o0UICrJqGNF/WSuPyJMLpOsAtrRGivaC1LoTjTUEk3aQxkU+GtU/ptZi
mt8u0RBqJhlvI8WdoONHFQ7fRmflii8n6QHQgZcZw4AwQB4R9iuo+xQEtdZNiZswzpMewuny8xXp
1LomzeU6ecJ/n3GovUMNJRipzTbJTUXcpzLW0rJYuw52DnLhp0gbE4PowAjWVNRWJijUGsaOPMkd
Kv/unkTOEFLnu/EUQJPham88VEY0lhgEC7i4RzagBG7g8SFIltq0FHYDu3B2F2JgIqTZEv00r2tK
wvRQCePHZ9f9PhQYws9up1VxNYWL/Db3zxTRojHBhWySTkgYIMqwsyJL1NxT3F4Wf1GwXjXB4nv7
C335zdVOrioZY3MGZstKGu96ow+KtHIx+xjiLT3cw78NpiH6goZESN5j/1PDVYGyJj/VsBNlg9Xk
I4ARcl96mZTPDINA12iQfAJsk1UqFIi4jEmKvKQ3YNhWoV2G187JJDxU7VrU+q3hZLkPQJ7PMP+z
+051+buHAMdrg3RSuCLkUf0YCYJ3HqKofUtn4ytn/uflJDbEe/prteQEup1L0qt+YiH2X+bSxz5p
1CHUSZ2N7IA0YGtjGLzmGmz7B7d5bURgynZEyXDDnEDL4Ku4PhNPW8+kGhW8mHDPv5CMMcF6QG65
0ylDl5qzSQOBUAjpXjUXqURZGbWRbzDp8LyHsio7NLIxR/DDGWOgwdeNLnTBnnfemjuG8lLZ9Xf+
2SKnzBQvFVADQvZZwe9WKxs0xCPYDQo2BFOZ10990t0JuMLK4CIhhc71fioLmY+rn+e7/UIDuibp
fFZ7V83f/MtTZraWYh0wYVB0h/k7hlBt10J/BuNy1KiiVgh5nMuQsN5KtVpJF7JWbgn57uTLNK9f
MiLDHAQFs0Y16ALWIedhZygBpZRFm/26ozRbHLxaKY3h3ZDabHGgofUoomgiCtZE4/hqfi+mXTtN
yDTSaJnjZm7Fs+9r6jaYlZmtjkV3wbAoOtqWNHqwwC71uqXL8d9hU/E0C0tzcEK+sfnDj7r5gI6g
e8KiC5g/EQGcAK8bt0uUZOTJb7GTScWngQuez+pySfJtC3Lm7ET5+1XIqwm6orikQG1Oan6Ii01e
KOFhbnxJAw+s52f1bxXIxthi4fsPhJe9Gi/hh+u70bPzFaQ5KB9Xjk3EjVyF/8BmLHkmabZh2FpM
tyjJUc0tl1wOth1q8YUn5jX0oyGlNQWh0Fwol0lVh6MaRo3bSQDT2HcYYNoBDaJtUlgkF8+gqK/c
YF1O3y4k5k85l/PqYt0FbKvItEk9UYKU/mblW6fea9FbKsdfOPX4LF8Ej/4zTRNWzYnUmzL1xnlu
7PzG9YVMdJ20i9Hjts3rtrUdoff40PXgUHf3rUM55tObHSSC3aO6H+zX7dvXbw/ucy4P3w4NCAcT
7J0w53f7q74CfGYvrv3Ctso6ih/3/5HQNVfVqoNuoawxLSmwyR8/JGu/eZrMDOAAXo7x1WN9XQ86
8Cn0R4JJ5HQm8cSMJ3u5ZgC1fWljPDu9kLCEdBWXg/wlMmBl91v9Ylc+ApGsonwOK4B7PtAnGIfc
4hCvjIZtJsUS0vK1fyMnBHHSNrE5DknxYUQRT/Wl6vmYt5PgOOM3l0kj8y82cmBE+1dbR3K8nVQf
OO34dXOt9sHfGu9BsL+1nAXvptiql6CEEYfCeSD6XEiyL3YRDxK5jYIHr/YmDW4FDKv1U8JPl1Je
YVKIF6Poo5MvE5xJqoz59O0GJKIxxKwQfGHlH+r8BjA+Q+QCvEY21h0BrXez66vkAbgSYDW9I6uv
a3V6Rcl+smmEF8jOyJ7Uq+VprGuGI4zW1ufZU+GNh7zK23AVRqybWGNJVyqEafs+uiSHxZ9nlO7Z
aPu2Q5XKI6+Dj6aU+HB3smAxQ3C2G3VIPwY7K0XVUpQrDy+RkYY3f+SfNVzMWtos+U5XwMTgPXfI
/mUHSk7ozZJAVo/C9wycLX+m8MxFpvTyb2HELFWxM9b8+VU7Ecv7BZiV/gWG3TPjdd9o5bOUoREj
TAkkwa2d7hKo+9VV1+lW1pI15gcm6kX1yY6W9yfaOBKQiwdYrePmJwjfKCam4AFTRmKZ0/yistbT
n/52O6r1NB5t1q8i5XxLgzGh6tDIsX63pu9zEI7aGovg73qDz+/XbkeJOwTJIZLkSD9KsiGJMDzT
clK456rai6IPkv0OpkNu0B6dPbt3O79bnZLD4/ZAz7DVReCNP5w6hO7vfehD4Xdig6i+JOT9BhGP
dTalByv+ekoFbIa5tMIwW6ZtyI1O4wOQW+hFpikOH7pWMiCgFsZYJE1CDx5J4HeusFGCpygnDTLk
oUiXrDf22q4Gl4QMyQvD0zrrw5K8htIkF/k8Dt6TAg6SaVSV7XcXSUvwVFNFWtHovHYkq5W5eg0s
iwLDWGS9aZTAHpuEY8FPn5QL7K9M8EsffCYigmkNJpckiyrs5M+2KN3CxhZlap0AdaG7fxDhrwXI
utKfzVPbkkVzVur1c1ecY54hfOnZ5iGUihppMEYOEyiq0SWIDmj3Hvj1S8JpUZIi6wxBegigKJ28
+4XYkAmgwzSf41410Qld8Y82Kwqi5uSz9BcKnYYXy1VSUABzjVbpVzc9AzDz7W+JKjx94oeXDqmS
Jo5YGAQ75+2SXv0c1s1DAzEnExyEMLUSv+2pzaOQrhlb5vbwcIslwfhSwZFdLQ3c7T2ER1KrPz4s
HHS363gJYv332Yejl8VuE+sKBJmNKOrNV5w8y+vRTXlw2hSyLq23v0pyYD9Iurj2NRquy3USaLhw
nBJPO+c+GeMe8uQLYxbbaz+5+n2jXdCfhzBtpXgFF33oP6Gb3wO8TsE34YcyYSOGUKDW2qlSZ6Cz
8n7gY5h9diW0Tzdp9JVUWcq+qpTchmVFh0JNp265qFgRMeM8u6f++Aag2uZsiZ0Hj8OudvYJxpos
Y5A57KZqVlqOKC1+5IkUgyzYeBP6f9v1+jWMq5PUPU2Iu58zSV/brk3j3BZtO2lG70qjlOZ6FTj/
xNB/ZqV2kQCEpKv2mzDfHIfgt5rrEOTDD7WZ0s6BC7J4o2Maw5gUqw9Kz7o7udIAuZV6QFbC/6kI
WHQWvbxX4vV02OZLc6/s1Mx8l4jDhlR/LC2HFHfIkIOYFlv9BsgF7E9Tn64nw3itFKqRBneC0McJ
w2yUFl9WVhlzpCBMGEYX0OCGd+/3vnOKPSAacsxIOuWqxhXd2BM8IT5EaMVBfZztjF04OvxPD4b9
SWuf8a4mylIXskySzD6jtnvrfr6ztC/5S4OZhYty64rTBP2KrD5GRrLIu+L8mSYb3RwoEKnGWtXT
emZP4jTayQTaARuk7OKKDDF2pl0/Fgfpf49qrQVOM8ou3U/6zT6d/GJr6RvA0N22fQ//O0dXDfkP
5Woj9qDlG9ZoPHB4c+GLWqN7KYVygl7BK0fYpCq+KW1br8HiCUZvVQ+h21CO0Of88unABbhP+x7/
S80IFX3b549k7GM4pkYd6Z2KQ4yuV9cEdTzaRmf/BgX2Hd3GX+pfUv0XMrACqU214zOwKJPBFZud
cNwTeqaEbqXvfQuZ/nwWnN0IFsEPXpp3TaAzQJSaphZsFgTAmTJsHU0avtP8iGMkklBhizuWTw3w
HJR/urhA59tgGPYZw9aDt0n/YlBu8XKTXDmmK7vsPewYjphKq/0emt7opa0ajBQWvs0o4LLO4VYK
/6x4dPafHnSI8o33Dg4/ZhpEGMkAtmej90nLhHyxzt3GDFxWlMkSpJ+3C3Vll7jr7PlYnnTWSJu1
oXU8CiEpypcuoReuL44XZCq5faO8iREvYKuIWsfsXJN/mJadIHHReay1gYJ94dZKS82X76nUWKuC
uk5iJfbkPPagKQJgqjmdRcnCiXQGw+azPpUomaidW6HdmPqKTQCyswATgIag0G7fyxgc8SuhmkhA
J0Arbzt6UvCuKOJ9nhE3ZhkWUCVkOMeLxIyxAruyU0sEXi1IT45IK2gxZV6ofq0gwX89DrgrirJH
hXxU6qfETpR9K02F/OHoACGwTcrpmLoyvVUt+tXisGW21+lKRcHHDYCLzysKHf4OlAqDF33C8pAy
4Ajxqh9LLzCxbRgbhPoe0OZJq5cV/4lrPt/xS3SxGnpAJFINGsKMxPGSAYWykqNBuciZPWCs9G1g
MvtNhdCYq9jsa8MSSheKzBKdK5z6FeS6tcDcF2lgN2d+MRgKD++okEHKV6PNgz4eiPCpz0QjULiz
PdqMVsucJXy5+Fw5v5NpgifA6DBye7lmSdBX2vPcXMAq2cjtnbrFolM7wm9nbtUPVqG1blUhzEKe
LImojoD/QHaDjUtLjIek3hjlXi63UvuZptpXjiG/4TduJNr13NKEj/aFRkczzaFk/ek1YEmY8H0b
UsKThWrTFvqi3FaNzGkbe5Q26lI/GEh4xgDq+dXWAuINsA0Wa8y6xusV6AOxUPQefA8dNN+HSXDf
hAmMU3+2HTIH4pX5Ml/qvMOUjVg+jABpSPl8dMNj/g1e/5blYeJQa3qFQ7X/L9DqYNTIif6j8jnk
oIgMn4BVD8aAOuWum1S5X1tQRVvr1SBO7QeVSS6Ci/nbHk7b0S3HA+OimPf9vNkNHXluFozEZ39Q
v5k4ZOd25od7FZBq1NpBAERRRXdhxquzUSBglGSc0g0W2JxEzcsBvTtHRYyxof1bvDML58huGKY4
MF3IT+pQ456HeN2BDPG2hFfwQu36+msBqHzAltSvEPBxvMeGcjVa9SzJxT1KnR/lnSx2akkEk219
OC/7UCSIigLRc0rrLMJ7pLgxQ8BKDC0q9liGUof77ZygLab2seCWWeqwzJLvlPJIT8RFkysWKR8s
8jD3SjjEK9yIib94dCHKi1OZFTj8P/Z13XCzbyDPHqNffibg4uwS0Mxr8GU7Dj2l6KJkB+utpZ4M
lSZpwTWJBv+JEwHZ52LcrIRw8WdfXvsUImZzhcINJtSyqeJr1yp90pL9C4pOk/Z89h0SsdQg+nPz
V2DUycjFBb2BO2xkXtdhR8NlFAKkFfM7A96lDJ0Zj7CJruclL1RedybwIYyWzTWWXqzXUX6n7k5o
LvljSEMuRs28szea8E3AGYsYtwYTsF+owafZg+zj9C08xh3zVSc3erT657SJADX/GAIq9GbUpwwV
k/Bz7m3q8trLFMpX5Iy+Uh2rTROiQ5HLNzKrHKgIc9dUuge8NUTrjS+20leptjaHsAnQgtpUdXn7
uTB5N8zWxRz3zBYOP5YgGUxa81nlxybvTJETmYw4nk4gas/mBr9L9SmpBZsOuhOJUmkPNtMUB926
Mdu3HSshliJiYe+Pvg176adC54h8lM20A9Dvn+5zFwmoPMR+OprbccYG8QBcY2vARty/iVH0XWs0
HH4daeXNt8P55ir/3sTTAIu9x5PiwJ9y93cDb+xMO1rHuhQMQ5smJvXRMQhaYNRkscPnbGMJu03N
Qx7nqCQhAEvNIvz5Qv18et6WrsjkQ3uOYkKyCzr0R56Kx7DYPP0zPqHxmncHokDbhgHQ/E+hJEZT
gzJJtqKSIWvJOFf2klQlbfLAcbFSPwAVtRC+unf16wnvqXw11MfByzXgu9WxyNCYSCexhoxKieAx
Kz4ykky+Kx3Ptzgh9pQKT01jolL6gQZzxH9deULca2dNgHP5pokxcU099cfgb9z4Wji2ojCSzGsz
xyLJ8xJkkzEn5bFZOOgzjwvJKdh/4nQ9KmQpA3rNBkt+jnVCp6QExds6//PeiTM1Wfve0dpMcNWU
R/7mRG/avPYWJ/Bhg+dnWhA0W6k2bfysd1iY7MI8SRoS+vtfcmrocL3vEebxmrUcW/RjM+I+QCxx
0P6CCNXxTD3YiLsTfHRIZ79XoWmv9Fp3tJpPIvzPJmhJsMl5tD62JyQ26f4HtupYMgfQAkm7TLSK
3/PMnH7tzZq87u5npO9TVpmDZpN+RMyWQbT8SUkspiP8KuWNTYtAMsx9uvJsIqUmZ2F+rb7Or3Cp
6mORrCCFYtRHYqet11UGrcRCTIN7glJIgkUjxR5LVMfLdFwYEtUAmMFDkFwaAlD+zvV+Lz3JseuI
+VR85ixFf+CIK4LFEUmEidQjucvmyLy6dLptT2eu/9G626z+BIepCB+PdLmEf2ma8Te5eOSfU+cb
BLyj06TWlgWrMH6OGSUmp6EfP21moQx3jfzkSIKI/mSBb4JFVtzfOQf7Ake98hOgFWD06lRBAYdV
07XU33/97pluOFykdAibF4r3Wb2nTexMTAuqGdwlczzd9ifbIZNeP1l0tXMf74a3z5g7zXE6URqP
RISoPRqk/jgnyVt6kPmsj7IqjUulYuVO5YUUFd/Lur2SqO3/9lp8Wohdgf4QAEz2UqhD7tGyfaCV
20/zcxvtfKe1v7HyI5fjln4WgDadysXd9l7rIm89aZx0FhWH0anmbai9XagGORsHEAvGZi6gPwwV
l+Yxsuntr70m8sg/EZenxzjpx8k+9zl3uYaBSPoj661wJAeuM24cZjwONoehBMtSSMG99wFx1GbY
GgQ+yIVPYXSN7fij+0MCuMRoR7hVtNumhh6z8n7lop89qGRWPxLJJsF80vE8pw5zWxSlqaWKK+t9
Nsr1oMXWHjoXJrB0AiD4195K/JzRbV/3D3c5gSo3RHUNCgdGGnDKQ7oGxbk17J+k6XR/wIY1fmEp
/yR1EM7lY9z95N1UQ2ne7ulGQc2wvztXyQdRSAmVCl04mKzxHEwYpO74oO2uOsBHysNxK634fZv3
bkuflxvGKGB+/f7fQQ5s9WT0NPgpLZhiGc3a2hT59zrXa1cPx0Z1NrHixeXui+ldZmcYRnl9CXyQ
/rtMNjHKK1P3k53KpCbYhB+qStX88Iph7//4fs7izvbwZsVl7UIjvVzsSoq1Rc8j3/jqStXUhd2F
gP43T5vRe4frzXxpfTmWidvcuii/EDLOU5Xkxvjv+eRMOxrVAvLsyYIyHhnpD/l1FP1Wcswr9kbk
bxgEcHzXaLvHlOxZEIAaqzfQSggLodxdo7fAtTp/yxxlOChqm0vMpCkz1OdTDeLsrYmMx7s00iM0
CYBrB84ekB9n6BN9ZKYAYQ1Il3rIDAQ76U84kxYyCEvAqqHhBisdGuNV07T5LcH8HUfn/CNH5RkA
3n5jxxnv+ko6IKrga/yxmDbGSsAdZ0PdAedv1kG9Mx2dSTML9NsR+/XbYVz0CNwbyPt/kF/CUCkg
MBaLGwQ1yqjFqtuUcQjkUk4qjAD4UyluaBll3jHriU/4j+OFTLgQXRW65uBdGhYwwEOVh7+6EvC5
G2ZYTEdiL7Fr8SsSPFxPQJY1HFbU4jH5WwJ4OwmwsX022BeBLX4ZhI7HAhlb/n2zs2qFxAjt0gLE
swJSIiSUoM6s02JYVs3vguSgK5mFI1tyo6HsRuR+NmDkwvkbhz70LsFNFn7+6LF/3I6oFrMirfQo
XLyPs66uFu6c/T1/E8syAmpcFDmfuotZ9mfQb2GfMV+OlFE6lCCs9YC7dWiH4Emm3j4kEByNUkHt
ICv+pbJZChMjHjP242a9Al4IZfWgRxVNnZZMc3rXysxKSb1ALZDO938+bjascUkKoHBdP3/Jc1cE
uu+1sJEhOFnOc52W2HikyOj8tffXVOrloFWVH+sw+XoQ/4kvzimh3N8DI/zn04M9JiTFqG+qtwm2
5f/YOi/8HD/Ksy6+VIaZNlngY181KFeT/Vohn7uFMUsM7JHokCwrMO6XgT+JefAMJPrAF5fZDAry
Fo39lsRTHEzkp0v1XDTgYDZYgTFsH12HrsNN9mFiYQzNrGVV91IDRKyFeDgUi8DZUjAkoR8RAuo5
EByYuMLfM0Phdrbc/75Lx/DskdgP6B4GlE6TvUzBRhXAw4MIs0Gcv2RLFWIliszt9WKm9huMhUPh
mWqtNltR0U4+5nzHJDGxT9ifNR/KTTGgXQtpZSPir8pVCva3x7GmGXKE2hkbTC1JSQ+N21a1mbUA
7NRxvqBcdnzJxE+ih4WCW2Qi+T9urEKpkeyBtx48QgZtrS9Qn7RhS8Y1QjDHEXWE5d5y0cHPdXg5
zmiNYFWa10A7MMGxh4EP7lpWXlFC1P2Ts7ivVQ1buktEiJnVkNbZYPCQOHxTtInzBDo50566ZvHl
/QOc9lgiMRtAUB2t0ob5caXNKTht2tEx5jbAFusCcRmBvL7s3AaxkiF4IVH0vfsdMWsNlMNj2nLn
7bj1IElaq7y88WUHf2HIbz+nM4oNQswmgg9WVbFaDm+V+YbC3wR1wHGS3a2DxD6qHapU57X1eMVW
ctx7o63tkrjHmFukCynhuhhxOtTU3lM710FzKu5v66VxSrdCR8mjX1FJaSVJTnUC3pI+hLauLuRE
5m5S8vlpeyVhAIT//3ohuXgiYzyLOAGK8hNVarLtksaCoHvpFT+SinlZD3PQr30qI0Qn9IIeXPg7
BFfwKk0Skesptj4qOnIuDUGjOSfv5UEEY3mF0CXoDEBB/Wfpp2WBUW7bl5DsloWXEuARJMaECA9h
hXUnsXDYsK4g8lDNWknHgCuD44uIDznpU5GURwT9U5sGC1usm2a612xC3Mz7KcCEu5qcw5h+eVhh
SNCuenBLjTjuA/dv19Tu5y+Ae3HgsiOPid7Bfd3Ioxe3VJYnY7ee+RWVkj4miFzUco5AKXahn1WY
mCTxjEjcsVgUs8vRuQmh4KJs4QAWNNHy3shAE5mOrHQ/UhJtqgJFDBCPXSOjfNXrSp3U5XVd8+gs
1Ou49M58NG/9q/eIDj4FdyE5bGGtLE6aLuW/cjNjsNMLASSp9GjyKzha9UL9Sa/hGr9l8g7Im/p1
EZPDp39oPz1/8wrNHC/wSeAQ1O3H/+fyqVC9KVuI5sZcuHRp1wb1VhAJ7+L8fpvIOFDzvcCn3gIj
duCKTK21aEQR6mdluUsC2hpXlQcMzWqH6nGj7IFxQz7++oEU0hpHrA1QwqR+HXAjnBGpuh+kmlUG
O07TtVqHBFI5+fbCFKnACZcYmypRQfS1OycTYQvEiJZ40GtoRk/um2A284ZRSwG4hpOS4tPgkF6w
pHblR1SeW4+Uvi+ScjYhKMnj8gWgN2jLSAlesE9UQsmEMVLFLqftCsXzenJBqs4u/vwdvmLugfMP
BEINuHYIOaE09eo3GWCV39PtTJWlNjBVNBO58bzf63dGQiNot3TZGDTj5/9qhXfc9x4/jn0jScKu
WV7ptzV1BSW2k3KBSFk+5H2ntgEcva72lVvA1pridjXdtOrpBFEVl6SnNsxHcea0xRAj/5qrIjnI
mF5GgdYjIxmCaUrJOMGY0aALIK60oBiDyLCMqdUMT8ZiqRRhjSKDpgnT5TfEUEYU3RPs8Cd33mCf
+NCAg/2ur6QaetaMSwEvJvolExPRrfko6/qPtnTUwEPgKgTXF0ndL+23BoFWksvYTFqrZ5gQHDZt
rd4BC8wCWlwGIocKDOXG2Hhn20pNwzFTF92RfZOcK3r0it3qlWWX8ZVl/5m6E3b3SPcpeTaCbCzf
Pc9/avHQLts77NUiS0XtXkF4pPGYk0xy1p6RI2HrZKLghOTd0niTlf0qMTc3cNNZtZGXLRuldkUE
5VQj2vCEWCCUleEh0udav+0dG3egmt/oZUlgXmsNYUCosm1mslOU1V4OFTWoDplntIa4eQercsSy
orJxNQwaQlYOhBHzT4vg+6vTaYRoIAxO7OVFmr/PKhkr0hcbvPyN5/e7Wtxj2vrv+b9RBKO6TLxR
NUOONMc6E8vX7FsnAgH8ym16xC4co0zRgyYqbUJJykojhxnTi4xgsOp2K9yq4lMZ4tmssBVkRehn
JFz7y7RxPYOZbDTwZ4aq7oQnwVxmjD9YVhgPZMMYxVr2fD4WCIIdIDhcAckn7PQjnmraph3Q41Wm
NFQKdbPrddN5tUmw9V7dJeQGE7XOLpcJfL7m8Beu2TLg9cTzMgh9nKNOAmzHxuZKMYfTJs703gLR
w2KONAygsFZrab0hA3q5bpDWpC76TI0DyR3tFois1Kz4DFsugXPJAw4MWBt5jxQ4gpve7mHlGZX3
BjBxG4cjWdmR7xc/eZOjfqbagezNGax/SBVCfmu7AsVaruJrll6+yD/rcfH8KFhvzvqMQPAGT8mn
pkFW+yqG6X9tRCRL8QDyb+wpmSya4Zn8xsN2DRh0ZiC5VGxxyKhE38p8b8MDknYJweuu9428Jp+y
Pfe+N+He4NZFb5jGSfti2UXr/hxUMYRzuXzBs6JeDrQD98TOAuprmxBqevlgEPwaTPbO2yaQLn5T
JlT4l+f1h3MXZ3nrv0A1EhjlomrowtjZzOAnlmtJ+nskYXm2WA1HoYYkwGawT/jMpn1QXH3NggQk
dOfrff4vONOwWu0mVQ2pZHJkQ2t84imEsQcIO++hM+zaHWhgj4N+RvtwSGLLjgYuUuOP4rGeQ5o2
hxgpzfve2CIFEAsfSqO11kJ9xwoycfPk0ObgeFvQeJvv1LaTgfCSTr6sUoDiMapTascQF0Lq+q4H
C7U2KqtXed7yqQtg41ntHQqQaSEW7F8TeVhUebxvGUipQHMjd8LE4lATmcbDxceq3vOsu0WN+kWZ
nrO7fbE266soeR8A7SEc0lL9Iv596FlyQvgeVf1Gia5Ix3YmLS0mN+aagbSQ+8st9cJxjINvNZY/
KRkut2MI9Z49bDs8GCTttWDu4Ud8WmQoa/DKBAkjrAia2XWQMAuICV1q5yw/r5X1C6LleljnoPH2
acw1eOPmCPN2nYQH59mlelUmlgwCQPC/OwAteIQVdN/vkOypO+yoDO26lN7WGafemSVriHJF/NE1
z3N1odJjDN0FRp+8OBUxzfzVDkO++T4PC2L9eCxTZ8HlmDc7vaaxCFnYUO5eTBiqZIo5MFSNOMza
DcHs+TftJOE+gtUj1nkkLlT6zTh2tjcIdBJHfj8Z1OPZNhnTUmx4oCh0QSEG4L3N5eiD32HVYV5U
U1p4NtXj8jBCa51MvcVA8H0dryy+k3zz4tRzW1xfN4JuHJYtzJZaexvTgSVkljDTO0wCh9InUumC
FgMajK87wuwq2yq2DmTSaId9AgJPBGYbtzz2jJGIzRbFT2AX3AsNUiwhcpUujDmFcHlpn9BcdA0j
DkbeZ8J4R9n2x5Beics1gTF2C0B/En4ENVvA9j0y8xcXuat2rSadVe03U7H4CdZdwHmqQUjcGeQT
crUa3+nFGi+12Q6S3kkdzaQY15n5ZkyDotyyiFITdqtsQTW5hGX1FFWP5zFM0Aq3ELCngga/fay3
kqg8KvP2hjvRnvTtnUaBDlVf16g4dCp2JCUxSmQbIP//Rt5JXvXsGoUBHvrUp4XKmq+i4K+QJchO
IsKGvhFMe1k0Hapfl/3jg4fq2P3j7ZuvqJI3iBQL1t/Yy6i0hlR7awjD3+7ZkyyEN2Gs7z4ZT3nD
tQ4BKoMGztjyXTAnqtX6z+nl2WWqo9hN+qYH1xgtmuVXih1x7ULhBzqJA4eCDqMFFO9N0VFDx7pz
wN/OKCde73K3R7EzFgjB75QXdzaNKeDSprX8n0p3HKsGm2nAblXwqEk+mQunWCkDJum7nCY5a6HQ
NwZXgn8oRb5Ziu69T/zb2xAjpGE1NkfqJNS712NcCLa6m4DkTdvZ2O8KA8a6bLw9lIv8NBgcqLUA
poQ63ic2x3nbsJFWdmsYwcbl19o5lbK+ii9nlK2Of1uvGwk/UkKoSj2e4V9ITpDlvL7p/9e/mnJH
VmApkcguMEPDeiYPr403pS/SY1NPH5ds5dDHREAnfJBwilI8XMYrB+8O63okhuGFf2NpqHjWh4M7
VbC+ftkdryibpBkeO2NrruqS5UicnlsFTlZdDb8y4rQ/n7tgULfX3Ill/d2xiYBHTcTvsEr5k7rM
tJREoDqQsTvOCixp1weQzJXo1T2sOFWAX8ESgmAWsFpYIvQ2nMSCE7kX16nr5HdGQzbEAmPvNg/f
2ExqySwTkdejUgF0ncyUVD9HnswRmU9dbo4G8QD1snwwK7Foch7Dm088enm36TEWrSwJ/HNycEOW
4ksG5tp7EkwQBhKbOqCaWGriCyxLEUkMS7MVgffaABmuJ1xKDIPpOhgm3KZuahWDhW4/5howsIpr
NwynGlx5hSVkbKNjZMZLgZkTxnNk6M3VvDu0e9Iw3IqDP97+sU8Xvo0POWzce7stwXYrvPSVBeyW
70uwmRqr036Z7SFsGbR7Tqloe+w39kHgS4QqSpcg4c4QvJGM08/ajD66y/bsua/W9swuDwVUlTs/
JxEbNiC6y9lBt49+eXj8BZv1gY5xKN5+mrQcqycmp+rstYCUEphW2ZtTrBS6aaT2JUEVfQncBEQ+
xGhpdZcwPlaG6Pqdat8iV3G6M+bXg3buDqmhchLukeSw9aUD6BLnY8C9qY8AgbgZ3vbjQZSV4aqd
hw5dvQgdUjba5EbVcQTzvUv6xvm+ChJj/8Z9+03C9++K7Bv5y10c0yFgciDSmFG8yhnE6DiiuVD9
juv6uCt5754RiAJTYO6Djv42TcEkPrbiIbEGd9sbh0rYTCIb1voFrYv6UKKSk4K6v1SuENSNejl0
NI3rQzxM8sGY1oIhSSe/VrTliZSd1ehwlJOYRcmQpLoh+FrnFWd5VP/8wDTZ6B6LkfndWjrsThew
HSECuj+UqjMxKnGSbe8Xfl4klTfSSyZqU52brrRwwgoyCa546sQY+DcKJhQUAEWfthfs68JfEzaX
PDgwAP9Yuc0RrzZVIoASQi1ihA8Hqs3cqAnYJeKBBI7LZ4mzm7/DSNuKo7c3Ir+scOGr9DsSoJxO
vXmWCOaO2/GqQ7/2LLyUIIq+vvySv3SeumP329FQDfTeyrSeX91A422ydnWsIiCou3uI0eJcOWKY
ih+Itwn82uyyHU0VwFSQ9Ydbb3pMZMdYmBakkVIHVPVdPhRIvK6ZYqGV5VXxFZ6+N2UkcBDYoiz0
G7mwwsfbjG56KatSCzpoUT2G+s0EzTnKxQvtPdSgiEghzEDkMVUOOXwWlLDScQ7e0zUYBJxqliRl
FWzzY9Kd3RckP9+oZbwz6YL2nK6WMJtBnLDsFGP2PJ/RKCxMzMz9Od27dh39JWFS3JLUlOii8LWi
ppcyQbnmEMLlQQRpS0SfLwa/wdFIHoUiquKtVfnotKNdvGOMbNRIusEPpF0A+c2dqcePKtq7KoJH
F+ADwgxezG9gV03X3kXNUTlP4h/geYDQnkg2eEmHnjojs3WIMIy8TbwF+lp8qw58XAcfrCaTTXid
J6BzQJYhmzabgKJ33EjK0M4FaIeopoOQo9JvGzj0wkEWfM8eGw5RS+rqvZXNkMKux/XV2jxBbKte
c7Ia+gTq3umj16fPYGxHl9jOV4/02LypVYQQIc5wMgKNI+gU0qIvpJWTWreGYNysdoeH7tZBg51H
MAdgCF9ZBuBcn9V5qzJMvUJq9eHx6/QDn92viG7z+ZSiA9+t1TTG9LMHqc7p9sRyTWt1s3H1GWqh
GrfY1AylwjK1lf8142Xeyo1oS0MU0S7ecrJphs2SqDRIapBJ6QxoKHElbjy535Iz1F8NremAiFno
CnXVeJ2F37N/DsfjVVRTTT+a9NdMz6AoilHfU+kqaQbWP4SmqlkUa2awjVIhgYA6+6b/5wHMeFzp
jtW/uiAfl11P7ca9UlVc2ibIPxXHtktjcsuZMwqeFJkheJ89JInQzLUZKc15beilTIuO1C7330Ks
r3wEdill3usm6L6AE3gEw4DIRjYAblH0FXMRIJcJtv4jXI/ko/KH/0zKZ58z2MkTPgA+M5Dr+6Nn
upp6GMWsLy8RNiO5JfU/q9QGHTNVhbojQrTNyr3lRN0i5QgBsWlRJg1z+/W5MNNR9oYDwot6+qdT
QQnqLW30vB2djq79lkigSXuLttRnE7YLDh+c3V6WSnqDo3RLZKCMMROqKKNrfVpMjBdNxMr5vc7g
zyNLN8V1NGlsPmZYoj1FKYUo3yBRudTgkAuvsWV/E252JDqw/SV7EYyiIHoX/xjPFKRuuHUz8y1g
1uiQRr37fSrvoYJpN2EcSllyMZsjZ+e4JgghrSSgMIzq0FlZDXNYRSRxD//+tiBmf7Kpovj497F8
3yNm6RDWojpj0Z6rlZwq/rWhpWh4O3gMVO6VqYzSD5YiSg7BhcMPwY2qR0867ub+lBRn3bu6k7KP
oUxlXnlMprmbnaQU3+Z1Rr913WcKMbwxq/J2RaOTLPXtJ9vlRLW+N/TaA+IJPH07e4il0Wq5FTqb
dUDrp8SMSdIyVgP7R7YRFbcuKjTcqP15vWDs7e3KmsvzkAdZC295WeHAWn0d43nkWlvrAmI+o5Gs
3l0wp7ZjVHD3GPxwjLlh8lTFCDbpIC3qE9i40QIV0cJKYrpXUkZCr3mtGSMLGVQufny0lTyVqiyt
ffScNqTFyr7eG48yLLfXlU+hXPQyrSu+Pqa5c7DHHPu4bsUPKwBKxwAe2bxeOkuHw5cPzRCD7fv8
30JTEQ5wboHSo9hjCG2tO1T2OOnQaUfkayqe5egXHqRHlJt9QKsNw0PPqZnFA8bYQxdSquUM1f3W
BYkWdOMfWoAXRTfdoZsjYiRlHZvUDrMl0PgyN8lUjWSyOmWJXzv3PI8pFIHRgCrwVciGTOm902qb
ZR+/koINCYwlKHTkSavRxMpk+dVCq1tEXxmxAgVKT43NQBbAV5Y2JxIEluFVJgLCKZY+bWnCrFnX
4m4I2+NJrJ6662StcUh0y1lEWP2ZvmlFCCtFjM3HinkBhf4rN+wy9blWxjn76ScuSl/auis+0s7l
hrkMovq2rZ23ymqd2X09iI0GOnEErtKEmS/FUCAg3LzWKGSKZ7AlIc1Ne5E4Z7yZDr2Ir5AxkmcA
gAXx2ZVweawiq3HRUTaPKPsvOov9TeOY1FoBxPLscItZYbDtEZGdaVC4ZHPtcRZInoYazLWFdYqZ
/sM7NFNzZrY/2OmvDR+mdp/YLz82Ph3SspdheYDIkdxtF2H7EpLZcFusPq0XJBtDhSj1KAoXUYFZ
QtT2tc6gWB/C4kZadEgfx7k058ITQ4ew24p1jWA8XW2oOAr6RRtAkUmDhapeysEfGg4v8BBUIVh3
EmOojs/Ack3Z/9XRrAObqu8bjEdgQBrh35sWzmPQVnvY+ZLa8QP1qoIEzBM3IjUOVs3j5fRxQGgd
qGQoNWDMKLC8VHeOpufQqPtxHJnA4Ku/FVxpWCtYNAWdrEia251eBaRzFvNOo8qb80UckBNZxqe+
F2cJjrHrZVvRXLVkIY+64lDWRSridaHWA0F+mN6a0OdsXhEnqN6SWegzHwjHNZDeIS8SKwhRw7LM
jHYp4P3Q/WK09LQJ3JVx54JKvrqHrZLoUV8GHbPMUVQzEeanW92rZddFrOAHNOUsI3C1XmA5X/Mi
OslAkyFZ9bJD/esY1ux53D4mIF7MxdnDJefPJtWIGZgOG2BUy11Zia26F5RWLH1d5/V5ub938bBs
EKXE54Xrt0QmdYzDyLpa10pFPnS7sxxb5cpcFRK/nqpr3dop0RobYR2inPVIFugLiLMuRnQ+IKie
73HnGI6cFlNNr6Vl50EQ0wVhL5rvucElbPAHtvBDT4OmKV93dOSvurvvBG4BayK2i0ObQ0tUs3W9
e2uOL3Cdyk7+CwLBsJZrjtRpbnePOU9K0RXdGukmH2wGKh7oLRZNeDy01TvaJe8JIHGFBmtYDcgt
+n5iZJgZqUgiVD0zjZGKctW4kcbtCwuQR5JCVUeJVQuB8/IYW4CCM9JwoRwARIo+23OY171KTyhI
oVa462098HoeO8hPGOt+DPsHCJdnFcgb1cfZpkXbAAr/DqQfSAjZqjLFExkwHu9SVElSToVtecj2
QRNdEpmKx1u4niLaYyL+6ChZE4l8VPufTMPpRAqbHHvv8C3vpwrtg9k9+lb7iJkgAcLev+81Vpic
trjz40fZ7HCIGONTFMtWmab5qqWTC7RABegJBgRV5m0FElYOCfc5DLiUisADQ39Jo8utoLVB4rds
o6HDi5NYTvXiX0c/YDROAx54UOquCj7ysyRO92WBtwXT0JElqoDA7dxwFxwQnQ42eawl/pnXAMXt
Ng6ZfLOSzPQBUW0GhLqxuwiyonva3kZDbJvnGbXcnyln+zC+vLARDMk+THLEFX7tNRDqpz8XikFu
cMgIkWP9zsmkwWjRsQG3j70WGiQGwT4YtbMsmDPYUl9gFwwihCt/52PZh+IRK/4sphSWHVtgvWkK
GenkQBf3WdFC/u8pjJxCB8IWjeRH2U7RvB3x51z3PqybB2xMNMDDQn7RLevZ6apZCWD0NDmC9Sl3
HMuaKvlaXycLKjjQmDaP24aliIgKxFcSTg5MpZzSp3MppQQhy/YdmH9f20MoD8HivbFtsiwLBoKS
P3w/+6vsT8YCKRoEwABjS49aB8jh87P74Wz1H2YBUxoVKBMgwb6i9wwcg5s167qsjmi+soYxByu6
mkGVsE5hnbDAIpWbhwCLIIj4YTRirAApJZ/KIDYaa0Sp0mnXhaTrDnHDol5MkxhjZvFw77gtl/VE
qJQWW7Hg2kYH5ofe9uxnKRbG3VAMp8ULiuQ75twKPPpyW8gQn3dp8sIfUUqpEbMZKo7IJ/7a8VCN
NgnvJ4De6h5e0NazpBTLc72roYpA8m7PzWykW0q8SSLePnDUtxoiPhKlLE4yRGSDEqI0p6x5GdWF
9GawV61qd0m+6zTv1daAlRzUv8tFtvhevqEDEK+h2YV8bQY9Ac20MvElPy9w6+hMTz0Zcssvk6BR
BtgE05trt9aH5dF6mLe6YMoKkArb0kIjQusaUAW4nkbGQhiRAnZDvM5RYGXRkiZSDPgIJlz32I5J
vZCa7TmQTVDNSfNueLI+ejL6YQ9cOGT0EL9tPmHks9opfE32VdPQDU8BKlkP2Qvp8UwciCJBEbsA
CXcbzicrVZcJnUZr2U6sIj4QZtR1ll9X1oQqly/d7xMe0NJhqPFbRgEizebuBxwOVj9bWTIamWIk
LyrNC8pRSq27VCE9x47AiVcBwqiH1VxrYSsRSL+LkA407GGpYKrWPypsQRCuHd5xMoCZHGU48FlB
DkS0yeNxedpW9Y2vx9uvZK+6nMQb/HPPL0TAq/jYQW7dXRdSX6YJevK0lfA4h+Z4f411Megkm3g1
6u96w0bX2BlP38L1rww3BiowVmQJ6OUn4f6NUPwZsQCKmDt4FRYjJTSKJleLYf3XRhZGY4V1GRwo
cKtawK9y55RNvJOqlvqqtVqjfzR0io0f4OuQ8i4fnAgl7aA4yg7CRt+Mdmm918EVREvs6Yb8uLpR
NoUtmbuh3cMz2OKdn1A1xgww+ogw/kR8k8kB5HoonQa6ZfMv+iOEBcjG03DfRO7TqFvQDyAiYfAI
/aQtx9ER9F63gfncZE7w84pXklXlC52A9C2jfzE4Bppb7XPEQ8qCWExXr8bp7m7JkW+XFWGbaeUa
oXn8Vxf9SDORocourSdlqBEILEDacTz+UW3vbIjchFJ23nRDbHjTsKbZ5UX3T1LYX5pA9wC6wu/8
caf+XHSL/k+iycLYAkcTZ2g8L7JIjX4wZRNmwiAaarGJShDxuvJtd3mhVYwXoEYPxY9H0UNxCAJa
eSZNhWdfjQaI0fBPUytaKPsiKeErLhuOEEiEAVaSxCbXc1c0uJk395EBdk9XKnUeQflHIZWFdq/Y
U/Esq6Ap1hzg6rNcjrA6PtBAv8A6nHuk0XmqBwew/2spXjWBAEptUv2UGnaO5Y6PmpnMoIZSUDh/
DpoM7GNGuy+vr95iBvE5xhAiIkDgncODI+j2qklxEqRW5+qEkPC86qpwG15DHoIoMIgN17ZXnA44
7VOCGl8O4WEz5VKxoSgFFinftsem+72Ap0tznEMZqcrt+PV2kSc6M5VIWg9WYwvS8xe8QNjfIlKp
DxSnbHhwVIlBB0dPRHJZlPjG8CMy9uDGpphSiLLuOlXgfLKIbzdY0VnRca6jtAgH3CZCO6Dru8f4
6HKWI6cd7f1jaRDuz760WqDpcF9hbNaCAfFS41y0aw/qIhKbVxup/1aTkDoHXthVRKIQEw2OnIt7
Nt/urY6oaiXAnZgB/FO0KM9HKsY3bwhTaWDusijIzb70pEXQEhpz1AoaZ/PngusEDC4ChUlz3sRj
qXTQ1j/UE0tLSvhNba8TqUv3gMoFcsOe28+H4h0MAbpx2Ec5ohZMzgYASWuKXgbfQ3jqJCornfle
ATsc1zXMb7WRhfs8SKnunumy8orJSKp3TZZq5/n8OFbo7Lt/0g0z+h6XqHuaw4VNGoeKI59aLR0L
U1Z+TDiZBCYAtqPrmSVGjnDmwT3mBX+4LU9z1XCfawp8wgIHmrfKWDcIy/Wds4dZubLRN+RcrNX9
TCoBp/2Nu909ch5oLu5qcSDMr0Dr/M3jdLaO+BIxDDtN22gVI7v233gDbG2iVVB27bLzYdyxDE/A
9mJDoiwHyn/mrWNg730Q5+CkrxFV5IAcX84ByBk/3MlaI4/MV8c5c3kVz/sqrRqJDJPyylJaJcy9
/8tocEbspuB8g96Z/J6a/X9aSVkZOrvHq2bq/X8WcHCmwIARZhDZI3Ifa9dNSmaofPDGZbEfMMm1
xeQFZlRsGCsIQgq4owuKe3TFVDH8aG/jV/gzky+X6UZqE/oe8XfBIXLlncc6SGZ1V2twwwp4RVAS
GHW4AyiZZTYaOiSw28xrCIyG0NmlYNqW8C8NZUGzBW3a1nXxgaXdGFW8Zfx1pXRfaiFthKB108c9
yuNpylutOC+01RZD+ZpX+MJK8CeCzw7H5H6l67rvQbl3roxUrRe9U2rZSBckVCxQqzQsCv+0I+nv
IPAX7YHOwUlVGb9jeZKFfeSYb3rG4eI3xT0trHHQNTyO/XoI/CWkigIgLGOAgxDfJEpJfH5nYWqd
txEXvQ5OKQNrpYTqDK7pDdpWnLhaBd7udBjSEWHeabfG33HJLnbdWgH4dH08wt8/AAYOPJuiW+JX
GDTLLMPWqAstQtDMD3xNg4ZAEC2sPa027AmIX5ERKkv0TP447od0v+QmWiQacNCVMpSRRtZKt1on
/SyOrmgIBMQ/OPTfY0/xsxhs0AzZ8gN4K1PkLNzhh5Z3BABtTZNY9UY3sjBQlBLOrn+/S2GW7XxI
wo9Rq013VNJgP3E22wX3bH2OBdouGfgNDYooLIOylqlO6fDvPtXbtXf3hmtdHLlBegHCjPrzoxCi
yBRWKiRQ4eA5btzx0cQ9oFKwCJeh7j5kv1Mfok4KcDAZMsK5uCf2lQKej/7dOjDsYNnbMTMSD0px
1VA6p+AqJrTBIaJ3+s2CveODz0t7Qxu/CtIh/T02J2xNCYSQ2mlyhq/vd581XwY5VB4Gs3LOlTC3
bdbPSQmK6Z7u/214GNVKRfeRwC7JtuFcIkXT6l7dTJhuImzSq7ADexF15gDKLMpvgqJh71nf8FGH
RS5Dne/NuLSXgCXY/gh9LTXSnovJ+TOXk7MpWrDTU2Wm/cGzdb/NAVGF/J+qqljXnnnmU6Sn0NO/
zvz9cHrrJ/xUbq5Lwf25mGrsyu3zHxJiGN6CU8xoT/uJvJgwmNI/iaOLpSO1+wySZD46gkEe7ry+
8zy8VJhm8m7eqXs/8BxFZGGLoyj80xTZeTIz7RS7XZl/s+8Apu0iYnoxmZXwDqa6mRZ5efdnVxVq
r9mdXUvCnuMSyiK0n75N9qpXZajRjdB5T3ltIkSNQJwKv+QhlTRdlau5uivvwE1gklenKuzqWolV
pfWi8jRT7wKQdEFPKrUn8r5DJNaLINaezmP32DYLGzeQ0iQxi/4HeM3DGwH1DF+PjwuOd55cTnju
8h/dQnmaZzfQ9ENjQS9nJ055lgNJqX0kbwqA5fiZTor8J097NrndBL86guKaHrd/L4CiiA0FaRbX
uLjPykv3zGEuU8fdSXcmL4VneuuZq+hab7eL6XYXgGUqi0v6Q8Y8QbXN4wPO5i0+wRciWDy61oEH
FYpRNBxwGXjMgUaTaSFNHfcpHiRGKd7kgvHPsevxh8fi4wGGmXinDXkbMVdljoxt6Mc+Gfw9WJvg
GwOwTqzSIWq4u2vEa4ACHFtp9My57BmcEh49grZYyI8zU7tTSilgn8Ps/AjXsWwHmdOgFMhyJ9Sb
O+bNM2I/BObLbcY4eMsq8FiDjavHyWdcjIf2Sm6UyBpzseU2llMQsFFcWDCMtX279BwrVQ0PjBGC
cUSnqG1yFP5s2t60zB97oMutqm8zAZkg9JOgbo6tFDlgbglOnyWIQXZGswm1t3zllHoVxAtOd02+
zhC2iuJ9Djk24wGS/0k5MQeFi1xdjs/+EbPnSgBfUBU7R2Pa0O8B5mAg27WOif/TwqBzyYpINv35
Vy3DYzrPV2PtZgRtAqayVQfufIlXiXvDtfB3/0HfIW0nDRIi5PjmrdO0r/7sq2pvB2YelnMg+VFT
CkpH2d0qWmkULCsMjiAbIPRLYJ6TQy/hvWu1u2wRso2vVfoEgzm62JVd+zzTlLI1H7ouBAUZ0DuC
SoHHBFXOxZrQAZsEwpnLCQ+b91YBPVVuMR++gr+FkraFn3Q6Hyk9uS+Za0dxKsrcnWy+S0jFH/sS
NQx0f4Mq8yDHFpX/FWeZX0sQAWu0/RwP+oi7mcLxDg8uofQhI3rK4JaZ+9pfxiwEOUUWD13BUK1P
oWGScH/HlsJS6y+ZS7RFQDBjkq3speDrYNsr/sMfNVxnaBCWFqI7jZt8Sr9wuZn0MOd1IU1lwWJH
eetBgQIAZjb4+QdvKv/onNHKCOE/bcvw7IOY49Y0ngh0m32LM8IZ9KeOIG3iIBgpuz7UC7c/oFxe
p8Q87p/tWzeMZSp9asILH61vysRfVfCRKU2pPSwXIoT0ix6LsXE3c/wWvqA966+Pgzzvq8gRSCVm
6fbbq8NjJldh7ztPsH3NslhVUkbJbWi+DA81ByNj1xcwaM62yQwABjNxGtxz2fAALNiUEEqyqYkq
dCzO2/3kxoorznGjiFVV5a1UwRC70tmAk07S9ME+Y0r1wTE8Oz6lDAp82W3YGLUri3oYDQMtT3/y
4N04anvccV72Kd5DLuGNPujI+vPXOdR0hbmmqE4l4dOp5hhmCfLWyXxn7ATFHn0IsOHjwxLxgyZ8
j+ZxGG8tv+9u4oTeKvhxchutwtKm6ceLcdGPCZuc/RmIRSvuCptIfyFYnp4KKeR8SczjjYwCKz5b
tqTzLX2ENJ94xYpQ4Ui1DDgWXAeorp5LW4t8cPu9a1q1ZlNkV1XYDRQImLjuYx/fip0GlsdjWFyN
ttMeZ9VBf000lDlLBooLqPSaWBREdALeT8nJjpVQcRuh0CcF40XuB6SMNbUVZw3wCg6oGAa01cxw
gIAsYgJ/qq1I1lcQzboxF4wxMFaWp41UzdnEZwz2utHprx5qJ5eqsm0C/pHhYVFyZBErGgIEO5DQ
44CZ9LFd+R0xHFTqGKNdvgDFnJ4DbydLgwAIc4+QHP8tD5681NtUM8uxM01eMQ7dZoakNNUhvYj1
ZJUU+a3ICEsSF6TOPBmKLlgpiSYQkhbrGlUuPm4K98L8MCaahP8laSTC/BMXpqWgygzl3XR8aAGe
8AVxHgC1W0NRKaXE/bA67NnQ//TU46iVngVC48Onv8bOZL1Nr/8f2vT1xCbEAphvfG1L1yCz6pa3
CJpUqDhSRIKlE/IocyVOTaDGrQpsZPe8OJeOiUPVY0HuwOH8xYuSwcy28Nd5YI0HoIiVgpFfNn44
+cYRRyP9akuWBdwfMi1KfScgecSRxWPVPP3SAuO+IuxVVO2er6VanDgiby4rov2n3fXV9Dny7VjG
+58n2DXx9fWtsMDzbwdIe7Xmesk4RiPVxZ5tRS2PcwWORU6VVySvIAJpkP7ih4kZbJGhFHQNctkW
/aKyAzd/J3pkhQ0mla/RUbF9WdHSuBugMuzhr/k8EgV3zpmqm38bxJR9mvJ6Nnxf0RVNOhyy0Y26
cfon/ut8NXq1pEbU3ncVhddCU9YBxo+S4uOjhVsblKOH7sK7MSsfhNrkHgkisqXzD0TbmiB+HkZ+
RJETtaS/Wt525sfi2A6emOkwuVT7wMNtssHttXaaL4XKy3BVZNBB2tbmrNk3zofGQzGFevqTreB0
zdmwzCiJ4vbiMu+/33UFKoIyVw5g9NhU8G82avNp4evnPIWSSxzmAniff52Ai1A5xztYuQOy4NWS
+37GRqWFPM5AIYqCFNAfYISSlKczKTiQSL5ectP2pCVPm791NYTfsWQbkkGLCS8fl1I7xcrATMUS
7JP9T7dBkruOEYiD+tbP4zUbgFR2k4P5CnY2tWczACDsKXVjIzEjHf7yJ6osEFqV9pDi5VTK9Z/t
obbJ/jAZk2caXuLNWA5KJDbU5RSBq99xopFEvQltGMsx/vAMdR/C74rrmCCwtPRcq6bpBm2em/o8
zelldPe4z3UrM9QTQPxc4IXX356N7xYdKIrIWabvQgqRzeJZGgnUMGpT4LRUOyIAne/VejHVKMwi
m40J8FNDOjcwzSO5VBFDXJj7Ezb1uQs+J1+p6SX+R377NsCMrhr1Ce8a+YXBErbvnN1Y/byxZHZ2
cPyQQsKow0mXtU2s86DspQUCc+5uXCclaZV1ONEDciSmIyLPhk1+w/B6e2E//fZm/1TSM4yytITP
2CFEuOH+hGciWCq5AxoWGfgsNXYksA0peU2+5BLGZ2jrEvSQveLDnGTehJilDjZWnxIV3bqM0V5f
eIbwvoUDLmXvf7b4X/elHeNmb9YZUqh8oKUtNaUuToWpk95m49p0uRxKlw659/x3T+zTmoC+jwLe
q7BdOky2MupAfgbrufEqpmRr6uBpVVI2NqrgcmgtX8nVe6dQxUTKt6WA/SgfLlL4sfdt37BCnPLh
9Gca2Rmc+V7ibQjrOcf4knEr0iRx7HkLomQMElPzpHkiGMW7DdIpe2sl70QttYn39SAtNL2xrNAD
YmN3d7G4nKLthT57O6ltdrhYeiT8iZxe29Ku8fVH4U8f8f1rlkQS2tHEGLd9y6k4NtbDflzs5JEs
qwDuFvJqISOz6e7tbjpl6RyY6aEngL5WNAB7VHuMNUv+ZOdbfR8LLkiRPxC1JtwaM4pmWPWuLMhl
OvTFWnmuI4u3cUsEM/RrwRmOgkPgvXa8oM7mx0ZhYDfE3kabbNd85P41rnvoIYuWAuiQUGHAVKoF
xcaFS+kJNepgShmM2dSeaPIv3X6TwJQa8XdIaWlOB1nErkb3tMhaSKj6eynSBP7VQgzyQXMQqmPK
Nm6OIRkIdn2tViW2kAodBSViD5w8MhgSO9TKz+avd0sgbWX5iSdpoytsVUAc9BRRGPDvpDrE38Ae
wNwqcDl1w45Xr68qxgN54lUZQbrIJPv5r67OulKpjKXr1x1qjPrpPmY4SwYZ2S5fEzGcDUm/ETkj
J4i2SPIIcArTvU2EKnhmtE4Cx40rdkjL4KPC+L5+V0PpCV6GXIw7QF0v6hx4yYsKk2en+gjSM6wk
hxPbJKMRKl1xFZltRO8+lIXdvzMBxMyffHI4NJlOjpbjf5bu1aQ4SWIFT03iJiVqpFWuVlc4/dHX
57WxuIaaGN98pplz6eA2Ja8RecKblzmN9XJ51BOCzwR4v1cr7ebIol8XiBIcQasptXRNmjPAOPc3
9ndnnqE6rjJo++GQkx22hYDmUKWbTn/iFZDr7zjEThRD32D+R3V4rHQ0bQvczANDZjTA2L0G3Xfk
GYFeIrLcVQF2gfrkKr5qrdkMubA01GQZRFiE63VKtlpPXobp0kqprL+VKKHHQM/e7pQx4/VT4pCx
HXfnfboOxycJZ5n1RhoJpYPdtBmpMC/oz6sZ9x8f6LBuV5nL9V+nk6m1+EVQlJQxtkTW0W0XBist
+VKYXD7Ct9fbtWb482cIoHNPr4qvi0jO1Tuhfm4wWqYmOYxrQIA9WSp20GzxjdrxnW14+X6tvA9W
z+0H/T0rXz6pL+4HG4TMSOAOtDH34goKTtExfHD/c3NQ+yCKwq8aSvqCr8biYvobUJpBZ3LPc+K+
vyqrC/1zL11YmvYOZISwkcquOwNny/ey7R8tbpBSBW96hIj6FQTAIHQw8SLMib/CR209Miin03gH
6tYTXS9QCickyt3bva+pIYbMX/LWKm+80R2QOCmTZ22l3TKTrSuGhWtfRlYQZYYCemZnNEuyy7q5
SLSoGH+uDjNoSiBx5lUspsQ1Iar9bRwHpBgTEOk4v/jxyRTQ15vDP4vWu6coqquaUTx/NUQ0/BMx
0tzYLViPH1czArosDfFLhoHyie+im3YIya23wvHkD679A6Om3Xj+buDe5TbZIg90kk1yKvV3BH5S
v5bzSOUDDSIVmGLbZNrmqCl4nHqsB2beYzaZzBxK+b1uX0LcZOPrAawNH6aOVX/noZi4nIkIHPnW
0SgFWiCk8jSGruayjJVW728EKJcRlm6ZuYLcidXRN9ClibWEdVweCB+qzxQn4205rNnpGsYB7HO/
moG5O+FztsQB/oS2Z5+S7EraB+kiL9V8cFMDWIiIyJdQGjf2tV0ZHx7im/oQfxMJgW+WTp0hhGZg
YmKbWaknWAzUB+/pSKx7jhHUYJ4Oggy59jzGH7WRIqxPIU9qIrOFekByQ9hmyc/d0pCHRpRmOmwV
gz3dUJjhzP8Yz1LtyJG9t6llDWttIPQNaPeB3FuHDdvsg12peE6V4aYL3DilcJeVvPyFhCt/UwUL
a7hKHHL1kHmgXbEt4lZmUy+p+LFTvLCSjkYQshaxq/PdTfscMAeETZvu66ofCF+kYqilt0IKhjyA
4mWnPj7BOUDsql2oUTrL6hOubL8nxaHYNE8AoCxt/XYs/0UXcGId/lj2zlWXudJZGmPqxddW9jkB
6xEvbeQtOmkDKgYc9NGHQNrYB6CgzfzC2wBECyYkyqeA6MMVInVsWcgSBkUeqQWa+dzGOFlzA0Vx
8IOKE180HJ2fF7Wg28MUpKBPwr2RzMiP5rYSUZ8SyFmuvV3e2paYi7mZiFcmIDlIAi6z3KVbKaOA
wkh8NYHr83pExZ1iwXhVKU3tGMtDiY3u0fsIUrDuJcMtAcvqsoKXFFHH5asxt9jlPpFojSMRYog+
K+YBZJA+X9xLZv9A6SMNGfU350Q5H2jbKBUVIIB1laWQ+2A2xfr5LL7qsyvghxdC1orZpKwOgPfy
yl5yB+5yEDmL+9gc8tu2/AGyrHG4tmDPSqmIbkcy2F90d+uKm71zEQ9wMgrkNQtbUvS4m30UdsgN
LkF8vsoshSaj6ft/QpQCuSgznpOsSwy275cFFe7Cq1pwNue2qIdNNuAvyHoWZJKZDs4hrHPnlxBk
uNMmyAY03LMGAVXfztARbWC8xjcYgCNPysTDEfjSHAXX2pr6OUHo2DSyq5hkiU75M6HpkYoSY0D3
JFT/YlyK8jjrRaadLJw3JX5wMHd9ktwJ/5H75NpnfBEA08Lcx3FsjOoV5fPNR5rbJbtmhZoKy3nY
dAlqG4YWdNjYjAZCbgpU4BFJQONzQ4P4pRX1TCCMbJPjH8L4c/VQcOH8GDX8beDw6GRNsavC1MTp
y1q7iK6iHdDvUJFMsAWps8n7HK04MDRGxfqMIeb+OrN2jvMTIoyCWWajuOINBhN6rcDnSw0A5Wjk
rKzDxekcRsBDDHlka2SQu116NfmD6h8UltITawSE93y13zkEe6OBFrIlUY80AvJD8VM/1I7b9vo0
EBTg4aFI3R81DWVZi14ixRSRe61FCgiqqr6GxhZ3OmTN5mFlOS2kkukytXrYvpzvZiKvlgjPWeo0
5TwbJFoK2VXck5KWOG8OLfIFuV9I6qcxr8yda09WlJsGw39pC7dUqlQRy7UUV2spD1TmMnknjy5M
UQGg4d8lFPCANLT0r+kWQVmrEQVZi27fpKEHs3WXa5LohTE6x1HIU7KjsdlI9lFxfXckvaBu6cCl
IIFK1noVCYC7RzKVWmsZwnF/tJcl7frWlewYPtfyIZDcpDs1xUTuIkkVKAqy662p8+uE89XAlYVe
X/ElPRGDCgB36SuELvzCl0Y/nJW4uaQx5JKmDHhPZrzkqGpgKQF3SjMtMhPUaEDr/DkvYlvzRM8J
H1R0BKVSqkTTH9BA6yeFrUUlsu4xKdFT+ZgdR0m5gDA03wrUVLBzGW04T/GmS3V3UI/asE8OYS3M
0CFde5nL2s36ewYX4BVgHhdTJph8OVZ4UOVfeVOSXlgyCkd6FBJ1LVFjAun09pqbndUTcK2Mc6pB
T1m5LsUUh+mujvvK578H2ZrwiFuwin98r+Sn3fP2bQ+kWGdiNDZn8j3OHz8Al+JBDcvzy2dsSLFQ
3YVjR+p9pXOawrCVzVC7KQEd4q27AUDCh6VKBLw5YrXdJ3snjZxGCeUSZ/l0Le/z5YgjBDR1n0xu
pgu/PskHHquh+vRcqYMrnsZfifVBrD5U0rVkI3lJDpE2Bdq4nLk+kZQJIjfOcfYV+1iM3CnInsTB
yJGErIxBRmKd1VpOGs9IuJgj47zU8IpW6VAptJYDwxy46a7gpQsPZWxWQyIK1GePKvKh8JWZcywy
wsCsHtuSuPwI1XviQIOSQtQ1JSmHG2NJZ4fOWR8MokeD54hsY9XR5UZYCBK/YLNOyecLaJnMyWGp
gRJmV9u/IJnZp9/cXuhjixe33l6ilSo8X2pFBCCHBu2oRmPTETbc46JExpnuIDgYniYNMkxpErts
1vsMmu6grBpT2ZTG8QVB0D7mlHkBH040a5H8Ah7vjte4R43LOHauPmZm+r3eBT4BBZ1Y10ePGEEt
6tm+kF9UVE00At+JGI4rWW5B8cmzSXTe07PJCqE8C0bDywnoVoOIF1RsaiuThQlsFZrMO4xxkv7c
MvyoY1AzCQyi7Pm2yCCRzcbjVuDGG8Qv3huIfM1tk+s+BjkOhq0XZ15ySlyZo1TxvTzcqU1xQbwm
z8wR+nRldgvfX2jJ6Y22umHiGV3MWCnEotHUSAbEQHBYZohnaUKxbhaKs+AHx2QbdRSFwrOfz5z8
XDyN8OI1jg/CK4j/UdPl6p28bcP99rNvE8SzPC0XWjOyecBiB6IknuG4n0FLTO1UIJND1le9pkY6
gxwydi8AFHthNgccP6cBn0tZSgLSq+UUUCHNGgFKhU6nFLZjTCm1EpU80vDnHwA/MspG1F6OIh1X
1FRfhiWhg1KoCu71EwzZyrYs897Xu9qVygA46BYpQP+K0zdzYObnLr25LYf9TzjPoKa9GsqfnikQ
me9LJMHkaUm8x2KkbXVetWu0iOm51jfqNhd2FLMiu6uRjhb6l3RNCqcvSSiJGoy9pJ6lUWOdefPH
2xIo1aQnfJDpg/vCPXJhbnllNzotBNVV+6Uzyxi+YAQX83nkF/4x1yBqrZfLmO6cUW0+xOi1qVhT
947gzGRIwfris1x0op3oZIa33/HBFl9AadgHNSnAejxi4aEN+pQe2DfLIz9V5+f+Crl5ifwCjuvo
Nzb8bbiL2IKoqhHb1OBiO3YZ3YS5nnGwY9vjEacabSSs4vy441M8+VGyTF19jZrDDnj7+dRVF3A7
YgDs1McmRTqIp33Caab92ssD54/XgHcoaQtoGwZGHok+aBxfB0JlqiKTkz9SCSOwaCbAfH/WCrzE
sAZ09I5E6h8QwAX8GqWLDj+KqX2IBfXKdfLIw3iZpLLF2iPjTnIdto7erIDuI6+bI6CGP2KjnluW
MhCnxSsC/qAFPntzxFu41771KaEVd2fPHm+vH+3KEIUCg98Hf7fuElH4RRnUSXpYchSdnChNP+77
KzTBskVoTSUblMX8LZ9hODxQX8Wkltt6UI0Be5PL2nlOTyxp0qK2vmNmt4bkvN6Ty4c8Og6ITNa4
uD1ITknOrbPoVQSbbYdEottiJNJ4zVQqD1WaEOtzDYdTSeTiGyuOVguVc7bvdERE87KqC/gyn5ER
5fzS36Fg/gF4iD4uCHzsmNHP2vivMV4mZQPGzw3692/jiMxOkhCqZy2Z9dgF9a77i48gcHnRH6Vh
n5BrtZK6woO0KI98GJSDBoHLV2X4Tge9RcYk4ZPlXkE7HvdO/UBjIMKOCE2g4CKd3RGSYf3Bn/1h
9Gx7bHSNEhfg4K6PUBD0wuR2d5731g7MRgWtxq3K67MON/guRLbAiUanmbF5jDhUjMtLL6CTmHRQ
R0086bGdQdiwXUYNpa1zWkKJD3PSkIxerSuMn6TogcKX1uE8EVjOn8f8XWolQdeWXs9b9a4/h72e
OD5awsC6ip/cXUU6u9xFlz7YjAfqwYqL97I5MEMNLK5PN+uJX8NKSlL9Nx5Syq3SjyfE8jF8dZ0V
amD1Rg2+oI97BAYILbkCnnE2bU5KnlC/pLydcU2nW7f7M6pfCy6KFDVLsWH9fTvw/XAujSuTkmzN
UcgpxOtLG1cxoTOeK0iAAxFCFxkXHjr8rYpla1TREGBydgsmg44j2J96iAlZ8UjMp6mZO/FzQN7i
xiqWKbOvVzXbB5vG9fqu10EFyG0C81mzKQrbNmqCp2HD/2c1iDR00wBrIYNjyAP9ptDW8FxnQGcw
1dTJ2m290Gt8bpZ0eE1P4Gie1/54T1yh5SEoB8Fyiu7Vcsa+TH6JI1eEyofn7K58Y4+qi9k3MKwS
EdWfRWocTfXkTuNDAZZDWFHePSnVoTNQQzv6pePhj0YDV2X5qQZeeZxxZnR8AYtTT/XsF+uEr3Jw
dAeXBhMQj7RkOKU2aTbMZJyoJW8adSbx8rndMPB4qJhfjGFKhaqhhb1fAs1KvyU8EK7k3Uma1oES
5DqaRUhaaslyJw4voUNYPM1XZG1HVhTRDeeq3jiAXholP9/KH2vVCzSlf3w94GYzvfYABFGCycvn
E+NKZaejFPzRa4ts85YVWxqsWfpXEOAoq7rd0hqh9nI5WnNNfmFJWU6CmVxl+ecxz4k+p46UkMfF
Ake1aCt9XBcKOfHsOlIKdzSfaCla5j/80Nxc/hbSjBq6UdYutn+HCAMo6sQpPh/mHF3kESb4ufWE
Oj8q3iL34W8JILgJt+HIGVRwk+mgwL2gpwCg7uLTuyuI4E08xSPCFEmvOe5OpUOVgWmkZMpJSuW6
8zDeOu6fWPsiayPVcTuIrTM6TZF4UsDhhHi9fqMKhp8rgU3hgiUC+UYu7PKlEUWqzJ0a4VUKIWCT
ZTQztv1EZyrq2MwLqRV22uv+fQo2eFakgCP+ICpc2zJd4cNgyik2N1ie7RYvRvWWEIt6HCJBeZmo
ydZ7NExDSfIdRrNO+O9jMij9ITfs/9oGIGMNr/FZzVMlrpw3Zhj9UaQcRBM89AzXviRaJkQi50Ai
i8RIVR8negTSz6Qq/A4r+ccRrb8veGjyGv+Ggu7dl82bEb5G8t/tsx1aw+xUM80zVeIRUyEqQkVT
/tGFbSfPARGJ1dObzHJ1DgVsJKca0JXThllFVIA36QSdH+YoCz2cZmJaWTJucfDM34ow1OBDXl+X
O3xlPONHjIHFrRR3aFAOcDNEtl0c/IKsHVt6TQFvfrb4ehw06hiqi6TqMpGATC6GUA5NK2r1wMK7
78F3fsPMjbqgGizJ1/UEQbmCr6dT1bK4G1IAYMcmWSfeH9+bU7UzZHJCw8MVIwhllG07X8TDyF2j
GX6rXbcG+AX/DS6tb3SjfesrzGNT22DkeFZkx/WRZjdIfh1gJkHYTY3yjEJGxMt9NC1SzuPv9ND/
En2jMitHpAJo2aSFUbw4QpI3Cb+MlRkoxv8zLdqUe0Wrz9Ep+BofjEEsX0j8G4jiInhyVYUN2bGr
CV0QCpO8yzZCW4SByjyLsj9VyFP+cavUPBp+Wgdlx6fRc4aKIvaTbD/9ccopLFP2aPuICV/2h8Aq
+NfMLR56yyu9A8UEU4cicwHuM5mkYD7VV7YiJjuliGAukw7ZpJoauyDx5my9YDZJBCe0c9kIYVSI
fQb8WrYMGHbow939frQfjs5LnvMGflH/xOmAc+MAUb7qffT8qjtBiHsk1UJri0SaaGrqUbzbIxum
bXMVxwIXYB45OC1FaDLHM3U9Nho/FFmXLZJFEXI3ssxg7dvp1cUyaWgHEJGlqfShP5wvzvzdw2BX
v+Nufn7i7HaHndK2fmodzPGBE4uHn4EQ3y+JwmLYxVLRzrtOuykUQRv4rnA0nhkc2egIraK6RDuh
j9sEbhpoy+QY77axLM5vmrPmDxEM2r/hHDLLpxMTQe6ntP/Zaz5O1tji75EosN7yp0tTfCD19Qre
W+DAU0zF7tv46fg68A2HnSdzcXZUhI4NXxV3LmmFGSV63sD9vjyvwCIaqu7wH1W0gGN5kWJXOzR5
lfpx637LOB59AvRy6/UyQxLqKUU9nN/FMLzu+x/1KyZInCCRCGUNRQNFEO6mgAY12DlULuDNZwwr
cRrMLIizED25n1bWBspryY3jLfTUHvwN/cqjRMoiIFpPP6N2us0M3/rgCmo5gVzNdl7FXzhQtSzo
1zOjWDbDuQfmDdnc3Np+JdTuwY1UgNaM8zDwv1TZpOqAAcyVUQR8zvBNmI7jyUoqi/BuM1rT5024
HdDpnwebDpjOIf5t4olKIwKg5NqfXXiTkLKKVEE2wJeM0FSHqEt9VBp56QeBCXnabeu8TSoXUywY
6EviAXwiEak85vM67K3dhZCt6AjGIIsANgjNZ4IXKICS8o+MwUtdSkZ8rZ2kDuKnTSvKFoufRRZ2
oxIqeFFCbFDIZ4Na5phWJUtuMMlcMr1Uvm65o5Z8zTxYOuB/0x7SeYyjUvQz2jcLD8Wu3JeQZPyF
717Fpk3LdFqzjYFGbFwGWp8SomCkBdt7ii5fgTgydZHR9PqeYY4s5D8mg/uann8qrYPeSbeK+/YT
P/DefRkAnWFuvOgXQ++vgsMma3uiOAuHwt16ImHceENT3ZNPdLDUyafyI8b5/ASlDdwNvtkiEUO2
N51Tu9k58YsdwfbOz0EAjO2O8EFtYn29p3iX63LFu5d7z65UKKGMg3a+tgIqI4sZmaeNRyFECydK
ZQBriYmOnf9maE0R4Fl2TmbBU5ZYQ+kqBLF6qvpomixfT040SW716gw11GYh1+2rAay1lLp1iGbL
0xgj9Zh0SlZwnazZ5ICKtSS1ou2Y25kq9r31u1B43LQQvQSKnq0Gnd+fLzmDPk/Qa84w6zMqlYDV
SaJ6m3RWapA6MOKye7nvBJ0qFWQ1I9Y5tKJ7EEs4XL8Gd0dR7RGqTP7GdvkAqQSK7LhtUeDAw5IL
rlohfhKNhwuM61k+I16AxI2vk4xTYFaAmXjGg0QaiKg9pU+sPqV9q0oPLWYakI9LuSDUuAOISEs9
JTNt+hk3BikDtALZHu/ozZjBdn+4mXdEH/vERc5PFx5y94K05JOxM7kO69pKKeRKh9s+puZN3AUG
pGRo2VS0NXc6kkrX0gJHGIRKcnl90JFwMxM4Phq6jky8A3EvqTYaJ8o+0vSy7tFzN2NkrVVs7Avb
y77V7loHpYQb/edqV+0Vn7rXznzP/uqSiwYRpFsKnsAZ3jqgfHng+b7QNykTgJD+bJ6IsY6rnd10
8aWW7SO2Sae5cAE1hK8bxgvvRjodWCoCyjxkdlSV3nwOs0tm6WQrC0f8mtUeUJVFx0enyyD9LzeL
zfWxWYOJh8FzuOqNwWZMFNmggqgqhtM9zb3Ga/spa8vobt2HshoEl1XeIYZTTRXON0QVh2uNm3Zq
b/f29aoqtgdu/e/+EYSPFP23of+zGgepooPJA3fL/vZIPzxNoPDLI0r9S/v55VkLeNfacIGD3del
IXwLhYcOZFF3QKec66A1vA9e0vRHpam0FlILh+kzi7qbtkcy7TWF6GiJh5RbuitsRLfI8ajdVcAP
AnlwD5DS6GgAC6HIPp5ul+n0o1ZPJHs6Ez8QxzQUyiCcdQO/le0bK1N4J4Clf778yVgbPW9nyuiy
ANiMsFzYoDQOUJP59p5Q2haiBmg+MeROblveP9LjC2JfiYp0wMJ9trcQKh1Z7ryAQylEZUPV98fH
rdmcFUXMAvDRYx0F8MtIpJ65kmyOcmVCEOmHs0cqmyxYeoXcGc8UjoRfrjpec6jAuVRGn2wECyPn
RsErxyqExaLum26kUn1Wzl5xGn/LFQBqU5P8f8wg2ahNi2CI+Ujz5WYcEj33eIFh9Ymbl8nrP5uO
gJU8YTG3FVZLtKryu4NCOeeawt4CM3jL/xnXEePNLFJzkguvanTqXBahijZH2LwJ7ZN2v6+n+orM
eXv9/OS/Z8fbxmDzTcH01FzkUgezoPm2IrEdhAG/E9oJfqcAT71/w/EC3u2zM7tDAk0BWzeM3JRK
Om5mYh/DkWWb2C93laAvD/9RDdzkpyzHZP8LPiSPitLc3aUeCOj4ISlYDWRqUWyQqgVMGpvNHnDw
/nk/+hqt3XgOhWEw6dFOXLQ+fEXx8yfQDjDmBzsYOQESrP3COQnZ2RBJnyqc61FvX51CIJIo2MAf
BdFmAUzF/ugteDlAnkYIFvN1ikoSpVjQo21vUX3dJ4S6hWjDMkG4H3Mr+MepjamWgd5Rcp0LabY8
pB8UW1KAWomOsqwVjckwYNiMZWBicV45LF7XAVJ7/BPteBSL+MSlUfOs8K6Qz8HyCRyY3kfbz3/n
r3goy38slUrC19XxTMUKydPzqr3rZZLN3jCdEB/3dE0vwiFMQbyhdTP2BxurJqkrCma1NJjP59hU
P2fDPmPU+c6B3/6Ppm241BKUd1608YUgJ0z2FzFG5yer2nAityUrqtJXacivbektfvo2IgioxRpT
zt0Y4QW5XRAziQsNwT7KSyqZrO15xh5AQar6vyN0RPlGIqDOQoIyLgFtGHrWtVZ/aiBlqluQ4Nvp
eQoWKtBt+E99Xh7wfwGZ+ltivBfkFngTB+caqP23afwnn3r5XALwTRp2/T7SEkIvgjU7LZgsK8ld
TM1s3zfeaT2rxES9R7MlJbpJqYUi8IYauLS2eXEMvYNXW2qQpETxBgaZy1KXTYmxYfCMBmOT8GzJ
KDMsPtX5pbJlXifaGTfboR+3A4T+L5/8yw9KM9wp63vK60RAbTnfbKWHACCTRjBIuLSyQds+FKDw
dtgVHZ4qNfH7dkA6J5pgpQKLl3z7HL+al0ns1F8krOAc3mkTFxv5WTsUvzKyieIeruxeSmtH+OZX
J8A+pjkYHVwPQYlCcUFCep4gUDciS/QPv5hjplTj90dyiFK1EEly2tilUBR121+yeMKZgQ240kUi
CuJ+3s7KaHL9dlZTG9+6RQC2Nj4bhHZ0cmAXvVGoJSkNbOq8fxqIU6ubJ21TjEjU8k+WRtm1MZvy
577q0a7+SfiDxQ3SxA8T/7lEb6p3bgPBeAlENoAwJbPoiYhAMCSTulKGgMSWKCf9kNSXEZt8NaDO
3BAcfhZTWqIV4EylpRredB8hRpo0aPHH/RY7fzoeMqTmd0YVikeAgw+FprQawMdWmyakkSjSFhOu
tZkntQclj97fBViwGzPAJf+JUwASnLd3vV8BChykhSHW0bO1nKDrmgoDceODVpLefNuEssJqqIDX
n1Rt8lv2lbAioCksBOmmupzNMkD1MJsPcYq6iW85kFfxjGNUbJVxSYlQUrE2R0j7R4ADCtvWVsxZ
QSP+hO10LdPE9nOUGOjImTVf30AzQjaCGtq4/yJS5Iemd5kyDwb8HiF8mVHJBfyHoMae5aT+Islu
zOqaQY0iJypLGzyAZLXGidcqmYvSF1ayWohhluNPV8t4hLZ+CV4XbMDXtqME4xQ3hRb5Ztv36nns
+k0trMoUn+LTuM7VIMAONWcDDpHjs1dNF7I1JWYoS36KuFhvHnj/wzPFVzyirVBQCBGVAfc51mBi
cwffV4X+shctU1yb+EGig8RcwEem4BwQpMplHdsE1oBm3Lh8xVlz/GeQOYMesiVIP+O1Q6irkgQn
z3EiZt6QkWH/7Mse1s/mxM2gacaW6AVH3nwSiYtijAez0dX5VW7P8hlaO8XvUY9rKHVeJiGKgPKf
EkR70ZqWhwaGRv5p7w0FbNcXzFo4YrrK2sZRUdkEdFBsIFSbI0Ozhx9ncsv3UJwcMjP76atZn7d5
kImkflODch5dMXmVs01YVWoMgVE0FnihwnL6zb9WIgUnqqOAhDXsZs5VqzeSq7bfIobapVfdy4lC
07OaruQIQU4Cyeu0jS6CFjTwstkPT8gYBfiUifZrJsjCQs+LM3boKqyd21D+ManLsKQkboqS2itw
1pK3vwLgU5odnURC+XoGkWZJlgGbzVKsugNpPjPahKHtdganPVI5kf2GuIjUmxMviFT4kQATwWEN
B4rKCDtS9iq9QErjmg/ZF0ZPmtMIqVlwDVE7EUSJEgGJ8Kce+faYRkoSnUE/uhAtQXAeWgGUqq61
C/5AiRVO9vq1Vms7uNuI2OkHCHtWGACxAyh39W8wit7t9AZlsna5QAugZGTiKF8Uu3LFOC1bt1zX
B5fYbfFj2Gjm4uLqPeAFCcz1ZnjtXqtdqR/foVkKJxgqwJUhNTHAhTeNu11+e22uaR/FtA/CoNGw
ARWdkAPdWQaCLmPTNFnv19z/C0IS6LpfIIz5EB1lSzRdep13mfxsMZLACA8WhCyVrab3IIfMNSPy
J4edyG43RtDDdg1jHdSuixXvE/5mPuvy+mLppRIeVhK5+qrHwHYiSTlytRRRQURoa5OsTBCRxSK6
zW6rPhrGoV8SZN8F1cJKCWexA1GbKGoDN68o0r/Op/labOvIBikk07MLhBxJW7nN0Dg92BRh55th
fk1c8Dxc9aUOHrg+sSBrJFxRGv3sfj78f0kJMPzFX3bPXtRByvEqQT1YwdyWYfHwpa/QTyz6tpUw
rbqPg7XCq+RwlbL9zJKXdMFriCEFkNnA5Tt2fjofk78/0/CE6Cy4Pyv+gIlxPP67YvAuOJO6ssJT
n7lrer7FWUIClqwSnUfnDhwnIuiZ7Y0pYDbwFLPl07AaP2fuqfCF+BL08nA10b554+kyhxBLsNaA
Rjn0aSw1sdA1mb6YE1l6FHKhN70M4xzzIPthBrw58bz/MYwX64IszQZFoSvRrZ2aYuGriQ3aQfvK
+QnbOq2qIEkATr8X/h2tlbsCiRJ2XiGW+YdS3VzgObuilPeuXOe3xVrF9ZaDCT3FwTwG6gIsngmh
7voLR1mXS7et41joAmIs6oiniL3iB2l4uYc5ZChzXb3ROvSEba5g1blRDnIwBzlLyhxomYBS0lgw
cUfU7pAWhro2/9Ba+2nGj58w+pMUo8cBxtajPTvll6LejcNJLAUI8BZlmADOJaT4AEszLfzIJzjm
Fb6SIBijk0wP3NA1ldbZCSfZSCnA2LWfkM1Wn6ALGGqjF2De/Ugd4RTBkuaKK7zOPyUHy+29mUUN
kH8v3Bt+MarCpOYXhuU0Mr0ynVWuWFyvjzXveL93FYhsBV4Y0OiCE+xRO/uGrF0Y2lApyfW3x4Dc
syXa3jV2Yb6I4zvk5F193swaPsLmw/93mX6UQmu3A5iQWnFJLJNetBuKE0twVkk01twgTMT1P+iU
x6L6LNn1M5+feMA5RrKc+ESjHV2xGlgEmOfqqxoa1XfFyhmGTOciehnyOlgKGSixruarEnlBT4zP
gdkPuZ0rg8e6Cxe0sbsB2leq2MKWZYnTMFN86ky3nD0IHQjpyYqiP1mZKvo53d6trjcbD+eZy3rR
LWGwE5dM0sF6uw0WknguDSVthhKcMU6ErfUb42h3DKCFu+9m8/aS3pDaDW6bkGtQ6t8tL6hIwXQE
8Ja84GT3V756KRZIVHo3ihOzCfjiuH8r8v2UOCGWyb7LvSV8ZFy4A0OOtwdjR7Y/Hjktffd4ElAE
Kj0tnqGu0Ndkkxi/oW7MmOG3t81AiAaD4RW797SceriwvmMNRHIhgKsSbqZb2ycexKJ+DcpxbA+Q
3bUcoJK5F/XlJWTul1TxS6x8qnWqHOmi1HtRBV0l0oLjnBSKgwoR2EQordSvhD6wp7YveusYxp2N
xs49kkoRJrSZi8O0HloPcg6lgUngWWnJdz/BYaTtDZNBZGJdecBVNs2ZthkMEksORGgNPIQ0QOXs
R9i98nt7zzoIjFSC+5ofwC9MEWeA+lNgf9A6AjJCDpIYmM7sqsMqnjYCJSepmjm5bIEH7FtgOEx5
ZshghGU13xx5EXi69RN01aPz+fLA256Xvl4ebSPyme1aaonIDVY+WAkU++kWMVg/l59Ig6fV/Zoc
vURoYVQDrxZ+BdzsYR39HTLjN3SlvOFmq0CMAA3N9ekPPFQaRZQfNKq8HNpJIWkfYCmpv/UTVSsZ
xAkiLy6ysgNVqQFLe9o+X/Xy72LY8w3T65X/mI8hR8gg3dYXTcCr+xtYxsa4qvzY40XshoWv0aqe
tJf4xABmbVzqvROc2i5sTPp8Vwe1R22e8+L/GF+0hsG0sLGqQh3d8RQTBAOkZ4ov3eT72vcST5p3
iPb8gYS8+FZtiE2lkfxBvty5KBJjU8wo/U/TYw3Ic4kriFB/ew4IQknuPXcP2AvgrSa1Un5WVBKw
1yOfhi5O/wgbzZRYaTumxsJmo2PiWk+EktyjWMgVH5B4mulvsA6+xnALvJ4Z+5PFi9Y4R5nGYp6y
VzsnyeM9ei6WjWL+vN5mZMSCXjhhuHyQWHRP9rhfQGX6go6b1fCdcBHxyRdDKalK5tiTd1Oy9Fq9
8iE0pXftR987OefV00JyzBuLeHw02XFXbKEaGLpQJTcDagAajAvef7VV0Pj4xtVgWNwb04KIKlok
zQNzHG4uitSNuWlbuTvYDFAGmUfkNft3zxSEsMc2/9rLsUAA2fs2aFeosjBhuokL0HkmAPXycKHJ
7sSSfeCieYJ6dmpIRkRVW3GmCueSpk/a/YaZzW/OEv0Fr5VhBn+cdxCNGhJ6Rw/LbJWto1iG0Wt3
KDBWCNC/DJ6EXgo6Vv2VwQgeOOZHW6kqP8h3D3453J9dFhEcOt5VZP+NJ/TuIpPa8qj6GKXKfrHE
vieLSQM01xz9E/YuUEsYkkQ8zxV4dgRvZsbsG0trtLvqA8gxfsh8J4S2hBZFpAoz/nHuESNVuuoB
QbMmUJgZZezcxXwHlGBRwseOcquTlO6f6Upyg91o3VutrSZcI9XsgraKsSvjCdawsN+gGIhQtlQu
Xv1gLR8y0eHJGpTzgIQN6Z0fxI6h4RfCLhn40FJk8xIEKOAajksA3Gzk6umbUdoyDXLoqivjgLSE
4hDWDtxiLaGThxTIZsbJd3Qn9nUc3nR8v9NunPWqRTy26Wu59lwcOOsQ2VSPSpAIwc5fApB6A8If
zTdrGH1RlsLrXIe/sV5txJNi2UKDa2cPMHnrpz5EiTjGtAXonsIQHY1pYc+jLD20SPxDxkFJEDBV
sDWtpZudo9w5nNwdpDaCkiB2hCGBrgddMI71GcvSgHoYVBq+iLkv+zCFbYQksf7//9qvOwpqMve/
TNZ5BMTz2aY3cfkJf1wEkVD3fUvXyErE4bWNUS66PoXbEY+PQgBAZGXPmOiRe8dUuF00q7hi32VE
5OFPhNJHLRm9pgWlC1OZKAs79Iftds4RkmOK5C+pW4Iv8LG3Ir9Z0nVfIU2sTGRIJq+hU/jgE+HF
Pc66DwMUaYZu1y7qIj6oSMLDxl0ktciXEGAeNIna/tTTjjIbMBv497orGXwYImxIVmZGFn0SlolV
ELYjxIVWRgjMf1F1MsBkwqqXS3s8xRyp7RPd+t0r9uglkJ/QD/I/Te67mfygkqF4T3SgCHyf2suW
HsuPAi2Hq6D2n+KRySoG6LTFJMzhWynSDawLQVyDk+Uxoy5fYMgivlkoQYbGkhqX+QznZ9Qh3S96
dXNOLq3sMw0uACqsBUxRXSCFu39h3dLyv5cAOqnWby7VKE3fR3+mRlmjyjOYWGuEfICe5Agxsmn6
Z52QvJYaylGT8SP2n7OyczIhTFdlxlwlxb+/1gD61jJE9KAHQy1E4XzINsZDv+DmEl6exa94v8Js
CqglvUjQWBH5aMejAl0X78zHm0lzExw9vfyrlwzgZ6cxFMtSPe/DcDNvxEw/Fk1K5bYeLb829bxa
vSgwwkSzwAPZ18HWCATz72q9OHVF+zuhO7tJkbPnXgO4DqsrMObyuIMSnQ/ZURZ1KlQhJtva1yy5
uC2rY+JhE/N285Onx7jVpT+72kEk1OTry2cS1cIKxAf6WJi044C5GIt3j/+/LZ4TnWOZNhWNQPcL
ylsfZKyAO5pF3z7G6gSnlFwsuH+zbB1sO97n2RWa1Rm/2TEbHJPaVYu6L+bK+rgRunxlWfvzecw1
2vzSnBpg/n2a30hUhyUSNVTPG0wgCCTmnLqf5udhSLmohVA7/pncREy6NvV2f+QOSdXNgyK1wspH
u99DxJB/lWWbJ/B6k1xWVgKUkHPrJZMhZPm7xt8aR4mGCYYRiWqayNUQ9X3aN+Tm0nWUrQQ1p1eb
EE9HTqXxbVOAXbcoj35/DJnVSPH8J8IFcxsy2pzTOWm94LSoO5LoaLvDdI0IKB3rNsLibd/SjnRH
pHF6+w6FAddUf9ybf0EOQcimtk+NORTFosnsxxOKkuZ+xLkyIFwFnW4npGzB29Mi64CoDLdKWpcz
cWgyGADjp4YBAX/l9uI5CNjRsxjZA2rGrdEQXvqE7nEsJKnl0kvzYuysE/FwubcQ8nAuNguQ3rFJ
xV3Dr/O+TPfp4ocgPnleUfsRk+gfew20e1hoyMG0/QT+oJmLSqK6PuyDQmRZ5o5CaEeRvp1PhKfk
erAHpUQBGCBEErhCH32Z7L2AyQiXJHDPxeGCc52hMi4PqGwyBRTIS3kWgxuCvql1Lf1EHdvYuXwy
b9qYqdW0/1KvHRmUYuVs2jh6U20c0mZP7UIg2APUqeo/cya8pNBXOe997RF1qBEiHGCOx/hgsIeu
uYQJZplvmq+H3H9Qdxq6ti81Da5E4l48uuSHy13L9tSObQd1hneDI7t10Z003NlhVVRMW2i78IH1
xEygS+BcqxMnEr3tI/vN9RF7ZLGZ6eZh47YJ1p3HWA9ygLm78rTEITU/5qPIU2ENsuWiWiZa4NHI
YJwB7mbLQtysTaJGw6NzoG3RMWYfxdoQZMc6kYHewPJIYYRF3Ql0zfjfwgZds/0iJDkxMqLnxzJY
jb9w9dn+nFZL6Qf76Hegr8GdTN4K6sJ9miOV6mJNLLOXuuENmpZTZPThrkckPG11aIG4qxP6qRMQ
CZU+z/DmVJfC9+rvB8mS5S5e8elLrn7AtLKwvNGVC+wvw9Ty7QeSQPFLa0LoUCTlrNleJX88WoN1
dV7eakXOR8I8m9lBRQQLATWSldiP56RcLJ4/exRpR6qd8kUpmFjtmpBQWG2evpGkNJop3iTOk25m
ZRkpBJiSH5ujYNbwdHtNGwvcn7TBK4IjnvY0cQsTmcROt1dm14kDzPwyaKa6MOAbEckVzJb0zi2Y
LMIYegUD4stJgTq4Ecawe5vo1AJU/uSXhvWYd4QeSvFs/1cbulvvn8CptxmAYkY5vFQnI3lgXRdY
391Aw/3gqNF8WHw9brKfFqy2wJ1S4x8hrtCwqQsphNa1WrenGMIWqL7JBi4fkUnfa150ziQWUJQU
a5fItR+1sBGr/z+EUadVVUpjyiDWIST82wVFH7oDkP1WS/U+SnIEqanmvN/NE6i5mUbyuwLRGD30
co8y727akVLOde13QdmDvOfg8JYi3D9QUeA/7QqNDvsVh1VyM19sWeKyp7oJ1THE+ajVmi0giPHO
IAe5culDlUJu7rlyUJFDpJUZOZXM+Odf/+yyHC5lhGjA/ISCxT/CCqe8KkUtRf5IaXIjJ3fREYTs
I6VWOD6vw7DcEEGb5p4nwt2eIUzYrCAAauGzqv0YGr+BrCvo21Gm6xO8x8gjmOJSFF30mecynihv
yO8WzaB0D012Ivj/WcJwtmaSWL45PGmerVmwAsRYD93h23/qUVBNoevwfj0aIbvMtVbFkLR481no
bzYUaTDxThndzN66EhtZcNqx3T7KJLhvGcqlbvzpqDvuv0DV66UaISpHYbG/6O9UhJxDuYJ5ispG
GQLdE5ywuHp7OZMekav400XKERI4Bp/3nlRUZ2vbMdO+WxjOrA//XzU+DtqtYkEtHUHi4iuYX2Bq
JRhoiqu0+yQZQJNuY1LxKh3FTyMXaJwTkVfQBQPNBCmpCGmy9PDRt5oxWsPnV/r3iYxVBJMfpwRT
/MRWK9O4+5nPOjdmwhE0KQ0p9+oAxjJ4yi7iu8wDJSFT0FrJn4hDUg4wqt6LjFbTUxzd/FxkU2Yt
ybOaWAFmFe/RcokFsr8//q0RkJbOAXCvP5Noi/Lf3w0HI5Pf+lF2wfO9MgqNlLWha9V3AVQaKaJ8
w6rj0JoEYQaIXm/rCy7ujCqIV1Zt0uDdyC3ixuzZj6LCHv2kCHoGcH74u9cCTu9KCc3M2cKXt02h
ddXYLLUYPAHOVfVIrcty7DKhB+4nCFjLDc99VcSTwuakOYjsmRDnTHAPo4+Uz0f7NdRGV9ftQNT+
rWpObz3JvWxr1nd23P6tsGM1MuoxGPqeo5BuOw0+mrHal4A473fC/n2QtSoMWstB7G98c6Ylp9k0
xi4p/W6U+jGoQt8EOcRaD3nsLsBgZsvV/PHbQfnyDPxeLF4hKXbgfYIV2EkTcIyWqAfcJ82rKbOh
mugxM9EEXlwku4C13nsYYBS/1/Jyp86wxdx+Q79DSa82OAvQKPPKspXRBD/UWLQmvHswj0oyAj9U
HEmMSKYIwh+slhlvxlNTtrVQkMioVBtK2g8Xl/4A5QnQ8ewvxnjGllLBEIvQThvBhllaxVWpwU+M
oHThCcUm2mZgSHH1fYFbvD2qXwnUC/MtyDuxD4O+KqM1XXQ7qchocEELrElKmy8GxUiIcVu1+zip
LpBDUEjxNwwJ6H6rJStncqqp5xhzv7if8dhMV6AK5ApisHHPAzhMIQ/eKoFiuGi9MnGS4lJXkE/S
qbctDK9WqqtE8KSSxLo0+eq3SoasF098jzBRXD9nOfXvJzNaDQq2X195wZt0f56e6aHwkcOB7QmB
5cuOgXtsmRv1hAxnq3ImPdPPmxl/Zbowi0y2ed9B71f1ftBV+7IYmiarnY7esahUSsmrf3ECMC3/
hX9LN7pZhKR/QfRcxoGypihMw2PeRnxpQAtWa5VWSHu+Tcr0IoiT7ETsyQAoieRwf8lEgW3rsN/b
ychhWO9rUdwdxZ2n30q1ztID3byYrucpu0W0rBp8KmXS9e/O3VcgGFHilsOhPgoXn9HzJictGgdA
Q/muieEv+UVdzBXqi6EdKYh7hU6x0Xbzm3Sqlfre3Pa4r7EjFnT6BZosVed0794ac4KgpcPfnZkj
UGQdsvhjE2VJd9HkYymLuJkZyXIM/jEZ/8x9esZGpQlJ1jd4ElmhOtYwwR95OyjFQmK8jt06XICC
5iiatZyZRge76YsKDePqek218kNfYnsRlyzIri9EEEQsHMrVi5uJiGz68W946adbjDcPQ+p9Z0GB
XsBlN7I6HsVasY0ljfPJOjrBiiwHEDAXA2bU+3pbr8oSPRY+TzJJlEibwQfwcLy9u8qrS6qnV9Uy
19+N4DGKn+fgRxoSrSktfzaKm3JGVGPeyITMijMv2Ue1ZCKtFQIUrGAyCQNatYSavh+IvpNYxzfl
74l1gs+Z0sA2UbJGxaRcI+LqrzEwwLPJuMzl+bz04SmP3vB5tnmMY8MPHP8U0X/29xBteEgIBhCG
B0EF5E7mLG74br5GNoSVLywRj4NWWnMycTc84BwGhfCNEx8QiHtHL/qqUpZPczXL5UF/ZXPF407w
yCMM3ZuWRpEXCf6uPzE7y5muZ3QtHW+0iFJNJzO09e/04t1cGDGhDK6fAKIwdNo8NJ+tn92yo9e+
lPrE6oyDNBI10VVksMt1stMLi2MgJ+bF4nm0ILE9NfcHcp6wMF+/JArgCFs/BG6Dxkubru4BwIUk
IWGHJ6TQ3UKQka7V6QHqQV4vDRM3qDdOGfGMxLZ3Bn07qJFPkqdD7ueXxn4lfvfrS5nVexVb8RvH
zDSGiK+zQIQg/xd1CGrabSVGIyOhYB+LsBAhVgJqDiLXGwFXjyeIBpEGjqYZdMuonQxQ6lXaPmD6
ExqOfG2fV1Quh8dI32Au6/GSuJG/35a9ejrbUZ4zuMNsgzpt8N3Qx+jOzSinCgLMuD5JLxBgP7x4
bF2VAuiQsz3pdWRmpd8Q1N+GT7ZUWufNZz+1W5U0t4o9FNh0fmNFP1eKoilaqVmIYQq1cFxrEgaj
ZQRP8ivlnuGwEx8SVDi4TJ8DE2IGHcKBjt3DTEkH9rGCY+6HroFVHRKk2Y0SaWqU+2uHmyF9KVwh
q+wkHYx5fxBNk6OsYwEiqqpFDVjQTupAJEMtqZYO1suFX27iZFIB8HNuS9crpHm+Bu3Zee0dbXae
KAFQ/I1Q+rWfsTFcmu2F8pAYQTsiL3W33XjU0ZxEM51bxLXe5YzU+aBZbU3G+2rgv0AfwWYHqIl6
4LLTxJZujzCcDtFfK8+j1jUGbTygB0So2NoUzN+M+6tAlJd2rWC1LcqB61hRCAWwsi/hC45d1IKu
UyqEf3quL77ielODHsIm5qduDOeVsnflyksEe6u4wUTJWJ1ypo8HH4mjyiZT/WQ51B+RYwZLD3HM
+fhbJs2IblbIPEHc94Jsg1c51DOemuEOAmPS2nSVm/LK7ALu6q6wlZXJ9YtdyLsdY0V2vUjOIjgJ
ylOgF/QVtAO0P6/EDksnVbTEm850OsIa/sjWG/sUPQrNH5hEp+rhc1UW3KlvIttJAs98V7duLtsH
nXUXKQ1FQYg34dwZjJt3iqAiSKrZTcJ4rpvUTsMBe1th7mwsrFJcsVG6i29bmF0wLc4TI0B+54Ll
W4WpgxPbbMZ/dJHmn6jvtVGx00ikVopY2hI7pkwVGWZMiyvXlB6SzwipShZZHq0i4xGpMTyjMfxi
62BOKzR7qQM0Dkef5hurq8eGoxqTUdVpOqnajjG36z40KR6mYrTDyxWOBZ6hY1xN1IhSaTsXlbws
9r38z4Le8FPN0wjiHdNqfG2SFU7vfO+tPBufVcLaUMC9OimjMzW02uacA80lF3uSTfPFeYUi4ZR+
cymwjBzVTObEmOcXma9mrLs6ncv0XE3jiFldzbItIDAg8OJbm+wn1n8Cz7/PZORbJKzlap0HbeJ2
FPvqWhBqBMSlp4t/B7vxikDfKiIYlGor07QWKF92JC2tC4y9d1H7LvJkucaTszsUTwkwxU7K2EZT
Ft66nU0ubdxx1huKsilBj3nqnAShgLvcjkphUZyNGPCABd1vEDczAZR6r0HkbLjJEmdQkIO5Z024
2DyfZuyA7M066rLF2l10HuGYH9G76oJo6z0x0835ymcaQyOXtIkqIoPeS0ToZf0fVgQlWBsyhnMX
XNXLhmIrIJAhlNSeJtPmnAhLLKT2r0gdHEFPXlEcekRuknJd6cNLNvVGXx/tM66wZYzPTbTMXRg1
6RmqjcIeZx59B1P8q15+wjaJHhVy9qoG2WP0eYkJScJFmxqTRsaZjmJPEsW6Kmp+J5o2bQWR3yMJ
cdY6QTAlv8CyMeBJZChEm37/JRzAWMOoJT7wNObxZB6Z5YA4cEdpGdeTK1Y+26ZTK6cmvyS6NFhJ
byohoLshupx20F+QiQ33VU0d0B03BaYFrYSSqykyPwFBxcbUoXlY/LRv5T2zsVdgTePaO6qHAFru
Z25eLP1SsSjWqFGhfmWhKuG4mB276GCojemOaZukyxNw5SJXorvmkbk07FNqeGCUi3PQAK5RKCkS
BTpilLCCHan1WS01ZgM/OJLuJcCI+gJaWe5dOsp5gOq6DulICpeU5t/qnjFXwsCoSei+e/RknMis
g32tTvIwrJEf4fPwMjT9I+w2MXD8yKGn8kwVVAeHouzD6rQkYAQ0a39138Ln/ZbaoPH0Zl5NLIVf
Izk7nrRTTS3WecM5ZwYICIF2N1zMwVQElZIxziSOYB2RhfpO3TQijXbfOmsFbceS2lyAhj/5/C4z
9yA6gUVatPjUNnT+KSgjCjQOLZbO4I4TOmNi/5EqH4NZGxim1yIJz/QA8Ffz7yWDLlKRw6+AinB5
LaOk8uKRpXv+/gj6OFWTVeVRyjPD/5AarRsR26ReSvJK6jZdZChkNgJjzT99eEiLu8Qa0cCeNcof
i99+E8yoo/PwtMjmeIMv/MizxwQNV+2tUS8jqy2SQrt3GdAvSoa98tn8TVlCY+n6tk31iG7UqJrO
9CZfHEezQXYcmr1HkTL6ntaJpBv8PtMvzW3FLRdlsF6Zu94xcKSHsAFp0aOLiXfOqxqcWhypbFm/
wdDvdKH5ou4G0ICzpfbIhEI4ruwOPGBwL4Jwp1y/3XQFM8yrXW52XCdFYR0/ZKm1msTa8ZOnm0Jc
ksiuz2DxlqjIgF4J3AklZ5Z8ycmkizt6fzo1vWFHZH3KRBnf4hcFH9RhKCS5ttbw7z3Y2o+2jQzl
Wy6CsHnp8b52zxzhC8ZjwkDivILNtkiAg5j6YFpOrKpklSm/oIK5Us9WJcKidq98stayIWu9z2r2
19eiXw5rrftY5otfuFS9XkkbWHuhXLLxBjFwuWMpwk10SYfTq1849UhT3TEFPHJ7OZvICEZ/I22D
w7Ex0UPaEoyhEVJ4D55F7j/gKCiFQogHC/zc+dKZa0cqPznyezn/LynI7AGT8arDIPK0gRCqgwzn
tObbytK4PEqMiFJNi0mhus/bcLytFsqrfuK1NVf8/bvkb++WypIv23C+1KsFqdqRWDjP3B+5fvNj
NYpuWOepSr2yQYOnPQmEg5WWfuwFJ65QOiESini5V0kqKGo8AiybgUylw/WzCvJEtpuDbICTRV8i
/C37T8p9RAKHmW9rvxJYnb83LsjdEUn7TnCxaM0Nf2kUsNFECd5zYDUdQQCuvXi17A7snvTUTJfj
9Xp2D+Tf5ltH4KBzI2ax1ZxCPTagwsQA/kwUATiJEFh52hqMRxVFCq52N2a3CEjW3t2tjobO/PEY
jrZ8CUghCxV//aN62DtWozNefzwg9Uqh77yIF0O/M4YiSpMBTdEVtyc3pQZeXmDF9eAI9ScG4pTB
s3xWLQn3kRQo+GQ5j5R/dMSxdTd3bVhpGDTnmWu7Vulfnmqs8S0V4Yy9CflIuFnbokE5j/cskoYB
uUNwLi8+6M6wlpZpO/TjrkL9gc/N3E96oZB7Ep83EthbYDO4HZ4IcdcL3mtxp+7iNkojOFeSOCXv
4uGbgqtqJVh+HXfxShSBx4QagPgkUgSrYVFj2USQZMQy0UZfByKUVmtIFxu8ZnrOnokkst0zuCnl
p3TBQxUGi4OOVEkoUCbJW6vKcGv+WIbKMJleNdiX+5x0hzoSL7MIOELU+GoMGHmsAUWxtL1X8mc5
LR8tjFdWnYiqBZfe+hZEyCr1Fp92GEZTQ1XLDVDvpS/TUvt1RAshFokCtrsSgZ4813bnDwLRXHtT
7N00IoNzcZKsW873Ml5YSHfQ3wBxHB7dRAOhqMMRtPqrSRDf++GfVt1dKtQPNBuHPWeiAq4p5h5C
fC/fL5yqpKBX7REiEEQGuuWTifSTzy09awiZWaHjskxXD7RQWSGZx0p49fapFP3Y6vikGA8I/ZCN
QqVtlbnMrVRHOGl8MlkUVHDoAdrCYnilr27y/djoYm1xDDzM8MQgpUMK+fgwpVYvMVQqTQABwmKp
Ngu0smSz84LAX7oZ/hrtiHp8gPzQVKqk8Bzr5QN93ufNh320YqRVY1Em0cad1kG0orZjKmvw5x8U
Xjg25J3u8seSvVhflTUYB9TZ0Gbf873rO6PTLt70X7c6pIFvokIzXBwZ67454xJmrd/DxvBvplBa
POzZ7g1CM6h+yAHLMXBlZGTNOKTOzZGJQ5fOEG9xpGYYqRqQLC2p82WQJj3SbM9HHIvLEOHz2kyZ
o4pmU3OlBo5tPpY0CueKGfP6FgbhzOBHfqsVYG9n6uLpWrYtEAAkbujD5Wgiz+xHYBuY+6DnF7kK
HSNbsotUYDylVMCETUC3LvxkbWiyxMYnbCeXYjVDae+4WsZO8e5QWmloPRj0uQk+jBvl+YAvOHC4
P8h5bhTzLKuPvhtiaocfgy1yjJVYXKp1HBwfh+6Cux8tvPlKSAgmNAvIfd0vqw2DbETADX7dXuXD
HryTqvn94rH+ol78wSKiDgcBP6BZEsswgyG8E52zB5PFehfb25pE2lOCzVphGPgUhh6OMb4lBBP/
revQm850jFTXpXsBrIY698NJ2UfXzvMw5YTfkvDtOcvc++Kni9+G+xnfOLL6uL/XTWWNLrzDsg6/
nVKDYcQMahvbj6em+S4/8YxuWzHdsr4hFpB766kezM663LXm/PN8U4yYdAm+olH3zmhIz3HkZc5U
EnhSRldvhvVhYuvpJbrXEdUSRjpPtYBwX5eWfdjG+We7fnDzX4+F2FFhT8iFwXe6qqk516uYEcC8
QCVXM/F030YVVVGDbTvKdy3jPlsQcMpo62p2ymPWG4H0VCT8i4iROgIIv47wBe8gjmN76CWqGme9
CxARCiYe4lmIHK6OdI1zJ19sBQ2xJL2a6E3bQ58HGBIjjCcnBxiQBLpoLU8mzibgKeMEfLSsmDYJ
ENQl9B3Tld5UXW9msqiCwkaWQzUmnK9fA7y+/eLyZPDNgow/y4YpuT0OaeIfM+NsjY/Cpb2CCTuq
7wQfRpUkrCp67yA1uHxOTzDD5cfwbIjT5unLT2/gfeasYFOz5vsrDj8TlI9sB+4x0Z44mjMhlfBy
SW+Zo0qgoyn32rK+AsL1YORqmdySFYLYaVhlgReJmOyH+sVQc86E5dotSEmG4C5IofJOiCNgHf0G
zhHChCjKFsnvpsBJ+z7Bmw/5uh7m3kgrf/sukKacK4E7zweVty6NDtqx/ZRGeEH/+WiXBn5+tA16
fIp/E3dHWijoZAUqMxXzxN7POhuLUNGHrmW2O0irqEyksQWTlWWwIX8KSXYOcOBbcOqLnkPu53Qb
a7sEY4NxqbHTqPFaM1v7DWIqjmnSPp88YZHT0/XYT5dvpVISCG6EeCv7koPpYuAcihdHrr5fQIZr
6PLRqqo6SQsSGMqJ5lOaMefIV0FLqqQ7dNMNP07TUtsGaKh4nOr2yu2yLHU22Fd3H8HS4biR7bLh
DPH9w+xRslPjbroA/f/R/Pu7m2S1XCfGEY89t8W2WEX0uo/Uj6/E3HjqeOCK2Kw7IX3AqodMldjU
tE74f0kJDbz3adSUBBbJLCB8v4O+gfjKdMojIgAcHyW411SlZD2f7wYI9jXvyQLg813iM+yYAxsx
NsSfzAoW+unUYpxsoRFW59ZS4czEjBo5coBigsIucqUvMSWdgglBPESAomIhCOajQF7gQrTC7Zyf
xxRaRZmJ3gl7Ea1zedQ8JD1a2xN3u4E5MCBBXCEt9ZapLOBq2MuDuH8+RZDHmx3ifMqoE+srcfAz
nUJwnNEYnyDi2aND9IW1WmrJghW/Yw0IuHC4jjn/jNImEL4tQ7BBOuyamcujWB86GrypO9MeKz8o
Z+xhCqvY8kPhnZM38tOL0XOO02LP4q/D1eWtxw2AmwdByPmCv5+gAINs/xnyWZUmKUSPnsWuVX3R
EnI0VcF7r/YbfBxYD1u+i/hZtqPPu0ImRQkXD5BAYOLdIVoaB/9OeQmkh+DBmxp2PoVhcAWTN7Cg
nHKw1GKt76pmQ/8od/w6wgNkUdu49CfZuSQG3/kPHh+tdYfxAIODE/SK/Au3St0uqDc+Ab9khis/
t6VRXsxdi21rQMLEPfaUmxBLybz/izi3TOjQDgLV5vu3UxPbhUJOu1/i9leU88N+g2QMV83F5FC0
sroxWVPKUk3UyqiuIk+mA83Q8K6t527j5o6AucL5jaVeJVP7d7Sw6IfQ0gCTxY+xQu+H7vFu8Q2q
weoC5vImP6KH+c72AVw8FJuyk1qIHmEciHyLtwwgTHHFr9ll8zJOc7zlA8XmLHuWvhP6ATJDI4b2
CpBEbxYIkleZQX9WoNw3AIuc7TVgdltexDBvX/m4klyKdMv2JYxDajlFq6n3SsrW8kiTXWK8+Ntd
U6EC3am8okaFR3c93MssY98AqjVSC3fLbKrH/OE9zj3HnswzfHbE4ldrJ57rAk50s4Ip3RrssGEj
ttVAieos0vWPBG848PhZsEyqX/HTZ5xJ2fY82/JI0wdn+30SDotatnutTD8HOy3lxqqDI4ixasEb
S1UinKJzTXnuZHHrdu91QXn7Vq606nNxEsrKBbC77didAznNpxMrVw67QwiJvjkCTg27vMgHQKvd
R4IYr/64VvEWHU4aVaajjQX8uHO50M9bKac4YCQlk1ktvQXwBAmYdGbtnIDjLInZNOItYFD9POFA
bAN8+eO/Hl0iLai37XghqUhAQbiJyuJHVjMfVLbmUS7K6Rr9AS9xC3PDCf/26eL9u6FOPiiw4PsG
iHSVD9F8AJzC6TAcym/Nrn4z6b1Jo7e6TfDfbOxr9g4vz7MRK4XdXar+2XbU67nZ5rkERZWcUboO
vpXEB4GzmD9/lbX2k2xgWak56RdqJQ7LzlseIdKbQQig7UGhBVXpkks8AonGPzycrH3RLOX9B1AQ
id9ZVOS7FlzWbxxNNzNrHBJyPVm/eSipWIxRrF25l7OpIp5P1X2aCmoPasNeT0HwgQEnWlKLSTbX
sIMDLX+9pYp++3BubYcKmTevbbUaqV5rUQIsOoUpX+uKotPBt42ZPvwIkrUifWoeOVsrB/jaC00s
Ww78Jv/Lz2I2Xeq5QCLLQy8Omzj2k3Td8D0pIGMpmOY2NcefuyMjQlvACN11aiFprPFh7Sy0JTR2
skcQJkI9J0u+unYtPTkQpQZez7q5cIXjechkV2Z7e2MQ7uC16fDcTri7GtkeXkYz/Q4eBmJ0iK9I
cvaa0c39NVY9tJDuHAUKlzxUV7lVbYG2th2Ztc5rNXWLJah38nmgVJmviBIK96nueVGwwAJv/4FI
dL5ArbDHWYK7gGZnypSke5KrCtcpr8vpyxsiBU7gwvxMWUqjPIQnWN6lrHWARB0rii6S+YZ723ct
Y6AG/iPA3qgHvXtX+5qgyD0Q9FYUepFYWuA6CFlHNsQPo9ZRvAc7BRP9Zg0s676zzOd+WJ9kc5cd
JIP8OZCcDg4+SvXxBZ/j/LjUca7GnISmOYrYEhu7G0kEB5hUqwKTTXffPGECs/sW8idVuQBEwprj
5XKZxhhHzC4R+2fR36QV7i7VYwsI1M2MDSG34+Tdm4gG1bbvth/kJwz50qhjlQae0hmRWNtV+9Tj
OMGhIWvXIdOB48Xf35WEo+fK2uMhyc3D4oGCgGxjaic91MWQsxUvtJfcdpetj9OOE4BzBfD6ehaX
s5tOdNo0d7Ezkg99uzMqx1liuIekQIey9AywXndRsel5N8TAaU2rZtzfdJ5hfHpu7iMBV59l1joz
NVHokWjxFXASdXA2RF34ECdsGZKcrlgtoUH8B1bNhr2sT6D5pNqYTJL4bI91pXNakrZQruahdzKx
vSAQ5ipG0oEGOL99a11Y/NbyToOVBviEEJQGgQgZvbAm3XIdLwUPLGFXUqHML/h1KPGFhwVgr9X5
zV2eFHVvMeYYW69o6NdUApiFI1o2XMawAxDESRgdc13tX2Hbc0FSWFNO3EWEBwuD5La5pT16G4X5
1e+cDBwzDnjZjJkJemQsupU8+GnzR6EmEfW/cQz51n0hvtm2sRnMpcveuIDEm9PqPOuTc4ddYgZJ
tOSWdxSgM4/UlGbE0uZoSLgpXZ5CbxJXUghI+AgTR5ZKenvU/3oW5HVNqhGqzJ8JZnC5jT3AOhMF
rfHNCRTOD/GwQJvz4l/rH6BA5d/+8BfpHufHmMDxnb5kWfLhlA52WIqOCtPEOUyFOIhnAJ8IJPdS
jhcFiMSuNleEKgiIVjs4THW+Pw2QSiBG2HymWC4tGEB8XHJhkAxvV/1YTXvG0QMYYCWR08b5yMpn
GkjvU3nHWHjSZThV8v8GM5Iy2waVHwMo85tL8TD/UvPpVVuvywHDr7mHS31KZX6ngOkdKpK28zjV
8QYJ1GaOhSDwO120SsNvAu5E+Bt6opfq0Sw9UTb1LYMkB2/pHHl1LzojPg915KjHCwvVGbBQJV8u
hN/eCEvFarJYmgEpu02su1iGdPDGpEXGqI0E1/77xrAD1NNo5WUhJ4TgWrP1wktbD6O+rsmIJEwj
Cl4NdLihEPfz8I6BDaEzkl1M7UBsCyTOALVHF30v4zT2beGCCTtURHmzoUJGicjPo8Abbv7/cRXp
DD04YuOBAPrwAkU14oY+0CiSd8eDtyqcetcKjNYEBca54GdYjzcFMXvxHHaUtuL642ayjgxDk8vR
EJlnHLcBYuU7U0mv/iK8VWXlAC60FMU5yl0iLkI1MSzViFyewH2JsyzaKYD7/vrV/oLpGmjjTFWL
B4YWf1dla6Xi8ZdsNgogXrz3GPf89Tms4XxUw49GdWnl1Ihfvgn3Ftv3nd2Nvw96wuyllMcjVVAg
YfVP53jghX0GoLLtrbyxxi0LvjPHQhFJNB1sbFc/nmSMCXt4y6621Eko+0nBYvzW97JfdL5rTeoM
mSdimimw0P8W9AsxEz8xtYhqZK/2InDZvcHs+soaFbz1jZLvyIpN8pyKUDAXqkw8T1luhi2Hkqry
48X/Omgv30/7nRW/raQjeuUpIhXhui2o/zRPXDMIkna374+5vvZZTNu+u6QvgISjBLZTHqP8miZj
lIYOuX0DTSAwd8Bd77chJMBSVSZWA6Rx0nUev70jzcrQu9DxWzZvHWt3m4VBgVqzTQH4UfJa3mgV
DP9Wk/Fmi5u4g73KPuLkpa7yiikvWSJ841oXb0AP94lVvcY+3RvUV8Xb0g/lml++ruqE0XjHGq5n
uqTVLLCq/mPtOQxI64dPKmXZIn0LnP1dnKVwkb1lTib+beJlYn0Y9w++DvVErrt3bD0OfrKypt8r
nuadv26hOcSy277NXboTgxErjkm6w81XqU1JILqIxdfUaGdjWoVxeooppT+KEli0h/q8T5D12cqM
ShLduZu/h5yvvakhdYB/EsmUATH33ivylzd39vZOXrTcGEktmFjjQM4UTt6Myf0Jb7I4tdKoffQ/
pVFiyf4N+dk7snv7fgz2f4mllUIR7/+NlOAr/YKDG8k0oGlzG1nQUgS63p5MNzRnYjMrmOm0pHr6
6ScZ1lkG8fxDaSdP7PtPpdhoHEOqCCZrU7N1oaQOeKDNWrKL1BgqUTsdTltMFXYOypkPbuk79n/h
E8q9bsgyzOnxPB9biBMlyHvvttf4FUWjEIcaxWSFJvi1cM5Q13v4oUK7EVMWqKSikQU7jEtykKQL
1dJWd0dVS7K8wkF9F0srEQGKi3vlkjI0Vch968gcbJL0WiXEGJy4SqX3QBUbkG5OUP7vSTKXz4DT
Rz4KZ30+Hx2eLJ9nMf9TPkKfJGTLFyeO8fMo1LRfhMf7NUDmIwWaewCHuGPQDgNe0wjRgW7+Ya8u
1/GOao0Y+DrykNZl9XQBFa676xwO+L2ljMN4zltnfXHDnoy66tgeF08oe9SfvMvHKzLzOvhmNJ27
PVbOImZjPRoVBSXqbicDQKqllSIYMXaRWdXsy/gpkq+l5iRq4LJpR12t8Ma3j3yoTvPSKBADJabk
xrpq4sNy4ao57b9t6kcB8XkgY4odtisJ7O7wVLfrMR7NJVn8zcB0sRNMlw0QvixUojOEuhO3HA20
biSsLgXPNE+B+O+QgDvJor8OW2RLEWi4JsgBxGq6pLaQbKC0n5tyS8ik0uKAoeduJ24PTdCuWENK
1zq5aIrHh6/+aXjJH2qoeml56tDiAYUzqiqwIKlOeFrsFaX7QZqjM5Rqz6da+0G5U51GSD90RhNm
xyekCm9w8HJ9VTpi6J5qUjbp2RL7+/NdYtEwO4CDIvAbBk1MyoKpOoKAEiK3/peU20kvWIWGCZFV
RZraefDgNllP54xlI8aur9pBgOq7g1yVyZbFUylwT+Mu32w61j3dfw3DaSnFeVVquRDlBKQkC8er
zG1Ga/aNOh+g0dnboEu3nx55mskY+o6vaqPAXIhenbiwIEcRbITMZhTH4/3Im5CjnCb6xTgRNbKO
gMCiWvotUz+nUPY7YNgZJvfzw+YIuT+VqMCbZhzvfqHFDNph/YbEnA7e7B9LibL4dVp9gim8mFJn
oAj5jEli4cFO2u/ncjb4OMojVur/GPwviY0i+0kUWbb99nlxulMscq8KjISJcfg13+/CSj1VK5gX
skNWh1lLYFEnuuMw2XYBBztBJzk290I7oFobuR4sBk6if3QmyWhsXMsXICKNB8YkJa7rHBoauxgK
zURR2M8Q4mHb8Fz8IAokdGzYH6jKuyyJl49FjGCWHi35QJLE3CNNNpKq3mVXw+fly83oRwqPEcCt
JF1ni8rTqaDDEG8NM3fSK45r6+NIhozDDtn1NC/TtsFYF6UK60J9TVWL8uDjSxKwAiRx8HEF7pIR
nwCuFouOBnI0j2WqwMOmNGYYm33UPdY33i3elpN21ZGJAn/D2lrCtanx6joE5wKKLHBY8BU3B+4V
WpKHeefpksaX+OVXQhGjWbKIauB+9BYjKD3bF9An8R/bJV19OUZcifB4i8Sqi0a67hm1zuH/4Wrx
adkRF2geKHMGKmSko12g48Asti8LWGn0zl4kVWnxt+q7lXEtZNeKxG0CVI4WGN5vmdbBBLdKAbUO
5zz7s+pR9ro0l72UJuY5LSDJclm49Sn43dr4QB49oQtkQ5ARVCQRQ7ykQk91JRP8NnLIVps6xkam
UqvD3rq3ku3HvAdA0h0uGapks+jpd/fW7V1T+ItyVlq5JuD8yv+71hvctSkbe8jukRIWjrlaKbw9
by6KHNP339q1KUAQOBcFd72RSL+OYOWGEqfAT6nH8IY7AUpeMLaGSaDocUHwpIcUtkXiePgL765R
93kdiTs05M3FkPjp2IDJxl1iqLOophyB3zXbfU2F3pP82Hkw7wygfdx8JPwfu5prb9IokzL139te
ZFWgcuZE/WnXv+/j0jCU5AmUNahrZTzSeJmu9VUjFhGBD7HXIAF+Mynr4mE8Nsk9scJdVHLEeH/0
sdtxvGeYPOhU5Jgxua2s2q+11PIlevRY950CUAVkHC/Tm4xTZIq1/J9aE6t2ykDOxaqtMptwJdWH
gGPBFwnVnVR4oI2kIEbIfqDlahe28rV0L12zmW61I9l92+6Asm98Ck00waGBctOFWnT0UPVWcKvc
w9IvRr5hLZkJ0l3CnBHKmpTJMCzfW5NVGliA5UBbZE2l49HI0tydiFIm1fTbW4yWoaDOMjfJeG6O
zdwELsDPdTeGwz6B7Rzu+QZ5CQ8zNDrMWO6Fja0IxFs6b5Be5LsKdEgd2GJeLh2yF3VWbyZ/m5o7
oSLOs59AiFTJx0YpWJ+tuvpq7zngGugkBwXaKIYiMyqZ5xyTHcWlpklLycEP5boCff+tCPUuOSfd
mfvTSu0VT8eEgEw3532C6eGa2IgFLGkUa/q05BR7IMrGIMj/ZbvcdmpJow/s1FldX9kky/M5khoj
frCAO3Bxw1F3evenTDiMfIdWywA9qphq7eWdBMx+KQeyUN//Dz5AQJODrEYhbKAfVGWaYohvEHe6
tfLd13dCAf/ZoTwllTmgVJ3PU3U2hZgQmFXVlFfVaDcfmL6eOAgMHjs0gtrzkcQIzeMQRy0AoNT0
GOl5uL3eqNjs8ZVTx2pQWkW2iNLqFyTqytpKXa+xXIU/TgtTLu77XSzCSpfDgJcWM2NvGhRRuswR
MrPxGlPK6yqulsOqSo4ddzzno3TstKNIkScwkRdsMF3fUHiSJAmIa2km2JL+N+C6+jjserR1NCoh
qx0xhBXJSNVK3yStzO7tgr5C89QWhxYHf3bZNtebbdoVK+rA2wZijvaqgosxAuTvN/YTa7FsiZlw
Vmz92n01PkYGmtFNqDPKRlv+eiR8fhNxdDL8psA+RWl+Vmh7SPDyq03lvSIH61V1pOYFNtYqmF36
LNAaIdxPGE4NMMG6xwvPr/ha3TDp48LneIBwXIaVQGJ8nF5WKwnpBWtFCTd47G8q9DZMDRxc7F20
a0p2FGrypCzHXQdeS7YnAIOMHppLeApJ3lOQb/NtcaA2HlHZ4oBegnXQnhSN65lb8Zg+A8LGihAG
cJJzrUUy4DZVFaDKumFCjSvuSOMJbwAq6PHAhDfg5BOsvS4JFmkIq8seFc8P5/wP3ik2aHc1BCFl
Wc6I0YEE2UA01+xLqWDeZ1VtNJPgJpdGlzqCSbc5Lof2mdyDR8+lylm3p24G30pIj5Tmc6dIXO5i
rSh2fIKiRpTegGDyD6auk5+9/ag2r8ah5upncJsECFk8gzx0s7U1iHbKSb1hSoQ9kJOePJqyDDSi
8JGKRBM7MJE9FFBvr/YOY89DBIv1IJk1wsyucQzwLYxmgFUcOlHJtBkFIZ8IIegv15n6I6AZ+L9W
0BmUF5kyeBxbu8keITCNhqB9hQG/xWDi2Wyi3DoAniGEr1ZySIqtUzOpLWejYMoh4gJUDvo5LU/a
2iNHSxLXCaKxmSsL+T8enFKM3QHxd1HCla0bw5oFGrO2yrOXvRLOJGbwnXBFxGJ7Srd6Y/6ptz6f
Ysy9KoHFbWIU9PwYv+zQPG7/mmJ4MpDMRLAhaOwmJOPg6C3VJzD/GsYykPP9USCH/MFw6hDKQ72F
hDay4nZ9/jmbaUsP6ygkE+SWuHqz7Gz1AGLZt+37ukOfhVKBml79NafAbw7evEprd7kOCbsrlNkL
CkXVv9ZRpG10X0uUrBD5fxFz0CXdzPKAO0MNN+rixClir9Ap33kEATOvDjmUTlwbO7ZQ05fFtGyM
9AUFrJUJXqLjzARjBjfholgsV7N/6oEdgP0WLB4kUm2kJcUXNoOu4jjyCQJMpFQLzuuIu/AD1Txg
9Gq2D+6dB2NxdWL6IS86Mouwpy4EVhvSTrWMMf1Tz9G6ra6xM0pyU/ScvKJOAGUVHcNrCUKrqbGO
mZyuvqmrTH/4bd58l10RE5RKfdEnCLzJVwKn9Va+1ILUyOxxbXN4smBDzqDSL/wujgbX+FbNEyJv
tj+E2y8Zy4JmKg0IPsMX9r4K36U6oCrrSK/CR/qMAkyngRTo+DsKzWFsQlv36X1wklshQUH8nFaS
WrmGHq+3uv3I0bHV1OA96HYf81dgnYF6tt0DZg37wjkwQLkQoKSksadWaiu83ukpWUGPxL+NiuEN
wWF7ruS2zBqTeVhqF+T+N9ncI3LAEFjv0O2K2qvnSvfg98jEmnc7fHxbX/DhTqTqdi3pJJQz5P3l
DOjb5J9YiYzO0HzFjdyKZOtpJcb6hNc0LG50EQHZeWXvbGhsTCfHStM2RIZuZvctCKdH/ZPj1AgO
6xJu+aqf6hKY/A7RS2UtcxkPRAbF3IPNOY/+OTeJS0LJCUF4Vkv0or9TRADCqXN4Pur5kT/AOLFR
zLlzlhrG/QTjdS3gOLNPKmwMh7KRcCnR21Bv4IykBtXcqax0J+3nhiPALn9tLg5mhvbR6lIHBNw3
8qbZqH+/zlN37ZCNCzqWrDzeUI1lZEifz22mmgK1LJxgcdBn+8l2xJ3j24570ii7PMETmhbJiZtF
4jwhnJ61EgxQtb3x+bP2qoiUz+8yKMUj9knd8ggRFlUKC4i3yAPdEpPZwqzDa7V3BIjkBMha0y2L
AtBhd+WSdZGEWuHbAz5/0637NHcuvnx+yQjlolsmpBIJL3CT8sUbFa1dVuzjZN5wSxn3xHQsFyVV
wjiYHnr0RxgfnYz2i+ADggeymRZD2RMTpgSzN4h8y0J0zUzktC2U108sSrdSJ4KMTe3V2nzme3Hy
/tGwUiWUo3NxpUMGKS3oaEMuHLDlIMwtvFEFv3XT1LW0NWSvdO8MVwK9NPjiWkpJb0z7PNnYUR1/
Eo9OpS/Ro0IA04aAVaZFAGcvXO7Vc3FVhwOgSrxyMmmcujlSYXAqw7Zyw8iUQediIKb8XJqU7qqB
fe5/wMIGR2c18IgdLV5VdYbdL3xlOGTNUagL87JSwGLbgR4sSyrfJPP2uNAtC+vw2kySnUZwvza+
NSkRDnGB1t1AQ8o5X8dnYDumvK4NbS/kF+ljn2kGFdb3zFbpM9G/tdhMPTttumnvxcvp9hRGIjB/
hi1tY96l2yisn/wrlgLHY3paGS9IHz9kqYC2wCQAs1EN/aMfNV/gpul1OqVf70pBxjIvTML81KTc
KV8vI0ZMePV0ZCzwhAcA3mbkvhOei4XGcNHcrclf4kIOFPosQDsaTLpGyMiBA8lYqwc8KOp7VQk4
NXhh28VmyFJebO/2/cqU6LiZEDffgF/hPP6Inf/2NnA0puIGhb4oihyJTwddg8ikD+dSszzNjAlP
e98dF1OQW40i9Q+Dq24rj2NPXDYD5v0/YbQ8U7cIP+gY0xSI8toUy4mUUUmSofn/wkZcuPF5Cy+l
JlPF7qGTHeoOCQiMXClKTkXPIjChlsCs6OIlv/7LFH+PzZLNmgFsetrxjcfXupDv4m9TlStCRqlq
fNysm51AQoV0pWP1yo4X+Gk2vEiUQAS3Btdvqucf2m4SmyW8XaCqbMj84ctIv4hjTaNvg7doXw08
qDGBRe81K2tvIzrYpue0JMNXrW7T21QTYXL+Ff+8RYyFGEtUt/LvSuoqmIzR2B2iW86nrUnh4xep
UPxTIb8ALKLef04RMy2dOLohuO9IoxKxvosJjw7GceLWfTQxLxxiu7nQUpxQV4zmcB1/wUwk8a8m
jCSmVKMvdL6A2WAda7SF56Ow3ioL0gEkN55RNkT6z2lKzvGE48sH3JQsd3Grl7+jFYSAJroVKmXe
OZEIuY15z4aujk+9B8qa2TS0FcxIpvC14MqbT2yWmkH4LsSHxbmxk1iH25S0pncrkPmA76qRBjmf
Um8fimcY8zTU35dN+2EezO+KMiICl4GJyXGIBTODDRCvNIGkLH93SpPFaLkhLHlHKZUm2FDJQmTK
vHQLLOtWljOtSKbRxOVVgxgHWLC9oP0mG2oVWA4GnOe83P3PlR/H+YcnD73Mydof/sXkJIwpXB2h
yJF2U0F0zeUb4s7BKGbnqRjqIcb0LFLxBCcmXnkYs66VLeCl3w6TpBfVD4hxtai8LUpVntw2k3sY
rg437pdn6n3pYKolIyOTnUI5RzRm1DKPjyFqwN/mi5Fpq240fohQLCD9wdPUPr4dAtyBkqQAx2Zd
Inynsk/ohnzvoVUtjVeqTw80iQqyfikWgREUUmeLcIUsTvreQ0X6iflshAIAS+OdfqW34u59ROxj
RA0cJj1I99IEfU6tzZ7vtkh3sDI/poL6rPvk4AbNr4FtBwAQLrzOFl/+vWvOezIgxETdkp1KCIlO
gsIDW3K2N2R2K6ZQYJZVCuNg2XKeyZxwUHEJaEMRskMBtaiVu7hEPYxwxMsGLS987pajK2TC34JC
GKiM9+kqM8kO0Oy4QcCvo4xJL+nIBBfzWjS4Iky2lbkLtIfPPJatH6levBfTnzV1UOkyEk01tT+N
6haKopK3O/GJlXmzeXO3FoMiLaQ56yjdfKGR49wEmJf+fclIPKe1PK//dcvFO6ysZIgiGj5TvJme
yjZD96/7Q/VpBMW9Io+opkcTymZGYMqyYHRugVWUPcE+CTA7t/ahCZEt+XtunSoc3bazC1kKl0ke
34NELR7MVZf1K1OSv0EF71TdeWfXFoxVgV6xIXCDYavCkiHZdS2p7V/lty1Qn+/KwcDwX4DGylbl
0ZR8zQDpqpHKZsTPsoQgBqYuZS7KHl/x4ZS1Uy+z9qXe7VmiJhympdF+cZFFh/ihWpSPmzuSaTGE
9cHAns2GGXgct/Rvec/Wp/mZQAMtb6FrWyIw0Z4UAgaBNQAjg1xsim7QGNw/cJVaKXjNB2stIUbA
gFxc5ve6mSutPgXjfrXeekt2TLhqdER40u1bOCNkafqqJRoSDRmJPCT1kO40AOCjJQV545vS3VaT
QdB5/rYYlga3zSf2EgT+VA5z56ndnOY9V73ShP5c1++E3F047SII7uD30EjS2/hOhpA2jsmMmHCU
FpLxXFr/CNojwHKY2eucXJZy6qjP8hupnxdCJHnAxItxRFmAlQ1R241Ly4WmLHB0RwuLbGHOO6LQ
/Zt56bEQdQ64aSTySf6hkl0VOPXT8dVHthE4wb4tBk1rOa2KMNBb101SQDRjhxx9U2hnkkpgdO9g
FeixLMbZKpGbFdjqsg/qZINs0RuTU6obmEzrVin5eD9urqkiwqhIwGgCAskkj+ZjnzcIjZuo8BE2
TPH7/sMYaBJNdbfipKX5+L0A6YANr4PqNQHwiEgH0tCr9aWU5DKAuLe1U311Agg8KfIjEptTh2ij
cBcRC6NBwBG78JcrGFDECquSqJP5PgU5aldpO//L+wBywJo1FK4gUiutYgkuVGfirjk0vfvDfvs4
0hHN9BUMsdmE39jW+NaS7ZCDqH/q6xSetgBbjlhL0KklEtbeOH9or68jp9XbUK61iwRJBUgc0G9g
mrRP1ieJSEpqjkLlDasJ0ryUZZpUGVU7lPbY13AsoeYdo+FDPzm42b3cU5vSFACLMGD6pjYoVivx
TCMi22irEaJCNTq7QVy7gVG2iim9ZViMpifT37voOs+/1DaV8PijYX0lR57Pq2zZQbxyOWKtvJv1
EyYIyONIzeg3TeqBGB741t2CEHO6m9DMcNw4lsAgSb09XKXamW+MHy9KM+bI8kmssjUpRbbFMRkc
y8PoDuy12Q9FZeuHoDuxMSukE2PDF4mniEGb4kkjWvsU7VSAlnkFqBxkRCOiU2+Ap6cV4rv8uCjw
xZQ/5xYWeW+KYG4jnLqWAbGfevi2YfEUHUWxm8MeLeU5ln2NGtjjk+kzxL2Mkog3fi3dxCJDLHio
0+Lo8aLlKAsrNY5LdLHpoCsScmhkEkzMrI2bqGgBeJB2Cg23f9nB+c7AcoyqevZw7vYDadtglV4P
IUgUlh42pE1xJkl7kf1dMFvwLC4/q9oK/R7PXQYOHl80FH/bvfuXBq72dyRfQNaF6mEB0fRUY1jB
nVpAKLZ+zS3w9aQGAhV81lCIUsStPiW6KAdiALjpEWiZjpR56VPOxrEENnNfPXyPLDXVg3Nn0e6P
QDZCLjCsxupcq06icpni8CNfXFBf8TgCQ+3x9pav5t1XTs5EKTXrXEf5tPKzlX+6AaQyVsRSHSZQ
PEeSaEE8TOaVaZyHsb/R/4F1jw+j5cWuQxAXi5valu7Tp6b8vPOjRZu/oNp7A+MU+vu9MVTKMAYV
009f2GkcNCtMmNcD+NU722ubffiA8hnbUKUBSLIrt50lytaH7T3wuRROtMkY2S0g8NhUBxvQw1BC
ACdSfFQ2piIfyEzpB6ai053u6WhURB6h1dkE09LO77wxPavKu4I8IhFLNPVoX2/GdrsRZaHyROfF
bfl2E2vDLIsbboqpUU4qCFvEhV3LLiUHlF3Gw3ZsJwkA/w3k+ytJnsPopqVoIOwoBdlYp68JEwbs
H/XhYVGD93/PArNlYhtyRzxwFGINmSWoyVbUSQiQvvpfvFvwXzBKU+PCTKVwALya3q2mDfX+iM+L
lX1jp+ylcA92pSuFby64kA41C9tydOtTrhnUrznthHwNxR59g0Mb3Ras4juStz/mAA+akU1ZtCyv
lTOIgpHo787spQrZvJmkTBS8ZwUcAYWpznTYAnlZtkS3wc6PZuiVFt1vSqSGL704FxlcJnUVUQTf
c4lqo75AkQUzxs6OmeYPLSICx8I9wjC17B9NcWPExUs1O6SzTO6gSNf+Zno7SYdEPmC1RKmZulXq
7doCoztlMLav0nk7n5042hhlnn1VAHj3K0qT25uT3RVlbFSWYSbHtuqHJIdfjQnQGS95fI3oAVYL
ZU21SMhaOhyMPQ3S44rHxjwSinrKdHn+QZS7tBEJBOlSjQ5xNkpFD4ERrlXHuaTkKYsfql2ICaaC
9zeRREr9Wqft8mSfx9l0aj43tnCtoWO9lpauacz+/DcvNY+zY8XUd7aJs5YKEKB5EIBDBmO1tT9K
bj7x75OvdHJcYYZAm8b8/ZSr8kKBliVXrxZ6UbUbqPhDF/jt3raHJfF8kGHLcVvXEGhgNHa81IBL
mgXu6YVIsSCCxXgAox8AkRJqfqyWcmm82sPJ1voF5W9ZVM4pu5qSTHypKKtNGzSfZ4XBwuLJW4b9
tXg8dzDURWEcaI2iNDFc+GHzL9dAc+dwzjI6i2K84lTOt31YwSIXdvm6mzrPehqE9wSeJNldb4Lj
4jsR6IGEXAlh5nzwxBtDdEqfnBvqvRqG4KZCmKcrYuADmsg/KqHzkgD4gn8dWikQoeBFoejyFFwB
HNSf+ZDVxWRzfdvN4aoRN6fp+3PVl3BOJ8bM+4juN+ZSc9Mv6KNC1R/CfQLQePyFCj46mH1TjaX0
pLESaUY7+PbZFdn1lLRfrmPHqlttJbxnfv+4wCQbY4/NEcnPVp8jqPTFAG9+p4S8noSxmiYvkBFq
UnRqN0O/TK+Oj7Xbz+Kiguk6IL8682bxa1atWjpjQww2SKEl/o9kpNEX3iiLHxk+169s2+2j2xvY
VEyGiPbxsjfDN8uvmQQHG8nyM905Otls2+zdeq0AZowIOxTre6sYm2i8cGvS4m5uwLFAsapZCCnv
S8SmbYQRB6CIsqU86I7UMD81jO7ai7nKlDU5LXqdve8r97SPQm+63IqQyu/ZXbtcIJ6D/3UDQ14f
eBDHqoYaEVB8iglUiDFgL3BX9sHxygSxAbnPF3ieFsIGK30E5M+oMp1sayAlhy8xePgOleC3lZep
DzCpVwdSbQSYvLjYpEYAReWt5I0kCAs+0UaOg6CNjiT7lhITnE5+LwNfCIr9KunP1xulebZs6oW6
4hsgEfhoZ1BaY6zwT4oes7EKd+bWu7MF54uPcaw0dcvgh1c9OrbIiK5Eb7gx4P+vvsUKi7RFDOzE
zP8R5McGvNDvjS/0yXp7JKvL2P4oshg2Ed8mGhjlG/2iffdi538+alzUOiMDuzVezeKeY+w5/pK1
GdHXhzENJFjPQU7/1COf0/Vq6jpZpye9crZm5a8WtqQYg+2vaQqQym4F7eneT6m4syoEdY1/DKGM
AMMoDgHH7xg+SnHIJ/6osyY7gnrgGy4j2QpMN1UWZQd7loiITZR1kNqEs09pK+dl0WwWCqdBIM7j
9O/JDtDnEKkQ6MEt5s4/P+pHDqOUWm4LXohunph53qoFAj9hvOHwP3aRadBM46XGuG88yxB1LDli
yvZvocskm6+muE2Bqi9p0PdJrUnWuHFpZZPwjfW9WG6kidtvchcUbhkHGUkZD9PzqZ9Q3OYigoJD
2GunGktL3zyOjFiGb1hSLG89pAr+SJtkwGmhgxdJ/w8+rqhM2q6bWNRkDVOZKtXYAtf1N7JF00vf
2BzU5kwXh2DiGg0+DoC0wvjUiJRBrSSID9a9lw94rCw5KBtBv7rgPviIZlpo37/tWfeK/oQYRkE5
CZe9WtpWFaPqt1VhEZFEIOiuwxJbvniV6mzhq/JLdAASpcSQkq2UjGS2d/lMOpry/O6F0b72Q4do
Z5lTtXOTQnwFfrwON5/EfniPUM/I3BpaZGR9AHl/2Nmknd7EBurVFdZLhr56Tz2KnUsaoN8zLRiC
7gJmGEQBsdI7DB34pEJxu8W1Ul/TbTO5XbtJLa2RT7XKtugoHho5prSeF0qxXoMMbDZMqvhlB12k
OETzxfi6rL+z20+0wbBb6Eu8mYkQxFvU3CD7C7XJtQkeKH1NglmqQPZVFqnY2XB6cAkhOMTqIpHI
HAVfMY0ou/Czi/1cN0GeUFlxONJGfRXeclWweOAnEHVyqq3ufjmrB6+QNFypG9Q6OmquGi3QiPSi
AIghxD1yQkOVZDlf/CzeSqRGVBcnIfmAqhVt5LAI+zOyK+oMxrgBCjTu8VNKTuaEu/BGloXo8maT
Az2cPKbD4gf37HB9thkhDybo0vWLcDQZETQZ26LShPx4ixt8PeZQ//KPpS3yT23KWbFVJC06LiZZ
NVxji8KHx+D4zL/+6cIQdHK/hdGWwncD6PKDEZvHwHhE0agC/553eqL+dYptio/1p8VqpCadmEda
RfPwS6RD1MgGYx6rqd99+LuKn9j9QDlP5L8IBlGr6hvNIoF6RFk1jaN7URQDIpf+RD6ny4UTx/o9
MiNk5XjGIf4H+Q/ceGgMKezbCvQR8alEFZjhK4NXKAhnwC/d6iUXBNIqIJZpcHO5fqs9DM0QtOD7
byk3mdQcws3L2hsUsBZQuwXQ2RfbbAmJXlEUBkptMAZWv6yIYScYdsFufEAnVDcrjnQW6uB+L4aq
36qN+buskBnHF4PB/VdQBNNBSWjFbkcx0x6jTpnx/cv5YN00d7EYRLq48tnCa0dchE7eyi3tE/jA
K1EnQlA35+j6/JlyKs424ElQtoYs5Hdl5RkRtJhaEgMaVw9adHCZfvaDYl15k7W2/vC9Nw8pKd2p
cWhO4b4wRXKiIcPBMgHjvKnK4MRtf63uFsx4fssks24EULVZilCFM3xnnQtM3falsJoGYa6Ddafj
qu+C8i2/YOyKbdoYJywFgRwWZ8/QiiwcYNijr3ILbScD03BQL7U13xkAZyeFf9mUflFmi7QlCk21
TPLSly71o8X1b1T0VlXiJ7MBJfN+1Pm15CSVpcIJ9cSv6wxXeHLUW5Gc82UAoXEQaYjtVC+UYsIu
UakEtIQv1fJDaDtk3He0+0gOcC3vtphc4iMNDBNgeg8QEYhJmQhiTvoO8rDP+xG72h6F7AViJ16l
ScKNLMm+6dhvTrBee1uDporNBkGC04ABA2L1UiR6vo6bBCj02zRXtrD4uQeMTEB81qD945HrwCLB
I8Z+FzYXApqMzdFnNGQ90GCWR87ZM/Y07i5prrVE0BJ2q/hXj0vW/NGd4QgocHa8FC37NWwUoYt3
tcLIJoQcvstowXBlnOhLVUdkg/PN3uWMLzlyREMIULTlL5KvXydq8Z1YOLX3x+YeTV5ylWP7WVZ8
R0EPbEWGcILVP/Q6N6WK/mSjYnb28scIDUdB7cBjrAUxHPT4UFOwS9kyDyhp7PrJCaBvjzXWChxY
Juo37FqMFcfG3xwlQUMiefgVZsHn33xY5m9NfJM5dJ3k1sdIYNi+QsZZ6FNWIe5Z2/TYdxx4K3DA
oVj4FODUojicrAE1/vs+VJ27L4XgUBeUCQc+FCz9Xs9Lr1gRdmyY88oF/KN6lctp69vkZJ5Cw2CA
0UnRmsSJXO4RejIMulOJMxvP3qmnM1KLwTDL6X/aqVB3d1x1ZJykzzmSR4MTv1Ze32agSEP2Eztv
MYumlY4RlQXs2QYnH/j1BJ4UrJl67Rl2DCQk7uGbw/21OBX3JuC7kcaA7hcNePkWJPR7Ggcj9b63
EigBE/e1RWZ91Q8qVD+gJgZU1ofiKlfuqXzyamynlGdzEcD0a3ldyJx5ski3i4TdxHgcD369IFRk
SKTXliMlBkIblYwbzAkRMR8qgvMUkW2l+FyVnJvr2sk6o0xKxe9XEq7wi7MhkRgEgv0swWYNJef0
m/cUbPRRM5Isu/4BLRvQFzHARLJ7DWwCD/4/+XiZZhwI+fYINzYNl7/5AxeIhq+/2DWFp2bW7sLD
9wtbo9Qiu3YPwj+K86H1g0Vu2iwtdZY6JgIEfX5ug1VvGXCeNjnKlkjvC+AfCQVugv+9b40/6YbS
SqBiCORPFJ9rFOgw3WHzYYJ/RGoh9UePRdZ5jF7AFryl+PnTI5uP+rV7D2gFft9UHmoBHlTfVCiC
yVdXHJtsyYZT20GPGtJr69kL/UQLo2TjcI+FbZqZ5/nl79qvb7JDURhYEB16q0upbYSwVPFNUk/N
7pyYNwEO8tcnhdy3onAWPEIDYiEGylx87dXaXXvJ4wZxwHfPP+fwgOcFEXCcNBkeo/7xIpFDfj+5
jVLc0OekEMdYj+P6eOZxCOfFEq7M6khvWD47ryBiz+3ZsiblxGGQzOMKgRguvlZWrVy2E06P/Ihg
Jw1och6UzfkAb8Z2v6kIsDpdzRsyoFRHapQaMo4H2GNdiSFUIRABTHAWCkwnGMv0EbafWb41IYdh
o6o6UF3t1jP3DS8elr4hH3dJdDpuCN1+BLO2YmGLKl704uBwLgLZRe6U5l8NIS+2lEAOx2SSD2XL
95kx9KvixQivBNeX1I9HRBYfAOGsLLiAPdcEfjAWaN43D0dGvcI8DJ1QLGS6hnTixfuvBb2yjm0V
qf5rQwk399A9SA47zsNkzvx+TtWLJM5Q18s5cGUPWVqU6B/UC+xa2P8FfXJfkgUnPFgbsf/BvrN9
Oqycd2FfMYsSArgMUR9Gtpnv4ZC3OkZMs2EyWEc5lUr6sApg2kefINJTCuREuhGPNsePFvh8fDLc
uLLHeiySrbYQ+Etp4FGXubZgUkANNc4VHvFIk4CVYHMFis20E1+wUPhUXic11sECAniloUKB/oAf
C0I2vcMPNb/6Rn/4BOzB62FRS7zkfUWcYGcjBqFsfxAB4x1SPGSABKua4KUzu2KjiyaExwN7pJHS
HaXwtaIKGmDgj9i7ECDTCfLrNG+rgOGbzUb757A9oMGHtUYqlV5TrZ4kZVT5zmvMWRPGknhro4G4
yNsZo+hPzce58nxmuRYXFb6638AtppOdeSRG0PAhqDCZTFG2wthO9hIR4jb41DjCD7lBPsO9+QuS
zEjlTpaAlli6v0wv+9W4JMkPmEhSNoIX9EMc8pPoAz4WAwisOYEm8pTbrnv7Bf9CWWoGFXY4NO1E
JLov9V139r5401R7X/8ItLF1Tiu96kKrG60M2p1riujbu4QPLikDKJISlf8U/JtPzfpa1OtAZkE3
2ySdzSN2L1FvtQp81FHnqCLn572sQkTSl7WxS0K8JPw02/2okMoLmVdvVoL50Pho3sF6Jm/DlGUW
G0g8/ojxS47ahO5d2iddgcVjIz4xXLjbfMpVFFSbIOQ+yPqMb4j/szYoi1g8E4sKHNk39JQm+tu9
InpQ57FJQGU3h+NMIgAyF2gSVMl5/S2u6DbYd0W1gZ2s6R7ivEbI3pD76zz2Jeys3mJA2kXV++G9
aJG56BChyhzcubmP4m+btxMtdNVTyQJFW8raks5XIeSnAdl7g9hnPGOCsKX+i974jhBZSVXb9Gd1
/e9K3srMX3JUuKf35r0/PA1dPWC0MqhRLS5NOY3Bezu87aa54MJz/e0lk7ffmqkJHaaee+Zwwknp
Lxq+sJdICwNivLeWRegrp0m04Rzd1DFjNuzJZu4iRm1cqc/V0zrGwOOx/brRoou7G4puaJlTV5/n
vaXEXj3EvgfnTg5UWttxl1fTjkZAvw0M2eWIRklJBjKWdZ3Kj3ZnNy3LHI7ALrd1+gGWV5txmRji
CRFfPPqfcSQrynI2oSUgPWfE5WJfbe985g2LLER0ocju7T8+RBws1Fo5Lvh1jg/IZVsEq+LzQ3zy
wJ4otDezpWnUiCMO/INKSvPHsU9LeBUyM6qLgx+orkOUEOBDYJywoxRU+eYtzh0mcD1aT9/iUO1B
YYMkLKa9+0xNVzSQsR5RQ5fLo6GplVduNqsNKqE+jSoiFQnCaOsbnG7t3rRVp8B3k5lP+jJiDzMw
y84wQZoBuIVF7FAkZUBKTDCNL4/9VgKcwFxR7jDqzmQInTo7aOI5UDnuH0awEmAj8aiX3ngxbQE7
VChmF9svqa2bzAIU05krKrlFjUcy3jZnfMYmB5YKtoLvui7CUvv3bK6sER3AvyylZKcjOlZIx8yv
L6sLPOB1N1MvkJWmEy2U0D1glPhyXJ+a/xdW5Ckw5XTy71F7m7PC5krb+ALmrkOOS1a7v/xLGLgP
uRaBXmitjGKQLdKUiMCJHQCREDsv8gXnKZSkMy+IUCpObaWP714CcwF4EIAB0aGuYyJI5jttl3Z/
3EZwxaDr1N1nF0tWnK64SqwErQvC7ob6WNs4FqiVsO+Ddh+N1zKyjUe7FWwtCTIKGrlvnpLVM1uT
5gD6LV/RWu5m/a+G9/jPjgAbuJuJBVvYwkLmYLophgzP/LXKSPdzfH9gQZ7wIpvY1Y+PR+CM0Xmx
lGG9IlQylc17EA7Zoq3d36za6F1qE8428EyQnuNk6UI0bJRtTaaIxNEQ0A5sYhPTXnrAUIX7yKQy
USMTwEZW9bPDFFXR7fxKZu6K0eulHc3LsYzuHtudKTbLnI34cI1rDuoFvdmGyNf7MIZTA8eZEwFJ
vkSdPuYDBjTCZamMR8ACcayqliYlgggiPjncaQqJyZn5sNZtSCWKDXGsENunH8D0xMEdDzJ/5co0
cL08r5lBdEh1AcEj4xFq75I9MiALmtHbNXOAc/Xmp9/AukVVYthuEWZroRdfUxCIKmnEWuLn+YgC
nQ7cI+npHk7EcY4XB2fOI0N6vod053h8CH8/cZc99Gbu/KTDoEUfIpGfrah/e9Bx0emRtN7QC6n0
FtIbFd5xpnxkjdpMeFV1y/IfKyZaDQkNtOQ4w11zTFAUPvRmRFhs/I8wH4r40MBWhm+0lYVYJz3O
8+s+thhSN74qSYLpGJfBduqYnWns76yIaHQLE8BO2pjQdU+aHnv2HyYYia123Zl1Ba6adyLHNiNR
aktAUdalX+NFVhTCDLvzAanrxuA7yQrmY7ZT6i+V2QUh1N1t1RrFsbylwmgTRb4076G6JpgH60qu
LZGQQPxT6XHFF1uHfLlOkbek49OABycm4K+1CXeaXJXhelYdIPieUbw027XvHVq7ItBQ6rc6qX5z
ZVdb7bmQOCYUa4QCUtb9Y5TUDMjLxdPVBQ8aN7A5Kc5EMXwMdr1k7L92qVeFJ+kICL4UpN4IIV5M
M2Afa6gKOi6w1Qi7FirHLtjzI/UGB427Zh3Dzjh5A0kanDzJ0MYsOLoXGXO+R2qWCZfTkuGaQbld
kwtnm7wG69t0kpwbowWK2gXP+ZuLfd9vBovUqOJ48I8cIxgY6iqdRjB2dfTQVDW37TBpQFCp2VOE
CwrWkiG+DAHa98yw7HgzqVF35vEsM+S0BJ9IlbaJmCwovUcQGqb6vlkmIvxInqA150wjT3cx4Rc9
Aza3/z7LUSseu/lvcSY07N/SZ+xnxq9N+rVvRlz5E/wTEoP059Y4QonYRluSjLysIaF2HaNl8FYE
oLiUhedN3uc8/v0djxaiUo1lIrT4sgMjZ6grNdIGU5ySPmHp4uSjqNQH1IThQN+gdUdqSROFfvDw
MT3WQc95/EJYgCIBI8PFzHbuArUJtYlJ5yEvhMmm8K9HWX4NIR/vXPNZd63eNwoOcd/fXeGjb5/3
SG/LBYSGu9cHzJsJB/CUzMG0x2sYlUM/88G5JmnZrzqLjDjeHMR7Wl8rSHAEQzVOM72460hDO0FZ
so4Suj6a02GFtxcWjMamB3bzoV5IRE6Y+wKIo+DsJ8AXrTFa9gwhT+PIkULwtn8Zq35HNjOeVrMp
46o9bLFks4QbM8nNt3oK5iBTyR/sDIjixVPS4YfIxT3rhucRXo4VH43Z49+1vpBIZZF3rmlKIPZh
zOn+dKJ4+CD5zOfIfZipLrIk9H13isU/HRS+tz+W0KNKxxXJ1liV3//roUZbs0HapA65lrKNSUF/
bFv70tGWEkW4YaVSwQ0LzcrhhHTuWhtzCv+YaB11gXg4UYlSTO10dzjrlYlNMK8qyaUkj+IL9nKV
amcwz/q2ZntlF4piP80m5UbDXu0q/w2kihhTeEKdad2PDN9vTlZ9Bsjd2LkB4m23+Ck654t6X8kM
UzoETlnZp3W4xjO4NkaBCZP1YRg2q0pyjOiEl2zMafTvDp5bwjCiQ/NcZ/Wj1WmhdO5/dQsfPZLw
RxidyTPOcLxLCo3YLeoyZO9Y3QG4yeR3lv3oa9FXsyfQQbH0/aPAqCSe4NwZOsHXyajZXj8LWHHO
JZeo72kNzbbyCxcIUB6wOIuX7lOFL4AOH7aZTPVfi0EIUwwsGPFDrm5ieKHSK9nbPBzeo86AUt/v
SRsLSdWD0VenqvmlX7iTmc/fPJGQSXAXmMK/ysruZ2fi657A4rjzjNecBgFpBCBhKHM93EHHa+29
H7z2lXzXvu792kAohKFCXCzq+Mn7rGIgGq1u7UKe612q76j2Cf1qdoYCYd5z/60afNnKgtiMptse
RCvXNwFdWnspPG9EmwJviQ2p5Y6aacfna1QGYIhR9riSN+4hGkicz7IrtKx3IE/eMQg94Ezd0kMp
nTtV1+bpwHA7ArG6s3xqHIMY0VjmEmhk8gAckjWG+cnuHFI3SQACf9Y04/tHwpaPu8YR1deLbHgQ
PoNmWFyOE/uEwnkqic411o2C4/jfeKsDnkmRxdGQdF2womMsIMG0qCEZRu3a5bGqTcEBbOLCtQkJ
jR3vs+Yl2bwhoEJjyFuWYUJnUGM2tLCtUc8hbXyZ0eoAvclGcgsGXZmbh65kxJfDsoUUSHcjBt4l
x3DGHt9215e01OLPr1zliudnhtqNBjbpp7BAHpAvAE7adnkD5qG5w1Sb1jlStBl1X7tFixoAu17x
jO7Du2RX52wPYHdlpN1Ftd4cD6zorqarQ6Qu2ka3CdFCkcEBLBeXPdHvNF/6n/AagD5iG6dBqJnr
lpTVwGxcQWIy8ASGkT40KKuqsNHtltrocljK5myxNQlVNsk2B9BEjImiM9MHjFXwQ4SPxFkc+1J0
7yLMw4OZGG/XsBZecKZZjPVAMpw4fIO65bhfzQo64MLPBt4gfVZ6Ssv+Vrtyarlo671wf2ii2/hF
p+CxuCfaTUf+zOQzI/XgYGUPHt3wDU3e4xwwQb4oH/EBhEFQ4cny3wFMu39ppZ9ieJM6uSBHeUqc
ZPhMdNZs8b6FNOlv92Lsfo5tzlLk7crwcXgTiE675YB2dN8/B1LbCfSWMAwZt0+stMiRl3GDm1VB
SsxtBnAxMBsTNkRrcIDk4nJ+s64PPOreEPWd1ui8hGfUsTWHyJl0Rb28e4OVjKXGx+ou7q10C+uR
0QyjKa9aWHNjmBSkslHYFXuxAYS83wNMYoQORipG7Nf23mFSCPCz45piN5HMqhmbS4jqhZ+W4mX0
6CPO0SQoLLWOeO36p3t4Ju7KyDq59oTK76zu1eXuVsG4OwAh4lebMJPjWWdRKuTpqdp3MW+rvQug
VEPtKQgHfgD20vXARRAug1l+MMrXeBgY/BfTQ5Rh1NcLUMRQf+/Otf3iLa3fFZU+R3LGopK5E2sS
TKbCWgZJw4iPGsHv9h9YINfcIANUaQocCUUevluDtqJotWVHfrCjnrkaDb0kwBhmFhD6/riOUAK9
uGfTMgfWxL59p140OjeDzpInIuq+cT6nVvAJU6lHNAwmWdmdBcasrxTTRjEOB+42ZUYfVtnRwaq8
a63IdsqArik/+Xv+8uzXg75o46Q5N1CVl0GpaMrJs7RRSEBY3rQXxFbRuwwYMiRd9973WPMGyUij
MIYtC1eCOkk0iViEXm1HjCPmLYMo602sNgZK34raVDe3VmqRsoItwJwD3dhDkTLi1HLyMKbD/wDz
Tdt0wwTB9cfOtofJdXi3PEaycvvtp/MYUCAtjF85M/pICK22eL0KdWysV46rJaR3YSfB4qs4qfQh
TiLj9H//ZI8PChw66N3T/5RT7agCNi3SK6EEN/odQp5/vIQJ7tO4/hswdEY1gyN5mjnVENL139ee
0ep1SxP8ZP+wFs+6MWPflKpYTJoznu9MHPaQ93GIcx7B6ZkjaUHJmAlInPziZ3SZZlDrvkHofzUI
mOwkGhOI0x2WDBCvqtOFuJQwp6Qc35ZGTyA/7WcfiOoG0YF8RPpF+Txe2xM0fDyJlkX41AcF4Aon
1qJpYSRjaPkNbZWQCbjHLvr+XCqGgfxdcazXOIhDHVNWoBoW5nPrfigt4G6RO8RVyaittQAfbphD
oYiKlqnVbBcWiGcYXEEpQekG89bp8LDQF5l07WEhR5KljmCoVDn7/tR9dMEIg1iGOmWJYPYz6Rhe
ZM6K6woHcWifXuPQMjaOW954wqeckuug/jSayBGY75cg/4iG7xnCX4J2vLzX7HB4fsb9/NOsFgBx
dwCDbr0LVe5zMMiXDq5mFlbeO5aZS4yH1+JL3m6lz2qUyoiE8LFWaXB+qgO1C9a6Iw0MDLJGpNGI
lzpjzt0m3Tyq8m6qOH59NYnmjFG1lXvhpP1hYrwyY8XaIChm36KuDTQD3uOHBx/bc2QOnQ3o2JYY
vw81shz1GhDgyfzcdd6BGPHk/6PVPkES01QBxSJgG4HYX+WTQUbKdOoY/Nn5IXXcRXQvw7twCxe+
ida2z8SgoZdLoPrmRA1AzspTp3OxVMnmH4PgB6Aov38yJygT280sCBzwR174HxAmrQm+0qVK2Orn
i1FyqLrz0mVaf7vC/SAtBnTLbVEGXr6a+8oiSem7/wT1DpSA+sQsllhSRvomHqxaB+4JUzn70q+X
k1chA5LGrQu/9eKb6f42WiHv8EVhzcrfNNbcux0508XvIEW3yWS4durcWa/9StMGJXRV9kR4rWxL
wtXIbe/Rl4crFAmpS8D8bGcT7qfKFjRo+loivP4fwzS2JnAHPlzSiy8hgdb/yu191XofH1Ttc6MH
4HA00CPMP2Voo46q2WrOIzzTaSY/anRhhb2bBChhXzi4+ktKDiI0vFFiqfIRxA30jXOiQrP5oWz1
9TBmoXvdKxdtLar22u5yUYr+RORRLdnaBhv4TNBDntOOGRiEykEr/qAgnIiRSDnEj5zdNDeSJkX3
ipjkv+rYlNiYuBEnEsjqdWKXzkihENLZLEVrdBIwinDrJF1PGYs/FMD5cXM4CfvdjRRRcL3WIu6c
ALY/swpE9zu3Uz81L5bnHZ1OTilK/wWK3vNXgpTwRlJd854yqHWbiUpK765HQc4TDVXVw60a0esO
LCdcV2va4wL0ewBV0e2n07ybDwWXR1tNd9i5jplg3NV2XEETuvmelStV2/6bz5I8bvlcFUBi7brB
NhPK2E4izgyf40yG1/kaePAqr8VlBqqCs95q/cV1xa53P9LMbmK7A4bxOK1L4hEdkNPtcNSk5LC3
1rIrrqan8MeoGlbXJklniguVv9pPbZLUisxLKz+XVxt4Ua9RRJ/R5pAQPv1XIEfeKKAXDQw5BiCJ
I89MO0nGmKguXnM78uFmUJoNrt9nfQ8Ngl3zekRjShfuDjcwfnpuP8JGduYrWpe4TX3i6Pmhp5oc
OvZYDwzOUicstJgk2zvXPaTjwpWMnuPHepy0JuPQ217uwgUMZMHJB+qefVrGXMwcqybkihsPSGY3
AtH2AluFDoHCmZMeeJFo6UXPsWLoBlUOAANZIzWiYkzGgyj2muIA670YWoFpXQ/fDEHCT/TWRpx2
oIsMNZzSkC1kWKkjMiVOX0GPE164oDGSFHhTfq/zHg3//U5z5++uWIqprJ4O928R9pLqGwdhFyAh
whq2iC68nvUQSqJTG5nnKXS7NmlnkO3UTbNL+5AlrExjez3JabgGcxRNvQsjhTV+IEu5M773t7l/
UPT29Iwgc9WENSD8s1YwELBEkGlY1yhlGH1/JPfrUi0dP3Qyk7EaV909D6N0vsbwS6G8KJHCoRxf
ShGdwEjzWnaMrfFivA466QvN69QNKO16crKrmp+VNViAQYtGMFpfg7WEA7PXDnwCXKoJ6A0tFHqw
eMe+9uOulXwgPJ4lKedpY1dhDqoZOEB6b+TLVUS74Xl7BErw5CjJUDH7TmGIncRVWESO4dHTvqUr
giUVSQRUWXY5KCB/a3N46LBr1KQnkaPGtcNv6Y+m+G3hSQ96qL57GG3NCfKJG3XPUfXzN7mKuake
Z9NH+t/i6+B8fj6voZwvaa701RDDz/nrjcRhiMNx+yxQU14dsnzSxhcWGS+NoPKZ0XwdDiRNL9YD
gE39zVFjq/LjdeOSyB9k9KlNItLA7IeSc1tjhvxy6HziVe2xgl7qAAKg6uswxv6F13BoGdxouRR2
n2N6XsztK2Og4vPnhCWz7QGFNuUTwGa9VD/BtJyvGuhyMwqQckkdZCgX77+LSbdAHCrbYhiYw343
GmKoOwfD7Zix+lsTGzmnj2gfc4fXvztdPvE7RCOHm9AStQ4zRhUOU5pmBnWWEQKYWQkZrew2w3dF
chAeXowM++Vfl1Bi2FcCgwOeiNn4SdFvcVvMWI3Axiw4+4IXCO86Vy/6eHdCLzJy7IRcnNZTvjU2
WGfBBnNizAmGIvMeg3InhrJlep07KDCspsmv6PgaOMSeWNkDfCqyPsPQ1iU2n7na+afboeJB5Afj
96wRb5zEaMJWf8fv0ghRDY9Dnpj4uru2IGis8cIo1zFO6ao+wRtMxy09OeRMFcqezyWNG7FuU4ZK
0ICFMOKLha/DzKfn8P2NxiXU3L0D0n1iD5m5Q4oK/xwdNIyVXz1UEBNeTFYMe6mEkaQLrSAcoyUK
W8QJRW0H1rLENS0C3n9MfHfYjY8Px91WyIIO8etulzwkoOJg7KoCJ9at70UzaKgtma/cboU0CfON
DLVgR0EBB2SPvUw+i7rTdPn2mgidT/Mbr/NMCsuBBWqj1g3Bg+1sWBfIYjV1RK9oezFGNBq7wsXs
T1ushyPhOc1egg/e4bKU462TRWQ6xJMGqGuytUw0HvsdK+LLJI+SGnTHyF9lAu0x7XVuHND2Iz/B
UD8lpxFCWLTTSIcEb7Df4aZAFDuZteQjmJwKhtHW94XHqoL6Q9aftVRkPGyrh0/byWsbrBuLgxbF
wFDcqRjxPxQhdZnzqwMitSSnuCEk4Xh/JHeiaHGuZiXTIWfWOA5+ZVEneKMCdPISQvm8xfmY91cz
CPfiDet6B45BYAWzWvKdzSYVZq7Pt1PytxkzSvAjROV5fHBdJ99T3lHUI3Z4tqPp9GIYhPtsBcBo
IVzLuk7bJ5QrSfeyOKnPEZNZ96b/yAuGHrO2ltuey1pF6rOXs0U2gBI8Q++rs/6fYDNC7SCu0SPI
3xDdl0DDFiGPCWwueLzuCkGqo4ywHc85aj8eUED7f7MhwGG13j/Q9vCJ+ACLyWFeo3J4dAh+Qua7
pyQcQYzlUnKiOdSSYqbOlOnTmey4IZCAAjj1hO1CoFmU3qNdu6j1XI49w9AQMWT5trXlkrJ422Yi
nHkky5DM09K7RZZ1uaEhzvjl7+Q1EwIPNSOEpYT793uMgpOA6DYddqgH5pyv3u2Sq0eWB2ZQLeb1
2+khSOAXFGycPqrEASqQHkufYmqSKxdu9dE63bVX4Pq6kJb1wCx4WGs1g76BTFjCyMlz25AczdOF
YDl7fafOVyIQ4Bf+7aiPtEaUND/Miri5meiCVugWrOkFQXquB6ABzQd0qMCPXskNZsgRGKBxUDsi
Jczhxke+FuR9JFEU4LGrt6loMg4iRsdTh85+HsNr6MDc61HLxxq9LZDzqcjFsQyt+7C59drSAFrw
oLBDDfTnRnGuwB4aR21B3if+Bg7xe0uUkyohx94Hfax6Bf/C19gH0cHidFRPqFhz3L77r7d3vssU
afT0I4JdNMukykOhgHaZbk3xmD9Hsh864I1bgxtAutUUXY6JLGpSgw+I0vprNxZtM/6ZbojU22gk
cZ4yoYblkX2vfbhUhSIVSJR7k1K6ygdNDBu1tohOwZasxlmJCFZ6oBtxH0aOwWgTpR0M4cvXDNEW
VPpOmX564z6mUpaUCQcPaGSeZepBpnZuuFOiGU4raVr5fEFFo9r6wo9/c9bCRn1v5LDbAjREYGAc
0nz8O7xN+j6EpXhdIf890FyOGtQhJeVHf13FvOARq8db21vwkUfKJ6DKu/DzQNBAL4jBVVMp9BZR
1t9pQVGED7m5ATaU/ZVBlk5gz6not/WqErmDQ1hQTfkmApbkp3pmMfzyL4gG+DOyDWWTUCr/ACOF
z2xcmh/mthfNmUY78Nh5psWnegicAqscK+hoIwmVajVWggK5fbJASoN8FEvtuS09QpyP3CdJKbyj
qlfH7NOuQa1PlxWTNrSzJr/T2HdCbCFOYlYsDndggLlFhijfpdHsFzZ7ThTR2dMGYDfios4wdjrG
BHAykXW8+UwCdc4w9MTIS9diTPNp/HOCZfskKGl0hwMttzLBNoTxIWfU35FABDWT/ph00Sfz7jqU
ckJ4Z+XZo+Mbv/cFjU8Y6StjC/r6suIE7FG96Hb1QNdmA7pKZBVOLUx/9JWdPNV7kuOnmUhVk4Sd
zjeDKASVg/i6ZgpJ8Dh3GsKNQ1LWuJbz9wIJ0xZpOj+LvWF9cuH/KZMhITqjSLA6vi2nkHYSpdlN
/2JINt29ox4UzGCh/BZAulrs8llZYDe4N29zf8RcFsosIuKw+46eCE/3P475aDLzOEUd99dGHxDu
MA/Fzcojr3DZZkGuRqv/kXWLkxk+Munmv2KIsRyRayq/8zlp8Dpe7WZZgDjxlw9oFT+MRXvYchX0
pjoOOzIQfDF8QJLuf5x6P4+dEewnyzj3CCRSPQC2Dkj2dLTKLH/IMSq8X2eiDWnntcozu35EmmVd
i307UlddiUKWRHXu0EnlrrNRsiG3vQAygpsOuwKRkqHV3zqCTPNxohVe38RRqbI9vGOejPPjzEFm
Bf+Qx5tDEIB9vaD0bLoKfrJZ32Ng2FhYM7454S2OvXF9CCC3JVSIZ7fNg7APD7haQZzDu5lB1UvG
BfS4qZSDBcB+9QuX0BeXwf6TaCly+fK5LsqAGLZ4WNQrjWS+z4ExGPeLMLiLoOpiAF5+vekK+KcC
eH0V53ZGaYuT5wIZ7f1MdMGVy98f4FnOggTMIukTbVbXUxMLHh/xpMxpxP7A7PbmN6rEg27slUuJ
euKOaorgpvm9PAbq8a2EmRbUhA496POUeUL26Gj2ZCXh/vbZST9o/tXTEJO8q1pSKLlWycCTmSQj
5rKTE2EeFqXJzrd9qD9osuARTw7oax01LpgqHhvXQ/QyFOl8CWxVCiqdO2zGiN3hzc1pgFtYlE3e
ny6vy+wEEcDIIyCJ6L6lnu8ffW59cWesVezd+8P/dXcds3QKT7il4LwArcc5kp1ei27SzopY/dGy
Y2kBnPOgr+StQJMDD9M2twP/kzUQZyAJzlwMh6P86a3O2pQwhnrkS20Sg5+ZZZNhhgOSe2jd4Z+R
yqY8LK82U9gHaTlI3NcG1U04wICFhMgj8jwpVwDwJEWBQisbgSbZS0R//Wz1xKFQPyZWtmxo1YGy
uOJOJ6tJziFOiJWjkpD6f251lFmmDF1PLH24Jp874DRuykwIEiAnc9HBGkxKnAhVN6iaOT00ACnn
4st2RgB2tviVw1bZ5YJDoBXDc7L4JGQbBPGqjzps8GtollW5sWBDqD/M8D8YWiG9KViApL8vMJjP
ywfp3joXGl9FKmjtd2WMfOAbqoUNdC3gMMmrnQbxAi1SrIuwJEdNCWxo5Qiapw64ydQhIM4/ZqcR
gbGS1J6PSMZpqld1cPEFSmojXjUWExz/axdQiFjQKoMKECXJhUS0EpqgmUXruf0raCC8fT7uTskH
oNYQ2HGh8t/z/9pbhMNduawHRTf2DGoyIXhMJydsnkA2vVGB8eX0XpStm/tPrDx06bVI3gJdKdJa
5XGUg4wqrVt4acIY1fw28cVRLNli9P6qaqFMGqbrjxnZHwv/TyPhNEnSSIeJaCyzc23HML2/zXNS
u/em3lpDETg2Mu04YAr7nrGGD2xleBRdcfnjKFBYnV3xXgzU0I/wkXXxkqJtZGI+/vxCcbWC/l8o
Vpt/GmsRsSvfA11pVDgrtR4mhYNpb2/ZsGS3XGzfauhClcGV9jMLo6CTLfKB+8i+/w6HDIA9t5z7
+jjs/8lg7UxSgtvnPFokO0OiVNOe/gJuc+Igy+FCQ7JQErOR4TcJUTCAIYGyhCWLtJ2NXeGlLxLz
Wfktfrl/UStixiNT6xCUmkhEe4oTpr8oktob5lDEz+2PXeYYPrrUlaaAqaIk9WaMJUuInGBNAcBi
8y4+tUB38alKQc8gWqfpd9l+wctKt5/dukICuhfOdNg83If7LjrHTdwPbM2/aCj7KISw4jiYfI9g
FP1Ynlf+OoNKJm2a+Xf5NXI9Y5j6mNBDzWYsY2pMk4WwAp6M+CtUZkdNmJE4Zs+QqBDVdO9ah7/a
LRBOFqn6Mik4sLLymCMNHOQxjBGzK3MHiBFRvcIx/x0asM1fDG+LAAP23yiHFSe+RIb8v49mNTcx
wwrR0xV7o/TcGBIKNTdNQDp/RvVA3va0+JGk2vz/3qg+XHc/U6o3q2BWAcrtX7wB73d+ELfdMYEb
yGpj0h1CWFiEIWgjv+GNMlYwFcQWIM9t6Qq6axA255D8UExd60Nl3/PE2F4RXv9zeMZimQp87wCZ
4YhH+QriwknScmEnqAzzUmhqfdKSR8cS/WvsbLnTFHVHfoZYbnfsE5OyFqdtvRLN35zjrFkwrAYp
XNB3sObRkdugQzJCMwyEAyMjv9fuEFGpI1RWE+jNRgbb0B08lJZssWWFZJ3w7jDxPmD4YRIZiZEn
mzEdRAE8AljQcWT0Y9QDuwvNoB9Zi3oLX7OQ0DOIwrtlaQWtVk3BgsD3T8m3nrKDEl4yjWrihNlz
BkeA9+jU6+97e9+vPCZvkzg5QBFBXizTATbXe6ljw9/LgQ0pRJ/QkU0LTbpwCarEWeL3YLcPWSxh
EYKH6ow/rArAay82AOyC/SOJrGgktPuHsYAtlUVg6uaqMFnuMeRszO30qCosa87HmXGix1qKCA2H
Jd/XgWcuSZd5f5eGevemM6g70X3qKNVcODzFumMAYrUPAGs+Ghvat6Gdc5Q/J1tQxXK0cgU6qVeU
/7P2FgrCwvm71WZ3edabJwuXkCX5kGqsyffjdqU2trKp3HPDd9fiRi9QwuGxqY0IEjGUZqdV4Bu1
7uxlcdu4mpqYOvLDQpxJp+nLP+GWwMM6K0b3/OAKR6GVocg7na7rsJFE2+QxS6uu2XFjOHK09ggI
6Q3IyX6TS9avT4J0sT5T5eB0gEoi24UcacZeQxVNie5dAEv1PPZ32WZZ54Kw54GATfUuO6M1p5Xv
VqsDeG/CHGhqRBjkGIOCm9fbApdbdcF4VklETrwtfZSG7YdrrDh8FrOjBCNqw+7kRWufIOOkFT/W
LaFP8l5BCbPBg4qbfjvQQuRvmMym7vl8v8y1EC3gCl3hRzjpm9gVk51/KI9PRtX6Dve2TYKV4HhR
UW35m7lrEVwVXSX6bkh9jWKbMA6d/QVQ1PDCqO0y5Gss+9iCMCo2tVVBKsJHHWe6FF3B6OjOmREN
opqppsufBAZosM/xIfRaKa4yDDMRpI+QOnXzd6d9fJGw8Kzxp75xFc7f6O3QROq6CFDE5Fphvpic
FSQZxi3xY9t5F1bL2wYAkMFku84f5oMWRXIpUm8wi0Lwj0YIOZrCFANrdjmsAkEwNhKEv4biJ/M+
rxb73TBIPblE4RhpEPCvcktAlfmOLUSmHMrjDYmxDfTe7feAB/VnZ5daLIhuxgscnuq+pYZ5ynLs
tMGF6c8JjrS2LY3wsWj6A+vKi47ua4NSmLK5V3ueAGk/f3PeiujwWJZObzeg6TVE7ZdR1hXytBOs
AYDg1tbU1QCVg7zEZvvTymvqPuOzBk9f/lXWIE+p1iNsxQOgE/KFVZyVFuDhUEVkMmngAEEClSZa
K/CVAj7zVDW2+r92AUZUhPb/fQrZ0JAvzbeCJQffPstLnNQw7es5n2pp3WcSpvVqQ+LGpuzSTli+
Afhvku2nv2RkxH8nTV4N/mnPjDzGFkLvlK0ejvQ9RZpRemC5n0F9Axcb4pvYIhRgRR1vy21CrXqh
a3I2l3arThzD0TCru35d/Tyoc/jtI7D5bl4YtyYQW+4bkh52gChwAx2is6C5LQhUhGE7I1DsxIVI
qMIFZY5tHaOkrZMfqIfEkuFJFd2lbQafyVV9/yg7CwCLtehtFJLoMUSFmcZr7hwYGWjQsxAHjZc8
kXBQAdMvrHHivvM8LoTBvcVvlKryxrFfOlueH5WFTFC2Uy3KYs8CBmaHGXMzhocjbv0Mpn7A22LX
/KitE2z12WnSEsJYfLbgH3V3VRgE3+gr+XuPR9dMjNFML8CzgyyVpxYLAwJJFLJk7zq9z3RQjJAg
MjZtJtXNzTXz9DTLm+U+kSgaXmO/pr4/b7rzZkG1HAqN2PTiXYLBVTYrdzaIwACORJiAPs4pLmSa
1lhzNDtu8GpEaKhoGON4SrGUB9LMyxfZXYCyoFWVwt0F4SDpRguwoVf/cZn5D7ZpUQUbCiUg9GnU
w1OAILI6Gp/i86aKpZKeznNrb8JD3rDk05XPQ/gz+PNx4e/5srK8/elM6zyV2gRTR74EpsTGRNwY
QCPCFV2DbukXdsPdubl0KucFICeegVRMlot3/KBbgK65x+D09/A2x5v8pbDU66gBCkhPE2+/3Dfn
vBrPS0eaQf0iw/AZUkrHuPGTc9inK7SbTTymDTUXvyn8P/LwXPZBNmOb66vTEXTvrb0HzlIqZa2d
RmaHBEcUau3XmLdFaOdt849b+mAjggI1ufa8HfVLTHctAN7u9JvAnQRHxeVetDJKZ8HWhcKg+odZ
b6FEqBKso6y/5lB9Jxykd74MhaQZd9ZmjjYILJjGVyBCXMJ+6yRua93dhuPrvMYeErR7ql87U60j
eBg8csbiZrpi2v5YvTJcVYT93KU5zW2i5dMfKo6qh9GaXAyXrzmrneNVYcCCiYJBlZCrIo7RihmO
nF/1Mxh3OMl3q4HNU1U5LmZeTXWGG8cUY0G4BCssgl9RXqHXHNgTYMm9iHLMvfhMJDM5OyI2JQXk
juqJanyPmVfMkjUQgWtYy75yCeg/NEjo59ImA1JGQykw1lvn7puvlonRn35fi0Ev7+HMDk6sf+Fk
tdrpoto1RvEGft4Z9qzJayCZGJ0kFDBvREMM+aT4urKhgYexJCYaFj/SOTHI/G7YAPSlMpd+ux8V
198IRg84ktwPQF/PNC9xrynYdWniKFL7OXyGWOiE5uTjPntU/S6sndlxZ105zvKuHgZZc/mcRI/1
e4OdiYiepLSbjev6J7AapbjRc/LVU9Ga3wh6RyyfznrgFx2ojFj7MiCxJ9b2oYeDyGR4fbAKN3p2
yofvbTD+YB1fh3c9/ri3CkxEI0ek/FVAZ2hoDf/7UpZAVmQB5/lmy6X0TQ8YYjiQzwmo9nlQ5Cn4
YFXessFuex4Wqm4TKqXOPMaMG9Twaq1kuirkzmhMHfeBbPSCCMITusPgAW7rZrN3l3ba6iJY0HQI
EJW+fAuorSAw/bwS6UcOoXPJgnevBmf2QeywrUrl2p54QWfYB20+QxmhUgGfO65EP1a1L8LmW/Lo
IN0AClvd/WT437KATW67n5NIiuJT/grRzQd1RebEys0r8+dV5sC+0pEp3ez8CYpn2R3MjSode/54
RBAQpwP/4QVWYITtncn3IiaEaWrSd6vbBBI+eKKId5l86toBL7SoqNWxR5l0RkcQsh5EdxjiRTBF
o0004Xe/kevNHU3ShXbUpRcq4jYMaHZJ4WsvHJ9ZMPkIr7m5wmqpxmT2JhNR4mqyQYj7R76jQ14A
RAr7QTCtAE5G1QwshEnng1o3OeizVd0ydNvV/9vaH73qEkOlcLQKD81x6bNrBQ4PCAXuICYST3W9
KN7LLw/Mu/fMYcQG80VuRpN71Bo7d7zXO9ZZzDh0PMHxqtgp90838dp07xJxmDCqM3g5W19LMeru
XUBf8Ums2dIwFm/zt0yIZNn0DMM7T+fy1J0Fj3+CEN3xwLL0SqDf8OixKfhjS184caeaA+O4ieWt
C3m2L/ykWaZ2v8oTmthTvYyVSsYsoIxUhNuNnqpfUTU9ajw/eB357FuJ9hVBARr8AOlc2lxnkY1G
1rBT+hjE+MllJTsKWM7OAwW4nMIIPxi1cQa6Bdo+IggPXEe2mwhRJKr5HHVxhzDk0LJ0f9IdbNWW
/2LacCBuI6ORiBc5ka82hTDpVn6PT1rwgYdsoezJ9jVd9ZzAaDvl0gnuW6Abtix7Z2K8xaFtCKMZ
4NVF81AFiar9zTMoFho1Y6FeQj2tJYjgd7UMMO3VHRsmBPQrmNawSPkgiReVBcYQz1NqVQSWWMQ2
kAiQbkEnQUaC2lQI/EljCtZPpm25HaoG+gaKru1cOM6BtdqGDCy3l1lf335rl8gOZNpKBHL4R4bB
2FjCcZnOvZhVgmkozR+SCSxvzKHnsJbHkIVD4Av62W4IjxtKFCL8rWFEyaDmp6wSilr9HLG2BCSM
ySmmJ6cRuKwsUjVzLIhcjYaxUyNVH8XR/eBwszRlUld1IWKlHEA3Nb64vVBBKGkhJwa/T8sUvc4k
z5hXG1kMt6SZF9X/e0DbxdqvTpKlixWh1ii/HRE82VZRzwTxKTAjy0sJwcUWAOAgMlRGwhWB8izt
OmgoFKrEIT0DJWKnJC87sFsS1HD5tzDeobdVqsqK69Wn7k7kzWtXInEeqhK3iIcy42VDA4SSqq6M
eta2tg4uaZp6PGDPhgkCjJAn7119Y05j+ddamlPovfg3wwEUCfOpu+2ac48cDaZGKooRj5enJZCD
7OnH3PD520ifKdhAV74fS7XzRBfyUyYp1vttzi8ZEZvU+Nm+GLEJmhmbzVKBodXKufiysGfzIJNm
y7vQb6xIu9sGMDRANPv4EvzwFK+Dlr7sYlpG71NvlPSS6YBjlezKOYdgMRVB9v4lVke2epRNw9Ww
YByFpJPSrGX19DuQw0P0sIdLcGakAhP1AHPVlprjUjsRU7Z2tPBK0QUXAC0YSEUWK17OTeorZFJ4
EaUbXq/O2b/pybvGm3pbR/D+sYdyBDDMgt5p+staIYUhKsG508Gb39e1HOe7hq+slTvF6lf97vL2
JaIiIUPMQcDHkn/KHdn1thHP1J8dAM7VAOQtPIvFS+zGg2ZkxojKu3nf6MHRN84Hl14GmRJMrmbG
MQzmxH7jEpbsrLXZVlMJq2xM4dVvFDeQUQYy1W+JACsuRk7d5yZv4Eq86dXFx6fC0nO/tAXLtqXD
k+RQB8hMMJP/yI1cVYCOYAHXIm7rlQ1XTT034A4LxApoc4czj6QsfGo6PK3pZxWXbsV4gfPaedG2
NGCcwzKVeaKrwmtFL2qIJQ+CHVVylLP/xZIgLW7vgW1PJ1wpqQrgJCFQkLJLR7a0yL+tXjNHHVpn
J+UnXoH7yQr8gkFlra97IPKeJYDwjm+VCYbGDghLwcximWt6ia2NYX6Vw7tXARwBhvdJJE/r7wnB
WF9wQwa1H2LeexKKVkzpu16yZaIvKaz14JymIvPGQIkIDkDOjRap9v9r7E0BfTQUEitoN1RRfRK9
Zu3kZXjM8UnVs9FeppbDHHXT96PhSG6+u1uABuiBvXE5UtHf/B9dnc1vLwzBQcLeTWY+zgjPSrPg
VzpVKoGIkO40+8BZkY3ukiGDrAgfOfhtiYjHUpa1pdm+aVc+eyUH+nTH1/EelVzxSVmBdn8VtRmb
snttedHtbOop+IDBDUAZB/JqM+R46vjwMDooGaR27f4R7p4OQITVEiVJibOxEQTQkEJTLMzxMWy/
kRqfcDX6byPLDgMrGtShomckkcX5NXVmuyR6mgLUhaX1pufa0os6Ifc/QY0hpgfDwFGisE3iv041
++2a62ZRRGhp56Ctg7VRjN4doW1FDNLGbql6kbfA+4rnwcpW9KAKJBQ0DATuqNdjjwosvFCfRV+P
fGz3lAGH9GRmMOtYDNNPKSbO+L3KGWdT0flqueTGIdeYQtm4FfyJN4rMd85FnWIiGnU9DDbjLGpr
NvJNoaVVyAUrNFBZA6Xn4SfaT+lSD+KbDb+/C5i4QWY+ejt87jeXtDX8nPdHCE4c7wXgkxtl64GB
NTAPKrZzOrxc3gyPLAx7BTtKULXnE6EgshTKXbY5iWrBRwooz0FqXPUCkX4ATAUSyNTxrPDDON7g
HmBsoeQ3TlrFCqsbCKi9oLiIBQD3v8Bd/zklyhdz6cStCXq5wr5ddwd+gOrLhDSmH6n4L0Dlx3YR
CzcwWui5sGETT3CmlNLaNG73pVmkrXeCSVfKKi+aUjWO50aRm7acHXBpkkBrNwrJVTB/jzy/wf1m
UzlU2hJBq1qlT0ZX0qz1LnXhzLKZu+qg26dNPd5myQN7Ov25lEuFcEY567eSXC16N7SmH3FybLDT
yDAo2NS1Hyi5zPDo2vz9lHhU+plCmCyUSXPOmb4TT6EW4T4lgSmLwa6m2M1fk8fTPiRhi1enniPg
X/pbxW3k61C7hgel1IYeklFrOaAWdV8GbzFHhPhyUgZHdqSJWaFh8vnsP0KFnVqduFhZwkfpvkfR
0MJMKzrBIrFW+3swOY/wep0gkifvvYmqra7kBxbyxaBshVuFaMt3wfaWVayx3g33QBfmE0T+aol1
Tpdqns7kWBKis06nxyI8Bb9HZ1CEJD9eAKtWPkZtkfsSilgTlFZT22J9qlhMMdysz7H9mWmO4jsX
exmrZM8i6eZV8f0lYP2n8px+afa/B4lfsVNGO0nL0dgCPuv875ZlX8UzOWaRGYkcgnMTSbtGku+b
QBJ2v8ucUzUT/DmjTOmq5Uxd4fg2vS4p9UDzb3mIx+mW+p0Op1EMwKjEyt7tCwbdE8YvyZIkWx7o
Lig9O2NipmqVVGdhw+YmTS/Ig3KEg/imtP35atxjNFZIknwApk5vKoRJQ1NmocXLSE/iWXFgxnvM
IHLAsRFungZ960eDuEXlwpCOQf8Twnnpyxay8yYTKmZg84UMRWPj95Huxkh8bmxQ1xfqFHyxVN8x
yKfApWNp4tDKMTDrHIArb5e7CxtiRsQuZYjtoz+nrp2OXw3OTAS+QhoESBLKf7bg+9yMJKso71zB
KQyoy6oqV/bc32JViVM8Jc3mnCMfJzzlM7717TrT7X2+9pp7s60rrnsSWHWQfJc/AMD3pp/OjBkJ
bKlhsX9y2Ni8/DmOR8wG16zVan1DQTSeabAnVwOAsZQSL9ZdOluoDJjxtyyN/ZVBv5+vVpKRSQ78
CkUzBk7F90v2av+02tw4zU7sm+RpHyjDGlxJblerEEIr/KuzIy/BIb0L3Zw25inXAkVAx4D3gJ4/
W48leLTJc+oNeJkr8Bf4FGxXs/CNpJvusx+V/7d27XqyvRvfMEonStvnCEy6ZCUpZFDfyUiOT8Wr
VWdHE4DFH8txdd7GDtM3BMBtmnnC6Zu2p2fAQ8dqG2O9GwQoys9TvK40a9MoTthofjEClWZR2CxL
EhLmt2wNn6cZixZbREnQfeZka1CG2DI4WNFlRHWe9VZbTdYsFA0f5yyXBZoFlOTmx7vxHdQrBhsC
+e+4mpamBngWWbUj9lD1eLGPNTWslZESmVRR85g3tG7lRAYY7z0skfzPg5HkdPCYwk+XqeL0ZeNs
Li4s9rrONTdZSWuuxaejwFBRGtdi+VJ82uY1U8ZeMTKK8qOX8OiQpx71yCci0FuEIWQr4+xPMCpO
QTeSNInlBiolNvXuvBg21+EiEDoRtlD9C8onHPnaGPRQS+0BasRDTQmO+Gu+30HWdT9CELzfxKwb
cdc/YD/AEZtW55ZDMmhCyFwXsGIk+Jevh6f5fb1Ua4l7/Y27KtFp/qgwbK/SDjk+dZdtjvTvgEBy
8nqMWwFlJenXDZtXjAJuALPJln/kHuL9dCWNL++xWGlepFnJZ5B8nZzRqB5cvboq4EdQhuhNWmYc
fGwywozXUpBvdp2rUfXRGkPd1Nkb1y0nJ5R6NMYh9uqLvGG8dY1Inw6qSQBLqiOLSSYD4DjSwo/S
xMvmBiXYANXSAEPse5u209+qFFog2PbURUTguF7e7jnYeIc6p7EB0/imhsKattm14Zt1lUPymn4t
gxnB5P9MAZKXu9JAaLM2/Te8xaqrvzkWwr5YA43K2nA0TGevM/w6Kc8jzhIy8l7iussYIHdyrYnu
4O7f03/hnu+ez8r07qLoPK5OWHyV7PwB4eD+OFSmrhPmxofovpPvheEGisE+m/GFTwNs8V7rS4bz
KRyce9h3DOHAo3BqiYJZ1nNFNx4Z0JVTlw/QGR9jqQiV1fgaDmNg33hHteJtW66ujHt4+G7RqL0g
ZZu/3/1cVGLD1LPWi2qw7QCPcKEJ/9laosCLe8zfRNCKtFlomVuesr2VdaLxTDccS37tEdxI748J
+lW2VMz45sgqkdAzPGBpIies+OiFS+mtomoRekziX0dGEyPZInQ5EX6y7bSnszYG7jcqd90h5TWM
s8oNIjQPavpODnQdX5vrqtA1sec8cwcrPBz32wrDh/MEKTEu4PI63qXa3OCpbMThOqyFGzauFVDX
WID3MizzrYtpZZeunaFdZLatIJIdACky1wm4eGRsHfTp5ysK5KclotyVfzOov5d8zOKOGvyQ1VCb
kVjmKPCfCmI+KSFrO1OY8e04552wbHKoy8B4FELXXkxh9sgDQw1FVxHKZulr56tM4gMO4EOWWrD/
Ec1rb9uQON9wIY7EfPlclJJhWpErSpxd4q7zZxava+imiAcFGdxhXzspyC4kcyQzDMtiUofiAwUl
IcSPxrxdIQr73+2IKOSLf6RGE7EIz6XH29YWQjisTbqeubmgbO+J9D6rOLylyTo58XpWgaupqlFX
l1Vce47LTpz4ZkB8F/tsNrc9W9jbUs65X+jYdB0ipiHoi0WOyXbmxNucI/YpQu2GjeMr5ko5+PaU
5sPCW8X6+GIRjhPdgO8Y4VgPL1H1+aJAD+pJYD6slTqsPBLVR1wAJA8ECjPyP2mGbzr+8bXty0ZE
DPmgyVzZj9RgvSN8cXITU/ifkjjZPj0ZZFzycY9plE3CMlQmx8snQsI+/NaWeJPHnxTZra9EmJF/
KXe4zHmezyUM4nguMBk3J2m3TZewFEKipeCXvAU9OVcbSfoSDUwbg/W2Mp0425UMMMX7LgTe10dC
CNGFLr6Owz9wA/uHpsfXtpL7oaRPgeSLAhNJC/KZVUx+ifYDu3E9De6aK007RZQlASHrgb3UL/SR
4K1aiO27F12/TKZJ93U/huRuO+SRijTIst+GwZB9nr4JzTlkBSgp9hAzaC0KNGRhKipGn4YbreFC
BdBovT6fuYMG5BkpZFxDSdfMR2zj4XwhMocTfLB4xiNMCYU3/tRK7NyiOylK35THhO8qtyWzFqbq
7QejOTb+R2tpIsuvkObsMrAeZ+0y6GVPYIjoge3Nv8jGbJ+O5oIhHkVyTcHFHRjzlkY9pWqKTN+m
wxBJoa3DolBCRsOz2a3TC5CTRPgdX7b/wt4iLdG4j628q0//gJuFyqqEiPd7iJwc+RmuH+5kp2ra
6UBF07IbXnsC5cMOrgBwmTaYWmETEBG9f1aFoJgps2Hl2wp/IG+VtzCxghcTP4F0GedXpRhwJut/
uyFxVToXJuKWUMdwz8m+QJ3kQU4yT4gtATl1SGqsFgUrfrmbsn5gYaqIxPm7YEJ2o+D1fDu+ICGs
3pqEv5CBACfjgWC0wLcPmTs7Rrxg+k3zNtLSydyz+i6UpQGz66eIhfGfR4GqySHkisTsR/dEdt6I
L719S0+abUktUOBu3PfK5cFqjqtBfCLRfkzNXLMie5mfJg2zovw2vuhPSf5A6dBCKnglmBrGA5n6
DlUp0XwrN0xuRv/d17xHEi8vRxbwrWTgAtIkmQ9BpvUDEt4ZCRz/rHvYEgz3DuOlAI/0i+gDsNCs
kGbflfuyVJ17eqa8tyC25j5GVhTdS7L6mZ+rWJzRMOXV6KlIPap5d6QRfuEEYL+Tb0+aR/ZLtwZF
upIVRPIbyeDJBp0jwqAWwB1RxIEYc2PuTmmUNP3LFW1EGArcj70v8iFvv+Z05ayfX7PsPQFfOoI6
tQ74pihMWb4h/J7iE9Epiljs0p9wbJpNtpkBWZkRibRfKp0R4V1tYWTTtRVGZ/Xz83xWFrm1J9Qq
YmFHOIy9xqb4N6908t0mAKcGpbXTN74yWoaWRnCZ35D98vlgIrFv4B6podoPzpt165u2cIY5Fzj6
DZ3iaCyUNRSXxS03MKe3Rma1udqYt8+SKwGA0aWHtU6Mht5XkCysKbAmjXfxp5MZOLNbXG2ysAYy
dugns8xKbEFw/e5Kcuwcqj/6Q7oklUbgqm2rkXZE4uMwybFqPMHTplfFF6mN2v0GMFbQDQ7dkiHg
2wO5Yo3fMEyU9IIq6+OcRUUTiZ626cqs16EwLkJFtl15vqD5d7E1mE8ZEQFUFf8VmAYM+vlWqWZW
//o3MlxosQUcJMAlAhjHYOgy5aOA/Ud3d/PR7sxDQrwVci6/bE4BVEW/933D9amrzEKLbhgmi8+8
6+m3aRWOFZ27coswXWevk6A+4d+NhkucnhdL6Lxzg0GwqiNxl0nxBW/p5wxAaPw+shbstYWwJkdo
01JxO9aztDbOK8Nx0+fKCeNnenYZBL0NocEwtjQuvqGcjEH5GHWwciWscj3VCDdt+oD50JcaCSqb
rYrRxUbJ3WlFjjf5QZ2SC4q7qrbvWWIitl+JjSSByEIq4Ab8I4ZKcelgmGohn11PLWsCYa3vY73c
RngN69TGt/DXhS7a1IDnQj8ClVqwzef8RFSchpiqy4XItjg9G8FkA3YuEtyk3lkuhMFW/W7vyrLz
zXWaYjKT0vmlGDAaPuzxHKYrguE1dv0M4DI1UVTm7ic9Fqrt5mHMj3Vt2sYRoLnBfOOBnEs65lur
hICuntqQaGXeBrZLLqLq0yxKNbiMiY+7yUPxTW8Kzodm4QvUKotoHhm4CeK81i3+GdOfPVICIop0
0RFxOK2LLyNGbZDKZNqpZTO35ryf/xqQmVIJZwTzbFa2vM7tYPIDCgW4t9mIyU3gYzEJlFo+V0ev
no0veNvVM92BPDAWmmXA08d212c3c6R0gz4vyFXa22x/4L/KoGQoRj5HFRMmdatETatgg8jcMIqs
GFCpuuQRNrT2gTMNWB6hvHpq/o/W+38ndK89LX+Sjsq0jCiDkrsNqulZL1PI0YeYmmpGciM5Ge/K
rzio/panxhk9Unf2Hvho/+csZcoIwnTOBkMfvty+f9nq78SIxvU/GS8E0J7TgxlOUQ8nEsOXSmzI
GCL6t+hzjaDxkjw5IzWIHaLB25GC9bNRtTivm3Z/PQHwl+30Fy26yvl62208vmiPT5BzjEq5PYdw
R2UiANl5Bi5qXhkZzcgrZAjDO0ehMhWnMsMYqkkSaAQTAP1wZrgwbx/0f7SM3xbZ5bCkjFaU4xQt
HK/IrH6otxXMXBvyq/+Ql6AYRT2rGrIBnrKSr+KsdsNrp0M6ZsUGkrE1opE/UQDQJqo6tTkNqi2E
Gsfwff3jNPGKXCWWx0Fp/2DWAqi/GoOY1Yx7Jum7V+8eJ7qATOOu0OWeXm9GoYUZ9T9Q/sHevgah
YPz0av2nstZc2dEMfFRgepcnvHhMthi0BWSMzMkvgVQvAQHgEA4mcxGhgz2iwGGATr0haQ5j0w2w
HzUPUjcnAqgUdy4c3F4LOtF2hy5jVorn14vVmFRsAVWlYYMVV5rcLop8hsL22KHSAoB7jqu6i+70
KgoygWLl1VlDQA9jf2hklDWy4hC+v2DgjXsC+CuYFNvpwp1Ojt++sa774+lRSJvUy7cJxQ4CSiUG
c4p47diFh05+zTbTmt3XY+iBA+k4N4y00eDIR/wZsV/MxjIwyxkA3qu0A0YxFXz0o+JrGqRTOk12
naG6sCR9bjOKxijhQ8TeC/q0Uk1+bH2k5xna1n2pRXmmEYa8/v7PWWHvKR1zM4x5F4UBkaS4XI8D
T7ZMssZeFSnxnugbp566bwtUGiKybXLWBmj5DWscwhreLnP+HBlq6iLXbgnPDAp40lWfNwSMfjra
4okl3J3oEWMzxUU/ROFdP3OqDLgA+rIYaCTEEUGPVLwxoaluX9ttwRV5bCCGY8/exSPefh5struq
EoF0uYssBLWsDthzUx1n2zxY7YRXHhNEbkIZsrUySCm/dHgJ3dP4ALBxmKymSI8t3yW+UwLDaP/H
b9XEUtsxcCPbwfs2/ljEC1Zbis00CtrhU7TsUkr0ghhWrhwRGyHoAQdpat27M4rwFv95Hk0pgSJ8
9z/GW7NOKwJ53fxenw3KQS+Vvf1qP7C19BJ0z9ucgtpvubrFbOzdS3UwY4ZW6HrF7x0Y4LDtWQL4
ys0P8ZWRMer4IMXGSKB47ObBKLazj+xBUOZWMEaOASCwAcMOnm7F3tT4GE6jMNnXTp5XJoQmDb1y
raQuBUWWs55+HrP2tcHdmeazLqq56zClhZa29splHpFzbapHjFa0RbSxyzGXcdL654Zhr0EwiWwv
Q/bNWM3lszDkoyuSz8OgD4+vD66SbZcw2LoMJHSUEU83RIfvbSLH5jkjWyf71O6sNjIZL4LagNmn
YQPHl7GOgD9s4jyg605sscgQAnGA9PTO8jIaPxcC3PQS9zrDmbEp0uWMLkE8gVYM6c2oBh1a5Bd3
6cyPXlsZSkVF5+qd3WPfumeT709bU9CRg0Jzf3jnYsi3qth9NL6rwxayYBtCMGWUuOmqe0i7x7NI
jNXpqMRWqOzc4G9/wWAjg6J8/QIQ6EESKm1d4I7FpkqsTeYfCPdYOm2ztN/YD1bJBrDy/ggKM9CQ
X24DHnf/CkO/4RIUWRSPMgFr6Mj1c4+Z0UHNF4xf707LYZpbsz9fwUkhrJycfMbjfhRL/DR3qneQ
Qx+rxxsyQJqBgzylemJIculsArCf1DshAhAg1+kdkJY7ic29KsrZ0E9NfT2/NLlvCdJsUIm4Putc
t1bITmka8qxYzuzui2zaZDVoVEGTJbjHp8C4thbJymiUt1D8LpZ9oVSCYsrdexf1PNDSIfC85gLx
nJKCwMDzHUKMjMud/2Jns1lr/LudxrDeVo+DaHI/CJvkONlpXJwBKLVP6HKdNMdyOZQgtdg8h2/l
eLIBaBviUms4cnVAzUojkwN3SQP4XtXlMHH0nWZkQhzGr+br26fYEJwiDeoEFv4N80ThNQHbIX+Q
f2NxKGS77vbr8Ios36ueDyjGtL9lxL8UkevSH2KJdSdpLgNCFkYwgtNUHvS+IfHJu5UnEHhglprj
aH5NyfhhC5k8lI/gt+WRCUCS4P51Cilt1uewKy8AwglQI9SWJIwcWkF4AYn41Tapvwy669yznBfJ
bvJ74oHW9cDRx8t1eWNPrDIMub6ft4i7d2mBYlIPaNsoauS4KCPEpN2q6HHeKKXWLOB1jEhur5qB
QPJYWB9uBE40Yx//pQo+qTwnRLHitDBCX3nuZ3+uQQij0IlmLE/P2iZ4qGOKBh05lTt9Ohq+o3kq
y6ooFH8OFBoqE+FsCrVUGtzFMLJE/jnkIH594eoGiyTwmwApzTn8Jp2UdBUfAo3R7ptIbu6O+9jV
zGlRMC09psky0j/E222N4GOQms9AM9m30+JiVxmiwhecSVwlqOzwwucrB8bp95lRT+2h5YC5NpxF
V+PFmdtJFBn0NxUha6qdwuip4ocI8A1Ro4s2JQHqPiqrDFZcAyDlh1dz6Ch4hm84b4vTNV3Nlc0L
dSrp2yBDzYUaQuPP8yQa/I36QjL7OxGtuZTKFZsaL+QdS/6BFbWbuZMqhOGkgOQ12L5Lt5dthUZe
nqfxXt0gmRgTwj/yxQFe4ERatBT8pnyPLGPGV4Q4kiIxmLkzqRRlIOYxV2YKdgIjFa8HSVP6PGx8
qpm2ef3Uue19EeO0jJzyuEwFp2bl6wAjtZVLgj2ybxfW0S/UedBCB7rGPUGR0C5BKf4wVdZJLF7q
y7FW/HfhxzHQ+K/kFWV+kTMP72qHvzIMmKXk3wmcQNI9yzUSBHzyoZSBP2z+yeHlxCadkyOfeNxz
rg25ypOFFCnvKTHRHGg8Dhhj9NAtwTHtAFPVw4MvIOsLlzlhksFtJaycglDr/s+bu3G1j6rp2ren
7vlpz9EezuJFEXOi3cYk2x9Ple70UNjzw+fuo3uFZSr/WZ3FSjL66wMxXgmXUNnvViAHK9sqxM4a
qqYtLxnumPxjGSiKLYh+z3fhZAMuakwzJz1/P8UgXWLebNyKcul4M9Gz3X1gRFkk+UvNK4MVJAqe
s0tI17nwI/Fd3BlyZXYjwMhke/NI+TlnGOVNOzRPp1RQEWxwaGUX+Ken1fEAgsy04ZTPtAZbDKjE
KaAOOKuwROTTvH3dSSaW3Yja3NieKF2trwhUViIlmw186RSQ5oOi1h05RdUR49rA22Sr2o/Qzkp3
GAruGs83zpfFS69YPsWJJvSE01Dr8JnPL+spDQq5j+sNYsVfpLRWw/QMkC4RAUDpscuwk8BXAUh5
bKCgZm9ZL5IN3TqRV0uROZtAYpE8yqBa8qbWsaIAAXfQoNZZLwwI5MhtH0RBCqgwYk4GJyAhpq9b
Bz9PMZSWrzgfLe0Dt/loqrvDZrwtCWaOEpXPJ+/mM0P3mnFK6eFvAd9UeZBI07VLg5Fe6mru7pFv
Gqx1BpunYHBIQO9UlzU85du/W8sasBq+WV4GGbZo/42Kmq0ufDS/kJtgzyvXC8v0njvAZK8ilheK
i/owsPkI6saHyz6Q6OUFaqCXdhW33GO1SFw1Gz3srNeZBGKgfOdPEVXFlvMJ46P1AVuKJB4D4SjS
40wSeSnQw9NmpM+cJL+fBvaHU60HskJvBzVViI8/G3W3idtAFh/urRIiLHqxxOkbvEDOUn3tcZmH
jDPl7TTZSOf+lQF9PHwEJYoy3ao6j6JGhH7xVbetRJd0CQlhNdjtWyclEhpiY2ONdJrwwF6IU7ZA
CCyVg04++YMFnDCBc1veyRfTNW9BnTSU/QEtQEVR84zWfUZWwzZKAb225WYHhoYFsfqddE3+84yX
m+qxBvtUMFNu/UItSr/DAcy5gSkmU2LC4fBY0KxO24SMCN3u4+DNAyxk3HphWwPLaLyYID4POa9A
O/LsqjATQKhaFKnbWRZoYTxwWzs+WwbqEd9saarX38E1KyrvT4/UcfbMJZp7hgp5TTC7JOIxG3Aa
39ohjAHebQVsSywWiBdTyLCxc2xQWKFiN+q41yQx6+CZc/YyCxsXcwKKiyY9Bk9rzck/zVAY+RGl
1DytTS4Y+qcDWWDz6cwkfrHXhgLgHcI1+3cy2Dx0Y5NV9d1+NcgNTa9InXOb6tpBowDmPMrAbdNS
3qr7tYfqlLdlEmj1X2uX2i43/71DFVIJa+XpSySR24cE/KE3ij0a+LpOCIphDE8pMpQaakgGsYmI
PiVhZGvfDAoTEHlTP9ZW6IyoOEZVrzAlgC+MMJimOPDwTv5YPN4cfZIj/lpUkL3OvrrPtOezAmNS
hS59m+TjEO2FpqaCtVDEV79FIpHjVLdemOtN0hzUZSm+P1JJdz8B6SYOvVdvEL/h6kB8X+6YFm0s
wY+vuzGrWe7417+D9ZzG7vKdd7i8SS90e/k165BA0oeu9JOMKbUPhL8TJCGi3A7svhr+ATMWU6Q/
WKVaZ8Gl9Eew/PTLg0MQoIUOnhRlfaQqSwklFyquGYRxQVinxcrJ8aICtqYJYavdmGIKOQoevB31
QTHlmexDKwblmJFKYwudQnjmk55JEGNWM3rUDOqZ88mZWxCH95KhjRCLvqb4a+ib4siK1r1AtZo7
nnYVGc4v1v/2HvzfriCkURvQobbkNP11/wCtDa69L7mHOjcDpcEgQOhg0932iIN4aHxzArVu2C39
2dcgvT6QjXB5OnrJ+FHCCms04tbPj4Sz+WKWTkkydYEN986G+WGIDLfM0pqN4DBVPy9ytIPbSryv
qO+gKhOsaJkvs6hk7BTKeOnpZQ3XJi4Z2BEwCD6YS7FJHzKgyPYbEMPxWY8OjkYnmnE6OYvwQfMa
KzOfg2xvUyu1O/dRLVnkRtDNICQUdle28c2zRvF6746sIdiO21lQoxRQDSdTTSdVdc//qkRvrMMR
T3d3aUDew5AK73chDrRRIBuF37YGPq7EXsP5TpB/gSdP4TXuYZkDYzHTm6Ug2v+CAwkqtIZ4sZE8
seHAuDp6NWFPBAes5FOXBTd/gTITGLYUNYXShOaolknmC5ODRqHQJR/TTHnZOfmtA/kESt38ETmN
XmjEXFGQIeDBibzPzBTDt62EC2n9DvjZTTtukKZkiU3CPzuaLH1t8f8+pbJEccwacnbjwjQV/5qL
kWEgP+eRUpYJicCkVE7TmIvwj0yNFZSRgKicu7XVN66bIgG41NeObLM95o6qOr0O8F5EV6GsmVWh
zyzL/z3cgeaufUuOn7cT9Aq9kK8hnBJs78wb4tRBbb95GcmMS/Ix32PwlYnCyY7NrcAbrgRYBC77
NFVXhqT9A1BN7SAgeMUAoyYPBnjfoq79LD32CMpTL/1/nH8D6I66ebiv7mET6B5w0jJRE6dEltQ9
0FH+cVuhNOIv2B632tCwY+flKVeiz9BcJsaCaw077xkM3/Pmh0ImdDYTln7VZRwKOQjdDtg45eUp
EfuKoQVl949Y5zEK+1SvqN+E1StoqD/fggtetNEaZ9GdU7kkCh3gVyMDezb0XhVl2Q9L3VI12JmV
ewg/ETXgNsOxlt+lUBQwujPmhrvlbEHTkcU2PYfeyPfksmOG20yUuMulnYoghpzY7dmO2Z3knFZF
C86UNAy9dQa/kIMdpDJ+M58mDvxhID9xxAyVX4cW4MP4PslfYqsBDb5w32Zi5/LwWmPl4OlMZZTR
y5bWPkUs6XGdx6tvWLQdw8zwKVgT8uPcA1DuDzbVYNEkWUCPpqzM6QXGTArPF/dKStx+LC3L3HZU
VdNfK5NtS9s/Itn6ch8EiG3uJ/MuLJSQ5O+Er54D1EVKxKzfbWdOdwJ3GSvYDMTZs7mzMV3VI2TI
ZmkiSHde//a6sehHBYtxfe0MG/VcOGXg4eMv7mFl907hdOkaBNYvCtSYSHLXsjivo/SpS7S1PQV3
+tAEUxKPKQBRyx+kgbikS3QYzMqQU580GP4GDXDzGxUwGabtw29AH2+Gp6eEiNHnBqBYX0F5FTxa
sqv1yG8absMHyY9YxLmwFE/xqNgoCCP8xnDBsk6tXE8GeEWbFB2xCYLvgXgDAlvjTHKjI+7bAlkh
PE6wREsZDJjvT1tZG7NLNb6D7kC/saddgBQQdhoJ0U1ftiZhR0DqwRf35MUJwl1grxL71EpdLyou
/4iX0WHKX+jWmT5kpKLk33FoXsZ8YvDtnGQd5vcGDlUkfEocu8dmQ4h7xCnM2kBwnetPlogmsy+n
NhdvXBa9PqgDq39EDla6Kd22jSDIvnlHiUtehioBdLfZw6wiTwF/DdfTWtw2mCtA8+kFqbhi1fID
C//jOLH1TKvbeba5jzEzGtTIulZkiGq7bM7D7/9IHkrLQLX01vVnMfQtUYJhKtu9ITlrHCq4PcMV
5UWlZYM+zkrBVmRAPsvscVep8IO5+msv+c2d0aND8oCNPHKDn/OoCHQBbYOc+JfuLc5kgYU0VQ+L
FP8c6x0fL48yGpI7v0GqRyq71zyVpG8bRsPdE1/AD1i6VUtpvzQU8M6YH459STRNhVraThrynb5q
fa8B/VoD2Gx6PzYIDTfM1MyDzjS+hCmvNwj5RrUnDmtbN3ATl1CqSRbVPmNct5fsSg9WLdTOMITY
e7/bK4VsoXHGXUpIirUy/CeKZ7Gsra0ogYPw6ELxSshC5/MEI6Cw1fwXH3fq61F3JAkXyGECxh++
3SYRu07lCnhRbwRx77Hrf7azMH6JHGFpMPbMRCip8MVSLjB1DS2lIRUQR1P2Vs/HmpT8vr6wYnJz
iyi6W/9l8+RDne5JuWgi6WapJkWfuYXzCoe7733b1pLqMu00yNQp6amxO6GyhOQS4BopFiIKL/5W
LCCHYJXsyhCKeBfI294GSJDpHk9HYiy7yaYf2R/OvX1mHUh3G9jR5NCI0CJ7bhJc0mu6mLyWo2FK
SQuv98kkQGyYOG+VNLEs2dDWlYw6GXnI7YEHG+vwVTS8pHpLTaWrQeLj0D9WeNsEuKiCn02YmJ3P
8wrePYtQOqJmKk4HgGUNQ38mT0qzVi62KGn1F7clk2YtLlrtd3CiTs509/wWtw4zpCxDrpika6k1
9n+x6ybCPDeFkvDpRMRxVFUTitHWEMndNindkuQbKimtcNKgsMwnqVreThU59zwRdOBK2FVm4Lyh
8MBNw69Iy502zmVrJgMDXdpzi66qeSJJWwthVGjtYD2gr+lH2HvRl87jAFEexEkep07JyuVKKqP+
8cg5JkZi6Z01Lb2UfTEuAq8vf8vZeXDUyOkDp7mhXzIfQYvuMkj2FpeVHlvEx1TQ7uG0KHNbgvCR
k8renT4+FfBB+JXJxq1nTdfvnmfosHgrmIpFSVrQ35O8E2XHMcsw9RL6hWpT+Np2ZBJXydMF/VkL
TMIe79wVAN+9sghT83hlTpYPK1YPP/V4E8B9Nr8dq7lOXJcWyBgLq+4+kCBM2bKjqOlZ5bvVXiuH
fZ+YCTSzq7mu/mjGYDEQ0LQf+kuJdHI7GiAVN3hW8ziPTpcz3INI1S+jVvRs+lHHk6Wb3AXcXC2r
hwzPjSYHvn0kNbWh2uEabLypUa/G0+sW3FA4WGi75FtQjx6cr02fNoPMlTtjtQC+phMwMUizEEvl
n6Ik6CWP/9ThIv9kzZu20MP+sb26X7xVdiUx440PBHc4qVmRXw9mnhWDE6kquYgW32AnMphxl+Cr
K6mYWBol1SaasWSzuTT+uRe+2Z6viYInIe8KTdS+lYipkea2AdigmCaUw6jrWvmY+AN4+X6yOz1p
pp1nArqP3eV4wkTCjb0sesXP77abxg19RNelY5N2XlWpTUWlkfIGH1maSFF1ZHaES2hbvfNbYpK4
rkT8A7pneZWqyu4y206CWcL4eVAwoMNgQuTnL39q3O+emVsgBr8pmJxhSaWlt0Xvk5YSNLCvpFlu
ymbRx2JTcpfKPDvr4u/os83kzmAtFeV0yHCNJmFDTE9ey0mpsa5zIAAiijUSo4i3wlG9kDcil/7P
KDfAyV+ZxnHzkM7qqln+k+uT8+ePdwTZLsN0jVSlzvVGtTjinQfNVaQQI0oqSefIPLa+bxaWMh6I
adqcOBrQ0QAChqBdey8LNaZCYpk+c/WDcEyXGAfVZs3z0FEagZZ8ZRAhurr9OzwVeahiEt04lljW
x8T+6hj6vpNo5U22o3i2fNu1vPJRG+4y46YusM8x1w/pyCRGecKb+OvqG2XTbmAmyzkyYOSi4Ipz
70QA6rY4YCeOL7458kM2coPovymOmyvoVzMjFyxcd8r2MmZdNudIpaWA+Ooiqi9+RGVVPPUK/yjg
ops1YI6+YeY8aQMhScopXoihHd4JdU9T95GSgNvrLXL9BGcyaCnmfv9yAtms5IGHROBgSF2YGH7Q
ZC4uZg/xOWQ2j0OULLvELXj/xS1pQL6amYfauwYUhfm4jB0eScbfQeQnZxLWqndQ3a2/jdunll9n
EH+Sjb6zAGe65wX0V8W/bJjx1IXJfjC6BTczlHvQuykgRuP54Sc9+z4xhCkjCD/7t4PDYhKJuao2
S3ehB1MBL3Iqw3QKoyvw+bJ5gnzr4wBeoHVL/4k0HvxdwCYVo3MxCOfsT4lY01OzFEl5jqIpOyME
mIchFq6wPvPC097B6Z8xM+uhgYIpqhUTU+sImgR9YaRFb8skj2baRpawffM/oeTvnnkXiEo19Qr6
U9+L0vvBxsMQflfQKecM4RUdPgRwCMNBvNwSjT5W61mfBvRk4cjj8sWMdyhqNqBTSMFNijConUT5
SXlpo2lL7JaRgIgKCnXM7NlzJyUZvXqSTP5Ea5u4DZzewm23qvm02Q3N3Z4XmH7W2iBeS1HgKQ8D
MZ4irFiy7GIEfzFPeW/4mzG+pLFRlNE+TlPJy3xufWJs55XMfOULCz8fes5hvGu/GNwQYF2oiNpM
WKUh9n7oFgAlqjPiQkOpp/n7S2mEuNRYp7Qe+Ti2111v7E7nWfiqHGYhZ8cAf5LkUGfiLeNvt3QS
BVl9ELiwY03xQGQOiVfJUGqZJNPePGovWwTU5dGTjqZi2MNeE6xqQdvCVnTaiedjfXqx/CO/3Egd
qUQEdLO0nZYAKJt1MOlKbfKUqCgiLI9qbKDmtFuKRQeJXY78W3135aIkpCwgdipcCIeOoCa4cDrX
4GqiV9xjYqOfnLYp2D4ZtBbejd2iDELUlUBxEWWw0n/rh8+i+uhz4hcehuy+ybZmUneUI99VDn0y
hMsolA0QbPcGlWSQCWXRJ0d9zOZ9iwGVVLAx9uhcwPp1KQpTZAFoATWHepTZbBNy3B9aYZ+83dPJ
13liJIKhqJf4fZcAryOOvHLkJE8ywK+PwQ4c3yIrVqCTn5olVCAisetdyjbeK3ZyEvl5r94PzQ4C
TivNPjb3ELHXpDXXnpWTD5VUBxW5p+MCMZ2QhlF+my0ZMdzUgQgFbvtLKmaZqfOvPi4blG2wr8d/
rzGW/yO/K1RmsUXsglCs0icCgGJCoRp82ZP/OKlxh7sSRNAWiHTUkGzWaBbLI59PVb62b39BzAhn
fLs8i132DZOtafXRh4nkCxwmJuB3Ta0fjiBCTuUShQkpLc/zpZFypDL9VwjSmEVvz+plZXwxUIHN
jVHYfL2iOcuTnSMHd+1w/WjLaKvmbaNqfkeMMp+7usQtWwL3bT9miJolqW+d5At4Qg9pd0WpD6eg
lLSAWR185GYSYJXJvK5FnBLCJESMEEk8Mc7IFGIoM+y1wdY6hKg4nf/0DKw4r7dBB7/TmllbA9XS
gbgAtH2xrtsm+isc7BLTln8K/1kSCN1XjngSPucAZkV3loRKY3YT50JE4JvzhqufhtzoJVU80RU5
A4V0o1C69l161e6kH1MtrkMxyeZqT3WPC/SyVzLw0daU7aLCVmhb3HT80//0Z3Nt+6RwGhtOkaNk
7oELgZ10hslMD3EX9S63zXhoxsz6bhIATFbUmuAFb78ryRm0jVWK3xCzSeDLe3ZXg10n5bfpOGTU
H/qwgNn/SEyP8bxI+GF6UESrwJ+v+JRQj6SIH/AJUiJPYjzMT30LpwXm5QI+cXFqSkwAzMH9Ivlj
yXqnmrtixYoqcyS8fKd5zW0oKoLnGzq8NTbLjb8ul1HjRufB/cNR7cRzHf4nyEqRW3XfDzbKpjdh
6uqKJURHi2WRpNflxqlDvvfB6hpXnEdiFOqahxN1qDZHLFN1psb+u5wFqt0aeiRNe3vNi2s5BkL6
0oNRflzKVrsvHxeIu4K/CtUMthJCx1it1WUWY71ypvsU5rs4MJi/nUK4nLdbZXS2JJY3QAAfZqvn
tmM2pcXG8JNhb4D+TQoeoNlYCxaq0bai2PBifEaUtQu9ynjt3DsFS2/LTgFHPD1ycWHwdvFEWi33
mg6kzLZKiiOLdt5gMe771iJQdFZxQbvn4vW4uJCxf9VWdQjGANyBlA9N7AiCStcP8SUflfp27H0b
PkPtW58n9WE0xXcJFfWw+Q874ZQQ4RUv4+mJOY8ClD0Zolm64VI9dkF2wNOiqvEW64iVibikePum
8Je2CtOedRCytpDmP5nMiiW+MbmEi3DFiMjvVOPLeUI/eJomTyfHcogIPhfNfpAGOsR0iMKHgtAb
s+fZfVNm/IwiLZMtTpoeY/WY2/IKRQa0Si0JnmYZsASsUVbgoDWRIIbhMccaDrIK0bGn7kr7s5AI
Bj1BbFeYL9obVuqSfxGTRUxasJFccjr7vSxhDe70vCq/+kzzpnFJpwNznQJwzvZjxtjEYzFmH9cF
Veo/ADjpcosw3zzfq3+55HaSaqQMbnDkKa2l+jV8mBPiPsCJMcSzd+IKGvCGJDsDGf+46ysVuqRK
7AIiwjXeivVxzHMswr3qZUUsBWtkaOZlqWUZYW2IeISrcbk8zVVbjCS98HLY4tiAzrXEuVZDqqeA
4o7Fd21Az3NZs2AaqZA2DWBbPVGM8SJWYiBwIKtkyGqRVNc0SB8nvoT0tMc29xfZWQ5gzqMCerwT
TRdD0qWHi4FzrQ2T/3vGESGgUYvi6NlTmOQTyx3vniCWlrflmxR0RbYqIaGUQDWCqXZ4PkWf0yev
yYyKFCfkkaJeWtFScpWAWvNjY1TWIElSU8oBbvSuLzI/0RCgGKR2CcTH1yJIqIq0QOyhbVJW4ckw
Mu/XrBJ8YjtTLFYr3O5YIbm3YYzGWExYfPdznowQfXYZnGl1pW3qDn/o1ckm3O6S1oVTpOhmcmrR
E1yF3Jp8rlvm8c0YFW3B6YXysvwBHudNQaJM88JGEHYW3CUkaUq3uLac3NnsDUoNugd+miAUPCDh
XlGzWhOZCowpaFfRSXLw8Nq6phf+pdnL14I7QZRdYetRWvqeOw18JHIqqot2M4HYCSqWr9tAwFJw
Gky6pIxaq73alls7ZsBKbgnnXKFbzKKcICPslJsolqxOBpSWV0pZlvFqa+gV5RkX2xZlziUUz8kv
JLbjCRpwpQDvbRHlEH83/LWO6lJwkliBoS++FOPKJplbHqvUKUi1WPWYycwLGAi3PzZJ/WPdj345
4OXhn9Q6uqUSlGv6JgpIFpwoBHEeMR9xqLaEpdnmehCVuVuucWs/isInDaFjEtDgZr6PqoPfKYxD
adh9RbdGx60oJXs0s0JqRYp9z3npv/hhUp51Ody9oJc6VeQyFiZoaTnMXndy9Kf6Q/2jqAWcWTE1
Ui6yJDf7A+ztkr3FFGv3d2HZuATvEsBZGhAbHGX38kgv3WzoFUHnkQoQuvWbGuuaeqolNH4zeFge
DqpTK3cpuY4U/mTbiGoWrEJeQTHDdE5bzDvnlv59hOLSrPBWZUfQNGR9ZDbPl0jOngiO+9+HSLRI
4bqfVma9YpUIocxccNjcgfc8bt3YKwxG3rWm+kyHiVW87orkd8lnKpy6hsZjwYkE4IUFyyRnTrfG
ppWTY9OpZYcCgYQLDG1j0xv6wreA3Q1sCsi/b2MEctju8is1BzS1ucMuiarLA04RyWnb3yieuc1E
l1LDKwM6jMujDqS8r7pnHLRxK6b2MCOt1I1/BW4UOdg8aGQ49UbBLy/uuIVJlv2QDtyRM/32bdv8
ViTUGYUgISkwkgjv7XFuHM+Cfv8nlkQpgQdDPehrC5JaoE7m16PG0n8AhAu0tl+1t8SrYkC2QyKO
bxnbFwl3PhzdO2BAZDGdmyLUVDLsW0ZoKWGfcfAagmwHWCytuIpla9nygYCBJj/6bk/m0IeFb2Ro
vOxtC5xv32KoomIU4LWFA9vMV3TnVZzOVUKmo5PJLr7gRFGtyhOeSx2Kk4v79tlHyP9ShfHCwGDq
X3FLohLCnNX6HZ4iHJyt6uq/VDwsMZeIZtMaeQXFp55tHfOUFjs+oN9fTXfVSAhoUwvBK6ZelMdp
Bq8CJy7QvM7jEUzSSzdMz9YuGAv25yeQvMn9O1MhV7VmPoC9KMjCAjWAE47FL3AZKm8+/27KW2Y5
htr49DqQBTvZxjfVNPCWuKSlzhURbTEw+1UZ1IF6j/FuHH6jN0FKn19ebxX+fVvmav91UafvfEdG
EwxuhFBy0/gTZW+mg5qQyeDjL7MZz2jp5sZBD++ULenf1u57Ba7ncZon4rDmTmnIBNKvftJsds9G
9xTus7RyyL0lIca7P4MslNn0i97ZJCe6lsw1LE3HjtKR2h/BQEBtjXmbmauBjwsN2BCToKqvV7Gk
2j5FrNVfwUw+yw82OJPqTGYsMyXrq6togzGdTVBe86gotbvxmwi1zF1DR8L1Ly0QYOiKI4O3JLBg
luBXPGMvR63P1X1uKm9gt6ywW3ZoUDHb2MU1NNztrBCO5BH8kEjTyHt3H4InZUoCV5EuckyW+I9h
kgixDKL8Dw8erSVw05yXd5j2R6d0vrc/9SfaPwzhq+0VrrfWI+GgzZZoz3lVfWOW+tGBaOz2i2du
CjlZh0R39eQbqsDJ9IFGN8LZJVag0Y0CWJi2uGIZbSmq0F/rIrgqWblqTZwf/D2twthuSMdwFzSL
IwlI1TojjzB0s3B0d7ScbgxVHAQqATkg+wAWZTROhEAUu/33AE19qTex6qSg5OZhGuYm1FU0WDps
SaSfkhQJeCMOQ2hkXskFdv8wb4UBFCK8XPQ8lT11g9L7RYxLlKXSmC1YJH64uReceA8zIw2T0Faq
yhcpVQelgWk3PyOztLGiNxzkSHAHDnzjSPiVbCPmIKJo8ZFtonopGYR86e1yYpSAK8iUGs2EMdHK
RyTYPxBk0BK4e8VfI+hYv7f+ZxHcgrPw1mZdNkH+p/v/tcwfcV5dD3l1j5hsD92ctb/2RWZq5AKa
P+tLxtLAp6mzby3psOThkobknhVOcV/HLLnRw3FGY3NUPufIsaRzq0NQHzufK7f1FJ6C1oLhHGHc
mNpF6effUvmBB/SFSoRaPD9/4M388iImwkcyKP1f4Ya7dJqRi8XQ4mA6PUpLCEonb2sdrHU28FSH
lHYhmtlj/u7bDAfi3rXNJE6O19KbyS05AWQhSyXSXS3YF6XyJh8lEPTA1VOkIc06nJe98PpQPIxL
9j0qSZCB9Jep3PpNjsZXub6mBahzG2JtWlrY1oDwBbsPfWbLH0j07KUObKbZ0TDcAV4EwqXc9SDn
xcazTl8HoeNz95r5l7ARxZXQxlfdTRdtcrL9J8oYPIXPnUzPHLHHzV3xzPc/OhvL+cSNcSG2v6N1
7whc+WqCZ9fKPOrWseHrMZg2fCguR+1LFc5+Qy1zzI0csA98Gs1dzsuaW9pQy8TI/c0YWfMh6gzp
Ef2I6rSoKlz0sGpRcEB+B925XlQIvPbXTA5mHXGMThkQUGE4tmdoUr4S7fmk+Xbg7W3OKAYnD7Q6
LZgn0DNv0dcaB0V1qNxla6GH+KkcGhZHEqrceCizkTmdZjzXy7C8NvO7RF2Jw2s7rFn/WzmDnG6Z
vt16JqYP6h18f9Hnw6b2IqJiQDYTIkxy25Hr8NhnDdR3CAg06xvQm+/XJiIk5AnM7gHKE+9jJEnU
x0fApvGREptZ09K2bSub+pOOKeiIjWbfY1iqfGielltgucxzhwn7a3l9M4UEdMQZPbHkL0d5rvCG
qBAWqRjAb6/ALFy7M9kztEseasgSUdJdwy8iRACjqrP6E4L6pUcihsVRQ7rWq8sq1NSXHh+10F0K
XlOtwacXegjweK1RvVztzrMI81yiIu6xPmAVxqRotaaorli8L+fDjDEpZRxY/FGI4bIx45GkxWqF
PkVdZbWdtd0qwfuePq+bSzqQFNvohEd9i6GIz3IV5xCejskJQ5Rb55eMDEB6CvNO/LMEd9HlK6GG
RVZWQWWektQQC5oFVnaWiCHLS4JLGuc53gh/YZ0ObMSKYafqxeQdLsb1H6FINqU86/LsOcLa+FW1
YyLEiCD+cfwF1MdRQskJPuhdc/5jA66SkQWZ4zwnQJ3RxY9VyMBph6qQkQLIgJQlNQocglMdBpmE
qAd9lZHSVdqP9cfI+yM2aZ5AqJ9i+nzCNwQSh2JxeUpzpzzJyFGMS0jIOEoAW4c6hSuxoJnt3dVm
V4S2N2gt4qb9v3JmYh6QmVHj9mN62qjUdVugGongpl3DLwnW6bNfBRy/zhTuGglaaMWfxsbfnQMV
oNHgh59ijc77IhdYySb2NC35FyO8qgb4lSqS2sSwiIGXfLFGsVpB5oFFp8mAXnClZOHtoES9bnp7
VJOLuvTR9syyaHZ8Yv0yqeIPKc3QNr+KbkVUU1Moxu8yf91sP6lmi/iZaS/oTsTjfpoWDBh9RdIF
tUsff8FGB5uVRyOK4EYrzaNNId0zhnC5KP9gt6oBDm2+bPtqGXeHXfK/BadPlLyeFhDGIgxEjRDy
L0GD+3NvCUPP4LfRQ0WLkQsI3dTRquuwpxWDeroOH5/bwo5Y5hy3CKxdxZX6C4ZOKHO7/8YrocpJ
DCUEsUfaZTnKx4i2SgMnPkV06SeaXCps5IaxT/M62kl0D+Yv3tJwa2+ijm1WQSjGLZFUdw8xk0xo
SacJ1B2bHJGUtQHJy5rSMqeTDGyDw5PG+St7NWL7B1D1nZl5V8FsaywEAmE3Ib2movyHxSezTIDS
U8Gii97aX+ehBUN5qQkwEhsSjLQzIty0qAcJMGflDbt9zjr7D/pOkNKbJHOmT0TTA1DHRx4CZEJH
uYqGJcnxVFILYf97LjnjrDh+/hPIky7VRghkE35aFn2r9+PbaJTZ8XJwjNe7f3jI+bN1bRnkUWHg
IttkFSg/FApssUbLMRJOlvEdKxIliOSwA7i/APjdOYYFXN8dofp+ehiPGAsY0P0mlWFeCr+4Px4r
IyxYaJ8+6GYHP7sDDytq8ab3E0tblanVqq1UVp4z2rh/VmCirx5cBz0iHd5QxN/r15q+Z0jh+YjL
UORl1UCAfY893IQeZi4TzOD5B5HNS8J53rOeT6Bd5XULWsNhFsRxGB90on7BayXjj+zdD9A4OBYe
qgecu/0LKIcfeBQsXnXXXQYlOs1ixHD0RKiNVzzmzEsUOb56QOBdVdsC70hnF0oDaDsTcDu+Wzex
a7jFSSyx+iRfP+AODArnOM35rhQbB3FQb0he2DUG9mw5wIKFhDJHpMbkM3GLyhDD5l39W661XgKF
7e8kx7o4xJT+f7q+xrtmOrzHhnUd1VwzPhhDQEdTjivUazzFFsUDdvbHWRxTzkH2PR5wMcPI+ycS
10vDXKBLDwN20RumTRcIoDV5YZ7NSMDYcImbV8pZCwIhAFuyl85Eh7BWxFCME2ASFJk9aBr2MW75
ME2+AVcYviugEypryJBuCN93wQU2kyDYWDKEap2dPJeM88p+DSlmhCF+eYzucS7nB/GsN6qwj7Rc
av/4FXAKlw+yWRFagbSLZW9P6SlyW/cRxFgjZeSzb+M/wwGWtWBPBlqw0z4dDTrOCUKdGJbnkTj+
QiMOGJvbrSHxpYVHd78wDM5a9oRRYLcNmvoLU8ljhj1GbJQM6B//8WR4WcwOlxxYgiLD/lz8vmRL
coM9pKhG37nGSCeAhtGqK7TJrSz5450ETEYc3AFoXadyIj61qGNvEvmAm9GxBpdUO2FNUw+2GW6N
YyTAC9UVkvKFHUtSlfvmtiZfEDd6sO2/goD+CNo2QawXVwr+X7sXgD95SD/PrIZsSXB4oJzSFZWh
v0a9X9o3y2bveDDLeVxCCT0I9c/isRHN+SygqSSBNq7AzOHbb6TPCoJLD5bCiaQZsksrYqSbwYXE
0FJUv4bV1F6hi1skPQ/u/T6Ztc59/AcakHvY+c/Y9TbnjOOLUfhy9cbwMoLAF7ugqEa/9r7r951S
A1JCshYU8tmPlZuZjkmfirTK3yPC/jqmy6O/q8qViSORcQPTOcM4nt/NNPpWVJiu3uyv6OvrEF6s
SFGTzJ6WKuWnRL6ywrsSYtit6ul3dbv4aNtcGg1uMKzqgFHIk0paCAdNceov3dBgeLBLMZl7ttAS
F3dewKpN/zzaPVknC62d4XFhjQjlSNVMv2IBDLVEl6GGepl2Lne17Y6iIr0TL6qwi9brHIJkOX/P
WU0m1NpCKnjpRzLJeJuraVQUin1GyU4cyrodSoSws34PjYf50zEXT3rPjmGtVb3r8w07nCU5B6PY
9NC+qDm9U9rXhXqTVop46iDK4cqz0B7hYhKUBBiXctlQTRaUi5LmaKxllOr0PjS+lWQs9nwFFyNq
rZjfoO2pug6ctNc7vPSmhnUBqQNYKrgv3r+9bZeswW2y4Nrqi+GRo3xo43N+yyLlTRMC11I48j0J
/e28uid/8P9HptWZEctD66Nzpmf4C+XM/94HrMAFJuzGirScEuoWSycHSYLldHAwL4gaeRigs1Ne
Km0KVVPLJasc4MVJh/iq3WHBNg9fSrd1ILpMArBnB6N4UGpoJ7LmkWbyf4POBpuB8KMUNTGxSXII
q0Qwg6azxJq+fgXKvEq+qoFbjkUFFXWPaX87ZH5EjZ3b/JiEbRy4q3nBJtLmq+86hfyQecobLel8
ACAypfGjUt1U9ZxGHzHoXAOEqugms0r1Y+rkv0yU5l5pYhHbNqJX/EG3HEwoB97Nuva9ravrzf+i
p86SIP58fynayA/gL76uYHRJ5ssmQZgv6Mz7q/ilxLDTwsfBBiyQmL4RtOoeZeyi/PVdgcJ+6L1E
lxGpMU9jcg9tXqrXd6cNtFkCaldKPIv3UeenTOlmnyh4PIBYsUN+8uS6QOaKf/ifcGfdUq29kVPy
XfB5AqpD04pUzb0b93tQt2EvP9miufMd1WoP1XZ2x1PiyzZyespfZRQHBFOOU1pnif5a6NTxgXaf
cuR/mEyWHbV+07JhX0uWfxR+94j9fNYmfTv4gr8zjogjAZyOFpke8D37yZLSb9HE12thXD1m2iQM
gk+0iihG+pQrQtxmoa5k8hYTMAPj19ZfRmCcy0eMzXebofJLLn58m197MvidAyDAHUmRvb5kOG+R
stoUtRhk+fcpjHVEuNSF1B2v8ls7etAu+NakBf7XCdgGPJ3TUZtdTLikRfSxbRViKS8qa+jo9oA+
34WS3yGKpVE4Km/u5TXpQALJNqMyo/ihc6GpyWZc592fxrZ2baxrlp40A0VVtSTyHkHfIBif4IBf
kBkCHkr+KhmORwsCpvEmjrf24LNtW1FuMPgloheEaKryiqHiW3K8O1jbi1D8287rh691XU0TU8p+
3umPNHJqg8d4/lB8yn6dHYEqVRIVF6plaAz9gM9o6Z/y4Q9W5S8UJ5lMQg4oHW+gii058J1KhCWF
mZAK/Qp5an4qmu2QIesptQOSn2olCYWe7OOJ7CBG/w01eO4mauXu5HIikC3bbvevRszTjst1MKHq
QvjuDaMwd/nHowCB+hElpmw7DHj5qxoP8aS93MSqKUrORlNJScMxaPbfSxvd268Gg+fuNrhJnbbJ
gXrPBtLIfpN75v6D9P6+Jr2AnlAUGyWLu7nU1t9ieV4MPsQFddY8RpDX6yuUCj5v3tRPLldoW/Mp
3dVBXQ2howD2kD5Rq7CgxvQn5wc5ZTzZlMbiaQrAUJQvDj47mLhrIMO9mJ9FQMJtKNe6C5pH4ffp
D85nnM3lZb2bM9v8AOiLYDDy6g777WN10tiQgUDW7E306fMMh1ijiHCEUzXoYqw6xDFgJFGko4ek
b2D+bhTJ+9Gclathc/TVh+3+csr5rBuo06oJRJUOLVym+VLgNHnzQuGozHSPCzQvt1b+RvHvsRKz
cNhwlBD5IGYFpvEifKWb4nUDIcUX1oFHfzaACYi+PaeQfWFg0yBkAGP997wPFuE6WRwhHKVKp2n5
foS66qAJVbYaXNua6OoCS6IVfamzT5wqlGjDOmUCflMUYdQ9nPDHbJtI0Vvvn5zVr+xEZO/lmkiu
qZyp+nnEjQubtDXoFdOd/SXFh8xm9lPkYEfsfwylWFpdFt8n7hgDmyHcCgASJqcikDX5TAShE+ML
wcELrYqHgkG+YfhWM8bEQ/SzS4agBFj+j62hCvGpNRsm7sfT0z/37XkhaIjBT5adFOGYR+gZ3FBx
TymOFzU3N/qR9+0xtNfQTTI11IC/aZdI+CzCd9FX+OIXX8wVKbhonMF7fINyvsDAdDWVCXNKiKPR
pY6gXNaTnVRf8PnISpOXuIaXDgcJBuu7qadOMM51WfQ/dsHbybFkfD9IQU2484fZ/fPZoHPMJ7EO
F2ko5yyTaW1/qK7vPSylP5uYvYIlvB68ZD7TubMboq/oGiungVnk/y3POvigFX7daiVf0f0SIwbv
8G3tslh+uNJQBHa2VwNVGrl3luCVnzvSysX1Uzq0eR5z/fx57aEKRM/n4HX41p3+fCU4PEjwZUJK
HZT0NzXAq9HQrSdV2ve3lKz5myq2xQYuU0xBofEtgvVpklxaHoX7FihMqtrmCpPtbDpBUuMYRnrA
Uu5sUIGZhnOaIwyC/R6/znEiZxkYdURqqhMhsLpVnaoL4R49cNffrEqEYI85XLNpTHl+dleOqDtO
DezL0DXwYSdiE/WSLsXmoyWTgCTEbvo/AKXCAgvEFWfs44IeRzW5nhqPooSEoLrtyQtuVCcyseuy
/W/SPBrPOp60D5Uq0CmPG0tnEJCLwr2OA4l1eQd4H4wk/xF8nvupCRgjF2X2exsBY7tqOFQ8P2QN
EVsghZ3qsAlvKbrNsVTA9a5Msa6NJ16T+YD9fwl5wVAZZcJNwu1/0vKt0UZs+qahCgSCKovx3GcB
WZGjp98Xo9nm9R/PcVP1AKS3G3RBgNoorGETJO2mwpbSHT6q2tY5SSSXJKPdNZq/i319nCx+TVh2
BDR9Pqr7wmEMzq9Wll/of0/a2xRcv9YULZXYKAAU7R48iBolaqVQfHG+IfD7+5prL5MgNIEhyMn5
nPwes+e9EswXzUSPf8X2MGb2uIcQbm56uotXUvAE22XDWm4/4ahc5jrfFZWEacm120+e12ytNUgd
F8Pn6LJhHK0iq4VFBWxoFewXnNXTBbZZnHfmdtB0kZcCfaCt/IlRSdfwVuZyBHcKkTiArJ5Khor3
fMTCmziWX2Dpt0nB+dBQGlZteTP47XIQOSXfrrDIO1GEeJY9LP4qkLZ37gv7ciOoIdPYqC/+3EFF
Sm9/vQVsViv/oem9micVvAQVVUiFSszuWnXdaQ67dfrxSSjp1Xo9EjEX74iGxSxmfl8FsCxKiYjj
uxb0Vtf6W5GbTYnQlJnljjbHqtUpA+wHhJtYMUz+nTv4iYiBUsKY9/f3va5gTRqUzxirHBCoh8kD
LTXc8ISVFBTrB4vKHDTWYiu1e9hRuObQF+PKd9qG/L9hTMROUP9kkP3nNhKdGKmxikCDWEObQSkO
wcoxKqChZWJ2koZVnCIAGt/4reNq/z8mWCsBLLIsYWPrmRBnkNhPcoe/+v+3a6NuYKHeh/fJQXAe
pZWcSVtAWK8sPaDhf/YHVAG9JGJjdFTzjy6GDGAJgi770yGX1NTec95+TAtopgiBwBUMrPFelOgk
To7k13q5J2Juo1S7WTPUm27u7b5v3+PlS0KviUocF9j148dBw8fCUm9sTXcXewERGzOZKlQIIQjc
ZYp9MClvWFbqex9nzKVATZfxgywBwaLmOQB0Ew3XmyDwW0yVo10CbIITWjzPkLOexkWW1kJSRYMI
nxOMTUTE9Z5KN2eFbnpiMYQHSZdT3+G2KHAcCvKGtb8zStvP9StrlcbDDo4UAcuwnG5HAKSA6WNB
vfRHFb/6PBn0+RM49bnk76C0+pJ3BuHimQ7/rV5fQfZ810aHP5Y1XdvKSlAuEqezTQJkLBUuNrmr
RR6yxl4k+z9yviW6LaRusIG3CupERVaRY88u4cww/z1TIMbklSkyb3ZlJgayks84f4BehZG+c7HN
RtrjkPmGseck5FRCnZRX/Xam8MTeOzdy01sZ31BL3MczGo0gWSHPiqzQ0A7Dm7DjfWajeT4grQt4
dB0QNFcFTrZTV6bfBPJpkgsw3/8ObE09/bLI2/pKhp7SIYq8MwfS0LjE1LmnVTUtHRzhQYQXgo8N
XfwPqIIfALMF/POzr6VcXzEqpyORvfIU6EcYSkPjjiKeuM6skyw+HlAJql/kaM+4lV7CB/WiCqn6
AIsJXeqqzGpQPZQcqp/jBZAC56jqepaJuuAuAUtAdjt9BhwJG7XWpU1wJsR/7jIGxxssL6jegb7A
igqQLy5I2sQr96+Ip1MDUewkedG9w7z6pwadZxwjdgGH9rNCrrCn9ojR85MLJz2gsemtdydv/bzl
qKNmgmK6ndScs0ihdk4+5MJ3cV0031XmWIZ9wKa4+bmMGEvh1zUVeLEBpXgb6C9tiV3SrZlbVNQA
PEBndJF9r0mKe/1JV7aYhyisyFxreR7P2AU6rx1mdm8t9t+UtxmvdUJdgoym0GclAQmEq+oSs+QC
QDnEFd/4yNLWrjet+uDeT6vBQ8zRIQGozOOamNGnO8nT2uCQfsYtShsMV7kzvarv3NXixiahwIku
21Ymsh/Z3aeOSVI1p+saxeNvT8MpEqo2MM6+QBYH3bmfWdqeU/FSFM6z/Mm31W2bcZsmcnCJhn+0
ghotddyniaVdesReWLiR25s2OGdqS6WK9pzhUHPahZMVVkl5JpcHK8cAGcizIPx7Ht0mXtGYk5xQ
Edod6UyZzh3jxFf2CBpoLHOCaNnN1EdKzz6TMi/5HtC6HdaJ5A7HIMJPFbU0fj68Uo6ts0TwBI7V
BQAllDAgFqwP7UvnUHymfNy5QUMTyS80I2+dHBo7n3EOD2TBgCr430ZchMOimQ/jurYBj2absXue
NO07n3wOt26hJix+CTj1fsohgtT0cQFZZw0eEn6XUtU5T6v1nb75z1zWCXqYt+UHlScXDvuMGVLT
pYdKhcXozQi/LV+2VfsUbHYLhGcE95rGYz7aBJpR2xAAqTA9xq0lIYd0CNU4LeuyzLLO71GT3rOI
pvz6tt64jiuac3+ZMoM6ORfCh9tBnTFFwjoSSUZCmorWyF/Ju8RKXEoizXNIau4v1RwbjNz1cVoe
kR+xbYRBU365WrS9bRhQrwufnKjaTFFwtL5IjXPWPEdkheUQa0P+LRQ8HF9+tBh1ZxU9XUn+Kemw
9bNKFFBBZa8h8ugqiBl45SIl+/aEdIwDo41v27iYGk8TLMJYjapXM30Hg5twb7Fg+NnDzhrKFluh
WOtWUKTSZgE/692HOQesj3GqTceJV2uPEWGJ5NKg7GIoF0y1YJqgPwPQwE8ALpTnBLedN6R406xY
oGn4dbyiv0cjB9PCsjEMHnlspRxEipIydudVP69P+0fczDaCDw4Gi0GaQEfCnF42xCMoUvr3D2sk
bRFFzBCqe9IluSvYzEYjYKWNSMm8ElhgBCAC9MtkU1+Z6RMk1HFJ2MvBDZtw2nA04tW1PsMvp1yv
hXQXfatZqflpdGmzd2vpbGLGWGzybd/w7Z+8FabEijmqJmxdyYZ8hHhbRixiwakm7uKxdbjofndk
6K5EtXnSdHS/cT7TJYh7zweXhnZEAqfTe+ree6kIZyf7uLdgvKlY2wOXIeSsCKm6jMIzHgums30m
NygJ7iQhPAwHRrkd343cGm0LxtxPa8pXVDd5lGPw04J3FaDrxNL1sXB/+FKcErpOeT9u0qe7nytm
NP1Q1/2WdUeWzWVAk8vLS71Z2fiPZv7JP3a/9PoqO3iOGNCM/rIgIif+T4PYfjI377T6b7cMQRen
48o7teQutWnxk4vmKVJEaWqVQA4ZhgeeAVLOK5XoFrZK3/fp+LqohsJOcKJ7iOP2N8/gAEfBiOqD
4kzLW+t8Ki7rYjqjyPeaPR1Afq7wCjF6ioCoTgo75pp0xw3BL7UvayhYKFy/lIihMYZ5W1nuTyLc
2lLeT6qQT3Vmxf53y7+wyLpPEFYtXMTjK7qd+jw/5h4+NbS/dVHByCyWpXnadzI6aK5d3fsu0tRl
h2/GUKVP0p8eVbDSkNd/2/XYLx3I0bH+yd6j6bEuShDPukBp33h4Ce/XnCviqz4XgwJpoktn8KTC
aPfs4R5Reew0o9JKDrFSu0cqCwTkku2SndGTAKpotgIb11fekAtxMhujDsHNcdNefj6ac69oWF9o
Kb/x3e/liN1rMrDPDCJbEKfFfiyqBR5e3Dy5pfIYOuL1g+/XiZJBE+ipbVrarVB5tWo23Iw0iKvr
YfnO19V/y1zeB3wtOKRmlw0k7RK4m04LCPDnDNzpd4h8VDF7/EORTwlZyG1kJ36v08x8+iKsW3cU
Cd7wiMN+Sgs2D9zJSPpt1KZIOZLt+cZgPKcknb4vtMFZhn7Fybc69hdN7FlCYY6BaQhUBOpDh0O4
ML8w7+mqLGtjEj5n55+u8vmIWkKiLITuR/dp+QQ24lwfqS1amnFUpF3cEINkfuv4qrNMZdaVpXON
MnSRjV2SQJIgCJrY1hY5STPLtEhRnh5UdmbUJDo7eNWFa3SGjNp6DfU58GopKzclBoZowiQjicbK
lT0B4VVTepitxII17L9wjblrLHz7ua9mt8v26hhQe4IETT74rE+STLsPOfckTFdFYDMNE+jQp8AD
VY30N8BDFwcyc1NsbF5Ylsnfg6n1DHZ3TzrDHEurZvVD+koQbj3jbppr8L5S99GFHyQHFMfHwt4J
8b26nnQ1306M16uC1kfMkvB+Zg37pkwdGAn2w4a03Qpm7XNuXB39zPJHJWSLEnhnqRRt2/YIA6Og
fkp8ir7gC51uChavpBMMQ2RdNE26iDUqSEh+xt7oNTgJ9Oa/dn8GiVzsSyCdIb0qvOh0bJq0FnIa
Oog9aulF2tpDj/eZUuSEtKq+B2F3anvs89A5/L4KRdTOAl/2lwDk1Om2bXI01dnT/iYAXZYUmnaf
/PCl8D28MfPuA0l07gnvxNqmZuYWDm5dRnyGYeMCTtgEFyg6Z0kv8T9SZADYjEstQsLnYGThwFZ+
YahCib/79NJHsWSTsHal+GqXrjeKteTlo/FtT6L9JAegIBOup844w5Vff7zUm2GFuD/QrQmd+9sp
Lc4Bi716yGAjFkJkfOzWFy5YKnSNPDEYdU7typfAcB+Xw2vIWhuXaHg+qMa5BOA3cX+4CsIaHlUZ
6WIpZnmZny/iwkUSWLgqKA3L0TQ3HFJVJIUvZKmJQ/XHyB+Pw73SvYK4do9wOPmo9JQJuRQZEgZ/
8MxaXo1WxY98egmdQ35qfDNjWoHcDO4doc6LA6TEgK0zxJEHn3R3GDC/0LxBtYRg0HKmholPdfFt
REC9NjWA/8TpQSpkiA81hLT+5C/KisMg00yxngfIdyjecQPJhllJVdY0SKqpmaD8S8oyIs2dN+3m
JpAjAS/FHD3ZsPWXLbkTqOv+bIbYeraJ31/ZlCDsdxnWM5SB0CVyMw9N64G7tlstKyvVV3KrQii6
WVsZHLDzqSHk1MRW5c8UJzBHNSe7EpIHMDRtO4CVMJYc1KCRXbMpfYwhGTqzVuOH050Dbh5IF70I
4xLGMhxBfR3d+azgRkHtHjCazEq0RPIJ4iH8g+wujXEw27vm8u4WzirCRyAR0e5ISSY5FzFMG5Pu
XyNzwLRwBM/89esyyRF/KMOkFNo7gthXBk4zjXQSBQafaHndp3H7l3H92/sN/ZqvA6mDR/pxp9vO
xQh1wsNGIRZigckp3DjO7sCYvWMvRCE925S8Ek8OJGNlJjT6RxfRYs/+gL2KLDM/55KXjrCRr7MG
74KrqgFsVbhqFsSfvGrGHxzAf16petamNq76eAsoq6QkABMz+3bjO3T+ISHR/pF7j9Z5eYniErPZ
39lzlgN+XwR5p5h8FhIoBKk6UCnlH1MtIV3hlAGcTHS1xIjrwSEBwryH+msD7Q8fnWi9jjKj7M31
+oSWC7SYUtTOEXko+JaoG25epikVb5WpcVt6A/S9HkURUMhwGj50dX4aWAipqwy9gsMaQhUJgWPl
gqqPWauxVXIK9x/36ghUqr23JSw/jrNukGqKpOOY6AdHFoOyws9W68ygdqE3iW/toLN7l3SOXsU7
VEeOq2GNktc6nnL3uxKFt5aRxWBWOVKUa+VfyUGsm6bsbQbpUXpYSjnNqEa9+Bwh4pmE3yhvlR5l
Vu8T1+wa9vnvk+cUE0kWJzWX0OkBCGcg9c4PETgGnEAfUPMI+YHFu2oNvBWzxUDDGgBLrAo1lbl1
MCg+7+9EMSCR+7UADQ9Nw1CTj+4wxFuFfCt7ldzKEudZBB/m8kn9n6OuK5giZDCnpo2gmJNhpDGW
8QhglMNXzcaAnRduPe2DAQ7slGgT4BZKSqADtQ4mffn8y4NnsMoAMBce4mvhfuQDTNOtI5eRDw4s
FHA6k9TmKfwFJSFdlgnCgcwC6B9x4ejNz7/XWM3SbP0tfpBgfspPze73FlaF2ICZGyr+t7BPfYw9
u00yAclPqGd/qBVySVV6lAdLptxz1sKALhQJCe30A84Eklh5a5b+AR6rvVJ2QTmMmdOW0V/s4UrR
9qIs37YA6S9sTO77zLtcu4GpuQ/yjjLS41aAC1R1gPPIOFeyujMlJBaE9m2m/cRLAHCjfq6rDTXN
HvxeML1kAF3svzJ6MELx0soTJyArIu4hCsz83AT/EKbRNRun4fZq3TCxVGEl0JkdeD6OGD8titgT
XgjF57vMYtcLhUbtVWC0epFphMtkiQhCNgHcuaI+BG71IEgj0dmhB6YMPV7F8YbUY4qpDcXPM8Gr
ypG+N9jYct7bb51OoxO9Rx0vOV4ypJe39ZbgkmMYkhPCLUyH8NGylllTCJfJ494B1c5fnr0G65Dv
FSq+xI6w+aS4wptfKpv6jrClmUloyieV6v3UzbnhZr0zKnyfrcdrYrxJRFYjEF9vC/QH5y0yo5DW
S/Ve+oGDz4K4E1UkiVVddrWLYFG3QrFJu4HfUuxoe//XVsXhGu1MltZNL7gO0LjrnYxo4H1eQhQO
J50BDeETlftTsbndekrvnLdXgEKeNUqQKSouWb3L68i3Vh9Wxzj05/7qP+9wNilQykLIx6IeFNQR
SGxZAOjKpvt6106NetrMc3dpxAg2gqzhYGfjEQJl005ptF4AiJcbmpEiDRx5rwJ9x6Pb3LTTQWb/
+Y1tubk4CngwPZXUDHq8MYaySLk656coFPJTlJASstOEAEtUlU+8x46MdJJWCPDlZItJ7pWzHZVY
TOH6lYOtcH6FzaGjZ7Mkgyk/EE2eTVZdivi8YKYfdIlXpdQkdHhH76n21vKo8vMTphcffJ8CgM7X
mx/ca2mSJXyZlrYH2cAPhNPoIZMcGtujc8lGaJFuraBQ1Cd1Hzle9eoiUmX1FA/L6RalD6jC/Reo
sa50XeDse/5WbXjNpAA26nKtzKMOWkMEMoatRRq5X4zumSP9/Q64HTAD+bFWqQ66M6EhzCfc0bUs
pzGapf/K7QnDdAeqlarq8wI7r90TlaEVSvltD3llDReLwk6xDhEuLXVmmMns/l6HZXTTuJE31Q9N
V+OptwD/KFunACS5XSiBhyj7HpY5t71zuUkznBY3J3LjCPJXCjaUqaC+ZXQp/7h0Vk/K1dsD0hAZ
/Tbl75CNmeN9NYIqLtBZWbExNhkQJvYPCQsydhC/YqWyuz6FRdHL/HlFalCiU/6qFXTdpe1GSheY
iNlBg+DD2qiOqcOKdNgr6X+XsMsMQtsMq/vysPAt4BGU+BYZJB8ED9Y2KZT9dbVXgHxVUe64uwSR
SvFKhPqisMBYsdVwQa83ABcu9piPn5jKfb1YZMYvsbmCg66Kcfx+Votz7LVhf8UihNo0C1cYX0R4
1v/6pqlqUF3wqNiygrJc45JgF1ZEonP5oe4G0xd57AKEhimhFkLvQwwzm1LGdolU7rwaYcljZeHw
YqTWERo2uA6/9tofQcGqbRSeF9CQTgzDOoCg2sVtrMdQZ8tbRmcjlc9vCdRL8MFJ1T+csR1HvvxL
/eZUme1UW7VxszI1BZUiem+pYs2D/6rVvKGE4gEsRyq/agIiIZN8bZSrNtXNqbcOMUZnwwfcrCeH
CRklkvI9TJiGUcLB+7JiDddDSmoasoXPtgRzNvJAhWvlL2rEZ81Mk/elQAnDBUkefcJbQg4W2fln
TlGDsLpUHGhFA6cq9YXXzq6zBicPVW/qOc9U24S3MhvJGNrIRNftukJXReKp7nYUI0+xRvuzJUx6
/x3lRZNsLbmsv8IhyhfeAZ22aJEXqnYyL6P1DII4LPh09NjGRhUnjh0JwOij2luMSAY+p86LewiD
yoe6x31+97LyXJPHJ/IS0IAjzRUkILkjW96Y/w7n9t3wxPY0mPe5kpFyXyVFSdesbD67/ng98qxY
Yq5mQPQgL8C3Nsn8TafADFaRYlV6HYoNIbnxmdmewA9YTq3/8LL+AeWjMfr/mTwlIFe8fWhFMalR
0r2SbuQGzmqtGp5CkGv9NWey3iuFtgOEcBzAD7c8yTt/AwssLMOtXBVmEdFfSiJL63gP+/qVv+RM
4fMRO8QGovaVXHx7lPncU1BMQfIeDkTcmiySrCx/h6CLD+sZpJy80O/E2w0Ff6vIlMOMTIxGF72k
kwyHfVSIcbmyVEWC5PUdCgc502RQnXiwW4Xfd7Ss7glF42Es1HRmsFfTusvHD0Nix1y7akQCCg48
MHb7Vyp1JKpBcdz76TH0v+Iyg2Eao/qovQbEe2Y7MlEKwFIIonrqvdoRx5SVd9ZLSXdis06MPllN
6flPxIR2haTcmj7qJh67qSEm1L0Ip9/IAEkz6NDH1I6SqxpNlF1Rm8Fi6FbY7wzdbDc+OoD66pZE
z0rm8Q1m6WKjSWNp8z0/5n17GCkVX5Og0X1xmjsEcC8vR2pw1fUZk2d/wNZnadZw+2yXM4YP3Toh
jmWgFavjNXFYi7r921TLJA01EoR2jhTGumMFqWZvXv2thjOoEUo4qVLl7dixyx6tEl/+vZqFNBIq
oTbCkOQpajkRZ2m2SdZDXWsXyahBSs3V4dQCrZNViPXtF02UILKkedvbt+3b/57wTxoPGOpZ6qFW
TVaLcakkPPLdBp8jTXV/nwjSKmvOIKzPog7PiFcWL+WclGIldARAQz3ftb2S6WVm1Aj1GuiIN5fE
vis4QBbxbD3PC95WGtWhQVlHRH7//boWlBZcjUmX2V1MqaE0PyAIzZCHLv/ovYky+KCqWrQhVvky
2ycXNwg7NiH1stuQrWp3cdilCoosv6iVZrDwgMs8Q9IGMX6C4Ae6f84jh+pyQ5q6fVnuZ1Hz2Ohg
6c0i2TcWyHOMwhgfx2PwH5wvgsbxnarnoGSSa9DvtbtJ9BBx3wfMpQV4OQGvneSRZymThNn3gWLn
uZeE+xowvC8uDQlNUdyDGaO1ld1hZhUWFLxMUt6Bc2uiYv01xplowGx+78HeqQtPwlX/oQIVrvdk
lz2Drgz3dxcxsXB8HrhjDFQeWX0Krh0+QNqalBTKUtPSrF4V9whtdWG7YK/LSmosodpZiOh5MA3q
gEQhw2rgiv+NsOnMI4BTqfxjVizl2o1lnji6OG5oatgGPSOR2M67E06m8spyCJiFLWFpFFBEf7Oy
rdfm17nSryMX+rUFLSInSIOXwqxaNm3FOkhgHttKnAN7y8h3ETNu6u9HO21ZJm/y/X37Toe/tWPv
dfG56NsUsy1rWuWSombvOmILc8KRH1bhjrMNCnXg7fr6LTXt/rheNNIsRvCKt7dmc2vq3orB0saF
teRySAU6qiKy9gZH5A9hhp/Yw9iPuUji2sdbP2oUdvv1J3nxYRIIGXThJbYHSjL/UKGrSZNa0IBF
bzhtIG9wMom0fQGtNw4yU7hA2YvlKQICJ0/I+AI2XbkmgnDd/I6nacZeBu2ZBl1oboodSNUkp+yu
uBxg2FLs4NqkZwPix/ZBddxfjZHXiefAMCl0va1zncNDnRSOFDVJ1prswwg+vIg5aRHiwhwgFvvJ
WL/ZD+hfYDRhDcX8XvCUiTmkw9HiO7MmL5+xYoidPJEjiOqz0plsaXLM18+suVPhMEPZIXzaEVhG
YlZ9bjiEatBq9mudqmm5i5wq06W/3rswzg8FKMKD4CzSQsQpWdUPytDIKZp2HhGg9HMPiGZgKc1t
W0q2216bQ7GHFgvo1qGX5JubJMVefVDlSgS8I/kmYi6OEj3W79rIddI+avjTcXh8IxpFFn1jBMno
LBzHgQ1p+y7lbGBiuKq4D6Jqa62t1W/Zsfrpd778gKCHCwHr7ruA/sWXwuLVN3lmlSya8C8JJg7w
E8V2cunBLE/AgHASJuP98rI/cVI1l18/ZltUc+A8zbrXU6SSUMUPkkBWiaXrmW/7YqWn/sPiO8X8
XC/KKP+lhgPVT7Bf7cm78t3nTOGm6POWySJzzuI5cyy6TOQIXtxbp1Eik7psF7NKIxMZrN5gd062
KZ/9IkVJTUc9i+gD1Js7DAQNeslndOxMu3pQ9SqQoIclANbKmNmyUsj2wmH62HLmB6ZXVaOfYkoc
IBZhlKgrb6oDPJFyKzt95s/1NuAlv0Em78yjT7njkLAur3a5PQn4Gm9FbXs36TCrx6NDHmYc8EG/
MrGTdAJN+sXaVQnc9PTlx9bcjC2tSWFQjAlRxAovvMXdBtHRotkG4TnfDSkdAPYhR2idnou02W4+
05SQiDXAsPHWQ/v7dXGRFM8WIAoGp8fsz4BPK86woZBjEkCXrQgKqmFtrthi2iKUu5/ukwF57C6E
nSh9v5m55gjc8LBsfwju0NHGvonaGOQ4KX5Vfg4/NEnKpE/LnUtfxqlxkiVYCextbenfrGLkE5b2
6n+aQMYGwA0HilGr4DGLXFbZ/SbdwYAtxY9Nu+n4Awie47XA22TaNWwUvfnMIV8UI8VQtYsiVF0W
2URxA+nwv++gKozID3D46cz1Js/eHCw7dLcZPCZkYIV2J8Z3T7GPsplje1l+XcY00Qa7D7fPoyfp
irBSW8bSxe1irci+s6d6q5t1O5rXr/uBsD89UwgYEH6ZRbphiBAQHEn9i937A3f2q1tEgPV2wFMD
vXJwdTP3Q1PPh7Q952EXUs0RIXJQB24i5u9zDD5y9lt9grHgIxYmvICUYjjQ3c2AiGkUHSfkv+mR
xjnCTk/30m5cCNuJgpzpgRtqVH5TMATUUKuzRRVCSYgp5c+srJX2irossEbybbuxjGOmL6uiXbwb
7zGkAx5Km/2ZXUP2/CmzMq8X1JNen3GKOxbUfjMHlkpeg2WHyg8ax6EiC4hmDciq/GmbEuvzsyeu
oEe87K9ro47eMb5KI4Qo1wQYYbK0T/fL8UEzpz2Fw7DXmd9E6tNIG3GgQ51Zizty/4jUSJA95AzY
fo7VXB/hjNIkY6CGBqRqrZUHr7bYDmuuqD/EVZr+GL8yOV+P9rroQKdGdD3mZmCyaTyPW6q4+oxD
WoZhnhbO2VUPFgzFIwk6LivAi1wNalJW90jTKKL8DTpJXEYM2SPJ0lX8PrYBEkyrQVUcxJ/bsDCG
Oi9LK0qLeObIo+MAkg2ADZH+0dQsIFupW6oY8A5BXAVK7Nbs279i5WJPuNAUsEH0ynMRV7e4RMt7
NavrEOt7+tDLP9Q7G0owD6QxiiJWZOrq7fNHp6z6z4Up5f7UiMRse2aql/XfMnlubG2vyR63or0J
meh+uMS2ulFGgPt196+HjKUeq+MQM00yes0/qjjxbiLyEwE5wikXHkNTeF3mm5FxQt/qBL8r2s94
AzQx4v5YwDfgB0+E1MHLyh1ZBud0FESGg7tBaz4YSjXQ0TH3x5O7QUESWTyIetU69wlgBgRJxcPO
rnme3NOlTkJBCcr59OR6a+vxrgiYm0h6Y/BIR5/fE++cfZN/oafwxGDkH7fPwxsQLmTeebRAcZHx
COr2F1nJa2bl5Psm/az1mZOkrs5InL9h+v0zgt1uLoKuS2EHIXP0y2GFp7XDN9oMsf2jdIimrPdn
WbFExeT8QzXd7RGS1Xg1xMaN+IO/XshtfWT7ZrDKLG80i5p/x4npxWh5DoDrbtdJVwLkZtVVAlMA
PvO9Ntg19oQHEk4nwHpiPsiwDQOLr5C06GpsCTNTzWfe+8l+YaSbpRI9HWA78rfc7mL5imQBuyr5
LCOSx5bjoXmyX5X18lfrpSnfQdfRHLJVf85Ot12y/5rm7mC6Nxk7G/TPRtTFMg5UMDhPo76US01v
abdy50llt+RplFFbL8aj1EaIXyoj+f9C0O/5VBwbsl1ClU9t+4AFjxBC6CKo9bNR7MfK4lXG0/l+
BrAIkhryQtBdSOKfjXhgJmWT85HFskZ73ccJOrWlkvYu/5yMgTgtwVDnoGr1+A0Gk45wrYVhzMPV
xilqHBIE8Bkx1kb18c4RLBvp+oZwz7SFscDn2F8bUEh+j2p1Qd5792RWKtVBFi94ZmnJQ7NtZn2m
+VKv9zZeS91aR/dzqGBNPWVur3f+N2uelz7lWPfQnOBLf2pMDm/2CoA6/fkWyIM+/dlNc7pOu9B6
VH5vJhDFR6KiTfzOtRv1C01cLhdW/X4Xuz2PV1AQJg5VoUSayNUccbz3vqyDijLkreAcvvzW+gsC
cW+IEmAsocidHrBwSDdWOwby4fovCHGqu7xuVlI+K+7vSKW391dtN70Ag6nkzQaCxDghdp1X4LuD
NVtzoRiVR1Hygxow/CtD+AToTUI1Mxvtst1hV0Cb+Glzp/oaFmEQYuzAxygTFFNwMQkAKCaHN99o
nl1Prg+uhINa50s7BvzkDlV3I6oRf1syJjaMeLyaUPnVWGjcKnrcD+FI/GxHaPOYuUjhHIXcCMMK
qP3mQNl97j1tpCIxwKCeMDGXsu/JEJMNyfWL/VTx9xAUDvwB8H2KJvoicryJR/wh9WKO02IcgQ6l
jNYzDStMXsqC4K7MOuqvDQpVgRbdCwBcsjTU005KbBMjejTp/XzqVgwWTbV8fEDp3iybw1ZA5sBy
pySLqSuQ+Qna/GXIn1Yim5EhrREmYGKWW6T3VCzBxkaVvCd8/jCSpvpDwsTeP0ahARPqUdlKVKIU
bAOv7DBobgiSqtmpzDPapuCM3ZDYPYvyJ+FAHwcmZaxlH+4rscM7hkZceNB89semrO79WjaGh8z1
Kn9/8mJ/Rb31hhnYEVdQJ2xDGpCNby3ivbgTjZNVeLT7/S9pLak4kbIxYcY6nmxRn4/C/r6jzCzU
q+XcR0f/YUspoHnv8uCRl+32HakqdK+RPOQpOwYdLTAqHHqZcmL5b4TcW+O9AyWNhEdz+GYDyztv
K319vK1c3HffU/w4cKEroWSylPHwVTxmJsA293VqVHxKEigqpdhmCEGZpbBFZONHcSPyOCjZGRV9
bffKjrqOH9QuvOFjSeHNArnXZ3BeSEc2cI1ALJWr9QqF9qm3MOseOrGL/BKpEHLIC0TIwR9P3P7R
8p7JvwB09tzkWuID4CHJkYW19JX+FxKuO7L8j00bNQER9AnndbatbwkRiWq736JsjsBnMHEGKA4M
uYR4qO9lvlVxhCkoHQp6g+kFhPmeIWVyxY3uGIUgXYGftBqZaXP4Uxrd0vAGpPSMArUAf2nz2pKq
B67B5HLDAm6/C594pKTitosFjdEKAJ99Hqf9xWxN9WdSrLBAAVXkgUItNgFxXhd+DwlVWlGIKZFs
d/b/RCnkfRm9nq91QMD8RJ2K69omPJTM9S1rNotHlXtxqo8ymQkkPf1WUjGJvNLwRtUqX+opHpfH
4KgeZ6QPjnYmSrYQtvfFCviu99gGvh6KO0DFgWFCHXU97/TcMNysamC4HhgkxtrHsNZlKJLs3Isu
Oea8+CfeklYFW1Q4T+AOOOi9+/fY7JvZBqyy3avpOdytcCknashBhp/a6vOJxEbVtRZEISuRsict
dE/ISosDHzpDs2+aB1p/extCOA2WdM1YMz9aMqqYnbVsTO1XqoHp3qty/MJmH09DXy1goJUascni
ucmbErWtHQkcM7+pFRYabZp5r+YZKr/lmSPxpMk43N4an/uGwJPWKbuzdke6v512ePS0Sg/lc8E5
Qq5eIY7fiWl/noqOZRhmT01h/5ThwVE6TizMhoj6e1GfryDaua1AouujK97986UF5lZ4d9733X4M
B6escQs7X3ZFjMvnTkckI+yvIpAgrx3wFGj8grDIs2ha8fecE8jfHLqzJtJHTQsg0lNVimbSuxaj
5l34aiYMTC4RQhr/G5eKJhztA3Gllt8tPOJJM43Z+lNQ8Qtj9+RQ8hoNsk4igEUGd5bgkey6qvtw
yCBz5aAmeZfortylin5mVLDWAbDY4F1A75diCLpYMn3IWhsm5SF97qDyc6E2HpjFxqd24Buupx6q
I0nP5D35kUrrM4pW/kznf8WPfklICnjU+eJvxCkHhzweAMrZRw+9OF0LYXUB+RCfvsP/A8cx6+98
uddURQL6IcMX2Fa8WnvONOjXqbOCzWtDk84if2oIUV13zHICzN85OuHq5zPsQmP1EqUZEEvqljXy
lQ84YTUT+KJsjUOGRJ7nUf1ebqsDOj5Imv/6l6esOJOnkzmjkvFJrn1VHBCwrkMvRW3oCK8YQ1+o
aUn3WmPx4E9s6vgCGMTHxk/Q+BXjp/C+tyeDsH8ur0TYxg44LM81IAc53Xu+YuupR7Akq/PNOJ6I
EUtkjbU4mIGAyq7biOBieog4WkbX74FR+1qflLnJ4p9BCQNLMH4TO9vimKngKAy18+ECIgQEB1jm
VXWJJi6wf+QHx5kFmnH4sGSnn29PXnf9HsCT1c24ckAWn+t4WYG4lwqYs5Sv8dSSGQhOAlGhO6N0
pl5pXWhvX5bsF+kVoV4b5ogPB72153AyWsUc8lQeWID6E3ZR52PkYxQODKVhpNLTQ2x2p8BpagDo
xgEPsSk5qa0ZHDDiBt41jNZ45hq+sb/79RUDbfcGUhpOjXLmnziEbcXXCBDLY3BnVEB+0xXKdwY1
ye9lBN1yBurGHoScqNZtlPsSaHr30ygMi8D/I8FOOs1gwppFszqZbXmeZRlRxJoGWNccOHspQvvJ
X2D40Zgw3nYJdaD69kXSD/wq6Ri5Awr1FGY/jOWkqfxK0fl+W+x2h85peWhvF+PKIs0ojRaEEhVr
/u2PuDTA0FwKiHMhBLCby08q903wxfixtsrH6ILICL0B6mroGfnZwvffVndwKosXLfXnJMjYANwk
ivHNZZm938P1YyMnos8QKrdn11rV08K+KrLhSF5+Ug8L40vGgkc5dNV/pFJIDig4POvIMGJKXt0m
efanhI+b016RxZKaew0pbgMaPjGNxY883ODEHXWbgTpMWf9ZFkft1cSrbQ+OpXquIn40BeWvZWpN
6y198j8fKQEuhkTh78dP5lNwH59j+sUuD4Lt+PD2jx3NTa+WzKQlyLy0l9gE0xB1K3cuheucLOzu
tVwbVoOXGixrIHKZny1UU8iF5otSSL1A7ETnZ28JRnx7hSdOgQZvY3wpadWcvQ/5QU8ulh0Yb6Jf
nG/4jDeM7NA5jMYYBlO2jrWtkiU717n5c+dQekRI5fq58aRkk+6CM14M6F6QsLTACdME1JhMnG61
qJ79c6zmY4aw4LytAWFZHnUKh+0mF8grx9EpNrZuvaAbRVh+PTwWN9LLP5n4ON1elWo8CwS41PGZ
+fFy9m2Ox/k7AYlacAZu6lgi7yBsU64HrUrhuZJ0Slymsf2W3ICCy9y6DMMFj7rUVhjSewvqgQjc
8ua+d8TPVb5TcmOqh3U+JGn0jyOY0HuqFvV/NwuxEC3Ab7caU1ogApvHBqXLYYRtL19rzzorMKmD
qZHT7F8LBhG78I+PU7/tr+guxAtnngOEwaeRTGgU1h+mVlGZFElnlbiSbbDtGuAUyTuKoFmJLun7
I5AEREDD7Kpl8y/hJIbk8URVzWeuj3qE7s8qgDall+trunUX/KdhC+xCXPzK7d0iVK56dttfLF8y
6B4TsdcOz3pyaJ5euWkMgk8DVLmoeOdczcdP0uSs5GcfcYUaqm39NeEBOkVsB/0UIwuAm3YEnOUP
FBlfIghYTKxGCkan7blfjdDT/kk27O2m+q3fZOITUVzB5FKiypRr757rOpfg3NNB6k4RWH3qq3AQ
dQPQ8wBdtvvkL6Fatg0xlkiS3ThLgOwXOjS4gShh1eUAi8J3VAzV/2WJHZ0LG5YVpquXSccREmVE
BxpBbU6wMG+VyIW2GNjSDndmhnsxOyFhJ3Q9ryWhPUAoqF4pkqQk4mbwoPmFnBRND9g1JrXNIh0F
cxhlZ7jekk1baVgctMdLxRrbQXPIQq4Ha+pHi3QNEL4QLrwdk9noIpXs7ve+RlNenZFpnBHfl81X
GojrvNDhtROllwIvtVclj78hROwcJrhAels9rD3q1fuPoSE3BosGCQtGbwKVHWydgCL8PSJoVFvT
DqlU4qvg/jmkUdySIOB978Kpc6xcJV6Ju/WQF/5pOUDuT5s3XKn1UosnpxIZoP/6/F6nciONcF/x
kB+4g8lECXO6qkzsN8x/0ahPq+UsfXcPqmUcvzS+ptkFYQQtjIECItS0/IINeBy8Rbsl/OvhRUDp
l3coxT26714xIFdPKIq2OEbsEEFwFC66xThfQkVO/ENKqD3dL3YRquuCuDcCMbZYeWZ9049X+1aD
MDCmWQMWhBe4pIBkwxOjYgPqi+hsCvbiRJTFrTA0xsNiVyiGGu4+C7YoRWa3qmwDtvwc7KDddwCX
UAJ0tfYwhIbKZuAZ0q5aq/6mIo+577yF56uqSaFS/CKgP0eFEyP1Knka7q5e/CGcwmO5Sv7E9GvN
j+T5CVwPcRPY8YTqH5m4i2fNwunEQQgGq06uBKkQYm09i63Np5ejcDrFjW+cVOA35I4jU7D1SUQ2
zI4Z9WQxgNoJOnNp8hFDQh5e949wRTuUVg33kyzpnFsOL4rTVUPFfOO5byRI6FuXB76PxRQKHQAX
4UM3tlNj89Z8/eBI0FSyQLcEYmV90qgrWiC1jR7IUlezzZkHlHbJpEbximNtnbifXyaraW2iXN8v
IOUQt1IrBqBnS6FBcHnIaXewFSekPho9B1W/4DML78m1VAAnATSPkl6niCXhKo2z0SDWrYxam1WM
qUGlDPXvW+u4b7xD9WM4v/0bVB3DZKvov6lKFB4tUC1odU42zm8KP28cVieGgB9+tAbnPK9aGtNO
XnLdtbOIfb41xH1VB6wi5l8D4+ieIgYMkz4xBEH6/uC7HhvgBlWuW9/gmD2Q5p5GbsmjDXA5XMu0
naaoZGUUGHNLxII1oifWnZFlMh0Uli0TobJCH9dM9b1zWZXVtrHiyhdQi9hEJcXdWbvLUvxoIAry
FKunrwWc/ksiMQCLzUYTRcyI64eQs8/MINJ4tyz4G+x9VOyYb+Da/8iHDCgu71SWc914psMwxOaf
7wzXbwpEbNRt/LXVs81Wjmg06D1Lk+Oi2nV/HSLX58keqPdNe3I9fIRAVez0b0m4JhQJPu5hQaFk
THiqDfQJ93uOAmgPCnV//oGJclVgnzhNJuGET97jF4q+peTB134RypvSOMySgzPziFXWXTOd9+FM
E9TEm2mt0pf7eUd1Qoiw2MTgomxStOuZtY5mfq4prgSwMR2pVNH9cipOWPT8fwszBVw9toczF1Ur
YwbgPY3wy8pXt6Smzd8XGRgFmGv+35ySISrLT7nWNFhGCTPAQsDVo6FxlHjIFSqg1Ka99/0eVWjZ
446R853Xz3cRVbPbXJGIm8dn6tcIvs1f0pdqLDbuw2Uj6OTpaTcQQ4rjPjUd1v2RV5x68rVhSyKQ
GQCuTJh1vARIBtMd32FgBpRv/iWMt5fYizKtJ5bA56HbiBVhITfePQWkMg49Pk8S1bianGOYkfEB
XiVjuX02/pLKC5V+uMJ0o7rgaLtf5aVwnLHQd0GCAACnFgienPaDGNdPm6GLGjp1nq8ZG82R4vbr
rya46wWrxnnqa9+o2jQDfmld6d+LY7i0kgj2gruvBEX7WxKrmpu8Lrk5Jrg+f47bpf5z3KC4x3kI
n4vNt/VC7h+7i8q6V0v4vXHyVZiSchkhDgTwgh6ZfKuNpL6GqJLd4WHmlvWVLJauX2hbhasnIIfz
vY9tAW/KnKe5In9Eu6EbMuPQKYK7o6KNqtpXwzZSRlsm9U5h+DEwXQ46UYxgTUdrZLeOy6eXZ63z
Z3R2RDJvRDj469Bv/+NrhNBSX2laOsHmGku4M/6NvhjY5rKJ5IIPSy8ErMYA6LXOaYd+sl3eZBbD
aDnPldCwnJCwNydK3fVqGcU3B0eGMStD91WI4s3ccgZNizSU8nDkdPsKCcUN72qf+amzRt9UW3ao
yZFR/snR17qwCyUN0t1GTEBqoODLg2W9YyXP7WW5t8mnhU+YBpDYET65HNvfn9Vq5gq6FO/8CM12
SIiuYTMxHM4QLtYWIl5EDR0z0mfXDQp8xqeaLwmXVxkaVonQ11iBcgXh/dtw9D2eCN962o43mYES
IKzmBTQDUAJiuxjRfhuys/RpgSNfOtl6AOcw9dvwfl42mPO+wlgZLYOVAVaBVhL2cTuSIShVKq2F
dVrceDltjJAVIF8JtKqvqFhKfbovYHWXU+Z/NNzDuXKYqWcPWQV79qoFl8FuR/sjLfK6QdGcHkd0
3EsPZWD9E0gUPjAc8z8PrDBM+eleoVQso16IkiIbXVIpC3z3dBDGH3VOrjDjKBpkRmLwu2P9bSrv
+LDMgVt2k7E6KI+RzCm3XJgBredr4MnQit9jGz0mtmlWlzYcE8s7a3nQANB7g416WkLL6S74JYKd
/nwESFqPMUGuGpCj7bvx7B1SWA2qr/s2SVre4drAuyqOJ43ddzrtD5c0lJDEQyRNrE2v36kWDzY8
cDxQbzvCDrMO7IMumNC7vtmUciLs3R2sqYK8yS0xE2b+YqKN7jadTjNo4BM39gT+KjczgtMMgQPj
xbZsaGsSejWQVxt00Ne62TCfbRT8ZfM+H8mIyVZDUVHQ+ATZ46D7I9pLkSRRrxcFHIBBWvJbu+tT
EtDw80+DkBQusVg304K5v7sCndyKV+eQ8m9/vN5ODiULYKcOT6CWPsypeebJUq0/mv1F1lkDfw35
odzyrQxLeqwYIjw1NYpa1qplzW1ziTBQKx1Bfp0JkwPO2ci1NTVP2mFYaukVpHCLsxyCANUa0Zb9
PKEWKr0+DnyWs4USpWmznlHKsNXBoeF1GOkhEma7hpRFC9SH1R/8fYvwMSEZ6fBXmG0j7jqHkp3x
/wnWtmmL/bUIlSeVw2Wzx4WZzS9qJYcVoaRhBRxmRK4ETK8c3tqd6cec0jCH9nCF/8Of13f7Sigh
2vW4VKuU8W4hoMfQSsE16wAawOw+4PbFT4jDVMxCaVUf9r03p4w+UTCcxBEc+7YGVc+t9/NyXe/v
1O3xoDq2U8GtgCGxPNEFHABrdMJoPrujpEP2lJUKsH4A6f7J53nDh1Bre347Qcwzr+O9A0asot3E
IUy4CYlrqu05WmbaTlrArsLzKahB2uMa0uVsFen99htm8NoR/lFY8jlYzT04w45T2l35qapLniks
WCgtaeQBa5oKTOq6vhlunDZJ/FCC9JkfV8n/XUkyNv7Ey50Iu1xeQWZ98k7xuqwyw/XVPUfm7fYq
kzv8ZD9par9FrbQefUSKfd0o6m/t1oLn0FKoEzg83JKOrtmI01Ggnxg58Rtd+akQljxSxOQ2OkUh
8qjXo6na41IKv23kXbmfG1Bz3xyilQRUAiw2u8e6Z0YIIMLujfVGJDGy00/a1mGzyCdjpBSmH3CR
wYCxF1ylR44yPFugd1RUz2RH2sSytxGYQg156Gz+hJiGKc1TPQkUlY3S2iKjWCbmwyowaOt1yTG4
xkq1UtYRk8YLMAUJTc9yiDMg/ePn4w0H73D7rKPJ3IJUPPHskubbbqfJ6RjvCHcdiHZRe4jslgVU
1yg4ZjOzqrYhu6y51be6Xz3hTKcEhNHWyxGUMv83jvgk0fcMmz/BWsMYRXHyv+7EN76Y0JN/aNb5
1IKxaKwnivnmKR9acwj7WKfUkJK7sCt/ef3IzhwenBUJ4wU3qNvvf2rwrMsAfpPzDy8YGXBhrqUW
ET2S2bHFRLF0YdZLKXuvVQH/Mqhj0oofpWUAAIxBF+JQ/Gv/M+/gAlBx4c4aOADi6kQ8tOFZNrpF
jLYrp0r1HqBWIcB+gHNY9vhTAaXTXkaQ6YhxGYxZrrMbZFTqbJwFnK7o5G/D6t0Q8f4eIRaHugYv
KcXj38tLh6pxa4qPsl8SLOf+ikzx+QCfWUwAprcfBcua7oS+Jo430uFLNVi3q8rkyL61X42SCNVK
kxdHAe5ipndQTrIqNQ0vhm73xFj99VhPiB9i5EFslWIaLXQeFpgR11VC+pNVsTlsoH1utdkL9Feu
clcNLOHxXgxhoi2eFuUkRc+syErXtB4z+EfJXbKWnlaNd3obHKsiKRyOxkwKdi+XaFWpdNBgF8Oq
vKi+F8SJJF/fWFQ6sGaV8arSKV0A1hdLa3+mV/vVPGkFUxwgyGnjKlQsEzzF2PoODRfBpEDW9Bzz
InO4jMuadCxEwf+mD+7gTL580TIuj8dCQZXDxuC0ytJNeCDGGA7+1YpagUsx4S0mEY6e+H+66OVB
ocV0uhDMsuRKd9Jmesau2iVK6PL+c2BcYecl2AB0c7cAwjLiPAIZicKc5GuHNspYMr9hJN6WH2Th
xwx4+46weeQaQ2nGACgoB/oZqrOqAqe0cKEg1CPnbyG1c7OmpnBk9ggSbHK37pl9BzMtthg4gwWp
DvqVhRWdVf/g5S9xyIgfCiMy83/63vCXcpAACH17MAZthZ1KCENzaFfiTOH9V+wma3KddLXx20Zo
iNNjkrYAG7t3VYMLDfgwCYlTzpj4d+0nmw890bo+ahcyvpDBxP1uejOol31P5vMB8RlsItrPTL4G
cxsu0VrZmRawYiHdyM+5dj9TGQX4NJUWceHELVHYuJOBN/Tchjklbul8q8pdrK8bpYfm89sIOkuK
IszRDHOMGuGl+9BdFbxtuAhX1QuDrMpcsoHzUT2/hWTVtk4eL4bX2uo9LOjdYj20QpTdQziXByP5
BPMyTgI0yKbr74cf8USeAWMRT5KaVYEx5zKZv7zXAd7V8PHb0rX1hRrFn/3xQ5S1BivLXveizxUg
56Oa+H+g3xsnZmj8/u8NFgVL01cFuMxSRW3WQmS7I5YV3E37vq+SNUip+wfXj/MJnpQscGNJVoXG
nd2iygglPNI4bhiw4K5pVV4n6hjF1ufw42y02h67sgo+vvtGCuSI8ETd1DQ7CVJ14OL2Zfv4ByZW
3bD7wfjaDqddwA4JhNSeXdVzjNdQGd46sQuvxfobGZanyhvLAGje3ET4ny0umUl4mi4U3UwIaSKN
krsFWOWMC+brAoj+hDbLTUT4eKy15VZuMZNXPM8Yffy4j7rpxrg44cplQg/PAo3KN3LHjIpaPcJx
L9JkZ2WvTRszmW0rC/IbXKG1L+RxGn9rNZHbFW2vS3tDJkPOwdz7PGRWU0iH7puomrJ/+cAWnFFW
Pn+wsOuzSpPLoUiHoN7LNkEfg3EebzNg1DPRI5MNy/bar0V2R4zoY6Oiy2vB+/0WTl4fVVGdzewn
AX+YAxx3a5vP/xu3UHqve+q6Jp4KOiWbs2nvykJ4jglNrrs50vZcdiPiDu2JmN+KO+sE1nildTOU
Ii2m+Mw9WSknYbJsI903apSBmOgDswUw0oFPS9zPuFD7VExIg/OeiQ4Lk63XebvZj6eN2BxecOc0
AIHweZYs4ebzJNXqQvSNOmuhPIMkL8ZzhprZ4QfqfCBjR/6z2MqNn5Znd5ILaQV8sKCZdwxMvM6f
yr2oVqOgkwY+FTn3hcPZcp0FT3GDiQMjm023/NhAo32LIkZ5OnsPOBunIOawg200W40EWXR+OBnt
oOVg7iET4VA2oBPNHANRFgRbp3tMCCJrtu39hG3Nn5U2oczYD9A/2vD1+SYVHpWBE5Mn9O2ddxbM
Q3hDenOW9PndgYGuc5CzjDeHmDj/PqRgD0h/ECfSNPLkOPRnCvleyEN2jK8BeL0eJqZsxnY1AJE0
47U6Iwwa6IWMWyCHGkEoKmsExT+shG/tYj2n+qkVpzSikwygmMg7pyQIcK7vgmbakSB9RgsqmioA
9cxeX47rZdYWiNTLpyDjx+tn4IVJo4aU3/uN70Y6T/tdZ4oB0AlMg+HVF6Orvxpo10hMPtAv1WCz
1tKpF/PjOWxYSt6K9PlvzKVoOh+HDe2dG9fj2quXqX9PIe2/kvzTixB1E4m3ZRe55/FxXPWm5Sz8
FUgNIlru67P3NMI0UwqOGwmEsZKPfI1kUQCFxwEJr/YsWw/45dpWCOeqzFQzr2HJdgF+3SRXX36L
Th5DuVnGMmFj3Tu5gMQ/F02N1bxca3NV3lNug/JhxebvMfae4CnNahIgf1HZkbEq6YF1fiN3lWgL
oODZtRpNTKgQC50QD+Pqbl1bpLGBqbCB7trbaNm/jUpEfhckC8wA581LVoEk8eGcLjb0ZyVPjODs
45wep4DG8B8q2SY3lOBojE3WK/gswbZFrc1Z6xZNnbiRAwIEeXEDkhZSD6rCoAzXcXh9ZeC8B/il
JSE+HKIfOrliXWkeZfLzlw7vQl1jxRlvFb9mZvWeAJGc/SD/ri+0fOZwXx9zGtI8GzNmOzl9rOWo
oscoCuKkroVQUBbHmoWTpP1xq18UcaK26N4QcuMoSWy6Q9MMWGdPf1R2nNClaK+BmLu0vs2LnRB6
piyraAZC3tpXc+ucsPZssBNGlUGz7o9Uek/IhGCGrmCjyHZsf0fRzs4MPGtQGPlbOTvrBthrnUng
eQVkSHrh4LV6F/2MTI8MmyEm2ZtpNOVMvsR3+m4gtGTh+Fz/QcO1RDI4Cj1b7v1MLlxtd2fG31bT
xaEF/EQbZFw12+sMvwvS6uHZVmlcEhq09AQeyBgi5dwg7mJ1rGzOrKaHD4qDOT8QqaoGff2Svp3/
Je+nH5rFTSzRar4vGqWWiTW2RGyTuuaDnr1Gd9Aaq2MfaVkhVc4Y0MJoPRXmLUg8x++3dUAAJ3v3
oa3XLy32GYIUXz8MMcIjL/KYM7syTSj1hwg7nl7jB+eubYi2Xbdi5feFeIZuojYvQ/n/r1u/X82I
1+S8pwQVrhVQWc4xm+eixw1as9ECu8YPIXqF+J0hvxAsA84AvsjAYYyrKZuR7yd2aHsOSJQpr2zR
n8z495k56qCpE5p7/r2z4JIROzx5zEPiDBJ7j/7exCeY6v5gxhqflv6p8LW935xmMIhoD6Kd4Erj
D4B/mjlc1lGDaU2UjVVhbmSnIFdvkOGYfriNweGr74mgTv6nHJeUIaGlwcA3sRGvAy3fFR4rV02G
bDXu99MtTkCkNWoO+tMdnBcq5hL2KqEeifizknDXAGECBA2lkCDG/HxmRQwMWh/8gENdwO+zPts2
4qJrdyOil8J91mVGa3WqQAvOq81sYRFmbIVqIBz9aoPxEJrco6QlizaTVH9fwunULwth6SPe+nep
nSUV4Jy5vSE9gsbqaJuMpXETZjJkT4g61hyhDcDqkg9zUtUvPSZgAEYXsH8N6/JHnTderWsA1JD3
f0ATEJGumE5byxs/msyP6NATBDaOSvl5aoFTw3ifdPdEn5MmiM/UHBGDcUFHw7xe3vGSzHt3oduB
Few1Y4u7lZPu876n/6eK9HMQRoZtxCuvvxr87AWUqBqklEydThtwJxWN4VuWh4+PCiGycu6nsvsz
Lb9jN94cqvn6gPh6Sup2womqFcswbdl1xzHbp2b4axBewGy8fXlfNCemf5+RqDPHEkznUjU3Ufwd
qK8iYnsQ8K5WfV8ZzqPUIwkUFcqRUeF8ICi9UwoVbOmR/vJaqWUC0hyPl2RoFu+zpAXmnx30SPlu
4CJu3q2My8uOyVoA2MK2dr53JJJp+SGg8napf/Y72q9qfePDtRl/z7pTQEzNSNp0lisJ+JRqB+Ud
18r4zZmkd9MFSZGqCxARruk81mufBOHR1vv6fmuPx/sQ/GKCnXrfiPkCppMfMqvCm+oioYIJUYS0
/K6zk/0McvHnvItaCqFRo6T7Lz3Xw/+yh0w6NBzkYj688uljTeGTkpmFwjR1X7F4w+OrGRdv88wb
NvfbrzrI6YaBxalFYj6KHbrb5jtPiqxk6BuiLGJMK+7xGENK3KX3N2swmYZbZRHKDamP+Oa0AQ6Q
8pUfE8n0NB6knnJpHORKuXFqRLzzu0Mi+W5O3jfc5ZU0iDnoFmKHE4WT4BbzK2U7zUv5FPHie5TQ
70sTKkcxhm5v2qwMhHZjLOZ1ndgMm6S9KaFKTdq0sVVJcKxanM1zTQ52Vi34Mi+n88Fvb2lruV0b
FmW2soBifq5+uKa3h9RutDKbPdu7+AMSw1bS027h2E6GPm8w5zyhWEznX9cUy4kEKYnmRJXs38EF
/BYfROutruZtsSHE1bVEEn9kIgrk6wSZxjiPHzJyxpAEJEzVZUi7fUgkGmuBreNx7dFs87Cm07KI
Dr49wCNdxFBsjvuFpG4B3gXZUUkS+lnWU004KHjNSf/GGbL3HYc9EmBdPU3ChfTyrEfdqY5wOVzU
0ggyBR/4M4i/IHdm37SxXCG9GbT+6GO3DBw0DInktnw7CXBgxh+H2Je37E3rWfJ0W5p6Gl6O6+64
zWev376xu8I6BO6/rLk3VaQ7hTzkfhJDy1kcSZHCpi6Tih47e4tn8kS6H8y2QeCegKpLC1ar/Qhb
eSb6wx7dkKqEqfCJzXmqimB/C7j1Bh8QBn3DlxOE55tw1Tvj+bBjNiYsGWLsKWtVgRFlJpjV8seH
eq6FDFL3OjfD4ngSQ87CteE1S193uHk2nJTjUXGFEVO+Coo6htMp628BaInXyxhvy0trbTd7k1l2
9e5K4UQuA6ls/QJOZTZHkD69VVKm5CvYOtA/W8koiZkdUA3fh0Wl8owokeVCPtugDtGDc6Ye83vH
Y2YsuMWNnCGmLhIhm4gEp0v/FEalcYMo7dcep+qyXb3utphy/dDv3Ev7ssYiCTvLkIqFOg/nF2DJ
6C/vg+iXRjVS15Jhq01D/rRwyEH399u1id/u5jsENg99dEVyheNNbKKQPcSnQdNssgDjdS29rJCU
tl4V9gUM5oOy1HwNqVCCVrsrn+nC9JW7BtRU46/kKllt/fRDw+Qa1TytRxuz1pjuqM8pwbGXFwsf
90IyYTz+Mm9wBsU35KHf4ZSb+InBR+xJR3Gey/bw5Sm5S0eaXkas2sHYGKrHmAcg8HC2EF0mMFNz
0AzbC28yGMNZM5y5HHIDmwzFZt1lEYyKOXbvIk1WnrWYhH31NSWn2OzVKxub0So8/GH3foK6vYmI
tKX1sTiMvCaOpY5rkLAy1j2su4f7WNbE7aiJCBXahLHMWEeyyvR3PrTXca4puhfTG5W5dlJktnY/
gXKzxoFnzFGspGzmPUCoy6gTgLef3WP6vHKjw9SIN8h1dcT/C7u658fyVzWS2OW102p7oIVfruKM
PydkA2oIPe9KB+aZAcXLyVy3lRttb6fm9A09dchzvzCQGpPgkuvON6bCmyVpxokL8+hP0+FQQI50
Yuy3qEBV/kNfXmvABjRPj8QW67ThsB0doW0kQHX6+HcOjjoPieiyiH+1BRVeWGwOCqkqjy8tMEnx
oVDfVoyPw4SX5DexjjOArlNMReWNDO4MhTjvghBIqTzzhBCPup0pNrVv3PksHWq9BZL6jYndLAZd
xjGXzTuV4hIFgKjj6qfRNaGNnxEnp8MiYmy/3y7gJcqLe8zE8Zvj4X8Env5Kqg0QHLTVSc6WF64V
sNzH9YGDpX9s9lemAxFH5NvwL5vFI7ClI1vNu+cs60/PuLXXrLl3sLqlIryRx/jkZYDbL76cjLxf
tKL4A/4cx0X5pKbQQK1VPwSknza8IlxhoBgkGMkKYtc1xThppYx1IKa4VpiTJ1SJ4OWEdSXqtPyt
icX9NBJ739MksVF6KA12PYHvIB5dbJH/vWsFpLhwuOPXn5MwQIHZ1iRpk6iUBTMuoVDgQ1KYRo+9
7D5/Fo57w9SirVS8CCuL9X6iVZuZhtmhp8YmhK5WORn2nrUVs8gbWX/WRCMyqfg+7MUyJC9r/GU2
ElJZqG1Pe7Ab66Dhb3l99mfjDrom9EeazGH+ugEDT33gqfpCAFOIikcCbzM8LboVZq6AZLhI8iPI
M0VluiZhve49CVnsUP9yEuBQFlkP61BcjIb86iYZxEAmdNkc23JNMeAPKQWY0QvF4tHn87eOUuzd
KEdp2g2LR4Dp1uzqurBRUW5syMIQ+D+pDjkHu2PTMCqYrFA/0N8sUl5b3byQgmU6Olw0dmk36PwW
64Cn16IPPdG5pTLMBxGtZVeAwW6Nu6reHeZPaPUXf65WXs07XPWUwfZjQ3yAC4EWYmnyNF12m6lL
IQ1F/hvKTCTFqV0+GYTv3AVcQYFIf/glVVYy9CRtPiBBUzMfSEvFwLJIbaTEewsjMLPFnpqOBuqa
lUrxW2ZH6cI+XUYBGpbqIDJuNczpfGDAePF1iPWt+ybUd3aM5UXYrqGvdaKYWdVbBCb9DaV9K6HN
HLPYM/n/5esE+iZ0aMjOuHKm6GIbvYeP8xqh10gkcGWAIU89nr4uGK7URJAxEyJ2wvQvW+DJ5r6c
pvlhe9NUPujAAMczbgRMzR1B7+K7fhpxElc6zp1DjW+q9UAzWF9fPOxbH09VxwnMZCyV8QEQuC35
xIN0MU9Ne6qB54ztdUOmTjOL8NL1G/udChxNjlbYhqWYxGWs0C2CwbiOEwp24+3Fh5oF7v0I3JiJ
ycdUuRZ7DbARRjFeAFzWmVFALhTpM8gGHyUGpYe1qtWhNdYEpDeaHBhUCrgwN6h4jMxOoPMYeNqp
hTrJ1neZNiQ6PzTNQlvmMysMEEq2VeL4/RHBO2WCRW9MWB6TxVgR/kBa8xRSFl+9P6mX+5xETYro
PRyqKMc7pr9dLHHp/SmOD/DFWapqzKEES4UrpWOtNmM9s3uMKXwOkrUj5IebVvkPQ2jzO6W641yp
1hBCOf+Fp8iCpECPrGs48AwwLZfe2JFm6buA22GfIlyynS8eTjHQUlNz9dpoIp319bgYC8Fw+cK6
bKFDd4LuEJ4SEtVKACUA5dcx6jX1/qxd9miWoU9jxIqponQjL73vanVZnsVQMu5B3QfdUxNRqMJ4
SIqzuaQLO2w09FTmVT3/GR70jIPlGg1sY1AcTb8ctYtD6tZtFaJxs4DQKqFVOu47kkNa0OYCTCQ/
xpwifoei6hX1mVruykUcmBEBlWzKiuLVvS1geCCUqt7tJL6BaGFgJo0KdWMebVzzk81lMlJSMzRW
kSpdzrBfinhGo2iQFPvDcrZvqf3ukVYzfvF2e2SbRD7aUps90Hv2MQ0wS3mIVP27Ov2GEtdnsMS0
BoIaifO4SVtA4W3x6Pmflh22/hE49IbzvCWiVYtS5XPzYvdIrcFkAJoyChBL34eUWtKrk1PgCoQw
b1MqlrrbSUL8u1G64zhvNZtc4s1OM38pPSgA9vVoGqz5mnQ0TyHtr3DqivxqyUXoGPQe01O/Oigw
1Ym6YXgqiEFZL4LsD+A2CZvC67H46Q/6PvHRufasDcXaBQde+IvOSr/+zOzzqmYipmUTZWHc+W7S
4vL4pYDeXypeg2+GX1fHVZdYaF546uEV9NFA5KblkPWbTDxUUTv2ucPv1KKii9sNn31bMnXKEtjm
wQ1T7UCqEsIh7x+3cvCN5rSH9KvNkT8F72dIikZaU2q2JgDXT2kKR1CN+dKLK5ivoeBOzqMbkQFB
W6xaXizwOPktOBKfSFC/e7uqD9Jo7BNLgDrQg2Cdk06cn1tJTm9C/8IeqCUngHJwtMc9xmswWtfo
fSnKvfBRJIX1iFuUoDuQ7O8UL9lbBwh0ec5QBfBrBWO5aswhyyqSyVtEwhOfJwKdbR/wQ0Y8G8ux
Jf2eJN+0dpwS//Qvqqrbfa4hWKhdR3+E90XW3ECiyW39hWMaeiHD/G95tp+/XgXxtsRCNiNkZO3R
CgrLeRdfm1o4GYsz/PxdXDr0dFx4K9Nito04PknDszuHHaKRZJF+IUR1HiMhYQLnKpcXoBfwr/Id
853nb8BAvJwJaBeXCJRJKVZylI387bvfDCZ1ZD/EALeAsKKv9WDrgSzZiIIiHQzYPVM4aRRtcHAy
EEihx5169VWMFZ42QCvB+Rk4A5wp5zOsAsAucl0uliedQA6VHlwBwTWHyeB0i489rqHqLCio8eVC
UIiqNiC/+ipWcZq3xIZbZz+yDtwByoaNysgtLLNudXVETTauGWescMf2cIuWTmD47goW3fySkYpc
F5tNC7wTOcI+QAQ0AKlQnyatt3QdFsbkHNY+0t4cAut4Hvj4vW7EaPJUYWWfZlmqy5srDNRUGHxO
4Z1ral5ZCXkMr7NBgmdY85sf3vFim6umSQtBreTs5UlpshhYwElikRYBWA07l/DZXaclxabLIjXh
v4UTrGACiri/yjD44rf25rbrpmGy5MQxtRjBbE6aT2qVaG/C9ALrv8omg9Kw56dN5lKE/93LfXX6
elJn5OVAGZZ9a72sD0pRSZFpqgDnq/HLAoNtdORgNUPd+z8n7hLGnjnzex0NlIR3Jek8vqQB4e/N
8qZnKRq7fbA5XgO/P4Jz9YsH0U2LAxJ/2O9zgHSoYjfzKDosQVidcEt5XQBBIAojemBodzmun7m4
GXC45Cp7O9thpm1AqgzSP9eyAcNwBMgKtm4fLnZh7yADZEs6yAVSy/2g1HCR/pQQd7CHTsUFJZEa
m5yllTK2/lvXWQ6fD2ASNH2DEviKBGL0/PQFt3mlEsuOpCODekLTQgnBR7za/x/d8Zg/dAGem2zM
7PbZkrE4a2A2RZJ+pUiHbxo9pcxv2MAf1vzCl4TrV/yQAAWLyG65L7QQkknpqCaBB/YHL/IVwZhy
qKNmBXomBlQ/I/Hdl46MrXE1b3RR17QawPjB2YxkcMS15R/Xtj+ihj33rItdH4vpRTiQh5XqZEZA
diXpOW5POOBfVDYjlj58H3HnDPR3QY4WL8sSSKUh0iVWcPws23Wn1bNqYrJqut1eJm7OnfWyVFjB
CnqZJmPKUvh7UQefawq408PijUfJJ42dZ3m158CzoaJGXgSgdvHbsqJNKxvNuYZLyGb/pCYhqkrm
OBIwwvPSO2PekdhCA5j7CF/XoQccLitNvtMpyX9WNcWqt9azON38uR+c5GeHANIdm3aABmUZEumg
WgIxKzoS0UJ0mPZ+nnLL9XVRiVdfd1NZr5lDxmYy44dHyuf5fPibErSa3w91loWw4u+vEI8oJUus
/ERB11CD8/RTBD3WCiKdoMdm4D8wBslI63APu4zvWuqNGWfeoioN5wiFnaJP8n498iRcRIxZNBzT
sV+s7M8fvFG033H2kg74MzaZLLa/AMQZBeuywDJ4BVpI87KRVivXEEi5P0y+95iP1GSIe5WsJM/u
Rr6/piHE7oX5t5gyaJ9bT8CUcOovim7vsqw5G3EzbbpA5XhTdl7/7me4Y1Qh3CyCOOLl5wEbQrAu
Mf4wb08tyTVyP/ElH8F0lTw/bQ+dhG4ULEZCbTZgUrwsqVcMOlJWMXFRKWCu5ovw23SwCgsoggRm
5T8T2wM1eai162U2XA8rARwcqiqHytuZeiSZB8nPL01zEw72NalFg+hTPGVGTUujcYA0LwG+qzgn
Xlxu/B884xubwBu3RRfnqkuiwWSzlZiO6eS+bAkNoI+0mVyKwTmRSzy4JTaDVZbumnWxr1rg22hc
d4fdXk640ZDDnOJZj5NPeBTf/brssfH7cXrAtETF27Dd86v4OzxV6xkXIotsEYbFrYb2eG69styN
t588m6ApRFQBUuRWau56+O9a881zFZMm2D1kVwSK3Nl0+Il6k4/IpIIctQf1CTd/l8GacO11lztC
b1AJ02GM5LlWMSz2LMuZyKeuViaybuX4tK0qX4tGcJi8yIt9XJOKIYwoHLTH2WtCs+H4+3L3IRsc
3qwxiIlw9Pkn+qbAA30H5avs2I3/dUbIUZne489riR3ZLFftGCD5uunHbgmaF5vAdDpsY77NJAGN
tDhUlUexkEqt4Z+YIJBnXVL0iw5jeXyTL1Hxs+wnM2dlxaVivVIcu+rv/2tf/Y3wTDrQWG6P7ZBQ
+k6ecLrfG+S5C+s6wKB3DsMh3Btw7u6hAToKAsDWS4d4Dds/XZ2uuzQ2LM5Wre3czcJNkXSppVQP
99zBSLwXErah66xGNcIkJlVfpSR90FabeYSt6+2O3v/BvVt5vcJ9MzcT/BjsqredzIZMaDp/Mekq
tqHz/2ANM+fhdVsMrAtIgBTSBne/kfJhXKWIpnG17PVQQ27ph/3fMSbUdyDbhdVmSqSV0yxFRuHL
DxH9R3it2Z6P4HfY+aJHwwmTpmTeFM3+K87tqcXtbt9UEBO5mdzYIF2ALcjuDfJPsE+kj4xsvxxW
QUP6A/8BBwikAtYfHDx7MnCjWF+i40O37W8CHeveI+Md6pL6t6KjpvKLA1zdQRum24AiEW8I0w1l
R2i9/Lx5XTMg1fCknhb+7AbM1t1AuBXeZLihart8GmSM6PksbIgdn5fU8Fg/EDqqYE3GoDDgIo07
2xJmFLkyDSqFk4vkxtPGoO17llT2OMiI5BHnFQeQmDTKXeUfAPk9mgtfkBPLmv/+Dwl/SsK0XpY2
JvfOgRls0YXE284h62uDVtJOFP4Hklzc4GDInew+dE4WKYF5eXf/m+wvbPRcEA1YTdfiX7BS25iP
euZX3FrWRrrupFV8BSUofLf2uPJVaEIxpO1aThUckpNFFqN54iMt3WvnedTQxWF69CXs8buhtznL
s4GX3h+QmGiIyt7MqZijQEGrJzSNcZX5oXj9aZDKt4xx74sDAWxVLrgGEbO3WQyiN++9zsVGLAG4
i9ZZk3OwoLcBwimkehvb+VZYRyozSZMLwM6evXsMr5mg3hxZuDMg9cLfiT1Wi0okQX1+sAk10Q1j
/+q6ng29Qc6ugDfAgCbEUoJYZ5SvQenUI63Iq7fQvG4hF3Pgy1bhrgWwrGe/x2PBzyRODEU2MMEw
1XdymUV4H1t+6ZM4wDnbJPPfh8fpoUrW+8tyICJUa+CwD67k1KaLHJHdPwd9C5oiLF/ZDHk8DhCR
pqfP+vp6v+HZXT2nDHOfL6RZcaMNLf3pDsk2LTsdonalmyOxI40UmbnCS584UCxwFfvQmBRZT9wt
rTCladUUwJuwnKEeySerjXeQiIiyGCqlMN6hlTA/84r/L9Zn1h6hjNTxCC2Q7NoS7ENcqsJxCpSB
dySfzQ8kkxstQWS0lvMYERG9mavOsCY+UT/tR8rOz7u5oYzOuL/YAl8Pq5fyoaGenVrhtyQJF/ui
p6WhbCNKvVhkecMChjC8n5rQDknuzKTZU0hCSYtfLtyQiSBKSVP+CVhHi05C7BvGaOxrIgC5XQlD
26LIZY3R4oUZULbJvZ2wTxTjGhpk2BeW5QNqnQ76RkVcipaq1OzS2QmVJfUDQs+jGW4GWK+r54+9
0SaPEY1fzeg7Nkdg0M4mh9p44eMpOpN1/rEDHUcLwNDnzjBn9jQVD1Zii9QrLxie/F0TeMUHeOK9
csUXGIWgrnjyCUj6T5bwPw+wA3ueNKH/lXxUKtrEnqXalECRw/TzdVNftw1wUBpadEY77TWqGXQS
uSgKRMlnB4rB1E8no7k/VIBjeaSJAD+N4O9RDfTP0yc7m7Cq8SvAoruqHKjuEV9gLch2yh/okjGi
x5hmggUXFukDnBcXydC05h0hKFNsDLllLIkJ8gSNiKALQZQ15YcA509+JUE6DzmZeslerIBMQiD0
p8E9EIyrr7cHAre8UXaD3YkDXDc0dtYbuC9u+FIImhEXVkSXnD8XQ79rUB5C+6My3L3GVvqajBBE
s1nK2d3t8hgfXJJkXPFpF8LhojL4t2r0EzTcYi6cQY5M5G5lWbrrGFna6gTmluRE0ysMKR8Le/kV
GGti+NS9xyt20iI/txrvVKDNnUT2ySWPuxUEvl/M1InZjIsilbnMJW9z5S9cKvbHvZSe6KuRjVeq
NBgJ8b/0kE3oDn1qZ68qOVVhhy0qJFyD6YpCrllTy+waLjTgj5sqhSGIG4WwEGGx5RivQAX8iSyh
INQ5W2ClHRZptc9Wu0fGZSnDfB3QMzKNxZIP/MJ0MZ57rDdkxygURnSA3yiQYsnVlS+ZxQ9XdxLJ
Fpn6ikVKdfrzmgpRMIe+xrjXcg2yem846BP4dLDyLiHAk9BXVfv09dZQcLlkl04s9rotSlgDNx7j
xaT1YddacTDr8tH4s5yfxNCvF76bcIP9h+xR95jWkYf+TIK53QDdz5tX1GLtso+bx0mlF9fYd/t8
8MBHvuQr7kakxua9xxqyTinZFeRZ78TrejYnt1LLkF34B4UPNauzzSlNrTL/t6IFsDbLuaA332DF
5kttWH7FDAfcE4ILKvuXpnyMWMQFrv+P3J/rC6kLHGD2xKHypCPmuGHInVrM/M4c2NH2EXt2lc5F
y5XkUT+7mgBLO0PpN42UWin/daaBckyyNqMyOIgMHfHvMOoKf4mXJ9/dHUVGsDhQRkjUfBDAC1FL
oyaaGga9eKZivkLJ2/HChlcdXlZWt+188BKVbQcyp+UzCMm1RVXtnpQJkJOok1LDSXBpLjQVlIJu
Z/kr+XbfaDNH5VETIJf94KH934EKT4/IeztzgB+1cJsqgZvh5ac8dJSGtASlhW4SkXmv/FSWefcy
c3Yyqshg6cmS+R5MHYYQFVGrXmyE+vEYDDeCuROsWxPyqcuj03PcZmIElUnH2dTBQI0KwZdxqx3Q
JuNDCwarU2TtZEBVOCy/lBikkzQs2N/KcKGniY80Vfdh7MghZEI+2p2mAMCHp9E4agGqhKiAFLbq
rKgBi2UCK3opx8GuCyu0AG1vWYXzYzEWlP4Eu0Fvs3Ar7Kiu03k4TBGp6YzcFE87mo35+EPRICc5
x3Acn6EBk1i3cNt4iyeC8BtwQ03b5IlWdfpEj8JM4kPLcglHSe+t8riXJ740SEIp1Rk3Li1iqD5C
p3a2k7HV6Zbe6cC85W6L7AnK/IBV5LiRnOtIa6rqquwnG4BWlUsPtN9DTEHZMid4AJxdwXYsqziP
yqHCjiTC1Tz1i6aWQbnqqWY77ipBKdJjdd9aGHqWvV50+yVbmNBYyXEt4vDyl4BOQj9KNCJE3fMt
0L4Jo20STHD9js6r5atNJNCx5hHHqjiD5RqudHrUXKA9T8TVW8w+gq3G8CYyn+sDcWaEPj/z9yRh
Tl5gWwUz0AM2HYMqFbQaJDIutF/9Vm8Tn58+gqiArSkUf+oRw2XGXsMb4K8VOtFe4+f8RCp4WaJ8
R6Zx7MzHfqiyoAs6P5MsFAkehsZ+4nnPAs8vp6t7FViQ9aGuT5oL1AGGdwS63LMC6/CrU8YH7vun
7ioYwIjqra6O8Fx2QdCUS9TBMsHLQ0DTXgZ50lIEoqggnckiXUt4E6DlA6BWqrJGIVShBMb3o5mn
3yDN3Z6CwpSAFj6tdGr/MbW2ugSzWpOW1CflcfBNTyaQ+cd6Ism+Xc3+V2vVbOswf2IUiwvUXQ20
QlRGkYdDKx/wqpr1IKbyrkk0o7ze5ZDVZYXE3CQVqL/CdKcBjcZksDle4ct+TQ6rNRB1UtdZHfkq
ac0x1iQG9VpIjYM+AloRwP8lCjgdlNxTGsNgzDGegdVqk1INt2kVifJuhueQbESHYRPPIySsBraj
TeBZgz7f5mSxdeiTSlsTaVqX3SKNob5C6eMqVWw6pJD3S6IIsc3uVuuhrkMlvXbTvicAcbS256PL
o+t1d+3UB1wsKuHtgIKiFI85GKm+LphncU1sxps3hjcGmom1A1O+nQ1QUYdYnRdTdNlUp5D0aO6p
SKKFfrE2YdTtU8uSET3FC2V9CLjBuUml24zA29rT51PTzjbW/UxOe3neuJF35nbn5y52WzNR2hwG
gjFp6hmWjzzi3M/Mh//cgq8dWljuyTvi732lw8DAbsT967YkaEYFczVVMDkthP0aHNXsfcUgT1f2
7eexL260mJLiptOuqpplPYmDTIATYXLfXBk9YHjz7PY+HS//nX9ta1a1f0/HB0TBmLq2YaUgHLgl
gmBV/NQtoN7B0Hti+wd/CW8/NHZMvw1eQkINVnP3oRl1lvEuhIRO4KaRcPz143rC1pBxj9X/5aiD
fNV5iztEhk7PIFqZbvJf5k/tRsAjuVu1aAYN+T7XGW5NOmVyTazON0ABEmyiUXA+aNGH75UGNGFp
u2+6IojahVH+Zs3vSRi9fFswjcuZ+LEXwSCs9yl85Ntz7ZdEc5Kd7JoiPgrNb0jvCsnwA1nGyscC
4MSWOdfcR0f6GSVx79zgoah1vzUmnBRICdPwdeKUvXSr6ItIN4BbNR5wycPPRgNfFwYhObA81lgR
oKwNRP7Z7b5s7BgXAfHiDGIc6cKmTeYrO3FIj2znB/74e5nsEGzvMpuH74PKWOe6zRLcr6Bf6emS
0NkfnaJ868ZvlXYV8a0CcPHzso8fqD5LWcHP0Z/eUM/vu0CqMV5hCQZRnZRenwF7oORb2eog2Oi6
dS5ZBKdW3KkFmIdghL5uCEsK6HnC0iWA4kjCRLR3ouly8XI0oc7B8vdphZawYamsDn4xjnYAVe+F
Y9ZkZ9EPhw7FN8mPCA1/tVkryTwO8Kp6kuUcMQPMWXMh9QMIhY6ay4x05WgyEZjzt5oDCF5linAn
Qdp6DN6ZybnlMbT3clMHET6lrbOtmAIorgqqiHpyGTQq4iaHgaJTCYiRpBI0VHpWVVmSSgsBRBya
hj8R257xahK7R1qYftWGATYJGD7z2V5b5rDaxxt2thqvvetyzmKKCDHLllP90FZqog7NadIgJBPL
g5wpeWLszvCJgdtdvP+7gPzfM/Ud1y/YLR5VhMkqMY8Sf3eL2I97hAqoe+KwWu4zpgi15GPTqM5c
EhFacnwnAr3gPoJEKO3/jzF6BffqPrV+wPXnjdGnhHt9GjwZFoW/gEShnGZF7Xl4L6G/dhTE/ZTf
akddH1qxL5aCe9SsA4e9gXnMp9PT1Y7igojuHxTSrjoZ3Ldm62dzw+8iRPdb22xkGyVOW5fgqNcw
bkOrcu5Jglxx6vdnarabt6REOPqS5B4ZtH5Jf2kVyQg091lLYdrgTZ0V5QwLRU1RQJgbXM9BVf6Y
yvqCaThD5cq+kam8mLY72nAzOg7O3/LBUx3Kb63fyTuDl0vQCmxYlkFP1jSDHOthySghJtbGL3YK
c7LCFm6sBdHShkF1RPs+o6yQaKluJqLcbztNhauSs17mK63AkR35NprINC5io0cOO+eK/XvoabkR
EROPk3w1AGJ6/Iof0JKM5UDZq96EGeNOagq1CFgO/JvqpaUsj4X6goDry3LWlwehdvZrxt3fWK6+
Xag+R9pllt/vxXcpLtjUOrlgfn8wxTfuZPzfdN7t9afj9J1qHEjwnGq2gibqqupesrOgIVtY7dqJ
3rRETkoU2kMBUj/B7pJaUOxwkBYwLVVcX8vZm7oaLPRLF3la+hLZ+sPcXHnybG32XSi9rVb65vej
0E1BuE0Z9YX2vBDbk0lTQBmgh5q3OgV0REr6H0GhgbOBblo26KbZdO/yF0+6gprbFuooumDJvGRk
mFqFzOOSKVmAIuK7lRh3hd9n1NKYDMTYXmc4yCR/Rys8zh6+Ch9gbdK1skOkFJoXcvpWzPkEg1vs
Tax4ocxp/4yqOl1EFIkx2nG78pTcAJ/msl8rwr8jXBYphU1UlvO93hOHg8KHkwZuA1C0jLZT0xL4
Y9RXKB3jzrMJLKqFIww71q2gWttRBCAenpxQWaiAzo0HLSayy/WjwOAtQva4CWj2t+gGr5lP+k70
HtLQE+UANOaFcucB+5oCQBPKNrLDwW1AdPnaCF128H01TuqZvjIbRF2X4RhzKoB7wl7tz9PgRSHX
sr5Ji+q+j7RLFGOQRIP5ac4VKCqSQq55bgUZslAOQHLC8d4mkQBFimdPcPQedbv0LxjEuMnLohch
5yaZS0qnWWPkbqcfaYC4bySdyU0jyF7HATzAkLw8KehNB17xFRRzEql1tzyMW8RdxO4fIZWAqW+5
UmiQf0YM7Fw/sY7HtvoVxD/cIZYeCG9kHZWiI5DO0F9RCOT6J50wEcgvOzCs/VAI/HPHBSzCkRHi
TIyRh8T6BoRvcyRi79uoMh6vvhzJEf0p11WgQgkBm4peI31LxwJWolvh7f99ogJ+ppehx69eYoqF
DwU5grt6qTtbreOsuyMpYXePcYJzzpAa68ikPDdwU+7vM1McDDB31UgYCUdLztNiGeLRw4i4ZM4k
6c90F+7b5GCo8JoINrDz4sReMSuDK4GbZhxBb9KcURf082vrXEVKvP2RjQ+9NMUawvco3nNdIzyM
uf/Oph+nuJCwAEJAtLNU9+1gBUo/gxbcCc7zl/kzs3CDWUqWa/+xwzaWkckqXgkKBzgR2iQML48Q
FE2ImYxxI4fI61nZ8pdQ8J3aHW66MMEwirFdOlLqAXhICjN72mmo2D/Q84la1ZuNMz5vH4RVLxwO
CUG+UAd55IXlQehZpoFBcYoA7haD6+dS1GWxntm1MW6AuWAFk9l2WxFNeHYz5pBrvduei4SrpBkC
hgdOtySEjV6Clkn8TU4tRdkDIcUFHOdS3Qys3mGiVs7/DEXE+pcWIl49xG3BiXTbJCe9WOvCLiVQ
bGUggKeWFEOJt6/ymFyClWXkHBjaieOhRj7NoLyUT6cbBwLahvnzRGdFpGfq0iQY6jehR7e+QVp2
5oSCVj2mg1vD5bQxVMF3AALmNDsfv3dpl9xYZSSP39uJAB3ZxvqlZDnHJzlZZYMJQxqbIjcVKmbz
rFHh5ek9LcM3dXI7+i5ZQfDrn368yOOO2o70cnlm8h04RpYpLTVRodwEiEtVCYRh+jVP8Kzlgnud
vmZ1/vcnZnk6G0RzPBX5ZQMoWlCf+h03GBIjHfvcY8x96CevZQYb7xN5ewt20Y6Uea4GyFCqxJlt
wxtvQRSeFoJKYXA6xTcUovRJQiAr19X5hITx0JX2l5kG2AaLY76f3ciePNPzYhFs+LU6KTioJ1KC
g9eMAQjtxFaiYzIEU/GCdPnYr9tFBiHiGu7EwU8ZHnezEw+RWdZMYavu4Luuz4M0RFQaMtQRKVWP
ZDL2iknA2cw9INgXS3Pmyw9q4biDKTDKRA5yc2HqBZ9AW3CH8BPinPFJL0wo0plDA4oj4SqOEfXk
nOyaF8R5q4ZAur+Qwdh6F9WadU1pqjxxLR7Kng+9aMwgsOYRzgAYdbEA1QG0cPIYPeoOq7sx5xY2
N/uZ0NzMlt0ivt1S1XqaxLOHdfXFwDjO5xEdUfwbGyI2tLq4r815vZ3H5nbUYF7HQNLy2BW+dsLw
IrR+LfZ2sd6gtPheyZVRu74tWKXyRa1QHSdTrYEPrDQpNJsuRf5onBp1Nrb8l9kWCCfITYb+a2NQ
w2TLzVF8SRGw0KZBfDLgK4vz2f3uzkeIxp+HxXey2LKovrc31KEpec1ASt8HSr/BtBd+JWq94ygd
NSZcGVW85X9XGkgrCFUgHh2kNjZk3Wn/ePJyxmRb2x0zqlapP1apucdYJaIefz3O0g99XDsb4HbV
LdM7DDUwMmI4ptmElSVQMXvdcbIUqRmdVNB2xrY9T/NjTrYk+DV5kIj+ie+GOCdjnE6cGsk/TAXC
gKVJP6i80HVWBf6+p/uRsJTWi5Rv6dwoEUBoDCPrRsOpjcgQKKXH9VL0tllLRhoU0MxB6kz7xFXW
CVuxV46tEo6O6SnDRNRfZdnfjJFT2WY5grX0iYHCcNivA2+Y2jXNziBVu3e8RPK0fxjddmMArvnv
iojrGg94zdFgRUr7qIjGkcjg4i8qSs9AIJNEzi+V2bq8yWVF7HSeUHu+l4leFuFgo5lSGxHzccd5
xBiGAwOFKIXoGbWGAYkHfiYdFSvsAdTUUhz/v5GwDgOl+8XXypas0z4bRiAK/Ih6D6wrkECZxSZp
E9CEGfKtBSiuu6/d5jgKZa61GOeoNZGU2yK789e2xwxUhTnbUCAEcBNIGezLMKb9eAbNuDQza0LI
NxX/d9fta7bV5WJ0oixaDPOZXGNlNt84mBEtxcROzbUIJilYc/r2jpz6Xp9M8AZhlC6d1oX3Vvek
+0BTJk/GwQ0QU7iqoE6N7Qb6qzfuFB8mZk/uJ77Yr0QFWuGhxG9nocPCKqIWljhSbkyaH5/hrF+n
HIy2d/jG3HqcUvmfbPKEJD3ySWKbSxGhpMsWBp7EDdjJfqpINCzCIbB9rcXAUkTRr2vHTNR4LCwd
v+zBtRz6KN43tNFJ1U94KqgL9H7C6johoWZ0yNiPOUfGdYweIOsGl1KOOOHmr3TY+MxUNYrfsJ1C
ZIirULWI17RZc4KkwdyARJ7cz2WFrqAdqLlrdb8dHLpgfcPX0l7GMhHKylVI0taOqpqf6V+SJmIj
08lhj5EU20Q4gOaCNtK72to6h2y2EqPq6L7LMQblyuIad+p1+jt1Ru1THZzg+S7iucTrXV6/x9xD
JjLAyRrCUCCo590+ciDftAOSLV47TA04StkvD3ph9jwXVH+IshjJxGpceZPwf0QehDZffnnYWcjL
xJYjut5On/kXYWdWPE6YKEBnJUIgD7CSdUqIO1Q2hKFe/MDRa3K1x3nbmwXRSS7CIPRD/m6Gmxvk
RE4vOLmDH154YvFR4g8oOdHqGADmXLMevhweZFA9vwOqaDnODpSvhiKAgtVi9ny+dodBfTH0gLzy
Sfj31gD73mhWHTH9S1C3ZMLD3ftrVgWSqaIssyO5z5ds11kiUVUoKyrW2Ko9B/JsxAm18qO2NFQV
tSLyqGW8ErxjdStpfn7d4wk7Gdi+6K0LA/StszInvPbVVwM8qEGaMGtpgEAmMaCozCAuCofaKuR7
jrAxTKfVpI/W3HPceC566ds8QXqPtbepROjy6AXbIe0YlNGyfLeHJK9m40GTNq93e42Q9jzkAnIH
n9TfFWHGo+arg6yrmImEDsn2B6iKTwf171z61+2UZmgGN57XP8M9imKSOxmvGgx9subXT1r4c1aP
oYkz0zdqinz+057rbC/+krB44bucp37TPdy7OZV0+p22LN6H9fLhuchJyaPCz4As0CY3cHKPV/Lo
v0uNce//nvN9nxfE3Vir4vfWelkRdNAJ92oAhIIecF9oivLr2kQ6x14/6ztQ2ucp/M5cGRvNGPF4
9TqZEI0cfmGt/Dvg8+Q8UL8wK8BSUzSqcfvgyUrjrElwf5HwrhD5bxYzMuCzBIxfLofsK+ptEXH6
80qplOyR7IT1y20de8WZkS/A0ioeYL5fjDAmRl41AxegSt5MlG6iRc8Go5WFtZ1gqoN1WOvBecjt
Q4Z9MpSQ5hRLMAEMYAJyS/tjqYERdNFQXa7FCXHxIWet4ZbrMIocQLNrApJHGFT76j/uRfs+kkZ6
E+UveNXHBbaI4h0M0ycVnp7s66N/yMrwmx2TeoqXwBbtpfSEs+EjBSDDKmlVvvG/M+VooOLlhcBk
ICm/sJ8hu+HUWIFwYLjWu2AvwriAcVFFP+HLx0y0bFrZJgSdh55d3YozHLrV26hTJvNi2KARdJ2q
ApxhMrd29j3ZW66K6BVDnn2fYmXCQC44DPLKMszek/TleszQubulG99iGAq2W0nlbDfi/ZsEPYmR
eqC3kTERj3z/07KN81AQJUV0P9HBvas3tDIT+FJLoT+ROrcNfKenisqNXeuKlZBUQtagkjXFOP0d
QHsx/oI6/O0MwtuhEWhA30wm+Y4w3JZkcwd4up40vIpN5W6G+0HfsOXSyHvONoLT189/9/IJDHdM
XipU9uGZXqUOiKfl1VPGMdrCodh6qURAxKR5Z/p2Np3GlHy82ApoiqAFjNhlA98tKFMf6NQAmZFm
Ecil9LRJkEGeRPg2oyr0JJWEEFG6V8uSgbXCCnkngZhwubYt/XlBZ+Cht5IBrCy7ceOapCgt/sM5
PM8P8oKfKvA0PyKQqXnDPWClyHC896zW7yG4m+odmkl5MednexSVLY1uksr0N0CuA2tyNMZWpwXp
OqH++693ly6SwlK7zF2FUWgmfvmma6umRDcac4q0qop9wclKQJ9C/HYjR4qrI/FPnMjIqN3qNtny
GYlliHP4hpd2a7pvNEmO/nDYiDblNMXFyK5T3LcXHz65MPoUcoJUIJzCytk1nRpodRXFi6QfBhz1
7vQYuYFCsX13Mdc2HfV/r/H7HhLVRUMsEfra+W314ryi24Egr9HTIfo0fIw5Wb2Z1eTsBfbgQVBm
SdtCru5jFFwd5r27D70lGGY3p9+tOnUyIua868rdAJAXYB/Pd8PQGykKNMChJ9ae08NITYAvyCgv
Gcp0V94gFZ49Fly2gNchYsg/WmWFcNo830BvCEFAQpbLn071P7jcyYftDl61NLGvisxWFwcmNNSz
1ductVg5S9f/zfpdMXWMU25QxDQM+j9AHjMHm/Ui+mDmGveT6itTg3qOaH8eTpfawK2r5dBBAjaR
oZx1f31c/dZh6S0aLIJ7mqHI1XUgbd8JGxB+HJRb+67it6MgTNabltEeDsTxn+rtR8BNPm3kL61M
zVS6FJNsxijpnagiEGvQ75apB/5MbR9BR6P099YHwTc6vy3oXcpp19GOMPRSP1ZJkNWMjqeOpfIS
eblNu1pxwKByqB2hzQgxt5FOkS5kKnevZr9ldDXRwxpkYn17sfIZ1VqTWmn9nlV/VfozgKRkeXpL
zJ8Vks2ORw1+EDEKFnf4sN5DkkMFpO2DPloIrRLulRYpX1DhQEiwh7RovsOTq4oHUtJfHv/wFF/a
zfh3UgssiL2g9QnKlEmBQ56FAHPTacwwZe6RQHXkyb3WsE4zG1HMS3UcPbtaB0HGA7p8MGdakaGj
672XWtLRc24jH8m44udSiD0dhF3Vnnbba+X0AnuevCI/U0p0rUyrEY94dpvbAsQZXQHbuPREt14l
wPLNQ4/QGEshIni49TCe/CEI9bXTV5ksEL++gIUNFcxkpKyDM795Bmo1JihAE4Za/pcTKgnm1NFN
D7eU0gE39oZ2fUS0qAlZN4ANciNNPQSFmV6B6HMfCN47w3RAUZZ/Zl+Y1T+jk8CbpQqRKutDAMU8
q8RZ/TrRQvrF0uyFl5vniZRgn0fJfp8zT5sI30K0DPywZzG5YGc+kXX2al6NeN4UU9kzJQLUYcY7
ht7Z+DuakQqj+6b4l29W7WeQVUifEtm8P2ExtmORErqzIZbZnZlVyQ+M4Pq6n3xrwahuXpxGr6Q9
xyyvm4dpLoXpZMZguc1HcDGAuMbr8yf0dm/Svxw1B4PzrbthL+j415tADst8TOMiroKsI1YPxHtu
hz06T1l7+122YAXgoGy1zpE5eLwIYnMbJiER2u+jtYH684C94wmsjWUsncDcstQAoX8IDNeY7fDn
oWjCVqBTdWxzeZ99zeCIJTW5lvpeoAWCww9kB+b7vsWKVJfvcNNfj3e0WPatvc8sgTT4tyq+v9gt
9pg3c1ra7kYTnsOGYfwKg0Ge3XT1Adp/9/B3tUrzfF3DxNhdaeyihTJqnaO4p/AlBVTZtY7yDnyB
5RzdJg+svygNl3pZ703I31yPYC8aDGEJOpFz0ZVg4mbfL12BmkB54L+Ws7PWPTJA1u29qret3eHG
+4woVYHD8MgDH3b7k0AJf9HOWGpmGPzFasMLztcqIKy603P3uNpXvUsFeij0lBejK7E9MFdv0iip
YTmmOrwbgNh0PXAXMhXW900+e9PULUrInc0Ym9frm1W3wpDspjYL2NfBqXNnQcHIHK+AsR70hfjb
UkJ75HP5AMJZsbfox9tdgLMbW8l+97qRSitxRyAve4+KRYRRTgCAnCiV06ZtrqyeaihUdm/kMFHY
7vMFK4Mzpd+tyOuG9vFEnT96s1AUAQgA+PHWbQDp0jerKS7rniVRQkJ+6A+IIIJKd0Bt0gPtHEUH
nWekjILQ8oS6LGfA7ZSae4O4aJiP/Cv5ACQIXjcDWzBGjY7GrR6nOUKV/NpGr0zwLfc7MhtsUVx9
e6saj1jpeotbiJxS1YuSazHed3ufJf9SvTH9TqFaOGr7XsXj0k9gy4ae671nzUUxw6sXS+mvrYk1
ZyrJ3vfG/j39NPatXZTWZYurhUDNwJnmAsF3vxa9T0ceuekKwJHrOB98mT03P5+YafC45IVliCnA
OScfU5Qfz/BPzA7dBOUkb0ZHBSEl/auYOcNbOMMELEb3AT/We/ZBMKE0axxMk4ZosfLRRluyLicJ
sWLlVgMxXsZCiCWFHnuC3ZpgJZYnh85ajOJmasARMr9r/sZYGCqwgcKuRu7FT4Q3vHAuNCyL7VhX
DThfD2+G7JGtTCkAEJZhTqg0TD+2YRNQmaNXQeO3ZvH24u7uH0bbHN/glZi0yyN2a3d0hF3carHd
56ekyozgr+n0KkoB4nu/B99P3MTxyojQBiLnIHErKUkEOpK6G7hVEyIY3BsRgw/276ovxiq8ohdp
SiaqcnBJQmMD1QIfuQakdJkk+Mx546jre/PeGjoHvzyb0xLh1zQ0MvBg21YxOT9H6W+9KWgT9iSo
4DD5Fax+yoQpREs4cI29fANafI3CcVS3NCxlpxF2GHaxl2z15GMNnFjqCqiDayISSbTrIqo/zIdv
A8El2T64GFXhIE2s63akTdk+0ZXPblvqTRQXTGX8WfP6dL2h0voCh5NyVqFwfZnXGnV68vzzX1pa
fzBRC1s1nnpFVW+X4v8FpWi3KMpyFWqQBmqgVeiZH5C9e0Qz9E9AJ40sBqCX0+4tOajHFvZNY4C/
la6ncPRZ3zOyBWtzK2UiRkzdpF94bupxPsBRomN8m+qjEa9zYMf5aeQ9W6Bd4giuIxgT219QgxDH
aB7PrvciYkeFC8YYa0uy7VtyfbEFS9nOTYbN7kG1+Gb8u9prlnzjXtFrsyahC9t3ik7CovCNwexL
DpVcfeK1xQ5d4I2yOj6hjhHqHqMcndGarkF5Q2sZcjKPC62BqoCZzKh7Bt7ELZ7+27xTCtA4Whtl
hwBLVZzmoWkjSX0lQefW01D/0/y7XorNiLYepJx4XRlYlAiFiA8U/ToE0GcIVmPZueomJJp1wxEX
gWEoxHZf3izW+dx8iTh3vMBoKM+vtQoV3WDihqBmY51iF14QDrMskUNIPSHlWbFcDRIe1+9+vpxb
UXza8T2aeKoIBYXo+3Yi7R3jRZNWm8y0A67bUIafff5C8av9uglam+JWkl0/WfkoSuOiRNfXAS67
PNMkjBpTVryM/DKgZvOI/dw8+nH+6GOwhQb8/ujGJPlTudfWTYx/z1jV+kfcUZGA5lQNQS0UFwB9
s0sShioUBMeYl+QI3fBsLCxULREPxyS6WxSLRxG8sL7ChBd5wct2BAT0TUvVMo9WL2PskcfR+hgz
dPrQ4d4zO/7Qfslz0MGt+6/YuhRI9slMZXh15vb8tdXmBrmTiAm+IiviXkpzDbrGt2GwcsWwfcPj
8a591ocE8ustd85yr6kOqU5Ni7TIAPnEsBUMuXeXxpeSyZGTi505abcyu5uzDby2sQ4gfAKahOTf
L0jU2rc9ObWnBkiWb1OZXkrNWCgYLLtzkmHEZCLJFd0liPZwxDW83Lxo4LSBsnlZDczJzz0SOyqx
8VedjCwA/+2DuzHdozEWHa7iEyX8jM3g5kla2LMsljlTrfP3Hq3C9fHrb5qJ4rnjRUCdGAX664ET
ol55deudJvKzei7J5kwle23MzpexWLXHNVxccrPADMXYOiD2NdKnNoG67QFkdKWegYEpEq1D0/+3
SyyOh+Wxb5YOn/IC6OC3gefeb2Se1Y9TnNZs4lEH7/q7iOKxzaGfDP6Y/76pKu1GpLWtvaCDj1iP
Lqb6Hb4ppPN2EV6eIc+HwL7RIU0e1mZVdli2LE+ywgrSM8xmhKWB4JNX8coM0ppt8v4Me6jdk4uv
jPqtcrLT6W7bWCa3Zpumm+Lu3+28/GjaLqo8fuwJ9J25n2voSB57u6tFDnHJF/7umzRJ+bUhOwNv
ucj9jBi0K4RtWOIz3AnIWsditlTZ6DpjRq66I4+fmfd7qukfwVwmtrTcAiG1H74KMh9m4vmvd07R
IzXC6qsAgGbklLxuxTbkcvWB2SkGAotorYyDInCjFMYhm2kAo6Lo46Jkq+HkRPcMV3JsY5Rv0+ix
v0aohlArobRGs6d7GU8Y9iQxshQO/JiONKPcnO5QWWfCuNfNzrFC0oxCD+gUozuGi6wD1a6RApRg
8uNa81SsarV8anhr/+3qXNEir4fNPaOSVK+iwuvtBEgjydHwhW6xfuCdmeilOlfUAn2lFqycjaeF
mfHH23bY3Nc0/42YwIALVOAc6JZe+IgoYFfEE9l3UfDvZxZDvH2jdOajRIuRIn+aV16F8ND9RtS5
Pp8C0Cc7UmW7VHg+qLobmD9x6/5lJMsX50nw99umVZ8EKDdF3HAovtD/mehQoyeEJ8ZHhcrlq4eS
fJtjWJnZF6wXaYdY5B3U02RHIrzLn8GNMSW0GS0PW8gdw2Pzjti6XECg8OPdcoWkNLzVCkXj9qqG
gK7RkUC5ZtL9qrdst3ymP8HtCC29k5M9s9p1FkiBgiSaWInoImigP+s4Cn0exao3pS6ANQbaAAUZ
Yql1pmEmGaUiVZt3jQ5WHGWrDgM2cVSliS54c5HHeitPXyhPl7WPK+VXpeIFk1PmOY6ckio1qZN1
1TW7F3hUPfpVgbY0XwAXiBs00GrcvXU/fULoMCAKNlRss3qzt817ngj+4WT/YRmHxUy3FFjQG5c0
24AmOv+twZ6wPVfRnmsGTFF4UCVco2e/y8W5Lj9WVy9orLGE3F6l5eX50n7nGPJPSUeChOsVMeE9
gdxS2UiC5ir78BLvX9iCHrnVYjv2ig3afEYNNIFCjKqvuUGSG/d6i52fEatOo5z3Vbi5NeT2gf6N
PFKmG/boINlSSW7k0PnB/PAx3IQ2PYaY22OJy4OrFh3vzRP6mUdURCLPUN7V2NKdGJGXyJOWpaRn
u9KNWXMST2jg3EQ9caEEOeiP0h1bDR9fVRqDTPG++9XnKc6gPuXxUCIvZF+Idf/eFd0FhLL1xlam
7pFVybe78cvWIsj7dvTiz4pQAuzaG8E0KiSikhpYxBvBjW5iZqAUzgbFrOgV86rEB9JVEovPtBPW
49KfgyFT+zXmyvr+cO3f4bl9S6RJ55Sm1yuICdqPC6KAjlzr3Mbo05aW4/5+2pFMZV0WTyFDAYvb
I7TL+2tiPUIulGbmmz9RJUQGMjxtyTqdaJyjtWIClbOlH8sdnYqVjzuO150JEfZW8BSSteRuKyPz
T3/e0IuFWu0MgOepyZP0V5cps73yBCfU3AiuJj3Nh+ZlROu9PW3urhy/m5TntzVzPuobBRwp86nr
tPh8cIlrNHrHRPt478ZIgDuCT9qP85PockTrsehNMNG4eOMu5zAaDAVESk8juV8KefjKvEylQqnH
cQJxusZZ+5+oL1MB7i5Kc9BTFLZ4QT1qREaBYfxD8xmXLUWRvL21J60ELhEPg5dSW77MRilcmDLP
4FiYS/YxRvNobmXpjRATBS7Ckr1M8t74HFMOcMmLe1zcfbpdUdMOE0zpyHC9OtBnjmoO2DUOK7w/
HVvtXCdJX93XldOuQqFxsO7C97tOldGb4erO6Ht0XSaYmXN1Y/oxh23q2wVx6GpQHTu7p4B8Kpq7
yTdbjG+fBg04cE/o+YIG7tRK14R4x9v9CsXvTe2zDtNW+D+O2QbEZzi7dbSHYiovlHmYFymF/KDO
KacT92yAxkvwHJAuAVYg1QiJRuCbYpGb7r+LJcre7i7SJd9wUUQPMYKNNAmTnV+JNGueNuUYoflx
P5otjA3K3bs565GBas2QZKWTk4BvR1JTb7pCLEpPY58SQ981Hayfz4cHgkxvUNhnU2MV0Y5WhUyI
u7HZXQsitWSkgPQwS9jI9roWK3ZfheQy3LuixNzRr53/Vhoj8tRkQYox58QqIxhri+ViL3IfKgSc
OYoctHIAYS7oLb3va4nN7uHiYlCkoLNEA3i+0n9M0ldlDCmfqtH7Pg+yD/TIxpVZF3WqB7mTj13o
q1GdkwxYbKRIWDaGXfQtHymYoumlJ2kkCZBce6HyXDa9p5jDxHSCtgLppvcT8r/wTKcuPv+56CZz
glEWFcysvVZ4ApE4g3uPECRoqV6Sfk3rg5k3KsJ8JFGA9Oe/pZYmrYPHl8H38HZwGZfXW01ZUinK
TTeGy8fO520hVVB+Hr62z5M8ti35yx4xalKqPNB5kwYQ4MtXadR6J1sSp30dgd+SKfZ1hB1b3qAG
/dwDBa89FxkzS+L2iBimQFgRl4yeTi4o929Ly3IVPyM7vJGl5IdqRD9PX2xgX2vpaezV1TP9HTzt
YyONFFbGVnVRSZ7Wf/3BGtjfJB5p06ZpMkwNcSHVqBbfaY1cv/Aggi9HrTPpN5iB+TpV8SmeMvoD
lxch+LlMpG6vxWZJ+NQfN9jZmJ2Jo0U5hZOgjXpLMOS3cvOEMmAE9QnkdR1as4R8eqldNyId7Dlu
K7uFEjh4PrCBirhgPOBeXVHf2K6iX8DQ0oPmsa0XeRzRixwcR2SOzrSXB4XKrDoueWJJEvD/T1TZ
KuVPZ/fcZLGwvce/ebuycD/KSnoOgFot49SVp8NGOYmv0ws9A4mZyUips5peyJA26el+34h54WrQ
7hDyZ4Ub/UwHLgNzL32IEDjvmuuR37rZwFmsIdvsrreoKNRm2nkbQpp+ODE1LI60zZgnfzZ6JAjG
JqtBrOl0hQTBz0JlEDqKPrrcSojYH14+06sparImFXZ7usZB29qfzIZ5xiAZ2s3Ccv3L+3KaLtWO
vLVen+Z/uBhNExKwAWgA2CtfoVYU/sGcbrDAEMeq9jrU5YznMWcow4HDPFMneCBPV3+RXWhv17xi
WOCkjn6/bFTOhl3uC1kZnHHOgk6zRdJmzvCStacW40IX4+Aq/X3If4BFkJ9vQFPAuqeQNCtqvn7F
eWNJX4T9spnh5f3RQBgFTSq8vl8x7W59fs9b82lxR3Rh11iw3gvy3jIB/MEQEuPXF3THrP34GysH
8hlcqejLAgnx6643Bj3AULcBUVLmjQ4vh9NKik6l6pR5QQuGn4WSKoDxLqQk5ejgF/bKnZIh5683
GoPhwfdaIR6U/1pX7DJZSYy4Y225qAmUDaHpn5jwpBnnjAEt4Qz6OJsl45uDrN0bRxNmu9fhvhFk
hUqAvHcvyjdzSP+yQ2wVMtsrIpy39TGxcA1qbMItMOPwmvmmA7vb2BfbCqrk1ULhVR/Wx8Uwisn1
Mb7vrRSEwADzM9s7D2lILUS8ryY7mMqzZ7YrDNRvP8TKvRW1EMUh9ft1rDZitJxDcxf0UY53L/hP
XKo92ix04foFX+Tb3BtnJqGr6RT6akchKMsuy9P7TGh+VgBFkCnhAeZc4sRImLzwoBYGhBjZ27EA
9bb9PbM+ccztzluizfWWUDkB4Pp7f9jXnG74Noi8QlB9SfmQXMRGlmHQbSa9qlN+VjdVxSuZKubS
FmENpnpgcXldWQ6HfYdN90uS+Xp+q6rpXzIF1DHFqmguqF62NKi5GDiUuJPWnxW7Y2tOY66PX1ji
EzNAQsdrL4QvrLANbZDdzVQkPYv+/yERrmEHXAES1pAQKuwp1QhAzsxWW08M89BwX0SEaJ2e8//u
9jcJylHoKgCFArx5BpUC8+fjJ1rMNNUlkFG9aMWrgYT6HKtuyPW5dqeF4wZZIFxoecfD+HgDwNIW
Re1iGYEABSP3x0Sub8Rrfo9lgXzevyDb/Bwyg+kuktFRaKmEfKGpVKO+A0LZg5/JuJY4rL+cXVOF
7IU2iCT6RlfjoGyoNLE0CFzMl0bTadY3lnrtlJQDazV87aWhiJW+Eg9qDHKjMC/HmfDVZOZoM73W
klzFXtnVLIqTxAeiuyZJZ8kcZcyntkVh4l2KeBsJng4Qa72Ur7k885wiB/aaY48X55afK/TJRMZL
nLV5Wcj+pTmvne5glAaCysMGu4wUr2oqnzyiJls2vmUrk8OtZ7x+M0ML7yYQdp0iMFnvDi7vqFxF
u5BGBCTqyg/4saYKSAzj8kJIV42bBc9l4lZJ3Ov51ipXynUI5xx8ObrHhfjWD5hddFD909YM/1wG
RE2Yt0RN0aixK0eJvdIrhu4rR/JeVeixR6TWpLt6nP5xpjDPR5wcBxlPEtgByeaTIijrrDmYc58q
AJo95o/Cl1zqLWhLtJjJqHpgmiB86FRX8bA9ke2wWkeqkbqz0u5/XJpXGN5gKjcdEJ+uJywifQoh
tsKlkeh31ngeCtsS7/N84lqIX/Y7fIwJP2M1ojRHTHE/1jt193qBjat5sZ+3hKzJC75SJ04KJSlB
v0BAU1WR5xl/vIkkSo+8C4LNq3lbtEVaG+qFgmXilu+3XPQ7v0wknoHxwcMxr9CnUvKEdYmS7R4U
9uL8HQZXNeFDEPl9lRHfS1yRiRFMq9H+RI4R9nkNe/zc1Ga2Dc5S9+RLb3INR3mGk99TlgopkOGv
xgUNcwXmHUMMPBy5UW9qoLoAO8Y//IifL40ALy3HYwWX1t1GvmudB1LhFxoSNz457r2S9ikMq+m4
511uVgIkCx5+TCteDHKXqm+6xRP+tlfHxdgh5Ug7+MuVuOBTWWBbVx+joMEieZDHZS5/1QB8wtac
BZzu3ddZWlwVYbq6dwPuE5/fKXm2WItf8mLecJ58xzFor5ET81h770eeS85SUELCUT404Pi9HKSe
j200QRA0Ltude+fcgeCrFW2ZgyNBe/yXNPQ6UhlCSygglWgDdjPC8xSjqs2VGtAaWJBh55Rdzd8H
v3xQo1O0dB8WiI9taa9B0ckcdSRZ5fCJSrX5Rkb7jgx1a5MV5EkVqcEsv87tr5B8P70NY0SE6QIb
X+Y1rb9tekEnm+gN5rY6WQSzuHVI/H38rSJr8m4q61n00wYfJLbb/WJ+IhjPvTagiYVta+it2XKk
OoATX7DOw+WvlWsRIRQCXNJGc5GfZnqdpnP4X8yhoRfpITAsxrgL1pNM+RuP7anHt9aig+Vqmm5X
Ne6DqL/zVmu7baUBrhJwCBIX+QUycNmpBHA5YSijrQh/V34usJm5MQTQQerVLj8+3VwoCKvt4XoD
U2ozEmoX/wI5QTlJYCfXm/wx1pNTLPBovqxMZRitVwI4UtwECuGd+NO5bBsspX4fMzrlhC511Do7
iPKoK7Rzf1x8f9jPvtljkv5loSRKw4zMk/j/+PyRnH1ttInH+Efe3O9CyIcNmIlObVjePP58Y8TQ
oWNZnQoOabx6HMrGUBNLlwlONd9chiQ3pp3KdW/8g20i29JSy9K19OIHZ+KZ9J+EZ+P4BqBorLep
QHvUTl6NwFzgvObwdttKlZdagyvKWHg57eia+axlAjCoYIwNL32WjihuzFmD6K1/zn6/VM7nB09r
J93pgt+MfWjF+lENr8Q29KEl1gfdtHw7bKkXNewQVm2cL0650YaZdWnURsSwFIMGdEI49XlP5D7l
BuyUSpCQjq7N/5XhyXOUELD36DiU1OFi29XJQMzvx2uA389UTWSteAvhUQSG6Rx7qAe/snRrjh5e
QxQ/Cp7l9Fy6vM3jWTgCrzNQIhlVwl6ne6SMtv7J6cRDo3YQp6OhNY6CBF/wxMZpmqFKvqN1USn5
IV3tqZZbnmPwq3j/cZwe43a7P/k9pHMgqZZ3UMz80snoK9YNmybaKlYwI25ngpNsY9M3e/ZBdekd
36bGKT6tpM3zO5QmDodIDivPa+BGv/rkEpqWkGWtYt2rbXZ5rSfgWla63wOcFmUsYnFpzFKE5O08
rPOIl7/qLGOD0scAOD0lcc7ISVG4UfazV2b7aDafYLR9P9KgRF0LPZrQI6BlVbLg2fZm8zqSNuiQ
gumMVI3oYDnGKZWH0QJumJgw0sLK5Tk3EDZCNZ3a4O+OWg+gkViNNAFJC+RY5Li3xhbQf1pZsy1c
1vWjGprd8aR3PRqHgyQtfUagGA8qY68sR6LjaO/iWG3w//VGwvX2ntyOT1ndNM3/wopZJq8NpL7e
OiBYlFVgJ7l3fYwqBpNLD/X7UioAZvIhPqYdzDttiZr0wPhlNuNdCnea3PCG2v3WufWtf2sUGx8b
Vcew42jUSmlbrx08rV79cK0aINBZC4NeiwhDvnnZO4XPcUJSTW2Bg2ob6FzVM9cD89LWG9RtwhOZ
O72FQmAOp+OefVMad7Cva8UUDUoUEI0JCpkfPTcgKeMpSQa+UF6Q2rMl5bTuav2sD+SlCpXi0y27
ecrQAXCFslvvwx6cQy0uSDRIJLC++5DwXyN+/qXptjj3nHGE/cmB5McmswS+TsaujXvI0vZ0Fp9o
B3mSK0/jxnjg5Q5UvW6NLQ82MjadmL4WFxjz/2zyg4pZWqrgRph01qhzLlAhL2VNEKv7Uyph3n1z
T5vEans4od2eB+3rzA8WudaK7JwEHYvBbZmasXqscbeJwT6D4UXebOCuF1koFkOEtMxjHus/bgR1
zutDpuhdHmJDK2W03/9nTNk2beppQ3j/LHjPVJUd29H0ex0bbfBuIOB2T95eyWHM6mkWA/2Gzofu
0qX5mC3UGNn8zVFSwtmykL8b2+A/CtytSbDXx/TlaH24LBghygvAmA2vIxoJEgWNOXRVpuTuEgow
QU87gLVnqVgXgQyb51YNr92631d39UsAFoO1+yqdx40wC5wcUxWyJWs0dkbGncqpzA5pF0p6MdWt
3M3CjEomsIbPaKbTiBEz60PeusjM3J1kPHyHTjyFTGz4lwKh/CxhrOn+j3C2dxgrNxHkwD/lZHn/
Ec3GH+SqaRMQRXWc0FxZR5K08UfVCUUa3IgSVCMu7OuCEZPg8g7x2mxCMOoseP0hNQsGN0XvDFLK
y57onkGSAFAs2KcCUBQ0eiEgCO7cJ/DJ7EgMhxX5cIw9nvAg8pIZSHLWdIBLNA6uz8fB1kva+O26
e1iFjfqAwFrvzfgNuuVYp4ycaS1VEyohuxGzY7E0hHeDaGXOJfJ2/pl4TUyaHtkUUuWLEpX5vWK0
Sh1Ks95B5QgKEfxZ53cPAzjiCQGvvwRgAmO3mNkx/xeLCgS1FgVz6aLEXfp9gIh6ZMXi1ufxAZ//
uucV7/nU3hdmW07t/DCDim0CHOAaOSE1lTh8HYcHvgqZpdqWh3na1LSxQwstIPulmEI+UERkPsLW
QDPSI9Jxp+gxRQGiTkMuwMgSAhGkUaHH1Ke9riNesusuujSVUoy6bgZ39Bgyjn16rTklODECy39H
uwwsc6zuGSNY6edws3pETw1m2tgdTvRWKyksM914tukwp2Ua//cYOEWCZry8asFyMOJgPSaqEBGO
ttkg8QndOFmxYMwCnuQlzQ13xWzcmjgV3uHPUtw+Zs5GthmT9o0qpBkTPoYw6Uu6WgTJO605uy3o
mcHmtZWCUz7TqfRs4BjBfdYzUx2jkA9YX/+m0zpYVJrZHnWGAjg1y3MFKKBA9QxnCpkE5RPvBxI7
QtcfCpPHYonTB/lKxtQF1tXwPULn1yEkZfe8mCfg6UWhEgv+WhI+l4/CFbQQKJ1+/gcAk6UQ1Lyi
+uT5T77eYa23rTmHywCx7X2EXO+D4UU1/1Ct0tS2G2+heP/o9NBInXZYSL2frogfQcXbSSQ9a7w9
LpRnosoidJe4TQkFRoQKlqKeaHZ4NN/1HaJEGO3YK1bKt+8cI8T7iZJBe7vBOdlvAgfS+J7MGnN8
OsgzjrVGdtmXfyb9qQd81G5FoK4+UIJxrFqLVYN8SkmvA6cP5Db2vnW+klJAchuqJ+nrbvsibyg3
G7wCSinmeDMOCVIJmSdP97udfEqP/yxjLj3xu2+/Pm33hhfYkQfQ0yYf9avMtRj6dpLaANwkP4lU
Klm7fFNTx90+RI3jSJ89bS7adfg+mV60gmhILH94JQjuzpcYsSfNl8w2Hpvk7UKLW4BnGOS2zstx
cXBoNftZNLjLKkIdv/ifClTv+LnAmKlOeqgVemtveiDmLUD14tQbNS45DqoAevGdKPlKU86LQq/q
TzeKWCTnyiTtAxp90EFyrfqbZum+zoK+s6ugI0J6o6/Nrvq1rYBaCRAB9C3nBqmDKcOhpecyRVp5
59gvFJzbOZ+3K1ifSPjmk3CtQ6Md4hBrdeIdT8XvQZ16l4oM8pc7FvckS/rndA4G1Z3KIQddlgLs
pTJFp85rRlzdIwpEwoT2N9FtEdV81tmWVO7GiKxXL6EBvKZN8G3vubGQpR2d2xnXTfTjNS/nvkRe
s0D/jZ0TTPb8Hfeb8cz1H3f6bYr6TNQMOBax+8AdM+xUFYYshbqKuV5XMjX/BrhAOPLI6k+LIKTo
fnHL8meLE3hJ+D7qTY5cXwgz4mlIZ2HQdBytRaQDyWjqItD55bhI99JmdNDaX+gTRncqM+nlM8IQ
xmxI2XoJUXvtSbakNxxqlE+u61zyAIv3xrSnnoHetw8o3DiurhpjQKBbqTa8lvDis/XzDbLcQr8K
ZszGj9mzG22uh8i05FXGp3NQmFLyUn0KFFOUowzSfYR2DFthUjTpsV3DTlGsWOyPn21WpESrnoEb
VsoAfVZinCWrStEec1irXflDDwRIGQ6vZxY9uAXX7DsQD1otaSdh/XsWfsNZ8BcxP5PbbDvHS4Hw
ltkjU/Tc2zh1mlLghfYEAFXy4yLccu+0xyo11U3LAoGIIEKYvnuyuDUv2ihLakfVWWP43XppeVb3
e8CMIAE5h03UZAFvjkBiayUcabSfuD+JgRJngUgRFrgiNuYjjoutIYn5x9fecVFtCgQu2GlIiHfO
sUouQ/wEZrEYrk4nrbxMeULhREVyYJTY/Esv9qc87Jrv3Wb28w50POEyohmHkx4bf7Fo8zH/EFsa
BgwWkthNQCin58G/y+rmTCSrsOJllTDfOQ53APb09kQsdrkzEerb8x79Ci2evjajfJQZo1gyV9pO
krnZEu29lT7IvETcwktLiWZU1I1CjFZmdkfwEy1jVmyE4QTibScA1dFqGuiBNRykCv1ZUsjHawIr
zGaRj2UV6e5bYvEQnu8XzSJ9pGEDNsJh0iOoyuizAZQYqzOeA486xVaKungPHNfpK72+h6r4E2Tp
QlfNHOoBgZ/+a6+JCjp3anjbRvXxJBdQGpo3KCd0eTCyHJPcxUdggOP9+ds3rcp3ECJkdtUaGPUb
Bwjs4Mh5SXhrSSR8vzyzbwAg3g8L8hUEK+V4WSwoAmBcMUgva19OL09NVljG+/R14tvTUwV8Vp2x
kV1+Ytu6IAEsubVwWZ9vjzVrrtO0toqppnsKM8u8E6IXhHJO33E9ktggz+98xelRVSa+11ARLikp
bCV/Qlog84+n4meaDyI+fqWBOAskWn3JO7vPMN+ny7ta6/CQqXhIYXfNqXvkmC8gUcxZ/rSomjqA
+T6RZVLB4VcKivnuUlP3KIET2WLzVmLvddWE7Ka6uDevluJKI7g8HPHVMSOIOirbiJindOhIrDW6
3LZfF2LJGx56swiIxHQbhIUZPw+Eqci4jrPPdbHP1gHi+1JutNGKY7mMGgH4I5bp8WTCh9qVDFpW
6qgdWiFXyIEOCVTooy/WrQaBjw8QzrkMd6+euNlyxQJPqTnPtQObWLmZ4UF2B1F/mhxDP8uQXpT9
QzCfG2kv8JYC0Y9Ou/r2dBLCJlnRQ/kep9hGQpEyFKfIfMcPNtg7XhXoGHqp92zu3lHGngGiaEWZ
HTc7ujJX/suDRCwVzkuTBscIk4E7SAyOdP12i6JCI9EW6cowQrf0MzQ/s6DtqM6orKdPpINC0zXi
C1hb5SGzDTcOcZPFhU2XGnoLwgp5tjb2tuL+TlUb+fi2erzCn/Vel6Om+lb24vD6yGdvMD7e5uYz
iHL3GEBoBsLfBpS30qsA1yDuZ+zPcVN+61JvgVbFNYrdKBtMI9p3N4cnaz4NiPmLDiC47HzV9FAR
mv6pxH30XfeJWMs7AAYUATx7/5P1MpLd2D63sgaP6Pv2uF1ne+sMa90P/YGRNhMJuJtWxypBeFjD
c28eg0+5UUTF+ZFe0AXX9Rz3O5zOk1+D5oOsDnbRZ1/4tl1047JyIrXPBDn5MEYmnye3yrMX6Q7C
XskxHTLV7oLlJuPTIgzFvuIu5N2WVYAQR8l5RVviPOtLEymAZ5FdWBW9hASPdl1gYBa3elGnqI18
keRiUtfNP0nE674UqRAtDZyachIGvGxYe/4XsSkmjy9izec8QhNxhchlqyHOsg7V9bu45fLmwTNM
UCDHTcywB9yDKtsMbwFn4u0ggMgzLf8eALQrSrQBrxMYeDKI625fXnsp2S6Dvjs49xAL0gfoGjiQ
Lbz4JaX10HnxL554kAf887S9v6fcsuwWUy7MN+s4SohSSLMK8fkjwj3ZghMeFcBUrlVw9UkH0lB3
G9aShqHRjVLZzC3liWDwSDKQomcwqkdyPvyvcKOEx79+tIhh2bLyq9rXZT1H9Y/8RtWjaQT8arun
Dp0ZVYo/C7lKIaJps6ZyW7zOEjiDOy35sQhEhTIUn/mdWlF2vH91eiEu9p9GA2gvI7VwVM3QshsK
GEo2lN+Crby48b0YGfRfSj0OXiadpd+wLPXxQvl+Xz45L3fnk7gshg/ba/KiAmjS4auwn7ahh68D
hIlipvqZPbA7K8AyoQEUnJnujQN49TGrh1CHFTU1oSJRKp10UfhTFtblP+y1BAiEQE6SqfubUeWI
nbsh7R/9OGUI08/vhyhv/IjzgFLgxOAbUxru8JiLM1KorbzW0xt4E5YGIirT/ZQ4pqWDVcwnFRnO
7mLRY/ieHDTct5hKJczyGc4+LZ3MdoTuG+Ci0hU/bYFSqrJxM15WzCicuil+bUHo8I4sQryg+sX5
TaZBg7oEiRAhfhwmDbX/mefltPnbM1feeCuxYsKAAgGr+ES81sXhEaXzB3ck61ZCAcVv4ZKW9Hf7
8+gzd9DzZx3FW9CmhFQq/udO0BL+5opInLN8i0MgY2/nD5IBs1yeXnm0SAGaDLd7Ejvv95loaVzP
TmwZq98FP3U5XL3JYlqeHbASZa8JAws+xGowdotXqBDjkptipkKhkSJcqjDTY371NfRme1yMNRXQ
5FOqNq1Ph1Q5Uz2q+F5+q3SEEPf1koK/abNCXeOpjsAYAsxO4qNNLQja7gblDnmfd6Ug3FhvDIuS
aX58D6KC4Ec7ZUcTQq7JZwYdtmKjniFdWfc2gFNr6qGSYfE7QqHaUmFetRV57wG82Mej25h2o2xX
QJbBiw3UZEqVKcRAZ6TZ8S4TtOha1Rj5lgjEIJAyZWgKUYs7yAdMqFKDhNj142Pr35SPxfZZ0Yln
n/LuCXhS+RlkN3wybt8KN3peXVmu2hpD6dPOpxzAxtay+cVksd0aZMibhhbpOxrG4+/kYOf1XiKZ
U5Wg0V3tMi5lo5eO4xtBSukRrvsDOlyrqpvZoqFGQ8x6hpv4dgjQFIqU78WzCfex/msIMlT1PddU
k7usZhXeGwmsG7jdzITPAquvMCrgnYSY5dNm94mIXkUpsyUfXi28RYrvbFp5ZAzg9/RW/yb3xvc4
B28NqECxfCCM0DFqRMvyPm8d0LvMi8O3v/3kMUmhtMLb1+ZI2WpsVQ7yquGWr64AzehwDE3YxszE
aB2JLckT2pUkTYR0mIcrW1SwltwHKNgjYFIMp77wkKL62B47Ey7l2FJlRLY/onNHBFS/SdZCuvWR
Y5SVZvnNt10JBcWom3MNrwokobHD0YGYhJiz+c21P+cH46YGnYeb73k5qOnPnuiugI1XZDFW1FDW
5aDdA6glgFuGVbNeG8BhGskcyJYdKGr+Bzvz8Nz4PIYsyiJu6riGErYJ0yz+VkVt5n+fS/lP47JL
JWzMIPiWiAyqSE+oyCvagZ3/Wpw5J5aG9kG+ixLaEk/gfDQyML54c3gc/CaH9d33jViXk8L27pl2
Q5BtXnlBxgKP7Qa3Qk+Qez2MYGccsBOq1iDAbN2Rz2OK96UEPjuZi54Muhh1FZjYnCKaNwgNGFKu
awwpRwlt721sjCmOza9AG0uAqBlkSpXk25wHHnK52dYdAEBh8l1cpBYlbyRYhJv0siU6gv4r5xHP
7HVwW4brOfCbR88MCIVzRo9QskNpPvEIvECnp4Q/QgToyHPykxSljRYxKwUZEUhL5PPQKqvyDjsf
ssiLxSctzxgZC03k5+hesouNbzuG4J5RnDzcRs2PBYH7vVjPhVQ3WDOpj7RxealBgy1Ct+CCP7RD
eL1RIYWQ0NqPIHnEyw5tw1ZvJHjD9Xv/hIit4GO+GO5n0CJfaLqMChlw9UQBuKIJAaB9xRpt+/zJ
+XlSdQsTb14a2wDx1kjoaSp2kfuvI8tM64NTovoX5zRzG/db/x7rfCwm1ajhe0DBxZ0UvFxYjDYf
QZjaHQpBx2QD/SNstr73dy/cHLkbh/dUNIa0nqGSndboNI087QEP4GH+wRUGaW7BnwGsv7fRWufg
K6BqVubfwrnYTcGVs5HTlMJtahUiwSBi4s30pz6gniBSCppW/X7F6dB/OzaBSTZLJABAsnFDJrTT
HTk5C9B+METDfUHaZT/nVRBO+M6BAcbhchN4Nfz5LyAf9ieWkWRulhLaynK6oN6HeDPfmZ0YUKIg
sD66aIkrnUun8W9PTMw0oA9Di8x2xjPN6wSlzHzBRCRRhsR4QdDta53aTG2R5tf2WuaY2DqXLkE9
8vhQVYVOmKGCK6C2rcg+WOA7UEEA9yfuYpMfIta9YkN/7pU5nWlInYeThewyp4B3u5pPMSiclOCx
RlE3xIP/0eyyRKtviok2SlYh9EqovgyllyT8k0MHU/f7RsI+VQOlV2FAsIsq0aICK/8NSXTki0es
i6aVcxzRLB8I4VDpHTuQVSeuKjJcpXwM//GepQrPoSCymEBjV5x3W2a/fer96au7iqLFkcLcgAOr
6Hrx6RB0UTnoJmFNSII5M5RTXhKcD7IyebjfGojCmHCgXCEXGnNzPFq1l29y7qxMP/SN1NVyJJ9D
T7ZkPDOBYWJ8Cd8Ga5KKHggXsQFid0C8/lH1MRnJeylkiBRcJkXjBjXMJBF7VyM8Y68DhAGxIPb+
xg0MTHkm1wbh0xyWtSTNGS95z5HtD3QnHB2G9C3THblc9nzuoXJj96NTum5FfCz6oDpn38+WKBAg
6nmC3Lh5OlgUUlA31aT3CkrvT9q5zhYjMn07PSLstc0TBc651NzaLAPZWjesfEpM3akizWwNS7QE
VgqWnp6Fi/MQumuY/ya+bO401/za30WFAoUrEWaMCakRLEouSWQwOvI0JubdnuV59J6+oE52TemP
mkl0nlMebkeSNMmQiEAh+K5s0vH/pGwZDbuAPwpAie0ZnXhx9+VEQes1Bzlma1eMwlseTYQV+EQB
jOY9YUVXDILunptTISIbF+CDx36mFxYUJXvn7aaEYO2GEgWykQtzoJAWCV755MjQjOiUqDg6HVeu
WurvrSt3EpoM9kVb+o2otdYf8awAq2AWD26pm+A8dB6mUfchTQ/YnYGyLITJ0LAq4K8tJ+34ELRq
TSWDsxb3x+4oMKJIgui8Tc2TZQJTKJiLm/iZcBlIdQs2tlT3xJGEJxSC+vUKheC0PuA+2zERx+e0
TuARVJwk53/1hiFsw1oGkr7/esLMZGqWAp46b8Tj9c4mzp3f2h57tbIP+4H+UXIjsLW9JcYk3Oxr
qEIgUaEax23Ls2sj91V0WDNDxEGybjGAnNepsVl5czBDkL6ynlEjsBnBJx8Q5gRZg9CSHvjvyRCe
UAh5n3MW90/nyLHIi78OGZk5AD0LmNnBhWRd74beBnXgf6eMW0EnAh7mBlQ03Eir7FbSL+Ll6yZm
W4ix7IBA9IXY/lQgoC/JNcmF2VCQZkRG8nvBaE86yWxOt8/F+g+8ZuoKNC/lyqJMRbfO5fC3z0xV
w9acEFXqKwYX6ceKoeJl0f49sPihRRR6kBhnEGrwffkjrYdgaf70Gccerks6FcuwQPkt2eCydemu
8UayF+2HpNuG2tcYqF5LqvjCfue8O09G6eR0POjTuWfdLRF/DCHcHTEYZv3oi8oM5fNdOMeta+ic
hcEyCTKcMsT9XmyXP6G+KanzE0hsWX8nortz9t7wQwt0QGiL35AFwX7MxGrRY8ggYx92lQ91lfEJ
2AeiXgu2jIHjhAx+nOqz9dBlLhIXcWNMbQQnw9zq7P2jus971CaK2fFF3F0K1+G3U7fOrohh+n/i
TuZP7CpGQXaW4DdQFFpoDuriRzGaws1rallH4SngsanXBwxDkgfvBo0eVf1UNnQMBfZ9xj8ugLSY
2W4r/eDYCSqGoGUDhitXv2NSYVbC7J8WoMSOoLABaA0aebqgxmg8xlyiZP7IQqgGDHgicz7F6X7e
xwT54y/E9mmbHMjDZYNmroBMzE82S6Yb9qb8bQoFbsaTdzOTb+W26n0R5f6Am1AY79wPV/h3HDub
2ihu4snwszrOjcvM9p9RrlujOX/wEWxOuiOKwx6PJWzDqeFco7FjxWQow4DQMMNSj4FgC3glI6CB
tKhfR7/OA49qpPh9u2scjRhQW11DT41U50+UTI27j09Uc663uV71cEOI0K/3ptz3aNjrDjkki4T3
eQNL9Lex7Mam5uavxOB1A+fp3omqSPIaWv++PLTd1dgqAtGI5YSam412LxSFmyCWNHle3hpvJTWd
IGdWw/AF90uBWLE4mjGFxI2ppDhoGmcM2QNNh7psrQ6bE+Ls7yoiRn8ZX4WEh+a3VWLR1xsEbD7z
QwnCHm164zXSn3o1kwW7IMojMXEkz4VyuscdvjE7ScoaICZ3zshXstNuXXrBAbGt9MY4ih2BkpxV
tpfpBbVYzaDG0HSL+bJYPzXMswq2Jwst2I0isMsUh4oQ3uwCyuWJE84iuvIX/TwivqXG+pDMItIH
cAo9nhkotYKro+POySQKOWx8pAd5hn40WSjHAya9U1sjcfQE3I0Wqn8Jnu7jIVNefn2WDnmHktIq
OgCYauQDY1SE59wgdYIhoyzTBRo8OTfNqq1krLePxaKLvNmA+j0aTKvaAk8RlhJXn2iTw2wm81oA
ORoY4xkgEtkW5t7+Pi1qh9+57rROCJ9xtvvNx8C3QsJZpAksgYq2N65mw5pyq+1DwhScnSQ4rJym
d19nGF0gQeUD6RtguVHAYiI/hrfabFX46dhJ0U1FGkufIYU/rcZmX1Ho8iUjmUtdeh8LzgvBcaeg
b0DHyYu2Oxf1xfFmKjaxhioQ7lgtAUn0P/oE5ggkyFiVHea3F3LyKGvgTX/5vss/KmClBfcwo2Fd
nPSOVckW/1+nOyItCl5EEAAUohfzman/RTD6oCjo/ZE0SCT7oqQZiV+kVBvsZXDE9YHvvnPIAqrk
RINuXQ9aGMb0XxingUiqCl6tadoF0XYx/Yq3xELWDjPORo8VA83d9d2j8TO02+IJXjYloVElETvO
jFMiQ5tJGwCTGlJc+7oPzf37tM5memcLUzKS0goqH7lolpFbBHcEQxCBTDvLdMvbBs/0KknUplui
3y3nLuughU77OuaH1ULp4SJys3r4473PWUwYLhHOpfCZGJv81HWHG+GUtwlQD6VDrjlvuxLSdceT
yuWI+ILws0dpR1zg9S8BWRso3XAidpVZYzpqibeKDWajMOCg3JDtdvg09qVBXJ7DpHBVTdnKNiku
OibDV7ZCjJAuNkOmMYtmer80//MfYZb7DdF/I+7IISR9/Tnh03bjnuCsLQbn/RT0APbddBtSk6Mn
HrVpuPFtmi1wOLkdkVDAiABMSBbdnOjW8MttdiXO8/XkaJgMwKulMhjXkw1dNnUyawN4fiIG999B
YsbSnId2X9wqMOHK/onr55Q6OQ/jFikpFosMXeWCdG4+dsCcKQ0BDqFxBC9COZ7lJfTE01talrHf
FK51HOYhc/sUZpDTG7/sRm2TOd0m1mFQdokFWtKoi+AseQ7RP0v0qfkt/Sfh+2OtC1+glfesXpfg
M23XUbU/yAW9E2+QV/7q41aq0n4fxkgCbUOVMvyvkZ33dYGJjgAyABYVPPHW2rmmlv3IDunQVUFD
b6IwZhdNgJGa1pCL5UZpHgNuBkSvOW2J/Yyy9X6JxblUJmdKb3QqArjMDehNmZ3oYPZorIjq2Y+q
vEWTrkGga4GcvRkgzPuo6/erCKVq9y/U2lcAaCF9IFqycXHkaiNm5/lY72qUxUB7xTMC5bHIuHdq
Qr9RTECaz9BYFdth0Dw0HLPTNivfq1h1FRd5ZwEOjcHcxybm4kGcjMKR1RQDXiYrsb43W7zam0is
iKrc+hpDHBfpxoeBAWsG7aOCkE6hyzG/fsOtIhlpVV/ecctiJVnJfWYleNl2OwIMpJukNrjM1Ze0
2vTY2xhudO7JM1Ka7CykLLElEtJMPvYk86iNruK5H4I0xqO5dMZYLAYpnrXOmHn51nPYCM3uBgD+
JKVthv8oBiwZAZfwaTlxzBOqsAmHcnOzG4zjUsParHGr+LdsPToNQzHnneLkajqZd5ydbB636qge
aAYMr22acJrjyir6/iqBvqDHaJ68ctbMdCTG3Xdv+Vtn1OYcmAtDoUTRcPvK+OpxaMLJ/6q2IGNT
b9SbiJbQmm65QWMdcILrztWDkIiLtxV7ZrpjTHD9FkXvM94q2ZOINzQNYNPWgznK767h8XL8qFv2
l2ej0tTPxZlYU5iyHtpHIClVh9jDnnk1/pAtilSOVbXP7XQTshcBfHgGvd0xUnHzz52jtL7wkhu1
ReC9ctjXXl8VWg6tcc0K3iDV1OK2qi4zBoOSZLzmNxFFb8cXtzfSwjlzS21FaBtAg2hEwndl+o2T
PnRTSRPhBQsB/1DyogSFDJsLcRjGVHucdBhUPlaQsRVUyNQFcOE16xaEsbxFo75CWRF5znq3Nv7w
kQfKFbmcSTVcEDHeVgNGdGua6wIn4cQMpjor2gd/i8e2ifFxLvuqnJdlxd6h4KxmcK/mx+mYwRcj
FPKmBC2HGMPZi0DU8IuqPic4FiLdaNNpej3P6tdHn95fTsHwL7cc9v6mBhZ7Qa2O5Eg9amT161SN
zUjItz9BKGCY0MGmOmanxuzePvfYj44BEwKuc5nazYqBXy21J/Qkm3WidzTdCq4qLnsEaUxrfh1w
S0x+38Y5zJEuF8xpxEMQFSjALFLJpwAhs6mSUji9Q/wo99INUwNSusuvb6SEmsF68wosHGpdi3OY
39qO54kZEu445IgdZlAN9aC6W0KLeNrl+zV2biINOvmiSDQftyZSMde/9Ac2t3vury5M8Yfaajed
F0h1tJCv54PNV56RRFxDK9KShha2o8gKETuMzqN6slXKr2+D822iKoQOR6vRFzrFaQ4F+l+TUYY2
W+8avX18nrwQQGfo9baYVs7gc2e5ECNpK+ojYcernORLoFkWRQL7TmuwjIFH9Hwg6EBpdhGUd9QH
kyM96cH/UljHO7Vre+NW0EVrEOqphPgrqHXEgdmF/qm8b943ZnAXo0k4Qgkt+7UV5VcJ1tOqQ/mp
evyDGrdz5Tynl1hHJu+X8XLDWAKc+hBE5bwDF/QKBTBq6DJE+RDEO8/ucSgQTbkc7EMg4Dfl3CBa
eygfIhlyambnHLH0C5HV/e6qTQWgk2wamvn6AXdGYFOXWFJDrsooTeMrLjAJ8wEs7BkAsY6D8NHE
Tpnyj2HJcKA2m2TLzNctjKhS/FUo2/7EAg8Y3z249MGikTP1P0D7PxCM9eupR6vWuTMSgOjApBnw
+nSW9QHzcGsTlr7tFDqYKa09+NqQTjqEX/KvPPSmEiTOBmDsYzeu9Jk1Oiso8HxKUUgoUpJigMGH
cK58HCEd6qbWSQXztjoVy1lEGLK/cFFjhtCvvArJBKOzDxg5OK/WEuPZf63RuprMPtil4k9cYBTa
x32ul2uARjIRBKks+bUIEAM91KfdEgtHKr8qQmZ4D6Tqa9I0XXuvdFiFY6stBsb48scaitMQYBQf
AnSL2RLemYf9PuPd9HbPZ422IPsEdicNtPCvbks1+pzSCLJShNjvra2IBIIFHutqOlV9RX7DS/Iw
vENv8hOL4yJHTDZpfrwTSgn9o4WCyrcySHA8cOJTGfDo5YGqT+GDoZGzYl8pCXP9nWupBV8HeS0f
yseD+yEJwg4NhKC7RduspPvY9C1eumnOCF/E31wfvTsrFkPmSBlMriQJhuyU9RpbcrqESj9SnKna
DiyU01YromO1m4E1nPEZP5EJYX6H81oa84adEs7lxfnHAb6TOrx/fptFnfP+41ppXR62FxS6SR+R
2QScddZlPu1/Qde7W/ecGJHkf1J+n39hrNDPy1pHbzF5RqjIBumjlJGJJgZAJ0Fdg2jWKOU0wyqp
mjvNMcN08DT0KIcK3OhDO1RYDtoJ1LpvEPAkaLrBp8N3bSAQ94vxjhXC+tl/FbmgeZf1WVw3MW0H
kDryiKzXMgvqR/6GUVt0KOpCSptcLai3QwGq+aJaI5SDB3BSn4JPLBG0mfy+/Bvjj1CRfRXGMJdb
ek1EBJRj+A/+fhq0+Q1x6p+QH3yBsF6k9HyxVykkY4zVLPQgsjfck74uQhisb6qgyfNxYzUNbxcp
od+7/LDZQFq2srqGQ6VkFE1zS4TmuCee2urH95JzplpI7rhwHZUMNgA2xp2Wdp1Ojgy/9+1FURpT
JLA3EMDT5PICvLlMbDIXJ8Ul81URlYxGK+CCEu8HOWd61e5xWSZ62ykpO0DaSgkYGXBSqz/Yi1sw
09Gev1fpeJktdLDgjXyqD1AfsPn04GK5C8pSucKcL3bNivQ3GsBG+KxFb6x30NMtXqMROavM5LyU
lpEQYIC9YcYnjhJEfy6hjV6Urjh9VdI10koVK4AOHKrAnyV/PkXj+mIkqtK0cSHhSx5NuqDUnPzW
kubfWmsXBvhmVSWJcvkJG8Bn0ysIgD6IhgqKLdNcw/vL1Ku0yNNwLrSVUKg1M/dqAFCh5dzlaphn
EJ1JyvNTiK05xTBAO9uga9KnvZwPFb2WduDhlvcAzkjzCVp9GFfKk5fVudMXdTP9iauHtm7BbLBt
8E+fvzqnrl4hfhlf66e+WMk7TMJqo63nivzh0LV3S9F+dJVT2hsYm5arl10al3iDs+e6aZKQ7GJK
A2FZj/AToIFQHPkl5OW4Mjdc9WWP42BuIGcnNAnPAxkTWTcXq3NujL7eWEkC85hy4a/RK7iyTH5v
pluwdgwKZH7hDOJpY5Pfm0+rFstwTzBlxP63D02yAcBB6FX1CiPVVOTAF+J8Z82ZyBZaB+Fl0ueE
rm2T5cjfiHQKI2FUylvSvBEYq+6zFCLmMH9u51xs4ZVwXD32oy747/OIBnjxSMWIPIBHUzwsNplt
WKWBfKsiK0PlUHqop+4IlJBPShUaRAZfgHgF6UDXKPpxtM2tcpPQxeNBSjFHJfH7PRc2R/8j/Fm+
3oUVnLGXEBhrXMfTQN7gjtXhVPAypT47qMZT9i7Nf56hlks/H3BjpTCy0zagWhz5myvO7jAE/C0y
FUcSrWh0m/15VuZFhPqlogRpQonZX+bAyO5ki71KzMm8EKt2+RczcjyCWXx0bjnl/hKl41UrAvXG
Q74bMaT7NcXZALcSHG8c2pfYvxmBZ6eFu/Ih513gtcpg0OxaW8WEmDBJlInkDxJim95aj6yaWmbY
v1yweV4HUjh1h4S1HICcPMPfUrUP8kOnCX0lFa4/7egsW6c+mNoyrZ2MpMGjmarvYsExZyyvqAQ/
wZ5yVGk1ayw45jgMFjn/Cb9B/juqftsGgawsKNIund5pzaxxHutaWcuLqoS2oUM01hORQDqLlOin
gve6ugsQ5uo1xYhN0zrquYo3uTiD44eBqvEFwXXRrMwDCgJIohsMo1xsIq8iato+dJVIlde2QCSi
kS1ZPOCJO2B1kgKGDjPOv+qVGe9JM7n/h96wHMwyhh5mGcmNxQxUJsbe1uSVp5UAHBwhbeRSdx/6
PD0B/uz1X74w8bYTW/gB/xqBQOvEMQCPTHOy8xl59Dq5kTCHx/G/UnuzvsmOhVrL9u+/TAz32EhF
vzT5v/DK4JHD+EUWq0LUtaoLdmvsfyESm99f+RAr2lop30xZyn41H7HK5PZ6KZQKGZrtbYFiUUM4
qglcowtZ3a9zl9YMkxw3gT6w0XIda7yFmBwaUMNl90NHlOPdrW6K696DAkkDD0+a1sTPrZxd3cDp
A809j2K7vV+jzk9ar1BMvqNBoQI2g8Na+RgfxiWjg/yTpshLPH0X5Kn6ysiqp0oYiInnrAJPPNDY
DcPCJqw3/+vrGWOz9Pe0EbpaUSWUO2gA3okScBsSPj3UiGib0kHOtD+QqXe/Etr7OH2D5XdSUFe9
blq0g6B01wFcXG3/w7C2f/FMDuNl8ChWkIFijn+lixk2jbdUOcHbPZFzUZnvouyZsVOOcZmgMFdX
E3PSFDNFwrcdeIT8Jx9/VcRsCAvgSbzq8o7BHeTUlGhgKWgZRnxBt/hudYQoU+Nw0G94bHmdH7L7
gBOXZFPk3TJP1bvgnXa6YbEuLpz19VV9iPwrfCATQ9GyI5mg5pGdXfsAeBsVmTjvJODnWWacauW7
c9tv8Jw2QBBp8sF8NJxT0w9YDw6P86cg+kKZChyeRsd8T6V2S0u5JmLwmKfO/ouuGF+6m887BBPX
kC7WrrYvIqW02ExOWqjZkhROMOGmyvgguS3QMfiieMXYwNIfp9IwOhYKiSvHGpd7rI8YQzf+CY2i
KtkHVOIyXAsuSEaVfy57WpFnQT8xfafWSLBdJ5Ymtmq4CJlGbdw+JTFQHvrB7CA57IJom74n6mJ4
qJglrslHPH+YC0sRsdoQ9bZHNSzQZzJQ2pjKATAdTTjo+g/SRX9kWSD7L7CMWgLVfelcaVtHe18F
ZGl9wr2YMQ4YJdLcdLWucvQnkJZxvRXvybmbzk7fQ1znnXj4uXWfF90NLCsBk8+VA2E1hn/5JlCe
jmlo2P86jhJLEHmaxNX5qbrrCIfIiBCe1mrzcCZohlUTjHYlV9akFf5Qiv3b9mI1I5WOYLC6EYYM
2hmDljObq18uNhs10kCnF4qDMV150KSZXFRld6fqxyPoqHwntC+wyNxA3dTUVg+KiWvdpRurBgb2
0ejoiO1fp4K1cCO2tHrb+axrLbVgjajNoRViplbuFde8zVT0XEMAOzc5xnhE2nwC3fIqmDkJpetb
wapz6+lJX7JZ3Ssph3L4683f8vDeFOjpiAZLkGASk9QQkxeDvn+b5xIngSQFi56hC+8388nhylbx
3C61KvMdYsiG9vDOoUWZQ3mGDiyq351dkKaqCGm3xBrZDnjEhmZx47BzjzJ/a1ixTKJ5KYX6pkPM
HJ7K0OhA4gzmHtpxU3/PlJsNAD3VDCG2GpLt3//XhFMy+QDg/BolSXMyNHXQPX+nXkbz3085pOYY
mKDWArHRRiqEr68rjvuSwfC6o0l3fxthiIYrzcyHc/Zk1WQyoOP2kprbB5K4U2esTdthbvUWajQR
5YWxZWQuqXzKoq+RUfC03sR422tXAIa4IsyDuEbJZYVJGGplFbtuAagJxR0eGa/yScK3Mg1xj8BN
sBn27rErzNbaI1jHI2QcueIt44MvKnGZpjlPP0/ycktRdXwRNg9YAUxdpo3M6ohnEp1oyWz42siA
3137Fl6OAvu3VkgD5V0+rINX4clN+CE66hn0tkMvGCILp4HZQfAnyBxr3YQFeOIakRW+cFOP2O3u
QsyixE1nMtZeIVxCNWs+D23b79rCKnNv+UYvykRYnG8Xt0wQtY3SprbfuVbKaHwjx3Xjh5r+L+wT
Erg0eQFYcuvDPqW4aPxSiWTU3gZpqUx3+9h/bmESwyx6g/wSKzUmOx5XyxYr3jAXy4sJ6ov4UR5W
Xrm0Fky2JIsIhJ8osR+P8fm8uiF0og7GhKkQ6iuWJBLuQmz3SWvRp4ce/0fWyT6RYqY7lzjbupND
eXfeL+vVhspUVYBurilcWGUEdx3nLp26BbWqFIew56+Elzr03Ph5hRC7vGh+BXNUdeqIGYAKQZAd
//JFqCnv/ZxEa6H2K2Z6iM8TNLesIMoKmcFQFoJgt6A3XuuHWCuLAETnHbB6Ki8R4psG/X+0isFE
WNv8uj865PqPMhTiYFt8GPdI4ZUHl1JxvPorTX4dm7HFqprb+q3jszSNDvgpuoZMwZEXXo0tBFNZ
Dfd5Uf363DPnAq5vjq3vq7sdzIsRIFhKA3LH3n4WKGqG/orWVyeyUeY1TFWJku56IN8QX0OPIy9/
gygqTtmAX5zK5Qwv8E1Jyeqo6L2i1E4wtihHLDRKZuG8tkCuk/F8xzVDWRu0jgQzhAogEbDnwYa8
vCB8YJPpkhKcH7HMhvuWg7XzjjPNM1dr0J1KTcOZpqGsYmoQ4fteDj4D637UVTHOoAHjKSjcfcPi
xXEqeK69sB9r5/s9KwnoFM1PDS+yQXpjdvV4LwAsXmb+C30QxMcdtM9BJ+3Iht5EoE3hFlUvkdDv
cIUMD3UY63zfnSXp681VYv7bhlPok6gJtG3XrzZzcJy1/jEjx85/3RfdJr+RyMpFBwyk586xDqnP
WlYbO9j/xBaVpbMR8CtTNzrRu7Yp8H5WLfW+FJgX2aP+cCo2PQodzkmGz6nHNyTdfYg4Q6TyVmae
Wn4pgPQ5q8ifAe3O1FCkcObcUChfLZ88YhkRZZBR9XrJDSxN0xD4qr/+owT8dG8IZxFoUaYJ1OAe
j8gMEyNuBT5vO2t0JawcTT4k8Tipzv65EGYqDKYyRwJzp3j5Jpk9QK9U0MQ3g2oNhvoWvrM+Vi3D
sAAvVHDRZ9a1ms2eY2vFm5oAhf3QY3wWjnl0brBzK04oFcI/iJFKkt/KJZ+oCPusB1jX8moIRQBT
2tYKtW9T1BvJHmIbyXr53YaAWfjwEIhCaIuWkIHH1oRV7+1CBbjMYgLevnqlEjgHA8j89JM77ca7
flGM5vjJUPUuT4AoAY1asiSaBlRARaElDW1j6Ppvy95dMBtcKb3avVVkwJn8FEzspwoxVneD7XHf
Vo759/ZTbyTpREd3iBV1W0Kd0tfWWBem2IiAxoI4Pnp8UuNGCIMR/9Amh7GKwX6c5F8wOQtVUCGK
aC0ofHHmXQU55o3gZqzqLUZzoTamts9jnaHD2b7/mH8gZFUsf17LXz/rZlYtR5zbVhUrYU5+RhkW
wc4sPSZnSWgQZpZ0tTiwH24fprDnL0+xCKTUsxqKMoPc4MwQ3vITEXNMC+M61CxaPlBnL4WRo57I
+xmAXy4BvLmyWMHQiNEqGgrfZ1LCpcCrR6tjbg3JbcHtNM/LxZjmq0woXZXMnoQ7OrZAjGWTcWLH
N7S/HcpBon+WPCHuEm6QZ376eEmcGAVGVC9rCuMwNTbS5D88OPGH4Uk4B7utBTo7AUHQ+LrUmFAz
X0aNwfWyXPM4BfdRagrqKU3AzGSs58yejXH0U2Mh3uiPhvCybGwjML6BRBdFdy17Ccq3G2N69UtF
WdJsk52G12xL9GX8ZUHWpDVTFVQgndy5FlATl/GtWFH3ae4WNZOQl6xOufJl8ruWdpbnld5p4D1z
4Y253O+kc6Zz/43lwX6tpIlHRo5MiBmQRHBwCG3+Xq7sYq35Qpu+gZ0wQooj/GDr0GckYjH4xCVn
F3P+6xsFkJMduq2Npq3WodsC33nngSMSHNk2dZhGrndSVghTpggKl5GxxKUnwfYODYPiORtjL7lr
BPz4ZnCNzJoTxwuyPtWPhbmdxQ4MYb3LLdsVLPSDTLvKlTIfpik8B+FP7PcwFtkIhM4t3eZiLm9y
dwcnG0pFvxGV7aXL3zebtBgfMij4/4YL4xkdyI1oBPceW3mg9tLmIRtxa81OLX+05zpSxXmPViVC
tdHjJ2cur+bMz22NwfGsAiGdbgBZfZeI8CwY5TGMKF1eawkfd3Q4Yfud6ddJezkRnhjMT66U9tgw
ahRpGQ06hg/Vjm1widJ0lr6UpxLpqUB96Kgo0uUhCXT6GuuucT54BpeGTSKd5oBYxMi8mBw6dH8W
c9lIvAnJvBOn2V+GEu2E2+PYjhRMx4WDIx6OEsObjazwnbQg62OgZMVUMYaN/vEUvMAIs6xADdvI
219xr+JFLEAhEt2cvjwgRPysgtowrbsRMumIILpHGMzsXrfotzDl/FHPE1paWolybbaAI8t4TbDl
EMJxw12FH54d5rAnOXbrKIgkH61BOu4/Nn80VaYy82e4D5lRv36GNY3CpKrPs4jMUfgW0C2thvou
tm0bYeLihxnsm3kc6/f2z+Kq1jS2XyO1Pgh0vZoGN9Z/bJUnsZAL2y0sr8PR4G8gVQO3tH78XQWp
lMpTFpCFs9mfO0rkTsTctVhjdPxQmMnSGFA+tbDyMvta+tXJJU65x1UEuUAyzotNAUbR97idmQsr
fNrvoGCt4uLq15zNmTXEoroYr25kAHFGvV3MBngf3KGrsBUpkPqL0AqMQDbmF6hQhbaCLmuDI0y8
JaZ4FWkuc3oM2Q2PqZV2leTDlV45PXmlU8cHlzd0TdA1GLhJken7H2Q0edsu1lWmKrZF3ldUzetU
brbHOVYBm//PGxBDgX3VVy2+ytiBCm5ZOT1h1fTLDwt9hizuFIPbdsK8tTokJgwPymLuvruOokjc
dXbwMTnn4KXXrnv30yLSgS23ckj9MdmMUSa6GDIu6CawWH4dJuakq5HvI9tVNBe+UiaU18hQHlzI
pdKSPh5USvwFlPuHCXTs6UWsBrjj43+PaLVIJs1tADDQQCr/x9Xjlb9HomJ/kuZrvEE077XrylK/
8Rdsjl1cjOSiYfmFFWcu649GVmRljNd0cdG9kWRu6kVdlHK6YAZ5OACSoMX7MZyxSjy7PixrBxGe
jGLo73D77JUhnBcwR9uv4FhDO9i1bowwoWm1GJCQ/QCZdrlgGj8HjYz+RDBQEAZ1g4bjYvlRwcjG
tFEQAncoa3umr54GWC2hCjBkskpjwvgcsk5SEgr8z3eLQIINN7sgpoQvkPbtRyiMZFUXMcRKcfCY
+AotwKHLPRYq7Re+74ZZ3M2PMoglOsS0ZJuibY28vt8aUKioI6mrU9kr0S06uZcZUw3LUmvyxhfY
aRkM1t944Gdyb1ldnrQ9iZACBz/kK4U99ECcAEXMA0eBdV41Ih3WrlSbrSiqdb7VPWZF5Vwf3K6u
chhhN9w3aihtpWqeE2+vqz69SFBW+31MnTHGZpynGoHup9tHtWeGKoEdEUSGBs9hD3H/8KJqi2t9
tGmoYohB929UUmGRUQvfH6A+6nMJY8ywwHROmBBl/AhAVhwogbgjLY49bX/f95ZkFJysVG22VC6v
cP+B6juxh+rY4CflZRQMSU1bBEH7sG0h13VaURo/teTEtQu0j2ei7lHo3iwy8BndJF96auGvtZEW
Vdse2jlryjuucJhWKFXXyiwb29la5zyZHExUaENiqhfj6DLdAM/bH5Q03qLvcYChqns/Uz7roPcN
wfW46+qCQRZD+D0idQd84/52Ybjqz7xnbb0Zy1nt2QQEpC9A4kJpUIqHmA+/QzNdgDhNC5d2Vjgz
EysyDkrrgjnZO8Tw18O1OwKJHzEwAmiUF3yVh9EZQ3VciYzUMYVvpTZRgKr5rgm9Yv8QDh6PxHst
6AYrbdfNHpPP3Hs82gP1LzDGcUbljz1akpgG49qrVlvuwDBROglWdMBNP2XbTNmjOgbDz7+AjSD+
Ajh57NhuCDWTghOOYUZyGg+X7vCAu04cH+fbXdCrVm1ZWocmicapU4eXTi/x5XwheA//HOkd7QWj
oMT0MQAR6UwBRNcvkFv5lB0XQEAswCrg03SGWUzgHHimhx/cy7JOgBlm/T1Pvyn+4M8GGajjEIdF
ptBeImlMvhqhBFgo8Xs+uDyWsHrNyO0inZAxIzXP7E+/e0QRPz2ouYkOPgKWPa7Tc8He+el2urGX
xV7ctJocxlSs7YZ/gD/AxyiGcbfQ8kl71zkMkIa5o7IpdfEdo504cAIBNTCKbRaNW5xOs9Xgs5+y
5yXN+JoRdsTytrNMK26m3KcEr5UpeBIe8xHHl66wrBWGh3wqe/WvscElFbpmGdWSIg9AUt64kMEl
kf5lLI8Bhym8ucraPJShs84nwencJkguv9N6gIj5jrXR+YB5aCeRM7nn7t2b2F/X4kUoY6DApbha
3L4F8N7DoDcyZzo5djXB9kMPAnG0BEXLCARDoLyjRW9eIIXQU3oisBlJddvYAX3BBOPEZAdCDD22
ugx7L9jYkKBQfMSstOUrCdmiGicYqeCV7yNCr/cG6isyqX32I3KFOu32Hmbj4dJrEycGxI759rUr
fNIhtVFB34qLWS0hZaA1/DQE085cdNgrHLDdeWZjZsAciGuR1aAl2lAGJ1o5d5BQLImSA/SOpIZG
rM4pO85D8mw8z9sG4l1b2N1jKCrQk6RjaEP6Rzro5OwT3LfOJoVR5vHv6nCx73wknLHPu0/fL3+K
A27GCtdGi+RyCRFhpA5y0V1Ewo8n6lrxSqwKXNgvy4OKXQSn4GazcyBh9PQOFIQRe5z7xlXC+udl
k/kZ37K1ebY7Cabd77imas4axZv9Uj3jx9oY4ZweP39oNJVWiBa/gOSaXiWklIseJ/iqvTn5mcSh
+sj2CTRkg+PUqSJGYd67uVwuj+n39Zy2fqw3JTUSVG3mUOnb7vVHhi/6WlA7mA9SQwdvHYDYqw2D
moxm+V72swD0MsIqG5hgtmDjG5oZ6agdjEkTZ28XiKO5aIQG6tPjYMdu0U0/sMfuRa65YcUXMf+4
ZBtq6gIKqPU4ddZVBogEoFb8gTtHOji4y6oJxBynjfn65rHDjvWPz38iz1NeWJ0gYlMnvNLYbXBw
GCD3U/WhCUTaB+FctJ12tguZK2+Ug2aBiOaV6wnEwMYSDyo3Lev+G/E+AfHh979mQWmpU3vfCM0L
xEhPJSWnKOGwap4/De66oYF2LVFnu9APCgZ4VaVPFLmny1Bq8BeavsgebEh00tj+IIT7rCWYKFo3
3zXzs3hf16YNAknkKg76SnEwS4ywAqapZXYsXZ5zc987bGoj80Zl9IQ2iPSsWZGhN77HuSG7dH2q
sMWGnYf6NoQUZqQYzZUVTvvY1GicKnnaLkzqJVEtCqJbnzAQcs77QhuAHV+1kRGIps1mYbhf8wqy
EIRMdaBRjBsXTvRIbI78LrkN1S8Ff/YpOrsVWh0N2suAtvk0ojADcPNvYsK/5PyNAVOAZVNLndDz
JO2wS3wyUJ1IzMRy+eHGtdZ4NYaFxTZLngLtzeVlGFK7FblHX9Xa7UdKdPQ8lIiVLcVSrLrvdvjA
q6QNAjRgXAhfdBY4gdqARc0c3Px+7IEkCsFY3lgUA3mGXBjn7EnwH4yMJDu2ZDqijS3HOvLjrUyS
Y1E1iCHb9SF/e8fhTT/Q34gg8pUuE9fLMwDSMZA+vu2u/AfcVlanJBjuw8h2u/SigH4F0wS5XKWm
szDSMce1+eaGOp/J9JcSp9Cou3tWpdq9Vvu+f11mm9zFd57nhb7nOUtBIM4GVNatBlhlVN2osFPI
7x4grM6k9c6KzBj8/NVB4ZzVhbAh1rHna5xx5zQW/246/zLxdcD9kHxEYmANzs8B6MuMp5ibjaFi
eSSohnKXlM2kx7cUJiQKdye8O9bY6M9lj25TLwZERlJfowLRafYBPL4cmHpJunadHQHURIFMvHsk
nuL8lzSzX9FLLh1EBBjbMXnHXwuSnBHv6qSYqQcRPpZsM3DWd09+KG3XXy49zhAepd9inV2mgYd5
rLb5K6uKKM5fgikCX5m7ms3JI+vr8ZtH0C5AcgxJggNCCmmjKGfEJlPioaTkwRIlK0asNQqE7gpd
EKtI0Qt94beA/tVOmvaBriQdirrJgjNJOvo7iBqGpuxsX1KTXxOAy7UNgM109KiEHhF00rLQ21cV
6B4ZmxODuH3q1FoRcnOeZyi8PgAg04JNdLQkwXWTWii57lt4nEWB7u2EFeMTLlbs6vM9SZ1AZH9u
bMtC7cRed8Wb1lhcMZ+pO2nMyi5HFBCi+7K8+1HvqPFKZd/qxoxfzAiIOrS0gqfxVTx5DqFmegaq
4lKvqkY2lpPMqIrPJ+ir3dH5IFhgtwZCdkawhI3lZV49L0pXhpzWThPxzdGWdxH/DyQkLZUvBctD
CPtm/NZBaNu/ZuQe7EzezSUvXdDmkVmU3+EyBStPLaWSwDWby3Iq+8MR432m+eh+E93OlJFUGnah
tkmpA0NJfcE+j61trHhWYzfDFHvjbYW4UU218esq/U1+peX7YN3s5a8V61QguJc78ufCzpWvFCIW
G6UeoRZGynJtvr1WcGhD8dVV26zR+Gi+WwXhsNOOeq8SxkgwvClfNmeKAWkvyZ6TYKuBnsW4Zx89
3SsQcyG9ptdew9svYx3ICE/UiNAKOLaqRGjayX/rA2OOZ05p6DT1CFYCwtCFDeuCszDFF0WiaKRE
2HgFMeYXegXEtiY9OiQqKw+sCYMednQFEfgzaMkSUaId0E5NPxpgmqPxZctw3w7dUwqyfmjVhlPT
R5gszy7zSGXD3sfg7UX71Yw83zEDaJKosIS6y1bkb2sMcXe/gcUvYMpi9Qtb8h3s5HRJzbIHjqVX
T/jXn4xvex87PSApG5bpvCswnjnx7M9o4bCk6ifSocfumGyvu432Zg2I8PZws5WIcro00WVk7sAG
xkSuKc6jM7lqUv5xSIb24frhDB3nVhFJeP1XIIBk0EaIYUaVfYGl0bAiJUYg2VCRWEH07RHNwjoL
6fQtq/dUgTYiqRox+GBq29sU8mmcJfbJnXWbOZigQa9sO87O2HNNlQZwD3207Cvu5n52TzN/UvHt
d8U1LEMuRF9BkhUMUhdneovncTGi8SOCWWpKQbA50mTlvqw9KHK1puw09dqNbZYdte0PPTeT4o2g
cgVVUxlFy2rKpKbzlv34PL+K6Urs0ct+VLsS6H6Q5Od7y/VXtRkPrv6YF4FlKvw1IJodoIoahknN
pAsh7jXqjb6Div7s7TgwIAcG1UAaGrV3Gq10CM8DdHBszNKlsLhqOLqavUkximPYGDmzcBK7I6gm
xJG+11WsLbLelr47NI0aBD6r0jJOL3+W7usBzhEYpZQcFe+kEb9e2cU9S1KWov22tbMOFR2RnrT7
4GKanpgH91z+GLOuJHbcWQSzQGrTw0Ckm1/j+2qdsPVY/TlAZlQakF2CC34VVcLhjMnHi/Uu3awW
HGvE12gFsweFZNWrfCnMQYrrwuecQBo+6+YVlcW/pLHmEX+mIBCvn54tC29DF/gNdwVBmsICpiIt
MEUGcbbgFABYEymtDwor+fE1XucpL1bMqco07SOYKWkI2dFoya+mluP8C8cPBfq8u6PttydrSUDA
8XG9eIAWmvENF0ZDGXF8iKbsX7jVZiZijfNdpePRVGHHenXNR6yoXrqvPZQwHcZnnt0kJdpKIhMd
oy1JF32PUCdfbuqttFEPODVgkOoSyYkQA5q2FfpzhN07CrUsojdELpWstffg93mZvn3qbINqdUsy
RTH2kQYfwIivuvXA32YvyprzEndNIZVSkSonHcl23znOlut2xl9RU6OMnMPtYYYH3t+x/QC1BpqO
4EJZNWC7CByDraFsqCmIx+MwuuXhIvqm0kRcmjtR/qYd5V03RW02+kAI8GLdGVYCJLovwGuVKAFX
Q0OQH2mDeUC0ev2ObqPEPcGrrTie+MwUoPM39vk2RPCRF/DJ/tgKOnHYlLv1r7VzxvND/bOyBgxs
bcFd1IP6kDL5IAzLBBH8Hqaj0KP+92kuUV2uyZpODZ0osC+0obdQSRxQ1GjInNv2V1SVkFn8v9Sb
LYV+rB/Dbcpe+/l3WFNTE1mErS3eKhEhU8OOWYVgG7gF5gYsyC1+0p7qEdzGknWTrCNY/GSzz8Nk
QEWd4kz+ZA7ZsMw4tYPd5aQktd6o7C1G4sFCJNKiJD3mSUWvu2SxGrM8+kzlCBm4gUbTFl0WQmj/
QkeO0LThEz3o4ueimIQdjNs85rVvA1nRyuaAdvx4D4WjVJzoltdK3lVA8cL1D81eO4AWfAAcREGN
6N7ihwPnI/nOD6GzLgUR1asfrhQdfvEqv8q4R2tVH3K2nKPdBxXYmoQ/Q2HGyXllV4G6E59/77Zj
jnunI5JvbpY47UgmxLgFsc7zaQmyyDu16XRtz83yB1naXv5hmu1VCuLWZEzcEWebwEp3Cx3t+6ce
uM45ga8oSK06cR1iPmqzMv1PUT9Sqa9bWv2c0W7adO7uNLtfuO+hCe0GynPHnc+8iBJevhOuTvVO
gRHX+FGcPyI3KZeRh8qXvYDeU78AEwXx6Px5J6ZNNDfjCn1+Ir1qyLJ0ygGosU49LlteciJRJMiG
Gmt/Pcowq6t5ApgliQplKGJIqIVgFVSNym34rlZZM7s1eIgBu86jf7TVoxyQyvDukVh5qgaygn9J
3QTRksL6lNG6w7SG/ewoJb5gAlw480l1CY7wkHE80AwD7ztT0nvHG9iKqikNYPo8CEdsS3DV44cI
39nvLmCG1qWLDZRLhsKeapdRDZIHLnsj+XHUQOkPO23GE8wV07OUDfKEUtJrJVqCJLsG8HztlLjY
FKcUQxq769W4HmxmJ1yqt4Dl/EaNWUlwMHX/KjItHpdW+adV8wM0q9dfUcobF0haxnVPwTZVCVZO
pLJc9SGcQnuiiZ/YppavvLKgDKi+kSN3vnmSzpCnAxsWCux9ceF32GT4ke3uef3bVO/BzUkdBJWw
KaRJHjlFDdHgZdKBdrDydIIeb0bwnQB/eoZbx+Go22waxDPk1GKnfRggJTUpNgSdLPDmU30AC4c4
uPUxYxreploMNaECyhIhDBJ3k7vKIgiNqLvwLAt4KVe18/ym+WuSbzkQ/HRyyAAPYecykvRzidWd
qcuRmqAg8walrHibcUHNpdGrhJELs75IAwZ2uWjb3IZBistis48qmjNTKKwPXzm9igMZbJRJBRUn
tPj66VEG1LrjAO8vuSMVqifohT/IV8YKS5Lwb5NzbJ3GDMMsuJQ6mhr970DoR8fveX81Hy7xIDOC
4QFjN7Q9oyvl0wBWL82Li8RYhE+cYXj1eFPIk8gEJ46B5ysOaP7H3sgXST5YhisDuAzaHkBrKkr3
8765qjoQ31ICc9CKoshl/Vrbnc3ho9Iu+agDgv8YBqUiaR9IUsQVGaotKLbCs4SmwKK4qCMQpK89
BPI/ytP2g5TQtpfHhL8ex3fKuXjYzx6/HOHKvRpuANSGGogF1hbxtUDG7wJE8JEQmstVaWmq9L1Z
r4k0F/xEhpLp+u2EFY/fy2SBp6iebv3Xe79SbFQEfrkWZ/1jx/BzLAU/bIrrsNQPqc30wOmd+VxQ
5QG9QEW1lQxqta/eU3HktlfSShoQnSFfaAr00m/LVZNY/rMT4n/uTf0yfH8FwIJ2D8xQzMrL/Ghe
Cgh2sp8MNJKJppC73oAiM3GdYa4L6eu4LumpzTpFy5yOnkxcRK3u5oeJoAkUfi/58MBWyz98k2cw
kT/JrpRw1c6baTxqhM0YZQ9G4jp56alkctw9cBB01GfR/cmPqiNG/JkOAtd4wOxtczrgVpQ7LiKc
qWD4ey0Qeo8+Wepa8c9aEiJ3eWZRkkihPeNUl6kLsEhS4RTq/8+yicARfq1r21JdjuNG+TRu/vN2
XCeBouD8TjWv5GhQVRrT+mdAHjU1fGLjuMVDPvmbn4Q2EE8v5Yt3UXQ6vfEi20u9tNwdvBhkVhKz
axqKSixB9d5Br5KqBjf8d53nJChPSn+aM2F6J8TRx4EZi4jHXUjVqcy4zFfbEMX5uvugevELjzE0
5/mpg19a2iWq7WzxH/xyFeW4Kn7v6Y/vdZ8XdL6SbO71NlOp8tzwXeDvIbOMpkEUI0CSkVrqT+bT
AIyN8d+sEm4EO5RwVGO1K/Yw3dCuvJbewobCM2hlNrpl86fT3XX3aPKL9eUrbNMIKBeT58Lk7EZF
mq3kg4UDTmSbU6t6mGtYnscKAjPZX9Yyk3Wn37A0EpLNkbvdLtSWqn/IgKciLZRTEONSLJ/NkX/l
nCnp4gJ/c+FrHj0ThshnR0esRwSLlrjeb+2vDD+QdfF4Ce72i+Jb2lxZN1nPs3bjBPpYU7N8tz1T
JCXjyyZjbdPhnWzhTzM9ZlmGAXyd6lY3WRc5pNEiwrTDd4j/gh3Nd0DqAHwl3BP8QenLg6z/FOzS
R/WGu4L1kPJmN4raDMytwS9ioeUrKH7GhznEF8GbWYEURXvbnmq6DcPY+dIWcg03PImeWsAgufNB
thMA327jk294x9uoPj2sM0F+sjM0c7DxpFflccD7Wu2Gf9ksfdNEtUeWUdJHReksY4VauFKzorDu
mweNfnq6ATLnfqEtP3fIw9QNVY5aVYRtdqR48eZxG+xGO7NnECKPYq4iPgXWwdUNM643p7KKfHH3
7a8X/PikbVzmLNxin02tA8k6kY7BaRMJNP8VaF/L7QSZXhGpHmJIozbbjkPtQi17AXqWkC9+oEkp
nB8y6UyCLGTnkqspeWPPAUXJYEHliDFgSvaVTHAU6cJW1o2zuCto59NyZVUaS72P7tkdkJe3vqfE
RpOAovP3un57LJbUwAHIXoJTba3akVUMJHMuzOWVDVx+vIDpUHxpZENIdxkj8KyoT6w0NIw5wuFj
XfbYz1PASUCj0fX39c8arjtCReTgBQrm4be1oRq7aoRzPF1d/uyboMRb+1M++NVDEsvOCboikMOZ
EfOGZV92mfK3BCCWG6HnMvmygETqVOTnFabz0kyzp7XXYpXR4JuBkQPiwbOHX2fDlD0JPH7OSVTV
n5VY16Qyf/cC/kPXXgY21eMe6Vdl+Ag1v7fY/0Nu3/I84CJs9MPtipdFqpwM4MhUg8k9b/z2CWx8
oJkwQxs5qee5+r2bYMpiTiSXjz+klAMP9CUUGk6Pdd/v8mJxtSvznxe/oZ+Jy0Y1Tx4V2MCc/Stv
p9gmM4TzSz/r9xC+peCzGP2LfVGUgAK/MJHeJUyH9IZpm6h0KmO14yyC3B4gbcdDDFrhlSG/oK/j
WjM9KYT+QqhZ7jRoOaw7QrTIg5E9XK1dtSTGTlnquPPWEoxaK/S/M9PbkI9USg2S9EGXS1Zrgbgo
3wkEmElemQojPZhcpRIalnl+NOwTkB3euhpOhS4wo1HS/GzFQsewstMHM6Kw58e5t4z6eZN6gqHn
CWeo9TgyzhSun4rW3PN8o2oeNik2Gb25WO0FuCgZGhMICkYXWMCTMUCdGE+j1fut20eXTPG7vzLq
ZBKkX2lzUHbX75lxxSaqrpU2etyu4ZIqPRHMd0TCg9elFIFDjtHE7b6w5bYtyr4NG9YEOpNbneQ2
p3OFWDsug+bSMs/hmjk1xDT+CTknnCyEC1cvkTIKuKlr5Fq4prZFCHdtxGPL7iwL5YawIsxyXmKJ
0thwnQrvN8M157z0x/2kdmXGX/0puXsT8YvCQAnJGwLvy7xIFf5mFionO6uZc9sYJbD6vAea50IU
9k+CvcEwe1C6oVjCS+rGp4AJM5XL+SYfUBcc2fNQsZq4gAT6K0w7OZCtodJOChgiIXBRZd2vhb7i
H7y5VWbv93VtCTx5HLnySfCkDwdO87jNogRrDf5eDr6B5FmHt9S4+YFoqMWIclwNSwB5QZ8SETMC
XHEWozIitYSiHfCEY9a99/c9Uz0pBoRqz4rrAWWM5mwlom/LMp+putDSSfCxfgKGtkdRldNlo+T9
IQu8zm+ae7/R8DNqGriS/zZQzv8pLVEhk8Fmg1zs0v05f0kUJaKjDbWBCbwpxEVYVeWj7//QzruY
r3L6r/zogoewmqSoUbNFqIlexpPaBXHJvps/TthwmYcVgsp/8cayLTGingZWGezAn73Aj7GufPBY
zXReSwxdyvL07VwjZLYBbxYLbt5LdkaixeuH1KOrivVLKK+EnyLX9p9MRG+3k1Hyme+BfObnGefH
q/OlZrgQxvjBNG3gtfT/5TB8DTBXRguPCbsy29IjwIntT5OdyoGz2AdSX4mNxU3k62tNwzRQ7+F1
M100BFrpxJpY246MfRh2jTBxFZpxo/1+PgDBwEy6BgXm8aORYSzcYuq2Fy2f/L3TLBlgrGYAKUpV
NJehCxegIb3myM3/T7lqrTlmIUwFyf5RLdkiYpoYiD6m02cg3Gt9PSC/fTuJV0LDdhdERzvDkPP1
8sVQwNSnoYDJAV9mT3r8EzgtWgIJe6Re3Yak9Pk0Mwhbn8Fn2sts8bJQiptKntVeismjm+ry3HIe
1JFkVdU9FieWUPxZl8zd6K+FfkExgQkB/OnhNLbYjYHPEcBt93Fdos2tug99UhTMHIHijrm8J4H1
xCL5nA475KSSXqPtx08VQMMCGx0c8RU64AUxVHFVFhhH3swOnWb0NOwyY4dbC2D+7IgqVzeb51VG
0oJEJVHbMpwMAYmcdl5shGlzcdity3g8YKoCG/OpC9Bixhu3ROl4Xwww//rvcuov3UHNLR6gcPPn
AoZ5bGVwDtWRHXBmS8nXafmnIn8AVTbT70XF86BA0sk31b+BQAU7CrcEi6nEHnFtC/x8jR1V4qW4
1irBdCX+7Jr7R2Xu2oP3u5YZi+nY42+iSKbjRi0qaaH7+sm+HswJxyC/OlKNrpBWXRYlouTbwHAV
wgpzdLjthOXYYItIcw8vcKfCbJH8QQJQc/QpcyH0IZjIowDqQty3aN6Q4RzdPvBgkgTHk5hwCHvd
JkkyDUaDBe7NJwJjHpOhRT+IU7iRFfmCniKY2YIiSayihv74fsrCXUABD8ZKBpK/SfHiGMMGi4Yd
+ZgvNVVgbQ+sIGD5okbag/GVi2QnDE81W3aTsm08Ykrpx6v4mGDmMY6Qj9pGW6kdlUMl8dzgLtmc
Nd/aXTHw8ChryHKej8lnkoNeGNUYc/leqLsZhmkIUkiw0nRU7D1a0XPPiraUUvYCf+qIMueN0/DP
KFNNUlyT2P6baufDqWrQVE3O9hU6SBAnFAZAzanhZ6xzNJgtOJZZU6aT5UAMnGdslmxOgp3N+KX/
PFwDPTh41DjsS2+nmPPDc/4BgzUEVENkuI4bo+ym3chRFy+qjm09I5T2WVuK3zWhGjjUx9h9nia6
zzRIgCbf/JR3PXJoMZ2i8UNM0LUBkEdN2oPLG6/juiHyY91GW+uvhI3AYHJD0qO2hSs9qzzuuoCg
qDVSuge/fZUdUe0pkn8GLaygYC/pIo6JcjmkfXgCCMB2Ji+4kApPO8Rg9foV+JA7Q19FepHF/w/r
YPe728a51lUeGLEgID0N3P8Fv9lHNyWgXTfcVvrLXm95UE9ux5m1Zlt7xRwdQRV7yyixs5R4Inz3
cOUFMM5pawSt/m17tHIG99J38lOu0ha7+0Ea1uRvIxWmYOVyQCeBOkEvcT0MfdERPklZ0bMXFx+I
4EMbbEsRiOjGbm6CYGOTNiitWXpFwTRzRhqHp294WR5sf3ILaembgEisua/hgEQhZKrF5IRD0JER
GNC9pS8Nt8X2JEFrHIgmRsVCC8r9MXN0/72qipy0F48nZOtImvx1Y2wxrDFBNuXBkGOrkzWOlBlx
uLXrapdWVi3y/DggCdCu0cBWLnP0/hOlgUdQkv1F86rshx+iflCeS3UCSNwTn8+tPAiakIgtaoeP
5P+7RTwbmaB8cDENeohQiATjOJu6GNLbnhHC1183cRLy+rUqFyba6D2ElkTLQImmG6YzIZdM8jhC
eevAHAzQRN4KwOMt530vUfTzk2uxuKyVVIQi71vKJE8GwOv9Srze7/F09OvyPvpehj5JpAAyr0eR
iGc5xBB4grGmQ+yFG6kD2u+T+JE2YcevNU0xxM9Tm1YbrjqGRIriiXpayE7+YfWZdco3ajyIkMjD
S3cgJGPwaVOjhkEZAYkiGKg6z7ovdKih6oID8PNDZO/cVNqTKez6GyP+mxXN2NeKUn3wcXSa8c7m
JIovQ5O01+eqAR1A3V65gsRBIHP66YyxeO3lzPXU6dYI7sCHKpsUAeOdgqnbWp3YDXiPDulW/Xkl
rAYI3SvmSWDgLm6K3EeAnOIuNm2TgGCvdUQilb1wFTuotzy681jQxrzzwSHRshW3BRTxz3DypMCU
hb0Rvm0ybUtV1AOyftSIEXBx5w1eZtPB/GxUj6jZrGC0zARtxV4um2gPK/zPQ/cDIMkqiyxJZMSS
rAsHtmE+mguFeVXdJ2/zjiL6Ixn6L5nNOALSex/iBSSuuk8k/TnLXMbLavC6ty1bJhWzZQDMhPdu
HX9N1fzKTsY+VMoe2i4HybXt9wYdwBIa3LVsOBgVQfjIUgxFjsF+yEG0Ru/qKwaIC/IopkF+NF4V
Jy24BlA+24ZmKVRN0b47ExByKCCBHIY5r5YL3qfutfMTHIKATrjXLHKOvp8Oz2hInBffh1pdMvOD
BrbAlGzfrTUITOHulc76IV7I0Y7Y8q1qqycj6c0pJpgZCqX3V1/KSIXffT8tatRWdH4f41PepWja
5d2WmMUJpgrE8TtUQQ2pfS30BWLAYpugW0EpuFE7sUgc/sTl9lgC6KpETczGKCdL72C9l28Zd0yz
m6MLJ66UZ8XTutOJIsY1iQGZh+sh7XyehlJpxydrFgn8uE8CFYep/Ihy6DV8omaQITqm40PHVQLd
/zstAiqBo2yQ94KxjZFaI+rG/oA+okYHpKxxnxDgW/Tp4g3FUlJAw1vhyB6svAbN9eE1A9dMz347
ahjHmk3VTaPGhltaMLDMvDOLDbSSGXgK18Ru47IPyLQg3ltyLM5Dm0hbiuVdQQzqPBlyNk6TUnzv
V6c0rGmc8QG9BomV6u9qThWrG83Czru5+PZbL0Z7bvVUWb7n+UXfhEXHIEygKYQZUNpR+2d7jFtO
ZPDAp6bbrWY7WwaAmyJYdC+eCwVxmP1eGDjYLntxo6zg8IjZ93iNGNkpgTG3axqPzBXMcEjEc0wC
aQKKDAIgzqnlL5Y/cHxbV4xqlIopZ12DKcqYxUtpCa0PglugfkBlS+ACJ9x6Rdwwk7arfqry6n1D
TLBDgE6kbYBFCCvzv/kHw1RAIUEdB+k6ga3U8YmWm7i/U0oNE1kjZBZOvbPJvxXFQRRJvFvWprzy
NbErv4DZiMqwgDJ1emAgFkuIM8U6o+WSDwMLEqMuQzchk+g2COPlqcdVbu4RYZRy0iK9KEc/aiRm
up9BHUeveWqe7Mj+vuN8JzTzqGhqKd0pVraYOvf6oMtmOGwj3BrKnXIDe5sbeZnPeotjHuMX8Obe
mJG5dUtnXgdUoauwIewqkZshfUYvhxWUIOvP+BcajIrNcwRJ9BPUFO6YWMKTY6EuviQ59lIyBUgk
3LOSRxWLBJ12Re76dSoZxH714Q6kU3JX6pIfgAdIjhtSN4h26ABOa1MmfI9+9s0444WWPyscSZtx
CnFkCbgklO7ssR8S6Ekeas2BH5sxEIYLejjtmDFgLamAv39/UXIzqmqKTFnQCa6CNQ2Q/VeHw1v4
drWpOEAJKiXCZeAGOBLGSvR3v+hx+dr1UD754TP09IQtgsKjcPQTgkjCMl42gVRnmSfYD8VGdjkz
5ZeUc3l6Y8eS0uw2bX9B1vw3zQI+HNvleDyzXT9wW49q5IZl7hJFIkiLmw9bUP5F3LnNlYNmkbPe
rgLaVWJeWZ7/33W9MQmh/KNnNVexFaHbgk+aikbmWU4TC64I0m0Dl3R8ti814aTHqePcrdiaTgTo
FCxM3cMquxc3rHBsgttIK2hXj8kBD+F/9bhoJDgGrtAD8rbYe9T95A+cgTi0cqE01VRd6nvDULCt
cJCSW2navQ0JUbdT0gFsrBckhuqOt2XgGARuF1QVfr7m5Yd/tGrWPfXxmmIwHhDnGv4rXgsdBv0a
yjAzxoWDSCyCMs8RhGHbdH6my7n4OI9869UiMLoTzmBMixDFN05r9fwahqwMNqynn99Do6DL6uBW
0FZrmiS3Mqg3zimWTl5+7cZloDCxr6VhZ9qjLwELgPrmDkJ4MITSqoBEAg6nWerCIR1SDOgRrIXC
10k/UoPSvrGQZxwUjUTFIe0TzqHVOxmw7U2SppLQBIBXTLnRksmXjxsVhZOfoj7HL2uo4ZT2BvmE
kaXwbOaZo3ZjGeumrVImL/nXlSoiAuTQZNzBbPWJ9wYOVxywYhDB7xIVGhnqmmqc1JOQ4/c2Loq+
I9fImnN9kuBxvWuxeF4FIvKJ63Oos42zfCVo5fRcGCTfyGo5mAOIfRKUL6KeypnBTQD5Vm0nIdG1
lg333rjXeCKZ2Tbp851xupS6TfF+d2bhh1ergkiGfTObDtssorRza3uM5cZlFbjOMTZv+5jygZ2j
/BzAPEAnzUGDbj8K7ADbZ/mOzj1uZ8QhTgaw65n9K2UDGX0ProJ0TgW5nlkPq6J167OUOflNMp8c
qiyqMGZhfC/92oJ1X1zrRF/ZB94A/Oh4yxguAzOgQIFBUym7DSDNJhb3O/76Qz4HiyVUYAxBcFaW
eu1CTCw0o/3aAXuK+a5XMzv4F4WiFkjdqZfL+RQzatz+cb7Cd8BhImLp6n3oSAwRvQj/6grlLlbc
N7eM+RIaLJKSdKaQPK7pF9vI+7wrOfA1aPFg8PTDU+gW8BK334vHzloz8GjOZZjD32np+551XBoy
OMVMYA5kVSuPfDXXulTfg3P9Y8KPwTsICDScFaYBxaXeNS1Xi8cMwuDy76fFXXD32n7u3ST3oev3
Ggp/sBSdIftLb4f8ncKY+MU8T25v63jdTaVRapwM84CFHy5a/i2yv3VzyRU4WUB6GHqG6KRWBoE1
RdlLhkI+saX2eoRSLMZkzVa6DlWlaxsPL1/79ERq69vitr6qOdvs+dw2c96XZ/5SFZIdjpf4y6J9
0Sh+Gi9iaO6LfPeB+iOdZgTxJSww1BxbpUM7vcX6rL/UI2b3j1zHj7uc57idsSzTYY7Yu1gHm3Mt
eKzyKl+JFrtqOHWR8EPCVGn/pRVawABxlGV/aEkNqKrSwDXaVP0KQVEBxTBmWvgzh+0ObMpWwl0G
/PysP0WAvFdk9iGsCQDZBdG+wE7VhUJgSeJbbdHtwz6Lv+us2bVP93n9nVGGIl8BepV73Xx8zNk7
t2SuPRx28Kaf9+UnwVWc4RcUoM3B1w0bUs/SI6z5Dyr23W4pIYlqE9StNpkJyqckypMijMoZqm81
woLpSFmIb8bvcqN4HJx/habBaGkA1okJt2+rZ4s15zt8xRVnvP3Xt2Y7TIzTN9VLEKUqC/WI6mE9
kN9WQ3VbGlHeWWh9XEDkeXHD4/uLmKfmNMR2N8sFw81L4DArVInTaqUxHCjir9FameOlhKT0MnAo
FK6oiQHNKs/DlYxvqFTvjWp5lYO0zqvoPGJYfaNkxD/rfZ8g1mSJVo4fyxDIDxs741uCWL66Yuyi
X0vu+o+78g/5/2Mg6nEZnozJkW87vIOJncXn2z6Lby4pY0g0GHHpPZkyROyP1J+8hjIGuA2iTeoW
0Q1KNwLuAuwvpAOtncjia4twQL47Hy7wauJ3t+PJFazAwkPg0tRQik8fT9WuqNWT8WUxy4qxcj90
sKbOCkySZwoyzXOTEwOTCR6eWfRYqMqeNGsBI9AccuwXIWPALYWKnK9BV3nfPAvAP6DBXWoGp80g
0bk5u2q72xd01Tciif7lp42a1XffdBo1Ug1Ku6fukTF0c/7mGulnaDhezNknR7gVujShPWZ86YG4
v5okj4EaegQ31rXTKC24BlQEgF/EtvR2zisSHW8j49eJMGQyz0AmbFDTibW8zGBQ/qC3DLQj0Sgo
yO7STrt/7ogJSivwhxcx5YKxvS4drrCJf+TBZJXCQYVGqnkLP1oFBcqrphoKxtiPT1+wYFdo4DdM
xUmMMm+2J5MExw/RU3iF8WBGIAbbGhBiFo1CZ3kCrZpeApNkVMxIpJE6SnnIHh/6v0w3HQ60eQBo
XyuL+jmIygdOnmw0wYe9tt6f/moo2XS79Qtc1hCSCCGU3T0sRdCulHytvKCOzDK1EFMgkTU2+p6C
BQH35BVhVFPi0VCyfSvaj8dEoWLQwRZJldB1+NVuQ5ashCxIETEfjejnlfpIYDmOETsrAYzb8GLi
b5tuC6K9yRkcZiMSDDGlOI26iYpl77CPssTZfvTZtaY7OfU/9DvUfK4HTbegIhenhJ7u2/9IUwpW
ZBr4m2LJdDnMtoQy+xP08Qt/cwSwEZqez9Cfm+t7td+hhI9Dgadmp1P9FANl8NurMvc46tSF9ugz
zBAeX1co5I9jOGUKyQDQX+Xltqwwy3aSstdqEONaZhhdMFQlG3TT2aslhGP7IgeNYO1DDN7B942a
IFhsutnsUFnJpLSnkatP+8WJ3DeP1EdSLc835gUAhJARMYV4F8ib73w6BFecOTChR6kPmf6opKn3
rL6Ez/iGyeHW6cKcnlNk05EK2Jmd1DCQ83Nu4VRkVJm1dDrlyG+hwYFDlsK20+FweJ6joDYFV0gW
hhz9tVI9kx3k1e/f5pu+DjWjwIyUTN+ZdCZW64vkGaaYce8qkFnUMToYz0/yWDbAiNDK4fRvyTE8
Fi7AZTe62ApOKHgNMuHRxV0WAtiiq2afBTUllLcgp6cfwumOCVWc5gFIod67ZR737q8fqcOS1bH+
UCA+E66JI8KoE1LZPSMuASRQu9Tf1SDe0wmtnjdz2RKvNUIwUuNGmtzm4zWtqOWy1FWA7HvbSdXA
6EIOJqL9PiRgkv13Bbr0v5SSHDMaRgwOc98RN7DY0wTHY/p4hpAyXCH09HZcwhiHD4BSQQJiHpZl
GmknOSIEFC8803uyfirefsBID8ZAnxYGnuDvZZm3QzQoSNtE2bszvrd/izpm4ZP+giIOy8n3cdCa
yhykZ/MNv8VUICPPKvDIkGArTmGIuOl8TAw35MOZYlPwOlZ2w+8Rb1vqhIeuwMr/NV34KMKdRfvR
B3kt6lCGq8LGHpRrM+HOhp3WLpm5rr03D8ruV97fghgkLiL4GpRvQ9DGHMrTzMR9JUyIXXkfDPGi
KC1xiT4BzOe+JX6c4R+wQzk6F8kXQmgJkmlYv/EuzYKKtdetXR75++T4FkI0LT6lM4LzzsWcKbUz
3Xss+dKrrWWFBy138MiR2RIc8goMvAX1LoY61xm+GaN2/87Y1n+YQ5mlftuy/3kYfVsJd5SAkqQt
okj2rlJ91yAVcd/rCpP6ObwWBM1T3kiahd1OIWDCNe3iZi9HCKqJf4jRG3E1yP7bUuaFolL+YLV3
WOkDvnjfcRXUqc/ZbpQ8uP2MbwE63X2vWw1CDbsBMWvdB6HyylznHtjHhA3cOXElA2bEXb2v+ePg
ghe50nehQW5VAzVsrIsPRgsGYZdZ22spyYFuuaU/L9Bw7ZGhjaacbLFwWlHb0OI6n0tjj2DGLUIU
0ebu2Redy2cjdTnoHxLqhRrsAeMw+JQhvwFJh/89N7NiRdQnK2R7bhQsrP+DXf0MHIOWOVc8cJ8b
tywiNGMvbMPxAGQxtYh84FZnkRTkDhmpR9Zr5opOofi9g3G4AB+6sdYOU7llo3Jadf0QvtmdogUK
J0o8dd5bBNNy/+tTUQ860r9aj36cIG7ueuwKkmGiNTWtFypY9m2dDwCfVqCoJrR2onj6gV4Yvl/B
GDTjXmL9d8m/gTTB4WJNVkA44VIqOfM10/vWXxOdo60BQaxFTabrvglnWHY8bICz65bEx0uPzvPd
BCk4KoAApvuNKU12BVq+q/P7/cjgT5cLrrAKA6bEFxa0oG70sOsUtBPMWnVrwao6h9HJUJX0MOps
plPASMSBOzswpPK6He5PSMhw7tkCJV66zUwpeWVunGH22xqXkwFYaHIkMn1Wg++pw5SGxlB0nuil
GHWTTjg4BrzOHG4YjVPApuOJxIb0ppx2Rc7CUOieolxxmt2JE6fX43NnFzKYyKr/1RhfJDifxqCI
WfoAgTI2Uorl6QbwBr/cdrKKkwYjVF6WuhQyrND8u2ecBioKe6qvrYIXYQXEVD/e8Ob9WT+/PPlM
Nx/+FabzrZir+OzVOM96jFDNSIyIw3doJE6c7cjo68tjUgJ4OfscrrFxpccbHUaGvQZCg8m/Ib5q
3W5LiLEsxKYp8SKqRzXwxx0KSyCEXhFWuPZiT2yOVjH4kOW7OSV8poFlUks3L51BSbdY8NxTRuiZ
BkfRQonZRhZJlqnLdbTuBV+PjPh9pRGQZMsyUVLrxDX+ueSzlKWCeKX+VIOY/sXZv6PanGY3NpuE
W6FYAQM6SL3vT/bcGSy8kBUwkX5U/lZneSN/QUsA/QtD6eB07jJ1OKzNyYaoMUHfn68MYqa9DbVi
x/OyXat0DB+0YL/5pZjrvOhfxM8NfJCtPtM6rPkdHa5u/i8EYGMh1Xa5i3IyP96dApj42JocITVx
N+z/6/bslv/Zz9GCeQORAKOz3XyZqsTS0aXJxaVcmmN16yUEube/9+ZOBVaGKGRiZE5TCbzc6xHH
EkO1Q8zUFyJS5UpAgnUZxq7RZRc80Bkz+/c1QB4Ir7CkjIVejL+8PA19tYrgW3dC23RKKXUjCw+g
w19aUkBG0usCU8nALkpa3nZ7jwG7yYbZ+zJJ9sRgj6J3bBoQCXiq8zWsuBDRMgpgFg4Xw+tKBrPY
5m1dR3DB4YjwIFGhUJkBVsbAm/UQnmaHuDoaeMeOe8uh1cGKyJirzddXcVlxGdkensH0F/7PoxSw
JwaxRbSPr7NrnNN/Ohhd8HclhIseuAmtcCN3ylN4+rpXk8TDpWHNx4qCIL4wxizqku4l4/P91BT0
fxUBgPvGUPSFe2worBdK0dVGpJjvzTukyt0bX84K8/2zxigxjDTif5aykOxcQCRsn1BOmkhPn9pX
bsJgnZJ3CTwM1vQ9OfExnmrqGvOGFOGw1RIkYrEd9WhggQ2jD4tX+NzrBIVRHVENxyLokPS1jmME
mHfQSm2r1NZCd6G6KHljLKYOUMeKKDhV45mlTWP8ZJw4jRvOVU3XwcsdM0mm4v71phc7F9rTKYHI
KD//tvHDKdqPuqwUoXE56OclsQOGfx+PtzfztvNcElsy48lJI0INU5ps71fZ+tK09G3mswTVXMoK
BovgpnRphj3UmyaVyZvR3nCZLFhbwqMFKwWypa8zGth1d0Is4CBj5k+NezwIthpLzMP29MyjuEcs
FnTICnL1T108FAcv+6K6YT4yv3BloMqyX6ZyonGp6dKRuAm5Bu7U95l/4SQN0hobvNn0vu4WIujW
QCVYnxngXcnqeh2nscXqGy+3yd44P1W3VnFDGX5WQCYxessypVpQsW8RbAlv3eGJP8taDpApc0hz
pGsdzxeIK2hTb3ZqExI0l3jSBFeCpk4b9hE8eWh1QnOiBNg0gSMnrwBLUYKn2b4P2WzKMDHIWjtR
5KrVcbC0Nc96J1/jxu8lBqIezkyzvagZ0ouyGWfsbeR6OFwyS4lqoH1s3CcfYRcnm1EQ0tSZtXE7
cy3bAiCP4YreeWu9H/MOscamnFe9mAt7Pdl4pVFoIPljalbW/28IPSjXswvKDnyQ8j/wFVmG6Iua
jmGO/dld+NTvG/37OON21FwjyOU/IbEduRWdvvPw+MPYJjlU0F/ZDdSLXWdaFXVMfPlDyg4WOqU1
TS1fhxtRWdNkfUBEa6rDo/27zUxECfGUiqwcl+oh1fzjBvXl0fc9b4OYLi8icwzNSPMjIc35Hdab
Hn5L62d6ydThJ3T8GtZdNEGPgAc8GLk6/Z7jrZJqB1P752/p+Ko/sMDVZlmW1MXGgXEQ2rDrk3H0
eHau8vAvt8bYOQrkiOCYvjR75EyMX2KGF1OQFyL1hyTFaoZdV4xYtResTA9SxGF8Gf5QalAjmAao
qcgDn0uomHfBsKVsxMLXqV9BjmleK5MCKhi5ewZVAtc2b65OjZBKXrKbBlO7NZwHySxf8DLARgF6
PlO41xOKiQCtE43ubEFely48GU/0X/zJNsjnl15ePLgUngvkYmXle9WTh/5gEWG0lE/e2Df/Nm7s
PK3cLDsLRgMTRwa6IinVNWBM2RUeDDiNgon+NbSxsHFNiIrvAryrIpwwbKXhwDDHapf5oJbJ63KC
7JN+bvvpvrUSNaYA/L14EOND1m1HUWKE+M7Ez+toaOpCDwS4H+5eAIRVnfErx+1sV3b/MJPBP8tE
CDpuEWO5Mt4JHKn9Sc8mzOeu6hx1xJF/474tUBMhUzdeC2sLPl1CDbQU7gCTMxPghCj2Ry69a7we
7OHnx26crkmAGiGidqdIZAB57bNDh7RhydF/j2Ne0e9jXKPu4xvJ0w00MjdJ2LkXnhRx+XRT4h8s
44eldVABi+Oxw0n5JQGtybPlsN7zJlfWwdEo+q/npmRdEtsmPBhdcKXc4TG4QV/ECMzDLtC5ftCH
kltvGgvU9FF4nllPXKmxF00Ega5lXDTbg19qqdYf5sJ4Q1gmYqOZroa82TJ03qr/gPmuFiQhSvFH
bxOqcb/LHr1PjtA/GvVH4SRPzHGqb1lOJtr5EliY1L/pha9z5HoymvljWjqu8O2YULLS2wor+kgy
XnJ/5A3dmfldkteGmOQhmnSdnRzubwAHgUTCzWrpIh14qHsyrwfV1bf6oOXjTomPpWpgoPqM8sp3
VbvPrqygG1YPdmlVNiwDXCcDWwDzp5uiWl7G6/YWy5R/Tk4rYC0MUevlTsy4GFB+U8aHc7DUgIKH
H2W5DgoefHiLK/5VxPvXLGXRNFPYt888RSuTiNLktqoFa9rccCZ4R04AIQPEHPViIjyySqEnlmST
KSgBzmZ5O3fF/J6LprbeBL2piK0AIBC0zkEqyam6fCCgAQ/gpFn80liph0D+0WmYQSGg97DCwWdx
86a4WM+rh6LUm3nc+fFPzmk2NuH8t4yZ4VDxrjr4VxuFXtyjxvgKrfyExaRhZGVb+OoQZC5OCrj4
CmIrgxKzHnsk0HHOAloffpJWJ1ygdsyM5iBSAJim3cM01y8ZQKXFpXEP91oLpYgUvymH++LFC+s6
K3hHi07Cr0A5qPqCdXmkAPWEUsZk+z8U9SZgRWTj9hIFHtodsxKNKoP6g/Glke5OlfhoQe4xgCQq
V1flVUbWkrDaGd6QYGc5qG6ABPMLGNEDAVaEGdCJzMnBQUpT3c4zFsyUY2Ba5/C/TEleL3kf89vA
7QHGsribFuOfcmz9manQEFKkFtuK2lzZDn6HTODi9bUKozs2LhgotLiE1pB+6sKY+Rz1chd8o8du
C4L6Y3a69JvEXAdZNypErm9KIMm8orO3O3YT6KM0dqF/Cw+A7jPNH3WjyIAwxXlnKh8AQQUHvE+l
a119QtDpfERzKNtOZ/zff93UP45rYTU1NF/abYyuRr5HfWe4I1rYea9Ty2WLMVRDHkoIgWXMpi+4
ppjNmFRscyKpHST3EA3My+ZjzAbH+1+k4AxNp/YTBicPMukDVXPhoVpQFpIsWXi0AczQguRy0Xvm
X2B3XmZlWKD7ULZQhcWMNGAl4YNWQWY6wPAFMESjZDrRTug8YFuWuiptakyAB548/eCAWAVv0F+v
VL78l9Vyzk9YBZi46HdA54bkH8RyZLfZieuBGDUormQoFcB8r+d+E05SqsbBOGsIAU6L/ieiykcE
3G3DLU7dZ7Rk4dib5TwikU5rA1LZjNelo0OpAZr2sl9811EIK50Zwy3ex4jarCEihOZJGRHOvj/E
gwaXnHsJ7SMmCr+zh2dZWcum5jt5PulCHyxVQeMerMemFM7rMq0E399eapQt2n+36qpzhjmy1rhV
7QHonKhNH8zsAoFpfCV1yY3kiUHK9WQqqsIvzC4Igp76POk6uVOtTY3q0ylbt+V/xg6OwebdqgOG
uszh1q+1B1UpYx8ZzeOTDPjM/fdTq8GFBNY6X5sCsGyWcNpN8rc+EdjkjCTXrQ2KxplZJ1DITepg
T7QFEu0SkrUdTT3MHX8Y8dPFucOSKy2bFCOjJKK5kPTkUoDXzyXqD/jdQAlAGPr5SioNl0OECBXe
A3G9lGbvRNtjilIzNzZgQpQ/AaBaZFEZApqeMAPnOIywtP/lphUAtgn3gs7e3kRi8wARZnhOLj56
Q6iM53lCgG+mX5FzijxIIlt0oj9CqRXxBvZFdUlt2j2ffpUM0T3In6Ar5s9hanDoyJUD4nBBOlR2
I+M2GwHEA58ULc7OF5g4XxXDiF5cg+yw06bGnmpSaHFQdwlb+1rTZu4X5zWWj4s5mOIxtW4PFMkX
8fhAX1J/JXp0fSm7aPNfTjRhmL9/BLDZ0V01k+19RB8KP+LTgT9DwaB0E6v/J3zOf/VbjoNWC2B6
6ooFz6cGY+Og5jH5TMY6xkbD4jqaLX2ro/tUHkIjR4ygSiRPQmobq6Ai6cARMFlsiv+qYNUMc/2M
oqwVUq3UsuT0e/GOUiuf4aBCOdQ9Guao7RkLgsZGSboWDZ7OyFKccsI3g4s1Lc+BF/gdQeJKJsUH
sYpmuF7ifPD8XueT8quz2XpaE/thV0u+GAgaECZqlo8Z7+L3Z/LlcJTNfwQ/oAbyaXM1comFBRqv
iTOQPnN5x23u4Txak7tsV/zG29bvhR4huZxO4pZVVW8JexDHqU2CWtYs1P6AcgGh5pveqmrtnJCW
T0EqQ8B7K9/1xDYHDnXkAYbo+nKq9VhGVPU8VT427jZ48grvgqoC5PdtWAyyelyJagV9Jthqu6jr
rQX2tk9k0q8Chvc3ISp+QL32Ldfq4B5OHiNuRaOlXPCDDBWrV/QNAPqjoszHPAvqlLyW2QH00aFW
yshim9TXY/Ei1DFHTMrew132ORHBpCqT6JordGhgSw3KEw944h/x0ZhRsq5JgtLiaiVVE+TqZoAC
nvXy33CiqIbOvLQvANLiqf2Spv08TpNxkEi9XjQbtMklWZjpYy/xjcesnvPol3C8Qp1qoGTSg7gS
AtUE98P+IeHTpa+ufsQVrTHpuy1qSkf0LZWnahYTDpE7Q91CoOzTTq+6NlzyahN5vkl4zQ4SEx7s
cJQQeeN4R4zUaez4KuJ1LYHTKOoalZR9teL+3I9nDkeMV567oRU+/w53UivkQSykHmQGKpoRUjy/
ZeHXwLIR+G6IYL0qSP9J1cT44pJQbmZzYiTqyospUFukJ2u4uPov9tIjhw0Q/ve+eyndznOEXO0I
JTMhlmdD4DG1F7snMhEJCxrvIrRhUnm5dq7cO76UGOjmf51HJ83e1Ge0cbjsPwzFEQrvY0eilsHp
IZvnnJc9lJQquCjukjc+weiTUGq/wKDS4JyHztRwCZDS4P/uC+hbSloi/6Z0kz6XFBf/4aSRjkEU
a2fnliaSDPrqAVZnjJsls3t6cY81x05ho9WNGpyGify8KajLleTQtl93kplZfEBCex7e4Vgk+MtT
bI1YXNwTFg5V/ZPQkUdH0I9BQoZovJETS3MKyGc8abz1l3J1IKyjpKl/Go/pp+L70OYHql/yts2o
LZjuqlDF/FSJ5iJHiZ6EkGBKi7PTWA7yyjY+SUso7wLPToZmJ2fPyZk+T5sDKfyc0y3Mahf6IwpC
wKdD67ApawbxzRo0uKQxH8LKEcpbdPUdJ/yvMTyqSe0bVSB55aCJEyDpJNrfgSgqiz4OuCe8sV3g
J3nboTrOU+9p6e6EwRWfiVbU2vd/Kd/O3pjFiClgO7sVWAKL8RXKGpht8ljHBb4Tmat8NYTyMT5Q
l/mBBbRTrqVdiVQ3Edm5B/v7VbmozSE5K9TAYSBXnKn6pAGKArsPtgqvcX/2EIoLAREziLiZmyPC
Nt0V8stlHQeAPSfO5KL7867zI07wLDLutz1xwWeI9PzPavgEmX9MD6h3NccpD5eqFi65PqccCsCx
sj/Ku/VTdPOPyhRP3tK+8DQ6mhEHKk6qtHiajYVLlhIqE6ma3Fj6cmGlObJyTBsovxMVMpB6Rxum
CUD3ae3HO8W/MLfNu4ZY7JdFcLy+raRnNk2QQEFNNDb2FFnpBJkt6dIfdrrGHFtH1Y0iCOP35VsE
JgRwHv89x25cc/6aMPIRs3uU24sbOwE0WR0aL3CNibDoi3bCx76ucWwr2GZJ6uTfJYgAGsbU9Fvi
gYWOsMkkzLtlQb9MDUsInnLzwJSzydY9yhSIn3zzc1PT0rmVNYgZpR7qGgMMkYOC+xTqh25IwusR
NB+TP6UpD450AYAOTV2yUdpGHEp0kaAG9I64bwGPnVVpMb7uK9DPEDiW2YTYgSiPeUYnlr5IuDTF
Q6DevdYPqLbykPFkJvCzkZhYEGPgH7XR2z2NCUgrr9kpEkycT/AbbfXvDPvSo1kN9FER3q7doyUZ
4dmoBEuGHadjXm47x0kPPa0+5ccEyYiUq2SunVLRO7Gu69+5FbuDYsKWuvN5iWHAPYZL4x8P/FLu
na5s7ApFEMmhGFZkmXfeRL6cz1t1oSWwZjmaeZRiVeTEakCalyGwsE3ZYu73ueLbtaCBEVEWMoJ0
na/ABLKW9NKIsB2DTwjEXYpu0aLNp25TAPfSSdxzkCHSG/z59cr6YYOwe76ee2wYWKiIAG3yxeYW
FjGECPoNLKMA3yvm9Xwul6Yx3BfutstGOk1QpX/5ExfQylPjZNAsg35LZG5H/oQo13S4py0Nb0Cl
dRJDp3d3FDKU+9oek+6ADIdA3VuFElE7J9nzh6WiWt7G41wjrlkDCJAN173gb0Zw6l5qGSX/uFOF
U3LDFdyvCwWuUVxpOS3/JhznkBzN/48vkUesKBkZq7QlcD8CTVXZHNv13/yu+iLcHNwmKVnp+uSM
j1myf7UKXl4HlIHJ55dkKIAVNAbHMY7n0bJlz4cktyomY8BREMYd7Q04JykKS8/13Z/8rDBY06PS
eY2Guhu/zQhMjAFhDQ6/DnLlIylLhyx1kdD35eFtnnCsBb1R+SOeXVclHF/boNwyhQzg1waOi9iz
G11xt+7gRA4PSFWLGB6Fs7oYLwG21vmxUgjx+JdY4izOHty0uudfsq6H/PKJcLSVWZPqJMQOmjd0
j9gEEavpd/PAteMORNMxOjsgALfIEN3RTS3aYVOjOpCUoJAbeRZx8MAl3UnsHoHOreoLHFll9myw
ehKA7Dua77kvLtxvEVYGYMyuS7Y5aAKsDKIssJMh+MaQ+Jgv122X4iyUxvhVjQ9MY9SLJ3kgWJ4I
OLBDzjGOoai5821FHEZo+cjHTU1Os+jwQD4ORWdb9Bm/d84iK3r9gyyu5EsHy8e7XJHRt0kA1U4K
wWB6BUZeSepB0SblwkhbRbqblU0aknDCF9ierWr2CdBRtlZS0qnB8X/LXJtZPeH714RvRr2x4bnJ
s3d5ArEmLHUZBIxwppmjg9FhcEEgIA/A6SKpOPlO5SbKn77dQWYuoN9cKOOlXHillwDbzIfQtPy0
KyMzlR0ZrOoOuS+mRRB+NuZLQecr5/HqSn4NRw2WrVogS8ooD4AhM3+kfEGMNlIC0CDzRDIN44lE
1Wfqsm4+LOz/exz1IV/Bg2s2Riz2E/Fc33JGBX4tvJ23r+91vKBA6EYGv1nrklv+Cb/zMRH97orb
DRqw7iWL4C22Lrxbj39IxXnhL34+sNfgGWzLDZaBeGsGIZW20O3B0XJ94qI2SJGfx/5gZN7BL81N
xJj3iTDvvVeKZBvRIxhVV35sBkpACviAs5IwJz8hJusX5svjWLy1O+0VOEn8A0m8DYsMNokdo0OD
IGXyAUBbCJJEJQ6LPgLIqBsTEM2sGrl04Cd+2bCQY+HNhhZYZEJ/jeTFbZaHCIQbq3nzWahgY+ia
0O0P0+wgrynj72qQXRWn4H4g+aSj+uFT4E/FGXTGkOUoP+3FBbemKrENGJHhWDc3RMFVUMp1yf6H
OOlCoyHZtr+xpAaO5gblMMBOgOia8CvGdr/QWKW9v09b6KC8y4GBM9bibd9sdBij9Igs41pgz5iM
jbtE/ko/Ll12yIG+lwabHkKmpF/8xqQXjcNjFvYukU5Ozkr0OfYCyyEbHSQICgAMgobH0xZISJze
ROQW0nIO+sGUtQlV7/5njBkP/rVcWf/vNM6xU5FlbJShyU58RowgMf9gpp+Rz7/Z1W/s4QGIULWf
mwoHktC0bIw5teC4V3oUxlhg55Tka6DQaivxG0cuvPMHSQj0HThNe4jWBrUxNJoSt90UZVTlt4Uh
xy6bbF+PKDt8YK6V+QoPaS4rdPO4Vog6RjLJQlKtmom6O+W17wjXG76oHCiHspeF+ZbnRx0VR2qo
SEHfeSX8wbi8AQCBCTd/RdyqnjFbFQSILncOK1c8ipTIF3AqerPh4K/ypMXPfFz/uSHWgBXX2BvQ
AzMEYX58umpBleSjoqJ/+haI6XzShP05ZhF+Z8VptO3QrqMrJYP713vLBPO8fQP2vVsE4ziYU2DJ
pTU48gV1/hXhNEBpw23C5Yc4ABca9ugvq2yii98C+d09+3RZ5DobFWFRJawWdqP/hRKH9+JkVIYA
XdRyVKHYZ0GuUCfL1DKIn7Oxw1Kov90BKYmAVcRdMNb/pSwZbWy0zRTpjlRNIT5oNC0d/hQqSSC1
GoFSjMTV3hGYMrVbMCyJuuCp3DKDhYo1dzjCho2ZdX6Y6nmRXKy1SFYP2djU1L/RBYw/9pmoPuuw
fI3xGXmVFG5xRCLyFA7Ec9lNjS609W9tAz+YUEitsXBsNsQvSTEpha+SrGkoE+yy0RScj5lNJyWp
zi+9WN5VVkd6hbG/kpF19hJhbumd2aJKSqR5jmMBb/coGq985On0kuet8AKx01V/uNkAujBvD6Dn
zp0lKlfH738XjPdcnpOk/AmxVapr7tvpOyjtBCdkbvyGe2+QlJG3NOov0Bfhzo1Zj9LT488poyNK
fPlHxNr7PgEB15Pad0pmRFwG2+zPjQTFAqy/f6kKmgsj4YJhIB/TwoJhm4ZMT58qpy0TwghSuK/4
inxaQa9uS79cNC6hhZePXKTZCLKarESp0REBixkGty8Zh0l+6OVA9p2bn1qOGohniPNEn+AWsXMj
c94Bl6KxtsI6fhg1MjmvuiL/TJvKWtWRjQsKcASKCjomJNrEoL+0XBCy9GUfvARCTvMOvTVHorhJ
3aMf7Hn5QiWIxroFA3dcfuMgyfEScU/JmSSEydSrKeSn3raLTRcCxyYaeWaMPpa3nnWug2TdxI1m
Aa2XqiOs5D6I+DFd/p3cxADMmW6TL8E73BN/MR2VPbZpWFBNBsHOYORnxg1sCv4GNfkICvZjuabE
AhY9AIjr/Q9Xp55sNOTQbfKFfSNs2+ouwYy/AoJQo85LgVSxWs8tfTKWfAe0iVpW0mgVNJwAMEEd
zeKOzelmR82eeg6zn2lcV8vJHSHhA1NMfu6oMA+DQm4SxFccqivLTedxzFcevH62wSOCp7Xo03SH
g831gcyLaNTNLEdTD4w2dmGi8bif0K+jnn1Jhr1NHluoD92JtoEsegtpNKHVTv3qOjlxPfM/u9LJ
INEdiZsMtZoEqrmR9HzqiHMqc8eA0SExusUnT+rkWLyrMMAgHNWM184MFt1d9YNOQFuSdFmiRgN3
zacN2FG6A3gZ+1XkZ9AP3iHvPeOxVDeQZTvmJaHZ29FzQQMO6CpWrv0Xz6fhcCitk5f//7ISrLlM
flFNoF6U8w+zCZyIURqtUHrUv/vxL/LZ0rKEch43ck2sUa3c1iUmt2wFldMJry3SjbCLfscYHdta
3YhdKY6ON2ykIvymnDw3FCJjJcYFvlbME3+d+5z8eTcGkzldmaskY8HgHowfJTIqEm5728qlNNsl
xpQ4nplr2JlGBEhRYPqK7X+b4cGF66pcudAtwiUBGWjEG5V+XbfhliEWVAq2TZGE5y6x92b4VYC1
QR7/oINWQ1tLFjR0ZKkLl+poGrlUe6OfozqP+EgjrwYvZ53vAKnzYh+e3tBGVZ+W3/RkCHOf1gMt
jRhXaTw6UtKgW9Uf1Wgz8tlEMhrKw7jQSZiIHgb0UQvvCTxsVTkyf99v8aKfPhx9SnQejOCUH2Ih
DurY50jk1PtHCWFQEyLqyTuEyCuFkPS1orYPPbxITU6OjJ0BMCJSUa8k/N+VNffQPM+arqe5dQxE
Sha4ISqkwut4J23ESEpS1Wz6MuBDeBwPqVT2YFPl5U9Ep+dSkv5rEDrj/v9KLbUBTxjdmrbt8BEO
B9BQVdS6bC/eQfTiy8LxHw11f1GtHIQIjOJZhcg4+OJNjnZR1KGbQGx4/HTR5XXlwlaNSrlqekER
qu+51Uyv797DGb8XCHF/2jl6EHCumJ8Qa0YD25M+0hS4Q37d/GbushWMvuWVKI6mlwEXwpGtCupK
t94pFKHRvw2A7rXMbHGZjX/N/lANhioFIxxNFer8lXH1NOzVo2O3NcdEvDY+Bd4nP0N/FSq+DNUP
uizwyjEE8/9HMIX15yOCvR8leE+gANbaTtG9mIfE7SV+cP1nu+Safs+ZBWgkqxVJx298vSfO7IZO
Nn2gvZ4LWC84siSSDoLs/E0xoHKDi15FxzBO2ZyrEZBJ5iFaZlXG6TD+b8J7MEfLryNvOekYYF1f
0EacafusE5I6MHb0XUqzZEUnWTDQATV0jGKnAYTqoBCSN+46TlMyRmmBT04Fjuw2SN5SagLwu9OB
fhJ2trk/kp2r47O+rac34Gp6Q6rQym5AtM0NOUFYDhhXiJPAdA9m4rMT14snHMXWu9eJ3X1DhpfH
0fQUGg2BYaFtSXPNRvNjyRGQ+IQWfin4OCFYB7WFWgTc9Uz6CRldVNkXFHIWjPLqeSSpqSYxIhT8
/cplNtuPgPQdHxqen+gVH576bo7Jz8Emb3b523J7rP1YArrOS4xyNlhzAZjwayW+4e5BvQ52Nxgv
4CmFFVMYO8qSXSjNiQymtXlnrajQhTehvNoG13W0YBODMaEGONanUSsv3gymU9X855Wh+MnVpqJf
IEqVbHmgKnvRe42nAmu0HE4JHqwf0ZHnnG8x2UggxTC6hknxud3B1BTbQIRpBEg0QCQCDYYBLuK9
ozBwv6/1kgdm6tdRwabmt2qXdt1C+unT6Uj0fDAxSlmW+Y7n5VgXn5xkwVUHu02dAKCBYVgwc156
zKAWhjI9k1o2wPxGzxYZbXmJXanJ3Fk1prs30+g29MRzFxVIgnIARbl06BoJs5MSVfk3gaX5o7lv
zd/mP3oy4DBYx10bFDtvpVesUKz517t4rTtjMHbIGaENi/VI7pNFEX/df4WxMLswJ3BS4WW5Xddb
/8v3NxFAqJkalTyvlU2DfVBhQhdrVcCCFwryEjITI1THoA9B62CZEMHX7tAyffywpozO0NwngDXB
yY0Lt+Mb8xFX/rfTBLZVoAUfU83cTKrrF5yDtdeXf5nkw1aZLgeQypDGqEiGWYjsG/qkkU9kP8ZZ
tO7yGfWKROCO4hukfg/wmb2tvkSvvoKcENqXRWL0t8/UyfyaRI6nJNdLPwNe+CNTD0+76NBu2pHG
9mjHDKBab4OsuIEH68x9h1UUXB6RnVwhD8Eut8ggFCdkVnTifteuBXJTdesFSJSL1fajSNH2RBRT
DVZ/ydYyXft/7mzviUBew0erLZJIacfXLhKyfbzJdBIW2/tsRNO45gZl17Bt53JtR4pnMBtNcGRr
RNkDJm2e4Deh+jx4lEyAYHkg6Lf4K8DsmZkOAtjR9OSlmhJzcSpPJvSNBdVHHfs9K1qlhcIxY9PI
JG1KqnItdic186MgPNuYG6E74M8V4fR+9Fx9+PR/0BWHr9ekBF+Bt4m5ljdjXtABVCUlczPVNQUC
4QoKtKGoc8321CoBKO8BR+DGC5Rot6zrf9+X1Ll8ie5SRR8vm5QnPmBsGR5Bsx+mePE3XqleyCp5
YqHhvmYmJmT4axiQ7VIb7PzJidySi0a2SW+IMG/tSZwH0fs7poIyL6R3CJ1tLUZeKtGjWJ8iY3b/
dV1QoUNxDFoo0Q6NSXCG3HrkqXG5exBAVWEjSF2GeDNTG9C+DyNs66/77MxzBmp7tV529uDuReix
4v7xU00IlmK2auJv2cGLZutmCS2EimJikRGm8cWuvw/dM4ZvcWUg2SuUwRZfPRLGmA7M+RT1CHh4
HfsMrMMUZ2CDDlt6KIHCY4KVL8tVdoPOjlZyZb0+QDGNf+oXL4t+cW++5swo8S37HONSqLVF05tp
dJH0GZSMTjF3hWuLs1R1p3DtglOKNwrfjBBGGwjlM/yXrFTdFlP6arYJsXhq1ISvPKKSFFAcD6s8
CpPMf2+Xdj0trWqX2BrXUFfsOeWGx3mWcuUt8yR1kg1tFUUenIgRDD3UFEZiQUhhKp6JOVwbpmFS
9sB191o3WB1i/8StJGci7NEVn5FrcUOidsthy7e/Cg0/iQKjism8p9+lOdcKiqItLvy2mHcSAr0j
ViutmoGSuwfCFf5JgQLiTrRttLx+Nw2ww+y8AeP1Y0fTZtTZa+Py6e9R9gsV6vr/9IclXmF/3Pqk
PrHUr1brfQbiy2vjougYfDtOMqArvieHWGqmvR7y2hqGwe8E3D3wqbTEDl8R/GZ/6XG5k51baQRa
wwO8rnQKJDzO1Lwc4oblzIgALImdYKKrq0ZDJ0W+Lc64rbn0fl4k3u8Q6B06Gzcb82/bImjrCrO0
xBz5RLvU6rikgwkPippoN2gNpGY2VtRWhZlctgbJBBdDlsNQ9+Ki8EyqmQnWKmW14pH/BLdSshOv
Y515Jl8L15y0Vqt2i2PKIAI4Ul0ed1jvpx7g8UIHXH+TBaOXcU2rrwRE2V+bWHGN2JRl1upXxGDa
REqdKsMAHZHr/9PP0k28cIzODOJ1ny6Ajs98eSxIzmP4Q4hyj3rWlACp9qnm9WXey4nDJHNVXbh4
0Rum9mRdbM3HQRM1sc2n8oK4r4oDMVVF1AVWYqVBgmcbjZCv5fmIZdz3Cks7SL+thV9PWZaGikzS
LBltLRvIGO5uHHSRXnw2IiyCTjEy5XNp2fdt0TYirxkV6Xm4vHBIMVlLBfgzz7krZX5xeugHMAaw
UmoyslikLQN23aPuexsQsRUZNUnBYenn28h+sY2wSDcb/EUeUgB97MsLINT7pJ99VFSxO7taALcc
PWV3+57mysmeAAlrFEbBBDwzQY6d/cQLWEYMIxK2gP9H5jqxXcSrzS1J/yBE/IIZa53dD61IbTE9
1bXjWceI+IASeqVjl3/Ycex3yd8PYzJsMGgJW7L/84La/y74sIj+J6BjYU2vqDXzBcInRVlh+UbC
xDurEdinQAOWcJJgx5eE7bSCpIZYCDdLmgK5la/UuTuaYvYZJa4VGSqP3lJQDial5Z/22k7Mm8Bg
EacrCTnnoyau22x+GXgaoLu6njC1S4sS03ZCg2XT+LjZr6nNbStOYMMYdAxsoBTMj1HwfkpcJgVl
O68K5h3WZzzK6yNxiZYKScV51nI2KjE5/ll1qpTvrWDDL9ANMOCjqS8mIW9tEAA0UwyiZFTdfgRF
PWQmZeryh/OPe1e4uqexybT7RBcYXB+soaQuirG/WbcHyaY+pQGRGsRJkVv6TLDnolMrZWjglc7/
14IjhCZonOPjJk3JbtMXn1GuDn5syvAJAetP4gw+fIh7LRctT3ZKWcw+CUYv11y/pqAgjw4tC1MV
i6/HA7c8o+zRypoMCaogewSKgUlJ6gbXt9MlgTe13t1O3F6Dznf+w19nEitDcYteYhKUXSjFmKRf
8UTjuHHSk0UtfJsi79Wz2J3CF+TYFGAjU8gM/LGCg6g/UVyOLSvRLpaUO+19IWhTm/rj3rqXvXT6
ZvT4A2BAsbyuq6/IqTcChgFwjo/CwgMy0kZdPvtvx6VMP6KdtSPgkqFHFHSByTxhv/3541Zu+RxF
j0D1t7R3BLKKgpayejxEu8m0rtvKZzPMmDBz7V70LHbZz1iQcPCFxJ/6stfiqmbAYuLQuVGUb7XZ
m2id6BawmVNpaWgmzmDeBGlUpUr7w7NihcHDdK/sC6it0e+xYkgSNHCX0RzzJUTot72DLhGZLp2+
NgErpO1hhn/2PZjWwccg8BLFatafDkZT08gLknOmUYhh6WFLnUeHzN5CbVoVIjvQqLHbMwOqA8mW
cveMPil7a/7wIKflz5C1NiRFxZpfh2ga22UFLrYjLAcrxGdWKZNCjxxOLK0cS9ieNfUjq5kMS7C0
hGuUTWQ5eXtiy9lUD3wGhAKVIbWxf1bx00xTX72Wo3091J+ou7ft+4PcgYqklrYhb2kxoYe6Gzej
5za0WO5g+sPF1/TCP0lnyqUd6LOTiGkV+yvQ2RSSqj64CdwpP9WLHgE2MO7JZnYZvIEhTnib4hGW
R1NwWtFneejBFZtU8p6yy97YXtmzo5Qd86FoJv7Vtn43alO38mxbPl7hM2yy2B13GIvCHauj8DZG
6QZYB37AvVKUu168RAGqpOAvjb3UWb+VwF1xCb+JRNlvy0D45MgJ5NGUMmgYDZXwsQZvsE0der0E
tJelZHQSLaOAkWDotHivrjdPn6okhNnAxn+VFNPuvZZ1bFBRfnNJNJz9CLhiV7RqmxywppxZaHx1
aJNS/9jbHUFNlX6uDc+wwHteA26203b65MBxwkNIR6hhN9Y9xE2npFmrVyAL0aKoZi6rw/c1k7jC
E1n3uKsFHlLZ29U2G5UYPM3zdWtroMLsVpF0oeTyZmUb97Ywn3HaZDEchcuHpLWCT4hbu1E6vIGh
svJm5/frDzK44RksLu1bzpiIeoHBZ7m387cjUNPSq8qlfGhcqAnEHnfLKDHZM3sExkmv5n1RciU9
kouAvolmWvY0kt1eOAR4Jji/LtsiEnf3JZMXnipb8FRfB3dcVtCkiOBmB9YZAiPva+bjB62Fhvl5
XzyQTK3VfDpG4ATpmlGIqoqjg3dm3wlDnm8np2Cx2b8KczSP0e0CDHtGkwOR+lXD6cmJ/if8oyi0
Adkhte1EcMUIM3IoQte8B07CY6mfXz0DKA2syRhiODJHJyxpPTuulXkCmOOhAL8DpL+LKf8IP5fS
ZplNNOL6hfTLZrFFxtRVOKgtOc0WjKnhhoBfSQe66ze5DI0BAH0OlyM6FBd91EkkIyyrndkg6zmK
vxM3uOnx075cFL3lxsMupnQ4AIVLoDeT9MyLr2OpSTXJ/KUuUuvn6eDWEywSZeC5wGzSP6ZI+Htm
ta/Bc/WNdHs871gYqeoK02U24SvegpbNcf3oOnbUMElns5hMANSuBl0p7SxRR++QwUE/io5m6eyY
L0ygcX0WT+THZeFqmxYh8AiVE2SwF3HsSj9d/GpBnQolEN1EGISmT6ZmjHrhINK8D2Y9FuynIgBp
PcjJNS7wHoqPW7+xPmLYshGZZcQHYL6thz3mjgwgrnDMSPJC4WxhTBjpbNk8UtYwdgM+f7XO9UAm
DSU9ZW96VE3khSiPH96x5tjMTapi0/FhxLQGq2FCccfwm3y1lL06dzA57d2eLyH6uGIXMgBRHQKI
FuxDCgrSQwyBJ/AW1A6o+a4DnSS01q+lTofxwXHv6fafEMItWo4eOvKWe3D7pl/t7r4gcAzAn8jI
4j6qGfVjjqn37eXi4UwUokOnzYJjoapBM0EKOJgXNVwcVFnlC9LON1MtQ6HGz5SHdXX/UGnnPKX8
5dBLMftQI+qdnWtdzO3yFANP4vRJiTrtc8v/IDS9JfNbbMw5xrhuxkHtTSny7doRAeg4YgF6VhJQ
MMyzmmvNGasl0O/N53IV7SZoDe8GetdJwqS6fMhQdYF27EbcaRi93SfysGrI6gNXvXS/ZoT5XAgi
8nQve5bQ5y/MI/251YW3Ej0y39NfglqjYbmqOkGd2TSKTwLLT6XuXa+THXxd1LqE2bQNsptyZWAk
DHY3mmYeDD9anvy6USQw3XLKntccwGRn+kBuUsQDhkxPGn8xUxHQt2CYTtmiWuXLfo6tLpoC43HN
XeDGsvlyFZPLMEPsviHU5OyY115lGLCm4TisVHR6iD+awUx2RbVYYQ2sJr1JkbDr+AaBHIzFgjzf
3t9QFW1ay3T+0eK2bXzmdD7qOGBHsusZV2eAvazK1CYc09WQR1h8pR0MFebLuBQuyc3LfIT1OebL
+lfeKlPvrHhczTRLXW0ZD6ZbXgvMbCWd/zh4N53LaeIHdz4pwztxlfZEWftjzwHIfwiwQkKP9M/D
5uxKSixuHQjvhJqsB5wE39kWDTDmRhqsWaAxdiMtmQ9PHMYWXfSshOi/bAQVElSlA7ayAITgBTFL
VCMOMj/MkWBbRy0EUVKpKZPg3ulq2saF/gT8IdmF5Df3NGA/zPbwt051gXSd0ZQTDyeko2sldL59
Cp+kTA54kPIbC5b9YakqgHWv7PfGI0SlUGU9HdB7sSBIYiAB4zQ/2IDSQu59qC5IYcYNvul15jug
dFrUBR9jUy4bkyM4tUiOTPSgRr2Y04IV6oK2kJ5BVzprmyrHu3xzKXBi0edGBs74hfhkymldh9qI
Drm/iO2KcYopMzG0y3yxF3G9dKK4+0oSMhTbn/RFsIziYYDFFmVrj1P6heBufA0IldQ5gXbXHpBp
XyEDVb9Sy3X1VAGfUKWZgfbBYtZymk2e9htQ/eNauDqbI/CpYintTyAcl8SNNyGZP4UdYe27BP0B
UJrJpGIq5TkfvEXsPxf7nzTHISi8wtm8yqColXCHjrb8MgHnQxVpa4mbO1lLiTd9EgdY8266MMHn
kNmtnzUIxi0rSo7WDn2hWWwOADUHr8Qbf+RkQ6XlPSycoAEQ2RscX4HQqER5RpHwd03rptYIMRle
9gGPOsqcSK+w4UoxTUlQqeeYxjmfkUQNh5aNGnb9ROn+FioLi33utTb90ZzTvwCI8QCTkN8d3WI5
rRapi3l0LjmZt5k2qcjgCV+Zkfh1ExnCTvfVT7cEZojDnozWD06VLKspvh7Ivmy6PLaW+b7Kdx+s
71E7W/huI83WECtxNfPXilflxu5yUKotu+go2B7dS1GTaR9x6WpMPJFv88ZgNZrfUctAbSua4ctb
7z8seCEqB1AhamD9uACAraiR0RKwQlKFNMFk2sUKMlF3j5T849UQXx3kGQDCCgiAHkaQL0DYKTcC
BSz9dgtxcoKIf5zm0IH/wjb9DRgxqR9Q0uFT4u0R1TqrV7QfJo58WFypuMXS5+8FGrQ/6qarc7I8
xPXZHlyjtsNGGELW5MtywQS/GwTv69lQKj1/vEWjenAclGBTzOBypzLDBdBHT00QuCxSUN58vdj/
RfzXLFrINSreILepLT08b8f/TptfNfhMaLyK0+UtkPV9CXn4wAegWiPrNRjo9c5n1gkz1Q4zW+zM
IdoCcP4vQcvU3plZ4D/1IXWhWhW0tMydmkRxH76NlPsGfa7dmZOV4OjJd7pnNoLvO4hwaIeXyxnu
jY+4AlqmxLkhASlowk/ydPv+A/1yn6lvvWWlOYEKv5o+ZYLqoLGsDPaJ7LM88vm1MmOcRhAVIqme
55qp8bPcHhVUbsIH23LG5zGg6vzAALhOkiuRVKyI3hvl0IoltR4PzaG2gcDjxTm6kDKeTr+Y9f5v
oDCpZRj8XYNXVEkA6/nJwxsgrUGHWtuxOMyfxIvxxyhOG9LadptWoiOeCm9QD+avBXz/3i1+qjtN
NFnh5zpBIJK7c653sKXjAaZVusyegryd25Su+nDmTVvUofYftawDRsiF9EWucjmZDQhZ5IuybJRV
bbS9IxloGgP9HcluWaVZwQixd1MSBoSytfV6uVwvnMaWphZw4s8zr07IBGe+I30WLshh90yg1RKS
Kkh+4No1qnxGx7ZGYUxW21lDNnKCb0vFXmK0sNsY8tSACFVea8EJ6tnUHagG3fQ6h6X+wH8A7WSl
XcbqqQ77RuKbIE31ueCHnPrAgSFFtctqVQIKFT8sQsH9CyeWh1pWH/Cw6k76hmZDtKxdxbwFSLvC
PMci6g6O0a6d/yj4WUwFTc7xl+w7j+ICCwf9FI12/GYCGmUpfxH6okTojO0aX3PsfBb3aytWYTi3
0e/c0zqRNbDsxvbk7W0ILaVs7+qQIP9mdgJbXZcfE1e9gIj2cP54GM/qy1rQxg1d8tvJtqRAYELg
TYPvaUlwBRxAhKQm1XWx+bfAqapufrRArhvsUhGRyI+6kw/qTJdzmEolDMd0oQIGCwBeJp+SqDbP
00wvHFlHWBbs/xVBmhvgpv1vRTOpzJr0irWJG9VNGbfTdEqEZF09O96/8O3uOsJy8U2Di4IyyLCi
SyjpO7AsNEhx6lnDWrYX5kQw0Ob9NyQ5pY8joqGQ1y4gtNl9MvqqdvdAMLSSIHkBiwmFnMZifJwM
uiYtbxZbaoVvGfp9u1xzaiSU/6e9NdE+733LhNxV/zIQDKnP/a+meVS3Pp0zTBtHQa81sTjxzHur
TeAa2sYoqoreMurouY3JqP/mXcQ6DreYtd+1dGbjwC0/3Ob7VPMHkXo0oovw1BagOOCVYNL+S8x3
pgxEuM70RoXiJKKFzSB2DkBcV4W15VFKWOXjQNbl2ht2/hc3jO/AkO+x10dYa2TDuzG9AYUYY/+w
sNq4ufdhrrxbvd59d7VHgY96fQUxqlnT4TD6g6CpqOtvmWLhFTBVVchOnZv41++qApj9wD5xyQ8N
ANtbxaPq9Lxhz3Am5Oojts3ySDHFQZipxKqr+WRnt2ZV+NLUMglNZMVOKpxHm819DBA+g/Kl5qlk
gd5mptsejHpe/RoMlhAf9xoGcmAR1+58rGHxh8VAcpoJpngmW7XMsR3GDYu4KJ4mFXpsFEqnaDR/
TM2K3ZRt0VkPVBTHlPuXsz7aAW3VeBYA4wKkTX+LqZ9d+lUKoM8ORWgqPAS+fETv0orfA9uWjHLy
+gbSRkQXflfYGBaUBvePqtj5VjWCmIdBpVvYDnLoV7DDgTsnPcDk8+C7NOE+OCpA70JjIVJ1brP/
DZfr2YaKToyDm0oSMFP1ytIdltB3khthlDes3fNYAVLZd/NeU8tjyDuor0YyNMH4Z1LXoqgMzX16
03JdYqTq+u4xpw5QQuLOIn0SAFUhnVRD3Dd78hXzcqUCbON9GhundbwMjKHVJxcpLbP7SDTE55ht
VPY7JVxUrIN1W6pwDmGHFKcMxTf3DBD/31obzxWdLHHU5qRRXsi0EFnMJf0lo2J2MhF0YqtVIjM/
pqDylWizCyRtafQfjEJQ8OyJWIryJJfPPqHsoudsG/InHnGKptxK6ZSCKNhQ6kRE2sbhMS54Je9x
aWy3i/Jtf7qEaPKosQg8TPIDY3rbuiRLd32j52Dc4NOA/Mi4YGWjjHjxn7wUVaee2yzqKDpMVsZ6
nCv7lxMrF5wOCqnkfub04M7YHk4yuinjvs9JqazcAjmqpFum0ap9Y3F7OQohDHnyBdNcXRiWAhkQ
SRddz7Qnfi6DgbhTDOhrTiR1XVK7SF4Yw3jluWHet5XvNLvu9E51Gd1uzaqz/ZkBHmSFsXcIFnjK
ojHpMuxnwcRE22wF7VgBv2La7M2DKI794t/1nKW8QL0Y0auheThBXq6HuY4UeKhoGfSqdh3G9ADV
tWEXQL7kctvArfR0SOBj7hd1UvIDkmdsaJT8jIrR5F1JSWAH2agC8uFkYlmIFfha3XmibvINMqew
09q9+Za6HwvoFzQ2nlWelbtZUYrmWCediducechXA37cvz9QW3f6f+MYOOdZJ2LBcRxmebK7vZ4G
kdqZgqNdBxnxb+mOk4gh5Wht5hAtwPa59wMT8c6GuphIhSYrAcyGJTckIVx88261QPC0f2P0dYu4
xJ55RWohNxZpVyt+1BAMfuk1Ykbp/jgs1sahZuSRfGONWw7aqaAqHYXt58H4nP+anBbhkXrIDhbj
VRYgytbrMCS+fHr5MreHr7cP0ItPTP4IvYHP6/C53JBLV2lHmjzJevxzL82+EIQvzJPdd7NDu96d
Z3q8QO6AdiOnOrDWypoKe1bz63y0KZhad1bjweprXA4cdBnLDvkhtjqZT1DsCjdHFbPjtPlXe7ek
z0nHfbjngw49Mq69/eWCMAM/hII90zEg7hDNJE7C6oJLsgJX88SbttN4kovAgfIB3vliPdScB6qF
IH0YopULGPXywlfUNhOvJex5k29Hn8FTGTrdZIK7PmfYZDp6omaG1yD8XAlAwaNN8Sam3K5kbq+u
rFDZXM0KIVgDJdsA+vlVXgDkZioURHsFdgPnCZ0gFTuBHe23oZFij/I2Jvg57en3u+OQODRHJSWT
5QOwjRpYwFBylFUm/q0hmDRI4bzE2/x2QTYnqqHedgucd70fOBNaDocRMVu3vWZCvtniaLUT2iv4
4fEuq6FaEVPNCAcLEDYMR2cIQrXD0piy1juY1rmxTo7je8jLeu8KoLO6F9XlEOX7nowosMntB8Tp
3ptmsSI98+8QywyeBv03DSdCW/QXFWV9xgi1FcU08v40+vxALLnu6R95P5asEHpfrZPg5M6OIRxJ
dfW78oEWVl5vhQGzr3hkTPjGXwolVP+5vogxlRLVZVsQ9GurFyGQmj4RrtWJQyxSRGrWz+oVqZPJ
IawLHi2rYph1zaumipGKhtXgpUH9MTSmJvI/6l0VWThAAlyQHqjGLbYMtjc0V8CWQnM+ar3aF1cU
yia7BnKhjfCBJ4GWqWuBEdvPgc54r4NLJugBV+BgSb4tjQWjKsLAyRL43Xt/BN4aLSSV1lfpJujQ
hRd2C/ffPXUMEYiO4Sm2YRk2gLQjjX9ZI9GZMAww1NGLr2LcQWWrN5ZHWyVPrBhckxEqv0hfa/6I
pm/Pjs7SplyscQUY8HsxBb5vHylRyCk9dk9CGUzsRk6otA7T9HgB6BW842PGDwuMFheSsQWPTQQB
qjIXZF86Y1IxLfOICnEImgV/pHuODTUUsdsK9NsXyNxRNOTyouS+duckdvIeQzawbqCDN9aEXAoL
MZSk0JoX7tFw3O/jloTpziyJwU6wARo5Fi/AfYGeecZ7EfuujHrISPZa3b721aaXU7x3cKRWTvYr
+00HPMw3GRvOwB97tREKrhvapKtfl8sCX5pVIV9oyynIUiUXxM1HMzENgClCIn40/VtEGoiXcLxZ
8Qryxfumk++IhMXJ7xMiLxud7GGM6FIwPihWu4ht3nahCTo5M6UwuA2tpYy/t+xvpd+uD0fMLvKJ
JpvxE8n16jQnnb7MiXOMEf2ofKA2Y7+/GifB+f5lP+U0Vlc7fmZi5J80VvO2i+ltHckrhpNeQ7KG
X9dppMPUpkfK5zZHSDfm6D66mN3F0jqOuoiAaiuPh69aWOOHIufhps3z5pEz1rJQyipDrxMnNWM0
gHLNK09hlHf4nBSHZ1jFTxsV1Eu4pjVYDMb63FiFjdRkC+l4dSpQCisWd8zDtOFDdt0X+sFkrQwu
OC/vUyBjgOp+nvlZ6L0RkXPrUNjJeq4GlOKXx1Ez94urrX78uGR91Le0T9Vhb1/6L11veh+k8imd
DIe7LnBM8W1ka41jIBkGAaIO4Vfsm3T/95LDt/afDgSC8sqyJUqLKEQu50jFeB8w91b0oPCa3CKX
5uMNfMQJV/+XPwLv835poqF2gitUmRqNGcaP5J2uK2KX0NYAJiYy/H4vYHFvvlfEZsa8PqHL/Fw9
zY3uf8QFYyrB8g2TnXp2dy8ULUdBwd3JwrqLVhRzo9o7PPwELDz0/COl9uNoXb4bK2cQ+vWdJ6EV
KbDCgTUWkohPYXwzJOjTVnm852VYRKbKWLQPd3Fan5Dg9PheQ7zU4qo/LpqJSlEyVfmne/KY8Cqt
cOjvLaRexhhCZeuLYCmLZVQHjOcdJ3J+uA9HajBLH0DZTYdFIVUeS444+YqzAIoN+EmIRWkXSiMN
u/2ppsYxpKQnc80DE/rxr9XVoCXK4K6LqNknA1mTDSNrbgA899Z5Yc2Gbf1qaKKBlevCjQ5jBF1u
gmjDYZWZ2Zy+VcjBHwEGcwIdPsxDsAE//eV3/exoIZACDHtCGN2x1PRtQJMf21MLu623J9szi8ui
BGFt+0hmnJcEdXIQTqs6dQPOdp2q7akwF7BPU/yl2EB8AWZmYrwjBeZc5rfOKNKKSUWqvCCnCpyw
ViOwgQFm68vcDe0NlYDyi2+lwbS20yZmVCirfTDdIAOjKbvaUbmOXWTWU52MBhVvdnTtFgTvzY08
RwQpTFYUHxVLDBTdY4SEA2EXws3qt07ZJxGzsE0s2/XJI32fHFLrP7h+QWQpxDnGtyxopT6lYRZf
jkCY1zI0q8QytRErAQ4iUvK7dYsx1YQ0YYhDiDMvlAa5rclI9AGac0T6BDo4UVa6uUYUAt3z18Z7
Xh3Y2o2+9uPOHSoV8bWd5/Bd/wGddxcW1aZd4zzIRgXPTBptPVE13vFUZ1/1AThGeT0KCx9JoaYD
JkFw/R6POODxhS/ood/4CSFJE928wOENM6JxIqaJKOhz3KGZkAsoukmb24wgdLrHbJS0hGa5osTt
T6DkpkS90hRxjyuYllmFh5ZKo5YhdeMnLdVyvxD5hdkgCrn6NYOh3UiTlK+mvUx5FLmOBUuowg4F
NPPQct7OrvNbquF/av7xgB7t+2EA6wNC3qr/DqSeaFAcgpBiZzVxwFXocfkhOosZ3iYRCZfkKczm
gyhtY7NzzVjsOkDQEGtkhN77MFvCKKRQvkK6xN1R8kwNvhMokzegTjNtdLCbmIbuMpARfZOh9MIO
uZqMMEl0aPFSvbZuuVEv+8GUuoaoITIWocXeLSeuGXOF33vDagOSH/BO2jxenXATqsZtlWqDokV8
4CB1nX7Gbbk6lmS7Ir/YCqu/ZwfX8lc7QZcyJM/fLiOzl899zLtw/BwEli182mwq0yi/Aoe95plO
amNEuLX6tnozvptKor7tAHC6JFU7jVhmfFaA9/rbAfFA9nGppRMATP8qjcAx+7fOHL0D4eG0iBTh
ouBU4Fom9umL1JqUkx1ZkY+VaQfkov97bR3VYIZup7K6jtOMfApu7KZJcvzDzhpXB1UBkX+JV1E2
QEbCNAgm5gBvyCjnf7PgFGx/XJwn3SsZOQYCpApyO3yJdYPx8cZYaWaHPdMASKof4Yw165vKWZQE
i9svrdtXk+qKIybqf84G19kCLvQFdO3LSA/g3HAyk42V7AXvpm09c1cuweSkqtey7TiHoahyoghx
N5oSfijoFrZMITWPDP4Q2fwxyh0OYzgCy03zmkqaCdspJqwdEPiiAWgTT8eePDoMTivwwEXjulFT
i3jc58u0zLgA5j2NktjnLjZL/vU/Dlb8ZlKD5POVD5cv2AWVoPPb+o0tvj9uzFA5VuZUeCZto2OI
aCqa2Zqu4vquycCTCiKz5u2GgO6NnQFzl0pLbcjWlm8R+0x3nzjCOV2FrQCcEHJxlMU3/JJWVOks
ZmQRma4Ar8IWTYvxWP3SA43eYY+jcDAtMHSzf4R2z1plXqbneFR5q2H/hD95vbF0xIJat6Fkhwq/
lPH0pr9kR/48Z6/dra6LwDsLtYpI485GifNvGVVUKcYdUzPee8qb44sRI4lGvJI33+NLlwk+uF09
nnkXBNCtiTsWFPAxomEuhuRSeVr6Ru4C45lP9sRQP0nAKtWh8Z6nCNJvDNdA5fYeKbe9s2cVhsw2
D83T62G2vYtBUnRIOfWRArFZfYXvPXdQC6OE6t0Yu2ENzGW8W2HnIUgoN1ctYmm33C1dOn0kPLF4
mpY6zj3kjyj5me+8X/ynbAovACNrBPlGGZcUvxJU5+qGVmVoPOUneqLUCs18GW5QZ/CcfEeIo+br
Odj4Y3S0WnNpbF9eADQhnfoj0qE9pjGUd+eLL7nmlFjh/YR2PMZrDLEqY3jdhb1WGKdeHV0iTHPN
56cQwPEG1AwBHIoCBen+I7Lgt1pmhSUmQoHMRSPZp7ENSX5yxbAV2Hti9afyFCgRI1Lw3pWUHDFL
eJMQReD0vIRLRLec5fdZpY0GPxivRdUa/2eWmFtepPu4kZWmpYgUrhU2FivrCvoKi8uOEAylPR6E
MZLntNkC2SCj/6KFdKgu2uehFf1n6i6ol8yAIFj2gwaYeay7WMJqFJvoRSw5SEJMUwz7ajuJBg5g
73D7fR7haXacAal7XpIv0+TLRJ+muVMTNiN5Mb8YGapF3QUAbfRxBjWtAtThwPnbIfl5f+ignKpZ
cIFRX0A9HeO5Rgypy6K0ImBlY5EJdQ4nLIdCDwvz9Oqzg/X5CJpQlZjLf02PHWzXT0jcdWN+nQfX
7OH1qCs4G6uE6Yg9TMfAl2gKOltA3i0V8Ndx5NXu3szNAwWgy9n7tzWWfqDMocHj9O69nxEwlMlL
/pSNxjF3jxM/ai6CTfM8IBsevgWrfql2xs5kfQw8vqDTouf6rZt4CB+t0Xzayb6xaWrBIcHnYH2m
oFaa0UjIttY2XPghflkpyS1VNc7UfOcAGxZf3M+Tx8Qa6VAom60Tn3OiaFmQ5eORywrAohf4QPs3
lL9+xzA1psQpKZ4j5LrM1n1VVj+K49fMYfbVE9JbC5q6Em2uedDfWe71VvJNZ+EfM5372LcHCghn
ZyOecXnge9w94iB9ebZNR1By02q/HHTG01YQcX/YJFMupLt0sRbJpiwOgu59AI/UQK/G7FWg2Poj
nvNrH35RliHLWNRe8+lHxFCGVUwNH35PfZw9YJzgsVhu0ZmNeuCctOUWV8tt+sX3Cu1FH1Y42ZIc
YZnzATQ6MV1fsrHCFsgrAg/FoDLpQXwb8psOPZ+ojiB2QiZsVLTUYad4EV87jyaqBqdJQg9b4Q7P
GgeG1YvGjAhW9lApQz0iu5y/uWZoyIqQvl48BrvcmdkP09tJqbCguBYGUcwNwy/3MzIxaF09dbOg
G6Q0iOm/Hz4PwV83KaSXtYykU4tH4bticZYVPMoJkJl+jsIkH4BobKAFzd/TKqNC8HUyKq4sSFkC
3Ply6lMVlWxnNXouso3/GScvnaEJg+PpCuBKvEUDDGuGX0TEjxz121+I4kGlSLybO5HodZ157mE2
pRX2qvdig5uGVEXy9iUMZG8ReF0xg1fbwTKup53dvJ+NUhc8MEVeE5FMsidj5FBC5aLkPL4nsg/3
6Xptv3Mo5HdfHQrQMpbey6DYNs6EOz/ANlmqxiu0LsaK/c1duRGO8NL+MYDVn+2RRXsy6L0YwFrD
Kr1TTfTTILQp4aJof3qdvdegfgQdwZpnG3gEGY4FyGp4lvXQZTxLL543apxXGJAckMZ5kOPApnsQ
hg+bX++Tw1cH3F9S7g+4CLrBOcAQS+uX03p21Z6s/2tn70ntxa9Cp5HCYPAzIMVMAKCpa/vjgoiG
RVhkhm0VhRWOqM3LnoBuiWgbsg9B23lfzveOuu8Qnz42AFyhutDONP0RSCU7wGJrOSsWr0N+6O4l
/fDXofu42oEy3VcbVje87viKOMwM4jbZ26dtO3kijIdtJKlrwVIFBcDMv5y+BIQBPaEYAimJqS9M
35mAZoTf2rPOvZKdmmhnXeRq7RWf9qUXJZRbO9nhgoBUw5OTSb7vmDm9fo9Fx9ne27zadjm5h/t8
sviwOgza8qkJhKTC5CveUaDOkXn4vAqy76N1a2aXz2656UxHdY8gAQ1Smo+3ZmGjpTPpNy7zlf5k
pvrkQPeVroMM5MQ9VQWysWe9ciX8ImNSX7vocEsUj93nM9H8egO6TasobL+VLZqvvL6j08Pzsqs/
PHlbzCwiaWr7osvGROJbarXOk4hwlrJM8I88566BZlSXGcLd1dO5bgD/aSpLIVOsut7W3IZ8dL/9
LeY7yvBYGGDXI5xZFzOkHqGiQeWhjlSD2oTnaO3MfyfyYxdVWMmtAG1/SQ7SO9uyKQVlH6CW1LNZ
NGrHqC3T+EOLzttMwlKDPuC4kLCuMkZZQnE2Hk4T8HQrSM9uv+Knui6BF28jZLL6YSLv4Mh1t3F4
g/eDrjt0bP5QUwMHtJXNanrTV4WiTBCInqioVCFxoMtFAqJ6RtqbCtQdgG9/0e6ycYlw60vbIpId
nCMLzYc+e3rXEtPVTwNra/zHUe7HvLZNH1CJ1nyeLCgl1O5hH3Gt4VSNKWBbPzYImWvo7IyiHZQv
ZTcuNj+Dec5fFjRelYflXYKOD17HVXLfeTqzNiACgQZ3mOZJAowAVd/FNMHkui8Z0qQthG1/J/zw
SKTtzqDslFtpgf3ZxzNh1/XdIUSp7rR25/1jLxryt8a976hnZYqc81MONr4NsRwc01YcukNY8qbI
PvDq9ibEK4AS2JF8Wh//6bfK/xb//JoYlxC0vRIS5RalVQ0wciEqW8lOlwK5hyfQJm407OZJDohu
gTtnF2qrrseQtYjPR8PTK3xPgqlkfz9Gw+gX0mgEnGzZ+DZeeieXz9titEEc8MT16mbJMbHyTe80
yQhBNLNxzmBVHoU2+WER7W9nFftnd1znEdtO5DK/UTplb0elkm8DiiepvGQcs+JdtN9Iwf86WK6l
jhmFqed2f6sdGeY3sT2eIwgeyaD6YXtMklvNXzRn7MJSM8i6yDcXAI/2iGkfJGfqn0obhCRMsRjw
OpEk3tZOWea13Xyaucka6aygAWfJlcDKsjlaiQ1FIrCQhdgl4Dh9zc/M9wUMAd5iLcuWZkCHUmjM
AA/OqU4+wK8iVGKvntgHWQlByQqRc6f0KbbpfdgHIW9+ZFw+ldFpb1ZqVVHRRL1ygBceeMKypPMB
QhzqwKtcz+95Ysi4w8FW/8rEIuY3ZekYigvJT8k7f9eZsTfALafhozC4PNFqt19K8Z6SLgUmYBq0
VpNxFdgPOTJZ77S7ylF9dV5FJAubKgz0Fkt73G2bLHOYiDn2193MsiaKYAGUkmsGoyC5ML7xVVao
At+2ZPCEpS7rg7nI7VTv/L6979PZRK/ffgx33cfRFZBPb8YUqX1BEX9iJUgmv35m8LZYRu5r7OhB
B9wJVniwZuO6rI0yM/XsL1xmORS+lyh632nv30Sv4+9huwn82nrmDQpevz7+xmN5mdXpQz0fIQqu
Arv1E4Cq+bymqd9OkAn9/wSUdOP64v+BKR/3PuU954da2x5ouBBfar1/gxuqQDRP0YMT2LwSw5GQ
t/k9qS+BnKmwZSZbpOZl3/us8ixXlCLlOBXfdIwwsUpNygprhXJGsDa9C/wTcNNPdxep2u40bZdh
7RtIzwspFmCIMkBRPuKX+0xN1LhiRDEKa1+yendabiCKxPJUAaDsTrECdqgneN7Q9ZVvzs4ufu7e
+rJJmXUensXzAJwoHv0j3REXT1Q48TW5GvJJ7TjREQWgLl1v6iyIXqS9ocYo40S5AI42fJ/Q6W/d
URMhU6lbqmnw6HQKGr8D5Mj0K1Y0mT6Q1SdY7esXNy8JoTECrai4kW45fi7bi/jHZcE1BQrx6Ypv
hybQCP0oEy6TrwFBOJ4Kd2bkhUIYpXDbldyNCDwUa89GgNUttqZs186Scwy4i6W/X61PsHp8um0g
9VfnjHWYTUT2RrBQfAjZght3uBoHPlUgvKPtVuhECsWTW7ZbgjRUZVpF44CM0qypncECeP6LrbnE
3i36E1GP5EIj1g0uBbb2dV6HRagppBhueaLaMhdl2AUzxStpCWuSMtTQKS/YZ6A89Ig6SJq1MeNF
XhrXMq8vFt6Xod8qOaowTX61xRRuNs6dGf470PZokujjJom7RBfkjbhsMIg/LY2/lG7FyAQSXd2r
EzOjUyHLryL/iC8rwGzisSsnjveL/T4TW0832KBS62Ioxn5AVwbmi1kjGw/QKMK1i5TcOhbf+x8W
XNRTvHARyg2foOWO0+SthzC0oKtsXMcmdZR0tnO/cB5JmYNYpfVN+UL0lgLu7MMtFkGJ3Y/ti7nM
hH2t1U8sRt4nueSwuHJp8wF9xJtE/XpyZQe+CtgSnKBVfv1cVio/mXYN3+4vrW4ae8D+oMsxP4WX
qm21F/sn33TZL3pBBixejJFs3f15kLEdt/FyzDRo7w+HQZ5dE1GqrDW6S/47mfNH7662s50qtOce
pfh7gPe1kpm8ceGyNM9D4nd87EMYlLhaRtm3sRcVpoIN0P2Tq3eA6X+phxQvOsApxw4l6qqVhk0i
rS8Wa7AyzXPQLo/LK/9gYWBscUgi/xdPpnc1Q9DHYvkKbID2d16Ub5GMoNLsc57CEpO9+VNMbYAM
U7qIw4J8YYQjeFsp11iJPpDv8vpS6+l3oa+k00rJTIid38Usc19DLot5YVOxy7oiIFe1RnnEAwxF
dK6CGY4fcnyu+jCHhZPQghhdmZo/iAXD9eGoMg8DgXTSTZQAjyd9D/cQwhcuKRzGBf84aeVg405p
RJ5DIHyzNymyXxvoWxGfvUzmvdW9AKDdhvTmsb2aIx9gyJeUyumOAMGvO0lNCQqQqYCh7RNVNPGW
t+n8tFoxkGb9Ru452lc45HDlGotUvq0rDTp58tdCROK3eVLuL+kCWlGIUWpRCk/lv3W2rBq28Gsa
weG1Ky0ybZ9Og4NSqYws0+7fFu7y40hbYi9xMs0c6kGPVjEmRS9ruoSSBaES8jJ04pZgHDxgeziw
gJwMzfCgnfXRIy4Ww+tCN96kA/6ESvc94mSEvEoAbyUjkC2Jdp4XDYnCEF8ysTO2hGHITiBxhLKF
My4Ei4GkXrFykeUahyUErJhDhCDqd0+FM5ptwThSxvtBF9I8egSzuDqSP/Z0K9RDWndZvltiur8V
PFtAEDFNgoFI6XZjnIEpNy5Cv4D4bfcsEckCVG1Jb1KiB6BL3rS2lM/d452Q5Ubzm0vdDY2p1bAU
49Ihg9/TGIO8aMX7uLt0PfYj2/LfYDRPDGfM1HN7QnvGIqQ+3E+b7wsp/hssOodadGF4uStLWnOm
zuqP0+7XLp0x0nn/k5DPYR9klXx/Jz+SuS/6hp/ae4zq84YjytHvlpBj0W6A+D48MHSziPTnXhv2
GH1GUZ3r5AtQZXyfDRMhXNJEnCvyla4uczqx/xTBkfjphWRuRcX197RPMT0zzVG11Uf3Dkp8xLp3
Er1PI7LTGbE5wfgzqMP73y8oCt2nZxc1bqLq7UTsFn1kzISi6XYuDxcu7+IA6ERT9dQrP7gKX92y
kRe7UhqQnGPiTO7ZgDY2iakWPrGYkuSrK10QKgCTGQaVfan9wDYBZzko4FRY6hvhNBfp7otU2J6f
3bADuuuc0Wdg/tsT4MQJjzLC/SxaLPxz83Ka7qTOUx1LAX3QlcoOQIxJ1ye539Aw8Ud+X37fPcGV
f2yTk8SPAUxXGofNA/5sDw5SOvFTCVRfl16Po7lb4xW4l2GH0Re5w5owEyIl8uDSJwz4747mAWkZ
TDgkSI4urb4p5YLxpr/9sriYi6eOtYDqHRUJkaCvXZGlmoutXDoYFTCuHHTKnNpJVr0iOWbrxjTU
FQzo58XpJZxSizZBd3dTVGIYQfRqVtCn1vgC+IWs/U5+i2MTcCNKAgFD4IzImCSX/OWF+DHsP+dL
FxKp+MI+8xvOKcKhw2TLUnWrZPduufT6/psJkw9KhwtMQd9nUAC/DKHkEHOi18M0DeCAO14GddOF
+FoiQHjbFqky7quH0ZTVHQH0pcSLfG0RnaoA/SXyqvFUq3JS0cKish/zbt9Cz+RZinxH8F1cU7Fd
XVB3z1X5qzi0FsRlIbhkgUFTl1uP8Yk0j6XBd7bxwQLENOArNIzU08ylG8K5UJpHnqlNpPU057uY
eqQJCKTdSEOstfeDr0zibi/D/NcV+C3PUWyGsFWnGHoQa8RCAd3Ng8lmZVWePZ2X03dwz0rUlzdD
EB3CXdjXr0uHGcneF56mcymPeX6cOISkGs99NSlSW7ZJznyXjtvYAlJjlxWSoDlct37c8bS1D5Mi
sDiFw5vDs7Oyk3wAmXzoyPyNX2l+cJLakrny1brI4A8PbQDHtUzMaS9OdMLzBwCMj6T593C1UFiG
delG2mhHAMi3XoLirvea3jTpsb9fOasnr2bfFtFXbTPanzWSlSZ3C3pMye7HaLkdD7bEzR2Fnm0V
lpKcWSyGLlbHncc+Mhw/M8xB1HP/Q/V52Jac42wZHy1KyP4X8EvRLMX14EkTWd58v5+GA5A6exuS
dRRNAtRCRdgLHKopyq0C9Ym+Ie2maSopHbRRSpr5fWgz0GXahL+8ldmADGoyxv9pOBYoU/Mtcxyd
H3G51f1qyMj3O2W3sB+QTko5XFE4ybcH5zWJCLyQkSghXrJIrW9wLw246dM0QXoq52zpBxel1THM
dNm0Cbj5+2DrZLVR4Z70XO6HQF4KopLq+8vqBo3xW6Wf1z4/illTWt9b1ybCgy7Uk+sKoccKfAOb
Ms6WbwGww8EZo43PThUcs69Xk4hVLutdHeri+xFX169hhpQv9T7o5rRdOg6YNztymi4N9MaH2mlW
V1yDlT/aqhy19bNyf5rp77ooIF/3YE3tOUnqO5wU3jvxWoOq2bILy0YGQikf4U4bsue24yFeHW3u
vuGrweYB6uqOColN8quZDcpLFc89mjLGgjTbazYa5uKf29KAPM7Rvs/+LXm+xr8+rsvWuKaOj7Wj
EXv/SG6Xa2HEoiXiNGtiWwfRrY7Y2gJJ/ztnDVVTLBzSBZtORlbQuUc389GnX+gxo8UTdHZBrM8l
rRze/6FvbB9c5qxYYo8JSr6RfO5SVyvkSoOlZw2+2CTr9B6+FpkiTpnu5yADpcUJV+QWp6FEuwf3
/gFS3qfP3ZXKEwiqmSyTRsjhVRrHg1nItAcHNiO5fZKnz2Hm51smXORkGbPlmfWjIEylKGVSK7Fm
yGlbbd/uASGoTnihy0aJmUF00iS5clUS4+eWfc0BSQBT9GBX+WhdrF3PJesHBQHZ0fy/0TYl6CXb
MfJ/bzR1ld6l1IsRGhzLttrTk28XuBqaz/GNMlkMr+WIMn4whdIhLGtvmkUc3stMV7rYSamvS92V
szFcCyzPDIm6jfPv4gBbh/Bflk2c1arro/iHFDhkZhUq4m+z0bJkRNxLa4xyNcs7TvrR+x1mhskd
wBY2aOI3TJtn/9hfiTnL/wnW2BTVrONlHTkbZau8e4/Syq8918h4y+dge9N8Yf4LSoVSWeOZY7TS
VE98t9ND51wYB04U1Vt1FkhY4Rxk5hJrJi5gaAQBzs58SXSUcH99TnaZLj/TZ4ZXEzUYjUYphWrS
E4i8ovO97SGcfQYKkw7WTss/LH3db+VSOX4t9HJbKYsmYYBOAb82GSwMO6sesMAAAV8Vv+uqTkUF
37hZyCaUn+fTpTNazCr2J0w7krEs6nG+WW4XVBeGERPVD/NVHTedwzMdX8eN/taLLHEK83vdGs6+
MPXu8EWJFIZftmRTX5o65MJUNOkarV0pLrWJCpSND67FH/qE34++Ni6LVMSaJqZaL8ELXYbjtkPu
Rrat3OUE12Eq4G3xj7eo2N037t8T06KIIpHUx34fjzihYT1z2H5VPajKmQqwSaNjE45EkZ1H2ZPr
/AgX7I6djDSyn3m+R+l6iZhfuViYFl3Q7ymcVQrNY0vRGJlLjihY2R5gUNrxW8plQFsmfxKlJDZ0
nlTEL2KcS8AUqhvUEhr3QlYAOdwQKvW5ym0oMz3z8CEhxzimgbBhex0AKfvw59vkiDWMsFVMVJal
rQJn70esJuqxKaldmbRGgVKGzgMPjk8GCAzzt9dVQXQwbKuLmk4PxCUAhPm80Ffej3Y0omJqzsuz
uPo2shzYx7BHfXbsSUszxvcVgdS1nqcOd2JkHNoESFXgk5EKSuixtDhtdvMGgyFAZfmYx5pc5MLx
+HW5o2FO4vWN63R1pQ7ZPIwcljgThq0Acx00LiAsQZY/9VPHPZZs6p+4yu6VFccNNgNiJ9WsdXQL
I5+ApMhaSmJT4aEm5XlbVJwrD2pqgPtaHvDt2XwqIhRjajLxUmTZr8dKhSRsS8vXDOvF6B2ly18R
EQH3QKeIyYTGXXGqCouCVKzYN92tze0eBKoZgQz8RBTTOkLthS1ZR05SybSO1ahgUgxandZqeoVP
OB+Mn2vESr8jxo2vCEIxqh1aUToPo2O3/GT5ZjrFtx7p2UJ49M/V1oYRm/mG60MMTskWjetHg0+7
SF8VMA7XVFBm9fz9VWckBl5puI6UCusLLFOutVvVDO3pXxszgw85qSoPwq2yQB9zwcxTAM3dGuEn
v0WFYiRjaAtWx0Ms8pEtWB1a1fkXmxWYood9Y07nF5LalnsM0WVbOedDcP6hAjMV+ix1EcbkGJ+M
2JVI1c10wV4G1xpQ70UT18ZavlfDdnepTTmqxY41OUM2S/QkEYyhSO6bZeV6/MoX72rDKOHhaWXh
m8ht8gZ2qrTjPcZiHzwZIkBpKguQyTNQ3gEzaTIotulhTKII+DkVNR/K74Far7T/US/rELwBoQHV
uvyQIU9gQj6lr57Jp7GkawbiVVzp37iqbzTMxjv21U5TGGLWYBa3AMeGKC/8voFbfC1gyXnQb9ON
yaEQbZg4cq3lGPXSEiOwHMN2qCFkZ4+YqEHgST8k8mwBnAJ7Pnt8Ak32MuaLLXyljedVFkeAztsP
mvmMW5syByAs4Bxrv/ditM7KnSyHRGwBwIIWwq+8nLzzOPW7JL7cGjFQD+jNZ3Du37nP/jXDieOC
STJ7VBYPPHZD4geFd2tZca1joBUxDiMXN/kWMefGRc9JShUyoKPFGwYdGlm6Dnqg9dR/oAJQx2/h
NE9Xo4eSUuDCTDCm//m3DEhgoGV+FqDTo79nn4Q9HsQ6abU7iEjBxNM/ejC3qyEsElkDdLHsfSDQ
TLW1D4pl4SX8llTfCunimy41vASEYXUjveiApEJv7goMWsYwExj76DEbUH7pCfrrFafs/tCV6r2A
2Ky59GNVj8yIHKVx/XDOvgHy+8VRZek3Z400wmIqa8tpi6Och+BBKa98vLulJGzj1mqLtJXU6pYS
hPli7zP3yFMTtk6XNdei+0OUg0LXvobKQciRNka0MvWY/DyXxKqfe6AjGMrJydcdb7wOxSFFczY8
ibfefSJzCTaU/ZEJrmA2Vjdo2OsWP0OBK3HQflcGnr/6rm03jDCcuI891OiYRraYXSbMQZMbpHU3
A0bB06IqaFm6sz14wLNSWG5p3HSR8+tC+q4lhvFC+iIgBCANtcjObWufKigeH3ZzHyGqDSnCn/tU
nxJphVWBE7BG5LzeCZBwcp9dQzRHU/dMdvUTWhlBI5hSGQGxB0/zc5/UsrFM9cSUFo72Z6e8KIGd
Bi/EI6BEFHr0vd1jyznyzelY5uEkp2qfgGg9obPxyY17TQTkOp0YtawAvKoSNeKyZnnKZKPJvPOi
lROx/bE0988mXeAvtfc60jZzt7mK2Fv2e89M02DPPceQ/77yAhVIUjTYbWDSsS6ZJC0VQw+a7mcc
vtZUx1eGa+AuQJekYYa3UatiAn4K+6QSa36hY7j0jpWG4yWRCVnzdjCHEb0kMJihbO2GOxHtImaH
XgODoyYRcskhzHFt0Y3qZMRywh2ZJ1xDC961f54J4S8bymn+9PADgaPcYA87Q1HPQwq50rPiwbWE
mIqh7TOYpbRT/YMKfnaoH2FzXvrFs/g+0XN9pvcphkAPHOKmPljbouPGt5q1+8Qxe9aUoYJDWjmC
dQhUTfj7ukHH3FxgAIY791BwOUooY9/VMEYCNNZtcVKDBaIQg1QkAxCpA10Z+1FrNMii9Yttq8I4
JCNZQ7CtNFFzI6YG4FkHWigGVw0lUrqE7kI4Y+RuF1eD+rMSJ1gGd1oHBAzOuhmUp1lNVkO9XNIo
zL/DaXNu0jhbEiSO9hdSrtrCTdz4JMtdYWC42fh+A0HtBQGNXjtjfy370EdmfttzLAw+11ww4+8g
tiJ0ZNcPO9h68mvuJ3avrSTsdTgkO9ZvnXv7bwvgmn+OQvinTbqyVpcv0pxVK66lR2pfDrDbqeww
bmsFBNuutKgYwLlln/Zh/uabJS3Z+8gn87f5L5c2YoK60mI0cuLZGHDNIxXDZPfT/mda/0k/xM4c
1dsWf6Ny5jCW/kUMu1tGDDpIl0DNoASskTWDKlCJU87GVQC9u5ZulYVDCw35zPXDsaxyZ/GzcNzB
Qvf2N/be5/M/oG27kLu3+3RqbhspzoFt7fnulG0VjrFSUlEhFFuSa/1Iwuoxr8kYNGXcnzlxVUjl
p5hHzS1rl0hp0NkDlHKUqfiminx5cfmEwnotNTyrC5Uf1kvZrBL1FqeUyC+/Z466vretpjsok8pl
tU9Io7cooHMp5KexZJDSn59mdu7K4Yy9nXrQfdnTN/U9ciaf/sXoCJcHpHNWUUXXMVg0F0mR1MsU
ZZPp+yZ5P7P+pOPO6hSPZuikx83A5qu5R1g/wCDfZRjdeB4xRDgLNuNZiMmNNcqjt+5W1f3BUXty
UAUudMl0scVBTJ3XpRtILDeRvtI93ULtFeX6+xZP/0gO94d1sHXz5sEAmCYWm6pdelycNDGQs003
f4GvhqQ9Hkj/WIEVM6dwNpiBCoz2J/szmVaZPK9pVsAqW80zp1wiE2OIrt+LUmop9Qn7wa7RQn6z
CoHaXRzw5UOtw+c8nwfGSTni3lGT5CMxewI50voYTgzuhXjNOt09HTyJ73/VJHbew+tWl7EH0HVm
rsCmMS2BOH9BQXBpWtaRwDVfTober1ydkJH0d2Rv4fZ2xumJE+OR9bSRCUN57ro8XipZ6YD07+a6
WuOMGrjubyX+Z6nS+7hrxG/RU56jIdpU89RFrM4nj5tWBN1zxNLT4uWokoU0wrADGn84K2fpmQKQ
pejerr4+eUagNdUMSiNpUShKXDWtKZNEe6m3gq1SOysrKjXdqblModC+EjE+IZXBoghiH7QMxdof
bMpqfkMPnozEU7v1SnmfvWMqBiv7dV0/890iFol/PbEjnzaHHIdPmsGlNvUu+Ey33YuJla6NBosY
GBhl+Q3n1NsZKmUD4u7w+5FjYyzTbP3BJIgYMdmeY10RXkgbV8stvPzwK/2PmvbFfArUcT1POLs7
NT7+KVYWHE4K+kHI2FhgRj29sIel/VG+rszrI0oK8OfpQm0poEKvg2tnVjhwJ2ysJ1gaIoFiA7r0
UqCoU7QORBjQQ+GBYdl1Jf6HJWC8WmdnQFaUTudJiJwYc6PfXXXpKWxl8a15hArZhW+zlEFCU9rs
h5SK3EOrAKpPdbb3FdOsjQUjniE2FvT9fCJI7sPw+tgsYhT2WLRhEADq/s1lwtdpYjiGExAwnwV8
4CTTZNHErDJQ3qMKVVmIAIXajLfi9nAL4KnKpC1ySim5JyWYcIOkM2JYxGXIw100QljZ6QhmRmb5
e6+H9q0WW/pUe8K/GIz+JNtZTAk/4H0anm8x9SRCGRvQZmsg0xN2QG/z8oAyTCivOMHRiHFPnVDH
9wio+YyrgW2RBKiyiqygrFiX6qCahbTzgZNE98Ed1pzF8tiJIQDuuXDKCGA+aw+s4XjlkWKTXZ5t
OrNeLgKKrkHcbwNa8XSSfxGbxqdqCLcrWipFFFnI+ReaYAzULfL/33JyBM8H3Ymuq7QiRTw9RRp7
tu2LWkYnKJB7mTrvgVUVq9twccraKPOn0YaLaqrTb/GZwx/qVRlCH+J4CkjwdTwXcSdEgPyK4qsm
HjqkXbhHd309Orhc4MiFVOG5lLe/HV2vbC843pY7ZywzB9tMLVi0ofa7B/l+eOOFrutO633K/J24
U7Jo8+QX4CGmLHrEWO55HMgzuMm3C2Qo54MuwjP3W/a2WCX9vdNBl5bu8xOUnoQjyHcM2H1hU4wM
7/zAOxp3MPssHNa+SHf0ZKvMaFP2lazS3DjCGbWsjSEiA8PvDwE9C/5iYdpAdBDvOk9muc7nkON1
sJaeu6Nznium8tMXJiSR1OTQXGRbubfSrf6LjhFW/v6qP1hZZOIql0mTqOujiIi9Sapdh43n9LMj
3+NoxuP81U5W2occ8Y4txPy21HuwWAI9M9ExZVgWtgP7FAZGwn2YnGBotg0B+xXmuT1uCVlbJ4a+
Yg6BskdRGPHZ2Ixf8TsMHwq4sJ+V5wUFOe5kOtdLP6Cy0Tb285VQy2VD3RTjdKF1dkZrfYpcBrks
sreW0dMW/fCc9Qkx40zY/96xEER9rhwZieZl4vRdnjMf8TLJ8WjtVRiBfR5SWRbd+HEvCTNIWVgX
jUfnODjBbGv2MULsuM8aAASLRVFPEsa2ZC+YnwyH0ARrAxG67Tpv7zK2w9AQC2h/J6NfebdqjpcB
KEpLJ9czE4qPtAzugRl0HDvuknuP+647VXugHMXPM1W/vyRNEvIGLi0WkjybnfvYklML+nt/DAYQ
eZ5AhK5TeC5PP7L0uwhIA0k+PVUfF3qrjRyhZaBqULejF7lcfG5lE+pFxEIJCcun0B8+tU137CAU
WiJLk01RsiJGKoSeK1SlDj4YfYqvL8W+FFignK4KtezSCsxFo6uIJlgD3iEbQnomryi6o8vWocQ5
oG5pVbumQwDT+CR5EuN/y4m+ppghaCsaf7QkJRnxAfFxMjy7MVKjzuh3BAMDhcLmrenzUdypyJ7i
X4LXQK0V6MCqOBTqzu1uLCuPvx8/ZSiVOu/WLf7skhizyHdJmN/X7R3LsHVXv8GFdtr/WBLCXYIs
TiXpFhm64SCPyEhCj1GIt0o2GHp16q8M24klUSLVo62X/qKcUKgCC8Vdp3PfLUU8hmvomO3Omu3o
/gluKM9ZjYDfoCNH4WMhVPHOd/nUuHJOekD+W25P1DZEJNX6/iPgmeuwUZPkU064cA0wHddEXNd+
ey926w/EXi0Ow7Qu0eQ4SQgFfpyGyDyPJPE/9dFsqQQ41gGiLu0LQwFlmEfgpmROWaW/OJI8JNgf
eHemESrlu2eNpPvd1Wl4Ooz1351o2z3DuOUXfGci/9nj4VzwGQlASlHlJVZ69ysOx1Xfc20ChMeS
sZaOMfio4PAOcdE4N6gnBaDrI1874KFs0YS9xRB8KHs2eNwNxH9l5jUho6L2d+9Najxk0EMt2/M1
s89yB6s3nleeFh6rGLunOD7KX7tGeb805YQZFLQrG9KsyYMh753ta/f0sJWIaA6rEUlrvk4KbR6t
BJEOPHTuu9ZDtrzj/aB8nbLw8lK7+XcyFkDJAIh1ERuikAJUpp+ukMvCpWv6zGy+mW56eEmqRrz0
oFnMl9lrzbddZIJMO4Ay535SlOPRB/HAs+/F20TabL3A8oSp7GH/vWDkTKQ1jbPsVLYenma3Az7t
XDpikmoifDs3o54zRGclCz/mksmchGdOJBpLtcaBTmEFQS9F8x821vtRVxJZSv3wa6eZ3o6Aaytm
XQhjrLuYz74gMrzuIPMt34f5yLuIDD/nKXzBvo0VI4WIZfjc1sg3alxAmPXdWRaNG/ZWUw4ns9Hw
/Hc+YlOAcNrNVTa0jq3q5jwQqZHcWtJMSEioDVFm7PLLUXOHJooOFkGiveZwsiP1gFQHFh4DMBMk
k8Ga8UhsFEunxJWVy7GA2bCERV2QMUYVyeNaJ+oKs9h8VjKA8Nzjci1AKaDDLWod6r+H8BDXjI34
VVssIsEAnQ7F1XwWF9EFCeUWkB0JgtuKkIdX6C04WfQkfYLOIALLiR99SPzph4biFvbEz/Ifc7C6
NEoeAQsHPfPvkFtXdEI55VKe2RFd4eOXWaUwX2qX11GEOEzOr+iHSZf2BlbJt9RiSwX13YHI24je
BsUufaV6uSDSRO7X1Ik7I1iLw97rbMapLeP4ags8vs0PGaF60OYCAnYlHVm8WrJjTx0RrYMFiLst
kM7K7bKgYEQ9ADJ8JZ6SrzKxo/s2l07oMCfZ4w3nB+MOVingiPFHGTuWqtlF1xLc/3TIQvhfp+o7
aHhCgjYzGcmnlHppTXpVa9tqtDbR9+NObzZCgDrd5wPlVBeEt+2m3IdcV47SPe3DOr3RY6zVour1
j2B3wYN7brgL91XGse0YWFQYWNmeJ7uNxIIe5gc7jvBukB0sI8ueaXqPJpsqH1lxIdf+ElMvVuy0
+uBuuXPDyiAXVpnHgfCJcW+vjfS2sw6yBcL9Lp339AHnoU7wXj6opxE5ULKhRf5QJdYmEhpnp4rW
m7k0mEELgjtk99uFiL809CLX997PiqcRii4nQUxwVSpr9fI5KH21g8zSUSqOLiRFXSqykEhiXMjM
oRPtPNBwdXc4eLHOaXM2NhqEnyGFXfGW9eYcBOO/JmmUsYavMaqujmxgA5BPSVHqKW+RQnVnOryx
iqEFRXYT5ticF4xYv37eiCZQ73vq3ZX+ETHAEJ95vpDHUUgfRVAzflhL0gPAtIAq0z1xO5WHVIHn
Qx6QwkvSWlHGV1pe2FeHaqLMvqMwSvTlfk665OkpLrcSZw1ISjLecxho17diORcd06E/ACTRNvyG
2VSUSTUyoFx5CXWFigsJ920geFUIcfrBWfXp6ZAW2HF2EI1GnYOa9wzFzTqwXSVXAbDzsmqx5GWB
9/oFHvbAF2q8qqugBWVQRN6Nm/sq92/utYNzrRrvZ5X9uMiCyhb4WCKqYJ/w1ClMWsBc2XGx+3C6
LeYxmxer1iJErXZkCw5U3NZ9NOB5bDVoqrI3DVmbi9K3dshFzXqTT3YV/9DAFTqWJFxILDIqdyd5
KpTF4g0PKvghgImQBEnLATys3GZ/UmklM6lZzvtg1qtmIWIB61TzuKZZSIANVLRG/ddR27QEvrTN
nEk4s5AOhprzlB4eSHlyYnTuFGp85JQBcRtsCr14q1K3qxFC+kTciy59fTgsst331bunae0+R3DT
gNnGH4I7fCwSRc/bmRIL3QxKiI8vAFBq3ScDtVGP7CqE+WkmN/eoQ8tIS/UMEgCxKMOksVsvv1R7
xqabFtfNQAdSWsMRTSFlvvzOp0J/A8UkXYEgigb0a9yMuwpnjMZCDENLJaIMl2rdD7mqLGtU6KiF
b1jWXq7a7p1MStbqDkWDVYwHe0hsQbZhnQn+4Z4DRyRzuEO3rfrDikUb7eXhUiauOZfmDk4BaNSV
gdzBZXwN+4pFzFC38bqx0tkwcF5VtLEYn3/v3LDGRxui69W45Ge3dsVhqOul9eRzr1KQiLEZRNTS
lEMfZNeZ4eSTCQhN/WsEBxtfxHVu3YqwRhKrlS2TcJzZcskkpkgZF5qrK9vF2lAS7CsMj95Pitu3
cWG9R7OD8YQY9/QmqORqog8P21g0FMGvdxeRWiVNoyXfTSyxxCmwPm1al3ygwoadBoQaekPVETDA
EwTIxkqlhtgFewPsilMMYyG82UfLmrhpufP7XL3Sdxfvohnxdn8Ov3RP3bUb/m/B3qmVNQWrWs9p
MFsY4u5rfCssmPCDYsCBPIaniLLcZVq4t6/lgdr5FQ+u/zDVFtcwhUY3S3QqOObgyrm2e+rH4HfP
XlnfMgMSXvkP24AxH9R7xTg4R8SWO6IFw485nYXVbwqGfUkA+Wm8iNbpGFLWE3sjxahH7IxBdLHO
QZk9i94j/x9Yph9QqgQIQd+DPLvti+S3iic8uksuxxVw1/TAcl8pu8WYh0S6xL2PFNDKKn+wbXag
+JZkTmvL9HN/jpdlr9L5H8lvPpZ8yVFrJr5mCT0PbA0xieeQq5oShojcuGMxr3ogy8AMFL6DPe5E
GVBDtHhDkK+b72RZxZODzwuADrVTuEtRGMXhpfrNAEscup8gxEOlRhVTunKoY0aFOnLjkHl9LI4t
E1MWxCa+EYZiuMSxJTiiFHxJDD33LQK1IO1l5YzJEnez2sfFcuKKXDXERBCLEodExCyWwGBkq4zF
cQ4xoAaRHGVH93vZp1tXJoHc3VrJQA0LYA2wORh+vWzotHsG8bbvh5giPC5Ovz2R+7SL1ZU8nQQl
0LdnVGpIuol1Z0I/RhJ9leTtlw+6XVZqgT0mX5lEfTbV/5PbGj5KkwJnn2uxcIG0okYbZnqYRcWI
oDvLN3dH58AKqqMJECIewMl7c3o9WBXAmhcToU9ellRNbqc1pQ3Q/HwveW62ce+7/Ir7JO321ePS
wiP2CRYoYfb+Se53lpE4yngH+lYIOVlLi2KCyUWssZVDFEFzfshdDQU4jp16CrTd1/tB2Pe1dGTx
f1DYLrE4MBFfTHWismfs+uT6PXl8iWVY/r3JzAC3n+ReipATDeD+4tWph1SN4G7UDw16LRNkchon
+XtXyf5S9Sgue2AnkHYVHYdK6A3hRmy06TuP2MHEpEplf/9JuhOp11LU3MqvtGngNZ+iV/6MVDj/
bpcXU9dopD1mWIuHNJk+lF3TBdMrEFsSr+n3xDd1tHg3L8tcIcPJa/HDspoJWYOfp2/Qypj7no1P
DCOVwR0/1GuH+MevkKWYPo+wSSR2DrTSAoMfKQh4EfrlimqnNBG/osdy7KXGRXJPDbaGeK+ojwIk
0itcN95EEUWynz4LjUvZnEFu1WhkJsHPP4Tx3DLfSUspjOtMhiat28n3CfHQ5QodpcnobG7UBl7X
im001NLtb1l7vDev/snIii8o/Ml0acSER8iNG0UrKuIhRiUkoTt6mAlt57Eexkdyy1wmcjsxGQ+2
uoakqr1OeJrhNZd8f8Tz1uX8UVmrvt/HhwKV/GEwpuC7Uz885MZF85pu40MkJTrP92BatEhE429W
3RyhpuHZjDQBRqMnvyQBcG/sAI6upBXslDygxuV/4RH5YHKOW2+Rd66OxxuWSorHY38ifT5dFgc0
RoCPWyfIMnqbq0wqsjPNFt+zuF4cgzBOKVq9qNIVeUYg/qlP2GrUZGzR1y1DWYXuRnVdkh8CxK09
ZyeZH7Ms8O4IX46VomIztTNu/sv/UBQSgtaNoif52aEb3tXzxo77My82S0R6k5YrOohKtnb03Bl7
MU4W3s8vZN0CDZpoGdno63i4uvpwm6e0WQW54nZXuOxk7X9QHWN1lW3k1UdWxnJUYqDBLpBkZ9HG
z5h3ctWSIEPeKBF4626I+tJruurGHByClEkavzAwY2/Zm8aZUx79OuosYGIi44fjVmIht/ShLGf/
K3yRRnneIiN5NOpwTHUiUO/+lj8cHpVs+e61h9JZVRILAlLtq/ogutOSRBH4p8ltvtExYaL6zmvO
KiKieJEjMTLNSipn69MR9Ud3KNqGvJWWmjeX4ZBoSX4FsxaLsXa6BDWbbLFMeHt295ZLgQ4kFg8B
K09m/hNE68NIHuHIFQmlgOQ9z5LWyekDnXmNkrn7u+1VD7pPr4z2e78nE7zCUMViIDWHwYRh7jds
X9g12RC6J83xh5ICvwbAg4khgzHfd6WhwRWHkpHMyYwYVqBRw0G/hZESKVdULqyd6oFnqm65wgyu
/oLGsdz79UiAAaD+RESiYem7DVL7lBBXS8LfFtodlRCsNYne28VNjWFEaruL/ZxdUh0A5OZeFbVq
NAM7W0bUpJGh6lYxg5GKN+MKS0TUGN30nrVylx+IhEuh/2Laf8cafGZY/fRZ84KcVPYsNrMcUQBT
LKI7f6vXHOZVZPOhRBTVldSBOEBYTyB8qeRCdQvDFp+ftCM0MUQr3R/6rpHyUFnlx8tdX9NAkB0k
8fl3nGgLHAQfF413pY1akijVthwuP7qZ+gF/aqfksqwQDvB2vJzBodDBCjvxQdkPVEwpBECAR5L0
UWDYUXxAilKh6Q5GiPz6C5ehEq6JwfSmdwFSNJQ6AHBo0+be7xqWb7TW28VXS5ofPY1I7o5rnfel
A5L+ev76MK+GT0WhOetk3p7yzlAdkhLbqob2eRVe6IXBg+r/bcknkeS/NQFc6ipJSXNQByUg6dHR
o93+tyPe8a1CVorBUzd4U6ep8zIBoyE38/laZBLWmVjDVX4aIwih3Z0E7WY5oztkfr7OWpA9EsZx
C2cWsneBtVDUDoi160ksTqW7HPGmSLcOJ0hLkn3oT4QXhvXDfHrAE4C6TsUnUPKQit6sqoHGVJ9s
ljCjlAp1PigeZeBmZROVR1HCMKSE59Q0MUekTWGpoMyUdxJ43XA3m0mcZzUq/L2UCcAiKYbHQzd0
dd8lNufVGTLM1ghXLx8kV0Ip/I5do+TuqxDH7AYxxerNuY+5tx2DqnxUvaQW/6GDI7sudHP/9jRi
y3vPsVLhi+bn79iYw0L7CjceAdWp7/eXueo9OKEhAnPk7fNMtRhiQ8ef2JHdsgAeWvTF3/9eyupO
qOuJ263qn8rdQvMa684IV4BOXIHB40AopMhR/qhNHUa7EvNtNrvUvupAjxt8GlwP00csCzvdjBGU
kN70F8rDJbalfkdD3ZEDsOpg2FM53an1tjI1DWD+vuPZkPapqQADiPcRoJfgBHWAjBweIfDmTjS0
OVI7qOTlnoKR3j+rMxMJ969d3Gemt9bNJacBI91lHroEF2adiBxOpppIuvF0wclkGgKtcO99aPA+
EzUS+zU0ET1iqjJEiXQjWlZExGypHLVpBs3/PXov3O/YinJQ39Ilz/I1CXpO/k8wjsS58/nFftkM
0i8RtD+VDaGZdMy0J6n9QZaCGMaxNR+KCx8hOLyG0T27c/liXpaRgD4fxnfx09Ya+IFu7h6ZnrcC
Dz6sBseO026/aMUWQoVkM2xPzRTT0Y1flp6WiWC2BwyQzw6ZGstbe5Tu0Fw9xsdw9s7Ub2ZOqDQD
KM/wLAMxCjhxD8hrGsDzPCL4ZLZBm5CNESJPSFSkdJkmV0N5/k1AgVhZC7glhSq6WoQZjqFTZ0wX
YKgnv4XDw294tS893739k5uGl2rN2v2C92Ee9MBMz9Ucpc5ZbynlTtFlOA6h7OuYUwMVeXLaOe9Z
IPAef2YzzTX8CmOUZRYfhBJKOU54YpERx7sdEUo9GgLZ4hfzKDiCX/bp2O6Sz53aU+YyJYlR4IZK
OhjUu2UeDnc/KIQ2W62NspxTwoxZqCXdJI2uLqXhyibfWXxSr0zT621z0qHTqTLCes6N5BLsyp5U
x3ebWWLzZ/20J3V89uPDUu03ifM6NuUQsdom70ALQ1DCkxS/reodBOid42E23D4v1vm9nPNEkfn2
pvUedj75b0ckJUtpKmr4I3Dg/dgWvNOyVqu0JhrhteMy1sLiyuJDxwz7UUVNLauba5GuqmZhbLCJ
C7FAk5Shu95x4rnajDxj7b/KCiuN3G6a5Dvp7r/n6NfSPxfqPv/qJk5hj6AjAJrCmUlnko0c/3Yu
+IXcS6zKCqy3dOpYbPpcWtYOjSNsYRLgUePrUTDqWPuM1ONt/B0ZkcDR+fCoUeZGpmmUbwJIZuwn
v9uOsEe2ui/jvJUG+KDiwmTkqGwwkjdC3yaMTxmtoovt8vqolmtDr0I/k0fOCT4x/12oqR1++v+i
y1lQLa95Q2/IctMHgJO9e7rA/ljMjmI9o+9+0ITuCCdAPIAN/O2N3m9eYkg+ens4Rt8vhCdKpYEW
xxYeZ3aYKEQT6HaEfFCRBv2ljgwj3EvuA1cSdZYhOm19R6faFi6B0PE87rXK5KGrI74nZsHQRm7Z
hWp4k41BJv+GNhLV4jL43yEDKZDe4TOxWuwgFlGH5HowvtNptC2ACx51iR6cQhPCXdV85FfPZkN0
XFNnHRuQ66X8rHF/h9qPhDMwBSIMuG+I5r13h49M6sClC5Vi7nYlM8iMg3Y010i8lC+SJNWjcYGE
5GHGKI86cIruM0rZ4jONUBTDNyxSgVEFonmgzQFqHVJirqaGIhACYJQX5d7ZJqXFQGKrRpCCyUY/
RvRic3EfPR7sxMdvsJwy5y+HtkvQf80G5OBXt3gMmvW0gcd8vRhYNQwxmEOGZ6RuT2zKceKy+cW3
VoPJ1zlZZJI2ymbsz3mKBOM4IoSJTtoKuizGlk+3ses8mVh89JCxkoMPM0EdIUd/dMBKGnV+X2Sm
mPEBEYUa8QkVIol2r3JVKN++yvFjRCmY/C74SwD6mHZyI7ppYscbJSguoPqsaSeGszAHDjozq0xf
B6oqQ0fYaBTdPKV1jaNotYXugFf8Ixm4r5DHxMgxlPJ8jKfKVPq7oVf8hR09E6Zjw+HxvRyljTEm
QCRm0gWiI1k86fJhlYJX22RHqp1felhrAvWINJ3DXzPwO7+ne4ZbneQhVfoSOVD79LgapvuonDFv
OaS2ga662905We8o2zbrWv66dwf4howKooC8y1i//78f830/WpvAsymvCEr+TCyYWIq+NjDtEdui
sGBchI8y4X+SiAv/6gf2Fu9Y4p7y8SYFSglN4qJExwG7MrW71QKyJ3sAJpPDSPFjHSqtqy0NRXAh
WS5yEoJziG4qOj942H66ireY4dFbIuQvchTtOgw1Z1MhxH204QaZ4E5YeOwjOjWr9DmCBeL6Yxl7
Q0CMyzw+Oztd3lvVoiAtvWCbKO0I5v32IfHeoWLlueq599i3zs22q+7atLeBqnXXdXoJsto8uzGz
Xu7Kq++BP6yJH/5/ginpHcyPbLYQdgtgu7GQ+KSrXn4FKVkkNaekF1o0D14mexDLJqfWs+8EwlLO
44Yvi28cMK82yq22IhuKqrS3bGdPk2wsTPWQdHhbpZFboZOZO8geyj5yhyeF/eUcMU4/Dn5HttlA
DYqbgCeKAX6QGzeBhgRAxILRONDOQlwRbQlWENxeC2YEGuIAfDFqFMLP/jiLsWntrtf443gUXUSu
zwRIbE51C4kgycSh9KAC5B6HTGbILbkfj+kiejWgxDNqtcqA/4b9AnpHQFsD6fo/C4FNEdktJ2KV
HWLOSAEvRxnjkiv1HEnt4XoB8wmr9LIPxZ7tVSlglqpOyFpKg8aHYvsLorXET12J+DtQy84UcWc7
PHkoEW0ZGO1LqY5IKja5UeovDT97aGEe2nDy46LxLpidG/UcAhNwywGhqA+zdpgHItCmY7Svfp3f
hRXTbiAB5nRZItieRENZ9kiERDqi/ysKPC0qOIbZ4EG4IOt9+6rbvOiw/HO3PIdTlEnSRbmrA4RD
Oa30KWOaYmqPihAhLV9iEl5fkJkNnyBzJAxMGEcDJmSuZOyTwndMuN+EmWM9LChYjoPnYGZtOsRl
07NatGE2ZeH3Df/5S7vSBC8bq8FfhKLdeVx0nzr8XGnbnI3+j4CWQEnzP6wbotwFz//oFxIAuxBP
6oSH70Re56fP14QanFXHXGfnkhjDm2yfH3QYnD6vkw4uFNKsbMDtXPcHvAZ/khcMlJ9BILYD7V+4
H+A1f2bYAH7an2p1BwnqA38nZTzn86bUN9MVyLIjN4fl3OBlfupLLcNbo5ARF2FGnvVMXJAh77mp
HJPfQd+vWnmVGtxakM+7dxz+1VSQmU5I8g4uGUcyaGU6GB8KX9FL8eWRR+N6HHMEoFT/fd/H/hUu
urOjr0tCO70VeUADYRtkneMtYq1Qitag93nrRV0hutzpwB0pmeTVrn490J+v8MwHux7JqTJd2R3e
fjmxrZ9PXrhQH2k3ACdZHTyxpscyLk6uH9SCRJnFhfVTFYBlOq275kWmvTiAkcvYN/3pNjyNWKKw
vczAa0AzUZfy3bn86S8S16xneU+tfKPtNUSsrRBo4LFaTuaI0dw7cqV6MKyx8kK4phpvBwMc1EMg
6TKJITtDNzToiGLrgmN3/CKTo1h2NhvI9WYVRper86AOmvRD9RtBAR1mc2BWHWt97I9cl9MeGiSt
tUDcyXIvJlFQhYdglnmHSKZlMWr7C+LkeojTi1AFNoqU4N0bZJl+eKmwKbNsnrXvf5Mtsq7kXlux
6ssPhqw34+fZjzknbqgMdl09SzA1OqB/oE2v1nyVhDb4SG01YTRUdWZelYkr2YC1ELSwjRmH21HT
1Y2dPAOBK1ZNstZmYZujiDNsC3XjXS1jYVgXzXgKiWJ2pB236k5bRgW/aZ8KMYjNHSu7cVOTdJcx
GZtod+jXHBoY0mBAksua2OjlPjfzURPUYtQFcv4+uUmhPszJO7XDYMzJiaD59YHIA1DZ2XQS/JwP
MjEYAZXmaZAMBAHrRiBnnvJ29PQFdnH+pkcdS4hem7ib9+qIobh4ldTHSE+lHCzwQI4Vc+jsB7hr
8QsoSVOVXAzaWnWugaczZjAkAcI2tdLTXG+EROJzq3a9xAJeMEKlQenRQTBxjXJyvs0ega7Wucnr
aTRpyt+nGH7XGFO+JSQWqflogRzFGxgjLGiUgiwoBleQCOF9lcRBsN9zpAxmo7m5EZpKfv9csMqr
ce/sFmXkH6lTa8FM9S6xR6uF8Asf3TCYAupy+S6a4kuEp4VBACVvPdKiQkPR3stkERDtb34gqidt
LJ8d9f+rESyZ0xfn0LG7RSTGPL92xFEasdT85w9hoR4MmaPPmgBSTMkj93qBcGnDuqfswxrfWLYc
hIIDH6texKzty+zJbDz7SequIbSleRPIkzw1twA9QJqh8OnBI3B2tvuPiJ+Yhueo5r62o978Vs+D
PtO8QLUjSyD/5xeRdm+GhzIRnH4zllTZ4Lc1igfp8GIbPy3ai76x/5W0m0F10xRhMAeMZcTgWK4A
PFl8e2Z/TYiI6c9NoB3uCoAQSW2TmfGlA/Ox8szJ9HfkhEfCo8QACWooftrVNW3dTlUxoZfRbJIu
5OvdkRkJadZVAE+7PwLU0t13LolfFA7rVpbg4HPGpliSQcAMRY4eTKSXK+7lnGlkCAXw/af64GC7
JvUYCZdUN8EbF50QZpZ/CQSvu1kjXsMGvQAecRMulkPWTKL+aKQhoy8ILceddVAYnTgcUtwIIyof
fixO/s1LyIfbF2x0mqrZcXU4eyWRh9svZjqJL6+OHG77W7Fiu8/BlE/qGkvrhclkHnvXg502/OyL
Q4e4sinL0YvbwnzDs2TEV2MH+THv24IcSGMXljqEqex8zLj+IwkdFoUQ619WISiMtMTXxKrHSW+g
RlLnIcY+w5S1eezexfupJIV1HmmPhQV9Q9cNuohQLxTHFd9JWNpgiLoDGGQRiapqPTNDinB6hBBd
8YvZ+TGu2T6KbTXlCjxdLZIViVpkt1q6KJ//RHgujxScZeOxBNM/mT++S6xQzw7wBYVAt8y+tFwa
+B2ECmajSOMgVzhB+Ob8X+W9+oHyStUK1pE+CQiY4dRz8ycM7km6DlQ69hsGeYtpq8nZrkx24gsu
c8R5AuDMQwXeYIUrzqtc8+tyy6ojsizus/6/3KQSil96I97fX/tYNhZKG4o+ohhN6RoPzIj3o+e8
rh6AdotJWgwLFOp3qKZRDUnxTmo7vCqJVE4lBr5y+RPAMEhwLkZJei1k3mEBlGBN8olkyK/5jiLC
z+W8EkWG3h6XN3hVZDmwjl7sPCNpPDpM4M+bV4XQs1UFMTrU9AovsIiWk8seVJhnfyrHHHAP8LiC
iX1H9U5FymPo0jBbeY+AfL2OdsbY9NJenZdqB5P/Q83E3IvyURENIs5sOjNDb2rnRgPU5r3OVK6p
sPGXNP4yXb++yn2iWVpDPnAMVqHyIYQD7XGG0Dmnt2KYZ66Su5xKLewJWYmipnMUNaBuERE0nQ9L
lZ0pgeT/OpLYCOAwba8XeXfN9z3MheTnLeT5xlAI3ke+KM+cUPVx5zBlBR9wsmRUESjmP6ipslAg
NpGZosisW4Ja6rLyp3Y+uSi0gYQmphMja6vEIPwzZpxQPqLnW+ViuB5/oaKxssXYSdFwKHTHNJzo
NT/+JKxEbnoBGMzbC2Mb0MgrtsXi9ujPWV3f0h1GoQvJ+wMlLizkGmGD/+WeJgdxeIKJLN4Q/fPR
xleikuV7EgZfpDj7AOLGZrN9g+Bvjnc2ow1wYSDghkZhNGEqyiDB5+nLGx0kTgjp4BkkHxCEEFhu
Sq8UdCwt7R2PFNNJnoWgWaw1jx5gOzKCCYIwBu8c+0p+gD8zXe7C3LXUZ5WEJhNiBS1b9ZTQFWjG
KwfHN/dvO4otDDOTYkM290YxI+KrsuUSajIvk1GmEpzyEuzMjHfTU2spS4eoihJke25WGZnjhzNH
qf+sUJM2iLppZw7UKShpIon0ik8AmV90Ly3GDR4rlVEYIIW8Ks6JXzbJ/+k4wtmtsWkW80UVp4hd
kkxRjY8NgHP4VNMHBTJmEA0dVnahYI2cLCoOyHT9BFDZu1GhLYvkk3j0u2sCI8icEVmga9dXrycf
j87sw9JbmkP+9lzEqbHTLfLymxUxvHlSm9Cy/P/v7Md/e8leiqDRGNxA+BVfpELz/A+LRw0AkEJk
Sfevg5fJb89NR/pKwIVUMpY+wylo+Am5foYt0GNuKeZhTUMm6NIbpPZOCVg/PZ2B4F6kSSlROj2J
W8RRkQjFLaOBjqwzQhkem2jFI8xM6luQODxHAeOCQJOs6SguMtVv3BGKlFLpI6GszjnKwRL3UV7r
iICuf+6sIHlF2BPOlZmrfm7XZU5ZS3Q14xaEdwtTnuJ/cX3LMnYxaanE+dXF1WHThRvq2yo52tXH
8cFLDS6AsjBX/q0PMcBRsANzo0z1OedzBV72rT3GVYBAUlWuBoRP2/bYqtilVJ9r1W5WMCTOR24J
N0eDyZ+7m/bJMbgAPkCNX/Mvn7TpHCM20oSJT6Pn2CvJfiCd9Q2X0dmsyBBQIL9WMo2F0ckRoaAP
ToMsdEAYMlavK05i51qpf2ar49Megqcbir7NDLY+oZIiGSdm58QzuUrJpAFSROdlMKFHIKfrBFNY
DGplKLegQGGGHoVkfy1BRwckxbhUVYK+c10ms44LNL0ctcA3qT5F5a8d4TbdhEwVoY0i7rT190ga
8ce3XhFoQkUU5YNVfeBW0yoxK5vWKYQNdqhG2SFIv46oP+krU2fxaPBcEytAhTcyfArtPJLj6MVW
ow1oOj9e32EeKgr2+BhNWwVVsuIUqf/D/SqvkvDezq8mPVTrOBT1XbI+SoXvTiwY68GQ4qvqXVDt
PLyX8nbsmD+oVMB9LKzDZMqvN9TkHLVmUfNwhvmhqAHPmoPVMhuzphy1aADoHUu/UOe1L4H22N1K
000rFRnPwxKx3QVGC4117LlWdd2cRQIjeEvgNMxw8E8ig12q3HwCeLb9zV811IhIHafLRV6osJ7r
GhWvcOD7c5D6Lk87/qfQM8zBPDTMOpy6Eg0uxtwBn7Gb8P6KpieDcVnbwiGsEMXJFT9aVTUEGEPa
AcCXgqYk6uX/FwMfSCEMrpF5OFVwKxiX+D08lW/EXpF+O4rgc8OwM5Etmp4YHXkcyy7Fp8+/jInG
EfcRHCirzgur0Dl1uZq9sWdxDBOgqBGzhOZ3+g6spUVxz3TjnKlNY5hX1eIA9s3NdnDOlU+bKDon
LeLYRtdry38p0QYBMyxp+frTUweeQpnc8TbUBgEVoCXxpux/eeWPnxb7B8KjATXKVwr4qVUAQS5L
mBL5GwNdk68YYb8nrs1lZgEVwJXEbIPGyg9dxeVJJclHFIhAyvWCPdtwia/gh1+HvppIVmm0DeY+
Z954v6zX5zmoqI+YDU6u4hofjG+bMJHTTllZAQ7BMo87uhMvqVlQLynWg6u7h+rGy1slWhprfoCp
HtePls4viP3KIQ5Gyi8QzEXLt6R7tOLjj2w5Z12NaX+8wuvaZror4z5TDSIzWNUat5PmedE5tQeE
4UXLcEB7lMbw20GdoVQOA5dK/5YkJWLzYeEkfjshh/IV6jClaiuUUJ8LM4ZLz05WKon+QzjmaBW4
QjaX33L21qQny/X6Hmt8ha+++TcAioW0Fg2rIQwIF5ayzfnNNAHuHpJodEDkcRObgGHbFMPy8+qf
6cia3Un8YcpNKPAeVphpY9s6juK1TNfNUdYDclApfrftoWoiaV5t3q4Ilgt3f1AzosVtfDlgf6Ww
wy6u3Bki/RA+X6WDETtmOclNREI4RjKupDcpW7iYeeK027S/7PsZHu5PN1TFgS7L34ubtA09sdqT
VtMPOwWuQvzgC0VoSgLmHW2quT4uKxFuwL/hdZ/wl8uatnamUCnjx8KVirmIw6/nSrBRQHSan5iR
fk8z/m+brpEbY8PwGkAnaVCu9TdftU7Dcb1RCg8xxEOBjnaUA1vmvbw5lsZc0Ij0JkxqZd4+aGZS
/VcMoiN7yOODQkTk88ogj5liU+x0qLnHH3zn1Z+PmNJAoLbYuDhVgoIPUZDIgsdn68CI58eWEH8L
KEPrYtSDDwvaIKue10BQYRp+uAToAV1gYSSgGt/QIakZtr3LPZ+TevV7uWVzZUTPERPSAvESOiXp
cfqxEJP0kMY4NLLKNdPrEsSlgSIWf6ife2VBWyiPtJ34/aDDnaP2V/GfXUE4Bj06Ixhag+d/RBml
UdX8VrJfW09lb1k4ab7lRkU1vUPO3ojdXsI1csruwu7YthXn5x4aiXC6J2QcrFQVDg8LHrhWwA7S
o/1AkinEqiX00f9VHjg6rBeeg9ZoWFYRO5WJ8qq+Scxe/tEFFcpHNBpbhEDmWirfIzSEG+kuHBia
l3amS9mJvKPar7OVoNtrM097z1L9E3mZHBHi+SKD0vyxKRo4X430dX4+sZryWNF35h9lvyWMHaTv
SgTLmcLfnT5hoLRtrx/CdHpNOub9te9AaR8Zr62tVD+6WCK9wT+zwrtTWJrVbLT3lb7ocwQ/eTbo
qrGLi/W3R/2D6DKxibbb6XEIdcc3HQocAd4mp7aTqlP8Ga5WP2yhFG3rC73kgfdKe4YwB+9WR9Mm
A42PXxi6Hmlbdwdhq5+P1assH3+Y30gb+VeI/x3ICHyIoYHjb23oiJib8LLqOdDT1HKnPGeI+LhL
fcVERk0375nBj+aA0AYaq6Nsb+pqHP7CSjQtXgln2/9pqnJKJERb+jI4oBMQmYF0vEog9+EGgRvE
lBX9Tc11/MVVkW/f2Prl6cY+tZXUPTjrzthMwHlJ8SNM0b4E8KkSEJEKJUOgGpaAZURuuyjTC2GN
FM/jtrqrBcFQwGQzEAeOrH3ef/Uc/FHVo9eJ7pj4LRV8AIwlDl8XQzEeDQagzHpmhuNVwQGcuB0O
lQxGJYr8eGXhiEhW4n5D5MnjrfUcF1YngEc8g8Lz4vq2gOgRo8xXorGMxX4CJm0MBjE2JZWh2rTw
3YcZeMrjoGamp7ckT12zs4OqjwEo5TN9F3uNVsfKamKjxEN8uzZnqmTUL/DTOZ3N8RdbARR3DjWP
OgPEekfuM244blXrMuv0LzSr0jMaDx83DuhULHq7h4etoPuS6t7Kw1bwF7aQJfHUzRJWBrYjHFK2
JLiosDi4yxY2JCcf0ear3QkGkuCsMKwpEHc1Q8NvRrGt5MGxrxlrcU3PceQqCzYPRM9npQ9zPS9D
j81gcVEpAL98h6QyPTyxiMD0We+5VWlwiDUqZJuBmOdEpzS1dC+MrVx8/JkRr61OPKqg0zo1HPpz
E7mArJ8ZWOhy5kKQ6uK3JbxoeFAi+9ohIGL6ZT9Yf3q1fyS+uMnqFN/X2sgP7aJRL0Y1Cfv4jHGV
OVCCh2CvegC/tlSWqt6Hk7ZVrbkslo6CJkrqb7gl0j5bLvKc0+H8W6vGcLNKWBLu9HIyYI50ye//
C3FT+EA4TqwfeG8hb/ip+AnXMlNz3TD+1PMIAb5oWdIN5TVUzkgcQyde3ocgTxAGzCqgLM6Jezdj
ULnq/2dD7/MjlF8hIBbf9J0PBGADhSSOsZZdT0af7RU9SOFdVHQ4g+jv+nV7sVOUx7pge+NM4XrH
wsP8qHRWAGswjv5aWidDaibX8jUSzujhUqt7Y4r4Rp7TRoCODJMVLgMRBORXCH1HZiu3ira0/pSI
7VVHu0cGR10Vq2ycqF3j0bk2OcsH0mK8UKFa2FPfFDHr5peRGzX2xUCr6fDmXR5vUIQu754QQAiO
togHImLs89H8XwNBzHO+6jr0kdC2on8xLWj5HFoMvdsBLK7wpuVNppbvFc5Y5dlKTTZO2xIObUOt
2BasinGUJxvq3MF87+bbY2wiTWvDYZnEOcJ7HCgkn24PcK9DjkQLRKsH3TneV8ixfftCX9l65GNg
xd/O5RNRe8mqiJlVrDv2sxO3a/RuGIOD9TSKsG09860efpihBtxZEkRKQvIO5NFSjptwbOvyChnL
whSUT/0mG92uIPZ9eB8RZassbBqIZP4xC+IzmEnCzqVIa7odEMPvlMtyWLSkHJELjgR7RpYqTdOr
u4r4SMkYJpLi0RTbya5aeaOcQoEozUDIR+djRpHGtgp+VHVPICRtqeRrqtyBswcJU7d4bZWwwmDk
GFob9iGrRcQNNa76guagT82Swg6KEfAP7t7lZIY9w8bofn0PHQc+3d/IBW8vqT4oihTGgx0ob7s0
Po9haXTEoNo5lJMGg2dWaSMxW4kLF4pAbNEXmRBtDG25WZqu3BJizt7oXkkNHSPxyMcBKezCi8wX
XMoyjz/7CZgCjcnbLeQwMdL88iIRR5SI9X/nZCJp7m2Wdfu7Rx4orQpwD6HlG7CKAWS/PzmIZc7M
g47Yiy4im8SSupbJCww6EaXUCV8+mILxAP0mg+z8VbSRyvAflAVkValrrOy3+LsD0UBD9m05po2r
4jLS7LGHnLAG7Jtv7FFTvXsYhZAk8WzcpD8zA41oqgl9h6lLoAOOig6mPqymS0BwqrSFn3W2JxOP
rwDXztJseH251J9715LFvC/cW01zxGS+PjhuGIcCyumZtornz8Z+0+09UVp1+MmiK3BbWBD8Q3eP
j/GHzSg9BPlj07wNMd3zvQ8ZzYcZc6wHT6JjessQQGAgIOoDTRZlmzAvJevxTafhItzh+RdqUNAD
RcrXlDBjABm83e46haysVIVpI1mydMlXqmff8UitRhVSh/17BElsXGiEOzpYN2v8FdQyR4kVeGZ5
Dt+0vmGm/ebJLrs+5vgssxsmIYWWC0nziKKTPyy4m25QfoHxw/CRVje7QyG1FpXWMPHKLYuUxp+w
WcRKTWItB7ld2psdq4y2G+4Ps1yb/ArktzE8rp9zXtHWx+QOwdXx3hhTDdRcXpWKnmtlcp3T6PAW
7SV2oVjeO7wmpW+JVqr9ImeZuN+KSR5mb5DfPTaPGX9uKw6mgXRTs3tWBp2QExJk008r1dL0rpp9
Z7NamHhp9koa5a542HswbiDqM4/gNFRrQherXncvl32iUGZ6xtpFLEAUI3j2JrtpBwbx5Ub6U90U
sL989peAbH6DkT93MuUqZ+h7brTYdw0MX4RaOQB+93ViYiPWbP90a9Pid/Sj6fUYiTQuMtsWiABp
wQSxFcSa64kHe1KYRKP62TngKgMvZY5txfppil6ujhO269+MFQOmq1OWdmZykejReg5piJVGWI7F
OX+fd8nChg0Q2Q1iWpLl+naDCn9u08EGDGHTZsi3NndS2mus81pm9cTylJgtgBRSRdGCjt6tnz9q
dbJige4PRo+M5kSvnWw9PRizvBIPAdm8EW8fuDnBujUzPyNIjN5iz5dFGvEhwszblM4TGaAKT5P5
A2MjN7+amQ0NOcN8dudNVZzdN4V21WwbfnhBw+4cb1p1pZTLvFPWgwx9IrMLMLDmRVEueCkc9kOs
a4vr5miMla0kZaoKKT6JVrLyuiAuk7Wo/rJU3j8F74Zh66rLFmk+yQb89SlDDascua4w7BbwNG4w
lnsrqKXpO4EUo/Vsjq7ZgLlWBQ1JD9kWetwS7qThpFgUB6G7S8jj9SN4zmntkM/p4oII7N2xY8NT
gCuYU1Bhmsu5rMxhwvYQBdl2QKTYqwzEDCdlE2UEFLM6M8oR2nBeCcuqVXDfAi6uP6/cWz2/3730
Bw3xknHk88y1Fpcm3SBnxY5HuXqCVHFwONkJMnz5Ip4mWWecWPNti/dzu274+ssWQ7VC89heG/Ek
t24n8l3siClFQLIqpH+DdjSvH22y5+T1CF7VC1T4xneQYYohPfYsNJ11xenbfscHDyiRw58TvHhH
kWCTF38vOwXK5hFHXDfjzq3HmoxqNn94flalP83H/J2gY0toAM+n3MkKRZalOe9uCEUCZSyDX/Yz
ZxnO6Y/RQ2PszYTphiGqC7hr4sAdQ72hqIj0wpINCrDpTNhQ93xHXshI6OyS0uO1eS4R/JzePTsB
xFLxN8gRQ4sh2vx5MXpfg3/xcm0KzcqrVhtiQraWJDfv1c6MFfrpA5Rm96WsFyp6506xxNe6NVw7
ycijbp7BcCP5nkluCt5ZeCSliSXfcUpaV/llOwDw0Ofoo5C46gIsFsff4GOev9XIBIUkrpuUpZbU
X8YeY3qLwbUCOvYcBKZ0i0ZBn8YdFBgeejlfY46h3vkdguxJ3EuXOtejDg+F1LaWFOVThAQfjP8T
sg+BTxTy/uwai73fJx4tQETqaMxaPnE3wVnoFy+icZgBV+Va2tqxoIwyM3sokseRL2IXkZOgoYbd
EHXMJENO9+3VbT/4MXP6mr5mOKNHMR8A8PWU/tbxbdxWIjEXUNHqD4FWPBk6w6zpt0l3YkaRJvgp
ysw6uQESVwGjxntytbYV3u1u55yqBachZ0FQ4rxNr0zbaV+L/KNvOJOZS7Mj/K5EcvHlGxUo27l/
/jVc3hG9zyj3YKqYScyfKrvq7UUOvfsC3J/kfNNjjiYXGZDiZ4f+IX/fvtQyI01mbG6cIeMIKJF8
ucEPZLDo6Stkm61Ya4CqTeAF3lWgTa6dmnzD2jlhcjVEdrsaFdSmgsK0ebGIY0WZWtN6TBe7UUwd
XCL3voLoimds3O1JoRcO8cR9X5bHknP82XgxzRA+fqOwTxqu9VCk1d6CM9MigpOF0XE9ZSewU9MV
ZxXdcrbrDTrdaHjAO0KJoVaCB4rl7m7Ao8i2dfiLVkDqqSZ2+IySDCKS85JVP46jB6oazULNnCdH
2Yjp8lhj49L8goD1Wg3+rmMRX2w49Ya5i9dqZgWwB8HFdMdk4nA2Tptql1VMaXsOyuAIiCgYfbnf
lfwAJWMVU0XtPoD/WsAySxUGJwvQAKXyXQ7CA6N9C4g5ZnPamUtYqi6BkydIWuqasv3dv2D7WTVA
BZyOyEy1nRTdxQb7DaRzMC5TXozB4quPKtkLIP/Wr6d+/bz2OWJQUA3RLziwwL7Rr6CxYLj+AabL
tGLlbrajimedXkDVII4vdvYFAnYo4DMKECGKZDa1HEruP4e47omlm/aqRzk9Zz5du6F+XqC+P90X
ucdzJ6+0J76bRBN9lMMvkyjseRI4AD8ZErnSau9vpIrVb8o5b1u6okS9/EbBk9sT5xYudI9hNp9K
lFlWsgt32bghRmwS6ZsEoKsl/Qn/OzHuJeckEbJzXtqbl5KC5DnoSuUdNXzlNrFpHZ6sZV3XuxMB
BkMb/BK9lcG5dWWOeiObJMgqWldcDB9bD0y/OWFkl8q56boa9/BBFoyOF87gYQpMVe3k6uMPsxX8
b9vUfqZPGp7uvufPiuPp8eRl47A5+LAnrwgXWHHwqU/+OqvInGjHHp1lYG/QCFJRo9OmmYoB4aM6
0rHJsOIWELBOAvCOclCZS/XBt0KMEziOFZKJDvK7WdTjLdFHYtpgisHopJkS8Q+xiDYDHBKPZWjT
YHhf5YOAnmKnse0XCKAv43JqNDwCSFhukuWfCuGsgwDkSP9kz0tIU2J75fTalADpTDl08r1tINmf
4xIrjqHa5G9wNUgvWDcng0hHeHx8otKEE9A0JmUg61loc7snBtBS3O5iuzJKZN8hRA/4Mw08jJkT
cxR+95Zi2nby9timcgsLUzkulO1Hle1Je82ov2ave/27yBunKN2BXz+/b/Py4hn3dNHsaIGHUaO9
4dPXzgnx1mIC/5ZwDY3KtpA3rUyFcsRxgBPDQF1DBsgsMIZfh9hqzRJim3F1OEu4dJWHYIYdgsjP
+nWGuKReZ8cxq46yH75PLwUFDXcCrRQh6zmmRVBhTSti0VUu9R/TFYYTjf1HklI675KLtHKfU7pb
o2jsJtV3iJFA54lUMZe2gVaR8fLYqvpsNFpGh4JRUwpwdcq/AEyyoweUccQgm0fNvbjIB6BkY4za
o/MafIe7i2hfgRggdEUoWFkLyRk/oowVMQyFcQ/heVezqEkiD78j0deFz+UEgQXI8c8zQR2yA957
4jarCqe2Q36/0k5mfZcOSVEi/UC2x703jj87T+jtPcmnxm8mhbJJhvcpFBWlEFRA4wpP4wySK3z0
3GvgXrHP2RwA6m7vkTINF5/XOFkc6KxI3eignYBMK0OHUF6NnZtgc9WmzZxTzKEeanYKmOTG563V
9krpQoHHSORUMTbtK1c3XDH6hwxRHH9I1TwEBNO6DGdNYqYfDdXcy2WSco4g02zhnK+OGOvna+6p
g8dwjj1PVlclD3sqge+YwTEzgLQnT13kNLE3/N/sVG1LQvRLgXIBN+Ts8cJLo+4Rk65C/Ye5BkgJ
tR2h9ki3TdaB5c70e982uFXwoRc7xpbYuFmr/jtueGwBENrc37rMSYSY5o6bzNICTRtubDJTgapb
MHgFhOZTYzkzfl4sZstQzAuuTh1tZMzlDmV3gQ6+0aLu/bEX5qxDSmIXNwUFzEbvRRh3BDyobw9n
mYwNkyiBf9VR2s1L2IwIbtLC9JEuoMGh/yQVgRd/0vhkCiTUujLr0hW1ToSOLOgUT5/qfu9cUJWK
VHfNVsJtsUDBFiZMk8D7FA9LNbHX/ex/D3D/1RpeW1hNoP3IuQaYrUYOtXY0zbXxBsN6Lq0xCwko
otSjgxGVB9BVDBsmAzTjtczU/dmou3yarWVBbggWgd5ji8udPOfXkiNjC12s0QhrxJv5Xj/Bu+nr
QmOGbP++IUv4UfNhBITFYSyLfaphz8x80gruKAnlXlFf4mzmtccFTGpQsm9OkXhHErwTXq2zbQkg
/1SrzRG176T7ZPJmoPF5R4VrkKfuZpwdS00Pn76WLWQY2Y2WI875YhlI6gompmbgXWlJs50XbL/y
1NqxZHCKFqFx5KJcBxn+8vYBPVemT3vbr80KaqZbCaAPmj/oTfeLPXNQNMOhjRUeZiJZEO8cxm+0
F68nkt49iVqSva1WMvJBJHyE+E71AEvC9htwx9ztd8ATfqp31gtwt7eQNUgtAIkdki/VNQctv+Th
yJUrMK01LeSzSFYCDlgTjI3J5OBPPANErQllWSVEQONsbNIQvR5au+cR6kpamKN/xQ5a9ae0J02r
VLFnMt60uPXYKQvrPT+cIqLg2JTVUOP07TAjIosZ+R4YFhxp6kJm9iMTWEHqtIo9DUmUDSnwO9gi
vy1E7xuHXzb24J1eyesyFplIc5qnFFosXQXOaCxmQ5MNp9Sh1Fsblw180iCGuw7RPFNdKT04IabY
uqottUE3pu4vlOMiPIPfPHgGiq2my57pfKaSFJ4TG7JO1cgS3VTzajF73yGJ20GduDu3yQEJIHZx
MZugYFNa1yagC20vSgyq1nCYx3XtH4PY2KX1wQBo860LF8z6cKnUY05uUN8O552ulBuF1n9krKN+
BmULvZQvWW6r9Vc9Lo3YeLwvl1Vayioxdy8myC2hqM4IKZNlsw+F92+lDL74G1aJmaNIa0i2PxFq
qQggdCqjp/aSyfIAHzMbHnpGhNeMsPI/VAVLpENLOnmuoy5egaqkKVUB4stqU+lSlPVPdZh5g/oX
qkTuYRh9xBsmD/rWGZA3CQumVO6rGPaVuxycCgx8wAmYQh3zEXF6yZESkkzITZNqVuevyH9FLanN
S2c+PySTLSHrLl7emrFOfW9rCA+YFcewg9pZzr/AA5hnhtwd1DoJ1WtRj6ut/3LjqSBLN6TLdMdr
8O80t7gduVPn6O8a8dUFeaae8OA2YgIOULHpkXkXTrDuvXRv8mXAnUaZPN+mysYuNlDYoUQGrnur
sSfHo00UxafR0lR+fAj2OcX0V2WXt53CA5tcwfV5Yld37y2ssQbyRc6jX0045wiDHYYJvw91yMXT
s/NsOR7sLaUNp9OYPhei6OHJ78kF+l5dI52kwhuAh2bN+2JrmKfdgI4xE+hWRoje4lnHcB2CwRUp
f+bp8rFZ+g2QduX07kXxNDwobzS3zUijsUWRb8ZWFn9vYWHTExjm+RJ6ZuqsFwcNhdQ9SJi24c03
daUn1iOzGDWD/zK4Z5HZtmjVkVlMlNGCxRrcW6MxMdHCKTCrvxK0bBFNFGKBXN0Pvhne4s3gnqXh
0qNRJIpV+01AOxv7EopPvmDM0Deg127IuQR11swZe+BkGY2mkBamvLrn22ejtP20Zso06dj4DhGr
IaIs3i6owkYXVzmVoW5WPv+fWmOli/hoyh/OfCXY040fVCdXectj+PFmTyA9RVU8U0SwGwvMBta1
d+V/e5p03QI7yvjKctpjDE6IxX76OpYUrbDxXX+YlgTtpCiNk3bYqTAlt8NpWGwnkXY8G3HXencC
LSW1GPD3GHOjCgLpkNOaAhKwRy2WEh028PPkjgHfLcZzID+4Q2JSdjYvbdmsHZu7XQ9VgAwV0k7Z
bZQp+vKZgX3F40LEPiFBWBVfI1dD8H8Sp5gaz0eFQ/07XKp3s3swaTspU3BMT37gmrqWAb5JPH0D
n8QjZS/1p42VMcq/nM9L5QiXL5XnL522MyktdiiM+ik83AaIOhHGD/scGq1zmS0C1HSgM/N9zLRJ
CWFor8rFqyYgLK/tNcB0EETTw4ENbqv2QICx/jOcD12PfJuJogZXAvgI+KdyAy1P9Zt9Sx371a54
fq4csK9MIZHLt4bjHKz1vciqVxorKFrx+8VE9lOT8KimzEJ9CGgtAyyEFpST3tRHWH9DKo2gUYLs
V8eElVW7Qlmxnh30lSQ9V488wcvGbHklUcMG+QiJPY7pbc1GrYWPEZ2XUVKdys8Qio/WFyDroBK+
91ZHlnDQlKt/OTNuSKlrcgqp1FeUOX7gbES0OyhBoNLmTvJqxUs2PHWJFybSPlca9E36h3F5kJt1
23Ppiu6MEY9Z2b/9l9ZqpvBMaGVs3xe9bAwIFPlU3oogXLz3JM2DOXVMLip6TmweSe5/Jc1pzOaZ
k6kptS/qU2IQ+pUVWtkh1aHxSzT8x9kzHlzpkCeNkIt9/fgZvFHKRHDcVwCVBoYwoVSGKPeU8LU8
SZ/9e5qmyqXldDe6VwLFbxR5BwxZ6c6E29UuDOBHhPkTG216UpkK3rBV6/Pe3m+Z7ErJoL94uzXT
7o++KMzGHVmQOE45VuApjBeD20N61A/b1WAQ0ALRH21Gab8eVXZeh1EKYg6OUCbgn/XxQNddFoL/
lzVIsd/1uG+SX30mMjguZk3lJuXiPkYOxtsvw38Hsjgfqru8K8Q2ONdbAVUtlRpsdb+wIEwfDLJj
hi5KCGfnfzzYwN03KpDfu6JQt9Ivi9CSEH77qWdD019RpsKFjDij6EPZ8eHJSQMbfiHc2eu5cIFz
SejLjeLIEv1swpV2EqGe/5Al9Q3CW2u3mttu3+dSSi86fNlsBabFKf32c2ifMJubAXjlb1K26TYs
Le4OWh8WgBFfChnNdhmmpO7PQ+LPDz288BRGxm/vltv0ILQSRU8uGR6wnfIgsUpfXV2UUeAzkskL
Pwn6883He6NreAd7S5iZCx9YqM+48hpi2D20ROIvzE0U9qwSWUq0mTBujMTNI6jNBgaZYWl62KmH
mMRF95kb6K5k8a8M7zudDXnErJAhMhzZsS1I/JIiAr2BnN55X/Ynz6kxpIs19jQOFULFUdGYaYGx
QkPnErgTNDgyLtN6yvM+lGh+cCqf7KARt3Fpb4IxQDkopnlYoRXmod7eBeVEw4Tgydve4FZpjkEn
WIByoGP8ps1XvUdDQ3VuYJPSFtXh//eWpSalgcjghyvra6Yz3Q7KR5IGiPG+GAdHz23hYQzIMgyr
aDgiHZuwwCxDC0ALkngDWWckDFXJrKJCQ5q55EATmD73Z+kj+/943yq7/khr+C2ZJ4UFA2e3tFKT
Pyasm9KTNuBiYgFNcTcM9dA+EbPnKMP1wRW+tQ1XnZ/cnosD1TG3FZyNYUQ1dev6nxu4sGOVXzie
lw6GqdM7XbUuli8QEDBMMgUSjVnkgi49AFUVlKykjPavF4AS1hSB6+1a/cCJWq98k/w228d1ZHez
EcdgYjlMGBzjiBQo/rqm5EgKXUXGtrWnOUCUbEPu7l7GfS4y12m+Tuq888wWawSvFfaNt2527bcr
gZQyko8YmgIMgRR7QzSAmewldLt82fG1VNjjkCNVRjFkuBnFTptvuLPRW7kbRKsyGlNJwZkJMi2q
WTa1eQEWRe41S743RJDHdPZnihGZxzK7EzdiVmznfF025uVKDLvgh4tgo+8r1W35idKw2lXk2/5C
UKFR1woys6/K+21QwUZdoUxNuVlpjqJPFiXQviPsr/rhHsxa4duCfUN2ov7E96IrUJUwc9MnkNek
Bjksbn0K6Va4c2mV3GFYMC2wCADL1/v9w6nYoVyU9521FUZpZwyx82bF1z9ZJoruEGwan1ZKsmrQ
mbGrm0bgXdgZd1caEj/aGsWI8r5nOxEo0YKmLBcJ+LaGQcpDMJw7w8B4j0f46G6oMlT64qU9q2cG
eXBYqF7E6PKV6s/5YH0bnXm1Sy9awOOkDpiJRp0WDtc8wpTYSUlKacaV59HoJCjdLH0l2iIkpKdg
/+Mb2k29fzGOQMEj1CCTKimcurlTcVamcZzpJ6pdcDd+oQHuS/6AFqzzp6ZQL4oQprdZehqbj9wm
SptoPT8KH4ixOpdljCo2EZmzQrufIaUp/QkL1ZMJ1wIFnNCDtIjn28/3gVVF11fIvzpmj74fARc2
EburlGJwlXHNM1aGQB/BtU7oabhyj/QWtwXLZSbRvIWZSO1nXMwi4yp7AQFsp/UAt+YIzIAwKUpL
YjZxyABKahMIC1SUY1nMV1aP9bCmHV2ZEvfvXqYodntEPb+qBxuHQJYpNfvR6fODeM8nOPmrc0o2
+dkrs2Weh5/mpfHZYYDhJ1kiWSTh0jFaDeYeBiolZABJNib/2JifvbY3+GAWwTh2yIJ9w54fpoD2
0ceyVCRNN3SeFY6Aq+UX2sHjRII7bwi3ltqsJiBkHQMk8iEP7XAo0/Rh1UNkBwaVuD7QBls37JAx
8Tc0Dv8nABCrw+HMATETnmKun5ZybplEGjb/PefD5mTqSNKbHgr0bl7R4Ey0dDlP/iErh79PeWy1
B5oMIiCmYse69ucGYJeLgBlG8uDcQG8Bsj/DBgQahKrqe0OiqS9nbnQUtW51b4wz6iEVYzUPkXZu
ffF6dsqESDKumUZT8Ntsb8sW9Rn1szHkNFmrqccf27eaapy0tdHpAtDp9FbeYdBcEyUYTqbSdl2Z
xODVutPCUkgzu79GpvFj9v6r1vXlEPBONUZ+TgWcuLCRnsLBICVqhBVU3EQjVdFtP89mjWrfc9Vt
0K8OtsU0uN/peqKtl7RU5MaaCoDjPvh+cv0w+eez+PxFM5bwYFEkdYWamd0FdKbv8bjmItgav5cC
HWzRUYGHiJ2Pyvwpj4YxSSqiI6ltbTGYdOdo0RLqDIcfeZvRvQxi7wHsy4tEzwEKXqbU7wYG4lrB
sEQUTUpWgayNY3vCDjFf6nVSGepuJkFSNc634xkcj+MhPLJ3zWIPbYy1mWC07gEYAe0XPR47Hjph
gFWVLynNUkjuMbEcgjpKEHq4LIcUcPs+L4iVrDi4QCgH2WXqRmkl/PedFJTsi9UijCkJ1S4Pqf8x
76LGBHLae0aMslscpzcwGsPKBkRipzMF3yFvoZBbbPSHL8XWwF791l9ukHzUyY6mZSjUnihcGtK5
uD4J/MlVxBN8mxqidSMtU5hJqWT81siPt7DzKWdQSH9Xo/XVylk/X4/N+czZ5vQADTywtxMNI3pM
j4yf5kLQCC3Bu2T7OfcY3vDaQiE4zuyTbJZmeNUQvv3yXOr66CZPLkLqdjAUFpJBF3IKFjV/KyyC
jEB7zkBYDv3xwVxHDMo97YRDiQtBr5W18x6RSJL78rUMAoQqv6o1PK4ACBITL9V1AnpXICxCh8Pb
ScIlnt3EowUnpE02fjNNRSBSDePqw4C4pz6OQbrUaBFh5/1NU2yZ3xcaQ75TFdpbZvacGHa1lYvS
26USOf/hdfEMiOqwiwVG0l45MVSpcWYsQnprLC7MFotS4ZMw+1muttWdepMBz0hfugf1BJ5k4IAs
pd6l8BbCdwjZaSOjPrfDPnznz9fuYAx6vqovyMWXub17XFq9u8Q6NIGQMP1QFkB6F4IYGQjO98wG
J2vJdZ3s0uhqm2usE/PcQ6Kuw3qQQqGsofsEeJH0dni4wv54ddJjaRIeCULnY+dsw8iCZi3bv49+
qaabAzN4Vzldat2E+aT7h7s5V862kmHvNogRYzSAVjxXEUT9BU1NMo/NLM12lWgu28iAmv+wjasr
sDcRh/A3hTy51TzTPiUEUQOLQWQH/AD9YjqZP5x+QPMD55We/3X8sURTsKNOsZpJ6jlqJWaUvaZO
rIpWPD7s6de1LoH8ZgvTOwBWgmh8PxmvnflxF/YMkUMuzNqcl2TBZ30ZjEtbUZJVyJQ+grqdKO+y
87bWf43pk4X+5dBbQmygfD276LGkoQMK4qec/qI8TSQeb5AjsNDDHNqi/Y7s37xCggA0fgpcZsLO
vy3NqAbYOQAPtGdOw+aLXPKVMqkK3MlyjwCUot1BZrxp24vwNRmJuTCOSjj4Xp2NRCVSsLI6bWLy
sZWYS9Dj8NGxnlJ0oV/gEHvTqxA6+zqZQkvXBLZd9E4Mue3zJzAGI5glhuglad0u/uARiVTRdj7a
D4dTp8xcCrXKd9TZxPWWb8UIdzT/RO4mbkkxHSsxS8rL9yoCi+3ON/QaLshhFW5LYkHKQHQLjxJR
2uWoztjavE4ubfpMlXJsmoXpqzMxCbQBZGkBjTmxXeYupUSmt1deJ7AiBFeQYUhhpRYDdx2eSJyT
cQO3zZ8Km9e1zXwapJBFs4V/Pha3R9o5qiJhjZ28HNHfYA6dztW0xTw5uedOSsVPLkRbD+9KNWpC
lUsBrHEpzLPkgFclA3HQOMn/vTENjRpfIWcOruLwJRlOn4Zdw6P+ojTZwJvcZjln/Epr0CTCxi9D
TIZ5zWu9RfuT4Pkb+8tYFL4XyIQ0fgtd6MlQC/t/5PBdHj5+N0HUtZ+hKfAvrw1cLLhOATN2zMCN
LDWuyHFnDtLthwt6osiu5vsUY6lwZqCM8nXOo2pYR2hiaeNYNwxxnzKuciA/E02u8v26RBiqIENF
wrl4cgTxe/UxKHwlFdrGiwmb1mu0+3WNOb29bV8JF3q6Qo+Do8g2nUdTJTTXpsbgk9KcuA08kUDh
0opi2W0W6JX0IEehxSHFhBFtXWak4HgDeY73Nh5HC156UiUDgCwFlNMflpzwPTvBIxMe47YilRHV
4rDXRzoAsd3TVp/Fp7MamqfNir6I+So9T8lmU50rGZ3IFyeFlPQ0I2+RkIkNwaNi+0RaUazLjPbw
NqEWnZav6C17WSLyIXQbHaMjap/PnWhz7RGIGHoMnQnBq8enhGQduiMy6/sNGnFl+XfiCwyCrR5H
0t4nQJJf8wsOjlR5uO4jVUkZ1uaYXAkv+xwgALFAmZOw9WOEo5FxECxdOtpkNieE/BCSZui8+sYg
RERq0lzwcTKaLRQ7uCEx4iHDvP3cS8SL/GKdVkxA+VVPz/hwtf+p7MXsG1O2aJJdXfpIA2hG8KWK
Y17oBQHqAHyDr7kIHYuEoRFCh6F1N7MdZ7MneUB2mjjIXBPFWqPMAWjxTLMy6BU97hX3l10cUZv0
RdyXz6f6i0gInphO4MJtHMMTLFNlTwSyPLuKzPNjPl1C4cXLEIFDpsqOst08OXSwTWL/9ND0xkDA
PnQyqotYj9k+iyzVbU7SSKWhSYNqFaUrpIy1TjBZL7VtVSAkQSFoFspzXU0m2g882dUFSmJ2xN50
Hz1PZk95CIJPtYKy9xHneanaqq6TyOr03mBGCbLZlr+iWKOtAqKCRzY4cwkoHYrIZHA5YkUX0Tq2
zmnP8d5bvKw2hVpKXVbxpRnvNtIITpQC7AbdZQ5kt0e6VjwPw3RBycR2PWXTblBADTfMTbo8TZdL
h8l8GEhHXg35WOYR7n5YY8zTAoarFye+gojMiRjYAxT7bYQO3QG969SCeQEg1AszgbUjhlVpnjQb
iA086y/wm9/mOkV004RigjXqmia9sdz2n5rQQ76/4kGJGyM5LUl5IW1TPKhxOqRv2Ii1e8271n0a
UJ+qznhDWN3l+eWYq4R5dfc7tMju5SsMWcEYXcZVlftmfJLQzY8AuR3Inf+c1TF1P69vtQmturhB
hCyzMLnxdDk8AyeBH1nGGh3d27luZ7ByM/18kNEZ6eVUo6f585gxnvirC/NvWcfBXaRpCABpfpBz
ICDHMh/TBQmM4MQhmme56wou80jSLOj2PjHYnAMQtiCkDAtbc4czzd3vme4oWeJAQy+zMVQJ1Dwe
/lik1frpcQ9ktSKQtn1l9Y2GT6TzxgRDF2DEQ0VFN2jkA73d3Kyq01LwVDbkTtouIY+HZ0kR/xUm
7okABgY8hoTmG3qXEkTWGzZWxE3i6hiiOPk6tDRdYE+YEgS5pj6QtJ/bhUOMR2RRmh286zWaR9jk
nkX3pYq8TjYAMuijphmkkty/M2boqYwNmgBfk9DEWyhf5WhVBpzRaNIvu96R+5+DAq/2YNEHb8ax
d9J+M4qH92V6oxsN9IaXeKHVv0iqjMjOdlCieYnCOo5pafG2/0fpceZjQ97+8M/3klwI7S8A1mY9
yjFd0Ly6N7Yr0X8ha6aYhwyUVLtVho1e6IYwL5o+edwVOH+TxYZEaBKKJ7arKEmFexG7s/rM5a/+
XWGJVmt2XqhaezQm6s5yuaIkMaSFofBCpux8Vyq3UREY6qceD9HZZQu1XQsxo47G7dHZfXtMR4Q3
tUlgWuB7ba5/ZKfL1ujAC2APxvYxAP7o9FUVVtC8BUIUT2Dp3vZRbs3hn04vFH9lVDYJe+ayQaDG
88fjoy/eTiu9SXrGYw8dDcy0z55ZD7v+YGrEwYB+OfI/+Oziup27empO9DMQlgz59+Y+S6m2JHD5
0jf+wzHC3SHiwRqfiu35mNuwS4rbi8fBiIjZCG+wn1aeSij4dryqSb8g8kd4mS+E6wFN0IzvIjCO
fR4q/WeBsZw4pmnW/9KHfoB8kQTpHyP+0ArjLfKoxuiZKeNt9TvFITAQ4TGnqou/4TV/JmJZzzrz
qzucgFmTr6zxxH52ennFeEVJA3HMoU5HBlOxN7r0RDIjn3WOwwfB5F1Yocl9U/0/o9FzEnD/SfNv
vxVN4YBek/0B+NkA8ytqNDKFlA5IrEnaBXi74CIuqfE6pZ/u8C0M3t300CU8MLBTRrLWoYCuFi+v
zCMKeWyrcGhq3CRyCIf66wbVMb3TsSJrgVaFqa6vz0TNd2Xf5GnxqjnzhbJnX06PtkaYadRQS9Q8
pRAwuE/acnIlM94rAFtIFl0i67tBx3ddBcbAce+asut+W+8anQ2m2+XZTjI1qLciobK5G8xvN4bK
vIi2aG/wHpDLt4YvNQXLl6s4A79EDfriL7iBdfw1DM52ZAEERip8XadSOKwVOCwCs3mnLR4cVnqr
1ErqdnihUbpeDMvDSaHXhU2KFwPttUstEytgQioSSnydNFUpuTxhYmkAIiq9bUEAgKdSYnPfBOTr
KvAwSTQi7ttJA6nZVYEH3PRCYqJUyu5OSxN+RVwOX+B2LbGEeWRmA+A4/G7X3KgC1qrn2/EWSHRF
DhTRatFxMTz0Z6LcJDP43jGDd3GVgGD7i/ly5k9cHSR9ujyT7JyLM6uhrOtG5Eas7BE+uGJi/znG
TS2EiNMJFQpkojgm2xpIvheo4wBlEdPLFZdFenMqUkYWfqN4JZEIMTFMUR7rP0X/cHq0d00Fac4x
yce07fTY7Gtkh3edPbV9bSVGrBeKAA7EN9/SsdcFpGImQICyMnaSvmgNZlgxYzP8zgG+DsYvM/Ko
E6Yja8uvo/cvP8NxTCqQ9HIYdLA1DDibuf3ibBSM050Vyd8kqJP+uoZNxo/htwu/+ElWU6OeD44D
u4vzodQe2Ap6BMkJwwqoT5cqUBm9PWymz1B4IiHXCsaRRxY1Q1FRa/7Y1bBMc+QoATINTcqY+TEg
O9w2qPSLhIBoGInZ5rpaIszx/rlju2wC68nySqJCd2iTKLD8cmWh0ePBtzTdo2+Srmq0sanMmFhE
Uif9Fx4fC9XerzygKpnVU7fvwuGw/YW1NHU5SBK3FtAjmIG6NcIad0T1FjD4AaPvkkpTstt01E8q
gT5QYd5gFUVx6stDFjczEnRsQlx6HQWzcYBCM9SaM/f2ycr+n9wRbmf+RKvJ+9l7M6AuzPhGhIuU
afRk4ARzRcLIXyo3A3cNg+5CjajMt09BY6R68+gmPmNS4Evs1c03dcPAJobXxT1/g5BhOXWnFWk0
C0umbcFLKtrlkiCqzhEgSv+C2pax6v6Ez0eJbrMSoGpGXUQWlnJCaIBMJ3bFmVDCLyoDZSA6ajhx
FEOQpWK/T9a/dXHyBcmOaC2+NGvLlx9pAgy+ObcWYfNtZAcYkS/2+89Klr1LLULxGNGbo2KnsI8/
Ub3pb/W1TQ0H2vcvHLELVZcwjrMgro0jivuJhDJzyH3llEMypt35B6VWHwc7V7P0XGiv7g3zPRZM
eyvtytZoTsa5K82WVMafxcF1kYBgz9y6xuEn5jFsVQ1QXTmI2V64yuPCG6CilyPPOAI/YhWTvler
+PAfi/kEhawe0qdGhPd1OOTxbITpNqDcXVbXQ8G9bVtZ0BTWFjSoxhF5sFbx1jXPGT2OGzKxerof
/OFJ+6XOCb8+4ZS1cK/qdbq35nxpG8R0umJBQN4AvRyv5x9JGCSEMDo6ycZ1WrEMXKXLh+bSIsxM
76nEEhilI3+IBx43uaMvPhpno1AroEFWrwkCu0QyZgh5300+SvOpTipM7B+/1SfMrupUs3+qSRAz
Lla1n340cVreZB8tivlZY/R3QgWQH8IDJMQ3nMr+jEVI0yCGcGdC8be3/GOpG/pZz3ZDS+z92eHp
/pwwCkzH8VdWfqHNpg5pp3iCRx/JdTrJQ4G+fFPJ1ZksDd/h18oas0+ZnztaV+2s+/tXTOnyKioi
ZM91aZijrvFh9G8mygp0QKUUIHx1HI8yzxLjYvrk8s7eN3RIJPnr0oBWOA/So38fvxTcEDaq2ABK
tJ76KahFNczHqosiMql6T2nzGec7v8fpTIv9TQYCVE15keVDZDzaeMCXCELpIqGe6Sn38peYDcrj
r+Q63CSK8ub6KYlJHMD7j1ERyVpcUL/fkiSPcU5nr5HWydwCbrcGDQ6THBEe1Z+oOkcHRSlSV2Iv
ktFHh95KFnzlmncxLLhuUfcQADQ6pVd/qB0hGGy5qe4NHkAleK3mqlNxgsxRkIhiwFE9Ag+A6cVl
OnzViHY4OYeSXJ+5oFRxpwHgeyVoEzT6in9dMfnDqU6yjhIr1yoOcHj9KPvYNOCuQ473XEpAZQdi
+FLQKehhLk/oaCqLd6V+gQ02Fkwk9wyX/Q7xu2aphDsepdYxptMPPN5wqL1OzegPl8u0FFvfoHaY
fyYhR+tqOrvb4r/SRclilFAs4EVjf/ZM5i+301BtRsBro+gyT3PjovOGAN/2OHZxyfzZfnF8Vn2z
5N89pPiozQYA6J/w73Mbc/9nRB1Z61W1hvvPuvGuMTyM5xatJY0xT2B2J2Zmqh3H6TdCfHTM9KDm
Fn0ETCw/V/dwRjzTsemCsTmPGLg/vE03pQoKDotKs4CpGYhkmIlfd+aE5ErGsQxhfM8MGdYeCZBZ
Z/8JbOwWwq1QPpTY3I+FTgzOUpMeoZK4p8MpOnC5tJSQdQrNWtqfcohWWXbhK8ysOjL6FRrPo+r+
1wOZwXDucHjw5ApGbMpdkvwYKSbTC5z/YTyg2rlZIuqsoBhThR6UdqXP+rMWtDHUx8Ky6ULOvHG7
186V77KPyv31YJUiYSqRtd/RW4G1Y4YZGK0ZLAfKOKpj4TNqCYcic/RjmItDsaWNG5Yn7ESTbiRH
QzakxQkmhSu2uQquhOlP+bH8GRUhDJW6pccNSHEqB4ebYQk04MRBv8rRCe96qY1NyKPvRhi7cCdN
CMtkeq7V/Lln1OfpSDIf80KQmODJ4Yb76LqNSfEmL4Y/KgEf5Um5kTO4Zl6qdkmwiSKnuig56MgU
ij7t5f0QqOtfOdYnHj/PeDYe/xzIOlTAbejrwJImIHlVPoo14QKQM10PQ47XjoFxBGu7cZNFeFNg
YPGREunHrd1S8O9mkFlxue+vxsb+rZOzG6bnVb+YNRTS5LqXIfP/OiMllfK+wtp7HRKdG562JUEk
QUSp5EmlNmOykLpv9ePvmD6pqATak7aJbP+Q0Y+4VgUYTbXMBDhWtYQ8Qf6Pzf41gTkci/4RRhTe
B4HI7slyb+MxQywjiivBOyNnsi1WV8T0cmLYHuaPgRBI1jxhCNjP0sM+EiWxwYNbJJDogk6ZZr2d
vfQoN+Ez3BroFZOZ41TgoaldnLKaIa57lDT8U7uHoAn8B8KJN43PSL33RaaRmclfduI4DQ5CTpWF
ZvNDBGUPK4uW9yOExVaQgwbBDevY9KxFlkXVkh2lUY56kyIsMEmH6Lq1SyIrrqNnZdvnRt5NcoCn
KfSCXeKdbWzRGusH9sLICa7bibs6zgK3zIdCjVuHtiCVoTXhnbsqA+UZ+YuO/c9hzKqDW5RDAcY2
41m4M08pNxdf6+SNSo6DUJ473Z+GKBRMJYGrmmcSJfYUofhSFw/l/InMqaxshyS+B5+6sfmLenIf
NGzFMYQy78fotEFIvFfj25DTKormiT9bUkZEVV+WqIcYx72iJtzqvgRJEwBVg+uSociJ+wxGzC9z
XI5UzMA2Tt972O0ecRt5E6Ur4cCzF7M9eZCU61dbK8VUT9AXYPNfaFmB5ilu8Y9z6F6QwgIvxyQ8
3e7TnupukhtOLJzeMWkWbJ4qCPiyI8J/QR4pPcc0k4KV8dATAicv85txz+Swpc6lxkCTEoO2TVeL
csxttMHiW5LZ9mgR9Hv4ijFUTYCNz9UQta8vcPI3qbKvyaOaS+F92AILuCcamh1Ylo4WJfBYfECI
5EUMjxNb/q+iqmYeEpxCdESWL7CItLQynzvuYzoIphUQBT2yX7tlSkJ9fN+zfsf+lGdlyFb5P5cI
bYDoV1d6cCz/IG1xcXZstnTwVbGfh42Zt8nx7M86jMTkzC4u+7N4E6Mkn31PUHa87fCbs+Jht7FM
XdEtIkQsA8G8kY8pWIKisC6xBnV/f4GHPvutsi5d8faBxfJ8+m/bbtUGpFiVa85v4hwXd9UA7rSU
nxRbb0mnl9ES002/TQAZABycwDBUuQjXfsQsj25pr3ellY+m4RjdDkep1ntDUFtlnRUGMgVtHPk6
hqW49TAP4w5Cn0Z6dVaZ0X2QwqEk4eHmvbRNvnGvnRjgBJJVsRPXRh+lB0mCUAc7Ffg4kW40m4Ab
IeJvIZH7qkwSa/kBtdqkTl16bmHVSo3Cwu0Jzv18un5VkLbOFTU/VAMd36E0o77b/IBp2Ap+OI5f
3F3geDoYHDoAC8SGI0sk7gyXxg5uj5HUF3iWgzA6M1vtTr5QKaNyCqcSWXDUa+9ZLNmE/AO87dQ6
oEbJrD4FbtzMJTsc9dwwa5zMa31rXKnJgV+lAF1ijsS3MEClPJbBdHgCLN3BnpwWbBUVZnLA4JJb
iu3bckygWMHoMbJk3qxD6m1F0JNcXuVyjc8q0CAlP9T5o8adEgjbYDPGkP84YEOeZhXg9Dyz/jn1
A0zWawgZSaSBg6KojI0RLpjM2TM+CcUBHhNqQhvTYoLrdyL1M4kDqVzbNIqVlWZpbhcv93GXOzw1
Rx7BADGlxtbkB7tqB5tmZFhksD17BDmpCGU4oARKIy0rq6lV6UuEl8Cn9rGliAw1jzZdLsvkhT+Z
Z9fqRQ0pxGRCl1M4IchRll/FAVrijQ5W6ryloAy8V6/FVSy31G/Ac3IuPHnz3jDktyNnFfkh3wtl
ZlD/Y+QhjcKGlqlRyGRJ6xXynKVn6wwmtKUXPfF/uYHZnqF53F40lJLRUWzod7OxyU8LSPaZ0Qbp
ROUvqHMNbpZu/MccnIuwRppRvglDon5GF6zA8k2CLSM0z5ZICJD25lhSnEYp+CUvPaedVLSEjWs8
Nz/B6UiJZHxq/y0yLoe3fU9daiOxBsJEwUeEvexWAucchipDBa6AvdquvgQpYXIb9SyGaph3p5b8
ETCgm7P6cW99i0Kx/eN0DfDaLLnS4mh6s2Q6OE41dFBdveMjTRIItl4AIHUzP5g33tv0j+K6LB6P
6r4/UXgdwbXtq+8Q5+CjbhUHtPu8/93+DWhr9nRGS02qyFa7aZCVvHYe9EkgsLP1GpdGqqCIye1u
O662LhDAPXXkjANlEj2Gm41NwGP13s+3TMEWWrdXxtj0gTHGcEQNq+Y2OYqWHrG7qdd7iL3TTuFw
hi5dn0vnQxnHSXD3AkwEx/Nlpe9Z6F0BRVYK4FRReCMChlleRnllSmuq8ZNXV8kTMXz3bbCX8ehv
E5c8nJLjyIt5AJTLem8uRLdBQz2QtLxt1d1LM5ubM7g4Zl4jVgXAZiXgdaVsokYwEdwXAmuckJNC
lY7p6QzUpyp6mfVEuzBibYjoDGcEzFEcm5tAr38FDS1XADvdpJCD042UJqUQ1XRH1C+p3EMenGFj
ZyDqI/8eFuQ3W51PR9f3h/Bu5sGy9YeY6ca9wy7d2ftfhuG5qDXRF+J8dauMbA6h8hh5AE2HF5sI
+RUlHHpgFejvQNQpG5lEBEOj4Wxc+sNzDpWgbgriseZyLq0NeAiQAeE3QvNjgi3/S+b/ezORLMMf
jyF6IIB7zPjH/S23uNPLk3lzT18wnWerPhOQzzpQjKdFzVneLbv6PRYckN2JJqpT+t5nEBbVJAXe
Any2qjCfF2tfcZFbfs82ENKVQTxw0RUbv2Sn03BVG8QkUF8U9vODz6wXo7lFCejKXIF84CMNtU0H
rvD6sR7WYytk137+coBNlWi7kjiKEJYG+9zCLtK6IwG0cSWW7y7ST++JFDs0XDaNHyRqQeFp6DjZ
cAhupnLcjE+9rWOjnwtcQQgOgat3p0qbQUS/Y0PncrVph6RuHvnsGcnOYOUg9TbCXhL20t3V9mi2
o9z5hR/i1wFv6Pxx+kRlb4CHwEOUO33S2tbiojRoxlk8jIR5a9052jwyB1VHnZ0AvxoWf3Oh7i+z
dsddyGQWfEKaNqOMgOUKSAr0Ce1nDtqjuO2mpKg2o6J7SXOK6mdju4y+CA2Fl1qXPF/kcXDIE9C2
w5wSn82s1Tav0lZhDZFghvd6lATb5THLjnNDnqF6HDnaPCZmmy5BoD4nJfIt6eUQ+uncc8DjrGVI
CEtqN8ogWXF4TCLguKI/AGt3XfAhis2tOpvO8NIAi/9g5lSWPv7XkQo/UX//m7GDJIGbVZAF72c/
/9VFsZ8w8/H+848CmVO7vgkFwTkMHBNmebjfaAD6L61U3FnGuoX51rXQBCgoD3FHdQRnyLvAfrlX
nUGaKwJt3DXd80ZfaoxveYGsnpgSakNFs/VKARmmMnNwmNjpX/5CMqeOwCLr4tIfSgCcaAgknLux
kyainLuuUYvUGosXYfx6H5ei57UAkfeTkm0HObnV6p4Ea08lD0DLzSersPkF5pRmMAOxteGyjeHp
FSS8kXz2VCEzUgUwju+sVubhtctk6CLr3i5Z7AvzzDJpU0ek/WghH2sAqMC/37HrLWH2hgALew7r
zCuu8MSzaac8LOCFHATb53oHkMqJHY3POr4a2lWHgtuO92HS5mPgK9SehVf+/i1bn13XIGdRmfuc
JB3qEf2HezEud9qz5OeWpWFu1gC7a8asm5OwpXnVd/M8gR+Ssr8tEfQrdhL74uw+05nv9KwD2kCr
0vsQ3aXyLPPLeUU9NaJ8CdhffqHokOhkujWd/Voypdqxum3teILbsZM6Dip917xew98itZHWTzD7
2FWwhs0o+A6fgWJIpuON8Xms+qKysiA66LH3qj9oyajsvF0mZgO5PBFxCXEYUnJAYsjhePhHEJKZ
HUB/x11d94iHUf8xP89szuvYL0YylbgZWyrMo1yI2G6wCOhCI1Nh3uDZYHECktVvh4Y+XEaw725Z
5hjUP6UviujB//7NJ/K45XB75hFNEfEiP//HHKpq3hKW1hOBezhQFFgWoj2QTcGBRSOiNxk26Y7f
4YyRUMAO9fx0l99v85FmUhx5yCYMgeZAJTv7ntdnb5hYDoJIngD57ogpTediKx2BD5Cor3hq6fhc
U5vCxYM2wOSq0Nx8w5kCIUToClxgD0kjKlSPpd7wY22e57W/xI7KTQd7j92syzoU8mJBhidSxbIA
gm5M4kxKGgwTjyXSBq117jhCoPQz0gTvVKbODN043KUmc548cuBdPgcd7ZBUf7RXgbwwdmoH07Jy
Io+/1OUQj96KhAhW19vnmBBgeseeJ659ECzMzf9Glq6G3OYeCSU8KYRlCrvI5Y7HCd1AxRSv3BO0
/2Y//GaIpHhg+YMNFJd7vD6xTZ/9ROqY+Fki2r6ZSmw6OSFtm9noiHV+hQgys/pPnQkdJE3+ocuo
TJNYzN9tmJhIGpItO1+S1KTjbyITBwU8aJ5yYqE+b4YjMlm7ouBTEjOzWHsuur20bQzdf85ivJAp
ksZlJt3TgvuoFemc4e6KxgmVkI6c4eWnONNs3GRAEBziZL7l2iFLrjQ7BFbEYUf78NzHpmgpFByg
ntHfoahuO3u25CT2LNiXl4edgaYId5+q0nZsndZJJU0/R7cq4V5x0CGdnY4nEyhHf7w43nPdtLXD
CYjWhraIQHdItssPkyELhGbKMGyTH4CNsH8Ld7QLxNen0IoE5xL7fJFDI1gEpIqe2Yc++rjzF9R/
ZU3KtS00dmoMgsfqt9Of6BHo/s5xGfjUclrGJG7PYPyS7GYie/VQNVO/n7hwZSKn6qws89rZSkbf
N3Lf0Lx7KvIAtJIPsQO6pFWujVlKu+H2Bg8UIsLhyQvAhlDXbRH4uD2xtFJ2pAc/kddPPpplz7Mp
R/r2DBXi6TUMsJ6E9oQs5i73uBXpAcPF+xfVQf4JvRpputo8o7sinbkeKSd/LJZlQ3nzX+LZXz/g
2k+nfxJ9RgHp0yh6qMOaNmvHi2ZsLK/wrmnfhzxd9iZZ2VNll8BzvNRyxilvwAT2luBv6czaXron
rb7VAG6+tkHs7qAA+mnI3CCLf6fIw++PGtnhtjd/fbJQ20PaXEFWC67O1TZ3cokxHLELeE9EC5Nz
G7vlvHOOH+SmcrQNLQ5l5Dunhw961I2Q0ks5RVxAzjsfXW67UYcpK5yeSFNMtbA3qCBniQppFfnn
zwcm+LBlb0OZNeZPkP2+9C20qouQ3IcoMzhjxyDPk9U68dnpPZ9AbqCWCdnZcH8WY02yVwy5Onj7
zO/1RqgWeV94boQMRME0w3ZdgQPSdyMRwwRpDYIbLS3rCHzIh+i0jxMT9POPD3d2i1nMJ5UmmEkG
FfWAHUPTwpSJg3giqaIViq24zqsqm4GOVx1QB5ISTmsR2IejnxcbaGL/kBiTHYBsswYfFDsym+Eh
d3mKtozniUkqQLlX2GHwo5if6mHrLd+4OjTpcGJq5jplii0FViYbRr47uHO5Vp2YuolHTcDfIfE6
6MLdBrKA2nqawgCJtecMKEarCi6td4GZ92cOeZ5R/WhA6dh0qZd5SZ+rTkCqhsGDl9RVKWEveXEI
hUyojY1K0vxEk2KHblX7jKxt6KpTUvP/1CEITmL3QCQJvhZdzC9sxKlifdzt+U74e3oIQ5SAVDOr
0hRLRNnqtzBOJ89j2BKGpDNbsf7f6NpykdeaNlqKy8+PeeDjODz6p9hjAzPR4bWpxKI1IVxueK3O
+8c/rqJoTKhUQkFgwXCnHcwQGNeYYkskbxqn572MJjPzj1HRwA2EWej+JUO7DOvpLQ7XldGBoLLY
8oepnkFhUGxXQDXXknfIALWqsktA1uMH6JNHNb/yhRqWJPQSdELuOFgb75ATDR+c1X0LHAPvOkyS
C2Zk7kIRwvguPApFm7tzhCXXZ7ZBeB/v8bZjittD03vZBO2bKrk0pNQXPwSuCd00A5LwJ1gzhhyY
cadDCqNrSAVMnubcGGjHEclaVeSulaeZ3ZjQEibRN30LSWmu1LrveHAlXgoDv8Q/a7ZqTb9wK3LN
e1auoF/17ZhNWX1T+uVEMNgyp3CA5C+YYr+8EJ+lueNrTxbfAZfJ6bT2MWdVRbSYW7VBNzBugg4j
O80mRTgpQ6w5POdvaHwOJTla5Ws8RRZAxLZzOAaJR849Qq+CuIAarHL0BCh/ChoBV8+k65AkjPJI
rSiI0kyJkRo3r4uhqaY0iV0gMkBSKh2v1r0ZkP445Jg81CZXwVt9kuMknWvK9T7Op1cAr2k+NP82
9P9+OIeO8D9aLYktrzgeLxwrrDDiP/MM7JDMmXUJnIDqLBYXnIER+mPVoIm/UGt/nwPKi8dT91Dq
kX49+QXK3rUWySClkn9dPcdapPEd9Hcsn4QCsSIMDwsDaA1zIpmY13V6VT+a0RQ0B+sZZ0sSRu5M
DZhRrR1RBYt2mUpZZUsFpAtmlgWtH9nL06RwupbMm+NuuMDBNQUSnuV6tuDezHxAyJPIgWfR8C6S
UokQkdH7652i21wm17l9MfFHLon6enOWEJh46iHpG7CyHjOvwkyL9QRH+BDZP4++mAF6qowNTw+w
qBMgnm+R8TAhv81+HO9wWXZja1OPdJbgFg5wg8WAR/JN/JT9BTu//N045AveuA6DOfuuuywxvuYg
wnuc9+u2jdPQ6/suBzXvj1AWEUnKaxHArlSb3N27aC5r48tmnG093I6EkRJBLP19RIJK2aX/8ksd
IS9uKxy1/5kEh86n6jN/xib/SlP2E50Wjd86zywFyeG5lGarnSnqScAs7WjjKor3wkyl04OEWZrp
spdgYNv3K0kPiLH16dTYoqN0mSBY95LLvT+TUiLEhIiNvw2db1oPGISS159aMzPpIZ6rkfPNUwVR
XarL+rEfegbovV9pECldheAi2J60uQOZyux0YYUaRF7MWHEHyVq9mBgN3vOsk13RHNVkKiRol2sp
GYYD2htFgE+VFMVZvBDXxoBhDv88QLfID/A7HegyDxjTHezolzXTzTQvDsKE0uD1zRT2W/cCkapk
/G3eHz3TSTTQw3hkR/GM6v17rHxwA76j/BwyEBhyVzw7sM/ofLdZeUEchvYj8QX76jUW9XvOBewy
45FSYpucir2tUQix+Zeblr+aQhNYYD9NYWFF4/knqXZYdUNVXLHQkYvqs7s2+xOgJvQITzG+SrND
VcvRs1Ils0IRgzx7IQaeIjQW2NnaXtToVQnRgO5cYhiCucsEbkTnTHTPoYHALMQz5Gt9EhxniT9u
GdKYnusn7OD/JGvfsXbVWuvZn5nDI14o0fiQga6QE/Z9iqyO+3Zj+CI60HP0v5pN9uu/IzonxP6n
bv9U9y4lJxnrTts+1bG2IiOrMbc6/9oWwZhuXjlxUPQHRSHZh/ewgCNhartr416noR8x47zVJwQt
yHTRr/IH7Xsg/GAaPPF2FzX12oxVMBYKC0p8t+uuI+SjSVYwSXKnfFoAkllRmiTIZq/xvsWRjqpd
4fxSJwQkB1U4t4lE26w78iNyqjH05kz8BuHque4aW3HylkK/qbwHE9tLxR/hJ0JhUbu8XShktPHJ
NrM3RPgR3HPWMTYAeTfQUBkpdLther7lblpkm/oTQD2YOcaiWaqPt+MBgdge62f+Yxoq5swlbMdk
3H7Pq2uMUWxA+T+6dijqFwXvdBT3MLTu92zqfktKIxRUuotNlzvQSbNYIULcwd8aXNt8T97V2WL0
+andXYcCtT2uQK2A1DAIl2B8ZQTifqYLF/nfxBRpLnXsZRiySe3Q15ZXOTGEbwvawzSvo5OZ4U8d
XRPxPebkMxA2uLqejgTP0Rt2UV6yFesc9Jz1Fmvxxca3/VM0Tm6Kr44VbpbYYPu4QnyXfT2FgF/z
SrO0VJ19eNR2xx/nQEGyPzJ/5x281vbBNpcsP6/KmuwIt5VcdYkOl0DMQuWFwYZgtmSIVin7R661
hFlYHjTlXWAizJBayPDx3V7MqegTIq6suSL4MZtbbLkgFYKNdGB0QraKdQqPhCQSHHE/b5cb/oHc
o5MSi05D1zqQ90V6TAOXxeP6WK57rB/w9VTRB+HRKJTmEZaA+k7482cV+dUEpP6NSWEdZbj8B21t
gUi3nldPLeqyMZm3T7f4Ax5DkMFgmjjBNUEI541UUK8jM+rJz8CeZN6oaY5ddQRmcdwOJ/8Lqrq5
LgSsFhG+O+ljPHPlSlxL6eN/6QvosPj9xPpuK6cEIocK+VgSsuvtmPKedH1cI86/gMeokc3Li6up
jzSNz1Q1RwOqyKWvdWzIe/I12RkM2WcvGUn2KUwS3T/Cb8Q+ITq8Qpws2cWOeNaa7Q4PQZLk85Bh
ITkOJxeudyhiZHt3bL8m/UEnybrUEUsG5tBwctyzP51fnUFKCTbdS3GNffcyIsdyxrworybRDNtq
3pQ09Zyo7JDcNWS64SBlXfROmtZhpjRnHEN1v1nCKXXUFFE1EnmZxsx2AVPr5iVCcjnPKDYeuyy+
tt7kpx03s2Q6sv2GFJ2i4HbEeciGCs+AtK2CyQ0CI/aLI2I+oB2d+81SX8in+v89V1QgHk6M/zrm
kMEey92fYilCTr2Kt3baB2W0qB9znr+lek5wHwN1pDZIUkW8PwA/dVSmDYUBIcKZi16Bb221BpnZ
b/CxzsIcOwrsjyd0IJeC8ueLqFhDWq4wgQkrkoQoZL9lWtYcUvGNfPl1PudZsiwPfujUxu0bI24C
3bkHLAE14Mrf7w8Ko+mVoMe+KlpNBjcK7KEpDbwoclnmAqKDqByecviHTaCqZO/fnQoIzRgzLwbR
3nya8pe9sx0wrTTCLHb52Z57YH484s0NtqkWrYvU96+uZQy5GuU3MfGooeADDuAtP1gnpyiLoVs2
cRQ/EhY0l2jKJ9gipikkE5b1/gFvflV+Dve/LDvOoszg5+JsdBGKm8FoOcWRPUMRrY6ctI3iX8MH
zFietjz8THg/3puK4/LMDf2/L/fwTx64UZsjx4m+t6bAx80Nrr4E9VJlw9Yvfkk9BHLN+8xsMMyl
hT884NXza9mO/MeT5JRX0t4QRDuxjTPYjXtj/7jqAybRhgG2Byg7ZbHcfAFNd571VSzJvWtvq0If
XblXF2G9AHt3oE8NWCXiwtFOLxaXXiEYgFhjKxHJ8qFc3nrAt8xNAyOfn2mF9hYQrwFvKX2WZnG6
7tht7y9k/TVJ6YNxZxi9W06GjO6IeM3B+Bzaz/kB+mc7AUcpLTpsDFynxs5poDy4T/l86VZP/3um
Y8fSNitTrzQjIds7TRyurKliMr1ZAx+Xl7Nivl+RuHq581RvmHgBKKHTJDCEutn0sZCO72h0JZQ4
FCPusciG7xi3mO6p8Ja7lSkXSXorX5UXZXACZJTWUlFrzDmq9xx8rJdmqNkDOyyjytq1LUI4uKYJ
KQ3VIsuu5wthDwlHY5AlIbmsGp6Pyi4RU4COVq1X41vIUYFiIGjdYLSdK1lziitpJ4+KFk7VlFkL
2+ZMjsGz62qicXMpCrFYupYZIFqsFHJFWghpPOtVvuqP3QQ/OMIyt0Q4etNv49puD9CwioYREWlE
LYSB0JPHRGXN1G9NlHF0vRmgZLJ7c3j9K9HxRKiAQeAJvE0p5cESQWBHExVgyu9cP3psDfDElSN1
tT309xNOmEgYmDIdzcgtmXGYtA6kJOaSR/aRYbgsZotQWszPtdG568Jr0U10G72weWwm1/+2Zbye
wbaHHplGugfOxvjCLyUYNGKkHbd6q3K1KzVgyS4fo0qqM5AXJ+wqEgx5AgaRHTo+DaNX4R7mJBMu
O2Y8ceh7xI1yyXUQZ34ekvMbVK+d7QaaAJhsTlOFWv0v0hBfaY1Xtlws4AuPritg1w9onAqukI0O
Q5VcpPseJdn/9qkIeN9uQi9AByom646BpTvxMn5EU+LttXH64DhS9y5e+FIHEzjyHNSNqIk/AEDU
CZ/3cpSP0o9xzNMLseH6XwWGQrVAgPhhQCd16k6aLtfd+zfXReMoo2MelpiYZ64l9t9LLJ1wyh2u
0Bhgxee2R5l31PcSE86VgJZg4IbMnjEe2Q3pu5Dmxx82MiQ9gJYFR9OJ5YoMmip1jTgl1XqgMVxZ
dqOWQnZOlC95UGbZ4D8TMhQkl5W+BF7Sn4SK+hknU6iCXWJRBFC3uk57L6leufK7Kle7vnuODg/N
GryoLr+ziW9b7AvgHRD6LCr+n+j3TtyCkWn7GRxAVYeAERtyVBSUaYE000LnmkD78dmbkGG6nKgO
qbWd9kOyVYYB/t9mbImIblq1J6nP9QDCkmPhYUC4wVYgIjwe7KGKiI6dT/WnRLDNZ1B58NU1jl1y
3yHumVyO2W78eA4aIm70q+nwfD49N4pcrofsewUf4l5Vc//n98oid2rTn10Ot83caAum4zNVMvCs
ToB6jOjpAI7nDqVlWghReeWvEK79PJCI7ze4wk7lHql/PVMd1VIA3Yg4PYjErE+P6I0U49PsKwCm
YTiiMkrrygRhPaLIwn7Wm/xNc9q09hH9JyQLd65g3DCkWVit6m44BjbX/FNnBkhVlAt0Bxrj7qcC
U/EbJTM27o0p9QfcRde9Q6tzEbuD5ldwLaGObdnnSiA0EThhYb1SH2L8yYSPvF9CBjYqKajgS9XD
MofA2Ej6y1ZfG3ypW6NHUPxanUxQ5g16r/B6vL1j8J0g/vdRdrurWC1fSsyaQ276lveGtdYYZv0Z
r/R5JZDeDJEWsJD8AQGJDS4vTH2zmNWD+xVLQ6YXf9TDYl8dh+jHLWODIIiy9ZxTnhTyv69srcg4
LJ9Q+ZR25TsDbK8pv9Sg1ANIQcnrU+rEf+zDBBSlEdXmtlwtumW8gUA1kC+8+X4HDj+Z2Ia65eAT
QBtMYZMUbnvGVfsItEuz/2m5xUYdzlIorQ+5dTQkmGWqD/jenS6kL8KFM8WvMZYRrTzK26P2s2b8
j4DczDi+wOk19OQC77nPmMXoqF1LHVCMmhmpsOtX2+jf2ljPaB4nf3pSI8e/rdYC/V7hXfux3Uxc
Uv2lsHex30X/wrfJ3UOHVAd0G4pLtu2VHycuffXwJIm0tXdhMX6wjIeh59ZdCavL/C7w1JJ3Yr4b
cUQYwA50CKREcz1igqxLynYEEDDz8IofsXXfnQkFgf6R+tawPmqWsqft8dUUgmtDOO+J7dBxnKJK
81EnI8RL5KA/PAonUCVdabB1LSb0h0K05ifYRje2JGi+8WnLS+yGXcfF502vnHydAgBJHqAFDrzK
6GeonYGKa9WDXBUG95XAX6TA5V19VLnv1X3PFWApUzmxRL65sLcxkT01ljkatV6+aywNPP4R7l/3
cRFocmor8GhI/lPBMB1gaDw+MXLuKDW7qfNeXAKJTJ8JL8MKZ1U6nmF8HO8oUnsJw1GrHCrg2yia
EyRGjXuFjgssG+nPg5EwvvopZl2F/OrbNYt/v8AShUcbXp0zBeESuZods0v8kNOR4FWVXjmgULgc
9joF3FLKXnZT3pOPBVwZv5GsUU365ahGIBmM9n2SNn7czUIGZi0pzYOlwJX8l4Ow9w8IJGGiNEfw
jEX8SoFRP67avf02BNIKmB1dxJPJHvZaIF18K1mhDrOS38orwFsuEenONWKLeiM4LF+LPuwCnaIA
+s5fBtx0ntn1KFslRBqfjGbgAfjjNxgaG4SSjQUvNYwJu8reNYp65JzQr0zEqFhY5bSqkRO5bL3x
J23oHn6c8jGQ6FFhEqDWjQ+TKNZE2r5Byo50JB2uroANcL2KZVi5lHktB+yxggOYKQJZ2h+/Ti5F
3fmwE0JHE84v6xY5LDLcAqMqbbihItRK/AObQldxuuCBlnCCRYF7Tim7CWBc7L1WFxaIIj//ogA0
H7B6Aq9OFlwULW+1sGnmN+1VjglIpJl3QF+RVynWL3cIsVJE3V2F917cakzbf53gehPcNF8CY0c+
IJQEI9tIWAhXEysst/RG3zz93F0VP9pb/yhBWb+v1ZCOSya9afNxT6WoWkJ0JspxSx+RGMvOPB9j
7OeaU8U9GMyI2Vs96hByNG1cn0Gl+JZClg8noFtWc6Lco+KBiJjJ6KZDa1w64aJ+ErM4sp/KkJxA
y7LN3GS3/ICsU2KmVOOr2l+6CEQ1Bri79piyFL+JumXX1EqWd720CAeIVMBZ6zwrycz55FeYQCdj
i1Xu8Z5FVXsvjOarr97KHmUDL50BQheWOvZu88B/bPDvuC+CD3K5Y5eosI1wsjH2uiW/1bHGw2ap
EYr0tboQR9Oi8tUdmw/5HEzyYZLfSckEvKlLgWJCcu11MnZm6XSiFV6Dw5E31Oi8hJeRAFPlLYjx
Q4kuEt1E1ivinQmcetAHvEjOcn3Rcva0kypJtZfP+/JigH6F2AxYfqW5boaHdl4iY59MwDjW/+s4
mSbH/md3eArX7I6ahMJ12WnqfV2QE7tO4lr5FVs90s7iX3BozTNK1t4HU4ljfWEZbLRSsJH1Ampc
0Jm0YjS2zfoPBk9AVMkI9rycppDaa9pOKdqg8F7J1R0gkto+iCeVWSssT+nLkDK4/9MRu3HwYdIc
gtAwdVSfBWt8Hs+ug0Is9bjUk9SD6rKiLVm4f3vWDEg69UxCnmja9ZuF4YONHFbqO0b1U6ggNC0g
uxtPTzJ3gOjTJy8rYR5qB+4ovmscakp35gOCpvFJgJyaLZcbY0ie4JBTVznnMEnFBkok+lmSRzy6
0Tr/1eqB888rlSY1GkLbdyejE/7/nVdTN3QuAzbvjs6mfpnlKRLMjh//DKK/ccu5ESta+dHBhSXl
pqSr9n7XdO9TG8WEMRZODZjwzEm3q52e7w38pdl6jn0htZqYOXSqiZHlZ/PLcYtNKDOJE18jkycd
Ka65Ee96E5169V5FsO2otkAR3CaxK+JAsRD28W5W4JAIvcOqIvATWOgxn9UuQNDDnEemR8Yp6UbK
JDiH3gfoP/pyJV9VCHHjGPyta8fxsOapvR8ChhbzXvPS5/CzTaHzTSDwn3TLxjiIZg2KYPTjbI9g
GtvFO3+tP6ldEeybUTbdThb0nQQ7AWL050Shjc7qwosxWT+X28jcXkeWcUzGXzyx5gTHRhgAZZZR
eY9QFPDKP95ytWLItSEezjQLoWfTOGLJ07Ks4YMxVky1hRYUQn9l6epXaxuG87JgerxdJb+2fuaJ
JrEPf+qVTbEvuE9TEVmcmuRhkL3U/sseNYH2KVuNOzNW4IWJBRBW/Kuw71EV2sb44gE+6mdQl9H+
Ondt+ybaX7hMz5kRpvt+XEnxAT3zBgzhHsS57rcbqXkAheNoKPJMlYI12Zn0kDRB0MMThYtIk2Qe
F8o+fy6J9NKYXr+CJJsr289WfL+Fa1S86GHDzjXYjnlPV7O9tk5jjulnbTh+HyDuOB69Ii46MEke
KxNzVQ9hQtzrBcpMZnSHOoPVtlYLXGeXzscxyzT+vaqf7lcHOvRBO30QG2cEOxtJ65tMIy6NuQys
kfjLHobEJGtt8hQd67h9pDuCPNZcYSrbVM4rzhhaLwWIvyYVBMBjNOcGBrj6T/N9lfyNG9bfDcUR
YNOaTofoHLd2ui2ZAysuG37du0ZFXfHFiDXAZQ0vM9PFizbRO5eeqpMOQYKAy/8Bn/tLHOl4w5IE
+WHeaZUN7gHY6j1p6dI2wgMf3H/qdwLykphLs60o9F3v/zrLuFhrkSzRostPD1VnN5rhqD/rA795
n0OFbXInI7lFkTdXcb8gN7nXIGPrz1GJe/kngVtDKU8p557ImYZDPpxNm+Kz0LPcmvgzyO+8n7lv
1egskoO/v14KL+Nevwz+1sEUmOeuCq2Pg0hg4XDf/NLAOOKR7Oy7lQ8eNOc2/ZguZl5NrBBq3WmK
3soyl6F0Vn4usRTC/MwEeSHaSR6enPbjvZ1C9+gYTMviJ3+SVQWlJixZTiuMfEQoWyuR38T/Gu7z
5Xd3h1kfWsaQwY1baTChjm8H27OFJaM4bE2GpfKatyUpNWBEj1qFLwI00N/SLyFMIvFHM+l3mOd0
udvBkP+VETnCzZvH07MXWKC+tDxV1GOC+3Svy8ZKA9LlnWe4LNDsmJ+RSVv7wfvUbYL5d3d5jY9a
RZsmqhT3YEIQLpSHiSVuuLDF/fEM57GYsjZ2MML53x6noyGcl6QXfJ/RLwn1TDxnCkNs/UkbLnuV
V4wf8Y1bnOYMqgISgprBxrxAJ9Q7/q/pY/fzGqABsTaxfgjoFmclPMypgthsa0Tgo6Z3PWxjJqwn
kvFfX1yKfN42M3zsp/Lx7OzlcNKlirQrhEjpSeX96Nnoxv2LHEGyHP14iC736cWbZftDUE42SLbf
RwzaG/iEjITW+BnsHfT4bjS/+qDx1c2UtSiABw8ljFMpg7mbBBFL4OwbZRvzo44WdUtR/YxwxJ/Q
BBVBk1zRnUAgpMEaqI1sv7z1KIB9pgls7uVK6bcrQmxA9ndfAjqjERBHtYWnMR2EMD7v7Iv9/uf3
kwuYRA27KNljUhen5iC4z9AhSUncUdjg63/qERtpjIjDi9lx2nEYBtTUg7ri0n/RLHZDse8xXigp
IfEyynjYLOW88k1B+Wz2zjBQS8tmrrNAlxCSeMQJOYaeKkVSF7lFgeB3J4v4/u/Z7FaYE79WGIhd
f5hc/wdG3TuQt0sl34h5PZeQQ+bOSUz/tj3q5JGcbRzS7tFqlW3ZwB8RRTmrPtPIoG46oV4ic9AJ
wZFrGQ8s1e1GeNDZ2ZV5+RRg2MTXssEIBDqGv8rt2oavaOhT2wTZYB6P2MZHCysBitWOWjRebPH2
gK5U5tUfXK/I0kV2JBf+SBqeHG+uoRqWWXzdPin7UJxq7FpnSBX2ih66cDsrE53xqTO7mHcIuQds
vI+KriNtEn2YVnXh0gZVy1Oi/zBVkrBzw2KNU8fS91UIXum8loxNFK7L5jJ3PS7vn7SsshRtIYLM
EJn3Qb+bqbTqOvLETQqY07h8QiXZfvQ8X1H3cTxQo2rYTej4ZRzEVo2oSTQxRm0UsH10tchi/PWY
lF0vrtC0a+qzGIL3p/rDQMVfMNJtSPhRTzlX/KKjx5/SBE0uz3iHmC5+FhW+WqTWXb7eHqBmo5vq
1oPMDApQh55l1ahS1TsMpKd4F8gCxwzlsF35W7SxivBhZRCvQYHYP4iEvKSEitdVfXxHROHhuUF8
Kuk3j+8luCnhnEiDEE+5q3U+T9VODI7j37Wr2Z0YpHFFOrsfHqUPAkhxv2zhxlB++VieTlcp+qr8
oDv6bEDjyk0NwpEEoWQi+LzpuLoRKoqfQ7miDv4VuPdlxT52uYz+YZF4TBVMXAPRBY2nmfhi8ddu
XNlGF1HzOq5ThVjr9j/5jQ8EumxBBUpSZM2BAs17GxWalruF6nIksOG1HEHdfb5rbwSzc+ANvOe2
5CM7os1lBIBduMMbVKLRITFSSCIT/lgT8kw81cwSpmTghldhakbAK2e7Sr2hxVMwEmcnsU+BjU58
z6K/rRoYkyZYj5BCEPoYIvITevbzpzVgxIcMtnV31b0WuDzQ1ppNpyJKpOvK9pxZcBXdXhJKRy43
pMbZbUAMVCMOOpuPLg6gjkWdeldq0Q8ZE7/QMK35tIMHFoogBIFlTpYQBEpw23j9hm9I9qEUGDbd
d4lolXJ8djqWpfWClHxjlR24ZefjwRGDH9zxuor3JtCIv800gNp5sgGa5f4mjyxkEVmH35eUWJeh
R2TKde2ZmwUdPS/UuJTVpJTbA50rVEiPp7TE38ElskAmRvhnQ1TdGpWZd3+PUtzWZb/Iw4XRBDwK
0kUl8IxIcehz+PHMNxwH6F+SCU9zo49MWdLCAarDJq/2QqtT1p3dVq8BOeMwjoAj/VLfztkH4rk5
D6Or9zZVVqmzZzuB8YEb/6fn4EoCvSpemBScDPWpQ32oMhELpTVRa6nRYRyPAxfEF/1D6qx3VIqu
Ebz5B4MGdUs1GGY0ahoEK76q/p9Ir493X0f4WrV1pfDXxpTcKN8in7TlLrrgxxavqiYyQmlLoeDw
7qR4rzn+ZYlw6aPFaoszagb0x848Tb1AhcsWiqYxV0a6BKqLC+oO98MLbI3tM8jq9QpTpdBMAXto
Li3L3mXtshsHlDkGiI376G0ajBpx5BqfvymZRzMJE3bSAqedT0euPU8muSRX+PzhMlFtkr8FbegX
lj4SggK7tYb9L3L1ZfTiRChmAFWNbVWWrIV2W0gJ+dmQneYpBB07M2w/9162AwkKRwXNcJfLbHD+
+Q3KqVCi/xvkHsvuYgfskhxAkl0VbVU14P7jdxMFRsUPF+LoWElec2aLr7vWpi4o311DleZ4T0ML
z/bhBlhqQn1Y6RgEYKCoJn1Wfn62jSTueeXCMWSSZPPBNP7Bzbw/g+vLzQ1Sty2iSvqohV4As7DU
kgToV7exou7VFOs89nYXiIS4rodlAwBIJWRCI64ZJZJQqPFtQhZumOaDQ3RIVoKHPqJWhRy3PHUs
PcTIMM9gTitGKz09tPo7IydWbhjiU+JQHiJwi5CVy19jAjCC16WP92LNdzpY9NyMSE18OqRs/e8N
0f03/IIrgxoRIJCUVmguRvJVvGWtxp4E0pneFKCqDzrZ7nz3z3lwie+Xkd73GcZDQdBha+bRuIaH
jza/H4NWIgtSLGFfYVSK6NxkF/Ky/L+WM2P/O85s4oxeT7UkSRVnunE2rGtw6v6EThSjyDj0edCJ
pMSH7ykJD5A8qy2umf2YALiRP9J+rM1uBx6/s3irT6dsE3Lfug6arDBxWFu67oYdL3u/AEzfrxCm
FM2SnTYQpLUvHS4wDy+6ElkB8opYVjqb37/2b39jc1QOoHGJw8dgdic3PY+nwaz0EyYn5VevYyLg
qf1y6cvhPkGS+2fy/42I9BqN5yL3HrohVb8iX//negHamqECu7wxvcvYaAzH/l+rxZ/2V+Qr1cm7
wTFmrZ6qb2e3nRhk3eREMhRm4R7qV9fTdVqkQhnvlY6T6zQyap4fikFiD5hsurJgtrbnV41ods8i
zc+S19V9TvxEl0dOXfQ/DwTd2+wgL3K4pVbEcojwIeZNy3J2DhkWmw/HxCcgJAex7xlsmNrGexD1
Vc3o98rpMcfxLNLVEw6C/nyndSxij6UYFEEYG1kizd+P1lfIf+atsfKo9egBNTWxn8QRYmGWoR2Q
2KS+PcploSpo8JI4VeqTirjkFnqoY02FsxsYH1yNdspKEpvrr+9DMCwD+DBJqr9SG0JcBz7h7H3l
tyPfKjVJmgtT3HZ3aOmCr9IZ3aWx059ME07fVo3LF2/yaWFdOkwFcMRo3gvtXLMz8FGXLna9nBsy
KqLhZlDa1kOgvDRk96yMTM/iKI8OzPuhK3cCojaCpTvaS4aFcVpuyyjdsz9r8NRypDFFCyomuc82
H6U7cMVe//ULZBKOlZhH1yUjnGXNKn4IRHK2m2lhL4LENMVs6qIdheEJKSiStzu5hBMQjXjC75j5
fLBWFw++X/AaLl33KBeBgeC+XMUTrRJxVVtqfO0iD1a2uglLHxwk12JQOUPGfLUJey5Q3r9frlKi
6cKV/g/Vv9znF1nZr0ZCM251b4EJFrGtjCla0p3ScJCpRzEoejDFircBsayAMRvaahAgnvCmSfEO
WnmIA6jvHrmi+dJvKOi+PJiS87+XKcehgTw+bvO3itT9nda/mqkgKK2ITgnYMN5WEbhgSzS5rMFV
LK559x8g82BGpfk7el60HwX8DhqfNI71WFoMpd+0KwZhRTn5X0lWtnps/o2JESZ0jbVKLnf/TVyO
u1oRK1WNuInQb5SucScq9BHcnVnmkewdT/84TgWYekLYlxpCzbIchiMbuCJCYRnIGkToNJt1F67m
Es0pjlWU2OnaRRWizy1h9q4Z0vvgjY34YoTlXMCAa+H73/xFX/q+x3/hziGbhKPYjxpx5JBY3u3v
2TJhDSnxruK3CyQlNyJYchC/JPZ773VYwjMDK5xp3PgPoLpystKtY7sS/K1nWDFd8bg9SUu1Uetv
bk6H6nn8x4Ycjqa7lSVuhfO6CXICpgrDbr0Nd6QnT+dbf9DJb1oYwqQBBtzt9vazQYPjveGB8PU3
/r4sDTCNpjkDQ4NGnYTtcaB9cDgJMZtdlYjY+JHj/7rHo+UnDi32XMQjrnLN6lxU5OypFbnCBy1u
xfeme819FPCEMfAK6JocTIXD/jVuvrurfttKmcuo3+oPp74AiVkXa01NICu/4f8Xf1c01UFYEjmz
/3MuYyuh4cTHEm5p391eiTepuag/JdW9NRKUlQaJJavYJmqjRoqjX11Od4pbcriVldSrpW5R/cr3
rc5aS7ZVkWsB4PaLGJkoufySzmJKdK6Hl9RKpZgZ/14c0L55YJ36u6e6prvxXjhfb9w1I6CqzTNJ
Bt6GK748LFYx3FN+F3qgA5BZ7U50JR5Gf5L1q29duI5AW3arAkvXWf6wK0+LzvcAkV+wUxy2LPZu
3cCRPU0WR/OgFefZWgOB8LFoqXtyDxjFHZxk/Bqew4DnM0XzsWyxVUYjun8MqNPCaSNix0afHy4Y
mzlzhwLsTJ/RvCeebGg9bayJVGepzM71lEB657lTgAWNi5x8CiOTAXMYZGxcOyPSpJqrQJgeALqT
Xlm0sAxABufBnBCCduZ95D0e8Ioo8/TphLSFm/C0xu8TghdkLHvqW9lIpQiNZ/UCmwaahq/Izv4H
NMMjs1zxMVQFl/DD2PeCz0Sjkp+N3k2ys81nHQa+xrXAb1ZwIm6DJgl7MNvT8IFXUA0Mq+knIMin
duycmEbjlOxsjE1BbXpYskMdZP81zSddZ3QBP2uH/dxSOhFo/m8MjO0O4rKEZZHN5MoAHL8FSjD0
pQuMG69HBaQS1ovHsECV8EailrQ7e2Dx+DA7g8nZOJLN8YyuqlFBpJVTdR7eLIj98XvR0yu3BXbo
8f5Uj4mFsfKaLnl8CcvpzNDqpt2YPmdnFkhbQT/PTKjUAimQlCG1jYernNX9ff78fqzLpc72q2Wd
5XiF29t0q0dNzg2RE5AHYmIYTSWLxvAOWqC8dqFFVzp0IpqeNPeutwVeqg7v2cGEl8JdgA9izu98
wdzl9D68vgJHzSMdq6ln/KBfK4e71WYjyvQ8tM5Vpbr4SfOVS2GnlBDzIk4PYsN7CiMrMW11+wK1
sG8ewD/ae803pCG5cvSxr4bkWUurvAYsgV/ddWc1vRJ9EvTjeYJv3FP0han1y13yh2A0V6BxmCt/
+vVKqWvj6ZHu/+MxTwmDgKNSoWuW2wz+Udky/YNZUqB9/ZZXBe99TJM7tzVBDAKoyCUXQIwLCSJP
IKIGKUFKbpRTrcq7XlsqnuAJ8rb0uAqCl9xuWMZu6tQMJPgrb+AOH3nsreD+V+3t/b2bGX93MzE9
ac8Dw5vWk/4xV0w1SyKXadBxqoDYwApKwDChOY9GJYDENuZHLbVGmA0X9iOSXyEXmynYrkRbukM2
qivlfTe5otv+yGcEjnSSQZeZE0zRABzz0TWcnTxdApvqCpWflHv724J214I5j00bjKdPzDKWv0v6
51NPjvmil6XJktKmsNXQ2s0AQ61Vf2nNCa6LW5fGs/lwKd3R9Uyf3E8GebDUDYDhPduyyC2VuQwd
CcSkPZ09UQyLV5zMey1sP74g/OnaeAaQMq6VESCfygkZkkuifMHG5hXkKuHAgGZHsuowpu7rnwmQ
sMDRi4o1GImzH61w1/XL+v2TZk0n9jrrNcJmAWOY17osIfk+1SLmqaMvO2+nhW6YzvTi5vmC8RKs
B3+ziUckaBDWGD6iUz3oYAtwG0a4/M788mHVpCNnyp1znXw2JzQ4A3pSlt+nnWkm1QrpQqu6shwO
zioccl64uZI4edoeD0yuZvURzNyo9CzzsetIAGdUug168iIrTH2p2ojXKhcMEJDhFSwssALCeZ5u
ZUqpubWZsVl3PJWd2sq/3WvAq+9q/PUDCvSFd8BSy/SO5lF6z1q6TIz+b4zp1kJHWP8PzTaegB9T
UoVfGwAUD7+hOEGmvOUCgqXn77WW9Ve19jTPQY5SC5n9Y3l/Y7zI37/1lOhrOSIOwMykH/ZHfQpK
FtYKMhjhcKg9CqnRGZNWiT0dmWhnCTgHkfVw+G+lt6a/tHl8yRYQSbpVqLomKoX74e2Kj8tV+2c/
U1AHY6JITFbD8vixHM7GoXvGaYGvNxJeOXI8E9jTM0NKd2hx+m1YmJXPPo95P0UI+z/eTw2ecnYZ
1Mhe3jzmURy/nxRtue1tE4lWvVyJn9ToSDjv52VuzVGslsoouOjPLZELyE8fgXnabqTsfEQkwMwP
9t9mc4CaY98DFWwvMY0DnvvwIEhS52sLiBw6S44KgR6V/PLMwhtdsK0Tu4Ia03ppYkyG2KyWKtCP
etBi/OBiSLUHlClCQuOvSGWtcvx0PK3BsET2+KPsxu34hizLi3ewkDFTIl/m2NGmcHTcnzaCcWeT
gCXUTRwe7Macd+JIdp5qALe4unkeZLKOVOD/BcI/jJvBF9R9LUUDHoterDg78Y1jWyMteExEBp84
Xri2cpX99fAyjHalC8RMfwJHewxp3badIpbpFNxmgA3ElzWiO/QWpkXDlgSqnqFpoL/UJC3QWApa
yUHGzK5OVQV6PSeUDZ2IRgZ2dSvzexe5rS15tLIaqXB3asvT+OT1ib+eUcWgYcgGj0lHzBwwTXdh
NWXvaANHTLxoOTFhKp5OdIfdjDO7vQHdSuMFkw37sLnUzoReQGGm7trosFKqTcgubuXRMp6W+264
gELwbF8ondc/7T1vPiFwQgE5I+XfzwzGveRQLejC9VAIjSbwUeDVsyCnD+JGAcvuscWDV2hqvSh/
hx9lnA1dLJp166Sby2ubPcPFajjQe1AE4Wxln33FF1SQFtBZB1k5lcGMspUhbiDhcI5Yhblc6U1b
/sGyPPjeEI+0JMtsompfoGnOAMny8RidrUOhFqob6s60hQCq4Z0ZGC23y+Bph4xY6kTzhuOX14KX
RJ8MZidTaRbIC61tr64AIrg1BhCwKIk5i7s82jwey0WYS1bno8zBkc98VZM0Z7wua2IzGW5Jt77K
20YJoa3zFlvJlqagcCHzTAlgQANtkAii/cQP4h3LJOX01n98GVXUvG9DzE7pcHvUn+7qwnRkazd/
jvor7sEa6+OhUkZMFAOw/fNv1ZeoC8IXSXeiAwMbQQo4tAio1DT2KiPiBF9/+txFH1WyLhWIu6Gb
ydcmsluV20sGHXgoYWN48kdP/W/aeWC0fq0OMKPEjuQjGajc/9r75ZEqg4ZHQ2Wsx0V18QibkYx4
uEYf93xso87gRSBJUpXlHvoRlW9XQbPaUn8f/wM3EdLWkugKuZqpzvxlvBe//J5g8A76mw2Pjrf6
bZZKsGie9/kI0dQjM2OATAcSaOohyAZd3iJtMhWpUUQZxreB2cighOHKiDIjidNKxoc4/8YD0aho
WZa6qeTjyQH+2lKyJRZ36bZFTGWhJK3JYG8keCy4of1FJBRpWLHyZgL+Jg0oCfmf6zh4GBdYLsLv
vv1/OjtsYJtmfLS7+++xVnhyMoTPdBMZdPMiUsT26uBB/w7ev56Uo9y5DtWVoZyzFWHpBrmeIQBh
MU+TZRN6J9I8j6h3kYArOw+3o806YsBE8FgRG9FrwPzqqkaJ4myiAFkL0Q0jSWAKcFgTO2hiCN0p
TbCdH1qetW+Dheh6pnhuDNzZkqx50N+xjHqw6WV368V4mqetOc7gYeNuj51n1ayLu51w3Y0xA1YH
qQSHz2vVqjcGPfP1ittnZcO6+z5DpGuqCF1OM4+/nt5vOZ7yFrU6QDXtcsF2g01dGh+2mzRNS5Bx
MDp2VvIJXqS+dV6qqupENZo5RItVVIxdRn+KAM8kAKug/0YB2Dgoo9qB0apXlbADbLlVEzim9m7G
AH8dRCogfJ2Z0/xbddGoBGU2W6Qew0pcCfmu4P05Q7AnjAoijsAwLkce5vDixwsntHc1xOc8yEnj
9tI75jZ/3RvE2lsBSSPdtGgoBhiASEhdj1IMpzkt3itiE9+zMW8QaaDmPciyzBmAQo8Fd5tQkwvu
VmuVD0vMsNfizOXW2RiDH5ZhrbwHS1WwnPbjdUuNvTiakDqbBllWrGN+vPlGXkiX700H96BBOdnZ
d6uzh/k5hYQHaBHFOTnWRFzHhp9SYdHaO7YZ0VBXTYi5axNnpQrCE+c/HWX+/eLX/4s0acShWFAZ
IZjZK9UQRB+4oqHRDqTgMLd5UUkte8sYldeRTz/EgHVOGol1U9e10wMBeLcR95SZ1OBJA7ru5O0E
lIhuICeALE3FcIIrQSte+ndGVIfvZH9iqjfj6aV8BlggjZWq/AUeilSgEoh9N6/Bd+LOmmLAJRGY
ghbT3B0ay2VHvEttNZ1H4WVmoWd7OUh8O6P+XJ6LpkkQ7IsS8Wzrc85b2me8uSiDyzvmGA5evbHN
godTxItRFXmOmgQns5DW4co5oK+SSH4TxENihqI9MRLl6/9z3bD1AQhM4aXEClgxyC/iDHUHxZMv
pnV7xm55AZE+oNB2Y3IVxLM1SzT9nMYHqL6vBnOKz1fGtuE/R34gDNwYDa1gUWb0DnP/qjLAN5YZ
cLvTXvoC9PkbPJEIvd8VR40CmV1ifGVTw1QeiUur3oRdoh/h/X7PPrcS20Ume5OmChdKNPpewbPr
kIxr9CZvwhZ1CVWrUYbL6S7a9iXr5/sSQQX0s+MtSSiATx0rdSGxGgcr2dQbWkGvmJEwSZvn39rL
KwjQVMwSkTxL7TyqbR554NYJ55UGJfEeimNBdc2/p932ju+J9YQ+EG7g4w2lBhAIQhrd4ykrEhYh
rojdtQ3gtA/K35NlDSAfZzmDnIN+TPyZX2nlPCmOQucdipgzWOs0fc1IOx5rv1qshpvUendRa2rh
yoMs8pO5CeNudT6WFBz2u0q2exJrlDbmOZHQdg13lvgQU23ue9jObZ8v838OAALqf9XL3C9G+rud
qVhDFPMF6hNOI3TjR723vbdANrL/2mXVuwr785WPW5/qsPFMhltYs7tdXckPZgxWa8PAL1rMt7q5
WZkKqf3WfOHRovrmJ795mhQqgGjGLVkSmES5QY7X7aImA3Yo18yhSUKbpVv7Hcebbvn66c+GQUdw
MQnybO9+S/DM3H5/W6J4HI4H5h3AdnZ0S1APnT3f3bqOJAIcaWUVCjBGiJTrjdnorTosK2truT10
hm7N5oP0tvbnu3HF7qLZzMKCAynmO2jOrU2Nb6+hHziRnr0lFk2hBPfgT6NjXW53fDv+mt6g3q58
rJS0Hg7rk48Xy9BwVhK6g2F6sVBko01qTIyZUre6pAgV5gQO9XXZH04hill+Z1WFZCWAEMsUsxhF
/xaDaT7oRAmMTK1b6K8vAjPfeyBfFfKKGhuNM+BZ3EueR8ICwzei7LUPUOzeZcHQkROWEjWB5AFC
sxQC+r3HWD1A1CCua90FBfSChudR/238emUE+jpEvQjp2O38zYpNYhmMaf8QysUhXgZy9DKGQ2Oj
HEZBQKvqluyDC4mcFVNKcCCal2kG2Sd+QzgLX/27zg+rilutxT125RdE45/Rd7TGn0/2dVseRfGn
g87kzqztLjIlI0Qst4mPD8Y/5E4jTyeDcOsfKP+zGNi89th4PAATGRzfn7QzMPPFLNWwCeyo6ICa
qtxBeK25LKYowgbqYuKsxA139ZuyEozCrAQmdecbJwpkhkgT6hH0hv4E6dKJWD+6arLhudqrjPML
B4RCVL416sdC9sN2w0+t2PQFCF95Fa98zwbcQ0YrDEh89bwuARdlMGe8oKpBmVAttAPVM4rZG8wE
WIIj+AI6IbT2iS8I1IvJDTlw0x73E0GPOYJlXVMbg/jLfA+/P6H3LuB1Lw0LppdewEeUH+Jswf0n
dkNE5Xu8veAXeQkbFiC4OXIs+S+CNcc54TOZUp0QLyKfVeyEWDpSqnNTy1K5bEocCKojS9OoOkir
Gaa2x8qcpNhGbs7JPnRXUjOZ2grzVI44E8QqK9u6Pjga8/GBLajr3gszMhoGPK2zzdc7Otwo1ETV
p+C/dVPH1hRvNq3PiaHmY48RZU5+WTC1NQiAgGacLlUh/h6NaZjj/veST7JgJ0cdPdGj/E7nusfp
OSHrSkx9Px3NpMYcf23L51jMn3FwXDCFZn5Spg6NvdT19VJKLpxGT2cFfS9yZPiCCBX4pDTSjjGk
wKIP0hZVNozCZDr0OmyFHtZM7LqwaONXKnCqa8Fa/uho63tCLZd5UNKZRs6flXTh9ses4ZtHO15g
LlUZjrrY0dwrxbDjXGpN9LKnP+571EKweTzKsLx7uEyTBfEoObq+Exydvtj/AaTBTl+/PZ6XQJcq
f/IEDA0mEmZG6/0ayF2M2iCbqXvBSbyeqTQP+7kqpGE7IWft6fB9oHF3v1upP9uTqNrE1PECRJtR
U+s7hW0+hgexDrs32KtFnEkFI9V99Fn1N5FAKzyxZ0iA+bN0E9FZclcVHwVtcjwHb4cxqOqUkgb4
+22kXERCnswwX5SyOIkA3zqZfO2VJ/pImO9pVaHO9P2aH0B5G3fDe2N1H3BgsW7uOj4CKKc1ojIU
RDDY/lG+ZDXJKDPkFfjCpQdHWGqtaSR65IV8CMhDIkOCieRUdOZulz4XvSXmPrw3g1SS1RvkFXup
iUB9+eSVU5wjT+Z8n0BEtJWKmr5tLqKLcpjzt1JWzrQLCJg996VdFjRNim2juGoqbdB+CH2nuN1W
98uTMEvKxZswCQiAV67p+cTeVHlIP0hEr09mS+4ySHLtG3oe0nHscOUwz6MREmOJKmFBZXO/CqwH
ViYNXfSdSYCyNtVs+y/Bs98YEExSm0rvJljai1Om7xFvbnPKCrn/+kOPQEHkw/XXCE06a2SRcmxS
O39JOeWUJsF3G8yNF56iSOp7A47EqrzxQT/nK91FQAqoWRN9KDt98vO8wUhcgpRoWXKBLVCy3eDr
vj3MiaM+duMo4G+iTdvqFAIQC90BgW7qZDMM+XUZKjBZamPVuKGDbz9+ld5ffHjAnSdZTCGa5Tvh
ihMFhXMPc1SojvV8QKqRxeKVeC5C9siMWZWb30EEB6xYqxVumh2N/eWnj7XWUOrMOKB0uIN0eIT2
kmigtoLOY4tXPppX6ngKDaKKOiquDVRkTlpr6pwYP142nhR2sOBmpuSNo1N9rlryGLlVGHlfKGpv
5+iWdzz+H0uIR98gDKSvkJbb2vxBroqdRU5/Z1Jqv0vafLJOM7ImIppi+trX+MCCUAXWWrQi7tHr
/enmew7FF1hRcsWoP5w77rjY+peNcl66/w6CYhUxJuXjRTnitvTxz1WssstdF1+wt1Tvmsn2hgXY
LQgoMS69BqmEYo3vqgq2cShhzkV358tUx6FK+GygYwx/qyE4y2UPcybBYIZWm6c6xOklm3UpMEdd
WyWf18W7fLZShpHiGell0uKm6raZ0SuMtDmFQCqeyXileXjSbG6iLXcm7Yi9OAwdReXUhWKFLlz9
eV56ahiIh43DKNGJV8Ivit4qjSAR6wvy+Vwgb+gm1OFpzKL3ay1aphpAKmeeul+z6ThEhZ8HM0y7
4XSu8okBniTKsZuREH8O65rLlPYgpwdGTPeUfrFaWnQ3gkMG4KwoFfj6OcOgBnoAaoRFzKkRM2rA
9Tw2s6c9NIuQxSzJxX4BCfvW9p0lwlAnck7ytX09pm4zYMhcgjjimYGBtujBuKXKfEG1nRGb7ZQ5
PU/SxbGToGvTeznk1jorRAnEl2PsP8LKqUYw9L+iXQz1jCSyXDnwDdITi0JXwR/tJ/DZUQZwvxMp
bepSA5dFzkGfAK26uSZNY/gFAbwIY3IthVrareYCpyF63UiqJKhqDcZwG5vHZUL1DhRQP/Yy/9CK
Ud9FZmwCWdeX0g0+JBW7jt2tW5VfRCB1wl4Sipc+HZb0TWyzMIAaut9z62NiuKCglL3sVFDscHb9
Z7LvkL3eNNXQVK40nqxLs9TKCcTKBsfVF2geigcCZ2EJrSPhL51dAPqk2ceX0hcyOuF2HxRuPZbo
c2xLpVp++OajB56W27r4xsqqZvygS/b8WoSzMcGOmRFDfEHtJf64gTzBUNZdA5f5vrU3VcZ6x89n
ZFp/f0Hgki7qn97nKNhfdWXjQUXvdnq42XJS1hTslXY6587TvBuhCfLPdkIu/z6z+Lf6wusAhCS9
NoTNzm/5YxW2wwI3pIoJ3Fp74qXnN32LpwCxYg6HltX5m7ZFXaY+yKdTDf4t+USzsj85aavhxWxU
N2/EiBxWWH8K/9lFZ3tkIRnWv7b8Pj/kV3UK5JvruB+ZbyQIndM1TPKLncNzLgSbNoSrfn2CudhK
O/SBMM9BRWuO47rpFnCx4lWa9CDZYHX3fNOM8RR8jIhWREGKrCoyy4k5u7gR0qSrWmMrI2x/JweI
EZuIdMwrfKTsgKHc4655eirfptNSIgMr8H7wqkD/mxEPEhdEMtE9B/rgMvstrPwlEP3sR7LWOcUR
4YJCoX5ptk7CBzFW8HJgHDhPvqeceAi0D46LVmvVfUk32r4078H6XtENSxACOpHSxTFs/wuC8VgJ
wDkNhI2seWNJmrRPYK1nh5teCabvcLwcYdwCcpyM4f7FQGz8pTvmGE5GZ0oT2ccQPFYzfcs5wY67
rKq1Nx5yPXO4/q+Pyfy4lsGzvjN0Y2zgRLw4sflqdaTL1ewpkEw8K9o2v7B6bNMfQWEnTddnuc62
9GFnQC2zP6aGUSA3+wMHofcggiG4kOlj1QG/zSUvxvH11fVEE9VeJWrbvqqt++goS6xXxObCXMpr
mFdEiErY2FjfVskVEse70SeaC2xdUS6qeda4qt1i7u0B/GLQK6blupB6jupsditNTFXuddkmVO5Y
oHytAbduJ7APvgcu1t//gRuX+sn+OGd/R/HFmaILqvq7sQVzjGllxld71Czg9nb8QMFrvhNWHsYn
UD+MsK4USjy3tvtanfOUaLpMxz0usj0XSc43dK/DHRQP77wAQRgRKK6NreTvrM5fpX8Kt3GCfdDr
bH+B3hvd4isWJy6vOKCpBcjRWdT9m9PfnVlQKhVHp06ae3dmCnDQYUoUvXGbeeYSAuU6FzZGByHj
22ip7+N6Mvmytex74/y0IgJb8pCIITNvWFor6UAN31vDTHX6joI754r8YDp6Ae1PZFXuKnaQCum+
d7wn9joCSklUnTjcYXMpVNdWpAtghaIQlLawiZ7dhpkpVIdC330OfMRUaaSXFZX8mljH94BgrtzS
oKFXkyiGGj8QlLUuUV2AzZBh0q4Zs8mcpfontWIdrTyMZY5HLrl70PnNGipCnLajJ0JKZepGqORr
43R1p4MTrTdazapFUCuG10Ry2b1d2yGD7eDxZam5QTQ7PqzMkk6Uu/69g502QX0dy21/GLO8+1zh
oAZOR5Zjbc73GYMSVxafOMt6nkcbyWELp/r7bSWsmnDYmJHDhswHrMkU03apgmkKFIqzXPYaZ6W6
MpGlwOcWcdr6dxJSVevmZQfM3oH/CkLoZhq6XiEeqj1bK4Ojo1fRYRb6e01qWI6ymnZVPBons70I
gV6M0Fst6zY5Uk8N/hbUU+HRjE51pR1GijGaV0kNkXk44zMmcYFA9q7btFvWHZgkaBuDm5r5c0Lt
6PrIvVFwc2UE1wtJx2EnEw9nTajQdJ3aH5uu2+QR4IiCdlf4+AubHQvR0Y0MiGZmhXI0IqZHRjqq
JJDl2mfg5NcYFc/xH576R0mlyP4HuWy0eDt9TcqulD2WZhIWO1BcRbsl7+Igw3Ko8VCuEeAqr3oF
f7U2dwq6l8f6FVALKWI35OVGINYrLwWMwyseWtHJVXXKkZV6HoUcbpqI8PaXDw5yZyumowxPb8jl
W+75LX2hiY8FdAFwjfKuFonsGK+aWTIUsP+KaW6IMyzly+7GVsMDJqH9NiBwmcVBpnexT/UAc8Ix
a8M9Vzbm8HIWYa+eEomqlQW40A6Zh7pdcevh+Ux8nd2NZ+sLVMOlTwjrRjZUfz1tWY4xqLrKG6JG
IGyGi9b3+qdhSWD0M5ogTgFFoTO5oXJX4aNASPKTbwbyJCIco1U4x7Us8xnjuBxvZIpYQAtBx3MZ
dumAsnyKD3tUQk3SdHlp3ZztiY+UBI1J85ijecLp73s0PpiBnuna0SywQ7KdTPfB8ib7JhGMBla2
pvQ1HmbLcxg1Gz9hdh71veJYI9CxCYrsP0XPI4YqWcKeTf2RNGkgiE4X6zYaz8bYqxZ400tg53AS
xMnRkJcMO8GHDtrre8g5UlSH2X22fpH0p/qh6sLVY/L4EoRfE4bH1jf+cZp0ZdH4Pfs6M4fPnUs2
h2ufPOCDWiXajR3LgyguLtlIVhqgUZiruyyNduxMHTIK61gjA8/wAX/g1f+xrZIoy/H+QAQjjVdY
HDWv/lR/kiWDDxoi786SI8n96iVN2mpsC78AdPeGVHmAPgHeVFhm6Gc6hxeG8vl4nwWbzx2Q9NtC
BNkVam7J6WHbcgJ9apQORE4YTDzPBtNK42qxAXb/WRcl4bYwgMqGlEQ9wLFw6QHqR4hR/Nk3DFUM
IeVtCpicdxkZK6hTrtzYmk+tZD6ijpatS27EpQyChhPzkWpjZT8f4BnQG36NmKtAmJ8CFsTXAbcJ
iAR1L9khum3XNJqagqj/Z2YaNny0izVVTQ1zJMz/kpIPoc//ZBgscXEUwqPha7aWfQ+b1lDHpYlt
n3PSr1YusNGWFUPexdxnTh02u/vP73ydvEM8knOVkGBX6S+hxOi/CkvdwX+VITS+binOpa5esxvi
I9aLOjTF0jQDw16gPQXup5zBRU9D1/QS94gkzufRXWlSuZa+t4UQAj3weMM8y1vKQWYzgBLvECF9
RizUYk9SFpnhi43UOHcFJTPnKvZuiasbZ05tz6+SFK1rFhZfJFL9vgxheMFkLW0H5Zc8sFX2pejd
iAt7/0ayapgIPBr453u9Vfr7/0ZdXTG3gW1gJGIcElnS2GfKKViIkd9OoBBsT8JPhGzPjanv52tM
j7OkQtbwSC3nU7IXWmiAiyza40JBzgPd1/d6w8EG1b5sznQ1WLeLU5u5Whb7hTXF+SvXCQ1fAXq/
MPCyhBXfNe7P4mOdWh1o0UOetpUBNv+sPV/xrIHkQgtDeXiGWIDxEYZDR+ufTCxhfCQtw3DHrp+F
8sff67S6564zKnBgym3Mnh22Tj1eAJEVZXWiHWzaCcpqefR7KojpyVPsTczBPrRJobsMIpYBmOS/
0946fmKuWMvXA+xJCixhjXb63qBzIuY6zV+LYXdqU1CGqwp5k/mVOmwjxutg/6PRq46DeF5egsxQ
5oYqsIInovQhPkjwXyE+4A61uFb+y3YzHjPo+4i+ULc+fTKZJJ/NOpQVsTbsDEfwNVkyoXEbYZOH
nLXkvploKFIvi6bNMneTsDl0AaEz7rNw61w19SRPHAatcI3Wsjw3lTkgAnwOElIGZAkca17MNsoE
cGBFkhCSwi8l2cmr2O/0W2B0d4FH2Z3Kfk9re17xFDPAhBAfTRaMNVDmeOgKDhtXEdR9QG6P4m6E
AuxEcZ6Bhv3gK/ul77HwFRxPeKGf5eW+q1mFudYtxlKa8oOr8ocrUKuD1PgV3veI0EdEY7I1fo+A
sT94eOaIUJqXbjVlF+qvIPfm1nQ/E8LvI2nzOE9R468NFx1j922Q4TtbZD7qleDAPo603pLR3djF
CefAr4t0l9u8GwcM2UAxvO9ad72OzsqlxOv05Eh833DNeU1EtC8B1DaShliuRkBAylWLCPXy4G9D
DsNGUkzqTGqCNOW+vFbcBaTxOaFNEqdnkKTm5LzDw1VoubOIt3T7ZGzP8JPtjrFT7to+zSGMLNQV
XCagY8soP2eOJ7iXmrB87Kemh7t8fevIf71LwQJM2Kks5OFFfNNG0vSMpHLOBRAextJ7PoAxEkl/
/8A3Or0awJv4pd236W2YAPofb0J4BDkd5Jl81guAj3unQViN0IFiONHExQvJySvY/QvdC6Uc5pws
bAmYYj7aKfTU2vacJhVQE7RmujzI594OD6B8I7EqtH5JRujKGesrAjrdobD7G2xNXwjjJW/5MjEu
XA67l2HM1jsQmBPe/GaqHaoSldnYFTunpGJv5yrbLNj06ykYonAQTYmSpOOY5yEt0O0+0c5+LYT+
k+pmP2/nxEtJDvFjXA5l5opc+QAu6p+vcGPGA6Ac2ZJFbNFrFlajWJKAvNMeS6Ak8KQOXGjtyWIy
prvJjAi7ZFgov9f7Ued+yfPzDOarmIp7dBFBoWfwgrb1IC2qK/8Go4IyAYOp0RmwbufmPrDO9aDG
CcAz0ha2Sj6+j4sxXFjoatpamq8imkHQOwVGHbo0heN9n/2RxSwEi00TBNrnY9B8sbhnAOAKxIV9
E7TSIR+AULhVaZYzu9OkKIfyQAikEBXB+X79kCL4Ru4D6pNXDiOPJJ/MqwK3Xxo3CoZexb+BDIgI
cc5a8ATFdCxAmm6mO0Zql3hP9Y0cxMHFHBaSpVattdaw0x/K29EdEs8YegeSmHcQZuch883QTCPR
VOqQMsWfVnQLzyr7+AkafdB6RCSv38959UmcSxpOp1Tm+FcBQxWseNAcaNDr1VIlORuAdu8Hk91q
EiFCECAww6r3hfkuIHXDl17LC1+yP54A6oMT9hxDbZ3QknU983MlYE6sCWYuJLnUhct9CumNan4o
IdQ3s9isRNzxWf7ehDUtbuTcXHpJ5aBR6WmhNyuMfwmfVqTjwM6pgLZntoauFeIEECkxIs2yWkQV
ZNnwkFnkOIm3EBA8/+meMt1D+8+DqKjXB87Nq8dyLjk1zNFayJR694JOlBSWGU+UwbhrhVjZHcWi
Z5ulTBt73oYeKEgIcvZm466noh94E/KfxbsVNgZ+u670yjqK3utlGIomKelboBoMm2QLRxctpO7W
7Xx9Sbb7dcu1MecjaGXXu6IQAmuWQWs+KXa1i2L/Pn0lsv1jdr0IBIwi3leS/HBiI+wSkzmIHB+i
KrlUrho4shIsuY267/pWR2Mbo4kmXUQrJlrSJDFCP4rsGr9T72Cmvd/hTrVdX+qXkcD62WabXC6h
nibKBGhRVNWrJdr1LlevI+QMn/T34TPU/1HRF9DoEjvN3AAJ0LbxRy5e3QPeh6Qh+93bfvZLhipu
6JiYRnBfIVow3bKs+wOsEDu4pqGZgncUaG7XOj6dhowE9SyusZjpVjruoT8IIIcwkZljg5fAm1O1
TFLAQZ4xEg9pVaWf03h3mYZzHDmrpPMdDyttot1XgWFPkNGdDturV2d4d9MLVZiLW0FZQnVeABrS
nqCuWB0VhBP3Okx33Y5VpwSRPOCbotoutGEDxLCgHcS2LF4iKr1ajatnifqhYCblEyVw7AiixIwS
PFjVSZ6YfAcoNvnSgg8rgkMnHo6cS2oCaj0x2jBqlfzDC0h4btcqlraL5RJ1w4nzEu/Y907/xpM/
yKOMxUzl64fso8Ho2OnyQ5k9Ddm2HCbugS6Z4AAx17uiZ10/kzIlnaOdUjjIu4K6B4G+rLuFmZhT
UF49YNQzBsR7NBzU+IMzYSNqbL0rzJD1yi190yF92fIK/cWvZYcYABbVrRW3qC1HsA41JxR5BWYW
p9xmJCWX73fn7lVM8pzO20Qe2d18yonaEdENlOmp+Z0LCBhbGVE3xDwsL2wy1vibpbLHRvgmxkBA
IG1WUUuA8XWQQptTl248i7Ok0I9mUhU65BiX/m4Nvb9ObbxpfotH9GkPsOoGr/jW684XQY4453Nc
Rz4e9fIXc0HZ26qwobCT1KLBLm6Xoibwc029gyuNe6qU15M53Vl/Qqwpjc9Zbz0sgoLOSB8d2LDz
tSvjC+R0G18WvHQOnX0xCtDc3MgX0xtODCsZCcDOFRNahj1+Ht9yNp4va8x8QTZEckCUpOYqvVsi
omJ/ipQvdnEB6fe0I/6gHea0oQxTp9Qy8bX/k2b7sheSbchM4yFdjpA8WRqCA269GnKH93fIKNAO
mUQOEtsyNEH76bYaCb82iiPtx/dtFu8ksiv7ivdDMKb8Iz4Z+JV6ZRLYB+6kkk8b4KQFNFJrh93W
GCSoZhG9Xvdh5HrGf5Km8KRdHuQZX4+7hHjB4PK4iYY6qCzzYG6g9P992skwrXJAqnT/MEWZocQo
nPsV9asD78uaQcCSIeG7v9MnHtSPK6u3MQ5RiUT6H0keqB4BVxRgSIEQsRKNxedf35/ZKl0kAou1
BnitPl0oWOEu7gUEc53O81FbRWNk0aT4+vuXQDDQ7n0E/c5AIxqAOd4NG5kxrxBysu/TtRhlAOol
4Fz0BGbBQl69k0q9f0YblxgQ0wPxYLhvFPtLA7SjX8b/WqWA1MPlvLESn8uuxz+rozb7wThYEP7V
W0EPVKcW2tWl0WADMRgP6GDJ2ApyG8fKcpkFk/5xogvvsBeMKxgxwNrtxKf8WW2b+QfPgcXriMf7
dUzSt5f9QJ4I09gA5kMuQ1fnS0kCilPyJfekMvSkYhKNC192X8LyU2TV0hYFyf8AEKEcIjXrwRnv
1wWlCmZtfRuiwUR41vE/bgumCeOvivuEFX4mcO9rzo10T8VsrbF+svLihpf0kS+Vh0YWTz8c4d6X
GL+aNN+OQKaQ8Gy47LaHwmE1+NCQMbytGoxehQmA3Ww35r2HVVS3d7MJYzi/WfNFfK/NUvFiMiCI
E9fcDefA3P4kzAmYNajONTWUTn93LQ3hk5O73+5CZM9W3dclneE9Rvc/yZ1MgJkV7hISuZ2Y3WqU
v1lgLkWEpD/pZ3JzfSXNeA2yay9i9QlfKZ6QWJaEKFtKQhYBnevDtN8Zbx40GhQ+QmOvI7icGDwX
b52ByIYjhSD0OX2kMbKrHXQ+OQ+uhR7WadJiGyIX5aRbW0gdFSJbrytJaPJQbG0d4WiJbtOjJY25
Pt+v4+DcTtt4nIXHOuc7EWxS3OJNVo8lhmkAiveGGuA/Zxi82LMEJ824JmrYf6MrlyQgOMT+N+r5
wDf18ak2WB/+djoxUX6QaQTk9R9SYZB6Yq/7qwBedXywtSJoYDdXCxO1tJm1n81+7U4eg3XQS3mc
amJ27nuGKnW3EpCUOr/c8Gl8idpM5OnVtL9eNfELx+ico90UjBj4Jd/NalP+4aOoHLWxqBqKxyrt
Rr2poZE6u2VbHGnYfRor+HJXYlBGxTZ/qqxUFqIXMqc4kJVcW+BA7QDPl7zj/Bqe0Vny1VcsGzb/
slfFk5zs+N8uyG0N62nIGE1WCPabEIJy8ZqV9k53y/dX2DI6VEeuFkYDEsNsEKa0AobAq4wLdLT/
W4arYS5Ik2IKTmfC2SyNo/0ZK+JMVpjEyl3eM85uIVyqsdmd4BTOF7y9OIfkCBTDovLHPWOhJzrl
dGxvBu++O0S7kjRz38m83Emny+Fhuof7lps28MQP/WbQiaGcC0+SajIVZaIeqwYMAtB87QqjDW3g
8lHl/0PhZeXAu+X+V+IgHCG1WbeU3fre9ePLkjLdPybjnqY8UngYeOOL6qCp56Dnish5jdWAxztr
Dld0CCt8Yreazds3QVjF/sYexRa9yRFRueh3eOji+4a4qjTyEgfZoVjlZeu702bdEu3mGnLXMbRc
6XlKTuA0TuwQqiFxLhfBiBSKx6zanZWoYcCyTDledNoeqRuoIBtTNeO6clEEJMjUJ3DGi8tuljFx
6p55tY4Cb+yQkgAzWST7d9REcpWIdSR/dFUT8GYImoR5Ptmx9mEAuVnVnmWvRq/u1blQ0uNovtqT
tjv/x4pEUfFMgddrnW8r3tgphIaU67qHp9bv3VOsmBzlbriD54wLYRCsN8au0OhPbWEg/qR2N4Vy
PcJCdwzcTbZnTtyceLJAkJhJowqX0MGpdWSaxL4ZGhIJGfV4qyf2Kv5gkex/Hqn9nSOaF4h9B54H
m8zAYpunWj8GRksYG5XWkFe29+MeZs5HaSBBU2Pma6Xy2gpG2k+0xwZupYyFcc66zvbKkH//L+ZP
VjWbIN7Gns/GDlD97FAGck80LmLJ1HKXQ8gxqThvr9B2CaUva8cw8a0XHQaZJCHnYec8GKaCGnmM
8HBW8b6eoDtVymw3kbnUuQt3Tdhpxq3ejPn8JZCEEg7sVPds+tZFCXW+d9acOowDSyRJDD3+i+90
lXZk/kZkEkAqTumB0Zf7lHdBISAdJ5sKRnmHYoIU7VaORGWSkWnG61zPbmpeO8ekc2rCy6ndq0vp
7K0tNyF9iyl+l1srMsAl+s1QtmDXJxh+Yi070z0FJ+x0RFTEhooAHgDrmrPLrm1aeT07pBXAVoNn
IqkOQxSEzULB/RLjf0K/4hgPPl158ITpjV5a6EwWFdmyJQKFBOGjHlLglv7f1GoCgZJ3popAI+k0
Y4KMxeXGtS1jyS5JxvetrYGMmH+DxiulmhQh5fr8sXIQ8ByK8QPgz9ghR2XobXzp+OFOpLDlAZIg
Bbrcmw8ouLhAbJ2uWFIspogETeXqPsg+IcdI2yJHnx4aTV2p5N9w0jbwpC/DJ1rWm5ymWFB//s7x
Xh4TEMZqUQpYL3Qtx6F9CY0b2g3qR6JPtkeBpS7cJ34t0FW6JxFDp0ZT8xKhzgWQWExglGtgbwyZ
FrYt26fNrv/Gnlo2JaehTRQQhf6oCDJuOZpo0M0MtfViRLzwmihXHWCP3r6MMJjogrDqh3L9TEVH
SoAWr+AOw9sO8oOaOaFazjtkYAHL/fS2+JpvMNEawuuNLm0uofC4O6fkKSNeQzuH2Q1xn4PcgEdJ
iFhgZPxIwhEaluVOK6XtT0zMwpcmycL9UhRejIifqsyTFPkuWrHoCQUR1kyziTUPd0crX5UXQgIA
WUxzfS20acEV32US8e9VMrpR6t1hayz48qfYyRZHHl+RI2QbnRuJVnxU5UKB+oAtlzQ8cnEgyQIV
sSjJxHJfMsmeKD+Opm9Mq6vqH21XrYmJa3u6ZyZkvJIzGLuhElXOHrX+IWSdyqVa0rlyacxqwBIi
+ZbzHR9qm9/F61Nut0Bv903t32Da3paZTTUfvocAYduknExcG/KQMltolH/iX+50N/fqJLr/2Brm
edWdKhKhSESQrkQK/73Q3pPbs9JWLQaMmzo/rleF1WaET5FrZzEsfvz8nA5csChsoLXx5RkW0wmc
mD3+qxm0ulGfeHYLpbQ6jYqjSUSVo1Po23tSuHMbmiwha1I/fLk36EPQXtfA9IN/uT1xcwGA21Ki
oVSL5lrw6/X+sNZWceq5CSoc4wTDAcciqupJWIczB+cBw3M5GvmUJMYtwZbGv+vg1t98DXgd69Xd
rCirNKrJZKUgdwaB4vh2osL2hBwx9Ekz4y/W2r/CHaq88uW76+yeNjc347LmERzwWysZsLptGc/D
xkD1AL4h53yuMkz9dA7TgTk1TcfYE6wy2w+78j/cRF4EOUeLpIYGVOXQwkIYhjMeptfcbB8lSR/G
seJIh0PT2nI6F3t9Fev/NmdGk26ampt3oU/zByTG2wj0zPfNFEoo0o74xhkVwD6DzrK3k2QlzHCr
/fSTdYD3pScBN1fH3XMB+OpQ/v1G830A2XBJir8nG3qYxNEfbTYPm3fFD8m6USxpQlWbFUzMuSKj
uLY09epWtsgDqeBl31bB4UQUE9EOqANgTLdlb/zDB2og/EfQfohHxEHds1atBO5IG4PEsXTxXel7
vMAX9Xb9Ud2yl6q05NSA+MsFG6Xxr8tK6IjaD93nb0N/EyhSYvZUp0iaeJwxsCx6A+YGqwdyyche
W0YJzeEMJm5nRJGAIeRWbiM8Cvhk7BYtbTravZqsFJCqaefK3CeMVKBiGIAsQytxTT/TdyNWAvhr
jt3cC8VHDFMwRnrdqmR06OhdpIO4kdg6960sNS/2GJgOvhUOLlZhoCg/GoKvt/hvqlzZBSavuVN/
9mkJ2O7As1RwWIRP7GVirpJD9NrX8o0kVtZDRt4UeiVoxBnKmzXmMoLo65oUAKRzMSrsGoa8e+WV
yCsNVDiHPuc7eJ2bn7GrATJP3jnQa2HLzqplUTuI2jNP+/IvnlgGKB89VsqzJmtDO/lyo178Twty
4ReRJUawBKDITkR2bVRv/6bGaIz057MCHkbPS16pc5bXfjRApi009xIBLCjYWeu5HGhuj4fwqLQL
UfyLHyrD5JrAsy3iA4DWc7CwxVHKuA0MKyUx95JcfIV3ps0LRjUodHTsie2AUn0NuRbtr1kI0I49
2C6M0xs6hnSeTbR4HK4Jh3PflqzlvOO8jZznFPwNV4tiyb3HU6AKAYLcieNN1Qy0gBKscrZye8GE
dSGlKjZXO4IK2H+i6JYzOWLPuShInbuOV5guSu7P92IidO2Ec+4wPj3xtjss2T02g+7U0+T40oQa
QujN29Z0wM6tAVlx7/lyNetx+taSyMPOT8dH5YhC1o+UaZDK/1ARrvQ96ynRVwprDPA8Z3cQLlMz
CMycFat21YhK96qDIJjmVqk8o5I+N7H9XVh46mTDCpFE/eqi5k8tDvdjXS8Wa3SFjBw2wm0/IfuE
l55DBl4oEIas4alx1PnYwttAY8M2KiFV8bNYNLQkg4PB1Ds42gTJv0rg6nvXbBGrhpBVpj+3me/U
rZY6S2il/93oQgW2dCCD/v8y02PfFY25/UFwPPe3TcIgezcbkHI4t3mc3mxhVzood0CqD6kUQ2tf
eF9qI1pHFGf5tZsU1ERW+x2bgp2u6wkDCvIzORv9zUJo0A+IMe7m96h3V1bgMYWtQoKI1Z/ZbSnx
WNQyq+8URbmp+uwspf/mb/5jjg0pPL9FvGaaJk8e3aCh8ttWRMgkcMVMRzyEQdB1C7Y793ZMMdps
RCyBbVXCjhupM28eh7VOHeZP00aWWx+/vp8sz2z+nS15FE5wjexnoKdjtuWBmdSnXjLWY5JEdI2r
blm27e9sD9HX6pn7xBRrl2C7yQFwOydbOGf30S3ZJN+WBfAEj86wE7hlWj9a2d5VUJ+oqtq1KtAJ
ph4Atks6KQhLVKeH9YK25ii7sUOWRnCALtJaFZxiAJBX2WqNNTUKOU3Uv/xTD+YF3CGsUtL1WGBE
0yeED56eGW4BjotMAK/zx5ig15z9UouzIqo2vV6oi3Eg7fvPaOhqvrmyBRUPvXId5ETHmYmKVyE/
aogU9m3ALZzNkCMDlOkC4976VY33z1RfjxfWA0uyR/EUGyYCxUIY7e0VzJ/YTBIjKsPWtlkjnjo1
eYi1c8LYormZXBg8c/Jyf+6lTGqG00o2iiBMhU1sf52q2Bo4dXP9CjP0Rd4rNPicD+siIjklOdrb
eyhspVZIHHHCxItsQxBq7gQUIJvUtObB7wDisi3i0n3FCZclpPDouDBAnlvp1DF/fnBRVVCZjzp0
Qx7vroqLHqV+InYkzGA/tqa2hlJae+8pgNPO5fAZ1EopWtVEJBYi9NAfDI1eEZFQfFPKhPAcALSY
xFPenS1GCfHDTXZuuYJ6A3XCFIvGJX3hfZn/j3owqddMvDFNc2iCmojTL0tkHubAAk9cKYyPL3X+
1R75iej88e6X8fToB7xJVgfR9ezZBH7y+L9N+GP/VzPCZmhS/CAORgRkJebcuDKA5cWqd0UCta4S
E8gEyRy257YhG96ukhKjBuZvk2aHYCoZ5fGAOu1xv7TI6STShHPQOLLsPwQKolSSoqPm63pL0niH
HAgLAZOgOn1XBLf/Vwk4sTLyUMs2gG8CRUrrq65b8+WlLFu+mH+YI4eBmTNhAUYTx/4dCoW+fx4M
SWcaF+RIMOJsg8UI/MiBtZQMpleDPDo6R3dG2uzIW/dvV2lesaYmL73nJ4thy4uQSywn+02CkBWs
NeAsFJpO0MKSCeipCe2RppYA366TUkkhQkXprSy073iYZ2mbuSULxh3woTkUTulIeyCzu3fa1e3P
/gL6ocJnGpbSWoKhp7LeBbE5jtQLRz3tpP+Zu16ZkVOk1PKuzXctDgli+sg0g8ru8Q/2fnFqnbjw
+gkl5b2u4EXi5y3ToTTNvi+WANlu/OWYcY3cQJ7tVb3O88Yn8CM4W07mW45JQLQCdNNhkSdWO9e8
i8bbgRe/roj2HR/hqhS3QP4cFvrFXgaXRwswwkRM9CaQPwjF4P9ZzLqQUjB0Qoq163t2pPFFkejJ
SRGGUWK5IFY1TVGYbh7mvpQx9ONHzoKV+e5n5zHwPhLHwBddZRSi3K8pAk4ntQf4k4p9pCdlkS+U
3dMcklGH0wYN7YUqum9xTGQdvq/mUZX8qc8XI1Xd0fTYpXPXdFmmk/1pAWW+9AZrJXuXew3fkP3c
MUBRHJfkHcafRaMAoYYJJDHTO7CC5f1UPZQR8+VuHrZcZpLqgaO96zkyV9JNAG2GVhb6ia6zTafh
PR/GS9/sKYZJJbf3O79n/OYuSTwBcybKL0kUpiWlHcRRiS8XHF96xyLtDmnn1xRUzGbc4MQ7FEdk
YOFODEqPjvAJGhNMy9oX6pxfrp8nTZ4fXMrwe6Fty+lJfHAV4v8zL5sfoy3zJw8V4DGBt6MTMnbk
PPcs4nLnfXlncmyB9HGIlAlGxwLH1BpgdPuM5CKdpqlDH88iSk7kPShFjNAiFFzYfGJRGgRoYwld
W3ObOkqe72vFPfgasdiDr+TrT2CrDl5G8RRs7ODtrCQF0inUgErMmGRKyK6YQTR/EgKdENcy3aw7
X3lVmn8ZDInyaDZd5h92GfxbtvmD+wONv4c+j5ztTXV4DbXIez8K4oWYFkLB7BL5adlgs2kup5rE
u7Qf3eTLI6/ppzjvTacGBtlvv/XaSkZe8nwQlnQLTBkGuyHHJ8xQ0S0/niW/ama8OJ+58ywcYsYR
hhRjaaPIeIOZyERXkkuQyAkFGZ3emDUUS099iyUbwzE8CFl3pleAAa4+uP4+oeaC55srdlcd8eyT
eFmWus4Ds6clfkqw3LIZiB5yAYyO+ql4/v+X09iH3Tdyov2wCCp/jRnRi4PFe6grK6MwQtVjGd29
mBjYWfpMNtsRVsVG7BkL4EN6h+YXCEYs/zhBswXjH73KHh23QhLRLzROTkRxE8oeJRrQ+GmOtY5Q
boPTb1oT/2LKXPBwRGiVosYiryMKzzeLZ9GPCaByYWJbj6mjvDK0fLGo2mbODUikT418JgGxQrVF
JYdBNbJJ8D5H4zkgPRqyLQdpfcY/ga+Ctadk+YvxHxJqmo7z3d7+FISxkp0HIvGo+vM8Z+VyCM0F
qcoGO9VTAYXqZ/LFQm28/ulRgPYgKmws5AqvR51SkQxvDXFQB+ML22tpkih8ezfFlS2H1UGKnT+0
ZcoOgAnng985RxD/TiV7aUoHOOZgStMXNUOq7r9JY3DVtBteCi6IwSTE7IfsZfrsD5eDuF0kgRFV
mTL4qDAQdX5Lb+wBptzyAimjXiFCd8wHlWUmxoXmUAhIMLpVTWbreJUWl9YraCEZk5LPDZr1QX08
IqfIE3SguiRef9tANLaMHE3UsulHeEuQsrzhW6Agwe9eqZBkF1/o76lhuuCgE2tAnbB6Fif416J4
ub6DAGwK+XjoCt3Z1hdUKd6+9G5KODC8ZhcsAnFuAd5ZupWBKDxd/iY3UyzJrd7EnGgkGHhr2+Sg
/xymIvmsK9c+gINTc3UpedNm9QpmK2nbwaVD5Iv+gNhme1CBoiLhpu+P8BXsULS6+kyTAFkUIMcn
yVJaWUoK0+MgYkEegxAaO64RPQOsCdcJ6oORBZDAhH2QrN87S/o/mt9bolnr6B/3/sSDbtARY8NK
IxGhXomPU/NWcVvutqnJAllxfyyZT1fdXp/UKz4yxCqMBiAc8HC0yF+xpJ63pCzUcHv9ntDRWQox
c6YHcS+T21EyUPg4LC3Z2GroaFwelckSm2NnBugXJYjHudiJMW97upMkxIXdEdzZwLOm7MAMbNCs
OlOmLL6yYNshSIuymq/kcLKpWBud4VofCUYehQVGDK2cXt33LOGz+3NG0BsE5Xo1MuPuLDT+Tuue
5qdveLDgl3A/k/6M/BVLio5r4mvwtdev3pvjgRw8URkZx/C4vj5QFh8tF/dZ2KfRS6BqknXg1xjf
x7gBOF0Ij0jkoTKxfxxvJyQXVvckbuhNK/pcTY9ghWy0l/6/Ncr4rEOqdnEXPOXuBwOE771PqaoZ
P8FcIyvXaYyGGy2rgS9erP9LvEMHBqorLavWX451KQczFKSJtclmKsni3+VctQJnVBM8EPPk/b21
3Ck7TOIHUNgTv6wAHoIZpTrwayJwNP9qg5AgKDsupDJz0Ef/Efc1WwvXKTMKuEt7xCPTnbw+T+Yu
1cvc54xAQywMeEyb4BVMFF7J5+xoULJXRX2iILMvC8QTDOA3Xc+pVKdCJ4djkIDLn7Klgo6e+mpn
ymYJDHSTHXfqh7c+PW48zfkl/p7ycmlS61tJQa/L0wuFxJb+n9sOBmNPAxKm4WgEVSi4rGeKgYKY
wMWXaQnuvdKHdK/Ih9lYDuuvjkQ6EYbBtvY9hTj9Cz90bDgB53NnbFWWejOFNDEHj/pRfdHx8a93
ACrKo2qFuRIJQ6r3V9s27wDsL5SB8voJbKtSdWEgOi8MKzpr4QMs9qDXtSsstDoqrn+ImRXrwSiE
SgJ6HnQmKCkbvWbhVEUUTfpPmYiiF4lTbWLOTiy5a3RpkO3+hMwODGf4Rzoluc8jcegIXYv4/P8E
+KiWOkLRUZyMTC8PpIq7AQk2ujF7MWlAS5wa8dr+Gh6WdPz68rfy4SS4bPN3I+gBwbiZtEtdfJ1y
GC3KQtrPyikrCs8s8fDtPufOb4VPtGEj3SA+NBGqEPyG0z6+1aamULeIajuB0fRM1EtEWOdf4IxB
TLLp10QlNZWBYcNOLlcwx9ESRT33B4GQcU3hMaMaOadtJ8Ehjp1KoIMXLBAi2EpDNcP1q8rfhR6E
0efqc4a/H4guCGF5yiQbhTV7pJ+w28Ljeifko9Fk9M/6dg2HUtJxizga9pamw5oc9wXCeCWJexJH
uIBcglFBt99am+f3KjGLF02NbH2yrNOZjuCaQeDF/qryJtZ6FzFRxXweLGTmHjmht/x+7XoHRJzc
hvgrVGs/ImxBBwaiuuDsnjqx6poByxzq39MO29ZvYiHIpeNAANG5dhkTeU3aElkkgQ+AbK8/g5Eu
GCR1fdsOzRJBSj9flI+Hs7hHVdlqbRtxRpGugT8n5AM7ZE8nMS1Gmlt8blZlZlgYeSUGp5W3e3aX
rWzA2QKlDjQ1U+YYQR3Ys4ll/4kEijvXZKQe+8qZ2l3YRJBuyXstNhT2YUvnqCvGORTICBvliq+e
mgOuEBP56l1syfHZveahWuVOFg9AABG0jkz9VWtB/JxbKGuDI6MK/v3y7Prr7SqJD5EAqO/QxX3X
Pp740lpT9DOf5OwbF7YCWENDf7eFLdxaeB7mLtE8lkPEbx6HygZq51Tmqdvl+iMwK140xgUYD/rp
j2hphK3R+KetRb78AWBFNYmBG6oIE685jfLQx66Tdt6W9WA2kuTKe8DuATfc+TCoDGewulOkJ/32
ehqr+g5VFxhfDqOVeAR/X/Z8fEZVBnWrybCIwDXb/wOcMIkuMbq9tKpaWsHWiLVK/gRHXr0Qd8KF
Yn0yDzKr3LvHAxskKMQqQkBG+agBucPEGn/6g95oKb8IAe9X2hJelPbRwIrcLa/CSXjThe3q8BPV
K7E1msN9MJ1xQWdxeUNx/9UuUdmKiT1DmvzPlZXsOg0bF5y49jf5L3WWdBDT+VySLMTUT/BMSprz
O5VNATykKF7w+yBotvWsq1lXdLwxs3N44xr07tj3UKaJOgqWzFmftSPLQWHbs55D7qmNvnvtGSCY
UqHN2dCrht8H/oCbefGqMZyEzoS4OX6IZ/Nl5hytl+2hgzgKKTQUbpuvPozAWPYB8bVwigY91BG0
fx9hucFsMRZtNGhp8zuvLT/rhJ6MoECRiNcYam4/NmRXiUj0evkQOU7vbOEy7ZG/Thhm+5WTlD+i
o2gvNYcEB0FMWDHFkA4NzsQ6JpH/H0xXLRDT4MaDQtA7LXH372hhNzZYueKcu5upbhXmd+BWUA0w
zI01+v4PU40eb6bVH3SrKEoXsTAeWCKgRqoOuB6M1pba2IUk5w6oir2cZ4O4zS5IaA674Wm/UkVX
sJ9pz7cbtaVXh0AOmOTZ1TVQU2wZmf7mABlOiNjlcG2GT763NxCq84HGpS1N0z9C0tiKN92InIOB
hzzRWZHu1HFMR2HKWgvzzkaLJfPr/ymPtHVFel66Fn1uI7obzZ7TB7oU3liaQLwwUklhdqpcg95t
J9rKiUAznVZf6kj3c9fJQdWBATrF6LU7t0qm+sPo2iGB6qoBovVnOZS/q8sztPd/IJcuCw/N2X3v
rFbpTI4JoDe5gXx1+8xWORSbFoqdsCiZT22sLQq/pPOnOdKzBUCJxU1nzNyqqXL4/uO8il8jhvxL
iABbSNp2MNFVEegwz6Q+ZExRkDp3Mi4rDOCoYQJKfTzRgeJU6GMJV3b5iAnjIkt9fSBN+ccXMrHm
aHa/4vrNXqdqgR5pP2WBw7V/Wm5Ssy9zSUwHo5RzFljokAc4xBcwLTT24FSBlCcBkIW8Re1Gc1Fy
xjRDyo9Fhzh2MNSHrVHgInG0UIy1iunei7QddNCQrO7utUWUiYLtK6J35yN6lgBuxRPbq8C0g6cX
wZhlMA4snYGnlgv+k2bw9yFT3ugbSqxcKHBpVkjcXtUz7P9CEXZSvFttSd6HcF+7J9LZtW5Yrb7a
XxH5ivYevrcME/hCoM0kup2OjjciWUEudAsSZhqwbIayBQSWNL1TGmjCoIGo86MzCICzNs+BPniP
satXXaZFzJdGi6amrhW1YdKzcvWIo4p7de7Ep0lA08W1r8w9Ua3pvlIkWIaB0CIEcBtFA6CgKkAu
xAn3TYZ+3hFNMC24Yp9m9+nEeNo0LYzk64/x1lo2r6kF1x+o2xHAoTl5Vvg4EfwYu66v0fc46ymE
BJDAzUpzmUB9eVG2DjPT1UDt7GDT2+7dNCgFP47dnmk7qS5Cq5dZzgyGqHlad1SLgIgoo93rLnHA
+t1cMQf/es0/CgZMycxHLjT0ptfgqBlrFtDPzMW3TAPEh8sgc38C6+J+2tiI4N6VLWMo5xKPkfDm
VtuiFlBN2wmh+TDjh9BmDDVTIuCPzhGf86orLHspIbE4/e2GmEckM32sFMhLxP1OXa4H2ExL/fnd
aBvHMD6GcYN/iJFBXVM4fPx/hjUWrAE79tB/zooq0WeXTbKpgL5AjcWlKZ1R0CquWhQkwS5wuoeu
jh2FfE+g43hseQsHK+FQsC+ODx9wru7EhKVtgpygEe01zAXqqq9LfJ8OQu1Go4ke8MEJ8AsR/sNX
bZKzf/0WT1TtZIAFuWkXqrVcdF1z5vL9VSQ8l3Eylq1FKFuMhg7pCPXJfLzh+vQDkSu/2tyEdDm6
ocuSbQrpLKgrAEAmcSwOFpyuh52+EQP748GV/QETTLwuZSm4TOgzBgRo+iUAkOjfDW9s8C2JlAFR
6y+uIUmu3lEsG6zJKk4+W59qYSyQt+jgrbOdrPAsTYXSaUrXvTfn8LePFZQeF3AHEHL0rF4cjrqg
Jxtx/gbVKBaE9Z0iAggXqHipsXnmxgzTEwPtmV1gqzVTzlsXLI4Ci6Sl2efCHY1WCvxDNht5PiVl
Nxovao7ZZYRdy1R/3+S53QdKJuXJ+wJNdCy5eBn+TsjwSCHrxoE49cI9/A3C/iqauhdkvD8J9xPO
w0OddA+Qz4M0F+7nEk9f/BVU13CaDuY+ca+YNqAvke1O3S+u9ZC/xRRmownvFJ93+isZBj18qvz8
GWQDspEZ/3Q+49mXb2IeGtZTJzFnr8teUc79Oqxy0vXyingjAXJvClVGGADZb3A1ZvPlKLNJ+B28
9weJrnhzVOK53jR/Zrvj1EwWFSlqzRXDDMZCcOoZzv63Hl55XjBtSMKqJ19WefaSq4VcJ1Rn6Mm7
XN1Q+4gxRRZEmbPHcyH0fNyPgVfk9vzN9I8iZFGKEKMEpR4RE0k9gA6xLyCSe8FfjXZwVIIUuryW
vdl175dU3GODHBcigwxenj75FCnV6QEr9L5bURgxAKKqRLwpx9hBhmzOmxDCUB+BocrYpXVP2k3N
2MRtFQpfe8Cck6w6f7uvFWR7+wOmoU1lEi8pk8PCtNNlWFIdqAoW1/t1fa9eMnNGFaVGp2QxNGPU
+cMz2hFbOZyByv6G9ewNfsJTaOUQjrTGnqV6n1BcDdEbKIWAyzmKLxoUioDMy3o3OXLpbAqgTAHG
9Y0eOaDTYV7wiO7W3/AYdh81S6KlEf48qLdcFplI2DmwMr6X+7E9uLxA/ciIX3RNnhVaW8cLJGRK
2suLM5D2iUJh5oDH3vwLlcRdxTa6dgV+QigQMe4CcHaCgrpgUzR0YB+0JEOHxFxnuVsO6NZjc+VZ
PCViAPe6FHKuOePBuFDBXKld35XSTglC/Bfd/O+rl+/RMSShpBK6iA7chu4wTmtNSf1Qa0oAF0s9
w6b/IYEM2bg+yBjoioXHHk3yl7m6o1eoV+2nfWGCtYQ2MOF0DT7OuPMZRRlMPDHGTg4xvTak+X+v
un3FYaAH5x1RIPuZvOshkUaieidmXfAat5h7fTUlTQNVbAjoF7qP/D6T0dID2y4qG5nAkA4F5+KE
uWFgb2P9aaYTIvIdnYZuloRmwbgcZzJ5w100UbElfRB/c0pcwd4Xa6fLEZfXUq13cLgRSEPM6Fbe
F9mrEuq2I6OiW/3/nWNTzdqgOUZq7Tt+sgjN+SQE4CaXPn3waT3V+L9cDQMOS98GCQ8/Y8zmSrCi
yHsg7tuMCZenFCFbaINIviez9vz/MI/r4XvSwfVZeXkmq85SuH4A4rB/oXRiUVSxiA0Frp3Rq2kG
6QehgjJ4DI2mJsX6zmSfz5lHpkfo3dEjZfkuh1PzFcNBY83pPR90V6y9Wm5WmeUJdn2oaWTKYGij
Lpt5Li1aSE2ZcCK+2oEKn4HeAo/s1KmQJBko+JSISQJ0W7Ix5iC7B8JokH7x5F5eidkeoyi2GLQV
L+zMDopa8owympQv2yUKwDiWmb8D9uJHqRc0JeeKVQwiGB0YQaOlOqW2SNooIxe2HDSlLLINAVgQ
RpENZOe7g48PLFjT6SuRItDg/qhW9jXpzLwi0k0/3Nv1lnGRgewTZIBToub4mr7Ufr3ztvadF+wv
xvIZ3r/+BUQLDYTCqINRCb1aj+k8HqBdesZgCVqwNc8JzyDSnSituJi6XeYSzwrnBTVlZ+Vuc/2i
xrJGCKxfXVkF6BTgl4P+VavPJRaZButszASJE4DlBzdchPWakl0CJU5lw1dpYCGjIctBCYcMGAKV
TbWc8vhQHD974k2YtklJVJdmkqaxYOkdbL1FpE1TR1AP9zzJMEF16zP6HMacyjtVJAJULy/sDMov
fQnm/oDvXPSGfCKHeLeDHEdSBadpRp9jOHvNK3yHT6pbenuw4cyX1AuK1Q+WKyclo1srK7fWaT5H
GD7BGSjAeHKhaJiXEMKgFtX2ybhH9zxlq4hQVXdXQ/1vYn5VSkc56YicB6mpD2rCB/tg9dLNFGCF
leHriYdfYpEnfex67yFzygwNI5ctR/IHGHx22lsCFxrTT/kPgHpGb2I5WVsxo7KRDMxhdFI2DCrv
yWvqFzw7WwDwyBdnrHn+LfMtJ8VGXNwDD/ZjsG90szgb0pNX2StA4npw4ox5p9VBdjXUp4YBCiMH
sQuSIqyuyiQObyyuorKW8/uv8TQXbDULsqJbHn1dSIP+Y1zAz0bs43O0ZoyUeYaKAHXrDeWxilPM
lJ8MtcABQgniU6czl2kh8zuWr7o1MnmpuPQ0GufDSmm9Hfsz9AsAoJXRHm66mMgsXZZkDqX9UCHw
gWhY1B1Xvbc5wwN7Zky1QTf5sC/FZJSharQE0ib8ucvumE72mmbb8z387aSgxtqqj+/uzw1oK0NT
/HP2iS/wqVJ+4U9XXQQBniAwxSd4cLj4Ny7QgZiR9JcLKKN7SIl76wpTAp5Gf9j3JYJkrJmAaSaD
oPg7/DvpUgyldX8I+8y0ka7MKhX3lpJjsUyheAeUsr6CwrAjYo/S1/L1bzTSWBZ8eqLl0/KJHBfn
HUlImtMTVG2LblfEqM+ldXVuIUnQEOw4rWKUCtAl7PcsCs9wzvVMzxdRmluMdjK+MXygokftkfMh
W7JJ7lb7s3mzLDBhv1bpW6xtRDN7xyt7eF6veko08uKEwUz/6pKAqDYHTug/aPsq/aW8g//plIgm
UnHBOWmM37QYg7LkPyr6BJGnCFEOazRTzCtbFceyQXFZ6/n2qqHlBEcW8g0mTD1mymWBhCTDUv2K
m3bOfzfULQfHdp0JRN68QQX7ayKeeaSVQALul5jK5mRY3zOoDVpP18xLVeggA/mCYPKIj7TC5xwz
vpTzfj7cJqmc5BxyS34cxDTXCh9AtESZSJP72Yh3xkeFwfe9dCyT569A34e2KztqU4AxoIKj9UF2
SNtic31eoeAQ4HktXDHqRlrU85j8lFTW3ynn/hOgQoNmy0f0QxFUeOu8vVUEnoDOxZMMjo5XF63n
0Ywux8udpxamtPKXWBW08LQ+KqTwFyB/H0FF0qBXLH1Jx+lzIR2UrMm8JsmgWSYPb6rv5Yzmss50
v5Ua84Os4TX0XJ4Rt1RTSHsczwBvVYdJfUyrqWX4sgXAcXWgtJMm8g3+m4D/TgZUVWq461fO6c6D
sUGmXN8Bf7UuyqsUU1Hjfp4oRVK+8XOtQFU0uJBdSkx0UUtOkdzNJrVxjrwCD/evwf/l1uLY36ys
BQmdMA31RA4N+EfiP5QthX/LP+aKqqbNjJb2URVlN58blYOZ1hqwek7gSI5A9HbqmCrG3hxEr7Sv
h2HfIj21LsRp9uip/TYlPlhxUQb74gaOUqqgdDvVGJyhVbSsQ1ehJWBwKy8aVrsox0GrTsFpy/CI
e5TqL1jeYk69oLjRuQ2Dur3sHM25kxIxcPQVZcydl0RJl0XxgDubEWqzhlzrPem7m/AbOHU0wP3D
4qXrwJeTqjaruytmcX2ox6SwTWk3xIxTILx4yDESQFa04SaT5jYPvHvfpY1vVg6JLLDlcuxLvGAP
XQaTHsV6eDkTOFejhtK6WngfHrr/a0Ho6gjGRWGaF0uYTdo8no+h1tvpFLZ/UhVLna64KrDkp9rP
RZuDa4q2X8WLGdI9K99lHN6BWJksMnusSBIN4ZMS9EBT5D2AAsoDklwVZZuAU7+9V90DjyBMRny3
QatMISX7sENst2WtW7YxDxYBgV81U7nrdpEzV9PEZI8BqHSRAFMiOQMMzalQQU2tuY1JWkQrrM7N
Jyi8BAt5MHqObEGFCXx/p7pzXD0sWemAs2WvHvawWZdR+wYm9Ip3qTPxrH6reKAuD5tztZ7MUXqx
fso31SYmk4WCcNJjmISOFbtn71V6kJc7ZyGropestRUuGrpws3QPjmRYJGyNJtAGAKMSd3QvjEWy
A3urogWPcyDdESm1QzvawJYC4NOxP3WnYCb6MG5mF+N7hhWHFTzmDo/l62dcAsruqNmWfTgHK8fv
yT5eezfhVrP5RNLP3Xt5s+hQIYR7s4r6S4lMQJAob8c1Ku7qOD414Qr7gaWDQNFEpdwDNj/pd3s2
91nY2MwsuPPFE5eherlvokAmk2NyrcEl0tN+T4W46uJSQ+sprUELPdtSxMwLvXtfTelB8S+J5y1v
wzT6XVJ0iUXKARK1MKwPYXeNsgpJki4NoIlUm7iMDdtEMoQckMHXcQLZ4HnAebIQG9kzeIvAxmLC
w6u/qntcD1Gobul9/g6hki/zLQ7+1p3zRNBA4v3vRXr3oKeqx7nOKgUZemSgaqkpwKWv6AG6jRYP
LT0HDpi5Uexmt+TiuWzkhNltJyMHMlj1GQXCDv9tmKjXo/WuuQZFz95HsStAlNiJWMmXqLsazias
M79OoptPZ7wHohIucet2ZlabUy84zRpGtBPoG0J8dKsPvDfOB3dy9am2phf14rwtmIXJk+CwB9O/
doo2difEDUWB4RsnrnnOPoct72tnItXoWMw0cZl1VNBkYaakANelRAgK0GyM5An2TOSUJxZ7n6cL
nodDfxXBGuXERAx5Ig0d2ZrKwSnMUA4FuxgdWk44ADp6dtPJMwF0mN5CTqLQ9STzu03Eu+cBFWO1
6Ml85cxwAb3XLaUyB1gWzUH5e/no92dOjqSrsGrbGeOWbn+c/uc1yCtfjwW7rEjnJ+3zORr5a4Lx
3qmH18Z9pK6nPThVyMyEO4/brNy73CV+xz5P/3/lsf9TujBBYAUL4a+tVN1eBSQ32icRdKDLIqKr
9A1FOvFspQ8vTp4dETgz18bI1DB8YxLgltkWd9LjVB5fYPzo9kWklgFuBKLWBOLC9XRUWwn4QZF3
ZkSJCAimAtLAR+wWAv1qjGQqEvLIhall/Uaex8w9w7b0jQB3QZODqnmmk42ia1uv4mx2ys2SHJ99
ytVU31tyEy+rCNqVIUvMIWbS8VpIfU6axeJX8bKY74/YaDUVdSc9E38onLyacJ6aH9R390jmgOxI
6LVgJyb/vyz6ISildAi5x+GUjuBdm71SADYxiCv8B+85Y/uXEbfGyxH7jAMhwW8PxW+Py2DU7U7O
OhE62TLIywO7w7ylE1DkAupOGFEeHhrGgwJ9fk5+mnuB8LX9sl/eKwpp+lXKfyiniOx2OxifowLH
F5a7C/KX9zemtZyeasQQpdqUhym4Bkz7NAeJwIyO8txsAQs+rBF9u/mZmFfcASKJXFYn7u0I6HVS
h4fy1CPf5amoDHqR9GvpevQqR86+V49rGP3Oow3ZXyKUXyjudzvWCwtBLeEzkZ+0Eb77Mof0hy3j
LTKESBkrl7UOqmQnGsHypVYftYx/44GpnPnwYE8eMZln0tRq8PUi5nWGOVZrCFy1F3DEb/WZvtHO
mhDbJ+wBzmsJy7BwGlAUlPKTg0lUVVeaBcTouszCdtnaeGHr1Ma2qp71XrDyNce+eY9y27Er6pau
Fk2kouj8kbVkFnZvGzUM86KAh+/hzGTMwdEtDkN1n/H6wmnYYnwtSXNbyUTHO49trrPMz3q4yfJa
e238moGU8rgU3fydsDOxRZVdzZd672o74tNFcAa1VP610b/V+kdfRT3KdQ/swDDuyA2OSnPx+uHq
6/tjZPoAxtLmARkt4eyi1cf4JCIFNcDJmTbY5xVCFkjy4tawNuSijBSH1SJWQ2pBJxVSswiyNcYf
f2Yf6qnCLdzFmiEHbAQ7wedMJCnv1vBBaGLGNZxgpWjnfhSlDpRdl1/zfviVNfx5nkx9WSNLA/XO
+5on6cwJLqjrz/BRy+knLhBEwoP42acWa4wUppfag133zdwvz7E7kUSayMjeC/sg0+pNwhskqgrh
nX0AWJjR+8wXXRwWMg73SrgvSR1JlnuPHKHoRMZdI/6pJSMjr0jkSicIhmLwcUzP2FrOURrsYPtY
vGJvdXaBtUi/hueBW6LwmhuDR2esWXjns33mIwNXjiBQIgaIb3U+kgxa0GYW5SDrNRuLaORWC8zd
a2tgb2gkTFwXJGPC+VZPCuWOXT5iPMQc1noPebcuvm54WkDmgHcP59LD4LhBM80auevvjJtQvO6K
zdHFy9vUHdokRTCYRhfGhNg7l/d1+/UMjT6Bc4oLwe7d2joHfvCpooD1V6qmOACjyo6djDepVLD9
FhUChTuG1Nt73MzTq2Oo35LK9Ur0pTjI11WuUD0AD1SzjUIB7tfuQ+OcED4GA4iOK40bFyUAojkV
oPZNhJCOrFwpV3TF7ToyhZAiI2QqG5Lrcu1mXxGya/oyucAxQ67uIcMKvmUxsF8NHcTbUbR/Dfgf
0i4K3TFVLJbopsHrD3tIpcCNZQUMY1/fcqOoCj50EsppDiw5M7ipeuCMFU7BoepJauurnqETGnYm
y5Zn6J5W5NY+GKkeemWqNOBB2/D9amGR4Eaqj/Rv9GCiJYn1M2c5YxWmj+SB9mCTXbofcZDppfDV
7w1vR3O17IPn4AurtAdsaWIO2B50EaeDJF3e9JJRYY66G7E7OGTu8QaOgKpTiSy/o6JQj2+fdGAQ
2ap9wEGAve3xXdI2kPih/Rl7hw7leNSuIiNfrGMpi+aQouXBjNnr2AI/CokTe6Rswry/3i3YE17c
lAZ4nntOD0V5mvsYe9+8W0h3y746qVYvuLB+lTjPu6x2ZHOsnTSymlpbCP/6FEaLumWK/bzOdffV
H1YIpda248e/Y5WMTDg3RwgzATQzDPjdXlZwWs5uw75SpVyEkYVNYkFu8VicWy7dhZWqnodlEmVQ
t/iz04snEu06MqNszBCzikuyHPPPvXJXeNpPDd0zyrkuYuN9taDlOyxiYjfhMnal0c/LLccXhePn
JnjKwxaZumpzoLl6/MePzNZ0Lb23pYnil4KMVt/LD2UWAIzxhAXDYFVtRuMBZFq0h7atLKQUZuHT
pTeCqy5LXqk7Xk/n7pYhEFbXaLcJfEdZwl2nuPITB7YPx8E4iwjIwREijnMBw59iwAzfh22/HpK4
pDlTUQupHmm8dgHHz+m1MXGIsSJTkNGE0mrsNq1OmViq0xJ+En9Z15+DO7zhc//wDUyWbvfeyP3w
GbgTvRSVIRy3iAKQh/biUkulYzMAkV5MFAexJEwR11oWkMSyhGOh2cJdf4eqW2FRVpI6zrfcfUF0
aIoLpgJFtscUCUUdVmZMk81wOVQbCc5yR70V1lu9yWYBjw2NhZf4AyaQtzNSZ6ihywDneaOTbJZI
vgSIrJu1StClgYDcj2NO83kPRoQmzQzZO66PrVevtx5mXNMHYedyo430Xu4e6huOyUMtoUdSUJ6E
5PUQvinz9gMgTseSeRv53+Ee6nkMqNkBPpe04J5T2FZe0dWoVGqTxVeyIcrNYUspSQBDeIumSmLe
kmzLsCrTjrtAWYrFfBOTQxKDvE0wY5wdFA7LGEdvU9CzGgx/DnL1suTCRAeZq3xNyvz8gmSYknic
BxJGWAhOUFKAt5qrm85hxHnn11BrxhP7nmkxFCCvjC3zxP6JxrN3lYgMQ4gXzGHjtG7ve2Tlzv6e
/FhnG9qC94bfhpGGQ/U2HXK1ylFBxxAmdaMFIgLyCBkKM5aurUqJYeFECUjPXJGQh/VjCu5OZvwC
iCn5r8rvKlx/lEOoAcM2F3A722U1AJWqXHR48McsDr4wJFyTBJqS/Gs7zHTPboGfCO4hufoFcNbQ
1jVc6iGYUEpwy6UoJFGCGcRvkqKT1dW6IS/qw+2+il9GlbvitvjU+IhS4M95wozcR5q9pt8y1U++
9Gfn7UA7yK/h14c3RQ8BwisO4+mT8tDuK25ihEUPzWZvd7YoLIU4xmXwNwy30qZwop/9vSPh3I18
mstcR41yrfXDA3hB5HfU0OhE2BwiApE4LDNMymPv3Uq7XbN1IMpF416KAhoDg1OMviYM/Lc0d/c9
MtrVzXctrEj/cWoWH8YvyzyCyfgKTaKPX+penMPdS2dslqLxvkkSOFLTnwabFfPGyRcU3IJxUwqX
0SqBbOQ7J/uOwSYYsfUxwTkXhzlxc107yvP2S5xMvNBTC9sXOz7+U75JHbeHJwEhJlOSBthFi3mz
cdZ9zMMtke9gYU43r3AN9WQYlLLPTASrhVKwMBFP5mnafUecBrM+1nAPSfXWjkGm5DiEa+yOkpVA
8gSyaZmNjdHj4WEd5KOYR3sZoAMPw9Ymrm0NcP7nWhRJ1LsczmdTqDpwIHpisRFDmbqz9K1SHG0o
dF89i0TJvL+owsr/wtxbObFTBRYrkOqM/IBNwCnNA4rktRUIkSNyC6zj9aU0GQ6C/ivQ/S/hu1hC
QxLNYx+Nw2TcjvZA1cnweG1eds92zp48FMlBeqCbw4ORcR63xVvPAfVauOMsfJt2awZlSN7sGOVE
YCrKH9W7S5SKqW9lVkLGuHlc2298iQso76K8NDdLBqk7D0Kl08zVJSrfXgdPuZlUGbnzkulfJUbe
bRRH9BWs9yBo4cZqco5xUV5Rjy6C2SySx5LypVfDItIPG557IKDbbWiiG7mQq5SqlguDV0C2odr0
/UOftxyi+20KMdTgWE9QWdIN6j4pOHpBlqOi1s4mPeIq0dwwFZJYIw12boB3gucAtdb3+YeaZ+t2
wk8LtHS5oFEGzNi2reeFPRdHdkfBtvqpI+QA2At8NZTPjegknAr7fFZPOyIS4ZMO5hbCrP2KFY1V
wCL/vPDsmjc2sQJmCezYOgrdNgg+2/TrjrpqWrCS4Jp8utUfp8lrIQgwZ3s0kjvcTWmiQq1/h456
dm48SnCVSl9rketVGa365A+Pnk87FBcpsvvgUbEJNqgK+TLp4lkzSNkEjdyP5dfXLuk/01o0ZlWR
4Izde2lzz+oRq2GhNyZzjAU9JWE9Kfq/jt/r9q6jQxE9t75sJp4oL1EBAgbfQ+PiJdhlTpmGws/H
B5SSirhtnbyOVCTvNb/lf/6IOTq8DFK3G/1J+Eg3RpF7XU4ulx9CUbGICxafGjZh9c80POFyw+GS
0VRCW5PGyh1eXuBrQYxb6JM8G29HL3UEx20n1pAP3L/1I2CjgRPQ9olEOup6V7xqtJiZn4hhA69a
bU45fDfKDITPJbiyrrz633MNElJe8atf0nhhadJilKmDpUcyLEApqlJ8S0oFhVuG2/SuDCbCa7UT
JJePR6E35KKtvqYpjJ0/S2OzL093XYuIj+Uhs9Xq64bHS4JInAA79WfsgAp+rgmvLQzRUtuDr9LM
Jg1m11PUAd7Fq+o9VU4sryV4TPH177zpuk77mOnzfyj8tReOjfj1KftRc6VGbgGpL1NpaAaYvKrE
jCvVvkVMRPTn5LmFzgqEaWfeFlxtCz/4F+5dSpShj6Kv1tBCS4ld0cRX2B/AMSNpxvH0qd/Ei71G
FtoTVHaCGoBWtFZpSpPJk8eby+3Xv2FlK2yRhSHO6dkaK9ozPBA6sS3eP1q2dd6j2zGNGH4j19A/
6/U5U10xJwBftRIvc0yA2MRi/06jsIpjg+ulfTIBLHYap/3WvxHjYVm5MQZztW6WNO4E9DwCxTjW
hADnOfF4jPUr1Q9qI/g9QCPtjz3/TEBaNUKzUq3dRK3RPDXdTpxvc+zAgGgMz4IZmiEsucvnVjKj
m193RCuWquS8yJsDelAJOEk+CcCyl4bchE4AT3IUHtOIfJzOd2/dyHKw7XvHV8wF4nqqVB5r7Ujj
viobw3v12EM5HOHl+YcK6XQ9udbbzpGfBh7DePZzOtsBe57uWhPRQl8YeuwN+v7cGuRYtBHHtePU
pQT7dIcsQnhgdlOSugU7n8Z1E35riGDz9xbGiAMXLfgr088NKhCGB5y5g4KeJVAqw6bZunbQea5S
e6mlcM1AGViA5ueSYPaojD/LUTImaeSw8jtIavV3bruOHmXGjLwmavSAthQW4MCpwXAIrFQc3Jjf
+i15F+LEIxp5h+x8nefcR4h0bHsiD7A6EaoElsx2Y+CkJAKw/gec76qjesgccF/z0x/hP8K2Vrgx
75P54m6j4JlZ7BOrKuA4mVxxiNAFRorH/HQsxIZRzG95/DrbkuiDCCT3bGqs58zN7IWxLGH0oDhy
Dr1uQ3Cu5Ko4uzTGEXU2yOQYLE25M1aI6nOyT7cLtVtgQ8/rUfIsQBow6jnjNORKF6q8xcMnUiIF
h8l/SXmlphQdAk9yCX8DlVIXStVEQgvrNgEi/gPAMusNmqwZBFmJOQ9Kz+W0ihg8qTFTOSftKZXL
kWnbzIvx5K0qs0txcBjNkoSClnFqjsyq27GjshdWePQIXS5wVG1jW55R3+Ch0GUpSJDZiTwctI3U
f4l207BmBlDOcdFEQnvLvUd0QLZti7GAgvVkJbHvlIrjf4bpHGYIY3pHxFQfqzDUtbNY+L1AdFCz
6SzVDotTS5NkU/fDu9QGf+kpsFZ2wh8/QMfwSP7vRImcydaYgW5j5W3xKQaqHBAR6W0hyjKLq5ii
8S3YmM7vEIgoNazpuI3dHqo96oRBqjjxCnFFzcL7tgU9WpryqLH5p6UP42E61lM5aC+HjMrlOaPD
gJMWc5LJ7zcvp2fN5z1Sza1yFqV0NYVS98sSgg2+BHIhUfK6/rtoVj6pLsF/B9grPtsvCOj+IhuK
FNtX//Pqv0uTo+i/0PBChXdfV2wQaCD12Dwb0oYqj6p1/37CUXzY0t+46J9uLggjdqGVCMsN+uRT
fSIztvIdZBCJ95ANqGztDlbsdSlyzj63DZ3hUUsxTeyirjL+nziwToLpGD9j77aRFLMPU72HUNvg
qlT6Dfm2x9LYv22IHRU1qPQbYzyvj6EV5Ca17pyn1yA1sr6tjCsGXuzRfNHEoMTS0GjDQB0nVgie
W7gedCDqwkJLvi+P+EjQe99qS5R5dphgWqNsHr4ESMAWHh2atMHp+OYkhD6axq00wuVwMvA/LHiN
n99oYWix6eufRFk379Jjd5YaJPcyLv/+MpFuQhCPBpgYoLz6hQmTaen/rWty4Ede3onm6WvNvLfo
iOMTegmElY2TotnY+2VGAV035TI6D1wP9E3Kr4Sa09b1U/L3Velt6r+880UtNUEPiQaAWYPcBuc3
BkhXiXexkOeATRlma2Nurx3wv1XnucgKb+5UIWOTpPF4Wik79gwWYws44YPYJzdWBBCDHp61dvcK
6fCK0FJbKNbv1Vus5W9foblzX1FW19j2fzN9A7bCLCXR9gLvmSDDCskwN9A7ioCUOa9wo2EiohxB
7bCo9BjeU1Loat2XKeY22TkLtd2BOlTh496BgL11fNM5sQfDg3Oha1F5RCSbUMbCOiaY7pXsFl0b
2588DP13IxmwEKnzbS1b4iHrccwlMOCj95YKRABbTBxNOsUNff4ruUd6x3ipYrOcquKmad6+gtp4
WUm7aJLtrnRR75FNI8DccxZF2VgcAu52StAag6hv7N5pcInAlEiCYrWLRDNE2sCVrQjDp+knZEd6
Iy1JK/Csw14WrDA4P5Tm5OGvgni1lF+jKdk/NfSGzuf6XaIYdQ+PYQQQ+nFXmfwZ6FAcYbVJo5ry
+i1yYVFax4dCyGXTBcfrMVGJcViXhKbctt39NIO6Zo6ETmN7UnVDyKfUfeZ76RkcVz5oXBICajMJ
iYPPtXYW+3FsGSx96Zmk489/itk5XU39CiCYDVeFjm36LZDa/FTyWYmlcUOljn8XnuduZWD8tHVU
IixNx8iSx+5/8D1TNBeFoeKlOzK7kX7LRgpPUa6Lk5Xgb7CENa8bjOXyjhfgfTCXmLbXJPZVOKgc
yTMax358rODCZi3H7S2cnAwUy8wcgz65t5akNg7xd3RwS1sjA05OzW2RxiQgPfs/erlNz9yfU1on
q2dRiYdis00gOGhoCbLSY7snwQol+lY1eqkhEx+oBCYhfPTI6ypZVUo9ahU7klZS6dtt/PsRYzm9
yuJK5nMQjmcJZE8hO0y2cwwmwlLXyYIZlVwDApgnc19vzQoIrSg39C3FSxx6E+MIW9MsAkSfmDwP
SZXhB3yQuY2POKHkGwAB//ZOpxluZn47o17APzc42+uDpI9MTwcRwuv8AwPOURcS7Lgy4jtYHjJV
abs3wuy4AhKReOv+GwA0IVqF4FmrJ9WQW8592sa8ovLZyI9qv/ovlaGRyyBE6Rs++uK5i1xNDj4A
RmfZZ7nHLXou3hZslv2koayXuCa24aDG3A0asCyu+hoKST7HkbQItNv9odpmRhORembeluRPsR+K
ZvVy8iGnAzz3jWl5vhS+gN918M36PXWY3El4RbUEvW/1HRSjt00aUJ40DTUtJWl/gEfy5MVZPsPX
VszBy3Jj+BONK048789TBNg1pU1anB1wGGLj9s4ils3JkFN16RVKsdjgD/Wg8Op2hV+0ZyovwBCp
kKulw5pZA7jIwXNr/7vVSEtakqVT6TbVDtHrrKyP5C94ycp972mQTp6ptlvYAwD97EObE0vHXnco
aG7Wnj4/ncEPfWBewxtoDcpngemsDLf2+ZZJLAmai8icIcADaW97bFscUpEd3eeVTMBLieW9Ty5T
nZ/HSd9dXyghu3jykikqJ7BC32qh01P6kCKHGWEeOHSNw75WFhYWlrKTPh+lDQpCMUoSpkRG92u9
p/C6zXzKcobJtiSF+PIArDKIzG7b1sKOMeZcm4FUeQg4czcyACsW59fh4pRsDQ1zceohWe41xrAK
nfp/lV0i/nTxv5m0YFkrIGfvzGExFc6bKv12yyRBEud+OtepSYT/sbyTrfpVcXTCA2T44kg/FdEF
+EsWwVrbcK/aM9TdKOaeg4M0JXa0NDM+ee0nXxCveSdDmD7tpJTehsRQRu7fOM8M4ybPcrsqV0v1
ww5+kvdA0IlrcYBaQOf/OvdGhdGFw47T+5RPjRj5MJj8bhjcbY1/ahbmkfNuETHPAOKYTNO5dwqd
RmDUgqxjXEIn8pAn1E3BOrYH+Y2hU0/li9BJtbiVo18KaWVBTUUPDr3WaE+ZI7ChEosL+1keL29W
PXhw2nQjWuDyfMLlHIRQuUevvzXQ/SnAGlfuJpxmQ3C3jfXnR8QCAxS0J+u8mrJhdOlpuJ4ZsrBP
S0Q+ALJPcWHcwuf2iTeiAGN36oJLGV6RFQffJLk3UxvPlqMFMGXCL55+h8AVZOomayQb2tBA+QYu
9ZabWi6KFB+c4D00ki72wNBSWygcaRJQved2L1WOXioVmrhKrNOT/+lVVjc6Pczs8b0f3eo8AMlP
JQQjKBX0r+EMXhIe8dHcCjSCh7uB9lPmYyhs5oFNdR9TaSp9EWP8UekkyxZApxWWX/+/wgtrutPD
vnbs3XZGGTzq3NJEbUEDe1LGDmNIk9eH0Vbaoq9bHtC6XB+H2CoLWXPPljDaRif8o9BbwaCYofne
eGHfDUd4g3BqruUqbtRxsIPnmJwJsGq95G+r9r6rh5rP2/3vdcFLOvL4eNrX9vKp2bT5W1jrCLvX
PVW7tUlC9MMHnDYXayQor6JrRARIqWGODcByzmRUcK2ZTrvVQ12+hZtVCPMtqdJ3NToF42j0aIuu
5WlsglVUwhpjupQ6CNpjBnKZzOV8EJ8+wvJ98sN7ZRCOp7FkrMMzlBaAnuhYlKjBTkySgDIqaERn
uZDkrsT1ftt9vF/5r1acnuWiuuaW+3KW2rTgWGTts8HAd9+6MZTJnLFVMhOkLDN7jzEq7643FYxp
+S+Q5XlvKqkh8x2mnkXP92ns6QS6+55TmH20a88/3Tr0zpys0biaj50PwNnEpL9xxN1+7fsyvhgD
qsTqgR389tCg+8QsM2PVMQtaNCTh5yuMDOEesua1Hg4+TeTSGbw4WQIBFC6EkBrF1g1hxJ9abHLg
VG9Uvt0G+rJcKVjDyaM8kESl9x67GVHAE77/nwxepZBQ+5vJTOCkdnuHcAtAFRqbunCRn6NyLIj3
qBqgAeV0SMeBNshxeHwOu/Xj0deU+YwrW8kf/K/zXCOb3WetGmPGdEX7f9NhUQoIP8IpzMTT7REd
hfEqobfIChzSozB+bRPTVgtgR2tW9D5gbY3tk473xe/ce2fpgGXF6d0troxlCu/TbP6pUIf2XAQf
QEFgg0dO/nlHu7htaAhykdf6hNDhP0o2Tv+NqepWDqLJHR1pDPZTbjPOm9mZZztTZ7xaPxXtl+5m
rM8BJYnF3AmbDBbxzkXm1jMpd1BstAZX7+QJBP2NnVtnpnHvV93HojqzPQdpEQc9Dq4OhE/uaIbr
IxToiKmcoBwCvdsDyvCM9CUo0x5w1WFWeG/ddoluXKsE9Rnc+qSQyA+ACD2AXXRe/C46jilIUPG/
TfC6wehvvcCVMPhab9oLJVa75h3BcEaw8ZVVeBFYmXS1ycdUNIukCkuhMGb0TcD3YZN33Gq8HtRz
I2AF3z+/9mmQFe+RLOuD7w94tPAhNbiTi0AOd0ISjyhIxGV8Sr3DGw/r3PaibZ6jTesZLENyJzyC
IEpH707UpMP/Qv+aabkZzwiVtcgbwRIh2JuiVSD7q+pAG80E+zrszKCqbW/jrA7IzdsoSeOnwpJu
1kXJJZgMYrzGTIWDGakX1vWHUJS1yK5v1NQKb6iLNnfTCSOhfgkPIFXj1xHt0GCb27gKsYEXPGy5
Da8DneuVUo3mfQccqV6/N40MypkK/q+Mk6l9xLhPPcyUMv/hCPVBiOJpwrtc5gCPOHHjogLuIITP
yFbGmynLKZLVoh9TS277PQrJ1JFMu3wwPrbNJ7e8vJkrTgSTTPUPhP5QFjYmYUv/t4IeexTcrMy4
4gSS3eS6havRTWtvqwUY6A6OzwCn0rFryIwuMHspe7j3cao3dJKD3Kj6KiBKIxmcRhs6tO1FDC6W
7lT8F3zTlprx53+gwicGxIXND3vmK7satOgTBENFgYHh68riFfcmSXvMFq55n8JE/K4ttq65B4ql
DdpRqNJ//HkbONwYQHqDI5CauIOtt1vLr4NSjaDx/P0JmMXuj5BE907nQUhU2zF4P8/u0ENq7Z6O
RTomi/LBg/MyMbmfy4ogbfeMLoOPbjzB1zcpyCW/yJ0zWmf0E780jBAzgy2CXoVnKnaZ626b/hvi
MVJBgDXa4w6mQyARAaiVmRCnHy0RmoT1lC3iS4SvIYzsWeez2D0FJHDz94H62VsEgj7crlQADw6t
ZQjfDDcx0iWcABU5PXR5UoqBiVbVfedPnLnzakPCtGY/RXAOxOeeE4ZLEv90ivkyBBgtpViImK/w
SHfmzKFez9FcOL0eEeE/dQy/XPhArNwkPtCXj8YQb8SKplCpGMHw+DIPJyQz/R1pDExdsx9RUaCp
bNPgIKNngGVMx+eOeuAeCkopuDkvcUtUahJC6Dqf6s7mZ2M0wbeyenr9wssGHBnrXRlDfbTaXCJQ
XnME79CIxhFMzFdDTWNFeATPopwEtSHAtoe6X1lDv6EDSUppKpDX6CW8BUcyFexvvxRI6lSqmhJX
OMoSC24NTB25dUM0ApkAI0ZAw5tpgCQH0lKWo22TkKaO3hB4Z356y/jKcyVbG2aZcoCHuw8sww3r
7b9vj5bVJIb9JAQNZFLVjeGAXYOtm87TjY8uEFH45yHU6A7Bq1bGjunlKfuWHpWjSSL9jvIFc3VQ
OJNKkuCy3/lUagqTTGegb1z0b+NKXpVIE5mRXgROVXL2uj7mSzQGkEJS7q+PKd+n1vX42nQCN8kD
v61xOEfzJP4DPTDbBgxpfbzqVgcHQOd7cP0YWLx9YGUgh8AnGlRhh5JBbngNCRYdKaACeMSB7W6h
8MmCRXUsoSwY0nJR5BAzppwn9y68gohh7ynDGE0GSMhKYI3hW3LZTCng7zI8CRvSd7V+hhV85gL9
YlBKLDT8SsaVLulgxRvDi3ybiOzItdciex3vZzfKKuZIcaIbVhU2mmed6aqDBcs1a1vaGG/8TEi2
0hohHHegzv4lXPA/jqPawjJjJODGEyAspBfJkiqNLr//eKlkXGIeHFfgtbC3qdAzsuc1LfAj+vMO
e2xVW42nURZZSdtIpH0A6XhaSY9+tjDPuG3MhuOWRrP9zhVyqFkEqjRuEK0gHdoottvOLNiFkMnt
zhcRMk0SVZZl1GSNLmXNIbZmECpqFZIs8p23+Jjxg8+DgMPyNl5ceiBH5/+vnYrYEcV3l8EmxYme
HnLWVORKXp/UzbOP/mDdZOtr71GQdhu3vz9X6EQnkpGLSroqEf8d1wY8Txf0tD2J3C3/UXGJizIt
4Iv0sBgP9of74/1eRsjniutndQ9PU4nRtDNxQmxB0eDG5eKQ85M0BNkF5+I5pHFYKLYhC95FkmCS
TxsS/DNVdVKFPB6aeIOY+6Qp/bSiVYyZ+t0Fjxr6vwQMmX4eqz2ASGa4LE8JVR5pTMfJKCed7+Ox
Ixvr042520nB0ocJo0iGiIhJZUh/g0I5CMn8aY/dofA5XJpQ8jMGF05RdXKutfkskeE/w+9NWK8Q
p+zQr1Q2xlWHbh1wiM/8O9TM2bgj05UERKLda7zyrX2cK+wdA+WkTcyQpBZoHM75nMAQe61gbdJ9
rNIJ5uX7YJoxcMH3ntManebBEIe0IZh5HDBGQHojGlsavhvz+K8ft+L/ZM+h6TrT2zTORpZXKm3w
n51XnP8PzIga06BjoEIGsRuyC/kiT8BCZEK8FZrqhFfX8wx5bicrp9SNNVQnpi/Pi6rt3RBX0f8l
LMkAXhn40xoHeqYVLORzR2xL6P/XCL/byDUOBby7G/j2fbr57VShUdvk1yI6J/tadcsQhIeo1GBr
kipYFKrp5563dZZIFuR2mWOsbPvzv2pb/p45tjIZBaCxxdSsdUPqrqQ+gHsnxvez+ZQ9RXRakZk7
GKw+jB78B+KGRC01Qc5YGNha6tqdlfDJBY0BTjK++mLUiWo8T5b/NqSsQwP+9p4set1B6DHRhwTD
iJ4X9uv/wq1kvU6fEUk/Z6SdE4Izek66hEqM4fzrnttG1/7pwhH4CcRsqB8DfwtBWDANCstJ/qBM
kciF+pT98zM7RUUtM8ut6KKrt4ND3LE01gU7jMuAi6GDQ5ERiFEHWYbyUI6SUK0/c0Bjimyjnskc
QceWOznI+cGXyW5ilq+e1hrrF7Em7Ie6qU4C7WWoFM1ozPa5Q8KPX0CV6a7TL2M216nQhsMouLEh
7wfUQ00Gz0uejkFftSCRf/+/t7VaP1s4hom4vlAK+A0w1p3D4CKJifSwvcdkjJs1p9ZV6kuaTg0w
DNiTBn6qYQxv5J2BJeg93KghgVv4C7OvcP5RiVQKJQaRf1hye4v2GI4nygNZ/Oc01aqBX/I1hwSo
M8mvLTlTzG+Ahj/LsYvw2eb8umCOzoG8TMKgIZXEz9Ip72A5dXIX0xVw8X4Ag63X0y172EQdXY4R
xkDu4lQ1mn48uvclfX6dA/3Key+pIzR+OpbeykD+t7flczX6s3zgzI51JmndAdz4g9GydeTFgHGw
G6I3Qgo5tKbpNftj/dCf8MURkHvzSg/kBHOJU4TGvGPdy2iyDJyaMUQARdPpXnd3osv0lIgRtuET
icgE4FAl+bSaVX1lxCz9TMte+X78tBr+nhP2q/aFE6HmMPOE5Uff4wx+rZ1/HX/3VRlNEa7pX3Ti
51enQ3GRyT3clUuMEiT/t25tqs/aJrHeqwrIkw25Ucq2lYQU5Kyx3LXK/QE4nzO5SPjafDwwKvA0
FD3WwrihATWlLZnv0Nk3zjAIyR4ttfRYw4nNyiByewF0HFkiPDREqimqvZOMaYpBjvzBak23wbRJ
NSAPsp4JwY25JSmHciEPnhAMjBTqYbOvfkmBUu1Rj3FtSrHiFPmyU9SY0sYQqD6rlR7PnvqBPqiF
afzHtyFQH9rbxRgxDVGzq4kUj3R1XtkN1TUiJ5078MISu7Pe1xnn/1PHxPtZKjKKx0UvaM8Qirpm
d1QKqTl7avg4bZoIg7LKSQMaeIdC+ZXACtqw9Ax5OEJv0xtZo8hvXcFwPyhkUkBRMKSraOetffiA
+Dx80gPe16MpB4LmjkRN7oNX8YHsLbO9nWi8LgxHmK5GzJHNe2tDB9fHcQtaNplhUPr+f446xHiK
cNt7A0KFYB+ZfqSPoF0zTXuCMwItHvXWO9IHKP/OOQPgjfqXUAndN7QpFMNADl8lqzfkQq1E+dvy
ogxHfmDjgGH/zOS/Nu/sRQSPGY0KeJEotyqhlNhLPi0CkoTVRV5wRukZmjyeOtn9tuUTAQSTLv7J
1stKpDPsxSUVwlNBIw9n+iFL04bSduaSDUYCIyd9Vowq9qW9ZyVv0eZXMtvManzNkAd2ryKIVH/J
OjBFFWM9ARJJ+2Aez+ZuLGZJvhl2DFcIq3r05P/Qx9BvNejVWVu/xBsshaPWvhvHtjgqYSs+LZ+u
nwVOeXNR0y8mxz2KcdndMcn/IFuJ3mi5bWhD8RhQ22AR2Z1Qa50tf4H57m5eY9fiPbLbfbQIRdmB
zoKO0xx6gRwNU2A4YHFIheh354eqZfXjg5p3Z3YKxXifIt2rlrNMRAkQl2VoMRaG3nuoUCZ6L04m
dk89vZF8XYqQDd49dqXumd8C0k4jhchg7o5rvP+J/CxmBXp3+6hmxt6RyMTpIjS8R2GqSGaZ6bP+
AW21ncc/0apoPytwzJekUOa/TOL34nPTPgdPK8iGxplU9OREAa142rLfFFo2IsvlJlJWZeHBhYjI
Cvc2GbfKGNuBKI4zYF4b05erRUT8CO7B86cjsBs3MjyruEcc+wzya5UqsILDihPdwXwXY38KxbSd
lrmyTee4QZWso0PKpEYAaoXsu1C8HYtl05BT1OQ/Zcc03XmBLq2hbPtHF819OQH6ugIrYPzJu5g5
M96zNZylujJGi1q1KB+jxVrdaFNY71ctl1Y2c8ltbvVFfp4BJJcbYxz+OD0yiizxnZ/3O8mEzeX5
FF5gvCvFDXQiVDSIF67AFcN9RCxeiaeNXT/IcUWLCkQ4zKcuEB9e9+yoEemFyQ3l5dN2wjgFKXBM
8yndvKxRg22tGNlgS0J2U+BqJ2C0qD5RBivfCv/2fZnFkbru8ZP6W1vPLj0u52ol0+0bIQ624uHS
LWwiP3jwjdjgdFOr0u5/h6nkTr2IEmBSFG0xc3dxvBS+jiM1GqUlohFL2paSCiKbOMlzwon6ugfr
Mh721s241/jny+tOcmg7244YHHcKIL+IU8vuIWKAJYEAmk4PcTRi/ipqxe2Tyy0i+QWw4j2iikmV
Lsykmkctv5jnlHTwQtZ1nk5dKtVx3ZgDdaiVfSyIZtBg2STti376s163uG4rNJQeoTEjano473XX
84SMWJ/hyJOjvSu/EBR7YkhIrjj30NxXREWQL5Fkn2gr36fCC0qnVKbT/717Ze6dNBrXjFes+d2x
GdzQ78HvglP7Db0FZ/cuwtx7HbllkNS4EauvO2KcjqVlycPDwvS7iT1qWa64NTRm7OdvX3G508sn
zghvDvsdYo6Y1baOQSqBpmectCs/snegS6vZR5MRElJPpue7dQIuHjJ38gY/ZHM+3AIxZVGM8gWl
k2DFWqRgpSRZn7YVak8KyJpanM82S1xzc2cdpECMbnWK/pV4KphocIsI7sjQusT/hDePxm1HhXwD
chpvTD0dDOjtVkZjMYoB0atorQ8KBX9t7CRn7f1EAfQ9l4x9TDVZgMGriG5btiJy1Y13P30OWdxh
BDP0TpW2i8VFaEHBQ3XDYqolEshIjqarvWzTjqeYrQ2/h4DpJagk3AzGeS2SdH6/zs3nyRvjyPeU
+hLHhAXFNuHDxaOFydWMh5hMvVLzuHM2o12zJl2fzbZKci/IZiRc+LGuFAEW8u0JbfBsk5bp5mBF
1I0b3KIZo9DUM+gicOpi+61wcWMUGSx1yZBt1eaDNqYFnTkfrjIYAE25Ro+EI4kpOJbBP+GZyG6t
Cz6yn5i+e7vWYBhW9PCPmbLAqmMayheCtS6hLuUQpVfA14DBk2ZBlrnPBCoGa6wmZ1eIwbULfWdz
S+d37IYsjEUy8sY35qGdMAm/rLEx/sENa4i+i9mnQWIQeHtxurVMxnyB5VgTC9XGhtSx5brYTKPk
++i4w1RMtCFReqS6UzYKFH4ELTZWhWL2lDIHTiBEzv1GuIBGJyPRuDgvliTiunPU5RlF6kyOpl5E
UiKPhmK3ZO2F9O8D5HL443W18kP2+GhLI85bfk+DxYBSEfuxubSLUnBlSGjWI71Rqx9fWhK1i/e5
9wVDB/jptRYLrJ8O0x39Lgu2ogL7FizuHAkx6IAakaVoWo1oud/KgblqriDaT0zh2rqM7tXcnIzm
da2y3KknG3c9yTbxZed3WvM9THz0VubAPq0T6a9tqFNvu7wjOVVBy7JGuZTBAXQDr+FYRnEJr4/m
jyAy3bZiPG9hGTuKtWxWNyFfvTrjWNHZ9rnebC5xR/AAgN3UOQHdNYtFV71VdHbdKaf15EvOZwHW
9Rz/sMSlfBgqvWYhTt2rP64wIW0A27QSKuZBsHgaLeO6xfZ1a9u8JyE19uacV39lAGucjqH4vcwE
5hKVBfiqEkBkQy8nm9wDMDjNsfol2e/KH12R8AE61a6FW10c+hhobr6vEsz7I5j2h8h2OaLAN9Ew
kz5ulwo4zjfOk8yvpXbYepZH6WvwD7dT8nHw+zslOhJmstyhcZdIEjRqNnh4X/RdvkP4QQ8wpRdh
IG9g82lhUDdAsOVT1TMWo7SfvM4jC+vaQJDNgslfPVWdnokpjGSAusodeAPViR9DK9eaY4j7e/+y
I7GLOBCvJLPiElbD3GnDiLLcqXWNG1DkbGCwTRL7vgmmNgD7DKBZT6OimO9BD2eHou/x8LlHtEbN
mGC760IE07nlKe68ux0FcMyjHPXJ0dCjzIbkz8zSX4qVV+lQIh4+XRkLtPGJngN3aQOAIs+7wUNq
SVQ+R1OGwEQ1a7C7SgOC05of2qSRzjxw49SivQoqlWNiJ6YCeM916m2E5GqA2Ln9SkaBf1IWs64E
GiKPw3i63OPgP67BRtyFPwvPuuISIwuQ0R6i9sRxNxP3x8I3E9fD6B3gZ5UEGLn8Xsw/A8afdxjG
SXsyeO9cZmhacWF9jmeKbO4a7OIY3t/JbYTOnZhfQC31HLgbhnB98MCGY+iU85NrGajs3sEg3BcP
QrbBa6urVcfq7bRF6OPJ5hIe6pWtt9nn8diq2c5LOiFKLd/+dXA62POlzFWmMuYUKEGa2VwvM24W
T/YmdqTSxYcD6ilrOyUapyIzp+4jrC8K19EOodOVsihiFREGJTQkdfRar01UMrfygsHTSaO2EXTx
FeTouMntppjySoMZmwH7Awc7JE6j8+Ua2d6bZv6KPqZmlu6JArh5kX8LQiSuoosm3fafTIFLsuJo
2RkvLCDtgUcVsNEODmnzkRV156Cb7q9KGKT+wDjoOtdH+FtqOj8vmBCDEsrgr+oq6jyP5DdmFUC4
qJLZxSxP9CAlfp+Xyk5As7bJNDajxsuX/YKGLyMw6crpFkhrLDywoy+hyE5wbZs4hB1AzCiCKfE5
Q147zF1hldGIwe+MWW968eJ9mvfvZ7bVgbv/qjh6mjXK4HDFbHmWCuaQK1/mwSKzstqsleSIzJT7
BzmAtjQmEKdXfJgmyCVTSRbWDH3zR4rtTITM3hhfzQOIzy0FXGn8ed8rIc1vHqiZPCo0J8qQd1DW
EFWjM++94CwFtMpk+zKEKfeEQOHF4yeNRVQsBcGoAvzic5YhnEpja2H3TJdRdnR3pA3af7kPYTAR
UgZVHw4UjTccTUveOcgiQzJgTnBSQK7kInS/fYFQ6TpNqb/4ErI/EW+tPuMwfNrg9hWQStnUgshM
XgW8EbVHa6bV+/hlVrKMT75ZzOCjMWjm/1QHPnD8kpO1OjDFiNod/Kqsbjm9fmLpFfZYxVbLzsE/
IFXS2d2wIBesa/afQWigKIHiEXXTDUj3NbrhYFQFbjqMd3Ds8mQeg9v1aC/PWG/LDuPToWOTK9d8
ifNOpSt0lZu8sKDcIctRAGH7T2BZwydSls69sDg3bq/l7VVg7UZY756ChdZlBwJ+MhKEhZJLJ8DB
lkGQ+juZENcYEeIyAFhIMUBJZBdP/LaDOuwN2G5tHVMAGoQ6qq0EGwP+z+04BWHAALxO4Vi7N9SX
8Dw+GwQ89zInEhUu+yAsSHajRbHMXJjRXQuaxl4D8pdtzgErMlKZD2Av9G6pRSPWDXI1xTcfAzpe
yMmmmeRKcEP1sTidETYxab6LAKpzFHqSFNtaEq6PA8FAKnbW4UhAzfFtPCtlGJHz0fTIvqiwocGX
q/Fx0EBYDtTqbqcRvNlT8vyELbNH8//lRDwdozFENsAv5fQlO2HBVjYCYq/CzCMqUSEqP14/fuOc
xmM/duaK1nvZTfPa7g0rK7AHGgLhy2S5rpPoFHqmsBXgDcWLbUIRz5mNIXsTKRphMVuj0n+UtsEa
zU6gWYy9LQnGjQ0uJYyfdMgYDFWdM5uNxwuKBIem7G3JPH6NCf3NsBQTpKTjDXBa1mj4UbxZc5oj
qhAcwNJGJwdCHnO1QMUajN990zHxZW6iJp5V14n8AP7QJeBI8Hc4spp9VtvUgV6AOXEfoJrIPV6N
++0+xPAsgB8o6iuOpf/Og5wpbXTY7CoceB61lbxxYDfEKlCWOZ3Es2pvKFAIRYLvOzLt83IPx031
iH+dX4V6a8tpOeUTXluRsoI9dnGfYnW0zpAd245FJoPlP1oLIX1KCV4YE4i6EO0reG5ETaRUyLl+
aosyHSNhgkVISr2fSuJRQsGATqi6hDApJ9nkIlwLnqGfDrG96JA/7MdzWskO3RybzlfOWKCbBU6w
1kEJ9NhVDQ54nVSpiyqVMYJ+1TVQUNd9UtoGyjZOiQVlsPmL7yCgbvVKOhjYndvfvCeSk29LZKZi
rirA7PBRUvpqi+G+CGF+ErtJ1/wTDofvAdhdYanBmDx7rdcNCvjFUZNfLJAHHh1ed6mdA4Sm+5sD
p/Px5XTMTMQrcqjjGZ3sQJR8VEbmAVBKLD3lAN5zWHJVNSanT3mpee2XR3z+E4qspERdwwZPUanI
m9K/JoSWKg7S+lg5TlpVvqwPxK0EjsMlggjH121em+dIDeND7HsYnAYsc8mTy2z7xbOPSSbjG9iZ
MEth6GrCWgDpCTJ01tUApBNr0ERKNG7Jst1dQWjF+wDdKdovJT/FfbOVg+YJeBrWh5Ex06RLwj1e
aOfcTs019tAkOGt/piscroljUQT0VoeujgdVHP+c/ChhFwuhdOos76yQqQy6cudy/G23M490f2C5
3hZSNmUxeTzlL3NQVV4OPdmvdLFG1o+HkjltDlr8IkbWTeqY+e1XOoKH5Lo3blcdu+TCwU9Ypbwq
2M8ptSRLFQ1Pw2a1a5DSa7py4BGWIuGJjppKv3qrJjKIeNt++cgVr6vrHofxMWQWrEQxHGyFyasQ
iAO00s79BleJbVP87Few9idpCHCJ5tsHaif+c3cFoYnNltegMN7Cb0uBtO/waUUQrCNUmrFnPAd2
ZPvzwrIkuln70aaAegFC/mgQ8ExjbtRTW2/YIAwMRpdDvzONdMqqy0qDV2OqJPEzE6MY/MlR4LoI
9IviNvwoU33PH473jWxeTMmgrRFyjSuXJNT0UrSE37VXDzcQ1FqCU+Ef0KWFHvu77eHLERFu849t
S1fwgopoDDBO9Mqh/0gvA22DYV01U1KQLUGzYrwwGG/vZcTqT2paTwW3WCuVNrDz56kGT/0dQb9q
24UdBiMiCg2VI4a5K2KUv1tSl5ld9Pi7a27fio6cdfGlwFKDhL5vzPPWn7kdiEYzVIsgjJfWzrxa
PZVEnkPRUnekthIijp8UPWTBXoysyBoX4QbOoicdXHIXp13Llsa7BSmPScIoLfQ5VVCDwEO2B0ad
KvJXGVDoHVd7gpP+VKGXUmSf/NbEOMIITbStRw+5aoYgoiFbeFqfv/AaPBq/OtpFNPVuYX4vAZEm
Socejjr6Nhcc+ElPt1AQAFEzxvlsDiKZKVHuuuOsd9DQ8J6VbmwEt0VujqplcHvlqYEdUkxXXGoU
Rdq51FEFcGB5Y4zmgmueiybhcg5kBi17a3eAhukgZuidyztg+fOOw+x4yItesmY16sP8wiyerpfc
FKiWY2AFM8ne4GS1TwnyBFD9H7FfW8ByfOmgRrrdKU6FV5yMcqLDpsKMY+dHmmh7kq8K81onZAYg
C3Q1RTQ7P/ZczAM0M4FxobwvTQTqQHWY5+jrECDzYNEdW4nfRegEMv+Eo8OpOYAFR6UPPnHlwdpS
HWKgrpymqws6/9b3EjQHG5NhZKwzhS1cY5xPgLSGNeDaMvKH6kpGSzHHQ9jR3vAkY4PevfJyDuXL
eyHeGXlSm7mScAvrC1kzfbnwnPVS6BDXEJ3emECAAG/IDdZsWFKOnWUEYA26LmQAf+C5BKhtiQdY
MX7e/EQghTs3ahCN918qAzEjH8BP+eKS16KGnVEehmy+ZcYxHdfWX6eo2ZMQRvazQ7alRLdAhnQE
TuMJJBVXcouhTwDZq5d3oPu9LLBjV6fUeWD9/OWsYgANM7DqRaC4IyQzEpzdr/+rLGRjMbKcoEj0
r/Mh5q4JEdz1UWuwUQ7wbLt2ivW228GgFCmwnoFpQnSo+RtHytjKgz+fpR33MxzNXm/60mDQtCR1
eUqCzHebwAAEAWAedTAcP/rOoxSe+55gmfyjeY+Hc0DFrEL8R2LVj/WhUS7k+jr6/EwkOEh50dqe
dsHR3Zy4cEgu0FnOBqiVEjdEqefeTUDwZtMBfbuC9aeO/tZEox04jozwsKV69vwr3sHS3Dd1JHri
hq6uEx2fsjxZVMgRCUwTRNQLb6ycXYWIaw6JSR0BWLSv9JjPj82m0BVquKZGwwaFnKYex6lLdu1G
m0PfoJELIv8nOY2Gg6cNKQ4jTqUQY/axqOeHvhmiPQ2v+/DV2Dv/LsWuTS00fiZ41p0v/huRJBad
vXwQoD8r/x+M+IEYsvLWIhSNT+E9rLU2EjZOfMK9YUX8WhJLtRa7EtGK05+9sLZyRAKN6I4fFqn0
xoFfqisiCSYZqNvjGBz0cWiVyaWag7DY4hqY5s2j7ZHhTtRDmDu26dG5lIfd4/cxZpMo1TaRoH56
FmtrlllyDHs0csGjifsCrgO7XvehK9OTkuJHKU7vxxXozHu1lTPyDeqNS15KhM1NCEwX52hs53Mh
MxBTZ9ALxZQaMAaU37TyB7ynfbb9BudDZ0NBc+jNqeiJvEKgpi/t93CLQoW9mbpVGRQNL5CWTsSH
YwQI/bIbfIYMbVBydTuZpK3D94+hGZRRnD3Hb23GA7+VnNmqwT8nJMZUWpZ1UrDuL7eieGm0eM1H
VIZ+6c39EZCRl8GzMMqk60Ax347Qx+gcUhCedZJ9tiUHlMOmytOz2SmP6HXbDwr+u4xfA9vGcpra
ar7TYjbhuDdaE+1bVf1uIhWHQnZ6wTc/lW+ZogAj9v9TOG9AX9rIIj8n46uzdhz29Ihj06OMFzD2
LKCgVOaS+TuOfjuBLp8v2ZLbJ7egOZ4nnt86stINB+Y6lb1rw6IYdq5oiGiQKsWYbUQ+nEOTnFrb
ttQS6olO/YhM+NmauqsDCalJO7oCMiC9/ij6XDNe68KbNCfR4m1NMEkb5PdFR8uTYPA9q4tLO35i
gg0wcYyo8wkCSSmWBvUBGqHQ+ZszzJK1gtm0yXmsF4Q59y3wfQUTIzro6Y5BZLE0c+5JjwhGtVoI
ja8eqD9qnfIqfqsp+MGYaLdUrLV9Wqi+MiRKQJ5twEBVq0wFf2GmDBTbkEoc5XJNS7v0TO/qKQK6
h7RNKVY5BDfeYs8o2uwB2lR+qQYg5ElsXw+vAiImIEXEDbNPmHLXEcUnBEOCr36QRO6Yc9g0F1HQ
MmPgk6tmtz0YrJa5Fr9GqCCV2yA0mxg3qJNbZFMX7fk/wl9MKq0gS4T1JbOiVLjAFDPcw1iOBWbc
Jx/4dn1CCGwh/KceSM54pDVH/648fooei0o/cjv2xncMd43/qd+VdAal25Q9yxTnsPi05L59Aiyw
qYkqVyjTN9cmPk2tAvLxrSvLV158wbBYXuZlXPr5w2zt6YbZtdhrmjE0U5KNw21bCg0lRUxUmbYH
l6gtAAQ+ILyCzh+q4YD5nnoruihvXlMA9xzvl5ANcyAuXW40Jq4Uv2ghfZ5b/UeK49CngS5I700b
qJ0n+O3gQhpbDHq/N6FdfJaB1ivZritQCOj7xsaZYQW9lb8tNDM8ywx42XsX5wdei7x+hR7kpTS/
6QLBuzdj7UBuioPLeiNdFvBzOqj+xtejgN8wp87SK35ZZVdvNz8MHIFRDf9tn/tV0LcCq6SaiWqm
WSPqvr6SdNkOJyY5XVNKTAeAaM1MbcUGR78QBIY/50krHa4Ql529kjiGOpmPju3WHbF16QzX6AK1
Yx2tGIsO6HBZZZkL8iEN4hq+LYfbfAopNwDjosGl1+JFiRRbt7nqIPCv54MZBS2ZjEYJEEaB8EF4
OL8475v2tzol4o5XCkFtM82dX1S5TS7ji6EH85rkw9AnWiFK9s2xiwt93+bTSGymAx8PKDYn3Pos
UK/hFRJFxkX5yEgpaxgW971iq/7pFVszsN2dGA2I5g+Mn7jV8Jg1/U1anhn5c7e6dt/aqMPEtz2+
FvMRqBIRRprN210lg2i/Ar+Ed4R24tpU+DvkIvzVPvRQXkVdqKtqmhN/3mYllmENupNdvq8f66Tv
ux0GbwgB/UxXvtq3ozzUuxoMlGzKa+K0PHq+ZrQOdsjRJyLz8okT5DKBL7hLccGXx0Q+kTgr+Lwf
BFRgs3HYL4SOnvk8LJqzDbHIMGgPqwuzOsavBH57BhaW13hOer+lUAjglmlOYMkyTyB8fDchIwh+
gtgq87YEzFv/n69lvE9OEsaFcJc1+wBTvj9zGqpV9e2cTYeiB5JPX3nnFTAa/uBB/F80759AlI0i
B396FYD1ZAX6vGOrAJQ6x8iabhysIew27Myyj1fN2WVCdT+s6gK/k3LB9tb6SNoY4NPRMmdMDWgD
pdPMoHxuHbkdly0zu6prJw7qTfAKm+wj/1TrXm0h7uXzSB358rJHeVOFKQ0prAVOpcnH0qxBKGg/
2Lutv3sGx8MKTyBbCIJJZoKeao+vGbAV3wbvTsZrk6EkQONq+QUyxVmXghNMbhJxS9d6mLvkRsj6
sJSDV4wu8jQ9O9yyjKHutC/9ivdcUrjOR5m27vS8DcbHzWYP8uVd9HiVaO1ze/55YM4WWyZQSBk8
El7EDpY5PK48VolNEPUj7/8PZUnZHwTf4cfk35LY8ggxDo5rFIRNuJEgYdut9Lv/TYvwSWfZ+xi7
dT/HdAx1B1BrFsZm5ShLZjlZlu9vb98FY6jwJScj1uiD/eZeIWKaX7icQZJ5lDhaQ0Gq7PKS0ISO
VyzrcBisrNPq/tKyN3fa7/zNoQI0gUa2pLDaJTmcKuT8FACjsJxROCgUnJIyvD2igY6OrLTuuoZ/
catp7BZoXC6LzVUQeiUwqmr0mx55vmF50MbEIO/shExVhv0GW5yooaNAozogESDJLy2N76GV7Hqg
WC5+95pnmfWesKS/QNyz6pIfQl7Nq7G0FvRR5P+5Lp/ViALGWsNgEwCEc13L+KejDnfeiPqi5Tqi
vEtGHN2Noqg5eJJD/QoUOxaFmWs2eEdWtOepc5hCXea0YtAhoWYEcOQXW8VtxC1hQmFHPSCeVi3Y
/Pk1WbfPGHnIg0w4MX6HBZfgebI6fjE8S3Pp4WV1M4tuYn1jSpfeeDvKWu5+KOiHjcgEI7n875IT
jg+rzGRkgoPOpySNcJKdCdWXC67TUBB7T8qeI5XopdweXfOZ5N+rs47dpNVpd+nJWrM1sCEmmJyt
+FYyUnBdM2+3VHixkU+hTHIvYGQFlAXz8bRF1byrn8UJykbAGhD/wojPkZslu1Wuwqd5Zc3V6fp3
5H6/bLFuL/MuDZxU5o20tQlS7BpnWrXQNfRjDR/fHZMu/W50H32H2WpJCrNN8ukXnQM1QNE8hY8B
kQZRLeMaoXOPREyMv3DZi5C/fY9B5rPg0Co0wJv3KpsV6JKEMJJ46q1nLRBjqWvkD9C3AY7h5/4K
MOWNTLUKFo3ENAtaet/gJUtS3oE1Dsqe4yUb4Uiuvbo4zVuGyyl4iyL7OX5jupSNA2VgktW1Db7v
FAVSPn8AX8ktAR+9OyqLiUdF8Rs1WBV58ot15YrBp7VR6iwJQk67POPMd7odTTTrDcR3lWaiy2W8
pyT8TBTgY3MqmkAvBSr9JYCZEI36xDA5d2Swf+IbepOqnDcqsXF6u0QPhUZp5i9GWzEH1NNzw3EM
uH4epRHjmD+fWj4oTGYd9doZlwUmrZ/tmff0czepXfuu1ADzdEZfUF2HQZdM0C+lyyVwbreE9y17
yVQEsDVeRklEKgbmTC9juTuXYOwEjh69HpEBs8J/oj3rCZf7J4IOahVFpKAeDbLJioQUgc3zA1Dg
zhRkg1y8ugO7f6dOvsMmwboedTWtz4luHCVvj0lnmSLld4ZzplzdoC+kqllmP8wzwBDwldvZxhRw
F/qH+jthdkBL4PipuCHo7yZCmJ0ccSVBxfNMok//c+Kn/DX7f+OeKnUf/S7xT8oKRRCaIOE3bU9v
p7zzNrtY2iShNjK7cuQkY8MHm9rN+jB3qaTwQ3thS5rrx5BNSQMmz3aAAbcDPRa8RhAXYfvFlmYV
CheJb6Hc7vMzg/XFxqFWJoCUWq3laibwCj6ICl9kMzs6DvBpV5xBY9p9VqybxShh78GKKVLq8LAW
wh+ZdNDP/yiZu2J6l1Gxv6b4QcYC2Ep8ys6jEbtGnbl/E9NTGyvfGWHBapse/xTs3XbntVidBLB5
LNeDkGyxIPPMnM3Je4PrB5E2Yx6dJyUw1ci1VxwWxPZzXEaQR32tPsYq0VOUTIMKuZJgZ73jmCaa
LG4SVoz/s1U5gfu2dVXvYKbp7bP/FIshweYn9UPHc1CJ7I26UTml/V4dwYBTeijD7RGNKQdLFwWP
QY6Pi5eOGqMB30NUrfYpp2GavnHsRQhN5exYuxMtiM+1nM9uWMb0vDg8NzmhjtzLDsSULd0C9hxH
cNfYgdRfx1Hj1AWWlJnJgoAn0sErtPj8g/XcUXYe5w3iUb3BL8FFVZdjmkSRfgR3641j5giVsuvO
InaULUHqOq6wVVLktiX1RSj+eFemcFkTx1YMoSXSyvqd+805hI2SIxSxsUQcXli+b+iq45E/8MBT
U43nDHzTgcD7qIvsJHKZwdo3yY7964xlfmmdb5G5ezMjktQsG+eUVTMGlLi7McTO+7zw4F5Ylw0c
DN4BHKJnzVVc9M4DFK76LmqrQgWJBnAj34NunrxVSTVaWxIJXzARDKAJ+0lmjGrGuQ2A0pQtiNm1
VTtROUvRdechBCyem+Y0E0hJbPwwFYnY7SnAl/aCfm2cZgzvPCUT9uLFL1bnUnRK359yFcoY0wH6
1sKms+bo9GSncIAJMki4rV1j/4akklOae6Pd7i7FobRrjdIrWUVBqjDLY26D9NIlZAVoIJKBH2Px
NEVZ/7hHJIqHwIMcRG0g8JZyM/HdYRIsLMFVpQHGLdcditpZKcZiZGc/6yDBxqenp7KIs0FXbu4i
/dIDXv/BflXBjU13w/gS033roCfV9NDTVyKiJPYhqLWxXw8evf9d52kgSxZ0jil6CwC1LZLQ5aQq
OyS8bb21YJn6AZf4VPe/XHaUgjDj6SoMRoi61F6HYmlRzfbeICYjReF/th+3xCN3fsZ6llUFj5m/
o/2C5pxzrdiUMi7pe8EckZYfE4nTlvqInqrdQCVumUrxVpZSUTNsWS6uN3hKtmyxFG+eHGpjSXeK
1dZc8Xk38doRyzE/aRCk9Y7hTIiF7VFEwgpQfs1CNAjlfSE6AtclaQ3M+AoxXbVvw1GcNm5NsCLc
omyFiiPSZ/6HXtEDqqaTvEIhDUn0nMzMteSJjlhcFyYAzueM5wEme3iph/gKS/E93JFgZ3NEShnQ
BKCD6vBYTxNoPb4fDh9QSQHPyXIdfeVxGizxND15GvTLrYxzeHtmUqZB62xan478cEegrUe8Drlt
Plgu5cmC86sDZOQfBItWDRT15Y7oBL0oe8Olu8SPigNlUcwl5PuW02KQ6rRfXLCPndSUSwinttsG
aCt0BCT/6XLHEcYrnM9cQwviSRtLtAmRwsBIE8sjnse3x59RbaUY8q8jRzCXdl3gRoTJpAm1Qv++
JcnKahopgFvdhgPmu+hyPItPuajEOSGnKNAFsFG4rL4+pySp6Rzx+5jYFnOWcorP8iFYnc+vKe1g
gq3DuelkJKa31XekgpkSSba9vyQ+3rvrsqg9ki5vdIxNtF9imTqViklX4QKPWOnl+0+df0x2BqAY
tUPEE7mNcuhDfm6N/AxZ0INnpSWFajOwFhSuH/MszQ4SJxEBmQ7BsOhquAxxXFbQgvnXdfi3Dmnf
GjOhsvWSR5jbKDPeHYPm5X2JChvfbJ+H+/sEuL2VDqVLxghaz5GbGPPWYyuRO48WKgVVTWRlK37i
002PrjKW0alAaxJi2NgeVsVHxDz92Nuj+JRlkfzKAdMDStC1k8Q4/bWQFee+BcsqJHwERg7l/Xdx
pwLQhrh2L7DBOqbFqmV22CeApvWYwZ83qnDf+W6njFDJwAw1PLmJBCr6XxRtmLIj7Ro8K1c7F2kv
9CCy7GivSHRWjkZ1PQNN7ZAKoiZji5O6b4A6lqd0TK06C7Udkn342nt04ZJYI91H9E/AYdj/tAfh
qxvKnzMQxlCDRpa89q+GT2por36/33xYFf71gcksd80VB80VP7VPwGPjnjRGII96FK9sKkYb5p08
Nanv+2hGsuYywwNwAen0c20zoA1vFm6UyU3gvsKwxALAL5k+uMiUyWS3niOd+nLwQXKbGjB162dj
fFGJLTvZB0Jcu+Yig10GtqA/aeIKKCmx0Wg1+ss9gTiikkd3b3YuDOJrSErWVc5O4f/b/ElcePb8
qJUE/FEnHt8PPgyTAmTq5qe1xkdknc+FnwIXYvlG6BP6RITbHvcgyw8nGKxmaQJKkpJ6w7ncMeme
pt5L12Gs5wGJ0dGJL+Dw9rF4whUBbc6mE6FkQIL5d+DH5j191jFIvu/LyzYanly1dZVb2ukz0+jq
EDTAVB/+kNfnhmX8YGWJDnLQWyDuZbRN3+V+UnMyks+JdkPpfT0kFMxoSIEfcyJUnxzUAtO3XDtV
uu2TUPkuS6ovevoXJpejKHPR9VO/H/sSiiPz31oiILWA7PJ8PstWWAywigt7+WYQva0ESejsTbCg
ZVDMkiCpgi8Um6zU/U9tKWh+oSguvZdsUpeJgLTIWV9anx0aLKD0ds1iYNaDk252mli2DnImX9D1
et0bpr8Sg2cCwdACsB0ZUrlLxI1s54XlkgKok11VdPWoUPmy5rg2oBbxOYivnj+5DbtOrnfILF3E
mFED5S1ZEGFVbcKctPrdy6TINMtXaX7OWqKH7sD7ytfjRjulXApuXjvQntCqSMp9ygCKjyl1TuRg
8/B73ZLab+fnWuwTZdwFrxKkI6/Z1+53ly11izkM0OhhODNXLSK7TN53/RPJ400pc55nr3w6f9cS
lAxNUrzSVU/Y4wBC3xui5/0a5eI25JuZConDRWb8sI7byUYbr3C2UWvQj7I4c8tKNRh62bc1Dv8k
0lao7BxzNVGjWODcmq0I/H0d3GvLfPV8Btk1xq8TCo8t/9j0Cau1Fs++7YXmL6oIb3FAbcPvzWiH
l5ZGuQXu/2aPTT162yhP/ASt8U936ZjOlgzotddlEItCcQDqoZwNgTCcZhLS2/9CwZRJ2a9HqkSZ
eu37RNpzpNIFsYOIzgMXde4Zss2wiGJAwC1iApZ0X2DJFJU+TgpNhvKINR7O+C2gFEbKg7pthtD3
Wfh6yvcVunHb02QYo+OLWLcdP1Qj5EhMuQOX+MuuWGzlt3OPIvCJA3Bhd5gjXa+mcBD0XLQXQClR
NJi7vT6VgXfxisMx/H4Rjq+vcfhY3zZE2pvmY4Kh/1H3fxlP4EbOTmswTVJQtJgTitBVKcF4lQd8
I52S4cniu7pL1gMYon05VPGdaNJNCoXfLXm0o9eRb92q9PJjsByKC7n4y1l63/Qy9cpYwdyE46LI
e3iIYHXJqaW9OvTBw3bd2bEigU32MAITVwLE39yj393jI1d91NsyBIIHUevKb9sRPgeZzJodlSjd
f+onEqfxOZVyvq2oFGYK5GPYZGMhTEE0iU9L/GN4mE4lru22DMr4q7IMYzEDsEg9FLmnqpu+LqhR
M/fPjzS+Nx+6N9lRUdpPm5bDRfJknGYuCUeDtkqgJWlpSwE+keKVrmSCAgFmqddXm/ZxiRG3q7kk
nCFG8QKhx4zVW04mNeiYmSjYNtWbmSZ/elhpsYB2yKfsxChGeWoNoTp9EIVRTg8+mqJSRWuZekKI
6YLk3dVpw08aCBsOhJiLziUAxZRPT3uBHIeAMEEGQ100eTpfvizbS+2tOuIhazdAtdewbkrV+y5w
v0ux+EE4XCJNAjjGt7xd8iNUNSYosHsk5jQZVs4NtGM361eoV/xNswtnJYHYZ7uTfQaRVfyVtysN
VAihp4qxLitqlDQWFCChdv7CcyMJILOGhLS4J271udB1FZ/nrts/D2GRTqJdL/5lghPNfRHyX31e
Xfmq+FqIr7om5anUQPDbXXT9644ILJjBnIyTToIl5KEs67XCcFD0IkH/38IAIVMnL1XIR6sXuwQc
bEM6CpvSIfg/pIgK8K4FD30rkgCJyb0UwdlW7XAepCPV6UkpFU5QewOfOeNfMJRQTZeFSorDCBzs
1fqOtt814Qf2HlkiKIXWAG5pS0ifUgMvjhwB2540c1lLL9iMFxBBLeuq74xD+uDC5QVd3rBmu2OU
ICWxq9D12nv0FbGjoKpwTSB3adVA72ESXrMShugfGYsdIFP5AbSDoRCvsAueQzKv25bhY8QoPU7w
SIAB1DGtIQfSGk6VtCXf7sJDxbLjz8fmIzPL693eq1rVzYz00rPWwiiNBmHezomvFDC5Ln4QZnid
fTUzXTF9L0eAsEzNYWdBhekSI1L1EZJf8/yyfDVH20L9x+Ux210uwGwFjf8K0n7IfRHiwlbliHzJ
aULrEJB+8tLsdt9Ao7IlEVPMuwhNpmOTwXEGKfV7M3Fs8fRtGovGInOWMZURS51Ck464zCszichL
Ev5jO2zT35QFwMb1ocFnvwu4OYbd5UUozIR74SzlPfYn+vjWwZ0/qFAQB5guPKyd86rTjAc4ZlqF
4KW1F1Ya6qeIl6ajit9Z6eLAD2VjXRxiKAaGyXXyO5NYdOpS0brzTlmTY8BVNsKbGjudDSDorEXt
jBreCk5h9SCyBNbCSuKl4tudy8ZAtCxUmLSrVYmSucJ6vm4Ud+5QLIh8CS53FfglUvG1LmxMGVwU
5csxb6iXP1coO0JtxJOG4cB8kJCkRef2JvASdI3WULlGtQPcuIuzUvmR9R/zvcoL7zGLH9X7ElkO
5yoYKEi9BppU1T3XYgOFGLG/xJEuSuCWxZ4hF6WYkvK0d+dtyF1jLJYOxmYRi78h9HVV9wnWifZc
2SARmVLu++v0xtYOYNHWQAeUc5Uyy72oVjay+AgXKQIujfbDMQJoPi+GZnOyC/ixPGpgRE0/iXKi
GOShDe6SZW/x8W5l/tMKdJAvDKiq0oAN5yOfo1mNAkct57ardytYl4oxaGB5JzO7XOsCFJooj41g
m4mkykWHSRPxpU/1FocAkBWqKAITXWP6rRVyK21sc3lk4ch/l1FlIsesGDp8nsM13AFNKm0ECIpq
zsX/vC2hit6mR/Z9gnDYQ233S/8xZ9XIn6RzkxeBMqiKFIvuhllRxrpM1T3cYmgXXivKkmfG0ORX
eYZV2TmLm7o6zlYd3F+njJ2Z1UqePAcPrM9cu4s0Jl5WatTgW8YkpuJhjsew5AP2Sk3YTUvr6lx1
RaKr2juHz+lVsld2lGf13OtQSg60kCswMtc7jLkDo/iAYeKTPvhxjvw6IGJf28ZcvSaIlWcUW0Sm
QIXTa/35rEmBJ/3hN0/EVBXgOw4rocMxKXVyxQj0aDXmvszMMDB2/EhXG7LXiDLt4PSvDDL/QYhu
QQ1VyfeyNXVmOT2PjPnwgM4Xuq0dUSrvgax2HyB2tSSfoiyPaFJGHP87C9vluxJ5bKfOqHnSUAkR
hSbERWD6l9hzRlETHlpxYAZRtQ7K0sjAUwmfFGPksHn8kURwCCM8cgzg7dmJpzPI2OCVtrmtT8/H
imP9UEaSfZa+lApQph9Cw42yyJVnglehkeP+enMQfsQnGJRjZPTdijA91ZFCboDwBsMLJYIgbIGs
csQeI+SSMtpVA9nNyObYj9Dzl8WdRpXgV4Zpi/2l7lKk1eLZJDdGD2Q2/3YSTgmUVV3y+M7QtLFD
2EWk9Vq2DTATZvbGjWIZ8TjxYbPWdIklz7Ddal8FJpS+Kof3IlRnSnQvQYxBASqiIwBprirV/CIT
tyrAFAVfsyUxmpoeBZSbYKkIfWrfI9r8qRW33t0bSu5ge08vldcDR7G5Zg7nhEj6nnjUkmAXSgPA
JYNByTFa0h0w3yVVQQCQKBIQBNL1dBVhL59VIPwkrk2uPuEbGR7re7xW7wYknl/VOmA/FtjPalRf
pr4AF/33iujUYT9JHLoB/l6oPa4ChovYqLAPP0nDrqGkYXmT3ZR8MN+0HAQS2IX/bCPLkCM7tYVE
IwYC2ccrHiVtKL7w/ByDwpfu+onzUDNnbIVWlTvILZBi3O5h/uvpbynoOoD4YejCIxDNl1Uc8Mz1
Xg/qLQGzoVcT53W1HyY6L6trrRcCIUfssIdU7UpUrcWDR2YCG4GFOA9w/0qOegUB3LElJ9YxfN5A
VpDTYanIrpcpA158GBttS+80LhTSaxXRwHomXcyhOfaSW+qfoFywZnAZ+3IS4sTk4dy5TEiLVTmk
I2DGZ/qc90RvM4NJmJ/xInCDL3Nwi9t5BjRt8YKGPFSz4ZMS/sIRkC5rFM/v3/yxYIlgM5hfve63
uyFc99o3PFzfuuLXFe6xNLs/8GAinmVBIn6D8v7VZu/LVAwA6Y8nkyKnf3WjtlaFU8tLVaQlR60/
g8eNLCnp2tlUBgEIZFwp2LgcV6Ro+yMg11oacGELuppYx+pbj8fm8i+llO91U7fchuIusejaebk/
ovnI0ZkWU1uQq2GTdB1jNS2UW1QKtKYCrsxpPFmp0s/3kBsmZTS1is1Ub1bDAjM/wNbSguA/QPWK
zUdJb95M14DTi3a/RvqSGldSGDXLVn7ygfT7lEI5z3AmRQic6lu4RKETmT1qJrrwMknvp1MLxJZ4
WzH5FdoyzqLN4wV9yOWpC9iTVH7h7NAOaWQOjZEA0qYcVU5FuWZKXJkvo1naRe+UgbtHMSFDAXPX
idS5aXzkHop+zrYjIb8YxAEK3k/ULCLl1cd5Q/X2vvorriq+y2uPTH4hjecoIqElAiU+Zhnz5biv
k+aKHny8jjQ+IzjFse+1czLbl5pREv7zSIG3cyecBjVDtwoEDELe/XByW6z4UBrOfpip8S6wZiQw
gANgOQvs5QXeNy30ct/kZaQxk+mHK4eVJ6KBQAAKDVX/DnRyzBuRdQJTv3GMSR2K7j3rgzLAhRPO
AwGDNLEo6oI1+Jenx6J781sM5CpYnlPBHvy8QnUOLXHlUQgc48VqdHjEwEosz0TwlU+G55u02Due
VQoslfnJcC0MPxqOpkXO5lxsjQWvLG+QiBluBfU//kL+oGHkVTI/slAmjAOsYJFAvNOaABCVf2PM
p144DGPsGvtOZsHwNurQdRcL7nF8l375i3DLxvEtnkubWJbU6TIqgCHodGwW2+UfUxtgnE+NKKhC
uq/ztWKFembsyS7jwFVkDSLwOU+pvgQWLqfcLC+dJp68iWLcuY0MgowC3/VSzJ8CPmmx/Q9TBvvB
MmONymGpQ9HjgfZ4/OKEBaC8SfTf0CEpJb/6OnX6438gji1Pz6G75i6M0MAgG5BwupukgTZDuVFp
wGCsehCqgZ334s6DJgrPzpi5r28ga6pwFqx+bwifd+mTo4SiADPZAPJAoR0bK5y8CzNXor9SNWxU
+2yzQWujBubhBZjYwo1RCHuiPKFMJc4vIw4Op3wa6oUgOvOsCTx8yTVbEHRmzDpSy/Ew4CadKo6s
upWnmawXDnnEu2KwgX3H6BfBXlNzoVCTu/EF0G9gHJopQ8ilxsc2KglTQPpC2aRoH08dmyLJlXmr
Sc6hErSNUq9x9JOXfzo4sYG64wPgAej2XYMY9qsBAWQMCKpMD3gbVZ+lDIrrtt4SMVCrnn/b71qL
8gHp5R+TC6YII+CyCZ9411857JuL0cjnOhdX0+umBAdtKJcokOYZBiXqN5c/6oGTvEuihmnIWwkm
tT8wJtuvPkjWZdM0mnmeXEsNBBkAI3W/1Ep0Yy7SPq0xvPAztHp1Z4zCsTc/fBCY2etO7S7zPNvr
RVB4zuc/R+fo6XotSkbgI1mLc0EXlXB1rBEHUeONS+9M6coLMuz0J+/m1w8ob6Wvn+tU9A465IKq
nmHNusbft8DeyfsDUsR7a8MP1PUAlsjf1MrUUaLM7gpDTqU7YmuuKSA9XgUlMxbEPIwMzzEvDpVw
TFnGb3jIp+RUoPpBk0bt5/AoNI53wSrK/+uko75BeEMYiS5Bqgq6D3QwBfNxzD+t6jm+G99eDg+t
eKUtfXWUYLzrnmaVE4ogoTIUTpgzpFGcsSgz4XixKd1Duzax6bp5Q9euespGd7uY/82UjzChjhYS
XCK/7z1ReYUFPMu+ZhFQSGhztY2SbDuhVNsJsDb4vxlBagJM9TgcR5qYaXGZEmfnHrs88rOphtcR
Op6gtvhjPrK5LuE4eGKHcCojo5JeE83/jFJpli7rJsU5nPATCDC8TTW+wBc7RocZU+5/U/0nAhmY
k0phC4T4YVc0uSc1V8xv2RoGwR8x775ZQRBMXRXUCHxUkjx4toLiopOvwdYnLFbCwuJUu6E/8dp4
F2VF1i2vbTSRvctiLybQiZf2xVSLR0qxud4lWlg240fpHTgV+6NFDfBsxpfx5uml8SJeKoky1b+t
rQeR4CMY8zjnshhQ+hEZCSiq+t4aXC0h4eY9dE0HAisomGeGZTBl3hXaqP0KWQKqHCPXPBdWEuPi
Vm7WCZSjJCzInnZh5W4Kb1HemIcWpcBrM/K5c3wOpA76Zcwxe7EP+MXEAMu9joz8Vcuj92axFFZT
HJR2Kw9pupbq3X/1WrtO/AEWvk9f0A+0TakYOKBBo4+h47xC4mpUbgOftBQh5xbjHtHMpxQaKnWw
wgg5/VWGOSsk48p8Ancfnniui37RCcDABkG0LI0ddr8bwb5wcpueAepAMy4eb4ISQwHMOimCLYp/
jxbof8g4y9z8YRqI9OQwqXtG8uZ89pMf4ksO61VdP5bNc91SbZ9ZtJb+dn/8PGdpl8dDB3+22PKB
YhAIHVacqrGO9OECRzqgY8ddak2uf5E9jYNzgLzxo+T8Wnc2CN9meVVSSQ47A3J6sNkIdtaAKu1G
5gCQqfHW8eReX9eRw1IKOfy2n1rsbH7xYivYn+DjL7RcOlTcIAb/vT6+X5UxhxBamnET4BAXIiw9
0IgP6yHp+y4WD+p4PWoGben+78B0MDTohNijeGwzB9q1fXm6tnpzMdLeEh3XZUOLLzu1yNYsN2SV
IyOT4M5akdPmbUNpLK+epT5EinGIIMbOqAOuSithhED55L1ujgLde4EyW95v0KiTVV5JQYlJhTUm
86yiast3NODqoEMaByKVyeGL3VQ/hUBLiFc8IxJ2G1d8khs3vs91o5z1qIR8fhaI7fly0zHi6c63
Scvz/z2F5KbIp9jKfX/90auqviSpdSe8AWmmt9HvLh8qwYYW+gDZlxd9v0gETD3e8hxDbqs/RGEG
1G8VDgxTI7OvL8jva3S7ertHR/nj1wLg57YfAR8eUtvh+CgGGSsmTmklKPe5sZ4TEg8KbtPqAwg5
sMW2KN8jkEE72LFBuDCJEPPWpR6G8JK5C3lrHTGqWaOq+MINOsbkKb/ALgwZra5tgoO5W1VTziLC
TNEtXAOaG88mdQLErkJ1JMMr/lWjsxDgHzGtAwyJa1WvCkU4eUIShYG5QxN0+zlwmQGHVXHqinSm
5ozt7iD9vQYHXLaYntvbcL0S9VmWqXMKTUefIdzw2+1Pdd7U0z83Rdhu/9FzFad9XX6pyuWLZaTG
ayOUNjJLlspLIKqwPxJufpk9NfaJXsJqLmpgf4T2exFGIqa0/4jw1KrPb9fcLltTCElnLTJXizNw
IHSuO6hSv0F+6P0JwPwofL1gL9r560tP7Ljb4pgcqaaeYZQDbJD3BTQAQ+9LLxckW9eBTnq3szym
lhitWUf89nhlHpwVdjWjydv+vl+6KX3BeWimrX5XtmmGPjdJHXfT52QXXE+408tch+e9XXj0r7wh
VMQz6qyi5Z7tRjtd+RUfhrlU8KC/XlGpkFUVijOHFzD6UReczdazrVCaGMN2eeX3ugTj2YYI4AQ5
bHmVXAwu9fvKBVjE4Vs4Kt65R+W+IC18osvi9kDt9MErRAcZ/ZBRV7QtE+PvDUOZ4KKPTRn3FHGf
yQ3uJc0qdDJ42vPDI5ALNpEGpazL0vk8xu86Fzs6Hjsc+VZ9TR97TVFnsFU4/jCn67kib4QauUMS
NMqe6PTNlZZcCmVTbHV7IpOiJat3wYBqF9AGxb298yfb5IKYuwRB1w3OhbYm/ds1GO/KeBalIovJ
iAJumcCXg8RHZ9SGAZH1J6g02xxOmI/KoyQZBjUnP3JZxvm72cX9FZr6GVKk8dc5ZnI8M4/o55ZD
0fkAEV6FJCbftEuO+lcmj0bIQMopcxhu5lW1I2milfwtFK6bBl2cJ7GxPAlxxjFbnXSfPq9B1QQf
bcYybg2DzBfVuiWBOrcXms/DsCM7fEu0AJ/Nidc4MUIP4gm6kQdP8gusCDF7Sc92kF2iX37J3Cw7
fS6jGfwkXz6PGBXDPEFXqNKvex/WYgvNOV4DihPzHWzXkSGttV4RoqX1ChQJtZ35F9kmySNdwwK4
GY+eXa/Y/QcQ9Ib+m224ZyJydSQBqGBvLVx//yR68uXjEB5y6IGwdYyyh6xb+j9iPPXr0s/pEGn0
o/CSuNbenSztvbIS9V3k/K1ae1K3FubwRMQn3xPxt8U0XjF+AfAq4ofS7X+Eqa9hdzC+KnoOzh/2
7+TvnfUPC/YgIyNkkEori0M7+CTvr0koLnGzseUONsVoJARiRJzWToh3MdkSYEkGHQwxXc4ikUFX
rmyJBqkmbb0yBcg1LfTDcNQIMlWqrMSQeHKMJX4g136GnO9fhjrMhxpxPXaRH0BaFXlf7q86RQ2b
7MBqQ3H+OnzRpDLLiaTjf146mRfRSj3YW/SkHKZ8q135FE+6bCsAdML46PeUpe6Wcuk7UGqN1A4O
q61qbF+bXVdKtmEyCKFRflWEW3NoedCPGcbf33EbAMQBQSsF1zR0KudtPspSd7BfCVwr5GAo1RRU
DCB7WS8WLDxrdz/H2y+Ms4ClMDwpaEOkVwWIeNd4rVYHRYFOMH2HaDjT6bKNAHRzlgTAoGk8gwQ2
YH2BFBu7s1JmUTuZo26f7KjZ34VG4rVzOoOHihSyY+D9j+2EFrCa+VRza7gQMzE1PfTu0+0n1jMT
41X026iKvH5UcrSup458SPs/uIvvC1vcSjilt3rqwDfxwo5OBXCevEvS/ClXrGCO9Rptk1QoWU1I
9w8ByfvmjbdYAsTTs54MwMjAVNjyc6SKw+T84j7eX/fKzbrC01PUwL8voxc8E4ZLEZJ/DJ1j5bR6
2K9XlqMaOcjw4ndsHa1AlBe9jWtWtr7AK3NUDbF4srkmkVDdLW+4sDpCeKhb0pj/Xy0QEE2mCPl0
sjGXm6R/zy0MrYqXS7O63wOAZOkEBE77qcrf+4xVyXq6olhmy4mu7yW2jQanKQz24oeXkF7yXFXd
SVKo3VYzesmfPW4cV5Kg0gZz42F3qKTIJky3vlqnVbLhKEUlu+jI7r/eJ+baVHXB3DvH1+9DhE/P
qDXNsxoltGnjJkXzbPTpfKITrgnntCo3jazn+UTp3YySMsMt8s5SSfju0MKuRB7R0XrCC7b/I3nS
t4AYzT5VxqPZ+pUw24lBKzU5UI6tNgvID46wsKuAdetO4OEJwUmC3JRCTob2lopZv0LqXZL8r+o0
tBOFLfpniN4SCrg4NVX+cQuWS17S6aDblcsDtY634SnDgC8y5QHVK9rAQ7crZOY2Gqij3H1L47gJ
Kuh9TfgMNaZRC8xvOU25MNVjn/FeiVXH6Pff41R2JxHckgdsKOssRc1qHibxI+07Wc1xB1LBsDt0
csRHu8Jr+PfPmHqN6AjOP4Tuasv3muTrka4rDYDhpvq5mML0DdQy1EbUrMpxexJywxxlFH64pz4N
Z6cDwja/y8BmK/bAHlZ769yhk/bkZ3EjOjbZO3Vy+K6uwjMBOAqdzFWiE0uFeKcBvY/OvUB26s0H
RnJr1GXwaQTY0rjPeJvanAPtIudzpt/NpK1GbmTb862yDvvhl4Wes8I+Xu0VSAvsYPrcQhSy1kGH
NnDkvndqoOau0JnNLtQok0GzbhuEpnWaj+QjYKg1Gg/Wk0IVpL1vqGBk1x2SovMTsqV/7ycxIAGf
MlQd0rwnkA7x5lSPKsysMuECo+3OxC7bbAH7zT18FTD5zY+e52dPd1wDnRdzGwaCKDyMUELTrP+x
11eLyFVxkwm/B0lB0fxyRGlqSY9k0i9WBB8zN+glRZ1nLX6YwkoXbngL2+NOVgmXWNUHbjWO0qc3
aosow129/AV9rxSyQ/Xdk+EnVzJ7Nt9J4F/lL381oz0wP6hwS88RghPZKpQv5Bnss8eU6HiSU1I4
SAwZMEXw6BTBKDqHORUPaSbxCAd7JpAxUP8nml71jtyVDwISprF6/ytHnqx0qrkRdKr9egyVv2Rr
/eYM6Cg34QCuyAIn13BQiFjh7iHI7OEzfdowMuXX+OpqOk2KolhD9SSvF3T3/08A4mEZQO792dro
cXR6bTHjyshzSsmegGjzlN9V42VPV/AOjo01jQ0QEFW9s6mHCPRqpissoRt43QNFUIyXDN7L/GUY
CPHesEU51aOCapH3mjcXv3V52rXB17ZrxHQiHP79o05yO/bLutzpBc4ahcLpAKfks0Eeo2gTuA8D
YlkBiFBYpMkcjrgADV/VRlrKBpzRfN4YzKm0zNw3BnXkWb4y0SpIJ5xcwRtXeUNmw4bOtUfOEJmo
zp3QBoytZ9pR/n90fmpQq4GQd2tmfBuoPv0kRvd7ogOUZmuGzYEPv3PHkBn2Up0rL9k43e3dtRvx
UrV2ke0wMJj6FTE63BS28YekfpG1cO5r4ifGamyg+ZSw7tYGv+zyqZWct2lItA2qbtHX9AXjrd6M
xnqWvLBVcKTos1MQAWI10quPE/Jb4zLb5jG3N8x3gCkQRhe+xan/i7zgCTLtbqS99Dw7rq9N/vsk
A/yKOHXqGipwdeh1AhHK+dvhtt0EEUSIWXnKgIT/1T+cWyPGqYF57lhnNktE0i+D2AgZi2/18jzm
fNXwo2huBHiFVrSeduuvpr8DhQdAxX4Bduevfe6jC4Zb/ZZ1ugFevgYf8cJxsHi/TXguF9bTi82c
/KqMBH5MQA0W4bPs20fNy1aTQ2TZOr2IGt9HaDrdZumLNw2ro2eWH+rLSc8Kmx6h6D7HOlf6youD
Znm2rr3UuUYCgMdi1CPpZlR5QffvmRO533lRl/+mcbyu4fcwT5rQlKzkab/ji13k+wZjlq7ewCQo
CdY8rs3hQabI6X7KA7s4BxEXt7LNJv44JNlJq0rvnEcgrP4B6YEgPlpFaZ245pUrcLmMBHsi8zae
XhS0SuY5OlU4rgIsqfH5BahoyGABg/fKx5yUFs+ozjcFfH91FJNa2BqAQ2cAu6pnzu3kSesc2LgA
qdXLzy2fZULbkI/f1zIBr37sJHXYTIy0bsCVQ+3MOc8DaotBpG8FioLTXsBK4LfyShWrO4BFXeim
AvoXYPcV8UQOsIu+MEmVEPwd+0GjLZgUkCoFpyyG0rxgPyuymGvpN5Wmmmgngo/YkI8nq1bQnvuz
9XTZhaTfEuGCwtnQwpl4Kz71se7bHBu6uOTt88T/7oSjQSJWUMU0L1z1zuD4fbf6A5aPJWWsJkkJ
QKhiPw/LJFJ/eQ/huJNZ/IRpup5eVGfbm8bJYW5txSPWkE9lbNynaLwyS0RQqCsHlFrPiRLa72Sk
p3+AKbRV4XALRvTOZyhnZUKek68VLe4x3KJK7pKD6fCqlDncvUu1KsBMeKFkWEkOi6wehSalY2C/
7celrWiEhuwvsdrvpkc8rDk3unrrQy8ofBMhcm3lXB0VO5SNTJ/CgeQjN3bEgKHK4MfuNSvGJGLi
4XhG3A2fSrGuBAzUmdke7pn17kbf0H+6LBDBCBOE3gXz8NcJfP2U0osfF5gcpP+pxR+io76EFpSo
3gWng4wZTsoy7dtswdNRlc1+51NjhrGRGuyiWxSDF+UG4IwCEehABBWjAHUrQcr2bsNO1m1v8AJP
Q41fJ0NjuPeGrlV7XJTukURJxvaUO4+10cif9wPYjJX5xl5pPbijx1sD0v9qrwAAU9mcfr1LiA2G
U9v7MSyd/e1v8ng5meQ/28Cpg5YpHOm3Th4me1q9Wf0z+BQrpJk0Uwi8a08uQR1hjz42POMUQeBX
+G/UgOf+2J3J/xzHLYPn0OJsZxVukYTh3K6PwDNjQQOqI3plv6aOzcrtTGp+ZiH+WmvWUhdbJZU6
i6xA72Y7U6J9TcyRDV33s335WmWCgSunBy03WUp8ef3fncVlidfBVvxHwrlsju+Xby8j1QDSLDLh
pMlgMu3ujSSnQ6heDSm+J83sv7+xaU4buQwZj7tYa0JINaigl1/gqiiU4mng5FJasaivsU/QsbUS
JvOhFIjd+BW4EuqUe1PdraXTWd92NYyshBry2/7jpJ87gr2vOxIMwwkmK4zEDQG/oWMNXHBchvrI
YxuQJpnnxsRY32m0XuulW94intYczyPPG50JnHxPVPXD+fxkSJBIFnjAloyWKAggEcfK4DzyH+Xk
oeZiAEKaKFCFTPxNjwX8+NAlJ7TP9sfszpsqrOdZix4uFLRQEZR4oODS43p+jSnP1Z/v9csi7Mcc
Vo5VJIcml0XTETcVa4LkMxbNHQf0R5VdIBzIdqOMck6iQAVt9OKg8fWK9fTiQDLsBgKIU6sje6A/
7IgnpfFB+Fu0oZO/I3ktl4sUNw6vBait7I14sAlPuS6wml/kZv8mwRwk11t20JT2ivCVmvbK/mPG
CUWTorOQmtHHQRPau+zqI+VAjAY8g9rs+5FhvDe5zsvVP+YQQG1xYOgeBcBTmXtTbgVC9k75TJOJ
CyzcbQwYwb1E8kWmShScDAzXpkPV/lANWLg0FIwdCoR1bojjx639parM0yjYXAyOzyrffNyBFNol
4rqLZQ9szeTBhBD1KqupEte/UL+4K5jwmDZUrjaPJFde/1VSXhCjiP5FhYrPZU5dDOW0XI6tJNci
jgjh7MdZirpTAwX5agMCywFp8aTNqTfqgkvAyH7OtqJxU66hPuwighLqNJk7TiYdPXW/+sKXtGkF
k72zf/3I7eQCM4gfQQH0t4KtqLEpumJWMA1P8hLUj7qkgkvxObN8fsWShU6OkHR0OqtY1QWDRDDD
vkMFPHHbqvNFLz46DHwVhcZgDJVv3VeOb8jt8lDr1ZHirS/lhMrjGl6Dv6Isqqj8Ndq2QsUm/vkw
3Ep0bM49Hd0i6rU8vaSisgFtiMedntvfQw57uKTFXRZy+3Q25aOEEDZHA5o2S6w5BLaHHy1sAuS+
L4SetbqgelmM1lGdh4kuuD45buqe+ASJQPcGL97CGosqyMlY+bGdjDQVlEMJrekZqkWGRvF47JsV
xjD4GnCeMj6YiPL/atR3htQ1w/GUeoAl742vWghP5xGAmePHhJQuGWqkmUZgOPg9IUaOM//P1DjA
j8LAJB5Z7tOB7Yr+A/IT8/14iip8IR2xnEjWBl3ELRrJtIZX9mKdeTciqGPiAfyGyOgGJz4ujwI5
YuDS/gi1u4tODm/nBo1yfw8BR9LXmUxylHHTcftsQpgw6iPufxhYMa20PC8NrMGG0Ho7aGS4SFKG
E6W4JvQJen/nYIrsBYDpY9kgz0l31Q/VzT3omiV0H6cfBDdMsyHcsHbaTI3PDnlx2H4C+07C5KbH
Aky3PsbCysEHGgxTTyn/8gkuz7XR1kRBEOkicFAyffOCsNe1AEJZn36/Wq0+Agq2eWZmesi6wURg
w0AVWAjOuBs3/rV9mMcscnHUnlROqdsRPWjJjJ3PUl1hzMqXzQxoNrfp4Vkg4aFL4FCiw4etNZbZ
IRpKNiwKObW0lZinyMrAKpHi/LtKQGDs2kWzhC+jM7yH2KGSTZQ6s+FinY2lHZ8Ng5gkZwZWd6/l
4+xPiRp77KXWGmnG9eN5yO+/WCR5mIcjrGcbXyjPSc23BhrePN5qbUHogQ/iN1zdH/60fP9U3NZq
gRmfilg9zLopA02aJBT4zsdZ5lXmcf7v9rQ6PFYxJ1bhCokkwMt0WSq95/UV5vHwa6si2CFwT+ak
W8ulqVKkJXHWxVoLK4iIgymEA2G8wgV/KjLWeO5cGkeB4zZ8SD9VoJXVjB2sguRpaCu27g/zJeJR
6Ixhjtv9JTMlLTOhy2NYQ0Jh3qYdaW509eKWCHDw1kJDDNqpINCDt1k+8NDNySvjsgXNzNOAmzcJ
UMMnEg9GyBrS9tsSLBBUUCHXykJwJI4WvXvOeMpffF1CTqAk/1zK8ORxqqgErtiFlcZTLRwU6wCP
fGhn2DGZQW2cvrowo/PJfN1uCOv4BpR6CJO6Z0Iz170XAZOKjq6XwI8csqhillYud9aLthLJG6HM
5xft4h8GCKgzFrbtNmasIFJy8FVsVgHfhMMcJ3Nh0VOSJyXohDcs0/b3LPLeBb7UPpzanVn9ALFn
+9HqAa8zneLnJuplv5pwwPNlxg3km1x5TuYbGmcsC0Wgtga6Jocs19RBj45G7EnwvOLuzuYbxzdO
WqjFVAxIDtsrZiwiVAywGIjATOZ2pU+iMyvN+BNFOsHDsCF913cLVbRs+hul72lsaVDk2Tjvoigv
+BmMX+zDyIHL7y5mKYVbTkj6UpLaAWpw1MQLMHWGuUmBSCzNRiVfo1IVNm3pvPCNQHxh9/d9Y9JV
mCVYZocf2B6xvFqhe0P+1OfGSTc8rKsS2DeVTosqtNS6Zez8ia5Q5T55tVpXPXYs1CjlbMeb12BH
epXrAflxC8XrUpmciunwUcFIz1u9WtlN0B+DRF0eRxusMQLAIdHcPZW2Wpx8WWDDjBKse0jpEO2E
PZWX0vhI7imdrtMpS/mP/9PKrI7rL8yALfujkUOIPTtFumKIffiBLmbJ+JiIUnw81w11S2wX8FPZ
W4HqLeFFVjfjZUVGCLOqtlGo/OaCzpjjVjAWPuZGwQPM6wTA9fX7cqv+filYxIVB0jzJFBFFpb2n
0e9hjnmXmwYqoSth2HvngVkp+FuOkuY5f38K3bWe/4Of1c09fGxUF/Y52jtO6sYkfU8fJhRYtUqa
EiMMIHFqddFImLugBYvG4iv3FIkmP8e8MwjhtxhJtAaIPDyS5h5tLBcWewZlvraZbPe62+9YuW4M
BDfipRhwncSyTctVhPJojgBPNz1/d/X6DF+TmkdbuJ5t6MiDKkC13vz85W37KpWfdVBmgrErCptR
fBc3iz2Js+rseYRGyzrKi8mB32ruXvy47ar3V1Ua0rnFEjsPr6TtPCZ2JUZc2msA8cGxgwJXq/Ng
WADsQlSMmeouoEC/v5ESzII4s3n+jHik3QhZWM0LAZd1jvY8E9JIYJ9AEh7zQkO2As/rzkQXC3wX
keEIStRyrqFZe0hlIuSg7qfxxN4wvkPAYPn6q+RQYxxE2rCmQAFdF7Fo61kmI5TFfKXUfOiQQA0z
XjykbaWe8WxF3Fdl7dkQ4xj1LDuSGfpZv/HWD5UXC4eAPJZnnodleevL6jAt8bb+aoaTWKG2t6B7
GHLLE67ls/NOVsKhkU4XeYH5MIpSHhmqKdxqgArjx4SP2HerR2DR9iedweL4HFsBpBtgsexbJQrc
5tfK2nngNzh8wohdtmr9fqxJY+yb6P546I9Xc4UAfc+VA+rywF70mEtipBPx5QYhBz7pq+9zmvPw
D5Jbi3oaLuq4jQbs75OUcXiZ1lA962kfYlrof4ft02d+78ZZfpgxLhabCUbKYJxWxl/NFHa3wCht
be7FQVLwHVTp1LUKLZ6dsgI79Rix1hn+hD4NMEBSXQ0hufG5BYbaHEKNG3oUmMR0BYI33et/b5hb
A7sALMQsa+O4dT23X8GXCsnbxDQtIROK5Q0k2w+GJotJFIBzdCtbZ5ZeMQSqzqyXTAZY0rTnxCfk
SwnVXZ/EAWWNDXsdX+v1fwpY4g6rjAYjtVW9LUzYOJrTOeXHU0NuA5JQXrkrB+fOxaHd4o/uwA6A
CZBFCAN4WWrM8GT24zJiPSu6mUOpkcJ6jpnrplneX8cYvVE9HaXgMzjSNEF9Pi3lkdTYAc7tRXDa
2+q2GXKKqwjp4KRGL0jUcssCGyCZw4/7v+r76I4bvpfJflGR+zBDJI21vEa62/4fWeSSwporDzl5
+VeFG1jpWBVbEqQXlUaCoT9Juq64vA+Kz0v6ce5I3NxCjqvbIzNR/iaVz8pxzu+XLpptNOEvHqz7
wdkJZvRSte3nT5/WVGyyIZG2j+0QtHLfJNn2P2HGsbs+u1cYgFwc8OXQ2GveGNmFJRoJ2jHcyMsy
LJkm/lSpJucKxduuZL7jGvS1NNijfJdcXlEhJnqBS5kWPpiodOQoa92XB9Drq8nXtEH8m7vL4O2X
RSjytAiTail6elmd/W2KaHC2oUdNUzkQ/4kAc72kDGZI+SicSwDL/DEWFsewGdEl2RORAX+sA+Cg
Vu5+zZM+/Tn3QIukZRzrAXAzlm0SolMBn/xlQB73ECEySHgBZbaitTw71xR5SyN8ealyNAie58MK
KRDdgwIZXyb+FgBAkHSV7cStfWi/51JWJAAgFT2XwKJhqaomtO7bgi9Im/mYJD+UtdXC5F7i9bcA
k0z4G2XuIumuaxxfGbqcdhnB8aSfQVumMNV8JwieSD2h5uqB+MHesqMfJSoZAATxPA0Ud/xOsVkD
tLgxMFm9Ovaq1Ssf9L22jLBhW2w/UjTkyE+N4WLLtwqEBF0g82ZptZ6eOlUBcWOhXM8jDqDQ5hl2
esAfDGs/dV08fHrerANIGVejYKvAM8yK8zRT5YN3DfWjXvywkyZCz2m1govU0N//mH2KE82mXkH1
0zA8lmalAGkQswXGK5N7gO7C1FutQGtoM78zZpIrF5LaXWCdNErzwgpiMiSd7xMCPE3SqQ0jogHR
gRsFVyjGP22IAaWIdYc8FCGsgeUsgLCygTzCfgBIzQUPs7GuzhWiYdzTBD9gstxWt6rh6mYSEh+B
0hvGRfsZoadttqSlS0cWlOqFU7R7Fp9DVEaIi8vcAMWvuZxVXhWLe53KrlU15Za2dIR0fsombXh6
jYmSdTYu4X3zPZyCROH84NXMkoI05Rrw+bmkMtHsWb+gQBMFn6Swz7HvbQo6aH6B2OVSIXBv/v5/
mOZNrzNnrtwAZl2e6pXWTkAeMe/6Em6oxGPmic3trRwuRkotWFm4GD0glvjQ11SGd1YWQ8jxJKVu
1eJ0gKW8PTFR9G8d/D334CTaSB4U3bH6pNDgfs+fkTMqFMp10wuaentHtPi6GFLOjfijLFZCjRzK
ztCoIwmr6dz+re0BMTt7SXEKd1qn4Y/COyjctDPBYTnS+0/KqrkU+4OtPxw4UMKYJqn+5Mjiy6zn
7RRYeO3UDViM6Le6V5MY7QOnicuUUYGtbcnT2yxMwTwS2KzMDeZ/jqau8c0hIviuVSeyEVCj0Ob0
vASbdxP+EdLd59ii8meto92rnd0+rsUvNqPeaFFjsIqRRZtzw5Qz3a1rMsoB8RlhD+JVecXtuCBj
KRuA/9AQFNB5EtbvZo0pWLIEa3rVCvIRiF+xOilywPePDqD3IUzRDepb11V7YAq1Bb6ndpPjhHdS
MlioGgWpy5QFioTNuqKbuEw5tC4oCDDklYkKFG9K21qHsecgqfGND7FePnmXJpqRcc8OPX4A0gfX
CS5+W1ha+zXAS5fP6Q/9x64pXa49tl9jWXwIqCa7mHKPlOcp79wKSZdo712F2vLXrO+qpfH0zODA
8rwqH509RY0dJnXrOzK3dNM3DlSTcZtVcZxgGQSzGpnIPQzrVzq7IPiIM62SwBoa2ayrwEiAQRBs
A2jz9X9SqOWsqV835y4ujLuUIHWOUH3LNyq8HAsUcplOIut8VEYtfgyJcg50RT/zCiFM4XrvI2l3
fgx19OAxCPsRad6vVABSVmrhueVQuC3dy4E01RanlAVmEiSWf4g1NOvRrnZgnxZydNP9L5AmUtLq
RjaljlaDg9icoRXeBIzgoLXBVh9wVer9NxLX/8jKEfSiMORr5gNe7lik4RWg2qvYSnsQwehol8kP
jSqwoNyvDG/RZJDm0wq+hnmAH2AbiUbNdDoi8NEitccvNYImYndfe7IO73GpMI3VbF6CAvXKoDFu
KKFgWJbnhpCSuqCvb894IM1ldWyDPiWqMO4/rxYnfNQ7Yn2ALr9UglK6RUKoAiCgD7j+60qcaYoM
2Qa/ueaf2mTFqk4hUVR1gYPJsayTJNXIMQlo66BOmoOI5UkppGO76xHJoMZzA70kvKqA+Dhvv53E
1evuSciBpU+T7WtZhgEg3mkc+np16HDnE70RjJnba2+3FMh2H7wW8ktGxp8SVNOQP+XWyM857H/b
PryDR3v5qU2cCDwTwyNz8Mtk80AvLCg8mvffF/wg4aMwnAq6katby+5F+3lpivm05m8xsKcEpCty
Obr9PBxJmT+3Rs/8XlOpuOFsi3XRYTFdP6WIo/R99HtKHwy8o5+Zr7yayWsNeS+idXjuT1QDs7fw
BTjdaPs5LuVSyEEw6Rqdgw4RkTNgsAtbkmNDdwDshnEEWWclxw9TlCxXoHIBy795GgjQDnjehZa0
rLjUWe+iSbP4Rvc1yUU4pMu0kGiNGIprrdvrQ4ozjCfAjILPNdhFvIUY0ZQnXxYCdwm2dvgAUx/l
qmPtAhxKbMhNmymcA655gxMLf/KH11/0ZQ4ar/h13aJqETRDfldK3CVzYBU/O3q9/K3BJOU2S/MR
Io7qEBGSW/rQmIyoBB94vIsV6FWZW2Q3gyBMqRXsA6RUKXNMiNWFrO1BLqMxeA1FoKb9F/TSbvpy
SDrfwXAjrdkrZJKGwXKfv9AeY4v5jzgm+v9e7n1c8+06lVW8F2+ro9dtL8SU9eTEwG/AIUw1OWR6
0hySslRpjgd5XzMqX1z8dJyqGEbFfknNBJtC+n429T7leaOgzOq8yPuyI/E/7tvpuAoK/FXfz0gf
Bbt5kLMsmp/GR5Ki1JjNVL14pSd9KbBWiJ27IwnbQHm00Xc7e7+dtEgBUZ6bZYYFi5LAvdFOwtV9
4jPj6U8nObHTUlG8rAEWNVw0ic69KUSa3rXs65GO804l12KcFv0LBOgM0SRK5UdCDYluyYv8QkMV
w2/mUbgkimZHRGI77LCq4k9h/DaKXU6lJWsGYoBuPPvNOKDHdJgQIs9BwOQtR9ZVsABzawl+rbAs
KyHD3Y+74Jd0J4nV9rL2Q3iTkF4CwboX7G1P/EPXjF477CQEDEo9IO5b1adI1We0dP1lIzIyXZXJ
eIhyZC1O0OSZi547B54Fae6LXdoItbXXmzn0HlPGrCB0ih7GnOsQGP/0WskAXDHw09GbckUvy87d
6HO5xu09KGHyR/uMdv57zhVMx1uLyeh+0p1iYEpyNUy7UDXGixvAhiN/xBaL7y+3yuWaSCyeN0BU
WBEwvXpuZB7tIaEv5xJWU6pRrCkbD9C3Z2IrperoiAfyHIqXaqOtf03ktOVujmUSU0k1CA96eCjN
UzqBjI54bq2O40ZD5AHHYNgiG6M+iJC8tZM8HvZUqacd01sEkUnkqdgY0wi6lGD2kX9O7Ih/dvM0
K+Qsti6xhZWpwvBe11na5miBQTj2P0fiT9YKwScGSdS9PkLKOng5/6Ab7ESyGLV9jERyclLoJbx9
2PGq+vV7ZsI4YW3DX9jsvZWQQnHt+MsHD3KY9JnBlYE4j6OiHt+y77hEmo/tKb0T9FT9ZwpbsTW7
4r5U6XWk003Kz9sNSOGg5HTh0rR/LCJMYixaA/mTnGgJKborsOKiyXxHRGK9dYzjL7sokhSz6l6R
Y/mkDwa+LzlIF8ZHsDxhOR/plstIP/yXm50EcRD88sLJxJCSRcNkkYbSWPMjtq62J9x/+3a/lokD
o2HAS/nIyt0HkvTi7XigWpiRjgtr6ZyMzvipztTZWGNjXrCyWRsZIpLcXC/AcNcmR/3d813feiLp
fKKw0K60/wPTO0/DWs/CnIuxgNWm24nzFZ/L0YzjMMwdiUgc9ZcPn+iCyf0kajTaNNib3Bs6aXY1
lyR1YpeLF37YyV2t/yT4h3dOfi44sKRCn/s7Q+xqFyJdsXjl7JzCKI0tagLWeheipP6lmqk+nHXm
82YrhH74XR8b44FvW5vu7bcbBGbyYvNwJZuJWx4Hx8kUqOAiiHN/W3OqlLQlgcKDffhdf761MJ9G
xuLuFIOvtyU3r1UVA1wmwpJ4YuCQp/vY9sLgbm8ptbpA5FXAt39RLNAu7GwaXnBi28TOkIems5kE
9iu2BxrOYD0byR4S3DKZPMHbpuSljjqrMVOZ7W3G6X6HAqeSKPbbEkzDdq4g8fmOnvr3K+uaEMgP
8hJJvs/6H6ONL9mP6gQf5DpamovU2L/uu4BH9ulgk+uzS1UUrh9sshejnVyOchd8jWmVY6vRk7zq
t01O4XtPidDxz7bPI0GYh3UWWEVz+y3ikROxJ/l/4tvBX7yT/SdgViipygxEKWtRkUUHsY6ufcPH
bTxgId+Osm+H7GFvkB9YIEH4vGtLGQoAfZJjxdzjYRjZNDXsru0U7QsA5Z19ihWMbcyPyuZqr2Gk
xb4Lw4kavFXgqGo6VuhaHuLM7JivWlhS1jVzlgm8J+lZbdOUnU5mUdEfppQgvk1XU8or/5jeTov7
3bFcqTxRd7y+9feFsm4GE3I3ZB1Vf94+xuAzSGSixfNKZwrU08NO1Ldi7CaUcQNcPxZ+wHm8SFdC
iDyDcyo5zQJdT/DWc07DRLCH6mRypfBUdu1oeGxloHzVGkZTxKHbMRcksi/m83KauOlqqsazFYRk
H3jlu+Zs4ynHr28P4MGbY48HRkvXjLnpdYUNajt1vmqVLeoPOswgf9VKwE03W0RaGqaaOQkizkz2
9jCUhAW5vJCWrRXfzvMccP5RB1KB+x6UoZ1+XBTvttXytZJqSQPndiiMbDvyTNYX714SYRxKyx5d
3d+FemMcBlvDb2c8/ADvhiizKcEDIr47ayiduGCcvVgYOadfzKhPscvy+wM8YOOT8pPOU2ojKJTc
fJsCVZ6cV1QdnQizSugI9d+Nr2hsBjK2RinYcNIBxfG7jLt3Tj/KpWUkwbk90A7wGUjZXP0TYAHV
8n5w3Krm1obizEcNCza3pyUQ9ntB9A8TPXEFszkga+0gO/xFoZetB4uF/ue7IdiV+1WaUdwaI+P+
+R5Zd1OIM4eE1IYXnwuEXxfRuWQMcjsIxduYH5RLoDb+YBW+TN3OwWgmMrKAJXVHGt5kZoOVVg0p
oPAo4WkwJYKEkDlonFjG+CjqJLfZEvN/b026/l0AkNE2bk4Wd33vWVKnF8yPgsfotoYuq4Z2yqjk
tCemi4o7rabGEK8jkMIaoWInaBdJDUcCmD4UqW6GKwwFXSfkoK70dB4+m9buxtXzOLIOy0ROWz1X
55KkuYimpzaCfDp9tmL9DXSziDD5k9zzAJikrz9ePFj4YrK9opiQiOsYcveBUihPvrkEjhuLh/SS
SqGcoyI9HD5HJlQYmjXcZcN2VJgAuRErb3VUOtSjclRNiI2tLVCBFG1LfKwdA64YnYPahF/3G1wO
gKvXk8TjB0yJOiidrW4ICUYLfQFNOnIr/ibOF+Q9KQkG1D3ffneNcVtKsudRvjs0+MbOx0qOY7ac
ExTSs4d59THBKq2K2aSWWQib7HN8IuCXi5S2P8Y2w6v+9GkqMCXkAKMp9lXYjSu2hGhQ+9x56eX1
R+4R0U3WEopluEfwf5WKbq6bJk6y4NFe/FCirdgMg1ZB6RV42K8Aq4ogNDGtEs7BaH0452VV2QGK
5aT3fY75XI4rZjCh8BnmwPzvsHafdTdHzphtbYJ8jpaIrz3sVuxAAWZlJ5Spd8MGRl3RSHUoXSDA
PnW6AAHBCKC2Mg5KSNKhYH82TEXQz/TOPHfx0xqnF97+RWKTsaMBCcVllKahZ0RptXai1JA/dm8f
gYEMrpQ4jkH/jsG0svwLNR1EakgyqfZfEE4bZFxxPRgQh9bt+gh/ZOcNLbpm962DDf+gjJaYjJjH
hh0/VrTtcsYsBl91qFsZJPoph5+F8R3kSX/onoB3sMEs/TwLJaaaA16KiZrBMsYzC+p9eb09p3em
mIkvAKI2385re9/g/G8Pwo8JUuB9hwJZxA+0AjjtgZkjDu0HycnOp5+diDwtYDQljcu4sF0YEVYl
Knme1rYeK8oNBgkNlVCH5llxjE8+TRAvojxOriWxQumG+nHs7lb7zOMYUolPdnA6++c69YdZnoVv
ZO4f4GxoV2oO/05mIBcukyu/AGgLKtyGOf5MRKgbqLF6z7ETeBFEHPJEYqAGJIV3jNyjRyvNvtzv
WGKA4gDBrLff0dBHp/4cHIoIC9vmPsdAxH+62ccaIHnjzHgGjzknd8lJ77vbMBhN3wJu/VAi+JbN
+sM7+kWYMLJKSrK2wy6u/ohYljAaKmYTOF81g1v4OM6RarqETeApVm+FvnfkrHa+0FTnsB0Nk+mx
PqdN2YJsihSOkW7qtbNLsl9JLrn6QlkHm0Gw6T5mojb4NCnrhxCbtZCr/K5Ish5xAR8H+M4ve2mM
UA8zekFKaIb1cRFShgnL/6zi04zsafRBtwgmidTgh8iogrrbLoiafyRCoZEkIS63zcy7Y4Xptgj9
2sufElnvXeFhTKgMm6xIh2GQFfhYFVJ14VAUN0Mnyyc91FYWKi0LMcoLq0U7mmoiJm494GIdjdvM
DbdtnF6rNe1MLcrqQyH9HIdAg+QHjL04DHeXl/3BFnf24efEb0Uyh/VGp7yxTDdg3zYhdvFE+CD5
BGqwePeVmOLZejsMpu6xUNb2ujKKhl9yB4NfVI/hRgNYvQ3W8k/08Aj149x9TX+DIs9jhopQkzT+
6kIadZFYNzNO+th/uxEebb0zaPdNSfDTXhHuUpz7kuqssK3+kVQMblSiAYOJxtJtz7GmacfUwezg
fX5ycCMF6L6ex67YkmYG2VeEvw3e0aiLqKANLbsgP8QkzU690b8hGrLmrk7bUn1DAHdLW9q+Ledc
2QVpyQJMqE6+UKWlDGlRmlPQKA20Z001d8+3ZBtVojIkxZ+5/V27qCUcNNm+i5LgRPoe8LAZoPuR
2KyJommWQ+m/h6YknC2G3hXTO78Whhe5pqnk1M60x/k0g6cKAVwm8YPrIwOQAJIcNnF/IirRs1b7
6SlEvn+nxnLTa/vXZ8AaFNpFg+rRL3pzpcWEVfgTVn2/2V+ykidJWnCVm+cuS4iwSiHekd1c0Q65
ErI5zONAmhiNzKrNUHYVzAzDJtEinJ9UjV3qZcsIL334UWYCZIinHM2kUZ0MBlyxcLmCNW+wclq+
XRjYKfAJJ/rpCo8Zxw2D85pbpTP9fNpW3LiKbC+ULeB1ADyo587ZU8tp/GpsOvWBzZiztUv/BCKJ
t2pjZ/ZtlugHpaxaRx6m9HR+0Z2b57ZGofomgX7Vs89o6ePDbgtbN7cZGqT4uNXhdULW3+Chhwcs
PBnaPuuThVnVgNGP6SPESY28eeV8OorjBb82uevrcxHGAQxRNsS6PESvTRG/BRZtAJFxee2x1UY8
TrDoMLMNdt6dxl7NBmcLNl+0mkRacp7CjPc9tnK6JtMIWG8L0LQxYeJYOmtiiRdeTmtT/tHC75DJ
V4Rh0pQX9iewCbvR6XGEL34h4iKSOSxtncR98oMsMXP1DCnCmv/59OGB0URK6qBStBvdbLyiiCsX
msmF+1N67wu6yDljkVgJJt5k8pBnBGEJWFP2ESar5e2xXoDlGgZEYdjDZ3lCWs0xUWfujtl6cntw
cHb8Fq2fr3TJh8xVt9syv6KLcDEjmWaOfrpTm740m+hVn/4w4yvtpJ0mrlhCD7AKJ6Jeu3UwoVfc
GeyEGRCa7lFjAIUeHyCQnV50naAmeFySGoyItadKPcGL8JHSt2R6sLzFHgeUn38xXby0fZ08Rji+
Jg7bImDWfn0mNfdLyWs+qlksIxkjmnf5aznKvdtmkrBl49OOS003RAyoXzsxOzdQivfYtHcHFzw+
Zn554+eSMb0VbSDcgNK8lE0+fRzZfAnOsVA6luuvCA463qZkWMoCDcM9daslSSULYcUJ2UK5Nart
W+x6ZSdkIyGq10tmMWHgigyu+pw/b+0hrU2lBi6uWRc+dlDJYrlia0OYVAgDln1Zllj9oKWjWhJL
isF0T4/YqbVA3rI5i4Vt8po+XHneS/azA/wIla4kOrj+UwpyHMMFWgdw55rEJ/KVIk+/KawfN45X
yqhCMRUxuytR1claAcRzAxOJp/YOUQwCzXfRwXIIaT9x4Jv1tHQsPS/wYL5Ctpj9UX6sqznRpUzR
BEU2E2zm6Hcf49dWCf4D+HreVU390/h+WXR+Ac1ZagWjJiX0Tlw2951zTocZ12MPuplkiNnA2y+o
OhT1qYEQrei4TiUaC7rI4mLq6dmraIJAvdzODlnRVKdKAIlXJ/qEWCIs/Y8ZrMJGteqnfw6lP6kP
OSWFa7Nje54QwdHYBhlxrXvdu/ixOZGtiVSIJ5m/kCaMYkyl4Bbb/AsK4sv/TCq/w0YQbT6aFHr/
BHsQS0rrRbLQtgc9J/5AmTFwjYU61mjGex1A2ifZ+vHc2Q430GYWvt1CiRT0fsTgqD0RfDQmwyIb
n2GeRR0iS+tC/5UuNk9S5PHViU2LwCRyQTmukd6LUA74BoYkp9yH7ouiwVl1H0rBXw/+am28oIm2
hOjJNGyMwaoTuh2yldQyZaGyjJsZTHnent7DRDpziwnaBHbrywoqIT8/Dv5pFsqBRkBXEbGVvZjx
eJjgNPtrKDLDd5DxGyD4D52YzKGt2ALOEDxeISpnGEuir6lyxC0x5GOdcdk1+2RMOnuN3P+zAFiv
p1N36A8+yFohO69+RMQp/FDyLlSk5nwqcWLK26mmJ9R68qYeDxHr7WtOkxaYO24UsQDj0ZQedslL
64sJ5GATOpklMoWVTqOLtepBHQpOz5H+V/Nknn0hOhCsM73OQRC8ueq60NmJhIW+s2BEHUmhv9my
4zlH7WIqrUdFuFME87aBX5agcNimLDDCR6EWe+Vs3MK7GuWUakPFZWv2b8AXrEDGc9LCYr4hfBmC
qc7kZE1DOgYtLkwcQ+Z0VrP2l6UOyL/fVauZjfQdMjWjHP/k6UIgDVO9+mNMIeo5wC221U0+iSDm
SqOwEf0qDtmBgIytcXMF9+hS9I/93fdA+2h0JjnKJX1zIZVA7O+IMni9edvzaSuMEvIzVdvXOx6G
1OhQNCI3eLlHWxAtRH774dg83CDnRS2IPxEZW10iSAvBft+XePmpozmRjS7u3lOQ1PMkypFDX84v
HIf0Mi7cxtmqaQzkYs99GMACQaaTdFN93Or4ER/lAWNj6KYjGSlhz1jQ+piNDOFPrJyb67cUFt4u
Eco6LUkVTR0oe3F4MP3th39JwEGtmLCEhp641MPTH5ZpEGiuuJEl1NeXy1lrj6X6fh0hDHN7zc6K
SdkO+dWvstrJFrHOws+t1P30eL8DxKmVYP0lfo56nUkRLi6yadYCFdnPrJYT1s5jb1EXtgA25WZy
UqOVLOtAhQPfRVdv751DGhSTgQcS4Pc2HTeIGWHkZI+eZlLGWoDuCVcYXGKioR9yUILS9dYG38ok
F7UE2ojaALFNmhVD5PU0UU0QWL2VzvzM2lyGvjzzYY7wy/3qaI24xmm4h+Dva+DA6+gptygLG7YK
lKErb2zjUyEgPhEVBWe4YlfMjjd/efG8wflvZCj15yyOPxlvAONF/04Sk/Dzs8080X/w8NMEVg8j
usq2oEnbm+kvTO3dUJNQ8tTQNVlEYb5vm6+qin0J3rK50mATk6d0ncytpptSSWtsWw4eCO9meoAb
LP/Kifp4g2xiQ+/GuLyE5DjrxbOThEe5dX/R0JIStI551QgqKDgUn6X2RG/O1q7o5GAzUR17Q0G4
RE3tgqMGZEv3rEUKA5EfT1eXO2cgJ30OkKgsqcJoN5yBIvMgDiLWeKE3UzpB3zmtRF7CNYQyuvxP
cJrUDH88YSyCwJ7U+/81cNCrVXbXcCc3fmENBZXJsIPCqL6p1sxCGJsBqhttdiGDeQhy01pijS3W
8anDdP6nWs9pgWP/vvY72XSgWRJ9n8ZB78Yla31LcMko3Gi4iKRey8vRhttcaXsIrFhQ++T96BJR
JOlf11H61HjYYOVrZCrqn2ukmrI+Ql71aMifdXQo21T1lRgc5l398FkDs35E9lCWfzQ6SWP7Vw9h
18MB03wOhwdqMVl0Pd2S9M4O/1LFwDErHMsm261+jj4rH26l8FpgkalE+FI3xu8Pf/NDcwVKu0qb
tQY+f6kJjym/qwxoo/p7FsLxWENH4QV/wYT6ZUjcK/TS2O9v8VMaiga7tJbYe4Ler9OaYziVKhDJ
p785AV/56ZZ4mqiNFmsU+ud2blJ7CmeP7EfHYktMbAo31dFvXC+p4B1lsPHJdYUiHkPQkGD9EsyK
H8J0qsoPIrHKUubqQ4pSRJiEmp5NSWea2lUdfPgeAqapwTk9eYltQLU/aXTn/jE24JZkmLSlzN2q
XIIMiYGjeYhiI1K0e69/EI4ivdxFmBOkdmYKgng069D1+8Evz1ahD5sAmOOwYL0gjXd3t9Yc1LpH
qC8ATEwRdLO5WAwtpg/XXxs9ZzVJQZQelISroK9V81OAoTnTukvymBN2dLFGHVF544Jje11+s6O+
RCIuivv8gZOrvTaSI/TKYN0kiimrrjHTeEFDQV/w8ZUSLsLAfy3ekkHDmrYEy1GxpbeczOiWNU7q
/LLuzFDCndQbTXNLQ9x+AJBXyJB8MbIStmtcJhFhHAytyXvdp2OnwD/yypQbYMfn8WSF8pyF4Rr2
lZBJfm3PfV7OzD9NhbwLUaztxgGAQMSO6ZYz9cZSQY0m+N8tTyAlnxjqKlXJs3Q8DadM0bm1rJkx
etNw75mPXVMqedNZ7BXiiifjkmhGjNm0IkL0Fwi68h+2mE2HLashdgp6L/SRsfV33r+j9AVBeOyP
7Owk7WXiOcAHWgcHImPxu0GoWAHW6Z7YYPl4shBa8D8lwjAd006ikSigtdy/hDOg1JYKYvcHOjjz
BwWC9AXrTlLuVBpBuRW/lL9t1MXhfG5BBVvX7ZrERJ+8lWBw+5RhQ36B/k1Z7oK5VV56KhBO9xoK
6PevGh7EBOIjVW0EbLe9kttHpmg5ufmyoMuS5iwYUiGaDQnzoVJB0BqWeMNuwf9sg6t1fr2DezAN
7XbOM55ggbTV8Zkl0VqsmcJBREF5ipD6fdgxcYpBDYduxd01JkPC8XGZ1msl0X5ywY1LZvmwfYFY
+7iVwMpVVeHMkk7YLBRQzeYasEFMLtl38QoTJPkjsclGBYuMfb67YR7Oe1Sp4mlC0DM9d0Z9fbdE
Ujpy/T5yaAAm3PXcW222vGW+0lvnHoBREuxXILniFKp+dlMS84JSOxEEXe/iClCq/Pi4YYC2FBKa
FiqajkQy471CrfSW3kd7toaXWfIa9n4EkzsoTjNhy0a9PEL524AqGhn3xcmLtGiVvmgynRzosgZR
C7Te87rJNoKLVEVak+Q+QS8NSOTTOkd1lXqNj98B1SbQ1NTkpNJnR6XUPtXl9Yu84xPkLMd+Eacp
J/DmjimJaCEGox3lQYDNgxLq6rGz8JW6cuq+f+m8MTdEvvLwqu5hYiu6GkfXMKeq1biFxEcYbQqz
0ALh79DR/KH/SIVtjxoCXXXEgVN7HaCYH8/K+4YVodk2sIgr2UPaX9NZhvyStKfG2ljDBADMY8/p
EbY7Lw4wafX3EbpHiVxIK5SVnjR5J3AkatWgO84YMSTerrOTtfmmTs9/eWk3wRWTppi09eoeCXzt
4tnLM8GLpOqv3soTkFNw+3srldIEBYp6KxdSQAFeUjrk4fs90FW1yhTZTvrcbWIg8KadtwjLnlwv
JSPCPezHrTQlz1lNVMWfP+hOfy9kc7T4iZYcb7JYrqPvTRVgDWgd8SDLMpLYiQvh67b/i7SWpfDo
8p4DR+vgnnTqrzKjwK1TogUPnWIpa6BPuk53kV8vH6y2w9fpqOfCwtp91hdqEU+l2s1mF5eXnli3
VkMpqEbELyJumyHfrtPUIBxMAMDsxRX9mI0so/0qqhngunFuGDIDGK66Dq7wd9mFVgnfbaW2piNe
Z7EdAyWmbXcQsR+5kMjFY3hMubA0QCj8d2AOKEmgsMQdyFj+exx/cSD/MaYU72A0HU8NLuPNscLb
uLzI6yaU+XD5UY1dR9QhOnLqcmb9wIpQwPI3xYBkFOn3uM23zzDJxeoZWfwPnjGH0eENMR2u5A4+
5oBjecvhHijUshvzaGFQKarOfOhxLAwxQd5+jRxzw5esOXtmCZqe4jSARtroK+XbhF9Qg/wnZ2rp
qEUcKmdFaNdXt36SVOfRltlKq7/iMvTluDFqCTZPLj08ASEvFBLx6iU4QORuu3ZnZgPP3H/ah+zE
ptLXjTbiR7ee6RwxYah3E+9X7hKe+qTgTmyg1MkUrmjNyU0js0NU5ohZktroc3uae/QIhfVlAzZy
FIVma65NSu9gAFO6hBfU0gIpOLMPnLDZrzLG3YrPmIo6+WLXQuSVGJaFv7BCM4zRZT5RpUE1uBqJ
xFFW/9Bsd/IoqfHajTXoJVjtkaoJD4vjSg/GWWVJTJui/4/dHB7L/c0fgWJkd7gr5m49HeDPzesl
jPplsmolCWUzIQhR/FqujGpRZBr8y/enAVGoipJi9nQ6X3lnZSNvNPS+nxMhaD7NRlzucQJ1/uvi
vlJyXr8wijgfbuzWvtq4fCdOzLrMSDxBINB+eX6Q+pQeeJ+1DLdpX2vAPopXnLvzAvYACHCce9XB
IqL8cIMkyBasOhkIOiqgxxZogBfQhJphUbfzASt9HKEVOhA16SdBm+NiEhVDqNuYCC7Imj4RQeaE
V4LpHsx57PpdxeVIbLpvYQMz+/7P8ODp2hCNxe4VUU7GYYTUfhS56lorJYTHkL8oTREQ8NnxWLbD
63ZpWUi9mrNG/snEZTLE9oUEsh/Uia/5r/JTgqyLk6co/1+SkHvHIiuPw+UWuXunfAIYSIxLyCHm
7n2O991NveFlvy4CDiKJBy9z5eMFzuzA3s1IwM5kCUt/a6h9oSkNx0enwcaerAMjl2fHmS79hb8i
9qsRrjU0WsW7c3HU7BlxW+pARHu3gwKysukb7ylidWyPL9Vfvjti9jZZ5sxCeVJ8xk20s1KMrJVK
0jW2E0XxagAQEYYN9mmHBRUa3q5XzSiK8+PX33aB6j1/8ZosT3nq7+O2iaSrLEG7nRt9gojbMNqQ
UPePD2m178IKwFdmrK2T8CQK+k+A+5NihZwVjbEPwGi0OeRet3cPKM0eRI4Xw46y0G/we65+Hu8T
Scm1RyVhI+zPuCy+GVcZdHQYi7+uDnW27Xab42Cbd2alISWFPKH8MW+gTt+DUWC8rrVGDaxmStXL
AVUzFMfvPhD2eq8luB9hsv0/LYUamrwscfc7PZ/RUuIGdGPEDRtz1tlRFC4FHHyLB8DYSxNTqPCb
h8plTKElOUp4pn73Vb8dCeyDoA0qaXNXAlYKrRJycznHgcNnLDF5LNW6iG9OCgL1Tfu70qANpYtG
hSMwrV5l6jBQJ6O/RWEng02tkbRtZoNHkO1DOxpZWTW+HmIFCgX+QnVy/P88hWMdXEcyduINRt4O
T3Ojnc0Ksx22S9bqS105vURRmlnnPwKKq9RnpiOYmiIaZhErR5TksOyTtSLnmtT41dpQaUdeeJ73
zMrWyII5zSakSsBorbdgEMwbQ72WsrJQmqxJ9qw+5qoelAQX+tj1ux1672Mj7Ruz53XgFemlHuT7
651eC3i4NNSWp9UrwGt1JNG0rH7DQaCEg9YpW/+yn2zian4L8r/DrIKctnlQ1WOZjJO8U2i/wL/j
Y9j2n8jLYe/33c8hBrNSlOLUqITJLkR9yK7sUPU+RA4wze4XTpQPJweCfv2wDDe4NcUoRS/DCLH8
vxLWPKgAQC+FO+7qjRci4KIUI6AhMV1WWYr2sOY3MUYiQc+WPWCl4DcymUUcbGbZT2fLDmTY600o
oGKpFlYqz2JVpTqzqriIiOKDJqriGG2qOZgsVKgrfIn54Pz7x2nIQMCS/EucLkjrrPY1fPCV2Nwq
PUeJv4f9e/SCLfoavLGvk/NZkqvkLBqxSVQJdjJtwWymcptRp3eynEti4PP8C2uHhdx4x+qGxJMt
oAANU/kXS7YygVXXFWKYTTVrvRSvSBH7NdOtQFnuzGrfnfequ/SfH/fBzmku5QlCXpD5dMJ+SK5u
vgAzpFIR34Gd0wFomnha023eaGLaUDD3Swhy24mZltzrC3azgEumk0lx90LRKLw3kd+6W/0AF13J
PCnHmYQjs5Jek7ZdX2EbZao3eWKx4P4tV75NNFuCW6r5FUyHlgnuhLhjE4yRjOJX8UXiIRaZO9GE
+a6kMl1JwOkzS3mRIYqhGoC7u87q+ee87hr4p8JBQ59I/8O8WgCE3eCT9Yc7X8MnKiwExJ7rbrEb
MsFGfs8qA4bg3hfGHebXrFBOgCCAesQRRA8h3FzLTPMbWxJypChrKQz5m+Y8jNM6YW7ZlIv8zc/F
PksBbUZ7mDwK15Jm8PCq+oTaVE7wG3UrNfhSQRtXgPHlXYBxdK10ykcOCdaX6iNKp+z22ZtKk3+c
HnvBnfsOAus3dfyaxpuCkRVbsimeeT3thqFEiWQc78gqamL2amWD1QE8Rh2CUzYWTV1TLedhe+FG
/RCsu4Of9j0IbLk9/jd8bo5YdUsck+uFyo8HloJ7dxrVDzRsd90avjfakoHdhtlMZcPFsKm2t718
jGc2MfJqfc9y3xutRH2ZpX4Npn3GiujubR0ySvurLZ/DU/OQoQywjYNu8u7YXAty66H1STSwtxgu
qZMqdgoA4vCY9y4WUR1YyiPXbPVL35sxBjDtELHALLUG/ZCC5C+k9kkXbFcXLoJi/Ff5tpPZ3KkR
G2Rxd4fpYdPOOJH9NDElR3mU6GOgq3vd7+zrTMOhn1K4w0VkpqIZNQMfxSZWr+k99PiLOEVRM75U
wnfvYEqOZQ/6c/LsyhsGfr9UWrHsPewR0Ilb8qUemHpJI7xi3p4nj5yJxDySN47Wk9lHKs630EhM
rbtUsEn26tTw6R2fNyoH29AjvXlZ8LZHZqKoBwaicR7V5lV79bJL8qtYOsi8ATTPgRvc2zODoJpe
yMru1QXfBWphQ0oWzDDeN4sVIeLcl95aJMd5S5tRfKSuhHal6WO14MnYs0f8cBEqjpqRtJhmRWxn
QyaKBRitqhvlIsYEE9Sdi70qRHhhZfwoeexBPBrX2//hLCsfdfb09LeRT0kq8RcVUSGmvsaBHZic
U2fbdeePIlobIi5WYBIy2CK/YD1gPwwc/LTCCld859sUeIwNLD7reLiEjagakaqC2K/EZb9/USGs
pKYjBzTt0exQLD8cNpx1NyOirmtqtlQFLs1uEPK4JqxuwXrp45yv2AKeEU8iA8LqVgJaSCeXoGB2
d7ydawqaQwaw46rriX/1S95HAAVU0M4NXmJQn4XnwMop0AI4NWsyVhIRKVJZY5/qYgMyXCJZCong
K7+RooI5eOLk8kBlPUtrNgFBQGz8w04gK86wuVo9kEi6wtU3VqgIAsFiFfewxa2Wb3UOBW39A1lY
2rtDO144cl033mPNIVXR2UEXd5r89JJDgGtrPDgDKfs1BqwrAfl+LbJXsKSGIbjw3bOzVu5t+KtT
wfQosQd4ipstpelR51ZM19G7M9x1MowQz3k5GuXMquP9IjtVcjOJ6sh42I2uB94GC2QzbDrKMY5+
RG0rxikmUA6NyfUN8k9EdWmmdGo0IoclA1QE9KZ9HlwwDKhE6+38agfzGz/vsf4fiRyYMPW5y2Gl
kupsTRiGIlCsk05+YxQgpivQSUAfm+QslTSxt8+tc5/L9gUhHpwcqCV+ebOv9Ja+A738m7C79mvh
xE7QqdxQJhgK9g+vgKpLjxeb9Ju9O4FPgRdWLObonH9aNqnG+641lcX560V/tuDDangAWK9kUy7D
ucoknfdfXqP7RL8gUFgj+TXGmBGk63UK7a201KK1HPaxCupbg7g2OzkQuRsLErTw2TDSkuXKKt40
45QD3MGRgqspNepf/rwfZSVxtGG2gvIW5VE+RLhEISLlev32Rf+YOKBuVH9miC4LmnCSvBSU0BbT
ljDcKtI07JqTUbRzurEf57+/MZT+4Xm/M6Jx2ndxP1AROhsjQgSGphK1UMAxi7E7/YqMtcvv1Ze7
4wY8zWWe05NwpmX4aR2z6v72DsmqmjGkmvpKs+RcSc+wnNIm+4WegzU8x5jEMVDm3xff5wT6YvK1
UL9avQMqXLJyQ+klsojYdgi1VSls6H81s1+VngO7kooFSFKrRxSzDj+FwwY0HaWGQ+13Rj0NAM6b
2+jXkMfDjRNnWdELuA7M8R8noAX3wHqFtSqOBrW29MLu3AkPV73ab+M5See4l+H5+hjIbSi3WiUl
gvS9Ey5Q6YrIB7Jf6Mr/bFxHSknJ265Mx06OXKMJGtN+4VUsA/IgSkgCaMf08MyGYq+HI6LSDoGc
2q+S4Ah190an/OUyRJS6mpWAUK1FDJ/j2g6kBLNts2BHOBeZvyFN+YFVN9V0d+n7eL1E3j13hGLF
pQCrHA9FsNT98Kr2vtqfutZlvrguDxdZ9aql4IqI+kjD/ihju3DPVALepyrLS78GivDgOp38VMy9
HocpL0Hl8n/hSHb+hNdMRioYWxo8iegAlsF8esN9HG+WGWXiqeSHOjUsAtFkXTh72zItVeFB6L5k
X7U/aK0M4CqRRp6J1UM3uou5Q60fhDKbjkLAcrMUOQ3It70UJYaHP9SnPGhfpxp6SBH/hSMbfnDX
m/OFUdnhxnbvX4qjT8FBFCAQtnzaopOW0YTHE4tn8PUe82nYpxiqjEyiw5WzuPTAXyfOpth6maFk
Z8neVEzYSeSXCWwQzfF9My1eYHk5Gho/FORzop9TpLpJE6ro+XJT/2TBu9wi1VvQ08pjIowBHFOo
+5PHtNghcZQmoLSYNQTiZ9uCOkkqfXRf4BLCe3/EMDqBWS/8Sk/HqCkqfqHrkRlhY7KdQQQhiwbh
/oiIeNhSqL5V9dXheBJAiiA3W+yabbBIh0Jx6z+g3maajewMAV/Q0MYYc1/qUlpbFBaowajQJfp7
qUWAPvxDEAZhYjcoQcEYj0fOHiSAp8DoFzdxMfZo1lH8dy8FeDnJL6Btd9X8Vl/iVTPkj2SHrU2n
zQheuFMu/0LN348n4mEf04mKQR4LhW2SQoXijm8oZgSS9GoajM+82lSPvRQo9csd2UKHH1WtagcK
/0YauX0/1W0zYE5VfF8+djo+sV0ppii/miTbl0gnl4WtNNDO7w4mGSIcEPzDCLJ2vYFu/17O/9Xi
ntrk0mVkrjVhuSjKyaamBYJZKqgTv6K1TWpz6Y/9+IaabxB6uBz/eYjrL0WBDxhvjEMoFCRBPkID
/t5pDuO4/peJHguKC9bOR8LG5blneSHxc4mKPaB6njT4XptQZyDm0dPHKoEgoak6FHJk0XP1OCwZ
EwX9XGU3G7NwB8Fs69BQ4PRt5nwR0M9l9L2mdIsXU6ZrOW4V05RJbLrGPThu2hHXdhXnzXXyHQIi
A4QMrAUtnYbcD/9NQmacFW+nw8AwwQPXGpLgqBe3cAuG4avdDUxvcon+cZb70ZFvbCZxlHyOX/fe
cbZOfnfntlKhMW6GaWmdZvgT0gAy17a3k5DjWdMNcVUBHkWX3xAURVGpPIEgyqcgD2SkKeLODlqt
29cUTyoej5BJvt1+ofM2nf6i78vzMpN95znBVaDWiJtiQzJ2Vkj7ecyo4wpRtTk4t19kLvugdpjF
HU2bMNkMaMQFHRy4OWEhjQlYhBQKgZr4oVY/BJ9ZWMO+zybU+F1N4pP2pAvo5EmeJKca2ZctZQmA
OgWuISIXGxtnaj4dXpm6Xd/EdU9yatQnCtU1JGsi5ZMo6EfyzdXvso0zTFQ9p7uKIro919oRApwi
Z7ibabLSbrGrM+gufRsxdr2WijM9e/msdZzKNYLjSs80TYtFN6P8SuSpMWOz+yWm2SRE/f31lJRU
HDEgh8/HlLf6VxAQkd5tigdGaKOOyWC297oSnwh5GKVbMPma45kyruq3INR8wXEKR8DQHKo1cmEn
w4ljQctNOs72J9LBjM/bdK6c8HRFOF8ayxYe8OTNcFzPp9O2HIOOhCeRSSAo91aJbEqnKsMax6AQ
sU8ntI4P52ltPxVnFcJSGft7yPqe01LG11ejMXLcesMEkBBRQ++E5T6ef/QHEks+gt4LVrkKxPgd
DO+YxRvIGeg7eKbsXOCbxb4yNwpv+MGfosxx8hhVeHslKxOfFHuWF9hGc9nHl8RO9pbNlp1M4Pry
VPY5LiRTvXgAQ15YCikcI3DJVS77BrYnn2XLNSLDQdlII+eJdL7iPfHH06P1wgu1k55nenUsya+1
C9UhL1kqyks51UMMybYVcOwC6HUmNwBvc8hf/9UeeRL0s3vGU0sofpf9KuZPJXcO07PNbog4i0ZX
uAFZ3f9rQO6OPPQoIyojFAfI50RGQc1HmrWMRC4i9SUiEO1Gq5FS0izWlEb36oUYKRbL/dLWCi8E
9XesvWoCtGxnEspeG6a0CVAgiV7oGyJq12iNEwpW60O0pW5Ii5OkLZQ3lFEE1wjIKb6c8N01BoFv
tKdTBezaFxsLcmR37coYnWhfyTVH6x1IokprZ8UU5UxysQsMqeiPqypHZ/VcudmaTxtVzYO+cDoF
P5oIsKRdONk1xI7psii/09y9HboiDuWvj8ADd59T3FBrzEnFgQ/uOG4dCyZAhaZ8o6vAIYl8WBur
3FnRi+J0WFCzzL3oGrHBWtoB4e33CnGLKLii0/wtv+LWUJbwlAn2uqdVNlnVVljW4i6oWJLTj1Eo
M7UY14zP6MuwrXlenmLDHPxZB504zRKNU9VF4dvzSlMnsgcDM4AeqIb9141hofANWzBrUJUwfe/X
RD8qfuHR2VDuI4PkcHieLn0ltFRWvNKZjuVcdqayYVb9ZOKVHNR50sAd4HDJxuzsC9ZTgZlagWOq
yXrvj32BbpminzC5LPg5Lhhg/ktHGxGkf4kRwBDjOld6fBKlo/brKsHG5Zg46kioI3Frfrj5Qo89
BlOpAK1SQQsEMNhf+fn8f66PkHNwbnEJSOUxBfy2yLKnvj7qnQy3GVbzc/R1Q+lMTg9+ZvivgXfl
WtRk5e6MSVoDsm1KUbcF+qIS+xe61aXCV3Xk/CJf12o8/8oSJv3ovCWVUZI8AdaOQu6yzmYtWq3J
aVoIxajI8Hu1ufM+95XN6NR8hpB6xxhHxD55dmIzXp/lGlTysjSrjJd2kccm4+F7xrphdgQCBCva
GxJg0YwHje2Gkqbyo7wzuLkWX09SXJnFT7WxaXfOrkajdeucKmlSCyCGBERgrPo/i8r2lxqF/P5L
60z/Z3OOoe7j0W+5TpsqmmdSybnhQURNDgRkwaALgosuuVbcl1a4oUT25yQH1nWUVnMhseGbZrFG
yoS+QpL0mmxPpRdnGw3VR/ySA7YI9WtdovFXeBh8cEqn1hMRZcZnruRSTB4TnOh7H7G8unL1foL9
u+oxBeSTArM6z+6ZeaApz1ilF1o6MyVzOyYI/vlP0FV5XGLNM2yEeGXUbl+rF4XUm6WLjTtD+s9P
dCyrF+R0s4AeO/jJETX8KHAYKo4XNY9+3R/eao8lbWbrDtiWabGjSuavKFOK+yHLNP9X5/1b5EMg
UUgHFzcPHsVXF8LfmLxumlMZN1LXCDhUdLMFbfyW6tj9mOb5PTJnC8C0DZe5amRthsyue+3AjW55
u/NrYJlobUYp63xzaJNRcy2PI13fGvEbPl1LTBOPqHZxBmw73LfeaPueNkMo9mvnVqelO4GGtpsp
5aduAlN92GBgqL5w2eUUR0C1u7v72tfQpmc1xFoSs/XYwPu/f/sEHSWMuV5COXAgZuc4i66SNsj/
5qEasDZrzNZat6fKhTyeThdVqxOb5xo8tOI+bF58g7o8X/ueM66+t9Vyqi9GAkPR1eJscZkCKjxZ
BdwY7nBtOh+P5+rh5fyyPjD7aWRqOU+Beb7IRzC8evTMS64Yyc7adHOQhauLCjH8FNBYi+opVlxH
j6R/wX0XpsVnBoYrtcvqJpeChAVtkNLt+Q1JJ3+GZybeKgm3rXorg3XD9hOyx66nw/XzTChQ5bf5
KN5on143Y3hD2LcKZeRmvTxZ4bF/m4/cqBhL95wmw7ztOrKoLDpMNSfVMyrxU6IPeSyUy9w5qVWB
HWC7QYmeCwIsYkwEuEJxEvBgrQagDvcfFRoStadymM0kvkOSFGTZM3htAkDoAY3xu4GjJnhGIjqf
Vy9j04R2yckNsQCt07JZxDtTBTo8lcct+6OV4605eMvrgEUhZpXF9pZ0+z0+ZDOnUK9ltEmtqlxw
BzC9J+n6r/9SMW6c0xieDzQhxXb4LEX6GvERsgI+niIpUsfZeqqBGdYndQuUa3R8DIedQQtWjIhH
/z2ye2wT66MnqWVqbKq1vaQWypu0ASJ0hS3Q4CuazqIA7TBvqNSWyIFl4LTepCeQH/amgg1Xjqna
vSjnN79OFqQJicFGh91KdkxWQHZRSTlY4PqOrwXXpEywADWrlzTM/khn09QP8YT4WapBu9oKMt2Z
k+PJ+Ftix29TOwUVTxQtCH5cKP5ZkOrf88R3Bdpwgd5aBIxJpNZRT8etaysqDbqS1b08EJmFcmPD
dmt1bWLb53RI899UMYJA9tr2ecKtpFyeQtkPzTffUTTDqi9kc6aQIVHg7nEBELo7ngQWSA1s5au1
yZ63On38O7s7WyNIh90JHWtQJQAlcUkQ9KCcpcylB9dOCwaV+hQj+bA0P0eaYX6NMTFi+e7dboAm
HiWsE6SGba+dJ1UdiLxC7rC/lAZ7T51DG6z89Lor3XG5oIjAGyqJqGRce7BS1YjiRijY0pRwP/Fr
cx9QJ4vy+F7RZyb6FLhD92W+IlQVDY0qh8fFPLMtHpukxWmd1tURMoC3SK4iyW+G0wuK3D+rnMCm
Xa3YUlU2hGuHpVGXcAYWqaAGpr8cRTi3jkA/bPUdo/nBr7JSGhp+gww5MelHZljpqoNfWcTgwqb0
OVnsPOYBA0arjBgRau9cmI3oZF8oNd/3QSM18vIa+ZN4v3TUJCwSsQKCo6iQiY6vsaxoBS7FON5U
xvG+wntvyA+ISeM1C5jkNkzOj4sbtCxPdxuqlBCAJ69PDDK5DFHxUA7lkEDGPve02qfv9L8IgTJM
6JfO7yZl1HCAr6BmUqNcx94ZR2PzVK9AHMRx1010eR9IfKaau7rg/tlQFyBaiwj/Bt/djzkj9i86
HnJrze5kUOFmucDYQEWQfXUxVy2U6qpaR7GyQXusEB0OS5h6CDg297M3IimkzeXKsprgXnUzx1eP
4R7zl3E8bJrmjLtpZ3vLujkoVy4Qe61uqcK6cOt8YSkugl4C76GGS3No58IebmnbxdE9Wu7dvWCW
O/HGL5UPoln/Tmxo9ODEns+Z+wSzdYmXacqrXfAbeg+VtVit9d5F1SPdhZH76Ah1USdMqE1HxwVW
nHpslqkKbWMJZrVH9EezWSkxGeC0up6g6P4lamFH0C9YgqQkOfC3lc+PwMDVv2Bd8GR8K+fR3SsL
zhEZ2HfY67Twnt2skA2VJmllQujd7CRyf032duXfpuzfUGkw7KUS8i2SUr8OAVLAJFEJsjGnn6om
px+kzpJYMjYrQMSFVviwxl/Lla2GeNI4u+FipJjh2UlvczlNILundCYYIC3sbzh/sIiTAVpQOX7E
h9YxX3vABF29lktm2l4usiHaKxs/9a2C1ojYpbA5UVchAuWAz/64a6SqB7IFA33s0PVCxJdSJnDY
dCn2Ym94AY9GgcwifhSQRNf9MbGKCGgpgE70mFLmGmApkw3VFyI5SWrszqvBnAEtYNh4mXT9wjml
WPTU3rewUJGMUfwd50O9upQgpFaR7v7o+o4Ts3h/1ELQGnGcTjtz8ZOsHjvnKA2YcN+Efg+/qVYz
gItno8jcdYSZmuebIBdWRytvKndqr/G/qc2oA9C7IMWx54WLXjrqRXxw7LH3+Sq2fhLXTb+Xdicr
5hgItkmchM8tO/U1I5/5+VeA9sRw7OWUfn0x2ANk5uC4bx9OYXO1LItiQwlrfLK+BMecdW68d/4m
zMUslU83Yd3YlG7NeztDTcHfYB0SO2GizL9cXaXAO8XF5Y5QT3eH1xeLOpI+Y5UBDTE7MCLLPr2p
0q03PMc1f3RgG/b3xTOGAg+y4RXY4cR/fFiPa1xk+RH/isChSyBNN+2LNvnoLCzxvTCI+vXhjMcR
vZcO+NnRksKK9Bn+bwU9baXzLne/NrIJJVq4zbUW7LF2+eutXGRrnHQ6JRiWGt4c0Fj74aGNzTGw
3UdMTrTevdr5lgf+2NpF7RwDPuDNsibj3ZKYCEwgKAv5FGpaZ3723Y6J+PltuXcjVipecPFnzCCh
COPQmlplvIcJjHip4wqCeymgiaIqCCyZ0cy0PUPRDm3k1eVBYEh7+Bykiwc8sggjBVe/nWbBTSEc
KgX1qp9Q0ziM15L3+PHDFapccbfB0IoKf5njkIfrNL1N4kY/Y78hNFrziQyYrv/2l1YkSGqW8jYb
X90kRLKqoxkurQzWERdHTinwiCPRV4s+zQahcpA5DrmPUFbhGURMaUaFYARct18vXo/lit30bL+8
nrkXnF6mDI6zRjmhxBCoHY/DMyqOs//iWmI8h+ErP1xJKGMHJLDlJH5FLvS3ywVIDL2o4Ae24Wrv
yagcIVLS/AnJbu3UDB7xr7c9tdcEI+GYPb3nVxCNr+EYvw4iqaw04hwsuJII4rkH87y9pouFGome
+9k723Vf5+0WHGTJ07gdkKLS2UkjiYx9SsJlQtl4DPZ4cyOSfBmC4B3tr27Z/mGXN95/xUHJbXWd
YbzJD0joIosUxMLiQ5LxZ/JzKKrCurHbjVh5h/FD8vvFfZMmS/ulcwh2/sdz5L6MxkBc+tF6PONt
deyNtsmtJBRVfef5Rl33UZUv9B14u8jD31pc38YTgGetUkIBFkNV/mvZOMrV1NAmj7upwctYqgE0
FwNHlwOxmdE34C9K5HT6e2SmMp98VJAls9PKXcWHNC63aOEbCPAMUIF/Spm6kJLTFVFA5XgltvF/
HlzaGgDn/ZueqetMAXlLB/URL1+oSBqW+UTsy6gxv3uAwrqhETiRmiH86wzChqKy4GlOGKHoGjm8
EK4rgvUBn32/mACSvgG7nNnzBY82Z3svvd9arP53qpTDSaw8S7ysVABrfmmYu5Ds8ngZnX1SlDum
c+1cS+TeMVXVs0AktUOL8AQxOqVpAmN3tj9jTawmgw+y6IJEDWfKQCOaQ2P1qcMZkPOlTxGxoRPt
Iq7W3J+XsekKq+k/49ZgFYQYqyTiuX95lMew3NHvAgbo4K5tdvjgc8QWqZtpK4gOdzDVMTMITZNv
s27g332SDMNsqbOG4poAcP/JMN8xA0SeSMqQYKJ8JDyqlT6g4o5YzHe+/UKw3hFxYOmLMIJ46JlZ
2cFP5lOyxSpYJIAsaOm0a3b4bNm7JGf08TFCDOUE1zDtaNXhq4VLlfujS9d6uOsLDqZ141fujCXa
2jC8YJIXXyAdyJq2R6mE7DiQT+PYG6Pxe9nDhdtSLAgEOoK0RozfcpbU4g1W3oUI6wwzNlLpzXbH
cLs5Dq5AAi/8BBa597s0v2w15cKOqpUvOYXdHEnO/zwnip+9OGBT26IOeQ7kr7OFFN/Gf5Tm04p1
WRUaBfcb3IbAu/ZY06qfIbDUdTpdhKkzWILPKDeV2nPuWx0KMeTqqoh2cNcAnmQJlDaHf7WCXd6m
FOpHDxIhi1wx9e0ur2bU6mZrEptYSkmWLTKhQnT7KSwHxV8QGH7eLcKKsMlQekV2cgvjPBAiilF9
0nrm7CiDs775iBMnFurub/EkD0TLPUrK7DilTsGf5quE4ProthV6oUJxSgFSUhbRAQZe2eZF6TrC
cjJKIi7uyEFejHYEuWpvGsTweA6RRvRe6OEptQjwpTpKLKTItqj1XAKx3XaiSpg5D2uOcgQcQBpc
7wRBWiTRqhcpBmlBvnFiJskGreu7Ke7SnYJ6tSSvRgOIf81lmvDr7JZfgc70afiii43/89LBeM6D
wZLDh/Cl84gbVTErY3/6dDnwAPAFc4YNY75hVVRo5qy2I1Ag1uF07AhYa0YxCv34LPo25yudzkBj
iOuYtczfpVqrE48mWJt8HqPtT+sQBin6iPJViBqzwY3nZKZOan+oeI2Gs59po2kuDOUdgDqco0Ri
qr2DlxKnM11Lts+Vgt1LlH45IHgLJgNHbgKXdKsQg0MgmggY/B7NNVn7+kyd2Rxjatg0DEIalTLP
5nY6ZDumgJ/DP70l9kSlT9Y3yjcrwIoHE60yqEwjF0VLsCrNO0rQJpmFDHUR4fV9HPnsYP4ZtPk/
i7GtEy9qW5O1/E7LPlkqqs2PNYpnErqDybeFt2onBXSafAx7ZET5+ioHf9Kt0oPFrV0wXEseZNwj
ItgBL/6sRJV30IMZeX4VTOFQE8LEpq8G2u01I2wojTSxtltIPm/lZ3sAYzv7Ppa84H4G2nRvI3/m
i4Pm19qPrYOKPDJj0ugJ/5hQF7tRxUbkBy6ZSiMsvvyz1vJq5a2sCe4YkpX9oXNOegegJEBRY2uS
SZjAAWPiVj674rGvJy/gN9zTdHaB8eNXyXsQFCQ24pXiA4djFhTCTh1dg04v3r2CdXg7Slc5mIYv
4m7plj2NgUG9NQtfwq4fhq8pLUPlxM4jD75shJObBi0gvZnGFCiyvy262LIlWcLrEfblHi0NnAGt
XbSm7kzLrQQpRQvuPT+EUuxRKdZSGBVu9DBQYdknnZZ+CeR3zJTwATS7p+rtZNP05JyLwnFNneCk
Dprh+SyI4VhxI72g2DXPrRDZP5YKjOBjz6ORvHAJ3+i+CHzkawpY+q1rAgbslvo1Hi4y5zWpblwh
BuhZyYaqV8KDj52ybfwCuyeBoS5laUlpMsxL6lwxEfz4i6CdU8zNU0WaHytkfyDSRgu20KpwWkUN
Hn0WM8Mui8m3MibKkX10za5b35MxViTO/1qfq8V/FqKPxdyZ0cjMpEGktt2bevPFc/GmvsLULHYG
aNKNHNJxXpecu3hUssDbT6iEwUw4YkKbKj9Uxo9J4uWnfVP8ZM/HB6+toNaDkVj87nTn1LRmJX4z
SNuIX6go9KU3jk5VAHfqJf2ARftnti1s5DddXAW1aOyhoNkNcxxUDcFU6zjctiJ4QojZRNBuEmCg
MR6RHiz2mOj79I7acQzYbfYeyyKuHroluI4hTkDgext05JF3zVP4+ZgPlnfy7BkZoUx994Z4T+zX
qt/N033tU7rHdm/lq8xlyk//LB/0rLC9YkfKH6wTMU63+7YV2MW8n6czLLPAUmfPsghiZM/vHX7K
U5pKvdNk4KgsF0DRpZkyRsdEknYNRdw5DhRUUVy8Pzo7x2b+u+ZSym7NOJ1Kw98hb75VJjKDXwUk
h/KQAsZbcqAGuRff+w19oD0oOjxjva02iD3hsJnwHVqU9g2sJ7v9LwN7dMtMYWj1AT7i1udZ10QY
k+KL5WFa5ml2fifwFwfADUCOLdqw2LxjWGa0sMYkrj15Ve4imJ8nWViaG+52jFQsRwReAYwuRGdS
SVRFvZ50Xsf3RBg9tOBZGMFTatjs4gOqYueUWb1FPkW2t0V+H4lidtI2YAc9Zuvo4zqY3/zxNfEL
NJStOzR5HJhc4ffmtx/hza407STsUeKqSYxTwKarCq5Vz5VUtBf3xc2/AO8xCSJzDfUO0i8W5IvD
4JgTp1E+szBcKqKnJkDnUfv79p1V7ldSg1vZlfKX76DYR0Q38ZNFNp2S9GNJr9vqd73M10RstiYH
CphvLPjT/PdOngGqamctsUoJJ1fVxX+NYIw7RM/sqVvG78tpIQ88+Lk1oTcNLt1QdoC0A+524q0e
2/bgjhm+5dbrsZvcgu+EJBqqfFTmqV2/HvldS5P2POSqu6yCDNEK+zh5w+k4+VzsOvi3s7v0UjId
rVFY3XeclMCeVPLCct2sp6JSJCoC3U6OWsDDkac3hSN7z0yX1z9TRg5ipqoHVB+J7nMkyAPngUsc
m61QA+d4qUQ/sgiSXY2lQeSqlFXmRHqDUSJfDPwdCzCuVc+P0BeXhOek7QUioCgcW9+xiJPyQUNP
BhnzbRLwTlVKdbZXbBx83zMsSM24UtHB2pmUJge3XghVXtQvspwP8RcIe1pE9Kp+G8accZXFeOt/
njD+d7vzIZXRw1e6r9FaFF6h4hPC4trP3QQQiaXrtpvdouOKqy70KXvuPGZzo5wnsE8BkJsLg62F
A1gETyb1SNK5AFeWuoLpya/hPgkMnBCjROS5PBNLh8MB9Bxl7ya+lNOu0EgbS4hzMqYB2n+X+7K4
y+bnW1yUSSe8kxWKAg9R6iZduKRWu8xlkbXxgRh1Ih63/+on/HzMNefk6PbJAWkfrnREf2rRS/f6
pzNEnYheJ8HKxI513/evZj+ETIp8vl+Pdam4CzUSKDwSUvipbuiazyNOlAPkQYg0QsaB4B6O5XqB
sKAEiCqHUTLvohA++8FgaAoMDouZNrDw9OJnnP9UbrQgiyeP1247IniXM1YiuQ4pJH87lZQlZ6Pj
1C3ezYq4aJQYRSa/1Gh2xV6LbM5zPeFxB+jTnDC/ksTz4UOaOrZbDl9nq7nWBWOOsTNaqBGKB16N
U0EKJlosWBDoiirZGXQp3ZIX5oA8EzolJikNNuK5LnolpYQWz+vwlLa1XqZqauolkEWuJ0G40SU+
JJxDxfRYkZ+ve608QY4TrRnAArUrQQ7BdBtlwngYzPOoTmpMbBDJrcd3lpAo6ujLprW1M3lDwim4
xYdg5+Huth7VLv38y3LWZ3DjPewUWk3dgB9s+iHUvLjaKQZkgXYr+1htb9OSFFuluzxioLhStGmT
j3kos9b0O+tBNnPLt4wA+dqylqQRHG2HzZaPBuR6qMHvmmo5pA/KjiNSC6LX6SrMauVHBSueV60Y
Uv0YbroCcbwD9LeMRgWr1IVHQtLSGswtsHTz+eL7wwu8J+OgAaO8uuBqcb7qPjeu/mwGWCuGdvdF
Ia9DWAq2Y8Rfm8hrXBT3dPdYMDI2zBAtMwUZNdGuy6CgQRuhAd6hYZ++U9zRKU4c+a5jnxPWXaOI
uEAqL7kSrqIYPEQ4tve/PQgu85Tardbn3hUw1ztCwzU1d/3sAZHfmKgsqiLt6vrFKKfKXWmBlPuf
3uGh+U3aQWz/VeGrUzB+zXbE9954nBg503ZS29WwhFVY2PSNcvH7E0XX8ryw6E3eYG8mjwCNE4qv
tlFlMyvaQwKtj3LdpxOuyKOo0NsT1ym0E830siDMfPDdrteJzZL2s/h+Bgo1KNJYL5/T+dXYfKMA
VMc0FttiKSc/kN5rIOz8JU1yC+J1XFNz/a+TRfGtrWofWIbrJoSGSCCQaQ3Etfm1xlrx3+Si8Gly
PUR/KxDqFwSqC1A1latgEZ+SQeVWtRvpZU9ncrFdsdoGtfYACCRXeMrRHRdk2bmK+akKx6+u68oO
TdGtPhUvQyUDtMDRijxTFLN/Xr3ypgK++e68Kbu4+9DmlILSckaYJmR3wvEZ3orvBW16YEMC1lQp
GcFAzAhm2ByJkdz1HvCU6eBWVKPxESdcfDEoqwddvuXSviPSKBv+DQFvXcgsvq2206XzAGxIwbxp
WFVjgq5ftHhDZtHywFHx8FlB1oRrTSGsTQMRS626Mh3deDwGkPIXug6Jg0K/tjWB+RVZqlLPBXLG
kAsZmyrEXbAw5lZ4y62c50DiLxNNT1Xsts6o+gL2Tkn4XgWlvaupLYn0XA+f9ED6rZw+5VxrZQWP
4TXJPPliwcYmyHLj8svTT8WgkrRcf9XQwwaE/Lfn467z02rv4q2ea/Rj/wBlI+Cwj02AC9d6X+OO
EdRSjN5b6qA9vyFkV47R6LZ5nc6Egzb/txoASKfHxCX2wi2MHRBreR8PUKAPRqaJf2U1ILbZL4Tp
xN3NdRq0AU55v4u4s3eyGt836wH5kcfP1dgZsZfHz158kpihEmcefyMuMAavOWB/936mOdO2aALp
Ff/z93CeY6gddeikXxFaTscAx/Y2lwumczztKwxtFwpA3dUVtxsdi3qdqV2U01po0foXXgoNALh3
fw43G4TW1FUi5bOpHRkS7k/TP8NYR8kle4r3Z/Ad2/Msp7ZxsTJrS+MMsxa35nwJBGQt0YQF2O+/
noIdDrmGgn2L0F7MYlEzXh2LsvZOsnj4+aAx2d+wNp4SgKhTc7Ouipr/QRZoKIuvKisOoo+FBly2
cmLmHHlaRWbhuBmHKMXUrU1BpdPw259ia29YxAzynM3wP+b4JfgF112NGSzj7zGbiD5o/NKtoqzt
FaK/g9LZmNY+o4FbQ6UfWN6Y1pmkef8RJsdYngQ1t43JhVY416GpRz6NWTFexnmHhII239OD6oig
5XKFTNhQsIl0AG2WLMsV1L84o8qIntH8ayT0wPu9XwKlZiZk88fk3gTq6AfXQQsRXqbpI/8/VSKG
wt9SLoq49D1h9ZgvLPhXRye1HIhTfIfUSFPa2h2dgv4JjeW4elUnW9ovCmR9w5DZnae8EhoOAWyH
MsMmRXJYVZ5iF3lImGAjtN/nD+Ll8z3Pa48PyVy/Gxkfi2LDMpx9gxjOItD40gwnE6OjBudpDrLM
5/Rar+uhhYS2TXX9vqLbZTJDMycLDBCO/YR1CvoC4WjsNF5pO/AOuJ6zctK7nSnCDZ0mEEIbwci4
GtNdcrkftQzj8+m4MpGgTDEVbuJaFAJLsIeHbBMbhJvHO+bNK3Gcil12DFS/Dc+oEOMGNyADf/FY
//r1N/IMpOlHFxgDvQ5NGoJzj1zjZWBdhZTfANGS4KC4iqJttmtjBKxU0d7AsHr+49QydMREDZU1
K2MzuSDQMI9Q2puSPhJoAQRLWxs6VNvQYtStmuN7ySqHSNa5irSyDwYVftJuR5NPeJYcFmsuTxG7
sP3Bt2ziTiKach4fItAm62Zk2j9Jji5NI6ZYu1MerQXiy6ZcUfb7BV93q+kpPZ/fKAQolVlAk6yU
NHOBSA+9Eq35fEi/IoaXWVJF7RN8BMIqdjX/DBnQUE/NsCX2HxcBLL9MbefDgYyEfm83u9zGxvmf
Wa4G9PfcumZ97AMFRsAG/Wi+3zVOBoen3bB/ry479Vt1BUZcBp/KAoiO7J5Z+TI5vOi0u2qTn+P9
iaSJlG8XNoX+LdVTaa01P2orvOmmHklFwY6L5jeY8b9wPGs2014PY/X8wkyvm9GKl85wodQYnVu8
xngQ4J1rXcY8BP1iani7zcrA8ac+VQxsugJoRR60XPgPfOtYWNPiyCfpdnla9nUDohSD9cl4GCFQ
S2MOQuMo2YiHkYAwYA1RnrdbaJNuvFAt77RhaW/9jcG957lHqNX5AGkxvJfwH4EawmMiNdcyFP2W
ppeJbGphojTRmscVl7FPSC5Jo5hYZyDANENobRvMrNtpadLcDL3KnFZ5cln1MtgWMQXDnKL9vQFK
lmnVJYHlG2y7hwRpKFIkYSqfhTN3Zjp3d6Q9JRLnmIxOD7AKGQvgP1ijLhfV9FZqewVvi40CYdSR
I+u+m7crbhgbXjVyQhK+eeQuc2pFisSf+3B4pH3PceNikVJPB0u9mYwB34tJPLneHQRcnI1UjYzn
vMWPEFruxsC3HQkHEHAK9YTPDG8Bs/ZPHEshVMXzA1y+zMxbd1Rws3eJ9ILRdRgwLnPgG9Nb7XIw
7I/4rEdF7BQNWuNrW4VdcRXoo+trMgMT03XnjbDjLUpOs9uuk0cqwoEPujfwbZD4fdNVdU/gtH4e
qgnha9LcyJYUDTK9wopAHhZd7Oy6DJ5sFEx4zTN0ZnoPLf7mqtoKiLwdy08mAvLXK9pN71xSW9wH
C77kPK7Ads2HKWh03UgoMhYB+AS0jGX4Aobu7WC27tJ/qG2b7eoWsJlhr3VIRnehI+tb4eIg2F8F
rAn3It9s2OJMTUwG1K0yATLAkNfBl9q3MPMAHWWIFqop6IIxGGL9dxcDDtpDU6LsGikwKUJwQCVj
a0MMQdQteXkQNscP24Zdj+o0WrbE5201uGzvdfzIDncvUG69gAB3KI+z1TQQZf9kLEsjfCgtPAwV
JJiOK8vusisWoLfWK/gi7at9/6rLGpSxCi0iyEP8Dg5nVxsEMe1F00kqJ2rRM5etaAcoz2oNUSZi
jOfA943JhrCY1MsIXBHUIV23WBsLcotimhWMcuBqJEGHBxnicCgrtPSMsSMQ8z4RhevOr97I/Uzl
DxxVELfxhk6BysNOXOrGrqrh8r6lRbXi2U+BFwuS25Bo+fhNpmz5FQc3WxWgR/LlrmLPX43Yvrxp
nh7R2+Ng1X4WblPCmlDieZ3AoQGPa9WId8EkY4WzEbH+4pN65hGmcifc4BfUlqSpEFON3n7doaJe
KU7TdnuRYk+0SEUy6zelVmSI+Hwvtaql/hXEx8nEGVaRG4SJtlNa5IXW1b3l8/OKTzKNF1mFtaq8
0+xMV2pJ03HuJxaRVC82xBwJFiN1fFbje8SBAjorX139APWSpO0FjyXdySR1RHi+7LGFTt3h0OrK
qu5Xbh1c3gpNOTyTAs+pGGF4PlymKA4DRMtWP5Od6ZaEcvi5uCeThEzFyooTvS93epGstnd0LPTj
AJH/T4XyiOdhqCCn7IdXi9BTZ9dA3i70NnFkI9Vp10+8AJUw1ESjQ0mOEjeWcNZCiIaaFdvcwIS2
rpt6FuiIP64lU82agq6mPBEv0ekDfyV7afHbHPClbdS7QXCD+m9j5HtD9mNK7K1rrZkaFiqgAdvI
DaXBwEMCZ8ortxtfaxdVwuGu0Ocn7Qmz7kFhsZ/iiMhExfh3w8pTrqlk5HxUPbRHpfd9Eo7Itlff
B2jj8+sRRvAy42aClhh9IRT+4MSpXGYK0bHoAHBuMxcRQvT4i9xBLV2pvfQzP3cngScr6QC3DpM/
ldE227SEn7rXWapCup2lgnL9wyEhY4orKM1Sqs4YqKpor9Te2TM99W1IrwxnM4VelnF9kZ+f1TFG
EG0JLRuV9k7p0o5CZZFKmEpaNEgQGs9Rci9zSHxkJWawDa2ArDZgXTg2Mzj3h5+ldxwHGPY/WrgO
8jYGDSyZd3R2H7NjPPD6mnIkXaMeuCYVGHfHeira/GWpZvG432yWzSYOE7v2Vm3namTztZOZ4esL
Nf8Vum1PUsUyyV4DLtXa32bgmX5b+5CWluiUydZ8RxokerTANPDabnCfMx8WhMlkv8EurTubZkX9
VVml+vC2YqPcqunURn1ZlOarvp+X3/MBs4bq6/ffIb8PsWjCPHJuj8uCKuPDLXCt42TfbXSpUQlX
hgnxZygmjikWskKN8PY0d33fnm4AgWZ9p8QimYYB+ZBPlM5Sv4HtozoArIBpg9UopnL/DJsBGxG0
Ro7NnvNZhm+CwUotzbWh9RbxTW37fzgWe1nYEZChA3o5jOVk92ryGjiDQdDEMXXyAPcqUX28S4tt
A3vuWvI1CGvW8Z1xbF2Io3yPakgJzE8HdcQ1DYMKPRPsa+GMkM0xQuwdgX18hD+/OrwCMHhI8QLh
pO7563uvKAhUHUpnmTIyNOLAunM5R1LF6cuYP63ucfCFO1iYG+ELbN3/GYbTgP7qCdCx2Heo1Yp/
W5dhkwHRvRn4/IlmSabwpxNRszWcpNte3mIOjLBxAN4KWUHUSaG5isAUjLTudsI1719vYjPLJUtW
dE4asNTArFZM2pS/eZIZD/qOgPe53J7hPv3E/5DJC5+XtFmjrxHTBev0GpZXUuGIbHibTWWjJuio
2UPZvyauC3Hhr15KGToTSr60OKkGkVZsfKWa22qvGKWbwMfWW7ltkl4KxJR42nAOLrz6mtHn/uHa
OLztUDO5LTU4eU2KjWxs4OtXgeIIcuwIRBzuBNP2t5gn31BrL6rT+3+XxUjKQ5t+kpEMKMlKwWat
7sqoDsTc65QAKH0YDzuHGIChxLPXMtVLEzfi8WJlH5SX1efHHtlTT991viSbkwS2BIwP9CPGA6R2
xCcShnO3ECodoO89h/lGWHm2GyPJvfK08T/R1PDK6yHZuX+aY/D5rqEVSTAs9/I+l2deOnKid3eA
d57B2EdHtJLtZ+N6mlw6Asz8CazigE7ExWzrPFmDOrYDC89j2dY0dVZqXgUOuXPXoDjn5EHf5yto
6wdmOJH4fIYS1aBGk5YD6fEYgo+OnXQIWkZF2ZCA+XCNzXy9c7b9A7MVxLe6gRIzt2pO+hJNGS/6
o8gqev9Cs/7WRkMCnpZG7tQtVOl4vz+PnQUHRb+HU/BOudcMnA75P02JfEo1PqLsvp3ATXGEvAXr
mbtqlcJR/FnAb7uNF+Zeb9iEBhjk3unp23jmeJ/LYJcaiwBrhO54BObgjuJEqG+x5DZ6MhgHFtCK
BwW8jG7m7i2LOx5MyVnA6A77XzpE7gnZFQVEpFnII4R5JjuWUSk2ukGJj0sAmeeXspIGNjK1JXbX
b48MICd/BMZshF1cCIIkD11gr33SZoE2biHiJmYCii2cKLpbgQNej3NkuBXfxdX0BowBOjhiXXdT
qjZvFrF/ofbHHrvKAOE03oSWViBCnYcbsDuFjKtzv7yjl1+Xo7V7P4/5jV5e1gumSCd+dpYUbtad
ix6QWsiMJ4w3SiWLy8zYtg1wbbdvzvja3JJ3OawVpDv+7gllwQrKEz21c4i9F3v5UGeRSvFTwHQQ
b3lIw1XBPfpNz1Bsl2UWyrdhA0s6nH4/gH1Yx7DGbpiyKgqLw254t3DKF6X5CPlrlnDGqPayCpvD
VXT5h9lbNBTET3E+Er2EdyvD+yT5S5yUhOXryQ5E5QCAMdtdo479gNAkjIwMMCwSWX8EA20Zh3zo
IYavoyAN+oKgQqbtU1C8Ae/QU+bM+LRK4leNMyXJNyARF+o8QuTLW05LfOI/LUOaK5p3RJsbeP30
3kSHXbwRc2oGXRhPF/Qvo5/848Eo8ZIKUhFmApaAY4UsQtSkc1ITH1Bg+YTAsGCy6sBSuSPK5/nY
vqnMDFFSchh8XbJZMlsBRsS6ExMPNGFrJAZbMGE+Q0XW9XapC3lBx8mJtRDDnfaDsTB82rslLZ3D
Bl0M2cwp/eEm8H74YIFGGlbBhOTfSlynnpzgYuWnsiP+lHuWZNyxN0dNeOxaTml+jQkmqeQiOCTA
j9PixevORdNqpB6zIwVZTR95LyNrlTdpnwmj+0kGulzVBXii2EacFAG89+mszF8RPLB/YljqtpcR
ik2s4DQva4y9z4Wl0PvD3+l5Q3VTwQyAF6oXJKpIZbQQesP9Au0C0hX5RJWYQ8HlJJI9o60HzIQj
mQz2ZcJU0OSo90mdNTCkYEZrfox+d7I3Ias+M54jfn5N4w+0OgUUNmuDwecHlJD7UoDbM5b8QZFV
hVjvwjEeTK/YoCXXKwPYS38oaCQeK3JMIOicEXzHWadITrVWpUj+TAjdP+mmSlCaIT1dNXg/263B
1ud3PNpoqVf91oSBJA2MmSxfsEGcstBSIzgoR+6dmUjwRuihTYBGDUBX9kLBYn0yzX8ClNQmYC85
cDGdqj68HiTa5dSx75ILmwFE4DGJnc4oSuHEUjBqKqwxT8mw6Kc2eNMacbA5PSbHxbdtWs3r5O+R
JxUZ9jtw/TDwa8aQRMcl0HCP3c1JNgCK1TlMHasL7fZ1hlxoLxltV260/txWp0Mvd3dErd5YEVZf
kGi3ivh2JEiALdWCmbOdtJW0AIXhTPsDKJgmEuYsum5+vLwHZtlg4SRpFgwXcBjsa+cveVdGVL3+
k8AdqS/V8fEHcZ2H5o7pvEjBFDFV7MaMuPL0dpi5FBQIn3sTZTP0tJgkCHGpdOrzBW25WmhZ3s+L
o2QZ4qqIjcj+hQXEVOfGgg4gFuY/HKN5hN28zZRwVqJFXGaYE+mXI1Zbp+2DwBLyLtM1u3oI3v8M
LvzUzJTTD2Uai2kATmMbzJLMdhUy72D0Ep3/Xywj2SklIT3TsPVS4LFNr10PrbVVKGPmK4fZW4X0
ueHxBv0qGCZ46Ophplq00cJE+91CXuCtC1QyBR2AAIwKLdVJPTy7VJ2GPNwq2sQflfwWz6ZTJw9J
pTZgvp3A5CRlGKoVIXEdI5xRgox4aK/lAo1bdvGXYbM7PbPhghTrKhlipuBVa8LuutU8dRRl72rz
YhUPWkwSJP/3BkhuXPMr7B/nOIcOEpsPOz+xuP9tlSyjLckeqhq2thZxn4IUdcPLmylUpfxTLBdf
J4S5pkGHRZ17ZfBG57/Aq7WQeXMQ+C4ZK2+2ii3LRrrZGOL5bhu10mm7Faqh0cbCbz/WE3uyqUnf
e20BIQFKIU0CYtgQJ8Iw375RIqGaoHE0AGoasz290g1oazIVZUoUwqZd+s7gp5qYAepbrulZykd1
9x9Mx/jAhUmGJyVFre/FOYbDHzCmuDBZIRmYrD3j83154+eKeQ1uUlxbhSkubIOxH8tu/hqZ3x9F
1r85G06juRLwL8Bb9wRSCqxAhUVj+4GjuhKBPh/61ROapLu3Cn+QWtPwKaqiyOZUJ/wHm7xP8LLw
IyZiKDxt1YPe5hIFiEm//cG5zY5hYCdBpAwbon8QQTEgL8xtp4YgdNnhoRkHuJ0rMxMkh6xd2i1I
/5++s2adbYzbLXGh92jVBQlPCSEyKnpDE1Chn8nY6EUGtvkNsH+nzik5XYCk/XgbbaXJjBecsJFF
tGcpbBvtr7fCA3tPSP0/QofP+1J+ajoRPNwuOQmLV0A7PO9jvD0dpOlG7jDwK9L737gXI96yaq9K
4uXmysPBM/ulTGB71cNvaPami13w777x7zvCAlBbFNAuKL5IPDfvAmaqJQUSO3x703z0216MV+Su
+mnAlJ3SY56DSWRlsya/xr8ya4E2GZ4M5Ez3QZIkXEtOCJdksAtEsmEJaD1lGFNsYVM8tpjNhqok
AUXGG7pbVsLB6x8SYoARsHWOLP4Du3ZL7xFZUnJS08HG1fxlHXOWgmLp/9hOElySvOYwkqJdAZbZ
qaQJb70bnDMtlMIHcJpd8lzU2Xl8taBZa5MuCFN/zKmRKlQxxKHLBmuJ+4pyRJhzm5XzJUORUjTi
OUfIVfbflBLyaLbSEGsRKbSa+aG3u0W2Yve+/21iiMLDckHgefMAdyJ+BUyD/WOMb8I3nsYnvmZJ
pu2ontgZTlhgaDL260mU9HFQ1DwRxXU3pq5TcUzNJevgPwZ73WipSJNd5WnfiygLQMgmqkY9K3nZ
Onngm885cSvsqodPFAyI8Nbd2cooPsSYX8GQK0w+9CDUdIz70eAKigdTIhgry05EHYozWwPXn7zA
bVEzZfzfAYl/VDM1x3O8PmyyJEnjojP2qhyi96NxIcY+WzFnx4Vy47DuDD+wVi1HzLv7anJukuqM
QO2D8Zmto2wyIQ+3VJY7CbbiZcXTc6UvBBWVPubx3YpZff9k94rpyRfU42GKJAH6Rc2pBV7CeQcX
ugvELuhb5ftCPv+v9/8JDEYuhw6rIk5HKz5AZoKO2Xfe9Qy4iOJt3FURfA5cc33kdq8LE7GE6Kru
BlWjMc7mjcvHxB1MsCrj+RClWDdm2irAZmZv1ZCkKVDqJND86ANWF/H2j8bPh5phi2FvN6rhl9pH
7St3cxbRbVfCLhtUYnN8HHPoHd98tqHqNhTtNROd7nv9bsSeXmBhywCuxppwslf8F1eVYAfeyQmG
Kxe5o3f1HNKTLXv14c3sbQ1hwXAoqyiiA39z0mLtDw4niZUgX65Izup4gTjjnxp24XpwIGdX6aUz
cBxTDmPm97YI2oOSDMA2//0HnUsBZ/anKUt+O6UdZQq2UK0RBmSRiB3A+A4hTDe1IkrcndQZ5XlB
T/7xvPsB8RWxIcOdPvKuPc8nvjlQsrsU0kGKO/FBpTmzQTFVTAAsu1v1h3JEQO/YG1BGITKCseVq
fRDy7WGrIyiLB3W0FWKF7rUxRNHGObGmmXltLhuYkEggfdwDFGs84WdtbuAOC7oZuhlq+utKBlUA
kShHxfj41grMsaIAz83cWNNGeKPRtI//hrvotuSe2POxzkIcXwJ4sS3/tHifLq+xfYSaERwG/gRG
Mbxu3FwB9lYNS5dHl8bP1PHq9+m9xKhGNYV0RN9a3XAursuBOAvu09UzlpW5QX4TGnUmRfjow1sL
PVmc2kZD3flyUVNSsZhTOBiGrQkgwYs/Rgs3F7AehTcJULaLXGmhsvc7bvbqcHHWldLiSXjc/0l3
WUykOAQqp9aRXvewVqCcT4jxWGoLaqUgJIPFcKzbBq1bgtKuQcVZ41E1ipp9pbfD67gJgoRrCXpx
JgeMQ9PM2f+dvkHpiJTmWebMbNfl0QHnWOgr8ddh6E4HKIB/a+4ccYBBZGtDwYTefV+BAjbl8Slb
VK10j7ZF5/OvOqLxE0p/JNZBQCjWV/srYBX6scE/KLzoygeS3zSGOSjm6Akt9hbkS+IAHUtrwBa7
awM5fsbr5YPhTG4jqdmtt0Kjo77E6k0H16LBJMAT53QIMksniExJjeFglkxhOG6X5hq0NDBahaZB
/+iMhyaKxL5QyNc1bPzWEs/VNRgCaCz/gEhwHyZi6cAGKkDHSWQCH2jHDUyKVGuD/Xp8DQxA0nU8
uPCaLKds2Tohs1PnYUF9FAo4Z3VlLafcW585IJnKb7YPNt84G9EY1maMc5WhKAHZ6zDginAjpish
/hraWpBdtoGeIeKFSyiolOqHpWqfpBlM39mzQ0He0QmB5gvgPFOvyx5nAxI0W8vJ2r/QpzvjHAdS
erGp8dSI9WiZa+y04W2BUwBiLSSangzLuazXLOrDi6pznxJaJ/cT7qx2vBBrE8p3Sq9Vxaho4c6x
Dj7+pvDuZwgIBVSNEmdz08IaQIFu50sU1B2xzGIjFWVq6JWMs9tuEVOgH3L1GwZygHaAbsTjXwdn
Hr6dq4WVAI2STIq0FRuK+NKxH+jpaviJ0leBTXOSmKCrBfeA6rbDf/Ka7GJd5GdejMZi81ZGSIGq
0wwur2gqE7eJ0biDf054lS8Pxa8OFImY2LjZN/hDio4GUSoWuS4F1Uvoh6tF9BLhGrNu8/8Y4hBL
J9Em1BSWTnVXacjT/U+vVen4tPqNM7gNc5Jg3dskv+cjLRlPrIJ1cz0I1ncAEVPCjwiaMhp5Cx/n
tZ5dDijbrvrAe6AN0pXbAdJ2Agu/lS764LE1ysFcxwsccW9du8Lv0BvNpKl8/qHS3phqHEQua5op
NKu8xMkqGUNzz/LMz+XGTpJFKHhdRq9UN/F0BnEqJYH5wDvYEJuxgTnIKPuINRDwn4kJcEpMTZvx
YRMl4sF7P/HToF861Q9l7UbdSnRv6IvZNk8Z3dyeqeB5QbCyM7eOZ9fmXGHTGcGAJQZEuDgLTEKd
ncuun6xyR5eIXwLDw9aU2YXucSmZtQ1kE/eYAW6aeAcioTHLISr3kcyZIeAWIehwdeqUVlazxuxb
CsDDOjcQvOPlvoJ18q+alWcRCWHfE0Cfw1eoNa3FEFYBZliOKOKiJ3z+1+7cjNdpOUEzjpBKTMlI
A9ij543MJoQ2Nd/1jFbkVGcsPLMwtWsk4tkQNajL506WS7FjLsuiErGkircKs1+lp1agOY8xqc2w
nxSj/I3RdRpgBlI5A/2z3ZCsSEfkbEDw6wOnnS0ukzT7u+AMpUB8wVXvawniYc0/Y+wGzIyPZWXJ
QzWdwFSS3cjbpC3xe+Pz7BNSiXJMrgnKKegtGAOr5bssgi8wNhITk8vZeKqgcozh6LAwMzz4y/VH
vXBqoH81WXbODUElsVqi7AF200TlYdcVEVzf3SNn6+JGUKXKCZQKuB7lvkBFOaXnVheGuY0LI/W7
N/r+VTba9ytA1uGlDqIehZZ+brqAjdleEvDP2jTiz4LHbQ8Ozdl+Mqz4s8KYiZSWMGtLOg3Gw6cP
uXtdnPCo9kLBeooNLyeaza++tOQ6d6f3a7XKWjLPgPdecoX/Tqyt5UD2oAD4bYjjp6f4R7oP03VU
1Fl1qznClYQ5R3fofliXkBtUq7cpqiXPo3KAxwqvb6XfdcJqWPCCUtx3M+3Zjk9JNh0+o9Co7pqO
7zV8ReyuurCqv5byT1o4+4LQKkQB+U1rFPj88HStigYMsp8XgfyCYzWEu32uWS/ZAk7C27art1FW
uw2Szv64PMUnLryYiJyDrZiNTYSYlUXar3eNh7/Bl6po/wZUnPzVBBAbOIV7oL2S5ALrbVqPCwX1
uZ60SjwSCJi7ZXvCJD8Z7rn0YIDLtWRPXGgGY0SoLY8Qm9+L8jhUEpJOVvznVyadADYycD7LnmeG
UwLx1YAQLrzlYRMOvTD4OFEv8Zz2cryRSPkJ0rbMYfHkDGFuz28fcF4lKzDEuJeUrxET3L3b/EIV
tg1+BBR935GbMY2YLUNtZfIqTvQ6Ya8TGmltrGv1fiFuU3YBtp4KXTY/GTeMKfJP1daDTds+JsyA
9fkwhcnlkzoTFYIOwr7FQdq0IYKy00Y3TeT/NXs5kUXy3ZlxMjmn/lE+yVMP9lVIddqckFe51b/s
VZ4TGDaq/nr4X4oJCC6X9kZMV8WDtOkf0o3GgemIw0Zhl/97pTghwcQtI2ZpCA4IVbiunLFNImd5
blkv69QMzdV4656eVdbHvToS+JOftHgE9TYP+JZVQfzAYNe3ehTbptAqrrRcqTULsPFvv/mab2qN
XPWzXK1OyufBkVc512/QBBCGhLD2wHBwZEvSi58rSPybke2us16iH5YKa1odl01UpqZoR/z3Q/r/
KojRzzHQXmTmznBB4Uyzu9bC1HKe4H0eTeTCSq36V30E5LOy2Zn7wcR4iigKl9aZdIXBfXnMQ+Rz
N7nhRrHu2kBjM+mRSnmXCRHJatFu1+/7lANTzq9aMrf4pDvQz3uJ1oUi3Q3A3iMIKoYLvOPcCcib
fkEcDj+IObO8jocfhOq3/WPpQBuSmrGr0zZSE2IR45YeguVFdic+DL1gRxWxpxrI7XsXvM/GUh1k
vYu0+VYEzk4IUZHkbzMoLpnHpPZLbFhIM/o8eZbEjF/rstbb8GaoHKF8rui1/yrR1vhtMx0q+4vu
6UuUsX/wY9hWkpRl87z3tMKI2mCM7gN+BOnuO2J0EV7OmFevr4lWxJNbNV2t/6Tz47Zpjbn+79XF
P/yKNvXh3hndm9T6oZIy77jUHRI3oB3sVQoAYJnFkvCMAtu4YsMGLsrnYlWoyQbLqxhP1GY5J7ni
plvFiL9iw2T4x/6bB9IZ/lF/e10/VJL0P3NOlsBp834Rtb8Yj5bNBfgl+eMez9flXeH5ofWTGbe6
40I8lvONScT3hhNfq6kq4Ptv/+Cm3eMVg6GYPy2ew1Ma90/dT6hXcBDMI2p1AFH/UB3zBmJkTeKl
E5FNfAO/u2maXtkZIQ7V+pkm6hAYNKr5fcpGv6tWax2Rs8JK/m7mC1IvlChSiavzGAo7A13zRqfG
6Kuf48gUiy+kuAiB0EZ6XwpYm97QnYCtUYRD4L/Kk74avkcd2pyNbby1znYYYRaNemikA5wt5q65
gdZnfpXU/QH2+chOTGiA/nYEh4Y18pGMtW3Z1T0ufETtX6uEWhSB9RfI8xIyO11rwmMeEvrU8B7K
209MCBh/VXl5gXKgkI5+nMktTy+s6sNw/68j+fHqfXC3QdkIZ0KkmJi6dDU6eICBfdbGti0NzMLp
fq31TdCATMdZHS9V2VgwmSHuPE08lCL9JN+p28RJj/jnD3ZKRGWzZZztm6Aw51hfy0rrY2db1X5W
B6S58uWl/KsGa7tdWUku+EliGrOGul/LT7gieBK3XFt4cXNyvXUqvN+rk6vMyHJwyZCmQ8taBAsN
NxUhsZO56/HVAu6h4aNa5M/TP1bKWBFqJYOcekJaRCMfIcJQuMMPBtupRHKNfz+d5fo94jGlIMzB
nmSMif8R/bFZjYJvA8V7ZYjqJaEB54c1KP0HYl098ELiPNKg7Jm3t/GdxMdYCR1rZBOyqbPtyoo/
jURx8hTS+UTve4vfUGQLyaXL5K/jwHow+HCcyVEtuM++bsvQPwiXVMz4VyE4D/1JicIJFsfOhtKX
pOeOsOybMo7q9lnzGiwN1KrpksnCbTjpkRYRptbLt276Hw4RwYHoStW9K+N++EtdZKimkPXVJH4W
pCZNyiNGBxhD/oRMqwlwgAAy3auBxVxuj5u69GKT/6EswQ2HXtWAK0hDV6X1Q1efRSNM6ws78ILS
itXsWHO/9sOHMM39v1QKk9MgMEzJhnvpkBWxbPihNpGsMbua2RtcbwtrUq4/hIpuCZzlJ9i9Ug7v
vCwdfkwJmhH66D30m8xzyGdyCszEqseiAq/M7dBiRpT6XTla02z+NUaCtgGpkZNRJUABomCS5T9+
Fl5DV3r0BqUTLKbekn6KCZ9w9v8IxnLCe1qbR3CtQmGrSSXBQC3eGt5GB9b4fnMypbh3b83NNKCz
erJhKCfVKejkLOZ9iZuGLqbW+g7Mktrre2lDB3VXBDHI2y9eefaS7BULsMKYk74LUMtmdO5kHaNo
tGIQeVImKdYzQ3soz+FfII5lVqb01inbWXPL5Fc5LIL4fPOAuT5s2dfitvIeAdDFtShIo1jxkTxv
SY0CPO6pVBoxBKnovxrk3C1XMOlKv1bn7kSfD3EoS+Bk+u9bePv7cY5u/GB42/tSpAmmVmQ3sH/t
ZMVONscMLhOOCrr/FX+LYfeLBMRu2GekARhH+VH++CXP0WbvEGmeBIxT0jdIzcyhtqEI3Fy9m7MW
ptyAwgk1evQdNkZW39U9DhwyAoX/eUeE0dbnxDakRGORO5uJD8Ri8W2m7FxpjmRiMheBOWbgtkgk
AMOyCRbFjv9KjRJH/A+XlVt6CLm2UBOtZfobcoLGrJvlYoJDG9ACPm/77jHquFXEpwa+0ddmkflC
tKsBAz6pt/+H1RZ0VkElKahww5RPLTkVGvsf+jhiHM+UXT9R42kvHMkprGBnvMM4mGNL2OvThPk4
B+jTULqJ4bFFUWhiccWjL0fbvOVrNFlX0r5isbRmkxHQyZVu7sPxJ1ZQKrr1K8mf8AMLMk0Sg7ZH
j0gLFfVM1+03iJ7VRazo39YGrB1YlfFhdB0tceF3JMunll1z+/n1ModUo3az1Zc9EuUNtNIB3qdg
sn7aVut9OsGpYwO65rpLoRPM4FsnM4Mia/dLHmNRzecW4FzGKGC8RLmr1CI6KBN/MsTk93HKVR88
WIImzMciGF160JZf0/ErlINCdG+aK8XltAS0aW+L+B1SWeBLMk28vfXLs6pcPuAsrhUI8K+kdJgv
OhyjrM5p4sro7BYxyCaZm0mpN9wKMa1lyRvLezBMgT80MAUkpDy0HcPJ0O3upaOkpUL3yU2fRkSy
tq68rCXuOYhhxmVIrAQ9VefSUbttM7k+biryEVKK3uOtLgjp64gNgAAC7rXhEjbtoRI+c4BoRziO
JgsW9REQT2RPIrC5Bz7GLl+Z6PVQQvAYFD93uIITu4jMVi+V829sHqRzzTOVVB6OYBaTXOOCxB41
8Ej/n/C96sj9ui0RB4FOf2VzsZWfKord6IdPK7Ydq7RLCOcZSaImoyX39PNb6JRKE8rO94QGgSNE
3EnyKJY/fWRSJMTPmeO/gHPZd4Fz3IhUA/GpTPFXytX1dCwbtZoT9Ufgj8HSgu6Gwo5YSiznDCk5
tjlbWiQtFqrxaM0ZDRbMWM02+N3XIUs/eydRadqhnOAYsYLJAG1CyXhDpbjgRaMUOBEaxuovx+hT
w12wCuYNO0lVaxpM+x5muMVZ/18VMnlZfb0X95Ft4TUPopKud/fZKyfbjaLHNpuaDVcbjg2hb8Fm
BgaidPiWLrfQu8B/9m69moNTFUbG4easVxqEIoZ3H96hpUQCr6TB/JiytvQTO5KUEBg39NgBmrpo
K0ZIpYK4eNUaL3q8MfusxbdK+N1Xwm/LuvPBETSweeWfVwQgaTRLFXUFENsnhAXbUInvRrD0HiuM
84TCoPwnY/wVFPumXynmFaI0sVSXw2X/xkgLMFx1Gu2UkNVnmL9DuBoteibK1Js6f8H4azIirmWc
voEzqqrWYZQ4xsbtiNMJsnVaQA63YKWmfdtaeoVzVAc9vN1QTnWdaQuOQHyUxnCfULJnF5o75s0k
KLDbwClaoCXqyLCf1Q4DvMYyB4q9EBx/6bITx5999LTZ7QcuE9vz112kqtU6h9vT53KjvMmZoMEc
AHzWqq2dl5DlTdue+DqkAmyJoKXiDnSOvsTV/Nims1Sk+Piyb60g/UMGJM+lsgG02TJRuga+o4hX
2Aekt+Zrp7ueYMBBhxkgaZ5lEYcx8+UUz02JWQ2kb6wCQsDNIhsd/siq3bsXGqexn4njS0MnnSeN
QLQS5fRG14GL9ePXuse/YKcxx/woubHjVS179J2WOXRkhJlsSo1DXv5o/JfuIO2/EUFd4bcGc/ot
9kq5jd5eGeGHAQ70NcPR96gKNTBVkQF25OQe2tM0l3ljXkrb4UDprZATWHKezDv6J1FTRHjJLP4b
1RwIoTJ5lt4tLqvBUP7ET0URS2WejzPv/nnDZ13m7eMxRLawvWOEU63am8QZ07P6W6cQrgWtAG98
Xt2/tWniUVxCSCzIvUahQidr9J6O1buB+LGU0/7qCPr0zDzd7wfmfsXvIWVWUiq2c2IdOlVs7FfS
/cF0SNCA4m7sXasJTasJ1eexJJ6sRJICoYmts0LKjls0s5/155D2uTKTNVpGOIsg6YfsAEja2NUt
V4qf3Z0PiltAqoTfq28pH85Ta/FfFze/6zKi6+ZOxAfoh0bx16+JX6nQHKxe+ccXTw7OakLsbPlF
xvMiOszGF3/Wmjv8eD3TAXIYyjNGajZn3v2lbDWjtnABDb/GWFs8QN3UQrqLBU6+uoIVi96V0HJD
FmTn5Zz3E/ncw78rnsWlHm94uxqM924s9tdeSMbhoWalvwoSSJRouCwdOu8+BXeg/fxH4dejGvdy
CadTx9ULYvHiahu22ns1dq7nZpAEGa58lLgIfGIZ72o2MHWYqyuGRUqWSiozwC0lCXmqx/NlW59X
d3Q2ajFQKdyOLguJ29zPKERdN2+4/H4KDvKkMCch9PdxpjuplRIH0hOvfyjQ7JbzfSx8ZmJW+GXg
PXtdQ90NTX9VP9+ZUBIbeTP2OiuzQZFkQqUoCGsYgLbPSwb+SCxIsUobPQ6N86P4WjgYeb5xmMY8
yKymMiaD0wJcLoSwOnQJGHi2FMNeGUSFaNaPBn9aq5zQTX44un2obZdCZ5yUP0R4+qobYeZeEnbM
rg+w4d8TonCtQj09Tpur/mK8i4/7fDpBEjSduDhOQjV4RbPm3T+3fc0eFmW2z/niOxBZt0RZ7+Xq
R5nFurH67njM4ChAP7OIq9Fc2o/TPGmfu1CT0+2B9qVU1ABhg7dQEiE3JJBUZV2r+Zy43Xt/Lc5P
dJeVvt5vUZRb6F+YX+U1zLxItjX+snUVwToAwwo/eraVpSYjuWkK5sPLJYdo5bj7cySt3RiPeRCb
7ZBwt10CdjC6Pa4BLKgp1hNyB4cOECHkPi5ywVP7eAu2NQ17ie/BuVtltgz+gBNJcXBLuWnEkt/A
H8gMoB5wXCEK1LLvYOWfBkk5/SEX6bq21VbdcZhWq2OnUVMWZ/OYn5HjzNOcgEakXO3bveYFlcFs
03B1jhwLiYUGt6/sAIin7hFv72ioClP+peh0JjHNeMCs2vru3sgaOx2qR26H0HqOva85yZhfp+JN
rJKqqFKHdnLkCPo9dkKO/u9Zjp501sM7Kl4QGIeqHYOkktX0XrhM7ruke+lLiEUzTjjAu4/Ab2S4
Fj5CQHVYtrWQZXXDDZ15oZBGcXeLdp807tRtW79VRlgDobPz9AgnBej+hDRBvHdgRn1a49sRchds
L8oXUEgusEyOTjKShXhmyd2uqzdaGEBFoglOG/o4G0ItV7ExtqSf9SWU9qK/U1vnxjqNZFft6Cbj
QVFxfWhsUr8Wv834VTRKDygFAoZl0Dzg+xFZKFv8Qq/9LgzRob7yyxPw8FOljkxTVlqmINW68U5x
oRAITUXgh3hsm8Nzh7kOKCkoqDebPRJm+Gr0jjaJyhHzt4wXlxDK7A2R2e36xtkL1qLap1IWBXyU
yYLROGwL87C2Lkl1HX9Q2b7tlq0T9yz4kKGpvJpIk4XwPf6ZP//xzJsGUrA07I3uO58jfddy67vz
iUi+8iicKFBiykUAZqy0NpLAjd+U/DlKLYJ0KdSjKod9TdStIj50w9GF5EnChHCvBLOZRPn9IWc9
U6DwEIBwVyp6fUx21ccAqGgxJEXOyZy7aL2rFtNTjzWW/s413ah+7Y3iXM2yLHjjZzgjYLKsrXip
brPDEThLw8lAtZeDYcI7Fh2djPu5vUXRK/ZkZp80uCEunl47V+LVJS8qy5HfPeNHe8Pw7uJxk7wQ
esnRtuabmF3y2hJaAC67cv+Pq5VU34++8yUdJHXrWhV8S/Y7qFnWXMpix220yMJRuz448eIvmQeG
9thOIsu3JpkQz3JQ5cX1jvBCl7ubtbyHZ7GpUWbWw3cHoObwKK7uNB9k3DfFjKGTgW8JpMgq9ymY
CPalAuCWNYozV9yYmhYvR5HWyJhgRMeVfdlpQLLz93i8ELLVIjnhCRGgSbrpLCSEjqwWwG19xDyh
Dgetqaf3RNTqkr96RxG6Zg+jBfXJXxvSB3XECTEFERhhbu5QZbQOCR25YSlay6O97aVd1NR6DGRU
FSrV9+hs2kIn/m9gN8DWgRPaBccQvjTNWnOCpDWYucibqFAahO9HLrhEg3J9mvEgbKMYRdk4ocyB
lDemQ1TH2+AawiveTFChi49vQtOnkXMBYa8Jkkr9tpe+/2NQJK8AUAwxOH2nMTVq+2fT1kyus6bj
b04YS8SU0r2yD0feGWzJ/l6azDDKPZ2DAIa5zxkprPhAuvcSobEgpKODMSpBMa0KxT3Z/MLjXa6N
S6dhg4sfM39Y8rMazBXAIjsTqvns7Vc+LAhLIXDFcX2QpFErPAwvZAkOPdmAtqQ7sUjw8U1g9H61
B3sj4cA+kI+SlocbMwjoAffUnOB+CCfC9gX9J1aoqKzeIlghab99WWgc0WS49rUXHbn9FOVAwpHq
4cpieZGX7jCRpk9bR1VKrE8denHjw/lHCunAzIgAdauE+G2h2Jusnd+rXKxcp4zsKJ1yEbQ/vKkF
aAcyC+zFQ44c3xHIsrpfoYxKJZeXpSco2VTN4tC6O4gCg9VKe1HhulB+JiCt3smAwnCzSvIIptJT
x5rNX9h3rUrDuHXOYka47WDPFcLR2HOsgPqpeR56vVZGoC0GnrhCkmBlk1N0cZUlEXxYKq5rRvbQ
c11rI4BX6pa+HuIz7Rpb8gNl9BOEoFFacWW5BevdiQ1zGhBwG+ajf1vOhQDw+lhiHVw0X04wJQX5
EqlHTw8UIDrnZMPqSI8voWt9QT/5mZ13HigyrQUAO7YKK8Gbp+0zsijgP0ZCDFbxPHQoG2/4qbEw
WDKkDyoRXK/7n9tLeuocZWCtLWKsdxEGETeehxnTxbBAbgadZS1ksMjs7u30+gl/LGojtDodM/rN
hvx7jqoDtpVKQKqsJedprQgfRkIf3Ct+oTpHeJCQpVNlt+AybQhDQsvxlnk2ILevcr32hXG6gvh8
66bdhZ7YoXLWZbQiNfQSmYZXdmRleKp6gHHTqWCw4WFTeiWyVaZ6+5uxMTCJQukA6fMcxOmni9uV
Nscdk3HoGpX4o35q2xLpBDMxK5FhIiGSGXbdXRyC6Y8QOVDwsYIAchUrOT2DnY9xSBvr8FFshtZJ
/YHhOGd3NgfzFQk2r1BSHaqsCW5/rQ/3A284E2Fw9MZSiXK/4Ke2utAvW52XucwjLka39oDpbtSC
LyzMLIRBbz/JaiBb6AMLWPq9VUTHJtaLkeNcsL8DnFsPCxaqUH520HxktRCeB6cA5irjfoHDj8Nk
JhbQuJ9aQsfkjhPe9e63cu6TEIddQYIBnZVYc4Mr/PLRrbWnEeNO8bWQ0AYuIgaFajawGBiwX+PX
j82evna7NC98dzjoz3ss2eReSIwIEtO+ds+Wiskyh4BPZbWIqaQ72HOCd/2GF/O5CadmYjKNfxr4
ylvt+Z1XYSk7e6enSyT7vq/dZiX9lzcO2Xueq7MA0YipDFkhvuo0q2w6DFozRxAEgzkYt9byfK4Y
Ig5uNnwt2T93ab4CcS14ok3Y4wWJ+LxwsEuTB6Ejp0wGssqRIMSVyOxAMB7Vh/w0nFHgL0g4uc8R
NIiMexyXx+knRJlPgdmYQI4ObTpRyjAWFlblL4hMmMlJBbpgbTnJRTApbQ5Oe8CT8M753eUJjMRp
OZY1Lgj/z52D4WPpZimng6VBne/fl4SOt8pJU2o845xf+sLIeUfsHP4P39hgrHJpT2bvzkFfPmGE
9m2Kc2upGWoYXT7cAtR6JkqN0p7HU2jMLpIXhe1JICjqDX6YWF0En5kcpvW+Uef3PtzG2B83m1pB
+A0/FD8SFJ6wVKjNk7oPU2qEsxWZ9WE6Q8lJ07iccf7mop8RB+Ogmp1W6fYshQWWAHYFkzdwogKH
RyC3XIN8YHqrPj8xMOT4TXe2iW5j093l+7PNJR1TMykkv6DUlL3aXmdQkLB8Q0zNwe7i626Y2s3y
SMVG4a4qcyn3Y7frtATL1pz/1WJCEXzTjl9ITCeLOa7Tndpoh3cxjRdyQdO/vEG4/Inh7+eyTVjg
Bli9bftLz44i2AkQfZ1pJD9ANqoT7gGzPbac0HQGXdzwK37d+bU8dZ7NMlpxFGeSN+XXDFwbhEI+
DJ2VaYoeZHj6HbElUPv40/7bH0qiuppFXe1PHZSU9ZUhxuhI9252JoGIcudpMBIWSNfnLHvp77bd
DsJHgT5Nd2yD7pzFPIJqFOC28HQm4qQ1+07/TgyI47k9FW96z/ENhSZtyAvRvQ4LwqMjfLHu5ZdU
DhPfn35gEu8Qhabck9cQCK46gN2u9FgXgO3N04qyRuzgGbc+8uP+VzLyUHetIudh762SOIzs4zfI
bnZoGMMe0t98XGCUPajbYW4ZtMoPNcilPbzaLzR1eoOAqPMoBr8aL12G+zgpTFntqdqdsrPWzwoi
uFP63NaxuYKhMOuQObiyHDtwOXEeCYlc/KbnsUaLpEmeHFheMbzfpIZ7iCdBcDkJq5rx4I/cQLMb
YhIbdeN7Jm9U090KRl0SRB5Zi3FH1QafOJW12IEkXECMFRkR+4lIbwFeUSNKbBoVJbJZ8zbO2wyW
eszgr9lJrAKSHScOFQeZChMT3HYCP0Kl0h4bxLqRpnZP/+aAAWioTErVE04FDnFj0+HaVLc5Wzxv
/vsMBmXfM9tve3kpZW2E2kjTKn0aCldBP+59UvjJFQnXcC1gwwEr+BAhoFoulJ1Q8oEEaW+lO+h5
bN0+J6Nf9mi7ypMicGJ/c6enB5czBzPPndnUQKRq4Y/sqp9wmoWwcfizxmOSP6UaSZilZTH4Iw83
lI/iFNzbl58FvH9GnltvZNkTOp9sHW7sZjbz2OAqw0LVmha4mi8S2H0K1IXHHQZZSsw9/KUQowQC
5MCTfYYBdOIBd4SaS7v9KME2Edqiz2GT2rBEngiRaVO85oP7xQaLRtbKsFU3O0xfStxNueLkSds/
klhk2qyJUjjU3jIOWqEjEm0RAN0j8qqz61NLzpG3NpmJx7+YlVQomK/sPdbsiaEwt0spzHHG4A+1
tDdBfdGsujQn/PQsdN9hntuoN1Fm8qhY3wAuR72jIfV88+UCIKIm2HUCcwhaAVp4ZqkiM6U24bEz
RV3EELEEsnJcuT4qCZVsw1pPpdORCXy7uokUG1rNR00G6XZzjTDfdSAaupQkVyM1PxK0uQyJsCYr
JchMENCL85g3RcLUILYIHrjtrAjOqol3NfaKlHILgNWcgmupqFSJ+NM4azMkvFxt8RBH6nxnESyv
4gALlkbXsKxdnLFaS+aFY8hldXMx2oVKZ+QqM3AoDTod0OG/lGuoRyyZwb0LCR9e71tXxGVql4y8
8vm26xt87Wc8m+PRMB3+LB9UF0YVVwjQB7EfHvE0IGJQgAGu6PUy265k4GuqsgnQk4pHBPiWQ//K
28gngOqzou7MDoabMdGkfnxaHvTYONN84NRMBxziC75RY0M7rFVS/kvFZuMH4E55GWV4UIxKVZcI
XzliNUrv901EiXf273oR2cS5J/82KuwlVd0i/rjVtTMBDExntJnGu2EkXdLrxU/arm6ZqZvcdKu5
sU3vvBLLKWXx0te/rWCiMGXOUwg1zRmla4IaeziOKWVWeR2UNprcIiz24bGqDdpXhGOefxOxsYu5
lkvdUfe/qUQXeOt7hAM05Dt2PLHhR+3kz0azHnKV7RYN0R5CK3OqeDMzALdUKPJUVGsAl+6l4pTv
C3PKWm6z9aILgjvNy7/gE9BdU0KT3WsF48WWufDOh/rLbtA30tf2xcmOfpxknZs4/T364ay1iouf
40BRzv17/Kyxx4A3CBvcBtCk6C52zpOh/DjT0rhBvKd2XY1CZbJ6hwde5aS1aCWvjenPeUN+e6DL
lVzQG4+toYjpBHgfKI7J3C2MLCdjFASNDSbId/wSGUQre4GQUUZaa/2f6QOk4dPrUM8whUFzTOKt
7s32wweUW5HwryUX5oMqjJG6ISa3B2RFp+0Oo4WSQbfS9MJoNXWGyAamxsbPmo7EhhNiJfvEHvwc
w1up3UoojQf3NhTyD8Fcdf4G2ikNCvLXyhsEkXOt0tVlATEKO8OVqeGc5W9LTBeNQMznWF1MADh4
KOhWNkH9pdUssDbyAyVBx1VAWuaL9P85Mnc1CI3JbQjO1LGnMVno0y04lbF8tR5IuGixQs4tBq8p
mZl2wqZBtVPPY5nBoHsNSHKLMtsWxNmk/UlSChMnHqiVDRXrt23AaMebvja68NY8mPFpGYcqzryV
28/+EpBGG8/DQGnx1YGoEWgRl+6nDvXaJ6s2uL+H+uvtdf9XYzstQLWcbwjqnEbxmF2zo8t3bXrF
xidtOXRcgFEDipd2tJ0mxAmxxc6CtI31ENqm4x4dBQ8qZ69jkKmmKsp6nu3gk9gU81+ruNLca2he
6PJ9+RkApGRYK8MdLLiRMRt5/TlY8EHaOhDs+wcuAlZ8DPR99MDrmZ4mJ9/yYozehHzdJYm+xUkl
US8MIQQrfY2k5FRJs6Vjc4eKvgwovD5N07nVT6mBDTAS+I9V2gNrNQMJCng5980qmaQA12CJIHsj
gGknsuEuDyLIyrgG6xcPBFt+DFIuOFnL/Ou5i6TzQavliNAkAmklDwp/UwD6FY0RmJ0H3fIuu4aR
yiLIPRUb4ojLKeeb6Z35cUNYW2nmsrXaDTUlx/+ebhqqOpTJNwBf9O5mhKsg5kL3gHDomo8Xflxk
ghfevshbd0eQGcpRJxjNTDgwL3xZSh4JJxJl0Wfu9s8PIiTu9NSR5W+XC59TADVK68r8ZGPscCJq
XTWQGCE0WOdXJB8J+lNzRKDQ9zWTvOrPfKA2JT+kC2vAtgDlM8od17jg3cVj3DfAYaUkZnahft5I
XuYuZZqnYZT256sAkPcXi/3vLY8R8CLTEVNCJ2WoyPJgFZKFtndUmxYgB+Gl2Y5Kl+ZqRdfcjJ/k
tHzHqxMGMssmFUzrTEKcb0CZ+yhuaCpVGKBEnajmGti5RwgxW/i35D8514KpcDO5Ib2YD0LfdgAv
qZAzz/BjBU6oRqVQkwWqOkcIWWox8SQYlHTHKeMzvyz0DW8zih95tqjam2Y3UTaaoceO3KGR+Flt
sOJraIsoN/lEgprkW0qXOojq4V/thlSGDqgt3isr1/TmvNUck3hP2Mmyj5cniKaLwCi4wkDvuI3+
01b1no+W4AhseO2jj/hidYf5+gnQRsuC8nknxQi+/aBOORDU5IHnxFdSjrr8XSP0EGrzPvFCUFZd
s5wD3UxGLfNGqbJPIncVhoPk6yT5yAJgxPAab+AUhjRmZIfAM5T+pzX5sQAMpdke2osFGLJqC9Np
F8DnM6+hBghmdLC/TvWZaUqWZtZpCRIBr27aQX/WEGEfNpBBO7cvvDO5YQ7NXOmKRugvnXJ6MvKr
k2JwbL87i/sQi7ESWf2U2oWw+aL1nee/edtHAdAd9A9ayNOAtxp2Ki64cBPgqdz9Z1s8snYxf5PB
u4Tvs5qyufxhLJ/lzWvfwp5I/bxTCJIQA2u3TOLLtgIZx5OMck/2hEu4z7CixVHlYXyd3/pcR4MK
19Lr9aDv45oidjhnAVzGCZdxt61RtdyBJbGRLu3q+jm/wpGey6l7354iIht7shBegTSgFv26Vl2U
0m1GjzF0CyzPLaeOqRPL36f4FUeIOg623Q+tLyAB30Rlsb6AgrdNMvIlYoMkm6SUlTZPcoStMVmq
riaIBvVfjovzwBCTN61Pl4DX1oY+rU745q37J+9Hw2ju/V1G6k+2vYfOdqrKkotqzKvs66BHyojh
x5EuA3oD/4HFz/+Z9KWPQoObagSNazPB1xdI5cLPCIoPyWvXeOv8L/to+StCVCsU+Hp2FdAmugWv
6USRQOrjgCyIMGvvr0kw3tWeY5e61+cy2L8WAgdi7DiZaT3Q5y7FMrC3rcuo7ub7K35G5f6LWhTb
tBUqDSH6Y6quPe1fyBIJ2nHqUDMwo5/1L/A/JjTLVzsTl0FwHxN1W1HfumQnxoLvevA3VkKhaE/x
2n3K4GV2/t2ObOVvpM+s9gN6gPfhux2zFYl6Ke89RS/tadGc6b0pgEm5X94Kv6pPmDbg0G5Ek95Z
fhuD17xUKlbv6KMqS65UZT6YaUlDf+w0ei3DW7ZXz7RNK6R0L4oPoMJHYH6AMZvM25fOfvk2eDn1
Oyqv3WnCtTJVhxlfl2w0ZwlmBTbpI6UnOT2pgVGYHxI3Mp0FxHTs5dsrrIXlSqe+lbaFRCPUStSD
/3khxxXVNr0LgX4uNiLyWSI/YU1WfcKx6AO840h8BDeCfPAOfTGqX2ekQ+5I0uMtlCbS4LVaneEh
VL+myFzA1M90pit8YM5CMcl709tcNrnHCealhqv6tvdhjH6QOQoclptkiHpHWOOi5yxMe0EiqPhX
xtc8txJxS3yWwQUa8r1tvvDWBXLA4q+Rkj9hVosLRsjmTLIJiU04ZC8g79kJsnQyBbkQz/lpTQyL
ZNI0EzsXVeKYwWZ8Cz3NgcCWRxxAfi4O3F34ub345LWvIIhN1tyj1pRtLOksd7DgfledPe1Ojdml
plmlNnHf7HJ8Ke0+mPN+PwM6j5A2ESnQUOs57DD47oLGRVWHHMYCPa4ohYusOmf3DLxXNQzKyOXs
uw2fAxzyKE1J3+GFxmiTHe4i8P8k3VkpXW3oDaibxV2+nNpS2yG83SAZEhH8sCDb77sEJ2PQ3m/i
b/RDJIfsAXFktWCBjL3bG/VraqS7ukQ+pS4KlI9K08ChPrMQFeTyJnduCR9xOyP3sFjeCxqB39Q2
3XTDR+MWLfQr0lpVWC7RK8pJP/abgRi1dkJ1Wi5duuaq011eBRgDYK61ns8brjmbpzM6tQ6yVo6e
jm3jbJL9dR1PFkhvs74y7CCsjkRCjMf+rZHtPrGDY8P9bkyC6nIg6jN+spusG2O/MspElmhLZefh
u/8nUA82xNKkM/CHXgKLiZLpeOaTHbxV0qt7JfuJW1qazbe2kDodHb5S/X5B8oxKqhUnyh7Fznvy
OkLasvRhKVihBz23YMTjoAIkOfzJAPx5ofHqOnPI14GaJ6LVO/XeLtgT0ZWHJ2A6a/q9lOMY+0O1
lW5r4o6JH/DMOMysUTX9Tl9OsiHeDbMEoPs7PtK7/Z4ngpCRGZIsLkFFj9Ek0nTHUQOzVTWrNpJi
IFBtctVRYt+vZ+rKxaAsqyjkWT2yx4tykgD5m7Czdcj53MXQuGxdWrEFTDK9orBZee2s6+gJ/nvM
qbugnN8bYa4naywQ6cLUnUNPgZC8NqV5mqElJvx3niwYIE4RupthcZZCuhGetoDctm+GBPTq/9Q3
IlJC2TcX1HzGp5s1IzUclOpGSCl2fi06hgV4adz23NwJn673eRDjGHCCXx3QHcr7LrHBa/hU3oI+
ZLAxmndig0XvsIFwQ1p2u6GMTRfVPITjnmi9PM8jMmFsT5Xl/R2zG4tWu/4xDqzZJvPlQWaBzV5b
SU8xkc4FMfDkk/m1pXZl4FcOlVDXr37Da4umcYhGcatsrFfW10ZAYSUZ9zUGW7xGdsxRS0nOMrPY
n7tV1hUMfEaluUsezuSsIUAysYVKjskxTgUDgqcqIHmlL3Jco0iGsKyagjdf6eEMNeIyO/L9dP4Q
ZZCHxp8OmPiyXOT14a2FpXXtaf9CsjbMSaBzOk6A4gDpNHVb/zNkz5OBPghYFoEbFogNp05TIEOO
QZmvSWUv2JjxKaTUx1cB6FBxGprPYdISqUCI4raLFQaptCxARM/x5bhcELUBU3XJOyv/GQaeqz0P
sz+c8Thvs8Hlhnw2P0noRezgitgG7xOlk+4ZCb1bNAiW2NpZ3nIer6L9YfnoiafnT0wpk/pht7k5
hUNZSnorkmZ5Gyer4N8PllKpGu4q2L43c3wyHS66tcspfFlVFjp0VetX9uMZPZNhczMkbCAokHH0
0HiwbT8RyYIS+53HILlMmkPMSq6d4MwYTpTr1/UfZunD8MlbF2yBPRJOouZ7DcaRrDo3QOOPAfct
2OrlSx0xBFHiSs2UpmNfWKithRf4iAdydEpbffy+DBbIFCt7OsSA0xc47/gQLGNy9vgT7RToGxqY
foIgg5OI35deAEjqqGqj/Ld2OsN8PaRYAr+QpJ+mJNYm6g5L+rBxVMhKdqLA570b4dKgD4RN4jPk
2F2rKjtYLj95RfB4Ot/4526RFrW24oMNcw4Z9ojzTmN5PP5QQHP1CDm/EReyzZvo6mWTQszQsofo
/yJ9fg/fKUWQdY+W/RMv9sZWE0QZ3DSQT2f8zQm5v9uJyOklBE8vRjnKECp7ukc8CxFQOtYcW9Ig
ntAKvFwyLyX4VPwSIuGo8/ok67h2rWfzfCVj/31XxkwCJHLw6jEXAHnzLQNjMO6dt7g9bzqTP6Le
8OZic03IL29y8Mlwb/b+w9ty+46xpcsvWwMCG5uLxVILudSDi2/wVMbmBcw+x7Kp9AwniXNgWunZ
i6y7lu5TmLNtegJe6qDT3z3f1TQfee1gb5L3dUBTBHb/jGxIAKNEM+ft+FLZ05kNEYLkYBjN0NXO
X05bE9mUc7dQfkkqAsPrUQg+kd5NtWUQdGVM4+aeX6KfYqxbbQpESQ7L/uALiHCU4L7p31n4PIQd
rQqczQkQracYf9VRU95e+Y4MctLiVd+zqxwtlwx8qvFqC4zs+JQck/KG3mNNUKm2o3IbhcR0C5zd
AYye8N19ALE4gmlqF7fmBbrIDgj+VcVCvLoLrJNkLzoMMn3GgT9bQ+kKskoCdFYFTWrP9MwUJ58w
I/YLAMkGeXnKy7Pd2dkzbu2fH24YO22nmZD1qSunsV3IDO5in2nz9AlwcCOf2w0J80cJvUn4KBxd
VHS2pCxar/A2CACxFFE1AUlMcrxrBshzkqpsmkFnqt7+hDYTfqntfMieCIcXk7iLEcXe9jc8CKOn
uWOldYSkIDdHXVp9CfqAQ4t5MjJuuWQvsQEiVBLPofy9Vwji67i5G34onFZO924aJ4HiyZkPrmXB
rTXrxXqK6NOKR9Pbdnd6zqCqgTMwDC8kg6ITQbAOXnhYg8vzXEFzVlmiApC9AdMDV4GZEMn3Zlrk
SekbYCMvbJ9c2kdjDOIhfj58ZNTb8JGAcbJ2S9IgHK68UM+AQNCJ7TFhSDgI7cZze3OznK+LiNam
x2DJyaAR+KLZw3UlMugDALH6XFnXXJOcDx/jOLmDqW94Uh6/a2nGD/HZXsrgOwtHAzAd2FRR3oQm
wZbIhlhMd05k7LTZM/JgEZDm3AEerxnQKSjJZ6ir3hyVB3e32Nm6RPcqaRXAqmyjfVHfg3ynzqUm
bdCAGlZaQ8WpCFoupXChFzwqtma6q26KO71TzcoYrZdI4pNB7038QBX5XpAzoE10nvVQjHq0kRqP
mVa0vILtEEB8SEbx+ZhujYJA+lMPnkquUYcXXYCKMbG25/hjmIdwmI6DhVrqTpRDO4fkMBvYAbY6
sAcEFSXBZVUDYDa9j018yWZmYdYVhSFZHG2UW5h3jK6b7EOoSdMnFV+6yaWdYJnzZx1THUxb2pDh
GPyGXN+XmjFMxG72zCf+ud0eIj77EjhYpH8y/29PSsRfGqYz/S4B2R5ngamvd4c6fehaB2cCcZCM
dO1hrFy00s1GhfD920/CFVi9JTqoMw8U/YAIF49MKvW5oRBv2Ylb1RAArRVo6jQXhGDFv2q8ZEgu
/X/vAg0vIM54+hjaA28lw3j5xsSsyp3eV75zk/x3553r0Uk+jEmjUahGtQMDiLfOCXVsWXbRmqD8
dcbqHZaERhats929+AtrBnC5GQFmfiTykOi0gCmmagJOrFXSvD6A4h5kn200A4ZAmSTh0oCgTyLM
KV/FQtH/W6f0kFwxn/mFQqMptsj4hGjbSLBSXK2oBVs/c3+Xmo5KGsrE3/kbkUSbb1VzHYb9wdgX
XYn752U2kvGVRb1TNrwY+Ck4ADXrg78ZPInB0aGi+za2oO5G7ChYfs5vbiB9GBqI7Lh2rO0qRMAz
FAXtvmKduxU29WvKSHyHrAhe1Uj8dB30DYfoGysYx/0b3WZbRFoi1XGnDRMoP7BHvy/IKT6lsA1H
Vo+wvi9NJ9vhreMPxTwzHJVgcR0JkO3rfZn5sdjQW1a9JM701Ssq1oprVHw9i1pBM2BzkvygH5RZ
Rlb87CdkHD0ZGBHJRPRVTdOFv+E5d5a4xKUkZZjPgS0HZjJWBTEDBuD9rVzQe47584PGjJ0oE1rC
x+xb3ynf17YILRABNS9iapDXAygp5jvBJda033kcudkrPkY2P0Hdq+iD+Tutqt5oCsadJWwH2tQz
UFjeA5IdE4aELFAKt0+WGvncWMDkuBnCGpf3uL1WgonEDnw4DV3A2qxfPTvXsjHSYwfQnj1/9DYX
bLzNw/MGpgXWegZbMwa3VDul1fq2p81UAN0QlVG0/Qqvi5AUvCFmjOopwMqOSG9nmg6mwhGln/cF
rxCsTv3gqRZVnoCL7iGFIb5OCucaq5OTJYXlcBUUkezM4rjf73CrQKUIoQrKZQxleXvqmCVhF7H3
cKH6MXdbB8JEyyDXKXqcyWNM44zdlpRVpe8Y246HzTVlx8lS4WUvZvRDl7LYq/CRc8/8G0+g21Sq
kZiRDsAFzHw1uFGFQtCBoT8jTSx8DcWKhBek3cbEG8EQZZ0YTOlnJy+AOnftu63la+Px1xpDmBu1
Hv0uf1s18nJmNEd+ZgR6iE1wjlqP9ZofuWHlix9thrVtkSlkVcB2tl4+/yTTRb/u4bIfJ53bOH4Z
NBSA7W367mmiHdyZ0rnvUz0WJrloiIi+LTLy/Bi38CO/iiqcb3EwbLv6FDMVbR0R2u4mTbT+sx/4
m+R9s5ftfDklizdrUKXNK6MODfdRDYrtAaRCDF8fuF4NdmziFVyIhDxXT2yZf0F8eyUJ8N/x/jlE
lwTrjTnabIlkx8NmPTLCmtfWwCGPm3J6raD36PfZGaj9gNrT5tNWRUyO/10OocgII5CBxrG658eB
yLZgVtITEgPL2J3EcIZXy5v0d2/frdSBwnKyUH1nvdDHygdSDVugTWtMuQnVfSTs9iY7HT0RPwvv
z6vzms6djMG1Oh1xWjqoRjRzp1Z3CDaMyup+4XMwkUPmTQm7fmF9mXKH+vGM2R8+E+rjf+dmAXtO
lsKhgjEZ9QZvKG2RTzy9EymIJpAZ8ndoxtgSkIcxf6D8nhqXnPnPVYWuj2CubTZv/4uSkZc30UqZ
egx4pEz/re3pLXxJLg8gyyBUScQyd7aEHj6xJ2wSiDKh7Ik6+xsxPjQZRpvxXUHCiLOwpYDcHyMU
6rqOD53nMV0ImJCpyBl50LXGte9AaYM7StjNqLbgQtKCjS9vLpsr20hx2CBTvA92sFQSOBYgn3Co
f+oqA5lZTfvoddz9TH9sO5obb+rpL3djL++Jhg094U87WWtSQBV16ju06djGBsvUZkpmSVCtnFBD
wV9rkQOx5F46SW/5nTfLb4jMiVy7xwGOU3DPPm+oRMCfeNyVpUdFua5ABqN0CRfqUvFyPx9yPA3d
Iu2HAxF2MdizzNRhfmhd5Isd2fmnUqHB6f6nldWFrvlZea32PYCNaqY1WXwgDlLX47DesmdSA6Sr
7n8OGyN7oV6ECCVLg++srVMNC1Uro2idNZNe9WPN6hvzH1lUtcxULbt48bK+uhvcyFK4vY9xWids
FVYY7oNlzX6aV1oxqNFiKm+POopK0+RrhJlrkjT9tQTVD46TQPSaMsrW2JsuxgnFwqqXhLvpegQb
przK5Mm389UjmbcMgjST+St82Q3t6U09XH0T1xP2zgopDFnWOjrlK/iNNXqm9K9vTaH4kUfUCAlC
+t3A0DWijgfeaFl4Cnx8FSQ7o5X8yxn/Pps88ZCnmtunnZ7E9g/Fn9uKjn5bRltFN9kMitT8/wAv
H/YPa9Fx9Yoi+YVrKPDCT9C71amkVYGwNi4Ab6VVHk1SfXObFq3KQCu4ssnjqKU78B6BMtLkk4nW
IlP2nlVqOBk1vlFBVcC9YUJU3nyrdQ6JwT81HZ/Q/Q9L/VSk5GmBq5GpxWgFMM50vr03e8BPTynN
jb3V9aKkApGVMM4crG4wqONi8Kn0+XxpmSdek1eMyPe+9sGbqMWz0Z59njQ6IfSSYNZI7aulehwg
Uzw+G49tNDeA/1jqHJ33ZFApYxJVRasUGvV8nfIMMHs4iFKSDbxArukqfCzgAU5MlOxJY/L+Vt78
r1Di+4rs5YAtPiicBN20gSfcAODZMEcK0BhC71TsX+yA2QhsWeox2c0US3YCOMJ3sLmbJLniQuoG
HkGnEx45oyvtLuc1oNUzsQM/GMw6lyLQv308LVfSZi1apNVAUNDBCCvilq0+LD+xoVGHSr/Ij1h+
GRXV3Ps0HhuobB4O22MHHM2BtYXsO0TA3KfVUO1Bts9NXAnPNGU4ZEerDA8AdEl0t+qCRll2SMFw
IDXZ+n3yKrEhCNpy8F4BwQe7iSlwuXDO68nf+QMyWLWE/qeFy6ozuSv/lePBV2PEbHIvL0k50iJ2
zf/b+CNymZkXGMZmqbBOSuAY4KQn+KD2+vM4dgZam0JjkMdug1vGPEmvGIxb2JyAWDGR+T0aOGOH
CLnp1P2EDrQGuV42L79jlYzASatb0zZjNJa8ZAZsWLonRgiFmMEjbcdQ553y3PrCS6ldG3awEvNg
xONRRXc8YMFOP+TXrPBBOt3W/Jmge6W9+UBYmiGWZcO87840ghD6GLLaIH8iaZRABO+UCcYRLvB4
3Bo2m8gk/4FP6esVToG+DOoWVsu975MgwZQPJg3AsoOFjBCdCBsPIW6DsSp3cxxdWSVXm/UukFnA
YGzjrdRFpdxh6PvSy6nLwGnbydK2oMVWUrfOygdMz4ryt3+kJWGauGdlTURj/Ud2BaTix93pzKM3
fEnJgV/XahA2/paBalCS9GiZWycBjjS1vZHzs4H9+LXg7GVFW7fg8ZzDn6ozDH1lws7vImfTzaAV
16P36O+n8Ak4QgIIW3xK3hzsZXAk4v35QEuhMMp2g4NRh5+c3dQttWQ73twOV8stt/vh7ratsrhO
4sOKHZRgG7vDF0OP0jAP7SXw/m59wDcNn25DHJNCwkzIa8Nb36rhbbVljZdEpjjNq1oUkTq6FExn
LydlUJH8LSAyk286mPXaQLVcisRpk55ONXktUeO5BBJpRV0F06z8qLsOQNLZ8bgUxIfFGq2V7tgZ
LPQSdOKZf+63ADpHKNvoyS+/gq16AESf9Y2jSNz9V0JDB55bw4PXJFXTnndPyk/Jr5Wq+KzGi66X
WlUJ/EqlVteG1l2PkIo1/LvNWSl2Owx9Hg6g3JvjxIAoHEXYVH6BKZOwHBrb4VYMfztdSKw5FdNv
ns/7Y1rES5UYk4/ZHcH9d7R325EEYR0ATMZySQUoMp/amS6iEj4fYT5PiIR8pgT04Y1AQVBTy/I1
7eqSbXb2XYYbq8IflnDWK9qNsOg0t+Mpn0ll6FpfuKck+xOYDY5R7RxafI8W4xVGBx+f42I5ds3y
Y4byTbKRaElFQ5PGkoldUCRqER8+qxKZeh2A2E6mjUU4YrZZmDCnMBHsvFOmM/l3NDSskPKDTsWN
sq/CSfCgixFzob0BoYqqmp55H7T6rfJZpDUgRJqnfz+Ewyf2aW1Lj6NUGtgBObyGJGyw3nFIPwlE
8Q45d4+VqBEVO1RjfQKrV1hkL6psuskPKAo5tbQHgioV6ra8DpPFWxWZ6Tp62wrg/5OmnFNLZx2W
C/Uw4y4pdjO+NXCdwcQVCu8guA91CjCm44ntZBl6lJZVeqaivWUMvkXYD8orD85/RNWmCpdN0anw
O3oZHtsOpi1h3heQOldR5RInIl1L6ieuooHXlrkkc4EhUI08b4dXOb3XEbc1zHBtKjwStATNg9fu
mdXb3OkZAIjwpQ9uUYkEznKTNfe+tRJtI76qEzKnS+6OzoOg6bjwUFQOkBx+FOLxO+ocV+6he+dI
EBDzPb0dTwZokIq+rE50aDVeBtNR+JshqFtgcUJrbED7LoFtMJrBOZC8cyC1rwrGFB01izIhocxF
IJ1jExKML2IlnqzwD2Q0ckI40fTZEMXdDNoOi7jl/OzcomT4spaJFT49kOl2vjy6R8aB3wTg+Gv7
zNWuGES52jVgJV1XIHid03RKuuCxD6+Hlnus3QvaP424T6ITZ1nlBFC9eOibgT6SslPKTof2Ss7M
3gAwtb7169W2yMecjF9lsJMsh9kL04ukE5hHCzAs1NMMCOYAoRoyr7KE7v1U28y/gkF7ydmuW2i5
kPa5FlpCeK/0fjNL8wUjna6cGE2phk3q5dGkzwQk2O+/5+eMnOtCmTOiPNUMaU372u7+7CmFftuu
33LPgrAH9CiZaa7Kbv6ErQp20J4sRVO3LRqSvEXZQtHc4o5FPAucmWZLqZSIlxE+ZB9hLmnVJhey
/Wx+ZxDkFmU4vUxubfIWAvsnasF7YO+DDdCIcmpHBnZZAQSqh6kQmmTgPgmRcRTGKHp4hvHiBI5o
qE0G8VAL5sPCCVnZB55IBD+u6wJub/uso6KMeNH56Y4JTIwXf/2z08WKWyPBO277MT8hAqNxW3BA
p3+TIiTk/Y4jv50eYgXmZVJiyOQdni6daHezWwCs+euL/Z8sCJ/gExbxMGuXTo4dEvRL3vvHcxhg
nJ4jkeswpqpFkufxsRU2Caitk4Sda3zwOMX4b4Xby/naMPfnrN2AbHmoQfhuOx+qIsBB0FaMJ9ib
/mn/T5JcF+/KrEm+AAgPNxVo+atX3dIerZbQvIkzuKbvi1/fwuEekrKOt+58sNchIHS18e7uB7Qi
Fy6laSmPPnov0U7h689U2kIPiT3f5sT1eOVKxMAqebZ1O2uKI9aoaYqkygmOPpMsPH27LUeJT9Na
DKIZyxu4BZ9hrQd0ZpAmGS8Cs/YzWrE75vNjf61Y3lLIwj8oG5FqbXOokou7NeWGJz2CUgmIbCst
WVCtIGzhKn+SYck9tuq1pHd6P1zirfWso+v2qXuGrDEAfwvEyde5DII+NhiSd2/3NOHcYbcZ4+ny
GP7GYc0qQvp2IKB2VFsfCbZxSMbjDdr80jgi/FCzrx3ElrcU9XvG8ki39eBVqus0QLff4f40g/OI
oNHQrlXI0JnAMJo6leeJKIIEdByeNndA1qi+o5m4LkcC294g0uAapBncUlqGd31m9/UW8OFyBo0e
LCTJPuxbi8+GMgOBAmD5uZMEho0K1374bbMxAEMrY2IEatRdYHF8UfzkDFqrLIPqitKQs+wkWlG6
rx3LtHToehJ9W92MV2zoJafhqgXeXa/5ZgmTeWkCB9zd8rJv/qp2AWjGHwUIW+srycX0AQAxTL/o
EXrSqDzgPbXCeZxbC8nMOs8PPDoCMakl+ImUpvsqv+hLJ7nNOhbRaX+lAyrRWsOHAn1x1wXmuGva
N172mrkp62m/4XN5XZmamCvvCyUWeAvqmNAIk2nBZOm09Q8pusK/7qixFiqhY+ER1tlzYOMmae6/
flNx6HEPFt1zzeBI6bmmtGxklWjj3P55i1aYdd1VEJhBKph4PPnwdLubbbiAnC2qj4/YFfevxP9l
x9rkxrIrmgSuDywQPTqDSZsGTOwsk86eYeE93y3CrGH931JVQHcIzn2KkNyyrOexHD62HRq/fL4U
Y4FU/NeFA/DGP/T3WvpR6jvB1C9H4A9PNsAI+B/CAFIwGc9gvceHWD2uPxkv0CDgBAV9gVCC/LKn
2s00WJf//gpUuN160hHjj1WzSuriQ9a0UNBZ1+AvROY8L3kypg4yJl8fVLro7xkZqglbw5YnhDXF
ZnYzQkhEu1mXqDeCPfVj3SggGga223e9SRj9FiD/dUT7QHWAwb6mO1gEMJ9cIf+cMsqH5YGO6sT4
c8AFUWaFUtWli1enjRRKMizWFpxhhrh+9wW1a5YVht3ovVdHbA8wkCvpYNkegfmoJOqEOIX3PAhI
RETymtWf7T14AdoxxZ9nOytlFQdV1zQTtfpt06rH+mVhmzPs5tQ2zuSa2dKZAM6NOjatbFlmfxWH
1tG0/4cLnR/pHAZvMDITl4S1oFHjf7PduGtN3GxVEbvrLMwFdBGl06rDnyKyxrXi0/L8upwmHoBU
0mOV5Bz+ZTe6oAR2cEZUJpT5adAvq4gmIJxiXUXJn8qYDCEa44mfRu7Hw/UMw314C3aL2ohW6MvH
XfltCxm154Y1omg1y5DjsGFxOQmcdQ4jgIgcQu4a87bjlWL8K7H+txo2lFvdZxqSHNuKaJWj7jEG
SJBf+1sy8bufF/XOm2HXxM+ioH+oCd9kkXfqOmsH/zzYiZtA5xNzzhhgC/lrk+2nMi8DHYkoqiq4
uE2/PILiDajzP9CR5CPwbKGvRq03WCuOdunZUuOwSdAfkhm/RoLgsMwTyCBWONgL4cdXeROt6YmA
FFUjTXXEzTRVhTv/r6Ys8/SqRaNoyVmcqKBFg5GKJFY/krDqtTygZgxEOuZcPf5dwd+cHweGrMpd
RLLt34V+3IvpgUF57WRsNpCG0zAIIw2Lf76oPky7/rdQYZModUQkzQ0ZuGwZA4+pRN1DOGf7wcSQ
mKoZJEFYgcHu0q3/guaQKhelI3Iy+34/JxkYD3xMOxJvOOBaEhcbW1kcnX+5JBM0OOiokgT/sD1t
RK9CkGo+C/kn9KyrnK7ApZ29y+fy9gVjypaNXjWfGR3BcsQUQMWeqadOJdG1rd58itup7dwUaEgd
OB5+gfLb+VUx+xDIoNodH5pHwTnHGSMtT5nFfNYBFCgC2G2DM5vWS4Rjw4r14JBruttbJMS+SBp2
a7vyP51u0PRSh8iPmv6Rwf82aBdnlGrTeKOIZ2T8wLSNKzjoOiMthHKqGFWjbzepD4Vin3nkHmIo
8CLoi3LfbmM9j9DD81IxojVSSp7AYZS7SR5OCVEy39xmFl40fc3nvtqXS4P6zPHqpAsfr5C79a9R
7p/5Mc1BDrnu5dTPtC2eKh3lFrsrxtDKtg/eKEkKoeMVEtc9+2vyAE1DeL2o1aJhXsU52vLVw+g3
G27DfK4DIaXx7vpXiPpjXDmNHU9vs32aaHgDd6MrVaLfWRZH6WPZtgS2gt5TVb/+4IapF3fVPoZ2
ZtY3vb0zkss6ltg0rMZWteHLj14YbPgKlEtGozGL65Y5nl58gDfVrrzlSXshPeEdfAFOJMqGzcR8
qZ9cuqUVeg2UD1MAUmd4h5OWeLmEfc7GSYEO14JJ7Xwlnv50jRmPLBzKs0u4fRmdRQXUEl75rT4h
Fz3YbC4d2+CTumxLSAgdeQgxHU6cjoxAlXchFdfs3dZqPlmMrvdLret4WE0R6p9AAJ4MWOhlfPm0
Y95pEayrqiySsFRYyXhwWbvQFVvczotG9zrN4y8S8i6686em1kaFnNKX3ugnEXu8CJfmj7PPkgc3
ce7/7aFHR0hgjOEGfSallU+492N0dw079uEi7tIQclW/nsNXvFASByQ7qK0zWZ3i5fSQToo7x+nw
PczVOF84RwBoCs2S6GeW6gEPOaqO3PxsGzUEk71JLtvVMu52dmKoB86pYn3n5JYKaXw4qsGx2Y27
viKwPqwZgMT26vkyin918jkjiADspfpgkPAIhB0lGNYQGKPhECcWYvANJ6aYQGQwWqRz9cDD/rGr
m2R6fobqHRZhUCzT00TPgUQdutHAVtOAtW+HfHeJ1oZnOPv7SnZ5vAvBZK0/ftGIW2yfLFRK9+jL
4/91rlwx2wbFbHCmkHn1RwE9tGnq1Y/WkvfJbPwcta7J69kas+vf5L4PQjzEcQeMNVFHyhF/sLAe
jpGon2iFZ+ZN48wl7hg1hnQjJFvH4KxEB0Za5/F36NHz9YaEhlDBJ+mMol3J3CV6D/DnRG5/+llV
+b6EmWEkFJHkus5XIkEX/0plFODC865WgwWReQA3modAjt3KAZAKcBjRdwF37txixWTNwFAfdQRq
QawJhk7TTDNmSIRgMrkrwLNvr8JYJ1kjqIcV0g1OLBT2QRMRUVyQOrdiGxXYM6RVjVLI9tffaPBF
oinMq8gTak2gAzqsC94CCHg8x6Qh/XiaDJ2usE1sYre9Is9KB2a+Dng5ahpVyRMi1IcB22zmRXgJ
qBqFQVfOojsENg8tF37oH9xlAJuCRGvlcqSwF1nZu5CiYXsVYK9zPB+OwB+fKhmVMrTFLopAo59E
0G2qCE0HUTZa+LpvPW4UbA5WPLaYLfVxOgNVpiHXNkOnHB9NZwNd798sqzN9O4TCAFX4a350tU0Y
UWSrtxh3HsdgYF2RKN4VgsQfZyEKkA3m/1P4GacK/y1bm+hd5KLovSMbGnhQQoxkSqhdN0ybYmf4
A9LRkuwtwESDOO8uIeuxx1J/aX5Jb56PJf4vgkBL9ATC66wQLH6Gl5Al5ZhbuTed1hUPZeapTn1z
fz0vVrktjV91MnZpH8YolDeuWvqlDt3JgeKGbSi+5QQ1tjZ3Mg6ykGJHSARibp42ejj8v04K162D
7dIKZ1K/LLJnZVBK1GiOwOAZ9XmZng7sv9qbrB3z9Cs0aAeVJS/ECt/xsWaIBnJ2993oTo2bN67x
CH6nLHJKj5Q3LJiektXNaM43izVf9J6VGtDIcQAGL78+8TyCeiAJhVdH7PFfS/PwxQpsUvc9s6w1
kzXwB1bVQyNjfS2HIr7P9gG0DPOmAhGtqHZRTnLwhy5B3NAk5rw8YZfhBVhuEtWZA7Sg1/pbESUL
iKt51A82Q2WqaDa1ZBee6YwuyeH+FM8xdyxZ6oWaf8m358iZ6RzwnG+AJ+mBND+A9TQ4zGlvtQBg
P9F9qVWxNqBKLSR7rGL94ZWseSs4QmBl3ZRHrDlih0x+eLAVjEkE+P6OCV5mb5X7j4K9NP/aRcaE
2UV1p2rAHxgzfbaDFj1ob094LwHjQpZ4wEBgy6yq/YQ+onAzLrJHULJvzyAjM8/gHPCwnZsFbK1B
CB4OqLyTfm9G/KfBaztKHnF2kKGGirfOF40jgSm9DVYoaWnazqm6Ho8XbfNsqFMH6y8UuSTC1afq
XTnBZT+PRhqEccanWkZpnyBwG5NpOeB9hLzGqX7iI3j8QoQJkRvbaAN7WB+fCq+OY595dGf3W+nr
+9P+fGgqBuOsoKmiOytK0q61WH8Nn6Bq7jV18WK0ykSFoMUK19s+FT5XqFj0SX6HYrVN6yjrZzR7
jRs77WWjCal22NGarDYfF4kMxzI4964IHBgi0eQQLWtlz9n6oT4diLrRAHVCoBs3RPW2qq80ScqE
9Lwg94EW7tF8t/w1SAep3/QIuc8giO0IriK4WPsqOdcd4QenEOrcZHsNEmq95xEr4tFfpWTScXAj
3kx7DdGSpbn7tTgh6psVlD651jgS3IXsEwRsI+HwXfkSv9UyfDYpbRLRa+3oudzudSGMbH6LzJ2e
neqQygFcRhfU821O+mLw+5P9P5yCKic8E+cOa+SsaSQh80yb+4oIXPrpdu5GwUfhwh7zqANaH1KY
8g99bMBii/Brrvg/AMRhHKb8sZrZXqJICesbgljP3ywiriA7UhCf3NDZjygEQrotqgB9MdfeX/YY
LOYlzNjIqK1ddydIe1eOvKdGwC931cBRestjcOjNUNRRhFE6YF3EjqsMKRftwG1WY9yezO0cJpnE
F2yd7D5feOGGMSv1iIl2fuCRmsrsh8dUeTiFG/ZJ4eCWsMjIUsTPfdzTCRkruNguMdpT88b4KUnp
Tz/K7WxyuO8sivvE1pm1vbqs9AqMWp48SopNn7/ySuRMTtvEOe/wYMAE8N3MbJs27cfJ/KMOxWYa
mR0d1a6TxzanlyA7S4nep1sbGj217Jvk4VAy7bkopXvT4ilfY//+wTpNdXhPuL5rBZJw0cdxfR6V
WsfOohB9LpjNFh38VytsbUgnh2nCiqTBWMsP+y5ePe4gujKbsiSx3+H5v7j/q/vIIev2Aml7mW13
3Dn2SgUQQluIJBGrUKvBaK2r9Qyx+eWErcT7z8l/SLF92cEPuQK/Hqu+LtdCjGchCQuc6Ef1mxGS
+CZUlV3tuTgU+dWBHBVVwvwKCZfRSz5uJYBSAVsDo19aXJ6OZPKmtasVP3XcEs3zjkhLHzASnY+v
Qsq7poDSLH9ug3ktSGJhhIQZNtkpqwjZWUDUNH+OyzPuoUu2k0VxLbjzgHAJGyxNgqpA5mX8TDNR
WItxrVVe2ApTgNgh7SrGHGSt8EeqQtd4AoS8bfxe/8IVjolWU3Yy4ya3TBThRyUtfM8Z8DOtNeUc
VyiS/UChKU19ZYBg9JSc166/IesNG3nbpDS7wv8c40wozJhBIaNSsVUzBpxoeLQOFfIpirpZ+azL
PmGlX2AbGGsMSm28PEIat1v7VYPdzcaQBdvHbJTlLS+FFo2qf11ILuNjvLrJNYZafyWJ9oYJQMnq
gt/yhlSqHapXkohwOZFQuhYTHCLY7CrndepXxaj7veGsryw2y2yAFjK9QmC4VLz/rwgvSZfCMFgC
Weto3TqcgBvefNT+Spss681PcIdn9U4Q+xItj49INIc/EIo2F3gt/CC2x/1pUVSbcZCtnix4OB5t
TRGHG1u+QrJBExzpwJ61XpBGjsxby3xJ9HRUrp1z9XPwtvgo8JF9H5RmVxW5FKTX+H4k2N0pXBJr
KXhSsjBmPkLMhhJDalZPqR5AYcxEfbSC02dT2Stsxbhy39ax7toWwYFGxeKZD/ALlKWa5IcjTjtT
tKDuNOsXO9rSdvyolO4RgwOdeIfacxodnnu7PZ0iR8QeLOBchCIK1pGB3qY0IdtnS+fP9dqkfw8C
udFEz0mE/wPhHhfX81pUlSWDu9Wx9e/FqC2PUb7lH4vAxoQY5mUwA3LfRuTq4/fyVt0YcZrpyPuy
aeYB1F6PyvVfZHq2HTsnWJM+Z+eyJYN1aVWsZqeNoYiE2QmiLKa7dEMynAXksiBwnZVFlnCdvpcu
4K/eMkK2x/cZjfamgZ0lhgbuSKxlJaNerVTOwXMSQm+sS9vGGXdRahCy6GwIDOmrgCxqFK71B0+M
6gMm31gov/oOHullnxGRRAagkbqLxo/XF3iPhijTFlAO/0Y0l9DByQrXxOMbaTbnZcDhvwCS0PLb
Fe7wfJw01RgoAtqwbg8YZV9rTkGAR6vRzj0p96Ts8UXTVHr8DxakDusQ6DvBPIt1QJGOqrLiiegh
NXI5QUx6Rn4R/5uN51QD1pJmXVO0un9+Cd9oFV+R8/hZfLa9WqRgwEk99Jkt+WSZEdSP+HhFwSOW
J50RF9hi7fhAD6NUhlXTpYDoTM/qYeWrk16rpFwEWY7L/jWkvXuFJ7AIdjmQdBgJv/rcPDg0BBgj
qBbq0qgjI9nV5gjC5KKWfEgjg1q1uT2OBxSj/hvGceZF9D9sz6CPef/ZqDjTg3V2yRt0g8bveJhZ
4rIV/S50g+BGGUfyx4S3ri0XMm1kXXXm9U/KjW535mEg5yNSc+EB2zR+BOLqa2trtB0/9e2NrzRX
xBaaxMQLfgQoV2133F6+dHggXcBPBRadQ5nZ/HmL/tTFZO8L8Dr9oUIA3MLMastvyHERz7Hm0/mZ
AqrCH8phyc2qdojs1B9lTIDD++2QjQpYv+nQkhtbzTRwTqK9Iu/9Q67IA/B0gAOdbb10cdyBtICG
y/VFZsqKCOamcoOJYSjxW4EbA7owT6EnzHlyNQZKxjHckXyTs/Q439rL0wHP+dXeifU/lTNkj6bj
8l4bF56B4b0P8hHrEztqlCmeVq3+vK2mkkTrJn1ujIoUCtdacx7mvB4G+iHJS9pJV2aAFjwaY2rP
GfflwO9undYNXFwv4hd7n0MSrUCwz5Qt28JCV5RTax7n9W7tu0L9SICxS6beI4JwLn9aLasIt7GT
LBzWPeJ4/jcV81LaqP/pipzcj4vv52TA3rn7PLG4CzgfNJQEDDeZCXFWlzMBvjzH0n7uWJlOg4sx
+orxvkPNw9nb/mY7z8brUwEo6ivzakAIMtNsuOdh48A5ecFr6dOq181sY9orWkT606Hz+Q37Wncv
fvBSEXh9BQ74VrVPuMkSTAHB9YDvpev0uaUXwIhU0Wc3hOcP0/biRx85z7GKI8E6Y2TbSBFGiZV2
vqWjcVXtBzv1xrOIzNbs9fWXDj3hjnkU3PfzyVAdfaGJhQaipYYzeYswX7Wn5e9hW8supC29twx5
j60kd4kn8SyATZULlI4xd9lAiQJCf5uKtYgb48P/Ny9/4rc9fjDZpYvjHGQw7HVnIzAmRP7aj93Z
vlUegRgVubzidaIaPBgX6ekmB9DPgRoGZTouUfQWsYePDObVdR/+mKmAfWiDq7/wQzAnqHKmZbAB
1PzpDWVBmKMGx4IOh8u/PCKDs+XxVy3oB3s1nblbM/ieaHfEX9CPRVhaPDVIrIyO6YZ4F6uNesGY
+cRrUFK0e6aRhDN5N9AEGCXnEnbkDnKa3cSpZgdWsROxrlY4iphDGi2+sN8PAgcPpcoV8C+zT2My
dYdYX+svahARBp110HDZRk/xSL8yNbuQPgZBFWnC4nimsbkXugQ8ASZKmJ1Ynahx1+VuhuX/rR54
Bnc6izvqBbkDvDU0VurY4pXlWoGuW/QUvpDeFqwwAzQv9eikEYb0AdngiTI5zefhQY6922f81LCA
6DF1N5hBtmGIDgWlzf57xR/tTWgjxv9AgBc3CQv8LqeGG8UBiaZofF1GDDgyIIhoGW83r4I7SiN7
qERuZMHHtZyMx8VyKvPgJnBQnpEu8aT8fS6tWhlkWpNi/jAVuNGcSif5pzJlabIRkTerjC1dTjeb
flJ9Kj4xTYkKy2xDauLGks0h+EAqQHy/ZWPpMuIqcz3mtKCy3lm+WODQA0Vby7Rdg8nXeqZW5A2c
GdlOSRPohdbftUtgd+22nVSOkk6N3zKI4FM7/tZJfl9HCZS/ICh38DkQ4iQUpCErtaKpu/OJD87Q
xixfezz7R/+BPP3TwMtuMCBcAytI/7M7cezAjCM5zKDNXQCBWEc4C+R0PL+W6dqoW2kaP4BZ47QN
IL1ih2G6BqCbDOdyadRuUW6RH26jvbgbJT9dLknWAFbFOl+f314jtPIS9LQIf0se4QYtSGBop/uO
4ZQL0/LSaJOU5pj9HEAn8PiEyYzoRJMeXAmhEiW45uc0e5eMa8xUuZ7di1HYtpSXzwVzIfgholOB
PFX1pJkoUCr/6yg0nTWxKL9kGVNGjrE6aCNfPMo8uuVQpuRouB8UGRpMH54zdR5+MTSNFzNzWJpU
OkxpOdTU3QtbY2fhJKrCENihUXhHAcWGmVeg+HddbsCWF3Ub+atkVRYUY9sTYWbSJesvUT4kPeSN
blrqXgMZ3Em2GTT/6cBUQUetNe5bVlbYvBteA32pUSyl/Kt8jWJSlNO13xd7tJdpL90nGsNNgWje
NiZIB/WUgFl4WvqvyGHNbxNavrgbx+Gxq6UVlLzA68/ExOHOHLx52gsXrFqGxHXPjSkkmv599LaR
oT8GBv117qBSGWebOhOpDwowE1Ywr00di2jDPf/Sin0Pxt9dyKSVWS1GZvjUyEKQp2Dz07tqy0RF
4bAB/X9dKN880aNSCpChVJClWDF3Q6Dx81oD7Q+P3mDN5uvf1GYdPNzmDCCP/N0q4OUAYplOjqMd
eN4Rew3siCSqp8GXJD0IuCxZdjtHXpjqEEIbbc4+4UwY6S0dgBqlTgQEX22hjLU7Okx+8OGLP08/
hk7wYKlZu7SFcZhfIIIiziF50b/a/12vfRohv8KFUpzc9MW9m1tb1EY0VcdOimTIHaiWse7H6ord
/i41KidObYKlTU1/mHqlPfmiwrnSk2MKOSKS6rkPa9/42Njkcl+Btb5QycmvD0UUWzdRrG0qlZXs
txs/iu6o/NFn5Cn+SW8MNThJcnwWalDyYRafrOFJwQM3RWiEOk9C74ef2b4sXmd4mzmMUEh0u0yn
VBEWwBiDOAGPjOETgx1zb8TP4VfDzW2pL8x2p4SYMjYiCbHPvY24XoS+JEfaTWwoG4HJxNN0ZHRO
8NtM6Aam9eMlEewxq8odsooAL4nZeCrhAIrCNvBzRRpylDGYPsORI0aHy/LMVW8sOK/F9l5ZVr5t
Cg9LrY5GE84cg4ke8bvopFQJIxr7bUDarj0aZvJr8ypvX5h/J5P1JH+9oRNnn/8m2mZubGl3seOo
/D50kzeyuoR0znSMKrx7A78tXlESnytP3MQqPaOETsDKmCCVknEyafaZ7Ia82dR8Qq4VZes5g5ts
RmuM633Y1NL1TNqUtoh8xiCGWuf3Pokqmvz2cz2/+96OLmrOr+ZOMKz4dGbZV6BKYfZAN0hqgRxi
6B/1E9PdPGeDpXmfpqYUFOsGOcbdO15kyMUpNtx74X7BYGCd9WBrXlmBVoLve/rMytRk7hhkTZk2
SBsrPio4CXU33YDgxHEeQTq/GtOFrxVzodBIfZw96FDgQbyCv00vNZ8t0b166X7LRsKxsy+Mdk3B
/WQK9SddRsaKvkh4vP16TTTqYWMKYQG4F4UwZRsBnWRyg0q+HMZyJeS2C9z/HMaGcrSgj5bDoSKd
Cvf4hawXL7IuICPdbw6gO/RgSi+sw3cHCzmadq4Yn1JvOEliuVmgRLZg7T7XeH5k4vuOSCHAs1Mk
zUe/rlNeIZ/GKfOSHjtJJZ3/yiNn+tMim+ns2ikue6MFk4Z9Rzlt7W+pEbktI7fGHbVW74aSrEqM
RzM4Tm9ynJu+kYc6+pAy9WiTU99gBtoiP7XIlY4UwYn4v5VRT3aaTYtoqpptOGpIel+DLCN/sh2e
oVTKC+mdRdru0wIPn4br+q+yQF/+Thfux9pR4anx/vu8vfnHWaxcLuVrKNNaCQgvscgDIUTdxL+1
TpVIgUmpnEqmOL6o8rE506ePTlBD2vTXZAzOeqWO0pZJZYUrOQ/tX0rOi32MOigRb9uHvlfWKt4L
eQ2/gnhS/ejEbQhTlm9or0C/MUzsa8N9VdBDfS/Tagg/r6D75QJCLC94D7Kh4Tzs95lkgvJulM5I
cVqi9WUACXOKDhL8WJpviknYj0VWSn+ulvW+BgfdGKeLx3Nl2IUVwixwaBSYm675wCNQgxlh7Beq
y016nDSE6p0qtRm/6e8EuUbDvYe9K2JxqKbV6qOeuN0a7uc9ZLd453gzJ0V1kNmbSikxhdsmBo5j
HmTHu1wD3Im65t/m712FupdxSklfbYD4c2Qn7mvIPBZKzWnDjmnbgcOuJYg6vIPq4WVnEvW57eQh
+iZ31Z5j1tz9g7GtigJm4zxfsakdc+bPDv4p5FoH8qrp885dpkTOdUB0Dd9K1RmotgZbePDbCVvP
5ma1U44QVMncedv5o9LMGLfg05tsUF+HbOuFp46iZQ/oYm73HhSRmDLKtytdwXOVYvfc9OxGDdry
f0seJ8Vfn/OI5InGt0mvvh1xL5t+bkhYftBVadj/Bw31MbM2cJ/v0qi7hzXe6uWifIvHCDQFCC42
xF0FpedkLOUfldVfoOWWOqckLBdtT1facvRxfC4oIY+SWdrGHQUfKgUYuDX9DVGRxhOgZJdxCyWJ
6HtoCmVqPNqGH/wld0XnBvQgjynd/8jCPIjI0JtsldhOjp9n3Z5jxkaWASJmZM9VjoVxznY040on
whVXj8xjw3i4UKbGDhM6EK9+dueqG1jxT/IiwJpkDOGE1pkfI6m255y3SBpMn2JrrQLaHah4nt82
/Yqx7TAUUMxbEg2DLKbwM+CdibwGsiGZ/+7dwVEmNyBXSsBnwGrIC/qtSHO8GwO/oBYGA3ilUCN5
OoW4vFeYmdrc2NMx5gksHmdS7jaXQLXTBFmTCsNcBbazXR1h3jSw+sXljgbWVT3seliuAcPHEheP
xBVH+jqEWRg/6btgtAk8hbX1e4WVGVav8lJAARoZITCmQzLIegMurGtDG/P3TrUfCqQpI3jfRWVe
kRpDM9f8TlxhD0tyKGbotk2wND3rds/bvhfcF1VhDOQUgnsayaA7EdtOJcil8WpbWDWglxBHlKt0
35sEWbQYfkrJ/ncbRbQWcPauer2mbxW63pwqeZiuW+IGWFHpZhA8XQm5ibs7ulOfLQxYCIhZ7JKU
OJEdlOZkE9eMeJ+TKJYBvAd/0wRNlV6gFLb3R3iqP8aoz0dZVcEh8HvRXlKy4dqh4UWlxPvKQbXO
JsRyuYMIvLxQfjTXqPjnTxLHOy7sTD5W78etKqQ7Ac2xMt6X3CrmdDjXq+b31AD9oV/fiI4mJlZe
1LOM2z6NGpaz/jb7sG9ZEM7voT72A5Z7jwQY4UTfEjNbzfriEg0Q8fab5y7TC0Im30KZpAYKrisx
Boel1jQmkHb+55IysuDC8duBsb0P1DZ41WR2FbWn0eDkmbxsI2TeBkGf/10zuzBTGGfsEqV2sqyi
i33/xYbLD7aCS3hVZxHjqex6T78E9nZSXurcU1poixvZ/HP3g6gcXAnISXsOhA/B0aSlw3/QDHDH
GrrMH1UsZ2cKJP3Uh6rchLomAU6VPsbggA9kJKlzk8hibN1r38lcaaLlum/LOa8sgmSAlifUUOcd
jusW7WQwdFulS12qvhstGS/R+u+JEjRCU1XgSlJkTmaVfj0TVPjq7ntJEU2OkycCuhNjhOv9HTPd
JKB/auzMdop8d7MOfKtR6KVUaanSIkFwku4HnjUxj6/Cuas0hdkfvOdsapwrQj3DEC+2GzZLKIFy
JVcmkVkTBgJcQXR0fRgZzpiIy3Zfnb8xdo0q1/5eY30eQVVWyg2O8Q3C5YslNCHJDomkZRqbsJyy
8kHgzHagcncvGLSThvb/YFx107P/F3ht9SDOaWCl9Xuxa8/mqiPfODDd6ufP8/CrjsNCmpr0jw47
raPeDf5bPonN7QB4ay0+eefQoq2jj03q2MLJvp0DvY9sQa+ANMvTYVxTe/0nTXUC9GIqPmoPKA8r
atNta3+txyefgh+I/xRHlG/pA6o5d2bP6yv/pfUfyV/cC/kU2FtWFXJtxNCFbkwLO91D/5gDuafI
juG/3oG42P5yAj8kJ0kDRzxQgzryAGEBm8Cuo1v7ebgNcY0EzsjkXAwMwU1BXDR3CgJdV7ETnyTz
yJ96a2LWtni5VuLg2ldGdzWM70ZkDHGTK0fG69kjSRtkP72wwkGLVo7qBKT8WSq5z7gRh7pgS5/3
Xl/unxUF7xjnJjIpk9JDh0dbJJrHGIjaETdDgMcBC+3GaMmRbWI4vAZ+oJUI6wkvAsvHLVGRuCwI
nHlOmn1taK+TmEo9n2IivvkByBN5lVG4BoaGfPnXkgc+FP7KFnMuXk8SU2NB7/dB4FkRpmnqIgVQ
86TI+lgG3rzWx1JsGoAe+KXELz8GUpzngtTTl1wL7tWQOMBOR1X1MRA0x0E4qCZoThzgV7dULcu7
ct0NDvaIzfjMsdJi4FHtLuVro1Qf8F6haoAJghyBOwJxdHWJTWeYfbN4sYhqnHza+eO/OFp4qljo
I1+u5ubrZHU9x2u+4k+tt5tIbZjcctL8x6WNhSoh3xhevMNCoYNa56AyM1XOm7auSitBYzjZYajf
JOWEcgwzJ6vz01uz8pkj6zFpWyy95jNNq4eZgo1u7rrWzLPk3UfrSCl/A3rcDNzGT9oAQUGfkQ6x
tVmp0Q4p+A+abzDyhpqoZN83DZ70Lvo+GVK7ERk4dCLY+kNqCMhdlC6rbPpvJh+HbzGotiuLjd/y
3hbzdaQvQNhBMSRMvBfKbZ0Rw4YYjUP23vp8I5dJFFt+CQYnjC7DNv3eJCX14w1ruY9dzbf5bLRP
e6bE7nzum2f78x2EAogece2yvjQQJgmLt3FvCThWEO1i4H/PqIFLiNGhWyUxMskDxs6OJwCBS6QL
eMUePPCzzaQ5n6J8Fgrz7O3nx2927zmmgIm+Wj7vyJK0F01nQfVO/p1QO4wxQHrve/3QXMaRuq4E
FRtxj3fUeejpzDz/2epA/Hvo9QqqB/2sRF15piPMRian4/EE+HT/g0yYDdE8n0UkSYr/BvFXpCS/
0bIPEFvH3k6+ppfKEhEe5JAi3nwiUxAI5Zyz1Y5UgJJOlEGLyOsXotx7a+DFUEg6aFiBc/oICKqX
9BFdq1IAxiTLEe/pmXGF+3CnrQbzYAY1JVEaAscrNmstt7QEWGhQZbwOnythaf8vA1/BlQ812Sf0
XyrPnp6Uwy09c2WD94CsfN2lmHT5U3PIE323DcHh6ZhcOZ6Vdn7UmZcnFe3GOZlM1aAMKPJpBrxS
Rv0VRwqY+BJlEG6r7csFQ9EYyqbE4ZQOOtIft6KJzO23jPNFac9Blenqg6g+UCpvNa7SM5y7Q00s
s4C2WbvdJqVA6eN2F6wPNggz2VxQM/ZsS/VKqxtv1rN3F+nABtc7a9XDAJa1OVIaC1z9cQCLgHaR
Bgrc+W6CeTOgzbFcf7hL5JEGZpU7YC+6u7ywNvFUwt9mqBc1Ppa9xPn3LL2ys7M137EWHhfUfvLA
/xhShFpIin/I1jX0CpaIF9/oOAd4qRWfTLgzhnYbZU6tgnWy/naq4SDy+kWCVlE+329/0283Qwfl
OjFCulFH/hLItH81YC2Ylc6L+VuYqY3VFa1FnDC0aGpSNZTPY/OI8xR0F+T5JlBsGu2Oe/2o8xjS
VJIyPfw8Dj4BTq7p6ZcIgV6mbu56plL7XHmhXv1yA+96x3kY8mkXU9Z9sYrDeadTlxtryEq8Fu/k
6wp05dakQd3hT+7JcWiYnxK5mf9N8HWaP0bile0UIMHNljlmP1mpsZVCg0f4OLqYCJRBjWb05Enr
mf8Pbw5C9zbJGCRcMbitksnbUcmZEayaxpetEs60vDLz7PIvy5pM8oTB2rhvQBHpH8HAOBDIjzcQ
JsAOeDnpXIX5+W5AgnGusN++jNDT8qaljMmPiUX0hLPC7+8CaO2FRLK1eluHk2DoYbappS3kuAFU
dhmeCQG0xOFJxgxf2kaSYrV1Tb4DyNjcPtlQtLNRmGSO0pxg+ZasmGzL/IDDgDuIKW/oBN3ELdDp
fftlAwGFbbmvFUdLrGS4oEqWPNnbBS8BtuCcaUlogK6koaQaKjDz9QcpDC3Dv1DBXdXZDsSs4EVJ
Uibc78Cx0AL9ULeE/zfOgEcYqbSAuneOA3B6cbGqcpqs8/bE8WMu0O05nJ+XgkaXeB+RaJqpA+V0
cQL1RLn5q5mSJ0wereUWVFnOrR+9VUwIpSf72OhFZSQZUK/moubvvmBiQPI38BA1dIZEpslfZHpZ
ZNIehF8PlvQDlOuHPt8Arpl2PBhj8a/KVzaZEU95J8Jg89dgW5yksymDwAA2MvC2RVs6ra3wRjSv
dbO+GS2K0PgK7vrbcVNegb5N3/8XSj3sq4k78yUNfE1rMTdddjwXvZcROUR2QQg1lWQl28prAvvF
c0OfYRaw7/MGlpwluJ82MFvFimijgN0LYfpujhVvhcyVgDnWxcIpIOclrcDiTy1slE43InHti3us
GDetN10HhY10/zSBjG3Q16qLk/Rs8jYGqORqEGym9Q6qczYK5kqt5jMpLisQdnNJCfrpVhnD12Bx
im/BNLoFrPTxIKkhB2Uu+NHhQ+0j23oSSVIUausMX6ozfuBR8O0e7m/ZUEDtaUpZ0Y4OYoaD75xi
PJwlK8rXf0MZuT3Hqu6LWfDVh5WHz8XePWSPLlLYFuIMGwDFQcwYVi5QalnHT+h/0FOT4MBbHbWZ
TkRep31DblVV3QkgEdxZoQJZMG9hq14QvgK/j/7tRC1rlLC8+qdRTylWr0vBePB8ZEtd2XmLxVIT
Xi8J6afu6gsn8sn0qt9RWuOp0qGxTBdIncxEBedYyPNeK6ZJWi03FYKXkMIpRXA9i3XpLbpWLkL3
KnDTdaeFT6wkJ/HSEBaVnsCKLt51yWv0S7F7ipu+A8vN0YCNKY8XNLtS/Swgved+1qDZK8BpCSdN
m0SOF0Bp+STotwepey+ZcKZjHJ6E2t5eYsIzoTj2iD0ufiM2z/6dd/g5mwQjks3CcweNqe7kEsIE
iYHs6VYSlSlvggwnCGNYhjCEseFjAVNlxiIOA7DMwOJEnJARQNLWm66D4EganHvOzUEwWjh3Ekqp
CQkIYajlYj9ZaQqPgn4uu3Y+7ZyV3/VGtRyHubiMvTHTd4j2qR31gwVJ2BzEk8xAlxC2a4ehNA+2
zTVR/Dg6zlzdMIeKnsaIfJS6JZe+B5xNKY7b/w7rn/ytfiYKVX4BakZAf7hNfrq7ShveHkarr5WF
cuxOuEJAZ0x/LClQW3Gv4chEB2RYLZ+EBZWMfeq2Iafn5BhV2rVduxdL9Gn3pGG2B1+medcIw7bg
i5HRQS09StOAb5PX8Q9xeDdoLtH4+UGlRJrRt7IcN6Lq1hZ41XP06tLa8GX80dToHWQYIocswvYU
nhRI6NsJTaS+DgBNZqP09y1+QKsy5fEVKY6XF5GeADHnsrwyQNeGSnBsvgRJg7AqKMibE09Qh7K6
gmXSbnrUi0L4DBBine/OvGsNXqyjGQL3/yGuY36UE9jTT+nM2dCoQijR+g970wRkA2wwu9mCwrsS
1mLOCx7ZITXnaaGX0M/nmiewC3NxBBlgoE5EnehEWmvcswGswknMlk6HkdJjp7AwC//DM3w+xJZS
4Ad5buqnbdiZy1kaTMjdNVNCP7OllfyZWrBZlVr8zFDP1GG+W+jmOOIwPiCnRSrKWfs3l0ugyUhJ
h7JIZHEp4O3wFpV/gPVWxxviJP3gZsY/2HF/AwqWCJ49Il8Otem3CnwSOOo5LuEpL8T/n6RTFHFF
ozkxRFa0zgAUYNxlqGgM9Q1Ek602ufI6ZYzk9BjU8b5/Bx0RHCMYKTmKzsSHQKjmKoQb5ZKahMBK
MkkVXKFvqwIPVHt/7u4ZvaaplWtH1c92PV6SVL2Cb4Zz751IuURZ7ZkWN5KtJIumvwWEAdLblh93
XaHSlfWgzTDdi2G0EnRJ5MSgBVLzJrxTb+TaOdPtZq/tG78MLDKZQyuVJLvxfZSiBuzjUF8JY9h0
1kDZLOKL0oDjEbXbBLtc6ObbNYvmKacyc88L1UPSjDtXrmfvSfa0s0CFO98TKKkWOfDSmLSXqRnm
Jr3DxBhPA4XDrwkvqbakJBsSFUn9FmfqPQUFOP4LnGKGjUyPQWQfNsKwN/BAM/JdKXkoRu57mBtV
ACz8/wTbyVFEjjy8LY9PMVKllT4ByY3lYJHFKlEF8Lkb0Y43uynHk7uM1N+IjnZ/mJzKyCc6r8If
3o66i9LtDq5cBIk4+0Y8KlC/0eEM6mRmNvLl94iwbv1rZDqYs34LDE1TYTHs0C6m4OSzWJ16669P
AUzrRyqKnNlAXNOt+QISPFvay92stt8noKVQYnAEeHaBy1JX92RyxHDEMiGlAZiPfE+ODboB122T
vVKY9vJ1exwSZtbUlqONDDQYndGaBtnURDtqkeHD7ipgnFgAm8Q4Y7SfaL9cI0sNS5m3yw7G9D5Q
uhSq6Em4bd0K9Mw08LypQERBgwThuJhxEAkki9MZh/pTZhWnA6WAlQI7F3KF1U/qL3f7n4evnNfZ
LcaaqEuCOGmSvL/xxnyddCLhPMWguPAhmVWJvHXh/QJq2OtxCQvu1p0HWSZz2hhVcu+7TIuip962
y/JA078HqSdGnKEbraP7L/NqAPcJFVukg7pBnEz/ISUZ9pS7/gEWWPcFwleWirB5KE1gmXGePGoK
X3uCyKYUX3ftm3VpLwwontlgzwt+lOMlTlhIu26y3n2L6uHLOKgWKSMMl0q7v0p1/lpyKnV+Pnns
SJye24lfmikLwNS3AJfWENZWScf5RyXB7VcfRAeelRXzjyo0F3Srfv/BgCwCCMwB0Ref0AcNTi7S
PQCNrgaTVXoWMBYWjPIb7vZg01MglIKnhMZFdUUHQE32TH+Vf5yf51ZWFJcySqsTFpsR4kTs8zyO
m959ch1olB07yh87IaV18YL/OHZkhRxiTZEh+FSo5Pd9HYQx8PXm7ZcVX7uRaudtiJrwZgBMD5Y1
ekK38u1s1v7wwy1J0moso87K4FflK5GK/INTCqUPNFJgtNED8SRFPb8oEjhmuZmxleHLmXgFCOe/
Onjaow4LvdRwkQR8fmVwBGH+t4yZloZgb0vJZXIS8nyvKJbxVU+hA6gJde5qHK8U1QhJyetvPXQU
u4H/Mn8nRosY8bHO3oSTNO7L7n74lLPycuA+sTeRzjj+YXdlDWR6fjoitV/MO+WYDQ4lv1ugCr9h
gZ+0dUGTZiKptZaT81W8BHF1OcrfgoBs04Xisxell52TmzRJnhcY0A8OnjTv+pPTyDGdorF1MssI
s49oJ+bnprJ0YPAqTAAJP7b6zOuUe2yZukAO38he0e8eKWTKzuGKoW+Cxvrtx8ST0bpahO/r0f4Q
U564La03+hJxl3JHDpnT4TgF1MMDZwmDjd3eBx46DHHqc7KMBrgvxDsDRn1VHDfK4hVRlZWQSLf2
TxLgOUti8KfzBQGx9UJLoudonPpjRvRTIeh+r2vS70dAQ6poyqkdvFSgJbV/tBa8PMrOiAIh2eUZ
5SUw4QUfWHyzBzt92k5ay9IYQnNMHTKHMk+QSpNcHw1nMC5WfytYLAwdCe45MppiTvEgIY4ECAOH
NyY/yw0kNWePOeKNgVuSXA9O1VmkAWU5XAp+Uk1QaKSjALzPlVbPnwDZ1R6cYmQouL+/qUwuNssl
UVsaRazyp2/m+6SymGmh+9cHf84k/Z1wlVAE4sHzQlcPm+1FUVom5ojjYGar2c+OtY7LAykWrari
6hbgeT/j55c57TDjUAMtAOh5PvUFJ/hF5tChNA9auXNbqBDfsN+txnrrfUeip6NCpHV8s+RihaL3
HGTXA6PkmnZO215IdCVVICAVGk77Hh5FPNmm86SjwJqc8iDQtChbygxZ99gZxzohZF0djY2U3Jor
4dSJT91WvMWtI9f9zjiaZ26f+MCCaMNusN7uOkIXiZ6nC2nNjxuTeMNoNYA1XOH4i5hHiqfA9ELI
BRQQ8gB5k51eUROPTuJoaBKj00DmD8KrWWu8jijmnYrU/+kFnt/7bGbap55+6G6Dp/PSFh2QfB9C
P6xF3IY8P7kML1hD9TmuavkXmRnbp9YiDYu4rTt8NdouMRkUZSBYvu+VRrAc6POWatIgJApUlIhf
V4diFs7SnZ1jgwZaLPUheIZYItrYyXUq7U+QosZn+cAiI9Vo16Ma+p3iEe6OiTaOvu6G2+YLrb0C
DQtr2pf7pqZ7PaC+ILOUYXDC9j0DAWdPqciEbJtBTgdfBesoqH2ppcczyj+EnoGzYaSXFECdd9gC
/CH0RNc8FT17d/wdKlxQPhMWPKx48qHmoqHzQ7zL0BrE9mHWVOc0mMJBb6Xq+tI2qcTYpEbhTdwH
fCmM0sd1jcWncMWbvnySUvnoDgNDWGbgGXXFpFbiJitoesjBQxZEtqX6moTj4D3pGI2+HHkT9WAJ
bQBu0Dmche7Udcp+0Xp5enbJ1tgXaW8wO4j9fukrT2OIEWHs02Sud2tGwS+c+fbEXOGtCvKrC573
iJK6Nbh9p+4i11yBIR0lk4FTNaRU0EyGXN51ONEv/sd1AnbCvBHQLOWYyfG69UWJRkdd4Cez9t5U
ynHOY1iqpowt5jhu+J+0iMObDsq8YZ4A8wPD06egsty8FhN0hJW9cEnKF47BsiRzzEWMgzFGLg4l
XdvUujOWn8m5ykJ8oXrvut5WTBnxDaog7puot+Xe6YwZvQcozdvvqCR/fh5MeZfUghgBoQSmIQ2i
0fvW7UNvssw2NdJZRGVPhBvekqMt58C00OOufUxVtGMFnGy+f1x9jCWO4Y81vhzuzfsMrGZG/82v
8Vdbsiogy/q5BxdJp+Ot9IJnEbQTuCa+OKGGZKHuk0TbhqSST40naIs41sJVCfOjCyvjpWnga9jA
G2l+bRrPc+1tHDD12r1IV/4zT9lMSSjR0U357+XAxehmi2gbCBdNtCBoTg/LIEyln1IlrMtgd4nq
Of5ZVPTJBocUE1OGvy2ciKV/Gcwd/gEXedk94YNdwOtT2L3khIJsyGhCZgszRTF0rLSgL1cXov6/
gWJnFKQK/bBDHa2P16t+kUlaahPN0sins6xb36EKF8ENIk+3NKVWCVgxgRQGMkOdboyx/wFmCHod
YfDH1bKnPgl8KTSyEstOwX7+LbVYYdkPO8m30lV1RX2T+rDG/HQcjwu3nQ39x5hm9WWbY1Qjr0UY
ykd+4ImwwRoDSEZglTNg+9ncEEAJVXHj3rVstcvfcTnAJN/0DNsB3DvTXIhLOzHu1fuLpkY9wSB1
sS0zSfHTes739daM/XPdpWaVHpQnClLgroVAWmZ/zPB2psdFB8mH7qrL/m66Prif97OmfpBGKMeg
Xl7lg0nkHC84KEPQAVaeL/1fqUI8EncJO7Up2cv2rDMYiUjWjEECaQJMpiR5VMANnblS2xFpI1SG
yWOUI+DuSGwrdSoSqdx9RT70G0bdzseWGcJG2ZIdgRR7qW5cNNMnDkmZZnijpb63bL6RJxfMSxOg
1DqYUnhfoOQ+cHI3L5b9DbkxR4Ap+1E2VROBoX5GId4D/GKLjcITJhCpxAupeGrAY6PtEv05SfzO
zNnJjm6dvFDtbgQKtOa75QsbQw3jon9fgNdBXGEK+YHR4As+WSIn2+N+gHKXHMCv+dyOjSQPpaao
IZIG4V5G7ApyDQJLF8v8vbBhwstaz1ykoY/vHfytCdmxKkuXSKdJB+//bnzq6kEXsZaJ7JDuXSe5
+boEGnExLVDSIo2UH9RjmEwRS+82QYV4ZIvMesIa1pHp7zg/CHvQ2fWiJDRVSSiLna5zOgFxs5hA
ICz95REixOgZSti+TAyKDOcObaAE2ukBAb3fWw0qYDC7ydOVW3x92cPfStD+TBxoqXYdE6sEipDp
US/shbTN5ALpfyQIjVx8El182nceTNh4IC1HUu9WcGaGRzzNKRnDZNpu6f1WU4zzIC8X1CZDBRdb
OsSMdnErkXJtFbzUCCKgzB1lHxoWV/HtseNhrMZU0mSVfuXmPocc1dXlbTBFWoR06ECTjKtPf4Xv
HbWysqMsAeKkryifjZ+i9nsfueecrtkGBokRShhyvsfui5W/8K8a95A/cv548MvpjTuz4QOCzzs+
mxWcCDLIXucf1YniOtB5dSMYFZXiBRGZk5XViTnYkkuRXHf6TdOk3KkUJkT2uUOFeX9ETiw0+twF
zL+30RhvdkerSfPo3U4VLivvCeJeCEV28NX9O/31+o0ztDv39Cl/QgE9wTZfAAIFg8205JHNGq0S
n3iAVAydd9O9p3sDEHcM6xiETxhjnmvs9/R2uxyzqtwgy9nu2RwP/KdWagFCLk5ZCsNNPFv6EmsI
967Js5V1ALJOMxTOqt7l0LrA0IVJva9bAtpc7tMyrwqHGk5s8dj4keLji9md8Ua+9s78gr2+zUfu
4+H2MhFIPF3ZEHHXMzcLeNKMuL7efgetIOgwy6kpNRlQkwSFtEJ6LYxyNRHPOXKxWJ//xgrylGXi
GWjv1zdYHj4a/OIaV4F4zJX4sxPigDGb/xlRcKVbvzmxN3lDmSNo9tTg8A2peSc0ojiiiuTDED8g
ZkPGruElvDvM0k8UtEadPHG9Ygley0jvvS2tTvE1OdyUiBlZfHRXtGV2QzZ8IAByg0MISz9rVp2L
IrYi8VKJjmcyrP6d3WPY/FrNzdNwcwACjBnDixZs6HZSg2iuy91UotYT3xB6R59+8HdscdT9CF+0
zq4CgBToqPHL5t9ZEJ6RFe7oChaud/1fVBpd8Ul5VGt6EnhI7nYjSuuAH8SV8+Ir6evwCtCiM/BY
zqwlVQTdlKIK4Ham3gZJeDiiY7AZTMkSLO3k9SVrKUtEZGUHVVlqOw4LmzTFqFQBrPciNaedJSWj
BnAoS8HMMyTlNyischCDDcq1PGL8Umx/niwxNpKAN/SBE8L8jPTp2eUXa1+y5jZvyqiGdnfxHfXE
56sg25AMI8Y1vzeXCaOyxqGRWQVrGSD8BRSnNFkYWFtQTEJf46e6YjVsyPDVWPlm4C20h4YfbslY
nVqDaLzmOOxNYQcubbkHIwbulgSqtrEuORHarG+AzlxHpJvb0aeoeN25943mpIdl1fgUvzoMokfI
z22Aj10ngh87q61hI4V1UuNeXs2NAWv+r4nCRlZbfwDL0ZUaPNbrYidMY0b6oB70HYEDWbBiEwpY
PIzW7T7DJLrp4HgGbGxy1Fw3+JGh1wy8+PgdnkuqR8Z0VBk9Q/7H1XwygD+gYYfwT1qPxHAQX5Lt
R7SyKwTGZvxRyZ4sqto5XDDKL7kzEzzRaN8ZJxDNoiGhlwmvO4kIRFYrJx+KWFyEc2/F62fNgcpN
LuyIshcr80eKzw4Hmxu5IOUowH0NuRDGnabHtwNoV8yTbV+PnSTXE2kmFQnvSxqRGyyk+4fdmEHe
7kFglnTTYcJFBfI06XFO3IxNbrkwglbd3hQVyhaU55bvVGBiC21rr++RalUZQ/mz2HIMonDpKQMc
kAQU1kUDphJBWSVYVSSyX8mo6ib18RpcyL21CKAU5pw2W5gC0VkouPFTwyzK2yPrgr/nRVNMDAoq
lP7/3r/x23r2mbT7Jpo7RK1C5LSM/PlAtnsjTr/A9BBiODTUcQKAIJjubxGyGLR0kplhcY7svrJP
mF6YLvI4jG5RFKxW5glFfaA6v3JOsoe5O8hiL4aR6BSns35ix3qH5qeny9xUyU+TNpN506rK2RNO
fE/MwK4OrlKWjTYyl5HAfkrYiHrCONldJ15VaweqsLth/5BHYtLPlhjuXmjeWP17e6237OlpBnRt
SGqyrmxJh19PKls++1wGSAfxc1+ebM+8e1kPqweYO8eA6WlXt1nvtbRAlrqTB59emBwDxua8XrWX
4F5GBshAdFM77KoWKpYbPNyux3BA+EPehWMBoIxxxDA7RhBkxOiP3YWUjLi5FvJxnl2/8cyLsft5
7rtAA9aYRa731P7OEGxbZ36PTRyXXTQd1enkULbCBRzr12gMfdCJ0AhcG6ZwRMutnzez/u4Tn0aq
dZ2VURMzElqkeGgX6bFJSj7FM5QI4Kd9shGTae0/Vxu+NqVmjTfkBYEnIR6gyJcFjIfRgrvToeJr
B2vAzMZcO3hZXMn2aVIpB1mO2tLbNLzL5H1mXOTUzP+HQX0XIzs4w2f4isXCFjnzuJPFG3Py51KD
M93jFMhm5NjZcJ0vZD63YOYbjQV4IAp7bf28zbIepuQ3+lebcX0WinpDpZ2dbuxAjWtavt+IbjMq
H81VFfGhwXVhu5UqC1Mg4bL3KiDQ/HGaPkydsqA/35g4zsCDIfUOOO6291ia1r0LvGHnf2pTvvkR
j1hvZUNbZxeSvM+YtXcrLIAx0xdNlCE1Wwi0HPV2JNOPnmrkg+gXxG6rXpYvbX1hd+cjo4qnL13e
IsyR9L+Nn6u4rkxkNXnpIqO0R7YPfyYghK1ZO3klujkK4Yb852ok69sgetDmQzM1JV6afmo+/mLn
82AVhgkmnbsAaZJ4IF4XQNIy16h/nJU49EE3+QqCL7Zap8Pc+hAc2E4mWfSU0360X4enF3F/ml1T
q/rPXtdm8MHOL1BImktj8pODQLgadG8UQ2Pj4dI1T6KHMIf6TLLAwtvVO9TLMZE4UmgQb0K/EajQ
6ruZDSbr0Gng3gg+cDzo192jluwkWxUSFb4UDkL6HvzoZOsWfsw1SYeF+5I+6Y4GBghKaZ9UxUrM
mwkAgnc8uKlqF4Vg7QnjgyIkyMUAJtw3b9M3Y2Aiz+uPLZ1Wj2fizmrrK9HPw0SODRLWVSYORZba
r7fNSYEZMn6fzm17fsiWuxIt2arJxqkzwl+JYpPLckkQ12H5P5GTLqQ3iVSryDfB5DyNbUr/wLvV
LrsuQqD4PUyN+nTA3gcb6YiSZXAMdWyv12MsZRvejU7MsbL/VanVgHSLdjwxXtRq03ANi+qSA33N
yc67wlwAiIwtjjahf5na7/qb6qd1x7e+Z0l28vMjvZq1PDhgn0p2Qd/ifcotNTG6TAsYmF4nMC5k
ZWdClVNt1qiutWW/5NhVVEUPF16s9BqxK2xMbK3fpz11+F1V2ctarVyqvWSB8XSe0C+5UNGMLuTM
BXJKTwr384Dl4/FD1qeuxlvL97FuVPKpjc6QyVR9rKBtBvEZEsq991aYQQQw+0qM0pRfjkAdoXQu
Gv2suX97deVMqZ2Snv179B6FA/WPrjNy0oziWDX3Tb8ABGfiIjEOHTcb7mLWLNK9DrpEtD84Q7DI
a1R9BDrwiVGQtzMQ7js2Ox/AdTnj/FWWuW+3DfFsdD+f2qDSn+F0L2i/ysrsQdnMSU+/H4/xhBr9
3pjK4dVRUFC/oOVG0kwAaHWF8X1D3YoU7ht+M82i2AgmbxNQlB4idMc/g2SE3On4PRd9eMbogbN4
pJGIJRVKfWaZ3fvL1peTifHqFX1o/DlA1sJN5/OvQQVmk3oPbUE/4vwcO3C3iG6VlJV3hw7U4qfg
hz1KMXcwpZwQP9npnjPMnnoSIq8rU5oIopUyaU7F/K/655XCgzd5S8vgcdvma4ieH/e1S8/7l91G
a8AXhQv0klDZElFFxK+jlgWjUxoux4ku6SCKFEaPS3aEvVj5Pf70mTaPq3/cQgFTJxEQxgWksoW2
Drtz/xLFSrcSWTOBJrOP4C71ShKlQLX/hrBE8u7Jh+s2f3seE7DDJ/0ORe+KhWGqHRmvknMtghAN
TRQgH1PIeBux3uH2Xx3dMQpp4HIDxeUc4J4GT8GCWIaMUSGDHDHOD2U1TALOanSlJOVjaeKoK1mn
a7oKcTiCzN2OP6bpoXtYaFpdZJGgr8Y2muLXiPrlG7pG5oNzfyviVwBK4q9JWglK1+RIXaDUzuKy
y21vjV0mjQ/g/eOWANNqQ0PyWHzXVG7HnY5h+l5jt6tSB5g4wX1e+9jXvC99AWGqRtbOQMkLbSPz
yS22G8OK5Fa6gfjM1JG+nUBY9cNcOFhMjclMUSTv9NPbbfgAMPg629XCp1T4B9gc3N+4OXYSf6HX
t5f+I3gM5XQgSPRHk9/nVI4dI3C5WkZFaR2ZB+KpOu6MBMEv9loGOu5cU33AB7z1aTtRod+78ZoC
KZTBCB77iBAhS8t0vROioGwq9Mh5NLLvqw9lT8DBRqR7UyXzB6YaUMRYaHE4a2d1neLgDyWpCKJn
xYIFU77plsbmBdJk9GLGqdXgXxouLvoycgJnwmnEmon5RmGr6pn6e8aEr4Gp3anRdJJ84b1lC8OS
7i3Jo4+qRPEcjPy3N32LxR0ZYBIzIozc2caxyLK20sUTHXsZmvVU2/7euITe1978S4+I7ziNQWbk
7cOcbyWKUMeClC1kmBbZwtJ2iHkJMviSGjT4+ibAW2rHRChjqH8KkVV3J2+1lyjIClnUpSmzHMVh
sxGcB/3BD8gWlxT21qZr3wuaQI8D+laP2aJFmY0ESYDo7WIX7vU0eZJWkylRrFso7VOdzf1QBiPX
JXA0vFANwJjrOsbbkUUuBs6OqAN3v1Mh5HBUh1WTMRq71u5CPLPsJh9k2bmnIQ9x3hKcDZWT33bZ
jS08Ms+w/H7CLqEUfzmyE+1t4LEUXOUUfpsZn3+2d/l/etIH6aMgY1gKajN2jsV8x4knkLWxkrXb
rIT5ujqtwKHitDSpjJjvO9HC0dtW5f7NGznx188C3jSbF4IlJDhNGh/Gxe7KAHFG+AbP0jIfG8Mo
BRiNjLIasNVwgc+NSbVHQ9TEKNYwe8dfW53a8xD7Ebypwn/hx7nTkUibttbT7PrOPBLt28+/8Sqo
UDgwjE+qpry9MXlxI24ASww8xlcUicDpFONlqAfFoCHrNxLLGTN6KAM0VH750WN3Q4QwGsQPrwMU
ncDhEUBu+CVYdLZu0EtULrR//6pZdaQ57X7cVhfV5rmIt/o+MYlrpxkD7XGaKbltESwQ9Q+tW7Yf
dNZC5WdXxrKVTdeHEjQznBfBwXJJXYdLpgy4LFqFs06lEgdUMsjPaLyg0FPfFwPkT+V/axBSuAKq
Y1BgHCruyY1aEX30S+542uFxQgc0NZ6DeTmhw1xJHzKhCl9Jfvo4l9XjskGcv75utPH/7tHH4LL4
E3SZKbAN/41eJOtLtKzNimmctXMsNd0p0QXTzNnJhC81bQ3QmCFG9FntTzesC0XDTylB7GL+SzdC
PehhwhV8Be2RtOICbu6W8F2kF3l5qIGmx2zmmsWQN+5JakKDnRnJPreR4ftNWC+/sVjm+73ePR+6
tL5Wct8VPUuhSGQgXKzA3G46gERKROBNf0AiRmqUfhKQ5oddL5DDS9x76R0ZEMTcy0dBnshaauFF
qDXHK4ke/+1Hm7BTmxvv3saFfDb3ekA3P5w1PIhLxGjub1xzFKAkowZwY6wCPBddifxYjc+K1SGA
lJ/ngzzWHu8Xr9fkgdYTJJkdcIFY3St80aQHFVETDUuNwwFmMEnZtCTEilBj2Wbr5oOpe+ldBh3+
Wl8QkQRalIDLCO0WltVvF8f2XyUDtoSIKcMcAtmvrpsE4ohgOKevscrWvbk/KztTxa9Ym9mU2d95
jYRqqlVy8qgKcEQGY76JpHoAfLjtec71dZNw7gD08kzf9+23AEgWe900ehH/r89p+zJyalxwE1A9
wDd9eeSJOpYX+/APdDyFapWvFiIb9m8AzwBRm0hwqxCzmDPYlfGHC6w/zD2UrC/zXiaWgDwOOeH5
aRWGQ5uUHxbsOH/PsUc6CJWBFrQ1iByHHdUmnTzNd0pPm+R5AMsoRtV7k1FMT/ZOKu00S0vi1auk
jQz3qLKOUIrsf0B9I+fPWYLFnY00o54zgjfr+pkhKlYR6PSj0MmKaCDCgo2izDIC2qsKZQa/Vixy
53RI5mHJdhUyVYrUdzEQ3+UkAuS8XbIGRtJfts0Kb3HQTHM+yjdX78EZ4OcClX1SzKy5Ci5FXj8U
TMEFGL8ouKipQqy6JOqAxyMMqdepPWUxOhmxw/fk6po/KuF0Ek/pA398qiSPgFwiX1MxHtIJ53Li
a3vgkYovhadzvU5ah7vQG0QnzOsDE+zSsfVwpyC1gxpMuiUr9ir/s2N8f0Vx0eTCZYwsCYGiOmqv
ykWMoFtIFwDbwOO3ARnX8ZKUoAEOmOCSJ/vbCSqGx8g4dF5suCG0z1Lt0T4s8tnBEn8+mOrhhGqf
9I5XaVjKE8DQ4oBrJhDdXq4h5ZlEhIoSLoOT8LmB7B1ouEXY5+G0ykh6V5LmA7km+rmWXLYAr3MA
NOR720qL7PTtectoimoTmd32Ql1Nvzr2tGeKoTfwrzd6S3gsxz96gzfuD3qDpbmxeNEqx34m+T/z
UAahpAMHeoXVf1W3VFkwyC/bVk8/EXoZTEd9R4ZahbE8qpc2Wklmnnjr8PitCCNrUyCP25NTgeEu
HUeGVWa6yl+csJupW6gFpbFDHcm32otizPPbUVyMVRBL0Oi9y2b78R01ma7tFrm3UtqF9nSoDbuu
oMnuVaQqMeDiaAfbI7z6ity3S9JkgTK6RY0hdKbIdOAEbbDGU3I0SEKvs7oaa26RFKwuq6WXHzWQ
4sqh72DPjaBCqTqaOMgPyYqJP0QHFH64a7SW3RxDrNsHJSYe6WsEqoal612K3/zpj3sqNWNhP0I8
Y4Safxg9i66VbbgZ4naTK/6neJwZkw9e4Gzvm8IqjdQlDhB3p2z+2ZjdQsXlraLGLvV9zJvYtBPu
mINt7Yy9R4SKYEc9LboAL2DGoDq5eZBCwrs/Tpi14z0h2XUvjFsdGc4qrt6xZzGeGrQHzC/Zb2RA
+4v+ZRzxD+n+yUYB2ofi4l1T2aacGpmfltHk36wmtx8FYxrWBfOtVPxWjlsFuMQ/oSkbMQ5pR6Bj
Z8WKdTps624+jLNbBwA2zGptxwH8LhM6LYTQOyBVMRylcdSX4Rz1UyyLPd+M3jZ7OZTqvoPLyWaU
TBHY47A5VmYWKDSWOhpTBAoFRzl149hr2hYYsU0wmgrIb73bLvfxGOlNxs25hokpQuKweLqiurG1
glq7MHBUn7Wg3EEkX99Ph+Y4JpoFZ0gd9aYWluD/WVdbtEXot9st3zIPVGEtctL03FiinRfc8kUg
1eoIhvvFjeW8K86KF0rlSh8z72PJvPVhBERkfT3kNlE1eTJCHtcRz8mXy+kZjbbiuj9IIG9K5+wB
EvwYp/PaK/Y522971K9dWW+2An2GX1kifWpLfOfM035/pVDLSeqKuF9moeqDg+LvIip0ET/PZquP
9b99eUifJRVNvIPMCef2QBMWkxz97z8cNBO8t7oAZd1ie7VnsLK/dYgdO5M+zo9KwEPf3Y7mZbVS
qzgsmIPu/iqJn/RpqyfMmtSOeWiEh0O2FuzPEbwv2oo93jEnKuiQbSoO+ZNcL7/fV+KdqWU2OTds
mNwt6HvjOZaxpY7yB/misCVxW8o3TLQW6wWW4IlDE0CL7ODZm3VE5JUAUigu9Vj98dOw/+Xi5NVO
qwcpTh83ZNqxcmkJWKOBlJQTw9R1LyXGXikBhZWQEuKkGLkyEiG4gzNu7AWcQwAbmc8cfNHIpytm
Ml0vPUNTuYDDON9tHUgu0zd76UYe+p97WOxSxuI1edAf4aY5Fnyes4LFm7Pum9pHOhmPRBhOpNUt
XN75wlCVoDAnm6NsPyT3tHJM+mMdVhJ6kF+OzgU/DJApTArSC4T0t6R3iQKCrT8fgL4imMRMxXcW
MoNSr7QgxyqiWEgm0DrFUKelFfMl1epyycTUh1Vp/kBgTsCPqKUQknj3LimufxF66+MrhpYbPt2q
uy34fGR/wdQHeevLnJWhLEhYXDb0SIXLYyc9xXOeLdyMCPhG3390ynovIxksDTb+kKnkkyXXsy8M
GEJKL73ZUFXbhjvIKXABi5djrclc6VY91MppgSIWGXYgx7FNx7/j/lOU6NbXxEZvAxP8758NsZnu
AcF0NHr9DoecFPNYnN9j9crfptYbCqfWKFPsmNwMfbLkr9MY2Dt+ljXP8XZAfjPqp43TUMnD6z91
oIMnmf15Ff/ZaqIZ2Wp6DB1xd4y3YqTcRO1LTmfX/kOb9uUHa5LvKG3/lhh+fGqfQgyQYi8Uc3HY
EbYUeKrr6596P1Zd9ky+cftIuf5fdlUgY21hg6Oos4ZvL+0XsEQAeMw6GVcTLvH60fhNDmrxGBCL
wdN7NPEqP+stxor2Qj4IrJiAHFZqdWLCDDY7j62jRyCScb3x6s8N7hk28CpxlENtipOa7w3+b1aJ
l7ZET5mZLuEFEq08dFYfvcRvl48vXcu5vVgZTqKOCz4Hxfo59/QyRbKrNIqUBrH+jotvXCAHaC5i
4sogTYD1ThRJKzucNVRGupwPmewxsp/Lpr4uIxc/nReR7PttmkVNcPosR9BPAIslodVfMcPOJy9k
gkwpwaEYMvdYePssQmx/9JeiAWSET86L9m2e6dDib6ADSJ2eWOon4pvpLOamC4KE8Rxe7HG7cwSG
crSodX3IpeAGz1gwnkmX8EGGpy7tRwBB4XRWgt0CJKaH15rCa6v5ghBd1g2zE5JuukzCaQTSflay
VStomUTMOn2UEWOxmZb51I5OnC+kYVlK5ogPEF0hI1g8xFH68hVoVkyGsAVDBnGgLOJPnJ+/ALwX
PK3yOnLS/6w0D+QygzYKGSHEsUYSXb/ScrJybH8eb6GaTFKM3OGeDhE94TBN2ZijXm7tE3e4Pqdo
PPn7oukkDwHZYF4ws70Z+/lWiS8wG/xfBd72HnM2W3+NgMKbk3AKo4apprU4ok8cBYem2fWh7nOZ
iv96g7ysylhP7PXkXG7QJhdpMjTF2Pi6ARFLKFj5mffEro2phYE4HbTgDXQ35799oHbMKBKgMgIC
KI6Vglgg0C9/ebmaNkXbVsia5tz/eqjDIw+YiAa4PZf6cFSwje4E8chtxRQWczYncV2quEArCIuU
WzmtxbX0jTGZj4RA2dgvOGy1G6is9rYzyU1MrVcXdLiphUwqDWS8nL8D7aE/W/0TCUOyJHI/E7q+
4uIZcJ6cYa5EdE3AtrNuqR4tfKBWU7bqLFAz/uwV87vh5hbJwehq9UaR0sZVWYiheVxEmE2zufbB
zSOIhfVK19bib539QisNNHoxhMXRC8VSfLO41t7XSP7qDtkhuFr3T95P1h/j2y21HcUBwWdgED/+
jLk7JjSLIg9oJoGoVXvU4pxhJIk2HKNE6Cn9Qn+cqExYfKIGq/IeA8BKfe8Dem3/x9SBXqYE3I5X
lWPUpSpjR6mOr7eE9l8CxW27mLJZwCpzjZpwavYVIhbeeV63pWZev9AwSxqJj7JE7t2ot943Utz3
5lHJq2ND/HFsV5oSwGh9RCalfIRibx75k5mICMqLGOZGn84lqehtvBX+KlBFIlrIwCw7VJAhagbG
TWDamIrd/d8QSDW7pbqv/HS9XVmBSZUNhAgsWZlPGTg6/pbRRgomDncmdALul+lpBTVEoBwFoQjw
FWu2D2Bmlcstnlne5myleuhTbkGwm7U7dxsJlf7+XS+7LjeAHjZp8fNlpiyfGRxrsNGz8cZRuCFF
XvlGB53N+ywNBbtDQRuyTmDREA5NhXN+R53Qi0PWIBWB/fdYp8Nu0H/Xy92K7elOiqh7yZPVmOT6
zIhfsCLAi5W/x3jjNRAyGzh6dyvwslHDqc3OIwcnvqU7FrWMkhYyzf6UpQXWSof6qfAkMooqOD3a
PwcpRyR2poRIouQetPh//GQGAChppS7w1nONDGxrJvq8BE6pO5lR/+UZCM4CeSszFm1KABkJXnfC
WqGQI0kOVatYR4hnqaYXsleYRAM8ebUtChny9tOEmcsABRIEvvZx0jUVSqskozIXofxyVPWrOaC+
lkhOV4yj/I1aG3S8qLeZPREMUI8zsO3VNoUBU3EKiA1Bk30LB6ddPhYXwebnw8/PYd7Bdxw/S1GG
4b0jwMdmGbX6J05EbWloTsaUlLMfiTiSHFu3BJPN4qb6AB+n2l7FkUZ2nozH4u85LAmuIIm8vLHh
MWX1PfkjlhU/nm8uxGkjzadcby8aRXDeGrA0xBSDGvJ62WuA5vvnJCV6/HjufuLZCO4C+MNlTV1x
lKjDcpUGmTDwHnw77igV3qzAZBorQPcpSkvEwVF0Cy2+APdWV7gbygQhrgQ1kR6fpAsN9nQTFWHP
zgpaDKacNbctckext3dIfAe5vdtfKzRfEqlRdSOJxkGcGEbFmAOwool3x0jGMSUWVHx+rSLaj3Wo
NeRuCPks65E7stBvjfC9ELco+kYYaZAuXCh3SXKbCbVDmXQqIqthwHOafH+YpJkxTySlZtMwNPDf
6hjoF4XGztrQlhs+8Oenn2qBpiq0GkZ+yKr2AZ+UotxpXqguwSQsuOZ7dQUyoBmsgrJHI/9BhqvZ
qYMQ/TjL3rJ+oGWdYItckGvQO0tIFB/8NsEPNw1mvzg1aLMXrj7k0RvVonYV8MYAjjqaB2v9nhyb
C09W6gfsHIiX++C0qNEvBawCSbcnR/9zf4/8e5USRUZiTeqFMJqigXzxZDpfvRbBxQVX4CzWOmW8
gxnnfbfDY5R8B0r4cxGttI4i2ttByiRJyQ29q+dwI0MGfQ18dPFSvqNT/ZfyYb0ECJ0aGptR+FmX
Uw3bR57nor4PmsNLYfmc0iDfEaC6PP800i0jEBLxa3RIpP2JN9BcZbZ8p4/kIjsd7x/31zOk6eq1
8owTAAGOjMFj+qz4KLP5L/yPzwLIq9VbcTwOUrMaj+0esp5Q8SCEp6pCvsug6AqNKDJ5hn+u/nwD
hcl/XTn4Odr1RHO7VumVFFRpZ5anNVNdAC0ttKzDe5n2HxQnPQ+a1Z0YC3mYFY3F9NSIl0Xx+d+S
Zph0Y5tjwh1ccFyEgvAdIrF4dyiTUwENUPnG0TrRZ1syi79kSqnl7Ynw6++5X7qtMJbZvWjQbNrN
2VyHXoZFNih4sJElvf86MR5nweuFP6de9q2wj65Jk9ByY8eXTEEDxFpSyiBPsN7G073LPi4Ad5Za
IBZPlQ/wiXjagzwpQNsJZalwGBJgdtmrZLcTxYmkYKD7Hk3YDOq6o3wBVdhqKGJmSmUhEQ6VBPK7
VA79ZUQaNppsI4+9LD9kG0oAGVDgYerWVno3kpmyf4lstqkg7wAEamiDJnxMH0mFld9cMaMqbA8V
eyVhYUN9NahP8oFaj4Bjf/ZMWxvw9ZvYTS2zb30+u+3jL+nFver1Cta6eKCKZ/GBEQPmNVHpgE/6
2Cxbe+D0J1byJilZ5rqomeawCpNKPcOoGNaoY1Tpwj4PwYp2dRc1gVZfrl77m1267REMQhDFYhlr
4U54xKXMm+RlP8AzLV0aEsMQ2ZlHh0wedbCHxOswdm8bdIhkvCcBuhD1CXt1oCOcumbx1sHTrMMm
8dalonWCyoxUoBWc5GSjOMyzD3ssXtzG0z5c4R5BZe2P5A1AZumm7ON12ZL02N3MT0oENZ8M4PP9
p2osCVLQCEHTTWHs3yTelgByWQfl0Cdr37D6SPwJT4atyWD8VWawDfiCRzGZcsc7kvsbBakuyqip
y1KHuM2/LkOLtUNiBWvh9hMKNG00eAkSTPttsMAWDRhnk+3Zwu3xWfXEnZFDAgzMPKgSKmcRaOlR
5++0ddsIuNG+xlgmYEFppCXnf+hQcEr22DsdxF2PeZXGdpkmthTiYErT31nWTz5xX0yMrZpyGNXC
QSjFyNMJhmdyn9piUrYG3K7f3N/dhGYPF339YNTSgDKZEkYXwFJtGqE4GYIcIwmIE3WLX0yr1tHZ
aXlL0mF+olZ2RvurC7Ma2VZlPhfDCmZmfcDORXot8jrG9dwROcUSMV/mV4AEg6bavqYXol8H/fxa
NodZwdA2zfnQk+n8galrOQjfPSAs/MI08txsjwgwug1OMtm0aAFGBV/GZAp236bQM3uhJ+eYpwGe
Xa74HXNSVZa/TXBaBe3FRrDmzdfOVE89WPp2kzuERl7omckuaGqAYjn01OHtHjpSSjSlhIjC/onH
j7HJAuMC+eE1kvPWi59MAh0hVKDERSvNd/zZmEu1oCBb9gFdTNEVWWA4iW6ELcJwHdT6iGF+USYs
YVe+4bQBXrTr2nc3jBdFKDYKEHl1a03Wv1bY85KC1ya0por1/zHs/22Hb6SzVC4Up0HG1pXcqrLy
YDUnnEUIX2vScrTdxd8nXj9y5pp+2qmMHgN8JnG5lR9N2S1lBIaXpjjaBbQaF4pwGHFbsXZeYNLv
GLMikdBHMJDaWV8pL96CUVr0+3CcefxfNaNUmyse6wo7Kpfi20w8Mf0hZyjbgcclQxlqJkS9cp0d
5qJe3HIiJXv7XIzcsX77OZx2UtUGL1GBVwtOhMtuvxqhtEnz7EPIFflQxrSZP0dNUSIp7amDg83x
2eNdtvWAnbvhxjAYSW7a2IQelfOXzuqKZEr6d1EiSPmgNR812n1DLWX4c2uMq2oQb3x5w5mek6xZ
/j+vG8s7UtNF6a3cjb+RUdGGkzcaE/CGd4nDF+R2X4Bhy/dqdxJ7f5R8vK6jqlRwTg9y4r5emt33
Q0jehHqYgy6eSoYI45t13H4aAETuJT3VdAXwR2ZBZCo6O5GSVM4ua1Bw/kXyZxlyPloOoK0hRSCk
+JXmIook9HnWj//ywV2E6oxsSeLlUyhJQh5Jb4IJfNFhkZrRuwwBkQntI5WUciQyLe1RD2U4tyZ9
sVn9L3N6zsZJaMg7eIbRv1o7YwjV3udtTCzJ8IGCkHfICBKIYi3ysI6m/bXYt0FYs6hqlnlF++Br
sbUl8Nu09AEI2EneD0tm8Hcvxrs7PvUKVcjEYGuSk7fJ8wzzAK64q+fIs1RIldvtjaYNxa1EeydH
d91Y4bNNczCWN21DXvXAX2ViL+7vQK/tkPONLofCVgzj9O9XiztLW+ZBssEayEW6CLRtWbHKMOdL
iQHYZkGJ8RJMW4RaPtpczeLCMFM844EAytSIaGd7Fdysj4T8z4YUaH5XSRNeN4+N/8vxZ+8wFN+9
YdAqxuToIwwIPfUqXdby28t8B4yIK39zzcQwTQPiuM1cr6VbcHMHofT/KJuD+StvtzPLInTx66y6
OCZBY6iNnSTBuE6X3IQ27EH6BgxpkQ7t4awFX+7UshgierbLDRFcrKkm11A/DeaXqS/1dcshnE2L
6FlwfhwG/4m6mNENMr6LDMZcImqkb+oMNwi2Cdn81UmlS+oRdkKuvDW8GNQEla6BEvRrsc7w7sN3
+4y193h95HGLOMskjDPAVyQswYGQSZyvaItnAzv/Tg8PHyeqNR8FosxQkKIgzV5hwUK1gxSjK9mw
xxpy/+80v3IdATDxMuG+PaBcHruoeCpOIdNERJtvDl59WWDHcdW7i4sQ+hlCMqeKy5F6W+8ycMHi
QhKMMceV7olEQU8JbAsoiAVqp0Nz4Doi2r16aEOpFbnfaGQ6FTseC1qdvMcAb+1sXWnGfRXW11jI
URKKS3K7TaMxdwxQP+WH2Jj9jpaQe4F6ls+hb0oc5s7epE0KJ6NxfK8JoIpRjFIE8q6qxoO4BNbD
Gxzs9N3uBxryIGAJYddO4Ir6e9dOjAhjIf8k5rXGuG7GCrGWuPXhYtGxJ5Tk4Uzh35j3zV4/SgDI
hoywQUKtKsnSQlyEw+Zcg5Wt+wSPsZ95QiOVPe3t0kumPT8jv/O4KNwiNhxvhkRFq2k+M3Ue4fZ+
OeW6AdU0SgqlBoapDc2U4snzGDJprzO/1TpkcxkF7H7xIhwTSr857lakWa5jh/jP1YhTtVTQdtpV
A18Gm2er4U6DahqwTp5XlyQmvNenaqSGWNE6iyLrNVEYueNOSbu/oP6VdKDs2ai3Q0rD5cznQGy0
4isS7OsdC6P4LtlMwKglnxK3Ni3xZAvJUYVUdSfHIISWeXZU5MhNAz0BzsCmJk9vy0Gf7OtVAGnq
E7hhtM7TRcZCU7jK1cHslTQ7CULDcthpwNO6dewYjomy1AlobLgDkWy4JKfz7GFIIcWAvj97yAsT
/Ov2kG8cEmcy33Onyz1gX4jlMCArPCX4dntz4cUols47gLqpYrJeqCkZW51l3fDhbK9LHDSJnkAq
qwEgHSydUvzSXmoEzu8TcPtzeYnvQnwPl6Yn2g6sa89mkoZ/K0pJTpO8khcjnwU+E8Wd9UdODlnV
l8ApwlYvRYi9GQ4DtWxscdHwauLi86/Gjuyu6Y5/wJpT7oyGHdDPEADNLqLV4Mqd1bso2kyBap3g
x68sjUys/z4EmcUDmlj/mu0ph+vNFxCLfiRnR0qHGzlC09GGgU9vKXBU2KxEovvmwouqtkp1JTwq
dsGAiljhC9qarAUC29HVDwHCuneDGsGYx+MtnGTwRUWrBEAOjx9YfWEkb1/pvZsvietZ/jtPbrWL
syt9hk6Q4GtYx8qvv9rvuYxNaqfcfvMZvzuCqHn2NHgUv71Sp8sCCKNX34jDel1alMgS2ADggrPc
61p5lxNjT/EGV3IJyCwfkCn1zVWN7PNvvY7/IA9vlMd9FJj7XmL3I7tvI4kybne5kJP+rge9Hqra
i2k/nVkrZurow6oscwGyAWVTRikRblI3T1i2EE7xkNzLPvEANBYwD1iVrqPtVACX/XAyu507RB9i
hUGv5cq7tRfuIN6dgAKmi3MwxDUK2qhxBSEnrRfBPTrr2QqXHb0mXE2vGdQH7XAT2/5K6lZVYf4/
BbSSZE+A6ruLi2DIf04jH/zQA0vxb0iUVk4fsN3BlVGvjJ6T8SUqzQ8OFf/mpK8bxdVu/V4ce38t
gqcRdv15ssTCXEl+Tjq7uduq+GI3GLTPNdLpxpszRSUlIsPr+PpZVXoFYveUUt7OdtU8o0KBCM5F
yB8K71RzjiboM9c39tqN6IE+0WmuLfpXvw2Zbtv3g3nsEiITxSrDxIJJ4uMsmsm9bfG7Xhqnpel5
nGcrTcTWIyDtgbXU5dIRnFr394UXaNeV37w0egtwwc8m50LbIt14f8NJ1hQ7DYQDjU5NgQdqqX5v
LyaHHxYJGzxrhBQ66b6h+saNN0RBppcNLxyyJVh9eFzeRHJy7p3eyeImV1iQOTf6ge6WGHTvG8Ny
FMPaIky+rxEEo4s3QpY0RFWpW+IHVrIoZyRipDyKUIgfbL6SOJ0YKvAjCx++j7155wkVGKglehQf
vfcrCtUHVyUKRN6fJuehDdEsLAm+FszcLnT+27uq9oS7sV+wYXUwG7tESB1nBtwRBmi7YIFcvJAv
J4LYN0jInmUBANSI1lskJuzO9umFd0bUK7jDVluT8Ul1oiSJ2/opxRxoVtuUhOwpFKgrgdedEXoT
03V2M+z6ul2L5kQfyPhVT2Wb5x71yWhtfES1Jl87h6M1d4GVsmRgjktUQdPF2sgUyohJ4jsvMieC
EGurgPtlRDRTCWxZTobqP2fvnIM57xIqceibf02RCbCUNlxJj47b6hg8l2t6N2FLcEjuLEh8epL2
YJEcZdVo75ZbZBgOkBveyNJIgMwoQb3bBNgG0qDNUcX4O0im8Q2kuiS19JKgWNK/rnviLtpAf2a4
4PowwD25p5TbkHbKp82eHVH+jDK9jziL2jXA2/5GndeK2kvDdHwXOVA3aZxnk+wB2KWpaHHFl6GP
YSX/xsBLL8LCi9p1yaVbVJoQL8smqVbDEWmb4Sxxv3Oi0U2Er2LrCdhtOOlzScUAwygJDxfBEdH3
l0rFWI+pehrM+7qoI5DhHO9ABwuzdgcZf3Yqk00a+nihfu2Nq00YjMewHvd9XUnmzZicYCr/PdDk
9/LqPQRbkZCbJFcbbFmLu7rKbPgAn3+G+L/Ws/enTmfVuUKcBQDyA8NfY+eJRAqdaVyfge8+ZZCr
6lGSPND15yxxhcYfmmK6hGkjaQ22704YE4l7jNS7sTVItXorOoZkc3HKZB6X+gmT9KzZkRfopOeT
cQMwhUd96p86JBwHzhuJAszjt78DJKXkQyN/6VI/v4duDCIOS0XomtfP3vbBfkJ5Xqv70OFbswuE
Evs3fKoyi/mW1QVR96WJKIaS1pLKMeQd9cVd/iLBleltbXJVleQ2oWqKu7cxcdTu+eyCDpEfGOqS
9fFJ7x2BtoCGwCx68mPiYVOwVrIKWIXbKnXqA8WxLSom8ZFaqyN1W/8T8okHRz4A9cxZuLS2Sc4N
Q4IDi0qMQy6bxPwsVIn2bnPHZhKWcE8z263ZO1Oq7/luSfth1MI6bGhxTvBVZXailMyCOnquyQn1
H9VQSnH6jlrotsZWhu5i6sseRxNOeAc9FI4lBafEvjC79EQy9mAn5cR6m2mdqlCnizy61VQ0yLZ6
NQ3mLGOSnPrcHbM3RnwGL9aKg+EI4PolNeHEvbXYN2GKlhWEkxn3pet7dtIrBuZ57Cj1clQLY054
HRWc9IqpeQevB5FiJDpC7h1VfAxwrAbGkkQ/6eUuzW80L2w9dY6hxHYuoXrKXsDFIUS6O9vPalg1
rzLq1N10SVLgUwDVYBnVvHyc10AW+LnY2UHQcJN1lFFzhfLQsyaPjoSO0f5QUNOn0b8orzjEfbCm
7qPnPT2FnBxfTbCXsCd7zrqxe2MgQM94mpjgyZ1C/tv6/aHNWSwIhVCunr6M++hNCedDvPhxyEZK
fQt9SE4lP7iVuH+op1cIcf5znvGWzn8p++bDJCf7HfPK5ivZqUh1Yb0+4j50Bka/cA4kIJmmkd5i
JGTmszsp91pSZf6cqOSlAXaiCsdzA0KSDy6rxWkW8SC8i/ZQ1bAkAqxG9Wwr+W9qnxB/pxa9O4Eh
ZMQZklLX6rsNsSYHURbuJnMNSbFHLHlRSKsBrIw/Zuj+57QP1bXTrsP3LTnpeYPwdWigToZcwlSs
dRV4DMg8gjVZS3q3uTM2ba2JwOdr/USwQQZbP1CQJuQEjViycIYA+wvK3RI1pDpuPXir427uazBl
pWN6msrsnB3kHb9s82pBB5DF87w90J/eAtmFyDphYoDr/9ofiV7Y44IckQNON7WtI5+Wvd31k9EZ
4P6Va270XZfX12vLnXzTDPdFuqYTpWRM5dzOOGVJDf6fa7+UcmsInCz+WxUbHTrIAb/QTUYnqkQx
r/Uz3f0zDxA91LObh14hnhxSJU1z+42dNOUXiaQ2j8/Y8gK/AMziDfPJo9y3j/Q5It4sTqGEprOL
7SMpChp9qwS5QD2aYABqKYIlK+LuQ+L6ndOrepwfTja1FaPn7WTgHFsVTJquB495Et8J6+9vB3LK
lSLtPhbV0LRtI+SYRHkikUKm+Vm/Qopp0X5JXyO4iObSxX67vKE6umOpqlgICDmJB/Fg+Y6apqI+
oI+ya5/VmU1joaEQ3DFfbhEGBxPU1e5SiPCBJ2i4zo2YCPnrENGDNcnvxfZZHz1ZuviU9z9vMyZU
2W6TtMBWZ4D8AwLJ0jYarEaUBp5ixEp/yfs3lhDS4y7iU+EshVWviXbpJATqho9n+36qRgF+8RMD
ni1nky92vrwcWg/DEwWkPmQv1P2r5ava/m+pbwqXiW7bh6bLprghn/sAjwZicTvZc/5g1lwfLINV
AJXi7a0w3OGig0+Xpy8oWduMNxWN5tGurrBcrLvdzujibafCs6ADSZzsATCYMxvcoDlQwidlAQrg
UimSzIItR5Wa8HoVnbH5sZ+rWPaIRH9ilmT76eDmiJCdFkw6uE8M+k+IqQxe/AyeS2UzJFceoEnL
Zc6yG5YExMphiUdik92WMtde99Fkh3CWwsV5nvvxRKFg857JYIYeIsVKaVZQeOVp2Emk0L57mfa1
W+eUQ8lI/jQoJWsTP01oHeiUMjydgGYIUgZ+ssrPZvGrdc4u9gu41bByL2iW9ADY+XGWiFgkBc1a
6xfOXDJhXh1JRSHxP4zw1s4ICgQ5VXEi4guOWVRNYjnk/YeztWBKY/8Aja6eB94HJRYmFJj6086I
hOmjfDFKL+4tA4iddqlRi8yiAUbSKT3GQZKAuIzJ1gOQeh2/e8kCXrRnHTXR+8iMbBjYV6PNDqit
GGVvbeBZKl1Xe3eIUhdKVQ1l5bUwZnp86Qee9VLl1YY1ewdWwA+2lc79Ww5xQWnFDKt5VHY+6QPo
VFzVS+2aCLgNZXoFlXqZhnkyP2/GJ8EFJ3MLBjHvd+EfSuJfl2CuFaaP+ZdgO3Neeap7iBwsIEyy
rohdasbCgj25ndyOA68H4OOS/cdJCWOXYpUkPM1hn1o6uYRKAWBjK6QnyHDbm8bdlc4vWMqisQr/
j3nIxIdQd894TVEx0MjLF7XygNsXoPeBeaDnHGKnT7bzmjoTZc6VDOt59wmMaFsHuaCwCk7Qlt2m
Q2j2wBxkkg+eiegU2YxOswiovmnr0vdgp0yAhC2/nf6AYuPCwTZkOnS6FLYLyVRai8ruUb83WhB8
gyYZFOge444Q/IIKQSRydfsSIMrkAuO8SWlLKi31OnhlR67rBItNJ2eHeqVFz6vj3AcTotC7pNeH
m3Q/OvcHfzoCWpV/HQwb/FQslFUggPxWdOZMlarh50OwCwNnqAvEOAWQW0zr0qtAYmjb011y0Xwc
b/MOPPMGgfHTGzc+jAtdPIU4r34keDYVnFj/YMncS+dwfgBqFGVzZ5AaNV93cPs+uETAz8BUUgHT
Tq9jj49dzA32ceusZB3s4unDgyCFEbT2rtQ9wJ1SeQ7FJLTcm5xNBNTPC4TXp3UAdnz5lkKS6OBn
SptvQFrqzBMK0jCxWvelvt2Bghb9Eyj2CvhbdN+cjB6b+qr6R9qBq9X3/HgyKk+acGYTSsMGv9Dj
ZQAHiaTmn/EJyXXqz7n8VNO/CHVB2iewAjIGrh2kHPtsX8fQ+ud7MCS0Y/CBQLdJMS0mQ/a8cza3
fs4VqIM9YgFHWEriQV0QbwZzScT1CsxVjMFY9L9vu/Yitv5n4nRWziW8LtET9Cj4bCETQSRo30li
bqN7bCwZXYOndwHsGSQ0LGCc9baESriBS+fwGC529+fivd5FxHQH75NRUZeN1kkvpRIsxZqcYF+u
5WfRPcsEQnjfrfVsLV/p7IYQJVVm706nymCeNhaWbJuSMkqZs+L0a7mC6gYx+r+JIGxePx5jfwP0
rXowEZJ5zc2ZUYrXosBDPIQex5akFusQm6P/zGo87owuznA7nBtSJ5DyUwBIjDOXZ17OoYNGvsYB
zbGZSrrBEzjYEfcmqmC5tZ6//g1Q7dJnIwIWp3DipWv9qD6eveqQ7612W87MYD4JtmnXBJOqZC+/
/SjiNKAF92fRdbyPahYeg/C/ieWsZKfcNfPPmZpbUNp++d/O0C8K6t5wVk2dxEOKFpYKgbZgnQFf
Nxj0A4LrC42Ec5fNoy+kmWaaX6EVHF/n9mvxb5Hq3SLP3fIgGBnMFpEYBq+J+aew9yhaQpJqUANz
sviBEcmSIxZE5FV5M1Jzh7NyxXTmsgN3fPsRfkhv/hHIJqXxeE/DVoIJ+fvOxSZSS7khDerDbflz
vkJM1GeVpXTuIrqgaOXoQNIYTVzkugPb3xnbs0PACjkvdIyQQZOw9uWHLaDGA7EHR+IPzAVJTu7d
WBxih4tD5Bj3bpHwgXSxLeLMvhfyErtBqocrTBV6L1P0YjR+metN35fKCpOJW9TI7Sq6uHr3Ejsw
Ic8vFdKuinBjXAuBV65CQf6M1D+AA7msfuvsOyxHSfWmm4i8ffr/oCMrhY5LI9V0i+6nyQDDMp4g
4mSThbs76aXOCSf1RwSsmnIk51MikNYeGge+M9gAu18QYNc5Q5WxUFTNrsJWfnyi10YMRYurNV7B
SSSbgg91uhztx4FLQPtPk3+vOAmtlYUfNh1ciFshKeJjIq2/Hsv8/tl5WyRT8h8M99BJIIH82bg1
QyTsho14lpaHIBDDL+nGeHjwW+3sb7q1+u2LiqmR7hCmIr7fpBubtToLgIoOYDBmNE+CwvYMLpwE
Miw4bTG1hw+9uBTWWyWMXY7a/yOTmEu31+cks2U74DVJwb8XeywumP18VbMTiHSBRrfMnuJHVgwZ
mdxJzBaS1W8TsVwY6i9OTE6xh2PP6Gc/CjsTwLEIHSW45fFtsUwCc7B5Y76toUo4LmDP3GGAlmc2
HI8bcOU46infDDUeuXIy3cAoJj55rdjV64QHp513B+Pl+IILQnHJxbVmFVQdEWycASR8d8Ay9aDs
yWGWgSVHR3fMd3wN7AUEoYIUeyp2NBtIMMFkTbP/S90Q75TGozhjSgQgsItjm7KLTMBQL/PMJS/n
xQyY7jAPrUkcWrT7QVdGhz7CflfXkUlvHSqcOfGWfu1HOzGpkF5QmbxBmf2i4W1vpGGVzlarqytu
M0dmQplBHtlgfkRHGDu+ytaxVG3l4zyfTasZn9TCDaEZrVCZZxu+mc8wkUShhsX+IgP0LBLaCFCb
msSZEtMuGrLwiExyDIjZjnFZykQw84H8Q0SV55CYc8T7RufogFQc/OhFVZQiIgO40O9H+pN4dMUh
K25Tk9V5HgRRWxTvKv4ILQ3tTgLREstIbQQDjtQwAlDpEDjTVcy5cJDdxSbNrW1GiFq50a5eVFZT
pDs+AAo2p6PERxZ/PjFgDbmz6nzEjuv80v4Xolz6hCLgV7avzQ7JdFEwOj0/OVlGXSG0skpIBjb6
GItxUQ4NGj00tXGCEVdZNs9eoZkJfeR/uAkG3xb7AozbF+BB6ljm+6SFeXqUmpQeeWJRJkjqv7Pn
K2iOywETXTn2AFzH7Axuhl9B+BEMiFF+5Uc8EdjBTfT6hci1ZQfGxC5cyFssF18dygMti/Frk840
YLgVICHhF2X6TC5McQsecTebVhxiucQM940BS1F5qjS+PyEzLjmCXtszmCotDGPoXvkUf6SzvqT8
QuCqvlvoTutmt5H4vX7M8OtdktR489UfoBxDl+nzQAJX2puHBy+r1UGdTCRli+xwuKZ/mYMnRM1A
EcwYafl7stAm4PD+FLSK8un2JtkXkFepzUQCSq5ufA+ltE6EC8/bx+MFGPzEg0iOg2tfJlklByJ8
IH2G+d2DJZY9yL6XxtiikDL4KZtNIWHReQuNZdYyUQ7lzFLK/hMQgqljdBMVy1ugnNZzmmRuvbOW
sbW97AwOTwKkDo9gH8mNFzDHVoRa65r/a8XoYAiYsr7QA764rFByitZzY+RisaaigsxMiB389idZ
1AgYcs9zVs81IGoWAWY3KvyMRCmXhBf/NUlKJylLfj2YuGzA7JewmNksZm3BpZDFJqtA25S3ZzVj
vzmwfM71wo3oLlTHwWW1y/h+ArYz33vcz/xMnsh0YPw78JN2L1pK6BFnuDQagYF5Ejz5dGQZmkw3
r5lqbqDHV4cdJYjir3FTg1WF1iikj31EvivHOMnkjTJB4/0wEXaGc4Pv/S6D2BzWNKYISZgj9v9S
VXXaOZs7QNUqvtJSnfgQtmM7Lx6VIKZlSW0m/CXroJ3Oh538CNfSJsDCeMnixP6O9YwngtwDGJCz
w3RnwXS7j8TzW91OTWzcEuDcMLTSqu4dWTJQV6RAtTmCbuRJn1WuEDiwejYbouMScwVUeCRxqUSr
9kRnmhyeJsNp7DgV6drN/iG/27SOSgSbR6FYKdjOm7jV7T2iMvDm0f96S/GA9Z55TFU1WVADilsv
0gczgkS6s7YJ0cjexp9Uicnfxo9nMgI3L09XlY4cZLSF+0qr6XnlMz5ZJfeRv7Y89vxE4Wg56e1r
WvCvOQ8TLoaOQPePKmEyu4Itx6L3mnqTJQTNYkreSAoijp73uoSWVjYE7baF7/KuNApTQSmW/nzh
IWb79WOQVHPSbPIOy7IcimAvxl5jzFJ45k//VgApJkTuLaMeX4unUAVuhbrvr4hjrXIdNRD74em7
5zUEK3IdO0sncDmh9ZqfEBZ3dNFbo5TjoYRJY5XJ0C8GYFQ3t3NEpIl6OMmvin2YTbDMJOHvrW9i
11ICaszp9jbBCIicUp0T4oi7tB3UrFyDsUxFGHxD8xDyWFaw3yeUuLRB7oXaME3QuRMyMGNgWeO7
DnSnMQNZVNpg2WFfVSSK2u2U2PK5mgXsKTz7ineqJ7/r3DUekwWDis2diIozqYLKXapyD3tu+eJB
yxUatHQh9/h/5sUx5V5eJigKKmpxTHMEchQHpYnrXBHjJLWtIFhAD38p7leIPIfzLpXStTHtaIwM
VmqUi+7ZA+8DwLr/13lXMpaBe+QhZgCXj7mlak1kxYlYjIQlCthKIbrXFw5OEYpVBOxSDIZxYZrn
hW/qyQKTMMX2zN2mHKD70iMsChDfrzmZAmHWJtffIi6z4ZuPUqT8vlH7yLN175n1q7tCEXDf5+sx
K+9rlM6ZdqmK84FeX/hS75N+F9Imi+WilrNj9uFo9aC01OSL6nqMk1fh2Sfulz99nQhhC7dsCoTE
fsby9gzH36KHzdC+l0ZiChAf8/2mMb2bBcgyWEG8xvvRzDnxyNy9NbyuyyOkjbLK6PhBvjmUDsdH
IUMlrP97aFQwPRyw/DjkWC0r190rrqAemKs+zoJ1Yi0FVccUm0tzGQ3jKe0loy0jo9mhVlwmptVW
PRLmp5HFqrA17Ec8kI83TCKFHANIU3j18w6Rvect2cGeIWv8dj0581aaJ9dUhuHZEHYoSNtZdTiW
1SrmGTbaMyjz7tF/8IxkTrmMLtccT1bVXJ8mJpC7ab8vlAIn5F5O7eCHxok0kKIbnY0w2OaencRU
klgndcHMZPtlm0lDI8w2ts4X1aL6AkNyerVJeACICKGMItPld/ocIkyQbu4VdS1ZdXecLeIRYuAf
q1tkp/OwlyT43WXlJZvUga0aFtGCAMxvIrTkipOZ/600o+MmbtlPxRp5ZCZpHkKoEN6FK2VY5vk4
acWXvic9pJv8HJccRFsGpEVTd7pY5CGFhtXXFH3vQHAp3jg2c39HQCpgoHcs+WiKaPBV0Y+dKyav
MyECpOW2i4cKg+KOO/6SOC4BKSDsm7bs+2moRDoDecrpvxaTnn6Sed+sMCbwfYgYDmh5izZch1Q3
gRyhhKg/zDm01v7TuaSVzp8Dt/sGy6iMmUHrleLVtL/4TBTwQB5GGDgJQTabQ9nnUyA4jdpimw7T
PnbyQb57IYiYc1tKfmAOTAN6qjkWYYhlVD0zW7e0aHL6SibBzNXZQVKDlo71Bs/B8VZppUVr5J7/
uMsJJ14GnRJt+GY6AaYNQfyoTaGLVsR6tBSE7ZeKwFJE3s6XE3dX1oMDb6bkIi64K+GcTPnGkDDP
VZaSCOAWWbxs0BvubvXdwMujEjx44ZE/yIcrV+5jSbY30XPYvVXgQJA9+nbyFwmbq1Uq7A9rU6ks
HMLefu4LY5yycMAjBBMhSfLGWht44DuR811W0lJ0DvxPPnklMxeXeCyEbA8NBxCNn7k+exYlKYe2
KD/P3Q0TQcMrNpCwaKNoXNCfWWAn5C2xPRRZEXnXA2RkgS6fYoJ6q1AAUybdOGJjYr+bzez73+Wl
4ctqhNPnZfiGv8o9n0CUnFkokfqQIOmxdpu7QlahEZKunItiAKjgFwTPDzjhc4JQgcY2Ul2fp2MA
YgcCup5PchIQ8z792z1VoziJzPkr4wIYuyzVJmAMsr6RAIUTevLOGJkkU//mLDx5JlL94mk68q6n
8ZNJxO0V1AM5KQYJRzJRxQ8ECgzvXBN7Hg+AdliQK+zpsnka3cb+78HDW+jYYlnwA1UD8J3VESQ2
f3IuAAr51hYJ2Aa7QkeoXwL3tzUIXunaknvWRVbsKj1r0RTnOYqY9zJj69P22rOt0Ez2wFQvNXdY
6HgE+Nsndd4CCm8EPJ33KDWP5xsvE/cA1b0X9shh+obJ6cR5g85N+mXlqzsPn6IRVh8bUs3Z+Dv2
SP6bR/FcWfM2D1gGfW/U8euUUyPTBmqpV6QE0ZlGk+ywbJ1p/tyzlKwoAbxO0/Cc2e3JgWXlWlEL
Tuarp8rnigkQuUb6ZNqyti/7qo45l5TId6TEkR3pjQ/JrcIFyCSDzCxTSg8/hz4x0Sx0mlhQ6yiE
KvVgllQdwbYFYoSAFLkz1dU+hosLQSSio8ZA5M26dV75fjiRv1iWdm8lX2ZliPIy8YpVJk5FG40h
mvorE8TJUUYVrSoAVU7pqbrgbMqMN4YSZjin5Z2t95A0zj9XdxvXFaw6Cl0cexYjZSmXIdkW/DvF
b2iuJokq466Asg+COOd1wGiE37jA3IvxEJJLttRa3mG2M/F+ZjSFzENLv/q/u8s0ufK3yCtcVM8Y
8NYq2eIDBLyTeN8P5NfDqtqGtEWVdyhbUQcRqPnaa8U+f6OhtrLtagmXxTELDpW5+V88dlvfQcUm
UCQlJjdmRwk+aPY8tCAxC5e/UHsqeRITmsrj7Y0Uw5EDdRG4geUFiD2jH6o0U1IwIXPJdNsegKTl
kSPcg7EuAmnQFfEch1baVR9C5XHb/HJ3HWsRqMHhiy0zasRj7Mhf/9gKseYiZSg6c+IDfgx9TcO+
MHMX7FZXZ+WBD5pTnuje79o+mewNS+wVUD20blsxg1Hy4ozq8XSIY6Vee/VB5Jm6hZG6Cj1xjxRo
UoOOeXDiLGOmi/s1fhims1XXELFkgjHO/uw+hZYszEYwqrmQTd08Bq711CPWB/j0eFz27YXf/QK0
+qdyauTgGrf13iBm53WnoB3afGHwAoW64o3TYOL3ny3pEwq7OSZa7u4mn5H4V1cMfXENYdZPfUwE
qClul/py8LLIUOMliAMoemI+W75u/t2BsEXMb/Y7CJ0xfq2Y8q5d2fK+fbtJHtBQCvTlt95wNIeC
nIQDU4THabScEHXKM2BM2+zm2mO4QrR8bjuUuaDk0o+8Exfw1axQNe6Y/GgiiBEeOMhOoVZP5G+Y
zs459AshMKyMADjjev0FJ43V4LHBa1WBhuohUEX/g/576ozoAUyuRsqnQUg/7vnMaUFRx8v4b+uW
K0gAJiYjm3XmSgFQ/7lhjcydPlsuglqqodaoYQLRvwl5f5TfopvS8cySBG6/krj3QqQpavy9FMXC
s4jKjP4rPH4sAgNpFYKzIgND81OoQy/Dl8ivmz35DJWadBjKaPvGP1wJHRjfM4cy9fhwRhC3S4DH
Ic5a9tiwDeq3qYqLDIVm3g3GAMZby6q/8RXCIsSFpQmKUlTPzoOPtstwPajO9oWwLuFZjwz/+Qzh
+/r7JUHWRe/VIruzJWtonhnIauOXYb5ZcTXbPOnweVWbNN00E5LHOrpOLicudx3FrC4UsMEj7QKQ
H7ZmPzWXytOMCkyTxlN+ekzrLz4v5HAZ47JK3xyh6HLBitkV7GYJ976DN7aTSBrRuS6Gi+WvawKx
jT2TyHPTlKIeSHXIznoBwqAAAR21hszTH12sQyAyTpOHzP8GGj9dcM+2JGUVHOny1Tmjj2flIFna
VGCwTo5kzh631Qq2YXuZsCzjJfySx0W0VUXHTRf6pA8uLshP7TdBIPs3ysLHpiyPXIflICfZ2Za4
yVkyjNLJNIeRLStVSU0ke7d8FQ6ycXs8tcYEYzrH5ZEV3dF+fjRfo4EZMviPdowVtRhLA5SePIsN
L6S37+8AtYnSrUsWQqc8nhiTrepI/c3/geJvtXrqa+/BBXVPR/XmyFvYQgY3wuL0Z4GgqA2lGqVS
MSPgTAuPBhF4rqoq4C0E2EjgPcPWLAZDbZr0GlhP6VQR1VuECLxDe8JQFOpHSBWqLFzRNemumHro
d/7FOc3PJwmLGTCJ/ncYY6QR9tDpjBqZXjhKY0ildo9QIP/je6s6dxLLo6Aj9u36WvB58z9O2AQC
kXjBWQP3foxOAeBHa3w06/njJizoUueZBJkIDp6V1unFjfrvx8crdyyLCFt+Zpbe8rykr/qhts0s
tP1jom7qNJN5MZATED8RZt9KXcIiZ0qdSABqCwBIop/Y9rrv0f6//cc3Gy0dFlziD4TSrWPMocPI
H+PkCGP3Srrgf35XBHVRq6Qm/2yHOhz+SZkqDU/Jb0VEFi1gBZJNE0GwSylsxwtC7XpwaqHMTQqF
rdGfHDKHwIYdQMi0fpKvjHa7VIe3uPoD0QET1O1IWp2UF8ClB9ae8/Z/eQFav4lQkJ/15yaZBdVw
6wWw1gW43tkExFsf1yXCO8hn/bG2viJ9NH2q2nMEaI/ZpYGsSJhJ2QI10Lc/Ska8JmLELruhbs5x
YcDgVY7SX7A8XlnPL1jOvrxfA4pOT6X7hEPFny+edqSmC50PqDWe0dudP2Q2gyulxTowK+UwjA/G
hFcJLElzVLohrswyG1rxq99xkbylSUsEwFXzt3E0mwYdZKPa+sySmm9BpfvEBKEwX1CC4oWZEGLf
sa9hZP2yXatDKrtsgGOb3us3lNH3YXAafl2v4KTnQ3USeRuVRPYd4/hnhy9t+8/z19FuGN/FgqUR
OQHahzOwF0ZydI6jNTZHKZ2hiaNZSjsERJtitfiSJQqdCB3ogBK3/1MnzaOQAShmKOqK0OO2Z4AB
2+POm4/nwruUCSI7Az3K62KWLf0RHpA+Pdpro6oMNGy795XZF+kkt8Mz3SZHTudHEwOdMolltMUN
N/ulnSAoCiLS/oJcEiXJtYUIBZAdPPuoONbFQADRzfXyiUVboui8zol5BiFFcf1NAGNSx2pVbRBA
/1uSfVlv70RCVJnpd9tMIJMix+MU4VvnL/KEwoBNhAWnXQwf1cKMDF5UGu6i6BSWOdOXs6U/QAFY
StAcifpQuDPtoMXXvryE+tfrVLtDw0UppcQdkQlZJ/lKWortGLDBGctYlZX1M/XMPKNlT4kFizqV
FnBy4L5KO5MEdaWCjH+U05id88A4VCWwUHhK+NAl9QODiCHVxAlWfJuX2dnZzAmSoYQs0E1JT/2c
bH80/lkN5eqfpyqiJ5/gggX6nMf5u7DCTv3TvASsz9NO6xc6o/pHN5L+/nJSoLuS4vjB879jdRuq
oBtNaH6IS7T6gSqM8Y15Cl+ZAA17/zYp5f2o7Kof05jEdzvVwbetVp1nIW07OO/m6Q6PGJ0oTb+9
jQrIWlIGbZfvDZmBD8OMipQ8+JWsJi5/g/F1iBSPsp2ialmsArWH8Sv+00TgZBsClYGD/GZT5BEk
1xotKwElSwRdAMp7YJDUMuhAjSxiUmMHr2xGDw8QDRbK90tRgMEKWRTcNt4NUN+F69JvW5+eAc/R
hw48fqTWYS7wXgR9Zdjl1rC/XtEbHK/0pb/Gw9exSY/mBvSHIeZtdBdIzEjQ63OeOdcbQY880u2f
ucBsMIIhO7aL1Ruc1/yEoYdxdAFWcw2CQMJabreeKLP7OMKSLim6f+BcNjDGgMLv35N5ggFLTQpY
N8kr3TXFOCAoVxp90i6/R8IYQXgpUYBvm9Z7mYqqRFleWK1PDh8zQ4L9gu26dk8o1pXz7kZcTe9g
AzVRi8ITH0ISH67wDFY6lvKK4gHcccS1K306YGrn8IElY1Kj5Gw85rVhOlrxuYoJ/h9uL2MPNniF
cH6gc7ugYAYeBX9ySlagxpZJZWZIbN3qAMUanvNbIRX+C0IEFWjSmc47WGIYX0Pd2nwVE6jJkd4T
cj29/NEStqlhYvppI6KIvlf0nB0iboY8Cvn5WFO8N7FLsAtwYx+IgIne1nzYwTSdCfZdNRwEirFR
wllQUNEZy/I7FWtm2OAP0HHmz1GmRhjp5eVQ4z+TELCx15kgB1RkgLPcRfIBXgCsPUlhbW3Sv4ib
2GBnmOXYYC4n7QkL8A3LdqdDPypJGLXbs8y+ScyESqV03xeTIT04WqRJ0mGzLxYAiCbsFWhUcNn/
rDktFg7HaIw086wblbcXFVEn73PrINb0PfpRP3xliz7xeDaDhhQTUGmZaTXPvk8VsDOCpE2BVXAx
11qUVpB3tzy4kU/3SE20MTTo957lEQPkyX6Zph/Tccyz1urVUQ7pO3Tg1i7lM3E6z/mFTjO5kKX5
RFrClyqMqXzaoQZzq04HPaQ9ldh2uybHRZU5yW31E4iMjXchaqL6ChgrtuKAEiOFjID+vxLHkx5q
G2akA1ocJInkGRdjfWT23dkgnxpVgOsxG0tHSHuj2bFyN75DnCp4LPVt8UVxB2o5SbHQI9NcQb/K
QY5G8ze436XyH2dLyT2a/I7G9OrE6s/98Y84pHQFAh5lgcfEgu10upbcmnNG1oTwIYoHnw5OlOuZ
UM0YJWVCUnoZ4aBWIIn9ACbTNnzvJ2sjWpbGb22IBQU8qTuTRtnmuMm869U2qB7ZMgiYdibQPLlc
rKUm0HQXgQa7/MVolnQt6QDpSe/4MUx0pNAVzZkkrnjjc4O+xtbWH27xYY4AqY+P9MkX2holvMMA
9u3c4bBkOogQcTE9nUDwaIC5NHaQeGZTFvqCDYWwD3QI8pMiJodRXSR1OcJ2M+7O0WR+X7lN/YjA
7MZlGZDZYN07WyEuG6Gs1Wu/2cW3Dl/nWbwpTuL3aT3Dn04dePCWxLHJLIYkVW4Z5ko9GQiiINA6
+pXQPYJHGQHkrZOB5/R5UJwosfP8td1VlNMD2tML5bXTKzkPRwKPUDCnmWlewPa2LHjjUzpPSHcr
MEYicRHlnQCTzXBAzl5ZGacBOEJ9f/fBN3AmGq+WmDetFEkXwmiK5VFECV506vXw6FZMAu4Mi+iY
ZeBQRMbjMtMtqfGbY0xcl+bRLMBWMeLsmxWoKJIIflLodpDLdszhpNIQIwvMokO/ahHFO+pwnWKd
ANaa0jdbSxHTP+umm78lNB8Difa5iFwLJlKoTCuOqRK98f5lLuZ1g2Ce/5egDu7C9J0wclpmVEeM
rknvAo9YGtCHzfaoaDItlvX4aneDwyITqAZYKPs1okx/0lHxOOUmlzaRG7WRG6nYRcmXi0qB0RJO
RZbDVe6XTUxEg6qZmdWDgtJV4nPeNhk5C/SiIRkpC/KW4uz7XodmRbbkgwfsP3mUzMgICoxwkEgE
RQO1LNNOGvFmN8O77g5OSm3MsrxcLnuz4MgDEyZNRDZg67yb4g11OOYI3xfwHuxM2kSI+DO+SG6u
86CV73qMHfSPfvWVhGZYwki2r7apDLBPx5L0bpVqfwfgv4i+EoEVtr2lZ0IQoUXro64bw2stEBpN
KzZts2Y7pIkNNSQSpqixGxoOsaZXoTOsh9F4RlGr7HH9BYKoBBq72BExPOFF45F191QkXbsrPnKL
ltE9QwFdKp3uQ/gXVTZI0HT7tQjsbCz3sm6eH/pF97HQCes003M/xmtgUstcu/2UCpzPqxqZW6a6
OVdxqbhI4odpDdTI8Jpibxx6OMbaZioWgc88i3G4grvLhuO3xXnmXjUCgZUXKN8cBLZxJdgymd8o
2ryIX812TKgbcT834oD0qC1qcQoh5OGsD2RDwghbXve8J05vD+uNbtch7XRAmSdNUY//metbjgPD
xwaRVEksoOABRgp8C0ObOPdoz3tXtP2oa1h4UR0mbsnGCJX/iLG3asYUtob/+zRUKY5UTgX1mDiR
LCPLIueWaVYArT2/Y3abVunE6i1k16YYp4WMooEQniHByxEwiDO8lzgCa/yhc7dvvR+T1ftuL8aR
PSwcYdzv20dbc3MsxhgiVtm8TtBuRAKHvrYsb4tb8Bq4OGhN5Ew/f4Ckqny5b4JjDZ1l0xg/w+HG
pH3QDmqcC50SERufa6Dm5AN7o04jsuj5oVMgZg5gXffqhPJ7EQbU82DYCRVYxLS6xy/rBdFpHxP3
0JuWpjaIXZyHRPUWrvAwJWorDU5MrHhuukGuEoFDixomn6u9lgHlYEWfyZvn5HMghJtOlTDArcdu
GYAUddeNf4yaGvf2X48U16ZD2lyQUqjmxy5tS5iRQ7h4QQc5n0X4TIDX84BUPO3HrSZFMmB3uiIT
0z2OFSo+L01vZpUcFMxICGZ2FjBJa/36DMwXkrMoyMmw5rMVfalEEqETC8K3U4ghsI+G/Now/xV3
VrwdLpULuffqjydsYEWY7ZgyyWvZBU1ccMZ4CROI6zE7WH44/S8zgjFUaDuOJ/YhCMpPsnF8epVH
5Py5AO2TtByXFbyKJ8dPNSaGB9563OFtLeHaC3ZZy4bSNO91UnujWtzm8nMNnEBcow3iCrag/zXe
6CR932elvwITmT63DbQYj7Eq5hpGd+ElSppzbf0PcmUyrAL1652AKGauZ0V9lL96Mm39RV0DUsev
w0EDdZ9MNX0ZcGfWPAzLmja/SlEUJxdKB+IcxXlgPyNuqMa6D/44RqHYFs7uwAUxR8onyVw8dnBO
W2pyUWQat1VAaNl35D3Du7TjRFEkjk3CTYTPjoLliVAjGEeujdRAy3s1UPb8ZeSafvI25axY5pJH
DLS8kNEiH2lrqUaE7LfmrDeU4EAfoA/pgVt0L739FWo2W9jdw2yiU5uX0ECbjtq4iEguwPMgmLzl
5RZfCs7ZsYHtlexGLavrcixHQOCoG+mGmtNtK+KTXjn7q4ENY/epD2pEQeUEwJbyhsb/DYeg3wdb
Ca1LvLBHn+MdKCctXa5wcf1ksGCbXLHrMmzrlt0AGxC/T4M/Ipa2kAGurItTE4ImChtK6+jngzyR
wmJN+M7BiXx8ApAet49rz+gNYpGjq7V6hWaCST/ijhOm1w1W9eDVRohC/Bk57e7aLz7fa7EBPDOd
7+uT0ZALNHk+WFBBfilPyxwmE/YtAxnAxzZcP3ghryvj7ZV459ik7acQVn2dlHhahCnS0uVvRM6B
y+o2Ibwv8hFxr6wzhfunqzgFJaAxS2AAkQ2VWwiEV93LXujU+xbXnyBPD6Tf8g1M6eYmBTRa6IJN
AsuAiRbesgIbwueSM8Cw8R1entj5pB1r/TgNhQQbmOrtiMJigxepPJ6gnTg54ztXfAenUsHt3X+9
yvrm4uCuLe3PI487b2RPWRdgrWVNaFSSbz1xA7dFVDfbIyU1fgyv9aQVqQYYIQHJyvQvKk+BoLbP
odp+Cib3e7Bzo6n40RfK0ZK4O9VvvQymsLel6UqpiyeiL4OecfgXP1rPk5V1FcV9PCGSHCW0/dky
R8qmA2MHPT2dgmQzeUm0sOoX3Gt3yA7TYvu2aQyTkPxGpSFbv/tTzkUuRs1HMNbt0GlvaS8vaTHs
gUwgtMjHBCqaTegDCuMhjwHiS6YdvNqsDs5nvHG/+ZHQA/oMXiguXnEznseYnqwcixZeLwLMSyQW
X2L+mJMSaekWvIigd3ENn5zomqLTC3LKRwbGWu1oXEfml+S2g7N4jZebgzjSiT2Hcr42PSuVsH1+
apQJP9MWs17gitHYyi/9oaz0Hv+IMyIUzW0Zn0bnkFPpLO8BfvTpUaz+F0JN352PQ6gv1MyB8ULt
IWhE/i5UUq1bhOYroj0AAEd/X4Ky39k5SKdtVrUo/wHvtOOSyanocwzMeAoOUQn1ZD3zDD2EfIMA
G9+dajLkTZSaCBS/wDestd4/hWyEeK34rddizsrXqEN30C3e7yFfdl1BEHoVjNoA645MjyhorgYV
LoxqbLr49BSYuoRXZ7SFsmVHytBgjFaL754JdOld4njcSVtaXEaNzrGtOnKAQ4ooOQMP/jIK5SNh
pi5FCXSCnlW6rx/cSBOB2bVfpEjxORZ6eMv57MUk//nBRB01ergorxfV9Y/I4ykL+v6rtmjn4neY
LBnt5G8caR0d9phXV/dcdJEWhoMBgWgzX/nS8ITCY4+ApHl/zNbs3idXF3iZBHRzM8vWI3s2gTtQ
re1Slgv9yQt1dIdOSVpJtNs1icDFY52iP4BADXFm6smxyr5jikpSAuPCtipX8fJwstGyHZq4YlN9
5/IVXoHulMGEiq0a8pQpH/78RYQhqU1XbrNBLMFmLP6OphTZn7ke3DsSFn8gRULRpqKNkdexb5Tq
gYfUiJMvOMsRFZFM0tafb0qw5WjF9JDB5u4rLhbcjostFzVduD8/vCFP+bp4P1rVBShGGUF+mgcz
8vXh33VfM9lSD3kzEJihnaXAVdkzR3fqYDKyobUjN9B4j/6aczXeC/09wB9EnsWAjZJjP5W2tMgN
qPxFvqIXh5+OwOAVb+0RLUSOpIIbMRIyX3PUC3i4ZW0/tO8R+uxe1+T5yKbe4bXHPD3BGuR28GrS
GSxO7HoE9/AX+FBh2BvFlIh93o0WYZY+DmHhN449RrPFVjfaQCkpu/gVv8n7fZPSzDGOeujZQB/d
Lt84A0xLumIFezbsWgAjdSDBoKG2g3WCPNY0vLsinDYr32vllrthn3VoSK5wToa43DGYMoRJ+xaC
7TKJiAnpURg7i3Hom9vk+sqvxUPQ+6hLYYmpR4w5h+2a2VKGatLIEM/LstCBSg4gbrCUS1NbL/c0
AspaUeCSlF7FGEpszaHq0rnfuiDBgwa3ZhooUEt2hP4kg9l6VQ5KRqrkWxBi4159T/doVQvuGsns
RnstQAE2IXaGTTNh9rQwAymOLy+46r90KLXj5VGRe66xU4cQhJh3TG7+YqwEkkqhIHQa2us4qeMH
G9h+XLD9mxSB8/dHFVS/1SmBsvz730uDBY7W55ZA2/aMyb8t3gq9/w+hPTY2NGhu8VRKwUDlwEuI
YsPk1fCWaJ4idOue+pzBMsGbPSpTHqh5lDAioIJ0Qg0uIzPpUcUm2hfNklxytq64NmlD7YqCP7w8
/1EnT7ZspavLhXHofnRkIxIvq7Y7Nvp/uYGgoMK/S2BVo0fUJQ/5Y8Glkci9XG+gsJlljyN9//WF
0ehk4t1zKeOm6FOMuMPkSSyRHLYzAYhdcVHLd19a8i9qG48mZhrZ1sqJVFbG2PxxEpy8hyxBiw7T
pbP5EffAHycxqYXxaNV38t3VUssGydg/gNyBzxpNXVHpAbWb+dAU7XGbvOyen+pwUwK6tQd/G9VV
Qqvg8527H8xeVMbPyB+wlNgjtE4tTQb1Uwv9nHzRqrX7W+EtiURxljlSsjtplkVvaEiebyo3Hhkt
AFFnKp28eW4P1TI/RV40M+OW31mPdyvfltHZ9U2MqpoA5Qy3gy9Xc2srgziiHF0pcS+u2KXJoEu0
4qZu7woRsA978FfmetXwWglpcbom0bAcnoj5VtnMmyRxVScRqHWhrsg0S354EPSPZ9N2XLIcgX1F
S+f4q9pMo49r52cmd82Ak6WABJY5j4JXY/oWTDZwxDJbhxUAwimmbQBiXF9JsYskX6cfWniaoraO
uwN7fKyWkORg0tgQ2NivFSBg1GkWi43njSCdSVNuMBw3644S/yIoBeaWfNe+83bscj8QBHtPd6oa
KHEY3PL9cAauybh7ELCOKQw+8BmB9JYi+CY1GpR71uYgXmXrOncAjDAiU1yk5wAxUYl3Yal8ivdB
eUQYYGk2DVXBxfy0I9rhQnCTi6gmHN1nDqdNmUFbi1jjciM7P6A438wf5TGFGl6XTuQliEAutDSc
D8zv/vy4fLUFBLcnnOZRW3b+vbwYIW28++Y8z73SbJXsQgETuDNS1GSpXnePUuH3si/SvVxipBRD
4jFtSLj0CQYgSY9V3jgeyksJn03ojYbd77ZhcPoncDr7lO4V22y7HI+KLbcWo/ZOCrtOjUkcO9EC
beguZz+5WAeCuQtwAZ8JRg241/YO3QqbplS4HN1BBsyMFF8x/lyj9Kv1jtjxPOuDPSCg+ncIpBYf
mWrZmmoEJdV6gB0hAd1wqvVJKDcwbmZDPKqwUTgrW5FWP2nLbNTAftAzcajosLiin6lAvhOA+ECf
mcYyt7nLUnnEP2NnNm1z3JgxNle5DnpX0sOrr7i4HSMgNwymHJ6bxOFINA/ktJw1dY7z0H67tEDv
kN9hmIoA9DYBivDTTtmi6KcZXbi51IRg2TjPijJlOVjKi/tkSQiFePbHmmDwIp7l5QNZvDZLCpFj
6uEkvcejGxNYfjDX9SrARL+jx9UcDvk3wLnO6aHIDfrHvFJeXvikD5OopGJOzW0Z0iHe456KOrp0
sUMXvN48az9tzz7iWEz1IBaUIH0TF4PZ40OysTnxZgKt2r4M0Z43E/Fb48mIDfzZZFVAmCVBFsjo
xA3w+Wcs7NeVmVk+z3SBEoaxwwPJ42dHlMZ5xFRt3FkPuOpmbu8g9JslXIfLIOdIM9PnXzoe34TA
P0fsOhEe4nG0+UUP8nIZVNmduS/rlij64cxqp9FcCq4WW+SlSbpJl6luinf9rkWxQfx98wx8N+x0
m4zQQC+lvrH7e3WbwaW/4cbDFo/HtdheaaXAN44ijx3IC5lW3ch41//olKEuao5sFCNE2dnOe02K
3NxNN2lWd02RvszKZHHETcCL0bS4fLsXJojzkLgbseTYjPWeHoNmbqW1jkUw3jJZgiz4EjVG/9TI
b5etVURUoWchJi2Rs11Z85a7LomtdHWIooNtt5RNeTcsEeIa9faLyrkH3mx5/PS5JKhkNP4uO1Yb
9PeO7/IPcz0r0PUcffXUau2KLPckNS1S20rf03EJ2WXQR1yMMNKrdwQQ7QcMipn8JrpDMwkSQh0X
7qptmQERcb12qBcA4kgueY6n2jX6HfGdcdoFH798v6g6Z820+Q43yaYIS5bLUDUFeClZGPGPqbOv
WJ9OvLegUinW/Dm4IjkUpLtv10TZX+UF5mG4eu6AL3J0/GOKjIzwNzlzpjPKMeV+IuwWjHqKMzSx
jp6S3DCZoVOKwkUJRSo8lNyvB52T8iRGRPKIZWPlaKCYkSBz5+Bc2Gwfj02WAF8kM8WjDgn5m2MM
Grl+B/a6Mo/QQOMwOLhtsLF5XjI3SiCM0j//xnxX3NaD/+IPoh80YhvDumfDz+UMqL9Q3kfvVseV
EXZcV2yYw8kYuh50+Uolqd2vbjRIKWzQwfDy27ADFy8NAMxRCOzfPFwp28CLwfcdyv0fBuWPBPd5
jZs0uFuMqoJ30UHXibHKi6lui7zGhubdMOv2e9l7LpuFOxCsTUO4XvIOwkNtPpRHScaXzgbYgsk+
9nzRyf44aPGe9cQSawj6Tm3bAGCHwR5lUjUnfnjWygHZFParAwJuBkJKAfvSOGaKgswCSeA3TO9v
KB9S7nZgN68DrGqXyQzxM0BA27FBEElOPC09Zjgvkk9vlCOZyGHeZezCqp5pafdux58CsZKNFS/c
tB1Y0laogGolDWoMyD9ZZ8Qu4IuyrF83oGI0WCLfe8xMiUhf2++rk3ACx+CkPS2wzghmSzJUdXda
5W6K96D4HFKpYXiNF1LrH0T1yQeXboAA6jvnB/OSweRM+6ufGLmNb9P+myB8kpLZ8gxx/ymnbUmZ
5UzZnruXR5TFeQGe7JPAACCU59hB+3v803JZ6SqEWsUO130jap2k7a/W0TfnsXrKQYQdcah81jF6
nKT0Mzqey995ucJGMhQIZ5Yq7DZqcf8giyZsJJE5781LpVS5Pkp6kx5Uk85CO2tatHPT4o7BLPck
VJNA4h8DbUI9wZOPufZmcv21zdGcVU2Md+tn/L6+BkDclkz4R853kcXyX5KyD3SVsJTTgvxYlrZ8
4qJm5g5z+YwA03Z/+P2HfwzSG46N7bxPlhQzjPjgF0gcMYW7G6QU6tsudd5hDRzTmWTHg+BXTVhL
UiQGIqjiahGGK/NPRufn8+ETWQigw5xhZR3IIVIgeR7GluU1sPNr4W8TNYSlNDQxAcj13Dk3SkER
l7qQl/2Jexn/jCEwn3+sB4vG/Sh0r+bm5alD5zAwfztnNsxY/gqB67BpYWjEYFYCPVp8AGUWG9Z8
MYsp4MiQpeujOxNwxPXv7CsB+AbmCsdK2g0XJq/vJXLmEsPvxwzKtiJLHFh2YEmZ7qB1kprUF39+
yB63wPeLwTUKBRtJbxydaSk4LFFXH+aiSmGlSvYOoO+ajOIHjTw0CHoR0CfOXcOnQUuRZf7Ll+cs
rvybOnFFONa7G4jb3KqPIjhe4B43Ib2nSKMxhTjYgY9Uabn9d3II6fCqMJncjwYBdrVkLUIjZP9Q
9u60uk4v0IqHxVxExHVhpVBvgsa372QCqfHXpYI2plAAGpRGl1PaMVR3y/ydSGCnRHs1QMT3BemR
v2ztaOMlpMiX2g9d4OV9bA9BPe9fZwoNK4fpaHqL0wEC3fPiRcl/oN8clDq9giJ0y+KqI2a8nah6
y0rmK103x1b9X3syLTgAef4Mydegu03M6YJaMmweiqvSsJr+bAoez898SeIgFf08NK3fABMDv/K+
BTMIRtCGjevkc2zyvnxnI3Lnfsm3shQWxchjxE6YkJnaerfhaGggXLzohiFDDIX2bVAdMPGxBVl9
4hJo0GKLdz51WY1zTitBYxHj5B/DSv3bWzX92OxI8IMuBDK0jo9CKTEzjly0ez+ATwzm04P/MgGN
6pEghRTwW9j05FKI/2Q/D8kRMluQ/DL5kZU3VbA2sDZZI3MoxZOdv1qbuVY8emcXBTHBqPZLVB1W
9nn8an3FGgrRlgfeaNh+Wbfphk3gex6o9CLidKcNrwPwIoGvjVCnRPDho2CscCHqXgVVYBbEHUWm
rd0+CcKRoM0pfESRHtEt7Lfg1/7Qy/12U/3+HULBmXw0tvvt7KzeKQBrYI5E2b+O3LpY6YI/QATK
kDEXOi5W2PFBF/l1o1LZti8maCa31dPkSxyU32gv/y09XI0sr/1es4KZ9k6g61/toPOuhL+53EXs
uWJeENAc1SlpFP8QPlDFPQ4CmGsqTGOvrUjodM3qLMKoc6zP65XQ3afOI6qMuboDcNu8HeA4Arvk
PeaxgMajraTQ5KT4fklADplJfJpMYNkGTQcotqvaeHzHe/lQwAV7f89gmwiYDtglHBrLYjZG6m4D
Rfd60c9xt8T3T6EtQlUGknHjTEaavYitj/Z/yr90V0dmYPh0dY1SjTOU2g1NxLqlh3JeeH2Kgiz0
C5FRI/FmLnxsrErAL33C/Stw8d+GNKqQ8DgZnZ9L7PWxAuoZ1uAuokuLzpLOOW2gZ62HdDFzn9yS
OPEbZdBtZCmJCXoq8kP6KXbfxcPIcL+FD15/1VEbEPSa6Tvdf6wG2FM2XxyhB0sa9rimojAkcYXl
N/qJoGqOQsJnlGjesdXSsRGt8VjIcBAV9WOEwnrMSRTtg0Fsa0I1aaqaHYPTLc3MxzSHuX79Ovhj
YXLbj0cSQIS3Gpt1cwae+k8pwwTvt8jHjsoNsQ6n0e5KUwLVcJ1g24J4wc5xHT5xY+wn6elO/a+C
7WybSFjXedJYmbQtL98NossaHWK27NmBsZvXsAfLH1XMfMnc3MGbf/SmFk+lnFc3J3sHQ/guqHpA
JYKvKE2tpnSSizaMljgkFhEjR2Nbnjp94DjDkMyfNTC/HucNYidCvDdfamQFNaCMC9CHCPMBlOUH
fkY01W5IcZFF9dXVNkrIJlE0thJBhVDbRIzyYwTFtp5KT8IK8aqxY87teheQvukbmAsryQJwsZmj
zesrqHET+OXCAJC7RFSJDBzYzODTpX+XFirJubzopWzAtwW2d8kt+633OisVyXyt1dgEVwBK+XaN
N1LrN+TR9yEVQCPPnoKtNh08YVuP7YtwCKYi9MMHF3O1jJmehD85xpMtjYegYvFLUBSmlCCBzik9
ARhYp+RwTuFPfYLmMB/rp6sdU5QSwQD4xnFE6vmm7zMjJPYeNh+yBS9GT1zKOd5w7+dSfwBaR9gL
s+6EsrBIActtHeuGMAuuXiJZJUuRi+EKzA2lESMP7gsU+mxqG0utZv54P+wjkXeacS1iLAe7kv88
HQQmz8kqL+Ib0PbyYHG6o3YO7WuemPJiXFHL7jYSUaTfatqF2RwDNIQsuwvcqC2T2c0DaTj+NAPx
XUFpid6ph7Lsh5bkhWdcicZJ4JLg5OCIQQJbm42E8O4EWp0hNiBoMktAZypn6KYfBWbOORtOBQ1+
+MPLuCE20Wbe836PE2WbbQu+1Y46l4+D6Q+DuH4HeVD1+k7dqFkt9/tJiKu4InwZ29jA1TL7vJzF
EwCBX7yC5+rAMfOt2HN0j/YFC127NkOBgRG/MWdgdsjnJ7mK+H+4J0MMcL9hrW/MhmbHXVBAVUI5
VfrYtbAEFF5ElsZbAs0nia6hg8dCPLe54B1I9IeCDj0uETPb1jihIluKLncWFQI9oBhxZFvZ9SZp
59v9tA9S9ZtVSn2iwKb+gkNHDOR+emd3HpEEG/cp866tDOvIjREVKUk/EydpyL/KfGq5RK73y4VC
/C7s7L4GL/YNshSzP5RxIHzrYi+hKioOnstqNB3jdOE/aDRjGtMqZPjJZDeJedEdlHf5t18qLW2B
mgz0yKS/LtQfUVYS0LAlKtzeHNoAktWgcPSrG4UIwB5JJ8kkTPGKo9y2OsYilutHDaZPNjiOMNMb
0UqeOHfdah8AMkZivKq0HzDWlgyxvquz1w+vg8W4ozx0uH3T/0UZK+lt51t/eMpEHm3gwFlTLQZN
AWBN09f+xEnNcRhat7LVZUyduOE7Abq60sfUDCRMucq/1dNdAkRF+d7fVDwYjot7NepAeAZ78ihC
/7cC1jFtuAQ+iUgxu436cK06tCoznH/2bDHeuMnKa42TOKZT9CyKPNVp1S8oFS7YZOjaF0xx8i1r
mI4xCbyV8dziCosvRqcZdxuzorRUw/TD9SC9YK3XvYqqDF1LBSvAVfGPzodR8OpCmCp1fT3eZeQI
mgFvgWvKbJD+tKn7hJSHPVsAEh4jZih1TNn8dGmxZ5KmwTZsDgdL4crMFIH3dOGy80WMVAOUKohm
6bMPd6GaA8jY8HR1+uLpJVpvsgvtfAzj/O2r6Bj5I6QynZ+gMezcYWbOcMdnvlbVvRsk8zEMXy30
oLZk+1eSfmihZsr1M0bfdaSumfIKF5zygOojr7i1deQnDGHMLIINGjqYB3PJlVVMhUSmfXPArSGN
fhF9BL5RaUV00gc/dSVDE5I7NMPIoQyTkSrYMj1aM4v2Fz241nzZfMWsE1ZcZZKsURnTJvI04T0U
3Q6QjJXxjoADnS8B4kgzaV8h93ofb+pgEb9jBebtNPQH4a8g18EmrsyAGx+ZX4zyEullFfJPgX42
oC7/B5JAlGSFMp0OldMtLOhTIijT831kA3lexLAK++aIIWS6zD2CpKh7iwa9q0AeNf2LCFf0YmNQ
08iSJZSXf7OigmChwMv+rVpTnwhBu5hQUOaeaQf3wS8qKRpvrduvFEvDn59/uFmnSABnLFwgTrjj
J7kkw0RpzGy0CyEhDyCYGc7iYq0jBKXm0T0cawW5y8HQri5f+ejD0kkVfYwoCJi0hJpbpxEMHRcH
hEXKfuVfblQymQqK0S/YFxvRREwJf3Jm2nx9vQaEYdDiTHWi0bv3iDZB7hb6WInPY8AOvtdgd8SR
MH5/6CTjWSZlY2aqlr5hBHPpA99p8GSCbqyKB9bAAK04OI+xNFRyVGjtCN2ZpsvRD7ldOsqCEV0V
WUWmDb+28EeAWvljHnj9k8KlYaDojivqzCk/C4iSxTmiHY0vF4aCXbB83I8WzntRviCW18wneH/6
9byELkzYlL08lmWpxFSX9S0M1+MKybG4g5TVbZS0MvqTviXgNOu6FW85u0CQXfTkpcTnrL+5LvXR
h18nKpEG3AcCiKzir2iKtIK6mRyM76BJLPQMgDW6pCZw56kHvzXER3DRxpis9Qjrg4AMQa+5Slxe
1orrjt/8K6HGV/yFyZELPZp5XmQGNZBYrxHzVO/DrJo6j/qHQOkJxgwgRc5lR53nSfE6PjJaBIIk
tLpZ4/UygS/Nd7OgG3GtxK2EWudGQCrLZBBDyN7/32m51cJ6K50vT4Cs+w/x4lZtJhcC4CDwCD4O
HQCGuY5N1qTlvqFo/zWZVz8O5EYk5zrvOnJzJqEuGUxlP7rP54PYzFZfurC5zjli6W8cwC8IfoTw
b8xaFKEW3XZ3YlC1TuncisGemgDt7maj9hZPNo+HP2CaEkW2WLk/0ewKhNND3q6oZwmQEwWDU7x2
vvqOJnxWDy9QmhDA3Ivc5T+/9gA3terysMkjpCVAPYujVBM3OdmPBpAyasd7gu/pdnzK7mZc9dDw
m/ACz2UI4Oeuw96nPLCmcEYoMqFXboBx4LU8/Gjpm8mWJAEKQWd+zOlPiAR8OY9IqoyuwSHJgUxR
XTxQLj3Ta29eHZJ0T/tmhvIc5hqpALkk6dP5AA/nBk9wdVpXeLs5fggBETLWHDS/z1qsM1Jduy+N
7hiUquHPS60OHhWpTsM4Xm7mjS9xjHNnjNMjj1iXGKwlzOQE/qbxQD8jL1+oPwv1i5gw6M0BFdFt
zakc7W1L4DnJzvLi7BYp8uoG7yME/OMpJ9TK7oRD4ZQjUSHZEYqcIUcIeUjl1nYZj4su9xsvi61J
f1WyyBbAbtvsp3TVOR2J7jC/0Gc89iYE4eWY5xGC8nDageVQNMLtuXjwz6hEpQDHNOicEAXRysfZ
MWwenE5CuqjbUJ2o1RBC/m1UsvXuW3JGJR92AKsYjwJS08frb/lzqj8E4GQi0XFr4QUsjzAis/Do
7lo25hsc6uraD5P2Lf6v+94aEm7klI1DDbkH5UXGbli4GeC8T9fyC8ptuHI0QtJ4pMkn/8wq9SL3
QWPyFa8vyOK/CQ8TD3Cdqgj4sojTcAxelyipnXFVofQK/CJzdLM3yGZ2+/Fn9DPIp6ECXKkD73DU
vbBCeFy2fUUpw6JlkhgjEMqse7uT7+JKWPEfPXLWLFkQ2KKJMWTInjFhEh07TByYan+VGOinaT7I
rCilX6TOiPp5Sgx3Ou+IAvPeoGtBpcDgK+yu34a5itQzb9bv4yW/s9A5xDSEhWZjIWRjN2V8PfhP
weDvm6YQD122ye2KYNCdjO1SFavO42mq56JDSjrwL+of42ivLmccexmZ1TQpgqmbVi+gJvFWYSCm
bRzzJAD+XQWOxG0EkJrLO5dOuQBfp1k3SwY+qyOdvt8HAFkjOGgbp35zI7Afh0HZ4tuBNXyaij7D
82X7a1vRfQPjI/yFvHw9wo23PKLOSRbtXhNbSQA+HkqR7AkZWvy9lZgwZ/jkzb/WDZJFp5rBGs+6
0h+xV3nQ63HKInqGRKRBPfxyOVkQo9o+XSfhp871ViXUjn2J4/S51xXRvXaxzwXrU38l6jUhN/gQ
E+a5/YVHNRdedkentLzi0d47wgF8MXdN6DiLpcs886ZDqU+JZgBvArDh5wbXxl5kVilF0SFbIx3w
5kTQqNlxuv7R2V0lyTd39HOq9CQztoanIzbe7J/vShSolh4mCZoZ6KlmD5iwf2TA2QncK+Rcv03C
aS/CHrrhOyUV6vYsfyxTsmGkAgIoeSOTelX8elKe/Sj/7QwkTke+1b8dmISRT/nszM67ykWU9f4V
yf38CwN9YDuQMI0YV4I0w56apceq0/kMvCTPiAkyncW4FPCwSyLNCTxpyKmXXiTv/0Z2ZgvgAQHe
ohVzkWvd4KPIEw5IFyKcTqO6X5AJb6nchKH2TOr8z943UU4lDj8CveJ+mtLuqBboy2OX+r1Vloxy
Aoe7tsB2FH6Tr2gqOGur8MY3izAhCqGmUCJM8FLppcZN+8QzBg8zOAEZ+ovKpGjBalPyofwOw3oY
0bg8F63PInft6OCr2QE+TOS8G6AKpNjLz4m5hc24Lf79YYq/ODbAe/sciWwg22ZFgnvq5mOi9+rm
F9tkb9Gjb3cKKQCawlkVl3Sv9xSdx/aIDDNuVuNbVMs7e21A9LNMUL83JILUXseybB0SYlmUkVM/
CxFNek5WPyh9s2Zo1zrQF8Zi72gYIBdmNfYV0vHLa/bIDxjILCCJPloYkz05JbTTBcIRwUiKiz2q
ts7HjPXigQ41+veu8pjW8gGT8x0u5/W6EQ6wTBO7V59GRtuvsCnHwV4HVf+mhNvIk/OnxzwcvQrp
yJUIhWSRCQG4n3SCYRUtwBcC+03gzynisQKGvlUSGl1HhxowmDN1H4nrk40f8jqZCc0/uIarwbjm
rwlgv4pfmLQsCJotgiSFpycsMWCmHHob89+J5lPr6YvfQDvYFVA8tSB/dKiq2MtPKiRwxDPB4NP1
wp+2rBKN5MppDP5/Je42jYVsrAnzwqF/wog6Xbmh+H6GUUDC5bXAVRBXwJMkKUejX2MGYZP4hk83
YGN0xqQTU+e6W/6jraZfHzHuJTBGXjHcIwbZ8FhpYhHWDxpM5VCn4l7+OVRRu+eLmbssf9ZsPOLT
51a1W76jMsMEWX/rHhJ8FyNH41LHMasp2jsfHdAk9x6Z2aH3G09TegJCwLhPhrRqLGwJw3lLqPq+
261rpqu8r8w90C1lvPywGOY4yQDVDY5q+QyLcPHx6SO8l1cCpdoMO+s7v7jTmC+xVjbO2gLj12AJ
DtZT1GD9AjEYEQvwPONDrY9qRtQUOuB2QGDMoAYcdoXSaB+FUsmHYrKAhGh5nxourtbyyd+yK1Ob
s0xqV+J2wZY3SZAiXIpCfuJvcb5K15cNDt0XMne/Q6fvD125vVD9BfNxHgo7SUZ7wX0itudi0Q2E
i+7OF/KpTsDqjMpf1aZmBm3Ws2RY6GlKiBqijcHVqo0nhWvBg1YTe3dQtNYCveNouvJ5LgL3J3ak
zZa9/qDsL/vYD1jHq8aF/DuXRArcXOkebnwQ8xvOUit5Vq+Ppw0J30AZAsBVk3kIIbiidd9pBoJj
6JMjO5qAy6G7i03AFPeb/o2O29n1H/KdixS08zpbSrxR5GDypkVNxuf0zFq8jkkOq18lJ95v6lgq
JLJc4rjC26KKuld2ei5TxY+wfn8AbC1IT/SIKYyl01CuQJ2i9xwY4+AUcEnt23Pjcx51/STUWAhZ
C8p2xyeiGN5qtGsNIWiE8ZhSdrjFaec9C3iv9X3nPCsqTVble+ruboAfoEcQP/FlG+RDiBvnxbJY
rDDE1yiI6dRIDgCE5Cw1dkVm8ffM8w8Rh92xML2tvH1bupWDFGkRlxLG1nCHCwg90CbMm2kSgJhM
mgrxgGx7WqCzGmhGtelkI8L3Ysju6v4UgvRSdA4qJQMVVvkXj2Dw2AgOSUaYJsywQDlv5W5XfRX+
EQo9nKcfoDsXoYJ7Ln/hEi/Nzz3BKkr8/peYDMKfLxFuoE9hBPH/Vcf10Ms7hE4TOpJ3nfpxPvVK
5RwUQtjsLVIAhe/ELMiWQijW2RX6twFVybuMf63wY0r3xviRABq96stbbzBjnu1fXV9I5FPx/AXw
yqY7eG1/Qk6tym/em/iNmwkSmxc3ivv93Z8gMjrnsNc+CjS0p8I6y28zgz4Z8xxhAhh5rpd4Qdga
uvi2AncX2ug3Kno+oY3NJNXlBy7/bZVFC13ODL/Ob7wXGd2YgAqH7YrSWMdBMcqsemDRHwLicP5m
HVvcHlLYsxy6DCDcWk/zF0LXP0E0paoeChXqUy8r8rt28mc5hDyPu0Aqz8QJNcgkQeFJV3qG1xyK
Ce0gfgUG7mUM4I+V1WJKlJu5TvmJrIi/lVpmaKKih0DUyPDfm0w1n6183lesDw4ZrGPycAhNP+8x
2tE3hwYS9FGGyYss7MsduUJvI/B4d4f8/3xHk75+pu82nBmkddbTfWQ17uTDhhAj4WI/ZHeABGb7
hW+YDWEIS1mb4LYSmbVfebzE5WJ+yqw6JfCnDqEw1o7wK1pbRIfSgIWp7Q8I2j6mzoDUIVQdLO7x
uc+8HeZ8G9opcZXCeSA7nejVgdNxdDmFQXjaGq3clc30Vtu/XPAtiFJF56Rz+l0B2d1dDo1zQWQ4
ZMY5MU1nr4xOPnikR9REohDI6nIZgUVaZDy8BpDoCBjxFOcktQtvxdtdOwCAPH9z5Dn+diCGfJab
7uLwptd7XqGWuPmXBqh9a/7Rei039Jz0XaiMtOrCt/lYNa0X9xliLx5LZ3UpQQX1d2hvcKB1FHn1
2ZvAxejnb1StbFh2AnPWyQksqPmr1r2V868Rci0dupY66sdBpdu0uqgAAZBqJ6WgapTiuHdSFDXS
2aE+YXhOncoXajQ/gSVpuUTtRxHrVR1CKAMd93cCQR7In0jFTIFSM505ix95zAE43l0PbeofXkjU
l6b4sMpJ2YqlINQAS9I4Lj46Qk3EKLzqG/SAHW8lokpjfgnXdKl/4L1r+tkxUq7xXYgQQj6nySu/
Olu8vLcC9dPh1YB93ySH8hW4GXdrPRgiUWxvvOjyAXGnOaEkDMFOcNYLyXkuxNtDCX8wz3433v04
7eDvU+H/QjYREjBoex2GOlthGgxz31E9Jv3Trt/8Quhpy5r9u7zpZx2OaV9ZqjKOCNW41b+7HHLX
wqP3d6aPjLiWn3G28SVwihj4nzv+V4U4SGsscL6JBh0KUGvkW0Yd7VG9uvjLUxEYwJkbh15/pC9p
DGEPAq76aBS84Q6yklofZeNXBdAcPfVfgbmCFWy9t1dLr5Wu/pOVKS8qq2dw7OYkUQcyJIDNkMSo
XprjIITSZPJ3HFgY8OomwVG9h55WH4FcqKCWJBNzyop8V+sRt5lb5b80q9Pi3oCrbRsYKorBewhl
ZeVhCgNK1l49oF7bN0n4xisr70+3xMUVdj3ZywNXhs/GJH50F2TZm5A4UoH+siGUAbTcx5DQB+zw
nfyuFo5lwlJaQhQTgIF5lrAq+dESPL3nIAMeCuU9qFnyH1tuJW3asxCRr9RWv5osRvC8wr/VRsEz
SicgVl6eTbOy9XUVWg3EUwAa6JuGAJEHGctlX+rf9ATrUiAs7eb93Mjc4gPGGDaqcLeLs6pRFtTm
vhMoxDU7o4eX4kSe3jwxZUJsi5l1nknDbAXSmZgiQMUB/OgR6iglYDo6rsy4Rh7/e3Y6Fyj8bOfv
wbgGkUc7p6B88d/eRrX9cVLYv53Q6ABLn72Q67cJ2IG7P5ixNEqoSd/i5uBYrvIYAy1JPBAVhMWh
d2ocrFwE/zziYwHPIi3xO/hSnKq5GQc+6bIn/yNwhbOxIkB4q/k/d+cTI/OKL3dPTaeEPICeT2FU
pBoKQeOPVo3Ji6qwLgGElm/jGECFf2mHKAqdnX7RjCNNlJqzeUC8od+xiZAlBDu7eqEujrLjIkat
75iBpMzLluh/vT2pNDz7ygpzUlA6Pmo/YPnWtzCMPq6ekYQzJYAHdHIXEOVkyCK1Qr/I4DxYKzAX
L9mG6H+UsnnVZtOGFxGGRROAq9lRynaD7AiA2AWIaixDPdw9aeBegUcqYHWwHzEj+vBq1VUReOyK
MLY4Ah48j7vnEzeETxEEid0SfNr2bifVvV4rxVtEys8OqGnYNTP0mpyRAycID8pIHUWADGa7mK1T
Et9DAokHFtN5JQCdi75zNGbipvUTgnL6TGFtwLAE6qDtWHIKHuFj27MDVKxmfD6Ia7j2QPL3/hSd
uZBx07D/o+L9C5oZD1z7hGj6C0zyANHt63c90b37BqezwhcYk8x7sZYKJSMuBy0GmFdPXqAEHi2s
jNd/10wey1nlhyaaRd8HHVDTdfNerWObn8t1CM8At+3YMC3KJjUUjpNeZrPuIUJDD8LP/nGaR1e6
MTAv+em+uoQdgjfTWVL8DuMHoS1zqE9XAhg+JF+sAY/QzQdwr8gD2pzOdbU3RXAtnjtz5jQPcmEd
o4h4c/svWK0ix8k3YvkIYRupfjUXOjj5u1oLqdcOgQMPzLn0KuNEVu+aaye9F+jeU9oVhgO+Xr4h
hKjT/ZNlVuS7VgohgUuHKCiobfeQfHd8v9rU4vJgsXcS0xUTyqI1Z/j+PCaHgmg5CU2TChk7BsPM
SqEVtXeQlbBX6YTI+3tfrt6rWmvlEL8Ny9kCuoHwFho6WWJm0mKcGrcBUaVZ7tui7WkPETl43696
vPgbhY8wdbqhx0QtBrqX5JUaRb3AzIc2UbILYlkHDzu/r2La8sgFtMWuTFzj2hvLneRYPL0Bgwk7
FMqHCWjQN4gbDHW0VNWS46Jp1CgLNVC/9VhLTQHrMS2iX5vZWMWPGl5wnMiKga/JPB9jpCB8CagE
ewF0LoazSsYelzF4rUm3k4f6TgTQLcSD0jH2mt+8aNB2jEvNSTtQXReaY66NSEPKsOCsnolz5OJL
WcstYjwewGGdbg6xNuOaaT9Bfz5e7+gOAkpMFU+gBENiFeAQySqgGQMOyienQFpDSUELpftdVqpw
rZVSF1/m5o/QWkzLcCC7Q7lPoJiTcIElwFCVlCQOqEn3WO1hkm9enRwadkGteWVIQgu4MJPMlUAe
ve9GXhmSuOpZiXrYkxodUX0owN5RXkBzQJ6yMUywokgqB0tCOXJnttAUuah9kkXnMA9kwP0BlEwr
b6EoUE7ceuFDH45fcUrhJF3mHr5BZ3HSsdbldoBjR5/nkI6Kt5+cbPKpJFPnarVyHHJQMvjZkqdq
5VJtywkhc7kkwPvkgS10uaDiPxELI1exRIffE9/OWvK4or9jTO8Xhxg2nKm8ffSP5PQkTSL/3El6
V6gDUjkx2wQdkZZyNEcme8XGq35spEnoj6CtApgR0XWNkDILUrDhG0IBbhMoslmWbyRlqP24LHqB
BxCPXm1nguqXahAMTaVeD5ai1SuA46Idm7lTSU1be1CYhLG4lbdWpWOezet5UQ4GrziKbBLnzhE4
boKQ6DhmCERi4c1ehDR7MzYfrzJotNf0dTdGrzbGHRMkhCDPsfM089lyKCAYv19HsZKEc+L2gpzc
gE4UHHK/bsz+3HIws7K8NUs10iqw8JSc5wxwXRYKpnmD4yUn4Ji4kLAuhAigrKWMzgmvrVmj7B58
aM/1uEMJLF+JooMnakk91subJDSu1mzt9tANlFi4rKtATsHlFRvgjwcNL4fxB/6A16z5RxTQM+/I
VyCrIdlrzPzXqZuu3SRxORAul/qzPcScmI4FJN9fHGM733Uk+I9xcIkW9YkGY+jGZkMRWsVKfyfj
u3bfO/RSco7qKmkzqtlwf/cPGTVPKoFMLOhJ12JULJUoBYT4WGZ1QSAB0vJ6D4fylQp/qtH2RKdL
wb7Kt+2wAgfe28KcT1XOnIXkTJFK7CQ/1h3TOtC5unbI3nKvAOq3EqHso9e2uB2+G3wO+vPVKgiM
ub3kB9bWbbvh3bQEEJeO4HqTifx2FNCgKxnc8y0HnDSsVMZATbmRq1T3vNavbzQhSJl/mCD4tVXz
jbuz5BW6QNVNYc7TwXsQjjZQo3qSyfeJcjoYMl6rj3Uzcj31V4ZbXFvZlh4DCrXXxruzkA9rNnvj
Wqn5yOWHPQgpvF2m75iXR8o8vnGoMMslu1Ntus61UbFjyJSF2J42X/mDyBNmwsydoQDFzlXaYG1R
EE5xQ7xde9daqjcoJwlTv7xoxlL05F+TdAhVTkPWTqZ2CgGjoYj3bW5Y96/iKdin12PMN/sDf4Gn
5r0pW43iOHBzFSS5bDt/SDLLCjq/Rz2xpSxq2BfM+MfrwcN44dTOcvyzWkAPNR896rsfvGLjU4gZ
fkJP+YXvvLz0QPfdYC4YzHrCgOHptJKKb/7iuxljOdZ42xK3XD3Ek7zhvPY85EuzbmvgzEuziCAN
BR74RQrODIzuwyHHh2COTQEJdfBRRikoVnrvlUTS9ez7VFjS/Z4Y3r+IYvPnWMC1xc5bp/A3lEeI
XJrnkrg/OgjwQK3g4BuvncVxflgjk11RKeY1STHHIsISv56uqwwMzTuohhh3sgF7CF2fNLVrRo3L
y0kXLPNYhslxIAGvqllmTfY1U7MXAvNQrVeHzxSRYzE72I+ScbudUr77D+oBy4IS2NQ64HD27GWE
teTTAcQCCoRIeUAi/n6Ebpx2VdYQaQiB8m/Lj2xA03UOonxEZfwx6f4VL51GhixrcXRSZ+MW26Ty
quh8X0b75mpGEahrofhB4JJMw6on+zAP8N1uD/X6qIBThXmqtHgIabRF0ayD46xm+KAk16FEaIOi
5MW+8CvIDFtcFcyVghEHAsfOTJBAonEEgX7XtwNTTX/WkfB+4b14gxn1Yf+Xb856CUooxzw1lkKG
B1mlCVhCLlUUJ6eL1sLL8KqY+DanuDeciPgsrtgcXIXu0eDxTuMvmILI70zSASUPBKv5HAjxYgwg
9au/Ke5QSGwILuzD9qxiI4mZ94/YR5JfFCf3eI0cnqMfWS+Jk2UHATc1iNzfiOYyJ8aIbFYSu2/x
hbrB4sEQiQGiC45z05c/C+LuiJ0ZtIVJmk33HIW8zh0h7+gpyGTdKV8Tx/hRs+X9mbV1lAq/38HR
Cjhgs1k88BGG7N9Y8v/sTOvBFbS3EUnKSPmfrocpKTLmfAX2Uvp/ONlt67IybyNHNxYXCgj3VGuK
Z2aoWkhhO6UFIpvEEl+C1YqzdcOPUm3nah/5gb3axrRdx9Ucw2ULiVZir/Sx9PgYPh6oCX+u+wkq
A+8cu/w8HthIygKz/ZZUmW+VtZuhQ7suK8zLxZiR9QBUGcehcWEuLLF6fPJ42ac6JVL/sDj5cj2k
OhJr14MTDae+myL410vDUbSGMPTzuNUfdBC93c1rY8mwMM8ofYe7bm6bJxY2eKInYtifihPuabfY
BGyKZmZjjDJVAfMgXW/xFh+/ogPFK2OIDU2Qq2gSEZTLumBs6Xqd5N/m9jNDakzGUK82PZykf2Je
p5h55h8GDq+VYy4WUn9FzM+c0j/S14M2eqK6ZoYY0c8XZtaRiteKWSt7m6q5HueWzdB8VoxqF+TU
qowgJtqi6eaEsWYn3pD8bpp++eAeufbpCqPO8bnUfVZ8Y56aiyvOAi09UE3xv9v/JWIbOHzOuFFP
Cf2px0zkZ0C93b0xHLYePsDnnZY+xI9xehlRq2n6ayxYdy7jtKmasIK4fOsgD749k3mjJvFsntgU
4d1kiQ55pELPA5OoVbh+sNX1dSD1dW+La7yVtbeUYZla1fWeOQ4aY7Vfc1Kib1qQ/cXiboZOEDue
SePgitRMZDRa9kkAY8nwMRL+3Vh2ooZaRo7y/jo1/Nlf76qgz/s47g1Zw5ZLSSafrVVr8WY3nZ03
oU+7X3BUb4S6RsnE/naIUz5uITFu+6bWWWQT5CTnMeJnIohNrhlRG4OtRPConO7mv+Zz9mnoJnek
d/ArGax1eU5XbGD5N8N5rVpVVEhSKYuw8uSrkKXCRj7HmoouVf1Pk2RnTAo5+eTuvCe7yEmwKUNv
qrG6qD5asVgO7fqwpHuRCglTEwf86uCKGRp+ZK9j1B0YInSRCysGzJQR6ZSD23bR2IzpVlIkLF22
ePB6zA9RKF7XkcakM2O7B5kAFlYUsxiz5iQHupm8KQgn27ista+f/Wmlf7P8uhMC3OB7wxWj/TxB
NaPRZ/oP/Z8hrZHei2J1Bm8kz6ynKqI16IYUpJEs8Zt6+gj4+7h803wbnhT7hJN3y5Ulsg9kGgSN
2uVEBhSTpicrAsEmppyUVmfb5Cc9D2sH9DQ6L/hzQz5jEBLnex6VzaPzDKbVYDoafKHV+Mvoh/TX
ohAXxaXm7Ne1pwK2+gnapjndvb0IobXsr0ydjaUKDSjt/bcoVwB214vfeV3zpuzhZGEiSXOviS7i
ufDGU33OtVtc5a3xM/MXATlxtzDhINfn9e9aO3mYrATAZoWp9N0LjDAWspuN9i0PC1qtkUj1lVJK
/x9UlWg8FMtE2H+RxlrKWn9GmXTTI5SFsWu3V49TnzTI88azO6cFmVGCQsycfCRWcyYrmLI8F5gt
jb0UJSj3lbksrzVOKGxzvQL7IeM+3Le0GZb9ONsKrDeBLnlU7uEpSIfKtsnHvpitDD3SXou8YSCe
QXRrVDGSx/3vqCa2sruQvT21/iA0tXlDe9cvK8MvrJic7P+viJHTaTL6jrF0B33TYBOb39x94bf8
FI39mDm76We795/UJ73NEC4vKdnghWZli0IP0S8JGGXMCZAgHtHRNPEG0UisRHbEmFerD6rqiprV
opsMTi6gBBFgH+P6iQ3SW9BnR7wmSYCRUHWerLfg4xwL+27o2D7Yxdt5C/Seu0r3hrzfF9LMhUCc
ya4O+FbwHb3Jf0hl9QWgQ9wAq9xkOOHx7NeXxjn9oXieTwjX3Q3jkNfXzMEtyGqQw5QKOoUZXqfV
0lC640yKmT7j4UxREpo6vSFLW0J7An4KKPhRoyTvb/nGomS3VMwR31WrVGfsUISjkTKreCs58dYK
lEFXWZzrxyf5Zf9VkcOrwN6FQX39JJeZSk9My5PWvcdRlunt2xakxihS0ai49Z0EffqK+2PgCv1d
jv/XT3BMMZkINewTz1UskzcRyQFJ+0PgxnR/o1D43GbarRteGn/E0rBlTMB6S8Kq6dTiV+iIMwez
9iBIwtpv60RIkwWzznkgI+yuN2wqpokv0+Nv4xKLV8q+Rf5n7PdSR40uPolw6VrKvY5tLTf8MheR
C4SEgKXVQ+aHmyvrSmblGMNnPbgY+tVm1lL0adn/ZECV0+FRLWxy/ukI8sDq/O/MbrNZ8iBNHmyJ
u4rff0PcmubXlqHPMM2skR7/9QTsmC5uPbrbTyP6AyM3QYXJCwyOwohaBBIGADvLF5gjM0dBgZ/0
/j2mBGMamidkpwFcKdgFZ3Y3ou37hEJ3a4YN0GC1ALasVWKT4DwrwKph7BbICdj/fkQLx3Sn/8zU
fnmvFsyK7tmPHNu+r1LTTO0EmdGhORRU/BRhIGcVEymFnAkgvYfqlD/u0SjBGmFZ5gM+ZsiejUf/
pkPVW5g6oQ+B3FyUjc0J0G+WX91aGNrH2KXZ8VQM+lx1+8yjj7g4GmJOwOW3EsqaG9OSAMBsNm5Q
hFDIAQ9yabQXiAk8G6Yt8gO1zEZgdb7g0vOIO6HaemO8otyi5ofG7IQTupRU7H+ikplNDUNMY1cV
/zFmsjg+k8m3t4DqEqTLVZLWGGpOqyr0v0Q5dIPqLI8nJBq77ZBADKv57qr8tUKpes0OQrL95O/d
I27SVCJ/3FD7xSjvPqGgkGYpufixwIu3nEjKxD/XRxIgq/ZzPI4KDsaJO900iO7hwP6j8tZRVKVN
nrta2dGE7yAIZx99+xKPd4tBJppfXjQzFo8av8Q6WdbUV4/uh9Hus3jVHXzLPcklqSci7GwTPyVs
lDzsnYq7dmgnLhqjd36qqtbn067n+i01DGP0J1o6UW0UZIJYPdokWSQZ2SQwq5wbCZvm72S7fuWk
aTPd5d5revNJhwZllNblqLHkItmNum9KeJkjwwuTgt0pTBR04SKtrveDEVqRf+yFx5YaRtLVBc06
cUhvPLNfDV/DErpC/VDkRtUZh4XYHeDsI2MWKTdUhqaVETdr4hWvbLmQHlVaMTD+Hmb9Qx0rk/JP
yP23mCmr3RS5xpua7ErLEcZm9PSlbQloyxDu5sgnz6iUYH4ypRI3XY8aSW+8inAsH1J49+LIUH/X
rvm+jHYADOmrFKXIUum2A95jl/DyxAfD6pOrpW4j8+Do/U+L7ZdQ+75AO9FTST70KewDvKtjpqRR
+KJYM/s0mN4CNHTRcK4bK2jg2hr/uZkhzujTzIHMC5/qEcXthTj7ZZfmQBrknNSgzIfYNFXSE6Dp
D9zWyUIXHQuaLYAc5B7hlP/nkKCaTROHM04Cei4dFxGSY5Xzl3oFZ6yurlnhIqjMQjZWhqLE5M76
84d4nnM5TiN+sbrYx4pUrf7snautEr4xL2cSbyIOputHpn3HjuAl/AmvndAU5yC8AxopwX1J28h/
iv6bl23ip1dEJTZCeKaoL5TrGrNNEAMOQyZpEJHUiWacCoqeDavprGKeAEdw595IETSzXBJS/Cor
/ssXHKqgsSqWe1I8Atb4M1brayW7QkcXVyrik6LWZNCnX413aTRW9XBJp5Z7ZgY1kAWKAcaYrJ+/
5FY7z7qZzmAXVjveS3R+fWP09C6OSFU7oeA9KtIEsjQyNRjC0ce1btpplS8wEr0vlWOlllkKGqGY
el/PEfjCfccPFgX/qZxRGBiAXy2//X6KciOrle49zHqlZFrJ1IdYWmPDDYJIvv0HHM1+XeBNOdKS
ky/mu7HEJ11lQzQr+MipHYcIzvlPFAYbdFhC+kYbr+jZiSioZM/5cZMB/77JNgbfh9bb5F2cazd1
5/1nIyQ4690XLS4ir/S6AYs6ygfq8XmodbMh9NlD/XX/NIpSU1taV4pu5dDqd67ixPDJp8ebjK9W
FqWHVQVwiTKdI9bs3wtC7Sl43+w7oZwI43OgJ+Fgar5Ul3AYP3PX/bjzxVRe22hbAoXPRMSmcjzg
hqy9DGS4Q+Gh35T3gKNtiI/VPwYWLyzVdxsGqnQf+4ElqRK1nXdbOi+hZklAV9vWeYhdwl3eUdc3
UE7M4prNt7ts2J8y4gGU+skH0r2hsDTAPQWL1434JYc6WrFBSRXQj4ri1Zyjvg2ZsgZJSGqVK4bO
AL3KScgckkIZ8d7s7mWjoW5m9S24ZXXscJYWqRyP1idOb4o2XrCAgkcuQuirie93wPRIgnS4LNaD
7PuMtO1+smgrUkZK0i7z5LjoUMAOa950zOgiVezYmYmeYRfMDEP9t/K+UKt7jl2FFr1A0JYZpWsk
+HCIC4HXQ1NqQYMp+ZXQ+3CwAVQDtEAYW6rMfPn+y/AzJdzZfGxaCLVvhHyKnJYC4gGawrzZjFwl
VDklzbzQHhYbb9dWb3QKEGWJIQEydqop1wnUdb6xDn6uxXa11Xhliu4PORVVEAwGX4IbIsS8/gRb
y6oHd6Mr1xkQrzxaA/PEo7bbdoIWmBU1WBc2C26paCBqv2nPuExY5vQIzvvhdFid0QF2WzLQZKzo
tU/dX9w41bMuRTVzGCkULRI7LsK0t6lL7ldU8Fk4tyveWiiHzjwarDJUeUwBHaBMEZFJ4868jz1P
1ir9zt07sV+BqiaW8z41H1vOmu9tlC8c+hG5euMcRktPx9R03WrS2TETM/suZlxaBnAxTDqHmplh
K4UWk0rfZrlEmB3MIjzRwH3n9+h244ywsSV4WeKb+QA4Zzj6HTPEaadEvP7jjn1v2fHEP/Vf91nj
18bdygh9RqRzYZhVIl12cdw4fN23e5B4rBTIBG0q0mhwkmY7gOhSzi/BLQbnLYFKCDYNogRGcqN1
HN8jVVVZ1dInwVsv1bQ2uyFgzhZYVpHoTgiVE97Clf8UQEHJv6A9ioGdREpVcnIA7kZPNPrpoWvM
NnrcV3sPIGliGpI2Cj46So9atBRpH6aCJVJozi5L3y2pU2QnoSwrC9zvqg3AeX++jAzYqGOZoGeE
si9iPfdSa8QM18w0qxavlo24txGpevMeGL1VI8LNBY8y2kmBTGvcTCzF1e614vLfwigzv+hxfdNn
C/ANeUMx0a2rxfTKBkBwwiDl6m8Ke4u8vBoHPFhgUFvG/3V5X4e0nu9m1MeVlYRKjZ4O8Nh4lMcH
lXi8Wnvk1mRiCPq0rpAt7Wq2/COHJvuIiiX00ghv3ieMsfo4hH8YFEEvPKz060idVZJRcMmc0boX
aBWJ5FLuyMVxElCnsj4rp56gd4Nx5R5kfturDTJ3l94o2mjOJSvcl5J78ij6rT7eE+xUHowrtKt2
eSD3pc/sh7r5Rkoc50g4z2Vw67Lh7dwoG5GCQDg9BBC7zfEwOrSgAekelJ+SWTRPz6SlWX8KW2wB
0FDRqAhoYlPY6qqp8mJAjJnI6OheE5IuvyYssNq6v5QG1kUWug5mNuolTTsbd3xRy6dgBpxay7ww
nPqSU5TfcMKPjlTobiukDcR+xwo2LQke49NF0T1X0biE0w6K2VVYLFmzA+H4Y4DcGBlyDendy6bb
Q6hl4/szWTROu4HXmsKSbI569NylRQ/holjB1k5w8LNVZEuczAQ1Mmc/pm0V4ruPDpcqU9lqy32w
tOab8OyyVTV3wo+BR758BeATFYRB7dzDuznnMtvur5X82FHs6RkP8HtzuyxW1DYtV8W+equfY8By
F6+uDjxAPLZZIhSno012IbumLJ9ZUcK7ANf7VlmpFVSdcVzlh/yFkuwU+jeZzrT6x7IXomj4iShG
Iq5x8zbAe2hh6NOiD9BoRXiCy7/PtDbq+Fi+C3UktseXioHgY13Sm4VeXZevi51rHUx+KNseLUQz
vvxN66qmT0Ff6pzRzOktGgrX9AbjuElYk/WGd11mNzN4CWduaNC/Akzq0ls5P6Zi4os2nVq/Pokp
EDIUNh72r9qQBz/1NmQ1Rrzx7qZIe+bAI/LwV2TR3zNsrOYyoiIHHRXojzfpSzAdafb8apeMnqhd
TlG21YoQiqo/iiWbhPYb5vxdhUa+ykn1T272x+6Mz+gjMedMmHGU79VF00anwq2CPbXgPtLe4AxP
Qw3LvmDUXTg9nnpuIclycQVEX4YKdZq+cuqYSj1yALyxx6DISOIpYiWkdnFMUnd14AdN9SsZOxlL
mTytaK/5Bzgb015U3EBg3lXcgrmuofjr4P8jRMcLOGFuASHEpX3pXzmbQBWXXvICYQ43wSoM9F9Z
bf4kXynA3Qs+OeiCHkQJ8zO+MpGdUk9s5J1sxD+6VGe573p38LC1ObaI7OB7Sg02L+l3aIo+QBkD
zTGoUYlUGKkh7FzkhWPurhm7Rk9el+ZvcL1BIQo0HqBQCB2AwZHyiwt7cw+ZIB/hieuEBWCT9X4Y
9tOot6zMkWI2nA49LudS3wTBeOZToKOVRK+rMaXxk7qUQRpzdfg1IEzcjdY9Iw5C+Sl2/pjAoH7w
cs/H9i8pdnKZ4VwsTRUo/kugqySAaZpTbOfYjjIhBFWnrG3gGF4DBhGge05+riw9UN0vQqyFsThR
NC80e1NFZOZMNpuPbqMnn2UlAvNTkcvrDJJc/BdtqhjFZ2su2TYj/7/xEGoZjn7SIGwYIAbPUsCP
VVkI9dgS6XEBmF4WFpLEhTJ9/qz0Kmcc6tvFFoEk5qJgLAUMIGJ1i1dwYDqKfmXs10QClSmWhIsn
xBwQIkS8CQxhPmmZBRK/0v2cdhkUn+qlg6vesLKlXUmwDkwuC0awlME42tnDdGBww7H2SYFPb4Js
VLU6JlKkasbGwXHuhWmyz/AxfnGSRdjuhOoU1KzeE2oIQP2v1bLh9BOW/Z2yYt1uablf+FkX/T1t
BwguwVXh7kq5ReHqSza402JVyKJMz9JWX1Oe73wgdPj2R622xUS+gA/RxwjKEeGw94nOV+5NSWd1
jQgJo0elI8TTtud3H6EwQ7713X+mIJqUlYKxxMlQ28JbeReM3drW34mMTXT+4akG6v8Y6atSV0s+
Q9KD1s2eEX9ktY7PeDCw8uU8VN3v2LUdcImjwo+n9TJHGG3jaMZd72V7bLriP48OOOlvcRB2KvO4
3UX0xUrd03ilyZ7LcPl0afLlXmOGNVu2xrjOGdcTiwbzLuVrRYVv5+0uti+plwcrglV192z97uOZ
PRarocvMiFPzwk+rHxyq3vMOQ0GbKAsLwdNsdTzNEkI3wUn9IozKOEekbtYqUOZemDO/jsR2zJwi
6OOUPl18gXLJDaeIIldqxDzfuTMY9nhvrCqgTFWaaOBTflLD59MYgRhXENZftICQrA8prS1PYn3a
szsIEAjwKl8si/+XqdHKmptScn0DPGOgHXwvHPoWRA//YongXR+f1dLeqAJdLXcld4s8pWKshPg6
gfRa5jhGLFTYMeCpCAlOOSWNmz1wKB82GRJ+7cubSqjM6IWjlJjg4+BRImpHfjY2ltr2wBoVE/Mt
492GL+bTVf3ilQizd3UFnnP2cnrLO0oqzTquLgnF2D2ehdDI4frfZz8UKzCfB0RzjT1P1gXgdFJC
2See+bkUtjr+QsG2cX4FIj54tPUp3yJNa74cUz4nYHQwKk4TQw148NjCSSph/dHt6L77JzIENzoQ
rEwhMC2UV9ckKaAACGI2h8Y/gvWhNVYdA7bkIxPEEKekugAFEq1c3Rqh4uq7AefkFTWiC7Z4D2UM
cWjymkOheTxoIGBgnLrF5Y255OJJwjROKMM9QepBPzjX2CDWD42qar65w9GNZ3OSU7jsaWucvCfj
uM/GBJ2gPqZhewI+3YnW3IfGNI5wViaF7zEZpECQKxLB101uiFI/6cKjpPJjUDM7h8fO5qM3tA3F
ZkMiq3GSbBGzxiHbyOJKObJsuWwKpmgNjIN+TGQX1lUqwpMyNjr8wBYSZtc50L7QdJfAArGJ0JMm
/cu+V4vX55H5jxasbeo2VyOItO4a/8Y98eDFZC7U7JOSLuJvVABRHk8XZTVctuSyTrbEM3JwBTmZ
SxwAIUKNrYtPRmASGnjKGCnZ7FqvVuNtBbtRQQerV6VS1KDK207LLES44V3qwAxRsgaupaq4q2Ev
DhiVHYzwDbVOH8abTLsbZxFm+TKL02g0KXVHfWzfUFdwc32CsuBTdPnoBbdpKt08Sl7c9fmkAyDp
CQHygpLwtFnJo7wa6HoLJM11h8CH7uvo8xmIsSMZdB14vjcCL3bmc/ZVoknUmZiEuW+8J+PtvtXK
OGAgo5HeZjBkG7kj2E8KUPfvcw/uCaphSHILxdIhleakaj+gFrMPsnYfKz25XZfgPQgRgyCNxDXY
XNJNnj4NlbBh+UDKfedZQkCjf2RIrphFRt038UnK7PTE4Gj4njY4BNr/1jhqnzeJSoTp2mOktZc/
70bA1U1nNu/1nn8A2lpwbPasEyp99rwrGKqTPDO4QF/+EJmqCV2kyufegePwRAUjmv9ctom9+HFf
vIJohZUNKSGzbpzC30T4UjSQo4u6LDU/91EIvUWpsu7Ld6rNlNwC2D7kO6F3bcJ4T+IWxUHqq0wU
wCP01kOU7wvt8MTUvazWk56DFd9xlelv1wz1Mp0hiGqh6hgdsy6vDTD9v1uFCHtv8tnFhtZA5exI
HveKP7YFBNlzAWX1Ro9svnIBgNNOKP6zcS6Gd336U8T+eJlYIrCXKGnq1u0wVZhPh28Vfz6/jf7O
MzOOtz4nx+4aCVeUFdDZB0muPH8Z/N362gpujyn6XDB9gJj7nKWUwJ4WqLcg8iTD4TR6w+m2wrkK
xZVoKgCK87tGU6hUHKD6+L1u1fy/lWEhIcad6RGCgxrgy9chL4cpFzcFLK8tZuxXM6z3xqUujHk8
8eYq8XmQCa2YIZdfDHD7oaEhKlw5TY+oCcm+oEUYRjjMkC8NMdM15NGr1CggdpHPPaJ1suug/3Z9
V3lPiccS1xPW8dY28nZgYqYDIN9ymyKwHY8N9JomsXWrLs6gIO8dGLCE26nf3TI36r52H5pkzUxZ
EUxy1w5NwJp5C4lNvT5vOA+vYqO6PMbm47bFV3FFGwN93gnrEOcckz6BhA2ALnE04Zk+dDWAlAH/
9QNON6Q00s6ZsutB+5u2Uud3gBlvI66u/a+ZAfPNvAPnED9czMFRD+GELZQOTe7+WHp1OYNyOXPh
5gAmbH5krjA/OaRT/42kCCq0M3tr+kjj2gX+TpjY3bbpt1yFaMO3dBwgX+toRBeK6fSBjKax5ZBX
xRH2QgMmC1wQ97LZ+uttNfxwYpyHhRGmJy+pdhWVKSMKSbwMs4S8nMG0qiWaJhmL8uygNaz5XlOq
TeZ7z0vfyt60odARrz8ODj+wzz6+UEXQkY6jcQMVj9PvYXIvwI2+5r3vDsoh8rsk4xqpFLW12sJm
CRp3JErSK8mgGNKdl85nq0Gl5+0bIgTA3oNdenVgj3BsOer78O0cw17egaNIZ5uYsIquReMDayI1
NI/K92KRVmVg+5PneALtsPmB2s67nuhy8ytW9Gjc8VaOQWWSjtWckoWyh8pxqqxNKCp0FWsymmfG
6k/41UhoOewecqyJ/zodic11kFI3o2DNgOOyLEMv/ijjreuhLKyGQ2hTMLnc/C1QzlETE3n7kQwC
3X4J9jqXUw3+cM5eA3y60HoLXmwnvM3Y2OKRxUxlkCZhpS8i12uY1xdRDwsLe3VK4ZeSuT9pMOtG
XjoHyv0OAHbrMbjQlshjd1Y9m1XByyeKaNP2Z09DULwVpWpq2B3FYdF/BAWX8OdrhpeuxP+1jfne
wEQv00Bs/qNzQlVc/eHn1Hn6qIHlCCWbm2i9IMDv32t3zksE/D8T6JjUcYOguIsGP+vp0dwxIjAe
IxD5hkkUm7S1iUSCf3rGcHiqSU2yONprEWWcHaYM4fSpe3/OyIkR8ltAd7wwJ01IFP4T1fRIkJgT
FnXjjb2cQjTgwOhRYHM6wPjOIjAoXRQSN5QWYgvC48rpJdJgOAWmaJHF9mrSD8ReOkJXh3rQq/GV
ika1GPIAg17SZcqIX1tat0tJdKdMyK92gDrFJgx8GtAT1IJn9sotmgyyTuGESj+xCPueOl5yZhfY
OkWeEY+3POIUh7U8qAHDXKxaE/qzLlnisrHVGArbVMSMfl3/WsQcqHCPY/MU5oJHlOzkgRpR53Lx
NetrF3kjmHzxvlDKUeOEoRQXyRyW/sSOITH4g7jQ8AdcjH4ts5XiasFqd4oemCXY2pNitPwy3WFe
ZBKQ4pGjKkUKRnO18+WTL01XA0FrfbyRXDqurqH4lgD60ak4EmynkGV0tRofoj/5tCdKqP0pTCbJ
7VkOetz+AyXACRsKvII8s7pYtAZNo2LZKv0cG25iKzY7iNuvi+v1ZPbsYHgjVdTEJmSOQT03E1Ga
pOySrYhF0lNDCvQxd0iKhrf1zzMmKVvTY2cKhOj+erqTLk9/8KYlve0e3m+jdd0Lya9l0yK9jAtm
p7hPQaXMNqZUaq1Z7jbompPsS8MGAdv0MLs0ePMm/jughKviKPt2qPEmN8W7WQhop9UynZuKZ11+
bAb6OXUB4eGg9Vw/8g2nPNfoy6FHp0jmhnz7dZ3SuASpgjJiOGDHQUU21Drh93xpojqHxbTYiJnz
At58cysJ3czlOldLBbefNVg81m/A5SZMpJXlAV4WFXFOSkJVlfZTcSwb0yvMZ3RoFt0W6pqTpqaH
sHuXwWJBLnVr6CUFJ1gGm7pJHNrc6sYATtMyEhGt1byU998A+iHXOEY/HuKT9lRnYzm2DxOp6p65
drIKASSMheMDJRNT7DMQtxW5eKMNGGk6DG+QL3r7S+Hoo6YeiAGF+yUhWj2ofHpnL/wL66JdXnuM
5hzX2AebCEX72u5H2gBDK2qEwUw9wJQM28WVsupyOno6fQYcGrNr7vDnWBXiFgGr6BU0THGBV6Zg
+c7DD1ndqtWRGB+hpkYg0E8IUCFSUJJVcwCnirkM98bjLvUYCdrQwoow8aBJBMx0RqgcC44pWEF4
XYBfDf3CYU03lhTMJ4Dc3AMpRekCOdsSQPCgWqpQh7eANSKDvHGpUPIHqgf1EOwJ9P55pE7MGAXc
4o7VA/CdEa2qt4/A4Phdy5x7z1U9GW0K0FAaePdOXtYEDHrC6plSeGWhc44MNd8g4BE6icY5rQ3e
P4DO2bWAEpFzYY2UupMxH2xWNS0stdsdkgaOrkcQNQch7lNYZ2MymbuXVW0KXp4hoIzjanxhffmA
5FvGtOqiMi1XS7lrmNpYdlaYGS22RB0qT5n/gUfMn3mXTdGou1dV2y1Da+xn3cXl6dZ5oviIixXu
MjB/0kThcgddSNoEREJ3lyJKr+h7Ro0jM5iL23C1SlfSx9RLVvV6nO5p1BYQTiXyUbars36j0aPa
xBXdev5H9uElQbaaULQZrURmZ7jRuEHNRx03lCmyfghfLJWpHNXekoH/96aF6a/Ve+c3KjijD5X4
mQm7RP/oAnGGTwrdzr61Z9tec49ElOikYCa9d144waZX5V+ej4a9wDSJQWMRwTdZIPC501A7EKvQ
bWkGbCz3OJOBQ7IgvXffGOSw+B7xkQaq2sD62FUwJbHiLFU1fWw0gBj53oo02kD76nPGJy4xQkBL
iP3oXdgplg2Q32g5ksmgyb40/FAnHwWOVbfSLp0SKiBdiW5Jq/zN2pzWX8C6Ti9R4vcBxiZKj23L
slk3tJBNnSpqufiIO+Hz62n8uNghgaRvv8KB4TSqpoX35ItLk9TfjSlB0SbfR+Alb53jtAzdCFxU
sAg16iLrNC8lIzAC4A3ixLRh+GOddI3UxusmNqT6Las6NF/vcWXssp7RgNEVvlhHCRIYHFgs8Xz2
DdwLRj9tPYZeDdwTtI/0HKbH//69nLw9aZATS5bFydrg8xXGaQZ4YbNvQHv8IJI4T8Y17qKUboUf
ny9s/qWWdydOrZodvNZpubZilY/swtuQ66n0alPfQ+4EZZ42Hnjj+UrJDzeazxlMXU5RfRcEkkSK
AvGuBsa1COvXhzE+aQXHmyhoh8g4rpXjceFUhe+gEHnOjKgUisnoCqUQBUhdXORMHeW/Fxegdbf9
+anvsYNapSBekoGlR3wqQN7PH17IdSrFN/Y4Cci19O/vnBmBNwTRj32oOcXT52RowgpWRTDkdkoL
qVLHXh5MBIoz8hL7yjZSNx4rPrQYOvl5PveKqjmkMHCsO4woxhz7ztUdoFrn+uWqMntXcEZUPBgO
sPU4dkWLsFpMOSYYPa60b1jGd2tXX9fdUBkq+qvZbRrWiO0W4USnWCzItaYKbnx+bnCZTsAI+CRz
D3CKMfomSxCSIVwKJOQyA8cfuDkgCQz5Vf4/wwE7M1jRpaqdHBpm9H5SEXrhoETrp0Urd9hIaeTZ
cINwEPDLMKLuSln877IVlAxToa6F01pUMeeLILLJ6u55iDHBEamAjRBjxcbYOkThfrG8N5V2QXuP
laMSgE6Ips3cLZvHHDOEoVn98z1XnnwEYg5TXuj8YiuNFEFpAKANi4mzhtweYxOCxGW7USy7/Uhw
mSRuTnNsO3EAXAKU/yi/8vfZAbGW0eHI9fjraPtoWgp4EMw741+qdjo+h/9oRMdU/ADLW/Zo2gxn
ASh4LT5NPwjBsuCtQPeK4TVI0YvUMkBUHizSbDXV8FH/IFl6ygTu0s2YgZ6izIlv6yyCn1UJpXBO
i4kkPpprqCtZYMokLGOPhhqBumKs/v/s9hkRNydYn8GexaSIR/cvzGehRmx5okApkuq7qlxnIjQU
c/TacQPvEWqa344yPdgtmzIhJjvNQctKDgd2jG2NY2ZiziJ4xILoxy7R6KbgXV/RLhDJ9C0UOGK+
/bevfeapZGQrSutXmwATAEhkmcX7/wNP7yqFFEVkul5Zr8LoPH2KdaxB+pQkgdWcN/8yRR4bNK3L
3OhZ70AoAlFV6rA2y82XL4K19F658S6vOZWB5RsajA71UfWIUBdM5RqFjARRnLCDHeFOlKjf6ZEl
nMH032oKc5oa77eEHYdKolgqSv9kYiPpYNBn0fcUIyJw//7Pr5wY0MS6raAY0UiWAhwScDOiBp0B
VNFzQRaD0Jl+vIrWi66qmtADOWJKw05heOBv52gicIITVnxWch7ubhzQURNZu0HVJ8xF7vSUy/0R
wDZsy//FxRTkxpeu30USko7Kno6svClTjk/gghxELE+XA3iYnRhERSLLfKQkpZukUB61v/4btrfQ
vW2yk/AHpDsFkGkOXLcxKGaZ/ptqM2IVXtFxUdQxVtXkoAt84SS3FEv48Gm4ZQI9W2u5N2Q0ezPt
8KZxfVA1QabagSfYXrlhwjAHsxJUltOrtgV+vSUBpzeKwZY94wYABDTOFT+8M+blGCp5j3YARyPH
J/sr+Srl0H231Q0zdw34SoX76R/LZ0td+sPMvdTuKpnP1Laafu+hy3NI07cLMhueRyN0rz+mRMv0
ZXEgx9ec583lzRZ54ErXj5ddHQpKXubkIXqUihxr60aFm+8xLFJN+gmw1y1qx9HoA5R0PPweFnP0
rKMUDOEGjUuDE7RsaThq2ppmZ254B4EHoqIhqdQOo0GgkkstGzqxPaEeRKxIi2QXcAGvuiQ1E3lm
EuKHHJQ7SGkxoedwmQdy9Fwf9eQR05O3IFDbeIQzVJ4TkALEiFRjtR+oshObFggrCDdqsi+p3eO1
VqCqCpZEp535l3BoFq4JVuxL5D6WiFlIhqTE6CKPQUV90ToA+0HpDKAg5x/8S1MYl20N4pStqOZS
jCNXcMLyfPJACGW4AnV3MT/DuOgQmRAnrl52ChoLuwS/8FeYwsKhkydyHBRPB6Qz7wV824AtFfXd
UccoYhn/QDXEGhsYtXkGfavhcPxdX1t028z8I7pxGQFygWfDRrLDqybB+skZnSP6PgGL/mL0g0NC
mxFdLbojtGlkFZRXCWvdq4iV2Wtjvl+Aj/FZWtk5IbaFZ7e8fkRfJkwzYxuoWl6X6qHKO0CRfQbq
3MttIU77XjDaL5PqBncpQltb0DemaSdf8BpqyEdKULyXTvB/HZQpdG+8tKUe2mOpzwMrh7EhIdvZ
O0FqIx4QeMiuLcHoTrXRv+9LYTK4lkOawAscJcHtocIYXSC9J6ye4dCI9jAn7YHFr9L8Kp7+NFrq
KZaQp/fe5Aj6tyDxwGqD0wTY+/7fGRt4l5ajvR8t29z7Xyt+7r65ZF3Pz9gHH+1Gl3Pg5+RwT3Tl
B98hxkcdI5B0YiHIxGQGf66lplrqN7t9I7OY8IrqQCefCIQx2D3vQ2J+wvVhX5erd4u3VhD/sX3d
V1hvcr8ca/QtCmZKxNzkhJVBGV/lyI+8euio1KtHujciKaZwQ4NlKmkaYgg+GQYIRN+p7F9hZd6V
TPxI1/jCw2K5iYIyW466KoIr2kj8QB9XsxqXL0BNH0PVSm522CWCdXzybbrrxNvqhLe4UCcMl9RM
HKh+muIum+/1dRY37wcw5TdbgGAZA8Znmq2rpYc4KhsDJM8YCYNLSi+9VZOQQb+MYtEbpEIpiOJj
Ys+XPECsDQNxAAkJAR+1wDMnAawJ/LiG7x7V+0sv4Wi0yMLLTV26FB5ypreweLY8a7mtd6014FHy
YSIg3yj2t/aqVQGBuHDmDnOPmcX+tFwV+7DgKX7y+H4gZldkXlLijt7CG6kq1fCiZKguTX4hcmB+
luKyTX9PiqEovKYuE8+2YkDA3ZKmTTQQ9h19VeSQYynMu1Olga/dDbjS35fffulCn1VfCheDfEch
W/9zCbzQTyZPf27Pq1ev+b7XUR2cWdEfRj9w87sa7qOPL31pFVkHL1dB/l5I8/kgt3DuLaJImqzh
3H2ehroUhzuFoU4komblB9tsCk/4eL0pRoGSTZPUzG37dsYJl0r9j68qCTp8Dj6Dv226yUM+cBBj
GnQOKskFyNmUBk1B7xseanAZAQBhELbWjtBaFnkqLB/8mF3PQfQOffVnh2wI+AY041wT2b3sFnDm
/ilZIkbI/aYlqeZqEPJx6j4DoKASxf/C36R38whSuwgk2wPWkS3xypKYAvVhNbjcdWYRc57AnCU3
Pd1I4BqJwWu4mdH/h6QmAGl66eyj9Ls5oj0RoLlq/l2cNuG+ErOjc3QB8nv9AbT5y7eeU1CLalw+
jj+YcjJvjU/5Xwy65fwMVolL7gpEDtMxt0u0awPZ5MdYhTa1AMa8xTRBznV56ajljN1ehcIPHqMA
KDb+lJ/ZuyVXQkRfL/Fgk9GN+yJRzWndtjmKHzguyyR0gz/Ld0MUzOzczHJHXw/lj/oeZY9KVp/t
TmYnCFgBuqMRr8iAcbEKcPOSzj46nHKzY/IjYGDYVzGMwRRB1inINf3sCL1SKw+o7bSX0mc7mR25
TwSCwR99+3wqgBDn1jMDUEB4172L/vfFxcPzwUSF48jDtlw0kJqaL0WBekmESH3UOOG1HqcdO9va
9vikBcZRE673peKLh4i3fNtDABYotxIHQxf+zFeOoO95YUfRCnYTVCwK7ESrtTsM+qAvtNu5e+lo
nJDLzB/aHmYCYYCOOKFg0Uj6xMB2b84nqGFHKRztBoe3+g44SEPeV1Ve8RxmySFjR7bgTZNM1B99
iQ+IOVMfFO6iWspHSd+sWSH0HxemITuFI928uKzB1hg4PpBFhbkgOOjFWhM/rw66UvXs6Cd2fbCU
iiQgqbt4hCAxt/hWeBeQ90TIlBBB16DFBQ4788/4MvUGbcWbhkqZmFGZbCDVTOLpHi+GqgCARiUH
o3plpevJCEt0NqESAMi8jUK0YewSICojM5ccYSTEB3EhgHcRNg1IZqF0Ek85INgjAOP9NQd7Hhsv
Kgi809PbStZ94P1Tk12g5ATGWOUy+KoJjYZpGjzesIr90c9kTAX6JeTieVfeYatfzbf2IK6ZPJ57
rYQ/fWOPRqPDVKIZoJiKU2ZQ4bV1aqyfBvVXoS83M5v2OKW8x8259Mp9aYesJpCNd4YPNclUHDN1
7HYB7O0aE107T7jv1D65BsUv8eqV9CQVHFGyn0noUxOmdST3d8Zeb8fJPrHlYH4D581Ipb7v2oGL
YvI4OiQ3BN5RoIZfU3rnYVTsVb75FbacndMN4qRnFT9j6BAP3iXq+i1PHAiVxHovPxJQqlQr4D2A
dT10DWmcIgxQIGA2E5rClHEUj/Uy5LqgBLjcvxz7EXrlK5kk7ENFWbzhUUQf62X349eaADwTkxMV
O5KZNcdnbcefg8pK9yGPdOK+FPbTI1PhtNJ9PIXdmVLt/kWKWoi/Kfae2K/Tq7WV30FeOFJm4AA5
QbtJoHiCPsx+O8Oy+J8x05BL7vrTGNZTVlaoKSUqOMq8fR/ATtLgJEH0WGkZgGJKCXst13jQHwG+
+tiKs8+JJR1tuHg+AFfpcoUEFDdVGWz/LpRgQJNXQzm+r/1y60R4zgXO4wewum57UnASLE09mf+p
+oxiN3A0BPYWCz6YnkyiibVTkQlhdeVLVWbMZRMowbdEcE9b8RwKWpqGE5TJ73ptH2D0KLPja/aj
hSwdhZ7XvnOo5dWtqb1lv0qaKwG8O1sCaXk+bMFzqPIe4TAGXEsBXX4r3nvlLnIxya38uUDSn1d7
m57KSBX8pmExXa8GFhYtORlIz7EuqgtknvV+NqRCVeYgSaAbZcVevPNIqGgK7skiN8pukikcdO3I
tRhMoNQz0vvdQG5ZNpJe8ZREHEE0rUtaqIUH0Xur50JaAr+wQ3QGahtQ1xS423eA7l6HjibhhnFP
L2GssbMbHBD/Aq8urhqmUepis2Lley53tZ5jB2QshHROiZNBxTk4cQJC6bKo1YbO3ZdQKVxPtO2F
NPCUJzGOoOpFphsTUgHMi9pNz8LmSRrp6uFZQ4BmeWTGg9KTbsn121J3+WmxbYmbX9A3zRzccQ7f
X+rM1xxDVT3ISvYM/DCJeoCaEbYpZnW7BXB8y7Y1ToLRQlCwN5bE5symDc6VZX/gvXymoDw3OtLv
1SlYeH7t/H/9Gfv650mQdGIJ9+gEONJvZRbEqSmx5EiqxSqPcmEPRUnx8X6E0PuMz/uC9J+OKg2e
eeEpcyEHZw0cRtJHvYl5iqmdysfola/AE/v3Dy/zv9uIg8NFKnmD7TzLVpLnTGwcFZaMw99PidV0
BY4wytk4t3+1FYkU/WCvvnt6N3YBcz3SbWCYVLCVEmTWDRiCvj/nqVXfuEJiLjD1rXdrR6b50/3+
psS/rttp7pxOSqt5VNBfhXEnUvKW0SDxbRJjh/WagxZOmBFTYxkj5WwvzR6oSBpAmu//1PGXbK+L
WgRF0brUeThdh+wTW07xkNXa1jxXh6VWwJo40zTuJQxlAiEe16yDsHyjj14zyDWDA8CZ3eeuAT/3
AaBPEy6ySs27oyFZA2INGaOKoDZuEaLkD+6qEOB1m+VlD3nbSi4uEctmYn52BQjrO/VZoqS46lpx
BP7XDIbERXC7I89TvQZ43YEUlGzPPTBTz8RvoUmGZEjQfB2yr8hwYGm8Tp/hsL4kXxf/9NR1pp6r
TIgB0wrnqShzClC+efsTh6vNQ1ZJIaLt8Sp2x2ujqmrO/9Qu8PyYR+49e9qmu1Dn25WAMtnkHprV
Ftlw7gZWQoLz+SxMBM7m8aePr0WCH7aIDqnAVug31P7Mq7zqGmUHFELeHKp0FqMZ1i3jVjqCzKEL
colu9wKS5UGM67RDg+7uFm6HwiDKX5W8+nE1d6XIKLFXV8/zdewIpkCCmgGSy13cizjqCbep8ZA8
d3D5eXSeNkmnL73VqAw8zJEVEc2Urh8xeNQFi0BP0KyNiKVc+trY7fuOgS+utvDiAP+lyj0GWgYv
bPrIa8stEFGjCuUMRNwSg0wZIO+388SsBosJppb1YRRa+DNezYHdpkjEzWSt3DC8sxTvGHLIcwHR
0YgJ+xsJPbXt4xX64BwUIuYyQZ+zncxj+qAejBcu8XDJ4R212E6/ZMJDJyzZtP+qpnOiLIHa7sIB
Wpuhb6qUh00wZgYEKT6uXi0r6Csbcwv1bDZlIuUaIlc5+mY7pvewT92M1UmgQYuMPfZGXhFvVbQ2
on+EATfl2z3VoQ8PTxSDdoGbMa0wCFdThAg1iFsuaL3a54o/Xvs8trV3qXR8vzeOu9v3Q4hTUVTd
E5VZIFdLygZnVNeVV0UOWLsuE00iAxeCmZ18qFSmla3bbugnxSNJqKPL4SNPBOCstQ4z5Jp4KSCO
9LQM6O5a+qJ4MPw/U/wNKA/r+gKyiEb/brLIpmzPjU7fw0jWu8ydzwAigK7vvig6GJVtKSnBS6er
+VBDMj1NaIMuwVkZAgV+FT2ef3r8pHn0lX//ALI38OKHdKqJe1yeRzHBaNWlQJyd6j/29OBJC4Z3
iVxMY6CIlAI8ZRgSWS5BnrSC1JDRjr2WPioCrvLbz4V6hCmzSMUS0Mo2ceUIEPletHiuRcKvLx7S
Q2S70d7M3Wfz3Ab9YLC3mzj7RA9E59iWf/ii3ui8FAWLH1hGqZTDdgnoP4Ql6ncQtsuhbznCk/Kj
a8gy1txin502wmwGN3KaSAt4qn1ccK0bdkuPzKZnBQ0SVXP71UiGHxHrrnBGcSBI5jGN1g3Cz548
OWylap/63r50H82PgCHsNLGzG94q5R2mqTCXLAICslbouC8jdrUygeRPzfrW83I5Tvh63eAjoMeD
IvG6Ou1LglSRkTYoXn+PXTxm2bjEfoDPO3Yu5t9KzPZmLyeRSotbFxOfTwvgsNmVRftxrGjTxvqa
q+Tw8HG5Wi+t3FmQjOGPnssd0rnCyIe43umh2PFy8Zhie3WhvXHopZ5ysVrqSVtC28IakNm0uPl/
h3gjSH3HdGXocyP2BnTUscz7f3JikpunIKoKwr1qPNvQondqBjLmrKhN5mUQ5J2V/8UXymxBerQl
ZB1GK1tT9z+wlAj9S+jbymaKxnJB7sruiO3qwY+x2lR3+TAhc4J5UoxTR/sbzeyNJha1kvT7+HCn
nT/LVD1vFV3tZ/FkWDXdiB/vkf34bsowqXPyZWQEgPz8TlLH21MR+I8h5SSCSHi67NYny+BZXAyJ
oFkAli0LOJKQKJqajpO+FWD0q4cvvZk3upW3G9cz34cmrdph5sSc6IJJK0KBIAYtyLpvGaxF1xVS
BQ9ZSmwzEaFvw46rUlw0vz+a/2xqtUMxpwkhe78ktxUP6N7jreZmGjZE5yqjlr27KB8fO+sqC8xo
R72hqmPDc5I1aRLdfoIjv5lHTIl+4UAtO6OPxdL2wNFVvWHASKmC8aLViiO2h6fgQBPdK/wqHV74
nrpI3+mzkV7kgf7sXNGyU3hgekdZ5XZcGcGrhaYWtCaS0szhS4W5Ui073/TW+5CI7BZ/PZ3zjVYL
k9+bp3jpqtGlWxiVXT5aTBBsENx57Q3v1mX3WxZR58A9D1aM1e7Ap/xuUQRlR1jyzqpIp2zlGWjC
z6cW54nyAmpm1o0YhDSaqxY0o0HL0KcirNWOrg6k6M+RKBWfmCz94ITJms7/Bu8V6dskEUdCv/FB
JhicSwBEHHLt2g/m6s5FByMynZ4Xd09j7r4EIqhlgDC8F2p2gBgNGY9U3lVXeYcsLvjiXA5WEwXZ
93MRwZPTTZ4r/+9lTzebsIvyjwPgpYBLKMeiAvD9lTPcsOe2lptM3R4TnF37TTsfqjSaQOguqFE/
obSNfKyJnDjO8UKLGfHLIyJn7oCcULN6tNih3g0ctS/d3FRIyXho6qUSDHredRV4OIR/+nKTfH5Z
c+U5hUQqZ04M7/DzKdPp4WcbLjgY5t7Pypj+QU5WPpR2/gUmWkQrtzr/ElfTQ9rg9EsuxD3eJbVL
g3G1RRDJN2pJuv1FElb4MXofIrdc4jq7rUsm7s0Od7/U922+BW0kOq+Y+T1wOrJQG1xurJ3v7gmR
UUAITzhNjpTI4uLo0+L1v1iUhGJPMrpMPA383fiegKGozaHsmZg8lOlcJnxN4g1GmYkHpK99JvsV
ag6GGRNbVKcyRnUNV94r4DLTNbIzfMDUE1IC4FDyy3XtvvB4SdevFXT2pxcNkQ/PhvUFpiEVNmhb
d/tSVf5JlBbi2BCzdfpLdQ7tGkMdPcsauMQMgfJPH4fD2HeMDtH5d+CpAtT5e1MQUcq5lEqbSRv5
ezziB2agvZVCrFHLyIHZ1WNOeqbZk7s3dz2dWGzueccehaCSsj07Y0gBBm3iO1/Pu3d9zoYjLMt3
w3vC4Inh0icPFb6RiVIkkPKbFhhI1Ey4fQVRA2l3rbhMWnsvdJiYCICk0tW2kPV9PAun5CGctVFk
08AVIPFdVwl+CqBF8nO8Ht2YDLOf+L34e/U4kOAKf+VGnBi8hhO/OmD2OFtw5GQL4/x0eioe52Yv
Glh5VXaiiEu3bfxjn1LW5P023IjAtzizya5nP7/Mjo/ODAdYzmnyYCKOvPAQAse2AxgbOcevM+ly
3KNjGlrVpCQwISkK8+RNj/QCIQCP1rF+L9EYeiZPkCde4uspXluwUmLno48HbCJsU4NFpBZlJwrB
H1iZJWQmxGB2j+cX1oizJ6pLKyUJASoKZQXiNd4uQ9nJf/5Hz3xzYc4zze5ksIxoSsZtfXqESHWg
FxqOriFWzAFXqE+i+UqINwjfTRhFLW8ndoizjJBrjTj8PAFT3qnRuts9KrX2Tau/A79aWwAKmqV+
cx3Vx/eU0ridKitmD7ZdeTTNCDD8Qepr5+WcJCXZBd2zv7rYLqYqZCUDd/PBmvIZZIJYNYn8JsG7
G1Sqjy1U/0L4nAx9QOJzBtphlIxI1jzALzNwn8RSOgTKsuBRiBbmdcS9ojSGvIfQf+euMncQ+2dY
TEWyXxcx167qEc/AJhZ4Ow841W7Nb8m2wqjgijdKb5sKzj5+lRp/lrVH6k5j9h6q+zjbAwySqq4Z
FBg7vLNl8LdNfR8eSpQ2f2Ds5xQw623IdAZQ0qnWmo3gOQf6n64BnO7gVKlKzJO/aicqlx7YH3RL
aTK0NfAaIWgmLwmBa/0a6BWVTYrGcM0n9kz85MEqBuR+vHwpYVFjK5RrC2j8C2xbykXkxtbLxoi2
tAZAeIISfCf/I7Y4go0oC+SfvHI6fDPx/q59VfJY3aCjcZLrbCC74ymuNwqcc6aSfs55w4/tol3w
OTUzsJGSdyVoqxM0hKHHmo+Gfxw5NOviIOpjKW3jvYdiFztd8sgLLguZBFjNCUoxhB+Gej019dZk
Ej25SfDS+OD9zx3WlNTfakV1VqlajVjo15CKuO08kcG64jJGOX7JhQq0S05FI4xh7Vhhh4O+6ksb
HTZ9wCvfIbO6bhOR7Qyqd3dtsopVehQxnSKDSYRxf/EP3WQDOEmlU5ii8hVp4yotEllfJ7zttQ0y
WUvJXB6jHi4wWaILvL6HgVswMKBg9Hvpot1MXcHctSzCwaCdokhXZrhYjyepPDLSWOY8qfb1axWE
TASdJ6At5CjAOdm1Vf9EFmdgFovyQwMBMnQCpYxDAQQmUZfiEEbuygOzHOMlwxcVYACHQkTH0Uy4
g7BHgQITqrEif+cKfOzwFpWgiUlA59bpg60se3IpAEFPDODy7cLSZX8OkeHCjjLu+ExN4usRFoPB
55LjpiYV6gxcoqPkxNR4Q1ZiBDCZUTqZyx7XDAwF5fXbBOiTYuOMK8snMqH7fOucGwNxlBDreUqI
SfbKz6vZkhIGiCejceXHVzpdlu6dvZ/8/fOsb8haLDOn88GFew/OcBC4w4N5YxyJvbGzs24EneUx
taO/I/tJ2hkI/TDXpCOMnKkia0Kupzq4phaLxgkzH5sW3jL3jsvlSyRle0bTXABif0QI1i8YD0or
cFhWT9i1p86jOqCwtJTXi/0KkpIOr/zUKBGeJcKs1jVkCLJYZ0eKUex6eurviXdlalpf2SbpwMXY
6gRwI7Q78Dyk3usEp6uXnVITn9wmy+QY1JSlHIDfOLgnwHsu8e0ATUnrZ8ybaQkquzpxbYTcmJsj
DaFj3fEiEJyhOfLAd9TSHXMbLutfBBQIQx2dDMfiqZSnLc/jbTNxnTvQKCqaf5Nezmxct257aYOQ
0Vk6q1rjpOkLZX/VfwHnZWdOeu94+06fCOxmBRi4TX+oqoan1LrSuLifKJ8dqFM4thv02MotnIO1
Mqwy8of5EpQ/6q6D2xg/CSAmJVpPB+qo0KtX4D/uNVR24OtdoidmMlgfecNhcoTOtb/WM7wXuNt8
fx0Ke9iSUFIfN1NhVjmPOVDHPOVbdtS3TaqaPODBHhMk2mvE1t7ZBTrhgQ+i/6GzU5i7WjRE+l+m
yP58HmciBP1PJjIlQmz9h6X49PO3nBCSpux1red+qMA88oZ17eIUy0WhXy6bsHWnZlbhMxwFbUrf
e2UXS/q2XOqkh1NDUEJ7lpV+duO6OmPFincRdbNT4/4nzWsME+0FMtAHq5v0MMuuIUY5as1Kpxyg
+IgxpYdMRn4y1xmHGlNb15CjBQe1l1H5GA6ydrjZiKayeEtMjlprdPUW15KRh1G0ZljsCrewnZZB
MPw6Y0CpDfu76fnVQda7Vaiqej4gax/eGyOKsBoD85fq2HctvaXUk1GXKKLdfCRTKG8GvQ1EOy9o
Ek2mW0zzYOS928LdePh8j0JmGGGM6N4cRGx6O+8VM1MdiK+FePr6HmIItIUipEmFk1CxFSXR2iU3
IOn8zuzQ7jfA+p7xvRHWsslUx5XYvch+9nxnuzxtIc/n/V9EqXHs62+BPnYeOtc8mKcyESklzmpu
/nNu8XdJlBXo4VoKp67Wyo4LYf0rB+32aGgrv9njc/bb/UJA3yRBaW2w8+K3WF/dw8jo4fsG/ely
Nhqh2XPE8iZo+wjNMGZ5/gOTQVqoFEeKHcaXvWtf3IO7eBAa1BGdCqSyY5AZrydzNZ8zORKHrN8J
z2ape1g43deZ4p2jqEP60rmsUECQX6mTVXB3jD0X7sPCEqva4Kp1piCGwEqeN74Fv7uEDkGF3hYt
d53tFugCprBexiwR2TuHqSBJQ5hRl60bLCGg54tX+gQiMtluU17foyTuMNqyKjsgJrSyM0dSdi1/
FUk8XPP+RD+WFqTGJq793Xj+Gc2XcNHFhX7g5H5AwKG0LiN4GIGPIOP+UmftOzqIw3oUvxa2XsP0
FlTPQb55ZFHQLIIqZqTpygqLMmCVogE94nHlpiD2SBlrkvtG76lquECsNG0RKyol7+9R6YT9d470
lUXMGMAkd3P3Rthx73UHCvgFYwFzKq9eAS7JtzWZuV9718QgMNmArhjdAs/oLM2QgijVpjdIe6Ox
hJ7VMJFNLNuLLhHlBwfGKLwx6BG50fM/uJpkM/bHbSvbIfApgezuAAylnCL/4mJh5EVo8K6e2BqH
VHtf495U5vTBZqw1YEd4Hyojqn75UzSV7QbTbQvex41fvY/2BqCMpVCD7FTsJiXdZEVVJJQ8I809
kHX7u000Z0zUmx8UY4FXUhyKFeEc/nIc/ZBtIK3mqKrY92ZbUESFGUlxJM549mG7dICr/1yEpxye
JxaT1c/y9aIVMjNBqvmeomtg+fSkvCMCRufMZpqieGTqZYoMpDYAEAukNUUZOUFvN03Zn6poiD/8
Np82fvKd/FZl7rpiWW+qIph/w0IekH+kVCqt5ppHdGHi5iUgZFXhuAqUO4smvgHKknC8z8xzQCQG
sudNDajuz6xz231QINH1Iq5ndMuMQM0Y1VOsKn/b5VB3BMfrQn+aBb5ZHMKMMy8S04vitplsyygk
rYX4AWat6SN1eom7i0S2mN+IE9Xf/edYxYofCudTPQFgJNPst3V8toWcnkoS5Tn4QEdHZHJ9fkEg
c6OY6SFdJeCkzAEAAgg6Fc/GlwjPqAdS2uWDvTEQ7KiMguAbMJAB/Y7yxdJWZOBjZamuZO0t8mt7
lOBP7VzW71IUVbPyX5foemLyV19ZVT3Oe+bCnPimfTp8y1AtaSHt0CDzBkvmK87GWjxYlAs9KTc8
hms2JlfVlCdJFmz8dP/7OIm73fo8vin+oemEffndGn8hswQ9o875tE7QLuDxuKBN7Bdvgz5ow2B5
w6hgP5UjPLWSS9F+tvKnKDR+Q5m6fNR2C6MbMUgbC4DVNowQFyAVV0pVqoDf+Tj6rvCUz9cjv9s7
xDyiPDpZ8jzOfqRSC0OyliSRKRaQlLNfwbr6elk4NGGeBqk5C0EPC7lyDQwNmc7LjRbmP+yLojLT
MnFKk0lRMrJJtWb960EW5V23gqiU11zHVuCUtYq2uYljtJLBwyxilZ1W08e7eprPNPyUOBrF+WTz
EMHfhJwvlZMPZ5JTRZjA2hrpfqw5uC5htLNBcLWhhBxPS+gyCgn2RKJ5wzpmHGMO8ijXeBYuTEll
mr4BMXRT0y5BiNblrN26a3X7Rnq8BSwUZ+rJkTrbF3ZWChEYLGWv6AGs1RUN/t/omu5nx6z+E/qk
XBapWtEu/I5dxl05+o3yrwv1ZWFgAJZlMZ+ydXmuzD7iZeMGTo7CVMk9bVgljFDdJvymWkq6Sl2f
nbpHKahb62s5S+mlTn3/pMpUXpf2h8QEMJVhPVZwXAtQnIa9TEYXOB5e57RSoOqnGfiV7MY0o3Py
rCxTi63KCvTXeBVvMN+f4O3RjffRbVlTBRcoT4ZHz+isXBZAIsZVPSLN39aGTBJiJfQ1mHTUmg8+
Ii6yP7IvH/Z788ZqjnqhoDW6/TMrtWz6f9S5ObemmGsc9C14q65u4rnLbIPRlWbk+rzMcGZnz990
h3qL6erTu9wNR6SHw7IhzDXuHujMw9346U5/Od88vO2lM3xHpnlrJJLqUNMTVQAhlgQE22NZtC5E
2F0arZMtThwQMye3KcXnNYYFPtpW3ZzWn4B1EhW06K0/XU2sUzm8JjideuUhQd4GwdySqHxX7c0j
vVr6m2Yeu4l6Z7fEBzxtKDODsWVet4Yy4sRGjj57Tdc4A1u0txDz0w3ea1jSeqhmOvv4jUcqcMZI
qz2gz8eyogth1HftsB8IRhAXoHwTmDmWejjONwz+40VtOWtytzOZxqwMwd4K8Oe0ySXe5zuzT9tM
BwPhs2nCzRosTibTSCjnOWLq6/IBIeorI3zhXv0QvoBYhxUt4ZYIi76aqbdkDkGAreu0BAk121oR
LMWmfLUM78gsxra3AfB9MYQj6R5mvwqgXZfEcfPIJS7R+xdGVBhVWzSc06EQoilJtcu5R01iev+9
Xzb9ERm5Z6qEkCSl5lb/WFbtPA1OgEqT3i5Qd7bSlPFTVGE+ARhApu3xCkcykC1ta7pNbMPxNh81
pT8/g7Ndmt5rYxMVsQclNuvMhTJsNWLJrcFcZ7+8M+RKvTv6/AY1A4oaA0WQGBgd9/CDrLhTEdpT
Ab0q2SI7EmtQSBiVqtsdntRla8rhTyyDD/sDgB+qw4kLKnDtUaBUM+IA85oe+fSmVQ3FkMXq0nDV
3209XqNLvR5EvI452s685yeD0KepqoOKMzK+TEmeswEskTa6S3ATQUHlq/WqgVwN3+QFrDZfMMtl
uMQdH3cUHoS0ayP/rVpwLuf1kknASiZvC3IbhCuZkBLTTLwMHXfXUVMXstNA5NnkF+XMsmU5lUQj
MMdUDUuxzVgiuZrQF/XUWJsb3U96rq8fdd/qFZ78TTNrw8hS09nGjMSPE0uGXdkMJs3hzCaoap6h
/dx7xOq4JzOLTI6L4iwJX4ndS5AKYW9DpNUvBq9BKBNJD9AQ58LmlhM1u//fOBfJrIHifUXu9aZY
PODCRCpplrobAqQ+EUj3FTy3BGBkVVaW+/GZM/RdQSzVfx1V9+N2MX73eERSzWuLbVrXDjYSGq60
vdzRjuyQI1CqHDR0GcFkOXkj4JN0LSKi7eKEKF06LGAtlVLbThAQad3Qk6cVbf6Ep4bn44m259SC
BcWdfmIiCVhuKH3a06XwXiK6rDkqDz4X5jAYrjTALYyKsWk81FiWqACEOoWFmXyxZ1740SM6Tvq3
w3GbZxIKVcraeGkWy5In3OEJj4cJnd6L9nIaMTTVATkT6MrDelc2cDfnfpvDvwyKfKKqfLW604yA
s2QVD/f+GarPsfc0N6vnb9wD9xHDrNSSfX2IwnOhk94Fm5wDYCHzwwlWDATpweh+4be8kWSmjXor
bbQOEyFOG/H2SsF7Za2Vsz2wdC5Hiurasj+2fRZsgG6aYn/ow8k4EiMP22x3hm2/3ufQ3D9iwJ9x
ZhLi7j1zWi9hXtFFthyZsNGb9aAbyQPNR7Me7fjeTWZ9WxNtOK2ncQAg7TXlrvsU0RbCXnXRCuWr
tFUJATMrzIHziejJ2WJbXdzwleZ3XUqTI3EarERszNayJjHj1v6dHF99W1iWCsH7MFKfyd1ckQ3f
s7pBlfd56xRZMvyXFAzObCjs7fohTk8mU3p8Y2rWqggxqUNKHObsItIK4NrEnI+zsSuUO61bBcUp
yLQTSR6n4rxYZQE4hY+UQHfBAtuGBI5DR9FrC+FtX1EKm+ZzB8EXNtbJMakZse1gj8CcBUhFxgrx
HIYWfao3ZEmEQ/14/idiGGTVUqPUVRqxT2KzmOfyzW05jF7AJXEKLm+YNjgNW2CoXzC2VyUDL/Qm
IDMoQzhzArdc8LylMoSSLlVsmulEFQOfhy88jUN8rfD+h+EmbnQaVFbYQb9eoA5J6TMvXx9rUyyq
JR5Tzjl9fCNmMIiiRmrJbKREN3Ast37eBJh4WxKLH9c+3gvT3tb52ZX2Cy28LD/zTbEOInxgiJJb
bXilZaOVxQW6MppsDAX1MsQAtm/uLX4lGt8k/a1oWZLZ1KsOp9vcCWhW3jY1Wu0ipCdelRqpeSXK
Ev7gWst4gPOC36qS1Uh8W2vT0i9XhHHLB6XnPqZLdp9guOO+lOUtF/a5IyoFel/1jnZPxPj1YbDp
/9DGOxjW93rjCeYdivcmWH/xH67UhozSlR7WzAsUB8z6WSiVLL9RDFEfuBV/758xWcF2UZ8yOlJ/
xmrkRHuwLUBk0OhIPiCoWLchIyVV0oiQ5OtYTTXGxi1FuCaRKgiIm3PXGCv0SzybIMIw81Xwj9Vy
f227GhvKD9BnsXeWIYWk1AIPREJIps9UpItbzflj5iWFdykdfw1PmDKldqt4eKBLmUcvoY7FCtRQ
5E1usTRcfb7NXBjAC//KHLJzmWy8bmWC5sPU6Iyo415HG12TciYv3jfP8fpIadCIUjOsJm4uk+Lv
DYzauDQbbbhayBkfAm9AftmxKs+31wZbUoPik+T0iM/TR4aF8qsm+k0fmVumlfxkWZB/Cz9t7uwT
q+DH508YfPsNxUxQ60TthQmQrHczgrR6Um7iGiBRChv0rwVygPl9eXLVBWa/kQy0v9LlvBef3TAq
cmKDgGxGgVCK3yiiy1Iql028YNP8oD6IEBtUus6n8hwpiRHS/LosN76LSEp/SSW268JOOM2pBhbG
Q/8V0gqT6djApOM2uT39TC3vGgVywnb7tLVaHF6PfU51SDaSNBmR8nC4X6t/eUycb0GYYAgMWODj
K5/f94XXx3ZcNGrCCCftuSQAdD0t4XcWHWSsTN2Vd18aUkCyP1xj0gqfgdP36lYIklaCI/ukWgfx
ncnS9nQruTtFmY+sczZhxORpxmjD4qP0yezdhGLPEdFf3f8mwWS5QJuQrkfj0+wrpaea37vjHSal
/CvxHZXaCL2enhf0Q56QkaJOqz3saDiB0xyPnXVbZy/jrNO93iNqdxCTSCB1P8Y/560kjDBAvWY6
wtnSG7puDY7Sg5MwZsOOJqyG/+iB6iwbFZ1QFqx6Lt3tZ9dnbMx76HIVBxRTk5TLD4VLMDznrf8H
Jsqf5l3yZZ4FFJXuRQDJqyYHfsp0dwl54eh2Yy70wqKnaZD5LIgsuZJMfpoeDPnZgZcvpJiWRw7e
rs0aLlNqOSYoAyyWHphkPTJFoToFhnalImOozqlNx2hB+YJyvvKhhpqYwYszRK14VKWETE6k8Ux8
DREpWeJWuCqhA/8AZKT8xVlnfP7WCDVrT3PI5uNHBa+1/k0awqANktFtalhrQo/MkPZrVYHb5Ko9
Sq0KIsq+dehcHCtvrmEOM9R2JVHGX8pSUHLUSWTqjmW+qs+uUlFOMHvdUEbmvHUgL+LaXTSqawtx
olhFdqBmKzY5Xbn4K749lv+IM1vkb5EuKHEn7ZmelSwtDt7fTt2T9wlbVOmlM++jY2XQH1kkfx83
J2RcUW2Tqtq4CON4Dcgv3ISw3xXdtRdC0wqdFpffgcj8QU0DTULrhcF8sotRgQU2k8PVKYFVZbM7
3OWBtTaHbs/99EoH1rCGLT9f4NsyfSZmrjEdFcTcD+/o+A6y2OZLLx2pLnCtlIbveiJDdlwZwxNS
NF9QmlanWTbBqpxE/7vOpHBBcj/PxN1b3yNkBI+CVTTH5iqeZk80YuZCCWfb7vO/QqGtHjYWUsyG
Kk4QuazvjVKJoxBY/nrc66thZGt7dtHKujJ1F99rkiNAzf2f0BImFfEN5dgyPt4u23FgNX2R+oN+
4fmHwgsUESWNZlLjexHyB7vjEIGX0OdxZc+vU2gHlFSD94DFkvmdy2Z4HQt+ARrLI+l0WUaN6fAw
xpZrqDH8/iE10BD11g70vuIa6GA8T4s58b4rtBmVAJovGChYeSEtIiIeYX4lnIcslQsxX0NwRgV1
1+suMGT68lUkQlI3sIh2C/1SR7q+L/5mOJwbGbPclFvg26hid8GQb+39sZk2nkPZFAnfaUD5PSgu
BuQywdPKir7Yovkt8pb4oOyGXhZvKWV+ZXI7CmQWw5ZltQJcxeMFMikc5yx9KYM8NS2ZIIjHymsB
z4K1V3sZoVJU+fDSeuJie/FsRARcQoQCWMHru6Sgw+V2hiXYmxxkarXNoOOojj7KZUXDgmvdjzT9
+UruhJKd5thNxaDDTbYR4tjAnko2sIvZA+oqQxA3ZwYDk5fuYEdOwziYNm/yS3ofuEuKBQa5BYlt
6a5b8aVVrSjJyQyXEO1PBJPs/U8d/7ZB4ItqYRknu6WYhsITOVx3i8b+85Li4A8YxgIooWMlJpGV
YUG+pn8r8SxRTcuowYXD0bKmIClAwiMFiQH/KyNjdPfODv31x8hrbiDP4IHNS5R3FCEsZetDoJ6+
vhhD38JnvzWUeicMenw8dtGgJK+uEYEQF2brKOKY9oOtRa8CX2qDj8/k6BdsfxCd6eHv/ww7WzBZ
Ih+qdmKsyw9cenwmSMkSZKvcjC3iG30hS/tzK1y0gSfIQT3/dKqWOR5Rygizsou+vCUdGoy/AGCf
pOq043jB7Ek1vXFdczoXtHYtS7ZbbMf0/KQmEClRMGxRplnJKYkRttBi3eA/QoUd4PG5CTNdCsMr
j2IeRZ04qjJxoQcdtFBWhReUdNdJWRI0yPlBhXnVesUS3Mxte5gTKAGWeqkd6zN/hKK3z/RCbe8Z
lXJWcQR9g92l5rOfC/319dVaeKnY3zeCKNXVok8Agqcb4SWj+0avP8e0pQfy0hiK/N9IUDOQ9mSi
rQnnZyMx9pfFaKNf9nc/U5Nni6KcS+LVOj0HFvzIDEGxZE2LbWANT097sVnQTllqSjxY+pZZ6QIv
f+PNBYQ//4wYn72mQvzRDaU4o0Hpu/vlCOzc4DYk1a2k6LLP56sX8QM15d4JFlgNHVjZ/7r4J6Xi
umCWNKSDDn2xIKx3wjXwPNMokIeE7NPTJYNh+PDDYZ1rKLg6G/xGcE+PtIXApFKPjJzwoBcebx8w
Xp/XYmLkauZ15nWOwZzdVHxnKTczl601hW8k+pgr7IgSETIqO+VJlz8vsZvGzk3wxXAxY9JqyuW7
cfmm03I9Q3JFiJeVOLyDmEmGuCrqQ7Hmq+QV/LZfLtiDnOTR8lhgR3IBOeZPUTpkDSpCJIwD6Jc5
csF82vMp3PA7fPEZ74RqmusK+0uoOdAXtGDBxJcx9zI3cCGE0QH+IBUYyYfGSjzkUl/mplM40PDi
rZsTnx0/XQRfVClWGvBYhpgGOUNShWzI42UpIUsrrpfnzJVsrugD/mc+RW+VbMu53cVca0aiYv4u
E0dC6UOUonQDQYiA2tnsDf2XnCMf8FoxHefdP+bYBoCQP21aG7ZuFBH2oyBcrJPVjLltnLKTkeZt
3ePoVV1EdVggMcdMzJ+usPVRP3bO8o/zUdM0MYH2RHDnmNt4CP31Mgtl962IWHI7Gz8xnPAZJfZv
oT98Fh4rY5NDRS6NB2xmgIuU4rduNJkSUYhTD9CrP8X+C2bVY50p3C5TIBzd2WvMtuz9iU8LPix0
yFsWStbSSUv0NAFaG/lOUqql1rcRartV5ve+sF0Q0vQ3cGkYLF49r2uWP4Y9lSk+t/dECDvY/IuO
kJ478XjnbG4ijdPUAN1dcxRsqk/wqMQVhxwseiwIiyNQbaAn282ejjye4KoTuHiilnfX34SA8Isr
cLjfGQdDxWeHOySY4UhaSXTOMvMnllmtycwl0yiWuE1va3W0omzMLDU9hj0IsjQbs+hYtLiTlTqK
CzMEj7IzO4dWi5KZsyAzJYr6kwnc088oau0gLavx5UmgNV20xyb6U/lsZblpZsh7LU/6Y4CCJooJ
2oYdHjGwRZuLmL7ByOyCVCQJWPHnYpjjpVMAFwPrQWsfQ1RJxzCZqDzVG0wsxezWpwKnQLggl0uT
PP5932FkJGVOikymbxIDTeM7Zi0LX0742VbfSVlDfzQE3MtP9s+iVHuFMRpYOBFzfjYwI84hJOUq
snzehfJ7gQEXbmLZAfvuqCIU3k3p8pFVYwav9rvEW6JHldKU0vVq7A74dOJdM0/vFB5LN6pyQmAD
fYhUiWRSM11nh0mL4TAYrjPrgN/QInHpur9EWu3vBxBtpjougW8eHiVC1+jmoGworCmoIG6MWgcu
VGSP0IvzT+FiXS6Mm6tAaKogJ9xVb0H8+xL2bzGMAwfGeltUq9VExKF8WMzzMNftGMQnDIsp8Wt6
BAPZcRCXTWtRhpDv6N1W2wrTrq7eFsfi2Mw/niSFfzpTM6WJGLVC4k+OxkpbMrTpVP1bQ32AK9Q9
iKOMSHqiZ/HcTofsZmL3hcwYOHxySqJ6pVLmBrJMKBCB2kwgAfB+QRSPjrGBBWqGLrgknhXzZ+R6
lnfQclPSJ/kOFKDklb+O2AsSSjV+lahHeRiGN+6iG8kCNUxnSy5UvHpz0JIDdlvEGveJcHDz59rT
74aUhqhjQjUxpnNrx8mmOUrfMUGF/u/4sl4xuOitT3dGdTyB/8Vwd1OIOhZF6xV1FNXWlSjGbyj6
nGseZMidnaMAYRyMQQ38tgIvcbIB4y4+ROwCB/9U2L+Y3fobCMKSnis1CsksGjUJTDZcrZ9XknWO
Qae4Zi6RH6xmNlELMG7S0lILTI3AhYO6XkEh8/vPGuEA0pVKAUTTba6JpfUuVx2kE/SuDvvd7VdX
iXmSq0eOX4IrFHXQwSN0vQzvbh1Tbebnhr0iyoW1G2GeRaEdvHtZiInRtPZfs4BIW3yUyLxXucAV
00dxf/0kuEtr3xKko5iFRVBhJgLPkqIPcB/BnfXW4GJiWL5PkEjk9UOcVYEFYrI1uhcebAzUdnL6
b2hf0V4tq5bpjpd8253ROpfUfGx4CYiYPTsOjJi54EN3oy1gNSPVMOUKyJNvmHxKLLL/jx8UqyZj
mZQ2oZWbP7PWewKyeVmz0Ks+ZXwe+rwCk6BunFkmxGI0JIqm70q0j0Rkn5vWY1esc0W2gvlYgY+q
iWJFNaTXhHL9e/foCwmqC07KpZCNh8MBDd6jJYiQmEz0jFRdkeY/00nrNsrLSQXek6qzfzjuRAnC
ombJBOtlQZCS2pjM0lH6R4wWZKf7DPqukKNGH1qAbIrsWiT19zjIqCQU3Ttq1unKRmNmxRmVBa+e
PROlGSND7REL1UY3j7iCXlNFBUVOMLz4HQgXxlI4Dx3cRes/NgwHmPpIqskekxsGL1/BLCs+w7Y0
msd9bNk2UHPXXdn0hbR8Joi8JX5etma65A0KcrtnHoewMxCM+r0EEFUDYpdCjSsQ6W5/lnzyTgmO
2p8XJOeemmj+D0ianOYhp7NmzgmPKjVJ9nzVfuY7gjwQScmiEi7TetjwLTnrWXsiBZzh/g8zzQ/Q
KrqAZQNtjTu9iap9aFNjSBXSjEn+S4h86Jnv2rMf8FcWc1AXuqwxbzyekAAelg+2SEhnrbTCCHx8
b18aHgg4yyNMXuYIEJjJEg8fiKwOzFqnE7gbh46RWv1O7wCwYC+RI3bz/cFECpTFQML9eKTweuw2
hbTJSPCdFv0Px87GMJGIYyVCcg4JLW1AHY/4mHAlEYvSTZlezjRrjQwPlo40ozFUfXsGywBNoudb
AuJeqd36k2251PQcz1MJCH0mG97tlVLNQzlclyPzP/fBnWwEn56tBjqgverszS0ZLahCnbi9dvDi
Rg1+2ggrXOGdN/JiB5JTj9e73RUjNyFRIGf/qIac9GIYxcmOGUOhwb3Vkrq+KaomBA6pWRhfkkvk
70Hu19ZIlFqA00usfvfhP1NgNik3fAyKq5DdMCsIQMVr4Aeimzmao3/ES0AGhs/CbJ9Sosy+dNgF
tp30+zFCaJ1oi0qVa8BHWvTKT78HgjNRh4MFXgF11X2t3Fvze+3LzbSI5DCsGMXy34GZ4i9f1P58
zKScX5Cp7VvgVzLWKpFWk1PjRyfJLf2JqVfEkHWIYumPpOsX7A1K++v30PNVStORozg6JjX0q9j3
Q5lZW3t3TP0tbIdNbLo7qQQzgzTTjJ73s94ejkAmIlapMcyzI9y1I/huCJV0heoEczx2ABy5tBhe
4XzOaPORh6DH4IL//jsBKUQybRW+Rq5W45gk+cHyJWJEJNSOSV0mDwGEH4e/b4L9VXMpuB6pw3W1
ACFqHQLt0hbPErWO1qh+jIcceD4RVS35WLUwyx/zaljdk7vG66kZ/eOi3Vi7unnHvK/A1hWxI7YG
Cf0RE/BrAkp6YSB8hsPqJCyl6f5bQZmX0fFtg6CI2H0bW4dqllN2jPZJmKzPEK392U1PXmKmrakN
DUq+TKCXreHdEQdihU5Dpqoc6dfFVif2ArJWgMOpVFXdDeUPyEK2TYgwZRCyn4wNFuicaPnbz0Bj
x2+WVizbureqsZaDHM2qsFBdMWmoejjvK5vbso2F7ciauIwuCxpngzKOfz0isjA3xTy1I7FkWwdZ
WINdgj5jLlFlM6PHyOzE6rJeMZ1j5HHHaTF495QDldVu85qv6hY9WwAvTEaF5+BtuEoBBME7YlaW
rtdcBDQyE/ugcsoFqqY+Z+tvedwhk/BnlqAxYc5hUIACm0e5goVKGI8Ltlj6bJCAnVJ9Rta650kt
GAdGdu07M/ovKVMgem1MkuZNi+GqTBT5q6TorZVvbiFUFEyOJEyVpDySZ212fYfR34OYSZaW//8Z
UzUyTFJm6Bvoj7gzOLMPuo+lZnLe+5j2hVZ+utWWgaAk0SIHjX0a24EuNr7nRVJUl/WnoPRKsNZN
kYT4C3Na29XXudTCRBv4hKPfgwyNgWfRw/TvP7i75zbhRYYujZhvgPDjiSJA0oxOhhRr7akoEU2c
nhdQis1WHt0p4c4qAZEfBONkp0qbgmz6/+jnR/xgowAdExPinMjbCtw1iuYREYPKS40SXaWr23kp
abUnabutB+9S1tPLm9/hemZmNGu8TDk3YggEgW8Z3/nlrkJWp2R4GabKRGwdxCjCwNkGBzP6G9Ny
itYOIwxxS+ojZxeL6DHrA4cbw8Hvdx+bIRga9QaCzmeCDZQiOCoyeCGWZk4BdJsuGTnaWcRmRF2m
4kFwpQ8KT1LcoBkt0IYmXYEfn/FyeewE1fQIOWyamMvKy6QQXPSCxciC4UInbn/UYQPVF5+tWJ79
dEEIQ8qwcaydcshI2J0MVvKF6zXPD0fhlI0IWfKQjmh9s1BtuqjjVtheARSku5YGgsLMqLvxOkQ5
uwsvGstb81tZYN/2u1oz1CCqIsq9wWgW3Olfv/DlrGqVdQ6fwQE3MPd/MSg7IPUkxOtpVxKyvLPC
j8yjlLUyoQ7Y8FC9oShZXCEjpGHgmWlLd0U1P87is/oLDk78fBD4CvBMSNS6TwzM4xBbJhpkE3XF
03APYQpVq279AnH/AIQvv2FBCpMzz992aaayp9dItkUIfiIoakA3gCURW0+B/12vXATD6C6XNbWA
i56x36OrZefB7kdLmH5bxJN+Pup7F4O7/FmksqJeSjs7rlc2wnaG2T17HOEZ3M5IRJdUpyTRQsS9
cdFU50xBcqz9OKYkYpZGW8HknJOxXU1LyLgbcRZPf1Wij3TkYUvMy66tMdtD2X9mi5z83z6sLMNA
K3Z5bgutW2514wk8wnLuEL+Izwv2Ec2yIF/x85AKhWsu8sAME0qJ8pEl+cDgwXv6iDwK18aXWBYv
XAbNW8jGuFW5+BqKvapawM2bby6x2az0TgenJ1CdTZRhHKmofg6KoXG3Kt2aPcPQB+JmEPW/jKZ4
ESjMhR384wV99IMJVx0XwMzXAy6UvR2781EJ1uWu4O+yWeGVes9hQd2Qev4GoMOcnw8OjwY6faq2
NJKEWuxHE3DgMbI4mJs157dQzpUxMNAHoWony/2OefuUr1mPykm2gqYEQ2Dm7K9dFts/F9fj3KwI
5cnklC/yoUUjKks7HHu65DrEToTtMVF/rTrkasFtSvVlNX8tmwZgzpIypA5USWFjaabWxDYAtl4L
fgo7r9kr8mBYjzjYkAJpN6EPuSKZvmX6aeMa0aylnF2J6ZBNrrPIuFNpC/3JWIM6SZS+5mV8qM2S
IRvUKSWOHgOcpBCzBI5kiBhA64oszgsD1/gD4VEET5UQBezLiKzTLJQpyFpdQtqdezpqIvcrjzep
aD57kgCZ95nJesLufpdic/rMPUTt+RXBfma1p/j7UBB3RrHQKdOC60i99k6JqZ5YnFzs/TjyrbO+
8PsCmvKI0XChZH9CJxv2ZcEOx98wtj9reMV2fiDMPiPf9AnRIEq9nJol7vIkxzY+uIL4LMgZz8AW
AnZkLgflLMQKwiZCcXPJ8wbw0ReEHn5ixNyNtmyBHGYT0jrSIhVLQUZocHPrWhc+ygw+G6Mrbja6
X+fLMkiTZhbKfFC3uxHFEjeFZu8ZmgLI04BXBz523/xP5jQk02wxfOs6/aePRx7TIODjrsJh7EBT
gb5t7pGhUuuriVJopYr3ceF56ViP5piUByy+VOabGSCF7HkBtyVDisRE6vZT4m5eX2AJoBSHPI6/
/M6aLsydUaF5sZq++SDuimg36dA68uva4iraK6JHopjp68JveL82kK/ffaGIslj6fvJqhBlUev2m
ZtLkAg2UnkfdHfpU59inqOMlO5YRBRwmFgYX8lAnpleI4wRB4Ivm1g3Frrd8S7bbI17IrRG/Z3LV
rHHFUeO8uY4CMuviNd7ZLKnvZFYfxSJOQ/vXnoVdm1bLZaNVr8uS1oEPiJX1r1KPLRlQ3DOIr+Wf
UrcpWS32Ei6rZjoajdyOPk19rNCCCei8TTz6lFWYc6vvP4nglrayVxyYAE/YbIbIvBEl5VaEEGqe
uhew2oba6VtPmfBoeQQjbxKggZMRLFa3R9ahqiNwvphZHv4AhS7JR7RBtGsHe3b0S6MeB/3D9Z+Y
izv7FjNnNSpppVGdw4edSAxMkilPkt8bbwal9iStUwsyDWEjoVxFCk8hGTiJ+HTCvXL2nPbeR+d5
qXvIbdMqoX637alza6WbczMf9wvHlnNRsUYCgU4/OcNcKS326/uTPVqR9Xe7NdSyWj1RSG1qvd+i
F2Ab08HehP/Pb3K+gm/YzFWRG3hH9GaNA2zDqXCwff4AuzqgBSAJtiVG9CpaYdpdjReY8UTF/5B9
XL/llq/vVZpFMoVDlOCD9mND5/mDrzeC+z5ZfgspntSJer1dzFcm8V4ox06kWk8FHIkLN3GA5Wcz
spVPr2+Kzpzt3C0DTv463Xc2BRBfb/GJzm8iRc35Ck2wRvZGJPJhxbJsRUb+eZZwICgb9QeX6KAB
Dp95Ru80gucjSwbz97FiTcic0YZsdB/pJD/MagUg5g+qhpcJlqBUKL6vA2LeioAr/yLvv7htBL2k
j2h1i30Pn8w4Uzl12CkkklO1RrvgvxIufAnelCd7GcAEH+4iIyXBdkcbFg/sDppVaRQqTFj4TN7v
c+6yjLcZmFSDGvN204XPVdvLQ+8hx3ZbEK3lcxC+Bhx+bc2IqV0pPi8FuUQ+YSYZv0obPv2YAFmI
S4umi74nm5RPZkJ2JkIpPI8KCeEudMmCg+UUTUots3yS7Y7OqYxzsro7uuh6I6VXGtHMLRr+QND7
usgLj/F/OV/SsaAcdZBJh3FJE6mbBXbFJfOQGRfhZz0lEwnu++/C9hNARRdZGbuAotIb6KKz0uJe
J1BrHiLFAnbgeSSZbtKpk+qbFATLa/B9ckdc505SOF53YFldGBlVP6gybKqTLdiyfPfhtF3L8Sam
8ZFgI4wN+7ALOMl4znqYX6Vm3SqEpdyYuccVZGcShNwkQciuJ5duDLvYSH1snFg6SWgG8N/GZzWj
/W7siBytVw8C/Z2gYDsN8QYsPY3aEd3neIa+mWKyR7NBvvvwk9ToKCo8Jh/0ZwBMHPDAAHFZFdwo
VEr/zHFYP67WzzmH/L+gGAWc/ea7QDz1ri68BJabKFzOGmDy+5+XE7pAv8BbLOUE7NyejoxrM18R
fc49HliOiQasONjquz5scDAVWVexVDMGJmIBUc861M3lHngUkAHTNAOS6ImiHCEYyqqRG54vRUWB
LeQZD51CPQud1tadEN1Vgg2Q7Vm0HKIYdcnMmbbDL+QcUFg0C2OvXbTYbntUbksMio9+FJtw3lCn
AkyRRBcGxyGr6XH7sTyHajFKKrdWSjyLh3Eo/RAl+9OpiqqF+M9SD0bz/W9YHXvpHqAVv1VRM0rw
q/qVN80whHXYZ55F614H5L3JvJhq/8m7alLiYjRAjkyJXwCZi1Gn0aM1SierPZuRbZUYxJcpANRe
WMtWo7AKkpv0LwPjVyuHF37vOd11iwjckpY4yMVyAtlN1EaV5FyBnHmMUwu2RiPj2Sh7HgiUuGD9
tWEPIaJxYm6kdfse5PpmmkiyX4SiB53c9rCV7RrkXEe9FDsV7iYYl/1crQis50y8sMvandfwa/V4
jp29DC8Rjh+nXLj654rKVtABHzp+Z4RVzEWoX4xAqlI5kmzGZE3vARmbstqN1X8CRcfWOGCSZY4F
F1dFwX3qdBThlZQtrXdqxTlN9lHHa14g8SGYLOYjFXxp8Sut+drM7Vy0HrbMVFD5HgdBTD1UUoJ8
jXG9K8TBWr51IuqIPm/4B9UhPBrcaf7F1wmqBUKSD5VulhUSLbIiEguvstDlZli2BjDOsLdaijqR
/Ah8/0s4/1ypHHJywF6So9W1Dmrm+Jvm3BUlL6YWwSsItYa8NDXqLCsaiNmOrR3sk/4Vu4ImB+zI
XZNNJ56OsQOWr1HlqRgLvctmjIk4077eC3c5hqONaLJpL0CmgayNBLoANySb6ooeUB42lBHzzyKF
ugKUdJyM7AxE35zr/3D3oRGjBZrCbXFNQ7h64n/HPHPpim2LSecE3BLZWvPOWsKjv9RX1tb52uHG
THCo/ZBjH6J7NafW+zVi7u0OCa2oLlXqbLu/PpO7zwDcqiqyHi9TM7N9Fs7PTMnliBwHdhxZICkk
Bbfm8k9vrYItMkCJmQR029jNmTOomrkODszFQfgFqjpK68rsMxVGfU7jn9xVASpoWmu++ZRWiLbf
IKsnTGCQ9dVEDGb/8n8HyWF0pkSo13Son2jA6POE6mq2uL+DF67xdSGQVmnkTXRLO15+zs2JfkJ/
q9uqZn2xS9bQGOyiB1hRDzjPlujDjeWUB8bwyBWnXraW6vQmEyfzW+ddBnOIVPpa0kaEUhuyW1LU
Y5Ji83/8m1vGDioB1eGIKxhru0h+uM45kSjPbd3mLYhf69Ux4xCr835WNisEJT+nWV9/hGVgCAyM
cqYTq5flCuE2+P5zpBYzdA6WbtciNndHeNIg6tsZuCxyJ4wvUM5ez/1+ImwZOhInPjdOcgkzKH5G
iLCw0UWcmX5oyf1fbhDE62A9S7+CXaHt1VVAERfS12K5rR38L9HvZJbkch7IaL1qwtcQkD2ZDiEy
fU0P9UhbsFcW1zyGFz9OlmofMejhRbrLs3hTDCTsnEqovPKoaEbtvVyYW8OljG2T0i8bpqJPIxdC
FbzEOSHCjNqH45/wObu6MXpYWm1P094OBBpQA4XQ1iit2HEM6IauG/UoGo4GWPaSiukzNm3uh8CK
AmHirNuG4wjjd0rOFihV+SWwN5/5gE4KP6HYEDy4HoyR9XBKjUvqVBHTz9PdWepbgVIu8yRraCWs
pZRZx+y3Qe/nj8OKAvpz6a4ZNlFDiznU/Z/X1EYZOyicdj2e5A0tQh6DbpszQKufqbCaOC8BzEbe
jzrDqdi7q2tUrBs02C3SoQQfCQYWzyr8WdPkhBNxHLzRQbH5k3PFE+NtCHpdvPyCSomscJlzMf6e
XORsBwLziwzh+P1d7hn6YNVoAlj55ii6sdBJWRSwXUAZrL/QjLH0ff21znNMutwwC2SYaokHXou/
Wtbv/lsiIVDzcRmQQVsIyK3+uw40vAy85KJWm0avAiph5n+6a71pUZAguAiA7HJKTTiLInXgD28e
SlcvaF239EHzyevasbZVPQK/OTzyOR31Tv+1RiUjD2BgZBewCjk8Y7mts0tpaClPjihwXLNURD+c
iiH0XhjGjxaRmEc/pt0REkxu9PJf6rgLEeid83Dly8AO3aa5VKSww66EMUZK9mAT5os/a1tt0N8d
Oo+DLoX5+AFpM9eQjgDu5eyUqEXDsFrnBHLHrDyOqNGTSuGvmr7UoVLIgKM5EBRJOKytA0K/vFl/
1gaXPz8V0WsmXSoRGpCPC8mOaOW2WwmbPNu9UFoU3KzWG0psMEEMf/k7UwizkVIKemSq7DZJpAMx
GU4RSl+e0tWtUW3ukYUz2Kn+qEyq/NmCS1wcZdppIJJ30cvt/PFFkg0rjLhiJtLZCua+iNflx5IU
pir7tNf5t1wM2xoD7NFMW0gNbpG7umtesxUtm9wUn02HJ+ypuAvMsXSoEhmLKFrgmDDUIpZGvT5q
6HB82bve/ar/qSrWHjtx8okh7fWYNPKs9u3sDeL8CdQGaCxo6rAl1VrEM8ZlYEjghDHF9ZcHGcm5
eKlMTTk/us6shruM2rcubMHPq5L4qDNLUsu6LkwdQzRIUbpRLUz48lpMTdDVLxumVEzZgCTdPVTa
BJWP0FHbhEGUQxBy9JdF65eQrjbXCXhhqzwPrkhaa/hVfzx46KeYNNXDOfHmh0Gau94Yb3fPKkjO
HEQF5unAaWWqZBqr/k6wnAgo1Mn6ODbljsYYe1W9lH9cGtyXeXQw3HYMd5ZEM6qwyPgkoIBD6+M1
hQGdiLTF+rLl/qALzc+KoP0ip64FSv7tGe0/IHS1je/sy65icIso61oFxtVhze/via6FUGReQCvx
9oZrIndZFx3zhtvPKdeb633IPnd7jK6bQ68dA/RmXx4COkpXUsNsJOtkUHuAVw+0NKAFw1q2NDvn
FpfFkVSwlShDOEhIzdW4RuEAz2AyeOPbl/glmVGvlT/w3qfHQtTFMt6een2BaNZdGYyWhAAnlQXU
Gw1VriDjeMDi7X8kui/DR/60M/7TLETsChweR8CeLjzzyG4/NBBE7mou8SjukHK4MSF+TicjwXoJ
sqzArepUBGm16QkaSV+x9S2fUyQz47h3gRs7+CAAHpcsRqOrleAcqC8ylwNLggV3en7vA1dyGk0A
EUz4tz+oBBpjsLnbG2R2ttuXuNwa8EZe6i35c4Cymv/3XKD3lnb2Qqo0I/x6CEKH5o0lWOQfHkgG
4P991ASUbfAqWPfNvqkXf+MkhHA0PkDo/AnRNOdUzawumdNKTo0AyDiv/5Uv8IyCEK71gge+Ne2W
8kiIbJQz5h/C4Ynbp/kl+3wdKLAlKzUWQz3fDHHXcDfJhl2DzDb38hf4iB2wFy9f33dsGS4sUKi9
9zkpfkpkZ+B3NZWiOKSiy9tlmZ1yIKjldN3IsyxTsPRHf+gVS31Cq8ybqi+++xG8ULrTcB9L9A2U
xW+5C1b8qwYqpmxBqtykDAo0mlVVWV6wzB6tP11clOw4KPqsyW0C7DV+QrxyyLDk/qlPqxL2IwDl
ymdyU60M+it59ia1sk6GV6Yvum0mkT8q/MFqyO4l5gzqsTqFHFaIjhehDvZy+cYVgRuveXMugQIu
B8C94mW2Mdp91D3GCA+WyDlF5c9uCj06b2TdSKPadtkhzaMoYnFIFYVLy2mKC5SbffaNLdZkGvJx
Woo5P2T8GIu9T73Cl/9AwQHLuB2kCFAalWRTb/xFSmGGLZsoTY9/HpKdS1IO349R25phkJws1y91
QZEq1kfJjgACC8EOYh3ZJRv7huwhRsP1+P3b4mnRh/IHFLT5v0RC5dfEys7vT3NrVnfhYiWaR6jm
QTIShe22bG3v+u0EIWAIAdW8sZkoxxK1edoldrmQyH+2zxldOydoqeHQgvhCRH6tc4g5DakNAqCK
3tqDJmdBgNmXPOShLkk50Nkqzt2BAr+ypi5qnvhK6LIVnIFLZLqNBs0Q0P3aC13qc+4k+W+9VUvp
LElxSk9Fs2QPDfYtzPmJmUqKaC8eEKbJf4hKYZsokfEr3+0fbFx77HmtdVTebJGYE9Zn9/0PlUFE
DVSmcAyoP3ADNKxpmiHF1WhtIKI8Agh64XDy2mfTYXwfv2ZQlnF5KokbaL01a5jA0J5FTW6rwhln
SOY2uu+ZjgUNN4gcea3jiJkmc/YTEiG8M/QUqAS/lAURP5u+cq96oJszHhMcmoJBcfoWBcFTnUR7
giOEaCaNc6n6nVLeNx9favjBxkZd+gY+DiRl7qMraoSc5kkpNR+u8haGir/4Otrh4OXYnPvs/N/4
+mS2sO8uqxqheRyWm6lxuPq7gbVtZhKp2tXkLua+WpfgZUNm0T+jAdg3sefMhkayHHm4BFKQlGp0
/kAptM62Cf/sW89sYQ51I8z0BnSHrgMdishw2F4mWZPKB8WtuRa/j+uirFJviEG//61Xj3YL7Jzu
8JNQyvvz+NmUhkpKLtwpOYvf7kacRFxZixFqBEcqhKHg4lqNuZIx4oUB6dpNG04p7IzP1ByIclEk
86xP9EpevE9H98tZYVaxbdawbUH+KFDMJQK2dQ1CAzh89mqMUhKxCU+mx1wEI2NliAq4XtcvBvWo
SeRh9PXwWWZREd7pnuZyYzj0UMAKssojg4X/0Gdkv8l4axMoUBWqDyu1i5/irxdUje6ZIG7pxtXd
5vWiFFC5jT9yzxPuj5MZhJ4qk2SnLXvR7oIQIHrJOO12bBqOKInQY2h9ZuAH8if358Vc/vzeVrsl
1shI+vbwCkyCf1Pp4/9bvnUDbq5elrEx3ANcK6Wh7odStO7VL1zhE7gsYzqIlOjrvNOoICqoN/jR
aXvWhb2/Pwiqq4eoeDpUQPscSRRElTlh6c18ZgVAw346W1mXPM2XfErAurUBpG5eF5BFtdbhEHMv
9FQvn3Y2duTtJzm4p0b7xbDjiYKESqixWxcRl003uwHXy3baeIbQPbxW/Vm43DKoQC+DzgYDVLfB
1w8UjHp0X1h4Tr8WxM3HCQWYvhoTClBsvfRyrT4TdACMdCCfn2Q19kalh6WHKYVTUvYOysTOIDXk
o88laNEEe9xIp/BLqBL5Y6BXjoPfKOhrbAwfO4wuEZsMUSAwauahOJi9SxbQGEOTzjeque58+LDO
YVpPtIzublxALCZWEc/k612YDqMYPdCCOEjJhGAQfmVemEUcB1R7qPtVlMC+Fs7P3NfSF/KRflWF
jhc45qoPeMDTZ+CxoW/gZcE/J3scow21dmJjxnKKmHVFQAckSx8se5icCsc3/El6Q4Plg0Kxqnmx
+sIGSdoyNpQhQMORsmQzDvaX7USQL+hRx5OKNBccB3D9o5wv0NpK6Ky7ggRl9gr6WBDem+WA8pFw
8DP/hRaGxLNWK0xUhTRul+iYDAHnj8JjfEW5f1YA4iKUUv8IwY0Gm/fsZKODZpUzeezV96+PsIbk
YyF0Vj7Uk+8Tft5V3DucUK5sK4j2zFMjmDxyD1vd+21hR0/af/6ucuRj7AZrqRTlAlCcBl6AQzrf
6UlT4FLzkuZLFbCEXeXgPhzI9kBzBJF8vCqaSGKp8tTdlqtqGDcveRfmoFaSe2pbojj2SKGwbvO3
qH0Okhpw4b2zguY+EknvG9u2ME8kzksTYd/iFLKtWpuIkoUXjfeN+Jh3BIWTuAYMC4ymCbmDHM6S
Z88K6Wjfom+tROQgxX+YdTsULRYDtxKkFq0VRIUZ8NlnVA9Sh4d9vRrFzKK4vNS4TkWPXr29aTiS
W+kkzFuqhzjm/bbBa4Bc+V1EprkptQo1cjpb0kBXi+80UJ1lSQ+X+XWNgowecprvz0uBYhRvG9VN
k+kl2LRYtXs+MowkpYY3UTNjKlanqMRj01W/266g3dUBD8ZT6TjGpd4i4zmixKx3Jsis7JrVLwNn
rWg3s4DefdV6AMXGx90sWVgJIk7eSNEcye/vsANPUbHwBQlsSI7wjzCo+EwzByNkZtxCYy0ShaeR
1M8EJuskxTckkTopl6WOXhhozN3m/1isutPx7umLVfIiyOE1eBN60+pa2dud/yAKK2kq4J4j10dV
qrpkYQkWQeFuC/F5GZIVvezuu8mgiM3X4OD4JMumRR2UU3xAJpCPPcmaFeqolup+cv9NEs+pQDJk
s7SFpM3C9AK5IfxoPpm22NvWSKSiqpyL4ZzN7U8L39XwtOnk8HqB2jzi0vOYNgrFF8f6eyIYyxmj
PWeiGnm/6RPpm9BblT74kr2k5X0FLRJF5yatD7MIst1/Lkg8N760yWUF0xe7vsf5NL9cuVfKguFm
7CT31b92BrtCjjvykajosRFwBIdWOFK21MJEEBFm2USbuJzGJYOSZTZB2Iabx7HaOT9RCv98bwzS
YeBxHzAO67XteJWIo+WZHXDUCNewqIHPszzSfPB+v0yqiK9RWzm7f1fBDh9qDZt9MY6DwM0qEKSY
Lxmp0BVZE4YVHt7z4iuBKS9tyCrivu8WK6FFgrrtCktPJjC1Zpr6mEr3AW4vT1pkSGEMqgQoSTrk
x3M3+9GfiFf6MrpEiKNqxHYYns9u1uPT9GzZZQKA0cgZcAj873WOpkX4IHu68THcTNqt0YqA6KbK
OQczhtO/52jwyCjzYJpSUkbpgHlfzRSuR7ZHGfZI1sF9b2LG98lKxbXa1+aCAZ/CgARxkR8uNKhA
EWU2q58BfwNEiHLnWrKDjQjo74xRu7UYVbeN0xumqp+mNiUhyMoGSg2itbNMyCuGi7OxJATPUHgQ
/afW19OrniRoAbTefwvPHHOvsTID0D6yTZcDI4vI6dFu2lGsecWCGZ4MTBFTqu+ReAfW2pAI80dR
M0W6dVejPWtJNTDEWUy9pIrFL2/h3vt0iBZ2t/XWWPlgDBwvSjisemfrAt/4qgIu7b1znCWgJVo8
7dDge9ROsDsOLHc9wk2jUXavTuB3nrOKF1MfNwMWXTQxEzgAwsH53mbMat3SImNUiJVBkBQK7VyF
IGFgogovgLrep5EZP/AWEGlYgTbGjyP+drP+4obyanz/8DUjUmfm4YCJQK8GQfyzYNsB/hOXs/ZS
ypL95vjPWlOrq/ZpsMF0zmQqnBScKEgnY1sVTMETZBPbsCMI5TSkxIcHk8cYcz0UKhmnGWmqAte1
vBExpOr698lh7m1gVifx5SPUsSR/Y95L9FbtuCzNtzlr3vUoYZWUaAynXyzEMJD29FK6CQwaJWHi
kzUqwE32KZe1Q38o0XsU20LDvfC+DPsOS3GTkvTZNrfxwmpQUmS8OIccNxVDCA0i1Ry/JnchBhRw
gNKnkHlTJJPJGcrTcBF04zjXklRPpvzkFF9BIuJ0Yt57LNPEhxNwTX0EzfvSswFkKP1tJSfVLmxO
hKqsBEdilGkqvokleWnAs8F7LWbEA9LR6ZNRcidf3rIK9cx7dZnAdHAZOoTMxcFb2pOJ09I7GpeC
v6U1lgYWdjTYjYRGrTvw7tx3T2DL9h12oL0T8LfyWdiccrDjIDUCJyMmyMjGkQnvAAuTINx2E7VV
1hUEYl+YCGXpFEYiwAfcKQcoeDYLq40YhKs592BaCUQl1ha3F7/zaWXlMy6hZ1L8SrRuzqCWw3Jy
C0lTKSenFi+xfU5Jcwf13yJaj1g8ID4HicwOU/qVw9nraaWfQgckgGw1899MfoVZNEAKfLNE3lt2
Z2NcDROpPpjDR6UIWUoUHFhsOhBifr4BTUqJvizvU/SvWtgV6MtOMZLNK6b4Ehn7LPGZ/5trSvJO
X3zFaVr36GSf9L2gsEkuIYUdinL8K9LD+uMlYVWyJ0ECtfbG7qLKXme0oM/viDmTDfzgNzZEoHaV
6YOQFIQgZiB6DXA2ppj3Jwh1uetsL5YiuTzljpe5tmPKn/9RMs2x7sM9+ky4ZIauBqGL2Q7a4kS5
xIp0JPppF2rsN3yhOF38OqMFGBa39mH3JxLusz8P0T/w9++SBHiDHbcXXea+Wev8DOrdmCjG4h+h
4M4rMnHAdaXuArQ8Ab6qXyFSta1HcjaUq4pOZ3Z48I6Psii2IFP2pLi4BIs5Lut37QH6iBcUWOqH
adUIbfVXacfM5k4mM0PdC8VjB1xEDnydrURWO9CLtbpl/gZKtO5GwUO5PYCMm7md99FM4wzr0rv6
dhM/9E03qcgtjpRlYIHUWTBDBkNXli8ZAokZuotkkgnFw0C76fBczNLbl2j94VnT84esa6fVBwvc
brXrtW6q6XeazisM04jOjj2yB0u+tEw+O5DoEyvlbnRafRKla167HUB2Z9TLEVzVg2JZxDReLp5Y
YM2xAb0U6UvTWWBt1p+fbzTWPeaV1WhZEadyfayoHSZznyPEuDYQR5w3drr8mTQ+p2Euuzv7iXTU
DReR2DbWDtGVdSw+8EcW5oimOLILmRmog+tPLvaOvAZPb7cPb0V0rb6p1f2Et0o3seyGE/drYhgi
+hjPgOotTROHqpjGcz1sbtE/GhW1SayqkjvqELPldfuEolHLwTzUWcWNrSOpUqaqlgqLnIrd901q
jal1aeN2uyQ1T3lS6HPjBhqkfYjY4gyKEcj3KrAfEeYk8fW8Nyr/ezxWQqgwGbdFuMhuL7Ex2gF+
pr+HMJFtCq9QLJCOW3JXQ+nk+JP5NImC9LX8zoTv062zmZ6IDmvtmacm9henOdlDInVIn0T1kE6E
OABcTSx/MCFqWHBtLxfVUCAJin8VUwQxMKBOmlVV5jgXUDOgUOmkJ0Jz3GxUqmUeHeWj9gQn82Dy
aqdfEknAlOUeMXwoerFU+OgcDAoZMXalIhgBbF8EKfZ/Ey9+TTrYjURcBiNFtOA9a2DS9yfby3Gi
bgXB131CXWudgp4xzyKXKsbguIINNX/ifXk4xo97RZ35ZXx2WH5XcPdf/osx0mqORjMgg6/n8rls
Ux/Uc16fkMbu5scudXD7Cr8gp3z/RThF7JO9y/W9fg0QGF9LGiON1Q4TJTFuiEV8QQfznyPkUYa7
goOXF3mkybasKsUiDlEMc+P9jNQGCnP+YoS4tPw2Bu/xKO8fb3c/69Wi4fReA7ILJr9xXTLfw4il
CEwzAOkHIL1D85X30j7OgnOyjGCKINtneFvw4gBKaT14FrrqzSMAlpgcOZONusiWi8jB+Cmx12uO
raWVs31qUv59I7dtl1M7kzmocksr+2d2mGSUGz0G1MicBhow+d7ZQ4L7nbqIaK9MkacBx5dGAgWU
YaLbtaKAy3bbYMfrnDbaC46/U1RSym4gXsZNwOukEtzRG2f2pheoj+stuaETonSmEQgEEgS13pNn
Ka5FT458m3rm13w7nKHgrk/Om2Q5RrqLKavCruVp2XIt26gD6qfzzPDX8FCE/zPQFZrKG+SDhXVd
wD1/cWC4EgoXan5dZtTV74KrMzp0tWgT2Eo9JXAl+sFfISkMsljKKv2YaTzUkjiq7135mrm6KFzo
L2kbSDqsnQ8YtPofj9uMZQ6D9Rdb0EJGr49PGssf3uFFjBeFJut7vQgeOaJ9b98Mf0LxEFg0fNNa
kNh+ul5ce13BALUArJbIWsE62wjoddiwZwLc9ZfzfAMiEMN1wN6wCV2jPH0Ffdq4fGDSDk0ZpdlH
uF1tbySExSQD+J3AGxd0w61b15LD5pOkx1Aya90gSRU8oGymzWmMLdyh3l+/t27tChx4y9RGbIyv
iAN9reugRZI035576lpndS3VzI9E9PuqX9nW9EjeXgpK86KW2foE/hriJhNWGf2CKzOmCPEKVCto
oX3/R+Rmq+I8Nk3laHqAuEbtKwYTGE1l6wLCc7v4cH0YrY/bqQL9jFxPvmkAQzV9T3MYL9SqSOai
1lrOBQdIpUcLtMPC4wpG6r3WhwOsHBC9AHSlIWDI1KfGY03vg0Yc33Z7dBTwj3o2qaiEMtTwawoW
75oeIRlkuACtv7FaJvr3UzooUD5/Y22zj84Oym4SoaYe6J3y0FPp91dc0WDw6sYFZgM9PPS1/aC8
tyjHZdEGL9JmY47qAzQtOh/YzWM5VmH4P3iAXnOn+HDw7eMWso5ewTRhS/Co+pukxZeaC9zMSQf4
DYdf4B6rllMhTJh0kOc4u1QC92wY3Le5iHBbuqOjichBFNZEc60WICaeehoSJac4jzOD7OwP1j2A
XQxK8TJe4GjckqKEwBut9Fd3qQsobPBrehANdRbWSKcJyiiWO01z403+baEnAOEUVJmJR8M1MUvd
Q+wsjJ5OAvQaGITE57dUQ8u+Bu3dnUAioybkeWm9qD+ckZ2ppiwCc5z9c+uol7W0c+vgI0rDHJya
AK8EGxpeYe7L2B0cNX1F0O03iTU25+kdCEX1enNa6s4xErXbCfryrZUpXgduBDgwXvDD+xofUmOO
r9SRoEQ7EVIIDlcPVDnJ6TsgjW4MrsV8Lj/wlVHFBhatxwA9uUDAzlvD6NG5t3N8vuT5pDZChpvJ
bgCigB/gTcEpPZMtqBtRSRBpFclz75hb784JLeMzrn841GO8PBc50fLLKaiClTv75oBgQ7iZnGDn
PEV2wUVnDgHHLHUtak7pupCNO7At2bUinES/u1DHAI/xYbRjB+i+xdfKjJJWdbY915Ewjfw/G71F
2CRiNFib+vbXdnBUsqeM6f2xA0+LYsJfG51xE9Mud+JpSEtT/1iAbqzWkaj4Gy2vNb7P1j9t9l00
f3Zk5T5h3hZ1fKfof2dDNYIM9b1It3G9/PptF9KGbdN7qzDMHIOC3Ti3Apdp2Fu5CFgbj1KPW0SJ
zgvQRgBGCH0d2xSBrw3rfRwvHNXkqgvL/XQj7+ppokOVw3VSKO7sE48BzWzxvd9/Yay8/rbVs5T3
VZvcKbMepUKYki+2E+5gG3V2Z02BW33OSSGApR/lgWGqcLHIEEIo4d5UQZDSFp8GUVdtripS9MHm
vlh6wNlPSAb2Xd3UavYp8zR9m2E2xiK9wGhUQYdwxgCuWplQwey9Fe5sEXbOvCdgS8Y9bqYyn4Ip
5kTEvbMT0GwiTaAJDaG+VWhqE5CbzWMjmu/1J/xigsNM7YCZUbvgLySqd/SgmpYVA5JIUIpUsZkV
5iaxMYxFyQ7yQpRH+T2FHc3mtiS2ltDvrvhvsDpTk5pi8XSjwO9sZ3AJsEvbX6W5S1yU4mQtgHxU
E784rmtexm1qjgxtCZ3X1gi1aj3xrtHxFxHPaPDhjv9fuH7eaPBsvp1MzqAmuCgavMdenzZyEOU2
B/Vdq0/v9typUuEq0DQO2F6yoNvC1xxgTS4YoRgFq4HaPRBuPpT38wyxrvChzsMNvZXGbxVNbi3h
PMXyZlooUFeJt58ggWMFvXbWQycpBHknQSr5eiJGAke63VEVGifrwbJjzLldRCvjJVHvbh4osxGR
ePSKiHO0UwCZmJn2pnT+6gOdh1ajNQ8qExiCkk6UCslalJTLpQV8PMwa2vTCN6SBv8hJOfSESlp5
EwBldZY7rZpS+38HxvtIQd0rd32qXlwUgiSbs9H36nqF4fH7cnkgXb3M1z216bZTxwC5c33vZ6z6
MaNaJFyPKLPpNbQwJN6/OW5y7wTl5zBcUJ/2oDEMRkrCeCHipoFxCpEiyHol8bUHG+f4y4KcBUsR
GY1zuuyvLA++G1fl9dTr4ZKKNwTe3GUBDGrt+ovlZsrNLscZXyjXJkivrrJIPKeMsHmxkyQrgEug
MUDb4RzARVnyZJrh50lGCfk0V19G4o4YKvX6iKf0x5iyZIGUYNTWxSVe4s7gIFR6jimpj4On9F3S
Qj3weQ4uUIj7HGdwAEOAlJpdPuQJ6XRYDhGmmHWIh04Dqi9Yq4v9eASTcUlEg285u9UuHANDLZ0o
coRpz7KsHoSrzNgNYwiduK3bMYEYLs/bboXLvfJU0b7w3WjTygx57tjJUxBXmKzdMZJndusYzzwJ
ig/TJbtCPAZzhnaTG86zKQ9mozlpm2jbu0k/zcaRe9W6+tPB2HUL+jTqp4fmL7uRxE6QLgnm6Oy4
lz5Zg5jCLblp4sKmT/guyUFaibMiKHbd8v+5SJFUmspIX4+t622xfweKK9o9Q59UQHPCymx2ygZu
cwZOjz1OIWyLWAPYmoHiFYxBjx5M72yay4BNCXtbxoyK41wcGjmbhe8I85m2do5lxLqUIe+nNgT1
eMhx0uT3eK44i5xNz0rx6ntXLz9/v9FhR3W/q5tOMSO041OqN4W2X1FFmiFutOQyG0UesGrU1moP
zIiI1O2XGa6+ranWXtcVX5yqX0l1yMzIZNGXh1VOF1+ImzkubYiV1AbgrupUqUqJpjNSJzSGWa5F
psZ0lrlAIm0hLqs7Jr+/aTd79M55MJFu2pRsJKbZVe8qxUpnffgZVvIqS7LP6XEyW7oY+Hpy0A6o
Ksclz9U1yQfoHZlGk1BtKVx4ZAT/vgyKVccVmTVbjMeeGqLMOQRu4o06FtHlD1PSI+iseRfkSz+7
ud38K0bkT5vahsdGVahr0/6TdF+1leqcvdnCYyu9+0uMHpN2I+nWiIfeK/K96XejwKx+UfLU6H16
ef6oinil8DA8q/2lvKLWLJH13/5KMp7MtlpAKgPvqw903KaniFfOWHtS1rx5l1rxiC1avBI/VcvC
DJwN2kO9BAZjVMZZczZkggwCUBBUi4zw/6YEDrNHJVCpmuwwptU/9DInYWKv7HrITDB7dpEEQLM/
lzJ2f3Zq5dpnWl3bZbo+ZBNKNTcPmqd2L1XDjoVwrQxEwdVvpdUa58IC1tTFewczIYT9U5/RAd3o
6yrFpNN5IrN4Bxx9G2kGB877w1ZH70Fl9esopEekoy0+Gab8iDEW8x7yRZGnUmAbUN5QX2XgNwgU
MqGBZMmH9lbEDqqNCewYzTm2C3+2oXpHgIdFlpbmJX3BZfnluCDeoCmcAi52AzmimEUUO3tXQRGS
WjUwd2vPaswqn80F6rsjPUQBedw54eHHNF2PJbWUgMx6+oi4qw1WGI5WHmSKRlWc3DHomJcmzvPJ
ln+rVKDT1Z4LwBUmFaInju6JBM5ftx8/oZkDqROOA6Q9QbCxl6QFlw7vDqYVVJ55CppTvBiZ6fIf
8OcEodU3gZhfht80Ax3dWpQ2eBW36/XQcCpANZqf0EwT7XZaxiLYFH9MG+wbB8RZYuSZK99aodES
IPY6VTm/hMvd8CytCdd/1VGlQsFWlLylSMt+Dj+1fB4Mj/eWfZqyNm+7Jdn5nJkK5Y52Ry0MXkFQ
vG9r7Dim6BQbHn+dmib0qwD8pqmta/QFJD41r065iPRWBHXZnzx52z9oa8JCZ3Mh156FbeQxKMF4
Vvi9U4wp03Qimz3fmNc1bfRTwLrSloHh3F+JEHC7igOu9iYjNCovqsMBGD4vSlVffc8kSQcJcord
YiaES6IcI1we8xgySVoZO/yXTkAQYH/GXDKiFIgHvozZzi2W/Gr8qDYK4o5uIsmvhbb04LeSGXoU
oEFMmwI98K8CU94eyWOQH7kxDMaX73Wv4msqaDAAWK9acmGJ9U6BqeRvvhY/ahsYKAo7P5D/e5jY
SvboezPIEQydRRhqQ1xq8EJdPMJen/LIVP+dg/nw6Anci4oTGyGuDkflTSQaeLEbEVlrsx5+c6k9
IgtYLr1jMD+TSMaQJzo4AsopohECv7atjIqJ4G8aNiCyeC76qQHoaBDYtj3VstedlOMW+4MN7+MZ
aDBbNCQ7UbrkwcSfuHMY1PRhhhakWaR7oizYfybLptIMClZTJk4Dscp0U4rOKAcMkl3toApB++1x
wzs4VEjQsv/UUvfS6Ci0ptaBvmlP9XyK6HAT3SJR1At44wYd0I/Mk5Xe9p3Wa1wNGCjNh4iwst1a
+D7OusvprrD9OIoeDGt+LOLNi2uL0Kdm3/lZHMDXoZKL9lzwfr1ygmtJ+tCaeFthKJu2cbIxJ+x1
5e6dwcXXQKNJtAi211Q915etxyUk8h6uQrEbVyGQFVIr0v4ztqmJS371ZcwiR2pu8nf+q609qa6S
p2z4AD/j2L07qpz2sCoEfiLhCr4gjtHhhaOnUh3kswdLiaqfIJofHIfEnIZOVFbK9mODqZBHXASz
EGJ6xIUThiDoYb1SM8RwWKnzxsxDlkKPGiQSdG50wfS1voaNLieWP5xCMgRmmntdcria6WebQ3Yl
JZFr0QxxtHPG15Bcw0ygnY9RpMq4qf12clL6sj8LrBIY2ura9/p3E4CwA38JxCS5VpLSOiUBqmhn
XVY9DFupG/FCjwdMWGMF9R3YztfqOjB2zmxE/NO9cgXKPSpNmsE7KbCpahGKJ4Wo0J8R6AqRmg9y
3tU/yPkv17ljktzb/rGN83qZen1LweyjQIVrEC5ODWuIHkw8jzYdt47U1zDzV+vgFDgjgrXRX+oU
abtXNuFRlbQ92rWrm0Op+iq9jS+9UFBM/rqjzdkPW5MeOi2wShg/6WImRp2MuhpxADhvh6z82qWk
pPS+2xqw7V3NfjTeqjxiUfzFWaf9g+QIH4wQHhmDSMtjstWAYseaMMx8CdyU5rjS3aiklBcrfRe/
U5n9VUq7Q18jLT1XhPYolPQF7WXehalU5YCQ1c3E+x+od8X5R3ZuNSDxwzEIvEhNSkU6FxirDDoW
akSP96r3KpAJp0gpEAWUebJfm3iVZppeujAfcwScbX4DR/XMqz0/0DlGkovOjcx3JaM6CI+tPhaw
V7fxgUzZ+0Y3pvSPxMopQP9MgAwDFKNT3TwMoZTktkYQo6AHz2HEksn6rIWUx/MkUY4bxWF6lRV1
1O47KUZV+I/N01ozYauv9H7knS7mT2LuoB6logFOEIKqElzE1ZFez06r3LNfhZs1gxWe/1utzM5v
RVlDZsUlkT5YpgDNYupwKBjOclfejhkHTyvAWuPWpLYm6y1E2og9nZn1794oHji2JxE5Vn6oI27w
5jOq8lxW4KJhxTgmd8dbXJC3N+XTE48RJBA7BsABp+Bia7hUw4cGmL0s2UayWLJuoSeVbMFjTjCQ
lp/QcpPBkh7TEShQsgqnjaKejbuxSLmxpfA3LFxr8485rn1MwibJoIMIbmh4obtf6vQtXVEOsiaM
UW4DukTSZ4YiKvxrMZ9kBmAi74mgoPD/PW5k1VJzibbpJ4A6S3O4R3VzSCc1d1iVair9bp/GG0pU
vdpxTieZ0uqJecsp24HT8FKIzHIQf6Cpib3uQc+Xts8fJIatDPDzw4JhLp52nRK7NjeO7Lmn8eRr
YNUvx9QkrXfCoItpKUCBiPSvdOIny0vI/WxelkhhWoTHzrCGP9bdv1blXsEQv0oEWUTY5BubQ9AL
DbW+474/GyS5Hvx5E9Ok0weyWCmY8fgT3niBvgA5sDykdVaA6Fs4YDjSbwsMMMMrij7bTyPgaSuO
blcGB0g4wNcJ+qHhknBRM2FbZAydOZ+Y4/DFoPLwEKSqBSKmoPc03xfw3SXuj0zEORhn+bLPoWgC
iqkdnNIZOvn7OciAq7hTNFV3UzlLs+y8/x5uuLVsSu3AOTJLxWslrdsfO2vfpentrjP+VzAu8//y
S7+Xd3KU9lFAa91AASyPEIG0BYqmjkEsdO5rhCvc4oMQWiQzXQ7cEba9EzRVzjBULUSrjqqv6dkp
soKAdIXOOuA3FX5jFZaXHU6lCe0LREdkmWS+c9JFYRR9Tyv+C7zpdIcXYFXUVl7PiMJj/ieNQR4q
9Wp4JWmVlHanEzv0qTeiy2/9QVRXtDyJwG5KoZuaQeBQX8Uznb4tyEV+N+B+5YrI1s2wJcxUL5E9
RfEZ3OavOHC3z6sXAb3p7zwn6mbwdyvwZvLHnMcBLHb9fxZGFI6Ov1rmL6Rsx5AavM5Flh+OIC3Y
42LcwnJLAWBy5gjZGROZk2raw+EbJZGvYS0QSFREYh6WHpf63ayw6m2xYy4D3kdxiu2iJkWkIDnR
RqBQq3juNEFBs8xp3UcW3enjLtiS9sgKIFGLw8OlOJpLn90axyEtedjpLldi/JyFo1tFdCIM4DcF
6GNwp6ZjFPHHVLuxvT2eyGtzrXnt5mWshMMMekSeylNmizBjmE0DYEymlrj8tpuOHz2ydKdFYkmh
phmoBymCZn/kdGTsVGFGEwHgOraWX/DQdYJBzOSSSWCBC/mbLRw0sqWxMgxZeK3ArcXRa2/bBDh/
OlLSSynsbTUh5gnUWGCILTXynxSHajd8r5nkYgBe9drlesbLexOiL3oknu2t858NQXPzaVSsLvYA
Pj72fBYYwz4dU7Gj0UxiIGYXPEIMM2LQj1Se0BzFQrMG/rToH+IuvkBoX8pHFNws1xotB3JuFoSw
7xXWL4K51nT7H70M5Zi/1oMaeB03qpsLtrUThMTY6QsRZLJRmdpp8tI2y9Z1SATU7mt7jWpdP53K
D539qPZFJAbh9BUS0Ml8KVabBDT/ZnipLgml7dxnvyLkd1Zf7SxtGLwfE4yqchufP2nOh87eDkcY
Mw/QYWk9xnWrTANq6SoRF1uHw0Bx5IL6GzMuE5t/tJw0QjOplb4RDK7Vjezdq96F+p7ovOQAMLeO
ETNCeHDbekzTkDaDT0jZbm3ZNgj7tLKmSK5TTIrOoc5yquNMjjspIm4I8ONpgN0LC7s0wpB7fl4/
wGTdTSA/9zalTGtzgzJBeLhua+yzYPh4Jsp3lq40ItcqAEpCZrR1CRY6UHa6NuOyGRI+APs+v1b7
Z3HkU8GTJk0JL9KMs+h3MyDhjfLKlU1nxNR2x26oXI140YcaCMBcodPq59T72hYc5ouaK2uQBClN
N8QzsLDxPLzGGR6ShtD622G+3I3MSKC18Fp3tvHaFyBEOwk9LpppQR5nbT6aHEtBoEQcGvwP7z8h
BKNogepAz+LWWA0ejVv6fDUqC6kdVorHWATkywnR1mtEOyMcDDRG74YboMqO86roNeivGM9qQcgl
e76sO5HfMywjm8QEb2NEfePw3dWpvq2sRL/OGcV66HXw3g9Tob/+0X7UoFZhzEM0JjL/TCMz/aB8
5asFrbtAd2Awus9dVJ2AZ4p3vXBq+19Hc4/L+ni2kA3qgfokwPvhYi+jpl0SC3DedxfDVlAcjmNn
ICvYpm7H4uHUQjne6+HrM+FFT0B1VMliOcf5t2mkUeoJEAxLCw/rlxrJ4b3Oo3v1Tm6Ty9lZb+Eq
HqPqG7J+br01tzQV5Vzj6KD1D8u4HpLM+S5g467rrh1wGk3ss6f9dd5aLfg+fmKuKM1FT0RhL8Qh
mja5GTz8CPMnVLK2Aoq+Q6z97m94YwsqYql1SuZttEA4W0bPIoYNIc9EvHP0X510oog5oS1N9uOu
2ZU8AMpHDOxy7Jg+BZUTAPqWLRKEi7NSDBgICq0b3aY447lBZEsp4pCT5T+JcK+VvMLPN/kPZCbh
mzfi43g6jFNFMZA5gcdqpklMVQx3FeUIDrLhQ+cmP/zz8rXQePAqGwb6LsHZXDYHwaqFde0fr1wr
pcSFiTqdG/Ruh9B6FnYzPlI8ZZnNh5Sk6wFwu2xFH74cbAskv0zkBi7urJX9KNg9Eizx/6OsFIn2
MJAgIhAMvzwHbyCpvd7Ud/fbsI+lzpKLK7ybA0Z+a/tTODXjTxDJHoXrSmi4dqo7v5iF0meS0MiF
+gKrTdYZGS0X7b8b0fJPGeVerCJuYCKQSWuIz04IYtp5NjkCFuo0JhPSjk0n6zXYhvX3lCV4xRjY
WoN7DliK5n5Xo8VUz6QMoUM2NfP7CI2HdmRT1l99PUU46PLu44CYCiIa5pPShXJHTC7z8c1eKNvR
F4K6lyBZb9RmUzliENjrL8EVl/Ap/2GhcXjKn/wtNWeSgs1K3W4YqCshnOx6cEMHmiwl6bx8CEUM
DIlqvAQKKc2MBu4/arky0xBZPID/MwKNnvW7UmFzV9vRd1lunocfITDgecU2fdA3YkB+aTXdUCRA
A4F6kWAkuOshxlz8AncIwKfYB5m73CJcGGrYCTA8x8/mlXr2uZEYO/wmr9GA5fYiWp/V2RttPH/L
bbIIc9J8FEodqaJYZZWajp4j14UGLmYO6jfpwvJvFlYaY3yW8iwv+AFuDNlc38dwJzX57xpIN8Dm
ZBucQ5mFQfXpIhh3M2Fai+HYRWzizaR2qp6uM2DWzCjyW0WJeTZuYqNjF0dXyb+I8x6VNGNcnOfD
kLQWLqjnZYZl6xfD/oLFLSMb/8fMoeuRO5badQMcRH3XM+i0sl7aDxEnyVfw1CnFrcSHYWfwVSZG
sx4JFgILraJ0qvsXyHxjoel/0fLwNVLXIQS/z1hi7Kn5IqkvdTvXDqEAf6Qas7ysQSiRv0Qr16Ap
BVbVn+BfSwV6r/DQ6aY6lN3d4Zs6AfTZj8zPcE0iaLFCztkShMFw1+geB2rFjWLb7Lhc/uln3Sl1
5oEFtCSYWsoEMoWD5YNZ5S0t+pFLzFXrTinlFk8WVxhhS0QmOYUEYY6JHohQUcKUWib4D/rkEnnY
HBvEx0912ETsxj5GNKKfk83auNANJiNmRZ2LAAGxGPwvYr2KWsPzpSxhO+eAmUXY1LHXaGsHRc/Q
dl7+KNCKkrVvwecqUhOhUi4dirpwyElLvW1CeM9HpyU7JepPpdxiVvduL2QnB0zHhJKn/QOM0EOF
7/5jgfbR+ejc3z5Pm4Cjp2Of7j6m6r2z0+akbtdbmfx7ICAfQT6q3KFHshQdCQS9OXNXTyAEvmNp
KbUGHojcgqbFkEHc/YzckoH7vI7cX9zwolGJiYxME3OABnjMowocw0OR2J+a0cs/0K+QAwrdDsbF
1/5BALS4rghdFtbExxqHa4qWKLrIx3vnt6f6Hlh8DC0U6BS+eJY036TJldAtKCA3EBedX62eHmeH
8bJ5nAN48O11bRiIT9rE10TdDl0z8uD3AkMwnCQw41RPp/z5iumTh5nCrueeSx+bpuEhgj7yuF6Z
3n4qS+/B/7PF/T2nX8oJHJ08ppLW+8wIlrbFFHIoPiz/r3r/UC8DxFBaPJttl/o+jnBQREsPZhdn
X/Bn89OhOTB6v6AhuJkrELOToPzoOVaCYgvM29FkrJ54OV5TDrwxVYfrrEBhscGPCgkPbrJMIEA+
u91K0nzSUOOfrurxXqiWziSl2VBvcWuh5KOILKBXI40WSXbcNyvBd4jRNmlLMUGvr+L7rScU7b86
ZRecPXI9lflR0+EZzD01mIzNqKSBpuNuBVf9xJ9s8cjnq9dELoIkiRhx7z6ADbCI+cBlFtgu6WXt
jD34CKYBSweSo9UvDmTz6oJ6U7g2fTlaGzQqt359d0gB7aLnUSkyXJ8to7Lsl1k+7CkIB1mpXEHP
8ySixI32DvaKcDrXR6bHsTYhi6phtITyWOcebHi6davN9pFt1EhKoStMxEW1Pe485/67TCfP/HG4
5nQDNbIjDNL5t/cI143FMh2S1bR311RXzyDtng+tHD4LGX0lAN3E00RHmrVyNapiaFKzpZYPq5OF
UKf1SwZyIUhWm2wCy1fwMuKtbvVvSIgTV1bvhYD9LqQkOt68Rq6US6gfmfFMwMbgZMZFKIwmuj/m
Pz5sAYEjoK1idS5piCd6nfHGC0SRBAT+uHp8J4DD/B0JXFcOvB3KXvPMFBp8AZKy+iCoWZkuWw80
nV8vsdT9Rz9vfJHJ5c6KFFWqwVI8gH37qsdNB0mcQwVfqTzhu23Ta80JqZGP/CmFINfuZfufVarq
7kh+5jmhMugI8kL7nunszVB+Pndi2s0kO10D0H5/P9Jv0/cAos56lxt5b11y63N+2Va2/3bAZbVW
SxruqmUFPiiB5cXpLIg9x6DcTFsfSgmTtIl+pydtkS29uUE6uFYhBRynlHIa7uQJiGOdGefWGD3g
01bpxJ0hyR9XLJELyVMEm7PUTtinRGYco58lCOTyKikQmaw5LbZpcyEkBVDJNlu61h4QJFg97b3j
Ou/LpSVq/i0fMTe/g5jv++2OxViEGdiWKgUH2jyhMsUOjEpxHgunlg/NlcI+Pz1S8mo+dtExOtBo
m1Ij1nHmr++Vvg0obCQbEWTz5BhoMyEvlU4t53RsT3dfT5AK3XOvTmxKIUFbYEW7QLpYbzaqn8H9
F0boBdRlAFKxAwnhCYnm+QdbYHE4WjT1dldViMyNQEQfLwZY37y7NRM/nV/MFWx6oiw3hYfxjjSC
XfzK+FGI+SfpwIf/YzTDM5sGx4/C0CKyML6vKES5cMc8JixiNIKyeZ806Qsf/+siRRaRLzWLL6nJ
yKkS1SYvQ1KW8j8/JPYYxJABW21z2n3ucabzelW98GGFW2MwvK5lCzg2a5gFHLiM4pAMpFcRKgR3
b6U63tNaE2zmkYj5tGjO+2JSZCnX8/4YP5gkjKqPKiJ6uk0mjP/Rzr1NryynoF09F2OojaEuZy8A
8MYBWFQ6UFJXTbtXVdeHeI6j144BKwQka1+PV9T8Ri7WxcLUKQHDXQ7OzCXDdQtlOTx+Wqi5Rh2p
EZRF3MZMTdfaAHwHaxIICwrlKqAJkGgZgSX/zxFf8iE+D9e0M25rh5DevyZnX/tkTi1i06W8ZuzO
2h85cVqLlqv/uJiKIz4Z10mG7yR6ugl+PTtlnzxv/bikj4XKDilwGokZLT9eqgh1B2S3Drwx6QWc
956VJYQu3wNT8365qhlAcbhN+wakowNk98knQVTpNsNNRQ/IBhsp7bfLh1VtJFw+Bu3zCS79hzG/
PjiTWicYFuB5+pYkKhKjQ/Uy8IJpOYSqLBc0xmZI6Rk2vOvoPCTMv2a0CmPXzFA5M1Sh3mfChkzx
WPB+L09ozT8lB6d+kliDox10wDYGK4LqLsakt0ZfD+u2vnw4FA+PRuliXuo3CGA+HLOK/O2Ri6FW
SbkbDzuDqugun5x8o9hJKabyf6vs5T4koHaneUMcUyNaoq1FzikVTq7Y2X67fGAqhFsJF5ju30bJ
cKybLmJeyBMF83MQ+onTUzBToep8j9MqHVKIXcDsyvM0PAp+1lHrk3fKGwS3C+Bhv9+gWEGOXZQ5
jZ8Kw9wYVUQmC0ksT4NwtbfwHYcnc5nboAYTcJ66ayfR0rNhw2uodYkz7/GTw1zR04h2sb9bbB1l
clszDkiufvcBRPSQ6DhPU2Pru2SF8COW96hUlLOqjUWOwEOpM/yqAxJoWVwR/jDd3A0cc8OVDXeE
dI13l5CC0nAIeTGwGV/tZW5zDglAKje1NsWazTfEzkpak33PMy0JgyDg806OZ3O/cyHSi8V03m+N
YijzJ8gej34vvE/yzOg7ZS6O+272dudEnfs7VifqH498up8KLdVCMn8TYx/GZElWiw0IT9hfETnW
cpZZ8TMhDu+rqZOttISSuStY7HsZB9Jsub1n7KPAaRc5XEy9ZFQonIh2FkRTE7gUuYrs1ebZmALJ
DDL8TpWiJ47yX7FjwEEdfaY4oBSohcwKRrAMJyMtTarQ646h7WGBUxu1tC7AE9AgiUHnD6PAFVWy
0bFkVxCQ4H+wXnPzW565R+cNdc+TEmfcnfxHQHGPMlphEe0f30eghiReS1YExw8GyPjyboZNUPQO
qPapqKqoooEqkr8fq7SwbKbwiA0T/DKtaIAfiM39na+BT5z30OLpXNSuXQgxiB0435WI3zcWFd5Z
Z7k8jTueYaMu8ciRpj/fKcHTAmZ2By2HNv8Ye9opP2Bnu2qijWFVdvoqzf0Y83rtQ6X9O/LPsdl5
ZJZGaQExebGlP4vXwBEvxtfPU9nbDfHXSbbCr5drv/kKCoXZM2IeXC8HTmO3mOL8IGK0hJKv0Jje
U7FMjehF2YYI0FX1ZYFVv9AQmiCb+7qCKcFhVz8KwQK7gDtu1AOO476Lt7VpWlOBnH/txux3xaBt
q24nnQDOf92DRm5kcVnFJl923g18TaOYd0VKHqtxAKT4x6JBzKJuz4SPFLeqmVpO5//PMAINQMhP
WNmyNDj1nNahPnqfkGd9DiWtozfI4EazFp7N9rU+FF+s98Tq8nVilNAgHDqstPRmpKdCZlGLN8DJ
Qp5nqEE9RBS4UL8f0L6sTrnPqBONU8lw3GQc4nrkRDLeyv1X/spb/DKL5Dgk9gVbhhkS5rhf8dqc
vKkNe4CYebw8l8oTTmXcsLWbtQISJ49REF3HzS/yIXBn/qu0eUCivXviY2ppMhjvxBsii0zlgx+V
77WqrcXcqcviSQ5xG1MwEGt7sW38eI8JFu4Doe0X9elHXRVnfU8dqSUtuUJOYSIUMA7GhrudrPKV
qUolfqWMMIvM2qJCbdhSvzXJZAgAHAhxpn4kujQfQ/YIxC9WP3W+sR2t0IcXt/KIYraqpKnr3jOp
ikNInnCAvki7cTEpNxtJvHUkmRS/Af5NXCLPLHrmK+M2/YV/C3DkA4BQVc/nR+9eGiACxOhT55MM
bbADFzz1j2zeXKuxEXMHkWyHwAi8vjem2xDwoEJq+pa/h1Puoh9qizPY28Obd/Fli1GonKE5ZT9r
FdQuMxJYars1bTChIDOIizV6Hfcycq/8FK4tGniddpV1snIqA6OtZmC56uwOSUgGPbzJ+zAx51Bp
PxPnkYTJ79RZWJnxGXP3DOuD130rymrSvJdJFXdPctvIFyKtv39Wjm/Y1SgL0wjS2s9rXVb5/4lr
9TwIk7wxU/sWbSIbSviU3OYgmRJPNlgIziKO5sTUoSv4CV9SDuKmIlaijeteZDZH4Ls+yLnQl5D1
vv8a5fNeWl0yviPK9/K/ZiUyWVeaKtWs99UwxJ7obNDp7XvDXvCgwd1xbYWyJ4qJWhi/ofEQqGNV
9ciZFQUCR4hhGSOQbwiWtGmaJAfAWd+d95Fjp9d7zU2nylEsh9T9gNUumUWr7mo3qYsKwIRg+MJh
BOGS9R7uO/76fr6pjlK50y+UxLBXPhB5kckBwXTfXTLbdHbDnoAkpaDTLnsMTZMBneba6ud8pD6o
phrAblD7q/ZRYKiRK15xW6zdqPYjse0ZPCc/+YWPdFs4q8ktaQ2o4OFuJkpvjhQmfp6gyygc0ptC
qGUEmiOYoybSIDRxmeAI2twzYeksNwMQjzCzpGjTlD3eFc5lkjisJPuup0Fpu0m5247g82vM3+21
BbFVkoZPQCid422vUh3P/hBuIJ4E8DyDwNWIVoGwbMVKcXfo1N3+P1mWlt70fTmsu52UqC4/mwbx
incBoanGzeeTCQUoKi2MkETbb4n0PjVLYvIVYqwmrdyjNV2xNWRUnhrAYkur8rnjyCQmhbJoYiiZ
zUfIPV75RGBKEFls7A74EcA+MFqLYlUiGmZE3cakl2TFG1GrRFCVFiRFIBKBlhJmAH1OZQU8aw4i
MMyY0M39++ksYFJy9K8bmXZOAXfACZNLEcAltFgRCxbNkDx78EJtSJ0ru2nQOoOfuvIIGujf12BG
9x7bS9Ho7TiZ3O+YqREWRmaaGCNmdfzteVqhn0wcFod97ls1uuv2eVmU/aSglVIlojab0SOAyvDP
CH2vLdV9nJpCuUKzVqgLYkYk7ziDeecvs4+JHaDmKibfSJjDePKV4ghNj8byDT/IY0mbfRpyRCB+
QBpJtb/xVNPZkDCE3UWUtSEf8ZO/aaQoOIXsdi2VWMz2YSZDHuhUnDkfcKQFZ6+LFn3Vs838KWkL
wMomwKFOd5lNMb8efZefWmfG3Fn0iKROnUDWw60HUHcuYAnaNeG3mEg695Wbg+7uTPhp2n9Mawp1
hfusC3qN00ZiLnIbx7TqjZ6dfXASncIbAIYP74yyV9gd14nOKKC/NKqMMkNEZclLHhD33FaQIvvk
eQH8/5z1bOq/Xj6Uvjc6vLinW9bJ2y3ZhPROji/OW8zpQhHCXjknOSDjPIFgAvXtgGPKfpZH66oL
DIeic3xi5/52amZEfIFhkW2YCI0+zTkm38SAqt5Nxhn/erzUlKuWoJ9uqUCnoOFA446Rih8g7vJD
gumJhVFMy2Jrrao+ALY25jyF864ijzgQmwn/imJvb5AMBPjF905AK8oW1oxedyBOgJrJVYrUvWOn
OQVL2ilMSQB81j9OI4QOpQNWTIbFdplK4JIf9hrCViDstCxpJnSddEXwAYBbB3DGJMXKXLIYTfSO
Fx1bjDliQTvooaCl4wjsLy0+Oy7fA/v46tszLc9Sb8sS1/Uhw4gKJowAEzgijUTaLZrCdJowaVOA
w90Bi96ZLvo+1a7EjI/2S4VLnljgAO1S5IOTrGHu8NVUNXILrehtqaSGH2iZLfbCXqsXjcMKFvkX
y0j9zm/qYD30e1uQ0G+9EleGF1B1qXg9NrrkNURq0CQCp7xnTB6IBaBlR6PrJAw3ZdDXQbGhtKEZ
3i1KHh4i3SzbI+Nn4lpHhhKEBipFhYcqCVFM0IkAooZX1ZqzuBVM6bfLyxbEfiZ8Fho76wM8F1WY
KnhKBDYIVv8XZUfFCBRVV5JdgQftlYu1QxpUPkY44OY3sDWTbDXSRfOaAYvC17zfvuOzmUS/wPa8
FRiQ02wujvqUGcZz27Ff0s16srhC544TzToxDUvFYJ9Rj1yf2w8zuK0QgA36Fcwx66U0VPpGHrlt
zMzk7ydF6U2QG7TYLOXC683Kl9uXOIZDD0yRjUNG5Y4hRmjBLwKLiCK3xmg9m9ALR7vCF7X2tnZx
4+qw1nA6kzNQNVk/IFWN6rUBLTTDqHKcKNoPle6Kos2/9FyWNQky74jjPjX/xH5XI1iCGn8aCFgg
2frr+Em5rrvCNvr+VrvlD7S2ZOLeKaCRHF4Q/X/rFhSTRY+X90UjumuXB84LOxo8X8o2QDVCjvLm
XlwnZEe8Dps0/Gt8Ax6pUq7+8SVuDCNaW3eTrJ/qKK1k6tfqGBlQO/Mg4SFk/jT3PIFMbRE7He6S
6+3bkrdttwV7n0W79gaM59I6rtkJtslT3j/6neCVAquCMy5jzNZ7DYykh5v0pqRrIpVX4MYjmJda
Uy3vVb8OeabI4RR8RoAQHPD4KGYF03lhyal0orrYvr9xEhNFt7g/wyOrnTzk3W0uN+ITscB9Rjm4
FWXhwTXtYRsQIGkeAB4B3K57EnrQrqzTEDUoNcZCQZJGHgyDD4dvtnm7oAkAC7/fWABymPbMN0MV
Q84gyJNUIsACy0EdsTixmlR29x8HDJGJtS1OqvKfjjdo5D4oferroozPJjBcsuW/OkbLXFlN/lOD
ynigjC/FkYDqnsC4Q3pABHjoQJU8Med/91GdfCZt6O8Ql9NpiGiKyLMAGrPth+ZwLQJcbVyRgvFP
ZGFvFWqoJcSjo+gA9uhYdIPk4f0iYNfnmb0YncpK9ysMcI/ES7VZZxiO//0eguieL2EIt4MZcIEr
j/MUdYvmVd82fx/F9/Ncf244xTeCXwYnbOa+2GNFReLaLrfrmHfjY5SCd8E6rhJFshLJkzPf79fR
uVW67oanV9iMDd9gR/lFpQATMIDCVd3IspzFGej0SZYrc4IF+uZba4R9IV6JON0Y+aHJV9IiQAwU
9143zzdnRmIiyAmQVQhEzwT8RRTvT1G8y4eMgU2zzaRyEwosRNNy/o+THgrebBSSoHke66Ubd4an
AA+smfFaBl5wWja8fyENh2bgRSk6qeYzUQYQE9PGZNqN9SJpLiVoHfn0q02rjD9wectXQCATDadf
4DWKley08GHtyhFxR45SSsE7SI3iEpVo7cx4Pzk3cvcRC1AeYjEHuau8+nxJPKgGNBUJOPGVicW/
57iZHvX8taj9p111pusE64MP72NPep9tIfSzYXJgM/OgqT2KnjjepCNEW6gOGtt4Ueaq07Ar8sO/
ST6X0k1c8PN8+w+jpxo2as296hpQcVkvt2eE/2+SAfmijjU4h0yd0+rp4KLzugLw4HP+IwftQaHA
zRlmXur4i0YVldExjLse8H6kgDrh5/m23Dxh4cL+5tUCOSEqgbWnNNjemm7EizGN0HKzlPWKpY8m
RM6t91wrtmgllOSrPPGracYhnMvW1vqd2W8sjTMtvCwSGSsr1tSpAZGMO7uD/kkgBl/lImtonsud
ccO0ZXVtbxqdFKMbrP7BQGms8VHnjBJmoVoKCq5oZAMp8PCxS0+6W2dqERO2Ppo2uEJeJ6ocoSn8
LMsaH34hDU4z196x18LMRPgUnCHSMvQymWvLkhz8DQ48wHSBpnUYyrAJuKPhgBgDCjyTcJK4NpBf
sCtDhuKGDepV5XJsiJld2oZfBfh2pjKcDoajTb41Mjytk3lxc7mwA/a79NRId9Sjw7RWqn1c3h4+
JkVV3uBJdmob/PF1z251nbz9V00b1SAfq3E4bI2Foy/kZ3X/2IuVMsfuMyumQSEJzrGXjJtPlZM+
K/9+7Wp4wP0iXxuL+lcWUtMC/Td1zYXEZMX5lBPY7xCnk+WyYVtz8YkQUO/WF8fVGjkm1uFjmK86
eUm/+0s8/ai7z3fDtVwQaJDwc/eOD+muyd2pVsClqDJE4u1rjoyBi7a74r364eKpJAIbE1qqyw4T
Y2ZlTavcVjGNLaCt4AMNEzbgdmjGJbSNH5CePjhswqS4q7TAfVvjRBu+1qQOrdY1iD0qCkCSTZfX
30ILno1qAjw+vKdoobFDe5jmXJrdYCLmyqupFq5SvVvpozrF5XXR80j2RYEy+uDFAD5ZdrBDrwRq
D/9v3v2ayTKqMB0vCb66c4+x+UeQrcUZmgt6TKc33W1Xn7mWE3ZXF4y6+yo+QCfEVBW/T2dYelfi
4hLHls0jhHHjBoPVVF1ZCglgqAey3wVAqjapo4KO7yEg1gsLbsMQrDZU9zDmWyLiy/k8+4/ydViA
qCEdBPz0U+SXi/lPVBF13ve7mKnodH8eqn8IgG4fXo/1u5haVnQMoOwuitDcg9p9l7WhehDfYpic
HACT0a/wyezEGXmhXv97WeLSWo0MKO+JWCojwRGC5dW2WX8yrgxZYo2Vk/8Pmyhc0WyeLSJkdVFb
Az4IHXqqpiJSDDg8ygRfEFpuD91/1GpFgJZA19Im2r6PmczpvkgKF9Crl3YPrE+hxccv2TbdbBq3
AXZSqpdqH52BCOXbetDltltmkqpve1uImlnowL038TrqjKpovu/jCai50eQaJcBEqm9alY/9r/jd
8KsHx/7a1q9F68AQxjs86N7+++AecWsy34kM93696zypw4R4FVp8amYaO3iNFy+mcN8YBIvZRqV5
8QezaDmVG91yGYlzabgLYT7tR+Kz02TZHF1fe+wcoPPBJYHTj0u7qb0w3txsf59h+hIY4FkWLNSX
ySQIc03+7xr9i4uKOTiLBYXaW84gHA+HaKKUbiOE5w9K2ZzMYPoXppAhsfgBPn5oyl4pmt3KerHL
ylp9djTBoXF1jJ4uborzCIIR+8xW5mBPlw9kZObHpj+w+ZWxOf+ODpdoDL0CTu6RctwvmcQxD6ve
B+CjtuhECbtWYREYQIozeD5r17hZO+V0HEKy2cEgCZoDNm0H2jrwWVFgMJ1rzzsS5Lr7QEwKM72N
n+d3wbPI6qxB6lvMec7kScX8s+NYIaPzH9IEkfIZX7nzlWte7ZP8PhlHWM0JGol+DniIeUq77QYL
KfdFHWhTe/6I9hAZ1u1jVzT1ZprN4kQdfxdr4o99e79U8TtShzq8rSkWS02mo6lez4JP5MHVceBV
Pwug+0ddxauhCU4bNJJ9kepXFTUmBXkJbJgJpmhc0rv8TjK0jjN1Sg3ZMV4hw7E1K7U7A5H79fMm
mVhQVsa4oDTHG/QnYGe/71DJY8IJb/hYyOOiiKD7jPbefkWoE9/3xdiO3u3pPjpUrGA58V5IGTN5
j40BztftHRodM+1GPlAy0UYdTubOPIX7f7gPX3Lz8+1iioc7/NYnl1cBmc16dKwznYls9h2avmh3
vQMIgx8Xo1Ns8xJSdFME1KYw4LGG1DHF8qcoWswP3duMNgi3NQfIdTpvYHpej6f0PkdusLxBlNHi
TLIZiKrXuyTri+hfZT9y2lwxEgJ81SmFI8mS+AjpbNRkFRMprFXhJzt4LcWGrPaLy+gKb0CKwxZd
Pm/IdJ06jKcPLXwmqyBIraz3Spha14Y7lIBKcFu//14m/xv9B6mMnSbYA+jTMDb3Clu0eRGFG5Su
We89cKGbXmHHv66aRBY6iQ5dPemttD4LhsGvXzIsSERs8rBZDFTA76dy5Nw0muPlfF5avVOrgtcJ
FEYvaU+R4AVgVv+wT69yWQI98W2Tfjc09YiX4ue/b/Qu4LAywfHOYkezkDqeGCox4+MOj03LJmvm
dubnTeprq90JBrP89UCTmt+JjXmvHOErHdR90H9qnvn33EOn58CWxwqm/Llqn6gW0bTsU/YXKTqn
G+cDCQOObYLaKhGIgCkNdwijwfVsiDoLYlSzYv/P+wvOGSTsXhGpq2af5bqCZi57OdAgme9zahz6
Sy5A5WCYV+QKwZL/hzH9eqY4IqVNzEBVPguzqkGXjk4TOSv0pXgdbfg6agEY6K9OTJJThFOVlmtR
GSNCFrzCUVbPoRjZdYfPCLO7oEM1vj4BsT7Q0fuGeNZYCer6R+G1+QLHtNbEbUbLgyRh82Ezg2vH
KirwscTuVypwkDL3xjeYlqOI7ow9rQrCE/PZgIJ+/yteanqVu2Ld6AG3AFqNu28mEJisekYlSFtF
2J48d1AGWshph6Tdwc/iEYFowIac2qNHsj9viwjgOt/QEIxRnQxpVJjAr4P7P6Ol/3N0vOWQkHQq
8QDFsVB2uV8ZvQvIN7hzbssgclIvxcK1cl3DbrWIskNiLybucDLPF+4aHHyqk2KjhlcIur4SU8+E
nSKZFCEI8Y7lB5DMzUMh0YCahkIezgOjEnGUaf9QHBBbCV/S0mYX1r/uEtRZewG5pV1HW9DwIf0/
m+FLizsS4YVBOTeepxN9D2DU8T9IizymrJqSF7y0rB9vHVxL8QEpyFt2BaozZu6Ov/oAYd+JQbgy
O2qy08vrkZ9B0RCthK6X+tPF9ds7IcrR3ZigbX4k5jpm84WfM93/Sby97HDpTeOLJ+dHmyQnOk2p
BYWcT9EJhAWwGhiSErvv6Zcz5bQ09hN+h7EAtGXf6Qd05a035Ohg/TwiKZItpDOV8aGPg6JWnhJl
UqdLVjkmLHpkG8y68j3qU1UhQK5aFMhpThzATGfzQrVcXM6uw0c7AADoqGvvcgnG+2bWqFv7cese
t2zxRzhFyzKlHuRGSh9lcnxzhPLFlHvFQn8oqSVfF5K2uHR1xaI6S9XaxJFJ/cObTJVu9LpXjc1n
d6MXEQOqyyi5fyuSemIUPkzTAUt6S3XfLQmtca2iUzjHfHRZIjuxeoRDOW55V67V8Yw7tMsRm2Oj
XfcExLVraYPsuWKvv+UZde/lJ7RmUSMWQBKaCmjFtX3ntSh0vvS6AgzLCKGaUhCW8WVlHfvoje5Q
oNhs70EcZIwnXiulZhAftNogT5qDW2uXik7tMfn7ekc+4dfQ1aO/LZ3IUtEDtEXm4ARLScXYXcsU
kVQvtbzgnJQCew4gtM1mxS9dL1VRYZ2N4VYi3pie1P+KbrGM5e0Lj4m3P22UgiSLgjojEQU8FLkr
R3kRnlpnekpebKDqA5Mu65AO3PEdrZfxfCmde1AJs56ZGoRePQT7hm5nScYjeqpkb6m4YLK2yGUC
pmWUmKbN/1ymP7Wxbett1kImuasRowIDvd+G1NbrCVA2OpBr3ZAhV0yPbvPz87D20zWSNx7ENVkn
3U0pAbeV6UBWzL8kGaCBQF7MwGHcX/YDQw1sHaQZp1IEE1rgTUOJ2Rz9ag/STTTOghbYSi4coZbr
2uDQUL/IYnUFN2nL1Fl7rCnnN/au7Fp16pklcvYDElATZDWfby5+1CkpEr3mgvScwlVF8OB2U3LF
w9d+Pu2WRKOn3L72iVLLMD4T772P4/k9P5GKcCRaRBGb0H7Di3c9PQ8XDP5lJdyrZFhaL8QID3qL
IknRfhEyFBRJTquxE5EbdcT4FbARGt/69t5qBG/KdIIoiGoyYMzZL7jLN5K5l3OMeLAwymzpwe3l
OngngcIyML+9PyKs0EYyGoDF0c7ZB26ic8gNY7bnuHl2xOq8WFiqk/7nVSQJxNL6gdT5JqKR2HIV
gLXatndkXCOAWzaUlJVWWS5rVtsZ6L8HM5E+Hr4ZsNH0VDksbYKhTBovTqW2GAdDSljUUgGf2Uke
EoQfsIuQs4dfw3jJOGJCLj+iTues7xLUUWhyXHhZtFWUM0kiat8eaDvaDzvsoOvmwFQkfaBdD3nW
R81bg6INOw7mKk5OfKPeF7T+M9ktj2bsUHrnpimf9NR1WBZMUlbuRNzp0kplL+A9F7kM5XJBARpk
7VOkH3XBgU3RcMsQEDVYGblxDZJj7JauxXceFGH7/4OzT8q5OLa09/fiK1ImqPahDYNcfjJzixDJ
aBvWUL6Oki3F0RvCbdL2P4UJ9MiwMlx3DMLilEoGhyhY9ySXC4Gu02cuGQuvq+YNT4NoTuTQlt5X
YcwT9uINRes7bkx48DS3fjjvrH0+yT/2Zp6AMIbUGkiKJWIk3aEQk29fpZXULT31UtIYfg0WxMvM
4HYVd0M2xwZx1aOHpvyhIMqbEbspFqlwmh2gYVHacyzHvGsWNLHTUdL8YEFiSZkozs1YxqFbQC5R
BDAKdILZXkKqOTRKwL8dBB44xKbGG94u+52yc6m3T/rKCrvEC+olcCHaGSHqrpFMYrt6vKOL6gue
BiN1KSe8JzCCz0hQQMqHB//Kfm3kCpPa8K8/oPGkkUzvXxonMdbvSALCXgfXc1JAGfrtNkV2OD/h
y6toHIQ5KjkMfnZLQ7JaE4Xc+C/UKkim9ypAzRctUZ/OKrf7UtlA6kgpYWim+fK6djMN8oxZdm0g
thiDACx76OidY9reu8xFPWGSdP5Qj7RzNsPTAFxnzRKIaMf0lwRfJ9g4WNuwN/eV6bB5p7y1qc4r
3CmgAZ9YBFgpsgxL5BatJzfE8brcs+ppooyvRcj7m74yH0X8SSNGQwwPq5BoWfTmW2N0eTGq8ovz
HOGYycQM5nVgz2za02/Nr5wHCWzTrFsbPqpMagiQFRvc+GCRpBraUsl7nnULptGGF/6egg7pGs+5
zlNZ1Cbr+/jIzd4i07LOT0RzWX6j0/66nKQG3GR1esqYkTH5yDxAkKagqTW4Uz1pYCdHZazgxBnM
HcOTiV8YUOwZD44aDSuHihIvsywazh8t5j6cjKWgVjal5rZilTdjslDvEzk7WUk5uIGeb4CcGBUH
n2/PyKNSjwMQ0M6yPTIPGYIEawmCQIpX3pyux6vdLJURROaeJVjCp/wRI9bHmVLrMt7RYwjjYwam
FWbcKFAd4SboFoxWrz4T/827h/vjcRUN7d5u+JDYlxSrwr3jeCJSzOhePdIYOXftjST9p9QJrUuQ
QFqQysKK2eKNB0ehBtMaZfXsdejJGndTvc8L+4npSd4BzncJHVG7VOXlpXTn5NjVKwkkfw6Ml0bj
ykrc6ngE8rc7VT70kXy3ZwuILTgCZzI5phkjoEJ0mgc9ELQvMbbKkQriaStrHILSkw937iQNOLLg
RCW/HO7VeHJbEae5Z2hOStQma/GP8GdeCTtbS4X65GudS7IwZif8TYNq5tjcAu+0nBoihmlfZCFY
BINNeLSuO2XSHrwHy0Gbo4taxWtQk8ATMM1ZyY2rUIovXhOUn3O1jzgWFx3VycAtWJrJofS1CZsz
2N0JAqJ7tYRmeS93YGh3NIHwrK0/AhOL73KRMzjfPKFcScCz31brgOxEWvoqYk8c6YXK8PAY8x15
mPBvc2G7yylCxuNue2uZU7iaYIk1GUDGCXoj0JooFiShQiXb0MqAMUaSsvX8rn9jRKzqRoAK9eMR
BUqkdCN/4MrS8cHs1lrDA2vX9bFIIX7Wz1pUbYwN8Kad7XvEHv11t33cqVLo5sfTEy5hcjArbwvZ
T/XtNUruzyau+o0O0nVHbMYPG5na5asefkaUecUl7/RuxWpG+ziKmQf/J0yc15nyTnWysRm0nut8
mxdjyNDHTv7BqvCaj65j7NBKKKCPRNEOkSxVHPogTXN79tOvOLC+ie1ybfUg50xt9wxWQpoSElLm
fbjQc1SV6JxTHsG1a8pS7p1pt8+F3MElg9GiQLcABqwe4PRzUC3U+Y6ZtvLM6dZD+GXBzkIHz2on
inLxkci1TmOMdrGZpJ6ysofnfQc/yRC4X9LzwUyayhnyl6fZe1DjX6pG4laZa4Zja6iFz264G7bd
c8axNSf9V9JPzGnTkPzAmLZ/uzf3MvqtRATO7zJQdM7oOCz7SGIZXGiPIwOF3j7F+tyg7Qksjyq/
ygSe1yqROEDVJrkur0fbBESLAvQmxUb+uB3EHddIpBUWcXzLnnNGy4qWzaBaXOSyNTjRuOYl+hJ7
voPXLO519aD+NHi8cbr5jMu3hLRbEmC6XEcDgmYXPOd/9B9juQSxkbfUUiW8ov0hvy7PTetf0qMV
8TatAWHmfwPckqz38XlytHBif8pB+E+DZB/PvspO19brDe+IT0pMxrThyM3c2mm1EoIIUX6RXn3e
kmstx6VVFcUddkMyPLo3ZSo6OUmbg2gdAM4eJlkPUwekZlgo3BoUWsBrLFwRSCVy/QhdJDfLYwHF
TORqkyFXfkQVP7fXQI5DPwHP+kHZiUlLG1VTeRoTnEmAyfGMs3w6EDZn9+m3/WPx8Arzigf6bHBY
72Wa2u7Kadx3m43tacE0zAxfdPHM+M2Ugl0S69JlOH0wkGfzCyikTQwg+zEJ8o2h5mGIJ02xbLAX
PVE3VvoNyRZo51AD9MY4MKRh5v2P28D/EbRPuHdDJuJOvt6TX8IE/69qCbKy/vpbuQ7K1zK4Tkcc
zgPRnN6s6ln/lykIUDW/8Rabl4BvZI4IVKg5I3nMx9Md/z+P7PXNPIcuQxAAAvP8/Ska8Erf+s2b
/bFVpFRVDegQX6X/2vNIb3Djs/04GqNlp+Tym5SfZPMmDbSVGU5LKQ63hT+VsECDWWDt3VyXIOXi
yLzIwia2kWGqPTRAWI1ht/xx+ZDhq25NcbX43hlprfzgY0eQkvCUkUnVQSq//sVR+o3qaSYa2zVS
JcX9n10K7D7NAkAxjs02njzGxtxy9mUVKRgiowTI655kbhQMuHdzPi3hnnGTMD5IAcU7eG/2x5a1
inTlQjy5S+69YHnaJgeQ8zl4pbTcDuoBvn8gmgLGsgQgfhuY6l/VRgQLf6NZLltcL96d7kkTEyvl
jeoIAknmngs1JE4q/pEsdpjRqLF3YiEy1b22x10XtkvvBtrkOPRylQTjV8ftdZR9V4UuTlaqfTkL
32yeJtWzzFW7d+kxoIVpUaM3kYJizlOOW8OQR+cx6Nh6eM+U4+osVDVLiuuYi8/GEvewzTNYsIur
W4DO969So7tzEKR6us/gvrvtaK2wIhe1z2NpMn3ivacA4ZWuo1+YK7RfQ01SNSmA4zMfQPsOHFDN
+VmIqAuyWEsxKmxtLOUgseEqG3Rdjgz9/DFsmi0xh5BrbBtyZekGIdDLARHiVs/5orjzeWiJkGzY
VtTCHdQQwQGsJUCajgzpBhfFJZxczqOS3Jb1+5+Z0IPR6kt8q1uYkvzQmOafvG391OG7fdKFHmX1
JbCI+Zri4Eo0Um5zRJ/JE7vTIJlniwddKuD+KB2dyVtosYfOov4bkqrpMTJ80nkx1ZMPeYfZ0CAW
uyRD+jvEyKFcoVnfisx02mHysW71bbbZ4kIf+p2bQV3ChbGcXpFZ9PllJExo4gaa8yjxHEa1KsG/
OnDQ+kFA2H5O+ZjMPj3foyOvteA/N6LvPuHzVZnRkhhcGl2gbRgvTh884mBTSKeprpLd4v4Zih1y
aXrkjNTc+8iQ2PV2UNpdYaE4zIVxq93mUBdBcDbxywnt0c0Ugrox6irfSrHiELVwR6x8CK6KfFes
M8AvpYaVd7jChWUO6MPGHvi0B8XoYHBTojL3UNaFJI4quTJKTY6DJ40gEaPzfwfELPZ9ZHLprB1k
ai4b5Ut5uNJmVbQ2OjC8K0JiNJqhFjg+D9HMNZV8lj6cDuCVOiRPpItHu5jQpf/q40C48F1QKg4n
jz+6+T7HmMlVwkvgUcJa3y2yZnkS42PoxopHkw7YAPtKHlQwfDDQ+TR6iHXfdFcvySB87CkN+Yg2
qyTZ99efZkufxl0zedvFfshhje6xnZS6uc6cJJ7juOZmTEc1ptatCHdw0yAQMAYFKCmGRhh6IuqP
Pg937eG2FPw348gPlYN1zST9jSqUUtX7bqN/J2Y+1+KOPjK/k460PE8AN2S7CCoEk+jRKWwvggCO
IHfmzfO0/giI366CIbwSL80H2KvHhTR2u1agvNJgpaKq5m+Mgw6MdP+emTga+QA4ZGXnzBlm3osX
yLkNy+BQbK4w/5W5/ObqhKhWKBxcIsw/26l3XurmBM3PldPyUpANmjnieZColMvnRwnyFdwS5TJH
5DlZ/PdDoL/dnZlPhz1W3pr7FIPjS3YTWFX5gN8/VqAbepvOB57I0RLbjC2IJT3v8Gh3EXcwF8pR
1UdgM3azzEmuxDK4l8b2Fw7S72+WYw/RNfP4jZ0E3s/lTjDcKoTMEMV/uwDAe+iaAxyhS2iYB/Qa
S8dZE0SJUmjjFMuqLXl0wERND/QlpUfdEgdr9tfGDsLu0DQDHjdYSiUy6WuwXXcIM1CJVjURHw6b
rvV5gbU6Q9fgr1mTskgbc+HP9UiigQOTsv8TZV/1dOby0BtIzV/kw3dDhoZ/FLhwMZrXyCNzLO3E
QnF0NMUcfhXWJnGyqAQ1fJk17gW2NaxzmpdgHmD6pnlprcKluALz+Ecz7SkAy4bMDLPqW9bcKF5W
UkUrPwN8PaDkKV+17MK3VDxHQC0sYjoJveMN8T/5CFOOyje27INPv7j05+xsb/BuwuqD3Dsk7qmT
NzQMIKWXSbbjcR8urCCJ+kiskdlJZXctUXYxqEbdXBuI5FaqRzNVqXueDiZ9Bo11XplCPLRuTFi7
Y6jTeGUH9v1AbkUeLq9iILpwXUnqL6vqQ2udYX9uas28jCpjKMHLYMwbhVdcmk5WWBTwApU49JPY
vPS/eTyTiVZmYPJQczTBvBw+TxwiyPxcRuT6r4WBcDEyei7OYvNFMeiAcgs0NxhqNAU3Xmu25HPj
2jQzMRxBEVNg9tyk3o8exGRxpCgxhpgiP3+JjVYm39Q3OzJd2yiIS9TB66doDj0abDmXlKph10i5
nLkOJgvTy4r0c4X2XKrn0MngcinwQVxZbDRE2MaiVB1zBepWNfLAmtdNIZ2kG1Doyoi+/MgNwo8P
yX+c6qFGchiWTsPHWdvEEw0kNQxWkzcIRcM5mpSVRcfQO2SpkR8lM9y44qJm+pXMa+nRVZt4FPGd
2LtcVe64z6c0M3reHd+IuSarZEP65AoJbSYYYjjHDbM2kFA0H1vyFVEojeNDImkJ2DLa9eQ9TUf0
gVG65Wc9FlJ607PyvWrb0osKGResQLe+SoAEl0gGOpZWzAA73q9ry54eBE9de3VtOvIj+fiqDqaW
TlGROj6uzYHsZXSm3pPK1WpzUrr5FGcHyhIm49F4CefvuDEq0/2u6SCYrMjXy4U+ivotrqL818N8
yKD8U3mQgvJ7NAdLGsh4oLlLld2DV5SOOXPnffWK6QByjcqAgKTZE6AgAz89foIgyzfaNNcqP+W2
vYs9FwHwFImHkA7JYHHsa0XTewtFfkFZsiZoQfMuxrGgBA6EoLJkYzm004GsRGwavUQkWQBeoq/+
+7fOFLfo/1TJTxzOu3z99O3tTUY3bnGVwB9oQgdVQFnnnqFmjiPmQws9mn4twYoakTNsDKqV17Jr
ZjKUu1WypfI0ocwtOl9kD2buTYE0vl6dS3dJEUK0vIElMB+A6kevkRz3S4BQ3xkQE6iM5B32omUW
fdO5rwPQoObqseS+aBejaqCVYzorIufqL4kNsSqram8do5UYtiPw+OB22NxriJuMr7mrACUK4HUR
6A2KaaFnYKiqAa32QqgJNi5Tg+kcd+D+XOYAeS8Ep9AcYVqlRUHIw4G626xCBbcAT4BXc9WUQHzY
/WXjr/+TkAsueSWimod5TnuWvg38UnTQ4G8pdB3ynJiWPVcKMdtWVe9la8ugHqZSIy7sJ1dF9bOc
Cpiwowko0BJjz+O+v25X4v6h4tkZj/S4ZVu2BPlAgzz39HWTZqjVpVXYjwycuX6sjOHPQKK6yRHo
Rq5ZjCqiYlNDd/PyTdIY8yNXHFynRNjZLbpSByHWeXSPAy1mFbkivYZVem5MRCtYsfwEpJU0Vbw4
5E5MIGRI7wH90uKQ9ybjuWeAz6Ddikbu5KKK2Gy4S+FapDfsj7te57LFXW/pn4F7aG52K667Y4UN
iqUlFLue65oSJ+c5jXg/FNwAwdiKnd6JlCD4p39Yt9SRJ9oJajrcPDLul/5bWM8vQgPKJi+d0U35
6GmCi4hpfqLDzzSNbJ0ufaDC2heCKc8ssr6SfP6Nm58vw5WIAdPYR4Zjnls1AOfpQxWSJA7L3daZ
oBK67uhbxjoF0cCi37b9HVWRbnuNm3hmnO7TkhDvHyLsOX+9Tin3UvfL4yRrHpNKS1g368rZo4Pp
kh6PxtyunWws92U420g+QFhrP4CWVOq7Dj9DFft5C1rmnNjAryCLTc2hzSLXiUfhlkodXHkqcSyh
YwL6TzQqiNAfZCWpl1YHHnmjDTgOovhsIiHUA/pAmF4af85tUgDqMIYU1jW/K74zgVEYyk4Gk8h5
h3YVvtFlJoByXx0t61bzKAFuzBKredANIPc0DZQKggMCaAtzOfZmRPfLagBTartuXLByGzGLFO2r
mXqWu7zXZrNVfPDwKIWCOc35EMIi4ANVqkVfE+uocQJ7GqwhGvVJndSgxt9mpyZbW/Ng6kFVTp9H
auA28r3uQx74cGKVczf/9lATvne7p5ZdEb7v0+WtHlBPeCoISBzqh5Rqc7ze+pzRq+bDkPnlo+n2
/Wbs+/tmDuNhgDQIkFytQD5RRQqCXvTjZsxByyX/v6RtsusHxQuBvSr85IL5geXhQpBxI7kISLaV
ck7W71FxKMMzurfroY3Rje6ddHtlXlhIS5SUV20imM7/G1R6PGBmhTk2OcSgcbtERQx0ytBGcpsr
JhWXymYHjSmVKLq+5o228HYqyVitH7sQHXLZLGSWY6lgFhrNXGIvSrc71ANSLRSrtmrbxoBvOyvO
unOwreJntla0TGy+c8lIzwHv41N19PtsR2DlFuifx7X6UMJka4kn4FKFwFxE0Sxq9+kyRgfADA7n
owD8hoPYa2RrzXM5r+2LXNamVsIYnr8v767x/7fHIroF536y/2vBk06FVbhszQztaOV+3IOJ45Kk
BE9M7if7qX2F0UPPiDGTbUqOuzcS7w5HbmbVHIfGUs/kNPDxbCDmEpugRq12cHrXzV1DjYS6DDEf
M3AENvqg+kEZ/vX8O3VDATjE+Y+piYM1qG76J9ufTSWyb2Q4LhU6Sw14dwLVYVL32mrbihgkdprG
6lRZ29OGNKoyozgfkPgILoax1WIc9HUvxG3pfBGCBhb954kbRQWH3v30fUl4LjTXXQeuo48j8BS1
lpZeCu2jU/Hr58OneJFJvQl24ChvHdRvjWpwsO5K3rF809OYB1oZkcI8lNosUU8YK7EIbRfsKMJ0
XMa9r4R9oUCRi8OQTdRQ49mk9zqig2AZyBqie3JCAvouYVmjk92YGzvWIgACVPRtKpKcUrLa4+TD
Gev2YHnj/US3Awm9e1xLrnpP/uBkrxW5q7w5kfiUVy+OQcumYuj1qcjF9tvyb8rg6wQUGB/zzZYU
WL5b5DEP5cESguas/ICECZgZ8gjMyEqLJ4N5VPu2Bzhniq8LZ+KqYzPIz9EfmvlPdkdST9kB5Vdv
C4gUn1ID9AWvOrJQqd6rvUggrhSQOBmFoNhZ2aLJbr/uK0ZQ945xGc4ePDUKuJpTQswo8F4kwLgS
J3o/ENsh3d25fbDn8Z2ObipS83AzVzHdEeaN72NbHSCFsljWvBUsalNtttrxDwzhDgMV55JGgRoA
+EX62PgTPvd5ZH+72tUMe5cTu+fNUmwAiLd9VS/0f9CimBrLJaeZU8XOupwMxuOTYE4TbNpVkS8T
Tk7gtW01o4Vji9N8fGzcdtBPYllXNtnLjtMGXuaCf+Sq2lLXDGSH7dKPz2laYoGe8U55DIYRSOmI
ZRpji/jqH4AuOEygHsazf8dE9+S/0wXk77thl0mTJhKwFS7RYi/R3yDGoPCq5XuHTQE7FvQlsOQc
Of1vTWJ8gH4pCCVpSP/x7Uia4gVHuZmOBWWu9SL+9eAe7vhu5G4u3MhI2eqvgXqim7qerGhCH+2d
+gUjHyyR3XHSn6HpyAH8FUPzAMG+JOgSTwK0mQJzBfeDf60Hl4lAfmqQz3GxtP5NwP6UhCYaL2cU
/mSEWgblXJdzySnFvAxzPthf3ieAe+NnoT3MBowPUNG+JU0pYpDWzBnjfsT6Y6jCu2ije4XAK5gr
slN21KqzRLAPEnBNNDkCsV6faHo2tFuJzxUlhS9SwcSPtKOCaoR6mF8daUKWt1OH/L6vEAQDtDOm
TqMUzs9ERLMLKenMZ5UoDjjQpsBrQxR5R245RkIfgmmoN4SeiiMOZ4K+ltgbaJGOrluTdLCclxmz
KKe5j9dRRnioH3d6hlFBBcDGTskJgxSe9i2yqrZaP2F50yibO08OkZQldRXD9u2BX4j4sH+5JxXC
pnCqGmwOg/HnMIJR0vWaiVZfh0qNM6hGkafPIglwSoLrd796F4whckFTPsnxrJLFM8wGnNfSzDBR
vAemilVgNTeHpxdYQOw/z4t9P3wwF7yfL6bxronK03lzyVnwDDqHFkvainTAGSIJho0IAKAfPhLn
/38C6eJiUHQPPfFCGGbSm8mmShighla//n0eJit7dY6FzTzJqErtSWzDiv4mKT/tPoQfCamSJMwy
lqudDNH96WvS3VVHzT5+UnVlf3PZTOwLCCYxXg+EDGPJDYUqXOeneSOlMxnBVw67vPGEYcXG+ymV
WRwhRjDuvU0Ml4ZAY92TJyu9brCpRDisyqCwkJJtSdXaaGJOFMrzQBpMUZgOlFVCOcVmK1+nvkTB
eSxArrSATLQyzwfmpJJ9uoXiRv3vaVCgezHv4kFMrD0dAkwl+yW6BCF4uAo0vzqUYU4VnMjGqA6L
fdWX/KJk9BHXvZFVPhSoOpExdoqYOBiUddHbfoA2smEuBw3YLChQDeSBY4u75lRow+SxjXNdEtrk
TtEzU8kBib4GzKVdefubAiiboqksiIc7JBXKQMXO14psQF2qwXESFTaenjt4qaQDB73jcg4yHwmF
dnwCK4N+QPBYHmEpEzPLcaK6y9RSo00P831T+RpG7gm/aQA50FVLQKj3K5LIgM6bZZaHE0sk6jlC
Y7Av6CJEU13zhjeF1zYh4xVh57RR6ldasXDoRGuwf5Y/UHTqrd0aHOtf35Q2YgsgsiBESsxh4o0o
ejW86HWGH0l/4VRA0I6zGlHW86PGNSyhyVFbCuysefev8pf0Uagp67u0fp2pZkCP8LqbJ76rkKLu
3b8SkiVycS5crw0gLBZI3hkRwEMUGsE6nQPWmqAKYgAOevNtoDi4XXYBCq+XRf/L+sGNIaDllhkk
AK1nAnxCxtYpFHRmw+YIaUz3YUKHjgwTegjgcu54b168UBf0DnkMXmagV0uPd9j6/iQLNNwKVkMK
6Q7AUuo/yIUn9rJTKLSCXMevp6vDkNRZEu7qE4X7NogIcLHgXjpUWgLWnqdHNTxEAwOvtY+8kMKn
Cx7+U3kjmOoCoN4ZAHlMQgJNtsHu+sS2bJNOo5Svr/n5QZ7HjGWSHVg8UFjbPzbtnc1VYdmIP781
vCSI47aRdnedeEjgQqarF6DeopIa/Qhp9pI7ngtFsfus6daortGqqUspRNk1tdcXUPrRO9sFnTLY
dSTw0uLwWCnHaXK3e8lSgafUyH13Vw0PGXbxTO4Sm7EgMnqi4c3GXrUveMAvsIZ6cXO5gOitNTQE
WSadFmppPuYvxXCTPplbRbwniszMtaTIm4dis8hoIk88BuNAgIpqFjRCGfPOy6WWXjhh0zIooTlF
0oINZL5ZroT1cIu99T2L9q7lElEckPX7cVogEDz9lwWWgihQk/rw0lo/HIkO4rNTLaLVOhn6Nxzu
RUGwjW2Nh9IBZ8RWr6G7Xg4h8ovSFnx8hXCRHPpJOnNFvxS5Ep7SVc2j6Su3Rib7jGoU/bWZDwG8
/Y/cGiw0wbRS+sTacFcOwapqUyY2N+I6sZqqrtRjEb8EjrqNkRHEns9632WMgQJaUoDGevkpMaeX
S3Q7u98Jfhgb/hfNTfDVqdGhdcNO6Tcn3H6F3+R+yxj7TNSYmWCPskDL6JS/U5G7i8sngsAo4PnE
43g4e4ApkjVn9frrHh3qtyYn1cOXqhUtw4CYpsYILkuVXi/sNCrMcAGIOnO9TFEKykp/S1vUDGV7
S7stlN6O9TDYn1ETUzxs8v89+qx05jIbO2icUuu8dIurs307L5/0WCuh/VN0QoUtP1ZmYEwK3Roi
X9f8b1xDWlUr4BhYwHVrHO+MjXzbIO3HuE7K7IqhyfgmqmDgjZ81qs7ClaNylQP4ieR+xx/0ELmo
odMTQoXoX/geWG6uFg8/1PA69GzJ9cS62CtLcIgRxl279kxg9ijgKv0f1XALMiNREfMrKEi0jqcB
Z8AUhCD3htffMCLWgGj5rkqG0bg/zuMfbxft1zep4gNM5GP5tidOLaKdVGSFM+hG6t61Eh76b/Ei
izxgNd2NJvIZGuEH+yW6dBlKHMk3kMhkHqeJmUmajfIjFuJg55W0rGf8FFn6KjuZY73QWuwoF65B
9x8i2/tvN5glTWLgAwqzt1ZllyQ8cTUuK74UqflmRLGmsnC28HSrpnR3Dq3jI5MhX5GeJxWJlQJJ
rxTE3AptDstbAqH25AhQODh9cpx/jO9tLaK3lr72doHmAteCCovTfWWoko/PNxETJ6vSYrk/vTfi
6k9Cheikn5YQBCtqNpO77653TZ9Yb9urlSemFKg0fOKTm+6nkVunrApjr6rKbA+P4JSfWs7bAvd0
NXZ34DXWS1cN+ND6rhaQykh5+byPJdVyH1XBkRzWwI7J+snh9Kejri/U7shPg0eZUBOD81M1zGrp
sTUX7m1qrrY75bDhwN3e4g11FMFtM4xQfs0qqzCRN4Jo1Y44AiYAK+Lm1dzjHqFOwCI3lpDCEakW
HoVtTBEkXBIJ9kcJYELU8b5RezrsOfxUmD7faUj5FmIyhrgpr1MT42JEY1was42qW9biw4lPhSiB
liQ7L4cu5cr++ohAWRVC01zV+feml/nQrKew4OIXf17AIRiXEo/rWbXk4cVMcCYk6Vjd6+tmr7v6
bTDGxIVAaewJYF/+pO49+mmnfznpStZ6KICuiIb1oF3ePtx6vczGY1ZpZ67qspXN8d3WnnHjO2uY
+jLvcivCKQK0TzLvsn8v+c7DLTW9q6oDiHH+dohFeKAubE9m0rrsqEfY0ppS7m5Zz/EMe4DHzO5K
8FOS+O3/+qNHNUxn7p2BMspDYWsFuLOQKfR4P7jM2ueIIEEJisfsfQogczX9l/A0QosVXKWHH5wA
tZ11WfCtavkwk54/pMTVgjePlkXzIa8HYLTKBc7DLXqDm7JDCaaMySpH4YbIWE/bqPwbs9NwJJKo
b+bzPgFonbQDgsNwI495GVTa2q7ICcoXx/TqRCuRxMKJP0hi1xfVLCe8kRpgMK/wBQlUxwqnj/+6
EbIhG0+k0isw53G+EAdjbZpjsOfhxdNJ1ESjAW83s5ebTTIfrzrzWb9qp9wExzIkhAPQBG0QCGYg
B/eD3Qo2e3FELdrJY/4yurrO2SjUK/DpIUcJf5kWo64YQ5m1NCQ6Fj3Jv1e7vXHSmv6xyrGi0S/F
+8RfTgXxnSsGMxSxkbohnSReDU1g5GqqE4Hi57CfS567EN0t8b4XPjoUsiDRVQ/z8iRr5EBGAgBj
zdmEuTe4Wt46ZfkMte/y9vBOfCuVS+/c3Mv+JIh7kkZZHbiFHWNnDSL9rEWrvMmbbTvQ/AHbrGOq
uDhyfY1byD0DfKTpuxftIWokiVTVC2cC0SSm2OXrUPdgF7NBtwVAfopWgdcNLBp7SvjGP8hZf8mr
UHIz+UbdrX0x9/MHLH2BnvREppcb8YBDhb+9AuJypIwaQJ3HeZ33751oaoKHLbTvMaGft3KRdxOb
pXE8Ehj7FffX7EGr5fJYKd3/ZjPiqZS3VU39aMs582mm+kHIWWYPV4gX76CBYFQDl7dTlHKxpolT
FCl6OgTCtAIY872s+/u9q9J1sup9yxVFMkBkNNl7ZhcX2e08s9PS+NvOoceibmMJZgURxFtE7syB
n2TW1/zK8fg1qez7cnEmBFaigaUQJz4dqiGujKJnZR0KolIDCvJ6hqMHrea2DuTqADk6yi8DS6m9
0sC6Mn8jKafQGGES2Nhwu8Y/N7Gyll9EhoI8T2p+nnpy/oOKbx6DNNJbTkEREcbL4SyTohT+1tnE
Duug57I70J+1BxpWWlKRL+/xV8H1mzwtI9EMN86VnL1gc8kjRifDeQntmF/JG5OnzXKaYEQOPjOf
cWjvexvNbLa47rwqQ60dvFjjiIIlznDkBNj9eEODZllo+UVuiWnKXzGTEHe3OWTEt/O32FMVRLbW
oAQmRQiESg3iEAk1PEXt6Liaq8uyZohlrbW1Yh/n/CK+De7LoMf0Kip6RNjNOJy1WbRGE/8Bc8k+
JM+EUBredWQibazvaT5dFbp0QX411/Jf3aR6QMhuNndlaqkYqxRif3nMW9ywhbYeVk/hHI+qGX0g
xWed8B9lB/GUMJxXHcCXmHc7jUDTNgtzBT2FU2PPCIT0Da3XdiTynaq58rUYR4T30TLMHJbzNqNz
UMbevdweAGjm3Fj6w0CZIGxLNG0L/IbdkZA7f3nhQ871JF+xtQY++if9cTaadf/AHgyJ6naEks8F
5dJakgVgMwJ3ztMHj4gsDoxzDJ4W2l+3NqzpddTW6UhroQb+M4a8FnazrRPsyWZF+W63+w3hlIdn
SkpbIUXAaogrf6m+xzAbJ8bjk7G0R4hqWKp+TdfZtbh0vjWJVeS52k/TJfiA0/t1AlStgSC/IlQ1
vM4voFdztOJ7AoT6C1IQwS9SLzMvb/Hi+EUnnxV+2vYAP2EIU2EE5rd/KSFSa4sFVOVh2ee4Jokb
Ie8YrFEITMDp04ft/zuwW73tqaSZaytJQGUH1cP+B83UAuoNZYKwR5ikmbB3phMerEBtSqo34Jc+
xlNuiwmKvXBeUueTgHQ4e4o3hj1hUhLAMBkSWaWpDmkcqeDxHZ7MNdZ0emN4OTI7Z74sWpxX1UVV
VlNZErsESx0LnyDLB2DQ80dQkQ+vVZX+Ck2hyxYc1/W8VxXy7DOdS08oiZbycPrDucapWgGo3VjG
4dJQ+aKEAj/raeiH/4I15tJkQj7Wy6Vo0Z3g76aBZ1fvleDM5eDRkM/KcUZeFXj9YZtRIFxxZIZ/
HiZ4pG7fWyu4WEY5hZ2OuF1Rq9XqHY87iJ4qubfsJJ65jXODCu2VFIpIq1gL9g13arbsEqWmXFeK
YiXU1exM7O33Ncjak6RfC5xr794WTNBbwfsj763HTFxiRdjkqDfv+6sqqQKhYpsmSjhelJYDAV19
IzgQ42M1sC2a98rIJXTnxg/+bTU3alumQSiuUOTLJkS4ZiLgE+JeUNahGZJBeffVynpA+dQZe/P+
IA0ChqAXc+89tMOsL0bL3bqDvG84JwrjiFSDPt2xoWiSVxymOKDExXtFSwiLc+Nx92tAIx2uV/Zw
5IK6bJR65n7gVSRvOBQbTlDywusFBMMBGCXegICoow+FdO6hX30xAjcbaJ7g5pOw+FZOkx70Na+3
0R42zDvphGm4oPCfnqvPmoW7hbk7ZLUpyyP4CCCLBzkB74c1BOfISTKxUj1t0wM0DEpcp/A76/nv
ZwmyL0SGsrUay4cjVsZrDT6NNQvKLjjWbhCVj8TFPSjfyFIV2pjTiBwhgksHBfBE8IO2130Yj6Oj
LXS+RJ/tJ2Ehhv6I2Lo0sbgN5tgonKnT122l4bozC96UdVrK1NbPLmAMCDdP4WtxljKuInyPPVpg
R9dD5cwlRxFL9uaeEDn/pZtq/7tMnWm0LIOuDQt2MEDMhFp4IxuSuB2IK0Xu1PUPjS6rfwVqqqBC
qe8I+F48FcimM7If4EeqX6rl7PJ7H/gJPH4sZYWy3cgrDXcAaFztpVfnlKLs7sTyGvXzaPF05hZa
r//y+U+4YqUb7AkmCjELr99csYOipIGW7so5hft/6VDMlCNigHczI3FEdd6k3G6Pb2DltiFCfQ7v
RG2nuyRbmY4eaRRczovZkb2pkSBcZnhi7G5X78gCWg9fuTIiDiJgS0XPT8VVINLxgRLUrwbRaOs1
FVoaIL+R5xg041YwXH2xJUXxcDBu2u7mYYc3XIZYarOCR1OjiI0wWp90s7FLPc5YQPtRBb4cHwiR
BHQ3G1pCskzgm1oxz3wuC3oCcTRG4dTvJtukLFN7etCqTzUQDH7cmAC4F59xFrM8/sKgZRLYxtQw
jqH7TP14dLKuIKHHqh0Qy6uf/+Q1U6ehoyiQmm0DW52cQz8jTiwP0n5IXdgXgr3WTMsbjsQ3BJfZ
Z5T3VKtXwtetXzN/MymX/Qzb7zcuslw2D9DNkmTL0bfT0CBWh+zFOaT6SM89V+ZMWHM3cmp6w19A
Ac24Suc1COF2HB0LwKZllOtun2EIc4qJZOIj0eVy7i6OjUABOJZ1EEdcku6z3sN9zad8rSpbXkpE
D/f5A2Tvqgc4RRPH5W/4B2j4aDth63wOpa57dz8Vakk946vj1EARuHdiF+EJeNSdTQkn1YM2UJ8z
yoaYRIq9/orSjcAed92P6+0utfR9obQLLRkdDNTEk1MH/tksbClLiJwRIjbog7VUdSkKml5LmwJ1
6yN4Ai/3BvPqSe+s5+KOSVj7sq1ydudFKBO1EKOpMbrCRoBo1d9uu4zE3THfC8EwF/huNteB9s99
M0mN7t0fUunwuipsCCg2DAlyL/6B6fgOU/WF642/B5axTSPrSuYJM7VxVNtKs/MGfkhsv2K9JdvO
AAtomEthMg7Jk0NjrU69pXTuAnTV/omaS8ixaspatxy3vt9hAArD+PQRH+1CrvNHuN8dFH85930v
ZDJY60ZA0qSrftVq9BBIMdA4hQ/0trpTMe9OttursBka81+becs80AbpOM/pY0stCWh9ABb3C1mt
EEXnZnSvDSY6EP5fOaXlJyV8L5sT3kDOgPX82y2Ivee7yoLoVG7z+n3BP/wn8NbcMn+mDDNqjrw4
BwDjOGCKO6R3BrB3ikwAz+YPIcZ/DbvXVmNrFZ1kgmpUhBKptJkxkws27Ldu7rhBPWH50jUPCBNz
wuB3j51tipx/Gffq740zv0FAGTtlW+r/ECMmAWIdsOEvwJdzUNw5dmA99QHoOvC0OQ0Bx21a0gPd
VXxMICcDag9uH1H8M2GZZyLsApGQ+2KPoBxX//2fF4HgJ+E5mwenH0UAM8r3HcFRzMHdbSp6xe0X
0O1r00cVGZQDU5FADGPPCoNAtNrgVprmZZvYga5sPn2F/QWw4NsWI2LLL8T3PWY1XKNejlqNSEkL
hQaywCpuiW1yKXY1vRQgmRYIWpRdwZrhEvFW0nBloGXOjesL9C+Lq5w6AYxL8xVZarWyjXlpMBKO
msfD5AVRzWV/dFomPxLeE2VHRMbYf1D9RjNj4L2FMoq+wkQA/xhITdaukc9qHm5bSNv+HKZu+EO4
Q8tHtHyAD7ia+vUaYVuHnI3+yNQMyeytmrS3LVvOex74f/5aP5zqHjt24DA7Q2uAOncazI2fDvHR
A/OXEf7MW5NNzekFztcBuv/fryvuCtk8rLvulJ+wLsmsokEs/MJ85a+zGa6ncMlGQCx0DXhiLxKO
sVZDFB2AVs0C3HtNCaMDtlGJ7HpdJNRG6zT9u4crr1qGju/A9pv3iqpjvQVuGtYCpPtGAsKdgZtr
P3Eh6PYplwFgtBKR3EbeZ6bnYu6yjTAvje6GEI99T9RydOxIemfG4wG+W/ElJbbPSNlMpmvS/VEr
5d+n0suFIX2sU+876v9ViJAZ18t6TRERRCfiF5w0Ptc3D6M0UPsq574XAfbhSD0Zpueq3sDtUyLs
/zUWTl/5VbMPJtalMDfcSH1oAXQinfQ1ktURp2PVzXnemsNs9HjlCn3U9p/5x17NxI7QgFOzRlNL
OuO5rqO4b8B2YetICTCj36WcksKrhsjiQMPwkga/478Hmpl0U1/uNC/DiCuV6Lk3bdwYUdryQaw2
7mPfH4fiHS+/Mfr26PjQzfnFZ4vUwl3ljyoy8xIPJY0DCs6mtPzi9yYeSDk/8lGMJLt8+CWkKN/O
XAGxC7hmUHE5p4yoTmm47jJIffG7qyEqFg3/8L/JM7PU1kMlmYxTDLtTY9slfAVF6rEUL/MHP5ul
6qV8Z1Be+NoHlAUZ27S+hpg1ruHxieHwGUVCaZvtkHWGyohKHfpRKGmuoyNR0qDHe2WBh7rssIVH
wjB7nMwbaY+QhhohuB0zy+AImpaQshPgy8/ey1tH+r0Ac3AFOIAszDO7lb30YKz+ZbO97IYKZluP
B2mP19XLbyp4h1upQXPs0r7i8wCEOLrJERpWBAE1Tg1xX0pxvSWRqLf+pPX5w8Yl/jumvfJklByS
MjKfg/jadfPyvJ17TP+ZVRbxlyY4bMht/CD/Z0/Y74G7GgB4JvxsrljarmVcQbrA+EvSB4K5p4XD
6cI1zsn4FZ7KhZp2P5rbl8b0RmAHw0xPEaD+zKxMcF6tZ2WTxzxXY9dnQLm6NXQkT3AsKcFnPkb7
SDBZoINGeP0u7OYiwehj9He2atvrrbTBI5xqnPWUvBq2HXrhI+h40FwLLyb9HXq1YlgFKkDfnDO5
AGPqSjQa2HzyPMQBoMqwIeUu86bxWKFd9SOenRtuxKiJZ01mTZ9WEQbLpliURyJwr0W7Ql/sUOvz
e3nofJZ7pd1pwsqS0FNefszsEfnyQG3Wg3TwAbBHnoP0tnVEfLyblQ8VQB0Sg4QIcfMzdzr9/CyM
MtKha8jzZcZ2dc3xEgqUas2d71UMm7rXBGeWdzTw3sJu6BxedvGex+uKnPV5PeTT0T9LL2IA0qbb
DlYxejcoGsX6AXl1J5wzjBBcLyrnP2GKRQKpnYs/He+242JGnwt39mY+0FuHEghy6ow/Y05P8yYx
pyO5zRQ/DSZPn8IzbpPQLnN2O/h2q7V64/4pYiDTnr+nOzuyR1dnZkbvQHZ0MUDZ55xQnwEEZeT0
wIEV5RKy+Cg3MonTJuHLI69VSyqFoHzqUmWwLFWHj891ahdYcnuwXaGR+zlHT7n0TrYvaz+ZIOTc
o84KMFtiDK3VyppXi2N7RZ0UqnHNPlcMHPLMlEMFBrg+tIvpd9rMLooC9C4Dp8JLokjQhdF9Z8I5
jVJaz2ovVsqbvjg/MJ3hlmhEH5aJJduatJDZcLs372WOj3Y1Bp6ClrqOPgmDNT/2Ok/M/jf2j/Ci
EWZTOc8sqS6ZuvYBQajbJmkZbx1avYcti/u5Jgj7ySxCZY2aUIAIzM+CHgNgXu3TM+3LyURIvk2Z
6XD6ncfCLkNQfYkZEYmcTK/jbOpm1j3293KXsuIolYW8fnKl4o4l6ulpqsfzOrUpU6HdnJs0Rzmp
FbaDUQ+vqtdKo5xVCuFGYcw3c7aVLddDNsHLlDI9uvppGk1QQl7VQ3E3RprL0qOM2CA4hzgxf92r
rw2MBQWZ6TmpLN7tVxf0702u9/jJwbzOEtoA+CERYQUncOgrRwHH/1+Q0GSDRTXpnhWlwI7cJswQ
la+eJQNjl6aaHJufkC92Rfk8HIVKnAAnP1zn66OTOx5jK168WfmaDY9d9kr+AGVgHDpz6kzY614R
4o8upTCCx+I9EALE8WZGIQ3wgM0B7I2TPny1nfh4NiokH6UiJ5uBP8ua4mQ7A7+Carf2jdpUVmwu
GSXVAsGkUymWb2eAXP/rTgmrxV86MaHz2S2OT3jHK6tf7zEWrdytsPVjje3pGFZXQkvzrZoRFgnd
V5q+buR0/T1PL3N1mkSyG9ApRIq1gYxUybXYEj29eDvQBayuwnF3F3NQ1r0VLPmijVzeGHyXbg5W
RMKVtRBon2HRhu4Q//9msw51d5NBZ9OdUOZZeSoAmeQ9EBHgp9xk5Xv443PECOpQJl4rIZzhrGX0
zeK0o7eIz6jDzgQmZJOQSWid18TSNj224+0AwqU5sJz4MFL+QdA2NrNIfWqye4b3opwInd/Wx1oU
BQSzcZ9th+3870/g2l2XeYYTgkvWIPcGXzds4YbGZ6pxfsTr8HK5ToMorfWKg9mX2rhB9lobahDa
dOnPUTs3SNiIektrx3XJmcvDrVauUCofezPFFpAkYNOeQJ0oIW9Tt8ctK1we19H1YEfu5v6jLZen
mJJoknMwHIxQLuZceaILpKrK2zLEmKFnzG61jQ0Co4BCKV3BQUxBdOxucaBsjqrC1Vd4WKqFnFpH
U8vPzZ7xe/JiS5Y3LVva8H9UiD2HIjPKhbVyXj6kcVkSiRbe3nIPmjeDxEH1RRF7irgzahhI1ILV
Z2uNsLhat0G6t8bniyogzYbTgdJvhgrHBYhf2FIO4BTd+9vmC3vhfcPYK+qPynmjfMIloCVU5yRr
I52fc9Cfp+BLygLeo5c/eVjQODdbJiRnr3wcamOiSN6fm9UHOjJo68UJERiVxiCzFgon8J1QBsJg
5czEOmR5nXGkig/pDrtNxWL+VyT9JsCpGJ1hhrDJ+rDgopOr/KKfMAKTd+Xzx7uJEHtUfSB0K+av
Nm9CCy9IJj+gmBGUpQB2PiRObA0peKe2k8L+VULexoiH31xzUvZHWXqXsGQryXUIU4jKI9S3rwFS
2ZWLq7S0TuQkyNErEgapXHA74H6drQ+x4EEP1GeuwrrWIGl3yL1gVkrutB9GdMBEj/NnPhONkqBT
py598rceHMddFvNLuLnpbq7DvPlV3G0ysaSX+s46xWFrxkJzaVOCJk4GZbyiF7X8z2n0A7kX/DX4
dlrU4RadqpZAh2HciuSUqMqr4CrpTrpKlEbTTreuJlLHIs6CpOKqmwpLwmND0qaYPyhKwOugOEbQ
XQ8C77NWEfHvqRFwhWlp1/pvsl9U2HS97u2AE4RXHCIQtbAQW3TKqyivLUOZSsRNWX6Yd73rE3Yu
4e58MuOqqLArYgSALAC8g9hh6oSdqxaUZ9j/Ls/ie/GQWGHzFu8CkcT15zE+s10mKCSHSRxunXl8
di+qEuPkDLC3nD3QPpvv3KLUOCrLwKGj05GHi/0lcM55/MOBIod1NSegmy5aisVcYUFD1nvSKrut
2EuwV6nkyr+CwMgyVC1JZomtvMQ2zRH3BU027b9VaPCRNvxyA/yyL3PsgjHyqxNIQAFR7yQvGTN2
sCjI4d0NnIjcaQqAEOoKSQXUrAgUadnKL2lCijux5BzNDc8wAnEn1NxZWxvYo3Bxa1/yzUcnyX+I
EOqNCHSFbsu2Cj2gP1AHnK4WzwLeEP2bVQoSSPgoqF9cLDTgc914J8YX87M6Kqu6+golE0fOvrWP
ghXUoz+TyFILBO9W0oVdb0HFFyqBbgseJcKH9JmP3vHxQTew1+w7vdiAJxXSFxopL/ziKTnsDqza
CKqw7I40S7RfiKqxIfj5tQ5FJfe/FyIqViDtDIFnFNfXblqm1fMXoFc+K6oeBrWPUcFSX9QrVvJV
aFXDnXKVBo2WvvrBOCk9meDefCbCqJcee8RZBuemy8qdtXs6V6OYTr2cCKM0DMhOXAdoldC0DVGR
Lidr5zlUKrEPg1PYixJrmFQV1d3KIyllB4iNumNtOBqhb3w6mZrZina+OMffx6o4ytyp1q1+YIXc
dGRVXD9Uv7djniJs5O5x5t9y8XHWKsL2pIaLNG/GIXtpQimhLXHSx/+Rqq1EKW15VE7DyZzd1jKt
4pGI6a7QtKYY2X3eYmnQTgr00hgv6LCvGWlUlZDMFXNE5HHXh68P1JBGBeVdaqoJV8a6EEyC8F9E
R2rf/dLQoJ+brJMCBu1a5wSjpT3bpQ4rN6J0XvyiWZ9f2ZaJTUw4izPSxOO373dREPIywkBH6S3W
fbEE1wBSwj3qevIZKYKrDzEThKooL7bV4hRCjh288/xg1gWhbgFHAuuhzQ+802dfaUS5/F29wcL4
FFqBzEFQ9J1QTYzAjcFWnYMovjb/2oUvmgYlAb0RqK+cxg/cabxiJYFV/l8cGhQOpfUq5YPTDMCy
nR6pp0n0+cSDpecKpbjZvB/LzwboR2qk4m7O2gCX/B+lxvxbY6KTIk8TuGw3VTOwY/EjOMcHnWVp
YVFJJ0kZ/6yZh7Rn3lYy8Jav/0ALEko6VQNrjllb+Kn/WDoytG3GBGiqL4THP2wxKU8L29w1aXjn
1vCuhSJDsdu7lnpSIndowsyeaiQkZhTHXszdbNOBa5yv6FLV4GopvY7czH7XCZTL8XbEFp3aV+UK
z0tR53WDeuSZJcbouVkOxgMfHB4O0RagsNrMI+8jVXlU3ZHlbhv2wmmixitVGggWX6m5ZDkYWAVQ
8rwPiB4EFxO8VY86DroaqjHVDqJy4KBBtp7PHuywpOyX8y2q58uaMTi/Bv0SlABq2sk2JLzp+V+b
udpWTt+9SIZ/DliIxj5P9fTFGv3WwK/zmxPFfn26f/5/K6MvKdm6KJ9tgKcHz8Uw59eatbkn6RUw
0/1v9Y06WhVHLhZeTNy6/aEd3iKI/3uPdNUnChSGHNhSf8Vp9bPYBqKB7IWlgTqyoX69eZlI519y
uKsV1bDeV4HQqYycr+1lFyxwKnebbNKro9zmeK3pwYhnMzr42bF1MDpfXXmdEYl3t+JSbnt7HN4s
Sk/bfYNuXhPrZWnrWzJP1ZXDvnTX+G02TAOt+SfQ7axRAbnucqwj1XBLBDMi03qOrv2fWMIGOkBM
vcu+K5sYfamwjamt083Jzw6jbb9/XP9F3D280c0zu5L6QO7S78LLv8sY+xD3gyIeghx+yEBF+DNt
VofTH/5s5WQHzg+zb+oWnWRdfiG388zdFFjhXGEfonS+EevR0ogvVMTqCbCkL5yDeLLXgjHmaW8i
n1UfJ2xDJcm21WAjEVuVM/sVM0GjmcWVwXs2ZKMr5Iv3uvHCEzaMlFKMlyAUoB00ZkFGDsdmVnDh
goMHLi0Zt3YIRDEDmM27QhNLRzTihoF+BK78Qnj0EwXpkqryJL1ysLJCNFlTd+P/eW8YzG0hRGos
vd9LvUe1qQMhZinN12SHs7fXo0jDGec8Y4n8zHDNs1OBiXx4g9IUO4AqAIWhpq/COKBd66uly4p8
tV5MQ/JS64nbNzWOW+DAs3/JmMbFct2dcAWOvQQhDHJYB00vdOW+pcnLJe7Sn5fvh/IbJvKL/+Bz
6dZRwNfLRtMo+zSiAgcelw5CwZu/HqQ0Gq/lYlN2SMSgBY60m37lukQD2vR52YAN4Uo/i/8JgQd0
/SEuhkqISO9lJr5fydQS3xG2JwFdEy+x0k6cNLPztoKwojGu1ZClmqEOgVaTyZKjI61onhJ6pIC4
uixWeXTWsKvKA/y04Q+w42tQpArr2ptzMGLWp8sgslne5GwUKwciXLnSR8uwvouG7wMcMj1Lo7qQ
zcKqTRSyswKNjhtusK/iUP1NZ2+XOfOLz/k9ScVKRfgqqu9aeKAwMQarqjU3iZNB4RBm75N7eAab
nPy4DgyujmILEagEs+c6Hve4Z2CUr4Qv+Pzr9cRAi6hw1duEIBm8k5Fe7j+43360vLln50kWTfxW
ylvsWGYsfq24Mr0hjlaJVucGLzdZfibOciE+ISH3oqT2Njx60F8ruXK1EF1DpidqKt7wr5SGQqYK
y7BvCGs030tsQ0+MZc3B6ZELybk74WJdiDpA4aBhX2oWUqpxURZiQjfsplu+r/fosX0kjbOjBKhh
Vqg62p30pw1hghnTmwqZSqgfZShcNSPwPlLJ9iC5bZcqrQif1wcXHH1/d1cWzvE8lF/6ZcZLOpo1
RXrhnb55+CA+IgrGyM0TG/wVt+QCmuXLsiRRRdTl+U+5QuQF4qwEA3OCdvzD62pH2doJck67PN3T
yvbxNTji6YGRvHOb5BjCQtzsHvih76Vgr8bt322fK7ywPxd2LnjDLDjZgou5lO8Yqa8tMi3j1U7c
lIRLnRpgNcJolLhMuoDdyLvhmqcTvAZX+Tya/qoQOXwIV+7+i5nBhmBzARW/b3pka4qEp/G1KDMW
0qNnMCE1kgEfWghKWd0I7BuYb3oXNQpjnVjNK/MjCP2cKXhXa93vq5Fe6Dm9BaYy2Hsneo8j4lpl
AQ11cXnQmiiqoyMuhIpj8ECEHl2Vco29/qQEyEmqgsJPmVpee19a/YaJ8pSULBflOLAcOZBFuOo1
avxm8lrC5276SinYEU6BK4DrCgsfa0g9OYaYzn3zcgJ9JLA7yk2t3OILU/AloKeY2V17ecHJ5zMB
TmNKapuq/EfZ5AaE6GsYaTtUH0hppu5/swH9lA9kKgN2lVdhveaJ/NH/2m3nbcXDRbEReCH7N+OV
jVLd4mxbd5RN/x0AGzzDOU4vyGsIBPL/tVubYDdpURS7HTX2jQUGExrXfswFJ5Wxwxx5o9ZsaM+H
DcMZffKMuJGH1xe5jWSplRmyqNVd294CLqcIblfEwRH1eXcWS9dFHSmj2jC7eiW1quBqQYVV5aA1
9yLkjJy4BPpQh+7tedSUe1zn4KVaNOCHec3ydtxWEMZJiPzvlj9dC3Vny8Md2XP4Aaw3HBDIN85b
UbKE4MvBltuzGscXDKvqDjeyb7Pjk7pyPjPn32Qwt4/nTgWWZ5uSv3IAVOIlIYDocNE0TEMdlqPd
oSfjPw7pdt5fbiEq/67OklZm75zY6jxFVYuO60GqmOTfhG0Lf9itwfLrREkgfPBDBIXD5YTcZ6ZD
9nwyt60QZS9nSndNzDiY8MJ+GamZyahtYYA+M0oG4BxxAmtJ2OPjCiISSbyPbJVR3xMcvjRu7EU4
v2iJ8CRhAqGXwvW2neDbROdBeuF9XfNwSgqKnY2+v6/y7FoO/FFS6tchpdNySqNbRaS+mY90Vg6a
Z9LVk9kd2R7QpdRXpmqnFd77xdK2Yc+/NXkXkypUZHeg8gVQ3ByKCnWOUvZGPhCyFMNSKghxQBv0
ewzm+VvcMO6RHgGKGOz+yjV6zedHxTievggG14yB98DuCxbJfAXBqWNirMLIoPxFBQ5dZJ7jw5Am
jDWhRWxX454WYmM4C3RFWVjjS82oneM66YNp9r0REER9/9hOOFXOVnFAoOpoWemchcBhE8vYQMfZ
+OzniSY0Rz5IT1PBLom7ADMecDKElQWdZM3Rp0htJP3SgPF5EZAMgA8fzvxr//g9XMr0ogzvIsBZ
zm1WgxNBmrGbkrC5uqXqgxYKMoO3g5z5SZlaK/2fXMYUw2tKpi2cfgMNh8Py26EB1EdpAdG9vVTp
r2Sma1IxvQUASUonlesqxCcjK6zkVkUOB9hqoVldR7wcaPiuSlywbkljNXeAPQsGI7N3Vpxa4X4t
OTK392z0nu9k32oiSZHpgnL8BbJz1DXhB+yIxavIOeeiXp7QLjt51d1/nxINjw5P7FLOpTOXyQBn
gKZ/ONtoF7AgsRN31bJ9FcF47OgUJsQoPzyDlP4FKboEbVEQiUBWsuQ0LiCfQWwuwGoenw8lGjZq
b0SM40JnZJR71cMQIAhXgK7XrcbHF5pGrp9V724sJ0/T7mgJ1kAjm/hLG9cFsKU0lSA8j/UEqe14
97tE/qwV+/ZeuoRVFzawwKDAQNkPQeqFR6i//86dBb8Vx7mnVqT8u5kkPZWqgOBchKU7Gk8pUYTi
32JB3CEWfI5an76wH4Iq5NjhD5P0A08+bmnS72VejqR8iY7DnPEmnbB8GFhIbIxsJr8Mmf1K7DA4
eEKn8U2oFM77bHCnfqdM+vgs5U5wzUltJzAUCESOK6AutS/SmPamdws0fSRJa9Q/r7oXMhE7vBVl
O9gG+Igf3pauua4xyWnDwjlvtjoLS0HLidlw5tRi5RF8YBnYzWPK4Lioe9UxiwglCOu/tE/uP4Xy
asyXKZjNrccBFENqdwhEiDfEVnGt7OB8Fl4dqzZ1tXYS+rylshQnW8BKh4Y/l0687Rv0d+5WCsw9
dFqYf7K31fkzZUhETNtQ09x+MyTxzjinyYJkY/Hf5J6ekD2vs9tO+Phv7TsetLSQg1/p1SKEK4td
Q/ltuHH+3ZK74KOcqepGQHxut/vLW4vbxmJbTXd2x9Qa776ZEiyPYuStBBG0WDbFLJanXgIYSipg
2jAJbtGSYyPbHf8nClCGgBVz/E4GnE2Q1l3ChibCQwVoR9xMFfWIdAA34llN8QiPDQpnbecpSsVx
XPmvD/+qwJRA8F4pgRGtRqC6aH0rpJCGc5kVHFBoCSp6PCM+mS7ueEiqOv8Z7oECbYHMzirhkSCK
SJZqt5k5wLTm/4Wcd4z0uUt4zZnyyz4duaLTmQ2PBE4hUYLQNBlHuCbVHiO219MS46lGxUuA10CK
JCGO1dOAUgPibOopppe+fhRNrzkNp9go5NHfohNM1yBS6qIbl3hHxYALuYCbldyWpImJDRkcAlcZ
a3csSkUvVHT01oSLknJC0jR2ERqLs0tkPD3hl+7NGmKmvKh0uH2FdhvPw+XbhOalA+gW58yJiLzo
vmyu1OC+a/vJ8h0QOFrjJ8XY6AlG+/pwivWr6hI+E5Ijzu5eZf5tlbw25AG0e6aKATlTGl91mYiy
mdBVv+ARPEKbZRCcf17lSa+DNLoo+SAYmtRoEf5LB3hrgl4VdPNU9d2Ohqb2xABOWpv/1w+ZXGPc
RuhLINW5GE34KoWC1V7JABPtmzhWY6L+PAw9kC6awHT7JUmHCk++vJR4Cd9L+e7uaMsMUPnKpeEv
yexaIf5cV1ucX0r0OzAfrnL6Vyo20vDv6dWLVSMwwKEHMXh3vfcskMbmyST+JG+a/ab/qQ/pl+JQ
eqgGfch8MKVf3h9I9vynNYiLaM+BAdhMKy2m3r4VXoRtS3f9lT0W58wJ+0JZ6fWOaNuV54CZ1+H2
tRwaRDgSzFl0uyUUCwurVBugIj2Q+GQDhIPWX2nN49SWJr0yT09iiuxOKyuIvp/+SqoA1s24Ii3b
UEGBFo/zyKiZaAItzwP/oGQinBBvzhJHGywI3xVeu5AF9uSNUMrnTVraVojZg5/rs+BFNPlQrloj
MbpKrEig5viuMKzHvaBEU8Gadr/icIKMpKy7ARkFqkhMASNa84jq1jVN6rSZt0GWy8QwHn4STD/b
6xHNB7G2KZfyeJvsrdyFiXA8KrAdFJd8j/7xP4xSmbvtSat5bQPILw8t1MiKyk3Ywbwzl1sTCiee
10xYs8LLB+Lm+YMp5jMyJfdJTsT8T1uVxwzZ0AzEipBBPYKBAgrY85HARjwdorIG3luaYQuiIM/G
1iIK+CFg3kHyEjjFaPBIG+EQfcXKw5InIhlnB3xJyGeJpD4Gy3NYNws6/gHRa38PFE90pJthnxtM
Y6QjyLBlK5+NzJPTBJAabpV4ZuGwwofmLHumpnbe8McRbvr1ocjjAYyl4MPY8PMf74MwvkX7rf6c
FGo+q5dGQB7cVdZw91vutSd8FBqbTCf1owQU8QejineUeNnin3HJ7ca3L/C2+WRjb/Gjnw1hBRik
KIWoV+aI2wUzOSQdD7L2tOJ+5FgETq9WPc7CsOl6tVNBtM/kf9p4UPRpJ8i5HAcJ8+7cqBPoPhmj
hWqY2//m+YiECaRl5EFF3wZ7ki4BnqvEq4Ff54ndmE2AU9s2x5l1Lf2ANIo/e9myfoMXtHcf4OMq
r4jOZqzbCdQXVuGSAS5KYDft6Xt5+PcyojVN9pbT3wAuxmQv8HzTHcOjxRnzYtgL734guPwx/ux1
74Qj8v9rPh5rwlUDX8+AObfF3u68B+8HE+Mxu5cL3zjjb159JM/xll2nn/CRprp3tooFy/Hm60lh
99mNUGCCrmi8ve2oeBJoiRsBPTmAAjvHF5Y0nhaD408hQ4tfvlvk+Bf6CrU040gawLzcU206V8T+
hCw1G/u1+OnMTxw3LsmVBakTKYM5AgCr0UxMvQJ29MKndW02lRYkvzJ5s6Zk87P+Oiwt1IOk9NLk
7BS2U8xoQJMJsDw6qtb2r+ZCz1Bs6bBFSOK1XDXW6KfXGWDUsNb1N4BnnEK6a8Yb+BbiLHv4u16P
9f/fQL1AVjq9jEQQsAkDZO5X354kis7NSPksUsPy41bErdvUk+iuUauoSDsW6Mli8B+w1RLvn+Uk
in0BAJlCPSaxhUFD2UxBDca4amnMjL5vRtmGZmV9bQEMpttWlC/7LT9iukZlpyD4bqllNIIv69HR
3sMsvCw4fBVn7pdY4sZDTCrz8XS36IeoRSIBfA3497C+4mIoL25p/MG4CdXKH2GW6l48folPxVe5
tOaII6aCfz12am7/rqJSjZ3Zh7BxP0tM3UzRBXbJr35ZzqKR3aA7rSci7JsvY5Ejam+ASJStkLD/
kv4sZ2V1zwOJNofCct3VpeynVSL6YnLboNRmjHABpreHqZ0uY807PWmtVR+hlSh71LssTG9ateUn
NBDNU/bAGkCJwlU/mz8RVmqVFAkG1L0rS8tvImLcJu+oa5J/MVSYYWJ7tUufo2BKhQiOERsOo0Oe
BIHwtPYduIRpfK8ER+epxL2dnrDj+UegbH97W9fuNKfU4FPoUbU42i0K5abjgriW3pHolhhZ+zjO
2FyLDAPy76OrMAyRcsulUjcThvtS2XjVFFhLGjBrsR4JXLSzuFlQwfGT0g+ciwYwdAM4+pEu8FeV
7w+f39u5axlQmLdAgLqcxao4hz0ta180um2ZWhBP9RfA7ZDrrTN3RTYiW3rbEaq++k4mviVW/QcZ
eAyrNxUxJrw80toMmn27kk1Y/kSw6G/bI+mZXhRMO9wGrCYRdA0qfHun9xt7Rma9ebCcACTDG/V9
R9LX0jwohnuh3nGzG0EOnp+IWbZp901oMcTflQTzdF0To/AkfX9+H80af9H6OghBWb1n+Wk/PAtT
QaHjbmXqqCr5ppRFgbURyu4GltZC2fADOxg86a3tljySW8NgWOO/Q/33YN7vx8yYi0R6xWt4eU1F
Mv4L7RvUI/VtiJrWgrzErpQcxL+WX+EdXJtaPJl8DuHSV6qvMfHEH+CBk9XK+VDhDN5naqN6vUrq
CGVU65Tnkd32E6MsW+cBW98DaFMH7L3VxHhcIXypTNgmAZPqrOrxFfijcl71x7MFd814RdeS/9lF
FH7BRAXQHWzXpor9Bw8NL5yjk5oZSYD81BaY0M0FKW7JpeeoShVlAHv9APM5I9ewyuCZVFW33RCx
+0qcDdh3a497KprWNExEtQPH5UqWlmntdVnGYnWMMkKOmKCHYrZoTglpqvgde9fX1N9aSRZ2VMxf
0o8ePiZEy9PnImRO38uOow0nqQXG+hT6TuERRFWHki8lPIyf4cGyzfFdJB4eh2ZOtxZiEfCOMIb7
hzLn1DEhwczVKGtEITb1VGUCyC5NKdhUNHaYPzLi9VzWrVGhPrhEoEhpq4fN11BeiyxN/Oqmt2dd
k9hbbS+5tY3jzsklyS6+WosyD4p6F/shbc+Gh9L/PJnCOf1BbeIV5Q5n1d0SIRbEijPCd3nrqiWM
CUV8LqGiRqpW1TKk+BzrmRer+s0qAOit6M/sbIfqaPUU2mrk5tMyR7muMmOFzbrIIM196KNZpBzn
lm8NkfJoXR902Pcsz//kSw0vaU25GwIRIPG92JT1SA+ggaIMjyPSO5Pon3spZcyRWU0HLpxdjBF+
qE3AVZgVkrVBubg8fb02g0lWlk+fePs6xpI5xSv6kEk4XK5siRQB9Ee/24ZLmYLrbDLqgcoNJXSA
nfGPEqx2Nxmbod9/4dYwXu5yZO/4JMgXOKyIJWCf2NdOPXKG9qdsqF9a6PsU27bcMCeA3sOVdrXT
u1h0oskJIbS8QUri6TDoD19mmwN2pBYmHqLAy6YHfE0e5yKQEYjVU6PThIMX1K3UmWbT6FLucDhE
0u6abHlNMSNolXxDaLvsnlUcSO9qspfcXWpkXFWZctO66w7ZuWDFrQoENp9/VshK+XHf3Slm5EvN
cEC6VxOnpaPK4bk/7+fUPIg5chJH9RMF6cckSsG27Zzp8n7hx7G72s3tDiv67fJXwJEdrHWV1y+t
EWnb3Av2NROSmDtCWni8LIVUSuLdB5P2cXIy8Q0lF0t8drP/gaahQtgQ+hZY1nlD0kF3GOJXWJ7i
apfDezriQL0W69J2pm+1vLAFSBnY+O79UNEqoIz243VwSMzXFuPU1zMXpd++l5sSKMUKa/tS9k4M
OrH8WzSxZngyRNPe6ULrQXEn8CnN891ZtxuCUULkvsmHD1PUS0JrJitxN0+MpvwziOoWAEiqM/Pf
6Y64+edtYcG26qMCxbdM5iS8ohyQdLPhDJKv3MF4kzAx9vBtopG7aroyFxi59xnebgR+/JJFQ9r/
6xblNtv1F7xQW1IbvCmr8EBQN2710NzgHFVRExnynP3V44zFdk5B/L04JFlj1608KStrj9fy6HVV
nFouAq4j9yvZnwiPF+f7eB0RpFkjqwknt7oGqfUFioTqLG9Y7GUc7wUphiqfdjodfRcAOssc0sdA
9NWx5NHTfCxnMM6bYIk5DJjhHKAHjLiUmJjtVIzkLFMSzBDU7W/P0tnvGi5wFCk38vjNx0B6HwvW
YIfxBDZHIc/j0oOT1tOAx83acOuG59AHpk6rCmJsbX1+i4SUhUNh1ntHsNFd8kx/VFirMkH7JJGw
KpmyoLXKYlf2ajTolFAZ/1TTaWwjku0TeF6ufSUdwBp6wHy045rtf5J4vc11qPrbXAfaP4X90JNo
b8QPRVb6fuImr+ZyayVwnobuXXavIKNh/CubB12EwUbQGsou0bD4v+DLZ15hVSMOsyS1pJCFpA/m
TAV/DHLweM2D/sHEYXYujP1M3kCRLghRJ7r4nmtCrTNyKD5xd43SwbRdMOM0AmmaxZwNRuAUg+d7
IvB/fVkCJYXPotTKV9PzMCetUGfPd75usf8Wca/OUqxSyjxpn8JoCeLISt06Vk8+WwC1NkDw4AHG
1yGexXAs3DiW2FgCLbtoWEblMDWxtd6W4LM+84OvU3g1NN0UQp4PzGbORGYtuiTyEi/UmEo1LaLv
KQViV1w53ZGBPobnU1bov3aN9Vk6AfCAKLXoiG9+ZjKSheNM8BsrascxWbquHdlxthrpIY4R3UwK
59RugSH29Ppl0NsNFSKhfeNO/uv+29JwCsRK1LKLGtIopvGv7c+YJqUBm3RDAO/Mv6x+y/D46JJH
3cQopx0Wws4fa8L7mJbfFIGoKuGToy8dA4j8SF/hNkbCwr2Ms5VFJqhxU5wkPWUeApmnYBqXzZ8T
tj5XLtxSCpFA75UZ9tj64rcGEQ2iYdbWVbY19dFVUGwQMvIpRMbBELRAInW892Vi6LRRg/ZQQW9/
BjJYjnxqkARxyZhsnBo67TFwaBChTM1cULcix/6eLkILyGAqhwiukiYxagFT7GKkETjgg6qf9IB8
X4zkBUvdXpx0HNqnZvjoEiQSDtWs3K5bRBgTgOEJ9GD/pMa0kWqruO0J+piXY8i9e99vv8QEKKlO
mKqm2tUjro1Ri/oagFBku40rcWFyR8Rxn0fBEU4pBa56A3wfixHjoH6RF1JCHYzXr/kmv57+KIQD
Ud0EzLBnMu94kWNULyRKwDx3KZoePdWdabY8lKXDCU2QKQ65lAgn4KAnHeIPK/JV7F8geM7QRAO0
GiE1lBr+pPn9CtN4894hUK+lmBVD3g9+P+MX5PvjfAFZzzWCrlVCb/pwVCccrCFunYBNL4zHvuvO
9b/A3p+driiFaP/5sGeTLYlD4kmIRay/CTWtyv0UovcSuLyqA5EhvMBsM8EOzXNlovpx/ZNGMkYa
KRIkP5EP3UWeSkNifzQY/6G5xXaMzkfbPOwYi2RPjuyFq8wwNw6W3F1PLlKFdIS3ENwN/TCC0aPx
cOvB+/aD6BHa619VdHc24fLobt2+Q9hTP66oFaihdu9nP6Dlbmp5WhsBdzFLJRrPJIOmvl3f+RG0
TvaXDpwFqwxoX6KO8lsrCpuvWzshbOLC2H+n6rFKBb29pA2NPbzWqvlFOkJcPcEDG5JmPZFuqWOQ
Gn+4t4SwTwRWCfwKQ6zvl3HN63T6QZVyUsuxdt6CmbGN8JJra7L/ti8RM2Y00RfgP2CUPcDefiRu
IFuK/g8j1KYWA38gnLEoWrPOVqimppIiZHMkBIKtjHmN6s/mKTUBoirANlY98yBvlVRBppIXa7aW
jGfCNLDVDTE5R+aVFpeqKA1XgaHweUy41a0WnCo4Og3xUZlOzwSyNP3fIu9mliexPsGRJwGsYaCd
ia4S2/F0/SWUN4s7NZR7WqE31K25cG5UDiTVHCZlCvgjSVL1LihOn/m2fSHvREjE3KgXAfq6oNLQ
oFKhBwyxGVLCezB89tx/Xw7cHLEbJprvR44jwXIrTijlkVupE0l9Gji4BzXWjTtVZS6YOmKWhrMl
/LV8kQrJ+HntEznm6rI8/oKwJwzvE01je0eX76FiTtElnjKheLd1/T35TIKhSNQSP2+VHgknYXev
D8g4FumHa5ztK7V/ye1wnZwlv2yj4RicGEqDdrrdtKJeKoze6K+DIo7lROT5UbURcnpV2+hJ65Ii
bgXA/V9oYV7YAVUcXgWSqO4frIPjPMkwK1XGVajnIN1CbnHDhj1Y7AdDEo5op8INycvR1+ktiN52
zh8OMav34cs4qjXJL9j1XLdPWfk8PX5M3FiVMpeom8/YYCOtJLR8nDXOpmBAkqKDSwt8waZ1RWzr
KUgUg/g+1wAVQzZGFa/dXViGHQZnHc6EmAa6h3EtIXPpRZMX7diDyszbgtOusHZrsygLP2jvAXq/
o92dQgruaRavwuMBssp3NPo78THKhngYAyYBrU40XSiOChrULfGTo67xf6qiQrPP2wXnHKAdCioo
fVps1gmAvepGGHbDiQF1YBPJ13R5w+e5dnt4tDB+szJkVbaD/plRNHY/lJYc6U4M4ZatSkGVkOTg
01Vw9v/7/r28/75UvaEGggZ6DlY9GnGLwWjKSl5CCLVY2TTefk1WHGc7eRfSTUScXqlCvUYkw4a8
l6ObVIHpqLMimpANqJE7KCktVgPf/c6frQofoYVF/MHIhmSzzTbh0I3m3c48ZrqzjAtD7sBWBc6T
O0M7xsaD0MjgllSMPVo9D0mQeJSz5R/wVY4crVQKd32tvH2fx/4Dyxid2rOEUzOazDrlg/54W/27
ln6vhr7XBUYOErps/xxe7Pu46en3uh+1RAY81kpSxn7mWVufugW/NsfKMpF5AY3EYpkmKUHR9eQz
Aiw/wj0/Ub2eWLRuHIRDUklM02O5JwR4UQMEO/6xtZij3XILKg8JmE/zB///J8QiPBSVZjSW/RGT
Jxygt5fp0BAkDc01WLY8IsQVwLWEfNa8hfag6qql/KYd1x5gkJ0aR84BI0Ht9BNryp9I3mT94rzW
pc/XFa92pF4FtBfE+wz7YfMsK9IwA1uBtyO6IqGpB6ORNcnMrmA8yZkT4gG2Bak9i1Wvl6v4u+uc
IQNkdUBGjBNLIGlv+E2G/jRne9m/rhDPF6DmRjo1xc6x0XzOPelcxLpdC7Tfyk5Wc7nn7H1PWydS
WZbMgqEamyJBA88eeRZxZn7vQMfzgHvnBbFCfk0Kq3foV6W9cTUY5+Vq6M656eu2aupmrTkXhFKO
RpK7BRMW5B7NNBIcwd/6g2TiSwEkLWGj3WK/IInRnLG9kFUu2aRm5MZ5jJSHgNwlSI00/K1UPX9F
Q9Z2ee9M1GcLUzStqpZA15LIqmogGZUEVIah6H2MSNlddPa43Hy7QVE6wwEwvjMMv1KB9votcqBO
66fW2aeY5AvKiJ6W8GE+OW2PvZyItTsNlHREBKPEg9f/DAVSxwwLljRKAtPNIYg6CoWc18b/B/He
wi9n3H/XIJQwGTssXq4UORpcXtB6FPw5NFiy1LXllzc+Q3hIvb/2KD8TH+UXYHDQwC+3VClcKxXj
rh/QJm+IelWm63DT+toWm9K1KemlAeOqQT/d2xd6PekXzACszjdvdmfLY0/PWQGB+PLlueyDW/S1
eR15YkMlTIoefpc2XQYEHYpu2F+8ZatOkn8nXqHPUjiJ9ub8oksgtnh32mkH9t80rC1Kfax1VZYs
q5CHYEJb6QbWcbROxUa3JGfcVF41sV5pD0B0K0VmNNfUpM9bkKuhchIXOAEcvDo1MpjtTjK+vA8G
CN8UWxl9H8zmRIxizT6JnL1F8WKodhSx36bBBs/4QvvLFEm2Pb+FQPdJfitWYHbfAkN4d5hHXiEi
2+KgAA4rocIzti5RhM7zAsxYc2tDZ66lgETQ4k/eFUjB6jLnzZ5E+FCJE+7h1OSKI8ChJZpqmX6o
wW+oRxpOzIz46fDvSZF/uQpaSTNkdGNEUWijUXcnSJiJA3YdNpBMsGfJKpR30/ttTuzrUT5Moobu
gilX0Isu4jEeGUxoP26Dd3xUdbmuq3ZY3rzc+bJTBhp/sZeodwxHwa5B/xBnkqTtPrIrPSLlQv18
yiWI84rpUXMr0WG9h25YPvzVh25rcbIab5F4K2J0Jzz2PfLRrTExGaJN7hlqKkbT6Ika2I6oKFyq
J9nXWZgDcXj5HoztQTl26leue8aU9exBYDU7BBCGoYZNzktn6s/DASK3ppEhOHWoBbGpzlVB3HeF
XEZGlLsq1BWSKAicTZ901JRsbo5thseylT2V6ZgMkAhM8RkuZpPcWXwg3/wogO4psbYfI4UJQd4E
Q+dfhpPs7n8K6ZLCJunJFhfUc9ebCaxUghDJz3OjWBFgxwCjahCO2rGhX2Qog7igiDJUB8KM/Jlm
XuT1CDMSTWu0mjpgL+aX2JyTl4ZVMFouAo5IFzVyG/HE5ivj319sgtT2+SlVmgJnQ/Q1X/xAem23
5o5owYpB3iWQm7c7UAlZCcQ7tdy/OnNnlO4BrdOVTpD2lLLg4msH2P5KBH2vE3hF87p+w8uvyfms
f9Kvcrr1evO5eXqQjwA+NKsN5hyVDdcqTqpeUSBZlicauVplvixGeQEHK7POMZWZS5D7c18SIkWC
ifwaDnrzs3B3HRzJwO2knlTdXhZbEbOdrqH3ef2qJ7sToRJbIbJGCyTWK3BNTO03/XGqfDc6FRAm
dsx0ojjmAqJot2WRqaH6bs2FuZrmz07/kB59Mb1lqC+T96ZymWO/vRgU0JAM8v1UOZpp/nHCV6jU
AHJ9Pw+AcGlmBBXsqEFnOKZZojRPh7Dig1CBD/gPtbl9D59pNmaUhMjmVEjsYXlPBdDIfJ7BvjmZ
/gfEi6ui7jpPRdPUXSccaUVecbt+HffTRJm1o8BcGcWDjSbZ5h+cXWBxC2basj7AYx3i/Eg10eDZ
5M6fKhF1h8HpwupfvxGkskUcw9Y36BBatZ0cPqOyS8tmMH+1AowiSvY3Zp10qQyJpgS46bndf/t/
53zr04w82zhwO/WlcZzlx5THT4o6T0aJad10ERlRh8GFNla9/wFGQxbevCp/eX74bE8h0pfWYuJQ
AfuZamP8tJRJQ0uJfn5jV5A2+TF0SEa9ye4x/xl5dPgH1cXjYvCLmKfpm1Ng3DT/pwI/AJbv3tMw
z7VeA7Zz6o8EUZyGqybJq5oeL7JLsMZC+8zcaputRjqoIoF+hyYUzvev/dnTiAd3RzRrORCalvcK
4FgtPBbkTWJsS1R7RIMACQf2QqD1vsYCrJ/iwpf7vwa7z4adLNJzMPVI8RsAx9cn1WY/0FJavOE0
pcpKtLWqGBqt7myXGxqbjHtcxW3AN7PLLbMjLypEZ/o02JqGwclppvzsIEtaRl23lvc/lKwo317/
iFx9xhzK0DurT3JlZ3Z9bdPxNgnbC0pCmpHdO/TChmstbH0JHz5Zxpxqi77KLRnpcEKMPHvr7JBp
lFZZMLcfCutsIJUd/OGyxWnUWL6qpwVbCAC1M4NSeeXYn4lCGNuEH1HMvwljRwP+w/8DCqicdhFI
MFrm+Mu9GEM1IX00u/+WHkzRmfUPWN2rbRiTZuDAo3qo27C1+dzOxJ5orfmmAPC8khL/cKXmaCOb
lXOQvHaCMJ0c8Ifi3UmJJuGb+MxB3xaiKnC/RsDP6MdVw807DCzOl4oGGfWar6q+53bTO8LaDBxE
yeOkeqTc+nNY2hzfmLKmzFpmKRw79lsxv6unj3puVJkcf3jBQ91jQUpgG37gbZO5t9oR0YiN+g9E
junQJLehadt1fa/qArfMa6pIhxq/ZoRndP+8u91D6afQFrya6al+G79KsCZPEfryzKMjSA1Ce0hS
TUpzUmwp+4Y0EVZOq7u+Rc8Phl4CjHQnR4q639fBiwj54uezJNGPQJ3yqGQ0g4W7O24qY4gJPphK
6MJ69qKdnRgVC+QR6usxejradN7CE09A3rbVXMDRIkGQJpTR4dfGiTTtOQ5HBDcIhijog/6BYoLv
ZaSnooaD/RWQo1Xo1S9hkDnqOFimuZ9dwU7Tl/IB3KXJrQ0oO+CUW3QltxmFiOMw+8FqjFlf5XS8
Wmo5dDQaEKViuNRhXAKeOM4ktktO0QU2cEIHxsLSFzTXGFQS1IU4DHrUQFU+kd8hPSq47DjkWVBt
KOZqpCul1+UokDIl0rmek88JwrGzutA/SrAyQ2/4LRuhdt74+SyOUu6N9BwLInYGjgN1jlfqE966
ioSICMpSc8M81Bl38RhI1sdDmyafEnbvZLZZmlb4rtYg3wJM3IgTLaH3xc782yq27CtOf7wv38Oy
F0oALHPuouRnjTDJD/7eY6SpAiaawokAFsWl4DvB/oQWtpyTv5q3YRF9bCcvFj0db1f0sRTYocrw
bo7qVZyHYrzT+Gi/2/FPkqub9coOsF4eTbr70wJ/GAtaFWrqB/kDcPajZJHmXGJk7nDM0Jny8wEQ
vr0moss7cHN66tFca9tT/d2oUmmqPeDV2iF6/2TS9KAebJOwSdGGHBiAkwcHRkjFlo+oEIutNWl1
ZMankg3B4s18s9S0SPLS9/g+QC3lbr38F6HyOcg9UViASsbdJ1WX5h8ze6KDL/+n34aaDuUFCmH/
O6m7Oa6ot6AQWI5l/Fg7CwBMuMwm8NRKlQ3F4Dk9tYbC/7YiLw/Y/JC9lsk96JXoSh3IaAS/x3gk
34vFCn9s6ZJY86x0Siydr+vJzMR0NLOkXv7uay1e3HfcnTGzBX31CLDpqmqcgLJI2rJHNCv22BSb
gdokeapANnDvxZ3ngEbU8BxIymRwduAQXm/DAaSTdG4Gf1uMBuvMHxxtTl8xXBIs7Dh20qFDhOfZ
Rzhig1h4XjxF5nTTCNWSnSraPli+kLLhJkcVg0gu83Gk4EUESKXSjA5/xfxpLmtmGO7mZopB0DTV
mc3u1r1EDMfcD0F1wJnpMFohTPy44bsesee4oBIzQ6MKrSWgh4ZJBwmlYJO6nufxBjolb/Dhdu1t
10gmaaB4BCmyBfZ/utFPfkVWSmgfKIK7HTjjEhpywfsGfvd9nAm7NgAXqyPwfNZaQOjyDfML7I/8
z9eogsgpv8Opps/9WvRHcEhkhiYLPMC95tlHqQ8wNO2rPQO2D2pEn3NzEkrKUKWyq0o/48iP1N7e
Gt+MCzzvtMm7ZGHvzqdL6IK/AXlw92YBYA5j1GznfQ1i9r4Gre2thWtYmCK3RDzoFJNENLja5c4p
1cDBqkem3bCO/1B3/DosQUx7aeHeKO+wq/2nvetLIy1wHqyiswgNoCG17TK/d4xn9BRuB1ws66cn
zE2VJ8btwqVGO8uSPj4bTW2ygyH+PuLMJUbihLjgg6+TG3c11LiwvgRPwJQhtGxlvxKhFBAK039B
PPvt+gcwda60HE1pXqUG6tvwEe/0Xp6XoRKjoWxUCiSGNFlHUQMiwuC0yuoC5BbYsghsbJBV4Jq3
KFKRQbPzMSCcIRzaGtHieotHQcVHPCBFU8CfMA6j6fPjxlMbgGyVLtGZiadofmxW176qQAoYoFh7
G3M5J3DWW+/F6TA0U9wKMsq3CrPQIqMuN4/w1D2TdvYuvwj2BZ1HeLbsZrf4Bi6K876npESumQJl
AXUlhWV6kB8KwpyPv+/6VsYRIUK+KapeD9oG7lE+BDDFGbz25K9COqPEG3zJoiAU8Ky5F1Fj+dO5
xWRPq7Ep9KSGmy13TY/LarW5yAqAtMSxrksuoxJGBuxcOOL+3tmP1ToLupCFYCaQ000zgp+I1Z9h
gXyF+lovFMBsAJNKQfI7a2btoSzDbDYDjFQDa/NaSsfRIjkp3AI2BjX/CS+X7e3HrCywKIRM4WAY
D/XzHxPIgC6qipw2g2Z+c8FoyQrKwR2DoF6SvFB6xyvVYfh47jBxxsvzzIS21HTy2sRMz3sPbNG5
qKPIUYR+csF/XQ8RJoO2hUP50P70YB9x4ew3cnG7OVgyR0EvrQpe/1KvYuwdT0fDqhw3clW3G+Sr
gEK/Id9mcjOJAgp2COfIwySHVX7elii4SxPDZBhWxK8K+Axkw9xW0Ier2y8JnLJh4ZfgvKHfoOh6
wXJ4wUs9UTgZAYYMj8j1OrRpVlg+MpkGi4KSKSHPVk9FuOoRBjZawwMt6uZleGRYg4MGJ+leIdvu
eUVCwiPUEcqIhPKS7wE4YS8gGaHtnWAus2zafJTHkiSOW6c5WI7pyH+UI4ap5cSUaQa9IrFArcs6
VIFWyZZ3DmierAPdZlDJyGRtlHRjIYyufpOMl9d3rDJ+i2ldzvJqjLdo7CSeT+3vsgmqQVyUndjW
4uZgvOQU7DibegLXR9O4+Q9/bEYnE+Newrg0Gan/2PnvLXJlrOMXAs0v38V2WZMdFBmVSFHvF/Ov
SlXU7eR45rnKTd39TJoSg/LmiSnyK7+Iqxx3iZIe0RMqKqBY+cHcJr1m9h7NvrOp7ekuhPIrRz0T
QeRCvYewzPQkAMGeHHMYPvlMkfBi23bJ5Ls8d9eG1EJYEXc+62y3bwIh9v5WlWUYT34trIP9HrPn
5EtHVMkeynBUYZp9vH0mtNV7194q2zx9TQnEmak6/iZXGWs8W5tzIReuxCRW1tP58q8QV4oO1RCT
MwYNvYlgcEnaPy2t+ebW4+Tb5Cb3iwjEYAnfNUTger9Dnza/mEf1yLZ0MRbW8Leb7YZNNIHNLODM
vdBEy6TG2bb/hkmL9WSMcMxFWBwgGBN/6KfGZ2PvcOEV473me1NPx93LCANXyex3RpnAUYVrYZFV
0lsAmZEsAY9kb6db0Vk9yXVBAudd66ej7YRL4f389oafUTxK1eOh5WWZg1XviiV4h93DnipVhVFI
/KPIQLZht/QvKxvaImqf3+JEIwId68tOcos48kEhHgGQQPaezacw3HqtMMNfm7q6EnZYnbyG68aB
fpC3QIFoPZgGNqnVFEQd6eQ365AA2GckJOtuInVAaKQnbeRiY0JgOBg6MrmRq/WpGiEZs21W2KAr
v6I/5bjpkCsfsY/ebNBwZi/hcES9MVWjBLgemk+qkP9Mz9iaSSyPaG+tKrpwncho+TI2RsNcc7No
JJRwpP3g3B6CFuotLstuCkG3s0K+d71Ebe58HxZD5m1Y0oJhFOw+pwyMrirxz/VT+fg1KWIi1dGM
RJJV8UFzJ4njwlNA+AQf55SEfMybUnkvDKYbg9VQ3PO1OhDa2n4BDj2GgcN4qpC+mzajyML94+KF
jDtjUa/lkXFP5WRIgqALtPctESYI+7oLYZk6ujQqNoNEpL7GGdQa9RgCbZi/1SGGB6t/VWz6+b7Q
XMcvM9BM3N7xrrvASnzazSoUtyB9OSi4HMd5abhz4Qwmli31xYQBVuRjfBPMRZe60B8yYUNuB387
1k1YD+hgFgTYTlA8CI3kWwe35PLuSx7ATQAE5VyDJRLQe2WCs8lDk5/xD4TYRq8n4b/RbPSVyaVo
EymY9nRNkAicGOdlSxfyeSwSzYaZc/a1YdjxTpJ9+AOTI95H+ExOYryvhO7r4shyGs7/qH5ZYIec
fc2zyyJTVCiGxNL5N/r1VS1cFd8hvzrGZLLD627pjiZxwfVE8cmUGMiHD546ugf4WV8hnlfmit+Z
OW3VjTN0qAJWM3QA+EngY2iUc074ZnVOWDbF7KZxbTA25MPucvIXLIzW/7RAttUXwYTc4uKw2A9W
gHzdxyOebvNYjAz+yNPr8Vdo2wvtrdwNvNnid/W9FK2fXH0iwY7l/IW+MIgz3C9qg+lRoHiUpqwg
IrqrJHtSSP2kVwpSdZ4zlZ1mAQwWoPTH2Ku4408XPlzF6mMkp5ncLK3THSk10BmEXFBnWNoizslZ
RJfYN06nNjr1GXCbYM3zuS3uUkGLdssNtlJyYSoX8LQD2pbUmtWmr+OVLivYRttc2Zj/42KbpoNV
GyjAEYhE0CUx8c+7sTvSTQeMvj37rtvcVTwCRN+RQp6qRT1VGoHPv/Qq8p+LulaxM+trg3qmFbzK
eWtk12U5XH9tP1QKCw6pvf9ITAiPV0lfxZupGabPB2koaaSTaKPT8x/59po5j8s269JjweDopeoS
FUQRgX1mSfVcjsqYvQB8sq8IFaigrnbXY7NjW2NI1okx3G+9u3EUkxdKzAlge/t9JPwka+iu2Unr
NlOIMeXDQ5FS0wVB0fEAZaZjecSDbuHtH3m3d1tm3dctNBLogr3lXnrP5HH13FfS3IVHeT0bS1X0
BqIkuU58pslH15SHr3d7eiKx1POOu5F7BH9BnAzAAnn0uVsJJoU6OudFsfTNigNIdIh1f6w/dHpQ
R0ZF2cFIlW/UH9VBGMnS+WDp5puRxEhfXIOtmVtf9JN4r9N+MyWT4wGLlPlb8t9Xyxkp+S9zF+F+
fVV/9i98Lz8VfUd37BRZL/ti//SV+q9yBQ1hyd1mD6XQGmy9BSow8Jp1mrkhadCV+Ci3qiq0ahHF
xxr5UPCdui9O7ulZp+dnYp3slnpvPYAq07W7+rgEC27HzQ2HgpESLMUKs3dHOlk448LVnU/gKwUz
KFlLqjO5CmgCbXgLgIobLgudGnGmJERKyJIqbq0+uTD1daxfOEwMiHzZsYfxtmRd3fDzrGYk9MJq
TpCCHs/0IKk1ninpCV0fzPQMYX0uIONuc4Rr2+xRINIFKRFTfDPkQGv4sQXLWaddAt50jRgSO4Gi
3SgMp9kxDrR/hZC5MhFZdzlLJVG3U6qIpcgv4zWSx5iOQ39V+Wm+Cvrck24vJAlmyzgKJN+qeSDz
SKAmlE3xtdJHyjIV0tJ217J5K7WrsgvJ9ag25utad7JJr4XOxoNwmg6nfu1Iu0l7WdJ/FrjH7AjK
UolatV8WaiDIZwb6+ctT7yXxCHoQKLcnAhba5iwQPhABTd3l9UQlOA6O341IFQXFCejp3LA1Z3r+
re2RV3hrJ9hWLJ+BjTtEMkXE/EglcYvbaFrjqru3N8BU9GNQmFTWJMumtthlxKSEWcsQBD/mYM1o
e8WFmCdvOo8aHNFfezGnNXrPorwMRCpRrRV4cksqWqU2MiLo0c/mzjfmMA8/cRODGELOiUxQZOFG
kqXyiXoLRA+GcZYOzi3tOo8JPMHCjqszRHzHJ8N9L2buwxSYSJzjbIqpYDLVPuUV5SHg4GqG+KS9
G0UaIadlTWWBIH0wXzlQv6VF04ON/eWbQMCcLNQUnoP+23yspvyhNZxIC7F+uDpugq0wK0W1yrco
ag0nJOdCoLvYU86ZuBNHXWxr23BPKq1WbD0oLISK/vdr4RIzzyP3nr+7+suDL57ShEoplf5BKknV
0A7xYgU28iqJNxwYaAWO7k7bOO2tSKmZYpN2sElHNIX5owtlLbXgeWg/JR04PTKKjbe4yJv+8c9t
PwZczqKd7ouAHCIHKQcIn7EFL1unqrNZGy3ucTneX4bLlneDJbZilvjFIP4sOv4nqw1e7kxM8NHL
WdHzhOrU2IMOWXkbdD9xIsTtVyN84oMeBctgg/eCRsMsbSglrz+RKpvyQ9gjBUFhR6h+T9tn5egy
5A+pzGH6DwhQo7v2yN/cdmf6pg24WiQNL3Q1Mx5jkOiQPCi5wec1ZMs7zruElbs+Czv//iq8KxGH
pLayVVD/q8o9ZknA/sh1Zx011+p8/52efuFP2NpSThoASOZ0kzWqFIATZkFaiX2uBz0Jl+vkMrN8
4nOeoHNx+YNusCCWfoCwkhM+hxsxhvFodHhu/xpyopYfimx+tL37yleZBu15tD23ocJmR6vs89DS
PnwysHRIBvZbqL6Te9LPjOx6C9D7IZYCCDwx1N9MtotLFdDlKxNcUWgHCY1owXc+/5kBfNWFfQvT
wAaJcu1sTl6/rcjeJ22fpq5jbQCRb+Yvt5+cnZQ8hzg+YS/XRwQOVFnoVLLMGDQ6OKraufT15P8t
Ew5LOQclRPTlEFPAAbsMc+nRAK2w3jMHWc+XZxDUInn3oXAW+6w08RpLOXvocRhHbGOCWfoIhz0S
wl3F8kunJJ1JcwEFz/0BYnn48ky++OKh68FvXx8IbgNldHPXMOCipdUwaEovH+35t/PSyIsISCh6
52shxlz6pDqahekUXkGoRJ26REa42Bl8vHcaYrzRbh3BpySWv1aJ/sNp6RCYbK2bIklCQq85hZHJ
YTh9e4kxcSrz5tEejtMvBuUlIkldxT7bcLZ6h2I5V2b2DxeTciltzVDR7DfAFbuqlSMikF/kkNzy
2lrM/+vSBmnLmcdtGHm6HX/zl1MeiohUFKh41gId96rjRBAusUyqWMXuVSgloJhDQOitJLcYvAsj
M1D3cHvzyC0CTIl1/eYQUeeTtLhex0+L2PVnu73FGqe1Dju/TQRhmi5GAEmEhhrZ5pygjAn6xq5y
WV+d2WznzkqzBpmdndNf8e0tX73fXHQwL5kXIHUa7RoJZIZ75jPziTSkHl6PMdxu5fKh+p9omfSz
vpiX4Sb6rAAidie4IswGffY7XEymzRuiz8Jxf6akPxIeo6i9YvTa6+UO54hINsmHUCkfXsTALr2k
B0trxx9OnUC+UL25zHHKMGFJ8kalBQC1VT8zE4S/fspl+6y0JSSlJ3J6EwO0AIN22mhHG9E/B615
lmzSaT1qRe0YyfqDGGckTH28anKKUCu2CkbTYwti9sN//xDU4k4QA7bZtwDAYY4JChDY3a43NCr3
49z3KimqCJvSo3BkJYe8HkRt0Paxb5xIp6ijoE8n6KjSnE9U4sus5D1GLvMupPCQ2hXSiuYeYMdo
+/lRAbJVif/O1gWUqOk/IXJGvKzkwZn0jumrw+/TT0/iXPZlG/pqt4uTL3YRvVPFMTdiXoETlWzF
aS33VqVt3Rwv/y91kHYQc0jjWVdi2T48Nm3HthviTQoorN2NyiV+Ct8XkFSLOzICTXtDvbOxhBuY
oofjr4eb8PZ86jAAjmUW8Czcnuxs+7JzX0Xcm4NMZdyNkrXtPUWCVbIGa7PwOFyKvtWgx/7axk0I
hfQXzrdCqyZD4YhM1qGsL7BoIi68VDO4Sck6nBHiIG+4BUNoeKKh8rB4SunEWJg8sGMn6S6fq9dN
GZ3Y8VyQhDA9ugng8/+epptxkaMeX/Aey4gvPRLcmbTYDEkqLYC9ARHpi4oBJVlvUDQsTT+U3Ud0
zAOYC5bHIm4Sx+PwwglvEgpizLfbXX0V/JMe10kY5UvWpylGGH3i6msZJdemkFHjF2wNzhD9N88U
bDDb5L9jZ4k286sCCwxdij9vy+KmeL8+bjGUwBvmbt3nCvz4Mlx3IVnXTeWySxmZbbXLoTycyx/r
P5m6qK6rup+o6kQ2Fta7c5QyxjxBZU/Ns5bhho55MfL1MM10yWhti7UOhEt9o992ZKtmkVVtuVNh
9xML/fzF1igzKt7narAE2w3pJ5mmVe2h0lV8fYnVdqgWOm2454etosEH3LLm834dQ37scjrHGF3i
nW54JfAhw60EGePm8fI4E4+7SKVDPF0N+RNUyxpz2XAYLMtd5ctrhFVNGsKkIJuVHoXdIQ2Xy2MZ
+RYomuwxAH7q72lvugYRPP83eCrJ4GJL09Tzlge3ZtqsTWVzL5c7bWINo5ex/SL82ykE+IuzdzV7
4/phaAoT55LCvAyDiDDTKCosz0NNRProAMfXn9nJGhpyqdgyscWp6TOv+RsAkGM1cMMKgWKl0BZD
SXDfE3qwg2iHH8fMQGURUC+VqykbzLEjo1IB9+TsqhovLG5mcBGQB91tcgZ8i5lT7W3YuG7pFH6/
7YLXr0oOXoCFaBdhwyi5oMxZzxpx4Fc7WmemnGIcKKQVe/50AZeGACP+CeiaNVuIETKEYYncI/kE
N+ATridvl23twRY5ZtsW44/UGrsn6bDk9MqqDYlRParY0EcrKCoFsr1Hf/EWpOyo2yplkFbRJA6C
pr7MdxHNcZKlH/MWWMCz8bBPppc0JQhTJ10hakFWLeMtQ/vAkjZf9GB0DeKdK12hpllV1p69ch2A
izzbga/liu5C6Nn6czCTF6p3gev2C0E+J/ULzFssjthHKCemgDAcIZesXCpKkeVJyIYG2HWmQxbo
bzugDm6ssV0pxKeJBsP0uZm8EWOWni98y+SoDzS81Ge65h1d9g6zxF7JEy7ALq0pZTaVQThbcZNP
lcpS6xNcX76f4A9de87I8p4KikcpEE+Q+uLYuzxVbEfLWUqyIsnWWCfwVtzcEsAj1YRzTBCUSIv+
jzBZpLoxe1ebSekrBjDX1Taz0FLkwqEabPyj3qhaIpcAMtCGw5cWeXbrWJXryO5BpS4pBfWvfmCl
/Hg80/zwmnMzgbkjJqIJry+zwSLHOAQMR9ng/ClwQlVRs+eKvQbXI0s+1hJ+aQhr7j1QVDs26oHq
AgGp5ZS7RijXUisV0cDmzdKuLhitB96vQIl1W5LTWoXYWbVgELNhj2PJAvJiNcg7ph5WUKQtsbUM
oNMmMjiF+7TJ0IYggUPq2dXkH9y7U+TM5OJDfcq1KAyctnwz+KRkLB9vOdxRm4SM9PUjENl77L0/
Pa/s6fBBiS684WzzlHbQA/dTaUkt7UdxGqmrTrH2FKLpHRm48lecrr5K1OuhholbpEjSmFQ0OF5m
3GwILUfSRBwkYF2kHSAkyu9nhdNOAweyGkx6X+HBz3uCWd++zShH79yCpakXYKojWO6NfLtxDx80
aw2eSZ/kpjV4au0EEg7BkOavMRrjiaCvoh/OkpAxNQNj2NfQN96rJVrmqLfpEECr23zG7Uaos+qc
pvBbeAKWQ0AcvARQSQ1qT1le9SK3qMnIhb/9Nb1x90+ONDmxcY2DzDnjtBMGDWaubZMUTlozYhYP
FV8ALmM585vVYSx+naUE+B+uCpsz7VFi4vgTw33oXX46XJk6LRK7n2lOskayTTmKoDcryEZQopD7
fgBeb64d2TgeDWyHfZ7do0I58fD1uwF3l/3O04h7nTzXuPH4AVxUprWRMvqgIUK1uJr1OmSRnJR/
EmyiImzt/DYYeEfbne638wL/l38diPkq/KtUGeRzvErvQ4nA+71wWnRuNpgHGm0i/M5y1/IXVIFY
X28tmanvDv4lsMIXJxCBXOVHYs1CSMsOIJxQ6ArsIr7bMmJ8KNBABcmDszwymveYIER49gi7Jsxh
AVUdDQQkddYNgfCbVPqlDTZuEqtN1T2qQ63qUM3vyhvx31VZ1nIFl1X2LksywdaVEHHJvRdgT2Be
vu4+GdVHm/gaYM+JxlhSBsucTaHQB8rtqG4hPccF9vb3MoB4NT/tzJRtVFgyzTycr9KeHZYOr0s/
++xrnNjdcSmSwfP4/lcelqR0CE4j4T/AQuFrsntycIlN6o9Rn0HjpbrBm7EZf8z/lpFrz+uVNr2/
zbk/zeiZWVbwNttQTU+GCzlqaXBJeys9/43Cygt/n/Q8y3mF4V73WCeqwgVbVrDI03MYBX4DQ8n0
HcQmgs/KaCppO157asSlHmm9O0Q20wm2DKkHsYcm12wpF946v+ucmc6cb1XTJiDjf/2FhweyeBU1
wPJGx3C+lYw0l6SKA4yACKpKsKD3gdn2QRBHnpHXmfmusJvTB++ZtLSDQAkGylSZLbD3LGmffIER
q54BR7mvQtXnho1tCdPB14xnbgmBIHeUsxaFEWiA0C713xJVu0c39jy9EeSrilmOwA9bhgHmCpFr
/JNco58lONk2It/OyvN01/rqactbzJRJbsTEhOXQuKr5cror5YfQA7knWkWA9zsA2c1gMHXNZhBN
wGAGKwI+OdRqnZDuqmsBfljByuFFAQDIntLGiFWhS5D9A2ClbpcHTfFO0PfrdmRToXn2JwBN1piv
vTi22/3Jys67Lc3A1HxCAbWcGHutnyzn8BW3tlDl0ZEAfw3gRmr5cViB3a8HD6MqeLI51CMZ2/bL
tBh08a/tp38hE3WDDhaUJQFSCV99A8N4gXYVzZS58WAIbUXp2ygtu+mQhnq18VA6lXnbtAFFkPJq
LIhQnZKHtCJoQdSXIrWZxWpZWS66yop8fKQn5T9i/VT7DMlQ+1qvxJHcGZADo9EU23ZTajfgz2Fg
vGF5bQ03RKNPacCu2tBKZn99sxLbHlHC2XFgTtbiz2u9BTjfRgVPNwdBD6D2ZvRhljKqYdgeJunS
+10ArtjTXUIh9DctwhNGf4kSZNyQMFdhIU0+rJepwwMthLxn15GAMl0rnQtUrRNnaa1OykIwxsss
a0NLrt43CI0/K5Dch4hVCoQ0FAmah/5LEJYZG78LvDGYjng9qtESJQuLCNXNV/PTLMk4Q3cGoq+m
NqoRHr1xYV3wdBgN6yI4OEPaQc6aHoTP5qed1EPBBt9/6YyRC6LOs+UHiOqADz+CdS4j7tix43Wu
LF8uvpSknEQ7ugtA0BzDqz6tHzoXOKe6Pfo9JfCN/kwWGOtaIhxvz6bhloiXNFZk+ZOpAoWprIVx
5fySNzraJZ0RcQtgdE/y/qPffoGw8D+YwGL23YdEyidWbA8BogEIrFM9ujTVQKm3ZmUV3Jup1D1G
QTjEl7oP5OoKOwT0Ufa4uiRaUP1NgKDglwjtmxuOBXtZ1HJW8KLSGNMOZM9mz6jjW5V8DFicW6yD
pDGIIUemuJOqFLvvPQJivWu+wuM4YOFMvQ1jmAnvjXWPLX+ghiBkHLPxpx/+uWli1uxQGaeVzxH0
wRukkWWIofpZtLu3A1WgRI65R5jhN103t/9gl1Ja9Ez4Q5TLmnfBXVFQ8cBMrDQujOd06e9NR7AC
w5jyfaHvKSh1wLBx4TQZUEDQqXXv0paadMhAZBcwyb+i4sDexjzZnYLHMAfpBVJZhjkmmOYvgRHl
7uDjuMQ0Vj/LsWqKWKjPAnV1pMz3RDbflbWRw029yLfr7cysR11xBvmO5QNYGg5YFOzzZf8iZOtH
g/h5oj59FEIix8LWtBax87UVzUx2wf41dphLd5TgbbtYaFecHPrFfGrzALQr5zyH5klfraMMa4Cm
VAZg0+HS6oW08t+khoTUBoGDb1ajXtnJjdtyHOCsOPnJq1agQbVgBoE4aMpo2n4VqLSvSrADtsD9
AxgNeNUKEFLQbww2kebMzy9igoRofSV1XkmcssjChtbhpUbVAKnV49d9MhyB97DLh6HYaP/vM/5G
Pb5mNn/CJaPnNdJaDkY3LGEBPF+DqjIbYbZoJ7rqefR0FtiMRydJGdSObfUJwL5BOwDGR9JfLrkq
ATyu8/hOmPw08xe8ZxWx2xSZfFSJ+Wo1ZOV1bCa5Tid2Ap8csO278/IQlTO3ERUW67qNtyVJjJ0/
/gIoM4e4FMeNR6i5qdL7gTguCAzPnCLhZZOm3dqbx3p3hqxgARViJSPgjE/muLyCjzWHaoRDRhI/
H3LkKBKGmW/spMrPqS4SMa3dVk82ZLx3fH9RBcZpodZTUUnJeTj+dA19YZeAfFpvXVLff+6kvuj1
ZHfPfmrCyrPqylR7XTArvT87Ji+OMnGuC7bC5/ELm4JxVts+1E5CJPurKMdWdWM2PU9xbS3ZrPaU
+Vx55ZMxOQWzBToQ30rsO4nj8eedWrOTY4u3RTQtX61miKyGJvAjCWKuFNoUfqjG5aJrJCrwjarE
w2D0E1vWluXZlSti5ulZw7cNaB/oEKXwVCHHGsd2aPW6Nbqfo1hg2uHPma4SVgUHEeEKoM12wmGq
mqgB5LygXikutPNyJU5fh1ORNqkVaVqIWO76bP21P785AVNayGkZlCkwgMwaDbyjP++Z0B+jnrVT
t3h1kfjH1VEcUJR0BAw8kdQdxRA4bcmhEUQzLyjfryNZtZKVixAquQvxYcPvSUbJ7EFgY0ChtagY
HagKl6Zc51tSg6ESvICZqk7D/Q5SvaNmmIoJkfzGcYKYN0s4aBtltjKip3qeYAnWigUg+TJbd6Ye
TQvsOGVsftA7MIeVOU25Xkf/V+A8UhI91VJYP5Celh6U7gHnMcYbuhJ0n8JE98Lnj7Y5Sn3hdrvJ
uuSgIK4xHnupJpZRXe1/0M9GU2P5QEUv+WWsHl3yYOtlSLXzvcNrLTXf2+y3c+4+BWP2JIJEr0R3
rPSlJP7HAUnhvG8qwOAzghcMjJIDhGLkO6bB9UVmqO44wee9rJkuD1kqElWZ8ketkduyHVvyZ/Vf
uz1hDXsxofAphAPXqH1YziboHl223YHop91emwXDb97WGk1eMpuCyx4IOyZ8v86QYZWYC7U4k3Lu
khrWrbJwxnOSKJRHEMxBjeJdtVdFCf19bqNf4MiXASpfaCPUlhlBbcH0mFMmeQzgRA2puwVFmMlE
iejf6xC0mFnO9RWbh0LY7tmrJ077kocQ1RRMih+OZbfqy/y9upFmRffr4GSixTdANhDGCC7EWQZ9
tUDqYqTmQKfRH6b2xrJb6E32oPVGJNayVFgPKswwl272GR3XPH4bcXjVBGXrRpC00TMx+V4fPL1W
f7gotcJATb1SU0wfynCA/ESL7bl+wDuaG03kPuWJFPm03n2uM98KyQ3N4NCFs6M25DWcTtOuH5ib
7UxdyNMyniJ2VRzWayhW9jYjoM2Lv4jhRAa5nF9yRP+/QTZxYCQVb9SzOj9X98l+s1h6rMSxIv0y
s0GHdrhZ4WERaQGF27zflKjtbHUeucRYrk/Kttoq2tp5dxrNbQpmTHaWUYzwgxpDMnpuCmNtQX1n
WJw42+HZ7+e7i2EUiV4DD+8In+PLPlrFlXozOqFzMi+2XFh09p9j+idsf3xeTq73LPLi9k7xDWrX
X3/2ooY8LGMsfTUYwMgMk6DuosOWpDaEC4SeIO1b2Qe+fEoF7krb0MWnVs+/u5NB7QmAout3wEUL
rW0PR6NtlKM0bvvf2E/6H0u2I8oy04Z0APPbCZ2d6E5XVoV7CyL7uIcustMxzl+n0UmwVq677psb
04BdT8NB697QT3+5hMDxkDPyBj7lPxe2UMP0W8HL4yMylvAU4atL7dALCVFyhX/63Utunj6uQMkW
QNLkxQn9WNcfqGfHiGc+0d7eWHhcHvPFqgz6uMhMUpvmsFomJBAI4HcAQJcxoz4Dlk2D19kPCP8J
v4t+FLfj7JceKr6EO/FEH737Ij0CbZO60UtOGjCBjsuY7zffRc/mGVCbMBKygg4Hf3bxnS//1lBb
+s2NR9HSqMiLiU5K1HlGyl+4aQEOWD66xB/iBK7E0bXGb69/5r8vxBvzAY5d4NRR8yiB2tRdk0Tz
axUvyviLvwHlKhKnumR334U8x9CedaMcHVxA+u2iQDSmAB1d9yV1CQlg/oixikWjONPm/3o9iEUg
+lXvUV3KkntTJ3eH26uAkYNv/sVRFl+I4XryrBaPRy/BqanTFOde+o2FiLBYM3Jcwb1pi/W7aMSG
LoshwsiddMaG9QTSATTVdVNRahMizFvK61qWjT4F+ycaGvsKxkxsvgbSBZ66YEJ/5+L/H9o81HPu
RSrltzmhc77jiaFyQ0qaVtcXvIY2seCSZN8ACSZj/xc7/TJ5/xikfNfw4N3+d62MQTZF+ZFZ5qq6
lNgsGqm2meAjJQ4J5H851mYwwTnm1tMn01y9R+KTtBZm5XQOnLl4sEW9Zevj3FhYWSfJabjrk3XG
80wXR43Z348ce5ubSaUMFc31KltaGVFB+pFFcUKpxMxky60UacAt5tMj8UMs9obkhqTFVkE73COv
Ld8G72tRV/m0INnTWBtcSzL5zcOm+ItV7cCNmLUxezmnBF9c8AW2pQs2kxWOzIGpVkFmyIGiWh7Y
pZVb7or4ny446mlvc+Gneipdda3mKLjUCRtcG3TsPYQQGe1M2G/08GmOBlZJLLRNS1zHC3KjvPHR
MDfSUMRneuSCby5cJK9w2/X6bkt1wtzEWW0D2tLpeGo+3ZGXJSh+XmljyxJYrRw19Zg30dQnWeeO
L0lWTBN4kRy4Vn4RksFPZ/4tjmjU6yJWvl1+uhpNc1wh8UZ08Cgsu51Tz2uJZFQVj/DxN2svDvR4
nI6KC7Y0Xt19HHULX9xeY3yavhie1fENV5KuYTd+bcy8g31Jb2CWvVAMK1NpSeQ/9rHWJi/aiIGu
MZ76ifMjCHhxh/26amC4j8soSRbAaVVWTdsi0CWG+YZnJFc4XBk4QBH+ZV2ym5LzlS+jU8OYIba/
uxexw1ZCdxCPkG5a4jPUpuoO54bU/YUSa3TilQOe0vw2APo6KcfzgKMJSljVo5kj13Pj2fz5GgtQ
fGWn+vhvZjupozjKErhyHRYgOQ5GdRc6I+7JjtcigwGqWsT3m3IjFhlTblpAwIPT0DRUTe+GHgFK
MhX6MEZM5kXlnh8oqIeZstxVcU+4wxy5Vc43aH+Y9/hstYgwMptE4oqr3zWQqeTiSxKQhA4yulf4
tPF8QFcdEYLajkc7KWGhnzXr2O9Dxgl9nUuYiCZ+Y0NJUkaQdgFDzTl94tXv7uTR9Gq93ew9tRJc
a0Q7XwOwFT1Bu7Hb8twV42hGICVSwTTZxZKrYQws8c9BffO63whyp36azvSMmSR2feuKuGaT3swY
/8T1FAO+viyAlVm0yLf5rvPha+13MKm3MT1fK5VzL9ayWxMzmJk7VxV+cVy4Ety6i4GPYGOl3xhU
1LDxcqJ0oKmoPMAtkARsNC9EvISJpTbuteEe+JKNplWhI/YNYtNDS+s26ByVbulx4rMRaf7+7qen
DpceAbzPs//sQMZcy55XVFvwzrrh80BzqxAoDhvVNbqat1xO83fb/pcXcXz3ZQKwfkwV3PoyOgTF
Gy3LwgCobRcyUfv311ZGR6EZ4Kv5Co1orSes3MtnwdaoyOe18EnTCINl7+9LlDeuircs1WhQwaz+
Py5JsBxTAlQCT8ziVO10JxNa6uebOqS6cS1mPHKPgwz9erOfVJBOxNfSN8c+AjmhOZ8J/P8a7gdP
Libx52x5tfDil4Lz6x7esAD/jN4LSXbTN/h+m1jCqO1USW4JJvNwsdzbvJLFjpZaXDNVTiicQK7R
MEfAf9bXOhSGFnnxDVIiU+RMHxhY+9SO2tokZx769asvJ8GG3XcYoP34l4PpofTpAj10iAWi/qX2
CXxHTT/TkmJUaVj0LSHU5DW7DF/gTWMa0i2t3ojbqlIIwElVEabPJUgX9C2rRSav9wqR6lhbHoTr
bMxtsvhDUUO3d9NyT04cVM5VZy0tfXqTcT+HvyhfTptyjyTg+CLIhnyUXsqB4M7JKBaXqWoqDTDJ
t2k5xd9jjPXmewU9FrNoWEZ58zoxgky0p8/fLOAFL04u1sgULXDXiO/BEbEus08kryZ5tAlNVtnx
35X46X1L1ZnmxSJLVh1BPGrMJOZIwYVg6Hih8dOou6ZqYaahAf6tSG8yvHwvhwzAK/qnifgOzad5
ZSz3HqFSupJESEjv56b5GqSv7/xamQygXDNxu86brEgCAdxDKpeCKeQQlyv3Ga5YPOOPnoBp3xfr
ELJzRLAA85/Mfg4L8bXgND0XtFgSHde5v5s/FQbduLqdA8i5JWyC0Flxavj80tY5We4VWXay0Quw
8f4WlATmB5JEYxoUESAlnWo4Ym1MjJbU5h+2QskvM9nabD15t97enXvNCbtfRQYUOe3owjhsHGrC
IwJqY9O+8Wi2rRIashV8RremXqjNAX2ezuCLng7oztFgXqNIM6rAJaBOFDkgWj2MMKZApmPjbKzL
IoqAQIC4/ByZmBj49YCpSJNEdOnLHw0HypxQG896Kwfy1YGRUIRTVUeZWByCt6pm9eS4eD0kTip2
zI/7OED9VTG4TkcKVCSYIVXcSo/YMtvapoFcvjq/swAqUPvxmJGdaO3NiyMcrFv3GNuhR0grOVzA
/11GsoxXSLXMkzgoaD+NHQN5DU1mEhHwHH0J62FNEPkLwBgtSgoAYljd+HOGK9onCDlu+84V3Kck
ZmZtoxav3+IryjAlbwWjD4AxP2DnCWj9UvWWyHO3v9JFJ5MvfL0wL7KMDjuh4FeFNeERvkBSxa9I
Cjp/6ZiUty/0VbYkbfB1nJBcWrHVOCV6RUXK/EdC1CUIzmrlgVEphi/atmbiGX489IZvCPdJzWAl
lyxyZ0fsldjJUdloSliaV0gIqYdf5ukNABszt5/xo6qAUF9enUwMpH66X8KtOzmXkrl2+gNV92lw
DEAsND8r8wPkp9/wnJnlQrlAC95wwY5mZcDBeDb2qhokpmGalJyimuSw6lKrq78FJg4D3+Ve49WL
2q7lxcss5X0bJvIoW11eQH9SX3JYINQHLRJRWQUnvPDABS1bG7x/jU01he1bQ9+hGc22dSrD/RFC
WeRD4EVZzz+Atl8t/MgECG8BDlQFGxgbms368Vq9bv6Lzp2LRHIu/GNQjh8NWOwN46F8m+8YdiYG
NnBcuj+TKW7Ztf0plFmUX/a4b5dIEhuW7gd4zHMiLTSMg7EZKnl54qRUZywMFJ38X1lgeJ+tFSlK
s8YBNzaBNR6Fr9YfsbN4fdpRmXDrBGyDrHPbGCzlQjshOUczHAfUMozt1j3FWjqtzPQ/gpou7WS5
UrbFigJxCeRRAWt1+9g/E/u/n9iAL9B2rlQ5YaBYxgx9OPko/Gd/u1f2H3mCW8//4hiMJ6jkVKNe
KeGA1YdPA2UiWvU3keDzLwqZxggP5wQ5mvPi3tadijlp3q2Gx5rXZ7WpQgjS8ZdR3xdEiYE7ZOUB
j5iKXUynaBdIhAdTxE+JWerS44kVjCGaaeE3048yiHkcv2uSn3lqsrA7ywTcX9dnNipn79LLeQyr
a1ksS8nnpURqhkWxaqCFPBtIVdZC1VbtGHWb5JJpcUxtlqMd2qNMYESiiyz8wsQ6gDlALYGyF9UD
MEuMGvAPhtLryBHCeuN6ZLLQ14cMsJQ/BX7l7rAkhwc8JMEIdpCsHFNZGJMxy4ycrlFz5JiB/ZU6
184CdXysk98RNmOfe4kIRVqMxExs1kJMLxIZRM5RikWCsTlzBUa52IDLf/IhfQcuCxaRfkXiFw+R
Mmw/N4RyrewK8XMr/Dg8rSA7AO/+5cJ4/J8u1a3kynSxXudB58fnhqSjmlvrsxwqAK3o624Huc9M
+TQ3kEBn1eiyOJYTYtHtAGeozYJgHI/Sy2usFs5Z9OPmi3h4xwevV6FNSnmTNIQqhuDLHLAkaaKP
2t+82SCaCwfbr0OjBLtTRsi5GuZ/5atjoBm3Msw9tTdICgw1vwjlNVhBAY5Uz+p11msG2ZRaSpQQ
SNnry5DYh7lvGpOYZ1toHfcD2OF6h+KaoWJzR8qMGFeqlY2BboQJgnHuks1UEpiX7uYHctnvWEjT
tXjGqjpHg5672/U8r9OmnyeJkDw0KkH2bgY/GZVsXP9buPlKhMIayVm8rSwwaSqrLVAxSwcDLmjR
JTqYo6mMBmITUpZANeD52GEQ8s4UP96U/ZOVcnbIKMgy0hAwrXOKQlhEVJnaBTbTPTsHaVEhg1nJ
fOqys4WpDtQg8vQyA3Mb0j3IhdCu9I7zwmJ6pn4llRLUzDBcETJVJGi806qJ0Eueq7gE/CUCT/Y+
ZTw/RsZFUt/risZRESfuuKk15i16M28gXRb/Ifvxmb5Sg0R7vCnOq4o+V3BzkKthS7LRbdXjSgwr
ntHSxJsGLlhCt1O8M2rK6OlrGgyYsq1BvDYOti2HQPtG+aVubJn4pR3WSFVCoSLzKyqa2SFxmrCl
HdiMcxjDLCB2WsNhvroZwqUjsJ6qsTHVTiZiQzI9yb/bEwqCx1o0gRda3sHfgkIsiGjBlvFP1VkL
6gW0ZcRLzyANNplNcqYBC8bCGZEzGOjLWc9jxQRusJxSKGkDQxQOwqS2FYcSlEPpfm+5VOJJk2gf
LMarYc1EGFPotaLl/aD8oJzbeb3VYzHRAOfymVpSVkRdH1Xb2tVL/3cabDvfPOtznlS4qG3OhU/u
7cRfVmqtWlHCF84ofqf3/9cDfSNfYVzRfwoecbyQk/Bl8hFN9HvqABi2Ys7RA/2S4s6Ix/HYhMQo
dEBRzVBhQe5sY8TZCmz8yj79u/T6xt7qQa+VXmiOxfYT3otsxQu7X77YzxnJRLY9v49UpXnpbZv7
olQr/zk4o2oVqypt07/cyU0Z+jawqCwSZwPw0SrqQQOX95Zx0ManxKuOrXetA8jMsp3yVHJmLuwl
s2+sLLWdT/NEMkdioNjNXli1Pn4M0Vxf83ni6T1KOyRhuhWsAKVVjbPgpkEeeDo8ihIBkL4n2B9x
a/uSqC+65o5SD3K8nR2GsQpcFq6o1I7fsc5V+jaG4aKU09qz7YtyAtRNB+RY7ymhO1BmlCfRKddI
BzyK+O4nm/9+8SOVT96sQL1qtME65R1J5/JaF9eCLEvQDEOHwDmieH/Q4EYjRt5KEf6MJ9fPniTa
W5RCHJC5dBmQ1seLZb0IRQMxnzP5/Hwl8UCUx6VmWfK4HqIr1LI4zFeGPZ+n6m42zSBkIYagTFWC
w5eiEFLq0wxHIjWTGMRM20AgqnaRqA9p22Uos3jv9yriGQEh+hjtcysts711jcaGdkyV3tNGojUc
7rIkoEQqYr6kwuyiZzgyqO72+sagFo917jpc2M5bc+xCEO8OPoHTTUaPL/usaw5JTQ8g7U/tnBul
95nCMyxtPyqp6x9Dd8MVu4hksNI04ZqezWap+EF2qNK3z3K6nLK90wN52+vkCQiebtsog/q9OpAq
BOpU+dKGgTekWFGGag3iKFOK/kletDTuMSvLCpfCRXpFcAShyjA8Zi49qCGcCmr9FjXucSWp1M+X
49J55G1jK5zXR1NJ5g8e0cHSTdjljdOPUKVRc2NWeOWU2ZqNPqSHk5AVkbiVoIlcTT8RWvwPuqKL
LOupptCC+gIbUMYwPaQkKjaYZZtrap1Re3jBSGvV+iW3EKma3lyKgM+fAzpFh5vw3JDD53FuEztx
0rc7gVSpSsLfU5fbmp76Zr270TQWsf0fESDQFjTpsQFC5hDVhlCrUEmnevdPAt28urRPdbHu+Jct
t0hxgQUuORG2sJvZuPToFEiReaeoTLvoudBzXtIdk7KEXzV0+IXttd7yXdpfVN0kiduJSV5CvTlr
FO4cCjlV9zdml/tM+/HIl8yx04bW8B6NXFjLOhFv8IEG1bx5TgnJLrn7dNO9ojHR9hBZ6B9sih31
lHMd/tGk6zsvt3vqUgMTZDGG9xh6pCp4Fue5M3VD+KVm2+SBelRvlmnGLuETg5RkZqqTqTK0XjzG
fBSIxSrGpffOiBqzRSwNcNPZ55ZNZrXesc03+69vFFAUn5ICn2ilVfTd8oANMvkqZ54tARIVyxnZ
+K3aNhCGuCTyPp01SomeEQBGAH1Wdbm+gMzDVBx2nHf/UQDl+sBFsnQcTP8f+Hqwem9DeiuI0SDF
u7vJQp4/dyzeLQRVJRICRTdeL01vDqS0u0owrO+ww40/dKCio7bmJZv/conW7pEXwLVF2SH7gqsd
FWbNOZyK9bb2Dj0CsCYXDdUvQxwldndRPBcPXk1Gym+JOvgQXIQDvjW3JRFr+6uR82ovH16MZeOT
I5mw/gfm1a6IoiKsXrSogMHkRhUh4BxYVnU6qSn7fQr26RP3r6Z05N4VgXM6yLff/VoDfpQk/Akm
P4QcqD6PPd0d6BRsQ2WMjcMnvc/E13zF4E8uaL8KixWCcq6XXoQtqJtxw38O7bCGElqi1EG5SY+W
tkMWOAPzdk664hpVom60VerVPL8EqeCDk+TtidBHAS5M4y22mqJ6ypf2QPvZ0fBq76pwKPObYZ2H
3+QAhiDPrPETei27CJVclsT4s/FGkki9EfEuuprUcBsdZ/1qD9T0nTHmec73p+iRlR8sy7ZSAOhM
y0HynMPMYenq/FM1BiN5fA89WP36HpH1SRqC49AaUiYvzIwJ6y368JluNwVzBpdrr9QxytytdZgq
8JdHsL+TleDkBehb14I17y71PuddjCQTz9NFghjPtRb2QutG3pG8rOcKsMqDcF1f5b86ARRYn0K6
/bwSxw6Lq6ln8JXB5N+OJMHWwoauE3JOel73JztTIg4AR39EYirWp4ESWojxF8P0WC3PklKdAMB6
8fzTN5HtlLOud32Rikbzsb44sgtF1z1YwtRjU4cTvMF2r/guAUH9uoZNJG17wx8PtzOvgp80cO9g
Ei/8aJDPDsQq+6T7G9TzOtaAVqexxjJiLKLdSjL0HXus7kdAuBnsDovOA7OxFHBSRnX49d2oSnjn
NNvxdAQPCRyo9GxAXFwyTV4U574jesLJsKX9416A9tfhet8AxEILKZ7auj3GmXMcNu6R67IIVtvz
VFyjnKnyKzxbtT/bD0IP6LnWrkibPbP1LgK0RG8F9D6nc11utsXWJf50fJBlN6EN8UGJlLfOPxOQ
qM5/j9KYIIrdLpU4MKCt+gtp8MaDUTQSEPruiuGCTTkL5TMMkgsGLCjfJ691Kp6560kUJ5A/aQA4
aFA3ZNpewu4nb+3XwvfNuPnec2YcS+ToOKuPRU2ikVJgj6NKUyyMCBdMevYR+wZBvGBJW4QhqV77
3tApZ3xjmh66wxSGlTSqFNOIMxhCN2FVkKdvuR0QRzOpoVDxIX19035sOoWoG/NbF6pr/2ZBIwiq
XyJXhE6bJg367il+GzKO5Sl2yhg8iik4WsAagwM0CcVvgk8Q1w1UknGhtKSnNMZZml/fLxVtCqkQ
XIDXWKW1HQ4eJmHFyHOAyXaa2LRZ+MDDxOIq6mxtuL7+DDkr1HAOCxv4TmBmkJ1YkO6DolWYBfTR
YJhNjsw9RfA3AhHxJZpQ70f4/8MgFDJ1oZZ7PhbDHQMNUC6a4HVJdYlIBVRRqhAqKKLdYDDN9PjI
N+HzV9rjjiZunKbjtGTBlaC1MYHXAMeuCSvR8B/1uDTbXOA1FV9mwLUBwklR10zUZiQ/unvSK9j3
032k6W00BABnB8cXaP7q+uCqBQzN83fZgOJq2J0k7lxsYS0zK4COnjmpVaHH84wziO3efj5wvBpE
Sep3gRlyHfvoU9HNqPdvPX9mYA2IaneL8bbf/hAGTFa+RCUis6+rskohw3EM74iZ8EocVAWf099a
Kx2bL470LJ6F5esyjGL8Nt4V4xituvnC6asGvsKbXON1vh3dmK77YFy/dcWq+oFgmyGOjEl7Ipfn
OXJVdfPBB5qYuSymu2ErvHgcyrHvkKMTV2hjY/8cVj8sYwlSoKHgf+b+zwyN/JHdUDC7bn3q4000
ufIoOSe7qM1B4i627OQAGyDwTgClbsuwpHxMY31ET2yWlh5GhJm4uv2FgZT++hpaFmsXWrV33l78
wMnCDpj4v12qvIbEdNQmkqFpvqIA0O5nO0v2FJ69g9ilthBKZ9NwvROIbFW6Kz1kSnuJKBagQkjs
wLdQhkDV7vCoBGba2UlZJQW5KPuBlf7/w/aakZ0FKocdB2Q7JeZNQbDKuMTqiq0WcsIFJ8ig6Bft
jcZx7DWVeBvzOd3SijPWKMQX/f+Yfmfr2EGdixlT3NWxWInhbQ1byOaEAskyUBDXg5VeK0nL9o+S
0DXg3j1N6hzP5J+FNr29KG9TVkTiYeEi2oAeHy6XBA0nkCPYb23R++tATUV/2HjWPmeHtaCfyvaR
dcTFZS5iQQ9gtO7cS+iwcv4Oal7V1XR4vYYzgv6HtRRoFZx9tAFfFLHGAgULMpCgHGckglLlvHNe
4z+poNdDVBB5IQiHo9k8WhoXQ5OCjNgtsWUYMors8E8Uw4e1QqEuALCdTjei9jDMQQjJ7MFgEwoL
dpANHt7aAxTm2Xv+SViiUPiyBqgM4IIDHSwuKB9PEw2yAUbs4eERmVyEVDsbE+XwORvzS/uZb1Mw
nHxEkSTjAbF19RAaNiPjI2UmRw1INWxaRFI+hElIc3gpKrBh33P5W8TMRb+GWY8erZL+lZ2txRrN
QUF7sNwOcW3iEYGAm6oje13g/jkkHhrKbFeT67aEV51DkKvsl3AgzybPv2gu3nMQHx4mEadaLJAA
sIpWCzlLXSXtpiRavy0P9d9k8XkBMGj4TjbriSu29EGXcR5bHjkOOhWI5lnxKpgzZkbgaMHz74x7
LUO9xSpwb8UwqQvmyiCD3l9JpETd3U4JpoIfUMHhnQdxthfiMxb3zykCHte+QtI3r8ytuYpjS5zB
jTiGMfQLQHxTCYjncfH2uBz9z2pXeKYeO02VR3WQqsrAmT7YgqtEZB3DNxbJeoqJqlrL4Dj4JsWc
PjCY22j8qOG6OuYfLFGSHPqACaq3rfC0anXCNMVqldfjSQMvph8C3RzdP1+AMRMfGyJPCSsktXyW
gFexZh50O9JzimBxE3CSsCy/k9DK28llSoitJqel0auKzYUqRhVrBTaoqbm8Av1GWPCll/bLHEle
/jnfLnFkNUEdSysQygQZZIIE+U0XWPhi5TbW+ZycxKBmNNwdqCnmrBW6l5/T/Kl6u3TWZprnfzcB
DTacXqjgtBQxqX/J3yVATYSE57n6OcOwZ2XhUNYp8rnpvAUqhXS26Ejzx/UMQ8Zg9lctGz1kxXcu
NCru8m+/jCRtIFW3jci/1liwpUKTtmTUalllxu4Z0uuq2JJ90mp0Ifrih6Vsv/+4awuwx7zKxbl0
2i4Acp9eq5zJu6LlV63+wr/P2Xpd2Evlb/uBjvIvDlhZlM9+pyajhvQdSqO6ZSZBJCGEHmBh7WVN
xcuLzKarytm92pvOxj2aIx+ptfY68qAFe96KWlpd+ugrpR7ODA4nuzzkruqv+L1Zu43YzTJaRVCP
BKD5t6iD706CXh8EwQTYx6OUX2jGTkqkyP/zA1MvlF0gAXJH4iABFY/bSQX1tV23jVSzq7TQD/Jq
UAm+29qQGwXoApS5UeRxEOfUuVKLW5sSjaKGatLSE9LziI0vXZDAJ3OJt8bef3+dbIOCWIpkUSNO
kXN9Nhmk2k+MKE2YggTMK2lAN8I/i8I3aSqm/GZF5c/KSjnv3j53lsdjGPSUZMWKUXEndI9Zcz3Z
wSPicJpaEltQA4wBNZemGB6vzwmECvlhWYMIKwIFqsVh0nnj/zPOq3Q5Dn5k7j2Z6OpjXDUjHrg3
27vB/jQ6O1JB6uuomEHVhbdIMChuO2GpoA9HbAgvM1S/UgTn2wMzfIMuAKXqpfJwJsnCJJxCrtPE
RS0c97d88sEHQ9uujpLkfQKBHrYOAdpM49agop/TCjydtPKHMWC8w7MHGILV4dD8ceG9yvZ3rQgY
KU6dMvn19SrD1xrmCeSxcoLV4qOybYAa5K/f7mgV4O5MxUkOxI140l0n6CbZg5ZI7md44dvfqfiH
sWuBl2tPRdpqS+G+Rdqh2XfHTYrh+e91q80jmR1p5zmB0RJMulVO6UvUHck7pT6shP8UYj7ilhlq
inPoV94z4js93G3M0rDXLNrk77skRAvuTxQZEa3ovjpqrNoZoA7Z9YlVaPUC+NhCq7YuwCUbJ4mO
x8p+5yteCiWts6bGmtOxrkEQHG7KglYHogexwAw6pVhXasKDKHFX9OeL39c9Xk/qjpyY9YRuWzsd
gUE85HdoxKy1h9O6erpcDEssLFgXJLeDJoH6XIPgM0fgf2qllBULS3Gcn7Co20o8qbEG2G+yhBmL
78ymhPxrDwVsx01zLCOHf16A9XsbQjkyHglFmlKTna2+1FPAQXAd94Vp7wR2wlDVJONDIxW6RF19
XXJoWZ7uKihFNpiYzTdj807g8/dmR13YFYj3mzOWcJmy5bIL6Bh6y2HUIMxz7Ku6zRoUryWVpiJH
26O85Qp7ylwAzSDIjJb4mILpfF68yBJwUIcBncd38CiFZAJao3yXzjk+FTAtMC2nTkP43rX44Zkw
3o1HMoxMTVS4+Mp62S5QnTJTnvqS/JFw2o1+NdsZVygG4OiBXB1ht1HGJAv+RxChP6qDiRnWnZQB
M9oBa4SO3HNJK77hWFICLIiDl/1nIuhVRVQc5zHdrye8EvJIUkBP6qiwY3fLFng6QnVq6DOz3mg0
aEJo6bUG1eLDquflc9oLAWvy3pRDGidOFxj86APr/sWVwyg0dlg7q4zh1/gBW0f3noB7iQ+6mEL5
+r6Y1S3BSw0X37e3u5CWwmlzAXCNlqCINVASFvrSGrJ4anjdKVKR9I9iFbYJe+gbyeBoP2Gtohcw
4Vu7wYy4rBhG/bSzD4Pz5IE3lJMutD8RG48A93MyqltAtZfun+DDNpCI8nIsgS1Eq+C98KZtqg5K
KkD49r+mtJ1ILumIbJTwq+UaPfXksu0kLchj975J/BAmKFLJoRsz5VovR8rDN+evdK42K93IovVM
m24rn8RdokjqGG6R4ujYuR5I3AwgT177vv4v7U1G92MdGfUiHIN52rRSdo4t4PivaxasLElXFfLM
8Bj40gx1qkqd9FBT1brMzvU5aXZ9sQOX43nWu5qBEznXPTPWzHuzfZD5soo1zrinXnqoAx8Z2jQR
F3PMK5EVYicD/NbWLaiCUYvW8EWI7WWAATpWoDj5vV1Jbh/+pErrNzM4xxfNbstwGiR+6xJC6xaA
ZNUh6svgMQHdglHii5WfYCmtjODaZg9VYc+Sm1GCnpp0rYHO1d9AbAidFzK1quKWJI55wMe9S9pq
ZrQChrs4J0zO7oPqoU6LHUjTK1IpRd0w06MIF/s8J7Y0Y/ypZZTWdsWAwM5eOK3GBO/YMktVFcre
hFQVn9hnUovnGQh0ycd3WR2JHvMfrfObaSEeT/pfD50m0lSrG8ArSgLS7VhWuWxM+Yo8M5KBnm3n
F1UZ6KLjZbkfSOClzWLUGEcawZJ8BSpmVY4Y0msSr8HHExpw3NEuiuOhFfVlaA49Fh4epsSgfR9f
ezXo9ymOAKdEYiyhOZRc3JQXNl417O7MHEquyfzHqpSpAmunMUIIJrgHRidEWOcE5GkK+PIMBDWG
T+igZXLo9x540IGXF9Mcij+5UgxHMJk0krgKj4CaQ70MiyYS3HPsEdRtYX/4QkQjNhwebx/nDpKK
O5ME5ax7P+JDyp0pk5Dea8DLg3ANGyn5q2ZfqldKNahI2St1SLitDj5qg315JLoYVOFFM6vuUBkS
eo2QU0FBqiVD16bOa5AjJN3W9SRv6aEjx5zIf9809PjeGt6+RdPzrdtpxz+EpFQxVNArrme0YaTo
ga04w3HvWZBmyloJHGfA4N0S0gIr6l6RgzxyukY+gB1OejGRKBCrX8jgCyodGxj0D3a93MYnkSjp
YefM3v5aT5WYC40M6AcAVHgJibMOLOdBR2P0tRkTDy79nmCyUJY6gO/uH5xfcCKyqv+y8u+n35Bi
K42k9yjNJ20WeUdnyqrK34WCEDlbinx/mrDFcjnS/dWJnKgns3eRKfKYhM5z3pwX3fParBNvwalB
hC0H5cyY/W6u2l+N5+lJQPTPpUQeUIGsdiFRlzTdJWt6fHU1o3kOukEQiBZlfLiR9m12nCagFQGK
zotUITY1hhuT3ZNKhi+0lpBpX1j4Bh33hoUGZtWmu5rGIwpT9tzUNsS3yF3gAZEL4UiVPYAM8mw2
RyoEEW3QmdH/0dy1HiFz7DTLorG5yRB6FNrqGX7ii70HrYZRZ6PtfB7M4BiT8s+h/LGK1NKZRBmY
bxUzBgMBRTpTbrY74yoIYnKaT1Ex4CZNGnQrhcq1J9fQOYkCjnxwHGuSjxJtYVmQWevkdtf88PKU
GPnEMRAcKZh+JktW51EIRjrdD3eaz05Eoztj5cpZk7rT+0+QggejLTrEX4Bs3ezu5cRL++l4gtMn
3SzWBBQf6z8BueHkXZwfpC0RheSvE9UPvtOPR974HCQT+YYDiV2dZ5hfuA1gCiyPVRecsBGZJIOb
DhhGICB/MJQQ5rmD6cVaF4u6XcLsDjlabDiu45CGtbnnjVNUpGFmfUuo9XNbYj1WRxdN88mAOrW8
tADiAFm7yQuC/F5D5uFT3qcrogGaY+VR8vRU3/EWV10rI1vyC9wQfI+wgmRRD+szhD8p6NA8vt2I
dNBqHP4nbeS+CUN7wAMHDFNP9GYX7hC98HGq9feGN94pBlE0aVLFrd/5ay/VmO/+5zamjYkqZwrU
N0/0Qx9Xf4PA1x+v/k9FNmRqcY3p2F13pkJFPY93XzpuaYLyZO42AbbubsWppthZQQfJMBXQDcuk
m9jOx4tDMkHW9DqQfmZ/UxeNESbUMl8mvFJR2edrO7Ep+omS9Nxj8Kw0Gkc1w73EWFQYTLfzoN3y
7CYd97vZK61kJ4rDecx0edH5TsuWLAAW/3/AftwoMxvcW3UVX4VnkqzJk1pnu4EdXuJgPIyzq8BG
9qaf6uJmBTlVnewQfG3i2dMvdiZBI3oI3n6KyZBUVrH6nHXHFmqnr2pRRzF8z7uTI5t6IqwaQf7/
2Zno/XeQCzGD3+SSuo3kSmRfN6gGMzQTQYgDGno/yxq/J8Cx9y7hYjRZpyCRpw+TLTSskumO2Kao
lTnrsN7uKCD++3266dS+P5dhbSngRHGKGp4MVAeER6uwEHj8EwIF+pIu2v/Z1iUD8WA19sWaKtqo
xb1DZmlWcm+77gHMJ8XUZD6cSNr2fW2poJ6uoSbgKrZWgzWmaAw3HKkTbUFDBe7nqyP1+9eWvR9J
ACHiVrH+KI5k9ZEaxlGEkSYl3EWv5VoG0zYnVDVUrIY3KfxMXF9I3dEIpCJS3ErIowFlgN0o/WL6
Dal9i/LYYWPVJyRsxBM+9v+s4dFZwRk+K8JmuMwpicK0Tp0dWQ3em3M8e233nFutEg3YeGU4fFRN
E3YWJiuWDqp5toffceZI+KLV/vBYC377xZet7RvgF6f/HfhtYEjWNROMhEDhzwiWfKsw5HCt15PB
IpNj3NBbpdnu90jQiHp1bpR9DElJPu2XtDkfCyDf/fPTw61kCpXD5xD4UvCwiCw0DaiCAPXId1pj
h6xWELIT6PXKlNbYt6AYtW1A1YZ+HkJeZUatInCgom4Kvj+o2JgU3hF+E0W1Vh+gTbNanKnJOuzQ
Jvg4LDwjbtfvuz976iJiHF0sNsOxU5rR+T8il9AJnL+rQCNquMNq0mW0KfenPQoK1khVnOmqMedj
wbnvionhmgjxqiAkhEdV1gSh616Use0PJyl7KjE+iHg7o5olgXWUPPDWyMAMrNyJpKY4Uk/imJiI
SJ+/yUMzeEbDy+jscGhNVVFoXvLqrR2YaSzxxxW/REQdVxl3WJR1BSZQ0GUuVR5GwVijwcysvSUe
MW3Ud+jppTnEleZO3ZQV+oaWDX1eDdutTDH4+e4WNzQVj+T2SL0PPdT8jyzZUN/YmtGziaNFzF0b
jf+n5sKJm5lqWIvGblywre6ctfEftvID/MnOQn9hn3hkVtuc3I8yezrjqMtVfAMBVfUcxq2MPFeh
AghHPEJ/hgkTisX31tXoqCe+5fYN6ElLr0OWXmdyvn2ZRpqfu3iLesIQMG3H3i1oWph4IPgAqdJS
a97tJSP6OcFD+w5Z7hfz0cBTP9RUGW4HIq1uSups/Wyxg51i38ToVt+7jCET1JrKOHjTtZ4c3KrQ
4nzSm4NxeCQciUJmJ0cotJaZycMblMCxcMvhdNNWR/6csZRND296fluI1YQcrwaFMw9uJHfAk64U
AarmuK600cV7gxtsm6ZQ1oZMnbvWOe0ZkhieWYYw+5n7E7TMqhMYlFjStG3polN26+5nPd4DnjZv
XfmikEvxFv7IAe7t4zWyj5cDB/Cs2YcOaQwWixZIQgVwKViwM30zBb6PWbNUSMLDbQr4ffc8clMu
L7d3A16UbBOl5AVtVyi7pDFyIgmDKq3SjjPrIsYY/ShLUq40cj2OTrVjzHTiXxGXCJi+CRhdPg8C
eBgsJA+CFTuNqyCrZWDB5aIiIT0r5hhRz5fqbfhCmmZ9Eo/FRxbmVKOleo7bYfLQx1gLUjEcqtHs
uTnVe73gFi9ZCrFbgRU+qWzje9+uZrTgXUq+pCFqYz5eHgBbMY4s3fgKcleca+l3ljzvzYVAe69F
ex92jE0ViirINW9NMSM9DOhKxH8bwrbbx39hCR2SioYabkps+iQOdMD6iO3OaS5SapT02nHeSiZ+
EJRCuObfAk0FWqviPfwfHjREj0y6bu7lgL9uGQSMcUe+EmX8ciuZoaGCPurMNO4TUvCwJltylTGl
3EVphtqSnJgoc3GUu9jemw+TI8vGgWIToTTumptsFq+QYHxy84EUfwOlKhkMoRy8nXQ+s+blzrTk
V5x/mybaw7VobipHQ60yjOUh0AxqBm8teL79Uxr5ZpWYudovJVzy2nl/F8x9xTTKWEOJjBXTmGNK
mNVJVOd1Pmrpu9lbDTN4rgMYrTD2rnb3X8CHOqXfj7D1JsaR3ImhaxeYa/KHZROZfghH5xoICq3F
ZrprSvBtspYKVIPwJ2Vdi/BDXsQJxb6tmpA2Cen4vuPCfp/1p+QfuBWBkL2Fxsk6ZUsUJTbiWDCn
swAOBcOks+X5BltdICHPYQX2N24IJefXEzBE9NHOY9l2EZ7x6bWO5exMRi+gxcgOzGbGL7iW8rf6
1k+mVhty04kx4sRNeyi0x0h6Q/N2pXG2OJJ611uB/hgs9GaCDDCm//oOzGByD2QpWY5z4kh+5CiT
Ab2AkhsDxGMPfObpe8stT/nCSUGoNNvJpRuCRxVs2nq/cDB977phkcAW5iQL8+FynUOh+bYqJbuH
7iPDP9iyD+/+vhQ+QDX0t8EFPoTGbrfVJf7uhFG7Yq/r2pzg7tR4vXO11WBJn3nNg8VEIvvbeqrm
b1jCySn85o2XSxJt3UbKy+ZtuiHfne5AQrQN5Vz5cZBoPJjZAXNVSUaUnkQSYR/N1mfY+runRFVi
CnuZlZVoYzSsGenUYOdDNt0AaHLvsjNNWJwu4W4Dj9cBAy/XuT6AMml1MvIj5MKbbVDu48A4Xcp3
mRpoiKsySufIF6FXDnc49kKiDn4QroPeBJWITkP+2LQCM6fz6UzOeJ7+G2IOsXvv4QPVNdV75YL5
gqG28BYFORWhFJxSaqrECPi9ROyfz+67FCike48ZwQSkb67DJ137OgXqzw8rBZ9WnmLlyKAzcZsZ
WNu3TOEOTd3N1dT/45xwqPLlA6Rp2gr0H/g+D4MDaLnVReT7Y9JhP8CEFRlwEjtxiro5VXS9P0ck
Q+XS6nIO7WAIbFJ/+6Y1bOf4QhS4+YSbz6a6qf5IRNiNyO2etbg1o3053pG4QJKOgvMOWefrmDT/
Z8XTr+fLA+YaC858Tqs3c2OfEOHIz+fLHUht61swYJoKkitVujdgFRelvAbxIDIdbOh1PyjsmF66
sSZr7qoqp2COG3OwEoUPAqwOC+si7/QtTWZwMlHb3tydD5Wj/nuI6ocwYRavWWGc4X21mbif7nOt
l+6m2t1JnkVF49IGMHWwLlnc30ODcxRMjxSiIr/nZveSrN09W8wEqPo+lCNvzZ8IYrJSzkKZ6bgk
tF+zX3uuY77cwtYiLA1dxMNyLFxXNAV3N0C3WMGMUL5pU9HUVzSUXG/1/p6qEO7zI35WcoVRHtI0
lBbOL+61NRRZQ2PweBaI6liQbr+22lBRBlky9PMj/JGOn7p4TXULbwXA1zy5pTJUb40VudFw7q5B
WKzygFU/mLDWK4y0CH8y6FSz2W7NS3HKDhEPe/H1//DiveUdc+QyrRt+0m4KuMm1KE2VzuO2j9Fe
LsvkNATzlvtCHEg5O/APOjibtZhBCceTl0YbgveRUCJONZGVBQkn7sMzb6A8nHsefSDtBgkTjW1e
VeBJZIEuRrRAgHLJhePAoF3mjLNe2YUmPj6Dgpqvy0euqISnpz9FVRptcFHo+L1CtH2PfTaSGAwA
qv01+0zoCJTUq/vWyYo1dx92DX0/ubHxhWj4ptdQE1b0p+lXlmyFlJhnRpB88pEiudKZ1OEhvfJf
4SMbStA3/atr3St594thXF/HncxMVAY+sxVYGEdwKrhaVNkem5VDUsga2cqqylolxQU4EvIuofqJ
gtO2ylEMwSbc36l1avLh69wknp0UOOpoVp13T+9E6fm1+7GvUFc7zNa9LwURrGfxWyFDA3ZCe4ir
lHKI6VTIB2GZH2vJjo4LopCf778lbgN4p5yMFgqNS/roirnu4qcVM0dvq+28VIWGGtgcXRySSVHb
k+BN+XPMQGYTkP+ac/ffMzH2bpplq4fPFbHSI3M9m1ZeiYPvvlFYoZZO6SiC8HiZS7zMH/2gHsKo
Qh7tyv7FbjQojUlJp7J8cjHyK5SQ7l8EYyibMD9he3epWpRz07aGaY1A29npFdxajfDGfnZmdKqp
0fTgyMZLuPXRnmKscrZ2eStjgdVrPHz7x34Nn5GTv2rYr1oEENd81sJw6lUBV7XIATCjlWud6EHY
QYpI2nO2hYkgGqdQ6pP5yhfZAzXt4shaQ9sCjO05MhyoTEC/K9NLAVwecK0UZap+RgOS33nVa8Ds
aqnjQyxKP2X/Oi6oSVLTuTLUafzNrcMwN1wknIH3ThbGlO08300elSbI8ObZMfGiJyJnuYpZdyyX
a1QFUOAdfl0b1ZzOx+wbpCPHypjkucV21Qdjl+UOkxrpJ4vz3b4rO3KIZJcHjqS+g4SF7oY0nLyS
9hgdHZHxB0LUqI/JO6tSN9Mg3SIwdDsKZusToU1+floEeNWV6nKeusCQVknq28/xotFK26UZ2bVP
sCb7IPkzRupPgdhEM9tdCNMVcJiguYXn+EMan7ledEKhuuLL9mLmW99GJn8OdqS8spAB4ooqZoVK
vDZMIBkC3pYZDJlOwoHgWARck93CZ509aMO3Y70uQLXOwL+Et5lNzXKSyfeSTeAyOPAQ20kKgjjG
LYbKYFuwy+Cb0NWzqwjdQgpEodkfKGUkTG0qHZmmyhC/dhAj24LEcnHbAXcBrlwurw1ukLkc9ru9
+vVlPmAteqhsAyRc9hzMfCGJyEbqmgTSfMnfDkdtDvDArWJJaxRnkkqZoco3SgIVDsVekX3ahkVm
yL+t9Z6M4D2cgqC8ZzT5r5NFdXy5GTc2X1kAhpKPU5vCsb0wwA4NrmVVv3D1Ifh/7erBqj2HXt9Z
E6/AwSYW3Hp5t1BKhSIs7xY3qo9oT/JG3+3O45R8DXTTldg0BZsm3d1IgRrecvq1QusDE5QFr9RP
x0yI7uqy2spSaIF6SLY7RwxwfxXUNltUIlzCNf8Hkihq7wqDdUVFW3PjV6EJCesUDTtZJ2n9BO04
uMR2Arxa60mFgd3v/yvtM3JmE4C1KiQc3UbhSS0i1xXdKgVwARlgJ2izAgFGR7d3mxY5wl+6pQI1
oDQMVs/oXhwCxaOzXbIcrw1qRFvLWBri5E5ObnBqMqrdPd+nGuLyb2+cKmsV9X/iIJf2lTJOFeuU
jKz5C4pTVweHT97rEymMC3C8N+VHUcp880FCNcN2LGmLxAH9pbrYaQHwouQItdrPTBT4qpMyjDLU
iJFno1D5y8oEqhTpS1yl7UtWkerSNUx7wZDV+AkJNQhggld9J8Zc2rG2NSAYqdgtfgpziOfwWYnm
cq5XL2SHuEJ6wP1ib+4lJwAgx6x0sZjStSkpB2YDBwCjSOoL3XMM/hMDaXfBzWY89T1drEnKNiFe
MsqX2tzsG5vUPUmuEJ0VgKjtqwm8OyRNnx0fcxepXPEnmr/IRF7E5SyDmsVhbD0TfD/UEgQQyy9S
FwBXQgvMW0BkbK+LdNNqCiw0BfhLRJj50Rbec/l7iLlxh3lzzxqcvDjRAFpqOsj/re68VV5RehiP
opp2N76DfJcFE4C5B1CUDMpa4rEB01F8TEUWoS4GjV/dX7WBvJy4lZXidBQYv64+VRt1zrfX2twR
GQaPdfpYOuNnEeOL9f+dEtfVYAjpBYzs+cMuWGEnK68vOgQUAF23cBY+AWDqIUS8JgdF6IgArtBV
f040kAb3ZqTmov5QzoXf5OyoZPIrLQn7wY/LKyrIcDyxcsV5RMf+vIDSppmYqcr9AdRm6phvSH/b
ppbPVlTxY9SYUdzlvQMpHSwkqmXhRdR1vZY745u2OCSKtIbh8YAljebOfwZ1TfLBeVBkRjlJ1mn7
N/mJ4BgnDxztigzBH3pfrjbArUXremvdDKeHjuaVGY9Hk7EWevLPbp94kieTwcnAe9830FrbSvkf
pE3JLhApujKyv1arRuEhpr1e2qgXKlVByCJrW8ylruxObIeuM1pHFo09XrfBE30Y0RVwK8EgFj9Y
uhoy7Y8KrEv0IkhKrK66gJgyQLgz3MXUcWAqQlaDWf3LMagQC4Exv8httyd4s21c8h+CUC361j3Q
HWe6rJavJLNc9EZf4gNwQ5Bqkb4qV1mZ0lVjfN/9/OzDh6SjIXzRZQ7XdwzvpXrxqSANz04HAzA5
d1XIoWyZXSajAO3KjW+jbd4/rfhsYp4s2MhznvgoWL0AkSIVh8BJRwhGhDRR9KfowOvemNjFM6eL
I19kvuMMtZNMiuPS3b4riN6OgqIqn/v5dm14UPDL+5jlnfe8kRcMHSI/95XzQeIGc3ymSy9iHAzW
vdwyC7rmT1Cvf4H8/x/tdnleOM+PLoj6jOwOZRAPbnXekO4Q89qILRgRwZK+UAfi/wNsny4vWhAs
XbZvscTI7Psq0vMSrzAPWQozm6/JltSgpGKukgDexEayYlxWCjV8kDZ/AqNbH1F+WpVUUQWQ7Cbo
51qruE1TzjULXnwefgyhykyv/KsFa2k08FsH5pLE136CrZT8bnp90rXiIaVcjihAlkxMhfLWAs3W
pTBnpPmbOoVnfRQg//nXseYCn1NG4ug9GYCkQr97F5sxFsse7Gqm/zUBJ98qzYJ/SSUFCwJYPmp0
kbez34AqFxhTdgN7GYo3HeIHLaCsceIOwr9UmL5cbZUrX28L1B8Eq38RcDN96YIOPxKhCaWvyE2i
NAaYm3+zuZTu83FZd5kD1UBzUolau1ftwd/vcjHlc82LSb8ndFa7gE10EVSO2206ieLEymf5T0kj
LPPwkO/sLuIIKVs1WYM6Tz3QCiWDzPM2epn6etiTPP9Z72RJYs3LgSwdl1zx4Z1jbejOri8Ma1u+
eak7iJycahZRrWXu0QMWYJCggn2i1cZ8R5gjW8XxZ4bKO+yWoJEOKNKlIs2E5FhkPLT8vec3CVQT
PAEWGAdsQxeEGWEpqMm+lBlrVyXkLIUgz8IsLyqr9jYWM5VaMqICRUxFrlnEiAqs153C3BhcVIao
Z44gRq1BzkGGngINnENSOra6wWCEisXVDthMIqB9dTKfndTiWUoeOOtomMCdA6jAooZxUzaZDHy5
hvEdCY94+tFgA7ee+vTM/8AROAD/glx7xL+VL4+cp0pY/DsrfLgggMfeIRfwHbWUedXpDcV3xqH6
MCb90QN4uEgcEoYgtudFJ8JOa8Q0CK9LXHhvbbssFW/kjbF9l/0vGvnzxjkYpme1JZOyqeGdiKcT
44xPgxHGfeNeJ/iVEwSRyjQTMSzFWU9lHY80TWnFLsvC3ALjbNaVFCKvV+xwFC41ZwRYBr5b3zPR
rmvUzKNUoGQaHYLnBAYhPOEqKa/ALpGhtTGLnAV5FdUhCjKpujmT8dzIpSCZJJHw30S8CQwNh04P
KyFRfe6tiOczWzs9UJyao1bR8vBruJWs7chQz93I3Cjz4KawbMB5VAHAcAfzkTIpJY9r9hzjLAYf
dLqsFPM3wznVCkRDQNZAT9BI9rbZhz0Yb/+zWflQlkTdhLsVXj/iAT6vc4LnmLRb733LlsT6GjLA
jNz9J1q02RPAbMZW2iOASBnD3N/FNUSyW95upc3d8eDEf+59wG29QTdUBsgA8mx/afMjqXoO+kf4
99h8O2eAbx61eCCG6mYwoHRs0a3wtiv/gVvRc1xccgWr4iiqNF9W5zTIROgv4mZGg7+zL7tCHmv+
ZTCl3TMqYQ6BVqJ1MeVpWP7qGjEKJrB5HjjPXMmxiv0JqP3tvp5bFdMtkG1I89qzDG3fWfjgZ3gR
hTERtpzMDmacDI98J4CXG+G3PBKVZ11CRk9OPPX2T7twnFNAm86kdSy59uP+8l/678GjxY3BTpBY
jb+L9xgXx4orznTNeZuoA/HzPNykSa65NGBtDaNeF+FMyDNWqQ0EiNPOsR2beE5aHE8DXpZV/B1n
5svs4oEgUfiWVwpbnetH9/m2rdsxHkmvCdOX2jTtw/zC/eHYBQrLB95ZYd3pRrCu+jlUfw1Z1YEr
hvl+Wy9f35+SXz464Tb3SZAukQ+MrvX9yUyLWMHCeRfodypXkZaWbEt4Yq10AAwrcs7NwUPf8Fsg
T38XcWiSm5c+zpi//5shOjpf3qzZxxNM+Q2t/+WbCi8BgWU9IdeTw1FhFTGtcbzbndBjppisdMHE
9brnWaNfo+2Fi9E3VUR2NKbuQMtsK5Em/R/HX1Mxb7umbLwyjFtiUBoPUEa3QOVgOPeJqWJTVpT5
pwnROBfMns+OkknJiAmwANHwoykTdSSM/Rg4g+dtYOwp6WnEsGu3liffMQDV802G7Tv4Q8IDZBOf
19QYlrW3Ee+jrEyLKGA+wvMa5me+zP30F9FGjSb6IhxisvxSxZSxm8rpbP6mRIck7CdnNLQvaC7c
hTx2H9MVh7MBDcq1ISAbF9mw1nu70GKkuIn0CeBy7DPlqd/xKtjjGoS5kIIxJvc9PbijM3Pk33sm
kHmoommQx2Rn/KOdQ7k8irn7GCtd0vDQuJcPlfqsrfnftzLHbb8gDmJy6ymdMsjZ+d2bG+JxpTQe
Tsxdjlu0jrE+rkuJiBtw8rrFAYW86iMAqRvVAzBzWpywewe2MiPbUv8hFHcprVcue98TI/6k5TYr
WSSNzYyFVINPpUU1Rhx/v/gH/bPhNkioh9LyfOayvWQv+n30UXWI2/xxnakWw4JTVcc35kr66uWy
kNVLhlXa1LKNT5m5R0MFmsl4kRDbpZbyhkzdpxwn+EssbQ8V2KT/5MuzmWSfdH+9q6qzAMmm5SPO
0bZ7FjvA9NQSpBkncIPMYFSC6nd7dI0MBxEnPSDWJu4DYiQxYe3pdRdRhRB/OMOnb0UqLFcyfD/i
11P1xQtFsWF57cGFnomQZQMDpc+q2UF5qwNv77RqDtGaDA3sHx1UqZEm6R6MI66Grd8JRxhNJqky
PJxWX0OvZsWx5NuZB+lf1DNboxChHvy/1ejO98qe1LkQi0P2Op/KYKh5qpV70XNYKXn8YhLqc82W
lyThoILAmx/eAG6m+MBHR5HeOGOE0eDOB2o1Tk2FvNNyrrKO1MUXfxMuSMNmbeciAhKz7YrjSJ+E
tdAT6TjlZJFfppRSAH36R71nGtG2wxrjx666RJL1shZcypoM1VqEXv9fywBm2FolH8pAsyfPEZH3
ap5wXqvOnSIp1aczEUYfbWZwoXE0Oi1xyViK6Qot3bhFwK7jemlzjUHFAABmC41yUfaLhI7UA5Qt
1suiVuAFrr4QTisIugvZ+4ixTdqrgAVbrSjzj6Kl4QOB9FXI3ggOpNx3UFEfL7HF7wIjOSCinxyM
Um55LXxGPT1vh1F94VLwsog7w4hrOzJcsTW1OAbkIAu78TVSTBsv2E33JtHKGD29gLPiZL2WaPOz
FfRZg/yNa4mW2ra0fEHE/eo8DR82VvhnbcwesGCwFsHgdIhYmpEi0AlU80MylF/qQEI/g8kkOOrq
QrMmB/OgpbdP0GhqwzzqjksbHdtlyT74U5H8u3kgSM/QN3EFetajkLqr35eym4YV7lMGLmZwdqHa
EOZwfgFOn/caLM+OsJENGrInzQY7xE8ULqQD0CsE67iPcM90kQRWBmVE+RefHKHuEIPJ4jXL/aqj
lFRcG5ix8URvgbpxtQeO4aM1x42aWnqojbeF0K1Cwnhk1iAVQmj6Bnp0SX2corTDcKjizrGkQDdw
Mq37S0SwllWgdUvZAvQVzthKKTgecs8G9N/pgpRigIyAO3oFQNIy5upeWESPs1cQI6RVfLY2Jqt4
yZrScwmGB2ZwuwxLcJTNIjZ7x2ErjK5SkyHtOxNT2bPdI4/VL09MLgMAiLzTukZor+F9R3uxRzuA
PO/HEPRQ3nJAFFBPa5rfh05nay0U8yh2z65VQNxutMKv+74UroVfOyEuQWJbVCa5/LVs7U0fN/Ua
hFoYUGpKWxlYfZVYSze55ZMh2Ks+mvQ+Lh5tBiGUk2Bs2JUD3Na9yMiKpDUoXbGfw49syBy08lqI
fnp/6ZIgXCsxKa2Zm5+GRNvO8qyANXBnlYnwqSjKIUYFs6155FplfYqDQTSJWFW6rxIjrstc/RTF
FFh1e2HfcWU4eIdc4Q4hnaLQSkgWaSIcBXpp8ksIMpKwrcO5asaPLGO7+nAuRSVDj8gV7CqNq+WB
YzXG1EaePmV/uAJCaFOCkqaF0v4FhCSpNk9PBF6ivO2U5z9LIxCuyS6+z7AswQP/aXGRmDJKpO2M
/d4nRW1ptOnZtVBP8RDgGl4CA93CiMNN7YjZJfNFTowCTaE6r+MF/ETdzy16+HzoZujIL1zZVxpu
UkqIBhTq7/chgZR0ImIWQO37iX4RJ0kqJemDAQgoJ21/EbCccK+fBO8v3oUYv65EPCtAWLr7j/iL
SJPIsgeJR5KTJ8G0xGY7ZJjwf9LzloM78RGeAil78UmopGNlCjL+m676xIPPpqOXiPpjOu8+1Xni
n6n8CvCKKKWQNbZhjcvGodpa8XRl+e3wFSuI4k9GcQ4WJMOEBjVbB+GKWO/kfpyAaQcajB2oEDai
7j2/w5PmRL2Gw7OjsR4JmJLG/L3tHeqX5avZybcF96tnARbjbP2WsMUHsZST5UY2uq/FpgpAC2Nq
BQNGoGdU3weD5Cu7KcdmyCObjA2OaKgnyZhrySTDDp3pr6En2+ACrit7kTzXI02RXMQAn34qdqVO
BESFAv2uPz4OT9cQY6ym//oirYLluGeWlE9du489/Ho72Ji+ZF+Ey4OyannxQpzOwtR1+Qc70IzG
oJIyA9aBUelJeJq89L8iAYa/Sy0AYB/Jbk1ARSYQj4BnDJbLBSFDuOAAPUl826f8bHfNtpwzducA
RKyY7tqyVhvxbrzveOcF8ER6PGtY3tp1KeqguvTDfA6nUnFmQkHo573sM1Bjv+azz3xqCqBGMDvb
V+0uStyie5YBsyaPGSVn8QL69yE2IkFrNmenZ3vyAmNserhvUbulF46CzuN/76ZCGkNo+yAvn0RL
F8gvWt3pNbdrSUTcqxONLy1AZfOsMHWHCJBUf3j+tu07B0nNYYtAYI2fbPoIiqRkXCBaTtD1sT3m
0Tin4inaObN6BOEr/1ULuIQDN1rTNg7lkZ1XfOFwn79yeSMcEZrOHCvMoGy3jbNrwHLAZdu60D1v
Yy3rb8D8YJ7/qZryaze1zURgzeezK083pWTX2qGw9m4QjjwkV/+pU4KUl5fzAwrjCv6YPVNLd86x
7l51KGI5vPskOX61V0fozDt2YtwvbMHYvhyLTh3Bvz4ujcerVuonDmzkr4+CmZnWFM1gT0v2Z1iZ
KadxemcMWxoRAJBKmqpZjlq1LxtPkdoS7HWDkpU8fO7xmrQ7PUkhNLSjPI4o7vRFB3QDms33lDnn
yf45WIPfe0UKnu6Hpdeusoau8R7JFTssi5maG/31X4pyvemKKsc1LiLljzfdAwJklAtkiEsfoX9w
AgQZr0iRI6FD70oM0Efjm+nkcJArgNT2AGG1ak61Yw4wy40DCFo2obT0Jmv6i/69sja4KBPlJmC2
29jjNEGQ+OBvZ0+4z+TlLhFeOo3jYrBUerSjm+C1bmpT63UaVOJAZ779bKRtIH06Yet7sejuc+yh
aSxXxX9x/fYVPju2eevqdHJEG61gOftH6pS4N18ZgCwcHcJCnacLBmqCqmES8PujGcUwoP8sIQtW
HGw4eKVBnLfWPiLgkqs12cZlOoxtN5N4hRHcARwPuXO9d9cM4mbjQhV0UHFVeYtesOL0NFoB/T9m
xb+OXmJ6y0TzHGpjF7on1Bwdi1uVkqUJtDLd1XKaoKsmAyQptUHF19BWM6wx8N+aT6NzwQ8ohoWQ
5Myuk1Ev75onW7hEqLpK9lDVlJ0ZES1EqE2DbvQzBOq/3foK+h4NVARAF9EPY2SxsEnua4mdsc/2
dVnwFftPVv4yibtVWdgu3nRps60w4ZZcNLQgO1gxWL1VfNsXCZCqOHOHFt1seiY7ItwQR6K0zQx1
odongYnLTgfnHEuWrdQU3iCxc118iYLt2xxsVQcJljYdhInT8GNcQZMPTAZIVVnGb5AniLFFG2da
qUGjarh5GfXkZTVVCBw+fDtBPnuTc5E6UQresETSrl+2XPYvT+jkb3ceVgfo87MrM5XXmjB+juI7
rayGZTcY/1ahFOTYAOk3csLLlAPBbl7qy4h30mrZ8l+kwC0gnS6dB4s25KRI/035Q07TFUSzQXV9
jMo9LxOI9KV4v8qlw35au5PKX2nphyqD+9RbktlijkZ4moECa8d8yyVOsXjpp3hT07nLigfyl/gD
gf9PlyflXCK6VlbrRpQqQe5/4QtaH+793yWzHv6RdXf6TQv+pOZ+lT/Apfw2/WyFoZutDZvhZHbu
ArG4fZm5fvYWUKMiZr74H10Cow015/Cj6p+y3Xc3kL4BNlneNd9S+3brvedaqS9g2rPesE3lVCR7
NlRI5qKyWmnG7VBwseYGS5IAR+W63oF/pefaR4/LFJqpnlw5OVb2myccelGJHCGajZ32cxDoFjy9
SAAjVky4tR/q+i1T6mqr88ROXpQz3I0Jfkn5MDVrqshAYjjXi5W/TgvWPHR68r6h+9Y1Tso28nb2
uhHRaHkypD44K5T0js0IKMuxLdT1XWM4HCZ0Jeo5oFwFhLmIkPg7wLPkJuSr0JdjeuQNSiMXK6Rp
YtSNanBNHLU/9UirGM8FaBuJLAOb1LjqP5BJznWcsBWdz8AdgyiDTBIdQCUtecM2Avg8UtYIZ8kT
Z5cW9ii4fPNbHIyElZ3fyl80/9CWH+vkxez3J200xRYpSUiteEwzLn4fNJjPQhe4gDSwfcYflLj0
ETtCgiHzKiqMOdWerdaZAjVldR4MbJpyxjixqMTguvezsKMvJgXnBHSkJErbhB8vZKMBZGHNYdn9
jMnb6litfb/ageAlKcpkRZx5Tbw8iSQkw79jLsz4dHGiTj/Q7Y/6H8oWc0u5zKJYUeD+HYcHsS+m
eJhOhEwqSzqt60EU0aIKec8Q2X7jqC9ffwMWGxbvvv/3g/bu0LPKDmVNvd2mN3JZMkS6A1ad1wgB
tEpz/Yw2wDNeBMAS3nHjr5Mkp94ERZFmZ3NuQpXjW8Vhsgs2NKcQGUTODT23MdHUmSxKeG85lrtC
u1K4FuKxNFr9VOz5tHKPn7+Ej/xQ6vIFqvtzYB0dm7r9q0uwivRjwyH7/gM1QJI1isSkXRfjt3h9
oGdSPI2ku3DGvoItZAUxIJPqXgp3WnBXlH1r/3hK9rIy8U23IABy8zgceCNbR+VPvBmnUYOq+Mp2
jiDhlXH5qFdFdUt2Yo8P2zWN6Lhn6DKjUnvaUmMOzaPSrvpR/Ez2jMVIAWnUXq7DTR+hZ7VMpELZ
0/O63fxAAC4PhYdSf4zLTB+a9DEdvVbv+1jMVLywNZTaKydPBF67ADVl9f2Aza6jMxTf/p4cid+j
quq0hthR9J/VA0iLQQC/+/MjCL8EJjvuCn9eCJLK+HS7rvha8vuYp8j/HDyohXpSRxtLL/ywyILr
/fjFNqtr2thglg8QYQb+sLmFoyMK8qUtnXgeOc5levSGeyLEsdCBOp28zoZC9bvxJjj1sI+Lrb6I
gnnd/Yw8B5FjqkGQsJpmV5NtCw72QapUnwzZME+iLmWLnU9oj2SknRTGH4MkwIvcmdTn59yf1moH
d6e+/wBkDc/ghwurf1QuOadQWzib715U6+MrGrc09W8IZKaRZhmT7cDZKt8alcN/2Y9EBTEVkYyK
4h+UvvkaxfN/AXxEB6nlgrE04tFDI5H6NLeXotE3QTJrOeyrIjiNn1pj2AVcqz85anUTd5rXUR55
4MVafdS8YaK0B6JGS++Qm9qblKCceF5Z7vgVhBbVC7QcD9DCi7MtcuK7tBrsenYPkCJHirQh8y4V
WWKSWsj1jegHX6J6NKTAAeC1y7HkZW/xrzJ0HNaVwCd33ZwznM1iFHqp8mOZyUOdHxayQIe787pk
AsPz7kfvekzDI9/AyBROjqLxR6dfFobybRSvBdPTsj/eDRYwXcz0jo8K5wWS54zPWuQtukj0CaZL
kszMVoDYmHWzPyzD3F/l/VWakeCPFBAIAEOV+XqWdta9mqOkaStWN7hMj6BOJsWuV3JRmPEWG+rq
svvrMF8XXJFGcRoRh1NkBJaeCrFIcW9qOKmbvZHXmcurQNevMVgNUF1A2PcTMu9MU6oxm2IDegAK
taMGnHk27/o2mxASHs73Ga/xM9Ahlaojit+Gn+/FDF3AsniPallv6Z2gXKvR23BkHRsRipaF+bsu
VfSQKbycmDhIjwd5X9GCHAnN/mN/lvcbysyGhk4bCdz1RAtPwPjnpTXGWTJ4VCaYhlD0SIrN0h9S
y0zWUvEauwk9LCSCCBKi6aNjBxoRGq/HZINutPuy6qB29n4sWehsr9hzTTefEx12QS9iMOliiYLr
H9iKMMHnmepFIPCeefJdwPOlOki1aGwVjJEJ/H0jNL7/bUk4kzkLK4rHkSlk13Zm8/1jEaVWd5Ix
uvKz8X1Bj4dkxdKdqA5rnmQkqp2D1dDJzRNf2mFkYLqohSHCmB3SnyDbA9GNTB88APumfNZhRF93
1p6+owhhlMb1oz0aviuM80cIBlh5AyvHDog9VLU7vQm4uxVubwMEKbn6UlQJQy/tMfxZ4Y8ImLP1
/VvZ8GLxE1nfis3ZNjIPi1MnfPJDOZKkkBDVrsiORHEvMmJAKDGNFhHmv1iwa/RxBlqtHdoHxlrt
a5v1FWL70+t4cvYC+duD3ro/l/MF5xQKoUMP6hvpilgnVorq7esDqPMFBg1Y7Wa2BFSpGQPiRhps
cyXUl1oTpcf+zz0KMgolZcA3AqCE8umlzo0pYRwN6L2uj+JpTU/R7nH7xFLqsa7XLpwvInHMxU5s
Q8yJzN0C7kWbvMtvTJwm9YgTGu2TdTpHPhemf/kck8VuFcFG4TG5snWGKSdTYQq9AHb//fnkdNXY
FQulZDdm4whTBVKtJcEM1ccaZlsxJmo9DrZ69O0RCZxCtEG9CgkJKX6A9C+7yTTvJJ6QFijDgtAs
TEuWX2zxnVrvy4y/bVEJiatmMrlQB8C+FoiFHYmCJNMQTQhZeTGfnbPbIt61FIQZPT/M3yaTcTkn
Ri0zoSTJ0oVJ0aVUs3YhslCAOBlfaGtS6Qr5ifLriJXwofoA3BqUCEqjPvPbowVlYmgGyr4c4LNO
MHt5FmcAZljn72zv1xfOCOu/eidNnsJWUHPew/XwF7Zycao3t9OVhPvIu2b56SRS9JmyhRkHf4CF
YKyhf1MRoex3D8Up8/kJP5igC/Y8expxn2titUTyvFPA8vHxVn26tEbZYYM7e1Ds9U35o/zoyMen
6pPGLZdgikJKjALd7b+SW1WT+OuQfuEpqrjsiVf27cZn/1JATfHF8/Pv07WfVYYctCG4S/sl8+EE
F0wvkMEmifgkF5yFZG9EMHFrkQaT1+/FUycGZwL4SvcuN5KafDfb7qOjEVkl8wq0VGZ/zouJpZG0
JPH0AAEya1kah9oPuc8lnTGgjAh6rD2HUrFpfpVfrLiSjBEvzMbCYqUm5UzVg4iwnY8Xe8Q23vt2
HyxmPRqQMHl8G8HdIJz6JmWYskmBpXHhsPAJeTZqa+j1urBt1siTj45HBzH1I2VJtIpG8G5cJ+d0
o/zObGdhPvofVeP/UP4XpLhKkFAuWgIbqLH+BK7VQPYeO3eZjXgagkj/CYHM+4KtAKoj+fL5jFaM
QjicTNxQ9pJbbMIopLNPVLsiuPbc57P8KHm7OoCe5mWwGvHIV6jsyl47snA25n4cuAKWwJpxEsp5
bfhNyeeEczWnOT8dHGBlWGfcAkgBdnH6l6xTxHFJaLnml6s4ITUCCUKvzQmBCGfw8JOKjpie2VJv
LkWdYtH/MHLHO/qB/L5OImvhv9Ere9PjL45PEwdEynwGQeoYTAEEMWjYXAEsS7mMBSkFXuuQh9RQ
7gfu6KHTpNE6K8TBUIVJWjL4ZLA+hFloD5f4OoSk1R2IUOkrVAaMJQ1ejoqrPZcu5NLapRt9qFxW
kbjG1jGjMiZI/67Ckl8AulbwMkOlXZ/A5p3xFoKg7sLoTGue190waeaewch8587cU2k29pY7Zz3l
6yJeciNAbmk3f1BKWpLYF9C4duZp7kzELV8hC51SjkbK67q6c3vr9NYlgLFKJ97snNrn9aTwXlZL
zusrHwc3MmaDFhTrbm0e+5jjbxRkKwiyi2YjkthGQUS1p/AwjkQsuHc3bCMIMU4RMqEmVvWPaqFG
iWw2H+WBXNCqwIPjDmYNA0rkYRo4NLOeShKudCI8LTJRj+NuR1Wc+5p1J5aUgkz8hprHFJphJpwJ
7wc14WdiWW33J6+kFfui83cPjqxZGSiwCxeRX8dCMaIoX+WN1B8vpXLGZWDo/CeoKELe+WSS+o5r
cwoxDHESnOBkS0viLaLRics87yzmOrobQAOvHw80v6KcyEyZxEcZ+17sIGkNlMXcR7m7tTWV/kse
6XIbPIbu3PHHZTDuXO+Nu1crDHGzALsJGbmmINSo9BdydXPDw6/HavqQCE13R7k/K+USkosbhfoA
Pjbivvi658yL+CA2ahGIp6gm8+gqeCjId3k8XFkwF0GctmC5HaN8gLhmR1xygG0Rr4Ab2yjZKAvv
b1wBcnaPXMLtV2B4JxAOrlBMbJmNrhaW7VrN3tnojnv3xfYtEv2KAMwdlt89w4QGDMauAOt2Xjdd
ylVg0hPOwYoEXBiW/A3sqCKWcH2S6vQMY2+AZoN4o2miT9FTBVIviITx5QXvgAbkM9OCLai7PB9Q
GU18+ViemAnV0sETtqOy/gXxt/5aIaL6d5IsoLFvsYlA8skPvjgXHi73lBey90CLkbrykbNsAFM+
KHXdCj7iGwvXcIecJitBcjP7czjjvUIRQqLfT13H0UPGlityvnqFo9SUvf0xQDxim8yIHv7CxMGF
owBg8P3nemDzYvtxxmj+6rheU20hGgxY75xteWyCaS6DNqLn4kHLDyStzu6DCBsu4LV4ZtpBa1YB
D/He6VKSQJLAUQIQmP/efvEaVsMevNARCcy1Dusc3KvLJmYVIlDUDH40rY9Ra8oIPkMqmY73V9Pl
xHM9eGHtXVMR5vwAeYirWi4e4xfgeFl+eq/HY5/YI10lf1n6m+DHC1gyVG7Vf6ZhU5OKBqLV6RUv
sb01fUIyL/Vqqkd0pkXwOxl5HA3D6KvjLwk6h0Cb+2jY3Jw3q8vgg9i1Nszj9R9bp2tdyRtGl2u+
0PRd31SYFH2f4hJaOibWf9Nr1i20zG9eeu/EyNqRSOi4lY0YNHzwyAL4awcBvnstgvW/Zbz9lCbt
tafwqpvxvTrXil65V5sn6nA5iwihl6OG9Y6jET5aWrEN02bJJA9M+bJdpAPlyae7WLjGbPPBLQoS
IcUL1MtbR4p0Za/yB3TgPLnfbeM+Bg1+hP39CF5Gir2TXAgVvNDU0pmJKheHhJ0EUDiwAB71IdV1
tyV9G+Wzfe3Oa1RO6vjqW7gtMcH3pJR8l4mFBk4jNnydaOEKhUnXlY2By3mUNvReaDQIhWbOG6Lf
0+cU4MRR8Q9FXmv3t6lkrmlz7dYuJ81OO67TOG+czjh+huQDGAUnTOCC2Cg8kPzya/0EdfgSjMWU
J13+AH+Yx37OnLhEr20usLk/hYIGy/kIYevKfZovG/N527Z8o3o1uoj+pMF47UCUmy09eOnn7n+J
IAHRZT+n57C1wrnJBf5h8xSoULtLCWlLfro6HfCR4oPJN9OLt39OkWeFbH3CFYJhgv+zNBgm2B8s
o2fFGi3goyFKFG+A7Ngw0ZTzWZtNN+Msg5q67yvmxfD5V6Xl3WFTlsDJEwTiNs4f5jVrtwm+DNrd
zSpAp+AHP90YQU5oguNrhCtvTYLdJuQHnAJkoZGfRugUO5RcniVD/AgL/RlMx0c5dD9TqErWEykH
nIrK6szwClHvuNWy6vvjGRugbv15N48t3CEXn+TRifnJPK4HJp7aDJQFdsCnFyI3J3KXbjxn4LoH
5pGTBcDxUp6rVkEESnGvWXvI/RwnvzJB3SVbiCvzfrQPaZ4JODQ+SVgJEES/RpSw5gSYyYZ3uLDQ
sb6FlueVSNEYoswDFsyrOrHogSM8dpwKK4G+60lYM8NtMG5Y8Y4lTC/UsqbpSrBYI7wjwnWGebI/
vqBjWwPs0FMwJfEsDI5KzNUAGf8KcGesOZpE7ZzdlUfky0UUuWZCCNf2sGXO6AcJ//hhnBwfWE5r
s4tb0jTf8mmQP+A2kr5wffoRDIsf90RQw08+XG8PAHYR93AZ9O9O0jdEwio0hNRY/GzLBicWYeK4
JE5RkVzAf3af88jhv6hgHgqSJ1o+c4Qxt7OPhqDst5IWgdtRoD8/fGTlmFywxQd9WWKJtApzNc0A
IZRoKkZBff0MThz+/KVHrA+fxN/92xAO8VJXvZ/R3zN+bAIq7e1BveVVRZu0MmZ4hSTepyPyrGe3
GIym8Gf/ePznTI958blP3bovaffKDfQbBfwPaPc14sKu5ozCwXW6qRC5PDGHVqyianMvllMObg3o
x4JkV7/v8SU+4HCMb2bg+GsQ8+Hj0OGRbkCtBnTzzC2BvLoi2iMUGwwup1wo2/qRqSGPwasm1ZVH
HZgowcv0cv6Eh72Yb6cUCV349TWefirJ1qGNtx3VZfOZ2krKejpmXI7xlpSi+bS8cquD5VVTsHvg
HPHtNzQiHqiOeyGLs47g5QwyNyDTuIj9AC1gT69lK6Aov+uc1IWj8c1O+vl6RyCEdO50yXqWPxp3
mAj0Jr1PSGGcu20yzmnS3aGjON2SEDjZL+YQhYT/SpDsqBJfXa6ie9nmofNMIS/USdkINql4ee9P
UJt6LCNcKB92yZZj/Eh6S5sckSBNbTxb0obVLUQRmnjC2BoGmg5SCZ6PgRS+2NVBX0Lxj37Hak+b
gOmpry3TnKszhdyBPf7SctKPUODM8gFLzcDy9KBCDeZNzesPlwO+Au1PEgapHE/FHxHM9Ak4VWHH
s9IinNVA7KrnVuTb4mQkhw4JouvwvzKV/fDfUWagd/t+mHcMBfVG+XppPGhYvARRb6JTmMfWs9dW
eAmXsL2qjY21X4kTe+KggI26VKabxWfSjLrRB5+70D4vPFWp6ZxW31ehacp8u1J2S5iwf/n936mS
HOKfzf1E5AZg6buk2uAYxRdZF6QJqvwIakmvGPMqqSLIIrQRjrKU4gp9paid6wz/vEwKDZlVG3+G
Wkbs+LMEwunX0LhXkW07zgHXi3D4TgyvoOBjaM+nZ9e0fN+jF5XiA7ULqkjyqphsFHXw7pKofp/E
/U5dRpZZvYIEdO7Cpu98sU5JTCmD/xBUb3B7R7ncx5qHtraheqWQX8DT198OG1AUox1pAsn4NgQW
eviYgHE/uhmclB2SKcLoRrdSlWWJ45SerqU/TtL4ao/fumjvCCG5Fw/DiiQKVl8ivQYznjSShHgr
av9rkXpyZCyLE1qFYZUYqtCWAEj4WrMcgnGK/WC7DaU35lXyZBpd4XpzWezxJCbRZDNxgtqTcH+C
xbOGbzzXLi/mPqslu3A4T7CJjWk3rPfmtc7ld6Mw0M2SK963nBKiUQLbT/V4nwg1SFpDIcG78bQx
PI7fB/i3O3KphxThvW/zOWK7x0jUfux1OWJMCFR90NUTMjmOKYwhjqVmKi2HFx5avpPjX2qUIUsS
VEbnAGpxsNutn/yca6Rr0iuS+H0MaBtNgJG76bzgDx0kogZhLOY/lbHLtmsX3JydwnfSTUJiV52O
8ovpFi7gS5Ca8SgufqP8UxodUyJ5CZB6LxaifhzXOIsX0XEYpRiuIylQWqIda/wooaJEswZelQB6
Hm+nvX+GtWX56LKhNd05hUhNmlHcRWbMvdxCJYRqs9KiHSVzkcIkJd5QrJHZT6t0ZdGjRI/LvmdA
oQSmhVQEwTVCYY+lK9DH3DSpUQNC4MQx4T7DfAuA7Ia9vqswpFX8cXl2Jb9FBumVEIXzhE1EIiDp
1gJv2UWNDULvkZymReu4fQinSwM8egPWujzJv6PO5X/n3Y+HDJfXblx3cmULsptjotVgHjIj4xRy
BD64f06iqpV1IBMesNvZYGll8VMpw+17bCig+1EM7L/WCOJy8+wFaKYAQGaNGSJvGIP/X8RVFwjs
GrGimIA6oII5jI+9VSkEpuxcddzUVu2SjZpbo5cSMnKLqoq2Pruk7Sbr3wGmNI/qDOWlHVu1H65y
3PFE6t/Y2w+bg89eS26R5DKujVX7iC3qjgtJOiUjLkgs/cbD0CEpTvRyPP7oEvh8oCPvcfUCkQ+m
vb5maBSOpaP7E5/mz+LdnB/0VLMj4+ap6x6Yy2PkGyEli9dzDd0qNCllDwawUidmkyLOGK3LAaqt
165UR9n/aRcpdthlxbwY5Wb3SlcOgB0evudWUGFTxKXfTLH/d1lOs6ysSrFZPDGQ8JtKs3XhSWJv
cwkDr6xiCrn3C7e4GAVRmuQTHP12FPA7mDI/8n6Rsrm9J08k8iW+BdPPw2lcNabwxWcA9EVbE5AO
2Yz8ivQKHIdNPQfcJvaoUPfZ1baVi8GlTOwuHk5d3EH9QKK6Iwlhv45zdZns2uAapE1SOnl4SnW/
AH5frs3Z0f+/arl1nh1YBW3M8g6o5IOOQexrJPAdpO+//7qvwPbd++V/0sL1jQPMKa93lIaQ6tI3
jl33uIN/vvNFgk+EmvHoQqrtcfx9MXlJH3kPcjUpXQE3VM6GRT5AN4RKR3g+XuAi0z3C9EsWrDeI
HUS5bhWBZepbpXglmTCj6YvOCI2l7FF2EQiw/3ktwavO29jf4Lk07XmSMEMynJm37MScV5bMmIw9
C0H8FdhWWUIy4UiyoEinFp8BoORiZHyimn+n9LU9joQEKr4NoHOU/omEaVV8zKIqHXyqlreKPB02
dAeXxRlleH3b0IO8hlOabxfvYyyiNYgLX6PaWkcX9KY7MU2A7eDcofVp3zM/GN2WTtMIHZJ0rQfR
mPk+Yl0LZtRm6QgaZHdDXKsNu/4qdVL1excuGX2bmAZZZvmsEUgjuUqW+yb/ice91wcEe2w/hBsQ
sxLl4OmuoJ08Tv+5YlvOqAN7KPV1sdGKFGQ5zKqqAnxY7URSRRYUJL8wl+RJYS84p1Xrx6FWUSGs
ifHi/nPfnu2ALGCM5in/0C6HdXEsOC9BZUVHgQ0plArkKvvJKGU25fLPCVQhVmXao2XV8hTxQ52j
g5vD0/z/vJgchy9+IWS1BhpDZJUeWXrSJK9aPUB5g0nNB46cdcUNM0IVcdTqIefqf+4Ke9YvAE2G
n3+DlOHBiEkKnaJYFrk0u7dDuOoUyLB+kGD965Kh38g8jqf1utWGKo0B3dDtemrkt4UxOGtiNgjJ
LeIJ/+Fkht0j0vj8HPEdc2oZL0DKGSEsZu0jWgAjhtRJhBihCQubecRAKQg1G/ycGMQXJ7n1j6h/
mLeILDLEZ21SdvxFNoz2Uhucnr2c+J7VptQOfOGT3B5fkAq9Zh86nXsbhxMzAg/aMptFCDUaDQ2B
n8Dne7n/rhdeLqsfuTAQVjDH2o4az2r9a5/xnuR+YSxAhL6f2i7fcgAB8Gl9zgb+rjPE1c49Bnuu
TgqOelu4ng7I+94LfPoNUX23sW9BQp2O1tHCnbwUZgKv/Kd9Mrq2+6eXl8z9neEBMY+encpQ+RJ/
nnwlrpBydiH2SuzndUmSol7p1hGpBsdr5pT8Vf4F5tho8ctbymtYOOUtuGJ86Wj2CRCEhC/EMAsl
DqjMCvOQV/iJGgrXXmKqlp43/kkafMAW0Poey6IhQD7HnQ9LFji4C+YAi+hCWq6SS2Jk+sVSb7hP
Np4mJ6/M7xZF1pGCPfbFSTAr47qlIAoOykum2r9RyF+4QsAQDezWg4cn9xImH1vf2BH86SoiIC47
054gxagdq+iz5JiPpZBRioOekV+NzBTvRM1HljD5S/+0o54oU8jICWW9fDf8nOCnpWUpGFXn95Y+
cJm8BxbexBfQs0cehyUHMWjhHBTYQ1uMi+OW6Qn/CfUCVg9v+k6uBnpy/1SYctiag7OOT1cN1yqV
Ql82Gy5nP0oKWhabuwitswNZbEkBw+4FF1sEQAKA7hXh9o/xvy7Rig+zDADZgkymq+p9FIvk3g5b
twe8pQb4nmTR56U+lKe3y39Xs0djXK3taLdJqQcy9N/vWByHDGdDZB70Owex7eMEycznF4BQR4c6
BSspsKqu8F4rKn48iakW7yLimEcutgv1g7TpAOfv+KudhaspGwpYB1H/d0MSg5A9tDa8XOK63HOG
rOoe9Nr7TAtaA+6kVd8ssh9kNQrcXOqM3bSMGTxcb8GAWqOgZosl6mgb5Bg7MWU4Qh18ehQ9y/bC
mz50K4F06T3bWTOmyoLpH6NfJaPM9mJ30kO82Yyl9OPlHP93lGg6NNClbCNKS+OvFf9o3DB/BSpS
oMILuUKXfayYKFjgido9aZDMdODL0MBZ1Wp5xQ6Ytto9UfeK8UC11QhqIc7pUGcMJhlqLsvD4GE3
FNb9+GKBH5uMpuY5grj77zTFP+KuTOrRsWoD3o26Jkf/gAQAPYje5nYWwJiwCoLakUqB+5d8UDBI
2VxbXOgMCsQ+wIaVO4mU32arEcSPNqr0R262kidMuGkBo8c03yBnDe3imYBHCPEgrKlZWn62PcnY
zb9rA4KxQhR+m9Jq/Jj3tGPUufgd2R15ahF+QHC6cf6VU3Bp0oMmqAiqVb+rRrvAW7PaHWmUrOpr
NGoMskNB3CkhRo2vH7vno/99uz31V2zlcRYcHTumY/tHU/DfPO3ONPZJnwMnB6kRaSQeoR6KcOys
IAYN6ghlSRscJz9trSdfoPNCRHQHpwArr4Ht4TXRH8u6PnCoG4/R9z2uF0MKYanogk97fOYJE1ui
0mt2meqjI16HVx47q+rH5OzFzwRGMBFwD5BSvyKdyAWVIyiDdJmjSr0g3vxNjLQOICAY6Cnn/3T/
u5YnrDNF66cLXlIA6fZv/nvTxyjEyUi05C7nhcON2D0+/fmNT1BuMS6Zt/WWDfNenb0RdYNj+LLV
uAHjODYElam4dO1AVDOTOZiNHCW6RmpvljLNPi+e/tFiKHCDQ1Au/p+U2Xy9Yaxxfps+gW9Ii6Pr
cWD1czUaaxtMRrAe3KDriT0bG3Jq9gqChh1IEMRS2nPuq/BPAC5H3xqqYcDdnZr+v2s4zPzRbtYu
uGWYm0A3vFZpHDwS/Hpappv0lxwbq1f0KwVYHwi1Wu8d6BkzYZ/2hyznFPLkVJO+zYwDcEFxCnQA
1yM2KK7DK4yAL7okcRbNlBkHKR4szK13URz87daO8l3A6HZBD1i7yQDFlF7ES8uQLdcVEXkzJeJ8
d6NWZYSpsFTj3H7TUJoeog/9V9UmMNFXGk2ShfzwDS4tc6V1dylIka9pqY128J1R3nUV5i6/s864
+iirK7tSLWJGlTnhK28f8EHQrgHh5gxfDm/h5udukX+vwb3uZQjHjhEtvw8i/T1LSv8IISXoejXc
v3hZwbzqNhtJhrweyufQIpnXOZw0R3ACNXHDlkhdJn+2ZBjf28UdeS/nSWwi8+9BVZJGrc9u0yN2
HYuiSgTBlxx13m0ewJBnWCtq386vCNxdMRBdpQtEYRYe2gv3ZW5DBnmyXyZ7lZyor5jBk25K4gKb
y1dY7TOfpH9NMnEHh9y80ECb97WFnPylUSFm9ySOpNNcaI4wR+OCOTlBcxiFXREG+ORIItRA65cj
2KFai8pehBOerjdc9T6ZfatpO4fs2tRmffK9kbdhPSpL0esoY81GmncYt1SP8J9XhwF9Unee2kW8
CIyLFaz0s+MCP277Q9kDH2MCrXlUhG1doA4jx7J2l50AY8HPBCDRhSUN44k32IUY76CYfcunicgk
OFarh8mQ0VTJVeH0k12MpC9jxLlXGStB2kmnLS93Sqg928PdXgnV8V/2z3Hzv7SGhXtKlKednNYn
Dw9opOsTDrOSvmhqDnEggUwpayYaqk/Zv6g3/lw5FQ30cdScWx+74lF7uOFUOTwyyAK7UAe6yIK6
AqsAvHMqxw/iaAZtgFSGQlD2Fz+GGql2dGdv3ZkzYoekV/6wTd8OKJsifBdzGRgkXONYp76m14Ps
Q9U+SBcehO4wnAebtReUyM0+QJSBRDuDXMB6ax4nPcpHoVcxuvCoGZhpYdKggENlAxb1hI4lQJGT
Ugn1Wg6jV+VeoDHPTlHENuEcazsXrH3z1wZ5oM4sZz9XGRof1Ch1E1/F6TDRW8uVe+3A/CIhEAAj
YhEI5bX1XwHpDq+0MAjAUP6D4SZ/qBMv4RDk2X94uEOEFowrWgeGDEjHZTUBbxQ2R7DKC93y/th1
urCpTq0IvFYWODxfZphSE6sroUg7/YG2KQQg5FffVW1blRo2+Ft4r6p/1gIzKQz/5xY4apZl3Qd5
IDaacMfvuK8eGXGsqjuEAIUkClhyTCTbQ21vwa4YWrvMe7wqjODJfptoLne5q9Rd0LuH4v0OboYI
BCGZHRDXOy6X85LEJG4ltZHYWbtdkU2hiqct99AVSaYMBGwZsfPjJkfYJy/Iej2w6aCjedHIMO3Q
yJddYLbKAMhzxuaoWiGNi13Am5jIMP25soBpcHOjoAkXSGpsadXKVr6GXRX8EM8k4FZ3rt85N8Ia
j/rEplFy0t5FqvBtirIHrNJTPkejgLTJkBoouHEB0PUUTXm/PrshlE4FerPTfEnMZMP3EjGgZLEd
UDRzurCPBW40pTvckaNeLZQ4xsyUp7IH/5ZWjQZxiYUa6mLCgHjNY9pZt8+bK72n28x1ulv8UZld
KoOf+J7w9taLfJJ5Gcy3n27B8Dhmi9OxTzrkYOlGLf4cENqAdG5zhMxBHpAFqOZo8gnEjXOWkth+
XFsZXRlmKAKQEljSfHk5iJOlH9hBWb7XHYmry8zZDYKuN8WFBsmeqRCaVdFyF4+tPrkuQ2p3m0M3
+QUr1UqtRKQglTJZxMLqcAqdL1S+wh5tG+DBfjQnN75MrlbRuU1H822u6pkRiY+1N4NAUF5bSswF
rBGprkZVfZG5Y92lr6oWjU3a/08E/zIOfANJ7RdTXOMH9uAQZNTqbiJI0hCj9Z4ySmnYyFAal9mw
RHG28aTbCzYAbfNtcY4Zpg0Fi3aCqsqtIX4rDkVrdliZRrSLydutQ0VTRSNvUXb4gbKjF/tuTlCY
PT/k4t80A54kEe+IaS3dL+G5z+T7lxhbDd2NcyJT3t9UebHgb1W9dU9jGp5lSDtTVAL4JshvK796
O07zHp4mtXEQz8AVD0XGb6rbDqQ1fDDKNK1gg69wIc6V98X+0g4i4aBxNJm1unfjNAYQgEbS8Jym
n2nA+eZitXoTicTiTevptueDvCoAwcfoks5dvb0zJ+rk66M314pDFpjBdijGNN0h1gKD5g8VhHUb
DZA5usQMZOBuwsRF1XNGoXWHXjM62fqmjwLTafThSom9koYOxdauBqwPlGkFbBT2WZxu592BsDfU
TYIob7yntu3xGdZShoaRiHs9rUMTdHLgyVyGhgoUp1jyu3BykPG7WWpduJvxfNNe9Mg7sgNgl+oB
oO0NS84PFQVo7AD6rufRrlDLLtFUoRHiFbGF2NWChwbidPLiySD7OhfRZOlGUphw5+TqI3449F6Y
XPRRQgMjToQygZ0SHsZ3ugbHNzjcwLV5vuL/3AEe90LFRLJkDQpK+vX+SY72TMYSoIz+VUwWKzR+
p8v2s3xstcHnof9fUQYXKp3PY6PuBrcg5NEV9G5dSID4GeoqQtCqkzpMV0ewW+jR1vnWraWtEt/2
cZ5brrdTE++98ZnepQJRXNDpj6iI/U8iJUk5GNjH+ZQV2s3eXmdiUS+hxl9hTQu5DtWSjvhduQ+y
DB7GuSBlLdjz/aZPLpLj0v3VQ644jlMwW3rn6o9Xz40peenHfqfFHo+PqrJ4rN8Swihe3RPRivO9
c/yYX2f9Zqb3cmZ4CZ0YTYRxkmAjmMfwX0kZKBc0xBXvKv7vpbP5vwqciDZFMV9k3uVS7ZP7WuE9
vrwLag/PtrA9xR5YiXykWuolf6N+DY+nsaxD6M2dlbupE6mRcFUkUuyCrEKZ8pqI6Z/EKsQrZl/7
/mnDo2Gcx2LzFRFfMCE5Qjd6W90usQ7mOhmb2VoAn8EOoHNzyuskXtFSiioLigbKwj/uXo9Eb3Fa
7Lu03AUbQZKJBw5UvR2+VJ8owayR1BqMu3yOBKM36NYLYRCnXU16h/DUPlrfexZaS+WxpdO7gaGo
pN3AjiqCoPlUFqzEHGgUcVQHriU6sc0Hdc6yR1iJnQVZkKfPXR9NDdhv1GNnXa8kCa8VwMgSwR+y
r5vEh+n/0/0Kxj9DbOaHeNKe4tmOTP1w1jHL8SLlPdCeUNmouvHtGTumbbFj6GR4vx3gklE0a0u/
vJ9Nw7GHjdo6x3AdBHiWR4qCqLo/z02QR2jM3KCaCAkdFqe4CKQH2x/v8mMzG/KUVUMYfF8H1QR8
j5gyU5SCtK9UXurPSnOwguPwoCpstEpidw41JvjWSVofGmPDffm5I0QNigrleziQz71k/jBDDCzx
6pNoCpfSl6aLlDfKVHdgPb2sXiete/bo3oWOnXC/TGtLhfdipEC0Plv/fW/+J23j99Hqo6U2YEhe
JREh4TANC28ckiT8aQELMniE2R5uBacs428sSoQWOjQ1sLC4KdJvu29ijJ5nvgIBeBTJdfi2Yjc4
GpLkuWUQ9NcIZ41rW8HBdJxp8kRNq7rp0MRTU/m1eqCEXWA/9m/NoM4sKiqm7OJEJAOq7Nv955qx
kkTEhwa43xJ3BtxJ2FuwbcK74jVkhb8otBxqGUJmTU3qywuXIeUMEzemHYiSXIoy5n2pYyQ41ph0
WdvLmOSSSanzeOifWu+aiqj1FCsqStMVl4mrJDunclUncLZXnCpOcVZkAHotYE59RvPiZ08KFm7Y
caTK01jg1vcjRewDiHY2nTv0zyAqK3PmMHKUafeyLuslu143g8doOI59MNTvoxhiBTing+t6Bza/
gQr6sgqL12EgDuq0ioM1cy+BIt+sRL3IwjXGa1xKPc0ihb27zsLlfSVPczvO+0EvrJWsQBhAllpn
L+hcZFDv3J7UyFhSBc92XtVYIMRC3UyjwXyz41UmyEWHZ5rWOQz+WcgskcZUMJZMMPnvgVzXSN31
3N7Gr6FDcidQj26XRGNhwXewQ3zCgt7pTOiRCby7vt3/SbZYIYZ9DUPPckumhLbGmpiKinXq1W2l
XNF2G9hDfN1S5eeEvPlgLZFlbHzFBjlp1JstaV5g+S/Df1aXRA/1E1WHHiZSKTNyyKNWPFZbpVSt
v6+ja/EUAOJgTe4uXTGBXI1CFmA7EedidyVtFZdZrNOhdshyKvuHyLF8c74bWf2D3s++REAaQHpT
rZKsV6QjMdP/UJs5+/OTNTbJ71mywlGANwUu9Ig/ElW0ArUGInTZFxszaCX5uqXaxlEU3xLQnPoc
aF4QMcIs/KzGtPM49NnvBaI+oLeijmWVM7qjMd893XtbP7oQ4TKMu6CrFAQxdh+ioTqUrolx8M+G
QHrHWevuc4m0TX/SXn21O0DR8yB9hyYzTDeXPZtuwAcg55Cy8c0t7PJCEVBbI3JCGQiK79uXvPb8
9vD8WAs5xNYO5a6rC6FZJrV55wIc9x3bYqQED8G87fgLzvoWum+vvJNKAmNbhSy3A99YJTHd2Q/4
s8k5mP2nysO84fosqn0sn5q0pf+qJ4M3q30CPF7IQ7PmqaVCfEgaDEWKGfDNb5pvGvLuRJm7Xmo7
17Yf5zZfP2bwECRLpiAnb3HtA1bV4LPcdyomBcy0KZdRXZd8sAsB7h3UbldBs3GTpVGeFzom99QR
3tgIKa3fj+kujlaGxEQuANknHuYbffmMwgFdk7GgqIZRn7aWrXOX6gUQXiGR5kdxytlM3W5tvTrM
ZWfagyuRrVuXVaiGd7xKaG6JnjrSzZdDoenw0mEUQ4PBUJx4eJKGnDg8SLZxk5rJ0Ve4fdPU0g5s
svkJYAGJjK62Cbit1y8JyjDohlBo0aPqywr6lvzQALghDZbSKaMUq5x1YJUVd3sq7vUn/aEMeF04
sWvzNauEh3HjaZ5NBGoNsysSHTLjk0Yx5V3EelB4p7LdfMtX2wHlwJTwP6nCCNRdZQRmg+ZlNELW
fMFo3pENqTcnpEdMVli4RU5E2wjZktTjBgTGYlaLN04WGfT9jQCLG7HoDdlq9ORxIDb5svRPThED
/aPEBX9Oq10vD6Z+MSZbBTgs373aK/ThB9/Duoxi6KThN3lTgvRRpz+2eY+t28TYMHKMh+AeIzfz
1Myyt7/pzPXjISiFj2yfuNprqPBVs5XBNDeg11Regy5UzzN5VO1+Z7GBzU7E87GcG4yMq1uXS5iD
giQUHYWbnLXtocO59UMDf2CCIw7sroDKTKSzg2D4U1ZeV1gGkMkTiZ6Uyi78qHf4odfRVdixKUBb
silZESOemnReuq0wpL9f3twzi8ob7Dk6syv9x3KtLijd7DDADLXLE0MMpnEzN62OQKEAI2OhRa6E
UnqeTKMn3F94jqdHnicDxRqs4riwClMTErg0N1w7JZ8D9VjELavu/TmFl9ouJXNiGw3JrlmnD+hB
zgGCkGXQS5NpDZlw2Ah/tFUK6BOIAj5xs2djAfIXhURGrY6pgMhHGfVvwoVvZ78pf0nF05tMMRTn
i+u1KVS7bHBYKBH5v4dZVffc1eDEiBFYQMgTQM1izEzRlmuGijAf0EwRr3Xnz6dzCjRuC0QqXLxF
DJ9f4ibMc5oohOkWGanzM5m+eGD0+ZiNC4oK504Tf43nzPiXuvA0HdTV9POD3ttxMRTKEAsfchVN
ZyXFqGKi0OQRhUAMPnvsA/wO2g+9eU0yR7gTF5Xv5NpIaNjJ80UX7rK8H4o8qsqGQNdP4IIKU6bI
lwn5rmvOI4QGzewMFdsUX/bkt3KfQSonA0NB/G7ahAjGBr1na30BM12x6F1AetFNtj/99IsnNH+D
JKzgyjCuY5/E7DDtutfCeQaF8PCEhCNgqe8qWvF1LgKtcQbrevVEwr+6h8HbuFhhqKwQ1FNLyl7K
NACMUFfOrKnlg/Aoc5pWira5iq9Y1vldyNybp8kvCWSiICyLc/blBK9kIxd0zlIqX9w8mJtLopwa
ROboK5L1o86pLdWjBHSnsHyNeUb24yKUiRIZ+YajvzMtH2C/SPwXt+50Eccq4DiEnPFmVnPVn7M1
t4r0h83XuM6fMNiIyaXPjuWuooQN7BBIi/nsLYDdL0ENws/O09nipZgc7GJmPUIWrPJnvZpzyqur
K240lHdIslmkDb/38WMMc/ZAaNpwyH+LYw1TcCd0TWvIvUGvR2ZH6DkVuQN2x8DNlTWj7FDF5VbE
QaxJhW/Zzwh0FdpUc20dLWcO6IUjjmk7OXgqKZgIo6D7+1hricbQkBM0iJ1eVvByWjF7VTgnHwDL
bEUtdkMwdMETxnnfWYZd2gjfzKDUFdI0uaxKvN+0VZ6C+oTYmBjV3S5Zxst1QV3P2Id76a/3Oth+
gaBpzJUt0tCuzQ9DgLqOakG5Az67CjPsqmX5PKU5JXWftqJ4072fpWDuJlop0mtCQx/sB22NCghD
gewXt2IdP+YzZ7fFgNlhCXchpW+nXJbmvehvCTj7oAdQNPLlE1aTg2vDUIoIQvTStzZN4Z4ZHj2v
r+oDLXLfEb1hgFNvk5lr2MXsPjJ1hNFw17mfksNugSnDbmNf+beXd/Q3PnP1YoYPnWviqSmxuhhF
e2+jJWgsH7TGjUcF4yawQqxIxRtKmcKftKCZf0pkSDKiRuUKWqcHdhUihbGQN9HGZohlIGEedWrx
FUEvK+qeOchn3wmkM46xs7GIt7FvnWfVzTZVeynEX6JaPoD7jcDC+QKr8SYJ+HD5flu6BnNqgak7
ZU/7mVg7KmZ2jGw+J+YP9kFxoNAlAAv5ZmcPzcQirwugLcNsFi9xW7Yab/YJ6KAWKS3U9atggfkC
PNEREuukrE5aJbvAgauiRtmTS9pzNPhXA8DMutjssc2FKx5Xdvv7qSuDwO7w8YrunQVt/bGtmtsL
dFjoS4MjYFIgRIUP8h14WWsd9IFv02xxd6LbsEPSACOEXqjX63BPiLQLC2WCx8F5Eh/0euBbHlrZ
rIvpmDMQ05nYWqC5e/sDxAHpxLzjoh9jBTUUC4J5eake11ecUosR568ZUOp9WZkNKY7rcDVOldgE
890LGmdun5fkUqitDzOI0394ABvgwZxaGlCsOzRymL0NpXggsSxMTq4VjCJOH2amsdOO062P6+lQ
+tTHnZqb37H+IIafw5MogAjBy9ZnD006rB9m+fd7lVfh27elN5pSywElijqv9UHz6W+x+p9Jf2eH
03fwApmO7YQwPRuJHk94ZAGwblmc4HPzAWaPlER3recwQseh68w7gpLnT1QHeNI57M5rAyca2J6p
zJ2ic0wTK2x7zZ3JrWPxl0rJ3MnyzVUegYKrgF9dlAdrjAoNrZK8QNAwRF+HPXL7ZA/T7br4RTHv
FYwU/xVpae//w7PkI5Z0nFdES47WPvyZ647JJkdSxgA1rJyQakA7XdE2KAsTykUuWnualxyuS0Yd
XzfhjeJfOyeUycpIui/IdX2ewMQ/bfTnQa5JAC+L/1JB/Ae05950DnR8FszFG7xHmirVaiXAd6LH
ruDLVjTtgq2KEjW40lsSgGHClMErCFGuDVcfdLjPABi1WRS35sgBXbd8cjCqbBib2gysnu7LZL3Q
9dfOv5d5GXpea0xZFZMoF52Nyi+nTJbk7VkZOirVW88d1T17zVcfEB5dUtkDAKk2MUos90R2ItdZ
sSAOmYp6Uu28ylH3vnYN/9K7iXxpLuJgsMJIlR+5DuLFyT7XvwE3F9SlIwfLOtIH0SIdcr6OF26a
/US7f+9c/q5D9yDiWPtSsFvgymw98S1SyUP1A1UAiI6MpIQ0XJAf8gqNpI/yAn78TkJS/2CiLUqb
8cs5sZy0IukVKGLC+wTBE1Dfvt2RT/uZcRX+P+0DAKh/A8fnMp3uzipSTGz7WHcIslBjZWock6Wb
zEy5IDEAIMyOIYmS42yJZHV4vLORGGLY66dak+ETP+saYNbLyccAr99ZrOT5cpuiiWqQY+hZwG2W
CbxFQdB8kCAl/zh16HwmJiajih+Nn9U2DnOgPYJPVQjS9U5GiyYQrX8H2yvbcbNtY1pNOLqI8qu9
D/cQA7kW6Iu+4r07+5AJBMBFrjCz6KZ7XxlKP9HUr1fMnJED6E2ci5Z4e5SM70XkhpyZfH4ALM8o
k2NDZViYx9s2lrpIEvtXV/YvLaPJn42thMa96oTAMFeytiri4RkJBDHwIHy5bMAVtPWMjr4uh4j+
mHZIE8sC/CAKvPQltjrzbhQza62FIG2FsjNMmNTWKYIeEX6R5abhEDic6S3HQ99HdqJDXyS9GRRf
7UqqVtbiD0LbEZ8V7jlHn6+UfnYHLuFIcGo/GVrxy4Z3bHjE9Fq0Hi+fjrJzR65pf0YSEAFO+Vz+
AgrursGPUUgMouHAsxNdimE8jePKssH3bIiSr1OXVDiPcon2668g0BXzFRliLzztEhIhyfa7DC2B
seOQ+fa+B+uXQlmTmKCZdPJG+n5LwuTZ+Jw9WsYGwviJTHkGi4JSqyPIx7+BmtQIc3EIAqdfjQo/
lU5nAqadPQIY7IHfgiWGn7UzV8DHbB36+fcXTNQqPsW/QYGzUbuPF0dvPkgPQ7/tHftSxVWxWqNg
Vjk7QYE2UqRUAqkSgk7Y79fCQw+dDi0WxBT9oQ+0VFzCrjNEc6QJg9NKXgk2x2/u/yxnRQahfBBf
Og1FJ2C2YqKE51RkrmhbqMF/n9qMqdF0b9MQbsKX8uFYqfCzSrLzXMmuszRRjfiSvn674Xjgp0m3
eGv70520P62+TQ66cHyyVCr1Lvnw6Tba+9MENkfMuOUW2U+VYZXwwvyarhkAhcm+W52VXpH1S36h
JhNWELCl7wmUrUk4mT+PzV7NesNJRgnZxoDYekn3k2KVMfCwSggAkCz+5hvkpN4OfOqggZNiVqjo
2rhjvEuArwUbTNjMer+xTZCV9Yz7W5qVvBFYYqmfdvTdzQVOFaG5pfQzy1mYHnUj3NcHZLCDKctm
ETpxr6iVIePRXT2ZIfhorZ6cJL2a43oshfnGx4QxGBKTkzglnFwOvhnyZAR+uvqGYS3gx0s2v9Cj
CnlBefZ00Baqk3WdJVgnmbgyg0213acTZnaUA5DPKDCpSS/mW5T6xNQ4WDvokMIQwsHast4HavNN
79Zz2kaTXWUSKflDSX2ghUHywls1ubmVFwzpKB0EkNPUewsqP7U2W1SDtVSbdFr9Rqny+hxdheAb
OFqYpbI+Ts9QUflf/767V5rkTVIYdYoCq1te3x8DuvvePmLmURRIFXDy/NF6QERCkITm/WBOnJ4A
qjdt259lI/1QEvhCPZJLXbxYYPvj+zmBwoBX1Ss7Zg6cbghzfMGQeWSjlM0hFYgb7u8eGhdv4r6x
u+UVMfagtOHRA5GAyXZ1xa+lG21JnDpDa6dQu+GfYn0cqlgtGtUbdKy/VrqSUXZoH91clCzaFTX8
PGgL5k8OC3/08t+hL0UwrZzu7VintZRWjhgZmc2sW5HT2EAzJU4D9/ylV4Ocpyn8ihdZsJp8I5W1
iraxsu2OeSEDPw6JyMIIrVsKwJG5D1j8tZ7OZHZ8Irxa9o5lB0F1kf6+0T49dezylWMQjQ6fkF+E
4i0PPAWTW82GMcjNOn1dTzWcQY4eRERHEtx444uFpoQDpmXNtYo6+JGpHjbnbQCONGCV+53DuxKO
gi4xjkJDRBws/gVdNeZEZ6a5TOVc30FVLV6RTjhEmgh+WW/m7gI5WQHLK4Eiwd6tsz5ihWj0cJAh
ga8WeZ8jOvchBTrDXK+bVpCHxqCWCnNQ/3zsQzfnB9/Pnagp9V4Ppba1a3SnyrSa5QDcjtHb7xHh
Fj5edgQHOjDxi4Z/LFPtVl0HI8EXK0TV1IRqPp0LBlV3tQE/BllAD5NLlzfAtlXz+5W75bkz7Giq
w/9voRbMFfeysQNclUOS1O6u6hYaAMwWn5J7ofdVi8BVTvMAlAIUEUkWnS0/GOlQy0ze+iBez0D8
gKOlMgGf+g474r+4KoLoJqn0Ok69KPkwHEkC5tXoEyIWB1gxINvFM7ydljkn7IXr+408ts0u13A3
EUp4R7pXPFBFIIwEo4djxMQqRShXuNLjrhaTV9U8hLvJKaIpc/j+++FKsFay8OLWFBxtNxHhK3YO
nUxj41pTnuugv4IOgeXt5zplXILOaKX6GKw6onYnckdAvZ+jkUM7YJuLhd/+XKI2ddk1J3cEWMoe
Io/Pj32SFg8K3r3f/Ai8a+OHd1UwDHdSUWYU1Mlcjf1dz4fZeI315gW0bHJnuyU3aPR0QCMM3oEe
IeHn0Y5YW+/zF8PLI8s317lIuk0DLqtZPqp9khQuKEVKq2g9kxxBX0xadufzpaeh4JgtZZDIlQss
yqkn/YJywpvtCD9hPS1VvZySsL9JKJ6k+AvkKgLz9Lm6wmeAT0sBCwtO1CmyuFT0C+Mc5jBMrzXn
6G3trGnWrMcZ9oo13402WYNtPzW4EGZCrPU6Tn2mXkZVaKUSTaHOvYFb//EEuePTC+bV5bHP7R57
5J4TfGc6RGdO/gYOAzK2ByA0o8Umtbfs0NDel8vcTSr9hgDQvPoeoieTHzulWRkSRMl56OegHfHZ
hMioeStOWDwVx19EjYyDLfKQGCY0qka8SX46RYlOuGIeL/cAVyhLPNoGDeCv6PoU/yeoFm1YwKGQ
YVckkdIcpC2Ia4IgilH9PAuTHp/oGjbNAVHTR7fnwIbtGl11y5W5rhNMe/Ea1kcgQ7oFCMq9K144
3d/mDcfggoKtuCC00nbUpXA3N0R91gYOqc/k7SDxRnxVk623xQlhsz52CWWzjU6gRhdaQjR+XIAu
ARbIrj+pykOHCLJGinSM0YTYZwsRNcOVBttw/sydw4Nv9k3iAA05QcNv2p0wPxa1KaGWq0kra3L+
U66e/bjET9Um7HrrPRMoNU++jbgqTTCJlu2OVD2nZ2C3LMFYdfiF3DOIye+qIh3LCHqwO3gstR+K
HXQ86dpyokr74DTd5W3KwKaGf821voPnaKzVYPP6QFsebG1kdl28ke3ZMNRvP6jBhLAJXX/CuMsz
V0+hwa/Ed9IUNeifeCAWqowzB2607XVOGsgRKYzcaF+iRtAHK5pHJJaQ/+0+vaX5VJ254swZbLUl
gyZYbtWROvXZLfaNKp7q/ESPPNIDjGMtMaZPgn/Lrh78u7ZIBE75TY+VKVWUxSHDPnHEu+mawmQ9
p8gp2cAsQ8nUE/IHoh+/ADo6QbadGVwBMHM6C5PCa5wqEQNLrDcpUo4WXWyDV5+kbiQ8yqEjyKtJ
jduIRqGnINdtcGCIic0IiNrqIqwKI2Ks9Go7cgKETyIjeBFknuXibCjwxflOwdR2VFMq1B7Rrrbb
8iqgZLBKpqKJrp0XhSJMw8HRhdXVoe8oIkgnFongB0dyQNoOfESx/yiBSbYHkvH8NL9yBpshra1k
aF+QFPOPLhfmqY9V/L/AeluPmqEflnbRsfq3c5k2zGHpD5NElp8ywytwBom1f8uZlH23sjVbrZnR
VbKHse8MVUvPsP1qNB2ai0J0nxQkREuk3C0MeVyfWahdj5JpmufGgVpC1Rsv52y1RioeziON0j7K
TBXVmhw2daC7EqxE4gdri248mBkvT6qy5T2auTzErLIh4x8YGrgD0rxUUiQTjfge8pp5EtTl6OKZ
n5YuUQ4bjDhN9Nb7jYSnwnkMkYCay2jRpuQNQaH9LoifHXcVobTLaBcJtINyJ1RPzJo6Dx7heQ7c
ee+sWbemOEUvOh0lwqXQI/d9I+GluAefdY4tdb7ELt+4OJQ4DgHTC1PRqCc4ERet8AXHQSRiT3kr
RZAkOb6pIYXH2yevzKRy9OPPdLMPr3lCiVSxdcP8hJUYYoZX5j4QNlhnyVFiUOG8Q5sMKyrpz3oN
XcF13W2ITIROwI/Q4F6ENiEAObqLot3vnpCEMX+l/+rtAnlZyoHj4c7oIQuIYp+K6t+VxM+sb4d5
p1sEFFHCAjLiRmPA3MyngHxo3CGjBPPodZi1Z/Q6kfJZ/x4MpgwtrxQnYnrjkhk5a4E568Q4uZrQ
PlIWTH1NCkA64Ek0RYf+7VBp8P0XO0826p8ErHruGCUg4+/RfGYmtntzxNhEFVVt5FENPQJ+MUuT
us4bgML4bbc2w5n30JAa07APUWVaqXa/dGILWo/99CuustJYTfmqY6o0WQb912cCNwN++fiqaDoP
q9DY8IBp0vBr+06jHzt4WB4o50tX1y2H0xoOkSPTbFoWdoHh3Ilvgy/vO8VJnJgF66eiY9mOiZqz
PFajrj+LkqvJORRsHDjh3cUdGCKp3JZtZv/nlehxTp8LlahsqxBOxCpdzvX45d3vKP7buEZCkAfB
RPIu5H4ntVZ94aku2W+ZxQfrGhxuz9WC6KWqvsbifvYfsRiSS6GGRnz1KXceJBhNhWe+zI7hA6xP
H9qS45MmIrZr1PyAaePzBfJN9jjzXR0tC7NAMY3sWqNx8nLdj8c6t9rj/4vRhfp/0n2GHN/HsJHz
ut7A7qQ2cv/M9gCDX8x2KhJbyHMVYzLetL2M29IbUEoAxl0mexnMQaxIgr6Uc1aTZa0xfF+l7Muc
r8gFJR6QiWqFcEdF5jgE4fEHNcs/j1tWy47ahsOgGxF4RYPg+JUUfv3G/SvZwE7nfM8mNEhGfbBX
5k4Ej46HE5+LAzYz7EmErXqK0F5+GPgD2rC+kE6GHdW5V8WHBfmQMI4wQGhoTofowYH9AL2JRRF7
jBDLiYdN1lXH5Gpt6QYL3C2lzJlf52j2btEjNAGt3KWsOwXGvFa1d5YfsnUjivonv1qEEBV6BV/o
yiolfNndDFnztYsCdmd2jMS0KYseUxoTDLYABA96N1bH6qaN/E0T1ezIrQGSzaWHypB6vCd1Nbk6
n+NR6H4t3BguXigItHQfUOy0YT8l73GTfO7T1/OeHWdG7TfOad9TxOduv4VPwyNpkLwoxyfROuSu
cm8yThDBCSw+TkxMVbzgTpavjj4ArluvB4KxWx+6EENImva7R35i5pEn+qabINneZDIDaHbaJWZ8
IawXTjolly1gFN18EatAc/YuLauNc/wGNBOrrajNC0IRsx+FFptii+cAGOIGmjl8tBqPUJa0+QkM
EG6/jsa+LTYSxmJXH81b5zhiwOc871DugEY/pCFBkIEsaCDdkKOD/iCY9rAs6O7j3znTQvgzb0S2
SkZWsLepq4HsDbSne4SMC3GsmS8xJDLJCPT/AjhfeNkNbak93xgZr9+AM0Lhtnl7b1yfeX0d5c4u
BCWWfpojmS5Gc55DqI+MVuoJGmio+TjGkrrkQvjQ215u5pDitFR7DCXG7Pqp7EY2jnyACxnKb6Vz
I51JEEc6FBpK5xtQMh3YLgcapl1nuo+Kf4ar3oYe8z5RUu+CSbSVceOKqDxyo+tinc2o3W7gywXC
xzLpnmipOdnzk78QqAdxvkhFkIdk0ZCfMJkXiDutrtloQ7QQpvQnAS/JNQav3Nk1yG6C3Hf2p2Jp
p2DfIdlIicivFUVg0dKvPPfFVxw12yTvCxINazwXqD1xLU7PCv4P3IVJXXQk0hShUqui/JwIaD3R
AIqqcXCWaQTMk+5wuC5ocG1VYisEJ7zjoilgQqRPcsJrCcSzeYF+ui0O/TH36AliRj+cVUsNxPbf
DBbZO+HlWeIurze5X81p1keiEhi6RWzSfI8CryWHmBaK0N1RTgDuY7HYi7sXqCayf5tGem2vnqcc
S+v8k2gemLsLZKfjOQPQjI1fHD24ifRJGjo6jUpx/XWytrEGASmFRa358nvpeF+pmRWXZUk6mvhj
AUaXp/vGLmFN4OkyN1CJDTGl5BwUagubcwKYGbXIYQjAYHw9QFA5mn8xvs5mIn1VlG+lXt4/5QPb
y2d5oR6UhwLIHBLeAW7dDd4PCpkG9mDXPs2rVqNCxg9hmwELW0vD9hygiJgriKNjwTE32hATu/af
j3BlH1on1W8aKfEPitApLy9UyOTJqS3guTKcnnTQa3aULd4QayCefrDPWwFPIicBa3qcdpf9BaT7
6HpzoSVw6GSFv3GzL3XQbWOp99LpfGgiDgKeceRFPDOm4S2aU8uHwpMMd9OEVMDcQTs1FebIRhFq
KmM5d/WUViG/FgTSC7BojMBgJPm1OtyAXSTgG2xpJSFYdR+ZVIyngD40RZmqFNZolwVnSRjnB9wM
Cf34U+/aqy0UB+pFzWQ3x5wcaR5gmNzu1ZAqXIE2orCI76MPBZC+N8tJkDnqdntvJe0LmDXAWzJb
2vPigLk4q5m/WcAyNlRTlTRvJx7lM6VOrHAKZ/kYJL14UpH+EGRFLCH3UULTd32/oLf7BdqBupvw
qVZensvgrmmCGZVlevOx8ywaOjRdR7/zo49ST/aLEXPMy1/AogzwC+pjygbUirDH2XXforD47el9
eJ8GLWmUwlHXLalmhwqzz1HVDNp9yienQ5dbrehI3hQZwLQr3Ew/tM1GIEDu0iYJJVxqsAVHDvCr
dNn0iRSwROFz+4PQdrTdKpQ+Upv9FUAPXHNSaI9uSjFTOYtWxCLsIGIgbrUIYqy6G0J6X+7flDBo
/rhdiE7uhlF6iV0AauSPmPMsJL45ZAaJJdDmvWrABz/OhmJl01/A5j4RZ8qwJ1lecOdC2IsQSd0O
BCG3evfU71E3u8rP0enKS53UpHoYtvgFOAOJHP9lnNXiS/eDsOgLa6nUxxkJ9cMLHQHtNIg08D09
q7WnosZh6ePN3LfuH+dC2xA2/tQdBM4XCG11M26pjTdgsDVT2AygirWwaP0RHHijjN0MxBiDw68M
enbUgjeenOxfZxQM0/I17eqXZOZqPo910B9WLBIZ8QGR6UAkDiuskMmEa4piwRXJ/+i4i8xlPCTB
wM4q2IkH6B7RHsAFz44XgMlAmIToA74n4AMtSdwPJ2KkCQNp4t8nwg27Wg66gS9ts+IPOQfTk8QJ
ThRAPnmK4losTjoijxoIvnUKCJrkEOMUwt93jiC+hWAbodZ5N437tQ7cgAjaLV2zpFPGEze4K93R
6zfaZfAF0IfdhGK0WEGMDHk38UWMUWCYaav+MVWt9iw/MmPCDE6fGhvsZ/9egl5mlDa9f9L7oicY
WbkzezJhvUqrp5CJ4gZslliTFE1s+ctWa4FH2mJlG7k4H2iz+nRoXMl80uDAydO59OHlW4Y64zuP
IwtseiJeM0lxceHFqEDxO+ON3X1INmDreiwH+x05IdmrfLih7OHa8gmXHIOC0Y2UZttAVAKuuCPc
na1Q07m81MwZAhmLx6+En9wUezrTAKk2zQ2UDmVLqAkTYt8QOM/906An3v5gk2Or9ji3apVKs5JJ
BlruNQlz/wRLCye9Fi293MFwDSB1F+1aLbOQs3OeSn63ifdf6gl1hiCqigNLxW4uhQ/4jkLg50XG
Qsk7SVfi91bVk5Fp2nrfpHJfdoVEjOhqQ0XM+zEV6zH/gC5G5eysuLXn4aTc+p+lO07pUFnT/G2/
dQNxf7YSGsjJszilgQIQW9Hc9Q3KXPWzfgbaJy88IdW8PqosoiXkY3J0uMv/foVaJ1KYlf1tiz4P
DEzCYG0227/fM40wijYueU/JyrquPq2+Al0JNtogWp9u9OXDRnaP+p4WLKvWTY+VQlom0EpzWyUE
fqUUbB8tsBCnRnLpEq7gkspVUhgiHezUhTMO1z4HYINIABm5EvqB57I/Wnjybg4ciFN3JTsyl3yM
HmDH7Lg6tb44UMz1YNez9Wp/NqaTpa+rAiCvgphdJfZ3z7WW3mI+taBgzQUhtgGdNpUIeXxvORnI
AWpv6kcG6M2mkGFAkVsTVQqRFNNg2oyj8xg3lq5Pi91VpY0ujC2NbmgyBHjcq6yOXNRAQiu4zz2F
RfoUgDXKvdnFgqHNbpAp9BLK4wMLBIisv5wf8rCv0bMlzHoCSa3s3a1iZy245MIs3kaw7tU9gzu5
YuqMnVXkpnn/JOyyHRkYQCxT4kIzp0+EECEKeNaE3ge5/tEC0u5uhyNYzgbdUJZ8QJR4eHe/Ff8+
fGWSJvvuxlssBp6FCN5H4xE8r6CHjcfaZhOs1O7O/wcU1yNMTDZJIif7WiC0UtrtCE+5WYDzQnuc
kG01k/m/LiK/R2m3EDgAkFh5gQrzR0E+bCTb+UGUOBhbLPJwQJgswkFZZQSyqt7iPC5OSSXqIqN4
uNKbZjo8wjDFo8E/5a7zZBwsKbnK3e6jtKSGw6HnuNrXAwtTByX21oDUvBxpQqvzVCqfnJAn0PgN
OaLWivtWrgffjamL9KXz+moHSFKEjalJfbRVp+WuOwG8ZUWSBJFJ0ZMZOaOSQCemHdg9UlFLE1Hb
Y39cVycJ+1Mx8PDyZMrRpQCqSwhnEi4NkyVFt7/5X4+hCsStK5IEYOnlo9UUcgY9MuZr4I+SMLUM
f+Pz8YRHgvoVJKn30WELc+D/I73zwDY0L1wNKanh3pV4lx6cEngL0dgrvjR/AoSaOHaNapZLfEiH
Qkfvp9+txD52f7hgVg7id308QIKJ/3j0nRijdB0cfNFhZY8lzdKs611+Vb3qdOvL5d6aizktHEmW
uE4G3qxAh35GcilOa3HOlPiBTLoeGkTbv5QmAfT22CTHwUbZH7FxzIOZYrbCB6EDfHd10AnBij/6
NAmRgtMcVZRdo81d+j7V7q96UTY/+XdE8xjtHZZZ90Bh4E461iOnOs4YV7j+8P4wBXLF+24h+VA0
7HJlRnb+TgXPwNyJIsPx9Mamky8I3u4cpdGdzYRTyHDSVZM9PsVrSkVW3zfv4GicoAhU/5B1wpvX
qe+jHKyPkUUS2nsLfuVpzF21PkkEtyJ/fvcAiATofxMbODnU1rHzS2dPX3EPDa7MnRCHPACQyodY
yU5FSbU1fTW8PVciH2w7WhkP8lLGqgU6mES7qN3A/MBejXhCsTUwbeuT8RC8MIkT8bbOeG9JM4t2
mvY4bBAqoUdgCuT+9sHYCLqsWrUmRcw0Yy1uZ8n+BSUnuptXpg1pUwHnwbRfHfTeueb+3lyM3Zul
H5RTQLnJ0kQhncqPUN4+QkbY6EY2Tv+c6AzkInh7WFjlYpzBz7Fmkls/qNEnLCMgGtpKyLQqySQC
qWIMYCy316h6w11kjTao6l2apiVY1E5OqFnqAVTs6GmcZ8J+bdL+qHufQOblKzG1EuaTggv6E7HS
yHUu0GDbKc0ZUwahiDSuCYqNOimjmQysQsT8Ullr9Ey5s7I3ZQHzxF++mqrse43N/tghxuGmGh3P
ETPaeAFvn0elSeKznZbDvdGgSPsplMYP6hi90x1hK1oYKYsj/BSl+h8QLpjwW/NmZDY70iRlytr2
WVFuVIQ0bZuj1WOh6Xuec2yfxUSgpbUgwSiZ8JVd2RsO5gX4I+N6J6NOnsrtB8u+PA/hGhKFD9rX
0Qjcyifk6lQveklTh3rv5AmQsLwprCDVqLhwHQrwmVdlonLjzwc65l6opodGGkht9/DwWdbfRZyO
mBxhLxTBT4WWM/ezL8lrBf/EYXSMY4k5NIaLGEUzB3IV2L2uXp5f45hf+5+9u1090g9svmlGqP8I
ZmRqworZ61y8s5bT/eTnTKefOjpUszFFvMVwvEGWj66PUQ4x4K20rVmjOozHH4ZAMI+qcDAOSJH1
9mjta/JsojczGSiPC4O6pCOX3CrgwEzFgyfn1bH0vNrTshqIh5wK506nQ83fjf8h2HDlFqHC6XO/
YqZVxqQXdZt6JOD9IVSrvN6KRwqF1cKTUYNQ1wndQ82xxgavS48lGC13wqwWJjW4BiWILnL0L1r4
OcTgUfcqAss1evnnfSx4X962rkfFLSozOQX/YdarfIzrVUf+obMCjTaro3sETiV3sYYjvQrZqcba
lw168TCZoKkYgnlksXq5B2fdc7fo/KW9p1k9tSe2ZTg3NKsJHccDekwrYcnAV95TAnKCV77q/EWW
Gi7YJlWWFQBciZ+Ah8cYZCVVSJ7fTM6dkmXRO89pb7HTfNV0obUFrR1Pxy52HGgh8PkfMsawDNdL
TXmJyis1zHP+z03QzE8gorRxmaJJGsK0M9TJhSAT2ojfme26hIhEQ5KeI7XvzUEF8y2XlBEI3M41
ELcvfAJZOVu06K74koaSbnhEMbGrwk9YwUd0OEJ5jOsOIV23RRvB6ii4IxgIAwrrV4CXrBJbqQdR
vh1UjNX3icYa3UVEWEkSPOPCLwNa1gIwz+lVvRUjjT8dM2QMLBex0okYe2lTv0uKSWMTCaBNhyHZ
LciMh0Yui/x/HhgwiyUtYnVsSJWD1K6NzEi5yMBnYoJ4RyvkdpP1sU9nj97Csen0jDO8Nfp3XVTa
x7tVe0SxjlymSAY7C3p+aPYwJE+/a8WFRhJL98zjsvUU/9FLv0O9wkuWYzd/LFMTOHMr52Vj+is3
cPDQI7TgLd+PYas18AT0+2IBa+JAIOfC1F5r/BpKxxcY9bxWEHK5Aa/gm1SIyNYHvVmpWLxtPSNR
r2+qxYQ+CwE7A4Ku5uQVLXWPHcb/lIjWJ1+VZv+gk4EyM82EhBjS2tpkTU99y22OHgzWeaAEDidl
6yIdYCfF7N72DsdLVqpQCMyuuvfYSDNikc/8o7Yuapr6NgHWLrukEw0jhmAUHb72i1h7rgipPtvj
hM4rNK3geo5pof0lbY9s1J4AP3H9CSnomZboDk1TruqRK7oT8wbwlW2R/7lhWN+c+D3k4gSz6ZUi
GE4Rs8JursW2d6ioROQqAKXwK/1v5qUf2z4RqG3ECTUznWyADhvbMRPnDmuJZfJ7nOZZYHLppvLU
PSe4YTsMYIBu1kRJWBaDnb7namRk6M+WzOYjeQaivIbqP6qxbK3X7qnEyG5LPL2e0zGoNDA48j6w
OB4vv7+Lt+vLHubvmlMBmeuQ9CsTdztBi3msK2ZdtskAtxLmwywe9UBdsAuWedM5YncmaH5lBd7+
2HtcQMeow24btx9KGq30B+TF+3sD5IcWM4GE0FXLVz7NNZPDZYfUzA9YP8E5Z/KG7o7DzcqtJyrH
1OZ9mDKyDi2SKvxW6C4FeyUb9UHr+2CzaqMW/8zf1OO+E1W6TdiNbhP40aZtwL9x7fVcoN3hDPAV
MFtBshxN4Ufc1Gsk4hWi5TuVMR/5szouRsqk1QFepUdvfBOLHDNoKn0uwnWcinLaKmP5ooo2EFmT
pQoHuHDARUFOIJ8dKgFNySqDX5OSxlWHyH5bIJeOq9tcmwHZ5YPOqt/wStrHlNAlFIh+96y5YQln
pyiL5VQJurqU+RC/JeV7ngertQUfO41XGmqRq4CumgEBCNlzM4AYptN0K76aW6OoWolElcvGjtMb
NwtNiSm+L3LlkqI3+ILme3cc0E/OQJ8ai7fXWXPoKLEA9avH4hRHb/oMK3Miun8Qi9/8M5OiCaEi
MSrvcYMlo6DicM4oMU7A0H47Ilw6lUfo+kns69J+duzBiA1cijWqsPNnzAa7F2CIn36GOviTOTvS
Tfa0ysH9JybDG6aVUTn7bG3NRNru2pMDib/8JplDgxjA7mteL4iRE2BAaUe/Xg6nYKr/7D3IyofO
2o3Wn5JzKGeDjKt965mseT60e414Pi5hfuOxDWYTMPy4kLwHvud4FS3wwbMAsvisUKRVYpyomVVy
bpfI2vGNPnHcew58FLa8f6+VmOYuu1J+gtoIy7xhT7CVZ+yiUee6iIV1FuyvinHjQIllahy+5eNO
PEBphAaP4NJmV6Ofporv0fHq2FWYoNON653huTwOkcXqhLHuYVBOMvb6H0dishvE8AFxX7gdLWYS
VZRZG/P6rIg4t2eyWigoNxQALjB7wCOejy7VhHOAFLshkuCjKJKWWXGh1xZ1qDzKfufjG4QK8ncA
nWwQsJHOyOHDE057gGq94H/kRNmBFNe0+OojqlbTo9a3kQcG8zUKcmyMFRcJuqQBaEmBlg5a1BQT
kf5yAeSHrZcjvVo7i95A4XOSzYPOBZP/O1yStZ5wVW254uE9azbDRQt8G6qcyUrp+OKSoRoWoFNE
JCpd+2R5BSMMiateqPdzzYyHWk4s3UXdRXgDg50OHNRkdpVG5VjKqrfnC75QjeoJ4YTbirqxUw3C
i+IUMqiOEYbmzqbGTiHhdx5f9ANh5fUqx/Bw9p1UvtV85Gd8+HsLstJ6TUewEFB47GU1yuzUIFK2
Gi/IpHuRww7bToQQezo5laVH6bKC/Bd9zo+TbF6o3dAFtyzKwl05kwngdKwmwGBF0jTUdU8oBY/q
oxkyh4N6jwUduS7suvA8+bR3PgUnGwdVdVdhomnOykMOoN0+BzB4ldDWml7pC0cr7vb4Ui0slpq0
/fNxRaFTKJbV/jrC5Yaudza4WScOdLgxlUF5eDdW6ppK9xe+s0f91qEo9wYswyKPHvhcSxJDN2l6
O2uolwzKpOGXOn7czcSDEqncl4tAb83lY8GRTqMxmWsv/H8KCgkBW67752nGl1V/utQVrfiYuzY9
Wj5jKZp8dm1ewPXlJnUFCUd/NpczpZegFVD+vSRod4EREmJrg07sWTEphhVvfoECBh/5wMLQS79l
i8y8uei4tGBfQqn/vGFZFbAPE70X3jwEHPg6kWit4ZAAhxHXq+Fm14kU9cgpFf0XtsFYlsPpUJa5
M/yRJiXPLUsRwJkA7qRvK0RTmJklUuo2oKSHjB8UGxMtDSy/0pY6mj78pNQlCb99Pz4DQZ3Z2bRE
oLNpo15OnAgObgsOIhsqeaFHYIPGcoKD41HlkQLgUQgD4iF7OhlVu6XEeDAg0fqwRTXK920UnbYR
+4H1nrE02ZM9lj8LFswq36etWYARZ3YhZGZUteCYxIna0loLpXOpnkicgD1BrzMKOe9LdYf3DkQm
aGmDTSZiFEcaysjdHEjEJqXXk8JzGWGjVsEgoPdU/i7uZ92dHJJwOtkNMYPPxM8UxWhAlmqE6cIR
KMqsVJf1Xben/NC6XwmLq8HHO8R9EGEUjbbtbyuiNJkPtQ+hJ0gi0RhmR7MrqC0eh8/y3GhPmtBM
zIDjopy2ZK9sSzZ0chazhtDZvDg08BxWtP48xtOEET7uWUVoXFhXkVWHC/1VEvWl+m8P4CxDw0iT
Ps2LLd54wcRDVNhfEId+4wKoN2T7Wv4DHgilZxpJfhqAdJNtPVFh7hv5h5v8gxGxFDd1q5ZJ3lrp
7FH3it0Ibmcy2Qv67kwMGh2glVhrLmdB49M785cSkXWT1DJvuBmxqlQFBHQkg8pYrbMB5z1XR0LW
KTqJ7KnEaYR2iOdJU8r+V574r64LP9+uV2kg089PxfBKlTKpNjIU3i9ckaDg9Rv1MfD2QKB3xiKh
7+xFvr8NtmOCszouuqbnawme23R6O85mNrt1C9cVlYtPnqgEhW0b2j47ai7Mjn0gsrz5w7H22zWh
EKtO8nOEiwr1a7lWZoLqvzPy4mxd5jum1GBNe4czWhtL7px6j9HehAIWcKHzeWlmUIHNOgr4APBY
HFsYp3KkSCOpEgd/Tq82vb7wF/Biikpj0Nh0QWbvhjIjIINDmHgG1miIg95akBJAyGmNelsl3ol3
/3PXK6h2vrQ5X8gTkr+UUeAc23ZpYk43uZdx5L/J4grGVphH+dkLslCN/CBLswIK7/8X0Zi7t6V7
2nx1hIB4xyVeWpXc9YjfUg1jJNG5XR8yPklBQTUtjWnUWXpemTbvfPud0B+QTYjbxjzHGGUNYwCE
FRcKr4mvFR3OojwuDcR9zjqZfIW+FaJ22jq/0iCAJnlRWBmPOe1PW2jLY44zcWC1c0hoHGI8k5Pq
jUpfBeEECDAnjkTmCh/KdbW8gIf2cxw8kYVWJgRez/FGxpNyw61TF8KJ9nd0zTG1BgOykqlVkvWu
oDBp/eCFgslorQsZDouR7YrJ2U32O3p8LGcCcZfc5yueoPlhjm0UifexGjybmiH9XjgNipa+3C/t
A8L59NLQO+zgichygRqIvjrSw0/lMEovS1J8SmuW9Vd5yPs3vT5PYK6Ma0bsuiDfVcc1N5iBpHrK
68JWgLgXZqfS6RaNYcx97HqxxbrXKnnOJF0i3YmLTUAnB1aLT10hnR6W7BDDG4kUPpBIdN23DfqI
RPCHPycN5zkXidnk/Y2QJ0T+FusX8N50zns0NIZXmWLuZPDdB4wAlYOYwHyszEPQh0TONGWZzj1J
6A4i3bkxJHvlqS5kXhOApwGsrYc/pcjNrTTpwgOb76xVzOX5c++sA5f0BWyuYcy9h7WNxuYneC9A
gGfDCzKgEaqzAnznw9lOo4HTTqMjsjqEGYGkJI/FuIYfAIx4SQvs4S9Xzv7GeNuXxKaLQJToFBUs
a1yY0XkfsEwhOjpAGjwAb2F1rPmyLBtChjhSMFJ/4WuSc31Z38Tn7PsnvfIxHLTnyO1SjPYxvV7y
ZOwUJpIkqDu43Ts6Z9z64kl6updm5p3aXgT5zB0/KNBr3TY7SBIXC2W3Hj4cLfG1IXTTMMERvlYt
KaM62FDYo1rHAPcrWapkhcH7sQXTCi0D6OVIx72v3ejgqzj9GGC/qcHeOuIwtJYEJmrcJxYOmz5W
bA/j8f3nWox/VoVuiGrrRrtuFqc0FyROLPh0IcPxwsXKuiO2nMZmaYIvqWChnZy3C7RJ6vqXp1eR
1HjihFkOgGY1Lwa1IwQB2Wlaxa4IjV6c1D971hlMqbxs5at36fvaSOevLeAFcZn/gb/8Xpdz34hy
KlTNMmXm0UYqznUV2h2C/wnqsVB8Rvlwoa6P7IUpj01dKwvyKsvGuL6bY4TMLIgRtGHfCZz7lqgH
TgOXMEWPoa3MaLsZexr9PScJLHjKMLZhXlWU8ELIFhW7GXk5z7tgm9M+YuqN4enkWpk0+AuuQUiq
pmxqWFX1xh2KkcAa1aXxxkMLh0+v8UWZZ/v4Qr2MX+W6ojAziiRD9SqYJwXVmivorIPP8g3lf3To
GVQSgaiAZoideUNSA7ifzuL2IVtwx6mRgQAoOh0Lj3+VzpSaXQrxusimKEojqtiavT5PEIQuz+Q/
ad4MtI4KPFJGYK3U9rIeHNN771xQadGngt6uhzrePjS97BO7wrK9YXTojs1RB78RpNmLjaA2/ui0
EHg+rCoix2PSS/SuykqJnqFAGSTOXMt18e4gG+eTLwV5JduhbdSxgvWZ1nsh/H+vvDhj3WbyLLgk
elkGyr6Fi37Ht3bmHXiQ+u61Ce6kms5Mx0lnEo+vT6gO0e28J5rJdosss+LssKZN9izALn7+wWwJ
YuCmCzWk/oEju1ZuwVDJDclMAg5NB/Gjs67fh5jTnx06PMirGLk0F49CKNHgyxohzhMOhBKOAllX
taOvtDuEg1T3x3y+oqgZNKVkZTV5XpM+2Tsss/lYVqumi1Uo/nU9U514ub40FOD6rFFJN2Lp409B
+9K8IqpHD0GxvzRuJM1wZKkwyELAT5AXna02/3iWwkkH7tv2dX0PzkmvoKJ8mOMXCyrs78y0Twf3
tJeo5U6uPxuMyUTACg3S5sN4ULgQuO/7uSTD5VWT/j0LFWuMiKgs7XyuqWmbOu9MbQbsihEbhHMJ
+uOGz/eH1Ov5zGHaK8NOl463800yLT8uOQwHx2OVbfvWdE5dnh/14YtRRERuXH8P8tLqQHHs2w31
bLP2ba4rzSml/KeD6X7RX0fWrrqz2ZCMJkqPGuUgXqOUMnNc+NiF8N44zykTKwuLlsw4kXQ2m6/u
0l4ssnWkK3IVqir57sszpZKavpdNiZr8hTTKC0lVYq/crM1k7F8PhGqwK8oJcdwt1dOQGV4Sr5YT
UcX55dJAIIsgDp8xdXGTQCp0zXgE5qgLWfOuPd3AsQNv0+aOxv4Qd41TYNZwhyxdK6+4gBkebKFQ
VtVds0u2Op76dukAffc3I/ZeMPkWr/ekjyOjfmUA5kNP5irvCNyYgAIKZv3no39qqSsHV8D7nkF+
aNEm4hZGk6UZ/XTySxNW1PfZqhG4IMR8FuNh7GMZLAEKVAOce1zk06tpPCjm2W0XIcDc9SReZ1Fs
jf/plAgnSk+oPWFc7iDO00nexixKU57rLcZ+XrkSAquMfFvWuPszTnGwjxVz9IeuncbgmU6ffijH
gkWjTHdIODoLqtV8kl5oUSxM4KIypsFxQx0100VYI827sVNYSsYkW2OGIv3EUW95jzpAuzLjnBF3
42hw0nbtYYfItHHZnByNrCLDj7ZgtQVES1kjNzcLyeo61fH3BZmjjmBw+WqmTUIsMwzDvgdCxSOO
9c3bbcojztWHSQ+lhu2nsDvDb2EDzJ8o0P7mA9nQA3qgsd4Qi6cI1zxJK0+sOQVUy47BKFaloypb
b3QgQBFzftAoV0iuEjxxeWHKRRCbzEp9t31FKyC1OSGr8tFX4nZcDTJS416QoLx6kDg7lbO0G1PZ
j3JjLHjhvwlhmU90nmvTCG1UK4im8XhmMgffKuRmL0jZ0LTnAZATHwgK3D6LiKWJ551bKUE78ukg
se3IpptluL9XqPXFlayl1yJQhAt1L6dqHb6qd3bm84090DF+ghum7DEuPsT2eV2IIloAsKn8uHJN
lUKjmhnaTOl1t7jgoiVN8EY3Lh21oF5G/oLvO3IC/AKGCh0+nGy7hP/gLWg585v03oGylWMirekH
vYmX4pMSAH3qEWsiAK1ydWAUuVzVOaFPrgDXOGaynD3UMKXjOI2vijU4H2l6KC4HbNyaqA0aHf5B
El3PC+iX/C3N+DSfLwR7qCP1HP7IGx/T1RnaIMdGXV3tWevKQARbR/ItBezY0UkrXwYgTDJCxwRw
I0aFjQtUjVibGVwJZnyYm9dAk4LaoycLmMue3U3IjFan7Ozp55eLACDz0mFpz5jpAIn4M79ezv7a
reidKFzU08aINxh4cxrRVHnT7w0Hps/wW4Qfrn9LbQNM7LqURxJ+ZFkaGgEnNPml45HPvd2RkOpX
9AR7WyweqXljXKuZvG/o8gs3gHt9YAgemcBfsPp63Zilc/WmRJJvAd4dXpYR1o++3YwXRj6H6Zds
mIRffjAu5ZxW1TCzl3NlwijZ7/OLIykzhpyeAsVlwPR9EJ4yddSCbx4rIi7vBcnHyWaYSCB0dWPh
4qrumxnfv+FGgHc3ELx2Tz4yFecH4Vh+nw5IBgbiFEw6SL5NhlhPm/aBGT6YEi3px7PUYV3SNF0U
IpsYkNGGoiWErsiQo32YElknIREOhiuWzyNuNJeLc5MUKJL+SfgPhJ3c5cAPfH8e31nkiyTJ5gof
1UUm3SRr2X3gOR7x7F5U6lsqQfjBiJODbYILH7cYiIH5ufYGc93ccDqxQQUWRCHAvUKibOuHWDnD
gn99xKNdyUJyJEe3sW0n//QvENPmaatdtg19PasjvgWkODjn/T+NE6NRc8dZFAXL3Pc2Y7r8adHE
pONiGZuWpLhpaAaH6qKjV9rYGjtIavfERAXdYw+YfsBplAZkE6vsb7r8CmcmwbI1uzrf363mRuol
W+GDbHiqRjAXQjvnZMTJgm0nb0cNqtD+xm1Gbnf85fgHZkU6S7FjFZW2ouZw1bjdhw+f+pcxlPLO
ZGkhX3lpiSvbQiDxc0wIEGrE2CExI5opXbgxTr/jj4+PJpwRtrnHsuQgRjKfT8xxIuz8dbXghrSS
lZ3kQDgBCu91NoOFBdZ88Wj+kcTSfHRGjuuDaOr1grg8YowEsqxirIpKMsTsz14YCTOum4CYv5b0
9F4CyUDpteMdlDzHclcnhPwHnKfdAf9VdF2jCF+DQT0YIGZR7NJQBHr4dHlznT3GIf72KL3f0QbC
+vtIw+/V+H4OkTM+1srvJtrWzOkPN+LzkqO8PiRstbvl/LoCdsM9kHKxN+TDAeD/h19mP4oqh65F
SP2logAB8X6ar4ZXR6MGK317//IqECmxCwEZ409odV2+fhcCx3OCOc0iEulc5UBZCnTD7G6WJzEP
QC4o22rbyQ3mfnIViZbaFZZNu+jNNMSwEjh4Do/799nM6clzxJLVW/jCnkz1k+h2eqf7nG1c1aor
5l2bgx5FEuZR28LPvZX0j2trS+78XxZS9R2mWTF5igNJFiEu+tUkt6cmNwvn8hHxu7rVM8oIyG8w
4an/Hzo27CcpSP7Dik2HL14qfaz25cFZczzgCtb19KhNgWEf1HMFAcHRed55eo0RYmF5R2kgnDEC
tDwlXY8Ad1YrBAEgOi3lS4YgM+U7SOcQhkJnLlx1DDNmZAcHm64b7fucJJLuYyzUN1KmEKX22kxb
VQrLoZiAEBNk+p1mGrw8rOEwCXaC4kjr5KbZsW2OfJefXifYUsopIHCYA/u1R3wnd717WywOBhHz
Kg4rhFFUeP6ETrvLSk1TpBuCxEPvyC+NxS9xYc+HXuFgupIxCQx0oIvy9rF/fdun4EKQI99cyNTa
5qVDVqzBtXbESLQOVA4cBuaajP1qqDxAPTNQbnC6g/JSmbvwwq65A7YVZLWsPrzABu+FSf5s7Ly7
4gI5eleRgBberc72yHbr3QoBcChF8oYjQxoHOKsFNs1lyM5P+UV3UGQAYyOtCf+XbXSuXYFijrMs
B5cFrorm2Dw1R/17Qg0XkY5uVuo0B4cUJwZC/guM9+2LP1BY/wE8DNeDVdGC5iSUhAcNcSzSaEM6
n9mC/NqhMWpsnTsWoECYgtW392cmPC8gEzrk4Qyu2vhcglZg2wOt05BKb82dugbu3jh25CJTF05P
iGcajbV0HEGGlgLnS5QMr5svLu4lJtAclZk/AuSW0KkK/OWxsnfPdPdiVMRIMT7dZZJKUUGJl1Zs
V2mSNiVwfdXTEPP5Q5qDJeYF64O/cdZEY7m1jDky5qRYbYU+lXPl9JKwXAhbemISanQT/MQOuLrj
19mcAWytKCtSuXVJAGyFpaW/6+QzHvYIUMK/4XtaftpW41SDDF12Iy2hidaMy7D2Q5xtrGX/rjQ3
483dvmGJOubR2NtF4wT1V8RUovx6UDzTDPVKt/1gU3JaQAySuE8cQA/h+Yc5AwyPOlRTaL9pdCrX
VlIfwg64x/jrlrhiiiw3AoBU3skQA0BlwR60HPczR6G2srMj6aV9BsNumo71JVIW0JCWui/+32DK
ovneXLP/f/azUvkaOZj+2iSCD3wox8Fk/JmWvUy6G/hLCCAgw71YLm5vLeegC2Hi05wRI6M5m8/T
xfRTLFnWeTM+GTgMEunmW/SCUcfsgOz6LMi6D7D5DGFV8mO5jCGCXa+Q0S2uBHN/5GcSbpX9ep/K
vSum5Sr2zMvtZaXu7HUJyX9ffnlCpDpKRgMrtdrBDBbR5/aiKLvrXn87fu3aCaHKQopy5shiBs9q
aMZl/FA2SQ2pEwFY+KtzscpNU4FECASU9iM2CXnpRnav+rBSe1PF3MXXqcIDS/nEfAiNoeGqkNUc
MpOwlen3kMj4zrxU2kKC4TV24Lj1hFVkZwcvBgzeJObj2M2B8SQ4fxtTDCimB9NaLsyDgYkh0Vrz
GPaCWMjtTQ/Q4nxcF/Lm0hrD12WszguXfT20l6PmPaIKETyBm7cYLUmfYpVrRTI36gToOSEd436n
hsoAURUlyKOCiKkgDKEorx6NNTuPrBKMYiBQfWhp6SgvKMR3s8bpAJ3dQSGKMpobSXhsW43VRien
vNux9s8DEhl9ehNnvYMF5eVJIcauw+UfpC0jplg7R7Jl7CG4Xju4xAO2Rm8uFzgDPx60ts4Cryke
FTQZxT/Yv6v3uvJUXYIQ5vcmuvxhdJjcoJsLlVNMnX8l2//sb+zIXtBYEPYUE+BnoSyJ5Axh2tVX
AFilu/2vYcTjrVGFnWJp9hoZJwouhxZZBy2A5NIbY3hjYgf5cLzgOYUKGU1UZu+JDkaw/lyLoHep
zbLkZ7GqHRvNHICkwBY6kdMEgA3sNRTC5kXAHERJj1OWPElyi31at5J6Uhnl4Aunyzk29sj51nFO
mFzJaEH/eo8qaooGtGM7/wb/b8e2+JM1ji1KmPClVpSjiIJCZSf5gi19gYyGWoJvG4MAbP2zsjDT
avytQwkcsToAg3weJ8HgmQMr5PQQcD7jB+m/et481ShN274tqST0DjSuaD7yfnBMRxzr+0vD2iS5
JXMUE7JubVDKVyYJI2kEeBVLzm0fXfu3/gzaKzvIh+ZnfmRt1ZZyCDq/Mc27Fg1imBIN1cc8o/tc
PlETtoFJRrhuFuk4O1cZD7S3N2O01XPhnEdstfyZe2L8A9oBJVF2/58TMdsRP7pzhfYlNVjBx9P0
E6JOMwsFpuzD67kEfitQkvtEzz1aErduL51XC5rdEYzbefT8MyfRtSUVkJJcwir+cu1yxWJo6pAQ
9XjN1vUsXbpR65+hV3UV2pGpvqsBhFPMSTc8Eg6qwtilW81QF1Ib3VVQM8YhZZIGAuBQm9UWq7vF
HKAO3Glrma4EBvpb3Aig2W+XAqCvvzQ9LZcoETbuRryImTfNe7ttyhmfI3XQA6XLYJXtEumasWxc
TXj9MANncE+33wEPg8AV1v4wFbpbo2nGdKLJuazC3kyKUXlYFlXG3UGIyJ26/Dca2TRn95620uWb
KAHlW2z/bDRnS5KGEmyeEm+cWRBrkjSdiANbBe63grkurV3KQNYs2bUY3ub1WSFX5XwwqzJg8YmX
lSnRwHyZ5o12x9k+M69azOe0xP9mcBgDKNeoQUmaQGn/JoU9Jx7hGkiulemrgwptZa2gAtXsgLM5
sLwEwKufMkE5QNpTtRbdRMS8odFPZazN0ASzRQxSptTA8vlGiTqBP8x+VUWFNkRhpfpyER8s5tqQ
PXWd18AOVC7mb74kAVgP9EVyane1rTsK8eikXzt5syi0uHF4Vnc/51LEIgbZfiNgRw5+dS9LugFf
6s+/HKwDoN+Zcelbmrbs/omSQq8Mb6JJD7KAH6BT6I8NCBalrMb49ntxmQmXHrKkFb6SV50jP9EG
0tICDIwWgb29baiZAaXhbeQkkJdVi72ym3kSABFSTKwsbHOWiN5TDIQSzil2zXaNcmvbv9Uv7H4y
WbhIuvOpzzQZZygdZjwCE2CSywN57MP1VOMC0Bi4CAiV/S00GTsC1vk+Oba5qNtxSPlWOMX0fA7r
F1YOGqYaJUWlICMbJnI6MjhmRih7giosQ7jBmQzV3aFJxsOIYPGbiuD8PMbsbj+2x4QIlNuQrlR4
z3Zrr47vPiIll+CmmigHwPrLwnNQkMNaRVvXe4J89UMW06QGxQs+i44frr8uck88k0AU07c1yo0o
nWyiMoIk1WQpuyBbvpkVmfRJiO9eInFpLYjtpLeNliGvXZiQZLLkgM0QccVjPnk7g32TxHQc6Hho
/WSagsV0praoVCPoJMobyCnX97UWIAhNQrzOFLjLIHUQ0BRVm2q7YSsYDFnEiqnGaLBz8xFCO6nC
D4NpQQkpUtseWTGGel6Kbk5kZjNI5H7dhDn21iGGWMt46oFs2LJZUArT9OYvZEL88489ptYyBwGS
s6FOOhUCmu542Vn/n5qLyplLnGjGmObbVJJ9pO1t6ofM7D5OYlJKWeCQtMCyfuZC2K8Us1vk9QD3
sAhD9Pcy2LcSaqAe/qiBaYJl3iQTaj4+AzdSuPn2rS/pNyBs+nF4NHx375t+MgGmt6e+TKtdF3I1
4xxsfJYPiKJR4Z3tc3ZoMzFqkqcMeC2HxvEo/ofFf4X7qb5No45cYeyx/w5orgQ1+HMxKLW7U/pr
AenuZtIMD4CapFILv+gE0a6Wc2et6kJGjHH9+OLGnAdStkr5G5481RhNHNSVxi/Py873a+HVzUgr
UwqnYwZeFh27Cysu8iv/e6bw3CCj+pLJP41BwSl0TYgqaGlR4J0gxMU2xWtysLqXgh9wXv6/GGeD
T5SMY6lpN6LPcbaKybTgIIUIprpDG3c9lc+zuhUA+3hu9CBiQcnI7eVaPqKd5RG5KGGm+ixY7uf+
FoJMkc1ryumDQhDhoDhYIKjZqSQOSiFK7THZZxyShC9JD9eR5BmmaCDcabuEXEPuzL7/G5h5YPq5
w5VYI2p4fcnutUoVq6bRPPt5jlypPyA9ZL624dIRs9jUDedUgyjVJVI+JGZjczilosyPwEbePG6E
X5VqDc/kL8yiRPebMHVQnbZhGcEzd6c4nUILU7NFNwHwn6iyyvZklypfSKkRikSL8dFweu39VEYQ
VxzHb3a+WY9f0VCwibMCll5siUmiOCACNuqx6kHPHJNqL1CkyrnW8y/TYq0XNIKEUxWiOVat2Dl5
8oWv+ILdHuWiaFGYhUTQtPETdXAbZfLbqonD2XW4JPepSoozvm6sNcvWVetuDpr6vxh3TWje6vHx
G8SbLwMSElmDMVc5xbhr8dzhO5b/qg3PvFFjzl/6o2THUfz0u9O2reDj3zDhN7HFRhjOuIqFClcJ
3P17UdCrJbOaL1jG1b9rVQLmCVIqsX7ot09IRMMLIBU/VlZYOo1zBNzo5cV67ugA3Gkfndx4SzdJ
+eW+1l2NjW+6mJUT+nmWFKDLBvdQr/cHDifV3U89IaowGWALlAc0X65RS1+SRrlY2+xUivVFoeEQ
b87iFE9keUUfvJHdw96GQ0y9lvvy4DCDgMXYNvMyL911uGpZb8Am2G1VI6HGy0YN3ORPt86JdLy9
p3OdOiLbCiImPLp59/N8xrwIjv9ARg5yTJG+EHj3yehKcWXUVaCBDxGGaQad8zfF9WCazSx5drMT
2pK6rpoZolM9weY4J2qHxbct+U8TP4fTjqD4Cl70pLyBD6Nq0enDlHtTdqg74TL+lSlQCV6JWeIY
jRyVW5H18qu/Nl2tbSQ1iBxSKkiOWAam93iPufFgJJzn06l7sjYEinnx0jpZOq0l4cco0vQGYImC
oLncwExUOhNWtn+Q0kJvi8RLWfxD2xL2erjr7TuKAct19i2O8SqgPbjwSCoO5naHTats10CvBOBv
YwtJ9Oj/PSHDxLqMIRMc3L/BptawoJ+S8FVQc2UjTSoP3Rhsv6TW83btMgCazlCs4GeWG28F5Iwn
JBcX461D18+AXissS96fTcDA94NfPRTZq24NAnoVN9sszGGgVG4g7+X+A82OyYJvKZhCmsfbaPST
rNqcI1s7DotAzrhkgVx22111YHe83RRZclmqnDWgh4vP9pKAzRO8+OCk/fryZqFVBv71ZOKQd2lz
z1gTZ4OkfGKY2UMAqCvC5lgr9Uusdqbk9ZkTsjxpWJH26pv14WM5NJTxB05uD2oNVDyexKCwrhh+
43DIBlHFiZESCNVT85j4iWcK9QRWqOEDByNAYPkvfYQzFOWNXqvdMZjqsh2yK5Ne9AmazkQnnCrR
Sn6s0gpaCuzYdw7DMB8D0xRRH9f3TyXr0s5XXa+sOz9YMeMOaBqTDSWiB2AuAM+NGBEJMNPK6Fii
Y1U6Xn1b7uJ65VVazGJqOO+JDeQ6JIQ6Ofc9UwWcWAgWdCd7rF9lEoWw/qaXraKiYt36CeNx2PkA
seqKEoG2q7a0kJ0eBnryRZ2BvSM2PfBwKAVyaTk1fcAMmYLn1RZhPmX5TMr7aNcIjyvlBtu1ZKhH
YPMck5nwNIfVHCqaInf5gLBz8YsFmMNqWbRp1dlHCPvswkZ1o2nD47uTts07JVddwxMiDOTiMgY+
c1y3H6fhlOnKT2yhMJ33bT82S1zztBM+iEwtPCiuPEvS5A6+1SFVJ25ozTJJ6p6Tuy/5ChwUqXsj
1dYroWv2SnkRQwRZfuClYgDLZnXsSJ2VbHMq9MyDrKtLE/BlxH1ahstudrKn/tFtdCVPg3lZpX7P
0HqTWWOkC2oENS36YS/9psm86gB+vcPxzKtJwUIrrRh4SfGuIBOdYu4UW2ej0ANZabhzNouSmzyd
Kxrinx3ZTTWXgaS6/CVtAWKkcZ3PLylcLpioX7x+yJMwRRFdrS8ctuurKvx7bQAjzAuAhMTBYxwY
CF3KG7pPoPGvd5bjGyIRITbKro4428mBYtFU4CoEVskMmUISvWES/HxQsC8CjEvLaSnO6+F51RGe
NyRGHzd07Wkf22vWH+ijSzOAEFcOdDW7gd9X6tzPcdqhx6ThKhj7pSw4dyoQZEvVl9cEon5H3ywF
1yNiNtXCYjvI7aVUzebqMXu2Ww80ys5kiOY2Tb6pq/+hQqvJSbpuB6lAXgPwr8RijqagnHe3seu5
kL96MMRUuWj1UwS7rn8+ldPrIOCpvFP3/r6e3LczjUITiPAlCNr9NadVADTxzMlHDnOoY+b5D9+m
btWeBqq4qs+jPvQqv+fIOOgmv+6ouBx+Qy4eTRd8JU4BBbyeaD0/37rUM7SFfBigspDNgpT330z2
3MW94xmSdCByOQmd9LnyiWLN7Qm9Saf1McuQ/6Ko7bkbdu4xQccjPv5e1YFmj6s9yaCEKJfMxSlU
4J1OpCmdHjcarlUR0cJyPQ1OgucYPFr/C4reQ+V+z1Lec4BrfcMr1+dKZU5ECzwg2tJ5Wa7Iio45
gZAOwyY0rhPAQksG2pqsy1UAmRf51eIvGXrX/L9DCPQNv4EPt6zC7NL2+6BNWcbzN1sPogctGPIw
p4qu35xK1uyuCqcvPeQ6ZGoXr5WsUlF+JFOxLgOC1HVkYcyw9R28KELjU0iM/WFV1LDy0lkoY9TO
wrun0fe+pjkZpyC9GbiMxuOm0dCtPxP5pK/6GLh+0MdVRrq29Z9hML1NMFqgiDVj6D5Es5F0dyKf
yWQKkx+baJVa5xauYduoOsSlpA9Zx1Cg7JJ7YkPuJww5VbHDCd3GUc726DrHO+Q8h3dc5Diivr/p
/kJbSmLls8V43vrapsRVpg/ue/08MV1aCH1Mhgb6oJxCwQ8FLf3IHp2kTyJsszcQwF+CdpPeW/ac
eIix5TEpjmo9kjXDHMu91sySvQcVPf32At9JK89lYLiTOTgpXP6vBVdoUgp0OCHkewVWgm2rcEKz
EyfWJBlCLdtcgvoOoVIbAjmeHnBMrdrOxLBfJW5wlaEFyFDfccHGD/aYZPtblduGWU1/p3M+Tl1P
9fyglBTXjj75KLA9SLKytlPNYFN9S3ToXjTR5jiE5awRjc5UTV5EGmihB7djpkt1gND8LwQedDTF
fKHQ1S9PKvWCzR8rxW8x8AJayPoNSWWeiQ+KCsylccYCNAYa36zuRjuVtbKV2s341Tj3Y7T0mwxR
cveIwqGxGze9v68R9DkUhNQc5xbBEnH1ASgJDg6MbtnC3+sAVySYeecUZMuoPUh0cbaF3zFCmf2P
yftFI7jujuneaO2yan9DKNBlYQ2otelafAurrQp+ePjSHhmiprl9hSdt7c9XxRU0DWFQsRhAXtcN
H/Okqg6sF4hL0ZeMuMtET3zi0qA4YCuoDdK3xRz7p/vU9h65wdDjNXBq38aIvEGejCA+xyMtOyAE
vQUqHD9047wfj24GG60Z+kSK4TCarZhibyhYg1xhbOPTo+FQ9+vWtlmoHdJvf2qRYWc64aJop3Ga
9c9nM1TqXBKnQpU3fJV4ENxTdohZJS3Wm9e58Ri6ITniyGqhfcrjiECvx+ut3I1yHJz3t+xi/kbn
xQuTsqZH7Bk/CKyxeDNwIKxrXlPPaJxBH/76GpF+y+HbKOx2ICrwwmjp2tiN+5iNgsbyUDzxpysQ
OO4RCSrGi/ZA1ywoCFYp6KwhTSI8EzZG1c04+eP7b/OAInYPaqpEezK91ijquDLVY6EHtoncZ/1s
UqblT2EX4EcVD+B85gzcQ8uWhyIAKgE8wGyo4ygPeu9ZHm/VGLN6zuerc5dWnXinlJ8SNJNtFOE1
ryLSHTvfUGLWeyoq8yepl7AbBFIZIXL5GuQDJ3hfXDzEbXFl7DfHPAJTQoikKRBmegd2KtFLo30a
uxEBXM+6Rn7t/fNqhPw30DZ1G9/qJPN3cAaNXwcNZ7REh2VXRIeWCZxNOaKTGr9nAVGLf33Ru0MJ
kY/Q6rxcJ06u2wS7mUygbK1P+NVxBxzeb6VblKabxRdX+UV1IVuo15A2T7YyTSjgL+B35oMp6kdA
P9N0+ACiOTaBCa/tSmravV/qG+lTBZqBvUnaHcAztNF08IeohxlUWlL9xk58Ze/xqPkW+gnLCJMx
PTzMNVUvfRtt2fbvXbC2BYQIfHvlJo/Xcyf6X3CnhIcMiB9VIcgPBaMtTjYSAClAsEkVNTwufy9l
6enkz2HYF3hPb4GZmjNzSiX5I2AT//kgYyXl/KoCz/q4xLuwEBwVXMbTQQpxkRS6lRmd7xiyNN2r
f2COddN4F0wXxKNLRW4eaMZZdORi1tqB9xMwhLgTjB6yIVsyeAkjdApIMxfdQeHir+cEIhNRmC57
OwR0suggLt24b0wlXXPYiSoHoiZHcHcOoQRJp/EANzaXvZwj2TO3QDPijGEa2dkUaHOfQ+22prSq
a2S6vlf5HMLwdRn53lmqe6o9htM0XkUjEvi//8V93EBfGe7WDCzmaBdv5cMMwby9I+Uer9IVGSrW
bYFU28nIXhaWPE1VLUsUC2Rk1VG9mjbACYLpmOI3gYW5poeEIUN557o492J3JUJ1DB3Y+QjMOQL8
kkd1GnZgyHVsjZ7WUBoigEncDFs83HRLFxQZEXEIeUNHu5Z+2SVU+SMAgmqAdYp6cBxRUVxhqQin
+NK1m6DYzcNas6Pydnsabx02ZaCWQYE5krN8JzBh9fIOEpDCOkn+oF5l5r8T1OExOJuC/AtXN2M7
DoJrD+tMRqSr5Ef4SaEZzPuGJNonLtbtFroihjZppn5vs6/2A+Us68HrS/jLjoTm2s+0cEn0UV6T
acPI61Tgyqi55PgxTNivPkGqorrG0PJiLEOUbkfeBBahYTBwFgKE3tV4dzNw5gsGamy/x6wuN+43
rCccC5srs2DOqHch/oBU3AcZdqMONPbN9PaQcn6qED0Nk2XkBQ7kHfscQNyn95q5f0BIuAiYFkXD
H8gyngqM0kViOBxMn0mn/ddbubbzv+j/nuLgbs7+RzU4xP0jcwC8STxI8K3pvjGo4RpcdFkAf7yA
iEDmYtUz3gRlGiHXZLDo8fGzPAUsKPZP36dP2A37nIgK7R5NcC9QIhvyhUyesBykVCWIOsKMXGTV
pkK93yBH0O/aHSdwwrqotEENlyzRI/JNN1OuzZeAjGcML1MDih1lZ5UmDKEOUS8T265wGC2aly1P
xypTrzaNWnF73AJkchODNVJKziDvdOdIqqB9Zngn46DD4uvZD/+lcDKWhaXd6QUz4a9insOO+o3D
MHI4C+N4D6W7XFBNxFbumWCypo/TlDl1cD22C3eULTHo2KeLNaIzIOKHS5mFXf/6BLcH3kv9RnGA
hHpaeoMCL1H4PmZUzNtAs5M6df3QSwlw4/Rdp6YZ88TyycbYGpyQHVi0aGRLqfLNRny3aLGuKcEZ
1gkmH8+gCcQBxe5Jf6jZUlBlN+vnc+Tyb3Cy7ztoIY69wdH2+6ftY6XK0EZfRIPVByWAbATC0K1P
zQtVnRxlY4jZtL//aecUT2Nt4WmTeNlEIsG78m3iRKl95Q3FM/hkrNoVTCT4Jwp15BnR3M6JYZmG
ALRocJogspOvPImMJLo755Hdd4v+kKS4Zbgk0n5uaE85jQWKp4kwZAEWefxG/JEJRPhxnQdh09Nj
2OYeozy5oZGhVasAlVLbfl7MbwOf/kqJCgG+95F0zKjXxBOU9RH4lovTN1Ozr4jsI792zaVi9atj
fVlLudhKA14Vgtt75sHGsF2mBosvQHJE9ZHBsWjMA626DUizpbDg9AWjZ4PccCc+co3qtO9AWvmu
cy9aYtOWNTJENY6zdkiDM8A7AE+f7/6uEHsUsXlx4wlX8QI75GspV0PVX7K/cjRItsawRYWSeNnk
dTikhBbmBYCRHWphwmONZSzKiWS3Jw4dVGoX4tOlIYEmu9zC+PNXuzkEfJj5OYowM3eBqScoHbCZ
5z9erTPmo40Ln6BwyyqOPQKxadYjxeWlWfaynuWXMd4zvh6EMU7bl4E9b7OCoHUlSZI5I3ORFQ4A
rvWi5hC52m1x08AxR5HG6xy1pFA59VPqoUFBxFYZr0SYWPHS/jr3d6W3NvlIMSHDbdIBj3+5R1HO
gbNU4kduFfPcZcyt+G71U1vuKpSv6oXWCWGYUhVBdEWP5CJ7QxvoXfqrtZrbm1n8pJnpx5wM85rb
UbhqrVPGC+kvH+CQbzW9TRwcBm/1+iWXKn2SKf9IvliKl5wk4mluAksw5202VlYY57lLRci99VAX
xwdeICiNB54MX60sQH6IbuWRn9ymhBGveY2YZodIyjwwYqJNDBHhb7NTn2XHR4opKiJorTCKLHK1
ZTi4hMc/ySzfK/kHqLVmFClB1Qc6AW+r7r4LKM7kiomUv3sNmsZbKi6rJpNFW04TIGuyseEmjkS8
GvgiPf+OdFjE20+Ri/QDzAhYxpnLgWdiPOMfxvAH720pZoXT4Lgag59hYVWe7I/Q1XA+fAiNHep8
7KiODecO0VpRH8PH1X+n3Xtc43f2Hc4/eOORCxJ25OQ9zFk2IJ47oiYNgg07zLBtGHQK4oxxl14L
OTarDEyaExuPpX3A8OEKxyqhodI2iB6iP7hTH5yG4knVEXLwDjXG8jHQljZLpMDVJsiuOOw9hKvN
Cq2FGGlbq8Y/cejULqVl/YH7MlLLH422vOKtfkBRKZObmmY82t1h8lMVjjju+UAtcQBPGMDE299C
92kgWr/z8je5SmeqijRdoezlZSYCCagzpJIFhqg/YGOBhDagA7GmQr08vJ3BKfK+zRf6coHVOPwP
c4v0L5LtrCLFgl77qajhadUN6DdbkqbYuZqm435fHFBMd+CByvyUsndTRIhzjwKPRHFcGEfxvTza
4EHzZ13LVnhet9nnPceIxfF+HLS4+72lGlQBArYy4sM4uRYLKTB1kzT66QMCRe1HkEqXv+dDH0Ov
nPpE2Q5O+rS97XS/wQ50oie+RC2xPXor4WYBKQThD4tBx10ZwVTVCVSLtC9UF+c/qeWhiy406Tto
mEZOlAZPbyMID2vgMEVpJWnN6k4H8O3e/1MIspQFOwjiEOtiBGBmCKSDYbOf4y7mDr+Qsh9xzQVQ
ZCnYPm+26v7dxl//xQFk+jXX0bg1ZUJP9LV0+LL3DiQZmir0YnmxbGgSsWo1mmcgPac80ZKpd6WO
YZLXez8irXSxpxoqkCm5pUxm6O1ra7V2P+21cEYeXY2TSClAkI0vNCMrItozxp1zoq/LKLxwswt9
KXSxl+O22gbD3uu9h7qlbLmwBJTGdJac7aos7/41c9F+E5PjahE7VT6j0tI1q1iprQcH5/28Ru+2
a/KRABTJ646xs/NuMKzipOrt4j2z7pdAOJOkJhfd0fYK8x3M+PD5V0t1bd/i9EH+SRk21JNEISVW
86EbNwzvgdBQWDIpN8Cc58fZ8ZmYBxoCH1OTCA/Sb/jGNir1owvEtikhDnaWHKnxZH/AZ56jOoye
ke8GKdzznVFfiS/fzz2DZLiGH5C9NcNdHAErA0ky2DLVE9Z3sUZEe8AW9mTFqTh1NE7sNBlpxCEk
/0jpyraL4qillpdN6UFQGOs5GyVgqjWSz1DXA0p2qERVYRKDdiNs1TLWApBEUuvploICHNOsjQz+
Iq+PRPY56XrnFMhUwLmtrCOtxqo5UeibF8U9fdTP1XGCWlxcaWBn+/HIx5nsGnEgiXqA9Kk6YOH6
rAC3xeNLeeqFOyyyuXDfq6zRZbQRnVUoFs2d218Is8finCC2cXvRB2AxiZ2df1+Bxx5UXk5QDk4V
WdeZjhf9kRVhNEKRPSCRhXAaO0Jhwv1yaB3C7mN683SY+sQDvrYkBY4FUy5HJ18zvD3PaCzz6IfS
3dpqBgnK5WqOA3YyHfiiHMKtLcE/McgAta7TifM9So8r+FQqyn2q3ACs5lWQbTctXhgnFyrwf3uZ
HTsgnmjlaSC9hSncfQFaV40ixFDundJDTgulLKKgm0Rovq4KUSrDHXPt1o/Pu5ovjKIVBwPumw46
9le9N53nZch/l1Fj09FbDTBe7iVMyFqYF75Hzq6tP4Jz2hGrAqwjNcVpWf2pXpyxk2VWMBXJwZEC
LHEml2A0Eeq1GQDITLOvzciQQQHKi+87LoyTqmqTw+YNOKlvrPjXjj7sWf+Trr1dSneu3URELpja
Cjlf0RHER7OWpeP4vIF6ErSq7coTdVqwZ4I2nBvOUKLKijuwb0Nbp5Eofks2UF2dyK6ZbueZzrnC
T24FzevGddQBM0ynhLABkn+2GX5Hnls7+o01lfsE+FxYMyKPpZ5H/5SwovmrjTW6fssJeFz6B6af
cLuNBmp8eB7qsZ3ocqzO+dflNBYOzvbfk/YB2o0GBiBq+xSLPZyy6EEdPLvj+WnBbe/SnCtOTUU/
GWnGmbFMyqi+49vt+KDmmpyTNOm4vsOREDtpzL0KJVXWJa/NMQuWBcEZpty2EsOSqyweNHizUSFk
EbXaDq0TWWGR7JKfVtfuIrogbhG+rVAyv3ydTyQP024wNiY6JFS3fz78/jPwoRRXVhqGqPv1I6JS
wjPF4m5syCl8Bz0d168n5oZksWPW3pplJkwxQbNOLIOLd7qQyhqTBvwdyjepBbvyRgV42waLOqcw
4qTAenjYroIVME9KUoGLwPKYcT+thlg9TnTzA2GrGWndG07LTa+EX9HOF6ez3QZwxxKMrK2v+KNf
5+TL8yHD0SrK+4T84fFsGMz3SCJmRU93Q2a1R5RpVPxzOyG0qZH3JaUEyfHLrpOx65KWy62htCm1
AF43L2SBpBAIpDBt/9YIAZ992o89gjmlxfucpsMzrMwjrOl1QHlFjCpclErQXd15R5Uy/NjEoAJ8
yp3fJhuKbX/wKMrHZ9GKg1Dzu7oVcG50ip4rJ11KiFuU2OyKZIaIVIWWc7epfIyCWlKIRxotEhaQ
BoERhSN9Xijgqs8e8X5vNXGxu5mNBM0i8RUklMIv2Nun85rACh2AR6GSOIOsCM6pQdwFBIlJPqJW
6YZgpjwYidZponH4RtzBjXbocvbC9wOvV5De/P1LxEHaHsl9f3zrQgyxLNg9oOpGCXbv0SiWj+Aa
DP+o+94XrzgCOJBzJrna7HsNdkO3xs4bK9AoJOpv36VGVbFsHYh20fi2/QKpiOyIzAAkvVrqMKp4
fuChBshN9N8MR9CWdnQQRMzOOVtlso/6PIWIw1PeisIhKio8GpIMMPmHumpapsY+mMEJYmkQEiEE
TVtAYAO8N0uWB7y6gAtKBj9q6SddKmTJtbVHODJYrOjp5hmqxATav1PMFQNZqLTl4Cma1KmGs0Pj
AZX9K3gHS1ujmbPF4zFh70CYGgKbfko1Dd6VFKtlbUmsaOEVtx+tYCbGHPN1fHszU1NPQkVDQrPS
IM17i83TJlo6/Pn12DNy3LprygR/VGXaPn/f7/xegIREJBdsUKeLWIYJyj7QeVh4Wxr3tkh5Orta
eA4jvp3bsJqDuU2jbFYEpH86fdWaaBPXQqo+GGd9Ve7XNtjhLLG1TG4rmgPGbK2X76z/OKTUUQpw
THGku+UlTe0lvjv6DwsAzT6x3sX+l/9W0qti0srlhXDqQN4jx7CfUKv6JvXrQGaGkjXYsvtMfp1s
tuo/dyYatFEAmNNjUYyIK5iak+6Du7thN4d4fx8cAC6mNe4tSUzJKcXJ/UutKnziSYVJHVdzurwV
wOgyPF7858w6dl6X9m8RPUeOYxYhWbNadRy+6l3zVeoa9PTRjA5JrRXJSnOY3sQkk6XqtItg/xvL
D9ErsXic7RNOngYCNizS0QziSTcPVtyBeKjn2PHvhw7lDMDSrXdyJ4jF0iV3Lr4kqWBb8JzdibuO
B7swDYdcin6AKc0S/7xG09qSjFltTCqXh1jZppi5XeBdR6gRwrymMJ4/3/RSUybs1wnrJXEiap1h
0eMTa+VPbc+5H6z4/EZWh7PYFubKmj4C53mh8oLYeR0rJDRYqMMm54mvl7Gj88OVX53BSHL+xpwF
DwwDgjR5TBODV6nUIzw1OfpQ4TCmY2lhtd2/6MgY36PmPjn6SE2yEb9F0XJaGnuzAgEHrvGaFpWm
C7KhRgIgH1wkQG/w2Ng22EUVE19tjYEn8kQa28J23rx9qVvS3F/Tk14Iut7dd+iZyAPRBZVcUFBs
lR0m/LXlXJ7VyVj/Wuvp3WAvDaCCg8wNSotDsqA9XFyGDdXye9+CXTekv8RD/Iy/1uzkRO24xaUl
ZohCZpVc8qxMECaflLVM9GVmmJbABkZ6Dg2VPHANyhUNyuWakep5B2l8lnka58m34n9HWvW7mPBD
7fPHyro/Z84zbqYjF/XbnP50XP8N3e09L+qgE6hO5dSiVKQa6fuMMnhwt5zRjP84tvTIq+2Edvpw
3SiJoNjvxtkSux6x6VO+lVSNcuQYBh5y2EdJOHUQnkOrkcKQE3HJJg0UzZesA6hsbMLD+R2D7LZz
pcsxSafclmfrL8o43khnL5kCyN3KVufVy4uK/+A0xue42UJos2UNpA3MyXq4RfKndFMgTF/6FKgP
Yto75zVAnbWBODnn/XBVM7tHEvhMVgOv7Rjo9FhlpJmWdz+lgu6egnNUuk55CZ7i2fLNkW55SYLO
jmpNHesT0QS+7YZHrCAYv3O21dG9AJFuopYjjg7EoH+NePcDluRo3ZUmzBF4cJgbqoke2o42ol/8
XgPHA3IpUgwNhLfyYMgHIpQSOqgSs1X6xblhSz4jDDIhfouv8tCwhwbB8SKNVUDNMJnwc5tDAGt7
Tp0A7gR2af7mBA3Ii70noq5+Q40A1CdoUHPsLF2ZXT/Ww9H6SGgNyzSmxl9UgqPy7qo7RHiaokoV
LsbYb/dFOrCoBpjbu8PgYZHXRmJIKpnnP2CQis7Gq8vHordWgJ4Vb076e/Mp30MUCGokby5d9aQn
ZxiVQPCuZDib9A7zvTdrPLt8lH6r0E8+A1kRhe2n4uA4Zcpi0UvnzUz3EnRvZzIAIcmcDQMyjSn3
ctgQE/q6wnvkRDd/tIzwx+I+lEbFSjV7VMmQpryYd7GhL6toUerxIRpp2UPTwUIVfA8okQliwoYm
9lccIp9DqSTYg6tjReI3llL4W897lt42wu8iALsgR97QLWw+ecy9K50D5WUjokDZkhNsyExbmmfY
f4+4C3Lj27zFqG0aiKTX1aBrn/S8X7TekGCAjFb5zmiaN2HltYdmieD3iCI0wQfdVTYtqQKGakki
5CClH9w6ZM1hQAQtej/vxuquIB3wfaTc30sA/wIArpCDw4SddkJvJtYN7VsYEcO5ZMIV2z8QvwUt
Ew2u8/6VktQroRoYcsV+n2WIhSj3GxooFAU1UCIAbj8KXnnrrIiaxq1wPy96xPoHjOsKkXPXJhnl
sdBkETQmukI6ZvVbwMKSm5/E899wBeu4bJVTtvoThS82ZSkMSU8MBryQco9IHwc181OMUjxHTMiR
eU0HM2hO5DecSGHYpUtbkJ6/tHkNnbLbuGMs2T42K2uzxsadymcvTVVP3vD74YGMrqQsc5ETl6XO
+UedM+8IwgojdVLdipqbNW+Qh2UIWzxInACOTmT1eZAWK+Gw4RDn6p0AzA9JW6wYiIAyeZW2E3vD
ALTFerJ/FCYw1QHZXtgUo7onwMHoJxTQu9fTb/SC/9Bnl8cpXya16WgvysCPYyDWK7fzKYPxAsut
m69yqdGULivM4MaR72o/e54WF4YzJ2U/3j9rCsx8QrwV5Bmpa7upXjujhqchxrmPSFIyyfb+LRIJ
NghZF1p2ClAN2YU8F0FfK4YFTV1qEgu5n13PAWpGHg70WDxYYTsAfJqUrG12jt6W1+3plWgp7RaG
Of8UyV5vzDlyECPmxcepJbA5E0ys680kzAVfec2BhdBzeNGm32eBvI7uUst0PBtDMM/MFA5655jt
bTrFLPNnTcT/YDSpgU9qOJ1H16EKxqmE8DsOIUMk47vM1xMS48MIBOGUO0YxmdUEtbuAfOIUkYu/
ICDSldKj0uqplnTQmOb5NPu0Xjg4W43ACKt5/fWgVxKiIUmd0cfUfNeByWZ58QdSenvn1nNhz/RK
43kPg9gIEmKz96Y5SgGb2A9nQM96/2goTu/zT/gIfGTLzDq+RrEdKQjw50ObtaVGv9WPebiDqdUI
wX+mIR2fFUlueIGXhH/a95T2rfJ60fg4Cah2qdsDIDdh3sA2FBtRhHttUk+jmdNiaMkZXR1vlFak
bfIrUm9PT3riXR4MYSd1TR2egCrSlmBlauLu+TflFRBheNSQazCn6e502RQGCNZLWmSoyLccBBgM
WAxzZnxJzDRMDh+iLIsmSfHrbS0Fu4Rc6nCtrYwdp/3RuTYeb/Wwv2tkHS3sTDyltihL6ABKL3bO
Ow/IPx6kvH3PJ3dLGFCdJ2QZQOtVDe9EztvC7DZspX3EGumeuIaIUYwltCDqpHGCIMPoNqVT4KOQ
d5b64Q18jlthXo/wG7kSRhI6a5x7B9ML5p9v4UfBO4v27ss36fZB3OQ3Kr4754YqDumsdnzN0y+o
/genk9BHnLwhULk7j/B2vc9rCcWaNFzPGDZeFGpy0tP7TxdFdnAeA95e44sEhyu2wtcKQ/tPMlxN
5KjLYwqGxnO+7e7CVF/unGaHD0E73Y/uybEGZxEsBZ53yE7Nh3c0g9yT19SbL+VEoQ/xEQ8gPe5l
OLtOn2QQuTcapCZkYLrzy+/8UxOLmYuMJDw9HuaF+GKOUZy7cL+GIg2XPf0D59lTwCJyJLKG2B5o
0X9oXbJd0tUvD7MHIi30zPHC6J5uCU8YQvoMg4ybhK8ivpY333oTYC7Wl8Gd7xecF2YyM6OXKMSa
6y3Zr9Y34lMeTb+BdJ1q+8DUYR4uAHHJ3SRS0+bSke/ehlEsSXXXhLb3azzZSRYs3mLQwha1bDFE
NrXp9SEUGgLq1gmYe4rRk5mLTLlTgM8UPpDeYiE0+kJDbJP73SHmk5jZGEOOHBZPOywNniiXQamU
tBU7wQRWxczGj0iSuXEFyt0CgwZ3mveirtJ1oKyR2PBUWBVf0iGfo+j4nt1kVLW1VHHty6JAP+jv
fAG7No78htfYayRjgckSthTtEUFP44/3yGTK465Lz7v1hW8fogq6NkVLHdj5umdoRrdBb4feWFDD
01jHWPfze/HQpZ0k/TBLOwzW5D6Rxf4vjhMi7ReEQQ7FDETaD4d8aCDZPbRmjQkojDVtU0Xwh3ka
aBl/OhbBW+gLia3ip+24l8eYuFACJZ9hM5a6y7uVHoK7dpa/Zae3kXw5rE1A3eqP7JE0uf9rjjve
AFkTi6L9OcrhfCv/RHlR/IXrw+JISSoFrkaGfSEWVWgmRVJyc5gOjjtz8DI07Qsb8zxhtilCzUFm
fYpLpmorKofNuTKnn+rSov9I+C23aviYLBOhVre670q02RQep6eobQ8wVw2XzfYZqyO5ZQR5fVOE
7Pm9Lpj2iprpCaav0P00XJJd8zdSlAy1TmlehFJYRzYi5wyGwA963RMhx/s50biKruJ7G7VUHTyl
44EvJGgSYGNetkiqSWG3tX0dFwvAquFBfWSoUpJQs5yD+RWwoyeaWrY0BTnBZZYwSIGsUbqtn7yL
uUbhWqNy8372yPTYjaVBP0kCxCq4WnfsLc/p5QPh0BqDTlRX7e+IO58eY8h4UhMee0A/3Mfa11fZ
v0ZYI97nRVZtq6XHO29tyJZhgZGbjrDVQYV+etNziMcSJ/ytJYrPpCS34cgyKjd/7Tl2JhrGYEbH
TkfpBn95ri+dKbTuXFzV66VCFVkHEcieGVBxGWeEKI0rS7f/X4ftdfuw7gw0Mc9NEwXuXp2POO6L
OVZzMHyoxVFEuzoH3ereG0Yd9/Ev+Jdzca68aXBnpxqC3I/O4Hd7F8e8jKB4eTpFccugbYbbdER3
IcQMb4azHfiO3jCM2EZtvm3djll8CpGM2QgAg+It1O5YkGKqeE3Z3Mot5a3BFXf+Dh41vz/gmlCA
i4uO2ul1R0DXyEvmD2MT+ooIh2TPEDp1I/oRIwvxdoksbhVvT05PVpKLifRQ4Ude3ZVMmr4guAAQ
IyHVqZxnUlXAstAzXkta5aFrI3vRmXLrfie0M1crwRhOUosqzpPmlp9p8soURDABSJPiI+b92dRT
4Qm9xk+iIVzw30GYK/lg1wbCG58kDJcxoz8xCOB7tREkewrncnf1XFcbAPaxK3+4kaQ8qhwORWaw
ezgnRglbM8RIeKkI6QngSLsE1z8BTOWHhk/9aCi79cuzZbpFy6m/W1F2Jbpq/PFqq3kWZ+caGzwl
piy4pP/MClMrEW0/xiLR8DGISpERnjar5MpGQFreH9faIwAfAzkeCEPxVaxPua5BhR4GKPkCg8vX
qS4BRJ4LZOdVO7Vxc2CGPeQEXb1GrbAXdlduxK1i2LolnofdZx7u0Y9hxCndCtdYLcmRuJro5g/9
pfSHMWmKu5ysZhJG+2KR82hFbkJJwLsJD74OFnqmoXn/5r+gLZP7SKWytnPJpAXr5tNhUhx9BEru
XoOAky+Q7tTZ7ks6zrNyznGRJBFO/TFbX42VD6pQGDUnlCS7tm9tDFZ3XPIVWCUch/GzDiiaE4AN
HV9rqBoiB5DVLTR0NrPl2/fiZvVecS7SFw+hxJWJep4Njq+Tp1yg0Kmd6WTO5bifMXY5PBVzLQss
cIc1z5mIeXIguJFiXcT5lAm/18cFU/BYQwGoeMLPHtGAWvFXiCVIL7LOJvFS0ffU1SRprPG6K60I
lcZ03o9M22rSx86igJBnvaEnXY4uhSlZl/jyey9x+GuKgCErNrvrS3s7HXDNJQlU3oSjXWfS54Sw
vA/jc6Lv15YEe/kOmS4UgG86jw4fqaiY6twIiudGS5yH+a9ftxS9F9l+1WDC0i6r9N2e7kJTTyXK
5Md+s+LCrKgFIZUp51oSufwATQ0yUD80ipKLFS0H593qz7/7u4keMJgYmfzraViIB09fLcK+mDXq
yxEHM0WwVlWDt3TKlLoRBsTimnRIBGgC8fLxNQ6Ghoo9wchzUk+jo72G4M2SotntWFAkRD6AF0a6
HT3q11wKkE8ntp1HG9k8ZBPojuiNdp6NwLwfrJuVb45r8ryAqB8NFh2YzVaHY75pE+peCntSkCxB
tNYokANrqBCHmTDKjjbGBsV0QFAahwZ+LIDtgVbmDdYkc3Y/RgI5QnzWsomk9Ingccbyw9JiYgwe
W2BvWvgKxNyjXhY594f/hFA9xq06hjq8l+iyKZkLlrZCMDlN7/cJfeXnVZGOfUzjNsnAxkp6Y+Jo
WDcG1qqBOW3vzba99Ksslr5z98cNbmtQIvAKNbn4OuLxQ9VRkNct52RQcov8+IMXJl8JgL3Xo65o
uXXbjMIeTqf7sWt/Q6IgBlqFUKTPz+YGqbx84mIRsQhxXJZ4/33k3bXO0Feu6E+zmoEwUEXHWRHS
j2phTavY3UwiSt4T6AUSBEAg35hl4NxWQFjC44nQ3a51pcb26znLNQ99ePldK3uYgqAVPiK4Ml4l
MaFXnVT564vtXHTEB+6vixp4tJuvOZFcDc8aLMJxmIKRBu+49/swEUC8Aq0QIXcOMb5ENrJnN6U9
dxo0GVRZOb7iH8ULDV6LzYsyya5gxq8cJr6PC3t5IfjGtoeccHwqSQdRI81DmR+bszTcYPnbIQ90
7o7bd9EXE9gmpNo5FniyiitxIRAFdDnhbP4U4EpE5exRdvpTwI8xoZcKurk4kK5owvhx1j2fArCh
gC2ZTwS35LN7VllzbqPjwvImk42XGHPkUwVfM/SWVvOJRs//LFQyG1giQq2nLuVjIu2OONhjxaBL
LuF7pNenZJYblq+5//liNo1nKj4Z5PHf9QqIcwKo4nSneJvOq3XiXbmWhomXSxoKPUMVZ34Kc81H
hatnJ3W6Qw7EpT/X9jffzGVjWfauqWDYdkjCW8aTpNX+dQr6YEVFZiURUd7+xcdwhDiUkjTAYnyc
q9TahrmpkYt6QySOd11ajXEpkqhW1Q7SRSwkYf2Hst6XkKMqVLPRJ5NnY7Od6WtniD7Ppcn+vOmD
miIVeYx7akW639uaEXUQ6aG9omFrpHcolipNe2uxMQ8EL4cmYc7sQ1baraAkpy3yf74NqAeGt2Em
OVq5ZjTkFb8h8yRtotOQ2+p89wzbo3HD1yyBp+POjUU/Bj9cEK0vPOz56jactQLi5e414HIooZPZ
/4CwXvpHrRvg5AMc+YwVNBNf89sI0AMude+77VbA2Qn20qFw4Q3W6y33xyfVQRdWgSddUHD/PjLx
vKjIEQCGSXwxtxj0KNu87/ffwsE0afDWM3JXMOEJlkDMfUXHo74qU6+ffdsEZvqpL+SPu4u0di6g
k8RFfe1OUYBvyv5bA35ddxisMRLMwE+FAHgjygDyzbIUq9pdlvyYLiEAZuwPDBxEzFYpa6cVzvCA
TPknnK2nuJDOKLGVyyzyFlC0eGc8dQLe94s8tDGK+fwnk/cvFhKr4oK+HzNma/Quvr5FXrNE8kIY
Me8kjpJo2EYkEULeTgUFfd42QkYkmKU7dC0zOSdn12123B2mrFQqRkqv9WnxB1VxVuTCvARZU7o6
nLlRvydnspXOp0n8a70xeBYkY6HoNrgdakoSG70at5g8k9FHZvxF+xc9h2JG3FzbIp6KS6no0m5c
RtXx8Jiw4KTDgiLoMHx8lrmKpOx6bvzJ3I1B+SywIxhb6OjvVY9AfAohMFE4Q6qWypTiUIcx1edW
yqAuz+gaaCH/VVTr2FFP56PnkTb9sVoPispLh9JptMU/N60+6FKnZlzyzT/qpUq2lg01fBsnRfFE
5kJ7r88HhndWLmqk9618jfvZy/ucJZ46jHsBnQybZFX31g1qrxrVJvGLwHaqlocUvohiGkvhhuK7
mCZkHtAzaXY48KQeunJpImx6DAnyqvtyDr0vyoAuEXSGvbxzxz/D1+sDnoHMPSMdG3zyTzLsmue7
1EROjOWt54Whn4d5T/W26Z4b/YxslT6bVGjw66Y26uo0gCQb+5HXSCbIEhSdTE886JDaFWBoLb4v
fHqKPwLU5yVC/MfoCajZFii6dLxywib3mWLnZ5SGCYjNJz6CzEBerJ8Nme/WRIz1MNMJ8gYQqpQV
wzgA45gJjErif/aNgFfpqCwki66wz8Ieyik1FiGTuQFd1fTYYOEy+1Inc4ng04pTjDbMRuWKv3Qq
7Pbc71ZITRBp7U/D8znSON/UKqd84F6Q6Eu4sQiSExdhPbN3f5FkhOTtAYUsmmEJArTqNbADngyN
UWfS3iMOFdsNyXigiXJw0HL3IsG/xbrRjzzmJ/J2Vey/wv1MNUEsY1d+3/HNFjlL4pZC3QvyATo0
RhJL6Yh/TbFZrBtWxeh3NKt1MOapxL4OlmpFeNWc8xzhUZ/7Hn3G4gJdLC9ceUve8j0IVvUrwa4d
qNGFULbsugAifRwcvPnB/H0hITFHmBq+pWk2xtcz26g/h02fkgqyLsMYW5gFULEbF3YWBT6DVJN2
ZFg3Zfy1FIUBkjQXLyHdBvJaa3ING/88JfSssw1Pn3GHxEaYj6EtLntIHluPjhgOyFAZvOpJHdaq
3Lo/SCzCHxWWMv4yHvxZBhc/79A1Vzr9pZsRiI37hBi4pmv73tmYnjxmcHFQLn/6XdpwQXy72gc7
KCs8uroA9A9+4c1fmWRBw8W1+AoB+Wo9+dG1NRY1Ya9wGQuccmi6lAJD3xcnbgTN5OUSCR7W7yQ7
i4h6j7fhqECwQ1bwDEAukHeeygwyGuxOjPTHzmp/YzFU0aOkluLHgHPeYZwuwnc+F3LlQqE24fO6
qA26vJaA2jDr5q4fRk/gXj7SgG1YyylslTk3ZSZ12xXTKB8B73x9+GEjIn4GFvT89jSew3LTdU01
FUgM7OUtw2zL29HMIVXdIWL4AOe4PSHIjZ41GmgSa28pLyJGy4GrE2e1oxAIL123Jqha6GLQfb0j
hwotepExPIyuAoebib2yhWMfG4gNdESoZCOdN+1vYhJ28tpvYu3MTeKu6dUuiZdvqlSJyu2ylwcp
7ZzsHqkCaSeZTj4rnkgLGKgBUaU5WfTbBz4AcOL57GkST2oXRPey+223ym54tcep+AQ4utcfBoLH
Ib1/Uv8QuEzXBpZRotTg81XaO544xFDR8AknOI+tsQIZBBc6m9q6/VdpYTWu0q4cnkGLl0H76fx6
2PISxp/Iq7hwZknPHb2ipCYZuAgHseOIotX6nQfDElL2D11syUf+Y5stMXxNjly83RmGpofS2KRr
MizLq90KNLD/leJLzqoIrNbYdnjYI4LgDmTJu8bJDJ7IA623SoMEcMV0OiMMn3m5NkxVggfJgl+o
rZLuq59oXFV+T+23TiKd8IQ/Jls7xugMT0CIaeoyK+J7IiREYKPmh+JLCjofDXWEHh1WXKe4u0/f
os8GS4Zko4BVZBO3IrhTvsgF9PreOWdINgJM0WpaoT+ZpOAUWdqAsH7GRa+MtNZF+7tA0oWKMUwj
xGITiigVe2RxkXLt1HL7rNav/fldZdf4GB53/BOAZ+sXo2Fc9ODvu2SYzw/mA5xfxmMcq6EDVj/4
NLZzwrp9D4UFr04qTdeP4f9BjnaxJWyu8na+9OkBJ1MzYOFlqJOnx17U6/Ys6jkAJrV0otytvLKF
t+uxHAstviP96zIkKZlQBvRJCP3WqbWKc7IbSYPF/REAodcAHnB4hnplG+/wIObgpcaYvpqPTnvH
8aTJbZotwqjQ1mhCMmbgmcayXaRJSPG/BJ8+JXhSuoHg+x3URZcP8c5qUhZEmJXSCRnL3XdIvvEe
HfkTpY3ee5xQOtUDCsGuk+9/TtmyrdRzFPm9chkvaORRWAZnpvx+sHGTV/F3UltaESTO/N3zzXNY
FcHbw590v5+zEuNXmmmZBemrkn73PjMsegUdYA/2e2FgaSMI9ugLUyks/K7FokCt9gBhhnhOLmms
a/Mq6OpoO3OoeBdOSevJc6QGpzONj1t85zyuMEluuOXbClIT39KTgQ1UorZI8lk9joHrhmw580tT
m6aEzMutEhISn7J4GkYy/5atUBk0wIjzfbLv6lnjUdL5IxPuZEHrnr+XwaQseOJiMMMZiWLQuunV
EmJkOw9Ke1HcZY0Xw1p6a11//nvq4z+S2Pzd2dte3ammoNEJO6qnA4GCEq1u0b/Xr8fbiW5S5/To
Jg4x8m/t/LOaF+vi0e3iX6DjK5ZwTVN3/voozkibFvXhw5wQrziAcVS2DlyTfA8wWYptOUiMqI+f
2HZ0SftlYvLocophJsJGjOngoVHe5lKsmMdkniUcSEqosmwPsOe+CNDIzPUVPZmqjY5pMLSk0GTy
DQwxotZUGKYKcMTzbTN5ofu3NDgRzMg77eL+dLPLq2Zkc8akTeA8OSvm8r0HvTLDH8f2Y0tODDrM
ZYYYfddC6a9H0z5+vPeM22kmDba0lVX6S54CL7htL0LIM+z0dSqHum3xlYySoqJqNm8NGl1P61Wj
mDbQqSjk0dSlr5ECyzYuyKrBnsE+3Ba5nIhSFWm4iVCvv4ma9rjl+nIDpKDUHz1NctpCQGIfbkqZ
jebv88IgoR3RuZJtPZLsk+3zZvxIo6SLRKaLr0VGHffVAwwBHkPc4Zgd9iEYjkI/wj1AYtslSXJ+
S6WZjMIswsnhUJJuUS56RFa1HSIrYUJjskVZCNdojWNleLBZ5rARXXOzXJ1fsH5ipyQy4eyqfHN2
tSKDmeMLZselUzsHKi3v+RvZZUuZ1M0ry85+u0fx+xP86N8CjW0rJjrYkD9J4hZOa16QyleIGwWd
+gau8Ib4efjlNioz8mOP8xBzUqDjoXwo6Gu43UwlmuRdfVhBpNllGjgvTGjBI2a1Ga8uYgv0dWHK
OV+DEUz0/s+mrCPTF0KhZtviBBBrpiSr3o0NPjD4pRyjWHo2y0Nfxgjss7Ul/3RxBXP7r9LfEnY/
Y+fs4qebhiszkn763vv+4qwBb0vq2FkOizWuSBLrtJOlpLlf98Z01Hbqn4e0N9s6iftjgqndrwIN
v2t3mkoKQ1GjLYJr4VYIV4DxMpYM8ncGlwEV0JBIpmTk5Oe+SmUBmScULEKX7zE6TLYJoIn5+syg
9GxFU6sNN3cWAKIQpRH7y/6LblhFSzike4HtQhWX1+4k6OK3iSY0xI29jh6TVTyv4bs7S+tZvfYI
BPnXLrY+JduSOwChZKLDuCnXfkCcKsejSQv4ygJRh6YtWrm9xIKUPiFBXL5Y227qvIAaSqXr4fhD
xqSx84F/Hy2c+b+G85BBo7PjK5gZv9J/mfEVlDn015ambrnF4D2+CMrQA78hEU5EMNNo778cQkBj
T9FVd9ZHSSV4RfhMJfjegvgWWTv+IpmXSQM/BnlU8B0pIjkKqZ6vtbFhM0q7nNeb5i6tnF+msw/C
LDJMf0TlYpWqGHm8OxbnMYn8LlT/8Idydb0Me2t7JgAaOykcPIXfy5aHVWZNZTLZ3McHCKdl/nYy
bIDatTWQsqbO0iwqPwa035lXVb8WuLdJPCJvj8e41xI/5Y/4ROioYclX0JUIoefZhSrEeUA2sln7
1UpmHWFCvyrfv2E+57ZXfuUZr+pJXD0/cwJbKyTgRlYeLuDTp88awRaSo/Z9dSxXfWn2zerqjJjm
z28WfRSq+p0W5sKB5HDRfMWaExkrsuQEcLIOefyGit/d8pq/pvsa3qG3Tq+ll/ug8Qt/hYL9hTc3
B2Cx6HzoW4WtqlZvP+jZWPP+i03gIJZyU6YFwfaPf7GKbYlTzwT0wRb2pK/tOLWttbOZRKwFRXnq
rpz8nm5h4Ow7U0yqXa7ylsXkWC5/IijJCDwetreRllaBynx4wSVIDl4Qd5/ZBD1W/2NoA8YT+Des
EUd+xtXpdFdssrMLdHP7DL/aVfbxFNZxeVzqOB9Al1UAasxJ+NeNXYkYIsg3DjyJ4p5OXqm6C9qU
Xw1u+WeXqy9BsLISXXDmLHN33lviYiCRfIb2mSliAu1/dr3hFomTueLiYlVdI+PN+9vcui3Kmp5F
YDCNvRpcqkClWOPOaenZYdts9eSN73q3rfIi4D3bsm7zI1M158Um/LxiW5VjHaUQK4LvPNnAcZcG
v18zi9ZjPCilaeXkKlUX0j8cyDP+tF4AJS3TnNKVL4I4tWSeUqDGiUFZCUVcrbJ2WSGtjLFNCz98
yTzy81KCbhbdfN61AW4h+O0cATApKMfRi8ZvdV9HPBWG8kS8CkrOYl57t0DOi+ki3OyncbBjf48a
MCqv82rn3kchvCY4I44OLRk1sY2SF1ttID1O28azVaEkaNHkwHN07YU1thV8TG9/YjhqUeg8B4In
3J8RZ4L7PLFKk5Yz76epwN1u1CO72P4wgMStxOlWPScAcEFxYQC0NiecN4aabDTUQV+Dg9Bac32s
/cxvF+CwXSTZ/WP4ASwT2sY8+aMoBjl+F8qkUpojueOAkVZKdWD8l0UST00GrQqN3G87nmjsPWdq
y1T0EZq3L2LiGkD3opcCGtvH9Awi+6EXs51ua27fpl9LrbYyOt09TCOscwyexz8XLDslsmL/ikud
b6u1awkfSmIhEPGi2pxcPyZ10TtkubESCdaYn/i6voRi/lahD4QUvagyzST7yR2til5PxjmRWGNC
hbKCwh1A/IED7w3jvFlv1E1KeAVX19a3vtCp4uNYWULeJxJol1iGcDnIUaPA8OT2yiQ0n/Z4tHhH
ZlXzO1SOKCtx5VZygnL4mwSb8s58ybCCIJw+0q5o+O6QYHGO3Vz9IRfhuoCK9/YBPIsmvQZxX0Ue
2u0TvHHkMUVwjzNRF2aYc1FF2i9tm4Z13aSXb+Rvd5nwb5tjutNB1aHwH4maYI4eCChzpzC3/OhP
Qd61xREmR4VduwHhtbGKhIFRAOok6PNd8XGuCEM73QE8TWGPWZ+isPSAmA3DRWSC41ZV0B4924Ke
9ibYLWSosQe1jbnKlPLvjuHxkhtUetr+R5HEoV7blcKflIxhNlJPgCdoegQ6L5u3FfZ1/Lcjt3h/
rlj5wzOoWv0AyU3pggohbuWZg4z8aIMWpID6lk7QGPdFDPPIbHXX8QRzEzGM58Q1uNeJLZaAcQl+
quQ//srurUXN0Q20akr4YjUxpbaW5WHQ3caO70n9ivxpNUofJItN2wd/yi2TQiOT6JECrxBhro7+
HD4IdkaSOLKetvTKHXklSqLVfg8U+2FZ0h8j9OP9G1LmbNodV1CDCAxsl4RWR4rk4hwSP0ueHyfc
0ZD7IvN92bpVMBS1n1DVwkvvpNZ81K8Zl49v1kp564yqQDrhfGUsp4ea06Ze7OZdq5D7XemJtP2a
IRBntAm3GBwu59LfA3+W+X8bP+hOttDqQNZ7WoFBTbCb88JodlxsEaf5M0RU6l1Akhiw7JU8p1Qf
nbbj9W7s3s/klGclmk4fAr8qI/BMeAUpztZxhCf8Bf4W9Y5dzlET8A2oT2yiW5qtIXUeIS3zb3rz
/fUSFCgc0dedlmCm1WwpfGsXiRjepXoZgCFFswyvDpqzXY20SRbLkcWELy43f6YzEWEf0pjCOE8R
ZACZgtz0GCJy5VqLJYcCTPYCH8bctqWOb44+oZCjJl7SQaY0quXIy5Y+aCgmycvAEyTAkfN+MqXd
+9Rdo3X91+DRU1u0Jd9gpBP8k/V98M/POXF+4CV8e2HKNK89efogPJGmH83sLp/nPtEh3YPAwySJ
9UEo333NLdlutPfmk7edzCDbFqyju6RaqUQ2KHOYMZbO7PSompdwaqR7BI6TZ2F8m6MtYfAfTKXX
gAIz4AhIrh5M0IhMdzO/qr/6Y13f+IVK3X5+JSNNT2fsCGr2bdRmCmGyMW7dmRKfqkNHtgwFboU0
NTVTTLSoCty0wPNxxdVbZX6a2tZUMEMPLYJuEN1hG5mA60nDluxbPzGoRUhcvG4Z7PXuTWYl+yjK
++Os0/sv9eGPJkS/8XvY45Hga9swENtBv3eWX8Xb4fUOB2yuAJirexiVv45t4AJlZvYLw7cuwhTg
2l0HuuaBkE6+6NqJY6HzS9nIuFIBKWesSteK2PpW592OXxTIrci6IT3bxFuY8w/ePFjeOjTvN2gO
Dxxtty9r6pFy2HHFkw5zNt+k/2DgWHciGzqhzk9/euYc99Ct2xQM0hPtnRwp3zJT2KHmBaN0AedS
ja4CdaEF5cdIW83ZMRcyhuHwwLfQgdlCW+gUmyoKLOxnT1KKRYj5b4BcSiQsW6BF+3R05i0TOEHy
Ly1sef4SsEfHwRVxfIjgbEvi7AQZPM40W0CiN0uCYkK5ChrUgLvZoEXsTmRGSPeKw8hr/InLraCF
mrffpGhsqEh2xn5JeX960hTmGQmeO/64rTJY0ATAEqtCnpzK/6ECmLv7Y86n1q1OAOd3qCJspnDv
1NG/YIfm686xDVG7gcAg/pTN4B1cCmTmaf2jsMdVZQyZQZAeOYFH4UGwOuFIlSK0ovL+YYIlCaJg
h/E/xz6OawEWpNVFVWHLkIWjpSdd0YE6IDI7NnHtf07dzh9jNtI4OMvGpkJi0VmcJLvhOC5tGUth
oUHYz8em9945pxc86oASogyklBUFUrId2U9qCNvBlHekLCTJS/A1UZsqoU44GyuSNPyUXHOaInXp
n9hT8TNjS8IfcCQONWJBNR6IZFS6yYB5eWggkjNtsvBnbQBpmm6qRSR16QJspmRW0oVneJJVOf71
qLaqHyhbCO322rRE1SjS/3nhA6V5tWefH/eJ3j/7u8LcC5HPoNrVWyOetvc8LO5b2CuL0pHuMy3s
cbzbyMc5VrQH4t6L/TN9cZj/IYxlCRspRx8iWIeKwpOlzpblS4gA3/zFo3VJBdhQuW1XQc9DV2Y1
BwmdSZJAyHv6fDoh36QCSk+rRyIZ3bDI3NPdV1aLmWqRXh9mGCQSFeAFKzInw5HLdMqy9bt6dHbc
NkTGxT3K/oQKZcjuRCN7JFAtFNOfH0MNffJGgXAUQmts6l1wcVS1PZkLCN6HD/gEIVZia9ghbkPx
lp7d2z7pAtoFTOhq6Ho1kLuK9e1CMl16585c+kC8gK3RJaOvPj5rVs8mT03KBwvdlUz9fdNi0Jg3
/cYf8ds8mwUQuDIsdYVzBByDw0nLJsu0sSL6z8f498rNTBqphW51lJoAyf63cc5vfT0cvt+4dvgo
WBe3MoWT+44JXSwOOsBZ/HFUwsPiHFBirW7K5caoRUKPGslVwMiHSlT2z9SyCj06dJped4VeaVxl
o6DMs18shqi037mHG4I416d7DX31/S8hp1ZQvsfToFIT/j/Igb7ViY+qaMxPm2bsl7uK2yoRCCa/
iisp/yEP9OOi51u9YXCz28h9tgJrAUH73RZv58UpmwhwPgAdi9RTUEVM7fe2vhAGYlkNuU+mY1dC
il9VmH6kiPw/xm6FxKCfE7x08mLldCegOZUMrvq2eZpJoIUNUfVUfzKFHW5PpONXgg9WBBS4tlxm
1/AEEnfWcN5m4AZYwr/MLge8ONvi2jZtg2c8Zymh/kcDPS7qAYjm/qEscY9UMIdE8zqezHd3hI5p
eoeCk9crUPz5W8n26YlM2qMOC8NdvtrS4FichuyVNsivwH5ld3OljkC5Y83S1EVPE63+PopkeaZ7
4+NCvvN3XDkpaKAZVxJoLqkQEXl5fQjvjJpTAeRc4rvmHKxVxv3djLYMwNxlrYuEcmtQKoFORYU3
ULWZOarUD3akdm3lljDGfPBjNoVZMe9krZA6+Zhqncz2cxuetxPGciq2aps5sOZPMyFXdFywdmy9
SFrtbGZ3CtloWBaVxYjlv7OpORzhPTlxrt1+CpoE4yj9ByH/U2Pe6Syjyw7OBMIg2bn+GAYblB6a
7JANiiqH1/LbSzMLDvYHwPHdUbNuhdpAFZxJ0i0uMEAGpvLV77/qjj8BUOW96rkikEJsZhNQBu5Q
elsACZjamNbSxbDJKMUxYO0vORpvP2GxhKHUZO/aJYEF6nY5pgpCfXptBLAO4HdXkxITNGoGMITw
hI1WPJ6oePxItE4Rf4IkNNCVPkY7i0c9BpKN6iIvOu49DT1XPg9twQqgtxIAkJ5oy+UK3YOTWp6Z
sl8Y+cUAiuucWatbeCGU5BcrhXuXayo0p77BFPCVDSL57JL3XzUdCT6rJebFwGSOX8wXfqRO6gbx
UufatBHplUn6TB+zJxE8aU/6jYSG4xKpcK+xdvhIUbPhGVclyMqjKaz4DGjxT8FMiG/YulYWk+WK
9txED7WKXmHzOaoEiL957hr27kgTfocZOtaFg84Vw8hEkiMlppmRTjjkUJYxDOZWy0/1DDHI2J57
j3UnFLHrMZcbjEtgNujRnMfJcuFuAXvo+FDw/5z0sFkj0cIxofxREYGVZPkLmVlPE2/01nvuPlyt
TAefQz4oasE1JWKD2MywUkzkGfATI78XMiQ5+5KCdg8zqlWyP32pr4h29Ub8kU64ea2R+R/dgaXI
xNwvvgSX53l4/U6rsVJn7XnUvkkA+WZmByUT2tM7SWIwLw0/2BTmS5cZhcHiCbv7q9WT0JFsU/aa
eKYVY8s9EkU/dDmn09qUiwOjtHzYFB0WS2VFTMZpuVhcRqRTqYxlq4KJCxS5E+VDmfGkd+AZ8UB2
S1Fly9nUuTU463gKg1WtSjzWRlzSANR6fcywrcm62pIQiniZUyrbG48U5LM5oQjJb5sUcjsIG+ql
a4Q/YG1oLHN1gUAY/FVH1GWKXS86Or9c1NFQssxnp8p3KYD2sPlrwYdj8luIpK+9rlfwBsyrclhW
knjFBQvwKXNJMzwDaLgyvxfi0JkodflFCzD6ffvxrQokitto5cnJ7Z81hjqHPCrLh5jg0SS/B65W
v4VBXONLkFPujLeHbVVdoNd8QvHX4Z9ZdVl0bSyskfuU8OJE3hqqrWgHLEt6CpKEtkHHkQ/iy9BY
1VJhHZofQJp6y7fA43BFunMlca8ZY3R0oNrXFksUqaOwKk4DQkqqAOMJ3jwno4h1kbBvw4hsyAKz
1BpRZXlSK93mblSmjmnDu2QnIVFIiNNmeJc/oBqqBF2xV4bQxOPDgJm7xTB76quSAtpdm5QGcXe9
eF4diW9R3mFgb9MdNpeSJRsShE5u3zb8ojEFMSDUKxUxbgT8jhDGj/s2a6NibNnJQOQ8joVPJ+JK
WyxEooOiKFEZ4f27cTPthzPqC7SbNKgmxBCcPez4k+EfSMuYLYDXYUzmfOiK5ZLfPLVIU3LfObg0
gzcTKYUMzmnssbnbXwvkD0YmrAql7e6+BQQFiRugm7U0ENxy/BUkOr9oDVe/QGikKWxvIO2tAC6u
XSUrIJQ1rAunMkW7XH2Gws/AlTTY0q6o+UIa+qIcbskFneVELtEV4Fp+c8zO0/E61/qg0UvpXcRw
nfNpBSArGsPOhAlodqhQzHQNEGQ68a1tbxx/+tPmxBD1sFd9KP0SpOKwiz60Ulbrm0LuxYZYR0qz
o61OPIAtbmoyia7Jh8dKZDdK9wW8CjiBd5BoTR87IB5vNuIB6/QVcIKpn4u8ChC4ofZzqd4O0yXy
2JTG4kQalFtxwD7fPY66zyv2NdQ12UfUE1T0RzqNrkKtGHCJCp0MFDXXjTcyB/igp7ruoCfhJZs6
tKMrglMVR+MAo7YPzb9JMXqCrCsgBAUjBeWaOjDeXDFqksQ3zufzB5YQzucRuXOTAnMZQrsGK91h
qtYeteruJbKpwmM1m22pd807DmLDMfuTbdbp5aDtCi3ym+8ut2k1ePVguRzr3USmSYMO2sGEhhOJ
i+RAduhqeCwzs8xrvZYJtF+Kv5xEB3PR2R60RFIigyibfextafgJk1/KmUdIFoEJmnXaiBFWd0yR
9I+z4FPHlKN7KQlwlbO63+9/9b6NGOZ5qGCREHCNbLwUTTKcg46xpRtKMh24xq8N12S+VqvAQU4s
I5BLYc8oDHON6zpZKM4EbR0iTYO+9TmIEhNzqXcZrb9DAQcGofMDm/hDpYaUUh/4M25WhnO9vAGL
/r8XWOgw8OND3cq5uZ2v4xGFWsgPa5p1Vs8WIu8KfcdqD/aj+fssDUwc7spuC+6+bv4eQAAJjgV4
+oGP+mWCEKit0aLN/k2c9s/ty2uBfCBNTU0X84bvlJQYlnnDw++G7uj0kbjygLNJYbGdFPGiOBrr
JlUbjhO8b8RNfry1bpg6h9SzDlC5ptVlmwpZatxEjhbuGWSub/weXHZ3TZaRDzp15FOv3mW3Jym3
sO8YhqSHHX7oP15PsqfVF3CqdSaKyzdEfMY7FH1Jl897ezg9HAGYAfvAp79qRXY3WJ4rSeyWqbbg
jJ8QJLuEhOx6vMzIMNIQYTAm8Sb+Nnrq00pnKF8Vrd+EFfkTKvJ+Ar93wTDdJnonCjPaWlp/aRDq
4f2IC9fjSwfKtSMN4WLq9H0dYwfFzGHx2qcuChHcuPMEx1ddTgL1rQ/r9vMZrKVcyuMFD5VdwYxt
0tc6eHbWARJH0rpg7Gw318JBJ1Ii1FVwkD29vv1v7GyPNgPZ+QmwrsKi5J05HZDlzr8veRO9Ubwg
998gRoC+8oxQYEjCSYcKLunO1JPK2Qlq/Smzzx/j/zWaGAjQyvT+tKtpZHzgOgL0KxkddUsfS2RQ
4C6z6FX9l8meqOIjM8/aP71OM9sDwujTo0WIROvWGMxn74drRIRPDHs/YfmgRWLKs4J7mCxRSQJZ
x6HhdmIA4qvxpvyOarYXcLyUdtbdP6UiS2QjNponItsz+MzhHwsD7HCmujVyEDdhRwcZEgOeKdZ5
/8IZkckHITw6Qou3x5VO0hT6WON19CMnmnsSAQcj6/a1AlNH0sLkNW0EUyXCI6pPsv06SlTGos87
93iRDx12+vzWjSHVbeKXq46Ap7LuVKgNYRaf3neurf/CsuRcoz5Nv/scd503pWic3bP5Wfgo7uCS
/CHC38sN0thmAigPEe+tNLQbAxeMlkhu+V9F3hFSRNgMJVsjvGqi3eYp/WZ8CmWr0uEL9ySchCnu
2H2Cd1i0RN3UkSkuLDBh0SJuJXisvJnnIm39uHASVyGepc/N8TXJHJWUFXGruYYSAu0V3hHR0Cmt
BMQEU2wjX6pW/0BHKP9KxaIKbosqVzuGtVu0HetahpDOe0qJd5D+aPeIH2SPQXdTtzGRt9xoTlAV
iAT509smJu+SuIVy8zgBQoqiuIPgukfcmbOY0F197dF101SXh373GGaIeC5xGXt1c3a7EpupU5Q2
qCZLo1Z/WIeRJe6yYfQuYVIjgxP7CnnpFKTLWs1jej71xym6/BwcTJF4YBxoZfmisZjiSmGRjSYU
75qIpezfObsHUoL5IYwwAWf3Ay65dsbWqd7z56hSzPW/gUJafqxhKb0pQkCekfJ5BGyfGbNH9ct4
62BAH1frYLh4b6UgOa5b5D0jXah1jusEQROoL035aHZh4mVxpv+s2bfaT4hiw6Yljie52XgPq5jP
6ms3ioA+QM1+MHwoLdVmJnIWp5kdhfVjOuu0dysj26QCXc5KEpB8AqlJHMnssfnLE1u8qjpNZZyF
OWooR/SGbIK5US1m1S6PsAbBQ9ITrUdyiiLIMXve0/C1ac3fRRIhZNcWJbO6+n+8qG5Oddt69Tzx
jyKVDXSEY01BwWMyYWNVMijY/5nxlFHX2dVwbL5EjGNeT89LlYpgdE4UIOI48hR5MHRdz5893ie3
GTZaEviA1jaRg/XHtGZ5UzeW+j5bzjrs/aAOh0jnlicidTakKGCo+BTD1ZutIn5ckR3UirbChhh5
c6MH3FavU4eRCeEL9PaPZyoos8NG9AQqWmQGVWLY4fBMEGCiQo/pekKG06by3GQeAS6c+dCdTCic
AOJEd9+nrSjYw9ezaXXp12nJyCJ9OmfC6aaQGvPmMy/nI+nz0CfYye4DUoz9Duk0QyoVpLvQYQUn
WRSuQqYGl3B+s/RXLnE2Rke1oTI6kf4B8/kxtyFwJoCijZsbu+O/LvCHmaw1QzFcEIvmDMb3Nado
gvhefQnFZ1vz0Zm64JeC/Zjr28QwfVznVpz5q9kWcoJ1XAr3Hjf+TpZOLtsnXpECskheG/V95yn3
WmQi/PmX1sYONTxMGBrOj0FvFmLInQom8N+dIE8nkKM/jVz2B7gv4rUB/1jgWDl97jxd/u+tb/JZ
qF7Lgv5owZt5PVNOgCNZ1gqTSFbPxQBBHo03WQ9z8un72yhco8UNeYsEBvlIsHbqGrwKr2K5X1Xn
1AnAPqYd+K1dRE3k7BYpYI5kpJSgrpDVDgbWhSP/Jb2Lez9yys99DdTkAhVwClEd6MpG9jl0zdXt
BvW8MASwYTJ32b+PYcKem9JrbZ3XnMz8hQiQVUK2EI9/p9TfVTXPMLWITNe39SCiuonvxhASJnI4
7iiswCynapprhLPcrzKw/SgeHpZK5DiKSxO2Hn6v0DttxFHhebUADafoqUguKBGkhKYSD+epShle
mHFcSO8POPtjRW19LQ5JLG7nXQsy4IVPYz7OdAbGh5S+GcnemJyMRgmwzzUC3z9Ev0SxqGUuIebX
Zy+fRu8+dVry/8zkZLkArnog25Z6fPgrev4M04bq5KFGKbxEnHVGiDapYjtIYdlzjM9El8Y/bJOY
0x6SuuPIVlNwl1x88R7xYZ8iYDrFHQXD+WK5i7X5Njl14OBEFMzRDimkFSoCj1FZ2vE3bTIalLpA
N7viO+h/WLDq2OUwp2KcYRuCeKlLxZD27oo+FOeGC9mrMXXiSW1svky6bD1McFzmwXkhU3hu7VJ8
DCNbKp9BkTUC0dPS6TEGFut8/1gJup3y2VDx/opcPUy2OinUnGJMboJ92jyI6X6qel8T7B+ZwYtp
im2kJgpgb0ESy8nCA7IIqqECWK/fQPgBgFuhGYq97xZBQJJy6KVIwSElinfI944uK947urLb9Gb0
t/rkOSe/vBCYu6pccG9TPYq7MP1A16QY+nEp5oxERn8neqYOavsSYEmbtLodFBLMWKEq5Fipi+w7
GW69n7pRP+inxOXpnrLLzSn7Rjpy6gmTFQPy+CCqqIWllktb7YHe9lQ65oFbLe2oMwBgSMCPEgtm
lVjoIKjf6TaSt06zSf7WNBBW9umrvdlr/RKmFCpiUosm4VBAIlPI4KwERM+umWwLxPYkPG53MREd
YzXj/fgYsOg+fBiwUJVf9ungEA41NMJNDS6YJTb1bKfiVPCUliOY4h+gKo6rqQpum6Dfkuruk9A3
CI/kw3HEw2KZAP/g7SVFhmloCtXUYIvbouUDxz9KP/HTRw6dHDkaPoYdQPkPjcAMK26tasWD05NG
H/QHbJm89YaT7uX4QqkIUv3vY9IoUzgyDGQivOEXHjSkcXv783/hHNKGV9GGHm7ug+D9Je+vVq2I
d9DiaptqPOKY9d9jC61ExpvRiNZd67LaKhGcA4gqR0gp16Oe/d7XLC622iQ5ZcvEP4J4Lb1gzQKk
Ovv6mjd1nQM88vyxpiMNIDiIE2uKJeq9l7iWPUIPngQKay5XUYAD1R83kHhHuvpN+L77H0RSH6tI
BZZY4kekZZhHH/DDdFuLvmTPwLmk7/31/l9nhSGRa2qrtkUW3QiSdQfHqMlTYi/WC5xhUV3MlNyU
5TgsHyuDpV36rkloMoanylo+pFtWzW5ActxA+L1DzRy1Gak1ydjQhIPAftl/mNjRg65SziK8QwLt
ob1D4h0Q0VmAyoj05B7jbyvO1OdHoiZogLPZpiZ7HdhE5Sup0BjV2ntQk5rttf/wtDy/fUBzmaJI
kfOPjOJ0FA8hMrSuanhNbCawjzkDPVr8rI0CYJpxlhYwxARmsC5Mk63wse1a5m/J1MNCzwTJnMBq
jz4f9zilp/gO8PMAy9zlUZXvPUOAhjzrUT/banhYExMYCI261j7JK6GN2k6oLa3fy4in+X2XR8C8
i4OQ1GzDmh7ybhBxPzimKlW7R603kq1DA99GddMuVXAxKOorAbQ1d3DCXS4xs6/4rmEz5CZwzmCd
UHKww1sXcbHYv8i0zGZ5qDlM061rzc452OKoNk1FmyOZyAnacDVmbKewyQC+Mggp0wMs/H8OtgDD
ZaXabl7YHgtTv0vavAqzb7lxuz3i7y+9iqRyiQ6ZBNZFw3hnF7wJocxqZBYsBVvK/z+ft+pIugFq
VqewRTdQShFqtpdsKjroO0vRQntS1ca7oAsre2A14CBPBW61Ij5lnF5Wm2YVF2+ovTEo2Kv69a4l
0IWV0MgQP1bmxqolhAlX9n5ly2qasGgaBmXxcPhlmifb+kKl4nfJuVmUWGGNjUb7DYCC58dR56jO
CZvdqXpyDMOcu7A4oO57TevMNpZipLMfkbKu3Ez428/tAt87lxW0AzHqd+gdhfnkww24i01XlyV/
EMG/IriDI5733ta8va/lozq2iIRON/V5ssipGT4GTd4N1Qt0hFQw2nkXU6PZUpsFhbEy7xGDcPyZ
o5tockBXrZEsG7UqsWupRxLPS/XRZ1mmeKZfDKEL25pxJMZK8qqXHZOBLatm5nKUa8yaCwutsNb7
C4DB/HmfL0wkBZeLbkuGw/eyFaNpgefmk6z5hD38tVv1gF5tAfTuIDPYUAzXtHhnJMbcIyOUnnQA
BQlrxlh2fJakGjDVJNCkG/QZAI5y3Oi03LWlrsFGulzzCC6gFmyG2ykdFKbo1hC0X6gimFrfajMJ
bYyqcV9Ez1HQQC45hg14q/Ubld52oCymhITXS1ajlcgHSA9fDg8VXophJmde2Hi+A91+HOUpHrhQ
c5mPP1s+uqozbdJSLl9GFHIwW6z2oQ8xe1numJXj/+bSVRcA0EzGYVb8Va2FFEXHhDOkYFiZlL5T
gRG7auJGtCAWPr5nUUN9+XEADhS5DfHy2PxRhHOpNvcZFaX584Qi2ongqrmR41sfhvJGKjeHO6d9
GL8fFbXPkCYZa9dRARSXRYV5X0e447RsJFd/0m05MZ0yZrW/R+U/dAdrCCbou0ZORLTHA0TL3zti
lOeIWdMeyJyvPSlpCfaHtloNpPDGTJwjqz0NJdjXG00p5yxtwtcbRg/SZ6UAwAEbo1mgKOaIrdwT
TlmidV8vfpyC7I4eu75Ps7gyLWTphY3v5jB5alLxcwrwOS492gENqzFw/ny5mlencYIWMXF3iKTq
tUtlt9ooWVaZQBHQMQSh5pBFFB/bYArxZ8b1M5ocPqz6gJQocESILQw4znHoNu6DwnibHNMk5tIe
aoISxqtEYfZjmQC8LIUSng2k9snMshgSwxRQEewWioEgwSGGUPuXMzIBEe+DjCX4cJyGPvOCZRwc
07p0xCrbn6uyNAlQBhj5geBLKt+wvYvxfsAgwn1ZIgbuWzwrDCHxpzG4DSg6GAFbLcXs9h3128Cv
kThf+m4IjmoLV4/SOfBAzWABk7rQNBL8EkDtIKxVOYW9mFepSNEOsoY4VfmrQbJc16Ji5X5faL2E
oxIZRUNLu9LmXMQHGVv+joYPp8PhTCn0HbEXOLPDk4OnYkJmA7IACLXib63uaR89Z1wrtqpWc0vj
giWdOMERe5YblcYKi0FUK1fC7I+mHbBvOAMGFeynyO4/BnBDmhdyWiG+Ve4CS8njCS+BgX5lz3AQ
8DJFLJuVOlDz+IVwiqj02t4SNZToGHz520xI0L0gj86Av68SMsUYgnWc4vb9VDN6DNUSdNQF7pfg
GmxLT1rHVg2f6cI5xbhaXd83KnRfkA7iLZSeWnu8T9i+ddsP+cdCD1a44jaUWdMht1DCceXE/Cp0
ed9L0wKOCKlDhakKJXImLqRpOgoCCwT7lZNYBMCOsEU3J1G14mF8w83C3xe2rQWOkVZm8t1VwC+k
fGI/Tva3cxPhb60NtOJkAb/JZQfJXEqwjScIp240YNfa6BrG4oYskI2lHqEPTE+4wkCLRnHgbVi2
gwzDACIZBvJDB3ep5zcIpv6Gb0RFV4xhRjKZAD8yKnW6OncfsGhYzXlqH948n2c+UhY190IvEg5t
e18b+TFfx3cdRHeJEk+pdXcycQBqLvyV/mxGsP+DhdafdstWDPdyiOrUKf+Gau/1FoXSxyIJ41wa
zAdDOtzsV2RTt1mDhaNAdjEuc7DBMrfYM372d/hg4SKp9GFmgH2FDybYMSah2vr7I7SimXmJD3BV
1d2DUq3nl27A7xPXrH7dsXq2chQDHw83Y7naXVoux9P6kqO8htuR//+iYPPmtNf/rHTH1pYO2p5F
TuJLUNwyLRbH8kz4oqo9ClYoyKjv6DwhtVLFVRz+kjEGZYJ9t7lds7Ot5j/ucbMJEF8o2PBjcVOY
7McvW+Ame4F+hwrCiTvaenk3L5mpeLoAR083ffywh0vGZXaGT36aIpFMqv+wBnXmCH2QsNQYR3nG
knARw+c10MQhcamnxolKyqpVPBWpPsOKIj5c3NPY6FYSlGJffoWfkL5YRU7t1i/56dr7qrkfoV1x
haZlPhPL83v5BzDRhpYyM1+LFDov1rCrxHWxlrhDPtP7jn8fNMsV28u7xZHR1kAG70qNnkv4wQ/q
+uwkbwfaxrHMaT071jMg6oya0F+snsGkCZ+3ZESRZgONV02qz6s/PqdqSZES82bLXSU454h9cUhn
FO4UR5hR3+qmSOESDI9oUZHqvTlhcbH/51FUtbedNd0Cld7JrYcX7SSC2c7m4ysgkhHyFfBT8Zym
MTcH36lam/VIIfuO32uryulDvF9UInbod42dhdeseRW9AdFKSbDGwz2zpPs9h+xsEWir1sOv8Djt
Gm1ZFNU/gNI4LgO2vV6pRpgw6nFkDJNph1tfHTPnzhTKKB9hqR3qAWZ+ForFEdX92jFkptI7A9sH
NHl2VfvqUQfsn8PKT/1H0UQvF7z/0k9AE2Dv81VkPDGTwXXdIFckgKdxypeV63v3vKpt+2+IP39g
gXGiw9HDfyKXCvjRJ0PRDifw3rtP/4kWB5UDJxxqV9iInRiAm3Bhw6iESAZfuSFE2+hGVqJl5S6S
mJhg0W6Ho27+blPyfILcrGA5N+kZ24FkBT7JZQTbYyL+GVRKZMxDD2Y6/D3Ue0KUmZVy+yBymzYA
+wfRW/hGkF3NX6lR0V4ZzPdwQ6gI0xSo05ZYMYifcr5ZWTKrO1MUaDTEdD7oYaP53/E5AUWpexQG
+5nRXNkuh5Th5x8yqOvPPt5B28VNAI2soxrz7b1CtqP5Mc8Jhn/vjEBmK5ejfw+rH9rqaHGGdPtE
EHATUOf1i3yQEk9dTToIrnYg9knyvIEg69vohRz6+4ekra6fBveHmQfZqDuABm4MjD+2+0ZoGuYN
89qA3hOh2Cs/mHnKadnoBN00X8F0b63i1cWGhezoNyXtu7VULqTOvn4kIb9rXjSZlfhyicYWY+sC
0cp+TcwwUSs/q+MSAb/rgEyUbkoTbuSWSHylBTp6bK+PAefkKVFW5J5Z+xIO0LcktYy198XKD/xB
5GpNf8T9+Y5fbpJxnLNHQKPrgqE8nmCMUJD0JuzPlUzNN6xoJZR7r7UejDTLfaL+i5L/7AkaGulO
+IOSM/eQmQ3gR4Lec369oOhH0sy8gtyjCb+LpgEWpxtQKPc0iw/5eFSzkxarxSYqKXU2doWnMoic
IAtBB6y3fvEBHT4U72sA9ett4WbzlM+yTIylGfKVsn9qmZymTJ3bNhMLAikyWhP8LTYC7kP+QpWW
e2dxxFf4Zsv6WCvdlawa3iDzUsJAgRYstZAlUM3KrA57SURQUzHqJDuwdiTnxGLy4yLMoCvbVXbG
1F3PCz2o7AIgEbIYApPVqgyf3PuC9N6ndkESg7VKYcwqBFJ+j7WHy+uzemdH2ZOGpeEruSQ1GveZ
3VuyYELcQbPP05x0oA7JJB5x7xOHlhX4XjJJI+rFoL0lIl3bka/G/O0hbmW7fV7hNQWpCigetl6i
zPJuQ+rLfboY5p3NdK/aU0So3TdftGAoIEOyomygfuZtgmj0uP6gCOcjQoBS31krPsyehFAAP7aP
LvYm+aUqhar7XnwK28cs6E2Mq6wCF1SVkuJXjNvG6rqk0gNMyZz5alY1AOZTwDCe4ESc8I9uckUk
/EuorqKrOaMCJ+CH9KeG4nQZRv5hQ6DLXqeL96HbNawCgDt4kge0XtN+7xgTbDY63TxVodQNtasP
WyNszxjnAv82D0mUipGcOgl3wzpZclKGqkhlvcXmvpoJO1h8nAOiAvQVOH4tnHrFhxg2QWjvFJqR
XzblAFPR6mDcBgmHkKlbK0mJRewckRD5DrWiRdG0DLbfMP48uwVBSQpaEwemr7qr6/XRnXb8o1AQ
7VQcTwyAM9Hl61WIPrkgp2J/N9FJFma40nWd+xr+eIh2DLNMVFT+jL9lolGlFCtr7xW1YXdhrKNT
5nNN4GxTGlqVgKOXBE29/a380Az4GH8JYOGiLLCu3u5q2JGzfP3AJdjsT9nxRIZYzV1LJSUMtiQH
mw3ZYxhlfRpGbJWnSh7Ut3nMEXZkfHJGh5fKST+oLsPWIOkKROP1bwKvZDXEIIwRnZNK5oyo6+ex
fHiDVKjz0bCmmvjIsWo+uSonowwVeNjEjR0Py9e+rjWQRc8uDBsmGGwnT8+e9W2khj8llUBuNzGE
oNML7YdPINpc0vKZYOsQ9YQpjihQcj8DRuDQCJxELcieElTVLjekAJGYA7MYufti0VS6uWY8xHRp
haD7mFJyMomM9jGV/P0jjtjhUznX0oSfizC+7q4tRTpoOPFDsGbKW3fpcsrYhH3JBAWLucSYh9Rq
yadYot+4z7IQz+yf7mj5ec3pmbFAsOCpJxhf4Zki75x0AeudxDa4K+E3LrS4tdEFZhtPqbnV2ZDM
Ux1O4LOSW57CBbPT9BNSGNFWsY0EXyEDBF/xm8uLEdy6UiKgbN5qPzaddPI32isGSC8ilpnuFC6m
aejj+Kv1uNPOovSfj9jrYQIknnsdJva2YKe+85RmpDX5WwGAr1SyRQfP12vXYRLhun5UwbDDBEOo
eSKrkua9xjDbZT+o5glUtaCyLSkCvEEf4vgdMAtWIynwkRFQx5K7THIZo+VW7QYMBUStN8SFiSOl
n0F1gbd5jnfEX36RU4TF9QwdJOxbC3WLRihmosBQfeAFA9PcG7ZqxtlJ6Dfq9Cozw5RlSvAmtlx4
pLE8wS0u9Kp2bafjFUMXPvQPkoTPRCND7f5/JgObKpQ+j6Iv1bEdA0PWtZE+ByNVeJjHx/5ITOAx
Unk6Avsfr7z6hW6jfGd76h+BrIojCAnh36MG1x0bTn4+fbOXXIaKsTSerfbzszUO89nYghRa3krk
ioUEmFVA4uT9+Rf+YP+3E7FAP/bVy1e+ILwq3my46AJVu0ZrBHSVOsZllq6aylkFrUfSjUzJG/z1
ot2tI+1pIfkSR1X9ZmhmV0dFWLBQk8e6N7EcNGf+mRSO3LVyd56dvWdVInu83AuJn6cQ9Y7RXkDT
smYKGE4MqJ4B32p/qZWJSryztplNK10k0LZWqIsju55YGBU69hU5E2UfXDqfnDPjvg+kCt1fGwOb
N5AP0xmxEdWOzO4CxqgEt2p9V8kKeZkuQ/prh9r0wIJZ8SKhCtjApr3pjfcerNKOCJfq++26pD4T
qD31cvCnCY7Eoy8ImiJizNgry+f0sm3MOs7BsxGMTY+38XxLIaW8GYQF8NWlJ0uSpOPFiMAUqpwR
ARi/q9fTB/yyYUEpxdEc/JtpUhintYaCZR/Ca5d1aHJUcbsyAQnYkTUzZY4+oNkbK5C4LDc1w2fd
O5wlADEUC+gcnw/nHZ5q2Ttxa/4Q/6x+hlug5ybUDP+8mtXp5YaUxcCT/MMI7C5ofmWdrzOhEVYK
bvOjz8LbntyIGySa1+GPJSb5Yb3NHrEgOkNtEPXZDdkzrMkenRjxAQDVSjBddfVlBYSk3Kd0BY07
/PfdQJz628f4t29oz38UHXifRqyElkVeoxfZ6N/1kH1TsUuCGbEbi/ZHd4hsREdTwUhXYpjtengO
yCAXP5vbeAnyJjWOUXgrOdYWEPlOW5Yhc75p5rpg3UiS28imCgR1a5ZcLPL+jYnxqZbLj33i3Qp/
gJpHvh5uBmEYwTuzwRckTxt17LJlDCrrT2yLpIfjq7BHtg2oWQ3uvLJfSVE4C79BJKpx0FsNxbkr
qvtnK4cvO3vs9qP/v7SIYG1hS+BjLM+fEmGqYM8x3BdEn0spGWj+x5gTNIXqYN6PI12acdj7mS7e
MznYidJGDIVYM61+PhwCN1Jj/LfaIaORiPatx1HVI0fLMgGU67zCkzQrgda4Fbw5fgBS5eb/N+rI
X0EFZ20Gmc+PQkV+QJDnVmqaMl0iX0S3RsKqWMBBewHY2hjh/C/76EHxtc18fQ0MB/yrjnky95Q8
NY+En5+o6CrHjnSUNFjNNVCoxMjP6TVMLDq9Z1K3sbzjfrcKp6lQCK2+a2a6fIZFEfZD7NPE/AeO
u5/xXoubtxgbpfOZutxKGXwL5clZgu2Uqi3+dn4xNWAGRBMZFP24rB7uHVko3SsAuNIv0jdGTlww
fpHd992+Adg8UKXKsW2eQAqitIIJVUDkxnh34kIixpDta9Cxt+kQZdP3cUyNe1iHyY+fSueWXtvt
2g/4bLpT+1I7FQjXPXiCLSfK5VWEa+dB3bS1ilaNIoE7Nm3FG3hOcK4JhbOIcCSMJ0ZhDaEMHrbu
cbhaRgnYKMhp6XIW7d6OIyt4mWk67B7YgdgWWfG1FNdPKIBw6vSY4l+kUio0Es+GWi2q327mQ282
0iSN+ico1oIXBDu6x9yQdQswcpWI8XYNf7xPCfRx348/zzXiVu1tz8CRGsCf7qmP8NZpCGhbyes2
3sk3WP7IdigQXU6J9d8LWjHzpR4kvPK5fw9iZTLDabRDjFXhgvV7JbPXIa7xBvtFjG6L+brh6dRB
hDua10ykXVxLvKP/rMUCHSLXFap5niKKi0mvl33MY9U6Xb/EDgEhXTTvYOaJA04f0Md0JiFFpuFG
UOqe9y+1Mn8uBvn/SVQ5clVffHw0Mukpw+7avhscbGkfWTWWnh4M/Kv9OXKkijm47bjAXCWMs2fQ
/A4pbcVsynpPjhRPYV2KEXW9srnsLjPfnp2Gvn8W1RXWkwMF6Dexvl/Jj8BiPwPvzOSAwmisiuZP
E90DXvtqGagSscJ9hV3EI8LRJbELyZ5BiO/gxpv+kBVcQHBIqyeihq2YJFa4S4dMpwgYv6mYCi/4
u+/8L5RiNrCO9PbVOuVu194TRdhn8LWQerH8jBx6to7y1H8/96QVQF0zkY98QJrcL7jPzHUu9L28
TfpiZVzPQw1+wEdvpeoY+l4wKxyFG6Jb8KDIXiUHgHXWc5fMUc3hCRS+mMGKXeup/5j9HssfR8dP
MA3auzgOZZtkEnKRCuSvrjNeczR8UYLVOX/JLcRCAnklJgepuuAnT6MsCzkEt2nkufrMKeKwjnUQ
Ez+eUrUKQUsKBp4HB3PO2WUAgkAw0RensWSLTwEQdEncxgHmG0VJ2fMQsT9R3JRhaXi1QKTSqkrA
hbDCgtg4vME6i43xqdepGx8HJhgpcXICQhAVQQK/uBavjWFx0wP5EsHCbKRmAPelFT9bDubpO8LF
fpA8heJ13+0IJ56RCGfeLgvCffvO9Uvu7d/iolAWndx6OdFVit8Sy3r7yIRcCQYOJx7aAkqoYLvX
NGbF9OsgrUcojz0rkxlnvt0WFLxIaixNbJP3S5K1m8vXu5m+oLtRUn6knzP+G/uB7GpGp9rXcanu
MxhIgxKcWW9xLNWHzr1ffs/eLSabjIsVDsh52cGOy68GL8ddWslK4dul9dZ9DZCUqb37ayGE2uvY
DvUpA5Ogmg6ddcrb8BO/JtpVgUz/psO5bYHoXlFTXZMPesxE6UdspLt7djBYzwAzT/llCXJ4J7q9
8LKKQE+jk9rGoD5yMX2+7zDdjC1TDhLibIRV71OohZCLGyb7WcoN0q5BOQSWz+77bh6YXAOvwEc8
HKCFR1TIYSABD5XfQZcBoxhWZR+qiNPr/OJG5lF5n7PlGSOGf/CbPKWUDHk2gHt5Cao1L9+FSDDf
so9gYTDg8xHtv3gWtzexAWfXlfNsQ9yzhmv33MKUyEbkvYUxxatf4/C/O/FWzNSFpwNZSpfQrYNe
SqtnFnHWrHK3muAxi6e8VGoHkWnFPWRx4OW2PoZ+owVugk/5VhXSyxnmIJ+M6UHWvUx+gHlpJSGE
9v4VsFReMK2eVxaavJ1BHQpjK6i7HhIqsftc5K33l3nfoR7HYJG44/yXkPu8ni8mOeg4ruDKE5Vw
4lYhp2844Pf4RcalnmCv9bsoW7GBXrJS4XG+LTCflRLI4DCWjWHAynPvs/kdnmxMeIIUguJLomCX
WkmJhD4Bhh40m9HlRSy9Jhf6yGAtrJ5lUzT6CBEnIaoDWt0fYfpc1kKfOsthnLLx03voAetlCa0Q
638xvEf6Hnxt/gXW/wXw07fOB2tyqWUk7clO6h3zAAwMwSGWG/Q8s4grsG0u+vAg9Nr/dccbDBxF
n5JGPcSeeNOUsprwWzMg8RjvfQ31mJV0vn8d8sefr+9/hJd9JbrKbSRlPVoYPZz/BJR51NBDUUPj
fR/jb7etBzBTF0RWIGX3s5soxG4cdcX9tevbaxtM1HyYGXHKVxDej04fOJ6JhVMhxYmQXMNs0N3z
H7C+G0k0pivvwueiWheR8j0nAvMeGFVqGPpR3tQTWJGA8kSbIQ6mneSSYC74zCAIWol1PAd/wbfu
4hCatOKo18QrpiYg9pONgzVeKno4mKcaXiPde26fSve8SWII2brHuVo9flSIzk+b/Vl/H4X46XxR
0XYVv/Ng1KVVJv/TtrxL9mpnOhaRrC3/ryjxWUhRiC21cyuMZ0iP1vAptWq1hem6MZclXnelDPMO
8tbQU/r96UJ9hpeVwWbBPvvcCCcEEEfLxc+7/uzuiabS5/+7X1loYwg3W6h+yWmfFQr3nsbyayQk
biaDcyAPNT6A4g4m/LaMAcqLWaNkXWOaZDodibhq3UdzMlocGSM48iuszHtMr7pfBTVYO4zOh856
Oby/xsdwE6ef92T5jo+Y2PHW32xIIFKWRc+c3nG90nYOsy98w35f0aDameK4OxpjnXujiEOAK4ow
K/F6P6IDkb/v4t+d0jR6xPQDDAJbUgkXtuf6yhJPBGWlZTNYj1K/Bd0bREGHr1Q5Cvxf/DXhXJRY
Y8qq2qPfv9+48Cg1tH0CR0tMQCAzM0AAJsvYTTKm2lW7hdUWVZcpPgYBoIHowkJ1pdTFV93FhTdL
r7b6C83rSL4GvyNY40Z3ZruVvNs/rc61BxwJhzqaeC5jaux146cf3R68NWRW87VxrfxQBrtJkazA
qOyhZGVwGzJ+qqZVDj26JhoY7VQgSi7c8ZGqy9QjNf0lMNP5TiGJ1Da8vxuxf5cq0zbDVes0Z6gF
1aLH6MeG2Bzkn36WwLXosBkmCzqLN/TL7smE23k3g1FOqJgySJv8K6RWKxYJ98FZwMrepu9Mjzo1
v3kArqWek98fwAQoFv9FlUCKZsbLkemGzdy66FWFFZHAKa9+fHIauXt0j6NRpwUjDkMVEp2lwelG
ty6p/04TeTswCKXAdD4EFHiCd5b5slRERJEeKwK8F6UV0PuGce9KcYid21ndDlSSPSql2VXE+Ej1
VTzMb/S589o3ah3ImGazo+taPcoHKN+0agUSNmIJgb+E6AtBJKnNZav7u6N4115uWzQabgeGJB3G
Y3cVw0jJyPAlTifErscBQurkjohc63+OSfWJmS9eBfWJtQghLCnAafaPCMGsXkumovGtOq7XAQop
wMU0ag4hVs+clU2Uqq/JH9mcsCYUzzPyn/NFkhGauirIxrPIhqEQK1xYTpgoehlNm2N9E2tTqHbO
xgdjcD0Q+T1q0tpnsD3OnVuSwfBK8TzhEq+gGeG2P/4GwLLsSTU/B1CeoQncci4q5kk5cHyhqZx+
YwFxDdxICsNCV6y6cqMNsQdYY9ROqDffOkNGkw5bFNwgbM/jcwAtfrYixag/cg523PxLJ4xItE4I
K2j6JSt5auybK6J0C+tv0nN3IHZ7vZW/p3VCwVF5QjPjqsikV8OqSfa1Xp4bc0ZldxCfivlMmJmU
S0iqPuYqdtHCvgWdTjdXbNAkKubI3ew42ZooVlY9W60mfop5ASTvgWI8zx8yfKEKMx9pXrOPmZdZ
ek0XrY5FARULyDHwdgypfkwZ6Pr6L3hrfmMkv+0p8CBvaOSr5qDtEBZ2Nsr0Sp9kgW+6wTdgfBVQ
6LEetf5CRSbpqmbRJxcZZPf5BWcJBnv3AWnchrFEDiMbA4EPEDFrc1g9FoiNO/hdCDb+VQYFlr89
y0u2GJH99XpO0xqJboBIQdl7f0AkihWphUiKbAslsGKmiopEx7/Bz1msUMBZOo3z9py0tFO86dcC
jq3rLrwFH3iFZNKhPq/NwJZTtDoWIDbJ3oWS9YegjFBj4QLF4wtpxVlDjg+o2KijkvT0lC6bYS60
ciGRw2pFALjJ5GmfPuLie362d8k2fxQdAiUIQ5rkdy/ZLwtjiTRz5J8oEjoSb3c3QKc/tPjYYqAK
3mIHSvO48wXaRZWlD96id6KdTwyW21b2qz1MnkLBNdhR9laU4wFpgRHNMhl8IPCbCOHgKATZoETB
jmacGm2Ol0Utfy5WBmiaGYPsLNDSnJrVw0n9bWfR1NdCHCmhFmez4kWUK8IVUOfh76y6l1mJa0/C
646Zf9IwXT7U6LHV5gh+eUlm0xU1m6AlsjR1bgffDnDXDp5IBsl0IdpEubq3QETFwpa3D09W9Hhu
hNNuqhQC5euCfiOEBOZ3Pg1tLIvmcRUUPGqQcolhour6AItf5oR02tQuPEkV9G466K/UK74tCR8Y
oSAmZlTia6uQmPI2CNgL5XhnWzJ6ICwnxuPJGiLO0r0xwy4B7qfhyOkJs/0yb4MhNTHD6uYk6Udw
ZDpcD0PykKCXmYri71w5O+MB5NVzvaVBK9zL1q7XfBFBgQJeiEGTmFx2QJrWpygOQWmDeBZbL3fe
Q9YuRF6iioSYkS8i9c9z3sbJ0cyOxoEC2KT6lr4vFY7c2Xw1YMHJuNgG47jRtnWJLBRTqGYMp87T
ECvtsO24eSwR4MvmtAkFCOmy0VFPUTjMbOizc8jUudjpIX+uOTil3DxixQRRYW+Egy5wlBN1Vokv
OJa1bhYj0sKv6pagUnXzxGsYpLcTfUCtO5VdkEAS3rFWD8c/RzPDUZb+Z5I6yMVyUNBbfR2Ot3Rv
D7HJ5/YsLrQwV4stxmbXywvjzl3iQ+1akieqas8VKmTMH3RVzUXSPpgAmz3VSGRm2NdQXNLWv44J
8j+WOrnEfIB2Y2FNqA2XS/pssT8/Q5vm/kqeEBd+2Fp6L6i2eri2JCBwkCQowae2Dx83EhgZqFhE
Pah8qItr78WOWv72KN6iR+nSpzGHRvFTs0dNyWKMlES2M4eWdOhH9LZLMPY7N08Zsz59FBW2kyaF
WVB+DE+0yLjNFpg5gf1okc3ilgc63xtrBeu/8W5r8gfp84FPVKjxKT9l+cjlf0Gx5pWG29s6YSOB
B2dCpc6ankxkkrd1I3JnaMInWNS/b3Vk+zkPj1Q8BL+q5T7tUFO1ucHq4hNQmVbHLcMiZTQNukPp
70nx+PM9YeQRJfftTLsLUUdjY43pJfm1y4J4F9KxGqmzOynldzfZX0s8HUAqJViWyA3YIQIuhvTV
A79EUIa/LMKWgbxhrsucETFHmi0nBraoVtIKFwe5ufzJ88zbBj/Ik7Qq7vjNKpEtvhlYW4oObE8c
6keXFOCIh+bR80gEu8HRN9uPEVpZHFAda4l0rzebTml6PLR+J/ULe47TC9iInkvSHtMMLItMP03E
AQD4eY4H7Evf1kSfl3Z5HTA3IvXGUWQD39dhwJd4GxI6dFiCiSJNFM+rZQKED9zTn6vKJVx26IPj
jGGWxP8rFs4rBpSXDG2ku6cXCnF/t86C6rd9+vBu1fKVtPFnFzr6t/RcL0vkQkBS7/9RhmCa2l8+
8x3ScBUreOcvDFJAHq4XMSNDDuNJx3FWoyEKuIpLeVzK2OHzm2nl14+AxlnEJVBIXE0jK66KySTj
Qti9vYFOK5y4GhCbAJ/qy2zJwrlqzPEa+vi8y6G7IcioYqz9UDxVSgsYW6QFXuqIabyh5h1EQbcN
S2eY2N3qut2CM6UofWz4pugMsmXvayfBap/tyvLer1s5DOvdwV8vh8r34Z46t0uOO3AMJGZ8tXEx
/pDTY80s+GjGwIMS0Ic9W8VeUXMTiyDK1PNojpv28+QCwUpEal/gek264TIRAeUnfdTBByQy9FeH
5LuNvyREBa5kEqgBTzyfz5fCXCQjdZTb0RDOaMxapEjUMRnLTQjK+xdtBSXuCLwBW/RUWRLc8hlf
G1UfQV2UdTqURJjDHisiIbqKVZlAwxYJiMwKv9KadHtAjqkylN1oeOLiVQJBKuY5YeMaO19bodRB
ktR+sj0pIboKhOfC4jopov/xtQ3DcBj+CweSIUyqbxMFxMtfN4JKC1cOJ4QL0X/FDxtGdLQPnPLa
POSjXK7Wm6CbUSMOeHzNNlPsejB+e5g6sfmaX+vA6K3QFKDdoBO8pYLcAq8mnryB4GXJ9/JbJjrz
y9+u2JlQkBTeyMd3fx7Ex7VGXPHM7LwlzACZs/KXL2NuAak6Fz1UU6HXQhU0PLRkD/+AwHoGx0e8
PVYH7kOvIcOhBY/CScZ7nS6SNFHxoZM6GzL6D/Vq2ZR9Cu99U25wAX+xj6lzwR1k+15E3HyomtHh
rJmZ6CaSM2nrnMJA238WacporkPuKacXEvJvzZiXeVV5OzR6OSID5egZx9ZiOg7arFxbxLye8DNv
8kf4dT4EEW3MjBZcEXVSkPqwC5bPtKF4F5xrFfy1DeB69TTec+c9rqbTins2lj5sdVdYYRSqmF4o
28+Lpu+obBzHA56IUxRX4Ho7eD0DKPBwNXodw9dF6JxqiPPh12ALIw5ktpgvDsFSyXByMh6Km+vc
3P3kmjaTyHDhFOXWf5tsOnv5EpQ+zIDDPsdFKEj+/8ds+9SATjWHrCsvU6yqSliHWPprPxxLlYCo
m1JFzqrhDXh7knyaDb61B/oB3UKmA8sXuIIkHs5w78jS4UE5jyPPEy8XmvpUYLIXtW2ZTPf3syIb
r4t2SJNWLvjHuNZQFr8hjMB3nNbi16SSiRVFc1DnbR/yotd3Le0rRl3W5LTJJZZnLubS2IzZJpvK
IP7/IUoe6zFB0AgmHBH/RWH51pbQ++1hUeOX/u5H/ajTiEoQ1RZHqrylWd/9RXIVoHIroNpiZ75M
Omt+w2nxmHv891fBehUpRQpskg7RkaZB5HpXd2D66QOuDYQFDtv418Ob7sofodKJiyIMRAYcUtHQ
Z8+mvdDbK5S+5LViQ6Y9GMnA1ZOrPk0eCHqSuzeKuRCN9zs5HTzvM1x3DoNtI5nkzXMP0BAplC00
eQ0dTy6F/rYR/yyE8E72a9FVyxkXyvMgFjdzNVGIpyLvSwst5n6vLk7pHd7jRoFw3J2GdFXZ/haH
6LH85d45wGjAWZad5Supxg1T9u9gqkDtKS9NlYV5TTfWMFVr8t0acsZAVblZ7jux6MoFyreLtOv4
CGj86OwUON/lM2Zt2s5OJVqlBCQdDpK2j0TKJnaFrAuJNgrD9vw0Aa0K+jVwC5EutjVpT8q2H03z
ovNa3IYNTvxh5yV+xhEJfqXq6/s6NcP7XqW1ZjR/kN2EzWYtMAzAyC9hK1ZqO+Xt+K6y6R460lx+
QD91kWHsPcNewxkNIQ4rzNCQnSCPDfYHVARRz0X1nCgE7XLAt7aGK0rmGLFLD6uLBct92F6r5ap4
yRIuGCsWBhP4fHmvlMh9vIAOLbeo0L/0azhvj6yHDfmsYeVpnCFNqAjTwVoAqrToAAmrvS+dL4M/
lrlZ0ee7ExykXmy/aNEkUdSXxdh533BcdL3374vTyobSiS/KJAhC7Ce/sTg8uL0keRrs+4NFj033
LByWHDbT0qWsZClfJS2wD3zMxbzkUfYzIptJkz+mPiXkHvU4Z01gAOH6+c2XwVXuBhj72CuTQ8Pf
YlbrLQd/oUp0wz0y/o8cnvzCN5vSouvCVDKBKOxNWyh8EQykC+qFFp7aK353yoRU9SzJxqGtFNJR
OSS+1jGLFPknHbjvt2lnvKZqlhF77EDiLq1j9//OvJLMbndjbT2ZQmvFFqK8OX6yhh8JhwcZfSLU
EeM2iVUVJEdji6A22DDyIPirPKkBtiZLzqxlDk8mcKV40LCQMn4YZa3F3LizWlvhJy/iL7bPtfJx
roEvi0baRLzcoFQ7IBqyH2NZwF+jthGHdbeXtcN0jgc8v2oA4T80YtQAo298hv8sfhntLnio+HFj
6vbLvz5U5E5ac+7ZoqekaWUnP2aEWEYPhDehCuySAxx21DyPqaIv1qrNrO8sF8yIg7dtW9mgc+x6
Yq5+PnD2XfGkJ9/VEKtaUsck7xV1EXgKt0aKWdTaYD8N9b8jumLvVnj9eVn9b4nI0BNYMeAxDLwE
83QGXHGq3Q58+l0eTiIB2h6OtxrlBCwjos0jquIZTWwUk22q8aJmQAlEEJFqHgGsMcOHwStLWrl1
7Qgk5vo7GU5a2a3uhbCLRIyr7Le+85xC0nvAvS05YYdSTs/jxqCjvrjNtqS13wea/lf96kHMm1xK
2HPwKHrqyK0bt7uVYnfMRkXBkN4BINWmsspnLfJUK9qTgZLDAuMKMINB26/p2BfBQAOR3pj/gBCH
P9djKXVRxXMuGplUqw+Bn0BWyHorAvZLaZK4M3/5+atrWL26fbeTvhvw2w/pSpm2/mAGfY7pNcFr
kjmH/nCI/ItV/EpUzZ54eglZzylIaSmAL/vRQXUwKHJwNGR8etDVR+cY0bmVXLJ7LAxvAxyHFw1y
68SSpDw14ear4mS+7S6oL/Co94Gskrgk7eJPw+nX99Yq1aF0M88qZLi5h5Fq0c23A1GH7oxJdDv0
i/9vomsUK+tpXOfWw2lgqU7bV4UoJ+bLe/YNVbAjzYvLpd81DwPRAvg6vM9GYAYy/oIQe3wgAn0t
qfu6vCyH6XF/PWWAMsu+8P4TKx+EZOBhfUG5QfPoAXqLsWN7XizhJT+Y7v5lzmAyA6pBrpZYi+xx
TB/59tZdgah6p/HfOhJGAH2WUvzxQf7TbEakZlRtuz7r0ufrFxUWrdnxFnqKvXbr9C4WUm77hPu+
FiDjvsEZo/NFMhnkBbNEQ4jKKGAcE3zuv5SgPz/FgssDRGAzPhDzoTtis0lUocGaaqF6S5ncmzS8
GJhh9lnvpEIqY8H75zs4FkJojikImSNN5Fyft3iH9rvEQqCZ9uCN0yEXi6iAp64lJiGmhkYLrl6a
8BN8G9q+r3hLnIAzY8D/L/62zzN6rQN96CjEqqr8JT1VJYpuDfMiAYa2r2j3+P4xuICM+pciIXFF
mw2esyNLV6H5g6LS/g3/gGOwZg576aEhVZD+ozjRRWgNzqczKZDSj16Vbv9R7+xO9KIEy/LY08zV
LIElQQJrEc0T7huOL1Wrwgk15Sl+vc+GKwntcGSaT3eNNoHe50cyEfODPP5ygVvaEpD5tYBuTy+l
CJXluxpMo3jHxmfqU1l6ImSy7BA8E4ZwpoZriuv2GJeNafn6IhJCrTMSTy0oG/KnSflOgclCMnj0
dfmGsxwhnb+D1oWkJTe01Ri4gR22TwVCNDlK/bRB0jRrWay1RI6wJNaAOZcR4oPmLMxdKxShdzKS
TX5yvLXxeFcn6tGk3Wx4ggi6nCsApEQwqV+XZ74y5jNTzH9PfovqA9yaPU6TBjqmeDkUgz9CchtS
7+XoGA7VePli3EgzC6OMeEr/71UR9jwoWsvUvXyTo9wYzt9uGJgsqjDZ/wOXNslLr/n9EwNuxNlw
AWBS9dkfc/9Ba8edJYa+RKKHxT94xP1eUa/0PV7xudm2kTuE94XEkFDMe1dD6JfcnqlKfCkeQzqs
ThQM3Vf9tzgQbS833qI8inwHCIGeyVVgYgRIm2vn5NPA7LbhwOL0Gd1rOWVk1UVpkwlWefFpPGFA
2gXyLqgE8eoKrSNhr7jOqs8T5I3nDpHS8ep4ttCn3iMThRf7KW/KpCxtEATYcSafoFPQn4iT2YcS
ITElVG3jVLrFKw0otu7oAaJc0ljAeSOhjDI9EsLAar+PFPr4mWejT76O0PFhD9f0tLR47SjGXd8Y
W8+dxZ/L4cHNK+cgKnKcX4yJIkKUBm9kaWD91C4aCqDwe8PRDjmiKC7EWtzk/ps+w9z3QzXquqA5
meYT5YJ+ZogUKyHP1ri0fOyZEscfZQO8paprjTLOJ32zRekWFRlZic595ZNNtXXEb9zKfroXVRdL
ey11f4Ba9A8zwRG0XdPoQVERzxnFD6J518z7nrtYp6HEgc/mX5YtMV807X6JT3+ncowSzkPB1YTb
ePqrYxGB7/5ogGXRbCsO32mIvDROZtgWPtKwbl3QunjcpPN0lWxFjxg/+IYvTTndbkF84BcTDIon
k5IYGKRPbNvOcMwW6choV+IJ3Iv7h5HVm9nJbaVBynszy/GJRE/4Y9nldmHGjU38LVT9rZW+/qt/
59/7he8q5NNqvcNyW0yVz9RTI17XTpj373sLHIfCzh1OcYhYoW3krEJ3pUETga/EN7Db13XbFJhq
RjTgZBmReBei+fN7bW/TrRXBq3yCQU5cZS8s2kOArimBUYO872IuY/xhTb31g1UpaxWwGo0LAMg9
l21514zU51HDv5nRgme5emRg7sUOeQs5M90xwN9hyhnllOQ+E71dfhuSBvMWmFYZKdBl/N3cOPZo
RHzjaRU/j7b/kHhaKPK3gIuLEpuKmEjZS7UWqRi/hjEaj6TPlBh3CqPla5JKyE+bMiRiV1u+8bU2
vPEOaQwCigMbQUEcqH6ok33NmOktEzs39o1KdIBBGZdWs/nZ8DXIMNrfveKSD/f2suqeVqLSlYmd
R9ZGIfNVcIyOK+BH0gCJZ1NV+o0P6PNNqmpLbh0LryU3vBnCWM4QT6oV2fx0P2evBsrSsU3qLCMp
TTRAKWn0Ifg/glvqe1ceJCHTjVWaAbyvyaO/pE2qBnouxjfdjrnri0ZUR98lEKddkW7TpBUv5UVX
mwhwfVlfqjx3fopR32OhquqPl5BmZnexhkJ0J6PPUSmPRJcoSGZ5BWcVdYYw4I6DU+FAxzIY3UTY
SZGJUXpRymbTnT4hyqIxFI7bv7r4HuOKpSDwfQ6vy+/F8V5B/ZQmQBDypklME1P4XGSrv36mYKHI
Ylq6m2ctqg6S/ZlyPp28/UBn5hdfkv0/YbqjgAeWYjkbkslhrFqXb0qMvH7Wg07cfPqZoXZPJ2Gt
bIIMVVLtX9BPSo79pBgloJM4ok8EykY6P8+3FCZGQ4RSnTTMS8uDjijc6yvfhFft6I0zmdPZrz6P
u8EfBzvfRXwS+yWaLXVEH91eE9KAH+Gdpt2fVsE34HkJb9ygYdGOrnoV3fyHPYvO50wlBHiZSrX5
SMTHYAKOswz/Ec7xyoWAGZKFb9NA6+tFmWjZAqi9O5o+/Icct2jjLh+2SwycAvwT7+2HMBHTNOgu
YlALN63xqjKyqK3bHVYK5usKMDf/ATXxH+nbMQHkrTWIbyz+PHHDGtQWsh4hbN4//vvLVTw9QW+F
1DSg5mo15naASKcqWfrmLfoFOnx+7iviwnDxE/ABYVM7g+ILe2EmWQ0RarPvLlnEAADImDl3NDcw
uxZdNyQ/79xQP9OKc0JYzfNFY9fQcqoU9c3KD61wcsq6TCMZG5vWym5mGYeyXLn0UpbFjwocm2Li
I8Y/5I5F9g7K+4WIlaFLG61x6YWhf6Qa84qW7jCIXlanu65egWBgyZDfO9dui+7cJyhlCVDP68Sp
lvx3JbSA9MZrmiuQdnfzEviVqOeBvAoV1d1i1JzXjjJNUJkqb+uXwj90hqHjp6qIgsnJWomWM4P2
tNQXUunLk+Qd6NntZUnn8AkF/UrarW2wAsS06stn9PCROEDaj9KcE1aKvZT3y07fmoNWP3ja9cxH
+BBM57gt8el/addatyLg3SbGnJku02b7N0S+fV6zO29guCj5lVUSGc4CT1O3bsyloCujsTxTDmhj
RA13OBR36Wy0YAONvHcH1QmuEsPUwjGRWlGsW8BBYQxZLKCV2uGVrnUANDTmFL+Abxe6WqMCtsTO
IRfER02vfLqCYQLwI1AbOS4oM1pPWT6cD3D1iMwZcQh760nxIQHh5SYvLfSPraeJ2zHV3CgBbDDe
p5B6JNc1Wvv6T9ZTdv8Lbz8vD5fwhsb4us4A79ylOL3MA6d81z5Bq9SrJwypYZCwpm/102TA5Okz
HNuHRsm9n4Mb4TqzHuwmyg4Vm24XzYNZXmQofPTxui034XQ/5787KgqAwjTN5I21I0kH4ptXx3go
feoeW2+cvBkdeds7j8En9hlu0z8Kp3dm6xg6r1Mc5RipRQcr7ShCNPPNvbp+YIi4U0A4lrZ/ldlm
VjckLvs00P10E0TsgE/2yt9v4YEvqIul7d2Qfq1FB0tUEUuruqylzIZmwUJG8Hi23i9eyVAOkFBw
jCwBfD0V6Vmp7SXqvLpt07kde++nHRaV1y4qU/BqMuHI8g3BWOsqc30YRdsvewghrflSjvUxHQ8Z
cN0Yt4w4MBic161QQ3cZja/plbXLYnbrOkkl1DCEWVpif6SJf5W+Cllfr1h6nLhNqyCoLkwCpWDW
Hm81kLj40Aou+1kzSL1KSztcp2R8aX5sy6cDCruVaEZpr+lOcarR6WcPlQVrD+OV+H5nEbTLgDpe
iZlnMCWrKZ7VeZux/XxIWqAkpJBF6bDZP+r/cj1tx5a1/UgZPxENaBQBPGF7NLLqxlzYWmXA5b/J
wvxRk2eOy3VCf7UfvCXqm5qOEAiDCNDWwu3QRXxWEA3pkjPFHnuDduG0RIsS+qsVzg85dui5q4RU
zH5KZRi9F6LsYjEI7TGke2LkAV4JRF/9B5xiWTirJqc1iVa+BZHYu5KEq5Vo0HCgNZLU0sOe50xX
3Dpa2Jer+WZl1rfAU3jaL69+34Zfo+uGxlHXCFjdQsewOUMvKcxE1tiYjwgIvV/NBGiLifUdwUdD
6Qo1y2YR6/ksOzHQiEXn9PIWK//awLZnnSdqxzC+2RrZd0VS+IFWyJOHPKHSfh5YbMgbUSnaIU3J
ooN00PcdkLpkFENXVRh5RtyPKbcxHotJ/pkYvLniawsiKGBUJAWJYHq0OleX7yZ/yMDYaSvjkaA5
ApW5N03w5LCRwa598y90MlWM/RFW3AT4NhL6Q2CmFdqUuEDA3LqlJFcudhPfV80d1uiQ3CSFuO2L
Rpum4mXP7gQJRgI3T8h8qOLpKTIwYQ5dAMa6uRe/f1jXjTh+XcVaaX4DoxPPGPm5SRUHqZhCoL14
KzZAXMVg7NqpYZBEhWYwpOMvyDfhiy1s0EzEhokqabw/zntmw0C3BenlQQOcKULGIeIUFvIpZ/Fv
0nTEwTjqBPGcUQFSgrF3i7yybNuKAV00I8yPN4nOIF9iTnpFPcFSMQMOlcLPcmPNk1Kp9YTTeHCv
4+V9eu5i3T35VA1ALnikkohSAgTTAuG64bfY2z1H4F+zzgJDgUr4iHrb+jRAFw9g8xWwWEkzPuY3
on3LtWC0E1VUN0EEuWepnPtoqT4oVccIUtyXhJVys+LXIx7/7hjSobjXpjAO5Uz4E4Ke3/AqnQx3
VJziNl5YJqZTbOnR9nBLyjtJlmE5v18+bnwKWsfzTBA0k7GllDQTmH7uvxcPvdPVRb3q7YdrQqdA
YnnA98dUpN0USCzpKk0pOndlzHOAdcEHk9S8fYIvMbWF4M4QIAee5IPnxcPuqRAXDzbuBrIuNGZ8
HTl+7oS1zFqFnMre3EhX1PYpGKB+92lKWwu0ea7DwEa3e105P5JjZ1lYPS44qVCxLAyEZXeOcXYY
qYaw7N/qn33wZVxOocG+jv+6AqSZewWdcoQqF8x1xuyLnzSRYGR3088YTNh4qIw0saY9MW/3kuxp
erAOpRbLSSyUPTU5CW8szBRz0p4aaq3ahhSKMTu22cAxWDlxsKvlyBwpNnHf3EdvZJdRvsew3Xhj
C1jwk58c2k34MpfXsI+Nj4HTDAntlzEG23AX80rtrTBnufFl5BqYRIqB/YIt9vn9AGt6vAaRjFf0
uPXc8T7tF5xopTcTMT4gH54C1Plp/zzYwYJnqmdEk5lkVqwGDs6zGgeyUAaGwklTFfHLxzCk8mP5
DiH8bdkzZEBpFnRvzZa/TDD13WzNJr1y5ebr6JOyWWoXU6KsqaCENSjAkBqDQ9yD7arPYb0c2cNT
EccxhVt44og56pcHJnBcafobuyLViyZlT4yKhDguvyywh3sVwuxB/kW+rs1LB4H8XkAmh3gZnfzK
a0atFFKYC4jQIMoNeDG4Q+L0n8BHPxvUcZn9fXcLCgtJKRczyFzjSdp4dkwuZysqtYfCNw+ruMI5
Edmb1MKIB2Mdv/B/gn1yAQsvmUX2DjIPbUZjR2L1g9/ImSLZcrT2pTqKHVp4QRuohosyOE6jPwLJ
JQNaCQcDrihUseXAiaW0VggVAsiEwFD8GBX2BST0ey8aWlwrtLZXWjqucsVKuE+8kattBOhPYfLm
XaiDLK0pwe1K9KX8hPloVNKrmlWNYo6opj4dRXG6LN7FIMFRESPjAh07YGNO0Jk1O+PhqpnBLOV1
tkwKRPRMyBOEDjuyDU2GCUAU6FPw9GD0pfYfT9Ryzai1cuSjRfxdi66nd5e06jlKgAdKo1eIaBp6
wUWs/AQI/9T9JMSexPt0NrJTZypFet+5nLBVPt8k9qPRrkdm+PiWHRPKzxbNpN6TzsxxF2mBtiRq
roXduyB0E7wG+W0cWuLMamSt6s/vupP+BsQA/1veg17I16Z59Me+yyxATfhM90fIk/1ZY/DAoJfh
M8USzXbPmzSa0PAO2uPs8KgKuY8Nh5mHANRLr01FJ7X3O4FxTVMEjaXkuuwH4DHshp8oF8RVPS+5
74TqsvIQL7g6vtwjeYmwrUxGDa7ENw0BXTw/onVSq5WG2ztK4wBbyGFiLgxFcDuJ+03iigaKsPuU
HrkkS+3qYT9CMUhdPAlmlIjSoLL0/fs3qy4tGHX7g58psFkFO8SlGbZ9sBhdxd1HJsddQ4iBfhFM
ZgA7YgcL/6ugLRkgNetNc2lOQysSG8mIyfYpPIVy6MLX3Nvx8z3EVJgok0YvCNyeWfOWo53qqKK5
tlZhbbsxIIMHsseBEBUYvqS9ErWCN6iNmFbJfX1en6hqKq2sGyxku3fTcJHTSggCss4uqJmrokjT
/tJqM9zn6SubcF+J9oeXAfo5Wu0B9s07mVh/KSXjDGKq3pdsmFKQbWQVSDShkzS5rjdy+uCw9iqA
7tHdmp7DXaLYhIRlGCo35Mk1mKGIja65ks/ZbKmxZb3HJThYdA/owifqr0uxzYzWGeGXV4cdDZyh
PiVe6sT7zeNgOP9a1gascpdNjVAL2NgZFJmRZIxnmujjIaYLDHlMvnz5/jNB/gY40AGu6DeffMCf
/dhHdsvN0MC9eY0Gt3M710yavQ18+c7f+H5XoKL6sJIdU82Ar3/ynuMAmrOiTQ6tpV79jvXBqnys
BuDTWfyYBTyhi4NC1JOrDsQT5Ln5uZ4hNHOINz0ihUvok7zJe87UiTLgsYZmsPvc4ILXZ0QWppHl
UMzoessNqdESJeWdvlksquZPRDD9DybAJ1sYseALX/IPtVOjdQsPSIvtG9XuOjUfOc6A59+SmVow
OhH6ChHw90xSOpO1pqYE6AYGiuzBupfqSya9vgpWvvcW0veswtA5luHR0uyJzJW6k3F1DK/DipRk
eWdqJtchgbkyTIqy6J17b2uHfTB7IAJPKrcvMhoH2DN+xlFO2gmdPLHghlPdYfV0LM61TD5/HDgd
rUTTwDEYdVU1fhBaSWkoPWZT7lBVeNs1+61VhHGTWWDBpG5gj5vK6pXOdgNagxiBXcAByVC68cq7
qqwwN1RHhVoGLRwFqbRPNQT0+D6lI0baLYMrPaP/nkMFDGt4o4gMpekImBxtG81BklEpTus4Arnq
jYrIlcu+CmE8+x1lKF115Teb9jNtNDwa1aQaeKHiz0h2lW3x7UR+wxoooe6vCo9arF0K+whS8IFv
T/yCtP9rnjDN48NuO9nS0dz1AIY7wC8NtU3t/NE+4WoHWKHbux3fHhvONvK07ReX6JhrJEpdihKK
PB7ED6uXI5BNoM5qCZGm03/wUQAMxucpifQJxLTqaKdgRMQELiG2SS/HKppxkovADkq1ctGUZ8yP
4YrcDAhmU9yUXuwVpVRlRIflNstw1sIwgD8wMDFzquwvUdImtpR+jtTqfF9WRpRFUc3LyDNOUQTD
HWQ7u8HN1O43oyEqO7/bmbkeJdN288PpgE8Ab99giDp5ylD88IWGG7agh02zpzg+zVWv7YMF9EDk
q3cIi1nlp0VyUVKAdingX6tesLLxmHgXqTAU+X2ikkNo6fRjI9JwkjAed+v6ygUiUfpSY5ELa8tM
Hu54fKq8B0zImo9MQ3iF+Sywpw/sn8Trd+8Xn+aIE73m7mRc9NgeEIP8mqkJGOZUBgWeWSDTGvXL
VQgxaspsghz0NMCuIMCuU2Rm40Lyps7qNv4ZUFZNxLsDMGc0FZWwN1v1t7yC6YMUnT+axkDuZE0X
/3yD1M1B1azQg2LUCUNPVkC3cS7lkb4uwThpjgEy3LWESJ6G2+CU3wiE1bl0Bemg+shqXod7uY/l
XWBLrPUSZ0RLk/bVBFf4PEE044U7FV+YsJNaiVC9MayERcW8uAUr1diuBz2soFnrnwYuF8cbs9AO
b1XXL04LgorvyDhCfK5iS+Sv7YySLx6SYvFNXcTJJ08q860/j718khjWbnHJJbv7hXmn7PscWLxt
A5vaRd5mL9DJ7Mxw81FT4ymutWQ+rMOc0eb6ZBL4U3j8DwzRZN91om56FNzQe0ArHVKkEpqz/oR5
CYQo2dQRCt8zBV5XCDjmE3B1kOPM1KpBq3BW05yQFU0TCn7J7FEKDJQCHGfI3thCg5Eh00GolzJH
o3vrgzSSA7P+4C5QsLpljq7XoNlQaY0DUaDISd3rlIjZEoL+G5CBiCyQ8pe3isRiEeJ9VeA25w2s
QcEdT22UXOliRSQuKdB599k4fQfd0uPHD40vM+GxluDIHMcEZRe+tcNdTjcefAUPKg3zgwNV+xMH
Us3m6GDkeEHTaNoKg6dx3YrQcrr7laf87K43YMJ9JRuY+P7T6bDh6manw9p/haHbBBGvJhvaEZ1x
8NtgrEcfQDnCE5G8NiDLtIBCEB/CGH41pNOjXrLJ+NC+YnXqtUuMFYVQ+Oy+MruJYEP0QT8t3wdU
fCV7T/1DfEi/lAHL1ILP2Ahg2qq05vtGZUTZWffxKgC+rhW2svG18I2XOsOqYIYsmgyO2kTARIkP
AwObY4nGAuUEjC58kTMmws3xKsPWkzjYaVwJqEoLXuhJn6yDNUH0E1B5uCOTxA7+XvWWLcXnHdZn
KpAFP3oCJhLFYgK8Z4t00sRAmL3gyK2Ev2fmf11JGmU0e0nUpTg9kjWTUVWmlF7bKQqJ2+Sfh5UR
GdycXHctto2R6JzZ8aqqdj2wFcN4x8hK8ZPrDpKwkt0/WjpLZXT4RVrNO2ZWD2zHzYx8Sxy4sa8j
Og6UBXuKmCNzcg5bD2cQDy5bj4eybcKjexc3sUSwZK+09LDYLSMQ2M9VHjmM33i+Gz9J94lnFZE6
YSwwUmmjvGaf0YVLgznVuaiM1NN9wVIgADDk9Sy+UK2AvBe3+FKCOnf+jVoIZojyLdNB1sN7fKyL
BgIhA+WTUOGllJUX9Bc1PHw619MeCpaeUtEVwguANbziGcr27xZXAXrrW90J4z737hMx+euFYSTi
Hm6OVhewSjve3845VvBEJTCgnlQHXH8BC14YwZnSL2PN/gT6S93s1V2VMCeV5B8kxE528H2AqqTO
S3RjGFu31qxHhrcIGQD7Gpb2aHpUY3btRCcDi5B3dN932TCTvxUqWTMNVkbZavc41ctCDfH6Um60
MkYPqhWcoj0l4vfc+HErdXaPTfn7mqu1N9YoR1kGXP01yoaeqQpdOgU4q3z2VWIYZgChLOBUM4IR
XgNkZYqX1m6+icdBtE+rH9kC1lQUNk+AJPPbFvgHq4Ceo/tKdWePVgaOq1G8Ji5GTqhyiuRK+eqg
u5tVdeahfOtXDqzgeU/oeYwI6pN2swgZB12TKOa2f/RWCNRlNWdpBHvK6cNlLOLA7exujJ0dykMP
VqtdizHUcm9xz7dkt2uP/E1QOgGe7xY+UAh7hDcuZgFD4h7cQ3TOb88Jmp5sAXyeaY68PDCTD05b
ii5RriAi/0JrABCSwNJ7wYltCDvouxqAnn3sHNwmngl8gAAWGV9pI/K3jwRzeyv7yHuvbe9GP3gw
LfIa1MVsKM6ZDWmtdG69Qom6q5/AwDvb9uKMS3sKtbJADTXcaO8Mo7qFoUI1Vd5mzfJgvd1fugQ2
88Rr6s97lkoSkcnOSNHTO5Z3sKM0C9uirHnxX4jal3PWG53HW5wMablASiJnDvqVgWNPsir8QLpx
M1YqywlAw0jActh+hN1MSOqQU3Qote5G8afntysmE6w62YdfBZEpJXkarcMLM1iQ+hgMcpbKZDZb
0ifmGNIuqSEH2ojUzYRH320esYMXcxS0No2aNjZptTqLb85W7FqGGEl6/ISIa28Qc4REe7cV4m8M
N3583F/H0K0XOZb+SMU2loFj40YW2woiFXCYtLZTJxEb5HvgskRFwk7B69OH1pJj47nobLuPwgES
7KaC6egMWJM1yscPdHTSDllt+SSrNg3NIkvrnBJjk9U2UosdGZl4dorbZeqMQwqO2ycrfp5l2I5y
U+n/9C08YmmXtoYaUjQKXlz90nPcHXJoXr8wXAXpN0Xmxa4qf9YaS7SGhPy8rlDif24CfmOqt/lT
BxPxC6gIu9HRzgI+iqUeg1+UBofGkBH/LR9CtloB0k9RUeS3GvUc0K5hA4AUX8/3FgkJfdIpnYtj
QKxKXWpt6idx5KgPpmgJyDyk6ALZ/C4v+ws1rOatx+JLltreZgMhwY+D3lpy7quI2r8T934InU9w
j1T4td1+dEbTONX2Q2XgwypYEbO+cNNX7gpSSMxo1EIfikvjvKCMv1b9Vz+RiU0kf0KHCxYJeiB3
JAnFgwtXygrMSjiiVriDPH/OM0v0v1NqNhK/iwoc7LNLwySeGWGFr66E2Ck1qqIBNHz9ezN66g7M
AQDCaToK2bNC4Dow97U4otX2r/rj4KwsfP/qKG+dugotz7rgj+b3BZDuBxnKd8mkuPjV1UD2xIYe
Rv1or96G22H1LcJF4UH3D2XS0OlCsLv1ep/tsh76p/AdVPDV1CU9s5fNhBA9Cma1XMn9XFNFdpbo
vNF2pDCRUxpKPCgFGiYcdMh2lxqXBlSjWIT0xB9lAoybbMVMD+abGxGI+TdgLdGpgPEdtLw3r3Zc
JY8OhBIHjLwin7iTH8xuJQtZZ4hmPWyeXq8DgSM8xrYRIoujU4WiX+GQagk3TNQepsIoGFSrEnd/
Rbzd6ktCKBKhPygkIuEgMayRnNoiJokwr+NeMOLkwRX2W75BBxHBYBdg4zzoGef/Ub5E5jHjBsQE
CrtJJYj6gIAmgca2ZMifjfajmFlc7PdXUAeQ502TgXzEiY45xCL9v5ynHNiU3mDU9xrcNE+FcDKG
TzS7uUlzjy0KN8Vusst0c3uDPuSuamFVVSXRAw+ulJRX4dTcounqfIpI5M0qF2UUzRMxCohS7B0q
Cl/IlsQspR0ABR5yBAtiKSVOxEkGsWUh4woZz8F2aoUKQ0zAXj66VQ3tnAVHWMemxVOHI4u4ulSo
lgEqBTpKBuVgAx9voZdqS383HDACJozn50TdhEIvQgkJUBR2KJz3TspSDqXYpIGVy3l9vWStfZSj
lZs4dgVfuO9l1MdbTDGxcsF94W0dbfB1IoXUI0gOR5PO0ke2AZhib+xa8OI+MZEjQskMcwVki98E
yLe8/DHMIX83U/I6svOLIHfYPWdUr/Ifvw5bZsluxssd0RebUTyqStLum698clz4PUNzcAF713ow
lxYX5RzmkWRbNFg/VtkGI3yWVqJHTq9HnxNBXPMU64M/q03JFSqi61k4f+Ig2itCls5qa7FHeR9a
CQA22w9xBQ92psg28mfhnjB2JuJ5d0ZSohyJPQk6QT0v4Wn9fkgE37p63JFOevxKhSczvS+6f5fg
HSTvGNBV4UkUbZ/jQxqzHwJWQVnXZItRpUkJexjqSCHvm0VPQJUU8Yt2u4gGb9GtZHE8fbIzYmDb
ms25WJhXqEsDD2p2muLmQq9PXsX5fngi72/AL12CsyWeMTKFLYZJfaWxEWIS4gv1Jr6ty+gie6+X
Z6ilRgDt7/C/OSw5bgQJSutT9VcoQwYv1qkQDv0+SBCvDCPx4CB88njMkE1L5WarSZ3rbrRpfK7Z
/zI08pDEzTgHWDqJZOKpgmKzQgH1h9wW5ZaBg9mqdEXvd2uErciLRm3ihVNw5noEvqom4dxSjQwr
XDdIEqwbryCrkRCfiBf66J/6EedsxAsP8qaUxP2vV8/vLP16ZWWBC8wGeABB8bKTtf/1sU5VHhHC
EI0ytqp2WIUD6wW1A7Tj9B1htlbUJDoXTSo/Z/iuDatxOmqkb3xEZz1fnFCjqnL75L1ImHFpjmeM
7nUQipDTRDTmddO9AlZ9eianBeG6mNvIOeu2Aw2McLG+40tqsvtHsVSlQ/Wha4CzmGqOzwPB0xtE
9uiNjlLDKuZPPd1ZgOx7V+I/bhFw+4j38TWDBhUgQliEl6dfJOrQ/hItgUauultM0LqnD5L48K0r
YIxquo6VMu5OBttvSO5CvcGP4Ornt2KJTF6aDVpY0Yvc+tsXJCKRcBLSt/LHTKKCX1/Xp0Kh+/fF
orGuN6cUcTAqdlYCJx0XFU6fbcbPqEfBv23+7CBhbi2JqJu3K4kDtdd+t2SnDyOqndhGG0gw6Hpt
xEiy4XCS2DGoUXQF7cjje0MWg+UlZnGmnwAhqu/ELQO/WfJ55jU9E5twl58PEnPVPNwvVwHYqSno
Hrm19vpMcn25wBm/dfszbBSLMP4zPGLsxOZe7TKbPdAyXjU8xoro6ldPUjjsfFocO5YAQ/rNjW44
jafYZX3ymCdUhJoqWjLNhln74B0vR+URkmv9paFUvwsrPX671DrC89VAh3Fgx5+08+Q8PApNkZtO
YBNBxluflSyJZPr5dwl1TOoVMRtRwMvT9Km0n6jdaBrKqNoY0xzrtla/ybWAl8tM37tk0l8d+dLj
3fXTP/4e38zi6jq448Gr4syVhmzVKIeGB8L7joTn+ZfHlqKEpVxUny5eE8gKgEEsEJHdltpy8Al/
R2TrLrRk+FTyCYYubRMdUIeG3CODbY4q8LcR/z0/hj0HPJKfZPp1oemLE1xhKMFEdGYJfzrWMAfX
xoo/et9ZnXyxyUf7k5xROYmxlRd4wjk6jz7j/6BYkWt0S035lluoxaJ8pX1UO3Ywet2tslzVqR/6
5fflFMpHyy280JPe3iv0gxuwbHGJ+fV3qXdzUqMHpMp2M2vh001RbRMV47fFjHDcPCfmvNaw64kP
nvhb35nc/LpFQn3dTkubJzZpga9rjqShIBV25+zck0Z/QpSoZ7Yzpbq2rxmn2EpIMgt3cseEvuB4
SalS6gPYHQD80QmgZwNcuHLcLBZtwiJncOm+dgHrRWAgDFIUke0PH8+9NAjbSx6Wz+klYJ+TAYWS
s0abUmxs+/FZo41bOR4+PFNrVd+D8QKpPP2RF3J0MDp/jZTqp67sWqDPuRqeg2x2XXl7OD4quY9d
jy51TJSn3P48MJWVviV4inif1MNFyTcMwaV1pxULrZyLS1qxSTB2BXRsf2+YV73rqVlt5rFxB4Ur
vZL7ch96XWUCIW4YBwX62Bb9Qc9Vh/xW91ddMp8L1/o5qpT/cE4eh926WxxhHDsHYvH+ao8Zpg0r
qhWloi2oXo5LeNESaB27HoftsdI8ecY3jKwkQyQC6prrkQIRpdMzayTF3DigiCH6QtJXEsoKOYTL
VywGj3BQUhog+dQsdj/LMytBjlywW+frxvo8ht7Ke4uu0aY9Ofepb/rfajH9nloZWxwdDtdm7IV2
fvNrgsPE/9GpCh+dVcwp8OM1Ia8LBJBK4raWsHqQ4775IgxskF9ZZH3RE2J4TbQYI3t0gX28T22k
d+ydvIHFPqJi4cZY5E/8vqDavS0VSYqZMbmktn4HU9+tbRKNe5CPoM+zFgckVFB4e0K2/EpkVa8n
rUazDSMCu2MpcddQ3QbWBZaLMti43ybyBV847suRx05VIhy468q9D5rbPnEiPYQjDdBCn9/Vo274
OSld+N87hrp8BOnoaHtAiRZP7yb4mamrx6WKIvHdtldoCWQCTNlFbOWAXLlcTj1ByDDSgO8vW5qH
OpTz7EZywlvdqZGtCZlMfqio0b8JfIWxgo0medsTQ0ZheOiIQwEzC9OKYpR5NBn0xWBSpxl9ejZG
3HlS31Mc7SvT2yndCp8vv85puG8JOE2GBvPN4ZOOb60PBtZUbRvuWfnfFj6JxV8tewT7mMDyJCPk
TRiSwJAkLP3+ZHpO2pFGQDbKAUkqPbQ3tuwfjo/P+sps3KRG31qIS3E0Umg32VJefFF0YHGlVNpZ
g/aSY1W3fgL3/GDStGQ2ntJapPst2lQXkgQ8q9zjjaGs38hFYg/XFw4T651JmCXLnUCbi3iWh/5r
OmK/Y7nvtfXJ5t74xlDRgQfJqwB3/VcZ31EDzAmPrEkylEy9MgjMn6jfOMKOL5D3hy6aNzxniMRO
Fa63JkBkFIwbNUJ+AMpA4QGGBVDB/1pE3uNk/ouBrNdYy/gujnztMqZvoQaUdcSui7Ied2RL6mLw
39LMDLVrWFB3Fs7kf4PejW2/Ul+X5S3Ws4zjowXFkSdiXBkLZGb4Offt6cf8OxXU5GC3I1oS45QJ
niutWhljtBntfij5i5g4qePDmiTMFcvgXYu89Jh/XtdARR9vNDbQPP/nOi4orEoTWm/BAKKF/GZR
jhToLEFOIlzwQycUb9uHcjDb+z/4yo690NcJHg0Mc62a2fEySd/eS6bBbEgypdOHq5idzI01PDcY
BkFB5IFEgG3MR+zYKkR3x6ywqyqhIiN4WvafXK6hLktBDdlti9qOwrzlWDI3H3Vjq9cSh1fSmAHY
+5NMsFghY4e8DKtRLp2C/+GpCDApeSnLYPB2jVzhpFFzWjsb+yRyVEhdHMMageGUqG0niy5QR/yM
hw3pRkIb71533eR42JcASXncB/PXFwwl+yj8Qx8Zyskp1LjiIf5uh5Jv33LQKb6zyOzy9d6aPTEt
sbHW/K9wW5D0O9JlqAYyoj0Q/um5BHc4P9kKDDJ+DjV8mOtQrelmw0r2lVYByIfLk6bEmMQAWlKw
rS73UG0zObjoUiGHBJ+L06Nq1Rg8balPpIuIveiNmNyc6DVXOKUkB6mQHq8Lwdan8xOg5BlePkrk
R1y/rFnXAYAtu7pF97cbD5OjekIrq4M9kXdCIK2ch15CYtHSWOzCt7xv0gVkcVUoYfenoA3ZP/aP
T5sG47H8sQwKd7r7Qpwvc8fqLs6+Lwq94/9RfuxgS84KuWqTJS3hWOr8kn8IQnbHls4jeGpsxCpi
4EIqexs2EWuZZg4GRloFPwE9fV+C08kudUnPL8YmbDuAGZNxQbaieU4drsN87vKAdFDvm4kWAWHt
EqzYdbMIYMg3QX1fjxlkBIZMtA6jVpKs2FpEocuR51dDEOzEXazrQSuK68uiLF9VctTFc3YoAv9n
5vpTfwQlyuT2lm7jm1puScMDYRiRv3Aj5xrVHrzT78bjIREXjTQoG3FQFmTyK69TEobLJ/747J+i
V24nkoK+rt6seJCGO0ygOaSiSKawYbmq1K3y4qG0Atey6ea84i4DGJeHfeqXVYBd/3nShBP7eu93
TP8hCsxhL4bVQCNcHds4s8JnEtN6Af41MRbds2QRvxnJsoCWwcVlkjew+ZsExOQbusWiFgCvGJtK
F7/PXRXpIIcwjO8/qfNli/FhnSsRNaQdj41w8clJpQymxPQ5nyJT0Bl1Lsjy+e2Zy8ud6gti34t6
YTY8Gn60jjUStZQz+760RffSAq0if2SVDNbztZAH473aOR5Hyr2ctL6rVtHnnCX4ycg809KDuAHi
fv9mW2ubQpe3sUnvB2acoQWa+n0rq+2EoIMpW0h/N5oFDkmptaV+c6FUOHdyQGXzSGJgvF4C9Xxz
zi3U9wB5xn5YtjbFiOfdfH7FdM8uaVdvYQD0EPu9ghDuUM4ZaggZylwIl28dsxi9vAZajAsvMO+M
AHJT/BlWNtFMlgxfMSx+kzun6U4+d6QMOYzxalUAdkQmNSjzabieYP8AI+Q8RwoEdkW74eB6tmsi
EXxVxhqdXvbSHpMr+u48oEo93lF/g8GiQy+gE/RxBlE3bQbTckRaPnPuCj6eKk44MHSaCASHy7I7
CyAMSspAtD83PNTf5JsHB21Y+sNYII8OrsYDjtm6hyEq33h+a+hghpCW2QQfgPf3Et4GtxEEx9wE
DaEL9b38GBpizwfvOCXqeFXlrS/HBfv24ON2yNKR5ToPJmhK36E8TfIqkV5jGFgolktnCmWr3UIl
o2L7+X+w5Bk8krrUS+IJSFWHNfva5WAkAZOKT1I+8grzwn2DO/x86tP+mXe9jupbTylnL7/gpqX6
4ycPTjAxtSkFy16YMuSBNlGZIIEUgc40kz0DThjF8lKzBceHl858sKu62bsEb1PYpnGDZeDdbwNw
8J7CofQb8Rduxb2kkSznhzELq8qq3SCVCow/XtItGdBK/iZbrtNO71LzEWi8SrqK1fVVJpAwpaGk
j/3CnUJSSGlxH3rv3JNcQieeIkXG9x8+cBXyciWRjaOGjjzkmy5hkOL5uNSV4JtFunFTX0tYsray
VMO2CYVgzy5B9fkIo0/yFefEyGBavGiDFT1TbhpA4oRc7LUiGcelTUoqoPzA1tI4tMXQC81ZT78R
4m6d0hV7f8qQBrt5PvtoQInN8ZXS1i7zL1Str1gqNfW6FFPtqSMaxbUMzCvE/HWGXchFfeA7eW0B
jcS70bEXGTwOEjTI+Gsb4unHC06qBOHSrLzHRk7rYiRPGk5+kbAm00vbN/3CL/GQmbJDetZs7u5q
91FBGkEVZMogipPg2q0kJtESD4rz/uphhNRcWKFikLIIOGT/9xLkSi30TyaLe2bK/KZchh8PF2I5
7XONGUn7VYUTmfnJdqe1Per9hcgG9m6PY/V33O8EyNW3i0blGNVdy0JdMxLPK01RzCo1cUQMl1ey
mCLVrSa6aj5T1qBginb1QjlNXfmfFHnEr+UYusVA/pfrbLkZn+TritSDOfnz5fGQ0xDR2+1+aKfr
oenF2TC01WG7uWcYv8sxODofNOJzNYbBA9Ebw9zQnrT6P9JAUf2C6g2QtVsPoAqVBRHky/YiXhQk
DiZIeG4IAeSGQeysTTDfS1wAuHgTOmRsJ7MZnwUzpNuDpQeItzsVVcQpunfn94hlb3NRsnKBsM2C
qGJfPhcZcWc17KNh68uzR5EijUG8FWnDR/bd+2NYskgoISNTq6qpuWXba5uqZrt2vyet8p2jMClN
OYj1/0xq5bXrAhDjVZDiIcB4GvRVpnW5m51Z2K7ton7X98LvrityXLZ2cq4+G8tSX6lBpdryauV1
XcmFbDCYvhe5UuBIqS66S65tnIYIEkbGyC66oOGwsjrHsOPbh1LC0hy+vwP4KFAOCb5iF9gqyp9S
Vohnmy9pyO/Jqer8vLShWNO05dsVoroTBQA/s89SR6W5U0pyskSkJYYZn9atiGCUagssxK8BrjtG
4eZ7r7BWQOVqD6osiASTEWlys3z5ggCmkgrIoQSqCrT00nfeFLL+KKW6UXU22jmHlsSdvBb4aMg4
sZAEcug57W3uoUMtJsYLVuwKDWbsgNySa6rqRBDa+u7U5hH3fH28A+f6lxUcdz3k/5BhggI5H+Fj
WfUKDOTPsqjoobCh4KujnVjwVIUWFetFPuqM5E7CH6YpaF7WpKN8MEgufxoauhCDR/rWD5twOR8N
ogc14TR29Dd7DLR47FuKWD84253E4cUYr2bNcCIbDW2I1WGRmifvJ9l2GKDDe0cnodmhdWJ580FF
4/q+BDRNJ3GFd4hwCqDiymeYVvJORv8omM3we+kjHeVBjynrBDwLZPBUgFNPLYGLxCEzGbuGsIoJ
I1CzudZP0aVQcRM7yRFThClJ1vJWDEluEFSGgTZyQkBRONfiWQjgZhKD6xe/AfzUvCppBq90CU/F
Wp058ZtrHy5BrvTd7lgDsMTPI7lkgksVCaWsK4KwIikrCTBruR9dW7FY6f51DFZKrrehdWVQ3VxU
UmAx4kDRiAgRi8sDdut5Vq32qG1LOnbNDzYGObg33LncceeE/UNNkqRESBbioOYCM/TLh5PxGOhd
AhKTMrZQJIVVlG0TfpcXEOzTvTHPvnpHKCeIoD6TCw+tCfIesAr4OsmCB5dsf/sNz0sR5UsYUmqp
gr4RSQZzc5EVL4487wun/tmE9vzrv6rhDG7jaNp541mRi7gzgWIq5v/mMf5hdFF5fhTOhxTtraoF
9zGDTIXN3Q3qZfZr88g9REXiIHdT+zChJEaPdKhNyUjHjywgfTb/CqfKtrtZva3udXZt9ybK1/zQ
kAcDhM6ATb6kVpm+3l0AG+qjbBucT3DOoPqAl1p9DOVrdtUpfM+UsHIjYhnuXF0ND+7do3PWUHRg
VIjAX8R7VyrlJ7rhN8gE7qTOhiZAY7y/KogZk5xJLbpak1suhVt4Ig4M/4T/069u53C85Rz+vIda
S+e5FllmWqLirkaifFOBmVJwF9Taqrex7AaM3UYzG9Tsi785I/ahAjBRaaWzmfinxTfqG2FP42kj
Ahb30YcKyntpsThnp+h4urOMqIRyyfl1vVX1kqP7rrbNkLxvW4YqC0lEBG4jeeeasaby68/lfkDv
7PsAn0I8BG9RD3vC9S++Yppmqffm1viS3gS+kLm8xsS2pNk/RmHePG9w8NU0n9FhNG5caCYIrqVI
PT/MGAEVsuzW6cDGvqHhc3mKA7PiKMJw5u0V7E3oVrI8EPxMB/Qc5HCstOAb42QaGoZ9ZpPOKVcq
pT8G/cKfDgJQEc62nhWOX3nQXzQo+rMD40GXjJZWjUOCLdC3P+esbM0yRnT8WL+86JsMcPSAX9/k
rYWvY0ekNtrXzS/CkjC9RACpoGx33HIXmeRxBoDdxyVLjTba0ONvQxb+Rm1uhptUNONip/hknHLG
ieBLyn/KABppDY6jRyfUnkL2dz3iGq+iTahj2Q6qmQEKl9Wb/OAOSdzz6mw1VQc2Exiy4Mj6pu1O
4rO/YZc6YeIOq7/oGbDrvZxR8WdHo1uU99nllNp4efLnhloekfO7fKdp1Uk0sTbFV1T4PdhXySn0
4LZp13ZiJ7axRTgGjZOOnJZCc4Tr2kPTX/+mDtlWmt5eIR8Gm+C/sXc2OwpIbumyRB2pMoVf60QR
TLRZ2/f0sJU0h6FO06ujynB7PyvcT93iSWcgv1y3WfiyqnMOQTuJHHZTQWtq5NNw3u4yy/ltfXVH
txjZ/at578CVHnvowbE9s9iNlHrrfvxTbDQVTCtItxFpGcSrBoRco+NrdaEKRHzxx31TbI16le07
Koa3BqTnB/nqVBFThUfYJKXnSS46Iqrg4J7jfW1C127i5H/b5ePOSVdiT2Q1Uj489YqCJyAQdS2g
leCpwxHJcwZWgGEvMhNpbmZ/L7ApBZ0d4QaZCDT+xDsUnTj99elaSA5yo42yTH/wNNDK8zmSS6t/
VgNTp8OlbBIbQrftLK4xuV611NUyVGfNmdR8Ga4KIkCFM11LHuF773/Do3YGxAZDV70CB1PsZgm0
o2A7cZS3dieDVFGTRoUPww4c7eVjs2qusG8MHx0TQS2IdiEQc2a22JUzTzksS9XmyNAaL8/qIUsf
EZYkTFMzec+O6k35w3gQez9TxsvrgoJgaSIzqyaHDiz7VlpVo1SVlCYCJNgW+Ee1jjjV59TBkIyw
9Y+fUItzAvQXv2QahdqayYedyOG2lVd4B/mZ5G3pOU47/gNbEtnAsXTVWig2MQReJ42hUa+OxGHA
mYOxzB4GeS9aBmQ2dq3DV8GS+ZVEXhobChgTlI2X65qyQbZfK/kpzaO3RpuquXgDsnJOHwEtKr6o
ZdXJv8cRhdvCW9sqth1jNA/aJGcHo/m4pbbYi0Q2j7vPCxBFWslba23PQ/XW5TS+L6RvbMkHv0Br
Ke+USyf8YUx7DxRS+MMiIEkMeQMA5LonlZ7UoFLnzPEiHdfowGk3IXnp+u2MIiO274JyoZN9F63k
RGBlqv5D68B95DwlR6nldR8BQr2j38mXBtSKXtBI4BhV+HHBFrl/vi22Xqub31oUcrRKJZN7Jv+O
cZ4wu/dkf3gsb7vGRMyTkXke3LmlivnNw1AIV8ywzqRrrtLg4c2DC1Yv6auvqVl3euOgKtfTXNg5
l4W7b7DlIDK9nm8q5x7HlUR0IWpWjTTD116Tf1BS4DnM8uAZRf74tOIXyruSWCRbkNACOb8EDZsV
KoUSGCJOsx7oXlcJAMbxZH3QwhMkGgf7/14FIZIsFTdSRejfWNfjPGen4PlCSM0JSTuANn8kg6Fb
VQBBY9t+ggjMopAoH1UP5ykoEixTWlRdyEQpA32boX8P+1MVsppapNng2iNGM5zCoPq9GpGq4+96
Jcimp+ZuFhP3AzSyb5KvIHipPbhxISeM6QjCirFKrrQ2YawyYPXI75Mszp86XIFS52l1wLV/pa7x
8U2i0eHU+cvnQFYE1Bd4U/PwrXFGX1cX7wJTyEaO2YJGlsXrNUfNZ09LAo1KTJV9Sfw+MUgCTk/+
ok6CXwLD8e0zUnQBWVXNAUYymvYmglUuG9yHrIaeoNzqpwC4I/jFxrsAl3zPIVuDkVjh7oUWintl
4G98Fx7Si7JeW1fY3AVKg8ODl5o+R0o7Ctdeu/akNnIDA5I8gtZ8NrhIQSY1c5QAqpZtafRAhghm
DZ8utUjvcNPeV1340scE3ZjCzPPAzVNun9+dsfx3zu/NL2RbbHNqk1VAn54sDzT02N6BT414P0A7
CplSXDq1nG0IKQ0V+34UeOgz701WxUS9VZFiDVl43lCQcdOGz48ajYc62YH/ayrZZr7LrNoXByof
Xy8oGUbC41KSa4l0cjub+jULHl3yrePvd96NUBLl+dFzJtY+a45vkKFYajEutGQ49rdZ4+2mVwox
GMOGbxNNuneU86eIhOMQIZeKbJbWWjKKE9SfpVHRLUVtpNk2EjAl5pm3XHN6C2O94h0ESH9HZKez
fyQuej7F3P9LQvczrTDqdULnlr4QrP7cALsV6KoFo445WQPwj9C5Ohn7wcQyDDXvXVoUhM+5nV+k
msuqlTSp9QRdOOIbUlbkHXCp/GGJ73Nlm9s05asYDdTa2pKylMQ+FkPEQorW/YGd3a92ekMr4ihp
S+ASeuyjajDQ8cwQp4PSx/R7EeCSewVCciSThUekb1Ch1R1pfMcb22Jfz1Gtzk36QKXq3xHwAndY
6lyHB2w9aBabeagIZObRSP6AViyXFImYiMbv7bLYDiJoHfTC3va4PKYRV5ZieYumrNmrc0Ot8eUR
vy8CSQ/H80ZlUadmMGX0Hj50J1wvbqd1Yd3CobfMnrdNHd1ebg5tPGhuz2IG6CuR72w9OYo6awS9
2Cb+9k/GiEshs8SlpE2vxQ6B7sSm/hC+siP6l5ZY6AjUECZlngbfF4NfGHXO/i71LG19Qz02H7Wx
JYnSFUAyEDPLEFKuB3qeXcGTL/TALSXJgeKye6cz6+sNbDPgrZPN+tt03QhUT1pEjpOSIRR2zelC
ZR1RIt5ncXWgsC6wWbpNUEvAu3Is42mEgWZlQO/JhAucNYAZ3V6NBiv3Bf7U1WujuL67WGKp00At
9KHUzcvEvVLrkSWUh6/uvsi/BHLy990K9tO7fy6rbuV8T3Zh+90yBXkUSTHPfQerZHwj71rNnZ4W
aBTrMV+Lftg57Y3nwl+JcJ0tBQhsPOj1yMUGjnHAsgEpsd8qZ7VcV5YQiI//Vaf7mzF8Eah3sQ71
LZK3lD7dtSVRF1vNPu9Hza7Po7QRJpKlo45Kw30sEKzyg0rKDEmd5SxFKxnz3PjhyGrqNJaw9lgh
NPP2v75rbOaB7YY6FNPOec+YpCcddHo6zT26YM3D29tLaBaoojJMsXcOLxs5YYFPivGLq49Cd/Ne
MUp1SWW011A4vI9T/QgMFOYb3umAY1J1hX1yOgmf3iMcVkWDvbGb9S8djir8Dggyp2DCltOQZVj2
Eplv2tfFhfeU9d2ocODWAxSFZ1Zw/u72iuPZvGVzsGqFgXOouL0b90yZ3p/ddVoLYhWB+bHot3bv
XgNl8iUJ/FKG1at26OW8VLmEyyBOGEXrOfsivZjEG2uwV1ddvGiiVia8wxXqAt8oAvLRKM3AAiVU
KO7EXDW0+O3DdsPDR0VpFRLCwYUrqEHW9n1k+nqR6rbxLGYu+z3pvvGhR7hYaIarT9V5gyt6Kn8s
FFbITXvgI+NFgYjlbQgXTXtIpOrXdA1bIGG+gX1jzjqB+JdWhnjH6zKTzGLszPl+jU5P11e4f7ge
vYaktnnaB3p2dc1oY26p+qNTX6eXfzKkOFMWBDpxHAFpp++92xyPX9MFOCZx2ZUFlX1XwxNiiU+G
LWt8Q7Y1qXsynTUO4PqXVCtmiDOsKZvQahb/ADLhhd6GP9sye9eyNDqkbOlHjpdIzrF40n/Bg0hZ
CJ7XaVELbiFvN0nyhzakeAjLku75X0bZHngqOXPYhbl2NeBOaxcMDS9LGYAicuF+RcfuX53ORl+T
b2g4R0AaNNRMORV+/xXL5vmSB8DNgb9H1YtuYFC1lGzBtLml8ZqnHKQXu+tuHnCzZ3XQCS8QySiy
TpH8w1vZGl/UuTTX6LwfCBGqcoj5Y6WUptCBPggasiH48+AXdK5NnSq7iodHoug36/Dr62w8FRSj
cwu0puTHWPfJeqIj/ahmVvqhLcQgDuuCtB6OH2VlqPrS0raoNSv07hYGuvgQorfSEq3cCSCaC+hG
X3mxDHNBPEe/EeD3YaS8IxJPBw9RmzjunWOYkXSxqa/mELfY6RrjgTy1YH4WqT2ieWfXQS2wjY+4
OGp9fJNZIXNWFzr8ksC4ERP5iE6xaQE1cQMRg9tgclxdBgTzfprmtKw9RvenYGaIjQ8UsSs/9BnT
BBzTIZmGpDxkK7abaPBnlkD99x9pgBIcqFkEBxYUF6EJi8gRJbJ/LzcDLA2YFwzxNwQuqoz7tBFu
ip2rKXb5oexFtz59/EP/fE5rz/vn2vsK/WQIFR/sCF5YQVqdNS+XW7z/BK+7VFo1/r9r0vg8vHjj
BGQJsJYY6rtXuJfX59JJv1AuITS8bbJaYuECNH4Z6bjVdZvJlQi/4XUNjj7xc/6NBfLO3D1fNErf
aumDr+LCCUEd4xgr3HbnTiC87nhZMmxlVzVgOaff7CBNmlWsNYZVkKwFlJ+3WsTYT5tU29Qo7wB4
aMlOK2Wo9fdmYSESTpc6WqogsKtP12PWAu8SjVafHOjy0AOC42C7A3NNk2l3YdvU27aPnudwoRnF
29OKLyZ6XEELc9goxuUyky6rw7o2dRMfyz09ZH87M8j5qVh4FXwvdcTqtUSdBS7CCIxt6apY9O2E
GnVifZi2iCYayUM1+SM64HpXpPT7S9yk+Odxhp0NatU1CBp5sdr4CWMExT3++iVNQTqkv/23aYiw
rzsIeuOlI/3H23C2ToX3q7KdJhxXD63TbRBXpCUXs4iuxjGXVLRv0A3/SKBCClEndI2F+KIrCnAB
/G/+I+PpXSRKJiFKgPJbmFv5zQKJxJL40s8v2b3fX+IcaRe9KM/P8dsOZqDBLF47SnVLrpRcwK9v
FIznXqlu69o9TgjkANPtOSmWU7H8Mde/ket3XJw+fGudtAClaEJoqpQPK8SXWvpVPhXE76S0amu6
A1/Usa/EsO7Upmdw4gsDpBMVKcqyvbK9ncKiyzvtZuRUc/zUBatXXw48U7nYdUrz8uArMcpT7Hfk
0Mz2c+nx2gM+yTMs2VYAlJQSSF4asaxRoeIeLNMon0S/nfob22RXA9DRdac+gaZn2ermMIEpWyoz
a2Bnj1cR+LUMshXt0+XO/kpH5bKBgRA7DsXzq/+DrRJPdG2m3Ne0lLWrHhCNPi5KZFXnQRihfjau
WO8zVjkd52rIxXHbr70Rxftlgsxy0biC/t5T0Wd6rIWDa7kgPkDI4nP0TaNAvlGOTGNkgeiFoEEK
aNN4OAKhI/mY0zP0itr55w5jiVaUKx2HK9SZi28qpg3a2LkyB6AAu8b0e0m3/HOwQB08doWgoFI7
X0Hkw6SG5Sh5j6TGwR8dXGK/clBTTJJRrl18kY0YSsIVu/Nqvnptawabt0KXTPIqeOl1QbI1CjSC
o5eplYJRC6BkKIYHu5NOygzzzYUwo1K0GB5AUG71UqALm/N9ke/Qj+mmRIPgAkmEEFS39pa0uRDj
P2SGqoP7F+nxQlKzONdvPvrcUNRfL7hiPhMZW6VnHdzfKQggnWE6Z0eGftG+d4/ocT+HIq9CaNQl
zbejzlYyiT28tnSQAGViZNHnHRaut3gt0VbIyT0aN/FO3TMPvBmVeef1E2kGW85cKEl5dDqzbuzn
C9vsmX0OAptpsG5Hu5yy3KPd86RK9zvCJO/p7zBuqggv0t2ylrv16IjTxMJsQxGDE+4kQWszJ53a
U3aUU3PIGLB89gSwo6S9jgJ4ndr4H54PRD6U1YUeV4r11fDynbrKYeO+i2OsjatSSZ0WM6AYBHtg
LnL9cFp/xvdwHUE182rlvjF+VMeRm+99r6npjxr9CpME/3o5t/Go/d4z303wj2Idhp1p+vez5KWh
cSbeQlPZTlRMfyjvi5BrJXDb+mofpmRMwd674j4IqpzRinRiHd4WVh14NdSZXcl/dimmrTdqo9gk
4KoAwvcguuBtRpJvnY135jQO2YM8cLLQnK2B4O3lhAiX5fASe0mVi0hJYt1nmQOQLzZvVi8xV2N0
fR6zB39931u/iZcDMYRlqevPEdKRMavypTffZWeaKuh00U0/7O3mPEkVDQP8ewVhJ/nGnRDkcD7V
VT0XpWy7eSgc1OkKeedUZdY0uTk//T22Tw3YEBc+yXBb3+egE10rDc1ncA3W3LHSv8NSpuah3qO/
bD6JNrUhzl+z7r4RaNk1D9bq6RsQlcoJfvkI/tlgxRwqbbVKs7Jgj32D0NPwEgNAyk6hDPmwGyrm
WO8wJ8yoj6xMGBItna0ZP6gLpEyCc7MaMLI06SrActhunkm9hiy0v/NlwCDah00KT7Jud6GYGzW/
GZdopPqvBY7lmooOMSfyqPHkHyrvX0WNy2Uro4x316ICpCIxHTLwZSKrhno8JGyK+ZI+f5kvWOY8
5eeg7Uean+C1xwymIPSPMf5pYj0MDl9DoM2lIrqm6q3XYDEbPbwF4z3nzYWoDeUr33DhnsKM89ka
dCr1c+qVIXmx/ErIaNCULLLvoks/cJbnIgQ2dCgachM75HJ6r4+XGiJixp2W/6nizbkVOP//tHUM
UfvVccxM7DylSjGYREBxn7DDmuwS8HYXFtBrEfdifjCyDhAprbztP4iU49Xk+N9+lSUPM53AaS6I
BpqLUW7VazKwVxSaHPcrSCT73um059qvvV+ZLPHsK0sPndbr7G/ySBklM43ZopEt8c1BftupJcYP
1HHsnqIiGPGt96ZYTG+hL0oekO2DpcXq4Syz929bNwlkjLfNMNAU37NRL2/krIyatMGTgiiuS2he
8jJybW1chbZ/P9w1FQGvC5BwswCKIWFmx+Sgv1lMT7BnF6gu8gBndLFhLh5lPI77KLCTEf96mnFr
kx5vwDzh19IWA2OTcsykapxtHELJoHaKkvEUG2rejxUooORNbuqs3daL5QxFELQyNHyad1gAc9Zl
gES66oo35X4XCJbK0Cg/XYN7KIOjXKvZsPj5eeNMUo6xp9f7ID1UnYnzBjFjjyec2acYR3RvUGeZ
NCmtEo5aSheTg2sycuTphZiYuFBVkIGT4LKmEehsvnQ7V1x5FLsrd6dKxt9VbwNHrop0hKoX1Ex9
wsfIDoZ4srFQHKVbtmA9OeMC/9F03nnzQSAFl/AptFAPCNLPDcmI49COJZM4fBf0wXH1xm8NaABc
oGmgBoYPcIMrdpHmklCQoBzxvosRwLsWXlpbn995zzUxJcCVXy7RljQiEroJ+GqJJo1mgfQfnJiV
7S5RnNnQ4lWqSfjOmMBnAuCHaB0Vh8V5QS99u+DWaJ/7c/ZeuZM/3vd5kMMz1bWIryL1V0nuIaCk
2ywGwOre3N2wyfnYmk/FkhnBRCbTGajBQxJwF3qibaDvJyLyIY/Yc4LI8ei79w97sH9u4IVHY/er
qXSsOKDFyrcdaXkrzkUr6JKjV+t8BEbG83Scmdvl9W5BgudN5Cf2tV/sg7oefJdHkbvB387roun4
YVeA/sJ2B8IxtcmO1Ct/aq59ifSZ7F9IsvVIZaQ9EIAcF6Yjc9bq3Aa3joI9m2NIQXUp7sHcfKly
+ErJoCHW8YqI1HZuX3ghNr3nwo4FhMhuXXPzDYUERNCFZb5hW+dQ+jdCihi19Uwnc4jHObbOjnSv
plPkV6q7dIMJyVyD5xdKBUnRhaPVbHzqM+TRQTJaXyAwvBZqkSqFQ7JpgueCdM6dNXMsYFbmvE3N
VeX94XP8fR0uNk4yel222lScDB2lq+pwXHnqMKOkWmRG72Kmh2YR7DCDrLLoxlcrwqQ1jx6KCGg+
97m2WWByuue4q8PIj+Yw+uo1nB8gZIsP2OFFnR9ukfuBX2pCw2K2UNKFgoTXXUk/hP6alvSPNbJf
+7PnR+6hi2QYXjxMPvTK6xWvC1Wad0d4EDL/Bxzoa011pPLj5RcqQd6nTOi2Z/akYmm5j0nXJdf7
9PvaJEM9Kb73sPrcp09Yp2QbJeLqEa0Fofa6yjEa0JjT84nz/jBhKryFuwmiNswCSNbRffvN5aOd
Ru01cYKj0CfC4qw8Ebj1YxnejWowjzoYSaeC+SRsmqynfCRIzuN4YfudLNsMPSKiwSlDqIVZxRjx
azMOXwI3+4DKpXJRrbRwbq/qrFFO2ROH/z4YF4/2AQDYnZDk771i3obK/SIPz3PupWbxmtb8dR3+
tj/CbdKbj2S/4J4mnAZH81YmKfbxI6AHlUSmVt7zqmnkRKwd2y4Gs6VgHYndWAgcb5CEiADI0Uj9
lLdYIDu+GLa1BBF8qVzJp5yqzC83JbjvJ5ju2ytOp8dMrZiSdHOcKN+pgQERsYoQ1osG9yOzBNO1
DdUYnp1NcheKt+N0io9ek8/1SVE9Nps2u3W2CfhRhre+Lgm0cOIfvhMx5fAojBB6mconjw+XhRnL
Srm43RLK01pqk/4Zr6V+tKM5o1IE+hElXZMWga/bumPEmddcR1YB1uSC1D7G6H/fU41hgm89mZUZ
xSxZAwg6q0ez/2y8c+w5LMuP+AWmPYvnmo8nfM8bPutId7w2Z3RzWCntzSuqVGPqwTrI+hCdVrBz
KSkWauxr+yeDpyV9xmXFg5qT/NU8j5ZFh4rCMcAIVkG57ePyqJdrUOrFSJmnoJP59y8FD8qy1Cdq
2k/z1ejLkIvkriTqxY+u1yl7jjTPdhdwAuUjBSvQeRU+JCuecKRNCcVMBFI2ls94xKQVzxMPc5r9
qtJS4JQgDwP7625e+VrCLw53nPD/bysRunx7FkIdUraTei+r29FYpZ97B015bt5XQKRf7bh4cavS
F6VKBhMmb2r6nW9QckUTN2OaGT2OOattVYxHO6JpPbEk6Ypd5oWm/MrMM2wbg+DnkUbHX4Sk8zn4
j0GZu+Am5Z1Kyhl1u+42Ydr1QW/Y04Wyw2+ALGxgCQQeIaAPY7elFA8BsWtEfssBeNbu7ZQE1+Gb
1lbFtEtzyYGcO+mq4+WWxyMBYclby66+6p1tMuHr+9vAvJb7GoJ00p3uWJ+S9/KxTMKMNuZGU+zB
KGjmFQeVHnlIMuTeos4A/32gmnR7hB6XvlXdhpSJoFph9Ucq14Im8NgTME9FEfJT/jSWhS3vUdSn
NUKaupSPLJF57nD/R1yoXKizdrHHWe6f88pQLWzqr7Xzk6sYuAeG9WRGSYw3g/HP6SLeweNDy5i1
KSiLS7Cxr4vnd9MfVXx7f8pW+TTPfkxmaMz2pyDXHTGN3AnL9IIZchqSS2P/1jMMFobg8zomrJB6
QJDifXRzev319gZFVHd5N5hqTE/ajO3gJEde/jIMw6Kc2pl8tWJNZEH6X4uQOSjYhg8U1reIIlRe
ZFX4x4PwHras5XEQtVqCK5Cl8nC1XjO4ODDnvdeaQQFzQdXkR+EEb20GDMZgKstFThCYS03wd1OX
A/K+lcka1uMT96J7Ha9VGe3Nb0qUzWx1eiIbM8kkDsp7Vk3c1gC4OBIiONXxEg3bjZNXzw6LI5GJ
Px9mh6+bUk01ZbDHYuMkqp5WnUI0dtFCYthyTbq7rmRn93liI0Xus+2EWLcdhyGAmILQPfa5bWaO
+MNKQe2aHPz9bTkJcUlxUfiFF8frGhNGIMjlhbm+7S+SPQB3TRIi3NOAv6j3jwvpCUpNuFZXGkHA
g2MdmZ1STWINjh9uxH6hZArIHMzV2HeLUypGimtvoGq1un6CIdAqyegyrMfL3pEpTH5hzjqNdTsr
GrL9b8Shiy5UZuFWp8MLUQbr0ylBJKuYQxYb8SuarMV84xLgZaaK0OSm6sNa0m5y9km0QpWsYACD
k2+ZVxKpezXlKBBQFSSxLa2+fCZR87skGKikRunpMeHtGE7Biqn6eZY3cD3/mkwV0mofsW5nNiOs
n9fiIs3iUjHfrrp2QnmIJjYBSTDKO/ntPNP5TweXQ9OHtRYqrRNRzzSYOBriWtP8szTNbuxf8p9Y
CtnPDhYl8ZqPL+Tmq4RI/Vi93kKSUK9jJM6LrFQ9NusuZKXFqn0KWN9XLgozzyTDyd8+jPTCMCXr
qF8m3lhtyIO0qtF4GE4L5KvaK/+ZdIvLeZEcixuTjAQayDCs47nMubmgh0IcOmvtlYdtBccFmFIB
XfmajG0UDJ8AA4YSYgSA0KJ7sVFv9tUIRUt3y1iQUeOioLJ85rHCQr+SBZI9OJ1DplyZlaBjF+z8
J+YGKKj+AZh8G/A1tweJ+1XAehDH3JRCmw8W4i9bGmOLyDHV6sDX7zhPVEu5u0eY3bE5QROJKMnr
I3/ySb9CqpTZVtWYlmNSxXqCMn2Gk5uoQwpXYEcOLdR8JaS/ZJ/SmHudo+0FgYoEeooA+GBNDyuI
/yaDf/O7KQX+zCbx1h+ESLqxsOtBD2veu2NwFeakzRDzWfKGKG2OOp/VeokZ/QKc13BygqbjtO8z
1vtVXmHNqIJpRZsqS7HwO66nNfEECecHJiyyx1bhXFHF32jtBE9UVuB8xj1ljQswqqwlLcWQ3kcp
cFjRP1JRd5FSIw1J3GO8KVuSx4T0LrnJT0GJOCAwtJA79n762wW3wEFxmRcscMBJqHZTjFpHd9jT
T80pnpB8phR/Eok5D+Br4dqBRmvdak958D0RaicKQmcBi3SxQacEJzFJ9GhYC9evIJ/fSxkIuZuO
daaGJ40emoOU/SwmIFc5A+w0cNAhyuBF8x+HMRBZOpCDUyNyHuRJQi+FP9n5/3ceOA6J6yhrUTi7
QI6HvK08jRpyfUhT4AVBjE24AHfljLl12TSRIB6DbgKDQcEYABEELK+QzWBFZlL1N9y9VLo4NULs
fseqeGcAUkBdqL4khSK5mpiwhHHpP269ZD4kamzL0Q4iIIxe0Bust9OuQF1YH77sEscLh9cEI6Mc
MahcSpRrLerpFO+ms+zZEiZn7wNYVQe2OTi9tlK5eQ//n/kwZjg+U9Bl1lJXUKtRr0nLRM/rgohL
6iwL7pm1DB5rDOsP8zeW5gkHaS5+b1agVfbgkKsdV7tWHkBJAd1JvMCkE9pf1JkXc0YM9kbBHgIT
gHyE8V+m3tQSshxqWiRryRzSmlGHof88OLuNfp5F9s7yNislY0Ok38B1lDHGo4gU55TPB9Aw1JuS
UoxisMSahb/7azq3BoRXVmbAo6lH6798VahQ8iPpWvII1cwagUPEDOuiBzTYuDusWi/K7QOZ58UW
D3SQLXv1zsn99jYpzmoRpq5mM5d54PxU9fMWS6k/n7mkepYOrHh4kBVKJfUi9cbY/U9L37T+Hbb+
Hb2nRMH5uv5KORuo3iciO09yO8qZbIkGzMsEjUueKoHxibSdQoBpPm9MIEN/qKv7InNZRc8Vbp0A
4THCTO5ZZ1T4iVLg8WQrVo8M9DRHT61dtQCku2e6wFTOig9VFaXnJ+wpPUUJJCBpkHEs5AoVPG4e
+UziI5Kwb5jCFIZsGBKgUuoFwIjOLZqbNJw5qAMxU3ewRbS6hTX+f1e0OQvrTWXIokGzR7xcXxsM
P7aZUzg4FUrjX4CZLfaGTjjarPZ2/n4FDt3FMwezjqlFsP7w6eGaZNRc7Pc1oQLeTScTcHtYClYr
6LHic27H/Ir/mxV8kJLggpm0XbwzSvOjU36sTlO/PLifIufesFQpUzTE6af/DF5/kMIkCumKX14z
vyCIA1ZvpSqhvi7pLe2Dpn6J90hgypl4Pj/e1XNYXhZeps/UDqalQKx6uSd61IGYu71T0kDKSQGL
ThTq/G1FBFqHrupV91NeFeMopqoQs65v0+cC9NSwRgKmXV/KEJmgv5pnfi4bMJoEnWfgyg0THtvy
QCdr3M8ZfEHW1nukPpmhu6is8HrhV6H1+L+Jv8LtUnTW7bYCwc+EUaAxbUOHNyPxpMYhM8j+kSnu
+eNibxCxxx8qbhuczfKVUdV8eqhAi2LL/IXbgMSv9gKKVY1ignMUup5IfEAzhhnak7zW2FiroJYC
Qqq7yxsz5jGwIi7I9EzpVrOXN4MMcdblq4TH+oBS8fn98LZyFwecx6WQUxnFUHdXNYJ+WAspQ4Tj
0AcE+SGTSyGdu66Ew6ToWpDmLP4/ptr4IS1yhLvI/iTa+LPgGjAmbnk/Hx29n1s4kMXDs9z2LPjp
he70YegRc4Ym+n9mII0t775gGK/NwVndxEluK9km3e04Xv8K+ZS8aWD/PuzgQaXqgdCFdJO1Vl6P
rpGy+941XL+4WYrkJIIclJ6+3ApNRlchWVc3P6I+1mRL3seQ6hFTg+dfIsFV2VM7SuzTLEvY3Cf5
dGXYQtuRILwn8K6D0eHSZDJCYB7xhi8YkcDt1g7SsR9qIOW/nmcvi9Zut1LyNuB6JkrO1flYaerr
ec9gJO63/8MIvi085u06PKYaljIaKp39lEzQ1AnAk/FBStKmU6h6aZjLz46Eq3Tiwcwj5q8yOl/H
bka7v++1jcGPJKFjD6xSDW/lzo32jk5TAOHeUkR0AkzdC8kmTHFaMXzqGsCgDX+tD7JrrNrYSBPo
unMypVN6fWsvOkhNfxuQc1ElIqieoPlbSnPt/c7uJLwOh7ius/RGyIKG+ssTzsPstkoKEcC7/Fd3
Ju9rjVeL9409kQIA6h5H7uNBBExd7zKH077LABTlK7r2T1hMH1TStr2fJOlHpEGzJjeJ2T3Gq7u8
NtWChs8yajA7dbD6ptuJYUsuhXUnXan4lZMjohsSQYsQ62czWNjOcQ+1OaXZGl2riQeHSKtF0qVt
MH9RvfAxekvzNRq3BsX42vV3BjiXlxGcmBfaH0auRXODJwIuXe5y7w67JngkOdU6l0shJ3p/277S
tUThYHFg2rWnGuCa3CiYUAjfUeZitxo6paicKTmJ7huvaCetXDL67/a9HKfzt4Zw74VT2/Xo4YBZ
S6kjNcR7dLebpOPhwvVVaBERUZcnDdQOm+Ld5BBo0DMhGT8pE3ks7qW1uf5qacud2UUDFXGy+L+J
c5FlY0bF5+58W/557RjdRa36HxAP3rV6G9ADGzpJE6rlYuEDnL2bFGRRPDL0+PUQVvVz2hy0lNq+
3nKzAfbqcXg+X69rR5Dwq3kwGxwGk7Pju+06fyOg7AYEy7nJRxYOLL2ohAfZLjXWo6EpiuZqnTCF
Utj/+H5ueuguSs0KAJKXwmJpyT9U4uQN4S9UgvCOj3Kp/5b5nFlagHqXAIP3t029dEqAn9Jw4Cg2
UPm+E/SLuNgfcxkJegnZAVrX7pa09GU/gmiy6L46NBoDO39s3DyNVHY40AnhxADZRkN/oh7p20Cd
0GxNpjylxRiP0O3NNMd3apMHKrh3NWXml4OWnrDG/kbXbIVvJKPhl80qHp1Fy9yzMLGAt5ydHWAn
8moCcqvuQ30R9J7dBP0K72eN/TKa8uVh2GjOtCLNp2L+80Ro5S44C4br0P2GdUWnzSqS6E2U4xTD
GPwgiBu/v2Ht+e/HuXdrMREkANZu1Hv2e9CZSCrb71zPsuEExbUnzZsrWxX8jp2KX6WUs7kToXzm
uKgxyY4BegK1BCNAO5fWvJDk8reILSAuOZMGE14kI6HOq+2tZjlD2CSBXyaJQ4UJ+QsUTdIOXpdK
x0SY6LrXkH2k+UDMOQSn42Nzb80aFetoLdXGW25WMYDYlrs45ZgqoHgbwMXMaFRHZFSEjXEjxxHO
uxh3rk6TE9rlu61QwyeJBu5A32NtiZFW4RmD23/2Nft+Oka6BFwb7DN2Uih24/qJ6XiXjDSQgG+S
R3n92cSRIvBb80cwYtCxb6/rOrhwj/V/ActqLRef/mi+SkrfP1CaGGEJN1FiKyPOk5ahxySxrqWF
JIJIJs3RW5qds3zJ8nAUKT53gvbT5j8O1ihmgrbtPS0RMqibcP4BBUs/D+rvJrp+DmaGOEXaKjp0
XCXAuWu79hi4Z14xY59lI7Pjl8wax3dsT95mMR9VrC/qZpPLYtvs+Lzd1wmQjwpBi5uI91lUPbtE
Rc1w0aOQapgOjTH2bRZ4JLjXdataf31SQWG6wRG6KktwBefmhy8gq4+daxt3WukNiya4lMDZO7yl
XdvLBdpQ1bWlNDjnKGno+5OXGMg2GfVDkTwLFtlpeDAc89MVp/X076nLHQoE/Rw8m64Zz/kB90ou
/X6cMVbe00NbYv/1vA84vhlz1xNvsoIRccjmVINZ/xkjDzOAeCKy7inL993Df/STXgFaFvG8zPPq
t1zliEAAE54Rk2DUxqVbKc0NKHRAhVq3QjXrU1yx3m6jWypV5mbY1Cm5GexMMdlyisPNZqiPv7n/
JVv3vBVnF4IcsuEP6c//PH5E1wpEvem4pTxdWL5w+mm9HT5VU1ukLdczAM3NfUn+RGGbi57hLMKy
61CEgSK0+MvYL8wEi+u82cDXcN03thT0LJd68wuO8yhQz1HWqp9CZz5/Hfj0E22QKV4+tOfXSvSe
tJnfO95UqhKuAY2UFdQUHueWEfhfd89cjpWXQ6dcuxjBR1tTP3SBLVD1dVxxFLdwGYoZy+YySKyo
p6DautQbOWUK8ysQuXX63GmLCDf2SntqcQjfVoYjy+nr1+T/VoVXqBpDGtrk/PJowqhWhHsjPU1S
ZdIwJ06gncVu7/gY08sLQle3e7NG4MYnbZ8Oh7DLedjfsCfamqbSqcteQdRahMqCA6/878f8rn+S
b7ANwIqAiQ5TYLdBueydunMTeYo72ayfxCT9bj4W/8lUdAbyx8TqYINYxeJugDx/IzCYDJa7dezz
Rqp4iF9FDbqj1mYxDKc+zfvf3bCmDwZOZne4949XItBcVci1kS15/arw1W/VoHwdb5TWN4ynoQgF
YLgIfEUVx5YUyRWjPI6Sg6R4uPw5zIx34DLb4ANOlvSRzMlpr8EDmDgzlOIE86TAn6HXFE6zxmCO
JiAXmwwl7CTaCAMLzyeXTwI3foHfOqdxU9jOJkahkNYWLtZR0BKVVyZeQtgV66D4VHlCSB7/N/XQ
GCrl3Zlva64/apmYgb96tdUQI67/5CWPQWoOJ6ZmlU9X2H0JPefz+TwkjcB5X1iZaw3ek+e1jeVK
cQemFEMKajw8KRsRs2bBIkSfwEy+1ss+44urA+QtzgXkZ2A9xcfp5FLLRRkezKWvz+lD4T2/uYBs
OvqEwUSKbdn4VP/pBmwwfdHJ2/VaKyJLEE4M51oiv04Oiqabtp2QNiH6xB2RVveWplhglyxYyVHC
nm/43uIjrzsniB3hn1zgZqmIv3lUo+akpK2Bgs1p1HObKuZR71i+RdxvmSnQVAf2lY4t2M/NhXgp
UhyQBjP2V4nJssHKl7BVpDuD+sy6zdULmY/pw9ZI5GXLeYb+TyRK3qik7oj7+sdW+10JRZR09Rml
bs61kEluY6hj431phfI9pXupeYTBxWQL+FDDOhkHd1uaHkawKHgtb26OaRDZMEHp8udN/ta7LbZY
6tzzlB22AtysQY3opmT+XoPbCHjKAirqfOXqoMMV/2ENMFRHX7aPA3DH+Wzyhux+gHDJ70KeNVr2
QyMZDArz3z3u3FoD0Zpy9CNE2LsAXAm7y2gZq07uPBH0e58jTeu42XpgN1Js8xVXf5E6itK6ZR8T
ketD529s1bp6cAmIYIzGRPwuopGGonwOk9mTckcBVBD1C3D2MK8lmiTk1sWIJw63DZu0WOyxdd4D
J6L2luNk+ucG5hHPYR7PrSPBVfovgwFDvpEXbfl7b5kBSGMRADVE1dW5XzNwAi5/LRHwGsCTlcey
hjGuo7f9C6s5SU+SO8Dh9iUOeUpZSQw7E+iEx2pFbyep7hLizVEnJV6ia4guHmk9PR64NgGh5tAv
3SZxGH/wdb+RXnqFnnIDL5McDL8txhygHho7laqt8605o7OsBVY7am9LExACitHBor8BhArAtLuW
iHpu/dOt3J6ebYpxu0hi3w/YGIOnqnX8e3XWltU+4jNwP4323e9rSK2S5Ge10gct6KoL7a3co7zn
Kbqfv+TbUkoDlzvdmi9YznhGUkYDlEuH/jw7GVTgbxeouv8PbiGDRiZdG4g9l7z4sbZkFpcNiBvr
gxEuneTKv8yLIShFcQ/bTJ0X+lZvKWtIL9kBIs6Uahzkm/u5r+QFzeniIH3eAlUg4Yn1uaKJEflm
h31T+6s1f/DA3XIZqjjToY2tIH2HFcnPc3Pg4PC1X5ncR/wbak2c7SqaFp5PlYIqQgM24Kg2k6Q9
BKRRE0XXcvAw/RhqQzkhjbQbsyUhk+agz/WhD5fah+IMiF6pdv9lrLYC88MMDntpJOXoSwAvoZSd
/0beWQ2d7DjPEkxdiTC5XWiAczLL+cAXPa/YSCIETtYGsjSkhrOvF+lr/r+4oOiV+jlW5mkkTIsK
wTXC1Os0khGPiRZzaGY34VNRyNzihWRIGzkpWu02ZKJB7hgRhjqfAC+xXNYxsEjQKs/jhiu6LfBI
oCjpG1LerHBxJ3Gh6Pq0vVs3DpOFCIy7Pj7NuS/MZ2BnLCyFWVGlcMKz6PLiXhopBWP6AKzYtTZA
RypG9utB3B2wvd2yiCjoFNcynnk5LpcQHLK0tBD+uutaWudiH+GfK/opNxn1NcAMMkGPZ4Wra/5c
bztva4y0RtEo6c3/ayAAMf9CV3bILbzcqLq6A5Oa2hNFBSkNSun30MN9LQMoYAtzIIOpjKumghmZ
ILhnqQpzDM60URbGk6bZYiZMLwiGQnYzoszGjHqSMrovBALSwoy8+fCD3zzLlFEtTqNncmNtvTJk
70LdNXkqp9R6uE2oVxBxArvZQ6AV7Opn+84Slyy1NQFeHV7k0qJOVBgShFEVqGlBlhJX8RilUXdD
S28sPm7E2VKsTumw/y4zHprFgFBUGrZmaf2cGrvgLH2bLrkW4j5yqqRywCnm5j93LpGVPDm7Sz+Y
a8egxhK7SKVBwzt9XnO+oixY23BVZ0O2ZrVL6lkfQcMH/LnbkMxglwu08jdvaYvFK9M3kwz7yZB2
Dk9PfGwKQfj7qMeJ9zDfPVtAkyU9rjJGF/4oledVDDRBk1raCopa33UlgTi+VoK4tdqW4L4xojTH
BfO+0ux2K9GxFHa6rfFPBAJhfB5WlrmQrZ9jyRj4c1uORAAh1ryW4CgrclZg88oV1txMiBxTICGf
68wq73jNNGKyUhzgUlKV8+tweHz//eXPku7upwMNtMMFEnoHo3a82JW7f7Zap07ON8TqkD3usmOa
FcS0ZYziDg2W+mo2dH35beGkNWu4JZ83yjJZYWhJmgxUFj7Ptf3aOFEJ7HbcBe0729w27lK8mDgu
jP1LehVGAzLUklQ/U3BU7R0zDwCBblouQ/XF4G7Sr6NO9jRuMWWFhEE1Xp6pYtV+J+/0eHMDQtMM
/6LE21Ndq0KaMA2gpp/o011TTp8e67L8F3XEPUBIN6gjbIIlP9IMazfo70ysvqKhhZOeDMVDUN+E
onu/3qP+a6SXI46W/DMKHimTRMW/ARkMEhoTlkIMTF4eZo6XMeWvS1w/IfIwAo2Ezi9PnZQuf5Md
hd3Ahx5d2wSJexcsfjEkUkvb0TZCPBOQnYVwiiPEGhYGVVTtrQzU+R9+PxVnm0oYFN+xizujXGKv
EYkJ3ve1sW/lqRjEY/PxYlAEVcwwmMVneQDocRjCE20Q6KrQ6HWE9bhnsCsVhXzxuVAwgqi6AMr2
xbMQWAA657TSw9dL08WOg0ui9G0iSjWhpWW04UGf1HUgCh651B1iqLF8BtpxJXktv40grLUa3Z6K
ssAi0DCe0XlC/SPNKk0WmJf8xcVgvyHzULULG9Xjv2oIPtu0DKuwHBWug8nsT/Gca4YSR6RFLQX7
gdCzIZFbSn4uhypHy58lq8f+yq6SHY/2G9XFGXthbtPP23BFv4GNktDIcY3vk4El0Spy6VYGCqEw
zr0iJwKArJzZM6k+xSRU7CpCU/ZRItbZXmFNk+jcQ8tOh3cibxD0ShHBD3dkHSYJfdTID1CMU6gK
yPeLDTRI7M63KSRM91Y9kXDjHcFwmB4daLYwHQYHIuzVHDSEmOw6amjSxrIs6Bw7x1e/lmG6xK7m
QbuMbekTYVnFk/1brpPGMZ1NsSwhmRty76+abGPFBzU+XSy6IJdD0TODuc7s4kd1BtR/vGPeT5Xe
dajb+0bRt4gmxJtJJ6wvb0R8Osux7x/4iRqLhd6KGX5/5Is+E2CUGrJCcVmkNLbZPhNNGscDGGLz
cAdmh45b9pAgJ1+1qSjXDw0UPsdrCKmTFn8/E9QB16xd+lU4bnGMs1ATbOEEhzuirKYeFdGT/G0o
8pyupI2oW3gAdBkU97ka2XrT/CcSqF0zmppsqD9eBYAmaJDdHn1xaf9kHLoIXO1KAxk/d5Xb6VNa
B6EraRTkHdHWl+oEKQzNTfvBmdbjLW6Aay+Ff3KhlI9pS8NBrfQlH1FaeIrU7AyajxUBIJgqWMqm
iiPwDWqio5oLwUiWl6kxhcDy/37F5lxV4VmjMx8TAslqc1EzarSwW77vEOoj9phVUSK9MxxXSTcZ
+B9GTlnBv0j+6boxuvUijA7jndXd4fwwY7PX65eiXL3KiFoaNCRq147lVfPcOUgki5rZptReMtbs
7N7XqU3sc4YBelltFtPIVXQTMDFsTTobaBEcGUZKGUPI4OA5gOctGxL/27tfNoCsljHDKvjqIhLY
7/bxsv/KNa+bGCSLLjNVohaObMGASE9TY3RlN3SQzvVmYHRONq6Ka7IBYCV5KWXtiHLRsZRiK1QX
6Wziw9NMhe72I3kaH7lRAVG6A3g5Jz/7j85ica17s2K/sJReFfuDpigG9O8mRrlSNdwypmZDntqe
SEYMtFPg/6PZwRfnuBD0ATZOqoDLVOhfJefXnXH2AhNxIR154fQR6ZaOGeJ/GT1qa8DgLv5V+1GN
GeQCxX0MBfb/PfBi7I7ze8KQwBN451GS2ffJ2Mydypa7nKrnUuCgzKhV53Qde/UXZOJLd16dYMgA
K2J0Qpe+bD6+mIRf9RAKXmQFmyEEsQi1AR9wNC/S3ZgSXyeXU6NnXUeiyf/kx0Id3OTIkVOkfDMc
/EavldUZBtcJumsmTwfu2DTG0WeZ4VAk4XgUqMseELWpx76H1a1hhFMZ4oqrzjGD4WoVNRYnInBz
k0vcIRm/moXTpdUdklKsA2qoMV+P4UaK9yhlAcRr3BthJPcEf8dQ+lL0cSV4Q8qISdpUB35yntuJ
tXrIq+Ar37jGn0li3iOCDix3E2bgtxhubbiRjaVwVnOwDo4X3KIp5Q2wzlBdTXjLNj02DNnxwc5F
n4HjsqqFelgM6qEtiCPfS0Jx8H1kKbVXPvHD3p7p07JGT82+zyUXWDWjG3wxHbIErGPvcjak+16W
JFCu4GXDBO/HWfCr7MgDvbMcCQd5KhKkxvg0LPxiAIHDFRFayOsXATEkcY8qIJ2smy2fMm7nPdUm
O8F+KbQ+M8f8LlYbxbrw8iBkRhO1ZYRil4xPzfZ6XSCgC4p+3+eNx844s9fqH7tpdCKsfQayBJhV
CVP5TP1DzfqXeiauJs8A/WmE+D4KCTp6rOq+RXDTXnGzd4k8JPwoOdGEcZSPz/AlNlh6hWfnv+gG
Bz2PjF7944/J4lSwBvNsFMiaAo8iAQghlGhgyFPd9U4Q0TeFfpQ5FRmRJFvENiX4cHHLYoQPHnVp
Izi1AI2mJBSAZdIaAqfs1BBJC3llmfud3gVbA7oaeShgm6+IyX2hpNR+uHQqY7RT5wpR6REJsNcx
OdHJm5gr11xsoemJKQQ3XuS9OP9kNn+Ix398O7nT8jfUaY/lGL4sYrNrCn2z2673lYLHyrv3c0pj
QCnahATHOtC2szL/gjTsUNRgydL/NA0sp0t/Hq2QfEW8pJvZPznxwT2+GASu7AjMtl6jXGgDgFys
lQwHE9QrJwT9pXt1325XCpdeOjR1xADz2kFvauj16G5DGtlvWw2XXjiECe2Tys5KSbIpR9/istp/
QV3QWS89usyP+Fvp3P7yJ6iH1Z/yFS3EypwpGy5aL3Dko09cRD4Uz6Beq5X8iFZO/ouWd5DN2D2/
maoAGRNqVn/ZxED1NdudbOMTGshfVS2Sn744ml+9/ErCI0r+yXqjJU73F3LlDhjpkRO5CLxjCTRg
IYSCt2l/UQHscz24mCauugIY0PQJxO78DT9nFqRKG99rNSkygLJWFEXozi8VKC1rINP5GgcK7vAX
1RreQnf3FTUr1qB2cz7Zk7PgxR6rR33lKCARQbiW1TUneaByvfVkSnQWhE+WFqo+8k+JgjGBEw3D
pOQyUJTXzQDiMUn+O2P0oJVF1dz0JjbtHZapvpXAK7PgJbzcWgRfRQ1Pzmusz1sJXRQC46BJ4JHt
dF5EOU4eA9/g03xNmTMWE3xVG8ZT7XXrTcIbeIPXHkoNlxgJ7XwIsMc62/UNJYZrq1XZNLBR/MvO
yQeAe7ZXaFqLYm6Ir/6XOkctilBW43wd6hpxc4Cyw+OKAGPv/L/sdby+BhwsBjyub/Dfs25VE/JO
I9bWdJ15/VZ1yBrwqQpe4a8kblXdFhm4xxja2yAhU+kkLQWyS132FVeufooz8AUbbsiMP9CeL2A+
QnP/+92ew+D6Cy112ERScr9YZdMUbtukjf1amIIPgJkw3fJRjRiRA8NPuHtmLF3ISpAHT+8gZRg5
KLgZkb6Fs3ig5E5zgWSjCQEBD1rehGNAtg9Rh7gCcPhJQrltcI/swQAa00jEIVZ/Ma8IRWAihas0
cOEB8q+9Gexh4vM/N1D3iCZ+J3Vih9RLGgd3ztttAlhA3OXeQ6UTmqeqXFJczov0Z5Mw5falWUlz
mjZxM4bSYCoLDF/avPPGy3eNC03GT3AfpBtvN/oKvbj8rYmXbKutpcFRaGsSUcNxS7lWQNlcY52B
7UA0tR019t5lX6wk8YOqV4wotOC68hBn64zpGp/gD7XyiZ/z/uRu4pIeSTfP9QKUxjsvLWcxukzD
IBipM5L6t1EWDhkXSDZqZg1gVPWjD32cPWrl1YabEyDoxgwC293Lh2jwcP6xy2sFIfBSDCl45KVc
YIcBRk/KGuwZxM/DnldZRDRnNDIzu/MuKZ2abJqWdsVAQW6VFggIlNh+CCPfe3lRELSSW5oa04b3
KUj2uskJItRyiyklVEnAiF6IAAr0f8yrZMyKWLE/OKbKXBX9pf32b31wOJklcayvRU9GyZdVXlgb
fkzZsnoAZwZ6jbvAcrrfATOvrkbhI3zRRAOsVbhBukY4GF5tVoBIXe9NDwr3fOC/9ATLa322t7lz
0NCKLiDxL47Ogx8Z08S5y2z1ON2aubx1r2azGWyFpiJmV2tGVkDu6R7IzYKVtNINaNQa3A1UfKtS
hwOS12VCPBS7yl3J1B3AicxilOilNMT+W3Mj0cn2eshhKIBPUCWyYygJD5iUORmosEKuNhlP/o1/
F0r8fykIzRht9n0fq1duzicSTBP/zV5B6nrnCcLsa38T93dilLVBUT75185/w3DGlPRxfgptzw4z
GBZP8sw4TeM0CHNQpABb83Kr29Qqp1QhjKuNdMUSxxVW7n3PmBRPV+7b8GSJ+K7AJ0FdkGvJy9Ai
veGMqagUFbYW6nc9vX6Z+5n9hYsRzSZGWS/R/kKX00NclXKCQCke0R4O7/F2l1MxUlUHRioxYhLf
SSVumkqJ7veTbq6G3Lz9S76CCvdKODLqkrkobvDbzgHPJlBScWnacFx4JMIZrrJ0qkmy8346t/Kp
EL8DBJf/MOXte/TSQI0UnLGKaHUHPgMBRUnxNhTdevM5kuy+4yW4ql7Cqpc1zyiGjp6F2BNmhdFf
GiAte99FluIR+O/GGG3VjJvi2o4YoE55x4HykqARg+J3tSAje9uFdWCWG3KNqV9CrJghRusrVFej
PhbrbUxKCn/lJD4os35lbqA9rbZTttSVIjhOfGvXYFY2efolJSAz35EcRNBRVrwwboKSNQHcpYpV
VookNy8rMUdGbfLvuiQzu4p7k9dpnisWrLbhx+TmoAFb32HhyeNzeqwZLQ4AvbXnyvok7jDibI3W
a4CDtCE2LemQhC397legxb2LFh3Z4KwbJ9pV6hQgsDIJs+4Wa3mZJB1lZ9PmDbiwTKTlipvmDKVf
Ucgn1aQiscyT/DCvBQy0MyycyEMc1sii298VBlauyhQvI1aup64Jlj8pVbwzL1tPHypb3lVlBuko
6X7/6Tj0mhEFHoacLK10J2O2LtrhrMIgXtDIrfOWVsgvaQO52v3BL3drSAhi45H6v9r0DMTUbOuw
1DzD5AiMadE3gAcoJ/Xz0SutM4JeQy9Kf6LB3YS2oF0wNtBSWH1VsWmxoRc0182wFW/dlSume6xk
tby6mRdiBRrnssjR53kPjIPsrLA7SuB+qFS0S/V+SpJ8PBuRLbQ/XuD342PdrjKJeEexZ4U+m9v6
0XJxDeGFuQZACne0n9j4tZZvriwYfIo08qKPdhHkR4wTQ7IDUbYoWFmE7AF2Tv07VvDC8lJQ+i1B
B2CbbAbKElYxzeEtBj4QPtDEyfWZYOX8XRdZHaU747gpgdzgNSbEeH9LBIJcePKeb9lur8UC5wDg
GC4w5GNNwLLnvYjYWZiFlh0gXH6M7lQYVZOZ1utegXuvMzUDbnM7lR3qcAuj9kK5/hQjAzktLOwT
XlpiR3VXYfuuEEzCnZWtErP2YGQ7PSE3SXuZQsEdMmGOy5Yeva9ybZcd46cM1qP7Hx+6j61NERc0
w+36CR92IGCVIKoZ1gCYgfS+3JXsOZOVRmy5Y23A3HlxQCwhfr6lTq8y4lyWcz537Xohc7vTX74j
Icteq9yk1dMqE61PqqtwcKLdm8zYwqiS1+sL2VD67kGg85xESnIRahSM0qJXoOXxfp6HGRJq0kkl
CufiH33r7Jf+Yko9CA7JcRgxkVmInC2rO81rOnXDysRzsd8J233cle1uYq+3CIL4czKljyJ2Xm6g
4xLtw4e+8UPyKUP5C/I1ddUhhop8d0S9AGXugZTkmFWh6CMP90TFVcQzwGketIye0TDMMxd/fNMc
ZiLvtQnE+hbSp3xp3UbRYjolZSBZ45mDdC3Q0nXACZDOyTUMpbfmRIvoCAMd66pCN8W5hSZ4Hk4J
e9jLXfcAT4XQna+AZpeihM695WZK+q0cv5a96LlDc4LWEqYWVU8ijTrb5qsOfbUGsXb1Qt+Qyw8H
xT7hUm0lxMEV3ja6+jxXREQi+QPRukL1bCmp7pf/b1Zr5hJ0CmoMkyfi5h5zJSh2bVa+xLODBYNx
p1BUKtFlk/MEulJBO7ADeIRWfG0Gla9vQtnykhqE183TJF1ae1SzQot6wQro5/IBZhdggI//Lupg
/GFZfK7TlAk3iYL9V81bRKkBr9aSOVm/xk5qLH0UEdITxkr9fQ7D7J8mcOC1igOez8CdzMfj3sz3
W/bOkORp606zFpHqgW5qR2k7jdHGMAldq7hjebTsXXCP69j2TOMlhk9wfttJaOu/S/tlhXC7Kfy4
Y722wx6rkGzoG7Yhs8L798ltuALs1rjYMOWPYyte21IkmjSfHzsBcndhZ80ZAu/rKmm6VEidcEph
kn8UqjssW+2dQrlg/Nyz6HpifzvrxeOrwhSRCkES7IbmGYIvHn+7opPt72lvwdZETJDLN3NX8W8f
0BDuUOj37xUZZsiwuLlJaGo3jUQgtMdgfq1hdwxvatNYYdZ4ZkCPWREdDRsIZAipYqCfIVpOlISR
BQo7g+A34re3iXx4lREyRRccLNTlD91IwvcZZz7aZD85W8FOETFaIRdlXZaleicBAf/NsM2Yo4B3
EY321YpFk0nb+hAEen0pLmn75jmfpAW/5gSAs29dqQvLqeunJWyNgMuvQpGjWqQI0CgmAGLBYHo1
BqxTkRY8A+4YspQBoCbmuaIf7++dtsnBv9x5PUw0KF6zdszkgV0jMVeTdcdZ/i4abpVMUqTTLbsN
FOPdq3UgqJVtn1vlWc/HMBNsLXRgq60Ul/nf1az1SPT9yNvhLRhh4LUNX6YwvGLlbNxsBUPvGyQh
tK49ooVJ94ZUKq+/AmYiijF7TOhaZDmEX9ijP588WiAHs0LJVFpyCI5LQ6V4SgJS4LzWEQyOF3PH
dRuE2D2Xwc8uF7I+wxyWC/KFWekDvInKevLYmrvH62FT5IQmkc34tP99X1qoWSBtUobJf3kmEM2I
UFqP6aOuN3W/T5pO99HoOJnxqym3ydAE2jShb3T7wDmqF5H8Or0LJZVEDYWmMUDAiyN6CusizksM
TmTpzo5HaUC7PSa3acLVFgMR7Qek7CzZ7vkzNbeR9TOGoizWEES14T4vJPZHY0V1IcPWuBkZqxrx
5R06eMFwG6JWTuwUC/+l/spsY9lR/obOPqd/9E5Jr+pRm/t9RbZdTeE6S/SYxAcr1g+K3Ux98/fA
KWelV3XiN14/Ey2OO7lh8wLjh4ip1KujVa9oVn0V2S73wpaFBYUdyyS49oBwU6SMYmx+r8k6Bhe7
sA6zN0vpEl7l7WEa4OJrJnWq5JHtEKMZNorrKRZwgB0Bh0E4NC/ekmuZJVRrkCVIZhI6pLIr2vAP
ZnQH11r1yG430kzf3yb9gkSExiHUU5dqp/sZuf87z67j3c56MX16821MsLakKbGO1Lsb0DMH3ATR
dzO65AdqobeSDUfLVyAegCsVlxCpT4lcy1QZBc/a1flpRbd6p9sPoHg1lL07RTcXOPMmfED69cfD
vToqDp5vGitMLZGvrzDrWlm7AneUg/sNWpV15InTdlpj2jwm5iEdAvGibR6mbXU5cxR5lxwsuQTK
OhAcLoAwYxdT7YNzBWqQL6OlCID6iUjF1ntYKa8fJ39txZa1zT/IkDvUai6ysSgOfJNU3WvXsWE5
DE1xZSeKy0+dk2I+LPafmaMCl8o8HKLYTyehWipdzIYDFuGOdnEG4CpowtgQGKlpCXBc6QsHgu81
tguLMp7w8Qa0EMdRUO5R9pRlTEVnXMa5F31WMLm2wOUXrKpOTjCJbsR+4rgFD5SpRX8v82pqhNFo
GXiHKqC9cFX8+8RwlRFdpGUI6rFB9HeKp5xBfwFswDsDe5Vaa9byt+gBWviKkBgzF5fhDLMYeQ08
kHWjL/tuhdpfknPYehPP85IrxTs8y8+NPI8cNBTMCWxChl86t7RnTbzkT0hupsAXrogM5IZaNEf2
BUgwyKIstwuibXQL/E64YZ2U8RYTF9eZGGNTLyNrXmGLd9gfcBBzlCBJYbTX92EjEvFqvDYPd7i6
Ynla/B6EPLtath9gGRjesmHmOmPzgFTYXV33coOyZwGDVqJ/217amp2msfs3Ti8rhbA7IHk7md6j
PN0d2pQ/bUj953d8nleSE6VxxHIeXjEiAxJfckCMjqHYfLmFd0p5ho2AjnitnSqdKzVE1P9ojo6S
u508hiWyVHA2CP8jUJ1i66X8u3ci59Zg93KQ454g6HM4VkREuacjBgHRond1QaW/pBLd4u+fy86f
cD2/QQBvHLg/P0GeKMFYXwkhWUlDDkKjYTkbbehTUvIHCBETaa0XPL4MZqJ6JwFH+a8XcfeqpgX/
aM6Iek4fFQ3yW5RuTjRNWkFL//G1Ki8NsFsmekkqC/yrv87uaEPWbUQs6k5TXchAFsftex3fQ1mz
B7yO3eWjKAZFAjFpp8Zv+Y1qrAtpY7fJqMZDhLSzMM3lGthjDAaQys17eQF6yh2VzqYSeAgb0T9y
MPyPwoBM0T0aNhnH6y6n5367YmDZ/zO6ymnSCgbVgHFG4GVubEeDLj44N3uUzuDfI2WlOtwMNbJn
+CiosJ23Rx5Y44qmQIplkaveEvM87iZzvvvlP0Dqd9xo2yse7BQxP0Z1qb3Tc6t7hxERVUEbeqSi
5ju9PRXeSM0R2xH6msSfKQ2SPnILAwBxHH2iiWjk+vVFYYdlWcuXJackKbvJ+qgfs5rOo1BOcP2n
EVhpucVlzQkFg8u7GMNM1H/ftHIcqnvX40v9x+INAXfA1XfUwHByOvTDVNHjaN1DsjheXPSq8duc
N6hfHVMmghApxe0C1N5JpSzSwDqfWD9eVNuvrqo7ZbWMwza5FCExFRGBmirJnvWegLpVhe/TqaIh
wxv3SsvSs9YUf6+RjudYuJPTGgxqlocDhOXsZJz98PUGMZ1ITKInqgyb2OXv+jJNEpjJkzfetSOo
dcbw07tpq3/+HB+VPZgaHVNPAqF66kzlakO5M61TvWMMrHZ/TEUutt/qg90C2/7DoFmlilkTIFed
W5fsL8SRPebT3YdcsepQK626HvPL5zf8l17mRsn7JaYGfBFEA9Md3KIkIt6+YIEfF5Hq3NkzYlG/
7d29Ac0swFkShgBawqP52nRdMvXAPMVyPijOIa72q88DU7QSFLFBN5s21vGHMyJ+ZIrIed9Gx3Xd
uHrz0sHJ0NtLhzuba1HbD5zEo4V/SP5S9lHALiuPrqX6bfg7Ox8mDEQQFGB+Jbsaq1bIPUxpkhz+
3kcoJLvpcU9YPGaHDiOvBcVgMD/MiJsgu8Bnj6fFO9mq9W2T9gsCery5Ba4rgm2cRMTELg8Xnh4m
jaAVQJ0/e3SnWuvZfsyen2Xw4Q5ekXTvULoU8lfmu+olnsoiOsyESKcG0A5DTY6icbJZ0B66nrSC
dXZXm/p3Am/IzC2TiEQu3Fnr+uajYFv+9E6GyOS/QQK5Jp5AEtzkvTw6iwmM9ubS2wdmCNszNRMb
yQOosFTsrEN/5WFoEG99FHakhmkC99+gpTpkxlxOgfT/+9Lp3j0l+Fa0JSXNG1FFtoagkW9ylmwe
FOCjq2c3LKYpQlAtC+Utbzr1vPS4Zys5rdma82jX6xEh13NHG4yUesKu8DJWfmtcbcJN3D4JTSP+
azbpTKkqfXHmzg3w09CAp/vFpFR4evt9qOg/SOa8bRh/TmUI+lflz7qU0JXLotxHS+nk+lxD2xFH
tMc7g28YaQdNiYLpaN29ZmvS+pXY9pdKSZXw53tuZZzmaFhN8U5hKdd5ZRdROT450MaYatk87Ir3
xrnwglkzlB643luzWR0AhfwiiKbloXIzp0cRCv7Wy/L0U9WtUt0DGTrq/JnA6QA1OAwGEFVCRw4a
FaHR0sH0rjyZghYRiRcSaOGUZm2535FB483kHkrITaZfpiUhX4hnz4z22TtIGe9bcYTOHVAtkOaB
WKJlNroP4Gj2x6ggfR7jrKWBtiV0UTK9WNSY9XNmrgQ/+zdMjeH70cm4kY6ySHwMEQpCrq9DNcrx
wYe0iXt7p3Vijedf3N2mxfF1djNk17LcitfvSnOmdnFbdGivB4Xaz/Pyjuvr1q9xRb4lAedYsjpb
3geOGeYxr0pVVNQkTbIETfCGIkoerMnlyUB8NBNeIMdpKvolZOHJooy9HhWR77GRYZaWNrs5SbXv
Ixx3wjC3/APpevjiZD/5l5oy1b8X8Fng6DyueMJFvToTVM+4THoLJxZpGpReUrYX3oAtlbiXIBuq
o0BeigKnCtlmdzrq1OcXF3XfiuEw4Uv75Kxczi+B9G/X8mYdpQLb0kod14EtEGLQF6Gy0aRxUCmC
xlt18ZUfL+fYu5r5BQ7MH62rDl8NUHsJINHFP3OHDuOEPZGfK7JV8BhUySriDVXgJjAiuFiujkhl
q/sJNvyFUAWJbvro2YyODvViOvjrUM9BbFq0iKrjaHb3qIiwybGZq8A/YpRsHtouwL6ShTbtUnQO
4z9VjBbO/hlQQXSexswBmFzj1pZ0zJINUX7PHijPH4PqsYxqIuwltlwx4Vd1SbUyUxL3deV+WTJf
X7umHOK1LU7wUBQYKgYirOxkLM6DPuvEL1B0+4n1Kvu9sxcbBR2m1bR/XOO1La4ZejTNxgkRQ3gL
21i78peZViNdWVKwEpH07xbpVXkFn9EdScJwdPsustuSr8875zWcfRz+6neB1LiJdY4cZvGCeC45
mM2DCVmi3xjrlLCRBXXYDUHaGdCixGN6WEopwuDLhgtrJ5BJ7AFM2O1xlXz4EZmfFXD73PKWZYtz
aINR2sU/ZqPMqCyr3sldIg4c9LqAgS4Q88GreBe/+Y69rflnvNRCu/H6y2ytY93nzhUfMBmu6fcj
VdtX23FBQiWl/tfhyx8gAlQy3ZVgFY1k8l/fvWwJuluwKL80F/5OE7Przq/X/l7StwxsKqdcYVCp
xinVtrRLXxwiw+T9xy9h18Xr7QQnAeMeBh64eEs1qSwSEkqubyXQyu8UJtr7exQfHAZ+X8dHKGCK
NQwHZDKWFv0wao/HwITMaWeLs/mZKhfG0kXA9YMxYfxXdYa0ZnokAfUMpSyWWhbXuths+Wrddq+y
8oZBm+kzJKGhLDBtmnpHWzIJ+q77Iwm9dbI1Vqqaq6GKbPcqt3nzBMaP7XWnDiJ8+7J4mecCek9/
baBCIsIRIJ1S0qfYPTZlojuYkwvVVF72uv2JLbL/T7q1i37f07gTq9mF8lDrt1aRCxZWdcDHVBmQ
fnjX0MKOuESqoN1dftchN9552nhDGeeQoLmrqo9KaEFnKpRM0EV/yKGIZ2fruNYfqZgadsBoiI3C
aIugTejBiENoOlW5woJYoUw5RTpJ6C9ETgGmp0Nf+S1aU60pTF70voAEj+enTuzpIajKBfU9lfDs
MxHx7OOvSaxXWGHncdBK6ZNTUdxdoiCme5twJe3sEVe1jjH2BufHkg8CeX8sDBydYLhzF6+GMfLN
+V1TTLSiIS2noaYND+5QBlkKYCfz+CuSv5otAHfobTxp3Vy3clKOFt1aBDeuD7VPJKIrSnsu2WPV
cPBFhGFBQCqDTizVNvtkLmXbuzTbLQzL8a/t7A6oXqSv+fwN0AymFLsRLKjBCbFJojsdiJUFN28p
srH0xmior4FykFzRCTCTioryRdvyJOpZ957iwH0dwBZNo4SZnXThF1I9/nvG8A120N6RoIp/3Fdh
t2kIQQQoY9Bs41FKGpBrVl57cu+ZSCFdCjVwAfF6CMIuYAElkZRbJKiZ7HGzwL+4fG35a+F9oEQi
A/CKKUIA+JnFvaxcouvpN90Mddecr8gjdgdmMprhMPV+boWxCW3K3wdMEbWmddzWbZT+ZgQNUn54
8qzWu7kfq3DoQT9NuMNm/DEC07ti7l069+z70sEjh6VswvHeYvum/dmQcB1jbgUlNRbI8TELQUQO
hoCrscL0yp2vZIObTwV7AUPr88N7ecMB1SBZroA/4VF99fWOo9hyR/5wGPeH3KBMI8ovP+tuv2FC
zMIbOw4UsSm476d4FRiSRaFGDBXnnFs4msz6GrKLQbvTpehM1+DfFe3V9ufO26MurxzRgaOyDfie
90LeG5vVJWKuY+cojicBZy16e8kizd1b32ZxJUk94yPxz3qCMAtrMF2DpqEpUKvqPYCpiCWMKfD6
DhGnDseLwOk2SaAuHmCE70tr+EKHZCwex9iWFO0FZHIvU3b6C3Bz+RTVC3QbReT/MonAIXi3ZgRu
NOJlK8oyIwW0eBq64f84rgyLF//LA4im04VczNAd5/fU1x9oPBEE19yG8sB4kyaJ4zOX76QbcvL+
n0D7sJUcjMOnBkFYivF6Vk3K+UZ6MXoe8SzVKt5nXleFWMpXXh9r6WX8H/bJdnFt8Ch0yawWP5Mi
OlB+5/TqH/WEJN3u1ZW2ElJE7RwC3KGtsJ0Vfv83qFlRLbqoZUNvhLvWuE0U0m1lI2gvmKeze/SY
UQoN2MNz9zE3esEqTJUhAau9xQiweCnm0vf5WVh79HaRl7ecZK85DPeqQz0+j1vvnCQavKOmkMtA
5iQb69eMqWcrv6se3jahk1xBU1aIGjg0popq0XftqAW1AOF6WvXF1hnvdm+Q+eKUaEC6OBPYFzZ4
awuoLjGZmeVD0utrSAoqZb7Npfv0l3z8qWZj/PQJ/et42gv97J4BfumzGoExA95ftjd3+mvUJF8L
Z823svsxbaAAQh6nw8AN556UebIqgvhMIrBtiVM6zRSiZXoGpKI9tURVSptCWB86b2OYlrchCcZi
2slo+IuzIFkAecwT5ZMC2TCqpFQYq8CiNB7YnBjduLqSWjg9JLUqNmuVho+mrzTwLLpEXwSCrizY
Xflbl0KPyoBMLW0iu9cGB7V2ft0K/5Q/hIGhOLuKp+xf/KGZltkIPe0+Oe5ALsl2+X4gemlnk09z
Ez2gVcDfZirqJ4HnJJ0929FoqgGDvznTouEDmq36oOfRuhLmjHgCsWYGclntS/4WesJoxDK8p4rR
jEcpBT+pXj7zV/DWa0xPy1HUGra3+MuRK8JASZFwjcY1GfDWizUZCmvzubW04GpUqbw7kknCvD3Y
OqVmqO/s0YoNTCVDksqiff2uzkwK62Tq5kz/7PpIpCXd78f78aHoXXLl4sbf+PXdxeMNUDb44psb
KfFeJFY/0h8bZ0Mws+AYzgSRraH31XKBzzQMa7YenPTeN6hqL02VR2y8LznNBVixJJ9MhO5skbzI
F6jd18XusQeBPvS6PqoedanWS+IHmL0TJUYDyNOI1uvjexG++rC+3u7DxNPvF7fwC08AN+dOW0Vv
pCTCk3ekZpNM+iEAlfyCEzCA0tt6jzeLr9+I4cwlKD5XAFmJxdn4WESotFSSXqejuWmie7Dq4J5Y
mdzX1qxE6lhVycm0aa0xqWhXGeqJ1V8G/JJ/rwnTXa6z8oEJSGVLEsEK0dezz/ylYvJgy1TYsRzx
OGJapgBvErjvlgq7hdwZ3EDMpnwCUsxk/uFX/bdScmlHmac0MMxM5x0+WKoJnCWLCehfsDsMe7hb
ipQln86bVNotRLGsVB4zz0Pky+epaeMomp+TJF18QuiTMAhsf+1zy4lfVVr5pNdglH06W+rKO3/W
iF9cYOBzKC2UYJsLQqPM/UTX4+eKUX+n6umOpKhAAAcqrKDtYGjqz5EHr2PFujwWtB4G6vRF6wpk
Or8oFr0Uhpe7ZzSIszb+z3wCnheo9LGkiT+t99pOYTL0a3iPZXDShIzSolS16+arrOAqY+8KSS5l
wKOZUfg0I3ZQP1DwQXaWi7ZcNBw1te6rirzLhy6lqsLOH/iHcZa36Dnq+O3XJzLjXSiWb3Mt6oL9
+KxzJoo2YE23dXhkKqTidGlvxWeai/aeup6XPsglLLYvEIAeHI67p3Eu1hWxxijwBfvmslMVhFif
IMnQatew7xwmEEbEBVTvmE7bZOLPCJLW5BOXqI30aBThd9hstgX99rrWIczV7tDomxCdd2FOjZEf
RLas2/cz6e7lkBGIvn5iwyMsqgrwlzncyE5MJ5t6ubGS1x0GiGZEBxHviFHGYtqd/bVxPlJW5Sw4
zW9U/G+4tzCB9Wyu2b+qjO4wRsE/AGWzcTVnANZ7YOdZY0xB6uxflQ8EHKXWGYohGWeOSFBO8Gyv
ez3uGMEbSUqjG4W+ZcVDGtulw+Ot8EjnRWjN1rhPpm0hh6i4ho/arHUZCWGJ2DI1KTIDIHTDIew9
K5bZbYg8Jf9I/IJ7YX/8C8ZGkUjomQ6MIcir5lXcFsA254j0JNzM4feLoIokwlaCGDMnVIlKOS7z
/bLkNlbXc5w8SMetXX+3F0+haAilmWFluB2tIGJU1l/LlaOal3A0XiXfr031CMFhtTmWiESWUDO0
ADsUXPZ8RIvUS/x47J1OiP/zK7iJHPQkmtPkiOB07bqTcKHU72kvFa3JTLz1v0XC4x8UMppD/MnS
ggspAszopN6QByT9VBNyBATSwq84j6P+X3N4Pi/dJ/vQxNSVczlY7uTnfNVHvX9JcMKrYJFAuhGb
xeMvKFPmZfDj/iGm7rabLDDxbDTp9WekP7wWFGU1EJtiE3y+3SeBVJHGI+87dkBJWkAyJQoFgDpa
xV9W7WFk90IR0hL5j6lb5MJcRUZv6GboalsK8S3un20Hy1J2vKjqOE8I+usACndml5hhwFzDAjLF
3Ax55Yb3b3mCGZJRi3v0IeTpzO6ho3/DaPokuADv41NN8h2X2/1CQr+G2SIxVO0s03hOmcxtvh5O
BHYTDsd1oB1bVYjrZFNgYjP1LuAeAHDGQFa8WxUaJQFk5k4DPLs/wae07dnxz45uwGUDwwgV4CBC
sPAEapSyWatzpUyh3h/RNorkUESc1Fa8bxUyuf7NWdvXaT4PSlmC9BRFypWwIg762aOwRYT+xA6p
7vamvv9ycDiCHiwx/2fZN9bx8DRqezpkxkiTdTep9vSHmbJDXIooeFgTf3kYahcg+czLo5gqQENT
3WaQlDmNi3r5/1CBhvv0YEzhxpJX831jbgugmr/DF2I0lw/5Lw9FEaEArMpqbY5oGoctFgjNwtYD
Hzaf1+SOrO57mvZQ7dFvYM3tcApFfUQUnrlCx207w3qTjCJyuHKrnIeanqGJ2gZ2J1Dp3sstPpV7
kNTQuMzF0gHNGtKyQtBu2FMVWl0v3ZdibQjnx7b30n9PEWBgf1aaHHNYLUO94nNsxSfCypT7wTN2
gGYHxzPTXSX6bf3uzlB/UJCTccp5GFbhKyEzbQGxjsj0qzuOaTFwB/HckKcCZHR1BDqyeeLWM8b3
emTUdWRDktJEzdDoMuqwiPe7c5fw/W3rQt+Ks79AVVTiRRNVA4cv/krH91hi7naCDJ5vx0j7Fxij
F8hx20FP1IKFQUvGbXWJfrHZJ8Qu8F08KQjyFcyDlO8TIXOTK4IYpT/dIJk58WBoHoWzNgHOGuVu
qWdO14usAdLCZPQk/W/hyL2zvnHscHgjBMZPuQ0i2D+nFpqm+LQltzNOKZGKBsZ/sfnVQpJsjPTr
RTJLYnsluvA2MknqxcrNMULgrJG1iU69PjLfDExZkvcG331NFT85OGo4hFFD5iatPMA/hJ+lIiyu
3mj0HdGF/BFEEO41IX0wr2WSqfEBwwBjHiIGajeHI1XW6t6J7vQRPUyNEWWBy0TSq36wKQCwhV9F
3B1RGxIB3YuvZyWMvyVUH6BtrrZg7xdb+LwIUr/GvXkEuiOk64u8cVcxpNR6HETI6BcBttUYR1Wb
51vr4d+cShSjQ8qfmZdXkhlysOH+A5YVX0AbV4UhfRaei313gUblkyhwEOuWjsycX9PbIlhkCqUb
wkX8HARAi+Gpos13gfb44uluDkKGiOWYVTkhRiYNj4P7TcAUDZ5/+gHuRyIVD4vdiM5WCDWNpf4x
0bGqDms8YImcTNKf7rS+Jc/jdRcsWoKTGsdg/vxQ7ZhoBM73wuJooyECsFqfri7o6gGfw5bjTTD5
axf7goSTdEwiORg5RgS1UpH6qKqgScS6AVedgAcc8sHbLE4HC3l1YFcXOIsxGAB+Nqcxo2juwp0d
7Hu+s5yiv4Wm95ZWCP8QEECOiGotWNe4XWBaGZKUFDqDGo3MzZZ4/JBxL0C60ougRMOr4peqIVfx
+3AUF7ozdyrJ+VDL9FMsjiS4xVnYK2Ho8ZWtHwMr+Aa8FZsA7mc5odQk0hsDeuHPWfiJYc2ZmPSo
wIook18XKj7698dZmVhDTamw6k2UOAaCRCrnnyIdhLRF60fQAunFNy/B7wE5nXgUiLuONZ1KJWNl
qRAdHiwU2Iicym/e6azSHvZbib8X616StWysLmuQU1+DgH2tvk2TDKiIh5IrHrRLQHgPcQHqkQkv
xyqhb51Q22giGi1ULILyYJRWBrlrK/xrdju0PiKuPns/hf9ZiXlaaDlxo0byRqko1vhO4k3SYnSY
NES2UXRUtGsv9bisrRVMhs74WmwOBcYxbQtgwNqs1zy4DqE68I/IBLgNBYLHrs88lTww1+EGkDIL
VGUgckQbAL+qWFq1t2wU4FB5TD20Zf4eZMOwpT/8+IZW6+oTcCLnnm4PTfE5ic9unq8MhqpC6zCe
2CHCq0uM2RZbPxyfonzxJRtHzre//Cj7yIsNE4btKQQu62LF8k2yMcQdRrkMkSA75SWS+VHL1j4F
97lQpIWktc1nhrsC0JSHBO5xcLh8/BtshIWPAmTmqTyyJtR/z6lA5qPUTGuML1wWmIGJe4gt2Pi8
4wNqQHXflV5IZqmuEMz6pfTNZdzBZBa4/cFq5nJRj1sGMsiZC/bVhyeOpk+br9TJmHxh65kJZwSp
phLzzrym5iD2qAFNMR+B9HKXQJxVfs6GUFNdlga3eh6Av12lLuAxflJz6KUT6/gbAVydUZ3RCoNN
YewmlC9Bsi1H40F6XJbIknTJ6ze8EqGE0O99iLvoE1RWWrH7GLZIh0lzDjkQEvffv0Tkfd/dP3NW
E3bmvk6ywl/V+b9FQT70eqoQg4fAi96LIiKD7yHrj/MzkCjtBNypfciaId85TeG2bKj5shG+I++r
Zv1kFN86M67DTc2Ing8oj+5y9QH4LHEpgivl6GR0WyAWovMnnKOJutzZ/LqTzl9uI1+MRBvI8IMg
SyGrRHqFOWdiIV9BSN4Xq7RFhdO21z8FjDBzeC7+hTWFb1JuzbrePOF4YkqHWONNR8baSQ56eJoh
bc7d+IiPAU4BWCkKRw0gqXMvzerAgL6ZrdX+FaZbxylFufzVs+Yt1XxI0gwXkCVpF/7OQBYSZxZ7
oNrcRZIaev2NPLUgAmLKocI4BBTwPBYCvLJLbBvN+HVGl35DY8y5Mu6BVYP2VgvockCCariqBOUY
WHupid+uAeEUiBBD5XQjzQY09Ab65Zzrl4O7huMaYg7pQIbzvUmyF1nTBkYik6oDbf/HjtSluExL
KrN9vmAxAAudpnvLzI64CSwoKmW9F/lecL5S0rZEu/pdOm2lKGeRDHex0L0+/rp7SeXSiFTEfmbf
zMMqe8NEiSnCTtY0wjaxWW48nvcgEdFxlnTUuM7xsxxC2xKRwRveYHf8GENtBkw1jl85o5VotbNr
ilz5toX1fssQBKgQ8fINEdwlcMXV96j1FYdM1HM/az0tYn6dxg2hcomQSX8d5lmwUkfjmh4Rl63c
9Y2moC2gYpMP6hJLZQBGgLtLUgk9BQlGc9Lizpsk99suGEDLzaJ8jQro3zMdzCHMF/gfeSAdB5RV
Q6K+Usv1+CksB3204jC163ZRvo+jzlIlheMaO6eIRHk0X8g/ZM8IpECtUyZc1M3TzYoYJl6eIN0F
AZ5/5w16uPEpXICexByjN758mPd+UMrDEFsE8hP48iyZKANr5GN0bHnL09v1nQQWBHgsRFu5ld22
t8cuT7rCw5xcFd6iYOEN6DPfLxK1YWG8GgbrJUHRIgecyteg+fGVCCYT5bD71Xa+sycE+aWgv1UC
ohKaU4eeJ/kyjWGirXFkkIJMPcKdgM7w7/3CXyMbTUMF/68mxLH3MlghoeB63ohrfylke2Mxfg0x
uTW1h1kNdEvLgDZ2of7dnZSmU3oal/21qezIZQpDlTkFb5rDSx8FDY4X2qSz//w1EdNUshTcSw/5
XaPadqoVFKDGwltxu1yjYCgpwQBO68aMRze4hHAJI4e94Op2sytgpZtkPnDofqFGitXlx/FpmOkn
BZjbZ0bmN/TkYppWKo0ahxNtvGS5+kR1fjB3vugtDVuWrUOuSh5VgGKyyBRqPrmSGT2VkUR2nmiz
I1pBV8g9B+W+FhHuwfsj/3luMO1VzAbcrKbXYgl90qwn4t0uL4hEFgbnsDOSfHZBsFGFGFwj0qKa
fVr5jisoWGpnqHR6fe9dzdysTRPhbM3lauSpJTjpZiXcgGHaczdR2kLevxotm9HYzWWvEEcIYNRy
/xAabQqqxVukHUI3xKuA9UdlfA2dEplmulb3fWnzY0lMprgZ10hb5nudyJXbCDH3yyoVP9WE9LXM
a9+kIdImbvEE9dWbudluQIcKsNiThRmqISWjbOx9f7uo/0qlUoFPlLL9thqvrYwygCovvtpWKkBq
YOpNB6RU4L0HkYfEB4L89fgwM1SiZg78qOwXy+ZfrvoES/pZfVnIpP37LgVYrmmH8Ypn0meAFPOb
Ekz+ZVkJ/QVmsmPJgY5uKTaOUoxMkziRuSfG1K7XBKamvfBLwMQMwFMScw4sbFAoboR+rGyf9jgy
8GJW3I0MMT5D5WN5wiE5zynvQKp87h7fxVSjDl39TClTkpEu+z5ix/3GmmwlCejQWNomoskkOCBb
q4T8S3QoncyrlB05/EyewRrNqfQqeCGg5JVXSGKYb0siPrBADBmuSv5B1H45mOPJXWALZj4ahN+V
s/XBh+Hk2t0B0DEAprdlavfQ8IdRD2YDswIU4OBYHtKMYd3YYRefI3qhxNVWWFPwN63+oCc+XJD5
ko9+eQ/EE8R8n41LSUwsAvC3zRxAqs9CAeAxuu4h4rptcC5yj9XqxspxtjzDwcCw+J36sSmGoMU6
tldXaIwHUVPMHgyRyxj1/BxWrboiyTunKp+oulS5E9zSx/5NroKF+njBpLVEV9KxipBMyR/PJBwA
XpRMvpscgLEjYR59xTtpcRCnqlR+nO9RzHq09IYt/KTS/Ah+p5KYIktobe7a6mTdM8vxIfJuasjB
fokrZ/yih85b8qjYfpO7tlgj3RSRrDM655VDvOqyIGKje8e9yCtP+tYCt1dIG2Ipd+Cd6MqqqaLO
FuAQQq3A3fm2wsv/xkb/JXso3c3zXNfJgX4oAWHLIhgvw3Xm9qEOXCiJ4Ot1+bh1/MnwDEZhVldQ
PF3e7Z5GPIsqkGEckFiiCE6yf6HTcYhpSIeLUnnKYZgnyhm/9tucnnYUc05EvIg1prY5gVMGoro0
H1iMmj9mjFkmBxRuV7nO4049yGYa07r6atnY0xKdBemrHJywpOfUhuqeZ/+nhaerfBV3TA0FSTYq
/BmjBV8Ny4+4tKUbVOg1r1e8+NYCAdSEZfSjNfm4eqREL3Hk+rrG48felMLYMK0x6PCbQnvur9h4
0l1uR9NhkwNsxg5yer8j/D8ZHhQqJoWwLUF/O1o+IdHs2NHiIiV86LtO0JiV9beEO/nzvEe4HGTd
8GZYkoW+xdeqgjkumgPuityxgKipxrrUgRz73zl0s5SAWL/i9zedoYTSwgX2n8Ypifq1G7zhId7F
kwi1LKAjjqW+Ul2fnLX6K62wiLNu2w7t0Itdjh29/hKYrHLTlketHRWgDcGttPc9NoH32azXKGr7
Bl9na9J12U3HOR/GFznDVDCXwCb4kJSI6PL5LKm/qvHebGud2lsjDy6UAMaQ7fJOZEowfNvGEHgy
SpZSPeYUw1UJRx9Cei6gX1CjHIH3eq10GM/8hjPyO31oK9Vz3MZgZotyF4O4u8QFdYiO3Z+vEtn8
gwvZERJ0FUFpmcTrtqq8IvfXMhu0oeKxMhLvnClPTkGYiejeVciyz3mGGj8X5d0Rg3j54k1mbKjF
WQVES4S4H9rHqYY+bnCCK/GPIguF4BJj9/x/vmQV6fdRd8/Zb/omMysj8lf/3Kk2epm+GvExyQUM
w9MvaFOY/DPfhHUKpsLGMDl3gicqS4nLyjhPbLsEVIEzSfNVjB6hvdRmf4PvnQm7Y+w05h5hgtET
YbiyqjuVKOEDg1fCvnTC/tDOLcuDPQovkjsKEtyxYt5LyTO2qMKJ8CiWyFrThj18LeOse21UE2Yx
UxDU2qyPTdcE7u9JXHzMMBtoZWSJKlv/yi33lka5H6aAYJIw8Og/qcuUx44YW+TP1cqknEO4nUj1
uNmNjEQIsOw5Qi+ILXn94guU8dNOt3Aw4wJFk9kbXvPrFdZXX7FEoCzKnFOybPubyhMWu0wra6pz
EGfL1ELflXYSDavLmQ4jE3RPmCW0z2hAdr2pbYuAxQqLAasR/C6N88tIBAI537s/Us/hZMrUhPiu
VY7UJv2mPhGEHNH96GWgva9KTEYQJzKrqH1nEqN0RcnlBw8Y04bCVzfKKrRIIvlMer0YJqKKdE/A
WecFJTDZi4GIhzeftQ4OSEsfj0wvI0vQRjijmIj0bX983k8073TtXSYDmMIt4JTOR0dOGkWAbPaM
YFC2XTRM6dWMyjixRRZqP7wGNxOfLY6LVADsGzwNmatD+HR0R7rPF7RF58lTbEEY4u/CDyqt0S3l
0IojNLDo0/6zTKsQe6UivbQQymDqo5n2gkIk6/8v0osXIPc/ysEfxzjBDJZXAVIJU7oNLmit0uJl
xii9kbmdqClTGeiUM1fTsLaNpa21oMgA8XMQP96XFpEAMm87elNyVxG3LMPPUdrt+yjuTvFRFSo2
RUupQNEgTtv4u/30vt8xS1Yi+F/Q9xH/P2kWpCZj1Z+vAj+A7Wk0WLzBmA5uUjYSnGHUcb5OzwuE
k9hcL+hRqmohwqrFg5G9Gk21JmTdEUVnGRiLJIyqetgnYhPq+bMBEzA8zkpEZaZYgsAeuWPwgA9c
Pg9DmMaOBEElvfCzLxp9DMHmlWo5Q6CMBDpEbcEESVkmPm9lfF5v+byUMjlOi6qX31058OGfb2IT
H5qQ4Dk85WzvboF3XpT6T2LsZ8/B1UG78jUXy43ED4dPXz8j12YoJOIC3LiCGxTOnKNQbBVxzoGP
U/dAWhW5OM2xXdzry5IoK4566a6uFKk+LsIFpqKLnKh9s8I/URDOBaYLpovoRBndS1C6V/3hpprp
US1B4xW5Yln7UAug41MCH/Gx9bixEd2ji83FfoOaGlB0VGDPRmLV7YsHBdmAaO+Ayy+hbhvkF+/5
jwFK/kTC5Jt2W1I0T8Cxh0Cn4tYF/BPLx/q0BxbNEoiBkpGAsMgS/b0GH9whCaBthvJLtv3mT9/i
wtpQId1Tn6bbrn6otWldORURbpDaxaUb/v70ZIhav23CsJ7bKf/pf04si8IXGYBuUwJWdOpJ1urK
l1SLMBqIuv0l6QmR2HHNsyQvQXItDRSAXOnsKGLcB4BBrdM8IyubJZVhC5cBEjBzi7g73pkXZCQf
Vri0XZ6nCZOms4PaIpSKtdzUBhJxRiFlzyYznqPECer1rOScd/pDsh62Ote+0kvgt32+87K4W6Ga
sGZkSIkYIqeskWppT0qVAyuV/98tE0f+9PyVQCa4iGEW34c5wkPrgc9uTGgWCTfLQApPZQPFumxP
qWj1+UeD6f0iKVec439yuw/3BrbGXx73ZU8o1UK2FZABP53lYfyEgCn47FZR24SqsSY7b2uhZrtb
YnVE1dFEsqPo39WzBZ5H4WrtkrDLjMRH2skhxP5RkIMuVS3Qdq9qYqdNT8hUvY9yUyJI/GAxI83X
7T8veg0HVlJTQFIW19MWBljlw4Nt4+qzObvqmaOLa1LsST5AZnj9sDlutNVn2z3OeUq5GZNF0uWt
8q+ITj8WPcmqWcNx0NFvzsKrhH1kv0Yt99QEUwCM3Pt+AhwWvGXZ5L6Xc/zThnoR/Z0c7gr7uF47
uyWeNjA+jr7UnT1PJxrx6yX/Q9UodBDd//EbGoPvEEkXW8yCzC7yYeSraEqH6fT3czMeuLIy/V9P
iACHOAAHReg31uSVWT5mNjnvINXvQtVotoQ7SamXN9qopKqR1RYqbXqKrdobxnG3ZKx9JhFhdHyw
9qr6Gc1zZ0/gOMf6uql/8g3icpVEo+9gBCyDPX7W7oS3AL9HmcpUX88FbSoQiRTc0E/EdEmzWZO6
Fl0Rtfp8j3N933OkPvtCX/khDjznDICDeoH8RNhYoShvvFjzgVDHHvr6bSusYIgMVi/W8Sl6QiXd
a4qyKAXxR481p10gK+6KhO/pm2LLJcDFciT7g2WVFph3l7dH9IRElwWM6TTFguAGm8Qo8ed6n5RZ
+9Rk9miu8vbV+8BXFCGGa0/zdXYybEtInRocT9EjsxgGV76gYBZ2TbRbAJpJXWY/9UYqZJuzbBXB
4CLEzu1vwLA2mySgNx1N9/9+j5DTK0kto2cEEXSdPYZQ+DoWzidQe4JqgBEeM8idufed1VVa++SJ
Shy4Qepu5oYry+vGKL3rGdoKqTGX1DGKQoZvymNp/EtaV+ibyQ2Satas2RPLtLO7pibhf0xzDaAB
tYJaz04OOaLkGo5CHdvr34PXnNBUrCm1d8U8KPL3jO0UO+1SkVhE2HBf89f+/5NErTw8DeCzqmt7
/NY3cxsd/f+hTUwH97BTZobvpx3fV78ZM7OEH3EO7+UQ8vxXdSpZmObqmrSmK3swYFFhdqdiOphL
RUL2cCP7itEl6qlzLH4OBD+oDI9H6iJiYFDYcDcWYCmKCUaYXAvV95v0UMXb4daT/wo9IgmmhlKP
ftJyPVmF7TT44ejFtxqDyEfKcAD1RHvbn3NasgWFekmm/ASzwEe1ltZ3Y8ldNtXhg14s7mA2JJWG
tNM/f9JuqMt0tsoBmcQPKo+YA+rmWlK7GSgffVeS3jMAIq4Yxg2TIry2EDZ7sO+S8i6hp3tR1RTo
rDzaFKsy1lBrNuarQIQyoHkMWiZV+yKe6XGHChY8DOh24zBXHpCWPcxmi7bwGqFaULz37kZm4iHi
pFv27XjjqixA/Xa/azx7BlDFPpoVlFwnJxxHzGPqKsukL1+uDYybzkLEhz/baGDl4iY2BCh+qXe9
2jIJtAwx4LlL5Q89AFyiMTKwoirg+Psa+08l4TNp90yeVrn+tg/Np1kVVQ88V05Ekw3nDHBy/+XT
r6rb+gjQYvq3IatWg02rmlHkO3BExE2k/Xs3XFZ4AiLqrfqv7s80NDjt4FZ3BGZUFRV/lV1bOJem
r0082Q1ZCHIeU5ChctjLnn/SnuJss1YHJ0E98BPq6h//dFeHF1ZcN3jZYSMXYSSe+wJ++TMuj8u/
KqUcchCLHrVMADQvmWy0GBX/CCVCGZR3tXrQ7QpDAJCChWo1XX42wwZmLBz4dh+T0Sv1LqqJoHLH
v9b8kom7Rfg/7+LHd8GHr71SUEb7RcBEN6Shpa9j8udaD4d8TSBHGSt1NWT/0VcO1+7/7MRwYS1M
iXR3RXjNrCOlhlMZqnkpv7dTEjvXg2ZqnbNueXf39KRWoN8kiU9GjEy0/X1HKrP3YGvx4J4tL1fP
Eh8Re6Ozlo1RL23f0sZ+7xRVDNgwQFxOQCW0PTdW5S3NRdHXdlpDVZd187uT3vM8fKcdlyLbCEgX
s47VaaLB8Bk8Kn/iNS8TF5PvmkvWPVujY53ECCYXXM9ZkdmQzm+EC/Es6C11A7Qcm7+etTEHcXOQ
bzquR5BdF/BcEsDH/Tc3jeSiH8GTlULpyun08sTw24Qq705/G1y2F1jl5iHP+p3rvThiZ4hZsciP
2RZnzG7iwXLLmtdIefc3WK2CCNUHVeLsD3Md0240VsUMEVsKPwH34+3Di/JaCEdP8DZa5ZTmzpkZ
m9sQ26YHZJb/g+tLzDVq2urvm/y2s3KOGvfhm109YXuHvGuZ4jj2TJojplLYLf6ZDUvw+GbSLc4K
2OtD8tYX5D5Nwhox8P4ozdzhuKMZy+AS1nu8HNRjpDJNMtzmncHvo6l8P7RAd7rQyIllqfCb2G2+
u/O7GZzYX57/PT1CeoQCpUhN0PObVLw9DjMljcDzbgn4auB8unaogd8nwPPYv3TKo93lAyN85cAC
H/kfJA33Pq1BbJxBHrUM7epskK/xU0RA8E4O9YaBkdS2pgNcASZtQUtM0MUToxxmcbVa+inFlFIc
MlwKMm/nJUBXt4i7FM8uDO2A4qZfl/ZuuROUyQ+qJnX9FEJ79A33syw6sIo+eJBs8T2mc8BAN/5T
UPuylJQUfpbf5SA5509W9K73EpnoHxq3Vpv9DCknMzRoP54Ss1qslSGuyVgWTcXvaVS7Erd9ECtk
nnPGNgqeSUx430+v+FAw5Q94MSksXJ7owTRf/bMNOyfRY+9DdZ2Fxk4+2iV4y/tF/+SpqphvMMNC
PvuQDZq4E0wzzc8NFhFB+sO1jHh5k17yBIvQZDXUk6g/m5MnFFQc1OT9CVycIMWi/JhGVaAgh/Bf
Ug+N5SN2YImYk580m0TyLwUaUXhSu28Gv0HJdGUHLklDhvDOXxx/QCOvBciPrT4FdPhGVI51FLGa
b+7Rb9T/vtHwtYRoFrM2SCNjdpF3WSwq6nw66JHNUMMPzzvEw5U7sQdeYS6Lyf31ITGCAM8o63b7
Ixb5NZS3VthmzgF1P9VhOu3OdzBPydGG1VFxF2A1oqEAfLjzwPbMMigXYTW3cPdhO67NWvo0o8kL
W9kWPPvQ4L54vFa4+cgxH0eOGwTIusqkGBFJEwAeqW8q7i4VKj3acSvQLPZzl92/pxPa12duccDe
BjwvlAv844JaH5YSPWm1iUsVwUCp1e2k3/DcszcGCAFSJvE+hmOTUm2tgPuW9iCR8rg50IhpVcgm
8/DiJkvFJ2zcKW+bDMrq5gihy8c6RSR4svDOEQFWfnhIz3WoUR9sxbGiumbkdmOGxQn3ClM89NTN
LBT00q2ba+arIR7ODlAgqXCGWwSwFU4D2pm/EH5adWhrluVIIyCJr0FA52jYaudvIajvMkB0JKpg
wlhVz2kWKw6aHzW6B9Yq/IsJ6/nnhEFZyTd/C1384AQCoDKVuDRkDAN9IBxX7XV1PhwhRaxgF+PD
yPvId66wz03qGi9BYhEkkAdxMOZrq7t0aa6dcxVW10P7rOd6TOz2KBm7CC5NUBXo3Xn1clXEtANN
2+9EKBPHrhiFrq/7JHs4Z/sjl047WyKW0dg6L9XbnIUsu9Y+jJtdFpm6AdgDwk2CS1xOv2oquUsd
lrrSycFhQmMCSedgmBDCmbnwEiVEcQ310nRjkEGF8AciOe4n5QLzynjKFd41PifWJ0vcculy7RVZ
L0W+Nzx0DiiUzbQnOGRoiZmiHLG+Fj0x5oQFVJI3UK/pJ7NWX9NjoApNQFv0E8hyPefGazEyL8GF
5+dfRxF9VWiOHizVSBF6frT7SqJE91tzV/sgaBVDWD3wEHmbKPt6Hip6UrTpuXZPAnXCyVVOlmiD
9h0X/cSIy4LNOnWVZbCQnjQgAfwx4NGKDmeKKtefW0ztQpmx4kF0YfKN9IwCxWqdPxZBy+/DOPAj
qcO5QcQvI3jecgHJ0U7vrj4NT52DcXUn8X1C8nqeINJM0sV0fP7mWhKhK1u3CB/tq+5NInDJ8x4P
DFmne86ZC+SGFW3pRy+WRxLOOGbgztrbVYaP+9eeF+JjlsiZpyte/m2IuWTvM1ZLwcpXXXti4+U2
b58VRyhUQL9sAD+8DNb6QeB0siaQu4Su41LuNEtMqa8z+vTNiAvjYH75WPJS9P4kUrLA+L0ufO2R
a5cp1Mq06yCWFlsaR6MFik323gLnPs4uo5KO5WJ5VRtbZd5bviOeo8TqOmQrf1jplPWtOOztUu1o
VNVLFf4xydsCwbyUH1gL8SSMmcUxqFuIIXbeaDyOHMcepKfKFduVA1samJw+kmxxLfZ+aXg22IQU
EsBaLEZTBxZ7k4R0amvifPOwTeN2sxcHtv4kXDUWi0ds26fZLVdDAD50wSZ6hzCPJfdvibpxyMY7
/jqeWWNUiJYQJXoNs1RdgAVdpzq1Qbov0MMuP1IAbMmQJdWHRSBTtMRliw5+IIVI8Qar32bBJril
oTeYfqY6DUnadse9j5ZH51neynCPg3Msdcm6+hbrQnZoloQLo7Rt+DbSNoaoLkDYwIhsuVb4zk/M
3j/gYRnab7j1gtftuQRMhDMkq0TlgZ17yrXW6FSgBc9JmoQKTrAW6i1Z6fkxV74RM4uEuzlSOTVr
4TfJN65fKzHxrQ77oiCbfR3fJvRY0EipjOJkieFo84tld+sdpnIPX1SiG6Bc/8NJnQ5VYYGZXH+C
lH/HE6c2cXbYyQldr/MyERPKd1Lq8hepLmbCfyOTaHo2xKEx5ilr/XnQ1s2ipVNTS8wwz34fU2N6
zw0cDHCiwcCLSq7ssIFEZVfRTL7Mr3/RjyRWAoeiNikgE/SUQdUouiZNDyyPlgB3ZSSb8VvdKlio
I8hHi1DOEOj/SEli3jt90+2xm+ivlZev4Ju22+kx7m5cBBxxKd+uFgE3dS/Qq8XZ/yq4GzjmLIPr
zc5mOxfz0JbVPLrcwbw7XCV8MdyWa4NRgTkfl6Sx0B+taRe1HeELT5bPw7q12M9sjYSgrDMvN+fm
x3v8EZYiKeDpPcRRXAlBL1Y8TDjucx4k1q7PMR42aunsEkbbZ7loDoDHYJUSlJOmWelxhqDfWBFb
LzXSV7jjrCtpv7n8+M1WKsmad0ECtXls8QcTPwb3+kR7irpDQXDrhySYyWtp5BUUG1wVgz3r8xTD
P2YsGM+l8OngxbGgnRU/tKiV6p1F0k7nsJLBdzUW4EyEeQPbD253O9mQR7fgnbUJsAWV48q0fjA1
Z/Hz+yYag3va7CN2l1NuaTmRTNF+KQRSxiN2XNV5IGx1nfLOS5/sGBpNM6IXlpFwqnBhVnGbeQJY
lmr1GedFbGqDsNXzkRYRbZJLomyM0JvdTo/DNlgHnMn+R3P/t8C58cf1H9Uwb3XkDVpZGPuqwqSi
ZWBOr7pPbIqulsdH8GJZ49i6qBHNJPJqjfaCFHW/ZFqsuEtn2Cyx9Be708TZs+P7hVVUxYluAP7G
yUbJdY+ZpUlC4eOfE6spi4O788T4P7R2qflaMrWLIqtNc7ego0Oq168tv2fWOHe11BcD66St5l+v
HaH5/8smhmuxlOWbhC/WiIpuXiKvKzxeMOs1GW0W8Iz9t37ZW9zGPFha1JZxVukr+I9PER3dbLVr
DcK9CKLwWGo32mOtThZzm25NQDPeqhlrXCA+lezWxAUCXwdi5/Vd27Gcu4WzrkzQVHgmYPv451vu
A4UzdhQEigfvym9kYZLVyELEBPVFWhfJrNYgFlmFlYLoKbP+MveHOu/yoUh2c7J0fOK9AqtiZg7G
8avYzgNIXYBtL6cz55cQ30NT8rb7SbImwv0lcKLko1PrbK7mm81wYt3acsYk1TLdJAslLeMDmXK1
30n8dqpMKIMjfMUNmPWnTusGHbPnYXJgVoFZO7cupWJxk+ao9mv8SEsye74GKheWrOde4EW4Qezg
yWCsppbRaUV2WlVSgr2gQJs9RjTVavJOGu27o2hquOgHnanHbBHUq3tDx8y+Ofwc+sw1eC6jr/9u
VrqlkGI+SgzA9cgcrkvvg+ecZWD7hCaIu8DvcmmyrNY/L0paJmHZNMBbDM2SNpqS/yOByRu1n81s
T6SN9I8ZIY39h8G0WJhobRJtPPxzsWvHBZqDjR1ul34LsnC9VvfcY4fI5gWC3YXEgm7kyBx1tvYk
tgxKvYySH5GUKr+qQ9aEya4gbRzJOK5e1Ez/5Ojwm54WyhZkbAqI5DSMeOyD+bzKIwVjASiiuOHK
+KckfPGcOSaXNPDKJeYV4baX2024+CvryhBwNSKe3czseOVu7TvFs+gzUIdv1wEgM2Rs2mzhwwls
N3p9VNiGLpvDNYZ4MNIO7W3CNTGowHjKSc+5Afl1Wsv+9wCo+nRJ2i8z+/iuTSBTwLy7DT79YqSw
zq6M4YoGVtDr+29xX5HNTE7C2ynLmjuVnw2vC+A+LZ9nUDJ33XFpFZ+RaNb3HS2aZAbA+rlteUx+
45YoazictjpJJK5jOuy8t5F/gZ3flT8F8W8U8ITQv1Ezw3AtgTBqMXWtfdmJf8c4bfoI89UPw5+D
HlpZ3eY5UAK/YF+LoB9B5Sm7XF28Jbb70REzYCUBLkSEHkR9Oqt/FkR6HMcWoWQ8Iaa06CnXYLD4
qiVLZKkyajhouOF7o85X1j6dG+7iWXEzJnYF0G8Hx7sQ5QsNcuVTmTBf7TFgf6Y2jr1jTSaijS+p
F+fDg2Hmyir5a+kU4M1BaBj3oy8j2y8IkVXxw+W2yX9SFClOJAwFnijieezLgmuv0j1RRbmqCGzK
M1DyWaKXz+Pzn66V5FjNrXLQtM50RSILJS/riXEoMtTzNa+4FspdG6GY4anPfVU+xRPN/Fh0Pat5
9/9jCLw1mEpSCIdkPu0BZEs5dQkhrQINbF4QXrKW1WdtkgJAiC4vTRlq0FxzI2YOEfYd5Y1Uz54u
/3QvpUhLQAqxaiyivfPR/2E492tFT+8pzWhGL/RIarzw6cCxuxZzQNVNOo2kyahU1ixAvi9Orp33
VFhSxIjK1IR9PWHoJ0vXa9FpkIATo1EZ3VWflqWBr9Xi9ogI0LGhzeNxi43eN8uQs/JXlf/MvtOK
5AxoQmL+afauuHyonf3p/XseMN/1/I6Z7U3kxkVBjGTGee21O01ACQXZ83SEejPT66FzPcDXOFHK
6UHltJmoJF+48XTy6sk7fYR5KPc4myygHr5sjNkyZFrW5xzxjFz6N46CeF4mr6CRciDYzIOZ//8z
8NzBnEYvgHWzOsSzM5XHD11TAdD/ZEQBU8+y4nquTjX8juraK/aqsqicKN1IpOZ2oV/RQ9t9uoaz
UOFq9acftYGRHvrxrUjiXOcadeYFyloGFJ/1yX1RWL3gIYcpVJVRtQtpk2WDzxeEstCn3+RNwp9j
R9T8m3B/2Azb3M+DigXjJtGGFXMTglp/X5nMdfZgpfsYa6QGohLeOPbWOXMnFBcDQDA/fxqpUx2m
DZOuUMXM81xs2gFUhd4WV7eoeLRbdc5/L0ZTXq5z0fZGiNPsgIwDwDLh4bwVnGvKzBL/2UBlDQh1
5Zh84YffXsoj2IRUT0LuHhzXUVecdMMf7ETeYAhSnMIEV38SroBjnObp/bLW4uLxUtZnkeg7FLnD
O6yTnbIVezm9Mn9bwaVTNWO0UE95Qol6yBI6Ma4273qRK82FgxN0P5J4ZfANQKqduwU4/++0FR0l
m008Yh64o7zOa77SKivkRYhV10hzww8KyXESj+ir6xr1kXhWAR7oGRfqyfSivDALUutoQyIwadGe
Xh+P+/sXfFTUnyFcMuUJdPeVjDCV6mXDivX/kAPGfDfzcZGVbqeXvVBy9RQRPWxKDwCRP3PoKm9L
4V5DFCwlT33bJY52care9NSHPZxl4cZZcMT37JviXRZU0LvW3oBXSDSb4OHU8zJzChygFqqlR4OX
iOYb3/aaz+Mpr+rUvPU8ZhlkYdig7+JUIbhKBCHCyqeF1GDYNGi10M+b7koRaeMONjx9FH+3f+lR
KKL/50+bxIofml42VE29WTL4UNrtazO1svqU76uidLtfT03GqIWGZ2sA7fRgQLogLQNdjytj53/a
3QfSwkoq47lxGtZW/oQ2fY9BHr8ELVmEJY6kyn7la/RxoWiNDBR8KyMurrs/jZ2Tj5glSZDZfdvs
gQ3H4OWsoZbh8sEZ+lTzDxDhstEiprMedMtygzIpns2EG3kDdgPqXrGoQJQeOWpO+rNnx0PA2rVv
cYHEQXjym3au9B5pZ0X+SkJaRsmdamZTKP9FzVWRxRT0Bf8wlKp2qTKwb+pqoCy+Kpy+RewnKijG
OdXoqqqfA2K7laPXBMnpW6IhijL4gapLlxBKJnRVa0yImuRp1J1UWYrQ3hNJhNCr1TEARxlfeOBf
CYk+1iqSkzp8irOmBTFR+HPRJstANmbsw0X9RmLsGotClGFVYjzC7MxrJkJYme//lhaD8VqmtlbD
intoaAb8WNEQ14ZmhHI3n8l832Hm3gRfVCTbGVgtmzA/7BUwpxVcuz2N/vW3W15uMvPwjTP+ZI8U
GJqqADU6s+JCUlU1FWPFjm/uAYwyopR0Q1Lzhi7pEg8UEfPKKnOqq7Gat5FUCdUV2Ba1IgDcMEJ5
xCCaSCZqpUk877uetbt5shOyh3zZcmIjmcraSkFSdwVVZqVz5NA0yRrYG/NenTXH7TZJ0ARCqxqT
04yAHGRMlBcB7eFSc0qXn/6M4TWjCFjt1WcIzSefeN79FBP+xwqytEyQAMslCfc8hQNIbI9fXqg9
TuEEq9zcpOwFPe+O04DXYwwJa05apfBVsfQjOKgT+lz62HNkhDt4inQGaApucDbfsJm4OW0NzhFz
Sns7p8Yt5YHRVM8axw4AMwXR6hcEwm8G8yqtTh15/h6XrfMbwWQifXW5MzuRbsgdyKGZfTWPwoKm
jD7qfDrVuz4a7V9PyZTtJroBpZeGrMj2Y2C1VcugSTbJSpr7fkIK/yVtoJVzTqNTvDb4Bj2H6CJp
d72GGh3dg8hA5FFUfPWj8RG2Oi7EDVvzW5CqMugT27mAvoeQ1phxEPYT6THI2eoR8liTS70ejs+/
J+RShZ5S9qdpQy8s3myLu+5cKnbnAlHe+Vlm539ZIAKnwa8+N7HfDOHxa8AIZNhaHhFP5YQiDG+Q
WNJcfG9z/iWpfy8KRQiRPPexepQOY17oslnOS4ko7hq7Q0dhpYfYBnmg+6edlRaoj7ELTbSM869k
KLF9JCQ+D8CmKe/iCox9dtvejOFz7WqWmGongfX66Mh62yzk7K1YnNu+LbmDrlLCKZMo9Avnyum9
89ZLjh503uXwcoq7sE+giAMW1pOEaaO1mZodawvUBfiniylYNOHa77sqvAcMu2AGC7QITkTz63cB
eaRURfqQVVz9HO/+ONE3MULRiq3UaZD5Dqg5RQP4PEfliBksKVRT43KwycXMzpLKLv3IviGP55jT
V8Wl9gG/5nFYXPiWK9tfnbQR5fwO/zEyjpqcRfxHQ15T9kFhE6rHWI2zA1hzdmJgv+xqSmri5gGt
Ttn0BKxxVWg6dxMZsi5drMLyiEBhsJzV5Qg6mj3P/B+dyLIP515ltD9icspGZBOjMZD1m5g+jyKX
tCaaHqGcfGHcX+HYXdYlimsvtE9dgL4wyhvKCDQhr5ln62OZ1fMzIZGxacMs5fH50YxOzqzwIuE/
IyHe2gEc2ICDbvB4bwh7yW2cWySs69PAndmMQcjMYuhrMbPfHPcSXv5bnrUpOKLqCepowAv47xJz
pI//Soz1qj5IRaZ3fxdgrm3W3EmKaUx1WPQZ/cUl5BxsK44vqN+NeZArfFDPul3UbtO7kNcxBR8f
gJ3Z7pHETVrdEhFvpbVNnHLfkip/L6UV0NvY7bDSNS+fFeThHmV/4JMW56zosr4gZhn+5hBYcziM
cI/VP2/Pmw5NCa+Wcxym2JHgUGvD1PZ0QFFntvEm0XN+xd5E4J52YP8+ZQIRa9H6dK+Ojv7UbUMG
PmhUrVQAezAHzJyQ7GHNsFCOmoygTSXjUnvOfyuhvsnHCPMiGN/FR4mLAbU6EMPDEjd74IVhSO/Y
dP/h/Qw8GOIWQy4z5LcDK4hlvEkzQBj6RFkqIRl88WHGCBqyWEbumT1KbYmBVuoyE5jygaUPTUmZ
6mmkRvtzRG2KyCKS9t1c3PLhKnLVcgkw8qaOIbFk7Nx2Ab0ana0YJnj+TqHg7ucB1yOnnj0yvsGn
hJoxbp2hN6TKnh+0b64JhFYdLybppnWgxHyge6tICHn28KS2AiH+/jZIcL4WPwrjSLmDLBbn8BTz
nvF++vjoZfTHvyrUxHDQ9s9dX+zHb9urklb31OLRGYvRCDoIMLlfuF1p/7lToNwCGNgvdMKayQ8F
Sj+uaTnYtv34V93swpBaU0XjLtys+y8ySx3dQGwUPCcHKqSdRGtMHHLTLvDVuStd5Qu7KoEfgNLq
sfcogQ+8uuzXNs9ZrWq3TIdpd+e4V69Te87z2W7gCAzGAXvwEGI4iL1WWmE3PlR7p1QCe/nG6l7R
HPYqNNK0ERDfQDgRER1M6cyw1WG78YpfTgtGQRZe4oVDGoo9i0giFQrs9GzE6mr71sfdxZji4oCV
UQZYoQSr811VXE827g63fh+lc4TDT6+fPStat22iJ4iTf3vS46Fu0iDB+1BIBx5QPLNyTafcDr5v
CgTv77huM4DEF/O6JSohwBSqPyVDj5GRRv0arUAiWoBsUY4CmgoHYOZlq0rgGC3O6y4Olh+bUs1w
z5Pcm3yD2aOSwVErLbG4mfOSe7RXgTs9mlhSK9z3r6OwoLKg4Hu3uLNsSBnCqQQyuolNHn+KQz4w
hVnDjJeCLVDnX86VfgjfUFI6hffbJiDltkSz01O/UiZyTEc5kLdqdqg33wrJTYCz5JsJ0qFSRGDC
DenDOTsk9ubviKJTT+jw3aZq13zsjTq3yAPIbUvH3c/ly7LlNQ+xxW+3tOc5u7KPWO0J50zcS49w
Np0DzcR0NY5g0lv7NETthR27dh1VCu9cHpVPeMqBOWwYYxd8W4F9PpqZz2nw11sWtZR/m5iTy1N+
ZF6uIqf3pQ1Ca5FnKAmrrsRotinVi/HllRPkEjbTkCMUvv1frGDpqWUiuQ6S52f6BWNwF+IXN1If
fYRtt5iZYaXc0GLtvY74Jq5rZYy4Gdb3VxRtzcgN/s27MoyEjLOW1BxKJvKxNnzsTsFjfCe2CAlR
5LvPAtYQ8GIZmJnBRzX+QAlBjrWn5nB6IFQU/M4t8d7/UEQooPJ/qvlTZiPAyck5ogDA6wEhadZV
+iN1FKYeAuPbP/6rI6zTeCJ4KQg3kEv4rAgN0LZuj2iqLASRD+tkPvh5iWSM9JLTwt/1PsGhSyE2
2AAarY/cSxPL2kp1zs9T9FgQvuisLrEKf+rB54YSPIppS5RBWrKhL2NgiXurKgMzXVcb0nfl9ejs
zWeL5y8W4dN/nYh4vSQ8QA3ClbNjciNdaN4sUhbB5HHPBiHZIuYhe7wJtcYmpFAHJwOT44ReaI+A
ZeZjFKhyuwbr53kCqRHTjKtGx5Z9IF6R8htVN1MUjltkOE9v6Y03OPaF9YucFgMAed+Sfd1rpS6p
62QL7jYfrqvt9p9TwMpj7ELv463skOQJBxiw2socaribOkPRTvhzZWo+B+2isdIVr8LQzJu3sZxx
4wOJw+9bD5HUUbZqzUtJeHP/W6RpdR5H2xXWyVcPQMTYEJqxEKiVoUS7x4j9YUeUbnzFS+PApDpV
VKGd/iVLnsW5UMRGjjRBilBUCheZ6kRrLn+9jB1UjR1fuETC76XgALKmlxVA/y+Z7V63+0z+UXnI
RBgD/UkQqJlYNJVOn/L1exX/k2m2Ue2LdOYSs1pO21ezTIm4jSxmYCEyy5sq/5US3XtB2eJJQ84W
2TyU+ra229dnhMb4Y6/umRKMl5fN7li7eu8UiEBvUOtk/VkxMHnkPDbpNqgLHNMa5D9N9sho9Mg+
Fi1C6dVexacrgRuoF1/WNeGGGdZrtSqOVwMnVHBhQFktWngi501czKZb4BlSY42ewJkrrnXtMkE+
0JMFQBf+d4/5/0jG/9/iBKHRCJ8ug3fu77fVQE1/erxmE96dUJkxLmH6Y7w0ohnUo4sT3yYO7Vsy
Smhp25TMizttg0wPKF++nDwb92LhBvCeAC4XnOSzMQEk5fCp33MbpCqrSdOirHuXufh81LrdI0so
Cx/Bi6bP8FGeJlOr3WwAFyvu2f6/ssPJnAOmCR1zvOIHjllwqYF8RxK+vZROk7zGc70CqzjWiqRV
TzYtRx5ztHa1fwdxDrRm9JyHszzFbpupNNgVqpZsxwNQx0owAs5niSEPLJBX+JhNgYkwyRNo8P7t
weWnv+ftuEEGyCXSiavo73l1LiBEhN14aTmto/ug/cC5cJRT1FCLfV6v0tx+/EKWJBKaCWakUecr
FTvhc68bsyivLWHIv4dQ8t4PyKTqo2TxdHH2Fqy6bQdWU1LlXR+SH44tL72SD9glyYbqf0yNYT40
axyAzInqhn+CTFFdmW8M2AxXtqp4P+f/JctVVL2Wus/tE7YrXq7LTVdTgEBapuQFHdWb551l6HqQ
Vm1mTICxVWjdxSb8Tyq8wEJ9tNICcDMFnsrrXemaFixpneDJCME32lVjX6gifdsOPasvx0WbwFor
QOxQFmL0LyQvnK3ry8dT8hNAh7wKi+DqOxco6VPYDqDILYWlYU84YvH0xxbBp3DDne0b2vmcAF/M
llshuT6j37oSp7UCtQIiny6ARy8YyfK9N2ctw943fiFpwm8xHreSc254FiXJ3V2+JLEP6isaR5MT
GqaAT/TB88tqOERR7Kh3jD42lp+Pwz4oqtHdG+nixRV8hXBl00mdZ76x9/P/gboqfJk+qXiEhcpq
JYdaTgfwW5GmYpmx+QjvOosty7EvRh1NBUum2hjVyYQjcBx3pLzyMOIAbyM+M19r8PT4LbjN52Hr
9lSNiUF1v018Jr8rHgS34R23EwX/KyYA1I+/eSP0TA8LnI1ZEPbczLeJCQuYm5xFusfJNYK+a0T5
MrnLMNHL4QMn71Ty+NGdH0eUvb2sChHoI4V07wzXZlHHwVk3XfHJhHc9XFa3ZEu/A334ezoHJI4r
S0+oEWix39137ih1O+l45Y1LRSz4IQHgn5o9mXGIHb7ttfZ8KGPYZ1BckRLnIDxDEPLGGWauzxQK
Vi9p14WrXBwHsIj+M2WbNsBxVVLVIZQ+Y1UGbZiFg0kPcFGIByYrMxiSGDZ1kUMmDHXgBPQmrthj
cCqMxCMkyJwByWrSh/Jk6OSR9rpRdnFvwhY1gSxR+2MXIpaOTlYk/yCRVlUiSvM02mqwLweYCfTW
LQllqobEX5B6sdRWyhfUZlt/KYGKwy3LxK5PCtGVH+GSNi2JVPXChBgsAQv3zmoEmHxWtdvCpGBA
zuPoT+xIielYHcnhNmelxoBHTERKQTA1TcXpqnffqybZHPtlhaTc9IZsJFNAK1GBTelSPpb26m10
9uUpKhrxzWJzMaB4Es3MNq8WFVRceMu2waPoGJSMimqL48d9ibDA2tV2URkV8s3OTw6MhO3a8j4h
naHxhyaYIbsCMZ93sDv+/irh12mSQ0naGB+xARPE8ru5rCMuSKFGgx/Y1qq7gDij1n4F3dU0RI6D
fUjYV0NvT1jt8oXO7acbLzmAxbuGQgbdel7ky2zhKZZEmyeeEQCLh57y6Re+m69IJeI1TBvZwa0U
a/oWLjYvjBqdja/apW31rqo480qUitBEdXhiqWm45tjdU2UeB8LMxzw1yrH/jpeRo1HBUAnY/biI
ZoXo10BiPhJgaj7AWj+cg9HPHhQc5wD4B2UY1apECGIci6DKlV9HlNa6Rj0nE21MsMLAhKjsdjTw
WHG6uC/iEO5VL3O8kXGlmyK6zM+b3XpU4Vo+Vju3SXYiss0lEgGhV14O5N9hJwJz70gnJ3zzhnrg
SE9pNquqSXd5tOGbgmLw7Zn3c54V6fZ4ryFG1WyBvOxL+w5zr/VN6SN9+sYONRB1ECPnAQyLCrm0
9n+PF56a9CDVFW/zjbyTioYx7FVm1XR2m00M+xa4sTqCPbsaFJTCczPryoAo80/DaYSbwKU7Rw7f
9kOjuLNj2PZedZSPrUSP7japcEtlCEMOdGh/yI1PEHWD+758DRLpqqbY81pfGttkYClV3YiVUJKP
CFhA6k8zvCcSc4qWZGWKhQfJ4De/GqnFyQCMMUtwi2Rnz2mb3ZpjVoNGrbPhurYj8Ju7Ok1BrT9U
QM+3NtlvwrAgUusR+zravnruYbo7FPlIIQjR6rexD843KBnoQHvnbUSMCX1Edj5ntmIlmhE5BcSr
PFcfA2Lok6ZlgD3b/UaEp5qmVQz8P1RaB/8WeqEW907bxo6yECjeOVq1+W0cyOOrbiOaiZd2WU8K
yv5nBDGY13/JRIHorD6UhMBw5OWfWWNezrmU2YVBN5C1vSOgAssgWU02RTvdxYFg67k5gW7BtCYI
lJO+TTeSNhpAqZ/OyHRLVuzY9HXqKG9gIXkamEZKhtM9wZ22LMjEM07Lf4JCKb96b28Gly9o3szH
QRfPFS2az0DE+c96G/8rHiu/6+gAah88GvVKIEbq9us2AqZ3UlhUcKLQ6v26VwdDBt4lbjJDqVMF
jnilYVr1I6lRZ8P5pH7rR1J4MNOMI+2CFutbnOGDm8aDRI+A1kOge0v3aYautNFIamThxhdhyfJh
XfC+Hr/WgirWY29oL+DKuBrjrfipSLvf9US0H0+7sKZTmKr7TUrZbKwBplRG50kPM5jn8Y3kNlG4
4j3MQGadrSoqI9tbh6NdSEaFris8oXEMvCtLV3xifv+K81haybipuPkwqYTgB0UEFzzcfbEJLpUT
tVSBYlZgPEUFoydpL71LVAdiL2qdm3F+gKj1MUdTP/F19Rq8sR8vqpbSsxxkMCIyNROPupft0X5v
4fBnRyltq4n1f47nNTmN2+Bov1Rxg87lJwoO7xZURhfK3r8B/VEkZzpuheglQAilGOYAKDJveNxT
gvaRX+J/PRnCDA1l3GrGGhDnIsdeRgAoevfoqLx1/eA7BSSQxdl9brsNMHDYUwxTM++1emmrZ6z8
CMZFrOkBseTdkCJo07Y5mqub9Ypu8lFG3yzdRkbgvLefyErbhpoQx56eoZqBWASNTfGEEXlt8krf
HWnJCn2CA9R6L+5ivxdJiK/pRbiWwlWI4zFf+tBfbZuuDbFQVBRODXm0Va0Z8E4WDgKKFkiuJC37
iJR2T2JtwUXUH6bOVw05w+C/y+QrlXyEh2McOPb/bU6pqr7GA5chnYB/7rDc6J59E73vjQJfmYj0
vgIapopzTrsfhV6LsK4/6ZN3AKPeECkC7NHJw3Dw3HO5dR6flbNEGdQUl9gqVvi3V8OGY2dpDAZu
AUsz8MlgAPwo/YGS6WkHhXbnC/olitwQAOSpg9m9B2kleQ6RsXDQXueda0q9hRsnlKobYHYV4Y4p
QlynlTnl0Kdu2sJnkMOHhawwE46weDU0NXB6yYiwvpoZU9xHYIIJ4CNUnj6+3HLlNYxhmy0OmXjB
e49rqk22v/uxeefx32JH2G4lavnV42X7hsIYgLOMZw6Y7Iz1J8CahEM0DocsB9AEZHIw0XC57eO1
2GixkjVfirACvoJ1rK/ALM7bKcFV2ooJlx5yGi2B+AGB9iuuf6vfggGqyzqpC9Wyt9ZMEekzsAAJ
UB9YRHHUXsP+3gkkSVJ3TzCtNBZlJhZUq+4QiUxJ9RNmmSVxaRwi67L/4imBKsqY5vS7FQ4v+Qy2
S7cAGqFClcIY+IVGhxumMm3QA9GgVU4Tf5uQ5HepLoFh7YiDozeRsv1VFZ73wHEtmCtBWPlP0q+d
3w0pZRF33HUHXy2o4V3H5ZnzcCSSMbENYMVA0BwEjg57HS639WAXjkkCHs4mBdiHovQS3IHvFOpe
gUT1ArcCVpNpFS0vkso/r3E3L8HLPxt+dFrErYv4obCERGOSDZJsH2ySdUVrgEMcKdwvqlP5jFPp
Qqo+Mf3M2mm+4vZWMIOhSl/nNETLw0dImSRE54FIpPLwSCkkrZiS1lqWYhmxxtNGQ3UH+A1ocDNz
AHVCG2oopCObEpGTrGUGgpknxWFjjx4LZT8OEb8J3dbjkKYFg3G5bGkXL8M3kkEG3zf2MSdnmTzQ
MOwaV01lkZsCzAU+f09EyU3N9RNsWq0u6OdoSFHOzGvSoSR0AbmayltsgOnN8ZAv8HV26mHbHNHS
HlRwf8MClyxNWlBTL1W1azWKUyc5lzDCiHmu7l2V/PTbHZgywDh6R9fQYGvznPlTyCM0FHaILXAz
3XpF/l3qClkJOy7zSwVjy5Ed1j8Lyu/wz1KSL2rvs9oB5+yrIsRvw1lD2S6aj3okns39ZEu9U0GW
oQ2aC+JtdSmUv6rWkd51AB9MMIla7l/yt5U2YaykfyTBwMcMxgxilu+LXr8ldlkuwVSgrsxBcj72
MsRTOtGFQv8TckaGAhloT0aYuq75pbomfzD1jtgwO8LVgP9HEeblt2tSIRS1RWeqB2GLsvSgqWZK
y9b772732xuS68ppezk6rY8xbNTGukw/UTLy4Ain9VFX/VNTeSdM3PRx4KIsW1pD4gvYfLDJ59D5
GIXMbpaAeP2FGQUAgbmVmAhwAASmNjTXQe9PhVN8NUX8m7uJ6jXbGpougYZuus7fV9mcAUqNrTE0
3c9r2LslcwBrcyf3CKGIOsYS5oZ/L/ZNkSWQFFc7xNrgdq8Tq98fQk5t50B8W1SLnAYr/m9s8yhJ
6RXuL7YYKfskMAubURLqWdbGieEEuzE6K6/POv1/q0qBITUffLedqfjj8xkJXxfc8VtdLvP67yWq
eQXjaESSInTl+4i6UfWdKdtx4AinCOIMsgzSlHdzsjXEYv1aAMX5A+N7I264/Mk7y3XWBf00AN5Q
681xGiUK5OeR0++vDaJF/tcqCFq6QNgsgg2JE6mUYRQoHKWGl1zpBDTrYBFm7Pq9dlT9EK2L4W53
Sw0W/GrZFr6VpGh9OPf2XjhkrQBoGefxNyHn6HV4iePn298ksTvGANZs/tFvHrNBcXA1rXgWzwXT
W4fKXmO/kEOc89fAFaLFPIpHHdmkFl1NX72PSlbjqHuhtje+SCm0KHONKouzBNnU2OSyfK9RYnBf
VtXn/ruzQ/7jeCU3sgNpAnDOgItrsY5wLg+cjPOwadGUzemjGcfIEHaU0QARjE+YvakCtHbUFE4H
EqKzg3Aro7d4GDFbCnbMOeaV9cfc7OLn7oOImwkyzNTLtVcO6noUf5Ljo+D7jYPJ72hr05fPRMCF
W56auhOn58ZXuYxb56uq3s6KppIGTGqyQ1IBaH+AW0Yi+nLJsei1VVBz2viCW9nwMQvG5p7GW/tX
hFmOfemi1Th68rqio8OMxxA+uM5u/j8QH1G9RQcTMRISgDg/E2vRUqkKi6jiR+sC5oMpHTDT2zu0
qU6bG4TX+EYMJbKmu7r/K7xCGM3i/8ij5E9bKOk+KdjEJg6JvkiBmNXFckvQZaxbAU0kqG37DIzn
3ow6eepyFn/mgfxAWz3ACTx5k7OI5Hpl0GvyZp1yfAIjnHdyi7bAMck7FhL8k7y/BlYPwVKyausJ
a4nw5hcfHnrDydfDInf53919tD0Bv5TaB/5hmFlv0bhZduLdMZj1Byhzbmshcfs5iRapjbQzBm0Q
6Grx/3HTCBYugD/yfY+7+vKXuy/DxF4uKd4vr9HdZHLcBlSH5yo5zad1WtD3GVagg2f5XB8V27ni
PQJ+zoBPwe50CFAuU090ycfnEK7YplGN/CN4NtuaFM3e7RUvFJQWtn3XGGdIStoo+nJcFQcsfVZb
gzyEGs/upt+OuBvuDpOiF3DHXDt0625FxYGxm8WQiOOUIXFF4Dqw4y/Bj0VhtWivBZfu36SuTtVK
CGz6G+QAp0Z1EKhCg74T6b+gzKuAnJzE6Ll0hmXk5oXhNKXhr+lKK8Fkskb863QxamuFeqjAhu8e
q29H2sFRj7cRAzOdcP9vPKtcELhKjNED0sePGdqdMmeuOBhqUg8aMmIRhznaH/jEh8lJ+tvuJnNK
qZqt3YP8h2wGvglAyjPz11EErGG4rMdre8/M5C47u6mhSej3espFdcvE7BA2TklIekEDWOHB2r9D
lVdjFjdJ9WhXZoQkog9KbbQH0CZaDpA4W7dDzT0hKidVu9/yrsTgiNb8uxBCVeRopr2c1sKJoDwk
+d0emJrNX5sNhLV5fL+ugjalrOItBXZDo1WCqaY0gKUzX7bgfe9WjPRDSxmKfTX26zld33zPDsxj
CO3zBESWLlNkTmxXGUOL+PbRUWxMUTYphKnps43FhTYyYsZ2ZraqVOstxdn0/HVaABncbTfZ9P0e
DrYbsjzE9V/aXa1OCkDVGfEq8VPV/ee41/5ThTG5VDMB4KGecUIsylOJpUkworEkzTPLi4g+d3Vp
8rSIjn3Mna4jwFfJ3KyKt3vxsRCb6zQSDFGWESXQaHwFnjUnsAKh/zIwhGo0s+8yPNW5Rr7fntuF
fu9WctViMG8Tvc2j9YbDBk/utcBAGPOcIVTRo7Wm0DBy4dmQiG2uUpCTNS11NEnndcA5PQtLJQe+
02PlEeNkqYXfJG/0VxCeVpo/O4ftlLiLN0TBBuY+JG5x3TGsyhi6FaoM1ts8JFnWDfYpz1OiFv/Y
/W4VEkGOL13UBg6Sz2eTreSn81j0TnrbWiGShssvVDs4GleKzJWujgnVYwDG54gkipjhEHV6w6vr
6IZT/nXBKGsF6T/g0DZIy7zkZLUBMwdEigREXpLrAQXXEHXQJ2qqkZSsdJ7FsjBc3s+WyqvWOQHy
/SZbvRWoHDhqASYTmtAPs08fhrQJme+yHR0+hFX6bCMgR3bQBkctxD755Q9fIyPdej4m+q+f2Ux8
hPKE1TvA8wMwjB9cmuYfE2SSuHg1aqEF3BXlr4ahv86eq9MbzS7OBDE0+EwnBp3o8hwiVp9Mvvhu
cQduey8DRElQcqZ0yX4qwHMP/HFOdFH0GzzmJoT17sapL0ojPPGKuQQtBI5dWvJJLFXUmoqYNbUK
pWJFflxlR5mLQInNdUoqLrOlxsRuv1DYBBRoigRqQu3Pvsozlcu1s7TZJ8tHx/60RU2/on69D36a
2Gb9OZjGOdVGoxMGbD0QMAo5f0CDGbHjAQ9pquQx2eXxSIDe8xTZShpARBQuHLBV3NQ5/EZMKzAh
0dXaILg027xE6qr1DgxdmKDNc0Z3pTwYGE8et5L5lU8epyf0XAa+3lyhLRml5t1zy5Y7EJxk8TdA
77o7hSTJ3C9tVi2q+BNHvKjgSNZCkMk891VnEuM3WBAu5W2cSc1RsdIy5UI1h8ODWVuv0Bipm6LQ
XVB8gnGK57KEwCOo2GActWVACqQMlrVaOvwUv2LPjWtCrnKf1lcT7UAg6q+QEZov+8w02ygP3QFv
9QyGmETCn3YpEauZ8VwovsPG741GGmWqA1v0GzINppT0gYoJ418/ILoNb1RwnurZP3x0iSytLKw/
yxFZA02xh0lyiIvCLv9P2bcpl8aFY4VuAqPEgeAZ0zZAxFCC//9woYOwo1zK9WWxKNrluoor5cS1
56zHJfR4J+t6+NfGN63HmytjO8/M1mdcuZzUse6FnxKYPlmVWVxn7HZbHFC9CKIYVKU9CTlOwzXF
fAydSKF7TacIIZmel2338BU6KnmIDpTVxIPG1UqsKX/f38FxwWNicr7h0peXggMqT3JHD8l984DA
7BPc5ytDyEdDFnLrej303/FTj6xEpfOAbYK5KdwDh3MbOLch/9Oj7GbMKpYPElkcsg9vMB+yejTP
uz2AJcnNc9eKDhCzqIDPJyejrNWc49mJNpwfUuf+ZwA6qxj4u8U3JzEWsJPnV3Xf5vTaP00O1SEM
kZYM9W5tW+c38f5W2pw9b81UXyT0ZJrgV5SDa37E8fKuZDInDCsfN+qFvj9JQJSapifNQ3WnX/gr
M7zTgsAcUzr/XYK4sxoK4z2HeIDqbgSusRiE8c0unNMP/e85++W0X/HACHuofB9g82OTBp6SBu8k
3ALzk9WHTTv6qJC7V178HnN9rwuKHP2hjNcRbVKnXqYy9GmDD/SMhg0Kxu9+lEpeMzBgn1b5+PHE
2GIE8COXApEPu6oADJlGzuQ151ZHUv7ao/swcn5ZR5NbjClDE5YWgGJIRZ5BW3VnqjdXMmlv4hRT
5YFSLnvUmpduoUH+/cbjeHvjPEpXP/YSXhO+RLfQhyrNxaJ4t0VlzezX45RhX31tKFpQ93zImHaS
L3CoGRq3MlwCtffxCPs8oFhkE8pF32jz6fX3MfhCZH1T6FV9+WcFHVrfY/CLOw3tTlFjiGIAU5Zg
JhtlyZ0nXIPrkwydPGEQfrbtGcFu4sUgxbgRh1OxUKOLCvOJHWEQPUshnEQCI+yxZ5voxRwmlGr6
4ExvxR0vnHMYj7MNgvWfIe1T3LHTOIQnX9/1JvhiImfo4b3OtxsbE5SzBYpH7xPD6y1bthvMfv18
RArrAcvfOSXOx4e6kPw7SOp3iihanH0TZ/Bkf0/NO7kKWokyvfDadl8O16ODFCRJ1Nz9aBj2brKy
6XdQGx5kedkIKsoZ238udB3FAkf9BYpMj9ber3LyU9TbKeeYwR5rC24N1XgcogH167Nac5VBU2k4
SOK8H30H0WQbrx4YhOw/C7wsTW7GtH1vtP1FWlyoqiApsxb8iCPnR6n0CwZ6OLPcI7jY7AU+0nrV
5EVRM3Uw6/gyW9PJa0XMo6aQaMoSUQA8n2C1EEgha4p1gDttzpk/aw+Lwb26RwlgRBq7/C0QnVz2
NWuIGwsnS974KVqVEn/hfZUVkMfxENncMV1fHpw2DNKkCZcu9SlXb02RlXIw8ttLbiqbl0z9Sp/X
vtxTKk1WpQLcPwI46mt+4POzrsOwTy/idVnQ4s8kNouBwKIuL/C8nNATHpS2YIlFCojk0dOg0MMO
4Q32U1ZHzU74TkR90Z32LZupJgLRMO8gkZAkTB+wX2HDGN5ris35WzID7yk/8d1fFtnECCNV2rXy
dcZRMz1BvcDVlOVk+YCZidqYYqFZdRnJcl45rIjDH8Lqrps2dVxomU1xVrOdc/qPTBvzeNLYhFPP
PZDe7Nqga3xt0YNP/sj6L3iXIq6OzjZ6teEnJjwZiwgLEzReQxui+alnAnyMs/wdudENvWrc+Mwi
wjcEFbNu6RsCBzGr8hajdNi9AJ/A4YJ4eYSwIlyvmRkV/bYwXW/qAg65hh9jUV93eX1zYas1phOS
+mKi/z6fhFwGeCk0BGoVy0RJUPBhvWrjRY7ouF3DF4+M3sajDE2dMoW07UqFytV/VfPqktUbRc+5
rhDMdGP+1Ks2/cDGPR2jQ06XhDZHXgf0u/3BV9QPkwgQQqQUkxgtsToIVv/EK+l8d0SdoN9OwEoy
Egf8ChAkqZv2pWVAdCueNA9cYkL9N1DFGPvsX58HkagaunTaNCMH0tq+iEUGgpa/6kbZcWMYhPFW
WfVBzct+prAkpcrH2bNxxSrC5NWjhVuzU3ZIdVGd9AV5YVJ+RqQughIZ/DHsKY36RReyRAPL4PFv
5aI7Q+69wHNLcbwB3Pn6gD2YfDRiPqAAep3kLidYLypgos2eG5rPYY2OjFxMnEcZ7XhVK5t0VPk+
44kRtUAAbNG84077FvoJ6d/qikm6WTNh/Niu7CrFCG/TQbXlN7OtHsO+dSlDxD0L+zIyJx3tNSuG
kqzeibD0aQAYMHMqi01cN+mIqB2HUPBbgKxoSBN5XRHNidoJy4wB/OWQzlI92agX238+M0Z7c6uE
f1f5uco0dv5ymCaQFRBIlUk9hpUCcnjedkpK0pYAuMUygaWrGKB0L/TWcytoVakLLetkg7sHDhB3
+K9pZHzfwDmYdU7s7xdIh8jmC02LIveuam1x0pJ21uGCnAgKDSsa3UOD9PqCU9V+C3XDqytfpLKx
CAy2QjZT0da3+XnTO9qbiDRW/D6m0Sxxq6PheDZB6abVWaZjO1EoHeul7I7itDDYOZqI3t/iqlMz
yoZV7Z+5B1vRPRgKINNKtJjDkL2ho0geOL+HUbnm5X5GDm0Pln14SslYcYqLbDjeI+/wvrA5clBu
/sKls8R4GYgf2+pxOdNp+lgUSDat8N6OUp0jaPaIzFak2+Ecqk0+dg+JOnYFi6rtM4RtFldbt6nK
uU1QtWlJeGUKtRgrQATijch3KQ42wSUmz1p8N250df+9robKwLL7mMcouV5qRcQ3QPjMif6KYQzq
upBQBqfibb4VhV1GT8XbRevGI4+JVwW3nrGua/IkdoPTa2gEuDf2twvpifT/nGzF9/vt/yBuuhlG
6TklogF5rkba+XjxqGP7Y9t2Xi8850QzHhGr8vUbPKiJDo+MqJ443iVNneVPIWzyDSeD/gnNP5u2
5BD43/LskM8vU95hRy5c9WMx0JhUzqPTMClNgzzU+QhB/sUdKOvw8DT4+kv9b5fpDfKG6EJXy5jw
qpN/KTEHQ3aKJ0CKX94IbUDMMz+fV1W+IyaIbLULZU6Erl9zmsooeFqndVV8HLFaKHobyp73gUfQ
7n7rKy0mTnPv3nucwiprOZVHxqjIb1kw2K8n0rfasu1Hmhp1ii6FDRrd/k1w7zgMSvFsP+wF9GpV
c5rsbbBGO3CdwQG5Trusn7KU9L3sTR0GG7agYGH7X5aa2zqQXNNUOpUsNeROMyRG673+T/2l1ZHY
jlozsSQzuU2j14zo1cQtGd9TE8vjw4Yb7s5y0JYZWcFpUmkUa9Cg/UA6bUsjsfOwg/zsHaUj23rW
7yEJYtT4KrN/XboJR0RqaNa6/TrP7lSFsvfVDXTB/Hu5w58ucyVLlX2i+aSywNdvczdyvUbSbkEu
jfbay6tedwOvfn657CIOBVHe4S/3hFCdsgVT26yEr0IGld7Xcgtb2BliWgseN1rPsJpbDFaSwPWi
A8KGmvccnzfTkdi7/sssprk37bl80zedU+UzTtZgrn0GQFvPKZxbo4kHBhaHCQioreSSBMLjSAbv
P4O8ry+mWj5Tp3/vucEhM5+UpdrfPPDn9Ym8R77qrwm/Cas+e6JcJbhMQpBSdrL6LPEA238lyQvS
VoIOkfbD/hlHn9qTfde39E/6zkQlunxy2Rj4RYhF+L2Bue2jrrzisWeX+A4hyccciPyQMQcOzImG
AJ4JkT81Sq8t4evUWy7vt0Rzg331dz3BmCWpcI5pAeQrS9tHlnzmF7Hxo+Kl9ugwlxC27CaKhuLN
G5nxuV2RqsmhiML3156sAHKpfcpSpqvOV0TdokG/7wuW6ck7+xIH+pZ7gqhGazzG1wg3Xtkxb86j
COYpk26g8TFtZ5qOAzmsFcoZDII+Q52J+gSOaodqSElYewHcFYQNTS6diOlj3reykLEbeHHRxHvf
sYRlgTh2M/2wnw9mFCFD2d2WMIeCg+4ohErQp0y5MlfK9Tnn3+ynlrNi9JbEaG0fNzF+j+G24XIl
p/ygOVJYFZrYEvRfBfLUC2XmCsJbOt9DcJZSkyH+dxku8SVkh7G+6Cj6KjJKE9jwZ9ijDU5HEJcs
okd88ZrDh01Cp1tvKZT7O0EpCJWZyYt2H3Nsp7YJwYxlTab0b/4qxpzVMFSOO3x129zz5DGF+7eS
CUQhs0yXwAbucx4BjVwpu0ZCluahM/B6T2T6xrfa33tnaL3oS0iqLBjelJvrmnaWXnZgWlHVgdaZ
dVrIJUnx5SpAtxiediyJ1j1/CR+Bm8Hx0UMPL0LsfiHDIFkn/7hgb2xJve1mMyul3N0niVg3iE1J
nXuHN/Xqg086G+P8/HSNwayre/nxjErJIdD9roOnyDew6FttVrriJjd6Fy2taA9SkwllwKK+aqYE
GcNzdZaE07TUH4nyDy+YpuGhVrWHHk7cbJ4iqBcitN510kjNBEZ7MQ/dk6ipdfJiRKE9iWbWDq6u
6spJfDF97lkSq+82raHZUkvw4dZXDjSJzukAIIuA9PHzkrKQLOaqA9liW2PaEaXdpVBeCmydBRjY
H0r7r661gsK84keJeD+sDLmGn7OELxUdplLYUinV/QdUJWZZntDcr1fJhJUQEw6sYDrGenRKIYiO
Z9NnppvDTlRmu01npQZigzvN5FG6YDb2Fg5NN8dkR4V2fWXqzmh8Mx9C1IumS42mIvbLN2dq+BN3
SSXlgiFfBtEUgD7lGay1njMJibgDdAp201gB4n2aX8iGyZ7S2rPInP4boPxiWyq8mEq490AEATwk
Cit+ydFrqCLIf1nNp8Lk7+IO5CxBCUk4lHtQKsvsmmhPubl0yAAvyfR03FJ+nzeYB/DKIz+Hnhg3
OiKEZzpiajspqs/v8/wIhQ6ifKNhSC32PbvxoeX/lpL3DyFrhB+gXFK2oEfWTdhrK5eZPSgYcUJE
vG2zZQMEmb6i2+EjEnSR4WrobBLcyPgjWuSzk6iY5+LpeKyVc0mszp0Iu5Fjtxs1vUsyvudBFMIo
DFZEYra6BgpOlsVh5YweOKrE/YXoRhz+y9CpqOHxxiHXqQ114WcdIWsJQzzFsyy9gpFou+RzFquO
QJqMaVt3uXwW4giH3JykDxnDSO2cq5KLo126cQnJy0fN9gnb31pgNb14BabVcMGy42Q8epqSkiSP
y3Ta062Gybh7BhKbM8dIbBb4HEricn2pdmmDhS+M3ZUrYgOQ1TR4Y6Elzyijgv81T55TLl9g/ftJ
6cEg8roTfmW5PiF/y6K/7N/d0pOC28StlsTOgGqW0ie8AC0BSxG+ZLenDl/GXbwsaz3/pfCVmFWb
hvfB6xT9chHAhqBy2wy4edr8Q9X6lgauRW2rGX0BdF7lmyDdX9jXNRVNCPMFjwd+OfYcy18b1gDp
KTQKKRp2/p0ZzszAdy/stecZhW0rWOisKGdtxh9UX/vL8PpdERZ6t9dqvplW+8ZGwe8sEi7yUwWb
MDk9TlUcIcTcRzKy2S4N7ELANf8lsj4XsPwhausIqYz2TrNnBf6DQIrhcnAjCbl2kjXVNFUR49O8
tbxEoU+En1GTPqbNZwPP+e0wp5Xpy4cd3Rqd0fxvT8J9lnrEKXtKH9NndxFKdJFW3YxaHvh0k+XR
RMEV90b17IniwWf0B4ne8px2ed/p7ojI1WyYCK3VFGxvLajDYd6Pzs1HD83/fQHfBe6sMbP77MDo
/cQNvnwHH+IjTFOOrm6zDYA7lR3WrEV6HUpXoqjN50UddNdn7d3rdFCsNOrsatt0q/YNMlNwve+S
Wf7eFi0OMi8csey2OX+uQ6NT+/fhuywuko/c5MuaSpBEyG1plu3USoNPwK81NdmHvekVXB9GhXiI
1QYXndgyKUpIHR0YLzsYBSXb38AmmLbT0qcYncsL52HTyVSWm+FokEJFGipgy6oZTUawns+nrZxR
ro0GGA30FCtNl/X4T4N3mQ3Z9Km6CBagF2PvKDeNuWx/o8u4Z/uni8IvFJIIU/RlaxjNjloSfV2n
mvHYkgjO6lZ6Wnls+IVZizB4qrF0xborbGeepCXDNOyWLS2v4MqqfL8G7MmxOich3Jt4NB3J2pBQ
QaMfslG0TEtk0FNx+cg2rDlQxi0g13X5rh/+ohss5alIzB0TwPMamQ8p5M10fVpVyt8rpauKcfjG
1Dd6eD6DBf8iKWQcG7i2Gy6FyYHaQ6JyjPWPRWQOx4AFiXqg66PthhpyCLcDy7KNK8LSZc6V6phD
ol1+sFGI1ttMnYsdJNTSODCfwL4c74KGhU9Kw1s13pEMcGcNsktEMaHc200NsKZMPf5Z8Yzgep9I
55ZCPhWUtYMatWfr1ItWc6OGQd52hrRWZhfDAVwKomk3HtnL3fdG6SHsq+o9bTGM19brkwQDM8kv
ntG+dPwZ9qzChZjoiq9b6k3sWR55Foj0FcwhJohpm8N/OCuJQTwE0V242umc09R5afQsbYmmPDWb
rhoz1C+0NuHYyjBNlLZlCrjoWxzEuHGmXcRBXeIKGruExwlCMLJzGmeA6BOxgGTnFfLF5dTmYrl+
Q6aD8OsbfTv9xELua/H/0j32QOw4zWkaVBIOYvPmJwvSOUY7RhvI9js9NB8Jcx8oWFG8VQWxJ/d3
o2QXDLe9viEeLULcAyvNaBLyXzjAcVrIpgOA7gbNW5wOWHHvmhj12ECzXpkWP/bClDUHgF+atqjY
TVjHNqlfWT3wAcABiiheM7NwOIPUlmb7u7JBOHxIxMu5CC2WBHbEUZMSy8NY3U9Sz2iK/jOxebHK
+8Z4GhzbFvHgqJ7vLnGkcCt+3amDzDZBwPe4PAXUxrUz3rcIjhoqA3uHaRMUuOJZCvNGgyZ006GG
bERDUuMaT4QgH0AfWYEe9ie5CKgDeyYRsPrbnT5FT/no2r7DA7AXCUy537qktia/cqd64MAP3ure
GlgW5OWJ1cHmTpSCCIUz8/4hvMBL82MZoEspOfZ0oLl6qAhTn9e0Gm0YoEKSpHsU2mZ1selJx8ui
x7JpGM+as3kAyWktwVTZLqffz0HFEDRvpAvTZcRcDCac0b5OA59fzNRbww4iYnw8tU116UHYzrAC
myFA4hJAfy/7sB2CT5gpu0LtExumq6rSqPOPm/1s8pKdYBaNVg1dHE9Nu3xhPC+6KH3Mrn0Ne7iD
hwD/P33nY5vaBOP+Gua0lin898dvaomGPI+KCkrTEV9cskg5sY9gT3Jrhgm3g913rs5qGbMyFjzT
8tlPHZPdPJ+6vWrmuFvD1kqMnoaiUphMyC4bMxtntR4bJ+woMCVRKPvA71loq5JOoe88zFpQJWUP
DaRmQWkHyQf5AmA5qS4piX4tENti6e3U0w9XQCOQ75gS3hpN8D7xwp2Wg3e6muUVWVzM/xxagwB1
fK3bqZhVjvd5U/BXol8p75JYYoGcs60LuxQWlEj+ZKBkYft6yvmuC/R+G+wahWodyqNkTVmURESg
6gAYjjuHQgK6ZOGQT7qHTXOauC5Obkzx8Rd1XEafq/4D+d4rKNcMlPEgvfLwPoTVEMHSk/hfxe7O
8lJSsk7S02/6gl+7DbJ7AH5nRatZo/BD2FjyTs74CK+QYNh7mJIyU9IdTz+Y8EBQYH/B7+8jZNiS
+Kk7uzMam4gf6Lj2WfDg57V74uUXvr70hFRdK2e6c9M3G7GEJECZBUBFK3juq/xGrqnNiQsEboQx
7LGqWgpEWT/upCvZQskdc/wMSVcGcwYIM6YjRjl6XtDZi9/+YZ+KpytLNz0/RhDKyfb+s+RWtmV+
K2H304BS9q4HAHgyVLdXqx5udLSwsHPC48G0gbT+i0CrjmN6Fv6b8y2QvrkCZrX30PE9bNXq1JHc
OTK2Vvyo1LHP3Cy6bHu0tKDY6co6KS6XZs/faPZALkB0UZ4Zb3QqqVaxM0YMnAN5uc7zn4lNeSLo
YSBcp+NfhPSW58KM55+HLnuOfttyFy230LIG6MmYbSlZDVCoFJ9DDNy5V0fCV+jdewRqGPWPj2Dl
RMPKHAJ6CfQb9KbfLFo95X51h6/AigC2Kt6q0GvQlXRIkAH3YyULh8/kI0OIwENedTKYX6wmsqwu
irp/cAiUFwILS288t7aGBdbUFkeYj6OuoIe4DSIRTT6jJZtq0ytVW2rnz3R9v6IWy/V+oMj2DiBI
bWjPhreviBLuKmfwwztrnqTrEDr54B/q2GW7ioJGjkmxeLZJvVpbe3z0HxI9I/IES8iVyQd2Isji
OjUKg5QUzq6Ap7RbiAmBc+MBabFxHurFUxmKAiBRnL+aWcNa5W3xc8h73DY7VnZYGhyBCuWt+xih
ePeZD67dVF5L9WSAqXyV83XaMCK+qKiiSx1+y1GFsbxty4+7uHaUwDhCMrKBfauywu63DFJ/s6xx
+XnkkM9T3tEqzYg8Nfrbjb9fdkbYxpAcw+ZF5eNQbMmthYPY5sKld5QcwAUwlRaqxKxWU9fp6PDJ
VL6/X2K4oJKzAHpy7b2CxiYLwloNak9Jtb9XZL7R+LVh/WtmO0tkZTM1wfe4j+fChlbSvCatTEHt
9AbWQ2Z9L030v/BEsW+6F3QKtjTbHv6bR3HmocHO+JiMFTeZXUBI1dhYobCQUMmW2IpOMNyb39BF
NiJrr9Of3OqqUs64uRh1yuCVOGmGnLL5sMnbxu1qxt3OMyZ14I7lXPsVUZJsdzxRuaOE72tIn1en
mbQu99Ozn/OvDz9iXRbtM8NRD9BuqeTFEZakuyqMNr1I2eNvOyb+wIpllWIIcl0J592bZCRvU9q9
KtLBj8TmKFmuWn9m/3dBOk6gXakN96cooOF9nA8gEIIFMKPLelOXSI57Ygis2jaLblUrto9xgICE
3m+YJO6WuetjQJ5br/zyscWA0EwJFtFOOC2wiz6TdObABk60kNA9E83Rm0YU3qEx6uHdysQaNzei
wB5kqsPMgN00EDeh7WXMmt2pfabUzdy5LXAc2W6s+sGtEc7DVxh3xS7C9tztroNFAWWMwRtAJPJS
W9JsktY0+9tW1kRvXq/ExG6R2iEXDCbUXwDLuLGuWZFY6gXTuMP1WnnjAKQVEyrPsbdWupsGOxTV
zf09z3jqoivqtMCc6bu2XwolkEo+B0RIvDY0L7oH4vSIDDBOYFmCiW8DgTM5WuyNscg0QD7vZiCx
iYFe9wLpvWN99JOkKrymbmwoX2qTFdcM4ozQwMJdTGFUiF9DFDZtjosz+AQQE9hAupEDDqxBQYpe
Wzu+NSXLJ2kSEbtjK9dtcuOdSWzS9vrDxsSR7kRcp4m6agnHQ/TaE9oVUT8RJzrNYCNg2k137S8u
7DDThQircs9aQPbkWwLU/W0eja4cnLTA2u/zokAYxRTZnEWsBOxiJOrP/4Y6r4pme1+a5e4Ivv9Z
Ij6DJRbc9+PJgWpvBmYbdQQXOzX9pflV3x12Fz7JbssxIzHzDjcgOufQGGbmMtEQjAav0HVD7b0e
XvcUjxvuHBTonln4sol3hIQFYd1eJct6lrA7WkMBCHzc9XLdQbS3ZD6I9n2K7NxMVTiFKI1OcjbV
mEZSYzdFWhW0SB3GJyWe40WrquKJICH75JDBVjWjbJCf1Ly7KpjkCaibDFkfEmYec4hsTYlx0oBr
lycrdtrsAdIn0vK1UwxqL6muBrDHOZoVWf7/3T6XZPm0JMjup6vpaxQOwFjHq7WJoSFkhUxbiee6
5cMjVIgd2NXYfFhQSLLUMJWUPkmYWr6yAsxWDWQEVtz6INUgT41cQA/3EzrlAR+FWl6lBGARY8e7
6To1FHv/OUuB2z5EDl1HGyKf7KW+oe/iSuONeUz7/8QsL0NBqW4iJb9wTW2DwHiER+Ly/6UrRtl9
GO42EahRMsKcuOEsRAeojEeW9TCWBIKzD0vi5tKWimHdwqKJtNgTVdqvm9i5lJRMen2HXNiWGlzT
HwNAX2pyCTqwwc8f7ijQ7Xslh7K0uyWPWikoUpCuuBP9borTO/dWTaOGQDMUwM+7YktCj63J8MgZ
uwXD9MiptYZABkGM4siFuEuWj8Wq0sxdr9ifbC09vSUq7/i3bzGWf+nUoxc3SHJ5v4SlZjXXdDAZ
2BFOBKfx4WZ+M8bSELpqvOdQEEVAPfuiC7EpmeFSRoXsLFGpWqk6slFm/1Ey/FbKu5+JQ4RtrbZQ
/ZzcWjeuGEylNG+cqrgAwRgUD9ln9N7qJ/RVahLwj//uSFMLnWEFQZkkhVrjFmf/d06j1zcI9gp2
nUBstjOvv6+z4ZIjTQL43yX2kjWjD2BGM0ceW+/9gq14ShvGw5fZiaYRBgeb4vdy7V8OR4dPp0p4
dMQUDjQLxQXPqPQz2lMQgqXqctsu2CFQIpJxbk+s/hwWBlpncKwlkXsyRF8eMpSNvmfn2gAinEFP
mxDXfczMTfadr2yxhcRzfYRDjGf5n8j4Z2WAuG5Csdl9xtoaC/cAp513Oa6GNNR1SyBv6xJW3eKl
jkTfqjfA83tg8xK7wdMa67DRFhjn6mSyLWb0L3s4kFwA/JF3F83zTaqM7POfKWxqhP4qas+HflgV
J+ETRbzUVezGpVHMQTrdX4INSN5lFlM3kiZDgl0gzwldK/wRM/ku9ck8hg6ZNCs8ONDv+UK7LwLi
ww2kzi11vqZBo8YhQoC8WuDbb5YxPeXGMhkuMflIRjtWoyrgbZqx+0+ZsNIesTK8/WsuM8yFJlGG
ZGtu93YU6LSMAIScioKu6Gfwxf+KuufP/7AO82KAjqyjCYt8dTsuhgL2zTJuqyPwLrzQLicPwmyh
YJ6pweLFGAc6HFS3T9mDKdul9LkXLzPPDy/WUz6kvg52H5BUGmg5OFgIqy5vDdHwnIv2ZivIRHu9
YuhsIVkDYkDAVhoDLD9m3IOIJ/Hs3GnVaiF4MZCrzio2v2AGd14EnWCiBVcrlDvbM+eQMVryLjZ+
r19K1+zpg/4ooDwWkPY4oYyRIr8ZQhrKIKQMwTlLtTeKdSxTAsGVTB3DP0OAO6MyXVUFoOZ6EtPs
O1p2BuLoZ8LHQp/SFCd3/VlLZH6Fzw86ZGvxWriq5o1+e78IcKzfVIwE1S6HGtkIqpCy/qHiFLvx
HVA+Bl/5lAls2m/9DjG1qWbLFY7gNCkJD3LHxy+0iAWsIuqActFNHmOBpUrYpcyrYcbV1AzCyGvO
v0NaAdk5bhIkwN3qBReRaZdbal2ai+FuYL4Mwpi690bBvcr+E2Wpg4meCz/MUDXl/re/uiHnaYWl
IXzyeFKIe18j15ydhCg0hA8wV1WGKRznMP3QZcI8EhsAv2mwsl06O017WWSGJjJ5qKy8ZbwUL/I/
PA9eqOOxfU7BEoS+HGCaVx0Rvc592tUgEMkYRRWTyuoeWx9oL43D3svo2p4spFd39lpuMbptxEWg
22oFBBzSaP8youlIhQZniK6F8elHDXNZuG7h4w1oPFrtmR70ZYtzCBiv43E2E7WOuD48frWGpmWq
7tczYa2DYRYGKcW+06ANO7G/foybwM54OFCTuuFLuienWO4+ppBuJuHTpnOmB2QQrE0zSfOlto+K
au2e2TCItZRr58pbNNuuDxymlg2qkTZlPHDkET3xK7/Xj7fJlGPKyhkmUlv3w3vkZblk1kxClRmT
pjhobWbEJ3/2mHJmjh7a+T/4966zZrt8ZLc9OZSX9tqAS+Fd2sJeqyEUpnIKtTvDMWPdq4Drf7dp
5qyABnN+FzKPVvFgtD61TAKusbSLK3gseLWHmbcYXEgtcy+oIRF8ivUburqrq5XsZZeqXitYea7U
b691eqG6HYn11jkeRXzO3Y8ycWS9DE92aK4rk1Q1dgYqYp89P+mvixaSDZxMW+J6ZLm6b96c0kKv
gxoLSrUdh4QggxBbXEGeUet5+Kn+/f4S3+kN4297yjskGVPfQ+elhVSyPJnhlpCdNZgboV4akXhy
eDzfGp7zFflECYU2QCsUmo9EMG2F6cS/BnXN+eXOTBb2V/CQVJBRfqnLgi9PYFVNOx+aJOhpxNSo
wzpcPj/zlxvj3NQdLY5PbvvHlrwT1IcgN9hg8BHHA3Vtx059rDnlscPGKf/exr+W/0B38AmGYqY3
+FAzyEFijaFLVJT+iLl2tIdJc3va6qr1K4nC4eRgzmWWT7l/r8WAWg1O8nz0GhBvzTkL9YK1uaC3
dwGA5c6xOR+//fgMHXuB/mXn3Ibv3+JjkaSTaN2/92rvJ4p8KHvQY2q1e+7WdwAPLgWRhqnkGLS5
yWHeYZweDy0qutVX0/I7Rh9IV41ZieFzff8+6mhjBoiF75VeDPGs85JE+sbt9h20ISJfV7VVJfFE
6R7uFI5Mr1t73UlHd3n15v3V7SUUzZlqu0L9JQ7nxzy3x0aI7tHFUBzkLndYUXGAJ1rVKiLJj0NS
VvCF4C9fXZkvFVCz4yCIH8Zj5IEWb2uLcYkvjUfvqFNAj9PBBgy+97EI2P925uwgKNRfG2cTrTrF
plmTk8Gch4Px5fuos32hnkuY3dLXZzQzfTo6DV/YjYDQCGIoku8eoC0AvDun0OvJ+ofKoQgJBxfR
pToh2OAuxGXpatErip/dMKrr6UkvvN4DbBG22dm37T3xsLF2I/CfOgPOGwXnUSZGGLjcUbWE3LCk
zs2WQndfrEWXGh2zvjwfF0qLd7o5dBInCqzQLANKKhulkE63yEX6yROAVKNLVeEBxzqOTwefSQzl
Vp4v0pQad1hJH7gJXOMfqZx2O6+5h/2izauRfBNXr/lq5EMKkb0dc6o7HqJP1gs8mfCXTw40lDy+
in7Y0sqVe02vWIiGeU2g3XQ8GlFyRGwFf+79MWfLSAQYABOoOKWT+lrG/zNVzJlj4o/Y41Ub/xO8
BkVCKzESLpGX7Et8LGcmQsw18wJs+Kc8VqddHgvwNel3YY6VQZQV6TlGMLWd335Vv4VUv4haMpk3
MkPfKtPhrTrYGFUzYPioxzipZoAp7GTZVSWQAYBG6A26HxWk+mhVtu39H/CKEi3OJ8XJT3GCZWeG
JJQttPEYZF8dvVvny8Uiboj+BJruymdPgT1BP/AGBBnZfRnBHfKCiqyR2cu263TN+LbT9U3bPLP8
g0sDCvqtItHKY8SMOmqJ1Hqs2GFGEogiNMu9USblSH4SOgGHC61i5QTiKW9+/Mw2q0l2WPnt9iWT
14HEYw/6oVtklXs0NcKZrwtNmXBBBPdQtkx5l+dvh5HHSgrJOVWb7otUZcmbvva5H8a20VPQRuo7
p/iT1k7inMgjrxUaskO/x5PUUUEwpCMhwdN3kSe5ZplViCZg6hDezzTtyWimbyZT6zXX29CF0I+J
nwcP/ZPjKItZNXd+eGwkuf8fpW93sDiYocPiBQyRFCL9C+EgN7ra376ZKS3uCV9iPIqtFZq5lvyZ
qEnMswUp4wI/O9NSWPS6+UYx3yEvltK6WlaEd5NKqqDsGl3pvO6Bi6mbYXVoil3wR+5iY8qm9HiI
Y23oKtyXTWB1fBTPW8IOhzqPWLU/JWeCWB/xpDzC++VtB0Lj+e0fMrgu76O7MJga+yRA9L7U8xOJ
eSQhQGhDVAo3Q0t5oNRw0Hsrl5gvep/ykVVj0NVB3aio42bteTrvkJVXNoA0W4PyA+s7f2MK0rEe
Fe2poV7l6P4KQM5x+aXhcJNYG6VrcyVJf6443B3NoFWGZQlXrYulfR8cmkfxgznItrNi1OQ+XJ/I
koiX9bX+y8YHKhOib2holfAL6czlWiSZUbDkvD1nt/gHgnUruYdoVESupl0Sl18SuIWSBbj2Ms/c
MRuCGSNngWIzv8buBnVr/M6YqJQ7NeIRuqRiVjAS17rZsCD9lHNUfHigpqTbyW6kh3Knuts+acF7
nr8q19f195Yu8QO3PF9sPWLa41Yf3H1zC5BP7dzvlNstFxs4Ir0XvaB6yCtzR7GQZhElxPB0HMlD
mJlKVXnXFeIn9YPm8CZHs9h9oh/FGB16Y5z1xFXXkKjwMkM6yb1E3V+7w8vHH0T3zJVqIpKTLxZr
LCiGmdbP+BPn4KOrap1opt+SmG12x1zWViS1coyk72mkI+kw9yGN2QjGBe275FgEOzs9XWOXo7eR
VwvCogOriWVf7RoNsTYj9QfV9xDK4MeU/zXogM54M3AlMakLeU5tbCnFPWpZHEKZ/Y1vLCD6/HIM
wCM33Spkn/ZxkU8p+4SbKOplEV2vj7rkN9P03KKm82P7yt29MxfrCjw6Oa346IkjXX/JmpvJuDfw
lLMbZ4xmH4RBe5XEfqMoo2sUPu3Qjtp7w1gp32ic9jL3V4pHDhhgZQm6SQuNm+5Qhrdm5diY+yoS
STdIPoVKs0Z5VQA9mPiii0NZBRsZ/wMAznXBVM0sI9WoY39hT+iYEJhJA7qcpufCdFIbIF8forAJ
Y08qiFUO+4wJ3VNozVB9g8K9GBGfaxRb3RzRBxklsX9e1XTdQV7LHosUiYV53H3lh7KNKKLAZ5i5
U+3DP5vSWNkpS/1XcvUglYcYHTzF1N+GTlo1sEiiM6dRB6yZF2RE+dagp3Qy9FJ5uIL6HAdxDtl6
pvls5Vlq4jatnBfpXPwX7Xdlp7wSXKy3wGRjBRILFttJ0T9iUegH6jyFaXf11Qc08jrIKZLNeZWe
wmYByxUIfEpikwepao2t+yyHkQc9+EcYIouYMgNZuQWP5qX2TUZDdppEy0F4z9oJOPYYF6KFTYMA
1C6LXZQV1HehkjFsu70+TlpWsTbazx6G4MWa+ECfbgaWIKUwNqrPIE51zHEGze/8lbCwWCCChY1n
WsmVsEsJQzr7xLl2+7nP9POrmJX6jp6SgjkyyPdSQGL8cU68gu//pB3goc8Jp3JAkcyGACRFE3X0
ZvcjEP2zIUOk44oPoCQvT9iVF/XcxNJ2XpwgnmD6zarCEViTZRm3PAOANtR+LH+5mGISvcX/TAkh
T6GxKKie2lAmJTwGFMCPlJmRWF+0/f+/Ua+CFBzfVnrTXI3rZ/C3NArcgev5N6F09NObcjmHhwlq
np2xki+kdgUph/fYRLfEh8PHjy8PWEsdgC3cBPYrG9SEisuGXvkzlO3bxI3HBxB7ohk/R7Hl75Ed
SkOOo34/h87SQdbx/RsMyXh52GJkCWbpwtEviDXWuPpjbiGT6pvW4VD6z4UFmGrVg1ihboKny1ir
6/Ddis0PspiUvT4T2dBPbVX5QO6Sr18cJhAOsDC9PkjALLgLeKv8WhkSV1/0d8ngXX1z8R1jRBHC
TLDW0Aygmeni1EsfO+jJSbBr2LgvNEZDIg22lF5IQsO3WeZN5vNmpa4bppPANCHnE4UTzOCJYzua
fddpS76PzFptfD6aX0Ii1O/ztaJ88SLVxTmjes0KLYiiD7vGvWUT1uN1xduk/arD2vjFs+6adrB6
VI16z92BWJ22NKs4tdmj1PNgkQxwOLhoq6KA2NDAkSy+Pf80J3WVvcPBw/Q4pvmv6fr3xJyihNtJ
q8cIPD1aOhljN9xYhBc/4GSQ14dB9XGNAARrgCdTgUG/IGjQcK2tcphf0sBQxb7E3CZGzjzZvWMx
hAMeOEj4e9Kzkl4Uic1jS/ObKulVZw3Jn1YMQyX1oUodKiB+qUKrTPjcjF/0NzNu5+8IgbgUrogf
284yOfaRVLDcyPOiqajhLSWigsJ06+Nnzb4ded+b5Yn+7pwqPykxGSBhuqIrJ/lYtuOeUSi1PPMT
JH8g48WuVe9AHfJ8PnPMVWPgGnoLJdH/ef7gjo33J3/PsU63MYL+KJDVVYtAQqpEBR3hklN7kPBL
iwzMSHc7L1YqIt3PpmwY5K94lvc81n3khGRZVM7rM3oL8y/J902tpMRmJmBFwNk8jIBLaUohLjRN
iQ6q8SkM3Trp4lxADy6kUbZ7763eQXxmX0aMr26sSnz21J5xTusxBu6MIdjNcrDssIgiHFSYuJ/6
8lK00ggvNsfwns6BZd0hM1109G6bYGzMf7oeVDk2HTIUm1cYZA9zMjdh+dPgn2Ab32nnvk/qKXvT
os0ysvxIuWQ2k9afre6E1VWbPK3P1fPzx2FEQrq8hem7oMZxAyjapNTGpYwUva3m7+MEw1SXK3Fg
bbh1HsudyzJ0wU7afpVljpYvDwKQF4HhR1VBrZ1gFcN09NchsV7aaqY91EOWSURY0e7bcKI6G9g7
8FfNd6g/CTv6wgbxvmauywQkKWUXq7iSl3E5Si3bTvQ+/bWIFqPqFmGTS8RQTm1Zv9KSIxMiG0xi
DPqBZTMWTj/QYwY/BnQU29G5WnQgLql4ewcji/cu+YvDOMSE6wNOel9ecfw2YzLREg8jM/PJYjso
z80Dfz2THVO96lX2vX4d9lKQJWwYdqqwc8ZuaQ/2n33Qyf5D0Fmwu18mU1Fe4fMb7AvftLDfX5Fz
/M6n3FyJXhm2IXYHqraIJkm+o7VVlHPs1HTUfs+KxbDkRFNyAI4eIyb7hXVfm729DAgjwZmG/77x
j98K1xHffZH02m7Hj+8jdbwhgC8fxrEpGBva//PG0efhTAJxDY32tXq7k21UhguEx38x+KihnclJ
q3G6kslyXjRsrySqdXp/FiyfMmJcBVcA8vuoLPLRMjvbOASElcGzsycnl0GJz1ITe4vp6fppaZtW
YuuaqyTGfplo+bZf39Sw+sMHiyAKBDOkYpT+KNjFIizQZq/a9M3kYBiqdMU9ezkrAYAIB5R3v15T
3bd7kjwFv9XwpW+vT09CxGXN7RXUSBli4nCBy8u5q2UmYNDXWyobOEPDMbRTDfm3dnEO0JMF8lO+
Wqran4xpil1SXjjOOTGRF/3+1GyS9a2MVMaZ/IgNN4FYrH3BRS/XbL1DDrGcxN0l5P4lfKx8cr13
j0lAnjXWLSan1zLtplJiPblDjdRyOnxs03HQWSqmy1xZE0OIUcbr1yAddXgs3Lv2jPvZ6ZIkqlLA
UaX4gLiiTfjkAh0tfPtJtCn3dPj6NLp4/Q15wA1m76SsEbMXg58SeLncUKFqtxAtIXNdh6eADTpW
k+e9JxXxgpVnNnHlbIHJDfugaGNgqzkpTBCefmVRBvCgiw8kU07XCqgW7O2RJ37mvnHhHhwBhKVm
gy0+pzvPswgrfDAq4WBHddD19cX3pGINwLyuXXTZyxXKsDmZ7Ag92h4L4K3Bqbjx7XLdzCXhKkpl
1O4k4ScJqeVjrAhcuqWlCcSEth2Hzz267KV7QSwEKU+ZsMiAQVUAz//ZvRGZmp6FMm8vvFSD3Ze0
/cL4kweh7vgKcxVSd8D2FUCcBY+c+fDlDtulO3G9mnxjN3qWQP+rvwy2Rp1KaIguUShftVcfy0OV
xMYuwHsLzr4W1mF1TLrXE+4J4C2qZLtG9G97KPJX2SAvOghDu2uImELJ/qK4GYWzvEdlZBpcfc86
XplxC6SSKKPn2AIXKODSi1TYtPIFK5QykCIU6oCf7aX6J7ArjPRmQeIb16rC96/kZrkia6D29HS9
4r/d3WGutcIUxAGT3FuHaVQ7nPAuiDAivXDMS9ZWJuYskLnJqDlGOaqw0Jgy8Y0idA9zlYEh2ujf
cnxJK1uRSrudMYYUbzhaZl76+l7dR2jPxajEoqHP9BU6+MmAbU5OyL73Omrx2PZ1VNLPNBXKpH+o
JsDEDpg1Kl+eb2cto8pm0xKcHdJGSnJmTvx01V1ytMLNNooWyXfO7o3s5cXzm0FWqK0PSUNH+Jo+
xMXUZg7u1VeWtI5iMXDSWGlIYQZeJHPuEzsQ452I4INfl3TClVdv4ya7k1U4Z/ku17A6tG0ZtfYh
MySOP2iJLxQKojKJ8+c9Xt5DQ2U9vsV0NPAuWfU8m9I9SQ2+ShdqC09QaAWKm0UkV1V//4k1KSv4
2+QCP+EFabYAtFiKWyLpLyylwwgWAZ7g03cMfnLmXjaiz+6WtgJjVSnxDOheo/gV7QzCz1zRcz+a
OWS7SG0IhBcabvWD2wNowXV8G9m0VR4lG+Ojyht8EwqD3jdKBKhLMGKtuBGK9Cfnvfjj3+20of9I
M79+A3v6yW3r7Y2V1/vvKWMYuLGbHKxAPnNhziOJDMCxPCIrbvxPRCD157HGgIn4ndJTNSACo/nh
3sj1HgAzqe+/h8eQY5N3XAXp96VBnVhMfFTExzj7oNls9cW4WE33DTjKtuM7rThtzbOghDez9TDT
JUvh7UdVo3rJ+6mzE434QcRsnWxgHOnLdyHbc4gErlU9QPc3jo7cdktqaVzOQcWbfsWfn2cI6RA3
rMFHSlSQmdO4GflGl2XC5Exy6MQ3QPC6U/U1jsXEkgTHdtYYLP3n5yPO3CJhtmERhjuyfyVWOyrN
UGJs+UOe8RSkTlYz6sTWu4Qx8quiuX3jqFHa3IYxbgSeIgC5dOcDj1qu3eoyYUho+1jzxMgs0JL9
2R9b5OSOe1AL9h5ZeF9yRr597S20DEUZVGYHutUVOoiBHsNrsZwcyd21eCcV+wNBk5YkdNnGcekt
tQG2YhFKuCrqHVfl9wtfO49VDGA1AS3d6G9E4Dm52lxdxU1I+fuaWuHa3g7Qjay+6RDdaQrALoaX
Du5L1fkA3j5cmbdTWsJ8mNlYfx0fF9wVZYzAZhD56ZAWI6CEcClWSU1l/F+HxmY9e0ludi+5Eanw
RQ6iv2s66SIVqY6wk7kbl3zFGSdsSqIahbP2p/YdCGlpK7G1zpNzZM+sBw+HSC0tbRdWG+rwFf3K
X262MXxuMjxxFocfDBxYSTCFm1IdbM4IVszC4DXH695qoXHDt18OJBwdGaLStKHAIsRMc8qoqVTI
/XiYqJZDVtOm0zKmH/mgLB5JMq2mSgJWCtPu8o6ahullL/DqcsIUGsbv5ujtOhAV9vss/N2jIeCa
RuHInhsjLWZVYskm6fox5nsDG3U1itXWJ/l+LCsT75bJQPnMb/dl5XfdxNNXRuNJ5okvrDNf7WdL
d64FvK5kEaTgeDVsBe2WNekwf9zzoDWsu2bvVTLQpLbwwJxKZsPVO6u3iNEvLOvUrGGTJbuALzHd
87UPl3ghxN4agZQ/bizV7bxkeXICOpwKR6r5tubV+/bNsibUm+0o8TbPdRgT7KBnkU9SAW4X21An
XPBZXENrxTCWrOXKRXZ4X/kAQttISdDkVT4jBDWXr5xMV8bIa82vpFJuuDPvnOMtBdyNFw0CyT7i
b/Rt1GboliPOj8aLHwTHRQcAQ/bMIWWTh8DvzdnjtpCxOwW1454pfB36yXlEqpLiBoNRCJ7vXAVU
FN7KnkzvCrsscXAq0YH10lNWuj4t8HJiY/3Cy8TPdk5rFOQ0R3+ElT6MbHnWqRsGHvuXGP8WhSj/
ZgPbgQBThIKXqvimE16ApN05jYjMPiw/h4751W36jb+e5rUoVHQSUb87oW4nqGJyvqhGw4j4m/0V
TuTY05lZllz79xO5TMMEt35UCjugobXycIxeOIPjxoOp47IZ/3pRXOQ8WarJmAIIzT8W0NfuMumo
XL2F7Kd8rgBo8fJnXanFObAW6jtJ88NSInSgxmQvX9soWLkutW+Cmv8/d5cYPBpCq/E155Bgg5DN
HOZg9xC8Bft7YvzrvmFUVAucpW7iZmZvtHs6FShSylEjKnPQpDXEVFdScRsDq845jU8/tPDjS65n
/T6OQtYbIdIDqZ2rdIoin69b+hxWPD6KXPgPzgx3/98ES2dzKzn8901beBDzwh2lBz+YzGPpQ3GO
jxeQOkZCIWSY+VheXiO2QHdl8ZZAeEyxE+dDeTyUBIoPuUEp+pYR3Y0ZyEZYh83A1SrBBpuYw2BU
+T/1s9Gk3dcQw7b+z4cokaqiMS1PVe1iIDnlJEGvjC6m9Y7DA8X/OAgkSpITtYpahZpeRBi62Xx+
im2Om/CMHP8An10Kn0o5vUjW+Eq0eKRf7prl6UHvUMlR66mPwWyBsA7zfweBw1AfHP5pZTO+JK/J
GqnyNHpP2e1pt5/rFczeOBuwoDc9uQAFJQzs3pbVH9IWrC2YSaTM+DYfV4Lpv/Db4EdwezFOj3/A
SPHrnSS+321Y4/xQtfGtq3uPMSdBu44k8Dy9jyhshgMv7eL+kXGvS7sZOXKuJ82BQP1fG9ywPWOH
Yvhgs0tSj/PwUal8g8bcWEZoKp5WyRxKc9QyMWJ/0WVnvyckbzMHbyFRI8Q1PjHZhYkUyK1Nk1mT
1kS17U5fklyvSyxxAx2qehXrj9nz1JvyA5XOgI92s5OBp977VW2Pdz8h+2mmw5Pw9k+elAwgI2oK
p+CeufnjiK/L8Qf3uCtu6PKejndc8s/CmRgVJMpxHcbmL0oiWFWt84wrdzq0j3siHgc7SUvnAjho
x10oVJW1iy85xv5eVHLVZ/mFzQEnKeaXmwLGjcd5B1ZvjuUc9pYMivFqFvj9jB0wPdKkIyMrO3kT
SQhtISbiFG0tyOD3STHVjjtSP6Zn7IH5H+p4NeToNfTSA45HWCKvfXweZeR1CmMUylWmNlfpvZut
lEuQGtWk3rhcZ+tOqEL0+3JPghL+oqS1MDWwaDPn80uvUP2bt1a5jLqpKpH/tElEOArPdaCIJsvu
mmkdcelGUiDEfOoMvEKRadUzfIeZHZboNw3XrLkKWx9Z9lmr4u0HQbzJwKF4Uzr89+ktNXuGFig+
lpxf2PwOUNwEDzgn5/UAG1axnsMjIQqUNiC/7p1sLeZr1KIUgq7PWGWmlWJ4mMmvqjdZPblVnKPy
JlP8EAxrw6eAEvyPmlg1dtAqUejAjyWz/QlM9QwNrVhZxtuabNwB401krZE8hTqMOtnfV2W1XBkE
C30DH6Br+Bld3cxr4QEzJ6KUGrS6qmFFTgqlClpP/H0HC7+22QaPzB8+TY7UG7d0qYlRP3ROFz7x
n/gQAp+lfhXtLQ+YwqUGc9PsYXkvSgaHCmWKt0dJtw37JyOZFji+VQNSQBlyF660mSsqHk+nNhwB
t3rkwgSUnySKYg2CqV7rFJ0i1ybu4/TGEYFKc56SRTet8skwgWn6ixs7Skr93dgmXqJTUKYUBt4Z
AZrRhrexQSlwshV1C1AgCCaQ5/0cFWZ3WB8sTQ9qbDNVYMvjYa3WRkXoGfmNtsOSvH6IXik0l3DR
mNLaxB3fuCIoG7M7WGzHHgrxCaT955FclC6lPoeW2BOXBY3ZF0Ntrc1P+VCR73NefrNbazyEX+vz
lnTJZ6iN+TvyhOo2lsm2PB9yzeWYLsyhymAdOYqGFgF08kRfIYO/cCzSSI9ZZYjeXAkKtznVBpu8
I6ME9uyvi7BZIHM1dRQXgP/ot1OW24TRB3fCQITLSyt/mvkHoxynvyqGy2c5TlEsFmUbZA1qyVhD
0wtbhkT8ZaV5mdivtE30V+1jh3vS/BSE+sDMLke6CKP0TeNIA2RE1pPIrHX4/sCFSlAg2D8XSUuz
ddSifBEwVZSVgm8YKQYM4LisTPwpxiclUfQeCnXugqh3zDJjhhabBx4pXQSLZhNjNO7eWlxyDNHD
a8s1WYdXpxKBnLcc2LLJ2WLgHi6b1IvBRyQCNE8pOFtaLEI8bspvZeP9CF3cS1LX/Buu47H8BWCP
0GTx33DoNtT04HOw9mg1rqLZJ9BI2wCMEEclagMVyt85AMyCXj/b8KjpTde0XPGtP7czBNtaRNyj
28QKMZg+EsUwca5In4NzovjwdDxO/PIhtEKbnTWF7AgOnvwYyE3itfLbQ1pOVi6fGVTin+JKjHwd
kyM7qD6dCBbvikVXgeM7HGhZ7Cayp77xw0Ha6Vaa5haAxBbYJOVLMGp7PPgY9MKKeL7vB0gEkFgD
GvlLEUItJAiFEeUnZc4RAtjglMlz6PvIB2AmVjcGpWu+7V8A6ih0sDxDGfiHdKNsBuzOYtMVQbzL
seDQZY0kddCjPjq1HgLchtr5I+DpPcHcTOOrgJ6hRU50a20eC1nN4dzbTAEV1SvDcRPViK8tkOm5
hwKLBY+yVhI6++w6UegihrE/EMisZ2RQPZaSFEu4Wys3GgL7Wjbuwy+y2PT1bPqAtvpkNxS4hWlX
PwTQXxQsarAXxVuLUHHnDp6C/UZfzyeZaM7R7l1jOdDMK9cGShMh529Aoe4VkpynFxe5U3hQJpaZ
PObCo2yH3MW1EhgVfeR7KUvxgLrbR8awroe2iexQ125xsZDQgUVmhaTalo5Z2l00n1ImQICiV4Dj
s2NrXzBN9Kj0cHs+3xK+pzOTGxcwJ4ftCHRs8cEHwSq3Xy2q5edx6sn0Z92c4g0+G5d3zwzHMqs1
5BLHdq/IZeOLUX+EJaXqTm5E5ivFRjwMHjUChvI4WX7/RufVm8IB3bLXJxw3Np0ZyOJeGIorWDas
e5hDOyb5Bos8ljrZkp28vHfIroLmQnx5SnAj3CES6/rFZGZU+8ACIVtEkm7ZCfbL9r6hkam4Jg3i
qD+zxv7avzQrrw2xzZASoueGzhURBM7stkMrx3zmRPdc0zTQYeF0680WPJCt7rTb7Ciqs7HFBqUh
+prEdF2/ytJbtmy+4PDAzNfoUKRvxlzjA+3WbwyPA6z9ntKddU5Dcav4EbcXSRp63PiS3WGzhtKL
/+rEjbS2JHB8oV3BhucdFrIm1OEQb3cQ/eedX3lF83Wv7sjP0Ub4Sbal9OGUk6n2HAPPQZwxkLL2
gcc1+OxpaJjUldDcLrkoQwmFejy242GCRtOQz3Nwuu8ikIJmskWKjlsw/HkNF+krKnA7zJ/4pDel
RYHAePOAmofDZY2lQbIA3t6bRwI+ZLEJopI2FR0NNCrAMxHlqFihc60nHYCf3igdFiNOISb2CcDg
hjP4Uh1UCr+TE2aGPJmPxrdxhtSyTBSpJlMUkY1QNkaYvQFdac1ryBQDgy7UHJXnUJcUnuYtSRQP
PUTNzUSnUXwi75WHtwCvuBdoFY++QKJ0zqbA2bvkp8POhn4LGo+0GWId8KrPGVFfu6nl5hbRj+e/
jc5sT2c8SIRsAUV1F2Zpq8EuOSCeOWG3keidYVYdR0VPYPteCVrMLgILOgp5jvuRYa2bjcDFxIOf
EKEkXKQiQ033o5Ogeys+iTBzKxDJ+eyGeNTj5MKYsFDzusgE082RifuO3k4brW+C6cV2PCDtTxfR
tVN83C66ztrf7ssaCfa18JkYJgdxAmvSvIKDROtRsf4ZbL+KGNmXynnOvTElR4X7+AJ9Lwk6hS+C
rXAlmkzG/VfsCyRjTiljwXS8g/0roy/AoQcH+vzyNjDcvAMGYjWsAc7sCUamD0tcIZYRNYVzO0+9
/3gVKiuY/18tdvO1qe2c9KyBWbUwscXqw8yZTSOgV2M9xTFq5X+x5Pj8PBWaN+TEMcEeN5Hy6Cca
SqcTLA1U9TIpV+IBGWJ4+g3d5CIn6cpBhDJyX0biIlQ8LJlAXwTV6Qa8UqkYiXQcvE5uRjclhO/i
5V1JZW/hVpGUYnvVYiGx/oOL91I4QCxBrzy7ehr05ydyURsKCMG7Pa4FFaHo2DO+C0VADyoZM1wu
rvJIAELR67WedrMOeCiDd3fspgMFZ3TS3e2KDde4xpdEreo9rVc0K/SlGJ50Whg1naCFyPn5v824
2OvTmIBGSFgEB1QQIce2YilS4jeUzG9H5/mTClziYQXunSOD3f6sxP/1ImToAu8gLid/+3lrBft/
I+SLOwYHK/QUaNlC89wFMX8s9pAas7HdCX/Vq5r+A0BAL6VqQHkcKT/yo5odN55wp3a4x7k/dhSO
fmFlB6PSzRrBVIr7QfkHSOa6tLxyitOaeMMOPPuc0fb4NVZJpZOK1A8WBwW03JKfaokALR4tkOrJ
sFhXZI73RpI1g3rP7Ukhyxn+1w3yGo/j7Qo+HKfSVNFMZigM9RXVMR/Gg5bzTy98hKI7kxCexm/d
f7BLlKjc/bi6xP/lXzh5hcVRWA976TVq3Nq4JIG8eZwYPBpJgUoNnYR+yCwaVBLem5R/6xHb8ULR
o0XrqYkaqr5aOubRrsJ1KA4xmV0XO/74n5Aak0oEK3HgihK4/mdqfvq6fqqauREuF+urTRIGVqfb
kWFHNx32tMWT7IizjGG4zmj1SamJg3WoD8IP377mhXlG2OD7MHArHycCsAgvCo5R792ZA0TV5zZT
BfSCSF4R+FKCFahQfQ1CVu0fXmuOP4n3xqhdiboO29bHyoVrz0Relfo/RuM2fvdcL3BdqCmT/WQu
rFXb6c/EkFlwtkuQCIycU/upzrlAoHPegNpLZqpnOomo9fbuWJfWXUR6zRDk+MhZ/9g+hyIHdLPK
NWQLgwWFcDMQNGf7oUdYhzucZRdjuEE6jcoS3bjW1P+IY+6E5E0N1rzVIyDAzDu7J3My4W6LKiv8
g4dRXXptPrgZROL2IzGNDAbkdmmoYeipaFlnk2u0hbT8Fy6ag3Vn0Ezzzlo45bCyUUhvPg3AuBS/
pVjCefd6rh3MQD4o202tB+7inXL2/71CHA6ozpOj3bPdTkWKTDnKYkw2qxVsOMzqNt4VwXzvtkUI
YxX1ctgLhNDhIhLWjxb4HvobBFMiLKE36TTFod9qWI/sPLRzuRI6v0AsPOglGdcN7knOSr0hdkUR
u1XLxtRMNuAQAGZRIsTPHwpDZ2A54b1vxNe+6y6Y8O9uCPrFRhzXGnE1xY3RzIBjWNBRmPgzhNIH
Tm4tRjy2om/BdmdOkYDoSt3GhvcSk/w/O1PMd/PonB1H15gmlAclDpE6d5HW4TBm7SbKg5Gtqv4I
6Ag1q8ex664SXfqb8GSexIY6EkNiT/GVRVaRdIp3p91C385L2s9Unl/ka1Dre6aluVx21bL4yyAO
up8NVTIec2d8N9YYW4HjJllhYcqRwRrgUi3omKpaZGQXRoJP9xiPIwo9E/9fGhHt0QHvt7TLnWci
1i6POfFNJx6JM8yNXdzJAzW0W1n2lbVwJkvdUTgGZXWJmBOz2WaLPRo6TpEIIarD64DjNuYFgCRx
LjsXkpdSbfO71NhdHTUcr7VWQ+YAzcQrJIMCrqlm443rtv3wWLcmAOrIqOv0CTsL6SSDlH70dacy
K3xAdnohDsfDcNSPORevPxT6LMVDwCNVTBbgFB4H7Lem4HyaakT/PX1GM1glIZY8g05mPNkWVfyB
1hZet6OgpFPf01rdcqvui4xi89yogw1wkIzpfgLUfZosmQfwus18Jz0Zsv0vPMyc4ZD9mcmDg67K
qA2fWcgyqqPllV4EmQlW4uGCsAJ9KxDBD4b792RuML9C5OtqGrn6L3rFUadT5iAqHDsZXD12gaNh
DEmP536ZdWC0DgItQTZnvGYvv+6vcK0wN5vGQMAjzEgmFjkkVVnwS1JF9fTkVgrCyhUBy7BFWDw3
eNCFmuJyArbVbzLana+T7sFKbmXzI0CFA20vO32w6PWuK8F9chol5MFQWuZUqjVydri95dnUyYq1
++JQydwWyL3Zo1ZHC0pAgVHwDeNfp8osT/yWxQ8s3eISkNWNLzcN7eSM36gyKdkAPoRXxhwJWZGI
iD3EvjBFnSOg4Exqkb62xHfBgaCHfzmlx+41moXM4nEtOOZsRGFQ5o41JVJoogZmBGQa6JFCC6g9
WOyKvgeYaARwkYTvae39RUUNg7Xqj0TvXOhHu8cVw4ASd0hDcfjtZtrhClFLVyeXNIakPVCE7Jny
WQCx6ubBsg/OaDmeJgFVP2/nJ4t9URTqZS0Vp6h7nqfuQh3wItxkS+pncDhMBZ06ZN/zrtwPGD4Z
vwOemADgXDl7P73qYgyXWd0DJVnUqAF0A38B7Acp9AlXqYnC4WDiBymwJKETokPvhpMbUlFp2h1w
DldmmZDZRkMrYlfClDwidLM9R9so84p1vUXqXjM2M1FG/md/5IhqE+5rSfDN5aX7TONaVI06msog
ucBhrdjO/r0+8QYxGhm2I8/gMitol/Hfle4nAuVeZj+mZ0miNemAlR+qgkCf2K66Ph8PhMgmi+AA
6cRFVcyWqJLMp3buSr5c02Z/nAJTlyi7ykwb4/M517XrsJgTdux3aP+kx9AujnCukmIIWFsqVvMK
43VuSsqGfK8JZIZorzqS0jkGVKJGXfQcU+zOjHatJVZlHQPOeP9PETTaI1+9VfmslI5vdVZx0l4/
3mWhT9Or6bywuUs3sV88r839jkX7QpYGNBF8unFJBlh+97DNjbwA+og+jfRt0kxY5kBbkbO0ecVh
Pp34Ed408lmzFpiyS+DQtqSCZ4BlGGlu753dBsdb2tcLy1VL32IBXb14/E8UGgANI4Sgv5dl+bmH
CP+4xtqFuZn9/OGLFg9fiovAeGkxtw+SKoktdg9AqEnujfBxiugNm8aQAEa8k442iwFoaawOxis+
lUlfidtqGGFT6VfNIMbpuUhL+L9UTwkVrKHjQb+5GONOl99tJStpZARc3BVLhRL8uug6JBJ+1Wa/
DuZQbzBli8Z9fNMSjm5ig//UQW2+UDcujVAMNtxAuQn1QcJ3ZFn/xmPJ7V8eIQL/q6gZWqGeNFDb
tRxASyoS1T+dHzTldxwZAax3u62iMvubHCLJwCW0BCqz7jgJWooYaNj/Q0aNtk/ZMXlKVB6Lq5TO
iDg7QQeSIU9BGwTUZ5Vk/grGDiS1Fz0N4DVgUX+V7oNDUiCBfSAWzg/v98UoO4b4owpvVb4v9wBg
lEuId6I6whg6rqrYyCCYUMzLccDdcmcJ/ySd6FJZHhQVEjxgBUaHrV4RNGTgYf+iFQZbdfMVHr1c
khxUy6nY/Fj2a2QVroCCC3BxJUmxZfxHfW5d2uTfvDqGEhlHM+PXGpKlX6wkv0IcsF+9Om0Asg1T
UfkSRrz0cxApCeQ7kfSyAqml54ADwATzKqQUoYrSNG6qayTg1fLWQv4b57gj2oRJLnd18oa6m5k7
Fno/nh06SNAl57+M5tOzE3hrw/DjqrdeQ2Mmim2LTTfL5ZxYXSwhxAkmWjBbhtN6yVMtv46JDrzZ
ZEYlZ/RZH2LWGl/0mIUUYxrSk7uadWlR90/+88KHp3dcCREiKS5ZBBsLR6AM3E066K1LPT4kQCwJ
0ot9YRusOi2aCHAYkhqqwLM0dIHTOEQ+9c4Yr9x0whjI+mar3fM3ZwFUtX0mSzAA/ztbdSo3jRwA
Zg6B6Y/XSqjLyKZPX1gN0WIM6wH+2Pgb2N93f5TfybItgDRD7QsKZFTdpvWQrIzTCIVQ/lyUt7Z9
PZa/BoLCWEAb659EA6+H1IBoe1tKD920u3KsisChEVjV8qfP2OvvjIKYT8FDRXtDK77DMghSciCY
FwpymbFvAfE23G7C/OP6u03Fh90PFUzErqWDbdx6J7qSBiD2ZxNA93+aBOGdAU1y9H/NZrRttkfu
jFjr1uUX8SNLX5SDDfzHtJ4fIcF/l3ZY8sBKSsytaDEio9jJQA3vS9/a8p47VB7Bhir+crS4IO6f
0sMJo709cpdJ6b1RfkDo9ATyNVjGCw/EpouEV0YblmuxmETcpkkkx0XhQY2/DGdkEQLCgIVhGD74
QNSH+NgiN15RBJjcVVqd6+gbRkqmbtgjLqxgNs9wYsZRqmwyVVUiSEWRPTTyVEsn20aSRxkksHSj
Y5h5G60oMdA5NmwpdQ9mZfBz7LWJ+jRboA+WUtDBCmbL8v+1SMkwKRSEj+hK9HLRM6m5IL89aJVA
WNyyC6V4SR9p9XFFXKk9P7yprkgQLUGJTEVZRHWuGI0owM3EUZVP6BZe91szewbbsN7U4IrSUuPM
Zx5VphMS+d6ZCxRJOz4VvLk/ltusqcgEMXJN9h+NVaCnZkfCZkiQh9BobDTHc1kqxuFePOAQx0rl
+iYzlUsSd1S+ehJ9CeVcIWUDucq48J15f2E2YThUVpLLVuvnELBBSGWd9qGaZTF7uspjybNmSKiM
kJu0fGXMWl+czs0nYmLfx0SuVPaSl07Qdy/p51EPdknW0BqBfcOLUMwl+V+hF0w3pan1rvv8m+ca
tbrpkW11062KyHnDtptClZSNPSE+o31RH1UJsWCF4SlypwILNGjYMvoDsyvprdz/C+kpuEtC7yPr
yYme4WR0GvtqpsPAXbp/IMgOfy7hLfaQH4T3vO6zqTsEqwLqfkJJo6F7sXW0LjN36BBot3/99mqf
mVUAcZcKy2yUh+S3tcjX3GScjcBnUJWT31RyLR8Tc7CUjbrXcXst4806XYFlGEbduKLVt1bE9jDn
bu9GSE7MdCP3nvc8xS/xwHheJ2T8dg6AxTah6Ag6ssNT/QOUgAPERH5jW4zHg1fXwlo4dvoMaUGJ
HT6JCtcSrYTGMB1gcPfjtBpM/a5S2gUITNVswNM28fxDyWXEFi13oKD/aUtprvBHfopk/L/1DJBj
YxT1RwuzBJ3ofdi4vgYlWGHaH8mu8ls27PPhCQfYAcJCr161OPfARlMx6eH9kjkjC3z3VPWbpYJ9
CTB3Sm3gZDX4UCq3qArXALl8J0C+r1pAkkWG92qv8FWXkRq5AD7fVE1kTvmOq72i4n12zgpkGdU5
kSTsmYDuT2O1Ghak+ttJNZCd8KeMf1gWL0m8Mo9fh0sapF1OsRm1Mv45c6Iv3yTfGUGcJW/6btTO
bIPVN3DcwFFESO1BC0G2Rvw7PSM3FmGbEA4SMKKLR/28+AM99y/HtWm3Hpf9iOM6kjc//p6Rr536
yi+Ak/yYGmOm7yYjGfX8pEs5uHiz5HCqFgwIJfaaXKsn2Ne3dc/WjBmxJPIMZst8nLarZ2huYOZG
j6up2e8/1TQyHkdjGeWJXbwBODHMdNCEjDy72ogHiTJ6KS+7O7elSALlW+gVSVwrjgCrdzSaErQW
YdhHTzk0ZjxLrG1PrH8fGr1H8dWmXJBoJ8vTSlA+VxSGg0sKqGL1oA8/aKoGNa6dF/Qjwt9Jwf42
9MUrbqTrgJljqEXCAz55YLpRSaaZVRNSyqApBU1jxSK22N65tOldDaQQQkoNuHQq2S99rmlCGeur
pJimI6Kc0czVjBnvPqqJYHekv6WU2jji7IXM/T/VBUOGdElSn6ZVoYksMLugkj6NpvgHPLitGned
12Oc/VgaBE5lP7fD2wDFZbsxugc6gApRXjl7gp4S64vONuF1+arg7V0fuNZt3rw94wB5L1VuCb9U
8EG53COv/PTe2PAkEo6+YkUfI+rLmzglUpM4sv6iMFkJ9tqS3bR+gRF6HWIP3hBzEsahDD9UwCBV
VFeFjRuXsxiG+QiOpO64n7/pNEFnX7RpEHlDN9temeHRqpXTBMYyJoq/D/VpUWXPGWsGD6N0COu9
CDfBcBYfjhI/RP/fokgNcQhqBryVrn8bwKVLquD+DKGrA277uPvKILOru9JHf8o8UIj9LBH+HF47
Qe/fsM9dzJIMF9CBRb39e6w3247OktHuZV0+Afm1OnZIOLlPB9Icf3IYk0IfLWAotGq6DWKYz9/Z
zdWIHSuWmh95RUdZY/67s0QtwmTkUvtmmvL0MSzqJBzp4v2jyQPpQZ2IEJAY95djWdf3aKQcfQPp
zSyHhVZB+WJqQG0HF3MhQplfsCBFb5Xg4g04fwoxKdJ7c6Us7w69xNF4lvO0vGPpkUTDAoZ0eE+U
WLeRp5PkiscIniPzqiwZdbwBpkf9hGv6MdifvKMdc5nWlTSXmnKrvj59j2nVoyPCrHhpduZwhur/
G47KGv0/5dtRQyTdK7JX+wk+xBtXnZ4/g5+oIfMAuxn3YzhPNXxyb40jMYSAIEfAj4sHxBcm+guF
IYx30WGmEdJ5pLo3qSTy5O3IiZLlU1cBFXaR1353oxBy/2htJI485s/aFMLalHd96kvMmGJUjy4S
ZEpoYoD4ipYd5Wo1YWdS29UrYbEVKHF6ReAg/TOuFzmwPh9Xaz8b2NJ89OiShMwKFHuku4YNYGbz
vnFi1NmwxNtskYvaNiqugm/tG0qhSMkO/xpYtazA/paTktM9/E2ALMovafQ9aPqlt/PABMwzs1nx
8ISP1pmnIPmJZpjQTv+5w03QtTEaymkuvOOqq4mJCh5NlX29Dsh0lzOEQ02/rtNXGMGN4x3wR3fV
RK5tKKmzeso6z8/zzoN65xXTp4FGrRRT7RrZhG8uJr4bShTPcEXnIRZovZKKaCKYXU6urd6T31Cz
k3WnGjYewBXYJTcb3TieY2+LtQucoW07GLykSvTlVJUlasnfeymRDqnCIpZvY5OSEX58e7TZbDMJ
bzN6CnI8QSK3OSTduqQoaYL1boCLvcNUEEbqa1UeT4Wx9BNoBE4PNbl6VWwn4CPcCVF1uQ56LF33
v8B3oGPwnmBsyMFRsw/HvoltINcaeXHQLl3nj/aS18KZ4PnqiPpfHXl/ye+t7rzq6xKWvleCAzIn
SYdJIuj3I4l/SVtUDufN96bJShwffvxyDTy42CmgpryAGduCj2IogYPaqk4pw4nSxNwCSHPB8xTs
/ta1dUwp/xYXAigcCYw9sTY89xLgxIReghLuDwojdyssniJgV2cQ5H1OECV/v4eZFqEnj/6Vq9H/
1MkCm4zhlopnhD1M4Pp3IhmXbQ9XLBWY32iYI7/Y70zF5wNCJ1bpvWdW0GvbaWIphzcQKSiYWxVI
OYxII036oUDWzTuv1c+EZ5/Eg74TMIFs+2NiAAszpOTEUEO8AbY3xhQ6naZI+5WHvn31TTPocBdu
5rFKgocrlOTaeRufRkiwHzpez8z0ksZyqHC4iAJuOa4N1bLU7Dud/vCD7SoYwDfWKUtmSNBkApPV
Y0nsNEZDUbCFpTYMfZx7f+dsO6E8Z8sHhWFwC8DeLnzKJti4ys1oM780Qujd7lMZXeknZMWB0BHj
G2L0pcQrVZ9+oRNfxni47+lRjOVQYbKhCt+SLdnthudi9fzYlxNF6oOWm6X7h+INMc88EcneXNXx
B+ujOFN6dKUydLBGQvwVZ3IAR7IZ3JeHjYQ8DQVp05zm5t2p8raSQDwjAWDNDuRobsMjR3HLHEdm
B1uMton7r3+NT7UBWSVzznDF7OpqrZUA67SMsDMPmRTOWvPCFBDNhvCFSBd1n/Ay0N9NxoWjs17M
Os/TNL6oxVseZAt2AEJluMSxMjCdzVA7LjHQ6BwNaFOAb5BtFtPdsPKB88y9tvaa1J1AavkLyDiE
sCpnP2bDua2QdDK4PHtSytWTcSctPVotOO6S/uWjcZyAjZfOF8pqmN2Rymq/4ILfhsM37xHeGnO3
2tlMJriwIT5HMZ/RBhk9GiBFo/EoVAH1CUm1/0BWnh2Gw1CI8ayJwaPO7D+qMr9+HRYwcUqjjbzM
Im4Iw/7IRH9IkcD0WHHMX4XgYwYCp06cOfhn1mc62YL3uxw1r8bt46Rh7RKm7ZoOhnyBsnT6wf5/
cX6riGh9JCE7DnwRwLNDqj5j6TcjtY8x+4GETP1r4T0ndHS5NM7eWj1wcsUvWUDAcDH4Qi1YD2lb
YGg+lleaOIy0YnLWX2QezTaoo5RpbBdJwYhOxzhuILVNBPYua+W4pGanjzGVGKdYdlO9LCtYLyK1
XA6Rudt2V1ojBEwpZiS/eqd/Lrldu4H34sV01FhvUcG35TNxjdgHalNsjer0FCnR4472/MlO2zb2
/kshtRs7s3o7GXCCcOqw4O8Jc+8zY4e6x9CSNFLOfnZIBXr95mDShDLJVnm+RyN1KZSidn37WbD1
AvFy/PYGAHkstazFBC1/hf6tjpcu/fuTmzsK02X0h/GU0FLbiXRp/8D+hGzznBRksNhANdaq7qfT
g3tyKd06U8zYDCyv62RQUg8olxLstSnNo0VT3KlF5bbfTCPGTGbTBIJ+RiuVsSYOyypTsogI1ivw
Y8EP8iIORNwWDTH7ZteXqsi07ekBZyWIa4YNo5BePfUDp6ZghPyOXMtzuNsyPJJ96rG+OfxwcYxP
9WW4WJ+uGGqDMJjPT3TV3LRZGqp3i1yxKFDhE375YSeb+b5dTuxLsFAVWgVAl2piIAGDZzhoRpuo
PLlICXAuYiV4/8xtYaqnuOQZ+Azx5DS3iNPhGlO9eJ2otvVZ58BfiQAqRnM4q45h6WtQvJl9YGa2
lSfW/4xpqJ6MiOb5gT7Wx1U+YE/6R7ahai1qLvaJxX0LWL7R8X6GNAc8o1VqhvJQsNnfO4svmaRS
ch9JmZ3RpL0oThhGnqxCDcqhyu8HE4aV7pI+6LtuYhY4j5uBxl6qfNmPFTXcG/GpQLfy0wddC0F3
aZQxZvQ/j/dKFADx/v/YMtm/vQYokEQoemC37vZW+xtI7rTjmS6YfUsnVlQG/akPVIiOsNe1jkX8
6bu+C8lEn9MNK2fT0qaNFsao8x20qsMX6Fl8PrmTJr/E5T0mqfAYhhC5Kf/+fHx6XCTWZAJQl9yT
V2jnhFUTmweTPWgv61FQ/xN3lxEgY6u8PFqXfVPywvBjOVYRAsNDY1UCC0+uHR53iQ+lMNC6ynii
/dkl/s6n2PbziaWSoqFDJ4XGTkZkya8U5oQzMBoxCJm2UgQabVBWoQ9UK7lRaqZiLcI84BNJ/kHY
nLGhRqoqp+gk6OODZ0cqGWKlpR7wYl3sLlcF+J/Gt/tYbvqQfynPDdEb9tZaW3YA8giuE8C5Vb+m
ZRTrgjYej88XYHMrCRQlB2AChqm/1PujUureyoE9fns7jVacHS2cgRlisxnfG74kV88RiNBegZXI
J7qibgTN6GF/F8aM3KxEaoDkTpmpKI+rDAPuDNSsLbjSZE+gqIqrVOcUhlZ6HAiue3hOmyQ3yeAJ
77y76wY1JfTH4zSdAZ9ONdwLkfqFO/TJMnXhOgge03tyB3qseg1cLIBN1TArNpgNQ5IsXuHsH2iB
fM9LZXZRUN/liSkMw6P2bfZxI0R0iMlQzaAJon1ZpskEQOwfK22y0Hu6IDS3C0MmnXwq7CJdntuX
oY2Ekt0dNfDi71x2ZsnQPm/nqG8Fkd0jMsWLVFpOFR7Gb5PhHBO6lx0U1hzSwCZ4tYaNFEMOPog9
jtK9eQw9hhMhoIP7XYoIDWwWNMwKLVzw+BRhs81CDOSeRIQs0bIzLxobPTFqB1LOxjxLfccLH+Vy
fMHRnPv/4aLNv1trzsduFNZSrFXz4soayR4gJVzs7ZekUHSyfd4KwnPT11f9eKVqsIR+Vk2BOKQT
VJ0zkwIwPmMLItoGp/KeutCxzP3q+vYJ3G0dus9X20UuFTyba70zNr66bTbMh/MeKnVSJG9e99pz
KuXDO3TsNKugqwdvCXRTJTDarb4v97xFmRRSHlS7T43o8GOiKCtPcK0uQnf1HOPY/vfgFk6Eq7/e
38DDojgqO35yn3V+6VD/XgzDp1APqcvHH1NtvdL66zyVcyGvKqiE16skEIcTCR7/6bptX9hjn/Rq
N3kcINhqTJ+q1WWOKe43187jzOK5RFP4QfwAygSHCkuWVx9ohEszIeP0N1+AXOdFoLAzXlCvReo4
XP5omwGx0+0gmCVPmbk6NlN/aTbqIrHGu4JQeVHCRqKZ9YtS2ZuUDd1FDnu6xBW8Kg/au1d0um44
0pyf464SoRn2l2ynazdNv6bntMRAfP2J0qhvlnxgV8nGAuhjmGi5OiSx8gJ6rM8KzENs0MYoPWf8
Xn+e5krDWQ0LFu6/JrbMT4g4R2feVNg3mQCvtJY+QNcv8igKLmjXyR4DE6/TNpRq9PXNm9c+Ivs0
AjmDj5A9VSKNENm/dtevlfROThn9NXRBnKIAH13zczsL44NMWvYXOmweYT9ifWTFqgNBygWwR/4h
yNqj+u5c2F0OuvIxsvC9Sqqrt5sNjxtJGx4ywRCdZXUPLhJGBQQlM+hFEDHQVo6uSZkVcj6tCxS1
YzJ1DtfOh3kdELKvnTKrCrhCciolO+MyjEyZDzWwtayOq7v++X54EB6K566Y3Tnd2CvWr7NQ+R8s
GJ+Z6ejniMQ9Q2o9yTwpuugJ1dnjTAuCAl7HpVAEkiPP1Ea38GbQ8fxDWFFyIRuxNtHRNE5JP4ap
9H+qvb92gYiKP/X+DY2aRouZxY2uPoIS4aeyr8Fai1UQqGjcfBcfYbjmgt1ayJHOghtIx3cOCeXj
5VLR1INvyVZmiLNuktGFdR4BEvYJ/WzDBbrgfoj34l3SqBnZd7xLtDF3KXumSQhXM47KgT/QQZ/2
erPbjBo4i3CoNPz1J3JOSSwmXWuIgVgdKQxEIRWvobw5b8VKwP1rLc6Sfd8CsvSLJ77IpTYU9XoN
xwWzWW5qa6pKq1Ur+FV4QCRqh3roN9BWBk+87r60rhi2cbj7OQaPHO1Y5j1rfQkat5QkqLG2FLNK
xKx2JkDeg6oEXTBMiUZx071nRmwEFnFwCcfZzjp4lD803Q+GN4wgQCCQ8QLr2C8UhcXvmgL3fDtg
5U79wfTcx9M0U+jZBrgJPPi4XwagfbVq12B7/BdnxXRK7PRI6ndk/Kw7DTeTrpTVkWaovtlYHWtI
n+C0HZBwabYYmdTMYEzxzNnJSt6y5C2/hD1jy4nrzA7GAnbQ34PEmxQLUt9j51Sx9m3un43QVnBw
mQpeFxsrd5ftQcbnKuoIA/g+DbakzLEctaFcx3CvqfenQFfGUTIcXkeqTtVXiqp+Mrn+VETjDG/N
RFIuh14Q2fv3XSOd5thTfjKkzh/O/8Py/JKQIaFaOYmMLKAwWIrLgiE8RIOdP4fTlkkBOxTOj1sh
Us4w9sW6I4x1XjeN3BEM3jEQoCgyxUUo1A1LFoQVygpkPKcv93cahw5r9TxV7bUnx1OONALp0K3e
qvgzsjaQT2bUozBL9IkO+AkkPx7gfKC5OloECoAgMKX0kYQwemok5T+IlfnZWMpPJwxSwLK6g8Db
maNeBW+hUQ3+f7jN2yA4fyoq53d+9WIICSbo0myoSPQPbYIEUey1hcdRY9Pfy4RIUHdqsPJupWis
7BZeLeJj+opCtLhUWcIEjs6K76ihIquaKofX0kaYHrzVq8or1lukNfShV2IhGiSGnFhMzIwyVYgy
fXy5iAkM6b/jefwT1jhd5JUwt94h4HWAWK3IuR4Ban89NHbGMx46gr6xKoGBSKXySfmClNTnAdqR
1z7ixSRdDazFroXmidyf76IVdgu+cJ3jPw9HprrsDNGk/KOrbbMDzhB2o3wqikqWmTkh7Q0LiTkr
8mTiaXYPmneIwcKVNJMSmkQWbB4lJc31duq4HLwO3oP1W7Vuh0kLn8J0/Yf+AoGn5oMI1OVYrdnX
hQjcsfQVIFzDphYQb2DxrFPNsPGC9g9QYB13y2SlpufrCJ6UvmSPtmVbqd+xw20D7QTkplf1/3Iy
2SzUjJO4GVCvnkpF3+KGlnWjqq+dEUa/WvfsdkENrUwgxmb1NUY0kvzAPL5B68Pb4H0I38sP7Bcy
pwAR8vZhAhv49JjODJurSor08n3wrRYvlipFd+Kwp6yJdHA+qvHzfLc17sSAVAju/G6LrtZfDNiQ
3w/Ku2PV/r9IeNy3PZCux8JFORQaQuPAhTjwPqDks2Sl4k/8YHIhv7voPNasTXpljRKjmLa6HcC0
ftyX7m5W0CRkssgPQnHjeq/Cg5U1BFZkB7e2s3zUSf7F8UQcJWlmEJI4lP2eO0qjZlvtxHBByDrk
aBRX+YVGM3A5CNW745AgSAi0WShljpW4Q1N7rZ695mhU5IeOTna2j2pR8QtNpj8ctZ2cq7RuTtz5
n3wYko/Fuo37grSv/y3qaSs38mcB+juKtEP+rhQzHwxJJO7jIaA06TEZjGw+jhOa3wthw2fmGu0p
sqr3hvvFJIZjwUDWmHrrVxgqC7CaONx2KO/v3G7+LexaIgpNBRb1DugzexflGP39Wun/SMwHgEz6
KlNDPoFOlSd5l76ncfmugGwmZCSaKtne34t7jeso1O97LMPv0VzsNzVN51EuX5ZFBauj2TcsWlKj
4tRyzA4Hz/dlECKy+8kueRgAENK4Xq7tR1i2M7nVDZ0N2bvlOt9/1v0s4GVS3dyDQgedTppvAerQ
NCcQcALSUiFNrVGy13vAdnE9OqHoPIJB4r9hCmimX0VZ0uC5JWqL7w5CGNwUf6UvdLFmivj1QV5M
yoFIU/38PRIC8r6fGJVLCWpZ7Dew3HXRkTYQpcotJY3ii+uWKM7hQYlWb8nw2IKIHV/0rgF/OPa3
ciuzHo962YS6zmurmj/Hc12APt3f+VVDGqEh7KW8Bebcp6gguNja/3sws0TaLQWpfsa2GuMrOVnq
kY68OC/t4lLDN0G5a8HUJLw0fQ2rjCej0vyC++yRQFP6MaGvX5bqxew+5miDlzlr5Fv3TsPRdIGe
+09Vqkn3LbYc+1b8uSoSRq4XoWZ+aupga3GhXe2zAs0cG4wq0sLunF1SB8OMLJXjos2rMl/sFQZb
0U8WSDGQJ5qbKqypy3qBfv3DtjD3O+pgU0NXJJgMEQ0kTgXaZvJatYwZFr/5WYDTO/awHmMG8mHX
7V1xSh8QS3DLySKhqYuE7Bfa4g9Eqp7BRPsLxoxE38E2FkfHyChq103+GFy08ZQpAOg/ROENNr3L
tHWLhd8KGMyVKH0mmjpPevIBxPuiLGHMw4Waf5efKze+OFijxLdCMNQraekOtvvZLEV9Asosl51m
7gtthhptJrbMxFR3pXXTr9JLANNSY7/nW4D7twM1XDEzcyUlM9bpQ7HWiWsd/r5PQCc339R1pMyP
iwsDrVO+fbO5j0iwJdc24tED2tZfXGHRKsg+Fmd0x+g5WqiyKlFbAQKxLn4yYvJiHdmgQH/nC9Uo
Jty/IabKBSFqS8XKyIHSUOxAaqZ/aJq5sOxI+rCeCR/2B9wPixBKKFC0grzG8X+2i7/VAXswLh+r
rQQAnY1JBzV5CIssq22APW8mKRXeEVlF+iIKD3kV9/tV6Z9k+BAvjh6KcJLRph3Bbrudb8dkGeIw
Sk6xnkyKkqlzkP+/RM3S/W3k2Si1Ne8PbQg3UXwHqx++7zCR8XrT+3CVhAuXUYiRJszyYTJxIrjS
Rm4xvagJHRg328Kgx0NlvF84NfgidAoesdGETQOh1sYYyEn8LnEMamWMJgdcvLP55W5yqDdcFr22
JfOggqvNlCInGj4sHKnQQXU3dT1q6r9BgLs+upH/n0uD6BqIH0uAPUDoXaaw9MOP8zNI963BYg/C
KC/yYrOLTwcMwJElSgu0SmU+A88j4k7wbqlBGytTWa4xDBEgGRRjJ3O1dW3enUNsJuqvWzza3ixo
keo5flKLLRecyHph3R5lWdfXGvcyzO2LZqM3JCY8vOJQ5p9CkJ5i4VVkCeTxQJIVEVbl09EjGO3z
Xzdd4adlFKeW+jeuV5dgnrKH+1kVlcELDHKDLAwgZy+FzexzyF00qjVzIlPeQCHiDOdHHJpukDe7
pVOU45u+oeqB6UBQ9Pc/c2GTAGhYsHphQZI/hRs8RESeb4q01wiqgdX7Yt5uqbdkEvN47nPSYQfO
7+J+rRdvQilkvfPpTnO+4MUEbUDk+WlN8kbS9BafYdSk28oDjITXN7rVpZWyBTW8826IFgjl4ju3
miUgZfKQ/o9t2dpFfddZmRCnoujwpqJCYEclRzHqdS/U0kI8sNtB4u3wKSQJewHFNPmjaEgJGfJ7
vn0LBSIiZyGoujdL9y4SMTjns4FZf9QQ9B+Sxg37ixd++LVrX1gkzrrbY70VDb2FZ+UtVET7Ujut
hW7d9aNewioacYguS3wJBPNUPrQ+l40+NyojnotvF3h2Zvb29ygJ0LJ17+eDiRROclcNhorcX3BP
+JfdvpbZroeTsc/LSBz4q+TI0INAPyoJo24U/N9dL1SYSY0cR9JsYBFap9ttWeHLlHyf1Qeq9Sae
DP9wUrtCBzVqyidGF2lEghBP7FV7oZYZ+54F5yGOKbfObj7bJYrM6UA8qlSFo3hRi30ZNP6ZZRF0
7L5auoED09IQf/kB4Rje0O+7Wqn7pa+EbeQTOA/cUO4A7v7tvawhyE6GyJBS4M6x4s7KVkicNKEZ
3iT1VEmmetiU/hxP5CXp7GZppsSW6jZHM3RP5DcRjGCMMWAwgVKS9tO5XAbI16+NIPnoR9tq30ix
pUG9opp2oBHUWY7NmRHyBKkcfTspL7n1uSMyPXlZiqbeIWYW0CUzQM7Yru2IXiIq2qSbPQkbweXk
nljPNl22+2wLTCMaUbHDctioJLVHCzY7Rgp9p8CUjsRiSOAjDH+aQ12qhLZmkUzDw4WvABGsPiRx
mzm1eSI9+ePB+8JbIjO2kgCf+WPIwe4vfudrIY4uvbYY2kec6XJ14O/1lL+XjldevrtsYeq/nxeo
OVr+5l4RPY3UkSToF/QzgzMjLARPAaqzOpP/U8qK0cUjT5AFS8b5EVaIvlRIpxi6TpTPEOwbKOfW
bG+MRfZiFTg8dK5Me6UiSw7+Na58q0JoxvToX57m3EEEC73HGS5vNXMlIL9LKlI521IfsSF02Rve
tdrw+rVKF126cwro/f8wLr4upJW2DbFHJ0jXS0c3bmj70NMCEQsA3iCbuCZuw7GYiDiPbN2L1u9g
tNCSWe7/GNiZDhr/EOimqLzFjEvks/MHx2sIuPsYZWvVDmv77Ns6wYyac2TWHG023ItO07ECEltW
6g3WqMfCTBIoN+DMUiIAMl+lKy4C2PKWBNjcOvB350lv8Cnve5Y8sKblp2IJHB8NjkjvWjebEaoC
aF0MRbZwyZJfuLq3eZF/5jHH/ptupPIeYw7vj35j5IBfx+L27IQKWofNv7JLaGFNZ3+Wy6bm0wN1
O1xbhXsf6GAhDSozRsnv6z0145EmjR2pu/j3VH+lR81PcF1g49Qfg9JWlz9yJZyojjkPiiZoxUbi
pR2v8emS5bPrpMVZ/lf2PvLTJMcqUnXiRKwB3j7DE5eydC7ZnHiEC/jKfkYJKlrVPyISRInByLxC
/LoYBPh9h1DpVspIIHW8wOirkzfBkxP/w3tjGebUxh6+50v34/lPBfWP65fn8qwWDezx7/D+hz8/
Sf4iTmDM/XRJF6OC/ibFr/itzv+VlQ1baZ/T4M2YeASVTEkK6Hp0LHSoSAb1JtDI9h5qp/fokYBo
kz84fqo6cJCWhtamSyh4WJVjQxGCxWuSzfhBfCoHNyJ27AT0AD+LpLJdEkfNoAy+LN9V8Nle2q1G
SAz7PDxwCNQtdlitCin4567LKn0hII601XmhxtiwHCpWKlRIr3/Yl9TmW9nGBroGMGURGBQ8NKQp
JkJqu22dMXEa5JU9GNzhyEJW/9iJnnDpcHzuNK32sHGWfgNGcrLZYAqTZquOkgpkjbd5KeDTNUSO
6fZ2UiJMM9jX0rX8kS0S1AK90AuJ57Ndr7ftdw+CeJafZZqVMUfj2c+IFOaajDreI/jwgArxoTSY
QM0fZASrQghrbbqC8kw+g0pxnPgEq5ealvtGRBSoMyDxQvSJspKF0cnRdvbY8NhXweIwtkLAFL4A
rvh/21YSjOOVPX6KX56hXU9ukaFxFY+EkipP/D/Fgi+DSQvDiCZjnN9TRXLT8Vqw9zp7dJPMuEK8
mQ/lHkgT4LBoFYzeQgTfew0aYCJazSNxDYDa3q+VCehYIpaKlRgSRLxO7I7UT7gPfHulwO5mW8ne
Y83ERRONGMOk8WGGYUqdd+BK4iw/oOxqy3EPDKtoykzypantudom6XbvFdG8jD6YBQfR8egGmMNi
4JuXyjpD3qylH4I+0k2aIeZO47ZOhfnxXGfzCBJjLl6dV1Ttrha3w69d55SPRLzvPU5gNwijSLZy
VAbmMRqqmzvBBCX8pY5LlBpaEdgqGJnRGJVY6dDBD1WzywQINtwWeeKo5A/tPf5ODg7wffYXrJ66
WC4rv+LiUa76GufGLVVQswDAjcA/G43azSf16j5jHO7MWeWSjuy1Xxr48jYv+rgs7PJJJNW8c+o0
ncVdXkOIu889I+W/u4kzXZAx0tOQ23n0VluJwUoheU1xCcw+ZaUi7hXNbnVQUuAJaW4Hc0+FLpRd
1aTbEuTaGTMnfh/2PTPUFy4reWLwMGk7OSHIImRxVihkiROz47EtyeqK0BRJu86d8JuwGzB24E3S
m5wu1Eyhr0/0kc3pra9czCe496izRETFEX6rKt3bSI81yA4jmBp3DL99ZyasFvVAM70uYjf32GAW
IwjwUgu/J7wniYVwQX1woTFVqZwGGQEs93IklvZqd4hGYTp55ciceCvSQtUm0DWb2iDoNPGrdAro
EjkeqSxKInMsCgDtdqXawriMiWqUT5wQZUF2DlpcFFRGIIRVvpeQO8gk8HIsf7lHJTHDoOl3LC/g
lL3d8Q96RCSDw440P/iOiI7g986Fqmk3CHaSq+ssUc3WoegtaAhGyYruM2VFdzjcBXaC4i0EXvPd
HDBb7DgIt485Pa4ZDNjCEUNyVJa/Zokg5m50yP0noTgWLnOx21YNj8MGd6f8yNooikCY4DNNaRJ2
Uq3syiycuWxg92P/uuKDHeKbqQEn29l47TV6HTYTW75TSs9ENrMUlIxzltYU2S9JMoxKjCEaOsnC
cpGpxgzGftfTSFPIi+jOadJzJxDLOA3e9dyRAqWeJLBG2eHPuCaQWwp+skPoKnRowAxSmxgCRYbb
oCMcTAQXUBj9AGn5TeMlYLqxE0A7K8O42CmZd4TsdZXU+gsNLLT0zO9NuFna3SxiLbbI2PqMnUBK
PUu0On14Y3S6fzkx/2Ira//xGqKmc7zgRCHD/P9ZVKII9DJsu8R1KqOwY/QRbmMjbiXw+I7FlJpg
En55YKB2IJhHaJs1iTQfZo3aAINJz+IEPydMb21I9v9zy8SwUk+Ohagb+T6dkYC9/0BlCIICsasm
2uxR3CxAHtAQEXM93rP68KZPhnbJaO9rb0vNBSWPkZoACyo8fpyqjUbbzcbzJcSQe/8aEh6eg48G
yQjArqzeNVF22LA2c6ixCHr3jIlV4KaJX4cF+jHoAJf1bSdsdmvvs7YvWCcsQLkzu2hgJNEG5MGp
6HNzF+SdyyNlVhz5Vj7ogYYyCHov+mOB1frcO8cv+/dWjwoXTyei0IpxgOF2vadu/WvknNK2FJOr
uptJ6zCi5z6rzOJSmvwrufLa3U0y4B3Bd75md6SlzXw7bvEs7cgCzh7acmNlJFjnTuqAtYiKfT3d
+sNJJKSGGQQca1CCvQOjbuBc2fzwd0OvfRXx5pY7LVAXqnwgp1kUA9rzq7ogk/DfkYyJTT9YQmtO
olO73czJ269R+tMgpdBt/bIsZKcT/15Bgx5dNzi5HnK0lrVyOqhAv0KaFAgbTjIZZFz8d6sb0p2B
GxsitC3QFQG5/YUj64PU8vtbBz/NPeMpYmOqW1H+ww4ZmNOA9kDfi87Fkoyo1/ZtBg0YgN+id5M6
mNvYEcjyXcI0Ut8b3Z1p9tZGKCXYVsALoF7ZnB8AuD0RDD9gOJ0LdIqNks1dtELbQEhBB3MN+Lm3
4undnB47k6a800DGHKHugSE0y6o8jKVsyNpm0/g1vgFsuO9x8kbTgISXqd8ZV1b2flDA7yavx8Be
P0FN0SF0XANVF4Nnx1oSkOAgg4XHch2eJrC/6iwbMYA9EaGuIHJJXCHMq5eBx4L70NAQj9+5+rjm
VSnxvlhd/w7NbliSWyJjS6P//jmqe2tH3eiiVP3DHTutXYbF/SCC0JN92mZlKNBS0DooNbMH66UO
vLHQLVmiSDXZ0OxsOOg1zEepXy1HO/KkfNZx+OoSxOvt+J2KdEvoPpVitXK9WiBPQJgTHXDI5ENM
isRayY2bl+PvpuXUHpLuILT0bydaW7o2rl0mb3vDHwPzBkwh4ufwldfT1KsV/R5BWW2cSW0z0Cqy
zsLeHm/Z8/56Dgx+o57CF7g+oNbKgf/8dG1pzCs0BEGgvA5q771WLOKV1hTn8w3tl8VNMEGTzAfo
IoeDWy36aJRuCsTw3m/rYRpqcCZ79dFlCuYd9sygfcsZvkt+KkBnlSAxFy3GEccunlr5oj8/kwvm
r/Br5Z1Cu+oYNqVlleUUbJLd3ojquPOncdJgimuZCdNFznGbsHkD7Ft2x22PMiDg00OvdBwM2riy
3YH85GnVt0gUspteMDgvBr1R1h94cIK38G+ywtY2Tgn8VWB5rlZQT2eyiUzUYuFJ30kP7UfTmnJN
JYut3kweYpGCQc23v2Ss7Je6si5pj95MPnHQQw0wYztTXDp25Sp3rAJTcVm8cICCswH9EaHQVoPN
I4/ie2EvgmQKiehGoqKL7X4oXgWzPHtrIGfFwTW6wMfaL/1v4CQlpOuhVttm9iP86LlsqhzbAa/7
BIC02stWamNJVGIJBMD9tPOTdjl8bDm9dlx3AzmF6gb6g5nwwlhAyZJhxeNWd7pn3mWTzcZ02FwH
YmrCT7BKYeYErUmJNL+y43WoqTpvmiym3zzkxUimhZ/tK5SzKaDOCY7I8fFPbTSSHFfbigrsb9NQ
60fFZ+mqYcpuSvBBzoGEo7SHr5A/hwnuqR1/cyhdlAWbj/8+VJRDSfzwlj9uU/XqnXCwJx+kZpvF
Yc3AdfX81wTAwbTFL0nm3JHLZ3X0UkaX9Cq6Pz98PAczpXlx4WnNI2YNQs295M8nDZupCZUovDEL
n46ZY9Qe2TbmYiHMtycEs6OsAzlA503vzae+Mfh+IoIyMR8ePUFF4HmkiiT79iqx2XpwDH0XCU48
ApJ3+lXmJNHZ1A+7qNRH0mgNk1BjhpC7dw5KV9ywTKOFUPRgDFnNV4S+QILYw3zH428J6wXE+P85
X30v2JO/XxhizrMKAFfsm8jPwDl1T+HZsubiiHfll5Va2QegH0JMXc9xdLrQRUffkngPKm2zrzVc
jQrVdyB54mzdA7jiIZfsDyxmkkJjjbNh+YD+19PY4rAM/kT0aQ2VBeqwIQExCHugguheFZMcQhg4
lgO9g4iqLqUgPHYGjTXbZlqKE/FRPBmQleofPPu6SbzqRgF4SrobUD5lr73KIDXwhBiZZqf3tZW/
9IH3r6abUXBVKgHLZo1jHGZomH3m7+hmuUpnDQWBIUMp2UcXaTT8AupKxFjDvUOEUipe7/NcfDqs
pI1g5Gn5xACX+Ts4NyICO/9YSoD5y5Dx3//qqG+wuKQvGfs1APq8+B+eMGJybTfRp+iDVJ8nW3Zw
P6IoECleagNJMWNbz8u905LIDRZ/pwSos9BPgRvzK8l84fg9uf0JktNF1Q98jfeoyp/gsP9Tr0BV
KAoc5UNEsXmYM4jlJHeliR4ouJSD+quitXdtwGpkpJWTOTw3JMMPjnuikiC5TRPb1hY7kq6bsE/h
1LT2OAxdocc2LXprF7gGtFhox/isaFl5O7yjrkVUP0S2Jp3x2wRY2xXB3Eb/dh5ccI7hLyHedSla
4l1VaBGsb4DLFDNRgKp2NV5CHil1YkZ61PQ1ySXiCU7nS1Fi795jE+jOVohVRdBVlw/MCUqrygpx
4InBWUF+Ywx9AeegMmfGex3gbabUtCekv1UgwviL3nT/FrRn8BcOSPkDiK6niA52sCPArDLolrWc
8XHYvVw9GAG6MFrjmzn0U8evIEAafn+EeiJnQIX9jJ+kqEcgG/TIU645LQNtX6+ChQVMVMtQrtWo
zo69HLnRG+lLaHQ6w8YfNzstI7MYTMLCx6iC3mVjls3/oQeCkuBu/Ie9BkaTWIyh9xlHtXExNwn+
sCUdzxnhcmveYZwja3kweAfPHN3G/Gp3vMlfMwimsMfNLmk+NTEhTvalLhu7IA8zL94VBHHWmxIm
a/bLRjdB/uVBNHoO/RZCdTq35fRV/KzzQotjMt2AynRvoRLHg9jB2waJ0pL+BytvewuMBNb+bg0C
+tpKgba0jAi6K0aOyT0WDkxN2AqcmPRyXleLc6zrvgUVK+Vog/9rbLZPsc4WFgsq0Y/I3G5pCyEs
e8UpQGDsk/5BxjIXfdREmq4ZOccXAnHh2PEnAmwgKOxMerkcGVgR1V7uhk+tLHzDbZn5xfSlsfiH
fzRh++Hvkn4Q/VGpMpy+g/QLRekaH3ETiCmQWqgG9sNW3UwNEqnFmanqgLlDojNOChHtKEJ8D2Az
QiQ7yD9PQSR2HxF4lu62wThI/sOijc2y5TRAzRyrNMX0YxO3ov01rtqFeGGt+7ljo/uXoRSrv+yU
E4Vf4pEp9Lx7Q7yAOCmzZMC+TveXB+N2Yk7YBl1rffKloSh43LVzjDh8mDJgeyjrUVnAJBA8yFBh
dLGA26s14FgKtui7B9pVpdKBPYSO/lxyAVt9CNuySWN7HpwOaMXUzue+vQEDUPf8DTbIItZ4kg+o
41SusYY1tppNTeB9BeU8vmfoTUuvpGeMDBnCAWR+MrXluITvdsWrLA6+d5FWz6EpmaTc/4bZiTd8
H7g9gSojOlxx4yndbTE5N+iow8Ks3NnmgAAQGI4b8XZTilJEfvW1u967ktis2Hy5tY19so1rH0y9
F8LlHFzxpk6dhpc6XGT4V2l6iSybiA3NhDwt4PTsLAA09rVC0TszZTuTsBl6dla7vW/Jt+eKDUHo
8B6fR0C8iCGOloKH1khQ+dW3Kxhqqo00LCjexuG0Exx6X3W72QPiAIW4H3O4cb7MSn7zL6e5Lhkn
w4ptdZVETO4Z6vtTUUpXnVqC+ptEl3QF+Frq40DPYqT1HPN2nwX4IzJ3hxrLZkuc9H9/hqSH6qz+
4ADuIWofRWSB30N0Bybell+GtVuLfVUUAu9w0b+NiDwGGR46WA+8fahkBAQx4IKyVlAydZDeTSqK
hu7HcTrMCJd2sei3lUWARH48GQASI4yRiL1fiDSGpNHEEIb8D92+R1ibTBiS85RYCyczSZlDH2Rd
GuvJ4cYvZ/anJ3SRfGshFkVF6YWgsg/lDmoIOqJIiOXeyDV5velnoHlL6m2dvxzrBQE33YA4/k3A
YSp+FcXB6dmhassGcfB7hvdTVuZFqgMJko4x2JZ2LLfUMfJzFOXA1J4bg1viXLyww69eztW2iHku
8gmkWo3ePlypbHlgMg6X9tjtiuATmF1bJxkF07Uo3BZaEiMDJ6B2i0+ZLzbuwXgIvXoMO56V12Ju
wXopLli/ImdRFoaXB1UqqbL4i9QyejfVRm60qbIffxzHcDXQK43VYzpQcRE3/2jxc/0Y5Zl2PnUQ
ladmc6MpctT71l6cP8gJ7tfFsc8kKbVh/4gNLSUsXrX1anQmyjf2FraGb0LQ+gaztt24nOs1yuVe
2hf8THXdz4P4zCzlCpXWb2yfn4jgbwTcCDC8IPQ8bZb/B2HcUkOXATvp89hDIA4jwNm4Pq6WqsUS
MpyUBQGzJhRPo6HLBbfFB8ziI7aZRaWX480FWn7j8otZxO7nCcnV305EHccrzst8s362oihY2f3E
mk1s3sBM10CdKbbjhX8/llGsDF3P/IQvCiQj7fbizouyh8V+UxIoNUNHUZz5+jYdHa/dM5EEMlvU
woHDwWpIUjpvctsqWM9jnulaxAka4OrywxfzR15zbkQ8Pfj8DCR6f5CAsPczgu/vl8kNZLaD6zdW
eqsEdVMIrkhQqpQjZCuAmX6ohm29MVxqzyRz3FYdC6MLhPS0h5V5KyoLLB6Why8PMqmtnELqwdRX
mv3Jdm9LL8e32nPcz1bY8070RY74wXbO9Y45TiqdfMedvCoqfTk3SPthT7zSZ1eaJ2C1qQvUCKY7
E5y3QOODtLwnSUu2mK4cNeSkUHb579EzYc7gkbLup5P/ghpxMh8ahp/69E8apdaLl3BH5VVaYwhz
O1f/yetyZQWBg2f6u3RU6vmCuQrZ3vTQrBR5RQm6rhepJQkT4UyUKsQEUK9wX4dsvcFcBjf81Ge7
OUATJv/4J5e6BY6zR3YyKa2Il50bsxAhr8jQNzry8P5LNuXh+FRF25N6HJmn/jxZ5cFIUIQ9ifuX
L0Ri7fUMJwHB8VULqKh5LnaGaU39eeGZ9iQoGRei57zT3wpJRBGDsa6zK/uZjsxs3O6oCMCNzQl0
dOpl7iODOakAv08LOTMmp0Qrxj+bMphZ96dTMvddoPXbcUf26/s2slHt7ioskxQ50riq27GmlxUs
ANx92nNtPHFyBUytzh8Js/Hb3hCiLiZeJyffOAoMvld6IB2Oh5YCOD4Swg94DvzPbSaZDfSZLfZl
YyvTh76rqsvMKeaSR+z3frW/hB0StMxuYUu8nKxBuF/zsVhc6hvOnBLi/eJLTf0BMbU4DwAKWa70
nOQnusU9uz98fuC5sInd20IpJdIa9VVVWOxYNZq7EZh4sa/3AXgS1JLMbICSaW3XP4FLt+QQIoAC
D2Z42vwX7CKkCuPYkOSa/hTJJFyiwrqZl2Dn4KohFDHzNkoqUCPkjt91Lg5ra+7i0iz/NUl15ECu
/yTNGcwr08pktkXxAtcmneIU2dgnieHS6oyPAdqYJyBcEnu7fsoXuMc0V6FW1GDpJsXXyO92WujF
+h6mLdGxIR6N/tp5Gx8ezKnZ7c2s3QpScSE0vF5zTkGuYnwMXUMqPCT4kU5hZ5ApeIIcc+qkjbN2
Nqtb9TTjZb3VePRiLUA4knaSKq0Bam4SV5r2ZP1NhdE+a4egd/WoklOt5MPQlUJAn4uH0uQ0bONe
koV4zwWzAYvEfDBKibAS/lV+EdB9PAjepyrDU9yEn+JGAJCJbHtWE84miBDP9mg90dPQtoOSIhjo
BXLOrTg3LKKW6LMOXsrWhiYliwIaLX3E6JZjXYqKQEv76n2BlskwVqWxiEBqmR8i8M1SLPu+e0P6
tXLKsBMLExxMBH/0dfltESXPEj1KqFEbsdVXTvozXv5u3MTYNFwMIYQv/I/bEBOgLNYDL/986s48
+APpHknquchHIBq9r0eWQ39I0dQOUm+DM8s85VgAChM869KeijhqTeWW7IwF0Aj/IsWazoCR2aUr
Jx3psgL64ZqTsoK05TcdkyrDw45d01upsiaOXJvVDy1bC6aCy62nPXV2DUT+vUJ30Gr8QKtrq4h7
veVdp+YOi+LC05jUxvtVB6m8sqi8hKAO5SWaeN4TAuHRyz5OzT2WqLIzhTCvJQ7IHj3G2y8kTJ0O
9zn3Ag3YBNVyhSlE92xvjE/bRUIjt8JfzO4YevIdhCdUpW4yCsoqbMbcuU1nwPnw9YMBFYFQQ/yu
JMgC4J4XJ+7eaQevjMBGZDPFJzX7wP4wxgBy7SyfDgG7MT6eFBJjubqu9a1dIMVkVlVyibyTm99O
kwUGwVhnm2sHftFbPX97uc8b/E6k5Cxccw/ecRrxwoFifyyQvDpBnQbXb96InwIcyDVUgUCwrK2C
zFwXAF+xQx763xck5PovGz76NVn4L8THeXpyNeBXv4J/rixi7Xr6SlpRbvtKe7aUfYosHyCNT8/K
x56f9UaM8ru85Iln0CHZeThVRJepRLsdtPe8ejSNqjLQv/pQI1Q7b7CTGDddy2T5sXGGmEBBXDfI
UL3lGQlRpg1Xw8VXeoLbFs/PME6M+7IqQDJjulMS97GwfNraDO3/t1Cr4ultAMlhU3CNTXxO1kK8
K8f5R6mPGSol7/96uM12W+3+KXWDLGUrDwPprvqxOvogT3W6gHSK9Q0E/DnHxbBo0h+K9vLMpXv6
/AD5gTRrc10XF+Ft1VOsPruXemmd+JS0Z3WkR3sjt08IrJIlp66wCRr7ZYh/wVD6RlYGarpBcW0t
2qALAsrrF+HuoHKixFcOVnRwptxpt5veVtV62fcp9/8RXlj3bJdPh4MXE+j+Hu34dVVIY7g5SFia
HFp+HGHAT+NHlEgIp8n+Y8lFnu3vGl+fNKSxQa2GK+MT8L97AUUFHbfOeUhHupW0oaSs+df5i5lu
Wu/KIKtnRB1qHahbg/oCtoUVV/tZJL0BtPwFF6a2wTMQ5M7694nu55+LYXJhSBEIowHZSyGJWF59
3Ul2rTiwJ28+ZikGdaXiw3NrWY+sMjKZNcl+RGeUFRVTB+M3kSV4B2iHU9KB2FoVrdLgCX0MwBsa
oy3ghaZNG9CE6cLwSodP8eo3lhvVajjlaEslXSi29h5GPA5gNaG7Y0E8W0uTkYXnXj61lAbgZyWi
jZZSjg12wrikJ07AmLmmIUx8NPfO48GZi1HOo/X80zdeWIQ+nthw3iSpNH3Ajw/LTYrDB5ERvuFb
RqioeyoFj5E6YvICVFDl8Nxp3a7pDLX1ySoVeLjI25tflmN2lUIjaspvDSrSSmHCNBOD1lUuxM48
oqpjSqsyYSbZc7yZDgxedzKErXsmWeN4WxSArkvcwFWvlyqHsegtCQn/eu6TaCUQKdtMRX97zZ5d
Jc3DCYhlxo/KH5ZRjD6ZfNI//IrfXgA7jiaqfr9a4XgAQcpOmP8U28RxDWBNYYH8EZpZDxEtZVFy
L0XcfSBKzWBT4K7l8emG861eIQH/ahJ49dZllsuwR8hZUglXPTbMPNYX8UwAX/Cqrz/C2mc4uODm
LLfQ6iVrhQDF3F2gzYO7c+7KbUnsvKtlNND3YbqK2NiMZTaeEkxefwJgyN3C1Ux1CsdBxAIMNZh4
o7shAiwyB63ajY7gdUnPVN/6UiktK6PlEItiUvRI2riFt+hvaVbGSguWANCrnvSn6lejkx2ElMB3
04R4m0DNmrTt7Fe1aOy5GWDgR6WjHCBbLNkqaNiF26YJufy/qwx0MpKzSxiAlsJMvKUI/5JrJv49
6tYnMgeUVnC95PQ7pz57zvzfBGo29/KhLhErl4n9+8Ka+db6wiERGio/Pui2H4grb8QL+Ld4lc0n
5jZ4RlB9Qhxruxrexxw8tJ35w9Wri2wuJjEYgLObYzG5768dj68dWxxXVmpJ4Uk+oGIhXcoSNk7d
ym+cDNaAp26RiodgkUIPlCqePuRUdvVvQQd/45HpDpDryMzgMWYYn47kqDOy7EI6a/G7L0+P3w4z
x0j6OSGOcQW5fkDj76+lifk13Z0gIoMbyZEKvLG8EwUbrIvuLKv3omT6BvrKcoY/iay+guiBoKbu
8ySSTyqiNUAnkqPXtd4FsMCdD7XbNQciaqYZhFXQCXNlYC3VHQvNc7xKrOJI4Lmg6pQztMgOd+oX
pa0p1vn5OhX0wqHqeRhLuxnEZtqot4WqBhgfJ4tHSebXV/JWIg81KqDEsp3v0tdFkqedToqL7q/M
jBwQ2/gZofbBPQ4JgaKVgl5ubVfuvNiTxzmD6+OZKECXShN4LiQld29ti3Whs4BXCO0GXtHJyrwT
1T1/kqD6RbcMsHbklCgCdE31NZ1E+W0SjkqmwzXITKa7QeIpaHJfhgIw704bJIMlRUSROI+KsziU
JZnfLE8JwEGF3bbm7M682+q0tJvlAc7IGmZxAqfaSqbBLLrxt+uQu9gada+gNSCh08QvJkb8ZuO+
p9QcQWa7St2GtOrdnO+0mYO6WbqVuhK+YVELKnDiA3N+VrNhN6ZiF66zpRpQe4jZrH0OYJNqKmXQ
o1jyVHquBv097P4jw650JOGz1jRIG/C8o0f3y8tie9vkjp5WxZ7bURoquvlBuRXLs4uuewXVIE5e
cDC5ffyzucqV91fZFizCIqaMmG4PJOfipWSDjvyDlbHedEIIMwRnpk3WzpCSHPp25GaO0C0ea2st
O8YESnTGMNrSr9IBMMfHGCO8LMe/pw99VABQH3HqcNUeIJYkZog6D4wEZhMN4qE9I0REDaW/mhnh
IxxZTxoY47ySqK5aoAVPhJMlCRhfZnmBcx51JSzgpJmlrruBd2uFcmIGihAB1ylQWG+eGd5jKE5N
b2x71e3XU3pgbCZj6sjYja1Z2g4gjdrj7LFOD6KRQxnCMe+yOmTjQe4Lwt5849YvBNSky658UddN
P2okairwiJfwHbwsYzKOJWZ1Ewb5OP+uu1zMvnZVKirVulfUcq50rgQBLCmclywXstUvHZOORLpN
z+pCc/ZxEyxGtFTqGJwb4Gtu3+YvZviYHKFBGh1XQ9QHu8cHvf6w6HA2rdxHrNnavrG16gAD1G+V
5wMKjs2pLvfa8OFssLedXhLRVQwdByB2Al6AzdQwUkU+SrfUjABkmnVTqrtU5aTn8eG+zLr3OuX1
8fYipbZYiymMOSu0EeLwyg54HwPnP2gyRjwt1MBI+ft/jCR6+yPtxbUaMxctl06OOImaIrs0iAr9
bMUq5RE8qOFVHilfi/8WT+4iv8Dw/hLOnMFk4wjvpkXnk+/Hf7GsdCCjYXH4JyqWCitFzyHpH4lD
xlDGmqQx4ydWZjNSs3Hw+L1N2PkTbwODEYijiQ9uBE7jpkOGPvrH4IZFiNoc9WMqEp13yfU+R6ON
Y6nCLMtvuAu23QxLb5iRFjkwx9scS4ulmbHGRj0C0uL/jMgB9HEVQzNWl+hbKaH6cPgVQOBQ3VV2
gkPJ3+AdG2XewPRKBBeA9Q45kT3LQAcaCXz7LvhVIBPVUMl5WKjb/LjDyXLVki3NxHpqCocPnROd
yKeEnF767HhHgzjpv/wqTyK9dGBG7mJ7MVTt7K3mH2MaIuoykyFdADRdtUBgRo0xS9o+0XKxHz0w
QayeKNwYwUe0pTiw/QleiRQtrHzuljW3L32uFe6LBonC7iSXnAXow11uoEut4OV84La3TY5W0tMC
VZfN0Dexyqmhxv+gPr2i7R+6MeQARYVyN5wZfs+UhIuNoQnN/9BWFlqBrzCMza7Rhg4AkdpQWaJo
mb1uHjtnnkEh0SA/ph6Do8Wq1pRpVOcBVqkXdMXwOws2CforEDinngRYOiZodhShkINW30aH6wGK
OErXTw43IJcGK0UL59Iy2YcuZLi+dKPHIHgEbvo5H9jG6KpoAKvh6H52vFSkcaGlusjwXhuqEZrl
nki87fY8XbhBiqJeK/OYZ8I4H9eCOXlVGJ5SEhTdHY50pdy3e7u6GXWtGDzQ/hnXJXbatS0BUfv/
UKhLgsGc+9grslZuFPQwqvSUUombEX+P9xRh48uQddA+wAjjKIe8+8iWbXUPWjpzVVCNCnSxxnkA
WxWzhId1ua9SanMzzP870X53Atgc5TvfZkr6lWVH4NOMLk5WAm1Nfcs73uUJ5d9vZ4oEabTfVXgf
RfcCg2EzcCVSClzZLoIBexYK5vWTOLtwxSSckVmTKdu8qOH72g/K3141u4RBgkyNFp/jYaH5Xo1I
6Q2qzr+9JFfWUPy8fpBoCURYYjeNmjexpY3ahOfBL3MKzoImLL3lltMdemuPhFYWz/gr7Vu+qPh7
309nCUVWvBFXonp56nzDnKrR8TKGoYmTS6WkhQ0XxM9fZ7J3puwVvav7cLTfM3K67I2MSZPlgRf5
7gxCg8goJ9Od2CazUxQqoRXqT53+v62LHjiDwaS9g+2OY+m+I8K+NMr49S1fg1qw3EfuJUYc+dgz
usmRuDQ36mhsuWhJoGkRfuTJ2ChoaRsAiNQNzPek40BVCdy11+9ryND+OtfBNKBpT/QMj2IFOEJ/
WixuKxCcEZiQpUNQi0vYwOvKEBlo3tgU7Nqh2npIJjF60EvcahViGIyx0YN0V0RN9bQO6F5E36rI
QLycSAUOW9B8HsLixzUPHsG7JOHGqUSVvDTC5FPqScYp+Yum58F3tg/ajmRyvguGjrA0iR0Jky/U
VYzhzImFDWcp7D4YHuUZD+Gn7jPzuyFRCOvB3tG3YcZ+h8/ODvlGd4ny3uZzxdsb69K4RFSUieZN
2FDD4w+NXa27CNRK96BmgB0nL6hnF62wDovr6+hXb4aiUG8bai4cCgtT3bY0Q9LSNCriTafnCzUh
Rf8W5xxc3b3/WuQes18ea3XPT9WfU6048NTjkD482QLELh8cZhmr5fhCh5KD7azKCXfJEhb3rnvu
SRSwP+DS5bRhv/m699ziUzRoBSYwza3M5SfczqHUJH3aSFd40Ul9eOpDF1zCcVnSy/kKyFKWlxh3
P/xK//1XTnwp6eXDpIdGmQx2ydL9607E9P6HB5xsqcSlE+l/fu4Ktnfjz/3rnnlsj7mhYl+VKhT7
ULaZAFmmbTS5Gqb2scDhJKwIvjoHDKU68KWrKAQpS3A51hhMCazWVjCQ7zyCCuN6HN9PqiCuRHNK
TAouzhqLu3ssMENQolZ6KP83n1xGx9miWqPFVqiWIIPdBSU9yd7hAvRyzcvv+oDD8j3ekTVbCJHC
n63IiX2LKxi1vxTOulvTN/w8jH9jFo7Tly+HjPdvjkjBO2zvJ/IGVaAUsV0a0a29k3zNykzuJbwj
rnrQmHYWIoJlRMV8HyqnpCuKXoW/NqhXx1gUNvbJJTopfAwXZ4dIODrMDayXIuFhJ9VBN8L8VfUg
CeT51kAP/jpCRF9EvjSSM3lwy+bwVhUuBWAeXaC1y347nuCXsgmQhMZor6A3A6CmO8j3OlY4kWUf
2x/lmTUFQRZPKOtOJO83PydwL8/5d3FVKI9xlIW+ak3JGNdvxVlojpSJ8UwsSjR1sg5DA2rrb3FA
gTUjOcu4etj23pBePAcvgOOKwuW0fquPqn30I8FMA0dFO2pZGyj+HEIcAJ5iHxs80HoEF/qkG1Vx
it6PWy0h7/CkFihsuoiMQcSYPj5Fti6ee2fX685DH8jajX36MRqEiRF8UvRBRl+q7s/W2f8Ou0IV
LSVTAUWN/jQPbLdu5jcr2Nh+S7VNillWBF4yas/LrfdXG8Iu99A2o4L6O6Lgl2JC70RaFNTFKpSF
xVGsWz3ieXii01oSHo4swAfAtwhzH36vwxJUruTRlHrxMc9CgtmcAl4hcgu7MGkVPRBtM8egJ10G
EsqiCPmlzViO4jiutt1KDUzPvcIr00x2A/L8CImzQYH2ptPlzzXigLMMFfhPw/2u3oQg2m6TMxBK
uRTceA7vQcRicvj/34kKAyRwXrrhUo+2UgU5B6iOrNW3QOPciU8gx6ChW1+Jj8xIR7QwvlJYFWTc
UFFffompyf5ZNlpKXMBX26jej3fH5IkDQVi4ftyBtlD15hpbAs9O0EL+5xbXwF4HDjAXxuAbA7ju
Rz8Od7u4iBduGiMH2oILQ9nswWRkEOaMrb+tAJN1of6rd1uxekhqco+fuwzvy0fOsAFMWHfmp7zl
5XuY3fd059X/Z7xvA9lQOattPuPRN8kdn5pxxdcU5livTESBSU4cOVXTALvagbIw7+xDU89riCr8
rfyDDrLUiAEJxgurgzW2Gr9qrlJhiVbRNY9bTcDG3zwniRGA7zXwxGcdcCcMY2MuT5nzEkunwfLj
SsfmVd5RPbzg8F7IqU4gXUydNk2xrF+nFA8xvGeEy4/zOUP8irpxEAxFQRV1L4j59TStu6WyoppZ
NrAj9iUuccJaswm5AmkaLUniS0A7e6hjnZGckJ4TeNR761AStTUKt7qYkkJVKYLX9qCgafpyGiy4
HhNO+R4XJ6u8l5PeBHgBJiGfamp+yBRVykOWV9aGs64vKmfM5FacSOBaKlPQRM3SSsthcKgsl3TU
XdZe0Npw5aU0lxv0AEFn+/BUN7T6vZZxTwrGdg9lxj9JiS87LZk1fKNBYo5F1lryR9FXnyhCh+Ff
HeCZN62SyC90AwLfmzwE8i3mAaQ6m02EPUD94NXv0xGPxK6uUev0TxolylIbAWpTA9wf6owqM9yv
tNOeaq4KH8nr60YJdXgT0KzToGB0Q/NaADnmMHVPqS4NrrgM4fDIvuTsmTegAc6rWu1dMS33LlEo
dt3kSQn5j5ZuhMKVbgMJdkxMTso+fKRrGi8jYUZGbYZvIe21UEPyHF2A9wN/S/iU1jDwCmF7ZV12
9phOHMr+XUemLEDzequ8BxFS7qbJ6moHk9Zlt13X1Knhoz7pQAy831WFMnD8L7InOade5sh3tjCD
F2lsYJVefGZVd/DDZ1TQApUFiQW3c1nt+/CmCJezzvrPtFRx+pnQvgaqrWdn4satHuxDgz1gl6p2
XI0NqSNucjl+K06RtskBS3m4xQHVfOksGXRMK8ZoURy94SKMApz5yCe5svwRB0iCOSSq7U5q2buh
ZBS07hBL/ddxK7JaNb8of2yBp1c2P7uJoGhU8LcjqbLCk4SoxdXSMTo1zEtmXv9yHFuBQGjjkcIu
j2LRIalmOOa/chhY2g2VCxlxJzDd8VKo/xZn+w6aT5LXvSIA2gg5tl8g3M5AZHTfnprxrG61Npvx
MyxjYxszkyCRLaepLruAcZP4E8CUyYOGebYnLQPF2YYsaEzfd2ZOS5yg2rLuLywR+4HlVzFnqwLD
vbQD+7Zgh4Jiq6LEd3n7xugrNxryaMRPTHHUtnRV3epaWlJjWhg7+tXQzt0sYnmwwR+Sp3Rjzdlb
n1qvh5jhUIN20xr+gBouA7wNqajTW8yPPiRvQQctGoaQbjMX47aYJEgnuRIRoCy1QdJ7FbEMRo4D
1P29z8RGE5cKH1CwkS9bSu0IZ7vAtVWHk5DUoVv080NkqA3rbGF+Y/MxWbUeHJTbo+/IamixT77r
041H2fg87UrIBs9lF7JqC+VXo9u6nGBKoCA7AwH0oA+8ptpQtGvHMkvysJVzctVTaXhWtLueqsAt
5+YlFkV9fJ5DxsHWTE47hmSDDsiNGm83kzRSM2h0edZ2WcsMd+JSn7aVfa2l2A1uu1AiouRMRw9K
tmDkvEWTHr+g6HVgoWAvxku4GMPr0Dz5gzTmWtNAvOhmpkze2OHZA3QMPCsRqst5u9r0Vib2jzQi
jQp89G7s32Jy/XeZPjlipp4XUEWygP2fh/lo0P8/5MipQZXfoVnjwoNK3xlp5Fx8AdBwXdvgWB6P
yUscDNCuycxDGEgh6VhxciIybqFwJoEZ/QeZP/if9EmRDonul4Isj0nO5ZDgoi6xeY5uW3iqvLgd
y2feTejxKoB+QoJVjZhEJGJRSCq6+Or6+A8OvBmdzDWoFmnnrsbJ/QLnnjUqzWl/MzNspCN1g97B
cY9mvo01jZK1mXFKLuLN6opSCjrJ7UqhuKbPMFoXVQVRq+IHwAwQfHLdzxJTfDlrtI8UaIa/se62
+sUpckrgE/qAy9eFAFjnw23qvkjO8u390WsvLkggMoRUNsBZGh0KI+hy7MeUB4lplWua73w2fyx4
yYgaLN1iKDSR9jFjdNJauDJQ9GZC3/bl8jlATs2jgm6ONXESsEmTMJO5Vg3AjqBc8dNcXy7Nyh7p
rNsbvtZ+BLJRvPuWe3jiUiuQlMcIu24bvJYw1KYF82sTPVKzKExEMIBvteOsX2X2N4EoagVKalr5
Z3U5jBEsx0DgevsR6VvjdXeSIKAr4pE0xWIQD5xekbQllkyF/sSevGejNTo6tiM9wy9F/iujm+jx
83XoFf2WFyXBORdv0SkJ2INXnw0KzH9GUqDb17GRQydzd3zfIFO4I2fiIG65v6Hw5+GPjgbWx/Je
cPMc1ztJw0l4f2VV89rDwsGnwcDG8dOTOkFlIrqtcWz18L6zaKi9ZbKqrqzjkPlVlyoKf1IsVzSC
YsSqtFdP65dehTIkAlFruXB+LrUffqhRkrxovV7PoSEwYokLfXne1X//nWiApoX1LUhWn5gR34jO
luAcO9Tly0T/deS4oYaKs5mWQNDy/gK4gjAZTNpaI5gSB7F5qrGour3RO4C2WQuAm/Bf098brF7K
4gnIVwVDIHaCCk5INIR6c5Us4Wll+Vh4amuIK9kk/Jbr+3WddghumtdgtPBoAUZUOHh5rJzXTmvx
bSSirNfhuYnqiwfsE6nktgVx7Jg0m9lQPVfClBs5moPAW6/exFl+SXeyzofwskAYZUL0D74ROilC
4Ie+V7a/s9OqnJ7Zgv276o/A+rLn3p3pagGzp6p3WnuKy87gAHPq/ysb1K+SGdUZpORm+YRBPzuN
YD5H0sMSaHsZKen8o9T54+w4eH42es1kJwD+FG9vlBRsu4+fi05xAS2IE1wtpLd//+O8v5GucMvA
7HqjrDX+8LITTsoGxFZ8iYGLIGqqlWAXq+36epdzs/bPeiAfrPXMFR6wesnsKfNvwIknbvK96B7p
+KSYj4yLohd5Qw4r0x5vR7auHU6Gu1MXgAUXhF8PEZ6B1V5hn8BEqbyB4UsTgbN3Yp30xmAor2OL
2urB3LvTvwN1WH5PB3b9jod2jx9fXOSGApuExwRCpKgO+JiMh5EmPhYxj0ddBDhBsCDLm9lBMLyy
ue/YabOuAYinbK1htAJy3nweza7M9CR3xx4bTMtGtbhCMsnk5BvIyNah8aBCjGyf5qaADYLFMv7X
CfHzU4bIxdq1u4wytuvmFPVGBRoAJHZdWgrlMI4EYVMsQIW6D++jYC2qjC+5zevcFeZvWErj6lCf
hFXJKkCbKjoFloHQ7k5LXdsTO5v4Ex6Tk3RnK5fzac9BsMeRotGXFylF5UDpgathXEXqrdYMHk/G
zLvj48mn9n+7m7IuUfM5oW+ff2yNbgdvxhK4wdk8Z5B1Ln7Zj8CAldyFwZrowASjK/y88NBALY65
mSuFu3Gy5h4Fhe0uiN4c4Tz4uPouVeTMgx6i5P1tJcT/GC3G6SgM/ctbbk+fhh5EQ3t8IbcVVn+b
tECi/D1wchJXYVusf3bskBX6p36xwuilr/GWEUcUty47h+L2PBAsTpsXnvgJ/Esr7dOr81z2+/8i
WqnmvBGd+PRIw8q8lEpZvajvofrjF5K5QtBm2DyGr3JNJ0m3Ajf50Ih2QkaSEqBKWgBwanlTM0zH
1z5M0NJnHFSS9E76IvECGhgiNbIUIHleUWra1lX+96tgNtuheFJ287hKDF71DDm+vxf4EDVJKeRa
1w4NYig7vPSayk5D2i3WvDws4j534DvYoyD2w7bLh7YJ8xnVFDvcGxC9qMWnPPxnzsv1YXnP7nIE
hJcDqfZvRVZIx835b/BlUkP08Wi7+miwuVco0WAL/Zu2WtjWJyjQyzETiWlD8KSRM06yVC0leOYT
2EVwErKQB3NpZRWuYPnTUTc9crGrtzMWROcpMKOdq6oIXQeKhmqpLU5HVDwq5NiR923gxbnSe5qo
7E6YVii+a4qZLOXuwCz2PbsZEuWg4xbnHwOYgJCqUe7GBZk14ikxX4SnoCn3JIZimA1auvHZm7B7
HYXjLaz0zwekJm+CpDvq/N2Rq4LukwUT2oDuOWPyl9Et6NM4DdiOqZJFsFJNEpOmMbjmrAVlBG8f
FRrpf3yxIWgVJPLMotdlGYip+HkueOhh4IfwXIUMT4nVaC1vRMcVKBIGwhcDxZ30RBEgp+nlG5FK
zJ34vIH2VOBwLU/rAkOxvhIRMro7pH40R19qeB6JJ/uUxkXNF6M+l67Rd20UpYqfjpObTNyD5vET
xkugyVdxvwSSwXSA1ahE3CEf1GB/MG5roM6vwd5I7goFB/ZfI9hawX6Otqw5+W6JlddH9WdxX6qv
ZJy0f7JdIfe7tGW0/R2kKiHjn5zi0/6asTH//lBZYNMKH+MykUdlXRe43Ve86L1VZE0QjoBgNnlK
fw6rgSpT1revi7cwGzDnuB5NEWQkLD/aCnL/GEJb76H/NB5ZpL8ly5EyVBaY40G99dfVcGpxN/qE
Tk4z5P8Udq9NnoJp4JklqOjnnSZ9MePCVm+LkYaImKlt/kLrti13bhpl9pP1WBuLIBxEoORPF3cm
srFjCdkOo6PUDSrirlJac7o+01nhjRkmOyuOWEoGlWvSjkv05xh0gJefYuFTdAYSd5Badj0H+e3K
TVI4H0uYftpfEMPtqRE6N2Jm8w7XJTy+Y8KJU99KQC+Q5LstOqWkl0JZWA0ya/cAhOjQkg9m4BDl
JSnAst2v5jzvUxm6vJeeyo+YlMBJgY3r2pnNLcmwtTEzyqZ4WaR3k5tSjVXcR9nprGczjsAm8itw
nNTX1NymJhv/ZT0ftWUUybbRX3w/kOGjD7DzLFRrlGZ0QF5aEMynaFTLSB8Ro0AF44xullgUiKL7
Q6G3PNOAZ6xN5Gn5H/0Ub4pewPvr2Bic0boydnQm6H9+PItu6nuvWMd/Aa5q9/LpRAXPD0dF8Jl8
OJYwe9RrMO5Vrtxt6H/NHLnJ/4k5XUUJthMIqpCfndz0SdKsCCje0w/bLtXEUnDhq1Nmy9l4AuNL
/D2NG8OcOppDNkUtJQ/V8+gyvTgxJtng0M/IWmgt362IkQn4d4uv8SOMT5y8CDdmrrer3Wo3GhmV
8cMy7gi0WXMv6tfPnS/0koK18O8ScTHo8IfgOgtWSX4EIWUm2bwj99shxO4v2w/P1nLCUVx7UEVd
xwcP2LiPrNcks9zBmQG5UxQDoshzmbJf/jfhtENbKy/u4wPzqydLHUdlyReow37bzuCqGX6BHvPD
akZx+Sa7Yu6dkBivPBUqeThSLVMm5SJ03o6ILi9P6n3onS4EZOgDAnV0gtJ1DYEEfaBxrr/295wc
dgAihtdxEs/jCFNdpAK5DSmGZk1RW1YNEsx861n4TX/mvs9CAERSvAoIlS1POberV6uEb+ixk4wN
BvjW1cJL8vR/IZL9ZqGYpH6HXkagIbXxEoekQP7PyhF2MJKZwmsTfmKKCwtJlXyKPPlsuWos3ees
eDTo4s8BEARkDpELf3UuOQkE+fh0DAePFE6dISY37GsNP4kATqLQvD7IYfZTK694U4rfCwum5694
GHhiENIPawgcvgYij8OnpVkKXpb9MkhjwjgWiwEQvxCD7eRbxth6dn/yqeZexf8IS/PzFb/09pNx
8D6E3VA5EuC3k/1aWLjUuU8YGdp5woJIMXMRMqIntICVQQdAl/ZYLBvtZO2tZnioj0EyGOGC2Eq5
66/T+t4XLcrUm2wzBGcc1Jj2q4Ilqg37m/v6iFnrpCCIq9n/GjeAGaPreQ+CtzUHR/Kao1aUyXgc
b/0pYd/dHj+kcaMZFwCBV9hGx7+9OFciGF+kPLMMSLps1arYWDq5HNYTq7hBPJybcnujsp+FphS1
zSRgHE14TLI1MbZntcAl31cVPN4lDQF7tyTY9DENeYP1UpnsUhowPhJhuFa7vaIXxTah8paFEF3g
LeBeaSCNxTeZeKsPA+iPgx0lcXcDjvaFlJ7UjmqZJi8yOyYrHK6AFwwbjXJ19Ag5fOg8MJBoPX9f
DMhKb367J+wFJjckhrwrcxs6yXXpP9jyHbcZOHBb9wUMM6qa6bW0ZBtHcC3k+4Zni01+y5VTRui5
ssOlsyzrE6OnalAoFz06LWWDQNR4goMPFJ2qtoRpXvl3FcsrQJKo31U8dx9f9P3mXisgKCoJ42vc
/svh5uAtyZiYfuqWvcNj3FY3vamxUhVpafgsmut6OYkcBhME36Mtxxok7vTi2DCZx9UDAmhwb64d
Zs1BdBrEkv8qJFggRUjZ0pe3XA8C0Ytc4XGpNrSO7tdW5cHNkbvOyMRwYYmsZtw7xbSM5y4zYlHc
kZ89ebYhblgnu1CkOjPaCbgE+GIC3PB/ACbbw6LneozF6CzeSoL0PGDeINg8kpBFk9H8uAU3vLbD
T86KNNjvuhFqGNlZaVJJgumM5UXlWBRkdY7GeFeTtN8mknYM/RgKXv5sIqlkhJmSiKqcSsejnXx6
be/4ns6zgAHJANH4jC5zbi4P333Bfx+NP7gXgh5MyvCOq0qUCVfnOoHxJl7LADu/dCrPx7KR5kEU
6aLa9TKvue9k2chQAFLghsgyeYCtGLp+rGXX/DL6JC5o/8elzMuZuN1/7r5tWZTK5KuijbQOueDt
8y1E2X26wysta5Gr/3J1saq1llse+oA7WHa05I1BVEq6US2tcFXxzPMht+yvVRx8egpaoKIHRsL6
K/Ovyf6jyAome7bg4Pnz/X1Bn7FzUkil4L7l2x7pZFMenLE3KVTFadLUCppz52hFfVccnRAgvCGk
n99/ogePz3JxUoe2ingSO8zJNTLa0YeVAUfjxNGjl5jlP23VlGTTEyvAbQfVZ4c9gbpXKz15kjex
bkfqWiGpMmhYQyTTHq1la9Y12jkfdYkcAHXqJIG3/tcn90uRa585bExo/Oi0CA+W7qVpXpieuRow
SBXAy7tdAhor47ZumQnQJOs0iftzy489xQGrFN15oCxwBw+eT2ZQtfm7+a5u7uqjFt6zdKVun3NB
Btd8w//ppm53kpnoMwDx8hTLb1QagijWhFnSAw4o7I7qXp8KFdTj+actFGf69ONxJtCqQuXekzHk
zJ2zeeAk3YU1yCDYug3YTPaVikYQGpFqLS6ZX9muV7Ilgzb0S53EHRZHgvXdRpeP7+KmFMDWw5Be
c83bT8QWmxP01tLxXNz0PJnLrBG0IEZ4SOyc1dvf/Vmgdu027mGrOovUG8CRkMg96bv/LEswxJLI
7NfoCCVZyowJpgnahpDi8PoXTNUiCtXThoINALOgISDm0X57hLzjlpUTKj1X5KTFch8iEdfcWA09
lNhc6xg9A7JX+k22vyteNktr7dKFpFeteZAgk6AbJq0OxuO0Zg7IqFYv9F0b22eoda8KksgZZQ5R
o5LIRKvc24U/0LnCUd1TFDt3BHV5eTcbsFT+0ILEes3NXOeO1+NaRKBTG83u5dv11UmqiGHtKXCa
oK/Xo8l2v5mOSPd5eKwG99Fs0UJOCbbIwc82OZyisockKH/lcdFGhWR+gvdEbvFyJpNA1BJPBPjx
VbaKFfCXpBNvKWqGA48f8Jg6l90dPViTyXhnAuuXo3S+8x04gJvHQ+kUChWZYc948jiG1fSIMFuC
FNTP6YyAtRJvcGJvBukSVmBmxvmhvtliv6oGZDI9s2XMrAAwryjcXwx+5OSDykumMxX9DAoNyPVI
0RiUB3XFBQKl9rhn9mfjmT8I1MBK+wTdotxbHsu4A05XbvyDiqat2YWKbctIycx/TMQGHUE2BDpG
72+1dthdbJNFI+RbZ63+FtnOL9E7DiqS0TxoBtF1AiE+FlseBbuapNWGOGlBU4JWvoIdElgQSEyi
4VGzVRZ6ivdCqc9AifjgBiX0NuDcAPIe3zquXTkyKvRmWwfsMlmAkXP1N7MUMzYujmRVacEnx0Cz
BCXjM31B/PZTe9YnFS9bboP7BVXSN+9iHFDTE2DKURzX5BeqYeh/aTG8rNlFgmaqGaZ23LmvI/Kn
drTBRkiKtkvRXEEaXtTD07uKDwLZ2ApTZsGrhzv5N5FY3L0CAO/pXcpqZ0LASKvOQoP8dX4FMk7d
HOZKETxMGRVCQOC42BXgwNpCz6tH4mT2gR3tGYhysrqFbbm+t/lJLC9BRtH2pb41kMnKBfTiJ9Gs
idI5YTDhnTWffioFOSl00Kyw22kfk9bKRSzmUyKKx8pKbNkiianzcI90stFcxKeQSG3z1Ncit8RB
oXxVd7e1YFpnYG658Xk/X5dqmjKNzPkHS242/P633Sp3GVb3ka4cC+t0k+IHF3H9mFODHl3WBFJW
iEpFmThbuSN3VAVJg6MV6ZYcKBbO4d0hUSQIqfwilhLqMXahPRxjUOvyUurSa5nqrF3CpgCTVzV9
sQ447/gfs9iAFolXyACsiTgqx3G/QfSwMOXlASjXuq5fB+Yfuau3e54sliSMLaUw73TCS5pdt7zi
fxDcQLHg/5JkAlNHti1XvhgQ7U+27IBXGCXh+ims0fMZc25KW2t9vD47kj6+WsffkbhzT5KwoefF
+gLUqdT7Y5Kgv7a96OF7cncRLz8u2fnt5LHsPz8eqQGEI+Fc7Oqhip6phPbi8YKfL/Ov4feRtNOe
NvyhltISQdAqrsrz18lgofql63wKNz71+xc1HND/IydiKff5i29WV4yWbrBDiOFxrmxMMy77QR3W
PUcRpP9pZTKaF8YjwQxrwMWKUYfzGTV93fJbYn3o56YO6ttTrTU6DmDD/q/p1+MyIFClgTV7yxuI
XQGiGHvQuW2GBGwRVm0q9QpTfWZMN4KO6+18H7WdKbLaQqYBce+ILvKWSRWBatR7hjyL9ADT0Q3/
IIylz0iY1OJoev6TTADRP2OGMPWet8SEvPWHPna7jOpBLlV/eAj/DwfDV1jUTloLAHV7qHF8G75f
aLsj44BDd0iQG6bxMQkGHs9MfF9lJl375h6CzVGMONkE4T4I7ZTu2eReUeh/X/uw8wQevmHr69fF
TPNaaDEWzSkepzTgh3MgnQbbm8WM7WSXyXNGLG04/sfe+rL44tCs+h7jAaD+vX2xw3NqcptJKSbl
fFtVJyFJoXMK8uNJ3yLEUgHkoHQT2bkxnjd2APIcUlSNfZYbbBxqwSUYdIgqrGDSICWL7yhwPGxZ
J3PC4YCXJDJFUJsXzwCB4qMakvRs8cP8bctRfcSv0ngXlQUulGR+Iheu5IGnzqMogRf1+s4M4EfS
2ddD158Wdg0PqyNqFyBqqICsD9KngHA4ZOOB3zYO2LajS2IKAHJhbufmocHFtuT+MKdtCYWTThP5
2RiirsEUcv95mgvCXIp/4nRa4dgv2zSW1Z3eYpezcq0Avf9Qq1LbCgPB0P0s2OWqtzztnEOkSgfs
aQ6CRwaHT8yP2mTjhPzgQ0+8Fcdj61mdZHkVob38LCzk/PD0+Tf6SKfZZrFjeKFw7EaSyrtIu+NK
6plyzd83+Xj8lwrRXVTfsz8WJIYY9p9KEPMbONs7FPmJUufkFVl/dFeXsAYkXf68U3WYJTS14VPL
ZsfSR6yW2g0g3PHEqVXOlz0qoU6lLpKP1MEvBa8cPA5F8Q0c/DNLHYTKEoiM9w4nyFuv1qorL1qH
ZpFpVmJ8vWUNTlAemSAovSHfgesnd1i43DzQlRGSHmEXpJpeFcITJFL0wu8y9K2X1E/k4o05eOqO
jncZgKkJVSvEpF88Jo0SUWXxrY5Zza7T/MaVdiL/vzdNmu9eafoJc2zopv7DFBGlJegADNT4o1N0
3TwcqmIknzAtdgutdXm7v38V+0vdQYzW2RRiGxz5ksBXVz6bczF+uteWoMCIFd51z40dDRoLWHFK
9f9CY9jK+uZu1ma8jQCBnI6F0MAVV0VY5goUlqHhCbZ3p3Ron3Bn/auVo+jTC+j3DtVu7a35Bm/a
ntfKbOJ3KGwC+TlIo7Nu8fZSNZ/JyJW983z0bfrfo/am6J4Sj7WEo4/Hb2sbUZPIPbtjVvo4JJ02
qoZEvtktgSg+r3qCbvYVzU5Pt6ByMEP2tGwz0DmCgauOHzBuw28XfLJr7l8T2JSQR86IBs9gRbkD
j21DGAB/6RfEZbFKdf1jF+Zn52Bv2MsQPtXzEhDK5LW5SZ1uigaOSy5AgTh8faNE+6BXtj6eybOG
fR6MdNyhhj7lxAJgm92XwYmoYU27skyeyYZSj7+q3Sn6yg1N0Xu9Vw+alGs/FsuClu/nJbTiBa2C
injvfkUuFjRDuHeq/Wyqydn37HfXt3ETSv1yhFjd0S6n/lCE9ZnTohdeUSt+5vM0T1O+iXOa+fXq
WXulvfVGhf4dTaTF05QJumbHyLilyo3Rkg3/vlLfHuSBzXq6x3ioYnjMr3iPCwW3erwNkIVb3kVq
AOBm8+II6HU+uR8ySpiGfhG6B3r0HXrMwl9ABEEy8kbMxH0tWw61G7hDS/ugJOYAoKIa6x0f7wF2
hldqNZ6xptJk6hmKJ0Z+P0jTTCiRGscmhG9tevh7EVf+srkzC1zwzwDaFdzhXvN+nFIY3kCyeTLX
gUclOpUFTflN+RXbp+s/TfSrvxR89p67wqWKVgfvT2w9GDomrlQ7z9bEeEUILfrr0bYYlhaouFzY
Xq/TJUh3Eadq9hXWx1IMIX1X/ZzlghVkEqxguPzRaU02i+zDe1SFChE9xB9n/sYtKFoeJnhV+Fbl
6Fhf92/VFcNdm2eAVyydpR7Ohj1IJYj33wDnTNnevSVJml7kJ12J+IFYKXO9dTv2mZjhzFrXDXcJ
WwBmmUaelrq8pi97XiA2ulGlCDY+W4sn63LgRUOr0gcjiQM052UKRemlr1JrexvOIktCiSd9g/s7
c/HStnOFU5CUPXtiBBBVwZLT2/laZKUyvEPK8ZSZk7MAgXiHx57C6yvsfoQBXcQkmQHt15mbvrvr
Vo5i8MaMqn8+GFIBhCHTeNd49fi+HFbhjgAvM5qd04zTt+P1nLv6G3fbKupRU4HYWdWjykn10Iop
sg5YjQm4jQ9pWRfBBG3q/O+upalE5oeuoo8rUMmiQgQ5kYsQwkqeylurLOz3qAB2CyHUJorNU1/4
Ag98yCkKF9v6Vk2hDMGeirwNCFWxVK8OrCe1lEFZ8Ae96rojbA0SPvpuBXh8sRo6SQHyYON8SGwh
w1JY3PIyLCtj4kW4mRf5abiedqrzny+cA4QBfGvQerl64G/h0r/NrFCjA+oLh8jOYJ7/WNvSUH80
jJCMPkTYDtppAJPllzg+QLLViVuevBQFRb05Y8bxGnIb278qszKluNoTVxHQP1sawNfzdbkJBcrB
/BykanbzWKJFBtDM0eDaEflur8nwPJwD+D3ghxMeNqkSfuzIIGw8rKM7whFK8LLkTwvo0eIL5/4E
ZcIxTzA8MPWXgiKf1vpA0JYJgqJtLOBHDpfrABHSN2UD6dvayFhOpVgXuthvyJtQfulEMcPmUMiA
hZCDMJdHKC+Kvz3ZFToQh1tROED5BM3cGVrUziDwpIS9IP+owQ8vDNaQasMRnhlEhxMCLuz3NpWx
lhE1n106iNedKjHr/9SnXKzLKVrC0yxQhuMhPRMa9ICxz1ssjg2MmzYG/MdxWWQRg+a/GvP050XX
kUcqWqZTI0ryU1pOYlUT36hmuPPdP5+TbcUBzFKCUjOhP05QvifOye8aXxBaGdRGNwd3KCa3I9xy
JKHqjq2kl5hr+689l4sP45sDRTICaK8VKSQ7iHuKoO7rF2K56hHHQDRV3f+j8QwmueJXuOiazXPB
WqK/kL5LHwSrDv/f9+WFL2y16zItVNp1GUupeQLZPFoE/qWSpcKHKmX/ThI4G5UySQCYYG0YfMxu
jJA2vlQTzYEujOFijYJzdeuitLtZY71I2nBf+9J+x9eV+ipJQ9JfqjqU7raU7wVhQV12TumOcZmD
d5E5PmZ0I6jsD86kJ8TA/JXmWji1/m/wJWdoBIuwsHrZsC/sAsb8NL06cWy54r/jHHta11+rJWlO
QZWFJ6cc1bgTs+gw4NR+T6pgha60/C5eyN5laEyY/JFwW/MBzA6P1DdK924szwR7kjGN677SJ0lh
v7LI8LAbMGRrG4v6lLDHr4QNzqu4/yMncF9g1kRcOqkSpXJY5wZA1hofsw+Sj0t5XZjnSs2/xHBp
DThBJplDCWj0fyV65rjIPUTy9bqQn8TyEzhg3GerBJczfkyfdC8nr7FtyOCGq7ywpmS0QcA4rwlp
8pFialjgpsdca2yXIT5I0cYPtvDz0DG6xc3+kExGRxRNwfrQpk2/mKW7WH8fBLwFEMcCyZ/WSCHi
+10uTEkiKOJ8kgO834r6jmmxz9rtiWKQ0Qf9Xe1vAOPbPB1H1IWlpPbmzJlQJlZXkSFyqaUz6Wtr
7QFIB+EZZnbMJJF3+y7TWtGhWVYlCOogllXGgW49pzUY88v7VusAY2ZZaIK3ICvBt6NBJLTljwUe
lJOgLWkLJThTfE+LdLpbQOHaGTwMfhVxZtkCIgtBoi0z4DKVVwhp1t/731yaueg3gL4zOZ/rfbxb
gRwMS64ygB3OKHZqay49dTFwpGzOmAnkx9f1fBPIYA0c9DfwZsFHbJSXUF3tDvHiffe/QZMj7TPd
I1Ht6kFBfBM4kgI6e7JK16ZBLm3y+rUYpUsParEqzj0Pm1YCij3lfZxMkht5tTTXJ2n5Y8rJGXOw
zQcNOMV2jXyvO+3ke2YP8MgZ3Hu36sQxHzUqyq5M4ivrQcstihOsWFLxwyjThuwyNIh44VdfnyHr
BdZuqQtnK4GzqF/BneCKpIxhwD730UmkbtyU1E/7+pba14DOxJhIT0/t425WKT32gQT8Q4bhF8dP
L9piZA0PDlPLwSWSlc1uGTxnUBpu8IbO7suS87vHNhuts2yxug+ENZdsQwTni4sY94ELHNXgMStK
kiZ/tXW4p3vhwcPWP+DFM1xsy06PKpnAHniMQDDGZ4DJU1S95BMQ8vMSLfb1Y2QUOg+ibD0aQuzs
gntWYuU0mq41R/SCwvQDMUD4dQs+xwrrSN05/575/9Wof7BYn3py0gAOCAudEZHzlboRPThy+O9k
5Nd2b/yd3LXy49ekCOSp7S4X9IZv48UGmXlLjxQurPryPrdC452jAZptKAlaUGVjJp4G+c6Vl+8P
kosQrO0MPp6VmGFYl36ldSHvbjxsxYHJBtIVUBCghiPkgSPmkizHzC9vIF5odEJiR2hIRQ6FH7CM
0+PPyeSHs5GRgPTJJHzN4X1LsNLC/k84+O9wFRnDtOSP1Y8RIFH/dfd3KMl0ZDB0AhYwMl7apUuT
15WF2Bnl1pMXaBAtYP3GY4jtzhmy+nuXbxqqmq7Kp/f75RMcZ2BQHxRXfAkWzN/9VvsHvfYnkmNg
7On/TseMgpnoLK9yVhR+X4msON5gYITdnlh6dpwgilnGHi92I30Jv7cy5iUwkFHt05uC4i/r4wCW
QjnI87qQLLKC5T+KyDdZRYv3FRXvu2Qezz2CTVy0YhS8B2MUzZaF9hSoIbeXM/xoTjLA1mDg6qBF
zMbq29e8i2gBnKrMitpOAl4JMn4vSGwib+HHvlPV5rBccfC7fpf9ilOkIT6tgxgeMH+Gco+W2Rz2
HQMxJ40kPJ6APD9CzzbS7EAk+1llpEIkYzDgUVnclwqAbijOejsyHoCpNQA32V6R+Blj38U//c8U
Cr8m1Z9NFgtydmYeVMGY4VfPMkbHlY+7q1DcprP9P7NQshsU0k6zmLxfCruyNWNAMinMDBPTq+oP
T+ggOzwdnBJD4yIGpOWZaXSrSFMyVSeapJhgkYyI+i4YvIIXuwuep+I2rNtCA92bV9VD3T5//+Hd
B+iTsNXWRW9+GDbSEMW3422/R796cySYFR5nrehdCvz3BUDwfodq7XxzIBsg4e8xqUyL+ToLSylm
UbALPhI5MQpkX81uff8c+XvWFZnMCSnwai3VQh2msuyrazTPNWKqYkvUv6K53OFL9kyxNGY+elNd
jp6h1fqVndV2IrVa3CfXSopGqr/NoF3daXRbvBwnUokLS+A+ykTfBxuAc5mGpj8gc7/HjfN7TX+4
1cH4gwjcoJ/OSWTPKdVAOvZ8w3XiGucMD6S6SRKk4oD/BEU9cUrH3F0+St7Bn9cx9/NiptcLsv/H
i0gY7nMRNYO7QHSs2fQgd305Wk40SeeiG5IBvaiMjs/vuzxvOFC2OjhhXVRZMF6zMMMqX3fqssfZ
ZnedUZUv9q629GzMZ1GlBjv2UbOHeJriSZHzD7DC9yXt55fH5FZwiUZblpDEgkfAg7KhagMBPUX3
YfGYOFi6DWp5rmDcef92ZxjbGZ2dV7EmAY4muzAfN8F8mhoSUWYjA+DPVD6zBxA9xF/CmNg6Xzcj
/tdllJg3LR6X8FWc+rDGTORv1bNWUm+HzQAW3vgKWSBoME40pvsYK8BQixcBjs6fruMQOCeS5R0b
98aS/tD6x1jd9MnFlicp8AajXyQtVQ/sF/gxXeVorOsYmM5tVoGGtLnAef+YtRhgGGAjFQeSWlpX
yEOk5ra5nbDH6TuqkzK68Gdq+D/yhzdT+mjAUtaX4QskzV3cB0TOOdCMZldUwpknrt+7J8bv0J66
bi0zuaoXEnALOSRQT1cyzmnaMRkmzd4KwxUcv46niDTJD+PyklvNRtxst71K6hzEfFevhpVMMjC5
RNz0cKzYnia4PWA8/3MRUA0VK5x9yCWVMfWzRVsiT/gPZJGnrSh/7GY7CJuc3nFVBpXxpzr8iUkn
1U8h0luDGtqNIMWYVDH0gx3gAqLfklpYPwSVwAoc/Q54uPTtZ82OXSQLVguuXwTlUEnAEniun4Iz
BN9E3uKcGQrS4D4gxlcInztogu/eSPVjzVLO2L/mCA8Y5l0tEO6O+81LjLCU932e/d44jMyKHseM
9s1huM1kDzRoJaIHnnqmPGtZI/9yfu8ZzUTaiI6WhhIfROMrwGfU93uXpx0iUEPoV2PQLL2JKxi2
T1eKkpOdAGe+Q3SKQQuGsdo682jUq9Rn17jNYnUGf7ziFvwsAnih+QAIh9+8encC9r9bdUsmgX4Q
qGtkMPUxeTraE0rXnYpueNJyPtpAzhWVLNid+a/WX486gEF8QawCL9/kLqON/6VHTvSjd7PXhife
oHJ0QF4+UEG1eS69mUSdKS9pdiZuRe6ievKHLvMDRqYkEYlhN8jSW5gDEQ/LWXOIqnDIuAScHyIa
880SOleAGBV01y207e45jPwZeTKWiTi9Lj1HEYw3BlmP+XnVUvnybW30n2ipQSHBleuC1PqmbdsF
cKOPcins1sU6ie3KKaCY/ByLjxE/5ZO+Om0Jsr6jQha7P1phNeP+ZY2ZT1Nt7tHGn3h/bQ+8qAYI
iaTwGqrcKxoTB17kOT1LGMJ0YFltP0AIOXLi4bEi8iCJ79hNE6Ji3aWS1YNtzKkDm9ntD5RtPPnZ
qgXogPlNzse5qvSehVVPX+JOjKOOfmSQxHDYcmeSVrjRMCQJuBqIs8s8NeF08PZ1EnOd+Y7Vd6qs
tjX70qdnJHy2T5KBnKSuaAJMZX6EDBTgJIPFAXS+qkZjYSsab7F3V7bn1j/C1VxV4r/JmLUxVGS3
zoZVZLNvkqMn4AsEH3vuTnxr9jwjSkC526uauGnW0qHouEiLvbrh9agBM4EnEwUBkdvDN4d6TEKC
ObVuNBSyYnDkg2CxKPT/juPOY5/pFclXppeiQBkfccc6HGXVK5DPyPs2+X+yqHXGwDNkAQRlZyRe
BqrJFF9gnHPQtuMN4DabUKAaI8MhpnRymvW34Oza/j87DfEkBEfdDl5gJkXTamjbX/KYXTmUWtPU
tz3/YgocPf8JEzetoXb2O6YmmOdc8D7EYo12Mux5F/Zcgaja5IxBbMi8aQtWPipTPkSzpJDbceQq
hWk+XWJYoKtnhWzm8By/vOjamBxwxstUkAWwADsy2ALo/g7jBA6E7XDdmweRmRcR4XH1DULXarVK
PwJHpG70vlxmcb/mDBO6caCUxICDggNkSRK13T3yOCo+wCOdtha4SuUrco39qPjbZRt4W+QtykGc
T8/ky2b/nBxfnl6dem6fydwdUw4M061dtELOOwKMuVjpKAkMksRQ4kafL53MXmun2Api714A/0pI
0ImaGAkO38WDACS8iCioStvorTlgHCwkAQfYJmS4Nh/gpWDhn/MOxBvLNG4qx+x8Ys3A5h3IxtgZ
2ZxsBP39nOfjZ/lNqMR+TDQA0Rie1aKAdxr07x2/1oNUxwe/9xw4yMn7V4zC7qk6xZbEsHZuXcB6
/LjUjjTxUSuaViK97yEcFjPLlOJLy3iqh3+UlabPqPgZnTkqiVWVfFDtGjVFHheLqxkYU483NX8o
HLtCdWqcOjGRsXX/JN8Eu2OVVRuwnAqdQBADS1XFjrLprcugKI6n8EcVjGQhpUaCS0Iu+0rTRyda
WwVjpuH7bFkD15B/XR6BfD8RHG+9uuamOXlP39gtAdHR+PUD6AqDnDD7xX9mlq2K37cv//m/qFrL
j6YtjVDZMgPXhexLetK6rWRxRU3xjBWrgKayOJ8rhxvaIh5NwUAHXIyJYJy2E/9vlkHqTdTsOtoo
16a/1uFLZl7ZM3I8q63HEaJIQL9rLKdafEd9scVys/+ExVmro+JCdUxYrwAZQE3nii9tNRr7o9hK
QS+iqHO6XVqq8KNJnVz3pr7vAsnmsNMGOT25j0B7JmrPPiOccs0WoYyhzsGXEftXRNl6q6WtyPjN
VZeaArnv7Uu6ppNXvZHcPLMVe3lghbmg1lapk0uuIy2NuHXnOS6eKeDqmmuGMQKV4It6j5QxUdjB
v4DQzx4HPi0GsH8lRaDNbC1VQyNkzRiNwvMsehZUbXJDBYNK4OW0muAN85VTq52r9ROorN1U9S75
gId5zAposQ33wYDqqzrkK/U2aUdddgFqcPKT5Z7MJPADo/6LEFNtV+d+oMNUa9txvUXTtHl25g5C
8OuIIiYUgrMcluh3ytA9RUVYS5hhKYBBt30sz7beM+rPCD7yuU/cpkrsOeD7apCaBEa5AQqSOBuj
uqyMo03opdhXbTaxLXAwqGWJIy3+Ot20mVoHEEy/iZAvKspp2FBEBhEyPDXvuG3YIGA9IJWq1fQD
FdbDPL1HFtQruq+pmb1zzN1SguHjkCZZWi2iudjD3A8PrlKW1EZ3x24bBvBDGtcoK9GsMIrTvDzv
vAqVaJ+H4XfOhiJHvMjLTmAYT7awwd+xSS/n3geOZxce/oLAD1rriqjB+TIDfNe65mzbiaC1O7JX
3L/tV8PsG8omOn5I3Iny7PKRmPUA01uLCwrRH+uWJ99JZRgWzBAhCHotAfBe3hhpSvbjqdVl87ud
IYF8lJywGt7i86ehoQ0/MNtRxTNYB+y5lHAp0Lw/bZtq7BeY8DLnyAUBYV97bTVxopGs5StxiWH8
9TJ4jp/ecnWGxSTtDfQKcrnPBdbQ8HXPS4erFPl2ev00Hagw48TBBwEtnDQJgEQiopm8wDd/KDeY
pGTbOM2F6/S2lL8aFHhiHpStWMr+jePb0pBOP7nzf1nOq4ulOVzpy1ofTqILBndxuO/8EazLAVT9
qelVmzifNCEIFAltcY/ipcmq/2up/MusEO99UBaXz/6WCE4sazW1OOSE1olhyhLgAqSvcl+MqNg6
6w3kiQZqlq29u6Hk77gRTkNha1b1KfACt2JIlXK8+tf+qXHVFKVTKzsN7C9uzY4ZILxaVynHZYQI
hw/icfaRFcnR+8FC/8CQwPU66XuvGs8I1qh/H9zooskclRhlKqITi1vvh5C1mqKbKJeggkIw3UKg
q6IiUgTIXHedVvvDHRR2flwELaGbx65Lp32gGX0gQJ95sUaECo50bR3tPv8ZmY9PPbHGrCoeV2cv
yy5HvRzx2sp46un2Y3bn6xClREZ9ThaqG5EGW4QhfKfuG8MT5ZyDJ2cGcVmtCbQRe9DHMrYB2/h7
tspVyNww5wnwRK+vFiA0FW6pERAqMHsXy+Jt/WGGOVABBDDMrfMaRIwI2wJnIihgwvZtVJkZw1tS
0ZycuY970rtjRJ5dOK3ldoRzawaU8kbLIQgX3tH+aFVom4+E7YtpLVwthlL9unGkiFUU4GwBOQc9
PXz+JRITLJVE9N5mHxUa0q6ISH45wIOKDIiK7j1qAonRIxi3BCRa447HW1RqlQoSJMJMyxqTwnr0
uVz2BORzj8Lc6+NfvpFBYn9AB91+MjVlCfExunqvqwJ5261TAvx9ltlQpU79ZOcXjY5M3VvG/D72
3DVg1ER6AioJqAtts1trh+mrVUiitNjHfZpKZIh2N8SrZ5T64T6t8aYv9OM6wOaGFpUeuVTu/vJy
g76Y3APTHNeEhHc/MIfcXL7bkGJPGxfvipD5iaBI0ibmOsnpRHahTCvDCIBuRgEddi2IimOLG68s
hXPwjxPCdX2WClid+5wlWRBB14s6tLQC9qvELUXiFQQ3NspUpj/8aJIH933luuhuWlZb3GLS0Ixk
Ex75uTN6uOtY4o5i/3x4+zDd0wwuSOU0BK6ELi7HIr3vRSc1Ub8tDHpBreHSQ2Ehymh/bvOZFlaT
45gkEWHrFtMipcZLMzfDl27bBV/kgJT2KqLFDqxUm5wIE0ca18o951v8id3zP66kOfEGwVXoAIG2
3vOGGNp6W669tUVPOZ6nedZhBPh8mRq6UZUqPmH0RvcQ1IzUkrAOqfh1dCJMu9lK8L5GO0/aeQkV
NPeDXUdLzedLZCYDkIo9EAZ4ZekkOx/fooHFcCd3EkQtUW4jZhi9V6MplRMEc1EtW9ZRjZJY0SRK
+BKbpTyXXUt7JYqPp0JuC/VeTLWFu8ISB/V1csPlcQjNWK2CwFuawoWLjkSVKpT+pCIreUOlbtck
9GEFuqNTj/RbJk/PL/tbLnZLmeGkGczQZ9gcKEKGRMNd34wjD3pmIMRXo1OVxBwS/Law/MojzBqS
AYJbba4DmtBm8zKQyGvdGgUozfBipQ9UjlsySHwnSds7kei3e9oKzhA6sy1u6mCuKcKQT+MyvOsw
tgIcnSKwXe3iZSn17xMANuB+yUbZ/HZqee/Gq7AcOPGq+oHVKO97jR1ZvUnixzGRPk+CiNTNwvwV
JhTl3SZmqwSpr0nMClvJa2dDjMlqVru0Ivf/Rzc+nef2tLxXoLCxZeEI3mYuuyf3/WkHYnwYczZf
nuiShZ6K/4NKWiEl5GiTRSqZrP0U4do1mZ/nsIMkdx8d518d1HWmmh5yQNoSHlcuy87tKmpL05KI
W1AVlpjws6caPV2WJIxTxWB62wk1xGSKI7t+MN7R772E0R7BElJ4aI6dA+mbeKKGQ0FZrsEFOy8j
DvYvVP4Yi42zfk5MgnQ+lycoW/hj2hXSERKYX6xe7sFt3YM5QZN4+gJB2KhIyTGyh30fy+zEbaVF
EJO9yp20My/BKTWWXw9qB2NRHa3rxnwhWBUZwsSjPdEnNmUGIJ5PEogKE5X8FyfRGEgFtsklZD/I
Lfye64NsuP9CgGtIVUX21iPwjVTp6sGGWt/U1czkJNZa444yhhuhxnclbWmo0jrjG4rQq/OYF9WZ
aOQTjVreK4koY+dCCxcwfLoHTthn+N+Cc7t9LtshPFMM3yg1btcDxCWtL1XijdJ3+5P4qYXSUnGN
65vI4N7c4MlUe3+sD/RKEM6gSuEyzoP6KGFqIjMSimV4jdyw61yutr6aXM+Js268PbHAMJmfzo+2
ih1P8oi/WIdEqy4sJHoFM4S2XbtBfXV6lJBCJEy/O+vYAHvae1zYlA95J2p0mvVuJiWf6A7Dx6XS
C+aKv7fw3bFfzGdLqnX4u689mdGjw4aiQS0zrrOS+gpmMhY9bmWAjfdNeYjYaQbKx1G+jXHbO9Ky
OqeG61/jqq/Pwa+tz1mXpiAYUAfzvdFyneA3YMqPXyz4rBHvpR39q1pVR104sbkFEQEd2/fUEv3r
2j84ult+zmr9xftX85mgxvVWojI/j+pSipZJty7oPq9KOmEBdk9j5MzkohF/xqLKpA0pa5xRwXDw
H6+5R2LO+x9aETzkZ8bkU+tk1J44kGaqGYlCBt606dMH89x5Bl9RIpwWDfA0Hq6D1IlWkWwUFarA
C0rMYyRmGHJJwWtWMkbv+c6rimLqE3zW1pyh3v71XbPFSn/W4+Ppddwqt+h44h8HdZm5uh/WS40Q
Pdc3heufRSU5p6dtMc3g9F3nhY1oFa0YX8U4GFfw7TCY8lNXq792GDMgCIABYa51TuSTMDmv6umf
SHdi/VeByTK9sfkXGh0jeLitSbTacpPS70F70zjZ3OXj/jaXAFoIs0x6LB7Vzn/VHA39xEqcMmh7
KQQWigmeh7VWTErRr9WVgC+IEeFQJbiVlIXMv2ad6UCCh5XS4HqZdzU3F7JWdjPTlj8jqzcRF2Fp
NFQb7s72fMO2Hn0V73GwFAyANWnzvIFxAiLiGHq4AuEBHTGSv+TMaSu2C/eqJeUi1vi5RjTVlWhP
KZv5g3bZTYEh5H6HBLQxqMkQ7rUC/NffQFAaBkVmhgiIHrO6SrPg1j1KEOWOyly7+gC0QoHT0yjE
uyLKIzPTF5neRZdu6N5lIRrC1wMMv9qqqcUiRtZ8odCSTm6tvfm6Tb/gMBOyc+eAtbqXV5xxTVa9
w7RUxIohOhO2bfPXCimkwB5fdLbEJHkfVvaD+7gEXAuP9GLAvBLyqWLjYe8/TSnUp1un+HjB6RgB
QB9SqbDlVumKhQbGn1jK0V1mbYowsNOVYzbJ4MPXOpG/kWNiXdBfuEz9ZUPvr6TmhF+bFBdATMPe
ZfJ0gdC+jJV7gYMxVcLP0m7k/JHOUEwQWFvQTVZq/iGGz3y87MmziDdPOAJKu/pZ10jJgyW4Inj/
CnHAxPTDz603mo5MT+BzNdu1veTzEhsfyRWYByoNe5RabSD8KGdcqJmTF5tQWWB47UD86WuOy6DR
hb2XQY97puGx7XyBbLgMUbGUdzeoV1lD3IbWUjksE6Ncc60c4oUo6KOaNcQtqCbHKHYLmuAEHZwh
UeY9IlC/4CwODtC5/JVOHenujUeXghXFyTClY+r428lP3aYrDR/C8L5bG6+9xihTfB6bZesDRehQ
rjEe0sl3E+x/ZQGUACxMJw/r9geKRD3Qo5DhV9fcs38RFuNYlvje3p0d1+CocvIbWQWEO1gQH/s3
3y4p5u+wmik2uu9Lw4hNO/A6UMNRgjNfmHSOK5AV/9rebTCBGHYWUqDXEUtnMrUOp/E4dotiErrT
ENBpIr7rIBDgWaBy53DIXMo2Y7ylWIfxL2DhafUgz3ijFPVEsrdX4r8Nx/t1L12tjH3poXGZwqXx
PeBu4NPD+0Va8+MaCFoCE6VyhIfssPv78B3mMYtQ1wqknRAdGbQlvmDtxBGAZRo7JD3KTfLtpOsz
wiIYpSVu3CJWRQ4ukZ7sLDodwXbHmPaM0ZdnIirMz3z8xQ83AwEtPRPPHgrnNRgDsxQBs6uApPel
/ldPEURbD7vf5yp0U2stTwG/VE8+NsOhZVtvD4CxaCbdyyZ7e9K11GrbRAelHNAEWSixPC6+LsT+
/7KUIioCatW/lzuEzUOWL5hJYHlmHVk8xQ8d1ObSm0oqnY0mMeEEzIh4F6Umn+VgZVL0voE1L6Ry
8N0zh9dE7/skcXHWmIxxh4iNm9X5zQB1BjuanypL9dzA+NBjP/xPo0plhcFX1pA8gRSBwVC4KpoR
9rUTDsxIBmauevfOKtju8LXa9cm/QwDcaBEutwQTZrncFQBay+uB3qKAd/BkD9pG7y7jYSeEB4GN
wyV4GPY1GoE3JhArCZykFwNxGSHsOyCTpkNSZ1NOzipbO8pUOz1T96IUlX2mLuCBOxTlDe+rpLOx
LEhk9lILhKUtf0tcBdw6HbnIayxEeihrj1qhBBWLpxW0EETKHOMmiUb7ZSbLBi13BGZh+HP3kDOe
DEDGkAoPyFxdZcrs+P+cTzby4fcKLrnwMHThfFlajTDUBkYIk0xq4FZPk6kq9AoVPoG/PT//992Q
q6O2V8poVT6SKJ0338RUMNXKaw6W5yzWNcR6/uGaqIZgpoUHTRiA1vaFUI1bXnWaeojC3jj6FoWS
y8Yo9Jaaiwu/fH+HzYPtIBezkGOb9NRi+Ae8rrLHxBhs1kRVOlJTAHEeNQCvhoUy49XVw0NhlALh
Tq8T7wFL7Oht+fVcEpCmdzYmJkkNyDsRxcExrfhMky1TUleDFD8rmm19kWZg8M978m1lnOb+Chpq
Mb2TjrtjDUICFGhWqJJG2ehuMiHRi3yIc/T+dSHFSYjLTNb1fbGa1fc7v2WZk0aS9tI5HegjUv8W
GSbgE3hspZ2kIlFLVmEg2dneuzmvwj398xOzc9pIO1JAS0b+v+ngB0lLG7KxUUkdpI56zGn155QY
Dr5L7Rq/HyK1g5/cJOatw6UFJUR9nNR75r66LfLZwPF1c9oWOEW1G8UdL0HzSIdGggIHtnGFchA8
CLw+AWCHB3BmNpdPmF2VfLim0EMIs37WCrwRHGzqxxG866r+0z5qZG6YLGG/hb+FMzh3IZMsvIT5
WRtH3s/ADUl3gTb8eF8TIoy4Z9tPbb8wwX2xqIaKQNfg2ojfcNSFNoW4ToRg4uyV5X+EpQD4WRGH
8X/o6Ihknvl0Uhhin1U7p8x+0ekogo6eDxOG5UqTrgQdZi8OivxOYwvwHHrYAh/d84vEaz9Z0I7y
nB++vCuwWDrvylQ9LyCI4SutovWw6IRO2lXZJuSr5vSoTWdwyCo8WtWFnpUzuHhnIf+0aB70UTb4
tRGxJGkE2b2fxwjP14dVf++2i70rQ66rsufJbQqCCqi4OjAiSBw07azMSSfqdyr/sUYLK9qoRtVQ
yFi7NP5HUoKHdW9Sum3R57OkB0y3XyanwruaZI2I48aL0x0ImxOn9gC7ldHaV63/NVuyS5hzQZ8P
1fkHor8QkwfG7y4x8KBgBfiRZH9cYJuz2KLSNy4cPkiK7ZjlUla8G2edQy5gNW0y4qgf47fElyLG
QyLAoDeWy9FM4klZWEsb+i6qDPj3maNq1CGsoCnfySrvJXvAXuHk9e56LN1/TPZy+4ebHoJK6/o8
K2hSsFTY6xkEtbYbji/aRgxlMthT2HbA278ojj8PCjqFtjSunxfR8AY6NyaW+jQgtfxoouUNc5bY
fPu4VNdTtbP9WsptjMnYpEftEbSgE1g8kg8hdKNFa/q0gOmIyq1u8WkPzMIo08OiAHRb2fvVzFV0
5+jfATG2jKOD0dN7u4V3JWESYuLgdy9aXU2akpLkWE4VWw+rAr+DNj3opoF/rm8sabtfG20vVJOg
xK0+Z2LxiwPvg2j2VXFfcxNKFIHOSE6CZxMKlXV5xg6Jil1tCYb3QjoQk2yrIh6HUtie9MVepg5P
rwdnz8D9Uv9Vf71Sro9De6o+IM6R761EFmZ1WC7O+PO3S4du8SfQBj+vNd5ZZ8JrWtvrWvxA26Fk
JVBOp7QMNjoXboz8woFRw2ANMJPbFObjKp4Z7SQiDDcfgHitIwpV7YtYkjDd7ZX99FpA0jcheDAc
fWEvMmxtaXkasKl2IpfOhEy+kMRajV6rx6Og67DjH5N5S48KOCe0BJz0AlBjNMgIZnX8xnaBEI1V
CYuWlAArbgWonMaG4N+sxqzgRJFMyCoj6HfwhJp9pkftuc5IHSBRhyRvJovW82Tq6dmxSvGlI2Ej
elLWalaXSlXZTxYCTXcIkBOyeo3xmppGXyUX9PypQngjmm++G0IskO+gLThQTLOCF3ArqtgsoDVi
/vJ9F3ICOq6NyJucfndvc1fF9fcwQg2IwoH91NQ+BrHOXM/XXPL5wWnXzX8wLLn8sGzlJkS5Ops2
KdKwFLb/vahzIHguaWPi05+uyjIR1bO61+DIlmrLfmAjDoOrj8DRbIJ2IORGw/60ozJiLOjvtTa+
bd1CfvvuSYMClyB8UMCLagdBMWkbt+/hlm4qY9ciFlEpe4zykLUb4fCWlzg/kJaBy1Bl9jvwGK11
34ZCH39tme7QlCS4/m5WxEbUJnN7KHu+T3V+5pGkURYxc38qjhTwdfN6UvUyYe5LggOUMTg0S8gH
YYhP772qQidAnTT7aC+bvcbyTtz/6x6wziEuZgIDMv1NiSgnDwHHPNx6jMOUVlbWJu2PGuEWI6/K
jEM+s6xw7q/CcFKJsZHfNEfV5DPd8HtgOgMGGvsqhERYqflRDvemZy/OaJqzXgWL48vspLKwnQFW
57G0RwFRDuWkhjNpcUmX8H0aIPCh8X8Hm90o9DA4FMVQdmL6+FQZibUqX6BBs+O0ipkGqnT/o8CF
09Usw5s46Gtgrof9c7vz6yzmDbJiHDDdtGPHRUeYldR2Npzid8JhedaFJi3A3TsRBP90IZyeDjly
KndKWnppvh8oIMOhQSFOm/jIyqDFiGDgN5UhSfkv8w9CUFFWVfgKNSGwWUQRv7qgZQFUERrPQMpv
/Z5g/lOatTeHzMTOuiEXBcBXjHFFYwxk/Mr68FuXCSh0rnD1S6Ftumz9CJj0rkYUeuQ8BuU8M23x
SBUbDmyyg2D3j8iBRp/Rztv3l7WG71iXATGNyTRolm2KUspYA+R2H94VkM1+0DYxngqa3d1aXrdS
kKvqixEfvU8QiBsTJ4TK46QgR6IsWAnRrfRV4OOGtfPXmszZMLKRmGYmpLd/1e5X/6PFxGDZG/lg
YJJR4/0Hs8ZOtIOTFeRxXKUKzJqzR6r+3BlRSSQWz9J0VCa9sr9TTNxm1pruuX0WRNj+MetJytnS
/qNh1c1QsRAsWHp6PwwsDvdxMHVzwjEh6DiAN7HsHH8gW9k9I8fwPkbm7wgb5TpDJX9FrHpmg11y
8jdWU7BKrD56Z0+D8Mm4tKkXQJ/JRCa6DUsyj4NtpOZhmCElUbUrkzKX4JCIOFtRYEKXp4SlAJAm
es0aK0ZRLWjvCBfNeZ6Nk8PLVpYXjWyeny//odh+lrOVMfYXAop9l58ul51aFhWzLZc66A4zYmXt
VRaGJYOi43wiTCRUqMBSKPI1XfvJqrxdo16AR8mNqbL9D0HxNqERsusN4nDkZJ/klLuU/8OCw5zI
yiwYmIHjla6GoMm00+mdAs0PSI4VUDl6x6P6BcIWVHX6JXl4h+V+CetuuWaPclx+pkmD41VUKsNB
5MM9x/PoShUlBA4TlK0SGh4B7PeCWujhlbjSLHZaG4NWGbOL0iZRMNAxoEoAvXYCpzJ+Wb6DSqK5
mmVQ0fx0lXq74aw4lMMeOCjfiuPtLiQApZXekAXkLF0+YHhRqrpRevqe6iEvWZogmYq9gLPO4bMr
mxTYhp6KLZiXANt96pwg0Sp9o066wIHwKAWeYDI9cyi2Ft0ZExIt6PM9xj0xtvZ6YYAM7xrh1T/P
qMwFk+HE009czE9QlSeupUtpmxhZ56Mv2o1GWkbLFvmEBZa4bn7QEsP049qLI5lnAcTLWjvryyxb
Wv/+pp1vVbdClbE/PakQ+7hkc3/tQ1qqox3HN2crT5aGTggN2CwZzakfpJZeFxwUD5Rjnj/6/jA6
r/7BDBXiTUEsias1sowrVVCFGQnpo6Ab4FyxkPeyfu25KJ6PCVsj5vasrx/Slf3uqCscLw9+oQaH
UE/zeyLInIn5Ai6gUl8Pol333mlehB3wgmZXZDbX+FLI2nha9+bqpe4NRF+dI4cIHx4gJL6OR/Fd
+EXORGFE5hu0OAtfbaIvN6zA6swkvmEfIzj4twWxBVLY4PxBi4R7wf/mCN675JLNNhfy0BTcDpUw
+/t6jmLe1rl1MQ4WHFMzw77FBoZWVdiaEdH8wq0S7YfPNbBollqQtE96bEFgB6Tb/Om8834O7Tp+
UPz4AaBOEmYQkUbrfWghO64y/WZiMQfxPjoD1vwuL+dG8W+hnTCkfERDbMols8dUT8ZAq0jils9N
XdTl+se6d2Z9Q7GnryCQMheE3KXjvwjVwZAF9y3UXwguuw8YylTPXh92Aeb+eHarct2Np8UnmyzD
9LgXia4xVpI2VnXFYEME1Ghjx9wa0h8rMsEX9jpuwYndXy3osTqThFvXBj2c2ZMCYz9OfcQFjEvE
zSS1FKD8unjppx7NgLo+ZZVUV2tZVPVGbF/UA4PLb5EHnmilWUUZk6PdZObLGTMryPUYN3tzxWBy
ba5WQL5LHM3m+h/67iAdc+/S+sTWNc3ltCqKxWJSBbt7BSgaPD0uSmULL6YHKB0NmJ5NyVZ624Dd
GnPonB0R4aqp6JfO71YeWfJoXwpYtzOPDVW9NBsuICafM8lTKhPPL8yTHnYWqWVYPBfq0Unu0v5z
Xb6x/0jEYHd+Py8d1TCOIOUjSOyEwNzBv97wJI5u0/HbqA9I8M9Z8+hpW7h0s8Mq3JVWMVYyMzKB
pkRPCMim/FU2hQsLQM2EZuKGXEhzYZXUK//z/buW6MuCkTeLdUN/2Sk1wJQfNxye7mEfQwiJKmjT
qlVCHZMcFgsRnYrnAdFpPUZBcpeMlFFiwQuZnCj3ApcsXZKAu2KAvGe3EvbQA6/3noe5l4Vi76Ds
HJi3OWe0kkz8LYFIh0LNNz66FvNLLcAIbvoM4eh22cEx2tWwu/64sBbStFCR4QzhLnqp5GCPHsuL
TK675iBwUnZYBmqH8na8B7Gk98BOc11qKrrKx55LnZc+sZMEZqD7NE9BXHX/JVyw5csqs8TiNVTk
k6oARuel5a6jbsdnGmNmnW3NDnYCX+cxYZ8pldyKIc5dlJKxZY8EQQ7qdp87sugWm6kPEYuHUd3R
S5DMP53mDGbcZohhWX3lPTGj9a7Sj3TiLg1oCzo35VfPD0K3YWAdLq92iwO+unsYPbfd0EqZqwN2
9E8SWRZgB3WyAVKvbPQJjc3MWm5zFM2+y4pX++JDUqrMjc2sP3AqxS+S07j8RqmuXY8leb6hRksw
SsGXSAgUA1uGX/pVnbSLrru0t4YAseqzcSmS2il2yC8YlENLyu1ToXOMyA5pth8lLr8MJaMW+gC3
2hkKWEGaRHUwMbUI94l9pa6Q1BhVkwmF/VzYFq8AQSfYmLcO9g/Zhz6ndHoUcomGLkvov0N5Tfek
yxjIgcFzWpNEth31F3fas9an0nz8ZPt4kQHEV/2w7WesQRzS2qSVnOS5E9osZkHxOx74FGcC0edL
voUO6HavCH7ylr2NZagxhaWteBH8K0ngt0pIbp94arLWalwPP3valTXY1jKIVPl7GdERgNhYrjj8
MaxH1X+4c//XxSiZ1F5o6tZbNl2C4eE7fG8Q6Cx+FJmPDywzx9ScIyU+w+rKWIobW6ZixDme6GqD
8oZT7Vks9juJfVOgKH8kfGFmg1b7RQcaKHhn2tgBVZ6Hqe94kv8KXpeCHb1JkoWcPU+1Ze+dm/+T
pVcqYY97PtBKghIeeQA38tzOwROQ/1M8LsyWpJBf4p3TZHm73ddX9LEBo+1P6lXb+KkpcxCBF9/X
thlPAiv9MaTxDMOyjwXbRTo890//MsVcgyMI8uEAWdWe6+MuH4ClziYFAempx77wzkbXL69Obqox
h8emFXbPySsW9Olmu2xAC/vwUbbQk+nCeYCY1FIW31+MGLrm0uiOL56KBAU9CYupeBqH6ZoJf+Ok
CohdOLwW7s0phf+Hp+oQTAgAK+LhDxdNB+9V/HzjdEa3ubG+QGQ+1yRv7h0k/RQhobl8/XQe94fE
7YM83NgtoD8dgkYiB6u/ibC/jgQ7nZZF3ippTVtmTVXG/m8YOmEtPDMVUl/lOKmMg0FiygEW5ysw
y1KAcc2equNhG+UUbTBCtXFFy7Gnx9x0fwH/zBcA6Vn2JApZR1DoRJQiAa5Lg/rl0mSVUJr4VS/i
Uve3vwz3z/NC0NV+Z+o4Nf5twEvK4f3jX+L2G1owNtya0hvzjPDoxK+L4F+7MG/gAoNRVPw8H99X
ZLFJJMLch4c979dtFy/0eSlp/dM+iENCKH1P5o/0X79itNmK+M6qCIHnNS3Db6G7abe/hbltPpNv
bJozxzeG0XAZYEWI7jnXb5k5ygApjpPedrAEu/+O5Z5szXgVsRVgJrPEn2t+CA9svCvOPWk4y+DD
pSz1DWzgjhXd0ighrjTqE639cltN14hfjO5dTj7ZaAAu3DUpcKfinAnp3SPHlGLUPtOiuFcvfryH
kmCGE2n884ARekhTy/XOne7vUEGGovdFoD7EaOS4xQCnDFXJZpMI4GpIexK9/SexS8hzs18mHACW
vTxoZvr7cjVoR13Rdlmn+bGytk8h6LiDM5jNwKVuBnue6OiMurnZye3RH+W4qBId4CGrOJTmE3+v
Bz6yfJe05RmepA5qsw3/OxSv7rzeDPspu6019P3yTnyBcFTfXK4Z2GOs6kgWhimqeS0suCDHZ3tF
6B2ufWlEqOhndAtmW+tCKZ0J2xgQ0HOSLwpkCN8G52xeCnjVRfuf2JQZ9zt5Ghb3Qy9NMPfywk4U
eApNhXWupkbi+iWYAe+nJQeWpRkVrmeBvCbAlvM8KT8lcw6OvjfaKIoLcWoZceogdDQCWHjzZo5t
vdoF1hlOEh4W0dezV9l6aONTH8zK18DYODAavuE3Wwyc3tvb4c1KTDdDyi9kM/leaTqku/4+3FCV
HuBArFixKgKIJG6otV7RGd6mIDyylLbUcFurFUMhqiCz/E3yXBnbf7wFd5BRMY+SGVn3BBZQP1uy
6Aeo+A5RPzv0LXqk2vVAwkg5w069Jxr4zuSvv3XPLnHw9wEpzr52bTyluNyAxeuh8+/VYZw4k/eu
RRfH7ZTtR9Wf1HPSCH2yYLvSIhlHZOCU5vxae4vXLJwGyACqgZctkHZxEQwPaElfDU6TyD6o/jKh
bcLSQDGDmutoKH1BVhyZ0WmESxNN0HdVWlIFCdoXXnyGqMIRFzf4qCALiDNKz9g0oZAsUmAAeqKX
aHBwqskbm2VmXntjzD5QLWH3bXQU/Q/rQM2xVjG4b2ACFgFSGbdjdGkad4B9jAkh/iey248bGxg7
dRtc3G6Ylo/3i0T0I9gB6PSp17chcy1D5Lnc4meNY75nOHN4Pa1b/Op/dzVoCuVe3lgFTfPfEiqg
dLFABDvun2a5oVYC9xr9A29EkwCZ+ahQcx74fbEWXiZEWnP7CdowMk98ihU8pLiwEKeGrPop8vKv
+Whwd0D0xvuMbv704vQ40ezsywrA9Mha2ND534cFW1MPoBOjzCHo+E34NOsaaST2F9FwiZe3mSL6
CaO3a0v+DPxhR3R5FjCyMw2YUpqqWc8PpGKWPBviEa9pQxGWgpnIvUztyAFuIwU4I5NkBmlWarDc
HZLcEzCZuyK9Bc4kBVsOkX1fzXfJ0NXc6P0qky1AWQSsymKXrO67ccDWKz/wP4g1LHyKSU+N2qwe
n7yHk1NTqHHcOI6+juf88QbQpVV6TKmRRwa9sAYFrh7zxp4poPJ90jkkEo7nhJVY41RqdZeycjfE
dhZAApLfdPF8dgUNpFpL8C0PzWBvWn9z0c+rMkaOQyFhlbIk3O2w/IhVEm5hguXfIDjZRpxuMyKz
vsLGSZv7o/webOanzVU/Do8iGiSIPiysa1bshk28zDcvE4OSqB9vcQAQQlrB+mtIduSOqVuqhDr5
znYNHNbFm3hd4Meagb4FT0+oXAecnGB9hYMZMzgbvLAxRPbds0zKvXfGNTEbuZp+6D4VUxGPytB5
+7YCbkWzSjBIhFiDnFBVgaz9iEa3PRzMB5yNKpkrc9RwwjYUBARZkgqJ2N2KyE6Wmtl5y0dgND88
keRe9e0ltW4i23yCouT/sCpaeZ3S1HwdvgpAhzFlW7p7ehRdpz1xzMHmKlB6e8auHLWh7gmlZVnc
fjryz1OVzBgCbGMVyL4zcVfSGjFWVjFo+kWgUioMifD/P19UHmtMw5TgSQeQDFEBW9xPaMurZToO
d3xREuziiMZv5ZyZPFxibHaPfzts5KgckeQUWmxecMA4K83qAkfxOk6uxN8eOMjEipya0vSjqcrl
97zyQjYtvpRiCcFuW4QP4Jp9V+7cAVihB001vSprB1Llo0iIVJHAlLtZMv5iUEvR0p/Hr/YRtMYx
arAc7FoTwZ1hZLtt69EIpemp9Gnu7Zl9BVpMogAqRuSfD+gWbjzJH/Ci8e7k5uM0L0Yzz64LTBdH
qZ2Pnfjm4FVIO/FWPHoF9X4TtiILfZJC6gLyxaWmsEqFMpOh1IRviGBPq9ZVj3gv7dbjrHM+C8HD
Ufl2SPD3UaOwehp/M2B+wt4CuEjw58HpHpNb5pIvC/kSP04aw+b78s03YHENxFy7LDQxAgXu7bot
8EC7Z+fCMDIfd5y61BfjOPqn2hDOzdZMA0l52dJFLl6EVEItFWNEHg54knkjx0rgwaLKr5qJq9Qh
EAPuSp3INlVIRLcmwpjXax5Ma8HArgpwHKCbcUS6WxlSGIOAiZLS51gCx1h2VB59N6YZxGk3XWgP
MBBofbyHky1v8AhiaFeenzbknhf4N0q21DZxh7UvQBOL8nvDZ0PS4tCmsLsVaWVqY9j2akRAMQJB
62tfJRzBVk1DV75qPbhi5s7NABKsp8SAQ7OP8xoeddzXENubEYItY9K32Lrf4ewsuDbDZhXpBqoY
5SvzlJrfZ3EziDVLwRnM+/8J/RGCKPIGHTKNcOUvgKMTtaL3pfT+dOgRc0jS4TlAqpbj0rJ6Ez6y
zFjXpfrrfx6r0Scva6BxEAW19CNR09UOw6r1YCzV1iKVElqwqR3brxyieNEU4SCIqGbblDHo1pH0
rqoaOek7AmWE1N0qe4vA1j9Ae4qAvDwcvJ8LoM16sUgDOqLiSsdBjNDWegErlPwubwKs04Mo1hA3
B0ygV+2s8Bn7zCaF3mgvyHGxJUwNyGG6IfKdMVbJpxrbKrDDJm0l+sVsS1lTSvMJaRtm5TDhIyIg
BCw0v8d7RJlzh9jSAloTWO/gwLUeG5HST6hbnZzdI8e5Gr2l9v+csaq/xh/+KTqIagwC93SRPiXs
pTM4cLOtmSWzCT+3aM9HYXgxsIC0VhDd1izZvxrhMpHrGhyO2CnKOJlMLU/IzV4IfFfScfgx6JMu
5UhqBRWmhZl6DEHw3c1o1Yg8bqfO/LSnXt/6IeltdPx8qxkUxTcPNXp9jOTP6fivSpEqyB6ENjR5
xNTg9dIq7vJBTBH2SA7mqM8hVZKz55RCXGWYdA1+vmW7RLLUqpFJZBDouitM3daKr0ywBB0HidKH
jBf6MZ6C6o6+QOgtQzry8/MhGSiuPPm5n+rRsXHfvoZoZ95PALjxAaP1BlzRyFCKiD+QFMq7Rtfa
vGVGG9QgGEHiX2zbibRoa+AKnY5Gy8AIZIYM1Y+6n9fBOGl3D79KwrNx3TuAM3BXMALHXzyVsu5A
K3Vm9hoXN0trT0l1lSwm2bC4FrCqXMt7PvBwBqIHnSzfbZInYOBnr2uQAI00BhztBZ/Jw1dktWfd
qQ/n1Tx1rojzcJfhsmFzjujbZ2gFVHEtAuKPebig8IO8Z21ZMoBSErdebKQzA3MUDkK17NjszCbz
kA/GcpDOzW/hR8goakX3s0QOW2oHqf5mGfsycfV4R28Q9YREyzsXswOP3IpGTf9WIJPYffAJ9Whr
zMLgSvb0Sa4+l3izK1ZXO046xH40suVWVKXKwQHdM+00hGfV6GwwblJ0s91Dor2q3sdsOzAYQWdI
4AeL3d7OtqPuh578FblPN3+6C9yq/9ezrrKDuiJxfLje+ObK0IfpLAJ3RlKICm6FpJhvxydkekiv
NdLnUE/XG5D82aU8hiFsMX6FItGOe3oq0UQDxilFHD0NQ85cdNK1yWt6qHH7QJtQNZBXMJPQ2xuM
9teiWDBR9jl+DxreiP6DweK3PnD8qGXKtJJ66qQ62CyP5R9kkVaLBTS0TEG+4cK8+f6X7rMcYSIV
njcunl52D7+4P556eRvELkomWt7XG5IUmXIUrzJ0ls1xmTnRtT/L9yspwT/ENB+nrN54I2kyP8N5
RbPPB1bUE7YWpwWijmywlxI6Vl3zQk3wKevyqhCl9YuXbNs0dxa+fxY581fqHLiRxr0VBLLMtfrp
jbrgVBT/015R82neg4Dkvn0HLQvvlH18R7bH1S4tkwMN++EV8KhLwHEZ0KBD3Va1cJiZ14OXdkGj
F4i+f3/4V9zE9wLdyTJxF8O94nOO/JGNJ86HLh98oRSLDRyUFmue/T+ZYbX7U+tH5q8PneUtnqNV
DRpl51UwcpMKlQiUSv7ePOnwNoJPELlv6ephFFybY2nJNYhIoRppv6IXAcWutWrNSblKc5F90xF5
15vvSO8J5evUofOb2zInxi71NDW5ktPNna1kQxre5fg95PjeHGz10TPjKxD0/HWdjI7oJdQ+DFtK
tMN0EE4r9hO6+CkQrHRxHGpvUlQuueVWBt4QHoDH5UW4Jwahb1XF18WOuFv2Z9piAjRzOvaeDGwp
FmQKFhvLXmzKnzFTY07qLjX8WGmnqmWe1qgnUapc7q0j0uEtNYzV9LrjrSCqr2ncTB2nms4ahyFO
55uuktuIcncDloNy8/rUfbqrmwXLVIB5urxbkU9j0bf4hmELz71teI3hR9X8/oWeZ2m4fpeqLqi2
nNe5z3V2ysILEyRfbjrRNO8k7PCyZMW64FGIH2DxJpJi4efLqOiT2bTWefcTcklDQcBoW8p+YLAw
CjxJ2nwYm2VxuK2qklq8aon0NHnc1Hr68wbNVVxWm/iVt5Laeq+a3Pkjgr/BbbtvjyaKwIUgSe0z
ZVDQIlPMGJC2e8LNWgvVszyefEKRVzPWCGou6XIzke5UEjTdRuAA7r7hJLtlxiZK1XhzRwqz6npA
n0bYZT9IwiE/+8FNttMa4Pb+tv5XqtQLhoR7jbQEtzC2L5w/jScIliXLp6ttnDWRaDQZLSRcc7f4
v7lptAgijlFynGpOdHGU3GZoSJtXj0q7dyXJghHxzw+FmVXvBuRbOMbkD5YZg4W7ny5mOzaLxfLZ
R7okTW0W40SN6eS5T7wiWtY51iV5QXS9xYIVmMSo2P+6xzHSH1mt592n4KM7ooNyje+25929VB4z
i48vkEieLbskBFfAu+fFIgtx250VNcALtJUnyPy7xygt0rND0MvmwCwidlSmx4V22nXuNk5QcsR8
FtYM0g7CDgLUuUQmxpAVeNVLQzcLVW69ORP0PmajnC/6M0qfQS4Em8JesY6I/6SYVnGHVUa5t14+
H/Lg1G3l3gCFIIvBu5olneKJ3a44lkV6DakBBQuXOwjgzMLEIgA12mg9cQsTG7/64e+2ruOCLL7S
vrd0G9odyUpgPIueTTwEL/mG13lWr3SrmAqXxaa0yUfr9Je+YszZeAHWx3hD09/aoX5A8dIvrKA1
phS8TDLtJCSCbwCfWHk4/BJHRaZal2zdI5xR3ynfFNdpJsw3cmWSn33ThfSZdgrThaAg8UAH6mMU
IZvG0cKV688XJFkpzBudMV+dBbMsad7HBWWtODYdF+8gxPL4saweYDTmYJ+bFr0q1LCeVGD7RsZW
ttnNA6TjLfo+WTeW27Z4Pq2o0f8zNXpc76Pw+R7AgIwoDbYTBuTK56tcbWsEXz/6+XgDrtQLTDaS
yxU1qkH9Lr7T4bSa0Bfwy8IUAm+xI3lMVfkRJKLXqATC4l3xHJSaS1hHXYL8R3ceqMYTWR1TEX7L
lnlVkD12OHpI99wD1VkK8FnfLxeO0EyuVu6XomZ1sCDbLvmo7wThiOVJkCnUuoYV1gxYF96PJm+R
JJJnbNDqHocxG6mx8IDGkn3qZO+X5tob3augDzC3g3AlpCRqCxb2vKUp4L4p0S+Juz+jEzxjYWWq
Wp+I3OA/YiiM/ZcjublnduacjSvkpC+Ab3oTPOY0yKs8wos0DjbBn/DGI4GZXPffh5513ZxDbGNX
A707CIBLVn/jmJ2gpLFQAsB5J9fH+av0VN8ugxMSzEZ6TvNlXVW12MGitmcmNl3oDRpVQov1RSCD
iYc/+4cbGnenunHRNi0XP/ztIfFXx9ae8Ajyj9r7lEikdRXXBavSUoS7Oz+NBplkobA567b2ihTr
mt0CahR5FcpIdSFCvBEBauUnOed0XbDBfZ714aiV9bkGTCrq90rfj+pGEqxjjO9dcbE+L+CRE6GO
FrFcDAFHUBr50dlBJdmk8A73viEf00U+MNoWdWA7eXYO9pH9mcIFvMqMoPx1UORpGs+0cImpHXIo
hA2F3L6ApzTaab5XphXuJbaP1Hk1CfKii6v65RxBToR/aMYUrXG08hvNfhk8C1SdnQdhVIATLPTY
pnROaYkIoVJnh9+SMgv0E0YC+NzYIusPXe274LgWx8YbBZHy7GOAUiiH3TInGXYqMzN8GWAKVEMD
M2BZRFu/znDaCmeHsq7BVbq8zyD2v4yLsZYCUPO/bKXhjiQ/zXS1qAjYY6y348oRIsROBelyzh7E
zdr/Uo53KJd6nWzim+DljwjLnjrRfXeRRe3jYRfHeXLDWOCVEe9AqP/7pCFJ8RBXNhOOHqfXq/69
Fax23FxncHOXqhvuPgSZdKBrZOE3IJhzHInn5y3/wLz4Y86A13muALnflmKGMJ7a4w7K/Ch13QBx
y+LnrD6E87R4Qm7f9YLr6I8DFcx6h8FOY5AIsWBg5xnMLiGDGy0xuaCTB0eqO3Je5hqR89gDJPn9
wEypK/VXj0VQ5SjWy1kdxdfYUdSs5Gw1Pu+qNlCOt0vHNohi17XvRYv666R7IXxHepK7Ui5zvuT0
ixFsi4Y0111kPA8rMJZevvbpRLXKujlyL6qaVYwzMYiyMrAP0VtEYIkJ4Y4n0yHhDzceS6T5PO83
7rD7leJR/BDneeT1gZWjUJKFrwJJ7HLZoQpVKcrHr+Vb/nBX63PC/RBuDYHTJKi1ohcOoLkVnIkf
CsZGBR9g20bRkKkfRmxLz9wswiMsYw8G6FG9E9YEzonW5gBG4TRb7FHAoF6mjOTiNGETipBuhyR0
vP35gsGmNKrwzP3tv6OJdXdZXmO/walW885VcD3WqqWCmO9iGUNI1cnyuBquHfk/ZdcWlmmo279h
FpnA5VwutnLn65t7oJX59woR78AargEgNon7n7nG7GKDF+3nk4injJXFO+xiem8CvH5cHFj5K8oj
+Ft39aKoeCreR/vMyAL4Pz6cxCSCoDIwSHatVN6oqe+UcLsQ4bjF/4eY1hU4bunIIagzvpIACJPt
7G4TRUVoJnHC5mVJkA9kKpC7UMcKr96t83stFapveO07Ifb3UGjNvotKEkvZexu1ztJP8oaTp531
20uTDzP3rJoEbVk533EWyO01F2bh8u6hZeFkMvc+1OSdiKKaiHB3LlHBWx7AS7O0Rwf08mnYExNR
mwQZpRRTy5Py4ywdIWm1pu1y2Y+hdHqGXpCdGXmq2Mp1Lt90Nb5xFRpHZ2cq+yqIBDa9Qfu9ZkYj
ccABCLDNHL7NN1MkiOonwUvk2op3JOJMEIRqbLBjTkimiWgXXltN0w70ZCXKthN4TIfkt8/X0W9C
qVlHZH4LjPrZSs76W7g1Ol26/z0pAr5kPmeffta9NYiFajpALw/ulZL9xGLurOhQNPZ9FQ3FDq3B
sthXVcB/tEl2G9a8uTTCcgtTfcuaVMdOXoiyuYRQsUjzBRSYlVUIOc8++jqqxM9KGEZPF59J0sH6
F161HDNOTRnoO6ViJN8IjvcMkKMX6+vPUfNIVjM+TiB31/SyPYSv2MDvhrJQdi+2/vwNz+i8+TK4
TAfxn5sTEBTk9psT88pz9U5pBB66JwGpGqwWwMk+xixr+prBQDQa/m812o1RXMfXuBl9DTQactXl
QlPqyIchi10yrttObQro0Gh5N8om45sAyeKyqn/7h//IFBRcoceQ9GedkIqsQlIpicqh+D89zMJb
O2KAjfjDuLwehFKu2LjUiWOApLMsdk6Qu7K0mOczHgMt72Z9X6cYY0cN9LXx6EmA1B1XAVAAFapD
uZRSxoakny3ml8YNjYWUkxOkOoTkdgxe7b/31Bl/l2WK8q1Q9W6eH61IIVSduECwZWIIeIyxUtdF
2eC2qJGL6Y2F4cRuta8Vdo4xJ53PdpKALonPyf7KtKLO9+sOl2H+FiakFYTU0pAYNRoIk4/uxGYl
S/3w4KDCeVt+QOMUG7Ik9uCg09ScNEgrHjBd2kbquYzWvnHUVjduc0DO+oTWy0XCBs3+SwAuHrgD
mFAaI49gVr1yM0wvuPYrCuE9zGuPNkOgAIugGEbtlHfUYVtm6/jrsHZAGKgBFAm2N1Pri4l6MnZq
2iRIg8sx7xXH0JneZkRM0p5wR9fU85v2qhxn5RBAotFxcEbYiwG1J6e+mix/JNaLCG4iqWOIUeoX
eaRsPXYuOhmadm8BUEC4VhmB+gW5N7Id2ArAPPjDhsMKwNLKl6Ib68tzkTwMFUg6SFb4tfkE1n1q
3qeqBAzww/JiQuD44mip692PFvyPkgGpC1JxLCOacgH7R1R/5+OmIEPMH8daj1hAn8s+MfMahjIq
HEWx1LjLCW0sTYY2wPjhUKn0WKdxOXOF7DZV05Vy6qN/UISN14KQdK9NgllzMgDylepD7M9y+bJM
2R6UrJDqEKWPXNgeW24sas9CFcC7hHWGFaq3QfmYPavBIN+iaWxlYQwCPI2sO1rqZi7J8XJxpIo2
Jr/qB7usRS9wpAPbQbqeeAi42IV3PO2i9We3391n0SEjbmOfKdt4R+hcFkBanOhZyG91AA92GbR3
FG1RpytWuzdiPS0RSoGSd4EaQQ0XQV/J/7c4EQu4PDM7DHqw0gzPaZ8ePgO1PfVgBPE/sjAL1MJ3
G692OBJrKPrCO26/04fRdwWeqXjAd0M/E6c01O8oBIQbI6pvvSggGq3te9Xqwyu0sJ9nPb0Fay93
QbejecJw5T587UvlXgTRDH2g8/TOh9deFpi+IrdRxLoRbl5mYN5gDUdSMfHKYtPQmTPakyYd/IlP
YHT2yrSsjqOPoXlhvZ+IfF0mDSjViNl2l3PSh47r1Wl/a93k4ll4utsbhbFM2nQiIFjXBfnV84h/
I3/BFFnF0RmGCsTF0nXqQSJzZIeJ6fPOIdnDV/ypN3pP5wr39Q9CcMgTgnkcHg3oIVg9VKrHQFuq
2Yn2Ck5b/lcWoIV8QLrT0FpfC+WXZPTMEbemmxX7m3PUkwpVgBvWdseoRHf7wItMSj2MHq7gzoHT
Tizgq3MRtgpqB9/xfCcjnK8XqfF6Q20JyRjcBJABdeBNx92wtME7TWqJt0qhPDsHzS1hJ5FOYhb3
U7ubpJi3TSn9OkAd9T5vBbWEql2ZBy4Ce5L25WZO58G1aKSRyOZOqNckz6jaZx8I5hnve80AVAKE
IbmezNlRo7KcH6xtR6bFVPP8Pn+1yQEiSBmpGxxDjhnkz8Xax/lxR0E982nwlo5gEesudxXwgs1T
+sb6PjkuWd2teQ2qSq/RDDruPlPR0smyXdtVqKtjaqZoNXi26hl3zsx5upX0ZLLmRpvwtk+q3EDd
XYZ3GRR0g8m+Ji0q65Qm4cDJWg6qE8LxGmSqAD00NOd9K7C47UWn7ZPfeZ8zTb+G8WItexMwxlH4
hgHJyTQS04L54VWTYhvxFDDSVr4mi5OlE1LJb7oKDjGITqJZrtTRp+faMKgkx5Asm0C4ezkyy1uH
f1IERtZiNbCI0h3luPo5Kwxwuy+MCQ5o1PprfB089XapwHpHU7A+geuL1+YW8a5zgRCD4BWBneM1
b8mu14lNOOP3HVEmckH5UZXCnepnKDFMwS4jMHfsyFeLg6k9PRhsKJ3ubizpnadSd7TkhnyA989A
BSNYC3JbI/DzH4uLGrixIKQMnFjDSuwVIzc/USDJDcj81KdFQS/tW8cYpD9kWU5UWSXnsG+xm6ZS
BIv+Vr0VvtgK9Kv+lhC0XMyY7nlPzc0xOU9TMBMKPJ7aAqlm9dbfuF6c4GpAwZw4Zqne2+WYp81q
y1mEIpZKehP41F8VY/PnsCcCi8p2AMmfjuWArG9yCIu7mwRsjGcfo7883K0xrhnIOAbD0XUaRaw6
OHWMYSErh23aTkUstswcbvJ7A9MGArIx6/f7zf3sgoVad26+5DRJhsJQQe8e5Xb2HfA2ONK1dP9Y
j99WYwYoyhC/2McKhrIIXg34VHgPNM8t7vHoKhRVPqfFSnN+89Jv5vYR1CySN9YvnyW1DzLh9JVN
jbLTj0A9m4QbHevmnoPg+zaUP7BcIV9rBIPRTbIF8lWxnKCOFaCyWkuER/fkpjYfkK+EwQYsh6b+
nv8Z+9MECfURWjMqz/xkr7zgndKoHMa1keHWakdp4ISMDlC94sQMf0c0NTIcaQ6osxvs0QzHuO2j
akIUMe76u2b5z6qDmm6gvI8Gaoz9jjORsComK/W0N5hqGoNTn1owEh1o3BAHc8SRJpDZfsQP+82V
/1M+jTEaa97KBTw2OIXYrmXgryRlYauKhYVxEBcziZBBRHN5PzMKpz8gFXakuUaBHEKbW3YD6TkJ
x/N7RiwIDTsdBBpFMk2vUKlNyTa49QZ/BVAg0c1yJmfuJ1KD0OJD2h/2MrOB5x1DJFztRqxgHK1m
s7eepSFULgvC6lh6r/g6ALEEnuQcTytmdwx0hSbOwWZ6NDM/4Fj+fCSxCFFV8tMpz2sNHtc1i7Ee
OBGWKHvaGX66/NZFp16VA8bxZcPsPmbCRyx3FKTRlyVMi9tyGE1gOsJ8Kdixu7yzItuXMfsDjQ5O
N8r+BAjuUJByrQDlmy25weuhXZJSjuBdyGE8hpbgmEVbXkQGmbBrS6Gy0Z8oEkaK4ko6+nIA6LGp
ftfiv0+ngx+pooIALWQlswsqXRSmGkGRfOL7iGnEHX4BFUpsb+FE7lzYOValEGxJSMGYfOZ9amks
G6+MC86g08rvUNN2PZcpAPi+lPmbpgDARGCgLiwRIrbYScvV0z+VlKp9d8KOxmvoPY+4GSwUG9aa
Zif6uLCi0+cgUygjtanx1RW8WlRv40WCo9L75OaWD1CdppDoxe3Cld5mm2+b2xQt+Uh1TFD7QCzW
b4yzhL6/0rJGB47k1PrnFTIaN7KEKiiSmT8vnwNK4jXAQ4iuU9Xyw7nuLmBd6UDYr36aCA6Wb1f4
haSWCApZoAUMEIXHGc8ymBcADhGINeGhoa6uC5VzeO0KIYgcgcIsOZaalpAvVf0zF5iMetaP7FlK
2GUJ3EfDBilOb3h2322en3pr1YfsGhywhYD329nCrtJa6WRUTOiYSUbFeHzk+BDR3ioY7vFNyQ2n
mKS4YKVl4wqJLC9rjrILFy4+nB8uZfR07Os5FrWCGND3a3GTwV6mCOcEGjTV40f56rBGNY7vojfd
Tg5DzNXje1RHCJdF/L8EQ7WQUikfw7MYZ2rk+N6afKhZ6w3AGoNyFAUaHZF48hxEfdnFIWmXqTWB
dtsbEXAOCaUxJ8nzcVtrNuMuAM89Xudk20kQzsmnJsGvt6qgjtXryykNqlQIkIQYmn8PB6pZowNE
p9t6swdfob2zu6zbS2+gOvqTsEOO14KY6AiWbil4z0PYgPZs2l5lizYEpGmJ2E/M6wcLzvksJkIc
BkQ/go4tDccfom9/lEYkQkJXriQdR1EcpQBvkWLoURdGco3qYeBbNTVW4xnEei00i1d8n470PaQV
lQY3TGdejmkReFq2S1yQUGxZiC6poZuAEGUxyyf6z3sl/wheGRGQniaWVVBL/Yz6kU36TMwcUbWP
T/RCgA00iEphKG+TV806fFocPxDR4BkI6LJSCqFII0Hu4z3vcTbQkvuQkm8LMKo7sr0gZxo0reHB
4Fj0I/Pr7j0xDwVzaWnU56W0JTaSjDV71HOHDwnaQEfxKfFw+tObjS3ypNaYC5nLZpoKy7YADA4G
7tULS7+a8FEUswPLRjVKbPrjvbjE71cMT9MnW0Ekmcxvz21L6YCyV3cd1U+7Bf1/b92r1ut1Xiud
Jh42We5LsfJ1ik2e8iIWVr/JKUWT3wnRvM01j9pfPGu4EipEQq2ww7wmJkgrlk9xo96bCKQiDSmY
fwl0ySEABdQA/i3C3Wt1uJjIRZUaWmDWFnTsiKW/H31TJM4fkB7wrROY8o30kvN0AbrJtk8yBAeY
PGddz/JMOqxrXhx9J+KEYEpCVsCqhsxP+r26KIylkgAhmRy7cd8PpGA0e6EcomGRTyIDg8NzQnui
g4E3cH+EChAmyOEe2jlV51vCKHEgKE1mqZddVkz/qdAhQqgBdZuVA8/aS2yXe0Os8O7mUXdSdccy
MbQ1L2I8MrrW+4ofA8j/stqzXMy/kT+EO6TOp7/yQ5rOIzqpkW24YEZcQzrqbLO7313H02pxT9vi
tjS7uVx2hraV3v4itM2YOaVDAK9KUawqGs39+zxq+H+0CYJmWPbsq5KuZsGiIfOMOimFm0AmiZwc
0EzWvWmaGv2EgbCZoF1x7HTEBLfxqnCr+Qchfx61G94oA0cqG3y+1DIz9salEt04XvlanqXXSBaq
G+Z+wWUW7cWLfGhwKFrYeFcO5iki0+K0/tOfqj16T+9pv8KHYYV2bvQtHTrOP6EEJpbw32KDmAaW
IxglUHS7qCt2k63huPcUZAxWzCQjLtK0IGSTmsISLPpN6hdXBK0EI1dY2/9wQfGEie6uBH/DEDiB
tJMrLw2zWw02aWh9zDOsw4XaSAvNNca9cwO9QufV4d84l66Y2l6XEeyC04BR19IAo1+KSGGz7wi7
WPbS7GXZpoVilELTm0UPVqpQ3lpEzHxjj/6O55Og6rE5h0N5t6WuKncmXg0uyX/UkURl+eCqx6fW
H5PEcplwYZq28nP3hoM0ioxF64x+eQ+H1wUiEsgtuLN9DPXgb//rfm3osYyHvXGfxASZ5Hpoo93z
an7UJpbCEKwUdTPtDDxmbGW5dnaZXhl3kcHVGHCeGI4DlmSymEUZwr04Fea3gkWRe7AZ9Rkep9XE
oq7WdfQXhhQzIkrIURSJofEI6dq6opH7xst7r9OSyUdgMe7wl86HFBY+NYnqczD5bRKM5ajjWVGE
E9E66p7WUAL4oErKCQzg8JKbmKraYy5ugFqpR/dubW7wiFZh9wSAlsQ64Zv1tYh0rd5CU6LA6Oou
x8cNSORd6dFdBbw7IOJ5GsmlVoN2sCYR3bU/avG0LnrLcygtVSCuxfLNxIeu8/9O92qHUoeobdHg
roM+d9XY6PxKLjOc8uwsfBe7a31pEDKZED/WDCAPYoen3SO7MqmtHjPi01SspDQANFywtcvmeMqP
Qgu7ZmpRCXujSvyQZ2UQXl2e/PP1l3eVq3VdsAF9tu8TKM3bFFj7VaW9oH+/ALaM2utlAiPgIbR4
NM8bfptCRirlS3gfYMyf/F0ERknlymDcDEVPcu//e6oOFBdI+GWFaaquxKYdDYpioi/ZK4AiiKBM
rYsvJ/TJgSfopJL3/KnWsZdywyF5h0OuWzOQ3uKsnBVbOB8rzVAfmqqYACq5wqXy3rOSqHva3dT+
uD7P14xI0AhUryb32xIY+I1tErfvwNE1RFSnt2VoHe7cyUADdccAixr0h/+fuU78J+yGXpYcR4Cf
+WnV692zb3V3kmxEhh38VIzDRc09poEXYQ8ASX6SrhbKCLkeid6P5Ckuc8z0rVmSaX9uXUEI5XR9
N70uI+XH1Z0OWOQxy/CJaDo6XwJFX33quDNYrkQAB0VWYTnJ94X7lEwh0Sv7p/FZIEBI0uywc7c5
KiLOiNQQ9Uo6MEcc9+mN6x0t+9FqBaB2E6Rq7Ae54DuzddMv13NorFJFXBZOS3WktXJYdaHqPtDM
G8vhVip1lR3FrvlyY6Fvq35yzXfUezPsbMHFdJSVGXDcul5GhXegg1G6ZcYcZiczvqewKkm+RN2r
A1a6Nfh0ZUOBTbheh8AJi5P/ofaLRxlWXct1Q3Hz8F9c0N+qyIEFb/+rlFGeiJw3W+MKgtQ84KcP
TMGPf+Ynh4pYD/w1/34BHmR7sLXfxz/Egm8O7kh1XMnlY8aH8jKzfhgwAiMMdc/GdP7JiZdiZBlv
vC+GYSTaf3tP9I0GTHOcRBNETbpUfMWb4rIAu+zLjADli67piU5xFC52gZppm3j8TnKrUq46H1TG
xxaRFlK3JSz6CnJZymtbhMpEBedUUmHjEKNINKhmxv26KQLFXQ8vEPZpRMLSQfZI4djD0qDdoezZ
sSWmmpZ3Y0YopermuaoPhLRNNLpFqW2+Mx40ra9NfPYyFw5QjO2JtExSDICKiIfkj4lETuaHLEmX
3dXkWFT0k32bFRVQq0iWFpxYO9eukYEuFi6L8iFLUrRPP8VXuUVTxsTqXe6Q9to9FhBM++r5Le8D
mIobZIOZuHMvLxMgG0eaxWmmod7EJGySlOu8TA3mrQSdHc4itZvFmJxPeWlrGuAbT2cdkqtonL9u
NlwhZOYh46r5QucmNuFEfS2XTFXvNAM/DlFoLEBbcw6EzbMiyk68k6buoCVGqm7NJZXdevA8IPaL
CqImOwOPnInHap96A+aJHgUgmW4DrEn15szwIYPy8z+QvCTy424iPTxKg2v2UXYeJmDFSYKHsLSz
w+IotvHoYb7XyZ0s3vtWkUdVdD6j7Q+4uv8BAfcm9+x7/ubXzF82XARDm3zkl+h5RfaFs3x3/NFs
WWTpum55ZmtH9RPrZs4xE9V9RPeggKFIN/IF5KvjWuFbPewGheFP8TSg/Mvq/omsktsjdQQPrPGe
81vRQmiT65ocY6nJGpGBpxFv0GRDwvAP/b5ShOeeqInDk45+EBHbTDMR95G0kI8uUn4JGAKOGEkj
IzXNSALZ/GxuXoqK2ml0edaizumD597Nr5B7Gm/yy8LaGFFQoQZ3POAGbHjrc2ZzHG+c1Eq8OJt6
cz7otCJfhpBy4g48n+WhIY6bDOJQUa9v/3HdnrmOOoSbI8IYqxcsXeaGKBMiFJiPieWvsjaVEb5w
wZFhUAKY+adWM/kYxZ/Z08cSTiuS8DE1R/BAhUZjk5PoD9q32wtGmQxPrV3CfUODs9bScRPt7GNJ
6wH8t6F+o+jXc1nr92NGG5+fFzhzLASlKSBDa69v3yAJBPwvA8diqk1cc+Cb9lxwslWtn3J5rGq/
klXFLY0kqbRQw2+cM7XO/ZyGKIZLXuAakjBbZEWt9nNtSTmkyRpBuI5BuQjCQAG0pc66S0xqRDtO
t8qS/nvrXNZtFmIu3qzztlsn/n0L9F2SBQ5pxFrZ1QGH0fBvd98NK87efa6yiFQJUMlYif+6dngP
o+hPha2S/CuYJz0wadvaUZIX7HZs45C+H4AWEVDTDKx7RUDmmVRoiS0Cty6CaejZKZl6Ygoymfdz
fmb85rF4kBZLdpSkOHpz4d5+EuNSlBOscDd6ZmnE62Y223tRXbohAhYZ52kwISqprcFwBzWz5h3H
G++xDbpjeKWYROyd9rZY0gxBkoBqrcQrLWVMxHJMd/KWAf5dbuHis6l+60NZ5ouGcO1vEmXBpmc8
/7GSAKirbYmWfXbhF2gySSY/uDWX5SQ90pUsz2jP5BEAWtsLc7sZAYTAKNLxk6Bc1TNzI217JX6x
5yUknp9O6dyhp3e6FgMUUdEl3CarrkLZZdfjrGZt7B3RD6quE1hzLM1E5DVceIdhYtzvXfqWGR7c
ywnM1QiFibfDYgbG1v4JfGJWMDoiPkpOWZs9Lc9x5ivpMlOSf2YZ+dTMnJJh+9BWX9Kl6f4Exgd2
blfav5srr5Su1dZqGuz+vUjreqTUwwOgG9zsjjbB5lnF5Kih25xZzEOx+bi44XvIIyM6u3lsN0k2
yVxVC5azPmnCgfoKDzgORL8Gsvgulosh/pPgOoFbG4AogNk3yTC2hD/KUIP3p6+wTFLc6IKnOKIH
qAHga26i0fpk9Cy8XBuDa+23fv08X0Q6Vz6qYIxhEuo45QRO+rGr/O4N1w00V2oYxCFgJZ2Ruzve
Isyvf/scHPK4uALXiPZIohb5BYVJKzrVEPEJuPcrUFgB4gbg+TE0chbK3mSvcfXeTwzxeIxOa/rI
sfdjOFEdnMS1VzqQIt0SFvwa66bVCsSjFEPBDAt0bmY+2kkwPJVvwoxuqzYHcvpyut6umwgMLvyW
X/+QlUClLeVe0te5RYKOXmtKqcx5bQzaeL2iGtb5sr6VfSaseQ6Ky7hZIyeCsHn0QbyLzI3zVRc/
9ZgOFKE8mZZ/B7sc+I2az0D71sw+l1+/mFQyplTr3IG5AiGy1fqa+27DeUosZ7ISunzrVh7dlBBb
i1juUkrYcyrRkpS600ZWHfln/fknOEG4IG47OvNgEHFT/KNARMhiWq9iA7NZWfGcHjNAoc0OgoWp
AC+V3BbogzSztyYHqrx+vv8gtG8zxxvsophZc25vh9gwhLxv9gkftQCX0Ti0QX/Wa7rsz4PeJ1j9
b4k8cgqyQ84Ibx+DbShKUTrzpClATsddt7dWWAPS0fF8LPquW3U4pVkDcRASLVf+wV5outJNdESH
0UIkb6GXLzO06mXbokgZtJgKwB4gEgzhukhue1myetQ89Mn6fCsTmdAwp1xEAbdZO6/kK8TYrtA6
Xv5XU7z98K5sohgXsNaGMS783F4NBlpAPdKceb9ebxKPick5hpadcK2+ac9/5a++9JOfW73RPWwr
8keQgH2Ic1blZUzLbF1qz4H/k/3yYmMVqx1EIoxeJJK0VCGVPNOIz2vOO6m3mEE5e+wcGqSY7A+J
03cDMrhB74Xy58AZ/NR9olPFpjKENjas0ha4pWYX/guFPUS4p89fXxJihOKTpMOuqxcqV1okknc1
xelu3AgR8YUKrwrzYjhPKhJ8Sau7MJ50Qs/ntMCardKUKsWZUNJn9tXuwQXRRrcZYsHUDCRRCRSl
nic1WoahbqyILb5GHSEacw5kJSbm+0gyKHAYj+PSh3stQ1Tak0S2SlIgutBlfbMsd1ALfb7ppZKI
TAxha5JCBMTYduBvLVyAkLt1+92Amk5rD++XKqWWAxVnrXGzETOsba9fVWXhigHxpxI+7KsNOG3l
h+inPzlRu4rEVHEdF6aVUHTRbrFQ/ZcfyromUja+k0Gmv+cUEtk3UXLmfXsUlEMKR7zBoMFpnYxr
if6RoOQZGQamhl9cfRV/QYK226b+wOvNJqRQsHJnFwWURdYpEQw36xfkovmyhXcLiys/kdKzNYgB
EpShnyTobVVzuaPlV5fO2iXRfnz/NKzKkT2CjNdiEqMQe7T6DIFL5GXoN4oB2ifjcttaG5aU2H6U
/t71jgBW01X7i7MYhPWjc3/2S8Pf5Hwa0ZXDnQTNU1Vqh/ph9wwoP1WJAWvhXSwbO7YXPXWNt8gm
k3nneLcnKyHDioE0Q1UJ9tZz4LA3A5QjQWFEPbI32ystkHrHW3k63MsK0GcDQvvwMA8ZCJuE+5LX
P5/xQWyLgz/PY9DSkYwFKGdZ0c3bfXqtFaPbF6Ni8q7LMls6REyp1Af7BJrL0XLjhPVoN7odsO6Y
pBuxJqAnm2mD1e1uM8Sin1jq86sh4dg1v88EMQI6ELKUg/iieA7cvmNDfPeg7q8qEh0Jw6x7rh1Y
uX9Ca4YB6EqEEc/dTKICfU8C8m63r3z1+B5ix3uaNG8kgcxr7OJs9JbzAptAgqI5cLmyajRAs979
uElKJUdkDoHPQLEgRLK8p+y9aDeD3Ferl/TcgEnHFRlfNeJrLKKuyyrarxdm3Ql65ao9Oq3PSq4g
7JoRZMbfjaoWo99v5S9ooGcY5Wpkn2wugNcAuf6D6v/AA6qiHhYABiLfdE5Tu97773Hg0LjMfJEI
05uEBnFMZa9WeHAVJv7uFRhDZjhQ/OIDeePtYsawdPemudxV8yWgQud286L3NK+AQPZOExSOr7Ty
4zgoA6iWfQQAIGIUwUrgTBaHo2vo0tZ6IJlXyxEgqOjIc3Bj/D64w9rBevXWp9FSE31Uc+T/5cKz
jx28JJaaxkRjcr24q14cjO1DiplBtQP9Von/aCQ/Aam+dUsPb5hbSZK2Amhf5j4F1k6SLjuPJDkd
SvNvNMLCMYzf5QbJOrJV3U6RlKapiofQAqiXyvFtHK5JJa7z16BoW8mINsdDXHRuz/Hr7bJuppuy
XgCFWDZz55nsT8ue6/BdTmAoXgHIb6niTH/FybVaAQVxOx7z9jpwYLVl8rFMwlt/bmbeOSBZjobL
VJ1vP0wAlpRAXJbKYHCYQJYU8DODwp/tZ2M9zuVezBPhauA6WHUgSV0XclCTWoXq2bLIxrXqhlcD
FwyXPAPQFS9qs26Gh9xBDsadb1kLTF//Dyo/yScvHTBzkzPp6R7L9El8qSWB0ZASVPiVvEEXelPa
q4/Qvtv0WfCOwgFzqHn9HOhJH6KGvXbfhm6tNep9r+qMvzdgv9HyYmxQaaGZ7O4pIvUPlKtvn3do
xKj+EB02gM8IYvqcC4JskcpRauPi0Vp28V2uGgF7+2VJ5k7qqBn0bA1G1NT2gtNIPhjonXHIBxUn
3Ba9oXf5a6xkRTeGSWbkypmaUmNKlVa302dM4GrXsV6Vl38g3s0zkiE2nLyyvX3FbnCzr+RqKgGR
0jyHT9DAp27wbE+5pHPTqTtwrYEZsqxTWEnNhiTLv87hWAuKIV5pxu/CV2FPBrrU9qJgGSgELjP1
ucfMeVb/D5zUIVDWexB3yOmKY2EQq1Y/a5/5wwgT8tTV7Ts0sTO6PE7R7TL53UoEmmZ41cqjlYf0
CYyefjEwikDPgKyDHFN0RoehAWRvORTSU5IoTHyhvmZZEHWo6MgPjky8fo7JBptwldySoc8tvBpM
oD5NVY4y3CjPuTNtTNfYn91NGN8RCeU8JSNVcqBYurvzKd04AnX0vjkb+5137FDOuIV3LSzu+5Uz
FjA1lffA4tfMQMc8PpPfo0HDDeSD/I/m5p2aFdkPWw5+GNE5IxfGpSDK7Yb1Vpc9IakCwuUSrILG
oTZ9xNTc+pIaiQMSCR2VNhve2HamiqqpSvFbcovr/j8Vi0/3ncW/Ms7jMpuPiLVlh20NolBLdZ0T
D6zA3ZApN00ruiAD43Fm6C8mqPz210lwWK7LSLp5qn7hNB1ykLIWoHIZSE4OCsSJ4rzcYtfNrJQ1
NrVkSTp88pPELEy+5dmGV1TK+7gzHxwu4n0YIypn1TXtzNqyo5LW/RFBTxYK/+K7TY2Oj1LdSxFu
bPf6twnLlVBS9CBtj50nfHAXB8vm6dHBxCHna3pMWsnpqwNhSkMDCTqoSz7D3vTP78FcI9gluiLT
9aQ83dHCbn32A76mQAz6Lf0dL5Puxxw9o7fa6ItmMB9Vlq5YGDfENTPnFq2ojZwy1uBcJLOyq/Yk
zigz0ZmA21tSf+LlYC8lsg7hmZ2VVHsChhIszz53DoALLsl4Sz3rGqGep2BdqFkRQDFO9sMRbQ/j
WGVnQoIKkeHwFAqqMxqq7Ma+GXYn11oN4KMJnCh3xGyKIX/AGTVoep31YKzNsGqZryzS+u59B29x
fymc1J7+XjWF6hcvKooQc1qUNEyvssNsapIRaMZQnGiBXprlJfdkf7pxkUDOzyI83TRgq21PGHtj
GxGPr6Pc5H2ahmgJbdSUZ0T6o1VZA0V6Fsfd+I2OffYoez4mO5+6gQBCM7w4OtKuAkjt9u9s8hn9
Qk1f4idNVsqQOtj9C68gM2u5do4N3xXNoRE4h5lFctvDc/Fg/V4u8dvKKQCucNho0zAzyUwgVtjW
p2JUqQeCJsi/vJPj4fGhDKRvws1sDMWj31GO1abq5Ms/IoGmyjfQxyMOF0zCF3a+liBwpN/OmFtu
aMTlp05SsDHHtlEsBmNpz9Rrlprb8cg0zrySWtROpl851ylZA32nHiz3MjSbHsKcxbsjJGZ+34UB
2enUVAld8cr0jazwH23WiLXsm3j0IfRaDCCP47hbBnOfxNZb0GmV0FZNsXV3JXqs9Hks9sotP1XO
kIzr3eFynIadkM+Xuk9o6WAQzpb9qnLnpBcJ2Px+e3A6MzQxHT5DXzUBjqLJaTPXuV+ZYyVxhG/X
Tp6XQy3oBfFe0pDq0hjGKRZw8wj8Mj1R6kqL9PbPJGObRlM7x2+tzYOeMIrO8F4sWx7i/8ZLrVlx
1gDMqqA4mixveTULQLNUbZ+VFdj2obg4tawuXPBQw3cSL+acTlJl5+HM0w6jp1/tUjYaev7Kukb6
LNFEcp7HDHwkznmLSONpmv2bT0UdmgnRMUZR7BHRwyjfcNSMIDDtmQoksgZRDoA4H3LeGNYKKGz8
vcbBJXZnuoJNQrSZ4ta844B4OuSiRXZGS2yJz8DH249XFQIjGq3xIyy+Z/zBbDyi8K6+VhdcTT16
c+XHXg4gaI0khJjt4bcV7eOzhFhAPFsaVd6pMRXgjSvuSKdMJDpD+M4ce6ODFOb6yhUaZKDNp0UZ
WRomZZ3PLTPtzLMbruZO3vCev0A2WZGNq3mWaAy82opvl2PLxaah3q4NkQ/tw1UMz5RP3mCpqbtr
YggsVbojoaOSxdLGs9HmrkjUCx9Bv88rrigoUOPZQd5YphOuJKcXVp5+mwlzhWPOfgTb4iDowSJ+
0bLTL33JG0aScr1DG16WgWTaxhZyJKO1rWwCU1uE/UoJzpwn7okBA+Bjph0FkIi+Wqpyll9zTWNg
S3C/d3cRNNlsjCO3SNfWzv42cQ6CisNtbVVW3UsfeyzWHimgg046wllP1a2K0l+HNg8f2M8sm95/
tmckCAHPzTQjr/fABi/8acdG6qldLrZ0ncf/uMhOVQnkG1M1ofq/cdtjp8RQkx/L6JZxfPXbKNOx
2mo7nJJHQU74hwHYSnq7l+Y/bUBbyNkngSMjM/B2kwwcxA4e3+UqTfOI7117DAlWtlWAKdxhD834
WD4tQJltHJ479OM0qFpRkZGOfluHluBPS/PWCcCwpvx2Xa0CWFj+qKRi19WiiG+q246pS2j/M/fM
rLp2loJA3BJA4lYmCtRfEZzVZ+YHFcuenZwHj51pXTj+JW/5PH9KsVfIbKllxYt+eUDmC7GfZCFS
RMq8+C+tul9AeUvRfG9eHvhC/+glk6k1QKDgiib9gXJv5oZaBiHIZpfYMln7I9yobQugtvtfz4q6
J231XrgWL5MJqoUUBqVgMIfWLOeq5SzlVjrJvbQhZBIX9LZbfIXcjFnAtpJWvgIZDK9DVnyQ4Can
MpbdmW2I8YFnwp1w5x9Op2MEe3m9K1ElCbhCsW1ZqIllqkPjkYsB7VpiVQKGilneZ0DGrKtYvIjf
K+zkoQL/h6OLvJcsPoC+SrUeQmQAQ1kk0+rwYIUle9zWAhw0zaaRgjnM4Y5WmWgCcCX8gj8k10Eh
SUDnlmS9gGNSu2FAZ/LOGPI9/pG7T9MjLmgFlCK2BQb27sH7x7f7yftOCen74gSR08nCLZh7uUl/
d2H3DgAwH9L+mgah/VZFIotbnbdbOSptj2an3xaclFLglQL7KJNzgtQRFg37rbRiZ73dTypJKvz6
cSWnkB/5TdWw5FzQHiPboux2GnX2JFzZXFPIPZ4qZEGWkegfi9OHS6uyb82tuDmHolqBtk8zU3a+
9R0awY8qwebGecmMnNeGLVHLEC1JSig/IcIoYZSR1Y6WqyDA+ayhedQlDVEnHOiEq1ryaUKiAVwr
rByEQ/m6lNhmio8HTROqFU9LVGlCjk+pE2lA98cCQyWuEkqN+OcNZIPyzDC1w/6B2NRpe7Y7cfNv
/oATuPD+XoBO++7AxI9wDC/5tAjguXgVZrzFX7j1RDSqQXYyML3VwM6emXmnKasrVTIi7HWc1cUX
s9LlKGeRhwlOg/pzxNiR8VULpy98soccHl4d2w40Uuh7zShBHJyZ84tjAJ1zrnujfrTH4QITSq4V
Cz6cXhUnmXJ+oU8VOdGK1a/RdO0euWjsigrxz2F2vjB+zL/AzUeREAqeWET36J5o79NVlF8b5LZC
mo0NbCO4RU7VMKNpoUhTI4Oc5v/+hNmQGy+7xoxsNrTtcknnNwM4aJMXyDt3RygPs7vagH91J7Cw
gRYwHs0XLZQ4UpVny+R+cOMrviNn2ge7IhTeMdmXuZJGLSia1BDLpuk8wiLGp5gDhjNQXYtH/GKV
RwXuPC56FIm3g3laFcQWRvh2r5rCSElfZgGpu8rj41RHAryFk2mO7xb94RKdWW4DmkOCiwG6Jd5T
tVTRj9bIGcqnI3sBmGXwd8zUyED3C6cXZbCgt33VBMmMhFsFjgTiGTiaVbP1vUvFI1liLxrmMZn1
H/vL53C1IZMuFAK0ySJUXM/oF3msA2TIHTnVpqiP0BWApswly7PlfTujZ1ctK54KmBkcrVv7GANr
ZiTqFMr6YxVEmks45ug5PSRLIAUj4nZuGZ4FAtLoNlZxoOlH9VNQPb9+KUgFBlNBeLqAqHKQ4uOD
nToeWwnN6RFTq3RN85JaeyI1vKH9VlB9EAh9iN4O5d1iiUMZFnCbNId189lhhy42wOEJDprmYg48
jnH7dXZs+9yezdFW5sTTgbukGovyqkkpKv4d5XV6Fa7f3xq3JoOWDmcX35FalS+MWtlIxVRBUMNe
F2xEdzp97K2M6/tbDkV3kH8OmJdU8FpB58EKPIx9Sudh+aMCdTOGp7vU1Lt1jlRSWHGsbF5EFim/
x1emID+65Gg71JZbyZaTOtVsdayIkgsfaalLTOqq+sbPssaEuLR79bAJsaua6lZlX7DL23o2muVp
A0yKPzkLk+IXy1opqYtrMRZhhMjNIPJxehqdfjbyYOLmfXlE2KdElNwTLcXGS3jUNNZ0WSHebLbZ
znX1wSoaHaFb4/Cs2WkpwUx0p6jBNSi+VVmR6eDR0rBYZLnMn8I13hNiTxGyAQoeyR9KV1CC8hDb
oKOTRGQbX2RxrsN363hojMeQrz/zQKakzsJ4pJsi1IWeYKshnIJHxFKIOkoatuVGKR5QvIiZLA7W
FOcQGtlxeTf/ruhiUm8h99FT6l+94xjvUNS6ScDz1/AgCf3mHDKhCGdaZMK59Whwa30YyRdYIl2+
c2lQ41wblYtIj25nmqsqzRNopeawJA7ahfocBBCppvRHuvs2chtq0juvXH3RxMDAwFWcR226pBBJ
fp3pbKNLE6LG6ftlGjt4kJdrU7J0f7B+3SJpyO5eeeUStkKXflBp0kPed+aDW2O4MnApEwptq6ns
X0zxsotA57OuJVsQlfDa4jo/9l6gOO+xaWmYMw18MDCuxVx7uBHD22S/nt+tUe37bgplQafvxWzd
+czQytwYZU5FM/rkW3EEqEuLSe6c5K70a2zZiTK2YBIa31e45bWGx9nN/u/vFgjm3mQopvEZaqVL
YtbZfwnCkjdBipCgw3YDefgCL8OxRQzi+SWl8fADc3L871Xlzxb/eA37BKp3HpcClNX3AKX+kg9f
dxJZZOscPDBYjLsR/a03/Lc/ubZdAKHlx5pe+JLANdwyuWIAD5eow/1atNmUJFncealRgEO+8z4X
MsI43BSJPOeIAOiXkTkzQncglGS4SIFmgKQiyjZOUMTmiqi/0510mP6mq5HK1FJpxocdDR22GWNc
PgTOdQR2eze5ZQxm8N6PTXCwXcnNe/Ihpu/RUsRu0jeCpxIRKSJVO7K6rE+4BKnXF3lh6ci9AClD
hd+ky7NdySULY9y06tsuidgQfvTTKLw/5+Q2TP4O0iXPIXBxL4jyzx/7uF+AGeDusiWWIhAJ/Sj3
7Idx+pnnsNYQsuK4nfLj5nLjvnD4eErD/r75h4r1maeRzxIGAMRNYb9Bu8OzQdpIrezZ4RryclO+
2v1OSIqMeRoisYoBr6V9QsJdWZVcvfV5/sMeIK95fVAFe5oAXYcvoi/vCLG7esu6OurisAN/vjzq
liZNzL+VZAt3nxEnA3ZV0eKHK5X2rbqptTCfx8JqPaU1fisXgkaHmwcGgYOPYbo41PlTQX+Fjuhh
l+x05lhICTe4d04lRzoyXCgZlBpfl2UJA0wJzSlB5cl3Z9QZK7Mm5b0eQ3Tz7Vh6R2RDbNhH4cvc
J342JrwIPrRu6AMIC05y/tnv8iAgSQ8xJiTN7WoMG0OtWe54mr16o/BAzZ1909JWofYfKQT/hZdU
Hfe5VT8kDUbfQac22qU3oBCKJXxMBmDQ3YK6BHggD4jiUUsX0BDMlc81mDXFebDL8x/02rfkqpVM
4eXhC+kFBEm0icUXXpj/1B4bqwVpCnAZijvbzPtnm9WjXom9S580ZJPRcLpCH72A4TFbV8tVff7B
hoVBDfiqNT0t+f4M4HaQaNjQ43WYxOYQaur7TKXXexFQ+ZMQMVBa/CWrdE6cXzYSC6e4A4y3KTKY
dnZNm2ZdCZvDBzKTYYXBWZDYDJNDIR9A6jAqeCrlIqioVE+SeoHX3PcZccoNk+CSw78DmVvdf5j9
7D9ixmazih15bShMyGKIsKR6nPsxCXKXklK6l8YqwUgw9VANZJWoxEWyG6CpjUrppeWcNFBjebPG
8Z/bnfSJvqMgb4MUWHrYxV8bbtjBgSpJe2RSFnCNs9ewmvtuI+wgyY9NmcW2DhMbGT2liFF9A7qt
aWWm8Big7nWii1ORR1FWwg/W0xFyl9gXbcy8hp0pOcL9vSFdp+58bROrUDHk88wCcOGhg4wP3Y+Q
o56fuJgaEM4T1/SWFCOJeRuzgbcAWzdaNuZihjBz4TXGYt3xIvK9Gp9RrzsowMsaF7NPn8l6B+4N
XztlfkhUR0yEmywJGvkcG6hJy+kL6NZ7+iCrm1svJNlb7md9za6a8SexHGf2P2qgsfG0wrMzT8AC
eQHa57RqWAh+5kPQ3PL9UwZa7iAComHMNROTDTup8gzcaE1miEKcDgBTZXKAvrARqQbFiUkn/3ne
s8Qq7U4WW8hWHYFDC3iYpYCj5NOO24DJjyy7R6ykLEcZpHvw5R07ypGBHtJ1x9lBECrGWpfRndRG
Ng7JPyMdTZoM+P1WLOZNZzfQJafO73LJVKDtiOJuaK5MvwqahoKd8Depfroo5z1PlsgMSd1YRRvG
ymcPX1RGXkfH+kwhibp3mbIcdWsxmZtMeSmoN7h31TI7kONNxfJ0GEgyJ7SSmV6HpZuFS6xekwDu
D+/fFyQDQj5wUEapUdK1SFAQMMttmT1vhbxQLU71sTZ/q8Hf1wnrx44BP7WcbabV7eU9HZ9H84Oy
lNUZyYEzHMYZr/yFc0t51wFvHpkfnqGb1+11cIaE9PMVQInAhMi79o/AV3b+hLDe5nusSbxHAPzT
qHNkIj1AJnssEYbwK16vdgEfokEFfc2H0gd7nPWqb/LD3EYSfLNAGCIB9wk0GQR800a0cLPYV2xd
Yl+p7a92Fg6uZ3CrjtSKTl0EZlH0g9QlxXHFr2f6zYbXON3RVWUtymh8y2iF/oXn0SvCblXk9mOd
Dir4meqNHsbQ3CJwWgavP7MBfPZfoj34L5egoVPeFoyr2XGMwh36YSuMgNmtGAy7P0H3MLW7hPHI
V841Q0b3IfJeQReS7KHx6jLZyXv80EaRyaIWOrLLSPsVkEbVzI5bL9TUvgYgGXYUjwj+jGgBmGZ6
QL1x3xYzWJowykHZQaY5Xjlh1WP55HwWdNSwr0Bp4TMLaDzatlVuceKqo4Cun1u7vPTQvdrJzKaq
vDOP8X+9Znx4PhMVZSl6fSuFXo3caiuVZpoB54mXdHo8lahIzMoLTYxdT3fBN+acrnOMNCgSO7s0
mT+cY53Dz79k04eH6Ero8jFnSQrv1qUmR7bole/7tJUtLSa2BVWRTWSidM0FEjYjwKlwmy29KGas
L9daVvxVCIYXSZFMwa5ZRt7bLRVNF6Q8co73yhg5Hy9pSB5vqjQlkIzmR9e6QKODSm2MTVPtikiT
5DdACU5kw+FlOFHz6LSuZcCvV9BP4tlekd5BZjli4juYgtgm4tSb7pn3TlQJNXlpryXYO2W5DQm4
wfg5+OcXLZqHFlclpAbYNB3hJwvuDRDtW5guN1wtYYQsT+Uea5dramzem84PSRg2D43QA9km1kCJ
J0mtniLtvPcK5FEqVdVmu3p3mtD1p/mk+sUG3meWDdUv8MylI3TkQYH5q99BfyJMtXisYymQV37+
odD/Pj/1Db2+ihKqMeNPa2LKdwXhRED7OJktRxmwS0Zj1O6poBx11xoyI7DlrhiqXa3NldJ1vXX1
yb7yDxwZbh+cWFhODFRk2RvfR4KoYU/BPIb+4SbOYx3P7jQAG6ilCPF+RwfK6YJRMRKaGBFOQQ8J
s/IPF98iDe/WEBo+C1BLq+BC4923DlBy0Ef9MEmysYY8eB7fxgXyuHfSMFu6iPIGmtHNlT/xIKtK
CcN3EGKg7AsIecpbfqL7eovTzJB4NdhXpzkLD1bdYrk0TEQmqeuLt+yuIO/aJyessHYS/avoE+Ml
npQliSCUl/bgCfPqMy0v+ll7Caj5DVTNaXl2PnFlTdUPmNmSZxE7aRoWim0ElE0dWVsO+tSpqjf3
cYRc2J8XpRDRDux8haaNPxLxu7Xup3M6jBw52OxdTBJ3ZfnqOULRFtlaFJa+PxK0ctHGzMjJqlLv
KLWalFITQdnHpooDRXxCslYKHb1Ydz5iaYcpZ14VDk9+yjMgoyiplK15K4/jz1WBWjDHJkuzEBxy
4pYoOlCal6kHFoQjIlUoWyrmHbYlYfO5kc4Q3k1OIAE1s0j1rh0XKLiv6yXSK5feKMs+KWf0KEU8
MLo3L3ldWYM+/xKE461Vv61znmPUPwPUJJyVYgvSx6d9QDw6tQ1W29Z4SsVMwLQW94wdLqrtjeQr
AuQsS8omYwHWx/FDF/8phFV/camYNn4l8bws3LR3DNcxIIalSXSE60nNhvYdBQhz9tLj9Gi3Cuxf
feB1c4qhOhhn2rfcXytn5bootooJKoxHmFeYS4c425RumSI1jJ2Eou/3qEyQ57LUOafGsghvyaW1
m3DtclYL7EO+3lXvb6oNbTvr/D/8jJ+9LJdVL+yP8sdAXnkon2A3FsyZbbJADgKczNncd2NIdX4L
mZE3UOWzmnn1wpJeecjTpBIWw3QkdQ/HLbCmZ4v+AB07nTZ4OBUaFQsE4frq6JZqjL3f9Mp1U8YE
HMAnBibElFnW/XdKnwac9b1HDMW+JFereSBsJdQS3Su+VwdkPad8t3dinj8KCJJXCiGn1dsKf0oO
mKqmMU0rt98V4USp+4fbgpxk73/oTskkMsIFbUVghd41S3WQxV49crVlk+IIy0NyboYVIVT21WtU
tD8Y5zJOzoBaGM+wdujTbJ5L/hwu5ZK7+kw//5+eNsPA3SC+LE2VtmLX1ng+NGx56rOR8xEptHFo
dEk9poX1k+7Q0hEF3525MOWpHoEo3OdmqSmSn5XU/WOmW1bm5xBZ9n5maQJyas3K9ig8GRxCa2fq
IBD3rKZPYm1RXBxPsMFnF2VDRmy/bLNF/tM3IkLwh9EGp1054O7yCwQ7Ccsrsnt++641BakgOPS5
1Vnd1HQB9EX2qIJRP/Dx5g+LJH39soZmlDMSVcIH4URXipSJhkwnnBem3vyxj7AGQqspNlkw3J9h
Aax1O3JhCm8Gj6N6i0fYrhKdTeAAIooncmnf3C/LsWMWNoFL7yywIQj5tG8GZpD+1nd5w5WnPANE
aiFX0HXzg76FwyuVPBNUjcRMpLXVHbhjhjQK9D0RXAEDLAnMOQTWC5wU/Rnm9ykKc0yTpm1DCzLD
/gGUTc2c5+3hyw0E181Lb66PyBQ1LOgpjrsonxVD+9bY66hGgdqeop9lItO4kDxrGjAlO4cKbQ2R
u6oZBRUuXucpwZedfwBv3OMhl2s+1CxIXn/5JJ3Jsin2haaChYJKNpkuUShERIV3cIHg4zqNxMYA
aoqV177WcwFU00JBUVy+KDM2OafjrG8QcN9v6TcrwmPBURAgLTpKcm+3IIDBALb2dStmefkQcxQr
zetfLzRRRQuBwInO9tPj7GC4i49UF3V/WktieJufWo80I72Z566L0XsQ6fKO5AuSoF7ttZQz2n1p
JqsvIYWQ/2U0gt5lozs6FwZ1OabIdiX4TAgr5SwkqX1ORQJfV5h7YZi7ArmFwKbVlT41+3fZ47EB
rCyvf2K3doOg3sGWKKrWdkdr/5KpGSomKlBpWi/Y/3jNR0W4dFIVA5zGYHmJ/2IhxrXqgLHBQ3Oa
2vLCzuuBzkpexqPqW4JQ4cNC0/M1UZvvY9BwloHVSuWR8lPI4Wo3bkUaDZUjdP/36QyS6f9Nn12Q
1Kv+JNYxIjFT909SG80o5wIueVkxCh8npEVL5zLG9VC/UYHdG+Eygm47oFcHStCY2t8AYgEI3pMQ
+bgMrR3aStbpXcgK5gVR/DOEFk2M/KcIRzpiz358Ytj/X0YWsO4cXk7HNf5Yc3Rhc7yEfdJqP1oK
oe/8cR+or6LveGxDHK8dwCjql58HrBHebF3wO69rS8i8Lw44rEZbNGNzlvxYgTs2TcP8gi1bp1St
15ZaVMOLectQvLE04SWmjoMjqFCZE2f1GP/NW3yaWQksCkZwHT0WDC3AoZfQpN7oj4rFjZEEbnOb
mmLXDM2ww6gmdQ3JdU36OF8yVl/wyLS2POZltUF5DgSNVO7UzesEJQCSfuET2ot24TMEvM95/GyD
eIDc3pAnWEArY+esD9nAeDKiSNcImDlXa+Qde36znz1btkanwYwiqbvbUwwDPGTUJvxLYg8+x4Ft
nt//nYUVcn4aBkaSW6rS/GGy5toStBg1MqvIxGQ+ozni0oaBXVLfHcHpIbUwWVoyvr//NtgCd7v7
srcYHMLgvARFUjfovebWpItqtnjek3AVp0lDj2oT56tzIiMHHzNGH1EW6zpZtvmSUONDm6b67Jf7
p+Up1omiM/Skn1WEFV13YO/jkvK7auxIg1/BIFuSLh02baUfnsNkwzoHxOqqZJq59s0FPofPI7iQ
4/i19OKNAKOqYhdhDikVhc3oVFUiZdX8rPqbtC0pAkzIAxyFbHefTeOsfls96ZKdn8a0+10oAIRz
HtDLrl5QHVHQb6cp6QUJwnMDQa7GDEUqkfVu0RTuJVzIqrKZAFqP/iDdKCSEp4hxcAx0gdgh4GgZ
+JpQ57d139vryog9m8HAZ9Gkha6W9wMwNZEdqD7LoDs4A1UJHI//EJKqkDBIZUiVFun+t6Alp16c
Jesm9pKzRo3TtWRdsSgYb088j+uQkRtIGDA2YqOZJwbg0UTgrjCZ7eaLkvRRbLSCqGiSJfPVbXeR
IBRhKVSaqTrS52HPl1OQPFeOa3979za8W7RVBAjdR4cTvFX53hn3K/Q/4ipFQfmUrGE+EGXMR2Lx
8z2ppsBFgczguYeHZ0oXp1CpPRNWLSi68mYL7+GDpKRR59MmDRoLBrPsaiL5FzeU9Ts589Ephmv5
Bjk9nMcyYexYTNuNctnMNyX0HHModbFnTj4LE7ArjOaOSZ18OCGNkBVogdGSIjnXMyAT1Zp186H1
SDVM57LoF+LY+ReTDNr3oQoLwpnIdu8xjgfKGAgy9U0ew7jACiNk/ZenRm9YQTyL7r56CQ8LxonP
6YMc5SOwomRw94wVRkQkHcWlWHLCm/sgACxYPuof76IojgoPbBl71M6QIuJje4OwIf2Qp2BK9tj4
pGE5lSu9kW/gUYoq5AKCDe7rsfzzinlz25dYkBfnMWls8UHePdhj/vB57Ook9DaGxAiiM/0gYLp4
Ct6CHCYHX7++rg0LDWNZJACq9jRZWFJgPpdSJt1C9okucRtnqip8UiIFiDvE9DDaboVkFEtGtfui
cXZwGJQQ/3tLp3TLlsdADJboQPVD/sYNF02biKU+BXF21OJiP8mAuHKWcmLaMuGb7WIzdjDuEXfE
7LpWyx2/LfyKLach+mysoHMoWE65XUPOCYzGrMVTcn+vgamTv3VRAqNJyjnerKZV/jhuq3RTniSq
7egrIcnGk5lOzxlto7maCgbQXM4+V3bPSSorKy0gTZ/L9oFDOpX1BG+h7aItSDKlFlhzDiXW+tvS
34uHRqLhpm/pjh8c3bgQHThnVlOBOY/M56edXqU7XN+HtaPAld86kVORXkjpybcrC3+rTuRB4ikB
ItV3qqJPv2FZe7j7FJuSbQV3G1UAL5XLwyDFMxcYeux1YqcOj9PX+a5zqsi7NXWEmTpJMk8vY/bs
GoYeVSPCDzup09JxVG2lqL65JJ7wShTSmqW2VWwHdOw9q3O2QX2kuzuLWn+yGEYrZXKQzqv61JNy
X9ppv9CHSqC5gvzCFWotcIEZGIWM7LMekHJ7HuK/Zp80+ecUbWQIqCOxyBl8fMSv4MSS1ZNB7TI3
Da/pojP/XYCXwoHHKTH/lKoueoewa8qKyHSftKqUXnH2lXuoHx5U7Y2xBZOdqJR9G8eT0hKOyVt/
rRwCCQeEb5mu4kbkDzRL+w4/wh4ALCXwYjN6xRqO9fsiUbPLqw8kuZrYYyT8baz6yC7lzPGAPqDw
kZDKSpzk5eFUoyitMRsjjTjxcRU49fdWLpKY4+BajNcd5C+lD4PysWpuXQ7u8Z3Pa93zD2N8LoJG
mhIpgpzcIf9WhkbWyGPfe7Gz3UvN6A307nYdYwMkEfSn09PRx++y6oZascE17v+n/tKNHTeGL7Bo
kbImDOyuEw8OkTi0z8S4ODFZLigU7GfIhIuqdhEFPIt5EfEqKSol2y81wwgCECD65Vsvy6rjPfqR
Vu6lc9VpBVf6Rm37/MDayDZ4JGihBgTLMviefeY2sWoBaw6df11ujZEMulo8kecYzPvxEswpiXwv
nK3YqjU16V1/y5JYrqq7//Do1jyHeDqyISxgea9R9O+CmO/QMWaYsCsNmLDBMG3u/cfaIM8FT4k3
vFj3iYIKLvMAlhD/oC9bKKRP/Cu6uaWqUhaQeX5HHgzbl8DOf+fSY+hSenduCUCc3l/oJK2+ly+T
PEii/3YqJBQzF/frr/1eXJDTYm1RoA6JyM1pmePztUai7wvDAInmdX/Q8ASMZe1/YM9OryFjG3pz
Szkeergx+txjPoRBQ8/PcHzkr0b8nm+ZvuCayPa79em6KJyxBeZi4d/cmpR1YvxArLfV0xNT0Q5Q
KYvUT64nrx6nRCbh799KvnnsptMV2jRCcPIsn7uTVh5+GU1uiiw17eJ1qNG0Vm6wxXcBcAJqvjTw
ZGHiUiZIcNKxf49RDxq8WdLzENkYTmh+pCJv6VEhAwaa8TujMpuUQPrRraAsQ38Vd4O0NEWZtSTP
oCvb5wNvrLyMkz4rhiGDj+MD8Ay1PXMLuIlu0z9Gbzxkyf3VN9S1RXRg4HHNw2ioT97B27pRhWmi
+6esHDoqgH21vSUKYMNuCSzn0Q/t5M2L9mHw57cCXbTbSskV5dNHof/DP94Zl9jjvdqfWbDSR/k4
+RmBWUjmzWd6GxVh/Bt+uLXqFLvHCHwFSiNt6xBXk1aud6etn2+3YXyS5WfT5l5oUJJUQxLtp4YB
sow0s8mqN5kxTRo035Dx20Ah6PhtHo+TUe/L9QVwwfThUS6sSIeDzm0KlPWUiRW/6Lx4iFbmfmMt
ShfHnwMvbqHGpqNScR0s0MLZ50rcB72z2kPOT/9N6hs6A3hpYDMoTpNsmMmOG1E9yTR94Y761gS+
pBACKdXNe9GSL3lURB1Y1RYLxnEbpL/WesjmAUXaN2sxHFFMHgFygwtWSzGU8Eb9kMBKA1P8bjMu
Pa9oChSGOhrDVdsguePucYs0MBKjAd6+CUaLFj8sqQNGwzG1BqXAlOz55eowint1WPaDxOqzbKdt
3hggPBJwqotH3cdEatmwME37/QElJ2GF65hgub5LyH6yxmpQRAyrrDFw3QHcLfzww0dIvsod3nK7
D+yiDJtTwU7VjS6oxMbfOBzvcpeFngnVU5RIH7OelggnEnz9jra5RB1wNrQBi0bZcQhL00ZrIcFK
wsZxpWdMFQmD3+0zB7GbTtzxywcjamQ35Luuu67cKh7MmF4MKu3MpqnIbaRu9tbjiiE8H8JrE482
vV0Wz6hPm9nKn053dEeIOfLf8xNylvBU1F8vYI/uJdg54Q7se2PbPsYr87x0Z8NTkt14G1QX0xVQ
shr+S8QNSJTmJlbzoy6GHneF4Zm7SAg6fBUYltGuyIeuLIUVaP+6MzWGjcx4R7pf4Qn6hl4UTwZz
nOmbJXjTFFoon6doFCPFTuPsWDNhCyMQhWxozErIgbTaAd8CYpFc2e7miMWwS3NOZHokM2xN5dY6
HKa8ibvdI+lbE7MHDsiCEmMo3Yy3E9QMKJXvBXfI0d6ieFOgMcmwVlquE7vkNnc8mkn4gkMuSd8J
8fDyZQdJzMMKxkH8P35c87aW++CKv0Ashk64ALUEluU2HrFhj4MyTPbh9nAM4kMq82vZCZIrcGG8
+qiJSRQZJlS2XZ71nkzUmeKaXTWGd1NqV1QoFQOrqZiVBS6UEnGKKM9R+od10Gfl2YjjVaU7Fr5W
Xe+QskP9EfNchRk6D6T1KccadVuXcwLcKRmMiEP6Fq6bHqxfp2YFJtz+em5fBm8/K5BxFK3FUyvJ
XBcXQfGvfumPUEdeRoVKG7rfVCpxqFnnvN0ravsxRI0m9i/rpdbkFPHXQD0gzK9TVXVcVLCEqFT2
EWcVLjatXBy+Qz5r7G+hzXS7qQs5S1nuE5jp8quTnUe3iK4dKXuH9VTg57ROznBpn4mLht8/aU8w
XOOzpp9eCGeAb3JDAPVBNs7V+Vo35jG0CKr8g824N9gvjPjgQgVXHXj/uXRsCglDM8GmDqLJ6//h
m4CLpsgT6ww5fwwcdH2pv1dp36d9jNSsdGNgJ81E6Ip5wOMNB4CTfEAc/bqQxtacIBq9QMuVYSlU
mooVzA4WclQy+wpwbQ2Vn7I2uUNt4I8lwv4+t4XMVk2gHPhRLTHmulJ1Q7j761RRnI9cwU86nZG2
NXxzV5jvcBhp7YU2ts7wiSsPUZIChjIxNBm5ZYQymtIDjvKVwIH5oeU8HsLjZ5SRmXJ3+j7Uuj5I
whzc6yMdTggV7BrZjA0xhGYtfdjS0Fr9mDOPYi1vcu9LTldy8iUAZNlOInQc2my+h3fWieNEaa5I
Lks13QldScvYmx/mCS43Z6g4jVtvUIMk2WOT/BibIAZuGAMLNRUryL/FJdofYcZ8D8DvEizc8IMJ
spHsNNuC5kFLn2+n6QW9E3xzmQtQB2oRmdpBOuDiyobv5Aai/KgPt+AUpe/B0ol/1BHLiUkUwo9E
jcdJiLbgP+gAz/n7OmPOLG8v3kGn7WeR8NOANuDII/UsmO2OcmntwdorV+N87BCS4L+lBhOhsye6
nYk1uDGDCCl+Kzjrxf0uP5RPVdDqZ4UPT3RgeHtsH7XQhVWrSV1XFZfjpj0MfCTBBLK9p0hFEexe
ePCIeHmaF4w9i0AgSI+Ntz+BOzmngy73AGopOAvXivgbs8AWjcK5zo0TplAVctzKBzY+9slAZZc5
E5e2Bbxyix5kYd2ZUDGvS8wXX5PEetaEMcHvpgtk3AzOdQfijGI+C7bbXCYbSRWSp/FT7AvNTSV3
5Ww12Ws2FXurF6dLgy7feRLAuUNd/jyF6KX5ZfCSMdpfBrX/G5A/Ai02f2LoG3Q4GLXOpJnkm7TL
6sWiYMBxXGJiDkTsAqozJs+GpXun+sh1Wcz9O6+9ZoS/GC75tHCvGbmL9+j0s1hv5Xql7W9gS3yy
qdbVyHq0O/7PVm+FAQwW5FTCK780mqNHown6Ol7z0vN0/sZL6FS3E8g5Nu2ymGjca55Bvs00UTtx
iIpsyOajdaGyF4qNDX4DerLXHfVsbN7NotxRT18N7Ivhkbd8fwOXtG45RWEgbk5pKpfa4QnRYiAN
nNHTmDA/Qo85F+Wx/l6FQbCaQgFbRZjlvE2jY0TFInIg+uDsg0QmbGZRw+302h8od79nBVKX9bk7
kVyUao31l63s2i2SNw+jdHMj+h5HwlsRc/WmrIsTb9rlzfxFzOBTRtddpoohHn2It0lfLFWNx8ym
fQvww8Nw171x85TjxzlC/WCKD2JU5nWY69ISs+MuRBQPPGdOJf52rXwzNTm2EzSSI9IPmu0/eBZN
qHWKL1MszA7vlxD9gMmPpaUaml1iQgjuipHxM4BVWbBgKMHRwrTaI7ZkYD66PPL8jnZYqd9TN1z0
s8ziQ1gui/fbjT8YIF3OGxAOFjxcOXvoxyz4IVn8R2JN/K+lVgMgR1lGHt0vYgd+oY148D+Mth/A
0SJtvKIHaBfJAfoOJ/obu1sxKFSZ0Cfdewqjwv5OzQ4TGdkO8tm5pEhGYgKX+7V3fhDu44kvF+eh
PWT272g+Pu5IUTD1gMT5R6bSXiSekeH9sZby7gE0ymTkRGs24BnvAZ50ShQO7ocdd6+zBplFMnpd
ybYCuOKZ9jHTxAp5rbWML69DS2QkgK8LLCcApOdHVLh3DIUd4Ta9e8oNC79uWby8FdIL2Exd9A95
LZW3sDYLy+iDvvRqCuzqNcjyUcbJiQXj3RM9NQ3e7GR7p52g9oec1tKHSnGIP9JHqbh5oBTF52GI
hIYnUWjnXGjC6+7pOd/VDY/CaX/D1PoCGwse6SvepJEPde9B/lUYLU1n1ojewZ28JUbuaMk1uP7T
tIFU52+/+vcgQ5IrlZtda30/0FDJiRuE6o59Ygf2oqsnzzJM/9xzvP7/iK8X2ZXsoLRai01/fZSe
GGs3kFtJ+VVYXnMvdBiPmA6pQxbYefwg29OjlwOueFrAMGl22hoEHP6YiJNpkEB3P39vy1yq8FTJ
BIEA0+/dz8HZj/Fjpd0p8HOL+WvfBJznSa4sn1ui6yE090g6UAYdW/pX9Zqp1tC0JIvb8ZtI5XnG
SQ0RDzCaHNJWqIZi7mpVLbWIF/cc3dLR0S83wedXF81R+T9c1xVIXUrD0qlUy+EmUdHqmWbHDB9m
AGXdhhgqZkx1bgEa8SZ6hnVXcmbOqPemQ1s3rx8gtuhpO93D9lL10aTfIdF0teorB5s924zDEfDO
m+haedEo5yY3AS+sEcdCafr5PkRADZ6C2MncpFC7ODqJACA2cKJAtHmbMsRNIra9k8Dmanof01mj
c2zp5FQzZfFAoShLbfRlfx6TOiZAZULranOsUYJEJNpOCbC5y+UVSWcbLL7Sfh8+97Or5Ognn5lD
WExvApy5unf5S7CZCxPjkWyRQdDMZxgrnZEwsEVw2xOwF/4B4TsmTMgScXHkjwzpnKyhRdqRtC/T
dYn/YkEDD30l7nE3YME9wzHSu2T0dBXMzPPadeHvKnSUcye5bQMNETNEK5njKKAjnuvytQyJVd0D
h26lzTrJxx8/kWVk1lWMEuLGO9qPi/xLzfs2mFlCZxlaBIXpy0dzLSjPCDzVtIR0/5bnz1UWOgPH
CC017pXIHCISv8Q9iKtoXqkf2rRJHRvA4t411r0qpwZpovQ6De5A+5wGK6QUQmUxxLJ23f9Y28XP
3Dij6e+8euR8+H+mTAv9XOAIJwye8B/vUdqN3/kdyT6FrQKGgt6lOuRvynK5ed2Eq8hM8gpnOF5K
Bhkbe8Avssl5JKwUjoHLm4d7RFXgA2Qj5o9eQPLxsE8SzQRHOvXtnuRPJMu2K+KOvFlNihISmmGt
zZT0ioSUNlXelZU3PwwjvhypWp/Jj25rBLLwOv+QcY5TDOfiJb0TJAuXw3W8kPSCqzvBLKTHQF4/
UefZBpcaak0Q+AqKstQOnzv+8WPW76zlVByExu0ws3sKn3xxOyPI5a23EtC/EdhfxIIMp9cjKPNC
ezbQUIxx5R14u0clnTbl+bKQCl1hrvyVlogq0cbV19/79CVewzMfh0O9QgutMriwibzt+k/LwHXi
HU6XdcQ/L2FGcRSVGg7M2cqbW86kG3bKVlyFtLSMHJPbs0x4ExyePwgGT+jJZ4jppxteSQ9LEj98
bPPtAmVGG86L2NamfhC623SBFrc1irorC5xpLdaMY0dPpnM7dXwI63dgKOHISYHWl/D9iKlEWJli
KCUaoYKsFy972jBF/WZgDKIvBKWdBtsSWBSur3JodrlG7oY1QZ4QPxKRxZblIGMmLD0gekmAD8aN
k2K0IPl2klNEdRu5EmLjG2Wn2kiq4APT6cX2Jq7mtiC7ZE/tRz6F8n66KM9H/NkaIjq4nV2x2eJe
xaLLQn2MHNf4ZRDAkRKLOK05dDn4AmQulo7KnYynm5MI9la5sOD+zLBBQLM5MTKH1KOppgyiFabl
N82jQoNW24tTsnX0yt6i0HGts5OiRonfWwh79hmF9I51sOVTtHzwLyyLpxv+zxdqi6xCXjM4fiEA
mWQGtKCdVxoDko8NRXrCKAZWTPoVHOFMkLaDgf+8VBuhB2ukWIz8H1BOAdKXZCZEzH9HR4UQIfaI
CHY5FpmrSL9TC6ZIyzHlINUq1grhspq3rd+sKbUC8kjd4KTkOoqpmOA1JPOI95P80yvX/8CMt3eH
gshRthTJEbX+J/sMX/yevomC+ZW3YldJLjYWJmQUQTVZO7jG4Bdbc10+iGLEgVwZHKyOFmOEHkni
oQK02CDeobt7FTfYq5rZzG6WBdP7U9sSgdm3GtpDtc+J9g2fEUbXB6+h/GSUVR/jb5r8TbsD0PPW
I61Zt7tdUhZAGQn6FLWBMUvmraWg3me73UHbjfjLTYCbhGwtGqpYh0TUmEr3nuSiT55YjKgF7Ar3
Ixg2yKBJ9xuagjyBy7ZQaL9Sso7JMKn+4nOn2+u4nDLk5b69LRXVFdviglOasn/WujuijcWkWxxo
QS7gbf85egO/2mXdWVki2Enx8Q3/i6QKv+SPnBmNDmV3NULVYLf7MC+puftQk86Sz0Pv7+gOj2Z5
SzckOgA+OiA4xhB8/yNTSj2uopCMunQSHt4DDegovUiTuPyxr+VEG4+LQ4CcDeQ6O9yFEdQDyNVt
bevEMwGYfkAiqXn+cBKWEEsAh/S/mtqx5LQ5hPX/kw51Pg+sVhuDsC225NeXjvvTdbjtjIiKS2Ia
QX7wWHNXbPO2yE6NCESV3lzOqfb/WakOhuCqJ8f5ehLeM5paMeymhk9A/xspaxdPUHzChTqh2vCA
uPD/nNVz6jnEUT4Y+vjZVTrMgrtGL6iqGeWxqsRIAB9hFprf1t8M8wv8MYMabO+XZaDYJC3+AEq4
fYuKrWeVMMDsGUGxAbV7mKBu0aT8nZUtirlq3qndH6Y6F62pZi9+23ShZ4lg3y/rBOLDiDd28QwY
uMgtc0KwWv2VBsPTQtNYs2sP3CVbcvwwMxweEmt4C+FH5RUl5QJij0Dm98o8N40eRDTzR0Y2k9Fe
E5C2OI7Ocu8i4CaupfBLq2GOapFKHnJj9ORJi9jz81B2hvGTASe1IzTbG4btTtOEYs5hJ9gG+ZPt
V8ziHGJblOmcGo+hno9iiv4vrflmEdhknopLjGgvGS2UMbnAmnu5AEXmvzniN/1XY+n6GWJu++9x
LYEjbVQ0PchPyAKfGHejQViNLU0mW6ljRb6OMPaV6RXAQCVhvzVhWniKlcCqy9sQ7IHbXUN7eWbM
B0z+aTR4V1aZ+ZoXKRQ19u+y4bIIruOs2B3Q1TZ3G+1kJ2hVPTjq12aaj1BffxyxnAzMMg6Eh4pA
W5d4QZM/Fn61Gy6fBoEc8LLuuV0+YUS3s9y7qNDAlv0e3JKiZgcsJGDouavN7hY5dPOHUvd53P84
P2RNU6eEOv+Iz6YMKQOa46MdUV6qRZbWv8ZOKYdBRUZdXyPNrhasSCTIwOEnzhNzJl4grY9ZfUSN
KaUlQYzbQt4YKzRkmz2oCjg434taEofQfC1/6/O13WfPMRJ3TqiyHH3Si5zadqkAOJoibQohajF6
cfQkh8Kill8Lto3aCYkiwd3hPI5VcmCjscxqUzjDysZn08P5UpubGNXJYjKGML6tss2DEWML48Ow
ucyJpntRueysKu7NmTM0KOmNTvOUPDpyk1FtuhHtfxjhbu5F+leARKnWmzIO61NDuSqsixl5TcC2
iOVMuYxMY6WQfg1rg6nwyRW5M6o/9E/IWmlK0PrXrE0x7etF077mRXoTGGzX/VVLJMw3u8ihKI+n
O+mpy702grsTwMuwVwbpBmN7h7aDHopAZf/aFOOeG9VL5h2oLAPx5KzxGPbnQGS1OyWWUL3tbzVb
S6UH9sVoU9soUwNvI2bf0Gk8GOS2RkxXvqvYgS6WX8mlx/Q+O6zIIOIuEYiGOOdf7S4P+OSzc5qA
zRN0S8eG/F7tJODadxpnEg2z8IumzJXGHreG6z5Hkr+YHLa7uUuFJt7GSzr5tifhu403vkmaltE6
7coLQ8NSXR0YGpWNbdefOd5S/fFlyp6WPz6DyEwhjaipB6rRiEqurNS3s0tfu5mtUtTcNhgLTXuh
L/exJgNqbQd+Cv2m+o7twhHyE6p8Pral5QUpPNr/ULzxkQ354CpmQBHoUI1Nb4iNAtDPBXx2lA66
nQB98XzFOfJVbbkNP6dV8/kelxnzQFy6FqMGbhE/uHOfrTEoaZfW44sr/sYXBDx19GDKZFRjWlT9
LUkRkWVh7I46HKTWx45Jtzp0znIEpn0I8pL8z/CauY89B0A8Jmk0uJirmdv3Yjg1eocJBD4bCbZB
W4DN/A5NT/Dg8f2nfr767beCA9Ko8H/jmODbghcPBy74Z+LAjMZ9iPj68pNyJkKR3cYPaSvxfKZ8
7xygU6/q9cOPTvnX7FxIIYDn72NJxxFxqXoCIu8kV1e5XqT781LFtCqKBdy1+MH6CG9AoN1X5/0m
tbi4jmBieQpThGwyn/kDeJ7nZIIg6wnhifjqSrYyaSc63LEEiEEfFV1u/ePAhigeHAzykhGxNRX0
m/kHVEyvlMgfPBCYZC8vPkK9OZGG36q3G9NfJjoLA0mFwmRPK0XjlCoeAPAA5U8Bdh2GcwSpeWX6
VZ2TD8crU6eelumirbYvTIwpOFAU2i32tQmKc2a+xen2FXdB34oi6ZSL6t495ZSr9mW78NEy2JGt
Z+U96OPnJ/yraZzQiU0t52GUJ0MoqTztNV6VAg2L+4n+I9U7h78NF9NBOLGm0nyk7ce7p/7wF+e7
SO3Cni22O9OzAqIkq2W9QgasGo27JEP6lTr1Qh1JXRGgH2tO4Y/DdGkCrCE1kwxa1vrEiPBUelQG
ss3qltu/pibz8LKLwP0G7pvimKM/zuolBdt127VYBnWZox7ciThXac5UK7PbSNB/syjh6sRwzZZn
A6W7B4wddXxcDbQ3W3dtpJoRYm9YCYDA+GYuIQda5q0/sPSmGWoDEWfMdSCz21v+YKhMVCHKfoM4
cB9FXRtDUmBYWNrsFDYmaZ6IYvEH7snhEIE6cIGSsvmqGKzvLZumJTmA1i0kQpxRL76WZ8FCZqUq
d5wiQVLShe3nQDlmcoT0FBIWf/iHjFTg4xOwEoILn1i/6+Lz7BOQkPJQh12Yxeq8Kc3ENelYDk5O
bmMTQZHZiF07fyGv0wrbmaFTt1jkt9Skci0fNrJjc/iz1PEVvWOfTA4oTqafk8BpxVyPF4dHYBZr
/NrMn3x654Lx7kr5gBNGEKw1K1YRHWHc7WNz7MC7fr5ovq2+A3MhxyB7lOf84J4GFoPH2WqkhwQz
juZa0Z10ox2bbmliJYzCB1U7HYkLV7APMV4FwlHp7tWnRNO6nh6psBYwoPvF3VSMkJE3X4I8I/D+
f6VHb3xHETVkRSfCUAqO4DT+Vv9AXCmf7abaLdMSDNXDGh3BYAj1Dp+3QcQDJQAoO2vhHqiTSgkn
ljgFsZDR4POJQG21JlNwu8Zy8roUYekJL7LR6iilYqS/lEodtuj93ENpEZ7iKYge/FhvgvQA4hJ6
Cz+LQrHgiQSdiqvJvib83u92zI1+Zbb7Hz9DnEemLrvXVj9+5MfA/V5pemGS8sQO2Hvd+UQilGTF
Lgl4ghJiqu3XiPGMPAMp3sylZyn9x026hY7tU5QRtIhM38UYXLISSQWgnw216Wbg1Y2Xx4ijk993
70Ii+ZSvC4ONn20/7BUG/qDIafB966rc7n4ku7Tf+wvkMMGYsTfvBp6MkHdTWfH88k5CPu2F1/V6
N4UhfmJbhBjv49T1so1X1QR+8NXXGr1jtcT6r+VIz34PrcgdOeIwT8M6ejd9LtkayYepNiDSPb7Y
mzZ1GTSW+OppAJyFDILUlJgnuT0gi0i4z0q+uzLrAGi6Hg/uVW/5LScY/WKf+MCN45z2yPWjnqic
cMZTNtcrKiyNxHaUhzxPMmFcTlHwmqyYgf+PQanZUhicelkjQvxokP4wLl0fLnpYx82VQZZGn2yM
HMwtM9vja3yrG/7mbtfLHAiHQmV+EDhPN+5RWhl1JMuRUZlMR09vLSylINAY00yEJ6sLOcuck7ug
S4zD21/vSJt4/m4MRJvrKogIBDckNjpq50zpt0r2bYV71FnF6JUTREKCgMTTRdUPaYDK8hgcB53G
fVWLzDvIooUTEp0AjMVargH6pn5ojHM9GLQG50ESDxo3rkBeuXN30AdZSWR6I0y181SA+aoLLA6F
5k4WKeXY0lx8qnCpFYwKtKPDhOSpF4BdSmeaaeDq5bqhaVt2y9p4Fd9zHXIFv8WW/QfYfqrZ7Qep
ea16/GYVNiuY+RAw/7Q7mNnaQbGEqG81yRPBxjAnQObvd5BoJEYdCaTB/JebU7b4GooedsE/7neS
d+jFGrP4EsT/yhYS79WQ1oNJWmcnjuIh1XIfNFCiJ0yLvuctac8TY1Rg17tRqCMGegIoCVOEks5O
J1wgBuw9lqFG9bX4hr1Xx/pWWTBUle+KqXFzPOSkziedojOST6z1eq2iRQ4MoOFQlnyTf96Xrc5p
SxO9Td8Cl2IZsQq+AtA+rtlkdv4ovy1s1teZTGahJz7h0ia00GzX5JeAfVk1y0TKMvsBQ4H/7A0U
NMtmW7oVAlhiS01Js4fNR/mrHXE0Ahzq5b9k/isxZndy5ljv7OXe1bJ0t4G0FEZ5NpXIIjynZFYi
hKgGw1bHKEeQNHnnHgnkrYpWsn/bSwMUsf/Qfu5gAzgSz2/88ab0hVk6L0DVOeJD192TtK59ovqY
vh1xei+YNWwv4a62NUMX021m99jXTUul/B2YjjmUOIeSTviGHwn7Am/zgQ3wVuuJRZx8gizdr6Lc
qSBmDXNfOTOpxFcoyI/K6Ttuvo7cstM88X9PpmvntC4wSDGqA6AgScNz/8xsXLhZPSCcVhXM8K31
L+No095iyS7QYE2wo0f8FgZaHn4nFoQ4lT1ZitmJqPu37T9XLVHLFU32GBI1WoKywM9Qf+eARi42
EPkcl7cfZlsV4JGoDu0mFlO7659mXBFZ6gLnf5JpWXf8KJOSkHYT5gVDDhZ6Z3wKIDwrxfj0/LKC
caBL74nfWXmRZk2Woda+E3EKmRsfhMQ/q3D8n9KYW8RK808pYSCZY3DOIaqYCdgHb7wy/tt72Un3
7B5oCe6M9RRhWw2ZIgK1mzhxrJh0fB4oST607DbzaDkHRL1fLF2vHTEkey2WRXE+R+4ot7Be801K
0d6xmzRG+q3rVmU+2QtqpfAUy1tHzgzfoOSVXNHaPTZi8lU//YYnlw2BKDYfFpCPV2NmcS4vkasS
0Pzp9Ue1v6lQrTV6GAOohEzjV1IjmyqUkc4qN+f1qyS27XoPt8SJFx11ep1CaMhtZo7bm/yoJrjd
CtvV1/tlfdad9sg40oFYN2UPmWDdGHgfC1zb1JJHmrNgZ6QGKjxr74d8lrV7ffha6Ii5aDEkGp01
lmqJ+tKzIhMsK77GTX3uJBF/9cNhOO/EbPwhucBculBFbcvEX1WL9Lf2BDrHgwLS2m35sCBlL1rM
Sikz9QqOtqWHmXB+HA5ecrrW41rX024VeKExnxQwiOn0DoyBiB4+ScgE4MZ/PTrdmcH9zWb05Os/
cEjuUinvTKv1i5O/Sdm/mvIMM4crYPxlkwFPFVW5nuUGGfq46olWqstB1Fp7f1Z8QBY7yNLiB9DW
RMWNIjhuw4ulnaonRQZ4nJl3p6tJXTmTQmK1cVpcyDeOD0ogRRmpTSnf1+sEb8hgFYYFaguvXsvU
6XnQe5BZHLuF+0aL8XUtHTPpl5sTiE89Nub6ofK8h31aQ1GTFyyYhbHdYqf9c/XAgOduF/ee0Jch
pKBDTXYDJohnvNMAxRK0SLn+k3PRuK2a21W88Zc5sAOlI3FQwclxaDbbc8kML6dvs9qVo+lRZYf4
vtmQFCTrGdx/o3tr+8VG2eESJIn0JBMicqqOk0zl/vnhm/81ZyRnyRoL2sQqzLdk6uK6Wytbau4f
UKgrkmIIVN1uQWdPX+w/GtRswCP7lvct3jMUQKKXhGLq5W8gCxJv/zt1qT66lb5PAshrA3GSV0vH
VMXfBDOmogmdA2SRo5vxu+B+Eppo90rcEedTJcipQtTffY6Y1uCSFkOH5PBF9YpvBmRfjCkX5d2l
47/JKyQFVZ2p0FavJ/GsOTC2lvGcl55UQ3ASLWVJLwThAgms9e79T/xxJzXnc0W1Xi8neBbpOqHM
IFXt/4UxLr+0ZHf4JfZ18bnoKtaC4dySRHK7Qg5MVBiHYFkJwwff1+GSVBO+gwN5D38OFt3lDVG+
GYjoeqfbKNXtVRwFV28jAefYc3kVAIGzuDPljkhthcsqO4iWW36zjtzpS37ZxfiCjIfVCAxLFOq4
jGwFIUe96y+fOE1k8cogwFlPlKGntBFipNYj97q/dAS/le0yM3BUL2tOeCCBV9dupkW1ptj3iTV0
LjAFdrxuFhBFm/FDxLYFq3IIx4JHXH3eSo5Zm+B2R1JwsUfC/R3rPNhSRowIl3g4MwWsOTAsVEka
8813XrE1xQHbdR70xdolKGSemhg4iiDpNEw/BAZd6FUVtwmL45bSral5pFEJiyl1Dsfj9TvR2SgS
lLttTyLGZ18uZ7wVuo3t0ASWXYEynRCQggx05MOiwaqbKAhdm7FItM5eTHi5br0OqvcgeuR+2h9N
54sxDtlHgsjbJiYHxR8fWM7xtIXC3bYw5UhV7RZmB5dEEVy6FiztI+AHDo/ZHJuatYUaXIX1lcLG
htxXbCC6k9QNiAZAQ/R41hFCyF6ojcEe2VGEU1mUUfMJUFIf6uwnXghXU8hV9phUd5zMH71TNBE+
O/r5PfQiNGW3NDs6Uq3YIvBN2SxSkGOZI6/Mvp+2qyqjhpHB+bYk2Lp7pCM1hMRBxpRh2aAq6Cp/
ws9TYmI5AZYBPUE6+ryGgVIhnDj09ksngDYmNoJCZZ5iN4Q+DeGJxQw+qr2WWmkITv2XYUl2r9Rh
SOO7bXx3Lw0vlck7zSGuhujNyB2w1K0EyFT/N598XlG8oxxei5b1mfaBkpNZwNoc6vEOEBIRxj12
iAFQEWe19+YscdeSamjcXc8sOvHsm2iq79ApnqjO3mqksN0VYKDDXGqH8tMKAbp7HEsIvx2WfQD+
2xoBryNMHRSlHGzxxhWqOucwy+B1BxdmpOejsAfsBogxg+pCsWencL/93PgPV4zfWwwcpWXKlzoJ
zhFWgU/IBK56ZpmoDmI8h7dWk7nkSilu+clRXuXCZbZ6KV6X6UkQFgj728il0YEDjcxWRLv4eKt2
qpxfFUpqKvOGJ1IzUJORP4EzxLwhaq2lvlJftMYavP40mr3XjGfn97MqLEDawg9n7Xt8ABzL4/11
jd9yW/GzYu/A5FGJmXwBSCkYRk2RW/QTxz5u499DqhT6OxNBrakEpPC1AUIReC3oF3czB+OOMVZs
0isBlEN0gi1c4+U6GHAmLb/7IXLfHnslzcxRyROEnR2GSEjBfFYgRVtZbI6Wuih79VYtHEG6QGQw
YuiQf7effyM9pxmvJJlI8K7pHTg17wX+oJx0UqbmI7Rm5n8S7818rSSXVPmVdpu78CoIssoDXZke
mc8c/iQQkjH7JANy13BOec90rwIVbrX5KlSZdfIjN+dXZTpH3N3lqdospyLHko13hhglYxlrCf9Q
V8j0YKyHFZZeULHlPI8QqEX/fUSX42Hsz1P7mzeA9Px5A4bh//lz7kWCt5BpOhMlCswP5JVZwOyz
Nh63WohDAnBN1FR2PW89pvbQnEDHP9Sau6TwWKi7UI9Bco1ltcagBRHjrAzHMLmERrcfv7a6wyFB
t0JIXs7sQPVJAglXtQ4LF4dYm0qA77IiHDMkD9FvfwLYM8cknyFmgjg8i14h8ZWJhTpcdyo978g/
ArGhIJv3wy0caq2wRE8Bs9G+fhfgk+OOm+AEpGStt1XD+YI5Doiv/TI0e0PqL6SKGH/A6bpg6zPg
o6Kf8bn7M0bVV7JN31G8yLeZaouRm3bFy98YzDo60pnM+UEyFGr5IeTtQ030jtWsgbMTn1sjMaFo
zWJ3aXtWKdOPqxHDgW4fkwl16K6S2WjGabcgyczqi6hqjODbuSlNvkmd2ofoYwA5YCS1pXCZYGHk
DurQlHH1CNEVnHb8Ev8NSb30ujN6rqbqr7qxfH+Yo4lTht3HGRN3kqaRkTPUVatwXq+UW0+kbDDl
RoChnDVqklFH/PhaH6cOz+51WusJxUts0HenVzb3nCdjj8ksl0IJSMyj3DKbWhS7LDHz1XwPq+TA
CE+k1tGqnlosLLOoWxw8YWbOG8ijSh8PehvHycTNURnNVzpkqwqJP/vEpNInESCLrr/YO2IhhLal
qlPT4HwW6V1vjVwmsE4JUN+7hsvo8OASN1SzkD1n+38qa57RUNbOs+TfGNkx7qdQ1fGUWsM38FcX
wRSQdBuQ8xIPHpXZ09inuHCxSeUYlX3Mn30YfZcjsrLvnzVQ1siU4GxuW4bFsCAb7C+2NRP0NLUU
4+epXzlTx1cJqNWMRVl1pdWKLv6GmlCe7P1B7mwUApHhTb076Gjid2ZeqOrQbwUJEvxDJd+DcWWU
6OxPBlRc8I4R+EwfPpvAnRZpS/NvyqyspzVOzFttby3wYUJL2sXWurNL3FgKxRhvMSBhANNrE2uV
CXo5aBFMlkd+Q/ZmDF2vOlUq3f3j+HMDVpFaT7PmoLbUA1UnN4+toXv29gW2AYo7nLSXDbglaAgy
P68i/PpHNJsEODXg0L5y4J9n14WrRyNjtuVsN7BlbNlVWCWsNZk8ljI581Zk4UG7tGQhawxiMNsH
zyjtF9kb3Cwk7ftQC+8nsEv6elyxs8gIiyeI3+h5ePeiTlTLr+h9v+Auwd6uJ/jonrGpvZWz+bV9
u6Nn//OrpJu4AYlZQt8g2KIgzwmgoHI+o1D/hBuRqBaIt6Yaf13+QbxotZ8BbYCOwy/mOb/W3cHF
nC3uv6/6ji63+YWmfXTewiQ4jOY5s/tuMjfnvcUFg0LyW+1mnJaRyshBUg/bOAITPK3P340EKl+Z
THbrYkYPmDJv9uoAZBeERfXuowzyKF02cqIEv56aHY2P5KdHzqKWtHcwEXvJtCglqUI2j3L6IvR4
UUU4dhKJdwpGdmqVrYwM2/Uy/rt7InsmrA1o/a5Rq7frLENgFbgvv8sp2z2G6iHXX8W3G1If2/tm
R3npOfGrh0HB51VOe2YodEA5OsWx4ZiQkJxrlhhEirvxDio/HPmdy5d20QEjXtYsBJDWcV7oCIG8
OwcFVxpWFZxRvALqxVJp0Zc4NpjaRo++0y4Kzm/sxEvgzhJsgdwUrAqIO/CZM/TjaZZpNiSeW7Fg
I8L2GFWFbNINLXKp33FEuYkc+ft+AierJOfUZMezY0X/+D8UaxeTl9NgZM2fjrQuWvyvjRLaU5Tv
zo2KgUIqfP4C30GLGeR8KfgBcMUJAb2rmTEgY49h7jV2m0ew74TD/rXA3JKehsMvyo83LdIaHxSB
8tIebsfjmSa00CM7xmu0+I95ZQsNMZ6vNNP5UZJkw8R17YYzjqs4/X6oDn4AJZ6CB7EfHb/uTvJC
d6/s2L1t+FVOHIhA+N/U9TWjrU8jfoR92FYbJJ2Mq49TeHSiUKiff+KNlt9LIeBvtPhMN+4fKtRt
8vU6rZ6KnWwv/Uovnbi0RkdhfAOHY0FBHZvbPkQu7kdUTHaaiMqOaRXD7UttFmR8s6YQaVLmjJBs
X4wAHO9unmTQm8RW/A4X79coXt1tfP0aFvP/40fPPQVkgDxXDJmnIpgLh4AJBM9oW0zoWDsMxMzv
rgKVijDPo9rn1ym1sAziWhwPHjSFWfYuvJIljh8knmINSR1Zj28S/HLhAXV8w+wFV/o21Hc9AIjZ
HlKFRQVfLJkjYaw7g6MCXB9VZ6+B8eRygW52VDWWxL/oaAaQQhRt6RxURhpgYyWPvepiRsh04hvd
cJQT8fugNgRQFKxf9NvdGVkhye1vdH/ggAB3zfOca/uL6fibnkTQq7euH48vLhruC5Y1XmEgm2tS
BuShV408EXRSGbzRtM7GljR4A3goc1m7xS8KBqpt0A6u3scNsgKZz7/r7iyT/+nJSOiadIJkHPpS
QAnSA9l4gJo//7H2zrw3/nE5hNGo9w0vLNk4JnfIjBHr1gM/waQA+W/WC8AKz0W1ebuJz9XB45M6
YKRSvy2eoRcv0CCKdaHLbsEGSvMSRQ8+PJASDjFxacZIF/0JD/CXb9XmfOmNwvEMw2RGl6E9IgJH
4b/t6KFaGH8W5+u29XFeCoS3UmOIFmsY183zMdQ4QdPeGyVRc7FthQgCzC0gRfwLFVlToqMFd8Q/
/4pT1z+UEkV9GLU6i+l/z8cPS2qfib3AeEQPoYdfFDcifAdEsmNutQtTUxr4GwU5cO7m0WahKshQ
fKhohoHWCMGyPf4mop1OCipLCDVfF3z+Ku4J/LTeZGQLkKtLRsedvyJifLBzZBE+vSNDvAXQxyLv
85GxT9aA0XLn5rpjPZCwJZ5UGhP4UIE1mXYbsLAGT3O9fnpb5uLA1o9yU45r2GUTo5ZBGRj2EO+v
agOEGfjmMZjFpbCzMQyw9DaKecCn+NHF0n4tnBBt17MXpOkHSxQcT9Gsq8Izq7zaRIPldDf5LcUM
u1mKhU9o7voO+GAsgHhNPSb9Gxa85R8kBOt27pHjEyC57iJA3WmN6CO/PnKPaCj6+Smyd3DXaSBp
h8hrBF/72BAQdbgS6xbANHUgCGONKqRmHsj93nzlrHCeQ6AkWUjA3X+K9cxW9yOwioD6IpaQrUAT
TbKkY15SczkoYhy2DYt50qkys6pwzkMFRqkMIovEcP6ADLKXZggvJokjFCs22VuKS1EFhoTaR/70
AJF4I1biyAsFOpiP5edyocmcZVsLJKh7Q4Bi6gO78Yw7lzsGtL6AUXOD4ViwGF1EuUaCnZRxYJYA
exQtV5MAZ5wKBSKihZjY1JuA8tcqJ2lHKkUaef58p42jhJw+txoxCJ2uWgrfSIpiV+eGLcFaKIPL
9T8tE/BUq4XgpV0wde7LY87GL6GLRNlKN5jhZKO3dRve9GZJ3sitRKIEyJky0/Xs4xYkLjhivZ70
j52telz4FeJ6ZZMr6+ZaUvXWh5TcRe22duF9KYijKBf6zx09wEPA/9g/o5DsTngVX91OazKDqUQn
mjfFzO1FApMxt818zJPQNpTNqCFQy5RaKQmONtaLLwU2b2XsNhm+7vlKu9nTEF6MTrOUvY7z/4WQ
V3hMF7iJ12whojzYxbrF6XAX2NCoo75EZhNrh8NNJzzBVTEzlRs831qj2qDqCkNCgdSAbiBAekvs
/cfOmzGk4U6N5WUZK7gPVlcFWCmrQnKAiQmkOWMQY8gcOcwXFBiij1FDF1BuwhNhv+uICCkwYlZn
cxRAuwWYYUvnl50qqAL4R4/ufWfCZUpWk4TcsjcE4+W59X6/w4vbVJ90mmmH3KQkzvAPGTmOHQt9
fssDMxVkySa0A3pEgzVYb8LF7swXgouS5noaU9OV4PZn3bJe8zvM43soAo915xVWkxPRXZjMZsiD
L3nJe+007UrdpITi3KpmYudOj8ntoeT+X+C46AlZwXyR7qkUQxq1ZotiILFJCXJXgMLbGpMaEXpc
Yi4vc9qKS35T8IWX1Khp05bcBoUrvgqHZPVG2PMembCA83f0dw3nMrhlFx6i9oT0U/evTKJwnZ/u
3d0KLlgR6d2Qmlwypn4d7A5kfaSe8OBOIdMg7AXNEVLpkjNcoTiWE8YPYD8XCM6xomStp33Ff52e
QfDcspkqeY4xty476NEKfq8b7QKPgm3YhfYLISF8BZv1xb/skwQKmlBfGh7aDqIdAwasCXC5GP/Z
YkZhHrDOx8FEDAyrlN9S5M0nlAmeSU822MDMkwJKtOKQLOWdJgw5z8u6QUxyKUpHXSzSVxh/CUNC
/ZCg3N14kVUB0KCY5fnqQdMtTRN6E525E0obuv2thEkKHLJu3aLg6zh0U31dTQqeDOsd7+6F4Z/g
Hngo03DcV9ypGmhHSlngxASWdky5baZc6Bo4fqmYprbfTDaK399U/Q66X94eUWz6dKkpbqmNiLmK
m+AmnztxvPk9gax8ZtCFnV6rYLzWRd3Gl/fSPZlUaqRYhVo6OpNIhzxdkSDvbg2Bcc2z7braCzOb
0y4uSGwZ0uuU+ymc2SlJBMBAzTtd0nawHj7OA914RlRN5TtsgFsUJ84b3cF/bjHL+7cfX+mv61yi
whWFubaruTUcUoyFVEmPso3Vbb+kQzvgedaopP1juCMKy1TBt51cnIZbML5OzFDShl83iGBz7Kx6
2q5JvagrvR1pQGV2suyScuI84Y0IPyG6GMfHKOCixrpkwcU6Y7numdAd1ztxYqOObwvE3QN516Ap
mSYzAeWbfKnK7qXvX1SrmVGsZdFzfeIuq/jJckUvn09Q9wXcGsDat+ptpQCRFRnQP+4eRZUlTKJ1
zuTQsTJz5hv58bNpL82RdCOalveJp9TrlRzkrA20Q6ar3iZ1A++WuHX9q03vAOi+5C5Vv9lP9w0X
M7S1Hrs8qcvHM53xku9BJ71lXLTIVqEZaCDd8ydMcptICVQ/NHIbcvmFEAsaL5PJV35v2LMZBvbu
jaU9UsmRVAbuoNck5a7cbTu5csdIis9D4sL3RzxFGuIzAWLFK9JuV6SN5misyeQ/B5LO1CqvzdBF
4e3F66mFaLr5QB+e9A9sNPoWPPI5WVxVEd1hlIc8aAh6TcG01bPILhQLzuvp6DKfAFheNqBT9Vt5
eQngYtq47LVinaZ0nf4pGeyeZqwQgD2XE0G1mYmUIusRUvwei4OWBVOYELMSrBnyMKFFnCenkyNb
ncRcFEt6myIL42kgD+GA04wKw5+Z1qJ4xcyo6Db9lS9IQ0gsbIBh+hQ1NMW8JCTDyatbgm6SNQNx
ugyA7XZxQNyaDgDBr8GksTxBSU2oew0hruCpEyb/qYKwjx1W5gawq7gofqN8l6u2Qh0zujD9pI/2
1x5vjHToJ+449MPfD+ERBTlcjMulobXnYLlUWs1DVrgB+1nyBbCAezCj+rNe6gT1hMyVs2wciNO8
bOaXmIbI5GSrE5FMmIU1pW4d2W1WqbTteAQPzzc7yfKkfCi4LpshWxkr63PGl6Jk1gytnB6mA4G5
lxhqM09yed0hL+vsb1mkfXksr6IW+ZprnDc0gHkrLUdcX6lapL7GhlM0Q3SEMy7U7kpZqSeoNS++
SjUz+eDRYHSNxoFY0C8pStbWU8DeB3+ecMJSthpLNo2BBqG9QjL9s3lqoBZAjHFXqJZWNhbqtUe9
lHAIsGcIpweJzPepAzYdPha8Zp8m/siBx1StXhm9Eg7K6TfreNCAGBIYvewhxBsvZAGr2UZL55sG
DB6Tob8p97pxS+EFY34pwGIwykX0AiER50PynpMMcgnZ4uJDtYlWoP54zsFEXTyuG0711fHD9Kib
3E/Wn93lZ27d8wcp6KJC9EbD9a0OKHEUuqrPCNiYP+hlnZ67ANLt06dSyROcSK2cnvFxXdMRulF5
lDQblT7aJNonBzcEyZDRtCHMH3DjvMm2/8E9BVs6zvOjLNMqS77USaIoxDDy7ZkZBrB0q52e63ZD
K5Zol6bJCvGYWDBPJ1IlBIfzP8D7AxPow96abZqTH1NfU2qykH6ik6sbg1FIpS8uCov7yRUyDYkt
NQ9uuROPt/DBT6D2y0O9NdImEqiBdqpNPBY83w0Y1jEbezs/zoxSh22Da5LSD+m1b+2A/wfWrYFa
i3GE+tGrNS+VTqymP4FuirtDLv5tv42lOw1Ui7YTmTmUHB+PCH4iaMatWNc26N+Mh+9LerUkF2Md
nJBCY0A7kPnJwq2sHThXZLct5pT0TQxidt/N7xInlZfEIdrGy9TrpIs5gtftoJswclu/uQt9ySrq
/hcOTMBnEyMOYpTETVlJ5QIba/rbIuRJzMmpqnVA92164wwlIVpGMf1fpHw1kdwwGiE2C3H+XyB1
C+wfzCseMmezMSxpG/Vb7c+6Ac9/P3uS2IUL2hQ1Y32SovRLGQ6xIz+IDq4bG7eqeHNB5KpVwYO3
eKV0JJHkqHwyQeHXyUHH6ucjlR9luPF+cRmDGOsDnhkp7k/F/sbiZVZhcy/gttA/mcf0Z66RIHBl
/Be8ydr+P1yw6dkUMOhKpY7yJzWDH9jGGRF4dAeTcMVgtWv8Q/gg9mVA4rOWyWvCc50R9cNaj4P2
bBrQPXmovfWwe93pOji6Txi9848g/MgdWeT3NB5K/74wLHXL0sZw5cm1ARokSDA2qPiw6cdSVFEE
KWMdY8nG27aLkzsbTbqYREgqKCVeDj35gfn1RNmMVhnLm9A8HuQFs2iMO+k3t/aW38Un0VHvil/6
NyKIkOqgiHgswx5ypxfhYN/FSQhxgiGVHfy75p5bA4egZNHYDAB5jfmpkeZ1HxiGwdxjg+3TKceb
5/ymh/KX85wkIj0xWnd6L5Bexe8apm1dblxpSRahTrFnglJmNw4axqv2SKCnIRiWNBTTHsBoxc31
1Es5HK3cWio26ZOYgp0+FbwyHyr+BaRRwHdWDviYEuw7VrFWCzVw8xvte2pCxHR8P6jPM9rZlWmi
6goDafHOL/nN16LwWx5wl7XMAAZdf03ikU5tQX8zVF56s6ABDlUu3C/klm4fzwRfy68yfYRc4L68
N+vAMCr05+aVHhxifSQhDOoifHgMpVo5gSjbzjeLDBATqmU9ZFVCTJJMw7Es51F+naZj2n0GFuh6
PRF31RQxzO74ZU21Zw34Pr1Fd6p7iNyTBPxS3+oMx3XCGarjwuj/7zMJTvc553DQLPNTu8kU184N
/qxRuReHaucgMXmlTY6NXbs+BEOwMrPlPRop6O5A4I3/JWdyy2sOVs8xM7/NksbYvN+U3KzF7SvK
qilxcVydbj1GgmvetEXPU29WUJy9BCCMM5lteVCn/EcXwgwWfk1ZqfL3RgzqX7IIiMLr3hn94jXC
n9InbMAmm6wvM4aZudsR80SoD1azVPaNYwNdtRq7xcvmnBVPWyze1BWgdv7fNmQyUMFd0pLa3Ge6
MZb7sIHW6ODMjLrLoj6jg9CrO8N2+MnqEROtIQw4P1jXmTjUz3N//5nIgnphxt+IYrJGvsKFDy6S
kijkU3kojI0UMhLY7vBtIm21/+j6cFm1msixK/++KqpVfJy95XmcX+dDpDQ2LJILg3tDYZXwziTk
IwMalQxP4rqOzWvtg+ouS2XazoLKbUt10TbpbelMSU7d4v61VDGkSatQQT4WOGxq9QPPkD27Il+F
FaaVA6m3e0U2ox9hGv6abGP/1cTJ8g16w6S7zQs9EL5dpfqw04iF9cQr2CBtuSf4YcCWrGHFt4oS
JPx/BSzrglTCGkkOELG5eTypafVvZHP9wxpxczNxqSAvkfCWH8zbbdX6a/206+uGWoK+KWbb/Xhi
L73zNo6jJvDh/Qoba3JGhb8B8/y45i7DH2g/mlumK6qbW6yQqJrM33bPquO2yTPDdUY7AhmBDzYS
9X+f8fxzBVHuaTYFD4KDRKAJXJcBlHnig5nCgbEYTp66B6TuV2sbvZdFT5hqHXq8uLdJS98PAGsx
oUx/KV1pjOaP9GoRcSQCDUgZgUVmyhnum16Vqhyn+bX7ByY5CCNHj6pVPuJEphM2T8+r/NuLWQOR
0CWbTuYHLY/De/iOsnMLJr0CxnJZsyctUirSU3yUk9ugMUYNGKINHMakTelUAnYBJcmLFTQIxM51
94Lj6xexzHjP7EZr7aR2qDBPveERAJaqew6UIAjwL3pJSDJN3I3DAm/w5sgGzbOl6fYN+/vmmUok
xgaJyPdLTMBGkfc6j++Q0WoFNvlgUGIYg+9LwoC8DYnzX2bPbdUvdBYv1VBLoZEQA5ycDmh10gjK
UZvnuTOKsDQXBAE15j02FCQe9UJoWm+ahwlxGzxl59iH8/4OThC/MtXkM5C0TSpgcmycRtrKG29s
mug+p9emGjTfjXgSX5SbQ2/2ac5uDREt7A8BfX8bhc9797xe3OPw6A+tMkF1MNMvq4RdsQ3jr08G
D/XAzM1+k2C+Kas6RtQoSGJZbxhKrJHrgJzRPPh0CY2uWnq2zIN/0fHJS8Coh1miO7Pj+1NLTfCs
sIozb7e5o0VyeNsXyTIjR4UDuRlb+xtg4BXpIChQ678YUziIfXNKo/dQGVsXXLNE8slfBqXcSHNb
JtxECRwjLWXLbWv78/9L2r4mFvGpnCt5gjmwe8ePKxtUqNcnPlRvnklGIETSMLwV1DaDWOnGA548
knYHf3sHe9qDnAb661hDjVm6X+7i/br3itTvcvyg1ATwX99lTrLDalwC11nRFGtQnu34DmDDVTLd
wRyg+sYepQzyXH0aaJ4IsYoP56UYxSVgLgtk+L7HIeEkMvEfbDNjlld4c6ABU/rmeQpsL5P/Le1V
3MJlD9pr0veVhhV7ustN2WbDT3/J7MHMa+GM1q/Kw8BU7luGszPta13JTQ7bNNR6zND1YW6xOvDL
+y0YnjtrGQzA6iPuY/FsCO/cGnbrNwzFKXD1pemEj/2BCbBuBuoed/Q7xCc3stB2mDPNcQEK3P72
S5oWuWKyc357YQP0XJ9gdL7OQLvesSSEY0dNHf39s8TEyCLWl6H5/geOhU0uxERtaMDbMlJe4iO/
0zVzkLWFBGhfHwmEV0CPPehLGTdvSOiH94BPvsjd95tLRLpWhN+WTHw+1nxEyRxEVmHajdpgTOE6
VMBfndG8PBpoZdviuWahBkFwovgbVuSFsN8SgrD1nThsYSECRmy22o4RKKrtqygO7QD6ZLu+aM81
b2KHi4jYe37t6pXlQsPHM8bMcwqdjfVKLwsF33CwylXdSDzTQDLKRnb0Us79ysahDxs73/1Epxl1
mx2hVha53SQX4qRm6zMxIDNsncKx5mhJA4hh0D61yeQwxg8My8B4xDKPEMSzToj3en4k/1pLEr/O
It/HIPkD53Fzmxqp5BLuTDl+nX9NOOlpA9CiW0eVKW/WUqUWcWu0GEhwmS6sOxFtrurPLO8bWizy
3/iPMUWU/V1usuFxjT/yZjhiCyXUWJQceDvru/HsprTifmGyaoMMbvR4Z6qkWdlgyQey0FEgkCsh
/v+hUeXVmPs523OiDHId8VrcXi+eCa1cadeuvsdHkSDvmAsruzCKb393Jw99qc627Jp9qgS1DPTx
9db2DRm9obFqrOFGFZMPV8xswn1JZf4XEWqBWEzCWvmyFvp6Odr0fwfpGAq1WYcM55fT4jhA7Lrj
P4r9s7e0lPsoSpiOVj6vGX05XG64mIAmDNCKlAyA6+SZmapZMmUQVPUcUK7K1h3BFXm2utemPnG+
+TNlDQIl13JYHlohftdK3CPYwhgeAqGOmoqKndRpcG0M1gtjcqzIOpKh0V8uv8X2gn2kmQOmrmKK
SB01J8qR5W0SJQFBZoeUhXHokkxGExu3iuwcBpCp9mpPO29MRzHphNO8AvezPvnKcZvCd+2U6LVR
cR4ch3aaPCU/Acjq2SrSVeh0mTQhyOad9ibiVhKCodJ2DY9DUvCfG/CRP0OYWXZbLt7VCYkPn/SG
nglSQXci+QYG1Y+nlTkwFM2Laf9Z065LZzNQ8xndfKelXeS2ClpHmQioWmk2L5rrgU6r1EW0sXzV
bNzQABiG8lbc2weUnPKUpoko2wAk8d1UtIbtJ7Eo0p93Pg6IOwb8XbsnWA5V6N+E+YRyuvb0pzzm
pR7qWPR7M+A4tFYgW86Uq+dFonDg4n5c7T7/H87poNzjkBVeJbGjiWok4i8y9UygiQ5nsABSDyCc
HfZoZmaLpVYAF9bodSDinXPbYKcMjL4E5APjVJ3xr35RqOcd2I/0qk4jrcVulhQI9xVLpl6eRXJc
pQV+BeZwz9FI2WKXBX6QcQDwqTSnhvIAutS5I8UHC+vFLxQAzokUKcoYZlVw9fh3OviE2mOMhb+e
L07odlbais2HtySTMxZHo0lmpHjKMX0Nf7x8QGYta9xELMzodeWpP0iSR03CXYNgCLTh1f1SMT2v
X8zND5RNQcqLxMPrAnHP5RSqTPutYJQPIvoDQWDHWg+AoCdlKHSauuoH7NAdqyWgs0HTI89ZP2xn
cP/mrU5ry3GWJgeuNRpAUZ/aadVlLK8O03PyB4YIq67iaX8ofZaUdPE/BzLdaNJQu3Air2eXmL+B
2q/PUr6xzWAeyCKWlmVgEp8loQOj3HUQrNgCudVcTEIHcSAxvNPHNSpq7N5+rhehu7ocHiQmCDdp
lKZboJtGqIn8+9Y+upvq0EXBa4ZX9ZQ9ifyL/qm8QIl8zVgpdzdQHYffRjfFWjaLVpiYYcb5vYgG
s5FPLPWaEdtatH7x4efeSMLUsF68a9nIQ0e28lCLaRiQb8oHCllMJnsrhs5l3EGjL4ciAlJ6sx4W
Fl2JbDDJANsZTD/i9Dj6fIjUmQ/wZQMpfw9Rj0KzJILqSCYvK9uLxSFV5AY/newThzceEXlMTMT9
wofeZqDlaC51xKQtCRSUhRokOjSRtVa5TLhnQwbVe2vS5ayW1lKIWdqB0GlyyPhVFMH8Oxo8ZeEA
fHUcG1Gyy9gRhz8gWTAGP2JJdvszn0/4cot59mrqNjLuJBqGg13VwDQP6/BPVE/+dhphNOMhK5L4
jXGgWsuLbZmc5aQpWB4/RquTDTxEFJ7HNVJUld4hmmCEucX4LYX5PFB/5cmGvDpJD4qjXTdaZyH7
jOuTFj9PU3WJP7y9bPxy9MNQxd3LFnrlD3hMj4HAVH735qVQAx3DvgPuzW422goXT2zOSwENboYQ
Uu3Txzv30/IpEgwDa8sb9Wy6hJsPXMiFW0VIDjFEMDHBkFKV7OT5f7kVoUsxNwbjrh59Bs3ZHklp
NuZSj2Jiw5vILFccSk0tFYmytuPILG9NJo/hVL95Tp68S1cwI6MOQ07L3n+fUml+7rLyZStpiBUV
WY6Blx0N0BqIlDSe8OEjWIi6n5gzLJ+1Z6Rkaf/s6lIrisVga7AWgnhMkSzXIrxBeJYA1BoSuX/H
HccDtXJnTjBXm2HSY+GYF1CVC2Pm5I7lU6iPoyU15TXAyKose2jk8LQ4xUXbvfk43daVS8BLVuQG
frTpfSqh2zXyoMMWKyG9PyresZh5OhWsr2+ig4aWNGgd3V4IUqIZpbyP4droTYKST3eeGFO+Z8+r
uxSEoEmm8/YF4FOknoWfQrFN5k3xYhlWNB6WYsya/LBTuqVFGTLeyEUJQ2YGR68hece6chddsZkn
5QwL2/CJXo5w7FgXZ/I6MRz1cwuY35mof4ZB5OBA9wyuMqDE4scgd9cBMU5Krh9fc8n9UC9GCdeW
iLfL2GDp9zZlsy00Y+OMA6x7x1fAwoL3z8Ifg6uU7VUTooN9mi4MD6A49AcYGGAyNweMv+OZcnHc
MtM00RuC/6zhQIscooQWcWObam+o35DqYhulkd/B8ZGq/UAg6h7V55ah9jT/z5FBowlwtCUW5fWX
ZJNQj9mLpLUhR0Rod6CA5TeNTokO4Ffc4AW316isyEVrX22xliMPNOzL2DMUXGowpMC28gYyq1H5
jmSG2XT1xsoQvdNgLa2g6XTmQTuoXpXCEPwTI29L6sE0Me1AzY4t8vMlIk74bDQOFD4MBAi7MJ6B
5Ddfpqkh3/6Gn/RmSOt4XIrNAhuIUaxOz+rEMtFwUIfW+1dy9st8YSK/bUm473CZy/qKtacMCq4k
8dDLN8xj2nniDivE0cbyQOV1J2Vhi+LoLbp/98HfEnFN4BxKL13Cu9IE9t7B/ReC4Y9yuTqZ9xlF
DeLr2xYPGhBsMiwWIikHjrDzRH579gVNplyx7emyp+B5kyqSPH9fAx2v/4XtNoi6A7YUMAnaG9Jn
Sr73uzmkYY4Wn0apzYOP8cIdXDl2WbIbNYTtwg6nWULcNLlsIbUljRXqQaG4rqX6iTeVUZ8yiQnT
P4dp5vETmBmUl/elG8VYY9dSJChTUb3ZOhuS2B43dsgHlDyDliIiFIHlwzCGnAr2zmJhedEZDd1g
+FEV73+9TR1kDZU2pDThQffpVV0sqiwrk8bUrV7hvUDCZSKryff6Z7w2Qjg3Zme9nDI9V+JpLNna
vSidQHmzs+ZRf/1vgvWqIZ7wVGzGc0wrKbWcGFTotijfRJXDXnkXxfSwOH4e8jjN4+7J5bikBZ4k
G0Id92yFqIIMtPFpdPstniein0NnPCBelV6pLWJgN8K1p1+xYFue8rORt/4mXPCNf2ojzBy1X/JL
M4MSOjjpn4AcGWrD6pRiXdIGHNlEMFKsUHPK3vSVxJEVohFxVK9VQpzm7fGmJUWxBoYBUE0QkjeH
6xCMtjZmZAe7wMZofhKXEpVRhU2UGqeNDs4JI6v4u44h4Cz/1owkS8f56p1BUnNRxp/YFEt8Rfku
aerLbUS6XFM16HGUVqQas6obUUCwvTbK/ekMXthT+UYz3a5hAnpCSmIsi1PNd3Ohiodd0fi+H678
bVG1fZDTfE9toZ/3TZaRRbPaCKT9hsrl8JI3lhQiYAcesBkpauxP4NJQ/WCQAYvDqYzuUx0UiJrK
QubqgOqLvSdP9pe5wn02gw1Heqozw21lDbu3NvEy1jpyg6REg7BPvxmhUQziLctOgITlkBGhKfvw
0K5f7YT6UDNnSMZehZN5GyG7sUUdHmBeMwk8PScszvwNM+6do+HL/TRo2w94RVUM1HZkwmJJbXVV
78Y+f56CTtQgH1m5EHge6ZrgjGTDEi7hYxCacv4sa3SLqxGI8w8BJ6C0oM7SaeBUMw/2SA2TCtt/
MEouhh/LFvgf8pnfooN4NxhG5URKJcqosNhKKetVuxOM2WFGcISx9L05O3CrGsngFKWOIetNBCpG
Upx6pxhSrgt0wj3axEfR9x6It4fz1C/Ka0UgumPX0mHJnlfVavyR7NhJgoaSH+R+GK4ik6BMFZhn
+W3dRVoKpvH0Rl+c7N4h1clqCCprnkDD8b3YiY+vOc2MGJysFq7k6Es+K6WJ8v0CqHiQPpKRQkgo
v8sv2mMzNYuot9VuDE7DdPl5N+czHsGyw52UGnKxyepX7pizSWGw0NQUsq9x+QyL/lGfjDUM67Q0
HwuVbGmsOwVBjpVzUhlDGf/wPvHqSKuediDB+1PIv57U8jonbDMKbpcP+ZKoGdwVJGFmkyT8s9zq
nPuOGDu5ips1WNHrwEMgwXU0Cveqsfi7GDvzlwa2BGTJn5JXvYMX7ux3Jbeq/BGIGAPcGsiNTyio
ByJBXXhPp6kJuM8DOw+KjT6JHporfDgsdcYgC2wWFisjkjFpSrEQQ1z/6xd++95ajL/6NfoE/frn
BkBYCTEq7osIiccP1we94pg46n9xtgJRXUZGQBdjMx4cSnu2divchEm//TNxLW9xDMe8mNPTznV8
PwPBS3aRMGbFBLCoMJ8fOK97niFqYkySu3OdjPn/yv3y0j8OhZq9jSWghZIgHMGCUuR8/j/SCn4b
RVqF3rq+3reZHMDZYrisNeFH1VHXqWihNX3Q3hsWyFpUtZDmbBwPw6o0KpazaOjRf1vKEYbkGBUP
eN54liu2pmvgsr8xysn9VE5XnkDIdQI1H10+H1VRq+/yZdxcwD0FzunjHDBrFKzATIMv7lF/wvg6
KbV5ATW/970RXeBdJvlHCwMCMx71v2lD38gmRsB87yE3qVHfcH0kZY0mB1lzyW+wIxtWAjehGmNy
0Nj+zP2TDTxBG767cZ3CrpXkshQMFVl42Y8Nso3P7X2Bh0563btD3d9UyM0Ivq/1KqBKbddFmFby
fIiQ3Xfma9kZ2M1+hZzF/piDn4NKu8KBXJGaH92pLKq33sMunV0UfiZ0lbh2nCkuOZ7LCiWDzMhw
9n2eeQoULznVOBEQKUeXcKtWlzC0abQpCkqW8+3jkbHeT/V7WrrLN2yKYB7J2nQvLL+nsqRJlKzw
7ys/r6/kZAmjZPjPRTRTBBSupnT1qAmENrlxzVqJB7krVATyAyT68O4IrQVNAn+EKKigGlDxzNRS
vvPTiLAa+SNSOFWNM0+ouAZ7S9gxXLTuBvIL/vjibkrQZOHRjHEsoDGtIMHG/A4I5cJ+v3IfwCYf
MBms0ITHDh96eAuQGEpi+OmoGY+alryLdolmUQiixeZYzF0bsWj6fkyRW2UgqDXDx6uWvkamME55
QWKXnv34EkbxpBsvmvGDuVw+H1fonI5jGj1Vl/xMgpM4xbYPAobErlDF1b/gQbN+DDj+bKSc/HyR
uKd+/ISyRykscrF9Rn0Lt+EI4b/QbJIaBh8FnXk+LDojKDaeSAEjt819C4B8Vz/sXf5aOfX5AhUw
MpEBQnDHotlYYNkxVDglWwkcaY3EK3Hd9qMjGDeNCUas0c1fWOLI75PuRk3xDCEAMxjFzVnqpNkH
Q8nj2VeRIL34lqHbJE94knAyWcHT2FiSNQqClyyePpakTGQjUM0prwifseeWCtwGB6EJ/eZZFrpS
ULHwfZpuiThH+PETSmpVsVpq8+qhJ3H8qPkgaJ7dDglr5pgitAH4xFqu671OCKkOGFG5AVuiJd5O
3Uq6PdvL358guciNhhySqQp3nQePA7aCGxcrVp/STyxwRuD1kOurFz3N02kWAn4A1YAkKTfdHdlu
BUj9UewUk9gkQBNGlKNjE5doK+mNZUS1C+fIy60gt+pXpQprkL2dJ0rwTZG+IHhjwVmD4bqcvMyS
zQJ0ltoh5HBiK9cs8thIhmDJ+s5+UIB5NajY6Ch9PKxjfnSQqwAbFO1nyUqvA0ctd4IfBTuySEbS
IE5x+O7pmub29aE4YmcrxC9fARlMeITafvPxwpANFVv4sDi1OFnXXpRyOfDVOLzCBDQif9fn/BPm
DU/jbMkgdGdyFjpyfucpBqve8g64vqjR6kYla1XGDfrU893PoZf1iMdBLKBUIlkoLfqwSSXGcDOa
PIis7PAigwSJhukcnyHaTXcqJURuLTUv5MnhCb9AY9tFoU6hp6B28YdUUQ6PUX5BKL5Fp4jTyA+X
gRvk8+35ID8A/CZxuR++EuLScaH+QH1ThfVD5qHU9U/GhjJ8HH0CG6GBzCZEnTrfm5GH626vLKYx
Y8iFo7MVfSzaTolZK6DQcjg4yOL8KtcCRq+q8u/HekHISC96dkbOwCjb55MRr0+Rkl0WWLMAN9iN
rhAPScOmxoJGxvM6DqX5ZAi+hOEcv9HOrdYrARX99/NAw0WKWJDeOEtKTKbDxgOYoM+JAxJvjQef
8slVNdam82nwo6WAqizeUmdBnovGGb6rQWSP5z4D1VctBPpnWknbxadZFpjE0vTDwxtTW4H35p+6
eRh84BmDlDQWr/ThCiFTyzO4rGdkTSEBABUg0Ic1FZZEjxsq/w6uK31wbV0l40N+a1yah2nODEMJ
QH5zuLRJLG8y57hv7TIrwPv95Mz0TTsed2+TkAqu1OqWnl6fV1W3K1ndBGGsqPLagbhumjGWdqET
xI+v3Jdw0x0bO0FTo1j49aQSm6lJJDewAgJM/11+xMb6EbPWis45Cg+2xbpBEPAtARk+lHJccR/A
mlCqbwrEmE+shIg6djFP/ZikAU0wvu+kdrH/cpBd+7ACZOidegnWD9PwPTEvOfvyW8tnvAZW5gmt
cClrMLpIcjYpjg0bOh5ugjQd1FGxS1Mnvz9Fb80x/BB6LKW4gue9Ae/DX4mTM4MkmK754EMQWlve
m2LOiyvscd79WboW2JEhdxKMOmn5o5CqIGatx5SzZgsaggz95/vnuNzRqGT7jSRKumncQD+ForBm
6VztaxF3BtzAY3qxMrtgl2PVdf2UuiIs3mh5iMJ8bUy9977O1zlcKLdRjJX5MAcGFyyIccbtJGhN
LNIRG1z1S1YiQZV0flHaVg4bBHZbFqfJzZ5ZhO4ihN5cw5A7KGpB2muFlD3P9DAx4PNZDvxhNsO0
jWw9QtuzeriLDZXdbISQPSHJNzVSf1gXLbuYRW9YEc0fnPpxC7nx7XHwRG/4MGYYsL5w+UNG1pm1
1qJGeFj9KmtdP0gQerEV0SgZ09mr2/ruAGTijFaEzGg2/VDw46OtmvMSpxYrvwUAOlQgEoVKuA13
jd57YpjN9alGH6gVT5Zyda2Wtyj41PsDqIH6Cd1fxBzsKvaBYuZ07/ZJzPZ8ibr1VJ4gxcUaaWCx
XQWuWJAhYACCZCQJdwe35X1zyIfwvIF7Jcj50gVsATMT6O1dwIxLeTnnVEn9BIoVmyOMzl1uxO+H
RK6BW9KKdsInHvy8xQcn4GB4ETpKeA83IKfQp0wwS3lHGd9z8N6/uYCPrXaEgOxwjGkcUBbfSW71
NSP7fs4f1CoHn9m619pO4sGIAE9W2c7icLjBdhMoQdQI/ad0BM9s4ZUA3VKIlUbi3Z/wlcFBid1X
sxw9wbv0HXiB/mu5tWxCZMgtX02dHylQXibEf1/tBXxiunbcReZm9tb+MaUCkPx0oQ750hz87b3t
v9Re11hRK9dmginGkWlW4NIqYvQC/fVCbO0qVyEanlljuKteaC6xYCb5RSPoB/E1wHYxHR9+2I8P
Et05IBr6vyYprQ39b/o8heih1Mp6ZW2rrg6C/D5SneUeeGZXSjoI0CxSWKPauPVG6I3kL7vYd4gJ
bRE/icqC+kyS1+InIGTejNx0kArSdSluAQsS2QBB95XXy/4zT+fEyRLcMnfb43JtaMOywcESWlGD
Ztx8jGyA1xQgSFoiLK7EPuwYJZG766FTI09DGTRZrXSrk80MLsaTT9OiHkuEAi+TxR5hi7ItgAfZ
5+emrad3WFhvYzRgAEoig/f1nAUEsa0bri7I+Mfw8xg6qso23xeTtf2M4J3EVUmP9Mc4O+A6jtif
fYVjRJ+fyEq6bZVViu0T471dglbMv92EMawQ9bB4d9xEJWbWm15lMg6g9w35dtB89jkqIDq58F2A
qqwgcI5Z7oHIXarL3ucb8Vh/hGsN/PO5XEXMwswSD1410LvO0KRnZ8/dRfjb11T+5vJi+c59iTrl
vPtWiQxU0l97pccLsp2Hpvrjsy+9E5Ju0GIGWzD61st3xzRv9TKArAAXMTEP/UpgKaV7eyDyajiu
E1UDXH7baO6IJ66MoTBxhZGIq3ZKCVDm7ObpsmVFz6oLsa/ICh5JgjDbejbuD7PBS3pquWMEn3+d
6pXqW6ATtAFyKh7PqS4Y25xF1pa4oi7cJKmQg2LXnkK9Xfxu7cNnxBK5HVzIFw1vuB7GOZ5wP3zj
Eh9xwgc9/OkPPRGde++IenJSttYzqwEIBma072LLhScc4RSzohRRPzkmJ+VgvqG7vAvgX5magQV7
NEkloiMi6VEQeO6FsFJC3DEvvINZUNvMpDGYRhYXcYojfRMU7W+CZKxdku2Fz0ee/L6EoBGct4OY
2TB6vDpChCoQsLXiR0za4mgeoLtuBC36Q6y5dn5r9Jtr5uJRcynejv67szqFdUiG+zNSEjazcF4/
EIggvLXmSxSTpyouJ0eG/7vACPFE625NqtzuydayORv5Vxfla1ljfDhOHepfCdE+z9kQ6VGttahf
sGBPLUnE3HTSJCNVPvTvxn9doLCsAf0eBbYYkMBB9yTpr3D/OtYemR7bUBAFrPQrU+WuSvikfQLJ
OBFSd+JMTZE0d4u1sNxbZvq3lokI7+teQ7t8bMXTMcm2q3lRRxH27GifmmBTJi/JigJQtSK2y7T6
p+LAGEE6G92e88o2CWg1dzCLVL9WXou73uTi481R4UcRFQotMdrwUr31FJxL+GgdXg6DoScPkiGU
g7r6jf3LOd9VuwV9Ghuvm7zpI+nU8s1xWffrEFT9S2+k7BIe0QDKY1KAKq8iuGtI9riiOgq/u5FV
cnYByJ2GBCAS6oDg+ylnW16D02PpTHXZQm7nHz+akuMOFRBRo+hh2FIlXAR4PB7/PcOGc4OFuO3N
IweffmIFR4nOe2uSIuMmuaJ1by3l84c8PNPHeex0sVgEUO9W8GHl3mGhfn5bH/IWDBGYM7akRFxr
j163WpIUh7cGsP88bAByuAB1jkDjDonwEy6vCAZcfN6BiKnlWofRkWLYVtkkKiFyxt7jGFGkTYaJ
O4xwevXitjCtfm6infFER68C8I3Tu4nE4l7mz2rxs6rUQbVI3VhZC5HkqzQSfFzp8mf6ybLMK7t+
QI2fHBTcnCH55SCJrQLYXWk2YW6U3+ayeKGhnTZ/Gq5MKfhC/LYbzalZc3fKn9fyccH6Ot9wbEvp
WKaKuEXOO7S6ES83+iXGG5wp5iXCh6fVxneXqWhTzbK5aYyTWTSYv7qVsOZGueFO89M5pE/LOL9g
7kqPOriqN5Fy1u3cWBE+ASbHhBYCR2jq3+FomO+RTgEJCdhJPOSyueWU4KwEBeQNz72fobQ0l3Rv
nMjxkRmizu4+6E/kWUys2ZPeUruwFQOewoGXJzrztu4VRV4N1tf+0eFpy0d/IjF+mDRhyZjUos3W
bnyrzlTm6wF9565lnseyk6PMkHXV+SDbyQZMihjOX4xOG/9RtNaxde44cLkesLqnzMB3dLvjY3dx
fl/8SEPfNaV45W6NoarkyyW1qeD7CHdxGevKX9Av5z7Sxv7U2/lUUt/QqWAQA5oDehQl2qPJ9F7w
x1pKQ8HxY+0dUvHe4rxZGfSS3U1I6fFM57FWr8B8GNJSsEmOA1cZvr/WESIr8Y3eTw4b0801BVqk
EiUU/Cgqr+Dh4aZ7UirvY9tWLzH3n5WB/OnZ5/X7NuVcD0VBnQ83IMWQ9Dk8y06DZQx9fH3CyIiT
jZHpTCJjUGOyWfGJqSPDCXtSL4AnqxvkJheofWcMZFAV2x3SSxHFtx150KJFkvJ0cuuvYufu7Rih
RULphq4kccC3BBkN3wZoLuoGANv1M0NWUSvk+IAqDBb0dkcTRMegYmGO0jVfacCUHTAEhUOfgU6f
/It4RQRND+ZqFmoZIA1ei4TmN7FEXvn9m5Maj51rSS5OLwX0x+jBf4WzSbsYY715maOkqlYJEp51
6ZcqZOcnl6OkTJMl7A8NrCnYtYDwGNooJHx8i+cMe3XBRdYahgjoOQTaPMSLYdGvDpxypJSLXVKG
a9N3B/c+67tCTQvTviLYE2YwbPh0qIwop85eoQzRHYWwCcixQzo7kXQK1VlM5vYIjK7tbKLIevV/
s5atxqI/BG/0JyLr9uOHgHZ7DvRMhLAX4hSdbZfMqP3fYw+VR+iLJS5Yu77e6FVNv2BnTMOnfzGC
i45LG3XRPUpIzZMwu5ltcOU1xB+4Lex/Ch55uJJBSQSMnQMwLCXuvh5aLsGm4kdYeCQLAMM2Da0u
alrrds6BhDbESZ2KQSs3od/1V9vNZZNjbZSCKiyph0zVyZb1SsVdVrFTY+S1UkHDsar4qhBJ2T9L
trdRAZMnl9mn46QYGF0qAZNQvOCzQ+nOjgfQCTbKIjva+deDb7bv5/FoE0Ph+FpUqfDOrwrKJCEz
YZ95463JLrN3Ozz7+sMydiUZA1g+kb9m8UZXUQpw307t9EkloIFxJSc9eFGAGMMvQmfwjIVpchHi
+r1ioZ29KJnqltAlT1L33lH5OtgplV0VIYGFTXNTmH9I0DOV735Fu4oEBkXAHgVfXy7TkquXhPdU
VJj0VEq8okDvn3EbEjXKaoE0FlPDZX7eQsnCaGIIt/kkfsbrce9MSx0VJxr3BCzPZiCVfUnEL5T8
HIcjfa2N2Dbdnsbh9KEWINf6P5DFdItADQjuH3I/4pySeb9AjTxTbYx/1HaLBUowI/eDE1W/VKCF
6pxl2xCcHf7GQnCAszd/13C1TUBw4NFF76aeDlxhU2cEFAZMlw8WRrCp4gNuujrui/gfO4DbkMkM
LMGK3BrcGOCwj2o8mdL5lV4mLPLN06BAyHp7UlAtbcakJlmu8Iffh1rQfVARWi4ujHJS6syAPzn0
7F5lZ661myuM+/ONB+1cqg7vRUBepVDwMRblBoUqna1WxnTojlmstcWObSBefl/d9y42oz6DWr1q
fJ4WD3uY+Up89yxSdj9DvA/wnsSaM05HLgCBaAHO1+2cb+NpGPzpc6Z5TonfbqGG8YL8kzus64Kd
oKVr2xIhQD19jTxmYTEW8oeQhE1cf0xzIFcRaZZApiiVrvi5ByJZFFvipf8fxLx/+wz3KFsJALSP
y2CVnFfQZtsgbiuK0VCjjWJ1zWv1Eq+XQjZZiRKApL5uyman5lthKU9KnmXWlpiuYFCtk0mngW5q
TylAAz1H70OjEHDRJPpxLOwZjKYVEQfEinUU2M2Bb4MTutjso/99mCGm/Idk7Qz0YLdIGVEbX5dI
TzHgzr7MlzJtXlS7eD/+FxtO49lGj7IPb7anR0SelFXkgS4LH09vICAO8RlPVYQ8ViJZFplCwktr
pKuLDFCVjXHfVzq6gnDEBX3uaMbgHlUwKLaz56APsxBJzU0S4KfDRHf1H00zBuReKAdfBO7OBysT
/eIo19Rb/9RmOm4vaZHZ6SStwvPc3V8RgVRlzPRa+X5vGb2kkU23z7E+wmM/bZiLyKSecvT3ovIk
ZQGNCnLvt+4RnRzEoPQ+9EYPGa6hqzdD6eUA0gRN1EyrFpmx6NoEgWdq/hchygP1auWIoYik0AMQ
eN9c/wL6xjhPOpqIiIMZsAEzZ6kFdeC93ItoGgLejpYtTEUpKss9Z41qvbar1g3hOux/YSbw3xo4
yR7JfoFAA5h9/68Ecnso/8wp4rWEI16Byk5ni1RfsM2/QtHAM7UTtIt8xi9JoysoPyh+LsLVx3zu
sIKFzZpatJOY9Wwaww7b4QU9qVDGPMd+0QC7tXeL4GF7YXnETDSNzeA8AuXWRAk8zU6heWmQfzi4
dIogwzCzZhIEcqLqa2AmO9qiRFXEDEm9BfcMYzvQ9vvHAtmnQ+6JbsDnQTl2aawQT8P7AN5mJl3Y
t7puDktZzNlU/mOU1R6SZBe+XBHKqeeSL6q1s+4FeaIj5lwLL2lpTgzh5LRvCsKbugqmFs0EDO8D
u5gyqBpTL1MNziTL2Gxh7MrkLQQkO4cYchBytO55ZnuQl+POuwQ4SErvRo6R2TVqJQMYwSILBMH2
/rgco7RZWGuGX6tXai7jQM9DSUsaEelCTjJrNTnr8xuVO9wAPheKh1TNxr28zakZloXD/aEOXq1u
tP3H4OhR+pxR/hAV0JYx8KkqnLyvY3RXTvWPFzlo8pJg7BOvH0Sb1eM63YSbOlEZfoYngrqS6mLB
oTcU18L3WEpCMPD0Sc18Iyi9CFpGg/p0G8GZ+nUVZ0RTEtGsKMeJnaAIyz+nb61XZMMuvTmL6k8k
wdEdM5qAcb1m2mQy5xDjU7vgTWkQeILgO6l8mEBW1VynEaHgiV/xvGeMk1ZOv+Fc9EKMyL79jfg/
0BklJqSPumHWPv0bAqMkYIhnjIf6pqeZLpdRKof/nDIIvN1YE54pVsDko5gvUPWKBCpqlyCFy7wJ
5AvVsolq/fEVwCTFaevppZI2PhhTzFNASnEbbnV1/3eO5GR9o0Nwk8mWeAUwZe2VaH89PALNrF1y
5XvAubjVWORLuB3pr79kubvDsud56n3xIiGV6jrE+8YKpfsu1zVKHbB+ja8DT3y+o1cYIOYvEB4N
/iztjTrhbb3NBhvduBezOeF88g6g6mbJDkE8fDZwGMjrlAWpKrO2NBjrO7LB9i3rIPKRpVOaQV4g
WThjSuu1FWKD8pq/qlBpNCMfYXfH8Da+osJUJ4xdEEM9aLcfIJOywOSlmdZrXPyd6kbb1x3rZsrE
CsG9NmWVSmER1DUCXs9e8Z9ISB/1l3lZdf9/S51NiNgv4etmQo8prJ7DtuQWshie7Pctsgsfd1q+
8sJTwg1JrAgPmkQMJlo0GihW7sSeUkOtkonlgOKKUquWDKQb6tkPWr59wE7OhtqSXLgmZeANaM0Z
FOBCl1gMplgnK0UWpWM02BcY85XqZ0+YQY7qL+KLzM62mx3tIegTL2WJNP7xHf2uH2N0k1Zl5jqK
Yi1/Mo4wJoPfvFeFXoyI5Ctq2MvL8SHsA5gvZzxy2iH7H1+Dc49UaPclOeU44Johf2k6dT0ky9AX
mOsdrdVB6ywQ4rFQnpFeYREXUd928Fp+OnGAV9BLHXIqZ6tUwxYV58TW/4YUos1v6kG0Ri4fWgn2
hLSjuvqJ+Wn58enBD3J7zFgUxxyfDaQzTJp01Uzlz9D/NMXN4zRJgdzB/SOZioxodTe47La2DJ1n
gzPDE6hPe6l3SfOtlWFL7UEnP1psIR2KWotI0n/9IB5fTBmZOZ/jIHWwUmdDWy2qefliRyCT+JSQ
j1MbHI5SR7kcrVZUKiMeMI0T049p3X2nNwiglt/sc6yHw3mza4iyzCSuOZD1xoxQy+zpR6XPsYGI
a5vk+JpChT/pRCTB/jSkAXDFjQO6xMA5iaO5KqUnX7SC20+rrVpUBlzsNTbeAeaY7DaoAOg+fkTd
j4wWgQouaiRO38a7OHMpRh9NchiNCuVYLF7hv4tI7hKxE1SJ8mBNTb90x6IW5DNuj4JUyEzWzzFM
yQlJUmO19ZcS/y7VdpAYR4nIawajO0AXLVC31PA+2E7S31pSu0aAtvjM5+/4bM51VmXuezkesaDE
m5VVBTUWkSSwecfP+Wui2gGPG/cYayPrbEMeDof4HFPbQYZO9mN5p6WbH0Vh9spm4730ObhHJ56u
bTv/wEaVYDNpWvbCFmWfPhjXB8C6L3PHBoX0W3u9jQTh+rdOGbdG7BGkcLybtxqFjUWh8Ru7Q4Oe
pXpS4mogef/GT4dQ6+38OzkWd+2FPklVzt53QupTm7xVjd+BuiAWe2cY/CriZoD2gE9jKA67h6I2
QCS9vQGx7ALFoFid6Dj9lkTRRFtwAvjlx8+o23iR5Tuk27coJkx47Vm3H4DoHMlL2fDraC5gOuEo
sosSo4cdD0iIl8xb7UmIWC2DHCAzfV3O0GygxvCWBQCLyqIWYTKbo/WyOsBUVk6HH32oqTdwS+cv
+5ubL5T4i9AGhSgEGBR/SMZepkO57mflG9bKoFPwyIkdAn2AsRYBhWIcb5WVunHN9Eubb8mwviMB
CyEmym+78Tzg9HIRIhO9Ao+4w87vAZk0LIR1gGVmX6ZtxiAXedBWuAB/kLPf/571/ATtBHsK/qS2
BBbIq4IE1Z3R7jUBPnzMBsaLOtsPAvOFA5PuvQXeSG28fCuS0If/hx9FvRgOwU/SRNxek3OzApFa
5kKO4xkQ01IkrRcIBqdazggMZBBPiC8XjJoGcXOLYDl1Tp1pKEy53RwyfK+ZLJdfD0jwQuYoKcz6
bLpW9+BAJVFQhmjDfXCAkN5aytRa8QhYJUUYS0ma1bXBzIpFJTqA5ewnwcfFNmgASwOcD2cEz5M0
2y/jXdp918D39D7FaI6XSP7t+7SdGHzjNBxXAHMdC5Y6u1dg+Mt9wkcncuj8d1ETR7KteMDUshxM
RT8xtgzFSz/YAfcjeaGM/fypfAMXJrD7BxBWUhvtEj5zZP+p9SfSwCu9XnTRVM+gOIh2+N9PJWdc
lupaK254lQdlZ3xeDHHjABts1ab1PALoFaDLsv+kyU+evVlNRGYDHKkubCA2r4qU7vXuGD5GivKY
f1AwvTrokC8MLzf20iyfgWruG7bwc3BjhMdEr/SJn+kQUHMbuKDYdY+bQfWjD8rt5UnUJwE9nQo8
KC+soC7eDfgDbZoeiyj0VxaUnNZAPR9PBX9IOy2W/7s99QTRXjsODwxk/dmrFi6q6fadlW6mTDBq
tMGkEloqTO+uRJphL1n4ThePYEHjzLZ1xjca0Ndf/58c/rYSEm8cn9BjeNniaPYWfeI/0MFw0UvE
XD9lHB3Fy26dxy4dxoMayui2S68Uey+cCrC6NRGaNWeG5+AH4VgjoSqJKNE+IsLe3WVq0ckqNSyB
9wamzeDZijhIR8x3R9zKsllmKsKDYqVTjPJgBT+3UfluXZBRycG+vI7+1y69MaiagZJS+T/xfF3/
spuj5ZCpxLp/2HrG9jJ5pKoaThKGcaZRN3oUj4Zs/e1VuWLK0onCKwkXF3vutZKcfARH7+7/VSW2
RJ5e5nwj57jW9w/fmjfat87EaupoMqpmJsBLaW5muWuwuyZYyMl1TonVFv7lRRID5GJv845EB4gz
dupS/UMcWOV1ETu2PFkNGx2fQgdMlJs/WdzALn7+0OI3Wfh4tYhw+Ng9ax8/5F0NZbAF/4pLH9G+
Fwh5Lk3LPxMYT+7tw115mnrpoHU/9afgaFo3U/UPE661q6lPHP+4HrKMTyOiuGrvGhjE/Q5RxlGH
PjNI/61WCMAgt7xQdq9mT+r90Zt+omncf5CLbHeJGBpXdGLxf4C5uD8rZWXle+8MFvMvrrjDc2qA
ah40XujR+EqmKWw0qJxMNwbopHBSCbDEde2Qn0l119enLHYzMNiZ1M412UtJECXOh7w+FRRygrRK
2JbwPHw2BaHUH3DljS6aE8+TXet0iXo/xB1FdFiGyq+Txr8UTknzUqq5ZOp6/GXec7Lkk38WmLAm
zhtBSBe2uyh7IpE4FtGIw6jzqJIPWzbx+oAXIvKOXHkAPr1+j2zNHXx/qoZgwMZZ3PzsxVM8s1c6
RbwaJSZ8n/69mnxMxpmdPArDhvVhwyruB+ZLhIw+sXFJEEnFjAUXrdWEnY9Zx9w+MY4SpVI6VaEx
0pM5SmOd7nEnemVoCkfTgjll23WzRnoBcEZLAh+nq29We7W1xZbJtDK4uHUiuWzgSBmlVnDgpzO4
tIgrRe/Dl5oYPErEmjZveuMDarcxviMGgUe0yzntpSlHO8RNbb/htstK+giNehsBvXRxyB5p4T7F
k8cnTh6DyvJtv+m7Q7txYHtw5GVpZgqQhFQ2+228AVIHMECLCKVhPuWOnfFWoMTz7DTneBnfZpVE
bz9p7gL4pn34uESnR3s0Jd4LBq0KZ7SpGLNMK1zrlaJrp53dZ9dRfu+mM6rBHP0/O06J2dz7mUDU
fYPSD9AVeror3AOYt+CtzlRdCVWH1tr3CaGuMQ8lC65CBP5BBzPfdXx3Hol6YwnfD4v0Eh8qlqSn
+deeD1u4dayehDHOBGQnwuKCUD1PTCxj4/gBX1R3h1OHvB8iNo11pOE3wf5B3xYUGEo4gXw/uh/o
eSXM2/a4Soyt6N0Noiiskb5cnyBcLzOmWG05AuzxeFoI/CuDwAbTAuqcbL7fS1175oG2lAmIuqmm
3u7ghtVFTnBLDHGWAYUE+54abpiSROu3iE16n4PSVmXrXJ3/cJ4khE4C0Y5bzb+evGDSSlodeXB0
tZolLzEDKUcvWZmbrOQH0GQyX/M+8/wSMZiUURL0baPy4Er7GYVMN9K6NA9lmH6x4IqIC1zyGwS7
FkMA9EgCPXpOi6WjpSd89oG2W1E9SSyDzYZX0U9LxH3TwvpcfeK2aAoqEQTBAdn2YfLPibr3qfFB
niTGJ8dK4jL2ND+ANibPs8hz7qgXjRCHCcPlfIk+13nkt4SmLU6mU3U+qPeNhwJ3aMNSHhNw6B9m
HzNVrpN8PB2bDNnvukIljDxGViEtKoDoFW3QdvHTJumxE9bkJ4fBargA0yjAWxo0l8ZqWDkhyW8w
hLBF4w+Y+UI1EQp1NwqjvaJs8G7eSw0gzIgDdLOJze7BRZF5Up5zk951qSPxFMS8SYcO4y9vtgSz
hapVVi84m7AcuX+H0E3KLahqT3IchlleYb/+2V/t2WHiTccW/M+bBCXcBWPy+i0k3IWQUsZJ6/wb
Lb24VSD4t4Kfrp466Qw225OOivJbYP+jaMIWugxCMC75Qlkgwv5OeYtpNH2WDHBsanCuLzPqeR/R
eT81jGilYxFCJNZh47gTrt1Q8heN7wGnT8X8bS5qKhN99/mx3owSwG29As/dn2eryBzrYExBkkeY
VwJeVSBo8Gr1Wlh4CX9pkqOCUN99BSgr7Nokd9tGB67Bvry8NmbALKHBaq+29QpGRlQ6Jv/tB2zr
XiZ3TS80IXIBAYW/wTSjsqvmdFJUmLE2x+vo1zHzMzeRNSbG/7wJbVy4aR1kd7pfq5kGCukWQdoK
9/mAo6uemGeWbiorjMpbytetRaYhruL/RE8jvnI1J/sgf1UXuNsbHROOzQ86wmWdjDOCajsEfIhj
cBD73GPjzEr8WlxbvyjsgkZ0hahOn9V49R3BxLe5bGzQyJZZ0j8LBYFCu4YO/GWn6Z6p8Fqs+4o/
2M4hbKkuaixsWsSFOUZx0uak8kv0VNBiCCHBAokozQ+I95ga0gklZRQH27vrBQ/mEo5CJBmtorsV
NsTI32ZHzOwNhXJwg3JdhSTz1ao7GG1DcFl+f1QQYLhMqpr6nZP1mU9XennOBhkt+5sVDG1xVdT8
5Ctb9LRAmoq2VdEXeGe1LRq2IsMt9oOS4pVwpFk/7/RBUZ6YTcGnm792+mwR5rlvHjKZKyD7tppT
VXorTXrS9LKLgt3zBzzyx08UL0iUWKjNB61RZDmXuZZO5vxzQ0gB91sh/hlv09qVrzgj1UQwyUj6
UFRG7XaEUyfosWuvIvxcQJ0T1MDoAGRSWjQUosMwrPVwx1teevy8VssdXJSnlrpcv5hVW13uU3+t
QilDycC3e1DJtCWvHLV27pWwkXaZpqVlviTMMneoVif/FyLNmPBp7S4k6Kv4E1Q7JpqY9hmTrwB7
Ca3+oU/rXq8dK95tvaFMdhaGQy+OaXIrhMRXgwmCbjqUwp6nDFPfiGU6ikRu/yD4dorDDCBVjdmi
iwyFj1Y+hxDBJlsS8cmhitUtMz1HYeHAZm5Xqfp3wascoRrs99fEJ10GkYO4ni0BuIAmOIhK3lCf
Z0Vnn3rwf/o8zB0CPsqP9W42KaV6veyI1Pts0QbCcBViwFFJICyw6rwNJ+lzyH8X5Ie13oykvOD7
G8q4PwRmYFQNIScx7btGqdtbMxHjpr6DjLEFQft3JNFq1uRIy6pj6ic/A1lUUXKdgyZMYWqWDWPj
lQVA8snI50pgizjgSLrh1U0Fh0ZpNrKDzntPhk7+YlOJCvRndbMiCXa1lRAaKqjVFcqH9JSu9FSr
t3AmGYDeddc2oUOpS/JUXN1Xj54IcTT5V1AwP+uic3lrt1sMpTVOnnMlX8SAn8rmHGqoBFeYu63a
LFAiSyTUrOjEkqYgj0k68YPiCTaoBE+3ypGJgCP2D9I7r85s/Qy7hue7pLZ402PALsma2f2UUkJk
R5WK6ZaXu04i8POSdbZbSxZDCgIjaUGKibGCqBybmElykbnsqxkFMQUP9WWzMDnXMKTRgZGCPBAn
/s1tQz5HEp0u7R49A70wfOpUNwFK8EUJZVelNSEzJ5JM0oLtf17cIQjkV6A+pLe77h2LzmxCdVXI
Ez7OGDSnKCjuzGD4DIpmcuEyA60RBIQs1jo18uLwxH1SzblFKh4LWRn+pRJr9nALsuHwZbE4EO1T
UV9ThagXNDh70ASoAtSXD7E7UvSrqhcDl84IVCZ2hGqpV1H09VJy0Dj/a/2/OjN53pHMDUqn48nj
mEhKuDaEJ/TY+Hki8C5uiV5F/FAUCj1n1p0fHs9Qhr4RFNXaJlzp3/hpBWmnPsM1rQ9v1jQ/ekyM
xXBEKzmKSlceNmdgp7r7rb4UVEzM9bInZ/ohlqj5DDkV1Yf9xvrAW5OKPmvB/zPYw21k6Z2ZI5Hs
xQP35abJRGaaXusKlWHReXgcSrwIzQ/ampXW4ihxQHaPc5T3g34JJ0YLkdpICvs1dwcBB/1pVh8P
PAf42Zz8BIAIHgeKf/El05i8G73He9QMf+DMlmVYwBgoi00AbzCJCDYk8B/WFR0+zmBy/LjFG5zY
QV5DMS5bFA5zEx7AE1ODzhijxD9wrGK7eC+5lLaZDAR8Hzntz00dIz/FR3PgBVEt07mfhFYnQGk5
px+YB/uyfQhb1p+Zpl3/pQCT69ahxOTafGGqahpEovbYYW5tCrLs2PgM02Ww1IXuRrGU+TX8ovcX
mo3E8ArnKc9LMetgSeknMWj6AJwUcgs/nZhM6lXuf0nWvIyhl2CPvSn6gZBxn0JXQupE4Mc0Vl9N
CHoIgeUz4HID+WuVczwVBdTWUdZLsiXentSTGXYenRZGvA9pPiPEgkd3/W0UwobOBoxizE8keZlC
kJh8d1rbDuzlWQb5l2bra+b+a0VaGB3PUyM0sxPQ2RqUt1uuiLIr/Ohoc5pxkYMtoR3moaHGKtOV
v4o1Y/nQq+2jap+1/CkLqaS/4J5EiYda4/DBS3Za3HHQEZSoEYkAXZueoaRltB5ONPdFIf/S3gGP
XnInSWzCU5rRlXFb7qWvWsG0pBiWnii6IN4TQiS2XGfH3rhRchRh68X53eBt6M9+grL8WQRD2Lzc
tCEevlJJqBFWjOs0hEZQenmcY84qNpPGPZbAc5JKZ71qNT1JOI76r7JJ2BPfvoUgOV1lQeJv7OqP
10zn+x83s9zAYiaUPwll6CaK2vpCTNMIO2mxLT1jn7wbQFu+ouryfPMI3Zscxjas4qCfLhn7JwDt
2LcAP1g21mlekaKL52iBaaUI+gxloH0aXn68OjhpkFI/3/HNJChTG7SCCl7aIq+5o3xyi8wFrdpv
/2LyszR/Pjc1U8AngDQGXK5XkBlSx64NwNcmAZrRDnHzsQrzmaKR3cqcQDkBGOyHf4YVFyV/wuv3
sDFfNjieqJL+AI43wYfVKodZVBJgS7WwwWwvcA4cMRW3Xu6xBTSJT1A3YhaBzqbhO6+UmRQy+0AB
RkYa+6J+tK2N9FL3InFqjlhJS3vPaOmPlTbLha89GE4W5+mqWGrm0ByLMn8L1HqvmzS/VV80P5W9
K37cf6SWMfMWYnhKqHuaDuQ+VNSRYz952nRx6SIlSt4Ar94LzBxM0jHYvWh2xuR2u1cb2iMFQXsO
JIyNIsdE9d1JjVScKXWk7X3FFHV1qhX4EN9K1SO/izS13phdn2p40gtZNefCJTZD+fk0RMRlS7wq
WXihOEsUUem6WF5xIC7hhmUZzNM8yZAhcnsp4BJzv2s/G/WXXs/FNB08XnMflJKT4wEMKgkymJNX
ilLIEg8U/34UBq+iyf29C00BoOEZJgEu3xgThEriuJLS6UptLSxd3uxJFrbbMRnF3QC+p+WTTFKZ
cm+kn11xJqW65Kvj6ex7KN20G3KGJPGBFtD/QOtZQDN/xdhPheYzyD1JrxXqJrq7pG2EC5HXWIee
khOlD/eK6xRE/fwmUW60XVoBz7jF9QYtXMFC5gJIJj9kmxGZZTCkks8xwXJB071qrA9YPz+AF+kR
zKJv8pUJm9s6mQqRd2dbvggs4x6yZznMb7sr9v0DPOLpDQMwmTRb8ft3MuYz/ogUsQjwTaejTR3E
jAhkz10SOxPDZI2QYevT3jJ/dPxV+BPPZ1C+yXGtU4UMAWQDirhdIJZUTjFkrwm7AP+UV6cOkouF
vQxZbOJ84f3/QdteW431lOHm83x/5/EbbXIrnyCb/bj0jIxPv7Kb+HtPjxkqj+BQogaKM5GPlKeA
gJkE0BVpHtjoCZtGeaHzx6w1rKtpIiI8COtfXxdu8/FitStKDLCM1/UX8BLx0sY1ghwI2tjgZvRv
fiCqiW/ndbSxLoBOMXtUz5S7eT0wVx4nspTjH+3dSL0ZaUCK/P9I1kV/KJS5zGhYUXlHGFEB6M9O
pp8E1LWLCH0lqGbpK8Dad9P+ELE1JSaf5uOwywFYrsLPKovzjCE7kfH/i2WmYhEhcVDSbpst+yV9
RCaLozv7eF9VkdzchqHMrd+XTK/hESw6wrqOQy5RPUYoM9dvvBVGsURZKT6aS1ZL8Swx1VCqDe5j
YodP3w8YXJSzQIb7ghety0Kr1uX/9Hc1T98cq5yFENKFWuPFcUonX3HOZ8C5t05s7gJvEB0QNh4l
UL6YgpcqEmV3JKdAxctSolsAGpcSbrtDZ510qHV0D/eBy76fdP5gQtpx9IsVEKJ9bO9q/ynqEhWO
W3+1lgVppm3L4WEj16n9bGe1j6A6ot5jCcVNjvZtWG7bNuIrO9uwbv0INckizo8t59aMH0OStjLy
V3joHvehzpS8SF+J2DKPpJ13TwwBchKZVmx1RmeBCPaQpb60j2/5BOgW0ixG9fYJ6UiHd9u8LPAV
OVgkDhY6LEE+0QPp7IaCRYl4AW9gfirnHwxo7HyQHIbPXJV1w/IEx5yK8j8gdvhIpt54ScbQsR1J
K0Qubta0aUOzNB+P4n9QW4z77C8kYqBqHg4ZkXfwD7VambCxecUlCaZgsXIM+MT3Qirnef2lJrjs
ujyZhz+fqMtF2du0pMGXyws38drNpDp57U7GByrxTux4RPfUht50bJ1C6nlUWTbhARBF5W9z7Bix
ehQfLu6HExXJQq4WtSyHhZ2weTX14nrK60QjLYOH0AhKRFIOn+G0WlTRWWs6y+YT/1zb3aA9jeFq
UafLXqc7vzIDc3dTVKqQi2wOT6oqhEwAET3lABIJKPaiWOYaB1Fnd52rxBWNrQOhBJvNOVd8APN+
N+BEVViixmNgUxIeXuvNMn3kDk82kcTNFzSntzIN/YOnPfmo0UXmEiY5ujWrIwAOSgisl7wES+NW
xhbV8hm6mx/sI/404MywfX9I0KoCu4JOOO/DM8KMgX03UhoHT9HiyYsrZlOw//Hdi2/5BCImEd2V
1vvPBbTR7Y2vQLHHrrZQBAzTxCVbsILUaf/ExhYxOcRZjUh41/BM2WK/nzOPBzpxXGm6rJTyU5e2
adCx0vHylcacbInA797DRfYlrYaSbXc+JVp30mZYsxFtuPg8tQUFUoPC/wlRGVBopFZuwF3OgYkU
u0q/YJPVWvnuF+nfmdVuhTAp8j9HTp/8f5OeTAq0gnqLIRBVy7R60h5NfITG+UiqyBzJK4gOiXNr
QDIy0d1OF2QiKi/uA3c8HdS8MqNj+4HBHAvy03MaCk0aeiZmDa3LlnOEkdRkPxjDc1A45OnQF/aM
1nFZxuzq9MLQn1yHuUaKd9wFX4D/myA/en1N4CdhMXdKC9X8eQwGDzEDab9jfmwOMKfZm8j4gic0
CpQwya+OJ9SdBDXAPDVDnjqIPFbHtSRKOjxKtBr6JwTQMvO2+Cn2jD9ZDAN0s/GC9igqbyX2pX0n
cOazTXa9Gkt8D/PJEGFjGo694+yCgFC8rdWRHTCi9+glyMXvofxGX8He12zUuuTT7pxe/pcdUvcS
Jq5TXpWHxQI1nVFQWj2PH1/sunmmkbJNijUtCAkphBiXDgh6QF7V0WhTEMM49HgliKhWsjeTgGrC
WaoW10rukoZ72JA1TlHkVS8es1+z9dm53M546ff16vvqIasLCNTmCiMdMcvWSSqPHgYByWYhiA3f
LZJY9sg3pr5lCQDd+aFQ0laxWhnN2s25M7K5vBTuyMtrN40Wo8w3I76g+okB0d7hlIf5ONf/2dQe
3e4jz/yE2rtqRSH9+R1T/vyMNDTjpcq75K2Fc9DU0OwnGYpDuOxMeTHwCONompPWAnst+02lAQQF
Jnj0x4coQyVQr5SE7Fu6xUDLsWC88ic1EaxcuTcnUEdPWqm0SI9uP5fPjqlK49PzfwimWkjGVnex
iNtXeZBtD0yi3pR01rIU3M49Ger+XW51nf0Mp4kQs+M+ncJB3yEGr+gp1z4+XWVbrCoOJsvzig3E
bmC2tebKTdkht60CJUMXYsuQuwS0kmwuvFHczxRi+jMX3GK/YP/5rUmNnjw+gC7LySAUYgmBZPZf
zuDTiNDTSlisWKYeXVlvdqM9inJlyejp1VmbbeAmjpA1Rpaf8wc6dRyR41O4oCWTRFAqTbzV98hF
rkomCg4xGORiKRqgMPE6veEh9an0CWwch7DUHd51A4vb2Zf4FhZ1ufgXtSDOPCAN/VSWSg5Q/HVA
lQJ98Kfs4SkO49NPPRBXBVG2FUW1zT8ziYqUOyuZuPVI6VA1V7U6KBqcsKI3T7zuS9u5oI72XrFf
yViL0GGCYI+d7wWA0ZR9w1PtyWegFog182dlipq3O4YcZ9KPmQKMW6EtbyRjauUuNHoEkSZJd64w
KgOlF7sLKk8QYj/G8kezZEFQXfXrJ+z24B9uRqv/apJuGHoFV/haBkbqmk4wDozEsh0pUuq9x4f9
xPUrfxhmO5sKJAg11Hyr1hTSRzGSgUvzDOGIdOBO9p6wkg1TJfWEM15hVoS6PGNJEhuNGcUpN0xU
b0kJIhMRUa5EoAASYPKykvXixVMy8gnMMjUe/IylfSQmS2lDLoK0co1iN/+rpI0PsTzQQDfnSDYJ
MV6URLKw5ISRvz9y6lCZ82cnd/7FHbqCr7IyV7VECuY/5r3i/6bzrMj9ivhVDi4PhbYNY48om5uQ
HquBYJLZgtFA1/z6DdvqCuITBn6oH9M2zL4WD4hkRezVI/MoVW3lyoFwDAeEinu+p80vM7+1iE3l
vi6cUsmMbzXK0YUFiXbPpLti453BkrCjBBtzrHVqw/xCRGUVhN7FiUimOC/mgglUZZwY8VassLRQ
rDibemfuWpvGg7FEZhmvkLZLdCWsMmtkdOcu4gol37FIIR1eP6pbdBd0/exWxd2hrLc7dCO8BBLt
izRxN3LnfsGrScpktw8fE50yTl4O2LhummwO8J4icRIuYN0e0N6FC4JUg5JlPyYGT5V+qJRLFViS
nSuPgGKhteQMqn+s595pZnnuuQEbVrkXaxGqgQmQyWypCF7vhAoxBgEPd+wXwfj9zRyPYc3fhZCc
OzyZvLVjrgYiWzk96pmEndiXs0I1IjCbThvb/HzMpxCdAMLcsgO2L26ajgA0EOBRZZlk+D5154sM
b9yWMdJiAu0OUiM5FGdaxVwB7W7tqIJvAFzGHr3GVXMniwmQNMFmolfdPbuNaFaZAjbHg+Qsggds
FmRaqJxEK1JLErrLMB1wJr6uu02QbWjgKLLqLhe1LNIJC8G7ZsJe0MyxtGTZWlGVSDb/vukS6kPg
tI9a4wlLS1sNSmOsNswete6KJoeKt4LhvMhL+O9NMAwWpbaXjWG3gWBtmrRnK+w9AncFz8zGJgnv
VbEueh6j/asyOa4/+QuCw53qy11kuD4s99nmORGiUY4aZYoKk+NdnZtE4LVl2i+uPXiW1e+COB2I
/xZBdzqAKbDhtCOup2MJ2lI7yMDe3WUaVyRd7BedSsrL8yxEKSNCX/1vSr3Gt00+l6JEoMg9H3aV
8WBXkGyllYxEpSjA/KezAw3N6wQdYsdLDPTFdT1UOOTgEm6/x7iQzPGRBzsUCNh0ezGQ1d6ncLbh
wBcah9ldVg50GtoXtVxHKyKOtwa4zdxqPdn6WEtI5/P1bxzJqXO3113bt3Ob51q4Fi1QN46eHKrF
7BzJmpcaYTbp9vezjKokY74EdSLvXsO/Qq8/knF2TV1MKAAJ53lr5L3GNeMdsEm5NWJm+72z3fHG
00A5ktaN7RNEEf/azbf4h+4xy9iUTvUcozBzXAdQ/r85ezDJPWVCPakmud8LXGtfzxDu1b3PvoE1
XGmaHI+m3M/Cx9U2ZFHW1HbXUu8JrLj8Tn4zO8Q4Yfg83/DeBggp/i15rQqmCzCcMXk8l7mRvBDl
sPXs2Hl5TpfBEEY9UtC//IwE7i6XoTkmEwyKMgU0WLuKmgoGlAEgleW+/3cgdWSgBWIPeRL+I5P4
OuZxxL1PvFiqIc5MUhPrCgMXTjY6HxIoC2ZMG1z+kPE4rWF1ZM/H626cZ0+1G4zhNzX/Ir76mgaS
AgRcGNh8VnxisrxiZAWvgqApwOPmhJWwJBufFWKxvWaZ5OGs9MgFvROcw9QZWuYHUohQopgL/3Ed
IXrVg8CDIEb/PZ+kP41lZNeX7L/7RGUaEdc1c8KJO7BLXDUtX8IjhI/w4MOHYQSgtHTRLR56H98Y
Idc8LCxmq3MOH2rI9EDmugTWEncRXKCArJSm0u1y2OtnuJJvfnIlAlfY+ftEiyni8qvvmnMAsTJu
G0KCZ7eZ7xlFr8wOgkO3blhF7XeKwp2FqWQ9VWisce2SQnDcjjm5jcPJk5AAIBkdRpAIk2tSj0nl
Rp2lzaeFJ9w/e1BBsQZ7EGvIH84292QZODpBFmgAgW9bl1Ue8lRE2W+Fry7o2DkbX570lxoyVZAI
6Vq6AV9tl5YrK/fuT92hex65Fi2FATKRFRulerTU9VsB9oK85eGId9InYT2qOfHLkHFaOSGzsl/6
1sSoPKHZMSoocGKZOcFRdj9UfLHUxRX75R+oJa/v8Y/2tW5kje/FhjgcpGFXzA/T3gDrhtf53NQA
Mnab/TceEG9wuliWR74F+cWexqWaHsUCnvz5v92FARfiqRBDfMGX1ywuc9aOE/h20AKknAQm03aN
XxTfl86Yl+BDf5XQyJa9iXoTOo4OTfZPHa37x3/RantXYgAb9i6zFPelxOfGbhmrIuCuN8dYeONT
P2BkW9n3tUKmLKqtDBOjA+yIz/STpM5ZebL0XvxD2GMVJ8pB/iAjJBZ4gAiREWifXoAcG5APrgY/
tLH/9cV6MZeq/oXHDeoSsgsgfgypt17hhS5VwmWdubj4JNd/e2EUUILvv9sYCpPI5Wh4zqs8WmnV
kjRi3PQaaCVxsv4sR7iYXoiLlDj46HbrjRlF203H71RxJVy2Tt/9Eh+VuEC1FwAgvQnZ+JugJ9Uw
LKRrucnAXmh7G0kXBHVoZCHnPB8qiWldrSyi0Uvs8Gkdnt5tTy0M0wGl7asbYjBloLGhA53co1xd
9BeY7vk/EzS3Qhp8EY2HewfeNyeNf1WRyM1ye66s4zIMQFHE59pkilLD3Nfd1r6y/kQAqtHXsXmX
Zl1q8wueA5kJKGW1riIy7gAozG3fkGhUywr57YKlOowWtGJ1bTxI9Er+BHKygfA3Hag9KaYA0EOi
ZBPdyB/GoZc7zhhWUfXULHBhmJlfruNcYxza9BuuEXwKF7mlIJft4hBsSyMwZOOFbKQfHIao1u1Y
4mFrjGantFSo55C969nWQLTnV4sL3VIRHlL8Rofi4+7Kbuo+XIsqPv1v0cjge6Ax33cwOzmohwGL
8zbX75ME+9NZQDQwjppTQwg3B70BfKJ/LLmzLFCQZgqm7VaKxg9iXj9T4TiPHnAJSnAEBUAKJ9w9
LpExcW6rwevF7vPHZYalS1pGJxqEQQ0eB3rVjc/AnVOLXIe3apNw8Hm08mF5nl46Y3e5pK6sP7OV
Smwqev6oS3yF+AbwR/GxT85klgXQbulxbFcC2jXRcXt42IC+SZvLp0jZ7QhmnVL/ymz5DrWcRIYx
YN6ZRP4c/hB0wN+rEIOl8S2jYB9D5aKHRNETto/Eflqzz51FhCNYIblfFKycksWEXnQfdE700wQR
2Taj2o7DyGdibU1M16dfd3DhnZ0mQXwf93tEt+myAUIf24erqgBG7pzCCnsJXpD+qplQo/9xtkIH
iTgcLZ04WsRDrnHychqJJu+OU0BDNKE8ppsD+EZx2ShRmMIg3pT7AHvSH+f2fDZV78fUqmeLbxy7
jYuJ6oxeSM6xdX/ueAMEddwAwkxD4T9uqGLyH8u7r4o4nsAFAZAZRdbsh9XIvLrkoOHFxla8aOUy
RQ24ETfgVamEe2r8n3t9+kfCLx7Kdvyb9bmTXWpErki7TcyVwbF6AtBpn+QwXyPvE+eyZDD8MlzU
xescXB4fqPBpicteo9+gFee9wU5Gwsr1Ek6H5r4DkcMV5Os3pXFe4312kAqU8sukdwoS4N8D8bd0
3DREdHH0UWNmK+P1DOW1eccO0EEPEct2ln2OEgFjR8zP1E9FvlRyEhYLbceQjjdhpMpStepA0gwq
s7qJEZs8Skp859S8XvBhukk6otXbywYfpBayOT/Tkp3y8MVEnm01zKMAF0itLq4UsYsJql3tLh+A
oIhoutBq0L0ZWqQ0f4sT8mdInRRvXiVs6rVXzygx6svq6IRdoDhy9pEFtmzm8aqeYhMSocSUJgSt
XevqHIbcYj7M7vlr+wEVFKUintBpzDG9VP50I9jMFGWF5VKInDY5z3dT1M6zSIuXomOolELrOGkM
oYB1Wvk7z6tXf6BoMcHV6cHAODPV1ukSZq5sbUZva9vX6nJtNh3ntXj3jIdy3MLNkncGs7p8cDN0
hyChfkpjP+qitEWgaRPK0UzwzALKbG8BhYWcqRbVK28hMSB3T10WcE1cfVV78BSwQiJ1IJQCa5Nr
bD6TiyzHVZIN023h4o0K0OgR+NC95rs1DdNQ9La0vIdkDRBL0I+2HO/Qm/tBW0/BhOQFNqTBhZQb
Cx60EhpnUPVVWFQ3VuYsUrf4x1FOSHkfpibtTam7CJmdid98LYAuRhUH0VLcx+HbR7pqEBKBpWxi
1bMnhCRxPm/4HqUSsCiJvWe2nbJ0I9T85vte7IIvzWEi+c3gIcvFkUQ5XnoGXjXJwV9vmfBPqbcN
z94uvboo6dwruH1bY60tdBp0oFacsiSCSeOT+jIXi4JBF3h2WLy9gt6NlXNPBGMF1EzRUCFSAyC6
OxvOYQaF0GsRVqA+sgc4Pkh2lHgWRfzrLwQ1zEHsX5I++9NZcjpJLjNsbD+B/4/JE4qBoEvVygGl
nOoozB5lZQNBq9FhOPrHzQWEinZ0yTbg/AkrM9PQOQnFD3T6nCjaY9QLxLKJv/0M+kCm5Z8zxoKy
yjW6WXYvGqlU4JmGpu257Uutxk8B/S31VES0FUyLZTGh398qeAtd4w0dFRcnELwaJWQ+15zdxShV
iKTFh3WfG1CJjSl1xz8KDAtGMUEiIYx4Ybuv+FsKGoEgIe3KWS4JGhRfWgFbjPHYzxhzEfjjAGK5
XUTu97gKLLrZr/8xmNApNIJ9uyH7nRLvz/kFoyamFptvH4zGWALJlR+KFIgHx4L6J2UEEKip+p0d
hw2duoU1gDbDjzFD4MbKk2bWV5w8T59YSCe9QGk6fZ7tPbDRvnPZYdoUYUDYVCLDaiH1HOXJN6Bh
BN9SaZB3BiUIZJ2I/r6h3fdvfZyOxqbZrmr0Wf+P8vkkZbaidF9XPIZIgLNMCQ6ujpNntftSK7NG
/SkitFZ0rsgz+Y7eLTVtuk4v9tzrv0nJTwd3ceXN4TI9ni7McX21u155O3Bri33cDoUZaHxTA9jL
kZGo62qGo7dGuA79C4kHTWxo5O1Yl2VmY3IgM8TqtpsUB/JGwVTjOE7qeyo4PvPWbpje+pI/57Lq
/++mp4nkTYfWAl6oeUfgsaLw9qjiS2dStCKIoJ06o0VWZ0jdbg3EXC3WibQPm9tlgUIr3bN0Me5o
nykPkRdyCfXeuEGcEiGTJKgjKYNgehM12PZCt/QGs2nVsntVe0DLC7Zf+iwLLMk1Q5jMS3xAZZao
87fCFu2/btGwpPGPKvhcsN4ue1CmDfaDe5UfguskeiO5HAIs6ItvIRUzNbmmW89U8noiDAGBeohC
/ej43GX+8RFTsvva9GPLV84CPTRrEvKRhfp4YnkPPrgVuqqK77aiO2osBfKwRqZUhMFA6M19GOfG
K5i8SFgwI0qDA+4qhK+Jh9p/Jx5rujxOiivseXwh81zsowHNqD/fvOdoRz5JTZzUWW14N6Pmf2Ph
hfuablcMH+RvW8nt/YXNOvRHHMMS+T7RMaW4dOsG6l9llzi1NGaCB9Zp/cEYqWgwwel0m5w/vhHN
Nd0ahu9RXfb7trP3YbIKafMCsOImZNp8L+ukTUDs9OArYVBPbWyvx5iJ2MYFA5nivFyExL88Zx4v
+HSuepqM/6RER56BBwqWLQZQT0qORTR58n23KmMHD7zEpisEycZjUsB3PDToSgX6RZsRPaiZKdYB
nenX+MCnnH5AOvyQk5t+KU6m7W24vYsw9khC+NyX7b/ey2A2Y7Bds9AqNKnc7wTqDtSIt8wyhacg
m17h/Rr3RlhaWKOdtGxjn/LHSXJRmmJsSM17O6n94LwZLxUTfOczvExPGFo9pf5tCLrM04li4+EG
gj87lmhnry4aqyJViPv+yKM0LuYqN8tSxfRrafzU8jfB4RTXO904G21VRTnzaMS0xKMIoHJgoiJj
vlNL5gNoxEd6oBiufYCo5GiodiDIV6sCJlLZ9lkll3d2ViWMI8B6vk0E0i1a/kAA7mOkECA6xR5o
HmmA8HNsUETVvWSShTDQ4flXbj/AEW9PE1ewtNE+x72mHcmT7hUOosEHNu61JJM13mx1bZluvux4
1n/kggLUCsGnw6wYgaO5hjGWIskU70KdzpJAQSU4JAb2qdgxF1fGQOn3dym2zIxQZjiPrth6/eW/
daUTxMmlKxmwokDGyQAXP4hkfyjIoS735x7IaEx0lgYPOwFcF8nIyywnxOeM9lu6kziqZHVEsecR
vc4RWwpVRYMLRHveGjs7MotsprnqUFz/ZlG2Jj/gDDvVTB91kq1re7oE19X8j0fj+30ps2Yn0oeI
/yEu2NB0Q4WbBa2w2i+0Sh+QR01XHa27HPZBvFRcs1vxr2I6ULBaVZwJaPac47SGXJI33AmwS1E0
LojYlS6yb9sgkJdOoRTpjl7ofr29t+i3AzjXXU6bB+hgYVJqD/Pd6FcWYnSBGDOm+G5CTPsAM+v8
9ASbLqjDoKmrv5xMudZm2kflKUzM5W0k/MOVIcyxJo1TyALkmOTCziE6jijghQ6BRBAPQqSG5WDk
Hzf86HM+CvdmWmnhOohfsTgx7eddQ80C41aQ8OPbzfGrokacqu2JjmS2xP/wzDG2w88nFXWQgjuE
2F3KOaYuQg2b147nBZ8OV9tUTVgDnSGvqOQ5Bf37g6DxkNwdSRpm5uTKy+h/AMf2fN48Jd1tpBKA
5PUZCoLYojqDQtQ0wPGUeHNAopi97INp8cHJEjDV10fgN01SaUr4CxeRVNywJ1jwg2mL971iM2tn
/G9g53WtqLOteVqH3YJOYD8Lfn17vd6VU/J9ezUFZO5OV2izzwbXGS62/FAzdi8kjIRqKeRFPlif
vbnkbbxukC5DoFy41Sjuuto3AD0cWhZAiLp2q4Xdwl/KbqdSCw+EFBJcCUyP5BdMijAkZ4iYXryg
6U1wZX0ivZI0dlZ7WA9VlVwftxd8kUbPGLk4NJbyyrmP3l03NCsHyM/y8jGQ+01akMf93beTzfkK
wWEtZB5VTIyDNlQP348cNRJ2Vk8crXWd43lQsAxFXtd1WzZOR/qIHpJSoy96KByOgWNquUNEb4A+
wUIeKiJqwhCLREeNAcmIZEQzJMX1J1d3RA3QlLg6OAcjwed+b6HOw5N5QSGcZ+S5MRSMPJmFqsDQ
uY/PwhASHe8u1mOG+LFjl5IQzSxDHynbT74Yz2ADsnyq6sGrYWH2pQYhWSGi0yhAe7koNqFQ5rn+
Gd8lZwcfY6w0ox4HTN8c8e+ggq5hImW6Tmt3P47L8rmuPbWq/FvbAfpER9NzGFDfUWNMfR8+uKTu
Rb8n/nMukHB/WZKOKhjilaCFoiqABWqyISW2zJ1i5BX+Fn6MhrTc6Vq9PpzrxSs/rbAt/jgljIIu
wDY5/tOcfKD4FKmtmNVZKnn0+ZzutYwnf7kaBjS9YNKzyE+45t4mjz5T6A4KXnkXMQ5Ev+pk6Pa/
s21eokqHRMMx9Qaohorp0xn/TO+DIKqSrrJSGOrfLk6oCqjureUMIoBQ0de5oqy683YFtggr4Zqj
U+fKUP5HToN0uII/WswjhTiuic5yiGUxJDNHjJa82+IxbwlgU5svGNKnUho8t0FnAx4/huqGsw2v
IG4ncwGbwGfZvGVat6a6z9u/Zl86FRF3xFtskIfNBHHU02X0Ek7covaveS0skHLIllWPMzyP5MKc
RGetn4Nt+zW2pKyUqb0Z0PK3YdQgAvywyjtZycDz2qSDvnGKP6js+pGFq2fUk+fK8ExuJ0ocv/V6
F8M0zmF6cRlvwZ4t2t+A9DzA/DP5ISV7WTehVvf6LXmFmP97e6MPyN0Fgb4qtnpvQu6z07RW0tAS
vFhwyaLCbmZoqwytmIXpS2Ag41kN+MSoP4N5yZEveadJFqJZzPZfzMdxL38KucCZ91C4rbo2mBsp
ANMgkECY4/rpjurOA//SdXq1cATbSRLbCZXmGhOAPXGSHP7t1dc6ALqD2UyNA19W26yfdtOcKbya
akd6JeQwXTlq0PyU18RCFZL3rD0OLUg5qxYIOgwQz8GCsmSwgU0xFxqnQ/wxZ1NglwFmIIehqRru
pbAjKWQWYgXLGOq6EIEdycDnYYG9rtJhD3u7OCTPE70oqc4NbLhFAKk0XW9es7xXI26TXX42PkTZ
XIJFRd3Svk/0sf7uOicNZjiJ+HDIdNnC5nHFpQ2Zi4bewyBsTUQg9YIQ7lnNpkkxtaimrjAh+/gr
sUGQoN5eKHYzJJjmmWW95USoMWdkbknTNo0PgIx4rZvkdyY1GEwLRopSt9JTMc6zXUmkGe7ZxTQe
OKWfhmeNGPbyQdCc986fvmDqyoHlEki4nutGch2JZjeroH69nPp2Lsyh914So+EHwYnC9T+0Dx5a
vVsZg83VqPLpiiyQYQaIfM8Y1Cyq/J/tuJwz/jg6QSxWuhNOMWlt8Hm6/hPgFZ2Rrjau9pMi6c85
bw9BkFC78Fa0t1EOmBZhhMuhV0jRe9kOUjnNJjs1gsyoh8026JigOtRVSZ2ePFlbsqR2xeAdT9l4
Hpg6EUMIqMfVGYBItcEKMLizvoXa6EyMipwMh4EFUV5y4i5fDJ2v41PIGGS25P5vOzHXbtCRjG0s
PYgO2FzuNWXsvnKPSJL50NQrdRKQmmYopkCWP/UFT5T+DDgADAJ/HuOmODmaYcvQsR+Mx+zQebwL
UIyT30OLHz9A6jz2+g2xoFZkW55KVjuJLByMNlEvlAWuPATbhluryXblJm5KnqXjGy9HwjvEBtBd
EqgUVMlK/6eLbWjtw3d7tC1xYA83xKsp5CKezgr3lmsa44N1InVLNIUBZpkcXPkpY3kwol++Ubpa
OSB6+IoVyCDgZ+nVe0stL4e/Hvg1MXPH8WeG8+k5otG8fkV1Sa33waWSZJR0pr/aKtGhykJFywc4
0AReBUN7yNomUw8yDRmVuSPxo/WlkSIBXeIH46EZ0Aio2OyppC/m+mayuv9piP28oNtXhvYW1NOe
ZfdI0gkAcZY+sND7bs6teneMlVndRUfaoKIohZ6AernPQSdpMV9rjAl6lIIAEMjaW+Scq7KnTxXf
b/loetVXoSCCaUdIsvQjXjW8ZiTtRpHaZ6iqwB0ivij8PB00sYSG3HY9l/53mmGALDCfQfisXJXu
KFEXCOvdbeFk5a1g651t3ARXLmuEjnWfmDMYAfj/KCvcCcMbiXFcu/X835nRkCEqEwlIL+5XNiKJ
mYL0CYdXNl424sZ+jWQuvIDQAZfEWlDSwVcvx2O45SimrBnNvjjC3nTl5jqKk6Bz8yItLTe17Nue
X9Lziit2CBxNDV7/MNKNLH/ft+1jFgvmhGgI0As883/vsdQRl+mNAinzRzfXzuO/tnPOQrFFlRXD
joXDq5LiQwG4NP7ALRFNFqmWdS/HcmZ4O3rTgp69VYEYMrDzIv4rSTvXm8+yInTff/aRCOfRwh05
VmhOaZXDiJIL9D0kab4C1xBVBhiwLmelM0vLJUEIswMuxH8X/wdVCvI8DzF2sYVZoax8RLQNTRdo
WU38vomXc8ZzsuvofQViZG4t8K+FensM7vXyzfVA8Hu/+0qLyBOKeQKQ4qaTI9XmujK/h+E/atWd
crOiFIQx3uA2VeBo4CARaHQT8Ujuok6UCOOYrDFvqVC4moDeVqoPPKSv+GBW9YZYyjGPxdwmxKSi
qvtjQqzQYsMYRGOh4PoZmtyV0BawSugq1cZMk38OQYviRT+A5kgBxXeihyb1RAATfpgKpwO59kDB
wHGDMGdvRz/wLXVQC+NyLjIHeVCdLP8W/iwMJjWbxGLPtQk12u87lOVRd7uFR4GhF/e0PYhOJfJW
kMWN6mrSchV0t3K+CJfhlyhmfLMTyRwkFn7V+4vJkVQDdCdZRzkiKr0SskZCA1WyeZ1OxU0wTumi
Ln6KJH9qAIQqf2r+CNj5GmCG1v8W6JXxIHc2oz8Fop5Aa4P+lkeu8ffKDqZ6+b90IGafzFdVGvpS
WnDqwDuNGGcZfcvnRhsA9w35KTW4ZYHCDYHb0NUbUGg/jSjJ6k3Ixu0Rdk3hCOj46qXAy5Lv+IxA
zII7/zexT3gFe/wUmuTRUJoKBWF6OG6WCxEXkqAzUuYaGzPogbJQ5qMZ0vtH2+qrM3Ocvb7h4fIp
kkU+AfpwCkDHCiRTgyfk8L9tPcGOwME3Rnb5X2UrX5vO+gG93wZHazGBhD8LPYcetZfYhvKGUeN4
E6iGUkivneG0n7jb1Li0HbTDdByKLmyVwQWCv351sHGD2Mv3Om6uuWMiMb+BpH67lkq2XpNC8vb3
MtsztVC8hqICNmg+l4I0ozNVfF148j3nVN9XMc+rO7eWjcM4vntRI6fXNi4Wj6nBxcHIJ7Wsqqpw
2av1xYFafEWtan7MOKEgw+UkVezb/y8/IsSKMYI3ODposaOVwmWSUraRhHnMn3kQ5pyD61h8z8/3
0dK6GdpP6CxmyoRe1JlWWPFzK3qxi8BDyA27pE5TjVNktqM2VxefQbfmnOP901Y1FoCJ3MW3Bmwl
Nh01fzeKH1ghJc7Vp5rOqQaaoAqvYoyMZ3vPdJPukmJc58MJnOi1mtoxVsYg5FBG3ee6VDWPDGsH
B1pcibfquPp4QtUu3hrJ2mQ3/VujvLfKzhmHz66pyT4ZS+RA1AgH3WGiWF97GnZjpVZlGZJRtr9r
pDEIEcQ1qPFb6VTbSW7+E7a4i8nVWWE/F9mPw9AXtqEITYPmZvZBIigoeMZpRHELyWFoUrASqOUz
uQBZTgUxHZk/ea01aR65j8KSrbS1maeEFE+y8vIiqaxPrtt1fgoA/ivLmm3mck0s8wfQRIyWQ16G
/EfRf8bq/TYX/xrjPOyUEFAlXx49OJhD4/URTUbpAGotwqaMhd5658QohZPElp3CXua+xv4Uq7NR
vN40Pyf/G99hOjsIsm9xMZJHQBqGtGpqiGlbqxUvMORCM+oCF2Wk12P2Pa5FsQIWq7tHLcLGrBAe
/WDD7KTiwczuH+5tk90qKd3uxyvlFdsgblxpxSOgYe6zCXdqvFGFRgF19E1NfVKbr2Ab2Opq7hL1
BQpNp7xi5HT6ZhUhuCyxsW6TwahYosJrTu5k1Ig9RKM/pKOIoNRPoHhwMiYKOWycMRzX/D3Tk6ek
z2fEtl/l7ZVgP5Uwq6xpTB3XqlL9+phRUd44Y6Lx/RE3iyjoak2An/ekWUN743bDL8SbnDr76ihH
qPrFgStvFZG04Y0tyrC5TLVerKqocQsNIxwumyd/0Kb5Je7eQoP74DZqD9V0m9eLsirETjv4TKsp
HQAhDoUPBV1RtdFC0NPyfq1Pr3WKQen5duDtcUQW9A82hxZmDoJxc+5mmHGQDesMmaVrWDPeUMOP
UlFWFY8Xmbu3fUZDpN+SY/7ytTk0AD2eGffHmZqCD4e/h/SUrdDd2uZSuDJIsNRTacdVBgpU9oA0
gjOlO7mIF79uJHCUiv15rIIEI0lgqpfe+0hIisfKz9CnZs1cfb74sg0ijTqjnlXL5kLzp1m8iZVI
OouVeKO0kmdjbF6L9xUZGyvh+sVsI3h3mFs+ge+KY5619gP/kieNwf9mYmC5fBg+tf20pSA6Ot3M
yT0YjEhyRWHs7GEReAeUtOkzJtZ8lGhBHzvftzjxUmokNGPwQOGIQMdhVIc4x7B8SUU1M9OXRdjn
XxCyh/22vGsloGto2B5dFgKRHRc+x6e5Gj2pelkhza01f4wIX6D+Gun1gXUgsscH+XfKALUyRGQo
4w0kqYPaAqb/pw4MbzOHREUs4my0Cq9njtLN4nRHGf7SaRpu7uGyoCQl0+GjhncMNLDiEKQIQ/H6
nHF/8R4MTiTOdyppn2NEsP+1nJaJE+AV1Ic31PwAMEamXBGDH2hW6KZaqYpeRjxJUVC7TIKU+wYb
zoLcZ3buN9GL/C7GvTzPJ99dGgzu5j3DiE2R0YwpBl2ygvHTjomfqZO8xBIXGL6YzBuqgZOlQaal
KzqMqy+ok7O6ULILdSFACBbYeZJ84eUAxPLy5H9K9ei+fL9mRQY+klBim/X1LAfQM+Lo/+8Nhj4Y
wcQT0A2KbpLkJ4zY5uRZ/ObYBQpAM4FjUIOb9eFH525KqXW3/N+qpVBNKT+8GK2frym/HVbKpL+Y
3uogUeIIw+ArsNSuEdpXA5oxu3W9iHR/UpJn0BRV8HHaVaheMfa3BErTP6GQTDTlpd7ya6Kr1trH
Xfi7cO3RoMKk9sFc+NehrstoTSID7L4hAaluQkevsY3nfIX9eeQ+B4HMh/JbR6MgtXdlxNOK70vk
R64TTzHeLOInOu35Q7rRFfqwMhi1fo90yneFmQOZfgFJCBPr+kvuoert87x8GUpvlahjDcIZVlOG
w9xy3iUezRLPKZRdGMHZ8QWGfkesjrRsv2yDB+mMZjo/nRfSt3yl9gxsiPoesupiV2yZj1nzx6y6
hUiQ+POI2tb5QOkMltX1cGu6SE7+BxMOYm6mKJi2w8oa5f7dpxaLpz30IY58cvHuD7VyQ/BaQn8e
KDkBF8kVAtYVGpToDegeDRBs9CxPcatVrW4FJoMb9JXcyxXsVrOXsYWph1c1HdTqbNAQ72wybuea
Gp5rY8rMm0WSSrEHnMGL5qbMc4hye/4Zq1a7bJtGMtkxJtBsw3Dt2ceoumipBgPR2NyOmIXqxZO8
d6ASXeYqR2CON53WE8lCmZ17Wjk3NMmhX3Vo7byaRpsZj7lXrgGo0qZwi4k+PGmk3YnSL+sp0dUv
2fKwWBhX78GNyIQ8XZx6P5Ubu8vxZrgB6g0JEemEy5ecy/N6WfbdyhaaNkWWUIM5m72ERplmE60z
/dgOPYXKrtdtyOvJWV5jzjv0v6543ukZTqAVVHtrCSztJ60rWIYqfhws4Bl9kbK5hPIZvEvQE1Gf
DI4twzVq4gs0pVGkPX727pfXR7eYivMoQgx1Hk8sseq5xHvJ13Dy2kU6BK1Y6C7Pr7XRJcobLiBR
WYiFq7E1RSUDDvvPNxA/gdRib7oERWDBMYJkFm+vexpJkb1NzA0/iTK36WF0N/dEUsT5jFjVnFHj
YxqushdkIYZhryRbMtiggzaMt+HAItoDnwCJHYnMtZjb+/NRD8y1y8C3Jyh5D3pe6lHxaO0vUuGo
K5sKGSvF7HLuaiNQf0u9+V3t6iSu0pqT2ZX17SrIgpuBdcBfG2ORrlxTPutlRsBWk6T4gC40C26P
nXeS56PEksAF6zsa6jJq82qvlD5dmQUYbIOdOf+Vhl6UHrM8Ix95bekyGd3VvAkDwEn+208rUHla
62a9wuivhfEyhYmw4NWe8lAUn6Mqz/QiD6D3xIt8u1LwtkS3YreBoJHsVRckntDl3IRrV9JNi4qW
I0TYLu6J9Y5pfb6m3CJTruARMwndBzD5bL51nSgnAlwhe7g9PBzmmwD9Fqfou/MLbKIrAhkHl8YQ
Rx3H5N0QPiQa/WM77Y2yHlGoXXU3mZMayF1Pp66phiNATLFKgi+FutXBiXkDQ289+xbckua/N7EK
f860ham/3r8sQGkYfUnXWP2xeX3ytMWMPaHa8pYyn8pqGN032JQl7b+F8SXFYffGnq7cekdpLFkT
jZYSMoLr9FfAQg/Pu4QscugP9r1uzrpNlqhqw8Kjry5uVn+GPjFPe9PKwbrFxqm2LJ+xjAd+sPmj
hg8BvIJclUkls5kc0iJlGFeGBd8/pNWspfden96CNCjJDsVzyMbf/rSZXyb27e6YZqPDjzr5LueC
y8lIuf89ZhzLwQgMBFAH5jQ2tVM5VAGm8+Mq4M76DCIgpoOYCeW0oVDW5N+U1Kzrb6z9kpVKVIg/
ybj1kc7bgnmLp9N34NHkykNBizkQiZ4mrmJrrTqrnl9Wide9pgLQJf++061mu994VDeQKwURadmH
TQdzIMhFJY5DjD2FEOygaN5bzs2BIMxtTsuIksRY3C7KXklYxzzMkS46EhreukL/rY4t8JAdCRJi
h3lHHWrVXlWjTvgcRuhFTXsToVFRJoQxmBr95gUUAYPt7e5B0w6M8QupxYsOKVWSy4vAIj1KjIDC
VaDp7MxJa9UIJeM62eFdIc2Ksw4n1aKI8zHlpiBUxSe4E15J2X/QHGA/t5BaXx+cwoYw5yU7xAp2
8YLogXCYcGtOH/DzSd5vYhbNNBj0BF9xZ7UKprF4hW35fSqToRuTAT+JUymc5yxx4E+bl27EWJOn
4ANVB20EMAPM4j1ND/2x/Bf8t7QqB1GhMmyPh/mxQit1AaCW2Z35ARDxmZtEvcbAxE04V50OxaSp
FgSNfHOQyzS8ZyhKz0ZhTaCWSZhnEMCjSp0vIvJFXbxYrlxLXUSJQEbgMsmjL9mz5Y+C9LO0iMHe
74GHkRLGWYUFOMaSFtjRnwwHKLRBt2owrkhnaZvtMhUNDqsakAbPSM2ekzhxHfmxpV8aXiZ8XSO2
8FJQct8W5fQnXEIRJjVLPTl1I8lLxy7u5GJ7wZGgcLwTl318zFxYYe7RQJdDWXV+9GCaIlXYU7Lz
eNOzFuk2ZGRNpiq9F0JOOgxdHu78mFIey7UF8d82Ep5kqNND0SAhtpkDl4I57M6fwUc0yI2pkYu8
V8n5jn4JdfF+7RiUrkXp1j7khj8a9cENjV8VnHmPQ1yBGVx5a2ra6ZLsPHdJ/4GwYLrEheGx39iD
t8CRUOKjhHc4SwmtB3usjonFpa8w/iCI5kmeKc/A8ZwGx/F6k2HVp7gabgjhaJQ3Nn0fN14IjXas
GGvpJag8ePTnTE5bwPG2A7UB9jRmv12haExsGSPs6tQO5Mn59bFO29SG5ZQty7uHzPhW2DfzvuN7
sU5Q/lQ1niwpZMxg7OSHYoWfb3+vUHMnrkNaAV5GRDGTc1D5ybABiYSKZGXS1CFM8cny98G8/qKN
y3qdKSpZDqli2wO4EVEoBoh6AEJTsXuDhJcx+iOvTZ6ZKBxBfxAR8kfsD62rHTl5poZ4fBzRUOAB
D0+QZUIqz+zhXJOaGJRnGB5hsSUOjajGVHDiuaaegP1lg+B8gmuTDzTk7xjFatuQ5YCHz+J/ZaWx
fun+2QdN8ttBXRsQeJ44yhSfmNNGcB7ZXddNaLM9ZzNXkpjpDTWu0/S/fs8Eai5JGYGrXxfiBccC
P/AXnIYeFfSrlfhRfo+GCpbASXs+V1pj050vp3F+zLPCWenpfrnPE9icYDmmTAJqimksu2vvCs2C
ZETuet3rBno1+/h7ZeQLr7O6r3uALvrxCc1VZc34h3uKLEpd0Gn26obEHmZXxRlMpLytYwtQNnu3
UA05MRGya9KU6k8WVxBMYw826+J5+x0iBgPdrEKJMXmoAsmHd2xxDaqhnapzmqmz6ioz33hwLhrF
V+pKYKTFI4dcyOsR+jg2ZFKniD0VL5p56i5vlPCclSLFVjqsekrWIzForbjbDsRrfHvocsik24W6
ydCJgvteRL1tlLOfiPO8d/xVPSVTtYX2L0yk32A7Uf5n0b3H4TFhv72/jN8iAzfxN37lehzvdts4
IHhbgnXyGXkaEfxywdpG3uDpX2+c9QwV+ndymOkl3Wan33Z3QhhLKjqtskQho4A3SEsbRE7PSFjp
lXKk/pVw8Uqkf09brcjThzVMIoSDgAYwsf0QaDLXW1DTZqL+kZ1YdHjSl425MlzZQ/OmVFKRXz3w
jpICNInfwVIpR6cWOOdFzia0s7qcadUlF78jf8rR8n9jy869LyKquosGKouFgI4k0x00nVvbAINQ
hQAa8i7Tj9DwCmbiebKdva6ZI15ZrVPLl/Av4Fsj9dQDwH6ueNE+MthW1Sh2YFzxgUUv9bVMGdTA
QDOfzcTMIQ6vrjBS9lXvXgqime5Zt/d+9BfE2et2eun/7J2TBAaJSCKtm1OVJK8dO40+RBjrwEO+
sfLRcCHQ+fwmBxQpga532QbVmbKsoaQiHmAMh/I5kgPPU0s/NpkPSRmwGwwHbcw7pyRUb7Sd/dAg
2Ogb42E0KeyE6t47O6443Bm9bHMn+9vsrfNjgywMGBVn7b/1kPef5M91DHmeFfETgIBIr9OAyGAZ
hRu4hqsfPNcZFcMxbyhaMokCLDwgncsNpss2R5RlOzgcYFsaakSOljXsm1FWqZX+DLQ6vzWSjKPi
gSJtd+HTnFnJ0RM7Gf5uHjhFbtdloBErIQpQsi5P0ySujMNcyQn1QbKLPXG5uHOHihe1au8X5Eih
dp/UY2P13pr1pQr7bcNT45klyxD/AiaPDRXp4vbJkblY0K72jKV670FuXTTi/j9Jkaofe5AEGy0d
v88nEIkBcOtu/F2oHjAHVLRWPDBsToyuX6TOPKMOwQQMt8RRSUjC6TqOZNYRoR/H+75VA/npphz9
UkdV64TcK4qTHIgvmzkH1kWMFLJhPp9UuebJauvf++MP9712tQDeOIyHqwrUVjjiOGOJ71c4HiCN
fytmEtD2qJsep6FHW2GQ0fMG+ytAxYQkrO6c5TQmVAh8yTyu4VA7b/FSxZcw+sNSIb16zgJzUKbd
3PXvv7Odr0SKVvOYOUUGGZ3gz+zDbPeB8vp3DxRGQakDiwZUS0bQPS8oxw2PO8shkNpGFPLQ7X62
u6a0FI6MAMFOVXSkDY1ztG9bAYH+h/LAY39stzr2hOulCGgsy8MAmTTkQ5WwvxD7x7Wp72LbY5uX
TqfJe/JZNJ8e1k9fVaNvkSLgmSnM4+uXF9NkvBvWq5hbf4QUst4LjMbZC1EEot2FfxAuxYDTfpgS
L4pKTEzi5ZzqfotfTbeUDS2+K9U4/Mag9XqnmAtzrv9Yw4pfwK+DxlUgRJvhFYEnycLf76tthErB
PWFK+vm9rNZU0w38aJFeRVfZibFOM7QGMJD185vGN1vzCAkFghdMI4PCrBLiFdE0XcHOWUq9E5BX
Dk/qljX9TDvoimsHjvhrU7xLgntycm6x/pDHtb9NurIes+Yp+af8oFQrWFF3p+tiUUS9hWrA7YAQ
DNX2oVt0wS+tDClwsCoJ2hKEAKy9dR/fCL0H5PM5g2NH3WRLIVgMiPbKUR3jFGkL79XW8p2Lezn8
Q1e0jXsZxoltIAgPrQcW320YFdGaKJBM0e7zqORsLVqI8iShWRQDWXx0IrMJB0zrDXrU+fartw8U
YASzvPY0XOKP8sx9beqrveqd9zvPraIHwjh0cjf0TL+yxsXo56Zoz7FYDybDMqxFhevG4GEywjn1
sGxwO0HU1DeE5/RWPf96g2Desc7XSMwTIyimzcAypUlA+42cBtAg8bo5Uok08J1v6DM2MKQZH14D
/iITNL5vT3x0q5k0GKAN3OqQnXXOfsjo2ntprSb/JtmCaPSRZMP8UL8mPDwo4ctrECXbj17QRwYs
ILrT7BAr6q7FKGnq7cKSlxMJGR+Y4EaP/QZ+6EVcOaTF/PzJ/cvpp+QA60uI81ju1rN31O3v9/18
Mvy6tk8doENNjrJGJ3As7sPMtYYzoXVLXUly7/4rhwJ69Jd/g4H8ry10Q6Cu/frwiRCSoBc13+8G
XQo/uC+P0HkKhtEJQ+WDDjdEEN+1JYWwsksoFdkYpYDmdOSmiv8XxWyWMZM5gqsDxKFxHm2TmvFa
aQQSB3MM5qcLndWEsHtmvouWCa+HO7fok6AngZTA0S1E3JFavFmL+5KYqL3gt6BxiryQgd3IdLbo
MfQdTUzRhzerWrzfOsZ06UMBd3sAmnS6SMZZKNNvuo4UhZZbl8trllUwGlJXmvshu5+XIn0VqBDE
Ctu8fzg9IDnp7JegEBIYpV20GBepf0RbSQTEnxI9mQATXFGmcEgbSotXh4qKszFvlGxObt0SoRLc
LQxHf1igAt8BTsG0J2ZiQDnxgJ8Y4rk5TUjbwAoPb+9RPRLWYJvUUQXUL3tH5N75EGFHp9vBlbcq
XMEfZWbD1s+VVCZvE5EEjLDnSpjxxabAhN0BqhHPiKxks/aBVXeFWv0ZNwAHHCtWPl2UbyLH3wm+
epaCug3hXD0nsgv8paEvWm3jMYDXmU8SO8Hs24PvtY/NDfQ8GmVRHZVAvqchVuY2pLtixeiKGfV8
Q4pE55PLJHiQg3bHYFZy0AlIFh688NHMRjD4Zo17NtVga4TI+z33/p9iRblufmm33d+oadnbGRpN
F+yu/O3WcVSX+FW07KwwJoDWc5mq98iDBOvEtTHA2Ay9rOFYjosxtGbMSS7GA+q3jhpIFtRRhHxp
mkbQ374gFaOLqzD4Ps5Y6OuJchPjMaDfINrYiIWox3QwdP+6ND+SmlesB3gzcYrrZouriKDoYL/x
Pa4LIi1+IydVySJ3aAq7fdoNxuJJw+kuGyIJDEWYuwvnySySIuASaOWeCAOCv9HboZ5DXJNVkTag
eidd54/QfuyPuboeHNd19ZJjgYepVfUoSIiKAbS3ttqryBLQIT0SdQkuFJVERPBarsQcQ7cRQRDV
WuaifHnxtVvg4E/EOu2c5hTNmWWMAE/styQeo+ONz6ZpI9t0rZCFrdmkA1Qsnz2vRt7yzKtjcFD2
uQgekJazltHP3231qpOPGZAucX8paD1YEQR86944SREWjVkuCCSApnU9SZ2Ol/W4KFEnopUqrxSU
dKcjZkdd7e5RcCR2priItOAy8V+hjd/2kXQG7GHL8w0pdrrP11FDhh+KZxAw02sp+iwvvxWkZLDJ
0JMwzmGRcYRgfT2VvyXM9tXR1v6Udj5+taUlXyBErvb+Z5OpA/sg2fhwtbMGvT5NL/uTh5N3L2bC
EF4dUpeZf5VPjJQfWS7MePQrF98He8emXLaocQJU03G2cXdg3Y1E4wQM9FS3sbC7wYyaHABMlZKc
Kd1WGuWwaKxR4D64l3d6gyksXB8/zliedBSvum7LmZpyCLpY1he8cPI0x0SvS865eE2W3dHE4c84
w9amOEkuIB2LknpKUE3hYyrX0aGMPMnKDNB09+Xw/oHoSO/+o8aFf1yOiwzqxH5pFIM/g46bA+4S
SmqFzItvoO6yiIgtQH7Vzjh5MJOjnwa6AihDRoVQ+TE2SP285W7VRDtNNfcpx9XYXzYEyhbFmZrC
fzHqxIIqElEnA0+geWcIrH0r6qX1i+rlVNXXVVns1U5Kd0r6NsOZn0iEs/wo/2W3A3Yj7HTpucwm
RMEo9Qyc+NEOz7gI3Z5SkEWPyVk2vGLXYa+4WzqimYNGtWkutvWRElm2s3vmMn6qqhQEK4XPFTuf
La0mJVFwLMP9JT3OyPWBb+CJKskRsTWh+Y7l7cqOQI21DFQRxgDdV/zZcz7wTsLhmu0ByMrgonFL
0+pB99qc4DfeT2RDzPqyeQ0jMCZHriCT52NmvL4tBzSKtVf9v+l20ARJYuzYmUqwDftltb8h/ztg
G0s9blEf0PfiOI1KafudCe9fwOyUmnOosLDqWct9nQRds5Lk9w03VXWpP4Z21uyqENl11gj+YiT6
m/wr78cm+le+1SUWKUE7GyU4fGnAxiYdMl6zAFf4pwEYq+aWV3n1JYmc30j5FrYKlz38uKS3xD9L
DgPdYF2ZHvY1uaI8vbhBYBGZnjhQ4dNtQ+L4hCYsf4Z6K5TH34WRqbifEyBaM1g7ncrB7F8BReuw
KFL9EYAy4xNoGfrMbW0gTgY+8r2TMzZ7SL0upnOD/WQeCYFl7H/xn4juhuo+AlM1OFAMUuTpMiSk
Z1v53wG/KeodhabRlzUa2ywiS5hFlOs1Oa7DMfGuEtuRtGNfV3sEvQlWwQIiSfPlJVAoJ7/pYlYo
mhRw1kecAnJbd8xe+5j55PUCGJDPSurrd/DlCG3KB3ALGGGsBAXuOdblb7dATIFemVtYUbLl3fHr
Wmwvk66y9u1CaHbINnq/a3z1x15c3NTceMWfGy0/Gn4WGHFo39MpdRr+rUD+OvYtHIRKadTsVhsC
K2N8ATmRDmvxGPPwY6z4KUv/sc9TOQqRCmLkhblcB3wPpyeaq7xXI5WFkgJwHuXjFodE2PACEBnb
Fd7vXtLo85PjRjj7IzVFFMgbWi/soS2MvSEACBLisok8syUgl5KfQQOG1ePT8RmNvhDmMTCG+ySM
n+Q56uTccgxohJ/CqndsdkTCXh3x9QytZnRS6dwCpr4pU9uJRcC+PDF+MzvATmrx8DVe2dfiQb+t
8Q9pqqpMu0Amj/EoGiyggSJhdUtpMwPi5n2/4OxUmbXMsV7MTsQ7Shg2rvHNOpYF6g82FX/BhSKH
aQPgZa8JmmTnQNZl6nFsruPgeFPQyXlt7aHTRn/eGM7BN7amo/fyR8wiM+3w1k1nQ+z+yK56LQms
5BTpps72KZ/7hiAdcZyez/k1Pf2F7o4mDV4Yp1iwD+tdgdByppLBw4vKQbggnunCDHqaPI2ql8KK
r1IS+XDuQgrzSIIzdG+p9APsdP8Ifn2SKF9McIDGkxfK2LgGqsV7V1uP+5yc8XG9AlZJyRAfEdGC
IVqESC/kCa9+Hv46S12uEV2dR3oPUCfQMITzKMIRma4c2KlDdKrHEeENoavT8e1yKBOnNSXrnQFO
LW8GLotjmZuts+1NAVK/nFq7Vam/NkuSXZch90AFYFiw9w6/6TSZ+cNOwuXNzymVM2A/Y6FYugWI
qhlf3TbGJKiF7Pnb9u4avmGOj0KT3ClyP2Gyc8byRPhcWJKaFSO/0wfLOmRipqJ1akSfI4jW+fyV
TBlJz0PmxYm40FCKWchNkn08/nQ/n52assWxm+kvD6AeGX+UlZVHpIUeSihXVd99EQMQ6FcJ3RW/
l3A7FKpS01tu9lZ8wxmR6Ql3yUGU/m8M2tHt/KtFKp14+oEmUmN0MyPib5HLQU4aUcR0C10CD4xE
l9mRf/x1tGkbU5bNg974xI2Y5NL+N5W/h2hUfIIkmHUEJrGBXO+Y+diPn5YGbo9vNdFKdBhvGvzW
aX+C8YKeTCjM/6opF3r2db9jgrInUfb2I3UkaHgg38YYjHEy1/tV9ORWxkGHeuKglsvQGToBLYXq
ljGdFtG+RzesZ9tPcilYtPvR4VHqJ5VXxSRBMzmJRDajEjHkxozgHk2pJp5sl9x60sjDGFTNNLya
1ha7y+TOdPy2zc7YguaD2BM+sGXeDbsa99v7e79HfltNiOTr8UNMpGvpXqqwVbOwUxYLZsu3HcyE
rkQW/Njlfv7kLyazhCtDXBtITXXS7pCaFd+MuWeuG9svj1lBMHyW5MOCjYpDVyxwpNROrOAh5AG2
TNngwyqlX1/ujcp5eOMtYTHMwiF9ZbiLAfTbAMh9PXIYS/+Fgsoot0Oxhcz8/N6iyTXq+DIfmN8F
0123DWUgPnNOIDcqLdpE4KK87xRxHBwiJN2qsZZ8jnZbFpMY6NTJ7xfBTure7HkYCH1+NER5osoS
9pURsVEG4blbwm2U1q9LbK8+6Ro7F8cAVDKtNk5eYW7RK04bxJ8ZfORybGQ2In9j1ZITPw5pARsj
umij7KpTZVrvZhzPGrOKOoEcMWnOqZZXsnReEWDFk0y3/SiRhG+7xejVz5d13J9/n3lfdWgHPnSi
Qrre1KJ9rBwKWClzwhCBWCprZl5Xj1LuVyfZYj13pKVLHW5pGWIJP03kvk+wCteqTYNfbVfmZ6qh
9HhEreItwr2/FvOJBFyUFF/Un/xAx3dAXuFaDznETzgFnXXN8n4BehxE/twxW1FO4rylWu70f97l
60QZb/bOox77KX6/4E+2nBs3x1/apuFNOc86aW2hTY83ggoulZGhpBkJRgfG4L97gLng6W/VPEMH
kWEl4JMPha7zyGDpZ4PY8FTEc5CCzw3cAcggR5LBV+dFAOJtwyYJyf6H/WmBOw/s2/jlFNcH+3hN
HB6s1CNWCyKH5GnLg3iHjO4s1eDXjGZ+AZT9cqx1cR0r2A4HFZQc+1w2+UEMPAeadPJs4zTgmpUr
74ySW4O5Tnci29Oje0q4atCF8JJDP5gU1OT3YFCBUfiK6X89k9o9jC0yp6mXvgzyAkkLx661dXD7
EzxuJNtdARtxNOL9G1samnGkhkU3vP9m0VKDMGnCJW23RimL5P8HQdnq0Yaon6+6S6W/1BzEjbpQ
55THK0SnYO1Du7HLsqwzcBEZVMS9rSGqRsjvupBdzwYEZ+oRFZnoRcTl5AvwlFEBqAr179EaL61l
8PsxhyCtPc4af/LmUakng62wKHQb6jXEqcuBzvGH0h5NoFhhQ2dnmmp+WP0HW2pxHsJ+a2CL56hQ
gPpFkSMSsXkRBZBLy46kqG2gv3+OkZRLWNo0c/FQh/wimJZyu1JMNgUpQuA4uyXaGgS0g2A9u5rr
UPPp/eEbe79KT3mzWFSV/lPuVSIw09xiFK1mhLuKQ46X7Jvh1YEpxXbtc07no9qdkoJrDIFztv+7
Q4sFtZkh9ROphpfvGTP4wCJ3uijVR1OYsoEnGsg5KZecTmostSZl/Iucle6peoZInVT5TudS8vGw
QN3J7xS5K75gCsOjHY3INND3KpKlUd66wfw2XaHw4nMluHgLNXenm1QzDq1i5l3KImVOCPDVqgCS
LZxVMmXyahV+q+ycXah4nILEDoomrFS1zO5uJPW/n0AynbEkwK+UonNpcSzH1DrdvbwXDfiYz0PE
c2xkaGUiHBPPjz8dvd8Ieay4KhQ23UBPyMGYUBDTRG5oU/XOj5OI8U/8PQiJoPuZnTFIUYo/WTgY
KUA2NmQgocOGrTVKHeyoYT+hzmq1OQqXekowBTv4DXceyZbOQl3+V5+xEOS/T5xIb5trzsYXJFSk
AW9++sJxcm68OwINmoYCvDJPegdNP8H2YyGk+BkCI3Q7twcHzMfGxFWKzFkmFCXg1gDYO7CWgYUy
Z0MxSPTKahFzKjr6f17CdxVFVZDkIqG7jUIG8ShzQkZGyBFW3RDgNpTf8AgazV74Dm0qQx609oXx
TkuXX1mjndaUYYvp4FdwLaLuTWt2sQRrDd3FyStBUL5kmNhJAn82N6ssQ4xP9UWkzbeu/fM1LubA
70lCvxNJbFn1Be/vfelQ6n5v0+Gzhq8C2Zk/4M0rLfOxXWoPpfkEzJi7vmpLYZ5yfeItdYNcQ8fI
ioHirwk479GdUJ/sjYkkrvVpHtZwpTvPdh3HPnFfV+bO90afGqsuND7FZOTYZ7c+6iRja/7ELZt6
KjPc95pzCAXYIacTLdjW6LvXYHhOIFCDoFl8/tFuX2ggIyeTsKvP/3Juz6lyts+QAmVGPG4CUZb7
AIaVbzRRLdOLgsmZm3AzmTG4BuNDMjOGsicMr1uC7mIkC3+XFTCWSqPifmTRs+70uT5a2SvgPSrY
OGN0JXEWO+xw3UvwmeR3j6BkROj6Jt7IoLhpDGoUJxPcC2m5rKINlDq3aPbYfPlkc7XD1Y5zpxmP
o/oGGmm5X0B6L6lG5/of2rv8wTiRWiXlqSxDMvGD3+jr5O4MA9SugI8EZhhoK9gb4tmHQ5djEAQ9
ofhPb/neaqz88WOC8NXmrwieRGgNUM4HtCZ8LsFuPXCuEwa+uGnKEtTYeE7cwDRXrfDxVF0TbtlD
9Q2+oKpvM2Xt08Alq73Okbxf2gJ/BLd6DyfEjg9ZjA3GoiUwsJoknfHST2B6ZDbbTgl9nIGik114
S2wO28bTs1E26onigpN1ishvZU0DUOAy6IVRTnikzrxNplnlHSEGBkM5hU2XBAnhRCPthpPDGAHM
75SelWcHAp1JdT68uxFiVn/b4mJGRU9PNbSEAF4UX/kE/2FLYtdgHT32byOdu8ORbbnEG9VZhlnX
DbsGwlPcbUkwitwLLEOFnjE9+nJ/dBDC+EY+9Q7iaqVnYYP3Qb0N2fPK/c8wPDdZy1Ih3l6HLMCS
JauSBguZjH1MS5MhZPyigpFLy5XwttjH/gzhPfIfXtuRTBS+vhrkDKg9K9oqG+vGbEWXFrI4Bftp
wi5F4GBUWik069A0T9gSwdeuyJgBjpZ4lxhfsM6ineaxEFZH+YfQl7r4hxFOsgLTc4pnQ2uVt3lO
XeTF9kKEijokShc50Xu7KtMCatEznsOFdM6yYOJPLJsZgtY+C5X+3rJtcFW+laMXeZ3KI7qifah7
BKtp1scNSd2RTxpTWazcgePfNIWO9Yu4zazjw3emRIdMR3UcQR5/SYd3SrQAy5IoHbZfsezgtNtK
RB6zfqrWO9E6KqifrH5+/bFoNA3/SpPD4LXTKgS7sT5xe2gH8IHo58s/PFqhFfd/xJLEXUF9P4dT
U8EQQrBHw0l8XDWVb24xHgHhADrIvAkhmQ7PE5gyYQhJtc4uP14NTT6LAgaBlhIusuTOIsE8viI8
nGVDAdac6Mve2vd/bRno1komecWuFVYvnLCcFOpNmqt/G1HmihyRdF3Yd9UfqIQmta/Oh+ruXrvO
K/WNn97Ejcnu0Gn0oKt3DyYkMvUiQcIQiYzBgDxpfSfGBdlIqWtFP8BfNvFkyPPJEULfR0tHiHwR
cetfWwGAC4YzLVrGQaL+hwJ2weHmb6Iu8y+7B/7gitCO9UAsKEx2ElvxQe2+vOuRh4EMGpw0jni9
ptLDTAeA/FaF0mDtGfgjGEt0aOA8dFs5CnSO/PIqUtIX9wcRslfZJRDbCOVLfqC3okkGsmzHzKOC
Dw09pfZlMCRDJvxL8ycC8rmbPkYIvc2T8rmnmJ/TvGM0B+XCJ93vv7v9q08lvvZQHkU95rBel4ba
t3rY3L1GZ2iOpjzyHW/g6tJszt/dHJZzrlMWgYAU6V3LlQ49cAn05QwGpGZgrXDF95ZBa5Iw1IkP
wNvpFix79SaIMQ6bmYDDOMyvdSjW3whnt17mJPK0ZfGy+1Vxax8RBega4zaTxkKi5pYCZdU7+LhD
2lmUYD3ImXOpYRdERZzwjsm91sD/noCukSSRIjL7CtmvXWdjyKp/SUi2rlP343fy/vLlbLxLgHzO
RBc1a5IQUIos/dZtsRIBnBfS1X0iwek10FrYYV7F2xyavTG9nk8P+NHKHz5XHTSRyU5dMgh8IKLZ
P5bg4s39aQ6PYfrkRVEsOEtm8ZC/Pmjr9iNBTLwU4WCnus4xvvETG61W7Xe8CZzVzQ222SpElcpc
vLmNatniqisoRc0mN38Fnkr+ZAN0q/TZZDfcjjyzcGgKQHOSnmxddLeD+QnxafoYNMyN1Fk1X5RK
d07b6Y3DKbIqy/DPerhtY/rE65a6nbLpUHjACZH5RcHS1lAJfXXDpXocbRfrWJmSghjrYAAPwMae
/uKJ+vImn+pp32I5rGicC+5J/GsBnAwQkYp7t2FOOxDbB7xZiNzP7Gdq04dKchSQVssVopTlBxJd
nXVBsgb4kSliokHu7EW/yEzfuE7IKP4FdmfxuuWpI5EJt/+z7MHQ70CkkcvWFgVU1n6lB0v7snT0
dkXTEHJ6SQ3OYxtqwPxLrVu804ex2ILdjw9EOqWawMVptGRk60R2rn7RPLIVNYF6a1epMxjZN7tW
IU0Qk8goMlPBXEbxM2wYuZp14LVMneqIknx76wGxfukJOFsWjOClKgeB4wNinCpsQGmhKrcKA5cP
DErb+/U4WCC9InO47W7aVq2o6Mxu7LBXKYV4SV0r+D6M4ME1vqMDYKbO8cCHp8hazDUbnxCo8rjk
fkPIuPABcfxeFmRAbw7i+ASIeUcCbm6SfXIBOhjhfIOJEahPm6kuxKW6PvXGb6s+PHgfwcwgtUFj
4xetlm+CqCqbjgbWt5xGPHy2vJXrIo6QP9o9YsezmL3MsfbD11cWThpuPvBEJaXixV4pfld9pRsj
WraDBDKLcYACzibCszBMJmdC+bgVRC3xAygn0TGbMgV16yfvLqCg2HCMaGCs1Wr36M35MJYkALXn
MRHMJIzDTbH2p1Wvh6XLEQGfzj/A5OKptHU3YezH/VwmPdzUDYQVldAt0pTYGEn+CmeQyY3yfM1P
zQnj/LwdPNqyowVTBXr8H8fXfZYsPr4ixV05OHOFpfwftEbe8o3xn3yg9R0va90eNBajvn5LUiLX
+LcTppudRB0QTYRzQQaBFzKUXNJBLMbaJ7a+zB35WRpMkBv+y8Wgpd6IDGrZLkyAKEk7ner0Roqs
gHoxLHoxJTVf4z7IUiPZDCHgyCox5f3xJV/YXxzHxJuNHC8RKVybo0QdEYJc0I4mDnRiWCYWDtsM
cIzmGJUNougJUqV22lJ0IM0zMSibg9e3wNS1uGBgCU2ENuZoZ8l9Zi7vhklNiCQnuSqTliOfwUoN
LmYCjcnhfDquoeE8CQrW5Iop6ZwmsNflkK6m07QmnQ6YwRzT8FECVR8czs8lplsELzVuNtbNOOx9
jcnCUd9wLRZxFxtfAe7p2tGDuxYM1pMMPbWgMLqz1J9B2m7eYDC/9YPJnMk8kE8vxr/1o2KEv1H6
SnfSJ8e8PwPxKI+4RX1VXz7yIKwiqMvGr12l/qkBY67/ZpQiIyQDLG37wdXJ+G+HC+Q9qF6pjpKC
yH64xpVF3Y2UdUfrhx9pWSLs3sm8bFPQg6OitwXfrmYpCynMrEkBuTgQRpTqglVFr6lZA3VAXOmL
Vss+NWMeM/QiOnijEULrD4b1c61JMvjfJM2yfL8iUVgaXjYcafFd/zIyJDLgSKYltdXJCqGGADi8
5AvEl2iFFsqIgJ28edqfjibRrfMPhR7BmEFNUljCmncewGNltGsesuV92LgZVsFcUO58FMP1vAln
gTgU+CH8fHwDqXwXijx/3fX2RHWLtnvFEywkYlMstWBB8XrCRer3s15VdgbtuYoxCZj4j276ocyz
m9RYo1IwXrKv0F+tkvDaPOH+CNy95g0Kh8Oup+kHo0JTvOVP3qsNB+ab811XmIPt3wmptpCQW4IC
hTKomHCkEiIRkpNdkCSXX3AiPCQCguMj28gdGhn24EinhtDixETwaz5Q8+xLypMCuNaiQ2OlVfj2
dFdrTpzQ7iX6nkUEAN5Md309hvczFAkViO6kdC+pJ7Q7TxKZWUx6jfEihN2N4V0jR5mXP3qpDQmL
bTmendHf7kUqDN5Ydt3AEwN6uG7Ozbs1TsY6+daoJcz/AsmNAgeolflChK1yiA04CSB6fgphLvct
93jHNSFRE1HNGdqa9iznT9Sq/T5BH2TUdm+3WKlS+FdjfJ2KcsyNNFHZ8vAUQznUNLbhgn+XyrYI
tB18Z2dSOg59eZ5+pIa3QXgT6VHZjOFlgWRsN1wNIH7tYXI0+JwP7uZkK1edBoEzWoBoa5sH6GXO
V77knKSrjrxO0QH/O5+TouTfEhWPg5N/uzY+i9t5H/nlaIiYNC0wAuxo0ng8mxyyzqKRthRRHaMi
cuI+zo8HDVH5zCNkEnun1Bt4LQIcHzEj7AUNyJL+y7QlIu6Hl1CW6yi6jPxVcWWv5jPkI1r6tO9Q
VBKkTJ3Yo77L5kG4/sMjULDS9XDLbMCcky0UG9vYDB6T0/UytDsSUUSXyUCIX1pHiVdiJbNvOPY+
AmDtqH5k5V2BO+kTWM2DXhRJvwQ3G9nC3HxDrrkfcG/9iFVf1TQ73h6WY3PzMe5Cy2KBLtzYDC1/
0SWQeBExOnZ1Lz11vwbT/s3avm0Px+I6fT524KM0He5kUF7EP3kf1AHFXyhFZTp36mJ27zmHNtOY
FqkdVxvzPk46nXNmokwOCO3qgkhbo/cm861HFtLe8oKCvvhS9FR7ZVFo+ORRGe254tnHr2egaEZ+
7XbXkDk5b/S3bf2MUMGGf7cuQmWGO7XhnisJV+E474QlNH9q0x0urdv0z4aduEBCA/J/Imw2Eici
stKyAn+a820Uoij60eAIZidzywGvHp5toHb8otVlf1B5aSpEyKMYyqutLdgRjXR0nXI6TdHpd6mq
6suMfP11lXq8lnq7vAKjpu0w9hRVrZDGRvgrIYMHoLLArjD19XTg6CcXSJT5va/X85fixpqC4Iip
yk8AvcPfsH4Rm9SdorPg7v7DLrjg+SUjOugwAJ361xlae3o9khddvyUc+eNpPBmv4gmKnaV9fLyL
ZADX7xhLqHFqjg/zEBBwYqDIcbh6w+YbHjOMbfSvBRr29k4YpjuGunLp5btmtfRqQOUokmH2Mf3c
YcBF2Koi3dGjbx+LsLSFUcyQuwRLE6Mf42OYgPeX3P2lZDVNScjM8Ph7xifnsfdy0zGyu+79DzC+
uErWi+UL/Qe/7S709wSPQJxX9QbBYubGd/7XEwFyQR/7G1o85OSq9eL5tc5u1p6ik3ttZPkX4GLG
1bI6ES5ynmhBW0gCyVlcOqnmkOHM4YquDuZ9NK8MCNti7pXzvzuRFztFvRfvov7cI1Yu+3R85KQo
PjO3sA00oU/cWC0zS36DwyXcUch27RBqKYe/qlGw11++CieIj61VevitmNerBZiXhQo4fLbuRY2Y
slrI3LfXAq3qi/1d7IZem2rtzeEgysNBi3rt0h1xcdaSYV0OZFNq4yvBvHxxL6WuL+ucf7ADisfh
IOlYFE6O2t+gnWATsQScALRQwaCMqJ/4OcfMN4S5ZMKpkIIhz7tGjh76Gt3Q5G9+4lnmE6M/CsX1
198QS6guzbmB2zGo5HmOavwYEEsakJsZ2kLHfNQiOGXJhcdBSvC6N7I6JZhpngs0ro2KoeKGr2W1
GiNuAwEktW9nEdNrn5nrhV29GwQAiQ8e3cyHDcSaK4cV9n4ot31WpKlsdbS1Y3HUjetG2aVj7Vhp
NEqSsjwAaK0o03nbnwwk9fMbOWqbwSLh5yTEsSKc73AlYFoMQq8Q6Y3vg0RXFDKqg/RNxm9bmM8i
yHCqMNjimxZ1h3JtHI+33zylBe0/fk+0r3hJEesRFopQwZsCDDug3uwR8OBdz5VBJWCbRtGuZSOV
0o2sCu5n7X4kaCbTkq8S0oFj0RI2+OrxqRf2Hc9QhGOnmJR1IvWd1CJ54RcMw/RX66aMyno9Y0eF
4Oem3Q0pxYQAUu8Uae3rgm5MKNftwtCz3F+oUYJ+qq/KPTngRYC0BgR/AE+9L8FzO9Gdr9I7k+Sy
/NGEJpTTRTQDKAgG6tluKAbufSexcGEbnbVwdzEVCRE5O0kPkNa4DczKHlbojXQU2AH7ya6TYY0I
0+GZT3NB0Qw1Os80ZKLCXP9Ett/PRapks3sPZKSOof5ZmMASl9Pki7Z5WUXmpTbMENmevQe7IKZ/
dfLobs8hRTXXRj77yx16SZujDzjmz6Owauw4faAwJxVo0OiK95ro6cEf6muUvWmToHrIJfEDNNLt
ceffxuCtAIJWRVuXvIMYFjB0M1KBbu7BQyLh8XIgG1Q6L20yTbiz9c150LkVcG76Yi5VYG9GFZrv
rjFgqreYF6q7cDTP8SuC/SxqzLtWjlm0z98tPeTVWEAfdodMZGmTzxH+Fd3PmeqUPfBB4FHcON3E
eDfYw92ViUIhKhkVF1h8vwlY82JgBEIMNxHRf7yx2Ny5xNDvSVLEnopbXlMGgZHq2oR47KRcXQ/i
avPEjAf1PHiNon+MEIV0hkD4a0nG+xtlNmRFzZ0dyaSV4nDkEkx54hM+IXbMMFNtLPtBeU2O8gPS
V2k4ZhmrNIKvCe9PuAcd6Ifv1QQ/bSk44N1Fdnc7NF7efHXvl4+hHj3YdiGh9RXou0t3+DMx3fH1
YOyzbeW4ZJY8C6hkzuoRrLoHC+77KhrBvuwqJ5YUjyNUlAqEEXA0Ql5J6V1iFUsWFEBfe1QY6dcs
jeIATc9/fLd1envfMQv20KxNrP9s0ypH8uxbu5NOvkVbRqW9jDByl9wyjmlpbvIw53SPo2nantnh
Lt7fWWvIuLC5wDl2zTil9k5mKWowmfkC+aSlH3W6m8j+95OL2MxU1lLWVvjWLHVwJcvnHHjubxHf
IUf3u4GFBhmfDpEWm/Zrnc+Vna9WQgElOtqzwLIIi8znGa4HLgCp+O+1V8ecVRmkqHZ7kRfBOD2G
fEY/1lbeflbdrp+yeZ1mRZ7sOik4FmLm2K2BEkWamrjxyYckZhh7eN/5EiCWWSGq2ROhN67TYKbZ
1JkFHMefvfBYB/bJlygEMW5da32DLHPioy8cHqK4dSkfRyqIoRj769uPrU5R5PKgx9CeLMXotO8w
bdUar/neobc47pFdVUw7mxPE7dgqfeYstBl0Kjbu89NFByRRDS1/BdHPDFkRI55rKJKbYHokf9v5
6a5Sg452svlyzBQAx09fDSUfs1/pa/l43CytsChletAkxuEGR39eqOp1+8qW2C0klXKp6RmRGoiB
LcA4bmbSCyzr5e+VTaR2Fs7fK6StfOJZnFkPO3xuJtj3idT+IwH+KibGjj2krpGjqnIeF4fL/pgp
eOFjl+xgUVO3ygP2JVAhf/q/nwKeFxd+BIwUDiLt2pYQZTeDe/P5B2i4veQHI/6x+WINWRhH9m5A
9WEeOP6R+yZuElc1quaelpmdo8xp9RsaWHcxr2E0AoM2Cw2xGYewxcXFhnDw9dUy7AyusqjnD05m
NcWCIHVmnOafM/y+MZ6aRVTAg6/9wHLQWdZyJU5FcM/MORjUE8yMNDVfwS0N9Ed+Gze6eeUHpMWC
4R/aoxtCKtAA0Em6SucJBHrB0dHT8CvXRs5cMbPN0M6qP5cwcP3FYzbvLwG/rXKk7k25A/BPkKIH
GwUJo4IlJmzU4hlAoJlCnYfkl5nbhARUUFFoQBuEA6pP68X2LpBXnTmCqTQc+ZofutV/z/iFhib8
tYbZO9NtG641sr2x87g3JpgsiQwF5yRtcgM2venErTtDy5ZQSjvXdkonA4ETJmLf9Dw1G/prLvDT
N4L8vGQ1HyAOF+VBtjao3pKty3zv2RGi1/d7aq3/H4fK7t6aM1ooDEM4FGTROYoHUlSa0DbFjDX5
LtIRh65j8zBaS+ZMtlbC2HspLPDoYQQtuoKYinTvuWJgYOPS4CyXGFTEhpRcbrcY9sRWoEtNYes/
+DI7CoeL3AsPpcQiVv6MRV2N8v4q6Om+C8z5Tg+6oMWgBuRPR0lFBF/7SUlTPpmsaAJJGTqnBIIU
lEqP4LjAApaMOGLPAlXEcorR3gpgBXpMmhsge8Y2s98OBvFiTD7mWEuWT9xKH+Wyb9LdhZ0xA3at
Gd/3SIWYQRBymTu4S9xHJIdaoV61XQuxWaEbaZWL+BRluOm26v4Ds8cfepIJPLZ8DOZnykHWCA8E
hVL6mJsROPtaiXxBcX64LV8zHlvGgU3M3CVlUGa3nwv4aZoSqcijBrf4ymM19gGF6IjHXLSRVuPL
OUhy3wic7hw9DxGOFTfgXbqL/GcyiUNyPY7S6oN8h5ERhE+IKhQO48l1IjEGapY+owpoVaAWmR2c
hY7m9xCHegpLf/SvkZwgBSTK0rlLqCXsORm76HwClagD9T7iW5uyOLk8UWdbBkzieqsqM/wyV1VW
xLhn3EiD3V+CLgRyW8yLRDewteRyruuk59LWK6EN7IDEtH0af95uHKJwRa6GMxfAypd0kSf9S90U
HvD3lwkyPL1uwCEab2OF/N0ylPS6aTijJNSucc3X6DYG27eYsv7bQ0j5V8Cj3mnJw73Fxi4fkhVP
gZsO63UMuQZlHkirWNKA3pSyKLK9L3Qw2liW+rx5HXmJ965vAg9nxnEylDBO/LWOWMZBel7c0FWL
GHr04SDYl1rDjThR+W2h+so/nFWfZaPey9pX2wuhTW8amt/PL2REK7SYrsLAo9XTgNn0xBRo92ng
/Zct2V1lnkIbRx8GlJ7U10Cbkz1dArY1id2pvYB5Z/WxG6xPA3cnk7059DwuOeDN5WrVLLjDKDsz
kn0W8o7dgUpHp22P+/XrZpUIUC2OEbuI7xiL8sX8zW9xXoRjlL2Svr13K9/okzCPZTj2v6pdTkND
9TPBtTR7VbX1X7V1sal8hIa1mSzYWP1IHtrceLILTYPFHcbUqSDXMOC8PZDn4qrgLEFhNtoynv+5
zPl00NCC1zDZKisb9SncjcxoOWJuGK9urm4r2I1npbjTznFcFfRGmfGbElkeL4D9LdGQ+kXT3839
HGKsRotsglMEYNuXPvv/4nuzvD6t7Ym9CJDlHvxVBM+kj5mIM3X9qZhHOMYCzLZWIdApgy4NzYUl
QQnd1knJub+cGHfK9ek9xsa0/ttZwjm8jJr3k3sn/OMdN77bGeUks3DewJywslpR/wPhWc7aC0Jx
6zRcc5iQgwYrCvz1TXtNIQi0V8CPCIikaFnKKv7Tx7P5pUjAMQc+P0XsyENLZE5nA8dugDojwZty
McS5tN9iTjc6rn07CEop8CkcdOeaLu2Fpzl3Mp4wHkQ/zCZfnGVKGR76xOUBuQvyQ2CAXbpTVrJ8
NQW49l75EBw++t1iYnpIOmn30WOYDkGcRasogQiIVzq6p3w0DqS302or6A7Tx1JOe/EwHM82UOwb
V3eICVYOKaROJADloBAynI/4yy0nZxHQmieCuTskaQprgKydW23sUvw/pJf95vPLEVUrUmod7c90
QWGsp9pxKVHFIuJgvD0XACBFN5YNRGdDedytXfE5kogXdUIVWIWMBgX/9Ehe/FjM1fUifbj027Et
ofRj8GbnvB58ZpbX6mlx4KwZZQ5nyA2hPIGEJrB8SrpZ0MGfmdLUp2Ui5h8K2GGWlzOgp2YkgzTa
s8vCU2KHm1igsnOkFTkCG2/3lEhq2+YX38yDHsDSXBun1T7EPkF/gVHbmEgidk/PvXNHm/RA1l2V
u9Q1uOb3dbBQ5jCfNuKFmg5m/NZNxdYjJ2p6sCBo3QDS8/bqsTUbQ0oh9KYGLkJw6+Yh0W4aiD8T
0Qm+hm6u/Ehv79KT8XV4Sp52rMDjtlcUH8ADW9BmEknJXs48tVseEEEyek8vcz0zyJMU5zrdPhKK
ljMyLorccL5gRcHMIRp84M2o8K1lNvLfbUDro78HCx/fKEufLUXFeWW23Dg9Qtka8DkIkTINdGFi
WDem6QDTQkMZf7JvLFFCznKom7IDrSyfWFQzIafvaWNnrP7Vr9PVsaYhcRVR3hVdu/Rl6z7wSGPg
Mb3KPd6glY/aj4MQf0kpsN/EOR3hZiV5A+9I2BxDAREFTV/UxG7KMO8GSBWGJUnFuxL9N+RZgOiZ
VeEEsrtA6YTXx32vZjfhhUbciuqCZawwWvzIN/YwcA+EVRUpvLZPU7tIYeI5pus0ta2S7iosZdWf
WPqligmBw0wG1UCm2pHBmDz636tPaGDDJaSn4qFluKQp/vZIyiypF2B4U86HZQj7+NhwZ668K/TI
np8Fp8VQdk5g56oLiWnrR3egHcPsrPi05D/oUkUdqRiE/z062KKegtVZmHIVWVeh/9sQ5TBo5zEw
OnqsFPphhvnLoP02uH6bhc1mJfFbCDj5QcfWW0ErgyY20ZVO0eZQQQ29tHwIr86F+FUX9oUR/yRw
yXI/xuUykkEF3Qwnqni/mlNfOGZlb9d52KptpWRG3aYoFxEZeDNsXF66etj5BccOoSlttMXZDEVQ
MNCRJKOGRxkuJ9/2Ac3CLTKpOUPSc6AHprrHw6ZUfL1+wzZ0iLfh2Bf8ceGIF7Ug1gvrcNRQAtj8
VD/LXtbcuHOiQipzzHQ4bJnPXcKakDGpqy0NyCBVsEs3STQ4gdId4I4oUPEceQqQVEkcrOY8NEWN
SLDmYhrWZ/z5E70YAplfqJsNpvnrHqxGPja9oFDhPPPYLvyHSmnU+b068cP9g7FonEVWdyoc0AMQ
ty9L75J1d890OTIUxGc3+bmortzMxD25kizemvhNJ1+IqxjZji3HrFraV6n42sWFdkj/2WTRgiM5
w7cTwB21wd1evSMuEHSe7onuFN9Zed9lrdaXrrEvcr0wTCK3CTCpe7qxL1O3w4srDh3GycgCgF6l
MbdUjwVIMZzk0yE+GCPttXx0RezGTlfdEsIfQfnGL2CmGSkD5mxTilEMnAiEpoPvtD2U4V6rL8V2
cVGf59kbDeXrLe+JnWaQQHu9y54u1s+10TtxaFu1x/7UY3r1aBzf/DdNfh50ZU0DgrcKdj3yOEbn
nU8RIGptUm1yafQOILWvzIpzC4o4gqf6F3OwwifKihPWbTx9ntHR3tz9GMjFlnq3J52VwnNWz36D
PyrRtAUS9HVTOPfrodv2sb9b106zsTzuzf+ff0cFFEvOl9vb4Vvyvpa+004NA9y4va9ai8VGYvir
uB4uCmUM5C893wULgsSxInVfYOyZRv6Q/rTfanEpNfU69OiVtVsEq+1azy+IlfWXoxbYmJU1xwYb
WnC5jdYAqV+5uqBYPhFTHbKvRNxi0LviYN/mUjjHr/6J5HnlkuGVaKv7/ebTTJJmxOxDmgoA6wRR
AmML2umESvfGdQgDMXzzK/ZAhEFQLpXBIIpkM4elIQTrATc4aDCJ+a8GTdIBv1705/8IZugcTVj7
IdIE2J6V9Lcyu6xK+JZNhRkueIn5WXLhnrnbXT+tjnmiVskLJetQhJxZ2G7NHB/ITDfJUrrSz0FW
j7nU8caqDYWje5i178osqRSTS0nykbOcOcOQozcbSmgL2z6J+iRTNCC633cMdA53CfFTV3IMVo5Z
gRc3/igEEx38AEFB6r2Qc7WKS9joqut7U57UEh7ejw+fHAMvbnJeDNP7FkPvavzKKa74sNOY6zhk
Tpn2Hn/bjevk7LGx8gKc9kQ1DarfurFNA4/O+f8AAWbasIj6UpCreCgDVovrxP2/sTtszHhT2baA
qDICnzXDl8qxHGMH0MHg1nUyMHWAjeSUpzQovjDteld5vEdP5+4t9/9XziNUzuHWrBHXsR0ONG6s
sPGvL6FM50X9aUjo/sTbOUiBU00HeAbT73LmncN08hTTL0Wm2jrkKXPW+MSIvlx2gCCljcAqxP1T
MkVtfqn8La1Y0ITpQESKjxWJZhN3zs/nuaIPngqCpfglpKqN5DCk07fTpjIzxLCDzUO6LEtbPkK0
zhgi7xLjxnT6cc7yLW1iK+3uEViyWKc4pCk5umDNPzJouH+QHxmG+FobzgAjZHgihDws4euH80na
f+Sj2oZxFuoe/yrjo9K+ZYHZPTGsMeTDhBn46o87P9clQqOHjGpBntZNIMv7mKRCEFuJRlJEkP1a
p5F0X9dZ2Ixx01dWyxyKRLcQxeUzzfr5AaJySLPrJiOFJeaVXVqRr6lyJ/BAu3ccb6CkkAktFUts
eRhPWQS6Ahm9koL4XGnoU9Q0J80fJe+o3J9O3J+SdfQJHY13ES8Bd5JA2kjKHv7ZSGKcM4GziMgx
etvH6h9hLPIb2wI8GP1aig5glQrlftBMX1i2S1JYQsUfm6GqNsKztVVfKLQ9lezPPPtvTY7RCRvN
s3hb/LJXVNF5bkMBXXizymv8LUc4WoBOjXv6IR1hI9uvykYPBQrPtdWoiP1IKRbWq5nltl7w1fIA
HT3OZlkZfvkU+xOrsGeYOiEzuhE0zH3IWHsic7iLUTjGWV0l7WmLXeAQiJced9Rh86/9gUTF3gpo
KEN0VBb3SeLKc85D1F0tuUYi9EItg4UT4QA3qZCS+I3OXgmrppj4m649h+v2/7QLfz20Av8Nzguu
MhFIzKiRT0j0K3jYfP4DAs8INDeFJLzJSd5LHZ2IWLeNLteZSMVokoZV+I1MjWgfiSBBzdJ5ajA8
lsY4oGZMje6g/8Du6Y/2faDyVCgtIj04bXAJW8xak/7TUOjEe73dtifgVXPr7fJ9TLQomKCPKZB+
i0d3zFIeCk2EuTZZU++vVQ5eD4JAuz22mcXtLCNM8Ncx4cJqFTcDdyDg9jJAuxtELdp7CtCRXkx3
QpJT1xdWNKW1zRu66ibHDk6CYty8uD2uBF+sxImSZqHIP+sPkZzLWCKxhKdqcfQFehMreTsHOdz/
6fzLqM+DvGh+zOnVQLUun3CCFJ7z5+7kWSujkiVBjxcM3MXrsszvTAe9Lg+CiyC4GavtQEaBXNSd
6d/RdKR33cgoU/DuMORQoUM1Yza5o+dTXZpee09hJr3XYfNIOmjijdRJw1dCHbrYZQ31YLhr1gkF
DKsJMml3cN6IZNeXL0AejgTOc/zLNbWZ1+NZ8E0QuR/J8UWWNXIhe36rvtrb64hTt/dPja+lgxgj
HYS3CBrVHxu8Hvk6b+h9t/XlWDhirZgf79rSDA413waExYmNLyercDvR2lU7ZtNIsUdjU7TmfaV4
ppwq/L4QexD80lmbUPJT8cTLPzYXKwnRqBTVcjpSSpfx+T3Vwiy1OpIDxXmyfsyVCBR6mIr9vlwL
XQAZJdjbULq4Yf04XXreHiCekjKua4c8i7CZp0950WnVGK8/WVOe0UIsmvxW5+d2YzSl2NbCg5jx
5cSzJerwwo5tUXz6r3BdPb7I18iskFScxVN2cikJLdVlI9bLsziwyhxL3f01BfL/TdpReFEXFNK7
zOfLnLwPdmxnqa7r5SdyhBVHzmbNUFQmFrEv+0NTqTyQh/VB7OBPfk6r9vgGBg8BVTnfoJzbJR6y
fMwMKwRdIJ9VkRZCs+qfkC4xSG70ebyAyMEzjyjSoZwNN6LZ2g8DXl1F7Q59yLzCOyToxebFUuh4
K9totRKOUqRL6ZT1d7fISk+NO9uO3XCuwjobBaZh21CwfRaGrdUmxiZ9w51UJyClWWewsMDSmPOs
GPz/PLCOgTwELHR31WJzugqV2Wn0Vq4JUTL78A8hO7KHfhqE/Byv4v5qh/RWZ3uo6uXoqYP34Iku
uHuRVzHWJSAzDXpVK0tpMki4VTnIXf2i9lruYM9vyMDxavsF1Q3VLmkHOZCNT7MnUhuqk3GavBLJ
Mds8tF8eZJgtQqlrYdXJzVjcMloxtdA/UFgyRuPByIemQurf8CFj53SDnf4mTXo6etaXNdz6z27m
fIKIZKf7y8idwaz5yUFiPdPKY0nSpajmCr1Ord3c2+s2ufeSYIzlcxn9U3QlZbRblRQVLE8bz0Sm
fna//E2HzFcatAVssQko7XggVRjVISjtJkVKAnd6AwKK/7xejmxMtkvvDSEiaQQqR+I5tcoCCpaY
GLw4XZmjZN+G/LZDutTFQUDQ0Xcw6ZrhNGvTDU5XHrQYMrP+0njba/w+4dWVjSXs/kibdHQYiECM
oQXvhaGwB6VQMO8fCbLoJ0A5fpHt2ndHc1JurIDNCVnAcKHCmrTcADl9UEV1z5mF/0k3oY320gR+
1Yh6xhTE6YBPPKo+/d1l0o+saaT5MUJq9zl+TxwVqoC7x7SmE8yIAIfgpK8o5eE/HLMKmnlSQlUQ
tymd0Jb8K7vgbCRTBwqClabIKyEBgH+T5K1NQu1PxNKMkpzfW7AdhGgLdAIzcKVLP7sJQ/LWFF2V
nk2GSfluut+X57YfV/FNVZLUDI42RzQ4hX98vo++sNQcImBPrrtJuMUB/R+rsAVI9+i0b+cNU+iT
kJ31EoDZd04GV4UlJzHCdhhhWtYGwtYs6vvF4fm1h1IqtArFcy1z1LDfGqBI0UVk89iuPXTAvIiP
/GSoi1pM5xzvvVEDNgmaRWNZLfQcY2YZBiKT5WS7YNv0neFb0fBcGUTt12/azEjZ7kSfenpR5cAe
XolQ92PvXKBSXNTNLw7jFo4ticr9AJ2a5ujFqN1KSJOoZKU6D0H10gI+NeonlEmauEn20uB/Xk6m
DofYTbjJ+rQSQCU7M1+nHGp0x2PPK/WeHzhAV0VfoVEpcMi8P5Sa7+MCyFudykmnFeBXR8dT6ZXO
odWRClgBYlUyeqbYMeNQajWRo7LAk9bX9gYjT4tTVTrkEPXYXFmjeuBADHSUqcy5eg1Jpd2iC4tx
IT8wb4Oz2OZtmlK9cSVBogo5sKxbuuHlf/ZIW5lhkuuB2b0bK/msxGfx6fhCChOnD4Su7ItyCIJo
CQqe/v9JFwINl95u+3YoZJBwm6H6hPJxz/ZvMLppQdtS69yhP3MSlsW9k6nFPtsJJDV5JePztvXM
OZknHEdd4QnXcML+kShkC2UNtBpX+sbsuugKP/ka9z8yyPruF2P+lDt1Caeggf/he+ITR78kTf2p
RgeWbn9GiyogJrQurzOkvDluDp4pYOsCqLvVbu+PVGQng/zclcygRL5ugroUCZdGUvXDw5PMR9Ja
UnRk4twDSON5FLz6mWtw7tfpjGhDkRYrYgTDrmcKYwifYq3VrTaWP4QIyG2/m0ZRni6qaZHKj2/3
EICFNiW8f3wcNLbQLK0rJ//PrPbjnIvRC0XSjTWWhDh6vf76QW1ZyCLsV966hzVC3gc/p/N7XsVd
6xMFCASPt9EtyJD0sn4Vop7f3Npp320ISDL7PO9AkFxYi4E9Vrxkd9KiNDUSzRluLu4uJ7khI/cn
pBeRlHUgIO0k+vTwpmJ63Ynpt2Kiebmn+NG8w9IKBM2HB7WDkiVyqdfD20wa6MP7CdmXQfzCw+ic
NjfPnmotN32DbArLl9oWr9gOm9jsQUTH1Eg5M2nUL14yeoxmfNSKSEY50jwRDJZ1h2iMs4rvQXa+
v/GaziwommJxucRX98iQSU2we2He1KXQs6NcCxN7kn1gnJLcdwpdipM1NE0mxIaOtNmUhTsp4ifr
jQcMmWPnR8CQoNuIjTaNqLDObZuJO2CfXujE/HywW+bRjqcrcxs+cbbq1++0eJxiscBztzBJyccL
4OidobNOwkWJOxshr7Bt8NnYUBNWPl9F+Xorj/hk9fU5Yis706aafhOoFelnfzXdtIBdSCWXRqHs
pd4nwV8ijth0mLin5cCjYsMQya986oMiSk6M9FZkuOYqhiXHMOtNmE5VGlzyxskPPKDjwf1L7rbb
wONO0BgSDYwD1z6Gz6KFwTbZCMvC6Wyt+2SM11kV4KFDkaDdkosM1IGx+2qRvOD0UFnr4Ue4n7cR
iROQRSymuwwEXeHNxaJfngw+vqKDatzkPI/wfIsYfn9gPwrpOoBxT80CgZgT4/6UpmAekIWgrf8Q
yDD2z7bsklY9x9gmMzeMzhvFNs8GMHXF7LKb/Gn2svc4h3Lgm88zE+ksAGvsX0aVPn+NZcl2bBP6
t0JcZwj6XNL3QbTztyXkMm+xiKn+KW3nrfYNpCFA5Y1o/0iXLTScAKV9sC1tSgUYE2mE9fFxufSU
6PaTrQcqOpK1QQCKRWTSo2tTlvSOuNaO2xzAZfLgZ95TJMl1QFBlXO09AnsLkyhdrVVsoVH18TDu
N8JlS2szTAPyyjV2aA97xiqElHqs2FbZJEg9d89oxTtaHFqJlPNcMnB4NAveXN5nz21ajBwVRkJr
bbHBHSp1Rq1SDkDXIOID5Z0sA1z9tnTmpj6EWfktcaFD8K8tvzN5sEnyImc0ZrpMr/B1ew0t/KRb
TD8CLDs2rlnd2q306zEZFE+EOj/aJG3i7y9RK2xsEDpTgWvD2b/pmi2jSZDJT8q4wzAKLrldM8jj
M2Tyuf15Tl/n5Zyml7qPlutVDtLhBmYf/H2zu0/URAaK2gAhZn1hROxlDWGpaqw6kuGwagdFpn4H
aXavSLcYeS955uoRzxhD2hV39X7L5Bm2OwDWqT646VP9WKMoEB5XddpG34R4uXM87c/HOdWhkA1D
WMHYR0I1wvFLXF+LW2V1JDhHsVB9mhLZV2nSA1kSBfGaWXsQI3StRLqkgiYdsIpJpBkm+fIDGn9F
KJrNvW8DNKSo2sMpCfmUkYzfaQ9kU2eZrjwQwRxuOghdF5AT1QN8QBQH7t+/7G2QNjy5eeHFUIoC
q6CP1uEfW9vQg0Cfb+hqG23dqvZuMNLPa1xfbwhNeKU5+kK4YHmdXcQJHwm/J0O83OZQbxnk5U51
rmdc6Fh1Pt61Eky4WBl3qjzrxZbgI74YKWiDU3EfSg1z0vhAiQsTIEn4G7nyJdS+thShu3mEd8s1
64Lh+pygatw5fT+66UxR11jnOy2/qb8I3WYoTtZS4V3c2D5fmEg01YDocEzlgiTB8cM4+8FwHjym
mLZ83fRCFfiSlgFeatr3d5TxCq1gsQZMCk7TZjn5HNQMkB41BDOHTjo6hio2T0gxOzgKrNQ+pws2
dqLjl4WoIU00amJA2JIy6mC/aQADHwmI02WhZzGYQJ/Bs2dF71k3aKY235E3R853jKy7tEZH6JC0
XQZvngBWg9OaXyYTwzIKMAyMa3s3pr8Fvnm/K910ks8VQyTikq5tHZkwcHsgZpedSTES9C1Pas6j
+asiTQgR4EAJqhgjvn4L4yJG3RLxsqmF/M5jRHk3X2Zwbt2b3xDGP/zCmUWarbGKiUEW7doWTPLY
caKASEdh+qQva3Ii3QBo3hW6qekxze7EEI7XFtUi9fVOl4uMIJn9yoznskDbv2PvMpoAlpbn+RM9
b96Uad7JcTRr+LuLImkwSJ8vVP3VcbZestoCKahPFqL5V7iZ5QXY0QJTVR2R2kzXkQbG1zo5etLb
7zB+rabM5QjiugmARjpZcXI8K4GrrpiyY5E/o6jmUjrUbDQOI/t2rEYUivKwKZ1E8Kur6UdNiZ2V
s1+pfyddlER5/oedbtwpLH3prnrkw1WfWMt1eczXD910aQMbq1EdBRCs3pUp8+nIQ0h6VwxUyVLr
tJkiFcmOGtBCal4k/UfsMyM6+3F7TsJ5l3jJ2IfTC0VOuD9jixA/E1rLJ9rB7j/4pyEBovQXecBn
BMTmoZ2VLOuEOz0wdAYyqS2kaC0nJHrMWAOVzo6RZv2HCVX1ZbjmBOtTK6rKay6KvY/lbXka2SS7
iPWBhjIS8040DfTVo0+9shO/0RQJIG41UYS9vltoYg3cFqlQXgRsTabGTjnAN0tD7IU7QGyxzZ7b
568BuipPp67EORKM8MeW2POwsYfExOOZBMqe4KIP3+s8yA72fGfCL5mm0XfOQ0cFO5/vXm8nLynM
OGR3VPjZH1NBcUDjrzv0fCaKk4uaMPmK4N3AYKjZw2ze6mhcHqM7n4IKAoEd55kqMZN2hd6IKFi6
tNF3faL5CR5llM0JcXvEqs6rfFqVRp7Qe/Y4ILZlk7rKtWzaguw/YdsyxJ1Ze+3gDHiWjhGLRCPa
KNkpzIxD4WgKp2NvjheFBBXRh6QMTs1eSGxmIjhCKd5Epp+HXoYKmRjNDmHm2Kkc4yoW3HJYVkqk
d+obUd5wfFUkHCcTjfhzpsJTHMHDOKEHy7ijQd7vzrwCCH5lHxiRqBKzQR3NhHZJvBpgbdhfhF80
7I3u6usz5SNMuUi8nr3zcRWeInWxHFwvjQDqG88e+jp0+N2nTMpTBgA+A/R6KqhlpdApmVPsdsxy
xc4KQxcIPGlql6zBRB3MFVLkWcaS3YGTPrWlKFuxpfWqpc8R2a4iRVlVaAwIlyYWTpdGcnGYBr/E
MXP8vwypzZ67txEgsyD3yd2YNDXJWNjkPrw/2kQRRV1Zkbt1zH9pKxyGoUmYXZ4Qlr6pdpxQI/f5
hTEbEfFVcudbnRhBZmN+5dGAEmytDJjZe4RPj7pFUyf98DNfZbXJv7DJXXUjNqvcrmARhl313eHL
+s/Jd/hbre/gZgfyKjx29Mu+GuUe4UQO6SJlSa0PEA8q5L6ig1tA3blX6zkEQJ7iOEEJq44d3JNp
0OKBBRIlDuDD1GVrlEetRWj41lsedhUXvcN44fwEzBUXn8PHN4ttU66x06v0pEgvAmr2LHn1gPl3
i2HXJla6oLUUblL1S3Gbfqcd+nxPKLGA8SxKFyQ1q5Ix71dtOcEW8uHNgVcMSFuoDzOSzgU8MEra
bE1GWdjVsiIsPAqrMGXkIDtrexq3JH9qRp+AqpmMRX1KbN3G3CV4Q3W+msqIv3kl2w2MjAJY4yA0
5heDAB5aFVeWzKEubIfLOfkgyd4puKMIFT+lmp+SS9pcTiGGlMDW9y76mIfRsTvUdZUF3IfxQimC
I+9W4Yu/9T2/cm7Vzf18j/qHuFT5++pBiG8SjePx0FMt3wIdyIOzBEpTYvYAmo4C8MFbD8r5mhRT
EkNWO81nKT93JMBGjb+hWtX2gxasws+B1DQwNinImEN7zZUdQhElgsSePCXxFW9+qwBq3rZB/X/z
NGtYJLfiuN4gglcManOKMN/ki4wrceTLGYcCmoDL6PWBd94hTEYb3NEAsBnogVGWpWW9KcnZ0Ane
wDlGY87sCWtl1VoZH3nfeTR3y3W9/tUZ5WABL8Kx/MEyki12eBLpij+sHVFB7Js9ieuMOoeovP9i
lkV3kxThUfCsRAdtaK2PKJnh8+kcQBOzKjPCa2fK+A5FuMj+QJ7p1+UytnJ0u5j1ByFxIFcpiSa0
PUMarCXPBBD/on9NVv82bV2r2al+21R5aGF0nQzQ7bjipwlM/kNSYmMplxPE00Yq5/WysAo+G+r3
4o7H8WbRg1OvVJpWA1ikyiSYu+JInjAqzkLlLlqsmN0wSsPZixbH+sRL8C8kyGuzSelt3s1fICH0
e5Yho3A3qcZoX3N7zC6PRD5W6GrzRcw3VEHJ2bqK61Zr98sRWcu2YCQ7lmKC9I5EB+RDL2UQGSIZ
K1D/I4oGWFEnkhoU0HGFP23NRVFU/Ci3qhj7Jeu7banY5F7MvBWLa31LFYzYVFWmXsjkC0jHaA8P
E+huuTBqokd+uRMo7oh1mEjc35TnD80NUD6vvW4gNapBVWx+z8c7qmWcJk21iE5/zmQGfO8Lc+DN
EUXd2Xvc0CHG1AM8xWtejMbuKpNTaiMHrNol73YgA8YZTtF9XivR6tm3lN/VYXQUZE7NyTzdrV91
sE3H7K4ydZyaMr5aGeBXDAZIQqdI6LzJJNYArMlQKYRuSqjgleZznnwSeC0XzxlFl5GxpgWfqulm
FXxxPDrOk0KSsaFsCJNapqm/GqSIlGJePoddD4klfpZohzVTBoGayBrT/5zCoO7tYuDUD47vYHZP
cNItE+LLi2NZ0F1Y+SSAX0zA23EAVTfWGj1Kw1oNetjVMH7tGq9RC0YKeB6/mzGePUFL4B/FPZfG
G41Yhb+vFaeMctVG0CxjLfcZmo7KHUkR4wXHATmlGYAuaHt9XCNRbTIdGeRcICMKSY5DlNcpPTLW
BrCmaX3uaQpVvatLeYwN8jYZstAku06tLYgxwprUd8lnVKsxdqxR0F8ZCaRJcV1r3P5yEmpp/BTe
bWV+Ezc/JdoF2DGm9wKCklTcxiowqtrir7l74jg/BUr7G2Rz0COaES3uigf5CsIUttMn+6FPJtv1
iStdRFGwN8L2cp/KOPBoX2HelQ4fJx6Xj0v7TqM6YhfB/BPPOwnSfz4XDKAM07dn5U0rKqwvtQs0
Fb1CbVjJjziaZr7vHYmW26BfmrTWlY039u1BxzuxOQtg+pgDfrcjIdQvdFd+UbCbAmblnPJgQ01n
+odBUfceba0U5KkBQRWt8GUfvV5HP+4JDOL4OYNqcbznbF8iCvVBUMPG3feyDA9EBKFclMsu3bqq
ILQN3V8NrsNYGwEIaL3eVmTb6uP+6ONC2zpzIfBrGamfBari5Juxtp2J2UDLDk7gBlMcRm1Xoozz
LYMvCpd3fzeLWpEr+fsgnU119Eor4OWImK8Tflyy2Vp6bVERYowWQrwwS9ARZCJxbyYE8mx6mgNJ
fOgXwkO/eMuEw9d37Z+tPpvYV2dDWlshDJz/SvHu7buyaqaYdMQVJ2CB8Rgdc3W1dDuqGvjUEWDu
lwx8INwI6hEdxpzGPLLvjUnYNSN1IrTPgQWOxkvWNdLyl+loY3LsAGX7w/C5AvJl3/zsPtk5AOT+
mhmk+Z6K4w95cgvPCFfcxw0a5hVc0rpKMgp/k3X7e8scBprx92RhgsKoxRw9uvZ8E4uE0I9LqG8s
17MMLJxEH2z0Pq/fNztuGS1Xo9t9zvhRg94Qy2vHKXlk3jyCzpIWOojFqhWA8XGdr9yo6cXTxG1S
E9brxz+gp+Sm6XyadvUOCV91oaSk4lfE9yo5y/vJ424C0HcdowL1qOk7PSC3081Zx+TDGlOiSg0W
A7GrW1C2eYooW/HczycHr9pj71FyMZ4lUMIY3mGsFVe8tcE6xHG9j4eawYIYjSP7VwCIQIe5i466
tbgXtwWV5DoeZANx/xb9+LUtx9CTYoLutEJ7PFylnMu5sVWTq4aX8C2CKztGhHGATDYBE+CnKYdI
EJTQFzwR03H/KTV2pzSQsVqJC1xSOSLBBj/ZSO+wqk1R0yZA5HcI4h/KUJWQ+uvg55dj0WdbQfLV
PtuixbuNNTjQtljUzw6X6F40Al6QZQ4R0nYb5dBUQTGYZacpDpwjyhCQUMgSzkU4rbRhylGDG/NA
BES2TznAwyjhgmtAFK0W9qPH7UAeEZWSUToxNV0GZKHUNb3w2rIZ3Z29hZ9pWcZW8I6LUpqG6qvg
Pxr/rHC5m8zkzdQvlyhygAWrv2xDDjRuXC4uuDPCHjqmgETHVGH3Uy95Poujk3xyl8bMwum9s1hJ
KH4ZjF5BVD/0FscqAuVXXP/ShBv/CDOFUmmNzLriV5GgVw/BMEE47VtHB4gJbukwEHFkXMxV/gv5
gccFCAu6JCo/xb8iJ4H3smqITE9TRSBjrkzjRVjln/U/zyKIdUhultHn5tYh7xxjIv0+q+LFoEFY
ym9BOTmnuhrkyo2b5cMTqriO+Is8B+iHh27bSUxxAMJO1cQxn5/XrEw4flJ7N3w+JxawViPTGkF9
xLyuYeSUhxJDR+2FYE0ENgIQZHmANSG8LhmdU1ChjTbp5Cq9UiRCzVMnLDGrm5Gpk1NzYWzmwny7
5OBXByXsl2jzGPLpKaIUWEF1UhKLXEgdx7/dLfey6Hz/MOgFGdeUds/fRa4j/UPxXpqL0N/tqPS+
HzafV+y4ACH42pnBxKCLUUeyBsUOJOsSmCZGEHmZnbwbKtC9BQciidJMQJQWv7aMRZy3IKGlbkCf
uumgbqZnMB+sfHDNhlVv+2E+3T61q35dJ2WBD/mHjYreWrAnc9L3b5lefZ68RXc9zZT/Sq1G1kUW
XQIzZ1jC0T53+x8RbnQJ9+MfG6sQm0ss8HutyNx51OgHGKHtXw/Jj1GMO0jZxrx5teepJYO8DR5Y
+XVaTwOj3mEIPF3xj+jg9Deh26ViZq9xouRQb3kTXjM7YVOz9x8p0OizUsHfFixW4KRxwW2zfWcJ
SpRD2+LQX2J9gWAx0osGDr+nbJ3hFxmsFl1ovStp2AGNryy6bUzGQy1TXGSUjmnbUkXi9KIFH0V6
czoSWJKGeTtXZigM45yu8gAhAEs0EGEw7bIW2t0P8dh8d+8pBexIjzgUJVMFJHSVoiWt/NT3ukaT
3Qg95PBHxAtuIgxvE5R6pJH/H06tiE1m03x8IJ0rvHRlsb5vGT38Qh+xXCzEVaxZ8xb2dRwWqHNw
HjVplWdYA2tkIj41B+gcol1MRM2BN9Ib7P0tLCYy5cqQSxOuWc3zQgumbJA2P8FHQ+AktGzS7Z64
2Pmx8P5MDZDMqMwIuLBHzu7xmzeHRtfZFJ91FqafAtVukaXWMT8N0Fwx9O/xi3f8HpLn9cQGYQmO
2Hx4h7DFref0KMwz6koUlLwKXAVALdBJPnL6cu+w35bAMG+o55yCi1kaxdH1nOa8oJ2OzHjkXREd
9dULShV1OO9vm7KLM6oTUZKjiocrFK+ItstKNFwlZGRDz9ax7keOTB1CQzvCBAAZlLi/NehPvCN8
831u6NwpU9AtBgLBctuI3Ccnv2V9caVByV4vk5J/e4UIJ0Dew8jtPBWX6l13vJ14GnhZP145Siwi
nvwNX/Na2gL0gsMsFeQ/hdyierM0pjgduWXA4cz7uf2Udtvgtw23PUpB+BSsZgxLdiqa1BIfpXQG
fkdNQ3JiUBJoZyyiMPMgHMscU5uKLIRSM8yfHuaYjFJOnWjscAVwX8NRxXCOYHYGaULupQ8jAKbJ
s2uzDF3qKj/ZosqDEdWIOuW/5BqH0CLI4rjL/Z0av3KOSs9/ynJM38m+7qcndoYvgP7oBVuvXzZH
OpINRA7P2K70n/jXlPa00FRKVRp5XxRf9gRO/TrCqDEvol0vbYR+EJ2/luQICMHC/MrJJYwjm4+Y
Uoew5fRflRaSp3PkNtLSmyAUZI1BATaPEVTr8PzoyZWwOA0WapmiOtzV7v9eq+m9NWMFyNn+9M83
WIF7nJNmoxjhqn2BEKqDyegPr+HkIz4cTrgq5nAXbddu7/xJdPzrsqZerFGpqab0OQE61ITNX65I
fxSNVUPJ3yW4ldy3t761USDkg2TmCo5AABDm3R7ZL6g8UGRaqF9SNUBlOtQr0RsMED5jyJda6KS7
q5A9mk9Uz5I9odAF+4Fo6Pwu6RKTQZCx3w7/uVnr0rESqK6nrNgMVjaaBaay4/xSEbX0QcZkmbxJ
jWGemqM+Ty1DGVBCD/HB5pZHbduV4qi6G68LO7GX45YwsWLJGMxYLxHhmJdKknXkj61VL91v+TG0
t1P6xfrF7+JuumtVJQCODAxfwS6urk+8mY/jDtM7i0LxJZxFuj9FK/+FnNBXcCcZcqyyTI1JUzaI
Qyfeqt4P75r1hMCS3/eA4iPzX5SDNl0msdDCGzuQSwRK+IdkDBAkRsNYWg5zZRYJpz3+EFZVi3ZZ
gUDWLM/mRzahbQPGOCI4RmzVMaikH/MCFThewvDodI2WMLgwJJxPZ2cNZQQWA3TrfUm4fQTDohKf
YIjiTu9hCN9RrlaR6rnERHHtNkynb0jOdG586QQ1VryukKvJRJNU55Qx/vrjYGk+O3b9lnggL7sN
k5JjazX/eJzGxGDcyN0oQ3fyHb/QsHAGtCOyt+jdkyntIKJS5+i8Pg7GePLlT0CesukdqPwQlvzQ
enLhGU89+vSGdrTW1yjyo4DiS0zCiwXjs0IhwpCHFEbqSxrkriatBFZ2uH4DkGuxu6VIAGwxjYJ6
3fFdJMRS0fJ8mgNb3+O5OAPcnVk/wFol37FSdnYSfBiYeO4eR3UOwiYBae3gtuf4E1kgJqzUczDn
EAjwFn57Tuz196fBOeQXMu00mBOa2x2W6gTnyc9UZeQe2oUbc/D28+AcDTujLpWyrYPrizPzTY4C
I1PmNesV2IiSjrm3/nzzAZ0+9wK3dLsCpcIaTa3Zm040/31aGPEfyT8NrHHHQRM0zQYr45eEqPwo
Wzo5W65D5QGq05pRa2KVLZq9M7o1UTUlHoVX9BSU2tpOrTlknMx3Bpy0JEVlThfWrn0PQXTIo9Wq
riV0jXnbYnA+pJZ6Hm4xRe48mSfxk94xVYPMn0/XSouuJslr3GBUg5yqMT8d87go8u/slL6oRtLX
4QRjuIE5RgiE9cr/YeRy8/cO2+C6q2NdBu+JBTYJ3dis4kSs8drhnLQU5jgnm3K1OpxJkY3MUC1v
Hg3imIWbv9zIVGoYNIQM7kl3YTDjEYp47zPHQYbY2m0y/kCMLK6CbHKu5vnp6xgQAmyPfJu75a2Y
5yXiCbBMRyHKyL7d+cCy48qzWjeqzJTfsw9F9mBhdyqvIKwpoAdmfFCRYO5cTngGiwXZTegf0Hc9
Q1NhBeLGUl/IowQL7wFLmby7KT26t1LPz8saOEm90ZhxczBi95IBOPs5k7oSxuHelQf0Kwrms0fr
ame2HJUnhFE1M4CoUVmBwMFJS51SqwYOGZbXdtWtbwM0IMArv6s6SVuWFlCTB/uu8S5mylikdotJ
9aTO1P+H+FJEbkFFiIPEoN/ZUn8lhaCQ+6caOe7jAV/K/5YnvC5co61RwUDaqo80AYbyIkEgwHru
FRAIedMKg1fcn7oGaDyB99xOva+K2U5kimuJF6PxsSTQYQY1OUvXzodEq4Bpjn1O6Jr1yi29viru
InrR/1cDZPOQL7JQVLPDM+zgUHjn05xgdQRac84lH4SzbxVEJ1N1J08Xv1aX6Lh4tdnbfLhyPD1P
pFEHWbIraqH9ACFdkS+Axa1a7jIWL7h0/f3fWTSQnRiZmdwL5f2oNbhncIpc5zQDPB2ST7e1sgL8
Xqsz+3LCAI+WTLXu5YFr9sEsyRAlk3ukI+FBGYlJ9wnZg1BJnKTT4nOdBcfN6954CIGJqSjX3MzS
UrF0Bd4eHFB8VwPkvvc4fVwUT/asLg2/ia09t3v36KOAbHOwFyYOyhbBR0EBxp3rhliIM2NRDDgC
eA8yHUc5igd4bMD/SxHDxyDthjZYLHABHWrJtuBeKLHsgQOl38dAWyC+kyq7kM6Soqq4BF0hjm4X
gdTUtI8amigfqaIiCc6Es1lLBfr2IWv4MyVQNUU9rAGiGxhE78SqD6dOtcUs30mtUftBNp9+0UaX
jrvHXm5SgP8C//ZbUW+ULRgqRi/qftP0EgguFDearlVAitz1AWrLQZXu3tk/aS47SUcP2tK9bAHA
P3U5/I34ci5IRE81gVfrOUtLQsXbLX8RC0zJuEwctkM9/hv3puSFmI+CkMsabgnda/2XLB7AAAcq
rJjw0qeMcMsiqFUZIYWtO59AwuDjV+ymTesVHTaXFxSuOcjQvhvOIig9Zn2c+YaMw3qf1PMuB7F4
/yrKEWrxpW4ltuiC1xm44MweIEVydr5TZBiYw+1Wz0AyAs6y8Uxp4mQnRFvjyILCIsKxQqqXGvQs
s+1EvdhfCFZNst0UoWKV8DVU5UO7Eh962GawnvaFU6WIJKe5JM0tTNooCWXutyAWDniHmzcZLZ/s
QzpUTp2gbJdx0SwQD3ZOjq29b6EimzoE8JlxCMYk1ro3xQrR/TPezGLDJkP5+VprNkXVboWA0Z2R
crHs3yI0bpP5GfyyA1knEpTJhQ9f5uwSQReTxr1TlMa8xct7XP6DAd25ljzWpqjkkPrkIpH2U+Jr
x1gX5QT7EY0oBF4C+qWf15i7cJSNo6vwcIAPUaWEtKY+NfdKZBPblPLXIIvYV1GfwtEf+UF/pv85
7wL7nFOBydJXhlQDFQplfg8E9GbO/UsjzjAsiT5wUcB9iDw8BnhHO5WJA1NSAS+f4warovrBuU18
aSdKETUrGS49fL6bmpCWBNCYOalnXWvuFmx0Ji1EjGfuC/weYQYqZwbUh1+wRh8l5qBGEzSKxdzr
+mW2zpXwbP8Gh35PK/Tw3zavGBc3WfuF3ILso103Aqs3nI8Zvy5bZszXYQXLZbdMCVw2K+28Ncyb
9NBKT0jtAn0FMML8UIwUB3tFqzQh9Ewqj/l+nWyngA4hIpWSWb2Cbbph2q65OLOXY8cXy2fZWfhk
V8gpgMvhPMrCBeNIMUwa22pb57sfuTe4B+jRptOlPTYq4wccs30Gfe37PXS6s1Fdw9YMI3fWYJOy
IUzauQIMG9j6N9NiIP9IjbisJVRyE4TKDG+tBRX0V+Y+4iN6jZgCk468o3eBKLnpahSm8r4LTyxV
OC/5tqLODrP6gK4POIOK6LoSf6WAXjOt9ZH+B+JtPLbES9enGvYFJMnOouzEkpS25AzcVqAOYVJS
VZq84zT4nC5zzVdSrt8PaE31niOpXFzvFUhT6L6LaQ0H8sLNHf2II4f2+K16if6LGU2zdqM5BVaz
yRjlpZJF+tAVc0lItW1j+OAf7dhkIby2OR9Q6eCrwbMGtdpq2W7S7U9pYd98niRyjQpbfbQSMoeS
iwQQ5wWp2fMHFydSn/9wPIxRT2eaDqUfqTfugmh+kaVsF8f0UPew465TzuG+Me7Py4y+nDwDgbjt
j3HMc/9KPpAeBxsnbZfl6Xo5le8waNRrGspHelA/eAIaZaSJO71JCtssjOdds6Odb1TSo/yPedAG
RY6OiW0YGQ6YCJAirfolEfcMPnVZhxcKrKq9qAy3a9tMOAlmJ2uDzjNrkCaU1ULd0ModvS2rfcYU
m1+hzf8rXaWWDIlF6kWold+GYgRkq0a2CQn6oykAymHeFvGvGm7O3H/ZgeWbELf+aCTM4Ko7U+f2
/6QhJrb0a7ZleneDz3EZLY4OBeUAih39DGRp1eHYT5h78QMnPo7S88Nb75f4p6fBmUWPRJpaMVnJ
YBu4frCmmDWZqt11FG/E87e1AvHlMq/vGIsaj7JpTCNuzHazHUMa2lAK92fjZ4tW6/m0Qy9r7YqD
0GaG1VKQ5FHbx5gWixoBi9MaOCLpded8BYbAOMtsiy2IsAeMKmm1iPMcsCrwpPG9y77C0Hq8q9Hf
fktYzgkSq77gyIT6kWWF8i+CdN3Iut7CWSpooaHNYX7dsIjDJU9s97ukPdEonmm1m73Ty5lvZ4vk
pqUEJ7BS6XouZ+T3EzNCWTty4kk8jE+BG3iF4zTIXsZyLAN7D3iH135ABQLn54W5fl5TioDIUTJp
as9QORhX1T0GW96B8dDuRVM3ZaH//B5CENTL7oshgBYvmxnQn6RROEPGJnkZDu2JLg7StDt8YPvX
TwkNCmPSx9zJb3buett8LQJ9QaQ4ZXDxqpRgSd5lL+4F1GQvCjHRSfLJ3kTsKDAxncOPd7Au0KWc
YLw5cAOFPFGxvO35DVyxHZ0AhzXgeYbnfak16DD4SGxMSQAyP4SZgkeiwWfprNu2E6sQ7hOj+/rA
XbqU0ybXMik4Nn4RrntTo7rhjQELd6RskEAGVyKFa4MkOXbj0Ff+ooGSM6AmbkdIAssfPA0N1siW
gbO/LMk/imPW/XUDckJPIHZl0y0n8qmBL3hcP/GLC9OyJmMF3nuhhi5vP/A0WTxWGoSROT2TUBAl
GY7AFckLFGOdt25adk1HyT4V87HLex0psfaM6ha0ZsXj2fi8UvxK04hQqSfDIrNuBnbDfNTpC1vc
weXkq1M6n/eE1mgqUFq4B52ys96mggcCa+36J8nHboNQLgoYahQAfFevBpwo7u2SgEUirrS2z8y8
nSArqzNO5HM1PZhyyDCs9a8sSIeVS2DnvviCGmDjMS/DkssYrbs/auhbsp59RmOXSVHw6DeN+V2o
mPd+5D9bDZKptQhd6XheZO5o/3qET0khX+TcBR7tUEWzH7mqj1eygWuSNhDKHcmHx/qWoKs/l6wl
7aAN6cNwtgeIYJK5PGB1KPdIkNPX5Z7uuy+lk4j73B4M+0utspyFmDsKT9CtvaihTgr/y2E3FiI+
+grBoxDCa1zNjpuemxROp0PqwkjiBcnit2SqYQxYgTHPCZtSX8pPiPyiUjcugAPrZVQ9nihIorKn
Ugq/UHbtiZfuWpV8a0syf/l62jLIfc+dhqdHMq8On6zmJhkRDGW9g6nRZNOUOWgR6fdd0IVsOP+J
3J1eA+wKjIfOvHcLpGM0voLbWVU2dJZoWvDjeH4AxR3oH4ED4xHEpBd3aVxuHaFnKN+KHWCe7jwV
YFWibIKfvFTWeIr0zqzkpFp66g0Dg3D1RdTFlSvYgHCOsgk7GTzlGMQ21qpSAXM5OSq7m++K0uNh
uxYHbiphmHbphf55Fa950zvv/AHiNZ8gWtN7fz/aPQe2ybtNFRh3QZyG8h3+i6DVcUSOxxcN0PXi
nWWUpyC3kkq3DiCpKfp1Oldh4EBkMG876nT1ltGOX6EJELjGCHZZKY3gsXXXfBcJ8hlTKCPsI8Hw
eHv7dD0larK5RAJxpADLB8hFQH+/RWLxGYAWMCEQfBvpgly9ma6XmsT5UnvGNwSV5QWC2Q4vVmmQ
9qqIR27yOzzXXjCpgVS9paUOBaZMxcWFfFXGcZ6IhEHee9pXZW4uwcLicTN4N5/zFEM6nvNdIZt8
hEbnJMDFjvYK/HCCtMRpQF2lBdt9mdEQi6LQyXg1pBq09vPnm4r7UR0uoO9iOpXxWp7q+tGjGzBZ
zh9WsRZpMfeJSHY6A7yJrXgUIGouTa6RFornBDpZwMDwd3zok2zJPwtB+NKLiYxjXxAus9BdBl9y
EpQdd2umd2YzBUArv8iFZSPJcRXIoIYPnw28XIHLCyD8rQpWjg/1aW7uaQYyACdPk5z4mvKrZOWF
CgCq5Yp5iZUCLic3dYx1WwEyrTYw0QrI02hX4dSTtUxfKs5AZhvBXuVI83O3slhKrDAZziGyZwzt
tZb73ZihAqrYivaHkVveqX8+s2cyQPyKHccBH71PHVaZqhNl8I1wEt9znqtp7QUnSKpO2vtXBC3O
1FHBhzYnKDrIo6ItylCHMCYXG/qiUl2LsawQVYAUOMG24JCAmB5Vr++a0aPm2/PW+022HIFJJ3yT
vy2h2wlsRxyyNrIT6DwUiPRJrfzQV/HW/d/81gLJZkq7bCmgFjKknE5wZQIhpwOn5+CjTcqjSJaw
lBNHoZ+bt3lG7acCJ330RICk/P7PFkjNDAJjlpvL5o5mpbGL9SSCi+icypEzF7bV0w9Yfygd/+rL
+g+3Uv3G4Zm/k+xN6KOSKh2FqwXZE48lmjOvKFfyWkYlZAy8GxOUpNdHMw2CmDmtHETpb1vP8SQz
pdXgzC3oSX15GCDa3SjHz5WQEulGU8r33bcZdPdMScWyFOfovIIt0J3jY5Lvdv/PrwEMbXo9m5sG
nq0OuMU7iHc09BPE/M/4qe+YcKgPZIukyYCe4y8+lqYzhCmHVnkeG4cx+gLhxsCE67wRXBsoQbv/
mm9YqEb0GQUOtXWNVIh/namZerA7iBTdw+YfnYjZr4WCI+Mijx1MdTOMqzzbeyQzzov9tSI4LoVF
sbdpamUV38saLrmQpuRAUDdq5KAudMZUYgxdYNKz9radno5kSt2DdDCuq90fOowkhJdxYnexZv/M
4xvARoncsAB1DaErdUmPS31b5x9f+uZryhpoxWV5vnz3JNcLWafjfxuecbuBNxedjK3eV9MD3J8+
Zfq/FqrrGDnS9AqHlnu252zfEz4pXP0bsvh7iRvJbd96yzYEvVKAkDnPJ1prOyCclJB4KzG1JhwX
qxdXdWV1qFq1dESEx+i684QAstBnsr5zq/RadTVza5DtxKkCIRzr5fFzLj6B5cjUWpTVzxHqzhTj
p1QJ+XbRgpLWZo/rYNRYrplA2cce3rjCi85aTlhar95r6Nd5NWMFhtBL8DMawAMF/AuMbHWnUFGC
FVgs80zMnNnyg4q1DrKtIRGohjjYFB7J44rthvm7LZk7WHqHGKoJiysNLlnXEpLb3GtCSeoKBqoV
ITtRz5MivpCpS5rz8EXHfBA1wJnHPs63PqraRFwAZYzw/OsKtgnbFAqlUESRpiWFW2/kefu5NhtI
VYQxHKixAK4jl3nUny3Qd++TpOQkkVb5MHkvv+kX4Enq9XoY3oy2poQ9VaNNKzkfmRYXr0jGeaS4
uhDUxm8/Od0CvuhoVOmcOhqsh1d2ISnxKVz91aPEMCMcjX7RDL+n+y0ScaTziCLo7LXuSenbvoll
Mms2TN1jiBllIUG+qqlx6NqXUuRPYC+HhoYlCcCjB65lf1dXE9wJ47a8s88D03VZrpMbBBUYoWGn
LO4clCBW7kF1NJ68iKcUnIYKTDiVlg5swuj1ZRfUfIIoYkVc6no8S+S+XYMWeiU1uZAxVysETVgC
Ff/K5hEuL06CPVzN5tvpuRHKp7nl9conq5CfSOiTiExjV4CGu1+pPBzW3lZ9ZaXg2hOZfrEq/izB
T+Ey+ZbdhODGScvBMnCNLoC2pmxyTxupE3oMKvizyUsNXezMJjWUcs9OXJN1ojo51ai07yOYX7bn
o0Mqr/vfLKxgal8hEQ2GKNacZfc9ZE43KED75J3/rdlWUBtvi7x8nCmH236bkyIn4yUYPxz0ViEK
Z/yF23063WGiwtyo9Iio69e865WsbQDRniDi7jlN4XxofeCUMeQbwjIXpS98eLH8IuBPX3Y/ZjOI
Ia72TSBp5li0A9UkOFCL3ZWCRDqOjoJwBPigrdzuezGHdCv4GYRiI6BMG4Q9/I9/XJu7UKmGWcY5
bQewhbY5ma1RdaE9stRrIFBLTkEaN47KiiXUKEg6LaNKPBasgohyhQ6bDXxr656eit7O0N5SfBnT
FzGf1o8cxPy/e6CNxe9MrXnvU6OIXeN31H3iKas4edPEIEWjj9XivnKR4sCqYF4jSNlVgxW9A/b9
wu+hGxWsmXcmLvL47NTLmdwsy0mMxKdyOlaaNHQ6AwrB8zkBULHxVjmtuXnHiXhl8C9xj6uMzrgP
O4mzAafXkLPEaQVCYgLzv9xSIW03KZR2rKfIcHneEDfMDPD1NSkYy3KVs3X98ezmXSrEA6Gk7T0g
9zVB7kK+65T4vo/Qj79uGGlzzFAFGa8r0r6Ne+0p4C+qJ6y8xv+jw2L+W7e1ColcxQpGRNO1NYJZ
zqw640KPHi7mRNVwJEqLOziLN770XxQsmbXUtZSkEapqW/qhf2Yc2jEj2MabCPpfb0UwhCExL7HI
njeppnlUqJDEXOHH4oNjJAr/uHYkdCF35XdXGNbJT75ir+gPxXehfdSQ7KQGe1BmGH0XkrkqD/3v
3Ua1845wxWPEMcTpxjVs/OZDrALUz27UDnzn+gYCUS3JQoIF28KjbeI7mUyOJ9Wzw0bGVFvUAGcB
6HNSvs/apYR+jFuCzMFaFY0Q4+SJLZKFHTCnptrDTE2OVK3UftIkfb8gglW/J8sLw1hds5dHVjiw
TiIzjSyBoY4Ouqk85V8hhtbh/gcP/hgMXTlgkFGzueaCrIcWmcv9lX6QQXwiAk4Cbj49Q+XwKSEf
4ss/rsT7jKsNADLd/gRZ/h8aGoViKfHaww/9bAXlSdfKQvT5gPEuYtXI8TfsJfgjITqY/NCp/azC
bNsWJUD6bNYnv3uqj1+YnZx6lqcbxp8p+Qc7K9ZakRQ5y7R3jBCDweXPvp3vW/T9U9muijiQsp2g
B8rvLgDKiYp1TvPtMWJH2SOhiaxN6NqZDaFYAzVwB4vzbB553h5QemhyqWoPdFdQ+TyXjXjK+C/8
ccjjGTnroAjhuxJ04u7mLWZ6fdkYxwP0UBxr4r0Ig5T1pMeWAyFupoERvDTtO3SANdue3smcgysi
ntmnDCo3lJbvUhMjONl0YZi+sAP5xv/rYyD3qvvyT0hZsC19pCnBqMnGPMh9Lk9n3Dge0J8prlxr
i3HfP0RMTPB4uE92C+IGrxBgobk+aWMLfRhqqzb32EOf2xbcxdxiE91S4P+o65nR7K7gA3C4wGKc
n2C8JgcSPQ3dNnWsbYMdtBVU688fG68pVHDlTnrHBKETWD5xeEntplhPnkDaAWmi6d4zZV6KtXIe
O08vIhyksZnudbk9D5JczjhEs1KmfAT6ugLiegGbNpxDGFkLwlp3aKwRdrlma9OxrAFqjOz7whIe
wMO7N6wgbeen1EuOYo1whhSajJw7H4s9I3HqFhbkakz3d2gl2nY+61LJEWu3b98bH/oUbKWvZI4H
cGYT5NfilL7C59pEa89eBOn0ZA3whEvdI6V4jJK377coj0TT8J/2WaQKXtmTRsDDEE3vvlyDAIvK
wapUNXwpnfcDQ3LD3O9qWpM7oODAWpBYcRsYb2gFCyJPBst10ty8S36ejdZK0FoRpIpfPAv135YK
ESvyGGs1/FQhmNI15rrVzT2M1kdMh7zUiW4k+K0J5aUphG8bHN0OX9fUcohzTS00BzaA9q3vhcDb
N9RXnEDfzprOwrOXq0No0/qiYaQEIlUvtJvxGMAIpGlLXgmh2G82VkQ24msFqQqQ4oIOt3MH8NOv
TZw3JUEnfo3It/Z/ENXzAsRwy81BpmNLaX/QG3qdV+pPcLfgMTAqAHnf3/hglWYPqD0323W+crRP
v3kn6N/OvM9GWMZS83BjLZH/vC//GOw9MMzuU/Qkm4Nprw99wn+iv8SNcnpYeHlwFTJbajsFdvau
nM7j/0LspuN7+SRh8q7H+YaVAG/KUNkM6wmYjUEN/+QQrpwbFR3XYlK/71UFZwzR9QIdGuZ+ycQ9
y+xlla3k8ETBFXl8lRlfEetdnx9MYKE4fyrZOs1c4qp0MhADLgwQwAht8qSdyIAQHcylobq5uII1
DwimJbxzJYNI08h+U2DFNcdm4oEuYxRe1Z5oeO+ZwfdbY0vlGEPhpFB0/Tdh72uv83wBN6sLU/4T
X0xXX1D6A8tQwA81lqabCRlO2qRt/HvTYm1GaSai2OnEwxba1/ZIW20n0NgVr3ouySMTX8GIq7oC
bjtWB9KxyDi/yKhcI7uhaddWhKN/pOJkD3+JXUJ86WA2WOssQ0frXNRmgEkGJaCiIRU2ogVoZNu7
UNjm2TLUyMl2mTIQVEMU1EDYTkyDuMabbVe8+yzkRAcr58iRxCKZBXh0QBR1kLl8QnQezM/axfO8
sFTbZqhFele+jYLdGHC8O/dI5fYwV2Drla0Zamz6ZmqTWwnqVUIX+UBaPG+Fovl0YkAW3w50vEq3
FS7FMNhJrnw2mfcEJ+S3+5/1jipDTdW+GZEBuWTcbQmSiUYDvs5X3XLwnwFOC4isLe62sMDhGw9E
73tfi+PgHTyMe3MDI8Yez/w4TrA75PvncHzDrbLEno2Omndcm5vynXxrnUG8eG3smc6P/VCztLC+
PFF6zshNL33p43hTRRbliSDGTtgWVi8YWUOCbMUryut+JDS/jsOT76vcWfD3vsY44T8ynKcg6jX1
W7NDkPNFlkoXgCBjgnBlykWynz9iUCiDlRp+86JPWpe7HGGmM8qsoki1RRqKCMOcnQz+a8cZJeb2
4jm+zzf9cw/4CpNrEBTr0XBDhVZozIEZMI3thPkY7ZMV8+9o7oi1ZUrsHiuDXJ2OgDXHwdpjxvGt
/bObQjFZHq53qPtRqvGUz/RT8PnTuoeFG+ag4kHPph7AVMIUBdYZVuMV19LkrgZ4FApZp00PQy2H
7d2qQgncMKejdlZAyFPC0GQURvaXOoYkN2mep7O38qxMQFx0jM9uluttL97yz+whQT3tM00mVPPA
3FqdTWNcVDvpZ8PVBH1jj4eyYJoDMkF8zz/OI0/adt7PCcIfnV3/XetC18Ao5K/IdM1N6SFh5pSJ
6OlpEP4nVpPaMmSUwRp64LWsQEYqS+F5wMFWFF3QFZQMvMsrwVpn+Y+fi0pDv5vlTjXDwU5TtecH
MhSnSsXEp/emRkvBWVT3Bo+8ySu7OCbsnV7opI50Umn4MTWOjqvIXJ0ANchbjbA3Y0pfG5E+4fOJ
wH5A5FXqqHl/xyLnWJBoNUMAZCNvizukA9nMSVnEmuDhSPVpUC1yN8O5qIqyETU5/KVx9FO66u2j
GiL76J7Eqk+FsGKwA2NT0y5IbCg60OzR2I0bIBsjF7EsmeKOaXY+vzirevKEoHZu7oaTjjyxkYx1
4xZmR0PRVl4yyoXeF0C5mx13KO0UM8eY3Vuwue5jqPiF9tNg5NoH3DAZLgizuKI8lYEJ0ghcsgPm
wDAk18QCZds8OQy1i6RWZzfr7XKmdMZ8HsuiNSJiRoMDiThpeTUyua8Eh6ewhmAXnfc5us2r6E+5
sPfyd8pSH3gl+UHPmk9o0iiup3AWYunu2DXFuhQeYsUp5LC/gTWWlNouVWwhPzbVrHNrORuIa1Kf
C8lKYzvhhQlwaJ2K3+g3XLqYSitWT6A8CsyiCsp4NP+Eeig7dQcifqDdS8Zur5zSMyMfU9V/pf62
bOcRe8g2dXw+ctW4Y8c3ypW/lSpeejTSPHHhrIteCG4E+4Oe8u6F1cONYPO/m9GwOGdUNtGCw6i5
2LaE71xI//+y3xKIZGn7STuN+mn3mXkPjyORCpcDxeUnq5+SQiGIJhymdqR2NqIpjs96R0LJx54P
UbNWuhazIzhS3UjFpNzrzgd9Yj4GZDfYcdEVNjBcg247zniJ8fJTHLWy7NrOTz1BcIgcE6VXfJjZ
nnUy9rLrIBsCoWTssJuXQNLXHadSHT4ldxQf2yYaolXrGURbUil4JX1iB/Mj7mBRrnvzay6+ydZb
+VZDh0D3MrrbpPu5ubqpMira3ZQRmvjPPsaRLok4CSHMDknjE0lGpiqF+pPFymKtaFkN+gKcx22a
PRMeUujrT7RPIoKEqxvyFDFxDsH9VruvXQbgBKDdIHE1tAatjyTRtqWMHZygR06bqF5Btb8l6dNY
VYnZG/1uWPq+GsncFLr778IPOqisZ5iyjPfyO9+9UR4aAGAsGD3jpz0FPyAg/jZQmBW3ghRrrx80
1Wk7mYpjkehovY61rOqfmNpkEQNm9cQh2wQXONmFdchjP9+CWIXICWjmo5GyvD8YdztDyrgBqzJh
FLFBV3yEzD4ja2/CTf/1pkh/yFjzjQFoLlhbCRj4VrdDex4ijuzGjrAWYkYXSVs5V1SVOqswSH8S
dx1iTfq1Xx+yygumwj/nPo6yfac+F8vOoasjPVfPwXOHI7D/r39Z7j9FXrjQi5/edYKziMme8lB0
rFlMCk+Vp+8aAlttIng8EXp4wB/Adn3V7VGINUaWWCPImRtfDvwHZqwbLWC7tqh9EfWPm2z/63i5
TIkoE7ToxnB3WNlL7fQusjWBHPNLnzJ7uk25YjfXSEqM4pha3qLN1mdqyGvBwmXOsdMYOujpSfWN
XqezptMQthTzcqguSQ7BX/7KHHHDhcSQLxxK4roapBeXEUb4hMvPhKAKYCrveXIkKoX0z4UtyPs/
sjFclZyOQrekivyUPORY8WwrkkvgfdSWCMuFV6Tilrh7OG8GYRD48tcs2xb1mWndnDqngnRwkF+e
4p1XTmtBa+5rSrSsknUjcp9AXnnULDyJfFO2xXbqvM5ABGWg/rHyxG/PIGvFZlC8U/Di6UDSt9pc
16MMfGU8WQ4XfVIC83DR7lamcxOAG3MDsdiEtfhSqEpDt57gAkV3PPEB0+azWEZerH2aOtJA9/4y
c0wi6rH0Tf5LNf4arovmEFKj5uTRY4MqV1LO/LKZETTGC1BZdRfIwh7FWaB0xwwlX2ydTgvchEk4
L3OT55OnMq0IOFLTPW+UREldMPbBGeabatZ6QnyS+/43jebPS+YEF0v7BkV4UFJx5/zZvTWuIatN
zTxqo3eqlGs78GqldOM819KbkTe0j/Ld5Rhj2GNeD/IUcpeV8Nq0OIkFVCjPzWC2anQhBSUYr6VK
t3zCcbGC5gcus64jDIATsfFG/IW9IaEszQUMaRDnDG2BTAUG+CQxbykOPztWirPGa2C5832Jrp2v
BHibTMl+ulCaJOuLgR6/pIg8o/qOcByY9x7OVxi4EfJsXE8UOlpUkRlwOCnkEdlFBLi9TUhEzyI6
nraEIMIogud8TtHM+O7UH7+WgEsG7fj6CgLWbBUMcMEHNds2l1Rb/hOfyVvCIDQ20Fowyaxj68tC
whqajTdZc8wkI27mJv7b0ebsyh9ZYlv1T5FuJk2ZlNqa4rhJ1/IsjLr9fCHy56tQhdQPBMGEdIjL
jQFo8h+CTrT8h9EJUSDSWuQXfy4RBSOIGvtTC1jBQiE8jQ71LuAr/vuw+t9dJVYSMsygBnHwkFjL
15nx6l6gDYA6aE59F/6Cv6/Mm5g/EAJEXuFcQ473KNpYlxsMBuymYaKIfDV0GRhZlTZkKkRMyjhy
AzmAmtHHMb3eU8HawuKHht/07XyYd8ATasktd0nF2ms0nx+zqK9MY+G6YYson0KclQoIYV/xFU1o
Vn9ELqAzrAs8DPH6TU6hoGDCQFclvzZ/ly9rckwotk9Xm012x7UjKpSgKgi1vfM75tlJw7QHZh7h
LeN6BW3q7ThWL9rv5mXzOBWPVMJZXcIbe6Xznu+4tWXFXOJt92eLVE5moHWkG169BZz3GLYtEaXH
fvgJvr1jN8CReiLJr6VaJXry9oBG0+o4r65u+Rnw0ygnD6xDB3JnKorBihbZ6NL9wtSj9FIHwzlx
aAU2yJaVEB27j9C7DzLgvzMQqP4AX2RVT/2ez/blmI0bBKANWaAXobj4hWhN3Un7wBxRjHkJ64Ry
PfIYh1jwOGeFp9Tc6nND13tKnb0cWMrbWDbYbKqa88utFjjvVqKF6B0g50zCVbdIE/XiV72cq8fo
4uL045K1EMxYXyLHvtGLfZAEW2GH15DeKOrQkc7MSOx/iZQofMj9mpW3+6/DMJelwBQ6DjBXqgQt
5FfKU+3lMvZJeGiVO33raIIT6BZRthSC+fumT019lhb+s9kGoikGQWn0197r68dFB6CEpkC+Udti
Sx6GxnwOmzNKcFx919GKP2kniJ4kq8aH4P26m7lGzsg8/RpELrmY7NZmSiGaJYCIVmI156T7DYye
zL0We+epBAKL/TaKJrjShRu4UOesvXaNhrxs0w93laI19XE9UpN8ddq4HCmhGHd6kQ0ztWvNoSqY
BF3s1g02j5eu4DkiW3cwxZM8fbsRfFSkcVL6dJIduzH2w/7iM5HEHkvFP9+smNJPjn8tmB3MJAy/
z5v/KXtskUvjTmeZLMcrpU4Ghz/+gdAW4ztZza5G+7kZHHNDh88W0DvqebtwwaIrvlptxNRuavvg
Xz1ukeASnkSIsSnoHnJcODsYRh3t4U91vVwvRuH32r9xTBrZPCInC5HLE8TAfb/6CIDbweSVktfh
lik9PMpLUG4S2jTJxZj22CM+eU6AZAufzlhwqiMTowh/7bipONnNcHku3YRVqOYs1vyhP12MDr5N
HjPu2Rk4/Tn+o3voWn607pJhBJjVkmgsyyaIVPwHDZHzcHiSkXrmJobpR52fJbwJ/iXTMaPH/KfO
GXJok70Or+Wguf6fLuueSz7nG1fTm4l0w1D4AyPNCYPEHGKI61ps1hK6PJLx6wRyWjm0BWHlPhgM
N5zY0o4pp6eLaTwacTruJvpnx/9/S3wF27CY1/+fj9mbVDwU3wDPvZ2XXkuPibMt26zwv1VMR6Fe
RPdwTasOlbHeVg0UJFdZiOsy0gzUVnhCdo+7slY+RzLEvWi3VsFXRTA5Tc6xj3tvVXHBqC/sQtx4
0EQHFx+C9J7mlm+aHcFmPWbwKGdLpF77w7r2eXvi9TK15zs4rcYfFo7ns7tFjWqK1dcsrIB2c1mh
UjG9L+c/E0bqp0w/XW3H3YTD9K1FeGrAgx4iP1B7P+4bdV/9paqTIsxlUOLtlQ04mfSNAaRbeWE/
AOWAwCRpqemUcBP5NzKWcz9eqQMk8HZ5wmXdEhX9VCVGRHNYGwJjL8bFVpvVrP/614rfKQIkFN6C
6OxOoxpS6f0Sf4WKDgqwJitjKMQHu0QfdIdUs3piPyXMrR5buxxVDPXbbyDHAPfy4BknJO7R3Iog
s/SvVTnOgTUpPExXEfrabUFTzISp1MldvmeCT5I3vUxFwXP4QFEwiw71eSOq89Iz7kGPOkSsNvbO
IGyOsOyZjUQ1Uln233TQJE96vwVpAf/q0wYBeDrsyB6InKjgpceUhgKTnv7R7ax1iOY4ycunapam
GWUxuaZk4klI3Cj9R2TB/yCu4G8EKbl4Vvm9Ie2T3iqRjFL11f8PmA0zr8pfQvnfV1cfjKSVpL5E
kcl8DsYwugxgqQ1i8VJOJZff4Uk3oTpMSfjCsCLHPiOGQE7sHK5rEcqWX3EGvLuq0Xg16h1eAdwp
tb3Vxp6XqgZA4cXInhrCU8Bd13zJoldn8dDVO/zMUKTU+G+tgbPk1qWmHR2aCR1CDTb+Z2/s/xxd
VncaPLJCpE7iOvOx8gUN6n4h3WaD0rTfxTQUaV3kHq8vHOwr4zLMa/IPPDY6Pp6CbB3nZLJs74WM
d2fTszwZlFYekowPFQ0/7HeCbx1XBaO+V9XuT33FyxTvK+Ua6hiBqy2Cr5H6Pb7T+cw0U1jxYW4Z
WVOTjJZvZLFWDkEaS647uHI6FtwOkpIfL4G+1eETN8mmpUNlyicJJdlnA2x9C+7wa/hryZ9egthg
xYmG+kRy0eXbNmmAS1b8Vb0F7VucpPlD1AfESCILmntGWc+egbnUh5rTv/kO9mxaOTfvLyNQV/U3
KgLVia9RlZJSUdqm0g1X19U9BsU8eckFG93HKvWmBQIOHvqL5JuEsxPY9t2O6yRz7Fxyvv324k1C
y4bxCJPzk0wCyUmFPNKxdUGfKrIXh7WKDQ2dZaYLnIXKiiTRldKYUtjLxicIHJDTEP7zo3PVsPTL
BYLFA8ZURxoiLZ0qwsnjH98SezrzuFvrVPODBl6bClJouTyPYKY1zX+7q2aSABXxfWa6W3d0bij/
Jl7e6XOl1AVpMtfflUeWgkH/gZVpJOpHDYgJmMekpbiBhj5PREtlmkPoTJA3GGzV6sbMSnxrUlZL
SDYCd1qJkzb2NQ9LmFCJvmMkzQciiNxuGAFXYl2YL3NVpIybBdnrZVNDxKksUQiwE37lH/aKDsPF
Bfy87v9Vw1XKbZTyGUfkbGcZFOVLDyB72hd0iOEImzJV994f03ppXHCbjBl43ZefjPg7427h5hle
EIhQpr6ZFZVEBf07NK+l3CfE8XmUTDjZnMkDFGWJXsgSkKXU3i/mDv4JD9CdpgM1hzzQUQvVLMaK
AuLWUyikXojqAHkQNUVtxZtjlRjFRRV5OzzsHfwd/CUiKOgFvoMTCVWANkDuibAlLB5CLYapnK9Y
mB1s88ij+WTRfn8Kx0wdWfgK2dlsxdCTwhW2at4+snpIz2CqT5uuGSjxO3ciZPb1E7aFLUW7Z6ZU
IZBx4USV5kDU6cBYVEAuLGZb/ICHKd+6KYOFEjWMzhzehfOs/IHzmMjrrrpKftPaLGqmNaSCZZbx
0Fawzzl1B2JJqvWDWLWen1FLF0QI2bqM7wj+qzw8w+n6JSsaUuhNk/vpqqmAqAw6p+tuGI0LWPdV
Fyj5b0AkPDOOyBiPGXapUJW1FxP95aPCoC0L7nh58/UNz/tg+H55ygb8yQrlyHXDEjzOk/WHsO18
HwLbojKv0DJFRp6ONZ1EEwCBDLbJWIEVDLnRBzxM8i5+9J38YS5fOVCobZxqjFddGvYiTyngHeHw
G3x1ALbifYi7bhKxlfB+lZhI5wW9hkMopdgz7/26nijjVDqJizqnOxeWVGUL7kbJUuIySGe//FvO
ZXteIbzuzh7Zp8s/gyiua0OiZGeNBr4mML2uu4hjk3DgOIUvOt0AXEv7GlvOz6mJYw03pLzkodrJ
5aiDP6kGZIK6i9V2ujjUazGs397MsgBi+Px07Qn+1WTGdIsUQp4U3mKeUYdtFPvwNNhdeyCU5NN3
lIw57/hx7GQ1lNjTC0ALJShw7rMSSrop6cGOWCG8Jg4KKuoH/iM81zRuXMSQvkjWrwmpwU9fcCXP
coaBFTknySw966ZE6pI+oUvPleOuHEXJcnaK9kXZaZgWhw+tEHIZ2i32z7RrPkZ2RtZKTGVwxek5
mUpfKD7k1bi55C+z8ShsVYbRZesdY1HysC4DgHgbdfMJFL85T3/nxGUdxqGg3QIVmOREVyDXnajr
DwujDiBtSqaVDBwvOxMdLjyhe4X1e/7KEm7m62izoxqCPL1rAJiYu5RnuCLvYPRStZKKRAxbrwH0
Kl1EARq31WGRNSB2htihznRy+4jmA9+x6bzEDz36OrFzGuW8nrUym6RD394eKtHbvO/dVntaveVx
3ARHNFhTXFD5RHplyg48rF4k6SrLzmNmyFvJ4HvpD4n5MUZYjfBP19RmI30xkOTCzAaSFPqmY3l0
lUXz+4CM2Hi4ujyBgPZzGGLCRlM+8x4/PAAmmy+jmvdYtrc8PtkSrYES5c0eJAlqz9pFfDKAOsFm
FhumLJpvxBk66MN+vJvTK/LTV4zhkrSdrnki1K1VtrZXYdEPMfMzCqUm9YkZH/2Y6EjoeplV8YNW
rm3C6vtCmGBhIytsRWYWeGtQPmsiaFC2OwNcPqsna8FeE9glfIbuiMhpFTB5FM0KLGmRPGdf3HvQ
b+ntzjwkw/7+LZTXrUjtjL9FJZS+VU9lJY4yQT8DcvZrHMc9Lz7Vw5D6xCM7Sfy+7PW/tcmPJOQx
N7MltMVtS2WvDp7X5P/fZXzKJ3Kos+g/yr8oXcP66B3hHgLXlvd8Gt6/n6BLM3oNe4dvdm+adVnz
AKLqHGFdZsRVrzVaFcsZZwGqVxNTCef719uHK/yFsLIz69RidjcqpD81kR13oKdQSAOWq926z/qv
kk2UituY+8/UihuVT2S7773kCFwrUzcweormdvBHjQi7e2jHxBq73Z/EkgpqGrCzayDawxe76/OH
ky5YFcOG3jYoMvE5k4FFMo/aevKgJ/UDFCKmHoMMJLioJI7KrvnyJc0J7fRs7B/LirdOzGqp8KaC
0g/xoFh8tJZKxq4rkUrqlSrq7Ogr/BS3a6vV/hi8lsEIE93TMiRV07x0ba2xrbo0EGWt6FJkG8Q0
3No5xJlzEVPUm2Ra3TegjTTDceA/EJk8ZhmgOAXy/G4K/6h7Chr418PShSbR5p2NcgP9dp881dCz
syrLBwhU52/qXJmnyRwkOdICo/yViG/zpFIo18EqLB3jVAG57XH9dX8XJe3d+y8I0T8AHW9X+VTG
7A9T1gD4V+RN8YFYY0gqd9W3kAiFSMj8RJy20JwhF3afY1PFy//2/154ob7k4eTcf+d4vv2l95zL
NO8TlX/1rCV/M01q88tvEvhOeqiYTgGREFWCurohYCKISy0uCn06Fv9UvQYhbT0iLZ9eBiCxzGf6
cRZdqH8GVjEEqDcBtqccPqjsZUrsyFuQGGQXl4ETxljRRmXjpOZpvQEnkDEYx0vwQM+lJ1KMViSG
qgW/wukhpGwKeLXk4l5jenNyA5lY4KwOI3UpSEiNFKtO9BddVKbCgbLQg2P5m67Sy8qgaOiykBxU
XJlHVWHz67Ohjwjc0p/ALc04huc/T2vIl8CimIzd0Um/JmKCRGhbXxkUFrFv+EaM/QVePICLgOrm
XZR6UxeQeynJpqySqbHokafLNmCE+55WOXfzAM+vG8oF/bHMS7Av9RESAgzV6RLGnZjA1WrCrT0l
oYVWm5jg2sFKM06G545EnZoRiA3Z+2P6cOrg2uRXkNRCooXeob+6ebeK57HPGwNRnQeHZVep6Gck
+bLxZDmCeYOPh5O4tN+TiZFBeZNObYya4zDa/L6RM0+L6/V9W9Jrrwgs5MrbLCTW0GyKnSNZV886
beT4kKioFQfHKMS+hgX0h+IZnH7+OZ7QAAqJ0o2E+zOJ0SW1nz8lF0n8VNV+8vqgXMeBJ+qSyUD8
HK7OtI6KgT3kUxCjm1CbNbe3SpN2M5WO9sc70gLC58nk/jctxv8Fzor4nBiBUEW+a7gzYZp//Fxe
CN/yFjtliZxl4W9EOIE7bTe0Q8AAcf2lvq2QzqfOAqH8wQxHXqMO/6xANco2jtqvsKs4Xabb0Ahq
H+BVZuiNej/hZrRppxw7HrrZ9f1VZZj2nzljrOOFZJC4zPZK4L2GMRSn/SrwnHF3cjE2oXeHJpHf
SaWD6UjPDZMiclF/cxMTHd/T7zJxLlBYdnFQqzf2MWtCCd6UHaJMcvZIlPQa/UGsrQynztq6lbUY
Zkg2Vuxo562LyKuKAV/aHoyyI32lCN8SB3JlvFhD/tczhFSYBgPWyyOudQvO3YfFl/AwEKOSkXFm
b69UtIVHErcxd/RkBLA2wWfKfMTuyLzJGwpMPMP8eael9mLx9iQhtz7DevAhKzbx/tiBXpCLeKbc
s6hzPpf+8e9R8xWkuLoiOuK0ZIwlEDTHJAGRBwyMlaooLOYPQuX7dROkeALFQCPZJXjk4YNscsHM
2gZzu29/wyvZ++JX+qQrqzWdrL19UhkrWO4KWCtPNIYrXP/ysFzujP9XvPoeEpr0uG9YFqZ4jByc
zrsqwnCvAxDdxIBXDMC7r2Hv0pA+LUKF86r6p3lN6VGoGun1TDak4yzmeIZ8zSnZp4q/3lfrVR5M
fk/puEX3CmXUWjrKsnv54Ww4mU3HpdjLrda67GevmbOwuQuLcXvhItPBgJpVoCrrYdYO7KfiGudD
6oOxQ4bsFLQX5sRg54kZBVX8vfqN3qpTz4yrdTS8qeWnLuZlGSHPeC/WjPVwwRY5mS7OJzQSkrL9
uF1XUA1RfSb/dQCicd1Ec6Y9DWaLc1YfTR6smBTwIrBlZra/+E4GRlb7KOxFjadb+rybl+3TCcQQ
K70YjT5YYFPIanHqLDy2YkprHMc8czCRIbHnYCH8igmyvGEDKStfeXWwEqOVH+TtiZMDUEyLR4cK
x++o0GeFJj7hQ5kkFlMIxJW7VJtHhARdcyVZVYYfjy7IsEk+Libkb3nBWYdg9lsUDC3+aN/7ssJF
NLUYo96Jd1ARPU+eGV3tV1EDNHQgLyjo5kNsSYfYRybdvdiTEkc2A6ktMlWRWSxC4RQUlnPZqpv1
uQOqKOvcBqAeOr7YMG5BEe+68ENqVOesouBBPn1F0sgEePtLQKekPdEPfnlA2USYq2qepH9aKxjQ
41E2PsmlmfZ9vVU9q4kTcAUlDNXNY9+HRhQkSCKlK0zYmoiwuOdqSG5nv0xjQh1Ps84Imyp4rZ55
Gih8rYAmqMNE9PMGn9vX51xY0THDxNy9xdWtHiMFKB4JrSrvgRIOeR8Mh63Z0u6Ok5l3LvxQLnxf
p0MbJRbgeOtqC2uYxph/MTiPc3gC7W5uwzpbjgSFZHFCQAw3/LTyYpTqlyQMzeGkncuHaOItgQqs
qvuzsPsB9sRQnZMm23P8SGXvbb1Gkk7r8LDBguiLsOitJU6YpgpaY1qZBoDMeiehrKGBeETZHnMg
EsqEnEXCC7ook0JNJORgAJKIwvYrtgNXxfftV5BvNiKqZrl/NHB1qdnaYfxROz1Y67o5qxRLmLzA
KYDtqY145iQsHY1iC6WTDG8BiNZQ10nOdRaHkRX3YnNDXXP/uB24fZAz9Px0odf18fnq8IQXpzaY
zjp26EYlFOqH6nu2BDJ6cx53FQm2uJ6CzRMgR1xiXJIWGvmBOoiXcsmkKMA8g6cEh5Z7A2KoqbpV
mhYLkQXtqKV2zcFY2mUQwmhF5ZzB7YYiGIeGMc94xin6AZigMBfxI6V+lRQEWDZGkeTnlPu4kajA
fNKcJQvmZ3Ylf1Hn7BUdp/I3TZjLXLJyBF1fOYR2m7Iv17tig4qW6Zy2Nq0vxgMszu00EgiAVLwY
pnfSuOmwlBPFoCP+MXLGTt8jUM3fF7K5IDKGQN5gIbMMzJ2MWn6RSwt/WgnJyLJTk1lQA1SVWfXl
ssU7d5fHWUDxrz7AYbzNhDQ5PYG5yBxe/ZxNa+st+0hZ55TeA0z7BKuAXtx/9ypks4PuyzXmxILz
nis0JFEnsUOoYIJC9io/Hq7tSPk6ldT3pU3gaBVx/0eIxZRmMAlgKcZi1xk66D6ZkZwaMcUlOBVz
kjHXYgvM9j4MbF/zCEteu9z9ocDVlZh4RdkA+siPI+TgFEB7V0W5HUTMKfq91yRF1xC+AzmXbTZS
lLj4TTrRn6u2Tt8gzsIUAA/LgOK48fN1awWfi6Q6IQShBLPUIzjBy+Do8pqQHPcTESjiaSwu32NM
3krxlD4JbCShFTtbLihtUGfHx0gaQfBvXiovQfOGR9tkdzZkLWFJ8CP04P2utBLKibcrjHl5+ztr
5IKqwntP00GzEtph3l9SUjySpm/KIU1qWs/7I/f4DwPzxa/woJcsGo3ies0YT7idt2KzNaDM6IT+
xDQgEuut8HaGa6uYasHfhO2aXbOVAyKeAgx4JMm+uvGuIDLS0Fqk0Ai+eHdtBNQyfm1E98bc2KV5
nixlWZPjU5X/vnGH9SiZgmmGLYrXivm0OhH1Juy+OcDF/u17kz6b1XrofTnWjZfc24O0pErXcEsl
n7EWo/7DGmB6x0vrrxYcFlEJQarJ0OAGopc006+M+cKkKJ/8OalvZHGPF5c/c1IAPi5/XeUbiqJX
4gfLwEau7whBZP1qHsFyWryHJIX7RJTqI3xsr6MR5ZHhucIp3HtIpPOvxtbf5YtNBdsyHSIc/F3z
ZkNBR5QSbZX5Fvm33JcWXHFLVDs1G0r68wQiim5ErICko+7kTNv2148Sq/66562OjZdxNmMyb5ZO
Hmq3GL44ELq/jIziQgSMUDzeRrDpnymptjTqzwjvFtD7gMK+X5rPQmp+o9eknyz+31+4rQCN6aDy
SXpj7hInzF3khmm+t55hl8csQR4wTnW4YICiUUMnm6etn4nxqDDVidfomafQRLRKK1g44ltGfW6i
5RcGfq5h5+K+fAUJvytLhQoj4s623eB/AoLYChT2jOipynjNYAOJXum4s9UN4CFcFjhMUMd0s2y7
WzwKPfVoiysWaetnI1qrPqbgQyj0SpouK8BVOtds8Wy7zg+iWoJKm9yJzAtEP8mQGUmaEopneuOa
uq+r5449Yyq1ULppFG74HUYI8zDxheFbXCUt4oS5azDSaVTIUAmFFCh6e8SBxJn86n7ztQVT1xKD
mPYZyOWV9aFn/KGLIRMPDGDp/2WLCuVBD+vN3JIhROfDCmfzcdFozMioabmUVMl4FLQlyzjCpbc5
wgVVJNEjO3IC1jtWYsvLFS0HC5QCuIoJYekDkOazRcWp2X96GtwLpc9OQB1qaXztEhyGaV0VaOzz
ArnBbs3FjAP71RZFrgn3i/6brcQ9+YpGp2pLcoAOqJQMSmcSgXyr9rixVZWhHWtaH964y493n/O1
tXKtrwdfQQu5mVzh6LH7t09UVOC1WwWGw8eLtZ8ecfdfZhmmFjqDVxTXhLYZRz2wiNvb3I6NrQHn
G/IkjIe2Z4xSjUbBSuwWHJuvGkwbt0sdzEOkcb5yiW2weZZyxvTJqQ5yHOWowcEdO/Q+HEuK9f/x
hE1zD4RehfrnjwWOx00Ev36UQtxZ668Na/UcR2pEg5a9pKpsYL2w6ry+q2N3maSqvw0eFvGEkgaU
pBZ0GnI8z52mExZo1wQa6vZYdMnQ8N33D1LvckYeXya2TiJH/+zT04gB5xfvAEtftH9+Uq6CqDvJ
uSmajgveYyutmsC7TggxhwI9CWvi06Ffbaf+GOWiPA+mk7QBK17p40BxMvOAWFP+v+GOKsvA3Ifz
fV+m35nqw6ixBeNo/XzH7TD9PgmlCIdlYP0YGnuuBBP4U0QBVLHR7wR0fRsXP0CoFL1LMpaAhVAd
NSQr/4rCRAIrf3JREKLxQPgKoKQky5F0WaObpW6afWs8lq/fiTx2Ds2NFgPm54jmsvIai/oqVl4u
V7mx95NO20+8YZTtomoo2qzN8XFk8SkPBIvaKyRlcnqseLjEf2TyYgv2qX7FJhOHflX58s8VZpUj
7KFS/TYD0ZjtjV5aI4ZXLTwhuZq5AUXRZCsEY/8OAHcXKYweON1q9TtzoB4Q2fLS6O+iVK8r3zt8
dMhG8nPArAC+Auk09UMNZP/PxbuX1LurC7jU4vn7lHSZDqx7+iGYKh4bx7jbCpeXzbRti5VzVUOf
xHDJ4g2lex/IXXBrwNZlgtx3fQbOz6gzqjEdYU5pV+L7PTDltzmaF0ii3AsHdOTzARPu1+d5ou4B
Owl2crINqYTGOqjuJtLqXn+BUvhUWuSaX+8mZPEfI6EKJq2qQMNVoWKNWBcrj4VXEiPVAwuJjA4F
WoWVj0WNMDgTHLEj69u8y8l5G69e+WRf8jO60rHYJqo4BXMbDGRnGHyCfvm0U8SHZ09nKKX7FY0Y
VJRC6qzHNFyuVMScRXkCPulhhbvidBN0poyIYB51tHfAfYtg8htYc1HCvCgRX0Lzt6OZSZSSHlvV
MhWwkahshiGAgapVkOB/h6xcuf+azVwuHNyc1QTrYw3EdyTwhVrGeKm6P3ZPfhSUb2bOX9POLFv3
j8Fg9vhAogF00PnNpW3P90j1P32nQ1KG9BDtgB2+hXCVI9SBG5ybItBigHrZxsKWOYYRXOsS6Yq+
6O96gzqUtccJWmROT9wsgkNLuajM1LNEAWg+JdI8VBHOyBLob2OBfr9igr2SiAACFK9IthPVeHsT
07t774PmMuID7cf56J8bXGfjPGaMzURj7OUMSUqGrAm81VkHLI/ZHPqcqEyOCHv61VMCdAByqWiL
7m0qSr1iP1qNBjboshBPi/NxSmUntUVPc0zKXxo/mS4kA6FSRAtb3pQR5JzqkugHCPDR5iPikX3V
PF9bv4b3PPaqPkZxG40odMxBz5nrJvMejS1tuResffyW2/1LhC0Dph6SKBzV9cCXyEzwceYRp0Zu
WAF+LReGa9M6oR5aq8chO9iglEkmd6Ncjb1IPqR4+MXvqM2whmAL+r06yeBTUciWejduYqvxf6A0
4kTfwG7oH4gF/nB7mvoi91xjNpBOqQNpvwNCXsDLRPLFFsas1zqLVtO827l74pZgATm+gA9PUmV0
xMv0S5gaoZbgRJr5MLVxx4K4h2m/KA58sA6NZar3gH6fFuQWo6P9iapc73Ah9VjL6qS5GskSA4/w
X20hn12DBn/7wbRBUuCiwwf8r137nkaGemruGqF+hLoj2oflQBZElcdJBw+rpuMDAezyJsasftkd
Sqb4h/wHO3n1Fk8ohNili1jI/j58WCi878GJAy3ayvMPrd4usFYF7f1oNTjG9U3d90iUSiq/qAcz
hj9opdZngWLcjcGf41iZOZAAmsa8qA6Wf5ll7dpB1Cp0s3jOxi5RBJ5+XgndgEAllsiwPUZlUY7n
bf3vgZCwjKv5wEreGjMrC3MfVb1gJXh/9udkrRa04hRDxmbwXmJSUmqQQekQso3rXn0V6zsgy26j
HlQuQ4Fkdep/0ls+tmYuHs371l0xhf9qpPW2zzISRoXX61K+sPy68bnqW4e2DihNfEXcOrIvnMl/
cwGye+hxiXc9gvNsnVBOJuoWjFaBo7x5+Kz7DInP3JTosFFsdo3ishk+9BXaUmR35rgE7N4dtuMI
WFINPRHuLBtvnCj02iy1jq++0koTeTPkfU5kOzD+dNWloP1bZyPwCCzs4OogGXqrdLcL30xJl/PX
+RbnUNL5T/2ydBWTy6uwjasaMHe6fS2sLw9ELqsdt3LjUAjEJNA7O/6LorfCWnHPBOTEHKZ+JgLt
kB4yvUXwG1d4z83B7HCslQt/ZsUFH5luSd5cPGdHh92ni9yRW0VfzGRcOXIJWLAg6BKn8IkisgrE
wpIxV0y3KiRuInzlumIkmQaQc3SsKsQDOlhCMS85EUjMLP4m1ArzO1+DB7cZxnMHEm2IS9/e6c9G
iBXxqjduiDKazW+XIWO4ABw1hU05Zm9s/0/vdfIU0QLzy4LuSPIGg23e3Zd49SShUUt6KGZ3lFwQ
AEyvqNKkSQbuoIB6GckapHbMxNBgI2V2ewddPq9ngdwRI3VUPaxxZdrQ0FJkYquvm05jalOzvoau
A+cbgr1wZMmfTNiha+Ota2A9n/ptgAniCWkkGKnk46XZpgAO8qeH8mLZYIUrOyNBwQUCxeux+UtN
hO4FhssdMPzsF0mJRV2avbfIbI3Qq8802UzMgDaoLrBlriblQtiWcUkaURPJKwY9G0BQqvkmkbDH
NtS5IRKjeCvwrYC6n6fBa8pVOCakVEG53+PTrwTZY2Eox2IiJe2+66mdqAXopR/TqSxFvbq2DIXP
qG66kYPod6ZjOX6Zt7db3iGgj/kqD/gr/UBDUbLuU3MFdXJJARv2GhZYwBKa42HrzJK9dke2Nxzf
KTz/fz1YDKhWKLybGa071MdLJpf9n3FPTUt0/IguqLGtj3N0VN5KV4QQjehgRRC1rRc+cljGT7jT
JER/LA7ejnnUo6ISl1P5kKxKFacA9WZOEA2FpwjDybIwi3Euo0WI5nsplyFIx5ywKayKxH49UqPL
bN46djt+kkSMBh+oIiQ6G0KF4hSI5byahMdZZ4C/OvAooUTfuZMJjnPX+vWcT7qRsiQrViHIDs1f
VGbG1TqVclXyy3fXRtzNRHDONQ0GkE7tcnmrNNhT5S4oAOLQqbsXbftXn6+MkvZpQHZvFb4wozEN
R0gudGgjzxCeLimBb7bqSymg+kY1aQyaiMBw3ry2VSw1Jau5bd+TpV6sLjJC8wzg5ccN1vAIudR9
CHMDrF4G16c3PJor4fNz506OxqQhP2EPf92JrxuWV2epW5pDFViS78yRrMX09bj8RAvATlnojj2S
ubY32FYI7cqJG1G9N2Yc9gwpi36qDIkqJ7w9XUDXe3fGXOkW52sPsRvg+HCFbLrdHXwuZatql2nL
kiX333MP7yBdGrHrualFO4JEeiaxvx29PJi5+RlF5k8JY7aEhtymUcj4Me1T9dbZxOo+84hNeE06
8ox7fO66XJiG0ZsU8Kk745dfPtX9m5gRnHlbk+lgCdtguvMvW/nhcUuEZh6BLL9SaeG8If+3P5WL
J3EBsBI69iCxQGQHz/rxuIg5zKZDXyoII72aEL1OUBYgm7Evr/tOZroW0y+LCtPXUSen1jApCFFO
0rYxlnXxa613Pnv474qV2+4VEsadDAKHvWIBnLmd8MUZLSQGebTR3coMcLTEFDAbdtDxOpw9+zyD
IRAu2Shf97hwPutRqaNRJT1y3N7W7gyUdHdrncB13Pv4y/gEBrGIC8vtDKHOv3ip1FdwbvEJ9oY5
dP0Kw4QlngDRHrlLniVWQWrfzRi7W9W42h0uCtrAoFK7/0nxXsYAAeR9B2BYdcT2RIHhQiiNj0x1
ij8PU0zI0K9sspVP2vU6qMpX7qWERCML8EUMn7U6BJdJtyIjRZmm14yygQJRkAY85Frun+HlH9Lv
uxxwPEUj/kHXYjOT7jJ2vHhFFibILAzvJzJLnGAUCPB+CLoRmTy+c3tMpTZJ8JUZkn+oyxjdUHg9
dih9RNa17eEl2CMkW6HQ/5R8o6C1olHG14jRHLnq2UA7ykWKwzBr0oVSQuWF+tJQS9oavEHn6Rs1
5p/iNhY5OHcg9+2GrC7ipjKqPyd+W2kM3Nsd3Ndrjck+q+52+OLq+T9HYUFPpzDqkIoICM0PSWHD
xsZOkLFtTOZJQDHLlEE9BVq7XmVLbjQn5dKu//RsB1yF5aOmSAP2YD633XSQIJq88pBmE1FhoFP1
4Ld97WdlKt+gmDm+p0PAxlmRx5aiBTLbF0yapNSDIf6zxohxeBgFG1zLMKojE2szAAQFVTA3WUpQ
66okxEeIWqsie5IjGdSPZe68Hl31vxAOjrglu6K8MudIpJ74uVyFIGzxt0ZSc8ClNB7K9/Ok+QS/
3Bsenw76y3K0EWosP2fP+sASTTWi3ohVGEbNEFeZigEOhbl7dnsTeUqi06i0MxE6xGMSmUKz8leK
2gRpD1W2CtAtVobkb40X6f9wJY8rTWSxmO16iXWQ5kyTUSe2FN31yGAnNzuSfpfAaBXtuDz1CZbB
CIKVnFPfY1jAP2sT3LMj/gINlROB38pSHpa6VdAUCLIXeNxF+0ObMhzhtZfdqQ/4F44rF96YQi4u
Rg1bgCQdrf6l6FNANy5WjM9hASaeIwOWhJ2qmSXnqnkgdd1MJZrSdD/VTnf+x5ShkW+gNTr6EbdO
4W8ZA6dAE5eUkxcjh0TAGP6LA11Rb7oNZpGlRcQgsnp/Lb2dr8hbERgr4K8rBPTKXBi1S6bYtBlE
Mqftdi7YQuhx+NFDLfauuLh9oVm38NAvBELTe8GA8Zqwf8HeqQWkLmnnvPKVfYnWcK0QpuRdOVcA
BZBGz642Z0U3W9K7gQWCHLspu3B15jbEfccRC5e/LinPPZ/4SrTVI0NZHQjmuR2OKsQeUADz571b
3Uc/veNY0HE60anPULyRsBbLd9ScZreH+jvA0i86KwEijho7PlWp8k7bBmqhczhmSVPefGJoMrSQ
jycl9sqcPtdHt9ykpjS2AZPzp76Y8aqYg2pByiYXS+ITi1FnakpUTVd7qJxfr3GAs9+1SDuEwVF5
snGMJ+WikuoKWNElPllaugDinXolS8Vz7r66WDyWJr3fcS5QVi4szUB1v3clYPJ7BqO3a6PDq/66
hCD25lupVV7xC+UtGhkPrxHogQQyZUrKmSJj9UvE37DhI2hmsqu2LKUzrYvNLNkDGxy8QCyDeVyZ
ZgYXkW4Afyq0PeGYFNW/VEWZWWFuTR1R4kdbmQT/CgA9q249d38a89DIh6s3Fd8h6w7DQkl6Sz6s
bhivVa1BhMwp7vlLqNI4ykq4RQv7xrx4och0QDPxMIqWtEF2rMphWcRIOW7+bZhk1lDCR8fxxqIl
Q3j898HdaYEPmih0Xt0FQ8wCq5IsTh0eU/2rEurIX+1+Wxxl3B61Qdu6l/5OOvkuGTiGWgTlJ2SE
nQaJQ6QMRvYG2UKRgC/4YSjoENo8QeeMp+Fm2Csljhd2xH4TCk0ZmwpUA7RtNg/Ba4PuqlyfcAfH
l/3G5AAcoS6fAsZ4WrOdgwUdmRxbX3/+wf0gP99pcbseOZKerreS9XHfaHbsz+zmzkPmlSUS3LKf
PXaeZWFZQAMod9GFDpIs1Fvlw+SrY4KZAMimLhhf330c7YfC781ZakW6WX7cHIQW/s8kggfeU28Y
+OaEmDbXuiFiLiclSLvUstDEmjmksoljc0wsxqlPnf99kQVA71GYcOWnkqYHFM9rBpTVOTjSZmJ7
SpP+6AFyxsPjCZCLY4oBhhVaMxyw0wYgMoX+5ADF3PjmIwi/CYxWXsCjMjqLXchDI28IAqaeMhyy
Eu5JijOrh4f/KW/5XAIxx1l04Xl0208WoELAeW4fGpsY+7DOM7m6uSRl6tpygvfA2pyErJbZ9iWw
pkNK2S+830/HFGiyyzDvXmxL5u7ubZHlCeqbt2HQvfkZEPtUXzstcgTzdffnRF3J6/vPfGHiBopv
ck9IeKlHgIhzcOeYvJy+80DeZitvKAUx7UYfVS3ui86IUv2soz76q+Nmarg1jlcOa3EFTJMYXAmk
KyFxFIjy4x6Q+0EmGlcAfaPaKGND5rXYiBE8RHyf2GNHWuh28yAyCDEoa8kyja/H9NMYJZ5suDfe
XHMYUnDBOrAFDIIkT2mHUYo11DpkiXD2hfFYKPUvHH6w9OkrK8t0IhCbLN6CEeoREFUVFgRvT9Lj
tH/yq//S4NZnNxIRvZM5Hc0XLw0m8M6Z7oZQ45Onsw3VX6HO4X28TjWpBSLqDHdZ0WjziJKeRwzx
Wki1ZwUQtL1LZA0FuTM8tE9aR3XhFYShfJKWg0H2QMtVO5NFrMiNcNwAfqRN8CX6CUC9PTaYNqf8
dSgAQdjAP/BxaqHkvBmFcyDgCwU3sroqYt2MXnOEnF6JwHdud6J7f+3u0QEQqmaiXu6lPX4HJOXJ
rN0P6aEFHxQIjDUjnc2EUdGn7vUDrdTC98j0l3IbKESeGFyK3yprhcwdhT+Mk9b7n8DF7l+c3AjQ
MjGugMM0F7kckGSKyW2SRIiBD1Z96sxZp56awp3Rw5/B887zKdwvEkFv8N/tsN8iL7/23l0B7n40
82P6nJcH3HsAgxZdVHH0Co/toMGK1sryERRpJwfh+ndHR7cC7TD2blFICPyRO6AUoTAmo6DocL9Y
yX2eX4cG5AUbcZmeQ0usOFvgNkmlxN89FV2bpy48j+qXwR5CuCKeUitV77V0s75nMQ/ilxOUNm5u
ah6QjMPJcN30pLzZsA3BeGvsZLzBveoK/j1aS3A3rfp3IlRCGCrh4n5gU4LPaXuk5wCWj01p0iV5
rBKtHO2P3RNiYX5HPLjTv74R/CLhevab3on3FohP6P9u0djXu6DsLWF/vufIDLCBv3VExFuwd/Ca
QIFPhDs6JTdYhx4nAv8IUeJ+ihUtA7JHn6f4MHuyuJZhVQgPpyE/njPag6OpIjAnCT3YVjE8HzhQ
JnSf4ZBYL9Nb/dNp/prf5esOi9H4OgotHE/6TF8nCh8oT9eaZNbUhrNzX1LgNUnwstguGJj8Dix+
zC2zHBYpqHnasrrBFHupSLfFZ3bASY6fFfyFQ4qSwtvUGQKAdWptXgNUyciFfxjTg+mSv9L+yJNh
4RmYNC6nxtRQ0w6ExGbCbOhodX6lh8SAuC5kPxLVUK6HTH98hW1xcFvog2uTqcLzMHnYsPfFTFdg
hd62knfQPWhCQ+l5MsA1kPWe631BG5ZgBRfbfb1wkAMhXcwaFT4gPU/TIw+nkpNqkiH0ezLTc/QN
SkwzckxSBHszmqGXzoT7kb47WmNcLJGW+mK1uVo/DDP9S9riPF+jsMdMZ7Q+mC/deE4RNQ3zB/9d
wiXthRL9Lsf+GAOm6aIKW4jxb/Ti2cS+58f/ODk4ssxGMm2ngta33CZBQtjqequaIyIaPC0pxidP
ZUMBnT7zC3EoFtk37CVc34oC2vGex14PhM4XTslXVG7HxipHzsOjfEdgx4ykLDBo3n4p6xwRvOCm
1G8JnIF45/CqT7rSmUeAXhWzfcCorCt3IlBhLBfHrs8IBNAICuDjLPQhlkxQ5NrM4uQK47Otr/1T
wBsKVNpqB4Y9kvGkSezV54RRF4rrDFdjihSb56pswLax6kX+tNxBYNSeGb7ELREdm/fFwSuRZU7d
4uGcu7B/AtOCJAFxG1E8Yxu6F/acixDR0C9+lKHpZbczGA4YfFEXl30g5lIgKlcU4rX9Lqky6h85
4ZiRjoLlwTOc4JbafuQHg9vI2rXQ+9yPS50YRtkkGwmNfM3a5WSNA7+rZk0+Buq2VJsr2Lymin9I
ILHgt8HnFF1K28M4E10k4d/jVgVeeP3C6PGkTuEmVcITYh0mV8nIP6kg949MsIh9ErjijubY4zES
o7jHvx7TSnF+KZlMaJx5frISGxF2DoeAoAXB5Vsc4kgOvs6V0YRLNWAEwULaSNyj2CjOnf7zEgvB
yZbQ4Re+5J+Dv1NIWbkHOsc10wNhz7t8bj3OFND+kuQCDZ2iRMUH13RJdw1qH0FIkxgnMJyJGbMi
e7IHWuvLrGXkk8AGtB333bd4lglU5Ss3ooWzvS5PR3GYBDXmDcw8OuFOi55eHj7jiiV5dWZgiHCQ
QwKeEXHpsbj1QTWIW5oiffMGJm8/z7YlhN9eyqzxQARI+hDso840N5lN0AN0SaGLPxclf0qlhPn6
8K96EYqwQsgP7WzdzSfSREnOsNX5Z+2LPZv3iZv+yi9TN6YI/ORw/2zFZSIozZ4MNae1BHpDBJYe
prvB+iXX278kDymxeho7mEf7/tnguQ8AdWHAfXGYbWG8gm7v0lMxA8AEildqQQLOSTsR0PoSfohW
s0KkI3no/Nhnv+YaL1DHnG86DZs6PKqki2ebYWHYVKmhnuaO+lG2Qkai2AqS/UWJIJRTjHutXOQw
5FFRnW6ro0fSm09bDFl91hSUgs87hjcMIAliH6V3jxWh191OvICs50P20gbJl9cx8HZF6pKmtvnR
M0OlUzdYNqQQV5VCryoJ/sEEOJn6ytgA1u5b2buqIaDbV5csjNmc98lfjKYEBWR6Fjp4sIwY4+hz
siYdlERKV5ZKOV9y8IUbKCLvbBc9OOMcb0zjo2JZp80U/yZL/j5k0ZXBRkrdmT6NdsQhCNDV7XRe
fGicGN43zYdETu6m1VUf4HTKMJ59b8Ig0aV8Z62hqwKTnwQts2Q5VJ/3hb5ENVvdtuI7nLbtpKFS
b7r3Nx95klT+fz6IKinRbDv2wXWb9bca8PSztjxRnv1lH3tiyWa1+zoHyU0Pivc44yRzo00bvVwz
XlFOiEdBBojzQSrNKWZzWpEzS9gx06ljxbm0WmYUcNJOVGGOZswrxSAGIJbtqSuOEJA3MAi/1J81
xHsEy3sJu+Z+v0OFGfMxjwtvihmjgfqIe6QmPcD9OvEOgIiKA/CpPxXMCmT/K/UQpAfmXIXD1+2n
2WisngwyPIhh6k25JOy4GqXdeP9UuNVdsXPpxki6Ah16aZa6UFUbWTkVPkVGokXTTwAU2XGqH2Kn
ZELfSkgR+0ZXThL8CFhjeoKzud40rM4RisN3vMdDBeTyOkqb3wOUISc4WZNm+mLbRh4AGonDkxiT
mbRj4xUUblT00JvT2lGyAYDhZtt8hIg+yQQjrBHNJvvO9hAufscAt0r9cBt5tUfSYlkqdl5HWy6z
6D028HErn0IAmk326Ju5UaqwD2zXYAMd4kYc7hBGtZfkkpBEgygNLjbaquZqBDo8QPq0d3ZBBDTi
333aJVkTuBfx/qwvFbqzpZwO79Nu9gUYhMTeAHQoBEvy5FRKKIGhUBS/XVcHxyIqvd8lrkSr1kdM
QP9+T9MecnOJ8+EA5sYHzqTOo6nBn9JlecvROlomu636fp8ObyTohitSEhNBdk9hJaY8WaJTosJo
rVzHmuVypEjWSG5x/PkFAEFN/2c983R9mEEuhLfVddWIMRPzrHVvPwmWDhKUzvYbfu6fkjMbt9V9
PSdIpB+WKrfsPnOQSzZ/m/IHQF3ym++qpMzkGZetLS66skMOgSR/GCnv7PrJU6FjnxreNTJuPDFQ
S+r4WDAL4x8CsZicJXfuqTlHhDd8mBMius1B9XdoZXlUexdk6geZQN7MapOJ1UjNzOC9BFWvot5s
BL5lPyld+8FcntKHUAki1b5ldEZh4l3tvKAv9mWm9FQ83cd/HilUuEofsyoP8dRp6kkvzX+31mpt
gCWXmlOXncDvQRMhQ0EhqvoRusA9bY5JFOkDNNZVe1c4no9wsN1jbfxbMbsX0w14GeGR4Pd8GlEJ
o7QqS/vxPFgWsTG9GN2/gxjxgl8ssTz24AOJmsPE4VmqLa7P1OLJtnXgrd3R3kZdpG5QNsdKBXuf
do3xJed+veTJlpNMl7XeNrCLj3yrhqQrwtc7LWHwOXHDjC+urVHQsgmNlKSseiH+Q97MKzCAQOI8
nSKYwiK43N4SeM2/A0QxZRME5WFsaK13gopLyQAv7NfguK6KNgoQ3gUWMqSKfHx658ftHdMcWelp
F7VQGRQSRpvvPokPeHav4QjdOzHjRGyCRFIdttox0bPSapt0woaEp5SpbRmLF+rwRdk66e/ROZZc
JoS6TF3QjKrosxHYehj3C5pOwTBfYZZMrK3cJVFOezsIfyy3ZjuHqTAek65Dae2vtflCQCB67yhc
POr4owcqXrBF5u2raM58qe+oCT1aa9Tu1MPLCRlomuCb78CkpcqOm8yPHwYoZcxGMtcdDsZbR4VC
t2CxrFNl4QdhWt+pG1xiIUfYbjHQAhHKwO3M/pbUn9tWss0a0mwLIHBPbfq0zHcMO2fzku0dBtA3
Yq8RDKJFJs9sDCTbZjDZ2uDQsNyd0rmWTAXdYN4CLMD6Pxb7F8qQllKXEtgPDIGOgdkeeOrPTnaO
6FNx61ttZl4KckLa6vdAklCRmcXv3vYNi1Wnkuf46mPMKNwe/ZH3ks8WoYImfItwQmw/SyaKLdS0
TXBGQWtkXzUK3fxfPO5MougExbpiC39TguvKDkjZl/UMfUc6mY+KCtKfK1UchDSzhpsNTvBtnQgy
N7SaveVaehJsysAXZ6LQCmxxJ4j8/2grqiYhuha2vTViTuiC4Bzslp7QRCzGJGQ2Rj4Phnq3LUOn
RC39OT9CQqCncoiSr+n7V1+inEnIrc66y+zoX0delFYK9ufxrsTohRMOSgXH4PRlh8uu1TRTU4WW
NTCCXB1fQvoARp4ALoUUwOlYOLrJhdbNrL4r6H9NYuqqfMUBDpX2kHcCc0JNnM138jBJUxCjwh85
FuiYYbzg3R061EY599e8gToRoGaCmaCgBGB4RQnmm9M1s05TouFuRpcCVG7lBjBCvTMpT8IW6Vos
Ml6qCdv14y1EAuo9x8t/Z9eSTgneLhr1NS/1OBGgTohMYm1qvAXTXbdhY9bYz0QY3FIPYAEif+PU
yV3flUOQXrE+z9INjD6bH62A/Ig8RrVRxykcUSuvmtrG2E848fe+5xlmY8E/N/e8t7M+lT6Y8GlB
UKCbSBeieaeHCM/tLh4Bi9DtjVaBJxeCokeL3Y163J65+hUewmxZPMC5qWeFUC/pwnhnJRcPymXE
MSpcBC3nEDUhyvyU8iFt3OS1i7lZKHG+BsWutTsN+bqHZf/nERdkzlTBtKPY8pWbZjRlQX70jWsO
p92IEPDALqEkTTNZG2SSwmvS1X5OuuBWtt/Qocq+DPzAsfpJ2iZT0vhJin6GM+e0y2mM6fFryOpY
tz2K68s5Kwztz7ZCA92A856wIWUl7y4jUNwpsS6z/GyXIlUIWCl9s6+rc78zbdZrjJzKpk4mPVQD
db4/H85/m+mQVccGi6SkqIx5Cos/S1GKtDKGuErk0h7dkg5IunspOedQWJ1YLf38g5kZuGdmSsFF
1dRZy2px2WEOwL+FbyRICztzmRowdcD0nUNG0lBL+/oPFeLHXmtZCTowSf4XvfhEOAA7nG8v5Jkk
jExLl66Ex/LiY5Up4atSafPqXp1gSUwi7CW/aBdcn4md6rFFKS08RvO4pNmCNF54GQZSi4kmaRxe
AuSU87NBBjO4MKGLrx/ZJvQUgzTeWwlFXwbZFYkdiGicSWJpBu9II3/KV1svsAEQwHVYTvHx+a9L
wy1wldnGepK5TBFSP5HhArJ993txOwENUHNOr5BCbqzFwW+tPHjR503YNQyZpni6gLG2IaSM8pno
Ar48xm6+7CFeyxPiPgFow3G8XGLqHYJFgHTQaKqrdSw3rqXZXv1Mx2u266rRmWNZHGVTA27jC6PK
6ZdWTorts4e3jNx5ZPkkIJaLQmVbX2KXaDIwh5HMC57KFOTBKKlJQSPuHjxue6nt+nNYrKwPYnsf
q4n77/TdvaK101VPWbTkDVs1AGXthykb3tDQQWibBcezsdBJ4VQhmYp5rw8ZJ26a+CDllcan7MAf
p08JFiTUIEP+b+As3WFUB48pp9XLeearbBcdSx7NRBMHGHk3/zh2/cqJRr7F3oiK+zpfC78rSlh1
tB5b/oAeN6n2LdggEqfof3AocpFK8NRkSCyl2nF5Kjd49T1PkGPMTqFi/2okUhi+slXN0C39VERI
GrHXlpavwbxtF9lUXfltXQEv9E20AKyY+GLxXRJWtZVdMJLK6QSrSRVgF8UPvJkhN+p8yf1FTMXQ
Ap7KH8egreOxeCl3ggH5HgFaOHiPJUe2A2K1+GuQ+Eg6O3Z7o86G1f1yZA4DqMKt2+AU/c93Hjk0
GVTTdnbC32/qwIQzk89QsCwVyFfJwG+9aFBYB9GUlkYNto73ySj6ot0BQDTqoDrp8FiNWoZr/kh+
lZx3JpiipJvrzlJ2a370fnOUWKklf1qs/c5uNTw7GAhj9W+x6usjGbg1kxaAkWKGH4HqkaT9uHyW
AYEipHnC1cGwz3Tfu74jfXNMmAVsC11neA0nHlm6BMdkUvVa+Q7nx0lX0dk9UXok+MJAlIFSp1Vv
iNo563ov8a34Di1Pf1wond5kOWEwOukgnpQ1Y5TC5T77HunuLZwbbiTxHzMU0N1L5qKpTVgUtT5d
XCGgf9xnR2I5KER3Ft5ixLYRS4gwEJBZY/ftCaZ8mbD3BjzOkV3D3RLUcSCpXqAE7dybYGVSErky
T1VPay8Ml7F1a65VlBu4w/GOKe6QMiBHnELVVL9vobxyuhLQALGYFBwcrhArB5nSqZGu+zkTgRsD
sPQyF++kpDdF3LmS/umjU6z31EveufUV6F/T5fBkDYDpPcOul9lMWU6i3OVaipZ4Hgxd6rYbXtlk
zoyojEeRKgelGPlImBRv9Kyy/S+54Fdils6Yf/26CxxStuKN99Wm5+4AkHv5EPD36d3EnsrgvPrb
KgfjIF6uMMuCBp059M6iY7l65Pf54hKXvYoE+SpHYtQKSzIARLIbV5dteevrsNgbfsw21UJJisTv
n6PyQdk37ncfnQDGOBo8v1iMyaDtHyKJ3ZtwORZGuP80RtCxisiwuqhqviyPkuZNt9TV3ntP29dO
d54jomp5fI/Z0QOrKIKMlLnN6xrDbLMqHJin6mi/I29uw8yZwejK3QA74hEYxwuFH1qysiZJnN0x
a/6Cn1CcJh9mdj8S1RF6eXGR+zSbaOgLOhV/qYglpKeGChWANuauPgq9OuoU6ldWoMY3cVYMIoxr
2tKnVKJVxjMj7JiKeF/9loicLqCDrxILStWriAePP56z9L6uuloCDduAkAEBHaji+NOS0SvBZ5lw
9xhetrmxZdXivZMhdQLKkV99AOAcl+59O+NshwqCofDDjSFag5HRepjtk1PusVdnu+49LrzpziQe
nfG91UO3acJDHKoWgtqUqD66AvU0FOlxbgDmc8SZ3JmcVUU8K/jL/Khp++Ho8WPJfDhsFwDSuUam
1OtliCFo1TZVEHLfxFjoN35Z1TIzkzZWMEeRTB10Cxsxz+q1UrJuFvrw3AvKp5AREMI+ePPHhdQT
cYpNBQyUsT+no1tUYsYFcYjgvKtsBNTRkzAqr0azVYFwVJk+0KaBvRyeZdqwujAxtYHvl/N/jwLW
dr39nPYyqAMS8ElcTpqfmoqpMXDwZZejPpvuBNvBj3DPSrp4slgjSTQDd0rle1JDNmeyWsFWkPtz
83FiG+ZhBc8frfbGPJgGBYgA27Zy7p4gowk9Q3Y08efCs/22pQRrMK9xQFgVBK4aCqzyp3/rWJhE
iLIbH+p8eqewq2E3oOCuDo1UrPg0LbTjB+bFWo/QqXkGhgyNVanXPXI6lzO8Y7chgsEu2j8JAWz9
kQgX5nKYWHuPL4LbMUUy850ZIgeSDFZmMGKcI6QAtwSzcYxqa0iZHFozw3fT/SWaVtUYRl5DsYDT
3yCeFfC0WeL525AcNTWhHj8miUKa79Y9aUze/pWIUhQWnQ4Ks5XTCxEIWdx6sVsvz5SBx0Fs941S
T0W4u3o1xszCcC7E0zih84fph185OvM/0bPD5aTO+ihZizwofSPFL/S3ZxBi28UDT0FBEZMc11OB
cFrHS/Brfsgd/vFGdlwQtZXnghO8I1VlQnatfV+Sou1dVpvjMm17YTe+BRjimFJUx0CM+RqWQ0xi
v+tCRprfD+pDbqRw9Vi3rHEN8SFI2bKJXOY70YmLNxhxl0mZF9DiZ7CjXpKYbAdqKp69G1T64cZ/
7UJXltlj7QYrCFd1cZBsKBeoVPgi0ECUiCA1mFmmSIuxp/ZjQoCLwpsrGf3Q7HQNeWR02wuRRSKN
Hr8rssD//TyuqIF7DYAqaw7IvYshCBCqP5aSPFX+pDA6RjYJFAb4cgxdOfyoI3ltl6fYagRxPa0x
Zvfbt3umWBWxA28a4q0OyFuVIx8GFfHcbOI36W5Ycosb5pNV5fhY/NgEPXlsImmB2qRsDMfUk5iY
DVI0opshJ7Rq8rLUyg0ZQcBksnIzlXvVxZhclcMSysbrozDL6C5FxWji84kv1+MwQ4gDBzbbPT8h
FN4lc3m64n164ZzYnuO4jsakxzkvNlSdVlEo3UjzGLQ6eUP6ZmftbaTC5VNR+BiU2FG0yxqtgm7t
0+aZt+hXL3bgxLGhCmsdPtKflYlHXeLPgcqcaVUkE5W3v+cQ1SsrnvDlFJ/tjdDM/2joLuEyAS8c
y4Y66/tO9WEsD3v/8/cGu8MOi+OCdWFbjWGEa/a6Z2btuSFpaSDFm1i5CoId8/7gThk+U0d/VNPN
dwjW/YLH3bIIn5Ts47+oOaPCvHS5/spLLgMmY6YKA4y2/aCHibk0xwa6caTjeKfiIGbbI6jjXm2M
XCjNoxvt2d3SZNGnqtg+j/9AgdSIuLpV0E2RkZLrKP4rZkfl8IfV7+1XNIzd+Fsjz2Id6BY6JpvO
GR0XY0icwUrODN31b4oNhjOHLjK0cVidgSh/U1niUdoCbNO0cyS73Vr56toxOKoI5/a9wa0IOpnn
NogzwSUUXh/T0BzwIYDUpRgaVpw7nKQC4IJTfqq/aVaXwrsnJMywh0PO5smrEs3sJYDBYRQbkURM
DALyK2GZ8cULC2SBEu1k55HUAUlZzvTkfQRqVM+Xkrc+vyLDtFdq4qfsnY0VmDdTmrCyTwiED5+C
FGiGDDl1LV0MPeTJe0zc9AAavveqziwGbkhcbEaV0+C1AuQ6o9UAIfGTy4vB58QsMqKlMk475PvL
NTfX3XzKWLc4Ok/iMXoi/JZov4qRRx+JaqPPojd/wkGvct5oZYx9bECgf6Lsx81QSJwk1jIaWeIe
GBow/NtsSjpx9xJapRxDe7Dg5o/VrYkql8Fi4LKiZ0iNYkkh0meihDlPtO4gWi4uDQN2Ob/mehZy
7zQ75ptPI6YVD+KvqI99muM0nwnIu0hYyn+WEvfPeWWgrYYEBi+Yo6lV+BAnji6ydMDNoAnT1TpA
7eaJBc4/iSe3j+xDXy7oCSHpRChHjdcVFIkaI1htp3f7pfO9kMmlNFCUp9ZFmHiIenMW4s0fHHjV
tJ0v6fIBo2KMG5nvEkE2+FDse6ZwtB5r5LkANI15njYM8oBeA9wWHjo37AYbQjDTUoxaSCxRzSS5
661IMBV8lqocp43LkXy0RzopkwYXMrZWgWeLtKjIJtCBnAQgj5LTGoxt7SG4l7OsnGYZaRugsdyo
PHoXcYCg3Y9tYdlqYuEbSpnB122E2moqW8Rd0NaU7mIZQfcPXMnQ1n3z3bu/FFljEZTlmKkHZJYh
5v0IDXvSVxbywcVJRuQa4dIJ3/nQGb0/JW8Tb7EZTORSytlUjhxvzPp3TqWlxSlxYhzlv1u6sdU0
0Pyb6ADGM3hlrXF6jD5TP9dQcXLWWv1+YJwibrXPzlsWnT/YarBMME7hP38fLA/qHZrcDRrz7KJN
YufOrDnpXGAXtFViXOfCcChcUZ0kQ/nAru164FCqdW1u+CuL15XZ9sDfTLnv05OBOK4fFnkOfmnu
GbPtdD+08dbiGNfBticKvwAR0OYur3zT/74pxG+9wir8BvqszvGREfXCYVsfFzfR60zYlT6rGyUh
5RW3hmohqQuAPon/Qms3emV2NkPxdPqFyz6c1+jGs72QkeLpjC86CHmS3zu5egYaR71NlCOl+2cy
0niZYBwFm3VDq2Lb1g8DoyPCc3oYmkN+kLTI1yzKVovH489EpOK5LETX3vQOJU17RxufbbBBy5R1
0vYaG7+Y5NTGUPJoz4fNSlO2ScdD638+DkdTD98IhCLextXbF5s1M0owE9/8pLVhYv+TMYIuncAS
jVKOBZeMcN0R3kVulSyyoPnB6r8+Bzxl3x4RfYvc1vZ+dCshJYpu6XrX0ZMx2nZH7ClejJtzBU5C
oRrwG1uCTK4/ZUV1nRcQHe0g9dH2RaO/NIbMui8bb3yxyuRd+qXC2h4IGUPPcsydVrpMx0TZBhp0
rlS8OnmY7bUEGL2HsA8b+dgcTzDlwbWuXRHa7JGWGY4T4OeOBKjafrDmDlZ0k/4z+fO5LQAxo6bk
7DpAYprpFMq7+3bvkbxSif+J6Xp1djGquv2/cp8X6ULwTMIgYdHZgfEqu7ZCRCs0m+GM4xiRsPld
byqcjU6TW7SHZJZhsI3fNMpsqz5ThlqdrxA1jLwZwXphrkQ0qDMqSuWuNdOtW6PEqQL+tFR5UgOx
UAQznA08c2VX/nBppv2yRKjYW7buExBcjFPUa5AdAzY0WhLGfJlgHmOSkyP0IuexHbYkS4owKIl/
0ccJT7WADdtYKP1JFQsAmFIsJNdYTP2aShmKDSeCHj8VdRX7AGIedSoJROAIcyg8ZGZNk2XAq1oe
1FnBBLhdGB7QbfTUEP50JlS0saVXbvw1rClYbrgTody41a2z49P3L0oR3Hd8pPFtuBzHGSqCZXlo
PHcjCW9MabkwX0IzF998hikVwm0bo5mUVUBdCcN4xBpXpAoI2vmHGjb5rD5Bb17e3i6P6iq0eEka
VGenkJ47Q2bkWTrUqGAK77BPwhtl0ZJiSKm6LIbf+rjyc18VO58RKh6iAHcfinZXwkzJFpoguAOI
W0LvidBVeEfUSpEV3SZAIPRo0yXL43F7RwNqMtPJtgNX0rEgQO50cfm2qCGOTkOOmAN59QCLCtD+
xwJnB5hqiJNdCtOw7d3M0amUZlrZfcY1T7T49+T6zsATRwl2k8RKjRnwXtpgijfANDub9TgYSuwE
EBaOILVswUDcepcT1C4Y4YtZU1Slg+6ldPhnEx7028r4DD1Ko0TGvp7KLtedJQSBKXw+9wz9MBWP
z8H/d7ewvtoy6DNodmFEC9b6MN10Gp/BFS4rLTH7X//NzimZAThPwMygyStHle01FO76EeHi1Kkr
2C5WDdrp7TcSpnO9sgXUnQCnF71eqgkonkPiww/1mdZyOrDHbkqvwYbieLyuxrx1Fbp0jLfs35pI
zKQ4B+khqRxmMnNdVURByzviTjwkdYlJPUAG4Dc2pmGVKdoES16g9vZ+ZYJuLJVFT2Sts/NVfKiD
RXOqQ9Eo+ATd5KrD0CtyHC5MnfhyLVCQU9wIFYNI0I6a/R+cdsIKlpp4Rpp/6SIhE2AgeD7quunQ
SHWEPsG2sm3ARYF0nm4j5NhKB5k9fl1BqgFEbF9A2wc4JdmbU+IPutzIbyYzhEFNEVV3/gnLGBoo
syMqT1Wf3GDxtWk/QBmnHAWQqQB1fDoVqVFx+pMsL07x8N67Vwfuo3Uo73n4sasZPIGwO+NIsbe5
xAyT+zDJiz/aHmmQFKi0B9ema6Q/y5Yq54mBCUZzq79OAZFl7raHEKyJIlTDUf/d1aR5Di1CKnfm
+sATLZwqM4n5wjEHMFI6V6GneNFnHMG+18acFBzPSro2mGNccXcCNJuWNlibkhsZqftXhbB33AB0
BJBvbNSJOyDHY9TJN8ENI52RCBHpwWcsgZ7H/cpD9GQGMnChBk6yaptDrRlE/uiDI5HnBgFL57G6
ICylHJv4ms2/2cim1bI+DNiEGpw9nqfLjN9LBxWaQdEyELjVnn3bTHyyGcxghO+ET175nJCs8XSL
bb4k7EJZLf32EcUW5GErbX0pmWku3kg9Zl/pcatpkhbpTxZQAGjfEblQM01mJQPxaKNMhhdJ5Nwl
jCWMcVQHFQGX7GOqrMDyl8jBk3cJWMCaiJHuQjd0cjndYQfjeDyp4an65R78J+J5kmY42xpC3cwC
nni2iBydEcSbsmoznSCoBpr19A2gnlYKqrISDFNYZ+bQG6hoi6vBt3I1dJ0W93MGpJiV0Ptb4EPH
dpS305EKPfz1dRvPjgdwrl352Ru3vU6L86Jo0eBIuhQvnfUu/fxFs9QRjRs3IbLAvMAV+kJQ8LbV
vXcRFgU3sysAzUAWwyG8uTa9PW0WGEFauxCpaD5VKuOlzEMGfzwyby+S+q4xCDit7hPF8EWGBneB
ClMtmaSsmlXQoDKQkHHE1mcfVE6AnDa3PVHwiitvnwH5bzdVwLlsNhA2zjV6/Z6IbxqUUWij9Opr
54BYDBPTYbLHUP3MjcIcToP7B4Yhh/9hfieco9veeIxGlB3ojXzLjuSq/IQ7ZfA+CRzHcgpm5Wuo
jmmd12gZN0YSVoinPvksDX9BLPbYFclIij6vFNJvYpL0CDY1RlODnY3gvsi1diaX+sW9E8vnRrK0
ygYVvdZ7VPPgHOGFShCXm814+EJulQ5PmTzEf7HmBTkKVt0//2rqnBKlhsOodbnDsDHUzL+D+2Ia
Wk6ZibRn8egt8inq1tQo7hjWaPvDJUQqPRZmrXaDFFpil1XRvzimu2Z8n5MAUEyNhmzyEYhDPLBN
QQIxnfkS8VY+qBHEB/Tqd5+2NOFPMCaD9Ha0OO5ldzNjnGSanMliygg2c+N4Pt4B31sCEjMcUDEi
a6FsrgwXJZmdWpfepFGdwKf6r5tb2csv+5qGQ4p8z6PnRJOgUKrtts+vCkVpu2uAdYhwTVOiL/3e
1+Ucmrno76xGUEO4E+VgQg3qTEmaxan1wkbJrixQg8zKLmwgYcsmW6kUhcxCi69tpojAKhk+59PY
u9zgWJR7NhrCNwiTPlSrea2Jomf6Bz48oD4jIpd2fl7n5rLf/JxrhKkPf8rizTFnDkCBvq6cnnPr
ydAcW6SxNVFd0JLcP+doffLCdiMuHduLRY7pp8g1jtqN8DwSaDrlCj8wWu5oNyHZVIV74lIxGhRt
B7qQ599yMwkRfvvneQsW8U2w2OJlWhymHwnpd7vMnFIg5sxzNe3cFsoeiB+dWGEE4qGeFlOcHSvD
TVOtBbin7untAwSMnVTQEK603mzpJcJyuNJbNK+eDAxb05c0ojrKqrTTLq7RAE4GOO5ScQCQruce
ReYxdzbFMUwJQbluUCrTO5hbhZiEZrPlOmWYwrWS4yJp2zPvjMPqI7jK2fSkqqAu4mI9uD1SPy6S
AEZNTjMXheioN4yj9FzXYQVLkliP4OZnxmUfYjEclK26DMK+1iIn+nAXSI7vrcQlV7uAAguDrwSP
It8+dqvWNexAcVQ4AnMyPRjy8BxkrLKJFaMlWEHoUAD+ja5LDl8bVnl6R9yPeod6OtJrkfgXPvwF
TmpnFoXeQ9NORihwRX8G2U3Ikz1JU8wldV7/6dFdfruP3Zg+y7peVjuV8X5EVfEGuORrbKdej/PB
EBVtxKLqCJvVFzRgkWj340h7nKoiRw4M2lmxKCY62qEAh2YijFTxaUwOhJ1vHa0ZqYM0iXyQxaX3
n8wu3tUsHy3TKirFa4WWJd6ciwAQQkk23NsU57u3BOVKYCMSFJkVjZ7kW0P4sxRR6/0vTPUFswRd
J8Vpmub0kCvEWdeLr6yJ9L1YM+ruibLMZzHF9Nqz0MQyecsq7p30yUS+Asm2g2muckWhC25JZec1
U/yhd2etTEgswb7CiXiDPrqwA2ENHI3QGTZ1vuDPpDzxqLHhN/DWgcDKjHlndcPaNntjnGqag2ml
ssK/JHGsshCa3DmIhjLNaRD58t9LmSr+MyPhwd4rQcCcveSh/UxPr4QUTUSQsnfmn9IxRSoYZ4Pd
ZnDb8A8FWM1bm+4suU2nvzHI6KiD+KlSJLeJrJcGp5md+bx0jJ3YUAgiPmKY4ZSxcUtvGWRLr5dG
Ru8WwVNiIfhvUdnw5t440E7FBtn0qzNGqJM8mjlRhYd6Nk22kE88R9yXAur/9moKnAVamuv8i/qJ
LDKZdKrN5JmQOE/R736Y4WPi0pxHO/aK7aOe5YQMbjSTDs0NWoFxk/S2R2f4CdWckMraqFD1W+M4
mxxtipCbq/CS5DiuPS6plBMgkMMve2n02dxJRqYAvAbsCXdKm05x87PNfNtb07ir8/K7lrURC1xr
URnH5Ma1p5tosPl7VPd8iVGS6f9Q+iPwSn9+bRXSnPFWIdL5FqSGcNspB0rFCmyibExrrBCgBr5q
Bp6vkNf0VTJ9s69T3ka57QFZ5OchbuqFfEPtzxtFPL79LRYeshmyup4HOPBhmZPD6akGGTAfmTfD
CGVuqOhYBrZRvBqyikoVuD5qGOp+FMheJKzI3fBXbrr0kv4nXmsC3TtthGGvTpRS3hPfi9LpI/VV
S2UeWC+eWHUUfxRn2Fv+YEqA5hjG0JnL89arJI5FF9pWXkaNUnE0/8AAUslFcjCtZ5FPxclgPGIW
FBayKWwhzCSz6O4zJalrz3fYfWlsj1qyB0gK1T4pO8s8rkWHlh01tKSfpr+1c2G0pnaG/62JBUpW
YbfdN3ytXXk95VUxXIPRwt2MBCwjkpojHYnouEJHv2SsktfjeMX6Dnq4a7xTZNGeeP7kCD4GUpEc
7lwr0mHjV/gqowH3talOdaTKfGjsV0dfruEtRT7lHMAPvWvQ4gANItII4zrQnK0UoADyUfWxVmWh
TB/maWw4UNMyKOorwbFcSY3pzkRUXyw4S9ro8FcMMo1NOR4zhMT5SckiyRmUb8f3TfXjeC0yG9HA
8gMlpPf5LFEbTBjUpok4U5kjKVY8R0f7RfLRxu/1uylkv/a0XMib9P6B/DTFAedrUKLYlTtuN3WQ
hlfwJ9rgDTfJkhzgoQjCz6IBVbjtBLgUw87qqRDetgXLhqffOZ75IDYZuRpUhJ19jhIjSubue6lI
PKcTL6MdNrwO86dJImD4qUoMFXVgwmWXBgGoEbz+HA1Kt0kXzaPASF1oQbx3o+C72tx4qN3GNmyo
hxPq/PXzM0vZA77wbuLH27Rr2t3OpXbXswZCrdeMPLzN7ioTM2KeXPg32ZqqKiX40jYTl8YSdSgo
oCKi+7thwkNNQ3JqdzP3rkXPEm8eybIxcS5t6jAib2sXpxbv3/a/0nXoF3qll19MMARpUwu02X06
eZ0whJcGLpsajf0uJnP2tHQM7A/rJzyIVA9LxPAlpa4oDqvhwfmd2rplPFjIJsyK5V3eybxiEYek
IfCKleVq1mMkExXWHeu58eZs8bMAQMaKSR5b1Pxy30m3/RsnaLvrZ0o30VZwUD+nX1glT55eATxp
YVoSX603o57MHAQ50rx0O+F+tFc7jzG2BD4G5LL8ivNu7XlkoWmAbvwZXLu0idLdLP+KAUONKBM/
/BEA5IorED7u9GwN4SEgzYefSHnI1Ww/vF4CSzQIb/p2YJyieH3UPega7BDleZBwjIpoY5OTn7ly
TalqN2N7tQJ2MTCcIoVda24QVzT2fx7QaHEMGlxPygz9EIHvkU9JenkSLomxhNAXWnh8vKuc0WFB
BNkAWeHuoNkquMV4OJhTsEQfrxeSw465Bkjdfdt6KdFsjQXu/k0vrE97wH/R4e63aLASOrIuEH7U
/ByFI3ijUMrZuwhXqA6falMJf0td/RN932jITcF8ps0hw+hKbqvEKnyCT8cPtBiVnJIs340hfDE5
v2Dr+WhymLOOrL48PxOXnPylWBoROjBdbRBByZ9IkMCHyWHLaINiTtN9CQjEroTH/u0wYOI0rD+9
mbK7O4LMJT7H5VRP67J8iAVAHP9U8Ockj+U+uT/dRaHV+eX811PW5mDKsOVrmtkcTGXeTbmYldec
Jn9fX5dJPPWMacykH7ZiUQggsGtaJiegJu/Ppzt7nxlZF5VvIA6HKLl5K8jHl1HwkHuxdwT5kZ+d
jOxzx2KVh9CBMsdFdP7ylEsqvqA9TU6OOm417a1t98gtrnp0V4fI5ENCXBwh4ILJ2lXVkD9BFTta
PaVuQIS0dnKtlSIO7E9X+WaIUdDlXEwJcYOSVwn+M3otpp7L1pZDFNZxod2GGDqh7Nd6otsE1kO1
ZB1PomHwTw0BJMHHoY5FUkXCoOxhdtnj36GME3U25f++ZxWxLZ1iqxLypvuX65Wt/0z6GEYk6H1h
9ZhpHs+MZB+ubTMevE7hrzgXi/o/Ngb6boopfHYHAVgx8tr8n0J17gerYn1GYjY5wgakvoGcuxvP
o4EyOj8O3ckUEtjNEk8/Rl85Po7mqK8ZYVwi7snw5P+zt7Zg+g57/NTgYdwysBHIjm57ZycvCKxI
UbEPz9q0EmYXs1B61ws3bjbiDEGzVj22N8hmWLoWYV0b9Eqi5CalYzxZXGafCxtq+GSXDRfBI1hh
JqhmlUNWzhx1wsR6LlDmsnGMWQiapE+lYAE30yINpJXS5+fH3GuC9vNGapoin/CYNh7b2MmzSC5P
dX1DFxxlk58EenWB87tiGskwSiJVrDCGYwhkkEdjPb5Hr1C2HfkI+ZfWMyOoMJ+0TueaENH525mI
AvOsw8KCWDCspNRjQMv0Ih3ndR/XGqWatSK5pVQJCRrr6w0oi2LLtegYLMq0mdsrKX/p75GTAdxv
Acb6w6C6LyODohMg61oR64BKrPdl18tVszGeDmo0bamkrRI4bwLiddJqsxo56D+VMAuIzMdPQlf0
IIQBcQFl1cRXgWiOX3R517ZS1QAz90I/GztGmSNZWSF7b4XTtlSWzGGGwY+Go6Ql7SewF+yYrn9a
TXweWg9Ut3Mi4Js8S40xZ/1QHjaTorFZyRZRGF0UyYoRtuBRqEnBtfRZsSogoLXLSu7rQbaZS8Et
sYZJ4yDjJeK6jPwdP//LQkT7Us52upWKJVy3cf15SemH+ZpNeT4mgzVK8k2RTnm2RstfpBFvFSVq
zuuar5WEt5Dv9BXG876KCTuHT6WeRgTX6wHHfcSZAIR5wApkQCpDGb9JWDyq2IowVcjVrYRRTTDt
IrKa/I9JHKdTwv7aLdKVXzgW8nuyk4cEJBC9i0+2NyFn/q+l4oa7JQIV5iVYyBgdomhY78dA10/T
RKI/WIMZdsWOLUf8kfTXgcZnFKD3RWLP4Cq6QvGn0aRXzNToL5PTFKLZNDuTCLyhXHkG2Xh3qJN/
YY6YEE23jOFj3dB9h2hLceAMQOORrjrLMrI10PaJkDH1g6GpnUmt5KPnqbT7RsokOXla7rjSQl6w
LnUzs7WfwDWFNKdpfgVI2qBnnIT2mjLb3AnhnstMReo/f7D9DWJDAPDc+sya/LOgBex2P9PpGia+
jXkHC22F8brmKNWpeK9V2BQFJWRFaEMmANk5XwxPV6p5AGdg3AMLLJey3LAICbraKqGT8laDjRbI
jselwdZe7U5T2jXV9Pctv3AdBVoJNsmM8SYsasE5AFxkvZI0sreORoAC2VdePAqlvnjZXm91ZJpg
OL7jkFfQNMvzoDANS1cYehA9qHlaeWhTgfW47W3AG5fq73LTD8VRQgjXzIej47AJaF6R+ejUbs8T
OmuKRRdFNbKxlFZQI1GQpo1iGVbJ6AISpvrEyj15/QiYzWlyBjYmh2YY2+WP6LmBWVhjlhtPn4mS
Gbg74iW1/Q43tGKhcxqfIH1H7w1cum7MU//YQrFkMpvWJutGOakMA1E0GgqMqgGM62LbFAHiFTd6
EPCkrYOX3gzUyelz4M+lggSnJ7WZayqpYjgffM/In+ItMljB1coD260XFfNGlmu2maREWaQCAh6A
UbfjX2g7F5/M+H5VLS+1bOM7/gsq6N24yBMLdz99j2xcprY9ycGAZmd+fkTHiJCZbW2WHJzDuzGN
+A3+pObbZmWo5sFG95lNXGJJbfu/C9OZjcTYnM1aRwU+opLFwIc47X15Mp2eG6L8imUiVORYI0Ez
UrUpKjnIhNTWpxR1x3we3wMe95v0aPWnghpQpsnJAW4oVL90LtYSbkUxowJJ5ksMce7xh8OqeRQJ
AUO2z3cGCg482jCHYmws3D3VsuCG33uwz6xS2ZPWbHofCwZVu9/e17ZGaz1hyskHNOa8iS9VX0An
VL85tvKd4H3NKVDHhM6Ws2HfrWIEtC5jgx4BhJX3G3WlIh93heJ/XGs8fHyHf+/p9tLEzL8Pd5Bx
PasK7fgAHw3aE3uUuXEZECEw+EihsH53qVr8EZI7qKHk85fC3im3w4mr5oCNZW87y7z7T87y20dK
+705v8aEhqFQzyKrapewrijj7RB9rkS0wBpB2mFBQSSMdV9thMc0c/ZOF3swuD3PtSkSrNefT1Pz
YgHAYx6BlCDaXlIaR/Lior7y0ZDvM5hvPBy1xV2n6WvjbnbSebW/lr4kpouhtoQSsBpVQqyyhsxk
wG/77x7YkHnPXeWTNR7pb/MYKfnYmwlfc+1k/mNKaBcWzKdpqPjhOt34CLtt6uA0/+EVSW9mHwV3
jsINrGb+RG/GnD20mHqdL2t1TFBRUZBtRdlhgvEXsg6QLfgf9VJi18YiJwLFOBidJlXTT6XKXHfq
kAkMR97C6l+wyfNqmaiWqkoZ3zqNcAvABguHTFeIYHpNW7fgxgrjKTx9+Pgk2d7edmofVsnBgm5m
LVWTFJIjcAsTqdAHLR+p3tahadtoiweSVY+QDCYLJVo5A2HYjB9U2WjBPsE0nZz1cr/FA9YnSIbp
AOxVjczlVuQH5bCSuoZo/ohjOg1sNyJrjT7E3j3vpghkFjAKYYirS2Es1IkHbR+vaWxDUCMsfDnn
qn1hlSOjLsVw9cuejuzvDce6ORTqzMjjbpyJCE78eF5PG1oAK+207mqBCOJdTpjdQSadIhCmV5VF
6qUQPbrOlEVIwaITfV6sFv5/2bETm5soQZ4KTsZKFAs8hRfaAH76eMZHtjw74kZEQXjcQROoIXrM
6QZdly65Saa03dEUv21QuK1IdphqcP9I3M6tqdgH8VizpO1aOxb0hS9BrU6Nlrq759UJ68fIBM8n
/vjecFMKAv8LVEWxUkhN8yeocrnDGCbjNBGkc+4Ukdrs0i0UWEm88FzkY/hTCOxzOM6A5b9kgWQq
kVHoQyJ2LEh+gO4mQVIsoAM/DKkAQIWxdwNe3qdwT7svuav1yA/kq89FztopVKGFqTy9S8LS7bnD
KeQjhlwVliQ/yNQFZCCyEiU37piLGPyX/W4i+7xInnUzw8zLt74HlaHLIOnFr+NOKqOajJ+smlqf
GTKjE0U42Y3i5QlaG7u1JiZBy7TtlZwhTv4b/SDPRVVjAwxALMm8ggA/i+cmJJtqFH5hDKiAkVKl
u1YPWgRBbk/DI9wm+4ZD43vpS6140gWn5gpyQCLAtEvKIKPR6O+fT0uO9uKoq8lb1wp8gI9miSKV
1hkaCno+8JmOVvot8/FVENPfZPIxoFXsttiIbRE8EtRQ0iqXIdRI0Hls9+/iX1t5m/spX9ml4Y0F
uAKon9rmnSpHVXXK/0v3yy5gVQDsamw76fMCiuIleJogXTFXuLMb16gLt8zV+GYbSbeyQD28D2ej
t3Xngg+7thIXGVAjv7tF9fcjBGRbhlAh90I/29+30wzOIBSKU/6f9N62GxAUwr3il0U8YCPMB71R
GCfHn0lBD83yUaDVv7bLTWs6cldMlU88+4d6rHXFGAhQQdOwJpeg3sqzeOrdL5igBdQjITJzO7rj
xn82DkRUCr6E6lBbs+M3uYgC9BwAjxjYGJjbuDZnE9bd5ActK1cfKcUYyfGrCSQJBchVE5HzCmp2
7VGraoc2S/BFOggH2Vg1usuwdJdX6NyGmnbM4nqvspP/IBZyyStNpxPGZqXrXCgP/q1SE3cXXW0g
5uWRNEAI1/hzo8o7hc3jSu4nwOzGJNfgtr9x864NC03F7HskLGhBEqvsfXgZxrh0/XrQ2+xhLIbE
8GKwfuSWdTRSv9rPVcqfuIeURPfQbEgliTl351M1SPNPxtZEVJyA2aEizIWvQOsNr/iK4psdj1k/
/EvMoPw2QZAyUTn/44mwIKw9+Ai1BB9VYFTR2EmkSOaIav6JePu9XtIGV49uk8M2rztkIlWH1GL0
Ohr65y21SDlf7stnuIi89y8j55c9cRGgnnJaKH4Ow9YKQmmSdve7abePhE0tBLgJ5Td9BMMCEyo4
oz0uoGwBMVwh1O6Ppzw9xAxktD1cXke6L89V7UuwA7MXqqKZ5Ooz+qlh4uyEijFpn7gHGHt5Itta
SV4/oWOz47DTxbOWOD+dYuIaDfCLVxowuzOvWAcGM1LpR+BH4Wa7qbL7sGnomPNvYyvS2Vep8U3E
aqUig97dzi5fjcR+FiBGGwSaGur0r8Kzi+SjvbNylo+aTQ99W+WBjvysMRgKyDrA0qKUY56Ha4Dg
CU3iiZpTpssTAObFSPdddmtXIIA5GLtTQ0XA8T4rQxYlWUWfRCmAhYZnmVG+NWGAbJ8hR1yCg+JK
onWpdnserLv+enKoIdh7WoaoJGmenqiw2YKgvCLz4McDcMhgg/3dagLnqutKAWXcwidzaeplapBx
oViQryAGBk/JmZHOERhAFqu4xWwoLVFxnuBkqkJ61HO3LEf+Z5aZGg9FnCbpzwROPpY4siSKEQyF
TsngfQJtvZn0WdIpYYsiVKa8iGVV2YlIh9/lUo+Hr6LQML4FUSh5FpjGB7YOfzHeFPR1toJnR9xh
ANE9NBCzUPfKs98z2uL9Xa1wl4nAem2AAyVlVJtS3VJAvSCm5xPmdcXNYFZbMoapYMtFfQjg6DLI
OndAytwh6aToFWJM5NI0Vrsj4voWtTV+tH16zEzfgojsnqrX31cdxXGzL8pP1kLNouEaJbKAmfuW
LW63ClLsxR9bigwcJ5M0uN80ckBctuX2jzMrGFJlqtdF83eyeT4N5ZM8iRYinETnCkJW5JAMO0tY
5VeYxL9r7RVfstfWYOeNvIxyXT5LBdijMvGeNUhhN0txczWswiJk9U+/VX7ShNFGRMfbc3Gxb0A8
TSwX620T332boBdr9GELz0SZAjJKWcHCgQUCtM79QGdraqTjE8sUb7GZo9gvZ9inDZLnYH+L+zgE
g7uyxbx+C4AO57Nv4qpLTpLRCe/0+Fa/YPVF+ViNXA/+AL6fs4Mq2JJ+2ntNqlX2kzXiCus5TC3l
nRBgTUax+WX2NSdyjILrsV3t+aegmitfZYTsAGL0A7rC6KSz5WPcRQAGCS0cMBnrViGlWthU/S9Y
+ZlhB8Khgnv5A9VK5PY3kx4GM7glL83/qj8/QeeAJUHwtTLZKc2DSO9htu6Mhr6pZnMT9mkKkCLK
5SEkNpbTB5nQHtAOnqfw2AHdOC1jLELvUXPf7Rgvwqd6cCMByYVtfrvYSmjOtenFvNnXeWCUzE/o
H2zwt2J9rCaiofOPmmEnzrUsc9xT0mmKoMbJYEsYLD9LTM4wr2dBGwBkDb5uglhcdYO2XgvTMgJY
DRajEI/io+es0FlNRBGKJN+0+zgymT/udPsReCrjQYhP7q4QFDEtWmnUkCj2GeiiKGHQt0U6n+9J
Guuvz8mIXcqVmQsWNDu2EVoE803UQgeTOLEp3fNofwGJyU4RjYHwjRUi15zPgKrXtN2P81nf5lqb
/8WRb9WOnsNFPeNR5F+GQxi9DCM+NPdGb5Fpmm+YNZqk0VyiRrOkCIDsBPQAGk+uKdg/J9zYoqKL
FVE0OX4LXpxG3h574WNMV52eW5D6o15DvdC2/ySrOW5upv1PeifdE2JXtCy0omc57G08eoM2p3pa
YSTEoYq9IohwXHCdc6AB8n85PsDUZc4erxhXW+akM6ZbcTZe8S1SkPh9+K+GI9VH+YmKSsyfwdt6
+w9z4RVoYYqndwf0bk+yzHHoXQnyoQQIhIIpkG7O85kEVlkIhR00jiwUehCrqDLM227N0rrbWmYQ
zDVKSGAay9M9sy/Xze56wlo1DGcXojbvR61l6Gm51NqgF1tOcsnqXfGxK4dtTfGmdWRAdLTzZ/bd
StUJY7GztRm8V7up8y+97gUl1OVNw9110+/OkOwYrOaE2NjPBoXus+s5cEJpufbWv68EkpPJjuVY
m4i0FrCmodFNULcFMZ8XN0dZgaGNZAarkQLbV4xqMUN4ARNIcv7ERAoFvq544e0sf6QeEITNmBtG
ODJa2qkOus/EsY1TCAd0dZ9G/PicJR6ol+8rsNYZuc8y8fUV6I34e/ZZIE2SfMgVU3ERsqiwngXm
Z2oMVB85XH0Nfo7yGmgACSyxoMd7Zz0PBC1PogKG9sqyG3XmYAtHm4GS0soqgAC62LQG62gOSv01
a/MZssmv47fi6wRi8cWuXgBIdMpSAvIpD9OV2l6JNUqcRObT0DBhILMf30IEAw9QcOyc7cNJD+rO
hA0K58ZUwGOCSFx2NxmBpm28/hphVsAMGyH1fhg0iVfxdjYL+MRAzbZgj14N8YGQoYDDMAB4TgOV
YPqkhiVIkPYGRsh098oYus2c6kLbp25uilduIjDCaBPXwj2jztzimMWhJsCMHKtlTT29iNTK11F1
QEdIWHd/InICz/ijENyNnF1XxAwJvdrsOwHyF5sFOCmCYJdtlSNyATfGSWfJ858fGqs2oaikUCw4
2PECOkp8RGUBDuCpZBOkmnz7Pl0qQCq/TBgHJb50jQmo0kkj+Dz1dwR6i6rcK10188bV6RYT4ZXc
fpMiG7axBnmwxuxfYHGMshPbVffBvfTfKBZCf+gpmw0ygAbwi2oDhE9SzWJY19jKTc7FOXX/1gRf
AHZ3Q0rPAsmFwMJXTxgbIU5W4yjerHW/LeIuVWHbavsBM9KyMuh17HgOY4SXlIYJZpf+d+TtLG75
gyx/98zh1qxZjVqXMCDoKiL4F7MTXt3sr+cZehZLWM5NnfZV6S0ariMI+AjjJ2fNU2Y7b4BU5QrH
7PIBHs7lh1eEW3YCh/TuaqJgkGKFJzHB/IfvrACsg39jv2xsmHXMW13MUczWfnbMS6/Ix8Y8fzlP
ex06m7yVfMLt9tlFDvLR3DQrDOUVCfZyzbzGBZYJ2SYPsrEebiueHNoFIp0gnduOwI8269WgkIXK
VJ8PMqnIGedRw+YX/LrzdQifJ+vV9P/McM0DZhqGM9pB0LPmuCwRLDQADthzroMSHY2zDfZfhpu4
gDnTXYDWu1OJ56ybLBBCB5HL2vwGeVGj43RAb77mBe7mZUXOWS4hbURYjC+QoM9rdqGOB8zFQIuk
jpDcEDJQlkaYpQql9tKA/qmT3hjmf/0pNCHm5ftC8dwTDG3m6GY41qLy7ZcbljrW21pplVF2gEPG
bpvVwXn1uDSlNqOQE4fRtTSZcItTLok+rE5LXEN3eB+MD34amR2GZvEWlKE7zliZO8m1prSx87hB
HLWSKdUrzL6FKTexCDZ3SCQ3vIzwBNq2PE1kMJXILWxC21Dwl1nEgIDvjUW8F2VDYmtf49fUPChV
8QmMvTCVmGQxla4EFOpDDTxpHQabCs6zyX9JlmcrGNxrrqMROftnPOxhbGiSAL002RJs9npaAQ58
kzkBxDSayMCTi2E8lxvW3dJKxYDOTSkpByS9BxcCb4YjPsdXfF8Z4QoUEN/Jss9XOp+i0rq/11xu
Vh5Vx8G6EVwNeHGfPmW4xchf/trHxmlRBOsVY8o+A8MJZmj556zw3kTRjOyXzVaqt6ziFSg63YsO
pP/YMJCAPx7V1Tn92N4GNfNcS006w3MS2S87Jmd/9yxpBk8fWBtdVF7tb037T4iOInBcpcod+wZd
p+kuORoZYsqAes9jng4zwgBLprg8wDYp7vFGy4IfkL8M6Ql9Iux/VD4K+/sHm9exrvvOXGO+5Y33
EFjq5Ci3d3yYJNCFahOBFWDtP5Mqv/CrDC4T36ubbJMwYCikSY1iFD89llherFVUql2aoOqcETca
8ThBQjaxBfExHyXqFgkhjkqY9T/0eFCm4WjYlyjbp8p6fecu9XaIsPlAhPND51GLgSV+h7FTj+wh
GjIqIhKgakNKIhDRoRlqYEAVsXA0ZgJ485+tak1roINNwn+EGRUcI4vSpEjsulivUm8wAK4Lo8AB
0GrpN8YzZi1DX4nFMjHV/eeoPLIcUUhJ6Se3Vxwa65EIQy5cVPPej8Y85mrEI3rP4BcWbt1b4ufX
vv3Dd60rFYFUv3XOUitFT+gh6IkPXi4dGnBmdFsFDMe4Rj1Zg4fBaeW/on75qY2z1je8iVu/wluU
OtqfEnmZE2qpsmTBixRXEGDuWU9N67YSZGc3sg6QmihClO8b0zachnwKGq50xIc0IAGe8Fn2Zq/J
GXiEw/j2uAeT8Iwn4erjRT9fnnVFt9sOPqZODO/QiZbCReQgtC9uiQg3+m6SgyCDJF/7i6a9oCpk
T3bM4s4N4eTutOPUgj2xNmHlE9XTxesctGgTjpemsgFNRLGMv/v5rVd4MEA/IhplTex2D2eyxL8f
bSHD5fpV2li8JAD9HKcUFL7yktxMwhKcFJ3Y/aZAqkQ2crsz7+ZW2Xk6AAPA32pPzKejPsxsFqht
BL1cwZsyqLxWxV1Th1ZowM+YcFF+C2sAMBpD/FkH5n/xzdgVAsaoircGM6f9/BDVoYqIFzGI2lYy
ZYP6aeR7byMNUUm8ejT5sPJNI8HGkDA4Vl/j7HfSCwBLo5Cye/y7fl6NmVjSNsUuIW/FQ19t58jK
YMQyAoRC+EP+DmqgTKn/745wOVHoNadW4SadykwND9wmxK4WsaXMY1g6+0WL2/6CknwCDUfPd5HJ
lHwd+fJeeOYcXVrcxgxbWWu+cISgL1C8Btqg5vvLerpyk+0+63blLIWUyCW40eKpufcxv2/2nwsR
pA1HuSuz0Fl0KxZ3IljqLt+9BB6bsSWhFNkJ0WDRZ9e1P77/Souyc9Onl+SHUK0gd5FQH/6iLDcb
8FCfKt8FY4USVyf7Evv39ohrv+iijJPGGqryzaVgQPTs3gzfxdFLZ/bdg3x3mgFmtAxcaSS+hwJA
e6lNcQy/Iky4OVY5B15Nehe9g6yv/v95oXYFt4+rozJBdBhHYHNf1QJ68uaoJSRcFtolAKFog/qA
c92T3VnRjSujM92UzLwwqo9kGXy5PBjwKHDwnQUC9PGMEBvCEBjzrO2c18CgHnhOCBCyx3o8Fg6I
jjprsa/JmiKyjYRG53cB5dQLj/V/ZotZB6xkguuqOt+65GL5mgiGDtj736Nt6UsgVBj9Z/12p+gl
pP/jbj08AVVbjqA6PDuoSpv7MBmk514aTYdd9/DYc/clX3dbRSOhsn3vkCj/8vE4TaDfdo1ZWsrQ
FfcGc22ZXuEFUFoBDZgjs0OX09nbrGzABXYawg9IYuLNBDn6wGxEK+02d/0nxMjxVHeB2iZvViNL
vYMKhrkC7s+I11Yvceq1obKKRlqYQrb91lQFbD6pB2KbZyMf+HJDjRr2VXfbK+gkG5q4oLo1+20z
PltRmrFM/D5TEe9pwul+Jv7iJIlOnoTCAeMXBEPB65uf0m3xd60NflQZAXQ81QEXAenyc0imUvde
TEW4XmY7264D6d1vhS78wuIoNWFcQdq+pM0qYd1BdAvDSuDUvfS03GKKUbaM05LvQ/PzgbVRZRIJ
B0PpBI6tIzztSbCu9JdqX0F18CuCgN+IeQUvRP+QDk+qkufhxLXms1sP4uWznZzQh+IRnQ1ucKEe
GlaZNJqlKRZaYS3co9OB69reJuT+4jHq3J9mzdahYrgtq0lDB7QvlTbx2A+vincfePq5tQTLte6U
SDpH3PSt6Nor0gmFy/iufibROhlxVLyXwI6RksH4KgyAh18zbzP9oNoRmLvnPBC+MgNn+qTeQ6fq
7FPsKxihxwF/HQoAY1sBKGuP5pjtRpRq7qBTY2Dr7ofiVu7iXvJ97E0TPFvVYRZ8darW/vpmgR+7
B6H0i8fFMXBNRPUyf7fqv0vbD+GFq8tM8L9uoDST+4aVQRu1Xa5pdh9efughMcDeqFWjsN7BV7Aw
ZcXdAze3pFDmxFkFeqYk3kadQcwunQelOP9h8hP6hjwj27RxZKJqxaMc3o3yGsuRMzns7fQ5dHbV
WQsmM0IIncStKZhm7jz3W/rRy6nLwgKApOcAHLxOk3llz2w8ggmCT7mObkLkchpywoOYTvGgU4Pd
ayefHoNY/QkAvAmln+i0XVn4HR6Wl9RwPWJiFllJKWzlS2xzejdhCxdhaPfdxZIUh0WsRkt97pzD
qxVxi1vet+6iFlf/C8jQNS/65FHlkVEaCXhcpCotlZe5WqccNS4Rl1rcpn4bhqCx7/le9oMp5IIx
CNi9816MozEN1cIcer8woenG9EmtRB21I5nGX1Qq6u1w+rUiOckfymhhlw2peDq4VpWwFALLX1PF
TVK7+Q/fog93OZXxOM5SPq0DsJimYVzvl0coRnpUNMhyCVDJdk2Pnn0iZkVrhMOQahRfyKHqmjQ9
lgXgN0u5z6umgPmhxhhTkFeq34qXCLPgSb3rAOzI4xk/eCOEBQOeHsAeOMA47bNQainZZcvQGFEO
AShjYHcWg/eoEE5muqb3TEQtrLa95LSAF/H/N5J1xxS2try0IZu4iiOd3ciy3W4ACjznsNNfd0g/
0wKp/FuzJgfjBBOF23NIC5MudgvK0vdXwcuadXjikgc9ZF7LCxF/U4YXJE1OrHl7yOeGQQzl9EZ3
KLZCz9LHpPR1GsO13Lk6Vx1u4TM8AXIrR2jO01kY1wrsnpasmIehdSz6d3McA7bsLy0erp9TuSdM
jAX9Tp3xRtVrRmeQB4e0B5vJ6OFj0khk+qxTpYtOphUnDXUU1Cu4Q/9LYNQUIXXnnV2s85cgNk5R
XWqsPnzEF2WoOHwkhlQEwuCRpSXyKSLBOPPIefkebjfahINLKU+3wCuMf+jNqAMExkN6h8ym2Fek
23DX2TJVKyXi/W1gFgKUJjMFRm4oH3pPyJFCsc/lSdoLeAsTgFJ7oDu7FjKxeQxlo59EUJotPUGp
5UGRqNFcAFWgUnPasZf4l/bd0fq2PWozwXC32vjEI30eYWQ2SyrMj1T+inyJjnu5dbgmy7sH0oKg
Usv3AIz3oChqSJyAs4ey27hg+SzKX8oxZo9qCHhhJieoJeyOuSUkewG7iVdRBqr/154GZKX3y6Xx
tDrARgd524sEm+pEAWdnU87onZmNzYEzZToUOP7GpWffeNO5fSJGIMHIGDEu2YUnhUL8OIHCm/Io
gDWx8SgARBG6r+8nBzpTkDFn18br/ZKPV3sfrIYwV2bH5bmACVvV8cfCTAypyF4kYuntL+jsuV9b
RTboPjaEFVKGEIsnFXgKFIwTVkMLsWLBYjpYKQ3plfKtcxbh9SWPYPq+1l31yf6ko5+GjLX85jq6
hKcz1tymauQDvKw48VhyVhsQru4cAr/jejpppzM70A20KjK/5ZWTnv4uzgIPCsJSZk3np8TDpXp3
bl7fBe75/Qa9+vZhZDI430lk7VNGfcT+pi8fxYB90PynfsCB4zclYagDhdTqgIjdZgDFmNmMPFPF
Mkz2EYDtmEp1YiiMQ4Mvg34gQxMHqIRqdM1KVf2vdG78dwUMERC9em4sjTxs9agFZdJm8w6ybi/6
yAOe9Nw7LoVkN01aNrW+yuajA+ehba4O6NLwSISO7z6luTxlBIUU1/GWVxhYZHDrdEYlJpFR5dYo
1XkfIpyQ9SJ07f0/QpLeJtvevIkcoq62887zf+iZJw13fAUeXor9Ii6xRm8HzN1PVmbNHDjGDLlw
PNhMP+qovSuGDi+RV0QUnBB3MSGkSrd2T0ESWubLCyvnXPKxsWRIjq6P+nhrfkRhGU+I7wXX0ULk
rKdyY+cxxZVqOhLlfGzJSKewPZN7T7nJ0wFiOM+Hx1fUM/7VrNGrVRq7igAjzcU2LrbBLibB1tyi
gKpcbrYGUkMpL0wSNF5sW74Kt+qKfTQezhPXHtp37HqiaznODZqx80ZTOHC30k5VrFWy7J66prXT
XGEtt5f6behUGZCQ9lUiBlVu3Lk9rBLqELbpWyvLahjwCfhWsWc2sdZ1dM9bAMJhc+cNlJqWuTYI
SKP7NShH+k3MRuY3hGBC00xG3gFM6zySqZ6AYOvRkzr12JJHVL4MOkXX0XZxUHFOl7RaegqYbWEn
cmnHH2d5WJ8R6umCfnS5NoLcrrXRqWyPYcy4FFk2/YdeNMktXGAZiEtgvTw9mvaWzOllOW+XjduK
yBPeGvmYGAHf1EFc3dDta1at2bXB9N3jiFf3gZzGcxwOZpRrhPcCjMChov2eKhz2nbQkNZij+1SD
ffgIyk96ygboj+A8T2QvX66APaqnD2SZ4RORxjYqKeuMrx42F8synBeX6vKMb4mrdXVXycLbWoFW
gVg7vbhzLQaMYUAnrGxzTRLWqRUCWv1WengM6Vs9pXQeCIIpEVfRpqTHp+/2HOU5ovI8hhnwzCHG
4yRvZzmZe3aN8EsNl5eb+2ZniDdZeXzCH4sMa57cHaM02TPE/eMROiRl4RCI+NJc2XFoETLZwLMq
0ZR3XNh6CvM7F9VE0JOpW/Gs8Ypozr9uN7ohXgS8IEFeL2vD2ULmGQD0Y1hWlmJOjHWtwEKlYSXB
5vQ3qz03bZDdzqN/u/Qqic6xG/x0f2xxIAOaEToWEnRDYeh1xVKavhOO6HIf4roRknQXXRyJQMQ8
dr5rPND7PWAVrAph7gXb6mvn08CGDLlaOJYFVgZZTuhUIQD7Wl1uM4SmY6E1A9DFcNGU5QopjHoL
VCHyg4kM4cZtff7hcFRuhS1M4J5dyA3sT3SYxLEJl3+EOnHeYoBhQqho1K1FQ7cbnc3wvR9OE291
MP+w/1PmiNT6mP9/xAoSXuKEW75TM3wGmhn2zQm2rIHN5eiYWQk4K4b98UB47KggNBlcKW3HrIeU
3cr4iDBvjlaEmzFaEWeODk6E4oYH2FQz1HByW7sxA6XSPrfJkzVFuRJhx8d3bV+KqMearhYx7YKt
Q4H3y/JW/PPehNyhXoGnb3RXKyKE2aECBt/RrZVUhuxrhijUlMDKbbzO6sjX4XdjurNo11eGoAl0
QeqxGVbd6YgCYRYJMyytFZ1YNaqli52K6w78UAFaUoY8qrD4WW5teywpiPqCpSBsxrCQAJDbeOv2
0XXNlLrDb951COeN3ZSyc76ZQKLyuO3zGMmuzerswHvDsulR3HZ7gRt+2tm1WiQS4kLQmhRYu8RD
kljBDQRzEfgqQjVrZJgglXMXQ7YZkkgK96OVr9dvjxqDbsGuk1yK33atp03OBayIfW2RXYkUlGsp
Nj9pQaEeqq++dSaZCmkTclvxkHaVFGkXKZQaNwPThGTs0E0Lq0L5zDZtInqR/PJAof83bOxq5i/2
jTU5hG0nwzcBjUt7mEpU//ieGsoqXqLKqdagSyiytIxvpHZ8h6oNOWA6MHSRlzLXC64fmRz6V8lk
lDMSKtOota/HUyF7angyRCTxra7JCzHLB81ECkIpI7yaXw3xhOQeNRQv8WOE2toI4VME03obijz3
smgS+q2iNP620Xkqhe5yh/5bJkFwxTgDKgW8TVcpOtMydREBLk7Xcpp68AZjlQiKaNlJTQH5gJp1
vZO9Fi5XAHPxyoiCGDdqKMWekAV5D2DEdjPXXCZK2ZA+9TiCY3LBO4hzLDkin9s6siBYFrap60tg
HqvB5ODbtqr6Q4QciQDZHiC1VrsDjnyo+wJ4aPW6DxXNLq7F+ryfzaxO49upxCRTGP7Q7F8r+FJk
vzfY+GWVfVjM4fjP2BLLeeAy6SM+Jy6VV2rp5sG193Dup/nyjljhesFKgu4pS2dgeA2xLocVCaRk
taQ4V4rCfK9mu35iwfzcgck3Vh2a9ibNIOn5n9IIqD8MSHgI9NYcCBnvVcUn4z+mxS3+BQWOJ4/B
o6TA+I6oaeOaGEGTviBPzWpoPnn7ykBmvIuYYtPsvrPyj+Rr6awtmoaDLeMsJXapRmSMUnKM0CxU
92fDETaHMaGk1u3cVDesaDZhpL//dAjMUcpkEIZSziK5zZMosr92CbXRzwJAjRhkZ4Y6fcWvlHDe
oLN9mhQqnMPBt3k4rR5Q1HAVH2IKOS52dU5Oayik2Ci2XRpCEoGvzFsm6RiKPjw4uGzhOc2fw6jK
9+qNK6Q2f6/IfXQ0wSPEJieul2/+wUYB/nkD6iSBf0uDZCAjeRc+jzFp0MTc7MXHRt36V2B449Ym
BRuW3v9Y+Z8epmsAcThUl7rqh5UtWLCsa8Zb18VLMkHYD6j6NkjYC/X40s/m9juAgO5QOy58xKrL
eqFUmsBuKBJfZXsnmvImfQp128FuX20rBAzBgIXz4sY2DumRBBU7XCAQaw4hSEB2tEqum0AqpMZ+
BI/+2LQWPxMh0HSBAQ04gJ+GK8hmUwuar3FixggdeeWHwO5V2kENRK2DJdOexfriP01EygVrMK38
kl7iw4pWDr+MIfQsJ/FVURgQGfliyrcXSIDT4k1UlM1D95KW94xxryxH5xI8cCmaW0vNBxU+Toi/
4UfvWIwlWxgIHHYQNbd3sMjVBIFiBzlj5pZO03kZAkYX+Kh6OpUahW/Sz868UaVDUx12WdXUmQDV
Q87PJfoU9dvGWBjapjo+hsFYShDJ2fq7x18ZguZVj1Hmv2N3iQqt693TAX/f81inHnyR3oUG6fjo
UrNiCsYcakfXDlItKnhoJQDz4vuKkr7HdOFiRjmZM751EIGHwq5I0c88K6omKXrJWG6E2puZ5YL/
FGrO4/LS8QWW5IeEFSwPbfYmxIcaqDTYs28O8hF9vz3Vqdx2vWrdWyxCdHRJ6vZnJx2PeoxEU2eH
85dGHhgWIjD56yKUlQvDXAgzz1pPtkolpQup8atFltf3DVjDMn8/vYf+foN5gNKcuLk0bEMRXd8x
8svWhlBFn9J09No05y2+vM+CGC+dOMUwGLkJZgCVTRaJbtiLQr1xKaqo83IiCeBxtCz/5lG7jVq0
Vba0+1K8xqoSHAv1JYn3lMIFeAfalldFjdn3e0FF7irctOzw+8ty6frNslT4r46LQMrybH31FGJo
8f01+RHCdwf0RKuPPYbVahkoh6y12oS9+NfXjKivfkHVxMGAa4gTgmkK7FuxVEM0EXVbFwy8xLm2
7IVWpB6ZBBOezcd0PKLNxCeBJgJKyDlXO69ezJ0bCflku17DUo7YPa3quj1TacJZcbnlDeIVFERC
sVbE7xgOPVgMCcUn8AUemosZ7jY21lcIucV7b8s7utke8vtEM7Hd+FhSFTzQNFyec5fpQmEtUOAE
RUgVjNwMeVOsWUrDbXmdfAKRNoeriQBGTCNJAujza1Pu53HoEsRkQ7y4mou+CXAPnhnfTg/5xunW
Kncn5e1ZxeXv6rYrDAScO0Vq/h18XsOZrkq+Ve24669hDHL001iU2AAKEKYpDE7NmjCobCxeJrAZ
dwGjlwPdwhYSv5cJDeV2Q5pwOzaSOyrQueEGWbxmj3YZUT5JGkAA9/N2wN0JxzquZRh9a070R6c8
lgAK610SUlXnvzYts1QAmMlqHsOjNnn1RiZDkwQcCGto7+rsI1QuCglO47G9XlY3hMBTYgUsiL44
5P3QpLfFnaTaurQVtFir7mR2QCbwrcD9sef9WjS9KCa6ESdNn15wyR8OaQazGxjEgOJPOV4+WtTz
DpXy004hdtHQdQgUgC6WhN1nZ6a0MvUXzJULC1wb+P63NlsugXc6bxFIR3uOVcBpUTRNJVsfARNR
mTxVikjjPlMMnZH7WioGT1dJAUMhZsydmr0YhsY6tv9IcKAP6KF81ukWYDhZnvGyXV9Pm/VcrfD5
HapynqhydJkjqlEPxL/5SA3ptg2T7Xet+aw5YpOljI0bJF3lXIRa10URe/XrkmXO/fkPGOinjXMx
5J3R+wb1CLZ+hm/1oEJPS+q2hCh1PpFBjvJPBS72RqTxyxjOOChDbGkCvbpSwz75M+byBedviVKD
ixQKb+FnRdpV6h0Qk79nTwB3N12+6Ej9cH59POifh2oei1tC5VktaiqHsqZV/QrhwH+3v6vzfdSI
fbXK0KHrRziVeYit6O+QfkoVoOtbYdi2TX57nPcG69U4UoJaSnDN37cdT65d4ZgKypRwsRkaHBIk
741sRizMDhIUE6jMcXxWoJo7aRljkJhS4b7egX5dpq8RVn3c4ZENqfgUQjizX2VDIZ9KGog+gD9i
IGp5v5y5YPXv6ymMyKBEEk+9sYourTlwInS5c8Sw66zFDfgkhcIzneqmu0xDm3/V/SCYbPw0wGoJ
aK1gPJl9zND1UOmAJENgW5UvcAjygOXy6aFU6ouLTxIN+Ki1ErNq9nwgBfsR84vOFTvDM1ag9IxG
cH6yLqGovdofOnVI2gQx2U+uamNdsRnhUDuvf7sTWT6jCrcLyB/PqQ/kheq/QsAFoh2uCf0ec4Jj
fVfyMOdqjf88PQktlsBcSxzHifXYsNOOhRe64v5ksRXMerRqJm9FDSZ4tyzOCfVhWjzJSlxPiMei
Qn29+eClvqwbew4r37SnQEC5iQGwKgfARf29yNJg+7sQ5xYI/jqdRQOiX2y/8HVTV2h+EuqorL6k
mmWsCU42HCzTVh7cTQslc3J/qMFcP+rSMqO8aozqdUdT8M54p5TzQDOuTiXUC12TSrbnTyI+qYmY
Tagh06oNnulegkHEIvMLmOgixnG/dYyrUOWe+52+HgU5jz/DhsXBAT5a9th5PbEkKQ8VQbr7wUH6
NbRELGNhdhlQITH8zyGjBrNA9/tyxtt2uEM67+HCOsI02hC9lbZTD2F4xzwHO2Q9ig5OrqR5cY2B
gyOWb5NYA7tByUXqTryrJLRg2E6zcP7FXNKi9yoanLkd6tPwan7kqDVFtS7+3FSahpSJxVDvw4DI
/8MZbyRGA2C2mEgNxU0X2Q8Y9JeXpr83mU2ydIDsAsxdKpP6dYuxmj/mrb+Tb4V3RlupwnIYf03d
7wy70iHY8bqU/pHV9kpBuVdNOHJ5hIG9w+uwwor/eaEd7cspbIcK+WcakVXxPuW/K1pDLyAVKHUS
SEGl9YC5MUIXxpoJ0zz+CwXec3gxFxmcoiOk1aNTn5LP6o0uoQU3GMleX65Zkru8QsMqpktPfkNv
fyuVL5D8XPA3MssLPFO60hyEz5C1yy4FJPzqpxnYCboxOZBtKb4RCug4lih38BYu1kjNzrf3jkx2
r7e8pFNPJEjP5TDaoYtwO9KeHkrztjgo8WsGRxPukOpNpSukTZ7NWxC6uQRtaJvQmD1SwPT28TLG
ZCxXWilejvNpux1F6pyu12VItZsc3ScHaMuCHagPyLQhGtOQ5+Odo5zy7J5jFBxfihWy52vTmcZr
5uL/PZ0dpCWSJU6NDH80N3jrfOoD1AS3b/gixkpFbsvbBUNnIEtjNgCIWUULiGTkec4WofY50hYt
nhG7b+NtEJHfGgrMIeyriPD81od/rckjDknG1mc0taHtlISFP+er23deZDm42PMdvDBsLaZKmQkx
e36ylf9zNCA2hReTAlYz4UwusSU0G8jErtMznlic15sKda0V91Fnlo9h/w3e8UYu8h2KSUMER9Ry
gv4o5WC68J4cnhDaBzhlLWGYl0yvhxk9yseSRfNskWfDhyXlYzFHgNlbrI/6KG46FHNFisnHN1be
IZs9YfFlLIw9HWpEyqkp2jeUsPj7aBIfzx+4cYGmE6MyeoMR11t59Gk3lqb31kSaQ9aQKGBNmihu
N7qkMqyvsVKSN/g0WUJ+90n7nNaw8EgviKlTF9e98CPpSB3VJs7qoKGw3uqq7hjfO3fxubsIQ09L
w+mcpscTSOa9+pGsy5tMFA/oZTdYkxUOGjpxnCwtmc1B5zxI16gIH+xizZHK2z/dE2BI6iqwqRi4
ZFzvpt3IJJ6F4zkxALCwrno43C11ILUssJ7JPXDu/jK7SZqS36iNVC1KAucFBVC9hcKcOz040YS3
VUtVeUJi5rInB70YHK4n1zv/ZbOdidAYixWRX1L5r7XRMsGPA7BpqzScgWS6avsQvmPMcQTdR/gj
I59iWMtdotBsbn6qsBMD8356J2GigRYRQUiaq4Na1cvXjkXFLLPpVvvZjeegghZF9fTTZn059yAo
MqmiFdhJto6EKzBGil1c2lWN8DcUQOV1WklDKdVnkidwYlM/0NlEgQ+zWqufLu4TRkaGail2RpS7
CTq+bfULVd8+Uk4ceC8wAfp8/w0wled7JcmEn4iN3FCXYb5bJIflgWUFtyVPk7R+Oq1BWBuBJyIM
pujxIx+k9Q+47qYDzsNeMtp5Iy2QmrfoWxTWJ+9eQwgDcUfCjc2R527+Gdr/ow+TJg7t1OhXhp4C
3GBYualaiUtP7lk+PBSBnGsvIbiBN9e44POOaRgkJYTTEGzwgthBuV507gcufvbWKEQU6yQQtM2j
FcLiSPchPotS6jElSIbmTHz7e+Wr+NFa+8d0hgVj+XTuvLyPgoY8jPnAjBtDLC1ODJ5opRBHQKN5
LiOgs/1Q7g5WaT6pDZRTjWadz3aRGLy+nEjTz7m3Wh2U9EIgZutH4f1SehOJZvhNxEZ147YNzbTk
0hFviL9r7zxqFSzk+0oAVTIXs8MqZGLTtv0q5OqyW+KHcNwVdQSIOOZh/TGiA3Zxt0NURcCl+N2w
vX7cFu3IMdoUjQRALvO/PWQjsru9kfsvkmFrYLK1dOHeo4IBHQxQbfej5jmVByBf/tlIVtXGad3q
8Z7mKM0rlbRWgyLiK37Wzwm+OUeaeT/uXhVM5gzFiNO73A5jPjqk69CJfakkD1E6RMAQTcwMHTrx
VaPF7VDG1+CqYsYKQqgojqk7q0vXv77KxGtUxCw0OXhBl2CVeWNQWuFITita+Eso0AngRo0ids81
1GjnDbyWF9gYcH7fuqFCKcU38vvvsfqxibOemwk4rfj6308SntpAzHu5FkT4XIyH2xQPJ5otw3To
7YQMs69XXyZSyLLH823FsThFZl19vW4msj80g88H3Yg6ifIDPxD0HjOjEdv9TLf9CqQhi+tGJcNj
8zckxnN2G/Xl1ZK8na6Y0ZxhLREXXhaC/a/Wzl3NiWFiHN0CuPHD6Vb825kL/Wta4uFDuvLTgrBy
gfApZ29IokkmPblhQIMNm2tsDyI7Z2HGqTDCTL6bN4bj8LRIrSxUn1qt+wo2zb9fsHB1Tv30x8r6
Ehbjzc0sOOOk5MrnwGYukGbh8m07/NENxX6NuXdc/mhPThcREZuM4wQ3JJghkDuxlAWFERfpqQRe
m6BCWamNG6UY0OZqAuAgenq3GAbnoOuUzHgGoPa9aBnKNb3qsU22x9aQYmpwbLxyo1Lc8vMXWw0b
dwDNvtcKfTOzDq3lqZy5CXULvYsIHDnphLRQuYXbgqf6MU/utS8qswlKLriudAyUVxMWYwBpBbe6
oBN+r2JJfAhlboKEcEYV8GUKgIkDV+vL28UVAX4ZfIZz8+Tn8ozI3GFA0te4z7uDCfUk3frfvhMz
sLxD9Y9fiYi1ZHuDs7fHjhk/eVk45MnA17XWLC8TFqXv9YqoKGhv+28PmCePxQOxKWyG0vV4bK90
59pmDl12RbORD+Bx2pMxHA7Lj9jvM6OhajPPfAHWxfubbGz1lj+ldkN/wFdRZn5hUkQlfaAcAY6B
WH1tQxGxxRD9k6lSZ2m4vpczrM/vYrp96C5BpWD91PFP8/aSGPCZoOHb/u18U8gpuuSdOQqUDzlg
KKV1YH4U7ACrSuBm1bNSfUWSqJfjq53LSOHan1s2dL9j+zxvUjYWKj0r2AvqpCWfW/VvhP8G8WVz
0rA8AHPysbDebT+3fOWqAvSDVUkr2Rg9j7usoGMMfLumbQ958X+DtC7548tcnjBrgBe1F1ZotHuY
NNdxRXQmFhujoIN4oi/hYWSslYsiT/vVnQqziVQjHEPLav/WnhXIj3ynBxNAsWi1Cj/ID2PXgcTO
JhyBEUVX8X9E+3v2JGV5w3iW/30LQ1C5OSLnG89sGJSPetP6SP1g1pGrgA4aRBE+tjavW1u1P4BM
7CNhBsFhRix4twz6fG0qrdbQwBfbTycMEAmlFawJ/8Ajc1MZRQhLEXbmKb5qDZA1kVt90IcfO3w9
4+kQPQifPAGUL7Em+tafdxgHkZxcLVrXHMy7bsxh2yHFS751V2LRu0k5Q2Um7yNbhQ4wj++jQXtQ
npolDp5wamZg5VmRr4+CWLDsQpt/12qkRghloM1tUt9ssKtduEJNtrm6HcT1lqaUVzLNdewzzLA7
SeHXjdduHBtnHWR9wRZkDb4VAzpaFXFJs/t9thnO8HmBSpl4tP9iqoIelnZP4/ppH0HM9lybEv6A
+SqPZMxXNzgOXzxG6ebdXyUNLbg7A9BAYyfVFuFM3ICYK2VzYvDriGorjjLmCXkMTTd/mbgdPAvK
mPFYK+t0EaIMvduZgHkawB5PolXvR22OKFsaYmTL2jhuaQ302VGBqKznDXPevaF8bzvBZwon+fwl
9XrThayPEellIbrBf6B6uNTXZoVzBzTE4xylxXsuho7/g04M+D3RgyN6bSIMzz+exrPC7aFnW4CG
nKri0Exyr/mIS1hImqYiXWGoZ+yIUR6qzFofR2RuiOUzMe7MlgQ1W0ZPORXlw/L8DbDg4qZNtKYP
DxUhZp40jA/jdYZxjND7E6NYaeWChQM2cxckVGLZrwAKsi2gaquECCF16VMHbbKjsmvDodu7BB9S
K+qvnYruIW9VUzjlr+RcP8JdcG4s3ylbVi7WsH7RX3rXMxwsn4PTOi6AQiRMZ80J6oxMrM4t3Olv
pSqVRf0htpAEX0igXjwhwQzUqqio1QIuK0vdxBC8ywwxXdxOTEJNhDxCSjq6Evu6tZN1nSi+mnd/
6hQdAqP+jziAseQrDGcte/GPhHnVGoMO6ABRUOwaA/Hm9S/PLknZBQ+eb6B0WdDmYtCJlR7UP1tv
1XfDYXQY04HO0y5vIqIdIbfRlsmudUffizUhcAylsdyv2WaRGHJcYXYjE3Xn8Sfjo1kSK2zFPj0W
ywmguF0nEbSsZb2nWu4+o5q/Kx0w1mT9o4uAzVrUd8oktiseLHigNiurCdpf23IWf49OS/4vNoL6
NEuMRvZuShf0MFE+bAdvHEuinjdhElm47XegUzUYYly8nkFpsfLzdU584UVWyhY33JSuiOZvQDxZ
6w8Fid2gyiaEb761fG7hSp2igCFg7nT2kGIL1WrxH+VzE96cdMsS2DN3RW5UxPnnte9Kqnqq+PjD
bj2HgVnYwm1DVwps3kkcwecflWiuTYcwIgK2qgtVIJpVdZLDhvx4HGOs9b7PqfVRQNDTjbvM1Ssj
aLmx5FP7CugqqyXFsCFhsSSIiyXrR/Jq69HybZK32EozCHHhDetpwSe6IRCqcVCRurL/Lhbx9bGZ
CHvYELq+RNQrR0+qtrrc3mH2RECzAkluXC8MDpzNFgpsEuGFYZHRE+IdrHek6tq93C/2QCmna03f
6Ae1cAalR06Qp/0cXwGAYNGpKzlhzlyFNnllmUPDb8A/j/0Djqcw4iJCiANnk5yryHFnqlUr3POh
il/N96K90F6oGfawuz2PiokMI8GAeHDOAhhv5pIaAPWm4owXXftluu1AXxrh6M6WptrCpGx8p3Ad
+udP810agqbDaBcPTFOLb4gMwABpsiR1TGIdGVhUeE6ayWu4MKHyFFsa3cw/jYE7xjIiLKtD2I1+
QzuWsuFfOr15WPVuQYDH4SKpKbIrk5ITjHcmi90UVsUUqExw28SN6HqalKoqbPK1Qp4sUGshnuLt
1nA4bLL/VjyqHlNH4pwrtjnj0c/OQVP30RlL1dnG3YyKQaoZC3uljAZbh6CLiXrOl9TJ4OKtmZag
8vK1EZpJweUJ9C1guh1HdSi5za8+j3eyopjhJDpaA9Yl5w+C9BDH5Xar0nihKM+jr/e2/kZRhly6
mvL1o+10HrapyokUTLIK4s3FOrn2yOpqtUNRWQJvKBR92wFYvYCzTPntIC1/7b3vF83ElXDdne/Q
2lQXp+qDAiCv/D1tj5GnRfud2ja+xqu19gSDRNLfH9StSFaaaRhOxj88f2iObicq9MQSylBxgw/U
oPib8yYVCVl8ChO0oQv2OwYs/oL42YMhlvNXBbYspSEeW0/VtrD/MeIBGE+hJ8xpndy/366UAKce
gbPZmC7pFPqy78pBMa2MXnthaCe7BG0LYMztUv5l1E08MOFCPIMijjqTH+Kp6fz+/UbKQf5TejK7
IgEONAEjNUC3q23AUPOR0bE6taysGo/l82J7J+EeemgRqHiaVS1Xomxpq3Eeuz82A38EHf8lX1Rk
JG8j5A7nBsXzkFoHgoHkR9sS8iggkVh/V2jyl/HH69q9uwI8kSQNjO2HSx7PM3PLA4Be4I3DMaz8
2GFr80itqc5zassygvDB230VaKzChizDGwfga0M8OMCJhnsegClDw7ux/CXNEJFEdN4fbtNWM7Uk
+LDAcQtzLC8A+u5ufV7qgPPf4oWEr+uaEtvlxZB0AUgVFDiDbFsQ3NwtdszWbQSLI4VUtiWsARzU
2UBaXt2rr4qyooTOqJLPXLJ1k1MrJf9poGvaMbNVI6qgZvMNUL19f+a40Sg8fFEshb8S07fbp5OS
h1Igx5UC7quxQxy0oGDZ0ngn4JvxNY4nbkqdLcBXZeocuSpvcstiiZqYNw4wcvPymeY052nrQB7M
vpH2Q9aAYKAytb4JILyuf4/qE7IVfYU8m2xUwzw5w4Ui5/A3DvkSv9FUxa8rzTTL67JbNA9nTDd5
1nbAElVhQ7k53CRcJSIISqx+nNBAsKJsLcmzAiew1ImIS3s6HU2AVMs3eDtcTEcWFfaO+4H/CG2Y
RLITAk1f/P8dcHkqg06zX9nnDdhkVAiKe00dpzBtSeagQ14kzJzGt0jIlGzZoHZiueDTt1lHvG6W
HtJE0FNPwwElrSGzIIwygZuHeBRpXosZcpsV1K9scqxDEzgZr8INx8/M/2J+hSFYE0seZtAPF516
WzlTHNBAoTrGn6vaHx7uaXbto6TNqusJ7MLFBSzo4cIYiIdMEZPlZlHQ6+jWlsOkEWc7gpf2IqcV
EoutEy+GoutH9QKC2pFvO12mSyJI91ebWwM34DcDTJ4oArnqFA9Mr7vEwqVLWHb1KE2aXK2UxMWQ
WjEEZ+EcH2lnHmkh0aI/9e0ZOFmuPKqo89TFt9jTIC1ZHflMabzSW1pm1LSBuyZezJbR6OMqbT81
5wXZzR1VJ8F2xVmKxcCD9c4WdoedbKyBx5W4u8xSmcNMUWBmLK8sIIwz37qNvBcw/2ICB22+3Zuv
H1ezeS6jqTecCYu+rbXjvih2Fw2qXMkUsvN2WmOgkJ1VWbwMQ4lipie05GPGeH7p53eAsaUlVsJK
F2puarkTHtiCACseZQmBd/dFAKJ5q0lwqM3ZR+Gu8XZaRUaOR1ix6/bc7+erA1VFfD/VUVse2bLH
uzKkrJtwTDPQY94PIozjsKNyBhkCs4K59ltAuQfoSUxRBxefFSx9UbjdPvPzCY7l9UqzcI/QzT/p
ybP6liMVZF1q0RIuMZaWOnRKAKv7mImIMZWwdY9bxh5olKeOtPiqsotPlRv+2bPJW1sg4vvBfdmC
kXRbRR64iwSu25II1XpJc0XjsllnWqliBHFFIEVQdMvDsH6cJljE8J1rfZt/530y+uYp+9LyWlOf
HvYyxOuHiprJRFzqqygZKTmD2CWYRx4/A9VkgnK89fqU+2VbqdHNM9pjVKLk4f9Y61AB8tz8dXln
KKbrfj7lZWSqr1WvdBwp7aLXG8ZYeroS7HWI/XTxQrzw8M6cI40HXiWf1gHoOtbCPqcR0XBDyi+O
6aUn9dLo/Vzpp38iNBV/Mj7BNJmF1ML0iqtM/ESkzbqNz6E8CG1vCpPyo6Fmumn0yiOJUFo7lPo0
zkDieJuOgILVAWcEXTd7rpzPR/tzpNDxpJz78bjZvqaxvyoWSlkMwC5EUPXpHwAM2330T2vo6bcU
12TlWGReCYQdA2kjF1ndju5SNtGGH2jOhAQa0Qz6sa29UsXxHdT4tUA3yNTcwbjxFDrE4aPiqK03
aQRL0qY75R1aCsEySFw3dEVMw2sDXklcgojxa7ihCVAZJhdCDXBUKeZ8Va20/Bw3vHfgm6zu/mDX
y85mpkwAQaIAkuj55NUDP/byDskmBXuWGyi4iXZgQ9CDN641pCmJmdHYXdLTbrUUCTlsS6QUikhB
8wNBLgkWzfTWcKEEN4+bS6SO7AA8G6mlIwLrVws3PtfrIxgsjwo1OtLIj5L4LyT15kMOj7MiQfSB
kXF4fJuunsvG65YzmTtRUx1bK8YHjeJYQpaCkmHCE2BGtIM5oqF1o4ffCJveyeEhddRrZAQtPlnC
Q0yY/2aE3BIAEuRmDrzlVi1MbGlNr0ebwEfsuvC8rRaDkV4rQ0v1FLTpjRcarGlUoCieiD5E6t58
fDoIrcSq6wDE6bQz1bNLhG6tl3vTsks9EWgpAae+SBpQP5NHF69kEFuW2XSQZxU7MY+Og3tVbs6+
ji4oxsFQr0WC+wU7iFWgZmKtcoevi/45GGAYtj2onLqK4XINRWfdpiT/9J7eWxpGQ/0sf3H1f7tW
uIYy22psZZPkjDA81BkI9oncw4LoBHXAj5/cmhTD+ZCte1KFhXIL+G/WuLxg82lYAMsvKlMZyW57
f3HlfHQr1bb61GG9Yc5PnWiROHAYDuURtF6IhLypggLAOVrFkmEL099z7jC4huYjQvnWQFZNKLNY
YxciYEDCXgOfM8Q7TA1dV44ooSQOY3ngH8VtG13hM+an3qg0SlBpTnrk0gWVaUbKkJL6J203YkNh
KOAHOOpAU+XYu2wfyYpdIDHdhRcYOsgcb+1ja1xW0P7XBZx5ips0XT0crP02h+KoxACEN2F+8taP
6+HCgZvPAjpPJs5Uu3g9GvkpxQFhMqFr9m2u0KL2fT/2sb/1RoaFaC8qUQXHSX1HzXkWnP73/5ET
9/5cp69rrreD0G9Z7fz4zR9YetS+8zpGt+Kp0gbsjpFdh9x3LU43A3cUqRsDIl+gLySZI6XpX+c1
LqyXFMJnd/FbfTgB2fyOzyoXvdFUz9R/xQ+Avt23F/enG1JlLqrCBUdrelGbyg+Yff39zw5Qx0dY
D+sWe5TGjf+ErcG/bjrC/aYljxWzuUID2IM1So42tx8uPdmRtu46vMB1mtDWg5KlXSaRApzmBjp3
/43Ahd2nB6mEupFNJElDQOzOi7lAT9L9WjecVIbnjsblAw+gpF0ws446f6aK7p1tLgE7UryLUzaP
XKCC/g/jjnECNkxHk0KlzIwqKUkl9VQ7OArytvW5bLH5HgPXcnEpslRr7FBKa+/qWhCXLy9yP9zq
KMbkNBbjwuqYWUp1AC76/pQac+oElqF5p7P5/Tqqbg06U7PThkXaBTAQpnDHnuE0FsveclhRHFOL
FFGSqZorb2zLXTCl4uc+ndxceQzXRqpdv4xFQ5saNgYG2jdebxiJrYU7F8792/xsUEpbbx+JaHoK
OpTkHXFQSo3WI0W4rADjL/5kjD92F1wXp/96txI8FMhVujN+9F/YB/Z9gsPnKiEQdxQd/lYgobR7
hqKQO/k1LRycOOs4Dh91XsrERmk2h1y6A+DofKEL6i3wdb81lvVIUuyX2px7tCa3YDu5zP+Jrgwl
UH7iqYfXfu87a+cGaLiyg/Y5WkwlJySfVyg4LYhJBjOZ8TaD4/7sYjFELhCz0UrBa85V0o5VdAWj
70EJVo0r2a/zV01KbcZe7sqzWsRKeB02hzOk4Y/WZ/pBMvM1kC797OcxFLeszQXv+WepOriuSxi9
biSQw2qPYSPVq7fRJts0UBledG2r3nx402bzwVS3Fz9WeL8crGTNMANQ+sOEtYhKi8yhKNB2JDxp
qgta8m1Yc5UaxO+vmc/qQO3LgxxyUYDk0B8QJ1XOrBoOcNCs+FbX32CkqH8QD6lTvy+/sx36DrVS
+EEtHaQkIaFpQN6X+T1p7iM2rFUPMCK8DYWmuJ+ZTC0wx5hfdIgF7Nh+HLUcnBDURjX/1uSji6AL
eA9UKAfzf12DrSdze+yK7OuiJXlwvf55TqPCUsrk+JwEIUCH9TgmYweze0qDOcQ9vtWFSIhmh/rR
UNU4UW6GtHMAnILzJWOaClukFgzF0wEm0D5UIQHkpqMHVsYoNt58aWse5G5fopcVY2F1lMCvUXtl
C5eSCKz4wiiWgmN05KTeJYs4meiX+ntXHfp1nQ88Ei32479V0fJu+ZL6AxH77mId8eYOio5zIqAH
Thwhie5g5w/+KYSRumBZlgZ94uqFgjNz85K+8ozqO0PUoQY8znaioVF+CKGV2JBXFM7H+8AGNuql
CJHVsIlm6gRBATO/g5VXVmHHIpFBORGQKg4VoEdqxVWA/JcdbaGShB9PkwX+eQmyfNQ015bucmaS
GiBwYBByEEnYt/5SYRd9y+aeAfxwVt+ivFjQCeRUKFxGVzmItUk0MArfHnadiYoab4Vs/beQskOH
OK52X/LpemHZplX4Kb7zzqLDErlak59kkhI+ouXhiqPQ5nHucdexHIit7QrZgQ8b7ZFKTjO1bDVX
rnONJr2l+WP0KKFwohn9gRc4RvZeSCiR4yKsbkjhrHltQzF2I9oBTuGUEt8/Ntb1p7f3w3AO7nCu
6jJcgSnTEuFXj5sYwo3futk+liypacN8FUJ3FTt30y+DGBcwrmBUmXiQmKXQPXy2/6mWHblYX3Tk
pKbA7uCqP0JLrWx17sKZIVGVNplA4iSu1vspKFq/adytouHNcGkkNdO4PVoIrM2302qnGhwpI9W4
uv2dLLZV1vnve8WKs8DnP+21h8rhj/hza24KE1ZK8ygwXf4+CslAUVzaYTFZ3ubFZ/dvi+enpVo4
is5aSeylk7wCv/6DdU+514UyN2lJAL8Io+MRSn1DUmh5nosRMMWDG88AtNT3iSwsrmdSi4WolWba
UJeOB04tsP4qBF2sPu04IyaRO4xUVQMYVFX5Q/sm1lQGvHIAo6IDczLazdWit6doUq5p5DEySYim
LkwXRiFTliHUrpMz+GOK/dNKnz2txA6CzAQQWbw71C2KpD7w0RI63BroBFth7XF7OrNRFSJzl2m4
CdZ+60WuImKJ4+8vBBOehAFhoFN8473lrP8lX11QmzvGwfMipOe2phktcglyHqSx5K/Tgo/iL36c
4QzVVPUQiW7ys0smIJun8s/auUbEpGYL8odA3+lPjlBtgjf6R9nvsuZ9uSMY9PZNmZAkMacGrhfe
pyt3f4NOgfv5fuFQBwVNJnOR/TQR1lXqy7AKlJAjbBEe/G0As5LbE+3FsPiRtXbvwspglvfRID7S
DIU8PDqWEmsdo0BK6xqdV2cjd5cNcA5jOXHvJtx3IvOFneDXCW6ZziDMpG5zrzXA7IJMuPxwG/jV
oaZ4qxzyHfCfdG6n7f4gDgNGKtJfxXijh6Flr6SlQgCFqc56PevNtbR/hPVpZQ+EPH8kPvD9ft3U
SY7v5U8ezE+k6nIuUPCa90EfYeBRxni99vDxN915/TZ/Np9pbT4hFU1wMZUJ5mgYk2n2EEZzBUMH
vfL4fJ6FxOXthfnlaVx4ya2zT+BWMD8qYBQkG4jJSF0Od03QrK2Kf5O//D+1qeMsfErvKY7Rl2Dw
yktLrX45q8UoE3R6LDZheFlbUDQJ9biURyDRyG9CljXojDSPu8cyjPcQLpg29cYuzICeX6CawPDn
im6qZib3BLa/xs2B2phZ9Cs5TeC6P6tjeeXlt1xp5vFhJ2AIQss1TJBUekS8G5j0ATKnFAmzmzws
cc6z3mEfoJr48Y8kpFGj2NBn9locEWeKXvp/9GHzD5BNID6Tovi9w5ZM3tb44rQEncPpJO4Ar0Qp
u4k911vYTMrLLbUOPeUTZ+b/NrhLxnmgW+5EcgYV51ZYFPwOe8d17jpznMMFUDbBBP6dY/3elI39
z5cPD3zbWO7KzVCoDZfeLWeHibtt8RiHmHeFCjy0JTadlshAROrehpvMJ20nK5FfrDa2pEoRgPvd
V0aOMMruX/uCpabCM3HyU9hUXAxHk2b9gEvm2F/3h40yW1qp0P+pFySmP0fnQ8YNSnVyKCfnhGz3
EAIQ+Q387TsoVHBaaPMRkv9J0d3eM8cMBtqREQQOShlFxkmejEiyNeY4pMMkt7E8UyINp/4+Cq/E
MgrwKOCTAAgxYw4hko2udffnSIBDaHMrBaQs1OXjFpDRL+O9Sx3maPsi1oae3VBnAk3PKBEQK3TD
CegOVZugJluZB4EaT9QecRfJ/n/NupmTa56fk7TuL86qN9716TU366uc2cmc4EIljXVa4Geh8EDl
Cbs4lAsb+/pvN06tg8CbmxFlFXs/k8r8faiWFauQCB7kjjsYV563m2/gGEjwqxf0sZ2Wc1NsqEH8
TBDuM/OsV+Kyp+TKyuoka3Oc3wahs7Q3ydCQ1Q0+GAPyXqvxrmFmXg/uuYNW43eJRCmi8WyFWQu7
iSzzMm19oLJlxKbzGgF3uFfz8k0Gn9KPBjAXrQHvj5PUFT3I40CTDWROAf13ULSMZGk9HLlF5FpE
UDps1IPpjv62c47t/psPgIELFNNLA82eVNYBguhqK3BVIZzQNXcHDz/5/QoJ6512aicBIoETUFN+
M1g67VqJoFeq56js1B5GvM9JFpIU10I1uiiyQ2950C+3mCpavCGxJI3WPYKOgOs3XQPCv/daWnm8
JSWtdj5EfeCHPCsq9abVtv4DtxWfgrsoMEI4gIajLHlTrcPA2M+BgpDyFuphqXwR+HeZFGxjFSgC
SpRGMR4mwSqOYbndERAfEobva2QiaINjW3+XKgsDb+0nznslO8zZpiccO8gkiuutuGJ48oTfIgA+
OSjt6dDBp7fmFzCFIq55dKrNdo7ZTpH8UENCr5EpxOc6Z1X4T6HXEGDL5WY1tHRT1to5ZI/nnDvA
UjwgGN0GWBxQ29JVQtDzgq2xBVYgfijQeAXw4bEccteFp+52MKZRKHlkKG0pZ9UprWxKG40E4QTY
SN8CmwYSmUr6B2A4DieZK4S9gDrr6NguTuTMuUwI8dP0H8B7tic8aReqDAHCPCaNQ0RZKq6TlEkv
Yzro/d8uyDEmuRPhYx8YbgA1PGOzvXUGcvavaeZtirTye9mD36F6/lfKGjtSx1gk80DhzyQMZwUs
zSjmXPtAyG7uM7KliwIPSQ4Q+Us/dKUwaQhB04tPUgghZx5tR5/T7G4yrqXRkhivEzEYtl9KXtFL
zNWem1vWnRM+f32BM8YN4/OX/C/uFLAkw8hbe9I+2les8iK0x6X6IC6Smn5V3ZZXSWuerg3P7lRn
f61D7RNARZ4lKbflvWv0QsgdJ9TYqzewDYpa6IT2IfySbTWv7X1L+rOahYQdEXTExJv5DLOOHk4v
J1f/YsYLGwwQasBwPPVSZi6viHNGMRwG6vHltEfu4nBgFKsev4i061wnIsqLCa+SZFLvz/rTs1SO
CckY9Qg5x3RBqq5odgnMGxgoG6ryqISql+MhEI2qSam3WXLiSOUsIF38Bz+KMLtWXatfl7yRVMNr
zMpsn70n2Oj+9kGA7+LXU7mXzntK4VwIujX08rRzQwrH4uHugGGP3KTM3gZu+Xu6J2J+cbEzt6PU
Nv5hm2Zw0hXdZJSBmwbKkgRUZXXzfQRQyKSa61S1bibaQKr10A/8UlAla94iicD8Nlkbzd1UBdDj
2PVe82HUUl2VQ5FJQgclndqblE4ZzwUPn8TWw/fsmehyqIii0wjdUUQS3e9R5UpYO9WcumzOe8rv
prtneptUt6Oli6q70DLGcIBgPKb+Ce1cL0mbgu2oBj2K5q94KLiv6Nbw9RiA39QWjsdcaAOb+shl
XccZP23UhiCoCGeFH8IxCa4FC7FjUyR7kCQ/c/trwSdGMscMpka7SzBG2mTXTj2qtZWFU2bxApzT
uFWxSe5MtdGR4NPD5hJfAsb2NTT9nVcPrd7l3P1cRJb56zHe60oXx9NIcGA6auxbb+pY9nCf47Qb
2ce8vgpPWNr0lnsO85/Gh7iNgiEuH4cTmSG3+S/vKGDVW3gyBzW6ThiNT8tbbdAHWo4DYMan+dQy
Kd4QphrqRhVYJ66o641WFzuSPEMVDmMkBOjFeIOCfacrr1vvP33xVJFxJJYNndCn5XUckhvQ/3Fn
+V9exEPk/Aks7Ca+I6t1720r1JfsW8ag2sqM/hzVFgZCNCGDrcIPHOIk+4lvYfl+rdMSjaU4Bgis
N2BFbJ0yaGvorXqXyeN4F/5Ir/J09mNDnWZtb64Onl5wu4Dju9U6gYnP7e3WmWiVxqCjWkabJLBt
zxwuSyOhiAZty9zehGzaIXFktBalP3AzbCCjnwYSeLtv4lJ9iLeuhgQzHvX0iHCSLF+kVnGr6hxU
3QQ3Naul+3NgWzb+U/s7hTFXQCOVK3P6JDGVftquXtw+C4MMJuEnaFxXWCJba5MvY8STRAygcUZ9
8WzKnynM7JAqX2jREmvDN0Bn5FNH6SxADzcEWPNi3KR9eLcpOY8/IzIsRLc6AP6NZvhT3jbK67w7
VRuhj2YZZVxZ4jxSpJD1SoKO8kk1EDD/lLVy+1Mv5lAK+YlmknNwXSIvrSioQdcOECKdBhq0tjff
qrkyYCOVqtrZYkHsoMUgemtvgob6bvMbFZqngeGVT2rRIOqoUzGR8WAL647+GlyL6vl+tcHYwwMn
1Wb58vfcoxfVFi7JywT8oRC9p2g7SSTq4jZP2TkMGH1Y8Z9wUr9Rr5GabwT9H+O9Az10+YMKIHox
ki/6fQDQ3Xni3/oQoBlYoFqGgE3ckvDlVxivFnLibG1WyQGJ428rgk4a+ilnU2eLCp2AuEbnPrxU
JARpjigFyTYtnxuEXPj+gBD8VsvOiPe627l1L9/zAyXsfABQ+7hvT3riuogNtqTw9epewap05kqi
EGKsSo5K85NXNNHd1Jy/mGIKUwIAYPZewRGNToCYxYKX9bkPDFoTgQ/HMflwKE7WZ91EUxYYPYKG
eRumlR5fWfdpnGWKtgZjcQ+jjlCTYxPhVdnagsj6+dBQK+7Vh9vNGAWE5wL80uTg3zaiOb2xQ9up
Q0orliWsqJnDybDnG4tPSYu6pGPA5W4HW0kks4F32tYJYNnqlvrIkFkcOV5yluNqYuMEWRaqmzeN
V7pekKnhd2iF+EC3QVUdDHCm4ebrdYSi+jfWtsvbK8RIibQo9UsH7R4qS2wsNBPue7+9JqD2Wvga
mS7loUExq7h/clJg+couXwvDMm7etqmNm71sRMFHC8h2flJXcLpAaUUC/x3Y7S4olLEt7M23/Bax
0nvuH5o4iFW470aD3X/babCsqnEn0tyAAJg93ZiOAhjiliPVvUeAxbRNgM48QsKe4n1zfdkhHJSY
VJ4mKsCNTJ4NyGlPlKyRVpGlKftY6B1bgf8pZUqRGKdQdjqdyvM2zA9tJSyXOSm3xyfqaTuLtyX0
X1JlYxp1OVz51rmuoOeirl1p7LX2yKUCzLfILLup2HzJXS8fEN2UthCu419IyhCM0FtF+h0qvwAL
aerPVIgP85wd9iBdgH9ksKLrn4qwRpvtBZiGfWPwp3pOkmPTOZFYllaYrGqaPFFSbbiZDzBw8pma
zTBQnZbsCdmk4MlAZw/Nt9fWvDnWbdwoVhyKPHWXLQY7o0rstHDBzDmiZw0kx0jcpqNwWBIQiHK0
wIe2oYULvfYfiEurzUy4090Rt+XT3EJ+eRGXgTEcwpKxOYdMND9KOO6tqLq1S2nvzLk+7g5TUwzK
3Sh01LDKlm4NGZXqkQxcH8YOeKRlCWlTPs4j8e1DmhBFFrv0KX//0OvLli9ACGS9Z4DWASEWPnhG
GYWgi4UJNz/ouKaYUCC2Ab6NgoUrm+vV+MSY4kyRuwAixwSS3ybU8djjtJhbF5crw1PJM5yLmOR4
iV5Sc5Q0u83tD5zQo7oKf02yR9gd+P46IXtu8Hb//iIHfVd3I5EF5bFFYeYkhi9yZDlrwoJAXKH0
FS3pfE+8aXOiHUrBH3x1WtMqkEHTB2C60vQNXdY6FWo0pO8AXRxR2C7VZKR3s8it6tERf1TCw6ow
cIR+B/7SkT8Kyo7roxUTPIPWfiYQcOmck/RvyEnRrvs7YgdnlkZHRLm+XERMvpk/mUAaCKJIrVRk
Rs079ISZD8ov+8ImNtDPsdiznvW6UjWq5Adst997b2lK79NUE0KY641ZNl/NE3Ek8tP3wslh7NJ+
MobBjL+g1vdENTydY6mxm2EjPjeOFl/ChoYCAv7Q6Ftn5Ou4NMhp1p3az+CfmOePinwBeIMT5dst
Jr0pJlbCJI7oL9v8kVwvHrlXruhQ9PtRlUo5/E1KSZpm95WyUMBNH0c19i2sMJ1JYs5J/Umt9eT3
UB2OSdyffX5nb+yhLWKC/yjW71nDezgN+4TSyLuzgqdzFt3jlTaqMPEHu6cwo2x0tbo2zivGoCkz
tfhqTskaNVISgaSjpJD1V7+LZNKlK52Kdem8RroQ4W4aflFtEfXfFJv3irnpehXHgjLhOIdI2t7s
ChUGYJlC7+eHpGtf4+2eljtjjcfJ9fOzSnYApSYbO8B54z/cS/X+yKzlk2S6NJmEggyBjxHpIzPH
V0yLEXJ1LEdthm9E65r0Fc6WSKJz/j7/Jo8iCDVevQa5v1UkKjt62W6f9P5SZjzsI2eo8vMAkkFM
Cp2eSjgOicVUS36iJFDQe7ErnMc67ytqE/qu741gIAASV/NfKhlqYCKp7Q/vEz4Lzcns2nKiczHN
hkSbPdiRshluGlLpoleX9qfXzZdJcwrYbBU8/Ob8M/idOQjU8lL2s1exD4xBZ5bdsN4Ik6HJ+67C
aMx6TIWCKgrvZ+HFWNUqmhXRqkjFpeMP4s539c4Mb0kQHXKMCOv/OPz4iKE5IcXS/ZrFQVvWVQT+
D7H1msml9ewgMXoeYmq7h2zgq/fEXCCZNIjYQFJ6KNjNEfupGDmKtLEmsW9fABNkAXxFdGlhddvH
LDYhAlT5hM686JvSThzP0rhC5O7p/514gmlk7trWbaG05bPtswCMDVaqm61ZN17qcfad/c8xh8Jw
yUXea342nYyAjyOSgcY2A+4xQLjU562iVXVA8tuqdY+KPEk+e1oycXoOUmKrJd9IdfrGdqWbvlKn
j6S14/E8BDaJjdRDo778GUgXM4+qc5Ruf0T3lcW/NCd9Ur1yIUnXNZqkSEaO8W9YBBep3DF6Mj+v
R9c5nBrzp515IJlBxwmfSl8xa21Am55DDCWNMpftCQiI45/JHJYxgdSS65Bu/RfIBUxGDXecZFzX
X2jM4SbqG5WFY7RL/s0hbqPpWFtxaz8flXc5l1NAxiLr3eiD57LVuLtcul7YcILDGajdLwfF5M7g
BqMs450oHtPzkLzSxoc5iZ7KWKfn0V7lMOCE54QuehfS5RxGiKide7Ih+nwbz1tohHb+p2FfapK1
Vj6Z7N0DD3/iXJ54ux1M5n64Pe3iOjnmm79JvN0k2lYw2ZIKW7W/MKFkmxYT7+fF0on2yH0fy0wo
+3C1ROHK5hsLmxXTdIskTqFsyqngxPCSdWU3Z/JHCvSjBn6oXnpSeCOasCFjoJHCrJuDqo+gq856
QfYqpYqhhKBkrskyF4WzpGjipLrtH+feKZmyV0c6kD/fTgRYqxCvv+WQGkAf29D7uydtd3SS0vwc
HmsVqqThGteC1tFPtpZlMdhNUI57XbD1u+e4SDUa7MvTH9TbLmGeGFjboBAjaX+U+/3ukpCldT7a
oTltOImFuOSicK8PWH9DxszQjZXUwKONF+P2p+PedtdZM+iwjDiL620PDqCg05Ch/SAwNwwUyebM
Nqmxjao3YYGDjs+AogY6jUD8xP8lUDxQm/NivMvrXihKZZRFwjSRWDUwhnmJMEFB57n+44x7vsm6
VytKU3QLzFw2xl6VDWpjwZFLHCXZU9aK+kYolD2Gc4xKx4lSW2hWzeIIMZMFqpbUTlYTl4MG95o6
DWoQocY+qyE+5FuIMWPERMuS9IJo1KmjZtuY7LQ4kxhb5A+0uAyU6Re0zM1Bwptq8nraY9Dw6BbA
NOAYETqy8X1SjIDtX6ocL9FRF0GxKgUbgiB+YdSxIxFaI9eoE1vmfRKRhzsoxHOTGq6IG8I7QpNU
VqV67OaalI0OV8L6lHfutvc98Ag3fdZhOoydho9zPZObDpq33VyoNPDDHBasLsu6WFL91tdY5ECn
A65mI7N74T6NIWVQYPH1y4M/barNbcuJT9FccEDueZEoQdiVFw7TpCVbmgCn1sPjm1X/kH5ZRCdr
xweU3+QgXCWmN7k9BMWTbJzroWIBCK1u4fdCjif0fusgZWHWFeNb3ICerIJxXa8uyq94n3ZK11r9
6kO7zTbsz79Fr/TT/oQteK79QLCAecee2fFepPB8wS5/nVoOv+VPtYqoM/yugkywa5KdSOQxT2je
ePvYEVbjqh3lqLVyqDqtHpNcE6KJFGkP/s720QV+oI5FKbsB9ZcLhAO/9uPTHyqotybtB6a0aTrJ
ktfVFaF4Ht4/ijLRG4i3c+RakaV49Znj/z+YziCEqfuNBb+ebfyv2YWM+JTqi080Ppp2YoQugX4R
oPFtEXPbYEcte4+qLa2/4t4NvjH+RZz+OPPvVYr+P1Kqjiu1GMqgoippFBANwuchVVfNd6D48Peb
NSSdfkhH9C5pAzpb+JOKpZ4AucStRlzcAgiSCkI1ZSb4h17/g3vMJd8+SK/mYEKei3HGAuVWWjLr
/H+1p0qcA4PfYopAudl7QGA3iC+U77HiTNwu8tdMU8HHKdARlrjC/Gx1q0x9LkjCsFhlcLLORM2L
rW9iQG88YuBvwC/jT6ThQKQUlEPpfT7HDI5V1+je0fPLPl815rYQE98jlCaGD5cGYqyLlmMgja+H
9NNKvF4rOWOxj2SuByqX2PFB5GBp9HuAB370T1cHtSM0Hoekc/l46pA3i3asbDMpoujgMglGiATY
/6wXZGZOfCvdHQFSP4jQWdadvRRfyrrhXuL8QCTMY32e13aks93cDWudaLex0SvHzGUGPVUmKNYz
saTJ+7jM5PvOyHdagUWkHB7neRWlxDGjBGyIP1rTCCUla3Xws7wYPCoRXVUgoNT536eNkVaquOBO
/6sMBS3Q3vH2LjZbpjv9nCPyNOCKCEkh3y0tqS32T4sL02OqamMWPhKmkDYKmNSLLVC3wArmeKKr
BJ4KaU6MxpVgXypBYEQypmIX+WIr36OlmY3yUuX56W+H400nJnTh4Oe9ziTUdDpKjny9oBEI2nUa
5wo4Tx8H/iYYu8AMbTGR4Imb8gwVWds3B/FG9eT3zx7uT4KezL/LflwXX62PsjDGFk069aAbASb4
mLFXCSYPJahvwk01PBn92m7datsUnqzLchmouW1/Wf7GJcRsXEW7KLGnQS91/2qw0KFCb0uGCGAE
1OTImNQdWyo/MoZXeZshOdQMbAe4rmNJyKIE76Q81DulyBJvaOw0bmBsYB0rVu2qNkWvtcgg1Ih1
mkgOFQOhJuukg0XOD8yREJ8FA+OAlTm385lcGa1uappPRV9GHSDDC8/UpaXHgDrBV/38mOkbB1/S
sQx7zZoLP6DUGDU8qD9LTgMZrHnoFPYlCXhDdOfKIWcD15Kq0P/P99egEy71aIVJPigX0k6RQWBG
ck8q3VQTLkcC9wmYNQ+gwhpvlBXsnVBsn460AL30EIGTIyHDorUbi5XglmjYufzpnUXjxjP8BwEj
Mio3ME9jjmSAlaCry4JNYlsymSti2ODoSE9cyTNwiyzmDR+eD8OOJ11RLiLYBjhJOV6a3kebb4cZ
x0eQ53J5WxB5u0AYIaH5JqnW6pnUmVk+xeAXuWWRI8QWyFWKXrwMCPcn5JnXB133BVuFu+oIyC6y
ZX1kLaEmRv2o2dEyMeMEjVVi64nudCVOj+2+oh3srxXdLfGLa3iZDM4DLFhTkOREW7ca8JhvTWHT
WjvUj4AN5gCSY0FeLWGsRzO4WC3zvvANOSfqSS261k7G8zx4v1G+siEW1RUudGAxzWX0qcnuyPie
wLlWUM2nejiI2OYeYw4lk+G9NgNUDLhcBHDzvBgIsd22Xslr3sutcuqDbcMMygTXXQ9C8gQqohCI
fw3WCsBwQEmR/1QZ72CplGy6L18QGcMMPYDzgBO+k89nHENbpmMTKppB/IjQXVjwYPyj10VHwKZw
aCGUlEtZ5B1ksBjBjmITxbzh5XkGtjdAOhY7mleQN8PUHDS8YzPIb/25WxNU90DsJ/FguDI6lTSa
K595aXUccbIorF/Nn4yy4hikfVj0woZSj16qxftVhdnI9CVFgrNv2s7Sx7+AHvGRCzKDAGCZ36eo
nEy15aROGGLUn98zQWexgr5B+0545NQxbWk/zvq0+i91h2zQ9YFN+Ws0HpStaRKtu0rXvUTtQN+i
NArtL7JU02XVTYutv1N9o588CLJpRegeFW1UDtc+SiUIBtA7H+TY2Z2nR9Hhbno8Yy7biVq8fU+m
iK+pkb6o4lMK22ORRZkb4pVG6UnbUW5yJXYwgeHeuPl437AeTBF9XG/XOU1Tgh5+7W68J3jjEtiJ
V5Wz9v9HajG+CHiJCeMBb+RBBZBU3etUXHm+tMBkFSOXsQCpyztRB2OW27wPYzrAhJM2QwM7M3ST
0ReeejpFd57JzBt4dxi9P+eulUTSgxcYNOhBHDBH6hdXP1+iCbXaAgNq9ht37TIF8xP8PCm5n7ym
l/ZmTZXOcgzY89mPs7VgWbLMNBuSNOeaUpkpiLsTVbYKAZcXu7fy8fOf4RrVBFlUll06WKKTrpGi
pZX7bcqf4gHjNfGVSiesJuuf9g2unVqp4xCLC8hCmhzodVQ+HcbcJZgaRF68KtLR8venP6Dc+vu+
fbVwBqY0WGhmt6teR3064b3NmTAsgZFOvfC1afgct/Y6RNXK1Z4TH02GY0uUOD4PyOAzI7IxQCKZ
ioyh9RLXK24hq4SZ8+DtGM7hfBj0BAw9JCrL8r6xr5YSwNBJ4UdCSjA5oAuezXoqIufoJ+x6t+jl
/YDxygBuBrOopXLNcucxz5G5ZlTaTWK7FWi1PlRTGfgEXsmUQ1dCBI6GNSYA4fFV6kT85YC570/x
jH6lX0TDFz9p1mfzTnA/cxiv3Xdq4DnQhESQ6o+c1vwEiTkZNqHfQu5sSQD5UI6172ppkGrWZXVk
sB1y5rNpa19S3FhCHwrPmwkcgMr0x0+J5bTRQNyvBrBTeiHj/fUivGtsmASNzGDiVgQKYUBdaiiX
kNuSacfE9lEl48cR29Izqvunmodq/NYAui3KyOyPqzyQ7snqzf5VzxoKMUT6eQE15nYKrxeBXEWX
BEqIl62bHn8iZoynChaZZZpYISj95rsPabR6mjGVdYGOL4SDB/BIQ+wIk3pf8HA7UCBpcR84pZbs
0+ZjS+FH2eqL2NGMy3uxa+3kjjMA++QtGH5ZI4k/GuuDGj+m1lN1hkW59V/dMdxUUaENsQL9ia2d
pJvxZd+INJSVnvknW8APpAMsPchWgtZUxIJ72W6Ty5tIGVmAtPonqSgieZl5YdBTD2GbGCXA+GTS
hiL6e4WTlJJm6sjZblaa6A+5TIK3AstYOoUPzegc3epQh6GtQWOQ29IG+icgK109f0SpP8XcDZZ5
tfiLblwZgE+0XiV1bMphvK0pNYeC+xozezfhol2iHgt+RYueQMabrtrxOQl0Fl9j+hLXbf5iemYE
0snWKgG+O5C/3ifFcvHisG7YFRilesVh4ijKgtmJTNpXE+PF8TXBZ70mk0rZmqYd04l5qJaqXGmi
SNO6iNk5Pc2ihoPadGd8PspPzj8KGB0i56BAmJusfy71nN4Lhk5Yslq3OMfzBBlZw3b3wOMnmdwG
l3frCqloEF5UqZh6W+w6rGl/MVcoC0WiqeDhOLA3yl19wzPuyyV3ZGT4PPQlF0+pU/RxQ+FIO/lD
9XItxYAV6HD9QHDCN4cSIFSzYYmG2CiOtU13SM+XOBq+tG8FrIh9WCwoDXruntKrhNzNQch0d8YT
t7VAxdE9YC5+kS39lCslNi1KCC7sY0kQVExvPdS/PBdbjxoxvJsmFpwTHFO9G22pIUKAsRGNfVMN
jNu13I4xjpElfMX3cBSX1tnTAH1GXGuebnHK/+YyvLO9jVGmmHmcCaXrDy6hdaIZWRN0DEaljNGC
wugmNSwYR/9ZNe7WgJM0q53dXShd0lq0c+Ft+XkBzLN1cBiJAWKEu1AMF+bEfmlmhvo1pIiSEgJE
kgVIkUGUFpbes0JDiTUAZP+v+MCJX9Kj4g9UPs4DCrPhtA29TPMVIKX/Qh3Js4iMm/ixbXWGpP5x
FwtDi4IYMHfXVQdD7nib2rJc4ujhY8RRBscp4+8aZoQk9ggA90YWDmw6rQzBukM6V/IJ82Hj2+Ji
FQDxFoCTxnYimQH7db5OxNs7qtDTgu52XW9tA4zOPWHqtSHeq1XmAAW41UUQNCclJ+iHETJXj02L
hqtSZYw4T87Q+5x8F16sCILCpGaVoqQqIMYZ1gsaign5MRCy/dlV6H2oSmDxd6BSZrWKIVUWGag8
74RGtdmZzgFZS1D2zTK1DSKjkmCuhjAppIN2kRitL+ocpRMgByEkx/YOhpQNjay2z5JTz7/eXyVr
s86vjSSQAlKFUK352VV2m92E8KWIoEhmE2y5IRBkS3bkP7Hxs/d0bQA1cMRTgXhotPIVQyIFE3Mj
+glndSXK9DeVHEzcNkYdLV+Mm3+OsuKXOrbTy4MC3qoVqas+/zz9vmot6lwDVY4n43vr08bD7CGI
OBvwwcExv9/EsV5nt1TuqTk8r9YkOUFSQA+xkuStqrnsNef5xcSh8e8USsGFkhskugmli0gjlXPF
IJtE3RdFM9AwtsVL0izgB3aA2OM3ZZKtVdTL1gzdW7RGtX6z4XSflx+/jKl+9UMXhjf6t5tW/pZV
C1usFcnJYldCTqhT+0thOGOdaKaG1itnESNQRoJ2S5X9HdHrSehBzQNm2Y1wJEG9qqLYOsU3ah7e
azi2OwrBebZe4FxVpYL/uvYYSlxFhBm1lombDOAN9Wj8pB1ymszOvwseexNDczt78R9gEw6SmZyU
4DcyHzs1Udq3dmS5dQ0aMRdCPAHn512c4CCqza1Jor4V23NoWN0n3NlkKksTj0SsszG2Nwss6xA2
28Fq6ESqxFh9YaKOGr0/NsggmJXm6gfq6ykRQa6DqhIIEM3RDqMkMD7YiNiKyq8p+ipeBJ0ycV01
0uPWMMlwGmv6TWgIMptFJP8dVdix/VvKHSmyE6ojg/A/UK3X3XaHP076ufdLVoOtiRprZ0r+n+BY
Cbpdcq8UXIHXOcC+of5spQ7TauCHZr/knUnIDNG/FZQRIYkWebfFNDRPMXcnaV4GG7HDy3YESb4y
4dLlqbY0lebbC7YNo3l7s87gqxq7I0uy5b0JDM4wk086P5GY3D/UAa/dOiVyy6qQgs/gYiVmYGWl
nbKBOWNrI0fxsUvU34M/9Z4RgwRmC/yQMmukvjp84xw/X/ONAnGOC3YPT0pCXXImeteDEV0EPMyH
q4VfgR7wJsbZfIp6h/GZpxg5XIfLkzBlxDEU4u5hdJpFuSZEKTydjmbDrGqFrZYpybKkIq6h0Sz4
belSqu3ZevNGs6dRsT5oPKNeK3bpxzbkQ+ZuT0Ewks6SVkRZ1YXP8ECMtfxjDZB+mwc30+KIk9Ay
cEcWXHtiq2iARr9xXRXS+SmC3Cou1D2TVjEgBXrvYqj1qoF8aVYKbatYbC5Er7xJw4YPWywoHb+F
7dhV4qiuvjxgl+SVfqAWyhS1C9MZ9XTlzP/8wzxf9C1UyLtYmJlQdEq8KDdrjUfE335iIJWOxGdn
7g4M9WdeYnBnDedrvKRA+YDRL2VwuQNlCMZgtNgSRGHsK1DJ+5LuCl9NPI7LDtXjbj2q0tqQez6h
lLFxhYMkKfmStnpE4WiSQsdU0430GyyHUou1d69oaH3BqvFAuxnd8GSKXJ/L4zbii0eoNv/bhFNc
I3wtCOgh1BbWtN4SC794MV1rGmrVYzNeqeQxDBVJfhB8zNpyzqYludTUNysSnUNmbQDdQiwgQU20
0AxpVuAw9dL7+nPHFcnmhIBNf+x3afk3Xq/8xrtpAsHnMjYa7Bw5KWg617XPKQKmwF3/fSIwrTDu
t7bjx4N+U4s6leYT3QabF1AjSO04Ng6/LmJ1pMU5pPeTavd0/IiusZAz3XdShLN6SZApM8tO4cGQ
ss9Z+AG8hWiUrvVU+GGyf/RzYNRubfMcvh6mb0Fa3lUth0gLtvwr30xHvPzD1Er4Tyktihip4pzV
pensFgW1dJt8bQPWKyqu+5M1jhwxRtsmFT7/FrTYEnGJxYRBdbjRRkAFPArNbuUq4KukDHyJMWY+
LsXfRfWqXxHYFWwux+Za6Ojdj1rGQhOS6x+fDxivGRnCzbzVTLVmOCQtKiOVS/3HzUD8Pyc3evw2
3Rsrvj2imP5CA8jgX6GihYseShuNI7DeOk9g5UXzXjf2/kt8llMiDAZTHsC68SFrAr5UHL+py3ei
DP2wohFrevA8eQd4kxMog08j3kDyTOKPkfnV9LHxHuomSMfNO+07nrUFNDmaYiUxAZXZE6V0Zfxr
IStK7AcAj+qfY4ZzOqx4Kdzbm2U1hcYRW4NLsgEfQZXgGdkVsNfrAi3zJrqds6iUTDMfu7Iib+BV
HK1DT+R81WcoBdbCguzXHEl+y17FDkHi+7Rr1/6cI/sKt6qmzzCrZWYAG3njqiLl03/Wco7vai+/
wsdx0caAXcSnAGRG/g1cH/5B0kbykCUMx58cyWTX3QuIIlIh9Dg/VoDor7Vf3bE6vaslLDvogzrZ
cZ8ECo+Pk+G8XocJ9ek99pZOOc/hc+ibk4N96OF7ValFupPnD+8cGCQ1OGG5tPoNqnTO5bFsPsyz
XEoGrHqakyszCKWh0NxIgAeXRn6NPPB+V5AIbAfcuWs69lnKoad91y+rc/L3TpS4qFNFOicxK7q/
mROEj2SL2zfObL+S5ItIzlWLgJ2XpxbV4MLeW0K0F6aLIwXtFJ0stYpJybnYl7IPAqaHNgYYe/r9
AQTxjZpItgIHDgkOUV0aA7Xneis9EwlAc36ovfuPt+1wjrD0HjiaXOLLcoJa25cv3okVoHAOBjqZ
1i3NjBQGkaGND8HaC7nkvJTzrtePFAmwl8WGGf7zC5SN3p3SWRnMUvaSwhX20GyZOKEDwQwsdnjU
j2Kx/iKaj7LQs+a9f0xGU7yWgJOhMXxVb4CN8OH6dm9EvM3/CBV5GhXcSKZzYgI6lDTkC5bp40oF
hV/Vv2Y8u/fULU3WGvpr0IkRZasU4B66ew26w0f8f3Weaub1DHAFApAULfPy2un37Cb6QgVGmc3m
5y7R7kbNY8hlGnhTP7clf/mV1m8/V+qi99UVAnIhFW8I7xeV+fTobY64yUISIg6GlB2oGElfANcZ
1RYvDep0yCu/3aQ/Dzo2r+d9vJyj5pLdpg8/2KWj5OTSyVGKRlsdkfNMsWIBSZ1stGgc9Ufj4Dx7
0vAAa8jnhIfP2iIrnqTYuwpkZx5fci9nEtC7VNnL/HP3f60PuTZH7l63hcGsXboKZQLrEvo3xSB8
PoPMeDFADuF509HHYnMCs8r6v1SBTvOa9lMei1Oih73WWwJolfH69phzU+xhf4QSSlB8k5+uS8+8
lmttXVuJxmIRkIHx4TFsPVymn682fy7dYTYF/5BL03Wi+Dd6pTpU9EG8sSrQbBbduW8ZD7BsVkVZ
lN2NZhKf4I6zwSnGMm2mPH+Pn0+GEVoQrgkUS9p1Ov3kNz7B13EUBOkb+RlJ0cfupXQsfjGfnRMJ
7USIOdkK+eR3OZiZguEg5e+sYt5Zv3jrmFXL5mbp3pjgszd4l1LE2G4DKG/P4wS9E1y1AmtT2wUZ
Wu+V9yH0BGgybO4fK56tpaP4PBSC53oLR8e4iB7FRCnGJUioYtumbxmN2YONlz7GPA06KfBCRbmT
tEeBNmx7Vw9yPHR/XkoO9Cg9LW4tkj14sV4scj768UV3Dh/MqicTGs5RkC7bsLfUKg62kC8g4NQw
21KUwvFzklEG+aSiYo64e8ODG6LWfaOYa1o4Tl9cTMies7FbOCN+4Qwj4++3HOVJNzltfQVFTpku
LyqQnWjYgVPR5rZhXPl/0jMtq8uP/R9/H7YcPJoaGywBm8DTB0YuRFs/SWiNQs3pMiM3JV68yqGz
Gi8lKUJdZrju64XAAHUT8dKh5RSodjC45qt+rprarixIcjhco2qHw7ruMjvOPAKb+RyOv6xT2h7B
5QvnrmWWLeO6MqThxu6Q7IcvL+XwTSDCSJFccVbVQmC1BTD0oT+AfiJjrk61GRpqRWuMnncJQYmO
CEtdjvP/kag6EQbanywj/x83yZqIQ+MFMsQj4kkSqY0CLmRfcF9VJXT2N7EzUQNCzkufuPX+mlmB
iUsuSm1hnNui0OOyXFX2fd9ezUjoohysKtlqOro4hpnmVRIM7TmuCRlOHLN/804pjw80oDcdoYSP
lpZmQei7GXLdranKlPRe1o+iJ8M5QwCIixBFG2/kgAqBeNftglLClIzIZPIoUpEZ+D8BGotUXf5n
ss6GuQ/5e+zfrDzmUt/pBIWFjlNU8N3/6iLq/r7BXfTBiyuRVtTH8Qt/ODs9TGWlkNawwrvEurDM
ZqgI75xZLhnKUV/0AEKBYRHYKsScOB37oLyolsI34rxWg0IJfOH3ni7uO56+FHzR1u4Op5pmipwY
dUzbj2CQuPygNHI/58e6+XC3ZzUnSBz7m6C0WoVi5an14VqCXW43S/KJ5rvHcd6IaNy8HeEW6OSk
XFkZ6m8sszfNrbmy7QSDwAKPwu80EPPN/wk5NZ6DcTVCGWbsGtI8P9fXMLlgmYvPwybqCdE31MOZ
F2pm2zHqz4Jgm00uxNMw47Q1OQhbkM/e3nOSjUbRGjlJ3ek9qrUbZlLBVVHbGEuA67gHx7K4ojN4
U/umUG2BbTsD2ZfP8dmKI/C6oz11HQwRpB8xz0y08XOnPH7JC+dv1+mseAGHoiwwhGX8WJN46o+O
t5fGKH39C08k0XIsc3hTml6Ug3DqZwMRFXahcHgjqo8AyXR9iZOAki9qVgHGrq8tNf+QuyrB65w9
tW1OiLYaHBCifBUMmjzWjegycXf7jJK9uCe7xLDIn1bV/VjPn60xxtNZsE+a0XOoPYATvzGqMXhh
8TJ/U6THWNNb6sNXiAApNbasm5N7/Y8CCZrmFIEsH32/N2CCgBQtFthzeHP+JUMao7sqk6OL+dJ+
zyj+8LCnU2NQ/Ox/X44IyhJTyU3mSILhT+kkCEdqVTmHk/5suFgfJdYXIOLldhjrycRsT3Si+rA0
xgs/87if7L4g7MfQcBv2eApQLH0rmc3IRpWLtnCMRah7tm/16eHu4UpFDH7h+lJXbJ1uKF4ANo/X
PH/3myISHa68YuowTRMEqKgTEFaGNiMg24TU8XcsWRr9bPlN0XUgoCAInpwkEKgmxhXzQkPK9/op
a+YQeueshzXfOePeaE7GKjWEsQWZlyp0Of1Z4CfFnwSNZa54gW0HXM9569RXTuMQKaGyoAKWOZ1V
KrXAM3TzRp5PKisIr1YI4FUxFHzShl5ajO+nWrdkqe13JubABbPAqwgy5yGVaICrSYQPgKEJ5Qvg
6rjO3iLHL2SyoJPDSwq7OHr2nWOindu5KuqF1kjMXFjYDrvl15l6D/YR3bZITAnPAkC6gYdLlk87
Q9ivVhDlATfVBPhUw0xPmjE8LgGRMJ5jMcMDZCu7YpkTVk6nglQZrEAH1Wg+14091Ul+NMLuj4Z6
PmSI26j/7O18dC27dDJNodnWdQ/ygoStTuH8IF/wqM9KdBeGRJBOIWTOeodrQMaoSoNj4K+7TUp5
EaG6LhoBHsHFSw2H36cQn3rl4x4FjiLtXLA2QDgD6GyezHYWCx76DEH/ey9urMk3xNXDtXnE+dW7
cX8zX5ltJ/8NKl5CNjUgHP2so3cM/WeeLByoa61r1DeEZfBVohG14/200QQGvF08uevvY2aYHJ8E
90MfR5ZUASZPb/Zgh5xDScyNLVHX35MPfdzNDI8mwXkQRkB3O+80F8DFIgAqtcPlK+A3knGtMuOO
NEILjXw+oC27wgUKcH/lIZW6N8dghV+LzPORvMLjI4VhAe3WL++IWJ96Br1Zp4sDAuo+xSVNtsgm
XtMX77Z8GGa00MijPdkPb/FqEjtU8ZGWxHjJ+YiVXVNuv0+M+BSSWCz68rB+gBRHJFkkHqud3GvY
27GLE7102hYdaTSHYEcezcpS5yubQfR6up/vLbudFTcGXbliv+7QLesInRFUW67pmkkvefTNtDvS
LJ19OEB80Ti3rqmsspAv8LQx4DY6fFXFZ5JNz/rjPsgf74G/9LJuIZ9OiRl6ftLze06PcefTuawp
nQ0p0KDx/8/4EMQCdV1z4YwjRJDnMr9/Nc/M7Kl6lopjdqsrB/m9rAv78Yhl9q93FoBWr7mjcnWD
SLs53JROZ9sCbr6icz/DEfwAHQ7BQS3qs2iCm5CdC8KIM70WHQeVLPzRund1r0BXFQEst1AVF30A
PFlmH7bO3+wwmVZMa93gfqqFEaLatDXcLaNWmlqBaVKTDOpJbD0v92F5USE4f/pwQUH5EPXDEaz7
tDOUdC5AKab/e281FsbuNe93qM3+J/RJFzz+5SjqtAj+GVO9yZqwwRGjy4y1zhXBxNImHWwUIgq1
yeZ8p9+d0NT5wSqF+s9iaILkoStutah1EHDgFCvlWdX3CYgUsuNhnuKMJdPRyJkzoYxvBvpO6Kkn
PXCnSZEo0qm/sa53ONZiR4+D26agCjxIfwyVfLC2e7TZoiR66px8TIdoXvKV+7nFO0i1M3y1gDlA
RRpWa6iqxvtG7PJy3o2738CniOLP3yneg41/QwWVEqEGtIoBMppkN4sTk9JZfQv22qpdSM+++TxN
HN5QGUx68NXRxaaNLPVKS9FWZaxEJGbQY+BeHRw26URI8KJsE/O/QXsSamteFTmAnFKkhj/BVvWT
zjudI/n+T0IZupkPvoVp5Tf8qans73TXukcHa6aUW66oWt45V7RuEUsWFZlJr6PWfCyaJsFrmNjM
/E+BHZNLSBcTPYfqfpXdAKU8K6WFfMe9vyIP/EZqjxUKiQxAo9aKXvPIYK2JM6psUWJwDzN2DSwA
PJkLz6KcTd8Ac+amGvYRwi4gOrdHAG3ouz+vMRn4yrPq21V6zmz+0NMElApZdM08EB8CQnzTcq77
NKpEtA20IUFNax6Qod+3z8HdgwJGLcVeTiBTmnEBk7Iy1pP1+z5U5Lqq0QoYnZcL9VWasWIXYzWW
UV8UfRlKDeEEXqEouEpYjEBGumEdJEQyD8mgtDLpn4tsYfdTDcTKXfj8AOQsqPRD24dV47rOnuZH
gZmQStltChizrVsrT9S2XPuV/408etps4KWqe9yAcgikfefRaPFOSn+4gAdxYpNGCX8/WyCPytSf
Qb6G+XF1dOa2omtgS/KJxbniUzzPRDNIQZ2J9vT2jwetH6FRNV/BwDKxs5bGirwEsAcitolrZM9D
i7Fl+utYBXuMUDoRsAc3ajZ9V+rBocNMdWfre8X15qAPhBNixJYvXQ/yLhKEKdc43gdRf6MD6kkI
6XM/fYbqOJ1sy6yGJ3dU85RkIue2CD4KRafxLt9N2BW+56g8/2m33RaBePmUFBpSehjkewDHw9jo
xGHI7PpI//OQYlGvMlwSdnPg7kX3i2Lr7pwHHzF8e9+XoaseuIJV5F2Qedi5LzO4T+4IGLUz+Rnj
9LdxdttR+CBAVTp0dolKjYkmcXFfmCJFGT33NfctwjahMi6PltH2r4i8c6SDGkqtgbEHm9Xlc71+
wn9jmCxKk5v1V3JNnA8TtmzvLu69LZooWuUitfdkpzWgV3GdYKW8077x0PbKXqexFcLQdo712EXE
751hzc30mzm1yNDFHG1phN+OzAJfMvZqiVe/ufKO6b76C7X1Ozc6/MV21CYV2LWOyFe/K75s8KDp
Ai8RJevNIVjp3PPoIMFy/j10Sy5g6rdkI2ToLD4CNIdjzwpfKbFCGMEiXQJnv1BXNaJ+kt9GsuvL
44mKWTq0j0ts/VoNhWGxIneeXSpvdS5WIBo98GGNZSl1yo4nLIIcizyFqs1krFKFJOyLeFwKSBjm
/PdvSLW97Fxc4+GnbBtl01uvX7avRF4blPOzwbKK/mRG96AgSKsQcfzlsNgY4Yu7iMZnrSW2jzwR
9lqN7KptZGq8XofNLan8++9Hv58cnPxIbN0jpe4XcZxe0GLvAbY71BNEoWOe9EbAr+c+O7pahj7H
uVWRfVV7YcDLLNCUxM44oWLLmoLEjAf3VQdF3OyvMy5kmBCV3cx945f9NxkO8yNzwpzNhnSHoLyB
rWJwrNGi0oSh/HKqmgAa4EYH+EjKr1/s9tgQ7LiS18ee9sz85VoqaWQ9y4N4WhbcPrle2wTj6Q8u
b90z4Jb/JbZgkJS467V7H1Zau0woClCEPHexPWrhRmxlGwnjmMmfYu4X399tz4a86NJ5PrmYMkXU
AUcsz19Nuzo5OWR0KOV9DXUUZeoGXa6gLBk4StvQ/vQVU9ovy9weM/BCBVEfpRhliBmSxJrh5Y5h
d2OI0yRgXXrs1ePItG6VdR81Jz4hJbf6SBB/bS6ZNhuYeDhhK2rUJWq45AU/4JGE6Y3vRAYLBXVL
4srN/TQ5A0vIbM7+6crXqsB4rEFRHumY3wnJyxcL2fEtSjcoXqpNPwwKSNYHoI5fjCGnMV3rS6rB
IK6bec5ushKGC6WONBN2fZnaUtIh/ua06RsyVkdUQhpM6FI4xTdVsH3ZYp39toCg5IWUjnEK3qz8
PHS9MxC0fPpc6+kms3lQRgW5nHDtsZ9XGG9EnyRnaqTwS9dF2+NtqbaWoNNbPx2CrcJ2Y4VqQqMw
WCOl6xnQLV7/u3fbvY5hcSuYVfVwmuXNNmdDZ8vZH69H4UHIH4WkR0V4Vh+W+wbpUUVySYYZZBMT
Fi/Nw2HUOzeVQ6oqe/0duTFQfmSPreXQ/Kwq5NpwauPzhYY2f5rY1DAhK1n8i2jRd4hQ3OtAf3M6
iq79cI42+NgyfQckDJr0xUwRDlVmTelt1BImeCz27QIl+0LVBHZx5izrU4Q52V71EjOURT9aGFW0
aRfVySYD6+LLo3fj00Z3BpNtScyYX9mY9LXlOoDXCtb1mZxqJyI11Gh2bgtOVYgb8a0aeOT63xhd
5NTCupHD95Dk5fbS7+wyjEUS3+T9isHLPxCq7AA25iOsk41hI7CedGVcvBlAGet4yi7hjvbbhf51
P1bphvB3rcP71ggtXLpSCIIK9o5iV2bmsvtthooI6BtFtWkSxhuqlf9K58AsH9pLhiW3kMD9ffvv
Ikmbg2puS2buL98uJOzjRgwo7llbBpnHgDJHaeiI3hXVQY1QsA39dcWBBeYr+WA0B1RKnT0pStf8
bopEVZPDiltfl/1OR4Sshd8EMwfJueZnnCsIk8v5or0ybKHpWo1xfTEdIpebJYksYtbrjkO9dcd5
tvvAROCUld9jrXIeOPimHa7ABte/IGOYq3Qok6NItpCA6q8pv8VCdT8zDBqH5jxUjefQa4ZzMIBi
dtgtQWmZQnQp0dYgfJW3YTRWjzjtSxRLK6vIFH33rpKQpdbKIZ1uCzga6mk1k0SHarcRNq6JMZfo
GZR3U1ygJZAVdJ8S1b0uZQMvA7wDzfeIERerBUAMbmIdLQ3AZIDp6em6kmdF/sq5cPq5fHPE3rzh
enaQEfcFKmZ/AvjfxGG5CytdBA9bOqBI5k7/Y2+w/+T70F7flga+FCUT/q1ULvZB8fFpgwb0qE91
2NLYnwE8/DOSpaNKXcEEyZyxH4UkyoiP4IQpOZembq8r6WIRtBavozQh7WJyVcjoAt2Fe/lcg5mX
VYBi739jf+vkKwNhCuk8ikrugbXgK+q4NCAHpeeUEJ4Yu+GDYAu6hBIlrgFIs3UvEnlVZvPADZ3A
k5hLwvcw0ZqDAm/URzXgqQqGGXqMFCY01V27fS199MLqtJBBD07Qieth61wKVuLdh1ODfLTpSWXg
oVsGKIVdOz5IJQaN0/AZEGvBwgzTR8XJ4RFzLFNanHODvruYedpfj4IxHjIntHjatmObSKNrwm1y
AM4GdYjiTdX58xyl67btyRGuuQtuoc1mtJoKMSHv/DiwneyrGui4oB1l8+9qUEctb8BAHjl1lnbs
6OoedvQRTYZyV97n1PPn3tqw6LJruVUws2P53z6oNmr/pY65W1C0xmsTFInpIO4vdof0ZncrpmzR
Qj+rb3DxxKtlzOoiOwC4dXf0p7YPiZc6XjsJza01qMNAjdq7RwjXKO8zjD6uknLlp/cd+AVRhgSr
1ST3gpRoXr0Bf9MAHrjctzkwloDcCsSLeVhv1zZxiMihQzndK4b2rZxokbhUtpHFNZDObLqNFveB
m34ZYSmTBBQexYs9knFbrE2D1UUmXsG9J3Yu4peGKg0EzDa0iiIeZvY/G5YPlxLGlvwLVWQBFvT7
NtB5VvB7sBPyYiKxLVHqL3NyIHucNnEdPo25xGLkmYm4F30u+Joscj1logw+ZccgUuwWD5gPRBEp
JGKzozrPxx2Knh+OlifYhUIsgx+IrazaBkbMg8ZHTMRmdhQOzwRF9ekpSOCsAhNBJxH+BTqEDurd
fyRhmgGqOCZrYr/DQhgYG7IUxHpQdIIYkF6ZvzQManyBFqo4uEmrutJaZ808B2i9bAephnitMYPQ
JRFxmVfyHEoA7x3FY5GfTnJL99DW3uY5uE5EpECSDsVm63HOhri7llOso4qWWgOE830vo1dCKCI5
HWM7qy+CgBdlZ5Vz7JudJ6DFXdgec1tHI1aAiDKH1bssMgoOlzHB244tKFQ2+2cc4nEl82w1Yr+X
lRVq1YK5dw2KVDoZuPTbWkBXSXiEZbbqNa3Kb4Ir3rhPrAg4JlfRp/13yBpDNaLzcdESxDXkwHlH
hTAlEdSruXuvpze0Co8p7oiFghe/SwGGv9cSS3GnCD4eY7nyOi3o2gvETpF+w9fNfCSRJ8/Fcq9a
mr6ybHmBWa4drpti0C0TPL9gzioJZU1KuLaZOOcZfW+udE4YeHYT1M+XMugC/8RVcxcoJ4Dff4Ov
zOrVt8alCvg1PYFpgRP1UwIjb7tXiYJLoExKdSyP38k7+rXLc3Hq3MIiO5OL3p+D0e7O6oIB0qCy
sIy4nkb+EeC1cpemS6lsvzDPwRUI1tvuZ3TUSkQGtsvpSrRCgmQjiPCRuFDRwGVNvpkp6t0sI6Zb
Ld7i3+09DSD0ZAe4c/VAc4tCmtnfvvnMXTKOdrli8E5wSN8x5FwU/R88etYFVtLu2gwHmYwdX6/O
FfmDJgrFJXJj9EfAFVhFXU6RWabSfvLB3U3Ttp/BC3mQbXhiUqwbd5bGW2EWl8bYhUVCi7QPRxDN
CHytAcQW9+YerUYBn7dp0zHK7vjb79J0gXkE5nMCcFhJfmBM54L7bTS9+ncdDQUfKECObOZ8iDQH
1sQc0loycpACiqA1zhk1yx1erggw7ojC7efEwDfrSyDfCr2J/cJTvuvMc+/5vCciJ0IRPWch5SDd
fXBiASWFvobGb6jGZQSBWf3b/NWNQPi0qhqI0ANtAShOp2a9Gy9hiK7w9LGyAaMogLendLTwWqnY
2S5FPEMQDgGFLrej70SNWb423c98FYKdU1hjPhK3SFKuwFton3H6CQIo0R+9J6d6ZoIS7n39AvBd
kWc0BL3oM1ryiCn01s65W3stL24OuSCOrDDepGd2e41UQu7/W876AuM928CkZzUUHxrSuEDzVPvp
bKeTLjSjgRc3KR3cLgpxX78DTzYJyPtOU5WwSMIJzEcq5f5kTh9vHPp2bxXGvt6l/UJ6nhI2iwaG
eAIc/YdZPvYdeQ+sHGFDFE87Oam8a2lW16zVOgmIhVd2b0CxzCW8JpsGAvS2b62/RpqawuvdEt7W
YkCGPPom/s9L4/Lw3CdDCsIXw+j0saxCuSBB1WNVFzW7Twkr9xKElfUfBYpr5JytfoNG8G0e6vCv
4U96a3V9/bOlpCJu1CGp/aBNKL0a+zeVNugjl8SSLv6ytUrkLVswMzHzpo9RUeqeuYsJaRvMF3TY
Giy6vhMKy6JDjfbruWQ1N+gJWPOyMMmjPn38I7t02vieIpWJk07p/xGWVEhmiESpfMQ1o4OVfIHv
D9nQDV6e0q/3MZeFlsMCYWZNLU46oU7w2k65KyQuIjnzEIAmc0Gmb5ox3yqHu9Q0n7KR0TY63M8F
+vmiX6FHyZtY8pm5pk+a99Zt9yUiIEvQu2D0dzB546aqjRX2iUBJSzI8NqRf8KbnKrOEyrWzZhdj
zGTR/AmfyZ9o81MRj7DVV5lw7OSegUHRs2XRdpj1SKE7BtDKQ0irpX8U8JH+nHNbD10rUTmW9CNQ
d+pH7xMKY40aFYg5My40HuUoedyV0E36vwCCieXrGQ8XoODkuVPWkhtGO6N6yGjMzZzg+nBjcCCI
O9g7fpdD5YFUWUzMgbMF3YOR80FmgOLF0A/kwgMfqcwo6BYB3PG3JHYmYbg60YbDDkY7yXT7QSAQ
T+LB062LS3ktQsKAAf3xIuOVXI8BNMxZMuLQmTGl60fmSnu2Nwsv/nF/6VXra0+EqzklGiUISs31
d7xZEDWbj5PxpkFZjNnOvx+X9pYYeVE8OiSnpAIslDb1LbV/+b1PgsBlUkR95QbgZIUFJrfyXGBM
UpZbWo+6bIrcZlfrz63as5eTbEj5jG30TOx8HEjDa9sz7xGDebuKUOGKt7ZLfsThvZLCC7CRLD/8
h4rk7TpxBs37rnaXuirzLL5S9RnzTOG4VPxrdbUBALtMwc7cUJ6mA+CuMYBccC5ZkIhCTm4Oe3ef
o44gcreI2FBMQjNusSa0SJCfkLBsx4GMR86GBFAGLYXREfZlwruZvNsvqyjAnKOPmYbZ/qrtKKFH
A4ldG2G9KYPpngVhNbkqNwYbaggCf9Ow+CvYXJHEAluBaqGJwmci4c6z1W1MhjZIc2SJeTnyO31h
EbK3DfqTyM+xF6QLlOmDq1mU6bzr73KXE2Xa/94q/akdN2JNkC8WqYcnXWBEuPyxpQoZJFMpJZDB
tciwX754u4Rp0Zinvz6CPRMSuwj8Saqd+gl2sMKcWl/tPtRBC+VD8gOHrKMpDVAQbdEa4G3HC40T
aWGXcAbs8SsjuQ29GMFlrXGEbY3Te63kvTkD30x1DFiyyJ6ElTwSFPVLxY0dBvL/NgkSvqXwLyHe
PEXyF+RhcEMFOVbj2jfwEM9G2RQf4PweDmOyqydfwI/mz8BcHdpbkxI2sfpHamrkeeTIl83xh0fG
S2fTe3/UZvkdkmeh2P0H0KaLmAMwHRGUDDNzs0eIctH0dK7wAlS4mfiUa44VyYE3xQCY3Y1cxVlR
I75/COEFCLtS8g4QhWZPlS0JEKUicCzDCcw8hVaIQbnRPpbpyd+B4Pvy0JMWmL/BcKx8mhM7SMOj
CNc39pwA2zCNHU9JnLflYhpqcT9Ok7Jft/HZ2BVZgAEPMMXid7wzcbxO7OFvUtAVlofk4mT7AQsg
nHp6498OFcV3BClvmZMWPW7UXRtx3qYOLdtI2b0/ZnlTAZ/pAZm1gUZ9h7Opx4Sz/od1FZfU+Bnp
/oI/arYaWX3P3PYQl8d5LkULTkdHnJwowgR/PLvzHfr7c5yq9vy3dkpFVme4BPOcinSZIIaNggem
VRrekfRfXMbCMKcEVutlV9+rQOg7eGAaxBpZJ6GjyoWAmDp7aX6+Hmdc5Tnlg1Wwn6CVrbf7WF3D
g1KmiJ2MgSWIkFcy44pDLiZSc91eB8cNyQwEWkWOSphC5I9NFtwMNC+MPejae90S7SxOmWVnUXTf
zo8llnx7MDFv/yfJpBVd+kbtJgNnpE0Bs5ZZOq7NU7x/NGJkTjnc9Xl8w2rsrt9Su2hqd0dxfgh9
fYqljaLgwp58ai3inMZgkwuBk1dqwsNP3vVe2x4wKwZ+GauRnO+uyJRMKmLdvyTehRrhIaz6FhOI
hzZ95Z3Z9SpKFgbLmwOv59wa4UFCwgQ5sDfB5ihUGJw9lYRjZPbWQ3NpfnQwm4Lz2S7jhFXyIlpu
3eexKPOs2CJShT+EGuKYzpK/InERCiEtAV/+sYc4m2A0pENkEG6LuIBJJ49+bj94zg42LYidP8XF
C/LBs5V2n6wUk1201BaVUpr9Tjy7Qi5N80ijU4fmZ029d0I6kOtV8GYiNvRRxhPKPUkya7hcXAy8
jUtEsO/LO6GEVqoU8HyzNi82YYKNXQg6yTXfthFx8FQC7TBkALyxIWnrDh8TfWPwelmtAa0y7cd3
ODrB3y3DPP6jJ4Mdx5vwA7GZ6jGo1lZqrLGsvRQ+yevlnalFHxhJed/lT7xCqGbuTQHpi5xnHEMF
k/2E9yfl26hpC4DA60AQwo2P5C63lha++Hsmtx0R6ewZEfiKrJ18/pKu9jP8gLCx6GKmTX5bA4pP
zbA0jv4aOD1X3v1QHSyddrC2Qd7S/jmRMH9mBhm0v1SE9nyfuCZq+cgITUFkKtvYShjUVn3xSqpS
5KEimTX6EIJiHptR1wTXCZEdNTQEDwtAkyu8itQ4JxxzCy8hyCR8X/gRt7V+5xmygVoZ1Q7lm+0r
eQE+fytQBznrIKo6YnkfXUDe5xzE2U+RvbnvfAJfX1UtYS/YVYD1/Mq39ywHdJe7ZSlgaQkMzPi/
+dfozmVnX64bWo+ZJ8WFdt0Ro7CqD42FE+W9n8jVE9sStKny48dAjEGzKhb/rTNEXB2apcvb7rjJ
ZjB7r4HnUM1BoJQ5Za9ql/76AQdjzeyge+FeZio2sA32mDvYf16WdegXyPo4PKC44qfFd1bjuP90
rOh3OEQlxqo4Ab4EqO6nA9Uw3kXlzulllgDtyYnnFzy1INg2qioHRCd61j3OMfs5F1ENWjkFF1/7
tV19U41KTKqJuU5kMQ1/SP2nW430DhDMjioxh+0OshjvRROPtunUwWF/iAP8enEkHT1lkFBA3W0v
dLbSjuFgfCEHsCs+ytjO4PcRu7gG1l808DQX+mZBDj3pswODNMxlGES+IRGYpaMJqFBbLrnmmwZP
LBAldjpylQU2NJujebidvEH6D7G4tK68bGWkPb8BhrtZImBi6wvVDsb+PZAfdr5JqzNp/+cCvdmi
FhST8lqzTzJNIIsh3MdjsdNzxTAGpSbK2NPAhFqtik8SFko1tKm88Q5fXHBDeKTFqwRj6+cruVgQ
yQ3LQw8n/En/sIFWGAFJfAuAR9mTQiueA2tdNicrsLV8+7WhEpHbCUocBNhrNhyy6It0wBkQmfMl
t6pgY6c7lMoCrjB49MUTH00+hdDZiBVk/lb+BELMFz+juSOVimhwKDAUP3MeT3QWGZU3JwCs54YY
IachKs82KJscHi6sxbYXPhqMopv0Uep0YfxMxrDKFjVSS9kGLCeAB0XI5HE8uJ/DrtRnGls9UMB8
5HLtLOs2aFbZicY3AVF5CgnIbnNG2WKnOjQt5vWM0caKAkfE5foDhn4fa6KA9ThpTSr9+VkEhyuO
VSuPO0WZOSoUV6wmV6ifl9zlkoTxxN2byPJmyKf/kSGJntvHSe0C4AHjayvAaDmPkZSXf/bKKwoU
bP/88Yk6qDQxdbHERc4nRj8C1grEQL2qqn1z2V/i3Ut8WFwCktN2ogOap2xNfziPI96+ccXUd0/G
QCwPH/0bAmOc0kcGa1ZcG6lqkOWWDrCq5hsz302Jrcld96+E2FB5QMLETc3Vh/Lrcr4ppWV/Wqx8
r9xH/iSXW6YlEDUpx6NlfhlcqRplXcnGofVW3p0Bb2lAhX5A2Hiy7Skw8Z9gBFTss1iBjIJqiyc8
CKuf19EV7bzRJ/UpbyJEbV++OgbixDrCzIRCT63WVkgv3yQg8GHNVOcctq7lfJPzNVRKutJUAA4K
goYy4kegYwYqOIv7YOSi7wvd0E48YnWuujQ2e/C3cUgesB7EepH2iKHYJc4PeG2F/MIciDl1A/Nf
cyjwF4ocprDgCdbgNckleJrH/Z/feoJ/hff62stGX0mk4Ofsy9GQVw9gD2/htGzEiWFGH/no04sS
64yT2P3eI6D1cJgN+rl2T7owciTEKWSr0LcKnSKb+Mx2BHcIGRbiPM+Amt9qH7obXG+qunSnBm8+
AAhFv0Fa5hhEzZbHkX9Ea4VxCBuu3KzQf5vOygRu5w42IjFEtcHFG+diyX80Pe6ltwpJg3lM5hC8
pjcKS/YxRmOKcsFcS2IhsPvQusMKT+GeGBQymvP6ml1jQDcvZfmMVf5cV58AEPQ213r3Vk0k3OdB
BIfTEsCv+ALGDKm75Jic+m29WoW2PKGdCgVOolGgcaR55mR7cZvYUza7BrgemYL1uAD6+Sp08GTN
3XsMlH3+k2MYuXm5/zAQllRKeIekhjPy4ZhPZLIJeg8dMEN9SgC2JSyAfBAg5RTulqg4qlZS/hYa
UB5dDNKJ298hNEUcSCp5awyzq/Kte0FlXVV3SqMlDccA9NmA2SZP60Eqi3WamwVc9QJ4rI9Fd6z0
zPu6l19U6f9x94KEtIBw60/59q46Rrd1/ssk3pidTo58GHxHtJLESTrvf3PBaFJM0MlEeeEA6TV+
SCceBtks+7Tn511YCF0Ec4rLx6X64Ac+43vmC4CuAAqzWXM0WGFBoDFjDzk+5vwBPbR2FsU7GrKY
3RuMjAg7MIu3XWnwwJa2Y0smR2SOq9NZJxQvqyQavMZgj/4OI/MpHvI0oVUjUWIuObxgqf7cx9kQ
UjkbckVtCZohP/+zy2jsAGrH/VMGA6GzZrsMQoy0IsdVPWSjwyNx+fqujynt0sp3FvBv600Amr4w
zCaFVQo2BUppu73gQ41GdlNjsZtxCnimwDq3qvtaHtj7sMfnlogB2N1KKO02L2okvJIbdjSWr7IJ
k37UtRTGnXkScto52PUG41pMh1GZCChNJG0VmRh4P9OVouzCIHuBuIWyg0xiK/ogFTOh8/ESy8AQ
oMj1sY19+bqWIScHY15OrrrZcrDz8vLn2SfPAOw50J5OBYJcCeCZRcHRIAZRqngI4qqAaoriHO2v
o6mbHHSVcJs3Svu6RCG/kJwF9r08ImeQwVZKx5mtA2VMgB+mPk5WcItyQukMw8yH5XB5Ogid/af6
ZFG3ya7kbI4H8vjpKooZXeWJjUrC0CZfozkCjZUD8ciRBf9XJyoXI9/zXDVaw2dMMVMOVteT/9zP
++Mmu0AqngcWtNFfblFlHdAu/PFF1Db74Awumft6DZuPssIQ/JS72yilG1BPpWdl05lWISqwwdnh
LZ8u5ApuMc1iUh+eLuy+WH76HQd/cTEAy0kGcIQe9r9xKkUo2UetYoEf6Wd5vPfUeziCLCCDOr4Y
71RYZsLFUz6+sNO5XnVm3OLVFgualGp66pUZIRPTCFhBueJLD24jebcAO6czpr3uqkjhKZXoOT8a
RDwX55Jo/+rp1rylKABBb57SANuPc7iQcngGGMldTSNzysNcBtKzbi5PO94eDxwin3MqV+tS08QS
OYtM8Bd50AbzNuvpeSZqh+JcjIiTvcWfd+on1q2OmRgrNF9d8Pg8zAbj1qIxAMqG4ymjn+CR5xOn
ZIg+VwPdc8KIFRjGTSLJ/hp4iYkdOpcQfbz+b4l2VwVIEjrEFnrRa1WEZkrUZvbcFH066YsYvZVe
9tTjjOlhPtHpD6cILyZ1nP7z3yX0kXOE6d1PTY2uUSdbhNlEHV4RjvMeLhugD4QOo8q0MjOLYpBO
bFqhhB0M13a8h1WsUR8GA6GUbF421d0iR/BFBm9Xlvc4c+3eGYIAlcFrwzGTOwPKXsig4XZPPi9C
dKydM/L9+9uDgHzHiEvqe6rCOPoZSJm4EwqMXKxEN8f85gwElE83uxNcpT4chFizaDusfEabELdV
QvELczZeCuekhV72BD+NC+aHTxum2VICNkNVYNDh4PaTkjGLNfGtWusqNH92hjTo27+ccIZa7iz8
nuoOZAu90WI+x0LHs3Df4w1I3tgef/qaFa+b3y9yPHfQo4I9U2gri3N3iyhkKyyRdejFlhtaXtRd
clbPrhE1fvvviRrRohYHHF051kOogTyIUK8pLS6jpmZDDsKGhDrYrRWzpeYR/B0l9daXBmQ/UpRo
dK5S3YZekZdPnUz7n2OzzTDFzMhPvgbwtVs6RAmAZYR6dUXb0Fl5eG6Ne3QUUG/yjDiWit2fevnH
kDq3QyMAeSsF8DYqM6Tj2ovXmlAP0Q9iGpsHKPcx0yF39hYAG7tFZ4D2MmVs9extmNOyi7OpmwMV
uSxq9a+otVkUMeusHlZa9rRNGMAddmFCY0fxh07SLjpoSkzR/2uEOPXvxRX+7PQKV/ANnyELDxDf
DU0pFvgrmdIWJhkz7EL/ShyuLSe33orQn8xEGz9qDSbZusZZ8Jynxg3GSMscwp2BUiCze2aI+ELq
9GGjKktYPhyeckl3TpQ8e+aR64mDTl5q6paln9MrFo8u5uPkuhkwFP/ORAjfI5HNgoC2PqpvYXUc
UR0DW82Q63udTKY98uiwtXApiY1rzXFuQXK/LPer+5PUzgpiFac8DAYUtFAmMHxuKz4ljU/I5Wfr
UK2NnMBO8EpHQld9kf3xtxv08mXhapkuyT2Y0hrVNQPnOaIJ+BvTOWHmioi6BCPd78rSIOgH8aZe
RDZY7lTLvjEC5nz59sdWAxNyZsHFhJRs/FfO39GaYQVWTtoIOHqvObWBnzzmST7YimnUmpgJE7yd
CEp43EJpZTD4s3v1buOJyVDiMiv/Jhi8WoUXuBvkermjWfY+15h0vVCw6s5Z2DvuHyXvHxpvtVU8
elmjJlZyOiVrVVi7/VSE7RTs8C+z1QGMCZuUx2bmDcaNdDl5ZuBoZxWJRd9au+p8o0UllDL4E7dv
FmK2hCQdx7mS2TGDkb5AmKcJP+TlT9VsfhGrbWQT8SU2IYAcHbDEGIZTVS/UQ0toS/jjlv2JAixK
5AfdyXWuagjLZsQwjUNyuIZoi3a50mA2rPQA6mU9EsGyF/NDrvbiD0snDooV7WGululLcs4hJIa+
z5YSt7ehxvQ4slT4bxFC50QnUPa9mpdYzqsYSjalyjqAxKKERSCNi8dKawzCLUGSardr1bYsvlzu
QRfkOgX/2z1NW5ixd/lu89Q+gV5URAwxU0dt6Essxol/cbJLfhxrlwVR8B0BEkkYaI7S1BMzalz4
EugKOc5IcZ2hFpzB+f7SNEgko8cDwC2oESgYcvf2Lu0kuu2vNK930MuhCpWWHUYido/0KyIPdZU3
KTI9prPK4IOU64MqaEZbb8zjv8mJ3+FBMs8glMjRZM/7uDKUU9zhm3jls3F8nSJniy7cKp7CG4kZ
g/dZTKRs2OFNatmd4IV9glPlm1RQxyavEOwmrHKvT/bQrHqLflYcixJRkS5MAVXgZby3a1iQsnhC
RVuHb3jPLJl9Ara7egqsEwUKE5hBI3GgR46QrDcej8RId1TG01VPHY1kLLHaM2u+E8jQIH+Amchd
vCt2Ysm4UB01md1ijvh4YgYepkwlB8ZFiIMwBWoJ8CdCoFiA6+dunLWpXLTWQBFYP4V6fhtPvinB
pW5EUumKtduVw8kxObnZOj89B5rWwtiyIq7MUUQdK0FlIs6JtkBiKPo7sPrET+bU0PfvJ7Dsx8Sg
DRZjg5QB/IKOahgOi3IpbTWr7y2YWIK1SrtOWZlIuPUaT5j1O3vNwsjc7LdkD6bxxSlshSjLwOb9
F9uXFEq54Np9n6jwB6vVt3IkIRJ86H5RHWy+q7ZvuiHvuFXjkX08H6DeSX+BaAnew9+qZUTgBtDz
hEKERgs3eRVVgtKnec94My+BA9xKGgqlHQuxn+cHYePaMMBLQnYKQGjfjAuH/6lvtFqgbg+0rL+/
Sz/TrcOgdhooOnTw66alz9PRdOc4FDXivCzCz26MwnxHfoCmZn7f6pbvqIooiJCg3CUTp51x3WRF
cArYK1+Lk+p/NdcRjof7brZyx+I/NvUCTxasZw+1oQetTVgnYaL2LNHnrD4ol1E+eNwLIYFAGzkN
tCNZYFQCSehw5m/zi1RRowgtjQCJAd/J9OliJizJrqywCFV1nYbZmILFZuqTuBUhtIVfEUOf9lpQ
meSJdQI+cFK971Tkts26/SFheE5RzU+UrJDje7iLFt4mtZi6fJLRmReEDbU+hqkqb1/jrN1aufsp
Exl9dszrIB7lMSp0q+sneWfoDSJNYZnYNws77F90PiUpug0bEorPdR6X5e391OK1zjgdyuMLNqGU
8vFCnEXrjOdN0xFcvnhlOZjU6UhUFeQH1pz0TW7MNjJvWJTdqUo09z+JXcDxizW97DMPHpS8jBrG
1PnIFFIiFCz7jVyKc8hBBbFiTcodzN/UCGOXWubT0HWBwJ+vaPQPECdhbtW+7OrhCHZ5r6lxEoim
tDvuqV3FgO8IvGfOKSi65+YuJSHzUF0BQOsElZTrhj+UmmG8Eh4m9rFFKWZfgDmGc6oX3n4aRtHF
6vftXw24yo3YfCx+0Puu/R/n9H9lWP701nAdj1iTJ1lDGgxq0KrCviFI5MujMuE4brEgxQxFhV6X
Qj9LvFJSK0LelQdjNkuu4NO0pd5sXIpScwXiALAa+1owmnLwralYslk8QA+ITADZJKoYb5Q1n/c5
HjexCpfa82+n2Yu5oV8nxNtvyK3h+g7a3t213CJcWDVcZj6Dwg0JvyKTH0z6QvE70ycS9g9z1n8J
K+sunzLyMbgwpRusxdsK/+/pF1iywmU5cqTQjdFlDjNcfR9Jjwady8kcNnsOtQ/E21gWI7ZSwPmp
dpj9BfiaV17RMoWCs3Vbffp9io8tk4DrySRIWQ8kGRV8e/kIrcCfijGrYQp8e5jHNC1NPqdf1Hoa
C+c2fD+A1GqkLQcEfLjL6xCxR1/3BClEsymH1WmclKXr+P/+9MvPJQ7lCFhVMVnO24uiCkuSoQ4z
nblhO+HKWSjVl9DMQtsESBxBZIJDd8yz+NEFJvvQhB87s9FeIXYyiAz13RkvxCofHbR9tRfEBKnR
oven71Yag3Hv7RTdPKfa4VQcXob6WragBTdoonh7yY27wibHLqFnTyXSTdecj1UqzZXKt4yabgAh
KmsR7GiBFWZEFtHWK+Oz6IVZwTqk7OcVVdGV29vy9a1sAE+ZzZ+IAzQHggr+b32HUZCn0RgRDT4b
oC/xHrqz+To5SRlxHNfSbCwiBDVB1QL4Vd+EyDnRBzwsJeFxiJi9pQ4GJoeXRSGKbovtcO1/x5Nl
e13kOnI5zX7qRWZ5OU260aScvjtp6WS7pUZOXypMBQfWeDoGNGAG0Fcs32jlD8Hqmxwu0DA+nNBv
JOdqdJx22JntzTXETRKsw8i2mIv3tAa/Nh07Wti+YhLG2O1ui8qRNPSQ+GjDfsJ3SHAmCTygDYIP
qJ/MCL1pQ/Zz486Pr6B/b/+MGb76Ii3cuR5XitaxvLrOT4hv6+GnwsDGbVD/nTaLBmZVSZ2JtOO7
Ei26fO7+Q1HmdCytn/pf49YYpcjr3ZWug8UQjIlZJfTE/zNN+5VmVLhGVsS4SH7u405FIcIdSHvp
9Vdl9snwJP8JZ8v7shFIHYtFr6ULeQJm8lH9QVCQm8Lw1DCHPdlBJzY5u5DHiQpoLV6DlA86R1rw
+ijZ0gOMipC1OI4SJttrhn+v6FuumJdWz0KGwkpACnbquo1erOmRmNdc8LLLcXc5i8KLQ1oNhV8d
6dzXv9fmQvyuXlwZXIdCBItkuHCWXH6jpxIgNJl0gxqSWw8tiIu/D0pBPLJSz03ISwtvwrmSQK78
uvQ9V+6XZYx1XDzDDcrPC+BoAFONP8gh8ssMHCWNTLD0Hbd4zXHkiyyYEYITaUOO/kimL0uSyiYZ
X7G+zyidufiFqVzj7xEGqBqGzOYEvonANJSmFpqLFyaSL5+AtX05eKz0vaHykWAmwQLnVtLsZ/a6
Fw8Jn7vPntWZqqSCZ3rsbMlJeWWQPIeVRV0KHE3kxkdMEsSG6JGySyLm5dWiA0PVwlAntjivjmKt
qMTR1XxyIyFN9uNc7c+kN4bjH2FoGAcBI3SVT0ZbWiS46rmjU7sa/TbyErhWhV59CDTEmwLg3biR
qrc7B0wIg83F9W2o9fmGlSjXZ7Hu/7k3xDM1WwSmD8+m9R/02re2R3yC+isg79EUoYlQarMD7+Cy
XrI37msNV+nM6kACggMQvO5tZ31PP2l3qTm2S6rAoH5kTqtBexgfVy9MlW+hBhBxX54EqXrBtHPt
PJXg583aGyKihgiJp9BCqEObd4YJ7oT4SqOx8TyovU0aM/i26bwMgzKdwd1/Cwr+731HM3VGIz+G
XicJoaSdOC3T81Sopr41EAkI8pI6/S1Z/Ht/2N6i7PmIpK/HAWv1LwyWKIyzYYLicYtRguijJwSv
HK6FdrupE91MP9GdsYQR8eRchrujjj+uTdlBJOkrcRkKdC6Ig26c4nkxGNshAAcm3CtI8+LizPhE
kXmIu4CWcaMjReHJJNdAiLAzG3zbz55VOIjEoIw4AeHInHXrjmrq3K45tv33KfpzcCuA3U8e7qZM
b4wrxQfKPjlOg79M0Zi1y0AXNXJcv3GEX5t8MZho02DpcmQ/4F9CKiyDJkAfin93TgwJc3hNLw8A
TIxXzBszFvfbwzLg/10rd+2J6J25MIOIylyP6OCADXew9vFvp6pB/XnQAGqKJxky92GumDh17qhC
qOHfaLTUp2B7zZVBKf0Yj386EFGmAdGnawyi4HVGdWAO3ZrWY/YqofWgx0ZXQ1wY2n9kGdRSx243
WZpHN4dHD/tknHxDWv6sUjSiB2WbR0ciWVqrOyDsHRSAoY6j9VJOgmEw4LNpZOAqU1BM1KCPIDzW
0emHeclBg3sDYYdTMlC+BSUEmdVBbxp+ASRVZn6/WHyaxvPAIxtj1DO248cxsGzfSWWL7E7KYP5R
OHlVfY1BPpbaASlyzu6AUKuQ+oaKnVUrEMPBznroqkCnq7S1EryeKOdJs9EgeQBMu15JppFPeVsO
IhIb0JdUy7g3i1K8xOOLi5ObprnbwOyahYKvW02kCjilwpStGXGSJuGhHTER2nvlikFjrNL39ahk
daeQl67uCK2N+vcopqwfzgyByotvZj6OStW2lWOsSb4SXgBvNmzbiGFYjMYPVqQ0BkSZIpjL3mLX
liU9UIsayIxu/4zD7tHMdjWk1oA7a/oTk/MdGnu7nMoBI6dABsZFFneFY6Lpf7jnORLU39dfeoPo
D2XFu4l1wGqamF+EUOfxV1uxmD4sbKiB6oWq1u4TfKQbBrgjxqdpDYe+rZtINTMu/JwVFbX4VydP
0HIV6pl7U1E+oStJOXXvxje8D8MFiBntQ7/e6lacAWwT39r4RkNu3AByLgC41TVlrm7c8WcGkDYQ
153+an0+bbXjvElO8NtUc0w/q0oAC1KB12kHfhU4AgmKUgTnMNziMjQCPDA2oQlQdz7HNsRbqCcB
7TAXh6VeWMMYwHEH/SdgbkUcd81z4jABuYH3Fxv10wVb5bq0VXngnyg9A6hR/VhrILUMxOj0VOr+
c5hEbRw75+GRg7K2aSuAk7ynoWjArleCb68MA1HAwAa4dktjHVe16Fq9LmyhDRQVE3Yc01MsUr7Q
PuqNfSSZcwbbcN315CDEpQLBscYzbL26J/5IEEwFlLpQKVkrfdz/nTUCD+/B0BJKLSTHy+Qhz5+o
8+oyBJaF6FoUrs8xppT2KD0YYYP7B4XAxGiL41eb201U+tcfP7e9uu4asRw/IU/j6HFlbGZB7hKZ
hoGq6maOih12VVfZIGwAF8YsMB6383euChxxq9rEu4w/n411fJbXHqIHsYqEShLKEKysJWkOOyiZ
V0SwFD3sXYlKUuNP7w6P7SMQfBFCI2yg3m880F6xuGe7KpRcg8ZCmdtVd+3pyRIWkJeSqI/ec0dM
yGHg7LgJK9j2zFjZjCIdgtcYmoasEOjMsYZhaTw3CX3xC6qwmy6/9j1SE0KOrtjlGPw7B4GlezjK
/jyWfL7Dy3ImumxiEKQF4Bkubkk32r98lY5h5ldGaBu+52+mkuVRuz3RbHHTAc1WwJlUO5nQ3ULq
1xCCpptu1+2s4TN0IomsU9O3nncExTLogiftOIIxpUOi/l8gNlZG1tj6C8xgQKQxWC4qEhUp/iqC
rCn+ZuYbgQ+DVVd2nIsdcjHvPeGBIB6rCYk1o5dA9Wv/DA5o80TBs3IYdMFBXq43N9HNr6o1siBF
eeHVrjW0BqHuRUAybN/glTa0H756zzuqTIG7//RoDdGMnj8MxMf0qdXEpMyNCTmioy1Yeo1S119f
H52vD90/4NgX5fgt1h8tpM2K/gKGc2MCAlt/mOd7FVSXPHrwOYH0MDugTE3Rhk7pZgFmahPPB2pG
GnFiIIDJW3nltJF0fGrDAnc5+IJhkYMSG/+AtvoatASW8b56pxFMQgSQkqeeMhMvWk1PckFOmh6f
fr3VXI5fq6Dn6dNQzaK+cKJbWDKFwma4pX3ZNOQYgOlyvaTuNaJsvJuWA98+P1Oji73dAugKpORJ
GK8BbRooEiRaSqiDwfUpfV9VTjldCcnk1S5KqGr5nMpbuwmnGswFESDEoXC3/KxHeKPPnMN9/sqi
7Bbf1tNLuKlqV4qpqrYDcY9dCqJmfse+yiPzxq/1Yosp+6/NeoAU521IGGR7HD6Hz1ClywLwPEa8
N3E/gV2Tm/v5gPBpi87D0EKIO4/tcXjRYFLrg7bQlL+/SwVK2KxsvnXniOYB+rNpQOPstiyaI+Ei
7gWK6wIOmG65BZBnkjSQhq1bn21bOKrp47ISs0cEcNy0l/plJ1urQwH8usmF9fiZ1s4kBz45WbPS
qvZTSw8iFXmQgUWfgJJ/lDGKE7Dls4JKoKMgKm9qSBpfxOA79+qCMmaNqgHNc7DEHAwEHneGDRxo
8RSJXO2Xr3HbEMAlsS58o56F3Ra02UVlvpBFKqILguCu4ZHyX3+ePPM5SSyCkWQQcjRXqbfMAk1S
Oh5VwEg/U/07KGjN8B29lDgXYTf3GIoO/kBWeZV3f+atV0Ru2ZUdcTfcYKo3mrfxMZez4IvSrdHb
dn69TdL4E9n4K0VlZ76QGh4FVka0RpAbzacNFx/IQtn1D2tUit2NZXEN0+CMoLAe3JzZmdWJulsP
9hIlX83zDL1v+huY4VLPrFkP/cHJ+bOmpXDJlYUev083Egj10MN4SfjrxaS6/d281GW438YsQ7f2
Kg7E3XboOhz3ElIKhwT/+KaiOE5QYSZrQT+WS1v5ts0C0m7I6vyG7YZU4nTElQFIBUtD9l2Re1sr
YGwSA2jf+y/rJhTxjjIluG22tUaqH91Ko4pIp03LJJY1rEUk2JXNQb3/MB2PvzYGEyOTGYljHsPn
20vkAszbqk7ticjyAvIi/JamtuC6E6hUP1Bbq3SV3CwhdeOsJDWVbf39EgqFIVOnZZ/eWWu0t3mX
QFurEtpGU/+OzxIBPO0U/DowASxGkwI1JbrWJo4eCOiXLy+UqFPWU0UdGQ7tTFtY7GB3iqPcJ/hL
ImbevCMeWHGa3cGE9WFoaT7OF9dcSV4nItHhV5A6lMFzIM7Pb859ti7/7DHuRotA+c0DlenI5Rv3
jjeGo/xSasVCqXZ/SeROt0xBNa++54fNm9z7h+KBtu/Or3r7jIaDyNsQzSTNG2TJJqYzXn7jafZc
Lm1YCNgNy3VMd0iqdJuICt0QIx9OLxs3g7YotPQlJr05f7C9uYp14bifVdPBdLqR9o7EpxPAReWZ
cHVBrn3CUDhNcRPndZ/LmHdy7wKsx1wxL9pWRCjYacfhfLjly59TTWOu6NZBdbCfPlabSM24ZtfP
n3M1CVz1QsV8SOnWMQHXa2fPDd6G96TtSkCrJCTMw/MYbGekAQ35fFbEABIvKkfMAozwf2WZYFRO
AKLPeyHd2mrX1LynKv4B9EqO2Rp73/1yqnbO8LDeoY9X6qhYhN/WYz5HIX6BD5ZxRb67JjSNunbD
EYRmLoSs6xMpFurEylmwkWuRCXKvXE8qWw8dFqemXe5qYdSOZ6u4kyYvKXg3xPHoprn/thPyojED
8Im/dLwwLVnssBvUaCVNwiMV9V/r2vFlHpEjazO+C6v4/BiZEYcPFmvp0HH51IsWoX0DrE3TeL3z
h/vxj7c89TK05+o1ePybIsXvx0bOSucw7yyPVyKLWet2Mj2oPJmqihHoyCd2DJa+Ab/qB7YzYPeF
8fhwUZgT2tECn/s4QDIIEhK13EGH6qM9felBnt2Alzcwg2TqlwScXqLu8om33e/RXA/knzjKYb4B
xlMqtdlsEB+0UeMSbcwn0SMuhLvFLxgXZLyebPQpIpgkAYOGxvDmhbjME3p76Nk7v2FQJyvgZOUG
Z214i9ME7MqsBxsN4hRkXf7h7C8qDyKkHNY7kgNunWggPMJvbWefA5d9io5Zs3GaqdMWwr35Qj9O
NGCLeD3MRY+QtNKGyTO/+StoeDmQhUe5McIWgdsJwAL+SdEidIJuICHJ89TYc1X0LYekEIqUghpa
Vwmyz5UGF6ZaEm415hH4VOAwm0/zieHn1dCPZYjeVwPISLjzlBe5JqWX/QSqTaFHCrwvsW7LPftB
ABZLjEFvE2WBdaGzhB2P9MaFGw8JQTXlkxPdxql7kfe1wLqofVyHg3t3zd87Uy1q44JkNOOVIK3Q
Vmj4YSt6J6Yp4hMSLcJPBXl+HXttqAYMnIAs0YQ+ucVxj1BgJIlWKy0C+yyrN6iK+QNebfrhQUv+
K1suZDWUuZ8xdDCa/9MlsFfMV0EFXkm4XRgFAZtZw2xNYzRjx8M8wOzZ5QvPO3XTWpal7LOvlJxu
XUIrgSTO8WEbzYVgrdWDab4hr+kMqTvmS4l274PL9kAMwfB1CHEkgi6+8H66TmGyNI+HdnU/lq3d
RDDK50hJBP3sVuSlBwj4fKifHiDDjZVkzrwHs6gB04d8XSFr/sHaFfwR8bfzVVnbeY1ONcZ+/PM1
h1XjZc/32nd0glSYSUgYdna75KnKzKdYIvmQXtS0BPFC1XO2N9HWexn4LOQxjh0z5J24Gfra9PsM
Uz+YcDkNdTGjIYSUFYcvK3w8viJb30d3yOjbqLHxDRjmbfzyIXZphjjPqyr8r1h1C+bKxOM5Xqr1
XsnwP6vK1GUuW8TlojbWMj7uPDj762w4gYiacsF486SQGmqPRHX55SNn97yAYTlgDkAqlbpEJ9Y9
0Cp6yvSdvucdpYOyYKb1z2vTKFxOk3SrukxUo+07Sd+0uyl7wjhAM6hUvJfwnxecjtlbkqRtTtjE
grcFSb4TqCD0PB5zKQuWaBmvzGhmg0ylIUS1S83oiiSLLXXQzpQXN6ojzxt7GsPPaIglibPizwUp
8JDLWXALwokwIgw6z49e3a5Lsqim3NyDWuFp1eGC6qGkoimkzOugIWSQNY1yaY/Nd5IiO6vTy0mC
b8Az2CnB2SsHX/YrnLTY+NPJWGMf0u9cIjns8eZ6MyID9ZmGMmc2Q6VHjfGcmnFGvjoJDxrADN6n
VKoY8Q1+eyUEud7xMojxy45lSsajZG6DPrPAx7TZovhBTNl0o69mDw8nTxSMO6WCDDmFF5EW+fVT
bhlKDqQVptdlK8FXPS+81M+vPIeT4u3SDJgKfcHY4afgAr636OI/0qCkWRsjMq1RqosnSX/tZDiA
lvm+xbZ3jwHGN9MsAVB4Kp7mupLMV0nvN9TaCWl5c5BtVrGABGQwDLBQOXWuq4uF+WkU7w3ckE7i
TvsDN2PBQ4Q7ovtwlAZkEF5bb722k8PpqBwnUbswz7rt6eRlZ9c6ocB9CDD+3TVvfP8AQ28Gl3do
RpZeY1G89NrHDjSA/lPeHAKW2Gmr8IXVFGwuH29zs+GjyFzU7zyqHJLg+R2ylHzXp4M/SYGm9Had
aLGM8zOF05zMDcpx4Ve304odVGIQWwp5kMJbPkJA+hRGlmlwX2ITROASB9hixIk4AX3ALQp58PSL
B124gm8hd7d08X2BwQMLNSaTvH0i6ZlK4+eWQpqDNIXY+5iVt9TnsM6hfMJ7WN8bAudnHuSnVnT/
ss4enMyL0BeqsrEovALKPO76TQMPOaz2J/CTk1Gd8BCKZpthBsAXxepFQBhmUzKxiJcBlCYYP90e
wdZZgTCYSLlGNGgIkIZEIgboB2Do5v1kyvezEOmyDVS/7yGU6DiEv2N8p09kVLEFWl75i3/S4Csd
1BeMNpmwoaPoU0MWigsDCxgljy0P6wgaBv4hicusO1oh46gP62wAZ/fOpOYFgEFoKq14nJCM/cPV
vdM/ZSU9VJfsxhsY21n0JckDvRs4N9Mw0oh+QC0A3/gbgpCUSVBoLpNvsR4bpN+LCrEqBz/gYM1l
8QbpUxRsdw/ZqQ58m/qd56oiv/4JQI4UVduXtZ7P7rJj+d3vykZYysYt7RAn4hZyuDewk5BzX/8L
+8Wh5lHrauPEBqhxYjm9G1dHUxHvYqGsc9Ctn5MLVkeq/qXArvLBR4Jz7M0dcTWmxGJpR9E8YbbW
wyl1Bi6dk6BfcSGvIxfnzrbEIpmPcweDssa2r6Xb2Ajyup0sbVc4fjJswvXyUZQi8qfj+lKI41Ap
OBDt/XOk5m7TbUxwjA1fSoqGIqomSbhKMHCYDxIqxcUAho95fkL80A9sbDcshBb2zwQvQ3RG+4m3
az5DYNzQx301rg9VR0WRrm549kqwgcOJd1GWtJ1V/kLZW+Jd1VLBXhWoPduwpWg46msxxNXkzzt2
CjoMgfF56LG4HXN4t3lF19PAl/7Y8UX/70Ly7fGuA2h1vvzY0VdKZWshxkfWwNaAlUgYUnH8Kw5i
ppn+Ki2UYJPpD4HiSzFg6Ql6QE+n+aD5RSSOUKL5mE1qtIkiGnot4/kU/KHIrcJDcdwS63ccyIkY
G0bWCSfHDTx+I15Jp8UBgqljFlUWuLk7LL3/YJtsimiMWMIiWN/rJB/eS29ktrjMIQf3x0rZI6zQ
o5spGwGVwa52o2RCC3/46egyBevmCMsRGBb9EFOojYaao0knii9Itsb1FR+gmpOmIwmCfkoV4q6R
/a1tyQkDbhGvDRENIjv5xvRM7lErSv+FzsQTVDkRg9gniBpe/YWtYZFil7CSUfitHeeyI+D0y4T4
s3CloAsANW6TrFzesyGDlwb/u7Yn0HuAQz2D/hl1YfN5id/boSY5Jie4uchHfpVU7VDQHv4HVNTi
u/3MI/aihqDMSxrOLXsK81l4pgqPvdxtNFet+or+QQ6vj8THJf9DNheVgP26WYvc66wJ5zLzXuYm
bCVE09Q3P1JaNWLZEUslbVTxWbUMWctG7YHbbFxJlnlWUxJ9Dz4+se5kVurUuFo84qfuhwUsg2nU
FvAiITxwVI9ntM+e16mwFzb0jCIksEn3a3iiPCTyaykowlfI5YjxLiTSldCn5Ijwoe+q3PACosmg
4FaB+59847RaTCfiUB8XdFBbQ1WiLgEwpv2CtAZChFPJnKtngCUJQwkhKZFrRsw6tDq6INCS/fN8
TjuX3do9dHUBwx/915OlzQAweWsMIW8bkEToCrT7MYWWU/c2rkG2I3TUGgzWz1+k4q1izFmHBOxh
UPhBi/1QMx5gfWqW7A2nK8xeD3wQYhVZumyOJwb6AHHPPfY3V+oOJPU95aFW2llpcOjhXrqYzxPq
/T6Pjtpdm4tQwuvvcsjhIIwXBoz4QCAauOb/Wzg6tHqNb20R4CJpdR56Ylr1MpwzADashHrl5lBN
YHBQdEKH012WZOxL2KwsaXXtGblsrdjKO+k0D76RK6XMq4j0PRjrYygkTg9fIhTIs3YPrkuFcDd2
UfP9ubiFI7moCrKaNnPyfu2AdrVv/qjRiWcYiPChU2UAD+GVapBkPk7TYdbw6EA/wM20nKOdIBh+
XsN3+S6Rumcl2B7cVpjGNwhhxrfPxNZQ5uQT8Xo/HOkTjdgI/NKbdFjaMCfObY68W0+3Ef9UT5hp
er2++Bb33rdT9jV6XlWsFi/iR0/FZy1NdL1ZOxDAbHDwkL+4L4FvV1eU8+/YAc8pp3vsp9Mmdbtk
NWk1jy2GubRJ6sDa3jAJPNnDSqWScFIjQmg5HnNXB69OVsuDyaHU2H/byp3hb6DzIbn2zq+Hqh7e
pmDUd418Limgk7CykR1H9Zk+3zaN7NxxMaM13iDtwh82zFJ6TGfamagA3imUfxqYhpX/37pcbpAt
G4M706cG5Gh0p9OU0piVJvKwdqal1alwDC12n3xldzTXXRVdLU3PGjgQDZ2hIqJyynqpe3MNE6xq
xPBnnxQezH2T6CHVqH9dnneWOtvSRovb+00oZTy2+Q1o/mcP9xRJLDB1iSiYxOYNlrOod7Auyj1I
FdI3zy5xJw7oNEA3atkMbkki3GktEgXcdHyrpazXbWMg+cxRQubzebXp7ZzhTPi87y2nEqg/2Z88
j7zYn6/vjeD5iu5gnK/qnZNSzv/kZyBcKzRxeoONKzGECEBjFWjLL+qPqHiPWGHuPQMfCLpNqA93
1frqXZATZcGXK9NU1heKgPATA/vhZpUVcDSro/Nr5K0Snqxhlefeq4l0Mcj67CVXxsiEvAsOvzZu
IVi7PRzO2jH/9oSbbL5tGxXyG1EQe8U2vCC5v20szAYzP8ysf0vfCWG4OdpFJmaG08w3uKEdpLs8
E+YcHf9cOhPSXe5EPRA+EYsQs4wA0WVeJ4dEwycqx+r+wUdMRAeLs8DG9wZuxShfF1OR5w2UhwZV
cL+APHFlQTs7IsM8W7E7lnhJaSAwPexiVp2thy6NZ3yZIpAw5DKYQJ9Ah78EdUXTZ/30mK/oPjwa
5Nsq7Lg4EBUnt9RvXkZoDn6yPAOFeLo7blloEOCTCH4GLTPMEM5ai5GSC4OyTF6V4tCXAVn6a3M6
1cUjmSsXl9AnJ03zCMl5eQCkMR+eqeoF4Jfc8/swePcIezpwcVSMVHOrwZ1frfQINz4UgrEFikD0
eECtF5eahVVpbYXjj2YgkWh3LimzpGVOdK3tL+EoZZAHl6BJfybL4Z/JM36Sce/Sxe4I+G+GsbBJ
lyI7qMtE7i/O26pDENCa8V4qTlbRCk1SnrDD58Elkrx7TdZArxpDhq4DNt2JOL23ahvCCk/F7G2I
hZ2Q1xj1hNx4OAhhrZM0Ayu5mLJAYek3sfCJhog+V16BUohKy26Es5J3ZH8JiGaGPXHlwC8j5/5U
qDVsNzr+dLcgR5JhrasJaJalbO+zPa9IawiQtbjtaoynjP74aNS1XAammT7NQsUSgGHbUKGDc2xQ
SP2+FbG0wPADML5YgkKEC1iQmFQhJnOcBfhQHdqy8lZxObRzs4FDcGR0QZgcMIdrjT4CrJ61EcHa
hUksetijBPgh9NXtA1tBkXAyX0LhFgCMNkaF+sVMnC0RuJKfDEbogZWIxOZyDCbdX18gKylYJH6c
CSfm93xSY4tU8VaLwfz2cr1en2mGEBwqeOUv8+RaOR+1xj8QDnZXZfcMLROFRbgW/uVysMojjuEz
ebrBBMds3Ox7eXMD7OEWXCuNvM5OfQuVj3kMewU6WCuSH7Q76evxF/DzFyGVDfBFg3VfCiSq3FM9
J5PYwrO9+bCnfXGc1bzrv885FysU9ODgyT2XYIu5EkcDM0Rbk/CzIhog8K9q0EhPyReOtr4jSMV1
4NGyb9jdAMeT1BQb40pXhobwZQYxvs3p8OOqKkfQUzIOwKLFzolyPY3WCVj7ubS+HuBBpIIxFBPK
z9Uxp5WPlQdj/mzTqgAUqXQMMO0B9/TZqNaZnjiRfcE+oAhr1XgmtdQ814Lyf1xch1BdafJmlxRw
JEJTNzXapMIHBu1dmCyY+pl/JrpM2k70a5QE8JWgu6vK5Blfynl6+emSTrInLdP03la+hHLzQcnH
TI8QN2ClpkSjIw4z8CO3vproeVijquXBu/D6k8wWjpsvrBiDz6IsHCHR15WvSzJkJ/tauw1YIpqa
kQSalGFVPy5ZDapF5R5piNElIxcop7XM2D04MtrD0M+Vxs4RIP1uH6Jl2VpbnVJMgrwi0U3poaKY
vtqKthN1uNTjWFkC/4eiG0z5P4E93t594Jx7h6T8oaTRBSoMI7ix/hHdt1tjkY1NqAdn0ceyeeHf
Zd99DFaDjL9dZ8P9IWCqZ9VvQs3e+MiMss88o9ZUf2J80KmE7IWk1ObUcDmImnJLg9LhQdi7tws4
nStsckl2pqsKnqy/EEeOE/XvnPBV9fog8pBXxOuJ9vNWLEX3rSMEC6CBmMaYjkM/RNSFg8QibNFl
sNudPwnA9aJqSNH1YTExgvzn5JAfTSfFErFNGOiGINs5vhsZXEpKNtyILa2ykgaC+38+dfOfu9MB
6XQfy/kcXFR9lk5CuC5zBFpBsLE8Py2bnOIbehk8B8UseYUAlQuCkjR/DpAnGz2TzRKGWCJHM1ne
pfA8WVfZusiIVGZCDsRUV9DOANXB9u1HZYVGCkGHooeeXbgJ5tEZRWDXojKAeiVZbb/aPoVgBlfb
3AVH/M83I+Fh/tLjF3v/m7yWjZnBs/7z40ENmdHjKPsKK2SudN5jdu8jZKg0z50TpU8duXgWmNa8
6NMkVUDbP2oVOLyx9Udep8WHWDd7ZwOzfnK9TaitSH0jnUdqdyarrBBiFUfL9twT593JaGaY0mZR
z3I3JFdC6rnrqIg8hPi2YSXz/LIIhXYOvYpHHBK28oMk05exeWKUSMWhgHA5vIlJftculvNzWeYJ
3BpE8ivGyvqQFepUqDmkpCdSjmuWqvJsnKHlYhTSKNZVYRoxlCUEdZydcegFRACrPDNIg779isaC
Gt3RrO/J+3AKOysIbUBJLRNWAw1ZWzM9X2Y6ccyBIqmluJBRrllheWEVknxG7YJLsCF+xG8zog6c
I36DA4xtzlVkuS5B6XugbOdFL43alpFh2LUkvC4KxqWqz0b6pHyavk+HuyC1uJWI2MvXubCxe216
MFL34Ce/D4zDPVd+bBnCEmxiHs2cViyBKdXtdz1dYwi/YaILHkn/8BFJtk10+gmGVimRCrGA8UTp
f43aZAUfxYuFNaEgw4rVXuNjwGMQkNTNW+JTnLgEO+HGlqztuDh7+mx1OH/H+3VmiwHz8GuA7gIb
qhsgJ/mPP297u//KW4P8DobVmBuFWdv7/9WGtY5jmnQUVNENQm/3/gVJqpCfbp/Qr0GXOjPK3zko
354vk9QZuFpmWWBGidrrnA04oY+uak/9dHTSqcfRle0cpoaycV76Z+Brl4B09LXDkhd8Llk77vse
NsQPxj0quuS1RVGWs8NWzsGjyngOixbWcAJRHR4RGHsVLIlhfSj7E06A3snGSB86Eb2gxmS9gdLG
5XVy7M9tBTth0yjAcF+RomSRDlohyVUtGJz3j1BEHnjHOB7RrUvFAEpiWg/GiQTMviJJMiZy2rrX
RHUV19UHIGLNEtgma0g+AH4BlfWc+3jMwsx6Z6zQ+joeJMKcb0CTn/CoapvPeF0bBtN7pW95c2yq
141pscwjgoIJGK/PQJ7X9Gp/sHDWTKrcpsnuBE/sDgJBYbnxEVFIfDI0pLulnYSPt20d5z3wOGTM
9pLtrwSvW0mAPSZovusvPcMvvmtow/jkfpSlKQY79oUOlQv8J2QRYWKW0OzhYp4tLWmxE8+zYSVT
VspNhArAUl7KOvhZvOkCOSeUokTrI5eJtreMkpPrz3BkavwRPE1d6nqKwKuZjQRS7czPBA7XEVFE
1dplm/d74yluik7WfldcJEulpU9YthAhnZwW38L88Sx1fVBgB4x9IuDARCDuHk9a0jIV1mkAB2b1
n2tD0GDadV9kt6MB/21mS0Cd2z0dNHOftpkCH8FsZLRHHElUqTHu4w0v79QSvR5Oh2umjBW9Calh
eP4Ja7IR4Lfa49ibFxwn907c5vGx+hByVU5t7V0XcpsFZQnGdLZr6Vws15gDK/xGNgrSNmByT4Gf
iDVrxZcgq57lG2/7W8lKpCHsPlZ0dx+41Pxgj3a9zbzNprrPzBpD5MvdKdxM3mnhnEU5DTqvyTls
/vocr2P2prsNGEmJOVLogrVppzFPQA/h+5+I9f3yE/AXhNYl1GSlz2jBjiOUJPHQCmm/YKprSkxK
jvOqVU6gY+dKLW7BBkWba+yEkRZU3MyrxezlYDI0CvKMaqKqmjzfzWuR+Y81Y/LzjN4glt28/JCa
kGlQJZSWrHkiJ0+X/7US6X0t0ZOrmNk66EdZkZkuRocAO6NWI0cE5tUj4TR9AhrIw0XVLsFb/MqZ
7hbntp6GZuPVsHUb+CQi9oMdk5ewBWNlMB/nCU6NeKB7P7FTTvs3Adz47kl01/vRflHues7bOx+y
ENT5Y5dMS7IsbEtykwWI+mPgNhSqfVL/8tNx42UUn47H4d28qd1hSF3XHOxXN//RilOS2z/7ItVC
SVVx6a0q8R/5C+3g/iKZHjweEjOXABcs+uk5k0fYthOC2pL6600erAYRjXzxvPt0kQudN/ksytSP
SDTbDmOQPsZxbONH6R9ZZGBP53+czyiewCi/sA+nLdPIrj0unJu00T2Qpjxe6VPeSqVqa2xm/Lv7
nV4QOE3sQpBGjNhbC99FeFTePPFNGskhTACqer42tMiR+yC0/32DB0XpPaLxYzFBZVRQOOb1indx
Jc3wnTZQ0hkawy17mSbkiaIKdeBaaTvjy8MxekcQqQdiHyA+TEWVbN1UpgoQcTiLFdmpjdNFYKgp
bX/x93ivvLX+C8KG/e+SMKfuqXOPcviQVzpKYxgNDi2Q0L2KeSOturm8yCV2ikwV0rCRDgyqZcPp
BLE5VPOEInSz7EzrOwAT8T6s2Xz76HZijQr/78dBcA4tGFXhbwjg/5vn3FA6KbwUFDEmg2SfH0zg
x7c7A3mWiz8B5PxaMBAko3Ey5HkJ9beYeHHzUSqsZowKSTN9pih9TSim/oph0W2kkf7FXmChrMl+
wnwydtFUlt70qxVbjBsAutGERBL3Z0ZC8ZF84NQUnyBKduBpLsWC1ymfu7DGJaw5tAfifNeLqrSs
eItKgdiBlTsTjLrhz9kQMlS9ppeO/DQv+sdENJUNC8qBs7nxqMnrlfkwyG0wEFKdycnFfovkL3qU
xlDYwbrQZLAO6N1Aod8AvbpmCqf362MOmGsjy1gr4k5MCOm27Aok2HY3Y77nqT00vDpEmchylYJp
f/74gnP3gG6e9cZAsFQmcbDWye0ShwDJXWr4LnELaXy8JiATmXxb+aHgnpnV+Hhfgv7ZhcB/ieQ/
dTNQJvEb9TbiIapV8F3yE3CemLXvxrQ3Y4uTQwtielpJlTE4Wve3HZWMLmgVau5vDug6tdxq28qM
sfVIeMXHeAEypTTJQ6BfAIoTajnLNN9I/6rIZHDBD+WZMzumDH7DN8MlxuSsNRsLsKPVZdZxwcr+
7QS6b0p+F2eTF1LHe1MUiOasL5vzOX3fhi+zfNfWrjLmUkBiSAu2o72lsLkubkEqkH37GZmArqSe
uIvVKGC7ElxOVCz06xKxtdiOBTZ5ZpKUE4gq+/Quf6wKd+k5/IZg2edvDhExIT4Z46inHjBVUhLj
JWx+w3synT5HFFs9oQgb1yGDMO9MM1jIjaSfa8ZQ40r5UTpXvrmQykmBdDW9VqUUQT1Bfk3AYRBp
D7cBrqtSY8mG6Ko0KpZqJ2oWIWMJ8kegJIOHLlUYeF67Z+uLqpXleIml+nAKTPxXgzREqlZplZoU
HbHYY+Fchajz/lFsozUXK/GBNGcRARNgY3b7j6bupAb4MP3ILf6/ToEPqGTf7hC94QYLDh/1p2VY
qhiOLmTwbaA9ayyOKc3NIsEttQTCo16gYMThnMz3A86NpH2v2r2FEqing7i7t8OI0DQ8Qc2li9qH
POYsqD0b9oWBf8pu8n5f24YdUNvt3K/epuWxyNfEj79wcf2vep3pW+hCz7GqJA4R+j8smxmNcU2J
JMlu0gYIgzV1NceqUmbiKp2kAqkpx8sEexlPf9RB2CkqkLUXYvJb4yqnTG+dnhfwi0RsSQ66xsgH
ze+0c7K+fclNGzOAJy3th9kxzSF4ouaXvMWU7P7MLqrPXyCxtk12pLLHTtF88LtN2pSPCCdJUJa/
+Ct8Te5ff8rBQDkThv6HQ2HrIn8vtObYDcRI1KWtHPZG4ldR6OwiyubsFAdoyk+ORzps1e2rkgGI
us2T2QiLTZK4OXSCJvzHzqfMO2EXl1s1y+5bwwj4LF0jieM2/dg9TpLauollB1suONQtF+MmzKRH
IsOvC1qf3volHTZtOt+NWI0XWT83bKcKFkrt7WftnS1712vZeqphEbUB+zwSVpew81Cj5ByRY8gv
Xy5Aoi/tlGzosJe3a8PX6V8MBdFQBXeMsYyV0dyW4ugYmDJ16jQJCECVogwvKIfAg4wZmspNfbwX
qLjz9MUIl5LIdjbiQBDUXD1AjvZTZoRowy9WiKy5DmVgUqTBmHCJ/ZNbCKu1NgbzfAPORhlswpRP
cH9o9Y6mCSh9evJPNCNdymMlg+OQTc97UKJ/KmDHQGojuh9QiiVSzIJLTDpMAQq5SJGs4XpXLunq
pQQqWOD9dooKu++AaoEMB5eeokweTiYMERKQn9DXIQfLHUhSIiKCkNs1ghJWmWGU/5lcWsTRz5Qg
GPX0hBY6qCz+KcpIjQgQkUYgViBE1i3StbHkZeStsB8/Z481Njrg6wVlagq01rsh0r91BSNBN7UE
uRZCa4lnSKZ+aBe4CoAuVJZrNlqG/0Pb1DB9Lvvu6SCu53YfGRNoj4KgdU2vrKtozo1aiXEAKV/g
XjsyNotBFslrQy0JQNM8lAhPOLWKxNeLlI5YWJ1USgiXM/Ylgi0W5UEIwU7Y2D5kEKvTciSNUrQy
rRPOHqfOgI3FsuQw7eMg/fk2f0oNrl5KbppXXFbjTlbMb5YxpzjQiONUkSgPNl93YfPX1MUPITiC
VCgosTz4Bj2jGVEfY+ZCwfcsarKWK9UvJ5WSD5xeH5eRbfcvDGRcjNGtWssD2mJR09lExOHFkafG
BsQRY9C+7iXsU1ysxEHhk8oNEVahJ/2japAGfhatyJok/mAzJgxLe+98YB06XKpGBbDJZge0ovYu
RdhYRg69GUu0zil9SQShEkXwthvXvgjA0fovvDygknnQZ8Imi4vbn7Y0s/eNO3P1MUdlhx11jnAZ
GqYOHi1WFxFFoVrbuz+6sIBDY5i76XS8BTHMoGKEoGAQRaPJtq2XPvA3hioclDfhHAxBnmBYnaWW
8Z+O3jKtwbPWMMWDYHpkTdmWI3y+5WzCGNJQO+D7IQmCgCaPHMHTr+6emngwr7p4WtwJllkMNg+c
+ns66IsemL2m6eskup9+0q8/VlZcKMOFnVXkCWGZvdKe0ttEDb+QijRG1pvrBxeH9v6K5ie4gVVs
5vrT/jYTKqKS4MQH2d/O6w4X2zY6x147H8+xW/sMV6CgRfCtUJVpeoCdWPrD1OZTIq511A7Sp4pj
rUy6U51qBr3vTTRspW5nYW+Ytux8c8iXf7L3N6MZc0zNBNCxkjEb5vm8M43IWaTcgCPlF4Tw534K
Ifq6TAAjUREjrK3CwG38r7o+4q4gLlwBIQh8sG5I76ytLX8TdW51MbuwkO8cHAAK2u4GPzB59XAv
Gxv/dY7j+Vrs2qq5tfhaHxjDtOjxcFSp3a7Mzo8eMuIKKy1mJepCdrxXjJ2hJ7EWhH30JqTqILAa
zHQopFpuHlUm6fJl1v3oXdyCrQ5/YmDY5F97gCL+ilcK25iXp4FI3QpeZxEd13ZSl7Kx1IhTfedg
xX+mrqbROcbU4kCaMs0Kwlw5yojyvrsrNtc69R6DGoOawp352eEdzEimBlMkNf74ucbj9SCjV2H1
ryotDvSD0FZCSBSBD40YrB+iJ6EA15/+yuZv8SRK6x0Vuq/0OxThZk81PGnVlorTTHNtsi/orZXl
gEda20s9/wG9Az8USJibc1WdY4AYwqAGaX4Fr7gtoYCIAEQ2HBg8nWMvvSjn8fUgXvz5JeSbFjmp
leQrQj5fJ8Ia/q0AF6QrV+lE/15v7I3axKuI7OQPPYFhrziLazMTA5eIkPg9G4rbklBPXQKhvVxm
8gUxn8XPe+OTkmiiHKywiuvBvHOsxnvbfuzI4C53xTUovwO4Zpr35WfiGrezt/OEhp8aFGsDcJGw
jhvM3Vzr0pT4/mM8ektf6yUyEdYVH2L641gwHSdOuRojE2T65ZRs5rQJ8jaUMqhdn0tORUmVV5eJ
lragPBnuoyvdr524G81bdPuL2gqz7gxe6AE7hHFmC4jmt/jCTfUlpt+sXr03ZPhXDJwxLSdk+XyA
Gk40HsPkE18C00dT+ePMkJOB0hoRVa1oAVw6zJOWql9cITWegsRPuE3mDQzDdidQ2u/Uxx3xpbJI
XLoDYby8NncErBlD8MTXmThmdtneWJowNqGtDQq3ZGPDyk1pSnGJquyLqOPvSfXedzhlPnvBpO0Q
/yi34kxy0IkQQUuz2+nqVnve6eXfS9TY0/QnqCqIPwS+qAMEHkhT4jsvu74130+ZkA9FwKELgq34
ohzlgBYrBlIObpJs3z5kb1bPQZNjudLKxluoIuZ6V9V7b0pSBQQFm7u+mPq2PoI+wjR8+SRGfOrk
2Jl7frY/PLzie0CO3eCdtvAR2TlPwRA5TwiXY/OIiatvjLe9+7xcuG0GTVGOet3YjBr1dDNo8Nbi
pGc559a48pG3Vq0Ftf7uQ0ahbQ6Gwelkz6i9vPwtnXyk7QHvehSyoLY16uwhUvCY3mjrTtCFi+tX
CiGI9K8pcNikr1aplfRXzzf0rKFXreGmjDd7CxAnOk1CGRHD61LyrIP7LknfNwwBPV/k0/Ky3tvV
ob2wafn0ctkNyG39ltnuckT/3M0LextWpbTYTALqM9Uj0f5YB4xoT6420RF7pZ8a82r0JXJA8n3q
9DGSiaXVlGOmrqn1VEDGWG06bfH3zBscKYNfeWrw8ddexjY7SsAPaSYT0tgGhDc9TWrH7mJTIQrh
WDux0Lt6fN4vq9jJe/ORC14fLsc9DNXwQfBU/ihGx+oKPJAijyjGyDcvH1xawwHwYpmWo2Uy19S4
HbsRfKH5xR9pliy+p67yq98mobnICoR9shMjylYAuBGzC1ngD4hGDmnRUD197kecW5yXdXG7zjzF
Pr0fmA73zCKHIqJZsm3co+BapC46HVM0yBB5O7i9+C3uS7BPTwobfoiuIrOUm2lN/OBpb5wvPrNn
FHjQAofgVSNDW1RmhIO6CXs3Zsix0dLcYC662EwuZzqy6MmciBNNnwoJjoZ1bEVDU8IJH+ci3uw3
uWnwK8UibaRH/c7RwlVUrSyyRWiDtlCQy8pyTfObr5WwxGOj/+WcNtMWmnXMs06QlkPsnH3fShxu
/mGDJcM+FevnjZ/xJB931dox1XVbPomGnbDrApTgwi5Oy/IUzIIMeLKyaq/+QaIOFi45NKnCoXCE
4zTN4ASQwTmQ3zUim51An5P1EBoaGxZsyAT6aKgSZpd0LPQ6CHvlDM4gRIhFxiT4ZAmGs+P2G4jI
Sg6bqfVZQwZPq5YfOsM3xnigqbop0g3w82KPx3q1pcAGRhdUpLy3RClJtSHSUeFMrs7Sb4/Xi+0G
y+TgbFPNNLtPOK+ZCDuRN7vD32Gqtvd5jZsv3R1fKg16K9haL2KRLjL+ua/+l/Jf+XWlON5bN/hx
6DNakg4WjaGnUvntMOMUHmU2MvU0DktFGKz6PpXesGQgRGyN0hVh+W7LXboE4o7Q9AIZtgHrqfTp
Yn0PZIabe+dJlIP/XGG/HP6vLle/kEb2Z96VLlSNfMpfXe6P1GjL0Ukzqlx7nauM+wck/0KRgNUN
Cq/PUVr7MrDjPd/rjiFIyh3tRg4hV0GTfOqgsqlS4BFRcer3b9cxnijsP/oQ4rClDhYb3y7n4ivQ
9a9eshxoPcO5a1URyoWGAW3niiAWnpqWlmCI+KlPx6TP/mOzm6qcUmMUZ0yRFoeUOfmkncudqfDt
6D+opcl66mFd/KeKdeL4byDDfSCogxM09Qpu/sjwVFqPGy9sA0xePu/dlJ2K05w6zTSCb7ZTrGMX
mHrzdaxvijuWKizL9dj1rK8AFAr+P4XC0DFdDfFYSTHT5I8xFa8vbaa0PorTQ6jP34FnY4RvboK/
rlpyuKqZBA3JFNi3wde4z5tN27s0Wjqqnr0oVuFeW6wT2W/s6eAuM+gsV2AkHSRYdUC1rr5Y5Wkv
KJAR+x1kLzlkDhzipD1J/DHl9G8orhBZAZn9KflxKWEKjBQB3oyWM7aGsum2heHSqBFaBNqFbLVX
cyoZ3y+2GPxSEapWIs5pA4mJwGUBHx9WpCoy27w+mhHcfz66JJnGcqcSQ3Zn2wrfXqjRGunCH2O5
InTCy+5o9+HW+omAg5BLRlvKy3v8ZI5yzhpZq9I4q2FYXnt47+pqqAPaE+T7H8GLdRgtOhcB841s
LeCnYf+Nc8v+iYQCoPKQRl0HGybcxhIsf5DpOP2ruEHT2d61aH/1xsPrRz4DFOMN+FhLvgo8UKxJ
yFAcV3zuSbEWXHRT1nP5xRdc8aWsJu6BdLb135P6TAdOdYDc9xQjKE9X878aNfokYRfD8S4T7znn
xd5yEPPIM1g1aKXlVvlNnTWxOVjp62RAhmPorq+OWEJBMGhYGmiZQwmtjLaayXJ2AfHPO+sYlgjz
qm1RbqMFiXy26HU2bYYJYRx/J1KNoNdz3CQsuHdV9TTn9GboNRomsLNra9xsdLJ0YkIYCSVPMWSe
G7o+DW0VCTm3HZLqPZFYKYml+WRhoT3Le3ksDpqaOJSpF/QLiIToHbMYmMqZDkbQgvPZnyFOF5oY
MBuVUqEOgNzUZphUnWV+tSAHdh/ahXYfMhv9hFZxfqA78KjxMvWe/pI8ofIogey38JWcFMRXvOgj
UN6+RlZmN7IAgQ1+QBi+Vbk5wuWW2uLBEYb3YG8Xa/+qMR1oVQn0i6gpJcbCGAPMMjmRRgwMBco0
aYlzhe4np1ecs90/k83EEE/VI5OrB3OIVjOWlPMkL6oFgOD2N8DAU3ysqD7/TaIR7oG0DDWF4lmt
cM3ZX5fNm4ugp3Vgov695+H5liFzw5c4yOpELANmJ3j88+pDGtCPPnpX8I4j5WeS9dimjeO0soZR
mYAwTlSEW9QS+gThvP1gMbGF4lqJ7CMuECpXJtVZwF5ZwaTMIJGNdcMO6c3OgAzU56sY9mm1uuMu
WPsMKv2FHfXxjk1AKMLuno4qF2BUUNri4Uuu8tHzgY/37glAZkg5y0lix2e2U4LdlSLtNXRMu76l
BjxbEf82g58MuY4wdi/gp2jv9/3o1qx2vVHcTFh9un0u4PHjzLfgKr0c4gXmyUiWnYHbiMvNv5g7
n1RLnFuOoqahRnTI52J6S7d8L2kqr1qRO82U575VQcR9nB/4wkrHGhT7gJaYbQn86gU1beApdq3W
pEILX3AgqizD5I3thg6culNIDmcbSWHB6BeZk8xHj3rJ4/OvPCfj1C6XGGmvAqsHs1+9AX7Kglgu
Xc+ySEraVN6UPgJqsh+SboAGzFyoVKGOnicx9rGmn5VgltHlUh3h7/kbvLHt3zNnMQQiN2WStnfX
N57op+X52LTqaMZ4tkh5E3WHG5jka7HzIccal5Gbyfhyw+xTJyjK8ZZ+bhLXt3fiLRaHIH17nF29
ptsM6LZoH3eQ44NTEpG4by8ceqIJvy5mhNYtAn0vYhqdhEeo28V5KqUoH1ct5llYS1gzQDXzjgJF
AO8SHwg4TmBTGHoP4Y7hIFbPfVCVpt3IN7xxoO6y0/csLEdv3xEmdK52iSIzk85FLUDiqnl0O479
DFw9OANSvW528YqG3vOHkma2L2CgVjTT8KPQPL8SQZtYuMHTLoYOos7nyL8EdWLbce7Dltd48dP9
BB8f/pO8Lgp71gXP+IOn1bOxKuwwy8EswFjeodc+1XtEn9EUVd9uGOV8f2GnVxvtsIV4U5hrC9KN
LSCZnJJ3koAzuuSm7bcFOqDA++O2pLDvngt4HYGyWEjZ9Zu5UGL1ihuQ5m46Sl7fkfzO21xnFuKS
Mr4p0sXJayhFM572rGyTcGxM5aREiw8RaaO9JdZ8m7Txkmeo+1UQnjX342q46lJb7aTi2cnXZ+/+
JhxkehQ7lwkV1n/gTcZ+z5f7X5bAtDOuWnv7wR/SBqpALlu2rRoWXiyDWODFLVBEkko4gqvCpN25
5UdDLACyavpdaEQhe14J6lnGuMV25Y8IVI+h6bP+r3FQLh2wr2LvV57b8eFC/dtEw/7n62vUMts5
13fRqR8qspnbTKxN3q2g2uESoa2zGfE3uUnvxw8fqNlsB7iww8Gymm8BXGQJv+H/8EfH8g7/PhQH
wbN2yGdGPSGfaI/3rMy6Bnb8JruQBFEUeHJb7sITE0ePFPpalWDQerXQkQOPhR0NY4okqk632nYJ
iFOxZ5ADuNnYDG8m3KiruoTsTnsKqnJQYIg15cKqan+6PHiRNojwtV5sMOW42bTDv0+thml98cxa
80uCjVIpoXqrPt4FBPmhX07wQPJKcxW3roqxHSxzjN7pNkSZW10JgqwNnJNDKMRA8bCLqjbyHPRY
kHTUQAt3E8N3UIZat4glxrbqbMp5Omy6e2FVcxQbZqbOMh1G/ZNdkSAD3NHvYlGoyz+M61zu3tTG
a92Ol3hwKXdryumdLpcBVwp7bVuwwjjetHIDtvE0YrXjMxSRgdPzXGLVsY8cme0Y0QibZctnia5l
zU6wVB609TfRyaXPtUA2mer6KoieUARon4R/yvwHdrybjrlsq6Wxty1Vnc9UVDRH0MQ/adeGQqHm
zCLXMoVWvue40VmlXZMvPgClCmHlliU8i28X1yBFi7zeCO8/6LO93E/UPeqzeQA2W9oPOdjeFivc
xjFH8833Go7cNSH39ujg7rH6GXRb8yBnlqRJ0sl8dfGeue1k4F6QkWaD1RqW3csxOSnl41N0EDn6
mB9uzWC3NCC601qKaoUpV7Vu8xlTxMYhpq2aAaEuA1cvMtOj17zu6MapPYNCN6QvMR9NvoCslrbX
Vs/rkZ0Ly6sA1lY5SzWkUEnUErgVwXu2E0JbqqYU7rj2RjKktr/uprc1yyRUPXB/k0vtNJK/harL
2d8HzYctCzZP2ijOc7459riJ3Y8Y16/myFUoDdQYIQ0lksEnDVTsVAgFDiTctKsBCQIAidr88xdk
gO4K6f0lqecrMbiUN7XI6NQz1JuMJzPJqeoGbHCKt5vPL+2E4/D04HP1TZMQiCcjJVGaiutgmf8B
TG/9jnLeGDSIg9ckdE42E9dL23U8L23ISxdqSYa0n6Y5VHZDRGlxjjk16pqUAFPKbu9Q3P2mnOtV
LHi82pW5i0T8Y6ObD9ZJR2ABhkk32Kq2IeFZwF8nSqt7faig2J9AWataOi+3YMzQd4U/DecqYeaW
rUlqXJ0siWyOKXyaGhA4UfZcaIqKTt4Eo5yvv3OopuIIxavGqEKIWO+J7lWp19CNmqfgK26Tf94o
WKnc0ubAfpmCTYnaILTpONntY74nJAwuxPovsRf/sxVrliHpNTtMtdg0+zebAndTUOlbz6TY8nIi
ETSi/K4MgTGAWtHbR49eAoaweNdNnqG7CLPHvqCBMZy0Jbx55ZT0m6ht8kATtOi1w/njCEH6AbJZ
N93Ic+3IslQD41e8WwxZ9SoLdOskSJiKEmX3HepjztGWQ5qqSlzNNjDRDMEfDnUm4ZPTx/+IHUAv
D+ZyZBCvbPQp0nnqLk1nZrgCFNDVEN6kSCqBNI9uf/zr6dkjmhwJXLa/QcSnIKlPhyEKtgzzfzpO
vsFvc6rTMK/BDtcKhKkHwojTm4w6vcweOny2y9kiwjDTney8KUbhuvZpxPeBqCcjz5eltEQqX3EF
CRxAqlc6Jpw531ClWEHw8ieJ4mKznHv72qCJqNVTsOzwbxaMiLuT1aW5mJZ7QgnQ1N7nJoQM6Whs
GjnGjnk6KshLXxAvLD4+c7UBzLBQER9y6X6gK6QbvBGSn9MA4EcWardvnC2vUL3/6Mt181VsV/ry
Qp8/lUl7kRKdEDEQQl/AOoGqINpHJyHl4DTYJglAIk0vLeQU1v5dkMHVXpTgv9PBdtCPYs3DK8Mm
16oUX+aqa0ijelq2wYP7DvHC1x4fMhZ+rL1rr7SNYeBn3b1s75QlQCF2lLGhN6DIwCaQQxc+omqf
GdsB1kX6Iba1AMw68vojrziJa1WSiLRvxLJGyKHZJXax+G+E5h6sz1yw46Vvq/LLCPcZIcsOokpd
IXEw6z9RNcLMfU1LRgCqt5+nCl7JBLUzS4lyeP7FCRbEUaWfSKMzeOV7v6SAepfXy9sonhtREGrX
duhmg67ynhXwtsFt0bGwcspWk43lMVvbu4MVHay1JZu+Dry9Q8b//ZsJxfPshKiG0STAzyPqDPr4
sngYTDoOLPLpu4LoOmiNQlnnSWtKJsSkpJFIH1mscndDR2RrNJ+TJOB8BEv/9jFniWvwG+JGm03i
qf9Qwy041k6VTty4RdjLlmaqS8Y8nrs20Jv1SCLqNqMWqBd5DvFcYl2amGfGZlXw9Tu/aVdKGAGL
j4ZIF8fAbmde6UVvbq/3B4ym9nOIWTGWu7sU5OuoCeHQ0YUyHossEnte1dhJ5vZFaeC1nq2Bpdoh
c22i0gmO5Q1ZhvUSrIlLe/g7ZSC7IPUMVRrgkuN+tUbCK/bdhPlzk67GfHkP67WVSBsIsrmpYkYr
EAyDad4uTewNXxILNRJYWX1THPDlXCy7HBLVHjGiFFYD8jpxEnuwRHtv6ZJo62wNKe1H4lVGYvAL
vS0jIcJTs6CB/7p1DF55S5niKqZVVCxhAWGWUgJorwyp3n15k9hRL9w5CM0o/2dBs3kUYZ6z7dZl
EkbFM9NdjwTj413RC99iqWEpTFcKktpHmCVOxHZsaPinpNHCMsYcvzDiO/Oaegj/H1DL+bTPKpHm
HcEbZLg1bHfXZH37CoMQ3ZUZXH9xWMGNHyZt8b3zIMsAOyxQrowuEP/YFuEh9m1z+lmbcQCS4iZ9
GGL1CT7rqseNuIGmzYGB5wyourGEVYxLYaGJV47wZ499tKuyqWr2FpfwypO9oaVA83AcI5HThMsP
FvCICpNMhJuisn74avJ6RnAhQ5yfcGw8JtqNrBRUX1Es8fPUGYnpn1B7+yMzRg7dNPM5GLPUc3af
IBmtbaOxovBKlWtnhu8kPclOssJI5H/rcRQFWF6OdYuk5C4jPBoEXQTe2JbZNOcreP6XpJULESml
euT+0NFkLGlSVbA2+7Kzs9VYUmgGTa8I6puO574lxG8tY8zjpZpRJEB+sFErPp4ylWbBth50wKsj
sPFM82SUUmvfZs49TUpdzKB3Ftq2KQr2Rvq9VWHY2gfn+lJN4nAiTXEPBD6zk1CKKtIRrUQKyyaM
76hI5OvW8OaTUTmgjcFTu02Y8I0m3ws0NHyv5m12nH08u5w3O7FAlPYYhkazyhOKmMlnBes7yQhJ
uqMVoMWGxdnDlJR64fnaN5Bm/xCzMTocwjlLKMTzIqnrA8QCGQMECF27GcG/bUhK4rCBI8tEgfTd
P6KvO9HzD/ZzYtrFrhnnBHQf5SCK9yh64MtdNhIE0TYPr3xJKOdV5FTBQNqAtX6n7l4KfrabJDqV
zmGSPTsBE0aOHpMcs8BffLHAvLpEsoULrbWMnOOjLGo4ao4t6wQX7DYtHk0g7Pi+OcsCAmHm7RO9
zpWGghbWVO18ymHpRmwVqgE2VsSRd5bFjFg7Skyn9NUKTss9SUwL1FhcRiSkb8aYCEPNMwHNrNi1
O5Zw5F5agViFysoU1l1IwaQXKEb2aZHD6asI2Iix3a/oMswzr26fx/zfuOeLs1D8X+k7RGh265LH
jNdHrG/D3jO0ZXBxEC9vmz9IH9/inc2uS4KrfWYsPwSVWG5StmLn5uc7hpHMOOmjRDcyz3ZvteR9
pvWT6h40ZWXud54gmSzXgba6dDNZJ0XEhwlCslZRUCiv2oAXYg5r4rrAmVvNSPCj0pkI5wVNkOqb
+2QDI9GhPFhXn5R/H0vKWyXBrE2AsDkNKBsN7p7Z4ye76OAunM0Z33Ha267GvhfIXUhJuDx9ndr6
5foAYOHpGC/eS65LqP84WmjWjQTBE8F7ox3F7/ulp/dYQ3aeTgQ+ahdPNwM4/SWxmnswTThtRO2Q
799uNRlf4w43s5FwLG3NTrkxbj3jIbwvnLJwUepLnxKzTzQEWa7CJO4dllilCS7duj7UmO736nEp
44fXTltl4hwz7xMYW1CizRTbQm26TUlm1MxGLgfkGuURJXn0UcADKQXSt4tn4hsEa2i+5OKzw2Yc
NhxnUM1IfKoJpLyhCoYAfcTKskYMwSFBOzVLfd0doMtEWF3+jebF2wKlxRoN/5sO26H28pIgFRUg
OwAaoS1LoXsjRSEm5DLum2qXDG8GIIpdI0P+ZcrOIljm09IcszH7svcmaSXiyQxYNB40LcGQqRrq
URbQ8hgb0+gLGJZEFQM+iIUp9k8pGhwG+LjTdVKbp/Vet+gBDetaw62NVQGwUXc1kdUx3lI7mrLB
sGJKtcJ4TOteRol4D3E5QfMyZc5g69DFq7biNJXm98OOr1bOxY98CVoPQAJHnn6Ayw0IQXdLTpER
5lAnAsB6mesNc47l16TR76eo6LYi+Xdx1Hxf3t2nHeWlHAkSYV5/V5YpfDo7ZGwsSUYOWjatFUXv
LjrIzzn2yoCFT1g3/Am4VhNsVRPbl9hzQRb8fi+Ir1/vOzWHPtICoThUbUSJnrQS3DTJQNI2uIpM
6yMTzadZyDi2xFZq0ONN6ETTEUDtP70qTSYZa+7Uk+Epxhwn1PHshJuPeEmPBAbmkMAnJrKC3/OO
3K8BxD2dKQFnpPU8XsapqM22A0XxnS8KtfaO7ubvpNUzEow9QCoKcmNPcWVwNYXD0a+5ovsfQ9qI
igqGhaJchKYAlHEjq+wEw0G2pIM1nSQJQ+AFhC8z9eV5jT9gbASgEQu46iB8MBNRbCef5ppNtVHt
Z0YoanK+pbi33/SwcBMJnc0nRexrOwE3zhBNIhNHt6z0020lYqDWCJ0bln5VMYO3TqgvhIOHWO4C
cXS/pgvebWtIu64dXGoieZNo9jRoY6I8bpJzZdnKGoMe070cO1Ql6hMPLiFNG/nRfY+R1uzCWrYx
fFVrkxbSoBP0ld836F+jXm+QX1KQ8WtK3OTjPKkPpWNb/usiYgzCAZGrlTF+cTmIsx1O6tzs6vvr
LNrB//qhX2OZZ+IGspJkfSChzljPhzN8chAoSFWXzbMD6DwkyrUWyj5bWQzbdHmeQUk2pMlZsTVY
OqYAlqbFhFab74tpSg+z+lCdPmGLbeBR6vF8x5THZlL6iCW7Vh5YG44kF/Atr+DsydGoA315Aqzv
PJ+KLIYvF5z5m/o8wvZ1BAb6lgd8yZlTUOP4g9EKeTUmZYVIzD4EUqsEKnOXOw6eZbug+SuOh++a
C8QP2XL18juVh+Dy/j6a4/AYoh8i2zqtOQ6luTl08emmxlrUbcoF4roYl3qRGTiZGa/dxi5rhm8x
0SzvwtLCniTVEKK1QHzvFv0EAlOktQ7MP6/1FDxnlivyjjTGPWY+t0CqfzQgFN9LeXPVZlzroPua
o7+kIdNpUO/p0E9UnN8LiOBL9dQ0evLqjA+dS/cPOdyqDQOGX2+j2F9Zv4+sRO4fDMFbNxJEspUR
zh+pN0cr5CMpj17N0rzo5Jo7DfR3xmIVs/l3atMfBVvgbFGsmwax7U+Tx6RP91vO8DxprURk2vIM
6ggME2/TcBzB/jAvgHGA/xYPDcnbj5Zr+bHjh4NbZN7A5b2Tg405znTXGpWwBKMZ+wA3+3g/Usx2
IpsHVLpBKm8egzi+fttTa8MSmI94sIMWqGhMQVGGU7dQYXwoXqLtYWMuKc8dstGweKqUneasAtRW
RHzVeqJkZ7bj6sqmO+/3Z0YgyRrLbvHIdHXXkWqEbu9VIT6Rrj76Yuje4cRIZ5VTivre/SobGbUV
GmJGIj8elul8IBhq7XW4HTLQoTe0HpI3c92qnWZVx2JiFI+irlcFK6UhvtYVmTQqz9eOeoTTsgF6
jVvYG6kxfXqboANZmSGps3tVaA70wTco2nQJLs68au2M52rIj3ElEx711kvrD5GxtGZybNYGDhcR
nQPK62JB/TXsELq9hrw3djWR9YmXX6yQLD5Uir9XcJExDvxpTJ1kKXo0OKUOYMEDov7PIvfTYXtY
Pqe0x8zrA6DVF+Ow9Cw0g+LLZA943SKGAJzLPniUrkW/U6s+173KeDu0h47gQ57Vn8V+mC3iI+Kj
HuTHZhkHdNjjlIX5Xa7dDEE24kN04hqL1WSBUhq2hrGoOwB2H/olZh+4gACb9jLupDGSjEFxFsIQ
qk/BZ06YsF6Ao2R+IJwryEiCdxfKnwro7bpkOR8sPT9DYw2h8bUYWSZ/Wt4j05mwxYDGAFhr6Mtz
Y1QOGcU+THaAq+E+S1hEYxU+CF8VKAXk38mFSoUakNqb+jWOqcimudeOx3nhCYaMWT3NTHx633MY
LT+xIZDpC6RNoOx3p9ZFHhz3qysBcwpjZjdJjuM2ghDqsPm9a9ROnNIU2YX0GziYtjJ5KWrNIcpl
me57WrWmGTIzPjt9R6qO1xt4U4gfdrfRcgD1rXi1WoOrlIe46bLM6w1nPgR990KXGt897hLjRpka
h5/JeoB1CqGXxRmn0t20B+BumdKGXIRnlfta74zdD/rkN8cGuzWQcoWbvRH58D+U8evWQDYUr9jg
MxuPMIgWTjqzlcr746o5rhKQLHkCsx2ZqUWcxmeDnW9FBsU6pvLqudm8jPD4q6ssXcT9FU4GWoRT
kWyyEaZ8Hjx2xReGNPX2e0ycM3PIjOAfHZ1eTg/BNGvq8aEfBiT5L+j+eEKp+/NUQ5fSMJQanYa4
1EEoonFt1Ck0wMtVS4oGYY1Du6PLgoN23iM2HU5WR6b6l08kKJ0dM5ekN9MMT5aTyIp05UhI7p+g
3LetMSwbdBDN6B8cbb7Qwq1eZhQdEBJlNEtdndC3qmrdimc98Cjw1Q3eCoojGfML+kgpvpmvvTyN
gEMndXtRydh/LXbu/c5DlQ9Rgwhq68PtktCC0Es3JrHrrtp/xwO7ROKDFeHT5qZkqt9hKsX/oBPB
J7c2wIgS0wpwUsJS64iHvABGbyftDxXw+sdW/AmGfWrV3nb7r9/5uKNA31w27hvS++N47EQCF+qv
oNoBH77sJ5PGbXoM+C+Wo2t9W2GK5y+Rvea8JzjHMe+oDrq4iO0L9niKDMds2lBPcf1OmLZa1pLt
/RKKFcsHxK9UaXq+HOf3ko9jSNSCyivV/ECTNXNbR6KJugbuHAcdU7W/8uw9r3x/LeewY/Oylksf
1QMMTb2wXpYM1P/1Ce3iG8xBU6CidUQviHGXECcJ+L9LqK6a2+I+W6QYUNE4e3O+NuX6Zuf+H8lW
oHC6iPdG1lTzrTz01cA5o1kDFC9xYFw2LZ3KxmDRpCfWDbPL/r678B3a7qGdLnRm4+Yb5clI/omN
vxRwRl+DiZZs0Ob7QHsw7cUXPcv53ymvOraGyTerAiwQKN90+1bnUB8VHHU0rwY674Oyh7vvLGr9
pRYIRnbWOSbCg+exU3FY7BT2IcqqSS5PR/xjMmfI1TnXtqdCPiBsmq1W5YHqVtft6gsZc6RIG3Fd
qAHVWHH8JmgpFNBSGogAGMH0oPF5lzkjGcAfixBs1X3PNib0IdV+AU5A+wdIXblCchKqm/Q0KbIh
iEnEdyrzt2ll9Z8DTdb/jXiyyH8E0c5IozYs4L3qCROKFC2zIkHoifdQvlNc4OLfOO9McZ+dNB2O
yaZiiH/UwVKgxLJMxD6CRIzEcaeQpb0Hml3wAhIg1tkzRo0AX+aMKWaCK04LPPrCG9fCq7g51RkE
MYWdUN1dQHgTiwFoTcfK17HEN5LQiM0EyYsKkK8XB352ioBsn9KCxRPrW+0+Ipl5/isAgN2Sr2I6
ieChcP/yZI7XJnsUA470Bt6nmWMqar1NeVISlJFAlZ47sx631TJPddVU407JRpbdkJJMhwUfJVos
0cdlDuCK6MGSb1RqL5eQW8Om1zVPtUjmDhYt1a0p5v4tE0q4XJ2anuQuj4IVzzgA/9RkGuz5GJUb
+1vju48GFhOiCh3tXtKhy6NxBEIZOtjYe1cMMV5zZPHAxXUwrdVHL3AxpRdjgwgo2XXXFdf0+7dJ
GH28siOhFLSblVyubX7t2ioU6KNgWnx/C+vAugWl4AjSfPuD8AZ5+O9oYvRU16hgDjd99mgHl5+z
mVmSQBuHu7kM4tDBDVndNvpbdzlxjNCXNgXMrvbXMnbh823C6n2r0HgZdZSEPiCGmCEpabfD7N39
LdAsTVClkTfvjv9qZlzRhGl7hKYtQI5ilbeLGg4F15sdjckhO/mwp+mSUugKVBKlAY1OUkFH7N0/
+0MbQVjCcna3bm1L1kv8WlSc3sD48gZAVOreNSfFDenQCtKxAOpQIn7YXiQ3GfunptcYMQ9GyvpX
78H8hEofbdfh0pC+lSpE488ZtZIaT1eahW8BOh+0PDKAc6gUdarljFuu9ixjil0ykBPggbfbHhvl
HrQVb9SMFNnCa0V2gPFApEa9jmF2ighIeeWI60EagP3vSQJdJyZYiel/B4GtQY/Vncbhkr5s67SY
r6+64grQUyoMDmCWvUfhW5V58saWQTmXD3U0g0GE+pZGVLiTx0rWrAXm4MuHxdwKo9AQXR4Qxhka
e2zF5mJ03Fu4ZzMOiK2K8fzrvMKcFUjTs+Blfzfx8TjYKAz16YjKGqFTf2CIzZUhZh/1kKKPmj+9
atAAJ68yH2qHBkm+xOloT7+m2LolobJDzLzxFG7oKH/F843tb+Smrma2Bg5vZBE32VKkqT486yqz
Vcy35TomET9+iuCf+g3e4dLIBB5cnrVgaHuhHhqZBTVAdVj7orduXCrUeebq/EMwjnU3hRcIrqcL
7fTfYBnUkuf6RCr85yAO7UaJOkzuSTSLOQ39W5U+C6kDShveRbho8KGKmBP934K/3no7++Cum6Ud
mKBCshiinxgIxoTaiJZ6zjP21RH7iq9Y0m9vfnPjmrOq8oOqDiRLtHf0mgLWI8ib/kVqMsYzJq9+
1T/pxrujkUjXh5ifxsLDmpy3qLFmqTYfIrTK5aEn7/W3ZW1uh283UMmlOxyNEt9bgPcEd4wAgGjW
XjCELrwz6d62QkLPtGgXATbiCvZGyBF53BXnJLBz542HL1nHaEjmJW+xvJ33h29yRXnfN0mMRE83
jgyhYer2t/VNql09sl9vPReIgIS1vUb9ocADipqIWvBz7x6WSINNOCyYWYk/GKEukD9Tznt2LK+D
sbNBBhiKF7UNXo+WmoKkYTMScFOGdiFSi8JI9Qdfmjzyi5TWCUknH/iRVMx+TL9DVVpOvDScbiQ5
SbnH8SJt/9KJVWLKxvTbjDS5QSLHgnTRJpMbSNv8BAr0nCkvHbo5h8+uICze6DaA/9khb2I/MWbp
noW1JexfIfO1wQuwvGHV4P/PVv34Z0w95QaoSpUVYaLuxzm6j4ARDAwez9XwJhovOvsC4ERthz9B
Txtmni7RUYAzJO6M2FLPu/Yyi2OUnTyuyKaoKKC8F4Yel2/hKgZ2KfRW439RuTqjdGaTOwX+Syy7
97jyqibFD707KTY0Z7kauHgHzk5ZqAOiyrx5Q1WH7JAah+dZzZlMk45fbijlXMd0LLZ7MtoRRA/n
jeS5hNEBkpe7m7LNb+z4OkeCiuz1KyLWZtQHr0XYFWMAQxbBVWdXCkUM6RmdbbCPateZoT2ifsCP
6fsAffnrsYddWYBZd0eXbjgp3INSp7+DlB0HXupdmBssC/eWh/atrIDvNKTVoLC2AE15XNVEfGzV
d8aTytesfzPzMXF48DEbgobq8akchylnbdxtJyNzlRz+DYWYFE2tPJw1dfikLqiub7h5XzMLSPfq
XeNC6WPu92qMZ603DaymrTJXj3dnocvltbULwsoxKrDTxslnTQN3I/PuCCMaWvbaSFYr3OzyIfN9
j966X+X4vRYy0DPEcfOGAALIPbwYHmjBdfL1CQaos57Mz/nSmt/Yn7OVR8PRH4bhIJ3tDUX8ZjM8
q4xmXlsL5HPm3lZpnwmTb7hCpPVjhtHeYcP3IN2gb2XO2HkUabUjXUoBo/+QY5R3nr4XyYerk7m3
pG6kLqmKW1OSvybwMah3c75h+gf64gkBw3WYZ5E716r1EJSACEV6Ntdd5djespzAmsoJ82LJXtDn
11IISBHtwxsgNqIA8m3umxR4Kd1KVuzY0gX/AA/8ydSCg0Rd9L+DAuC74i9NETmF+cUcoxAIMmns
Rm/ct28uCvHfa2vojDjnni4/GOvq3X+gztu/352hdR1tD3Pd9ZIg93thECllmM3g3TblGfd8cqRg
WlESilJ+QvvyiDTt5VpXbO+aCNZDGQSZJUIX67pMInfM9WfpQCF36TGbeqLJAjzauVhJo5Y5r850
k4YTfAC5i6ehSCzGo5l6Y3sPpzJmsK3nJ8EfNj7xlCMlhdVNAW5peFdTXAiYbsnKWjVYdkcE85hX
ESmN/QE5oeVDKF0ZzPMk+CuBTsM+bKzsTWCvkCD2Gy/HfgGr6TtqmYb17ynTDmqSFbRhvAF45dDK
M5fgVKIPxZE6BTKo5lD9BGabCP1fMIJ1oEinRH/fdfLn3C4q9XcH/rGYeEIxQh3cqUny09lwZ3FT
eOpwW9MgW7y7pGDwmBKK96D9gUH7GAzCDMoKH2a6xEfp7jpmd0DFuAdBCpa6cx7SQS9g9YxpYxu9
Y3wvsiBwhGtYFWPbdaUwXSiFIJW0p4Nmc7amUIAttWWzMSlv43Dl5JAlaJlk3zRsN0ZqFiFzwneX
fKPBCka6pXARHi2cZYwWvtKPBmELf4uRKg6n1c69F9IrHzsFZWov19qbWB+anE4LDthxvsj8hhlR
hNRlAhWI2v3nk9I0HNnmWi/rulngGS2lfrSIahW9BSNJvPIWVQzaPahzdNrz808bfGcsq/9ybGzv
bATyRuVvmy2F3bYwMXu385jyNEz2x6E4/APJHYwZNlk4Zo8yjUDJQnUViqAsKOiAlskeVgh6qK/n
THROoUoyM1As83H3AZj9QSBUrvTlwZyGiJkYc2j+DCcRjQke1Lduz2sXC6GtkjKPnGM7XT4BIz6+
AYAmYpuVub3Sml3vZU6GuNkGyc9ZiQD4i8bWB8QtR4H0RFl+6+J/cKicsU/8il/FfAGXWRFtiw26
DrStoMJkSKznXn2KvGygdOQvHaJyPTMQabzP7HwiXI0uRztfF9urdnhTOXvQMEAlQeHqf2Y3ksIZ
lI5ZKj0wbbpiqnqHe3sFYdX7UGiEd/CCWhKVz52e+nrufdYLiuX038l9/kEgN5UWdokYt93j+tVD
PJHgSk4PCM0aM0vrwLOLeQoVImaRznwkoVZlpMGoeU0NGaOOPdDuMQP94CfkfJo+xaPzSd8pdaEx
R1wkkI0BKHg7DZTHoTl/41SvONAOwh43JZDfnZx6ZOYf1BzyafrThK/gSffarj9S1rFx+oZF/vfP
9u2QO/8bTh8U+izXjmmNcEoJLvmymWxkl0f2Aey6E56vaoR7K+ksUSD1HGeg2FL+Sv6psEorIdvy
DQTvtisGew5XO6GC7sjOUP0Hp1Z5EmUM+e2uHGtAe3JXqpOQGOY9xd20aD4bEi5fV6a8FCNPXFRB
v/UJGi9QzmT30eGp1bLQCQj0cUlkcPA33pAGcpPjkvnSSTJsYNZHyfMKMBh8dTdISeDQd4gDxMVL
Hed45O1JNdgETU7yIocDod1n8OzbFhpZeJNP7OcZBYHHLkIKke9O7HlYtwbpGFiuGSsMCD69hofA
6d/AU8uoh8NTSnyDe6fikAFsPpmWcPN6Mc+ih+QcqntV+vv7DrBO5B/W2V3WpY0a4T/RyMi8ghbn
gTwaSjCKG/RXKNEwu/CEeAqqiCZbXiC1TRKoCC6n+vZM8XIUAshg4fmDE4n3Coqh5ueeIwp/kdp5
U1Aq/U4Xn/HvehNWxH/+1Fg0zcTL05FeO+QRZBUZ0OYCssjoz0r2LAY+88r1dCCNuA2twBsIn0vG
wPm9cXssIIN1JCXncrJHvuidvj/AneUjhx6wJBybfwcN8g+hmQ/XmiDO6jN8JxFTosQgWOZ7/BGQ
kJw4WOf46bz/JLGU668r728Rh42EffVMyP0U5VPtvwxLjkqLyulUgDqWt7Ew5oFSZivMtkUM032w
sd6TWoJaySOazi7an/ojZ+RAxydj4rizw0ZQSUV8IJ4+QjTuVZsGS7Q0/A9+l86j565pRaW4sSHm
N6MmnLgfYSGK5LmFzHPZEE7p0VK/HqXXy8KMAWrrhcpJY4JsNxBx+ZynfLZD+sAPnXLgsCBr+lhM
R+dgfy7dr9qQcNch4lRrKdSKuwZ2LOJAQmRmkdOoAwVE9kc/ALo2Y8I3cuP3R8q93pXtatSPmNaa
Wjne3/3npyA0GqDy3e/mr3h1G4htztQUCGYZJcowCpmOu9uXUDoXCgCAyfDRQXYy8TQAgQYqDP+/
RQU8d7M5+XC13OU9DcXyWMyKaY00mXkPqYtUCXttTTVr/lhexrg2nnkaCzFz1Zv/yM2kJQLJfvJM
MS71i7y6OJlotRIXX9t5XxdczhyrCHUotyYFoPPJUYqgdUveBTJxPlfAOXbRZVGW2jOptuT4shOp
X7XxZ8zt5iImPMMllc59Y9RYjg1+cJbE1iB9eBkVS5g3J4LJJmo6h3bKL5ehm60dzn8VHfUmLJlo
td/YKHYUakHis4NibajFVp8AWae84Y2EsgpozhhHV0DHhLeuUMyHRZVQ9LbzHQ5QYIPSGvv8Smr0
MJwBHOpwtgR/cchTLNUZsRe/52Ca+nyrPYpcBza8KJz22F+gCDYlmXI8c+3lhefKy5HLNzM3NgQq
a6zHJegfr+YQ0sq6nz/kL5jnPlzq8f2ShAgnKey+NA+nHH3seWGhLzqxov1WeRBDAg8mJT+tzbaF
Vllp3zMJqHRfa/SHZ0Vx4FIwW5WTUYYvrJEe5VwWPg20ummV4ncxueDSGRYsEz4aq4RIzgMQPemr
ZbazTkV+orLmhvIbrnb2codMSMT3LEQYKfb62jlKkT5fqESssZERNbF/c14I8ToQp8YKK6bq6w67
53A3iiOstq4AVB+djFF9I3cJosprMNuSV/ihVIYQvrAThng/hHiZxqaE5LsoeS/aKKkNN+gNohcy
WgW716nNEyvDfBOaCbNCqFWxvA0kpU1/8V/bAUGO4wrNpNeVH9ZRm4/bYpce5BHyqt1LdP0mZHOy
RWBHlSImwYSm4+F/iem7K4xw5MEdGmbLR9PqDq9A5ZItR127R4/xmUXxMzlPoWwaQY7ZeKqIlRZx
INj8BzlDih0+gN0Q6koKWacahvXqqf411Kmbj2Rn2cHp/ZBLidw3AKp8DPJ2J7En8OB5BvXvI1tE
hesVomdzzqEk/xYZDmftwi3oigiTC5SZmpQc5fcY80umRrSv7HnjzB7E+vRhag9/yHlrMQMQ5k/E
HYHS843nyp3UdEzifvl3oCsyO+QUZ5f3qi+gEvLR2DYklJ3qDmzZ9z2TX8sYS0ogln+O/y11VShm
YxfWz+4CCpb4+dlT0QPrOdAcJCPfAaeWVu1cd1AdAuMzpLWKK6yN7CphZSmDne+znjlWBpIhhvqN
L49+9+UlhshhjRZ3RIujYtV7v7hyneEC+rCHxRNXfuQP6+EPQUXhsjoul0gOY66GAhSqNFim0TGi
NYaj3CiH4aUxyzK0ukF6wy2TUeTQj/jwOzLJzq3hGhbZ31WjYKR00+2tGb5WzSNUbiOsA57GSJxa
twzyZRCGbtS3vWvQkWCkFOXZQb5SXW9bp4mAHFgxnycTR9ahRaqyYHJ6zO9MQaFo03UzSW7sf/aD
lN6GnFbkAw9TpmDmr2hdCURXxS4QBQpJiDl/m3B+VyEUWDuD/N/IPKjKoeicQKQfzL6CnHpV7Frz
BA1YMoJP43k092zf4Ht6Ua1SNkgApmlcLQO02Zv3fD25UXYxHDPIanG9lUdI39vDt7E4YrXsNK7I
4zsPqTBE7BA+D9R4anAFojFm1dTAY5qbYlSAtL/erPhuvz8H3M9929PxgIGJrPwI0qvY1lafDBMH
gJ45Wju4nXHf6bAttiUYFfI5QBnGUFYRnh+uXAYWDCPIstZ6Kik5MZSbh4y03svGwXTtZFxkwgME
YEMC7sb868+EB2EZuagkKs5npi+Z1c6O8+oVtYceNUGZ/9OT18rXMfI2Le8bo0UZGs79wrbUNZKs
8caJV9TcDe/W8bkzJWHOEJzBPYI9SGegOVapYO5I3JFd2YZkiicDr1+WyLMM0pw+E08nMzb2Kho5
g2yS5yMJm2qkxZW7S/2hcy9fDkUA67Vu+bJieFM85FlI49umcwGbhRQLSlNpTdMGGEGOyN3bbrC7
ttC8WfJhQDrp/1ja5ti7O4tCtO2miVypr3T+m4r3nKdS/qcs1VyEdavTWZh1IJwRhd1p+DC6z+eB
7LL1EWeozLwDiI5dHA+dh6YfTEKOkBGqvbNp21IS6wQdI+HHon2/pCuvrtglOMct3hcN99fjR73r
1J6G9JgYhf/oVd5CKAnPH6JC2wnSDw4HCDjk5Lftbg3Y2+0E0WaAhdhV05cnIBFLjUiyL0ysbmTf
ZNuphrNBkzEjJo7bfzyTk9LJt7KzeeOYjUomsveOns8DhLcXRnpglyUDJ5c51N+G6lNutCc4Yh3i
paJhmvA1jR/nVgA+2ad+FineqhipkpHuENjlLAZ77v+WmpLhWog8cW9URe+9boVkINdQgW0KrzNM
LkM/wizCUxYKIXy3cB4P1Z5K4jnq7wUWnxr5mIdOU1RO7PBOCio0kCVrK4P/MvjCWB71CbkroU+s
xZ6ywiYq7fVF/Bx1un0qkEnmoPMl4RngjbQGu+3iZanrrWvUiipfFs1PCu/RdFN/ACW9Qxr1vZwa
05OqF7FilgSMiy33gah96uF1uTxEf/y2tmW9SMsILUKrUJOBkT4VA4Whzca8ed2KnusNQw8IDQpS
IXsYjIJ1EnExaqWSyIiXYSqUKH46mbClV8I5YZZLSuZ3MEYFO0975iz5ksVJiMzPUPOR4EZXbBNP
aqXigMbzhuEWqpVzactT7HuTQ+GPX/WKi47vSND2/h7HKUB446nq1ntPgl6TGyPqoEk44zdZ4fcI
uNf9qvZBMba5/4J3apZ0PHgcYsUoyEm97GxGwlIDV9bx2N8o/dQ4z8LUdHw2tUlI64Ei8c5TKXD5
UBjw1d9xJMhE4JWgCNwRgKRPmt8TZ//BdTRPUAkMwac5AcjMCpuHr4+XqDBACGjoTUsMd3uVFDM0
4w8VltNEtgOuIw64mJFUuyo/Xx3DSJ8HFJ2j8qDqphe+7YLXbqEWp9UdksFVKcR7GlhCBkBHXcdq
9ZhMFFYhqx8BZwgsWEFp/17IJt5cCfD05jmMKoKbipVAqwLxX0NcT3g6SBikMFYBl2W3/bPtogjG
Aw9gyVFJwbt17S5v5nw/vjjC2YtiMafaPqxjD5dG9SqNt6xhQVm/uss5RwksEZcClBoxy8A6oai3
BG3dtLFTSfyCXserbkwQosQyn90K2dXOs2Z7wGQqInHM1Rrb3NAp/4ARhseDFo7SrmUTl654m9RM
0n9kKna29VS9YVtLDX94LCrF20D127c3dCVUAGreB7kSI+/CYWrKwKPYSOt7USj3yc/xmx3/IY2z
o9xQm7YJ2uqy9qGAIRXe1m3tfedUR7mRgZUDAHzTj2CgAyi//R7xbNj0XaLxz4TZrLYroNn2w3GP
Ia80V4VG8tNfxe7Ax3qbUQOuYfLbT6+adgnpK1xm6KTgweb/amsH+1DU7gFQ99dHJUR2RU3SbMfL
kweiPpTaXY4xmpD0Mv8cIOSxlevq5Gl0vSnmQQroZe4oPKi5nenHUEgrUAAXP0t8q20xhcUQ+eVq
oYxz4dfa2/uiHoRBX4DmCYnmE56dE3BONVIrmyCBsF1OkvA33rcYgl30dVGLMQ3a972nz/iJTsNZ
MFwAhMXVwDdk5tJAjcGtkVtM8O8uuWL+mWO19lGH6cWO5EbZW4dG5GYscTlPqrnXS4fBaBoydNHt
sI3YazTBlqPwEBf8da8f4udKNOqX27Vt1l5dNdekRuPvl9Qv7Itq8GGRNSErBE31F6RrcUQJq/PZ
rK0T1U/xAHam7KKZSLDUB9vTAn2kRIKdtgyEmo8AJtA0S5B2WOjzfpiMEHhYEuzdmWVliUg01yPS
2NY6q+Vch0Uw8Rag6DUKPWR4/MUgUGtrcXTk/s5V28Vmzw450lAJBZnx/C6mfSI7ZOauVtqjP+kO
9PHtn5UOJbN1MQAduUpz9qMdkrnrdC1kct/k3Sysfwh+1JlmnP0eTkvJAXON3Eyd4jEeDQIc0Jqr
uSSJjkJvXefLhgmBsLWrAvDXBZ66IEbVnAfL8PmfjbvnXBSHvHH9fLFaxAy2CivgB3Q02EQxLO7u
pYMK900u0UNMDp0Ix91CKIXYRaez6YY9WDUtCsJP06bbaTp76ft6xBA5BLXcGki2CkKiR6u8jRaE
eqQTAgn3/48yXdzSWjv2Atgfzd9nW0hQ5yTmm4OwdiTDM58CZGntMRkdT3IpjQ9VfRYWU9WHtNSs
m2Fns0ANQl2iOFmxBZIokta8qRqYwYCV+JZf+Z9L7AiY9tFYadIqK6SwSxrQHZ7prmLQbr91rNJw
F40pO+6FXMvt82IZ5JhiVvhUwhez90kbUvdP1E/EqtvltIVvkKPymIHInDSiIy9/NOI+XSK6Zje9
YSTjSXqPTUQcY/71xSaBqpkF6eA/tkQ3Ewp0ZBm3CD2hh6G8yQJf7xbOpyOYDaAN7EDy3IYaoKH6
Y0vJrQqJwuUsZHDWETGM8P90m5Kxca1nC0RK1yLqXnLYDi1wBSbUkrT/iTW5BMOWRD0peLER1N/E
Q16i2pxHGeBnIxZP6Oauxv6PfEhAaSkhJE1CwTkMk9XpwZiJvRkNSgvFLzLKmbtgu5MUrpsKHjqt
g6gbsA1uQrJepviNvlL2+jZ9Ckf0dF6bmdjZq5BzRrI4jCsrJSdOAeIHdqMhvMb7MFxo+KFY71sg
9qrbSMkgZywEHbRu5iKqE4nImSmWaRpByghe5Erqi5bmQRv6Tc55qXsuzEuEbydFffWpskNsNZf5
Q35lALsbJnCfthHHzk/wcM0tqBB4OaYxQoZK8EJgEGtx8TfVqlRn3fLplUGlAlyUcBvpL0Nyz0eH
hfvOUcXuBV0jHXta7mIgIFslBE1OvW+u/i+LlbDRVJK4HNFfsgn39cS7jvI0wOXT8oBSZzYcl2v4
5E3bT7GSLoG7NQBlRNQXlzm++Pn27cPrOoENkNVN+qNaq8YzS+PqLI2LWjhyYtPb6JKaZd/FwAk0
S50wzBjJrvzv62mdA8C8Axg3bjuUdVSmFqZq2KMW4IM8ozlqaEaQNnXPSWX/GDZXz51/xlu/oFiY
3XHcShmeSX17JWcmlEkd6KHk9hFdYz13edfwioEVhgHb7Z+tzPOB0wEK8C1yMlHD+pjyl8PD6O1q
G9HK3W4cp5QUBwgPznoB4rKtoSwenKjazoozGUlCJwIYmgTkDq3yUA+YFYb6d8Ehcm2ot1iO31N3
Jo+ZO1pFJ+eWpy3Glf9saBqbx5fdgV0NayyP2ww96bShq0IJGeVbisHvGwPfydMxQ0c2iaO3EWlP
gUq8k3pSMlbIH2pAtC5Nsh86OK3QPkeU0YEcTNOjNQMMfI2iPZxAeN5mBDnAHohHHOuecWsLvUkl
xqQwInJvSyike3htn9myTl8T9xIayP0TMXrauaxTWkxIquTiMvhjdv5r8bRi4qf1tOzgz9ssYpfz
VlTZjabZgd/mhVQNM5AhZI25CYSvGyrfF38kCVhK3JUHw9aj111qhdiplapDBPEK8KTcyw6V8uBM
HoUT/lHa0zct4cCGK40CEmp2vORs3l5drUn2EcHOLzaZ2oPj1lm5NUJLtm7abtVattI12PJB7Pao
PKjs39+i6RzEyB0QTBTz24zJfZ1t3xN6tEiPRtuZbtPWjvJa2k7YcF6FEUhiqDcyByOJfbi23pzb
Q1k7rbXcHjHkrFClxY3jWMJ8NBwWL7t7JhtgNAyQKasHeF0TJS8BVQiHUGGmIGTtLLIEaWinNHR/
LPOKuerI65UMOontXTE34VV6SFKCXhqpz0vQ2+dbvyr9p2DC+GNSzDZSRvTMAsyjxh+p0lXcaRxj
FBJpKq81qsycXHHrvTT70ZoFcyqq030hNDHWONqNmNUvhI0m88pkd9xJKh96NPHsothTDdlUCzYv
D4fXjdBeBa1GACTBeN8WEEkw1fnYy5rWwUrs0nKLcF72vZYluUCLL35MbViDM/Jtpm11R4c3NsBk
/RSasI5g8AYiV/dPLFg+znTIbHUOciKu1NeZyO6JHA6M5XqdsbPnBYs8SeytaDTb/A2ZBFXkYc3y
iyoSgy8twefWVsq2j2GWh1pIuleHh943be67YBLUZqtspADKAxE5NCaXP5gxAXaqg0HhPV31l0Dd
X9pcYxxH5yF0tDstdKn4vBM7P4fmwc2QLoi+DAN9e5CXtRYzvfYDGuZNWQMUBUc9HVHBXPEoL1II
JNISmg2BJERntVp4QIk85OEGIjfgGLXCSNZ83Yh3LiQDty+DBIxt8xmW79kic2fNv/dQlRiSmML7
fcFV9jH5d1so+ZbvlvtEZwLWGlzCgFmVzGIDVN9F2E/zLiENpcs4tRZtThDWSM7OFxRNVZa8Pd/2
jq0WuZtRyR7T/HAylCJwv7NRsL+mNre7WTMLj2bFkUvnVeULLxlFEafrFZQdrskAFhzt82AbNUas
BFO83UrTTPHEncnWnxeHfA+fURpl3d8Pw6eavnxp2+ynWGYyu320dhdyQ0+mlzasD2MRcDcJzO7Z
LbRoSwecb8Z0EKnAAjTvY4p9CM0BTQaElfrumSyxKEPscWktbYOC3hoRWz582AtWWV1sJ9iXCsJf
gFgLAq7hvy0PSr2cYUGOtwCZenasx1TIX0hCr9crlFuqVY6VCdOfsk7THgTeu9kpETJWr3QLl6Fj
9evJWfr4Zs9FBwW+/Tg7NTZwH9g+eEjyYiQZIwLlspcpZHvlRq3bTybjiWllQSwC/tZD8qVMqJ6H
6sObYNk2TAAETT2VfNgqlzFz8vwf7CqPpiRh7r4IxnnHm1bo8wCSIyhTk6osc49sN9b6O1ZqifCq
6yBwiO1qbgBDwfG4fv/BhvgMLCk9ZJvqdqI//z8kFrjRuqHCW2W266Wxn2bNXxxp7wkS/mOeDJDi
4UP4g+AZVxOcjaKfQ27cwMWOBPGzJ9TzeCFGs6jAGIe0xpOjj/dmyKmwh6xQSzHcoWqhEkcf38Ox
fdQyYeQJjj3z2g3kgkTPhNJniMWMLsPA4QQFiqbCEUvP5Nu3cU3qv4B6JeYywMMJchAJZe44kgRR
NAi/uzTqSx3zw/KynFBy8uKljN6x8C2E8ghV3vXnrnT8qtpLWbY6fp6OpkWgXuknKrIXCUlHeVGp
myIWvKfkJNVn4gfzuD54JIe49ngOqCAqaNv7TsD6ruxW0IoTtxG4AI/kqmXumFTuAmstdTyHVzNn
2oXTmY4jzdFdeHTPWME5oaD/5k1HvquSbJMUuBSOueTgn3VWnSC1U/d2od+hhWgt0g1mTcFh7ojP
UZP1pQu2iVoLIXjmi0zK1ksD7rKHcodPPNjQFYkzpU9ujAqqfe7lwcbnWYVwKV/K8ucS9ZISkKs/
0I/Nh6KcKf/ioVcs+xKTZOlDapXF3KdZbpRY0VU8+GUy+v9DIWQnP+1qMYnGcABTuO46o6JLgykj
l2NMdr/P63yfF55v3CsOAns5hywHWbtV+oPyPiplzvkHRftviNnmX/HqR+Kjai9tc/jOyWTpz1LK
zt+5p6Rr+2OGFhCIuqIHeH4pVNW/OpaOIaE73y4TGpSsOpb5Yvg9avfkMevL5upGpqHD2nze7vwo
zC4YlQUdDuQf5r4MCIrk67WfPZ31DmKJOypT4Vtiy8K0gbQB3vO9hGmRDzT1Lc0PA3q0hTZU6mWe
rMyX0gvXZeRNjMOCVqhohLKjbTx+SfjEVp0wK6iD2h7Lx+2fS121fKRRLN/3tduZM9iCkWAFz5y6
d8zgrBYlS07VPbEoZb/MxU6uDqNjDacq+pVvAfBzKygR4YTBBNe5FavXk2XfIayNB3gKj25dDVKa
2J4b3SrJc0FZuuCoMge8t7QN9UJ8taoiY9PbWnLE4FLuqPXrH4bWCedAAh73ustb9xS0vlWup9No
vGsne4VhHk+Kcxe4tJrDuBov1GYYaPytBaQLn5EqkX5zHApKxWakjyYi0yWg4l4BA8l2lOZoWDdX
LfRFxa6Z3Klf6igbkzuvo/cXwHt9VXpFkMid/sSQOx5witSkj2jLIRuQF7ZXN4wmqnYF6M/7ir4h
QG6Pb6/zJbcrR3wwZByys1BLxSRnIagYOBLrB/0cmjH4I722E/4Z/JkZM2y8NCmaJ/QfhTBXQf0J
tSDad4vv6yx4VLe+G98pGu5dPSlQH8nqoFlerwvaheMFzsVD1mzCwqRsFfxgNwnN9e0hCxAqAVVn
7i8kNpVdRCNZs79/piZMkicijx68fHAIoZGcWjwaYsTc08JobfWhx8dY5Id+iCjtmwTUmYu60wsn
GNIf4qdcr+8qG1JKtJEeyM6vnxNGWkiiKRGQS6GyFM7p1Qjp5kHssNxdCYGvVhHvHwVNlcI671gU
ImNiVGUn97DPdsqSErUrge7IrHbBG9HFKFs0PFqqs8uTiP2y3pZqQhPHfemGFOhwADVKV9ig/nK8
8CTcjxLsWh0gnVe/NNhVI2sHVxJ0uPSnR95Gk9k0KTJcR5500HJHOhEIl1/U1f07k+yH+ggcMmyS
ivUx15IdjcepSkFIm2UoHxcKwSSXXZ+tNLPh/SG8Geu9hHZIpqz4qEXj7bf7MvIctxnIlsn0pvIT
GCOrnERcRV/lQwFgXPE5WufTtP+rHdQoQp6Dn0D3bSt9gl63z9RzdId9Obs6kpV/VSfIjmiOsQSe
TBrMvbbsIK/+26RCYP61t1lT3m3iksGXMACEWy1r63sClDX+973rQywALJoUEpvD7MVRujg+a2YP
vTgs3XsdjhXNSxyde8rxcvRQFJQfFvGJrjBRUy/yzH2NuzvDndb1H2WdLhD0V9Ove8uP+1BRHi/U
eR27i8i+JE3qIsrNE5tgdKUf+16iT+eEC+aFY+s7FAuhdKpTHGuy2dp+m4qegjbNQwlkMQmZeGr5
wzEsjtcpbhOV4ZgmokTyrIRnDuK+CNOuGKoGMBAaLEeYW3s2wgLajTMPIQqv2DB8WzlIRBjfKwz6
GNOGgNyewe55GzzCToFCZ1mm/JN/zyDV/nu19n2JjZmeuM+LfOU72JgMloCuY2BkdyTtuNv8Wufr
UO+ZoEaEhN1ztZIvREmRXHB15mW3ZE62Es99euj1z5ZNcqEo7zfXx8EMReEraH5G32+fjbFGcOkf
JIfQWj6+0faMhZXMNa81nhCxgLmOdNQVGni2mRfiMm/JIFlxJzAU2AT2AxuxJud5Tc3/bVtmXZJD
adKHCLKX76QPojjJ/dOXcBKaHIbrPXaU98tBUYygR3Uv/0wmTwFZUFWoXCIZ3VD6O7wAysDIhC+F
v/q2jD6UtNpxQCaNhINtzzEC5xJlyr1LbLHc7SazmCjjJaazzf0NISW9NDuBY1MTd4HD22waUW4P
CDxuguic9+HAhFo62P+/2cjSjXWCow0u3UvXyifCOU6mwzV19cgR5ZegGvfeQGs1wpGYWzJ8/fVm
ofcayEHajOntFi+6XLblYqbod456ugXRHbVQ72El3r8mHhEfE2eEo82AlSATS4XKblE6ablGR+FS
y/IIH5U9bVKy7Fo8ilYEt/snunT/PVTsFftY4qCbO6vRZveGy285OztMUiiMepFpFbCaKSb6OeeC
WuIdZZRTWjOVeliHyN9+udxrQbZkdyto3QujolJxEYbJFaDoPn6UTci3qiNHGPfYH+dOg3DGGPcO
Qez6YvP/CgjUCMybq8UFz6Eb588E4H4t39sD4+yCsdrA4Ajjg2gDQd4Aj38BshFj1CukpkgbsFNC
i4jHv3k15jW5VVhLd2T916uXNmUA11lOC7Z/JmDOJv+f6wVttbV047BVObrkIqDdIT7c/hgzwDKk
OmnAw0BILvKXdxxuQ8ZKaCgX+pihX0GOTw6il0A1K9Mu3zV1AEVopQD6jfnXb8lk9JXdrFCvc5jK
wfgpDm4aMP8HgWDhEM/i7OQWYjvmqZX5KvGWYMIdxko+XAsXRiY7kY6DxAFH3+arB0RRBoVZ3+1Q
NTMpasFP/28GvaX99O6vzRl9hh38twjzP/7fSVcurQvaBHmibM/MrwQ7kDRyP4dTaXaNYQIanmhJ
021Gj13VT9O1v9tEJZ8RjQsTwcTrz6KafxdUGc8i9g1m78Uwh20nKTxDIuT6fofj9ehndVhUg/dc
J4HLSp76pAW0wlqsifmvGpsNO3eSUnSZhg+ZmnTyPpNOwtgHuoByzkqwZf/Ug04PuBxKUGQ2uWd7
v9KW/Bu5KG1hhBFz9G6HBh5vKRMUBNf7nIhn2DqS65lbmZ16zBS30V5g4fsHB/ZwpHU06lwxYpXT
Vh5Ynv0mJR6zcBPSx9EAFmBiWsPihp/d8/Gj57IEi0U7bDRQg2MGjoxYU3+Z63WLoTlWp+ec6atI
npJjw+XR/sqTVMKeVGaeK9CSkOQBhuMH5fpsH5MSvRVEIMRHD7NUE9jbt3yu74UXr8k9R3subDbQ
YiG9jQtV0jtTzMh1GfA0apUeSjD6doOxtKz8boexP671pNFOkwm5tZXIZFzXsarIvBbnJtCn78Rc
H/nGgDH/BrBGB4Iw7corpstGdWXowQIJG6ecOF0AmK5/J/DgG7y5GeMNTaU3bkuYhPIqwzYVjwsW
Z4fjlXxlMO0CZb94/StfQj0cffnt+1/QpiLscRSP47pONCyx8Qgz9dioAf9Qsy0YAO/aGX1xAu+G
wGaKhMdOw7RPkg1/TmteNVAL+g+sTjLbFMU5NowOYGxGpkf8ISSNmvR4vejIh31F9IFHMCaWVJn4
yzFXP0HSom9iS8FxXElyza684LtHy0q91fpPHpFatDWN4hk0++gL4yWtgAFoGLCx7zTOcFe2Yg6L
+Txf4Isue108uMntsSfWcdyoQhpqoKkZZrAFSZ+SlfLbKcFbLmIpb4phwbMoK80f9ucW+9U9TTtB
UnTo6iztLuf/yUAQ1xhELtrQPpcM9M7keSjf4pdgi0RymN8j9/zLOBA9A/0YaPlkAJJDCIx7Vwfu
DeaR0JmURGuNCtboIPBLQIlC+CLtQae2G5zq+uO4hW7KPH0ag6iMYW3jc+stx67YMVF8myCV1e5Q
Fm9Q73WT9KlXEOTXsyfdbPSI5xn3UY4gJCq2ptK5qp+q1Su+ZnNt5o01FEq0HKcUtgkuKXqW8l+m
P/69Kq8AM7TxgJATTbYENTdmiEE2P98MaH6ieAyrxGQRWDoStEMpsAiJvC3aQ0NinVb6zItRoW3F
OCo44xDf4CESBF9lBRH00DEwGBQeuOBtCSbaMghDuIlthttQ61LhYSTrPLYzmeUDXUM9NI1lPcjk
4gR/CGpcAlOMLJ6HGiSAaGZW7ApTquo1Cp3k/Q2VAl/NvwQ8LpHWVoRLu5b18NltZVhqt2W2rbtJ
ISAmrIA5b20/uPKSooSPVcLRiia+JFzO+UbtNqMsNTpB8m3SxOi97PXv0+Cil4DY0f7zpDvNNiGl
j1VG3jlXu6PeFLpZA+lv6Bogy3JZ8B0PMVf1aVh/x3yXx1jbDI8wHDbhzBU5XZVOpueIUH9tEbF0
YNC+0YjnWfTUeBEryOzMXOusyJxIiMFgmcvgFXn3f/pALS4/xWde28ZPzncGPdfHzRrRvIjSJZhE
sFYpUJgCkw0OLLhpBPVMDPYU3rOLVEha+TcK5GMHZkbG1NXzpbXKhlbXq9a9h6oTC7ie3FXwyYpi
H5giUV4STjrfeCuWLj40UlAZrXZjitpG3blmyjy4D5gTRdSk2MdaWvkdMsEgKPz5jTmk9nGk43+a
1XjVqJ4g9Qx3b4+8Bf7HwClW2RIZrdUozs/fuTL/Q4IbH7rQP8K99sx2GL4Kmg/uVaByXXUHE/5i
POVBnzZ+tqdgtAqMM15GRep42TwjV4eHMvu+3G2FhMM2JYviwDG8Zge1CafU6ECWzaW3MzRN9idv
D9aAZC186G1CK+y7u83sZ7bhYhBC+YdQck12oMTuujWoy1T7hQ5XPH+Mj6Qt5crfeJbM/0vZbWOM
uvoo90xy2UNXkUpn7Dpg6xvPDCeXzKBsLI54uSF6UkuBStt0hvoMyJEAyCwLgGII1gvJTBw7cWLA
N+vv7U9slAPqQkMON6WyTVmTE9+ampThHWR42Chyu9cXoHxDaNtxCJxOznaeOLlnjlTGIc8U7P/D
MIpd4q0LkMwwvwnh+cVHfWIkr0zfRbdi0hxTupeIPGdqz7S3QzT35fGDLU93Ef3PDFRYx1q+8CI9
Mb7VbzrSsgJ7iSz36OB0OOg60tEyrhZKHEyWg/OdpXFRXBDP5CX2e5djwoY1uwEv5dO/I+Qoc2ja
wSm0969Pb5tpU/2BRg9p5FzLjVYwI82pmN3xEVMvt+6MRSPD3F/Tj7ft4ketAwVZ8Y+zYRo0As+d
e9vqzFNbgvxuIZkPnEygZ8gfneTUnNyo3lMBg6EYn5gmK5WXp1DLNo2vNmgKjH9llUqiBav8cKRb
i3t09JOM45ploN+jxCHVmuZAznHazGlhByTcwk8YGFGSdHIDF3FCK83VWpvsNnbHPYwKmooO+1xc
xYZWExLmcP4rnm35jekbVgnwzW8R99L+5N76WmYvvAoeg5o+KL9zIDLFNg4siKVXotOyl9P7MJUA
lK81FMls0vTdih+J3bD6ImWgtCBr56jubBJCN8WY3HDsYOKDkT8wcwrCVx4+hjQ724rnnb5F5U3R
S1f3h3iHymuX15xK0ch98lbOHQLWQ9WyMLN57ULXA7AGUagvD3XYlApVdEzyUDHW8WW+xp4/oC79
PUOV60glCLw3vRY02zSxnMOZBNSwyjVTAIkhfbfTKz9TSlUrVTX05pUdD7uBxc1aY1I/q0HvyeX7
GbK7VGtlhRxb7ujaX00z/j9wIgIMVwJpy2VIZmGFyj7ZLVAQdQyW1EurvI/e5l4KLPLwmhF4dz4X
On8dD+L/j8qhwIcBxUkR/VnRcNKiuCpIRM0LErhkfpXEcUu3wU2DTJohRUoZwLjNz/iGqcpebPts
Y58ekop0bV2qe5XzkCMG4sFvE7/4qUEsNVUQIWIbQgsu9IsqIJDKIkvMVmzlwBal2Y2Jt+2LbFVp
Kms5QD4XD42jlvSrd89GJMUiA92aJX79EipfFgVK8wV+AOxaBPC87+ecUtK1+Al0UWbVZGn/a1N1
QL0ozX8SGJ/b9yN7XlhJsV28/9kiaBmLjvi2xnRO7eWTTd9ZILeOPpgGHz0NfMr+wyo+NerQaTwr
IjB8zQ8B4/PnH2EgKFGszljZhEJsMhM1nARiVtCY7zNq79Cto/DpazBKya38rnP9A6N3uU8LMwtH
Cec+yAzszwyRaC2Q1+CHghBWsUuBBtRDgDcIChdItNPChdNlQItF6WOteKbBC/98z2Dcf3/wnnUO
7cB7/P3Bj0ywsl4V4+zzSXG0yDQJM0zuLBd5EirWfdqV77lkiI28rPmYPq0XJZ/X4S/il+xwo1MW
rq4aaFPeIanPi6q9AfWTpAyjvNPHKLFV/HT6f3gXzt+gztWwQpj6Kog+6BfyWgfmSc834AR6QMDH
MK1w7ltKqZWVM1CXIffHZ4DdUrCXU6XYVSe5tkmY32fpqWbpCzdzcThHxYUTFHC4hF0dFFjkUjpe
fXk3lAuXynMQfMDGqh9wY3GF7kgtPxc8urN+BZJGixdbZ92MDVAJoRFfjwIun6DYoXIm0kbvpJ0G
WPJHKSm37czhfnRtwQ50KB+y15kV8HRfIfet+Fc2n6PV3Fqds7Cm2xjWtPQePcT/4X4QolNMuSOM
S1k3uMk6BKxPdYA9VEXTHEy6BOsOXhkukIOVlw3cKcUKkov71Ljnn3Nj13/nEaay4fmbArB18fWH
bOIS1/ZAM/I4vTw0z9A9VKxlEbD2rh6Hso0yj13ed5I2DJPD6l56Z1jEc9xJLvvVf6ND/SkKfdz5
UsFPFavUZgIXeIGUYpiAmjinjHxf0XUnXFxjy0KPflqtix51fjLN9LktCW1qTrP/mVRxZjNpWEG3
sAOV85491WBVfP3y+k90Yd7iynaWst9mi+J4J172k9+agO9tCCuJ0WtOjy0qLtGy1rmKWBOLPQIJ
ansNgeS5fZEpQahoNTTVKOqNz/HY+CtdAaziUZgO8kX+C/15dzSmzj3mv3cnKOHNgjOVIBYGZFmg
nq+0swek3P3X7M4I9C8C6XZrjE6LSvLfo+Lkqhr5DIcGrbpRUC+H6R2iYZiyuzfo4stIf3KT+T9m
W3MzqflE4qBrhazWj1zC0S5D1eZKUkbiDCjnkVqtAdrUSll0JqclbhLcORxnb7/U4CQExiCX0E34
oUfXOmE18qx/J+fuhswvOXXL+5mtlc65IeaWlB/JyM7WMO3q18wfryP6Z9bg4LxmtPYk476dFheP
nAapAx7vDBh5F/QCQ4q8oQSUmYynxlRkpUbKihDGkma0Lzm9jljV8HVDkr80R137ECYG347P4LIo
ZMdjcWQLaBi+X3jqKVMtaRIuYTbbapPGIh85/aHYngM/e921kkAGklQt/ah7a3QevWxcXFaF0ItZ
mFvlVz3FBq669QUsIvvJYoL5r37n9NZ2XEEghjIqgVUCX7cFL0D8hHhEWPaJ8ohe9w3zpNFf1Ltp
DnMB89x9s0gjycS440aw8LTnNlvlMcCqcXPKkMRyjCtg32m8NHCBJOlxc8dk3alGMxlejrlHU5VY
XYTnKc893H6EvZkuKY768upszJfZ5hkKPTid6N3k1uE+c7jePuOUZQN1MnGXNTDHIBZ5JnRFcCSp
BTtjhNJuI06Pmwf2Sw6b2puanZ6knGQxa6AIqn0NzK8owRLVS0A1ZWrxWhNMSxHcKb3Tp2fsydQN
R0YGoJFCi5cvsdrqpF/ZKvsd7aLfZ2Eyk8gEvy9GnjozB6o5zORNFBFkeSZz84Z8awjNaNzfDNI5
Yksjg7y9PDGwWyP+Wb4IZn7jwIpYcPCvusJY+uybE0xBcSeY06JWWj4Tgzhfuo446NK40/eUHURJ
sjKGyd2LdfAnQwnqXgQKdOlfCOpgF/VsKYoVxMWkLHkEKdg5F2LGy1UzfXgR118EsqPXV+HdAFjY
yHEqZE/ApAs2aAHRRu1TPhmmulkZ2yShrwlXxR0ORhnTHe9R0vMOtc8gJYW9ObbCWkSHzur/1R4F
VAUowzKpwZlfePdaDuPGPVvv6+pDJV0HGANj8yMJAweu29uhzOHyEOfBcdEe3tMwrkCTWetty89o
f/s0pWXRCgI17XCRRCRVqNnt5nMCoj6U311rFTLC7vFT2EXm+7VChfG7F/K+c3eZZih/VhBcYctR
mmtVCjoSAVZDtondlPH0/6CFsvyJp35ER/J4/Hl5WIygdllZFgw+/L83LgBkrVStOQQIg1Wsr4UY
2/HBmS5ZggR5JFd3Ok8bBpXCozgvSitLPydXWKtBsJYVUVsaHl+qsK5RBGr6mSOiI7TUcvPoDTOC
2LmtJXroyhjo+Z840xhJLovs7Wo1goIak6S9tvlO/j7o79tNPwG+cdqo2HtZsbDgPH+1ujQrT6xa
TJfY21a5kcaolQSzCxedHS6AvxzrygicMyhu+k2kLceDWm3XDyYznKhllIcZfqntgUzQDd+nbHF4
WvyQ40Eujxz1746KQhKGXhqET36jC25Wo09a/huzb92xBxFOq+Ybxd8bVFC00h21t6lmrqHtKPGa
3uQT6IGu3bTaxr5NhYrqmZ1Y0ruwKtmsLgkfh+s+anPKxfNKlpYhkpA6RIBxOHpbo0ue9qnNbWfF
MivjpIQ4IwLanR36VX0NAwC5K6dG/QBRLKc+af7TRweczH9SnInX6yzwunnQusRmGRtovgh71895
aq1XG/OWQJLrsyLJbYBuigaK41A/xfZaEWoFc5lJk/dw4AvGDXHZHd7nkFRM5xvIfNAsZ8VlgfYg
3sxfRVX3RezublJONF4FSF8rqrixqCQHQV5Vb81UaKkO6hBYFAszID/htqpC46jIPhNsR2hH4o89
QoQhONPAfLXGj5y8BRfZnO2F5/p+5rAKhYFltH41jkeLRHqRL2lqN18wY4zdmyYHHOYJWhWLCfHS
PGow1t/2fCg2VilLVOliHo8VSMNkEkJTWd1Wu7GKLlXzlm0jXQ2/qMVacqM7a+FGO7m0pelFh7Vd
P/VMXYXSG5G6YQrC1T/Ci09SZuRVdtgTlRmgj1+YVU/b9eBQbd5IwJab/OtfWId9ar5yH94bR7N5
+XIA6ygakvBYSAXu70YS4eOVN69GZXMqUZNzNUR1DwEstOarEHsXPCbRax5k8uY0E+mlAjEeFE3N
b35NyTUXwougpbp9y6XfmkSg1n8so0Rk/sFGktF7trj/K8JrQgVkT9fP7Rau/rgS+D7kfXy4WjV6
t+NmsJgK8DrZ7lWvFc1yR9aTHZmOB88z6ct0dRplIPZmDhzmr9fP8UbVpombgxiJKv1aBPSTArqI
yGbe8e0Y50Lg3r2OqZtjKLSZaZ5uPjFFUHRvXggvSGWwtPNui1WYXzw7ktIVlmLXniMnX4U6UUQu
VePDFxaA6gVZjqUAfIg/t4h2UioDPD0Ram7CY1hWjVOkxWWW9YL0LS7MCPDRigbwvcKJj/15kPa8
4UcUbvM+UAUmu7xymGgW6Yz0027XDoT1jZQBqnThv9Yl2WF+0aVfSDBY1zfkIyJgamLF8U/41Rvn
2e6E3/twm6mLvZhfIL+PZXIjolcgloc6F3PA+bsiK5GWbYfaBXRxgRJNyu8jO5LWc3gjN+WT8sq3
t5iOSf9wggO8pP0xXfkZ3tD8NLY+yA44sXs3naLgMa/zNy6oIPEPY8fYPwNgCiyLn56rNTtRrfuw
WHCRw2iGEf/Erb0P46wg5343gQDNSLyGocG5EXDlZ7Y26lJxM5LwLSl2jOIP65/tFUqwSWsJUrj0
aRm2cBvfryuhNPGL+DpAmLOR7cy3Zpb8rq1VCK3fMM8W27eDXFWmx6icLpWzchZfeEUcOow/N7pO
97oZ0X2bH8pke6S1rZ+cPW1gqJK63elNr4Fcp6HsaEisgR0+NuYZ3b14k9wbEHjR7kGELvqn5Suu
ox/p4txNRXGAa5/U1cmW3U8wp+BZ5wlyT2zjvZ+KR/HWPEdIHX9MUiMaGz9uURCiKE/j8N7LMGJx
IX75/j48KHIutMQt8SBlEpXeUgL74yGmugu2WKHLiEGOBeoQH43X765BX/slVQ23rb2iWUFRb7Y7
5RouoK5wcUoWu4fbcJzpsMCaQSV4tiS7VgEKlwS/ax6mF2pRgXn9IYyJEAOsZ21ZRVPrzoSwENOn
6ZYCEeDvKLv5P04E8oiquxUxQuOTUeiR7xo74ocv5q12LWzP2P9ypheGM3pHoN6/HmLWPVU/C6hb
xuYP35GmO7eO8Y1T2yAJcr6hiyHaIoNC311vc5OeqCVCpC5Vf0PhlF7DHYW0Ox+h83fPP1WKmsVA
+OARnkKqjLC7BYFJ6MChhKPowo3TFsadDBUuCihrx7SisZgTqTZc9DnvEuCKjoJOJAuj80vkeZBQ
jSKmfWuxIUDnBzAmmoKt9nxKLTf7Kzh97htnwPStFzI1ujGnr7eWTzstFBZBbFBOSN5hMBMeVKBs
oSkmOl8Hdfw2CgaM5Ky3rGmTBMCh+yZ3zdF2oNK0jn9LZkFY6AYYODxPqInXZc1Mlagsn2qqw7M5
cqH7UGPKW5/2bN2XY0onm84QwFh++OC1YqX4YGZhA4eRpu9cclQ45EpiGe60QeRQ6IseNgOvwcVi
MK6mNlErhmxXSGnJLGdzNKaeQbsmdOsxfxzxy+pVDukANyGNFzrkhQHRFNMakYyTrthjczNHdmrb
uz+yWnr9SjP7g1DuFyj1rs4+T+qNGxeF2bgenzkXuPdriGVdZPQZ3XbEzGh/2pX00MHbVoR8g0U9
KquSzLIwUqRvYAXrp+uSQlqPytdXgovegPFOxLjOW2AkPGRPFDRNuA1MVXVTUUHBSSMW9vEI95nH
nLlzOOIAuCOr7FeWkkG8YavCSNhoIqwQ2iBnA+ONgWO9fEZtLhFPnlv0jB2qFEl6Wk/YTOpyyGuz
Sj01EMAt5ai6tvv4FkJSX092LaSWjk0uAqTEH0raSxPwfFWeRr8X95j8nrlEC06+9wac1neF+4Pm
32AKqJQAFCLP2oGoZY8i83XapKzdlhYsolQl5XZGwaaN/4xVQFsa9JW3i5FOBKAH+5tZLZAB/0f3
ofcvdJ4MfcULcTari51hjoAj4e+CcEAg0v+7Yi4ihFo4xMbxwaamTci6LG+nF1fbkNji3gxQZs6h
QyuET3r/OdzGyvC8JFnZCrm6yodV8Z08sCbvUt4O8l90z5EGvWStQMxkxKoTMc1voQ5F7Xgnaj82
hIL+lHfKNN811Cjpx3jGvcbriHlgy84BxP+IYS++9ejhMK+EdHW9x5Iscvm8xfoiLuM9+GHwhXsL
QKyuqlI4RhJ57b97K+q8s6jHOwzqE8ZG7/A7VJ0ZhQE8oUf7GTXxl/AhapPm0VO1hwlvh+S862U9
XX87IujxYbWiqiLWBqaWKPU7rP4whykjEPBKL1C39uZPOZGIB4XI4LnGctgrk5HCs+mGWC/pr+xs
frOZqYSBkiYMXZJpV+J9tDLx5maTiJzUNDshRXqogC+6bBkcqETL6WPBEn1uI90jyNrptMw15aXd
HB/lT2/BziUODLqDEYG6vT+9puIZ4YzVkBfkl5mpSxfALIA1OD2ui2wwRQykaV/NoBfCXV+cfT+r
5ZYblyynDg+xhEKH3ff5WBjGjHN/6EZHYheuVs2An1xub4qNy2weJcOeAmH4JNVVs/2hZw1U+QP0
n/Pk8LYjIawRaq21CJWyZeMGYsgBq7mbF/1w6UAaqQhMQKdBgpmHoTGiJYNF3IsD0fQBhmV6UzP1
WlcPzfbbEATS/4IxY8yS1++0CkdceDiRgjxWYfsoB2GwJluYw41ggZ81lgh60Z0G6iecF/1E2w5O
P9Ecfub9tlCxNFRb084zFVhkno522UuHnCVjsiyZW/GIT3dHTDb190tV+Fh0h/9dfrqCa9qi7cGM
pM3lDigLqpUZVhpqFPy0N1bGeXRxNg8XcCDIvBo5KfPyZ+Eq3aUezCXx1diz5eFOtMtDlmwjYM2N
j3pE4Rqzirw7zSxooDiqbHUspJhNjTB9oLWeNiXsX3o6feyMq+AvKrD4MFDPD63C20xLCjbx0M2Y
Oj5Ta8tsopWiRe1WPx0cJ9gGfIFvsEvKBQZqN0YGRY6+dEchVS09wqDtRJXA202JWe02Gxd5TM7S
QecKplvsNyDUL1UZKpJVUHGRv6kHjMubvf7RecCV6yTzo/8Zk1y+abf6CS9UtCfXg50yP4pxvFs2
R27XfJq4tN7UHvIGOy/LH8mHUxyXLlHoC0X5E2Wo2AiSPQwUakoG4EOQ7ejRsg3dJGU03hSjYTRp
hlTDyheoI9PSWTj0dDAjLiGW6pNH0uxbLukmcOqPqTR4TjNWzrsLVSjCP2YQ9SsWyJ0fiJYx3/hw
2h5Xjk26YVh1ZSflqOJbmkYR+mWd08Y9yE5Uy3UnXoKhYCBXBAixGmPNtcjicqSyRYQWde2PJgzs
Q2z33+pVj0fZjq+NAP0alTVIvOV3xl2l6uL7rSsGWc8MsQMU7qz5M1lyWKAIiBa6ZRC6tleWIrhi
KUKMvXgu8/MexNblF3Kihrgzp+dY6StvYh7I3joME8TCuzwrCp4hvtJXpznJlfZ7ybgCQPxeO1Ys
nyiOellyiIp6i1bVw9cT09PiwHK4ZJJMeD8kSsZY0DVT3dQIa/tCGbqbHjMy/T2oHzJ5gRWHW9xs
pYATZyqnsP2IhY64bXEkU2/8gCE3fbFLOph2RbfwILkrtKFWHhU9Iy1r1EzxsfgX22TCgPOQkTdy
r7LWc2GFFz9pGG3ig3BZ8kAsJTZoXH3K5QVBGJZbBQ0EgK4jX3cyBYkJL2Z5fl+M0raorbeAINTz
YfCkcgWWGx1Buo9sV/pKVH0dYgfq7aO8olURRM63PrYYJHdPRPSH3xa3LHUkril0eQYocxqoclOn
CIKhl5Kqq83oJ6LSfliyednMYr6WpbtTtUdVp3TwKWgK/bRvdkpwhOFyXKbNruPJ/8vXvMQ2S/Ww
htY5tnBOkuGZDyJj0N7W4GJcw7eSi47Ub29WTCOVOg2pZ2RaAXvgVI3yVGrcMK+NX0DxReauRB3v
8+I2H3IXLqNWjfkLRoc2RmDj6u1qAuN/XPWUuKsew7LEAlvna2AaJ3oLNFoUSX5lOF9qhV+mFbOa
7wuEuBYzG0/DtgxTiiWksATuMYkHyWfeYo9ZgP8+MVTqL2GBRB7bPUODJYxdvnAmeaam749ZZa0v
5v32NqIRW6pfP0SK2oclYrfIN42SfDo81sFCCUfyyQavN20UsMDl4BsgRDlXkCM2Mf0zj3icco2c
zV2pjE1yUtXqN8MTVML5EdSXd3E6w/5hduMHHAhxEZ0k+4x1h97oCj5pskXzGdA3zE/dWLJKbZUU
8CQ8f16lIa37lzDsZ/kMczIgyUrREKMCKi/6ZSkhWVkSGxRYpJzdSkEMpgAY3wyHZdVD645NP/2Y
00QdfEw94bofK/RMPMy+8imuKcMvTWLOX+xZHU/wftsiUjC0pxPiDN0jc6/MpMCy3fN+oEoOU9qn
OLLXcvTO/Z6YBYx1m43GFQV/BT7EGXJbEjkUDiqyiV9JZOSqjilSwLoTcQr5/69VpMBkH9Ey+Lg+
zNv/RVJO2ZxWeDdODeJWHKgGnWOlGrdayA828AetUs72W9CD+TyyICEsYbdq+5fi+rBWek4bcoP7
PSgkT81B5dd7XIsooM4mNxU/DqUKqxN/lo1xi+9OiaaZRrCmZi4bun+ajDnWUVyv6H0BcJQI8gHi
5RD4kukKxQVdnCHCF90efLkKy+bNVWv1mqaF/Q9erQwal9oHQTnFsWFFyQvMOob9Tif73S2IpfU3
4/rz6/DQk+FpeSGp5xql7TohWWRdtSxcqUrPeJqX0mqRyzhHfi7WNqMO36tjZgOBxepGt1LnMi/u
6tVKGS1S7ayxhC6TwZM2a9HTqGhGQjeZs3+yVj1+5JhRA4zzGEJKG/zOm0C5KOzV7/vt0Go28a1l
M99nQiXwS3adnFNXJPe7WDUlgJa9l4KvJacPNLVy4434BJFEFKoljliEcyfD0g7o8tsZPsC3qeIo
3va1sCefiQbderqzSfS8eOBvoCmW3ommOqLcG8uavf/bifmzj4eoWI1WINM76bdkhTuCd3iZSenr
aYc6I72/OSfvh/oMCIAtJjvAo5KaijRdO0KcTOsyysOzCpKu5kMrFblgFhDz9tVHMuAIYZZIoEch
AX6PLujEdNq8ZH1QkdLJAhk7sKcK3ooUaFjJMfzeqtnLCwtcKUtryJIWjSGrYI7IcEWA6pnwm2Gi
b2au6djlgF11giNSVieWcpar0oDvRwhgbCWYrNzghTxCJYxvQTYM1/nfhLJoT+uRtZYrVXZQb65R
i9Fgjg4jg7V61onjadmpC8DxuiqaQcYInvymGbYHRlHgdqZigjeytnh5HOMe42yJ6xI5JPyLWE75
YaDwFUWpFq6haT5UABvirJnvl16n8MscgX0pbshjuof1R3OBcKYNqUKDBAnSJ1McHamrR4ojsWZS
zSW3bGeiMjm/MZ1ZE1Zc373CAsRt+xy/nntm46lvQB/jM5TSM/fDsnpGoxpwkXn008L22dqhmiNv
dZI9xTQJcay8PDvnfwo7wZWSe3blExJGYokedj7EfKcd+X6xN9mpwnmXBymDLvzD7X1OIQ/iM/rD
wH4o8rMP28tl4NQ/DBtqADazpSDkO7sZlRanAMWz6CzEatk/CdgRL/OnqUNkBB1O8cdttH9FmwSa
tUN1CROFfW2genh2Foe5KHrLpjCPgW8wvFSjs/zcZQwUCjP6cZHdwCT8yJmEu4uZ5AfPZhaBr5bf
E7BpUsf8R5MkAPHkVBVwL6o3LEQZ781mcLMsY31ecrxaWtZHITNZ5L0prSxj/Syzy/RVj8PgrI5y
BhZhH4Knfq1CoFwK2naY7kj2a4QyqcAH4FIJ4U3YO/FDO9agKwFsxA2cuJh81bXWtY6KHgRrBmUG
g8sO5hpc5M23qU/5x8gND4ppQxcb8I9ck6xqEYoRDg9lFiIM2QfNdkcDAhG1FV0ctvAkn/bRB7Y+
jy/0084Qw/L4Ubm/y0JVnFyknxpOAMkjHh9G19cCap/ZAT0OuDg7+qeKx/Jap/pcGuAoIJFjirAi
dTE9o/HrTvk/W9wh5wNIT98YDme348uo9loHC0vcR9XX6SVXQ+nmF4iH5iWz++upLJqR6BXtfwbP
yxOcRMG0JQn8eg6epsygxHhXBFUjONF096sYwNSCjAw1F6a6nMciarX8IiKbvazpfsL8QnrCE4t2
V6Cy7IjSNbUWIHzWKqJzbUv/cPwcq7XmN5YM2w2oVmsrb2yUkCltjpoVlvlGkcfq4u9iSdF6FvN8
+u17qNeSUmFKnOONLUgTmP9u15mhGGwduyqMwiAVFOQjzMPk5wmQIM6u/DTx5ekLZIKZPrMmkAGD
t43SpXQ5lTKvsuEhBNw0aEFO5yG+MOvrR7ETFy8vIsA1iP/a6Y0ANznmA0TPY2We6LKR2eo+VJlF
KxwG7TyDP1PfTj+00WQXE2CSGt8H48cLMfv6CHOUejRYFCoJObizVtG2imsL+Tuu7mz0nmfyLE66
4jTuiIuW9lgSuskrHFUeHIidCIpySfGmYU/k85+d6M2dBfY/bt04c5vIlcdd4UnstG/ZIiqId0ix
sNcUtQL+9ulF7n1QBNbE59wRTjjapRFyXkFWU3F0I4m8pNi2Chl6HzXQmh6iMA82QP2UWYBssh1W
/6SJ82uysDKYLWLTi3q+7rAS1JULsAIxP9AkZvl0lYzHFGGw8M0cFlpiLr4czfBIbBl8WO8yAANk
4STTcQzAarSLT+taB0w7rw8llWBS4MFTMAOUO4yCXgWaL7ZnNq1kyflYqzhlf/LPrnIJhzIo2kbZ
4c0Nwh9b6W+7mXpSMUlnDHbRuvtwImuUWlCvLHy2dpNBNIWlSgfaLY5oiI0NRQZJJyBncI64K16J
xRQgFCn/vNlsaBDH3N92++++Zec0jaYVkrnBgj8a7ucMh8WR1bJqcETA8XQb2i4sdwf1OJkZwBkX
sGXt8FXaVpdVR59K/xkK0ko9wWnfnynRngYQEIkb5QKw+p/B4erllTIWisq3E72Ucu+57ySM8/f5
sNSQVBNlbI9wTZS2G8hzpT55ulb94jQlVjbc14wcUm5+7BuS7IPjYlYe1hjHCQs/uiJQdqB76cHe
5uePHBy9h20lYI87+Z4aWEYzbLMb8T7DXVckD2y481Cnv+WO6kblVMTOFLfKqdTdeBNvnZH5dyVm
7FvNusuISv69QmkcoX8aDIEgSnPLZ63VD3ojKD+6HijBT9ZVUuR/57htRY8V2hmnIeYPDwLNz7Xh
PkzX+8MJnd0VzX8tnCgaDryvv+7qz34XdBZ49K1zy+eOFuDoLT+qNytcbOr/zloh6m/iYkyRHpKZ
bg8b8dn+c2xSZgEgLMI6HL1T2s0++Pkn8M4IjdMNHVESUIHVgVFjbZGpwH1M2vMhiCFho0C4LPvM
yCt8PyTr3Ls8d5oHLyj4WQImzlvrvbKJQ7+rT0gZMMwGg3TpoDYdlS3FfZyXcTPlq2SMUWrP2uDp
d0mrcv4SXxInSneQN6K0stxQbvy6szIY60WZIFr86TjgdVLIHAJLUHgPJPHnHDrfWRE6QqTx5650
G22Sj4e9qwu1myQOA64O/qd+VIURD0UA1ydrf58qylxFXc/pFNcIVTTf1SH+So+SgoppbW/phCEU
SnQzTIF69cd9o61GiAlQl+a0l8th2GleVNKCbO5DX/Khm/2mjbBMa0MgbHLcNNNs7NAO30nc9K9M
rBAZFkTOO0y7jKNSuVGvYz1ORZMW35J35PfyHGo1KxNc37zQovMfFozLkWn25QEWguKh6Ri46BYj
xNkTBFFSeYdqbo+iAD+UG8c39HzJLeWJvb1mmn715z+njghdBqp00Tf1cUlZaICQkuw4ejXcDh2z
h+Yz9MynKm78U96uVVK9GzenB4POP+evCTb01lP2+V4ADvXVm0ZYe16mkT/K2aurjwpuEgdS5XBN
kTnMC9H6FUNDu6LAEaLHgYLfyBiICf+FfOBe2uiV1mRyCkYXgcCEdV/htnf2W/j0qMHFNwtv7OtG
m/L9pojzn97e4898NOu1J0Cy4e1u6sVVGqgscPaF59joZ302OezAO7rcaThETgXK2dlwn2oLXfOK
K6IedCsfCislerP8TQkPIfzlnufpt9aAyquOB6OYWCIlejTfaL1M4ZJZWffdS1CDFvbxYjQbUq/S
QS3VAoO9yP39ZKZ299tQHNpBm81j4a0aIWQFDZ9wvslZF0E+guSoOecO6VSqrgNjjr4A8cH4YU4t
Q1ZgvJhveLu/O+FYXH98/QUUPC5QIcqRH65Vdk5A3qtDQkHuM56GbMytb51wYx8S1gurtMTcudlR
OYEXelbuEu4X949E68KPymFK2Ewpq5nPdul958oshztCaSrXI4XObqJ1lA7nX3PY96F8+76Enfrl
YcwNqk/zJAhTn8deS1AuxK5GEc5rSVQ2ijttzn8YBwSAm+wT++c7HAD8jbyKigwzX9CtwT/SdLKW
XqCzFUvnuszIlZWsiW9lDkuck1QXmcpRMlwQzsgk5I195Qf+/07Kc0CDGzE2tHw8dqKZaXXV40XH
KBmxZbQvgl5outOGQIZtwzmPt4yyjk583xFYDmFJ1EFj8lc3F8QLa32XdeMwTBiw+ig0Meiy6K/E
i2EmZ0XDj+duwHvZm+Pp2Y15rFYcE3rx0qGkUHjwDddBZFqNGEwrgDp1wgL3qBPPm+A2qDhf7oj5
crSNwdmOO3vpqZcQxCyCGKo0W6pqUueNzh4dl2aVNm46oYEXfKLGCUd1sedJ6y0tN3FZx5IspQc5
h6bM0VbpSmf0J6wXxskarycNqXmUy+6bSwV/h9QCfvEhJt0ST2GTBRCJX2J+/yYGyfJV4RcbgcVe
QaIkNVY4UJPK4RhYfADlrJ5JZD8iWsgp7dKzPFRfxQyS3dyl51T1ifoqUgwEhC9MPVaZQt7mw8gp
QKdVYXhSfsGxZ0B1k8ApsUh0pywZoPiD6n9qVgP0sJ9JZaGlU1uJvDAzcpXc0PyzvULHKIPNGSOS
XqY0TGIanyMx751mmQrr15aZImgw4c8AMkJTTWLqYwpFOzM5WTbogrDc4XLz/HoOmegSCah8VFQq
sav7ORr/PS37jq2pt2yenqPMEUmuZtVfz2mI8OSL3VZpEJ1OF2IxD4P7i7+5um+tsjbqqjC1Qh0r
m5XKpPdmKMAWK5rZQsdL4pzmwJ+L9OvlIXkFZr24CQqpek2pFHCFUXKwCBk1DtoHaoFifCiZ0zKt
u0VPh9qJx+JwVfhrw8bC1MGROcS7EagF11NTutvJuExj/X4NZ0mn58K1F3PkjqpNWI8FW9uBlk6E
K1zDsHqbY3cbZ4GD3tCbC+/szr+L2W5f3CQ/gxL1XniGI6F5sWUFX7Wp/ocVHFdwhFWUu8ELVc7B
noOjguAeB8QLg8Jf3tq9yz+3qsze4cIRAWhJxzChMOA+BGXdJOK3lApPdBLwiOlMg/eK3eYGzmiq
5xywzfr2qSZ3JvsHTxTbDuQlecSD4cxj1XcFbKf8HTkEpBXNlqT6DakPwYHrCzvXbxP2LVNfO3oh
iYCqfrpYRNUE3tSwSDtRRzut3MD69uk7o8Rx6Je/xHOBPH1+1Zj3AOWPdVyJw5ZA+liTIqb48pGf
gFajAWzgY+GfHW4fjeEG4ICgOQVS7fJCkEBNz7vqd9XNqrdctD2TwblqWMUXRy3ySJnp6V6uMFuQ
l1Qu3fP3vz8Pgqtj6kpHrvP4pWO4Y8wC65hzEtl+HgpshN8jBWAVxD0ZG+phjtNmZZu0GW6Km3uA
oZsClrpWeEj0VLyGb3lWkyFdT6r80/AsCvQ0E8pfWDvt6COzWtITL3hxDMXtsP65W8t0wn9lpT7i
gL6Kup0/3XCurYV+Bp0hWqx+WpJelvgmI/hTYj0rH8fCcgLpHyd55L8ma2Kexni1K5sR4hrG//qx
EjUtOMNX9Ya9RtQ4/dDcXPoVB824WDhapZaM58ZbxTvgHUzSY49EkTo3qqhTdhu9JICkcH5Vg8rm
OXVhUwDmzIpjxiGQFpUsqO6+7Zw+sj8xMTh6n6lS+yDBzoGtos3cajCvkh4u/FNokvmduTUwfhid
mNfHsRDMCVjeTK2mGuhx9kl8Cz80EQb3ApwuNJm75OFwPxLfxRGJSxecU30n0KmmqdRJnLWU6944
dAgFvVbYOGXcwUJFzL3C9aSrRYaAzlVI488VWXctlJy41DrLIX3eLw4vRQLkhdvInMnVDp3CJLGU
4zgE010k27IW1qfFUTbgshj5F8KF1pdwgc/3mSM7CFplgpQOInzFBIJaguJ4VSio2EDzom/ksJXr
PCwoE8H1ECjI+MsH3bBpfc9DrZigdFHPvn8BSeafydPXMeXn/fRGma8zRMC0Z8Dfltg873B4GdNf
gx6AaD8E1006vCed8eqqXl8q5IzyHD+DtwN6y6Ix5qVfmIQVCPjDdvAlmhLI5O3FjmBHSyxb+gcq
dejIembi/JNUhZinc6pboIfQpLeGw3JgEc1c3c85Yj8uT0/OqNP3q1MA83cXQnf+MSTggxFdzO4j
eoSCsAdtfnB/enSqS3RYMcfZX4h1JG19M0xtdbWHOLVtv/V1hYjgdWA8BQmN6OZ3Y7ISvMAevM+G
O/jDqm+9aTGb7PIm0nL+knBxpQy8P3l0+ANwz7vBRFD2kHG0vlc+zDFJzeVUutphCIXR0ftQ6OaI
SoCqioE4Gs2gNObiAGB/VsOMlrVrz4HJt+gaCYRYNlmhZKGbEri5tEZmPJaZqSWTrmi9EyPNePbu
yXsNM3sxZXmI2w25xHRNCeKBF+H81VQu1RE89jm5/WYTwaJqFqgp7M/+zmtLIUBRDzu+DEKXGnpH
ogNF3O4jr25tPuOfWsH6wBAXaRpt3HmTQCxTsMyZZU80jhPMrW+JEp8DFSEXRu7UWL/8hDf19IsI
Qo2dxNvKCaYTOVKChNRAWmqx6a/gtuP4rpwFTpuvSJMWjucgaBYb5nSw/LL6IXuVNxw5xVal/Zze
lxrxJa54jyOpQXQKfqrd6TOJTTvr4mmZQvz7R90xifsPsiyGOekbkLRpnjtQRElHC3QJ6oxpgxMs
7s+vFINy5XfKWWTzIHh9hjuG4xVNqopiA0QCF18wUa+kXW+zsN/Us/v67Vy8C9pDtfQeLTa60jfc
A/Ev06STdzkghEoK/+DdCjN43C72cD9IGMDq3mV+f1rUWjVBLEcyh0Fl0R8mtSShKfhvS8BNErbL
3cS07EnUw+ShPihfbdAVnNXyEbnsDeLeBxOhU7pHTYq9f/ksi4xZwGa+GcVtaA3cBzyuaTD6efuz
2l6IYw3ovPHw8rgG8bG3f37p6XQng0wl2gGX2oNrhvWjnVFW6UvnWGxBytcgi0/DTMQe37G5x74D
Db6kOAHabMVBzSvubEqkWC/eZaS60QgX/svaTTbCJoa7cWWqjcO1sBfIpHan8Q4TChDZcM9D2wkm
ZbHR/rQeVr0rYlNvm4J2+gmZjQzzJIIK8Z4Mbut4m2GgMBUtVDZNxU+kOg5I75UvswmcY+UCQiK3
Gy5arLXSY/BiUQ5A/yDtGm+3Bc+ozgw6rV0HeWXb1Gn9m4N/i15WbzFQ4ZFZTBTfrMH+Qmi9B17b
FZPUFzhjOkJNmDuwnDzc1NcBsoBjeg7osueh4BwOKngbxGk7m4MYivD8R44XH5KgWyYwqX4Q2jIl
cN9wc+pKelufIQhhlApzgHz+Kvs20D5XaT1QCUgX5DguXwAen07UinmDMp9q4+OVWuXsquEFl3AS
cwiUJiBQQK4xAkT2lWIfA4HbPTs33QuM/Pt3LSz4JAM+tM4RO7bvMUnmLsCQUN5HegUH2K7zHHhA
/0+AaqlVuFPSuqJ0csitnzCMWjiF4dglkAbLFKWS/PhiP477tLWGMZIGp2DizrtwNYZtV7J7UCPY
eqFOkStlW+pKw1E7oQCtmvqbNkMg69+m4e8g8HcsvE8PM44m7dZNv5w14milyYnIazKSuY5aMprg
3Zagwxj1pQ64FjGdLJiWNN8wfHO0zoYs1g7UbTTikVn3IDx4BUzpkBOmv+9N4J7TPTigOcBWmEqi
TOTN/29eeVy7uAgKRhTSzU+I6aqYCeHDndl6keZtRCYgDwQITOVmBawY+iKMnhwTsw89lOtDJv9N
kPzPI6QteoJSEPzufWdAFIcVkrtb4xFJRAz4ddEAPT2ofZzQGvxPVdpE4mxgdEPPAz5GIfzsOVQi
W0me1807jIbbhWXevN9kh0U4Pl1htMIzfg3rATfU80ZdKcx4VEV/A/hHuvV5GMQQ3hCbw19Rl6CG
XMSXmMgwOqvN02Suo5AszHEM6HHuZULUSu3ftToYzFC6AxO3Sue/m/Gf1dpiXcIPKiUroYO0SXSM
QBDTM1AgOxW05Bj2FFk/0e4zZpCOTEvSmOHO9SUiT5RG3RK2kJd52kqL6OxRpb7DK8ZQicYS17PB
j20vhSaZtgB9JS70G4VafLmWsg2XUj7c8JUZfF0lbs+JAwXPUeB99WnAYtB0+FUKhP6J0P5hJwOR
9UbUwfbpDQQ8x4DjICwRVsxNG63LcgGR1mmTXlpG1vUJ2bFTQwaxtvQFdv+3tdKHaWo08QT9pHkC
1ghwojWidQ+/iltB8OSQnKxnfF85003G/pv+Om89wlkg2z75mzUNR+EIQhtibbXjwYzvO9zQkytz
tFMjH3Zbmu1U1Qm5SSYrjqBVZXmeYi/6dM53mV4tay+9A+PQhF9wlOL87vZcreqwMjqKJenKRSKf
qDxTUFUUrwxfFfzmyIV0O1S70Fj7L2ND4E1Wrt297qjMLU413M9F1yxH8Wz9W+SMfeCVgXUtreYT
UQWBdWM3pnQIPC42r3uYhe1qtmYUi/j6mgbHYd3RGmEJcuqN0WrZ732vzElCUQjFLA9qy1gT3pRu
XY3ohOMOvI/Rd0bJadCj2PGQKorbra+i3gNnmR5GgCn4C2eGA+Trwc163rkKg13VSMMGtGLbZcbo
RnJp5FId02L4yifQ2qtCydrt4LO8YNrNDD/JD6F1O7uRT2iKl3HskxYRx+tcSUh5v02jUDQH0X7Q
ZrOdY4KUW3AcWUIJHlIzwLC96Uqf9U/1fywPMizr3sSOz6UoBBF/A3DFAIyCYWgIBn0QvQyxOjFh
do9bhkpTkF/Us/uGkTlLWp1cEG2xfYzbALFHNjjEOJQPoenaZEn15MXJ16GfRKC/dx9P5m4rAIMq
7XYdGupqp5yKr0eUCduwhVW8aBeiNzbiFlqFrfXUPQNR1jYGbKxvN7Nk4lxUzvusZE2rBU+psso3
NNAnMn6yCTIyJUDIUh09EyaTgy11gXGmN2FAE3Ixjjo30yuz2DqI/NgIM9B8YWa6r7Wr6CedCcMV
VrbUd3DzBoeF+K53QBh3nf21G2aqsGBnsGBwtOzd+lwZI0Lf+8erg4DM6Mas9/QH68Szvs1P1oCK
YGZWEhX73Vr+DdzjkQt5mXIZL4bh5RFHW4Cr7ZLK3Y0Lq4x/US7gNmh0O4hG6y2FfSYn88/ZtTRm
VufUqxdbCQhyKKHLXlFmM5xHQg4AreJpOJ0nqSdTz8Ioj7QSF67pwW0foZaIv9wq72d2e8nBGWI1
+6wXVICx7z6+lTz3uMvjZxCSbdi2gOBDbUyt6whpgaINRimuxm+S4CWAuLyES6Ef1lcJ2EY1U91b
I3Mg5s+bkVAPawtaO6lU3TjD6h56EGHKzENWoynDm5+JLHP+fdeVk8yC0uhBJjuN59SiB0wC91gK
NWUiLnXPAzPtOeeo/oWDMZUH37/TDi8uCNxHOyQV9/S9pdiL/Q8bXHmsVS5bBk0wOskfPPq+SikL
y0iRlLMyDGqbQUXV55qiFIFZJYSQfQer7Ix0eEc5LFKuBiC/J7HA1c0ZbZeTuog2nXrCrUvRETWH
C4XqWE1xQ4Dz5fTclJe0S209YS0EzRB4O86PSyvl3+U1nbldFeuHnNC2w7OonGoOGHA6eKZKDl5e
d1nlBuJPhOrFQDH9Db0L+vAxUgHZ5tDI+4C2M91+eRXOBVdzj/hs3NAqB7WWY2BjNBqNo1Z1nHBJ
D/RB5ZDPFwoDSvOwdAyv1JdlKdlMMow/Zh4m2cF1etfSGTnGHyNLVC0KkT6Tx9CwzZxK8DFcve6a
uItP351VhGLPRZ2EMrvBiDR63f3ZPm5+CuHrG0zr2cjlM17ae0OkKSIAuwpvRrOe6BhRhf1DEwbx
hpSJedTzqtaA+LjPhhYJbihoB3guCHbiejbmK9/UeRjsSraNmFOKnlg3YTjFTSWaqu72TQzpn4Pz
AhuogqwvthfsOXxWaTLDg6OBwXEx9WVJJP1/3kSOzfZr5cZbBZmKr0l3TArRhtL85TOY9S4lgLzz
/FScqACaQtrtDyFBUs9ULmKPhpv7nHsGy7FZXomSU51Vyy2/I32+YdZXPjr0HSLzXXFDgG/VEeeE
t81H6A34H+Xd6f7eSaODrW8f8E1l5p0pwDASla63dttV05S0ILXfDxWTCiORCm6RNN2ky+ndYVO/
Z9ET7z+Lr0AnUWahj3DKp+S60tzX0hYqs0lDfIUK0j96wI55PENkMZjZPjO8RciFWJ2llP3ibAQr
7oyY7/px8HaS0aqSLnrELC/gtZxnGWWQBaQ5Eg2fb8GEvc3U38+pftLeOnyQnrRmn7Kz/QUn9w4z
MlVU7B9DbfXoFE4dc5/MSG+n3nRwq8WikXwZ6Rn24GXhFVyu9xTbMhZsH1sjbTIsLwn4l/VMY788
VMZnqjvfRqXpSLyZ0sPJUbatYFxzFxvIiQCy9UhUebOUHnLXGOYjPOxyZtVPY1lgssvgVEackg9q
fZdtaBXEW1230sdLTWSjGdUCfVlfCWXG5uh3ATDifpoRCc/oU66ejbQaYejJc6WRtEq/kFBCRjeU
1CaN0hnpPujf/TDqqC6FCEzDcBBMNMljh1n33nlgD0WmU6EnznFomc4cQUImxPt8sr+vtE7qyutD
rk6tz26C7XI+kjyrXC9mCqwai6HT1Dp/AerVZ+AmHnsiuO/7TA19EX/XTpfPMZMNRv0Iwq1r4+of
MivMHM0N0OKE6l1DE84Xv5s7jeVJM+UdGQHCTKiNUW2Bnxre0h5mK3t0alPdLFC/UePiqyeADIy3
LxQH9nDXwsMc9gILSgayrB04cx6GmDBGs9YivUB5j7vdFdel/ZZBueO9f8NpWHCfWBI+ZOEJcmP3
SD39MQRh5AkUNcEcXJRf1VPR9YeC2kZG2I8BsHX2PUlA9IbgChoB9LCFxklvW7LpvwsYfFwWA46q
v0Bbankb8Tbe5LcJdPfkpaHospcxfXu2oIv8j+FdpnmaUn03URbQLlQZvfT71eQUkfG+B9KG/c1m
HN7Jmr1EVsxrXpwwPVIvUrQRX1yg42y6VRbeBIZbjau1s8rDorwAqAFU6JXQgtv3xVc5IXr1L1WG
5tekmgboJYcqvgLle9bohbT8rmv9ZYiwWoOarKBu+PC9OKSIZSx/Ya7l++Fbuj0ERwctOPXh4Bwy
ilQaPAPy5IHXEtWWnc8t+BWgA++sEZj1eHK6kjRwUTLM9MfJAi48glnLp4gD30B1ApVfAbseRreL
vmpdG/yUAsbNrtqgf+RTjVhDqhWCgqVhNTG0ZZOiJxdICHoCqsPaeQ2knWiTC+ev55MfL+WBHrTx
cknryGqgRBV+WMS1X2ZqDayfL0wIbTWaBWEMR7oZG7+D7ChD0lAqupr7DEgPBQlsvQwKEuBPp813
EwlaZw0kAXWuk5UB3JxyNFZEKxini2fMnIOOyABnZk1K51umEPg3CUuL6HkXKjXrPIkkEO9Gzkrd
oKdHDFh+CAfGC4HZYXbSdmg7zkhXZm8qQgYGHtrFzi3e/e+Y1VXi9q9Gfkya6U5fCsFNYNkkzkgC
GLGvEUio4hZxfMkgpy11wVh7itlpfaULpkp48MMauVGAUBlDMNrfMAiZXrrkcwq2xX6ghKe1njLL
+S7Qtyvz4NRu8l8wFaN5vW7BXHS66qjdTyf/7VgF2+qq31g8KW03UTpx0JZh0Vpu0ScsrrePazkx
gRBXAeWgTvjUZ7dbyPj/iOX/UNe92WMOpLtSvYIFtIMBQyVekCDVzpZ2VXF3HZI+nUPrV37Z8nvU
TxFt6ZfaTBLe5BZ2jeOcgWk4XRqTFD/u6KtL6cyNjf3h4dPBAg1DqQwJOw9DdKAS8e8AWJ4PVcui
qFlQF94giihc7pCUI73XLRK6cuueKXBYFIkZur+sSv2tLnmIGb6x1UB3RU7oIFHLOUkIWhrfRxbq
6i1Oxpufvk2hjRxxaBr2YT3AC1mt5nW2883z68QD7GiUMqiWlrB1FuNxJs8qnDWWZqDzQSducrZO
qlfIX9jroEsKnCbxxu9hCUwneCTJ/sC13S8UowlQzaplDfct+vl3zNhwhqsHtmlXvQd7oIcyCZnG
pb/558ws3jmjBkObxBpdL7tiE4jBvKGYKC0YOKPXzxSSYCXDfR1y1I/ybK2xYLnMgaF3t4fyP6Wx
5O6twGQicgDNqKi5NjpU+0REhWjxP4cp1LX8SJt44Qm7DiYmWbySpaXdQkIoy1qfDybC5HP1s7RT
pEQWXXl54gXcDsI1jeOyZeK3ab2ub/T6TIE+b294rwGZm/0ccACPTW5cXuLLhTx9Bp11WfLh4t/b
DGlSzjF6Ow24SCIMHSc7Y1VLkabVb81YU8CUSAgqi3FeX19oF6jhu0OVIlVPWoOZvJstAvTi+N8P
V7t7Bz1OjMPsBH3TZFKgG2ZpH37DGBeyC8zBYqNjAd6/kFYTkrt4LIEYnGtss7RSF42JqdWa/z5w
IgBzDApDAA2arnYrUXWQjJmQFMJ6x1+ziWOVcorPLYAUEmG/mP2LzfU8BmdpnAMWENINC9z5amlL
+IXioLTaPN1lMiLl3A1ws3jegaEziiR/W3PfbV5I97PE/9I3NSNQGF+jakNJBlfFuM1cUg62XD51
Nlsgqii11nv+0FYvNfSaSo4BfUIzpHYHGzt649ukIwYAwK3ZF6cNHXpQqFxPO12iRkodsXFId2JT
OxcP96u7k13sGEAzTFWWQSYJARnhROhyv13E90ywmYqkqcNcUu4REkCy2BIC/Ute2Mx2DbDEWBDA
XY4md/Zx6ddTcWJRncEHqPWgmREzGwH27vAxEIrhtS0xfOuRUUdi8GMT2AXmQbLet9JkdkVT5BBO
K1C1cTY1X7paOdwgp1FmZXOV4v9Vb4Z4JLKGd9xSRgonphZaZ+Kg6D/80lTTz2IZsOuLgnecuSZK
/Y2i5onhGgklQyXGA1efIZR53vzdHH5WxmT3IadgZYJkXlInlC9C3Ehy+STs4FrCg1LVMw8StaFh
9Uf9F6dIA40965LEh7MMH1Y+W/0oMHSKLifxQOjE2D0K6JDlXVEGHNi6WkNYbc66koFXyHqNx3NV
JZ3ik70/rsxp6x4Jebx/RiwsLejm0S6QC6mhzmVmDVqsFJZwOEsf36garSiM/rHHXaWZqR7SS9FO
6r1/T4XJn0a3wKcEGcnTcAJvGmigfTa5Ml/+/Cy5cxyI4SF7dtDHTuCr+AYr51B2eEE4Xjv1tSVW
7spQFXtDHvMODO8DnvQZX8+xMc/tatiah1bXtGZ2FYe4FtPbzB1evR3bv4XUnwe2SF1dH702DFbH
tz7rg7U2TrUsgpSC9XzMLyvfJI14gD+X6SLXha860f6WQqyhr9gOvLs6DmnUA3NI2yl43A40xiYb
UDlF9sXGYOAp4gD7TgpYycqPoKxXEIQkIcbElWlpFAJeE1Ms0vJcaY6tqOxs6Nqrm8W1kJk6RwI4
4uzZZDJD2qPGKpyX4Eob+Eg1+ASJUd8H90Nu4lY2U0+kcbRQGKdPwnCAqMFjPJjaq+YrGQKlSU5/
cPUWGpd1AQ77b1n+VtNQ2ojBnDE0dc7QBf6ZfnW1vEByg7BNX8D7u++9RB24T8gMALaNtqN4xUrc
Fij/jHP3Cba1/mcBvLd93TRgR8PnrqUDNUkdZ8U1ZahV4fNAzKJM0VnCNvHNsb50W+qHd1/Pzfz8
Wv/eU4Au1niLjQvcWK0a19GQ8SmZco2z63NJVdaYF0Mb5I6YbETswpDsIiCCFTGCA1AjALKXe0ey
3urIfMbe5GOFqsHEvVs8un9L9BbBWnIERg4MDp+niGxxlm4l4gomBBdbXyvnjzTLmpYnauoU/KKP
5PPW8QtTOH9E45EHxRwg6ju8fH55hMB5OGgq3F1Y0qqknI6e+69JUXIMeSFLhGUoluqm7UjR9tMC
D+b7aj5c473+U8ztvi32PajPWYZwn1QdMGEH1dJQKB5D6YPwevra4LpOMhUrTfBvcrMa0XNtcqGi
Gi9CLB6qyUVWXZpPsgvvaBbkYgZ+euqZf3tp2Ia9irs+vTsducJGIeVSW8owhBy3sYU22rOR6x4o
WAqPiFytTVrP31jh6NebhfOZMdDBmDAGcIK3NeiRFsY/SobZHRKGC5wmLoZBsN9CbV062EnyoJ/q
I0Csw8vvDLLfQR+Z3pZHk3eDfUGW5nHDZykPR6DiYCLzpMUhMm+3Ak4D3XAe+r5NyShlNQukWEpc
FPHVI9SUUi3CiQPccjSQ/LwMi4ZKWQumGcxC68Vz29R2HxsBb8gny+Tqi0fiWKba/0fZBACjSjbQ
bM5iCxXzkVU6bxSUbOIAZiJ/zxX7NucHFrGEoowiTmFp9gM6gnCq5/mOyclGP/HTSwBIxvnvT6cV
NTxFAS6bQHaYDCxjB9/nvQxbuZIe3WY5go36TGUeIMGelg/0e5jo6lqD0TObTNGqRJDcqnLk4LlP
7JnNVXC9luY4q+TzRsIWcUJFxLU3kG/T3IDjEPcgn/1ADW+YGQ2AqO+bvPMAJIHORi490THImJZ0
XOw4V0xrudrHGV7BNgyo7e9X/mZJZJbGtFDa0TnloEUN5KTWYNRzIWgnvA683Dv16Pc89y8SU017
2ZUyqyZrkCMaaGY89ZCW9ps4camsdDh4be+KoB6JPsSjhvGhGR8hfu8RnWl+EP5ASSNfS1Upk3zx
SXwBni8C+XodrhMZOjUGck81Lfb3AyUubic0IgYqt2PArZgguUnmJxKNCHBhbmQYARlLA4puVPcg
xP+vPyvGk3deKWsQ5j7SQaQiO/lEXVkl7lqC+Pz/IDyhDP1RBGyyQvqjP36oIpPNZrXshLNUhEGQ
ca/nrXQi+ma955/Bt9fwOTCwGJ5WJN0NIqZ7beF4CGI/4iQzNcP2PslwpCnSh0oqLCXBgHF0zqSM
ONPiyMQJtFAt4N3j8XGKzTqVpTJ9Y5R8ZW6UihS7sBxlDuuXu0/kWbfqhWYQttS2udAxQuohZQ5e
mTBDdBaI5lUlpYJxD+144U5lQaZGlEOpxQpHIUV6VBFCnc8rNylcsX4c3Gl+k3bff9KohwJKNdVl
3s6F4wo9Y2FxzHW2PeeCQPJY7uymvBHc+iaEbYIGtrxrBIzlSd5Ma7mi84GNvPf4nRWi2/q/Ae8J
YK7Pm8G9FZ7GBS48xGb/S8nUP+bZ6Kw9GM8Qhn85em82CRgnLcgdPlWlBi1MSamA8nUmHG4YImzY
zfNNUg9c4O3c9nUzkoUm3qRfNOL/55CCyO+rTn7cv7QLPV3F0caJV7kZdLw0Z+mMT98Mu2R16bYA
bJamPGQPwX9iUGmEAA6EY4alX3PE+fwhLqYVhjtE9NtrWA6RUj/6nt/TfmnMvSEZmZcU6BhF/2gk
0YqzvY0V5DGyeEF9m/0PJJI4TDdu/O2z+Xaxw88Vk3Ka1NUYq97P3lu25tsPRbkk7MzZdbJ1NkJU
Q/Epn7dDWaAs0gP92dmU2pd6IxcXyCICODsERDT5epbo5uJTSyTa+1NY2KkUS5xO/Kel7heuqPfd
7/UAvMtmDMkN+cpMMvFw0boyBqBgU/NsVWMHw76C9nRjn33TtFwdYefxLARji/5ncHe8VxUvtPo8
O6OfIB+CIEmk1vNhs1Rdf5oDR4VxvVO+J7osuwyFy3dmLMH5DSWI948CQq2W5cog2Ifh1K7XiiYa
pv/g3fjbYSAtBDAWmrlmCwBhbhMVW+wroVAMBBQD/II0eYCC6u2CQK2FYegKqJG6SamkDB/Exu5T
jEE3MsmOX8+7URhFyLxQDxpglYwtyr9anxNb7zaGDu+DwM/2vfr+ppww35GNK5bjeJq3kRybjAD5
4cjVmh2nV9tQ54gF+O62KgJsOTdhStoEmlpVsic0rarkDrLsEtSLDsEfdJ0cKuHFrZsEn9tCbQWf
u5hso2ijeaZZfdcdXXfGkw28LSBWtTp3qI44wAM0ALR1Hg4Gv4EfGZu7/g9NYvF224zwE1o1n5pX
/Xad5OZPh7eGOWBvGOXpNuRbPrfR3AWPeHEMnFt4HVUvJGTndFcEEs3PWLuLPtR2iAC245OGnlDS
ZWwQ2D31VhYNwp47rJXKXvKx0ReMzcuOYcdU+gLvJd+K+TjJy4vfAKjmq616UKzNWkKApG323z6v
RPHNov+bDgfjtvrRTLMNLIH//fWSYuK8mI0QNqOMIYeH15IUjjslF7C/4Iwm5Wyrjjk2BWWtM/oo
U3ij5+zRngIYL9pnSTR2T+dmbkvNIPvAr33xvGeYjjKZvAjRopv8f9nzMxq2OjLNs5QjAg78e0X9
if8S/u3vikgJtKVqQPAxjhaCeAdJ/7uW9d5wibQ9n/fVkoWYpDSVnuhNQvuRmKZY16wKPugYkt1T
dPsX5WsizN7h8QDbMDdNPf375QhZS4XM8QsTs3LdRo7mfuJGZmtfpLK3qjMJ1gIxl+RJiSAjxG42
W2dgmiAXOhkekNsr8ZbMzbU9454i7GkaAfuIvc7NpUtxsrOeO8KNSPUQm5++wzlmPb1G7QZ0KJqa
LYPW59ZXTtIcfuQ2ZjjwO5AYZv1Dfq+ktMNG3JPWmHIM+0ksyBVGRDbXP6At1DeBOuH1cVBgekGW
ABTa5ivKU/msOkmwtcmD9tlPItWZ6rHoimz8yUEqdmMbn8K75dGu5ENJilRQZcux54zq3FPUMNuQ
q25huX6eohWLWUApHVFGNsCFPPXHJOiBFAWMFtJ7DiF/3R4vp/xx/S+ge327Evl6iCE0U3O14Ym+
8sHEf/DBp/GVL45u5qP0MeZiwP/XUU/EtkeMY/q0sP0FlUWMH3f3FLjxXSK2pIHO+q7tJTCTldjk
XmokJ8G8Em7F5mpQGfV9ABnZiUjYROfHUNiya789sBMQtIPPYUt/NWJtn+TZSL/IZRVgojJPohlr
Jb/quPeuwQ3kiGznS7xxvIConuc9EOhg9tmnka/V1BY2EY6/W/Uo2AB6Sk3nwtA7eg77POMqEKvh
AuSxtFN2q04bMBGXteWFNeadW5kXN9QL/6995OlIj4lCY2AzyFuAmctH4CULbyo1WxYUmsjewSqw
PMh8Bd5QCESRUgQwG69ikcq9t3hRnh4YYtzdkHcMa6WEnIP/nEJcPP5Mt3DA209MX4JzDUMGkRMC
gxndZSkwit3mrN6V3tLMVFFKRL7nSOO+0oh1ct1hsYawLZRZYVXT/uAEZuvKxkJczI9egHkpTmQK
83mcooVoiWzoFGZnCKJ7BdVKUbcHvUFUMDjRNYnYB1OZwiX2pmu1n387UELQDCEPL24x47j4t/Za
UMtPYJA5rcW64PMiBAkw7bDKE+5rmKV8IDeuv9WmERwHVbzdCVFTPjCzANiiirUtNVTXGFY/6nbW
Q090ec5UmW1Su7bWAFYP0t47zSYYag5J81gtMcylPzYflx4O/8/A7Di9LHM1Zfz83r0bdLEwL5zA
bahD7xyGtwjudYCruXPvv+h1LSHMvrTTA0GeHQ/KPLXv802hShfr2WsgIjK+DmeffrDHcU2KkdLk
e3FrOclvZJ/QfltQRScV5kg94vYZYoMsPKn3cSCvXwaOYIZq1YNjQVIuLjklK75eJhmeYXGsLtuy
VKJvfifivDFyN+tFEM1AzuZyOAcxLHY002n4gRirWIFOeT5sSNcb3f/B/4nQiIWsi0HX7zVtVBV0
S04t/elTzu0nhNgnFkxS1WB+s29HiopGkotBLnc6MCVmn/QUEct1fzrxPvZAtLlXcPhn/zRy7DKS
Od6851Yl5fccu7FrwTnlX94+V0eA6AIdtfbrnilLu1c3qtjd5iV/d5kHub6wP+E0FeHW3ZCFPv8H
YcKpq6IwqI3Gdc44br1JFahEvdYdrLRH2c+ReqxuG+7jmttF64XEcbl7ETL/lucEvkeJPc0UJbNU
KbVHxZHBxJn21LrkYThW9g9TyftFGAYGFOjlS0uEBxMPthT0sFg4Z3jWNOfFzAvg5iMz4SRFnftH
uKcfEVJYWtF9YITE7HmrvKX7VILDov1I4z1cRwt71//L7/n/WkYdGeSDSgV2FAux6eebKhQD+VMU
hOjXNP+7+iU4v6PNEEeDzkowoA4b+Q20eZDtwZhH+clkOLuTLEZsK0G5X8kTVrI8PDLTG3hs3c90
MDnUBnEdRpMuestyl0Xjyd47+a/NkUpEl+DwHhZmjDo59nzNozjjahCleDW9E9+2X/DC5R3gIHiW
od6fLPYkmiqbBixaYeg++NnFjLNDfjiG8dtc3BvtxIUUxoYKKt94JEEFpVZIKUpSsifRaawLGyZR
qo/N/4rX6+0ggqAIqoQCwCkxNYWfnlNzoAjrDIM5vTAYcxlt+Xxu+DtzmZoT3Y2IKr/6eW0ZQO5E
Egzp+dk+JELe+d2xZeRMrRdI3kZT6rUiU5NLwJyg9H2ETkKFy22lhEp2xOd2d3+ACG4p2UROwfxP
1cfB87d76PwfASHb2SESoKGkC27alDlZKbsLv6qAJ2sh32FRPA9mGambHGG6xjuPm2GtTpZ6RiWK
YLIjL+wjMAeE8yA65HnwgSyMQ8xkvhdeb1xoObwDZEgTav8pegpsVzKd7rSshLZGgFurMZFWqtDe
yOwHhuWIPbSgFBpvZvbKs6XT6PdQvFoG/hVxLjdUPnGDl1Cu+n20M7hq+czi/3HG4/gVfV/kmiX8
tJPHvodGJyk/NVySB1A2PH7XSRRrYaYtdJEVumQ4LVVGJkc+UEY9Tt0ywSFIDiOrBEWF5Pcuoed1
j7oS/0qQtRisD180VVgbcvqmSNuqUh33RG9pl4iNY+l0biLB7A1lkSeVIweuoMx9f8m5zrthov94
BnKY6u1LPlRfE00ZYm08PrRREOfhPOpm7mHVGmw7e2oQRGouDlJgfBH0fW8mOQEaUjGc/tsGhSjD
hOy85ZGRxkG9c6JETUM2b1ql5/SqqHfiKubYaT3YqCHkkWn+SKvyYsK1hFvzWMRUYsFYpSKwZftq
UJMJqT/7eH7VZqHe/FYbS0MdOD4cCHmS+8Y+WnCuZzm+Rp4nEW7d/vrrp9/2j4FF8C//pTEMiBTJ
VVBFo423CkMU6p2VNu7WK2VkGXN/USBwJTFM0lvZuqUFhzl6ubmfcoeTDUMILdg03QmZHOdm9x+C
yqQi3KPfq5sELGsyrT8V/KfTKjqgLoWnjEL+68JgTGbdH0q6vZDybVO1lYw1myQ0J3iiMmVmSf3N
vHaj/PvjwXwqyYuUpOokHcsF3QwJhhwoLNgysEfjxYkbEOS4EiMXK9WwO/GlaS5OmILqz9sExMK0
6H5vBiSO1iN4+HVHkQxHE21hTNpVHnzDBs3568anE1qj5xPa4emLyhlqWq0nbpbBLryos2owRyai
bRTqTKHWHFK1kXPW7O/JSZ6RIqAk1h0SHYD8VAxt74bB0C+lsISnLlA02zFzWeUr/Ok1jw2wny+5
XR+BYa6gh4l/qP2wUI7uqukclZSgc7CwCopTkQcfF51mQuL0Nru5753FL+QKOgptzAqNqSbbrt6c
et5LiI0ivTGvdwsCmajjdttOT7D74EZkyn84tA718GCxCoCAjetQbeE8udSeZunPbIGIdyaLiK5B
H1lG4wZBlk8eTmvsMHq/eUjjT+G5gLwimz32bBu88cp8ygk0fTG2bXW8drpSSlpnPcddQG75qRsQ
nYmXAAY4b9QxTuuy8cLVtbz161W1xgeMMGectLHCihUTwEmMS2Mau9vzkHDZPcrJlqeMo56GbVZF
4zwbowMRZkdd/zoLbE0BRzl5w8tDlMADxwBF+91kFV8/4c7Aw60VTXMJZBCEQHADY62R0OiOKYIY
C/5eTqRBGFHdSNDPLbooj+EwxMm1LybQfAEmZBchRHIzDOBiU6oslP/vx5DED+DHfB4D7AaVb5WN
N1SbfV+h3paMchFfp/sc3iR8IM16lvBPfHRXY6kdtRFdEoc/32RbeKOhBVLOqTXp5VwhWpluJ0Tf
I52oj1l9q93xDvcC6qqHfKeLDqHULobCxGRSY+28FbxxRlcynpzITefVhjJlHaDJuGuFpgFjMax4
UZ+XTjVxASa5Gj3yIOhuPr71jJTbRo1auzWhVsPMBZtWkWsc+H7pWueWRGO/rHh2d6cqj0jbn2F7
WshXwEakXjDnnSs1x5sPNCzi8O+s4N5JEXWyThYoRyJ/LFvfpcuCv7sLZK5RLssWx8Ha17D+bVNq
hvuTSTxow6078v+fy6xvXNaDx6G2lXrqwMxuPj4yTV/Vt8828ML3B85KVYYAVC8gJoE6eMxbzz6w
dMdhN4Kp0OtQ2utzGupOZAm64TXqtkBwvGfBETqiJNWQ6edPIIwmozRqGMRsyM/c3F3i2YjD0zBl
9lMueEWLk69ZdzeI+mLIQJZ6QaITO7Fe+fso1keToyza4HtUk8qvAqkLM3AKZ8ROwOtMu2TvXanC
Q0TZPoO4Vvi6YgHTiHqdEGpTkHgBIcBGQJEmCPYwAmqFKWQE1gTxlJ3n6t+Z7CXGKv21fkq/nGki
z8xKzxzTOsTXabwfmr2vcwFO4wsh0kekfzZFABRTjJVChhZXCmjn3ttY6kwk7Is/5g1Yd5Tu4fDg
obMN8nvZxxMqbrnSFWFGbw/50A9ktZXEhL4FsrYIQuBlS0y6l5m1smgiDUXBVIDKfuZHjkBCJpQQ
PK5AvX87fiF+HcI7RoOqzR/9HDyICWmZ0UHUSJ5bdEvpJycsMuehZke8JVlsCz/iz4x6V2xK5Xwk
YR5NeiQW4boarlrqfRPTCeIWRDyDQohapm+x2LMW7beoHIKZYFHoDR2P4EEh2fhOA08KCIk/rZyI
oCUhnXb2oqfXA/0wf1wS5X37qeWLrW2VT4ZV6T8z5eFeueZWzgbiiLkwkFNBkGKYL/qCO9OhJaG5
gJXdFpMe58CKjOYUAC2vsCd/FsTqOGudgTpVmQDq3zP4S9x37NFazoXxFuSW+YAvk+GX7IzkydHF
8v4UQPydQE5NvdC1lxFnJJJDlgA1o5fsoFu8H/dfZsM4XvGcEen5bCIt5rLIQzz1OG5gEJOESXbO
yNEE8BWwt90fArskKtMAnFhlACCbA+XzEDx9IjAh0GK9axGXCFFGxvrEV6AZamO7UV15LmkCu8iX
71xW/eooqy9U98+xynawLqxd9yff/dECgnfyMWQ7N2BsKp9Hnuo3RE9lyZXzNorzABXLGdegFgg2
2rUaVbwKUZc8moy33+wNYiF9pHG9BtpFB8v875TEn6Z6kYem5SBREuHbv485x2h8hw+ieyGYeURp
Kahba6Ug2WJAPpMJjXHTkyhSPfuihgUnyj395zfeM8qmx9y5KuafyOstlryqBKoZe6z4ni2kN3tk
Z2875e51EVmhuqjDPz1puZZkxzzfYccd4IQJ+VJDbQauz9FQWwuIvvUUedOgprvOdgBe7AsndUgi
FrBQWsNwvXjlNJT6zghYBs0c+COXSxRkxY3HrTdiOPC6VmJoBHemuJiZP8df3mI43am7aE9KQNPs
igZSFiWZuhB9CyGBQCkv+BfCZua8dmT6+1rMtE/EkQMumKoXAVlCNKnau90xshiqkPLN2/6y6eSN
IcoPqWQSnh2AD9gzb9uckVQiUJBsLO13dNwBkRLi0Oi6ntSGwg4TN+6Mv8j3+r4C0NdEN6rMl2kO
5QitHdvD4aOBtWOxU627ZJEs4TveZT/3Gpyh1ixMr4lRKV/5Ma2/pjHB6K/glUW7MrsY/nXgbJ0D
ngL7IF+o50PLBKdU+IQxMT+ecsxKgT1hD2V+sgepPm7hf8kBVPM51L19fN9kFs9Eh/HNHmxzAEWv
JWEDqiXxfpUKshgTW9Y9h2s/1CUi1R+6YKEWbxvEM2ehJply+Ynod6NFYJ6n3ZHXcTbOevTWVkUs
G/aAeqxEcE5ehQLsPbNhMcYSaVkwP+ps7POH2lxlxZoSfV9SAGmqbXeChR+kkLmaqfyTFNBXXp6r
mVccYlwC6Q0jFj9GJs/l/aBQ/VqRvSTWboZeeO3ML6AP3+s26a5XwxvyMr5nt1GoloInd7lZj4ly
DyY5ttDhiS54Ng2cw13VtwUNFGTDXpdonZjZK2B6iZieEoFG4cGqf2UBd4M6YHYfzeWStRzJ2zAi
u9h/LYVRCIKc6mkl/WsmPXEvUlfTSi+fGlUAQobdMgCH3XnzAwOhagd69qXM0cSrj5dSdWUo47bA
aJXpKoxXq80lYE9M6Oa9bDUVWHUQHCCq0/wLS+pvIR8L8RgHxJcT5thaSIhPkadahPRf8r/bgauP
dwwjyVFiDwDv6DZPIrcExfyt8tYGpZAzLxru9aIcSa4dkLserRV9/1ptXE1ee9ff1h+M7cQwaRX7
Q1kWB56xkGca5MicRJn5aFDLut6pmjYoLA39lKSI4j4OB4b2C3wFa/99vajylbu4lylmZgtQcixi
4WVKCisLV5rZdpAhhdTwrI8S/lvVnh3h9u1v3GH7c9RwLaisDrAxVTjZ6lsjHLq81ubZQM7de5t3
1si55WQNxsrnqOh5aKn4ZKEEI/0dcbr2agEAh0NK0a3VA0mwl5++hp2wzIc76SG1xTcoJ/0+giJi
NcjVCrFaOrG8CarnSSLx8hGF6Kl/3GMdO4bc3BHB1nTvC7JKV2XxffliTeXtcNbSNbUTQ2cwB2Wg
Nnk4HE6Z6fM9ugF81xEvp7BO6lKU3rGh2GC2KosHPeRnhzr+ZC2GW0nyLd2Yxanm0b7xkoVtbMNA
scapB+sZOWixOdvRj6R3APqUyji/PPiX+XasEHW39IWWoLCajWrmPk7Y60ZxWwKbJDIz7UFX7nvo
vYEMlgL9cY308YPSgAP6SHNJsaionsBOBFPQ8dzd3yDDqC6+dFIEGUSiknO4TbJ3BUT98CWS9D1f
Zq+adHcuIpxZseFBEJ0a7lVH/tBHlinr2aIJHIy8SvxvtC8KFT75JSgQYfYt65yAIkP32p0bQWgx
4vmXGa6ySj1lo0CcSugFQpLh7/U661swHPRgI1ZMo8grwdl7Gd1xL7qBtpedaHbtpFO0WQwFkDo6
27txyA1YVR9zbMPh06UKOoNO3ZlTPBOXd/8/u6a6ySHjWuPw2uhMWPqzi34wnPQztu6EQ2hg+kC7
iGD2HINwBsCM0atFnnrbd9I+XvfO/UQqDqYh4OREr4+0Q9UwScmPoOcpu8q3ax2BAxiZtQkMgd3L
fV9x7wMOOuPWsaJB8Y/WosRnNvcI2ZJ5nRSIy5liao3Sk9y5Rv3a7EAZrcCU3hb1FaLHXuuEkWPe
jUbJnPmMsh6IO9VfwLZ8LO4lye6RnCV9+y8jWA5PvNJDLpkBp5qSlGFEcnKGJJ8rwcxDSCwkPlTo
0Db0nI2U2eTQhfh538n8qZitmPQMc+pfqHCBzSwbmU2dPfdIfnRfKcJhRab/7WmVMCNIn6+2RVRw
9nq0bWwFdxiUbqa5KE7n9qy7j+jaVtB2A/UxeIqPvJFuPZcjB1H9ATth9UkKMSx6mQ49DOsWlbEZ
unLfUIAt9P1C4PIutyCV1RRptPdSnjP5QBDZ9HMR1foc4wUFs4LaysVULChYduwRlwZdCD1alY2L
pB+HwuzlHQjDhy7HYZ3syb3qVJs8ZZ14e02AIz884KjayGJ650LE3H4rx7ePDQ4K4C059rGLW5xz
9pWmEQYymbTXi1jN6RQWNlRDMBuePcwPWoovhAm10bE+vL+A50YDnE1uy7RvrPPMWW0GMdw/gLNa
hpYf3zR8Ik7v2TFupoF4PUvaeeCJXvCvmb0DWXTk/3gpYnxA24vxFDyEbzq8JjvkrCMUZOADrOkH
saR/HWqHqfKCW0t2d9OmpxGLqhdIsXK8DMicWmRbJ0N2tYuaZAWCD2BSUfpIyDQMK/SdOuB2Y8fT
PSaIhLvqCN7Hx94tsQW1aBieWdtdSTjx5Y7KahGqMEJCvv9/99uPhNr4zVkFLml1av0UMX/z8UsO
W6+obSMV7tjhPjp33TxaK5C3shFQ8aCC+Jb3o2VOsie+bYa1YbTn2nv3aJP2gZCkqSGj2+wvbQXn
1V3tbIxa9k53G54tVyaTLXpIR78qDYSN9mGFFamF3VUL/JOZl8/xpLlw3nKG0qJDsk+v3+zpNKE8
C6H0RzypAc4GDZ+bG6fnUZH60IZzwmTwYSrSrwEh6gbcx6KaAzYDWWrnhHi8u9RiMf4q2vHXkKVz
QlHahN73zCc3R5D03TDdGaXeSGtu3M3CidxJo9U1qvkSOU6GNVByWsAgHoeD+io+IBgizXT2Jga6
iRmumigwpSG480Bw6ap7GmT2X5gB1mWuF/zixOocPtNpyERAHkUhXF+TpZ/RMTFxd7zIzT2OusgU
2G2iXoO14KqDbXCg6I3CYaUH+zdQrrfDG5Ptc0rzHFMNxH5jbPVNhoY/cMsaUPc/GZFD2KVZVNc4
FkaUHSk1EF6jDcnl7aDRY3ASO/ck9+r63CA25rnSTYloqn2eFJzxZldgXVvJXq4NFWGJfzwsXQTp
RBD/61Y5dNHpoyGKKEgqSZTTvVm8Un9F//yWqyDwH6WHMSPFuXpdONm2zICtcVQK0nl9EA6Zvi3I
ICBmByL8XQkxpe2iGwmHXN+odhSKfjz+rVBOgNk0c0KC0Jn4ocE/DzCQkpxhIukCjTfcaD/mYjP7
5a7+9supTEfW+M97rsA2zcowkfKiOWZ5ga+EG1XC0YNMDQAiVE/FcZ1lO83QIBBI+AIxXuh6vl5V
hWoCFBQGQF40sNaZpaLNADbFWxJQT4jnfUgqZackiL4ecpBIpkc0IiBoDOEB/iegZ1hQ1yXqkm60
SzP7gRmYx+xBXgT1u/YpEHzoc5h6uHUbwW7GsR+oFGbN81rItNJFp0DYV4RdkDJVUDCQ4GjKeP8e
hj66r1N/udtEhPza2KmccZ1IwclXLvFBosLL+OwKFy0nJoM6Hbat4RRuk21X5DT5vLvwFiztjMOU
X4DeC3FGNK2ypFF1qHHZbrt6cmxnAnvF6WRBbpvUEQgSzQs+oPRZqV2tG34qpCzsCggkXr3OzjRq
SII2UUGbPqxpPo8TTiNKdaFKVbnwjmf17vCOKqZljnTxzYpeR2ArWFVRm9Z46eitERdO4bve5LS7
agxGuQ5nsB3f0Vmad1NhF8ZI12OCIICC4GePbERB3ly40p0wabryS2ToC9vTSQPzgbH+jrrXvdYf
ufcEura9ZHU/kv15nPN496GkoKTtg73BJ969CwTrMWiKriqRjdstEiLcmeVyazRkWeYB044Jg88h
zp8Y3b01ESzcFfVdzSIdLSesvA+bLJX8sReOy62+Q0Ya03PL/ZcFz13ZSUzMSovEmLEuP9jIlZMF
8akOkj9xlu6rLk6tOIvuYIv/kPvOZegfoVm7smYcLASo7eKrQfPJ/uTJD4h88Ub2tEftHYX9lmjM
IfLMP/20sZejRSGo7d6aIs2HcOYekrjBhgh1AbDZOC9aOmMu2FrzLkkId54Uk7wcFy0O3Da8gJGm
h/DJLkmpPklgMakXnZa9YoKxCTTRtFVkeKSL1dE1c5t+3OlWYsgNWo7O5oIX+mFS/SmqenHbodLk
l607NabpB2/+o32fxNWVPoPeBTSGebSXKwkTbGBK60BnRfZ7Caw21EPMw6AetUksmEQKY8p+a7Ny
0KN+EvDoNZhQWB/eruAEFyKMzB/ll26IRPwCsCDBFrfLvbXR0Qyp+NBEUEgICNshtH7BsA3TnWoD
ZHzjVqUN1SIFf/rA8/FOyQl/MpWNrbnJ+oze8KibBJisnIprVcXG71JWh7sEm30oqkwVVSVrPZc5
CxOpFniFesNVY5AeTC409BA9xxeldxswiSkGjcgtSvVBVjYVD/aKm/vR8fuyXk6iYqQK6Xm6jVTP
cmYDpQksursD0SIcQtBikrBTBccRg32n8uL2Mwq+wb/7xQnU3hhdts9j3xzCoxpLY6DKW6X1qfm1
HQWR7Bro/FUQM9DHZNXvZlL6x6fW245ZILK8GbPWfXLMkJCrlmpDNlwU33CcPJ7hRcNB7jcSa9I3
mddIEpFfUFPKLK0fV31sVFBIy7JIg/x/cBmdchzSbEaJJbDurV3vwg3d0o/0OXuqtl6EQeLT/fiQ
Oyvk1HwWsR+XeRmQnBAZ5kkZKPvEQ3MtgiyvxWNWPNQUdwMUqUmJSW7naVlK1hIcOvMX1vFUh/Sg
ftsVG/6SRTTIl2FeKnKtyvRixnXti5laKu5ntPrlKd3+LWiJuxjM2hcesvUL8OldCRXSo4tqLpE7
QGG1cPjvkCMUQ35/A8QnfC/jfvMTk+Syel7A8JcPRjrkACnZ6/bXmVYJOou+UZLuxG4V5o+b2CAv
g9tP6sg7HmYBHkRzGGj9HokgVD2Lrg1c1cyEOTWKwYnqPtuHopNim73GMRYf5vYXdMjAvd4v/704
/tDXOLvhxd3EK3P2HfSiDWFViYup+TtjpvDYuVKyFOxj+uU/QdXpddADMFAwoJ/RtIsvmwcDYY0K
aUzPSn/T4aoWe43ReNUTk7igZw8kXbq+2xcET31dLYQprb+qobS4E+oPNJ4NU+fF5nfOSGZNygLv
DIKW+6jro6OcyaXbCyumb3fQRcfM6BU3zF9HnZWRDRZAkizZkzr1QaqFVzIE0IfYEKqgLaeymqnB
uNk+yQkPDRWF0wsYDNkF91zyd1O70cG2Bd0colX3LIlx2nTiofyRiqpm/U5X1NdO32lLz665QZqb
jGbY3wCFw0WH+1kl5WKh6mXwjSAi6v/70XZWMkj67vDZHCsBPJasXwrsjxRtGz1PWgj4eAq1P0X+
XPMfeyjEwChqYy82effB5M4GmR2UFE09sa73Yds2LLKZb4bCLvaZ+iedyv+2WogJvXxHx1Bmn3rz
MBy57Wq1MLXsdr9680gxWrakTfISGrYG6MeBV2Dg1SOHxyTTl3Hfc9MPpoLHR8YTPLXSqcuKjZWq
Zht2HoMDKbZHJq30KeMHk3YzrUrqJizsSd2+AZoOzfOehJiA2rtgOYwolKLUgM9bRrXKsIfGBs9h
SGcvoFoY8F39rGb5LQrR8R5k14fpHQyEjbMMwZ8U66ygIobRs3g4futzJMdbc6XlKBStWrGQOBRH
x7eVdelhM5HlKaLE2GMa3X/54LGaduLo8laX1rCxjR95FPoEvlunaVapTFL/+3i0iiEsOWK4VCoL
ZztbiD0RqraIeA0OVmCOyqgwq3UA3Dgo5GmF+jhApCkIXKxIioqHruIE3z+7y5Rrawc2r8v0MwqH
HUBBHJLq01n3rl+v90JQL6MeyymYoBGP6SCptFNyCMhyz8shjwwXNzptK4s+wcY/Wtu/0aMhMvLN
6dm1F70dkMHcwm+L/SkI3uUfjBi71m4y1Zq+sLvTerzu842EqFBnrMZAbJyAUqwcbWy4JDS5eXDC
kbxidpgua0GTHEw5X0dELQAlCLNFSn3eqR+cyFzCf3uKU5AHf+YqXb2wKYM4pPIBQ5tf5MKwL6AK
UW7aYLUSh/8IgAjI+89JtoZTFx8Hp6pSFc1HaeR6fiq0PfSOG9iI6K9i+BVDPUbTKr8Dc8J1+Dsi
59AvX4e7BCulhyHKwLwdM1QCLcJh4XNstVwk9nYJKRC74GMXhzpp1LfbYhQ4iwE5IsI6mx1IQbuw
xtAMv54b48V0msW4kns4BHys3YCVa9wQSHxGa86ZLSk6a/pxMu0/YIEY2li2x/OaDuClHkC1WHcy
ad1cILT9MrUeFuLC+aAWjIpBll+xnIFaH7nSjpRCfun+i7BsqGh4U6oOUsTjFQCKICnzWgEw1HLU
xDLuWDNP+2XHAozIzohe+PMa4tNhjCvWqJpi6WA98+F897uBIwILJ5NL6G1bwTUhP8fQgyxJptDG
EpzNog4br2e2Yv3sBAvdqxK8+3tgYWsKh/7R/7bq5YzdZ5Qru6jEgEozXEAnyGCKPb+7Wu5r2P8N
vXkrrPzWc1RavW/ht8NvDu7SPsA4iYYoobWMKEPCRazU0YKkwEs4NOtr6TCv07EnRxR1xvAmKKc3
7Y5/X4rNHs16e6wT+vuQmmw0PZrBNW5VfTBsdSwYpVodI0iYc+nT2KFjwAe/G9LGoesa/NZuol9X
3h0NUHjTE7FMrJblECPF+pvUD2W4ZC0OdFu2p6W1iazjY6FN0tmsHlhTUX2HAxtgST3EL3DPjywk
4HNwpsA8PFz4JBPFX5hLpKdLodf79KCyqsTWJbP2mxz7ab/E11hUub2YaIqqW+8p7psHQVtP2Bdu
SCJHThT7sIHwUUFjdw7QLnsymSGOqBpgb1CvRXw90JdSFtKvCN3uUN8llkPHLiIsH6rwLFVYLi5f
FJ01dKummK9/JtFKvtnmq5ZHvJ/pszecgm1rYU5HBLXUjoIzhHvD1lG5fnnx/Df5QLO8qCYu3w46
91iOepopX5le/iDJkmTDdlCCc0ekinHzKbBfh95TwWcr41Yev6yEAWBroAQpIB642Psv5+aylRwM
iAuvXh79HD1T3q5dLTDllkbwRiJdqUfd8Iv0YGCP7sR1b6qMgjPoJr6vnxUGezWFLvphilP69svG
BoBMzkgp0If/owS/mws7mksbTxQb35loyzUvLGVmNoyVo+r94zfouJs5Mh050bbEnUaRi7iJZuaB
EF1jD+y1vLjlOcxrFI3MhzSmviDGMp0C3CtVc9H/Gs0U/KL50Dj4M39k7K+bU+CcXm0Z0PR1C7qE
Hlm62yJlqvIxxxc6RvpJokEODl1rCYJ4KPiNQEyQOfRsgQgi5xiNHYeM8BdnbZBqGeQY0SQHvdfg
KlLThDTJa/zL1dnDjB+eAqUoTOUQBqp/oW5dKAuIlb90woWsLZbVkLQ2OzIKZbae+dTMqaHyZkso
OwGD/728YpwUU7Q118PHyh5NP5iTOlBtetng48TCJdNdpjmeNmlr8fwLmJOskWZ9TbeS0qCp404u
Pz2kQUDDwXgdD0yFazu8ELd413Rs6cvwZBVkvIqjuzzYTapaiKP5x7sicKUHmSfQGFugB2U0Vo83
i4pRQbqT+ejJzigzr8KZWE4eYzOqpNTH03CBOJMhhLQ4KMDwYDtfM6gMvVzSjITdhLsPrfG24yAJ
JY5/NraJoaJs9P2bw2dpG5VHOg+e2Y6G8zidRfxWrw+FRhxjY5t/HjFrg9pOXZ9G62djWcMJuhwH
kEnNbxICCjvb1fNDzODrhR/ASRK+U+zeAPn7ydYjaZlNFJ4G4BmsAons7r9SDDQ/JS/lC/uZqQ69
2Ki2IuwqxOF1ddpKlJDOb1GtG8AaoRC7gGBEQljfldWdaWEeTcPPwS/+h2W492HoxgSvATgtc3FH
Bh8ts8CEXryWG0r/JxyDARUfwHlHOJTbkiylIstS/B0AsMXs4C9Ksl3CcZjuBV0OYWO1raHRDKRX
WhuMRtueJTUfmhDsQK5ehR/AwLQZjACL+vb08AJYOe2TfehiNqtJXFKTOlxI1FXbF6E6YNdmZ0es
sG4qb3zYS9jloWfRidz5lb0IPfCXmsHo9+wvUEnoCmqYgf/CYbyPRN4CSNfhOo130+k/1LIXo3eU
jJsGAGHj/qmRjxW4naqzMFlF+Y427s6u18zUKSF+6rytRsUDcu2Tj+LaxNtuTfuN+s3+dgVCVw7c
A3J4bAgteRUnG/i7oVD/maNQl49gjeZc83H/1xl0ciVelqV2/zSvfD789lqzqnZVD4eFOSGClRaL
tPNvR2JEM8DhP1ZQYoZiOx6YxSRUjrEyQho0S0tsusW525h4s3qwiZXEL2efmzsrl95uTlI9quPk
EQp++gGBR5pVA3V4xRHTnaAIILG04PG7raB9iPeGKdQ3n4KRN0i+S8Nkop2PlpWqUxaJoAGG9K7O
wQ4HJ4MOSB+Pot2kfyO71XoKR+b7ZwYfREuu02QiDvnbQFVPJEfKRY/0riX7vQQBbIMulciNIuSG
bszWHCffWW40Ptpjetr7yfwE0EvAVxyEyFqEmKCr9mCcrHFBxup2n1wjIWxvHM7msXKDkqnP20B8
BDfOum1q2ft+M7o4LAoaLM9rV+fRdpYr8bo4vEb/zhUtCd8fS3YmaOGzz+XdQ25gw+vjn5URUIoi
7uD70bRBjUCss7LZgnxZxINxtOUStcm/nzb1BM+P+F3E9hOidHZ0RA4Apv7BnyWky/jRrFi92yzE
d+oYLeEbgsk+qwSQCbE+3Fz6R3aZ2IvAU9/79LUteft/GQglBpGFn+2I3fC6oGSjqkplaof0y7F2
RRRA+Dh6UqAi++CQHcIr3LqImhiE5JAt+K+BVMI2yEiNdBMzaWMAHSXOX5lcP0iD+vr2F37LnUbf
iw31rQP4BxMbF2A9NWObyued98/b8XWbJDdXSf2iGpm/L0xGO6P2wVSIK+heu5/oJ07RS+xJUL3H
RxOU8BVbnxAKoizBItk52/uCRHS82G9a8raGwkc0lDgBay/+svCMMn0+TGCGdh/S9afrCp1KGJM9
ZfQKZF9IqGfxJHGindiD2OxIimkxv7Q4LAx9qtYnkYM2sz4Oz9siGRopuK/FRZdz8efPQOORShDa
0FVrzoS9ggW2xRuwmlh636Mj83/yrQuMota4jHgfodcwu4EiGcXMO3TTpRqyQ4NxJHinW2xCPshW
OEZOlf8y6TfTeJRD50yu2HwAmE+RG7WaR88QWV2C4aSfqF5raHkmyFA693qxMrv9m7V2RDZDpunA
IvXC3ehQ137/IdqYSRRFslGYOm+vTpHjBs2NY+3KWo6HqqOVMjVDo8j9mLKuiVdwYNDL24clMAmo
vj/rYztsWASTcWMrY+bStnL7N44bhCMCF5ppz+E7sNKDlgFrbB7lFHj71vhTGa51g+nthqa5mw1W
/eRmT1hHEr65t0c9juf6WgHwHrP6CUuSoTtHuUF2ydJsLxkoSwZdcRofYrK3+p8ILSy6FNY4osfK
CE+ILt6d79SzgFiPQt/6h06WbPHbuE4+9EuIcjAkjqcIBND+Qd+4WdukVSUkHCd29YmVOq6nHuw2
pdr1g32ifl3/yp/JH8lkHCQHbavM04tNU0xk3gFO2NSayl9+vF+19nRseeF5UxZoTm4h13ARDfzx
eXwQSHmC2ipSC5PSzjRtNzqwkPyP7/Dg7PB64gM9NDWbUYWbeXflHc1jzy7ygsHu+6KTYg9/C4ir
tUJRWFYCgjQ/JsX8U3eWaRrX+VplnLF7bmmLr1Xw0B4vppR9hQ+U66bfsdSPU142GLKN0/nKvL1/
itqC02FeYWRLgidAOAhMJ5+B3K7c/woxrPACtXJD/fK+Yc8/c3kM27B1ok+EpSsQCKGQagvSUvKj
FuNpJAuV948BVjTyBwl1/cUWaSFncxxBNCs01gAjlpAkcULf2VwszfOKePknEN6jSKmrm0X1ie9N
m0RR+oGCsOJVdhRtPLaiqtH85Psc47cfZlCvQcdXP2mos2hYmq0pOyC32SZqAnU7pfBonfuXWB4K
hjfNmCzfZsTXYnF1VBoG0sB5VoYtclKxlwD8UG/oyfNnFunvjpYJcI1TyXZxkgTheyHSsSSLQ8rp
adCkuEvHHa00aJqFu7m0+1RZrKDiWJyTRK/Fk1HFVeL4Uu/vv4hwan5ksk8LQB7Q0sIWwkhZGsa8
n8enJUs4xJur7lvRFP+LftdlGiVp6r/gABFMcxfErQ+E4ZRYfBc5rmwXo3Cmq4KJh1b+TApAsFoG
I1hFN/KqNdyUYZURR9Z7HtyQXTsenzpTzuV5xg3TOKBANyR1qTiW9hCOZf8gfWpJhda6mnkMzxxe
yzOjp2F4Fz/tRx3c7GttvOIODB+xsLtChQ/ZLBAeO66x2FcliPhWUWyKSGj52NKjbojqpTjqGWH8
QfJUvqu4zmWJZP7ExR3D9o2EIa306CtUKH8DGSTBKLQr0JFw1+hehJ+Tx5Q/dk6lgK1hiSszqaSW
VuDGJqFCyl3vui9xR5WTfuyfXX+E9f//xUyrvvKW0ftrPgaxXKkJC9qPxGsu9oHwmAH3V7E+jWil
dfAqkRxxJFpL7uQ4ii/Z1aUcHwYUxd/dooozdVToom2khaOQHVTL6n9SOLmFtp3k45+PczXAgBJX
T7n4V9pLJfjrrF5ilg3vfR5cM1SgP8ULcbQVEdUshahbU1x+KYRLgUBmlVB2eYCGDyQXCrPP8Ulh
1s/anFB0DrVyVHWaGSPQzEzboU85Es2toJ8lwOEpcdn8P7yx1/Bkgc6JFW3IkgbrJjzjFckcGxhZ
8Z70JgLZSCZnF2oBzVQGGqEHgQ6hpJ67GpHCLMR5ShNqO10YMViJWV7QOJ6f4wLv0rOePmfOvSbY
aGmRWS+ZcCH5SPOy6Y40Zl7ktSIchBrypUpdnqrtVP2BYVyiu3hSRE+5V8An4NElCs3Ob+xngx4+
S7ZXrhslLpSpAeAJ6rQgi5IcMUjjtTR0+2gzJARd6W5HlDXv+VBBKLpLDCOIVNblAbokopRvcTJO
aEKfL+sfTW5MVtazgvAP186WBS5XZc1jErxVs2P8JDVABKhEzbBIx40lI4VDFFJEAjT1ay5bp2dm
x6MdtH2pdU8J17ez3Z0p1UmncosU5zpeAWYCmPh6xiaHhQBz6aZyp01dVCw2yIZpv+JSUknyXkRX
gCIk0w4344nCHcjETI5AxUhkEiGHeiTxhMvaDoVNIOtjfM6LBfb17bG3DxbRp8l1MSYuyMskdR0d
c55noiDeANP2LYEQuwoJmUlsaglNeV4uEGQckuM9n72YcbLMoqcSuAl+H6IiGMkpCHATkJ0XEOsm
h7eAOlYeRdxRb8N5SHD6yLyeiaEAOok7NdZdZrYg63h/KB1HZ/h90Ru4HPTKF84GCrROlngaq8OJ
+dVVDrnMjUu61Z//wtfpH+l2I2Ill3ycyFPqwcgj6TSdTwHJOU0xzPuUHK6308Z9h8rlX30sMTwF
K/W9WUCnsyrY5Gb4PqViteC2J9olbC4LZXuYWENJv0k4E5jnaqALpIALRcxE82L7KT8EPUMESMw+
5XU65HUe9QCbBO48Q4UostfX4jYNn+UbBRgl293RXuAeWbORp3wYojg6oVML3gYrBWtHlw6Xzo1j
3I8jBNZgao/dcKdgrIyNBKuw7qMvANm3VUKNnemIF6W2enoyEkNwIVl+TmOXi6jPhwUxHxwycJv0
Sr+jQhynFcaiqXq4HjsAbv+DVwThYl0zsFCtu2ll0CwakLgcBzd5m4TTr1tMbl488uqCViBV0Ryr
qm6DuW2TMUb+QznLtscxarGEatn3FJ/hle1xPl7ddk+WET9xfaIjiU7c8pQWRE7mc/kW2LNCISib
Q2FdEUpXcDwCSgs4+L0hdYXi9RjidzIhxvlkE4rXyrqJ3sJwI/2nDXw0cck0PgnFaX09U47EboGn
eL0Ue17kzUEf9DHT1OV4tCDMfhTPIqcKSFpLzaAS9+PsTTCHWzQo6QDZNrcI63CIyk3Df3M9KCYx
e2DQ/aaapzvj+zofQho+p5lKE6fAlu487Ir2l9AOXPJrlkp7mBBytMkik7AXxfZs1LieRtETFdOe
CFG6+zsqubg0LYcr/XXpEc+gi30yS7wx+rnDsRnYFqk1MzDCEcpJuvu/ZaMLeE2/THlQAvMhnBjA
+91R0VXsEXJdnHVmdXWHThHgRlnNuNEwcZFggA6v+mxg8nT0NJYlRNwfo8btCbl4xX2tZss26Ui+
P1/DnCuYJ2F/wUdZjNe0UBSNN+nz3UqM4+sQmLlv5rlPDwawXBpJaX/0dabgI+qITlTqo4ZbfX6h
aUKTeUTkSGgMcrTIcw9ipvFpmlsQ1fN38XJcgaHKJMZxQaKvm4GSXb/t6iZKwGxl8KxrAukVavDD
mS/HxvcE/bFYYHZ+nKf98vodKLOyU0HPTPUB73vX3xln7C62VfPcWxDS6MUvOa0U1V2KLQenp6/k
XJLJEvEbrX9/Ta3if29GcU9KEzAm42Hz6F2tVGp3d3fdLA/VWDxr+61yyGiBbXzNWamdYkeNHtHO
Lic1BrLWTU8ptuGO2RtkCzcXlYxcspVUA1cMDLLP9EGUklAfEDPaUxZaiyc3IMtL7QvFwl27inJy
xh6mvNlkPG4GJaKMSBEWT/FhrQ3ub7dkftujdLfNblAQvMPcJzzx/ofs5uDY4N8BDrtK0I9GliVn
890F4/PQM8H/Ig6G6gbKuuZ2zgUxJZd22mo8N3Vgd5WIBWQ36L5aRMSiHfPjh5MN4/DZGid9w+YV
gPMIEOV2ACZrwjuNkx89w4Yk7awZ7kBeWrz71Zp/JDp2F73eT4zCkslAtssiet0V9QCGoZCqBY59
s98xViLTohHoxUU1kmWtXcl8QK+Uinv7K/IyBDFbmjhMXpfLArihrXOXZjNEKUoXM6NGlQiFKvjf
7LTMUQIC3esOJOCX1B8eURRTQiDV1bBDWF2XFcXhJl9Li9qn/oJ+778Ccrffj+5k4vE3pUAOZpiQ
KXDsUasJeiEmH/mSPB4hIdwtJCRYUD4uWiJ63BaEfkvaVZDK2z1IqHRJcXRtc5o5N/RERoIivJUH
JhxbTvTdiVZseCCWOlfhvh8YvvfPxV4G2IwtU7zP92FJwp/Sxes26zjHyTTxPsnQ5dk3VrfJgwKW
gKI8pjPXs/1GPCWFJFLr0ybjzvn47CUyIwo8vcuH9yABRxr/mR7E/2Jn23MvjZcwxSHbmtOubRpg
7+DzdLhklHE0rF43Fp32P77X/Qtsde9CdjroFYNbKKeLNet6eobXadnHdbtwmr9mw58yo17AdaTz
NQycwQC5x5MH6pcWRTvNl4nHKUKStd/OuaOCGZUfGvaNXGjjIM81QYQS189Q1vUZlvlZKByxXN+8
7vF6OMs9CmgAGKh4nkmC2f3j4CzU8iHLDsoyMamsHgOAlwyqhcD+LnEE3fBVbudqzIgS9aIvj/mm
0cgzu9OhcDtsE6x90OVuAR84L0T0Wee9P7bLsTsdiyBtFBYBtlU8El4ALtf0ULcJwuyfjauVD3iQ
cZDmZeKVw9qvChcTMgiVlG3H8SlHVbsCqoqamMQ180dsMQGy44Pt4mIKZXUDpsqRJSFNYpYQ+9tk
dHhGCLSrA/A7culZvC6vGoO4y8r5+DlxdNwr2DLTG91qUyWPJmp8jA6OYdOLAgncV2nBdS6OVOhi
ZhkjDazGhz3OoHSwLK8Yyj3djMrEuIUhA3+wjnb+PqGE+32dGCASiGlR2nXWHGscb1WZnHkKHq7l
iIgAjVwnspL46oZAm87G2sp5HhaXu+4heDQ2+dy1kR/i/uixT3DOV1apu5FJ2OdrkFHv+rPOh4JR
i3I0hkB67XX/meWYI11G8PrwBMW/UkQRa0Q1HdgkfgN94A3ilR5f6V8MMOGNOIN48YR6iOjxP/Dc
N7c1VPVXM3Tq6JQoVWQ4PNl7SZfl1r4hpsuFkVBRiSTbkh4DG0GmIz3YKaEc/iSoJ4ZbdFUpMl2U
XeWf2//Sqe52s7EHJ3OQGTSNs5FcMx6vwS8P3TRhNcLHWIb0nCDWcQumYuoRJ+lVySPN7/GRU63g
LIzc/YHSFp87SUs9tl/jQdnOhDiWZzdOy4+4ptJow/YMPHRpQIQGIfHbz3zEsErOd76lGWSGAqDT
FB9RDuoj9P9dIf8n17TM5qPsrrMrrVk3dMtIjt8YXGIHib0pm0U5xvvPp3LqGC3YMGqf7KSdwtxu
Z7D4k7eul6oKiMkzah8AeIBokuggvxHogAxNx8EEuDZSFz6t4yobrhjxtxqCYsUdJOUGZgrKtBwf
ewGGlbiYwZ87jnkUcQpaWnOuOrZSNepZHCC6Bnzx8Dna5cvydSBHvVXZI2D2ulljiBuYvAd0YoS3
na3Qiy0S+nFIaidRRYlDc5V7yYtNTMOBPIyC0x4RbjIevv6EhmEJ3/OtgTV7E5EaHXI9v50l9HbF
JiVYuXBzWEDlZsgUp4kAoP8z96sMSG7FfWdYUTIfEFIaPAcNjCThpKIGv8a1Jmup/VmBWMv9DodA
XSf34pM65GOBuafNw2q0zSuNxLfKhrTtEuexj7TimguszREUs8Uuh/LPSNjxYFsD4RXDbKfNwCck
DHVnYzmCSG1ySwyNMzdrV5IE/b4U8caVjLcRSp5gXZWQPl6c5Ov6RzCazq51uGOECMdFOw7f5m+b
T66m1aNMVtcU4ebsku9Dco6jeKBTBAf4Ki9kYx2AL5ooQOXKF6m8jYTvHLUcENe6BMXE425zqXcC
LgN5DtGJQWfkvhM3pR1ZsAlLto0vjXmLd3cPRSrlaER2yIr/O4kDDBsopO8LLORQ12FywE8041+k
Ncqb16aP023/89HqOIF1UvKxQWABw6T4TqG7Wy9JOIuVcKYHONbG2+xv3X57LUGB86mhATeZFjWC
bgYulmLWWqmpdhCHz0qB9pUev39efsyRaeaduxejndokecxNESQ4AeSBP1Soq7FyatPIfDUsgKmZ
12vNPVep6PJL9tbxkqfoDmKtZhIPskvKRclWJBbdeHvkw6MV/R0Y4gGKEmkk7TPDkpyWH1IBjPqv
o5KPHMEhPh8QGNQq3iypNmN9pv7La3+08UhvTuwa+GeM44RGuBJDbeS/alh61AOZl8SIswig7xs4
FPvpCSZh+nxEpDUO8veThgE/odaFLtL4K3FKwjhzb5u/TW4S4+Oc+tCuPQ7LcG4qv1NIQsYlDaUS
HdQDH996JvRE/z3Fj9Sb9cQQQ/OPr2JxWYo5Kchvjpqc+PkzbFdRtj4foq/PF4FvEETqGGNUT8PV
jizAhnGIhYaTzRXjfaxy+CMpw9ijxCDvPnN5TM+l48YcIU+Qd0Qkd/jIKlr1XknHI0YLmEWvOTpP
boppmeFf718jkKqDvlBYI9fvQm1dGCjEK8dAF19DLHrNS+vccEVGDZGXCBjJHf8sv6MYILLmR27C
WwLApcrscO8/BN1ze1P1Edu/+GQVFm6q1vBmkDsra3wL3xUDfTf3CajgBY0Kg+Eo6hpSEKzAFqxh
5IjHYFay6h0vCErTNYAyIz5aXGKOqygn0XjQoVvf77vhAlcnhS5mRs64Uxdpu+4Vkcp7MSswyfU5
KRzyLWMdeSltZQ3xWRvz8jNtv9KZLMPNZSbQyTkP+/2bl2lXsHK/YgWK63b2un9wGEazzL5H4ce6
CJ9M26WxGQEfM7IqQQLZNvk8G+XU4tjqSVm/leKHRj7gARYHH4aTD8584vNqrn/eiwrw3zwHqJvi
aW76HhCCJT3yOwh09TDzYcOqI2doJMCMSZxMnRjr5trEKQbhIvsldSL2Qbxijg+ienuFA6Q3JxVD
VLqNSSobbN9sCX/gCQHRPeo7JIqmN0aT+PdgDKfeHj0g9Pe7VvFAvXEAnJcVDpNeoDqFkp5DKUUO
PtRMpF0TEElDtqy1TayejTChpT/xtLFA1Vk7gr5Qq18K/VHWOHNC3ceq4DQLV0Kt5W7npnuK1Ujn
ttwwIBZau9vAiffGN1s1TkQB2hR7AdzhRVI+IRHyQdZda3mmgxIoGAJaeigfP5op5zJCSNrfpKtL
vP6bIQvximhBpb2oWpsB8uvz9Klng1zb0IjObfK06SvWAEZUFAvogHB0SBmejf+4wyJtlzuakPsD
SIOzfl2sguYY8Dfs2ZlEJnFNyQWysf1Wu4gJjVp5oc+TraFN5JEokQbvPbWU6OyuQ/LyI4uM4x4W
np+mNcIL1BNSzPURKXSe/D5Dqvcm/Bh5TFm3PuI0131fdspSErzOdOOzPfWo+hDnYtNe0lF+K8WE
A09RBYtqHCtHD+CmDGg2N5zMxWxx3O5Hzz2w1WxsX4o4Gy5oWHW40EF2KHbcJoFMIG+LpOJVACX5
4+J724VYh6lt7rx0Yu6iplkYBjOtqYaqySqNLcRiIZM3zXAO1uuI/G7O5x0UT3z+Vsu310wS4qMX
peetLPoKr/HQzh0WqpsM5BVVchdrQvG8fUJowSbE3lrkIIxmEcOgeOf6oOPXU4FNKbMYZECakXTu
X9m2BqhcQ1rCnM2LfcubTjCTOaGMvPIqirgnqMITX3ocm3gQcD/Y/jZJFAD0G20JP6jey6AWtBnw
CviZFHEcLy9xzGhB9lAG7gfP57sC9s+iOnO2HCwm0vq9oCk5F7qVV6tQ92z0BD8VMjj6Saj7lr0z
5bSdFqeUBYYzJ2k3UU5UNo8jyZX4p7BFjGzgH7jPIpnGBBoKBGJ4bxn1u3rS2oba051Z4gZFoT9E
NRXTtOSwhdA0Wn47qmaHYoMaRCy5RwjR2iixXfBhkaP7LUBXhgczl/WNygSoQzx0WH6W2lMrMtpa
DTyOM1V10GSS75CppsI5K7W3PRHittORSRW5zrMinLIddpWrsWgw+V/xmTh4IbhlCZZHmMpTdYui
0eYrxMuHfY2gyz3nganJSm/rd+8dQt9ZOQ6+aiB1dJOoh6yxuzXscOxAis1Hopl4b2pYFoXzZ9nZ
e0dbchTe2NYz7GIOkhhjZ6yz5pd1D4pG6pT19JBYFh3zetpEjBc9rG9xIEYOJfKiJpvd+O/wOJhL
BF9/R1FupA02jmoEqYmOcXaBLo7ZbGZDTwf3EtT0yiguNHXBTBKxQFWmMd7tHskPwkkluHaRJFBC
F+frrj650o5zc5/V9llnsNE2unYMoQbdMbfvyJnyphNPl3eZzpt/VxkwRE2+37sQ1VfkrOhUFhcK
Anf6N63uEeJmRTlidcrv2iVmlfEAj5qCwJZA/+fS3JQTeVWGjwAZUGLRK1E3OcznkWSgul+M/Jic
SFYDAZkSOBIFSlJE+X5ZMm1LnpzvFw4iuti0RuMD9/s8BgZWP2PKfpsbEgjtZkTXOcnYPvUorb3v
g5rySVEtkwuKAHIzIsZVFmL0OiUSwdquA20pUjy3F1A3CwmvNnhEd2/dPVtWj+vyuQZaJAJgzvOJ
7jFiOrw4o8mT5O1VQ4M5tv6zJti8b32p+jizWJ4hKY35X9I6zz6mRby9VkFvbjh34UXVthehKzdT
zG+WU50ZuRpi6aLskm+rIO4VISVH5mc1Kd55fMCk8il7up/7ftc+fCcDMRQwhhNfxTZvyVeUT1YP
GEdQnk38sqccjXemB5Dy3F/LolkmVrDCNzZ6xQyxF2tooEZ9D3PwT5Ol3yfR5rWKUCYqMxb4RdRf
LEn9JVNcE0YrCG153KcF1MJ+2CSV0r91Y1QP0epxbndKOBjdxOhPk//BhmKqb8zkgj/aeVsZ9YUY
M7Bk01JGrV5WsWSlJ8eByzEhGFA/7dgkp1iH6kRoIwkWrSi1hlf6unyZOLZCj3ElIMv3CZD1fLXm
sbNm6zY4CvPKZOGt9ULVzh4kq+tUJWr3NYEUh4IC1ZKJIFPAEsvnOfl69rf92SUFeBLpVOFODxv8
1I8V4qtsDWI5OXvqeMJifcGadN2zo8TwmVHfyG/TWyFUiyyDYKae16BfxiCMKpEcrDnLmRBdIXdF
5cEKThacmCvwEyAQhNJkq++2Q3VXKRcI0Se5XK0j/nViPcPndCxFA7ze3ZchiioTl8XVEFNAqtJf
mgqppv2xIAsgOEUvT/pevspZuo8ENunm5C5IdviKsuQB4gygETr+nAUz2dttXQspP4Zjg8F56UJo
BEucaM7+QBwyD3S7lX0d0eBmTRUGJJeQNT3dpvsExahshZ+BN+sZZna0NHakUqN8vD6c/RfAnhel
S/DtrkGsYbJvlcteSrdxgZBX7UcdMCrSIA9Xp5+vswT6bvr5X4HGXlFQF841ZAnDQwb0krlovv3A
02tzxj7yanuhNNke6d+KMMfJuIOlcg46aB5/MN7gm/e9Ti8uPHOXhdnlQCBBFIcSbECdMRbUrf63
1LgggYFMFHOnLsTVgpN9AZbvaQliK8ipYy/2qpDCL7WW35H+ZHh/+uJ2gQUzL1F/CseLpnqOEfuJ
WAuricUe+SIvarsEMcmama55P9JgQ0ISCTvkPpWgZKiAaTAtJ3mUb4ORVDY3Hb0UCHUeHek/mGYO
O1UyqMgdkpQrj2xVvTuMu83ekjefU5T02HT691lAGYNV6prTkLTm1nRPVvwNgQQkta+xhpmCMn/V
dWr5TCM7+14UwfTX87GOih3QzP+sI+d5Q/r/RD4IUd/YZkNfrH6cepmlcdyvWQnxouonqkUnJK/q
6fj3n4u2qJmLKwFzUlzCd0b9xmUQIhIroy5lK8OvDBq9p9tNen0mbc174kSXR/p9m4UBiFFkPW37
UNVm+g8PmzflnZtU1EKdFggZX9ZwhLyr8cdKwwK6rzMSbbgR89NKuhCpU7zCS1w6JnCxN8F8NUJl
tndVf4hwLJRJ+dyPchh7xqQKcvyafCI1f3GQVeGe3wDTHijgVStBqgE2yUJ1uqU3e2blV8g4nR9I
WW8CjZRgMPcciL0bd9HzV1+WkOSKQZTlTTlUFyGN0xF0tjYMLVcGqbpDt3aNYx3AOkLW6C2E5atm
DiyPLW2wdzWWr0fzCrOffiJLiMenpVRcHX4QdD/HaBwxuDS3VpOD7v7i91rdxUADDK5XVUHPHn9O
7cJbU6GoFDS6vIiOmNnmhgFzx2vkqsIbrr6gLavrHmDKlLSecedzelxmimhYF3VpWcwXM7x/kjGJ
/2xj7iS51iI9zK617cdxjpeJwRrtMjtRvn5papPVeSitFPT61iDE1+MzbtBJDHUxDWcT4fiTKV1R
RxHXQQFK7mj0IC4JYF0YR8quP34p9Q6874xPjsMKdwynIWBMbf/Ai/foxaKLjwEK+ZCkr9kzYcF2
Ktz3VA907ozgmbfWNw8JP6LkWgPYRCg9dno+CqTEoKIeXVcIHHVDR/4u0nzPvh0GxGt0IvQI4/C1
FEV9tRCXmMAbYi8/vZ5pkMjYcGO4ffR5ZYbLqCtbKb4252M+bl0hkud13rMLKoxe2RSsIC8K8jLN
rRRHjHv5sl8UjSZfcw7kH9M0/bdGyyTPP3ksTWv3oKKsGcEIoKc3Y2lUtVYY8S/V1z2rOyCksva/
x5PGVkbh7hH1qnrdULDcxu/4Sz7a1zT86OM2xjXfRRfnT+ijq3eVXaLDynTwMMrXRgNhOv2use5C
oD69q7osQ6YxEa8trY/cRo67Y/2UkAxVwwPy9/DBzD2ZjDqjsg0RYgh+S8z/Lw3i9Z5ePkzoDfDu
SYTkcPlSTV6kwzm/uEkqyekptCOKCiNW2KMftD4IVXsuAm+k+kG7ufx9VZKxfdpsDfVtfyVNHlKJ
v+6d2GYKDBj1eOQqLUC6PoXxsiXCJk9/v03TeeCkiE5r0scNxYXC7cH48LiOqsaQU8RoCpY2a5Xi
M5c22DV5E1W5J89DflDmEG7Kxj+/5YmCtqasGiXkKSQe2RHXxh9QTTpUTroeZV+sx02OUvJRuKFP
e7iVV02Gh1ERMgmEXkBvjaHI4Dlf8FNJd3IdsYK5GQxtULF6mGhQ551HeYyKT97W4rdu4h+NB8qg
VikUoW9k5KmBJlAE7080Ml998av2u3el0SDD4V6SyiPRLHqAj2RPJHbCHyXUF50ENgEdO2zb017w
bck3kM+hmBeezSj36ys5Q8QN/thakYYsJDFSbtg6bcL0AS/BMJ8A+lq0nQ/2tPusUCpQwJpuISMM
71uKeMV2c7mSUjreMV5vr9wZlvEjN+7fPyU6NyyEAxI4rcIJHn09GEYCkpg0kSAwznDvXRWR6AsT
2IcfKI/usgmupykfy/IeaG2b+G20sobTscM24AwtIMU9drLZv4RbtDagmHB0hXzay/XfQRLWso3S
C/f3JeSM5OFs4JsB73TI8F3pF3gU8Hpge/fV7+BMs4OpwnpiDu9aEh1bkVJKxrxBNk59A+juax1i
lMMGECaNLuYVfiYOLwgScYbUCLKx5uDjPo3e0Alfv0dWp1c91i3KhlTCpc5UwHWgM/pCVv735Anz
esqWTFBvi1MJ528N1or1+BkiOzPoDJRrtOCFQhcuaONb4E9xh+Mhouw618jNMfXaA/g9SRJMa6Mm
RxA2dhQl1NrrcduKdYk4MzxFXDmpY2Wg6MRKG+mu0MSPSWOObupL8CeqtHJ5VQetpAuCe8+yNsUC
F5XhIwCmgFLNNdAWxqtmkqtIW0kDUuXMw1RAQBVIxxP3m94jy2wWrhXDKXYUjAbXclCsxFbDcyZr
vTWhkCxxXomvFRr2Qk06usaJn6BVEQKvUhC1xGe1fK0b1M9UqXfWn+sRx7CnGhLWzZCqVtTV/UMm
8poZwaIkjX5epy5HkjLWCOxUZ9MSZrQQzToqx3e2ao4asR39w7XDy/HgU0wO8bUgcMs/w7/Y87n7
9MkQiZmTFgx1khN0xY5EKcfNW4jSIKGcoJdJGE9MjKPFjoqZOqEDBgPIW1T8sZzVELI/jQYcHuHt
j4DFB0+im7tx+Gmd24UBMHWw8Bhgf0Xssk7bgab9/gm1YTPF37/qc9N1FeITo+9nJFwshAoiX4d5
qH5fxERkUDzsCQkCJrofhNbzoflfGbuirIgZL7tozhEu6X64o+h+qDs+fjoCvMWDF8YT/vpMxA3Q
ah438CJkbWaCw6JZnToRD1ndBA9lUoDXF22d76kvXJI0LQkPTE7vQV0harXJHRS6widztLECkgI2
MlvV2bb0OgSukFwENkHUTtbEbhfYbMB1egQ5HU+SFogHlrQFM1NHyv3UTeaw5exVJbXGPUpoA2nG
naDJ/PigbAw1G9CgDpSPkgFpVZvYhC0f+Qj9KrJk+F5LnZZ8B4sJb81pXGOVAGHx2GWTEwYwrMxD
JcBvoT5ki7hPSxvmOrjVxTnuJf5SHu4gw7lpPTb9Ujm953KkJK3H8HG05XHh1L3Ig42ofC94zOoe
FkrR8I3n8Ey65T6QmI0TjGs1Wllm1sc/tFg9AK1izgsCHGUOANExPjn5r1HdGxJ02nmlrX2mXhKN
NiFmu8MvcFK4SBJdZ24mfUqII5dBGMKP5NKnv1Nu5z0debXTQLUO/1S1KFzVQsvYWofTarn3mc1X
+LDBeUNG35yNI+FYrqtC2mAjy26dYlVCiUsn1B+y/KjVXmcjXXqnpND6Q3pGD6sh/OI9rauwdH3s
xglqqFKhoWhaB0/B91KxxdH8WN+9o9nj8U/mTA+KIjvSni1QsYg0c2HntzdfLKVBWbE1GFGOeKHd
npmSv1HHuZ5U8qa0uquAkZerkT0nq9TDDy4FNGBSM1BYjIg475i4Efs/aG4P159Jmm4Y2xFirJ0c
1boDUynsDmuLVslGZrrzR/+49PYgRu8sP4vN+KWaLz7lV/AyVHBpk9tj0oZe/yturHFLrPKCvMMV
tqPhS+bu72XqhOk0WUeCElXKB4rNcecrNCcyzmQZK7jOdH5N+BCx/+TkVEMPUk+ZSnuf7+79aS+u
nhrmFJEVBe/qtEv/unqxFeHCZvKwKsRgQRODvwscvavbNmoTEgFyUXKe8Smq8Csa/Ajtrd+v6Yno
6zE/swggiP/gW3AAMEn2OiWPfNgvJ4dHkQdzjj7HpsaqeSsh6mayOk5f46Iv76HajTtl0mvaBl4+
bu2RkT+6RInfUFMA6fSrorl8OF9h84fL3HG2ov1niNHFHy6QhcgRBrNOvdFtFJl1+t6+SCaD/1YF
WH/nsq/EsVNRWvv7RtEdGJXc6DALekoIqpLWL1Eb2Hp3iRI+RDMoSNOqcEq1IMsD/eLThrQObATh
ExIV4DRaLFX2Bjhks/52U59oft8d9p1Yia0iLmXg5ZTike63dcb9ph1cCt0jH1lEiiHQKucXXXsm
Xiey4uRiPpKVMTM5Bfpm60+ANCOsxIdAZXn2TqxMQOphfKu0CHlYEUHR00OND5JMGgH3HCEfBdmN
kVe1JxDqXnvDhR4wea+jafG8w49ihF3Sak4cBz4w2c+UI7L8/FryufxND/IYO2RuTq4vVnpH570m
7RZxODkHdqaV1ziKqYEItqQw0gtAHDv8+UXfbVzAXAEu0scxY83RswvYnfLQ5nkThQ/bYREcwsQf
36wWLqD+icY1znlkRGJpLYILmK0evIMAUZBfKOB0ksL5oYkWvxVOfi37gsS2sLWKGpqw7vmK/x9q
z/gIYYT90mgbHRzbwCeBsTceBk4QzjS3OA1gSAS4sYPupPK3T4spWUamO4fW3jj1Hgk9JdnNV+62
/148hkSNSiy2FAynLs1fNiDqf2ZCf29Htqr8t6yJwC9usHgyEBB4mFmkDozcicFygc4exwcYeXWd
5y6xFxg8uRKPIwmP9biesi2wkQ0CABnz030CMIOkPX8xEYEQqkgci0Bs87Rctkxm9roJFR3bvNN3
4ymNl9vqq6SnwDRBuckGM8yacdWgFNnQWqxcxo9qevVLjwIciI6nmYMdAzkraryQs7MKBg6KErNI
lIaYL7pLbhK/CJasaBgQYghXNnyJvgSazz0id6/SOT/6e4dG8t5/bbbMLMxeH9AirhGrEwZMQa3d
LElxmIzQ7LBUOwkDv1pDJrI9w8uINbYM0wK5gN/LhrCOrdvQYnjj3Z+Jn0uImZoti26gSVbTBNME
4ZhwRNI4B4btwYitHOB2I7/PVUMLjH9GRcBgL75cawkwqFt/XgkmsQbUA6QUsiJHty16POIePSp8
5YK5MIKunXpUbXzyP6b7eM9kfjTfdCwWRPwh5rv6uZqSBt3ZtNpXIUDiOIBcWuJK9+koYbuuXzDz
uf0rVoI3Xfc5+sDeQhZ24zSxEXKgqYs6dH5WcU9GSASVReclCjvo1XZtLsKAV9j5REXHk/4+VdHK
yXxJseGBVtsTklnI+rdui4YEaH7DprejQN++oWyKxlFHdLd2jqF430PDK1nuipGWat0wCejhGxa4
R2GS1GZG29lw8AoGrbzujBs22xCJ9eFV8/WkkkAjnURWk/zTo2ecDOrw8bSfJFXZQ+kGjza7EFb9
z/Sq0tpoRGQmjkEroZhJc+SBOijYvHMSf5bd/eZNPac9VmWRq8o0c/F36BQu97tXv1u+NQ6sBGqx
v7dcIbBmDtj9H5GjgTAJgfuyNgHJdghhSTTmYqQKWMVQ3E95kw1EBZt6De3ekUlE8RbgfQer1IoE
cQ+sQ7eyMeYEeSyg5O/d1yZ+ExmpB3u4uA0pXCB0rYvnicE511WvwuzLzw/lKDlaxkgVjPFYGFUj
pPYaZ3VMrCUT/PLq9+rVQxKgt+tFNyjqludqd2LGGHY+OSa8J3zFr09jCgpaFQi0JioVvSV4ZPCz
1GVlVX30m7PWRxufryjuQqlb6nDaQpwdDQ4NkanIi5tHYTafVA/VMDFln5j9MwTDnuq2H11Y9GO3
fohVt//vz4At/t3vW6O/T3iiM+0a3A3HEr/6krU0gy0a1QIdCC1KA+N7OXpdCObxxy8GB1BmtqLl
gvOHx1U/FDS3Wd+4hJoxL69SjQbVIoNTXblDwaQZasvmqymiAxtDm5HSXpCnoMvLT0DfTUhZXkak
u2GVSt+onL6p3benp8knFL8c8NenlWDL8A94HPop79lXV1jCZZ2Kcf1JId5+3Z7duvvGG9x71cxY
TPCvheKUoT7gjhYi1hgzj1fcmPkVAZ+lsjpRDiIXcsQJPeVsrW7JMNheQcGPVRnZZHeHVIn/XIfR
S+yHkFRroXKvCIyvxNXiqm9leyTbs1Qf2hsNioypnW37ftNcHYsXlDoEdzd55PfciA3ktJqAFnaO
7IhlwvR5BkT8RHr5eU+9/atfdqqARKaeHjt/LEhtIO/iMoQ14wzM+f/4uzpmhYtcAg1Zh8iysYqY
V70cOk4wGKVBo2QGFRQlWan77nvdGiVjbzrP0thZDX4vMoac9FaL+CJqjijyAqPdS7WUXjwjHoex
Wdvf/BbW+2CCLBija8fT1gibcfbuq0renikJ4OxMhsotMdMEXgjW9SyG7P3Sisc/DkfGDM1Xoxem
bIUJ7/+jIztfj4v/6o8oaiFpw7VrnkMaSIiBGUVznEeuG476Q5mqhM6k5ZrDJdfzuOqbRDVDhvDZ
iaOupRNdw0QcICul1asUSdg4fA0QxIO1uoaTT+egFN5Dku7KnVqrSIPX+QzHcaxfg8hVsANUVTc7
JditJtH8cD2bKLg2lsytY0N+1nLT3vpYf0SuHydPb+IG6doHSfYKfZrBr+/pw9HTFIdjnPkg/Mdo
ctdooPt2fAlbBAV4xnS1kWECM6CqHc8ncN7vmVFYWfBM2xVyFsag1FbCJD/v4OdGsNCioKXgtm62
Puc9+Ha00yuNkpiuaxTQNaQXGsoPSNTv+uwlgBqxU7QNQ8dfJg/1InCQ1jSZ2YqOdlk0juY/bENc
N9fbive5iPV1FQH6FtvQ1EN11E/iXcGBIv7+mdhPYGlMNtzgZTkShQv8yOB6UNza5SvP48uioOpS
GCzQGUKj8pfz2BQVocOGLjTD/OJyAYu9D70UPe3VfrtPbDr6BPXr0yEgfndDaf8/tECBpnJMu9CR
UlaUEaIrl0SpWhx8bQiLxLMuY67m1qW2jR//2mDDnBfNSm8U5YMsWEZZiAaU4+AAfHddmF5fk499
yVJXr7y/s20DpTVxrVJi4ICzS8tdra++1Mwug85QX1mtx/cVmXd6nrYnKtm2IJD/ahXAboaCC4nv
1eb1aaOMz+pVGwG5qxqJfpKvTmzF5oXdg/BQl/y4BkHUJG9DAXHhhdLCKgjp0LC14oaQainOhGcy
UZrThDOFmR9k5xrFtscF4DtkO+9kWcc5Gk/k1tjvf0a1n7X8PRjOa/OGToWvQwOTJwr3/we+xLpq
IKzzDugVxtNxYYYinFRQa+4xoDMHtspgF/2YgeoqRhTL4UYo5pxuqsXoHTRlSrQhU/TOzqjrdZ5J
ulsUMMilamFKd2m0f6W3q2/BFkyrpmP7I1JQ6yXVlhm8WuqPElntrnrGc7mqRwO/mhb/pVltrR2e
SoWQE87wi+grvFy/iYJzR54NsF0pTJtMn8ujhAQJkHOL4kdnq6e0mveSLZcBkSR9mwfUmevhG2gO
WoJJfIgWIZwCcgOhlu9wayXzZTNSqNlNft5ND3xkvFXGgRJXd0vHXCS4h7G9/RHmxLkENbpj3gL8
rbXPXchPLd2a/O1ZU9yoVhVsy8L8pNqvzZ1huSf7xjgpXoTRt4/23g+NkA1n4N064Hbyw4FbzDVd
O6Mi2Ex3awRNHQaGyk6JZFde94xNttWB/21OBcarWvwkSj6R7XUq8CJtepK3xS9sKSc88PBvP+Xa
81cb3rWVDkyvVxbwIDahyVWtXDdtzPrcOyrkszgv3400vRyEbuIo9e3gFFtH5U7l0aceLK2v5Hi/
+aMH69I1fQwQ1RxCcGWGypkLIVUMkKZgubT5LZUYsUXkS86k3SM4uQ+tMnxR4joiXq+1BmKAFBV1
EiyKDZnJAWI0sywwu7wBeH7AyZ8MG0MkiFdDmv5rtatAFAR0XMBoieQv4a4vEfQTYIHP7g0LRQk2
aVaWMiGAz7iO7y/URUMlAirxKPt8aBvGw2/GeM8CYJuM/fEOY6ihqvXMZH0RDIX3g/0uVaDASDWj
/MDfeWGuBakqASjOGC1AtU7CXWaraQZnMTW7GIpD60ZUzr04+asRShYdSpq8IeP1aufdiEUrnR7p
nx4RW9TBSiJv5wGNG3v9pIIqfmHO/uPWjNvbwetXlN6xOyHxlUdXp/CWeBLdR5nqww05GD93dQZ9
PIjDirXTlskhs35pSEpvsz7Q838vJqS+y0tuUOkOw0p1+zqeB39tMNTVxa89qz3x5F3uaQB1eY7J
NcKZ+V4W0qu3WsX9fgrbgLbMjTHnHuI5qS8OgGkwSKUp0T7U7r3k1/Ddi1/z6VNvyrlb7KHmccv+
1v9/M05IECFRUgZm3zdCJdJ3/VkOinTZAl6DAZrljnORqH67xoYoarILKPjjJ79qDCneTUFn5Tp9
FzgLJyk3rd/QjjzP7CXaz4b4EJrzu+aceFp2CgBe5Iebx+8WeAoYmEO86bLA/lMoyLenST1ExIHV
WucxZT/a3hh3sJN4vBXpwQ8i7mcFDAexRj2zX1zma8PaRh+cRCam9/PSZtS0MH+L8aGJA9S/jRjO
kjRksBUc/JKx5KudlwuvPaV4eAqjdbs64ZPuqhQNQoQPqyH8xQAgnJkQV4hTq2qwNHeLVtr1T5Cj
Bm7ARj0dUm3eVkxEdJ4okvmGeTgCf3XHOumgabOESBU8gug9XtyDbVxaWkgTAJsGJva9HGVCpBuT
+o3XQ71sUUFHTW1kdbs5fBtf1Nlo4QlForu0eom6v9sp3g0GviAl2SBbcP0WL9+BGn/NSDvUeOys
5qY2MJdfZBzcu5YZrswGiAHa/bnTdvsnRL0dxqXm3w6VvAfjkim165dohW/t5kvjX64kYjUsUN0z
Kd9tU4KP2RsbL1PIw6OA/VMBlc2e98Zj24UtsAGivtL5kj3orWEQ+CzoKRxtXQPRI5FhorlateZq
ml708AMSt+doLT4vGy7O+7k7/aAMxQaOsUNOYoJ8AGvGR0Bw8h7BQiA6nJ/xGaM9CYyFQ6X91G+W
vdTx9wPJXGnY+t/AiB9dToQFPyuSFpt53i3oBQ2z+LjdOdYkA4gTGfX54nVlIkVFhFVRHWUPCvP9
GhHqo1kI49kgU0VJpa9T1Jh421TsFcRmTTYfIpTnxpwkktkbzGFlxVML4dnFhCpyQ51meSuZOQ06
2q03VezmTIIXEupoBCpKjNS/ScnQ0+JWn7lxwwtA1cHYFbVyI3ua58JcRR0mIYDOjFZ0wG6tOjDt
7Fjr80F0uiDajRgWDfFwMXlO3OGv2UvuE6+seIs4/ZM1wHoher7ephBzstgwmO9dQJsRVwF9D/eq
UyP7BEtXT8chDitBhrsvYY53Ge459oSfaIm9Tp/WGpx/IuBaH/18fPhxO4jS8fXgsO8lgEYAnmNB
0i5qZRiqy493bR5IPXL/mYKmP+LxgMgDDv1IoeW+uOYqeSeBjKzS0EpIrSoWAmhTmRWxmS2XItPs
DnJPyT75YPGyH1HjrYHFozj8RVVE5MUgn0E9IeYDE/6MCQMAAdM/h2ER/a0tp3SfAxYna9xV59jt
NspEbBaoF625ZaXweaVcitiQighRrjTcDuNf5jhmhfx1KfYQQwpYuOM1me8kOjXFcT5mv4SWFqPs
Hh9yZr6b/6v5RQiIGK3ceyZLGiHYgT90zeB/6DY3LqzfIJKKQdOsAYkRFoIMMRjTnV84Wj3B74xI
8AWSV93v6mgYb/oW3TKjvB+9Vpxqqy8mXY/IJamK4dlWbT1tRlUf1POwmmuV8CGjjCzS6DkGvCbd
JQsY3jmwND8wcH+RVR/aivB4rSJfNYbh23XN1rGJYgF2tcKGFFfnsoV9SqJT/jNi5DO3OIU9FGyl
yjaA/acQA7wEwLm+zhTMkFl6y4HNuJQfWvHy0a7hSKcTCMaoUKk7+1Z+oWJLLL+MOMTaC01ae+qq
YsbvDzhnzYFLyzODifGJepqYJoE1hN+e2Utay0q5Ury2IWs6jji9TPU4ETUQ7uvRjwfd8vE6Tm3T
XRqSHG35qLEjCvVPhaDoAwmnBcaEAhQvbTmniEj5z/zH29hPH4UQB5T7WvSJXJBfoR5f8B6hxe4Z
vHhFHmV3LDou1bv1Oey2SBhx71W04V6B0jRMiRbg/fErp4r1yVPgvtz13ie12D7AJKoekUN/lJLL
0qCbiN9yQb6OhdXc6nOUMR+j2N0lZ0ObvjPZv0a1ayxV92Svsvlvj0qRHKwzjmArIEp2cfD2psOZ
NvDfFiolvL+2tWnN4PBZ3pWLtbDdGMcZt9euhsdCuURg1/t9m1dQQG+TkoaTj0g4lL3OOjwTRshb
2HQSe4Nf6Dy3n+zCDFM4FTyZgHkdmFAsuiEiRYP7ErSPvKVBnb3CXYDMZT1Gs7iAEQ9EHDClzSYQ
7q3SgaGIghZZO6STL6hAZME7cFomKBOwkReLQkNwCfYuZ84K7J1dccETt8lFaHWV2LvoVqGyPvgn
8Ta4J6PcWFlMgDhm89ikl6p5Lkn5ykpn5TD7+ePTj1+9eky127aUL1/S2vB4DJ81omqv6ZvwJest
TfGpSPrzL9RqDxi4/RHgKspq+ggXJ4S8dn3oiTWf0oCBnbv3AX97n/0Cix8IWO9C/F4uR+rljS0/
PGip6+Ng+lWLovVvt7cCUAC+YpqVvHGTa2tKHt7EtsWViy9c1DzQZ7Ff+umkOcd3ePyqXvKGZfmQ
6a+TZvKrb9sb6BNi+ARQs0s1l7BfkK9aoocVlgm5Xfae0hAzXxTnGEpAReIDEXb3YcQHoh63W0g6
Tbb4jB8pwpWBZLoobW7+8Bk2C5NL5U1+ku0YTXKGSFzg7K6Oxj7XlJTnvX0d7t50Vv4fEmnGEkyX
3Hx6AqOwwXLMZoy4caUhySHGEOMVobyTN4VJosFVAbriW0TQ5XtCUdcwSG/e95WHDeZle8C3nr8f
UJ1uLvnrsQaczDMbSMMSit1qkFaYm3lzaynEL2atfNhosPqQzRjxV+HpBwqVQcPZCFEs83GJ5e9n
i0VJ9+iSOBaALxHWzOCl5P8wC9HPFReT4hvm9PWTFLK+QvglR1Mf9TRqHB+5BcAabOsfKtDHbEg4
BvL5z5Fzu6wjIg7wt62eX1rlSBC80Nr5qswb2BFyc+qfC+DYuvXXO20zM/uuqvFLxGS8x4JUaxV0
bqywZG0qiBaJvcS/Pkzc3h/H+BhiHeE03J/emqhMTmM3SKM7CJ4l9AQEESI8DsuDOBGFO9+FyOb/
quZSivpx0VrJpuRaCOItSWRqX4M+7f8KEssBe0N4R1NoO0HCfP8W6iQs1PcxUvpkQ35xeSXr+0Wx
RE3H/M4+3C4DwanV8F81hrFewim4nOVIbnsX5Lu/hlMU+A67xLUNFKq+65FW4ChFnd63YBbGip0z
MU17AudAOoDoyRsS3jQMAioX1TW0V4TmvveYQGcQTd9gxFc1OXXm2QT1c3vpkTD8syOa3LLG57Ua
elNTD9aWpYJrIDxmYPEQUEEnKZIswK8nVc7IdHCtHpwmsRFD1PSE6HhsdwKi/aMuGQcv5v94xLfq
orv0JCs9Lwi3WpkGfBRCgs9HPwKFkXNPwk7a4uNMraBQhQVD3+eWSzrsF69RmZBz+h8t0i13CExA
bqQuCrbspaqEeZrekrzjSVQjxk0ZJls0rXd8d/wbvc1bKG9hAovx4+TiyDrYW7m/8zxUjDVXDs/F
YPL7JBGy8fjwEvU9AmL0D82usrm4aetmQILXKHzCBVUUjSlF1snHw+rUvhendvU/huL0S28CB9eL
q79AkFACPZE00IYsOwPtDW90S6MKWIxYPQ8JqdhWcYsch5MMtumwg8Fv/pRNIu5HJ0/efDTodd1J
dm1n5KMdMaMI3UjOhsJrgN1xT36Etm8rvlvjr5WkXyNFLlR40mg3aE1mUxo+ov0+sKzm06XNBF9R
ZbqeZ5FTvEc+Jdrtw1ZfiSdWCmZaoUUQqYlVHH5lofA79KqQ4nEVSNAHomDiOJgwlbtgPwjtKiU6
C0ckRvteIV6tqYrUM1nkFbbTL120rYwrLW82FsWP05ynaPLkMqF8EkSCf4Z00W6EgQAPsh8Z8JEs
BSo21rJnRnaFNTL/++yzrtHIrikTIZP5Oqe2/IS8cs2GoL7OZOOScnjwk35gCS279Dnp+BV2Jqn2
5zHzf8MKuGLU+fIoNov/XGSqzDD/IueM0s0lRgEwzLpMCz//EIvA0WW0g4cSs6VmTw+zGd7AvtF5
D1nJPmaUg8RW0h+lHzqpf/tpnKPi/PyM7wCcfGfzqjtdXC4kElJy3sRsUZHxzGCBKAmtZh8RZRYu
8JDJTg2uosZYQ34aSUj1Wgh/3Jra9MVtq2yUQ479/MU16mTCL2E+N6XdSGaMfJWYJMEuWj/ZS+I4
TYDBFawZloPC4+e6l4H7LDOJRuVgjh+VX1bH7GiKqYwE+85dTeYM6z+XwdlAs5fkX4XgUU8kE2Qr
1HdM2u2cDAg1adLcjNKKAFOk5OeOqj4YeazAbpp7yaW4QuXHDxM0tGlVG6CHL5q3z+a28iTXqyxQ
fMLidJvQ7O/41rytHJpitY437Mec+SXRRr4j3oO9wsaFBzybI4nU13TQPGbjg22kVJi9dZB3eGsl
DUk2EnUm/6o1XwPP5yYbFN7utAn2gXP2Z2qIelolMBDY/eW0RseEX2tnFsf+EbM/7yiwy6ZUJTbA
zZQAp18MYR879kve+gMv7M70hPCBTSEyFc30yuz7sBvfMLJji0bhUsp/DcCAkB/836WDegDowPn7
0onnCnAGW90bklhV37P58k/9Wsxfw0tQ6up+znoAF9OEaLKl13/qH2sVvlortKMgSG/Eo9bR3L2Y
7arLPKlvKDny/05uFMugEWcRDhnyO1n3JYXbO3VmbYgxkZYz3V8YMrpC1ka+1FncmjM/5OiEbnZK
D7E4jfON2bCjHbXOah5EtYaoUVfpjWsDiwW4XJ9JE5ERKOEY+VJ/Mrbx455MrsLO4zwJ1817EWgW
fTse4tp4nQWT4ByuIoWrxCWGzAV/0U7WJF64ChYGc8/iHHNRngWyWXwT16SY3WFPk3jAl6DwYVLE
PesQQyaZgriTNJMLwh8NGr5Htv0msq45nutzLoNzXIpBoV2+jzUA70UujTC/3CAsAOrkBpsw1dYR
cvq/1aFd0F9Prxs78x4z+cVAiqdlwmC4czeSIZyZ6OancrK+KRGT8gGoDKAiIBAF41SvMgnxckKv
4W9Lh3Jn6SbFi9w88pqoIZz2xc0t1HshZKmbb5SIcc8ojVuGJDpbE0Pk+3yS6KGARvnt62nmgZwr
zNUMWZLaVdaSoFlnU2q4nchtxwtc0C7t/Rlwq645wQUwhWJwudmH9m7oQfEpPTtrRi5eLCMPjOe2
pEHgqwAwnTc04g5tJuIK1DYlKD2l4r98lgLm5mknczwcFb5Zkze8DgjGgMe+rrXXHLYNbVELNEJl
yKRXJQBncavPjnV5Jk/kDakBGDsqebA1tBbIrVlRnL6p7hn414zR/y8vT3bfB2i0XSFZGeh88TvB
bKh7NuXT3Wt9iMW6sfeSR29anlqTnERvtAWaHYc06jq72aYEPp44ZAIBKO8EA/E+Q40NASRprD0E
3u5yAW92hisjKZShk406lBebGVSDrC4tpuSEzN4keHu3+ZsHo3chne1cdr0ksOjJJ/Ut97gdXb2y
t9UNy7ayM8kg/x75NkBUwk5vv2SKQEla/NfTmuG/DAfEX3hci9vwwDrnDiBkDWzCpKSOOV0t5MNl
AoJI8zds/iD3mhz4mQjs+S7oSJ36kwzKv9akAZWyJ2r5m1W9c2oIT+ppWjloxhW7h6jbtpZKvpmI
YCmo6zHdIwgKUHcVT23OLbB94EWz1XKp851bNR/aXDs03BFY3hkwdlUMlxo6cpjIBXDZo2yCbRsd
7WhlCwA54ZtO4Fj2KlgAoRMnj5TdahO0TvnDfecD7PoxmccfssJKiXqCsBQFT56cW3CQXrOJjL/t
KN35PagCj2//zd23SPzT89UXuwXwG7L3RD1nj83goGkwclzhHvcWvwhlvmH8mjDhkImnSNWCGD20
yywP9WG0ULRSfS0zpGdMmU9SChhdnTTYAoVDH+fqcZfQhDzOXZm28pWotZ0IOxRFK88xi0M0YbQO
qrPvnYrtqHorUgmzz/lqYB8WVkdxQfJLrad5YUaDUULKEjHz/c805B/oitALRDIy6M6oZctuGgRA
I4dzcPj1uK6aOchshOWpokT1/npVJMoWr66HCRQu1lQks8X1CTxO8QXW6plv1JVrC6a5R/Hf6Dyi
QVS6VpxbAxpeEYBZQ7ohxmOcUv8D1qmFg840QEt2YYRZF9OuiDErEmbVIMVFI9tdpCsGRgu2Prs6
s1w1zOP1VhcRCqB3UhHfLUGBBRtLOH5oltmWPhUgN2T58bXN6WqVcvQvIFWqjkCduHEPlLlXE20K
myxn8HpY0suNigdvO4mm0iLDXBewTsTj15QvwNCQRlH1av86Uhbw0JMu46TcnnLIJcen/JDSbT85
SavOCU8xQ47/F3g8RQIflpvwEU/m4E+k+o6sbzGS1Aw2m0hbdPcAbpptif5hEi8Z5943biN/+jv+
0qMwfxFQjXn1QduD8mJ0seOb979jqQeJFDveTfe5IJjzwA/2+QahcXqbkNF6JYeljdfVHlB8y1HA
7XDyEHrsyt3qrWFZReIbMNzmXsqbMNaMZyu6LdSfnBzRyDkSC2zNmirMj8Hz6+y3qjssR2ch29eS
/AdixogZtAg6gfEk9cYriS/DoL6eJfrQeiCG9as8xCsIruG887EFKV92ECrF82i8ZLOV3q0y3LE8
orWPy1WrppWFL/Yix59UL/ataimHfaUSrwyYzUnx1ss0MHwfOP/EFpMRPX601HLM+VsjL3c2iHE/
4suqBd7csCGXAGkpZwwYxV13CNXRUqTsTBkTlsOrGQ0KPsRl3nL/UjC0xGjjeZy2WKsQ50UEuLEK
mFNBfobWomrG5kfGf9kn8tppHkfRiSdSXsctwhhAFiET0YCZ28SVTSJ1Ri5wBLeyV55e5AXhnbRj
qYpuvbBZLwk3hasJlbcVueY+hhWy/6XEcTEnWGrd/7Vq/0Gsnb7Kgi6S2yTsWuzjLsCX81ok2hi/
xMruGG/iyiO+H6Z2wLy+6mkmq2FhxJZmtM0ifPyui1qZTcMkecvD1cj242AcBRlWQk0OLHo7r1/2
dqPw7pssEz3KdDMeIw+PhxvdzPn2Rc2i07abOvK6vRQ1E8zOuPi25LTy0oBBEUkENvmWNYTFywqX
z8jTfYlvSFjQz7DsyP8vlybkPh5rW+/gKFPagKi7iRHcS9eJhPFTqTMKlVmATy4AXsKsqmazKABr
XUqh+SOry/mfz5yz4IYuRDg+o1U/CqoyEGQbSreoORO7ZAXksZ6kZuH/wY7wFkcOA+QIV/MxXlYy
8aTcTQ+BnUyYYlJuY1J/8aOWzjPQAWMHiWbk/U6u6fDVubddXsYVzx1/JizfFqLV4W4+TWPnPnYY
ZR5MAttQ/mI+eizlkY760bDDuHfFhCFExh1R2mtQc4E2aEZxH84doUUWJ2xwKz3usGYZy2TjTr2f
apfAz5HFfz76bT/L1CFNXJKdbUck4BOcr3b7/V9TWIRJ3DzCoHmDcFlEgNymsY1BwqvYVn65q3b6
9OwiZXPDPPamgsDjIdxsKNNL90ERO8vw84ur5P8TMe2zMFvIj1AIPQyENXt+3ZdM6ElwVdfVpczR
zKapBHhBB6QR2O6fwWWlY8jqBIc5TLdQOR3JDu0/bIszJuQwhlY18Vb0SforHBLOVTKUoQTlltmX
hhNgOAqJci1LY7ndHnCKEl15FygWqLEapFeY43At+JJjZ3Jrlj/kMHDn2UruE5TWs8B/A0IVfvGX
Jlsq8QUaGRtaPybbOUUfKu6taLu5IybIXjXf+pMqLT6zzn0Sd2IlgKas5hChQbYYhzUOBOpiuHNa
jsWvz0PgDNabSxMq1h0Ue9TUsLPW4ATR3syAYTJed+Q/TNvTptTA/GvJufxw8wczpkGkuFd7EAFJ
20x9GMqn1QST94pfpZ7A/gJTGymOKSu3KKWbxP3xOMuvSsBS29QfVF+l0xhxq2WojWRc3fBhL9q9
ZwPTX210cg1uPRRRpqZQ6Wr2fdUVPrAc9i+HxwZduNRcPsKRTlXm0X0fCqLPRVj8LjGO8+5Nglcf
ghNts3s7AIo/NqUjkYFLKZCIuG0yOa7/hENyKIlhzk8APae6YpXoR9wCbnfLUA4T/eK4ndN5g9jA
LQ3/SWTIKznSnjVnnIX/x2mcPDE3MHnhS3EdTcoc++9r3lEUHXtuivlpBN64qYLSCNMNPWvVUEQc
a8hEnS7l0TabZfyEnktjqPMZCLpYFh0qY35NEdLNeK9405laOVSXoapBruCumVY8YF3mTgr0/klN
XnbUnR8qCAxeTTlYS2G89fVm4LlMMTzeeGgHMysVFnKv0scY5yWOK6+usp4f3Hem2kLuhNdS7HHI
hyAmLxUPpq3SNHEw43yYG5YSFuatclJhaiDUUw4pBhRqeq1IAu/R0+pnZo0uIFbVET/Mkg+dXMdU
Ft/wDG4au3Vipk9Bva8WzHHmhm6KKhoE0J2DLqjsXOezNq0Z/18r2TDaqWG6yehLgLmrTy+PYJ6y
BapgUbI6HHr/6wULmjIwI+sIKTIxSYIrKl8VuzFVbZccXleg1ev9c0OAUze9CMhZy0ZJCfpO3Smj
bV0LEI4l+YbrlhPJ3WI5/JFkVpoHkdV8H+vyycVU1KaSMgKF65AOlqOQ1g0/6P9VBRyF/ynH0grL
pt2+jw0pP3GuRTdDXn9Umn4jPg0HNdar2Za10aagnvL5yNpYxBV7KU55jLyBPnRdIh5H+0WNSfYS
4I99Ey7/YvBXztz8husziaWtZHuLfRbFKFag0PHRYgsAY2FLTWDg4mDwEa5klWFKoPTx+39BOg2X
ohOTqVPRINd4dTP1/YyOO0HiNQjL28nvRnSTG5s/GCae9indE1ZkDzKKJgetF27q+lkCU9pWImj2
gljpbFt12K/SbMZRuvs2SR4/qLPPSmmTJhKFvHAv03hGnfDOtfbkx7hNtYpP/Ffyd5SVjZSj/5fU
ForBj2fklylTcWHpX7cPrSKAn1OLRpw4Otq/WGoCIzZxa9gziOa9QM/Eb0ri3N4CYdVRj1+dW/vz
9PtT0NVHxaUYyLeJsDYPnj5amrRn6RQnx43e4Bp5U3e8JTRmIzbswOxtb/Ff0bP6D7ra+pwxot47
dc7hV8n+4QxRoTNuvTKmUVmQF+Yc9RyRGIiK3OYorUjIGFQDCzfkOLbBM+w0EpCDbahhJB01NUuy
JkrE+eBU4noBY5TMNL3IJ3T4wqzjQ/7zZL7Pb4vpYtjfkdItsy6LTUPq4Kjlg2J/whmpFdZGyU26
FwTb99VCJgoKErn8Fpi0tgUaMTIJE5peHPzuavQqbPScE6vsbH1XczeG4p5HjrEX9aSfjXrIUW9x
uUyAN2xw4jFU/hhFEe8absqArRiXSjsUqN7FTJzFh0i8mOgNYBIc46qXBcnJWDe1nVA8/FXZ81n9
VgDWYxno1JJHaNhECK0D2ijJ1hUp7Td/h8cLgh3rTDQzxdtqNFR9uekXDakBVyWFvvjjSnMNwubJ
yyca3MBqBErJVoOTDMLDD6L4YbfVt9KQX9ubj8eftmo8f5ERLTyiRmvo+Mv7qBeH420ZF56JWn3A
RpBXFiS7CK8emvlNr0UoJp6u1h2Xbb6u2yu+M3lw9ipi0ttdpftk23NLciT9FXpiLp+OmU3OyOvM
Dt8I6EUtmQcEahIoaZdRerPTcgHmrMm/erLLTyhuYSUJFw7XpFRaIUA23lHXC3C/Et0pDUhb2glg
TPhM4CaOQ5r155SKqj24Pgr9DdyW6M1Rm0AGlLeowdwLEuekRScAky5WwuKRDFeLbTis3OOSIZFp
F5P4uxZweraCr8Va8ksC7OUAL4Zlb1nVaFHNAAvm42jiSxVYjdnix7Vqvz3ccTPwYeHZm9X2pabk
QXYw/S1ydn/girrruEaorQ33tpijcpBdcOT+cLu6RGHxdVI3hLNRNQKYY/DllCl2yi6+poTIf7DN
AoUtqey5Zo2/d6t5PtYsWg2hgMN70SsZub/iLoNHyJBs2BuMNBPHwrSk98isRVhxB0ZaujJ9AD3w
qQXxJABTISuPFmJLagt9lxbsePNFJTSpMbSrg03k9FBWKKWdnVYdEYYvUgTTg/Krl38ENgHFHpJ0
RUEocNwO7y1nBKvBzp4Uu7/+gSBN2BBP3CrnyH3rvvG3YfA2ZYxfUX6WauocU6nqYf4uIh7roWtM
IkN4QJnimSgpKhT/IJzHY4i3nJJ9g1y1djDzKhHozkNGL57foxIFY7Dd93lW5p2sQV1wqBC9Kz8U
FzK9DZ3j+hC3S2vfxz9nNza63YMv/M2KDmW2RFZj3Rr4HiHig25mQVWFSB6ewgDQWKPnMQhs6Ryu
P/rPHnRsUdoKc+5GtqzK9PuPx+8p1U//zuf3vq4Ujg4zWbRoqXeMAr6V1vAPn7KPKqyv7Il8usgH
4YeMx/x1UplaRn+oSeqOKPLIR9A+KBxwoyvHk7n1x6LoLEETr+TuT60aNAyGfZibZU6Dpfu6d2xQ
adLaqDk9cezlsT8W3bEkpz3FY/eaPqOoe0zFc1Inzt+2zh+Nt7Zj1uyph1cypL3eR7ZvBwui7lZm
mGwjuU5exi8pHH5P4+8R8LIlG4C0c9wAvYIuM7XPJmwR34qyzZAivlOgFBmxXk4744b2EJxTNyGc
6DQC+8fzXttvXFxM86sA0wtLPZDvcl3OR1KBV7ZTij+2oZetQ05L/crAKDEmKuQGxCpK1t2I5rhl
JZr1iL4DYfgYFJUYNcnWm37z9HllpFF9AqYECmwdpUiQJIVPfkEsflnkifA9ZKkJUt7r3Jv2hASO
HcCoXbptzXRpewjnUivznld0EodOyPBte+a+7UpNYQH4fA7YASPRnY819R6njTzeC3uvdpGpwLDW
HcR2K4232lfo2e/Ut31i+jly6CWt5nplcX49cdW2Ln+kiSKQf/sXs7Vx9W8JWKN3Rn+k4/c4gxhE
dbCjFiIJNV0UGjdxofN0Xbb2i6lnWUnZMbOUygZrWToWTfIVeAflz9YbEjTLRtLC3u743VrwNYtu
TMlt0GfrCiO0Ix3TF20gAGuBSUmpxLCA8s/I65J4Ujdk36wcAGHmEzBqNgKt9iP0vTnspkRP4JlL
SxXPToF83JItHPnFdmafkVmxlt/ByEytoqXehAqrCyuPrWgNdwTmwJs5LFagdMFbZKEtnPqxQeEo
yRPAGpDIO66GKCnD50MvZvor0e5Pr/9C+Vt9ugsm6ondTed0JOaSvj63JDHHhozo9vdd6n6DuE8v
0QiJoKV0pB9A9Jw5lmV83cmd8kPmSC59FT98wSTkI7WbEdPw8pjOoI5e0SOGuqMwzNhfWqqTO5wo
EpPwkJsZbjhWVO/KUJxhdlnmYpO9KGX5sUVsSylpfvCVBNhA6hk6XPhDri0kRSpqE5TrooAROCxZ
hfjig3/NtgM+wHw7eSF6mpiUvOImh0ZQYrOStMs68YgkgzyK8b/R1fKPOKOuKJrWbNWqHzRyxyrB
GB317PsyK+rq2V65BfK6ExecVsg16QyVL8PNv9eNzNoqz3tm8CYyHjxQI4Y7lqwH7jAEOhQTzy93
Yk0C8AItaV8gLo408mRVku/2MpsslVQcIm/Xq33kmE1RgSbmKiv2ZdDICWa8AHAvBpOaVvDWu8/k
izSc3mB8C4GCwqK58zh8V5NL0I5X67HS5IowRK9mSxT5VSmv88W8D4yP6LGxxcBnarU6aWzJEmnR
71YsfdTEQc+lUaUQ0pV/jNLVDvfmqPcryvY6/kMZ4EPGZWaAGUrfHKRqK0+HXcQKaDFehTYtZGBZ
aRU77/6gdil0k1o08WBgs7GPJKaAcMbcnhPGh/SVPPHmBK4h0X7rIO/26UQtoYBUA28dysURVNjQ
eqSkhZPBvH9MS0l+5+BdF8OVHrW7zkCO7AjpAMQpPIuBdbDFl+lsGm2W4Pn067USwi2h0/4YycJq
fvANTRMEV4eNTiIYekkQvL34HELcDVv00i/hWnlknN7LzL+GGOBh8vOTKUgzsJ6zTMAD4zTW4+nh
6P3WPRRtJIUw23xO9YTZnROsilvO31gMA6x1/jRdvTvIuKGRMmjHc85jErR0R7WP1IY8zXrmpPuX
HzDN0MDeal2ODGgx40Fm3MZprDP2WCW48nKwLjjiEOp6KdEaYv2IQxljMYrLVdPz480kA5JLJdqb
Vy16nL05LMoybWalJTgwvNPlOnL5vwy9hRhjIBBCMj0ikzanXMZ8zexiJcsxvx+g8jZdVdYVpmF7
upKZf4Rg3EggRG/WRxVgeLlfq7lGB0uY33PEPn95FoqWumoJN7j2WQq2B+JzOkUs1QBebrCAeA38
xa9VcNOaLyTTWYUctAl328avQaZB+ewMFOkcKwwTqA/g7qknt+u8odciQcE6TPIqy9Mmld1qtRsu
gf3SjJSiTYoo104iNiyk390QO7AvTZY7dm+fpemntLW9Ip2wEr3B+ALiwTjXH0LjheO1I1k+zpMB
E0Lz5L4XQDN3jNHL5cI1cSaMASeUxJPc0i9htQ6BX/mLLQvdPsaAIQnLcNfdqRMbhRVSbcTwOBM1
kIHZSKEQUkdScMGQOtXjQ8yccSglGIRFuLHo+iYSl0mZVxVYCFOIrUWw/CtSsU1+ksKuh45J1vMR
mhqQTSMBbK4AOrMKE86u7h+v7xjT18XcN1v/+8tQgYqMFp13CHFm+TazNFJeKmQO0Fk9PVGQpNsP
vEniK3iCmbk/ZZ7Ev0tNyrs7zhkICZ7liGLCS8GKvrcE6bQpwa7gWjOXLOwV8as0fHOkPHwllTD0
TIHOVwNhkpMDvEfYmOTunZsfkh4UXF2AR7eTsyQUpItdqlmBUlg+fWfqy+6HK76wEXCd30PUu+eP
JpvNAyvL4WrOSAIQMzXM/fhe2xzQeHoOn9m7xorAGGSoQZzFhWf/lP9E7kiDpC90yTrV2r8GBVXD
pMvYEpRh8sxmMW7NOFLTJxXMEM4JDEZgrmIhpk5r9whJhpOfDDo+sMy2AfZRdywS5ZprLca4jh+w
4f9g8DGaQale2WBmfuIZ2VV8BCViZeX1Hw+x3rBOB5UG+sdhiecEQIpYJ0ftOeK3f/W4xL9of17K
eR1IZcz88Wt5cadK0AaaF5FjB8YDVkUYKKgRlQiMRRi7daI3gY/Ub2ysoOJe0RgJjFYW7X30PWJM
6W7zeAfoUxehyxwCupc+dOlfM0SRE6KgL1j1+5WFRF2SCDzmNUMm1rd+a7ElKShf40l/2jEq3Uh5
3LxAzWwFLCmfQn3494sDiVtX8Ex0Mv4F5GQT2vqy1r7DKuBXHdVVh95AP9lUTih4hIhB0HiXA+uF
Gh5iGtLOr8RTb09UEp+AmIIkmb87rqvBchStYIB2Acg0NXdfvYeveuRWs+BIYzXth2evC73aJY5y
x9Z56H805c3LMpvojCo6czXAPPFklIVVsnWTV7uHYzm99GsdKoE4BbcAOXdXJT9emA8SzwKTGa1j
uYXxwPEn3FenuwaRJ0RvM+t3b/dgxKAr9AO71gOy0HRX5jA3ZhlDpoUxACUVEC84Q9aURTLYWLot
4l/gWr6fseAgFqsCbWVNLPqjC2rG5XI0XD/lHFxg3kOittIY/9qAKfCawQhd/X7kHvyOM77Lx02V
dNe4FLgj380tfaJYr6XluIchic42VB8shBKyps4vnj+7TF2cit3yRugos7HUETraqQveEfkRdtot
NK5hI5NsMMM3ptoF37qLR+8zPiMNRfbCB2WvC/xkwWCt8eE4QdbcRbD7P+hHWNp72hCPsKaA8Wd7
/VB5l/IaaCUdZMUUDJnXw+wFB42vQs18FPLzILA6cRqHuhzwB2DxkTyvlUMfACycXPxOSb95y+X5
7LdfM3gzrAil8A3e80jD3jNifTIv/n3orr31nXl4fcRtXjDpf2vnO+HIfRzYu/fRICL4MN9eNRkN
hfRz5g69jE7QHOGe2gU3ZYwf2j9yQrUfQ2C0aPE9dwrj8RzEs8VXHvPwhJKqnF5zn5Vqz9ko+bOh
YvCK+zYMCWuZB1FBkGp9wJUKjDUnL9y5R7zCvikRykcCgG6WP8nlhIYj6v5TqNdJRf916AmToFXv
BdOym1W5KTchESQSKJ9pDiS7amNQQJjs04nYDbMXkecchVYyP5izgJloGOAZl2CWqAsubKFbH/2A
Up+EzLDPeaSYK9dxIbLpPUkLWPVlsffX8Uh1YB2RVbRLpxPrtXf+GsJoOuSHdMteQTyjtVtTJ4ig
RtPXTpggoLTsETU7idVIKr7m4vx7p6fXKUGxUFBc/8S8Ttvh1Q55AUgz/NSlrShnE9EwIgy6G+xY
BnnYssh8cXgBrCk5ohXhkBGKA02UKGGtIXwleC/5FwQc639/US97PT/q4WoBp7x6gTIbwi3ZlWfd
to/swXGdTbHah8/yWRRfPXASykdAKcncs5FLP6Ztojj2koCt4TaW3GAlnT7G4zx1E6l9R33kE9Jr
wgSQB/aVuLZkZWzpR6FKpPraE81mv8XDep/lQ20JYmM1EaS8ndQx5Rs2thEB74kPCvM85K7U/ZJk
uWG+B88tAnZTUGu79XqO58GKGX5jQItBwlJNEbnGzPVSRf9LbiaHmhzmrxwNUbfG+0Iauk+IpHbJ
8oOzJ51YWHe/4TK2IDbO3j4K3uJ39mtAgGxCFEOLsQ7BL7ZGhs5CHEWhChajVL0RgTdEjPrDwTRn
itNOA3j83H7AdMU+05rUlNhzNYeebHvHl3r7F27tUoSTNvHYQ3mOGmTIFVcQP/9QQPYiZwQYx4lJ
Wb8EUNFb6MlesLw0OKB+TWd6fud0m40OX3zia2lBc3WNUGQCw7NZO+0lPeWgyUkHSN5S4KKW10zf
8k2Kxrn1/4bvsaMEnQrRvBTq8b8HwVfRT20py+Bmoq0hzRrurVDlaRTEo80gPA6R1GrqbaUXDRUh
TgYTyUURlkliAVUtij/PO+2evsGLdCk31YZI2e4ucZTYrUXD5GV3YLNSqCiJ6Oxh+6AhQYu66nj5
NT8v+VDEWNHbjQLgHHPx7sdr3xK/2fpVNzj8ZGWwWmN/9xbHAnp3OQkudXOql2W/4mXsrGqn6RzI
gg+59yX4XT7JxNQRBRjfxR5QR8h1dP8l6j7/u6ava/OHDH0hOvY6U9PaNuN7ggVlbXwdKHiF9bT8
+14cRXfBxSOF7uv4fYFnYAMNJ/UMM7AD1BMEoFMNm9+By4bhUTqNpdJSdzAPufkFIRC9dqMtiD7y
ysQfaLi541+DiaDELCCl5wJjUWqz3dHGUGZkEp4xOLnjPpsLkbyXekqxDa7E/zBc8jnT7MnEwZPK
vkv4ujz2FpZj6JQdax5iEWZ4WguhjNEphHBvLvmd9nX3KhkuZBqz52paOucK5kbdpYUhtMLX8JD/
dtG+G1izdqUeUQP6N9xHYhwNrHJ6zfL7D2T4rW7OpynLUmimo0LJTl2qOQHzPLMug3VVQ0HbmGz+
HaVw6TpHu1gimpWiDfb4zIPaQ9Xv/ngXyCn6CmD3jD6DgUUy5qPU320Bw3om94cPsnpfpV0OgsCB
9ojRJWmKLT9e5MNYHwSx3J7Geux2X2P+hWrLOTEJCB+M++E70BLZhBhqT3tlZ6GiV6G9Iy9hQqQL
vyrTEmnyozdUDMVP3xah7XJiQin8avPaKSMsO5cl9/fiDeemZMJLYcUAn2o4mA4ipKC1bNJ6OObx
1ztkYa/s9xVFWHh3dSM+zeqZDF29LHI74AqLy7QonEnNwKSrQ26pqb0ZiZEHdcPxPllRrDgNl46f
pMoSmXVBV4JDQXeDaGuGbHL9HWnJesWtabX1/TTTrIFYqU+xXuSdDid3CD0oiaywmb2sVye3nXVU
dhIgwhb7Kj+hzf5Hvaj3v846xA7/vyqasX/yxEHdB4IMxuZBOYvKkpxQ4gyCIy0zPOefBlXLXt2w
HcvF9nIy19Frd18o3skghEWBwvy66fwpt7gjFPiDOiqgpUyYkkibk9zIcy0TJxMw8B3VCKH21oQD
nbVICaed7yeaFItM27TvAI6IzEAkN7JBnAzfAP9P0KfSPl5OIKIMFYIu7nRNAGxq9hX1Mcq7xM9R
R23C5/BTOI9UuMQAfQ3aengkXxJdf6mXmD2ZzeqlthKku4Idb1epYBfiDRLw1HO+sn3u4GHmWrPM
wI9GQ3wWZudY7+ffd8jxrh/N6EpdD12NDgU7JoRnGAVrKEgXAkAhLbes2hQ2pA/JxD+zIB2Hv7p7
RYhv+56vDufAPgIsQ51ziDMRNYyv1zfAa7WWi3KpfEDoe0ROBPnx81AHXw+/PQoECU9c/YL3r7Sh
BtqgFlXc138xwNdwnrgDIvKEkbVBmDZJHleCDDux+pGMVWczM1jwk1YbSXwxYjsZyI5X0+yE2TQ6
fDGmRIRk30zwxjtROFqWbBC1Tf/XBd09VFAiFk6ZZgy2ag/H6l3sphzmf5pLho9aR27M11ftWe3o
lg0wVHb5IFH2ZzomXeDbkCWBy8MqR03RdzxFWzXTdy8bzOp/AOMtKq8XQfWp9CNk1J9DFVvMLo/0
QEzscTEziogdlfFx1aYalFAFXUQrPxSiZZBcZWdba372KYf8jzuxAdN17BmVjdjz9sWVXsCcUvxQ
oKYbZ7dT7t+lhAkGd38jNUhLnF2bEqXSTpUj8ODnhFYqQiFoDdlUix223zS/zRLdXr4r1xYdC7pl
U4VpCWoG+amT/fdilm85Q8n2VP57AX+X5UtTA4WvCAaWtKr5YyWIX3oDBAR/9F0euQhBUIMIQ3GO
cPRClpX61IqQD7ge31toqg6v3V18yDUGcsFukeEp1mhLsniq9aOPwDGW3DlEBaxjoJ17R8FCi0Ea
8Pv6MqWigmm3PTTlMFJF07rvuiqzA3cwnp90vyQku+53I7vlerojnJucAOQJ7wuSS/cNtkTEUBQU
oyKaM5ZLgepidVoF957gNHyhviC+NqtgRBJpDdvS5c7ckhTrNgflhr8nDiq/3q0Eoswe7y/02F5g
tmbql0Cd1wfub0YmiDEwATXf3a1WfCcbJECA7NeauS9ATOfxDkaa9b9/x0c3c9XVjMyssVC3NpRF
1IDnYCj1K4jvZFF/mHOjwQ9dJXglr43p6wddPGk1ENE1+Mc8J+U+lu/4i5355EA4c2UJdreQAhK5
RFnyu7rskEePvT0E/hRfFjx7gkT4DyjW2bjHk4L6bGZM2T4uqk69G72cvGSurXJVe3vpBPvR0dDW
rg9E1XKe/NPC8Knuh4OwUUH5AnQdjmnfa58zeXWTHjL8R5GDUaApBtiH8GtrfbZUjSjlcOxpc9Ms
MYBOwvNGkPyyc7WevImVSuJBsRf6EdRR10dyOT36iywD16nI/MRgXn9NmM6xfack6T9isiOEuxDl
rnVfn/Y0PKOhuSB/QWAde7zB5qh5I8pa+HZdlxe8nahC9b7avtgqMp6xjwZyvxAqMX2v7axIHR+O
Aau6m5w+4fIwXlAuCa8FfYRjxgaJcpLzIkPYq7YntK69TaaO8tmJnmIzp5EVD54lK931jD6iKwM/
RoHq/ew+8VWYMzIyah35RGgPBzp65iEgjmZ8MyAU1MTrlmStJz7LJiaLp49l3wX2Gth7PosQKwtw
PzIwkC2WYJt2Gt7OAzKqw4Wpw4CfMsY3EgUuSbE5zDTUvwNPaUoihGUgJg9zOF7Mu4x7iE/pmRKG
IAnARd4k47PetYD9YTq4/ISIYhE1ZVdjQXAh8tBVw+cwrps/v15DeAeT4huLeRQIHGhke5LwLurb
i5k1PYcQGrYFd9jQ3d4crcbyzaiWK1N2NZangl5GTD7top/Jzrj2ry8hDy2dsUPTYW7rVdiYmq7C
W58bFMGGbHCXYwI4S4+KK5dnjfyneCrgSNqcQfOYlXDJ4Zi1nuKodCUJ6QS4ln8tNxmnqMEOG/O7
uGiDi8okthzJ/l/dVHIQ1nAP3vxiG9swNCL+TFK8fl8gnjlcCrzzF7yQaFCyQ8Ex5pWugfWO2EHc
D7aHVrsNf9DfYZChM9Q92jfXsUkhDobORPYwVhTComL8uUQpPZ10XRZDibYP3ZV1PAVescVfov7d
gO7YJnEccnay8spmLP81I297onBSP/+ql/S7r5Drou02q9CjZ58N0Teku+FiwWJMA9FFGvkiVznb
9h5eJ7gT6+484GnvF5AC0VLHacg9zHwg7HRKK7C3511aI5UTSg0YhPV1TW5+gnMKWekemF9elbc8
lYfwGNrb+F+BbqGVdlR/X6Fn0ksfka01qV6BGLmGH82Kx6PgGi1IlO4xkAwHyXL5cTeIzOdrRegV
TfMTvIdyo4IO7bAmpmWcXCQZI2w5Ul+NLRPGyLMvsxNP8FjJ52kKomC9RepUp2KMSrLad0M1BP9K
6zrPo2PxMApoawA5qmNesTtgrb1WOSc9QQs/57X9hOLhvSkREo0tlnXcx2DseTf2NmEn3Wb3nvgH
nSGZhRYDAS6+9hpao4TlKqddK9aWo4uV9mP/xS2RodIEmUyaSUledVVFDQaALEuQTGlrKJiEf4wv
we2YkIQ9qMM8SNINWNrklzSVBZNM7lDhmxpNRQV6SduTETSjLfsb4JmmCm380EfQ36O7jt3wy/Mf
9DcwqW46Rrg88VXTa2HwRShtTPkoUUwu1HH9QA55QXb4sJOQXCrtDAgriPKpWtnl29sSY5iTuAqj
XIdEEcv5FG5+RcAfWa7udmPv1neQEP5EYVKu7OYcOFVf2m9/cGIJXQea45lzubGSMvwBBKlyIs02
4esNlqSSNv97iQ2TbTEmhDo1SZVkbtnk59otkcsfrJq5Whj3N4hkB1mQ4CfdIpKCxhKQmJKuFn7T
wGE0w43roQ1+vIX48k/lk/XakAjeS6IxljEwKDslkGFH2TkWzRj01+IYQyo0qfel4mlq78GfUjD/
6i8hFy8lniiTyiyemit8usaTyutgzPB+btQqdCItXr7As9w929ilYUbPGYvOr831OVJ/GKIChlmN
hMB7d8al2bdZIqzdzQRr1V8zLJBuesFvM3dA0pgsSrp6lPuqV0UXmJN/cRzbgihgMGLn+oxswN15
1djuyg6XBvCaSVn8aNorpbTagVU85tFSDTLouVsZ6AXAMB5gyFms1GMZ+O3Y8j41jAxRh8ynwMSw
PH5kf8U3/cjSNgsuMndBFtSYNCHqBEo1KqCebkWsqeWgEHJ0Yx5MObquylvTD7AViTOClDgcTHDy
5nhxKAWuUng+ZOvAUquWBPJx9cr92YF1qVewjBQa/RnjV05I1vQFtpSR1c6rlr4/im890vC47aVj
UMU++SZNuY0rFt8KnJ/xqfUB4vNvapPx1wfthtmetqkI/+y/93FWtIjrcM2Gtg07+JpSneVB0Edw
dxTj7kpQjcRsQkl9c3a3paTufH9z7aiaeagL7KJ7jPnJ1Ggtuzrx49ZXC4NRP/jScSKAcuF28tUU
FFhEhZPFWxuuG9MU+oN4Xw6DuAFXWS9ogeSWpXDzCD8X3Xdy3OmG8Ep+mknK9B3OOUbWcLyNej4A
i1O4SBrW0N6vWw3UDVfLnsIUsDJA1caYxELIj+pm2tDwuradh9HS+bHkIfBYkQ088ODLoEptkX+N
D+VQRmoRDaVsRXElzsxzBU5E7ebKisjZib9zjc6c9tyMga+JPFUbCTXIvHv7HIPTd9UvCeygLfuj
mZpZpYhbshgq4keREKr+jN+IXkG4n2g+4mx94uz+EAraOu5QMB5OsZbWHnLM16LY0aqLsFL11H7k
Tng5vgfWOxmiZ0/Vt8sPfCKzvvIWt5mhId8EGQqop5vmvoIRPaz2ukR+cQx8zR7LF/U1ub0+Xziw
yR3eL6eqZCMs5YMovbhadOlBqTv8r8cozbhJzkWUDB4Is9l8d7uzUl/0zJVQaW1+HlV9cMIvwd1J
/i3HutUKHTtsJnsYkmccv6WRux8CdVcHX7EKRYkBlob1T8j9pgRyZLBBOyQydPDEy7Jwb/IzHWJR
qUBJm80r5zbKrN5FTx3nlgk4Qq+SBQqSdKDtLhCswv19AoHkAfp3AXZKA/yt8fWo1dFc9d8zNNrS
OmquASDtNXuGaX/w823e2zXW2B474LFytnljEDbC9KACkQSIGHbdxvTsClcPZOqC3+QVgPRk+ldz
MIyj/F7pUwFbqZFlQ0R+bX6BD8/zlSHYVVWYODMhZAFvhZTdA3ptvbGx5V4piK9kloJSfkV+GYZr
O+LHvytXFjTugjy9hAp5y1vzsqfCo/7lvdbf56uwzVnPYoKLzabhsd/4tXp7nzMs4jPyZpP43zNX
fpvSMrUy/rh0VxN9IsouYta8/FqOBgj8vqYKy56FGe2r1y1mDjeA0m8h9oZXrXWWcSjo0qolP9lr
5iXj8piBry6tOGKqcjNeUJnLREa7BkcVPAQyPoIBn2R97tCQ2ENWrF3dobOXFfEYOVGTqe5GKjh4
UvdiqX+USHMUyqT05pC17SguuY7gIY04JPvJ0+KlP3w164YB+L2Sr8Qxgm8jRpeHI8LL430/1CbF
K/NQBVc88tUTglEKDAcbBUNc/Ra5uy+ogJDkGxS1DStdfIW/WBwT/PgoWavdnOajcIE2T3dJYTIC
qZ6Wv1z4Ely4bpgEGBz1kMTr9CzPsdvMrvCICN3SId2gvjQz2Q73YLf2+OVSPFC3BRbuAmpjiWJp
xZohGALM2G1IqUIjot4zZHUV0Gi/RVOkbs0S4r9kVvlRRAJSCA1GsfNR7sj2Emw3KqKvK3GgEO2H
x1d5WJCqO42W1FU6FmUG7sNe0vyIr6Srb79zesqKIFI4lGPi9dd+wYQ4tYd7jJVwHOoILf/fMXHr
olEqKXCNTOx9bVbAivFn9rXSvBYocAZvui/EFslFnxMsZzwxt4u1UGzK0QAvBgZjtqvOTc3ZzdmI
MNpMiYVsA4Swn9JejGhPBac1yZJz7X8qWLAgm+5fSRD4KGGfHKuqy/wx2k4gwUjVpLuNAiyVLiaL
DV4rOtjiOl/eczm8iS4AKYmjxEHcFCIRAb+5932IfX+3QGKEXYqxcEJ9KUvs/F30DEX9PClSL7ky
b1H065Fuh/JvNY5fNh9qHGt7vDCKS9TnLVl59Y98NdPHoSfebsj+7yH96jzim3b+dgQiwpAhvz3Z
F7papYhF13e0mkzmfdxDRGUZQrQzhluwlf0F+rwn9Iez+r/UEsgReIAWRGzNXp9aIHqUDoUlewiW
krL1gqSuTkeMgPQ9CdYdidQCfi3gxbair0NUbxcUMOeo5Jx1wgXF2H9rm/B8W+bdiXc5ax3Qo8yc
vdePYL6zu3Usq91N7uDt8aWxpnSwu6WICnK5QJP5vcRtwMP6pZYzfKWnMWgzsYNeGXfl4Wr+ukQR
nw/lECT3ytjWkAaY/nweIkdZlBbJnS9+gmShSs7ahfn8yr6jTt87uPn14R7PVKe3pMW5zBnhZeMI
Dqwm03Uotjga1bh19axoSD9eHIK7VOIYNpkyFmHUoLRplH/pFZbbg+w7xG6qSmDczl+MpjH9H6bh
3fXJU5wDElgfuoO8tdW4wZ0F/SXH3UhO0ZOGydoX1YcYGzf+atXNyEWcADhglyCNOhZFLYQekgc/
BJ3z73S2pfi6547CbjPZQQXa8BjF6UecwDNtljdcY855elUXxzjKB/qSsN5M5JsUHuNACvi2HwQc
FCP1PN18Ee0YP2N/qfoHck5bxEw+h1vhwNhpz33uKKlatuddQZsAGg3qNHX7eWJBnaq4wu34ckSl
0i8PJaFclKbWjrsdykOt+HLE9heSOcdicMDv0ti/Yhn+OJMc/fchYhVX3bTB5MEdZ+D7iwuTb5Vw
skIfZfqU4/ft980TGvzxfRT+Jtmbu0e7rLT3AghNjcZQWWwKO7ivK03tsazok35lgEGr/8BmwLaQ
CPZ6Cv6Ekbumf6Yt9lyY7rpIozyHpFBC+Squ5COZNCEzC7YdRNmG3n2np8I50/vSh0pJYAsNFXRh
a1TQOo8R2pB1xxLrcQkXtPuZrVjTCIT/KYMQzqkqRj/YUu/9Yn7mM0kvL+lMO0b0Q7Y4xJ1xNyDn
SSrrDXb4mu2f30Q2xiP3lTqDsTIh/FLSsVwo3x8KV80WX7xswanF5soPfh2lDroej6hn+2CjW4XM
Vf1kX7vpdwruEuZYgFL4NT+KnRICBpe4MMtLl+9vliqpSPL85k2u9yOYXyY+mmwSJNpbah2+jrDJ
2DfaJsV0QjFo54wfZ2MkpWE4XO80yvU9sNI0Ci4nW/dPY7dcBwrGMpJLpjSfhL9dM8n2pSSxpDXj
+a40aDg/fDZ9xutvjzj5UUDWy6s7WpxuZ3qbPQZSA5CTynftAUvBOB3CD5pd623ugDM1UwrH2kLG
lhMXwnP0y43Xv/TVQ/tZWcppDy8kE4Gi9b+T+wm8efuG2PDvkDCGu6JaBnInKJjrrJyOxgNw9EaQ
HYK3etwlw6mmWMrQh0wgF+/8XPDiqMouRTOtvbcGvkxPg5aa4bX03dcxofcgw68l30b/J6rNKg14
P+aipvWsj56eBAmvqKpCTxpJ71K0zY8YHGIV7LiR3euqqW/L9D/7ME4cNwJhgF3sakha3YcXwZWV
vdLR4mv8Fa/02izOxdbbQebhFWGTHC0MLJXIxmyAXA+ckqrt/+9fIpVBVZZBpuGiz73LAafTHslk
u5uLGJyUQYZmoHA3YEivv4vGqXesQL6HzVcU6rXbB41xEwGw7tUWgcBY13uQl223XshQLM6s4rBj
DrhTonUE/oVSehKSgyhZKfG/G8NFz+bSnF8GpBjkl+fCdSmyZVxJLX7AUzPikL29+Y42S+uCEate
QTDIdbU9elqAdbvLWUuO83/kP6mYXMa771BSOIZ73XnBTjuxTyfziUWRah1/EV9hAglmQXWY9Q02
ctWBwG842Xsyzo7cH5J+9toZgq26KcKEV/v6pIweWofnuly/SEGMvqGK3sZbCWl3qRx3JghZjXqz
rAiXvM8POFwSQ37YJ+5gU8VMgnhKlsB7SLBd06iQq5+M3WBozI5zh+im0IlQQdl3FUq7w4g6Z9YM
KV7hlSdZ0NxFIOPP4YloDe8zfkzwVQbBhxUxL9uNeX9xgOueYBQF3bXKTfYync2KF9Md3h62zHzM
Rsf0UyeWesaOl5wfv7dA7RCtHipyoUcQuArY45PMuRPBxjisI4CMxBL332VwG9H0Wf/pE32ZbqmO
aK6QM+Katkf7LyzuS3lEousxah/k26jw/8m6Q1WmeLgUZwcLSBZ0vvLibaQ434FZChp79MNhav+p
eweyNOYVM9+t9U7XxCJRGbGc6dh3uw+hmlXz6W4LA+3Ae0bpsVugsJ2QPsJ/3wp3MdkR8DEszUpX
DxmSHJXr4onMdCXD9a4hB2NB3wqMEwxTKRiaoxXFxZ5hVjlsa+FAWSyLxEuNM5EG+odA/uvbdx9A
rj+WFkAHge10zpVWMDxXHltfnrjmyOR5gtl8lY6cIrdFaKUzrlokcxiJ1gn3TFAfWIVl3D/jDPvb
L70OZWoyv7hgRTW6ZmsWjL6m8DIiUduL61toLZHtoUXgdqGqE5rFMOKycg1m9CJLCbQfK+h6AL+8
k+U3VnPzOfT6k4Qwa24wK4S0jCd0/+EkzTZGhzhIIVSReWumLDJSDiCRwral7T1Ze4oAMfjtZt/f
CKsTzetEW1M0YOcCWEnK3fsV9wQ098ZQSjmHlU/YMYNHNutcUcEeP2Ee4mC/0SOh3qAP0DLg1id1
7NCBOsAXCx/ga8qCQ6MBlIUjm9TQAtjhw/8chI+Bqi1mMGtjLBeEgolb2Rq8wpTvSI7Xt1l8q3Bq
Hb6dUkQCN4BXLh7VYK4JeeZwyR4k7qB6RO1FzMC0u9X7IlKIiLb3Tv7aGr3syfAAKx6Q6Q/rdcWh
ikewjKR7z9A7vREboRYBjjKZmD7xVwmGNrSE3vhG32pp5bJhfsBWF1rJ6MoBjjZwgSi/XCkbyZxb
KRnnPNIRr/Qsndd5R7yWKEJK1wGfwCX88BmlU+pxIfAbQaXiuOMxWFbb/beLJDFsvMyULy8wg3Sx
ooH1tMRicQ11MTJ7clukZoQVoga2V+TS9JE7NpPBBur8qjUvOySpZwdFVrzib+M+m2mFW8hJukNX
bohN6QndoNUY5EeOE1sgFsiEW9232ShCw6kLPx47kH6UvZgbjWcfmghDf4c6PbWtaVtfr4mqrhqm
s6LU743C/JA0G03yCt6rrZOfEHVUOJvqO7SjbvlP2anRdckOifNA+xre6pmyFT5U9v3BL9odGu+2
VK7+L7uJxqG8wI9ESiDcJP3wFvWILb/UwTTK9AlNTlM0B9OyDZve2Ri0L7Y0f1Yy+dfwdaPZvfOR
lEd8gPxaaEe5uzl2zxOcXT1z8SNiQQyrQt1MNF3nWP0BWLerzGfVucltI3ezizwE/6jRlOJB+PLi
jmm7JrzQGcv2rySj0KEdptWXoXGLF/A3zfZDlIaKVn7MMyq2mnImylnB89yrsnzkuAvl19ciqekH
uMzmOB9uhwhnZP/sgI2/TDlDUy+pAP5VnGEZ7Ideiy64O/xemh8FWPg8k80VgdM93fdJaHkshnIJ
FnZ/p/ClSsyYMXtAZkqIdg/dZnJxZmsJqWkKFPeDV5TUmfY7UTyUQkmIfC6fnun7+6VEmkhTeXOz
RkuqwRObSwjxnbR2PjrVG0AVBZsxR3IDa2gl+3aAIV7D9lHiLDkfGCp46dw7DQFgXagIvXPdLfEF
PCzZIVfi6mfXjKgrZsLyoROiInJAMy8W8QaiT0h5a1Y9cmgV8VFaUMbAOtlIH2sDenm5kz3F5tfi
9eC2mdOBrGOyqrG9okyVHSvMF8TUbNibCczG1I36rUXp7N34HZCMpByCY5WTkQBPh0eTCnjkbMHh
Q/J71f+ReTjqRdV5Udqr18pdrpkKNxNnwAG17uviXWz47N9XFfBau5D1iXKYt4rSGK/untQRjCj8
JV7mVYUZ5WFvYuttDOuEWm5AFo1ir/FD6gTQUln9Wl7bPU+LsjIPGMR4L+pEfPXIJrJOsWIA4gOD
/ZU2G9P+S5ygZ5EgFJwZvku13vQT2udjZJPH565zYH8PoBjczjW45Qpo+XMKRGsT+RQrFb1x0Ejg
eR5byCeyqLpy7YQUlYqAinyQbS0XPiFutLsiSDTpE1GwdMH5a9xA8X8WrIoOjfhglvNIvOP0eIon
OWrq9VQz4wwyvnDlPhm67PKDlcCb6TZP8uaFOdwsOtzh8Ldwi4ydmFDIOAWLbMLb71RIYc93cq6K
3QffgnGGhXq3Pqs1xqmMC9h8FA4pHcHKqSuwXOFkuEOD0jbmTML4yO9F2s0lKZwlvDk063aumgDO
balUYK0lFCABJAuwX9XKFaK9HjRYzcCa+QRS/E9RRNKSPUxXb/IDsI6MJK8V+y9bdPtqUp/6knGB
ph2nw4ejfvB+MvUCsafAdJ+Gt1kUON+w3reXKZWayWJr+f0p2jxezIj4IZ0IF5hbzsbjEmNA4arV
1TejYz25ssk0YLYhHZy7Y9fQqdPfNsM0qPURpEpTpETeqTg44n90+g1Ur1oJteoQbAkAwhszBkA7
O9A47sghtbnLreEmkJTek+BVBY75oCjl109KJVYiF0t1fBMK1pVCG7SOLnIVjiCnu0P0Ec5UvT8Y
99LnnqBZwyIicyquYhQsNmj+Fr7Q9LehIMirqgLsqdG4Zgl7/nwazvHhuTlwsYQ6i4WFJUQCPLqC
fh/dllwrQzEbnHDeOT4u9fOkwCn7p2CXI6eElEnfS1fqDBouSt2mgDyAfnAJw4p/4vPsc8nbzMx/
vCJBTaKsY88pM302Z5+0t7Cuqnb7r+SRKoaIehXE4eZSBrLzTjsIPT8215lskuEzOTXmvqtTM9rf
NWbUx3NF0UUTvaQBdi2WDrQf6dtPRsoxS+2l6KkB9yez65jmZ0E7zVbBtGuS9xCAAg1yxGrQkqQn
W2gEEVtac1j8zcZ1y5kQBpBfQ4WILvN2NqAHicwqE3+fHl79rCEJEdtrDx00H5IfjOCBuDYt3yLE
AFcH8HA84KvzGBxm+Pcvk/pRWh9W/xY1RZFhzsREC/b6eUQFlt+CZtimGXiEM7V0zgkEH+FaG83V
vRc+hRFJVaYBr4rHUjwVNEC0+p+k6yWI34jYdUxMnZXLxgW6wgfd6i6YID4Od6jCEA4lJROvnkJB
duvh4c/p1VTuWol3VE0Skok4rGcSVkCkcuMvT/XMkGMYe+dFKK0v3UX3QLiU3d5PfS7M/BDKjQiT
VbaZZymDNMiE2fEQuuwieQWwEuG2enYLkulsnvafZ0FzqWI9rMX1KpMeT0V9eplcT8UyKCu3dVlT
BxKsEAgg3CtYf6SVGENQjHwcTo5mQrw2M2XBReFwACpJ2cBQK2QWC/9m6eot68j323eRgBOd9kEc
b/6nt6vNOKGqqk4qt4w/3J+cIug4RCl30mVAMfbzE0qnjmvbUjo9b7qD8E7dlspnb9ZQf1YbChuL
I/d89/nHVaovNjNhy0URmCFdTsG2rGHFTtceI7MjWcuvNkCRKlIYXC4+7jaB7Axec46V2qZ3n+IO
e7BgEhwjK2S81AGd9neP8P+fqeK/Q9Tt6+hLTJ7FoBfYEFD41nzv3M9jAdHj8i6Ggofp8biIK3O6
UhS7S/iFdtSyTjotDY4XtY0WGjB2O4ps3BIOyCjYNV/ZHmPb8tM9v7dcqTeZbci7ia1ERX4i+8Wp
pKdwBi0TrZo2/6saTyf0UTC9G+SSHNEeKPA8YsgSiyESUUvy+Nx0k7doVorJetihsvo0ogc+k9JO
B1zfZ6ADw0kRL0MY0LnglG4L7u89Q3TRIe/xZCi10we7jBTpx55idSeVit0X014IznXDyWlBNRrr
pccvXCR03T8Fw5IR4sI65amHa03gZWB3XMvZRFq+IqpCFIN/ROUVoT1KXNRRc2qxUtJuWZPTND0z
Bqa0d/AQRsUZ6IMHtbkrPX4wYuDz5m6Y7Pcq6wTJx4NfFuuu3R5Jy/FdnOLlZrjAJHhZa1B4Snqn
cq3APoC6b6crTKbrtgX04uYwTzo8qYmBpAtCcqJkB+9OOrPeJuy8HGnbcVK/E8lkMe1t2A2Ts2kD
IFrOZbh2Y4MgVRwLHM1zl8Yfq36KETcrOoGaq41moAmXX2ltAuLTfN9qjdWBWmsi6LH2+Z5pBglI
U49OGhgJHxqrfp8SLsR9Uv9oN+jGXOi88uTP0ns00Mbctun2pn4juPG20crPqZUEQT4bnnZFnjAN
uLFKBpWhIWXc6SM/fvkGZKcXc9xUhYQ9nWRTDTD8x+xQO2/8ea3yeSScjKsS14C8VLDrSDhjGw10
nTV8yLuIJ2hn5bjD1m8S9nEHl70l+J/Qb/oJCx7Wd1KTIbSz88/s7rptX6Vagtvt+cZ8ahnLKAoU
e+KEjaYNkv10k3DmDOgw9wjRlwAVT6ArjVDv4bfOIAwe5SQP+9jRAFzG0kvsGqlHR/hQHP/FQnKM
qsGo86Yjn6RMjm94JHZFiXFgwZQeXAvvyg5ZsxL0PtAI5eE2hB3vVoEDoH2b5egkl/tLb3lkMVu+
k/a20+4++19Ab9jHVExuxkXSIg4HpRiXpmxQ3BwpxXUGHtJoTx6ovXFjJjuYYKRVvU5vA0G3kQiO
pYqLm9PPFT7jCBqekhCp7vp8iCrAgfICiG313XiAyx0/jYLWn8J/ovwqA78ST5Sfzbsc5+s4SRjY
RtSdVzKmGaWVhO3oCwz7SlNzB8JW/GCOcCP7+EwZ9BrABHtajQo+e9nke94HhQUiJzcR/w388jOl
o5/TLfAJ0yGLQ+x+jZd2E6o4Vbr6y4MbjI3g80KCSwHc6/CsZqhB8bqlX0cj+3Zl5FCqpiTe1VPg
m4BDSNqy+WPdEBOBlta+ZQrLcZSpUYO/SVSMizxE444RwVYqQjEKuHAd8tp8slUNoeqA6QgrU0ny
aUpoCqsTafrXFy8vrDiFmuK+2uE158Cl+30PurzvdlPcQtWZ6LBgNpScKrUU6V9rIGbUui4kORt4
2xS9Gzkk+UsdWQKkFesPHIK5vkK6cCqvgTzuhZCiBwhvBfkIiKjanOimBEAjOGnT/HUwrYAZdxBv
/xtjR5XsWlS5lwfTB4O9VBQb2ckp92MyLRK3BqI6e2YTmmqjLHk41vPU+kk5NsCj8/fkDRs8GeTd
C2v2ywTOrRMwnR7SjEuV/KhqRlOa68xywb8nQEet8mn6IJaJ5m/G77yIrX50VTKDqrysK5KFU2sw
30jH8vq1CGHNQUKfpHUNMiJ43bhI0oKEzoJYhKe6eyCLEXTbOc3yXU4HXg389T6dJt9uSpY8+eC7
7ZrS7XbVd08xYHAweUi8XULUiVh8WATvt0Bvdt1ltkgzG99d4zVsh4zySTPV5IwbuwvaNOLmeGC3
u06J6DcSoeCcQF9CrWPLRUEzduPVJgLz6cgGBtrJiZG6jSVqOFYlXMEyexdaWMak7gSjdN5811Uk
tHeQnRnIm5Sl8g27UuHzgQ9z6TcRY8BPUI10rP2gHQGi/l5N+pOomHSELjGkZWZXiIiSKMJjBWI4
Lcuom+OUdkcfnla1dGD7M7SNOw+vq6zTBTw7Lrs+ukCRwM6H7p86JqQ4n/W+ITThO1JJ5FYfmggJ
mWSL/YwkxcIGTROs+ShUqb2YO3UMcK+2CIHGY+y1Dx/iugHLq1qTe3kgRDpCX6Xd46tVacZKfxmK
dJpfdThAXRHa0ntGeq2zOUe6cAfMb7UfB7NMTEhBdYRV49DYT+HNVkOjZQZBSlGjX0Wc8SBnT6KF
UPgJ8p8J5GeQiU6wrVLzYzKBw8+/xU2LUkgVnU+HRyb93TYCfB/HWj8LzjqGOJNnAj3z4BTTftuc
jpId/dbEAFuBneIH1ays8IEEPYzr9stbA4/ZSeRorLnpMM/nEMIV6bxFfvD5Fc1ml/wU/2dQCkeH
TfPe6amkPprtCxthL/RchnPJOMu4eIoA47rnxI6KVmokwPapY4sIULN46Omja3FICv40moObY3nH
jixIUMWmk6FzTqd44DAatY6OnYrttDguZ2nvyd46i3ZoO8CbuJdFYD/x5XR67hbDpyiV/oWPsKQA
iGAvUJkN7BZ8XPhvGXOrPSgBsZz0NYrD0T/E6Go0YcASVKvCuqqO2wZGuVCLbiaaVFu3CWghOzCU
XiWPyxgI9stpd4QL69WuSG1Mp+rlCjpDV6rGi53OAiYqkNTsDJQVIhb6yf6cMc+beGr/v008qtnE
WFvDHCmK/ndbL8cXrKkHeBIy+1LrJeA5hZBqS+x+PzGHGrS7rTXsR+JXe9zvDgkgvopl/Ak6w+FC
9norUWWq2bZLXSWs7qvqIOM/HkDUfhq6ndWzcKVJRe+O0t2POpSOsFNg0IcGcTVyVlrUGGZgRkbo
MbxFl6c/q1pCNhxUn1yRkN08WpDUjGmuZr5qy5WaVg6AbmgiQaCONEUXiZnXWXAD2E5gwjjbI0Er
gWgRMtl1H1z7OwYooIR0ns2GtuHYY0DltYG2+pAhqiCy+3qGGDSqn6KxYe1oms7rYr+1HsZanEXU
LVwQXQYXqrKGESOGtFUJvAw+icAwB8yN5eAHaShxqn8JoXEs2ijsDQXTrKaJQI8umulCioWa2xfE
9V9y5EvIz0LqEzyD5rIZaG3wQ+L4XRWMAsrvcGDN1mW68RtZm5geHgllUyqAwjrT9RhUEpPorF6Z
dDHxY2HCzwzNtFCInYGuNI1x7qSZ7GomLFeb+yex7j6yTo7hMsmo3vtRqN+5/Y/GYoG8USDK2aew
l/ISa7rCafh8btEXUVZXTrS/SuB/ilvi3zBDqsw6yZ0wH7q5u7shrEmcKRxmigj/e+NE1UPpq9WT
JRf7vqx457CV3CcZ6BpT67VfQ68DenFU+bjYuSTb2Z4/k7Zo/CouGE/GDlVGqT1lQ3QjWm/slbKu
RJpV4qv2aWcKuaoBOX7uE5NDqr4yvh6sr2kQG4g7Z/S+E6ObH9bnFsgXFdJ8ai3L+zxtLW1WFJZM
5KqYjXfLRppBZuAdKq5rKemooQ+iVDUIK4oqKzPzgxTF74AT6bjtqAUrQn+8qcjZyMQtQnTSCzgl
QXPoV3zWzCCuNhESfse5pnCuZwLiaMc2VegECGcUwQHa6hlKT8on/xufiL967OWELkMu+X00aoHk
ZL7o1F0PaztRSP4Ad5xlvJlcFPOr4mR5C12qggBPpHKsi2YNw1i2GtRt7gp8kTLKS45AlYD1woUm
jh+1iakB70cAn/bS7S47iRr1mlxfC4rXH2n80qunOA2vhrVEDOFsM2f4cWtoZBk1qqfMl66f01Jv
Th7Cpx3OU9HR9/SzkT1jINEgL3rYlRdF5nzBheUgKsZQxWfRs28LHgGiEGNqXmOG5iHUtWNup0I5
rqRiLXp0wKC/lBhgAORy1IoYMIeAXN/WBH2D3RvhZnNql7qHBv3LFMOuPDNJEozzFPxWgvLU9sNL
hrAbWgo4yxUvxOd6BWPlFt6pVcgLxSso+UZOXFhNSgPNqVaUTfKyi0FtU25WVw1GVTIrFxLTrYYi
45N/wwrYR7fjdpHWu8JO384FOCFqubwIz8XzWCLkjypIp7NhTtgQBDzEI9Og12BUUar9TqMzuDy1
A7ey2YdPHMjVViv0ksH827IGCfN8j9hD5fFLOX7cJbDcTFHcHRqT+N/yBqJU+PlN5wInNYBQ5a4p
aDjJ2I/cHDV7TPPJV60m9N+50Ir00vkJ+jYmlp95Gvw12c+9x33OjAzUwXC7dAXYPl5V7Mh/9iSI
INLnweRfDFQtCknJgHymTNYIShleZbYp/hjyU6KhgK3r0rqRo9fopugJPrOvk8wpNZdHr7wv0WOL
QvJJsYRFYFmJ0Q/ZHnn9lxvFtCjJ/OYr+P3ng1CB6IPVjZqROQkx65f67AFFxCaZKYVUPfNXkwDZ
2pXgEm8spr/ypwUizM78izpFEzGqqNnOXuyJ3nJKK73diI+T4kz3juAfEt/0swUZZqjyWmumkrwg
YZurtvmCyJPdozqPD+3XIb5Tupg78efwnvuFIvijIKdD5VBNJ0SnAU/HpnHz6gSYxb3Q3TDvzwrS
fT9G5wd0U8etWHO3v8+V93gziqPj1WxX71DTa901EItgyaxGx+TuBLVJ/DEV+WDZjrgnsPjXCbXi
L3J7QgknEgOX54xKoq4OkjYCYB29dljZgED4EGNNGxEQUsHdVcqXpk3I8p4Y+uqMg3ovoZlD80Vc
1em+qiHS+jMNwmPKAoIkm5tuMr5zVgXYAjC07Kp9YpqREkj0CG2rMv1ZJ1Kta+lBdyV9Dfp9AwzT
rVbCVW2karQUVD9xn6n8Vy9eaG6+O+wxZzE1RUhRNSaUYxV9FRdkG9vQsjhsxvtSTabLVX3HiZY/
PW3oFdr1dFKplf4PFyvRLacc2gw0HbShk/ExUcLsaIr43k8dDBGHtwu/4QLArlAwY86tXibtYZoL
0t6lLtHKtSjgIBUiwmW6D/bjhuCKOFFOz00mPY0Y+zTCut1PNjfF8yCz2ZVgaBg+MoY/a0pqhYoo
lXvuXY+6G1LwYhXZOratraJ6SmqFsTbzjjV3jAzZ1XvqV1PPFZgmzkaj9du6Hb6uXpJ1cP+5vZG6
vh3MKX0ZRKZUxAdArPiR3ZJ4NBU/HamfwVUf0lPMfVtRnjCtMXIMVI8IxCmShIpfc+bLai2sJjd/
XCTlMS51tEiCq3+/H7sNzio7Hb8NEnpfyMEvmi8+yS7BRxoF/NLniS35q8FlU/XASFoABlLd3rIv
nKqw4cKXen56bk4EPMq00UBQYJfHhGZ8jOs8VR2BVUrH8Peb3MW8eytB/ZtsIMUHSsQgfdFGZAJ1
lQpXtesleKJ/pytSsRTcRxf9E1JvASp2iLWL+mHjC0H9LRAJKNczvxbeeZtpGN25GqGhsDpFUgVQ
wrHQKwcopxf+t9mtmQz2/Fj5s3X09O0CqywfoHIaprHlPBiX8R8cveku/T0Z2OiPbfu0AOSGSoMk
R3O5T1etxOihZPnDnsDIiBt99odHaiU3A+0t501OzDovyny84w+lLPhkX0bjeswulwe5ExqSujLO
O8Dc69wSR752y8L8djswdlM9DQXXjCQp1Se7S3ghaWLsaZHwOs3OLUo3dpcRCpQpuZdoiBDGXEyU
6YxDFUVjfrc9tU6YEBkFeKGNo03U0p3w1AR4ia5/oU6v+1machgL2tRVcDHyzbZFxuSAlN1Dc4mF
Yz3ji/gLKkjNQnJR0x4J5+qnCd5CJBsdjhdGKYLyX3t03Oesjqdxqh7taiERwzNFgcVknFSbJflL
Y98NBOp7ziPpf7X4jZV7cq6Fr2dIJ+uY5SypRkAgRaEsRBKsnri/mmP5VorI2cOF1GSG3LWyKg/p
O2phHR3IeurTOTqDK9Hzm+suOHcHOY+z3n2iMxICnvK0uEglkwPQnqq/plkxeDHMaOAwRc8d8pyH
kThvfQWYQ8ICERQtsaFi9kw7lg4oWj8fpfIDW1gjA+HFoFs/PAJSGlw9xDPV+P2kZgYQQxuPrtz4
psRnNLqZ/33HqfpCTnJ74RiXJVKl6EziRnM8MlyD5N/U+rAukFAoSa8RgPEFmtgaYahupAvVdQsw
cdcmGskWX5EhXSQK6rufKPPN8NbDtNmfGcZ0V/lt7K1TkPU2z4mHz0YBP2Kl84VBnhamA6GNUENB
XNGuxpU15zl5INTH+mq7BPyekXMOdAiu6XbT2j3Vs+kTCxNNT7tyMMTXZeaaFegFg12zVHn/HiT0
o3PCpCTFxBmLIo2X0PDPianqNs8SlmkNNs52lA9dC5EZT3ZePcnIZ46P3U4FM3v/7Pzoj8Tjv80s
4oYMuhA0msVxuflhwG+RfXy/Jhw/SeV//epN8Lq2f5en06kQ7nU8bsKhKPegWgIOdSzcWIArHC9A
KFq2yloCmPyEdKha8lWFxCrGfF/tDEVhCLDjz//1ov0f0Fr6r1ITnnW4hFWtuF2I+mspgrgGSfWq
XfENSc18KcqusbeOmWVjDFri5AA8dsCuqIeXbq6ZKBxTiGPfrfrP2IdzVv2ICl9D2rrx2zYMUSGv
txEdC/Hd49J0YXLBrhLoeaBwzieRVAAcfT4ThYhs2ipFllUvZO3TPN5ursZ4FKjv6H0WCSDc+4S5
xQhpSTq3XcWpKSs7ZinH0q+1YUKxSzF4mtWnGAcqACCDw6iCWY2/xccxxQA5h0kzC8WQ1L7HavPN
Uy5JgSPhK0VBexzTmvW3yUmWim8mmZ2BGViyVRCGmqaO+G738REQgZwuQWspEIwbGERmk3YyAlYZ
2znwpKloKg5Hg+Dv57nRMzxOWhIj1+CNiCuJzvFd7QCmp/82rwQ/htsCPDsDmFeYCtQ+BWB7ozxv
Df1RKrnYS3obTfzjWIu09IZ7ljws32okHQNDljd1OJkarOUHSpUuYeGqiKkchpt5wvHcU9yURvDB
xLQwxnsAV3CxMlwW0CPbbNP6PjtNMsyA1Yze5znW2JmNHdb2DJLMephYd3r7cw6Y43NRxa3wcMrp
O7RfBAtvZU19BrfBLKF/hqg1rDpWQqh6CwOJ2yP/axIQ42UTa8blqhZNpWAC8OOjgzAXSMan9SlF
NLbkcDV8FAvjkBTbxqj4V5/QE+g0geX1E+hd1Ej0br4WIfDDIhCpAtjNhBEbsCkRRDPi3kZAjEdb
eC6NBwCy4SwFG6kDQIBtg/tlDmZO6N+0sbNSFwaqMz9RMOFANxZtgSiLJuKOqFbpamehDOZRYbp0
36wSXAX4SiihCWKQiMrUgGKlL7CaoU4AyufX6F2NwCf6Nrq6d3wI7+aLXItACyeTxGhbbsijacks
xLRFQj3L/USVhiJCJTK6yNGaHYW3p3SOgABxxO6/3jiNCW4ODT7/pRqhrnRtj7yKqJigv7ZBT2xY
69ort12EtblpIKxGHjifs6zG1devcMkklkVvegU86j8pepRbllGZmDFuBdXY8W/DnqNcjCwKGVIO
IoKgwY3mN7BQL2taTr2HNzspQM7n0EoI8UNaPbH2cPVLxKlv+BKdQb2tJMdMa9kPaUBRY35BTX7W
jUoaiPCuBwZWMphAnOtbuBvcFghiQj1Mi9UAdYJgxJF+XjuUoaXvrkkYIYl2TE2GzBnyooU9svtd
h0cURXJ/rrimrDEGwjh29mnkZRdLnbse6KEHIVmpJgCJSLmacHwSjq5jSCU76jfmhyEts0m9SAUB
wm32HHX2cb73dJF5EYh/hqI5qFXaEZR/QUXcL25JHRzumNkV24CnzAO8Ow/XbTVgLwABeA2/ArGn
qcF2gZdoxiDMvlYf78V7x+6d74lZMs0ctGomMnJaKvnNpIXE8wH/CHdFkocpH7zgpB0PLcBJ+Ush
74jLrnHWqz9gBddNn3ZtuwLmNQ9HhtYrOS+llczhZEfCaJfc95U7e32fDTWJql30Ecm79kjv0ZRD
9Iy1ibJD912Pisiqj4DnY9RygWJlWEDTbNIALq3N/VjpcPxfssp3F3n2lT0MP2WuYvh1HEve9m+D
ingHO2oDSXeHcqWAHuxwXPAAtkQxJ0zHQLn1fbJMEo84p6t446EN9sIIwaRwbc1YBk8dLFozbb9k
VogLJ/Zzvh3XDkLmjqbc17BqMpwGNq8VA8UYR7EwEA1+iNnkG2rYTPtwouHJ1AQ6T/D4yhj61vng
/ylVrxkI6qrrNXE8nIhDR7LSyQ/OzdOELR9UOPCYMp8oxx+2AtGBrgpaBpd/vS4zMoWozL3FxlrT
m/c1ZTFdL7NSHdrGhJ/yXFPeYGwmatwZgD6Fynf5KnGL3c14cMM3OPdk7+o7YyVsO5R1UoZTt8/c
qsk26hOB3XJQs6KKjOrcc89yKAkAZjo6ul275673Bca3+3mYth2iJa4VwLyei5tQZDsCD/Bt20o0
RWF3nWQECazfVi3xNhYXWbolTpmipIBk91+rdlTGBcdspaDiZOhxWryFH0DlAQngK76bIA/EqsPl
xv9pRdyvCp2nRyNP3+KTgqN/tZUJ1TFffav/dE6sMBItueeF01j6AsclzvaTKZuYhAggGwOun2Q/
RhlcYDd9KQm1AL/UbCbSLbigKhpN7TPV1Gic3O33+kqDNwDvwG1gc45WahkIJps11alrB+VCYL+8
e8GRQW9PnJOVVRtJJV1OJAfOP7IV+i/l5k+K3OGNwwRgL47wzvnIWzk8SPoNyhmtfRIqSHtpvaxX
RA5bBZ8TplNVHnBtScXYiQAK+hwAtyfagftlTvqQSMA8x6qfSS6iYpx2nTUJyUu0V/Bo2QRlGMqC
itEztK1unHtaqr2jlFzuUSVqZquTHDjzNx1k5LFRQDWp7UHZnNxhfyE0KrlgghIx6MX3iVFUru0K
hqpzSaE3yDvB8iWjRYZT6bAX/m9lWjEJOlmTr1T6fnaJVDRR+8cefQxtyh+MUnH/DEkgeOgulcCN
TH2KX2fSmOFn/Lue5UzcRYsWALhXz+oaTjUPZEXbxLcsKrLv94yAuzjkXer7OvrWtFQE6ETCl/t/
Et86fylMBZHJVg137jbjMgEhcEV981FJjSaYXNqIMNf9/S6E5GgujM02rVSDy6aKoUSQLOehjR+K
T1F3eCdU7nQBTh4RMP8/OmHWdQFyLAm7JtQc2bgCfeF7JSgwgCsPtiaWPBtHQnQCvDCoprLyby+N
rwxe+FtWtxvdB41LudC4luuJHAzFm6rQR54QnQvI8+erVrdd2oMwYHB1Jo5UzRnhy+FOwrdbnu/6
LbevkLLXXbfe6Ms5ls2AazOn25fn2XA2FMl0l/1YfB/gqSv/63ek7Tl5HqTCkwYouwrcu/sVfTn1
V+JOTzagWFyBeJsca+GsBVo6ScRGVX7frcPidhXqfHRymdeoekHWK4TfwaqULUKpJ/eAW5OySy7e
nSctaxohaHZRoebMbV5FXDPGDlsOP7/YoNxQ6ZlAFsoChYpbgWGhdlDaAX+O20ROfrU6fQJTO9OZ
PXSWm/mo7tFrA5vBOaxbdb6dCjJBqnQNFBbBl7uktrrAHYv3/+jwvJc9mvRhxiUagLCfp6+OGybH
Mo0cSqzJsashDO5UgXlOIiai0cgZr6ROmDuO8RYOXCOoDhBq19sqgs8Hmn4wuWRLn61CKOat7nMh
d0YqTe0Wi2jrLZf61aMberIWXcHa0wTaj+Bp6Ubg5kOKubZDRU2FGD2oCXO2Bhnlzg9hidHahtHv
O7juiuk0wF0GtVRcjaCyOkcPaxAuKQQI/spRO+42/1yugGPtj4WAC3/n2EUIJet4z9Ph5lDLmByf
xiOxHCWyTQ9pUXmzsoCth2R5Si8pbdfNMrVJc5NedEpiMrh/NJaHMHaZ12nwwn+YZKRE3ez7diXA
22dNGNGan6L6A7siYoXcocWc8DGhaVsvwmhajnEFo3NUH8JhI+ruU8hXYdY00tI5CGPldR6+PaFL
bEueSVM1XCLGkfB+iwHVrkgPmuhOxQxy8m2LGIdLddV+/OafKby1WhW1RszPdnYW1jTKC6wXCu6Q
axhLrynekalf108GTlvNQO7OMbYFzkAsSyT5GjsixxedOP0sdQL8B8k/hD8UgqIWr3VUaiuhduZE
VNyyPWmoYZAwQn6WNDrWznlJTzpYx7As72zUVq2eWVQ/8fsKcFpM9yVbIz1wdp2IihFVA9PYxpLd
Y/SW+7rswJSwu6poYm8/LaQGhlBMCKTlf2RBkSI5bzc9t6gXRlLsSs/EdeWZ/4uS+ZLAThicN8E5
1cqZxi80xaHiaBoPQMOgNyN1SRcX0cDRp6Z8Bvs2Ei0TjGOW4VUWgLbRNsI17HsRqxQV8NB8c7t3
AOrPv5GY1PN4xGFV53fef8Pd4el8zIwPknOY5wixo48Besgn0F1kcp9wREJdAmGM3E7OF+xd1yMY
arVA2ivMO60RKgYaMu/lgxn9ofshPkI4UoyuN/su+0Xg/iPArSkVPg47MaLMDnFJhjgQ8BATLJB9
wOwq045dFO5jTpgNqLB2Jqs4ycluhXBOharV2MP+allCH7T/2agNiUCOXX1B9Wosiw+nNvtQzgsD
xoBo+Vtvv21CV4r/awGBrhMP3+5dW3z7ib0xXLihgKwUjTfHKFX8Uc6Z/X4Rk1zAhwZ0RuLH0KxR
/YlZzN3fZ3GDHuC2mANmCtzHttsuHtY4spP3q2Mipq3cU8P33V58ixHq5yH/4HNNcC9T4JJN7HHV
Tqd4+6h8fhks4DWaKIAIZ+ikgImObJpxaDYu4r1M2D1XBLo12LuyNieNWAKkpF9iiIr7ycmo9DPP
dc0BSsLabh4VF84A1Vdrj+bsQ4w9v6t8EZ11VzO+nU/eANwt+Cww2kVzhmJytKWviVVW1/U37xjW
wCNjjgj3SZSayWT/dQU2GYrM7z4FC0wqjX4pJyXwYLp0tKyFsLM7m7I36uoqKFzhGyl8UiYl22Lh
VYwPr1EwBrnybSNLosjyjEJ2feOVxjp96V6HX9Bmc7P2sxY7anMaktvWZc9eG7xOut1lCcfKXEwP
G3OVyQpjmaCaGmTb2y+g//673QigjYHFnbecmF41G/H0hHONuvl86UXpa9wf9wKXmYQx1WCasH5a
m7/7dzmbmPIAr8Dg9O9KRN19r3Nip2J4nf72katpf3dHq7DrOT0ABXMPgrRJ/M3vfO4pvS6MHREE
Jz2x103kfM8t5TU1ENRZi1+wzEgOVvDIuX4RxJxEiOpMIH8/l/JcBOOQ8pI0PGMe8etc4vBw6tHZ
unenJelAzx40NfbWdRfZGFE7nXWE7OIbDfN0KBUvk7adintE38xggHdebNJ50fBWSACFPKTNS5mk
3ZQw++ZUg8mG6a21Jjdc/BEbCTxoFqx1NXxAwsmPjJP/TjP07x73nzFrjofiPHy39KHQwvMubCUs
kcIZ4miF6Rpc9kuRu09t0j0GOsBMX0Qjjrd0gMCwMNwU8P3Cnkwkkfub+JELXBxmoofuuJ0LdqYn
nIilztkFGBzYD8qYSbAHHRmcNoDCgG88a4C6GtV48WBkJ3G3O9iNoOCf/BgubtkxJ3t+Bu3U/f17
JUCmI3ZA8HsNiXeMb0yOLrHADq+ueO8VkRqrWvs6sItOlfUKHRjyu2TWrL0m7tqRozEuSqcynjkb
kQwjbLQ8tD9nTNmQyna2Fac1mKtBiWEBmmEEp1b2rIE3I/tFwcDMwnN/CedlOwyw2wrmRY6w8lp/
xBKokdeBrOIFuY1HLM8oEyQ21EOqdrc4XLaqk+/CbqmzBF9k+tjFJkHssh6r5AZ0rSkjCF3PltOS
M1UvgCVWP+PeY9hBI4jTLH03SNHm/JRzkhHJ8co4iI8Xdb9/CZIGP61u/Gc0yQgytuATvEeRS6mv
az+WcFifaYwea4fZKdX8PzYvzGInDmnNPi1K+SQR9LV6rfac+kfOn+tcSCTysGQdlglAZuR38XY+
9xn9UOM2zJ2ialF7UShP6UKLLq/1AZpoKtBgHF2iTcjPxE2ct+wkFk5NHJEtkBckPKKrQAWLehZ8
CBMS/uWcxZcS9vEYVPsYPRzxEuy2jV5gJupTzGYxRxns8N1ms6EI+Bc/RluRb4RNuvNXvrKeCp6c
9B7uUXvWhF7/kKpDe67H1STt3XqI4iVmIYcXdctdqVhfvETq8fYcI3lUh3XphO9H6GAEfu+UXZdb
jN0C4SBaZjTDIqU5G88je97U1RwIcqV3bwYD672a9sEteFZLLSMY46aiNLmkuUbP83e1GjHSrRET
snfCWYZWnX4ppDnhmUGV+9Gix4zBDbttx+zTXoUat8Juc0hdLqhUGWFV1hyitrLqQ9oHAcTB8hDv
5UeiM9f7kPxvy0ih/lEH9Q5N63a8owJf0m6qOWJE/z50ImpUUEGehfhAEsnRpym99gOM4jiTE/Hx
TO5uk/z6WjiEXLBs8AioPqV9MhAkDGfVtsCs5UrSP6Sd59++5vyv3voZm6FoMMkW1XwIINSy5uhV
8eL3RHDbH+TDOQZF5fjsdGnMhM9ZFztU3wiSSiwPczRPfNiExY91MCFabaEx9FJjkuL376bm8VSg
TCCDn1CvrZpBZHhmHBpAJtcx2Vn66uZaIh3+3xlBJdjq2asumi4QzcO/iFw2PQY+jZvTb2+hI/H+
1RJC8dtJC3/0GqUgAJA14nG33yun/iL9uAYWBMAKT58tpqhgjsC6kT4Fmb3sKpV5Mjhfn4f9hK8/
rB0zQa85ujt0SFAqryUWG6KN6up0WZqEkE9PImo3lwjllQmoRKqfeyG9u4Xnhsmc5LNbEGWOL+pj
QxGV/3AWBsPr3nwU7s04oejZJ1a/fiVbJsQWrGTe2m2rtzMihzaauVEgYb6TU5rTqZhBDSm/YFxR
nX2SFs3JWL5V1PrF4VxI97VATbmD2+fYOg40P5JgumZw2WOL4zYn54kRTg/Zn8wvyGvUlwlQpYKy
P43EVZIWobwrIzvVKhUSUF5+PKoyvak5ibEKnfHKmd5PoThJNyJm4QhF6UQW2PwiingUBpqIGP1I
swr54cuera6dNfy9K0noVAgi4m6J3G8PDteDed63/UcxHu/JVoA6GgvoXg6SBZrTlIWHUdnCPyFz
FTI/i5PI60N8oUK11Q0sIkt2iefTAW11jBuOmhi+jTP8DioNLMsLXq0kdYuWCMXF76zvmsEbix7c
OC7gZZ6Mv/mR//LI3O/mzCLBk8xODxBufY5lrKEAdjdstGZBpCf1kXNqYXSpZ3KeKRu8jELhK7a9
kq3taNCqHhMpLl8f3OmSsAfky1JHkmnVSWAZaxj0j8chehyjk7mSEZ+S/+Dy9KDJUwR461WMKXFN
LoIefkiKfurGhIX2uNmKPNMCCo5Y8YbPAHtz5OJnwfAhwY36VtvTzEx2LU8eKiaumGetrLR2HXKm
0ewbC9pUVAgIwe1A5QzkMUD019ScvIVff6RbHVLw1jrZ117wEpxFAEmfjvwRYLCtSHaryM2az3nk
ozbnExw5ekMXXiSkkCtEyipSsoyltUjkKPFF1qgPJXX9Q+MUh9/HAihjfyZiiynZNKLeslO7EuPK
Et077hkftr0LQ2Yc9w8rRz5aDU5qEZmjttLjz58WIgSFRGDnW9EMWSWcyOof37321MB0VZtGhqUF
p+CajuHPW7TTExXKspJncSjOO9HhY78onswgkaHC/OkOjPjhOXAICA1E9KlMLU43IuDyb/0kQMxj
4hpMjfz7aYASkqtkdb7KP2KDgF+TWVQMigSrUgAhnhdrrE+snDOPEzBAs4qd3bLY+huD1KiZxD2O
W1zoOT57RIxf1dkdIfM0pLM/lkyMcTxnZHyYsk090JMJw+3hFroBWuLB2rg++09hvz/IHxNMgMbi
sDnkP7vIgFGBuiebOBu2kY7SEcGRl8QCXJ3HJM/1bdfUfm+i4D6gmv5QbG9C6S8UprwJLnHpeeIZ
GCCM4oQoi0x90O6kAhCd6MLGwDDEG3lep9jm/k1RnmJVs6LVYg1tBOKujduX4+KvhRcDLWOz48H4
FCKVGsE/r2wjNhp0S4PQSDvAvxc4z6RmM7n8o9hoT+C/eqC0LxjpbOaWiqgCJrytjIHVtuCBxqb3
+FVVXwHzOCxs1eozl1J3hGaAf4MDiDayXgY8aQYGiYz8wx0TNltW9lOWzEpsd9bOlt832HKERyBE
PaM2SRQ5QLz422Z1W3c9HdDlsw41fCRykx4m3ye5pH54JXQ2Cc2zDa1f2JVK5XcWikXAGnMuDe3Z
0Zb4yZbFBfizIrwPYFxfc5QYeoY+52MLgQtQq1iEW1XLt84XF/rxHTUtqoykapkbGh0jc5P3mSYm
XOCFFJ6Aso2/De1GWLz7HOHyIdOaBFLoielFRZecvguYtcMRQQZuvYADhsFXM5ftMnC6HrhBJ24l
BQaiQYZPLIDLcLVZXfV5/cYtBHIg6y6wxOgz57fXfNCwD1ufzzkndewCpdBTdl7P1nODgNwYRwrq
cse2im6s79XZ2ybeM26ja6utq5mbjAkXREawY4Oy4vohTZ+sJiFVThu2HVIW7ikrQjyVqAEq6a5a
aOIDjmbsW5Y7nSjnRyT4rt8v5hH6dvEjgPPEUcZZ0CxpHe3x/4jgFkIQvrb8glaHUNSN7al71soJ
mMUDU0XAZFnstsdjgNytv31/DCYtDJyTAhM860SpFGG4fHcN6GA2Btz8HN33ZZ8vOtszSUfktkc+
IVuQ0xyAdzqq/HMRq0NjQ5dKCXApErP5vTU0Vi6Mq1k4SAfBvaiX1k3NLkipfZiQimyu3KXGtsg9
igsgf8b0jPte84d1DxmjfRHxcZ44fp/OZb9oOTGRdCWanyYCPlFXpw2pyxvVsgDLegbT5eEKq3s9
4tVRwHVvaIuc5nKropyL+rljXslALOnsmsyj1438buoLGETC5ykIwovQBJw09xoSNhdUBEFsZ51b
O26qn5GPTayInYAmMGvaUANNypzSRtxmljrwb7FR7drbPiYbVGUbtRhWFK8M5ovWtMxisBh0jqJv
aTDNVp/xPpoL/8FMIhXCKQONqyuGPNB1BNG47O8hiuOx7EGySzMSdaM+0xqLOE1y7UVWT1BpNPvb
tdFEt6I7vsZi511UwUOiIxr4uMNsNw/Ag/MLt/H3p3BS73Wa/v7FbPA4BhD5ziKR2sUILhLN/HKF
e1koPI4mCRPLElbqSY6cbKl32vYipBqWi7yMrbLlI4W6Rj4whXEBMGOkNhnFntJdKTbj1nTMVLse
77IOhrjV/pZNEchdj/YReyS2doYP313OhEDx+AinIhptSw3TzfADhLmltj0940r/M7mvMy79XTPb
6qtsNOYojd0hrxTBj/7sWIvovPY3rf02Rn7exuX2YbUh4vnae7e1A4/AvNJA869HopclSu/WTeNg
lFoMDXGlW0yxhdmxrBdo+lOLY7jIz59Ph7AQuB3Oi2Se3WMrZEfSUPlJznsRmorv93pVZ3PoyHbN
O1dJZfLPTaGbTdjniD8cyGLFDJpVLCH/gZcMMtJMDPdGZ5RwfZIU5oLRGWzgdAZz5zEatsTLYUmH
5ySiVD4UY7FhgPzs0Sq5fSztahdl3k4esh8nA2K1WRXnlyq2loa0a+FEpmCKLqU4Wk+48YAmnWVI
jgil1htpwaQDXcR7hhQbdpZYg6D2QffnEp8oiT/HZ1XSxi3xycYOQhdLsyz6w89x7LJqZCKTWBRq
TbXR2YPWJaih5jv5nZuyrcZCcGIkUdsVBtbkMz61xighUTr3ofX+mnfCQYJRSDamXsliRKAWeQnE
b4KUlOhoj3d+x9hGAYH0jUeUHPY4L7CpCltx/v0vFcavhGQyzNh6a9IF76k5OPS5DYDaUr1cAXa5
IV8PmpIenNtLj1c5SZ+aSls6LpZmlaesWMCKMBMLcxgzl1IgYNi1DJTyq5NH9i1n3wDRcD+w+qN8
jBdcpqi5CTJEegmzJ5Aj4EwzeNjsXAn4CfP8eGjkHu4R8OvgDbEmjBHhdBPIihAmMFDPXJyr94IV
11UOphW9gEZuQhCd447H/YIH4M/aoAH7eNiFJs9URkaiDFpqvuBApCx/qlDS9ZTfVXUmEZDtGBy5
nwcm5JcjZNz+y2xvChXIAWKgij6MbL63tZfzOjkhhZNMI5jyfbfw7vv/5+6L12G+yxx2G1/J3w+y
5U4Xz6HSxSxNbEsojGQw+lv4h/EAX7dEQJhSRfIF7sY/4WOiP6271qHKnftHFJoH1dCHm7TjHkwx
zXCamNqbFdgw7s4uX8VrXQ7KIOhoKrClLg8Hmrv4WYzVjpgY71q9lz7z4DOpV8me7BHJtYRXAoZd
x8LTZ+DxfY/U3nyGdw3vf/cGGKkvBFs97XiNHIzejFkM7kSmFAOoEAmvxDTVKgSlArhRZPjVu/K1
p6q5tOXYl35t9HfpRjpsnIKHpXwanC19TtTjDSk2CbjK46tTbJ0x7NqoU01FXfNc/8Bd6ZbNe3DK
um7KHASRy/fwa7b7rw6m7RQQMXpXBenLI+22keoC7rCF+viZUwm7uqvcBTDT/2ipiGAEt1IuMoUd
td/+DTiyq4ReQ52+XbHaE2G/ntNPvafmABTksl4xkA7OSYwJRRwnV23x76u4MqGAGChsVqKYV0A0
cgRbznH6Ep1mKB3G3FgG/HileMzOq4/2zpnS7IB+HQ8G3g1ovyCX7ca7ep4WXWP2ysMxHuyXDoTt
sPQY5PrsWlrbgNM0MI+bgk1Y6XsFnWw1UugWcTCVpBbQ3Jhv7F9ABYfvBc1sJb0KJhJ9ZWZyyNj+
u3P4cCAzBMdqF8Nk76BYsn6JvmWGH6rVokMOKfw4jsdGmmqhAWAUjlGhQV2YZRp49BDS8l9oOq2Y
gLM3+ZGrL+pAmr5HiU3AdHS3wOylFGdDtAGMdb9W6YmeFVwiixKo87UzxQkH0KxtJ9nYLFnURBch
kbJGyUIoOwHV9+eaJdHeF8izVyuEG85Qh6v1iThv/V8p2h6jXab8ymBgUBfLIckeKG1GaD2wwk3k
UMuXlCyz6OebxDQug9Q9vdP88cBz4VC6HVF05G5EwdY1rhZbA5aIlUL3e035SA86PUwsHge5ORxJ
xJlmL5XVYneX5dPSyb44Iu2GYuWXCU5abCtmdFZbuJ+ZY/v85+DjyKm1a5icxmMO8DTxa14X2Ntf
iX/f1X7xN79XNr8Ktoi+c2E+N/ToJlL41qZA2VhaFdCjjj6TP8ThEmKtVjHrOy9oVxGbudNoYgnX
B8qpPGN/r48NPLeTwz4lDAAaGgVrcqL5Ne00VUFlnaCW6ulau3ihg6mdhVU0KBOpjxFG7nSSkWmP
3AYbJqvQrRcK3OwP/soz0Sm1hpFK/VoWzVpZNbHXZHMI6CJYO0x9QKV3iHQAxpVj/WUFJG1piULt
2K6uarg7bTTCdKoTiZpsVoX8om6XS32aNrh7iu20eE34DT5ppzmKvx+ughqJBolnszPpPE2YM3Ok
XrO+94qmuHE563YfxjPcSZ8ykExuYlBh/uiuDrL0vLh5vSSXGo2BMoueoMT8TzOT4n5dfbitx56D
Zo6BWw83Vn+yAM/p9aqupkzNprWpBikea5n+WxdOyfSEbVARQ8abYrRafXSQHxG5vXnCl+wurg5q
9YnPDv4MNSFCWNzfDHRiFkmK4MnXiA1ruDA2jGPCjxYo7VRukK1kEzaCT/DoTPPDmoyhJr2c1Anr
blHvVUENEJE0nl17gw/zYd2H2YIDQTCGn99o/9j9mOBU/ITUrhSLyjgQGY877qqdcXJPOuY77sX5
u6cmBh7zkI3LIh6leYCDNhRrUkvH4nWvHqGPCTtyDGeuM32l70nqHzKcIMtr6ZCWiy+bBb01cdO0
9gEkPtbYibFvMLC2fyxUyMO/voDMcQe12pTET20OCe9jjTC+MP3zE5fl4IQslw0LcBWAlhPQAX2F
Gxlo5cAVgDr8y5c47uRH4UUJqyeiso8WOFujy55HQaX4W0Hyy/wqax1bDlvrXhJ8rOblcNE4ojvA
9CUzd7sLbeM/1JS2GbcBiFd79ZC2u5u28Dmj0YBzx0i3GBy1jaJBeYXPzhHESfUXbXbWo+V9QGKf
8LB+jch8gmJcOVaoK6JXgGPugkLPaqzp8wFnVx0/K3msJl+HkAfJwi1qx3fWGTf7cZE0DKSjN3VW
9iO2r6rpk2xbrtcn1Lx9VRasxgjnm4Y3LRugKXJX0d92Iu+BQm9zpPW7EhBrIeYqVKmeBFHgWBLo
5SD7QDwOM5S5VlJ2owQZSNmluq/QR5CzWZ9uMC0Fsn32MWJ89JiHJG2dWZlgDjev4OGabHW3c1gE
Gqecq41ocS3NEeOB/c7BLIlTQf/Kvyr1y+C/dzR8JG54962FNAfEKYr8AQ31vn9WSFnv6HS/gcVn
g1Lck86z7OYVUds+NVHwP47+kZQlIXMG/aVZS1LIknB001bB9LV8u6SDqAv0EVDPslJ9ksALbkBG
Ym6ue6GpZGXfNZKCXjvpq90b9UCmvOg1QQtPbHpYPrKQnHFdTRm+u+eiSks/eO0oqv9H6CkutooF
goOL+9DA78kAtx6Jymz/+mhkkmCEA2tME2RKn4vDthyUdE0JQQ22BZbYiUaoqUGFgdNsvDt0BTqH
GA8ymQqj0fGdpDeBNumg4ybpeSnnM8E9Wik6nnAXyY7YAlMgPA5hBaVGYC9aRcUNLlI7XZpSXUve
+ur0o9TNPh/5Dh/J6CF3MjHYt+Mt9NULunQs8fwPLc7gedq+tvv31RiQfefjJU/XWM3/YdfypWgD
fICauKNWSvMmQX51eN/TWcJa/sObr1zOC6qkNqvrtyM4W1OxJvsqOKm7o175ZlnkxYY9oOdKFE+C
Q7YEnFBZwGldoCz14yEjaBOnF9fE036+GqUTeGGPjkbhKGIJuxfwJkM8OYlzEM4zblDpWGIMHXAo
f5h+Xq7eMioafSYsebxkMhhd5pEo4FGqLijL4bIkc3hqN68P/O/Ub3wXqjCNxwlMrKLEgYTmO/9t
4A1KmtTo6ZYUVCHomQMSTpZgii/S7b+3UJENut9y21CpVA/wVbnTjvM7qq4g567oW+9WN5oOLhQs
chh/CxSRcYPJn7jtAqinHkJ/eHEskjjFsI9JD8mNNMaWIZJZVE8ClNHCszFIzLv1H0Mgj9pgHXcm
iNZqM3KBvTYJs+Sv6VepHn+rChLRnBXFNUIFljvFpM631D6Xzj69G6X+gkxo3yOfPyAEYPrmNayL
v7sCHsU6PzOJhuOt4Yv7PA1vTjMbGpeDPMThpcp7H+8La7CyO1/I35N0/ls2Sql2ng5iQz6sY6VG
RhKw/ekn0IUxcArH/VSVeJvhBpLR36PqJoobcynO5q+YOeuG3cYMbMGDlou54EVS3S5eS4ivRk16
ikS+CfiF3jpM1zq6CUs8DE39UO2P9acPhF5Jmcx4nulGMzf8u2dtpfA1uLEMkwwdXR/DhfcuwEB1
bqvn0xjJZNPQgwlFFUAWgA3lNFdv+TsWmRruIT7CW+AfeyHLUYTZWtHlAOHESZkqLX3QjAsl09xD
mhojNfJshajNoxVCO7nmz1/e2aaqLv4HjB9LOEW9HKGbhE/kOjK0JI257tTYV+uR5cIO444b2/vo
ZU6h3riBTBNRQuFItG+4qIKzorQIg8kLBQm6ZwTCYsTy4W9vVerxhz87af6mDhR2LNbfrAlzlzID
f2+3aF047OS+g6K+68w6OaRx7roGYhSpDEElavLN7Uc2KpbqG1+Y5C+YK8bWaNrs2DsYYbNYe7E+
rw/dC+xul23KjH8MISlhZ8c1by6pmSGfBD1oXZsIAGTUlfaSOEKP03/tYi15n/TWNp9gWiXasspO
D0BWtU9TU7ZlvwC5fEPY08IkEgsLzLw6LoFYCkjQ2FZolgZG+5ErlGiz2BiKCwgnvNxJLmaV55oI
jVSbOuUEbSugs/Pf9y6ZdCPKoYQHoAaCdJdUOxV/fr4TV5m+JOnqIG2b5cIDhCCtvLoZYP4iQvLt
pZCMTBzxGrvcJW8SCzP69q0sHF0tNZbVRQZN0k83W3ARRMmANj+kR/0xgXb/+7Ar6mB+XQRNAuzp
3SW1PZ2RG03TiLVYuRhE7QXLdFgy1UXYcm31RBx305/8liYSFivntMSXkfvZC6FppoyV27Ozd3qG
yTxGNQAoI6Ap4YvmdUd5f3Ms8Kzj4gE6grpq4+XqVIzj53YBLfYY+LY+dtA+oe8tDNgYAXKgCbJK
2TlJkErv7DJpsqjhop/PgwniVe4dBpe7dA7/CTlXnyezlbXciPBuNrEwAI9hPR6A6WHdj3rDKEWF
XYdD0bPCFrffRHZGRp/JWQ19szIkXyCss17pMVB1gN3cIxRjxciJKhW3xjukCyAYAM/JRnvHWsGl
FdxOPk13toCoSpCZj7XRfhT/Adv4V1j6Y8emmb9LQsIDnYEm/fWJdse8n8eXnLpwV6bhY3ewnWA9
PmtUyQsArVfV+GtrJUqhRimk634N49flUSNsTFqsoANSQkPyAWQPnBtkyiMSNMq3fXZBBRw/U5IG
/ev+40yfrS7KEkxi5wNJ6bATt/I7ddsDgI74Tb6qO3LFlcf67dKJNM6wRBECH/J5CuG09aTaMPRY
B5k0VObQEt/w2Z/+XqmCAz5Sikm+Oqw9SsqJ++2EHF6XKVE97cR6WY+Xeh1ME3fc3zCUGCU531YS
K84Mb8KH0GMCIF+lZisUR9NsumMfG/6ZVh8yw7eG1zdnetq6kX7djSjwxwXdMZIWt+ytKzpnFSSR
2iKF33rvxsyCDoWF9WwihJIRdWBpNBefXSBItNY/dpbLvoFaz195srM0Nh4VRf+yyHnCUxgWeR3a
MPZad48FhPy0CpcdHimD2clQDQ99gP/mhhC6LK+69vWs6oT+lyIt7H4KJggmQDoiwyoTw+ELhAki
4Ungb3cQZwdqwCKQcTeu7aP8dsvaJEdPt9Kk4cddfTrilaXC7bd4v0C1ovEvphjT1QtlwCZbrs6D
265DATid/I29DBuFAek4A8/6j9UgOfy1yCmyniL6YcYfDljEehgYAeCecJsywFZq6kq6hg4mrWPe
0Bc1kd/Rn2s9AgxzGW570pNtLI/j4+Z7yekgJYM2r4taV0OT5+QmOLGsWCjrCYoZcIjCf0hRZX1G
mFiRrvVMF4o7cptdYJEB4nHQPYsjcBIzt9l/hhhm8EEyU1kwDAGgKUFDoGAjgHRGcVKkGKVVAjkg
DoveNNW2oRok859jAL+kz5wcX2tnQeIBhmOQXdCuFCQpYEjSBXBiXAQ3VbVSBpnUreiC9xtJ60Va
SjcH4yi1D8t46xpDyUjUl5xs3sEkbU1wTBxdcPisk2vZ6BB3XkvzEb8OH6cTHLPmF6Vdx3BtnfSe
+B4OpvCG4i9vNEP9rTfa1L1wnhmGQ3Pjb7P8O412G8swfm7LY4VIxPW7SGfnE+Ie69bS2gkLZvUk
IhFrZHsm17/bnnrosDQBSZaTv2FnOJj6RufJkaK8jybekmIFwB9jXEl3cN0NBopIsms3BpfCqZAu
wMoVoAxEQVSdvWJ98mqJzRZ60WO3tXgyyb1H+FWFj17SEhco3rO6Y7m66cgN0LfGFxg0mpzsXXcn
q99ZYGdofOZ59HZ2OlegyT5CQglfG/cl4j9Yl/QJGJ/7dJvcnjtZ2NxURDdrxAPbesLn6bAA5B0T
Bob6BmZJwwEj/ZJwfenF7nq9sfup9PIcpYcqI56oE2CWYT19Pfjp33j6MJBF4OnWCM3TKhpMGcxG
hjeDcEq88lH6rT9TW8S5zCnUSDTR3MdGMxsAi25RVOBK7FhRrnf+hrgaZtXBwn+FTe6MvveXfErv
g9frwW7tSL8B5gAb7KNob4vM2fU+3qlFpixmV+A/HPDcFKwWao216knwHfNeP/rhkez89j2MySTr
ZVx7jU5h+ncE8GJUVrx+vLCSWTunfLyUSLlPcJwtCBiAj8lmMdzGzbZMWio5X7NoDWVNLFC5eAGq
D3M38ILjYAwMGzLh89ZO8pKCTV4IZsdwQAvCtpz4m1rCkJ+uBUGWg/eh/8mrkXGr5WR3GNIOpYz9
F36RTDCFP9Bdfe5aPghR0eMLD8ytawGG1m9w4GLMID6EgGLRWH5RFsMuERpWZXTWV/e0ua/ZPV29
rhtkFIf7J8HrQ3vfPKBiXqc8H1U8/MYZxA1iYII+JlgWNQD/aVqs7aBlt+B7tVHGAeF1mfIQVhGP
xKuVei9GjJoLgPLFsEOXnbOeTs4IK6/bf+xkwbASU7eSk7nqe3Iqhw1aDHvIaryKO+VQ+cKM+nqb
CAe/l8EGms0k3vdRROGcCbXaM7SzZYqX4UIQUB5u+990VvNMnVM+KjFWFMcZxwEFfLhnHa70DP0g
9W9kVCpZQ//P8fnqG+dDtBl40oRTRTKAElaHkgApwqNl1vJIO3Yb5fpiuq5Sl53SH4JeyqUdGDKT
R6y2ADsrUtHxA611l4sPhYPFHRyhcB/wzrPCe3hT/SHcccjaupiFHKbEHvjlxHTQiJvzBu/h+CRH
zv/gMimOQzI3seL5gyzGv7eFuLLxgsfJVDFq6BdEDYXrD6vd19eaQebLvqEf1F5RVdNzF+Putyri
C3SHBe1IiFgcrb27zbmebxgbVYxfTERzgSgRcCFdnLtc5vs9GMALBMDz0Unao/g6JM3v5pcmfT9a
QViCsqm2zGNf5RVJoYGFvbTE6ubNOgJ7zqW1REfBCY8jhqfEsYfB3+Oq7Uc8gbC2J2vymd3Wm5sg
8cw6aHRCyxOXah5oGTeocm56yzDtqsBOMCtUgC9c5xUqPe9e0rmZzealzddKv1J2cjQb+lwCrFGW
Zi495WXtOTEVT4ocpsF1inHCDDWXPAb44Ty/EeBW1myVH+cVobBDkdV0QLTuwObigjl+ddcSYXZo
RAl0jIs+n+Z/tRwu/NC9y9dOVhRXYcC0EyBZoRVwuPv8zqQUXn5F+LXD2FSBNdC+HMJubOWY4SYA
PH/aXf1ipHn7XTVcnqupm7MDx8qMA4nGBComO63OciP5HQ7PacmBHrZV5E9EVL82GUJF29wHOIfW
86JImgiyk/RIB8AL7RhXqmhpRi7egtEgrGwkq3ZgTlPBPlQwXEvuPdlTn9LS6hvtowkkSEH2aCi1
ewA6nOptcnmQF0DqDXolK0aw8eUQt2xdiVGI2MNgeLeTlqlY7C/YibpdFF375xvQxQMedp/PPjrE
x2OzxnM/vLYRsZmQkUqpgIK4moO4ZBKNWFbi2FTvkUY1LnmMjWkQoPiltZfONU8znKFeiGZMCmHy
Nhu+hPmsASi80zwjLUVezNP+LRdroUPbL6RFSc6Jiz8owIbw8gfGMF78Qe9n2gPt9ZLOYeDePEjV
JdEh3gbT4Gzhm6FBT9g/IO8IHzweakS7FH2RfaoD58gI/CEYypaQQj75J8+DPN29fnfmGyvT8atf
sNIWa2yleAvKVPN0kMTkxVfYWgd0StIHxa/4qFEFMG7KPSIAP8R8jMSpxbgKwIlcnwR80QrEBjjO
ffgnrBu2mhOhvnw6EZQIXLfc4eeM/7CKPNZ5RHB/q/glmgCJTBaY6qX6yuHGHV6GjrATrQfmah3o
3LXsrnUjq8x0tSmZ9+IAQlqzcPBXQhM10wDFocrQFnud51zwh8MVfHHIg4SjavRtzbnoVmdpcq1h
wCsG4ZRypWtu18FLxKPFwQoH1Ncn+/uFdWqzNSOvgCswOCGvXHD+Ac/1XMThzagnXhcvPAP7bq9C
KJ2B9b4ubg5Iw+cQVMoZUk+nWNsa1KwVm2KAOP6Mc0DTntZ5KeZQ9yGaSigZxIKVV65S6BidU/jt
5WI7MOHjWTLj5p+yh86oWjnRzAypCaWlWxuz32L4SqnsKMzenfo+pBD/riGdokOpLE9CY9ljWopL
EtKUT17TsZ3uUfX9U53qMd+NgBAo8uxHJMLEkaNaVPCPQ0UHaCSa9ompaxdrVmDuY2MkYoiCbEvl
g/+K+xsZwcwSU3SG95T6PrNAAI1lEyUq1R8k8g59aOr0++vZ/+gJe92U9qLji8ebNr5zauJn0d0F
CN4UqBpcn3f1YYdWrZ0B1rVIEoHxEBueMo2iHtq4Z8gdnk71bRRuhlhd9BloQSvtES2JO/punsJy
gNDt7NdNzm5FL2Z3I3OnSYX/4F/NF1MkCe3jfqpegWBQ2kaMDh0ta05ChNafBZxmkIfiNFhlxkNe
lel9b161iego0IfLZgD1uxkw5RYxzNl+7huAnQMEQt3/1pNznuKSWlprMOkNKW/X4lUWwihCTq0g
LkrHVMghp/0qgsK5FYpgffl2aGQ3gvqwhbTTfnZELzcbLCR2dljW6Z1+WDOM1jqPKRkzQAtJedjN
Il9WYEbhf2MZOF3oAh4sgAYUHiND3JYTVhcThyw5s0ggUmBrpiLN8xjHwhmLLsVaB6dJWb0mnC0c
C9hUAuuIS5K3orDO4OEg5Je8d8lY+odFuvQqfvoGFkrIiNVKxPm9zt+YjWhQOb1ooaVVnS9Y8azM
eD0OUsGBX80jJkOLBZ0plPWDRuQ2Sw2djXxB7JC6kPY2AMWpq2UiXjAJS+K38YljuEv/5NeA+LK9
HN6VF60IpbRyEDtDue5BHOmg/p9RFaSFhxvF/hqwlFMmfh9jo68qS1XI79rQHdJ1847jLTLy/jZp
BeGfsuNWoxxd+XHbQlJgKHZIVcY9Xfu0DpcMwxQM9IlSCuhS3CXVKZ6SRCCW+aozByVloesTfejO
YkgCMFhXn8jBoYfFXfE8pDW8bd09tXpk01qRCUq0k/urZWn2SD8WnJshb7+DGWcDN3RYAEtxpkk+
6DJdNJGdzPc5U22bfWoTrhR8egcljsTYt8iNEjJU1/Qb8lOr7X2uj63HJg58gYW7/24fa6nxYs4D
3Knsma62p+JZ24oWSBvTVJLwoMuL72+mrf6EhmjYHlKUmRWSOUdUKmr8qeBPmdPzTMddN306d2QU
HcCE45sZNWTs8sx+Y1wSkUIcfQvmSUtpsewI99GepDl2uKZvGwsm0BaxaHYTijFYbe/IBgKBD9Aa
Lzd5Bmu1tatjEQO+BQe3i8QiGQb9ipDCtzx0ljl8e7V1H3Cl1pde2zxj2B30wVjN3Q7CThIVSnJc
Ot2fhq+7CjMGQmbjtTqPc9hgdIMQWjayEBbfwCNyvIbzMqYPaKCZiSrwFlZjX2SHQytCala54Yct
5S7pXKNWJAyHyk1hRbHBSmvPvGKDILrl8eQgkNGnTlT/FpVCSC/OOE9czdhLnsQmT3qTMPekZyG0
ITQ9z8b2qK+Eu8UtP9uu7R7nIcClo8XJBayWhs4B19aBHyKkmeO/qr0QPJTQVz+NUij1xebAxBuh
q5/iQ8W0/flgv5Wbrs4qjUmq2F+GgKQstluOHUEPu1VldQI4x1RfVLwffLXGnGogOFZJ9M9ZEOKt
kiHEVbPGnERjbASsGBQ0JTVIRPHVrrc7+eAjihpq57PGRh/SswAzyH362Y995AuiO6PBb504UYiB
gvfdsxlTiEfTCrcQcu6NAAYmkhINPrEkka7CKYeOeOBC+Z28sBlQwVuQa0Gl5hB8Ff85/FqAh31i
BCrSAR8f+5s6mlO02cPiJ7teQQOif8EJz8/tboihffd05Nrm+IPBMQ2qAn5rs1ICpTaYt9q+85GC
q07ocLeR2k9N9xqIKr5Le2HCW9t6dSUABErq/kQOluozWHZfCWH7j633x3zNJEz0obge+vUodAUw
7qNcSWE0LY1ilgdTrwwu/Tov2CMyw7k+t6REMAy9ZbNWcu3ipKhY2u1NqqkfZW05pcRIvMRjYkm8
0Eq+Z4EjS24WVNp16r84FAyHXnU5sJz65JjwtxAVNH9/8hownza4A6zlNXeZQQ0Nki3ALelPC0Iz
7mmHMWx8UKFwhM6/R4QzSVHkX/bBe4TAu+zLruT+LytWRMenCj2JdGxqDcMboeKy5c1X9fzLdJya
NgV/zV0DVGx3UO0V9oyW6g0q6FAH9KlokLs//9AnAJD2C668S3umfTrGHqfPg3tlnrDTE53rSjgz
4yt/8GRpCiiToQA0OPT2nTPbABruGNhEXWshpKtMNG/Th9OiTjuHOQBxYfPKUJ0fXKDHdNXGRNrA
ZjeNzq6d2WTm2iaug0kjtFvSKNULM2PZqYeeQKfDdtMQMURx3likj1Tsh8xmnBCOpnCCg0tjTZFx
i8Tfv20Yxl5mBaQtvGtghp0z5FAGE4wtzdJY3q5f4qtxDeJRUfRAYxC9V7FZWOw5y3LXBsmgoOSn
1v5geJMjIgu/rD9zsx0wkg7LYe0ZAywjdm0hmEY1xqWAZXWjg0rrr8EY0MnsB4Z42lSE4R1XYXHN
kj3YX1HHH/e7CEN/gRt201GXvFW0Lve3MZoRwIMmVIEhPGTZygZJM+a8S4mH0xCAiBZFYy7jMegG
pjA45V62rndQ9E2/vHXviLFUT70Up8bAdkOXFO267VoEtgVOkyQVex/jj2HI2U5msj8KtnATchVN
6dOwQdobU7QxTKz09j2Aj8MXue6BNNgMafTAeLmSjvdT1RDM6ccTKwByEJUe8r32fXesEoDf6C4y
nrBz/O+ZNt62TPYJJx8nNVkrY79FWs1i/x0tRf99FLT/s2sd/9ZYAuvfYPu1cdVTCE00fCiiyZDB
IIH45hr219jN7jM8QGcZA634Q90kaaFWNh672adleHuJoY0lnVYhNhwgHWahikwbQWGVPXxIgTAR
tpBIMyD/WPQ+KkclPh26QaPLh8pXhVbMgKM6manv1eFDC4kELDCNXUO0wJpzO9gt6+WcQ4OMvqvY
FmEbKWIWMUPSuatcxfaUNBDTdYr7Kt3trWnOPUMwY/sdo5EOcGqvufMuQBZhkBRgEE/8rjTds8NV
dIkr7oDeHZzvjfPknYebYSnAUUcEt8fD6mArLpRG3zDYdEILtjnOFKZ66oxbg7pCtCyTlWhmrfF9
PhXb+/VxhHtqh8Ja062/LKtl1TsktZ8A+BSCE5E3kNI8GGb4YTlEdYi4gTYWBJHQ0iM182RBsbEv
DdcebqCItlv6+yNUNcz6xfvlcuTlOYfSgmKlxQJx6eX4C+BEK+kJtx/jlG0HJP9umZ/1CBeRi4KI
sF4yFnRYVGgzgbTxTnp3xiGUX8dnfkQ6xFhc3Y+MpvLwS2GV76GZ6vmcRxJp9ox/n5Jw7ywPQz+j
235loChHV79YbUfdJkY6gxCorj4H6OTxdnNq1oQ/L+TZx0yJZb06TVTIuzKbL/oCAV8H/ArD97k+
MB3QyifBJdqxRf1hoX2UTMcwLtaqSoj5HgngUo5ZLLjslFiLdKs0hbpAwIb9XulcZsc2EruzPK2D
6VIoAMlNn7D/B5yxTREQp2Ckq2LkDukv7w8MO4/iaHibd7MDOXbyn5eRDYyKfzvsGAVQ28xh8bAf
ytbSmJLQxOTGOAoGew3Nk7tyKltLt5+R9iBRQeBCPsxNf9k+yLyByvSqxZ5I3laGKJjT/yhJxWxJ
kvOdcmRzl1up1Euxn0j81SzwPesKI/BIDZvWl4HzJ0ru37EusScMsVS2pUv8/jiUASQsF89X+Cm8
aRh5vQ9MymgtP1q4bC7XdsjLYJbYTrzmaJCVaEGeCWiRPoP3UWkCZSqhJuU4H3fzM1e5hJX8gAgS
x8XnakKOxybgmP1g2UqcYamDdJHHftK1Tw0X4InKlHzubqrAOC9c6PfPp3jPjeAoKsgG/AzYsOG2
1D2NErY2z10Ozr7TW0H6WD0sOzclks+2Pu2wi02M5ArUgJOyiR7skIw834C2iYMpuWueBQhDce6f
Yepbi1Ci3ajz5FFkwc7wpt+FNtZQV6uJsRGI200tNP2oo7dG/dkEvLn0ido7MP5bKDPbq8H0G6EJ
3oBZzkrFfGHkC5+W8axpMc2dJhqNcXXhKPphDcKm2cu6xtLj+oI8ZedWcWW2fM1M4f5YZioOr9sn
DjtZq1+VY1yybKowr4WUC3b8Jfx4hae/sQlCaoFas8bXZdGYUkCTYm1WWJZUe44WTmlWJZUGF3aj
LKPP2kqIYOJuv7/xUPLHvW19sI2rw3TTHWDhk5HUH3ciZB0cvW+DET8n0pFzyfbPVYzwbsoQlzQO
Q3MQ7UM/cG8gPeX6DmR18hZRc3hLMoKCL5hNQ/esNsYE1wBwLd3k3XXrQ23yHjkO9LO0SrM3e6q0
UaRKMnQ3VA0R7D7dOuQwU4Mv/mM5RJ2rEuyiNQoFPmOCTKgxaszaFgh5fgnJWTTgYFbpn7HZtwdO
1xAoJnZe6DmyNuDTnWFXPU3jz6n93pPqMUawF+/Yu8J3R4hx46lpLw9Mv9JJD4/Z2A4L9pD8ZiBR
UUX0hD0F3EHvuIsTNhOjSLXAEy/ZLLKFHDz43fIof8vhkqYvRlY8v3x3jOu6hqsUYZTofiqNRyfK
AUZPtSC0sEBwsKJDRJmh+bjO+KJg0nocJ9RwyFYPB2GDG3G8r41Quv1nbFflVsDdlg2CtI2TimR4
W4x74rc2kmalB2QrsU0PiZj7fnR6+V/GK0Yoh9nUUoBavavHx/bbwK+rfCnlUl7T1YLX7jeFU3kx
mtH+2c/EsdHcQXvHXUSwVjTSueeYSrKgVO+nnCrUXoLtKs05bzghCL9S7bLkJTnfDpMnGMLrku3q
pzJr8cSnTxH1ry31+skXVZP2/PjZ8IA5+jF44kCkgPVwVovde3aKajbrZP0bU6/GaeDR6B8FSUQ9
mhoxmV8unuiVn2WRsgM7C7AQZy3Jydokidox/dnQAJ1UdQDQr2Sj/iIi24sfsHyFIYWpTPi/6bzC
0pV7Ouq5geZjc3udxdnWqXXd4nnAFj9jNoqHN0Zll+U9R8JvXjJel8H3oW/nzZFy8USrZTEfD6JJ
xa7JmlEJh1J+QdY2hLvmyHAIJM1CjHcjhvX46kV/ihfJtwExzfh5jjxbJgbr2IPGc8cC0JNeMqaX
aIPJPDnSIlO4mdCz6yGTXB0uJWxkMX58voyq5qaHCiCcCJ9TZmR8eMGIeQMjakZuSj7r1UWqJZ6N
v4qKr0ldjRHch0hXpUDLefUUCyy1y9MEhfXa9SsdaUsSlhiZlHipA9/YngL4WG8Eur4QQVVGgz98
cGCUFdrwPv/kf10ZH9kanwqk2LPlEDW1T6iGF9EmbevPQyqxKiyFwRcSdAzkdz+J5/seEQja+yO7
k+GD+LPEQySAkAdSXQy9waxYMRsj0YaB5AVJ4Hs4knFAKivlBxfMJP2TmRkGxTo3nzDBIS6ymCRY
0C2vHaiUIErQiKnmit+Vz/CHCSLy2sdsg2wmFvY4rA9cFyWzVtjm+/Ywrp8HDJ+Xh4DR9WEe4jyD
kEvb1w6qmfJXHagfR+prsRz4Xtw0Vq0+I/eiiHWddhionyv4zmOODW7gXVQeV8LVmlqT4R4b8XB/
muqt2n5uUg4o/dFXukabFTwyDBiGt0Ipn9Q6ae7MWWls46xajP9HVp8dFoNsiHYP6P0jPQIztcxK
DsZexPMKYasSnrnhVsZliq8MBc/TQmLA36MDVBWYTmLYxmtPH//XPl47/z8iu3WO5JggkZ2Bz6Jn
Lym5g5BUhEDizdKmap9PUrHnHrmlb45DWDcgMnjuYpARZQT0uy42jEDMX6vmf6nEQdQN7FmivIA7
tD4HmLmDTmEEWbFIR/Xw+60D3u11Bc6JCftikky3xEBx6D0/4JGKNs9rTNqeiWyzwjypYlfkJSLY
95v38vEvvaRurGfHYQMIJHhO4eKsJRKmPqjbXrwxWnDB/ETaIKkftxuXMsaMF/5D727qGqs2jb3E
fljllJ3Apr1tFnw4Hr7C4Q0tkpn4z2ir/1HnLoCYH5EF6h4PS/UGFqAbA6nWEGiTfAjuWA7aNgOT
0dT/zGvUvO9Qaa1OxvlBCtTnRbuQgKq820xU6qWEftRTdl5BZxTwvKyTo6wh0PsN8yC72xs5O7IV
daGi2h1kT6uNAn/DWLFqJAIvldp74fFV1mqkIsHw/3leWrDq3EePFHDuyJaQ9WUHBA2AZS2TREth
9Dpa2PapjYYb01H5KnmLP9ty6Zu2OzJWppzMkXAwfK/dlePyWJpbNqT4KAph8cyk6xd8M3E1tB+R
WJ7Okwy7mwEMotNgIV5G4LFpolDQ8shMw8nS9+T4CDS9Q2MNXcv2NMJxkLAaaXtBk4lQXXFSULyY
jae9/7q4Mh6Cmzt8TmBj6NeJuS+sjKtTbJ6eq/dXnzqNW7Z7O4aUjdTP4Em9FQTDaHq+7NpqXkR7
OGsIi+QlBKke3ppgZ9Nj528klxJhuUclWLS9I9+o+2vwWcWiBnXACso+GPZpiU2qrultigmsB6PT
hz187+oEUSv82fvdMU8Hx1lvnB69pN7xNbzalQUpkv2IddHiQf8TupmY6IJyQRWxI2Akxfgp4r2m
VhP5ghJvwSczxBSupy8/G4yfjXX0XxE9zVDHaRxd0K751TPZcOc23UM9+hJzgwdmkidXrIy0pauX
YycTtAMjlcMz7GjMS7FdH0/004QTPNbr+iU4H6xSMiDzg9vpa4qk6LfGNJEb6P3TwBTc/OFRk24Q
rx9cSncN9Rg0kXR9Rct2cmlBQ88V/DMkn+9MubISbjeIlnsQGMkG36tkGDZzlaR7oIA7W/zzoswI
gRc51InOwzHBMUyaVVe1XegPHMHnrZFfr0MOerWaiCMd0hL0VCvWDWlsamY6x2KY/NsVlSQG7LKU
nYOOPtctoD2iwIIxY9RRLpz+MUIwy3DAIvPPKhd4xaUVz6WH5rDITlTs4T7xBhoQbiYuK+LhDR+n
+s7MJwqxHaQYASXO0MRdKoArAlfsgbd3zeMHBJi+Hr2lFiIAVHAV4pufwShp5BA9d4nbVjagLKpr
J1AmF1wJclyp8iTcjSzpsU614gmIdLSLlx1gM3LgL1S0x7JLuQ2rBntgS0yiL9F5Ik6tiWmwZ0o7
F0Mk/B0nmLydK/mwoLAlSVJ/YmiE8HcX/06zvNxIbHABSx3GGxkXL8l0gjFO+u1tHGzuNxZxb2K0
NjHVvhNesMrHvomaRI+FXWms8cy12cLZM2lh7+bUWmYZwxtNRZhnpnUgaWZPZCZ9AImXRzkpAI7/
EapD8fGZP+MHSWNEBdx2OvcOG1MOldfDA0CjpnMryjYlm75nPKOJ5akaHIrK16lpJJRXy+wfBtVP
ESinpYqLxo+tYB8qDFHIr25aSJJqYgcfU0R+fpzWFjeqV8BCM9tOf/TmDexy1Q7XIj9DuU3Nrh1z
hvEmGh5rEYbIFt90UB8S5JpOb2KjxnVskDyK3+XeIx9N9yKYfnYIE8JEPsLnPyhjKrQ0LeNPljqH
LIn1xEsdIOxEm1frFPBSoLy6u1th7/SM0wpN29u+wYFwGe3AFlBg8iWt9SspqpfQBKqC74DyXxgr
EPHXzY8NyOXhpFPzHL0IaLN8zox9cY5pR3Cirzc5YUuBv1krpfkjoCyhU3B5Nf6Ct36CIj8l59W4
kqP+6BMRwSDn/Pw5W47N1x0D7Dd3fWOmgX3M2P2L+N1yJiAD6QmplV/m9H2MYlPjJHsSHTqMglRe
FPwcceVcYY6lqpJPTHR0HUSCntjWSpcU39v+1OE+KIpj4+sB39rES9lP4GIlXBk79QuDFwA6dzhN
xNUZTMHjg2vYVuOGRBcnF3YjhR2IO5Er+z/XzqdnaoYpJ46KDMx+1vPvOIv7ZQ/okYkESIumbSXp
Xe7WlGT3omJ3PkskYDm3v3+UuqFJeKQdaoKnoxbZoW/IhHs6pCrc1eLK5cGZy1oGWEMiTdvXTnJ4
vIFT98CBZ9qWx1KIkN2WaxC8kY1YUbT6kNd2o8kTuZwqRQYAAYIh0TYPk6jkg7mQM5QF4ICeMVoQ
fNuRCLW08Q2tiisO07bHID4qwK7F/R1vkIlP3+BlkMZ2d7xBKpoNkkDlNyTrM/+4LecG/GqDqogJ
VECUmITwELlA9DFGlTon3591fIWnEkWEeF2jjFiXj4PBlZ5wvDpC9sGi2HUJzbXkk45cszCwPpUv
+MU/wVlle5KPz2RfhnG5aUdgjgA3pUWSO9OdZarVqxsLfIRt5YpGU5tFe47DA3aBOQyCDlzlAvZQ
ryCLqj5psmzO9514ifm+9pfZBi5bV6KO3+T7GOWiNqfaGQl1xBWOgRptg/ftu/JBhNLyq5E5EPqS
4nxNdVMMGIW8+y8xUXDydmOFghQvmaYgU0UGb31H698t2DitzD1U21TX85MJTAsZiAeTtMQO+T/q
jNJ2Kvc8g8uzj1ZxrSiyA9rhHOIJA3qgi5+O8V9fjl6mj8uNsCIsBKq761sKFnHF3bxHnhgO5JAq
M9xn/7zv+JoOa0a5R86EyuO6w6EBqRfqUqAbh3mW45r+AlrY7ZxwhIXRNGkDD6wyDNagex2ay9Ol
LoHx7/gPImiy+efyNG7283psh7bT6nHaHzuEZCZBqhn/SKOd+EZ+c2vZd8gDKpMu/BnOf2Z2C0Bd
v+9rVVa0buuY/vSAjv5m9sUtQCbCAXFXR5vwHL86gIyFeCyKAiIcWu0bCqlPdqNJRRxsMInu4YtR
vP/CeW9v3JUO7dzLgi9OL4HFYVZpHjeS21WurmeVnw4goQ9EvuPI79uXyNv+PwDykczruQXg46dK
TMieZMqhU3uCmc6o5PuirnJnaO9KDPBYshlJPD30O70r3w6ZIUui4lExU1UA/8KEFXQGEu5GW7Dg
AwyZuCdmGPsUbxOfdqYnE42vA+UhXKKxzDNNiy6s/Yl4GTTO9wM2WQs0k4Sb/kHEmBrXoOQVL7FL
XHTw3r26RPBuQArTZEi8OMyq9sAvj4Xr48si5DhXNGgY+VM0QVwVmKi/rgjlSESsSBLuJR+8IAhz
YjHKtr/TX5b7OZCXmy2uqi+Ns0Y7PB4FpncnUmef1d/v2SKwBW8+1bFRh93TG3zO0J9ypSeco9t3
b8VpKz+dONZlQ2QRONbOV3ndhX2e8+uRB8jFoCFgypXJD2tw25dS7c/Jm5AYW2YVpIdwxf6FNu7f
Z+LP6eRPxvFeJEYkQHIKVGhN77z1oaLDowt3KmmP0ys5OIPYxXhDojtFg3DU6Ki+CG6jwc1vodWw
K5zM+P3jJ9NtOsYoM1tz1wA0b/Gr9jZEzv2Phk0sWu3p5KI0ueqU1NnV7fx0VkV5STOqDkXgbvtm
U5AT3SFvJlakcYPDl/hlCcUxtMMSqr/HYbgKnQ2x/Ytdx/zTYywxjLbtZSjhQ6bQnZDaZnj+R0+z
8SWpmBFlkbeRc/YmqPSLbd//Bu4rK/2uJviIHUoiX2jJ2+/rN5MN+KQjogc1zvL4XVnTmcVyAdkI
O/WEd0NOPxOBMJxgT5EHceDGng7FNWRSYf8c20VNBLVYjYqleszHxWLdS7uKkY5nr4JkQkAdW834
b+p1Xnhja6cbS9JOiKtjwHIN9ZjLe8+Uuw4DfQP9UN8FUIbZkh7RMcZbIu7L8vKve3lK0QaPkYis
faNepIF39cJ5Emki0WhV3COYn4AwGOjj9d29gtY2RJ0SzPCQyTZtRF2f5Jp51Cku08Ewvj5QAwXU
IV3nEvcMg8F4FjGkqPepegchWsZXBZxcyC5nLXLpREHEYUVEFnk7Apk2JC23Q7ld3E+xfiO4jAlF
66AtdDyJpE7NyADlG5daCOzfXRDFdMt1FDCfKHzafohSg0Xmrn+Nme2Xa+Gcv0RR/PKgCDueSsw2
/J8jpevrBKssy0gXlfOkCsrstEMZTzYu1QE4FP+nQHUrBnsDMYLVmep0Kb8O2WW6hRdHIEh9TKsg
esfVHndB3QyfCdrCHqD9iMHRrQ5CMu9rxT36D1dWnmehgyCsGOd5Y2Wc5fU6g3uMAV1OGTIE04z5
O9o6YhRaeLhBQayL9ZM70g50KgHOcjeVo5neEfaN75n1UF4ZiD2jt+0+b/AxSlszDbor8JZRgmSd
uPU4xoxPaj7zjxSZkWIdHWTMPncyPdXXw6VhPx2jI8MKLMVekurNcDy6eC210Cr8ke3DCw9Dc+6k
WarJCEBkCFJedJ23NK2ZVoRChlxJxmOQ6/rvA5sihu/vl6/tOE2rwq2zLwSbcRQqfQq8iCIGjcMq
eaI3KVulKmBnO6HaJJB1aGnvT7+hHNmeEhStI+PFlcHHIRaVwAotG219XJMcaeFYAXCVTO9LW1Dt
zM3WdcS1QzmWY7K93n/kCbEg4teW2bqe6IDmokw+mkSUxMNYk0eREG7jKFi/ljNEUy+nzGBM3H7g
yBQ8Ai3RxDm1FhN1C5jxnAgishq68ciCSj36EldZzPjDPTMBhcIMR1MGpzhMjLwN3WO3Jaj/3IuO
W7oWYyFCOQrwJi4peIACNwodYnGqwaU8y3jt/qnWypde69xFCXenXsRqieOIpd4gKuViNWm7f5pG
MrbjL+/ahXQ0aYBVwT3V7FSaVbNntOWAC1py5P9TbM5a6j3YOjOA3on9Qt/azmk5XeAY8Q1FZHTy
Npx03piC91RSOVENx3AqJ7EFq+Soeph0Xq0kFJHvFjswbBH2izSITU0ZsUNg/XgEbrvr2lrpZ9T1
mwn71i7jYll8GdXAWTC6hRIB2kbrcp08fz43MsTGO6diRRyDxyi4lW9IcTdHttwPiuIulfbHcHLU
igOqv3GVSesQeYg0JbI1VHKpRfw6gRFug+AYgB5XP1/1RjTMWvyz/wx3GjIP0C65TSVCMC5do4+W
ctbdElOMWWpdlgBDxg2AET3onf5X5YJZHeTwq6wv3TisQOO10UDQEVOXrSSKl4BpP2DgEcfg92d/
jjb2gUY/eS6CX9W9/MMOas3STxXdcfkccaT/l2GzqF+3lRkyjZ4oSVgUI9X6rDbJUCQzMhpl6d+5
JCSok9JgzBrxDd5tkOjydi8AJNXFTKLErOvaohjn5KPHTKg5CZ4Hq3EQI0zT1TXFwVe2VAgHK8f+
syccfw+/PBOM3gLqBgn27RKTobi0Sx4i+IEiNrAoaqBUndkQP2Qw0CbrR+p/H0pPDE+zJD/+s7yw
u5ubSF5KoIpivPOZcazvoVlNcfxgUkKVDWOlJZJxw+2WRTt0GtvHVyCewVi56iLxrcc5d7+TAifG
Vz4WMpsH4nxv1l/B12JqJZUK/SmuzmmCOYCT9+XZt+EQkTSpEOTKlM/RXHcj0DNTVBfrFWq7CROV
qs0c65RAh9lIdwjwelq0QS2EP/vkhfyx4+a6V/KVXC/kGZRPW/IGc26ebhSU9VjDTApOJzBxp3E1
433SPMjEjc9u0ezUVk4hzdbyF4XfLj5K0bZVFk14TNmjbx8m1R5+agzjBFT1VO7SZRcLW73S/Bxy
PjQvl98VKzSoOwlMQZ/GMr7PC9CWvSXEV9v+AyiWBRgPw+hyQEFZN1mgz8NvinwwNtx4RrNgvLzE
ZXavpc7mcZb3ykuBumBVJtYE9ZypP+sftBWEbyab1jySX+z7GbL0waDqS0bqMQhe00oHNqnEjqez
EwukT2D+imikqqbRGdiC93cv9O6cWTC6w7p+CqcVqpCsmcdeqeMJgmtQ99YbcucV8VgFzdYhBpnV
67A9GLAZF1w+1MEtrYDeQ7uDXP8WNGtDbAnMCsckCvyl8UTSrykt5WRi4EWbG8x9hDEQOmKG78Xa
nPkR4M+XhsOlYPnyxyCY24ZKqKv8S+LgCNrAKMPABHOmLEuqgVTHJsQGio35Pxcb40EYcyAmn8oB
Y4ASUsFs1nv6mpvBIgP+aD8t2HAAtire3nQjhZzXCumwtKMKKcPgUVet+fy5GJkx3sTaJirrcb8x
yURIQrlQZgTUtruwQepL21mxsiMY/Yt1uiYs4ELMAv4fb/OAB/mTqQCjmz2lcjIFa/XQFI2oyAj/
GxXjPFyptAoks57QywI0FuKMtVoWr0ppkNEsnO5TKY6lJnW5ic/n6wwCNCC4e/REpvgXZL7u158z
bdk9OVoyban1Cytn4gp90uc3c+ozH9xgQcCttgcgiyuONk3++5ItG8UCbIfX1JOeuk0vPXYKshNK
NyvRVsxDkFWe/hs8dzBZ/XsWr/xl0VtFxoP6k3/qR1rFWFEovq1o/Oo1n1XpuDAeRMT2AY2G2q9b
rv5y25r5oyqq2DzBMrG8hs+xTNicBEu5BROqttdnC3M+9Owtj0EHJz7ubrBZ6FZwmFUlm5OIYZ/h
fY/RhXxTvk3hUb2lhCeEWvxxhpgeL4Pxmscn3yiVe1cBykrKefJO5hvX7Ldr5+XbjObzYOrxSnVd
HXdQUSHITEv4Wc6HL1M5BZ3VTXtRSYNLcGZxmy3mj35KKaA8FXgcS3JhQSm5hbRXg/fkkwPlJDcj
sI4384ikTy26C3ICpwW23tgEh7gb31wVLPSbYi4uAfiIyDdrt4t6ozMdGxKS6fGTpPvdlJThwFIL
RzPU69jlIB3FrctZsZ7Kg7D6MKL69kSfHtWSOt/rhny6q2KymPNSBIc0SEylTQF8+M0adrMxnQC/
G3zGpduzoWhSytFaDfR5/vu4r9ueeOVLQgYsiNR5veSP3cAQ4teAX6+ldczPPWzP2tabaM5+bImi
TT2OTo+IikRmYYoaGuyIs7Lkc+0sM29NLiFls70jw6qSgDp/7W9d2YB0vt2qpA15M1AVWLsPXgSu
32WJ9HvfL8KSNICHIuGgxWb6l6O8V1Ri7UIWA9gcdV00uBYuddgLpU9yULXXaYc/uHCP9YdGMQEK
NC5k+yWbhfwyqNPNC74eVDr5iZ9PY5BiBjMqyL9rZrgpRQ6QuoeG+1ExM/DZa2dIsqXf0u6VdEkX
afVoR7+TVLar15g0xGZotDBwcCJwRKVKo3sZU0xiCjxFDx3M0ofkOrR8Gajjj7jVquZ5VNxp+y4Z
gYacU72hsfIKH2R6SABn5Hu/PA+NPEm44Gzhviiwnud6ERq4tc9rm5sM5wZU+Kn5Fa69YX27dOV5
fWhZrTUuD2GSSTzCoB90bHO4v/Fl3EvI/NeYydQAxtvHHjGNgENL6N3C4Mgzp9fjXBE1VqYqQla4
iNQG62ixbeqnaQyfPtqn2TvqYGvy+lDKYxS4Q1b2BLmy8IV67w+1zB4TCOV/fe9XnQk85CAM76yD
jQp4J5TgthsW+ifQlDFXZpOK8hfPcS7cTpzU8dMRLUtqBpLqw6s25lwxXf8+NPcarmuHfjcgERJl
QUAThyWhrjoK0oGX5lMjIuAbpaic6wPTpB7oZFOd1vRlwj8tXzwiJqEZhztZ205Xswi71AjkUugN
ieaR9j6vRU7+/MhjpiQ5zrBgOaRUTJ4fRwNPaqA5OCaJ/ONXiiKoBx314zJ9lDw1x4V1L+a6dqvd
F98bfX9xEw5I6wKXWX89wTo/EJCTOspX4czRf1uURx9+RcpisryD8l88+TAzmDwJ2GnVW62CJ6NX
VO0Vc5UBqdxQHAX3JpUWgTZYLxwiZ1/4sPjQG/uAaipZxUdeYH3SP2aaP08+R2YsF2LrnzjhPNEy
4csJqARxJw8TALFpw8YmIcViMG/SUxTvwHgypPStEbLOjGfhc0Lu7eisCLCY/3HuZORh3c6xo1Df
KRJmFNeR/H4xJTwWshnNAPqGE9gzLYDIhO38dfi+EXY+wKhU+lfpRXjSC0rFY8bAzGmuJadqbQvp
cyG8E74rG+7N6kKS4RwiL5U4sqQbDhMjo/8MpPxNwqTktTJlTb5x6/QYRCKoFIrhtQ4++vSWVAYr
IQbWJVSQxm6+/w73B2cCfnbq4WhuS+mQAZhj8OtqzrYx7C4Fg+ZrHdgvsjSC9fO8SWPS/nSvJyhK
HbB+6wtUMTj/T5uFQWDdNt6x2e552eSqI6015EjssBuAb1J4H2lKZPkAvCuT6UgLLuK94HZFeOLs
zQGVNFGRBCSU66X2HxiEybOAP5DzUwbrdckvzt4p0esFsLx1syQ8gDTx92y8mBBmnt3xpTkpbQ/o
IB6OEVUHJSRpHaXxBEtgP6GhB7cB+46+7YfJVQmURs5GN2fzmjebMANptxzlZZhhXsMqnrpzR4k3
u57a72s5HRDPT6XoXrtUSD8o5J/07DL4W3iQSZpQ7fXHmuQfaNOhQkx/TMLqUCL+wFy5R3DqQscf
Ow6MH3egRPE+q5dDQud69irxU0qX0EIMXDIBDZomW3ItzhNbxQH4KPgJFZxINSTJ4hCUAAsJvrkt
RvfYppFLHJP/KOgurQzeysCi3WD3o2FcQ3rERH9mMVh+3rGTtnu6mrQFFFEDrkNMYWB0r+mqKDpY
0+fclWBARpUmpSeqreyTBjdwsX3O75or9KQn0OlMf0vu6MwgJm3bpgl7MDO7wXkJ/n3AkE+hQwH4
J4CZu0ksjl0jUoGQWve6oRN5ameVog7IQGJUJa16y/IwWgbqTdRjQJiQwO3YMqF9oOwnq5suh+Kj
iU3bkPbz28+0jut07imEAh8LTcfOHDLVVNkFcobW6V95eHRrWvRYL49lbUJ3NnXZSxWDyTNhFdI6
v9a6Vvz54PmV91XvT/drks/tm2KgkW9dey/tcJg6U0vcqDckQGMh9CCgCeibQMMpvJrehV7AvGKD
2L9QyPlrNKpddc8wQtOkXpskPU2ztCGePbxV/VEXFey4BHsIe2wC+BrvWlJOyoVsCGCrFI5HxPac
OrOnZ7QRM84+xwGteUks4TYjNJMuZdD2anVlKy0HYZTUQ2/gfWpqaLqgNfV0TXLbR/lnUyxZQYTs
kTeqDX+GbuoMQynBgAlIN/F34ogKkJhkHlmSFny8bf2jD/UB+DI/U32LwY8cMvS9tgqKNlpVjxov
lkumPNnnYShbzTCPDvOcDkcogMmNMNbX/GoErvT87Erw+uXZBmMVUZQKmqi2TrbGnYCzPYYBUkGJ
t+joamBrMoTt0YMbW384cKUnQpQeXyNzJlBvrKw/6691xI5iXMb/WlnHCIrWYkvR6xkiou88Y/B2
xpAtp2s23wUzaGBez7H2Vvq+oLA0jIT7s/QzFESZra36xb9efsbkGZi4b3/552hwjzplu0HKauDH
ZnzmxCEmbb/kVkteT8mjzSb9SBnTZXH+QKQpZ/QsPpLgaW4lwp4acozFPBZ1dCQc1StXWQw4ifk+
PwCa5B0TX8oSzd2cB9dhnKSR+yCDvkCzkd/ehg6IiyQfc0At9M3sGNGxxxCg6qtnwzGu2R+DCQNM
9dETAndXBsidmmFP8ZAfRQEgUjAuiKaFp83Yv2jPgZNhGEC0ctDH5J/BPUe/g8WVddW29cj2+joR
kqcRJIb2Dwoz2kfA0WgNg3OHo0hBOzpcIHod7nyy30xRoPyvJt0v/f2ZT/0D5I/jlvdOty9YAqbL
pBl80/LGtr+HjEyep34tpgqjf/zEZLMSoAboGNgTmSIc/ZYPTrFjKZY6UGyqntL2pygSYl6KCXYO
gzTeA5rSM1yl+5uoLyl/983IQgoNoOOjGDJowB+uAtsrjKfh+hYfAAOzVZf9gqKX8CQa+CzmM9Y7
2vrddY5Paufina9RQDzIAqb9bI/+AVy86FSTB5ApNprXDIFCB/1EQOMsorvQ2cx3pW43yiDiprgF
6zkMeF7/p+oWca6HsvV72JUzEO1fX77wzQ0lbZCCab3lGsXQS2zRN6HuCXac9hE6EKt1iN60CL9Y
R7H6YXczrmoYKi4m08yPxKm/ToX+XtNrdTBMEnY0iI/CDmWc6qfMf/T1UMy8aCkbu/uzsG0A4uqL
SrhaC3/BJpzrag737sY5zZVa/WedI5L5m+rtd6l3w3Rl4Ng+xhUWfVu56U/MAgHcxp6m0iOeW4vr
4NY/haOHYLzxlsCAOHBfy6QcYnJgb+fuWWskAUWieJnd8GNe2FX2zOHrVyehXquaFFp1vR9/DD+Q
VMibVO+cpE5E1klkYMlzZkcwChhD4rJRPP/13ectcIarh4950Ucu2/ByxZfGayGA8vfjmE+rBZoh
5TEj0ayAabDg7TZjIdjuxX43iVw2OeREHJZPaWBH5RFKUD+qYJouhTDqk0fJtbSLBa1tKWBc8hT9
B5S2TTY0LBXSY2i0vWLcNJgO5cY1IketFQU/daDwntZX/l4gLL4nR/YPd8iUhjyPTpdzr5kE1d/c
f/wKDEFYcyaAwHWd9dAECQWVTWohFeQpF2Jtsp2ZwM5BUb/HUhiNpKbgmJ7EbWcZRG1G0saJ85wk
jhVh2NvaLd+hsjykdJuuiScsmU6cjhYoZyucGwN85QZ5+NTKkeA9tXqFDFZ+VTUArX3zI8BxfFmI
M9kw67OoyOO+mGpSlfkbYHxPemZeoj4elLzcu0csW5vK1PbUa6vg8MT7n7QXmzfPow5JfoiTBlvu
N1t5/ZFCiUOOKWaP7nPBZl45JUy9Tmk4NCsk6MkgbMEFiIEEEUAb+Ja+uMn9F5QuGoJXdegl1G8R
rhhg4gTRWy+KRikngRZmHpL2ZMVSzgOCpOi/kPKfnmxn5CQ5TwlGU/N8MHTkavgT/riCPmd00zgw
iOmTaQFpJa0lNxHP+LOvyefSsNwsV+e6LAIhdJZRf2RMM2aVzWVcDAwwiXyxuk1E8qz5Hi7Su4G5
Au8TpwchAeyGPkooDiQiiZIEFQEvge3SASZrsYMnzCWwQtsoLa/3eDZBnLwwf3lummltaux7W35O
nw4Tl/kDVtHrCWQHMzb4W8g5AE8DG9duc8C+yD6qj49YWggU+QQxKLeMN+pzF9KWALLdYwx7BUhW
dAXKq1GEWem03HvCSI/jUfr00egJ7dpEjFwhGiX4d63Zms9n3UGBcWTmjdEiHOOUOurgRSyTot99
xOrNjPKGj2UTTUMnncuzJqGLiqP0oYNeni4E814J0UeGptJG+hj+vSW80wq/DEFPDw+CQEPHGcOr
1U0L36GXdnqxlUh2mMGWVsT1lu05huu4NICX0SFuPKzhac4+/wUAjZTygWMx+Yq/rqQHKpHFar5p
v3T6FQ3FA5972br8sOHN+FH08HkPVFXdkAgI9Oxq5DplKZLHYY1+VI4hAgGeAq2ZL7l3eXt/wSWV
0a1gwYLBUEkVGnrgoLTOsb4zXNp5CWb2+1cMR5cMET5wUzVMyMlem5Tz4hrg2NyADDZE+TzJccEX
o6MU+ghbxUm8D4S9BwV4hlAct+lbXQf1+KqTplaMIihNNlDtby4K+4YApcnnwo57BMCaBIOtw0lA
5n0Vn1u3dZejibH9AnfTF/mfU0CZEgRUzp5W9hdnB1igwXHtYVmqCKhPuZ7ZTjWvWLdV8Rk2uwkI
P2tdqhc0vLrpcxxjhBIk/e6hHYQc82X+RZxILxFofcVCsrvM7nZQdzs06RuS3CuF2S/3MhEmT4R7
2MZytzzxjLn2jKWFZPH9TsRQVRJyuaVuI6xfrbUn+32YQtSui61oaiU6KRH0+jugerTkKgT8KVCx
KvKb1AMJDMt90o8wRaIBTB55JbagA+tFCx+AFDtNVSxbrOlvs5E3ff/wLvg5A0he05wiV/b3By63
6VkdSzetfKsKskMha4HG1ESsXTZelHeAGxXLLILRL9F0aX50nptxKcQg/1FQ9T1hwQbxal2TO3Yo
+C3mjRZI4m8LI1kAnSJjmdZU0optiCxGsV0yw3Uwei7uGnD8WUMixTdUz9EAWN0C5JEOBpSu1uy9
gk2uBjsZI0dcQlvxwABDmmX9oFzue7VDhG4jbp9nLkmgMsQ/kAbJy0MWZR/nr5EBv5jF5YzwAMhR
nLSAI2ZUWrFMHNyncV+pYYbnxQwGyaB12foeKH2d/sTWiDgUsklf0vrTNtLh6MQPM4yAt/T6JVD4
lz+d/N+D14uqqqc0T4ePPp4HxhTvsHmequBwLcWmQW5vV7+UqcJjsT6AYsmI0LDbtveUEegDtXLk
WO34OFzG6m4hfY+VWFxxUwYqDe6+wNMC9+U8LFDgtl1nSVE1RbKQ3aDNeNVB7ig5EO8kzx0Dd44I
4fbzSbrb4Tag7A9+aBFlaH8mdrGcHeIy5Bf/JO01cm9jtpegFi1Vw0YVDswrqa3J8CPg9q10ziek
5fGwRLt3to5jzIXGrXmXrt4B8ffdrbumXocAyceC3FD1HO6JkhwgCEEWLxDL0AuC45CVMdT/KjRJ
k0JJlKVkr9Gc1DcC0IahFPkPXb67BV/G4YI6ZywZKvjG5awhIoRCi0Htqe3FD1Bl6xUl4HCFxTgF
CvxqD0W0Ngp2kQ3F8p3a84nTBzEpQ5a93TopurTuvSejEWJceoPtCYqbC8QdsNSxdwfQtucoxtNN
3CEeZWha6QiWJR/l0wCVt3PYJM0AUculpSlISv4oVXvdQ1FmHxILyeXqCWEnxW3vqMM4nd+Oh6ul
QdQkkVQpoZjwUHKaWNy/YVd2qeoTViEqbtX7MQtn+Tw0tJ7P23YPJpZBeJCdwiw8ywPDU8M09rGw
IdhkXBpPjQbBe4DM7OO9mSKEQSN9cQYnq1ElCtUeEeOUbazvVwSpGWT7BfJ3MENllcMAlcIbpuP9
XOLiFe0inceIQWTcq5DtXBbkCZAwb/LFY9Dr708x4WUayJvaKtzUTTtbYRSrDh+plr0/KDfM2S67
qo73U6Dv5fWrE2h/8FVHTpNapjelu4SFcFD4unN0LuPbejfzgnhD4+ajEYMXFxDzhRqjVIzTeqbB
HPjhO5Etqeho+i4VY1Azb8+l2CLDMivtkibPjl4/6Kgno5KiCmP9AKrdGhAynEguaqahB2dXi9xr
3zkpMUTd2GwRPG2bJ0BFRllCXEhPrxkLv/JwqV/OmlRDRl5ppq3Nv2P/e6x/KIxwjC+H/DLQioE9
2zDVdMg/eM8NTZUi1fMaZx/mXZvwSuBaA5B+EKasRcNou+tcxbcJJPjcQHVzN9jPcKPV5ZkltdRt
wLXlTHYLwA2zTnKAs+1jFuPYhQ0tO1nYkBd2/COWQ7qLrkAlYqiHnaQECaJeg+8A994hYJxwT8/L
2185MI3z1l1O3uQeQyoiC9URRyyo5R9WednyeiT4jeBC1bTLUPZUrZ9CXORwrswuOrxzMHCcoJqb
3RrKugRz7+VPzvgD7ZSgibdztjIb9VccN8t1+7SMB0rNNBbOmD8SbaTrmCaEb9z4vC8iX+JnYAC7
GnHegkPg0Y/wW26+HH59MAMBz6BCCw4YFaPZ7+9tkKGZR84ODcupAsMcv9B5mmXRcLo7E3aCqJU+
ij3iC0Oq00MxnVw4w0YvVaT42huhxsURwtAxyvPREiNINlmmtam90bgV/CDwxPHn2j3E+4A+vfWY
Ek+s/Z5NED4aFuZcg6Z6/LRLO/0gYbLWMHxze7wnpY7xWY+7GjBscRNHgNoWGVGolvaGCwvVjMQG
KLDTVDz5W+cSozaGWv6VW2Eyapy3bJ8Vt11fuLD6Tw8pvRAvNr6Oj0N3HGht73cH0vbWpnUq1lKv
zoKy/hxlD2e9kaKsACXEV4I5mFfBKkgEJUvFIVChKFPlPRwHOpDwl0sayKRtRg7S34N6f5U+gD9E
w+hnGf/YgwZ4P9uI0MoA20yGqyN5FdgSGbl27mY7tcx2EvML5ya+UwO0u4c3pcsONjQwdvq49qWD
5Q2U7xAiHV5BgQXwUJDXh31WKoeeu2uCg/kaJsT8MmRgAC0Kh6DOg1I/H6Vz0kM/meH94ECwYa1k
ZtK/Rkoy0ougGI0zakRhUGQKsbzgD/NdZSHeqKc+t2Pjdp62P1QBNef7dthDiZrNslITiHQ3oLqp
qLneQJI2lnriTbzJupGOzrJz74qz0aC9YMf6B/w/lRwayotTkL7pYeK7Q/HX0K4NKXICctsvaTxp
7a2aq5+ArrbKuBaLkO2En97RoO98urjf06C2arbmhmlfnI2AJ1PQGeFLvBgCT0bfjiBqI11XwizE
QJw+dRJaLCewRqlK/9FsOA9DiiS3stSE9fOTaBuXkuA1IFd+QiM+PerflgvfWG5nkIHXxieNsM55
ZXMeC4NZjeqaY03F/73Ny2huq/TFG84JY/+pLBf4lm/F2ID2lUHfHbD7WS9cofKQwMky0EkFRohJ
lv8aXKRAnk8UgJX50J0EPUHKgh4DWCVCuyAdBopDcS4wmXcz7N19siwAL17nfFrCfTkjRXqQRGhb
hP3UWCD1aDhhOcTZaq1/8r6Kbn7dUcU+ApANRVn+l/SE9NTBWqfE/YDhQs+PP7OScCKpOBKI7dCy
AeH8wgewg+eyfd4l77OoFOBBldBzWgcDIm/IMp9u451bu/SMK15iiUDL9zFLQN/2ziUm405NAMDP
N96OBIJG199q3AQ6uz5xOlzAhdQTOPbBolrC+z6PnVhplfRyH4vMDLmlhv3BEs5VzxkOhrOi1/3r
NoNzkFxRXCv8RByHfdnkYIAXtNa+kHDfjSxES/mVXeGFbM9znIwCMqeF+LiE2aq5GYkLOL5bolJJ
XAM2KczLgUROII300yiqpCe3p3HIr5Kli9PNGi1Wn9nV8VCZuhrPkRW9EH5asy6vOeVk9SYejIpG
JP6ewcHiq+lr4Ppxptp/CVsqVUTCRa/K0coc3wDqfsWoI8Som1p5FJsaEjWVodVSOJ/DcrInxMU5
tJ16JYChujwrfHzpxkkMf6phtQarTsktEwf1UARyO2ZIKxRT+sx3Z6ulzzsfTVrGtCB858zGVRbm
xsv0ldCanmkNydytleZkgNlqq7yG4YfHO6xY7UKOaPqyNHP7mPikvtWXfIR7KVnzHDEjy22XB970
FTkEkFnDgfr+84Vp5pK8Jia9V1pVPP8RrirYbT5o40XouV03tWFp10a3V7BegfqQYjE2huLH1uYF
bBLNphTWTwR8AGudXfRO7RVnEP7Ux/Tat4nca7uTs2FfqJeDt+Oevj3nOvIEk0MXf2BJufXDTyY+
D2qKbnqsriHJtICaEvzHPHl6YZfQXi/J47NbpmsOIi2LNRezy/OIlQwX+KCVBTr/1GoC/UWs0mIo
FgfTf07Tg2FnyNHTTd2z91G3tjP51Bhuh8of7GFvYf6RhaGZqOqSi9nVU5yCb+VTLxE2yNAfWfev
QbLWay3bk6EUu/XmS1LMjCpglJznHGjKDp3TH4ImAzq5sCqaRrZe0Yl3wGJxFwgIiiojAJJHnY92
1ergAnxbB2fXNGXSqkcyo4K7iQkF2yWzDEzweP3Vh71H2UklrajAHtlIEwRmwfgyYjlZDdmakbn0
cCZdJ+1+svMZvqCbTRIYHq8vhkvafv527HFd4M6j3Xx0ozxnBg+FXUt/FJkSzuoTsY/mPqEc2Iuk
zJ9PAKHFG8OpGhxqr/fvRd6KUnGmLGdfy0hmXPqHwdevCfPzOYRrYwilBiscnhZk7M9MHZfA4XIJ
4JAMlkhUimsj3iL3BntTpodg11dHO79wFdiGm86B1naDR7mUJLeywTDwqQSRBj+pan8KcG/WUBHq
dl0fLELbAIwQR5mgbOOZobBNIObP6NCJcwaOsiuPcMC+ZaSVX6IxaeMmP3JT8AFvjUvs7O8RsG54
mVnEUJQtoupiizqsdg0askyozxUxqe7cQpTMUDyUwIxbBb/BybOYQpE/dquvdyp9q0cmVJBSuoy5
JHL/tILvKPtKzGJDbtxhg/MbiXkPD9toSyELCr4sgPQlD1Wsdxku02cBlCIyRsM6UswK2EOVYmXy
edOaWCDELmoaJA7h+hwZHRKNLKkHSqvynCTLuE9grhPUCzBg+Liv0jcXgQYfP3wU5UPWh2s1ZMHH
I/OkVQZvy2gVktbs6Py4KgQMbh6+Rd9m+xDnuP5CWiS5FYIO70jdI6RRgasxzU6Wmxkjut3d5e8i
xwtRcVDg0rmNi/hckd8rEEXJ7PErdhi9yBR5f+s0P6uAOFaZN0tArrGasQTpUxssU0KTXmcCxquV
IqcyfemLEaCSgauJNtQqpMpFt1pyVcKoVm3Dpv84FdlqSlKPI17bCag9yEhdq9lWyBsyKM9nDP4a
N+0ilcGVJ5LenCHHa4OxOeA+Phc0JwM/xuwot0k1nF8uy+2jmMQtjZhkXsN4xn/idxjXOtUv6F68
itUBB8V0+mKeF2/tvPkRsfrQQCkbNW0Oc3pVu+sIWXPyVaPEqSNqLEg7GBlwRL0q3akEcZlLGQco
xZVJDZjCT0yr7N/4KMo76CtGLTIzgbcFgJVmJoi+L1u+Cb6l9U9HxbZBUT0vpGDBRQIsy37jWv/U
+0n5c7+miIWL4xb7ZYCPtqHr55FwtZGrOUiLJ3ItUhXYf8fIaOyvvlDaIdQPMxOkmVhk/SZJIkqe
5dYVOF5tlK++Mn/3IFRE/TrakcoOxSTlo8rHNXKk64ivSXo++Z+yPMXeprFQJPsrB1AHGPIt2gCX
Vpayb3ZYrYO4TEsfkVTw/mV7Asjf21KDoGTb7Kd8oLcQTi//8WJY3FB2yqR2umcksyWbSnvsg6Fj
+5rSTfCfOBE8TLPbxuUWXELlEM97pJNqYH/NO3csCgdSmJoOg3iU/QGNkrJJFPlBEZSHug6YyE+v
QcbPMf2h/YZ1z9wEdotLsRnFOIDPhK8VfsWzRbyUGb4vkMmv/j5k64hk3DgfsdYn4CnaSBUbVy+r
NZOg6vBAp+TCNx3QsAeKi5nzxZmXwtWWZbavY7cVYlo04aSEBmwJRTSZfN7i1YZbsF0KoIo6yVDN
W5bQuLhtLo2rTWNStQuhu3l/zHOQsW0nWx3x9HXO0lVHHKvbjzeDXTYlvKiab/pcKctQEu+OJvsQ
4pyWuzmHSvAkJYjwLiOkpJP/Rzxu0C4SE/Ky0n4QDU2Gr4GASXbJIHqfG7aVs14buHeP2PgDUYkn
D79DmGaTcsp1oFp72T5wGJzI/POTIgjXyESqBlTImzd38JuR+QtA9dNt+1qtVSAcsKk9OpOO4g64
fGV2PRPlt2q+gEdXkz3cIDjSECcVh9dk0EhR8TQZr+wNZWSD8Ew/8UK3QVGOtbpvaxfFDmjxto6i
wBriar08FlazTPrAusjpYptDYllA0CAivCWyoxxzAz9Pw/QvkNtcvYKQxx1FoZHyodf+3Z7ZGDoY
Nrem6JUpGPSZB5IRactkME8FOGG4ypwWUkizWDaYDll/KxkIm7QV67lXQgrtqLDnVu4ZGqOIDEic
9qt9/aDkTheFpPLwOU4s39BJ9VjJllb/rwqbMGdkeR+9n8MDr+iX4uZoL/VRDhMv2HEAi9mnJ5Cz
Do6NVoyFiEgRWXi7Gw4BbmZcZZW0g2m894H49kIkP/Mjymg1y0G59LmMMrxh360IX1rliPygaZH+
nTrgGaywGIDkYPiPCjyDUrMSizkPhk9Lkxv4wLMX4D8GgGMZTQR7OkpHYuVZoT2eUsAidOWl0Wuv
id+Js8IuntGP8ZLYxpVQ491eTVfd+P8/eP3KkwfH/9y7m01OctbBy1VMmmB39xhBDeIYlj3hRvV4
+2nRUrzn2YivtP0lhOo+rMcv2xY6G3Eq/0Vf2UVsqOJKk27xWkUlaWiJ+Z/uFr24lqHPMjk/RqtW
hUUFwjew4yNvOUqcwGsxmOxfPDRtoT2nmfDB3hJ2OfOS4BNlrFeLNZNNXn6saJgO8Bo+nsVVKL54
tGpTPJjfW7bMLaNA3eJKP+lP5DAG78mCWlZnBffkYkHr1uHgc8RmYJvCxbAI3v+IjCcd0M96gbXC
gkiUjJXSQKZktNP463jHxST/3VwHHoDSUbfu582N06MadGyAie636v8+7+eWDdUbGHN5KmqXFGh9
lbP26mk9cX0kjl4TBOal3o+aqvuQCbo5icS3M0NH1bPQoRTA/m1AAxEzVk6gB5PZQExai+z6b+UQ
iKG0t0hHtW0epYrvcTu35tDhRowC+mOMi1UzaCJfMmHRTwpWcZGVDAIf/wti6v9INgzZT8VKxhYy
h+Upvkc2eNdTMlUr0czEGSwCHbZaaCEWJI4yAgTe3BbVmIxxlmcIHlP77nDMtktcW+Dmqc9PLiEz
3sMsp1uNxaeeZ4HjMxiNb9UoE3ZV6vO4zi8K9nqlC/XqEWtTqLMoy/uBRIUTqqZ1Wz6VT1GoawYw
IoFCR8IB4Id7xnZAh5Wf50BzJxKftylxIINylI++c5MiebSO5DDl6aEZkIlZ85Mxtuk2n8MR5xg0
B9OUkU24s+AizaDcgHAQY5hkzpy8MG4h5heOMNLjivcckUcuTDBn7YRR2AYl0SpsFVj4aNf7D7Eb
5x1HXrsNlt9rKW8WREz8QthjhtgX6n0m4ZgnPtRl3sbFLvZuEeRcG+uJycnEB8ZwXNuAlinKvgLy
+zkftQMYx7cHuOZTcE5IjYukPKvUDBqGwXX7AYLi6phWolo1YhzcHhqG1MvTGkI6jiXyEvyozaZ6
mKxxH1MV3Pi/fpBB9/yzwW1uLDg/UsPC8/aG0ODj/AIc5WXykVJ+UVr/XuevAGBb4gZ+kp7o6eeH
z1ubY2aH+y0aGznbzDZubU8jmNjVDe5jajiartBdLOsVHyxVSeeXig4akXFuXFo/f3UJLIKp0oLA
BaserX0l4o6r2PdKjrmD+SnRDpWHUcdMjhZubNt3pfZuiZensFI+P29d0lXR0YeutkJXUFrtA5ov
yi+j0+pV6Muo/7tprqWHSDw8hWKR+CwRAR8c3Q4NfPYYbuiNiY/CcaBYtLlwfE1fqvF9pkRWWZiR
MZS+P+SRheHvgHkvJWjPuyhE9y++v+/h8ELv3t07fsUvEmarJF5Wbzcj3lkS26TEU9efpIiHfMpi
PELEQBFszJSvaTrXOU3Y4aYg45goDw4z1LH+TRdsl+Os7sD3+Nu2E0vq/pBw1NS1uYnnX4e/CYTO
Tk+5/eJ0fvUiNH4zIff+J9DOXItEqSIdZnhF5OQzU5RykBrMFYO7aOKD8Zx42SoO2gWOw1+27Ise
btpm2jVknPlsGi8YhewhC9gaIVSJXrf8rUCdUu6OAYQppgGI234Kw6zyDfwTp9C3eGPfM3v1x3C4
zbXX2F9kT+VZ/ES2azHmdXBI3oqUi+rVO35ULii/kKAIfuDI1wo6S54asSyTPlteROcc9orveuzp
FDPNNWUixCcaIhcsZcGYhlpRPNE3wUXrfhcPropMqA37CTBjDg2B25z/TLHHdBXPHLzxaDTDKtyr
lkyWPdXwZUcXw9EV+FlQFL0PM9mBPRx77icqG61AW3icP9Chay9YlxZ4DM7JCwqilSV4xxNuaYN2
q9+4s55XTQH7Le3gkJL6IDlEYLubcnUcZ+uZJOeG+AmmwPy+uyvuaOJrYR0cnLyQO9dIW1PMlpdM
vK9vyqAc5H2TckjwxPKU883wYBFciN7azp62iHAUrfEfsbz6sJUum38jL27fuNpn2LzOSdjUQuL/
BGULFmEYkNgcey855nIw1tnKJAx/wInDPbJ51ZiTdjuaVu6KVmLjZZexoChP2tzQgW7Jaf0Yic/f
Z0M50K/FxRJoRP6Qx8XszFBizq+AvAOKXA6/7ewJd1bv0YjSWGto0+2JeYQG9COBM/bGQa9Ma7dU
Dg5X8hIn70/4rRyKvnQ6KDckOYC2KLUkwFg1dllxPnXSR30VapdIozMNZU8ugv9YjhoAOocbmtIQ
mEHMCiaj1savZTxi28yxZVrzUOilvAUm05erXBC5L+B/FWGxf1WT6omtlaPeiFk3xAiPrsmdmVBH
VNMOBvD1128q57Yw0hwze6Dc3Q1T0KB6W4swamgKW/89dGDowFyhiA7Rc4Uxkeo2vMX6BWJYhS0d
cNqAQjgb0Hj82vC+gsqqJF/xgBq2GGT4EItii2TX3aVd4Wm3sOP1aPZJC9VWEMvtcgUcNn2ChsRX
OT6Q9JZ/90cq2bMmDrqq7iIrS4j38ZPisO+oj8VtnoA/foLa9fkR8bggpfVFNKhUj4C5xbCBr+Y8
6gF+Ga8LmzHYM7dvDjsU4S0KGpnfuPefvKg7tYJlR9wEzylsrTz2lkEIE0w20fDA9rXhuk7n7UQS
7QpWt1j4aaGWUiLn7lhsD7MrUhkIt/bY9mS8iUGdJWsXaWp4F4sGv0oKHa0rnj2p+k6WVkiGzTh5
OtyvLamWenAV+3cMMQQ/GNQXqqvpf+TgKIiiUI5nFXCHsAVKBzlCbxp1KpYzIRA2CAli1L4zgyGz
6szlYJgr/bES4cRNztB0eN4YjO8oiGZFGWp90WiyO+AJL0BpzZiVJZ5eF7Ppa1iLYvCvPDM8D7na
nz5X/ndU6yqFkk3T8gtdeX+jTChTjAI1hXA+mi9dJBjOOMidp4J3io+A1E7GVbug3i+qLuEHquJk
j6jkQ9G8IO27AYu9cDaR8Dk2cD9ZeHfg++rYW1YQ969jUqcvmxoChBMJJOQJ02dd/MfGYI1Ce8Nu
JtHNeA34wAluYMdZU1t/FG/6uozngdhoDHbTaw4AC5seQW/PfOy1D57EredC7ouUb60F8/4l8j07
/i/t01kYZg4eU9rO1+jc5pWcasdiev/rBNqRWgZonSNyYe7jRGpBpNX7RDis1bJLF31b6LQTssW0
QRjtJsjX6cywoAtjDourx6x4l8aKhj9KMPaxLbOtOamrIMBokALbyPbAuzIVdFzejHOCpjDN945j
pGQ72ohNkIOpvOtIaWtBc9N9YHrEa1FvOsZyz6KQ4ng8n0aIm/Q6XfWhGsQjDr75ADHAO5edoFbl
NGb6qvx8zrU8Zr+Jb7TNcxeqsSwKFGDq9ZttBO/oOj1tOxndK2ySVc6GTyMayMZdc7OvUOERNpwl
XoXGLeQExUqTUKRdU0mVqEGEmAP8bIwi0w5KDaFzFHw6iRCKL5l/3ESLXyQGDwwDY8HkEnDy92WI
sojaJMcgaEEyIM8i+r7s/+loWtf7V4n0GOb97oj9wEs72y6MVgCLL4kH3flsKjlwtvdBnaBhYVTv
itz8J55MEOH7tbjjbl1nkadNJ3+5HvrprK4vOuh9oZZWX/X/X800wDlb1wfunjqLVYxyM+KF3Ay+
TZD1Qikizz6bvFLtHadCiSuSyCjuqeBtWSjaMQjIrPwbxKQsV9UrLhUF0UpJs7laS56ZCSZaz392
uwTbSuotCNOlx9NRIpAmsfG2nYZ9S1F+ITAr3ooSCt0REy4c4969rqurjhblgIUeCSjxNuXepRUF
MOVSW3a/+sBh9+xBm8G0Z2H6f/TkxuAD9uCsVOypp4j4pldA7HLUHhTDUwZly+x5zGUmol7+N3oc
cRfFS0WxAKtYsFKVFaRY5YZDtyzhFmZdqan4V+jv59eWVXnIrkgNdDVrnu2b3qdzlN7YWSLq8DWn
EcTNFi/M9uIQf2ZIU6B1uDjBRtCbPxNin/2WpMm+BqrWM9YhXKE0nA1YTC1Pp050oRW7h8h+oIGA
B6Y5hffV97PBeFpd3eakTwktgN9uRDmUoYwW8247FNFyKJRdwxKYCudZzR5dx6O/FmkvwEj2CllO
0foagCCBdbQIvcYaizc/t1j27exHKBtHnkdBPpwOmszHFyYrSuLoOpm7T5jr9MjZF/65jig88v6c
35UX4IR0IdstlYRYek8iD++z+s0UwifGHemgL1W+wuIdegEn7kNqTcvHvE5mX5oMzpRQN9GDNWy8
Tp7W67zvYdZqmQTyZo/7xbROJYKW9/PC01SGtFWASKDUr6qrdNHz+af0FDBqdBVt3llIBaKNbkv+
V5n0c8zxnzkaFK7/+OB5/ImS1hDT4diJ/9ESIJKI0p+h+scy6xVsUpsjuUNu21FUpiWpqV/4Osxr
4prWpz0cfEcNylrHX8i6amOlH+a0+4/673nTz6Kq2qj1BIaC20DMJdCx7XIVkphs5Wj+xpSiBld7
S341gvxT5O/r/UPjstusspKmFMY7IxrCPP/6xTOQoxSFOH953xcojt/W9aV3PtZ9LmEBKOwY9uTe
+rs4woAuwk5GFSMU42yIT+zQrQXYdnLEYwFAw400XV173v2sRY4mjefEMErIPEoVl50dY9mAqo4U
3qG+j+gARs0IZclMCZV1MTYv3p0H2MXmiEAs3++99fjy18JiK2Z5KGfMyAHXRORZF3NJnh9ee7BN
M/DMfee2sxwAoQBhCsOK5ik4WmNTugWzJfw9GwLVCL53K0Rh9QelbUxXHz9tdDnnSnRwuX2NQITr
CRT6GPVd7oHOYsbFY9nfEWalU+KByqiDKs1O6rI7731Z0kINaLAzymG8HuN9cl3clQ+G9SRa2UC7
CXOfhjBKbqsstEIz5UNEVj6cs3g0/GMY31Pc+dr/2kCl7QNjQhdI9RNjBorapyIo88iJmncXZldN
sL/ih/bup00+5K4zc0o9uAAJ/5/6IHlI2joJRLfQnDVp1yfBRpK4k+Dfh1xpshH2WecObrSia836
4zxuf9lr+fbYWwCQ+0DwD4lcFvgUuQyrDyFOS5G+J3WkbTx1jTT7AaxqDd/P1LQcWrtLg6lPA6iQ
CdAfyeVuA5Bo94HQRxGxPV0HBnXzmQoB5JeTDH4/gq2aSCHnvA/vW0VZCJR72TzSpoT8A0xRyO64
OOmY7lk8aWfiXj9CKhwD0JSJ1LzBGRlWzsGW+XFVRVkbjEt/D1gj3RKi8PgtyBwBTxeylzYd1LqY
zNiSdA+VCbgg/HDMh9Y7kNQCV765I3JlxhcLCoGKbB2sUTME1LaJ/oV5WccQYAvxkeMfruFOmpAv
UkIWsKDLj3yyaEf6wRbaWpKtCsS69gCz9bEbtFZq2sq74gJ3Z1NbjIIW9nhBiz+J7yKrZ1exYSFq
EgnEMEX4Q7HwQ6fa65XGWqTF4VpA5PaWOsASgLbBoxKYvqbZG/l7nyDXEqbFyW+pKWVzhnFgLloK
7b1oHpx8ZFMcOC26mHA9n070+QA4Jg58pVwHVeBYz2wNMMTxiQ7cf7ax3i04MUMWsbypboYNZ6Rp
zndQmoxem9y7DVCftxDdinqwWo9sp5rY62h/hFsHWTQGiZjr9yJ9r0AZupdpLL7PXTpyxP4+7yY0
OXC3zLdG/9tqZnBmQofHSjYJldT+HADU2AcTG8OA/mYNhDWruUypXRw1tkQpLDaci0ZV6HCCMyQG
NoWRVlwrmglUDa3wBDiRTOZeD3JxS2zDUwNKVE2yjmNUc5YRPmIdXkQHGI1Z+V+o7sAjq3bBW3GG
86U1EAR54popcOX1cSUeTRh2xisg07ImD3Rp0H2bF8fjO0qOOBQs8AD8WD9k9lP/OxJgQSiZIKEl
bI0Q6TpvQ9lG89n7+zFJqS99JMireXnsjLx4blWcxibbShmvTT22EgrS2eF3j6RAQ9hCliKEV7Bd
UQdeHH28B3g//wk/9jweduFjbeIEeM2etMUZ4i6yzyy4Mrd+ZOHdMlPLm9mgt7d7xsHUGXWUxeTI
OSECXMGsouxcsxl/adrddfobb/g5kYquasvCFsAwHQKdYc3MczHrL/xekhsYjO+jU91NiHw1v4W+
nvj8sqY8Uusk1EDwQJSnIRgeR0MpL+WkRlcKqmw6d45A3sFQ59DNUt/7cic9EGeGhYX+rPFvof2n
kIUEPxopWG3KAldUpeWck1PeXWFN5hgQHxokBB6ig85jXtKdm7K8h+meSp3rZMv28Gacvqwf/Ld5
CdVBmcvYYw4U2lFCLez+rHTx7fTrhIO7/7aGhEzHlF1bTRvlcNlP8gGBmI2CYIT6uIbdP9uKbbnp
P6WdgEOmYPB02tEfkc7hBfi00KRtkXI8qhAZ2DSw4l1kxGodoqCbQNdL+jJYofk2ZsSOO6t+Qzdl
uEepohAKEONBmEEfh0fVKSGvAfSTp0q5hwNpydov6y/AcyzeN5kkVvx63A7boCHPxZe55TvDm0+n
2iVeZf6bX4kumC0Bi3KXuAxkK/oj4JbEWzlObNeXMbeWrzfnKLMfAVH358iQ7pjtxKhW+V3s9OLT
KQjZ8T2fjC0owJEgpv4dGj1CL3D5XEMxyZGydNabncGeQYjj1L8o12aQlPpvWMtbsnnNF5Cx+Dgs
cRitV2VBqB8mgdB6sgKVdGhk5T3zsCwQdw22HYwqp3fAxzPFRM58l87H8JkRTmCislBKemhxj1vH
YTYQM0uWM7DY+TkH8UMYDvAL6q7U1OjIBupcYomy4f2DXGjuq3Yqu+scGmZl6nsolgn+1nGLzuG8
Sa2WC4O7gqMb9OJp5xctMV/d4Y1FOdFyNcRv7ytwINlxVKAGowPHHRhupTSyH08LNliC7vaQKInY
spoY6PBF6I+yIyHHPfiC9WdO59W+vcrA3njf3RTwJLVTBTCdAYEUYmQWSDy+G1Kswhxtuv+uiDKh
EOL8d6qWrsgGw6Z5unfu0iaJjgVsnYqus0hfJt8pCXMRPRFl7oPCw1XpU8c7Eo4vOQRxxjmo2cDD
OOjwmuqMMidBkFHIUJl9KxHSqQpnFMpyxnDFMzYAS/uExzA5TvKeXg666DkyHp6QHIAPmORGke9I
qOXDVPFrbUqhNTF0k97eroEzzeU8A/Pl5uhXOsUutxI5THpQ8seF1GbHUoV09bT2KyryG3Y//8PV
YkTlEOou6aa8O3yAs/6trFGHWRYbVNHbvZ6VMKPR5NSqqpKbms5/7ZJ89kPn6lLWF8ZTTr3aHqcp
dNgixWqJM6yQQXD6FHEO6iQyFC4lEOZeBNq2jUVj89R+zaEmM0PdnGsjNo5Omo+JgvW/x3ZB/QvO
83NWynRCwHgvfDyyB1UDk2ibg1pb26BAJTPEr9Nm2KfCCY70axYdjnNjsx8UaG6f3JcYFwpmPRW9
5Lnu6bH9pKxyBjRe/rI5Efc84Vq7xE/zg7ZaEtdrRYR1zbQvx5Jl0UU5D+dC8ZeJD9bcL3/fwh8/
BJUrECshTHuui5taEbBNutHg6LvAg7nHpxcyeaQPc1aJNG4T/jSbmPcLjICTmkKGRrBdzklAKlk9
IkmvZQgtic/y344VUNCVwTszjPTrFhpJzH9F8fkR0JE8wEy5Z4GaLE9y73dgd7SvBDThOmatLaRT
4AF3uw6pw/Cs7PB/BrfdPws6ajrhsE749//CKYup6nEMF/Q2hiG997rOMs3Jcuu514txEvX1M7UU
zxIKUqFp8anGqff1Y9Q2kctWvqsqGLLTU3HQAo0YuPRb2XKkagBVdrPCj6PaAuS5dNw0ptf2497z
WDN91Y7PEovWkUNChFIA/XUFBUlqiRAFaMiLeCPFzn3pfUif7gZStyHezNoLO36s7QEXscVuFyps
29FF8W4YwVRLHVsWzSlGTUpI8DkKw0UW9w8MMr/BNh54aE/H+QG5wMlcl4Gt3dsv2rYse627XTuT
ykfs8qf/9spNjRbkRVJSDp8bTrBJ9kNJ4RUHOday3Wsyxh67MLQ67GPAJSLpo/wO2RALHq8Rsyme
EfjPAOxekX5iDfdR8b4R1ruhXYiGiWFYfdObl5PLmilfNlfmkp59OytOyu3/wudIDrTOEICHDmZq
giDSX/62m0GCSC5Q3W58bPIuGuyDbNfMZRyX+8mGA//b68jwB6U71Co0fPLHYZvcqy86TyDAU/i+
1ozYJXL/HYEhFU5+ciBBOBSiICNMhfZup/wSqOH9sKcInte9nCYvutvt7NaBEx7uWa8zr2NZxtlo
NgM6hUcX1nLwvWOr2+CPNPuugmwbzS1U0T58NND9MY6gynpebjaC+BDkzlazXbd5gix5FqnRRULO
cBpbPn3aCykRDCGedLqgAYWsWZWA+XwNZfiz/IirxgSlK7Q3eqCBSijjEqZuAgGAHShvhLZGoy0P
V2OKRwtTY8tyh5GNkfGAH0iO4hP4FkgdTpJqadM3Sm+x3e5TjCvBIpDljD91NR8NR3yZQrLa4gem
DQL9/38/7wDOvc1TrSD+wc7LhwP5V+hW8GqkrDN1TWhonfy4YU3a9+E3/VklxKEafmAPNKDoKYBi
KI9ZMQOvAGwJLi9yIe5w+HL5g9ewoEiIB1+e1ppHlX7u9g5QouM8Au9Cxk3y4mF65Pdedu2N6j5p
X48zSfUdM5d8KgJNR8DO1l1/4sn3mg7WAfxOcmYo4Mdu0rfRS3GojGEJ35/z7E96otK3nN7tCvCX
zS0Q6ogvAM6qkaozlMOecJIK511BLkf1pZpVYeRWcw3I49/lat1lrlNbhi+r2IpY4SpLT9aJwojm
B/J53dAxP0XKu40Y7E53uVCGdtsb7M1HbbfsZFesVJ6Zvy3jsqzJyZ7lWYlg9tsuDxqsSBI/k2v3
wBGTxDDb/RX63U3mp5lMqs16eExI/OzidyR6ikcgm1p9VqxPWvDWhaVkVCCfWq2Mys+a//DqReK+
bg8huJWV20+ZLuGIxCVX3mnbQffV9GR3bvqnTqamLn+TH4eMPXWJp4nLi5tzOTFCOPVTMtAAoMHf
1gDL1xFZCte2tsSC9ou3E/oSBBd54+G/rExUOtwpCqtgePBH122vdmByGqmZZvdUAlBXsbcvCngT
Wvnmf0wCaIJ3uooQ974vSC2oc9nipVPXTK1xbVt5UCWKjdI/H/X5Qr/qW94ijWrLXm9t5OnN6/Oq
9C5FSWeXIMwCSpIERSeHn9ZYITy429EtJdG8w3WHyPWkwDQqzcrzyJHot10zCPGE4Pg09zWZx/C0
4FTodIfRR8rWXsFEx+OzASrPFRNIr+zTFGCeV7znlxn2fZEJIyQ2Ky77/1jZ0NiCVSC5eaotxawI
ip1+87XDPQfOdUpan/XF3KLmffzi2Av1sRKMkriyxG877Kh3ZUWSM7Q7HoXWngkZqsmsZuuskD4/
KMVY+WlDk9b0GoJIS/yBeHzxPIEDbWn9mwK9z1LQSiFWHrMnPJ2wZGBWifclyaCia8OUPQWOkNR9
1gvGOV53295VGJXjUmH+hShBcYgUnAtDvasK/BNlS76AreNzc/6tregL3mk3ZMSs1d54ALVXrGVi
3OrINbzKAQnV7K+uiS4a/EaDeiPF6vmllGr19TbDa3VY6XyrMlld5L2qPPxHwEFIsfGdt27gsEbH
6GNwIk0+e6x5tX/sObLlHndDY9n/LlttSLPZRi6v1f7dBPuynI/GdSw05VfgwAwF7uqKvFL9evBt
tuii4wEPXr++l05gtfsQMEi5VQZn5hXFg5J3A36eSXUWODZnMfRvdFhrCNHwZmuIbZkfXyv/n37A
3m2jmoCmnBkRCoPRvCMHa/8eJQBpC47tMUljG73oZ1h6SLjNj5FQnNlE+WmJ7xCBWQ26iL+OE1V7
+LcEgQPT78wPxVCI0bYDoskBkPY/Ey+DsgbCkczU/hlbrjou16ORiJmJZP/47jcPPu6XPYbEfBwj
+x1Qu/zOAtgcHp+IEw99iWg/bP2IhxjyezDP8ZVbpCJMnXZWlg2xAJLmsATHdnwGfk9IkxPAXyhP
unaRwgy7m7ePrwsHC5dJ2RF+31FILT7rGNoKfqHDPLWJW7uAwDZ07NJRz/aF4Jp/uT94AlY/qtNl
BcV9b+ukJcYHB7cVlC8PahAYAZZlD784QUXrGAYtD8R3Rx1W727XafzglHEHvjwpa7tTskIQr+Zd
h2KaVT5MYEFidwW8PjjtcD5QkTgBtP7dlRtpa/MSP8io/PduHOdiW/XbkiP9UZeHrpi0mOSVMI7G
kNLDW099y5Q+wO84UY2Ygtcv/WCRyZPLkLZvG+uIMLYGFt5ZhDyjXmjoEsdjGo/m16D2c8u1LXqK
J4n59/apceWISHJnh/LhgSIdvRCepmnTnUa5TeadZdtpdywREfJKt41jxU7xij7kzAwmU78egOG6
3AhTT/jCdwGKV/zA8cmyBBNXu/eiH2BndQla5lWVnDlK8gpJy3u4nrfFKkKGxYlNx/3MwEq1csny
PBnSQ2jVlvflzh6vmmJHpgjdL19BsIZvDhVPPPG8xzDRz4gJhR4xZlKBeX4IN9y44AEJyr/qhFpY
4DMKsNtw4atqAxNi8F+D3jFJRtiVlgG1+9wKuD8+kqTJYOgw8Zh13CNfUwnFNsSD7R4NDKQMJe2O
c8dGXEPAZgRyOZMWiaTkBUaf+EN8S/sTwPU/gxwA5NLlHNNaqi8WR+hV8dbfk6YfzuE7iM0ADAZB
TkJE4RIWHxq1PAv+o6lfyBCgitlO2eAzeiOF7QoPs++lGgg8pAnXSKoWFXjaPIbZSOE7Mz5H6v6W
aAhGGdtzTL6AkD198sxnt9wPtt58pEgXzDYFrLS1qT23nV8bZfue2DTwIkEcS/2mpdOI25WnYVRZ
m9HmM88p+1GMbS5f80yNFFdHy2RnqrJEIvCGbtKVWMWBUjFaoUZXEFdcC9sYd1uTqg1b+eNXXo8M
KAu+J7kCR1NtLObyztKzPxbrMK7K6p6ZzzGwsWgplTwnI+mG9uWWXSxeg/NxlYFXtYPKfBX+p02v
jPjhSoPIAIqu/8/8ikjQhRBt6lGqpUtZnhcS0tknpTXpRr0s2xu8zqBqYxThZzvRDi/3HclFukPU
vFWA955R+BFJ9E7hFo3O6iOcglO3rBBTdjhlupDdgqa7M+QWBh2iSoyWZKoop4+Y54y1UxynAlRu
rPPIw00IsDTIYXRNJ7vqEGFinsHj0uTWGDFB2QZtSJ+xJzflnL8SK5BWalpzB06bXAex1UQTOt/W
djeGYX2wJmx5HazLRzBjFW5q+pmO4hcFd1WJqU7NzCa+sPVVjts0cFE51mEdbKv6Blr6vwOdnCUT
4dxzmBDbRMKZgQjQOjQeji7Qgrdh+pG45CdPsNiQBjn8jMUGLfpb73Vm/hprgftbWXgVfsoHFTDe
4gHzw9iL+nqRxuK6GQjFm3D5H7gkMjjJhSMkJ/0zHv2El4f9pWhVtmt3VAvB+TlzBVW38XKsKPr6
a/sMONKHwbxQ+DbtfX4lW8bBzmQKVnQObXGyFGa5dxf9oYo0p2gZ9ZhWQg1FrMrGu+ROuDZddadM
PXuxaRjkfM9EJFqENLL3R1bBFwzYs6kGzTVvUdox1Dd+atRNh3Q3yXZohgfqUKphcBYBn5Rvwnzg
hApR/ipiRHaCVlrQbIAf77nnAshav67w6RK008MnsupBeHWmzu6X59vgRzs2hzts6SnetgTNrV1d
PGuHKRvw9DAYK0NhwVxM+u9iiGLgLJ7YT3BvdBwnsZrbeUvvybQG1HAL7kkY7TwPZiHmiEYhpMgC
39G4Jxp1imT5UcFmpxX/x0yIR0d49blQMuEr82OCWSaSn+BjrB5joxKZddOlvc/6ERlFJ7OHyRo2
xxYAM9QhfyU2ChUf6fruFwp+sYzWJLAY1u3eHkghVCgKDgWSlLAmH6ZJW676BC2lZbVr7jUrGfW+
e+QYVtejlG3cFgmNu2p63j+9wDpZl95iwGIHPis+xhSTYwZ1uoaQ7Embuz8UxkMenNXxUVUU8jFa
2HYG7t9jIK6G3HBmkX60GQbx1I7u0agfp7jB+slPgDBJrtA76Ocqhc6+nsgsRzy7VqobC3jJoPtT
B0/VzAasRHCcXt4sFlvzpIOBO55pCn6m06Ymcler3g4L6spYHf27N+FzGMDW6UcG9jrYW8y2mLQE
uXRiYxWy2pmKQL4greepxVAnAgco/UFGufsqYD7nJNEbymGkO+iXsNwNiOMLXg1hG6HxZFHTPimw
DEvJSkdP4LysisUCaYAi2U66ZVOvMS6g0UDgtBreLSiy8D3l1plBjdDz27ZtTDRL3yrhHaLCnNkU
WcI7SlGpWfnGfW0v+72QcJAzIaGaBrCB6ay1B/BCLBg5Yx952ht7fnLMpw1DfpzkiHe9knd5aWlq
7e/1MkCTAqhyvQWa3/NPg7a+PO8c3qFXpq1ReriW9GJzy0VKdkYMrTd5FoHqRn0J/SvoYxnwutzn
wVfn5hipYrh0+OA5O18gzTA3jipWGrHbNf8TPKNt2ngFK+ywYQIfRSn8QEs9G8HBeXWy4l2qBVOg
3vaIZuHXdEK6ZHXQytzYlUh8jKfazCwHopziTLuCFn3sPRIzBT3CWYqOhsdg5uKeHVaY27jIgxC1
Y/TSPyN28oXo+3fEbxT/1U0MlqjCZnG5f/WbQCHvTQAGT5gUlBCeEeCymwj03yWFQNdjiwETqe5G
gwDdQX8q4/CZjTJc0e/048Y8q8hvHsBDDAQ/AfTOyLTSwnCIZbV+gFutym4iNMWC5/AL5e9l1tBm
X+SaR+Z558VTVkv9n4aDVFaESkylq1zaGc1xogNV67YYb025WPrIXWa4L9NGtfe/EFhRuDfOy6RE
jTFcy5VXO0u+WUnZWbI3/YN1BxU4YWYKaQ5CM/P6BvEdG4DRB5JWp5Rma+sipJOZkPT3t5tqS+wT
bPMvdJ0jcMsf40oPsZCUbJONBNKvJsMf36l/8Co8dendFE5M9EmJWiAZ441vv/5+WLR2rOw+SlvT
LXn7ahRRxDsYA4evoWtZCR+co2TNhrGbsvlvbMRutA67uG3IjqgTYzhRhbG4abVcLK1OF/tGpqmB
qsBtwSAL0TPZyJvyhN4eSG6QYwiq69htJy6NSsoexOvCb8HPdZwOZedhYqD4bebejvEPwGS/4vL2
W4aAdWKVe+QtjwFgFLZK+BZ+eyKp9fOZBGOOofAhup8eDwSb7/fj7u15XKZPRHSqioJmZ6l1Mmew
MYZcWR8Xb1ZNOSrtYrVcDg+OUHku7lg12QtVHZjasJkwUvjVcxWN5ROqdeVlO8GWbjDT/3E8G3QY
7LY0lK2CsI+IeoNBq2dAePQuFdmnLgtceuIEQQYFbE7IQgdTGJevzNgdgiqW8nHWyb/kBeydX7bc
fAproxlRYGFDcpMhmJ4+6/N7XymFdxtxg6sBkRzTgn8OQSbOaQ1wj4gwH9b1705c3k4rY9IcVoKd
zLAVrDCV3LD7xVhZ66IieCoXZwJs8W/+jxsBBUeOuYltiPrR3eXCpU2WUE86dPqrYJIVxo6EBIsC
b+EYKlZGcc05UuZFPL4mJcuhbTyc200wRzOebXWA1FqEtwhGHM4l7gcD596TSF32h1YpsZxjk6I2
Vzq3r9knKtkNe/8CZ1Cs7F7RRr0xmpfTiaE/VoBYSqBbQE8R6wsVkREjKUFr1/qWgxNsxwid82Jz
JcvRvHbO0we307sy2x2eFvE1MmXit7jbU0pbpExstwph6m/GGR1jyDf32wqaKQ6WY/RXCOMEjrrs
dp6PoE5PF1/t1sSl5L2pPpbl0jQ7QV0fS27Bxr6f3HiSYbZefw0iyxAu5uIHQiIxSwM49V1SLKcc
kZGCqw54x6PCvn5WSGUdEObGU1iS32kpXAGuAjpn0g2z7OZnkzp9PZ3UGs07cax4U9sUowY1WJMi
FIA5WaAydez6Ls9404UzZ7Gs6zU8262JhhS03rtykz/ZVCMqI+BSTmYta1zF3gUafnRiuwWyWEQa
66FaZ8/TgrxKb0ahW0NAN3djZJQ9YLs4e6E3cjJs8U+HnFyq/c2xFnZ3GK5Ao9LZ6pG9wgwNjQYi
S0T44mUKkBvbum6C+NKDcYD8yYvgwbwEQ5XdyUgUYKA93MUuDlsnQrzMbCR2E+b2FDZn8RCRraEf
99sFO+TuKrh6ZOF2tyCqqTGqKmSZFyWug9WDdqCV+cDDJGaJ2EeW7L5Fbt4nUqfJQ6Uz9awjvDPJ
49xPSr/zeh3e8q+JmibeC40XTbSr5mmxTORh3VeJLS09nxd3q3Ae+yqpME0inc4imGvHNGISUtBV
BbC2jVMX4GrlGhXAsPqYy/j+VOutRajVqFhc0kPvnvuormKog5e6ObJpRAabKdYcxzDjEZk/9Rn9
xd/IkjTrOjyE2RlUBo66G1LJ/FE+C6LskwuRUd9hh71mhrAhO+hh9LPRsuYxBZaEszDqosgExgzr
fjZXEjIzDMjJ7BPvOYMNHaOAgXqclk4nyoxFmVAQl4ddLPwHHbuNl/E1AyUdTQsl91scCvkmE2YL
kHOy+N0VtsjmqnUm8MPxGjpB7V1rCTwukU1DQV3Q72isFWaKIX/UIQQOPDKPTitpi7T/IdrxvD5t
TbZCT/i3LuEPhu+TDqWE0AVOI48Flf7n43qMMgv5v8Vcb+6+b0B215KYxmSHid3Mcbu0LfzURloj
bofE2NAN4bftQ7ZF5nO8ppVetZjSv2lWrLtvsn2h4nRIq8qcqsSfBtNLq0tUUrkOcDYxDtayIzAe
nOT0Hhfea69XpolO+NM4hE2zG+K3DcHqxKJ49G1A2TM0EGtnlgRsYdYDC/0McCnjlNmNXmCGGjNx
zHB+PKAHrOSd4S4KgHkizwErPejGOGxShcAAzEc7Fg36QkN91ZI3PHbeBWUEhZ1MkvZQyxHWJpss
YC28EBSa/PsavwXjXC+FW0pVHOvuqgIIhJ+cGrYYJiicvWq2FQjdjFe5PAuL+8lPouAQznVpOM3k
OWu5ML+kbJSrxS2P0zQ0uHyBWw5k+KssVEhQ5CpKJ1kZyoz3j7JAwo2Lr0o8TJybmFU1nWIvfO9y
h6QfIMgNUtRUULDDaKArkGFnI6PomG/h51Q1DcWFWU4oIMhUisS1qFbvjsjLHKxo2QZLMQe/DS0W
ogjGb20A/AifMg7f4vEUtwH7D6oSYQElu8gnecGvrcCMvZ+I92taM4uKdy9ncimTtCFWqXr7YzRb
nvY0p/pwadzhHxsLhbRBtzBSxoFQYXOmlBVyM+OA5D0MryALzilIq1yViFf1pZpNUDobn0l4xM/4
iUhoMiCPeOe83HA8hm/ghCTj63jv2z8C1Il20S4xKoSRd3YLqLcdXJmKtgP/cSPvElzbeOsayJMl
Wc1UkHpxacBfPPFYMUJccf+GTT2FOde+Cxnm0K6+nlAQtKDR5iFY92a/i/kdC5UfV45ux1GyLhck
BhUCeEqqaokihjQf5DRL5jn6gBrCUICoX97ZnkpL+2pHy6EUmKq+tvjT9OOrPVRo58MJTY+6lc8f
6CI3JuSnbEk3eDEtdRY/vuni8Gxva/JO+jAjkOzOESJtvtE5ClGyMybN/XZf1qV0KchNoyO/fgeX
GRU96I5jdRfTVkYFOu/wn41Csr10YSQDhBh4GzfX7JbHVei3ZmPnQd76VoBHj4C0WFPRFkRH4Jhm
2gkfJAGEd/jA3NQI/o2Tk18rZ7HvERsqXZDMxMbjj1i2x4bn10mpn4eK3agjcd/dMbHahl1lMktC
3c73k656UcBGasZrbUrcbIiLf2OqEndvAf2G6yHVhShjTurngtlbk0ko3ucGmsJIwqE/qPsKYgJi
e0zeRDYLWGFigWkMRoxLx6ruHlyNUSmEQYOFPRvncSCN+5262/QKuvIysUEwEW9lBg8+MtCl4mL5
SuVi3rSPAVtBt351QdnSNtLUjQW79cLEaeDUpgtjE2QPPZIpZ1MsOTC/eHeG8VJ+O+JglDlSuKcu
bH/YQWgNjwliqLKCu8mAzjxQ1WFZpfmYzLWfACEhSmYo2fmk1R3hMP8o1T/hwLVdYiYmozo4Yn7q
aPlon0MerbfImXjqS6gQE54x/ZNBUE+ZijNeObdKk69wZL7g1diu+cW2EpElcl2tsNQrQ0xnRZ18
BmNlH8UITIRtYQRuwDGylHGagCLlVERBUoNGjqEjaWFqZJZVKL1gycvk39USNNCqeXFr6oEhGvi3
JJFlC5m3BPL6AWofqoLOIu2hfKsK8uEZrbO4VoGz/SBYU45EPWKRcjEckYifXwWH/MIk5Mix0dyU
tVBWqo52e6sCYuNbCgmlajH8A86taJcXe7DaaAlpLZoc+cOKyj3kqx9dAUJnUqhSdK6maQVGuaEI
eGiuDlgLQ/rO7SZqpu+ioHv2xw5lkv028UZNbsMIpsBxn8sJeZsGkS56IWMzGLDaAsgHmveoy91d
9kcucNcpMfEuhjzOpMLOZ7363VrV0u3UoTok/EQ6AREZQEqMglAgyw+3ymg5rUWi9+IPMCLwt2BK
TAZErePzZXL+0jPYvRJShtzX/LsOd4wdIGsDha+iF6lDwPSe0/Fdx7syVPSk5tysdvUHQdi99d5A
XDlzuzeg2NfWoTVs6W5P5YOV1PgFddIC2xE7nVZlHYsGauugEnB839dZOgoXau8QHDnn350jVgbp
nE4rWqkXao0f7GDdSFmG7ZpKRbBC0V6gMbKVv6VvKUGHCggWSxe7GXxkQ7soNCmoT+h+H4Rw4xUE
vIk32lXHDjzkZNfhmsIljX63kkSqiY0PR+QTFu0MAg1ZKEeM4Baob5J4/yalgP4OZgF/VquXJZ6e
AP1O9ca5d/jGa1mXviaE+qejrsVVDQubKgusa1F3tcXDWK5sPAqL0DPtVSuDA/VGmdIObTEwYu7x
rGys39QfuBi7aVhEOMyitndu8+ikUxf08zlc17Nf8Kh9tP3Asl+4NKDjWd/d0Z4/OE0N8IW6cg1n
bOME2lXVbcoS+pjrW0WwmxrznL/R8ms1Iwkq/O+awchpKQOBoKSDf9N9Y03Bw4n1DhH8B6O7QX2N
qVhUzZhQb3N9Vc2+W7YUXoIOI0aCRskGJoh/9s+LZArCDvUJFgyVL07l4+y0DsH7KRBD/VSKVNP3
BownBQj7EN03zVxy2MCACKZjukHGq+bGcPxd4T9RIwmjO8KEG/lEfOeXDZdqIzMrmQQWzdKwrtaw
2N/hDEyNcryHUXALOzL3OFOSxuWMVxJZcDWnXioOcoJTAwQ0mtF9CwG6q1s/thgZVylBVoYhRtos
osLJrZzJeX+KTBen5t4ofmDGARmqPP/RhhnpW8hgYTpVnFGANyavHhRbH1tLXdCHT3Vkii5C9Y4A
fDkacl88S3Okrg25k8kMFKJ+OvSu+VfWotyASiU0VsceKoNYDj8KGZw5W45qet7TlsUf0fqz7Lly
JFZS23jbLkyL1GDYOrLjsvqaMuM1ncGGAQ3/b/DfJZ0tRFcuQtAGdwDVsASoX1FV30MT/2qFCET7
3m3PItOBsTc4Sp5057p3Nzw8VMtmQD1AajoL2BpzuXnNGRhiwIEA3JrtAggYMCbm11tgOAjQdrMb
AaIBd05I27hx87vabSHokk32kNZF6s9vwyihgJvaTjC9mUMAkJzT3G6DkDNm8Rzsn/13d73gqaXw
jYLg4NefFljJJXqcKLFmCONXswfps2ELBc1plh0Tqo680RpFvnBflf3sn1nN69EjrTEo87JIlwOT
N62MslojZ/WySdyUEP9hSiKmLMAu4zJ2BzM0T0KALP1WFPOVA0ZFe0FwLwfaq0bXe+LI2Lj/KIvQ
JyvTf3DedTP1wXlTkXVkuu8okPKcpxIznCYSeh18ReDrTfi7KXWUGMAE4aYzEuUfAyHX5WMXOCXr
nzXLZDR9SD4qjdvFCarQlHJGdf0vhhpTXAaZwRaZJ5x8OhbuCIOZZi+D7wPBF4fvclAkZWhCjxm3
6BzokbnBPpoFGgUkm+ptQ9EwHBcxNnDc6Wy0ltxBJpppOy4bDnUfpYM/3qW0kmpQM+/xOHpXGzah
SG/HC0eKYsFlSkv6X2iDIyuQmZ+okxdQXrueaaDQjY9ovaA1c8UbHNPq54wOTQtfxZ8nNaoW+fB+
OBmt3NwtZipafQM5qk1RdgDjGDOWYA9Rf0puAnA2YZXdvOTSbmnoNeOa//W3MQkcKSy2QUKbWbB9
EJOVMm9CrlWD6JOAHOgfuo/tD42KX56XH0WkbK3UpZKm0ABsKFb3MQHuDjCA0oUsYvPiUBZU/agW
V50caYKNX6lsX3eb6qCmJNJ131ZtqoPMWz0I37i8NVdRO7QQKQXjKI0SwQKvASD5EuKqTcIXYC6R
xpprxV0LiYI0PgIziwrlYehFJip3P59tQEzW6bC5o06F6KKl1IxdXWWe6QtwKIX8Dw1BHPKcVtWE
xHrnGw+QaTbqStKMw+gYhcy3dX+qvz/kZlv8e6DFdD0VbN1WKb0TUBPhoOdtkpVGA9oplEz582Rc
udLgBoWnVZsv/hEi5yMyFJMg/o5H/URDXr97k+4b/fpOXRYMQTgKw5SRkiCkaVz4GYANzQo2OQa8
TtD4cl+bbBdtIhxpC2+kdElLrkhaiXQlMxhq7YyUb+M72lbU47l9L7tDPcXbw1965890lIOC7k0A
eFot0mfZryiod9DQLcaBDYN/wbPdjWxHTGhYQS7soIoBHHIO3bOvRPJAkJg3+lkRuhdpnfnh0JOM
0y9dK2aId6R5Rl2Dj2xafLeZ255HstEGTPXA7mBBLDhHOAEZtNuI1SacWEVu8uBMXLNRoBF/iHK2
8P0uOVsjEvjeQjITjwsSsMbgjpL2MmrshKSKFLqTTstFEW1Wu4anedVnjK/Xw5r/Nr28fq4H3IsA
cD+IA/EaDs0fI14y/o5BtpXd7xhm/uTdzuLuvJFqfO6KtGrgTJK4aywlxX0WfuboEdR+ymfO7XKc
KMcVfa1u86NZ44phXI6zx6PlUfVUFmuPg4qxcS9i9qPqtUzsDu8pkqOne8Jm0+RxA0Yz/O6zae6T
zXTZVJQlFhhuQdesU8rLyewbQsneCwalq5nSv6tGbx2mqzoWFDlG97vh2XvY4al9JEX6hRDVizX9
UZKKDnQWL+KayimVg4l4yp7HX2P5kG1qQttFTSnFWQnJ3F2xzVj0fpOWKEhSkyXb+uG0C3QNS6SB
5K+vaiUmcDQdw/+rVBJIh2RHi+xGeXsDgsxRu1jqXFZVu6Lofj5sEsHn8ZPVhtbGZZoXatzT1J6Q
FlqTiX/MMTdrWY5y26x4YO7k0v4ZBayiXOpvqd3AQ1+5/XJApuq6kW/J8+kQvMWq3DiFPSO8kzgv
MsyjJrsvhCVcW1AnmUOE4gbPLocPM2HG3aRhLjJ7D+Rf+UmcFYbXQTneTPmPqiBLGQ0w5o+y5rmB
0LBmXFz/vB/XPPx6sOJhdYRNKfv5fILmesGgX3gjzV/Dx6G4jgsol5L5UO/hFBO8a/RlvaA0QWlk
xaXNc7tv7l7kxNjCYaSbs4EVSUxlOOhJKlXl3KH1ySuH/RLG77mPJfgeQ9UxA3hR4uke9p8NFQtq
9zwMfRWxfDn+E/z8TLQzMGcr/xsWPSSk1UG9QtfIfR/3x6FF5+/sowA4u7+Y29SDZG6o+663ihL4
Y4oLFpSm9Xn9Pn9hiNMTI2ksYxymUuzFjqtYdWFfYaUoxi0RD9a977Dw6e6RCjNbfBdxvc1C1gzK
qqWvBbYQGATwLaT2OzUqbgqJmMZZmJbRF6YX1785gu0GggC0gHAXl54YvKST6RI433YYt5DrJ70i
laFTG6an108Fo33hoVJ8U8kDgm4ImzQVtXZnHkWTW/qSyprn0E0Rgah+rr7onT3X8DksCktW5cxm
tf5XSiJHFtk7temtz+W76VMHzvhY7z5Oo7ATHkFfY5aFo4i5yaWvzYeh/0U8HIkQE4JiJyVW+ryA
VWnLduWzJtEbuOwb0IahMSpitAFvAG6YQF+KqpCnIJx/0EF880N5ycyYDhkM8EhExWOlwGMKjAPP
q8TL9lfszMenr5HBTOp/lTzI/U6G+/FyuUpTJ43wy8xSf/26hVVp8UKhkXhdgNM2Orh1L0Z1venS
7FF8Ajxavp94CdXip9Gpy3vgiYPAigVgO66NYI9aspVOocwwy5UwmQXv9KiYZuZMwoZELPmVUtDH
aAtgzcyjoh+BVlWZWtIOju1XyotYXqg0uEcTKaQlxlkBLLZpFwPTm8cTvHSv86W7FcdZ/nXGxDl2
gliA9T39b1c0ryPdfcKMSwXC8ov9jWZOhAKVALwAXBPe9SFP0VbP3mUhzrq7NkouiNihBRxAzhT+
xm/+0g5aElHDeTPY1FujkvtTA0MoCDtU0vrGByoaPKdzmeG6X12+ocC4KU1VM8mwvphgXdxy2CVF
fiq6w9NmICIjq+1lYwFUbLepMjYtr3Z7ccH7M3mgAZknSbgmFfxgOGH7SAbbpPSEByoVYxoQzKmJ
MGu5SjukE+H49zMB6WuARu8u2bYzuFnxdKBVTnebEvOr+9H036ACUMwTDsF8FOFHuF6npo6cEtCs
aobfA/pelyocR0QDjsglu0x4734dEfbEKMmHjMnfX9gueUbsC5i0rjIhcHVtx6/AGgArnjtroSwf
vKXyMbn7t9TksYFpnEf6rhf9rOhY+rvxU52qTSmviyqS0eCC4HAg2eovZd2pShinn9AbVNvds/fl
roXC78kNTGHlDUPcKr+ag8LrUY76ausRd1hGYy9Q6zph84IklUm+2fXZpXT9NOS43TNDoc36WtDz
V6+npZr+/Jz21l8phUQHOGWm4Nzh9DZ4oC4xKYSWI1skcbhLJB6FvLYILdSWhldEPACd+yNcn3Bm
K7Bjs8outWlvbt/n2SST4q+X1zVl2Bhz/yqgLeBU97TA7iIRBy8NTXP3vpjMTR/Wg0aWoE2n6Ecz
N6eHCNXpyEDR6+YTtq/+91aVZWblETK2R5hq7AP+wSbuy7F2ScuEdxuJMhwfX+2Fl5UBwLEWrv4F
HBsfpByJ+GEMsuMrRzVt3Vn1T+4Mvei8ytq/e/rb1/LQQ6/9cSm3PM5NSehHiUl/T0KR3mwb/6hu
ZWo0CgA7Z6qoMHkjDHPu2vhPoPDXzHGBhUtZgpu1i0IH1w308V6b6Cjpu+CxmyZ2w46v9eOc1H3I
s/FK8v2RP4WZyzq7snsSh3RS9uCg7oytyRnOXKJMdO0ESLvJI28skR+M83TH2NlUZK7MTbHZI8OF
bqvp5MzvXoZrRLe8cXPp4a8IIM3JLAZcQKegiSC+IlH/pwwPRwctfLyhdjRhcTWqB7QHLipjwjF9
MGmqw1k6SnDVC85XkCpYeX51AOLe/fDWhwiDUgoQUL2Tst69Ff2RBrdXUhgLHW7tbWrZHteByFfK
125N7GnFc4j6Z6VsiSXr0SYYBEhQRK0MMUiS/fAf50qmgSpnzWkmhMe57SNBY9pST/Sry7jRgGMY
DKYPX7eSI7Gq+3zAoRTNbApxroCg2eLqqkOCNMd/SPfcBV2bAbAc8guKhA4x6BH7n0jjJFPbbpbX
Qwxt61FyaJmhcSH6iPEdRFxjYA716WapxQkBzVqpVasD8O6tHph77j4wxnDzZ4ax89dmdVJooqXn
D9mMJp2U8VdNgwHVCx6cCNnUAhGfZIkm+l7U71oI4IzSqMFc5R8Uh8K9K6gBSQVMuquOYjIt6K5O
WTiCI89kCT+50YHO2EMoDLgdV4M7KxQn0Oyril6qIk5gds1VJ9AtiLXfGLCc47y9AlhJ9EE+Qh3X
TfWsC17diZsetRVM7vvziKqbSV0ELACrobkp9TS8zNX03q55o+8qz2CO1galagDh6cUCBpx/aDHl
yzFapWJUQA2nhEtt0J0vYQudfPrp3Csh9TQQYDQn1vCxruIQ+RJxYMH5a0IqSLS6JkDihjdPE0B3
dxTjYgnp2r0YxIn8CY654c+eGgT8Oa1XtMjdGzvw1MEjrfw0H9ZyBxaQu1P8JZLYkt0+6JVdqMRi
kmExfYQalGzkF0DprgOkFvQfM+fWF9Qx3pUQXaT8Huo6O9vLlBmoN8ww92UwdZOaW9oDo6AjULmx
0fgESPpu1DxpmALb4Cj8PWlYmxbnK9dfIpzU/bNE0x5Lbou3K9YAjwHSeJkpDkhZlWtz/o0FuXhG
NDlP3dYl7lQWLKm7fFyyrNL45mmRKfBtK47GaUODUrQfnu+bHXgngh4UdcksT7ennoHK3rGFdtR0
uLxcnauLdMOOEAm4gaqVNv2H4ivlTApoMUvd2lQfT3AVq7iqGUIaKV/QK5n/p3SD9uhfKEyzVf6P
K9WOe3M+NDvYWJrAM+YSa7AsgfY8aZe6UZFJsUxc2BIkAISJhx4Ap+fGCh35dF3jPzOx0jsb+2nq
7fnasspqVAF0g1orT5u5V+hDRmW7a8eP8QPvfc4c7/4wkrkoBlJnfgnep/K/yutgjD5IEajWARJj
p5wpX2zte6lJX5ex3sfmjj1JGWzwfLAWIYIV0v4jfklFZb1k7HcEdagX7LF3i/QNaNCKWqlEJfyZ
Mr3I0JK+6+ZsIdJ5LgcGaMhs5b74pHHD3Gm/57dJ0n0YrUCOrfCBMShMTNaOsDNyA08c/sEUGRFN
sSaPAn3fz47K3M9aiu07f01p/PIO6NXZJM4Cpt2GUKyklHafg9uJyUxPhYCwO2W9BpfLnujCiEqI
09yu+hJfACK6LZs39F+yy+g+LPNgXO0j0RI5sPwHnFBJJk8odbaDxPZmmuBPyDaXA4gmYygkGqC4
Hgj+MsaTs72IOLT92gEq98H8yAw9WoDhhrSR8BfeogY9M4pqDom8MS/pvEtN1Blk8X4ZLf2XQuBm
NfMXw5l1rK252M65VLinoSqgIKeSQAqLJ27adzpHdTRPduiqyh6LHAiPfVpK2k/Ap3qUyJmBYVyu
Uzbezo8W9/lRC/VBDZmJBZuV/niyaebX2lJDZeCxxhIhbn0Z5cbcwtcY/2kKgfeNarZU+PkCUeyk
7UhPkYV65Ml8kePVu7x0/M1KsR7SSPEKO9++MHhD3s0q0xVnn9ANdQEGpdC+/5imcNc/tGro8xSq
n1fr6eSsHwqFiDkv7lTOMXQiWb1IdwVWxGCaNyXRK694P9Ht07nJ4FZO9bthyAuqTIsdqdTT0GWy
iZ6YuTRDQ6HxAOJ4qSCcxLbfm1X62XWDyN9gSKl95b4i+IXqf1QbKcdUYAwxGW/cpeO0nEuYVE2K
IowaD7xl0D91FBRf7sH+NZnawyVQwPgqBZFN+Y3hqBJiE+llQGiWSF3u0dnGolfW2jRFYrkGb4mm
JnZqikjVij8K+Dr+O05zp8wZ+PAlA1kZX34PGiK3BUYUY29pkuzuuNyr+kFWPFC4Mx2rftigBgyp
/d5MLedLonnpw9csvNCa3S1SMp/hf6or0N3ZnIQ90ybHyL6qXdK0ASmmMjRCpW2No5zMMP89/0gZ
S8g6Y1oQU1QnUnX9iFKZ3CEsEEKsO7hLVyQoNkHOSYC96tXt7YMu0jPkrW9eeT2LEo/kAeujBsxp
ToeOp1/CmT2Wb7c3HjBZwBnF800fOe0VtjCvLzrMVpB02RIGkKSytJ8fO/g6QhOHN6N12MRlitEB
ZNx6fSV2VzFzaEcRTG8ssmfthue67pdTdwt1VguKIADL22am2ag8+dDnl6CPlyNRKcHEL/wJ+Zo9
yceG1tRGAbE0zgeVjCm4VLmzRJ2sYMUKjoNIcYuyGqa2V24h+rifqttIAnqVsrGXA3ey928WqMwR
0lO2UD478lo8fy6HizcZm9KYi0ozl75kknTIbiqzGvEkKGS7WxsALCvcz9lsRFFm9VtHusc8PDNb
szRdh8goDlLin9j+k6GFWBCJyOOl7tHs1sIy4p4r1hVuBePXo/YL68lAro33bRJWbDVZmOObEDs8
lxZPQwFml8iP9UyJvgljIDoaZiR7J7Z1UgjB8TH/zooA9mYVe2CPJYplvwhDJmcKqeLAb/SRApiP
zuaDmnP00tSjMa7h2vT5XWeUSRCv6S0qcWXi+Tdz4oS4Cg3x07N2/b3xkguizazelNWp/NNnpwNi
hAaaHxeAvkoVd4Yes2VyAoQda4jCiQoGnOKo7I5McpA56xvNaNstNO33A3AFzx4r+XGyy2NHWSgy
CKlRLnnkIRX7oQreBVhjRByTJJrVgz7k8/TPfCvLoExN/8opzWXmwkSaNELAfeCm5zsi0UT3kTgx
CB9Ds/vGw0rj3GZ1ymOdfe3Y3SsrFoRi1Td78DB5vkbfQkBhywcXRjWPr+Uvj3uQ7nDvaMa9x9uH
8CyfqZUtlniaxVgL+oD788a+YxpPDDL5Ci6lHBYOj8iI8InQnyB6UHp2TYhv9o4ZQJFu2a/omWQU
fVQjwuobvFc6LySdJ9ym1zI8NeKzdsIpKEqBQWDXtnRRhcFSgN4ZlTd6+qkJUHEQDZlTmJ42yOKB
1U2GMytBAXOOk/K4RypKkWbwlWjWhSsBQPGkcSyD0xl+D550qIMoBtbcZU8Rn1Tn6+bG+L0rXR9B
UqTPbsgSedHhiAHEVzI1ACJndMNXjWlbkmsjW/33fI0kkTBMpOL+SyoSBj4R6VmYLO7976Xfo0em
QI6glVNyFRthQPd3K8PJ/eqXR+jsQGX57MjHsPqJca7rEq0ouZxguUHmwd9nf6WRKyNj2/nsx9nE
yQGGaJ0FjLyAsBi4qfzEmgM2y4znefctpERp1tUwqBk+iDcUqkPXlP5JrHienXhMaW7opkAP2rWC
jQlmoWZZFwgdt+t9u7Mo6z9J1vmgVCFOXTQhl4Sv1CEBgdBcCRzyy9YSWybqVq6Ncv0Y0fYze9no
6TnAjEGz81vlnnUHx8FKedsK4o1gv9+PNw6sYGM1FNhdYtUC1CjtGH/N7beMBg9d+9a+bjumcnfU
m5dt0DqxqWDYOWsi8F5fvA0YaI04cJJY6YOAVlnb04nzL4GayTXKOm+aKKx7/YFduY87TCt4OJVR
xLFCO+Q7CSjl4Sx9cQbCKYYSxNqYDZ08GjwsbKK7XOg14om3Mc1NnDL9DVDe25iAZw/aP8JpDBDD
bUi8QCfT0EvKYBvcvCE6fGZlKPp1/3VDK51PIF2WB5cvEUdQw/TzRqJtIqFPLQ0uIFR2HyQYCja7
GuZGzDrHhEmDSK1IXXSx65IHGUwwPBhw3z6/0G4Xlarb8lzFCVXkqB/vXkzvjA9OynidcYJ1hmPw
6YaUskpXHPbkeUxMHweaAAHu0HVAjEMAiGFz12mS8q7HMNOtWE4JcKHb3TkQeaYO6yEJhII5UAy2
eJNYxAJ1436JuK5hut8q87ptSpSed6sVYI1ESUh2lHQMP5ZlbDHOwExtxTgPaqAXtf0dd2w9tPZR
tr3OuqB1sBhEJXzs8K8sgz6G0Ge7QWNdmcRoMltH34X0EcGsfa5fgpBVqyvaqGEuNlz1mpp9iIKn
+j6Rr3xRu0DIdA3dlYDr6UQ9dZi6iP6j0/5W804+WQUC+PlErJF+wVFYGSropX/uXlzE/n89v5BL
WoW2Vo+07SH/KXrycX0mtilsaSkOXo6kVzrQCTjJ/loyxDBnfvPTSuQksqiALg9JVkDzud4t8RyN
oLowhxyn+7sntqwJ84u7RJsR4MCJRlNrStoJXlsyduUtS7mn3YTs0yd1amI0+faBxlg9mUOSjJOT
QmwqX38cU/Tzc/zgB4VLpjnw3bGvscorkBHSD/eIlQmR8ic41DrN0x6gSGodJyJgVFuO0PsjqznB
tMEiqUr7YjBrON0aosGa8OgMmb5GT+HIp+YlFL9wlZIw87fQdzZbh6bS9YdY4bMrYkezy/4ySwBg
fULy0PG1CC0V/PeJVNgBtR9Wym77Co+jp3JxWHBWm9X+23wjBBuO+11rMCShO30lgAiBA1aHpxkP
V2smF2UpZYxQkVOrhTASaHGT/309EaR6q7Lz1avJfS/DVgg1tNomK/y3hzxEREasXarFSDsst3o1
23rYVUSO4loqZE04YfXHLxEz7NM8ayaAYVJNvbB1SProppsM0+7kKyBsi7KZBwxCcF0EC+DPGzb6
JFz8ZaRznxhrWAfJwuiXLJX06iJYfA9ZrOiIWEtKteNCwlgCCya6rbjgcqjQ83ihN9IDWpryrjpz
jLTfs/cPXOfqPk1SL/P3EKQZPkC12XfS0/C5FI49Ad/Myno1NvXoKBdXLMpJ3PtTlbqCxv1Fih40
Dk8uifbq1bwa97KiBJUh1vlie4ls5F7RvbOhWwrlvt2Lv8qlHT1/BePkkP9ARxuSfffgHlpaS4uV
ykfHzprIYUU5I5BI72V1hbGQpNZjHwipwE9oCyCZYm4oQRjuuQcfB8Ql2y10WnVnjc6SUXzM585J
qCUTdNSA6E7IrJ7PHEUFYWfklm+S6DynLs9CpjR8SMRp7Oxkxe/eY/05lTEA5NT5+ZNu5nKhDKiu
ISmt2tBy+6cdBuytcftnJkn0w2BL+LH5dPY31+IgikO1PtSlutpR70SP7IwjzrNiK3JnnS8xj8BA
gzYlj+eXbA1EHdTfSIcxz+PvEBd/0PS29MECrQpvevKvQqzj6RceVaVIrd0WzsPI0Qw8rEvL0bUJ
3zL/bz37n3tkotipP59YexmGW+nOyf9Ti9fy+w6EUaBs2AVADnodQwpuQd94wnf0GWx2oRJ46z/G
xIB9NOyeQFecXsZcLQMuUkiXkd/kjVfQnRnGOkj+E+UuwD9UMw5KaA7J2qryaRNbf2I7EitE2tcD
kws/qycHfojnKNQBmajo+lJp67soKsqHlOJDn6hpWkRq0qkD7noIfcu0+zlENfqBh9DbEFllhf8g
vGofhuJ+i0tM/BaPooC1O7TouVKZ3+eHoe0tRV2X+ns6KkT57N0n6XIqpOxh4gzQzjW3L1vI+08o
Ju5Z2TTfv2ZowOBwEvy/n5j5FdgjJeBocxvMvGZfpEpAsmbn9KtgT0e0RYOTxOVEBzchn8Tbv8d1
RIrPe7N3ZGfRSSKjHU3pEyW0zNjfySyc9zodO4DlWynaOQrypAiDmrofdzAXHtskDpmS4Ccz7/4e
ASlMGYUz6RZQv8lH1uXbqM9qPMXsBwwIyFtOzLxYjE79mPlo7rwmzjeBjhr2S7MWtXl6E0vEFrRb
VwCQd/RaK1eh4Cy9qUURdntBY0zsn24kLH3oBfiT7y6UawcAwA6K9ncGeZikTMmmLp5Zg/i0U+aP
p6CsfSbOivQ/S6hv1dlzxvUQHkF7WVias5hWfzHqtQc7ji8SY2EgwCoLnVDJNiSAPvGzveJ6fH/v
OnhpyfVRB5I1JaNeAKghE9XW0dXdnkxBRvZgx6HYHpQYKvHc4scpRvPgWPHqhruUoAriSgqkOtUR
aiuVshNPFNZu7cj5XzMUCwqMJ2+2j7ARAghACU2k9NXrxsh5rPpu6NdhC/Q6QGw2V4bHL56oAD5F
wtYxGjXiFXxPSG7IfIuocqWd3p9BdLZVNjMbYb6q1eka0fiNyvr638wk37yW0lhpG6uTzjYD2RJ6
pLKte7Nijxb4mMqROmMZxLhdBpg3kqfzHeTrFaj3QNvL2nmlf67TeHMlkcuP5nxcnDCMfTvxajjc
9SAYq3ARQNBflTiLjE3Tq7F07ETWa8xiCCMoQY6a7m089hQzgIFJi4JfNUaLe1MIC1nnC9tSg3/K
5TIkb8F43ZRsBdzHQ/ABxtnMWtaDtJTeaZyIZMm3s8zDdfa6ZSmKnh1I0MY9PFnUEssze4pvwKvT
7lcP6dOyEZvXAmAwMrIFhRqMJ1zL+PA1vydWX7h2/LtWbudp6eXrhA3VYLSe8214YKuodIoMDtNq
ZZxABBgtZZe4EAJaIe0eVvlrmeP+fFZdpcS1Xu1qVV2TFw9GTd5Cfe4bMTHJ++oiRicTKs5gKwcD
fzob/7vl8bl9Sq2JG62APNyFmLzwxhB0IphthdOx01RvKKlBYrtd0EosutD+m+xQNDL8c9rwsdHL
viAyiyKUH0/PAcL/she93Z0oVvG1peITUhTH2Xl1bHSfC9Cnoc9HU51U/yuo/lmtfAXOFAjP81CH
0QTyGTnvk76jOraJC4X1xr5Z5or3cvdkKhHuE7W0utX10xMpbzoCgR67As6snaWtUiZjfVnw/K8r
JbfIOYCKCWnBQcmJpZ33Lta/2dtyM1KfKRYS45AkMDSUWdQUM/yfrXD1ICN880Xtv2f0xsCUX+C4
VQH5IA7v/TI+JPoyjHzl33am1XDyBZVrLM0safpKYYRHyys1hTxZvcbj5jEgQ4TVy/o5g9WnUh8H
v8xaogfazPb8YucLrTmtz5iY7BkptO4giKpwmBi6JLxdwLPGbUvo/3PuWozn4AGlddVP7cMfK4L6
udqQ9yGgGq8ducmFd7TvVXGqLTKdSmGpKyjJxdz2MwNjxcHl5JV/+RoUDGSzQ1wv8iQR2Qa94jpk
MilHSxbY2c4gFBa4LUF8/+nsQHanWIN67C5bCiUly+my+NCz36yMzQH0q/6KDvNABnl7HbWX1lS/
oGiHmv46gXA/WWZ6468OIGYFEBD71U4F21HqsuVjcmikx0XmE1OjPP0kkpX6WK96Pjweuzho9SI9
7XMQHrmLqpSMzx2/IzUtrC5Q5oee79cWPV92y8fmG3BdJ0DZ1gzWVy/4ibuSYqPUran3GrWgf4GX
kqvClefCL8tv6+3D+HsrXkM38pycVGJ360b4sCj3mqxk6grkYXjP8P0TOfJ1M3ArPROXWb4nGJI+
qIbncVmgzIGTO4tDldEpWX+V2wZiHA2YO39sqbh53by96z2qzjdCFbsyC69Rjpbm220vHT3kobma
zb7UJC89n/zlSNNlPI+BPtkKq9buWY0FQadRLnlvL+06NqnVTYv6Youezcr4cCo3THts3aOTqnHb
EzYL9lVUN3VUoZnDcwPglPGY3MfnNP0k1BUsU0HF1EgEs4QD2ONn1lGZ+f3c3Lv+cnPRZ4zjdCXX
astmQR6UoXLjIO/HodpyrQ5uK5eDOQEKe4ysTKYBMBZuwxsNE1iNn1am38loCyjrihzestkKTmn7
inTX8Q3Z0MrkY2Ol+EKTfAI2o3WB++taNF6tQEpPnrZpeWZ9tKTitOG5pspTBn1ahNxkVD6nkSJO
aH53bcjzrt1VQrOf3gw4zFMuDd67dnhLXv3o7JqEi6LGstkuTzDOhOdlPvy6hkbTeiIowAtA1Ycy
uFStdH9T3VBWXOuXYBwJE03eq4S7xdxW9S6huNTikWjahklZZOZeVbUUSbE/xe6Kex31SRB8LUcI
sTjgM1C71UxHOupJzA18T1zNKFJmQDoOGTh9XAyt6RdfWbIme3RtSfiZPE6G8odTLFopQHf6+9d4
kIEQSo9zMawA8TAh/h0z0f89jPzoU5V50wOWP/ZZ41Ag7TDuf05+xWXl7Nt3KFD6636e0xQlB2vd
L8WBhY87pM51pz6Q80/M6X2e/HUnyHq8jCZauXmZAxNKtbl7k+FD7Q7KccUZfnIEh5h0A2eLiDMu
hf7TJsPEayDMDMtSowBiYMXbWQZ1+SEocnirGkt+SV6WLExc/iLv5kaig+owUx/25kLeMvQLBV5a
loL7c0cgpvhZcanEtjBQaWsaIMYjxV5sTTqxVVbO5jOixc0b1hybWPKktIOTcxJkMgaUmObkiYFv
CFIKZ6kz3Zo9LtRbG1M5z+vNTHoaidIH2wZVvHLxCP5xecHHYYaIlG9dkSEqmg30NQVt3UTsi0cB
MSDKpN+UZZTEx5WG7WoGnQQ1fwyBlmniZqFy1X5YWTlHaWiIf+tDiQlZrkurjg0uzZLHvhnQgEq4
CNvi6yk+0BCPJAQcw36+X4gEuY0apZvMbaFueJ+ENtk7N62p4WDcN2FFGOcmpDYZQEaZ/jd7Lw8B
zqggd7hLABwm3Mgl27jLYpa+aPzO4adsVil8WAVCN9oEsX0TfEQ/t2GjR1AQDOdyD6Jbb0WYHgF/
All3C8037bv9NSvyVN9ur7Dhgc+IQs3NO/QJZhs+1huLSXrd2QHnTd+KwRZ7RBTXApwStVv4YO5D
pOCqjAixDsEIf52p+E1Sy8YKMH6yPLE5z2QmvoCnIcaMRkAzEErEBlqmhR3Xc1HLHTV9366RQ7Du
HeFUCZISLpfes4LYbJawU6zGn9kv6wan6sMXtkzEmUAIQXfUrMt2761YTDNnXZzO3wBU6fY+5o4w
KZDpZ0Qb1WkYUjd5AC+OL8glmcN6bc+mWZUQrcVwYK4CCHZQiJdQgUtwTRYqDExMgnmhRo4swP6g
gZJp010z+BeDOpewljAfEGxEGFzj5E/kqfd+dE4K3mqj3qcI0CUnO6VjXc94sNEw84SfA7BPaETC
ttrycjPMv6um72oLEV7dgcaTFa5zm34tATO1m5GoLp7NVWL4eSEEAp1Y5ntx1Qb2Fov2zJP+gB85
3A5iwcIZtW331NzolDA38DX57FQbTJmQQw9xssArIbZ9G4hccDw3ej5D2q6xNzrEWg0AtaaCooyw
c+deZGmR2NzMBVwhMqTy7SCRnVhFrn8eNG20NAPinEwI2OQgeBC4djy/hpwfQ2FhLXO+F5YH7/tv
4X5batQ2ni2szFtU13ZhKteMa+/zyE91sEyEwgshNxJKsGw/V0iTH0SXjQ71/limdwWszBOMr0El
0/atr46NAJ26bwNTAsHGfaY18dYINJSd9Muz4yijHfmLx5xaOq1oy/NhCR/2YqEqDq56RHd4CeH9
5VWRxPdWP7TUm3s6PmBDSIAMw/pgtm9+iI8PvPbyVb2wlg/5uFVVWeQASQSq1TsR5DrKnRET1XCT
UD1xX4DbR08lu3OMJvbU0p4ivxgp714nAtgZ80YSUsDqvOhIaoTtnYyfUacUQCxMji4QKmzAYkVf
N1nxSRFr9dptqn0SP7Wua65d3TttCBsgjEReuJmPj3vF703j/5sd7mHZnsQgCp+JKvxjtlaEpXR3
+zAmenn7HCgqqIVHElkruOVUzeK/BVS1UvbEblWqC+mgggn4e3tFXbzeVwgKMQGRuos9kDTOPGYn
sGDUXumanKwCJh3bm3YfJuaHXzA0x8mDzX8onGqGDoiXrv0lSmu97dgo70gdgeEYdP5pVu55EvoU
DsbG32p1GMYUmH9pc3AdVKxHoqUyKSRx94DxAqZVsAtw7Mt2aIKLleDVke/cU4COhrbsRNV7U62t
m8yiM86A5p4gs6T4+JQuU1aNaha9LHpPLIWqkras1w1CppTNVhEdAR/3+5DXCQ+O3h6tPiYAPaSn
Y+aSlGq2NCHoYEHUGBquMeDbRYrNIYG+rOfwdrpW5UrnFRNxV8nstHPZ+5HPBxhOK/X9pIJY1PpN
Tcf7TjE7VdRvezcUbAEDwC3kyCYWUcYE4Lq4mWvuXmvtSZRl7ycr1vt3XCpIvHh4Vm9g+gyPAofO
xwymU2xhm/b79IL9KCLdxTl6kixA50V+bx5EtrZXnwvvJV3tVG0dV4Kr0Pw3yZ9BiTiwZlR0FyjI
ao9NixN8TgUNvghtC6A9Z0NnNTCNUXohp/Xn7rmGAqOb2+R8K0QOstn3iKoYeAMT7PylE4omLLgA
jqsLxV251oCaNexJ4ZeQbQ92g4AkjRqzEnsAe54MViaxh8PIw0uBCbK/ex0aFJQLUpe4Bh+xA0kZ
8TBrUX5GG5OLTWw0VeISxZ8joZTCf27qQa5PjDn1WIdMDZwCXIFjN3vpKFCCC+XVKVBFpXb6tDc+
t3w9jBrWCzFfNGXUZQvlt8cfole6OGW+EaLS4sna8PXEC2rBHABBaX8A2Md7JB4M2pAx0f5cWzpy
bs2X5VQo3CylZhTtRlxPzhQXLgoXAUzZQNzj8Lx4Un6RK4Be10EpaKNuSfqjDtMcCM5BaARvzBmC
EAROGSLRi4x+nQ1q8G30ATnwRxxkfyCV2UinMDefAGWKtYLb+63+6VF17prmig9JCsLRqP197kRC
BMTV8TDxfzh8ILM5qwHE2fjiaDhJff2I6tTNXKT8zY8SZeucf+ThMw1+c6MrTK6ncHtcSC0quQXx
deJys56NZ0PxvvpjgpLYg8zBiG+zOElSNKHKuGnm/rKIvP/opUTfqEZ7KgGdNqqOHcrxjbco3dzf
LFLsUHuD2/OrFT9p/4r5SpUKUpTXen/FSRzCF5fEucZDg/nnx9nnnPIMZpkL5FO/F4IilZAZM+qV
mpM3XDtBaEvwSAKYM+Syr093YJILOTJrb/L1h9fpnw2SuZp+AF+A5EyJmNDnc9SM5Y8ca4Uo0LAa
4MxPJTKKnwdcQEuZs+ZiflEOsYJOajlX4GK0g6ogyyl1TIo+E1HYfkOnI7JS5Arywu1dz7wP99Zm
p6NghCyZ8bLbLEyEI0A2x6fGXowgw2opBsa8edm5ECC1/b/U2Sj3OdPo1kE7AQnvTTxotAUKN4ju
oNfcLdoFSiKUBJhxyifcSGExt6L+yVb/Zen+U/R3BBIAsFD58qRD9Cpr+98wJ1sq2+XNWQSzIJ5c
XvLmAc+D7qdlk/gFuRF/3V+KSPfoJq7I8XHH6l+rtByJ15nrhfXIBT0v2VMKJsNke/Nn3APakQUI
IjHb9Ri5UzmXSO367HivSi0f1R3UCFu+7T1M6slF3m3WcPKAqP0uEVkiArvordM74VNbkuL24gNq
h43MKdl/Pw2ZWHR51EmLZYGlRvp44YwFPilTGYv6Qmy5oOuLy7XQXDO2p0elVcWWbnYpblwIe2NC
T6sBZ4rjwwIgGZ6a5pAayX5/XlWSShBTkbGG8qf4oHn/WzM7itmZcGZ9Gk36msHMzqY2g0XGQCAZ
ldEExqmXAoMPg+utVxRZ0cesAXgAfPqxcNuIVJ+tVSYyw1MKLqRbWrvmcyu2cTO+OKOCrE96uRWn
AfeUKP75jMBA5OL491cyg19jc7aYls9A655uLU2DcVtgI4HzvZm+ZDWOukQM9pJE9qgNFqaXp+j3
bEQI9PKlFfb66kDolADOu3t28JlPl9IBVu3a50iZ0EG3CZKoYsZ0aG3ScFNP9LkKKU/X+eOPN4h3
tqTy3ydd4i+BI6Wr9bgxFxJZCwTMN2Z5EA59hFCCFZLl1zeMdlba9CfakJBeNfbL0I9Ajrv6LMAI
DVy+UUIuplM7eoNPIRN4ST9XzHEjaQ+gZc/nZwIk+/sUnxfeJyQrYMPLu88bZQuajMAmZw415DsS
RgWwuKuIru/FAoqdLAWVRd+8ztc6/HXBEnnAPQu8vaCF9Fqp/EtSTejqxiU7A4w+LuxRnA/zmgl8
gYNgDTBNA378ryHt+Dq3pbeF0HEx/xaYFuRshizDywR3YwUVZvG4KjrWgiiLEtH/D2pjLAVsZX8I
mrQJnk1eAsyM9yvy0qeRuufPVOqUVOduQI3N0E4kod5ztdmZyVOTrjfIGp3ZbMbo45dmJ3521P3j
fau/Q4LMnCKhUFWLXBAm2l5fOXeIWWAAUUF335FHrPZVRXeQdKNtlZIOL+H8qTdaVjWlhO6Dnthw
23L4uxa3YKlPx6tQL/FroJEyQ7ujJX3oJBLxX3e3PfWmhdtZD+p8VHLuALePwhUQ0OUaykp6L1k9
KONMAmtFPGE4jgx988UJZy3tnMsjrRTtCg3gf+wrish3WYPMFtQlo9vcMByEjRkpAZyT7hrwcLr4
G+0vTIUhdsFasHTbZqKMNihouRNKVWmMRYxHbFqQVT8GdZjUcrwWfTN3xKF5IK9KnJvCboEkml6r
L/USxaAPDQKoufU0/lSkNmXFBdiMxAKEKl6enxFUT+/fKgHCBrFPwu+346ctW89cn5ishsv3imKq
yH5MPgQ/sn9Q4ok8NEsFXzC0QdndxbuOwaEydTaoPFpn7OL7lDAVIA7+SjrKhcb8VpSYeepoVG0n
bxfwZ022dOZjZj785AuO4W10eftZ+4qUriOecXMJ0wzOHv5fUrUm6hzE6o7ZJt/4duaH/lKvcCQk
car0wjOUumv4ar7SZqJExCub4+P23bI7/eg2mGux12CL78aDBIJE25LoSmmuF7dRwGU/qImDgWH0
nYnOnKd4/MUwFM7yKnw0kqmrmeg8coVW3hB0URlYhmfW+kV3uj4RDBxSFz9YnwedZ8U/Lt1zDnVo
kN/HqwsuWoyWzjf3RsuvOCnS+LXo5OajtKj05J2iabpDNZNqXl9EwXkUUxA+UZn6LwMxXTgoY9LB
yiYgu3Nj8sR8GkVZ+QHOz5ccvkDPLLAAoSvmmgkoQ8nucJTz5/m0uyOE/eU4QVHkxkm1fri85rkW
2kPg4kkc/5nD9gy79KyEcnq/ZBsB0qqVs0fnV3e+nTmW+U3j8xUlDm5Gzu9+ZMZ3tabZIm602DoJ
tW3lFR4GvYRfswbIY6vGr52O0NH2SuIctjw6lt6H1QP3IfPh/Qc9eLFZMQoBHkQOZ26UqgpFJT2f
/b3HMsQwq5NfbsFbZ/ktuLEvGGDsOpKAtAgk6rkFehjvxMSHnpc5H7ap7pkeX8RdM1c9YHPvRtGr
2nlbdMxQ7opxxda9XmXXicPuIY9Fvxl4PwYwYh0DhxGeb6HEx/9tf9ksbjs3pOzFeIJ5i9C6h1sp
wqMmxDFY/j7jBlwOGtdaDBUeELZKzbnsQKQbGZ5UMTszE2j1FcCHbuQ9UZLWEyubeu9de1K4nE0U
Z8n2hAc5n0cIJot3t2yBkVuYv68qFxo1Ls6QZIBGBmTC0oPo8HJgsc8OLD3Zi51pGIyQtzW7ikzy
X95cJrowjHnpIuubMF/zdQbFiMml2maXmzUd3JhtuTOumqs++QXOucJec08lf4YHrpkfHmN6+FrC
SFeyiCU/lk7d1FNrx17TMK0ESEJkybjWQ0ZM9iC4q24dn5kyjob3Mc0XAUcLSmoKfjG7AibPc7RL
c3lB/1Xim3Nyb8Vu2ui5YNaT1Q3+z+L7Z6rH+JNCnr/1Q8yXN5NYR3V3KjjtRYX5QBPFdclOrRZF
aI3hpTApYZQOBJiPPhfyRQLG8DdA39u85dJ1myiA9X+fZQtpo2wy+hOqjggeI+RBY3SeXhlcs9T6
579OpdMCnsZNCMqtO887fHN2CGeHyb5xDEi3aHuO5zS/YBqymGdB6Mz1IpSN79rocFCcucsT9EUG
d0DmtxKqL8HpJlo7kVeKjEINM22v8sXD1/bUICo1osrKWhbIGNJo+A8IhyO02NOy0aAaJRrs/kON
mCH7sN5CsdFNNqq9JAxoXFt9adjyuvPVwfMXG2F85nFJS+9j2tH1tHy8qnkxsX8XlOWj9CI/A6S5
PJPybbdivewf/NPfo2yEJCTcCvi4Rd+CpR8xnF8mEJTwBvegnaC+8QMbgZ+PRJHQS9UYa9Ud9+Da
vSB+ByB4tmRc/Zwou0uH7M1warSsX9fhNrpsW2pBim7dVsdwABUdseOc7YUCSAk+XZjluxpYdO2H
YF2tiaQ7Ao4GciPjAg0mnojWsW6aO0vg2Y0bmj47RWDM6Ds1s73Js5VahSGjVpdNFADc+rAymy8B
DeapHFAF++aUkEbx9t5DxA3cy6+ul5bhF7zMj3PtY2hnGOpzX6mA/LY57vrwKI3t/GFGY3VGELW0
A1NueG0k90NzD6fkzLDCU1V9O99oLqiV87xcNUf0D64sm/T9DWsYMbe3PUq0VtiGKfiHr0RTMGFX
kSLCon//Iy5mG1p9E2rSVUq2seG+nPxrLuvRd5RdiD5reHTUJZnmZ9I64XJKFRT4vv3f+1A/Vm4Q
MQja7e5fMP10NSOrjV6W8yY1rn3PwcUpFMAyyBhmWrcqyFqoSW41FuwvvpzSEwrgvlEgirp7AtoN
QQFpn3NdPsMfDuUl8//Y5r94EECulkriQjQ7KdAl6kB+QZNlTyxJ7DuQbW33ATwIFBvVR5tellrn
1uzmWaK0479HtlEUveyhGiJO8gn/xMBevaYI/T0vhRFMKsjKZwhcUaYPbTexA3Tc2w1TdmWtINzJ
PHIJ6DGy02bQRJ+I2h9Y3VJUITB2DMAs3T22Q3idh98F26Di3uPXEJ8JJm1xe1hd78KfjqHk5KE6
MmdbTLKa9oIdAyGGD1AV/XO/jLK+xLSzPFX6RmQQSaMYnyK8/dAPNY5xS64I/h52lGLItuQ+uAc5
tJq1xbJyLd2UD8+0/W1GcJ/o/fI96e9hXSxU2sMZTyPgOc7oTw0NK6wNsNWHPMRr9RQTULV6kymc
VYPneIIESdHWf1Rv4XZ8NQgHLDxTbfJZCgQuIrH3QUkA5m736Ag1B28CqUgB48fpC+P8N+Bthwfp
DR04B4TvrlnvJGKeSOPLBghJFhmc/7IwfVbVYO7vkjA34hf8j5ja9Vb6qVf1oabvEzdJvfvQ4A1p
e1r4oO0eSOGRlUjCBRqV+wwYRhJWlu8z/gpPQFP08MzJiht1FukX/xmB519WSX9YFWr8EWwLF2Fj
B3a0VYjvbxwT4UAG71fvyIMXFlf1OzFJCmIxVamqwiAFyQuHvEOh6znqPzBgp4ypTb6Vi+c5sGLK
mvWG9+ovTRV1NNbdBgRqs56anfB0OCcPw+5e/dIE6G6V0J/5bTpknf/3lsgaGvIvWleMuttWmvUf
rkcDjHeqjGSY0XYZK5BrbsZjW8fyPtOmFaqMAfm7893AfyuV9jL6aNIXxlyBMKeCbn1e2QhhPajU
hSuCLDhqA7y3JajqTl9HHGSQtoaMYNJQlc2qZLKPd6HUmYBHe1cLbCw7M/yK+Hv1TNnmuYR8dBBc
csJ2qd/HDXqttF1acnmAyqBbYKU2kOriBEdGiO1dFT2cBD5/Sfbd8Tf50CQHNOqieFI59GbPn75v
T6v7Ey4/cn3qUfM7rPk8l2vpkq6GDLfiO/e4bRTmiPU95rJr3UtQ1wR7FUc85qcOZb7WNSjCAA2G
A5eFuBgL7zm0KFNzZiSb2zXzo59WMSxkCrlB3OKHn735ACG6bBkb19qJI6CAveWzOdhNCNP2dLLi
ncVoxf0X6ELzs7bNt5JZN29EKKOOM3+p2eLQJk028uICK/EYoyvI/cT1bWWEHAG2JZxDqAEYWYfF
Mm5mg4+VVKiH7G7V0fTs5YsNVewkHtvEB1i5QqUQ2pwWGmNV+N0obzQuyS/zYEp4TmB/AAJHoWbn
DTIPOcAI810ijZ5PmCy2uX7wdcImatDY7NwwuixZlMyHZafTyMpaITVJsKVva/XoRctHYmoHTWu8
xwR0rKOcK9BrbV51gHWScMy+xKcfyajMVGAR45XBSy4BzlLxNmeoK9kPIf34f+gnWxpGAzx5uJM6
Y0V11al5QAGkIn+z573tlkXi6PxYiqA1xN0i2ixs1ysOnIZfyHBlLw8hHM2hNnonQW0UFDeHAf+l
qdOMe7j5q9PP8L8+ymurRXT4iy9Uas5ws9pVB56cGSZNTbbbx9nAPcV2ZUyr7inKKjqEEpwSbvn4
ylzt3yyZqSCPvs1x9mHgxLiZsKb4qHurRcgCQxaVJ1m7XuBdkaSR3mZbq+Nw9NFAM39rZhxXER2U
agPatkAZSpam2l57OlYSdOFEGCm8TNaUP0RMSJB7HpLJjQ8Pk3uVwJPe0kX77v72Y3jlCs7j9L63
7v/fX0mRbxZZMnfdeLS5FU7QEKoQHdhnBaae10yyi9qIx2AQyPL6IrY0hf7OQ7anlL5yBOVasfkK
4sQTy+tdBV0+Fl/vD6vAiB3CoFtlMllonYBzkOfeqdNGgEzd8W2aJ/EX2up8AHsakC3vGgQMAa9K
XvcWgKBCiVvQmqoB/Vuc10VXmqRr6rcYZteHIcpFsXkLECVpYqHVxJjvvcymEU5qpTWjOgbgCVx/
e+iDlibNIrvH14sammS7Bkayg980qAhyL0taLk37HQndC7xClgb2Yfi3vizZn56Qo9yQZvFOmj40
Nu6YTv22Xw4IKX8dQ4ONYe0TyUGVyas1JT7xU2etZCtkImeVKfRZrsW6iI5cOwdujmfXgwHFowvN
het9FllBV7lGg13l7w/TO7CwgVdeWRsfl4Q7II5TbHufA9uY3+ZsektXjM8FHdFA4oXzplGX6czh
Gdsi2+eoUjZlrFk+073aJLHO5JaWncOOKqno2JrDuwHTQJVTBSRWZ1xs7+YJYOcWgM2/nOKHKixw
zamRWq+nDqijeidiftFfZrmL3gh2O9ROhdu0dOExp/7iQsYoXeCQxg6d8QsEZDR+pPI61UwnPa0e
dwzEnNiYlOuubYH3w0SycSiZL8eX/TFeLK6xw5xkuuEZD4SGT2nuzoum3oryAZIrJ/3R0n4ho9iy
obJHWEZoPotPwjs2uJ5alWca+Sj1fscyFLX5y9ma3OQKO8AWxEZDlf5HrdnnY6rCr3LbeuBDiO0V
vKGD5k4C8lIj41inXNR1Z26yOmcBuINPClUvbx7a1x/YHqKTEZebj3NvvwtoBoAKVhsp1GU779Sy
AJg8QXEZDA3YqeyEEkgIq6XOBY7BzjtodhljOXJdab2X0FnH27y5AWg7qx2VwRAESOOYAyn/qngm
NrdlNWtBbhSGw4Njl8zhejOHs3pZnb91FDxM3CvyYtmQ6+uwX0PYrf9skzD2JXxnFbSPdC88U2z2
hp8Lyf14HPmBmx/GGR8rVQ35ix9ROQFM2ckyQ0Y1Rmk8EVAaZ9bC7FiJ5iN6odj3/WCckmfrLeZH
JFp1upuA6ATIHSPJ0rEdUfN/PG3jzt5YlM5d1eazYyv4p3MwqQccqhUK4re7ik/lhOdTf+Ki3cLl
POYmQZpRU39FAdGBK7tepsxVXEQ+hw/21O/JmY7tXKzRrrQNczvHDNNJPlB+UNqIQKFwQA9YaRUF
muza78i5DeCm1xaigzWKsLBxiVBaz5lcwslw/D9eb9SemzZuLWw5vfT70PXuaPkeqkXpMktI77ra
SUa/E8td5/4YoSVIo03Wfqd9lEj7BV9WexPfC19nGBWPKv2XP5rp0xvyarubjBvUPY4tRendKCHy
MLhKLGUFlgVPAk3HjGFVmZFxnq3LpsCBp5xOsXfJtPp1YS/3J9N0L14EzEPHPAmaUscevyoc2nzE
2DUbRza6lkyBM/M34p86w+0KXCFxqCVVF5/XmSsL7fyVGhFWPrNgDW+arqtPO0BfRzhgwaCAqppx
7j1UjyTA3/UsRcZPDOBtSweTkgo1xkCbBBReza6tCVezIXLl4Rds6/0pMZ41mCIXzGB+wulhxFXH
oODS4LuvNx4uub/2ZJ4DAPrdp1QDw03syLi+6hI2EfYbLJJLDnIRdDYz6Ex2Z706hpTnEXctBNCM
Yela37O/G/OVW0aR9gwed2zONL2USbZKmjUqScMkkrqXqBbpou3F3mYyiC2OgMXJh64dsS5PxxOo
Jl/vAvLkOuJ+uIqsfA+J9uI4Xg+2pTJxHxy1/pj94IoVpSqE2k7W0zBA337JWa8H/l8zgsBZpqxR
81rF75c+UBPYgeA15ZmNMoxXFq6rO23JtumvhewD9DqMDBrMFQJLSkQ7JhDZQUsqUVVVF+xUqh4z
nMI2YN8QPeLXlYK6TWxIObLSfkpph8oxDRzReI30ixpD1RDh3F2c2T/BulIhF6WVbLYJ1aIY/Cdh
sfUGT/rcPmViBKOr+ynAlmHvMJ71ocqRKN+d3ag7YXpgmxW6NK2PeAuAv9whcpejXc9YrMjKjz+t
TUFWnpz7CVlGiQe3jLVvaCfqmB81KnKSS/7MNhn9s0gllsICWzTRSd2PG2jVcWB5q7Zk+6ytAA4J
2YXI27OhKGjZl8XXGJoKnWqvIZs1zl4985zYL3chMC27v8G7SLs69PH73de1eOyr67uYY7oxp1wj
Yz73uVrFJx/G4+WO+oy1PgAFDXitmJ+nv0Ar9px0n6cM5fjtK541xzo/oqetLcVXeyrKjHnhSIcK
n5G2iMcqiBDxK4/LOOljYXKP1oUmbQsTZWkBPqxoYuCc2UPsbS5+6Mn7iMWX1gZpsfT1ruszk6Xe
iV6BVtGOF2dTNFEZtO7CzwxTUW1YClRLwdTq4dBSd3EhbhI6dN+kd3PH6txd1bsslEYS7m35Bl1W
NOJqFzB0v3tzWWYfXeh9+fNh/Lhu8HJrzCUIgjP0eySx8XHRsgYbNF6ZcmAiqGHvQg28REqqmq3z
UlPG0R+rwz+sFDqtU/h6Kev5VX+338v2vl+pldP3BOpszKxdgP/af+qjvb/RBxuioiqCTDBsLeel
q4gY0LwElY7wJQiyBVOpjki1d5+DH++Iq4NCvG0UrHTY0yAJOufqirrf0h9SMqvxESjHzWVTqHU8
zc9s3r+b2p3lqBNY6hvcXKELgkbe979cUUI/XmoQeHSqqVJJdkDVi5Ez7ojPlgrlV01as8By3JEQ
MjeEuA4JqSqqWew9Z5/bqucaWi7TknymaF8gyJJpzhwxp8QgCXLVklDXcQdqcKneDNAJlwghFQr/
kD0jENdVDoBYUxQpSQw/9TnYkLogx5NxaAyzu0oM9PbYUxa+/D5iTJ5A7z17lXr6vxQJJ5pkbhZO
hpwUO1qHkmBtRA34d0JR3Bxij7cB0Git6t7m5Z9X8ror5vnzwzhioNSvLtDDMl+3gylv5RxsnI9N
YT344A/KK68qK4u+2SKYvE++CROnpljhUlNm63La8nnAn5osz5EK/b9YYY7sdQD2W4gIzViVPW3i
NFI88uC+fs+iuuDQdUw+JMl+hh/c+cCJTYlfWEhAvPRx5+JyCav4Zs1O9D1CCpKDjly0JsY0jRt+
e7FUBmw3+Ave7rwkWfxO8axBCco9IM+6oUPNOAy9bofqAbiMBv9FhkKjBM2FPeFeQtt0sKBOo6Lt
b3GC9lFKiYCM58AvSQjKoZidW7+CUNXAEEcqxYU5hYOLDzLibgxfcbhdLArRLTRMxgKEDYtVSdBD
ZmUSdPWALRTexD1cBCfOGADP+/aQtAe9tbZvIH61yTZZjZeR6+m5fGNzIxgzw1hZeLs0MV54UD0E
msRxZb8gNpbtXX/Y+zpz/bixGO5eJ8yVHyZCW9svr3S9Ds95U9YuskTrNe/HbVs1l3BeAStyiuDw
t/Zf+qydg0UGwEIOp4dU0o5Kt2Yj9emFlWOICIqeP+wriwQNG+QF6vwMyWHRq8NwGgHCL8vq62uX
zBp/3mAQRwco9bKjs6EW669Sy4HesgaQQTJWGWLjSVemQWSLMlMwsECFt/wunTK77vWb2KqCpwJQ
WLWW6SBaCBss13Lb7QszXLYr9T/+tWAKy+/+ta0m3kEfDMXrFKK5xe4q6doMSQGEU8g0ewHZxQtm
H5+sUo75BxbNdOAAme+bWa0pzWGm0EG7kNLCqCPAvtGOaYjJ5cKBe503X+1uwREdCs64oxMoQXLx
8+c6DgmF+Z3WdKRDAtstwcIgrlc2VyAjnH61S5Ez5RPzKN3O6bGDdVPqTb7NTyaarGYz6QHbAOtO
wssxQ6B7kCsI2LI1fMjpio5wdRqdWO3GFhmxRZCQBiy7/Ijvw2EW/ugvKTFvqMBsvwTYO5Um7PFn
ZIiE8AETtN8yT0eYV+vRYPAL+4MraUJLI6JO7HiFsuBYMGWN31bjeb3fLD2qPwF3UXrGvbi1+3zY
Q7hI1J1uaw1ePg0xnUR1L+OL4a8y6UqqsuGyLaIHfzoA8pxRHWMv3UiWk+W5XY/YAnA+kSAcb27t
PM56P4bogntKP+bKY7FmL5K+Ajg45TTWCgl2XWmgZi/KeMec+2fFFxUYk4BKsgb7BC3kDYhBXIrt
bNgAvCFJH46X8GopJZNcCDzi+Dycu7WAiKRVSwj6PXnXy7tcOw+BIgldb1gm7ck2KeQ+pa/vZZl0
KfTCZeAZXfeo4TsxAMwVlPjd2GB3PBqnJIZAnRzBS1icY+Dwsk2arQR1wgpqO0QKJdkIUhxVRXm6
rQCU7lY/LFVyQDZS6A7eDN55n6w6Afj1cflgZH1VY7btHYBYSF3O8G54iL4ubpugBQPTTNVXjCt6
wuLfU1a7rpFmScUqrHLFvzzCjbmNeWFMLB1jOdzQqU0rcF3fUXQEqU14UIUEsZYAJ+PCw6QJo5wP
ONqhiuvObjGLMVj3o+xPOB+IjrYIUARwlAeykcfkD45jO1wDcGDkaeTTFDzMt8w8ar05UCAuP1hx
Val9rUW84UcEJsCF1oHj5FfxNvElX94BpA0EwPvk+P19vM+5sF4PDLFB6xTpViASvmiQElZipwEo
C2IwmXWSbHLazBqk7CgPTn8HUroJH1RKPoy96l6+/Y+3S6dEWnYkSUapvWA7oq2nF2yXgxdQBvxQ
fbePEdjc3RVNOu4QpS3EDlVcorIRVYhQ6Zgd0acJGqsTLiB92eERZDz9P3y5LToNlYNXrGa843Jj
iDEF2glCktYcbZqIbjlX1R+LDV0V1uVJQoSNKJeSO9l5pSHSoaNUm7dgDdbGR7aRCgjLEEjtgv84
03I7RXKSxMUS68FFQdp+i7xczrAZqp+jrEee46epTVdDMWnOko5RpWOpBDsep4friPqZsug5L60n
fX13uDX4GDEWAHqnIRrkovWW623toEOHxZcSSI/WMBliTTif32rOV6GAHYAu6skqeXaqSeJ9tiBA
0REiPFCTfI6uCbKuh1o+1/PyfujtBJftG4RCMfDHzjpOwgfkessGPxevE8k/UslirgC44EwB9sp0
LAsRoT4lZsHdBblsK3DMUm9MFxlCwuPdk1cuWgIZXqdPidKFMMm3VynFuukGU1r+/lwjKJx8cwz+
hNbrV1OISlG8zgmA8kTjKc56605DQiuIzovV1ovSy/EzF6GuKpVGL9/sqAkw2lz9vBp91x47K1Cw
WDVrlPZ8hiO8Cf3bGEZs3lILjwIoobGLZk5oRvE5oucrEXyJ/uP0MV+WHdv4ZkIzAgDpzRaumYV2
idYAeT/zoSC+pCdi1j5E8WdLiEhPxTrQfyTxWmMnlPnYdyztubQDH2Fym45gyQy+x2kyp4NMXGKx
YQRDTFcmykTGMrfoBSGRqc8vQh46RnneVx5jopHyuNCkMzFJujr76WBoGb2eHlJKXZzX+zeQ+aOt
fET6n4pk/zonjNxjFcSbMsYWbD1+bQh+Zet9ifCrE7+8KZwvqExf0O02HJiKghiR5F9R3KmF63rw
dAFLKVACyKdNulEDQJeVjP+d5deJgTUf3AywHlovkvFvyVKTR4sD95oGzk+skBmUt787l5Y26WZg
KctelE00j6LoNZ+5gcYTx8boAlqigKR5vslOD+4WaXtRpt749XXOEzZnWZmLVVKBW5h9IVPP1Tdc
gAhYicYMOujWLz7+aabjWtS93DysX2OUdSJMFOlX9d/KZL58HxkM8MV53uMIxqovFPGnHw0UdrHD
n+iSg5prezSFVDANCRsFRS3hu2DBQx+7dx2ufm4J2Hgt49WXP7ZM2pkNiUInLAQAmfeB/crcjKgW
gkBGJxYtmj3c8sEikRwxKRKU3QmYt1n2NzeqUnUWK3xayEL8an+Dn4m+Toq29rZj2e2VjQwGKybz
zTnhLZIVvBhMqEWmPdDx1nR3pogPg11gddZXQ/dCOHXvDgTlvkxKIQwL21X8S+d23qGf5aO++vI2
lD/b/Y/YzDetIL/Mk+VuYAxDmIFpbbmoDhHav6rZ/GAE1RuS4z+fwTNHYbDIJYGrS+/RPdLCx8lo
FBJ6kx+EnTY4FMT7PEXx4E+LOC/GTgzRTsnlvBwueirfUIBUVyzNo+1VE6eWEd3ez53exIyncSfG
WmBCQ0ovGsQryhacv6HHnqqAExRY98yM7ph6FsHIl9sOnZFtMvzvMQYVfpo61+nJv/LxEa0Ys22/
GFADTX8DCwgFArH8Ka6IyeCQCXbzPWdjKZ0jtFKiwqZ1dxN07ash6ujYFOj9gquvTywnTj8vqsLq
bBf9dPG+TyJNG3AllsQ6kVB6w/OJgdqSoy43qb06etJuKgwxjgDOkQBjXwoda1DRW2xx+uaWCVTd
M2MI/EWF5snJcJTXTJEbQr0onqcd7tQPt9QW822di0yBfjkwgMQM3J+hxXJ1OA7t8lFdTjd86u59
04LIBnHFFFkVzjDLcOCNpzYDrJ08cTbU/A3TJHjpNeYov2fFkWmbvoBXBNuBh+Z43YHaxUIQ6RcS
iUsD9+G9bbWKyFFB858Jrt6I2H9sBQM+T+Ma7wTiEro4DYoGSk78gFrAtiW1rP3r5mOKcoWuEN/Y
wRqRdJNMj2qIrmjK3UQf/PF9rjmHdD56PzaHmSdMvRxZ+QBYjqGvf9kM9siUET/+vwqix1Pgzixl
7FKonr5wTynyGc+Hj8xhpl+wbEA9YiBdsxqkE2Rj6LgffdlzWYz8TpeWq4QhKYAv3BZ4vC1oxikc
C9LOpyvKLRCM0C/qQZhpl8ktsJicCKMYsaSVjPxp5TRzEEn/LBC4uFZ5Gno3aSKnPG+loNlQhry6
rfDJxhtnBIP9jLqZIwzBjMYaeQ8iMkHI2i0YwgpK24yBNbb0sTeoIHl05i1JqXlhvga8d26OT9+T
MuBNwsaS0QmuhsBvC+efI/njsSnE7k5njwi3gLKVtRmiZSRXv4uOcBw8HPxgUWbVS/cQz4juj4+W
8ptmXOSEsEMri6gKnwUcBukMqMvDnr9CRgiYVBC9LkYaIzLrKYFe5j0zGw6d1p/swLuwEhwxQjR+
ZGkIlV0VQfdz3x8R+lDWeOBj4lFtNSlXVVCM3BpyoToqvBEusNzkk/mCCWgFgs+xN0/p/A1OwwdG
gBBdnKYPhWMlVn6mCWJjgxMxfVHzRP/V+YLgWPjFZekhbcaf9SetcL1Vn7Xxx2MZ9gKK/QGdEVTF
AkC4glZtycyXN4QzzvgvYNHKj6yzTFKaYO44HXGUkVCd0vJXJlu8PAiIF4eydZI0DP3scOXmYdhU
eUhsBVWJdgvpKiH6KL75YN/SyRAs/pSVO2P5mczyJCGlk2/Cw7lC8tT0SERIm1RV/5JYXSc4BtIg
TJLNHTDrTq7/ExqeQCdgQnOYeTksIkDB+A5KpAURt/hQwZzwX0qDZueYg29fsi6r0PFl2hud6Xlh
n12XCojsuSj+HXn7Dg+zXO00VqLRGFyEs63FiMVl528Mu0iOauVPt+Qvgi2k3E4RVuLOM2a1WPQr
HQ0ATVEycE/hPLftPpT6Q0WwCT9YYtB9hW2xyeboorvyO3TRShoqbRfjmAIaQm3ZQ7qQ4E2MB5ar
xaKhQO7EzPnSVKfAge9JwRFr/TgeqFfV9lBHKmhN2E6Or/NZF79/6/slvA8dN0miN0euVGeUgNXQ
PGhImhB17Ay7oeVb8EnC/u6usfMffut5ADNZoUxzxR5wB/vayVrbIu4ss79d6VZq4Wk+rrrzPB03
69h9Ky6bn5eM83/4fYDy9cfwCqZixGMNVQGQKGI0JuW7fhE6fuKDkNU/xcC/UzD0DS6Q/jjTalTP
S/4oBKLNd/mhF6n5eHaWKu4buTgZjPfPlbIdKWj8H7IKPNw3DEmoDQm1X3IJStIii5nQ8Ne6LB1E
uvk/BIgIxV+QEBuNTqbvy6iB9IGgVVdYjOX5CwvENSGRdwzpy+bF41bgojPJl08W1K2tlz4yOOkh
mtJXE7dLd+VaaJiNTvxIoXcKZC7iEh03unvZWgTNizn7esfc8bCqhaskra+5ypLYFMwofCFgffuO
+9rYOm5VjasJG+0b8kqxx5O3piI/zpCDyqUamHdsU16YLw1P/1FnwCxXtqOCe9Sg+MXDoaHh/8ui
Qil65yPFBRxRhVRCjLWpJBBJEBxYM4pBPVPEisofOZGaFCymrXFp9gHKGXd6M3lBwXS+YxmwA71L
5aBOAHppG+fJckD9UhCHiV7WVwd2JXhMnvw3hb9Wn05YMTHokF/ea6Z91FP1O5dU/IoaZvwGpeHC
2W+9UJIQmxw8EJ5ft5FxMdWO9jg+cD15U7FRjEHlVnNeM0cAWrn5sBYjFQpOhmMG5Z++v+tb+96q
9tsNq7Okw5JHFmTJ0eSlp+GO1KRKDUNmvWrw6uOmPtLRmsOh6ZkZIZ/3mUE52ysY/8zgfKqVPqBi
hMxKN2FrFs5Y3I7ovAg/35Le3FEGNmFG8xGq8T06Rhr4acxP5U7bIcx0T6A9+SZeKii7CYb503uY
by2/2Bq2IjtmXW6DOrCne4w2sKXzcG721xc3ulKvQ710h38i+KyBfU2LZ/UN/iVmXqQHRJTqGpLB
dnTs6TXMDwvIHRzHQU7RjEgiDMiP2aXy3YLQoVC/K6hATMrlQI72fkt3dDaeYZ403nZsyPALubdr
/DKF7djBIaTIgn0PYSfsMGlr2OIzf7p6O8xMB4/N0ExrewM+tq/y8DD+80Grzl9Avqjnu/3VGsEL
Gpk+UMGcurUazHRW937f8e5crva2wAt0qtQcnmT+bRBeXWJdzuWC5ZDRm9y6UKOvplySixJS/UCH
vi2LwakrHSQBU8HHNYkk20G44B++Svfr2TxBoFAMBY2k8v/4GOWJMtw2k4aS2UibR/DqvHVF9oIz
rXTycmzcHF0d5Ogbrs5gbMC+Cw2IBEedQ4YbvuiFlGqnh/mPEtDpgeea9MznNS9g+4M/KZeRh1bJ
uTBN9qUQx1ziM9uYftnxZA33JZlBVShu1IgbuMz82JLCPFet3hUQFHagFYyOrm5kPiROZ51lYUal
PXtA4SquZdi/2hFHx8GofM2UFSjCKIKJqbJ6+TQGGxoTWanlvb5gvdKkrmvqDdWLs1q6SCFIB+h/
IDOpl78zB9+iTv/hk4BbsAfZioHig6SyNNpoYe/01fw9gXPzRlJGd2NHkze/PQgTGhhQCSBFERtw
29EsUN6G+tSQjFlahJaCyukfrRClT/Lc5deKXqaco0v146ka7qjwlcMKpw01yTp+Y+BHVofWW1q6
o+2O/hGD14QggKj4EBr5w1zyWBma1Vhp7mCN0eUcRehVgmU+1hdSjse3YT7iAe4ph138dHGL5tFf
KlYTR36auQwVbXPIHqfIBBdLQBC9NuhqTVVlEQI+McGxrutHRdxcFrIA9oL5QAgwnYRjpu6JnzkY
FxiRnyyDGtaxc/N6Fak1HTGKw1iCm8MnNs827S/0b/JlvpcnG1pd4q/8K9zfK4U86SbltM6dnkRe
iDq7sT0+S1apxbp1ckGMslZ8m6MzxvP/FxHEpyGa+Y8AbmX7C2QDFx/DdMcGZPkffe5Yf50C9QZo
Kby8JzvgIdP/vP7gxTlZAhHpqM/2M/ieE1pEoSE8iT2TNah2vXj91GFSMx62CkEmCbh+WNGWqDCQ
MUIuWtWjtSoeAw1paI1lj0SDHczdF9bR6fezVDzvtqIrtmm8Up0qZyzIkFrsvBLtPNSd43W+wyTd
GmWOQCofSXwO/iasmU5zOfAkVA6lepowT4xbHLK/efWkh0skGjdr+/5RqGTl1HP7e5U6S0iIBZrM
45Rf80478SOzkTMZ9ZbrBDhieKYJNq+I/BCLLm7wcec+FTlhsQl2j/M3es1dsZz9zCFgVFu/VZ3Q
KPSqzPgcHiBllhPQcx+OijLblbMNaQ0uWqE83Sl6jqtvLN1w2JqpNIW0vhM94v2D5lyZucj4XtpX
CNbeT4mM1SgXa02FQYyTGxeY0Lnpf7XN62miSz5JgdtwHbKBKEQNFWuldmN2rzSzxuYpitC26XLe
QPn1oR98EReMXutN2VuEEc/JCqOZIdd1DvgjPL1CuTq6gB+hFKMs1cwdsHhUH44btdAvZLiK7N30
FPPf+OGBGTM77XyJxD2FR0Yc4+aa9V4gYcqI/MBmQAMfcLFxsdgUjC5FJeG/9KRrUAQ2qY4Z/ffy
LwVM4zfwkfZUwwwTLtWEmGL4NIzcKF7mshOvg1mPrYBBXEqPOOZ2q4XHX3yW0l9sy7AW/q6PcVp4
EAnmPcMVr+HbE/yNp7XG+sOyi2yFid3djTXU4D6gSSFV6LLkYn4WaWWRJCeetz/CjDgBBgIKeY3t
O5ZTezMT4yppK/N3DonSIubwiUoFL2XsYPMisi47TVm5vI2RXETydk3ReWTuSpjGC2e5kpEIT+GL
BUO8Bz93XBTmXu+Nb5kn8DVzL77E8hb4H/FanqD4MsQ46n6ZHEgWg+tY85Uw+jXDykg+/8lger8I
reZP+dvJfyPxoTLWFN1bP2E7oqZ2q91ljB3vnmd6bAMKIvSruE1to1oYkdpDsKE6QCKh0KN98a5W
hzaGbGhTssVqJ1zv4Vbm08moyqbjNrHLavW3X/ARVKSqTVQcYfqEO0zD0A9UqW8rudPzE5/l9C3q
Udq70aRhScRUdm22kcqGIl3MhcVKGVvUMFYFjL+okQx5sPfGtI5d4h/eE3+P4QaKozbETrIDSRbA
IOr/Ur28cQDK7K97lh339AwdaOjXu0QCFU8BcpK4+7vBq5qVNZ3OJ4dhcxPFI9SljFPBk3Qxap4v
/wlal9xVOiW2bA8AWJ7IaspaHC1P25AYko5nNsKI5pzT6wcqaefrogK+vn2AcOql+lP0ddTQ2iBl
uxTg8ZIvdJA/hnrdirk2FvnVa7nzfcSNWv78XPbxq9xv14oOsHv6Nx3wwFX0cI8HcsxlxCntW6M/
663LABHyqjuSK0ZS1w2JtOim6VkSdbLMjIChLAx72FTF7jIkix2ERAWc8ASMy38BnfWaFCrfD2Lm
1pilzG7fk5SMIke3pG5doyjc2U+L/GDZSDPU1DgxpMNxi5ODm3sXyG8d1CXO1zRnaCPnx9VtE+O8
8dxzyXoNeUBXZsn0X6uIsR26uSeKlskMGH3yQypA52NbRtW7zPWtLMf5fImDK+08FCf3ybl/sybN
MVtHCkibUarZ9s7dSqOI0/zV2IS35fPy9gKCbYW6UP5iBst/xy3JghDHooGLcDDpnOAW8wTeFUQS
YOXNMnzhx55CCUt6zyNnPFqdcuz6jGU4qkUP4ggNE9MmAy+QuSIXOyzFZj9N2fZOPbkYdxyghk0O
eWstJl4v/k3X3phft6PewnQFXhs6hs5uMnJhgEkuicNeF8+qUlcjrp/5SYKcCl2OaWzRAc7GPpif
7fw2w7jC1JPMIimNxMcAvMS989P3s+JU6eKThN8N/c+Q2uCUZYJLvndWevkSMcC1oM4WqNpC5Wb5
1KCddVmwX5INdDZDFDYG0UHxRT5+8+BivzcM7qBAFNKHwUmqTau31BzBsnYnnwZS/yX7m90DdzYX
XQqvadALkSunyAXwi7LzaAainDcqJDXq+bqgkiX7bMS0UUIpU25nL65KNsvwc1mhqWtf/yBe+4cW
2IdJb4xArONW+JlZ6NYQtUCDQn9RF+yKc/LH+skoDjb8ZzsE3SI5cwj0VOEWWXM1qrEVeh6TK1iC
NKCWrSu1WGpm1vnRJd+0opBOR6UqT1XWh/9kNA6/mlcdqxMz0QcbETxbQdUj8tmTL+NVH/hmZ4K/
/xXGrYhThxM+6EmnqNwyWIzt4tdrK1INVRp33KlaxKUbzMYcpYkXkVxzpVXwluor+5+8DSMp4HLo
0Q+NgnLrsAX/vlygSGJ+ytdP4K7P/jsXeW5k5YQ4Klqen4eAoLj4LuoxAPuqu8klYDiw8Zssq+RU
rmQVrI7DQ89fLIp74rn6LcbGWd0AJd6EuQI0G3usFeCwHEZkNhnyTBek63eHBzQXu9kR//9wK/te
Z+XdOzwP7hXfcpEtF3eXJHoK4EvQrPn+DR4GPVMJ2kf7xW0qknH/PyFZFW6uRfBqp/PF4FBSs4ZO
fW8Bt0wPtq81LP01ElGT0KaH8WKYGxGHHNES2iCNjAe1eJOrfss0wG4gzcN5VvN7KGQF2NqzwD60
tdGKtDHZOubHrYNmjQ3sCriLDsxtWPuTaSCuvqFicXKAwrXm0DJrzS6CUDcWo/pE5sYRkq5QisQt
3OgJjOIebHHxQ74pCO9CkL0wK355CkHIuGjjdbNl/7KrV9lEAnWUIomqwx9IMKRrTh9hjF70twgp
etxDuyhK2V9OMvKzDKGfLglEycY6A8Relf1GqyAI0Kgn3QhaUOheaOxLbG5P2rkSky+zE7exlaqB
wSPaabpeTvQiOSezKyiFCI8H2YDRv/SvzvVNOeFFUN2RBhwDk+vSLz15qyoIE+CD+jIAcg+xIdOM
uJSlu/TaRB7qbN9s/3CHf6jSVlIsEYnB0OXju385TIAoWmFrWuaTCzdhYNHNO9xdUw/cQ3QgDHMQ
42C8eU1/694urtRDqOXxXbKszp0r/+QToxKKEp07/ACxtyvE6LJucD9Q8gerhoAfmsrHah8rUYVC
tM6bM5hFnW1/GjTRovIsUA3e6Q2mIhyNQk0jcBXkQ8dImf0uZ7nFqTfcpFiZscTrvAA8ZZ/J2bag
liMGB/O9JC+Sn/kNY+UcnM5ksweQ9RYHatA8PqvvwWTkmCY0gesIPholJmRCBq04trqcG+dKaiPi
0f2A8B1P5Mq2q2H9h66o98VfvQqsSSqgCelJt4r+0nxgLw00EMkt6omMym6mphQbR2LldEftSPxH
fm0Ey6JLCvO/iSUc/hmjshcdaRla3WaChLYvmx/dW50pBxfPzNWc9u5w7fL5GoUDNauYFL9Mtit2
5ZgudjyZDbX41pJDkpug5tkMOHYOt5ggAF0zlvoo9AOPSnPp98SllM/PAQOx709L+7FAI47YvqJM
6rEosmtRU5bJaKHhglEhcXX5BdNoHvTbK7Rv6bHGXm+h3VyPiwbazgGKVTDjIDgF89lj/s+QvAjZ
QVLOIwiK9ndPrNmuHweJ1Tpdv6VlCKfdTOpjUUiVZBQyN6irdsebdLwR9uQPzfcZUopAWzrS31on
EfdP2nFJ2xo5ZqDRwgRM0Nu9eQVzv8oF5WX9cdbK6P4O9iPYN2x71lM+00GXlbsf8TuDfHYDrN4W
UV6ZrQYs9m8pBnh068DNJf2EchggpaKJhMQAb2jCZn0F4DrSppnhrYraxyMWBGH3gT7uBjZrvX2a
WgC3nmAuEvHSidV5su+wDLDHtPQJpzk9Ont2V65lxCre8Cs+ltsjZjVCEmG33PUiGsUaZdRDdshS
8O+N480N36+EUIxmSswVPrF3CVLWjU39u+d3EMJW0WUGce0zVsfJTyZ8PK0hnf8apCsxzX9lY3MH
pbdkwFZ4c2ob2F0knIJ2z3c/+wVvFEnOfdM+la4CfDs1LmoZn5ZDUudC7oQUgRSUtK1RcVFqJxis
jZqfc86AJpy01NQnEFE6xLJmpfuMU1+sHX1jNVaQ1spVxRRXLy57E3e0s1CbfGlWybmSVFo2a3bW
jtl5O8YrlrwzmFTgGj6+/0aSAqI/cMicffOrpC3r9AfDErKHQl5vIHPQYa+fpVYPXRu9IClYfNFm
al4Bt9J7jfiGSxb10+8GPWw6XH30ukPFDYJJ0U34vX8Z1DydMJu80yzuoum9pK8z/Rjxq5z8XpoJ
/g6Ec/zSARXwfaFLhzP75EcuySw/XIIvWKsQvHK53j4PFNAZdr9MjtuPMcnVGWlLvX71q5qXliAz
ibVaVdFUcrcoqQ+RQN+clgfV5MT0HfRRB6zBgA+lTmSUsdSMWSNZDazzpUSY8njrLkBRlaFR9W3T
37qt+cyuBv9jtST1oLXdwJaA/QNdIr4nowwvSXd2mCp03R4K39xWU/w8ZSQrsl1imDhbkTLZ/AUj
EcPS2oEeOgi8hW3QV/HXRaNSyJOo20te5GVy8PBFQHLZ+3AFabrXsKdRI+4Rl5lKNqNawTBoYjZ4
Zg9OZdrbg2rSNavkmuJ3qRcsB4ouvq8Vn3cy0nlgHMSSBShOO10WtjI2Jzue8NCx6V6ngCWutrvR
RbPASr/DRuTyKqgxGZ0ZElMeCNEoLjjNc7JrD14aY7PWBMjV2VkU9UZTk8mLc0oeNhYifA8cUl9A
YDStBXsa+UU4z41OqDkuUyhiHRLoOWeeqnL4HDEHO5fjhMp7VGxivQoPq0BgsXypmeff4cXvTdke
QGjdR23FP42RxkurCI2sB9UTFOwzu30vNKbmi6ojLvaeg/LBHzP3tDMkBaWhy0cPzVeArfsW5avP
veYBwbM7fbZ99tu7J+thesOUkUIde/oP9T/zG++KtBtIQxTi4Oi26YRlVeS4yzaHwCai3ycph3+J
k8UmC2Bto5aPrg90RubBU07cKMYcyf3k1Rvl/SOOVoR0mfqkikpivL0p+1yjGfiOHL4ikokWmm1j
CYxhv8jkHhEVxuKzCAIbq8f4+1c2/kWr1FMPd6ylcDFKPFmn8i3eu1YGbIYoPttiEiasCFxaMkGj
29SJ1C67AQbeo+qQRmtWCQBhQi86sQswg5H2WDR1gi8AmT41Sib4lorqKG9BXypMpZhNzC5UFt37
A/3n2ilkzUJ3HKsekqbXhETjuC4W/aBlISlAAthZmr0e7w0wAHZi5AgZclTd1av17rNR7TuLE5NX
snCV4hVft1EZXPo2onIdXrfeTo9DEjWI1jLrRfIAThKzpPidVt0ACgaRdJ54Y6gQiRMh0JtFwnbf
So2YhvVcs3nutzVniUNy+EDrKTqN5GBTryr99SJhQd1r++FifY728+Q+Hoa+QKJhxB8LDKsTFGcH
103UU2v6kkCoVKvoW05Ds44nTlmodKNBWTB+He3QiRVmfVr7grAZgaCeP2H0MX6pxEAsyRgeLyyU
rJPdMa9QO3CmRBuP1Fmcqta/dq4sL8ZIGirSRd+ImeDKZk+4ImNaHL+LxYCKvhm6B0sPrwT4f2lT
1w/tpAjbK1gPGjCZ9spyBHYe3KCZ7Y7PgYp7kfRdchnYtFkiyLOK4LbkIWtbbK9AJqgS6ecHQYFT
non/CPnmgr1uCkFCk+U+7ZcURWDrNgQYi8hXIVjtNcoAnWBztawF16mcNgBel+nzICm6SayHBfDe
8Pc+BmaABJifnH0049ZSiIch2dBFujWevDISfpse1UkJxXw7EyAkag4KfY/KVxmUDR5c/I6CwHk3
xEQN/2BiLD0yoQYbY8Gy8WUDbOb+P0mH0pOfWQAiTST5e1PlJ3ACTvM1lKqOWeHseNNT0RmYzRz4
wHc1THnvUs4+/CWUHBHmnBed+cyzRp2WOoBeWHHs1WnzUOtTAnjt8uJVzkv63Xj+0vnuAu+aGbTV
NIkU0EFPu03ne26cJ7pXNAJidaIOlE0G7iJTfVjmeOLJjTbkMndfRdj468s/V+nmtzyhPE67jK5M
UwS8SFp939sjjlIZRYDwx9LdRBvQBD7WMPA8AVYa+stSRHR+XKUKmfVFnkzWl7sXbLnhnrCTagET
6JGQjwf7YN/iOwzhmx0PQHEX+6Ri0752cPsYbQq/+3ONrA7UxAch+TPmqMp96vFR2qUjvHT6pdO0
TJ7/3ZLT4R597vlU/+LSvGDb9d96f2m7czQUv7RPGnbOxzmByxMdh9UuWU6WNN7kdSCWIFvrfxiS
IPwLLWz6YVRpqyNb4ygzXsWJkuN6ykkcqxo/qYbflmDHgdb1vbXGR4d3IwnoGpAdCkuNaDGEgOJt
VGsdjrAxAaeK17XmQ32FQQVktchLC1rCUT7Zb5YqytsM6MUZ8EOpU6OBdRY/S4deGgPqQSd5Pdy2
VejAudiAdra8tDM7v8PrGru2calbJ65EQMEBvbo3REU6+7HKBKe/WmCKRLEcXB7yoUAiSkH9z5Au
Q0fgoCGgpaWYBx6gEIam6dtd+I7StMuutvedkHmu6dTwadppwNxDc/R+g1hE9QgH2cJ09LoBWucU
/3CXz811rOJ840ikTz4zdziKgJPnGH62fL3Mtde3uwIs2PQ2bEqm/6s1aigB7rnEwaxsvEz+RrXO
hfK+RvrcMt/XHl9ayukt6909I8RzXr84fWMAZEdwLul0frK1aMeya4ZgTnp/TnpWWsFC+5A4MKrq
wZaAI86deq28uwl/Yak1EC4mqhDb6pDJMmxq2PkxICNQ4dJy6Q1UW7JHG1RxvFe4KtHj7h93xTh+
6zmh0egvWh4Ntya+W57SKQp+kVmeDmgnngwZC61L4MI4WaAVEK6uhUvHXC8cTj4Jcb7H126BCyLL
RYnAr5SjppEuSJXdlBTSOZaXbAsb2qSuTocFAcCXBDyQPsUyeDHPQFxyb9yNhHSkMlfNrpAEwtoX
DxbM8582O9XmCkSs+YiTzzMHYtVK11rwglmxUg9rg/6HUcnwEt5f1h0JPArDFXILtFf74Mgv3vyY
AkEjGCJ4tK8rVt6ghDvAeJJh9wGD+FnhI4iwSEGwYAt86gg6x8xmNhmo3WkIhU3Bo/VMXBTHax3a
pTsflQr62TDx2iyflxeeI+g+DJqKcsqWvCfha/1HbOWVkJZc42ctusLtSIvm4xToA5dRlYrPdk/A
1EskMi7dD5fgpnbnKHQwxwddAlOzBhhLrTyqShvDbx2Q6Gy9dSlEhmEDXtrzNJ++TkKZkmiva5XI
Lp0wbrVYK9ZtMb3U0An3cidvBCTH8Q4wZKqR3jSfO6Jk4Cwy7J/2CH9AdcZSUcLy2xprPOa4tv84
bowom8rIRBB1535TZnIbWPHf3Z9OL/6sUlieKloDxrl/IYTOZa0Q5WurBXian9TKW4o2Op01MC6L
qvuSQuaJKRE0cf0Go6f+QA49giTOP9TLManOHeV4aC9HDTE20mC4JyBJtCbIDOtD14kKb40jmVAk
1q8iXeTPsOdjtXtxwnDIWWHtIEXZ0BH8DtIyww5llRWEKToqYCycWBgqkGNxYFLUJieczH1POXt3
q9RaqC9GOSAx9diSm2T1pPCtme3WFs5t25EGK4KhT9itjPCo9hWfrgbjZpd89qq3I4FbPfwu/JHk
Mlj9K5FfhpVqSh54G1i2chftJ88/oBUbTH3yikt5YXYnJdU3HKwydFXya+SF0DVV3bfRuK1jvMQN
7WOsfgZozmhD93a+VscDW6XlDm41ilfa8GvWhw+jgLuF9j2LOdc/4y6xpyMZwDWNJ9JVBv9AaPhT
7XNqse9YaK7ooaxXs6C1Txtuf+cNp0+Evml5sHlP8M+YyCmzlrRkWnlLA2IAtO9pi9BmhQwDI2rp
3gJGs0coqVZCmNLDYHB3PkChU/Z6rsGNGkvNWFyD3AMJtzj6RDG9l3DB82vO1oLs7xYA73W8f4Tl
0vfcueVFx8hkLS3QAzFSgj3JOyMDY6VsoTR/AHhrB67qo5vpmH1dJqXiLzIPpZOLQGhiog+hy/Tp
UPaOvx7kzrAot/z/u0QymYtCjzyTP5S+ggdyDq1eOjDYiOP9B8iBBG5xvUxJGQTaee1T2DwfHOZ1
ESWOxYWvASdQAK/2IRObcuCZ8E+22o6sI7doHBkMvyUYZ3usjcPWmtcfk3m6gNcXQP9HvkzXV0yt
H46Nc5CgkUvEvVrnggBfDDav4ShkcoBDhPKwF3KAe5Pbf3Bv02EwxGBwGPNZkXas91pGfKfBtNyR
P9kW3g9zz6jLdQHp8/5L4xh+B7GbY2dveBp3LvM8z9Jh91ldzvU32D6jTOUlQ9zETkiBxsa6WFzd
JvFfK/VKrrizRhZVDti95+c3PJ7BJdmpd6WAC8c8sdXsUM9IWf1Nnf9wGnI6nrvoh8iXUpaBUcAI
ovh6QrV7TRR9VpnCn8CImiWX2uNlghJ6xjBkBrImtyq2gaJv6AlDRnjoU4gn7LQseoqo+lVY+lQZ
fS7LjIhxGRNwzufZOLhi8Sn82j+i6mZ99PxUXSQwzEDPjsWoMlj3Z4EEg6ul/NIAIrTPy0yK6KAi
5p3PrlLKN677KFzbpmnK5XDJ6BDaD1+LR31CQxuWbj3m1K0sxgbVc/2WOkY/YBZtrZYAhM9Go9fp
M3YftW1Lkv5rKf7GP+peEejxN6H5B6mQfFJiM/yKybedyN0i7zA0JFOtyQETYIBi0HdYtXEcgH90
xg5Y5j6mpwmL9vTx2boFbDIdZo77ItcHVhreRQj7cKcRGYRvcYJAYdY2TWB51MkqIFllA+gkNGCN
CLelT0O9WKaHpsTDQ3dTf1OjpE1O/UP0ZlJNQLEg7aIP/kpj/12ZV1m/LCzvhjxFfwnrwvcs7eNY
ta/varb9rJpIY4+EWpztNj8e76JfK6TfxLXZIgrqY30DYtavKQ4X4yEKoKUTNkGUzi9mlURqe6wc
FdW4e0Jd1AHnO1felLaCgk1mWmxx/ABHCpNDFkqneZGlLr6SOqJBMhn26s0ggZaUp/oIdNS10RGb
mpNS1Xw7qBH9ilvUQQpxEVHEOOnG5bjBV924RXOUB/ZJBjuyCw4bnVXLh/xBxXkuOqf+WtAFBbN0
WyBSTtf+TWJ7L1Ims3W1JCn0kpVdUqP3f15Cb06LN8guci6d443UqnlRV7/t+f4dnRjM3idWKDmQ
ovmB2nNEm22RpNAZpAJtxUTRKiJ/nxXdQOoIX9X2Q0GXP2r+RfMQmshB3RB1KxaMGS82f7CVvV39
ZNqGzTm+QVLFVrfc5clJLcU27P6GRsAWxjzCIYUDpZO9/MSMfdrp7iit+RTFfIqqk6QzYiqldO85
94psNGOYq5SWftPctltkuSTcCND1/7RH0qcoX+zCS/7ZAVdizlRJQ5S3JoHhv84eexGgwYIObomN
PJhffET/rA48MAxYU88rWOmNqn9aJsJtB5iR32OnvqT8JscnJ6yZV0kY70w8Hr7GSLknalp1+3cc
7tTFFib3a5zAEb+adJG3Zt5kQs57qum15mRPJdZnjcnllDVupDJbD3i5/3iSLrGEA67nbDZICcip
K6h8NOJtRvCN9gu6oNbQqwRnKCaVcA0Z61c3dADRHVIfy0esifUKKXxAQhBfYpJMuA7ao5uIODL9
Lb+nZ+o/eeWVPR8zm3SS1iEZHnIpQpC2duYGYz2yqIgpTRCNE3YZEzd+oAWtVEBAYAbksDDamaB1
TAcuD9TB16axHWVw7ygtyA8ySVeJbZBNkG5sqAv40xCkqbjivyNSNd9L8J1BCCYzIFpP8rdc8z80
Wo20jzvTIvKEviNZ91lQ4ZKeav1yxCy+5zGxVnHepvGRnjIJ0V6SEZVHA6Bclkskh9Ub68xdPhWX
JtvuJ3eY0RWGt5ybFamyPwsr3EI/NcjElTWVGc45OlkkVKiwrA50Sk6rvjZDk7te4BPOgh7chOBf
jA3RVdTYe6KvBgyag+eNFXMlqKedarbJYYoTOoJG7BEVjty3QTs4nRU6GaMM+tIqr4w3K9BLTrFC
rIPhmakdattjE9d4J6NjLnGzvNKwabMf7MQz6j2prgrgNmzBVYUCuAy3U9iT1boPPA5th+4Sm/OA
wPzARE5R5LUxjahb7bkkoENtrn+iYWl2Bqao3oDQy12ecMI/1uXPYV++ukKcKQjOx6kpVThB1fm1
s2PMCNAfcdZU6dCE68J8bKD7nRba30+PwHMHLoQp3Yr9+4iKtiDSp2+F2lYrAxW0aHgKYnJsqX3g
IwdMTat0AfiwoEeb2uVAhJf/7qRc6qHLH6Kw44a/qBaZ+SMBNxuQj4XhhdFC7vsX2xFBk/ghrS1m
xYq2ZDBtQ8rAvjYFrTzXQLP8BIb6aP/lmPzhUSZFixHOAHblpCR3dsU5AFC4dP7RIrHzrRPLsnmI
H9/nxQRes05xaA5xnpb7Y/RuL3YdD8T7j3JQBHKNnWz3LiE3/jISESp9lnZw4s4QFGb8+OUGfhGW
hGW7YmXo6Et8hO/6kuEVnm4xgGqYlt2YRgepIMIkXY3wRmSVdtiAUgnmCca6LumwfCg8Ws+8zrKZ
ldzMti3uj83VY7rD0llRrlMph6zxSdwC2bJN3f2o1IUIYokoJkO1IoyksRVQckR9T1kXsYL3fawM
DcNqKIqdbuSOmP6aqvRgiRMY7Ls5r6k3d4w0tuAxqovirGYZAsrMl6/GtTzj3AtaaqXMbjkGGFL+
P2YEYXMAY+6J0A2BmN3UrOKXobcSZl8zgj2N8/dN+TazCxOqIYO5RDuUPIQwke8g2vl8XsoAnyIu
hFlwmfj117XQnJP9UXwCtLHvbaLQKgWwzpCiND2T1gvf09zXj1rYWX+AFJ0JQbqO1Suzw86hBuqX
BqfexNP9/dPjtjx6JIYMu0+jPrBTg10Zr5fe0j60OaNtAb4Pju0M5FmbO9SNCn4w5RWiP+I4+Lkb
zisrpyPYcVP6WyAgVOxTPrh1YTubZbS46WDDb9VaWH7KPvBUPhlwCOCRv6g/2Mx6xbG1nHtbf78t
F0CIeIit12Epztg5/DR00zE2hzE8WIsFBUP4bwYo0uGcWrctVAJN9NnGnqS3Ou2cXYQElCd+SYlX
r9xiWnUpSITm8DdGmRTIusTXBzVB4TGBN2zKJYTqSp5A2YS32AozgB3yOiu/V/oKQmjNkeneOJ7k
TPxpZrPTGV8IW8yhkg5dXiTd2wS5X9348vSLOM/cnMKWl0ElTpCwmwkRtNEJ/bPnGWuz68sZhmaV
+fC4RClX5OPt3SLGy9Gmxab6b5qa4B3yNALKo3x4JQF2D6JX8lzNoQwwkdRrcJx2frKm7GMhZ0iN
5Whli8vy/AU67wezzGVrdxuj1HD9hzuXiP/XGmQivnzMuaDPIaBzplXGhqK8p9enFq9biQCvcKjw
QaEH8jAhBrhXto9TvHadzn1cIOAI6ENzlRJ8lhY9YVQH2Asn4ZyWv12xaCfHIcS/bJmcSC2rJ+Y9
iy3fb16vv59gnYwON9uP16dbhDfZIduKVpIcADD+8qSsSV6mfwJ3UzYxdj5D1Pt2bSQAuP98SLj9
FFIkPkPModEjY2v3oibxl91h+SvUZNsTN+mbyPJaeiMX47/NwyFJiKNVwMpBv7HvlNpKdEXuxC9a
ZRi14fbfPrOQyAYggvIo/udYdYWBCA32DpUNXNEag8L3B1kQbOGLyLiQ+Swsd6AbNx4QdQowI/Of
HlOYf3HRNXmHj+2TJw8dkREnPwSd+x10nEFoWOAVlUEGEjFEYaM4nuMqZeUaX1mo8tuhQ87ZJaSa
MJ+lQaBuNZBena+Jg82mFbi12V4z6aGUspHLYk7oR6ilIqOTejbGiMhg/56E0xs0Syymaei1jbbi
NVGY+A3dGKnd835TKVE7I9Nq7BnmEOWMhpdeD+0ea1QvmferQCQXV7cJmKZyQMBTDZwXD/lL1H0a
IoFrc2kRxdofHAl+GyyRVPOAPF1Dak6IbLxw3OsW7u7sndOy5oANtlu7ZTG7EF3vO20iO6B0ivbO
8+nzhemWXgacWhHJUWUpn4pH/iDETBrLH3w8hQganD9+9d+qW1i3FUiGW70ePEIF9/DSIMDw9jNR
KJSwTg5KsbONISLYtkdO1Wvn4/wIDoZUFo5FI+VxG89u0iCNpyfs6CEkmVDDtiuFg3Uvg1Au8P7b
3UWjwaFFa3HHhDjyNsR6AUnsMtdVxw03nyo9er/LQf9Fe/O9M2SkT512Z8vvUiU4xxGvshc5aTEV
f2YWGSL8B54YRbKc5jjveAaVW9R42sa7v5NTvYf2ywa0iwXQkPEAGc+/Ddg2z4o9++P4aYsQuXnh
u4sXtT1G7T15F8rEIPCmp4sdaQInDBKv/LNPjk2Ml+JL9tc1COUewU2Jk03c0yvvzVnc3r4LOFZR
ROZ/8u0q/uuIaUge7x6Odc8QU4roKds3BJzVHaCrouz6jCh0ZXxrqg0Ow8+TyaYKfYXQeLBiEiVe
Tun4Moe7yPM9Kw2ugNELC6W+zmGERyty9s+9pmgt5ukOnoQSLn7o9th3FywMFcmKHwQSXgwo2yjr
zACpPNsk/qr7/KDieL7YQfWUb/rO2bMsw5KwqLzo3EzTu6O9+lPSHpyjrp+oU2mnZjFY3nzcVWU4
/1gr750Z6QrvdE4YhP0yrAVf3tTswNJalFy+rh3qrPz3Ri2OBwWtnhq8G+XweOKG8tC99nCqA4DB
dOodsTZqs+aEhbs+zJqGFScL2ack7TvUJyGGfx90b5/xeCB2uhispxppcwELeqfNGEldVMauaUP6
Qsphsb9xhwQ1mwzpl/CNyfaxCdRSK79PJhhE+7n2xIrq8N62W2MNPGu5JsPlPLI4i/qEr3IMUKMq
//3tggcp6FqYHu7z6wMnAgC+O4vxBZwP7SQsFfURhVHx0zZt88Bcci6v804xN7eLQV666RrbMslu
wEok3owjxXbN7IKmv8tY7fHqu4YUuvQDkzsgtzw3SLCu36ecpo9RBtFu8hyHhoG67pWYt8ulXlx0
ATYh1ggdQ8Kop1pvesf+3kWHZVMWsZMakroSDejYdyHuFm2B6mWRMdM/Mc7iIEebR2wkrTuql/f5
+7mlBSFzipEoMmCSAXhnNN85shWv6GkKueLpaERko4bjZDAcZ3DTjg8sz/jZFJ0VzblccMOIyby1
nDprmqFe3YBvirpBKeVKOMuE60ABat/m0vdFItvVXfedbFthAsnHA7pCP95olHEz/w/kZLtgRByc
1qL2GlDhLo8iwlfh9o2FZIxdgDvX9/RGzCaLj+55qJKPAUbkytdKquxoz0Bj3hQaaX2GPL84Pjfo
03xY0pAU+GcGOl3vCYIhkWuzsXUNnZgiB/fGaMUHEtULihC7mkFbIFncBRzD7/LGM60u2Jw3h63z
3rIneIofP5EhV/0m7NGZDhmw22BiHhJURdnbTw6EIuuec7JUE8dJyrHHumKnx0nPkxKpvEIDPlZW
P2WY6epj2O21UcqSX9eQtMcePdpEcBXTYD0bukEYNhHGczJReEw38kd4ng4hSZNp+Ts2dEdWc3c7
aweafxcgusi958lIPe0ikrkV+d2M3Flcy/3oiCu9WJl+K61R/RVTT9zmhuWOykZiDJWmdFW+yDHV
ddItfAGim7R1q4FwN9C7g6j8AQhzX1Zku5Es387/ltQPWzPO8AW0yVwJfDf4fKh+dlOZ1NsDR8Ky
4gdsq6/oxK0XCRADDeQjpsjGtP8IW5NZ4Jbbl4lUX0lHwL4CNhJRNaXExRhECd2AuFgpi7wIycnB
sz4HK1D3gFuN1Mc8daICnga8s3To+BW5loaXvSMSVml+2gCZoxXq0bO9arykIhine5/uQGaEXhvW
LzknqKi8WOvTwrloGvVj96vbEz3vbFxmUNsAunv/Us6Dp4Dn1RCbOSBldNC1jOEaAOZRHV01ZGUB
Qcm49nCkqSUroUDupscLys+sSl8ICZLyrVu2KokkGXXqkpr5kGeRCMpYmfTx86dGWxalSemtkxny
tFJOWQC7l/qghzeVF+LkvfvaoGZ4sGjfQZGPRCki8DpmdTxLHMfGGaEqbvXRFbqrN4cgrA9gAryC
L5LlvGtm1kwalj1SWE3iJS+iFpLsyJb7i5uiPMRiKyXya1egLRrkJaU10QLU2ECwfk8D/yfXHVbP
E974+NGvGwWpB3SQh65/3Ca+gu1+Y8DL+soJhQHjf3kw/nY3CS3GlL42fY0VlsyMjcTivtaDcQMQ
YCc2EDBc31mpToCF1Th31OpPin+DrBqC6YlSvc8psoeaLKj2b2koIKKeXq+C16/58oLu7jECY4FG
tru4CRYg9Mbf0gHgH6f++9cHy3BjhtrJafQ6p5in1M0jUyK643XJ4+RhoQCf6aTOwV23RzE8E6Ds
KgYQrv6LlsqewkZC+svzCj3HkqaSp0eU91K/v3pB5azMb9gxOx6buE/0l91IH/WAVlgIJDDfYDg3
JyTRCU5IYTptBqpVKzszEYEGuhlD6dmLnT9HKNa2GCvMgQ/WWT3AXLZWiDL7M8FhLDSRuWenJhrg
1pZukIyrc4Rg1upiyeRiVyDj6Qch42/8PyOpe3GDxZeHGcRHHdC2mZ6y3dNyz3QhtDxnSMfCMMzx
r+8yoYBPPQCXekkfq1f0rjMZYuPGlKIZhqzBAG8jTz7VWt7cgJPmtWOzzdl0zYQWmBEnOmK5r+MV
cB4eLfkYNjWINMkaZ8Mv/wetX8WHtTSyUQT5n2UHIRbTspjCcyiVwao1unm4UgBzbfBWvOO/DSdP
ppD7UARtCe3Vf5BU2/p3FccTTHG+DCst5QSulkIfOR1cCE91VnM07jWl7aqlF6/jw4nMRtQ2Ogjv
oqnRDkjyWmeSRBzuvFDlmamVKVeH545TjEg0nLOtJBH74kahJh41yh6l8d/5pOdLq5Z0HUFQHBwY
nvjqLLU1k4jbbDdmzrl3nkPsV1XmV331ayTEB4f2QEQyShuX3aeEwUpo3a60eQhhl0VtFYo6ZuOG
5Acs99fHHJ/VTLqGOM0S4S721SiUXoxU+/LUAS+dfi7Ui0xVGc9Rl8wRJhGje6CGY7AaqaQ1Nwli
gbPmwe6nJAekMUFw1NmZKJdlDDwJaPQhP6dr7OkKFlQWuDhfCOaFZGqwHTzyYJggo/apIN6IZOnX
2t2qeg6p98PQtx/5Mpu55jKKVBsL3X4q/HSy9Y52xkpMN/uxhOLSu2aP9uS+yiCnFxNbQeYiWtx1
CzHpsVd+QzsmwoJ19p+J5Ein2hcgVAbO4cLs4SxUWIHINxlgdLVqGaAkB4g3Y7PfbBtlnOdTE7a/
+7hd3kZHnbVX929SribvSDoD2MNnzF+NFc0UgxAsaz30VRubzDEdb1Ps0PSE2W0ESMDStP6DGrIX
0fhciubOR4666IBwMxlzQPEYm/RdkjOatEX1l49a7ST384xP415xGJpkGakz36/Gzy3KnPMn0X9C
mrq3d3spue5U/zHX6Dyrsm1+M47+yf8C2qzplcWzHBdiNar/1uWZV3lSVxMuYH/siwI0TuakinEb
zB0hw6DUFJ5IoOMaJaNZlM8Pj/nke2gEN2xlp5+RPFAenXJDsLFZ0goQBDq5F4gAKgrIfHOHKHDK
xt/iAD4kBzgyQpMmYUkfsYLI0sN8a1Jdo4jErE11Hns6dpQFH0Rs1fZ0gt6jiY+igcs0apKmleva
KjR9gAA1bGDLMBtQi4BifANUOfykiZHaZ9f4/Ua1nEz7FYD8H2cmoa+vB/i3q5DvG25znBT/a/ub
hmpR+77oE8ajnDQGYTPr3Zju7WBwDpOcFaUk3dXrdlAKeMGUk/HFvZl+FP+Hyq4kr3cU9X7owG1F
wkhX3hhlFDer/+DT+fX4/Q20YSp3FM6NDE0S8oYBTcXFuWuT1R4CSo2U7Oev+bwKXw4fYSj5cJ3B
rLzx/aGsroJOYh1FZH4SalONOp8g7Yiki7WxQ6SaVBdjKpa/fxWuQnlCgArw+7l1V8vJzM2SQZ8G
jnqOUXRoWBJCDw1xBtsrqjbXW612NeR9aGh9ESKJJRdlGT2S9zcDPaXyb1g7cXzXv3cfIEv8Ua39
hswJHxae2KRKkLDLZ/bwZt9/mQ0xDbjWCOJlzMxFBpoJRB+VcrMQydp3pdDFEVShI2x50v8E2tTw
2O/pXzoNLTnnMvZz91Jkb1svELLp2OZT9+8TFVLLqDpT2zHVeP2E7rDlWy1znvQv0cS+7geLAx4X
V2xkui+9JvDhK95hffqhiAbSF1ltqM6f7puaDaAPJCAaG4ZvTE+/36z2Dw9G24SzEXUhumnLmteP
NGZskCfywLRZd5W8r+b0l7d5g2VAzwuhiXYquwgarudXjlrrb1XY3ARqfdOqiNFvdJ6Y43frN5/f
1ZUAU5I5tmGaLcXTQIz0FXS2LA8xlxZfIUXiiDst8GMM/iUbTqbsV7d5WaLsMzFIvZQxXsb52s6j
2t6mqTXqcYjrl+FLWHRPsE4kvZdCAm3yaDLt+dgCavGJrNFxsu+/yJ0Ht1u3JEdAbo6cKEGkG5Ez
lvDgUJwh94MY8chpOSVsdVGHj1+ZLZgzvxb++lQ4R0OmPhb3WlP7U6cpZOGMmderjho1ZVoc0DMh
yVISFiqni2fFbvcJHBROG+ZN7WDGz8Y6LUt/oM3xMZ9DdG5wwdnx/VtUS2/T1uX5IBKfpw18xsSO
CvdHPC5imjbXRIhWWqwtpf8ikySquIRyLwoKWi+mN70nxIWzyf40DCDoVKkndF9J7sEAaaCRelE/
s0JQ3NV3mEe4YyjyKULmbBDG7W09z49omvFse7iZhur51Av9ZxBHFySl25/WIrfoHJ0WTlRGY5bR
UPJOYCe57QIV0tsYz3Alt1a+vCmpMoUkzgulJ04OuzlpumWCpdcxobuN18h53r+GRdqNzc55Rhz1
s0yF1fSUxSSiEXf9cRyxjJ0v+atZzp4/fbnsNiv1l/U/2LA3lV4AWQOJZvW0+pldrAcF8k8Sc1l5
ySRkNUE9eye5VA5FsHciV2Lc2v6eP1raSVgCf2LIduEFYIp1A8Sc295KDBC2AyVP8cIyXTqXqXgB
RqARzvlWsmI977uUJFe0ZxsRfCZIvdcpCCP3YxTbID070OskMVrYi6jgI+gLmgK6NnB8IfgugCrq
MZb/NWvEnbZl/W1E0dikH93TghO47xr3LQ8Sdgt0CflzB+sM7w4cp8Lna1/rGvpOnilNnd03FaEv
VnLVbvr9u+MKG64eTzA9gFX+HaOgKz7PHwIXAwTDoipWu///uJ5+KatQB02EtLXFSqLa2fx4Th4C
6SOnwgnLsjgirzRCxmwWTEHbOMlRcaFTm2sn0mrpGmMsOHdF68pSwgHuFF3EeyIJ4UI3HCRIqHz5
EMWkU/DopnM500flxVUvqoQHAm4tlqNMepn529K02SsGTcnI06HxLiOoXxn8dcFZ/cuQ2DUd1iFh
V+7pqYRr81ItzNmzqhM0ho41N/D6dDlU+7WS+Ho2WIDPW1QCvaM5P75TqoGgQBulL56mBD8x1ULY
A8z6RmlZOguaHGkKQv7GlDCLjZ0ibejyIf/pjKkLxP1NSDY1cjBWtssKIBx9t3xBVG+2ryadXTg/
nPMR6I7K8i9D+rgEWFi0wcG9TWSsn++74w+son4f3LYsY7iv0UiWPBendnRK3pWEqWKMgthGD7RS
IBemgVbsTZ0OrmNpb0tEaBoLs2My7+WSmeafyIzQjqEtpqaMJUpRM9RT5QgrFZUhA+IENo3RoioS
khXYWUeLgVXz2DzpZcMK3UEv0aHQIkbrS8PI3oSm5pVPUDjglbTbU4gvkkl50Y2dX01rgZyNXLNP
RGB1lW+cR/e8b1YhH8IWVpPyH0I9g4hDIk/POABaLOptbSPzjFLeP/uz9vXFd9UkKWcTvSY+FaUi
rueyptFdBfsv+NHXTRo4JrQuKnA2FYZjiyhJXSWlvguU8yIT4XC7HKpFjJ1QOU348Ey9to/1AVHx
+yswY5K/whqPhe0fQNtwgUffRshNk81v7fyDuIwf0YX1Ia8i1u2txWrjAnRIpMwNLP2D+Afv1oB3
5JK+yZRPoQJTwFlvUFo/7/yt2NG7QqSKEByGfEKT0t/l2aKlbkat9AgdqHf92xuc8SCa+7ES//mx
faOM7+5DjG8cd8ToUjStEWYK0M8aFW8ytt4IuuJj/KTUV+ik/TTG0VGKbck6ACkdJOgI5UqUjXFg
m5UNxWGT65wbiCfV2iRjejX8Y8nUX4D8jL2/tl9ciPAKAwqnu/0yenEn24XPSKOZlwekPLvEX2NH
924mIRJCR4eIloIruZcP8HlFtTkXbd3sTMoDpDaFqSqjGtUzq0mjMKQsR/TexbuOQRNgBVnqtKZa
3JqbQG7/U2FVmOTe5JayRLfb4Zv75BNn6nyPvk5m+SaTaOYqReOecuWrESWR+Md7QuwIjbT2BZTX
MfyyWCucIbnPKBNvGqomCNpgzUjwsGnWHZQgdEJxFzPhrv8xgEW7Yo2rLRz/v0b4ouoBCoO2iHgL
JQAwY4dkJRf/HJzr4qXrKJ+f8Ckwo7l4Z2q+U+9ZxznzZJIystJGUrwgyckwoBGfoQCE8ILNVboI
P8m+SkRK4PpCaWbzqRcQr94tO8yU4JWuGlVMLXqpbkKYk3u14v1HnOzP7KOUpIKuHrFnmUaPXI9x
EzJTkPhLK9VuQku3IGs9OJng1HhveB244jK5JZD4SLJ2FaCjB227s4ci9EbslI6kwC11Bt9IaOju
bsb/j7de6LEGQ2dD31scL+HkY4jX2gGa4LauN9a69ae/WrUI1ggkqW9i/ya2bsUZOeyNagfm/WWh
c9/ON/2kMkP31NljvoSZ8j0JVDsV4yBUiuCe90YepRZJttuRGBg9XH0DiAxphZ6/fyuG/Tv41V2W
8BQuFJcsFq2v0Ga1IiqByR7/kW71X7GurQOgVt6M8X0lKMWi6s7bIskrdezLq4HF8iPosljbzuIb
yO8rGJeQ21jxuJjpUkhCnbt5sdarFnE0zcO+7NL18BcZvRKmw7Py0Q1/q5zwme+GIwp10WmshKz2
N9FzQ1cTb2Xc5fYZ5V5PAyc0rbKi4SJVu40g6K+zyHCZHVmW2wOfK/JnJW7Ozb1lWU/jTHAof7gY
8cCknjQR+q+3K+khDpx3V2h8mQ/eJI0+CSlR/gikQgkEAIg+rpjhY8d8qI1WWjwCp9e5a3yeCuRk
2vmHQpBDpOjA17UsflRUmBmCbUVU9+4BMHflkEBKoZZfwIsFlT0pjw4dhi3hRk1SJ/y8kbZtKloT
m35q+V7GkjtCHUff+FEUJ6SMBTB6+GANuUDNZOo8ZMIoFJapEKi8cnUOSPNtdc87rapNnMHMnprf
kZmp05G03957Q3SKPUqNK17NxdhaG+42naEFoxOVGikmZI2YZdo5hUxRMMODP7jE74RQGbpwMyjC
qM7ghUB4SDmtpwuhPN01xCZXHpHvUyRj0hAtybv/eQm2oMamZ2IrH1HF2abl6QJ0R/CPwx82GrHr
yV+z1EJ+LCNUGJGP4joVoTPUl2QJmgXf4dVdMcS7hHMMIhL1t7Xgd5KJO6JYFvQ1t3n6zGneMki5
KOpvTiOWdNaEXM4o+7vN3592maSpQkiBtMygH9U1ytZK5sC6/yH48m5xbkJf4bDhj/tbxPZpKo3k
l0icVuP6/WtJ17oUtRKSCJEtGOIHGKpkN+aH+me/N0BUrFGAg/SE+vPLHXgFD4wfwFqXUZbqMcf1
gpdl+feAxjjS9Xu46dFOMyXcwtpp7qbQ6uHzSBvPwMscRi3Yna3aI+gqIwGPo1AdUY3dcSm0Pjha
Fmyqxn3AqKyU8iOexScbd7GQKPVFsz6GOriIdftmMlAP7ElkyxJy/ey/tAlEyW7qC5MvWj+sTBeH
hDQ4chZb+vkGFA+NMjsVL5WYmfwXUv2crf3sioiN+nzSlLsz1oMQU0sVAO5R+IB2ZQQMP6/In8le
GJaUcdDLXpkXvm111qbVonk40kA373Xcrw1KNjGnYHPK5dveDJpz/CYgPreOVA4ato2csnQ8u8NH
c995UmEsD7FxawAs8FCVcS21wvetzMlTuUSsqeVTC8VbmfFd7PQe1DDg/uBWJ5SsJxC0JYOIW6ql
QeQJV3TLVWbELBbbYSnNv13/ckERzHzf+My/taOvlmIczrkzuHnl1Tk4I3eWpDkWfDN+MlvQN1AH
bO2BlHhPi694EJV66KxkwVdhauDe+OD8upCJnjd2VEjuaENIAhs2rNM44aL0S5wDCXvnJcwySqDm
E9bjjAdg4ZpyspW21Aw+2Diwr5oFUfmKW2rNgbojrwRSzuqhK5E5thj+3RR4MNVe1MgkXm29Gbn9
Xg0ErgK0EMev7U07iig0fgf4iQlbRgGub2vdJRFtLOgKF6IfYKqTPqim0DTeIikcw63zoh0DwtPp
u4azaVM1kknTR57XA+fUFne8hwNnoUC/S9O0fL8X3GczsQJXY71A9fzmL6f92E7Np4ov5JlWln6I
qj2zpo9/rWAlMFGrFT/Odw7ZIWZI9cxljeIv+CaHYsFw5E9alh3cJlpKKcxD4wpEU1GWZ1ESNhKS
50gTvutLA/Xf0GUfuj/Z+qyPKapi8ixUTcRuutIMuESJorPbmb65n6cu9vbml/9A6/u+VqrUIrU6
PA/kuNDUoP8H5+21dVt4zhd5cG9yKIZBaQAfWEARLp9mZ14ZWkK3anHjYs743JDNtamlyHEa+8t6
taatOMXIXI2DU9YgLHDB2VceNA4DbDR3v93f8ZZdxi6V8boE+VswAI8y04cbcNUdLpaDxDQk2kub
k3WQK8+q7HxlBI4WUwK+lbOuPvnz7z2KIV3U45APLaWqpcNgyqXE6VE3wvbYzsdchtHZbutJ6OnM
DJaQ/BuGIZ1OJY4lUXyLEHcEA1xR0V78FTr5FJvblg75dCiKNYue/860ybq8kRN0TQgb8qTOn3vg
86Fm8m3y4QWxIzgQbqzeDilUjVIm3yPBk4H3FUpIvjiGk3QO+SH1kI9lImqdO3nIKVnVezKUhPrA
D4SORX8HkDD8/RMCGl9r7YSVlJdt5OH0utVFBGJNoCHUsHngxCUMlqpNmhRjbmSzV9emUk9a89Q5
cSabv0GmrJiq/5YM7GoP1j5AG9UW1oHnAKTHGnx9yTzoRIbUbGvDSPPDbRWc9hZr5ILGiyumF2ho
E4crYYEG6ZBC0keNDBo2xkT32nhZTwAWkXzePVyelZNYgZkT0jOhQg+k7j+thq113VDG4qdCdzxK
M8b/0EG/zz2D88hEAWs5a/xedeo8dXZmQYroeIw0iOi2d4/lWZgla8Z8LfvRoNz7Wd5WiPsCUaL6
aGb+Z5ZizTGkVho/ACAMtaqv/nsBQR2akOWFzGoO1USJPjcX0mFGlj5vgIHBvJyHMenD/GAoKhc2
9rpPeayFCVg9qAW6nnK+2DVFfPnHkyMC14yOzGwJ8o0s7YRzXeVlu9Vx2I/+4MAZt9pQwLSSmgTq
2HB/UEZ+P75ysu5yg+941fY9XkFQNU+pm3RDQqpo9VC/ALafV/TJWW5G+vpTTvup9a+axu5SH6IU
WnDvPJUOvIVcFmYnGKGiJHOHehSsFRmPRTleWZ5fXS8A1suLeIE/jcV/eNoRzZAXRLRhDSJEVGQq
FQdgn+1H9WeuRmWTZ9GgltNtCwl6UHV6D8KC/v2wd5ReiklcLfiwZFIZEIGM5IFUh/R0k5zRJz8j
BeehYdtFRcTp8nPPjGvGIbtKATR/F8D4CE3H4LlndkG2MacpxeL+/+VU2DiCYE/Hk7lKO1MokIsM
kJ9PMsUVzThYm1g+SE0/q17zHXVD/PX/6NK7xN/enBvoJqtg1B6umUuau1PAVjm7JqwN32OeMljh
IthuW0ZB97+886pQIHawLz0turOxaanzSimmT1VCN0iS6LsKZIVhQUWzhvLacDpvusE7sw8r/OaL
lruWyHRvk5caUPOh8RiHrNq7LjvVXZQZTKpdp9w7kFu6VEB67tcpmbXVZeBPCCCkX3EiyqHSZ8aW
rROPBkoYtMBjh8MCRO2W+YdGhde+oyL3A9Ntwk0n6GZ4tuJwdU9sCfzx2w0ImqqMgiQs8t4MJZwX
LFlYvSVNFRQHUCyNIlwl5QdR7x5oAJHcqhH/rKRApYBxPHCZvW9O+VPPluFJtrwe6MwrAgU+Q1q/
yc2RoKjfJpxFXwBPMDgMRRQUnH0sgi3URUq3CLjKwMh81fdVzyXtBYKzfujNVdQfbkhfsTaZQRs6
S9ydVWhVfWgwONngdfY6OXS9lyyNbV5iCPDOT0UlaCCFIYKgD71ivKlZ9C/ZkNRMgy6k0EDBzvTs
mKUwzIWIa5N0uzDak9bMMggjrtPyJyFx3OYphT9dlWrndusnBZovtznIWI7xJyD1MY5wwQzZPUTQ
+XEoraX6JFsfGDvho2CKnQipaptuwOr96eaAgafmqYTok1T3d98UQJwr1lc4UYZ2E3W99vulYiyI
cCaykFLZZNv3wSuRZhFwHoe7GDnCO+eAeMfYhG9Z+P5jqw3BtpfZ5YF77kye+1JxkvPP+gGbPIQ2
mZy76jKQQouqb5lPVMD1imHATZwb/125xQ51mHGd/SmzhOEK+0aysV7j91GSNLEROZR/jWYkz/dd
WvWGIsWwGYVzHZWNo4TwhKK8gJiu7k9MIa9hi2NwsCkr477GYkoPidnpcLR3uG+yE7sgb8+oMofg
9Zly5134ba6rNnldwTv4Z+qKvDtgq0kFiKwkDJpLL5eE2nB6mWsTKBi8EM0ISkdDmruDdvw/pTCc
X/vVRkr08B0+MRZiGXcdtEXFGxwmnBSSWlyZtzNwiwx/IO6LR0ceDJ6+yeubiTfoh0cAo6OfcUMu
9PKoSesmi22fjY4BydkxlHwq6ESSyQR+XR1Q+nw8GK6akN0kPDrrngmdNLFkAZ1TLAvSDRWKl9fC
Ar3kL9HzFWP72OuJjzW0vO0xxbBWoMWysm5CeqyLtt5DEGR5vEhTXcJulBzHevyHTa7aZmeHX26J
29OCZgLaQaNtDkYGPgoCb0MfG9GWDUoGujnADBwXeUJWL9XCrlDZpt7QeUkpsrD43AN7IJz8l+if
1vwBT3VTh1MIxf8cBdTCkjS51yF41b5RWhy+gmZJ5HSv2U3ZCKEl7D1OqlI1d3XC0pKDxUmDwYPe
EXH5IoznI46c+yDRBAmF0jghBzI8dUnhnUZGWLRQ6LsOBXI3RIlTXFA3LFaLxVb/PLnHnddJr6h7
rgSYQd049TOEo6hfn+PX8Z98cfwSvKdwAfCYfQEVOykWjvlFjdM9HGv9VxNrTYqDECHEwytTosJv
L7X3G++mE72GdrFSlOk0/jMBjR2zAz2eePg3//dfOKX8X6Nw1qTtwYQEZSZgbtX6jgpxx95tWpQN
R+XcZpo9a8QcAYQaMqkBkdCagDpVsCkec0yT4jyah395Ehf60FJgOANTQOnjK98i5zWvCFudu9Tp
2NzaF5ETfo0E3wZwQzxqDYSYeU/rxJIRHYpXXvPlVj34S6txAFanJQs3Pd8ofJ8A7zfHeBI9UsEO
ZxYOOH8C8P5cE7ElQKJzQ4fMfCO+PGosYC4iK1BEzBgLGum06YEpq8/YMt1MV6qRBV4IZpQ2P3/V
NlinwN6G5pG+6JY6loG79xTTYbatMonf1ih/4ZVbw7AIzuWYG8RTA+fRZfYy15atu0xCr+lvjnmk
BkfXMqBL0FgjF+6idzVO4DpMoXTbjcqpUq1EijKK+XM8A8fcUc4KewTLBd4FBgjZudxKeiTtLqGQ
tR7Y2kKOyPr9B0DTXl5KG3VmS7Dng2VK69vgFx8SJrJnyMlnVGDRQXPRWmuFlB1GEZxgPbiCjmX0
Q1EP1QoCQc1tuvQ1Y3W0DHUlFheYTN1H/LINkwg99H2yB92zfl5uMxA0E5YRUwjOEtkLYfYYpr/V
uN57CUfk7kARkxhO+NSd8U9gADNjsnof39a1T5Qw0by4YQB3aduw/WbufEqSEfqfb+YDJaVXEnrE
5jB4+C2P0QmG17xw0pG7UXfWPRdraEX6t8qfCYElo2/LTOjFv5+WKzJOWBdCTI/bq/Mk+xyhj+qf
Q08Kzwd02UI6BkGhO3NoivZqlf3uAmncg4WeNVM55leGLOg8Gpsmli0FEaw+r0pOU3aOmYicc9e3
PRsS8cWzUSd3QLWOfnfk3F46E898EFHUpooG/xpNUwPEaIzbuvMRIFe+OaVorS04MTJBgqRk4RSS
LPlIiWMMVpJz+AgN1Ba11BzPxdP5GWRSKGeIzOmjPYfaaDWHvv04PIfnkHmaoJWNd/8Kv2kgnsnr
2fJLIy0dxSNPjqvfv92BSnfIdXBxRSwNQd42jApm+jCc6l5bnAa8kdWxoAOuFDZFvDzXaM1H41km
zGxpGWz9Os9X0gN/0rSK3VGHPjRpQc93ExLXNqZIzc5l7Kun+R3sem+wa2uyq3Sg6EWivgD3zvE+
zr1Q4s9SWThHmAHOQLMrwJbq5JWiYW0nhWgO+RlHXHP/sBFiH1RDUrozu1xAbdvy8jDfLwGgREsY
S0enJ3wugPSzRdPL53WBITexCkNQD29KbwmJuuZ1q4Yid6EdBKVcKfUMMFxGz9dOj3nK1W8ZHbKH
6GlzwiUJ3uB9HdPn0U2QmC4IflP0LktjoEVwXi9iOyHSBqLx3jtE+ACosNvW/gp7wN+lvn9clJ9K
HK3hsO5gbIZMhiDiUWab1qJ21029XFuCgTMqMXAHWWoU7N6/p84Ng/qt6KMPxLD09BNFxDm7ehPK
CcmZbVZ9R1G4eEsmhiik0+/BK0mibl8W/dIvHTn7zX6/Xa8BAoZWhR1zmYy4kIOqD6IoAlu3TChH
jjMDIydoP3XMj8CIBLR7MyX93IAPSeH0De6A9Tzc6pI1h3u9c8A1fDB4Fw1Rs7c3XZyaPdBQvJbh
a1kVaOiDSPlmzZJRjvUU68rEHgmA9riXPLTqBh5rRRQIrmAHfbKf1iTePs+XuLX5rkZQsvbeOMjB
BK5Gbf7hugDKw2tgSlZBzoWjWjLNpVrcJzFVpbqktV7nNHwVbBOWLkXAUXErZM+/AQbHpf3hcVPy
Bs0+579wYG0Tiy5Z4kKnRNL4gylWYYLh465x6We3V1gVsaFSKyP7deKFEF/TVfZse4kRqwZe7VSx
W66I2DMVn4cBA/2hZPbLsShuDVi9RbmVbnjzo8u+MVYApXVTKGDqEXIUaGN41G1LRGNO/EZRMxt5
+jG3WETHavLEMzCZlFsf9ZcEMZDlgjdVG6mclcj0ZbLNlbwcfWPAAvsZIDm5VBjZ/Bz+stx4Cdca
o+N4BuC1tZHVr/72htVbBYFvfdrRDUNLsI64IjWaNyXoUr4XK089gmWeOIhmvbNH9ai9+Dqz4XH/
r+8P/hJ4BI7TyiME/Y9+/1tNM4NfdPZUWnUpsv9Cp1njglU1cr8MmgBNz31TGUjMWURraW2d8Kso
cUjmSLR+DomDV33/0vz+xmTIJ/lawTl6ABKH7YDn/jMGGWCHDkZpoSYwxSSxYdVGrNq1pM7FO+Oi
2X2WkSbWXt63O7xKu0eiG4rQHTswPMj1A2vNcoHBrRTN4u3ELwLTo0X9rFi3X8ojl+cBFlFXcUJw
uvJBWLUYVEquB5izXHb6ctLkzIwrzAmoY6KUL1cWz1R5nD7EkhF2XHssMVljkyK+PFEcUTvxMZjs
fnn22xDP1P7wBHFVEDhMP6paUi+1YqzR1Nw2wNYMZa6qWq4sWFLrjyOVkZhPpWJKMeDVWrrPO0Nt
auvyYkV90DM0tWPzuMrQkZBJ0i5Cg/LIX+4FA6aPEDNRAN2yKq8+wLqLfq8Btwc9tEhFgR6KS7PW
Dg/p+r6dbXtMRoL1JRdbl0QmiQ08yJKAN4fuouznm5zEONH/6UoDETcXlzmvl4vKe2c0n0N9Y+Z1
NrOo3ivyCyq7OxJMMyUxa4fh0A7iHvSlrYFdME9lAKHV3k4pWtgSZ6dHKShRma3z2Aj9KZy46Sx0
fWcKONjJ95tGtxw1BgU7BTJ6/BLadjMusoCSJ2UgdssN3XrVND7M+siIUrpaMwu+jAWyGFk08oST
yNNzhIMw1ChKboVSdjXzUv/g2lrCbAbLzmN9RiwbaUXmYQe1PJ/FIp1gVIeHKagoiMvYthdTwbsW
9scG1SAgnwiLzpQFE2a3HKcalIPXmtvaaGD5XXUIuKnw9RWUlYkwihblnT2K0MeXgblOloO/BqSE
2AX9QnNkRqMwiOxZJZ5bNYmhZe9O/W2gAPmaG4ShHb/ougARodPtuqVA5j8AbC2l8jMQe5wNDRJr
vwW+HFfI6Mxrb50q98+RSD78vKiLdIkCZNRXmZOXHQPfv82rXo58TgUgNEKTqqSwaoMewCXnOxOe
eI99h94JXbALnlYYgjw6oA4BnlnKZgcyafLAy5sDUz2HxGc=
`protect end_protected

