

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WH/1Hfau3yp/7ANrlzYJ6lp+xOi/gEnoXSHu7RquVCgxmSwM+u6NJ87pS5P1rM1REfM6bC/4VD/K
djLzpKr9YQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K9OQ7UQRJNNsqlJeKiLZja2cTpdn/7D08GuVLJ2Q7YwPyOa9sKS+3g/15LJ/yRa/zU+A98tod3ce
QlWEn4ue+HTvQflEH+MpavwOpNzd9uaRdRTecGrueadi0jZCWhKDECPBSOBftTcItmWjS+iuOrYA
UzNSV6gBgTESSUMmlbA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rfuGizF/z8gCeFD2+mr9MbjRWuTPDiFayAy9W9SH59KTv32ja3WRqyFVDNKefGFWmFgyXwscsdSc
S/STQk2WVtfaxUn47IIZV3HVYpgEROzZ8tdQyrDPMbi2HwmCfaz6YD5xdrfG9Tlx4ToidJJ8M9l4
XJdd32TWh7NYEzLxqVy6SlnR9JfF+0+Nf5C57mxaFcf8i5qJ+wGXhxEFyHFj5aPx81iijRBXdTZB
X7F/NtLKVCgLQvWL22LQZOJhyZVP7Cypy5OtaouwesfLnz7akydXxvJf1kqXrAdSNY4YWjxfZQKZ
dY2m3KiIO6F542kNq0ktevUOXRqWTgZJhPauRA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IUtntTnFOD14laEXhqBklNwiMVlWXctApP9259AAx8PFHjFAnJ8PvitVWk2w4ALBNs1tWO3QG+lc
7ANJMKcNRDw3DKgO31xMYxIed+W9fGmJO2Vhw+W2lfZUNPYCZDcGN5zCsW0hJkR6oPg9+0a7K7Sg
VTgdoWPi0vZlEf9gd0Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NobNPEAvOyayp1TtUWqLiTt1wnKf7VjSBi0esOl6kg2wXxaycO7UdL9j1KzK6yLaXpPqGWArWcdZ
OHZWjNgANQMvd87WyNjFR+DZMXSGqH3lTJ+rUOlsySu0gV6nE+CIBmIaadzXmtjlUXyV/oEoRCZr
rq22ZdRXEi/z57ExJp2QenIf48qX0mmYi5gFLdknqEc/38ewzEWm4uHsakTPzO6DKZ89VmneHDI0
7Rw0KBtgnhcNeggKkHBNrVAExbuEzB7b9xOHs8SicGFL9UTrJpF8NFV5zuKj6z6MHtvPDvJ2GC1W
BJO4/x680qEH+0G3sdhClIkA5Ln0j075tcfv5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73072)
`protect data_block
6alIEceMDh0EOO1uv7H8b0zmY+IDdixvY5I+extGoSZkESqrlar0V+MFlDJiSQ12pYJVZz6Q9HFT
9EGj+DCBP8NP2S8jcgfFoso4tpfPO7qRI1Cr7fiPhCieuEluWMirSgHJoEwC6S9lqzEhbGF+akuY
0mUUmWJhmBtL8bM9cTLHsZ2EoKx/uG6wRrXfP1KI336O6XwgIuGrzp8Z2QgWIcnWmwbZOPZbDdlt
ubYfxxKDgKWmvEBlRxp8KPwSt2MgWShJadB5DFB68HEgbet8bKD1s5rCcc10i9fbYN6xnBLTwAwx
mctki7yngn0F+N0r4NHmXYgcm7U8ibRBTv7UbckXobKEBJXR6rSqjSdH6dBXXw8Wwv898qqxbBrk
MWkAiWVEi8HmVTZRZu7lPRUKNINIUhz1gtmLwIjAbddwkI8TExOaK1YQ4/IjE2fXiD5AoI1QgsW6
1eFp95AwLK3nIvnL99RtlbwyKiDlxysMWhDjsofYpq9vW1wqlsJiUZWYNoBpgb1tGyuDcRlUlnqB
3jMvWKk2lgHmCSYoPTIut1h2LZdPBkkiJjFogcx7biebQ8tg1YA4MVHzgZh6BU8MFRyVUBVz8z0X
+hzSnWDxBtZkYH7KKNXcEtXzIUzXDpLQOB5uflwmrHiKOQAb7oCX9IgJ7bwzpcJW/+TfihHOy8pM
7/19VUbtnGK085xFRhi096zZGZrLfr7C0HBTbIV29qDLNl1hDs31XSDAfMJcNtpD1TT2F9494n0Y
HVgiJJEWgUqIbF3YiC+qb+/0zV596zP25h90bF1HcqpfA77RwLd+DPR1/QSQwuhHGltiv+CmcEpy
9UHxIDGPG2zuDSOjYqx5HzdIhQhKMCSTxbXfDhkMz60opG/hZqkDNq3cxTnSixoPz5li8OyRMQN1
56enffnBoBFGhM6794SIwyCZRDK5kghuUQTamdwLoH91CjkS+Yhk0R2RykkPweJypoDucvWm19UI
SLP1qBsw7RZMRaw5FDwlwdhAI2rNmKyjkt+rNu1dWtnWoheQpN6C5KUKDLCQN0pKr6mioOHDaWlQ
UcOBq81ktFSnM29EbWQyr4aVGZyieD4J/1Hb6VsZeecZrQIDG4Obcej5JcLBnoqYHKVS9OMlksuc
ROcFHE1zTYqc+k3pSkiGROtThDp7t/HUC6imAH/TtRf1vZR6pav6Nss1bw2L3R5P5LaamspLC+Mw
WAS0Ll4AqBgnxEyhbac2vOSUHgGsY6Drmocn5QbQm6KBPskdtGSvHnm3peWbL6g/63xnOnUE9wAR
aepYWiZRGsSk3niEG3g9FLq+vgs54MVAoiaYZ7fVM8aL2N+Wgn79VRSvf6lhtgGZoxuzP0b8MTvK
905EHLcDhh2MhI8WnkeUdIg8WHIMDDecxBek2sDHBZeqUGgeQp+qtMRrmUOhv58L/yFi74hIJEVS
sLr+KIYP8iil0ycKN3zBF0wOsCOx9ACie17xBidc4EpzAGWsBj0ToOIigKdtoRsVxO36FsY0/tFH
zvtPBix5kBAmXdLLbsVtsx1P9nwl5ZCM4fGZjy/kTU79IeJ/kn0JYzHvdrD01v2Nw6ob2zVepHuB
FY0SV5Bt8CFmEFyhMmzjc1pv1nPZyuvSsxCyq0cDBxNvCvVN/86ZVD/nQMd3jru2SiSm4reYr0gC
AN8SPkipsk+/ZRd+oQbFObtsxTinBTFn7MwASo8GU/ZJYZixRhFmyAKHyZemSfdta14sdwGqBc0b
8+AnpD1vtEqTGYivktnodIVYbyqVwZ11EzfEoVW6VuWA4WIxDGq1NyRYybO+h6WLU+Tqf5RVzhw9
oWlcwm47Rr6XjBo/C0982+XYIFZW/knNJCdpZHh56YyAswV8MlBVJvlDPVDyVRwxMl5JTlcdSJEM
fz6ZagKQSawNFDjkWMk+YGMHQ5DGZhQPBzy2UnoNij0vx96DA10GRP5Jcs3rpwMJsNZJWRdpI3L4
pscglhE09xANAXUiZ9i6EzFv7ZcFSK/jzWH2ZG4LSXXXJBPJsmp8FWN9istW5zbng7OgDoPA+SO4
Sx0X0OJnIdevXZDQYK4GZJjcS32N1pyYFLgkB784ntn9zgIsAJUnqgbNNXA68xbg5BtbmuIEKcP0
8kP9ocKKJiX4AOBG87KkkQ6sy6gO+GAWDX/Lc0npjFp3PpzNLCxwknBD5Qkd9Hgmifb2Vt8Tmcg0
ttIV8QCgaEKNH6yYyrtlAbpSreXyaXFqMGLDyJitf6J2uM67f/ONvbTPNzuvjr/5f6R9PBq/NWC+
TdbTngJSPdWv9EvjSWnSZJNLrKVowLEqGo8QRDx9/Xd8Bef1+5I/IxXDjBXCgSaIAm9U/WmOEu8e
MU8p7ix8aUrbxKIaiApkkNrWXlIgbbQlSWy1+FtdFmZdjMMLdkR72+oGuN4X8WsKPCXU8tVyWGQ7
xqbUUB47fpfFWmOLQT13j45z1Ujvlm+vivz+jEFKZjMSRot9P8g+mGxnWj/d24Fmu7wstQNuMoNl
FjAHnpgiR97W8pQIzcO2WzKRIB+/4ndZAZ/LbnDncQ3g5Y5QpaJJSkCD4Jt70QJDPhHNb1nF+gAN
zRS342r4CPQShMzhOicIWv0gZYATVO0cuMVUQUr9jvgtBVLiFEP3Xw+JADSahMLc7YoB0QrkgFMg
rdlu5N++y5E9bKWZbF4UbebGZeUunQALslJpdIaGTovEGin1HhLWvL9CkagWCUgP4C1t4/R4HMoT
DIgmLY/l0sYiPCSRNpaoypen2B3XNXeRpt+7AHalWZH66nvtoOePPu8lyXT/7TJ5nuFJfgyPFJtd
M2AuTTXUd89ZDcOmOWIp5O5d/NxVXXywdTLk2fhAkS/zyCYTsD4vPJNDGbnia1P7rTC/W4qU28fi
EA2IPH7VIfWLaQF3V+4DEWWCahxA6IjCOUPHew0jTuebxOMn+k9metf4grsmW8Yh5IyVzQSmRP6U
1HT/YpSiBR6m8ef5AQbnhIh7/Hbi1qtkw+M8BQQ3bcnQJPuemfvRstbZz/F9bKT51DS9oSWDnodq
NmaHNTV4P1UWyRlwMg8IokE0H/Sng+6rQcFYWEAZWZzBsngT3+sjsYnsJmv9KMvtmcIXRpTlYDM6
VF7SJsz3UBKSWMkFeEoFhI5L4u1d6bJ+u1TgbeKGz0FaAVKS5s2aB9h6ihlsv8qgeoUJClUoExFC
SaEPIOb4ErKLfSOdqr6u0EJJpA0juEM2p1XpIvfNZsn6nX+hTtHtzdULhjip14uqYy2fs/uOCoOY
WoudyH2Qcwpi9sX+ikZccUDWmME9ZbTOkwkXpjXwK5W2z7AOAh6O9hGWKE6d5EznCpG3Z2Vw5scg
RxcDLbayGc9hMjzteVqEhs2ZGV4COmQ9BIJfViMR1M44lWlxfAB8/On9jN5Q7hYPBpDyTgwlv3nG
9P8yT4U6Fzv81Q/bA3Y461UgqCnmvvMObQnaA0GFuAyepsWEn6lSopLz2eCmVD/Zq0IdgQ/A8pIA
y4Dr7pRtaIJKaa03de82C8jO7pON5NoysLAUxcTnJBW9FOO/knaKHKwBMJ2CJ4LxmjHkp3zX9B/H
8SUBkjHNqcb/EhS6MCl7mgxB7azdr2SrzvrohHNsl+YpgA9gP+mk5SQwOS2ErvAScaJWpf3NGtZG
YnZq3Z3IQ6abUNxDrMfHO9Q7nFCtWAnBKGHGD8aUU04xhhln1AIh+hpQuf9wM7MLJIPNZkuRmRki
sNsTZIVUA3fBHDAOr2HLBd9KrYxe1B/O4mTDC39XwNl8wHe64Vp2YRCQJays951mJLiIBapSK1CJ
Rmw1/2dbXviEhuAoqQKayUU3UTK4X7hCXSrJYGEzrEqNz0AXft5biBhnnUjRzrUPT+ZQLIxXu+UM
qbHzNlhsZL23xa7pYm787gS0jmq3ia95HaZ3sFtQoALoMt52IoiEAaGszEtwCeODIzaGESRTAF0g
l2ymf9AxDLkrBDMQ/pG3pVB8HCctfKVt0enr6TLqMqXDnRWmPSRRkbn+RrgEOpJ2eIe9Bj7IORbb
4sItBeCrSF73d6qp8x6PXvJ0ln7D/iBBLQhrOafJbk4GamjP0aufLn95km41UsKqqwkptcIbZpik
wHcbCDg1KIJarZDe8+I8GWvWzO5ni+lMMr0x1WtYbdwSxTTC3f5SOlmYRyAqSZQh6X0hhKlRqt+2
0+k3n16RAcWMpYIhvETJCmA120A2ktkhPyzz0HHQE5LmyuV7xzlLdVQVvSMtEFo+GfqAD272z81u
6hSbrmWcSweUAcL1higbFUYIkljBvY7IXOA+SQtMDwt4lMUqNJMlbXAQ+VOVj7cEFHRQpDWIlvOs
v9BvOxWYdNPYS/j3hKrhBu/ZIPbQzuJOM22cIvwrJf2XhFzm/W+c6+utcb1rjGHG+5ehck/Gp6L1
8T2XawKaE+O/SsHlxPkN0xuorF/UbcMkYmRJYMaYIOc5ku6WR042FsbwKjiWBxiA9iZ61YUwZ6h3
FfWM1l4nzmtPYXL+w7u95i/c3lpJG1q2YIOaBZyA+il7AbL3cOgnD9WnCLo7at2Vu5A5MuCLqF41
l5ppi3kyOe/OrfxZbGoipXAcIvzrMqN47Axb4AxLklqe8alwboT/mT1ZFNmIjlyik0WfZSqRtPVr
wFdgkSnoesHAdEAjvx93Mn9a15zfTmjUSd0MskZOs443M38zyNBdxty9BVV3zJBTzaQo9OQG6e6g
vKvmdQF/vLT37mT+FQiWc40/ZHOuPEUaG460/SOGbsIylj+18+wN0QQqvQLY56CmrAHjcQjzNWUe
B++dQi9gfYfkzYyBK63LQIlZNNJdUtOa1pRc8EAYWQCLVqLFaTiAxY7wgsuaf6qK7ofIexrliC6x
Q8AUYJAuPwGoh6NmnHa+1cqe6FWvLy439jeVtuHOSUdq+BjRRfTUOgh6S4dLaCXOb7VUMydMyOkz
Sdu5vhgdLtfk2UCCVcQ+8bYSGC0TJBa8mY4bSrV3apOWvtEf+/5znQVyIM9CaBohBgY7XWz+KjG+
7k+T4zkhucrvfVayUSvtgL3K/LyaEKZQhpjfbQayg027BJsGrE4wmKG0v8QQ//duX8Uj/YMOeyla
JZ4ZTSWoRn3hlb9Kgq9E8NyW5LQpaXT4Ue4jMB3NHMdzmOSFvNuiv9DJ1VOjeWPrvWWBtFGW+Okt
4gfCcv1Bxedz2+fgjH9drFcDVpUX17cPGOaMVGDaRweYTuCFUQZwxPAFWWgpH14T+I6y1GG9+D7k
+pJI13Db381FeHB4chJDGWH1huorpBs6SV1LGjz9jGvDTSH0QIQOxRLEefc8F+Eq7M3yur6tMyA/
tfR8EZCt1MaCVSMSeQ1taWoP/7IsuL6ezwsh1keAhhOugo97SPF+sYmh2Jw5IcBLfqzNIXc0vK3r
7UveXQCKCJLBQ6BrJRXACbg6vnliC4u8Laf2DA00WH6VtRFflh+H48/0XErn7dWYw6QaVWQnnGS6
8f3LWVQs6ikiPaDkFhbngYdluftsbnaH0l5wGjdpCpApQ6FxpESusxPYClUEUB8gwIr29qHTHMXR
i9n5JHJtIeTYCc6Tm+VaImDrkw75Zq+RdVGCS7paI5MYj00HfPVC4W/7Lw0j2kwIExSpULDiszxq
+Ojs+h5TGhKx8piCpkO017AhOe5MW4HdbgVGKvhgcVoiq2o7lRdMY7SqWIBhLzS1kmy0Tg8EyOnt
AHqR/ni/61cBTjxa+5bVqgi63cBIgL+He8Y0ynnHdOItV5bzQT9Yc6BvmI+Xcaap6kAuJ8ToAosw
Ozcf38KRdeessRRHQ+9Ruil545ZSUmNlAh5E/XzCwzsCoKJdCuVQ5uYOa0mvTMBiNnTGQP1/9u1N
m+R9sPRHHA/x5RmKbnz6ntT59ZW3DQd8Mm3VFfMb/eSVRzW0zepi3gxx91nxl6K7tVhCcN0nYF/4
gc0wKvzeXzp1RaGrTksseMj/G0QMD4hb2qh6/efZ+wWbN72X9MZ8XMKjIf1vgK3pIM1aCXdiDJ90
HOBkwj2HRH7RAGG0jaO3yEeWCl0HsTJWQZVDds3f+31PxbjePeDv6Lve6IgsaB4y0VRGdx5uVImI
Xbb2iOHcTJTwfxiqpPed7JqYSI7vJFHLLmfgZufUxXH56lQxwNu/HB0uiepe5J90FQQ6NDAWrUks
NxRl/kge66ClnuQDkD36qwXbv1wKmLIrQn6nK/a0ev5SuQD7V5q3yVT2iWnHgJDwTgOZCsEjqjfu
xMPt498m/VnQIOKhkVwEnHB9WaDQYzbno0C2SmUQgaUcdZO+/aduyRn+G4aWIukqwnSLZbokwZlZ
QBYyKnTxzDhV/gudplNshP5PcraPSgLc9ATFSuhOBP0ZBNgABXlQ10za2x0Al/PG8lRTUmbkdeqO
KTdOmJKeU7N+lqUrkoNcSVMS8787JQAUEc9p6gUZCrYeKLmEFs+tXVGbFJSqfjFk8YN1dZjK4yrZ
42O1iSo9fjJZ3CW4QIHhw17D0dA4GSqinss5byRZpe8glEYZQrOzWe6lnYNj0pyb9Ta5csT5Gbzd
Ky1ujJqrpCzAZw9aTkCpx1wtIuwotM/XNxwBOIPeEcvvDRzQvAGEjeGkarE8qE6uF87xc2tcCpdA
v7jDvbiFJ4aSLcd9r69aFXniOuZCkGIVBYVpc7ZfMz2wl6jqQlmEnzfxgSics5GIYNJCHoa4thhP
ooiUlFtE5iqe5XEc1DvQnZxmwvpvy6xk4mQkVLqBO/U6HXdnYMfGLi2YqwN143AuiTLmtrMXz50F
btUyb9bl5FTmedtE+5HiTZQZNrut5NzrpLsXhCASG5n1yZ5XPm7iqDBRmqqISBcym1/y/igvA70p
DCVNsg/Qa7uJ2vm0y9l30Xgs3x9bTMhgga+vSf5UAKJ1otaflGg5D5gKJmeIITh+h6YS0obFVVp8
MrNzOi661hfzknZ9awXmNsOZj592U9VXtW0F6dodY5/+WL+LdWo/S4CkRAGb4q7HvEDQAQYqRc/h
Wel+39cK0l1e0pCoTG+GUZm8L5HKlaKAmg6/h6PlZHaqV6+/TtZV+stZi0EbqnQXN3FFdZ0Vhjxq
pCjBDsX0bWMmrscJGGEVdzIXhAqoe9rIfC0fOINkxMkJk3gLmjfL1GBwYnORw+qCiI5WGUsHmygM
ujey2LDL6LHvdL2dqTg6naZ2hZRTM+EvbFGZUhYktQ2OqZJ7I/6aWePSiqWYptscDjx0WdXKaJEL
ZG4Q2/uh7DHFO8eHlwbKtWHdhKiLPmUDcNY1n2MWrU0XYO+MNSZqCXe9R2T5LTVtwJond09tTaXW
U+0sBBtSsCsCbCFuYlVVbszlpAIhgtHldUsrzT+bn0GYGk1uyqb59VX3i1SGMrsDRC96HSM2OGJ9
KPGxZ6FsSeayK9SCUTqLCfjahcGNitmu8uXJlrpwTM3WxoJXIqOT5FD8x5t6A4gEfmbgw8kh627x
eu1GqhcyMfyxaDh1OeVFX6ykDhmKXz0STcePxI9HqUO7qHfp3gRqezJaq+uvT8tDQ0QQ8b2tAhXJ
RQ6EpcOU7qfWdxglD3lktt+4RC5qaKK+RjvifS8mvljAhvhw8CDVDw0nLLklJ/DhTXtZGxOGFIiz
k5D0UXYP1Txenn1ODMO5cn/0BP5MWUmANodUv7Spah4WPCPLPX8meRvm57z8OSsGdL4o/UFzLK8g
y9Zwe+lpFexAbm1YvacxM4mg4/99y9N4TM+lUjTnyOc2dwkJn3SAm93/btDRdZ/1cfV/wWbPssuj
bnYVkIyedaj6I1yJo2W6K7ebh+KckD9mCW9x9ldJhN39g5hANxmF6G85QDcKXSeSq3tUBGpeA5fO
4F0R1ipIzSiAPU84BvcMh5zHn++r7UlfS+Eschs0qtsABbHQXF802b3VdrmbJWUptCKR6LMEAgmg
BojKTtvugKMzdDAikAbqSDeqk39GKwE773OoOE3rJI6RLbMR+n8tvjr2KUfW8zPfZOWDIissigiy
3LKVSIgrsVNChge5TbNNPmGPnT0wgpb5Zr7X8/EKlP8h9H1g0EoGPuGiT+Cdwsj722pzNhkP6VaE
MGSzhXWt2BVvkLOugw6wxJVEwLwsVqvNT2jpDgsuPu8LgpWR2x8mMXq1nBo2+J6gKo+m0T2Bz1DF
L07KwDuU861mJ+ETACQSubzTbFBhnplCQi+g3eJa7idrfKFrxU4kmDuPIlMCyyskVaXqFGpMLE1S
UHqyLiAnDKDvbXJSHIaST00aI6n31DHMRB4UMjKc0CZCadf9hHgPuV1Vt7qV5ZyFzmnEAsVTx9R0
Kn8D6wtCistm91bTSEUzD3d9xfGe5zHUpdtL5SB8GxoIPfGwSeclHoZkJ1TmYFpvRfVwsBnbrPnC
D30a/MaSJWiHHETXSEirfZmjYzjqOQuu0d8A2yu6AEGwU1BxDIHdEmOlkDCDnz+8Sa4MnpB1qj2+
b2oLeMQnOt1Y4rZEv8P7jD7SeA8j59RKGvQzBgUeIAAuuXhj99RuEYXER2porBBGjGNpkOjTJaZP
G0zj3CFPK/CyYAcjHGY4la31JX7K8WIKZeSNY1dfN6pFRMhGdCjbgxpmIN3HuWGcWHGrVIKzS8hH
QcLSCRz8Y6SIV6ONr19UEDvZd4iJcqYEMieZ0B8CUMajbK+sJltbYYh6WDx5mtUzkBAcF3F/0gxm
CFW07dTNx6BluQ4iivGJ2qpCMnFMnfqwkaj6Ymk7unWwBiddSfB4heRzLiwta0C0tZr9VbNmZ1DK
0X4dsFD0RZ+KGAx2yNI9QqurS8VzbAf9ECkneAXuy4JfuZDZEmkJYx6A57uaFFQYaRDkTLId7lty
hSBq5SX4IDZI7cvSbfS0R5K1ATYOjvJyd/UO1MH/HZbXtDbWB9gkKUjWGtxjI892rXjF/NeuDLDi
spaFsVz7D/51u7Sn6CZ0frBtKW6b4of54YiW93FUwbGsTBk/VlS3U/SkIVVIDAn0fbu53/gneCd/
YiPG+eTL9XL/Z7W1cjovpKcmSdqmxzPoTI9H4bIeRCyGy2EwXP+XAkm7wQTeFPvQO8G1dsj18BRU
FUEK4zyv+D2MUjn+w8d0Y8oRmQKI6oypxdj7zfa9JGluUyQLdgqJYfk7p9LMbN10evtbtheHrLVz
fxJm9mEMBSJq0XWcVm8CUz9SQI2N83KIpw0L+IOMZDczHMUhv/l8ZCLXjLBVXbDvWfOFac6Q6l16
5GGXx6hCoJHuwrEKVjBaeTu2k5+vHAy+uQcTbw5vFv8ixfnwcPZxcNCDwLOLZ8Mwu1CwrCY86wj+
bRITrZndncEneenDgpoOH8tYQsEBwQlpp1PNZWY5eGGD1IuADUF/dJ6i5ZucMBFys06pO2XGFFkK
jfXbMQ3AZ4hN90KSYBPc8LdsOlF3i8j2XxGOqvjuEiWAIxf2U08zshf7nmecGrgoCh4ifcza0IbT
6yPwINOHUVUyEjh9y4HIrqyMf3oftYrdxVg04vTEMjkXax8er85gMHBmD0gmQSFysoRsd9iOYgTw
6EtBl/0UCd3RwMblXa+QFDbUAsDA6y4ZXWwyY3fFcscIXgP1dCXl2B6JC49KXxp8aOWmXOikKunr
Xyr92WQ/QsqKU3k76AWuG4IT+PGswthVaLEQUJV2jYuIFHZZNsy8P1/YuTGcl3KZfox9uagxyCcz
NKbvtma+D0/NpPoCqoo2CkRfemThAkhXtUOR8EaHvALvAsKMgr+nrmMfMSjC+QpLr6b0M1ZMTGZF
lrGCg7gr1uSVzoIEk8AnFjwr6uu52kiWCgMPNG62xnhEqfVcgNWAKzEBpvqlqH/Buj8NWHY4fPWo
DLqY4n9MKzLU3fP8OTORQmx6IoliKhvfdl9Evx19mNlec9bD7KuYa0Fg1gxjz/smgOksHqbKSSYb
VS6KBoqK1leM/1oV4LmYpyoH4qBiqYKXigQRwR7aB3r9ZTyvbwjJkNIlIQKfgJeDrYugklNWLIaL
oCJko5eq/osIT2fpeFpNkdAw/1/pQ9XamxdUDa/s+Vu2ebVtxsJpK05NIbKjKfFEW9PCtOllvMaO
Ogaez/7HrSCwMPmFvW6ns+hml64wqwTtp0A7PdXW4D/ZvwVfurs2o8fpZX8oP7rkTBnKseVRSnCZ
eKgSGL8pUTFEpU4O0GCYu2IMJFpeOaZLIlpqrkMK3h1a9xMB1V3nfH5HYJZAn54npz8JJIZFuAcW
FSwv6chYwwK5x6z4VsN6ssgPCao7ivXHXw4UU6h7GmjX+wXvfgIBWbxNQfq+c75EYpYzGJngdlAY
4PguYEdUCtDdd051x4lk72DcEwMmabZce2ynkJqsVCULysJZPu4kg/wlh57CrgHi+prUV43AByFI
f/JGE4mRE3wwoiJ0zhg4PolC+ACLjEsQgnM4if+tGKyIYHcgWZzxZBibBcyrr3DWfTNm7THJfeY9
xysUJdAuTRpAIGJOHI3j2FQlLniz385+mrUY2i0sEGEBJT5vq9eRVDW8oIt33PyEG7iMeuz/m+lK
N0Ej/jV4Lpye9EGS4jyhr9AU8nk8pqx0atSf5ONoUULkAw4xN94fvUScvjHEndX0gFBuP9mtcnLt
LitLEHLrUrOKPKeSQM0h4f1PcbCAEIYWiU+BdVDz1uGz8tFgw78V48EZYIZ9VySMSV3UsQmmJNvy
G3ENKmaZsCPuI9P5qjmyxm10j80Hcoqw7/WxoUdzEYBKk8wKZPMY1cxWScuYeGAn3mOoygL+K1JM
MA5NFBuxpkbRdroIbAF9byuyk/AKrSIWnHv/+x4yM3AhOY2yuNdDjjTu4yVjfzHmtbcRWtO0OeXS
A6u3lU/WuTlrwCKUzu+erVPlcFezai5GliGrteKkH9B6nkRQikeAvT0AagrsxQ2aGAgeK44ni83/
rnGO934MTvhboZv2YPKxMVOqi+546aJmQ5Wcw3OQefoMkdrM2dsY2bWyb7lHlXTm4BeT8Rp6PZHX
9KXTqXGIqpu5fmoG+zKJ8LNY4oIX47flB3683Zbo+rIa9W8uFfFjsMvZKg/gOriDfbID9RpLBBWO
0wHaWOHKioJktYQ4ktR16CFJggrPMYLUEDEd+idkbSSboRYhd9wQG1Lo6XCgvtUG24TXioaI5AdP
/ODgOR/CunGimgIuU3H7i2lh2jkfg9pNVHvvO3vSaMRAmTr7O7C/vpaF1+7gtAHSdTHxe9xfQry4
0K68Sssf3AuzKFhziduK7+NxZ37SbuipuEYFGfenij26XLhjyrwb5QKOHB1WY64BPoeQOJ3e7xIK
aQrs3RZTMcwj6dIaOjVOcRUleGE7qSSQCJOR3rmn+kutfYlhd9kTxNDys7Ok6OUgt4FvdmdlX8UP
j8bPEcAIOvryp2cok1dH9OTR3NufUwCClImljWbAJDMw8mQ3n/DnYdPBkVT/PCA2lnPmeoLuL2mL
F6S6/8SCTICeHUfpC82Ne9cNpoFy8VkaujG49wyRukNpVX2EQAczYoekqnySzZGcRXZILaTIBces
ihhutbeZ/YkRkWPnDlMi2MEm7PjoJoeClnavNqtlyISnBwc5fYCYQe/Gk+8x7Vb313yUWWbE2lrd
YCNSNle5KoEJGYfwLMnV4IpAZDMphN0bwrTAM+Bqwpzcbb6mXHrS7uiGVEAi33sDfJ8m5dmiBoaq
60JPPOn9AZWnasUp3tcjRW9MAwhWk0F3rsbisTWoajt+HaJdbKBz+BMYWBc8TFU9fnXPoT0dGouQ
9g33HuEzjgWp9sGjwt+WRnf4oXfF/yT0oHY+BowN3X9TXefD2NJry2g/Vhs/tn72o+8i978z07B3
Fr/4kDYCyZBZ/iBGfcyFLnMqwxHPhAG9qCZeYMbxBTonU1QZzPwv9JZKXeSgjlQWpE86Sfln+f6u
QhB3mLhblhZq9hWVrzQ9dfMnq1K2kJylVLxm1qCPssEHwcmM16f7LD4dFveByX3goHF2orGQGTeP
97VHxL2hBeTn/ghC0uOE2XtR5JIYsQmGT16Z6aFGAPbKGcCYuAOwoJfVtCoMjbtIJcFhTg2JUCbg
oUnXZCOVvOFC5GQhHnizRdLCa3TvFx4LYKGZtzpcEKNAMEIh39W02iEh28jUtqJJucU3Vnw2C0d6
dMuAwu6HO62UZ+Pu+r6kYh+OFgTNNAnZjlCmz7KQHMzaYkq+cJtyeFDI/N5t3Uh4NrpSNUqqOaW3
jRUmmJe0S2UndZHt6QW12EjOhIKy2ihFau9vydiHB91AYkJtkOqRJQ4jVB6KbN/xIx/0uarBC983
5FmmrXR1w/3eYbA+Dv2vooklyUy64aF/mqtZ3KBxROUsOxBsb0OT3VGeilG69pt6Vf8Am7hRTSCV
5r0Awo4wh5MAyS/+jxAZQDv5vHobCkZqtbOUoGA9YA8chS5OlQW5Zm/VlLfozyaO2j0CWWxGRd+R
VZCmXbo7XBfrUGwLgeuj07BGhoFQBJfsyrpyhg7IseD/Fgv8IfFrR88Ze8qkeDbQVSNOxTys0pDH
snqOVI5HWN7UhQSxq5dUE9YtkCxetnfo49OfNbHTegshdjE4BeG+1LOSrP6cEvoM6aXWicstJaN/
vfc9d/ppaGrGWh0eKqbdnXVGIVkLtjM6vWH4HAdghFS7i5yhwHg/jxNAuNsT0wlvmRvwkxBnNupI
tDRzdsov4p0vTHcUETA0k4OT3hiSFOgmtbx4ZX8QPHdH2Y+wKD1w53ABgVpS8pjOtelWoNOkamvq
ZLBkJD2cFLsoyT6EpLeB61woQjRNHD3IFFaIaBNqUY4S1bEeUVUtMoi7tVpQPMhdBICunezC2YkV
QrVfSbNkmu1IjjpOTeo/NVy7C8z4ir1EXP4o0mPE2R34yIKVowmu+0E+MzkM1ihuPRsM/EIVgMUY
Wl5tgcP2ydzf1bPZsiIdIZAnh/wBCas/zn5x6cAofbQtY0ojZKRxZJMjP2MuVvu3+LxZW6Dux0uR
b8ipnEsBccw2zCztQqzoXVlRrjQZfeHGWqMVnR1EMgfP9PCwv7Bpg2HaSh0X+R3NX6jTHs1c6eDY
O8nIvy7LYTnJswuMdOtgjNpLvkjAzuZtuUnB3/DSdXrKB36p2CpqAI6SrN8s+0jiCZHL3xpA18y5
6ABOQ8KyMhsLfRqIdfUUFybvdfMLYj/B+D0EAWslbb+zod8GRTRn1i7J7r0BZTtt89qpujAkun9e
VPM7N+8iOct4xzz38rm3gs/mYN6qemwFSU8Wn1hxjeRN9utftVazcMplpgWZmrv6JH/+LhgRBJG3
jNLV4oFNq1/6RLqB3NEmmbGEHEsk2y9z3lBrzsIrixcC4Xb+6ma544TuOlD4RM0MGlGfvl2uHKQN
cQZ1mWPnhmrzvvCruuoWSfKMCTWcr3RSridDyWVhjd+5ewaKzeaKDCuCb1n2iERpaxs9uiUZaF+E
44xd5RoQ/iTI01x/fMmgQVolJkz0g0wWixIhWfo1S1+E5+9NCqxvg3m2YDcmsha37xr48XWm+Hmw
LdS9PltwXEjL1HPr0bNedhpEyM28rtkrJZfMpmjksIQTDRAP3RmXigzYatCZEc1IWHQQ3Fl0z61O
pIQZB20irNITNqivBPJWmV9I2afiyyL02VE/qAHZ+Kks8SjB5dD+jkmJEnignwHEEf8Ez8uZW14G
TA0TwMWwkWO5fLbm5YlnYqEklSU2vdcCGbts0qcLeNg/yiE+gOeIqOjLFtmw6eSubyh5kSy5tYPr
FXvxtqj3373SjN0cwFmDWIaVCA5VJ3tJSrL7Mi32qmAGigVHMj+79YAQsQzsKng6ECbHB/rQIAcH
OJsT/w0w0icBnVCvL771VJfwTueuIJTmrenxqUTijg0LjEXG6vLYLHvRuguwL8bi90FY9ZR3vQdF
yfWsJIeGScNbDRJLjYJyn4YsHnTT8vCW8vDTjZGxdACyBVbAXQz4a7lq4AYpO9AGyimToVoxegXs
Jde/Gt+XpoHQTwidK+ZwH/D7FRQGY+Id7Mg311LOziqvIthLvtIC+KO03a45SNUuKaliAD/OVkwi
iMh/420XYkxBh+vLF1ZA+USPg60h4BmCQgn9XoS3YRTx5b/4NeXi6auuA8RKdV6Tx9DVNMqhFp44
8PA+8iqkudRPhqalyXyRGu+dBdP+ipgj7gN6yvD0ZoQdfokH5cvem98A7mFRKwfoN2QLPM94MgQx
gWpcbVakj+9nRgjoyyAFG34fUW4DTmSurL9QO7Tk6uhmfoca6xkoeyGuSN7GF+UZPOmorU5FoW6r
1PQa2zBw+5mpxTtCrGa65yxky7C8USeNTnxCCP9f2lZC532n6/053mH/lrFfb+eRFFTOMVqYXdDo
z8QDJQRGx57YTV9FOBFYG3R6TAOUHWxwFpH5jvid70KalUwqcqH5dQ+UCHezM4ADzdvdDY0H4Ft3
xajrq32sDhhcKPTA9VThK9cocWJJdYqsqFfH6ngOapC1b+opCVa79QFAeGX+zbEQ2bE/2SDSBSBP
VhV15cY5YCYa1xcRaIYVt8cARi5Q+TVal+3G6+7xfbi2PwD00f0+2LwXgSEbzmGJmX/dzTsjnduX
RaUec+mgDxeluDW56LjOZgGyTpEFUdaqQV9ht6XreHUHeajeOBYhUz32RjjFg9psJH9iuZcgjiHr
yrpRHHtJWz076v2jT0sb39Bav6OMeKY9omPmD3S/haebzJPWnWr3DJE8IUbyTXJaQzzLFdXer41T
jPbkiw19BxgO4TUCrEQKhEjnvUBcDn+k0dGTx57snNkbzQx52ztH+2WUH5/vxaCUOTPiuMU3oRgS
VlZbKagsyOt+G/uwfjBBpKIiz3i4pBwFHkEeAjAx1AuT3gueU0Y/vA28ceOPFLlApXqZ6GqCQLKA
Tkzi52aFBabL+ZzcyI4jiJXkj+ZA5bwY4XAHQYb/kHLT4GpSNIQbYnv0UQqbX8KLyKG3XJAS1hE8
zCAobFJVmKiSZQm8xkkhtavJzgNL+yPYh+yX1aJEQbAgDvx1V7m6/ajkk5D6aVU626LiAmWl+pi1
MdLsCq5PM0w6o3ZAs4Mprr6L/vkogKR15+I8HlO7wKzXNzZnq0WcnAV/Swsj5K1Zdeny2cNh6NlS
tcbktACNQehtZ17T0akq85QqIG5sFxL5r38L6NRBn0zV8uoFkqTrBWogi+kKlE/SmVFwBT/18dJ9
wflcgfSL/5x+eCbmwi/yaNwJx/ubCEX2RoZdGkHMLYnTd2cmwvPC1LyrYCJnnvqPs8wXdUPBF/4s
2p4RNPaCTOpj71OJ0XOK00KeFVxmBxStRwtU7gS7Qu4tOtCZizHuxgma8TldGCiVYzyw3s/4QQTL
3s9tij2Fmy4m8Wprg+3t4sqp3k8uqR5O3VikYn25kAMRc5HugmKerFaDca3j2Yfj3jOxNzWzJ4aG
kl/Psct6lP4CD66o/RlGKvbanS5twWzVbESFrH5CTx34XyPsl2tCBppudDqLSuAG6WLkl6yTVJmt
AZ3M5OafRUYQUqO29Z+yP7uf2UtChTwLnDk3xzwLYspqFtLwuJ+55b1uAT5XurO2MzgXVsFWKZSZ
af7jYq8b2InihvN5HqoF0TWfWajBucbPwzcyufGe44I210WxAv+/8SpCbKFaG0PEeGC7WwvvZB9L
a6oMGE0u9uNqIV6tFNeOmVAK7jjAMqgSu91xfpRScpLISPK1wiO+wzsTeXwJoJpX2BEZ704hOueR
j1m3UDismDnnuxHYHNzUPmTJRIVdqvU1hzlDpquPk/4Ejugp1o8j9SGFnmEaMyXwEG599bpEZSt2
qNrVXuQmttkNSUMFdW9FV5w/AZ9/V/LQaFBuQF5kJLry18ufehM4m1hQUDk+ykpNqhAENdFkMgdu
BW9PzQomNAbNwFov2u/OfcM7Dlsjf6HUPI3owx9Slr4FAy/0gtNRqlB78bmJ5N97odtvYPLYoHSt
cLsxWSYMgDvTfohHHZqJsCULrO716D3j0R8fb4sHA/wbfMrGSxT7Cqs9IOz3sVoogWWvUopULf5x
GQ7rNz835CAvgbCN21ocJ1kYfGCMLS1p5p5BjQt27gNrdepNX09CniQd9i9oMv24v3idRVQctiT+
XMWTWrJ13iXPVuiAhNP2NHL2FgXP+Ys6vE0vQoV01fp53cSaZ8Zd0OasKfM8vJ9K++L/+qIGec6x
h/d1FejD7X/oT5RDFgVtO/v6mcm4JrbEuIRsudNrSLtgh5cg9h55MWDJu2ZVKgqxOvfPlqN7OwYb
6g8A03nGyfWujBBVg29S7Ge64c0jevtukvxGPayUTaZ/2pAh+hj1fGJO3AuICkK+AOeTNbwXkdWo
nlU/iJgI235wvDFkd1Z7MVjeqOXY9HEWxWlxctKF/wzYmZ3bN0A+KsV/8n7D96IpBGfFOAuMlDsl
NFSsQbdYZUu6XT2FPNwOQ0ykn0k+K3aw11Cnv+P946AWqDZv+5WicFOdeAJ0sdiP86B9Ym7bWWR0
WVMy4+UwZBKkvvac6H8xeL3jiONBbYanbdzCjGE9eKNjfno8gAKtHFQ2h0SA8N7CN1ABHh3whyT/
D7m28PRgnMhS9pHJQiFibfWIYz5aUbGJT31hL1rMZr24yY+yQoYzwuAkdlm9dwVn/98aHKQRNXdP
umsKxwe9p8GKqYQpGbMVq74ZFjPfwejr/EkFCAChpJVPlLHv8100br3BkeFnMp3VQvEr4TYG8hh8
xU2DunVG0+RfqYbpN09b8EAU6VbRdzB7biJvp6Vt2SxSBJE2kK1feEmM50NnjyxdRayEwajQmLQt
xQX2bBbVEXbxnAeZfNj9Jh6Ang/43dygOMzL7AGKCrJaus6EVBIpkqcSqZB437uvABcIRnuUgF7M
Lrmzoyr++jVSK7+qZ2kgDiapc7HQd3FQ79Z/jCmxBdZF/Ko6IG/Gy/AGzyuaXWm84TjlFHrHYWtL
jJor2aTfQ5li+coByidC5AKm2+Q7ZighN3/o1262Lsl8vGJRMLJazuQ2l1BzwEuVtw+qc9le/tix
uMa/dEqZNi6BIYF1bOkvExmeFmLr5/lxxsiUBs0QwK/IAyeeBDY0owouDcuOX9428GY6M+tFFwwj
g7MYmZg9QfkZspLV98fBj5tjAmVHg1j7GjEeG6JfSWto2vb7iKhSdRXvd2yRp6v09ihdG2HynGt4
t8Al7XZMvZO0mu2dNquL99nL1ZRzwN8U2uCNESdAbkiT9uJit/9/ziXc11v3hbg+ciN5+3DrrQ00
rJD2SjymLs0qfwSxAR9+zRsTjWIL3XinkvK5VrKgHnVSS3SiuPzghm94+QuzRMF3GxH7HcFB+f4i
iGh/ge6/23gULNK9wPNp86xjc0ftwjcd7Onus5TbxZdVG6Z9iz+l9NAw69pY05yEQEWc6kZ8l6xf
8T7WCo/g68vG5z7wfPBlbv2ls3JQyAJ5J39wPTimm4yZBIcKevfjasjeYsxUGFvwPGRElxJezNzV
i6yGHqwvcokCPu+mTUyslDV/tVWTlfLgQ7+EKPAHfFfPYiDt5o8sdy05YAN2cps2MwTYCX+tte1W
OAF1VE9wiFyfvmqhTn84jMa1YOlnT9L6yexkDoYHq+/umJaG3sWFoFb3Ui4yDVEgInPOm2UC31PM
oCmwtnA29zF7NGObc7+RENZIQilYNucD27l0vawJa5llvRX7bjNMPyH5WbMfYG2TxB3vY0F1uxwO
a9gwo6NwzSekXw8evtQxGFFHYr/GYzxhyH/477/h3SzhXFVSHaDLU2mmiw9uIelXKyq6UzKCkV++
nj71OX/nSq031+NZJsjCanjWN1f/bZ98d/lGrcKwxJW0lUTJ6FkcXRZH2oHexrUivzyWoqSg68Yx
YgfroJrYfyb2p+aifE5Sfm8svkXD+nvR7zEnEOftjRn8jfd9zVvIW8IUMccg8MeqHFENoNOUmLRw
FAQPFyVaL5L+PgZuZs5WTxS0SMB1Pzid6xRcDVH90QXDYTYtAgXspK0MTsDgNTVmvC6wPBUwazMP
YriN5ziMCU5eSqTwnoo/CJE43TGr02lO+rqi/b3CjMfH8ct7VyqG+b9nd6+uPIh2YASNmY65DaOB
BF3H+ibD1HgBbKKR6hd9u3jO/WOlZewuHpgIN0y5idiP/lQQ249sNQd2E4dkZgZMxYfbL7BBYWDP
CmtzIu9tKbjygVCXYlJrgBDEGM2xxHVPwwjPVESGRu/oAG39jEsgY4zJ6NZpUmX/rZWQxSE7L3b1
1VIJWz2F7eUCT/wTcL/CklD9RYPmC0+VesFIBf5Bvp/iD8KgzRlgQyZXg/L764QGUKFRXdzdEKGf
zdG1IMywr2lm/oGjUx87YYee25H9llQWGy0IKAIC7vy7xxRoHZ+Zrw462TTNQc+8MEITO0H0JwyF
BfKxJ5Q0nbIbkHwX7jTS3AhYE2OlIDinfnfBll8exojaJFKLua/TDObu6ofiGRxxdgbrIbYBb2tE
NP8WSKXP5c41DtHZnzNBfu18IFRJXeX3V4xlja4gWwYPbjDSWmKZicg4V1P9pYE5iJwWbanjxT5a
Sp6EpZe60TjB0OLEQIxDPo9Tb8KnzwdQbjrrVYFPTagd5rZEbpKg5HQmSBaCBbPar/DmEJSfSvyk
QKl1FYIvebNeSITArG+pjOjn57cU/FjumtrrzvDucs0UcQTpeNVtcA0P/a+Bsq4KO/yCf7+ZbOKz
GM9Jfy5iOASmhd0gOCbP+bvURhJv1dvhJ7KfmU8kFVnI7YvMYYxXVLjlTyOFz/I3QZXhNH+zX77Z
EqEydCa2H6KbS9rEnbxeEv21xgG44CBU1t084xm2fR0UCMJgTB0SaIewopUhZCOvgmpzZ0go0ob2
SwunBR8om9i3qwUKH4LVoWrLWP5SIRng6d8sNUBfeGOb5gAnbiWIPhU2dL1fn1z5mGIMLja+qXe0
oEd3uOQWUBdO6N8xgAGmx9j9UBbR0U7n8TF0xckzmdBYO/WUoIITsdVVz6itq25wbk56VzNu2j7c
8VijOv2viw/pwBoEk9goN+IOHIpJV8bmSTrEnErSSu3r47t4jPerEhXPcd1MKDAjXaD0AcEVc89Y
hVS//9+4Nt0pSCv0NIdVVjmoDI8mHrj0egPxahy0UfFIRRK40AR9EjGv0oWEFVHBfBqfRTp4jhDD
LSDq9NNR2oxo82dXwrnGTvJHgffqaPNOEYu4vX5AbcZxbmjhMESx5ioMR/qQs5gdoy4RDb5IYEyT
96cpqHVYV5ymPKRKo/u7q3GROAnX8L2P9LObvCH0I8gIDUopznnsDkoOnkUvF19Yc6qRPDcQomZ9
pYS+EP9bOZXLaAZ5gTdKTWKGMDONzoCsgcSAxd1hNcXVUcR/tdx/hli1wewegt19ZxYEX8CaEvI7
Hke7l58UEPSOq0NN0k6xKa4Cw0m4eyoSS8hyfPwknhkrGmhgo73H6MRNAYtnJ0wQo5JzqrxPdxqM
m2W4pdIbDEF0Glool1KXlAgkWDAG8xWp4PSxf87wEaw+dA2b6GGVFH/66fyScV0dX4n8e/eI/2uW
PRyje1vYyJXLA+6OX74cdT1T5lzzLsoLdshu2sWM2AAMriIwL0qz1wZMK14Sx57kQGw+00Mnobl/
sKDKF37tVrX0Q+Dh1MWvelhBXwmnFA832HqJBcxsa53Zt+uNNamwear1+3KeIAqhh9xWpDpHos8S
HZpDvgpaAV2OH2VZIgU9GahxunmIBDLb9v/z44l+dtgoOiuyW94V0lAgUNwmNZL9vEOtzwe0XPJO
qctfAJf45kBTlIH2mgPOLTK158KCMbofuZWdT0VFg7s86xPZLjvJcncAggujIXqbab0Ddc6AZlw/
yuXJ5j9i7jgIT6RaRfk3AlR43J3E5hEQlILBNLH4A97NpBLBoiU24P9gEHZHnp+vFqD0oYzmGjpH
huM9NEfNnFxWZBNoECpHzNHFd6e3TAAyU5zLRtdULlf2A0+Hxq8TDqL9SVokuvnCmhEq1YT5/lbD
FY+fiCyQr1HB4IglvJTpLAy+AtFzfPDr8KPdAjYaD1lVVEk/PoB8TT03h7+raBzexekPQ85Cky9F
JVMfPHRRdbtHHqpMixD2ieHGcjU0KbvKNIkUS47MmifBHVjqIfiNKcgx3KuFWQU6s0xw/gyh9CSv
kYK+4kNWhuF1iONOviQj3pOt9eTiNuUgEJ3PI3jrWuzutfP2iviWe+Ov5D7LC8w2I2Vyxmh17+Sy
eD4lNoOcMk0u2do6Vho3shFwoR/Cdx9FtUcJ+owgfcL0ZlN7Ce/1SG/8FCMI0sVMqNVal99Y/xAT
4tZSwgxig77swybdRX53HhnRhE8Rf6HTjKONKzjKk738flWYv47mFIHD0cZpIDUIDnPbC02cJO75
gidK4et/StfHUeOh/FlWOZB5PPeQnjMVDYmR3xOWaCJWEeyTYW7+ZN7CEb7uYfnRYx7+FJn5dNbC
j15eVeZeHf/cmsOTQdIzTfT9LWnjZVhrdx/F+8Joli2kWgJMQ8ByO+Q0blOoEsNDINCNpREp10/1
vy/1sXeQw+54UtU0HRq8QfxoYQ1QkQrxjgDZpZumnGRwELXWDkofZrB/b8EVGI8MVNVb9OC7C/4/
sLrjD+LxcSYVlwwrYmQIMkBvJXhi/eSFGw50GfiC1/NHFLI4BnIRcoZTlbDeEdg7e/xPud+Dhyz9
DBaPc233iFtwc472hF8nMLdBeQsNxha4J4G9GdVANa4HyP69uqOKmOhIXFZFJIoOJlh4EdM0+ws3
fJ+4/WWDQTjp7HyePjS1vvYbwo8/OMFY5SWfadgQrvvr5kBsq3DILGKomtLfUQK8svgYpVwOcty+
8eW+4nktynkQMu6a0xbTFN04CFogEQ1qNlGWk3CRIRw8lZdCOc1F5ebQaanAwaMXkqc7X7X/OnQw
KkI9FpffPLnhfd+Y4sYPhXouRdoEDDcHiTqInDs5gkLXf84kYvobO992qYx+IP0U7Uj8Ww2pXlBU
m3FYnulpUh1R0RMJ8QetJV2yKxIUXbEvAeT3sa2FR+e7+CzJevqkzCApNoL1TNAzNG3u0e+JDxAs
GyTabCOuZ7nRnvwJe6RarIwnHRi75FP3Zr88dadAAvHDMrAzHyJyDWFMjm3YQqopZ3uZRxuULLLg
iUbaxlb1XmvGkN2VpIvrIU0K/B2/ar0YjfiQyYEmXmCQIOZGf41CC5aBqdGobjxhPlZ4f3/6lRfZ
R7kWQ+KD3sizhqHXYsQcrgA7yB6RHbOKLegzaCnG2JpoJLBb+QUyLgeJ9G0eQoAaq9FaWvQVAOP1
moq4Fl5mbQ07BgZ0HNVYPgOLTsINGDKM+RRnZ71dAhRNPVzoYgJqB+e4rymjPS92Km2LY+UwzTAh
ZzknDUZUEHsX5KvVhmP7z8sR9oWGsbNvYKh5e9IICX8Rq/Z+Lr94rWWaMZ8y19M+tjOxAd6v+p+y
PBm0YeGGRqqZZZ2/XiVJ3MPqBidi+ntLKfE98vsqOdhYIHW9qf8mJyWTM2TIE3i2ufdXH2xwCfxY
K3wnMCGIehq4GWxaKv7Hj9Y1znURwR2j4x9Sg1+XyUo7jVp4g2T+OrMLoo9pnut5/1HzUNWvwyAK
pwMOdc07qaiGfe2vXoj71Ql6E6XWGfrYpMunm2OsLK7+nUvaJgHeUL/NMl1SzDzcDe7KB3HxRhsK
khdJJRjnUayb9lGYEs9FGrR6saFSlizGOgypfDbIq0uky/w2ITZcC4vmod3s8JM5UaALEfp2SleA
7Cla1g027ofTuy5VIzPEDprKHma1EvR9V8LYmfOXi9+4HfXGidInxjXERN/byP4w1UInSEPJ7qyO
dfp4zEAkYO7JD0A/fRJrl6wNbyfvjDMn35heXhYmNhHFaJKK5FFtG1mw7I912MwJ9LMJLYM1+sF7
iFNZQXVvcGctv10KszLKgw/XJek0wKy58rYnz/TBOEr4oTxrq7+FRO/v6vdMs8TRG03CKQucJZsI
a+dDWj01yUF1hmi0Z65H4OHn0KEjUoIIOWADrgJBM7FLMRl7zMaw3lTYHE94fZPEgYNEoD2MjzPY
3Yg4gUiP53UfJi77q1AowSwccb4X56sRhEWM2+YyS615I8QVPhD+0k5gF+hiq76FxqO3BD3XgKw/
JKZvkEKPrFpnTHVboBGNGX3lApNB08Lc0Kvt0WMxFXDLeDTWJaGwR3c+6JG2lC/Jt50eVRZH2Fhm
GWhbZJdHcqrhyAQH9CA5Yf+aCDbD9e7Rgu6e2oGU0m4BQA3bkMW7XHytEL3W5lUq/uqotFr/BdSF
sViq0ZB+xJSbv5qmjZss1vgugRBPDBYsi6wiHzZf99b9bitXZEeyY002mlV+leK7MBCyGY8QGYnD
i30j/zk4/rpH87rygdR3qO0ILqPwVcnZOTYsFQlbd9DycsYU14rBTg8Q7gssb4ACQ7x5kJLfZSiH
RjvvQ1n9T65zGEXvIPE7W9aXkYAj6yTyog5FN1lB8VcuCOX55+5zE3Lw9AvfdFBYNe0Pqza1YxtX
iTcXMCEMpIZiudhtPnxZL/Rxb4metq4Kw/Fo3CWA6zeOyhiWuLtLwM8xfwHsJDqtRWREpAqDJ0iL
UoRBnyIgmVv2PVcZ6pawmjw/2SVAbsKP2yK19Tj1iQbDqV1DY4qhuQY5/sx6AsLZ+SchChEDUiB2
/8/UDYJjvcup8bausoLlq4pvbvG3MQiNHN/YOFrOKflM0PDbMmcJTP8Xe+KQwwtgRWSqidxcc+HY
dZ1YSkNU3b4KlX0eMEBL3Fsu4MxTR9bE7mY4NRyCisoCdA7iD9sVH3vI8ocClVoladVUio/VMexl
EwAZE+IOx7CarttWo1c5ve8wEJHZwk8rTJMWEjP8tOXoaUVayG8Dx2L4U+mhL3L7orf6umhl+cnu
10anBbu+aVfRWFo5c1XmnT7s5rJJoMTEqrqJLUI1HBNHl7QBX7LXl/hgyK5S++xCa1FZ11jciAg7
pVUNLCOTZRLg0KthTzC0q9Oz0dAC4swjl5Ae3qUSqspncqb7Mz9tptEanFJNeA0huWBpU+gHnyIh
Adqxzzn2doJkGmbqoidg9SdvG6ULwyZz7pygv8YtqFRBP8DDcaU06cwHHV7As3DGHzV2pFPtyYse
fsjVUdeTsDpsFWo++KZioRR2H7Ge0+AkUzzfLkgImIDZhfeIS1iTCyksLRFpCD2JzC+h1OBPjcDv
4al5Qn1yX/eg4GACov+bIi1ZD+VzglOl+uOfs5nlp6Vkp/8LLmeQCaj8ms+31QFmKcE+CFfzmwC5
j8KEeOYby9a5hGhwrMXbjjmiztCLiz+Hq0mSD7Y8Dgk35qw2/evzzAC+2airCatNyTZ6b8OMlPmw
gvGG/q3sjRUcjstrllmGz9ciF4vWueQuLZuhYdZFejkrz2MRHvzSPpxTjdE5HHz6RiLU7nSS9GDl
xIKbb+XoryDrzYXpHNTKHm2YJ2JZ/JE0kmW97zRnZ0136B669/SzzFZmTZDC4X2ps/jjX0gr6TY0
UFi/Hb7MZsM9fQpwJ0UXF1EcY06VDBsE4l6PAP+aMorPxHM+wn5FB/OU3dSbpw0y1o1Osv1eRZUp
uMEgjQPTCtWAXg5Dfw3dYMcqMqM1YxpokVwGd8lgcbQ0PnbtUkg2sz425lnvf9vY/MT6Kenj8vvz
tvILB3tI9f7IsAXR//OsXpnqcZmhbYObUgwSLLYH6tXuPW4U+ogmx+m6P8fpbNjMk4OcO1KeUyjH
yMayDwDJLZfc/ud6aXHEis7a1gbYLhDO0rlpOCITxfMeWASqEbgGqLuLZE2IQebgHJNVvp6WAiSu
X1/WaAllQCR6koY4Trmfvs1efp3vKhgJPQw1HUB9sC64vv0o8MecSQU4DhmyBSaYyPRBQQazWiUM
Bl3tkXObSTcdK37AwOwsMo/giZqSIB+Vq8yk4frc7xLDjW0otVvfiHbumPlUt9TR1TqkozSAxUSG
PZw/vm0JRZJO31CH4JCFoUxr9+fmckxhdpURNpvKfvY1DRYMYFvLLmWscAskL319oSKei2e9YRtS
QUY8F1RETnOE5rzq6gxD/lndHqvCPW3owwxkla2q0i0Lxnp4LT/FRkoelaMQ3aXto1tJWe89oPgn
1lTG+UAm9xEjwIpBf3oSBSUQ8XIgBPjk52EInGQiHfKi+v3TCrRhASdIjbSro6/j8XOzvTymh5CM
f5IA13BBLhj/G8mzgOmOpXT5HXyW1cLc/eSt0T+clvHnt6fhR+JylCGXMUkKmbkzGAL0rR8QnGfQ
ZaN5KGZuipPaFJXGY/kdRcF5T0u1ZK61P29Qw49d5dxL+TF0Pa0FO3ibTMmheSP5WvNk2nQoFBbN
W3uc1NAL+/Vu1Uh1ysmwKRoztPjcFHXw9ltZvhDXW7igSy/zPDfzuvXYgWDmm3hu+A6N7o03q+cf
ZhanmwIn6b33tg6R4dXkNzObOZN3yvaqyH/roEZ6v+iuNFr4f4Dh8je/HQHqDTlNgM7ZElzRZnLo
AOD6carv5wl2MTwWXkenqvfHCPRCUi2v3K1sU6UHRKQGZ9iWbgr5EVDd+MD2y+VimEKToYMvm8xd
RPCb85ndfO9iY7/eHIr3AmyilBXH0Btj5Us+f9t4a8hElZLpPPg0KoUdruHQ0Rqt6B/B4KyI6wRE
gb6EAjg4hJHCf5HB5R+YRrpx4Y2vK3sdLdLuA9t+1FrHE67ODHQD83rjLdqJcKCQJUR2ZXJKoYD2
a9WCk9b6nGFwXiqR4VOxtYNMqxzrhilRGbzUL7XSUGrvwT17H35BkVtWZj+3tp2xxTOIv3xEfOJd
hW/2IA7RmWKOy4MncGFSh5naF91B/kNp5ikvyf03euPVZppK68iwRHjdH1bdYim4g1nZAGQs7Vlm
dAvpDQhfmZ9t5p45GLR1uf3EBLbqoznSfM6PKIQwUG8zzAOfxG1n3bKorOIG0KOdYWv0koyshUbF
zVk/JC2Et4qu6+lUp3MQSf+Kfz5hkxQrC8HvbJp/mrIPmzauNlULrZyos7ew0EZujEcThIc1PMvD
j3RF9dk28Hjhjn5N03YmZY9AlTMTPFZuilQmFR7v+VoA+m5GYxwKadEzn4ich+mtEqIOiRKqIe/6
A8dAkgrIVnML1+X9GeV6yhSNi00nQVkzRZPQjrkFTstSnFeEyG2+BYKMsSY/bi4BKXwMR5hqgOgI
5BT1pOW9nkm2E4jXz5GP/+7lYPwY/e2Bv/AUjJOQ2VZaC89WZRsuou/HNF6pXJk3rSpsPxNE3Xwq
RtimRHfjgPWZqaWr4PaI6b1BGUQ/stcwrKeDdwsoGgMUzBibUm+8twH/a/N2cmWLtnoV5ZK2nZaF
0+nhzqSCYH/cegBT8Oxy5OjxjOIa3gPW1K3jFXk3xejGpVvnpkssMiSB2ZrGVPQtRxeQkIqLHJFj
2W+7VNJKU2pnmuL20kpyPJHwUQiMSrnizjJd/HP299+Gnxn/gYrr6982bdfPndzqPEDdSwel9KFw
EldK1eARGbSRBjpfBCE6fzOpur3xcrqVq/tzji2buYUjN/lF7e7z7y7SK4RuqNoumWfL4EbcatgR
iua+MjFejKniRHchYmIZi/7SLTL6oA4OvnnceDQ/pVsedM09c8S8WqsdgIlC4cG3EF+phIrcZMzF
DPpBzSWHLNB6YO7qXzuhV62FPiwh9lbhUcUmzg9wVnJVE2FNQ1fYuAu5u696oaGRUtU0ahPOhHEt
zK3fM+1oJFdBNnrekoFGPsOSy/y1RQIKtLrKadQ4MZ0uyI8LamOw4OTKd8mLvzXjtNMoir3FRexS
j0Wl/acoMNTaibgxuRsEpTs1aBO326bjDJBH2pdiOsNPwCs3up2Eo4OMHuDVhAexmrpAiIRNUMI2
l71ziKn7M1WAMlr9QuA/i4tIyqSjNC0/T9AjudsYph22jCx635feNRdJ96WQMpEvx2keoenN+fL7
UD9C5CcMw8reRobaLAd0lg0ert3U+vYOODrXGGIdbPdwMm1y3dzwYgO/CViAH71el39YyR+qZqF3
iE/ZmUqAqFGSMIftRqSloLuWboK1E856SORVObhuFsp+4mlmt5kyTh04jXNtmlPJnhv8nrb0oKLM
Nf9f8gTsrpzFfs2mVTqYLbR2w8hBMHjj9OTBp2ZQm7F7UVKI1XBc+lcHQzZb5T5YXiytajn5xrEU
sWv72vsfY/vKdsZDNEQGzo0jnWbH/tnqOPIzUqSbQKSbiQCNc2rB4Lh0CQKh65b2J9p9B1zgX+y9
9Ll10rlAdmXEakHJwyV3UzJjVVpwjZkIgP8C5SAEz4gbCBiSOMyOUVVFc/S8tKFO4IHqrfcaGaij
a13ajwZe+AvLZzrjXGYIPEWioUflSdmC+YdOeHCE2qtLls6WZhlVg92P9d3Ml9VP2LzRiTeD87NV
qd0tewA1Xwt0Bp/XsIqgO89uDDec94z0xg59gFe/6Y8/BBQ9UTllfI5kqXpG7mxP2fqO0xcxhS6t
5d0gIWLWekBpqXLn7oNiFJ9CLIdcEYXZ/D5H/keW1ytRItR2h7VNm/PZts2jaWfCK6WkUs3NkHxI
n4RIeO2VOoYoAF7VGJ2bGzZapUI/YLk2REG55KKG6R4pbzfz1VvySdUBldHrXwzfUajolk+ijmmT
LO1HjBFxuEpAyLq25WaRvX/dIauuvFrnsXZ6+qMyFCy6S/V4p2AnHAKHPy7E7Y8xM/L1aZj0Yzyn
Qz75K8m7ZRMTSNRnkd8g6sdI6W43/iLV37OTXiBWGpHn9XvfEIZ/wGq2IJTG2kIw26IhkQLJZ8Qr
8AJsLCmOyPifbsA5o3+mo+7XPs471tztjTMC1bq2sG40SdpJzF8AfQNQSaQOI8vCBMEJjJKBR2Bk
DFImLMXMM0TKMzzYrVj0Tvg/Y0mYmgwtDhMbGj0QgJalhIWWKbd6x9aj1SZTJiI/XLLQh/k6R0xo
csHTosm4r6PQoKS9SQa1UnpkMNpVcb3rPxFfgktMTzqzUt9zOGTD89kko5Gk4G72hWX1tX/dPEXE
N/ZbEBc+yaXCiB/ybvcQZGpcuIOE0pS/8waZQGN+foyLGhWs+89AHig5Ok2zGgq+ScRwfmxju/qh
ImaL0IOCjYP3jtZOUUfe50rhrXYM8BzyJ/MImx0QNHGtS5X37KF9mPDfIRsnpBvVKDSYgahRgV7Q
tk+esuytnPNZn/3jaDlrHtTFUTmJRbeh2q2abSAx2DnmhOuS7toaOgcdNmNaMhlhgWCFepfro+rp
RviAHiHRDE04LpN8WGm5ithWC8oR78x1LV4kMttpdtooBUgCZyutSvCAB3DZ36Vja0hV1owHVw9n
MZRcMQyIRnYFUK7V/C/hPNs9yhCFVf8nPoaxb3TkVFulM93qCgp2C0/y1OUwPM7Cwy533n4zUAls
z2TQ8EWuf3kufGZdpxAXd4ZhI3NsLzPVWw5AusigPDo4xR3/zEeFQD4aNb1gEFHxrUKGce55LUI8
Wp/CB/MgTSJ1GncapX+FGMnt/4hWsZ+J7tyhpaM5iv1e53HImk7lIv/qm+3FNtlI2lTQtkHsGIE9
fgbNpp1bk9p9epd3uf++rsLZmidqtE3zg7Xk022Isj3Yj07cKwWhaPWLNOOBLgK/+DatosDWHpwx
aKH0wNW7ce4Z1bu4ZGyPYdVC4q/bny3BSVwIMf0e1VFvCMSUcep9Xv20jGfRfaxOa1BcCjRoz71v
7EV0K+WsffvurU0S3CPIhOYMLL9NduOVOOP3DqVrGz4CDk32QEj6L/2AMIod46uIE7om9nPnNK2F
pRvbEyk7HG9TlBw4vEGB9nl89fAK3G1BB++o8bama51eOTACWkQtSZ8gJXFu7y8jINRffi8LVtJ4
oDSSKVOPfRPxCytWbSutGMlPgPI2VelFWifur1jW3W+g5ARpFbWt/xw4Gam9fd4/CSOOwQfcMm79
kVKERbiKa2bg4VyGapNRTtsHHblpRP8PnpRCMRk6g7noUPyIKJlBpVQxXq1a0RAzKmPtj5LsV+RN
kVsdY2T7jjMS5dd4tjr/avTimsiRgT7GizrSdlp8f5NCx1cl5ds/zYeQRdsG4d8uggf9wkFCkg54
fEL/H2hoqf78Zzfu2iKk06O/A2cLx9XYlFWzST8JR0PIlwdqzawiXW+iO+ja3Qr4S6QtEcYJaFgK
b3KoB5b9nP669+omGPMm6ClB1SBSYALt7iL4OYx5WDEDqKe1JK/1dcVxVhWMigbDHq650q+/zeKq
HwSf6fZ0dn8+hM4PHBQv8/pq1g+6nMMV4EbeTwTQRIt3K2OYBOS9SZCPot3UK77E2Q4S31Wp9Rzz
wTNPVYPIxazaKow+Q4UmASoai9aQYZoWNmbcfXH2+bWLIkA8HUykzpNieZGnFU0lC7aocToof3om
+UiqQQQeUFvXErx+K/VAZClkZQQor1e/r1rl9zif/iskQ1dJy3bJNIztzwNyjdaViILyXrazECu4
kyfpveL9H0h0yIP0uWBqcbGflly5GXWBZBZLLSlbJV3T7jx9mdhQHY+aP1Ep4G4/EmZeCkj6v37F
95/MiOG0xJl+G7Sx6AkbKznYGzLpkC2PyqPm3w9fZMl11YqywtANKAyPkIWv/5ARaFExU6W3etkj
3gTBCq7j+AjAqqephNpPesZmI7gIPC61ckPV0J9k0KUhXZ30hL6UH53C1p9csayR63kVC4MAc+Lg
RRCEq0w/I6vfNAw0Y6FS5tUdwavnrRz64lZY6r+qoN9r895MJ4rn8SO2m/nh7BBSsoIbWb1S3WCp
cGhRdW8njXGiTcw3eJJ+YNZddwV6V1qlgDEoNqBESupJ86A3jvNjSBRuZPVZ7kv0zNs2XSKA1mm8
g5Dnv/Pdi76x9gCGv3COtQlzPKbVbmU0+z/+Z6X+R3l1Qhpva/JNQuQbq8iR2jknnv4NZu5JfIGw
Zq7CmKSNTIRBJ2ETMxG6KOXNfZPfzp7gxyAvE/i4LcCi5DE4TzWVO/61wVyyd93ffLbVlDn+UhLQ
OJAHS0Q9E58ugYMg2hrEtkq6bMJbtiP3Grx/vFVku9pQDmJGPXV6B76FTVozPOq3T/l7oPTpNAP+
sMPNOaF8hj9dwufrib0MGYIELqS1UfCMlRDCY3OoegVybDY4gSwNFEHmQm0GzhNaO0UshwRVkLsV
XAYMkVo6kXw7WD+3leaPC5qIZUjsbagVLG+nC37eugwwgkeNxeYnlswRL9vPFPKGiO58/NfJH2pr
JOcO2h4Op0Z7kFQ30s0ccPLUMGPUeQNfuvusPLWPCJqxQf1N4UAD4fphkTt5+jzarVmPC+XGLw8G
4RzSfwzZ15Lyjwgw0nkV0/dVHUm36IIh1yfVRG0AKjDM08zdVAQ8cn7tQu0FkUxqBZKYcadkd/gs
fw/Pcq9OqW0jQE5N35wzLtxMVetb61dY4lMGccjBXPrJ/ZaKFHmpVCFeouy0MPyi70z4SmZiq+JW
6KukNXYaqHWtmr7o9+kI3fA/HjslnS/N8SCiBGTG4uDWW+ugvlcdbR/z4bBPhkW0CkAQANsfQhHx
W4YjbQdXdi8xXkO2sX1GftK5AUgGuYxebid81SR7EP4h93cf8sR/VimOAoPY/tlhpPARSExDHT7Z
f5L5ytI0kfzh8PF31xDWeO70BS7ld4t2+WK6Cx6wCoKUyhxUEw9Q0A5vE8zr4HLJl8Ix/2knIeG3
MRIFPO7GNFn4STDLNGF/j5bCdJAHYQAe/onNhr/Mg1HE8f+2v+5J80KHRoojWLPxE6zSv+ezwCrd
rqcJpuoM/RdWCswdjeWKMDJf0qqZ3kLz8aVm/9tL5qf9T7sna1AYT7208tipvv1Fh1iDwQy3q/cO
7ay4IXBCjZaKoithVFix2LSDmDZFx0F5PVyuKmbDHuWf+OKhcvaYjN2KqndDWXHqwyHkfHe0X3va
NJp5El+2/WTLb7JBuzwcJVc5iRdOeeZe2ydWUHk+VXbifTyAtLDL+n20Uhlz2rfXKPJNPA3eJ82v
O/zwqkMcfH8XtblaE1OVfyNdMIrNSluK3dv5OY2tbpSsRdP6g5Cmp0Llb2LPTEHZjG71uVfCHOvi
j9a9nauiklWcMf6pDplvL8/+DD8ZN/ntRokqPbgzXk5q5KvHxjI/s9vGRhHdkQTsRrkZIL6lVmzv
6Y6P/BFJwrYqbRK4TBuGHBIdzjASPc9srTivxfKgnpbPXpmmartWwQ4MDrAveK86NddjHC3rBEhW
rIdQMDbVwODGLqSvwvWKo0dXl5DWxRMKcOfo6Q8JORQGdzeA9ACM9bIr2Sacw3/hzbFaZGiqEwRg
dAFLohJ4tFBM5qU5ChgDjjUXr+ScR5KC3XllzWLdKVnmsDLgprvp/zS0sp0pl9ilAm5opaXgvpzI
4PIW+qq8OBdIhphcNiMmaNenVUZrO+xV1wy64KLog1AiiYZUt4Pj7g/mZO121Ww4VijCSv4unSP/
NyMie08jT0D8wfdRY6A5lT4DYm37yisVJRht7ys6oNQpFfPuY2aGweiRh8ILHdyzlQGiQgSqfc/1
cbLlnIZNM7k/i21BeEBisUQmQH04OOLqXORPmSduAr0kumdpJkZbv9DFOWpNxNZLLYkeQfFHfyqM
YwRDXO5FyhIEzXg+T8OOAXwYBSOPiaGEi57aXOH/3eEhk9B/q/J+2nkFsNZNBXmSxvt/kAS83aq+
9loll72hHTIPabnt/k8suqcw9KY+alfAnf7n3C0sc5nEyYHifSgHtVa+jgSEKEJX1nnU1lpPxu/G
5boV9YX8C8ZWjJG1fpRTiwy9xCVukkH/GaOLbejZR7hFIjt06sTdLHPTZD00sRj619NnJWR97bG/
uDly/lXJVo5FJuBa9didWWKzr+QSfLZt7hata32aWUd2qijPsXmOrZIV16SX4J13yCvuRun0i7SY
OvKdM8HICaJKqM9kthW7+pZzXm7HT3gS+HsuNEgJwtab//YosoM0H6SondCRv/54rpSC8t8NLmnp
LSCAzYviGp+SnCwFo0V3OXW6EZzhwcJB3fa9g/mrjdtJ5naatYaFXBswwc3IWthy2BrbLUQ43IpQ
I8HboTaLdN+LvVn8lcyXwRxlnO3MHEn1oZgbzlPqaWhFMNiu+cu0I3B11hN9X7T3d7GqFEM2Fcsv
mcjt9KiCfFsxYtasu/M/shWBmMYu3XXe76fTZejlz8c0fPzH02k1pDcw/lGUZMFASE22kevanWD1
qnpOhuG4S9Yfrsi7a2eAPuDuaMGSAurfvEIEelamM33+hEWANXZ3VE2lqnKcQYX19nI6rRP4MLd8
GJ2O4aoyD7yHUHXL5cmcoa0b9BhHWn7+yuunYjZc2CFWYYh3Ga4OJsO2LM/SgDRhSIvYw/iQjFVa
kSO5jAH1BeDSWQdv8YWDJAt0hPR6G4PaJhPdvTRcuLNIt2n+3AXhxrqtYgksXENHD5GbzDWU+vfv
T/Wc5lM0LC+KPUg57beaa4bRyit7/VIUyZZATOT8UBgcuahNznXVpccGwsaq799luNenm0pd8o/s
7GS/gU9QOzt/+V9CgmvvtYqm9RQoWrf/U/GgAXvCKRxHuBP2gwBeC2qIhOWnoacyXq1YEs5mL2fp
TSAdN/aRbbS9BPvpsqx47jX+gfObGJguXmF6NdCt+5ahpcBXzRFmGOA7H6JyJ/n3OfEj7eXDstcF
IAX35tHRqAeFKJCD9NgbRROnf6raRi8jRShbijPe/X+XA69Agag9q/TkwZIThxK/SRqCrz7119vo
h+4XOtyEZu9ZzOMbNtEtIG10vvvlXD99B9QF50hlrekDeO7oijibhTGK2ZRFAMWzdX6YiXJ1JHrm
YJ9nuGZFTEkYJdwQ+L4RnWFtdDAgnIuia4paI+DwMKvCuLflT4xmeBAq7kaHTxiAuZmCnTm31P7k
mZNhbbLHVFaZv+KNvtAfEJntBkRbR22VMqr+RxTT6DC7exR8OZ8M6NVKhN+FcMxETk8szdQSteKQ
zVhgtwUbPhrZgXdIFtHgfsWRVKfHvcYQTK0n4ik9w2unnELV58hzM+aBPOF42gLORccphquuOJ3R
ASOEvrvesNUOGHNfKlDZt48d2D2vpvpcAkqgclI3vhlsjFyk+JNy6zNEWAyg3ulapPyXJv4TO8Ql
F2SOYmjDdO/V3LbVMqVOdrSfa7rn3N5wstIFbYO9/34EggfCKfoR9l5oILCR6eFysE59ZFZbuB+O
UV+PiT4eA0b5QzFjX5D2IwLmqwtMrXd/q8MoKcHXn7/zqdx4meTuQa3Iyw6CadWL2r7WpQSJMsPA
BK/vml53yXPuCbKZ7v3DVQRBVW8JgMQzheJ6TnwyT8148hD8afP29r5U1qcsfE0mQ6pUsYtNC0FT
fVKJJNbuliHuRL/tPGuplZ5qmHPd7F+aMJm6E0KvEYuWa72ElGeatSVSVr4BVMaUqR+37kvFcp2R
VskPUXoz1EEEalo8VgYJ9Xat/ds42X8MHLqY7jilq2NdwNlQZWxpuw3y1PKjTjyPpI1VOrAMdJhC
acaBKoF6a8WTJSHcPIX4QpVZV4MdbrRdMkfenXzVCDYGpvDrxG/0tCh0WTaJzyBnar2uivVOAhmh
aUocms+z+gOev6eAdLBy29/8l584ZdXOhkVzi0YYSmoz44S3ZhEVhy4BTqGgkKvgCHTGYPW0MDEp
aNTA+df529MeMNh8RIu5rlyn6L09C2MvJrzlXAs0gIZTXYWrLjswrKmDSqDiOizEzTKj/yi4LHn7
wFNLKxaNGaq31S2GRGUzoxIQvRAk7p7PLMiBkZoe4E9HvMaduEzVBcToz9xZ3y/Rz+KK0K4pl8D9
+swiWhOOlKlqA8spy21qOZTMKwroQ8z1+sStDYFS51KZR2xITFegakI59no46nwTMPt/R6doavll
lqcJMgHfmuObjIwdUuXSEiuODVlpTadJUfuL+W9c3PexE+hoNfDy0B/BimQW1GOF+nR5BXYSaxVD
gC8/Rs+ljdNa4sJulOp9IuoLySN6IAu/syhzbF+7cFg81vh84YfF+nW+PkOFzCoE94OsqG3H/759
hrQRuJTtVaHcaT8nPlCCeNYG3eAAv4tXuEgejYgthq3IEpyuOz0NWzb8QaJvKwdh2rFOEEo4PUtL
xKYkTQyEAMn/cfV7PlEi3aZ0MM0p7etya2g+w4tY39cRzWfT3BWeX1tEq6dZAJw6xrb/W+69GV+4
IJUJO5eviG5Z6Fi/0LCIXqKCG7kPaSBU948Drn4E0TbV+qZRcYBqM7E5otU6cOYAmd2/R0PwUEAe
7TXB0XHRXmn9JTlF4fCB3wHnyc9qGrXbmMqv8nsyIkBahMHwScpH3/lsNf5WsQYkT/laTk8lRHs9
+kPDugGKW9oJIbt8kOvMT7sWscQtMua3nLBkZ7SycFLuzk0Sg7uZTBjFOTx1tNo6cw3WIIoAZxly
0qMG2QvZWjA1s1WTz/EL7l0szCPB+NPVMEBqrLn25kkjLpFHMYny4GWos+JcS3d0kOByff+UYR4C
sowa7rjzde6x2N/Zc90nWp1TqT0rssPaAXwS7/gVEbyKKveE0Zd8IPlgb/b5ZEo3LyE4SwuvAyeL
dfpeNTSytrT29JXwhDjpprL2vWBOMw0M7o4WYSCwUNgHp59nd0jvvki9Z4h2CgFIr2/CjbqplpuV
X9ru/FBQJkU88dpwXu+PSOMMTGCQTpSXE5XQA9cgx8WSLclVsys5cuU9bNADl14ptWT8j2wE9o9u
G8OgJ2mBVIGrvmLLoabmjVWU9iS/VBU2gFFYlswIpCngYQr77i5BNPQzsChPDPJo7qejGmfFP+nh
S3M8zD8SxwkNmRFn1WEDa2DJeuBADVaVxT0DKxDr/HvksBsexVCqMuc7IYeoLwbiuZzZIAQsXmmx
QLlV8re2XfdNG/B8c5Iam2a5MNeQkFN/yDrLNfYfWQcl2simrozaL5Uc4d27PxQ7SP/hb7iNKUMS
RTg6HocMD6F0irW3m6i7ikhGovJq1vFc7exIzg0wI8UkCDLEBUbCzd9LN5VcrDjEz/PiVxfHFouE
rangLGewOwftFnTD3qL3Jfooy34ciIwvnJk1DrGQWjJDp3UvjdR9Bp8efmk0OeItZ0KEmWhNNlPA
VMaQq7lfVMiTD1SoYTjYAxv17XJaLhisqmhHKoO5RyvA8wsLt6tH09yDaDnO0cT/BrXHU5C/tXhF
lbHKQTSV2b2OPbm/+8zd2LMr7Y4DZG3iEMWUs33KWq3zBd+RpG+ptXMbM2Ho1/5sWQkEvskXM8w+
5AUEnwJWfoZrJL7aW1GOjhTu/qo8w8S/rrgsh54MtLDxCP6qJ5qU0FlPdngyJLuaYO8pR6d9mPoi
ZkbAhNXiGWFkTOPxJVT5A70WwItGaaR5C1c4P1GFK2rvLGHC8f5++nPrt9hCC6aIAkByL8fh+RG7
GH8R9VbYiDNwtFy1aNkW3BOjz3BnIsdN/pDDg49JrnQYrxL59iLxQYn0Ejja2u6Q/Y4LJfobF8Oz
cSpqjzrW85UkzHIOaPEj2ap5JpWWJOulBayj/Vd4RzxhMOSzcD9Yg4IyCZaWF5W8lVaSYsh/3tCv
hY2S4gs8si2UV+IugGL7vWOmEecOa99lHo0eOhuq20B05YVkIRtlFq1yWuhzf/VESOFZkSQ9K2mW
L0Z1K8COHit0bB9icx59nGIGLtP/RzbCi54dt+2ddqRaUDMODJM3aj7pLubm9uPv3WYvIO9IJ5v1
5xjtSdsHb4KJuTyBI9yPFr9Fjfk3rxQvvN0lfBrn48OXOZfG7D2NbQ3JQ9+lj9br0F8GoHFEWM85
TTBIPUIwPLv2A+GGFf5XUGiJ5k8iGx5ui4XyKAoIa53x3g6QmlnylplwBSESVveEpeZ2fD/V4BN8
OI7Fz3iLciMOG4sGvpfS/C+jWrvJ5P4zZNIzlokXWX/xFfqkfJvx4PJs4r3tfyw7mu83fdGzHgtQ
jBPm60XnwykRx3GOcAI/uXgKDX9h/I4ZZVVLU79A4Mg9m4LhU9XbGss6x+7V+ZJCZ2d/KBFfSmqJ
7e7jkXNpoCvkwu7vhg3gM/hGtKMcQshdMN+YPlVwishw1QYPrERvEP3clw3g97kJohki5qxrSKsh
MItvRVVDOztOtF68WQA56OVQvN+3katrPDygkEzEMMizYn/oQ8SXufPz/cqKVqYsS8gNsWfczPo3
D8YT6dmzxBPYB5N3+VgcgyXRd5DG4kPRyZrYPQWpoxv617xFn8SFMAbwM0dbZQznHUD3cdihMjtT
a7UBUk67sb1fdiyPV8eo6S7R+rI6c7rQ1/iK+aovRx7+GIL6lnmqxPkZ972W4ffCbN4/7e04h6Xw
1tIDQbhxQIckMce/rhoa+N1j4ghARNsW6FJshrt5lyDO+2E8oeGLJOBpbJ2vQ96migusZKkCrlgF
98n8SK8ijHkEuVbZEowaby5P6pz+8gR+RnMHdfW721OgBoDxCjRwVZTlk1lVYLW4tk0xpqpWES9y
afYFNq4ycB2eDLncLh6qd0CswHjb5EKskfPMFKzgQSSOc68px7wRLNsQfjjAFalYC/XDhhTaEVLZ
LHYzC/IgiwB1QZM1SqOKsyXUtOiMBlByyuANyhfu1Xs+DA5zQl5sEciP20ouedT+cdxl1HXB1VpG
RQB8PGDUIClHHquTw+KDooOa9A2NKB3/beW+TQgLAcQdvbaYnmFi4kApljRP2ZjRSw0oxf9HyfA1
3FOsAvJlEv69t3mxeibslJqcN5O1xF4YhkGal/xmL2qVnW8wSb08cSa+frvLbHRZmVfHuJJQDI6C
CzJRcDqWf0Z1SZbJgmMBZ1KsojvFUNjiaxqGBUZiPvb46214LdSCd4eJnA6XHAXKOv4Vx8MBfuIr
JcjsZUMjS313iuYXxO31MLtreZtbdztHt6TAM0d+KUHiQCuJtJZnNOpu92XHLS/RmlOOoQav2c0w
L0Zav9sMOF0qiLqYJQdFrCQtJIxQl0/XVaFUjWXDUL6XGzwcMh00njrrVWb4aAr1efrK5lSRAm+t
hMY70bc238DKFcN21r2lLvE5uP7Z1NddBwu04lJ5xWwWw3P0fErmksX9ZcURcAq79TltKdCigp3n
+8RFnv2Lerr103vO26/Iom0G5cKuwUZOi11EfvD9GQfln2m85WRWSr7q2zIRdjreAU0OE7nvUazQ
GHg+G+k6Zep+esLZ4gV4MZMDSHvs+5NksXhpF014YI2ptK/CDt93l4+IczJAFX37YDPB7uXSpXNP
ZmPvcFDWte4t9Xh5SFZYiWIPgiwtluq4VuqeYaVHf/7z+TeHxFDQHOO7y/91I2/Vo1DzvuJKFfM3
y9dQWXd0kmOCovfE9q7KV+FaPRJD7r6uxa4qRczny4IFho2F65TSvbyKS4N7nrgbze90h2/SgwrE
3sYs8nrR/tjfd1YnjeKeeQsjAFcVLw3JmwqeYanxJfenKRyJ5TDDoZDmoYRmqPr+FRecUl0XtMBB
V1cYvPmWUQWgsRj6FYbpYB4ApLBIELoMXPxVMryDxxjVxfwCOVfGy29NBS/PFjl0IOIVwSK5sXxc
8xgDeAprbDFhuFy00H+qLOgC06hGo6liPF8QzzdFc2WW89U86NlAohVJyMR2i2UitQQf1ilE5fcB
p/r4Y6xMCTHnqXNUKdyrFh3DQK3oFmqi3zTFuo8UIbmiwzja+HLdFoMi5aPE711DKjFck0Ahdcmo
kvvdDntlR2b9zLH/gGW/aeDFmKUsusv6GPOAWOBHc9Wj0+lsZvv5HGOfqfmznQoASrF8r1ToRkfD
EVpcv2fswe4t//Xwu9PIfyZU+Buy4lCvQsHxojbAp7bzULuq4ucYpto+JqKdMF4zbT6jTcVROCna
V2pzEbL9ECAHYQVyl8BgeREDwi6wYugESvGA+xwXHLXuR0X5D/jodH3r+eTcvEmSvw2njXnPQZEj
zSPL//8LP3HkiQED8FMrndwnlv96qYiz0PRPES5P0pHPJAF3DplFsYeNT7oM1kW0E4IjMc7hb+FO
JmVSJ7OIGPwQ2aMKB/Ys6w1gmM/GB/eqfD+GDgGcge4p9QcMRjvqoB8RMrRPf8ZAlL1nuO9emfNA
AYJmcxo4X6pyDVHt/WwQRvAJjRyHTueVxLjjyQ+2HX+HBlMvJh+mPq85gWVw0Mu0+SeKQlHja7Bd
XE5912q8JDd672hp3mDOdlJogzGLhRoVypjKHkn7qVAoSwWOmX38WHboUlp3Yr2d6ymnVKnd6o9O
hqFM94r3u/GF6tmWR46ikUkfNuGRtmVIKTz6uPGdSmkkUlTxL2CtKszfioRtvNRMVMl43YmmdYa3
V8IVPE79WsoA9CTtQNlyjNeItCmUkGtjtNsT4xKTyB73ycEsTNX9ase4eTM/BHIHhMpbWrXrdWQb
7OMOq1NCOfiJYo2a0QRR9FDfU5ioBMhUxP5g6xH/G85ChS1HwjKZcN6ZM6dGzPYBtPclcz3Q9reQ
wDgIWiLpAxdIOFjHH2YD1jlGF/wjIMQ8sA0OI7WVhNzDJt2qgT/I0CnRfi80yEYWR3xQCgfR6gjO
k9oPix5ic1B28xrPTDMWZAcWsNwGkNvqzr367GZyEEzh/l/QPq+I0aMTTFNf/AESj1r+glosjvuF
b8broG8UZqTg9ZU36VJppZlzO2tYr7gnKMOLLdCes5uOmh9TTtdqzJX8tDL7ZdL4Jq5I7cKn6rNA
fP5mNFBIm4go2HjWLGXTazoPNQ8H9M7joy5QzJKO3U0w8vi8b03RNytxDHx1a4/YHvnDg4fW/lbv
V7brxDIAGl4/nN5h3s2kLsp3H+mshv5pTUNHGUGGSLjLIKyo1AIBl668qJDkMziPg+qqPo6k8nRi
03acR2h3sikhz6w1HIU7gO4gjaZ4UE6YHBX+A0tG6Qxe3KdDZb4N4cP345gHYH/MuBRtAxHIrFL0
qb/A/aJA2apCvrV8jzyeteGGBXrKR3onm6BFRqOdyv7D7w0jiNx8yFBu6WM2PWQ3WYbnH8WSHXUZ
SqQ7wnHdsYRRERUazHMTA5Oe+f8+Mb2Y6clKxL2dxv5NS62lP0nlu46AQIOmgAvDlPIKARKf+FM1
8qtEn2BtwLAsSafmScTVkY25gLFy9Enmj8eSKwTY3bHJzOYEnP4qqjHSKhB/yfpHkrRYu9OYvzLM
48AmglSAsnFA4OJuHARF4LKi2jVX8cM/Awpvu8Vymh9fp/6EZGG1JcvqOYaAVFav4Rdlmof6KUVZ
+++k3OhMoE4IUWwGpX5KOdCEOV7HtpQKfD54ZidS6eBjcUJ6DHg+LsTdoAIaXIc7j7QwaUDJ7qB0
xwHBxy0HVqxWPMS1KP3AsRcx9nL1p5zzaEa7LrqHFgcB8tdB59I8Ir9SscYJQi+RbK/dtxTG2oVu
zLIcTXFUdLVn+h1LUdrGP8j8bFnJ7x40X2yXgBt7xWrp/N2K5m0R4Hymu/Hr/ELUglRNxKtam2gK
ngEDCmV9nV+fCrurU/A3XkSosoxLzPR/NQ4J/E1pq0BpIBVem0/nMd0RIbHXHEdFjHX4d0Pc8oN8
yiJZjJGTBYJU1vrgNvXxOv9WZ4M7xgxfQtOTGWLntvAG9cIHuJn35L44TxuX+TVE/0mt1HiEMBrn
zU8v/5tgGYn7Bz/9LfH6JJATy+esEVEvsuUsE7u2QIqkTbc9+v+NMhU6rvuRHls5/fEpBQ53EvJF
niFmRsReYLDawVCz8sePBrgxhmMuB0Tf46CSRNRyNpcjctliizur7/aXv2EDcEN4hqrFWy/RnAYS
PxWGvqjPyajnTv5+JWnGtM5AdJV1kPXRFT+3sovnai/Eih4bx5ZTFfOpVvxV0y6Wnl8RxznP9Pq5
+FQgLl0knL/Muzmv064nNAFHnInhZC+ahMMpbnkZwUSf1CWPcCQ/uf21nMsptJjphx4JWx2LdZQT
/5HLfBfpuzhtbzQpWcjeM9OZn0rVpGCxVPP9s4KtvvlgQfw2dgomOLLD22tLckDFdkPT3fOWIVyy
Cd/pOU/PDsKJxxP2afFy3vYUr75BNjXBF/H3SoqnRDd+JkqAD2ELQf0Kc7AyTLQQUgsl62oL5Nnd
/WByMRMIq0L72cpGSJTo6GzZpTEHE5lprFslUT+CSWzT5tRFhYVB3905qRI5wxXXG0AaLMJV+oVf
q+KIUdUwCBB74HITwDuI+5n1qcJSmxTgFFyUQ5AB1JTZkdijsi1pryoiSUQ4iYTe9nyLgNOC/U7c
V43fuhQFSo3caVfaf4zemQI/5WRaXlYqzbJNxe8MZA150+Dve0+Jj0pRgZMv7HAvWDbgmKBH0aJg
bcdfX90W9NqOvAJj1KF1Fq7koXgHtyrZmWGp9NXcIZ5Rr/v07yPHPJuKRi2/0gH7V9xjviG0ZKXV
CVjcfBPMT4mT2I+yeZ6124KF4l8yjp8mJv8uOyfx7Tq1RN1TlIEcBwLcXTiPeVYEGgGLfsUNophZ
VaGwzRwJIJzpzteVu1GADDF/vQUX3RaC12hSusSu7HT4qQ26K2Qdy++JXddjNmMsMv7gxR/hUe7J
SVl7+IZcM3lIjsj2+VAIOXbez7o8YPuWlT+NHPAiZ7sI36MpyYl/VNIbPuxqaUb/YUDmGZU/y5sb
xnwGL+/aHkxYqAfuVfYfnDbN2zupoMqMk378C/4X6yi+Jpxp2CHHe8P/I8BsHMrlN5EkwcAlzrZz
OLpgqT9MqHYQ6qJPyTPRlbLiAIsFrNyDrBInqJAO6pbJRHZ9J/0wkyKweHHNuRE1WWb+OPXkEA1v
kyaL7r9wR2FLZSN25AxbV6zhpxkkQDNVxW9Bln6FmKjAKyrSFk1oVJia2DjRT43qUmQQzFJyxojm
Gps+4zxQorRhLJMgZJmnI4MAlRVRUjM355o3bzFJV6Nra4qRVn0Yt7b23bZeIZ2yEdO462GfP1j9
tuaQqYY/3Z/SAf+ePcCr3uylCzrQtVVqgrczifOKDX2sbYD8W1sRBvonxE5ES4gDooRM4Zne/ovO
7dIMUxSNiqJM6dnH23OklZBvUE4MoyLCEzNB5w0p19Wzg9jRfOGVhYac2c1/voPwzHjTxA0k+BjV
AI0r57JCc4ZZDS6lDMddrFUMBQKIH6taEy7/LkEiadcNiaFNoxH1SBFl+cqz9V0y8mG+VPLIQalu
DLyD1h0CGUMgK36H/WuaP7cL+anUvLLaz4Dc7GaosYIgqcFw0rdvSk8G9WLIYMf1vsjp9dD2Awzp
GBsuNhNmuy/fCwQbG8Tj9eEaCkuhzHr3niCVJu3aJQ2CamLXOCjG/QcngbdLhjyqgCKn8IFL5awO
H/Gmbk+NblmQfQmA96MFfuDglmHjp9uq28QLVsNGVQTpgJqmV+R0ci5Kn1Lhdwv5+h8/D55wywZu
5ZoQCN0cA4Hiu/Hhos6iRoRwAEtpZRrbYfq7GvC8T39syuXj2HW1w1S051YU11hcTPuhBme7ftsl
vgs91zwoKLr3D0XnXnKy3wla0xzrOKw29wLSnao29CQ16eypGlKx3ncbl5rGzTIemd8bPmpd3PWP
tz53YcQKZrp1L9hPgL4G1J2fhbVRPpVBq/hVVQxXK28lShQFN5pXuPIp7EWHUjTA+OwBwsNXz+Cl
GpuDROxDJGdsCYf3boWUlOUmQuCIxswDc/D7X6JBIzlGY5tB9xsYvzmvU9aMV91Q0UxbsbX6WnQB
bZobaIKdlm2HYEQ+6LL3fo9THTowQOBczewjVIxDeECDFRPtSq38YTYILG6grz0vg4t7ydA/MiRC
TP9fUhRx3bSosHmTO+JLtYphmAYSCo9I+nK/ysB0qZM0wOyg2hVp2sEg4ODcAtbFgu11jrJf2b4o
EpJC9IZRFx7J5M4FKq4TklS2i/R3RfxJdRdYXC1Muc6VtFsSBpEA0DtmbWNyHG2I64qF7h35zdPY
hSakGDTopUF9j3QKNXpu2QfGI4k0uGJKd7f8HlX81JW9/bFwfzdU8DXFP/ytz5AeuN2xXaqXhjBI
1mpjZjEzuxWRLY0D6gEhRxaGQ8uHsgSgQOX+ZCbr+4CWbo8tyfZuvHvH17dBI1YusWJtB7T+M8r0
6dwT1yWgSvcmLb2e0qLK5GLPxUoa7vmuVKN/8RgZKFI/0wZ70oA4XwbVsRyn5XjmjyDCzLBnLQEu
mcnHMlSojZgvU3I7kPma2mZBALn87vjjgSM9zSwY6X/rvnGEaEOZekYTcIVEG/+XaMfS1PPSvSKs
c99PD55gBPsrOJZEZiGkyoc0mMOzUgM14sUL6HzZ0DiZct9VqdtNZVkpzBcT6pgIiqrEpgKiU8EF
FGn7sZn92bwIEnHPZqZaC7gJfP2wxWeo6cqfL2ADstY8ZbYlJp9n9u9HCPhfa1Tml4tSy2GVYtqP
V1WYep673C+kTPjKk7Pfm7unluezkuTw3TcR+IDZUi1a2/jtfukccTBt0mfyDGwsSJyIxfx+sPAH
i8abG2/d817xqqgL891vawTWWA8L09V3leoAexIbTLbEJYGMEr5oTvWGWEOc/+1E1pdJQLm7HZv2
RvCKF37IVMkQtBwN7UEKJlz3Rp/WsEOf8r04q6A300Yj669fH1p1HL+qZxQ1Ngus8Hk+JNOq8dE8
H/T5qbo9C2EXbj5YcyKKc3ylDlJjVonKrRLFQCCHbu4ObzfPOLlbCroqTbmsUmYyftvK0DQPWj1O
0haB9s3vNf8bwGjafnIEFR+lHFtZsnaPsb3+8UHUq0B8JGfynlIXdyvsUhUmcFjlUZEQ1lUuJaeG
gHm4t8xP3jjDhNUFcj9lb5SB4VivAyZS8nXke6LwV0VwpYLDOv4C2j6GnykBYQoV+5s7VLLxBECG
frBy/Zg4YN2RO0wmdgzmWVgswAbKA7DHeoCBpCwCbEkp1xl61tcWiNBo0o336AQsz+QAxnplilwD
cD4l/WNNJxJsJ9a0nC4sDARbz4PKmcbHEcit0TB7f6vloCC9RnZtPh/yEHdwncDP8iDdwaMmvr8D
AVUWjjz8XymnpqbkiPcA5ACBO4/RkeXWc2Om1L0cvmxoDygU2ISLwdVIGOq68AIxEQI9DmQ31jcQ
7bK//HtReK8xpgLaxcaUty8ewlzpjCWV35KKOypga0dAiIFxMzcfXb7LaHHlZXrLdZPCoStc/AoO
ILnnMndnWYCCIq/LgIQioxgT3nLBJtgtMFkBuyJiTEzRGolg2DjVAFzc1A28n9wF2QK/dp4nNbWQ
/kKk6UZzr5r3GCEF4Osmfb7znRNSPjoWz2ZimNYAHdvq4FljgNBc1pdsTGgd8EqwFJx6t5XuI7oA
6Ntj9GSbUg0ZnBZJB3IY4ar/p3bw9eaIhWxznbMew8zQ76qyqYSaZGrdbj61OOEvPh71bisdqPFb
rSTb02DddItDnMCTxqCpQg7+NxAnoVEUqpaL9KjWYPYtUZvVc4pPNMv4zpjox0UnY60oaYQltFrq
4QTv7z1wByZXLcshauk+UGNJwOrr7hNsTDQvTqjTJRM+eE4NSk8Z16bW6bxEjJHKI6A90PiKa+NU
cDrxbZYh+MJLjV35VyZjIcLfwAfQ0Ltt9ryAy5UROFTb3f02rYSVpDvSQmPLyyu55Y3A2ujtSP+C
nQ37LhnGKI1I+8ABUHQiiWojsi1spe2Hp9zSpIzg+RT5T0YwnmPT/24XRydM3EP7vl7i1TJXcc++
uFCwaF7GDoaaFrmwnxpQvqUC3nIiSBS3cq6d934ZUA6Vl+F1ORf01F7xh3rCEim/xq1pZXmhjVJW
F2FGzvcfKioc1M/RiI3dFjbLL9cEu2mQiXhq4rt0i9wDgNouW26irHKTOLssOAw+YQa68lVw9ypm
QOV0OstJjv7vSUUfOi61AD4l7TYkCjaB2c9QI09T70Wrh+J8ZfsV3pKRxAEPlI+c4U2cxWjaRidF
qvmtCAGF7iBSpTSrQqCNQYb+0/EMCdzGx0bJ4tYq9oI50Dc17t88hUREU54IHRC7q+25GGSZKTvZ
cYGwvUl1kWlFJ5pIi9kSGnUNyHB2FIRsyOdkAHJeOJNFuvNaR3GwjS+XJyG1wY1JSla0ebchkQiA
wY/g3EdQnXhhDVUaayw/+5miNzCMRfq2D49w88AFhQhDnD2NF0pRT7UjQtV05uE/4GlXoo7B2Un8
+AZcqJCFVSrDx99qz7G0YUSQ0UBci1uvIWY8P5u6jcZb49tPvncjoQvg92s5Pi8E+2Qihr2uw1Td
KeT0ObctpH5Yi7+Uqv+DjeZ5y4HzEk+eHmWrFyoUs+ASSPkucjBaTxNTu+WoSlJJ7N+4z50BgFzh
DqMKXlWw4qfVxXIxU6w4uSI02DAIuca1CvSNE4OW5eGOw7XNeFGTBOoZSfXHAhlXEEx4FbekhwPx
obZzd0ImvDA69ofgH25W59BI8y+bN26zPRBcKb8d9SofYk4f5dyXAOHLq2cuYbUurLMfLkcZ5PQ/
WjW1jK2qZYjUdQvJIuzOjkFw79QTexzUT4Eod6PnyQGlVVztf8KBEMHDRi6iayaGNvDjjVPxQiB7
45m2J0t+O8yEJH5/s+vTXkbvYTG7eLPqse9UPvzs89BhXDRVeca0sUoepVC+0MhHJz4FGYLbnGke
IONqikaMKX4GV6gsAHT2Lu6XNL4tdYXpQ+K4mzjLx0t0HaXca7bfqFTjlVUeb6T7m8OmVtRR12gF
MfyPTwcSTOu5oU4iWyne55euv+VVIkhikAss6sbo6Cy6A0XGzsqEZhX15Fw7C+CpRWEbod3WkSzz
HpCJHMGikNGaoF7cI4CEA29GGl/42uFr0gBHQYVruvDv/PjnTKPOiDN+txtac+Y/jcmxY8FSSSzG
Gm5DyffAOCCoc/RcSpB5JmWapMqzVB6/UBsFgP87i3si4eFN++QabkRIMlc5Cs6MBPKFgYmMnGXR
a0L2yA9sLd+b2FHgfeagPokAUA5p2NM+OERvMJhWV+oco7Kh4OacDLuuyIoKcxB4hRX0PYeMu6ra
7fsu2JA+FLWm6sSStIqy2bdbAL7e6WHXWAq+eXDBolcAca+w2HBmhDwKkAY14KSaknLMfLWE30EY
vxHDywFybm1sUxFpkzOFFLX6nnjuj1S0dY/6MOS2WqlzgfE6QMrVwVAq9O+JkMLBEQObfrf8yIF1
VbMhtTolkQJRYx8tNwTGm0y4qOb9eSDagk9lAMk+z24GBtEYqYlmaRN7zf+N3n4w7IGYuR06ZzTp
amnMx6mPue/GAoXuAYv/W3LgXLwVFt2WZe9oCFHIRI+AONr66UtUXq7EE5bNZkROdXLcHdAmJj9j
26PVbgjZbIiCqjYINkJaNBfcX9En3RClTIp51RPdECmN2hE2wgv+No+Cdxl9eoArSMVwAlUF7svC
xJDRd8jtr8rRMa/4zwm38eElrsiyQl6VrZyUvhl8ThiSOS+aARRMom7+NuwELWeH59cqHpnKxm7/
u3WsUB5BoP5p+Qe6eZ00eoZOAR7xDX1z5wkP3Q8zRFtoMfxvv1k8/j2DyL/7qCZBb+AxUGPkv52l
HUr2C7V79lopz7cjBHP1voHnfQFLB6u4xSnwTnO2e1mxNxEBxX0QrP5kqDqzxE4Dbp3IPN55RtlB
oo6ZHX7WoTpqqywXJj591bR5a4IP8Kv8FGeQo1sgmjywAdlTYaRateZQtsNKEu+sL7LO9sJEv+0L
Ee86RLcQbuOAEJ0KZWbgLGcBWMOu4bXgBctBiP/fSDr//OhWt4R8booNNBG75PqRQCBZNtXntFT2
e/GE+nRBDbD7CX6uMXFznzyMzbELKM9MLk+ImvXMJ+JmfpLcpJgFn0cEUCyT6SRMbTvTH0lyfa5d
scWYGm0vQYYkhu7OufUlbLvN4ZQkaW5rPLKtd+K9b/l+iI71jUkmjlkOmEHzYVHnGsGe778KZ6ES
YjeXcQ4Vs/zQ3N/M7v7euXSuBGqPkAktad/sPqC6vTzJ0iu0m0JSRNzTLkhEWpTQFfTDsIPgtKch
zt1oEyQhBruipJVg0JYO7xrfZFcwwm1GbLMOR7b2y0CD7gcMZr7ugXtLdd4iseN+/UkbGsLOJ+gv
BDz6OpiIPXcP3nsg6YkPT30iFPZ3y3csKcUC50CzRBu4OZycfw8ILDHxCBZwv7i1AvgA3eyQAs8B
AUD5YD4I0ydK4aY7WKOuQR290zjz+d5xUUTB9gZyCLnogpQro59usyw2I4PYSRRW15APT3nduqsi
DqayD05UU7WKt0EzEiF4x/wvC1h8Vd16G2QH5q8oIjdmZV7gV8QTqpmWbv4LdlXXFYHNMYyuNXo5
kIz+FOyWQqyonBphYAw3QXVOZchwNIwHT0hXjI34rKiHtAE7gHkL7B/2mZHxWLs/18auZFp/ccrN
oJcvPVt3xt/S2dY7U3ciNoBs0y0n+F0rJ5VCYh8NTmFNcSxmfWZOEJ1HAg/S3GJuUWv2YHEZZtgL
7LGnvfFRxOXz/aAnIe+i5OZIMiOWevDmJL6GOSfGKZyb7Eq4AX4sOEgT3tgTQfu1+7rtyTQm9Yxw
OJWf1piDSMCzT5WQPjxfpKxxJas1oVDt3SMXm1FyalwDuiQsb5rIWUimSn9HZftvefdt/RRJ2tMJ
mlB7ODANHtExupXBWGijVXmcO83v+1+HvUSz6on9aArMVPIGccBdBQo+0M3GSDnN9dy33GffTXQ0
l1fkCqZcuc9XeC3ouvssPl1eIo6hOkFdiNj+IfswHv5AndXRiMmVTAU1Au/rA3Eh7gBVbbqvE/t0
XI/kSxv6qKaxNvbMQXDRU905ddbuoZdBDcJT4WwSzC4j292nsNyYPwsxvUBnRjtT5oWltt86wHFj
U+8tmRSWmzJ7GqRJmQ9eLcYtfVwQuZCLDA2IcEdXWbqQTqudSX2rfGzpA+qqY/zAtIEVlSQxN8Zm
VExALOqSzchbrb6kmfcyj1v8CbldoZjQ38QvIkXYMHBvSM5ailmiR0aeyxHpbGakuowSpVK7c5vg
r6F39SBKxDwPxe5MWNCdEzE6/P/IUuLqyNhXCS+EOapj/SJK+J6/VhxUOhOYWYfDqNobWk+XJIqg
YaTDyPZuvYyAZA+3N1kY0phEatxn7VS+Rg0gTCfJACjjxrE4NeGbyQ4WgYeQTsJVmVMoQUV2H5Ww
AazbF3t4G6H1W5qcQ4yWv/qckQzXmu3TAiornqZBBqkoQ7truD+wCac/2nCrP+Q7nFM5hfoHLNCz
RkAc2NrgNv3NPiY9+QhA2Nis7BqmtWRuPHYJQwsobA2azSkU/TPMblhgxBog8K1Hnxs1NV3Dx3CB
EtdPhG0wWAsiXPRmjUmf0ATZo7HCL/xoUsLWSul6WsK5vREDTsfczmz05H8gqOMTORZn+tWlpVYv
qzTfiLbNHOsyEvms6IoAByaqNSJ4WEse0rSOyvwzepeVfFA9OzpeloITdoYKNQVvUGiv+moagRiI
x+PI3qVgGlVhOj2QtVUz6e8oG5yRdR3f/+ZJXivN9vwmHaXuSNOUoFEefzWwYohTsNHOQq+q3rns
dBwUbnOJbHMOihXYYVj/GDbUKnuE57ze5ky8dUaPyMiABx3Exv3jgViqNRLr0lVun+hnxT4OmT6a
7fMaO2cuqIA3NEueJy12zp0QCYWQHKg/BfLeC8Hd8V4qx4cM92NRGAFbR25u+f62zoGMPy7ES1i5
Lhc59LrED/vUuxImkwizHa868ka0N18IIueWTGj9FqBW+wDqQzRRabHtPH49CPDIdO1xvRI+grMu
VpiYy2skZ5/ZtPRxKtW3vn1eho5o76JcOAaAUSbM7NyWQvBC2Cl/nm39+72sAvjOIH0pKYRAVSIJ
Taa0s/icGogaQoi0PvssmMQaRnB2aW0F9PRfgrbFBWT3zIHNdXnJZ6UEni8tbRnKRHgqBexTx1Sz
5lgB+t0LS/OT2amd/CXYT5K8ey/MP+2YCzO03AIs40HzlQlJw7zWw+aPIYDLMkMiYQn/Z0LexZbT
3I3FuRKbNwYwgZ/mmNJCplnTzhBr6OKz3Jmx0mB6V7jlwKVbdgGppN/Q98S/8eB4OljbCzCEMKMt
Jisy7fWryjuP4WVCvXnb2/D0oQjHboa9zmR9QOhGukIM34FERGEglbzrHJlvzLaVp/FHWI9dMSBt
Z+KdGqtFOD7X7a4C8Ar1yUb26twX2suPzzDaD2C0yrPjsu8OKh25IoIo61RO3ano0GtnoQks8UPp
6qnUTZEvYJf8h42cv3j7JnNkmq+e80Nm2Gi7kzyy63BKrHZA33YdbaXFGhgkquNAuwwFeHSBUPfm
TdHv9EG2q/zMpgUR0pLnseaTyodsa5v421xfp9RKp/Yc+9H1UD9mCOQkkC1NlDTT/ypV5QQQsFKV
3DjjOqX83JekpX89BJDHYrj0QjobDAkkfENzqFbUfln+Ze++Lwpf6mmrfPe3YhbCmOtwx2AcWrZf
sLtYXMNttcrc5M7exGXjTXj92oV+omlG5E9oyYipo0AknUw7wVwjKivQapBi1HmrbNtBkBph/omy
XQHeEGD3xhew6qw+SjDAtIaB/JsnnFhrmP6u0NVmMZqn9aBhE63d29Px5Q1eMHBgCgidQhT2T6Tz
sctSxadsfLNFZUuYalqqeahEDbm/7CUJzK4x6/N4LxdxV47XrTKhQpu3AY+l2PM9RlixA/Oehp5Z
4eSAQiYLJzoxwAyvAXVSsOHkaf8tbqsfII/AbQ3Njy4k0KLwP00fCTSd3t6/O7q8c7MKCy1PnUhO
/MyJ1S4FxIWCtfMVqCW/cvGD2XY92se7hHa1UkmFBhmsi+XUZcsOLlvI8CCF6PmnVZ1SwuqrLL4+
loeZbD7BHi46/vJIQacSKBtmAFOcG/MBSMyEO6XLBtIqTQQoEs6owSEcvqpfelPWImY9ml4ahOm4
L4s0YKet6htPT4hioda8KZWLxSt10lCw+5vsxbyWjzoYLXy1NDNqucmSOD45azhDJKN8Zlj4r+OC
iOxhArek7LgMp1LolM+wWIqN2OoheJWxdKbMfvD1Z2+vrBGffpH/EfpulpWAFqg2dg/gT/nngvec
MIeNZoQo7s5+wRyBRzlmZJSUKfk4d/ye6Frg+xN3cFqS0kRZS0wlF3vTLHcTaeVN4sGYlFX3x3cW
ynIQq8zKnsM3Lz8PKvcSHM5FnpXW4lPDKblp0IW8zhFLIFKIzH6LQitU79FyD7+DaW8lqzblR64b
S6GuFtWX0vMcGjR6zQ0S91x6mVpsB/L7zT+vGC39QwZsJyJsu05rb4SU6SRk3HvIYVa+T6L9LaFR
g2NPNwGZT/E+6vPEZrRt7p5BKZFtBiApTiChgaDstTUD/pbusmvgOfXQKsM5mBPK0LiONU6KCRm+
3PDEXeoGSTwsoh0m/2JlEqh6QxLYjD0aGlNMs74v6Qemeaj13oSyJHugNjIPfpT0rWSLwAxBv5GX
V8WYrgZZFfyjjdmbppfwG6CWn+uUnTULxfqIj9md3nP9DHAbqOqPy0AdpgNbQVZMVpx0wW6zFQXA
BL6nqthl/EscvHwRTQ3lXOttmhOercYGoaoYipISAobGfGfNGX6Ad/hgU6V56DaDmBOJkZN/2xGz
kA30JjAB4AOiHs722100IRSnZ4KUNBKkSAnUvdee1yydhBAiV460wLQK3hESf1z+TCh5Rf0fn5yq
IS1HPG1If1RHg+yUvHBN0OsfURpJJiLHaupUtdC9E9LixlVqfHVgWtmxmMB+PzYyUa/hJoKla9bH
nQL+L8AqPCw2qyJ2Mu42/lIfPh9IUSyqP4stI3cUwZRgRrjuw81r0W4lMQHUU7TE+sF1uG4TvLAQ
p7jXmDTIn9/2lyhhAe2ACDAuER0ANm8j8vO0FswhDbD/oRQ/OXsBu7rRoi/xKtoNlzYgQrhx2kbp
HhP3Ycc6611wUBKQHhY8W7Fxv3BNkVmEALfSHzrDy+QC69dXQERI6OaPEqIYLjsOo4Mll60PJ7wx
Ivw38NGe1Nt3A/N3lZMqf1OYwwu6mxoY7EM61bXXTKsTPxtxzveHx5Jw/PiA4QXtsORHctuvMubD
YTy2ZcaKDKzpjC5t4f6rQZXVXDSR0DVD3TAyipK8fgvsMcri2lnj1Y2TfobA0slSwGWgF4rd724Q
UibOUSPebzR7JeR/Pvkst2FPqAomXc3FMc27L4Eb8x5sg1PiFejI6A0rl+rjeQNDe0VXcRwlKB0f
omiWB+UQImv34pd0Q4P/XLggan33tXjKD8/8LuF61E29/0BJhfNoa/KvFZBbUW3tCs0GCBQZSpWp
aAeVqnjkYj33QRLRpXJmz9y75y25rss6JlolSaZsUKaHutEaHzmZIuxQJ8oeuZjVlkh8HhhW+XwU
shlNQkqJMFCiv7Oa3ETK8tueVT+OT/xNUEoXfh4JgL8BV40WH7q0aCJI8VxlLZEprGQjIvUmlQLv
3Mr2Hk0ln3LDnsSxWlVYHotXUDJKQfrzszHVmr19RRkdMRZFoFJ97xq9Ulo4SDgIxjukp1qxGKsB
wMZ+ZU6vH4xG3LVtGCPNyr3ZDWt7XLhGNOIwLdYUfMzyw7yMT0t3gNvyA61O/3pyKF5+yXmCKCGl
57hY63yV5ugYJTJhCejJrSpbvFXmYcK/hn87sm3nANxk4CuDRU5EtkiACki0RGBu+PU/wkJ6gdjC
Tdnszlem4/xHEyJdU0xrUoiHWeeLKyvge1MT/PtIch8sypzWxuAJz57z6WK0PYdyQl6lNbPSFUEx
z+LhYfEktO1xFfZcKLtMeXIz6Vo4Po2Lcol373Lfsc2OkZE+ZaqWOu68MrGI1JKuocD85CvRPVl7
hA023+aMVJshHzaLRCxJySw4vRDLEKv0kfcdXnOVyC7E2FwErNgmypSFxM/FdLPUfTpShNIlCUPg
6pyJQ38ThgONTnFc8aUY84cltMFp0jDHP8A2vNssWUa3jHdvLwCpCdj1I7QRt5XGFdupJfekSymF
lT1ev3n5tZUC5Xwjrtno33feVShiQ34k5GCI+MeRatrR8xC3mo9VHTX4yDbeVN9d44LODVWE5ZD0
/ygYhZDfAYORNVKMzxYLPISL41FEDNnj/VQBQpXvhI45ztwzbNaTrXXjHPQL8YXjlAxA0bOZ0fCS
XME8WuEoQlQ0jTAxo+Mss/XiC15cEcrTAVuUvV2v49EvjqQEzWvMy/QOQXEB15/RE1tUvhMHPN/q
7apuul1/lkgbAapDGISz0TzVKx5wDS8wqbwmn41vDM4/liAggMXB8h8jU3GGLEQc7pFSa+dpOH5x
765W5Wz03eJssZrrOaSluBZqAj9AUED0YQbvOWHAoUW3IBc6xGqshmyFRitLLdNpkjj/o9chYCya
RzluM3+B6d7JxJw2kGBZU/DWDIUAx8biBshRwoF8eI4TWc+63N8Uo/9vMoehOlnYYguzqAEGREfZ
/y8+lEu0FQBWRTG53qzSYjaoYu2K6okUYcr1V03RVELSWRUaURr9vP33A7K3+sjdZd11cPJIJ67s
IJ1CEoZVvFvoCTha4NHNUe+uFRRFXevA4IFboIHyC2tsr0hzT9a7A78qpe7vT+QLqcsxjSSHn8y9
umD+6LZM4wRP5kHe8xKhO83xXftyRVXSQ8xcGq/T1x3muV4f0GXXKmaz+u4R7ik4uo9P+yl5fQfq
qANLBg0GdfKkpO7wCb0yN1l/b5J1/2R/9p7/Ihdx/HTCvcyhyK1BK//PVR1/S3vCrOVlK1jGHnzG
W8hOr5/Tm0gUPQ3Jbtoy92PuUHoPYWW/egk9yL9ycWcUl1Dc5aJk+BOWjrpurK2VN/zWmcBpTIHP
94hu22fngex65oJ2owYaua40ei0ArOfjTiFgMLK6NXA3dypPtHGXKgUE6kaLBYqvjKOTAdrmzE+X
IvqT3SAVbut4ngAB01rKcV9bkw8Q9V9Nlyp0o4HINoMxYHVniLb+VCewI02j9jiuUwhHSh3+E+p1
4o6K1xUvqoJtv6eUc3dUGNMnnQtgG1awL6x8bNvUhJJsfjfUQvIl39P0XU8oMYl5+Pu8eO0l0uhG
TvvApwY40MRbyliZT4YuNJ/eQ62vhmpxmv0xGRLlUhSt8KzdCfbeOlTBmQ52SIWU6phKGrmjV0bQ
3wGtMUR6Zau12LWw83jkSh+6/9UqLyzz5KnHAxHKx+ZXu3Mx7zISCLDpMzOdfUL7j9878Dj5f2P8
1Xsopjy3EHdH2GAhV2p6jKhini8cGHZefeaNF/XD2y/c6c8cM3xaD/bKYwlgjNKUvFOtJIzInr5e
dVmbXQEXPs21Azd/rzeJRPFiZDpRyx5YIh+WcRMa2Ycem2eAHT7xTO1gsr2Ya0xGUjkKtVdUmlNU
IVTkxk2b+oCPMLDNU/yimcZ1ZgUPsJ9TkhI2Qd7f0wCiBpSAtE+Uua6i0TxqZ2K+GwePxQcrNMIJ
5QK7Jtseh2vuhUa5ouVC0meQHvQEFkypDUOmTI7iJ2lh47JHRgZCWb69UE2r9h01wH30mIqgQDD1
IqHogcTUUB1d37vzqr2MgM8MgWtRiW1rFNPYL2jSs0qs4FjzdWjMqKU34GttjCkWNYCpN/TMQUwf
oVQgO1G8t86DS6mNWSaGTS6VfPrjSv1mzmyv8yV4LJD6nSTEsuq4CFrNgrWNCAFgGc6O7H3xJ+4S
FBW18VvN3H4mjm2KIFsV4HR6G3TEmMnBFNa12TsxRFBhbmEjWjeCa1t8BUS2cPHTHTjs7IoVKeEU
C4B6Qt/n3N2fdEkSZV/65FW/RZt+xyXAfJV1C0FxDDgBDla1OUKFg/kYnyJf75lMbI/xp88ZdxMR
Vw7QS14GgGX759qP8TH7MG0HSFbnpEodJd6CGokGCCNT5ptI42QXxKvz1AqPoRgHffBFd0ohX4Ah
SonMj1t63X2t5xBuMX6zNzNV9EGAe1T2OX5nkr1RJXbSHovAMtcE3lqW9hOL2z/uZsnNYPGRjubA
N51iylwn2bR0Guz0t1tWnU0zUiLZeN7uJ0cEb3Kg/D1VgZZW4b5sJlK0PFJqXYfz3vZbhkWAb7Bz
nwUwalx56enr1o3cgz5tPxDJASyFvshG41BZC4KJioA5/6AXBZ9dFrcOiXuGlbcWmqywQph2gGoa
EIu86OVNblxb5c20+siaS2cR0DVsH9Z2EeYEnIu6DSjETmE3tWwb50dQlsFAtUya7fl0/6w3t8O4
FAzj8g63WN4MlAZwDwDNKWc0pQRKBaxDhdyvJmg5h8QBjT59efzzLpTonuTn0N99Kp2Oumgh6DdT
+nmKRlclWSLuNU71rba1WZ33WRKgZpG6vdWNeiY5zP2F/gj+kPWXuy4JH/gKn+evmslr1year9Bt
xW6BOevZpijqrh5u9uBWsFOd4GVBEQtJWXx36LQQgY0EW417Ul7H1dgXsdWhGTD7dYRDfaE4lbpu
BP42cdb/wEd9I2dYzxC40VeEh9eVVEzthUIFSP4o/xWphZb8VopUt1iwB+fjtr2YHEGVzcDIgk7r
FWy/a5+dzF7NdFFcF6HG9Eq2sx9vxDuTFTpy7nvzS54MdIsR91fdHAplskWGcOREJ7POA5RDWmzh
RoAedHG79xBvg/33hBOBc5AdbQeodHuIWK3Ca4tHBBB0737NAeZ6kUlN04Ljm6DFbXGE0r8Ghu6K
tHPpnH1KhGYUJ5WC7QDo32Obi5cSwzwRaIt5KMfHwUO5j4ahAzqlL05jICyhPO8WdFsUv3tFeJQp
OhXvRRsjySYf8swTPXIIb/S4V9HPC43o7PvB3YjclSJTjohbddE13D9rGLjnMyXszakz1oR/+IBR
b0luMO1Z1642Wk4veVgKFRDDDrTQKc1oj9GqzB7QxjxPyHbOu/dTw92nox4NKW99tIhRBPNNpL5d
VdK5oOyEng0WiI80bGVMYKZRCE7lYDecQB6qblr1uUiAmjqXf79ceuTLg3N2wKEzD28/mcQD6zs8
CBNwLTyjmy0/FMqSLzXYievIaTHXADJ0PWwK86ZR2It7HwC+ky4Djl01K5GXIXpyStLWkgkImMNj
tRRtQXm8Mj/phMtKTAZk6opTFN8IWgTY2MWXhSoPvGYy8Dpzee37is9Mhq7lTu/PgApbrm66DiSW
wsBlGTk0RA1O1aQHOhO4Bksf+257Q2PL/wgeaorEYIYHsVQbRNEY/GpG7GQTSFlJ/oMXq3hGNm7c
sJIRdWogTLNCyyJo/NZE9/4bMYZmgUBc9e24RHiqihLPvh5waIOl8Jau91loJj3YAawn5qehkhNl
dlUcnpqYEvWTRa6M3vKe1pmB4OCHVtGvxkAOlL6cUhhMAhiLi/gQa9QYN3MlWHhxZOiA66FKyhj2
TQ4iM+JWFu14SB0M/ixHy+aSNF1b+qPvl7aP0hn91bZ0dA1G7mQ3Gwt97juO8G7sx/HFIkiQog1T
+TILqsZ/oehEtu4uKiJaYw0WKJ77pQsDT2pS9lsVRMSMPcPCS0tnNbZtwCaforJ1B3Ss76lcOR1S
tJyFkhePoiQhMdsxQtCUBTY89ypieplB2TDOe9jxDND6V3li5UJFiF+KWv/jX/U5Utn2mS4jtPex
TG1F13hjEBG/NZn4eNn0LSI4rBmQUU8twalQoKl/PBvU1jT4LLH5LsgifoPcrt5M+mEjqKxOokmj
qXgLwiZxDUEExV3MoCH2stf3v8SoDadhB8aL85+0BNdDQkSa3rxPRMTB0sJcSaVJFBnvBqGw5hHt
wO5D08RylQMOnhQD/+eJl1tcAgUCZ0V+dOkFVGvB4MSiCX2LGwS18pnGALmNjcrd7SFez5cawBQk
CkDmflzcFa8WaqxZ1JAFzldCD3dJVRrNewqF5D+rkebAW3iCM3NPsYzNwL1kwDJxIvgbLxNTg8o4
Hx/j7ZQaSsuH+kp3uWVcrKTTAXEXGD69Tohqe0P4nr5cAFmrORje4lIQEcP30ute1bz24ONQkTXJ
ko8LNxMKDsvKQ49VpMFhEF87FMu32FmIbQt2pNTDJjzfidAcSwYdZHQxuL/f5jpXWVt+cJ2+otcj
uRhtOd8TK3GxRts24a5zYtSn0+N7hXqm9HBDqMmKVpX9nW9l7Fucc+n4Re2UD1G+3oEU6lYTENTQ
rSnneGwKN6mlkRO/rO+JfJlE7QD2w4ZzSCl+LuusqgpRRELpVHeU827J6r5Gco9JFfChTA8a/qsw
cP0vnmqZMiQ1oyV2xt6KKWes9wsRwKDCdYrYnhKNqO4E80FUw9uW0BPt8uoIY+Znt4VS4e4iyoSV
RR/7jZGbrXbWEkdQr0bO7SMXWSk6RbFAacAOaQRu1OupT+6kZt12q7Ishin2y8ecrNbsAuJomIm7
ECuMLTH7B0kn4z/laQVinR6W4UAnUOT9l4hTfHR4MGvcxY/4Zk/VTRgI0SIcbpfciIGwR/Pjjibg
W488aqS3C1RFz8M5xWGJ3aOC1oy2Vk+iN3pBcq45irL/wo6pL2WI6KlsKQi6/fKVLtz6+dSYqpkS
KKvHKj57Tdi9PU51NsmRUtZmFidfQ5rA01tTzOfGzS8peNP4pWiJ0sSEQkeCtJnbLYQf+e/UfYJ6
rlrKCbBT5ZnyULLYZXpD4inAAxTO4u/tp6URkBie+UKYnpsS/kwQimk5bSrWFATMcLA3SD+pVU2B
jQJbXmaGEcQV6XTVSIRZ1AUDHpDUC5HwYj5Q6XUaINhH4Q644jbcb5U9f8eYvPo5yaJ4lP2eIcwH
DVaN5E/WesbBo6nfFSdTdXQJkeC6z3dML0uAATR2xQvibnto2BrV5spO1o1IWrhjFbPWgGCKPcTV
hmDOlFg0vCJfvUxCSc92lxlwlD+uhZVGHMoao7Z1cXkIeIKZRqyB0ykBfPlxLO9qrieUcum0BYMr
K6GV9qdiZeyQ9n9mqeP2cdxuTeB40+mYkb62zY6kzTSSCWmH9S43MOzkHoH/I9Yp5ccNQOIQhGB+
BPVzLTOxImiaVju7+9j/iYvcYSRbw2XKjSmjDmF4o/vLGNRLHfQowGEhUZXuU3PjnTrHS8UF8L8p
CYf8TmW1ZI510btG85w/Mvoefasd77RCST2/8UJKsQOtwldcTXBoRi6n9zc1G4n2N/GJLRBFmEda
3N8Kbn2rmSNQ8vRhXBThtSdNxyDOb6swx4Hytk7VXVngyZJB049aD7Qk9p69urzFCv1clAVgOsy0
807bzmAYoqgLx2cIm6u+nXW9ZPnQUfYB2QnVlQ/mkc1EnKAl0/5tURmFDpRndCshsj6d1bybcil2
1Zfb7silFOuONQwpIinhEcgFvvMd1S3PJJvi7oRqpY/VTCQ8wx5t+mp0nvZFN5sFABP6mss3dDGB
08gqpY79juqi1nuA0eNaFKjYohEjiQCAFoNw7Epr1WCSUrgRr+cjDUzoI98cqHOx8pG3GUhzICjm
dipvCRDVYoRmW1TJb+SAwgqZYHjn/eUrkuf5PMdYWTmHFxK/TpLiHdhEfVW3jF3kybfYTGSAH3wA
uk63y/UWAmjJUgfL80jyA6fBBmPut1Z+1VWeSUO2mFVdP9TU+xDH+q8OxFHjnDcDPUgRrpxyF4Q/
OoLoXcM1rAOTK9bVC72QmoMqgFUJI64AQBEOm0l6vT1lAk9rb1YkHVQ8AuHYGmAe3GCzIZ2BU9mV
m0SUtrk0FruJC7XID/M93qsNDfaysxHazU+2dW749J2Hr2hgMzhyLAM/JLWbsLYyIdoxqYABcyeG
8aTlttaT1G06eVr7QWgPUcbiPBmsW2JtHE/7YsERKCjZZxz08UfQUGv1UHUQef7i5uCvj17Mzv5t
B0ZYlVoEz+h+LH8NKqsvlpbuuRX18Uq+hbiLfyPKxuen6C6Mh4bX78krnqe+Fba9kzBJ6w5p2ca0
CwepUY5tO0kj1yTVsWGDcsFK4TKfYHMwJodA6v+CYM7qMm8wvh4TRzODJKGYcxv4gtXVydzjCwAS
sTzcs5V8aEdutHGaV0Omc0NBtR/TEw4RQ7gTCU7KRiRhuk8uqkF/GLU2Dljndhmw6bLwCQwiaiU3
mDPfG1GVGgGJ+b56jcijWBa/29mQ5mQzK9oi9a1bCl5j3pzLaQEncZxS4EDOJ1XnikjfKuLhnS8b
aMLYeY1CT79mgAzyB/74gQrbJsGCKW+hdJkP0R3JSLxteKiu5PjXH3DWr8cXub+mrkpdwP16azAH
OWdMcElJOMg681DGSueHXI4xWkbWdfH2LOy5OYUZKdARKOwXswO83W0014JSoMsZ00HJWIC9RU58
3ocZv4dprUycBrCp6Oc3Dtvkayn7RoNDfUJCTJ2ST6ovXM0ZOCBtIVBr5A2hm/PgOknacNXQGcvN
TtZ3prm9PVlLGav1U3EpL4sxzjdvSfJ2AVoTp4D4xKCv5c3518FnvjsAPspXiGdDQ60MOYcgjfii
evLfOHLEjqeOQrhRFr6VZ3btQSGBbC1l1XQfaYC31nJVvG1D58QXF2sYTazDOqOHFxv3U98yjfIq
SSLjS3zVoOLQTORkVa7qUGMOmWrcli3efjir97I3yNlpmBHzx/RlnfcauNPJIUjAEiu2fJkn3DxP
0Vx2Wxi+pJKE13Kq4a7Vs5gyBqlOIY0b8zzaW1i1r/RHfYVHaLLcY0wvmWBnndFaomTkGniQSvcW
tr/kgfoEbDBswrfnL+yD5OjdIglZEqSxfv1ga2I0EajR5a8Mp1212sfuuKLwPMxnXdfxWLjkHKbg
OYLMZs4ra6L7u8igbB3rZrtr6Qmn0fRDYJ4im2FWHEADORR7kMLJUa884ZLk2IRyjnNc4oNwa5gO
6JCgAZDRp4b5ozbSAsIYHzh4vcKZeouqjSZ2B7sF1LaPPNdMk1HSplmwRp9urO6BzIZAMQVf9S01
JXznt8lf4KnEjYFBd9/Fk44vE0uxzGCtyE11C4YhxWawi0dlokK01gci0mlrLjTm3iz9ctmmnQFH
XdZHXRxrccEz/AIci8b6lotG42oSVh4q2XZjHrI4yrNZypeWLU+RjguiIuCSBP65MKOGzPEygucQ
2cxUYMX4rn+4iBG85wBXV6ABhMGNXyW1NlThlEtL62jfswXGaRahgn0iFdi0deqerNfM41v9198b
ScfZ6ZJnbpy0PIgGSRZ7KQvWDRCkt7B8dQKRRsB2PcGOEWhFqWTIwxoelUey/USedcY9Gz/WQsry
e2dJvd/Yiroz/VI5V5n5v3alDcpjqE1jFNilxuTK+ECuLxFwzZplNowR8cFC3U7l34nxXsBXcjVn
fLaSgT4wDx2bhSpJC0apAMGMtrMOSW8TjEqYRsQT6EHZpci8PIK/Pa8sqkwlNRngkyKSQ9Txw0OX
QNYvD0Yr6wU2PWlzbhuX/URyul+vPCy121IbJtGmg/IFeVjTZbL2/tbagTsC2xGa73PYJEJVh9MQ
9zPnrU5EPw/ABnQuZlIwS9lZxSrCRHCqF16Mp1MQzKgk5fuwDU92czTL4shzCp2F62E+LPGBBTnZ
QCm3S2sVj5X8rog20gpReu1wk/1sLFzXR3Mif/dNeBfl2On8GzHH8WiK80POTmqPttVMnbZ5QVol
E1lqB6nn2dR0oXIq8hJcKwy2a6vW+tjxLhGs/RVnYPB8SrjyQ9LBm2zacs6mOJK/dIZx84+Hiu1G
hiKLXuRbbxaLssNiXxstmAiikJrmGexVVe80ilFFa3orpHnryK56kzCmmCPP64WY3szFMWoFJJXI
y+fTtUXOwfzn0vLsxMPshoDHwMRWxcvBJDdahqWqfkv1cJ3EVpHjgzxmVDv9PbxPk5LXtw06jID6
3fhh3eeOfFvYJbzJMQOjrNFI7ndGYwAjVAJjATgHslF3B8R/9C3LY0UTDR3eH2Vj3SMxysBaxSOB
5mbQvec2VpxqEhXMLdrnaL4LZCf37behh1CWWkKYHUmC6jmoRBmEneyO0qL+EXTJ4MbfaAT6jpyv
jCF13Jq9GsuTAeuyQnUPAl5N72665ks4IziRFvZLMPkFQFhx+AKU7MWEuxh18L47CwgcjnhcJJMr
A/ueMKDgeyJMfauvHCsGSwpKzpsMvkl6QgyoXiDb4UypUZBiH6XraKYEIDC6+Lvv0ZG321NUCsbn
GnMAPaDFSfppIhsY1n+hMoos2WhqeO8WglMRNx8e63iKYLep5SteVepsefQ8ATpfesXVzWMPhQUj
FxqSSBNn0hyuK8EQuBURAc76BHbognN5VFXv0SGnEVJx22qi+MtR/qruf/yKQ1+xFf09bVUB/Pz+
Nchnj8bKwCRyHwrBtAXllwCzw2Af/UmPCjOSm7j6WmmXkUajiZHUnsVvLRMXxcUt4H8UyD6oKOvB
4TmkyWLFfO9HY5pNP0FWwV/YvxZoJqrjh/3WDiWURf8FFxzdZttw+iKKOMbIN2QCs9YEZV2UBwH4
gEOnUaRw4dQIesS59W7e1Ju9hS2ux2S+uMvOhGuOqHXMOC4E4Qf3hobGfrFPCu2M+meQXm0NfeJD
SbmUy//C9FtHh1UR1P7fSK9XzsCguZi/JAIF/tj3zRF38Th12DUhk8QMqQ9J3lK739dSos1NjE96
M5POVGaayRzftdpbQVnvkNVehmxAiI6cgLy4Z7FVVCyAsjpqyfapy34oXoifJbHdvQCqMwK9yDLw
pzvDVdqlmvw3T+Nn/Fyiwue2qH8f6OqT5UMjVaRvxfrrFRmUwV0OgBvjLBpKVERHxQaL7NVJvgEQ
ExEkXiSNlik6gHV5JzrmKAR0oBJzFEnzbtwoOn3XP2t8YLcnxzQNMSarv7rRk3WhDLkIOmJxg4zm
mqLUeq/f5Q/DMh9r4wHWv+NWnvVxP39ktksiYieHjny+jv8Izw1a2/e507cXKFUDOzW5N4RkmO1M
3dz/UwZb1Z4UcmM+Z4L2BDu+OofATDok7b0soJ9UJkbaBXLx5QcRYQMNJW6vjtA20gR3Hh+rrr8G
NmvX0aD+pvea0j/TRzC5CKDcXFubJHAnmC0QGirw3A9DPWYNs3/p1u4weZnSvi8T0XOVim/fXlrx
ID56dhviJ4BTFjQ4s6WuqUGa7VSYbomFla45P17P1zV00y1gKvWUeeLnfCO4hDUJQAMMZzAb1cZi
CKMWehGQdtGBilaJ7DVwXRToOSho7UtbgGDiKDH2kAmlamI0DryjPvZ5+UuiYRYUjBgfFHsymfB7
JFYxfp7Zy9ZE7Fj56g7Ch3jvN+QIZ7wjS/XQsDCen0uAuwHmNC3x5ZFKjmUOBpuAJy4ESbKfqwgT
5iCXnDhqtxsylr18JCw3x0/rqNhylDtVaA7A73E8UmXC0f4ZT1ZVCQfFM5TJ/9dBSZBnZO9E0xBl
VupN5a/drx6KT5Q58x/ssp3ITTr8UAa7Ac4/2jL5WfgcVqAQ7qTH3/Qqi5nOSTfaZOc8EVtatK5N
lZBnFxBFLHNOYePcReC1Y4AjicQtY8h3p9Pl9OpMdVc/4BibU/+3g6LkQH0ORMp348CkFXUWZiw2
qB6V1RDsv3b163IX9ypc/WnjBofB5ewuzU07sYt5lR1dvoOYWpADMDHBuuy4c3QbZWAUCZKMyC+t
DFSkV1oxj9bVuXzzP0sE/B3x3zVMpHIjWYf+ZOXiTCko5hsd8N2ohRgP8o+wrpn40ID4gJegN8Tl
6O+pWsCdYGcqU+8M33ofhMd6eGuERiM0QRUhYhZFE2pLYH7qSDNvd3AYDrATlKh06iwcif+2Li6g
wpgLsT80SfYKxVlD29yoJtbh+pRZZ1LSC3TenCC2rLnTGIDNy2ItRyXr+GG319oFUg5zCmq7tltA
nmhM39EpYWa9w2Q7a0isRxoxyNg8I4g4c81mGUTtptBTVBEFqpT/0xWEf7s7/VFAv9myARpMiowS
zzPVYJ6O5YuL/puaEDF0pMXDyyrhdqpqbc5himRbT1SR6PFHSGNxJPzs29UTAYxkR9BCis8NjeVI
luSCDUA1icyUIEqCjRCQh9bwenZhnNaAakHHWypUCnMkc0ubsP9tngnZoS8uSnyRmtMCTAcbIbpk
SZExlxnIHQzWed6nL/fKU7XgYvpjDKXE/9B3D50AjVlArDiayll7Q4TUCQ7fTVAsI1BhmhUkaxMZ
VlUjZyC6emcjCp4a1rPQ52yrr7X2aivw90TFcS3SGd6+MY8pwLM0HMIJeZK9IaPNw35W4XN5/Q3Z
2GWDeTfDEDgs8LYItbmOI6lOeMZnEbKn8K5AMNKSZs5eMkANCYnZV+EXrWLXKJWct0tOeiCpTx2G
cJskdXZxQTKRRot15XtBY5WycTepy9hUeOdI2Hv+1vosbr426OFKy3a2u1hsEZZxTzmc8h4OYXkW
76wpuXL5N2mxwRCkB1MjD+M7S+CrSmMkghYKY3hv5CFC6LqMP2Ax+s1b0DMETvF25Qm1UFgNeLfa
OtY4zrSxyN5TvzCGe4qcSpN/DWoYyUHXFQHK5xF/pTrPOt8yBx8rzxEZG9ETCfuP325h7i8gy4sl
HzR0dG+uDePh1UxQDvzx7Tr3ZkBo+XLKGSEuN5lp3oJ4Zr0qTLUD49GFAmxfxs2T2Us5LqNhvKeD
8+3tGOViQ2Bcb+Y1lldVA1zDLm4KJaJFDGX4SVdQEZao3tb8ieG2InZ/y6Mo53zxneQxuvd1Ek1L
CMuMBEXhPJKKzTUPmuZicqb7KhCvqcK4DxSTpnV3SX58bYbmAz75plK2ehri2FjwFoYca2LQCOMz
8zx8ugcN5tGBHEAhouwZEev2KONHGcYK9gZQ+rXAMszpnQiFzm+G7rAjd6wWkLVpqHYjn4XUi73X
BrwB5OAl8ZHZDFkyyzFlGgHEYnwRJ8149ZWh59SpiT8Yptupnl5T16dsILCu7kWceFG6XCfcqDMp
g/Z4CWY/mtQatyjWKuoA5Zexo+FD0tgTVo3aZpLOJUYhGRadYa67qxZcKxpl5VgvvTPtnpjb6Fem
T63UEZ9E1vdVRZn+CxKCwHoqCBErPL7Q0jKcUaO8o159i5uPRoxVs0Ckq16fzoAezRTvUctkH5F7
iMIeyiCRbQAjv9S5IS/YJMCT1nZlCB96Mmogb1Ii6HPB3Rqf9zWwehXjhlu11XUzO2NxWS5dVKUC
WVIXhpJFnQ3rLXoKnDvOnJj5xKJQzzaibezhV5kw0pUjYsr0/ERG4BY5t33k+MNSyMt4dO0ZjQkg
ME2rype2lU2amrIodrJexqFvMaxsI0xpIQ7UgIvovsR+32qmtwJFQv6ADDyM1wx6fy4fbF4o9QOd
dd+7ISH7oxFl97n4Z0w7XMzVkHYVhkefCGxupik2FHcmNZG/vk/VRRw7084K5w9WoIfJb+xo9OAd
+CGrDXIoUnI+/i6Cxt/DvSmssnJaNariaBKOkhj8wwjf5jLvDm+5vZEZBuSHr2RIxW+TtUikoH9u
T0Yme7MFsg36CsHIc0Zj/FlAfsSQpxPC3hiekyki1F2LqpgUdZHN8Z8vXYgOvCd5byJ48+FLhpYq
s8KvQ04DMX4MlZcdEwM8/vG5dyV2QHcSnoC31IgyXRqp/IKmKv2XXz+ZdgZVyYcykQyAiS7jYxf1
24prm3pdWhtniuxzELNpZ2/d0coGfURiWy1xvNiyYeVfTSe7ISlUOYRlNIMDzGpS/J1OhL1JI6El
R2uHHToGPBVcdjX0b0WGFb3zGdRMTz+w1OI4xvncnHIvy8RXWtvbaiXPRjTAQgnNW0Qs1Ueb+MvA
+1nsg35ghxK9WjhVm01tnmQ+lUysrfbFKilU4/j8IORQQCp+c9sEvHTYbmDENK68h+oLlIBVSswA
RfLMlE+C73TgUe8dBSPl4NbZkR8phK8bXu82JhVhIkOVGaCjiwpBMbyEr798UBhyC66dt6t4mfiW
jkMjpnRVLdqh3osAWCeV2FVE6y+QZFjAo4ZeMMRTEwLMx1Ch4xpW6O2OUmG9xUTdWTh+z85geaSZ
a8B3q3VyPFlUaTjKrAaqS9yahoIJqQcWAMNK7dayrLvwVL7naClqetKwX8MsQ+HDGiYYkFdydx+4
txjaleGvLVGnjJOQxGvvAPgG9kMSgQY8iExFFZlP/yJNwoq8sC48N9f77xiBvawZnxDnPpX7EEj/
vd3P2PUp0oQfH8JZtjrxfAm0zl08xoN62wC3GbmzqVjboBFcScBCYBb0DUvRC9h/D6Flupcb01ld
F6CGh1H/MGxO13mlDHKhqTNHspvqQ5mZBpq+N96qut8xFpNwvdxxkmUTM6jjwSnPdmF58gjkj4Kl
ymT3hEWasXwcybGOzZaDm8nPnzG0xkQX3Za41MzeUOyLZeFm++4QEuqMjRUgHgcO3mAYFJzbeqtU
U61Z5Sub2EU1jJ7GTXgUBO7PQDzetoIb6A+Ps/M2hpUz2776v5YtPN1iDokElDu1+vTajE1NBZzE
Pwfq/sGWe7bYzYzQHAIIxJ3JU10uhrWETBVOFkuEFUX5w4PXSY3/Ju2YTj4PgIAEsIt1Ut6RDPSW
kVzDi+KCRrz+KkutU3l6ge1/sHBty1pHNh7NwdjdcSIVmmSPXssMbN19TUrfffcDbXJVXWlCn1Xb
tNfE156slY2B5OvC5r81xv+o31pC6QL/quvuIUuppbD+KR/Umh/rGfdPWT8wZZh2k1NSSFxtITyA
EVDUCaW5AqYOFdMIa3LDR6AF87SvutyBadR5m65mgBwXLK3UZ07r4+4w34Q6pmAPrF0oNTvOzogH
NwNT9EhyI1WdxEtB13eOFEpgOfAlQ+iThgxP6VNVbrBGMdkag2txnNtuJ0QnAjnxslsQX4S/i/8M
wmop8pFIgfUapO6qdORNwO4VqvrBpC3/9z5Wkg6jn6irLrPNBuYcnIVrnGWesAUKNkol8QAcR1EV
CF1y5hRr+opHdMigwmykJYF50ZpoE1+/uw31DecwyJRTFZ09kfhUuAKySm7gpjMkALVytqXRFJ7h
lLW0wN4krvPK5bPErabIXBHbboqeL43vavc0g2HFRpCid2d3r5O2TlfgNBS/uqn0FAaAOmMhzzzX
D2z6l4WBK4bNVJcu8cxnRg/EM+pP0aYP9azJU0tJ7gl7xxcsa+CedSFAvbhyOEcWK4zrlOwzyPn4
W+Y8bA0cUJ0SQKf/4MVb+2UlUMgNd3iHYJo+zq/y1Mq4cbt57iE355svZzv6I4Hc7+7tels3hJeC
1tqm7WuwWV4Y1PxA9BkOeMoqAGkf3w4pPIOReq23eYiFP5oqhhvD0Kjn70rrL+IqLUx8Gz9gvaiT
NTotmvAo9YWw0Zp7jDupkGwZSm1FnYJUKOc43PUtSf4aaRdqvu6KLHFYwX2W8Cx/PFWIdQFwXpHp
CQKDFqNm7tAaR/T8Y29Q9/E6qalEU1DexX+aJ9mWMdVv1emZMe0nhgu2JJhYVoGYwhQ5pdG9CTmu
DrrSOp6x7jYaklPiF+tEcoLwhdpMLBgqmATO+d2Br6JfLkEjlNrOcknjV0Wd1XPqk5Zauwx9NGsv
gVVOvF8IBNnMpLVk9IqqS5UIdC7BhX8wCnbU2g3DW8rSZduMTqHYVoPM0KmPrWfhmXa5FEiwO27x
o7FZP+2VxLKRvtw84bwMw9ioBrFowOwNbuC5GZn8jyMP/agiV5oLmTT1ib+zb7TR7NwSIKSTHbj8
DQjkDV995xc94Aw8gjlufEmmN5F8DfSmThwtlynIQ276t7Cb+UW79PAKw6Yct5fpQnKWtVPFquo1
GsunFtS6p2LLKlnKpSmFl/elIvsjfFbxCGdHpbke1vAppRC3BiqjN5c6dnRKpLb1zB7gGzNF3AHx
fj4Hq20S9w+UoPeq/zWGi+Myrisarf7XX0I2bL+U+QvWZyDAw+O50ZSAk+Cj3lWlxPlZSYeEYJ6w
4emYGT2YXHwPLSUyYeics/k/bONi119HdFphGaZwAzt0NMhC5Q6niMB1qKgChemn6q8dn6nSQ7sv
xf/2R5OF96VVe43KD9wHtQuDOWvOi5HyOcgw1bW1yEvHJmW+cPC2MZV0To1kaO3kOgAKWMBCKbJV
XCan6vBop57erQwdVrKQ6sWcSDxWp49NHXmPQpLOakEwIK/GbBkjSu32TYhAKso1C+yBeJmVCrHh
fy+H98zA2emyjwiPn31gj8/DG6Xre2PTeoaFRNdNd2BM5Z0NLr+OxeifwECdlAeAVsdmHmiFqt4y
qQSss9h0cCN3+rD/A8sMexhju8ol9L4zkXvTnW+wScSEMwUSxEm/fZe8bmFDkCVwZI/F9BvSdC/d
5T+Beh97A7njvvwprxo4LOBDUrDte4AaiVzwjrnitiO10Bghcf0egOhagQazR2MuSPoovR1fNDIU
hOR5UDBjl2Oc8+7ZDbF/pcMxI2wTOiN6HKJo+hF6tjUcxBmokLzHXxlp45IgfjkzkwD2Fq2/5piE
wt7VqRhqWADmg45ia2Hm5hMOHyjOmcA23lodyV5VjNimdca3bmtMPVxGHBdmxjhJQG6Rc9GIpdGJ
SopxIVyYvb48w/4OmoP0MM+p9RluuPASMdHVVF5mPN+JvsEog+qPXCzxTHWQLc0CN8NdbvMBtKR+
QaVA6P2TbnCl+v/mIgJTV3sFt0YU2sY0twubomiy3kyHgCEa5QixpP6FeTabOtGaMMqIkTMkQa2/
4gr9wPavEm7Y7awxCIj3ogt6nw611smmpEiICM1dVH5FCzR9MbQrjqPHTQlpOoERqHidc2gPcR3t
h+ik0cA/8ujGUzMp3MYRcST7dAXarvtwKPXoY0geulmEG7yiXUILwDB5NeB4XfFEpkQl1VN8YxlH
EDVU54djCSUvnrZcQIzYm9HEBvTmcI28eueJ86VZn52h+ju4TuDnsAAX0NNU/ZvHrbwdXpp9p/Xn
k7foZyGE7StXI+WU4C62dyTAL6RgQmENaf1EX5Sctv7YPdSnXFACgYXdroaD7Hb4Gz57o+94RcxP
zF4rF1+bKZIj7bKU9+ghWEXrVRDmAqXByPbE+Dbe608YknHYDIWryalP9Azbaru5MBLGxn+WZpzx
rfGs2mgW4FqjO32ubOwP9/nWaIhaTKiS6Z1yrvkZByBWkofSdfgohrEVmdCL4pt11dlncq9gKop5
EFcqet/4h5otpPO4lJKh2y5DbAYOX4EH+KSTe64EFrY+ga3jNw/J8mlxires/NcoI3p45zv0SZe2
tr50L+UBRXvmbLNoNUXhMWqrCtKTLdE8+Xt+xAW/c4BGJpArpfVh7qjFhr3JQkNdwGMXxg4LySvK
Vz367RxZ9BWdjfgmQXp2iIOXUKHbBWiPKjxYfGTVjmLyAJiWjJFGDbaFU6eJ/oxINEdEDkWspgf1
0MtTTACbEDvifV8fjB8r+Q3ccsdj6z9lGeW0wWvtvzrcNtnw7t+J4+JYauzb0apWPiOdqlZK5eVH
QImXCNDrtK0EMXezPkWfSpA2obEbI8+FEI5GomDfqi9030xgZ8vcaDsdT6gCpW6Qq6aRr+fEw1Jm
hCWLDGqH2ZxVz5mPNh0dHkfOqsva3dmlGe1WrexDnCSIrn9OHqNuYjWXQSsWoDCFcQx45LDwEvGK
vt6ltndS8RpOB13ONxCvaJNueUTnkwsMgGUg09cu8EpZEIRIEYjLdSaC0/9FT9cR41uFJlxuCqBU
yy35KjAwLwzXy5pZuvv79+OCiQg8vO3vM3qNmvO/VuPNMnSN4OuBYktwH1BS8lEsj8wm5ZWDnNd4
dEpoStgsimFmHfk66sels1g2xJm9qvqvzA63fwsW+VRJUkj8HdDs3kGylvkyc54NVuZsEaYrBDs+
IIfwqEqdUCXSCWub64LaDz++F0cag2OlsllAvelJMKI9nCz8MQW+EuXnO80LfBl10Bzpnz9/Cr7g
6O4XIG2C3Ni5fIqx0tC0ibPmBN5g/kLznE9rX5g9I5S/mWcEfXOYx3xE4PvVof5Yo3TlFXw6YmFl
g5KeuIdIIaph/abd3Cv4DqWW7ZH9SgNhd3fenibtsr84Pb6eNgPoDzas0E/nbD78h3s7cJUASX1d
TsdELgwWrY9NMrD7MDWEiPgCPN7TDhwgFOxWlrJJApD1KQWvpJrckUnlxFnyKMwnGTbK8ZMwzqnx
uz6UMuZVHfMdLtQ6HtwNeUpPWhCbP09I/KTg4XSJWu55Bom7aGF/Gunn/Ot27XoeQPhY0TKfW8Fx
GNEKFP4GOfzFzOXAvat8Igg87CCny/Gqq/OB2nQX1tqj/owtDu5fKq1PzbT1KWoyrI92Wtpk6TPm
o7S1Vq5FuQ4QJy0ebZhRjjJgfHYEVzezrFeiut+ydXZ9CHM2UQnfcw3Pn5MKki5aikLHDzBs02qR
TgHVh/1JYNCkb8ed9T3MgvmiWo356eTeznRCvhkMhkvGv0rNdYSKz7fvnywwqAvIPwz6uFrHoE1s
pSG4o6niszmU6MBaHwWL8hBOAHMsrSjcMOCHL0J3U8Hm+PwzGYLdZa15993U3w14jkLotTABt4BS
4+GKKMWjKaL68EjuHSWNbtxacEmtVrYXtVtGSJtJXLSDQmwAOHW7yErpQvUxZ8OeZ/WygvWII1aX
mGYPr4J81Zs0V6dM4dh0wkgwXS2f3krhuObBW385XnHpkK+AW4koSxT7YnZeYSKQxF3B8OkhuxLR
y2Ng7j90XcHcbsUyOth7fYAyTTQVgceZI+rQXrToAkUuu/533XT3Y3haVKEI7dcoNVDhFy0oQY7Q
mJRlX4NcyHPqmQVvSGU1Eo7Svk5gukQeaCAno+e7pFiIXBxeGpuFumZCn12dtZkFg0MZycaeYr5M
roOJc8T9rDE3TC96wVX64SO/RHuui/Ha7Rt8C6wQEHOr89UifvolB3adAGVXaX521WBZqAJPLnOB
uyvDIZpqStKRhEtocoB28mPVkvtIEzSb2P5JoCEN/0FeGjhh6Z1ILPPdHxZiEtJfoYbXluhmebPy
K1xbCugjAyJt/gNWpkIkNDAmSMmsuwRLxMgAZ5IKYhHnQKXNkiH9M3PpCvx8omTEOkC05G8ZBZE/
3D+al8v09i1/f8Y/zjVOSF+i7zYdTtX5E4vCZGjF8RvzznhVmkWkQHlxKSeMOqYNtkcBNL8pajbv
2o3RshHpN3Tz2BdneQISu9U8bCgEFCi6+PaKk7+U37q8DtjzNDkA+2ptpp5/7bX904fvTrYRGckr
5SIme5A52W4tDPpjilqZmNBbnIyOFTI5bdgFQ6+bBjEdfLLan2wjF+0gGI5HfTHrS3ZyX4VG1N8D
gLZM3UvHAtIsbUnYO79adLiGHDDZwJ1bk3DmUksHrgUUX7CahX9MhTTmoNF3eEp8Xu4zKSmwpYkL
eDwnV4myL25a8OJne5R++64cyFyl1aY4behUewrzltNDynpPs7pzANP/pwy/8yXRKj7BL4Uu2lXX
Af6wr3ht0+1MgnzjhEVg7ZUTTAU9Qkt62pT8AigCMDi/DM/Sdpt9dVKOj9aThSXeRjJmtQzLPxsU
QXBiyWxFOZbWpC4Tj2BjBIcAkMubUsAnslxnLS76IX8Z46ieOlF1deFfv9wA+ETIMiq92UWdD5iq
m1Ok1NMwJWMf7WjpzIu1nEkjfpsWEqz5MDuWDnQE05Qh4c1/YLEjsVLzvBsdq3xKQOmqHhd5/k1n
vW67D02Q01ET3z4Iriy/Sr0GUXrW1YpJe1WaVWrPgIUbFeWbdUm67wW4fihHt1fRTcO5VcHwiFjL
I2jfKAlSvkbZmo46LJBGcxVzGqXGnQAsiVGQrCACgevQ0MT/bpei2HrykGIbMKBmB8N9Hvyxfdhn
7i8qYpPehwgHx0j8ECGcfGJVUS/nAGqIrAC/golgVoNGy2SoqNByFmdEbV9RZPNzAu0G6pM5pz3+
DLYZYe35zuy9K/6sBdN8jCZNOaxtid3W2uaQGdBOMXCoSZNQs3Pojq7nHBEcJ2CaRqgdt43o1hMx
9OTOoRzThNj0t9bTqZF0cjITxuOvsWdbtMiiZjR86AkZn1MHiw3wD5Gf7s2SWNXxToWRwWUNDR72
wv3a1NkEAwd7acYsNzP5U+hqdyft9viWSxffzr+Fev9xaiqCMbRFdsIXzqqwUy/pQgSsza4lsp/e
QIV+toHZOM23UapojeQPGmeJxhfPz/c3lKOO062XBVfPJbCenpUUBOWM/ULevKWTt0RAbn72Eypz
WhOEFyDdGXrrP4efXGOThrLDMZW7f1sYNGoBZSd3iWIywTmuy9/eBUG72IHzrOZ6sjq1hlRFMbuS
qxO8qOccBAJo6e2p8JhEoxXktpCnzegHwacFxeK4Q0y8m0nZjwZLF5/UMcY1Xz9GIzgzY040ljVJ
TYYLX4zR1A6sgsmFqpEetPRv0ICOeiunX/pe1bxn8KoeL42qdNvxMW8QmGP7bkhjRoDEDtPlF4/B
Zfkh6XOdAwudTDMO4nBLwuPLAEMaoDaTCf3PSY8deVKlcqVJ+q/Fxsvbh9mpl8S1Jd+EBCyEGFyC
ZOMuGSK+pbJCIYqbSjK7xSOPo2DfCMGLKhALe0Dn/ZmwBIEttroSgm+2kat4pKmdPIZVCcE+HMbk
RawlM/oqOQwaD96gjrAXln27PHfpflvwm62N0Fo6jW97/VMx1AO48uASPDMjfTEyduGBPMCFqHld
jtXojDkWQYRYyn0yMkiHN+ADNRPl4dMdKpP3BeMv9+4dfVvRabBpS44W6tCeaXSpBLUzvKwPobS3
wny44YygBkfz6F5Vy0NcmE11h+0t+Ndt9PrtFPtHW1Is2+1eoS4uRQxEl8h7jU904tijTnQaa//D
vDnpdx8K97r9HSeB+UmQNvA0I/l2QfQUI3p1dPJpFB7SNi6jyDUwZy+Ky8aDFCkNrv06eMetHZtT
Xz8Pl8Q2krT45DfvW3LsRG3c0gyekHX0aVduTbgByWL/sLRFOkecJt+EN0AVEgOo4TkABBwrOcmU
I8nMviLBlnLZyk7R2aaP1gkiizkJMDrrNjbfDFs0/j4oSCUb6tNQfzvSvePDsDPtY2meCHJf5TFC
m738c1pZQJAywv7TK8LKMyuyA3vm89/TOd4LQ1UiXOvaAjgxDxw2rtxJ9d0HzGi71OnlgTirKlNu
Go2OmV7QJzTVZZxZ+Ysjo7zyJ+aEXuSzyBJMjMNuqLayEdQqfsb6jdefqyuEL+3omHM9fOdfQJxI
MWd9ddE4nDOjVcnrhNbm+zzODKaBV7JWoqMVDHdWxVJWq1HeJQOX6ZKdf8boKT+CJt4WQnhEjRU9
KZcpA5X74RSdxyndSKtwgSyd+kpCKyNOc55Pvh6FsPZq8YBEToOxnqrR8myTnebeXBTuX1EvUH8X
flM3xBB7JWMLSiqLEDyeiZ8I5fwfSWdRlpgaoQ7PPzpfZXD4lQkCqDYwFNunK1f5XsdoYrmf5VC0
P7+NE/lvOesVMoXu12hpxEp0yWezdQu2ay1YX1Q4QFMpAmkTlW9A5FICruW1sAZSVB+zpuznLwlf
nyk2ExUw2BRtgxL/rp9lFCfa9edjMR9BtmOCuK+ZHyquwI5V2IyRFV61cLuW8ONO8qaZLCq1TI8w
4ltf6zDqIpKr3xtitiy/ROVNf/BqYx87hNOsJX90CnJaO8h60vqfU7FOlldRJ3wZ/10sM6B+vLoA
+CfMksbbC6fGEwEjVW4wXar6OJtpJUXsIYRiXONcFCbDuRdYE9TozIdLtkE1GqJhQvby+PUxnjbI
hMEegcfOfzkR7CJHT2aj2NGBh57EjpIw6HAxlCmJbdS22h+6WjdhbWoC/QJLpSNRmTVqB9wEdm67
TZ+VoPEXiCwXFWEJvskmNonEnR2ce/UnsOQBbMo5UdOeyCn2qdFaRr8V8KWqDyBSnBDC9oVEIToc
QAW5/74ZpNzNm4wwwUELtcJa99fZ1EpWXBDy6uWtI8N3n515vTZkeOakn0bmP69T5B90va4iw7lN
GS6nk8CQ97sBaLHK/1gPhP1rZg4GQcQACg5BaC1/td9NJZQtpAVkUEWl2lpkqQNv9WeT95JLqbDF
51+26E91kSKQlXN9U2Fs5YdW3062+bzwOPdqxW1aBJHbijrmEYmGfDc0M2zaIXGmn0BfexkpnB4P
3uyXSP0XC2G6vLMfwvB0n0bo4SodrUM3ZnZ6Wga2taL1zO5Nd/mOKMNqMDirbjl5lqq4697DSvLO
jc+NPn9K5o2GdBxnuuL64THfEE3cnq7ebVp/BJY/ER+rlOua7/gagQLUBRDu/IfuXXk9I8ZW4jMg
ZJQSdFV5HOEiLS8Ja6VtHktdk3DacGWKzHBxT5RDBZZzWAX7u48/LOAZjNjVQ//mAMcJGx7iskhh
yTvsdBoNRibhCjKZmiB6wroXhRjGdyP5Tz/ZZEvd4DYODVOznlUJ9/S+9w3oaBbhS8zuOFL1viif
YtgEJ1l2/Q32qk2H+JtVBA6oTWcgSyGUDSBScWyg8zGozVQZR9lsF/tHb4y4CdYAjLKhOFiT6y34
ohFMe9g/UnC5BOHTEBzienjeB4l0Bv/POY0CW0YD0Qkgb6dYo3GJZK1tz3Ybb2/E3QY1y/rqZK+O
ctRg+O94FtYutMsghz7d1Qh0hsOso1tCyRY/u0y+Jqt6no4RBa47kocghTtaDkCiLJWEWC6sYsjD
q4b137JnT/OLHRPSwB8Z2kDXFO/P8cj2ZUNUWwOG7UFWVziYrXzSlEhMKr+ja1AxuztdFERnvRBe
Z5b3P1giAkaQMkNWX3hLXyGF8Ijq4wql8lBge+l0NdNHKaXufqv+W0ohiWRlQpzC1NOcpZkEmFhD
J8FRKIqRlsUv2Ojh9BROb1oFgVhZuPP6Jt75PdzbwVH+1k8qwJ7LSYZBglRtqQikdt0Gk6hTaiA3
QpaL/+LU/WDQpD2iwsBop+K0GZLWdjig0dwAydAWluRxgoEv7fqJB/cUoeU2vHU1OtdtDBM6tpVl
jr+FnPdmjwlq0OHt/0t4agFV1I4ihtl1xjeXlcNOjCOVp+wdv0wTz6+HfK25v2JZfoyuvFtoanam
8SpvmLHwHQcgGYjGvu3GnaPJwon7XckhbzXIkPCarB4E11m4lCKQDjQU0ehA2mmV8rYLXF3Y7gRe
pD8rbYX5oRzsJkgMT5xiqzUcJe8TkvnaCvnrl+DPNobFiZa07SEA2yCax649ZRQXLLbQIrIOB6Eq
LZiRVMV9ddwk6RhAy+l+3snATV4ll9B9IOUwrO2bpCc+gJwzfQUl9KVNhPAY6pLq9pYhjNgkzOVX
MURlxSkH7M5isKP+BTWzmbtzNqoAHliZqJggEOFRoMbjQFF/HvwvUpbH63YBC8j0RJAvbh+5p1Jz
Vjsgm5teTAyrGwqGVcWOfHnZCKiGUSFH/F8IXhOxsRqIEM+2MCzwcZvzfI5VbJ9HMa2S4UT160Yx
m5+uxmxb4NNY4ZJv4cmZ18/yDr1o+saC1LWGRqxBbrdQ5gP2R0ghyTOXqulKw8GHNBLQhuE4LaOD
ZI5fLt81RoEAUMpJHinzn+rzwjBYNj83HO4IAwLYypBro5Mz3b2GHJSTKJtw1fgqd0Rs1RSun6r4
W6WRFD/uegm4ePNOgwWjXT5Fkx31fSsn+UUl+RFd2roR5KgTHckJVHE3bZFD9B6XLn3HcteE5sNP
IsAI23ap4OA0W5N2fRSCthbAKf+cEvUzyX8visA/Lqn0LWu5NYrYpOlKmAF3Dq6lX0ZvvST7/BvI
CoIjiG0wqLi5LATgiWkqg01dJm+0Hp4e1hYIg1uGPGrKw414mPimuVQg6gMmwcgEB3wDtZQ7PuR5
0pG1neTXCDkDuBPYpXaqaXgkCoOET4pmdWrBAxn2ds18sG+KtZg60jtSOof6TC3dFTKXfd4ykgFj
yfDLGJJ/e9JPouRFQOslfJXOCTGENVMxjJcGeTCS3xcGzoi1SfhhASYHMXzY+ioNTSTDG2cOBw8o
cF2CRwuv8IgH8HMMu/+xK7d0FXfu/B5Z6gLJZL5VDd4E4UCiRlSmIwNEZC/PPwImFPAh1k2mSFDO
gaxrPj91bZgEOg0T5ito6m3DhMPdYua/hoAN/w3xj5ZB1PZORvdVoCgn+BuTcqArNa5MhStNk9VA
zWNZUN2RWmxgG6aoDWvH97bFu+KCu8Jjaudq9gvah6QGdTPFPLFCZa05b9q+5awVM+6NEmJC68q/
7sdVGOi4SE3pgFp0UPsa5pZV7LeGaNz58TD743bj2ev4pwsXIdDfpZkKIWmsVYy8nNRvihAFBBu5
kFmWj4OoNNidhEhiTprz5GvAF9rcwomyKOKGl2haGoLZAQJtl4blQGTfCjibu6axV9i2t6ku/89O
iRsw0Puk4wKxzJCkalmeAw4AwW1v+pmFCOX8+Fidu6hU6Kvrks/kb3e8bzUOTruNcYV6bEHugVjX
+SznpMx9phmF34qp+/yDZ41Lzz7hF3P+7RI2zi0ZdsyeToxLwB5j7dBn5t2ruY5YSMEyjiMQio1Y
4evVuahjh3ENn8dA71J7Thvm9I5hDiXE0QxEQgVVXLZ2d6tTo5EdeDSEuJ3Sc19JSsn6qw/1MOU1
EX9fCxQKbjHo1dp7t9YPIoww1C+MBZ8wLZOtYsgWmdWUJiY5EsRbPkxlgxEkAjaQ1YwIPfZkrQWM
YC3/LFttUEQc8RG6C6rbnO5y0jARMlVlZ7SXLYqaOqxHOyDzHPvbgJc5HX9JQ7gj5tlOE0NVeDw/
rGj3jz9cfFScCT3HNlU69sR0xEGJUBz/AMa80KtmDtS/nekiD4w+E8cUDoudnZHo8tjeun6asoox
e7f6HtwV453jZ6BowgjbxAUeJqiugXzuH2pfypCVgPWhsX/alnzEwBsoPnX026qInc8aGMhv6GWF
o3v9DMjKsptiv+lwRwS/bgKFan5Y3+78huE4ZXVadP8Bpo+D9wc7EM1FykuMzyTAxYqYI+YW1pML
yv5bcwuaoQg2l48oGTip9cQNCdWxP6IIy4IY+rZzTOTZ2Crq6RLmXh+UDlOtywbcrO32ku4sEwW3
Byaw2VpPUhSNmLY5v2nM9f/7tPv1+tSWzX0rn79Adc8grvXJmXqwdpEYYrAViEzVe8IeRr85MUrR
P87C2Ml9A9MhyA5RbKtq6yTyDCq3aExOiIy3pcSWbmIFTdL5PxyxZapZQo85nEjDQKE9KKWlmw1U
QRAehKWct3+0sDqX/h3ifpnLiLtoG/LW9mNTmA2Yke/1pZMDw10DvOzrSwC9NwFXYcNEy0ML45Cl
KlNIanTpvgLOBdfTDqO3a5WC/weCO+t9ZTrxyjdIWD0cv7BbRN7/uYDiha93H8zsuV35sM+GK8zA
4GVJlbn53Gc5Qm4+sz3srGR53IS1Rl2zyqyzxqnOs5XcuAPel/2Vm94qLf9QgrqhUcA2j5SohBta
DsDFn8NoCDKVYZmFA27MvDzemuRGUXm5GP5Ag4Qq8tCVridIXv+yElPjZ6N+BPQzJRyviKb4Xst3
tQdwa7CeovADE02+oV4hqL4so3vBj6CaIKK2WNPE3pmPfg1boEhX7qO8NlhJyNyn3kQ/umK87AzO
CDxYKiK1zkPMBnsIMuzoqjgUluUGRdxp2I4XO4NbzWVta7N2eU3YDEYTW9DLTLas0Vzg6Q9I8aNR
moRtXAxBa/UbZ045aSBhq3MKNqAURY4Z5k/dqAipWx6fyL6HLiRSBUj3Tf0YeV1Z+hwfEiB8qyv/
gXL80Kt9wKhRApHXKjT1VdNAvBHrNY5zdjz55gmxGa0CO79XaJ20pOkovBSZTi2xrNHA3aana2M9
A0IZ4lkpcCkEb3pSKI36I+Fz+jFsxVZ9ir74+y0yx/kFTP0Cq68tIyuIbgPoYFttlSBCe8rwa1qY
Oar0RIoE2Q5bx0zGmK45kg2fwNWur68/5Md36SxdGC2dDTQj7WPEkJ3juRItz9PfAKtOgMv4EsuY
wOC6w3PTlyGqjhIttejv2Rua4KHKfaLuPuxNKppfi6pyySMSE7rnxezkvQBhIzOnlOhvfMIdKw5G
It1ZG1+FWpd65ZKmAwzRLIoNZUimuzaPC4FIfPGuzzmaeoREH0E4oxOd4I10z0NKH6Te6ev+7Qte
ucndzmviJrx+169cTlimYUzMbDmLX0gffGLWqS3I8Ja+Z2QqenIeBov0S3vc2hG5x15IWc7VciEr
g+7dwXD6sqyzOB2wTmOEsoTA09pABGSoljI9/OyUaajAnRlkDTip0MLJSPo+Fo9BXjS1pJnfcbSO
7DPaVnu3f15m+3hPjqOqmNsdLBMay27ImFlWDtZInLmLM9CGZ2jFIH7oI8PMy4ciq2gmPXRLL6aV
vJ5EMxO1XOyplw6on13PdJUH/9GFB9uk1961L2jvQKW7kC9Y/FhWbCm1CTRWyXJk09qAoqNsy4i7
/qEJOdkSOA2ZpR+NU+kn7pVLr0mnbha5L3uCUQLuicuZ8sOeGbWnSRUrCkGxfh3bxVHgGz4RIoyg
dsnz5Y85OFLfzEJVfkzCbRxv8bzatTabEvG032/zuLM4jsoRkhNsCvPpVTywyjAmxJRU+IBt+axx
DzuqAiRy1DoQ2JHnRYHNR6HZE6Brk4NNnz/EDXZIxtm+llHEKWQXwyTKAhL8+mAhIAlkp1xl5ve4
yb5F2t/FQIOMKmpowuIiximsTPT2KmhMh8Ta8OAs4Wa/3DyOazfaru/VJ/ZPhOjvsWmGoQnGOPlD
6cl2Hh1o5hq16m9cFo41xmSx00R1b8bfEqPA1ihTKdQjUfsDkqTL2CAlmWk5PFuzgXmNv7pbup9b
bFraCFeE11bg7w0R6ZabTdExcIQtp2/g6ECuFL09mHqjTak5I2pRh5LgbcSuH2e2Hs6h7HEBVrsH
QbRIHjfLw9HIuJY6wTcmzwu/Dhbdoxrb5ifWUABFyusr22CJpAxyltl2GTuYDdMotzkbpuFDsVS1
Ye3okhh+pKoCdWvImm6QfRxq570h/MG57sJojBIlZteOy4TjRDo7Cz/LBOtFD12nQHQUv5psXQqa
rsF4I7GBY6ycRQvB3Wz2ltcSpAl2KxuegTw+iHzE2ZmlUOJudB6SLSwAk2am1mDpMof8Qf+ZgCov
R3rOZlphDqtKF/7Yh3diTM3AHTmaJH448LXsq8IJLVlO9TVZCtxutgWqsAq45/QKZarXj4UqLY17
3OmX5gPfMD40I2g+MByn6Jf2bYhBUHmjoIGKGJBM373O3z7p08+dN9hLrB70cMdj1WIgraZpLB2L
yLMqy24/8ItiB1dMxAX1H1QP43Oy2uPW7gj9BzZITWJpWtAlR03h9Cegq1dNkA1+aueapnpBd9Dz
hrp3JB2ZsSmOWk8N9OkM1DcloASaWuDv4nj9c/GjyPRAGLuxd9G9ufCmwroQx5mkUBd906+7xsee
gC5PAFAGMyhvBRCUkhbP4dICPHE69wjHsMrNFmV0gfmZVc05xLYNkwl79lbPTuPuQXBnapTqfYaX
wlJFYBePlwt0MuXU69sp01DzZQR65E73PYGjd9lS7+tE7IiNWGDaQuaSpwRHMMJvNS6CieuhcBdb
TYhifJGMrfNfEypdsQq6cKYXWsJ6PgUXPsZUAX1auVEPjE12OhBl7N1uP2ayWkuD2+hyuHN2MU/Q
oM0BQiZN4F2wTfboYZthU3E+63Thv1Rt07wn8Oy7HB/2YpeSCK/tgajfFpmX/5je/Pb5Eq/MauIX
KTGa6tAri8gDG6jFKY65Yo/dEN5hFns/pR6YEHY2tb2HXn3d1TmDqvCN2epdBUtZo+zPd52letgi
5rNa8xzNOjQcFF2/ZgVOFO9zzfNENWm5wr3Z7LQWSO6mhRSSCUMsuqRcmJ+Awy+v3uAZHw/zgJd7
nfIb4yBlpNHl6cGQHAIhjqyNU7JloSjgmrara6PadFt1QL7ig1caTbgj1OKysoC7eWwVChHrzD+f
0F5ySel0YUsP5auyfBKzbYnxJBFcElpzwpMpZmjB/VR9kFTaOjnzY47Ni1u+QvXokb++lOx70HQg
QpA+7oh/y4z9hkP+uUJ2k5GRMQ4ZOkKRsnRNqHIp/DDm8f3gZwjjuQiaD7ZJMpFF5KDvrR6QvDK2
jbG0lKQrQoX8MPTnnv04AwHfyFaAArjnRcgGajAOR5nYzI6FVGMPIoyzJAGyU/583ngboZTQ+ArO
sW00XRfTrj0tUJg5gPfKZE4Q1RYrDWCbrlMqCxWXqwaQLlKUklGzWvbygZOMSqagNDXStjbHyqGQ
GfXiwbYiM4aVAkgS9XCcAtMLCLFadq34IcE0jI6oh9EINqfHbIVfrubEYSA5/lgJNrIHDvUQGuEX
T7RCbsJGEbEj+I+HxDZJkVBWwQxKp/poLWna0UxNf12X5uHVe+4vlySD3gj4se3LoqnK11jVLfJB
Ly4KcERqTJJ1BcmqvyfaaS+nhrq29o3zzR4Ml/o6A1ij+CU7smt6mJyMO+8aY+P+KNPs13zSIf/U
2YMDvILYXhgDeoPAxRxKtDKybk2MWgHfdpPRaj4G5gC2JNk3iJjOLtI3vriIIz1kuM0tCfkq7Rrl
q/3dzc0nl4WE3CCvkruMIEw6hLOqnlf1QObPBNkhub5HBacSOqVitQQMHHiOWkk4YCmvttWwx6+e
w1kvC1e8CwY+V8oqBkAovJW2QiwYILCnKzpNyT2yCgNdUsgmuItd7eHFV7i7FyFBpoZUEZ/xzl3v
WbWhU9YqIyug9qHMYyqB3MAQqsPk8GMSXWmKhpUPbwxvBQ0VmQKlfOt/migR03QT9eewMolLlC2q
gEj6CUBxv/GASH5dTHckQN2usDTWerRPnPrFE7OdO6J/KPWlKcM1GO/F/HACAL6WT/4XifhVTB+G
dZTQO9fJtgGgEcEffvqaX2RVPUgrun5f7WZ1ppP+ZvVzCj2YH8/Ub11AJjql3bDrI5DJUhSfg0u1
GYyS6x3tBechgbZyx1Vj9iI3K1jbfVmxDgyDm3byFDomFA8c1BsB8mbdEburrH/jmEr2T6T11aw/
XZT9Us9qc8FBmwgUpf3sDBcwCuQEB9nVvy0oGFgQdwCD2ay04ptSfapC/sg+CjJfuLf4ZZlSaWAU
lRrknsn5gN526BBwUiKlJpKGfYSsMj1WfkHJbP9pdj8qp9YaR1HqADQV8VeKJe+KDcEW34MB7XBi
MgxCwM/4c077PXfFKXfK9aBAoQOkx6oSRhdNRUbWnlYkxoVOm26gU7X1a2sZezjm9AqdkdG7VrSs
kJncYtIcvaB7TEU8HGFI1cRqsVmi1gP+RxGwYnaltaWZ+mgBEapu7m3hyKPc0cCe2ptoaNWs0Ez6
2G/VaUOLLdDHXc8LmANeqfDTNd97R/3q8UjDR858UvO1uInIB+COncqg6G8IbIrbsNuGc7gS4j2Q
Eg4BgfNwqIQfsz17HLP7LaoKTBT0Xtgb+lKKcEZPALiICIKg8KC5PMtDYv4VsmhD97b+njcvgnHs
PhOKCnkRtqWMX2UM2Gi8SIbK0GfsNCl07T6pJK8a5F7D2M7nNhsptVfJRaNUvqfCR2OTfrq8jKOF
GiSJXRfLFDYiZr6NOMInNHjYj1AKn47TLjr3bNlko6JKS12Om4IoJx+FyrVf7Dpec0s7UErYEnJn
mpzCmvpivqrQhTgsR7UKAEbOa8IiwQ0oj+g8F8OoBTT3fjxRMbhFr3pQcmAkQmXsumQN1FH2cVYX
UqDYIPzhtL0O1mxwIDXKw9+Wi84YKp4GYinHCS4gLsqO3RBrqkWYvuxKVualOOeb0ust1jwCSz4g
i6/LzGVYvwqlO9nM0wv6dMGKyjHnyIzfwErYt/o038C2L+MRXBArsQyUzSTo8TBp7C+VOBSOdW22
nAMYzkezW+3O5kNoboeTOXyPR4t+lHLU1tzpIDnO4Vt5o7eZaUW6xGcu08rDZx1ixlxcN49iAxtL
e8tlRz3mYgN+oJLg3KR0ebXFwo7uEfCVbKF71IZJMBlmfygGii7vrOx4tEbdtzWDndza0syhW92T
pCZjwQpROFyZM1SGeOr+OD8XGy6e33VH+ACzEdWE1hOQPdv+12zH7UmJWm8F+7tNAiEvO6/WQFqS
lZS6/f+K6kaGO2LgLt2t4At/3oFoC8Fif3iXBne2shD7teGkrB3J2ZOVZXVrfSUCXW4XGvBysy3Y
g+7SdeLwh5yOGTb6ah4uJ8FzoscwfDZDW3JiCEEysfOzDinnxLhje2fippCG/MVukIOKeVLeyfHA
DiH70MVHriMWdsWm5T+qszkC+sjypt77i4DhI7w7wxs4XsJdfxXpbAqdLIz4t+dOCXvPTlG/IqHx
p00RWX8CNfEBFC3kBHgiW/ef0akPase77GrGz5xsOKk45Xam3SAfx5dYC2ZvhsEeG+Igt9YO5OF+
DReUcNptAy51g1gr2OOz0FFv3Ludn2NgWUXO0xB9q6CUskzmAIwwfM416S2K27czKOZBcH99c372
BpHi9aMDMuW+RkshsHsfScYk+rtSAYJmVVRfjnRL3O90HLiJfQVcELPiOIqoNW9YcAIUhnHNYNL3
H+34nMAXdZRO1WIO9/B9Q8AGRdSmnfF48MLqXnBV3ICi80m5X8ZRzjyY3gLNS3FeW8Ojw66S139L
7r27LQZiqYIiYSkzOGXHx9tRqTTXWrAZSdUyfyCXxgDu54MtxqGKafXIS+jOZj9k4fEIKBOIs7dY
se6weD7N0UjuATqRsgY4SZNnmnydcLFAnbZXiQDvi25PTjxlHVkTJRcT0vqmTaCVKwF6FD9mhDbD
zOH5Ejy9fO5GdyCgZzvPTiubLhmlA1yVBEn0gmGXW2YNrwQJXweAv9bJcoAdpBr7oOoOv3rq/zGf
50BcbESnJ3hZVNs1hpBpY80QBCPOYHHKzJx1srwGp7ZgzYPCONsQSQbTIz3lhaSGlfA695wXA6RX
Up3k9IIVMPT9ZSQjbR6qAwc04oqvQVE7Rod2hyfQQDYLlhfnd8f+5E+fy1dogqFh9af3Watj7AU+
K0Sfw0RRiEUU6Q9DQLkRah2MmlGBwmfsXOMW90/n5nALCWzzW+fxCwIvlTiI7rzDyrUtvkQWQGCV
4XVOcWqeVl9ooZEzzOmeaDK7iTS4C7CFwSRrOQbL/h68kFsqQS35YdnJ3MPAogRDRL377JbBHgzV
3+F+bwriBZqtbAzW4BLVxLqw1haUh9v3NjCO1CKSiiO+rC+bje9cQRD9LFNy/X1jMdTsvDcWQ66+
6t5UsAz0L8KOzcdElZZdvM5+cVpzLIM4Spxz9F6R3UCKAv5w72IQb5uS+D1wisQPux3CIkvAcwms
etsl749MqLJu33eggXI6FDsPc/48eKx1dlIkK5mldoVAz2vkqmaeypLkxqygh2XshI3BYEwo7azp
J8fw5gP6Kupio6P2qSDg9PW6MQCqdr4eMU4VqPMdT5HUGNw3kBrKwOp/thFJJMFd7vvqagtW9HT8
Kj0crVUzkU1mfmGmDUzKVzG1odCTP4VgqnT3E+nfoD+BQExRYpFNvrOPZKZXejssJX8uFAdWyGE2
C6YtRu2T8iImepr5sdYiAyRGtBJqC2y0r8PCde+n/O6hO+nheHUTLYqA/Nibvn2i5CCLyZDYUuGg
pPMIjMA+m5khBDq2bSA/BtLSsiRDBBzEK0UapolLHwzRWndqS+eenO/dC3IrfAYI3CSz/6n+m0Xw
5i7r79r2yImI/k91YtZ7erFt83uBpDsVA2UDdNAzrrjTysWjHFDWjvXj2WAjnAl1lAPL3D0nlKAG
ozAZWVMgAcGvswLqCL7UTqpYoKoQxc7x6H/8up4Xq/OqguvbE6HtKB+eNbJtth4qLfrgKjXiVKT8
4ysg2GCTSX0a3xxunF4M0zx3LUjeusTqPQ1eX2WR+fczQHqhkqKADOIRd36iMalrMYAdcVJzpK1P
O6fG4SOhXNB5Z9pBXwgBw3SHJOgU57ieaLBWa/QQWCE9i15xJFJXEfpXJym3KJPysdet9pi6PXQX
zDLl61OPD67iNFqWhk7ozUFeK6yLGhb+ydkSHP7X+oZ+Xw0pmcgr19ukrE3v1boFET3NChpGi+22
vdnffYjrmN3HtTQm0N4pcWBPX76ObSlZOvrELH35b4jog5941S51lF0lPeaZUJaiMMQbv9O7domV
Aoec4yJnQ2RvBtc+I1k8VI9FI/2DCv4SbJv+Hc79O6lOVU5p7jV/oMNzZgA/N9YAbfvt65z/J74i
fNkwl/zCP8r6c7zXRn9rIdisRvF0urJbQxxdnhX9dnePOmrXw/jA/NE2IdFzGTPu/P3zvrEnSGca
jRe5nHFVIJwD54ECDhgx9TnhT2SFgnrIpTIeyFjoj/c2UJbHGxfEHOPP1h5st2p0jznEysYKoqtm
uhGwipC7/rdT+w+42vr6rjm2rZCDa0slPGmgFvoLVSlAxpQReC6Vbxegv1ZW6tfntYpNaWht8eNQ
LEL06rGSCFF8UCySntMYooj/xfEl4NNTSdEaC4VPIBB+ix8/VD18Mx4raZ9VHOE+93fCCI2FUXVC
e29YBTKT14Xm+c2O8WAm1NkYnla4KZ3i4BhSsX++sRFs4OIHNV1TdsSM1XE9kyYWGYBgjyjhwoKZ
r9Ztr9J4tMhDgbq5GzOHPm+pW3bs7i9vG/4rg97xX1IMkbysIhXsjnRJIT+x8XP/Cp3sIvWx+tvI
anGEIU1P7tCoQwyVwz4JFSGAbhKA7/CUV2lq+o/HzT55aDJgeWyCRvUirXbMo/10ETclcCqKp3z7
0mbQ9VpSPaOio9TNOifUZpat3JBGX9K97Ksi4h3YXXofLNIutS01NdU9xRJUQmVG+Tb+Y08DJkZ8
ttZC9WmJ6L5gNA8snHWP/meujlHBVwBBA3iHNx3NkqbcnZiPxG9f7ltKU5VZPjuyZQ86vW74xR1Y
nRbcXzpJz/UAawwU5oSpxBXEjTGlCK0pC6HLOakLQfcxM9TJicGha/+A6JiYV1i5upev/9xvU3GC
Ca2U6d85kp7U7onTPFWgNvFi+TldXBRHSYbnR/VtC53UTAU27MQ0dDukLCc9iG+htyLazeTWjehp
JZmVY459azP+5M/89YrBsclwe5KOXp7MvzkH8bxJYjwrbVYhAYDnrqZPsoo3C3O5xHRDQNr8FnEq
4ce8Q9uaWYI82zQMv4hN4sRkPZmVY5geX3wBaEK5YRuxOUOMEJjCLw//jtn20J29/t5eHfI0Sujf
4vdV+GNdadPYRc0LeTeAhd/0HJr7efYIqG2tMoHxQB8YG7YvWHCXEu0LLo1t9K+hXL1tFhQGF2uC
zpQFcHsUqMZk9yaI+hmjM6IQ1XT6dDxuSRxJsNPwiGNK0p78A29uqNrdNpdjbpnxNGCInAQStpQ7
35mAcfc/2LhBYoVqfujPB3TAh3R7d5BE0EITDIYkhNTXMDoxoTcb1rp0wB7+CST8Koq1Sl4gNW1K
7Xnz9fhWb2Z66mjz0xCbXOgp+Kvm2wkowrp2yd8yz4aiOaWq8A7qsqXbn7BFhfHB1qRQNPsQkXs4
tW3AOtmNQE7onkTeMMxl9+5LTuN9rsqpnSvCUiu99QOVQWnhfI26CIVUkel7B1vBLsh1R7j5vvC/
N0IkarasgIPTBFvzbojJXpHjqn5P5ASVdJgaAeQpFsEVUWL45bGGsFHmpGO+Y1MqaEHW88d1XZEZ
IqOwRn7OF03mT6vbmIBE6eRSLETOSNg7I2TH6DUNwbiWns2aNomNFvLiCtW0CzK4Vepl6bjEI5pm
ALaCGTwPauza/3+u7uMsFGf92+dkJElcOhPZCO1wDAYeFlUU613V7CWrRT/bmRbSZMsqaEqFVgg5
qaDV6gRUaUa6YUgPTC0xpIYpfQ1L7nF6aFOtSU2YGx3uMldAJhks0dBSl1NIHVoNYWykjY0SEek4
2uNhSE2z4ReNwezYWh9GNIuSC3CPwXdxsQhk32C3gqw43yXPH7QW/0x6tKlYdBswu2gf6aSTdkrm
UYkoV0bRHBeu3FAgN9plWvk/wbz+Fq7Q/MzlOdNzl5odHnaLaXWlNI2nbuVLe7LVdIRvyKI3r+MK
q/oOk5UVvYNhB5Bv2FJezeIjqh7Lny0bZ1yEzLaGHepqdQeKWrdXyVcd/E6q4VAbe/jetlOInt9p
dolZLlnj1priA9QYyFMyEVst+RF6ieoAo/wS7To4Oudc0Z8qfwUJUOhUorkqhw8nu0zY+Ax2FUnj
m9MbwKlshgEjMHe1EDOJP9Z7uVplD05sXZ6p3v/Se67X9f7pf4Uq5lrrp8EqG/McFokno8ZsDv+8
OMRaqvCWc7Um6OkMLRV018iOkYHwSQl9p/5E42C/x2uyRDz86rKhbVN5KKTjE08bV7uj0xK4hM6v
D1Ei0b877HGB7jYgZjpW3NIN826yHckPGaFKfTKNZvCoE/ZTNmbze0s5mlL1/7aDXYOE9HQFo9+i
7mBbdlYMUXzYRswzXlY8yjY3FUm64CYVD1UDoq1cYLCCmUs07qKsq/p2WrIqDPooygLCWX1S2ZBF
UYhLZl0Tx/puFrS5lWbadOS0mqxPRktIZQ8QQj/6VsKes4b1Qnxacm0fXu3NznhJ9wnxlaCzOibZ
j14exFdkuhveJU0aG0+0OnmyIGZDzMJacCt+0pJHZlNta1zxzZ+lrvtiIvCkAw+rgjPMbTHun463
1GvkMqW3lwQGlHxUNKUg/T0GNf0/tSHFuIJAmY7oRUt4+ttcMYGfxvaAgJCxSDhJen0lyfEIiG+i
NSN7A3hwrugilYEZRC5EUc4KlbrEO0PcKE5WWbafg52chK6VcPMiKC0n8dqHJA6yCu1LDDNZDFVG
LQlk/E3q2UMormN65DyB+lYyjwGEZMXUynuIZz7UKRFwkgFYAM+yR00LxI5RgHzPaC2HSrKaVmB3
nTmLWLMt7ni+y1Ow5owpPwQMnENkHUp+vpYkIj73yOaYWs1EFQ/aj4JFqGY0j2rAK+H6HQg4Ig8Y
V35vC1VW62VUq36Y3GxsK+xPqm8CH4PSMUqIC4xI0cZr3OjlV/jfa1zcnDD9zyU0x8VecBXeLvWP
s6Yq7Wasr5KxbDRpP02WSni4bYnjS+MJdhnUoes2881Jujn01IW6AkCT3sA9h3VPszPGFgwfHaqO
jOUBv6waIpeP9z+RksAZcx1iE1vV7hcHwQsuiMlz3Vp2jvR5TWO4EO0/rQm9I2oW49tfEmZVH+vH
npQFFaXlwhtZ4EFasD6qhrPoOgvMjihdR7wRusmhkuYx7qOCQ65ZPw0a+MrQQndP33f/nZQyoVp4
xriPgEhqGhXvVciINaG9F8LzNYedtg4Wh60zuv8MQ0yecWobxqij6JgYzE1/3ELX8xKSB0+4Ti+u
1uqoP8tlNhVFkHsWHU9bRCi8WLlJXsvu9auJuyRuLcbvCbOSxkhalHUUp+G1lcGHPXtAnczND21G
/gmKhHxZN+X5j2p9bjpSQjzObo+T+hfGC4XeHrsRLMqkiq1zU/XliWxiY0A9sDEBsfN8eWd15auC
DWbiLSHGgIVhQehXhP+gGQXX2ATvZQy6fG9ftD0YBieI6D19pMQy4eOXU2EBrFOGhssZQqw1+bDx
kraZzL7sc3zQ5uhxeC85AcJ1+sS/ezYMUa2aHhGw9rJsEsrnCgfGxxGwJ/czLCpiMGEZsEzzCOtJ
rMWEdOLv1yST4707ToUAtZ3Yq2U4GLIftnGG5HYeH1l9ioY4+h+zoaT5+t9vhCRyYQJh7r3Yg/Gi
7RjgKtUHiACMaLSoAitgjussj/38Z82HQJbC+2bfVBrDiOmMIbET3TL//rZltuP2It/EvQ4NOq2j
LMALOy39lWORyq4BjPUV2kMcLz1PLKSStv40hlNR2Gl6V+HtQqef2Xqc1faTT4bljYpMGsW/06Zu
nGBdzRuLr7nBP+NkUNlZMGJoF7/3pkURy/n4XXuCZc+tAXRAQX4q+IXuyVFtbip5Uo7ZMZ1Rf+2r
9OgWh+E+8nWAYtBKxlzJUXXTxomNJyqGbHrCiIJKbxeAaLhP2mpLv9EFIf1kq+HbroJdsiyFMcip
paZVSdc9AofatlAao+5zT3VENWKlOX27KwzrsKor7AjsVzTcFKMyG+XX3S1S5/FaP4XsTm1bNqpE
3B4C1+ZTPHugcT0G4j3JlaNf96pNLKmZGp9hGmaEVCVHXfBK1fan2tMoEHuJSTox5yRlmta6aH/L
PH58YpYHF7h6iou5zJ6C6Am0CvI9VafpFh5O1mHU69IsWNrj/9w8eQltz5dbsV9nSo/YO++wUmQd
vCCeHVn0Efg0HRA6QWXo1hmJf6H3gLn3+NLR8WVzzhpo7zIMHuefrfQ+xutSMxL+JmE1Qs4/Lybn
Z8juePLSnOsRCNvKzbPN4rpaxNZowKm87nNcb6AiQ6Ahi0s5d3bMMU/UArMTxJ82uZogAyqu/YJB
vT5FBOs4yAorO8z3XjiX/gfA4gsk9gwAtn4kfwR0VJOgpBCvNAsynC1NlZu05PeODP3xM7YvwoFl
HgglQB3w5pmLBZd/PKJ1szJCwnIZZRtiq2t/CVCOS1hui8C/SZurEO3KDqMRdmLRaBVwMvAHPLfT
4oVoUIlQKrFJoeJyboTt58I+0DH0LenBbRPYqiA5W9dXXBk2O0eZw2gSpjhkVqJhXuNXQwsyU7Fw
bgHLpfi6YxyJDXdiZcPUvf1oxQh9uw38Q2gYk1x4oqSDheTeipVOWB98RTgSxrSEt3AHuawZwjZl
ygo+EJfJxm+zFBf2WPtx4u9+iEuVHh7aHkFwa6GoUMXVMTlflzfIfqe145ebEWteSfenauZAFoZX
B+ars1kLPdcOQpUqiaUkLqo2Ma9GVhNBu/CSKRrMVK0XETilIQd8NUBEYg679q1rCLO0gNUm0ujl
M2Ks0J4Yer2F9Z16gE1p8Fk7tGOv55rSQbfeq1ijncntS2b/5iWZiQasB3dyyailnPu5SzqJOK02
rPZeeWc2Xzo785S0W1CX7tTpsIhlOI2OzOJqigGseb89HAOQhjy1Orl4T8d8QRA+ccMY0xFRS6r5
BaVxaleU37VGkRNSs+bnbdoPq4E6jkKO7Vi/6VwiaQ35oZnyKGMIJRucAE5BM/UIEUVDLT0M3ad1
uVUEwSzGya66LmbbRjfYAP1BuvXhm3RMhJiTahBmrlEhUWcJUHfucSxlOgRWX54gEC4BHjyQ5i2T
pFIrpLz9wvwaC8eJ6CN0QQtvzihOtrhW08cy6lFuXqQaaEHyJrSkXy7LPeOFy+qy7A2g2Gloa3Oc
KwBaNB/457v9oMeWy5muKIrxZ/Z4HWF9gXYwT4668cNJ8dPZQUgnWcnFIcOz1HkQuZ+Dnnzg9p79
N0bXu4+4kVgb7vO3JlsNi56Mc4tQSdJ7yx1pTE6dbKeu2aUnSv51QFkdMI8ZKHLAk4rn6pDSd7Jn
wArvF6niMJWplRy9/Tf/Ea9v0x3YaSym971vsQmu5KcRGoOuuReqESr41v0ElP86Ev3Sg8fDew/M
d8NI9A+53yOnfFdlm7DhRPZ7IsXAVd1yOP0YBJ4Ae202gmanrdq9ARzeg/ffYWesIQM6o/SwyDo+
s5DVhhAIwZaGRPSNzqw/kWYUXblbJYO7AIWak8hTkvzCGaG/l9TGXikc+UjuMNoojKJj+QhpaQSi
W5trUSm40UfI/SovMRR8CUwCbFFDJ92TPasvrjGzTBsJOL4xiJuhhMcEzZhmAUiqx5Ns5BqK1qPe
1S2v/bDB9idXN680dkv5bcJXW1eItzjUuWuVVLQPKRe/mnotJFjc7Ja1Tw5+hv2+eyNwSHNfTxUo
WaK1tfxeVqVgLPbJhA6+rdWYD1J3w0sl2kt9LDxUnR6iyvR+igurBt+vqgvXwMnazLbOrqquYkn2
TVPRXhTQZsl+BK31smICto0juh+lhfafQQcyKjBWY5XBPpRZBK/jcnkjCw9JdWbTmO1Li4+okPzw
fQqdaHSH2kKZF4Hwh2s/AC3iBFq+3Rz/vUvM+Yowh1QhPXlFJcHgC9e6Glkp21jUmSIxvzd4iFMA
wwH3YUWk2pIMNLUABPlWpFEWl/wVCvLXsv6RFEMkBeAPhR3G7rrjhP+yhlbQyZs1pP677EvRvbBW
6LxHSUQvez2CDJasi5ZGH9IZna3d0WkeqBGT0K97ICbRUTS1wNLx71vX0Q0XDokEpXefJMUvGqSq
Fjs1H4RZM6P918fSirmsbI1zZ+mIeqvc6hqAk+nz3Sgl+yamnI/ANnJVrP6IGbjQEz2D9vUiyVnY
YOxnkWvU9vhF/uvIRk14a5xreMeV/sdtATJ19zg4z653Uh9IPsTloO3tNfWhZBpPMncx+1EkXib8
uGg+sePCzhgLZLiP5d/eLPp7NnjtR9zajOYB4MwbQawZSyqFkDDSriQow36NtDxTrM71dw/FvtPe
Yta9V5+Dc6pygMs4aNSbxKxPlAZNHm0pvLLmc2lX7zkREqap2mLqlq/4WjEXV7gEwexxMAeROStY
1mMkdTa7Z3jx3upngJZ6+t/JkTE5lgSxqD4OZkEHUwnUAQQnzRplzlSVhYp3xHRfV7dauiv6aOyI
Eu2JmxdrJ+UFEeOgJakyoeUgfRRWjLc7vrYUmbOFOb4l3ieOGPWijBWMlLuHklF/k66ifiQZs5U2
r6F4qefRyDmTflgMn6XLJxjGvrtx+ONrWb7mjX96TethSeFrnxp9BfzK+K0d6hgPlbGXgTWE/MTA
eMEwSmH/g+cXdmr1qNALm3LtygYtoaJImxQum9+wEexe7YeMRP19zWqc0Kk5xH44bjWRnHc5tMCm
uTMCpQYfaxcx/OnKj5ERZk4NCGE4Txt4Zz7KVeXSfvRI3YS/8cPp90PUUL0g8qG3qaFXAoP+dTbY
EuOF9PC5mD6aaUPHDCj2lxYEbwTBPz7ywHXraGhvZL0aNwCXRhtDBsS4sFREAGhRmP4G7QJJ7ePR
5CxGZvouobCGmLvURPcnxlJM340iW4ytIv3ofPzX6Ii2I0UTcSKeL3PoMPQ8vMcwxOVtDXx4N06W
SuuhmVKoDMrN5dM09PxrMb/KIJeLImjNMgbR/oujVERfd2cuY/uMbG0YnFA0Itmpao5sOD32b0Nd
iGjosaA3S4tOEfUcTzLeseMtX24QP3oLLpiuyZrW2+4XHgnYT7HkPg0O7yWGeNY+PKuUc6oJcyEw
ycepEtT4zjA15izh53edvPWZheDoCiSwGlm553uTC5sca181AVKqUORLR26utjjI2lKtQ27/4E4C
QeqaJdAWWsTStw2f5ctFrYmImEKSoO1FVbTRbKyL79IWs6FcgNyrwOEo7XUUenv83mGW9PZCZAd6
eHHz48NkjkJom3nLUDx4URZw5LyvAFXaGyJXiZUl78rm7LPhCS72J/KRI7Ze6ela++fp/Fnax6Su
EAPRaP80pzVhAHScoXbsLKbCIFv0pgbKt6OwgU5kwBI1FFiwRaXra+DJlhWPCZwSzcSPCkF0s28i
eSCCFEqm/WGSoxY4I3kS2oLBNp0+IizjzX2MuiU5hhXRfqGDiXS0Ph3zbQJnIeEd/zfVxTcqvxMs
lJpiECp3VSFg3AsTXy8mwG/PPrlEV1WminscZ0ESP58Gswf8KdQtAestybT+vVcfwgGmZlvLXMcO
kM55V6uS38lm0mrFcJgR44w3LNBSbN4Ry6mJ7XqTaupaD+d7rmWskGWwbLyLV8M8HG3F/ec10vM9
QEbo/ynZ4dweHOVspAPz6eHfpNg7ieZSksEv8QtoqLh6txNcXBdRWyBSWRAeZLkAxCtDUlJnNhtg
uwvjk5xq/UWP6C3VEa6FiyiU3UWIHapC7y0H6QCKjfX8wMpBbC3D1L+DChTpX+LupwxkxG30KI+l
tnP8pZKqbGMn00vGjsRTsfHoMAP72UalxK0rLM6AwxbsV7GbxE6yBlXXt2s1wHMiIPvSJd9gc6LG
E24Ysu8gw/orzg4j+iIf9Q1xJLuOjovk3WvA0TN+8f+tHkZdd1q5yPWJ8MP1Z69psk8VO/zHjCKU
bPoeCXOhnL6IFXHVIxQEzvO2yAg0pCKHnsknpVB1ZtghS0NphCrJbEfr7uT2f6C/AHRr7UkxwzIU
LXuqSGaGfyGeKIWrEaW7ubNjhZAjZ4FrZDeZpmU7YuiOieIzWTP/a6m9lxYk7awttgxkD6qbCf8v
W/aq5JIHX86LHdBlj7rrrj5QfJEw2M5Y3AlDi2Z7oy+lS9dRgxy9RiHMVgZzdBVoFkNa2aybVdSl
uJv6TZ17YfM+5z3fXu+XLSsCUrlMLdIGvAEoN34bwjg527wPqGmFd/yzzSt6KpTHwnuBKnZ2KQwM
idYZMzIlDWzMr/RiVCGJQJHJJhaLRai95aHX7jxsjZJSyahWBzzlMfsHujP5/u2DQJeMcc1jsEwb
aBezC5gXxotJdpBhkaiosmaJfTMtHp2HE/1nggxQJ9aLHA5W0KE9EVoqu1R/u1Ugz7kZ6FNo8U28
AE5yLmgtpAURhPt1x0+b3pEXzZqO9n3TwtGVnx7LPT/fA9rA5h1v9rAiAwumVDBa3vwKmaJYYTXt
rzUiWpsOmSabHE4+APUF43LLTT5Kd7MQXO24DXMi4IVRKs6VT1alcPimZU582JTJ0bu5cA8IMYmQ
ZO2g8o5JV49KRz7Q6fUsuDlLZdHrGQBrBvqmpDDvTphpbHIxLwhgNiS0Egf2UPgbTfqGiu42mef+
iyPq+Z5iQBMAnKJ4U2nIR2AR2/S0bwz8+8a9sxWnwHiXBdVkJmbCCjdVVKNTlqwujldzZKQecY2C
2e0ZR4Njd7hYISzcmaQiTuIIAReRlJ2vVybNNLV+VaS2ExG6zrPMrjSy3Fz9E0SgddcKL38HnMo9
XrRhZSnl9swbEN84kDmM/BlJC7rGm6y+nCJYyPpDrKRx7BfZ+BiexxEVsiWxS5nnj5nbfJZon58Z
khX0Hcq0YvwZ6wAiRs4wcwJfdQhkoE+S9+Iz4wp1n/QsvxawOH9g9GgEGAbFZEktQgR4IkWEMdRb
aDqpMqv6MwWxLdS3TPlYrpy1Gks720N1ofOWeUv5l6+Vn+vrkqXRoyGgNVsdTSiBmtuDbjvkUspJ
9nGG773etHNTi9sxnnTHYQBPQBo9C28ephJCpu5bFaBZ2uIX/x+L9xSliHnL/I70keoO5kJugSbR
tguHcA0zggCmq4I7or4W71SaCGhQCk4ULt4hzyssPZV6KQrjzYkJiG4eWMzvSvGwOe/BShWGRDli
3q2WSVIMJ9Lw15s0ym90q5+P+Cdru50vUfWgvswi04DA9U1LfCLlUvWhSYmtGscnwCaW2NdRynLi
KDjcrQcuou8tVOwgack9ItwZQhk6M5CmG0dsxaI8VVLU33uRLQR1q5BL3zD4yBpD0CTzumqwBRQu
aeRFBTrmuBLGn9xsnKFiWTODMC7pZ851HVsAtuZmzt9yg9GkJfqzOR9hdxiTPMyfubVOi8qruCPu
dLKC72SY729Sg0ysUGk+lY2uaNxzgInfIgQ6guPKGpyRm9IE6478QVJWZD9uC9YFYYEAC271HFJT
vsvnzC48uxaUrYXBI/MYd4EwLPK7jpDCez0cKileps/lI64Y4IaquJgor0LICZTZzpx3Rbsm2bVm
tYB7K2msAZCDxFYLY72t5QugdJdWKd/3cE2GpqsPrJq2vUE8AOIahLc+x0weBpvdqK574kGicZx8
SyZPiB21IShQ4JKz8X0jFCoSMcVrD8YvGkmS7qR26Co8ZqiTWOolCCWG9Kt/NXNgPMBUZTehBB6M
btiMbnqCkqcoMcqSkRewOvkG7/tXJ99BLmZ+IrFNVm34p5LZ49olrm94CrHQ2nzC19552531UJ4u
nVvX/YNQ8v66XlJ02ojYFoEnyMEp6yzWXMIPaOGiqfXhsd2Iqdc8OovENMQoZIWUHA0grn6/k9QO
zLEljH07wtWvSxrBErSYVrzdNFaKBokKLdNWYEY3mwJhIS3l7nHSz21ffBeVzGhOPkQIwp/aVyUo
RKbSCKFO8WIiRKvIDDK0Tixy4iH9v4JDDCqMQ7WRTtlTINKxrMpFDkxbZNpXs/6qe5kR3eC8YIaK
RTz9rXPaQ/g2U1AWASU5fkHqhC1Ewc8bD8Cb6XrDiV67XUCKGJ1hl680A9qWuk3I8lO3qRRtqtEl
46MeItDexSzxl3f+O2IpA1E8leFhB5nGbsjlG1DiTFLVBzLahpkYyCbggAtKx3e96bZ/nrVQA61W
78U+Lf28YHf2rXNVKpJVez7LUDIAR9S/zKm/LtcWcFtu4AVg/WLOB3VeU5pr/WQeSDpU3MotoIGp
1JVj2Q5eKRP2YSmt7iSNLIQd1czT//3cqOzhKJImkPSUP4uBASEct1Mbyhanm/t6Bfdz+BEUOH64
6CraSmudBMLt2d5i/pnuDJ1ieKK0v2W/3B/hBfZUviNxiZL+LezBFfThu7Z/ca7xMXH/1FLP6FLu
gUOKegsMO+Fq8CqJbVY4Gpa/mXkq4YAswTHxcvda2mlnDTNrcnOlIwnd1CUR+U3Q8Isg0JumuhZv
KBcdjiQYIUaazMyJGghGvaFb1bEj+DJ6iFoLf50DIbWEQI/6vHV6toqHL9+K336ZhT7dcu2W4/8v
zdARsZspi0I0kX/M5oKDaMXh3iSXpSoGYbajV5H9lDUdowAvCfWPDior9dNU/eOjnV/gKwSHJRk3
R9pIBA5FiiDqOiDUPIvfp5S19P1+xAXNSq8guacNEo23rXrf6HBCqtxH0ZEMZhAlUr2x44mKNOIL
B0DIG3xS45pTQW3axjih7N8eHSjfyle/xXkGQQ5KPfw+3TMOWyTunMYeWBVDfI79n7uh1iXxdQIc
AOf/YDyOi5+KNzM7ZH8GN02Sq8M2KI49K3566SRj/SyPXRluvTaP6Qf773yO5P9J0A4FVWxFdysd
MRb6dNWr0PjsQ42dS+R076LQY5x1GtQXb7jX8OIAgomvTV/s654DV7QZVQXuE3eKVdrDfw9/kX5A
tttnVYK33I2kStb1k7Y/9d15YlBuRnYQ3t3YSqteKzsKrci9YOm9kzq3HX9QK754K61fY0uAZqhR
mCOOO/hkhCpE9sC05HrIfbrTue3ET0jKL0WhpA7MDEa+1YFLA0Dla/LSEdcaw3xxAgB+HtJEAcbB
L9temIgeM5vrK1XUPWPEFT3swRiDIkghzqehvKcBtJ0c3HCJFNK5XV+1xuw99ian3ZtsexXXOsfv
q9daAbRON9sLRyiWtJxjJmpyggzvuxPFDUAS4GPCIN73/p/ShENaFlyqP/SslnhrBrVYA0IKkl+F
RGQSqcyyG4U3RzV5jnp59dt/4iKfEXex+/x4zlPuN5UbYQQVD3xwg3G30AqV6qG5GW1ratkc4VQ8
/dfPmVCbQha5LUz72tVURuvvCj9bUiEDH8R6VIpOnn4LCfRO742Udgoz6bWSr/LcRvmIJzvcnZJf
c1jVsUS4zmXSiNj4Q+vrxEI5aqw4HFpapUKFTeNe2Ajkf4u0L/HX4b2lD2iujdUjDjIlT2P9NYv/
b1kcHCstyFtZra3jByRQ23l1aF5ZI1U7WZtkQNO/zCggnZ1SJfNrZQWbGFCB/1xtqRQWDL43gkOg
RJ/qLi29WOghcO51eqgLyrTy1/8kQzcnjAKsF5qkF+s5nn9TPgjQ9DYg1MVbRcI7wv+ru27ls393
h1+yhjIPd+IBXZcCbFLZMBN4FpqQFZyzXTINVMSRhTLU/QoX8bpID6ronXcmgxZJQCn/1CFxaE6J
Itzd9/wIWYvwbiB1HisgxWn7XsLLnRu5iqDZMEat6Rv6VQ6fBWT0kikgPN/PDXdgDI3XCVYmCjV/
5JemAmY/e/7P9+h9s9PIS208PYPxFIJnSuiJumT746UlPRYZmm8XqsMG52YzfWRDVnlPEPGhhM07
7arQZiMmL34D91RyhQpGyvtMFoY6R28HdpQRVa5LiUFsLnj6E6y6ifYZty231/pXxzz1D6KOdu12
LKXm6gzzyTxQx00g3yNgKRx3GXR9Lg6DfJ7MEWmXQS+oNrBuwJR3Bq2xVvs0x6OzHvlKmCdFJSf8
GDyqzUglEkxz1QReUMrIsJEkzD9NB0BdNVWGzFkVcbz/2aTzky6KtDP3GHea4XJIV8+h3WnRjzzx
oJ1i7N2CweqWrev1q9vTadnb5b5ViykcnFO8Fkti/6sF58Iy1ggY6iqoclX/FpBxhktKZKyYg2qd
4GhURIJnKooEO6t8VP8JwlOwYwRCs7nHZnRuPecSECjvbMQ1wubVzBSoJkcVkikfua4f9GMJIeC5
cNdTNXXzKvgU7O8PuUXq/nbWyI/gXn+V49RZaiFuUCyfr8qlvBMlBlNkDJXILzKSbOcMAPNN+Sn5
4ifYqbtq9dqV/ACEwwiQd4iY6+CqGAFQ7o+d/kKeg+FGn/TZt7enGgDV0+JdEBbsOtP3Tm0SQkSA
tSzW4YnB3li4/MV7yiVpK5mtsZnLRhOg6hTj0ChdAEl6aez1rmcwbEBtg207S4dcrIsvXieKzh8X
Qw07oUzrpSGMsDw7boNww1OvT/KJW3ZSAi5y6Os6NB1xpzS4cKlh5SDh8yRzQMrbUPm/O8NHqvhJ
d8rcq1Jxz30a8bMIHwJJeckP1DKS+LNg2UVXxsg/5i8RGIuVZQtE6ZrI9+yEbGRqbtkSClC7N+SP
9J1Nw26z41FNj4VeRsqYhHrEPoPD4dIxFbwFzr/fcIEHc09mTZ03paWag93RaCGvQt/GJa51UFqH
PLSkrFTFJzWN5YBgu++7chGCyeZmgVSyp2vC9pLYMQbz7D617Br9ZZIFdBMbrI7td7y952/smYGl
D7aELAgOAURqIcLck3C9iev6OdJaalf9QBfKYbdvPUDK+EM33nhqnJW9/1gVWvZlGDa4wWKUUuhr
h1zUMwgPNVkSX3p8lzzn7VYu9JmsyhlMdFjXJyil99eW0gw2fto5t7gy+LCnq7HjaVRhrAoM1jQk
iiqkg8uBtRDztgw3xrHhzTPE085Vsyr9HwSHnMIFO0hIW2GWPQWzadF9XnwEsCIzaYUBlHCOC9qn
ACqtuv9v0XRmhs0Z7aHSdOAGbBrarAWG3vvPkqq+FPIy0JV8W2vGMISX+J85d+OKZlgf12zpfy+y
H7UUANdYlm5pUr1v/nap4Q64dXOZmCK6AGG70QISsV6RrOLOjVfI5F5lbEcJaA7lokFdpTSzWpwA
OzGh5F6Fjlsd2Da1+10AyDjeU4i7W4bO73jr0DfHIdkuhogF/wJa82SwJqzrDVkYGnhh9IKK032I
DSEmO5CTwkEJUnFxneokIWPkk6xm1NnnPc9vh/rfLTp5zi71kgU28EhtFuT5Kx8I6gAdCLBFlpMP
+ajxL3aASQLuJHOa+BJAu61pJBFztXpnYi4T3we34hJ8WuhlUOcMl1ZsO6RBjX5CDrKsmE8PSYIn
aRQ4rDHmHPurwA2RdTJmb/5AxEh+edGjcZUgBTC7pYm4kgcIRsget4tRbFEjdi2gu03FlHaSiTTM
S7v5GErqVmyCBC/gFDrSPvh2JOE87RObia1AHlCJFyUYr+qyGzZUWDUwh7fI/LkDyhBsDkf1RjZC
qvV0ldCbSh4/RNAxJaSXiAEkzn/HJPNLqFxVHN15V6an9Z0F3LB7U9sheUI3ENEEzNnH8wkm+Fmn
C262GCHnUajC6E2T1lk0aadm/4a9oJkPaRFE1r+QjnTfOJ/SSVfgeTcToL5M2W59BfPSEk2YzuKo
qMJ4yjSrahVWZp7kmaTtRz4TaZBS4Jx8F0E6DYHEvvYicf30zlp4j5tmLmdHsJuDkYRkV40HRBVG
DNRGiv5egFrrOmxfZFCKs5j6OknzHEKAhGzn5xRD9XRXjcShG6WztVLVO/bZPAAzhCbjrb+XLs9F
kcbJWDkY34ILITBrS9+pmVIW10g5QBIFz+u/2h5OaiaMHMet8fhjkrXsYecAScS2QfjUAgcCV7vU
0FxaCQU7hr+kl64Y3YSGcqLRxiy+LDE7P3u9lyb7IRETIzGPlDk52Wcpi2jLIupGEw9RYR0bp80N
rtD4ciGMJv8ZbJGpRtvYRhJuB6h/iSY21FCyAri+JpSXJk+TQgmTuH2gV9akG4ZB8r97pjSWh6Wp
gUNB6F3Kk73ksA1j4tSaPiKnuJqjTalO6t3XRYfooBYtqzjAmFZxrLWD+hwktkmyxXZMefBMD7uG
Wplhoy4orFf618VaxLdRslWML6mP3aOCl6wpop/+puRaRtvpvqwGyp7B4yzc5Wl/SxM+eaLJoyL1
Uau+2eJPawc3EsvG8PuiV08+Icr6jdskyF6mHgsUhaSFvrKkwrrAyj/Xmejr/Ks6ygsw3S5yXqRV
rQm3IYtv0v5cuy3P5lLNyXlaXRVlThzJrfN1sM+w84Q8izzxNPCPi4WyoplhQGvzVl9akzPH/rWN
wTQgoR5grWAYaJwizl4jMBfh+JyLxPrdpqQHKp2J59wGE4WVIC+isbsHFgxEJdw4TqzuRWkKEC1k
Qw0VNlOQzqREotlnEISoScKnTSTkNv6jbHtwb8SlJSxsFG3ddrW42yN/9qUVXovRhRtLH6HcGEUk
hBH39ioNu7ABdbrrx9PgjG/xfUxh8GbfaoWftNDWUZbQNbluX6MWrMOsfKrmy/XVvwH3Z2KegnXh
poPjHGY60gKpY65tfAcQI3rLTR317Z69QsYJX1unQOKUW0J1O1Y8PLDvR5CRFOi6LKcQrLH8Lo73
YeDQcp9TDX81VuNZ+x99qVup/lDBnnfBdcGqr6nrRivcoevNSUzl+KI9CwxDb9MD7vKynosKkA+a
/6kCziaTM2p3+o92OgInMK20fz8sL4JQ9AGmYy+Z51ua2k2b2aMsli8Jre+ug89hks9Ecb/d+PiA
0XzySOYtMFvfZPpbzpLt4c1oKna7Ep58gGQFidCW3IBaD43pgbDwxuvFQC2Y2GcTZv5uw6XxQ8Oy
2zrk2h1Ezkv0Oj7cYoyyMcLCcasrH5uc9dZRYGhl0IG6e5Ym+bFIkPvBh8QhwuSn6d6eeuHCzF78
o5/JbncOa8VelIhJGC78SHVJYyZiOkM1C2P1K5DUcTvHTJtiuQyWEOQXkLiRilFdNukh5QimB+wW
qgCNLKirGETY8XM5eQ/5J7Mh3facbO3j0LTKnUWxm9P3GAJg8v+xKZ2NbpJH6vgfdj2YKqg8bha5
lTYdQoY2t2fpuGtGXBoPfpEkWT/aZuBv7u8jFsC2eFXFZwktb0GFI5bFlaOxaIrLMnvUJNmaxI6D
VzFZmMw2xF4kdXAKbRBKU+/nNvEurMJfwLCyV78Vrlbj/hINVlkM55AyZebRpYeJynjUvR9bE3RR
2U9yI1HfDaxghY7mtIj3Khpw7d6gkIU4RCUjKsHstDBcZkmtPO3jy7nfRIP3b5tKsCctSgTvnVEi
Ppw0z7lnHidD4aoGhmlrV+qXey2tj52tiw3OXP7mloqgUQcuFn3HGdJ1rhSPghOZxFW1u2/sG0zR
v/Em4zlvabBwcUtR63dJW9zLaRyZ5f4yaca+EvCvZcYVob0LEAh8WtHi4IgUSseEHJrtUjLZCj5t
xExtVO6E3BmPjLvrWDyGfxFx9h7LT/bP7q7xOPQX5SjZIsAmRmJ12KbSWV9PwMqsgqC6eyiVs9qC
GG3zAZ+kQ1cwC7kgrV2vf43rwk3XqFfdMZBicj1ByZ2FzCfhLGMbbfhV4B+srUFYzws9Uh/zGPCI
9YGagMYcl3+UxSFFn+zeU24shnbAIguKqNcRr7IEGpW/oFw30FwP7k+d14fD3VaQaYg5X2E4R/ga
U+CCfQFTj8AkBOhwvKPHey5zBAML8n3LpMDGL/1dsSQvIN44FSNc3WH11UR3arPX90JQj/F5egpP
gXN2wiOXqgmZyks5K3ERbnLumNPVOibK4KePHLgcY5y0rAtynNnVQCOjTA6Aj1eNW+liJabZG6UF
lHqSEVMAL1J5I0dUF7HJYCzT/Mdn84IR8TVEY++b/DJzFfD+PA+RK/0UEx3sH2zD0++mjaEnySln
bkusILxvIbzh7sK5qloF63Y1NHFSciSXU4cmZ1N7h5Nx+v5+JlxO9fzhbiOoLmccYE4nWEC8lRE4
fS422vPgLTc2pLJwkibJ7Ngb6fAG4RvtNL951F+0ImcwWquCTZg1UR1droqVfqcSdjHg23AsecH+
XrxQJXryG2kJMWUrFWtTUEF4ybjw0e1UXL1WIQ6nDi6JTmuimlcGjdOuoaVk4HRF1bRIC6tci1ob
Z4lpS+otjOtIU6cQjzgUemlqzaPl+AtbHGKkPbiZq56K4z8Eia2IRMhM0nIckjk3enjlRGWpzC7M
tzk+no+siETcHzbDvPGv+4nYudbRwMzA16cJ3eZ/6fAyprn2accJnx8v3h4/tW0DrV/hzkLtcYZm
TCCsdM3pO6mwiDA+TYJprRONYTVgFg+sHOxuVI/rsJrP8cTF17i1xkKMnwXN6XtWVsJbVGRVQjSw
IORlERX+ViSt6lim3D9iLiqC1ahMKQZUusrTX+RVa0XS9TT94vBz5jbM/Oqr7B9VFhnw5AUZJ4dG
ZW5nB1kxR0oVUBzuvpBxNM5qwVzdXkTkRTlLo34D1JNqq6WTgMXBnlXmuEkqgR/6v+MpCySkEsLe
e+SU14/GIkq7EPit5FKczMvc6KqLpUCvc2ut3f7VMTwg953Yek2+Uq/Ed4b8gtQ4qVrce6PzZT2d
Bw+d5GxO3l/10xiZH3d7LzW5lYDg6NFxVicaJAe6AUFJWkujN+a1dJNvPnf94NS6hYSnQbnSiFuA
rtUB1v6jKKXsa/7z4pURQ1B1HlXvjp2LH8SO7i/oPDJUw7HAurAxlJxmlL8Wu+vPPkmZPFiT7jAH
LIsBIN8YThfJ5Ru1W7Rp0sQrahiFYT9sKDNYv5bEs6lLAG8+uvpi2GEVaklxYYmNwIai+tFwi6Dq
fpRbVvJKgAHwWHkt773e0UHKtES0KB28r09rVYMLm0/JWROTWRax6ITUu6DvyMaE49uX2aKKUNgp
VNJ3O+caSgFnOvwn+1zJ6xwni9yUXTe3YT9ET5K5Y9mTj50Q55dfpZJoluKukf3ysbTSDyGDXUus
4rguiV42OrFDB7e4BrCtiFQ0BUza/xjkCcs/HEg/l/gDnT6fJg4Wnvn0EeLk0wUplXrYM99v/AV1
cQPXAYrECtHxD52h0pK+8JGdkI1ami3fBQLyFU456NoIj7Q5h2AooP/tw0EUZpvKF3gPw4Mf3txN
DJd88W2dH+sy8eLRBDQct/kdHd/nTK/SGHd0hElGtMSk4ffYd4Fo165nRTBhcpCGWgdjz1/Tzcuf
NzIypKeO5VRDtEa0Xm7LTsUjGuP0kQWitZnxDd++DSbWvipNHkaTQ8HZnN1vSa1HdFZZRqgpKOG8
CX+49DWeApkKtRv8pYD5tXJovFMrBUzWgBmxR+gkoJCJZB9hN1aHSULK6cdgLNGo2p2saAWvlvyQ
hKgkQN7AeS7N3FZVvfo5qBoemqBAeZ4TLG/+sZIJ7Kki9w29vqdHlrCjebY6VuYdIg3JE6ZyCgFD
RFIGgIZ3AMHENBbN2ph0FvLrONH86FOc1jYY/5pFYAqXNv78izP2R+hfmpn5cTh3aQ1MGMW5ZW64
0uaaNHpxoeFR4OWH6SrpSHHyr7GdUTm+XcQ1fHP66ttoidabh2AOMWWm9KPuRYOPHnxz4t+K/Qjc
rUDb+yloZ3EexBHOM8r5NNG28XZzo2EgP/m9m7JIhsVPtYy7o/MXrX9q98PLZu2NvAKs9OhBepZY
SV4a2giol6e2jCQCzcv+KUrKBM7Wgp/+eO3sIun9FR1ROHs05VFeW5hY0ClqvlPho4+ZmORcVxOH
vtHUl4rSZPAJPh2NK5HHulGbGiKktx1o5tJk/TRPJFagsGRE3jMl5SJOMaIwCKmqAnQ0yKhPMaLd
xzFpLvMRcFRtvWmO3mO53azG6CXPjqyEIJkuzsiHTF9fZ9ZOXLwGZP9ZlDstM3t98aWWqK17tmap
vpSERAx5PuRmjdW88uGCm8EQgtChRTXA2+Bh47mKmSpzKtbwlaLvRzROSmak8koFRJdNGgK9ZQ==
`protect end_protected

