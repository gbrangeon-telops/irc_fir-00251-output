

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hezhI5arYh5Ll2LsYr9SKRVb8M09iAN2m4JSbciXeqmprOA6kAYKyNVYZrZl+7uJ9rCbSy2t8SS7
C18wuehlMQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iG3qoWxeKUs22C9+IygRgNw/Ob9GNJdHtLxrQAtYdMzP86eceFi53EP4Epvud6QFqZ+YCcJAJz6X
BiP6+zFZ6SCjFFuXw9pefFKNSIH8+q7UF5dPb1d06lbHzIZD+3mRDkhnSZjrqT/zLAUZb/IQ1Lbm
Z5oVMb2d2CoW5etMngE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lCcH3M3hshWBn3vT8V7Ds2ckpLb00IXg/NREvwDTgQ0x1n/TYrAfJvH7lJwH3QNYGbvde2S4oTtp
dxVz5eb3NKybz4CG1wYBC2N8cyfQblBGlezgCm3PFTB/fb7+0CJP6o+JNkedc2s49uA9zPZB2axM
QOZ+WiL1UDOqHRt1CYUPiwYxRC9z2R+kY3HwbNnbrtScHXOfjyqwc/ifFZR8DvMU1CEJYRjuFvoW
cH+V2gM6YyOHMcuZuaYjA16MxseT+50plqCZJKvjkYTDhSYcuZeDAun28dPbdfRu3AO52/Kq9gTu
MLy1G+7O2B+746vqe0NC8W62Tyb+rHxVnOWRgw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NvvNy4fG+VCfM9NYumsm2clZ8IZDrJQ3Wi+cnwU6WbSkr/joDlB0ZRXsdo0mhVbkhlHdY0OhRpkR
3RYDWBuljULA6BTyF1sag+KB46HFjV7grhZmVLUbBkCWRKYz0xq7bDcNxf7s4evpI4rWpbAGWyJ9
TlfOT5npzM2PM090g2k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KN7EzciqITw/PNwj48fL1Z5o1AjZa3hMKXx25N37JjIMxkR/++b3PX0LoYvLH1v4MmFRO2F2HE6o
+A9StU1NJwej2oLxLD63NMJa+VjJBFCfkNayO25s8BHSFsZkhjc8mIC5S+PHU5t+p8zDOXzJvXOx
j/qM+zNzxFnZOpagckJWraMSJbbFjRIGq2RuUI6DTykdz7949XyxajpE+pE2TrgIaNudJhMJkV8s
PmKxeai9osJTVlAQyTdS+HOwcKIcXexlGTP+JSkiagntbBuHEhDR83LTtvkaJx0GY9b8oHB0RXsI
Jp2E0CkC4MgVpkaduxkwBZ7NjlyO6dFeIGiehA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35376)
`protect data_block
CSpwSTdo6/eamr4ITKiZKZXViVLsrM3JmbN9D6yHRBmmjjerEnp1S5s+3Ofjw/p6nmN0JDgQDbDX
lqVSItfpkVGlsQzjvWXeIpJZMBfm3sW5/3vKX6TCC8zqsyextYuPLVoNiX/KfM4t/7HZmbN6rSXp
9MOMfG2NQ9XiX+uKM1Jqv06envGrp6MUWqzlrINVmqbqGwVGhow8xYtxGxwIDaT/o2XV3fGG0FJY
RIIQhNBcQhJttOOZ4EhMlmoToULGSlb9gW862Po8s3ZgwIxqViVwJyEeohsvr6KWXek2FhPLkbO3
ASd6vWAGoMI85tbijRVjNR5HRBtg43YAWmIOBBtGs+T3NusMmigud451+vhCQu5mIjoOY1DE2G7n
VYusWtkOXptXCm6PLieTelrNVMENzut3VyGzQoqoMuT7TTEabS2Djps5RyCiBBM/X+MUHRsM9jD1
dweas0Dpbyt17pBg5Dg44rSkMqxR1vr/8gXNQ2DtD3g0sLoQDx1RfQyQ4n/bfAjo6oOzDodUZGEO
C0LB9yLdEioU4taCzHep+Llm8jm7ylb1FdG1+959/ghyZZmOK14STMjS9UkLGooiinu8LXRSlA/N
MKM8JeiUJusVnev/2LivcOcJcB51G7Yw/zjagKU1WdsCEMR0mLxqJ4shrU/Ox+oldiZW1hBcnfZw
qXBH7QFpFvIrcyhD1RaMg6ofAziCO9HoLuZxuEwglPqOgjC/R9NydDyBwltgjqKXf9XtoStQX8wK
KW0fesNbzyW+3DRlASSQQjyUIYK8Z86TKn8OzdediC5lCW931WL84FT2vjIs73uJ+qBvEwGcl4vx
BzTKLHG2FWDEekbC4uTMe5cSnMwdDrj+SZ1phRt+Vz5IBCxaCmb92TVg4Wi63UXf2vQs5zi2Ovl6
P/FsnNHogsL5ZgRPfkddNiFjcwpXb7cyb9WOhw4Od6dxHv0HCZyea4wnICuFnbGucQYUTcJpn7+K
31SSBYX8Uq55tau3WtoRHQGYolBVakf1yQFUljMsnk5QDlBb+glzqDYRzLPtnE9LQ9EJ8pvK5oXJ
15PRlIkm+ZLMh+924bdjPx8Aw8Vi9cuuAlRkCnMhAPhJPWUMvPf+1PD5Ya8uRk7PybEHHC8jdSXy
v9MB82i7NmEK5yYwCmk58oSlp3cEv4/EF386tqOhyhQE1X4wW3Fe0pb43vF8Pm5GcDZYLnhkw1Du
9xcaXMBhBjbr9YSTJ5zKxfaU6GTruw8Oq5JmIIAw/7jCmWLt40+/CvILBgitkCB2sJVmse/CrAOO
t/+vVJFsrgwk7UHvfJkA7AMmOQrptPzoKKaGZIXtCGI1lnadRDhPTmAl7PAjiWE6HFPO8luDc91c
rccRl95+dLVwWaKdGWGnzhXtRkCSvWLzXaBKS4X0vWjApfavZMKK8TzPSKySYMQDhnbh5xavFu5N
+zI0P6ROtPoNTgBfhGrZWefWHJJwKtwE0lN1iOe30sOFOlRErJFhMaKLC30uzXw8HSjKc3zgeypy
lP9xZid/VhKyH0FhmJOZQbAwrunm7OF3RSZuhBg8zjmm9mT8r33Q39Fj6aoBl0ryJpah/vqLs/Pq
MAzsP3/6+Dl6QqYfHC5s8GxiUoOZQBZOcxocUJmOgetWmEqoEVTetXaPK2NppEZ1WJAo1ZEV/X2Q
tWN4uVyXti/UqukJudm9hvqQxz8xdfupp2izNOfFzeq3A2Hl29aQwO5ovcN6Tj+e9f9B5fEn5Y1+
uJFMGA6+OdoS62XMFcQSywlfhWLfbaHWCWzk0Yi3r10DfObfTmrGG4KffjxFWaRQY0/ZxdBT/IPy
FQNQVkolo+k/qZDI3zzf/xUr2BAARFT9kBm9xh5P+SMto+2yidrI7iqBlbejIxZ6SE7N2ZM9zT/A
BMp+aV+2BMIyje0XGpUbdVM5RY7GHoMAcIoXVoHizghSZNThUydYPdb87utfUEjONdgxbD+gIAOd
lpBRGCmz/DYjunokbdAAYWWkiBKxuuUQe+KKC1e8sv8cmMGQIYxtwoayoXqNQ68eiHCxX4ieV3YD
6pehduAAbT4k4Zsn1yGw/XMskmzvArrQtR5n4q0/XBknt7QyXC++XdIJHprS8kMzRVrrcNIOPe9D
DMdCUaNotpHvceBTCOnopfLLs6ZxFxMEWFaAKHfldwz09Ij4ZahortnQP9ZszEgNCc/XiSdTaQTI
Ile8xM0FOGxr8IaLqwFrNrOpbpv6Fa8UFkxIbJdtaihIyurQvvrSIdGuLWVZIZa2/9Dl3FKaCxtp
EDiz+DcBgi6e2eJ/1alndjBPqPkDFepQl7HeUYSGGImYErbjX/Ql0R0nc9XIqRX2cIZzWATadKPG
4JNOGWPqQnZlhqp6dGkxlL7C+hTvwhPK8PwsASJxMJh7J+PgdmcAroktw6NeLS79YAuKsQ9Xvg9h
sQzqY89LXzGwKAywS2EepKDKb416bSObUDVD8ySfzN9AeptDNI9tXF0uLsINHra6y+YiJu71yvWT
2m/h+vprNMbd5Pdq0+6ahCG40J7gVZzkIYsHrtf5LSxNmFBdjR3uOkds0S14/ix49+DErbu0G438
4cYxigShs4Swp7e2aSgU4jkC0jhbELiQVc5VLTeMMl5NSxD6MH6wn/6/ppNFnOp2DIINsHaTLXqz
dnwj3Txc8NuFEHovL0wkvDRj7F71WmmcqT4pxpCPaoRnI5cqndke1dMiTDLO6CYvoA9eNBvi34zY
WTd1rd+QcQ5fLkiw73IZI++lsK1NXZMljkNAlUuZwoap1bKk2xsZmAghWIuEBkmTuHa54QjrfN0K
vJkdaoOsyYr6cydaNOTVIt8mehrI84dl5DhHBV1xYmXjyrDSEvw/sJeb8Muxptdcq6eJSGXFtO/Q
6ydB46y191gxj5IjCYu7nRQNyRKDEKtXTGpU+jShMdcvQkUOkN5LVPvQ05LRKFnIJ9wxkePig9fO
FkGZyFHKRn4/JXomdjMhWuPwyI8oN5RDupMFI8A36YyfgIHp04YLlsL4/FrHq/SkHQlWUoUKBIBX
zqvi+3CYPgr24JVSTyG2ME3og96mFitWwvbYNNP4pYmeQU+vRR7QCTGHGXUzwx13odamg41kYK0z
GHAhwMAUk1DFSFceJ6qy3yjHZNjHLcFDGliXeDcrv71pga6WYTT6ie/XzsHna112r7b5nJxIJEf2
BeWS654VWVqj5sfGKqKCS1lYkXJjYuFZ2F4KxMzyu76PTtHQDhPGEwrRHqkGJ/OYJMe1jUb337Da
A5KkANX0pDrgXdJjXxJPnJppES2ozgfMH740cV0+/vT8Ha1ke1ZL4Clwurfl/7+Yab/TOldQr6qQ
kfTVHxkWxEdXiMWGCbCFbOLbEt1tZBFZYRQauv/yIKkY1hikpXEE48zXCCBqMT0ScqNtpSoVVJDb
GWKfQTJqXsM9m3pEYkhJFA1gRdIezv1UwlIldiAiX+6og5hlCerBhATEJAF4YsszzH9s40/U3DxR
pEX0pX9iJpP+7JhZsFTHjfi/tt6RZ+KNRIuQ6g/M1RElYeBL3M7IgD8yWTDGEB17Dvuuhl4fbHVp
NLOVQRpo7Cszwb8pDfO9YLhQ/7oc/nbs+xqS/O3anaZ7u4grEPHcJw4ceOeQIjQvJ6lDl1H4Nhbm
xz5pAutfF3bU2neqNRGGmERXcH8TLiyONLecSjDpXIXopBAa9a/asT+IPDljnFBXSUt7xyTGstMo
37AcHFSZd/aGozRWFyuw/N87gSFY27V4GPGhZAi513OrkIYRp88+Eh8am5qmpkzyaaQJ7a//UpXX
qC2zpFFFJuel0M75s0kEgqZZj8RgY+79fAGOMurAmRT895Tx/Gg1B2HThWMWIEOMJq9Mmo5UQIta
YRMGED/Xgni/IZE79kSsDhoIuLbFOPlLTuoCNZwt6S2ncvS8kyLk1tmQsL3dn+N4D5vKC4cHM3p7
eoE5JSzwUR22WDKnlsyz4IaLT0s1ItvmP4SddqVI49PVMIcS8kJN/bUIHEnbXWf7ncluHfXMCOmM
vBlJETRhG/F+U35266myAabWwyx7GPWxKkK+enTOmOp6qTGw5yRGUJ9rBTMjg/yB9ARnEMIOqu/V
zIiyuOvi/9D+cyhy64uQzhi2yR6p9hw9khFfIS4UrgbWYII1Aj0hqe2n6x9//hFz6lbvqXNfdxDV
ElPsc8yTi6fmDQZFS7uqdom1jnNgq1YRP5QIwRiah3o8olM37ZTXyfvJOgv8TIwBH9ToTdFp79xb
YBxIxsVU27pczTm/IqRSvYj6Po5BCuAZ7q/7AB3qg2SeCQ9/RVRqypt/Ial6F5FDmNe+mB3m0EEM
2EdHN6iggyAHCWKmGuIInD+RU1g9Va48I3+6tXA3LPvveqEjE5MivUSdvQK5a72Tm+Fm42ebRrU/
hIvutIjuI33r0uZ5jK/XAKprf9apVZUTMtykT3Bq7BTjtMDGAToPtQFw8o9F3ng26QZdDSbGQZZX
OQRQ32WR3HzlfqehIZ1m/mheRuFEvPbuc1WMp08AOsbFTeZSJpjcV5fXJmof8kLm3I6fm14FYUp5
D9ladhGoHXhoEjrQSZeDCoteHqDXBVo3WKQTaftPv4D1tA+HXcO17MIzDqAaLTEm3v1CXxOBJ3AJ
736ZQP/m41T94xRke8WuddtJLWv0tK7+XoIcE5PsQOpbQwLDbIf21ljBUXykYrKN6IJJY90BE0vG
3KG0lo6v9TA9BUc1VIZLEvXX1IfMG4qIYJfhBJ3Tjj2e25ZB+aK+MrXHw04hdapiDQHDv+0Hb1rz
uHmFqOj7YrBeqPGK5Ub3MvOvy2D5sPl8j2lygwYijV19VtIoWwUn3PP+m3G3lpLDhWe+8eoFvRFk
YtM24808FCGdyAMjTombznwmmxn81gZCa33H/FXRJSu8dSj3pbVrrviJRZma5+Foz9pKHr9RbGrM
rSm7DLOBbasX/CEbfrAH1Sf26j/eXS3MCMQkI6cZkuj3Tmrw383E6LSK+wIzoi7YSOoeeD4NOWcI
eNcDemN8+cM7+Ng1+z0zXJwb4O73sgEF7NMOE7C1tg5vjBxsTfz6YQwa/IgHM8fTyeRFXHLfhU9V
5PfFVMm0k+xUJ7lFqaUFYXmQrZthY2kZlS8zrWC2jPRNMzbAw5+2Wn7g8dPjwH5RYwJ2UEZvKGc3
B7N1ugnyAiq9xmro/MlACemElUqpr9TMaHDxX6Ve+NY2+UWuzWKDiBAuEJp2+FiLfQrsDqYWPYLt
rVbjeUUCJt9Ojin1cumuEgzxrkSVsQLAS9MHW61LzxBUTGWIj6tLbwtpTEgMb0i/uHUiVDXERAAO
SQboO54kwLG5l4Kc41PbDnyCcDeICgXHHo2LAruBqh5onYhmDecZRYKxYqF8094J9cqPp2rEITmz
4XnanxIqQpnE72WEvs0IUglQEfUfHHU3QaXiVZuZ9o/HCaftB9DFNBEtCyq6qpi25ynKaPMN6Q5B
GOiR5JY2mvU6h7TuyGfcLwWOzHKhZPv5EuoeCkAt3FnWRyIUS1LlJBValG+5Nrh8xKCgit+mnAea
qxZGCxxfeSkCMBDJtYJ8fcJYgJSjNcgdwokjAo0d9dZuBeknk3WHdy4MawoQ7QXHxti+2huv3OTZ
tysEF6Q8qQ7YBa5i8VW0ZWZF/I72MLK/vyf9f/V2mZzcmd0Et4NlnGK74yNDwgZrOCgBAmHKQS1C
6qUBYRhqXsCqbu4GFWlABftQam95uUcQgIHFRjJebJsP/GKUp5AEKHWAAth44PMDdX/NbNziw7G3
Ld0281QINC+OTyhPN6kvKHwBDYAqECLJJAelTIJoC/eynIfurrxe4JX8+sMGcEHVW63+joDlhbD5
lyxLYaFMmC9P9+2G8U/UIW8rwkSctF5zyMKWrV6mNRa+E2xDNiMxwCy3Oe1mwNBLjuo5W8qFFM1D
5tlnHHZfwNqfT4Qz7c8k0rxAHEtjSBNcDQbGoeIcTUvNdrhdbZZyhJl4sivG9KF86GwqB/Tm3QMR
u3sI95qRCT5GiszJwIUSp4/1pnUJZvj6sQLnddD77MmIBVTUs59gUywgBm/u9d5rQK5IUydxtTaL
gEHsU5E7cnig+ehKsP1JE3c4n774vt3KxDw8BcqY6Lx1dwGGSr0vIgF1ksYbkQ9qsbbwkcUZ0T3X
xfSvsgbuH8qmZ1uXB/ZF4eziruZ9d0smnA7kROzhKfPXtvcQB6I3vPgfhm+3FpGVSDoaebHhwToV
eLf7NSok+NU7aoxBjhFwlRq2m41B439/7mMZBCiJ1rbVVbvv5Bqeijo0RqO4THEZDbSlbvQFBgXU
Nx65nGPr1ZkmoCH1ivNm5ooTTNaKmJoVwdWsGQ6bPGi+X+Izg/uZ/KOf4pmd/AHO+cZ8TGUgTqh2
72VyxzCe/APuiULJgfRVapqyY/PHbakWGssDG5T5Hi0O2vy2ClwJXxVddkVeHw26sNcir9n0lF4b
kabbiaQhMMwB9btQutM5hb9mtD/hcTIJ6BMogQtlfm1FJ+XQHDu7Ysc5n9nkhIzB9uoSGjtKbsY3
laLgbkJzMAphyjtnnkO3VDEwUY8b5zi+4NaX2EfnKg6mbBaAPk9q2Gd28K6fDLA2yCm/I15Qxxa7
ntYuxwgycdwtOAcKUsxjVPRMC5u5krCebE9FxKK1W9roImTxPxxD7U0n7aS39etNKCJkeWKH5t7h
kWDdS1L2tqXKR2TwefcGDYD2b1aWg11CQW+/AfJuBnKSoiudJFvAExorY9ojeKcnCIvRse13bWCY
klIbuc5qwwsJQDx2+KTTjdvaTnt/jpJSjJTPJEycD9NHvhf1vT9tSYmejxADTE2QsqxGWseali1G
mmRqLUccW44kNJx12VQLtNljfxLEc7YKh6Up1pg4gr8ZFEtkkIM6BxE6mkoG9h2u4qz3z/JAE7ad
cWp7XOTCSMBmkw4mIUpN2wiPkiTIum6k6j3JLX0OhpVNcbx9rla3yf2Ynf4C3Yh+Lnv41yIRyzZ/
sLv0HlMxzxhFSLuIyPyFY2yCjz84qgRfU02lMoFRGh8A8oQu7FokB63RVq6ZtQucCKPDblRvzdm0
wJY6mEJEvRDNzavgr+RcoCmj8DtSrjKUzz0k55BCASJZjrJcq0vBJFXbZ45HoF2X1K1iKfPAV6E0
EdVMc48KE6O2E2qa0X4tYByE8lJ8WAWG4uukqOaebqY+/oahhh07b7JSpzEB7VilZXS6f8p8LcEK
tyAY9DNGnofCdxB/Pzq6Z4tGC7Hr80LrPkYop0ShzJtfw54OMFNUdKYnoZnZ0vEGHk2m7QuwBbTu
6oqiP8CVXUewMb57noNRyoz2KeDSYfymd/QxnmWPgxdcc0IIWsragMJeyr6iXJcMAg3v+vLUdUna
6j1jU/+KgbYjc+Da//LC4IfqmX4wGOsLZ6dcUpbj+q1YPobRsTA0Ntgns3JDh8NA+Zhxa4I5kZtA
1xlUq8iFmmNAlKCSR159XudiV1i6Uy+z40caKEGGbKAIwMIAe1aOBOdwX1IS+Jhu9VJ3oYiWMRt1
PiU597UuLHx9mDC05lHj85ZxS7MBDImLlEIT6uKemFDojErKpYktBBhfCzEoN4pHbCufo8Jyzp2n
JBPooPsZ4sWy8sO3fRaxBfAnB7QsA3Uyy9OzgznK5rzH/lVO5QMbOA5nfnwSnVh6KPbpFSZxmifc
DRkJkHmGp6a9JiOhlc2oa5pxRz3SWhO3qYzHsM2bq6J8jvkacQ927ytUSzimV7oAdcyGolfZx7oZ
DrD5jBwDzPRcnAxRgjCLs1isyprX31XKyAK4VhGdLiHlL1cKCxYLkldRjbHElCE5rE7mvtVSnGa0
6aJjntpQmFUZtk6KzI8BPnxoRdm30QOkBYnV0fuJl7hDCMu1w/pwh+u/yLue7EaDLs/toiOh6ZeR
YaAuvqWmWYxpPvQ6/l49xteARVXghjGhOEiIITdcZOJ7tnHFofdarJgnySTxpcVAEtTRyMcMhq/W
lKTB+rarZ0G52MA0SLprN43J3r+MghrtPKObPQNAEo3hVRLkKP5s3kq8G6XgyEele4pGjjX/KDOW
op850i8DX3TZKXKHGGOtUbs5EeZSo2px5cRCnnFxx88/s8CoahxPyMjRG02KSFkkeB9EKlQr1Ogk
avgXFLiaoeQc05ac1nWj6EvQwrpaldUAyOTbE5yDdR7JMaSh2RdU/MKvXt4jsm1mTbyx2zewu853
SV7myZnhg+bzVP7pl6Rd3qwRJvnhfG9fWELivJ8/4qnmCp2BkC10qOu17ce9ELDwSZGbxSi/8QrL
memU7wYa5dCIXG8e4anyravD4LAlm3H9FjA78OEShuhUgX5lySZy4Vyjku5kygFQDh8GLceiaZrG
h1i+nM95U/CdL4/qk3Po7KOcti2nTMGbSqExNUhz8uyRGxpo2qJyY4uDFBFr9v+C3zNaJbTfEZvg
APlIGdmgND4xa2S42e/5LhBdEKCdeDCkELO91kLqfz0hVcxwpipIWmpi7R0jeCb3kQhUqpkwh77Z
xSxR7xMphaRvINsmGxzeYBHV7t7KpIi47Hw7ZzwZGj6lpKoP9Hi36XP3aOV4nJBhL4VPWDskHkZd
WXMmIyZkEH3jTSx4VJ23PeIWhJxEebUzdjEb+DmMh92kyNNjDPCwT2LJDcPdl++kUUpLNfaj4JUJ
eYcLfi8nvzDqKF4JBWh9o4CUrWsc6hSJDWmqHnA8xa8DJ6ESG/bDmp8ztELV7SkS+OnAhrqYh/JL
B/yGjjVdyCn6wzHw6TJ6quLM2Eh8+uzCsIh2p0kF/+RTlHXYW7xgyoUoe8rtETylcTuNPoLv7Evk
6UXZHFxKkO43EboNjQu3TZkQTtov6NOjb3eODAWOmt6hOvfK5Ey2omUr+g9YzOPuZ1TGkDoBJ63+
tZZKKkEeCg+tXLBg0RO0dog1EdoNpDx+bloBD8IjfQ/mc86jMbggt6ryZzsrw3fUjmgZh4sM3+qx
kLOCzU8ZkwViOPoITznIjRC6tmO24J/VdKPr1OE3Fq5IfbQsHNaqW5w9r7kvhWzHMhCvtl6zN0R/
4P7HJboiLoV4TGp9mYo419W2zV8nmhUvMRk9qyAyq1WeBol2af3PHKXkTSrEs5gOsRMVWItA6a5l
qeZXFLrbGe9oeCbkE/SC4wn5yQUGZyAr1TiIhTvY/cJgP6DqoMn40d7gAwTZzJCeX2NRms192tUg
z3FanHj2DWkb2CYHEiO6JOsZX8DLKJT7lfHznc72c/lyAsdAkmCF0FJyExPUgWdJC7U0MoKUY/8e
whYylkbAL0j29DnwwSFrqUa1BchgwuRJ1Qy47P5oY3nMeOjw7+Z65oegikHHtSF3YGxDjJZ2b7xx
sYy1BVWuT1LK90TlnsMWxtwQDD2Cb4/RgqPuwgtRI+Y62dQtohQh1Xs7E8TzX7SOwFYl0lLCXxcl
+nO28MA31zxHGwKoICwOczT6W1cQdRk7ipgUXI1V6vJM2Y6Ax+kdbS5Q6d0ubKmvV+9y7NvyjkmH
toXAYpaHUxuCSm5Jc8LCrv7viFGdHHpovKKHs87lW0IBoLbr9QrnOSmKNAOp4OOJI85GutWMLbPH
pEC450Ye9iawHxWYbWBZE9d61GLsYyrKu/zJYqo9zXXLMLihA4NGBtDzcjKBqaVTw014pgFJvHTk
6Q+3Ibm4rIFICi5b9uh9PSkG9CioMIbrppvuWfJ3gmBONU6IwJXc9vIWXzPYVwT8GOxPCWrsrwgg
IITEwtW/m0FAbPx6e2THgPsO6D0HChw4kcAS4cKVLyAPwP376uXjXfYB5IpoixhwWqJUX5vQmFCn
MKJ7bPzrieIWR72LMVFxNI6XdnG2VgwksMh3a5r/sCZ9jDg1xfvFjEj7wpehtaeBjkY4CnQnnVZx
Wnk66lBnFICnjKuJ0S4yYt/fs+zME9mKOluRP3B6EsbT36gMbWcaC3AC8bNhpEYQMWgwTNgivqUN
9M4zUg4wDYbOub0DDxKPZrgMIznHvfuAE7nZKKKz+F5PKr7I/pKjBhlrB3NWaG84dVSODjQEFm1+
ZKZUTnye63nvxVTmD/ep9rUsEeZzo9YaaM87n+/KnDuLI9B78eAuynjO8MNlAy2sJlTYokVM7vgl
nuKyTQRfEq6y1vFBx2AhCs8LMIJ59h4VFPePlLmw2yGDwaZbIDnR2peK05KHS+GIvT2eZce9Qv9v
4mFZ8CRccSqEPhw83eirhOLQQa0aQb1JIZU6cUs/XrwKWMjJayQP1juaLcNnlg2wi5R/zUx5pn1y
aU5/Lp40K+xNbHGEkdwADjenlYzhIY4sU0SPEYy0Qphi1JhlnLKiveAj5gFeZIyr8v+FqKscXJOM
1Auppgf5nEprf7Vw6bmjZ8yIuLLdWmJ4kTqaZADMNLNjO0qqmKK8Ro/CrVOvkQMUPHYB8GgVcT21
/ezZmdR+c5nzD1m2FRp1mVFcApe6/X2NJuHTeTXN3x764gKt2DOWlkTKt1ihqMZaJ1FHYkzKv16K
C92wBlxPtkPN1c+ULLY2xn7Zh7d/ZL0kh09vq2OlyKdInnx8m+YXE8l1XvFHYEeu+jB1GxGq0Sok
apHiyMQ8KaoHtn7RADkEjodqXbJmDFokvkjPeMUKyF0yiKKk4Vj9Hqp+/gm3kDquPO4keqLN2bW4
UCkQ8y8DhJnUigq5VQuyLgud/teMA2FFcXEvOYvvXSrpxkzV07YilI+6+Gya02ZEyWJyRdSBjjrc
RUEvhBgOn4AlJA8iuWhYTLi830i0pDGcYHMzaRlfKQYFq7T5nmsYW6ib18Oluotf9AZCnaEoVtyF
ZjnxMwo9JeeWsiRH899M4s9AMZiDzcNVQb3fRKQr1aHmTFMgO9HVadtSga17XU7TdiIixJjZD94V
Ceav89ZIIGOCE0oj77+4u7gbapuja4nu/gL/+ieE/pxb4gXiQslDymLkhVH053COOoh48ru8Ogri
TVXpEakmEPEXbIs3zJuZWbAo581BgoaXlNFfcEbb+BIY1/96G1K3rmrnAflwlPyiPGSH+pNPtlw5
k5kBCnTNRpzVO0KRQ+npuRITmzrMfp6QbDQr5Xsjv4UKSFhYMyZMMaRBGJAWATq4Hx+ewY9+xYKa
2q+wsvd2h1kYD2s2id4Pz3PvitVoLd2AXHWXwDXRKmPwD8tjatkj5ggi5Cbps9ibo3l3oW2qFFUh
udiXUaq13uRqE8yAYvIN92jcbm9eGF7U1obwYohZViCT36ZJmuVPKUZhRC75/Xo9P2ZknGAHXEAu
clrLzyTpkl6roAU5QWpIsY1cMj11vL7YhI049osTM6dnKQAAdabnZIsiPeuw65Pt4WoptASoLCOp
MTYA9PPjHK1v9giwDtCSSE4Mi09H+FGJhXCRi5efktSsOzayyhuQiP0RW6dYHbuG9WaoWn5heMiR
bG2pSHxVhB1aDcKDyBodEBFS6I9wVFVlwOkrTAh/iNlMjKNyZeKf7SYK0gq85dQKHGJODGZkgKg7
WC2GiasmS/CnBfrEbWLHAiXjeckYYM7ehKPXxbp+VojXo2ieEKHwhFY/YOCRra7yBr1U5diK7tzf
P3m7sZCLb/w20JGUbcvlJqO39Cy4QFeh0bCgJJgLqjZgJ0Cgi1r9S5uA/822LO43EAgpiLgVQVGg
PmbAAN813XDqKlvCVimvFLTNJ90Eiuy5mHMsIa72A2g2O4hN5sFO758IaYb7m8CssRinruXUrRLG
heDvEmGDTIjZ6EVtlA1g1F1EJQewolkNMCLdEURTCfqCsLDhEMBiCZ6s15ptSQ67JPIEjztdpRdT
Vioj1s4ZUMziF6esxeEUmn4a/ARrvyrogLDOb8sYFNGEbxzeJMaINnEWbAvHP+F7m4bgfeyBaDcW
VxKgaG6e/soJQ6WhzLMtHD/1wE+1u4TFsbmvOhxDa8PVqjhNjlxA3oNR/TRQntkJMhrUbIJFNhcM
GJX++HjMx5eyLSsmR+dKGycNPUYvk3LvNu9NsqmVJr3VUYa/iai9CIEC1T6F0pcy+Adtuu5cJ7xF
Z3BLJj8uxstwE/4RByLYE++dusSmXxFsECyV2o4jqTFB/zcVSEB+EE/Qh54ZDiOZ9swEtJGXJ0vo
G8wsRa17fsHQXy0kLgR3pF8u1XbS50aJMiRhWvxFOMced0qki6SEtLHWAYnrpg4rylHHLKYpaZlk
N+bUpscHKObKYvGLera7uLScBSHrMkNC5WV2dIZCHQLqzrPk9agQ4RqnJUErZr2JF8CsicmLrV8j
wDCMI+GWqN0gQlzQ6C66lJwQd6S8OFYEGfjStAtIBt0Q1ZwYEzy+5ugo0cvk7HVtF0sIuZUZuKN1
8jfCOIAw7vrhJEVYaWqLFopwa4ksJ1lgsuMpMaWVReLERNSK4woq14pnINJh9pYOKETqGLXssVWF
n5Y+e2CzWFgxOvHQc6MlU3kdRfUE5a2CjsIbUhHQcI8jVZm541j70UtgfEyQAZTOkG8eluA7eg/Z
zliQGYfR46dY811nw7O4X4XX8Rt7n3ZSh7C9fzPkUO2O5Ze7XWic5nTAehlDy8613nHFqF82wJih
J1rFNvgbZMZ+K0n+n8Paa1WUo7LfWFoMgTPjU4pnPB+BgYmt2tSCmslz0wUmqluOWuwAYfgOgwO4
+/udTeIPq3ot0Rtc1db73333Jqe6yIGQiuljLAjM4ut67cPqhOXlL2PwTU0O5OMSCGOmPLRxvYFe
d0w2PGJz2QAYJBniqiqkJFA9vq/v7yWIeExl6sOF8VdsYhHYeoACdQ47XRlpEBcEbA9K2yXNiXtT
m63jrb0yyA3a9sp7k1Euz2tVOIKlKyxagdKTOvYTlthw0p/u/geYn5u4tbRb8TRGVdhKureOyALj
pvFEvO1QocFAtFCizFtuSGKUiXu/9GoucMuVhjfgjpTUdA52O5B0yiwkz5+N/ZKlE0orxDyGAPwa
fIdE3PLzx31LPjt10+eXxW9vIJXRcgDm55cG1KIYNKoGINXzxd21w32llJCE+TI2iD1yFJEZexXc
yiOIj2A5LZ18z8zyhgD0xHB3rtqeTufhCBQGntDy9EutohVEtByXJkoTRlGSI6W7hSSBtfTKpH78
81yQlQXI3/Vz8eapAfNO70D3vYBD2R7ySNvgapKPBl6L81I6SevK/mE9AEvb/8mCBnWAz4GscqHU
QVOC6w48l/QKJcf+1Vr3WN9i1JiTgUIWFPUeWEeTUjkUeyfLEeO1eQrvHHUeSPsdVNKW4Me6HF9x
E0yV+f0NpRfBWL66ZuIlTC7cRgVEsLchNXbGENQx1PPCSXT4ntQjAH+iWCNd3ZRlkRG6vZ3nOljE
1GEdm4Fopz0KRyxfaiTR6t0yCerZq71CXZUHr5h2nbk5JlRPd5e59OQ9uMO7FgVNDfSKcXGr9oLZ
gzhaC5foWw6O4S0OPjiKXPPcOAH0t5KeCqnHBaHh96t2ImQju+4cJbArO8rwIs5PNz1Zh/gGHZth
GBPVofAguLNT9Eemh0BXXnvl1DZfdG8h87V0ZjgsV8pnHk2xaUm5BS9/wMWfuYcCyUZ6O2nJJtP0
40QA+Mh2quxDRzeLb04DpzGlTEswgPpYAkRRrSJCJVp3j1t/wOW0zVpVMrEACXBDZXC7ozbn7FMt
rHQs4DROK/3V/lQOBw7LfzLsk0TWaRcQX2MmkHIyAPlmR4hl9VMt1B8+HEva4muS9Tno8MpcJtoV
41WARTPH9S9eEZsoIrOV/yt7HH5GxgB9yQyoKeqEBbrPthiXbLCEzFRGii5qVGgJ20kkjFaXtnLA
ccjD9tHZYU4Weq0UrfaDVu9QV2ExE/oKSXaPn7r3dgx+VAgr2zE2YjEQGrv1a7vE8xqA9EU/up6M
/Ncg6f+PKYy3o3INNLz9KNWJm8tlSNs/m+2tLoYFqLIELmvVvgHL4wZ9I5/XltEgVGsvyu13SbBn
U/2eXNLIG4/cj9oWnpFww9wAlVd6P6F0Ce01vyDly7ATxczI9x5FtDw2S9og1E/u2ODDyeTo1qVk
EwmktsFPaHmbn2xOs5nsJlyX5O4xQ6tXFwgA9G8ypBXaE0MWWt2eiFL6zecsuaFD5JXHa4F03xnl
Lm/7lQVGlIVQ6/7x9eds35a1Gx8HS8m8Ck+oxYpfYa7CQv7Eki76KDOS0p1btOxec+OwXF/Vccqi
SFIr9osawo56xKk2yqLubQb416RvmgN6mMG2gKzbcVYQpmHcMM/KETCDGo4FkY7dCWdV6Uupturd
rjj/+w9O/gxtG1y5WamI0uhDy+QEYjzL06UBFaSwS65BcfJieX11csYEoS9B9lIHPCgJIi/x/06L
vb6PlyJ6EZ/g42w/o3JQK63lFb+y++5fSc9db7MBWtpWoIVTVuT2EfiS3XmGGOPgWgQRG7IlxeMl
fJcRZNE6jJxrwcTPN+NQ7LF0HcVJnShvNA5pOuSCW4YLh4aBZAhjx/SuHDNAbJxFM7RYDnvURx3z
zfj5pPzcPL5AhgmP/kgV7LXrT8G3OJI69MGUC/EyXZk9BrrVLNNNStUyta1msBLr27NysIT9O+bs
AKLZHDz++Luu6jwriqTAg70ihgNI98Wz+nZDBfDrVf5iGhMz0VQGoyKWd7AVzvX2MUwOT4iaLV2+
31zzc6V1HNOBhQMuE2N6aLJuAIGzqOkA9oldvvFZRjCagpecsHZtSY5HAmEEkQobrBvfQVXFNqdC
P8YLURz4JFU08lxg0OGO9eS6jmmPvaqQLrI4vMg8MyPsZSeGtzlD7sKU0pMeu9ror97Ygn637Qjm
3O/xz3dM8vFLWLdRCD6IzUPigXgO1HjLqMy8WQhVnehbuJ+l7vw5bZvYZuJzNvi/GM8XVf5egi1s
khXiwksiS5ehG+E1ld8SQY6cMezACJk51yIu+f3WSTfmlYGOHUQ1xMKx61c/7mchbDIR2fModJFS
apvIsMWfHNBp/z2iQfFtmPQhTp3hyz9nrpDlGFzzmzFCaIDIDXmuv1XhtxxofPsOIDI2HuTDvH+r
/5hGWMfgA5hebXIgNl0YyAtabwP7HuQzjPwqFoMjzRn223NLkjY8wGIr+3OVHZIboJDpALZ9iZGA
Lp1+hChYoQ3uVyQ1NpnXog+cRPLCSkLlftmlHWL4qFywaKqXgMXcoj7+xjj0hdqoWZ9EYsxbWYeG
m5Zcn31kY067G1KeZLsPkjTmo+7H6sVSDEo5qQBv6n5Qe7Z0nDjg+HmIUsDiKMgVdLs4EXIxFuEx
yvRhj0HNtArURdOPq/dlEXz603U7iOnLlsCjIImWupScg89erJNIIc9Az/PpQ7f84EDjnIeG6ctg
nBJ7srvGiCy3tMkK2QzVBD6u3kxCav/jbG1kFHGlZtzPMSrajZSvaZXyIwrM8f1y0FIlU4WmI000
23GZA0pz/qbCydTd0z9ypOzsllHqYsd4pkiWD5L3tk8TfcI2JY5sAadBFCOPan/PJznBZnbg3l52
cP0zWR7HEmPp57dHO6HlPUH6VT4dhq9zqtb0AahWvrrDQogApa1qbNYGhCs01klPjrXdXCiZogzB
qhbYtmZA+g5J3CLi6EbYw13e91bej5lu6pBmxmDBIuoCdGwZnfKEgJ+zATdMptzHjozyWX+id2CF
tP9jun3vO8PW6vf1UNziRqITZe24Vugv2hhaw+cHa8BEH8z+Du5PVJHyc60i5TRGhjRWBsrUSj6N
wwRU+tijyeQyS2IrdX9DW0vGaa9pFmY3M7XZJCciwSryT4O+W/FdEC0QFw2LHYBnGSywXiC9Hw7p
vGiqsL0tOW0E+A7elaMPml8QLKJcUZ7SDVkZFY72Smoo1ZB2AqopOOAW/vR2eqnbwVjckgsYZ6MF
W2ucr6B/6isvbLtNB9cWU1+hdxO1m4cp2hkycpbyaKWS0QhhFg9FK4GlE+tP6eQ76Ml7PcOMR8XV
lCJR+zBSudTxi5Xs7L4T74RuSmXwaLTWeV+peiqwnh+vK1xFKZonvbyqU7p2ROANQHWY9IFaG+IR
Hzk0IqY4fEbSs7WmK75d43ggX0x7n51pPHzFRTOfaIoFTlcVeQZXB4Ad7oev6sZIZhLbWpJiXmt9
U/x9zAGTb0VwPnxQLJ6BsJ/GPth6+Pg46bH9zvOkXAyaz6sO+20ZnP7iRukSSPWSgyJOonW8Bd5Q
ZxM2mURtUzu1LmTpsWDwXtD2B9lZww3he9PCWPY+hql6b0gF9yGlQlTf46rHgD6F+ejM7e3ahg1o
CeLVYPlRV7Wb6rVQ5rhp9WDy1ApP3dAf0egH8Hb8FxeqmcAP4Qe6qFPluAXLi4EIrlOEiiybXHOR
YBIeWyJOxC4Zn3wwb0mEMdUhwuBOrdcAPqD4qcFXbu7N1RIMJXmY5ZIdvJUwzmU6DK6adKs31xl3
E+qv3SJIlvROfZOz60SAE1bjenQKFyenin/yVOLhvtunpX8Rn+22gZlagNXci2WveCzmJaewXrS+
xtcZAXBr1Kwy1S4cHgwMKlopD0KSLo+nPl6hZw4rumONqIZl1TlHmV0NPn2cN13qMvwtXACOT+JL
1NURocoLNjA+6RFcckV42GlCPK+gkv+ry7zV5Du952jKtX6EHnC3mnJRnRefBcz3AYYUb28tlxpb
hlVcuYX26mBm0b7nKKzmTYFu6IazWiKegiGlVYP8lUNu8Bu9JO6YXY+eglYShVY4Ss0qwjOIObx7
cIrxupTAxmpnWEigzRxLzncCC2xwhTBx1EliHqJ89VFJB198ZbPHQyMDJSsG9DpAAvfER0WLNlOb
t3dPFylIXMb76fxlK78fVFCkPMePRsawi3LY4oZys2vI7tY90xkbImXc+jt1Tga/F+d3krHj35BT
Rr45yLHJnhI4LoRVbA3Eo5VCC3tA0FDQYcx/JZ3Yr0ET3YOmaFaZ2wMvE1NIrW4B9TUgo5DLKQZK
6MAc4nSTrSRj85QtvNHAXHtdAWc+zwS83NUIhhZ2tS+QVHivc9+SIMSdO8e7P48rdHUx/IN+MYPE
op1trVpruQaGzsFp/osUfin9nNhJBtdz3fa+B9/cnaKeaDBWz0wFUZUByw3MTRx96jVCNvg/BSOk
PjlZQDtFsJqBFnjmCR3oRE5KVMMPTzpvW+x1nzYwAZCWLigkTEscHIdjPCmy8vwhU91stBVu99xc
XBr8jbtbnGcS2YmFFM29FkUbTEYGPAURCHn7Weqbu/HTIMNfPcYnHl2Y+3AS0Pxroe/FhW6pLcir
KFtlc7X+iwR++BlVPsMmoAFjPMKAPRpDitvkukguHnqlpw7q0RvnHI1L/8SCFi/KVFopo6x5vYrv
YFsPaF09s312HdLH/3s7hntTABZX/rvgVfYkHeMuaiMzMkoNx1lvogNiP6Y5AnKk5wDcUPqvjOPq
FUmWfgsP/iOEr0vrioL7XFayru8k7XUmgW3QpyZj/uBjtSUEoysm+JthXsGdmBI0sOMoAI/Ba+Hv
ay+V4XNRyXnPph+x7/Nklg0AkAOq0oDWf8GN1bGUU5kBict0V9NJLCfb4sOeEHTPbmO7qlWf+fNV
xCSEjeuIeR7MO7PXXF8RIHbE1AXAm3N0ALkvBGCNhNOljvIQwFtKodD+VLwePa92tqBzPkrmjpPL
jdFo4SJwA1X74ejbtQgEjpNmxwJidOR4fIabbEd+H38K7HrkfUFb6FsNTooXC2hNTtGmOOaZf3mV
ruIWqldTPCAA8Tka2nyKHCp8ETMV8upVaOQWbU7uDKQ9qWPMs3NbzDXSNNT8D4nCU1wtryf+3bKT
9ndoVS0KL9GvqAfle4aKp4ubgCW++Sm3BH51d3TUqdQ62/mrAp9ZE4mFl1F7ZKk/O4jDftXGq3f2
RjirXtpPzKRWNk8z1sraOcSbxEaEDL1CHOO8jCa45Eh3ilCRG1MbI3tfJ7n4tQEwen6v3FqjPaLd
eSjoT3QmG81rvXpxSSnnX7lPuuynzUxInbpXHprTfNLR8OI80yvmPDTQKINVl65uHNlc2nT9pqMJ
J6Iz5F12jGolyN3TYJ+eqVPUQDUTYkp5+BdaDA1v/Mg5IyD0/0KmSrVfZHGa//oxF+erIdAkI3/z
h+4Juxap//cq6xPmto9v8o6DZr39r5T87tCk1Ooh79W9EMFMTCdkYddpiU4CjtftGBV0mBYSi8Ce
Oge5A6uijisha8uZV8oAuRo6xpvGz03D6abwdCUGp1VwVMnYiaQbZ5y8OWZUwwZMMf8vfNews0ay
RtilHFcKBN2cAFtSjp4omLEZpoNPMMPs6SZUueXIMEgIOpgITTNI9O14rOSy9IvTYnt2X/HOZSua
nCa2qgOhLoMlk89FhLm9DTKXal/ftNyBsVYvwzU5XK69vNf1wzuVkUF/BbmkhrJ6x5+3Je9IJ4J5
hqohcJbT2pVVySm6MBV4jBSu/v6KjvSXNQ1ODEEQoDxnmI9ZS//AtvxqVIf8WmH2TXflDlIMwXpd
YhuW77/AN4LksPao2qtlpvnIbW6bpE55fSUFs7mFQTIkQwZUBmNd6MbMo/qfmNw9JnwfAXCc9HCe
merxGgPuz7u7Dnlfxz33Z8cdqQEji5gIYIuaAVQnxj/TCCPUOBU2aUjDgfaKOpNA8wv45xezlhgg
0XDstCYDILjxHqdL7ukl6zIprakITFIbJA3I9e3SDNY/MEWAIX1XBqmd2pvPscSewmSyhAbWbVue
YkkhEHwdZxhFIh2DTTPbs6AfmV9zRAd4z/1j8iuxE49iRrlLm71Zspq80M/E05n3XIsNqx1Flvse
6ydBryia4u7Ev+XNBvjJZlIIISSE3su+qGqvI7efj7IEYXTqsH0eHxrHnYzFCFE0bvlIgMFlYX+L
nSslR2aR3sIIt6ag+oqiL1QegACGW3gxvUkc385uSkgqk3FYu1ztQraddCBTXt4kedcmKP1xdFle
X8An2X+wFp8I3q+TwLfJqxTVQY2PokG+EybfznpKjfSHTzHMhXEZDMpVoZv8uYL9SYErq+WH87eU
le1r3zSxaVqVqvZsS/sjEEH1knjJ0XgFUC7gt6sJ4wzXSONnU8H+/hOFoognNHGGJh+MicXV7ZO6
fiFPVpy981dNEdrgv8TRjWCX8EI7a/XFW0TiMWyNbZbGDU7gjYvANN78r7d+AmPgM+8AqJyjoxZ+
WJHZd/4zTrHC66hbQQ6K7DnEzQS5pwtXNG7TnZQ3sTP9fsBpcJiZWHoxdh4ItqUVKqUOkQwDA0lz
zX+DUGaYHJkIWFCLFKPN3TB3s2aBGx243t7LNnmF5lUGdJf+MjMCESPb6YKxA0muM1RSHW63h21J
not5OJavowW7dHL0bN3+eGE5bvkENIQym6m8eDZRE1npFAR2qgogGsosbMli5PGrV0dRoGIW3PMN
ASjWrhv6bSSFqj5Jp8uezM0lncqYfiUZKoaEpYT6pi+p1xCh3a2MXvqhNlLGGCJKbT32zLMiVcDW
ZvQDs0xLQtCqBIwvq+0VWCU7KoN5+oHiXWpMMFyONwT7JjktI4xZMIXVjcIn+b8YVm3lZ0oigaq9
AHNh8azwGyqBf34ByfM/1adps0ZoUPTCSRIflulnXI1Sgt2hcquuXCKCH7oqKc0bneDnS0oPtGjo
WX4UnznAU6rtMNQkmX1oXfg1RlvepyqWcC5XrHraCc10IKxxCmy7zvhWAJxskLzCFyCCrrdGCjVu
JQuz4EGdrWWbLybvLZrKgY9H/THtLQZprd98wXOHruGe0hej3+gaProoPYvh6h4uSi4VOUKZpQHv
lCnIIUXCwKcSm33zn8cJxZCelpX0Y+0LOBvLr8/x0cR8B38uB2YVw4prwlBQBgG9lOsVbgGpz2lk
hLJzPXYijLJVHBIWGgB6nXrFK1K/PpC6B28SmuFQBmUkr7wqFkHZi/zIhnhsc9BYvAV50hDSe+Ml
w/REOCDKteSs4TNMz++TZM7MOpGNvBxXCgB0qnormamm3HxejBllMYAOZTX0nJBR+xyfm1PwSRbJ
yyT0+ZBI+ZVKUCOgtHRsVsiUxokSZ5hJwbE6resJ7dNuN1LpQB8rV3S1D7INyPF9igaPb2XetOWI
LeHv5n5FHPo1miLl00mQJ4K+G9z3BPPIDXNqdm3UvUshsjrwEFfLdoihrOf41zwnZT7ZhSksytcq
Pwn2P1Nc9y2lJUGf44z5l7lbhF/A0wkHAm/GonlL6o0jDnOfEVFVWY4APXCqUZQPkxENA2Oxi/C0
QEkuzCYjA9IM0E8J6Hivv2yMmZfb8uiZxpHWeHfnsWrVwmiVr790c09iKWmolAtJiO4+N+qZ4CMv
aEOnuWDaXxvO0m8yu0D0IPMbfJ/XZ/6hXIpPI5AYM4yYiL99kC60HmNmYni61b1jumR5eMzMJKWO
blIyVvp3PcDgPjXkYjsHI/yklikVJ22g73O6w2Y2lIImyzPG0sQsHrT77XZrQnH0MqTpta1bfaWZ
zQN9z9zZ3OQpwd3pmF4wlA4JccR3sJ4WwWniryADWD8izCISBYWHLo+LFtNnc8AdE3sDufIDTHp6
bAqFRSKUrhYSS/0VjYxtbmAomq0nRMK1ecfWh6G+E/fh8seO5xKGU0DlTw7pBAYlzxb37d8MoI79
SHJMH0YXSocTGQsYGpch2WITybAtQuti/7rhOYDL+h+GvxK0aR6T2jSpZKNDW/uH5m6NFhu0J+kh
1sSrXs3MLqW9rr5tGj0F2rd4d9BtvWMYglx4GRxz1l6TgKpGtVaDBci1UDNgpGm1kFDeCKI7P8ye
SYKQ3w2MM3JNs9p9XomuDuGqmJzfPaOq/JmH6/qBT+6M7PqnnizrDn0GFKNJz9Y8szBAU8t+/YS5
EVPqdH1yiLhPAftzs0MjGAnuLg09oUeFenLsYgd9tv6WPWUXjsehaDXHNhgsFqBh47QUUYjlIpSx
vHK+HF2RgFSHKpAXtH7XlOIC0fn3hg2hIipB6TI51UGBmocsCuPJWjhEk4xmqp8Yo7A1LznCWhxM
F+e2iV/bi3cy6Le5A/AXKDljC+BhahWZ5Gss5K481dYePuJ8k5uN6B642TX4QD5qNvWK84xRdppA
fxpBvGYAHgtg0rszyEbh7TzsqHEyQPCrwSW4PsNiE7a/JrGS1t2bAn/bZOmNo8nUaBJKW2a3eYD/
UBlYZWRiYWtST2+2tjDy6JouIOmi4fmQo6XZXNGdV/mti/J/CfehwbJd/mEnExM1+l5GWndE4egV
RU89CdRpGfnYLHOsVdsbrepnjRDsVkVFEsRkztMJy5jsaIqoLmGVuRKVewsdImXGs7LYod3HZ4qm
h9cEXmyCJkZlFszsBhgx9aYYs8o6Ec23EI1F+XmacmsueeREIVOgInQfeXKmzMKV0IM41NDzQPwF
xdOKCNwjNOeT265lCgyahMnv2diVbbEO0CzgV0M0TnDEu+KTQivKTCfrNdhbfFjNqKMqiTJn/mGy
pTBR9GWUcH7POUWW4CruuglMQJnQ7dDDBHuNXz+I08RQQDHCnrso55ha02bSteMy5fHcdEHKPwc9
2Z/00iKzsFnJzetps3Rpc3qel/nUEbHnCTlpk2EyxlFUad2oFkXaTJmrIgzlYCht3+nIUFlXpzEL
xs7QgMcB9coC5ZdnC2LVe2jJkHaFQURWEgDCx38N/96VjUTHzCKDZqxIyO2VZYHI8OAWHKmr5LH/
E/Ny05To7pB1jtzgIFEs1pkfTq4rILeakgvoSZoKLLl/Mo5u1fUMjWuZ1l/pGj3oweShgCC3uh6n
/0IzaZXjqTBfCIon71jJRF/sAP12JR4AeTiQkbJA/5QSbNJiPybyDYOLzKzW26bfcG6ZqSP4mB/P
pXUmSbEAug07Sgkz7nsqYPYbN7eGb7B2NyN8lBJG1/rup/xBz4TNCCl0IioxeMe6bb1VM8rehZNf
JwUOFwNM9z1q5OGZNcp45+o2LVae996DVmi4uLfyWU+iLjIIaS23MCgsseOPo8Wd41/9OjbyDuvF
1oewVE3yHM4o9AxuR8RpoG7BobVT/aqIYDKDaq+hccrWM6w4Rm1v0a28zDSajia48W+jZZoj/kTg
g18VZzIlqorFCnhXEV1n+eDN2++aCYe6+9XjT+uht0qtufx3rThtyM2GphKVXTJPJ1FjKAFdqLEs
xnsmGB0u/NI0HAxf0wEh/lYwkQL+jArq7LhU1CxJT9IQljVkfcv0a6Nb6DJy13JYi149muNpTUGw
vBzbVozrwqQYi1FCSwHhirwVePGIrez26vOApK1nKRGv+1W4ZlgvdWBN/dFr8k6bsBB5OWPr+TER
sIFNnyywkRAe4D/w+NDfq/p2TYNoRlEX6eUAoUL/rc7szGrvqJAJ8V6RQvd0HUDn57A15WzKTE8e
37JiGNgSIpGusZhkvtKbL+XUtUOl4cJtH+tKLioYSHJdQCp5wtWL/M6Goo9kyotEbQ5wLK4HF+uh
bQwaSk+5dEs/5BARyWOjL8KcRxnGh6OXJ6B9jaVQFtwTmpm8MsmTBD39pmsoD/kHQVs/xznkPdNB
dkInsWjuojxwiOVqiTGuULTom8chuen8DR/zVLmM7/IbxyQp4dKOvkx0hVylhvNEirv6aY/SJL7q
1d84ByKQr1D4dEnT3Gs3q1DegjG/CKO2CpUazDl00Sebv+wFbmm5kwZQBCYH/cHeyx8LFnd4Tcs1
I7+0m17H4nTRTZbUtVx1nUNvpGW0mgo1iBeHmAsQApf5WbyirF2HBQqX8M8FTm4mqisXVntmXZw3
Jiy8S8eiRxKTzjs96LJUXw7nmpvACcO5j/RaaX9QzkhOduzqSQQi8ROA5ozL61OMlgDsBHZyqtXw
uTOgmjfJKv8aTz8z1cZ3MyhBSWATW6GQbZogzLvZj6jWWnplYdwR2/xyBaJ0tyvAJQ/QTCAqjetW
kKlu1VvfF3dtiMMiij25kENCA5bQEo5a/q12/k6wdB/bd/m1xqNHxFsh/61vbVLQs7FGLli3RjDr
loPhWlP/VJAkalmj+v/Xl3kE2vgaVnHahHhJyo9dG+DF4TTBNVSEB9t1I4CZFMcklc4j3ZllPA86
wndlAaqGB7tOwSVw+1TkJ1hKatGCNvEU63eaPvEpAsybjBaEcdn/shVbO+7QULymURxS1jtAisp3
ZpaOcLNq1mmHi2GGXj62e2NHU5znhftEg4jTmBEVlnicYm6awEbwGXCnleham2YhApTyCCnCiG/P
BJz5RuMK95j8grcW/RQWKIki3vVMuYRXcuonfVZNkRadsYKYRKYkTZ5pk9S4ZcLIIvtiWRjJbnsF
YhfEiyJlsCgEGMLl45kc2EktNpracPDCxHkM5FqDZJiaiVGw76v0jjqo1k6dzIqosh6jjdQUUWku
uf6G81bKzy6xJlCR4gqvjrsCWla1kJyBjrEm6BgAl5pTVWyMfHnvv7TbtXmXehv9mCzVKGm1k4F1
7+D7lJQ6OP23OqpxGEPWzKkOcI9YtyhOnXPAekYOmFkr0feObW/FdKDxja/RPaMgmr2zftl0799p
sVZl3R5bsEkW3XaxVqBg7SrPeowzbHHZvO6A8dFw+7lxKgalUptpfFcyTwJmbZDnY9DI8RHNuecT
OaAxBTyxcQh2wcBYHl3wq+eQR/qg48J1pFJu59mlKLB5uMYQ9dfDX+a7U62hTd2+3DdVb/DXUHeS
AReEa670OMocKtw1rAGwc7/R8W9FxPXaDC0Bv+SLTl5cKxgb0zEAhA2UlYEqeHeC1k5jeZZeFkyD
aX442FxKItBlROiXLDXK93uJYj8KQ8ln7ZHfhxmG0j1KpQFf/APjiU75meBloo4M26ITJy/0XFat
nLvbJaHpGdrnL3CLNDJQa0cmOfvc2xi9PFVVIszTLzvTvdMOAxewTjkHWX7YKWwpD8pm2sOKlDKD
2rfRkNExBqFTsvDbJEiXxgcM9HlGQ2K8n8jKPExUdY4QckGBLKpeujk8Y3dy3mJOP/QBw4DjGYNR
mMgLPya0N6N+3JVx6mTWhiPLGKldgFTmDrbcanDCVRtoy8SSc+Tz+NXyrtDrvi5b2zY0c3/P8Eln
naxbAjnA5U8zIyEVdneVmZNB3vU2rRFeHrtWsaweNAI8GARhF3IqCqVf58G8TjCuJS97tjRABbmf
SZ/9thbUKscHB2IJo7OMcfKOjgBcNNVnq3huTS35n2aj7VzkBW50abaG1cuepMU4zmoxG+JORECn
nCaHlnRtvkD52ZLXH10u9AUwQGusN24c3lJWByg/CkTw9IuR4uYixMDBV+h4XZz17Sy+4NKFww0G
wvdNcZdBNFqjYYv7xbpHygXy2qppLHJdedvbUjzHzXtfOqucFflhTJMCwca9Z3e2yg9sEwU1n94u
2QydPZs2u/2o3AJZ+e/0BsOEmrI9hIXLI88vaAiwjpHJ27aNIDF9pe64sYTT4Yzfj5ZDYZVu+BNg
4vrtk+RkKXQ5TS+46jjwLb5rRqWLKJ7fcn6sFDopjhvgtLU+w3z9tPE37FDyENDFm2Y0y3kDJ+qe
UdWmYP2jPC+31Ivdhm+jyyDH2/M/WQMCkeL3CcTfi8vgakzcEcGyRPoAjG91I/4fWxprZQ79MwOb
0ZmKbPaXt75yZPvLS0J7+nYJJOm1h+B3Gm/J9Wk4cBR8a05BeKaVuC0oKr6rS4okAqZ780sbmFet
FqOdBQ1b2FIqRqQv0v0Ij0vLtVGoemvvSsiAkBejkxIIiIJk00IQSRQWXbJd9F5Sk4WfAN9CvI/9
4fXdQcuUzQF07BSAFc3gOWaLiNg47gqaGizLE4bvD8caEtnaXytzSsPRt6e0RcyZcG39lYDuGbzT
m7Fr783mC10MQRIBKeOt6R3JeMOaphw2Vs8YsUtSj8ao2vohdiwwBEeoHgJiOQxfFF9t5klpn70e
ot9Af9FjTBmg7q7rRsyWLDhdqySiWG309FHTUrYN/wqQzyIJvfSMXr3owZPiwXYnMNMYAGarIQPD
ik8HmrA8vqmeRD6gFxvAEVCQg6A18hp5kbcIMfM2lj/EP5kHhftUXSRh1Z9N6tLeyB2uGxd9S23C
KO9zRFalxO63H8z4hn5G3tJTjAFpElNB7mrr6d7F6KzDEvR0dBWkrZhLdOq8++aZrqn97BgalAaS
ULFR8OX4tpylZG6xVmHLLdYm3ffUp4cFdprK8lDIlA6GTsZ8aQYqmeM1tYOVZ8tJ/9FmkOgCxAKa
ds3ag52JfhgOZBYkxQphWjJBYezMYbYVPCn6XOkAB0f0FoTTRV94V+viv6Xx0m97zoafOn7kQg2A
fG/Lpa4mC2vVd/G3nRU6XcrzzfkkPRpcU7ruQRbC0oAlWJx1un40Wt4OHKVkjv2yKZwVunkiTLKu
WeF/SHCJA8gJQA8bR1uRXadk2D+F52Nd4o3TxExwxG/4bGSPQZmFuCKM7Sr+CK/k5AwegeToGbkp
xMQZcXqIqH9mUHe1XkG8dC+y9N/12Wyr0INV2utCg3THM584ipflakY/XOybY5MmrudN7LMr0rq2
ACryOavTkahkuXdgKSX5NzHABHZx4FCI3nQsP3+wIoRMzpuOHe02N0ZIhSpORiXxixMSfOafQcsb
hLtKKRaZeuVyW/d/JrVFG64EIPhKQ3aNLb792QFmV7HWHemAPue5ZmW+mNVsEro71j5x5uFLM/zp
+Bd68UsYimmcYq/6xiNzvzH10iAFYteMgjg+ObMGF6ctautBnZ+nuX6pO+Xf3goy3Jn6uZNMxg+y
qL3/9jwCw9Sh7YAChrvVnlyI72prF+ilvJDAyv7VRr7sWsd88/A50vzGDGKxtOteezan1tYkC8ub
JjnOnN60iJeqnDy42diPlJ1wp9meMqGAM5fndxha/m1TY7n52ANWH3ReX+yEFhlJr62uVKE5Po7I
7LW0pib1RwUczupysV7pEaUr+s6k2v3hWu5eAEXqDx0K2dbzNYIO4lskQ3+Au4QBND7yGQZzFcMz
iRTFPzXMugQbMVdBpEaGh/U6aOeWwBTlCYFtYrHwXn6YdYYPOQZcdJzx1EYisY3HtMTYH9bNQnwh
Zq1o+Sbd/IznWkuJaCxV1vJ9T+jTWATcyNJyzVPKX1ca0jtfgVSgvNXmAe5VwTcb1/BYk5vFwSYo
/7c01ZFm5ZlQXISsQGU2mZ1MbXLHWGz9GJIRBphuTVCTC/IUwDYK7Tn14Af0qnFNe0e17EPnilBn
x1I5F2gJr2sCtYxFS58YSyM1IOFReY3IHMC4lgIJ+J7uBg02ybUuU5jR07FxPwVe4HT9f4keQoRI
O67rIorkZwCvuldZDj28JRqpH9HdkxsHjkt2uSawQnoYLH7j/YP3Boj0MYqFiE3QhJQhyjfElhRz
jnOO3p6LfjS8z2hWdLdiksQvH/81/hx/szloXOLhSrdsM+6E1/aWrv8zHKf5CJAVWeQIkcFQnfe4
yiu8XwbdKRenC0CSG/PuNGyI3BgUN6xzvZxW0jp2I+t5Y/zjmYY62Ll+Mq6CkxnYbcBhEtvKfBxY
99+Ik1frzzwa8wLZGR+sHi6/RAUhqfPkDVSZYCQ7ywTeH+Jbxzl1vsBNWjgjvozwz8ZR6tbUHjvC
3axrtvL/ji7SWxaVYKGTQxgdIgez4x+marxOkVT3WyHEKUjYgZUBK8otj/I0S6ffTkCQKuo9CUG2
92mH5SdVZAiUsnVa91itFu0gdkj04sXO4y6G5IyZs4RpDbdtO6CkLdS7uoajbJBE2Et5hJPLJiAc
aRY94rLlSlYeWhQUALqgQkpjOQsl5tYavIIOCS9ulPDtNzFTwSu/Fa8stUeL8qRiK+pvtYMJbapb
ItD/a0JyUaJ17aMuXodKF/esn8scFOXpEfn2nXBgn9XZOxbfLFZO357Z+Gje6/OSgwONdwIv85Rw
sQYxreX6B5Tv+3/i6GVBMBwhjS/YPEHQjqs6TLUXPeFecpWJLGysd12Vsw4GAbj57ib2HqvRQVqF
RCiVZ3ErmumxCTNk4D0MWtMm/GuCOZAI+CxXB+STHqJRkZWeYpilBGjwFDHQ9IOpWyqTbfLGf1Bh
Omv39sQ4AEyPgFwOfE4/04I63uU+w1GLTaAsRtS9p/SPiXtjdEzkuaY8sKtXwBjvTv4WcoVriFt5
5O8qToMj7aLw58dzJAR+BvefvHN0yVwfg2GVS8itdVCpmUcBZ2pq5+zQ18pCoy3fBSGOAOwe7PxE
nzwWu46AiOC63fcU6GcGezSk6e01d4svZEBvOVFZF34JJp2HYl8nWDjH1zXSqj6aqYv4JfX4Vlyw
U0voiVyC3IwSZsKQbXq5DsbTC4uJMFA37UQb3lO77hgX6YuCNlremaMOoi0Q+569V7CIuePJ7GUh
jmxmkh1Gx0LyvLZUGG3v/2ZyxYIX81pCe8YKtaSBgrx00BSkuiasRVeLNzwzSjLyCB5e52mxW/tl
IaYP1GGDwnPFBACb9k/+WoCNQPZAQ7cJt1OlEsgV30pAKjTMSe2CA7S+4VFdeDil+nxB42c9rZaY
O/ODEwUN0NxuAIte2KjgJ3b5B1xYj+lWDvxKorVItqCvororQIXWCAOoTPsK46wspk25WliAoleX
WxH1UMnVeLv3MmVp7rVqQi151hbxzDkU78gOSSZlwOgY5G4I5HpC/nsJBw/7wY/43jxuIJrGrM1z
mBWpOdyTu912Dk3J1tBKoceaP/DR4KtTguoHtTDDlgd4PIwz7qvsm03HAstkQ+5tU9TtXiEdZZPc
XcQrNSjOV2DJhhTjBpz3/ANSmO8cG21PFnx82UICcAn8Z/KdOrJ3z/T4pQ2Dfx9oD3NfpP7S+oNE
RDlMT+4nDP/skZzjhTqu/a0ZghiuaoN1Cuav0v9csXdYrwRNej5Zllg7se4YoTI5IZSO5Rvk8JRB
OyJIA7qbAoWS12T5qlf9kf4sHnESYDycgNMZeRmHzuX/fTcT7J9s0WLyRYmBQpF9bESvLuaUxNBa
1gTtWaax6ivA7frACUgUCTmceD4t9Z8MjDUhjG6VF2tVzqVn2d+dl8cBoDT/wvbuUlBNkdu4U/Yd
k5lbHgJKfd790OLpcQQqO3zul7PN7JLpKmVW98IU488p9vmKQvIEvsEU9GbAro1LjDQKerTbnIwa
3dqo2URWEx0aXaQ7hwQx5JAhvH1KPaUE5wsvTn1SbpWroIgBH1BDufpeCqflIcih5gt1OLPRNDw5
VdXPveWdFWwwhWjyr/3KSDrpdDEv2XjSf5jWRnNyTeRBvgehdebgKDlohkgwx4U3APLBWEFGUugB
dQrNIu+qQrl74/gdGFjS4Fn42+DoZ+dXLfrnNq8jIS4salUEtnwJrvr/rXvLfGq6eEUjH4I2gUNx
HTGwzvWyoPX2OOLpzFzPfyjC31JHiDNJqfh2mE7AnI9ighog03rqizouGqROc5NIs775/LyNAtHE
7tBb/AI6Zq10RQa+uevErzZsH0qdF+HMPgh4J1OXewfnu2mvuwov8cCGom0PltFg6fHX+2b+9Ols
HwzGQjCubk7ShxTw1yhSPhL5iIwPRy34fbLPkZrCuaFqmaNoU4p6h0pOAWRs411nNGcoo7zq8QTm
vMpHh8NcrQydnPQ0WeFWoWTqHooOAxhE1PgT9FvONECC7Lg9vW0Vtj3B+yvOZ5kn1Sxt8GD6iHrD
bUjWXW6ofnTYfifyD7ElatH9/kcpAMqX/DCeF1lTpXKCjq8vAa4Dp34WiXjb8pFpc7bbvwHgL0PY
YMof5uJdWuzkNZe+CudMZzApxQYy3tANc3P0+24dziZFb1JhYtcmMB+veiGo7WOOlPGVIaG2rk7B
GaX2Pxi1i3dHo0hCWRVMs3xOK2uaECkwfv8/DrKOXpIdOtgp9XlBO5aVBenUkfExW57Qk+gPEFjC
3ghhOOqe04vFCeY3gGI9e0PYK40wvn2QldLGYgzOT31OKewSNqfXLC+ioKBvtBxnbzPJvbkTVGsc
yemesG3UCOOXOHDRiCjTfsRkCVzx7rVt/gHZFK2Ep1yHfIAX/ABZV9VHK4YmrJSdVzHblCVcfgh+
B89wT3U1FzMMT/IH8e91s7N8sGQs+reexR86imMvuSKLXQwgvi4GciO7HD5ZL/EvoJuEvZrnqzFH
i1ZN6Y5tNkd8vv/dPaADDS7xurg1tknoR4s576t8ExD6TYiiJJanhiOz/zWGuAv7ngtT86AZ8COD
h3oRsUUIrgxXM2oPbzXv88ilpMNeasOJpkq+QBn6rC/e1Ik/Jropk8O4/isAuOwFoT/CGAvVGpaG
RzLJ3WArSBH+ljXnbXf/NHVRZOwjYQE7ee1VP5DGrTXfIPLJX/Ov2tqsnGlljKXE5e1kr09q9QAU
KAKggeq+D782isrqdh8p05Sg3aflq6+0/y/E0yMwBCy9VMztfXvwUhZLVhachwkeBxWT02yfZNeC
urrJJQ+JbtbxxOuMrzKwuOurh0P2MLVdJCo2scw3GQRj4lSYy+0OFsaSzbfryMtkGohaKMemBzuR
41tMkqJlO9REHji/pyzJ1W/1YVDmqAsIlQ8uRHLXdie/octZ7WjR6VKhzFBITfp1Hxtxyt5KecE4
FMJiazFC/9lHXNpdEhjGaKr+5GWR+OaCI23PTIqBzUg9utbMCFKmqRWghdwBEcz8QhehG7EXqUSE
PSzpN2zZIMcXYnM1DshLdn55msZ/HPlwQzyFEvyJysovVlwKdbd3jxs48CpCCo/DMWdPw5HLVb7s
IKw605tMIwXOsE7VJv51TCPm02RtzwJSLyFtT9Zac8REBGiNFpcTjdfD/Ux8tmuVKo297QbaxpxP
cvzTTcVOqnoBOwWp89FofH2TgMZV+edYQwu2shHqm0mMNaW5YhVdFJyxLzXLWl+RU2hL9MSDW6do
S2ySdqqqTYU17mEoGB/iXVpGDnQTxnnkrXGvrLXuayIvgqaycHTZyGKr5RjOE+PZR2XPACIDGsWM
6KRrPCKT4aF5hTJWFzz74XaAz+xkCNF1L3IwqFW8UUiA4uaOcXjD03YLMutmD5CXtgT4YOILRi58
eCOHhhTRpdOpopooeNaYHmUwNhuBe6q+mT02ZyeuDj5qMKdYXlXQNeLpZYDomJ7+j/8ueM/I7rSB
k2Kd65c3NG3tetju90Jhc0Dk76yUKGx5VD4NcWnjhyC06h1HchpDZhVACWQdVtKnBFMBTDBm0NYn
SYAEvZOwFrhRC0wK1CwuJB2mONlp+Hi/LF5ziq2Aa5Wo3PB2pfUwa3PORftZERha0jCjtSBIL22B
t5N6qJGeKwoLs3DhToW2YZuH5QKfCltJhLzfG9SQK2qmwHqtx1RWXxXOKJ2OAI/sNv67OuTrPyTl
UEhRwm1WM3uJCBYGJ3130up/EO0DfBBvaV0SUBImSHQZeEbKV1GZ+465E/vIgGerFAiQcgs9P5F5
2S9eAwOUCVKFo6flihGxiZSq3H9+11DnD+IQPLXYnB22K3JPwvQJGDCG6/86qUZeMbA0pGNSNWEM
Zg4dhGogIUHib6mfn++dXjoowq0YHBl0ORMnwFebuVWZfngUjt33D2UAKkLIKvPbeb/ZztKwydr0
YGzYItv9R3L8suGMejaL97Vyz+X+HZudVA2UOy5Nqw+1qt2ws13Qbtyx/KZhDywW6vW0bIXJzkI4
rpcnYVOYRbhLiNPRSI5tN9pX7s2y7ysWLusnYYgXfPYrvDb+kB2eCK3AbfCNEEpP/5rV4MPEQ8hK
lOBca0+v5UXSadj7ofY3euuc5xu7vsiZbeLiicfrQ3T1h+dhsH62jQGGpWFOyiXnTwWyT02JW5tr
l5j+Ts53/gWizD+LxMqBeOJsLsVdGv4j2U0IoT/Jm5z+bKDkJK3mE0l++xiFchQjLlaCKy3pkik4
hBqUBwcLIpV1fNXeyn8FhpVaCRAdwbWc90dC5Y2XJa2EWNV2pGm9uZZjiZBihxj2ly4sAWBoLlEu
361nsM1Btz02QaCxAjpqF4Bi6vI9p7B/dTdctkENMFhafc1Jr9vl+9j+RM3UwJH1tRkg5vnkpGsU
DWxsPNQbZ2VbVRi6N6THu2o+cTZD67wlXfXxOMsVaeRBxpIfHmn29FCTHVM2NlyQFLaACFdKtLs/
TUDqaraRzktDjel7W5aVd2cuDoYAjGxBQgUnUw+qdocgumxqofbGa2IabJrc2BsWo3450lLMPBB5
8209pdc9N4cVVv8b6jGmHlp2rA+6uN63AI0rLCIx28WROWry3PBH4HublQuQGasp8auRNvlQM7d4
/rCrhLCaT6WAaOKNDSRz/NpcOP97iMrhi3Dn2Vg8Jf97hcWQ8aVXvI3IyQMQH4m9fqWVqXnMlm17
I+d541Nq+uM1W/wyV6bv9hX87mwTUuEJ6RCkloueG3HU5twg/LWr89LWCNMHqv6eXAdL9XPvv7sT
Ud2kBC7sMa6Xani9shkgkm8kXwkCce18r6ynmwBdZmB46SW4O/OBa18zNXvoPg4MGRDSrGhgndv4
S1igxjhtQ14nJ64xqBgCRtrTM1RugbyN9pvx47fZehq0G8FTpbCedJfDqqe9xWZRIGjEZ4lKQkrj
jymvloXgiN8QUag69MHGsw+bLzizfopJue+1cEcq2zn8gaRfqBCxkwO5GzP1aGaxHnWPHrrn+8lf
KErYLtlE9HcwE/Vd2WErx+KmgvajDoSoCkTw8LrbvuUp3idnywow+1CTfcY2ITr/IegVbGkeK5YV
LwhVwpjWJsrF2F2mENEzXmFWQHas02/SP7v/sZBRLGgG+ltt7PhGZKnygeKBNNznIoM0Htx7FZsc
73zbgsbz10N07odaGRxnIjntW6jA7TpF6vteS0XZAUR4GPjLYMq1YMr6lZcVnDApsvsU846otV2n
/vnF6VlmlfkAfoZXbpyXqxE+O2+N+33SU/SZrMZn98rw9ois9U2jHdOqBnD3LlcqaKEOfZI6QXqo
zvqGOKq8M6IikmMHogB1wx1kNCQaN0wkTGPOqZOCbmx+th3P/A9TA8m9KbK8kqbHdHZ7WlcitR1l
jPVZLbgPmnVulm2SyZZzMrZpMMHR5Gz+7dgoUCeJ2FNZvmKXbCWmjAN36SWq9ynt3vA33w9kxbAO
cHEULWo8d/80CgCgS54hw2WcdWIvTeQqR+bSL7gTvzPuYvidMs6rBl01PFb+TYsKScytoYiTZFyo
1V2/eSSG63rOK2tI1Va8yfSTVwNdazLKGyoGNaGdI5WRIGi79/sXgiELrHZmBzA8nWSPTRFsMl7c
/CDGqPojCAKYqQoBXAIqexKr+oqRIOccdpfvZByBVVQPcXJ6uFOEHrTRBs+pvxorqO/2ZiD1O/wa
h4JYuV6x/yLgqwunsRMkAufCOT9diUCYsZxv+lq3+SaCstpzk/LnNVqAnyYZ4NO51fIt97POqN3t
+IsKy4dv76LDcBTjg0mRaW5WsUAZAIo+UgzGN7eoo58y8GDNAAtdQWgrAKpUpLgsvfe87nhIZSaF
eWMPt5e6QqqGgUKppY/BVLIfLqdkY67HdZ0BIYvLe8+HvZsXI+2bAp4WkPN3hAlhtshmQSNeteWl
D9OQBCiieFshsasL5FSw+M32MtUIqtLs1p48P8ZUaK/wpNRsRhiESGu3xmCHBpdnCQJAiS5IBrxD
2m2jhwvkBQeQ4ZvGP2/6nL7JWP+7NIObrwF/ojqHvHb3WsQeNsHxEUadaCVXdboOUziHEMUJid7e
XSwA+1pB1s+LmecAyMRNApxaaoR5cXOoLu/vj6ScrYx+4FD+pCWGJl/iP/+Al2jgs2OSN5+MyNjm
mOY+i8Gbkqawu6LatT2U+rv+wlvwmnjW5bPhffJElC2gK6BIU6RhODFlHdxboBgsnX1lesEZs7zL
MHKCeB2NauRM0Fl1QWNvXWSHbldU+NR+rLPqQgSwJWkwlW+KCjGcHExOTVwIPFizRn8vs7GUeOhF
/V7bTwijHRWIrC4syo7ouL0zORypXeAeTPsYj16Ehxy4VTkRLD6clHVfrEz71iWr6eG+W7CPS/hJ
wHgMcypk5YuMrkB3ak6L/mf40Aw9Uljxfr3/nKtQv5tqNK+s2ofDgBbXuFQJ9aNyi3WXvv2jPaiN
IbFa8gabXaKGDFHlbT9HL4uDvwELhCckdR6dJ8rd++byF1dgI49ozvgl/7ybJChMWEOL2Yzxm+mm
UxEcBxR6LDMJnNdLkiJ+ghWAb+/z4W6pdpIiKuTbuntwV17uFZs1LwZ97VATjOFSoKjnt6U+qnuR
FcJuutGMnuu4me6hO+S8fxyfx5LhZ56rwDw7X1/Qu8F611CdIkbE8RGZO7F926bm6DhhgHnP13ok
5YVVwf+stc/1hzFrwOPCKCZUIXC0PaxAkExT7VX9+Y9TWOkxaZmbJj4Vq2WoYaqVsd7+BhhujkID
XGAfCCRQtd/uAMyQZZSqKxVQjHZ6jwyhJnlQzp3AA4vfb0avpqiijUYBKm1wVSFwJW8cm72yxar6
nZs5lS0mAwnBo5gVr/ouXfvaqHaZH4qgIaJkhiV+Ur5Oad0nvIlYi+0WKvN6Qd1uNbFxiA6gaHrk
EiEYrXufNQDTldx+e9szm1cDA7XUtQHPjqVjNPR19jfySJuNF5nOdfk3k2ulDN63v+FKRgkznnHM
VqohdcYVjDpVPT9E4+PFYazsJBJA819i36JaHWhtWKoE9LdrFj/V//Cc7+Gi8auJTXXA/PP4hvvf
hE1mDhtsw7IE9i6ZxTAfR1ajawz/UMZGUsryE07rDQLqzu1y2Ic/Bba7Qmp4MtefjqrRE+wc/4c2
0SwR3Jf8D3+qsa//NL08RNXCdG50G0Eyatwc1zQANH4P+UQfNfhkRUvcx9Gkvr1UHgxbJJj7yBqz
rS6/17nL84DuvI/Foh1vckX3kHV8WTEKLlPWX0XPm0lW4r2SxPltZKTSXtni9HbEhE1Nk2Pz2VPS
HE8Q6o+Jyf89nT3/8NLSGwgdWtvKCD+b5szuCgn+4ryTOHzWGNpEzZh2T0stFCYbcY01H6bo1FUo
xXneqCrqIj/w5ZDTYKiX2N9FRm2QJcnU5wLFvve1nwqOags3iN7TiCjQRO7L84+HTMKMv59fivhN
ydM5WXK4VJ8ATPFa/TfowpiLHuTH/zWf5ek8hGnCnF5K/pwDtdWKT29oeDm2cF+7CUnrdPbTwf0W
qidfJ2Cdo/7yQnoUXpGckbU3gNpxv4J4OI5vYsSzMOCV1iDcG8wK95ijuO24ryf+yj9K+B0gU7w2
X5PKfj+fo/bNgpNT+DhfiDHY/XvvC2AvWxDiXv5eYNCbr18YfKY/CKXVfF0/rtr/sz+Z1tEZzlF6
V651aRWfIsONjTnapA3V9CHtIrrfQrsfeCDBEoPYTe5cZsUxVvN1Rvi3ZcuC4Acya7nIW4AA60jl
CZrPZD4d1qzO2JD+450G1KlaMorsdiXY5eK3H4r8DkGYiu73EvRQwrMjUk5DGtI8thZYnvYGex+I
c9mNXkSUgsxdcfTteUIDBIC0zgHOJSUezpGO5DKmUy6MyKJGQza0Uhk26Cs68MqhIkzLpOV9Q6wZ
Vj70YDP20J4ukM+shJzGM19ECBYW2bdqDyFXQzrgaqblKRMo67RzyReopKflO591pEdzIW9EMYaw
BGPWwt9qYwBUxUZFWCJPPw+j9K9nMhgQnHNqnCEi1lEv01rCe63NSWx/nJiw62pfsdIav29yBr/3
1NIfKXXqEx9fr2dMohJ1iWsqTw+V6/tzmKUkMGinxy6JDk6WPw6sVKfg5HLnodkvF7MukbekoV/E
3MdLrX2Vsa58GT2tJfaI2GOE3T4D+djmCJmFVpipVOq7dcas7XB4alyGKDvX+mqFUjN/prTDBqFt
gnf6+appPDFlfXCbxWCtinJvTZGM0ji6KXoYh+cVlIyZ/1Z33oLWY9vzTNVww9NpC5breafagKKA
SNpfbU/WFNwzO1IplubPHSw2Op+L1FABQUfa+CEpz5H0Kdp3KItPXP04GrxIsX87t1rrhyB4VVCS
Q080Z+6NZdaELRSSBVLyAihsi+s7MZvi/vLjNefPry6rd+yN/krw0YW2o1MYHnwl72JjQgXfmqzC
rbjURf2IiVORZQ6UQLhNouiQUHON3JNsqXY173IhGC5iG45cW9urBNp01297RxqL7yV0WOrWhOh0
nglnoutKYgqyAVT0REn985ZAVZHBETjp2nS34Oib9JSwtz/Ai5btcAeZjz3oeJ/8auYNf6cj/8sT
iony/txH0PA7nh5a3Vgle4G3Hom2a3QpaAWiEWe06nM78mjywbG5Ff3ua63K66AAq8YaX/KwUkjK
ECw5M0gr8ZijIMs2JI7Yi6bMd++0uqvmjBhuNj/EDDZ7B97RF7lasO6Ht9dP0V+4rnuITTyCyyfy
7YkvK1YNcY2xySPQyN1dqCGLHqgIbnyELPqXw+9o+5lyzgAsiySgUAKID3R7C5NzqyQ1LYR2Oj0W
QbTuN8X5Pi0lJ+DA0ELvKAXfBzGxs7+qLrGBkcjbFaCBQxp7LfbQKQqW9O6+2WTWUBmi1gzYmhrx
2CQuKNgZlwWMzt8itYCm3Ni4ZfXPYuPLrKs1Bawk0wywQwqzocMWEgL/mAGT0q3U6w1bNR/y+Rzi
fpULfyJM80FIJmKF0U5fTH8SjfsTLIi4WMjAGhO0rrf5Q6EnMrY+A4wXni4zdrn+YzXj+LDA9sFa
O3pgVqgrRp+NsXr0wkH+FqT5ASYs1/KUKCd5C2sq+G1kmcU4+em7yDNiHikVAO1i9EVsrVN1D5sP
jFgFjYoHVL34qxpnAwUMlHllTd3Wr1HzmJ6DH5DYaIlmvkjRR6MOHHHm/Q9hcq/q3hKV62/jt2Q7
V0ekKWQLPLvrZx565gAcdTlG4CnNeX96ig6V9Z6OQkYd9RrlBoSu3Tsn0AVHKqMpZNRXSZPHMGKZ
VSAOekJyuW04wzygqp0qL04MFaWOxS4YzTn9ON6hmZxxNOGNvCAHQKb/e0TLt6RAWxrY3pWRLC8/
d9wW6nD+aK/9rQ6LtVuOSvroEexZrhXR0cL/T4JLpWhFcOQk7Gv4rXw+8nUETHku0cHoe76jg9Gm
WTAH5rI69QLe1qDTTfZXxlA1pybxbuZPwftQFMMDf94UkYELDMtXlfSBn/VUy8mXUYq4Gw901I+E
ZohkGvNTR/pVWbNLU4SxxzIsFnBWouQJ7SdcjpLRyk2xo/WDddPDfKhRWgh1jW+vagg+bYQe5FBd
QYmyAmm2E9ULA4ZrLtuGTGBE8oHskRgtYJI95S8TDYu6UPWx3I/gY0n9QUrLvuzy1Z3mm4HG2KVZ
RpqpPPxTm8K3xIyCAr8nTPDxDRp8uY9dRTuGsLZuOzjD7JNBy023peVWueWr1VxEtERrLVcDNWBu
VxlwVUUjmGDkAvAGwm5mJvrpXNyvYgREQRZp/72eTTi0z8vjGqrhGs8jQ9ySMIZbIozuOQzCIZIC
67XkAMURmx87bwCOM5G9H5o+upnFOjPc16xdADYBA4+4jdTcB7SS5SYFHgsrWmiLbOksRM8Bqd22
i5/uDD30p/KzgoUkTq6dAAnSIE47szRRtGTJYQ/8gw5C/Qqxq88JFdBd2FLoku33270MwBUPWq+H
5pRhwTphLo9HtzcIEk805A+OWpfyNFSBo18kqDbExAuCxv7S3amxX8PF4aaAWZ8RE/ZFmJRZj4fk
ktYRyG94aEpfJKtwGZ4rT2zRHvOj96yiZlrWWUs+VFR14OW7aGt0sYGYpiKCFvXpLmYNcVra/TcS
jG6d/IdWhwF7u9l+BuGSOjOwTFfv1gvzmFna6Y5htpgSOi8+bTLPeYKFNEIg7Ve1RBU5lgXG82kr
tZ59isBjzcwCaVQniKH+FzQYC4qpNCZdXcpW3c1wNIRUp7cpvOGaEn2Dwq7dPcWt2CCgKV1jmo0H
2T6rFX05mInx8I862X8Sj4tpFdsS1dTbKKzJ/IxBQUx45j2PnzAaVpEky8SitZKWIRjlFN7ntgon
8n69PHU2P3TjcopIY09SfZPGC9AbcyI8t6LXFciDlODoQo5Jr65ZjaVBvTY0saKpQQgLfr3WzFJk
I7eIWdMK0Dwpri1PUqSy7BBeaJDb1CX5wWeJxmaM5Y0Io9G0r7ExKl4xiLN1GESH64Qt+Lb04NJ1
kJhgVzgFFjBp/cbROz5CcIHapxAleVt0kcZ/DjxOx6ZVey7r7sSEHv9CYjNCG/hHJ4IJClwqxwb+
ASCfUoq6U8VsXoujqAhaR5QmFfjo7fehwNHRvAC7+FWiMo2bn0UQTbPEngx5G8eUGOVGAcIZBTyH
eDwP3w3iPhehhLfuZPUymL7fbHxjEge+IFGUizURpQ+Ah3zY/Kta/S8EpP81YX8OBA8zUf6nQAxl
Ydpd6K/aKeOnOVdu77cW2M92Gl/UaYSq85JFYv8+SqHq7z59PqlADYMkYjI6kSCRGh1HUEQ8hhau
XjFkNni4pc/TESgQu6k93/n7bX38/taENy+I7Rz6BJxUjZCypuRmtfFKpWr9t/7VVmSyzV9+xT7u
EHRPFxGnmBd33/jB80cP01ByXsfBsobDkq1NK7IY0DR2eh/+jcb+vD4j08qAqNNH8V84q3GCpogp
ctvg0fLHUMCOyIM6jTqFhW4ML5X85IUMxk8L6zEr9x1ssE/CFHantsL0EkZq6Xp0rOiSp3R6i6vg
uzgmcqN5GAUtqCgkMovg+OXb7gwRF39hwMXAODPWwbExVM9Z6ffs23oEtBiVmuGMfbgbKhqLLHV0
pAQ48/uxeO/F651TeS286dtlZS5A+dlAXijcGUKuNN5prF+UlIGyqJQ36cn6Dx8S26KfyKuT7nRw
3eU6fLVJQAFtA7tF8cj+K8ESNEYLZXsEbGN/y5GtIgTru89fcgoOFVEF6bZIRQLVWAstwsuAPS34
H6K1G7NrNE3OLb0PCDx5L9PwaP784CaOB+iRV7CwjxguS+mA9qj9O5jVwBc326rcpYdDdpCacRG4
sJl03DIe8Tcfm2uWn2tnTUtExaVFoqaA/UhtvvVsjfhfSMLieifMBiw+9JVm+spB0nIiKacd7MZu
jB1kbC14dIY+oQReIWsnuqQOK1H8r4QrCP774nc3W7D6TGfIhbyQJBiWVn4Jb8rfH5HhrjNEQT4s
HbeifkyxI7L9/8EsbAK/P7KSD+zhe+sjPVYZNKAXMjh7LcY8Io+QsWZJ6CFs1bZBvlhOm8fh6SZW
JmBitqTPRXDUzd9HyklrI7VtR4Yi2hRgSTyS1W1cn/7dB5SiwYyXYi/bL5Q4YRS6XWU1igUKH4bU
AexEwkJ7zKfeEdSITGtDhULcTBnF3CGYVVBiDGTIwnJNVv8pLzCekJ15ulmKqqanRs7EzHbY0LXt
rIqNHd4t1OgrXRBc+0r7BH4KKn0DwwUPH4PISiobgVtJAHbSB6s0h8wqCs6eGMsQuGThHMtxybge
EsyVWnqJco0xf9dDhlErP7epBeRIgvLslN0kW2HMW8ucRUj02DiY/xkVR24HU4hyS4vre5Mdpbp2
SmC2jT8eOimnrQHZPHDK+WQpsKIAtA96pBTVYoLHoUvjhfRtzcji2HqGVYP7SFk84dOpIWeXcK1U
cSLqqdDE6XZiLLy89IBklX3Id/1Iv28HVSrFKWhzuKG5Nsq7S8dytkqutqdQGXeujP5UxZ9BG7MF
o2ub68wsO8S0hU2K4XkYHlB9AugrsWcO0YHIq5L12r/3tsIYDphYHDFpG6bMT4RixhSP1LtjXI/H
WrUmerVizqblrzJopw7UDMLIap9obNxNPL5Zq1ttk7SJ3NOF1FTTCGZes5Oj8Opez75R5uYh0spK
ac+K/Tf66pt8XSdI1bHMbOgEg65XVylw+iQmJ30XW5h/TLrbUVN+pKyhM31eR57hmiIkAEgQTFFu
4wcTslJLqy9ChpyGFsvhhoaDLkQNCYSIP0/y3zAgeUIBIxrMV/KRVyacuUhPnC9ieXPrExxDQYFn
ZC8T5+DW0udalG7Mq9rLQmtfYgewuFHM3FHIrCyiMtn6EJ83U9gphSy6XLjhsQ+qWWYiJ5hVnDzI
Yo7ZzG3D82BDw4JEZLuTDoUCFFl2HmzIMpq9aaH9xRTN/8xDw3tlyO2nm9M1S/q4//0rARhIiiOO
Z+cqbqbGHB5RxRrhqlPPxb0d2K2OsiBzvysfr5Cjp1UdJyfGOFoOspnLgPd03ASklmoHcOOZMpr8
daH/SeeC2aKI56yzOKbIaUxntVYnuBUOhEkoa/CF4Wr37iLkfY62S40lk+IgQvqxAYmi5LXptzhI
SgKfPZugNi7iaAOYOuRMGZCFwkQ8f6Gbb8SJ/YiKHY863ih2KL5iEH6bbwlQedXVezGp3MSOWhke
zvVAv93WvORSzG2KZ6PA3bSjyd6jOD3NqmD+n3RCAgjNhxIbo8UPnnzUQLab6Rc4ZqFim22woWoD
TCtKvTud+NrUiSMDKBen5FnRSNtbdOECP9FoWHqHlxsFn0k3JCD5lRp+WEh09bJm6ifxsRA0Sosq
te5DHUFI3mWH0JhV9BKMPp2su4UJqj1ehiGB+juo1TkEIlrwszUcXlNWEU0iczG6otldEMHDOOaG
BIIRhkazXxwIf9qTSW+rhGaFDfAPAuuvrcJM7pMk27wLZUwiNvAY43wcv2eFNE84fXcdwDxy5WmN
8uiPwnfMX2mhzcd7sBZTWI4Avc/kzZ1XC489G0aHivjMB6tuVjWLq/2nN8s59LV9v372T4XiNjOz
OFXeM7XRuFuBZc5HwthHuLWjLEykSiHL+eDWAslnsv+z6/R0gal/zmqA3UM4iS/ALrFODEyt/I3k
vvEwF03rnODxgRaM+js3bOkzI08S5WHn9tszX+HeSdkMTrmzwOFnqHluyfbWIqfoRWrmVIshZ/S6
LGy2y5lafwASlEoWqjTDo/lIxYl52HUYqCbDnB98WhPaioFQ7J7d5uLf02n+RySNg/W63j+Ao9ug
DL/Qtz/lm2bChA+C5HdZTANOcuJIPk7tB53QE02PUjyeTgyr1F25HY4YdukECb50odiu45mhM40n
OWYtZg/W7HbywmgFO1OWs6Fba/1VDEvtQjuWpRr8JXBF9iC0AecUHtY99q4S3OJlzCOiV5oBtrUC
/PW4+/LRR3ciWL/lU4MFQcw6wf9VkQWcee8Fgj2rh7LQJgfHN5+PuMog7pEl1bdHXlt67KqiiNxB
NaIspEWCKWdn7iPrOKpi3FnrMX9bHO4gPzOrLwahsoRXaVa+3kR6Gs4jcu1l8JOcuTVk0l515dVm
SURSp1CFFq7IMqMYlfBO9ik85GJ5Wi6CwOmk+5dTn6PZ5e3Vc1XbeEKwctGFqcDrOVtnaSc1xR1Q
RqxxOebKhjj5ozAvzCVvi0/Ep3bmloJ5UvrbSzGRmQlWPhmN7zYkl1PivRoXW3yIGeKSBJAi45+u
Z2LmK5K3p2xHDJ8ZvhmJwjnUeB9OBhrmccWG1Sam3MbRUGWIxqBAk24dQMesYxlWQX4QhuUOwSCc
DSbYjyyCPzUaOinJD/PvM+NSBEdq/TKBw/C5rgjtLUKMpnZcn9rGwnG2JGi2IQ8mUrVeMj9vUKbz
Wy/EUo7lVd2/wcMgNUCQ3Rq6i4QLKmf3sj3fQMckDGIAJmJGKHKbcas76/3uAj1PVPrw91YTKJ2F
SVTE6iMHGSXiBfPalXpKSykHc+15fr0LfiKLXu+wzv57V1Z+m30FYcG+FBzGePL7o0E6n+sfbbw7
bHgJqfr83NE35r9NTHTiFMjEXvkIfd0XIQsexmAXLnCT2hJeLAZiG2c2YCYtVyZskY8jMv1jH478
sCOWTVTWHtaQivvROZkycKnxhPkqvqskfSouVOgvXZCOks+JHr0Jk6XLtlu4ADh6nlmmByoXBe6D
Yy+SiV9mJi+85Rko0G+U9zmIt8tHExOHEbxck2c2UBzHDE8UfWGT6EcEwxjOccxZ4T6swhxpC5ac
jU4KPmPQesr6f4s+nIq5yJHeZRMCVhNSSL97FgwsEub6gM0mF77uxi8irZn9bUvt4eQhbmC2RXIZ
mcqhLrTaMFjV1ZNfiGA9kAOo28AaopeZQbO8ADQksPFIibG1TlX8qO6iei+joVPfWO9kSyAPnFqM
EVYQW1Fc3YqPsGTC65J091wOZCQG7psQLVkGVRnIZSKk0PsU5HU/iBrcqff+APJrTDoCQzYXc8/1
p/XPeQhquj0+pKW8GzOpZYkJRda8gxOMDQD1DTc2xIaaTomvLPeBo4YSkkyttHcp63jPoPy0todT
74meB5qTuL3vtZwyOPlYcyHMaE9R8x8S5V3zQQC89Fq+Y0efStuKDQ/UiiQvRhnprBPy6zDJ6Ue2
w7rNtjW/5nPkEkUKVWu1L9B2Yyfv/U9dtgNXizSLfWFTg47C3JmAwsoOWeHWMRIsZ3zpmxALcunK
ZapnZVxmbPu2+yTLtvPKLO1VYx0/EfPY9WV4U3o1kSJ/o+gB4wt20X8PLms4a1mqm+/CbIyxXOvA
WPcYkPhzJloR49t/eeKZZL8IzyynzSSmRNUTWdHol2sJMFJi7W0c4NV+mN1No4jTktyxarsliQmT
+m2QxSO87fP1+F+G5VAOHLazcwZOweplXDJympE28m5o1G4aH5tpff5VLDXV5jc/ikf3QpehOEDw
WtQkA2pyQmSm4JkBDOZVJKeHPNKKp2ftkEQznIIx6iDDSHfpjsrQb2Idue2EcO0qzibHbj1eOSHo
hw3idqV3/DsYnmAgspEif0sN/4k3RcquTDdULIcX6lKVyM++RrsLmA4EDbMn8T9VQq3uyC9PleSI
EODhQDZsN3bqhoZOwaXyRdFQUN5vXxbbM9/+Izox8V8tDhAgev3aHpYnGo62n3g0kjFXHKq8tmmR
ry1Sf94RXLbfsKPGA+D1xlEvP8Ry5duJOmm/zowT3N+11+DeX+a51peAGQWlJzazfH0l8CgccrPX
CKTBp0esvtVoouWD5AWRPhAM6AM+OeWJkxr4ehvvhUjcZCEB+G0oP6vyNefOWG+ntFnXd/+cwQxF
46ynEl969aOgulNobEuR65V3VFuJHDr+6YYfYyI/YPEGtS7V8CE8oXU9AgAO1PfWJlnzdmJAPzu0
lVlRT0rikSko19IT1bEjRCUAz73rUfr+OoEC79I3iEggTdEFvrZzqAIFG5tmV4oezyS8fl5i9NWA
nhRaFa6+NDCYX0LgoyoHzgxuGLCKLReQyfrVqF4NBbdhQgbU1MpyMN4pze7QyzmfmWhay4WHi81/
SChS/HwMrz1iWUNvruKWw7mn0Qr2tKJyd/dFjYankSMmMgjdpOfEvB6x63A0AOpxg5Z828jJ12eO
U+T9zwRII/dX+WPiQJBViZOXDe84v000vHq4k+OHbQSrVcGsjzHOsVHBTC2DNNhyeS88S1t068zm
RgKkQgINmzc3YTSjjL6bfiNm1qItDrzwy1Cz9xxtksGNSvFnp/xa9CnjnTfoPEOS5zaCmOAOe5i8
rUat+7rJHw6CvIsx5Xw1OSWjsFqBPMOCg3g/EtpUGOufdCJSRG0mlf7KGgdSVep5gpwtdHaiuuS2
YGNwxWmwm5zDpbI+2RvmvSFO3jSsSIxWBuZbCIPHwtwnAng5yGR1piwJPpek5lqVfeUKDztk3BFi
t3eEdZiVFd2qMgkvJ4kI3Oh+fxKnuIvJmb7jxRkaMdAEWcobnKw8CAqNu/b3HsAuXZ1KefUykCtO
YOtN87DW++c8hJmjCnJN5nNKFUBm8rtu5GfHMASpx5uTWmgBlRQUw5E90hXmG/NoO4xcwAB5sPnR
bAQmPMdGCl+7gn+VcquWy+EHGoTHxdiJ3LuYOYnnjqQPs8FRq0bJwZUHO3jU+UMjjgonD5Yf2tWP
yKNT6EFEB0E8HHUxoSbw75DWciYN/OVQzjvpXUIhcxJIi7r03RzCNQyP9qaHA+BR0laU9jbzJfcH
IHTbMTaBMhd41GhYCpZU8Vm+i4ldfQ42CqF/bUtRxEvPC8koyvrVtYjldn1X8Y7xNWN5eaf9fHRs
0P66TVa6vXf54K5a8CueVHjj2TXpwkrxszpuFU0PrDGqBwUv3cvZN33RkeXrU9kl60nX52rG7c4P
xLyclCsDCE2sgl3puTM+pYyfSYC1nQxCGsWoVn92B7f0d3l/rozbIGjMWt65bcTbxD+Xy+HrBure
S6ITstJGBIshxgYXT8JwI7dIkuKyP9O9HNQNKacC13raCws1XeB21WXfZ90r4r8a/XzJEukFpuPo
VLGPVu0JI4whHPmvQXslhNuto8t4yRCo2yBQiH3EW7EZ/sgXWQO+aJ5AFWfmJmPs/V0Pb1tGYJH/
1ZazoVoQlfI55ewgnWArPwwPQrpet+sfl4qt2hyId6Bgo9bBBkPCjvTNOaySuR1GQUTXxtsXu4G6
DHX3cCyziiutCfny3jiEZh2cVp0FtfbELpU3VtoEctgezryspi1Sbe2gCXYSBeCJDqAWLnyCcePJ
+98X5wNQeWAMqYoQUPlnILdppCim14LnfDy8FvUFxLdvaJyKXqKg4OKpq6yjRVQLPGioSSH2Uy1N
EdHH024+uPGWil6U/xXjH8btcoeHahB27i76+JQAkiZKEUCgbpvUm+H+vvvgV/T0eefUgnpwQ/U4
6SNtLCzO2c2yCZj1S+zbrwQxBV2O2P88FiNayUwy0Xf3d/SlZw6+PWr2RbwQ0ZtyHBXDGz01ffhV
ttreXVTJvC4PxTJ+z7cn6hzgXTgiNQadLFnfXP3bOQjY10H9h4QqHYnglFXH16KJTDV0TdB1Go2/
DJCU9G0OMN3NayRtII2Fp9z9KvbUrh/Cm+Ym9pUjBHJPIwqPVOg7fP+So2XPRY7bHKTiQM/8iIWe
26V+fPDx3WpoOH8zYxfpM1jz9MSNXJPj+ww1eie3bi8zhg1gjVAFF3IYYZ41BZFrdLeNg8oa72Fw
lWd8jos/iOxRUlrdxl+37nqRN1qw2qHRoqadEUvgHn+YqsqyAe8VmwMx8ty38TLrs17BP/1X/VDz
16acR4ai3ZKlYQJf0Msm2LusX7O4r6aZG3e2pdBWiEWq99OQN39skYzpUG6HEV+/XY3KUoSU9M7s
Me6dkp+PHnJrdFSLoarjTc/TmYgjrDUL+Cl28einX3Z3q8rtPFj2FRvZPXgQl8mSrllOP3xuq4mY
Npdy0xyjboBixbLykMTaNolniJZZMcs8VTDO8w/YHsdxlfrsJXAT7hoP5vIMaq8zWfy3r962zYMg
72kku2fVop8dRuDQg4Yt/Lm5gCEzStZyXLWYN1Kjn4PB5fwhJUwcMMsjY1Iwr8B8jbTyk/DYOaXO
yMNCUnwKTPofBmlC+eDOJuPwIuZnoQTpJZpHGeln9hnaE1rom2QcOZcve/yq9J4PGXYBmfD6IEOn
ZTLGxeWb5VDO+Ox6unaj7ttZlWr67/+oRFHD2XB3IEEZHLOfI7vw1k2bCSoe+W5R93E5rqR/hJTA
HuhAVVyIplIkvFIfKZ8j/Wptxf8Mzf1hssuom/zlVcEfb+c09JCXD1dKPxJwk2sOYX64p5iqf/Fp
es/7vbW8F5pbfzDVMIwmzBLZdDV3lU7/4gv0yf3UGduL0o5FEOlUBl6llrVzeAzjk78QDeKbHS4d
neBEls3vLJIp0FVfzqiRVMdfyYc6o1hL//UO5bLjkwYmdcOrYbFzc7kpmqeOXTDjUPtjBX9AId6t
+wWJQzF6IU97ULMspw2FLdiwEZD1nCvJLVHTty4AW/dFKcO14+OBNL5NOmY73MNZBsNEPQrA4lPV
3bTh0wjVvGIyjJq/ZpP+6pyxQ9cbAJzrXguQRe9PPHpN7CguPzCIBL3RAUvea32yblcWiPnGbjwk
NUxZV08Mm14sH6Vfu/juWHZjj2f31jQQHuJssEtMdg9SsuzCa+HYvxPYggCjc6V1DL/r7WmrgoZX
WvcD+W/HYbJv+GZXO0dmeYQvoYCSyANDRdXikTsKdXPhCM1C2HRjAasAO03EU4dZZuEw9pqkd2ND
sIsJB6RDAHoQFbJyYdAhYJ4CqQ3Naa0ox27NeDTS9fBaBZIhbVE4eGVyzwkx0xpjo7HrekJazbXG
kEh9gMc2ffc+nHSKIh2G/XOGC7cYgiyf1ZSDdAgbku1zUIozq3HTR6CkLdQfgICabYE0N2e4uPTW
67FjO+RLaCkWhNrhmJ0Gv18xchd7HVmrQX1ONIhCYaNeJqUwBDBO2w52DHRfrZoTXVKzme7tEj7A
aeMtQ1wVpOolZTjkZywNja9wUBZ4datV8nTUak9Nluo0CZydmBInt2SJMi8zL3mDOxruTh3qoIYo
/lAjhnZ2SMALYQVD/AcHYcfsB+5C/+oiJOB1fUutRUGZvs5GGdgDu7u+23Vi2P2faeGWtWxg22Po
UDvJYIIWJKgQRPaggzf/EEYpx6Y760Gz6pRA4MaTz04UcDC50+bazF4RA0+jnRLReDWBAlrtgnz2
2oYxJKC+9jUERhh6LBW/E7MnNzl20WP7XqTN6E35ZN+Dl4uTRhjfseEpmhQ2hB77kQhNNni83Wz0
o6bFcOALwSxxc6DQPsgDiFUBkgzjFht3Ejd+EdzXurzQK2NhsGElMCiEwJm7HtERr2Q9C0Z9ZWP0
iyDNeO9CtMUrwH68Up3XpWAv7OdVhg79LYhnc1qYgVkHHRBNJ3axoQAEdcCiLmUbD0TPlc6o2uWz
1txCh+Xy+/cXtFT/oqJJsx+BxdwqANBGjEI1Xf4P7ngzLdcvK71Pi2gXvF6VHBQ9waxoZfyPPKS1
7soqnZ3P50aTOoM9X8kxdzKbUzo0DCR/NQ7Uf4EA7TSTFbVSMc15M4EjqwWepjx91FdaPd/YoCME
yiqbucMpgAFE9OVUH0oP9Wop43rGbtoQexBb4iaSVJC9vt0zqilTSFOoZ885QNhNsNCXPhvc5ok3
zNSziF4pZ3kJpS9+0t1XSVV1s+IgIsx0QrMqANhv7u1LLGcZcFRFxM0MziK9IbWAvCj5uLEd5LaW
rPSBg5k/vN5EEk0eu6HgT7m5GU1wjLO1uRsyHl3g4pAGVgwkH0cnUWNrNCKq6j21kXLd/vt/w6nD
oV/SqShdb6uEpg2WLrA1dxZvAEmMP5iAOGmRZTm1SLOxlE6ec148rl9Mok0iiUCBizbwm7gYYTSH
o08eidR1J/sZuUEEiq6w3dL5ENYv/6WRkNAeA1ze7jY0kC6UCCGKm2WG+Ut0LsLIWB1IIqdp3AU2
40uQL6kZ3IN8GWv7PL+aE4T8DI+z5c4y4Hs2ZsGviav1FWBQUQQjnWfozqTpjfJTGD1HmqfuU1lH
qTF9lYBWsArOsBjHX/KaYs490G31WMQLYweVmjo9v0p5fnVA7+BzEtDlBQv3zFPkj5ZaPZzNT6i2
O3yjXgXudI8XgCu4G38n2wCMSTIIM9x7kcaw2RchE1UBE6hr0VucGX2acUoQo+gsxepaiRAPuUFc
3+Jan8M8Xg18agrIJN3c8MW7303yohbZ7KAozB9CVDEPM+W1dkNu04JubltAvLEmNeb7IrJsWJx5
cKw8Np38FZqVpwgicc7xIUNQk0z6M3p/mCb/C16QYL0ZdT4Xcw02xFIwFqxQ6qVseUCo6F6ehLyy
ooU19coZy31LI03re0FnbnpN5Ka+F+9gGhNU7VSH55NHIjfDntroLwJbmK0UCKp4y1Mcop2c/Aeo
5J3uKmX5/3o9d9qc4AXc0Wgooq242lySMi7bOa31aIie7knczfl5yVY8b2K2zzR6+x/5prH46D7+
+w05cysVdBSf2PT4nHV0vbxAVbkD3dZHEcJ/xER++gJvYeK21XOgA1l4MRNHu1T0VCCsPuk2Xv0l
+c3dyDXNyUeZHW5Qmtl9aVr1eui1X/KIk65VLza69G3E3nVrxll1JCCUSaVCv3BABrdfvNN9vuEI
Qrk+LIJI3vRB/QDAXoi1LZfSDL66MpLSuOfB+smypApu3C1DOeHFcVPTybqworx7Ve+hLq4M0SRT
NWLEhybR+pezcJspqjR5ji/KxuWv/AoAqsgdW9hT4s1n2OXJYdlj7vElrOUHKE181ZEfX3YngaTY
ULnNywjildrvHFFsIXz4SYQ7muaoZWVTMuG1aXkw5b426rLVlVoTUa6YNlCxVfXTmorD9v6+w+h7
pVYtxe0m+4f/KfIbAnyfGQ0mVLic9cTxqQlpGZEVb+Iq+g+tcoVvVCsR6hNsvaSzycRupKuc4Oq0
MvsE08URzgFYEJPKpToagpOYbEIOBOJdBRDysbiNlUeSTRmZlyc+FvSSFBW3dNztpASPleIH/4Bq
glTQd9u7VN5x0b9BvkmfiZlT2b6TRMabAVfF243m7K69Q1qANybqVtaaVfSGO6mBddDLfyPll9MY
zHcv1X8poYv/sHNDNcSLewiZu6kSfeLXodzZECTSLTuE6dGs
`protect end_protected

