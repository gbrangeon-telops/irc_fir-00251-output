

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
q/LTCQu22IewzFL2xoALv0V8R0cS+n3ZGOXTlz6zO0tHpf0bhYU3nG7YhbNw5H8bMFnHmKPTo6eG
UeGsZXmzfA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RYLOlBm3BPRhwpOnNgJH4Vt0qZdXkt6+qKeUVOFaD4rlCQUegbI8dSeedwyfmRhRBYYfcasAbBQY
SHt4NDprJvJn/h7vAd6X1UjRiIi8OF1s+lR2yqR+Y5n/Ai+CRx+BajVy1wGHxdjiCnM87Cq2Hq6s
UytlPbN46pRkluJe6NI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5Onxh89dWZfdY8AMW/MOzaZUaP+doVdup9B0riUkkwljU4WHOna1/K734H9kkMqSDTQ9ivkZIsmH
DErXjPeoJcAWqHloB9UX56vG6J+JtHhxXpnFa4rDUsDzFadXGZZrXqt/NJt/7/nP2AP1p1qeKRkq
ksYRHunueBYG/B5LuPR00cTpoZaaCYuJroh/pzkerIy/CPNX1RAKt047HCKtvFBXH7wuqo/yaUyk
Xkrxw2AQ0ggYgz1hK0KOdWT2JckcbGgVwPsik+mchcvmPUBKx8qFAnef+ZSGsUTy+3gjDznrQOsF
sJM7rKdsAjU5OLq3k8BWR36ur9hbMdk+lvFEHA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fe81XuZ9RrG7wwwI46b8GZQ5C9RFsRlLr0EzhGvkV3ZMeUUoQPwYfJl6GHoj+GDA9GnY0KeJe84A
xt/fhvb4h1DNhpVnvsOo41gu13r2msE3kvHyK8en6IodL/Mdh8CmalY/a7ZhDb0W+KP7rEAgisED
MHKHkmm4OWbTY9lIJCQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JHuY2RJ1GBIZ6g9aWOE7BqrGN8uQypqLnY0uHGFvCX6msmuceGWWswz4xbJBwz2/gb4ZfVDTzfAB
RXiuZlDm1B8txxWQYaxO0lZYlxtzCU/lUn47fRBxEhyn9Yc5lQx2oW3B/G9c81S8zCONQlmapnrX
y4OR/jDZXLz2wxMs0tkWUSXHisAbuRctLOTsTUfqMDUsJS1g+TDQCDpUDXL43sWg1LCRd7wDn0um
3q29OwHxtysopGOz0DxmTcK07ZEEnSJS89piniLxLQC53j2zOhAk7sCb4iRKccCVkkeasTjlcMTi
rJCab5WZRXi1gu1yWZ5s8tCfrKbGVSZTS8p+pg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57216)
`protect data_block
xO2OCx5Zlw5We/IjaMcgSMhuOVrX+4f+IwXtDHGgczCiB6IGsNty8R5IwsgnR46pDW//th82ABaa
bwmUHpwea+953uW9ADzA3ePqOBHpLiKPyPCjBUKa6K37/JGCSoF+iriexo1/D0EY9ZH9udYN6lZf
KVDr05MLJ50cW8cVslSTRSgbMTA+IATQhcbF/XMT6IYkxp8qd5abjrbmct2z7hc3a58ZpRNqtVKd
zj8MkOjfO5u+qDe+W7VpmnBm4Vv5lvyuNoOdFxhbi1MwIJeKqzX/ktbeKoV28g/zfNcCBgUjd7Be
q9zcExYIO9++qCLxDBJ6oMpqg9JJ57P8AMDPOOpZprYKV9y6AV5lRMyqeXRBrpmcqPaPQ7VmVqBT
Wmuq1i0EuJaKWX4Q02HG2x2zzvUcBz3GeLTk9QPqvY/dFl6tbW+fbfPmQg/jphgGOTjgtrLeW2J0
IMveOAOWKMI2wTdDhXpd2REXyfYOUu6wM1YKFml+PSsm3nHPLKF7wr3eCkkueHeHg62gISnoLD1r
4jfMySivayAJii24ZNbWalMl4NL8KutYMjpmeFQGIAss6B0iisarOpiN0Dyxd7WrT2KAI+d792bW
cjlx05wymhNfeoTstkV5zU153UFzWDlBe+xESkvBQJt4x2FhBdXcp9ciUKRLuv1OxgR+9luNEAiZ
6RBqV+eC7lv90y4SEvej9BgVijA3CYsP+oN5C+GJMbFY2cJ/2o9Ct2nHET/0zgHqS6jzsIKN1Rbt
AoJecLCqoAFm6d0mp6fHJ/440D/FiO1U074Qd1HG/sH6XwtLmCU+92/G9F2zYQcWA5KNkkfq3J2L
5CEAym0dl44CbYrEO5bNItRr3dDteNXIKSLe6nQ1HSGCwXVxI/QWxRF6iDROVjxt24ZgCC47g874
g7SKlBOj0i/8JxQAmWvwe16SooM1e3Z6s7j6/rygaWXpfm/tkVIltgOMPFgBQFwp7ZDlpboud8yi
hBD2OB93o15Lrbhy1SP5+MDAVzBUYVAw4HSWhpRW7Rm/3TE9Pt8jTjsLny1gd9RdD7lnbdx9l9dt
wLCUhmM2EUGvWY7FLghvgabL+pUJ0XVfltL8aFBPiTeWIJPcXpL/pPZdWzHfpV6ssBIhWVLZyRSm
xyL1cMi9cYhehh9ednK2DC8tddmx8Ky4d2VdpeW+Hcc2EU4FRvgbx8cTWEWFUX82+ZH8go+Abtfb
LELDheJ4z8adXIcgmdwkY1226CQvRuv+cGwGL17tLrRBz0s8TUbGyac69xJXkYRS3cetnURd9igF
jsfBeNWepet19Wn1U1Z72z+wI2QfrRsFQ/moae6hFdFqCCvxPm0H+6dT3p9Dyo6HzebP7hy6OXqI
6J/lhIau77KsrT1DXId8DnyPoOJj9PCXLE1KFtFohxWwD53IYP5A+nd3va6GmlLchVaRhvdIzIiN
Utiius+PmO+rOP0G443Hpzia2dmPw6UVnjs6cWoDA1xpLbPrjvYYq8s8noBmq3WbpRddbbceuP14
3XyJGVC/dMoVBS0j8pD4+VrF3yv1b6gdaDv7r+WCJgKlD5RLDRU44KlfeU9hysrmhIgwHPqh2Jdh
JeIr7vqklqSm+3ex0WJ/fhJjDvH5VwOxFD7YRp0EqyCat7UMVrgKpwHE0+pak18XscwSSTwAKNzd
7tuqV2l4rqjTkixLX0Togm0cveGO1ErtnVwZBcJT1mPHyX2/pDmY7UD9/O8pr+WJuBWN/EtHGi3e
4nOOt54/t6JnCGoPLKtT+xd+LhKcq/OMQJI1FrXm70F6kffAdkJEQm7R0AXV90oG/XtYh13i0xtT
CDwn+lzTTdW4HXtvZuxhOQhfwt2X9Sm4jw28JPyrOnme3hIPBpoh1QtR3w+ZxqO/AXHV9GRQrX3h
BpwjwUy+ZIRVUfiJdOZs7VivlGwQvXhvnqhe0mnMm1DjnFFrLmbLYtnBSA22xkxNhRUV/mf+qmy9
wEbt11mFBpT5oPDgbsNzq/wwUXRrmkI8SNqE1F9ZvEzMr8Wz+7QiFnDIzn/Q+f5b0DGy+LxcTVTH
/7I7dneeMdyskqMss16mL17W/vCfNM0ytFRIDqjP28SYzFXo4nbd6CGYb9bB8zuNfSPU9lyZa8UY
8Hx4OTMzeA0w1jr3BfXnPggoHHj50TPIN44SP/vjcbL33aU4BDN6/5q57I3Ri1oTsU+JlGpch5gX
RNXGFts3khfxZv/IBfKmsxWe36BOn+vR5a2i+RbwaoDYgJna1U8e3OBPO3xTPbImcJD5bLz0nLgQ
UFck0vWELhtUQ+zI31OkZ/aS83NHaBgsy7AnjkSG0NzxvMkKnTBf7/yzUaDIzYTwTgoECknwsibK
k8lVqhuMHpVGcNPb3/ef79PQXqDTJ0S2LImmemFr7up+IW3gFWvaGPd71xVL7nTsOLt52oROMmsE
N3NGPGYK2wnRUhiA7zWsgXNTJ6KYsqh06HWRJFfcsU0p/oMDmZpXXVK2HfP2yhHejXwxl3GcJkh8
iFe148yv9Dj3dKW8cnpBy0gEHQ+7PXfOhlBKl76UcneKPOSli93aetMSXLutYnZyYlNOpgl/CFT5
91kaofU+aaeB5rNCn3n5bAVXt8o7eQVznXetV8ng3QVDlaSEi7Cf3x8S/PYJw3NKxs3X3kc/B7kv
EL1CaWR1I3asHsYYGE9JXrntvBwfRGqrfvRC3NjCcMi4d/whq68wx6WMZL4XT/mGodsIJ3tz/2td
1hob74UAiCPngIfOhEJxNMjoVU4dwYhnWXvNvLzcQ2RicmiAtvCiZY03CummMqnnPx/k9KmXU2H6
oXK5OZtgL8X5I7Wn0KtlZPcpKrey8xuCh7vbH4e+JrRzodGQJkgzGPG7/eBiC9zT9HfYx0ZdKnnm
bnbMQEmw93KLcHiuoiAqKLhpwCJkJH+rULZUiQf27IjYCnOgFbJCBTlLSfUMtZVDhmyTSgHhkAHy
BOq5reiEGMXEZw6ql2uMTQY+2Tiu4fUebMjBKpPJ+TzW3Z7KsdMp1w3VdEoslpB1MIBsy1GHGTd5
qlMDmBQFxYgqwdrl8AjAFJvZtZgO27Texg2/9ILHVWwsJJld4NbHoaqtS7XYEGrpqzjbPW1SQjAF
2wEAOxkqbQyHB/hwYycDAqHttZVUqY6XDn4xqlYjorN8S/uMGz4alDvp7oygeVIUJwgvtb4WRvbn
2x85XYH0HeuE1S+9DYUMZqY8VGIGexDHrikwAHJjpdjcBr9Uije835Mhq/VwoKwYHxXiy3vaPBFX
2cVsWwa6jQ8sc9atq+hVcnhH0x1CZ3nAgpZWvQE5Vg2Op5fpJSfZfLoAjeEK6xbui5uE+g8LLti6
LdnZm/dZ9Lvuwl7qTuO3FP1YMV6I2HM6i0MqaChcTK8gfUIUXB8YDZBR83bImAJFyCigxGEV9n+e
KP3l/MkdilxrcBBGGJ6prj3b9Vx+C36pFhsmf67j5leaR+JN3stnwQvBwOYyEfIu4lPhN2TAKR3L
9gaE0qXAk8vkuINBCm4j2d7cVQzx5280tlFRa4NQza5foNdm2seePbLs5pZ1kiXTWwcfE2ssaKAC
eGLh8deBtOfi1N12N1G5MP2rTW9V3A/nsVFsLEGQItJWBK/dFh/PGL070j2YKphdbnR4vE6IDP/8
RwKe4ob6lfFz/RiDvq8HoKc1Ot6pAIxJ9D9Do3m2YRrypUcBL4nLFgS4kf7EwZi3oJvLGZP6JqTO
ZIMzrNwNMKNuZmedOWukIeCUydHt8pmttsJrmWYB5h2l0RGTNGSJ6mNiFWsyvkKIOzanGfFBt4kY
QzDvXZ0Akrzuaxny0mybxqOE31K6iAUhVnSG4u/EbOWv37rSsIZHOPr2lekzIk5Sn7rXWyvM7/1d
R+2VEHPxhtP0fUd6FamlM72S9zM3wguysJMOTURmom4oliI4lNNjNbFTKXSBKjKPYIaSUD1nelhK
//x56ZBk0DlAnouFrkso8fk7WXXa0O22+QjMC059/vIpvYR8CtFN6i6eoHOeVo9gc9XXuNhEA0fJ
fhoXlm3wJr0UE9X5W8PeQu9w+o506GVJFUmciussnr46crpgD3EFlYc7Hq67XtD93p3yhkF1oZ0+
93ouvN7lU8nO+H33LBxEc2bNzDQNDqRzOxWIg8e/E9BFMMGX+zad/s1zy1f6AnwluZ95bfuixSd0
iLYqy3SUGyc9fsnHbBY284LVrq9H/wmzFvHVf+RGxFTboYejPf9RoGINXMgXg/Fk2ncxZ+RJ37RC
80fE201fxaLrL3iuYd2N67gTWE4fQtiJTYBAtJi3NiGmzsaT4bqjTMWDaUGx2BW/dyCO/xtI+rVp
LMPhsuZn9AgT4E3JqpUp5W1jPUCp6Lx/YK/roIgztL4pQttNCFSHpasSMaNhMqHh+ancMjelQPY7
RFjvUwKs+MozvBpkzNzHM1NJxLW5hajt1QXmLSK8H56R25pGbZcUwtGqsRRx8aEVTjYZzesHUG7j
1o008FuVLovlyiYCdAAkeOaL1L4Ht2YGu7ctaCSwrLCcQOSc1RCLwUup+Fv5SrUhuY+cO8bEflfV
P/JvsD1v60zsV3CN9QY7Qhvqqb79jPZZFicXR2FM3CYMtddZ26U0lB4kkepMlLqxDcDbFhPEWqmJ
pDpsBqi86zYiGdJprP5pmwE8wd1yDGZHD18CZW4V01+X2veeH6XVz+hwfRTH5CIZP9OTMkB85zJ6
tDjg3fPA2sZtOzGeWL4UGd2GyVjAKLkqyZ0O7UpWzQ62Lu4J0JdNSfpgaP4g8BouaqzwDYzSLXfq
U6bKYaHvfXxO+6KoQWzCwHrfEZPns4Ov5pj3YMWbdQG69nOj3jLzIAYNKXQZCSQPv+mdrfnUCTpA
dG1NzC7kY0YdlH8LLlyPZK8wgNu448brOZlYz3DRrLexR7poKjheepv4x4gGeapn3m+kWLAKwdse
K9PGu1L6QJ1ifyxhY7fcJIfSu0UWJZiJumVV0hL4LeavFijYutvXbOKSguvrBI1mjA02kiSleCjm
0S2WYkbuov4MSC8jWxzDnfK3we4kCGnmb+uOfGv6ewJ+o1L3TnWh0yM9BaU76Gvme7wfK566nveg
V6Nt7V36FY1EczIsScc1eHCT1Sn0XtOOSNtAa+8ZMh69krE2BY+I8+1rEpaAQcj89kl1ephU3S2n
2dURsuWVXMHaN5kTQxOGBzYv6+D5AQKaAppzPdjA7+DFOWjxuhf+rp9H5nCR/Jw4kI6r8H5E5z30
2msSxJuEkiK7Mgz+no6l/ijPrU4NR+eBXik2NSVvSEq4V7JsDYifTPTixRgiSkjK825OltuVxn9/
i8sHpLMRS5o78N0TRn0IiZKdAvwPYqZxCP5F2xTsfXF32X3BhLj/B5nfm6gB9+NeLzEXqiODMX36
vZ2Q+OwyC2z36OiH5cx6Hr868AJ5yUVXpJ3wZLIs7iK0MgfmfY+izm6n6NSOuHtM5fuA4F6TPP9H
Ge7KIqevBFLNehpwoym1E+XgKwustHB16R7sbEw03ZGk9VVzNWD53rqpp+ghbH4OfpFOKYERq7iT
uufl/ckzq1x3o8Jua3eX5TMC7AEXkhMBvf0x6eKRTnkHCVx3igrRM3I1LYPP/J3Fv0cRShfnGQgJ
LrXTzNNyWOHYWvQBqh8+M9oC+7KkSZeYhmKSZBp9KJdysdFJ7nG026Icp5yhS7SLlfqlLr0i8oo2
0Yk5aqn2kKKcBYKk4cMj9o3nrY+vCwJ6ScPGf1FtwI1Q7xiFY1DL+C16Bt8oI+VO3AZ8VrsXoPYy
PQ35gEadGN9a7xdoyqNLN61cuZqAHcVm3d4AQP1e/F/NjU/EiJ0PPBUNvPnxAdKFB7YaDlLmBaLA
5R2aWfqPrgWE1/UiGM6cdpfGaUPsQFEW7JCAjQGOdiMPmOjNdD/BUtEKJ9xD7Ej+Io9YfFuw6Ee8
iHz6JP/eyAkiP+F575EEBIkcRvDEuh4o8tQDtViGE9f9VEu/cAqghqQjt2PZGfk+22OEHM+zkQw4
HnwTyB2Il4MvijIJUoig/G9Go0brHBEjDxrF1oEOHy00AzPCzO6DyDZxo7+riqE8Ombeb6u9mx64
c1J8IIyX8AmvLbjhypJEPx4sEmYm9wnD1pm5Zzj8bFJCwM3Ib5/5tmrh7+vzzCq71zpXT2QncOyW
QOz9JaoouUXc1l8j8hxB3LG95bF3Bm120OKyBDPTPNyPbwcxnel3PlW69+Js0U18PwHVgXi4ADZn
vTwTCgTkA07slD1O4AysJ1EvYUmALuwsmqUQqFYALLZaS+fpDbXnSjpvT42j/v+HbQQygEWqwZBo
1NEV6VSRH7Lw77+8kusiEhs65XWwlDLkDCnk+nn1FZRe8+blVx2lTgYmxPgCW1OQKE7v1O9VqZu2
/BKMpHzPj1UVPBHKXoNyUwmB1y/gteZ68+fPRG8EH2TiHJ2YF+DcaeZnNjxBbOOg6vKBoUw2jM5p
n/FTSxkm46dMEEM5cmLAQ8PS5NJq4HdGD2pvGUegXwEn8CsDmTTJG7N3A06sXoNWlDfzLc1oKQ2J
jsbZdxwd1kSBjurUtmZMTtJZ8UzEEHCS11d+Rzjl9xk7Ql3rnZRgZLHtW81Ky9oN0IV6kH7o1s/q
EnVoSXCe+bcaLPwF5Y+xY4gAmdOH6BOjx2+OCsrmXG71o2d/Z29KeKju4zqJgOkOhj/ymSgE9DjI
DMHg0adW19kpNxLdF897IFsDWYwfz9KBe/GllhzLE32MEFHDGvWYha68wJrB8oaScxA+x6FqredH
koK4bIL329/G3M4MqvYrObDQkT00A5TGpgYLCX3Qt8n0wIHtG9739OtYwHtRD2NE6NBDQZTI38u4
SorBsug5JMvybg5ibHVsyVI8viSQYj4TSbZ8gGFs6p7VvtVlPzUbOlCCjVKU1cBJswfLUnG0gm/Z
LBw143aEsifmd8uSjQsOMMrbAJoa6vepTLJGjp7paRj4LmnHOGIFomBTqZztExNGmzWAifcXa12i
eFVFnHYYF3DGI90vhf5mdG+xoFsaUpbe+ELd0qwxmYuSy3xgRSk4G1c2a7yi+aQey8gnepSpvzbO
KlKFnjx9jHc65+kajr7L7YirV7xZmvdHdrMRHSwlZhl/TLt6TejQqVSjrDmLKev4GBaQEl3Poa6e
FBG2kS0mSN6ts+C2koLxeGxS+tNNqKKMi225coz4jDantlVGa9My0zaZDiV+ELwGaeK94sIfdbTI
Drl6yr4Js9QznsBqRsAKSG2qqu4Jh1js+jOaWWUJsFbKzd3OzsyN7SteFrpSMFOeut4qOIKow/e4
ZPPLboS0v3cCez5UaLxbJKljZeQ7AV+C0eA5QLvDIQTKgHfEUHWHfkaIEuTHIhAjEtayA7YM4B+1
l0102FQtcn625uuJJ+eXJT6XdlxbVcmFYYs3yQRsSeUkPGRz57oCFcULOzp3Y+mMVwBXO2Bgahvo
ifVqcFXE23DXtHKOTX8CXokDX/fUub6/+diCTedOEpNCHmhwLC10h8yrJAbPZYCSqzaMiKJLbJwH
wa9DabV/REs2Qh3ez9Of1Q2Djg5E9ZQSLdzDJnoT663eE9CQHV/P2ozOvB6OY73E/O8ZXcJFx9Tl
WnpluVsW4DPv/7DtMXT7e9EL6iWsLIsWWfH/KMAX++5RqnmmZ2VCo/CO+z8Wc+aJOb9dbCCPXTs3
gCJovmfmww29wHSmU1DK0ivWCEyOml2rwuhcUpTvvgrSxcN4o9peOpqzk6y8ZfS4E+EIDJensKOf
G0Wk6Tu3hO9tPGpUGx0QHWfN90wXok+dzIlc5pPN43WTtqAismL4aMPRGWuhLiz3UD3ZRk7VR+Cy
biU9jAY/ysmXJ2LR3BvzUkcm9ygpcjjJRzk2evq05cT8pslBiAEx5ITGsNkKpsWgMvyc33C0F1T9
FkPOyWo9kgilGbGkKtKTuD0w/hfnEBRNwSCGaxTL3eum7qy9YaWOyYzEFtAfle9d7q260IkF6/r8
jgtwT321XTFDjx3a9EaLvem+szBtPcbLSh1I0FX/1JsWvhBtztK0TcEi+U6org1s2huHPCOhX0ST
N21otxIUCX1B0GMP0JtWiSFpdykKS0MltZGh9FKETQP4zCV5CTcTxaAWwzUIF/bbZKQKF9mmkUKs
a9bBb4Q72gPaCQCR4e8VH5GvVH2PEa/DXmErRDRvASNAchJBuoyGbaiRer1k3iDaO6knDL8Doqxr
GBY5YOellvjOJ6DRWN2Ci3fwwW2rDXWdzRQWQGWac+B6fo6DBYd84xtwOTzqUe9TdOes40/oU1hD
Tbl3AwRbziOvA8JI0qQPVXkC05wkuteuUfYOkGlWCYB+/vtfoquCFMXSYXuG9vZAuUtdaEP6s+ch
bDhL/T9+uHI4O0IzFymaX3inJfUQCnSBI6CdK7XjaQtOdOW0Lf8Auarb4HpaRh4pet5BkPP6lULo
vRh8oJlJtNchcZ2oOEZpVm7gciiFReDsiQaVOh7LeMicYL5la5bdOpd3wqpndo9pdk9CYaCPvEhP
izCNzT/lNA071rNK7zYKKFHDUqGNd1XB7ExtJaNHqv2EijzHASW3N1PGwyvBOb2l9Qhi3efW6Wvm
y/uHGYphLYF/KozXoHPTB9D3l55NwRZ3tCSBwPAFrPrntRjMnsSajzUSazfN7j9TswurUlJjB+Sa
s3ibuSQ2EAlyGuVv9deDaOOhvXUnhADVlN2OpwFLYrLR7gXbK4wUkyME103IkeIbn8OiAAXE8m0W
fonarDIkrWel+hiLrfxToZVFq80v5WCfYzS7C6bOn4hqCLY1dqgjZF1yw1QqOhopJYMFv6lu7U4r
0lg5lYgs2g/6BdqFXTdwQjztlNqSMBCqEBqjHXiqFXxEI+JM885DNYm65vXZBp82swqkfObxGP/s
C3pInfHJD5WATAsFPn9frJmU9clLGB3gL/MkxqVEwN1uxCG0x5u6bZMdavB8GC1t0iaO3KBAlHMx
pWag7EkJmpHAWGrNGJNG1SaQsYFcQD8Xgo4Q2Ncb4mHd8xp5L1BsWP6TcirYXNdVE2lQ2lj3DqV6
XLBVMeqk4+47X918X3CzNMNepW1dtTu6oDaNzop4FeypobWuk1t8L1030iwAr/FeG5MmWILd25zN
D4g2ALfb+0Gpe4LZFv513khDzOFC09L9xMrDkOwpAo33EPV4hehVjr+M61zmy0BptXTey5QOq35r
GU7Ai9+cuLz5ILvMRxbMH9cQ1QRhZFrKKO2IK5dch6lbuiScJJTqT+23rB0fH/7xCem6gZbFFYL5
euapXXVYX9hOhlG7+L5Fx2gUOSTm5QScfC4mKZc7pwerzRJjeRgLkxpXvw5vj90MN6LlUwE4AsUb
sSuLxIKGRqtM8E8bh2AKydinRFEXWuVXQed3rx++tXDsgIir5kVK1LAi0d4BdlOYxcTagF/UhvJ9
TgD4ZzYUnC4b9ViPd9Qbay1KfNnhED+5TfUhTATLMgyBTLIvh+OoVB84y4nQGORQcFwqaBV5qqkh
rNWgspKLCGjWYaZcEugOuwaFCdSySteK9pZlpC9pzchOHZP4JJ6Ka7IoX4ZhfF4rS3rI1y3qQ1DA
/peYFxWWu+cMXqK/2dpUrJqCiN9curIg/y2VcdVjPEoHDzPilbUaWfrYztYRTiq2VbtANUnlSDb1
zxZbLThNPpKJYFYPI0XhLXJT0+FgXTsf7eKX4/6b/EubUatuC2fXs/WXuH/ROKNsffcao8hQ1yFs
rrdLsDJgHp5sZtzYufyogWFiv+jc9XfrQVSXu4AXHiwJ6su1n13bW2UPl5AYDEtXt+D3dOU4IsMb
nf03Hd95ICQ+sqyy51euCsFBJez+p/WHL6MjWnBl6h6RCb4BzB00Hi4Ft5b0jcOAEDv36TAby5+L
dcKzkH0j/HRtLmu5MoQOUOkEAYAS3woY52XU9paix0ozriW/XEL8uKcHp1NFmCx7QLZ3LvfdELI3
DGQhHfB+6oD1SRbwMeuzTrsFxYDwSvap010P2kEHe8aF+PfOh78tBOO3Mq/HbYTNmXgpBDeKMjBJ
HKW8qfXw3cu4zz44RKeqljH6zfZIKzFUziIOMgs9F/e6Ha5rCbljndVcdCXY7sU9i7RoTdu9iWr2
yY5PcB7gQO1nOkxfestcpz9U+e78Rirs5dBuvbfeHtrfw4FMHEzqGDw28BWfEuCf4bQLk5p6bYVg
iGRPX+knmKDS1ieUnBKoL79I27jAGzhHtjdNprhJVEBf5zPJf/9u7+JBxn1ZGBDXOpJMP45hrPy4
PJpMUqmYboBmK35bVTY5b8wVyS/LQlmaNrK/OfmfgltW+e9Nboan6wVBcfSW6smDjAGxino8cde7
eSgxGkow9L48NqUNEtF6MOSXYRsiAEu7qUaiXEgbAMSYxAYYImTdt0vs5otn9SWi5vl1Ksb9VhPD
7sEbu76cbvKHSQ0l3a7IeBlcIXUxbGxc+qZCX0tOk+tCuEX9d9kIW0FXA7/7Grf7YNsp8pTU/7a8
rPoB0l44eEiLID1PB0059Qo2hOaCA/wakBg5GAipjNL8VNFdkLgj2UmAEW5Daz6GOi7KtOCgzG55
TuRV05wsEqh7CkKD1T5EEsO7Vr973myEWjwud9CbhYxPh9Z5YxlyJ1DlG3ntlR3ypKADqjl3c8IQ
ATYgpjCFiZU+kye9q21ZRpPdL1e3Oq/DKSWrVKuCNdxQhjJ+ghXpzOuiK78koPRu2Ylvd7pIVTjX
W/upI6upTwGYJKo4SIoIV4nATbebWjBbTI3CkxQ3NJbNrj6Z8xupPlR0azeQq6AK25BpFgzXNWBe
oChvUXWb8kQKdE5NJtgOSlcOdEEji3lRlPp7fAmaKCEJExo573Y3MpgvBkkDeL+uXrteWR3ZXpVT
ibdm1r/IcweC6jWNK8GEixCOuxrrBxto2nHadnr0WeU1MQOfWXf0xywdP+YrYSJf0gLUETvcLx3T
MGdadjU8ZoWQ5/MPFU2Xmh/PDZXNVGyRIM9u6dCBVhCgUlt2rSk3Xa94OlIiVGgKKpbRMugNv6dK
MG1qx7ihweHf3Hr2T7KB74fdSDnk2T4Xj/DhEcSkjPK41ZjhglaKiDsapz4LJk4p2DESC9lOIag8
c/1q74Ww51GDfx0gWVbDtkqScAkJOsQLLp5vC8gXt6DbW8iVXPjcqbtx5lsn75f1eprAzDI6fnOg
1toK3neJuOK74cehU47GZYuDs98pmntwRan/IdPnbhSrVFfZ4l9E76rfGPwanjPf4aQ/i3/4sdyr
o+vxuTPpE+BhMbHR+K7hDDREfBNXqjb17Z8SBT7ubs9qdkbWLexDDRqlSdAYvY8r71P2YWlnLrkI
Z7/Yk/zeJ73lRkmTwC+eis3f1DkfsXxk0dzHfFbJkNor8F7vr/DlIUvVq0dzf6BeCboeZrfGq5zv
YiEqKEpxJaRN/+5zA1mrJ0Y3SmPo9u1tWNJAkcCmshVMZuXmWZzCmfP1xc4LWlW/qIJ/jJyCbs5G
yX3PH7aV9WpwmvXzeQs9FW0azDAI/iOTNNlgQkaQxSm5dS07/f+52FRPjHU1rVjGH3hB5WxD4MVG
MMWnEWPdBynd+qQHBa6vlG+ffj90ZLP68t6cfhOeYWaeWZjCtdy901bk6BM4RAIOgv9fpQOKFMsY
k4eb2xZ/4hejJRd5Isw33LE4Im1nzjuTwy14xnEcpbk2qmPyBhUmTZtEr5i7ZBGeHyLVnf0+A9+R
1X7DcjKgSlP9kR2PGs+Z0bJNdLlsR+PkrYNYFZ4inMHnVCaxmCZQWPPrz8kjrr5cPuy+rw5Wu7x1
wDOTiyTPpWoayRjyJgCsPl/D+BRlff5fxP3a2WqnvfkORtfHppMw2viOP+CkWGGVZqp3cwyj2t80
IsJKKJZ7PhMun83Vb61Ie72O9B/+sPZXoN7SIQ+BpQ5r9VO5zn3KHHd6vLnrGNDD4I6+77io5ozi
EUqSii14X8MPJwJefphaSM/vIVLxRkBnZnvqHb4v42cr8ob4pbWZtG+JJpT81eHDy2T1e3v9c/G5
wRv4w78VVO1UavIcVQ/IPvK7wWm3BgQDMTQSEkMJ3YkQOeR8v9jNO0AMbpca7dAuRCftcJSXrNuI
HJmuJbtx5o6zvbWTVk1yOMmog+J3yUA2VNY69wGs3IIlhQr1myrhUW6e0QnCoIIOpVrzPgOxOdQr
AXAzZNSbywIMwz9TCGVjyZWzpQpIfoDdkb2CxZ11TrmqQCqVg3UbW/XlpfhWP0sTPXp4Rb7SD57+
IF5cnGsXgi3pWl5KIFiUd6YXEpJKpQdvdolxd1Jh9qK05g7kICxAEIq3hPMvGdDIDgWWSwjVGZkG
eQZ9XzK/Sr3o0y/lWveYmtZAsc0sDnj9de1a74MAUvOos/VKMEmcjOxQlvKiokyo7YZVJnDnLMMx
IFB302qL/q/zFWkHE3IFbxdvyah8ten8wME9U6kBniU3ahqNUElG3e1pxnX9b8Snwk/Jicz2fnJn
JMpCSOjcUFGx70r7LT1Z6PSgAxLGMblEatolQrJVGH7WfDXkdOkAi302Kw17mf1PfIfg58RjzIA7
kFXUfvEW0/UEilv550mptl6qTa/R65Nb4BfaXhJ4bKG2vUQzmb9hB3nx+ruNeAIukSn7jXge456T
EHyXRDXTxY0vTQjfx5WyWYYTd3PrGMW7BIhcCSch1k2B4mPi8Xr/zvtYw9O4KDhYNqRmzzDDm7ib
ALR2OYSeMKSUwPDSmp9dFhdSEq39PENZFs6Z0fFfXWuemZDKg7S4p5RNQwbV3O2vPqAkdl9lwASr
goHCIhvsHvcaEmfZ0Jy2s7TcSlqtwe89sALs7D5ZqJWFwbRur3BeTCkSlgjC7F/p0HYdLP5k41F0
zrPGgrQbtnk1nDm9cXOC3lvZrmZAmjxLgHBNgH8Kz/k/LNVVPVTBy2Td04r2y1Cvh/kL3j+adK4t
h+iUYZRUyq3p5G3yP2+16o/hYmZRJmnsbb0s15aroaulQgeZxM20B2ZPBvC4Eh4MoFGz2N3n9jRP
R2P+bFMOxG3qBpgutlSiEz2Na+GO9Vruob159kWs3motMQKnis3cAS08ZJFo5lCw+Xns2IwCeXVN
DvPrZ6ropwVXaNt6PHKtil8hgaGrqCjiR1RJap756nyt/uZhSWk9rHe5ek59tln29zK0bx+mP1cG
ZyTlRT8jba0Ut0Fd8cdx3dObL26RDsm0V+TXgy1BN0yyxOzcWXGz7ximWM6OVrq3FLC3Q+6kddMU
aQQcJVTxRhqSe1C87BAsq1y19AxmnNnnuCv6p/VLBPa6Hg5syFBN1BIw2BUu/rVKHG3ZI43OSOGX
DBF5Bq7/QkddnC8Z/y5r4HxEnpIj4ijyAxg+MjzeEF2yI1iheQDDv+vaLZUJEEe9U3EIsCVbG5wi
sGVJASMdj8r/Lvnsy6t+pzJ/4Vpl1GFwWtIPETRBr5kjFeCJdaDaGa7ssttMKWnEQ5V8njD6oSvX
xbESYIifU8uY8PDZ2NtVSwSZW0OxlBx+vklBcfuvRtuIvUSK+YLvkkk/y3sqCmNEXxj2nRUURXGy
GKCZAl4rFxo33zRLikNWi7QC0u6xjbaStocZ80npJtZWq0J3VnJ7OozqrgdQPwU61d5mtwxlR8ZI
GhwwWZyU9XmEZksndnxczH/T+ymyFRn5m497Bft5bTgldqY+s0V7VzpQO9jKwziciNFGvnCo3JmL
p829g/olt0ZDxE6YyO4gGvgN4N5jjnPOrEVh5fIHGID+L7sJ3acq3yJ00Zmq2DtWdy+DlPo1vMlu
7SFMcBDj6e9wPQheNnaNK9Vgh/J5K2YEudPuTquVZixpVgfufhMjUcYdWFRZPGX8UCG3w/gQiTf1
Cq+kr7qQ8PAVbnxev5Ers4TqfUxNJGsxKgD4D6ZdwVj3IXCQOWT7vp0133brgSUb8yFMK/JUCoD+
M9IOeSeEm9kvM2wB+Zx0vgYbCPq4++WkMVMeTKRrAAyRoJQUh0vUuPJbXi+qOUm2fUPuakffks74
v7ORy+FSsrIVW+OpQDGM8WZcwQuWYxQFx4KcnbMQuIP92Z7cf5mO8pSQqbrM64cVR18AwXIi5Ina
myyC+UzMokmBr7dL0snfdn6dZ7JjgvVOgS+DPoFNNuh4NEuSJ58WBgU+Wgru7AgMGb6TmH3a19aR
2yKzpcXeS+JGCotREBMoBlrsVd1XgwMXtrN4OnyIjEvFeNfiaWVh1dMGBjLbYFMhMBd1znVLZH/D
5RMeQdu09Gkwf0IfzqtFVoPYvvDA3TZxHT5FcBH6fvoHV+QRVkYJw1BQ71yJKCLT09mMymOgl/eM
Vq/7hiY+fD0zWAS3c6UirBH4CmPFNxhAou2oA1TDF4TuvqpzGpZD6fvulhgPV22032b9QD2YoHTi
vN010549q0qbESvRV7bHyiEdyz/ZfiZd74PKbtjdhrGwZv+XTUEEHCkUAizLxIqXI+/a7XNO94K5
IVO8JcJrWQOdVXxuiJwYI7VOZ4ZThIUEiNVvQM5Y42HVIOX20Ax6/CUNDh6HSZhF06lyeOYogkvj
zDMUgvdAacrr7B7F3W1kt59XPr/jzo+g/8a3+pY3FseiKWWy4l8desarKkl7bTg6/+id9uhhztYg
vV8sho1tMiGcZAFDzl0SGckOvmkfTEshF3pUr1s9l6CypWqs/CSZ26ipjN1Wy4GIwcOqyoV3hm6G
2thOlEkSfQlsy3W/zhsFEyYOT+J8vpscxn23aURoKWcRyPJRqUaM9ZClKheKoj6VpGp1FvY5nHbK
CRVGbpNIVxmewe/nJ1lcQGCPV56o9Or86qRmQ/h0R4K0NjgTSHnTevAs3HUCCpWyA9Fiy+am6/gP
yPp/2NyT4dH+x6jI2zIg8lyVYFi5EvbktnM33NDqvvlqbfNnSBHwj0MhY+cQAYF65mXLj+nxPLKp
BldLQTNDOOsLkmnJg/JeiTWwrJVf1uc+BtgjdpNgdTI1uzntm09hDAXKzP8WhH0mtwurWxdAn9yb
8XAV1fPLoz7LBUNLxnC4vtRZqfSgeTQuZsd5MATluzWtTPk47Y8R4XY0w0tHNtJsmrGdAVy9aKYf
sgUz5MiLPSPu+HNUdOZcFZe6yQH0qcjoc9BkK1Ffl0MiLXKRBwMbSr1Rkv8HY6U3b68I8hOPoO+8
zVnX9dAKVF3VTissOCfwoceMJlzpF9QQDM6yUSlsuCs44xN5Wos0z5rixxRtgO9WDt1dPK1pKULd
69+QwxBY+fTt8crWdfgo+xh929/O9yP2mSHiaOk1MqPbidXF1B8sW7VV1YjRsIWV5UGVQ6LmDwtw
fGjpTR6ktbX2F8hX7E3cJ/GlEUPKcKneefNahPF70bwg1TaZDTghjSj385vsKgFCGnnNFgQoVJbv
+lUjmLry28rlNSaAr3e4QSp5Re2fTx5P2iX6ssOvIMqKv4kwApdXRtXwiAi7u+P+7apyPY3Cu9Pi
psUQENWq51hMSsbHEvjlQaU4P1CrvzSva86+wz+ReKh8h/Y/+wJjE1vPQ6cA9m82OS+QWJZFODG4
/VOat9f+SYVvPQWzOSIBg7cMUL9HeN9WQ41B2ld2+CPdEbg+rcVeuo1r9ZYlasZGCoomSDwsIB1o
GwkgN1jFvGvpCoIsAhsL7D8RtoVy52LVBA9UNyJ8cPJL1WcYrvRGOi9GlXuKRMT5emQ6/SfZyhXQ
4KdpW/amcTxvqzQ52P1tZZdxagQG783P6SDCVxFMGx/BR6ETxaabZEA8UkX/BqiALPDv8anPSDxn
jpXjMZWYNei0iF8ObTspCXxTXXG31DSubhMWRJyntRcJMcZ+riaoFk6Dtxpz36Hc8iLV6bFoXr1K
vabT9qHVeXTqgyMYCILVCiF8R0buvdNjQCWa8ku4nNKn6+fYqzIRSz81+DglvmKe8cFpFsboideV
mr+HhgfdLsSy0XQuhq+liKaHpBpSrwBJFVl6X6NzFE2HlN7C2Xu77m8x9pv3OQLefcWIBxzza14f
049kjOUZl6YRAlSx4u25/mxF8rn6F/PidaQ6leiUrGvIe4yKFzSeZjpk/PCtklQO7eVrcA5OkNSH
ZoP9bdAdcxFLeFy7rbVC7jrnfC3wNKF/i0C5GyE+268r1flpoisyYh+QBH3KfFU4B1vbyJPjixbA
ZcleWvHD86HNyh0jvA/8r5Admg9c8CUYygGLES0NIlf8Oy826BsVqG9FCnhtbPyyKK3FTyzdgj3N
BfrYmUKIx0m0Uh7j5bRLijpI1VKR7X6x9N/ZsmKUAYQ3ZWenY3X9/pm2ZeHig7HHZ6XHa5uzx61Y
8wt3+A8Ca5ugx9INvjnDWeoh/S/fSzm9E7BFxgnSjabo4gtzBHP5876YtXyOxc5t+NbHUxG+13Eh
zsCHAZIkG72RKfx5GV7otCsn84wq4fRQKzb1EfWfrIkQlUSfLzEwx/4gpHBph9Ou2mdftberhwx5
lTtN9Hcs0Xe6z4jPqmC5E0SxnxlkEn4HQ0GPHMJhOW63Y5nLxNV8DE5PE+hz1WcCod53L8JDkwjT
EMcenMcNao8esOgMUhbkW7z8rAKcunyBVfKMhLsu2BOmbNSaXnipQQM85hX0R0ji0KvCrujtW1GG
EvUXRg3coJciw7Y51u4FoQK7f/2VrRt4bGuGdeqfeIyGzZvuxAVQLUSd0mxCeM1S3ltIG1yEAiua
XQ/6+qX5xfunDZ/vTTdOBFSGR5wilNfvh/G8bzOXA95e6eoobhFdwSzWBOC4pDBKVEX/afSZE5AW
yf3YFd1/BWuIJJ+zr1hqawt1E6dLqqNaVLhv4g2FQhusgy6nsGggGcOku8B7FYqsTU9a+XMaGQ1l
MDvH3bredxR8oftvUn2ssGvWX+o6gn5CgcRPkLZIpFdEbTfl9+VQiv72oR/sI9dH1Pu7Sd+iJcVM
Oan/WJmeRyIoayBnAO4RKnY7RsDgBSSGvZ6GWuoK/l52BJYMouIN32Wx3FQbZ86vRUKUkFhNbjk0
2On6U7WL1uKsr5WWB3hNfA7GeNt0gy/XSFw9Sw8FLPOJntgC+I8qvWpfHDlTXKN5PrUuHbHW0Zl2
6vGzmqedgiGTkx3Two4FgWSgxXdcztJ3yP4aLU90apWHbmOPqgY2aP5IZ3l+CbnjM0g+ygjevfPM
ieWXSuwmvP1rKQajFtRCBr2ZYJptJiuFmJ4Vh72gntiB4IdUuA4RszCOfV8i2K2o70ihMhOZ2smC
Rk/P8sH819MUZsk12H5osu56Sug0P9JVDJzJKzt0Z8EuJF0Fu5mxU9No+K+Y65blkHjvYtRfMEy8
526rsAnaXhuH9AX9XjKS39KqveN+jW3GqQbs2esWOWKCOzq8wZuS/EAR2H/YMzsnXd58S8UKrY4M
8S3oreqZGKuPN2zjz+4GvaVThEoPAAafieeLvH8uvHKhNhhOLVCtokcCf81V7g2lhpSQdbKx+b/f
mP3uPcchxInhAzg5CKD2B0OhtsBf8/BKLSGtHZUD0RUtDExZ4WPi4/v1swYCDZdXamEKQLhmQolX
f4W+QQgdEnB9a0mDI50qCB+M7HnQpPchaWPc8SXneUN9iGedYbhYkoZStxG6js8/euTZMcnambaP
/mVAeiXvUmY5H6Cs1BQrDEQoOv0eTTwP7WY6kY7Qlq5PKctshBM1oONvdaAcftqiN2JL4bVYzjDe
VTAPkMuwU9ZO6biP+HK2VOjHlXxrmJAq3A5Z29X2Kff2eEbPPCqSwXwEpd+Y2JzL4lyd5PoNH2Xg
do0oHCWvuzsMuYi2fvyB9nsDHEeGbEE/cmrW7H1wDZ/PKOy26Q9sSOVjTGLuvcz7b/4UpOzTjgqj
A6fVSh1lDrDopb0k3k+fyfJD3fG2zxHij0XMMqHSvTLKjwIO3JK2NnRyKyBfE4G6iu7ExI6Feo9n
/z2KadmpjSKIiXRMuXlGn0KOoFXP4GfuYxOk2F6PSHbzya1zc72Zz9QPfbUNXx0tQ1HJVODPnGK1
IfGXlnk/4DWyJd5nOhyX3Ge6Y+35iCzJpm4Yz37iYpzj2pyauTvc5K/7qkcNCsLB6KuvaTkbC0CK
8le4o0/EQ1Zs0riAjwbBQvF3vN9y+vg5uXe96Z9bt6arvv2owsxUzlLcDEaCe+KGuHkquYcmpycO
tXufljcd5G30PZF83vwVh5wVO5F5pmyAHtLhhtSUlko++SJSCSd0JW9mqusAtmgP7fHJt9fT7Su7
ttTucAGHlddHMfbUSHPp5WrJz6lgVlGj9A2IwBekPTq05X5JXEmidUNRmQQrqxLTGby7mPF5NW07
d2u6+Dp766d3GgqEGyP3ArQ2jbRfRn0PTlARBXTvov0EWzRNfoefqHwWicTBGngP8yf9MzyiYFoO
JTM0SwLNqzuxlzGFLCnLFjFUNehmscxHbJwPjEZN8sWAGMf1RBM5z11YL4rvPaS254voMSQXOEtK
SvOK9Q1En+Spp6djdgMhi1pSX2kZWcwSGr6CsKILZozj+9LJ/D6tbmMCU4kgQ8UO9QI1Xc1BwNRA
X0m/phJmkGrI9hxz3rFVpHw3aIX9fiVn7S6EFCyT3w5WJkQUh8vt6w79XBnfyaNqEQCfYAyTfiAI
sGwwW6msQ7N4zQA03s5NkwWI0H97iSArA0/w2LF7ypdJB6PuQJFZgW1dNw/IjcjBqN8/SEccq+ha
0X9XLXPX+fCtXPlPzpjQOrF+uowygbFZ8wYM+GDmM6hD+GvqsT3xSMfj7gwJRkZZ+WcwNkTBrZse
5R9zuKabxNbLs7yfI8C4j+JDekwxbsOETd5WPcGk/VCazhAH3UxDpevoB4yvcs2wh5yExqkZ0Mvk
g1byi5vV+krv/AU9pEqzGtyGKLaBiW17dNn6b0h+YEmgvUbn5nK8P1NmkAbwI0R+0AX8sXTHXGxh
zAwMGSmoskPqf6sdjAygR4+u3R+LCC90e/MvcE7MlBh5wjs7FxdS+EGxtI6t8aTodwj//Jis3ePa
CGzT8FLRz4PShfeA5Gzt1gGr/JtMRDxGOdZymqp/vZKTRIZfrKO7U1RlSu2VZT4eq8JIVx8kHr2c
3IKSU1Z5ug+XfpkTTZS37eubUbtInJ9oShN+SdzjLH5t9D4uXZg4fIskPyIy2b3qosbEoAJTMHU/
epIgpA3g+gh3U7OL42Ov0rUl0HokDzBNqJK3E5uijLdz2hMDKYxjD6qN8B3/oSglgIdswzlO2IDH
IwebS02aHOye+qRh/amH/8zQF/uMgADszMNbfB/acDL8TFH4VrT/4fjb/PWJiKvtLc3NNbd4a1Xl
bAtWW2Yoqqo+PdAZgR1ztrjg8e7EOQ7VNcqEADytpRpOhd82E0s2QHTAI7g0dCMqd+zl1paFwoBv
TKZVWpF6Fd5lv+oA/1+cA7mgKn2XP8eQTshFJhh2M4tvbq4xZPzv7D7WNlwJWQGAUqmWpcWSi/XK
O0cvdFBQgG1rfOW8gOO1ibQbXrB1FLQBp8XIXTxzo+G4CcgqcKD0z2YHaICwck+kwGAR6KX0EOfu
B71RLvrm/IoVpJ4CrfatlK4ZeCDF7i48KQqPJSU1o9xCY2Opbw+BGkokBiNNCjNTYIBt6N+iwTcV
4S9hEzOeL1/oelTpypAxHSudl4dVrQeN/pgCfzTFNtT6VWPfyCcerJubWDQWvTosTzB3eCN6C7Jd
4VlHkQD9JBPylZ9SzYikJlQfb5rAQQlwLVx4vHNy2qpJQqsjLXt9t6xS+M9/aNnB4vrWt4mw+ShY
IhzzpkUXdfzJ1BF0XKpvjm7hHrGbHyaFlULzekFllk8/MtrishBmcxm09/raiCl0FYkYM/g5P/Tj
WJhHbTVCQuiGMHXDNwxr/OXyqePq7swzrXROltQwvMIBkXfBFaKOG6wzOuAar+jX3X0zIG8X2qnO
jSjB7+8X0TxvDhllyPfN0YEdyRqSxGM3x4HiQv6f3GwRY36LeER2+zk3aaT+KxyuN4PhlQoBAgz1
+qADV9fxoHzX0l0Sna8ohfOAjW9gS0NnDg+WMpqL1bbHWyuLaPOHitE7tjxlx0hOwkCUhBemd00L
OfDfIm+bxZoDGyTuEJd6gfQpTr3QT1FGLjjE/oSXzqYIUfFr+If2QWeCGdexiLpi+E6HebxrPlTV
152iSrl48B44kIa2/kgYTcq2VWDdbJfLYfFxUYVtKpAGW5J0dkPhdJKZWgbd1P5GHhyqakh1JHfz
1reXsgfg7c8pBsf+Ul8UmYRrVb5RQoxAOp834frbX8wPr+4SSZ04fj4E37+QFfGY1arfzGNaM+Yk
+3ynluCGvNOTntqEentTwsX2/a8itUwy91BGcQqQ6Go42vvQSYm+l5bSN3aSEPYFuzA5VXKvrGod
8Vs+hnXDM4opnQZ5RujvG36uy2ii5ALL6ArVLiab+ji1rK17rIEddinHvRM5LLUItE3c4pe4eipM
LSXPnuiJgfElG7AkuFLQwmGJdbWho8TFpDUQx1cVFMfghCrZkQLoE6nNHNy1dhwuX1bGsJJ+o89X
v+iOyzQezCZyAj8HzNnZylcPIzajRWWtVVpd8RJfuA3UwhauJF6g8eV9u4G41mSdJyM7timSaXtx
inJkCcMQp6g39Cz+iVYBwLt/oBfZial0zCdw1YWVXRL8eQrRUhE8hyFnYikAdoTvLW1Na/exRsOY
1LlnyM+92jai8RHlBIMUckzr5emM2bqfbni5lrTkkEzJLw7B27HKMk0U04UhiUYgjfgHqRRf61fR
hVxS3CWPmxvmcLSYO3XZfAD0ZyqbZehjc2nIGrF7ZJii8QCgqhCTLJktF0hvbFMf2BcXag+LxRKB
zAydweFp/3rJw6dZMN1sHMSnW6ISvTGXUntAyKSu6VyRIy4zDtlcCDHNOv7oKUWt3kQ7KQB8qgdV
tQkrvAiUfZI/yJj+IW0AYqouXkhA+sxIkCf5KZ3k/UAipLcrdxjsYS+uBrho1CBK+e6pKZ/5rWWq
LxUX9d9xgZZsYO70GOTdrmg3Mt78IV8bszC5I/iFL+i4J+peFZ39fMTqZ2f6e5qM6TfL6l9TgU5/
Og4fm3SrMnIRGAwfHotZmBjMVF5q+FYxmJ0TE0UNRaejbj68p9cV6sUzwtb9JS2E/oWoWpkYFo8K
rwL35gEl3CNIm38+ovuOyVaSxBGRR4h7ImZLpOL4zrXxJSTEQHRCsAaaIJhvi4VVqYH1ZlzX9/kq
gCKDDLKeEdhpoGagvg71J31KOMlWR4KCMFmBHXGa6yJDSvcF4jfRYUW+/56eEC5Wz7BEbM9ipCPD
4SZFE7hFObXt2isR0vxiNGXg3nVxzW26TFFGY0D4mpZG1MZvK1blg99dN+bOUGuDLsOWnrbJ8F/5
jXJ4HIL2mqEdyNBZ4T/IJIzhFqbRlinnjkgLayytldTAF9KRHhw0QtYSvAoCZLtYi7Eo9VTQovqN
bKWkA5ixXIfFd8rUK3+pmfEf69eHtTPUMttdPjMW+GPHehaDINM5eBxGZgNPl+kWg6TCmBlSBJpS
6gJK/dVnJaHrJ5erQ8BtcUU27jhaUp4S2e0BqwP7cfSg0XhJly9mDCd1722A5LzE+UzhKYGTJP+E
cGEsglXnAmGGqP288hICwE90hbId/dtEnLCJQ7xX+osTE05jYv/9689CSKbU3/VEwUvzlpmqBsGK
3357HP7T1pxEevuUqsq/wgrphnK0Rp9Ai5wgdOLX9QjS9udDMzANlCWKvZrmZuYIM25QUuPITTbt
5PTjlmi82/Tes9r+gjwla8XzA+Eg5Wy32NLATS7OtURHEVli8gqLRKgw2XnKyPBYnaLPMGu7Nty6
HD5svvfJRFvTIuGTHBM2ukgWs5V4oi9Qfp9kIEm7K89E430Vg4bobSX0pZn7CuSMN9EUXGF5FQXz
ZJ3gxI2E90jd+FPo5QrykqO+rNKpe4D6sLFqsx/D7utzeIg6sPTTpTm+BXU1R3aEdfuKegUA33o1
DtJTMe9gKZ8SSYJMvESnkG8MOlHDQQ812J+qujGJcpbR/R9l68Un+s5gxgpsiSrWg9DJWlXCKKte
RqAhHtLtBwy1UqgRGGh3EJ5RIbzL7K/4CiUpAVR76k5P0rl/YiPVmZ7inA+uGoHcTnQthc9aLkj0
v+VeA4cw9NwgWUHJi1DX+3rqmWyHIoe+aT8EAQAwU+zjrlUpVx6AIWOQwd9gRPLfmr13jhwhc9YG
o2d9r2XXu3AWqHmGr2qYuTHoRsDoHpomP9MmASI4byTUqwD+uIFHMdwBAnKWpHhWPzKqUMyOXW8V
/deKGL9w3J41nIkBDmqIcKotlVYReCn+y0T7OnDIJsf2JArnfygRx+odMk3+dLsWVZNUCYGR5Yxe
8CAA+bNdmwzkUGsjv0CrEPqMjVOCDNioEdYAEmdaAyRh6hQZbvEN5PYT5eZmctFrgMZpNXyNpVMD
pGgB/Wc3SDHlAKYStERBcBGLEN6h44ZyA8Lj6S34dsHip4F7/8jswUluxqQEIa0CFcWNcAG5UyBF
U4uyDIi0tapO6eKvoRKad/JNHsjx2QaW0xVfj+fWRipjwdTaxNIqMmObN2e118TdHzXMsb8mwQbg
231p9Q45TNwQZOO6pjZrw4xJ+zHZOVwMu0Da9100b8tHuFSVyoYN4l5wai5krhyrN/F2YdVX6ojn
63T8DNKM+hAC1jj7H/FyLtOEv64o+WYJ8sF0NZqmvftgOEe+88gj5QhqsGIErNFzAI1spfKcGYla
j/quI6kPXkkYSvtHKRDsFoBnpMCeveaAzfT4nd7rbQHXTTUzUJbxXL2/Soxw0DAcSy67M24TNXOB
FwAiYHDhok7ikVNv19TbQpSkMorMZsg1OoXasc1hEzu9hR0R9qCZmEL/nVn9gmvSvNlglazKiAhS
qwZ0CLJqh7E0GzzFV5eE2U9ZBROAeUyvtIm0jRQpdpUTVLzJW49tn6yj6XESIIGFHpJshMQ2QCdR
U5WvoBbtKYSmYN95m9NvXK7yrjsYfEL6/do3hhUlUcBd6Ut8izDZVyaRjqb2/IAPZ4wSRzf+3oFE
NvHsl+AIZ7zot6gcegPk4VePbuiuJ+3KF/MkhQ337cBMsaXSlzC63bzKV8wlgcxp9N9cmsi6Oto+
2fyjPr/1m+zLEWKp+zasJjQOX5/KCcJ2qwd8DfXWhRnXlxcfLTbAuGkqiu9keM2Z8ExjPRwqwV2M
PWvM/8cUENw2CrLg5PT7OxnYTXQ0EDW/EbHXvrvJo7PbhoTwgJg2sctjryuBlyUpkUyKycbkX1U4
eN9yt4KWHPcHWfi0KlfpPOfY9KBqZzf4Byp89ioR3WP7GSrqyO5fa9V9ByJ6+coYXJgqD5dJ4ZZy
3XtcaNVoHqyO75x+IMdYGlC9UCLP8tnT2clLIeHECIHNoxGli+gIJJ0qk3Hz7EQH2/gxQQdMCn2k
vtw9i89vxqFt0Jc1/miewcrkuUDGEvFOoEAyr3EFygmVxgjujQGnXcBvppmf/J0VhYNvtI5NfI0f
uWMtSqXeNtrJf5TyB7/aO4vF1VqjkPF/CVq+osJM2XYkFqQV/nOKLvRg6g3OgfBrLLGJWKWVnbQU
z421NLUgKdEUPdVdDItz9WkdB70jLaFzAEIDcSigVrOPJ5iUmAHAyJwLLjYAc+hWscUGdV4niVc7
h7pQVM02CtVd7lxbr0r5JMWO+LekREDqzKPIZU8cuj/QT1wxspJBwZfSfQdDAjdYZtnzcxay2C8m
SXpq6ubtYoNe/gphjL3OTBcCnAYzP+1hE4ttCeaprnQ8/J3FBxSS7e+6KXR9n9k+zHO81JQ/7XU9
WCDS2/BvK+pB72nd3pm8TSNwmcwDno26P5QXBBVAw+uAPyt9pwNS/3E6UiVBTdMsMjcpevNU9JG0
CXtgdoUXITrBZ1NKmPHciCT7bKs0LwpwNQl8NeZBMk63LL2HzPSwhKwNEPnwMtNjkFZf4bqRpB1o
XXKjcOiDpCofdyHBT4+IX7xB4bGW3sZbwfyOLQdYdM4fulwokHFHd5Db/AzvdFWS5sSwgK3sI1kA
ZvwBssjpKym5Pp9zjSGABABoyEdkqCvH5aRb+APRWrVZ7b5gw0Bf4aWo5/4OMYLry2WXAe4n9usC
ZulEvv6FjlzxdGhQ219SSCZoY++rawvhbrg3wq9UbHLOI4xC1zNcScOwiBn4mnQk5kG/7plSCbCt
znjOBc0RDIdK+BNckIVVBq+foXK19WJlTYU14is5ACZ4cPexFVNdZV5eqJxN7X+IPXxgOlyBn2kF
3NuWHuZqylwL+Y0r0+nTgF4tWxpO2kvH9l/o7uGAz2ujrtIOcF+BoCDYlE0Jkeb9vSxZgnibVdVU
HSGNbBJYnmelp15s7cNU4zk3ioz19+2nnUg1oX+BqxPxepeC3EgZoJyZ2KysmjrGH2Rl98ApcqIT
EwqMyoNyqeueJoqRyNbEC06qOebh35wYyOeuBnrBB5cK7qaz1IhAzg5GMmfmdZDyslRjnoINHdVL
NXmXY9kJoYQMtz8cvNEqsyH21dL3oXT07aDbnPvRRmUOK2kiXDvSAw/PStevFfJyvmMn8q97IVnL
hIuiAUpaLTzcbMe2E69AVh+doB9d3JaQfmOTCPOCx+/EMzLgSTEmRtGWZc+Cny0ARC47rjFxphXn
1HHmi7h7O+8caI/sOfEdEoi1U5JwjLc/PEuB9tM2Ul2LW85WfERJD+DisiygZuTsPVHAPe+oAN14
Q89Trwja56M9QnSDhJeH0jcJx1sypgVTEMXQ2NRKgaViVjDOhOnOO2rIimRx0OsFuQbyjGOmJ99W
SjS/LEdqKPkhOXxrRrE/fNtzY35ABhfHrdgr7O09pi96LF1fACTLx8NBZ7lR8TfNEM+XMpSAp6EW
xmrhrAz3xOHTltuMhHv44zEKujjZn27ohdPSY3ww/Tcs5HrcjsMPqkDLjm5QHfKywZgSh3do1GR7
nt+h0Pic03zEuFgNU9tK3nlEUqwCUS/cpZdSxisZz4l1V88D1Efko+lDanjUStDtQHne3g9mPFuY
Kv/xea7wDqGrfY5E/MfF2ZOwR+xG9dLEN5YS1wurYeVz3IpRGkp6BDnmG+Clk/i1iAd/GH+a31gx
h8aFq8kQBY4OimtYo45zjAJCWiqxdp+HDaLjTUW30dNyTF2ojvdnezUNbcbgg9cWoYhy21ZqBRgu
k7a8+Wqql5hUG9w67g+gB5MW3o4Tpc3IObkDwyzSGCoopwFhxzZmk0QtSsVy80p1Ofto19jpFi/6
p8Q4sHlxo5dHDNHT+mjq3Ns/eOhCwsttM98iVZuAS0O2EO/DQ7IjBYok8YIuReo6i8NaRQ8anwFW
rjjA7MEJ6VVSjtl+4KWyVrjRxWKdVhaUxyLWQCGqLAJKyU43ZAWC60ZhG9NqerufdusP9vSYK6GA
1UhhdbNDG8gfDvdVG7ffeXIiezzE3YEMhKzqS+PTC3JwCCd+RAdAWIxsYIUZnoqJhL0lz4XiO6JV
M5MQnMvZ0UfhOqKUXbrhlTl/pY7YuU3Hfc4SrLnilIWlzUJJUhZWHIHlKP9+tpHqhkJkti6bcMpu
6LynOwqA9IIRBnZv6nebcnHJnAg/Fu8T0TlHcsa3n6VlbxK5haaI41lLA+E+FckTH4SXzxyKPGbM
g3YdeM0atu9bVYoqwiA5M1Lr18Viw2r7vdO0/j4XDLhbEifPZ8iHpWR3gjQOscMjMLmBdyrNUR4N
qN4DwIOkAhK6Gd1FOy9N4ZDG+UnKsnFd8p0F8P7UaDGsRiFkG31YurSVupv1Np1iUBsNH9V0D1oC
a1eIPKsPQ17yPd7m7BC8kifRTzzyLXWU0c/EpUQ66nvsqbmtDicbUUg+3OfVIkmhwGoleLMFO+iq
+Jb/FXyx5GBIVKlis8SPcjOTh2HFo7qNQYV6EMZFsuFPfpN5xeHU6+Jpely5ekXBIyZgav9d2JyW
UmtNo9D4Su0XIdlGj5qApgwEA6SGEccv2XSsqPpMOs7me2Y8nKM49kuyJTRuh1waFGgXthAdJjQj
r0yf+csjfTkiZOnTUaNsYWswmBDeDu5VPXAoaCbuUcXl7BdRBsMWaQow66md+XnDaQon+Icq6BGP
AYOeOBny/OjoCL9pzXSo/6Dw6EMdeWv7ErmuAsFWxIbBtzv7oM6taC54vmymFKYFYZ10rtMIpCtt
IvSp6pSiOPm1PVCHIw/powI2KcLP3lzEv6a9KOVBk11lp5LQkpUp+snRnf5HDgwAq69NB9ls7mLJ
68veeq1tff6vW1NrjMdTJU6AUlDbJHO9FzGwctZUxlN3PbmRzj1hBbYnFL5/EGoW51u0Xwv6zCIK
+LI+d8IP8g2q3ylTK3ith3GWYsjKNV8apmtLMSkJkuuRmJ9YlPhP0OT7PCFyQWwE+ZDVLp+yirGa
NXGILmHKdJmTNGtDHGFQpy9+L7VG2J5EKu/kKFpc6MTjwNNqWfHCS4fL6G0QxAK9m9ovFrI4UHV1
Gj9w3DqcPKUN7Q5DkDcGdi3Wi2KL/YRgqVsX0VF5/DBl7ltO/WJmHoTPMIZScjbtOeT2Qi3cxyF7
ftRPag0km9GwhsZFX0G9DXTdlWCZtGVnNNeGcSXDCSgQeGg7SwbKYaUkwU7QFDd0LcyZ7kJi0BjV
K1SJ0phwd4a74Fphdzaqi7fyiPKb8tT2jwwaAmat8z7Bw+eUjd7inuBvy6PMjVpy0zymzn0DbC1+
kem04oibMSozlt2D2vAqhte0LPN5433BAwLZLvbpe/Uf+aZZxmQAlvpi3NoTl7L7qOcNsI/FEgTm
H43XXsLyC5iH5vTRbxGDso+EXAVzPZSTqvm3Uo/O3+Se+g21gxDZJl2J4cTpGMgH/kBpgEm4q8jt
T6HjLMRHmlZwfIXQMXSYZXtuPkzNY5Qazel/119lr76ueBKaE8ACmPCGFhtwQCAstpn4rh5zZRHZ
FUQZpFbKcGVwCk7tiKd0BFIKyDZMI+kSoV1dVonb0H5H4qah5pLuPujc19SyMuZvQvKLXK0Tf3jH
8MasKY3lOdJHKsB8wStiI97aBKjWNw4l4Rqw+qBaexuQXRAIgqpX5KTS0/Imhe6OzhJKHeZ8WMDr
9FymIrC1jAnjxjV+YoG6KXyiaZJA+Kp+greHoSalogU93/D9nKFbl1US0XzLuUVNmL1qnYuJvig0
HIjkfQLMRGP9aKYLWGyfufvm2UBaKXJkMS0pjHQJAmwagDFoWup5QFviLL8pB1sM+yZRginKrYhM
to+C11MUlPP/ic79IFbF6srI9onoBFT2yUB7L8nxWPoljYgH4vV9gyLvdNDf8k7l66bOgrhCYH7J
kv2AES8N2JOJ+7VfpXWP+0UjG73zy4239f96dFwHo/vPgbJjgDZKggV0HAFbeTqhe2tCrJPCDdo9
BRnmopJEnoWafO9NowNuG3iwfj7hYO3lEGXHxWOKg8ARzeSYX7ky1g20nw8ajhK0fNz9BOwnVs38
bEkdXiciGuWdz/ze6KvLzOHn6ZRVKZeb8tCcEPSHQqmTK09Tso2w7Vdgy+8G44npv7UrVWKYLQIS
vimNChS+IibzPistnBIUrq4l919p2cQTnmlSVrUKaQSMuO0jbG6Zm/khxMT/XMUOXEsycI/TvVBc
eDdrFsJWjmQ7STKsj/zx4tGQt3fKvsjJOz0oQ9T+Vvy5SONCouMtMPIJNHRoP8U/5Mf3WrYFjzSt
xHyYj/pXiC9w/1Yfyffd0GfR0PfHQn6G8r7vdoPqZKrM1cymaVYrlcUZPLJK56XVPiIk5J43zu7p
YhCOManYeOF6vB0gIhB/OswdL2UhNqIwKPbgeg/pH1qhwAzIlyY4p2oA0DNbzHQgOzBEtnXhBWhZ
hsS3vzMpPShl7kNMRhCgijQxGAuOcSCdW9Yu0Zo8MWXkVeuteKxMK9A8gDxl8NwPbir1lGmdA88p
O54ql/XqsYjr3zcID2MlPoMjrLyjpdCfS6kEEFxkbtX/LryTqlqscHG40dp82NbajY1Lr5QZ/9UO
2dRXrbtbNSGu5fSJ7bCRH8iAXCpl04LH9+yPGUCWU20OWPJKI0VbiopC3Mp/uvOMJNeH2gnJMlgc
nwOBs9ou8cO6cKqLOB6jtNOUYZeyRwO9dnIbtnxhx1i57u3xpXCbhHeBoxwV/6D1DD5ANOKMWrId
5TV0UWEPKCNZRS4nJ4zuSX/Gb15rtEIjXtaeUTCnxs+nyfrY6pPC0Tdq8PpoK5WE1NF4EZWoSLGo
9Z6nNjhXEs7uJ+ggZe/6lpa1aIClo7MZmsm+pajRN8F/wFoanmCMnO7UU8HqMrjAJOw02H3sIGG1
CjYrl3tmRcVc6tPjcbHgTLyrEbckgy/56ItQ3ZknRYaYV0Y6yuZLK5pPMoicHhmJAHgiBFdTEJho
MFdr4q04757qxbh0t3NhO2pUnvtxgj4T7gbxrVr7GpvQNuV9LPWGax42apX3OpZWzAEWJvSsHIh5
ogBKpYPpAoQAtVoytI74ugxbn0E30Uhd+0e9fNyy27nOarXJcg4a6tVps8GKa96ec1A8q7iua9bp
4VeJMqdIPwYETobLGOvIxKCAUEBFgP/41ym33j3NOS1heoYETTLfeHdd82BqWHB0IoBKn3HGax5G
3dVBHzWfYDCyCU3xzDFVWbxyKZ4uxxWphZ0CsCByQNM3LGnNRYg+x6J/ZuQzfrErrXJNOOxnTAgr
6U3Guu/UUldn99em0c7+b4mF8Yu7SWl4JlMi5nN0hQgTzyHZ3uoaeDWK5yRwGqFlWXquOWAtcS6h
ZNJosHJ2sOwPkrSHxCvGulaUm6oxm1g+XIDE0FK/F4ZwtjwXtURn2OewuXxEUXHB2GvSbKAMh4LR
/Vu2mPPatt9VnXmdsDYoPF9Iq78QVC4pKKl9D7/8/m2mYP2j+ZyYPy3e3gCE5MKJrweBFGhrdK4b
2K5sxm7lHJWtcBRb19GRAXN9jHFGRKaOJWPOPyEFdS7SZkB/ETKBeeL/0DFCXyywdJVUYPTDUtg/
VqOOIe1zKLxwKazih/EXb+Zqkc8EnTlz3sG04ygn0TPWHeuuL2Jenx9rAcyqRQ3OwLAfwYXWP6Z+
e5mC3QKBuR7jdOzLY4I3umn/XLUXAh0nzTmnn3ETJEiMfWDhgttuylysP+zLUUADNd9knfgRBMy4
G+7IYqmUEH9OFMWm3351bV3/qNITRlWt3dIo16pcnEerlYWzmeieDrcY2hVv8S5frNjtoEh6Vopi
pCE/UmsKcEZsDUpZJFs6R7rNjhnq2nVHSV0jG4mF4MJC7y/EBeuLYZZsNBsGkhYrmt1jiJtVOp9H
JT/p4mkFVdaRWS9z1OESdm0qG3cVrBbBx1iPguQx7E5gpoTdZ0/jfbUDFqu89aXjiQKLc5O8s268
rhyjHeU7hrLpU+UMgIKdnBYxvpSlkulmf0amWSmI+dD8Oz+pPyDnWZwiX6dpDGs+x+W9i+ZRa+pE
BRVqSLt2QhT4PHCTkF/+Sx0aB7bwlMZ020RO74CeROlPNoX5NZaBftlh5ffmR6nZcZ9K2pqJrVHA
iXMLSIYe7d4LSapzUfhALnGJPmwmFlccKgntaBELePnHZVCA9dXu9PmQzOrvkGNPekzZncjj8Jax
RoYGXGGdWy/F9TdFn2aztQmBclVgCSCRZmyq/J3Zmhj3TVD3RXVEAeBhuADm2EStQE3W9u8Rv+mB
b+86nepSEIzLoKpxQdXBLalT52VQ9yCicl4kgwpG2RXwHmfbgZHumKJrV35Q5BrVvcEFUMcXO2v/
/6yTKH/ockR2ce5edn+COFZg9huQvyDs/YS8vUrnlWeMW4zC6uu3OOKVb5FLjRgM5t/ltcYlAGs0
ThkznJH5RVnpKlM8t+IZXqeWjpniofxQh72Lci0OIqm0smTokUIXdFi30fW5DOcBFrgaN1pJMHrd
nMuKtHvqrxrHhZoJPmx0MZ1e6KYRYl3lyBKRTTYvIgVIK+tN7Iutz/rFFHU7fapyN20y5JjM4LRd
mpbsVh4M3k30q+MKeglCBhWjHSljDHnrRhcBu92cruzeSiIGZv11HOhf7F1JKsg+IEs2+Yle3vN4
1VxsXHvp9VO0HOoi9FEpFX85YjkPTnN7g7EyeUBrK+0p5+26exiKOJnPgS+P6XrKzu7nhLDQWfVn
/iGNPuC1/R76mRPbZppaK5kdlmC2+6JCV5ALoF9p1xlA0wZgWGBbek4jLJkGa/g/5vQSA7Ftrw9s
uEFAUHXGMBDz35V6T62S8gCAZWGSk1UShpDUR8iMfHOjjXpgg5nDCmUZDsJftVTkt7geycLv5YkJ
2XDDyTqfU8eyKBes8nTnHzuWb2FDKXLa9swsKa/ktYSEGsobt9Lc1lK0vYNdOZMdN+4JwmOpcieI
HL6L37B7O+a6ImOCzUyUY9a/jWqeZcuas95F9Mvoz0S/MJIRWSNL6snGPimEfpdxL49NlP+TwUbv
Os7bYgUKTedg2GTZFXE+Dp3LU9iDtOlJA/xVwDg/kY5fGqFupSOv0p5QWbAHGBOHFpQin+2PHOR+
A3+w+Cmkwrx2yF0X5e5quMVDZWIKkMa7A7ex/sFUcHgMuiZGDNZ/bI5y/EiCvkacZoNkUcjDw3PZ
6L7DR8N259cc0BS/iBh5tPGlnANa3CPsOUtSfO9IF78swTpVKR2aWPU4Q2rV1FsqzqcKDD8fEsgF
SN8mh7inD2qlD16ZSn5jisk8Q73dAZ3TMEhIjBT52bEoAUAAYBu/1yiabkmzQyoWP7UzCF64Ukyl
S8zTV+ke8JrNiVfsJduGAG3foQ/a3xhqcS3FvSqM4ceV/M8yjYYQYBBegSci/kLBvuJWFhITnHzw
50mQ2lQzPVASfiXKisP4jHa9IZmDxKmuUxHHmaixZKbM/rG/bfMwLVBm10qyzG0kIB3Y+Yveru9n
eAd7BMbuiNcDN+Zml64QWhLQbA93hKYLxPBRl+m8Ne772IEWYJ1ELXWbc8iKqlyFMTSGqlSP3vej
UacY4uNDKtsa5cPIzS2WCz8Kg75zrsqVJW6M6fDtd7nHlutbyTw1GXm4rcAH+72jzO/brXg7wr9p
mmA/byi+eVDU/nJEX3Wpa0+1SeiT5TtB/TKKMREfPFMxajH23C5kspg93HI0EcIimP0pGPdOL7yD
wzYo6xg5CrWSmY5/P6VVhidPLV5TVPEMFN/7Ipx88vIGUwldIbtfJnxPd3U+X3xdypQ+X7Yl1T/F
Bs4GFMxDl36Pv8rw80gv/fqXFaXi0kYss4J3eqgUWKJ0P+58B0desjnVgkskoogb0Mq41e1Lr2DF
5ntPIbvWxLa8toO3oYnfZBLZ7cZ6shmIO0Q2yoZFgV7/chqV9zLRPKfGMZ3PI8kCFjojMM8Rr+fX
KByURzshLFLPiTrMk3B7CWA6p9IfTGr2sg1i2OzcuHdkt1ymDxlk6+N8EFF3WdGyt4OYyf4HKymG
mtI+mq/cHQkAm4M/bcixQ5iRv7iJuOmjc2dqFfTvL7VZnXYE+XCO124FilT9uRlHV0fjTUHHj94n
TRnylrmjY6RUieJQO4OboCGkt+MrG1jkC1Am8PL458nYLDupfb8r7s3ij8RFc8mkW0x7rZSfd7ef
dvYL1Mp850Og+SQ/478g4bHgngZgHy3uC8GAxPepc6LQXnBU/4OmdpPOkfXUkxfFzmPg+cepwsCd
MMuqXcD8aeYKTZgonfHwcEsh2mR0JrN86X/4yOri8AMnERgHaz596HsrqIgFJyQ1Z0xZuLpryswH
x0sFm5sDKuBe5h6JfY+/ruDHHVginQGjVgKEAHBvn31UNgrJsUzM0zFbVjdm8+q8bl1DsZkCT6fO
PzUiPNMrGJhEgf3Ba5KTKfwgmu8V28iy6hNn6XszXMt88SLC7uaTQIv8ZDKDFYp/3R6Yv9rLA8x8
UZdaK7KbLASSMYwAodr1SHSxVIqstV9qYPtI1gED6LJFqvsqpISZTyeOPHFV0ts+N+tcGpJ9oSBN
zScQSfQuthoKZEysjhPW+6W0qty+BVYqKL33K05EkmN2gXCTugOawudUl2e4NQJyJGUuIbv7uIPQ
20pJYj0wG/re+kdO2agUGHpdid/88rT4cnhl4nN4bhZYlH1gxQhHBpNtAz+/kszlrCKQo1eu3cKO
ZOcfEvsHue6MEdUi3J1o2t0ty2zaSr9H6attFsth1qiwPKbaY/TLjzyOH589RAu2S3e0Y9Pp1q/B
nwV+aR1JUYSIeyWmV71bR4lE+NrnCWd3XzaaRkRdvCwHddlBxgY7GcEcCu+3vJSyLNJfXXkWsi+D
R99R3BsXwoNdOSIXpX6HKvUyMG08/JeA6QIMTXGaKbsnw5U/P4yzAzGnC/QZUegpIqhE5+hfhZke
pKfo1WUWaxaO2AbVHYokF4zsZise4VD/2oOyUqQhMJG6BxYFsESjJj3wcQmbN/NmPTP1UwbbmAQb
BJMPcdpcMCnB5X2ARob/6hA2K3kWI+jq6swUV4i7Po3nAyqsPNSEJs8bfS63CODS15K+IUldsu5x
6Gvuvt3lPa8XH7sPOY544weOD4IRAomY3eG0TzzSnHJwF7iyyOrS+r1MBrCPUpu52IbNZ27WLj+9
zZJS6eoqPdzftDSmwZxcC9tD7Ofx3NKdZo8EPXBtY/nP2Hapuem8Ai1Ub6rdz5dgZ2uD9SuMchNP
yvgiNfBhz2Oy+bLkzR5G1d5FnmjqM8ZVZec+NcpICPl93MzQ90dTcMe3YNL0Eork/vAqlXOF70a8
/e6e28/XejQLo64gZknrwFKgAWNWkahBWTM+ELPp01bxLcBUt6SvDlSj85jS9pccYtKve8FUsj/P
1KXaatAHPEWyxoHWlCgjp4D7BQHSC0rf26mfb8TKH27wDTARLrCAjxKra8XMarEtglVhCe8YpFbO
VVjQHeyuz5YxLMGDg3z1hnKInXIUCxotEJRENVeRvvqak2Fm8bfsh3924DEol5TuMuFIA345be/2
y5GngctGGYUdDODxCw+oKqCaZfjYlFmwgs2TPHQTvPhsjUp9XjcARq9Frss7nHvbfyKue5ezYcTx
wJSsQdr7T2I90FpJjwdifk61SAE9pGTwNzZ6YJGDuqbyh5Mr1smGuXfBTYhnKz+Of8TOok5NLmoX
i4lYGytY1Ofa5Z7U2EB3ZyFyqkXIjGpcNeufAG1rus6LuYJZ8je6UqbRxx1J5DG/yYBUJb4c7QIk
AYz+be5zDcbdMr9o6a5HBEc8zEnGv1NFTlS0cGSPlIak9LsyaG2U5gDOlHmFZhh0vEPkYjVZSEHS
HvLHmrgiYMsfFDO2iqI+GYuFWhrI6i4fLfUF3osAtwY050XCIcxQ59zHMobpQc5iqerJep+m25Sf
xHLtTicSIBv8HgVrm9BWGhM00bAvCmiwCD622GuNPif89WiikZf7txFBwofK6m8BFSzX4gTUZTnR
8XXcDI3FXQJlbgzcUA/rQz6GcUMKIq9tr3hv99BAGRmtwrcjs1G7fhsj9w449odJFO2rU3c7dby2
+O7xhjmmTUwRV33BJ28NDiPSk1CF6jVzvyz0Syrk8qYqt2foRRH61ncQ8Y9X/yHuL6dSZfwVmohS
/lVv7CVKrogkHnnr5Flgti6wiaufQkGmuMw/cnGXRSrDfhyCc5ivrHl5EGgoTcKZMI52c9wV0luh
bS9mGrRXTTJem+N2O7cG9Fl8Hq9L/wZhAWlNhRxWmh60/XBwk9WtTRnOXcP6w6KxmnUmFvZP9EuV
ZS/4FASt2Hdp4/6NTsrrlEUcqEc3kicMkWPY+6WKvBu8h0KjEkmgrRYLsI9YYpiEf9OfobkkUroF
feJ9rOWRjbtt3IoWvN0ce3WfwM6aYgkCngK9NEr8bE9OyzzgVVXsJorPvv18AKeq3uRGvu1P2fp1
u7E+WBA9lENm8hAbUpJuOS2LIXYzizZKK2hEBTN1s60tEiuxdskmftGzUhyOkh1vB8rNOCnKKpKe
7dVpchRIzrlbFkeXPzvhKM45yN12xVS7KvsWP15inLEfPtxWPt//L9LxYIKADVxfsmuwNMswoYz3
b7OwQv05UlepGNrnAQxnm3K79Gvq0Ee/F1o9sEYHGPUXqpIg1YSKCQvhbbTjrowHaiPszYt1kdKQ
mzhQVP5JobYrtviqbkv1HKQR2RJZokhAYbc2EI7/kMpHF4PxVy+UymPzOwlRn9FQ9w44ym4yiXyI
gQgE3DDyAnUoKQJAAlABO7JBeEa1W0JiC6Jw93iKKLaMfwgEjmKiVhOMf3mkeMgMG1CPJg/LcLIX
vVCtwPMea2l8k1MK1IevuBOyYBd21+ubLeJeQE9bMP1paiLjpOUQs9G8WoALOflAf4G+rjStqFQq
DHNTdHUe1eYftXyCCI6RvyexURjR8RG5jWk7fN+TIJa0jKxQWcz4UIgOJQ73kNQhencrfGBzgdep
maKAtkP6g+Z2A9zKx5+OnY+BVx+DkkohvgwDeGoq+GX5yYqiLCVeu1UCp47OVT9sfQ7FFmpZjgP1
cB+OpyP4FhUHkqWS0qnnzFiwABqJrxIyQxtjDP7gQ/TKkmfsyns3WBwIiNOATSbGoe9TQxZWvZld
Q8Q2uajD21+g1W3EOoCkZU+V2TDs48vTtTvRl89aNLHCiZVrrs2mkh5+R5a4WbQR2D/rzQO/FKOn
IAeGnu4OqwhXGf1Q0e73tgh3SpgXy7J4ieJdS4Fvs04Ihfvbkpftyj6jUD488QASOz1Yl/BG7xB/
ZK7hdohej3HZdu6BNrJ0Yg9kfNNfMBhUJIYL02QJz9TGtaN4ZIsXEK/jXwriFv0XJaq70/RIAAs5
IFfUEjLv3S8CCw3QOpf1V9Z6JnXQgVt2a9uJjdJICOuCQrUHhxini9kP6BmATiZc6sYG5OHQ9B5r
Ru/3NEQqp8CZZ0+bVx34N7zjaZQHYWLXFtze2cLJR2JDY4GayV558lH0svUBq5EnAdRAWjp/hHej
6C8vPxJZpDRbo0nmolN5jMrJw31prWnJTL6YGjheSrTW7UWKLZSkxG3i0gPPO5Qu3LfGOycfv0cj
7PIcEI1WYca3CAYDU+SJVxMb/aUhxr0o6/ll1OZEeTAPURaE/vBXOdPdHlOxnZPvW3i3hX54Nt5A
QLDATo4CG/XP2qAhI8UtnaPdMWuVJoSR8I5FQuyZOrucvRwB5cSeHxSMA7wU1/ZcjL4kqF7bLvtC
RVjbR2BiKhBR2n6FmTdpvIi1VooZJ+t1MoSRMib9Tikzv+mGNecOdikYT1nEp252vefwVWo8OWKQ
jaPZR+ruOAa647Ar9vzgNnE7mAkVBdQB7g8uZkU0bYvL6xQkRmd9ma/BUQQ5eMYY69D71rAQISTO
eRuKY7QjpyZFTL6xgCbfalZxnV5nO7kaW5B8nygbc7+XlaTD9frfZmjh9Gdav0hbSYfNBrTRU/Dg
ebZlAAFxwriJ6G6o6ncmykgaQHdnYiXj0MTwc9oNCAHlIKwhYe7Ymnj7P3MaMADdyi6tgDqxt4oK
SVUNhMSO/dFbBG4qxHUX6C/4jmyCOJayKQAZct+tqyLHA10KaH1z6tRJniTnicK9CseFdTNgoVxO
diVrTuUEIHo//CLXPkxWicAQMwcm/rGCC/bgsd5vFkCRm4JHNW6W2IMrXAQeOfTEqWG1LmbxtN0h
1gPwgiqqJBQwOEHYpfn8wjwtEhwcUCafFJ1adER1c7H4PpyzcgdukR+14Edo7BrJkmiFpD9DhEvt
D/0NLl/Y7qRHj43Eulw84oe2yREpr/tWy2UaBrMFFgWtObTasLaAmxU1EHxf/gY8pNvOqoGJFXk/
1y2sTaDri37GjUhB75j+NAwjoi/t3aT1QyZW/f1Yrj7bJF7CYmAe1l0+33c+3nfgtPkEgOfJpoCx
Dz5fRB0uyYnJqq5Ksc5dbKz5seOiHiDg7kHJU6j7YTtWsw5M52YbJQd2AEnympLQ61GejFqSP810
Bu7vkpJt8ihA5PTkJqLz7Jh/Tz6U+7RJvD4VBXANsHmORJM2OcQn4NAqLAgw5fk25WMzGqhnYqWP
dU6LZVE+lLLLnVtcIzGHd+D4xZio/+nvMuSZOFsg0QyLpWDZBzj5hRG75BNGOihQRyg0uDtVyErO
+DkS7FGK4klm90KRNjK42AGeTpc2eQo9FuHyId6+I70URiA4Aa0DTU6FtqTSMNEIQ48/RnGMarog
jGUBz5tWC0UpfaDrbI1nldksI2yOwWW6bkqfIL8dPI+4PSteBlaw+sfbMbao7BcojMgsg2KIwZkY
0WwXBZ7rENrhqHIqLF4iNy60MAYXmgpuhsCwVI+VEGwQmsCTsS2LIYiVf4xZxvI78f4jUANtspvC
n6p0u5+CQGJcYxRWOrn9cNCeK9lTAoC7ZIxw1o7bMsyLOdYlr1u/TSy5SHqYuW1Yy/lhgqsmnyC+
oXZqYEEd9dDXYhV95TLmGM4+aaJqEcyOtKTM5jfBxcdl6c70nIMRalnYU/CJq0XmNBeGYyNcAdKa
h+wBOx+vw5I5YCsh5wHjUFdYpkaTqBOZ+pbLh5hp6Y9IwqkyADomcGNH0AKqWCZjIfuuYkuu/2Qv
D78cwdnihyYAwOnN9hG7NDb2Lc9r0gZHsHvEr68l/VNSmEWXY3CpFAStwwqRZC/gwiTVcIkS04QE
zSfikZ5aOXOY4/Pr44dY10KJg5vMLcUP1pDty+Z0Mk0RPGuIWEj0hpVO7Gk6UcwgGiPscAgs5t6K
/LrRF+nim78/liozdv+Z/4A+PlHvzNL3Wb3+1wETEJ9FJhvFPuTmRg5DeVjcbxqiHfPZUHo5xAl5
hx+SZk6gM5e3mNFxfca4EMXuLHKpXgsoco/5tisIiFNdl0gs/b6xd6/Ihundn2uEJp1XvM69eJvk
LylHXGHNahIqA8xhJQmYCdQjM23Tv0uMxy8JZO/jLSmuVaK/Ul0Xz1Re6W5gpFemjqUyllgFZLhC
ve7ORoBb73vWBQ73iuvDY5jQqDLTHZ2PpQiYIRpVE2+C5TwirgUh57k45C7TN7d+DRJPg+oHjXd/
JYf5hFPX47EEA4DpA/Gqc15PYNy0BhPkfCse7/qGey/tEHYnPrpzSgUS2tZTxbhWH+dPcCYjNa8v
tENI14hLoiBoseusOe1iOziXHUWG8x4BHLCEeFKxXIPnTYbDKZrdic2Q3FW4qLWsYzoeSSMG6p/X
j++8MKiJtzF/9yCwhZA0Q5LHpSK0Qhq1/9UCwBx3/4rkscNJpUCmIPP1Uk96Hxlib+Z8bT40MfZx
+o23Lj/Z5CV6PtmFL73IVh5/WSv/ajusmA7iLMClJ5ADdYfPehVl843E2NCxTfLGxtOq60vP914h
q70Eabr66pQT7vl+voeBGbRAoQ8GmMmkYt/UlmMfOly/JBBW9EMjTVsIF5vDWdhRtRZQejQw9QSP
hDKTYkeLp3/vrKdg8+Raxq1ME6dITqMBX+t+th6iqeewFY3Jc5sW35YiVeiYg2PZSVjp2Lh7j3Ml
qyvx0GVy2FHEMXotOh9BtFhQHhfdiIKvzVeAfh487mvjeZIUhSXROU54g5LTyiV3JlAKhMOGYAfe
8cGQRTyLVhNhrghXI1zvvn9vUZIZBAXhRqJXErvoI6161LSZWvFi0oSIY1yi2/h/2FjBkDkGX6p8
2vHynlg9oDr76EgHCDOLdDe5ApB3wjlmoq5Y2kB7CUcyXS4BmMBwEeYT6mCbUOZs8+ZNsROgvqBy
pyywqV/wRtak+5F9xbq6KWvvaVlCPmDD735gb4eJXdkRxm+NauNXh64RTo5a/v7zdo+iIJPpAnOk
LaAVKY+KRazsyyx5jZdxgJz8qMT4H7C40zS9uS56pSjzPz9TB4/icdzMpHzkdgVqvZb1xjomo37Y
43WLCG3O3ap3C1mn9Tt7Zzp92F0KqTAw0lbX39ZQcNzScT/JK3YxyCpQ/TBGejqR0onDypbvL9tj
B8P/sG9Ffss6kWJnrSkKUXrF9ldvjC5MOqPiza0ocv3/9r+Go7dzX2MdP4ACvEktECVzrRrUUu6l
vwgxYJ1DT8TiQSgYO7cHD5r2K+bJLB4WZTju0p5tFHUBZ49Z+h4sGXXPCy1NZ00zVd8iRdNQ7d3B
0qAPGbFbDppAJDSWrn0fAnK+iNLepJft6y913SprbNLNKyiQi40OTJZoUUBNvkYZHlV37sc1GC5C
2PDjBBCYeeaVtGLXG8e4/Sdp5qnXuKf+/K7d4COIDq5wVn9UpVbXJekGoCJxw/LO112hIkqjb7+7
zOFcYgQHhc9Sxxu9lHFVsUMooCIN0YD2YWztY797jjdgcJ3UmQTYQdcTKXkKJvF81XleTz8iHFEw
Z7BBpxJD4xjrHd2b79V3FhBnXHR/t9jDT/1+CWHCYVl4d7L9+5C9oXdrcz3bKzDWgzf4R4qpoNzm
XFrwAtunVLCPSbWFJgofwSTAwaKVzM8btEFWw7s/86c7O65tMKOhLLQbtEbhuvxNuDTuDH6YG9fA
3+d59CffsiQcWiH0/pVotAfnzzOuCpOOkScuQ+GCBA9CqtBrjOe/mTxP2CHLzvPur45dRBaswAMH
2Nbf7HpK0DLl5bJ7z3X6kZ/FysIRylZO9dqk6uRQUZaNJT5KYQ58Tf8vybFVghXjkBPiHYW1VJsp
BiYJY/O0dX3hF8sGdUJoCDUfPzxWuBmE0Mq0Sna1fLZRcIJFejQ7xhf27n9mOqZb0SNLSi+QusvR
pMkLdEduy/26ysZ9VIgI+k644GhXmfWWzajHaR+lfZHosH8HUkdhHWokvYJj5VxUFdl1+sGp/VnN
j58C7Je0T7ADsBdhZ9U2SA+khMFhbytcYIyBK6nqrnmhT6wHHRLSAmpZP9USkkFvADBhspBsM7xK
DBHstTOLapWTVmZL0sWWSjXARyV2bfHUG9yeqwwgrjk+uCxh6YCF+nO0w9mcIn2HYbkbwJbZiKZj
O8iSgzOW6ze+y1RZI+vOAoNIjKvpg2N6/Co9cizUIN4IFPAHu3s45ks5fFj8kxFzZWD5QcRV8GgS
9V6xw+eCvM6oIeHrkGiwN/YBrKRSzpCn2bhYydq2ZJXylRZnxLKsZKIfAzy3/O51SRqTi2lILIT3
ZJnLiUb+yXjruGmDk1yxizE1OIklP1cDutwu11h/rqwvj3ZI0RqKm5BwwVO+rUpQVko907n/ipr+
TG/rfc9n+hBhLOvv+SVfzWmZnxr4jUXYiH9hdQZusN6n2NJMD6zE41z/jwGWF8Hp3HCMy8c2uy69
zO5OIkY3Op8Nv0/86eA9FiNrmukOBFmpqGw1NoQnK7gIpXJm1gkJTSZJGuGO14mFYF0NZRdpvjFr
R7S1jy23nzjQ9zU+k6WcfcPDoIj8pMm1COwQqxFYvdzv+YLgOCw1dgLwmP09lSCGDke8sdCwjlI3
p3ue7wweEuqSI8MnrFbTWtQuNe5rlATkcXQLKB0CS3wTTd5U9Qc956ZFGRCa3Erk22TfV66xSjRm
R0rhJ1g0tUGijRyXv5AEVpqHiCzjVJvpuk0xjPxlYCbaPCZ1zkzPM1+x2Rmlx/QqCgaWuTdY/NVC
w9bWJ0wK9XwITWFMrF1xoDHDvK1WXUsVryB7KkqmY9Qwhgj1Tl4MJKxPTZtkaHqfz45Ja4y4Grfn
q2mBNhUQ4vMUnz5+pN1DWubPezjuf6pNMOU1l1IeRJ7gNk0KlVh6ka65ArT9FU9AH8Vlek+DMNki
VzxEG6nFxmyYY1d8CoEwxafWXPuPISdsi1AAhssgF593qR1WS7J9DiU3hItRIkGOUQaV4qASk+zr
bGSh1aPk3Oy7vTPmJs1Dd/5wM7jfWZEagjUws8DSalrrUUymDojgHvYXxCojWekysrt7ECBkP2KJ
EA5HKeoBC2LdGdB2FsJ2UXuzUIF17tDlxJ3MAzi7ShzUN2wl9qGHrDK4U5Txcs7kupAWts+d6U6N
mqRC3OoQJh+Puyy+majdfvoiBWYrrIeCysF/2QWoKhjcgBWa+xoED1X9qDAGs5veKab3m9KYUpjo
aGjfa7vnN+wsAIMMjhRKbhQ8N3Co4XdUMuU9FDR3bVPVNd7UW37KWQmyRTAtqmuYBeixL9OiGJKb
tfWGfo7PRs8/Z+BNkTbafAMFb63K8C8G3JljRrLC2g06L+KpO1uLWA+/x/c1xcfWB+q5GTPgsMV+
79uV8nJbp53d+72gIcw2wGaUP3QTC2lz/pAcm56JFaBw7QEDj4d0vBwexH2BQ10xg/1yINdLc6Fp
d7fNL7o1cjgZgEsv8BLkO0w+/PPj7hNDuM4KqAftet86Cej49C7xLcFzxUvjRmdu3ZaD6NkSQPvX
amcVZjkZS2fmeJ+9weB03GHVMhhcOjRTkmsI6tufH6aUOfZGlPERYQxQZc5eWpxat7+6I7R/P2Ot
fv+zdIZXISHpiEn1fhyfHY0A2ZWWf6loQSngBKZ7ptoUIdJcuZ91pxr2LEVlS76IfrqsRD0Kl3t+
4BSzevESnTLXMBJ5PxCJqjHcz36QLLRULJj1lyyOzRPgMHbX4Aka8UDM4BfIIM34dXT6w4joSs7u
R6KbgeiVrR4hf3p8SpzHAvymLi8/WwH3RQLN6nT9Ln6bpdwVHHBNxDbEpn85fcJEF/wrV+73xbua
s/mxi+jYqOzyPxIJZ5CaNXqvGY06psd4h3dvxnB45XiAwtmFsIgnEw8SgY1B3Hog6+3MgTpuR1PK
aeDWX7q7t4iXVfXkYjc3MUHjer5YwfdetKqWqwgaIPjwPGtzuWcALwzdcna9cTIT6K5NZyGE03lw
Eg00ruBd/AIRtYIVa7jPLJKLCT4IQVU5ZTRUiWFPTTOEyBFaZ+ktd99TuU4+ut9EI46d0eOmbK40
mC+DReFmvbcK2juqSP/IaPkqWmFrPvhDsuy4NtLZ1E0K/SrNjtKBjM2w2Q1tfNYmXbUza+Ww6GlW
36fCM7299t0qdWFNgKgmw0xgMtrkwXVfsHuWkfbZ9ytxhMovte8MJFE2cWUKxFkABp5iDCw+B3aI
34LipXynsfjYrdi7nbHM/zzke3QO5QwxinnTUq2fLaMcyVhkRhDHsJ+EP8aEPZD6KJJ3VdkQb9xx
9sumhQ47YyNYnO6Z9iLNu+XGruEiRvBqApWx2FV33xTBNukA6lb9b8GqNOy2nw4otsaErymuWocy
+Q53aXTnrl2Buy/eMpxeHSi+mfy9mmc2PGW6nvpdyJhpeHsQPN+MC6r4dECaa8SUs+25MSrz8fOP
PCIiMsKjXUNbIoN50AF8EoKGIaohWTUhWai4Pqcpszqt+o5ODIUfF/hUsC7IYTk01W9gPNojZ9YI
xuo8Nouk+HQY0ZHRSf6uxeWur9NBWGVUQc5leIzLKMUTUvKY9wKRC94wcizAwgX63vuFSaqps012
DPkvsR2Yna2pGU/hu6m/AhAJJVP7G3pHyYT594xL4Pzj7rafXLiWUBfL/Lff1yUut6GXvUtsB+wn
FRe8Jz8CE1T9j+oHRY1EGfoi9RQ6GZN+LURsk57gmrPuN6TOF8nr01KPeKX92XPj3RtaX5E1zOKA
8i3MPCCRuhDNlyGwZFu9kwgeoB4EquMKAvy2xbVVH0e4YOdnlcQrtGiOyxkSvck1djJgEDJplwt2
AjyHy4DYxxfHOhSj8j5hf5MM1F1qmEDEGILVimcOc8YhGonlDtZIBIkFDOLQSKcUPCQuZ9uP7lhj
dYeAyvOl7jGjWJt81piRYmxrp6rg4zq+ptBTYJkNR5qDm4Kg0RbMft70NszFKtKsD/MqNOSPVHUH
0m7CTr83xj58UZtyWnKi9ooBBwJ8akQUHaOxmpJIP1PzJ7rmf4YJGYS+fJkKEbaj242J+kdqCSdn
76mrvr4gQ20mpmz3PVhVJYZe1sZIsybuQKZI/AfdibKq3bjHr2JC2aXoLGX0JWdbziIVMcidgKzN
MAVtIgHZ0WF+Pj1vdglTzxyLwkWM3qemBiOoRtEQIpVfjwNd420YOI/2r8gm+agd1NG9O1Tf7iSb
lv0v7I9dTX15kQnTCI5Akl3WtXIci7UWph9D7sACgAboxTvfVfcLkUQWeicDshyQeNIsL+A7+wM3
VT7rj87+BYkgGc6LKSicMTHrZd4V+xvxNAuvg15IPBD2BMNI+ZP4YsjlBXf3GE0aBlpG2wQkBLjg
tIR6Pt+YigtvDyGlp15OHtfn+aF7HEn/zLmeYX45b7YhgpPFE+b7F7lqA984CgROLHeAHNPdOLsJ
5BEXmEoyHpsW0xtQHRwjNx2icXdXgib9/yudP2/OsBL8B1iDZGL2VY7Xc96okgbNuvHjMfy/yFOB
TX+MpcHE18UbpXuGAojJM0CBQSymTAwVurrZyT+JtU7LwyR6JgDj6pdXMoBMohPwQPTeSy1oB/hL
tpCJvAB9psqRtvL5zWofRJt+8Py/zZ05J54g4McT7oK3BvuCgZHftxiyiVoyKamdOMrQKRlvSnJs
3YOrDq9AKo+p9OZIejjKkgaeYfZkChXLS19qDJX3joW7k+lXpbHyPZqdtOvAOlASTwkyeK25PUWG
e2R3OGj3tYIzJtQ1vrIT/c6AamlgNV/MM91p2qje4gkKyzwzPoctG3/Us7GsCiqRpIdWwiRVWBZI
D+vo71VBdD+JHBImLZuem31vdNFQx54OJUiJbhpMS74Cp5JugrMpRy0pEYTXecQ6s+OgsRcGkh5W
4Q6/4luxUkbskEbXXqDpe4NRKk/5gp9kzCXBCgSDB0pd3ppdc8w/k6HyNVASelBxT1WmTv9wDVaH
m1x3/5Uj+o8keuGS5ylxavC+cDgxO1PzFuaYJi/XxBDgr3B7mhevxgnlpCmtGTZh8pq+lZyz/7XO
Ijqs2RVT0sETd0Ea/MD8lSghJwKkMo99UJAaJ/QNnXUXpRfR3OOw+wcIaWw5VowZXI3m9cEXjnBr
ZvQp181jdsX8K9TvU+8mPfK4NngDpSiP/U1kFyAMTWpThFuq2b8XYy8OwpB7uq2V6vRgIiws7r0N
NlFo+yfJR35iHlssO82KLKNNtMb+hogEvKX+M5VxDkfKMZp4U4Oq1iknxjExyiPwhK2YNZCWP/JK
Zv8gW4TR2pu1aUnEcTktCINvlmKtAdgiUoVz4Z7Nq1MwaI+FFS4C9mt9yrm0Or6h4GnT00PDdBsC
pmQCttCdmHSS7utHesvBEVPOYWYAkJ7N67fGj2HB9T0elOcMOcq0AjxDuWYIaTJL0Kn6YbChcrmk
gOOVOUduDzKru4aYHnNPNJx9qms9yN8z+3YYbDueHtOqws1IQTnssEQVH8qLrZzwkzPVBh+9oMtY
orhQ+FQlPezyUwlMKsmArSiShjBWTbr2veWij5iurFHNNIfny8CGmYigdUyBCB6mK+Nt73L+dsGW
l9YQiyXt86xbhg41E/u4VqaVdSj7AcV/Ql3YovCfICtzlvr4P7NiD9qsvnBYk6hqS0VNKozabGb/
MFQg988iCELutnym8INbo7MlYk5cossam3wI1C1obNyiQFUI4stsGf5FBck+Y1idc6N5+gIgtAxc
YpcL1Rc/0KTI8yJZXvZeK1WZiCZSrApW1KVn+Mp4AZJlTnv1F+r1lkO93CVuSghpAb+HDQ/v5iqd
BSofTozrLk8LPelSbooUSQn3SoxEQgenXYqAmj6BXTzGnZRJG9FEUgpIHr/tZ1vhmjFMWY0fSCZA
g3WeIoXAOy5bcf9tPKvXPrJz0vhU8RZS57Y5IS99GsC4KvC0V04hQ/T3lucyd7uhxOa8rEBW+Ds7
6RlJyKOdORdEq3n+9wh1tE75UV7qLCEChr1tptecCUTVnqoM4/vU9aMO8kAg/IwrJ377X/nn0wEI
umLUDbTg4luPwdQIUkou0aLE0YpRw0SBWl6ajf8f3ymHGdtd6askgpObxtdB//qS4xzHiCjSn+Xw
vIj0utytUgBzgPt6vbEOOzboteWsxd2sHOXXqXenPp1prOPZKihV/GqDssT2Baf6AllEOhURuFJ4
tuNRAyPrTajnhu/472DIUuxJ/nnSyG/S7FSxraC94aWVAPHCjOqz7zM5cXMVNpzwPf4PM7bV6Ffk
sr2skZzxGD8ZmjpM0UmQrzeKXAY0kjBNQD3A2WSlkFxjMtE8EnWd84fxkkBn53dFyvumCco1qnPc
GEDVLEuZSfTVe/nrYde084mvGn4eR2qkkK/ydvlA4/2fCqt64F0QsiH1H4yLXoIgolbJwJPUeVJd
RIZix1CkK2LhH1FT7p0GFaF5xWH6atVQlWoKTtXrEoxj2fr7hQLlfPf9O3oV98au6uaUucEtdOFJ
1HH1QGrDwT8rhwq1EJq2uw1NzB5+7fm3956AGdGoB9cP7djk/dAaGMnma6TG71RkT7O1xO9JWrk1
Bui1ehESGt97n0+CNE26uD1c0EI+LkzHOzZKwXdigL032amGpoJKEKfd8V1aki5v8JOXlyDdePAw
m07buwv9yX3wE1NEKl97tY+Ln8V4XaQzlTYPikK8kKwD8IJQi/nUFtuoQI2MMmHV041R19AyZrph
kqVwylAxdy/dWGhQJ19OPdIEafw0Hu4b8+o0CFR6dM5RgsIlHovsVcyCkw7o+CpOfYO4CKhvlV22
wdH67fibemhuWX3AUdxZd/Ix/nk9To2ugBYlGcQsrN0WLjNvM+oox06wx+x3G7LsS1UkC40aUg0r
3KlivaSJzrZpeae+d7xxb6fUhYWfhNirfyeKynxV9jmELz+htmzyWkQi0GAaWTHGFtZryLz8e3CU
HoQ/lP8B7wrLwuOlcWQWZmSCHcU/gJuyy+QGcBgtMBo6/BnkYo7pF3k8lPu9pSfNOgwQXkgeDlZW
D/7FY5H4VVrrzz6iU/iMt0e1xA0fkVIgwSQiTEMJ23mPEuQJS9tOBuQIwwc3/IPZS8DcoZRXcpVj
lSYroswxLIHtmbTj1eMeCUX4rEKk46ZhWFUxoEQPSAW+CrIMa09AfbBqljlUSFUETAgrK4RH81AK
Esa4R2lBFpDKtnNC6r4H3GylY8Kn1XLryF2e5HtbRP7fp4zQ1lu1Cd8uQhM6docD1OF5hLLWT5kY
z3HIbMoqHAGucFC80CZXqgFOcKBG5gaKUgQHFxmfH+HlO2OmsyoktLVcpdzkCPMRX6bdaxSv8UQx
4P94lEsS04g3RfAyqj6RYZShQ8AFpllayOgpRO1sDxIo9qhJaLKc/6abjWg1xmiqZRlKpZx/qJnk
C5RwgOlFcmrD0CbglVSz9MT2XiaRARd/uWcAkjXJAsg6Wkz5mS53m1ndnuZ8Xq1ABTIrlXZ7NwLF
RypgGkryhj8ad6idpQtufNGQA3NsMSsJVhR/XH3aXPQDKo4f8UaCdlLxHAC1bgRbOP5K+kh3nww8
RcZccKcvDGENMy32Zhivb/do4B+KY0V/d6I27QItPv9AsI8+IexkQUdAQZETdUPA5oxzD5laEoHq
CvuPD7Oja+jheWtv+Lul1xG1SR9r/ieM0l9N2fOua4Jt/ZBpbvXN8is4UuJpfL0cRtRZUWBow5hG
uPo3ttBG+UKdr7MZ8cBGsxFXGWnrQKhb6KypyzoO5Ug6BS3IEaqT4M9KjCNJecirQ0DzbN6E0w/o
Lo02W8FR9pLjGz9BFqc4LlwvoXBFbp+TLFL/p4ibA3TpuGxQFLBTE617bygk9R2hLMzyKB6ydg66
hYv2ctNubodFyXZFSUA0aQIL9yLDZeIrb/KQPhrWqZJmREddNJRUvVykHr3fuPzqZZhbWFXcCqBX
x2Auzxhby3RpPvXnGfuXABukUDf1YPMkAj/R1GqDos1N3I37oH7+TbrkOIEVilybBhmYjRXnGexD
2Qho9D66Mb2km+kESndpe/k8tdsuxvzg2jMpqdinkJsOLUZGwlqyD5EeTeb62IZfae038QiGCLfH
27MKxy8LTaJCMCA8VowTPMRcgNE3VwDQ7FOOLYEwBHprMyO1XKLXikWHisEYOPOQCAwstPkXxKu5
CFfkeW0s7ymHDS/Jx0tvMxya7WDKjhhWhbFrjhO1ClxbI1fRPQjtbgteJFIennB36WqxpCpyb80j
mDpRcIQyKaso3wlIbXzV7NHoV5ROIFYeWHQsZR/H3yamGC9f0nw7sI8hZx+D9JIDB4WBhQwwXO62
XmJ0vtIybl73bp3c+76AY9hWnbuGYLsLK4Jql1jeRrf2f3Ig8HmnVlfWHH5CGUqHLHUCv7oJpGaa
Tl8wCIrpkbki7Riq3PVnLO6iS2RWLUv+6UEb/Y61LmL5T/7N4BoRUN0J9NRNhCuYGyLvrD6qPmcF
pW0FH5wbCZUty+PNelnhKLu+9dpF2w3mLvFdfA/++UfADhvk7WQMLuDJs6BrL/3jvypltaZ1b3YA
JphRvaMiDdJ17Flvy/zWabpN3n2Y/97Ygn9F8cWJq1NrVPpOBrnxQNZ1ft279g1aUrsGCoviKPHR
nZYshKYsDLRihFd+QqUn6vZOTHEIfRPiVxBi/4Z67reyQSIddkVRfNP4ZJNu09q5w4mpMmCcW0Jh
/EdOEcdbXfwm0N9k9JJepuVXuqXgLU/W9DAcMYPVHAMU8cnL/Eqx9fBIkGmVV3/gyPEvFLGiNAo8
iGZ0j/dVspRx/D5iUetFZ1AUAqctJZnlB9kS4EBh7gQ8hYceDc5FeRpwYGa8WAB7I2cwc4pDogIz
ZI2GLyGdWnw6c1ZRoseRQtODGuNBNlTGD2RvY229nDg85mOmRoqDpSFOQP80WCpJ3VoXqm52uuic
OR0ta35dHDJo78c+5xaOdA/2upf3aF07yRUwpNOKtJEU1ClisC8eaYKOCtD1mhdlbgcyBpYMIn1Z
0I7YiTry/jpqTizZF4D3wyz4H9K50Gr8gREPfyJllQQYSRXCHfkrSyaGSZ0wca92B4TIBynfOxPQ
jhSX1vD9c06FZyemFWEWWopJ9aJ69bJ1lz0A3onLjJvr119yo8ZcE5vtgU8/0/tnFpzm5xyL/dDi
QZkmZflgiC0kx9FCYzYnc4fGXB/TH1YyiotRfNW3/aFWaJRVWYQzxnmqpU6NvN9LsZkdxTz38Gg9
RN7rQ6zNWfWwQkEzDS8F+g2An9WJ3edR4dKtZVI7oJszWa2synCaOerSRXX9uLjqGEnVXVeIN+M/
6u8yYSL7uXi1Vep6nIAUFAK+/wOFqcrJw72sAYaiNaOOw8nIuu86yO0Z1U9XW2msvAzYar/XmOKc
bLLnnUjfXDjj2xJ6bMw/+qns8C//lUMF+yEVc8DQbVhX149KX8Bivi69j6HuXRbdurtihKHMhwHn
2N6LrQqvNHNUP5EN1CpLiNLcpvsAa5VJq34S+MRMJUU3GIraONoE9X3BWq5gdlt/XFK2SgSYEVOR
QJGvpuDLlzPnFAKTQN6Hts5L3DCoFI+6SvDJeBKSJ+UvgPVX0QBwchjQo0AIbBejZGiT/aVsN51Q
36DbLakFR9Vo6aUp5GIcQSzRG/Pb5ES997gAufSJP2zLKAX/t0hJJbeaumbhQuVk1FstwaBI/woM
IR7fyG+4GlASsBI6urPbyEqoaWnPzyhUJRiPHZAUHz6LBpNiioabp/g8T4uc5feKFz+8xXY2AIl+
rcIOjc/4G1tWiOUbbVJXvuShpItJIkrViQ1PNDzIj2Y5+/D583b+/8JBGd24g6OGc64zDExx1dLD
bgjwgre2TEOzS8pbDVZ1RLajRyFoimEBMaAMjGTtLcdR/7S1iDOyo05PcpUv7wgASKShVb+HyKES
GHtdg6991kZ3Wc1w5aGQov/nb3e8JvjZ0yS1T3oexFlamS/SoqPMSof+JHSrog6WOYjD/VK+aOu4
t8WknkhJbr2uku+BQd3zWIofIwnQkN20aErxqrrpKtbUptaTYAOeVlIVAsh189urGIgI9u4GnRHg
blKU7E2PUOUQUzN2z8N+OKjpLWsuHgUEuK07DoEqpO2oMgxtvb0QtPLWT5cG3rF0mFllyt6nDfLm
jqF2eTae4bfeoEw8E3l02rymTaR+mo9KlNKzSL2WuQREj1Qlphxk3q148g0o8slN3IzM/kE14NOK
42cTiE5a3O+xlfHgkQ0JghksUHuSKnnb494f0FeK2bioc/CUgTeCdkgLuB4bU+qIWWho3ZlKR5Gp
G7n8Kb4++BmOz8+9cW6UJXtJux6AvcPLp/NxHtToERxO5NHCcTu7kfwcfg4Y5BhbvklbQdRxGJYE
sRUZ9HnOKbKdVndNZhU0MxtLHK7zT37BQgbYTS4ATRxmOhdSBv0cIXo6Wm7PlmcLIWqI0KUoNiPS
wP1pKqK8edHEWaKsNiZEJC4749DyrlpRHFtAeEnxMEjvNFgtQwIsNQLwKqum6gLMgQAqkaxCVyaF
Z/B6m1JnXsN9FRmZEaZ4hKvQ14ayknJ+YzgP94EVpvqwqRtRMK7x0g1XypEPjiy4hSNiZ0sIEvjI
M1uXMvY8ZwNT7XJyGBDBbGt6BmxzNSWUUQJTcfu9VmHInUCcAAWe26jm6Y6sLuTqZMLFAQaGyZdb
Z8Y4cvEUkdeMC15S7QhYbWwp6jLheqBY9BD3dHMdoZDY1o3JIeMkl0qU1xkha4tgg08/8Wx/pCTj
GJhvbOprlQ2jY4H7oh74sV2Gju2Z7hQGdEQEplP4F1eDmzwlr78detxQ3xANlAEWFCCRCyAihSUX
AhcmNL0AnrxoWn4JAuawAamWRBntSLMVdiNbQUFviZeCOqIFvW1XiiLYlf3tHLTWZtjPBdBUu4p9
5Lfg8JH6ytJbzeP/QFfpcnLDfZPLjiwficzkhKkZ67QPsi6rMc5wlZmty9JeBaG6Rhof7V+/eU//
UHitH9eh9uwcFodELbIn19qvmYIT53YtFy+EA3LvH9hiHKFRp3efgD8hZ4ysAj/k/90Yi4Ybm4O0
Ge4bMgf3YJGIqTR/9w92JPYVWdOT5ZkZop94+LHgzm0AwGI7in1KU6vshHDCVUirmaMfmQ6oogKT
Kif+xPIpZi3LIFxb2kGu5rUJC8bTT2H3ZuDFBx687gl6Jkfa+sCIlFAXntioE22b+RdePGvtTPVu
H71GvHOYBHGPZH+FUUb3X1iPXW2Kqi221C6SFinZwrG0Nns239nLs3sjcCfgl90wJGLhasS2i6Y/
vsialRQjPCfT3nTOhOWPQiY4Q3SgUO6jdtKeK6MoreFB5TS5VivRRxsmwUU2moQp7T1323yCAxYv
627l3/xgv/FOTkXlLI1k1j5nCAEqXDE3NjM3CqABZyFOFZxJWhMBLVXKciWxuxs9N9JxwPzwKQEt
AFxbh3/klfKrzf3ng14YH00CWE9mSEGf/9JoiiXJb0YdY3osZGC8v2qzyOJdudcpoTF2MT1jH1OB
AJZLQkpboL1McVuRSFfMvrg9BeNvS3GIUPWNEFPNmP4nArX8dC1EMVwakRgOjeeWxFWebFcBgH/6
aJfyPtoHAEkD6XcQnbpVsEeWtODgz3WGjvo+uw8fzGO4nyW535bvr138U3DoP3cnDs+lDUjPV81Q
cLRsSfFK4lMNntj/+KWkdpW2ebtRQzAhoKKg5JwMdKf8IldhTWMhl0mGUGPdUNvoggbPH2rAKYFS
0VzEZfEo4+ck1PSyU/VYbfoGr+XXsU6xM5fBO3EVg8xZm4X4K795dogUA8EymRV74Iljc5fQ3nmf
YjyIlUpbXoN5CjHD+RuHs1dCVm2qhijbWw7vQ6c55jYoL0ZZmEfVqxqu41+6Rzvdno3FpZ4sYYOL
iIxPK15tLk8sHZpQgZAEXsiulF+WnOwHD4TbN6gyBHymqCSEMEwXtivLgt9CpJeAJ2ES5Jk8nX6m
g2JurH6Ct8tZxqXZE3UCzcYiXvzwqFDDOT6kMkMW/7ogt8uPQ8CEmc/NZwyuVXZ8Mk3ywkDrrGZ2
yKbWp/wc7wykeqVlC2Y33XCC2jVX0cAj3mAF4INNqaW0n2VDOUJz5GPBzkvTTOX/4u4onxDe0khA
Ceald0jTilP/jMDHNmpBazkybRq7D89zblmrWWpKOkzzr10QAEKzc1ZZt7EBITZa990UOAKFrC44
DaHAUSc0VIFoJgrwJ6I6Te3aNHmh/p9/0T2MQA/LIpbvHO1iNP0uCccWSzWqLxDMQmm7i0Z/5Tui
AO1TBh+L17cIyg0vguEYuS182AiJ53wc7ArR0NexD00USVbi+CmGFVBHbe5vLJepVAJ/r4qT03tV
qqgfV3+NUVAlmDUuNmFOPuvcozd8cJVDRA0a3lgUdju0MQ2/XDckEx5aRiVzNYZb/dmnX5n3DInw
SG1AlIm6QOgoLbXTFp5l94OyRvcLxRNxOiW30E34MBDt5VbzxwLNEoRaFgaRivM4nLo0AjJ403iG
4+yxvHHh6syGPJsqTTNT8wjEIaeHeCYSdHQs8r+Qd4NJBvys/Y+ZH8vquBdGIsm9KoB5iwROOlB4
+WDN1YxXAG9lgsg8TdOp4pKduKsaQnOkQtxXnK0OpCZn7uLhB5ds2ebB+iKF6C1QLdALhUEg6TYo
M70pxQhxYCuh/GXw/L6AFZYEGKJMlPMhCXjJhp8OGRq5tYRY/qmjRXHVRpFHExBmXPeEXmOxyqgB
AdQuRVD+hS/hQCxFTo8/oXrD82klGn+w/bsV7dOB1j2jCUS3RtS5aJL8VbZhEk+IQfK8IRxHI/Gm
LVm+hOYftFetLsrtFhG6s86wRDCswR472k5kCZiTbC+Z9iH+yyXYS5VjuLZmoJBl1e87slglGaaL
654LhUdkT/DI0agNJfu/e0cIj6KnMMqX9cH2zPahQJymRK+UqSR2On7M5F3BuBVPf/9k5H09SyoU
Qb2OOIg2A6UrE/XI1nOXu1iBYJ6tovcZFdDJKd+NA/Lo5dWzMmm/YkRNRhtbDy1VGceTG6jtBPBQ
iZY2GB/HVyaJezaI2WDI2rD2Yl6LUwd+un10ElfIr65uqWQSZYOYpXKn0scZBuh2NBPsdnNx3SHq
HGNpoULBCWqjirRM81yMFDKUj1yUiofWICJaxvP4+l1fqkYxsRP+ybaBI4iZtB6HxZ3IdsBESzhK
BreThVxhDSsP5eBpOWU483PoazovfieSr0WH4gzlJ/GY5bf7KaW6sBuSjUGJhzGEKX25Wglu72VS
eZcQDEXTqw91cmXt6IHn8hSR8apnFsR1FwiHsOG2BjL7h4opQXEO4QtHTT5AyEhe8nSrtoAsudjv
gXdCtfhf37WTiGQF/HQTeTyEoefRTnxz2ebniHpEbKGXjKbBBlTB17v0Bh+akSS84BlAORxrYL3Y
dDERvyYYvxJPBDJnIWxGvrEE/KQ4kRrtYgHtvaeC9NotZLngB1laB+9GgcmZ5KbaA7BkX089eP2h
DlgkUIdc8ioL+XPy3yRDOC9wjoUz4YkIVAXrMibE6Y8r/S/R/8DjBd8Gw6HP5Ly3WKse9jDOv2Dn
0GTvxuXgk872PB+7aCUiM7cVDt151mUuiKcWOkK+i6q/jnnkxlsalFPSNCAuN8jqJxgIxhd2d5Ae
N2HDnLCgfcEoXV/GCCipLkC69RCjcKxllr5WzsCrOq+OatQ3Tba0XKHmxtSGUx2JQyv6mmUbFVbv
iS1CmOLTTZM12Vd2b9w6O/lezKeNO0L6lxrL5QGW+HUy6zykvCnTgfLmYKRCZ62sADMd9DsRpR8A
hISI7E58b8GP8Xa4GxccAuZlw1h6d4tFKctQXbCou2jaFGRXBewbVTXi1k0ZngYVV/6SqU+JaAUT
hkTudYswPKWg2vLHGIwDEdhGOxPFk/MnI+rJ8kefhdShD9E9lEKfpCIYJaEHMxjtlr1qmuaqf5cU
KuzzX6DTYFfY8VUICA2ohwPkoddJ4hG3PdMavwd5L7O6xMtG25E0LAyUx/Cd2/JhMYXqkkBT3Iuq
AJiqqSxCBVShUHxk101YKiZBmNzlN6pU2DKxGHDLUBSV/S2uI57EtQG3H6fRL1HWr85m4qXzX83E
YSZQ50Z0yShPxJ6b3RyYYOp67EySbpcMBUWuLNrBnYsHm/eHjni5rW/ud9fuhLz9diGRGiILOtcJ
kRVhzc2/2jyg1qS5MnxGh4ECEYzM1RmSM4ZESecjnF7ak7F3XwzouiZav1JfkcLbwZZkRDS5cZdr
ZFuqMsw1pK7Hlv4kWIBr+nVqB3fhWHwWDuACN5N6MKTGFbkYHekAUdeXl/JfQTJh+Z+GzexQwQ1u
fg3s7KVCxNFh+ClrGDRgRfFHfzJkcrWSIHSWNOVl/IhPNgbqh7ekWECkAMTvX9kK3VubBHhUZQsG
YIOTjQtZC8UmlBHWWS9+nG25hI/EVW1SHCYlOl8Mv5KOpYRIxQaIU7dur5l6BJigdFrkd1ORWM+8
XrJAwwJVhAWyZ6zdOG2yFfH6zwEAMhrhy8LmRMdVKycvfKHakCtlNZOkzpHQJToWxS3v7r2BFpLG
oiV538q8kPijhbFzQi7JnBVSYlBh/C5iUfQBYdGVcThFBNCvIvpVcWjlYzm+mNNJEOKgJInfwpuo
l3Hebz7POHnyhmkFM5Vo1mIp/SbvbSQTfJN25YrlLFPBgVF8/sk3AQFMyFXYEkdOdnCWGkBEXJ/U
xk+nuqhuq/4TtVbcM+c1kr9xUGouemZD/rawB9JE7yMBoDTZgnJrB5vc3E9IPzj9WCg66vqxlJMI
LbFp0Ptk84ObL+Mnz2yLdDAUUh+ihyV35RwuYenRO/1gB6IZANUMVGxyDItVTgV4UxnY9zOSyBqL
uIy1Kz0riSmPusN6V7H127FYMzp8s9sKJPgMeXWP4I7U0eZHqZ+qFUvZbOY522lZ0jFQWNnfz7g8
TSXaIPt8snAwhjpE70DEduIUqsNrrFmuKV9YN0kkeQEgVWBxZ2fwRn9EDqSlTMVZ/UnQqXIPmBqq
1Z2CaIgCfQ1EenZlqh3/RCENrLlQk6d+3T7j5N4Mw/GvTbqYzYgYqPymlYd4BkuiUsOP9hQUHwDw
AOwOWJAzFXujTmHvfndZqAQi4+4lYOJCjdE+HTtiuq2f8fTdLq1VW5Xkh4Ovp1yfJbvf6mD2b64N
GLAJt2jqDjLwZrxM41YuNNI/IAV7SyOpBNfro3P1fr6VOjoVniskmpGC70DlnQKQMfRIDsZ7tAh1
8G1oSu3nFkCpT2NIOtnxo07EOE3NAJy4M2/x3HJqs6RVsRsznYbOrC7bneMtJPbz+wxf2XkVeZKl
qTa9EtsSozai1kysigzVLXrdiDfOZ695a3aKs9YWtPalHwQSEhfX0Y8kp0NsrRvgp703gkaN5dSY
usy7hmQ1WJDUiS9bAOIR9RMlgajebN9qMroQtYQ14DKz4yRsvPxAL0rJcTqztMNyn+xazW6MfUBk
+W5KyO84xwcOFRGXILnKlwFqgN99zDPRBx4aICu1yoAyBysEfUzxdsdCabuPCcXfbKBY2XiXHgKc
wteZtyBHb1JF9xaIO+/gNLkxL3wt+fZoYFJ5CZ8HGnIfvZE+4l061zw6xWPW95LTnz3wnpI9e13A
ckfSgkvjmcO43BnZiHLit+0bjhxIXP6kJN5AIhuDJr9zKaODpIoTvi2svesvDpjSaHeRC4oRmOoA
bAnXUomLbTetwDOaC2qNP49Fkb0AhlL2hq8fJUc/YNvxLRxkiriSYMa65zGFVHm7Sg4YVSj8Ss/M
kt2qOmYhm04EUMJ3bvfb8nrc2gaDvCH82R0Uv+pVuoerYniEwraAlAkruuZd+c4tHj2kaH3GMJsr
uy9sLLAT7TQPgW63djRv/KdFw3+CNZn3MQET8wtMzxyJ3H94vwAb0pmopVZdBmhKreFGZYAHQ5wa
aM13VfMCBMiAKHQVTfcWak21RxnGRHElPbMDF++DrTeqtd/Yd88h9Rz8mAUrLdlgVNt1PyWmIuNV
LhzOOeWV784c0Mr1vEJXvUx4DmIUzBXcqOzmEf5YiCaz8o40gjG7O+DZxuYMWbANcQ+R9CAYv5BZ
/7Qq4l8CTwjucZUia/UOZlfyXaKl8EDe1UuMBywjgoUmt5+OKnjBBRbMwPlpdksL7fMcvoNlDqJL
uAkaF5jcSimg23n+yLXmp+e/LX4um/Rxv1pX3lV3U2lDhz3T0Wa2/l89CI26padx2g7hQgEp+jh7
FiJRIo40DNVSjH2fmaV8ZrGJJEXya6FwZuXeR3zR0p4FQnNfeZlPSWBnvSn+Fi/6wuPMsKE7Qz/5
ehzAngAWNDp0rFL6BJd9OO97GkUDIWdawRZbqza2708+nOEy852ehYey8inf7VVdHXZ/7ir2zbHI
76ZrKxrL7eg7Ei6HT/pdOzjVFqXG60/wNq1OAEtPG/lVkS6ASbiic4T580NhtJ/uUIZA3rmYGeYf
Gb7suOS49+8gx6iMeLuBomcclE72EO20wm/ofBP5jZXzsKyAWLZPs9+cex9OVhRrCwHpD8II3Frj
Cn6nK63Vlxv7EKlUCtRk+Qg/9hphPeHSlUh0YAmcP+QhhNwpFMynANAgGz9yfbrn6C4A77j6jtcZ
znBbIhES/mNywAygsjPBWZv3ola25/MKD8S6TiSRsaeu+BRhBBXB0PaFmTEtC9dFuJKm81lZq7kX
20JzCc5crYs2RYBZU1BNz/xp6qIvYtpK/RJsE6HMk2mHyd3TnOtlB0A4mJ80IyhbvOlD/O5Tgvva
IQprWFb7/ZAJ19O+ZJbYpBlYnz4R25pQWDNocvXxlcSIO0d06t1AVr3ZxZaHbksj4Fzu8lg+uGtQ
Aw/U2cvq4tnskzGeLMCqV2c8Nr3lDPo8ylo3JSse5BdAaluYCL/oHHwi4xa9qpHxdby2kU7ZABhn
4rqMNQdmEkGWJlXXvT0AMvO/ZHibjVczpm/4b816mc6N1J54UCc6luNV6yJysCNQcxHAb+JI4gmF
TZFmJvep8TStMv+J4QbLn8Py1vvCGBlRpuNdL+kASR7+wNoByfFIynfdk9QQo07pWK5oVVxxkEJK
tAFxLZBIO3Zu1awlEGhETY7gyKdMdPrnrfKjV9Ubdc3oiWp4ND616wlDjUdiFv2HqeRB2QIPUUtd
Fu8RVF6M6hrfx11GBXAx79zratUVfFgrb6CCcfYeNxvdSxHGDNFTAC22vt7cDoAApbdx+4jr9X67
R0qioPlhuMKMMiWcj1N6br1PIiqCvVDOsvOo8867uqACTJiVPkzqjIXCVtbYpug5vSCYilq8KXTH
0dPI1XnOzGlXqxDKPdEv4pssZLxCUZMbKZQaT0PSpKcM9gGC/SDNKSoslzU4/a4bFeldZCTzAGDP
7X4TowIamKjSnxPBBtWcUfor1HjrnBRpZSuganNwSdWPQmxGho+NmAoFuj4mnSOZfLzspMdfRvXc
+bYobvNhZb+UzQUWa7ucwV8sfluowfleyTPFtQ8q9ABqSfAkd868NlstryYvuPhrcFfh4AP5SUF4
C27TTauDxdc/oVZSTC1GTnrXkl1VDdYdiAshU/Gw4pYr5OTe4DRhNVKJGTgvkHVBBGtjybC2Zgko
KfHHGYFzdeYAiBrYY1kFOSmwnqeblcPeD5VqBF1S20HRQhCvgwqcpDHFSZ7XRc1YVMj00Xn7kyfH
pt4ZOBew4G3S+j/RUiSr0qDDQ0YkIimhtdQ73HbHZBY7RvgJylx64fzQaiEX5WnG+hxxaZHUeecR
tQlSNBzrmt/UzculaVNBGD5FsanBlI2vMT/tzxr6KQde2pGkeUisZLO7vx2kjbNu64WbHEjhhsV5
N/d4lI3N4dpiExzcSq2v8ErYnuJy/U9q+3qYfKjZxnTXtd2eVyW+dqpEJJtaitQ7mrihl2PS/WCs
tawSu9hxeGbZ2ChyIFMPBXoT7VKv6OfFsLO3Vfp1vTTbWfubP78Rihqx8HDooYycq6gg3xdxo2G2
FeQaLeeQrEKMa7stZt2gfv8YNgnrs4imvXhZqScFrQbnzGeILI81m6yu08aKw8rXfVSpQTc7w1T6
BvivjwLVvIlrzAJVyFtjWjkADzaLdLuArJeOWSHilluxGpWq5a/CMtGBpy6V6QsFLoDBbSAx5Jh+
X6qIDAyq+mL3G9hMjAb49RTUaIJz+i+EL4DdurJEaL99+VZoStraaXoyr6kGx7GuVI64KPjidR5I
h1qgSwHw68WOA6rui/C0vhtmgvzfn8gZj8zkJRLcAfCV+83D2ukX6Aju5tVRhMBB/AO9Qhor54Il
hKHmBkErXaWqjD8ky5rN6iibnverb59H5s4idknSTlMGnpZy732LkQyIIJkcS6Jw0Zhq5dzXwdHH
hEDByPZlB+2YbGWFsqwOt1epHRiEHoIaYDKJRBgz74FLaRjlLcxTb4JnWwb3zr2vk1jw0TaDyi7w
X4kU/6YQkA6Ac3+DIYOIvcS8jAZVtJM84KKAXS423pvaLp7psKJ9b+sxn4L8EYDHKSh2B6wi2Eqf
CcpZ5eh3gbVChtBJ3LOEByyO+RsxPTcekVCqq3uMsA8yQdCUJQAc38TwrS0u+kSSwOjBTjIhxeM5
OUC8WhLDRUorp9kpWJiuV9nRgXRhFqdGSqiwMhYvhvkKGrxBMoyNJUBBfrnRM8XmdPYeA+j0zGwB
UmeSdM7oQEf9gtPUL/WEhHy8FpQeOPx36WbTYEfme5NfsSiFZErxfHkqeWbaLiF43bG1439ryeMg
JAvqy8auC192tDQ/czP4Mui6eatWYlp7qtTF1xGLBHRYnln2TmKd50uS6ha+SpK/njkIyeNn/Wv7
hzedn78gRnIXveymWX1vrsXxlhitbm+Lxwz8TJENg4BFYchWNbrVvc0j8XXvdQUaYZXWxOwdRWr6
PmmXkhsIHe0zcd5Zyx/aIFV5hV5yfO4gKPuXE3q5xTQwnbpfyVb40Y7R8xxqs72/PhKbfbRL1c5G
TbLSwB5ptz+84n4+rtB44jCYMWLZ9O7+haRSXxENEbDgE/dSq36LavPgz+BrQwO2VqzMn+J5VxJw
7UtRdxumJWPZvdSOXMVHz68Y0bfTVrg8oLBgYmjkEf0UkqD3njEJnvtsVZtoAsCe5b4+NLL5cx4W
1kjzX+TAGF0zBXb2pUbSlGYXzH+uClzdbKeG9Gjqzwj6FPQSfDmg3yD4FwwRiAFVuFYkZ6Bwr6bB
BBEjnf8FnY4HQL+b7NwPhgDKa3NeVFp6ofqgkltL2EVDnTAuYw1B/rYPxGvPE+tEunTZoBafFVob
oEiWcUlZDpG+WUNqclrsX4az8Qgj6SDCuIpmsMWUzVBijghIKXnqA6hMglR9yehZqHObLG4EpuJS
ArciwBjmbZeGw8oTEYIjISoFdzuV6aktggNvGDSwJlxxzRsIY39yDTtzKfNANJmozWnVEvWTjRo3
+80Nm9hHey5Dn1K5tmsXSFh+XPCB1S7gMLZBClj3iWmy7xuC9BGuXZDILweI/bh1NIhq2oDMaYBN
itQ0zc8G8HN5kGXVGNCqwrUTxRQlH+f6CeOPjYI2Tar7P2bVle4PLlzck8aXJp+ufeuVdr8vxetX
Bcfg8elf3TM6lWVhsWAV91L/XeGkqGSRbh3KxR4wuAM2WOMqUyaSgcFq2SjozWVqvZveVfxSqojx
k0W/wtiX1m8sAAtkmu7yj3C2yMIUEqIQz4fwjTOO7C55nGAHYfZrtUQsKLKYX6XDOnBDlg+t3mr/
C2wX1g7kJadOdvWvvN8ReXDOMp2lf7mTKBHiWPPNjHPWBukW2zd12wExcUh1aEDtp5Aqtf2E4iAI
RoCwh+xZuy167Vwc/l0ipWLzSGwzg7TQq/4eFGTPYOgRK1fwecNE5r/F39sD+erHSB2RJc3z2TUG
VkMuxxLYBdqBfncIUkZLF7vcVR4TjM3NwAKkYAxvqlbvSShf1Ytym6/PknZU4BQmlESNK51VzRGI
CeHBM55xX2xs1eXyUCsJO93ZmPLv5sXBzYO54RWxLyF5gsJRBfO68MIcpRw5ACchGFAEZTkR3Um1
2KIc8a//LYC4BOqqiKQhTR/DOwl2bLupkr5uZ6w/A8HW3tMrP9DZUvIp9c6vk2Hpa88FohKduhfe
YiDTZQoZeNk8Ntvgsgi5foE/UTmiKTAnwyElGmAQBXbs7Ne7akTIHsaCaPUBJXhUuujGvtsSZTlQ
Vok15dI0OUdtSjCqhjy9fDBjs2bNz6w21eJK0P/abdc5U/AjS+ia4DiGYSA+gAZt4DcUCRNHBxK6
t6sYJQKGFbXr6Ps8Kw9lvaKSgAi99iSXBQUe/Y3fVjJmkG5pqfuYE7KB8XQif5XcNoB94qJ5uW/T
91pz+E77CWtZBcU6M9tHoJCgxuek7THCOv2EwQla3dogHRoMjQb/J7FZPAvH+r2y/T4zdW+b8uxJ
wlehcR7fEVPmeE0npAfrdRmc/osR2qArMPU+saOoQi4lYioyDfHkRsgSfyoP2zdfSHaJHYnnFoeZ
IYGcGh4JeoYaMt/NI60X/upiJfle3Z1L2S6bsMmmAXeFciCBvdt+Tr0IXG0/x6kyyEazDpKlghk/
j21N1c48qYtQ4MkC0ZoeeAQKI/asvke+YkWujuv/aMi5vq+X5hH6fhuOHeyqLUAsWLLRbVtvXSnh
TP6/2VS5Xejs+Esxy5UuACKbNfWktPk8eupWciM0W5/xSsu0pPBiBVyjulgAsPy/M3Tl11M9PEqZ
fLBWLx8bz7CofSnkJS1w56ibQR9IPCVUchRwYfmtuBHvUSLun3luXvATdGi7v7xXSX5BROf8kljQ
px/sIMMjsWeJ8nwa4jgUbP997NJAlbqqTB/h9I2px74cXcMTT4JYxqMlkXAbWfmx4XERwvWtUasL
YmiOgliW17EhNnXIB6wOtMyiBwEdgjb3hHHkTGWwAPt6rXebu7wpB8IzP5IWoRKJIF90rSKdFC87
aYMpgG0NOPJeIPesOY+mAosONhz/ZQUS3VNYk37o8DaH827UAIQhKE8uTv0X8naPFjsk2KMioLeg
I66ynsF3TI/pEuOrIzHoS1ELR/Un3yv4ovJ0vaUfe3dJrWhbjHQoQRtitS0+IEoMaMSdQeEMLaD1
ZljrHbLID6zTY0EGo9COZEXa0javoxF7RRK8Un/4mbqoAIpD+Nwe6MuqYUnTdubV3Gj5H1arjYUQ
prD0V+bR2iLRjKOUQYl6D88sOflEMykB6VYseQORDV7iuShgoYn8/G73tNeWqTG2YwVQVywX3bGX
VWuoZGjdUKbvCUwK/tk0NE48pFes67ghtUZ7r/9I9bb5BImTSdteHg41OVvEMzO9DTtAfScLwtuR
0eoVdYg3K4S4B7s5nDFeb5bDlfPU233CvoPOMfpTu/8OwflUM9Z+PFE7oaoaEQgmKv8wnUw3VT3r
xjfbaq7v6nB6670C3bv5x6MmxB3p5YXv2gqt81Uob2PwRddTZ+yT5YgM7izSQDGW6mDB9TBs2tH+
UDHtVmItgXdFy9aMpuscZpv6jExS+XzE82WGXMgavULLReHo+z0QAAQmMgcPb09fmYtoAkrG971c
ognE+BoCn1rFuyJ4EqF8iibLZN+LWVJi27+Wrv8aK5q3kE06cBolyQFVISPcljiFSK+VX5mo9o0C
GSX+NsxddEiKXYxbMhV3G7aeZfzWXiGZLj0k/GS6dF2CEVdF2jUorDx81V0jaLtZx2kUbYmyxLHx
E46JvBlb2v4M4qTlV2B3iiTmO0lJeRSnx+Bge/8l2iB5vGxXyPu/yd5e3XySgOo17+yV5R/y1n3k
cfI90cHqw+mQa8EkZJ/3SxLoeMmWc0jHZqn7t7ygWP/fbhFkhE3eP1Ha0a5weDW6HbJErY+EwBHm
oDQckluIoNmT0QbhZpCMYugVsLPvDlTNYACwwRWiQcqsY2y/EBJqvhrpf8FXRHb/3ceI8POd9XTD
whAcFvzFNUABG0ejdeMZx3MK2VAgHJCP3FbdG50CPCmHzbXxf9pjoi/FQGGzUy7PuAICz/EVcXyb
vrVEutz7XzZmFgiBkSvuYp4wtbOakES/oxPuhA4UV4oTrOtwdVGGHeCLy08EXVpkxJRV6fhnAt2V
yW+EiK64KV+iDkckaW/ILZFvQWw1VdduDh0hjSmmZChl88ME9KH/WjQEtMXGMIsL7BMQ74lJjtI1
D2MgAV7K7UPX8pzg0KHcuyqJPKcohVm9LeycvAO07k3TDedXzmUHGOAct3k7SfEdd2KY3QgEgtZY
u4i2SF54f41fKjYU59gy/Ld8Tr7RWv99lG77gWAeexvuH7FFsLg7KB55s8EVJZF/UCCcYlR48en2
KvZEPX06V5356EnKeWYbyX2BhOG5F9Gugv+KnHLD4e2beJw1r1Jby2eZbqR7l9CB51Vr5WENwMYi
/1M8Vgo5QJVCInezsiIyDRYkoBX1dH0qyBlMFfvBLnY7+x/BfICnFij0f0S6CExJH3DMC4d17oGJ
1HcQ2DdvTBhQIpJJs9VmTUX3dk45dPkZyPf+qjhKIq1e/jKV/+kPT59VczCp8dvu+3Uw/CiQptxX
Fc/IeXZ5TJL4QmtmIqx5Vfwv99dkJ6sP1jts7yRcUQuxVzkbXuuuFhwPXhi70tKvDHgFmafWv/So
hCKDHvz6hELsaeXHwAB9GFGqT+9C5aqXAFJMPT5vm7+Tz+K4IqB95rAjLwW+OXmZY4pWsnskocGL
C4UM69A1ICTHI3lFNAwjH1FinPkYw8te0FpPwA9lH11/VDBY7+jKA+g3rBtRIzchJGU42va3ycrr
euXDfmj3UmxeIYDlnPsdBLR/9lt4pn1SyLR2PRVJlNTlsHNd0Fs4IEXNhSZaugEWIkPel8WJbmtO
bVSQyD+VYtlX5ghbD/13zDqwTCCvkHQVPBxHKp4KsO0ZFxoGu8M+5FKBm7HoFvf+NQv4t9pblzSr
wmGRWJdmkQtiHLpu1afa2wuIwIajfbw0mIYow4rm0kDTmzG0euQYdvV0MWoS7iLpb1A+uSWiEmGQ
FavwkNlBpnVUA1xuryI31shXg0OV5yewD42LtzwBhX71arrA+p0VKKyFQosN9u8xcYV4bpyOYaSE
jHTswNmyy7kiBtIWYkup82t32QmptDWUYzW584pC46sBuPx6WLXiph4DEuakBVBzoWlG35KVqMod
tfgFZdkQl25DNfiK2dVkfrarAEkKOC8L2hEvtUN8qmSXQAt4cVzHLqtkX5IR3mTp5yFyVDl6YpIz
H5OKI8M8+Kk7zu/widpD3xrSLuGh/i4dGlWEy622/tZ+x1gTKktAfe7qGh4rqNjHK4zqCIEmiROD
7n8aKNlqALzxjC0lf7KymAVSLxJw2l9L0aFyAMcTx9O1U5gEUWqRB9i3xM5hX4vvQeY3Q7+gXUGR
lulHidpDOIz7yeSrYMrnHzZrHiCbctT2UrJiZmtsy/3Ds7tkZgaQ69Z2gfbtz2cEvL+b9tKddnWO
I52KP/h8L8NpMd5YX+v+5mkCZsgW3w+73iskKKVookw1Pk7pBEWKKiA6mf5Zg99W4h6Igc+jiruI
MJ+a14Zcdw28wVeSQOFlq96HX17ocpDL+r6Ii01lO0CUKeR15WcgwiNq8JbDHUQhwi1MnEmPYtob
Kq3/pE1jLJfF+7btwJDvyqcTfJ6GCmJbN+afsugi2LhBOKRaoOi5IFFN1tmBK7FCQ3fyrnyCllwj
DwQ1ukYNElXcmtZHAjP94Y1HzuhKDmrGleiLlxFxlIdUX63jSi24AR5OkkoxWo1sbK4BeXY4SnAy
QWRA1SFLV8Cbc9WX0jclwHiJPJT7MtY3KtmGnMAVXDCvpoYcYyZKlfXwNWo53cC9ZxwSrsHaRaOm
+JVCjrMG9uZsnNcBpjXkbjSP7UepkEu48Ht8obwT846ifUJPGicxeVgO6njiqb4Mk0pyjFj+Dcw8
lW0MHHQ0Ll1WBn806JCY/wXoSBE5fCnC+es3rDIVh/GlSvlSOHvbNXBcP5uKf8PtmdG2GMK1+jG0
W5VjIednB9ixlfLXeJCAqWfqAQrhSMBZl7DPKQScfiEqQiosJAyOMJSYO3D9dopHkeynm6LP2Gj5
QsBSULA84zP13gNjrfXPXlVHKBhhwd+iKASjcmH7zd3JPIFqR3CxWMrICOjFW9mA1gZKeOer90jg
2X7ds1oCXJOKvA9N5Sb3dLrfcsZCQYZPqd4VBM8oM1UoFE3J+yPkAJCApkfkwaLWg0tWoC1zNS1k
Fg3TyRmK1baQdBhm2KDYIYl8K2rP3+u9ymGsNYITDkWPokNagKjnLVE9mgywoqX8vihpyLx4HIXJ
uvDZWYLOB7j/N+SI+CydOnsXraUAyaznKOnUZdz7S80xYbAE+Y0Ve5YxS9tKooA+540jvRbAqHDC
6ZCMOWZF27nK3zUFmIJP+SZvQoTv00ka7p9A5C8bOXy5lcNiC0jsyE9twrH2rW8jFFRBwjFdkuVR
Mf/O3czQd6PkmwxqABJx6+ho6kf8fQ0GpEYJrEvhqDDmQynxgS9PfYhWOzDB5KMh+4uh5lsFOs/Z
/Or32M2ilY6pyHuxBRR4XYx7dHD3BXjkjEe/w5e+asASqwDmh3GmfS6WFocFE/uxo5JZoT3k6Ojv
lq/05LUaxSvIJXCTYlVi7Rp4wPNeoUE7pBtbc/0isV5kiWi0rO6pE2ganUbBRIYoaCaqCu2UrayE
hQ2nOZ3dAG45leQmn5V2vuYUvakoKgBmv1kbVcSDRoQkRHyw5onWvDDieMDpDi+lcPPEXl3fjd9V
6hnCjCunzeaCreKDoavc1q4ag9UcReKA/EFMEk6Ug95vvxqFsVtiFCzg21gRVRbocL9IlUz6ndsP
Yw//JKAzoXY/KTOfzV13+nb5KsMH70AnI2VOx/vdnal6yRC4Il43c2QSbbEylc+ckA2L9Qwn2SG4
nDdawzOPNHkRnIGOnXFCIFoEfZKBKDH+GEyOcrwOXHTOuVoW1u40RgMOKsqEtgAjlyJoSB5hAWNd
Zd6cuDYL3knbeagLY8GbrJRMgeHy2iom+62eTQhKRZXQ6f5NlTZ6OpvYyf7o1Qr/ZakrL7gDSXAs
pxPrsSg3ScwHVGbYiugeq4G06ZZTKXhwWyGmOLQMYs1YTWsINrHoKW+aciyWPgBiLJ5QAlouAd3f
gGZmEh66MvTYlVdD00oiPIkuv2WcktgbO4LNIN1NyxxqS3rYQZsLW+tC3/fkKX5hX7vjjVALF0Zw
rBx8oar9FUbTNoVga6FWQjXfPkLs4FbErn8gXAkLzOb3P9o8dXDJtAnr0xwIUxeQoeqOGn0bhYQF
svsv7i724RE0e501U/12j9D0LjvujAWaW0NMfEbLi1otRjKnoudOVh5RmT6gubDDF/sMpnHIU/2I
fxlmKcZnOrDPZ+kOJ/QmoBKc7tRNjA0PaMWa5tEQQWWFf5Vn+UKlHUaoXITsSE6Mot3la7cZDgCo
ZzIKyxRozQ6TrLVM3a8Jo4NU3ZpuaqaaQSrw3P8X3U8O7bYMtsTEprRBt4ONOoY+fc4XDyRNX/wJ
dqkTrPJjE9dYYc49/094XIisyuDQdR+q0RkhC5dvOOHI5DrxNMXM9MzhuuoRfh6Ko98cEIlopSg1
PXXdoByXvH7aeJFtig9GufCm719Ppey1PIBZvuXg6hM/MZNTehH51D/vog4rg1oOh/aeNrtdfkVq
hOVmcwM4/+k3M9aviWfCR5Gk84gOyn2tL3CBR0uGaURM0Xpf79/I8vL+Y2ExtI858QtS6Zqbmhrg
w6eLxuD1l/t+xQfkeY6VvPipqmoUdvhqpCl9p2redKYcLOg/d/izMxg7v+Sv2iP29A8d3Mx76r40
JdBRNha2eXnt2lAJy7aj0RiZFGrpXfYBt7mU8AtMv+Tg17uaGC4VuxAmZSEwqrOpBVCl0J4HTSV8
6lPLc6jJFUqk2t7sxekROHopoZAmC8HNJclvJN34/p561l+9KtNryW/6SH1kyCfVx3ifg1qFkI6R
Jw8FKvShHaPGmR3vYy/MEXBzfdUQitSbzpY3MI3DHDWImw1z5e2np79KQmzLaF/w9Z8ksfRRcPqE
DwpMGlO5L3F3vzo4xDSGFodxwF70KvSG8TXuzfhd3KKc0FvD/TPDXghcShoH+0954gIHTRz0SjYL
sMvazx86fmaGzOAYZ6jiPukNmx39XTWHThEQ9RfN0TqPYMRxAjuK4Fl4lebbDgLFtywLXqU0VvFH
LAz6V4wUBBGhAaI5D5SZBDPZtmRsV30eCi84G7CUu8MRXTN3mAzEY4ET9fZjQi8mzleCDBQ9S5n6
R7jSzj92bs9OAu8TGVDwQrruoF8JvMQpTnUcQQJrIm5S4h+OAB9+bZh3oMbC9H6xRKeVSXC7RKk7
e1Omfgeg0l+kuP7svfcF8FSfZKCJ2cxW/ri284QRIXZYlzkql9Rhl1ypUoWbisErUqlhtQPcU2kw
NrpdMhc1tRmGDoKQvnE2RabtE157ykCEXO7DjcC8QrE9qOxICq8JsC4l73//rD5itmU9qm+CRWv6
LxeGB6OU2ZyF+THS1b9fcFBCAarz/Zxo4LAvgHDaY+IeJyI2B8ner9y2dFPCKLVXP1+cHiD59vxW
g2F5K9XybamZY/h4K8Z6dpEGQ1jhPiHLEezSdcpz1LKGCF1mzlTXFTSz5XhSAx6nTTx/gTxl1b1h
V7PHxnCjJob/r3CRI+/kHrDGUYEMkqGkYl16il1hDpnw6wFnR38xQACbgrr+UBNNnjgTyPgIzX56
otBXJrCmA9UzpJjD2owewoZGBvd7qsxzz/01xoTa+Z8iwjBJ3cdCFD7jnS7GhDmdlwpRvyLL65Od
gwHI0IJjHj4SdOvukb7Bfpl5X7jX+yYIpLsIedMj05sEKoXZ0GwToZg3onLRddnyfgh5VPlPl9v9
+4pgJ8fTTPLfjZ8KNKSXZJezC5wuSDrI31cC70UApltklJlc+VHcXX8VSXtOigk7nuZLyWGrHn3R
6fxbtjyimxlwuMPQp92xMgZfA5Tk9/An8nN8InoM0kRtNfR4eI7HV3ngxYbGCTiD3azV9FlpvkSL
v4aDBF8ITbcwS2m0q81xqeHi3lfJ25GeVeFqrgKPwxCd4h6LGPIUXKnyRsuyluKySl+Euu2ZAOEN
Zdjri+XUekcnghQsdJ2S+hzLk1DxtX9hSruVoK4nnsrhIRhHNJgfqE315WZZKlB4Gs2nHiivDrtA
11hk2zhlsvnM0nrhT8EUZXSgG2K0VQatqmR9OS7rYX6ott/xJdhb++v5uWT5C7BJAoDIctX/Jfxj
OceBO+uBTYBj0PD5Mq/h14gIAMwe5WzoavyYyOBBElAZM3Nt/WaI/KwLYDjVwUfBM6o7+ujQR+iX
QFNLAVhI2B/pUs6Cm8JGTWiuF3/PAydqHxYFGJUqZRJZ/EI/pF/eSzPpaOGFdP7JTINz3p7a7JqL
SKH2JtiHS2Tclp9eS4YarQAW/QiyrLL/ceVYteNYTZTP9dFT7lvpow0+3BXpPcd5WboqgJpAZYVs
2qn0RuaAfoy+xOOLF3rUfZ6L9AZ/quWC7G9mrWf2UU+m7SBd/Vzh9Rjwo1JXcyKYdUXUW0qX28IF
O9SWEkZqAkcyZrBtCwUein3NBuAbnxeX3St1BQw/sNcOQsFDo3cyHKR0AR1aZ0DT3Qr1yihImq3+
Wg4+0WkvBoMO5cmgJEC8OhgExnJibbnYiEbkFmcA9HITpZnXpGHznHIK6SDkimxymCkM9NxAMYoy
vbHAz47zpDezUdiwlsM5LKifp5je/Uz8Jw2miOp7Hf69TjlRWZ1A0iSxmFMl+B7Y9Wq91cx+pU/H
Pq/cAfhHpbkU79Ibab/Cz2IlGYZwjnq1QwDhyO9++c90n3VSESxR979EbJM2SwHS82mNUvZKLmkr
++hBilYFamTZUDJVIn8kCdQq7+pISIirtQMxlvuHHNB3GQtoE/hXK1uRjtrghwLd4jb2DGBRMPmX
8iHb+4t//bp085ftsrE9pjMncz8/RFnyfU6vY8er8dTCwcQUniPMO8qEwZYWu733UaissDjGKy9B
minxlKi6bYZvQGwEjnJ5XIqz0Ydc8nhbDz7q1p8cUBVMPwoIGtseNHUtdzRrZZF0RyA1tXEpiluI
cNAw22KxaPDsMI7MaCaKqtKKzenX70+QXI8X+6JQw3/O505sSyHWEJoWmog82AUhRMC+ckmsC4Im
VysG6dxJpA6MujuB6j7tG+dyaP5K5dcv0bTLOvZXSeh34sG++hOkoXuQRyX1IM2Te0KZrG25o9wr
oaT3t36TzteMqMlTiBEx1QIjvLRszDUVWoudw0mm6JqeL6TqesXbylVyi8B6nkcNTjxeKPyOSoY8
2O89/XtNYLV5sqnhhj8/KpHNEpUwoptZBIkBUzrgAGVgRQ1d8o1r1devqVzeoCIA8LerK0HfCbyA
f592Z58258mlAWntyk07BQIYcr1O6CkTiEuWER60Q0b5SpMOwLZ33Pm6perc8GX9hA74B+pF7ZdQ
IxrLRHlDLl0EkfukL90CcKVZR6N+fIG9AifGfyHdcLo41hJmfpnep7JHfHz16+EWoR/nVGVPHjdl
m6HI5wcHZDGANosBsLpMHl6nvafdtxynSH3EesMo6UZddoAye15iAO2nKeP4jeW/BCI7zZx1Y4IH
9nzdSw5jFDbH6y1moEYYh7RKSzxWufiUnZ4QJceLExTtqg4vNe7Zvz9WAHC63+BwkRCGfkUO/wuu
jclOBBFnScK4tx2PhWwXMZhICwMrNaXM4sYESMkeV/HlvyC0fioUTD0PDAVUgCY9zErGha9eHLNl
YClSse6844X14GToKZoxTp5S/SRjzHIJJW6H4gvzIGq8sVFNvEUfXOu1YZbopHnuNUeAdZdiTXJi
oMjB4/F3IoqTH/xhbJe0I/rbC6mw51/uCvw7k3UnW7IdJ/BHNH/zR9e637MF70fjW8PpuJO0BNge
r/KvrWIx4/pX8GW5ETnFbHmF/pCXtcrGC/yhQoAJdxmA19iRG60J4SYiOAPCB1zOSjPEzeRl54mk
hmWYzjBc5F13rh9j5bU4Gm4R+QeNET8VnJ2xE9KpQEVqXGVPbS6hUi4ypD2StginTpH6D1nSQiNj
+KRdyy7Y7frmXaL42lQNmG72xI0wsE5QYO1lzEvFJqcR4AsOGRMKd55Fb4Ngo8wGJl+0qDk/buZJ
DLJwGh5mU7GJZopEIONf48T5XjPlrCieBUruEBh0hjRSLn8wa22/e8R8H8MqI8e5N/UdqPH6+Nez
YNFW8rwq+Sfxf22ayUCi5XMuuJadzP8LtJtinqygrsvIhAUdhSxIVOmFg0AzzgAuJId7kSdIxWP/
JqQm2n0y/sSAB2/SWYiVRjPn2u6jcgCrGmSemJkmdXcXg4gNwPH/9cgKchgWVqexR9dIzNKKHq10
x0GOx64qstGmc7IbmNvZqZDBAPl6atFW6X500/UMDSdVzQhy12ttiS6O+1ihMDQiBmHoPKZRMaGd
UmIUGA5Mg1UqFwzpDNbLnHqzOq1sHq39VDcjEbyw2mhwfwlYTbX5x9GBvVfpXNK6tdzEcSxUNOLy
GktQdpZWNKopAFFF0t8BOCdPoYpCYIwRrM9KJdwEy1/M0UmVw1B5cRwmnthD6ATUvVNbdnB9By+D
9eoonAnJ//neuiK3VT+VASLt2pkd7zhiIdW3GwjLFs03tNUKI/6i3yD4zSFXiXkKAW04Nga5rlJ4
W8MO4MUDh/q6PzmGEMGhSdO9QOznDQAcVQNVuVgLJ9y1GDY2SdixcVUFqZw9lkV5S5wN4yn7JVs6
LN63haHyaz/fgUnHoWn5TVs0kubAvQDvAFGbA7hSpConlGyMTmJYRPyk3AVdDhSH11VXuJ4JxPZj
nlVpqTUg3lmmJrl/TsMCvF+Y5lqTJ0/iZnZNGCs7Ncittxo9C3Qg7hjb+HS0r/eILvig+U5VzOqr
m+jZPBwBVsvRBx0AM/a5w+/wXJ5mxJ8v6FruGpskgJ1HXf2LRVQCMIhHGJXAKDQGs4e4atZTnibl
ONT40N+Q50XYNjwulzQOSjzLZBdJvzsj3MHBNnqCH1Lpu744W3M1AUqJTWy9C9x+WbgwSbXoMJYz
A6XQkqb1Yr8SFx1gOrCK/ft/4UDnAIDi3SbUzgUT8z0M00xlQ8xZi3OeH1EGiHAjFsBOPohSJIIg
kZ+pZZPLqALqsXzWBgI2ZormaEUi9XguDyTXu2rC2Cyi7ApEat9g6I42tUGqKe69Duk2eeBCAhPS
IPAAxXCjxn8V2yklMvKtwTqw3qAjZjgIcyEEXbJ5jbTcdOHQKXYbp8/TRArL9+vsiVk71Bd0GqOJ
qXZEZg/ckpp4u6/H210k7c/Wy5UWvpk/3XgFjjpQORJVze6zYQvVuVSMUzuLOZCyKERewxzqBUz4
LGC7wBUH7WIUMolxlP0EcHhH1VMDrjpC6FT+WiEuPmsg+3J6avQ8VZ/s2kdDvMO7gebUoOUrztBa
fZYE9tW+HH5TzLOQUZ4BL5HR28SQBm7VbbdhfdepUdsqO9m1RXEnsVED5wwP+Zt5LIUTaqcn7e4j
7iytSXglNeUJywRS25gdaedH2ZNkDFrgrCIg/wkoSnVjAyW8GNo+sIPlyNAQzc15CdzqO+Zu+Tnw
2RpeysBLqy4CKijWyjQMCrGGqW+V9h4k5nr5pUmbKNB2x6P/URjMvjugDyW93VyLD51nMlpsfU25
bXsOjBa6VrExPu6RzEqtozDyGJnt/nnTOcvCOEeVT8TgpbY6o2+Hnhl/j3gVGzqgtfhRmu7M/Q6T
m3Z7ZB/vz1OK3Dfi/GU90FN+byLB0r422xY58Nn5ohun8l/hs4VN9ES4SUqrcSwXqhWfpMM9dZcV
FqhVeAcwopDrpU1tODIAbZNzUcLY87CfGbGTILlKrYom00iE1UUwYJJN7/SPAn+vNobG8AI+0Bji
iCyOv1+zEuEXuJlveoMmlmRtEtQ3y3MVL90cTEO8fZpyXTMtL8pxqTCanjZ1BiP5Kt5bIWIB1ODz
j7w4pxHzgRucq8nnaI3LcbEJAaAb0eYzS919PwU8Xw+0wmCidxtOeHnMyq8FQYVadTAPzVFpr8uF
wqEWv6vvfB7AtGW2Cs9g4FrWZLknWBcjpEVOpPhS3b+oYu/0XRU0Rnry+Q6qymAnE9urMald5PWB
zH19B/PDIWvIA3YPrxJlGCDD1TZABi/gu7B5QfZp/1irWM4oxaLwOaxWG2f8b5mCKT+ZZVICslGR
YiLRrnId5YYDLZE8EhYOQSsEtCINWnXcqCAg2t13a+nfYM5MoLrLLSkrHJd31laHdX9QS+cvtrLG
0AsUjEK4S5Lyv31PKfIj4MMQeAUM2LQPS74szByYygr4hebOsZPkAhvqgh+zTVMOBke/tXSBNbuQ
XNHgucqqyEYxxDbm1XVuxhUKxx0NvI2LkW4z1mx/yAGlLHLdFIAQKcOeNiM7kG26vtTgI/cLLBXS
axU/mfjVCjYuyODSp7Z/ZEmqwlJ2a1yv9vxwmj3Hbvx6M3SKOLHS5t3jh/UvYuSQ2Ackk1f6Ldgi
J8buqOJdRieku3qGjwto8bMy6k+ftNGmOx/Y8FXhNbDcTS6wpUkIS1DLK5UTkat3stoSFHycyOLr
rR4Rs1iOhGnnfSlnw1+1f2eCI/aSpKe49t17muM7GrN/oR2asr0PN99cQqzwKhXEXlVrfufcpgdl
6f+b6xuHW5HGe8YXG8hYEutnYhQd9/P3AfTYZc5TgS9HoF6z9EXtS17J48mFt1WzfZt6AwEuhyqr
2JRTkIXRjJeTXndkTMnLvzMEXWjoHNK9cWbDtCYQHkM4fmmPLiP/AlllJZHI0nfZMhDJ7ZOK+FXh
gXm6xuypfoS5tInitriY7bKLl8zUuWiMf4DSHrmY3c83+R8meuwuwnujjmcStrPNbr5wE3B/aaAU
+vYtqTdqfv7UA79YY7iHXi6cUkB1hZTQqvRuH+UJcErk+dSR8sz37hkWeE1hPtZWhu6EJiFpSs4l
VaIvJWjSpJ9egAoJYArRTZGt5ke/P9btp+N1mz/PwZzsrKoDVrhVkA4S7Hu+DVqWIWOrifkNWfF8
bRWiW22iPUznjWmNAjKSxoJgPTPqA5bUbuq6BBLaYdNK9oLqiXHTXcrPdPRm60YLGGgx6TPsu0fQ
pspoXe5qzSuuwpKoUA8QSmFlmzjzLE84xSolRk8E4k6yVu1DkuvE6F3Ucl+DMLeXKxS7Wc3U/2xe
wxw0ebcho5qX3JUnlQfxxSilpQixQ+b7qRruz4uLjIor6pr9dFvEJmbRebdeEh06u+7CPAfdzxx3
HSIwEe8yNQ4z7BhkiFEB8nMw9rbvkH0W51AG9wIdPeAr0CUN0IwMIMI2KuvllQdkFsf8pDrzIdHE
o28hgLwBU6GmGxmHYQ4/AiZwTvJqnRb3XVAgz+DkGElJDLxkJQ6Z+rOiF4f/HHC0QVsxExTLvFce
FKoiI28jMwdgMsY//NQ6gqZWgeg1JFxblB25hulrECWbc/tj69YHjdZMWtDVQ/IKbKhiM9UuuNPq
D5opNBRDoRDt50jC5qAqsJL3QbYDG2Nz0snC2I1wj44EFL/s4s0oRHZ5OKTf6/3KMk9CGLrAIzHa
H/eQUKWTOMjVxYSHgqJvGLksptQXABWPjV5K5D5Imvsz6k+rX6VqhG4U5wAI8QTBGYtir9KR74G/
/HsL2Dnf1349BqzfeQEsdko3hwoYqHSGCDYGiIH5FfJ1+kRKujx4goGR5Ayjv2gaT7UvKb8WQvmL
kJhnIrZi2s3dSgAd94+usO91siKoSQqP4ZFaGvu209tD78ukLR48qiDflYmxXZn2vUo33G0bm3H6
+g+apqhwDncHwyvGxM0nYBujGxYUxrGlwUgU8NU86+EiJIwOOrxwu86e88seFIWyz/IqfzIDDyf+
XcrWflpDVKVtawZqCudHI5T2xLwgTSQolKqUwKR8v/bgMv6QeOcVDaduT0VAj/n0C+EtY27V+4TN
eoTnfl4S5gHTGd4s5jJgB42xUh0a5h7z2eo9T83VeXFY8aT+5EwmhgJXeRzdvYPFmJPOJR+z/hkw
XrybtEUp1en0wE+R2auaH1DZ1anNKmeEvNlwqsCGaj8KvGl6l3Rb3ywGf5ITaVLN651DUvVLXMxu
tioWSnKVN3JOIJtj8jl5QvNklZRYELCW2gBc6mUYZWuw1iK0hpxux4f/1R3Fvtn3zFtLgwHKYT7r
9br5DhKDN9claRPPqqR0CXp4IAmpu24evoHNTxMmQj9h1mBjWvbNfgXYiFtW+FRVjv20MLF+0MD0
eQ+KXyN0T5sPlwa0ZJPXnglzlJK62nuhkrosdDXQzBfaTVeA1DOyaTB2fXbRSqpBQklAGX6ZfuVQ
t/qQNBLbqzAJV/kYH3XRsXoyOkvwA25hKBzaEb/Q1HIz7VgSJIvsZr+nB2AkXXxHB1ARNDfXgZMp
B7mEvAAJHs4dfnaR+yWGXZ9h9d188O2CK3b2nZJoftsl6m9drvgqZT4mD3Onx2+f/+X4zkemG9hI
vDVY/h2FLpD+L1FS9jEB8j6Svf/I7ks9twpXnHIqmTzHs/tsGY2pljxw+wSg/mvTmO8toeCdh0sF
J/EcsBLsVuP8zlERdkrkjv13hXuTvyf1n0nKhQa6DZCxX+ncJIY2aPqSVpseuDFFWWFQP7EDc+g9
CH1+vjfzTjdp8DykPsxJ3nCH/wCwdr4zCbvpwha8/Fr1s/Ph8Es4N6IJufzQ4Z3BGTMCfXn6CVf+
fLdY0xlosd2C+iApzi6bpqzNSqCwR8Sk7dYZUhbjZECqgq4a4CSsoxkX1Iz/SYMPKZBB7LSr9kXf
1YblbCHfq8HlSBqxC+H4Lv/9djC+p+c0zoauLq9izZvHkZs4SQsDDwJIzdiahhODFTEbFN+IVOyO
ozKCh8MpS8Zx1tktIbqGuMGUgUZS8r28lBAv8F1hAqrujiqTBp+KvPcOc/EwrX4+fD9OhPpxOmHe
IRR1/A+NHyAVv+DAyuGK0qIyWnY4P6rkhIXdhAoJcNPCk65fTnQwA8qgaA+SgwjaXJqcIcn+Usc2
3EZ6oeNMqUyuZZvRakfbWP1pm+caoTcH0ghfybHPftXTdRfXaSYbeIbwg+eDee0bLepg6xR3Ruoc
eIi3ZOvh2mkBNklXgfU93inaT2djh/XS2lndMDXZylSdgDtahLRxdfJbriZiCJ+pmxDk6EJHFUzj
zejEh60KE391t2jF4fAzYwPnCtaC8Ou1L+xXKIPSzv7TR8Eh42BXxNplWfkJ8QzV0aH8mifNQzJC
02dcGykLBIW0bjKfbSQTQPhSbzFW+tbEpljv/F45UyaWNeGB+J4h9Oed1n4YYVAQ7iGXcy1EkbiK
ZCBV/RcJ0ldm1+7ch7SPaI2w3MqzWO15tbQ+S8mIwadic9SmP5Op3THrnbJfL6EPp5sNAC1t/yO6
63gJ8RGbVCFPuUkdLRrN6p+BwAia0VHCgyeGkc+ZOx2cAizdqIiglSBUN4tKHZspCULWWyFSOI7N
e7xp7RfgqiWyI80YjfoHqFmFbGht7i/nT+zIbxAripWn6iRIcdrh2xq1yUtaBs3MAVO0Q0fEz261
p3ww+tzmtpxOCxgYEwnNQL82ww6sJ3vVmIN4FMBvzCLOhEiPjokzKnezVZpYnV0ShtCXcw3Y6C0W
qXyQme1f7qbYxJtSxA/8gAW4WuIHoB9vL+q7lpB1TLGPMWrqpTEVS3f9Tz8sqmN2skLCtvEFv1J1
ONFYM33wXedBFZ303G84RtbXGhbaAeqN4JTE0e1mLxfvtxAXMbcsexXt1DHpLJdF1cWxRTHAvGFh
SXC24huTSLCHBZiCiwhhN11yrOnh08Togo4T1mDBUBcsMxd5ORBx0IPw/EXcxd1iiFizfcR1YOis
C1f6u3kdC2q3N2vT31Nq9stcUzues+txxESs0f8ExW1/Gnao/QvRXwntIFaiFVKskyPWWrZsByLC
vNAziOlnEP8hLYk9nNDHo3KjDBE+Z1eeA61BqE2dZwtVPrZd7qqcBzr8MuN1qhwgRswE+oh6q/Ze
vuceLIZZSUtsLl5sBRpYHBte53Js7T65odFObKnzDnK4RLD8xUomZm5O9LyFxM57BoS0ReCbxWfB
bPZSrxbqwWXgf8byAoiYEk7ucmPtY/ZOroEX0amUUR7JkTLqhou2koDxtSFSbkndaJJqRIajbGxL
5WBVqtz0rgVCz5T4mKloyuPwv55c9uHm7XEm8nuRD+rx1z6OJAF8qalFb+xGTa8eCaAO66emI0gm
LaU64B9L8mIYVT5d0SFnDqP6OaMKMX3McbtbWYSpehEEuJMqiZA4WRBCjDnyNBak2YUTeRiUWHAT
QP4HGkCoxsO+hYtWk+XUT182l+RnsifWijIiQuSKLSjizFWE73D2vDNGXbZyXMjbs+wRoTbVMETI
ZzjWINsum0Lp9vvjfP6ORBeCD7rL3lkQCdlrjcSrmJ97cBmToBrgQNwJ2wmqeOuFuGWUx3RV9Shg
QAAA/eKogkKH+4BXkAvfLrZj4Tt+spKG9ppdQ6b1zterHwLilIN8z1rZ7PBXxT3my9IzFVAzotZI
gKNDE07uEuKrJVIlBnNFR/bb8jyDv77oZnNz96zG/HTpw6QSJlgLpAjopzHVaP+34nXO/wmp9+l3
9Fu7dPmfBpfMeg5+UAIouGJSXe7E5ONs49VocjJLsYpsWjUH8mnyYPrrcWQfxFNSf/ggV0cqWKm+
YWaWW/j8KAR1SD2gLtEDU/+tN4MOUvwH1UZp1DxFCPCofVBQC9D8bub8WP8MYZFbKc5a701w6aoo
VW231v810vyS/orduK3/9kc3oCShWG/+b3KdWT8mGulnFEJVtHRImfWRWFYM6Xck8F3zg8zaEg3H
9hp+FHBIu4XfAZyOb01XLGbkWQvn/5RJ/NFQBIBbVntkOoYW/s9Fr9n9FvZGfLeH0WFiMhuLMkPD
nBaYnih+k3R0a3fe1ll2Gj2uyI8RTb8d7dWfXPnbC5/r+so0MoTGC/XhXwnz+muX3JOyIX6YdQzB
i/bLeYG9QySQdsTtml4VBWKLVb1SZ3X8GLNt/Dr3T6qjgz+uxuG7nJ90N8LOdyTx6ipROl+AF5ax
lKbXsmX5AVDIjKlf/D0uqPVoP08KE9Mb1feUzNrxXkffMNzdTXS2DRlhm4lJeuDrx34QOCkbYpE7
L377qgJOIFD3Z2DthiTSi5AKO0pm+eJk5FrlVtyUj394D309z4VonIRuRlUr/cPMQv7LhkzWWrrG
118JVMRiVoCgvCKpYShO+mXghRUjlWIBd6kKvv80v3HLLlWxFe1fGeYPlVI/L6pm9JNGvBHvYd8z
ETS4R+w8v8CP2XIUaHvPz3pK9bStWJoeyGk7GpXIhFnYApwxLNqgN3ZkyrVKe3w3ff4eH9wI8/BV
arHwX9WDm5/bTWz5tJrYMuLU6zlqJwa0MUvy0gYyQA1AhJt3xPp/egMWqGGfxkOoJojWH/vva+68
FFOPNmwsuBtVHefJm4GArtLxo8cqCmtYSV4k2S6ckxj8SVvMQtdp5e9DSb88DWQ/+PzMtJGJnyfg
YMndaRJntMdjcCeItgSsp8jDsnviO813/DAoEtGM48OWlrlzoQp2oYATeUdair7vfPkhIQ/rTpuU
zZv8PAD8Ob0Av3OSdD+81/K7ZeivxUcBLzFZpXqU//HvU300KBLGP9e48EuGkMM0lmtX4C2m7vF9
1Gkst8dFj6tGjQ+YxOo9NXo+fyb25OjIFJrXyabDeJ5vVa4Co7AthuMW9FNsDPLidoIFDxFGe/Uz
FAJ2bnfBRRhZca+zKaaYSnrjT2j2cegGPHeTZ+rkGXf1W6iHbXQdtOKGmBE4WDHz1jy5s263vEz/
JamskEwKV9cY8tX46TRuNI+X7H6Zf6xX353nKQYSP2eBEhxicyDgxZn/7xxFmCwAdwKzCgsXpSxa
X8IlH7edZ8NrsY3PJe/GlBmYMuo/h2QlYcGTrZ2STSGM8j6x0XPUdpe3C+DitY3J9sYS8ksah4Da
7iSMXI4lG+Vr756Wf0DcEwtpbblSVR2sIv5tCSyUlFJNGrx10UFn/6+4y9Eu488zYUUiN947V1AD
QDekJSjMyzjwxosV8dhJIgL674F8gji0Phs/9K+NX9ijwRYBjgIudt47Kc0b61hyS0zNXjKl3iZK
iZg/KWc1rIq9I6LEGdz1tPwfWo/qoMVTqaJlybJZgPaFkrubycESURTxz2VP0C2NQ0AVhpXNnHi8
1a99lKUdOZG5XEORWOTjDOZNQJDOe4RDcqgbTQkdLWex5PT0TZG4XocqJc5mSTCa4XI27qjjWh9r
T6c/Nhld8LseVo4Biv/sRg29n7Ph8Gy5KTo3uPp0iRxmgAuFo+kwT/3N6gIFpOqHYppMvzZbF9XL
jhegORgUtKxcawhBwb4zDkjIiUIDByU57V2XW5DZqROG1yBz+YzePMEihNZy9Npc6UAvwGqcN9cO
h+nOMLtQ2RTYnwwExhIdvHDdwixl7pGn+49YB5PQxb337paqywCf1N+aqpqEk11PUDcmie86zBWw
m9AORsJ/bckPv46JSaCB5dnuhjmwcRn7Nbvpr9d0sW1vsmasr7Ov2Ej5FkRzEBIcmGv8MhhhXlEz
59Fb5UOmeUvNHy6GkJnQdp2RpaIpoyAgGc3gl+PiafZWktjgk7owza2qVwh8sGWSqONLyWzNH+Hl
rEXDIA39oHzSpAWd9Eg4D4NTWbWu0lXDTN6KTm1mYvNmG4S65v03FYUzkR2NvBDZTHLD0DvPNxiC
o5Oe9QqAWtYCCIcHmO4i4e4yurOqjieMvel06fSdVcaD9ziH4CwZ98GZow3WANvZ+qFca+XQJ4xa
XK9LXlCxGG6k9+hVcVQjzupgqmiYVp6ztHfD8zWLjfP+hwUwv8jKKo6cAJiALE88exBHICuD/5XK
RvB+8GfrZzkrbsDZXHtYUyLovmG8T2AKHOadX5Vza+XFVem5AN/nila2VvqKZZkuY2q+GTh4PWBy
tcsgVLKzNLXUfzn9SGRKO4COUASndulFItqJtZmk0EdVFhBLjDzc1BpN7ViBG3xVz2fU8mCELGCn
WnCmylQ0Qz+Y1hMd0v7HF6WRLdMlfiaIjnLCZaxtIsVBgwalbQn/yNILpgnAzbZgxbO2uvEFXlMT
6TExFulhx38fElw/dm97CI8W3A3VWIx1t+OM/noV+3VJJBV0oqoNbz0XDxFHjyMpotu4zcLMuN/7
1ZhL+PkEJ0NfjtIpAD9mMiUK5p6an/l529AEGnDHEK5XQPxQ4pvdf2Bsk5R/OWYMhqlBZPWfucEu
ahVTOxFFy/hLpKTsP1vYG7psw2D9uqDDB55n7kx1+mhx2RElSqRDRzpjWLDIj8tBkro7Z6UDQSqq
AsciREHDRMpvqpFZBd12c5fMuSvI6/PdVmFzrK2jtROBX7n/FihbBNOWnnMRHKEaKQQS4KeLnw+9
QWgkFe9WyNFX2JoKI42Sp/VXvzLZgwfDAvFrKSgLwV7yZMaZb9eBhEd/RZkvmv2TgPitkf33xJEA
kRhlAr0XUqxgTM6O9ta2ISw6jjkEVKGThLW4cHdbjqw5CPZpavPSasDh6Z1MtQss6P79tz/vif7x
Uw+iCjTGHXGzT8ko1s4I+kSNZUeca3PSLsguYE+avJSaxGTvMdKDlPylDV4YZqIubplJboPEy24/
4VtIUZbcSI3gEC2Uxq6FXVN13Hkml7PpVbVLp66wEH11TkxH0NGJZOZmMvo4
`protect end_protected

