

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eddlQ1EVBhLWIw/V3Y4jUv/9vIqrPH4OG//oOzrJzxfxJoDe5AYwYtf4Sd3VIdakKHjGWL10tZxJ
4ECEoEAvaw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eigFAyj6GpLic/D0LIryLMG9xQfLbNW2aTMhx8nk48gxIwiUUV5O0RCi0c3WxlsD0Jm/PNvkmU9f
0bvLBoFrSTxK1CBf237YO6kwoV8FPGCIv6uN0rXS9lJQOPdNh2ZUFAvoavKMegwZ/325WocnFLGE
+YU4kz1iYX1mmK3UsWQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mnusdFYP+cjTwVO+sX1Blw6b4HVRZgRv6yA9tZdzqDv0sG/5WALWkeGj2iueXjyR4cWjsJaH1ItC
lJVwVFFXjpYvHwJ5RnZSqxv5F4MQSqH8KyPuaWJ7fxXpna2BJOvJUmLpfNOHHcM9ZtydeUw0FeC9
iaG6qychgs0JvDwxBvcNWeI54FWlrduydqedwrfELAOgz2Hnkk/tLLl8ktgdmAuHiBSlaAN8i7/7
Tmw44CbQzhCNPl2j2hqobn0a27C2ELHJlqNJpm8TlXqvKo4J8RYyFeM9H9JreJ/8JZ5Gf1n3ys2S
lY+Rp2WYXmq0OKzkZyIfymRWl5zSUC9Q8owcqQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uySJstuqi1YIYxsMDiwNUjJcaDIhlVqhon/QnlfUo3RyDfx9K7bIKjrz+E5jMqOrIwDUZDswr81x
cRDaji9FXOgh4P4INZOlQhXe8T+6WB7arsOA8Ipz2w1V2sV1eY1zPj1AXh27lapbQpMmsim+eCnE
1jY1XASKE/xreD8Glkk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l0UqkRkbyGn9mj0GavEkdTUw/Zw8lL7XEPhtCkfsrXvwKb+1KR5+77+E7EhE93Pmbk2awJRlXYwm
D65p2I5aXxW9fMEUNE0pZrhuaqpOOrPdC2bw4gaCcKb2BQm2PHu1PwR+8skPqiaBAqZVoUwFCZE8
LkMHYL9PggokRGZn1pk2O/ghNvl2eJ30v5gmurH3kQ5VEWU71s2ecSWfrCtyS9G29Ke80rPgnbMP
zifmkvX8s5FcVU1LeIe337473lbGtzk/tTh1neIkyiQD0Lkip6Q3stpeftQqI/864FlzKS35OASQ
wgYvGQgHNq1FJbrpROfsgNyTrijicXvjvpG0Gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37152)
`protect data_block
Wau7QSOO6Xh0XwGCqM4rssk9vIPBJ/V4TCe6+UK6km8UVLK8KDLdumC6cPeMOzQGt+JCIz8pJ0cV
Ex97pLbiBjIM9r83Pf7z41+RiBSS+UniCFE6ciDXfViqb0RoArS4WMNj/bnouA6qBvab/oBB/bVp
teGXfrm9drMsEvVJP0glwikQEBXorJZeA56+4Jh28ny7aqMI18S5VBG+62tdPgnq99/rFXYCE+gS
Mzgg7ezsv6lbYh4BOubTGWhl4bVMgzfUt5KOpeZb/CVGILE4xusoE4tMt8kJLcHcfrL7f4IiA68x
vat8YYQRftOzrGd67LabBTrRAxDK87IwbrgBEh4Jg53NaAyuH/BVQCZKM7jqsGr6VATn/TOPsAGA
kDPerfxPvldkzCcWdPUAGnskRLTE32OlrVdZJZSLUN0zRe6fmYnhYeflrLd2PINvsIvpVfnw7S2X
G/NENqOEC11mNfPnt3byA+FJm4ljGTQGOZSPulSQUqnrf3xjh8DtvXsFgjWw0fmbK60tOGuqojGf
0OQv12Rr9MnbfHumc9pMUKGTzii/fLVQly32kPdN177yh8S6r+fkFarYo6erMXPtgbh51LBhjnwS
9056oqjOMM8+KTI6LtKasGc9omdlA+9uvUxsOBkoSbxo3uue+CJ/3Dg6mUjDcwvcbaXpvbyfX1AR
x1rYff3e2rZMYTebg+rdwkovR4tYOXoyIZDctslpHKL7RJ+LKz79hII8TXx5SF2AWX/BumWfyQ6w
JdhyNoEwgg1B6QiaVty8AyCYP4dSs9HOaQ8IiFQ1Ees4KeRyQC4ahhuu+t/QQzpTKC5/SM1favm1
cAbGuSndGsNwTNLDod6cIUE1exF8WtRDax0s7axoP0bRl91HSMSmWZ+gbzkMmLv93h9X9n9Yx+LV
RPkhxlc+k/2cez6iW/fL+L2ka1voo5BUFU+REt8W7+I7tTzyaaaCLrYIpCSLNsHL2jZs+fW3jPGI
sajfZNrL+zC23/Oosqo7uu3Hk1OrFKp/zFDO6MyIsDPCGDuWdHA5/itQqWB2Caqlk3XpLp/bgkvg
LgrnFAPErnD5p6JEYTWJPdTwzESZBY11uWVW9yskktwiV1tL8P1DlsCBgUwLWf5bdGgGqmtU3uJp
YtPHnuIpuTDCuSmQzs3LOCWkpPE5WAwz7UecfD4pKKyDs5x7oBnZcGdb3NUL9lREnplvST3uOOuO
l4q/kDUW+DQn09YvyqR9gg9x+sHd9hDXbUqOYmZD12DSfBso25Ewt1e2PSd4g3+jrFY0i1IOxfRS
a/ohYpKLiYOIwy/AloTeDdIGBnR1A0W2MMam+JnimV+N7PsbOPk+T06Xc/QWzdN9c0MSvTPSkVil
yEFuDc6DC17JromMKhJYnzMe1UyAz3RPTRhXpxlLXStGEBvXRFdSS9QEd1IuUFIUmI4buQiQ283+
0L2Q7eKUGxBjO1sRuH+XtkI3yTbIfxceVkxGMf3rfCxjb+kOugwKK58o+Pd9JWtcofka53S9u64C
EtM2thTeuzStumXwMDmhgLigDj4q3Xybs8ztXPak85Gfm7/AsmMUZIrGIwfsaofXG+Rwm/qvXRT3
aiq0xjV0MOrKGzPLcEnzZpLoDyuMw7AqRSZVrRwRJpBTvrFGgLB1Ax+R+OvA9ctDurSMiadN2JA9
noqWYvuTCgrXT1qnfMuFkw3tq27w28dfEiVaNVaKj0aEBesd2fz0c+AKNJiDT7H15V4jbWfGABH7
OvOaUbvUYMssHsDsUUvuJSUjcV5wVGvWdZSXbyAr4KNVvFcLVa0SHYlw1MwLq8osFxtykfXmMWwK
UfPUCmTIic0pLIm1Z9nqopUIC2EU6TpBxAX0Oy46ilblOCRD3X2aCGDSrqpdp2RfdRc4o3Hav0Ll
iPCxnky0SkAuDm9u+6wuINSqdD1iLy1lzMc99OYpXJPv3XNd41lYCwk0vbGY+knkV4x9KpBylX7u
fZzhWTIHMfxYxceIP7dKR4NSik7Y2VH62f7S91A57SG/9TV0O9QtT5uKah9DSVBFvyK1lKE8Tzuq
CwrK+aasKqMJzxYGzmxL66RuXQR+9TlittYIKMF9Js0bCuI+67AXCtDQo+INChueTmOn0QOcwiZo
1AS2LO+UtwnwBktEQPiadotSQt7WwoLBKpl4K7J74u4WmHJvLakf8rFJTk7pfjXzR9BKZoVfYbCU
LGVzrqZcPOzIMizsgcsmKHRYG5RpGNpZ5c7O8a3yFVoYw3T0x7zsWN8VSTMwFbtdL8BtEHEe1rLs
Ab+ulEy85fIjJDU8jCwgk8JXGEbTeR7JlHhpN44eCqTUMgwuAGC/8qsKd8GDxc/tqvUzu0I1o+F1
mZiDyhXSwFIR1/TYXtmGzwSbVTkbJEfxtLuOk0aNE5tPTGKcJ4WHt+/1lV1EAkFx09ZIRrlohNBU
1gPk3PSA8x8xHOqrmaTcU/BZvyHB8OKmystYfyHfL0kvF4bjqA65F2meodRzV8YcyqZ6pOW6sr18
+PbjZ+l9hbLrD9wc5vJDSaEUpUHR+fUIywjNzgDUGNd3L2aFeiduYMBEm85uu5J1iKUxEBF3JQ1i
foiWoAFn+NwRH9nA7vvflE+G+af+MP84YiPZINlaH63mUpixpUiNwuQWqJeL26OuNWWHojblygHV
/BA2rsXE8I+U+KPTCsOK/QD4YOEg60ZUBqsIzbppaGXX42jIYOWZn+obHK7l/Qki7rnT06WmqsXM
VzYhvPtl2EOKih6IkJ89GlOt0RCA2+tO7wpxresf5RKKO+/Ni1MKBEVWrz/V15QLtykzW54/XRGf
mnVHY0aBsOyOgn3RYdHFWRNFGHuLR7vaOyacLdfRD3fPfMPybXV4Ht/JZ6MoDgvHeVSN9nTzoM4C
VgKDc2ZcLkQAKaWyOfmy1nqsYyjmk9O1juoGAj7z6Smf2l/x0NwNNHqZWLNuPM/L0a9W46UAyOdU
pgNDucjc/DPnA0Q2C4hcz4vb3JEEjgKQlh1hywSIQjmyVMxTujP4mUf+8wXefSh4nIBSRI3sYfr/
rxUh1B+vWcx/QVTGyZYh6Jc1aP7SMjSf7GTyPe5Ozgx5PW/JrFijHzPUCo97wyZPT6pTjEHmJOgg
kYADPByFyCHLYmZjjwztgjxPTHuxybBmqTFYMaaBVEM0jIEZzeXf0gJyOUJNJrZN7Ej/Gn38rCqW
S0oGeE5N/n7yKoqxjvUWcFLWlHxd5UlfkXRnB36ZUV02x7UnMhdr6e4s3JwO6JinAvNAPERBQR6D
nRpM7W0+O8DxBuDO1FV/u+Jilr6qtRJYr5gzmYnfoOXtXjmv7PH2AgsHBvRG7kQt54A/tCOoC+B6
8hrOPYHFMIuuNBrf4sdwq1L2EGo7m2om+At8xYpazEu9LQ7M6VRss/r+5wlLeU7oBAo+IXMXeVmu
vyDibTnD1GgLK0NY7oY1UOR66dbH3j8FtazfsOyuyRkGreH7H0FzeICrXqjJmyNvpIWwN1VeMbHF
Rz7e197FQZqhATI0lu6y3DFZuvNp+RAJY65bW44cD2I0eSsTiUH3cRMcEBsSJsbzrpueH8sWJoIn
sMJd2XK2LpIiL9DhO7XAp+dSYJ+tErCkrx+8zxlv7bj1/CbDYFCkT2BD7yOQmxsbnNxzXioKeRMh
Z84j/i/0ER4V8xLZN56MXL5Wy5Z734diXIdUGAsGQi8ENdwfhzfTOcDMMB/TukWX3fygbSltzNOJ
hSGu8hcGavwQ8MbCnDKuzlrM8Y5lQxmkv2WZKQHNNN6c/kWwTCINBADz/1wnsGQxKRuiQ5cz9J2S
DYWrFosF8gZyv6NVIyyG+ihPJ6BajDoICKGcqz0Oz45IQBKxvDd9Dash6tfCp5FcozZXYAZ52j0G
18OKmi6ehLUq9/UNS8hF0P7t3yEhUUZxrYBA3clpTA2Io6ZtGns4Tx/xC2/LgQCkw6A1ZBVRYec0
UXusPrvZhQ3irKwTil5+wUu1A8P+oNoPlINUvtglixJscpD/ZnoqskGiMqbxyuDubRvVtxyq/Xur
Ljvd38XDr87fxMvfQ0Ngyp0kVzsTKez98nM67ayOpgiMUUkTuY7KqVFUxYlg5H62zxFG+hz5FKzb
ODYZ1ZBc8WjmwXU2688IePrpJBA/XBWI+Za2voicBWiX8w67ns343f9S+galQGgSAVrgwJB687Sp
pYJA7GXbMZRdGFDckfqtldzSDb3G5Tv4iBelOA3Q/I7ZCqFrXPPfccv6IAoPHElz4J8ez2UKcg5C
3q5lHVPBJ4mhSpfv5jhKOzMohNb69AktmgjMJEkWMsazLDAlE71WRYB8GHJW9o3MQ004UvGa++eQ
xQTQxn8oqyHdT2INq1tXkanq7jWROMzZg8Cf5dAr3dl3tURRrAcaVVLf+FHp4lcLZajshCXoArQW
JTJgIMdlGIqkLv0cs6hH+vg+QgA9G38W+NRQgCC++xJKOLM7vKYKdtNByhzSyZiWy8DvAtGhamJq
Pj8fj9Qencv7Kzd2leXzXAP91RJ31ULfNe11qnx4GvKwsedcBcEEkxjJizTlUQmXF4kWLiE+j9fJ
oKPidbxF734zt2tqWOAG+okPFR309XR2kQQV6iYYYWziuJoQH55tlThyQ3eIblRYAjv1E7Wb2vAP
iRwoD/m8fHr0sz7nDmOH10KgH14mKU36XMGHdJuDsyDDGjwPDHxVUuntBxSlr08/5HZ8xFUl8iHY
+SmleQd8X2+p1pRLykxM4A+ASaQn/uko8egqVeXhAyZup/yltOSrrPSxYJqC31JX+VJSk9QtCckx
qimgG0VCbTvXjuzq+PUJ0rK55/2GB5VjibfX5HXRwpSXxH5RtLFtPCRYIWuRXNOTWUNBZG9HZI/k
WwRJ32zhavQ7pgogof3RtM5VL4STNaft1RoneesKifFJO4Br2TVYeLHQnKHg/sRzA4i8isteUuoE
eyM1Nn7aslXUDdz9H/iT0kRqZuEszjr5XJc+HTGxFG0tBjDy1IxElec3OypCkvOQe4hMubCdTup9
RfyMOEeAPPhh/Fm9JbSVhWgs0IWrCnfPPJrDC73ZHmi/H2m6hK4ssZmLpMbCNeNr3tJyDPPuSfA2
V6jTxXUyd4+l6QlOoBDQIgfOpjnchM3DMkMGq2s/kyvfFD7UVMNXvTXDTXchgh8Y5Mdn3D5qRSnj
l9IY29WMqDSe0XKbhWFWK38rSgl1hvD9jnYstNzsxvC5sThEevkqsVFGBWeNFwmMTt3m/jLc75Jm
XrtkP/Tl8C0hSdcFwTxXBSCWx2qNf97dDkQhKu7Ghb+ZSX5utJz1oWi6TMGlvCQg13whQHvYOjau
C8//w5iiXbLDyov7SNmboUzyj3odVTykWUPwCKlvw4xf5AOiqxFLyMHbGj22TMNyMm5ixGUDzX9B
owqxXBAPaOASZU6CdhZ/hDUwhpSyTVA7gsUgY6mFv1y+Pm1p+1YbcDMQblLGONbzjAxi0f9wSNtP
hR9TQaXC6OPhgQW2VffdiOSA/sP5X3YJ69YmlVQRRpTyCpDQRmFcVxVQa+faiibGcNl5nagaUdxa
qlTlNsQqxjPId4L+5qYuC5mMQV/8Znol8GrVzCfPQUJUB+xccDxoPug5EDWww1tdwzjcyePb0mtH
/i9MdFHe1orVlRW9D+aHf0m43gkVNnQTAnSERzEuqqXyR1+vpbKzsyjHM89K1jTBUBBNYUJD6jsa
un5r5qtYE7YlNZfddrowWA+uyDuN+skXqWqmmBjVLJ1UfjHy29CK8MHrWQJhBi0jrKLQhuiGCw1o
JtOpczkjil194ObnJ/nFqgQs601u4f0kkap1HEMtOj28elm+yj2KVf8GgO7feqA+BhmewYFhJJhY
MR19Bm+r1J3gpLkDZ0gWNtDRqph33HIBN1UgTluH9tHe388Ors5ihBp1L6yDkUhA+DjY+wWzVJrr
or8d/XJSJYz7170rdRrjr8VmRhGWbfmxHgRu9Umr4OMMumD+wsWe0aWG73p2O/Ky2GHe9WCZzIAf
lofUl4S2qqr5yMtGPInxHlNKj8sXRpElJhWp/W8QGeKtJh3VeR9Rn46SWvsmXN4DC3YP4pF9ev0Z
nl+JPQDX25HEoBX2hC8MkKmPNOXV35lc6dgqZuhV5Xi+7MtN+eN2GkzI3Jl93zWK0rxtlCTMxF5u
xw1Kslr4hU9opP/YBwHysa13vW1LMzi8rMUP5ZVDtPjEJd+/xJbgUA713/zzWgCfYgZCAwePuxsL
cIMx055m/VZ75GZfTwRWAUsbetXXj+j8xm/GQsp/uhzyMMR1Nm2gW3bD8YLDXjC9mAbnofmsv7iZ
ZFBiZx8Vh5gnq7ss1zNjc9niUJttH+zaTuCDPloP1v3Yn0Q/Cp5YyrZi04+RKZ2QRSWLhLunM4R9
DbgVScqiVK4pSMrZKXt2iMt+BIRq4pc5aYPe+S+IftSpLo+l3nX8CneBOoxxS5u5sgo9d3sH5XsB
ojb7d26z1hotXUXFjkwd74577GcqrIDtj4QCrPouMQ1BljlDmtmFi4GrgFvKR0hGOpLgvkdB3ZCt
6myMRYKVGDzs+cwNcBEqFo5nW50V7z4lUzeyNJxp3jQ1jzK9EN+sfGoHyB5ednpLoWsL7WO7MDlP
/DPjKPLkuVkm/+TGgS7p9B35ChVDJvlzbPLaovleYYTBJHB4h0tUw90QSNfH352lpezju48XrQut
kbGLgVWi1XyrDD2vdkDx27f1OY6gWjVQRDkEntTEnsKQs8RdZxUtVex+iGV2BXyWzXcuQenFwLZk
sd9bTo7Is7IW7LLbe4qRMQMZaCr53K8g/D29aKHBL2Gq8U97wjNIbqqz/zJZwRL9Sdc2MsyJd2WW
TXmw0CTrrCqD6UEOcz2m6wmKE/wiqOiuciDQ5a5FGHAPH2bgsy3hfhcBMR3Xg+LDeuGzFebJ1+Rw
CU9Nw+EgzV7n8fupLrs5Ft6q8YVGzn/EHCxOj147+Gm6TL1K4nVq7YrqzdgoSDkvClEZYwB2YQyU
y9yEuQzGQZbHniREdElY5d97mnrDDGwUS/KP7c7U307byoZZ9EFIlloLmfjhxcMzdeuFA89jxZgQ
uA1TKag3OfPXDLnQzP7Uf37DPEZe3OjUOgC2jpSljjoDRySNrqGYxy8uT3zmh4gl1779P1SJDb6b
D4/pC0oUQD1Ji7gMyCthjiSYL7ykmpjmBXGJIshO+aA+2ScTYnnndSNHIt2irVu/YOkhcoL+bmDv
vsNLVTjwzJ21WKZeUjnwdr/KQgPsFWksDWQfUvjquZpznOhWKslZ3mf4oZotl2+6/itYXqCET4cX
RoT2Jbnr1sdogSu7Fdip6QPB+zsMtt+lwXfE8BJQWaOGNaQUXPaf3UtUzkjDmR9/g/BpMn6SNr1L
83TFzkSlxBT8TkPOc2ju+eWffV8z/kTyit5evD/7kVJo15dLryNrHPkvuw0QldFf6WGBLS9ZQS0o
3GtWfE2cOs6TMK07yN+hNqEywN5hZW5dulhrsEooeweydjXBks2oXliK4LZptUn1gf0BQeDHerfc
55BEjI9kp7rm4GQpTyhi+IPuTjSXFmKCc58dd3yamTF07BgxFDxQk8zlCoNzw8SDvQXs224CImIm
5iA0mLVqo9TPBrIflAmPZzBsQ4k9nvPLschfmsEJld6rJrKA3FK/Qh6AbLGWlz3gxe97ohzp2ltv
9EJqA760buaH7x22o7jfVhNZ4DKMJ2LYoIvv/YFsNiSYbMFz+Nq+BuJy70+f470uo3MQPuklU/Uy
8Y2+O1HPA0B+TeS6p+4hRVQlR1qlSiZwtjgeMsFlB2rW17wHQvgwu5JrSOS2k6Wb3ld5oRAE5L0O
eUCRXiWhtcuqQQS9hMeevhVJZcbQdpYKq7E9YNc+2RcqCvEycu3AGQsc1XxD95oydNS4R4cS1Dz0
jIqMDxfYvYmRogSG1vA18ZomD/61m0jfUC0sqrVx2BdWI/PXhh7JrCHn2DBbhuS/L0lQ1Bwv3myQ
c3UvEBc4IBvmx/UCnO5XnEyXxWadM8IhoBjg7qJZdrla4oYO8+md1QolhXMSdPgYUBazvE+f2j/Y
UMBSlVFInwAlxenpSYRs4E+ikNVvnvx/5a7wb7yRdzGc7I3Ofge8EygpTIS6cntJIvvgdzNSJ9Po
u6BiSceemxj5sH1MC7Q8A5GO5gJVSZ6A+7o+95HPifjkUkm0i5gb0JCukKTv8cPFl8h4lYhlMGgP
rtw458N6TKEcbOA7Q54mMly/bj41yYLjC0L+KVVXcTa3uRRnDFl0LLMQHFcFdz21jGhdAEjUBoB1
6wfdpMDKKTrv8valvK2o0cemsuXtc/Ogk+YJcA9SFLvSzFHUmVUIEKM0dZVU7n8opIA6L/lnH4KV
pDu1YXOEMHutxyerMEWXqbBRPxP3cAZZQfRf2q+CCrUREBBRk0YCeu5S3zc84Eo82xZFHmBALJh1
9O0mUZCeJfU5KCIia5Nav4IVEZ9IfHIdw1VyCPFZ3A4VX2ZFpGeEgjBG0a4O/pehqyUryYy1EjaC
i3f1nsnOoY5/53TrB6NZesRLgbEhEUVC3m8qK8AWA4n+ktiHBPVzVwf9XwoiawhYyC3+NeRxPSM2
rCK8Q6CPZyv4sOR1+hNj6PWAm2Efczm0i+Q3cab+M6MtiYJLTuTNmC1EomIz5g95T2itVa3Tm6UL
GAXFXV/XEzHP8+rPtj/uo/sFMSoKFJT8CyhmZDDf/58LK/5DUv9j15p6pJIIMZKk109WdWhnmPDl
l5N6Fm4GhCi25dJwseRidY43/3CQPwBfdMSKNkH4sH3SY05UR+OvnwbVT8eA4a8Xk4Lj0xj/YNjR
8h0qInoLqDUA5Sta+g4K0867wyvmznM9V6FqzxW3R2DJn/Thmcy8lROLHK45UUGx3XjBMd5S9/77
NXQUdvfJ4N9k+NBgFuhP4+NjC9h2cW2cS0a+dcOAsDQhRxjlscEiVigCwqxfM4+UlKL4ISYt6gRO
8n6nYy18a/FZhXLtPrtSeQZuvzQNdBMrtkzeWHuLQtaxW7jmHj2JEWix6BiCWA826pEDLV01P3VU
zjEQMKc+PU2NCOzJ6TxAFSN+T4qpAvjvbdFzAMaLbITuLH7Oze0ijVi+rx4BUi7hQYSaJeHgR/oq
fS/tYfx46nLcpBskyrXc1W6mkSihMMXH+5d29oU4UGopQOOhkGC3ZCleDI9rZcvFqyXIyWgkHzTx
35c0+kELDjWqunixrm0itQRPHojyI+WV0ZOllsplsAwkWTkaPXAkfMXB6wi6GBAmyAc15BE4MshC
aRglE1M29nCegfUOAMp/UbeKjDD7vTBPVHcG60lYrWGFDxnZQgJZAomqSMTyBVykALkpcbk6vKYz
cqTlCWAavS5iyeRNU5lgWsk8It7Or5rDmaV6rn0R1Ji/ATSvWF61Jh6K6aS5SX+uOTAqu2Dr1RZ+
guUU8T3SIwugV1uZaTSyE2D3oyMC6w0AnyyRduHB9B4k7dQ+dJZkHOu32thB0d2oEmUJb1Bazj05
bVD7hfoGZPwKUnRK7SOY8KPv+CPjcRmRHzMS5Mfw4gIccMZaFt6a8BbAMR2cE10Gygowxne+SIZr
BVfGH//iTiHguDkee7hXN/211efIbUht6sSy5xyt5lCjFv8Es4lnlPFmd53HSIalnZXwhlUO30aP
bZJlTI1dUrmBVIq0YRboQ9j3uTtGLJUKZwroi5LQGTAwi5ZDY+GX4jqvqKBekkWeymcfuqtcuGg9
MT+DYR63VQaCGfy3p+6FzjeKeF9SQNwaKjtRl75UK7C9linRNBwItbsahOrR26boFlyMPJJ1sa4O
MSg2FK/en0sf5twCzKpCxAVIlKkzDJ8t1dTPqtwwOZdeFNHgsHOLiLlr0s017Xsyg26UbTn7PbQd
yptpacHML3hZdTxYveNzWq2PsNm+64+ZpPBWTPDCYi8sHpaPNtRG1f/j+YsbDF6BHToWQDX1ovTU
qqyVc0BDypKLFb5OyZTW1FuSvnN8uHlTBkf6ibMFND9yWy1FwiPiU9o8gVduxnKxJAZh9bSsOcgk
wdWX+ys6Pl/qLuOK15+zjpdXlnUIVy2x8PYBZ6LeYX5uwOqsVtJmg5t26HHvMB+NdCyRi/aiGtc1
+UybXR3P5Mj4yQLIqOf+Hl6Yf4cD/yki3Pnzi3szP61jZ87Z/aRiKxBgLn/k5M99uwI1RoWXODlI
6AZS5xfCikE9vdXl1FBr8eVlJF8VhQDflwTZO+qlNAApsqGd6hpbzbhb5FCxkuML/djynrF+goA5
mpxvEtMah55LOrT8dwSbvt0h5Mi1LunEHDw1fhVfjPEqhhGL4gtvdJty7fI1s5ThgBXX3n90gdJu
HbUj8sF3rjFcjHQnpxJXnX5jiH2xS+8kyXyniL+zs3TCSuB1iVRpE3xH+hXisyrC1o5tqvwSa6VD
9oKA22dkyM5oAJjW77rsmi0dw6l1yK3VkAvjbpC5zhfwgs0KDVOXu6B54TUogWp3+th2O8tjOky/
+mjKCP7a+EPSkkarM1mvr8/EiVIApZfteOa1qquRQrYFM0Wp/AUQ7GiyeGyrTweig9oOLOGuBj/w
oAXl/TguuxNtei6dV4sQr/d5iRrjWr0ohD98ACFVzqyOCsnrsMyfxB0T6EKkB0FdABefEmAJJNac
OlN21MJKY7IP+cL6ZNDDL8cwlb463sOCIdpJgsrrMP2HRHXMrlJoSf7/D4/6ColzqUDqh1OXxRbE
bEmMQ7TNjUnBA7HUnEpxllrSSWAbJ6jgXspH4pLCZuuBeO0eTFk1cv67g25gr0krD/2l5BlogSY6
Ogk9z+MBG78ipUTauLLkOZdl3uyWV2IDHul3bg3dFb8/C9tHBBONxCd62MRp5C1URE9ggzzu/LLp
RSSJPwxIRviKdLUEfs8TjGXm+Y3QqaclrY/o9x+Dshz1QSSe6EDr8DghNrdh12Izd5K2SLmDuiyi
mZcPuokgojjZl6sdV2FdYdczbSXTEBL0427Tw+T53exorBR3Gd98gk8z0kfLLHxVMBLF9rJ3Kz+Y
2cta+Nz7QZFU0bzNSEm9Ok6WaxmcbCFSkuWiq1kn/eWZTxfHsI8axlOV1T7NDsdjD2JeMwpqhxaC
yPj13ZjdDdnjfk3TaBUJ/PydSysR+zvpmuIQ5+bX4IhkLV+FSydGsYYaW2Zj+aRqxnVjQk7XHhLg
i6H9fkN9gqrAFYGGngRNQHOFcPPw2VHtsjDGK7t9OLbhTDxzf5Cvr9Ui6Gj3ekWbJwP1TKdWzVep
uv/xGmUQH+Oll4Zc0wguTYC2uXvZLDjICo25M7KrH4wdU+28AZu/TehpVVm9uFrJwGx2S4fou0IE
+ZmqZ/g2U9xkqvoTYRBrKhx6t7gE3WzL1TRoCo9zqrVIxRqFnzJVbJ1Z/ofVh8Ld8CDuqkeO6KCk
epIzkQbfI12qi6CCiYC4dz88DdUcq7WRonFj50YhUj3Zy0eS4PPpmTDwwVv64cFcChy6nH6MI/mG
ox/6oUJwoI/IiD7dyzWwYSwSL6jrg0ls2PjdzuXWSwXDbPbjIgmxj7maWpSt3DbFMhMpyo0cK+xa
fbuF6+1rWrZNUMDcnEeYxSFMDtePmLcucGV9ZylHxkuY9EK4ncATAdENlKZWjNsg+yGfU1N1kyso
YF6UrU/5hNwYLuu9B/9piPlhrn3gFZo0GS/2GrifvlA2LH1RS9NVdtPx9dEXiforvWSreZ3Uzyps
mA4slhl4MWHkwa1IhaobFVDkqdaeHKq8rgTk3NcQ18+rGBdWYFBFFjvb/7sxXhiCNN0bh72SB53/
I9EuOPOyiteu0DInmT4PSUPvwUMRN+jNDkC+Q26U7hV13qEYv6V8ZTsfqbv1ItFWQmKg7qLeVUFU
lPS78Vxw/PnKmDljNoC9tFok97/tBzFDWsmyW/FMvFe2gX11rN3c8jj5B+uyda7dRNDSVwQ0KNuC
Vo/VpngPg/oi1pj1iaLTY1QNA8z/HWbKs++bFg2KOFSALGcYTwM7uXNV1ef81I1W/xvEch5bVHjV
KuF4d0o2UhkNt6SCS3aAzqPzwwsi2Tj6M3W9bB7QYa3rBpA2SoyCBrrDWsFpUB1fTnDRFfCSaNvC
B0aAS8BJmEZbkf9dnOPLzdtgjAEatpqMmO3oBspPSeNHNH5eTsbMFxYYE/TJrQF4Nv8laQxtB1C5
XUQjlOAroF4NezfdHq8pEteIt5GzCgglMF8Q/dmC1qiFsCTWgh3RlVOz5mgBCMhKg7dSgG3k+GHg
lsMzNqG8yKI2OEXNdKSVlb82jlQzOL6qLf/xr5VDJCpVKC+QAWqRzksFcUQTjWS8JNwUopnMt8Ps
cpFTzzQzBTKFnDrNcOi6/xsfzz7GCwKvHdk4klfP9v0KSJy2MED8JhoH1EzWTsnNVt9QMwjVyUXb
2STmHLfZTVvcNatg3MDxEuWfEadYrQWJbMZlcj/b5d8pBLMEVdK67bUPgszlHbbOAsvWIvmPZR6Q
38DbF+wLVv+5yDPqXlDFuZ4Rx6VrekQgCfLOXP5VOnDBZTyFzFAbBf9wKAOeyrM462PH4QciuI5g
UY9VoJ4cCfBvSKXcF5c9lYmw5Z1zlx0lrTgmUD6wTsShn+UfclBXVRUiknCIthqkhxd51Nl1v0lL
YHYtLA17HIe+YpLgHEqyw07Zh3OVfvNRp2XGVsuKzeiiACPv8oePZ2F/ykIrsLrlpTkFD5PZMnsq
wYqBtauDi6s3/rRlf1IQ8/COp+2jsHAXBLBKDF0DwLshlo9r8ksfr9raqE1QEjUWkK+xCn2+NgPe
dceFsTle8i8Aqvd1ILSzcRGk5esxz4IlUQ8sHdZoaCYTR+/90PfjAimGCWYovHsdjKx/E/nX6vPt
qfXhNbuopyqzmfM0H/Pcrw4G1W8lan+to+GbrOxIagKZ/n5ADlWzjItRMg/h1a+Qn9cOCF5qv2aT
UYduyVJAW5NrXOlj9la2IB7MMMKNw4nw5CiyCUHM/emXfEoXO1Pce1LitcT+Y64LzcYjTcS+213h
e/JEnbHmGWOOKeofY4mncpX959S67JjIuQ4E8wSyM2YGPQBchNwf1iya2mY909DLzAPfYFBBWD3i
ePexsEGab0evr7vPtUuj9hUkNFOZabeC64iyq5KfyEudU18Ueg4+G8OR4QNR8pLYsbanWY2D4b+h
tQIAGeAC4O2SMYctXYEI1qUlSzpVQ7E85bsdvk0yCAAlsbS8vofcHfSvPg24rbQiY6JnkPMMgDhG
+3Diimbxytptskk4iPYUOT2T11RO6kAgzEi8LtkOfzQRMhqJynZgiL2y5DIRE4GqAMn3+WGR+ne+
eoXuDHE3aor5PjvGnppugv8yJzQVYj+1jKvcc7D1cqyWYHjt5ZDk9hIxlhvqVnCxEVObTsihD312
dR/UZ9fKKLOiRpnUQmw5od14tB+x05JAZqzSDBLDY6ki2MzZLQLB7IM5Dkz5GLcpMGJ62bodU4BN
4BixadnL2MJNHFMZEAIQi9wCKoa2SbV5zSbpr2vya9g0VA3hF4Y7EvaLkIo8qlcjTLpydIJ9tID1
rckp7OY4jYMJSKH+wduze0k/Pwfk+1+rJgFwAM0QoxbtiBD65QMr9L4nv1frmcqVeD1auQAzi4LI
qE8OTcuNzQdFB1/ngkMzZggPBnPWWORW5KB3F7uSY8CeTUNogrlc8RS4PgXcF/gERvnVYjUcT5/O
TpxbqjuhwGc9XoCMMIpqK3+0HHFwiD6nfUYSRJKDnRGzWRzeg8OMw2ncBbg0yTmVtIdY2oBJcaaE
f8qhAgBcGJlqB4XVS5e3Jve1srwcxy3l/JqJUQWT82SmxJSk8qKbGKGOPVAotXMcKBXmmKTIMsip
XiapPWE2Efxh3mwL9qpi9he0aV4hXFfKBFKUfq0ibseCIS53etBFUjKXXx/1ho91313RCzAVWCpx
JmJnR4BieXmK3n4Gxn3TxHDnvNHIlTF+QDYkFs+yaU5WXoCB0U5o09QBVlEJjAP7P8qHYFFHLSIp
6TxAU0rlK7pjXCrvUBZ5g0NWrzW3p2YjvY3Mu+edT9oxb8S1UZODOgi7574PopaTkqh3dNVMH2Rp
rQDjh8PEEmyA3pxpl34b0px2tYnm+HUiA/v5Lt0xhRonOPAbku09pQy0K19ARkRjgiLWdKRe0Yu4
ALIkPvBSmEQAM/gBh2Kum8XWaLMqLKm4tLnMOR53B39foDnSyeAigVMf+YZ2TS9mARKFRxl1e77q
ffiK9u34awIYfrNq+EpaDRSh761o8vq3UBd/PfDhfr/Ck+ONhC2Gqp7sYUJoNAhiKpw8368pQ+fD
7ISHgH4ZFtv0VdLh1iaFcI/+4hEMhpjPgK+U+6zhEk1ItVz1aLEtLsT7RM09yOmiCwZ9p5HosNdJ
j3NmjdUtVfc1rrV47y5pRmhFuK2LV2vnQe4gGA+iZYSUTE+y5FnodefPI2hpL4QGwRVjHfhedqh5
k7OIcW8w+l4G+Fg/7fEB4/dRXQRRvFLzqmUOA34e3BOgl0gI+VQlKyXHwwW8DDXazXe4VIh8rW0R
Q4p0gtOYjSOP4csHBp3fDDaCn+LRiTz+tWdnnY2CE20sDorlXwPC1D6x47dfThP/plE9b78tE4IR
Xt9MX5sJCS2GDlNPSov+kC1Ss3KIFeEFy1l/otzFyuiojxbOeJwLsLO9fr1LUgNADuurwpsfYijb
BKMNf1kWGHTLBQdmp/ZgqicpF07uodZZvZsYnhLwNc0takDYVQnqGRih72Q7zd4IRdrX1Gb69wlM
N3Thkz3C08X5ybR6Wtsqc7xlg47//f+QaPvRDz914rmrxzYmIyssrsCtVcarwAzIpY12prY+0C5Q
VAKbXOnjiFiN3kkk+opueQM3JjhgowgzV/NETJpBxD7aHqYQ5kUGuZsR0xIfZUWdWpG3RZKKMyvn
6L2jEQOs18AY+10GthI8N0N7XU/B9BbEHMJRHYVSBLjNzuMiO9LK847x+W7V3s8E1/yMFRRIn8cs
QsENnCd559H1xv4btM6XXWeKKeRfu1Ztta8G4+Usp62vKOxXwdc/RA7eVRsnqhzVbiqzN2pvzwrp
DCR8BDP9C9kr5JwF/i8N+hkj5rtveq9WjBT/6sbPSG80t4v08tlty8+5lLv3tO01cHIz+5CcIR6/
M8thwc9AqE3ahSeTI0MZyEKQHVQpMd97gV2XynTbdEOWAVdTloz/C5lfrbOnDG2jRBw/ua9cb+VN
CasVhmU2HRFHfuCDr3Kkh6pdJbk/c8A6gFDERNL0YwgdhTzvMzHGk3j/C8fXafhfQD+2IXwWZoCQ
67BeopvFxhQnZgTiFvYEbCwQryjD6EJ52thsTOM+GOKHUoaOX0fs1ywO0BDrDhNE3/8/uB4K+EDj
cQrAf0upN93z7IyvVx0y+PtakZhtnuPCr/Jltg41yIMB6XWBbXzUYUm/T5dum25vd/WzgIoKvIwW
kPFXAMtctDnsmfg4USWbUCc8W/WrwusIzktfMRL1CAaSEmzS0a2pG/KWYOF3oSyS595h6cFrUiSd
LEr0vw6di3C7GwYHTomr+4uSnUBeU5RvU8DX6EHJZICzgPWgI8nry+j58peZ0tpiRpJmr44fvTL5
KI3hCdu6aGqxQavop6L/jSIO2LYCtwB7Z6ETr3NR8ydAuFCmgBgGP08PJk2M17HRFSYf3R3o98R2
DfKcB0b7ukr0MFHTi87vRjmjZc6bzP9ly7UF7cKSxvCFChH7EpriYfctecN+1yz2Zdd37Igrf0PP
+c9ojtXHFS1Bq1o/KuabWOrwE+IkNqyyALUCfAxprpV6MxiSJ+iPnFR7iVeoSpC0ebifmzEPgwNd
Metyvj/1bL7Pp3yJvw0EYKi9+MDhdMYDYF2rl8HZQLU5a9dkL3gGbiTR+2G8izg/Y/j5FbylNqNK
vhCdnj31dCGi6net9PZ/TatYbMYGbDpNFNe4s+JQR3R9bAKAlfTFOrLaHcBNKpwxQUO6ud2s8tV8
4aUnZYJETWSf5GApqd7z4SSXHAq2dtz2OT88at0ZPRlfQZRmvYUjYVXm8sR7XKSseU8k44AH9MLY
kb4nYSFFJZmr+X4fmYSpsNIVU2uFJRdmVdXcvsY+3wROgWX8LKvbEd4WE8jg10cH5hFfu0ZTP3qt
3vWgnhcyVme6VDzSbY8Z49PO/1rUTT8JaZLk7mam9TwdKV+skR9HWGYvEqizu8eoTX6FKdOhFS8s
BEkdXYvkJgGtjWQg55bogH4pj6ouEvYPCeZOsqKK65KrGezt6eQ4qLc2EVwWHairO3SmpKev3zd4
+dye7Pzx2KEqnukkz0tMUMd4NydSgub1c7Amb/HQqE6qwxr85BBulgpQnu04bn7YG2NY0Lb+wky3
ys8XR0FlS7T3g0DGqB3C9NbQRFwL1L2iiFCL+C9XAiiUrOBa6SZBbeD9NL/6X3xvo5TLi/Lx4Y4h
/DQneLPjogzysYDz3Xzb/nQEimVgboxwbrA5YLIyJRhfOhTYPLNv1GyrJ5kKt5qhxyQolqV3EaTg
JP5Jfhl3DMADhsp3RETUqZLgpbgh2NaXpYrmjkZSEjPVTCspEgEfY5bO5Q6P91Te58g4FLay7wLI
9FSviRVFjXrmbuOSYqelHYNNrVbetfKzJWsmrP8ONNPMieXmCrTIksjAtM+nAlouMWCILpF/nNba
PX6kS1NAgIHoP6E2SdJvfkJc+GlabCbqzofG4iX3VHX0Hve0WrGgMUVshZ5vAxpaEU2kQBxe3Roj
6pcqGboQPaQZ/EHk4RbtsRvvoZ07KOemBzLWcyftVMGQhzH8dosaPLXCPXaletJM828sKp0Xp5Mn
5REX0aAQOIJW6zH12fA3ng30GzI1zUYV94HjTVlmULfxP0KS4LnEVN76W+oO1q/BadU5Re8d5t/w
3YrLl2kad8G054OeCtFML9q80iv06OW6NDGBWHyN7RL1zZCUPJMnH9dmm8pCaCF12l+jfS72Q53a
cIum5sklJ6TceXeEpz5fwy/u0N3/ZFn4dgGcrkHan0vpELLFH7CaUfcRcDo7FR0LT2qIy1Ikxb5V
vc3lR4XCBH50km/MF6pJt1DxmUE9CdMVrF/cIvxX8LpO6jagOITbwFcz/LMsWAjl0/vcBqfBQWYY
cjGQHK4IqLZZ3AQqLkSjgmrj435kAiG4FynWvqiCDg4VAziqgeMd3DPqIoQNCTzSShFizeQEJjC5
qXAvW7mMzvJbDJta8W/DtBVhwDRXf3thsKFw33UBmF64NHHhOAUa1XjsiYxaO6osSCJroX8d3m/7
JJI+pXWXKbk9+xEdmHPgESsyuBFMdGAUVGZTDU24CRhUylC0U+qHi9p9fLuwDas+7WaU6LqR2eX4
tfhonOCjTMpgdOLH/I1nku5PLHhosB6HAcJ/TF8/HdU4+ypSS+rIv3KFNSHx9Mcd0D0oNgeJFFBN
TlM9k0dJoyzHo55BAc8RQ8Mq+Qv/q8aI3pZnazk37Nc1j6yUYBpXyKPiUQUSwz7G5iCx/GitnEch
jWGYvRNKgQ2yNBCZwQRj+9XmisR5CXHo4qzfX3t/o6MzAoD7X0MuDjR1g8EbPpzSXHBBnRhlKMom
A5BxX6LXaxyvN4RsHcVSYPJ+Y5KCXiCMf0VvBzPRe8FNE+iMdz+aHhqtLNZP3rnqM1X1Vko2hkGu
g4avB6v7b67nuVckRdz8Cj9QMYEeg78HWcRxN5Agp01oIzT8FSbhfw+r5UEjnkZ7NcD3oCadltJ0
Ra9JKx+QmDHu0ac8R+2I00Ckd3HQBlmAaJIaoFQ/iHZA6mM4VTZmpk8CrWERLtjvDUEavd2R7xDz
THwP2fOR7gdaxx2Nga+YgI+ubrfEl8URwQ7DbfuyYc8qc8/A/emjUFARLJ7cYVKQCRu4GGcWJIh3
/WRDSOjdRi3Ia2knNNzazYnEedDu714DGJGIpPHFQ+Gx3T6wVlcwOdreFM5kImMerpzBE4xd50L4
a4XipaxHUvQcOCQkluPRFJL771tDzTqhRVJbfzvQqAAB58rycjn0KYj0fI4AGo9H1cAIRKu/2AGO
xII1kB6qmK67a8BebGni7LaTY3v0MkxfaQ69eAAeG13VzBscm5cy2on5F3kOdwl6+fDxyka0r+CJ
n+Ypj2V8xvCX5ISEpdCytZqBYetQJJMbm5iYCkSo8AhDSPAcoH8UB8oCjuLbLu+K3H+2fA12VMon
gmdO5Y5AicDBnqn+X8h7BlRp/dcrGWMgtHEZgwNgxhtHcu0LijD6gPrqKrsUhdGb1insStvVCrZi
cjCzv+Lu1119fgav0ybxO75cdTqr0psMwQTwhaJ1IvjqQu/juczKWjL4X9C9Hpsu1R7Z87k46O80
8m4pBcqFNPkHYMn9r4E9juLQhIrjzIC3PDTsQjXlQK9Ajf7nf60PutQKMDHm+oITUO3DkId1r9er
STHTf5TkeB4ySuDvbvSReCtO5MKbNDthlh71dEhR1dvaqu3o/K/lH1MeIjYnGPr7ePvGVx50AP8x
oRwqpQdmO2zUHRMQMQtNyRw9TYRqa1x36shILLQ6H7cvcf5DpLJYSv6VxnZ1ajk30AuHaZtaqfsy
eEfCE4OJe5crfGz6RHxxicAjstFR5ccv5aM0nD2eYvWYWegMsyys60CEdNa70V5GzXn8G+R9q6V6
W+Fgu7OT+wayt//sWzDjeXEjUfKrfeBrsw7gGOZtxP1QYvXLf/nh5mbs2RZePHPIZCtb0EaNyTur
ynNpsD2pa+BeaUUqg6qy7yBhR/YDphi70jHpxSS0j5vVpjSAFVgiKEqLtyYJ+6eYXoWGCIaUBGiq
+0JlYvDWwIN979J1M2rPljcgVHnZ7QVSYyDqFAAlYueWt8NWGkC+A4sPxyMQlY3N7uKhpzRCSVMj
fCPBEvmPgtnTDpv+/ZhWSITOorRpnoJ1knEueR1JkSncQji7CjoBSu0P9/kgk88p27phZOFpnzTX
CfR1nhTjZZTVQ9qgPCTdRMDupjIcM4Dd8oUyYWQJlXdURJ6qRTZrFzaz3Xf1CdRnhcpuTalkrcQT
LcLrQSBElUCKltFnj4sLeHhFLU5STmve4pF+SW9HwIJrkcuMVDotQJDT1+yU8cqdpzw+iXKnIaSB
Ycfu6Qrl2jexqGKbm04wvb9NI2u31JQfvlfyi5M8zzylTPLw0pQ8nmDg0pcGSJ8+9c+z6UZxEzDN
m5KA3ehDi0RTF3TaAJ7DSlfP+4T1tAB8E0JxHe9+vkTrMFz0QZ8nL923QtqiDlQraSi3V8YqNEw1
cToWkDB6HjtV1gf4sXpQ4g6/8IFwyPK4+KUxoWWYRmXUTnORR7MC3TOateq3Ogx1B5QR1/z9FOzF
3Jq7lrRwQ29qtXFbypib1hGSeT6X1tjRFkWi/7F7UOc/pnJA2sQEmZB4Z/YdFf+JzW98/DjPVDse
YnrhLj6o6vatJJjauNYlv5k3waj93nUw2lF8QpiKr/AQbHonxr5dQ7sLW9keWVHPLPQqbYdtycxE
NPpMufoD3FWXzDc989JL0PIAUTT9IEkmOww8WlOaHPlxYbGCnn8EFts0pas0izjiGHjNvp5DgH1M
1QNAjRep/vTUcpaL0ueJpAeKmnZPmt7wXGD6O3RfpD/l7Nn9bl1fF0cSrVdM4Z/2sqGZaYpQBjQ6
QMZYnmQDCKJJ0FvQuu3PdSOXLVbNr67SmTpK5/YvXeG3QJpPUU7At6ggR9CtCGzq+hcsewkvKzEb
QD4BEWSWC4PALla48wchRBmJxnZVYBEcWH8SMqq9cMaLc5GR3PEICMTn1tHfNP68x/WtjGNKE9Mu
DICw/f6hD+NxbqfMjN5xe6qJQXHvKdyPrOqV5AQvftpHTNtu2UrFHsF3Yxmx2jhEwiSbMmSIX2wm
RLRfiGEVPCtfaK32ZHwwsEoeuDjIluyKzbWjODs/yCWDETkyNzbYTbweR67urj/0ucsggkmIu8fv
EZEMsT+eoVbIVyW0ElwX9v2T6rSZWOHrkpdruC6ecpmyNlqS6vc1d7Qmtces8+g39WMseS6IBN/A
aePLrFhfJysj4cPF9rGSp249CVTW7+GBMYd7D/Y977QZ1JupkYN89xfn4pRQ2zu81zx7qdb+SKXE
d/mvQ1lDCvKAX59do6+2k6ObxJq2gbXDNuXndcTwDhwU0JrqNkfrDWKc6Z63/QWGqFvxpJMncdCy
4QuMzzbpzU6eEE0YK4F5ONvu8VQovpi9kPSem6z9oEhWqxgs0fUYMULbv+DgecDg8N8VQ1a+rcDj
qkgdSADSCRSZBGtwxSky/Vjdf00Z9cwm0rPhQy0lLvLit/RBlerpK6FJRYeutIALOG4CAKzpyNw0
LQpglIW5TfqZfC256zJjmHhE773m5QCLUgNWmvPwQbRHt7Dahr1E3a25eJuN7ZX11VrTx68HqFqN
dKxICC0oueoNjT5wcYaIXACXY9kycsAF50NAOlakOznwVDpU5z2FZXOHR7Yd72/HSVQdAPyK+gLK
N28CadMhqyLF+nSuwN6bDxapwuUJ4JZoEJ9wQDJ2SzaYn1hOZAdgDkuJUhDml5LnAUDT4gQB3nwq
uBsgeLryZUfTnLsg4HTqndq605t7NN7TsaRgmlEJnSJOMI9neBgzH0slMPCyVGkR2rK55DRYmOo3
R3yK05ujB2t+yCKCchi6rXJy747VFmKoZxkVQoLioopg8vZ+f8853DbJ5yNli/gvD1IWi6+FlJ33
RaQXpNNwWHT9QkMEwbVIf65WWh2m2sEv0E7m/A+0GrGpVYk+WZxro+SiyYJQd0wPJ0fKecs1xKgl
sQFonPmtxt9p25orZyZT64JVxfIJ/Ip+RoRR2Xp1/OufU4MH/nz9TGLguqNdiEvDHpPs1VaMrL2F
kVQVGB4eW5E2yTlbc+dNiLMR/bMW11ftK9vqsJinQftAL4UEoW47XKJjpCWVdRbH9hmkinonnXBi
GYBfKZ4RveIgYAV+MATb2vYcrEhUnkx1l8n/kjJGzfdEGhT4vUjHi6rLOfB8ODxHVOZLXVcpEhB7
xDvZVTjD9T3KGzboNLhdMiNEtD0NgGtkaDUuBHL0wSWZNPuY6e8K5XXdn8EZ2kcRz5Yg8Hm7pU6L
bjEH0XronaRxkIz7U53pALClsPEs/t+lzK+M6BuQuMVTOWuCnev85vxoILRGwdKVXl6FO2gwQNUo
12CC9+jTx2nCMikNq3B9lwBCqBkXNAGW50LxiifKr9uSi1+6dKj9k9BLdlh8nIFH/FtBoo5AofPr
jEG4Xw0yV7I60Fk34cvv1B9q2sGVWa1NMeVXs9a4YGfXJEWk6tP0/7FFPUUig0yaZ9X+IJHfZTNb
MvRsQVkZLvl+l9ATEzv8i4mti98qHBxijswboPcalpha1gSVpJtqMzLonYaJucC3uLhKApUHFo7+
BSfXbSxNGV0FVWRnJXtxmUzH9pXENSOISwaRXKrZNb0AfomKCTyqPORrG0UTCH5iKxTtO/mwUEHZ
t/dlMS2VnUAXz5sQlBjJ/gzrg7mycM+KFZavFo7Zt132TUk+qFmwJU6fhqxqWHCiNAtl6Wy9IMBS
wRPSA/nqQmIhQATgBvckqPorGywnSYKey/vkbs4+ic2QMMTN0CxMxa/bjpfCKUeJFrDQPmpP5KxZ
HHF96KY5mJCbEkLjnajqU09Ilvy+OiKO3zFstOJjHqB+fDwZfy1lcVuVxJ5elUiBhwA/BrQGUogs
yoDhSGgygV3n7zxQhgzvIMS+yN/QYZNhpKlSt+0Yq1JVZPJW9+SWQdz2D7crf0Af+Iz/JIy7607o
C+FJvu7w980fFhru5qx0sMWF9dfvAKY6T2D37g7YTZOPsP6pujUxNHa10JGQf3bGvmVKQyW1xDyT
WQLXVYlAgBGqWDzOKcQ0lPSHbUmXDMTeyfR9q0UGfPnpwhvqHD4o1ixHlSwjg4pFFaLEGjB1eIdQ
5E1E9EtT9u2qIr+iZCv3SA7AuqK116+hlsJEcfHs0r93QnDJR4y+14W/Dx9ACdm3cWzGODej8Sct
VJcKLCxALA6lEHlwla2JzmaDxN9t0EqWlS2Oa5rK9jPG/zgSiom6/LiCr/z2d+3bPDxoFJj8kGkU
gn0i1da2HZFAn1Xb/D0bij7YPWNMketCy1igzPQvMAGx7FBpxv3Op4Kd0Tg552a8Rt4aeiEAznxA
ki2B9Jo4XX8kOjqD5+0jTFq22lJOLuPr2riy2Y7awLak8pb1YUWBEViKy+ju2wXjpoS4QWxRi0r8
4atjxSqIRVqF1g1me2qY7Fchq6EgByTSHweBzQYogRy0sNHdp7eXpdL8TWC74Gc9E4v1d6++o2pe
RglE3kdaOTDFyTR7RiLwNfStkNbgOKmjE6GYNWeVTdBQzfoYKOLMSDLXNO4pZ7RwdoFojWAHkaX/
DQ29WQaVhs6SwKdYegsKPs9Vml6Zq0QRVrLMXLFPS0iRuVmJbuzocPf3C+EDSl/cLEs9a7VjOnTE
aEB2HHfHOys+pSdwwaXw8hh/XyGnes5L5IQMlMq4XvxyShgC6QEl4QfPwmnHCNcQZjTsGpZguUz8
OZgYMRbLs54fjw8KkC2JfRzaRfAzYm/FI2WlkMIDwW2GlXdMdXMk2HPsawLD/8BRJsVdRYfrAy2+
YJ7CWfB8K0JNJ/YlCqrYrq4gR+lmlzqw/HnteWsI7U1ovWMQXMmvstXxstBGp4Ck2SoRZu0wvulY
GI8hRdfhKD+NRYTfeo6SLd8z6AhZ1ah8M194NlRhY20BoO/pZpnlTjpjgd3lHOfY2KUmW8KtoDRu
STocofH0rLR40+n4+oxIptpOLQsaDsrcvC0FvOFLKOx3Tdtbp+CfYV6i4I84oc33kLTBpJL/bQLE
bjqenMT2o/wqUx22wUFRFPZcXiL32bguAAZL5xKGZvn0FtK+B45cIK50T7sanPxpV4mVmUURGQVN
ZCHRYOM4zDqgEookhnGjUAWmUjehpFs/Wb/QTpSe7Kg7+qdPwmPZIaIkVqiX9sJ9SzDXlfuo5GjG
KHkG/paW8ZzJImFA0i2SeGrupAGpmPrF7O5DKQPMcYcUvLWjFw5JNwOqYV+3ILpgp2S+wrRgS09G
FvcSArlIQ5uKDbkEEKQYquRY27YBUHIRGpmWDINT3FWDg7cgSnSka7clbCNCiFNJCeo+l8UONySX
j9C932A1lSsh9s6Koq4zzR8hKaXzqVf6M/3eCpMWQ1QFtJquCPWKB+KhNc8CNAm0mmIquJVttKOs
1w6a0HSwyp0+Vrv5KknVW27ac+IJRkXhk5hvGctOo2qEuiOUEqTi1KRNbf/U5Rq6r/iVZ5DJIjA2
tawMjK64wG6VxHqqxhCFD+HA9MwbOmoepEzjSpindOzjZYYkg3iOGgS/gYYUK90JJzAglunvTLWl
qzDssGXZ7K8PTcopJQuayXleg5FHbM+kGvNqlLRL+F2UeCw8JzUiWWKwt2UGin9ltsu8lp5vfPRz
T7d/AoD5DjzYROWUwVANt/bhlpZ8+msIjq0ANVyV/eddAL0/WBQBLGVsRa7j3bVqClyVr9P2EKhz
SdRCBRexI5uz4vbb0UZzU98f+zeYnYHsWjH5v40OhRme6no0SEO/PPXhKIq1nzztiqRGM3+7i3R4
MnWlzISD2z3TiuVcZon1qBdlUFOEFiseZ2+jYq4Nr5FzPmVXz7lm/Jtj3NgE0mgX/xPJvRIcdtkV
1IhliuW6s7JroIdZ2uJF0DfYcYAfosgoCfNH254GXSX+kaOkSs32GXBIznLqdnNx/66ktFOT5jIw
5OtkklMVqkQ8Du0NEhD5EuZpl2eZ5F0bmXgkg92A0gvSTSbYOM3UbcKT2oxbPqr26f9d1Vn8ChTC
N2JqzBxHPNbr49V5MGzEygG37iSnzNdGHthhKKbHxGT3vD+l/F7boQMeXPPmlXuPZ8fg4FLNMQBE
+f8j1bfZnH+xyvd9ofhyBcK+Rx6PWNmIbKgt3Uof1954v5PyAkyiCt8PCutmbTRCQKxC93SEvbgo
0ICUpXSwekfEzsaBGPqq/Trt0CRLXeqj5/zoJ9dGPWv26s5KZYsB8DtdHKnY1v52+TOPqtcInsgY
sGQh7scoXScEZmlmnjlox/4HCx9S7u6flxkOfQGnIHVPWekU53A5+A1a9vkQ2w+TicKT0/3ggT6Y
vpSTAtlm7GHjG5myl1QVcokfiB67uanuLex7d0regYTfJTl9P78ijhygWa4lKELTuBK+ahINVgDw
3TPdQC7OZ98PNtoBSg3BUWGrTgshCZTYhUjMMVM2r2luXfIfHRTTrsOmWMt0BJN4fDUomiwrxzmZ
XDBXBWb/k1oKpWrZQG84BIqXDUTGdge6svEvbd2Y513R1u5CLBLFJzUkioZZg1GhX15yDqdPBnRN
+YulpdG2STLCd1SvSL4QXL3tAYcGAUnGEr8VWuFALPPT+vCBvxbOmHpRzD9w+oLzrLHLxXYT9A0k
NgSkZML7/wYscWQKTpd0ogg770ZDHARxd/hCn3zlkyhKvD7kaXQvh9tair5R2SyjspAUScHQwofA
rz13Qotu4kXU37fuDba7t83Tyw7XiYq36wrkYTnyMKPiOr9hzEFxfknVOAVXVFW5dPkXOmabpy0G
SGuiTYnRv54QUqGXzmwOXf7momSMshYVwpr6Up9AWg3Jbw5COYhbJd0673rhp1J8jS0PN1ESEUbF
B/pQjkkYQ3ypca4LmkMFXiLWGM5SRHMvFuDA/tr6mxRgyYPTukwFc89RxzKGdU/a8j5cSqf37ZMT
Zw8U80C7ybN+SSkU5gfp77Q9CDzKv0OCjWiQ1NAwp3nYB2KnjK0baonrup/7PS+LRPupDEAf4s4r
kPbDcJbEn7ZkQoMsiCql4Vo5A2feXcZCpYufIaKeOHA+YYMbmrXoLo40zDn2ilhV9sX/bPpBY9l2
i+ORIvSZoCMhYvkvXkHAzWRcn5EBSVw+u51plFdlSPf5asex3nrUBH7Fgqb9g7go3z9SbrBrblZC
XGKk+52/+2LWBNpDaoAlYIikN8dmEJBP22ykDjxWpMm6xOzpABKmlINTQrRoYTJG60SJQBPLP2pU
+CpFTTtCXMKsit6ffD4PNggz2Xewl/anz5KF4zS7xLNQKvAuWTrJEolmTlXeVhf1GmQ+ItY5ozSS
oO80wo26TekvD4vsiFWNxoaRiYBqv+xCimfMigUdQRsq9ocLXd2Rf1f5yyMLQC3nvs/3zmUy0tA7
DHxQ0wuvgcJ0JItD5+826ypWmyFFY7a7Q+lw0Xg021GaAEqqR7c+SdNQ4610vQXTSZMu+vyQhHh8
eOk2SGY5zwfsLJYd5/GTdDgOdkm6Na9qEWkANp4mHWRZrxdT8tbPSi1ngvwUWX1adAtjaGYwtKcW
Ac2L0Wu0FLhHLTrwh6uaH6w/duZlPRlZEOPfe61jUcUszyYvW+3sluVL7L76SZzwksjQjhQAB90l
QdMYXMcAlBBWAzirzTPAg1lcW2W9qavTymuZ/T+N51l5h0wYM2KFYZirTRRsMdIEQF1Foaom6aSs
JrGzcIPi73Onxd/Pg/NNt1ObqZNmFQUEytGM58k+S5UD4rqC8IC20Ed9+THOi1Sgm3+dR4xyXJRe
nkh8kPUzKhsYU+bBbe0EFQrPe4WxDFXtKgr0gyfrnHpXvApCit85iTruu8xInfXEVHiCVuZ3S2Hg
EiSYy0YRBNRnCWhR+gerQbmyI6sUuYBGs8mI8jofvaWHewsPuLggndjjwu5J3QCTRBBliK14N+JT
9Namh6lLRv2jiVyT+2DUpa6O27fdDQFCh3cmfENvn8rEC1SybkTRw//xcLprRoRR2oxu75q5k+YE
1LFwudHIwHFWIZtUvOfuKaJudD4qMOjWpPlVOI5wrPLUC/NiQxxYxGbRP5W8R47PZbYUkNFlE9RN
5vdUEbHnskOxMhZMIeLvoL58laM9NAGdJFsKVLs1tpFBNEIcKKnr/bGyt6XC6yk9avFH9AlKA56+
ZtCghfQ3L1RMwihYE7w8+4EXVzvnCXCAe7EH0AP0CuX6a6KBGpUynlhO8UqnFGjLFp0p3I8lEcRv
J0rtOrKqQ6cjp9c+BMWrq0GbCAlBWb41kV0gP44lyPAM5TU0O1Ht6l36h7itpxPkqGHP7in3rjI6
zWFC5mDO3DiE2lCUzQEsok18zvjvOmXrP3Sj2k/TmzHIblC7v3Yq7aFSjcyPjNsxmsiIWFljrxnw
/osPse+uTPRTnWe1sltThISMR+r1v/yG8M9MhAmd35E0lSFHEuiNx3zkCqU4rWpoBA47LhPcuRv/
eFfWrKyIBPTJarCfAsMaIr+LrRS33yh+K6I21IOz44kERB9MGX9N5u5J8RaAw6e4TFqWO5uHtTls
7nmICuwycl/ug8g+vMAHSkYBruc0ke+ucECfJy3T3IQA0nfvEJh7Wzo4I6eZ+Kh2IDK8vTC17rSR
8N/iE37sgOLQ52spSvPT0ww3zmRM5NIigH4uxDrEnEM1DK5essyVnQzhvKsBnO7iKhT9Xla5cN3E
b1POU8lfNk24gJ1nLKfTtQ2cfU6ZOP6DxBHixKiCx3kpjOy6ECgK5uzzvksYG36dQTV0i7FJ+Y6Z
Yq47hxQTAl8lTd8CE1NaiMitBpvcFH/6AyXexAGQKGBirnKGf6kWoA5m9Nsy3dprnsEr63FhldkA
aitAFbqsAGGfKoehTHQZ0ZrqzfXFtIiME4sFiPKKyBrFc2T0v+wtljhEVeDdvu/Ak5lH5ECXskSw
W3RiQnT1oldmDaN7z3jkdqHWyVba+vNHQCO8btBLx+yPcvq8jzbt5sgwBdTcA4LfCJHkddESu2wD
cxb3n2AZ3LsFUwTSO4XelIg9l40Qos5qy+ZWmq/Zd3xtNFIfkrmbt9vRTbrSsWxmwRNx/j5Rxc9J
6FbrmCGAjk8H/H3i19v/rhh3PGFvs3uGSwWhzKa8HEZap9EwoLoERTod5ZnW9NyerhOjdwr5zex6
rFCSsh0pidtudR+AdJgYA5iHPul7tz1rt7KfKHUoHoX641Sq09zLg4F0L2V14dfQghL982kcK4O0
NM9WuSLtn+3L9t1HKTiUH8RuWFUItQ4UvE394KcWpGRUUjFoNTWorcMtLXNGCfpWL7WqyCcPOAtO
7JPJ7cYxZAqTo9feoqg84yU5uK88pEkaX85NjwOWu4a/SWShx2jH5lNpj/KFaa+gUD7sZiQfkBCt
wBXMENv7s6o4CnwwE65bzRXDbvZwtU/3+Xu94tqSz/fYIi+yh4PAgPMd46E3vZGkI7PMKjzbWncX
IQLKcD+MWUCqvKzznhLvZNguauho+Gkx4pz+ef/95Qkh1Zl/kNRLe5e0PFRHT2gRKXIGTkxwDLVm
n6EUCGIzPGWNW5hxo4qbU/ngEs8rarFmr0phm9FXDDl76YyFhtD+SdK0kvjxOp9tKfepxdeT5Jq6
g+HEAZtdMDR4pD27FIv/V7gBlRu2AMCEvrL2Cse7gtVqVJrRGSAq7fBFw1n7Q0UqnRHDidldPJUn
fBdXlA8gcMhbKV33IAx7Lg0NghvpOKTCaVAUHa5Mo7/5o74S9WsNy0vLzXWSV9nv47M0UudIcWbY
hnpPC7PDSDuJ0huHCKaS9zpQRV08vOglpB0B6Kbr0D4HRVMHRcIWvSlQJyZEFWDh1c4NkL2u7L/2
9RnwgjBGbv4RHLrLAyLo56MB5TmRc3cLWXH3kGiZCzMqaMimV9lLjE6jtHSkzXNckdgGWxVpNepr
FMfVeLdyFo9weA/oBNtofJuugn1wPYnsvngmFxV0eNHpSQXzU6FSdUbqXSVZZuqiwTt/cWd6mDoV
hehXKP25h2BHJFMYca4iU3WKPnZ7vwa/yEml1n1XYl88DzbjoJXsGbPPUweuVs4evhC3k3C/AChw
F+sFbZH/8OZiowrjRhbrvnv/id/qJjSaMLxnOv8p/WT2HpECciAW2Bd+TdR6wXustcoGWYw5Hjjk
mV+jQBci6uuP4LvKg11P7+CTwvomnMsRtP2XCwrN/1SSXFkeglifEcqw4e+JI7AuCQdLzf6d84u6
dZHE6dGd4FpFbQI4GAAviM2TgQqYQpAvSW384xICmBFdMhCGkBPIFCWzyKedC/fSVN39YABwRoDY
hdApJEN+BkQzLA7fgqXLXOB9REMFK8bRxsJuYC9gfsWuMgMi+aNjURXYMhNKeSgADi6jQiQnvp2D
QgUI6+Cdj6eqP68Ek/6b+K1Zrre1dXv/ePbEo1llKzNDrwS1dnR+liwQ7yc4c/7ykm6uakngE94p
an6lujBuP/PDE+vQim8oZWc/fOJ24P0cBUjfAieFKbT1Htqv+6Zf9EMO/GX01m+TB1fPHmiC7aDh
Ywe3w1cF9eCH7TUaIwCkc933OInveEEIRKxRME/D/2oHqtLyOXwoO4xAknek9DYmvyJUuXlh1RlH
62sRJd0/14qFmY8EvOjMNo+JlHK1891nly+bU5XqP1SEJ857PzARJ2giSddjeOOcK9HlQ5GSaJFF
n+8d/oeSzp6cWjtkwxyZ9FhBQnSIJ8fE5R90NVX5LNWzEcddEOYa8GqLluN/AYYuE2qgp88R5JQH
hJPew5YZ6ZjO0JJxJsK23VM9AwJNZqjtfeHdYZ9zDhjftXrhwm/4r0VVwDrQvenw651kORkejM2n
EescIDBOU6DVGbqSfeaqYF8rX+XRvFGWZL9dDsrCcPwkenOuf4/QmKt1I8EUMVP9HUmC9d/CTC8e
QuJpIoSHS2/0KtBZG5vAzgQ3Opdt2FsJB37ZwlnTc/rS0z9Mqpc+esWUKIWb4GNxe7+1o1mQLcrz
QZ0BqkIzCk06ybExXOpTa/53KW7gIX/oWmivb1ugMmD26l/oCPjZQDrjWkkiMKELgToczFwbUbHX
csrLyhqzNKdbhs3Acj94S03b6RXfl8mxptQk9/1eA/gVmTGfhLXlcKUJF4nEIteYjOcxhwsWhR3y
APHLxnfu2YqN/HHJv28Ut2bgNE/S9w6D9MRwaMuDHittpg9T0aEsz6w4pogbtWwIRaN+Q41v7XGS
55798M0Zt27LpiOwIwDTiKeR1goeWCLvnpF7jW2gA/jocPw94VRwLE/zzuqZbLCPvN+8SiXDM8r9
BZxmypOxOoD9Nl/fg8W56scFBVLONY46/YzoNA8CEi5Q5JNDKS0R6eO6XUTIJM5nWF2fRO/kmmB6
syCqpjpL7qqcsMt12mfdPuvPTd6XSBWiC+sDTOUdIf/wPvf/vVymUj/h+tr9gxkl7+VL0hBklptw
6evyJZAGsYQcAuOB9jvMM27uOqMKGNyy1xM2IjHTuXdB3gbcvEYdj4PBCUrS4PBJ9fmIRJNWaOoe
fenNyI9prlVsyGKk/j+25Pr+5jqdOdL1G0Cdg7j4nwMzObzvjwngYd184PlJa2PEUfkpi4SF2KEr
RuCJ4oCpqzO475Qv/CcSl4ve60tEPw8NFb5bR3qY/qF2X3672IoJu10VR1UebSrdoKbZZZ5D2tzY
xZp45wwE6gRgvrJXTTyj766hMAi5mjIZ8EUsmMQ8c2JtdutVAqZP1ilEbCD1P9fCLmzhgA7GFLPf
FHwoICHG9hI9TVFJCgI1f0pYouiVugwW9d+v07Y0G20e51HpOIlKJw6lOnnlketlk+ZC64+KYfeq
QH7E2tnKYLPgT+vguijoF1F7PVPgjDg8Pyg16/fyPsHoPoi39K5m1pTZZ2fLlk8r83j+82uwzayb
FYsCiqnjkuErW+RFZ/HaZEB7+yQs50+BJB4dWREX7FYHwzqfYe727yV4kGD6PkpZvg3OLK6gPxPa
UmZCQ51OpazoivCHsAdvfR7BZXlLS8sv5/DR7c7HMGSdvST/J9GSPUMahV3yCWlhHckNNd40XZsI
f4c5XytErHKcGsZfe00b7Yqdgz0j9fZmoydAUaWzuVM/rZKuBeGEaqAtGRE0gfFkmyq2cMEN3F01
TG4LtVF/A9vtB+L95KIQs7WYgGbPt0y9xpbR1ZjE0Eq+qdbhQsNip35lO6x64UsffprVbWwlwaXQ
uffQ35VPM8FngFvoMSmpjBEWCLB4J9cOuThKmRUjSMI7/SX4pXVHUsjsZS/eK1E5suDfWLaSSO/f
aKLS352qnih9f/Nt6jNCCvSmyLiYiKACGlDmikbR+l6m5Ly1GMS9CZgWyWYpGg7nEvmhrVPUpSTx
TJOlRzOhP59DeaPSzSSwptqqIFoGmom1eWmKFUy3mxEHcPv7K2lRwMw+19lNw6FUdizTwvTBLAms
enWLmF3qu0JcRPTu9LtgMRvDetvcX3dWNlQt5dNeDc9O+lpQRKnQPXPTu9x52MEH5DgFf+DTzfdZ
HIN1zhJKA2ORLi+rIxg+XChDq6OYRAO8TTXLvs+fn4yMdwVdTFGH3hh74U9B3AIRSNYWhc9eLQMW
mB23Ub6p7Cfqi9nsvc6RrjyCGsXIDId0KVvzqBwHTM1hgxk+HZH4J3J4Gqw+fI6q+Nyx+1cKUn1b
cJ0qABKCqToQXWJyd9PmKc44Uo8bD4u51NXs0RYT7/7pQv7XAtZVSsCoqL7bN5pTgrbkgofEt1JC
Sixg/m+HNGfuPulVprHvWcMpkV5fBxBOeSC94rJGGebtqJ0uIP8t2Eifk09uA8WiEliuJ3KBOE/+
Xv9nWYxbVFzwirDCRKNsPycK+NQkZFGMFEPtP/XpsjmkrtvcAPKrUdyIAj3fsMqcCbQACqknsO6v
igiGsnEFm7yUvR6CE+IEofQORkfzB3NxMNJoz9AOjfh7pX61Y/g/7zjKZvuk0244hhDm93y9n295
PgMGaCcKNg+7Aa94ouPP844yRa8a9KRpKzUH/CB38xM6mArGCsSSZHD5gVRVSMtlW4rwxdT5x91L
OpVeMh6OxxmundHLzkmndtE/4g2OlRkAcd1cgiQsPXIsKLA2ZyqiJDIQC0fS0g2ITmZgqzF8nqgB
rxuHE/HWxoEYIGpdFpMYAcIFYFuVBZiOsXktDntzln9QK/dYd5xCXQQDRXWy5mga6AC4y/s3Pb/y
gKdiOqrExRin/9/OMmE6G7rgnF6EI88nss8+2NJcVX6aPVPmvb5VJ8Op4lbaaX0taNNQTT1QDXLa
qo55b9Nka5c376BlMLdyLKXdYDy+rCq80iqeZKf24LudfemJND9b1EFZgbQAMJrczig7rKsx6LzY
wuWt+vx8Sk0UpY+dQG9U7qrSPe3CCSPLfyKss+MdcN5i/qUcAQokBtbL/LBKstm9/E1I5/0N+Bvk
QSl/XHofPtENcN7iSb1fgs8RarecKOAS086mw1ebO/nLKyIvcxEzDmJFGtyXIBrlUim3nxlvp5kq
uk1vB2p6V5o3PjbNP9BFHzozPfLg4Lq1J10lqLPFkiHVVk3rzKuxMnQmJHIM1tUnXNG51DfgxHU6
yGNEwmFJCco5pOJtJa3AWaKsKv94Rt5vxxaxSJIoPiwxvFXhYkdB2IRgw6UcwBpjGLyVUZmXlmKH
jO7ZuTTMqqpm60gMycTYUGmrFqx6sgZLzygjgDaT4j+rLareA1+D3QcN2FLLI15+34omBLV/K/Ut
dxqwMr16d3yIWBuBikLb+nE8/lb/1DWY/L+gnchzIFB2KocuiWMrfKS+BG7RQ52gU07RB+hew6vb
PJFs8BhfLVZpqcST5nYl3ScGyCTeTiEFk4xrnPqcFy5MEaCZ8uKO+80YTEFdPT/1DinjWkFFWJXm
s8FFSOfpt0EzstfSm4BlQJsarqTrOhQu1JT4SVNDZd0mZYGk3Ftu7CJRsKveYajEkAOD4v4D+3VG
Oi7d0mDRjgU01A1XQxxCRD8n6qSQ3jIuQ1xBRCx485udNE/a87YNjpqrlssd3gBMMNf/N3EN/wDF
uNewlAQtHyHM/hz87IN2qV3Uy8qDOcepjb6snoDQ5MJv6guGr8zv9RxSPNrKoOKFP4ww4n9rOEbV
uGw7QaQ5aHL/Oa3k1KUkGk+3FFyAxb2IKuULCF3SwaLNCj6V6FI2DmFtkKHSzS/HmXaE4qFYiYoK
4WjOumCIPgZohh7TVRZ8VoOSIzY/C2j7CqoCz5NRKc+5l7QAD4UWnK/yhByYA+bmeUodogQhrdep
6k07TfiWX360ycBDgvr4G8eAt2F59gdbUJQcXD/WyrfVnJCnTgx+o1PnLNydeA7WzwO85p/q5SV3
gbABbJf0TGrXPsilfampTGJrrkraNnKukkTvL9inyr8E7X3fnBkBS7N4XRRc9BtDC/aFgbKS4fy4
76w/L/d2ZO+/i/UBJUPzuNHmayzU/otmcWeZjgAT0ZHvXONYgmqxTh4bH3jZBw64ZJikGFO4cTjf
UzvXuoc4GdYjLTsSa65sNG+78u/4cXWoI3pWYdtT6+UOJKGfCOSUFGN/v9SvKUs27Z/Q7J1Pve6n
J5RQqvYuLu4QE+iLl453ZQGQdhKdRsKlqndTOjgYOP3fY75YFrt+8Ku/PnyRHlfbEuvf6iRpQAVg
zCVTjj4PxSl90si1aRP3czdF7pvcTJAu5d+iwutVEo7gvp6Dx/86grVHguctxQiy77mjk+IM+FKz
AE7+/CHdezm2PU/gwzTxTVX5FswFm+9Ivo5a39wEXsSUNUoeveTo09weQFiH3Z+XEpXtefTXoWSY
xFHWfKD2GCC102VLUcBDXJhvglP/5AsIeY4dZzt5Dg5TkAtkItxRM/4PFRQ1/Ydys+ZZHA9K22Hj
EDzUR00Z+7LeB3sKcXtiPWan29A3q6OESNlzRcg8kwzy4OoCVzlRcWG++1tspJsiht7Dh+/lbR8v
JvgbwTlv5lmK+4g3pG8CGF1CAw51iWI/DZin4am8gSZQ5pnTd5HPJigMLwdxNbzSBPOupgT4Xcxc
u67gEPCOB1q6qvSR6kI2Yab/l/oGv5qAtoXWE+tluoRtxGDipBNfp0S4BjONLMieZry39a7MACsy
Zwm4JexfCuH17dytqvkvUBgD6UYlbaBjbCUAiiOXRbRYxSo3cZvnPbdvAdgPQmamiIM3okg5LsJl
Droj9HIJrhC4RYy+ziYDPXVy/xdRVCbYAp37HPsIL411CeGF39jS5xHGJfi5xFtS3Hbm0hrkWJ5L
VFV/N18kBnYrtBWCY9bhZiCdkB38Va388QuevayjdI7svHvdbhvg2xmDAMePDEqzbqvvjI5BW6dN
1N6ZcOL5lBsM9Caz1P8sNQkfDFNi+8U0G+ahWdhdZHzaNMpAas3QctY9Tp+9WjVOpG1RgRquxqAp
kXC3WsVmC1ffS3CMQdygEsnJLyas0Sk5mgqZHaO9FBfxwQYLHtNvpW91O6j1+ptdMU52ZE8CWt00
F1aISD7aFMkNrW/o8KIV+clZNIJMytHbhMFH2pYBG1ZnsiynNJaMYz/Wbnjgs1Q5E6hfj6W7Zw31
sr95ny9pmnxEd1j6ilTTqU454xhEIBza2bieTUEwKGGO3uQGki3CwasxZ9Pgnj2DV8TQF/nyCUFb
BDeoPf+KhPyk3pZqxCvh+beoEhYbltaFOGWIH2/JxJy/v3OQWRPoXvruf+mPRLLDstjlDY8tLxht
wluI+fRlFHttu9f+DWRNN/DHCztdV0+zHcUIJD1n9AdKaC5CnAf0d5NLNoiZiPCgDR+Jo0awoKBm
bpRHtwQEtzop9v2GbSreJIj1N8g4c3MGy9oGJ7iGtOupjiw9Jv02BooUfD1RUbSTcgAruLLJ8QEP
3jBvkE1ejvQ6wFkR4DYXrYQ5BNFgy6WBbdEFgS1lSekXRbRR2U2hj/2YjFZdqelCVee0OT4IDw+r
6QTEI/HSvx8ul3npNpr9j6g67JFK+9qKKMfYq+pDW+qfNu1EEiakpCJ+0+TGTPFo30alGaR1+xr2
zbC6NiiJOQbvqGxJbOBoHONhVbtiXrnv995xhL/H2Mq91vKnVg6i62iLfbFdWcPD0vsW52Xggyqw
6YuvKl6UdGUMQYpIMSxO2YYy/OrbOs1uC3ndsdK1f/2+yxfsa+93c+OUMP2v2qGKEFwGtbhFtRkw
iS3l4pdgD6XD1i5s64Wpow6yXuTc3+4Mzuh81aUJeQLDdTDGFvsQxpBAtlIJ7U2V2YZouPidMfG2
Ncru7bQXmy5FKCK3rFojer4C/mPdD3B0dvuCalMD/5kA7Y0igOe/iTE5cMqra0Rzk9gBoOMOv718
ZwI+Tu49/3Mi/FSELI+R2jzlO534EOZXCp4Nn9qDhdRoAuXu7k+GIHCU4FE4PndbIBgO50y0Bh19
kgv4/KGwBoK37D4eanKFasRujx1kln8dBRzAmIR1sujianP732wrnwJnosCuEiuaIO03942BIRTq
Z8Ovd+cflvP1WG68B52imCdLT/Fl76YWRnAZUksDOG5jv8wxg1aVIDTPobrLdOU2kdRwGyvRzOKO
xvL/UPeDipHXqxB962oH+pPslcU99PcLPtdQKgJw625lGt6+c3cKuppzu0U0GviY4Av/bxlYxZHf
29fWGLyFMlfOPtJLAE1kkJVwGeqEMbhv4qCuBHp86g+lGL8Qq0KWyEL6C+JGvrsYoopmT8deDIof
3shbOzt6V4QLh2mbjYi+7WOjXRE+brK/fufEPnajico3YPMtdr01x8uTa+7otqOL6o22qH/siVPI
miZKVqdccYyN177BvD/iwIVHeyxGr+3EDHMBjFhfsRDPGfyLaZzgZievzYD5m2Al5TlOsRW7EECr
+4Gr/daXbv6qhX2RJqs/QucEq8S0DPypJeaD1sGT5Axjso1XgqojeKBI88fQaRNBqgOzk8wRyPFC
7G0ARTa3izFNv4SLk7nz/AbCD/nDfzRERkOn9ciR9JgDYcsNF2NJk4QG4MjPMtzn7T5MUxug+ITi
M5DCs4hK0QQ6T7rp9B/79ylSSQ1w+itYgmkK5N6M4Wce9/t2r9JuWrDaMpJXrBfnEww5RF/5wvro
xNEqC9Oh9HKlCF6/MVtgG8Jff6s74bSe2KMIoQZHGNymHKqAHs2nckR7wiH5dNg1gL0JNKFq5f9D
1WPI9RBb238g93lSUj5LlcVhtBPHNvf2H6t2U1XZ3kc9MXCkLJc9tG3sZ/LafEWR0G8nRP6YXrYa
rIiwSNO0R/iUTZ8WDPVGBrRD3cq0dEP81cty5RhzeoKyU7MxMvxoo1dFAqpRax7w031A0jfvXetT
BwEmDdUPdrxfuecEskrVHtE6NkA+sVACKYb+J4ogMrkxIl5qZq7OEpvXUaOeyV/pEgecdBmP6ahX
PK1Fz6BRoaghWyqIUKPbzKsJTNLrEZ/zBV4kS6opcDsf6k+Alc9aJhdSXHiiZBVfTYwVMd/ALMya
M10uR3RVQixQzDD6lu7wdCwyGMA/5BZCafmXPCNosQobX1Wc4URoerxA6m9AsLhguLCgSqfrPP+Z
W6KZeeGcFQHBW5rFOQzfZkbpn4RDMOJzrYMqeNm3DN84R0eoKDG52bVNxiJInPDc7tDiAJ04TOgZ
8oqDU+Rrbft7NFQ2xumAhvCT44R6DaLDBC0aCufohb6DUP4qj7j8zfqP09tGygL2H37p9rFbLUb0
C9xqRsEudtx1BizlbFNmS7wC8AS98dtwJKtyNoZ1CBeL6UmBnWJp69PmkutYXmRdaP8ybEsijD/3
sQUyQ8VjAcoQcgITyNlfWPLXzd1xa/gIH/wWDDYVcQl4AKy6woqrZEskONePU5ksiVIBilCYb7BY
Z7E4liVA5xqO0ZUB0NoQgJKh3PVVCD0b0cPuoobn6xRAFbPrC0gjeuyPGVGR5Ss1f0cXkmk98mIf
a/c+vIgsLDMgo4RLUnuo0+sd/lYQNWKm2q+MFCKGdNxTzNeUWLMdhG6Q6w7X2nWc6CglxvhURK0m
0xLZcApxd/g8CXWEP9bPEDraZX2AgOgJYxojO6y/TSIpvREwTuEZtlBOtyM4ixTCQWlq7kKrcP29
TTGeEdlW6ylL52yC2E5hEFVckF0ZKuD7kjELFIE0HM/NnAU7cWQ3+GrmVCjNIG8VXp/ZbMyGzvDU
K6DgROpa9mlt3jCWZQFSPzh/yBXRZVM8U3kjnpTYyVtZNMqBGHxHY2SydYqExKo2g49j9tALu7D/
+11kezkE/EjdyWrIBi6w3jXfsqof9TtBCsx1VFNyfH76W7+s/f5RtH6hd8Hog5JbFUzIDYP3Waue
hhvhnC2SpVEZ321c0OvdnTOX6CESgch/T6UGfwgTeMUC4p/rZYxU4SHptghQ+8u9QO6/yzQE41Ue
aBNoU2AGc1ICNDAhkucRb2WcdoaliCP9dlwjGeF/aaLV/uMLx62ZMhI8CVH229yQo9iDnLRZZClw
6MFwSbtzPS3STYGArr4o+Zhr7P7JHU7uMFK2EoegYXIZHgQdvRGoNHo06xSuiF2hnrZhZr1kVPaU
nNfDJM76895YeF8AG861SQsm9G52bdbw5W+W+pDczGcf5wymE5MubFFHt4X0SqNmAquOfvMypbgU
yN0mxkvUG3QGb6EDt+og4Oy08885pm+wn+xu963ZH3W7fm+aR6NU/r6ltP9YE4aios4/nJbQD1eS
cgMy3+5mByJGYTP85rXB+jotN9WnwHH09lzqch8a0WfzMu6by9/YW+6ihV8gHuTyoxBePrpcr8dl
WwiwduhEPH0xcVTC+MRmemHf9DXPohmelxpAw9zTS5/tMStpdtFzqu87SN8hTRL3LMVAaC90YBou
LCMneqzk1yJlHeAndhFMHyR0wQbeR+Gy13YGYcI2u2lZdqF7IJXCG00D8HNzfLJb1Qh9xkRVpRPB
qNYkKGppWNNqxhKxkJkQpHr7X66Bid0Fyg/u2TKRiboNGHS0BkpWTChxaJP1wGoT+yj7/AncLELn
yo9+W3LYqWRnMVf+6TRg6paYDSSRqQHpss/OBx0UFSwTCR1tfJ5pmIEdf2jtJGZinQEVq0FB4ksW
oCZuB/42iTj9EaWjigNuY7BpqjX6e+Ov3HdtMO+cMg3QOwPcpNSSzDEUiSSgwnMnlf+3Pho3YJkx
MzqPuyucefOgRoxQ8MNX+kJfss5fW3PFottvIV9l4KKK9FesVUZ9oOzfZxetaB0LGEF4mi8v2Maq
mO/Yz3l9Np2o++3RBJtAkIlOqXNEsnfyJ2iLxEOE1dGozpPY1fl93sDe1aEj9SF35Tg60TX8s1PH
5MJ+6PKIgPN2+RujTmq5IpeIJ85Bnwl3N1d1XbwfjM9Yq8q0NDZpiNXaq4K2vEddQd+32kjuQ3hG
HINh2qJini8SlF2spwWgKp+iMGthK5QpHj2M064GOF3Bts30PJqhDm0/GPSCcoMVx/swxYG+MaZx
WLIAvmaRBbX+XkQhpx0UiLsNwMnfTzpnB+8WNu8QDWrYSGRwvSc3QpFCW1DPWWFNTK+1JDYRVn5H
dKyT9n+xYggt0CfTNYgSCVhebebiJZFRzhCkbFL7DS/xnKmCITZd3sIAIBMGHjzG7WHQZS5uKbZL
7A0Uo9w4EgDnJugV0Buvhp2DgLHNaC0HrdfQH67xHHbbje6p7q5O6VlskHI0qczG4jAY77GLBf8h
mF8RwYBYbzTzIOzcheI7z+vtJTuXeh2HIcCUBZLuqxiFk7YvZqMKAfwLUEHAFDyZ9cnshgdUgm/q
enUQSZref8xlecPTUtwR4UVFv/joIJ49VDcyLUTm1nGLW6JilG4FxDHdphokPp/Dq6Tq/xAPp16f
8x4Hc+ZP69ihtD4/ZzDpkb9J2tpvPPWJqGMX3Hs3l7rHgYDMcJyXBAVCdpkjLfkxLyqE2SUU6g9F
nOWIC7GOBvVEUJX2fMv3i78XTPtVQtTVKvpfXXjukpyKFtt8HQyKvEuQ/7FYnA4n2aiUh8mUR2Q+
I+nGzXLEX50Gx7lW8mL2+uDm3PnpoXu8sNRcsRw48hhUq9SNdVy5XomYwgoObaqxWfBO5lxRaY7s
ZUMGbvURZRfcqjSnmgs44oz5nRRrZcuJm0pXlCBvjDgsZf8Ai/YQa+E7UymLo4bZEI/uu6fy0rrJ
EucZUU9Gh2XwbZ9UJ7i4cPEB/XodsJane5YGCuCTuUuHQWI/0D++Vz4aiTCnK0n9CI8n7KXtu2PA
pO4/82+xEkmUVQEFtsUIJ6OXFq7YnAjU65GhIRquvYwvy7A4DIfi8yDcF9pCGIJZD4nNVmBhkwfC
rTWdqUuSzwsg9OWVOUd9zBTyMdfrp0fZzH15if4HLY3g4BQ+HtbcH2oW9bR7LJvg0LdYDqqEtIrc
kxeJj84xoGtTBrQkS901aBcJncdQM3UU6GM91wUGBjp2s6lbr8+DL1ff43U6LXCMlE44WP5HRIJF
ny8ICQDVpGxMlH+q9+57GV9tk+Tfr4CZ53S+1nY11hq6rZJAOdh4MkuKJdg08R5NVF1uFOUR37nS
0lUYuf86UehXRXO3EAoPZTghnhhkPhF5gt1ts+wl0uOm0W9EyzdZe6sFvW26RKF+a7G+7F57tSeZ
vnn4YZirq3A7bJz36hDfNjcgvDMYH1E1LMy0mz1dp8DhA9x5j5zBM6NVck7AdIWxxSovZ/DG//1r
XCjh367ivX8gVlGRyzKWUyjLDltUYSfb72h5bVtTepnhf+bgQLEx4VzHMhr0A760TeguX2LT1gXQ
KWp1p1ObXgLkiE8TRB2hDstCnNpkivQWR5eZqSBacuuoBBStQyQboVdhuiXYdeK2bEeobbqghkxe
jB4catA5qLfNPgkJr3m3NRa2QHsVh2m2DwzuoqNJY7ifzHdmoQOZS2YZ+/IEodZyJkl4sh1L1HNX
oU15r99R2eewVYCKMf9Z0DSjS6FFjAps2juM+g+FJowTsEk9BpEhaUBHoJ5+dRNYecyykq9GICGm
2voALxcd9KZsiYBiBEDSDxxWNKtsckpjCS4j2Ttz+RakEw0PaEWx9bdu+m9M9fBb0vx1TjLaJthm
dw/qmoeryhxc4vrXOrb2VYfD89n+R/ssCRKVlxs8tqxWplgyewqUMVJlgT9rkhZ5Pd+/Riq3yz0q
qbwy46uj0xvxmKQ8du1leoTuLWLBRXVWbmYxXOzCLqgZh1Rcjwc7QiF+x/qPBZ4NG+cURFL/tsMf
J5OEKK97V/0lk2U0yWz9st6YAG0wo+Jlppr3oscihualkEoO2wCRNqA1d5UPRGc/Jlo+W9nTpNpM
riNDnHLjmOQy9CfupfiEsX2eJDiOo0a+Jt+2RADyqXn2bIq/jwoIeJ1f8RpoNmEnVA2dZRDMqKPt
4KaoQ1WnAuXkVTz/GY2MQeVl+LitSJvXxc7b4Yq4XbC5SVWVQfKoKm8Mu9y1KiRQVG2WHhhyHWjw
npR5ThlCZyVZSCTUl92xFrFJIHnLoLx1iRARLmuhBknVM4aivM1ox9UvcFuBJBZIaEOyod33Fycg
Ru/g0d+7vLru36SGEh14Pt6Zfw0v1lLlNsSk09zgqu53XT6ouvUb5T1gKRBTSG+cJdTXK0E64NMX
9bapeDA+uw07ETxPhEC10wCO9YTmmRLm6GC95zjkp/HQ5CyAlKLIUQs2TBZHYs56eWg3qFH/j/E1
HQqR660a4YZDzgWH9iC/3/QmFHz+YcbeUR/fmfNXx3e1qoLkO1xdePe9TzbpnnJs6p3nA76n1lzl
DNgRT2Un5z6GbGBLUvY+pfqzJJLEzNzu1GE9MPXq0Kh24W1V3QNRJ11k0HtduiBxZZh9I87AqZkF
v38V6oXMwJLd2fFCrVaaRdSIH3yNIc1kM0giLepJ9l1fxXVR/FjYZnpvc5LjXldwQRnZiVm6EKo4
AacF+nF1FKJORBZYphn8UmQSEEPd15bH6GhSfF0BCjesfxyxNYDR2uBPEotivchqZtJ2Z1/Qi0JR
LAY5Uxi2uiPLtXiIXo1+7SgupxhG6lcSAwFCVVqnNhDWXeZH9QZs3GmcYdQ/72+/wnkZyZTuiZiz
6CCX+2czgV78XUXzPQaj4srdDZHQA3tCGv36tWjW3hrm7Wliek8dD/XaNJuetbbUViWjyrz6HMxB
D7oaiH8LSWDn7hg25bdMYHZxdeqBjcxhasrcynebRIGVgKQh2oq1BaZs2Xo6wz9JC2dS4d1gMdCP
+DIBIzTbf7Cedgs9AgiHyEh95fuQ0wSnIZh+SnzTdwNHGqAUl0HCdIvqv15fQawAGfiJXUS0TLIh
0IeIfwX4FNgtvtM8MKFWGHkdjVvZZXU2a5Ffz2wSzRnGFLbjV4qZNJ+wy2ujhXKR1RQuRLWfuoyR
Lyhp514af/EVUYX6UyOlgozrStuMgO2NvSRcHT9IEr57WaKftu8C3nRDpvacOfTgYAn4FlyYay9a
oDWJvhNQhZYu4aWf/O7Ys2gp77YSn+OslElMaBDZyECBMA0p7JsuIpEZ1IVAqHgjkvKLu0PkIMnq
s6ewv7ZjIKeiCWP1pn7cchEAHirHLkGXZMhPEJxQXIt2/xKN3hJv8teMIjK3uiEpRTn9d4RnCOgZ
oxkDdiaReftxqW4U8mXa3DlkTUP9cwRAIYYb6iSOjd1krISUpNv5tEnkffbBf45lpCKHqEJBLTmD
Fw2bwJp2qJ3D4a5KMmZEaD9hk0lhN/DLxxeJN2vHw/z2MP83jFA0e+wFtByIex+ybwbkiVHQS/sS
6QgkhlexOMtMcfK7gOkdkD6xgqiku2o0OpoVUcNda2O3OYrbKsuAFagAobNr3HIBaWXWfDmsJHA0
OuxSowyp2rCPKUCs7rLYHaptZEYGhahpCgpAPEzdkRlpBo1DMRQDxKaxp9tWo6H+GwBlEU/Gworr
FTzhQJQAElyuYtaHXEOlxFYBfc0aM54gjsIlIdhKXdU1b6sSFh77hPBHC2Osviw7xyRXrvSbV4bu
thcAXpXJa0H+d0pxtbpM9qX5FB2253J4L5VrBULLkpmpjc8yCfXDsj7GihoUUoZGkNaWUvU6kcyD
5qeYq7V0eu/W6rrUEoSUwgGtwgD64oE9ryJdljn9VSnlE5hIVTcCCUfjDK3fX+gE4N8/P9iTRxKF
Vrxr9+Ud0s2JbPyHzmXxDGNaCR0T4RIGo8u8A0YmdGv3iHduOWb1fcjMHpjK+ZPbKlwMopil+czE
BWgGjKnNlnmUny+M+9+ZEDb2J5o3C60TLYncvqmxErrH4s9eBqBHMXM3DoxZL83Pk4/v/WUXdkXM
05h1jdWvr+QCvYi/Z6gvIBYWu1KmV0i7XaIZzOflcPLIoq2gG0eJDnKbK4FR0j9zEABBeU6y8sIa
Bdt6wtkVbG9cxL5YiKxHhfVeD0NM3dgWXtjr1eb3aIo+y30yUyJ0hNOO1J9c4NX79TRpjIAxem+X
BH6ioPHyK8DUrqzoNV6iyspq9WwTvCekCPPCCWGzmuoJbgDgr6gNf5N1Bd57qFb3BK4SMjLaXvlT
1XgQJGWFFxWNMobyNNN6FqJd+uocPr/9/hdn5+56OUS8lo3NopzbsfKY+EXKwS/wu62d8v822wRu
tQZWrvWPH86dsmfhfuoYRL33BZoyRYuOl5bHUg5TMLB13uWK/2aZAwZ8GFLMnQVDBaqKXlQctU/J
aGkKN/wprbDA5EOK8ieP7emHFtwZuNbu6chc2x1J7yahwspqcp2LKfpndzwy8qXlsTVFStp4gfGZ
xsOTE1U5VvMIiAz4SoT1dcsyBu89Hzz57yhGWbLT5wWR4Dt9kKHOHyDMFHoMyWcwR4MtL3RvkzAx
T24v/0R27xnUfPmnz20j8W0mIaO2Dj28JSF7kfLhV635SF5g/NcuKBC5XCBiw524tlhLPnXTLlyi
R0n0loXsV7xg5ItFuFs44N1xii5rKghzJmbNLz6l+QkXqziLsAlZLh24z70+98XrMLOox/UutIJM
b0Zrx+CnMFR+mRwMEyUMbIlKiBilg39MjVGyjmUW3G2HGD1y9d7J3TNy7vrhw360RELMvZGWo7dI
AYrGKcBeXnZ4IRiEEOd+fBths/9R/QVT0OeXUvi7c/5QxwfTbY7QA9Eo1e5+PtTuoqCakAJ9pHgZ
WvOBrEiNrn5vwOIjQfAj8b5O7xiGNhItWKzf7KclfUIa+cBaBRO0PqlnbQegnUYDDf3DxoxWt2jY
i0Qf1XnRy+ztoivAlLwOv/uxmOg+zjlRFeZ+vAcKEjfmpmSYrPYEQzkam4Lf5e0w1YVe40pgF8v0
8iVJY+lNl+qOd6AfjTSK/M8iGS0xu/ghRrh5FguRMeYLdv7CrGH8Pvk8SWngF9s59nwAmjYYap51
dmhd1IiCCGKJyhJvPLy+7tkWdiOfJAxLJnH/EXFwJXwQ2H4JSGwYg5NH/R0LO/daVmOUfM8LSHIm
Yr50u0gzPTFpMrZOEW9Ka5tZve4PPSiCXn2+1/y3OTw588bTazb6dP63Be+cXObZVZqjPVzEW39S
c1i4hNTWQaE8TqyF5MpGbEuv6aRSFAZiqb6O0K8AmeMHKAHnMjT/lKiQ6Lq9G7FDgFvcs0IsP325
TsQXp5vYdXOTHsP3CWUctjM6AVX5MEkN20Xb+PwWJqZkbXi+Ir4iaYOOJzqViuIjbmsT23sDAsqA
faFIeDAZn53WdSZ32vTfX9KUZgwUbjkmVUHnkVOXrnzuTLclUdwHCSYeBTjeWJbn34lbDEVL8ghb
qZg7T7aF6Bg1mVSMSpAObpv2dTaSvrGjvLzQDyM0TmCDWQ7pdS547+O65yyvTyhQ27PAZiOAkn8f
8dshi1vsT/NGyV8+EG7yNxo35UZpmsrl3ecsoITTYgkgplNIyhXkca9OQqNqzzue0Px6NDZsith3
se6ffaSMQSzXejfGUn2VZPhwT1wU+EQvoUKbiVr2/UjKiXhJjYm5k1KbK9kDo/1jDr0+xv0Y31h8
xDX7URR32wHtD2cHPuUtNhLX3VCerq0OVBtJ0AKblaKkfzegA511qL9qBSyvEOKx5oE+ecy6HRkv
Z9g+VaOrcd66IDPcW6r9XlPq5mvazuKVqi+nt8zmiZHZSWXg6iVdGNxti2vdMuWp8JZbT8JGVoiq
fQtwQwjXwzj+Er/AD88Pay9Y5AzyJe3RgFV7ypQPL87QKSvhfYEfB7ccMdZWteFK4EB/ryeCFAZT
eW4ZvSs0MoaRAijRF0KoVni8qyhyAkyhQDxy2eMT7Y6B8O/IabsaxyjejsbhGw+tylKLR2YH2GNH
JBVqhTVmF+LeZJpWpEGawZ9BAsOCZcCcZP4yKQFz+g/MiDjMmtmYa5hTrFH8BkWKhx3VKf/rBONp
gzrxBi5tmMZlbO0RsMm4YLCEpbO8zIB2vHH2rkPEvK9uOLS4NOKEd0JAkxJVEtZ5c4s+qXg7bpMx
JVnC4VB+bsZkxIM8i+/KvUrKF8VhpTRsjsNwagH3yNhODsa5pZ4PCs1UdAAoht/I/bnpyzMqPJCA
/VvQ9GlZxrzQlJ/UVPDn05GgIO86+UauwytbNd0kGy4vjPUgSpUduXj3oA39aDydMTHGBuncc1IN
dKJFfHnC+81ZDXBX0poGmf9Tp19fKcBNp4cO7l8i0Cv0ucBsoaDxSRPbPxBRorkZ3J7F5m/Kgj3M
pHWoqM8CDcj4tH68KhLxMPt6jLtwRwF6WsbmaG2IC2x/StoCcAI1WVMhXtVzjLmz83LMx35Zde1N
tqsotA4PpgJOXVKoXJACpDJC35rxsSi8knuBBlSBarn4z/n973JoiCIRBvgvX57hramCBz9SB2EZ
Eh156RfNPunBqLFEaZuxfuyL1xwW+8/UrH3z8Vd2RTb70ulwpHPSqDsrLwIG83wq3KWTyhayXAOB
tA6ftfPD9a6bR0dhQv2uhYbIZSIzBJsOjBJPbVkOn0ce62cHWTiUaEaQSiOMU5wxIodfvM2D3XEV
bOoAKKNS2k076zx5maU1RrvcUxdCe2yqYViIUEKiSPsD0zA/85w4uFJStVSDP+6YUHYyQ0qcWB9l
/Mr0fJadCp0Tq6lta9KXr4wo+mbWfRMMHYrme5RdFlL+/a7svz/+OY+7mhNDoTldsNZ2pV4d8E4y
4ZtkOEHGPqMx/pMzSVK8Qa5lk48nEeFj9dwo726kPkQOrJgvEusfa45YT+QkWH5MDQCGM5mYlyCP
cq0vB+GZzLp+5ICoydTvCxzh/66d/87p+9TYcpjn7iNn/cKxRlCgGaIGgVbO0DRJk6pHrxSXK+el
V0R27pfFyt5iJPj/5bzgqhtEVyfXNtYfIe/mfcOQjXqtSWaFOefg6BKP8Ke8lmBzg2mSbg4/T5QO
PpMg0iWVR01mYx7I42gb37JEYkNhkimz++qBAJxBUBzjBdFQCHZcY2d6rW+jTG+qIQMi6Pz/JKO0
zj/Ha1BuSXrEeaFJgtMz0cSdWj/Ee6SCRvPqC8E5W1WiOahWQzBVTZI8rj2e3CgGjiDRIbWZmpAT
WtyFX+9GGhvMbnL3gJhdaOSsBjvg1LbM32TguI0HY/BvIHDJOvzS0FOcL/6SZJ3J0I84+TbWfsFE
Cj+rut1mKaiZg3LNspcAjeem/i2gko3n1Xp+IEX2n3j5uGRyaffNBmj5KfajAuG/vr6QPbhejY+f
goQE8g5RMgB3hEar6mO9rlkOWYzZhStRPN8IMAQ5HsEg8ttLenFzR7ph7PeDolcyjYl8e5oBRMea
V7vcqiXzmpopjLif6dAHVfrVw7UoctYqWQ0zf+7dbRhFxY065UAckMqCu7rrlLGpyBdiWUJxxTgy
LFgTPjXskEls53Je2aW3JqWQkZOHt42o4Jj6xZUya+mEFCvvXG1uLsXaX4wH6w8aZB/fELJkHOrX
EyCCXePl2ejB+UhQ/xWTeSSmYc11gk8NK5OaKL2SKroCf/+6ZQp34wEOkiw2qVpcvIE1ENQEiLRS
DkLHcs4S3qWOXvl1r9w6FrBv91zi1d8QJ2i6Ydj7T4kUCvXLmSIrgduxZFqwnkl5IADspZm6huoP
dMgSiQ2HYZ9KUWfDf9CjEj16suq8EYktLttpelmo8SPBbPoRqkn3iFYvZqdxaYm9iXAbErPbSTfU
qfeCKWhl6wwC+ZR1yMrDWzrBxM+BTmeFKASMfRM4uvb5Pg9WvuKg/j1XGHM4yAp2cnHn6dBnHO7G
sGVgY6ExEZ5NGuLkVkP1wNto5eQXHv00IuNd/E+e6ZY82FEM97y+tidmZeVS39Zaeb6mzLk+yap6
IqCX6SFy3/yeWqNoOQCujFSu/PE8UflWTGRhsalcsYTccXKvWm9ZoalftC0aaEceXYEvjMmq4JGu
euN/9MTC2PQQI9tcjMjj7xvNCWxeAG8TDK9rERomOfZBemWU1SSjbDjfK0RyhXvTeNu2DsSaEzb6
MuTEQmow3Op8elraScYywJfVF/wU/7ui/64Q8OnNdv0x8kLccsBiuWd8RjUiAgEVEOdsCS9aqQqW
o03QVaGhNAj0YDpTQCWqkukvGslSf+PqKwjhKBTpggRwcDH9nWiok2rWXX/+TC+rCVk0SCOnzCw9
VR6aFlEUeowhzZmovewnrjiPQnUSPtKMgJkmsWp6tpl9YLjP8PFXCK1b2pC0DRtkOv2s8Qn7yyQC
ZgK4FEXd3YlkqSJ0p/lLtq5zi3An6cY2fs/XrCNZkwJNl0tEF2TOyAdHVj+vnZTvyY2DM1azmDKe
3I3zEEBF8xZNZXeQZe15619ZNE/13DONfQsvz+nIeh4vQaI4XvNA4QVizVOjgFFfbt53KJhPQW0A
Ou90lGWuGrCFAvccP1vckcI5KVtdJJf3FgKYWi5rPdniGSlpbENLAEf9Zi/a9zmwoAc7x7HL5Thj
qDy+JyGfFom1HXPNdtM7OYHSyG+s9wCoBXrLn0tcWw4ZHY2tQ4Y6dDx7I08qs9QJSllOtx6MYYRp
Oc06cMM/e2LcrhVQYAyzcJBOr1wj24YaxTV500a1zgT72DLyA+eJHPrnhwy6nZKF+xydV7XstlA7
nxflrWBeCIqAmbazpnBXa3owzVjgTovlwZFhv3N9UY8bLGdjU9DjWwXxQ/KIN9RfNE3kLcvU6K8N
4oCWpbYe5aDzSoHG8ml6gCJfGQU7XAqkUK1DL1WJw/kzgaVn0s7iSr1S/SeKctsWJXmgir2h/BUu
WRHdbm2FyWOmk3dgsr4pf5IT0budHVZlrvcycAhstRnEV1u5l9aB6N9DjNEEAdp3NV6wQf9nINUE
nR79vPwVfm2l2VfArg3nrQ8CtnaAZCuX/bh/iCWkSUF+U/l9bE6WwpN3O+p/ZhjaBRQ73wSNTS5z
mJHeFz8grq1HxSPCGIQtk2rNL4DestfhQQ17xMb1Yeiq2729oF04CpeqtUrHLXWL4b/sV839gPc9
gWwRU/ZG3JvQPuPMlEd6R8+H+Wl/uZmFZ00VVpqMGFZDZxSGvXYDCxH0heReGI3KAWoWw0ZXSBi9
AuD45Cfz0hTVlRJ1C+VtXEAEp1/fJbhSkk6ef0M34PvIdhfPT/SIJ+6qQKjBCHrO89TGoc+jRWVO
1go9IyBz0w0dDNZTn1qNyiYplhohT8HohfEwYgn7DOh7Jih5V1w9EjG46Fet0E10zryclBom+/9Z
ymcLpIgHBhCBJygObEjP6jeEjVgB5JbVZ70rgG09XCbbC5rXXfPxOuPqe5aHQUEZAjYqOIN7PsQv
VfS6JUI/FrowV5ps5JGn89xjEBjXhsxe7nDCyD9jcnc7CsI34HzYpll4mB7q9Z4KUNXCuSHfwa/G
YQWRPRlfg6MjHYhpqqFvRFbMHH4KiLP4nJbMpq7p7KRLSQ81bEc3TNC9T/bW+M5Y5oUSi6ccM9Nw
WyAiAG5XR05cS9HU/mNnxUb+uPZa343IhNAgNMMxLd+e+Vn+/us+LvsS7CbotzuLrYS8VnWPmz2C
I1Nj5kdlPXQGvojACutuHZ/faAOXHqi5VnVD6+nRNZ4iEqnePo/+x9o+w8FFBEwGARcDVkLMej7k
Vc8gw1LFTm6yn6ZeRX+FzPc9V1C0nVz3yAZhyB/bGCZrPT7ZO2vgV7D8nGkI9ATIq8JOOd5v3fqH
FWvGc2QVb188Bhkr1lZjhdh9NIgZslr35R/X0N3CHi8gkfU0pPXi4uNGJtRjcA2dK1vjBq8ylno+
NlWX7LT06Op5b+0pElfkl0rN2RYQNQsWqiDc8DTT08a0u0yBouFSgmsiJ2Z4bsa/wB/zcxehcbCL
NAPVc8PZz+OrIroGADv486TsQHy599Z/0yKETzKd3479+QauDcAhyAGg5f+qKhRyAAaTomZl6vaA
6xHrbtfVBtQrSb2eOrbx+wd21MCPCdSmtEFhIIHdDyZdjfmvY9SCCsAsHrru40nYF0B9eiv5LKiQ
tcxgJ8M+96TPdydm3Woibcf2wY5mzMreJbK8KlLjEQD+nua9cNcl6SLLMbO1Ij5dEKjloG+znTDS
KSUUGF5+R+r+jTtDt7YogJnROt7VEAmCAT8bUMEPGu8G8NOyddlSS1dkDYtneVjnCa8ELjjrJNxS
qubIX3xP9cFYsmQ/wivqoPcSSAscWzPCNYxnDlcRJyGai7nk6XfDF9c/bu6eBe9J6Nm3kYX1GVvG
Gafw65wsw9zQ4/Exdw9NjFwVahlKw9kpd4g1N7YZS6kXhnsUjf9plcpxHo+ruzu3Dd3+RK2B16O6
uptm80tixJGaFn5DTtV7OoskfK4L3xTjheJ7Hmj1wn/CwirYDmQA5/rAetDzaptlmQfzHyMf43/r
j9LGJodnCPCQ/jwnYdzRoS+ZqOSSUTty5HruSJj8f/FfcpkU4YWhN5kTgV+VMXT2SJ3j2IaQq4hV
dStb1mB2lbylVF6gENgg0J2Je6xLsoKyFyYRMHAkQ8nLJvavaki3ateHWmeA4Hb28nZQxHw/P2ym
fyFPOWJhUy3XIOsa4btikdJxeJWosOP1N32p3yvOnS9Ny221vvXrCHOb70a+p+u9usbSYBExdeGt
bEtnDiHX8h4L+R8weJxzLmlOWe7fCLCxoCxOq7qiPyYrt+Zdp1kPm+8Bq0XMrbvJLU7lBeHbOGia
Dg8YrY5uIzZ/z51Nx7sPdWRYCSDkRNPcol3YTWV+vuQEXJhMe53ydspf170K0AGpdtIkXE0l8t6U
zvq6D1osxG9cP8PQJ879k4kqdLGnYlwUuQAqlEiAeFR0S4dj2t5GaldTWL7EVKuhi+Kt5foPEkow
A2ToIa2TPxmPZMvhOaROXvt4giHyMtJY+S9fNQyhD9igbGJgolnPfTa7wThTCv0RqHLTP5MzBL7f
aSGzeMRAWfWZandq8LK7+zqqiSxwlEEZpSdP2K6JNaNowSc3uSRrQbIFoaxQiL6/zBKnk50QtCOF
3V4Xya9SAS118aNzNwbofH/pLLoGbZpQZeC9GdkcnpKoNGb2MwEAlktSs0XBCvjQGAtv3NZvy0Bo
intNBpel+8L/X09uOF3yLofiR37Ed5+kDe9fMxSpUJCv2jZSJdSfysoMHHVAqllB+Lt+JzXKnFvW
g4jjEi6sJSHQFQs/A9c2LvldJ4M6mfznb0ipzJcjRgzSbmZsMEs0Bm4sF4U8Sx12hjM+XG6eRnRf
XB8nmWDRpbNIpvNe4wSX88Fwg2jHHZGvvD+0prGsdHRqqyiF8+7a2mFusGd9M8SOADuNTbJfnDUG
l4/q/FsJ6xPFZCZU/LEdkJol4T/DCUThGt5q24IY92qaVWWtm9Ma80OtEkI4CUlZJloLqZxJ5h5R
/zdXbvBCIfUlBgD4MjKMJ2QybjxDfIBSAgr9hXv033EqFZgsTRJ99ZOunJmL8B0d9HoI8zhyuy04
vbh3XcynNa+GcqXs+4R+L0kxooJ1qMsuFLQucB2DwDbXOXBrIWIhw0DjUejLrVqya6SGraPh2CkP
+SoSkW85GeRUCtGOqwLLJSGx13bLmHSRy/Ni2Xdze7rEBiWgUv8yc83Ts9Vh3mFNXbHytRMC9eMm
ueXQcPBWUk4IneBuwpyWXMvI7vcq3BXCvnP3TJuSUxKhMEDG1wNEBo1aFnW7ggA5+L/qpZxI3afG
fhQiNA90teNKOORqBqFsHOK2v4jHgUw3S3DyaqeIOBsjpb0W1hsnhX9hFt0PexS6al5XcpXVRhMc
m6eqXXpMCnfqmCPTWuSgR+dvlMMo3TUdqk7KTNpVN7VhPTQ/XIWboFK045rSwnqyqmm/K4rHDHVS
My0UCHJNxsZgXkZDrsPwKs1H1geipb13qFIrh6T2hvnFps8Ik+Btf9tnrOnhpXmam8v0BeMXSdla
384k9XIQTs3NygqreWOEesdblxqkXKkthCo62P6hrk4lEzFQcFfRuRcPTPd2ZaJZ9JEO8Vg5knUj
Y8PwXCBSyn8Fh9iof+FEl7t1gTp6Irjp0dJHzP/Jc7XYPpKT4q87MThl24XdP6GN/Dm180sksXiG
wh6YOSCPu9g0DK8VWslM47CU22oP6xmV4ZMIYUXSMwZ5GhzGvDcwkBTy3ek1NQadu5t/bNgKn/xR
QqHDPq9VTEczghdG3taLmOTKicvTPn6WI0oRGd+WrnAnZi7IHNmIL2tJuxn7Q6FEfHr8F0gz4cnp
vFpJ1bO8PmiJxWQ2hvzIRlG/UAA+1/rYL/WlmVRVbyr5msaP27ZguotHd1PCfgP7zIBCwjDo/XAf
YkGytWkmE00T3P9m8kUPpeXfrZUk4g/ock+bRhxonyDH46J5fbccBogQtc6TrONBrvr4Rtc9zoKg
w5mSRiIRI6BeOjdmENPD/9Tr5W9VZdLDw4sqYbrfa4GlJngKWqaBgiixZ9Y02KrxDhj6QobMwE3r
mr5C1G86CJ/ismIAAHfUW/PKQ9H3WhEdt+BJ2jcC0WW4orNBIOZa8VjABu4q
`protect end_protected

