

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cPZ8vU4rKWICMycnP8ASghxteX0KiiSQpWJpCIK7voNSpkWhaLkY+/QNXKrCWexA6C73eW4MlVqP
U/aYYyUL6A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LGoeeEeMUHkj3xBumwl7JSHXwdKJWR3APWiWCdcCy3wVC6g0GScQrp7fjvXp784YBiHqjtsyG69d
mOZ3fy7Gj87kc/h2xvc4Kp6GM/IiHJc0mbPVp01AJelfAExlIEaVGoQkcAXR2aVikeaMxuRKkb9m
THdehu5n5eHx4/tJQjQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aia+xx8RLMhA3IF4tHoW0Vw6LtYVDVgU/c3FBWk9RJ/SaLw9lkXng6eXJGNs7uUJXmkzrbSEXjkp
9p7xWJMhovE7nwsp+7RydSgRQ0ttqPUbPZE1eqSc4iNU9Q/KQ7cPFMFwb6o48JfKidjAmSeXX5a7
n8A9TbJ98klc/V+a8Nj+tTPfVP1QI9dRmdzaW2w+actp2BkWAgSALKaGkzvCVGa/MpfN/fdLNjxo
VsiL86HW3arw5N+Ra4HD3GVUtLt9RoCCVRrMaYywuIwp2m+MgGVDwi2f2wZCZ3t03UamXKangjoy
PBei/XvAf3p1OvrOrKNUCVdwEg17DQWfBwZyYg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iSq3so3iXhp8LA8lrAo4ElVWkZ4sJhg+rWrioZWefLcgVs70gDbHsh3ghf5w2wiNXalSfMYzUoxO
skfS1+28WFbvBvygndpiSNMXeXmzWGrwBeHtNO1nR5azyndKvNsun44/B61XF3kTINCJNR54A+3f
0Ezm1jX/FmstQisPDpo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fHCdwSqtdLKfkpdCYo92uS5kFXmPpII38bIISEYuCqZyK6/BVCrCUL1HNVeJEgqGnb0uRqkye2CI
eX2LoUaDxy6iVejnRrRRAgNtgrlZcFVc3u1KxZQXk/12l8pxvVZj8jnWgIvX3TEsZsoZ6w/D41BC
6xhd1LtUfJeg6bsnb+yBYV5+H8NnHOqkZuFtJBsUzS1+4qFALyFqcNVJhhbdB0k2hn6z9cG6wZBI
hB8OJAFj6xON517ug+qP1OJf6uK1rHsG0pxYXoT6xch+UowAmLY8V/4+ShcI8rx6DLYpPvJVhEGV
fj/RQD4+HY8CEDIrJcGjF+Rpk986lOFjZ/hvRA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11888)
`protect data_block
3s8MjyQ+RRfcZ7ILFm4Rf8tyrojf7fJatd6j4Q244Wpp/dmGcarnMQdIMAL9NJBZzNvuddh3TJLN
3vsgVW40A2VJ4kYTPkrJfgR9Sotd7TEFrv5WJoSSqt086jtWLODUahjkQmfgwbVzRByyLkX4F141
rxQtVf4icJ9yhNndDJVa81S+t8k8q+uRdw+a9e55jbrk5T3B7JDwNkf4CKgmPw+CwC5AE99UWGMH
0LO0pJKyI2kQuLCfbJTH/aeYU0a2qK5OKMSR8jmSbRSSWmwObCTlDsx9Usg3T0tgYhyiimFjjmKp
NjOcAJCodgVfkH0SyKdwRg6wPhzx5nMspoqv2LFJNfQw6fuc0rWWaOzsF1tyEEsDJ6iQ/wrIXFu7
wS1aV3997xAD3zV/9BTSqfnzp9rQUI5oCpyM7bsOXaqNUz/NZNNYtvie31vDnRJ5o7WodI98kFMX
gDh+gipcPdmJRhrNjGmflVoPFDfLDxJ8bva7f8nuNU4gjoEhjPH2NSsQytfZQR6gyHo58Bv4tv/r
nqxE3i2VQaXZPfcpUhZc4m6Fm68NvG4Dn/+7huc/SuTlt3C+IY+zKroWwEcMFuDC35WAyuaih2lK
KxjQgjKDpquSWmag/gzE/ICbMrQNRqc99uxAxReg/A4fPoOHC8e4ORDuv2e0y9MT5FZzaf+lw2m0
ZkTd29ZUsflKi75YkPYFBIh+05uhMpJmtjRbXYZ91lpqY3+afYlcqj+0DlEC+GSTG3odWJuKp2VN
wF3Y41DjL9M26F7iFRilN/Ypz4JiPsguIy3FmM2+vGBWH8EhfCfQQHPV/3KzVrw8mf+SebuHmaRd
5bYDF1OU8BflMwLRxNjPJ46Pl9Ek9nj/sf/CS4u8JxPuyl040C08JhRjKAoGL1vLtL7IW17HNRkA
A338H2Mb5WXcqDNts0cVtys6wsNRlTaCsfzL7N8YXnxAEQudWs3ultIz9egMY6NLiMKRVlpWkU3C
607/gHUwsPUrLL4qLa4TyyrdRg9gcXbGY6RtjCbJ7xnOc3f3U6L1wxE6Fm7t5q64Hgfef7zkTp7m
4g9UQtGIm391PVxeCrP7ZVCVA7sfsicNFjrYDD8BzmPHInci9hbmW+dU+HsQ73xIVI+MxrK7bXa6
9s7tPEOnfGBkkU8jGJ7uFoUYqdefcz2KQR7W/461qoCjj7+HCL4zFZd4jcm8l2yO5VW/UqJAr657
o5S1wSp3tcxR9BbZQgooFqG+Kex+jUoVtnHbjAjuVWfyqepb67cgSfrBqZoaqtGQEisxEEPisqyx
qj0Kk2bmtxdpxTr1be9hc5vWeOJz+XychD82ilLONxnNNps+EDYwDO2RmcdJtOJ67F0pBWnp5OHc
VOYVpRmoY3waGRtGMtt3z38IbG56s1jERMKJI6iHLv99WRLwJiHdz93SyL2BNmnkBdFi2XO9Z/+3
NmMWJFM+mzRbARp9fnYn18yc8PfLyPremNO+t2BULrldXhLXbHQewcqeDIO4/5sfqv5IKxHZabkP
nwNchuXLT1YK9qCh06TMMwpCQhtpGvyXtMkrWB53E7A8Awf/uotmRn1h+6vg9DWG7gNDzhyBsG05
y7c7S3wSlz3stnna5mx5NPa2b1w0IbVuqiF/Y44/hsKuDr8+FEk4U9k4qBawU1ENlE8M6tHvuiKl
dFR5oYNQn8bGpX3Cg8CY7IM2rNPmDU3ivrsEyKxj+KNDYY4qS+olM5uafA7HltjoScsqeDQVRCQt
Ev3SSrscMPd4wVq4xjvlOGOorgWWdFCrQzEIwq3NxY8WO+xK7wt/yxV6bOZjaMIvjmA7NpYx6MrH
fb1Z5r5XWKdA7yPeAlLaEnKwonNsBffRdLDG37qem5436E8T+77X6mzrYVIOXEwsXOukjHnwWo/8
Zifv5hVerl5w7I6c96MByObWlGTdAcB3EtqGH8kOL15k3Yfatm/h3PJNUxpjze5i0wSev2Yg0824
Wvbv7wq7in/wSw6JbQt+a30S7WMYjR20nV67r1gU7Yvka6/lCFc5bSMG9nbpvm6UfVPITKe6j8BS
q6gLz59vC6VK7ZArc92LI7Guiaah3b8SU7nosoU/qq/xXorekMlqSWzJof6K5p42n7FOq49tQsKw
mZnTHnGxG6SbEYPfXqQYcc1WKao0s6I82D8uzIzDI0KiXJEzIssNf0UaPoXUnqtGnJIqAAWtkD45
Ah54xjWJKEjSzrvZKuTSf7sgjH3dHgovTFaUeBryyGBKIDbfATfQF+WgYblMBQvPAX7LlQe8+Jyj
Mhxaz7m/JQIvb36U7dLZqQnkXS+UBV/UXcpGiUlp7f+UZtev3bLoEfaIMiw4FaIk85Faf9tDBJn7
pkEdwD1ePgaME6xwqn3k59HbSkrUVlF5n+o5dwYQj7K7+kLQupILzTMCLDvMyUM2yUi4rwLmXaTt
qVXmK+Cbh1XgHG4dsN0UCV1vz68sJYpikygpSK+ygq2NhjzdlhvSQEOlgLxPoh7XseipxWs4JnAZ
3/9IeQWIE9N42pH+H27Ro4uH2SxCNMVinia2w/YiT3O8CPs1nU6P9439KZnZHVI/FBw/HY+/SoFz
S3EruSYJ0ED2QYI6OYtWzO//px2r6plMUZcL0VEcXBTbP+pVyhpXofNeOe9jY19HMmc+QfroJlxw
OI1wqix/0IbZ43N0ZgRVRrJIMfPP1IlRVTQk8vB/oKFdQHk+5vMd20W5w8hqwle/ew7hNkZc7ZDS
gxK/ttqb6guqipE38bI+fAVo5S3P3SWxhykqt7wGVnAlaMkfCYe2s+G5NBD7vponyIEW/i2Q0x8/
7pad+pfYcHuOn2r+YELEQ76+RR5/ygTek/zyrFBEUNd79338b3p9IrDDYlBX2NBKXGZKkFuAYJGg
HiNX0sCgex12VUdya7WVd01z012zSfstQ2k+BkmD66+ib+c7roeWNLMUz7C1Kjtq3hKDsriOSD5L
BKe4wjZJFgSWTlBwe5qtADHQdHyiRBTlLdaMyS1MngqncBkRiDNE+ZUBmGU+jcX6YbZdz4xEzybg
jWHopJTO8/Tz2/YRMGKokWMX5kB4udD0UQgKCuwpo50vZzQvFXnkN5IqPTac10qgSJERmt7P77LJ
l3bDWLPlw/+jsG74F8q831dgtJJNzWkmrXdO1KZ+n6pSOI9SwTJkHU42PFFFAEB77zADHqro05VI
SemWKHNWpRbcYbwPdKEaAXWUxPCsIDZ2GGUreF/4I7wMjnwuDEoyD0O3+kfmCBF88xEnCHOz13w/
bHTxPNJPir0pYjg5xpY3Yk6KswqAMC3az2Aj6Xik6yFvnN7R6UvUB6ZdeFApK9IQtoX8It+SJQSJ
fQ+SRmaxmmIXxYgd1wU7JC9YE0P8tFES9h9O1YXCzmdAg80eqAo0I6EeFVrwIm0w5LH94CPVU/sc
EjzuXYEet2hnlaAfK7KimAjMrV9XeG3DMtQjlJpXdoWmGQ6TlbuyT0kHJaWrxStNpbbVSzw+t5wb
P+pniE7bhnBfwT6lYtarwlkws59aFYOE2BmulvrlBwMyGs0BZ/11nss7ctderVDOFGiicETwliq7
hVb5dKsTHpX9TSY0T5K77RljSE4OwAdJ2mzO08NLdnzMgzY7oi9LsZtFBEPl35X8DkzjMqGGGuW2
TR28nLmPGqX8B9Xot61IxMwEF2/m71VxNVnIQHbtvEVc/AZt0J00+JSSaaypOhDCtv+1tRAXMp0o
KOwxP8fjGFYEWoryE6vntnIvHxyUN5EcmtAN+CCeuyQl/1z5RB38yycfE8h3qJVlsJvLFjYjg11x
yUyZolGoRfvULfnJ0mcctwPEc8aFABzRxhQlnqP9zSdbXD1aIXy9yNqx65QLEQNQjYC/VmeXaBse
W3WJgxl4OqZvPl7XxV7YBE9OWz0gcbZFAdD/Q6RC0BKPR+u9Oc1r45BJp/1D+k2U8lmwsGKbJU/o
2gXRLu8wbQy70xPl4Sx/4y9T7/tX8P6OpfpevzqVA6ZgMVDDe6N4PMk7XcQAitgEA1fLfncvMfYp
dRzED9o3LA4x/3srGskFXssTCQRwRHp6XQLjeeRT6QfFYw6AL2f37sd4jQXPTBqMV98X9ylDAtY2
Qb3+YEYoHjLxxwesxQUzEi3qQU0xjn9RJS2IssiPu3Cpyp3u+Cy+G+boFGdzGEr+Uz2FveTLaKCj
nTPF8qGQkrbuoDQtIeFOv4HAgZieHUO8ogSu6K47C2s6rRrcwpdRekh6n+ATZ+tllxpQLJlf592F
N/VR1Tb25XARBV7aGgwzzODQx2rzB7lGvmaRdYGPmCtw88PQfwWtHAberAL7MVPBr+dLL4BtQ+D6
VbZ6VU2/wTJjLqN2Bh2Sr+muvKbPTpxwK3U41OR4rZ8sg+VbjbBj8J0DFj1wVtGd2AlHEhIKFGr9
I2SzVgIRzZKjhem/o4SKoh86H+yfuwLdbG5PACJZvPrrxEWPg6cb3ZLgPyh5bZOHZMXNttrgOqvO
5+fEIdVFSNxwRp5YHMOhsPmKfL/sKy0E24jS1Wg/AJkLZV+/5QHnFcSqf3MI7ffuI1Cw6ShwfycP
QW74nF1tEj8aTQxE82A0TJoxfIDVsu64uDUwJmKWXGZKj2Q7AxN7aqToDGsD61PeLi68pN96xKmT
3x1kcC1VYinMt3Q+VxiELFFo29IRlKoE8qRCMNYQhYgt92nxRkiuRsnGxmWx3IoLAFP9dOvzaXZZ
7gR1S8rBNvfmbGtSMLO4SJB0IAGX8zBwCdu7QGzdENul27kmdXso3iWZ3pOysC34jXnKrTyf5yfw
lieGhD5fW/l0qCwY5LxTas1Qm44+4A7MdzuYreLgrzR3dBk1w0bkKmp6VKK4nnhjhJo8IhRrXfHF
2dU2CJ/BUxPimHULe1tskiSrHL5SszqvYiUeHgY/v+ZIO2MIXnxGz6Vo/cIQCiOPeP5xPCuCiaWm
ElAd0TZB3HkOk8NIxQZyguIJtkKT+SssNQtJiAcprwRhR1eReB6AL2LP+Q1Lj17Ej/+6iLEyrfb6
rlMyHTf9YPjeVh4FkkLgwF2aP6myDgN4bkzqzp1XdAfiRHJ+FNwV1Rk0sB96CwKnIeY+bFRv4Ttd
baarIls7S2Dhus2f4Sd8pLeHtxP7aLbL56QhLbShfruw3I8yx+jIM/YmFe6A7ts6PAFrZe1ys1kI
MsZcY78eCcPJzour1Yq2/eATeMqrtVk5cSN2B19xudSyujzFMTUSkqamEz09KBN2P3lpn1kot5PM
EVxIYXT/+xOyhQ0RfpIQNhvHYIjdmi3QouevAYFEp3EwlYkG517uKRvULOBk27ozCR6TMEYbuwtC
Co4umHTas+kvQqkto8b3vTDh88viOXAwJNdm4i1ixlr6FKZS61pEr2ZGAO6/WRkFyZtGLBwsHJBp
rOfXUMlVSqyF52RY8huNvhJcoiFZ15p8ML5MJ6/iMI2Bww2K9EgTqILlwTmAeIZfFlK7z5v2Pnp9
l7UujGHeFeVsKKAt2GANkb+zv6pUy2yMBzNyYWgj5oUkHlD1fM12WTjAHWr9exZaAFzzLhdrgn+K
O0ibXEPI+d5PZQiklXfhZczW51qa2bWXzi+r9bMaYFq5REsI71BmagSwwHFE0SkuiIhyq7z213+0
qGKTf5wqhJH5xbt91CcH9gKU2vkwM3uoXlqxOBsWD1+3hyjctIEmLzqRwkNt4GmcaJcy5a8LLECP
1ERNL8xn7CEUC9lYVqBJPZyfPBfMUO6od0ghtHlCYBe2JZT79mWRmEk1NfMIo/i6BLlP4d8vRz8I
eBnXEwsZyFYHeWprMQmIGNDqPanPsC9qINbITOIpn2+v/KPcEO/NO2G66qZ+wtpu43iyDGs96s8s
fY1Mfu1faVK3qABtVv/yfUADJRMN1Z2GFcln2XLl9iNfi7lfWgzop+NA0XxUcuRU2iwZE8Sfnnby
d52lJG0SJXT2zy7PgDBdHxWChKMx3thrdM62I/qemCEBHqttn+qLZR9c8uE56jkEFhj42EsX4vaw
W0YYNqfPtV1BjtQi6YsguVqzMPjdtycf861F/2pH8i1lQMsko4uCJlCVjy0NYcTCPYMmfcglgUtV
YZZ8Bco9VPv+K6z6FKz0mZwDbKyhBlyteiD0/tiuNh2c5MxrxmDhiC9CAhiln+9l0ko1pwrRPNf4
+FTbM/MZt7Oiy/gvW9LqFJ9VvYzGHxW3FlYvZywEcn7CTJKtD0Z88kSgy3rzjmm/ja5wIvktzhEV
VIKrTkQ1iMYtZ2WySGgevul9gRMNuok9uCA4F/sKOY44ci7YKjkXhiMlsphrCICEXuGWlo4h/6K9
Ggy9oWV1m/mlrShMA7cX/Wil32gkG4wYbzZlHy5WCZEGyTLIKhxfJzLn05RPYAYnhSA7y+iA9dVh
af/pFvzAtbSsA65mhdX2WBx1NsrfpoP7EZicPygI/fAqt5OA0y93SFFojEnAi73D6jfCfBaiANdX
xa4fAXvZ8k3RhJ2Wrk9UNgSO7jDCoRsoa/kKqBfovVfJjCqt/0kX80O3vihjQBUMlquA8OxCvbT0
WUVdi6B0nDRivNzcVGA8d3NAJ53oBmg0mgLLxLLuyiPKkifSRZnpa2zk12/LDLILz7c6Lq8gZ+pU
IkYB90qARJXQdSrQjiVpZ+iJaPjv7EE6CxwYDLkBmCBy8Rb+MHvbMY/xYCIbR2IrETExYexju0ff
a9Uox4v2QCLiw1hJZrHDsoRfCV1+I7cNgpsVaBnpNls2swSuzkxiEtNki612UGxh1vQTT3PNdkFS
Ju2VKG89qHJNkZiMyrAaMLZRwt+Udlrp2kusq/SE7YIqTPCckdWjnsQMkmxEYybyhQs/6BR6+6Ey
8iV0aJmSYrtmnabzWWUE7ekNGoOa3ht428eqzKErfoF1T7noqZDnaZMJ3rmiGG4UqFL6k2a/Y1l5
O6RROZxZ2gm77qSRFUhtsCC5sLUTeend+cFFx1tGfBIx65al31DjFlcMP92hdJunCsSHAFPjcmDD
HXQvxTaWLNB+q+45wa4DZk3JMWLn9Nj+9OY1VRkhwemWuS5D1NSlxL7UncdTVVk0JqCHedbmlEkc
tUcDdBr5/3vEG6tmpn1cNTDiazRPzwQ2411FcxN6Rv4+ZJw6C7PTfvpqAGtgAiEDiEAXizQ5ns0w
i+D3qITPTYbIkJGOYRjsi4dBKwsyi8cK3XmWUPxIzaae0+fDkXluBFbRHDMiXyi5hJmn+2XFkIj8
DTDbhuSTWmid/7VyAb3mykZZOY4DU8qNbZ7L1exsxDMRuJKU3URBsB0WVYbSZ41ixnfLqQTNrMVB
rWdRgBrwowGb51YR/UBlABwUdFPcliqYAVvmUPOUUUr9EVhIJAp/iAf+/0SuR0Ofrzm4Hudckd+e
qlvsnjpoeRuLHbiifgFANxNAbWdZICAawzHgtLJOLnmOrop7+5KcdZ0GxD9t62eZr4oljip7vzAf
B94IvGHoZ+dh3orafvr9BywsVN4ai5hTklwD5uA+CyV1CZcbplRmt0xX1V8GZKipJc37vY8w0jDL
e/JM0T2s6/wCORuGMNyTELhjVtQD3Pt6AK0JXI8wlMGYcrk+PIQZCiiUhYYTSIb1tZ9ojUJHJIGa
v6Ro0KztW4A0BLpd/0a4xdk0OguQ78Bz1FoRj9Hmg0t3jK+i9wcCVUGFzKjlEsgzh10z6we32zgN
tFe2nwh59nrvqk6ckPnsd8qN6lcnOOlJkdmF6sIOFJz75Mfn6aoclpPCtjaMx21HnfedJ4o/Wgjx
ytVhTlE8uxE7XSYG7YwPdBAid6JG4jWsqqb6Dbc3I/zi5fzqekI70+OP8K1CJgVHSDGqwdS8Bdj4
mwhdHmh2wkc/uJd9AYhCJEVK3ARMQgWqyyzC2sXxnxB7MQ/fgPs4zd6vjXXYThLgJE11/tUOoAYA
aCpQx0XgZRMZXS1EocPx8loV1IKn3jrgYdKKYWcjrHA7zHywT8PxoCofVazDZHgnJsVNU69ySNeZ
SHqmImj6fh51dUmNEGwdGMHWGVIBlbwwQ2mgV++w0HuCNF1mg9vqRg7GBo4iimtxs5DhasxA4bed
qQGp8YaV7OHyW5lqLg3DYAEQTan9sng++UbGyxtqeJPB5MSmdqMNgiS+ZSRHKa2Ja3oSDKMg0jjk
Z/yuC36BpKvrFLO+EaHg4Lk9YHKlLO9PTPAQ3gRo8BPzgADRKTICo2qD5cBeO6QPrLSPD6bnlxXo
Ros1yXPvMBJ8HvlzEfEIsBPbkEnGWOiPQjTAkWu89zzxNa46d3kCX4YuL9MyIoc4JjGlETKkB3ID
PRZbypjd66hOZXGHbN7NKuHDfflJbHq8jv3lP9QAVEz6HK8IOVcGmKCeCSl+FSxmXF3ODpCM/Orh
WoWYCqr+bmNab33UHd69EnY1JEVUq35dUAKpNOH7yU5iIdeyRlsJCzzPe+bM9uIxPHLHBlAQGrSM
kKnr4R/rOBTCHuITAH0eQPtXSo4u9MHGw4to/y7TIdFjYkLLIY/+JjuwcTox7uzUdlUhIgDZ8/r2
ROKiVzdCYNSp62Vkk/zn3/KvO4C69FzyQjIkLrp3aY9u9T64uGT4fisQKz+BnAoy6wavUfcITs/K
B515J5J8G/LyiFE4OTEdVFi/2DMfUH1Wl7t3laJcsNRS36MGj8B5f1DpITypnFFxLO0nRrCDlR5t
3COlshXB/qtwFVu0Am6U9Wvg5PoQa0+O/VU5mxbMXorVaLiCZzBmXifmFCcyKnsYuuPvGPzvDAs7
5E49c7AShvdXHvoaIutJ3N3rZrOCBAQS0lENyrguvUG+YrKC8JIOf5cgZWSv6V5iMNOazxsQEj+K
EFV+i1bt9HpUYk8KOaXsSMUq2FlwtH9VWC5JhH3Utzm2wjtcSNARlyNTG32xNx8YEXR2Ch3hlcGS
hoFsA3uCLBn+qMT211o3SG/TSyOJxe81uX4Ho1c8mpS8KwSKG7GHLt0QPfPdkd1ozcCsi/zXhPPK
mXMN24Lx8AnWmUy75CB4m/C1dfSlm7WIo4z41cP9tI1H16VESN1NniHeIdq7fdXcWXY06MN7B7sK
0I+JwjYKRID+6vr5+5xxedLk0vHoh6yU7E/8fCcw7gCep4SVK+Hl/5e3d6N6yNMv1+cceYXoOYAd
3dThE3L3DsEBJqMR1zXvdrJfeFuvCZwAd32cAfk+woJEw2yWm93YU9UgVXbBRHR/QvU+eeyxAAbE
+QZCfc7+5DuzhLUcTZej8XDlIDJchzKBwpNhS12brZO/oxqLJKK4fR5OSHBxlIoNTTih9N4T1RLy
YHU+UWr3smZ9rrF8Eq4uZGuICN/i31jee7EL3q2NpLLNYX6Ixz+FmH612iNh8U2i9gJwewtJXfum
qvOG0ajpBN2UzWyJLZZUAXhapRjMu00iyzkGOpXfZiHVThBR8ROevPlk7hsN+IZ+GaPEvtQa/9wZ
JgYmLABvVHIuKKPFNNgo9Fx5/PhaBmzpKLRSLEk1FtClforleZnmgx/9Ve33JO9dDMUbgGtHXZjB
fasCHb3B0oGgTLxJ3O/hRZgRsDXUYxrtUwBbAZW1iMMSKZHS78CrSmF5PBx/p1IpBmYXZ+48uBGq
rSEaUK8x+o/TbCh868xZZNpgUFkvRCh+YPElcCAzDvSveD3hicz1zDWZmJzgIasPOax6bt84BRPU
OrVapo2OZJj5YNuzm/jzyQeMY4rdYIPvE3mzzJjevOrC4nhqd+kvViZpgEM/W9fDAAXxY+bHf1ED
RKzGyOntYQOP7Fx7pmNS9AvvZlqMx/x9sLnrC00EdmoQhik0hMjRbDIaCp+ol3J48aHlC+QxCcFC
l43CSPiyk2sM6UBE+068LTUtQ8En3AlcUla6MGh45aelF9FRNG84W7TtWfK3YtUVo6O9esceJALq
7tXD91KLAJBqT6LOs86LT9lr32oOAT9RRvUJ3+e2C53RtruXBewt3eD3XaLKdsG6Tf7OjqZdavpF
UQcsI66jrxZnykxzI7Sb5wkINUecX+pK/M0LObdfZimbK/aHxLlqRaBZ1A2XaB6MFcd9U7sOlHVD
nvqkLbbRMPuCT4mvdp97E+h/lzSTwhPOqqMXYTZ+efvjeQRgmGdl/30HcyXkKTDdaqCOcpy2BQ1j
iKSYjbawiVu0/TEo3YCKQZMz1Kddj8JrZrU5JJGI4/x/kd6KU6AFOphR9cXBVN9y2nXy5e9ZpYxf
NEY8/1Zte9aNpedA2MGXF3DuT1AHANU1QRaHPsqHnPOIAWl4gs88G3E+4NQrxsiBrkWj+gEJrDPh
8SSBrVe+Dq42+mkZX3gdsKf0nvfPdEcDdQj03w7yiM+Dzzm0onBmBrGIIpbs9fVO8wZKAZl4KuxZ
rGjkG0bE9hLre6x2GC6p9CRoK4FKoAnlrRGAXxV5jDILp/Sx40JGidba/yR/UR2gvGZ92ki4ffOr
aObu1I1InjtYHi6WZKGXB2Xokx/31V3B2eT+JZRoorPORSg1u4wURPMoeRB9zPKzBMJiaJVrKGsk
bI8lQsHfpbHGFDzVMXaczZKgrGZ9TccZjjzyLUw1MDmgF2TvNW255JOOVCsKqrdHaW/wxeeq+Q8e
E76xgU7T1qpocLF+krkE6yFx7pP0+1hXVr1YUHV9TTqs3TwfkGEJNSrC4YIA55daGr8X1uL0zYfr
/SWdbzGpMop4FxtKl9M7rxLzX+9UVls3Mq9liPm9JiMvbvxcd8cHQBDGASuyvgTU4fbmwTPOReCt
0j4fWWDwqal1xaRmblWgF/SxjbKyURjM77k3WWnEtdeKgukzvX3HRW0HihhnTiFdEGdprGq0kDZw
YKW6758cA9XDRkvnsEDaWmvdLHpk6GBdQyTf29jMZ2vVgz0O8U0c32hRA93LneOOW3taBS82wMTM
MJ5+6DFrXq2QVejrl9klZgiJBCZsPY5nycI3SZMaugdse6DAOKEUc0hS98TU3B4Mw7ZN+Iw8CReE
iaJiO61jb/R0+MPancYerT+5zjZuoEE28UWD2la3ScapiehXqlYjpDuXJn8PZLRk6fbVunHvkWnO
DetZCkFCSHEphkTMIVlR3Too+ZWDogBZDvVPjZMT5wkXBL0ZnUv3nFW8Xy2RgXfhPwo/dD2dwW3L
eB6mazMt5SjGlhfFtDcqrzrI8NTjVOaradFNKXx62Sa0FMPPgZIViRiyewbKLDGKtHxaEcB1epwf
3ZzNl+JMx1UdNYYbCoQBZpXMaRYSCTfVqVG7cuZKlIETQg6n4JODT/eqqNX8S6Si+c9ab4f300l7
jD3fFQ/lND8C3o4+RMwAmDP8CjUZfwLElNyKCgg4/QKjN16CLUVAGbhrASV0HrbPBCxs9mBYUfCJ
C8sqGCVJ5aD3SJXXkGPeEiRpKczny5qOd995IjX1xIM9CUG34ToQY1WQfOUzHwhF8JCZR2hoF4mD
dx95sSl+eKNty0NezgwAniwRzdaydXNDfcqHGxBpdplsv4n60XZzufLUT4h1iwuO+M5719L5pfw9
ZmzG8b6/KeUGOSi61Q8WkcZ9ToGRMaYLYscgxgfGFRTKMEQWOxK7MPWn9IYOTNl3QLPfta/ysow3
PmS/vtVeD3SZBYshPtBJgqpNhF7u2a826JETuLUxnyUNrb4cLFIPCr2RevdW9YEFrvf7yb9TU+I4
RRTNzDDkwikKbUofVNcqGlIwIX0Ncl612TpsQqmVW1Vr9k+b2wbrPaREYY6OvT/6HRVILpkzriFu
VYdrdjQ1PCGJlce98V3wXfkBWRCLTgg3h+h0dcurkGnYDqxBhzkP1dEMVTQsGI19vIAa9qRL4JpB
gW37z69IAMKV5cAzvJBF0hOfvjlpkbQXMn0NhGwB1gNol5CiGBYHUDGRYs80d6/Z/jSse5mX8nuS
kw9cgeche+xpA/2OkG3Y0rCUCjmiFGIsvzP3yjNca6731JWOUHWb2pZ3yfgAV7GZVp3UEDGVT0vP
30aWJV06ykHCAsmBkt6BQ8jcM6jbQOIGLSRBSMW+vn2cFZCG3eG9z2e14JHdFh9b1HfYi7MhVlov
X5owAMLFmkCCqVnrUFvYZeNxyMrUw1+hhxnrUEqDKy2BXPEgxH9s7kKjnpd0DSDbFORJ4ppJGFDf
NAM3jMND6bjO6X5jkyM+cQMtcgZKSgM+BDBohDl0xt2DajUWbGf0KWUCNzClMQFWqdG6CMnsBG+p
zDdchPyuhZFB2p8CNYb4lX0j6tT41Fu4BwwhCz2OCLx/uksWZmtpNYed8ComBph4wcg/mCuFb4jz
HMEE/wyFR4MhD2u8FLu60eHEaH/+9N1GTAxxscPISHYUPEttGNxpHsa0eX2jWpJenWCMFZ/I2hmA
7uP33vVvZC0au87chjEZejX6Bb+2kQ0JEHi10FAKXsBu1e4VbCswmtHYnQ50i9BR/DteJpNBo2fK
IshHXi9/Q6y0Nt6QfEeut7mBtrDvfhjEwLmX5a/YtczeVrEl37UjdST+2Fv9RcgntiqjKVCNX0+k
oHv8yAwB012E2EKMwcjxzjSnp69SnW49fABs0/5Su/ksaMCoy7zsYDWR5OsyQddUzeHKiqGNc4Oe
cgayo26mJSyJhHctOnRvz9Eo5VLKgzQiYcqBkksUwwiixSulCxQ3o8ng8vV1V58AX6JxIHh70qZZ
+lij7BslSOQkouOK3Vz8hxAQOJ2Y0UC8xGpqE3BY0SRf9nw7nX3a2os9HJEvL42Xi4L/q6oUIs47
+i4xpK+s1kyPC7237SnGRDTRgECKJtpkYvXQkxXdfbePhAzeKETZcuREowME+b+SZ5DumWOiqU/I
pX2ETGwzAqhMBvEfKbe1sxJklveTfC1FgaVnmnDZRGyPA6b2WT9MYeln6SAnyme+Hq99qBzG2H7j
oulk/k/A3964RP/8rgfU5b5+XL2+W4n3pO0zFSIQqFldw7fRe+nRyCNVWHAUe7fUPCwmjW9mPSRX
h6iAEI5d4aFWjjF5ZzjcikHDM+MIs1DcO7Uk/3sqc4WBn5uqXJ1vbtg2o88RZHJGYvTer4hClpNQ
Bq/Yv9oSNGJq7DKKkEFljzep3MS9frvvbQuPz0mwhU7njERKXaa5UJ/Rj16dIsrQJXD4icgEn6j9
1Aa6dYrXy5bFvpHk6a1vFA7ZWeH9X/cut1sTHpdWOxE0DkfsX1Icu8hheJoAY9zh+Tk3s/B+Ds36
KNj4Qph4Ssmvy8kFqz+fKG84qUtMcuXYn69My3YL4tWcTBGNsdxdpaFjsnoabqcG8bXONZWdj+St
HorzN2V0YnNXVF+HKOgzbl30OlVWq0bZ6uu2Hl1VKS1+mmGWwEJk8UgveBPMiZB0ByRN4t4INPwq
yHEQOdYasdGqXzEr6A1E693TxgwpVN44MKv/HU6YQXEjTIXCOvDqX1hGoEZ+wF+Wq1paciR7u+fM
AP10hOouHL3Mlv96kCKjzLmLoqsJl/nZX/i/H655Oc2d0b0lA7OxfLuK5TI5sBoz6UNsSHgFX8Z2
WF141jlbgjapysF+MIUn5r//5B7NU6FEd1cHVUKWUB8G4imaq0ElHBdgqbcKJAU6Iz5Cz7jJlMd6
xcOMKjLR/yf63UZEP6T1felyfIbV6aVsAafr/ohykwi44EA0vT5ZHgv4imi+5u83O54uUw256oDB
vRqn4QMZmvZojkpWLGMPECmA5yr7Z0ICtODtA5DxxFR9yLWkPXCvC9FwcfpCwngz8oKFkIoS7IY7
XJuUtMVeSlQiLe6I/Q0J4Lcl6tmwV70qT19thF4LkWkVvUOWM0wYyfHO1QMcmjkRCyzEhoZd5aah
9hfZwKZlYBuW2HnPRcl0sHIeMDhZBA8zNav0me3HExdvGjGQgaQ9ci+hQVlyGyopcJMnEYrosUSG
bs8UQPdRFQgnIvM0Hu2Rq9Sze4DM6T1B8ry7ouCHURjiEpLpdXaHkT23Q8AIzsVgcsDK/Qaw0He+
tYfYZtUnZfRdwBi36dwwU23vE6Gg1qoWNCy1Zw7c7/MJDzdFIBYnIiVcqzVjNht6po2kUGG/98ic
0i2XUOopEhpMlqhPj4YLdaoULo/yJsA+Wsxhaal18tNkQX1bkkr2RApmr3PvDeeqhm6EWQYfSrYJ
0YjCc3B+xXFyPMqCWKubgncFmqN3xuNCOdidTo9lNRqBTKTxrj/twguoz9sM+3d9Nr+YwNtwiPi5
5BHhxFIm2pEZJ1cvb8zKwCNI1qHA8rR8WZiOfwWGN8nmiMKshqfrrrwVdEpZ4jmr07JeXlKOoIi5
V6Hn9nT+t/60FUwPrgmwCQhT9n/3cor5vIWakvIUfRKmJTs66Jm0UPXygTXayqOaQ7Gb/age7BUK
IdfQWohDsEctQJ5PnDT5t/tnrBHFdeRYIdeuWLKi4QLyjpyhbKNKDOvVvjg5Dy/ZBalW4AAgdIaE
3zSKi52fG4WEvEqvJU0JCFtEKWMYYB2siM9xIpM4j8SwYamxwSQekUVozSiwTrV+AY4pgOPWBNLf
gLVePEhW0lLQPNOLG7AtlToYIO//aNA6ArBfQD7s8DTJJWDDYJPp26XSD12tP756QJtypn+OODfM
i6O/ESQnB6Puy8xvZzV8t59SYfg1PD0BAxBLQn1zypvCeRTLLuvk4b3RvPf3ThMS4jJ7QDbySbKu
IISW1Fr/488voU34eeemFbR2zRyzMHoUVhaj7nxx2aLEU4qhVgf5WMev9v5vUOMluguOu12rwXep
GpHxPN6u6Bv+5SJQ+MF40XWD8udXoxhn9LSAitbGtsvr3ajgKlNSbzlxIDfL5gsElk3OjG2Sb+RG
tBRvwVpgenqzH0Kerv7f97e7fjoIAmEjYmDBNoCvudRP7I3mVm3/61rLC4+t4RSWlVwdlSUpRizt
H/7xW84PzFtVevxkj2tDi3RCzLbcudNDVYBUQSoO51CXRA55KnR5aY1x4VR0sv4L1FYlU3AzzVF6
5EUYofHnu7b1fCVRaDpjK+IEvBTzDCqSvpbI//6y0JpNmF63gkdh9eBQII4uUCKKCuk1aMFZ9j1X
rKX0Pbt+tErO39JOaVIf5jeQ/jrIFFSkB08ezgxrxdmrOX6+bdz7Yhu4KzUdw/Eft/Y3OgTws8hj
RvGEH1boBDX4a6t3dpgCTYlO2GNmcAxwe5WNQvyRQz9e9vvL3kyYtDKduvpBpCIiTCxGAA2Tpbei
c2It0r3/iQkDwko9fFhNCba153/ioi/FHsIkz0MC6DEMB5HvjdfTOFiZpUUBTWhTD3RSX0xUZTDD
M2krtnOCETpg/ci9BtZOwjTJ4OC+O81Z9UE8L9/0trwnkvRUPkFbA7bf2gyWnGYV+cvgjHyG3/DO
30l0BG91VueCHBbsULIZtucl+pA1U+/pSrbwiBobzCJjw2Es8UpopklyRLIUeVrD5z5XrxZy+mEf
hBfXxrz9Xiw8gupv6SxGqzzPlOxuAv02g9RDCFy/d3oECrkV1linG1+MJlNjcelBdPi23NxL0B+J
0UT416VI1jwZgBAHsiKBkt9/MkF/qE4kfQ2VbGBBgYBOEg22ISA1NpdH6W13h3Xfu6KPAfhlsQjo
/boyDQa4eIliOykktIlgBmRgd2kbPhXXXYS4vcGS7fBlttcxJcmnOCZoumrdOUPtVSCanCB/yncu
Osx4qzRSFrjSuyXX6S9T3cCP9CDG+8XqCZEFmbUbw+3BDyb25a0eYTnxZFghV2b6/k/SP9TjxseW
TAqhftiXgpZuzETvdjUcZhwS0BFjr+WbNR7zpFC4MzptXorFW21FEISMFe8w+dZIz6/d4ZrJErXH
zA6gPORdHxl8ZlzD8HAwD/g6PT89o76Vl3Rhe+8oveaCNXGGRF9lXIztwd8LVhZefGMr0WVP2ZHN
eFbLpcujx2EQgI+e/6jF8ECwx/EQf486dSO5gZdgyDg=
`protect end_protected

