

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PT1CWY3UnkDDUklMeaNBhV6BliNbBJfbhqNG4kOV7Gat9/z6WihgIxC6lRE+3ldfsLvMpYhy8uJ+
25GNPlskPg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UvJJPlyuv70VHT4mYaiqDRKTOeGm/bTLqTJOIy8dhI7h8MQzd+YE6IQThFVGwKNg1149OMGabrJO
oYkVzjNGF4B9Aleco2wvOpKfvWGZDwt0GGcY0bPwCYhgwzblbjwmCgPjWkv54osNVTW8DzqpXiHT
yqTtBlllC+UP6StZLKk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IvSnqjuvUH0Q1DG87naNrsoN4LstR88Fpjj6aMMwh+f6Fho6xAvTtV8qJudD702FeycqdNzlt1ai
QXhCNPnT2uuSCS75+mdCpNaXrbRjxmX/iWoxCnzawaHjNORHnFYbE5ycb12Je0b7xDgqmfK+x/mm
Rr1i9nWC3k0y2ultNBrqag9B7JWz2UiAxNLz9gIhkdjfo9uuq7n44on8tD92VMcRgnjXzhfwsV/R
WQcm7g2SVj3bLFjNpwKO0qkV9egUmW/eEov7KDZj0D4B6HRqmpo2DevGwrEmNSVhbBsv+hYHPySs
vJezY6TBoybQdPcPOmulaKi4zQJv0qMBHUSRhA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
N4Lf2o4qQIsZJ5JVKzqV74g/C10RJITmHA7UkLNDA0jMmd38lQ4sUVhO++1w0lqqkNK7gbVbdw+5
aHqNf15gjyNPjYW1ZhVXHrYiWWCWKhn1CmdTyUXz9OVBdu2lqmPJnjbOZQNbhaspal62bK34xeW5
H7uey4lH4qjMdyRPWyo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WmWXhlbOXU4TrFQt6FbjizC0tiQugH2eLLLRZI3zQRGusS+51Hgzx4mz/p2wkOrjF/inwb9EGctX
9EIb301sFgIc2+iI7RGNXRFy/HDMZa7bViPHFvPX6IIbSblSMhaUsZnDGZ9ShEIypX3t04pywLmp
oC8cxeW8KJ9jku9s++a0XQ670LJrlDd/u67e8zo+xwxrAToVkNJSGwQcgXMc9YDwrXqUemdrJGhD
qf93Ms52+vFz6ikE9Bpwux97WA69cn9Tx5Hhj95T7V3DeqQDYaa0G162sFOeOncPAYjRFsxSNp5b
cwcMCxbjJE/oLyWzhKmrRPek289fPpANZ4f0zQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45744)
`protect data_block
m4EZC2p8pNDCwZZcDpn+mheLKbszTz3s58njsOQ9lQQEbOJIN/HtrfNNHe7L1cern2l15GGH+PN5
M3Cr71VjvOGp4BNZSADmCYSY7OIClQ12St/KovF55Rg7/87BFBrt+D3PJ6rwW6tgvohJxF/fbhvu
lsiRDPk+vFhN1hsoT/n/+G1TRoFhD7k8mCAyuZBNsguOWQsQyXZ5V0yj9LOFfjSU69HVahFU6UR2
9wmyVP6XL/Haeu9b8vZM+gD/mutDkKhflFuT9xpJ6+K6Bu4gOiV/6NaOH7GOwici0PoqahmJm546
LW19ye3avNQcK0p7c5xyDd3MfvUf5e1qkr/CPpXP3ZybT6FI2L4qU5OH4CsKgwicIPLsHOO75hA7
RW6W45q+6pNEVh5B1pxnwaFxJ5sRe/oXe04sdqSKYDnlk3NoM0MaewN3NdieVY/2meuEu7LhCNAr
7H2njcat/Xd3hYP2cVWskZrCBaEEFlTJqagAVvqxCVErujsM98xsXsC1Y9cvdKvsZuN5cik3RgNK
jOzbwIzXNRvE6QoevTw5J5t9hZE5MAs88FGB908aFtBMc5/nAAGe5GxEhOFwA914GvxtJmnxWj0l
EO68yBAhtTrvgOigUBLHZC/al2U1BiAJHxJON7uBLHrGBhA32NPfMtCe+UIXg+CgwD/yVdbOrHha
5uRg3MgsXp1iVtHAS4N9ypKaZHH6xGk8E51GY2zaUAexgC5uXSIcHftL9G3AAUEho1tfUo8LNNiY
xrEK5DJJmGK6+1REKknCYZ8TxcrnCRXL9J06FQyJB+vyk0nJsj//03c2WeWkz4ZQiDmPeRrUNqAg
p+bLzoUH9OxyUORHlIIp9wCB7Y1KElCX/A899n+RLSzqtKYYXwM6vzF/Flb9imSYuhOAHwBHd+lg
Gl1APawEox0A6aIbbG2a0wpgQK11Wp48XcYlrUJChAgNkiTXHa3OA4fL51r1/nn9G43fWfFeAZJ/
NVCQeLYD/upOOJEukU0KzCYW9COMi4cFfT0K0Xhy0VXTxnk1n6+EomERxADDByt2VZOpFu2XM98T
xJvLqS6BwOzSeafwhFHb5CyBp3+/rwEUAqKwtOkv8vVHYT769qD5fp4O4zDFe5aQn0s/lQbHSpN2
zjcOw23XHrhSZfm6ba9wORdlJ1SUfgtESr1ggXUW6ZCkFtVwtKhwV18815Go+HBhBCaLzMHbQyRK
gVUALmjeqC4ujp8w1posLS7p1bXRVeLfCi3PVTLlQ5YKrOp6n71hV/Prvd6KkhZnFlXLar46N9qJ
IvYWBNnnmz0ak23xj8MdQjUdYWV46tR1wUNGUX5U7Swg+xAx88iLUzjOHuX9rvb0UVOWZJqXZz49
GW01zuIzxTVknUgpdwcmIMF2e2viJ4rWuEl7/QnD31XxtFW3Jmr4Q9f5lRjnN3AoslG2tgAC+QkT
k+4qcWWzFx0bpHtUA/sYZdu/bEg3aJsYbmCxambkL1HG7VA6anw6257nJWRvs/7N0dQH3eDWT4Fl
xoK6DfWs7yIPm8ppRpdDTdmn5GRwK+b5JY7rmnFnOKxUzrFIP1mcaVdu9oAlmUpFaZM3DF4IJrGl
Ejug0tNfnVHFLUrRveSZNhp9BCxLzZsBPahGcN4OPZ3G/LIjjX5sPqFxqNrlqL7sHDeIz1oHvsdP
i13y+WpDRFV0F6G+pZaUtFQoz++rRU+aVzr1avYGAEHuAPUqmoiyxV9cYHJcCw2X83pEuAoIWJEC
+pHas1DP/ryeab9u8twp7ACJpkXxUeConYG4EhLcQguh0p638rHcX0oUFd2rSqmzGdhkaWP6yF/Y
Z857qfP+fvP+B8J4n2w0rVHDTcBr54J87hJnDM7yG8GZh1WzvQOdURtyG4sRQTdmTycj2L/rya16
jUi2qK6T3Wh2guoa+WXfDaPbuDAl7asEuxM/zjWgcQAwKqZrD7OFS9Wnq1Pm6Cbh7ubDEEtTdLmC
xHAl0hsh2rt6i9AxualPP6cMZZCTL/6eSmsCubn1yGnIHmse1Y/GXheq/DjHaAVuVhl6YOt3wcOu
wsXOSR20JYLD/Lw7H99Mg6NJeu5ETZe3YLu4dFnsR50jxXHcNVMG8M6/VrgVeIlhGnJPj5rEX9Zy
KhOc/EaWsTbcwYk+eTps7HBoXK7IHOFqwyPnhCKDjTo1yEFGbHbay85jESaEJrCE1phhaQejfx6T
YjilWCa0nuEtmLlTGBksxqPLb502ocBZPCiZo5wr2CcnwhCY9Ypjw8QTiKrjlyn3O5DYHXR2e12n
YR1JAtR9pMCi6bcG2AMSmP4WiqLlRVwI5O0d+b0S6eFE9Z3JG36uf68MH5vQk5TZh/++V2sHYrKh
CLfUiz+StYbROwcRvbpv1QuWktUcxp5b8LXcD0atXvoTnsarNrriLM5MShrZ/Grz6XaTvbl0ykew
caN+tHqU8361LiNDmFKuPvIHPjVVq0ktrOmjY1dcKO9MIuFT6oDe4ac7PjDzXk5sTYeQ6qJoX3U6
sbprDP6G+peF9GYDuDGFXHup7doSa0N3w1gywoMT3Tg6t6DPapz28FfAh9CTYoXDJuGLz/cpg6rP
WSbwrNPLnLycqZVDDcSouR6oZw3PbG9zVp8siE53FPsEWEoEmn5DmA5kElvRbnhYBj2V9YSRWL0S
FqLPUUc26MKKZoKsWfm+wfAFOh0TcmAw9w/62/xSzGRT/K8O2JZw/rFAxTW8WGfY5BWq7rURll1x
1B0ekxGXR9/VNPq99ll1UFcIXNqgdE5jkHRT4JM5yRcEnC4ul8koRamrq/a0Ig+gkt7jzatPS/tX
mI6p4uXkQtEXQnU/OLA6WFt7hyW/VF5EeKDli/yfF0BbLdhImn/IQqoiLGV7P+qxXl5I7j0pkb+t
65AK4lHt3D+5FV+pxYxI1WMTjdchuMv/yE9OnlTtlVCeZ772GZUvXbIHwQbz9X0pqKYkvMv166Pc
TImdE8vup1dutIoPy/2bxewXalwJjj/IhYex6vN1aDg8tMCcVkWUH9kmLzuwxXa63Kgs7J9vVUk0
QkcT3Vf394SRgrKJRXZibD82xxkqomMSfBnVY+jNqXAbmf7css2ezbGnVcWEUdabFeGnGdHgT9az
w9utOe6ObIZyNqL3WnJ364wjGmXzcg+x2h7DpdFtc2jcC4/tp/hFQuOdGyuFPd0g7jnAKGcG/nCH
ackKhykWK79zPGORdO0DvWsdcD2dcnGJYhwzyKUUu2SRMRI6PqoepTBtoKPqcTyXm+BNT9VTZ+o0
RhPqox9JRfVUhsy/QSaSQRiNMt/WZdgoS/zXwFNGvy1eovgZ13T9TCpf/d1CqhJ63eft4xDjM/UB
ERXKQdKQRKwYOfyIx3fhJIkaE7yXQPxRzwOnUDyiIHSyJknSfebELaLOdVjAxq+AxHpMXDiiE4DN
RQFR1R+I2oDdUaNLK36vy6whGTmOougnZvmetagPFOQgiBWBswAiuY9ZnxQunKJWPUE5tXytGfQW
ms6WHz/yXLXBgm5GW2lgnlwupnqErFpLen9sVBvF8UqHeINPDfzQTV/0jAe2/2Aasvkv0PejWR/Y
ya0VpPVdepmWT4CEzZiuiNcSucGsT/Ks2QGaQR5960/S+1WTt3UH7mFhiRVh1uS9hu++szJi6v+C
u6ErkYOn+AUIcFdY7/+9LDXB02gfC6+iW/UMeomUurmQBDoMuoDD9qK33X4WnHlVgqPoQu/v7xEG
s+IzofRQytGW140BJ/KExscdqTQAH10qoQTo7DvvUEbRrC2Y5GmnfhoIdqr5iKogaFNowVv5meoR
MpYRXsWc19b40MvQSCf3MssXxaDb6tYUSofsNcqzzRpgQdlrg5smmz7442ZxrQSu4TWNFGnXFzu7
1WMqxt1ywGzI6059E3Q8LKbXnA7Ze1PYooRBae+AzDKPTdLCuRPPv3RrKyfDX782i43jMW7QZHs5
msw0pTfjV9BaJdnXL1+Jpk+JlhN6DFsiaNSupftUhnI9PCLfkJNG4AslhdQUMO+7kDZOd1YqZRBx
B31gCy2vx1XwXvT5e8d/PICTHOOqoRITt6fYyTAc47TU4IyqI/mb2zXpG7yB8sWlS4lTnjTLR+rY
g5u/9PlWLGBMP8LLFXHJAzKXlt8hv3/ufaYd4bDhjBrIXOg67be/5LJ7c1rVowOUL3+VPY1aaqtr
3JXDtj2d/aWLhCv17t6DjAq4jJYb+siEUu/hWSCmuxzmNBFWZzISQi+xRKcAGZhdx74b5Uporija
RWjw8Yt2fLaQMMVU3t9AUzGLj/XCzeamFYyFfuB76a/4CFz4ZiIC+MRmbWlev/tDWu9BN9FphovY
AyNMm20Ebdy/MgmE7HldGJoJhkQd6e5wygZxCuNQXxfhTF6h9bZ0DWoMcHKcXCol6NC0hizAzwrQ
3Bybjkzytbe4m/d8+LJhYVatnXzbKEd2P0HljdAkdrsKmDyt9uMgnG7rwip7qdtCsj3r4Dg/8P8O
MjCNQnVhnrs5or2qMwSS0x05uvqFN7K9iYX2uK9nLomIVvp6Q9oKfeV4WvrU6GyXLtQ7MmSEztI+
W4h6M6s4fWItjrIiHZeSZ5+iM/vG3FI8e3qh8UnFIfL3bXcl679mbaaVWhXCWrHclgwmMQaRX2wm
UxaL6Fo+witLnbzTPYUrjfgENZUqsSksH1r5dlJBQ80Z6uEi5n/5qHj7cBRSOfzFbJVEx1ifmfP8
yCABmoj8BQOP5qHbaYc4CE3ySK1wrwqbg81m2JvuIQjlBN6D2+bD3HjmEBCTD/gkBYM45wG07GYS
kiCgyRNHBIMwgsGHT4DPDMtefdZ4g/U/46xu1R2GSYBrXwfEM8Wc2xt0Cp6B8/qgbYZYDyBXpPgK
vLMI5/VLB2mDRElROZywVPYw95Ux3Tn+xQbwtRI8A0RXNkF9UruvDm94NBftL2oaRX+fQyRdkb0G
4meto6DpJAsRNMvCHc2jYBjEgf83OMBzcPgUExKmZq7qO9kwikLc0spn6jihk4IBqgiJoUkvUwVy
HtUfmPZ/cR8a285TalveauASXnBm43R8h7I9GDzbBKElTH2Kd2uBAJXUG64Hhw7J5lCPD0IfoT4D
wnzMc7O98MhuvwIAsRak7CuzrUrOqiT16CwqKpskS8XIUF8lZWFVLgFR13Hlks8CKlYl/qF7rvvB
8+C3sSXJlMFafqi8j3CKNTLKZcQNv8n/XmMxsRq/j+Fw0KsHwDLMvRxB0FPWIAmpFTDoDpBxPlLm
/XprhhyJRZt3FmPsFbN2+f9PHgt5UXbKLSD81Rs4klF9mxC5eeOgjJj/dhiWxZR7VQUwJ/DsOIOp
2/eh8zap9Z+T2VZARZ4nUC5KW241iNGoVyiGC6leUgHEn/q0CuM5xe7XNf8WbPkLAPE2k8bpSYMU
xwvhHXA2xhVlv0hBw860K8kYXp3jC0A69kEJ0dbUiGtzQYf1XnipV5UY1X9gCxMhjl0MFYrLEi3x
D8TKnPEejIV8RWjL3EkKup6FHHgKiMpRHIfXBl7uN5WIqXUKsou0Efv2LvcFuCNEI0dMVSBXmwzM
iWuFhNUSFU+QPfFEuQFCqGzOvdYaLEYKd3xWDLRDAPm6dQXHHyXe/UBKfnLltoHc854GAOiXFHYr
XtehcKFIuf7DVm6QSJsX1GytuPSmaY2Nj191IpijXzUpBovic24Gv7WT94XtsMr5b4HdIrnUlEBE
RXBrMJt4MCsjzQ+dn8DqjYUCfBjHfpp6Kw1uCWJxP/io7gSWSmuGfUACYqdoZ/U4BtuHSq29xpur
cYqEsgKKQnFuVMOtkTIhfxjldjMBERHuNLQTuE9bf1OJtfxiL3tEtT2U6FvmRzV79TdsjQvjBho9
T9Kbf7hB0x31oZrFO+89O3PD6Bn1hwOi4/Mz1gsqRV3+23fxMUAKNJ+00fHyNB42r4AuZhhyf5kJ
g+VQoblLOtbZrzbml8yYmI3ahfOd85taVkaIsIBKbk7DTytCdsOtnuE+OBtZqa3LK5Gx1zE0SKBR
M52gJsYrv7QDXYeuN/cEjdzIO1mCbKKqnJpLmcZ+qBTKt0C1hdsNRvuEjpsjOTztyj+el3vNeY0d
zeQbH8Lz0GJsb6uR1cqHOlF8t+0w4S8+imjeTZotjzGig4YdX8icvSF4P2Me9BNqXsxO40CIIJur
OLavjEnIogOT+8w3MjUdcpz1J8MEIzrTnNOymZLJvGLHHj8yxrfdJHsQAYbpQFkG5oezf7LcUNx/
53F+LUFq/fa0sm38S4hzD0P7cQOn0hnxRc33cGqoK1TSwN9gpNEMsnNpgS+kqdWP/q4tJMsxCavP
fQ5NQw11JPqGFb+Oy+wHv99Hy49ZCt4iu2L94s0njXLrvYk0kU3uwj0S1JcEYvxotbfiGp9RAQ2X
lnABMSXDf92+zQ89rDXD/S29I/Ui8BTpDkIzEfg1sVkSQy5jNMuDqYeBn4d/rxoR7Cykyx9gZO9o
YSJjx4QiQmO/xWuSFgZ7EvH06vIeqepxZkvNSKpRDU0tf5e/8a4HKumrwRuRrAqj1/vdxbyNIoIx
lMnsRYHiN8IH5MqP1761wnO7MQCgmxFol5zVs4Ecsay0IpVRstlVpWWdDX7lyuG4KqUZuFF4S8GH
YxWEli/SNuUZZBGX/C1iDriGw2QIRawjpnegeJjY2MapUubWMo2w+x8ijuufgrPq2ArJ8e8z2uNy
QHNiQC+cOGMil4IDmInqxuNFYDNQcQDfbPqBNe7d7Sl3jZNkTByv3hvyT2YXCSpjgoK9F+WZL/yD
MaUPi5dKj9zeJaOcLZzfyUrDSGWKwKwbjYA86baOzoGxzWQfazz5/XvW5jdKgo5fLozoiweyLFqx
546awayFKwtNCzCHv006dEmW3mU/6gGzLi2d/W01dQARFgBuodQHS025CE7F6yBmtbRT9lsBp9TE
JrPhmQV9nxHWCR9BGOzOtVHfc6Qw67WvgobCvHNIpQyUFxlE/DR2PZuh3BJNHIhQAtsOJb7BjHQU
HGomNKJ1zOSnkPHGqGlqjz8Qw0Y/fHYifexf6SGKStrD004xQrrGDOSIbYNw/HNPkcJ2DJ7AsS6o
8q6Z3x+7nIEtCtMtH3Yr3pJZp6LDZUbV9vevzOV0IrSRegEQqcE/tFAHciqdntPzO5yFxSllWF8z
Xvs4ZJ+51ZkS4+nY0JouHahBizZ70girrNJKq0rsmlkXvHgTHLLyRdfD/sCD7bZgX3J33K8kMdRk
hn7MeQ6vpjezY/BXjmg+5hCWu6joFKsPqPUG5Argxz47n9aQAOnIMTJ8m1HDjdY7tFMEIaNQ/Spq
WnfcUikWtPFr4YTd1ZTW1Dh/x7GAEQUylb15J7z1oqfwrcq2JZUo5s9buzbyCHEd1Na+QqL0Wkue
8LtqkjXBF+CFh2+m9c+MViUEN9NCsLNOfDhI4gN+vz/rMCSvvLJz/1CwThuEmmFXGGHrASSzcA/b
vVGeANCyMhETGAyygRc+C3nvuTr1fT9Gl85tOhFl9c8J/5NMTA1wjfA1dYUO7lNgT7l56vBHLN2c
T1clzv6jPGWC4E/hyVgmZ4sKEZoJC7xT0btb4LSeV7tqYcdU/eKZHx0zHMd3q5M2hRXMTJoKh4Zv
B8dcU7qT1jDvG6fCEvTe4eLti/W5RMo587728DwOIkCL2giCYaV3fDOBk1lenDVTBplW2Js98MiF
gmW8m7UBjD6+CB+PJ9vZed8AFXiWH02fO6wPOey7iqh1XIuPmU8Fip2ejEHSF/YMcOCwXn339bu1
xIv5/cbxsVEG1+Px1PPEcphc21S1IYc1z/rMfTjKz+oAHumNSnAY/dKQ38pPF8wu8QSMM/8hyN30
sDFsNRu/tGUnijC2lEsMeGStlMBzgD2bd9gzyGyG8UCInziBPFOFN7QJ5IW7oxUJLAJmlS4wXLbW
CBm7ex+p/QszWtVyLnTtppoANd85hML6oWop+tPMjqFY87p2jQb6gBtwYvFXuUTv4NV2K0eFqEL9
m/eRktmJ5V/yoIdTfdn43mHSJ9RCMhV6kmj9XHttfJS8HEvGU113HVE/FRmohhOOw46IHuMEvhfD
PJ4UNIXaD1pZvPbpLqwke9+IId41Sa3qWVkcGC5MeKyXyyQummxzUMZOsc4h4Tn48+Spl7+zxI8j
Oj6H1TRZYmm1+CEz8+Zvpw/IrSg7oW4/EiWoD65yAnbW72Xh+AbCtJ3/sbQlckAAtyWoOHTlxq7t
otDlOg+nP7XPEPJIxLAsBXQmO3XKjc9esjobd5pEa+kBKGvW8VHnW5ZxGEOLvv0E9eBGAmu8C7AK
7Q6qaQylQUD9pffdKtRvOVeMnjq3+f5+hLFe4Iw+X0dAkYScZx3tzlFWjlNffMM71GvQYJRNSDgw
YV9a/pWnFEDkl30WwsVyTbct+ef9NPe5DnaBuUaRq/mrUXRSKy2InjHw1w/qglCKyVH3R6NqDtRV
MW6vjr+5FXuje/5HYsc4eE5o+xbmqnG7m4Bgzq5CgON7oPoOoEFM11ihWLvtwg774yG5be7Ba/QC
ECUylRQxYr28bfIRx8SnpACZtY2wZ33qzFMqmLf+3aBSxvS+IEucniQJblTtie9n6LIMq1CRIG7Z
HM0DHregLDOkcqA15/R1hu714Q6rOzBIkoUCwJ8A/pdi561rMGr0SmE0JktPFuU712F4/OQAi6b0
0vb6V/KNJ9Vjg56DClwzURSOL9IlFLcHP1FFa06j5+gOGzI/lyHA5O4xd1HU8UqHPLZfGVuOnIGn
lKPiHXlTqofCN8ZEhQ5eyxOUj0XohdpjwwuvYaiTQUU0ivHpt2BiZDMl+8KLSE9K3pdE044DEbxP
IqxTCixTTxXP4nDGv8x0w8Czo1tOcqOKSS8FfElSXBURcLJsKJ1EQE87TZUW5YCKR77ivMLgP9EA
oNtT3+shjbGiAuJrX4llITXd8YbfKbPdLUkpYxhOArsZNJ4cH+Rc6E1NOykyyOxcMK3nCRpEQMBe
Ok88Cj+SastYam8TKSdsQzJyMp2tRaGwNL6AvJKRZAdh2I6OLIZHPhzcuYYk6aNu8cgvbEBKAG2K
bhA326Dl5FkBVAHncL0zEz/QGmqLi7g8lThp+wyPic7F+icIedrvMg4RwClmeMb6rb7EfK8fws0S
Oh2H/vx0o6VHp8+HD5ePqFjETGKo+iImpgYpW62QR8dYXheoe22lJbk4KXsLWTUH2y6VC/7dOKMz
OToWvBM8YdbFUYHBNFEkMZgWJi7gn9wxygFbSs4MhJcwcWETkVht2NuprUHBiQQASmCjyBbMlyo+
uqZjxSUBrotamXdjKPZ+tH5hbryaxaqgs3bnaeBl8yI7WbAdAaWwVcQoTamQgS8SvA1IULpwrdPS
jPt9M5BvyDiQSxMDOR8BKhwHnNGqdEHLlHZ6oMtua3R7+PuGjCl4Kk+5EZfCbc9YRxGlGWb3xQYx
thmke5mfxoj5ZtqAMmsPTKrJg7WxduYrZlIWy/X69O0IvONzq8pHH1eOEl3h0jUxMP/BBlWPpiGR
XvhHFdzzHoLR5ZXrN3h6qJpluCP9X+RhE2CrzMpXvk2xbbJFkRe5+tUkDEiHE2BSokwUSaoYBYPU
lAW43De1bqXJoE5QpIiImkrUNcB5Ydyg+LqD17uz3jxuhpxQGxglIPzLZ24OTd9D+QeSKM7Gy1js
TOebg05/fVgxi2Pc8D+ZcZ5oHLpIwx5UF1PIcI1TkrOJu6L9p2w8fnE4MMszhKeDIklKNnlng5Hn
hoNPRg09DNgq9B9EYQ2Icr0lqndOlPFPCdh5xywnwJDpajEBglwdMuIoVlkXgiTkxdzUf5us9WU0
lub8qiYal5K5z1+sXuRA0Cr/CiEHulGJCmmLJxNjW07SGk1r1Wj15FOsjVIN3LyYOmbillMlHbRE
nU2ODeNw8Xe8l8bXFqA2BN9MsmJcZsOywTm3RnhqiUVHOiAbmvVrakBfkMpEsFKPDMujQHwNJeWl
j1o/CFR6YZkTJrXWd6MQ0v5uJ3qqw71Q3O3umDMJlU1Kx+6flDkIkH+OJ3Ookx8UpxAeW87QcBIZ
TD1ViN450k1OwKrFl5ydQBmcIIpR6YlPF93m/ds7V4Pjm+8hkCGQt8ioCyOiJ1V3CP9q/Yl1lWNS
AmqOh5i9EDaIQv94qoFe8X9rfnZSH7jHT3/E/zTVY4PQjU4sS+pVd8ZC/IdwKzFcq0yZAOalfjPe
671oBZI2IriijEdXnpTL3vo0cbZ+W2HmNeCLov9dAOQndSjafmzq4M7jJMKg1mF6TigUbhGa+DlT
nU6wjsjeG7YRGq6ldha6H1qlpu39h5nQ9l6pjfLtrDdIc13bRyXbaZBtZzApqVubzisgWkmLocz0
jVLh3WkDKbway0+P5AHsy3BmFhxNMagsqfIZIzDDh7xOGrG0XinSjVlqHCGRK5gdpijg369qGIH2
OX4uFUbSxv2wGzt6QFd5jFEcE97PPSUvzQ3QGOy1bVVx3cnErr1RoGBABmJ0WBVbKTlhfm/Ft14g
yo9a5jQo6QKK4/wb3RhUMXjMfabqL/yrl++1V0JFH7dWeK0KQrRKTAeFBbauif7Ups6qcm+J3ulE
S+oAGfPVgw7g7/sf6qQhe56A6Irgeu+1+GqwO44/KMyVrOUiKGVWEhk2K+mu83UYx2V4M06wYTv/
u32ZMdo7qj9Nizc08mtYFmcMTRoDIliBaqJhESN65PYZzzF+tuu/4r6cPF29w10S4uk5GbLT3JTn
7uUSKe4RaatCb6jW1L78RPX/IjOQPCPaya7qQYfdnfj5USfcpe3hLZY80HpsC4tDBw/Y0qZaXTyg
ojhPCY+ImxdhjssR0hljtf8UbC8xGOSq4M5fPO/LYkmWUECtMAw5sALdSyuvli/KWBUXRM28dwm7
wN4xgzCRNU6wjr63bf+nTley3+OaF7O7teelppHAUhIKa95ViYgPAsj2DLLoYtF53kaOSwG8VZXh
GP1NU/LgHdU1AWjQlEJ5EkJSmqQGi84xpTj8PI0ZAxMOgeTNAIG9k9Rbt2MAN21tBeu01cTcXHUt
LfHqz0YJL/xru8Jy0NwFWSMRQqY4eFtaCVc6zYqxx6KNXAO9Q9Rt+GWHyZxNKiWIQxoyDIt/2FG2
Xz2Qhc/eeDZfB5Jh/5i8M/6gLqQLc/0f9KTj9ojfgHK4DDT+9jCcmSfvoseRK2iTOAiDQxG2VzTh
U3v49I999Zq1uMsmdHwJH0gvHXgmWG0SS+Egf2J85Vub/jJbsCyBcUUE4Mk0u2BqC6WRXYzlxkl8
lHiBTZepFkXDsBqlzZ9/I0d0g6C8wlHDGb/RZ/anb4bEImjCWn+sTqn8dzu/Zyju4HwqHQJBNcF6
ouKA6ovL6WNjy6pcTBAE5hxpDeTCuMha2o6FXidI/++sJLhLLhjcmB/Dk91zayNV3fPTodEN2uhU
OuNm0ouo+ddwgYsBbwjwZMNnAceE79XpE7cLcQFsR1UzJcgPcRMQ5pm9xj/ZQ/yESgFoS1mbuUOx
RmdGFJCO7mPzwuCDPFpYC24UHendRhzv524GisTlEf6gL7klSxi7CNwfw/wZD9LOyiR9X6JcAzdL
zh+QrHK4csdipT35YzwF17edwrjcfbKFP2wrGMcPx7pgWwAwCR9N763V+SviBbNLhCHtBCmGpjaR
rIkNpJ5GzZyCG8awsv9+n+pTh57zaC9nY/W97dNlu25iUjlx5894qxAigQKTOF4EpgSJBJ/WGnv7
VFmyFIb1/ZUJjTjo1ZWTGySZWIxKEuvFSDLuKpGJIyWio+itNNmywC+4GnT69D44MRCsCf0KKZFV
slpAOOVtwn+wiKLV1lFA+rQinhVPJKzssv7fIRHThmpoiQSv0MrNY8G9wZwjfNycQoiE4JoICqda
7niXnj9agsywWFjyH5FiSFXm+pMO6TD7q5yVXqbdeRCQzyNg+hSFZyBHu2t+d23FZ1qKmI1j5Vy1
QpyCElDXuUGvyk+9kB1811e/Rx+/sgpgHgEOtxTG2P91CeY7Miza+GWxDGiltOc9/wsitwNekuiH
YlNJPoJ0lGPB/1dc0yv7sN24FMW67btrPnwGeFAd3xdzEQZScO1Jt1YzkpKFbJyEkp8x3ZNwVf2f
nEurbQRKBtbgC0Md2vU7u649hacZVLFyMZ02p0spSkete2N3bHeqEAjFlQcoNko908WO7+kQTblm
DZfcHO16I/TBK7/g24xTSsWGyhyjHEoCQpdtd1y8kY1SIkUzHOxoMeyiYL4hoj9R87siKSZVG5VI
bE1l+xBYvfAyHGzua6YXBZDMr7vxcHJ6TL+e6c1DKou386hwUoGnMcJOKT13ZwKwcbPXdA98bn/z
bl5lcpqCM/CV05xu9VxwEVI44u32ExeKtrltgXpI5KzdUmSSsOhLgS3/7LfHtvPYT98X0mhdXL2I
RswmSrwkEAtFyMBL834MtHdB5yQRoUq+XdcC4e+Hi4edc7BeMsB4x+OYB/VhdGvEOOOSPoGmNOFx
53fqYa6/FlDcVXXbt/DNFm8GnlVGz0WgllF7JERJ1RQeLbFYrVa3HVNDcTz1cD3cAGbcsnSKNrgD
z2+T7ckZ1T/YHVCVpo0xy4ru4EButcP/SYTF/RONwgiNYAL7/y7a7Y+9SaITkol/BwcaMiUbXmUU
1fWGBqGGb2wgpN+GIC8S5QcQDlQJUh2yUTNO6YyMRkNA0fKUTq7p/SzPyYHdlVji6SUA4tkjjb0E
e7sbRFim0d+ZnIP58/FRr5TFlsFDkYGw1FGPMpsK+2bnMx6S4LV/YdQ6eeo35+phprO9AlOIg9Mt
UbJ/XFmpxymbY6HQQTeoa3lwRk4OwRAgMkEmX3pM419G7A18j1t6riWyQyeUEpKnG3fzFW8FLHWY
J5jqb9CGvXGNFy5SrYobZx97VU59DaZFAgyAfVnPXMKEi/gAR34hBSPQNYrQF5Yh64LBpX459xkN
pO+AmMg2d0bmky9N0/X+LareNzurN9AewpVXErW9gzZRqZMbbn0QKe1IhSjZe00JfeYUASsMztbo
r8bydDuKNNQunlFl8mS7cKoAKprYT8ZLJ1cwfAfZledKJIQDbvCTI61qJoHO6XoUCVkNg5958J1Y
v0N4KJ3alqkXfPlf0B+6buonN0XutZF4weuoSgk4vLWnIyVmMOuFddB448EqiWZdOw75Pm1+/jH3
6WMq1mZ0vwkHz4ly475eAfjKTgiPzD1YEheeyxZlvib7kydju3ayHsQYeUfWA2mLZHWEx09qTURc
UqUeNp6oqCDMU5nhbv0bDGhW+qGk1LrfGiofWTsY8h0eLhBJCN+OpKU8fbUJ//7QER5mg5dYOrP9
zjp9+sixWhnh1lm0XIuWAis/M3ciepDjocSGlaE1CZfZzta0IY1Hzv3eDAjw+cCPXyMrCpKWJyJL
Z/6esMWXBjYSnhh69edz7LSfUrnmJIw7vVsooxLROS8lKv7pW/O30O3LlVDgK6c7BHoMTvGSEejO
QVDBjtKBFkPxqlrPlZleiKMeCu4yPblT5dFaTRnvcoK27DIgkYD4bGnInR8Tvnd4xbsUvdYf8Oq0
97mY+E7QuueKrANg0Cc72WW/2EnZGWe2U4Fd7/z8qGrdmlWvABR5yiAYsiysVBbKL5f8ShOx/zWw
u080Z+ibS/QBQbQEkt+x9WVICsrU2yGsWshIaMeMsk7siTkzIAsfhniOfshXjawWiaIvEUKRgdK2
ruacvR/a3Hovea/cZrUgGqdCbj4CbQ2DBzNn5w1h/zzYI975Q3KHxqyQ+1pJaMi4MfRQHP8rPaCJ
klRC1C0O2VlypaqcpGKdJACvKarMtUYoaRaHdVuJ/2uCEt7FuJ3ssbELXgbbrhy/uMoLUa2Ky/3+
poblEBo7ghCLkNTWPqJVeGvxm5Gc+N9X5z5UsPDVVpIbnkPY+RxSIeagIV1F34YmqtX5NO2rX5E6
AHjektJ/4lxCyv4Y/n4MBBcQ3wL1eqfwPkCUyw1gbmy2ryikG0QfQ8Iqej0OIcoro/ACx/XRzVh0
YaL4oD1h0aZl25Wjs50w5LG/Xv23ETafWmXxqOb0f+pez9INEVEp3kYh6t6wwslc4UidivuBBUMa
Qr+5KzvrCA9n1hIjGQbwWAMWy2tew8gruOwZg5UyrcUQZog4f+RoxvacvPerTMNpM9+chYFfvN8q
LTz0Rq75DAjy9kjwRSbDKZJbgtydt8Yz+JxndqdVjMX5/PkhD2T4tX5ApfPr4+pVl7wvgl86fXNE
3vUYhlp3jdqi+MuTzEVPGmNYmbxW5eBl380RLUSpNM/L55g0i1o35Nd5pIWISATHikfCOk93SGxb
ouEkekstw7pYE9XnnorKUgFSGqFJqF8UHUua3yl3GGVJndpkl5sFRkvHPCGjxvYNicAZHsuANqZf
H15ckOD2howq8dN+IzbBYk1DwDxaqzMggxFLZLuq/vx3gEPso0KOIbIbSMZDktS59x2ojIwq9AG4
BASxfBmPtjjoWX7SkuZDZcSZkCghEOfblPbheVWfk3Hwfcw8pz0RHz6qd1i8bgS8d9WAvweQm+5w
Bn+ZNAVKXNcSdeES1FaUcbOJ1/tLvgtvex2xh04149i+Hqy6lSnfWf+e8KjVe09L4ADIj36eCrKS
mF7BhkS9XW+slu0hQ4VpwL98PhuiCPuKtJPWvoH7sILciteIVOd/05IohqnDR5iKicvNnlWp9v+q
wTZgucTxd5vhBEG5Brea6VcSYGieKiqyj3sHyd0rYekVra8okTL924NtVW4rYd2Fnpxgu37MAPaM
KRIWEWJmRmZ0aB7ndJu/Om38/SdOFJ6X51t434JBgNt441Tn8o37UeGUBzHB5hB0IV2/3sGSVEaL
TnsrgxAQEaB2pwhk2ADR0tjbww9v6K2ucBAXcBBxM9k/maakJkRFaSIPVFs1SXiiKLKrm8Zt0hDp
4/Au4gQ6108yoU9+S0qhqxxcko3PlQV0wtSYkP445itQbhH+YDF2kH/PelL2qW9x4BK/3wqmv5zR
OCjdaAq2ZixlPoMnJ6pm7FiVgNuMhn3KtRujsc1FlbojNGJalQ79u8tTKiJ7HmmvuiuhORZKsutX
8zW9F1X0KPVadbzmFefq9f+FwE1xK5twL/dKm2veTpgDQAQD4vt1SPRm0Y6Yjh07x1gJnPS40sTW
KA0+t5ohOoevsdoHlqqoNcQ6tb1iH09VZ6WVNKOIQ9CfbK4Kn2uqdGYMm3BNY8eEpFxIC6tSxJ+3
QNZhlrsaT7pTcrZjIHh2kZun+mwj9JFJNz2qxrcufi9OtrNTS82uzZE3a5aLi3e+9wflZ5qjqycA
7yP4CCGRyGCJKXhhQhAa9WEE3SMAWHwCw5UrGXiekbAD/wh/l///WQmjnhVqK2Y5otj9sJYXyz0Q
v1EblxU5ecEgyx0IGHlKKIFEShjBzpa62jQfKSIPqJ0NFITqfVi+VoIFoS5ZTE+fUDwAdoNwLQ7d
w7riHor/6lfQjVyM+jvE3/c5hmbpg8unFG5EaNbv/iExKzyCeqPpXixYccWJHro4rLDssjENNoOK
nkmvOIs1rv0bRh+6r290OSxqmyJC4P5hOMmCKNimqJ3uycLr6o5ELLpAyc4G/Ri8sRczL1qSwX8V
Pb7MgGRVvpGu/SYCjS2ePh3IfEiqfOrza6bQSZrrrBvv2bM+mLLYqOsFhXVp7b+qyHbuu5hRqEBo
ZrNO6tFiTDg2n0+uO6a1yHuwZsKfg74dsEnwTACGKT2mKn3DT8sjMvpaUUTyabIJwWTY4onDfpMq
heQT4PCtJBwzXii8Uen0ApaabkcxMdqzUjyYFJWKz8cFhSoV/Xu1S3O3T9EGV83QcFM3o1OpyoeB
+BHayUsIZggUJqSWTrz5qCm92T7uwmZl8EfEi2o51KNh194sEkuCSgdxoB0pSTwBxnpqvvWqRLC+
FmNWfn4Lue7Y2mbz6Rb/uaS7kRVy3lDs82zuMH2QQU5lvav43l2mdhI10UDqvzgoVqyZ+1j9UB+j
br81yOdyCrC92vAKfyeNKK0ugJOZR/dMOfMu+xhocBvlsn0rPLE/fey0IHAQ+hxe2Bs3rJhGz8Z4
O/Fsk5eqmwgyk9ydsreFTLT0evGFqy0GgD5M4W5jvNWeIayy5Tbk4fnzoHFu1u+hs/BhUbWmzEBn
AxxyHKFo0q5tKgETSpNCKuRFZkV7OSlpS96a4qgMQswnCIFoYUAHWupDCPXPiTeSvv3HKjdHwisS
1EFf7EcnzYRgyIiNoCfHGxnOVRNpci/WyqlVwbnnle6KWTZMVMLXsGHQViHlEBmMNsgoz0W0cFIq
p3aY3QwOo23JfE8hV/gw/MZIlhBLjEDDKFnz2E1qMr37bNAYYN1PFhqiLVoX95DxueTtc0ORljXL
IuzrQ5GkMamTypaQ40NcLyqSn+NTw6ZmD4QOn9uPAvkZjqczMlxAXisXok6ICWaQTvwsH3hy/uC5
ySmEN8K7tA0FFwLlIG/Szon7Zsd7id8O6w039vIpW/A5yuyBI/sjGJIVgraPSloDYY+FA7f6m4s6
bFhcm20k8YYaSuE41gsfY4LjufLXgDhndKQc/mjkmL/up0AqJqFRkN6gd6ZLI9F40bBYJW7ToDry
HjI2uFdXrx/Caej8LzxR8l5fMPfQTvBFnvc8FhuqjItD9+3VfELFgaaBPs80lPl6zBPqjPmd1yjC
UbkmRNYXYXxgkYflRe4e3K+vakw5nvq8D0MFYSJAIt+9/aCEjHB17ofG/SgACrnRGhGbD9aQkj4k
WBE44ztJ2hYhX/4R8Bcumkd3BFheRbtuFiU4wW3reFSiKa7Neh+FkSjhjBwH9qmMusn4yuPrrvhq
raaLyMjUJ88599UszktyxJ4bxsN2nmDH4tFN5Iy4eIiy+w77WSxQAiYqu0aoGo0A1Ad58EggBWhp
0xMpUyI9tAVLCRyTF93YnDyZgBZW2Rey3g1d+dB4Gq948yPRt8maDxHrZvm+ABkReiADv3YdavOV
ONMI+w23cvj8wDef1cTOBm4XQcmHu8wBWpwwOTdcMNmw3p3HdmypFzsDhest9Y/ofVM5svFHA7nD
ws9NmoR4IvVXuV2sPP9CkRQUZ7uzFtQNm0tmF/mZS/OTgmAkKLfJOxNZOoMKhM8U7g2eIrL/WuwZ
n7wTvPA/VlOlIQE43b3yDPM8cy234CLZ8ZgDz5cZCJF1CLn9xU1FtlJBrk4jZPls146L+AxvPbvu
yyvZ1tBv7T5rln8QzJG5hPLkBfKw4nXBf+gPOEK5leQpOzDvi1n3vW89xdXc8N+66fmZiEEL1lop
C2t9GptrCU+WSrIM7UWWfwK0N7jdo3c6mJ/jeTopi1jd72pamctDnVr1ip/NzqTG534yFeeCZPUb
hxxbK/iSexMBFSaRF/8Zyaz5CGKsTC8Ipmfcc08MvxUb9+O51ujUNqpPXbqIPxxjCgSckhEJHNep
0dffVh+pMtMcgK7XdYqbHZJNuxTvhUCpw65eZqNEBwWtOmG3VIhdNStpgLssf2c5aaocPprHzCJI
4fwCKMLZ3t0UXNeFUOs1fQQmjwfiTR8+KXXeobSbFPgLCjTK2kWRFHW+uAkBm6gMHgtSZ57R0Au2
tgzPuZgiZVfi1xC8vOBsiUUzsv2QDFkQpKbM4LFalFvTXc7uUT7emoxyjAP63G6+KMJSXFv7Au/q
EcVpOojzkBEOWHuHSXK2fTX7Bx+jb9qyFHhiv2ic+u3RoZlVUE+Kindji9tYwviembJT+o09aatR
0tdarqxfED4zgIR1UYypdOrQ8JVKp1lQBURuJtW3ypXFB6/4KbF5oDwRYfpGIzSTAamPm57BaIkK
XsVrk69ZFysQpso8w/dH9Lfa8W6ppAGVeYW1KL7Nq3UY7X3C9cgdrwz09wDMsRhXf9vrrTPCVlwj
2z976+3FYFAdkW+3P5O3PVUwOdPdBRTKZpjM8l3uLWjeEByDDVHKwz3bNE/t4xn4znPSOaBoLXZS
GsV+lFB2DX6yFwhlFF+NL/dY3nhCoM50bed2iIRmvGnxbRs+yqZf+Qr4ezp+P2j+qm+q8p2A51Ra
BwsOUxEONu2AK8Clw7cafv4Cz/4ctB1p3M7Rya0RKt63bdmrSOUZdRC+qAk2WY8XQlEzgkPiaOeC
7Nt1zxrNrNy+JQzDVAWKEm2VHNxkiooay0XhaFAL+d6+eQv0tpUjalLLMCWoy3HUI0efVPIm89n7
/q+8FBhWzIyVQBwpuTj4t3UtGeRLAmUlJ8Fna/slOJm503igGcPFB1SVjMOx5+AnWogbWvj2hRLW
8uRW+ViTvhG0BS8sgDF1mMuF6/rnImw1neze/hHsXco+dH93mSy6OVVDMWYJlJ9+vw8e/5WKu+jR
TWPT/fLewxSEid6n2DSisBQOgkG4HnfDQv0+eWVxt81rHKxAlAxmfz+u7po+o2W8xuw7QC504Txo
T9WqlTkgGfSfJ8R1G7EqOXonNlyE5igXqu4rvWe2eSb+VirHfD7R4fl/tbsABCeLVaOlOn/Dkno3
iqMLZ4ULTUhbsz1c0b3LD74eWyM3iFrkJePsBZjivDDVTvQW+VE1nee3u6yCFK1Cp+eF9A1IR6y+
Bsz4mQ+/CNmZHvZn0s7KtOqTYKEJKNPn529XLce07k1KPwFxiZHHVNvqOUejmvG2VhF9EzpZrJOU
TmZHkIag1H6RCh/p2lBR7GSYfwe3YN/HlRYLyYgUZ4uqyTxSt1F9LWF6Xwejb7lYcqXzoVYqBF6o
UflDRoPT5qv5RCSTCOww5O1pTdgjwvcM87q3f9m/GDILz8WkucmYI16gbRrx3412/m6jdWGV/8n2
qkS6DQc0x5U+n2u97ki1uckmSePNLSOMUcFY4ZUod/3ICGnaR29ODMOMy8U/CDYoplUEsFgslwbC
Uix2Pxzbo8ds/7+8SrCmrb6Pcku2YN9EzjqeWZQ8yjheWl0+YVXBI8lqXT2Xx15lvaY7nHGymcCA
r+LYCRkXg0J3xd1j6lhirYnnUVNT2UoeXbk6wtiL2I/GxPdkN6ksd1rdezbnWSQBaa0J+BNsZekH
rJQ2VWoXLSAU9CWprFTVApD5l2g8tYJxLWJYQIMM125Dr0MJRrTJUvKjLGF99bDaM01IXhkgAoaT
U9NrXIOri8Pzvr8BKFNUmGw82VICua5JsvrVGHeubrQ9py0XCXo9K3S61HqDubfs04bO4gvcQv+r
3Im8ZcgYRod01cEyXjk9F89RXdzknwi0YDZN/9h3fzHgjtW6jcg1zvT1tZEdXQGdElK42x+/FjNb
A+zZ//fesh3e8OZaPHCMtFxAXqdwjbZB9go5kmgnrLV3K9pToVqRjGk5g+hiPqTel6uhKZR5S3k9
9p+i9V+1IR0S3OAZV26nLIAImecqpssrCrb1XBfwIBSiyb8Fj3txafYQO1imuWyC11U8AFxwkrBB
k8DhT7EjV7YCzM4wJ3ywFAl39AFTBmrDoVIq7fPYJn+jkJedw7D+H+sawMCPJcw3oI1XMPX0x73Y
uNKrTM9Xzqpp6kTEGgeYV/WS6FSs+Ks9OuPNUMWJ41vOXsW1KsIZzq4TuiqKRmNQ1PfgWC4Lutcz
zfxCZdUdQh82R2C1Z+JS9QaM71DrseiWRfutujAL4nZ+8x4gcfGvMgxFNWh74q27cwcEwV4pY24n
TrZaC8BOfepXWcAArPqQb452Ckrk8cP2fcIkOoBpc+Cd5hJQpcLQM08oVonxsx6g2dRvNj8MfpB4
ZBOdPLgltDiiD6ei2wGd4nij45/4oxweGivMqqQV9gM3Kui6OPqmY7lqDXcN3u+EevaDC7W5qXD/
0PSyTYEL+UrvNKW1P9SslpcZrxdGbyF6GPBPtIV219b1fUcj8kG+hrDtZOSuqvqXNsWg8T5q6Qpt
P13qaTvqAEfbwKg2H0bfUBb5dtqEs+mGCvtOTyOZCwUjq6oTNPu+E+7xb//z3SIYF98EcGVKwZ+F
qjmmLyoSuehrKj5Kar0VpJI8zZX+0RP2P8c8AjWEmHjSEF5okcmOEumXbXFcWrDF1wMquD9kLsUx
oKOxBMtQKU1DESOlj4KYRjDjXFg75wlhqJQK5PUKWQcDYA28MFJ0/6/uF1z4/yC5W3zAqHAqTDYI
CQR9LDxh8RC4EFceg9HfPEIsv1JsbAUu9N0vd8+c/M/XrrvLLFM+ioqbiP3FfVrjlvC0kRxVh9tD
TBbDVdhWWamp5Ui892tg050Chjli49iuM+5L9t7Nnib9ykotkY/d4u4ywtmvVWmPXMc+xVi/BTuB
CPRSyNdOV6hhL8KL2HGRREBMN5KsC5GiARCMjkvmyN/CXDT+kB2CwI8mT8uH7X9NlMZoByfPPQbY
Pbk9OY1jpvpSINjR54gZwDZQuvJxlB468Bbqi0oj78XyeaPg5a2dtgcVvUdT8FPT0UOt5u1sx3zh
r90f2n/rS+gf/zJ1yt//Ldkw9HtGV31rSauo8Z6VDhRticfSG3BevI1MTdm5yJf5LAYatQ0R+yGc
mshgwidBMZC1ogcr+QO4jccALaqHRqeA/BVR3r6RcnUbahU6mbA2AgVwFjxXtamoIq2stofIb6iC
iYr7jbufNeqcEDOhcqZNsP5WM+RAma/9vY8JCaVcI0Jw2J/eJjtLBf+IV2HnitvIWmYEqxN6z6k+
8NYICIgiRldOq2Rphx8dE35rynN2UxcNTXXWj5slexqjJfBdbwcE0EYF8BlTuDG7x3KXiM/oYqys
SlP0u0m7BPSWgZBXU2PQWIn0w6dZURPeqOxG+Kc9EQCsJ876PJ2Xjj2KicuGs8GebahhcD/1rtBV
ELGEQg3ldICFxdsayTKJmpqWfNwthxDuzi3eHrWTauafH1sLgZhw8TaO5Y7+6iHrxgmAt/II/iZB
uFHob9qbJQYXMi+qG6FvDgFJnKtvWQTUYQVImpSQI6nA/4um7DBHinmXM+VCByLi2aAqdL4zIaxc
RPVvvp9Xsfhsm3raoc+GJ+GjUmQ7UYQLRLrAPHhEPcNaDjvjYyhfHFMnCYVIPk5ud6PN1kbMbJFr
vH1g601FjJ+A0JW50RqAZbm/Uir2FFvnsePf7qZnQwhNUwVOEROjG0Tn+ubd+rAn2rDIWNzfT1YX
KUSIclESWAlSO1BmvAOCQ4+2ik3PI+pPWiwKE2eN91ot9b4/iLZ78ceD+RdAYvMpMXMzmJnIiDUC
hxze88ROrW7jnXTHKA5tIQ2ezV/F8u4s3Uwe+pAm52ismZvst0QmZUKkzDnbZt0FFsdKvprGEA+m
jbBPDUX/NNP+tvAQvZDkr5HrcGseHr9XodxKlcgXkBlMs2QqIJpZF9uf0iQ7T9b9KLCMfRtDwwdt
Mf6VL21VdgLQh0XB+E/e6Bmeij/yQTh1D6n5LD6cOYp+xuVn/3yvCw3sevo0kQZ1QA0cbfJh/lQE
FUSIWQ/1rdy0bzoriSKqGv+mKWdjnHvGDrGeHzm9KcrT0lM1Q0jPC0csFWZttN2N3QhJt2CZO1+M
3EVRe80kjCSJ1+Feh0QHmcKOFPtgGyz3M03JxNaHrGYeyWpG3z112AUGXjd2+3Dc2cSffg4WQHMb
Q3pakIA96aGE43zERPypUgw5O8u5ixC0ngv63B5x8NO9khuBSTFOTW93c58u12kKxo8IXtsRYycL
nRJvmU+g2O9QxqV5jGVeAy7i/SFjRPwKebPRcVYNorC0714S54zOPJo51fZK5lNtmUCw8F4TSf0W
Qqg/tc28DlyPCtdXGpEvMm8/DzWdadIbIb1PyM17272eRTg8xYJ4dH2x7q8PLXOQTmcXFQthWhw8
4kVvzEd6d2z857XtIrCbOtX2hS8uLMrUgZcwwuPEvCSWZAx4/UZ9kar5WKUmBld1ul0KIp+WsgWK
uwsLhuRQ0jT1dxC1m70FZyYt7tMjdVDuJr9+rWnGiCuv6Vma0OXJz6tgMNg1SNUdw1RfqKhWZgZ0
+bLdT6h5i4Zikz6muwsnjE6WGSV5Qreq0G73vqf1yAgqRR+gSH7olqjQkq0Iwq5w5JpEO8V9Z+Iy
yQcWOLLsbIdVCYzMD0H0RAc3Bz9SXMM+yHPWi3o+Dy4tRxOg0vXOHyo5OXb/Y+3OKtt2Nqy44Yez
r6mSn911vOEDm2QvN/3T7yShYfzOPDGY9Tn3mC8SPfzJofvubHwPmBlEWpvrnjpExjZM0OoM9rVa
UUEpvBkKIVV25TZF8p//3PAOWWSO6e0rGavQXdOYy/RCO9CL87oESMJSKaYbTHqhj+3zJe5MQjab
68OffSSvHzy07Os1lwsYeT4IZLkEtXOYdcXisQNIAJuBWHM5Hlx6Zm7goX9Z3k5OFma+WUoOhjf/
EXoWYP0RU5Qnc86UEVaGZA5ozrGxbbeL7Cl6UX8Pr3iS7WHiBc/ljMCXqpdV+NH62jhSKSIp2q9P
ilB2Qm/nmi0+qG6KSLXiVyfAmJ+wFtbITeM9FBEovjsz7fLbWcT5364rnShtCwxpkzxsk6Bh9YK3
IiB4mnzrpv5Zrnlx4MaWAZ5hun16b3/zrDG9EPZx/NhG/9W+CMXFVmdT/gvhf+hM3BpHVJAhLVUV
qG29z/s0Udxunq1LjB7ubpQf9o0hMR3zeC+0EvzMahSq1gFCIJOqj3WweSENvxPrt6TT33EgwlKs
jB4DadIkPhLrVXwF5ORbw9rYA2IJ1k7sUwDIEEfs7XhaUmCSz4fkxJ73v6KOWt+CrT+5rxsndNur
H1aGIw/X0qSIaemfyNij6T/+vXgE5GfXy3XN/K9kMKzusqhvwHvtwAx1fBmdo8l8OP2I44erzcIh
K4jHIjxfKkzfXtXe4OJP8WOqHApH5n20iabib9DMEk3+DjRqsitzkUM/w24q0mSc41omweuPzw1k
Wiv5heUMv4AQ2QGasT+E9KcfJfZ1XEwd4M8VhZUIBS4YpmqZPxVMr1kmeFM6G2xBfHxTItuCKyXC
gIJk3y8OLBMUunXSaE5uRbbjye7+Zi8oysTCeiNfz41JyALKZ/a93mamzvKecO2mB/hqCalg2T0u
acArzA6yB2LRKlHOpZurSfGQsu18MrE6v6b49QnzINktqSr4vC1hbgDCyQNu9YXa9qNOuvnMDB7h
Qybt/h2NvUGCauxWq8Peimag7P2buaOcZZj6uac/273eTXHVI6SDQVgslqP4rEtIzQ+8G7NQqKYg
FAJrf5ZMN5nixzmla3wTTw9CB7g4KQYMO5dxaK74Gx97/bqMNCr9WIj32vl26nsRDLEmsyMAJ0C7
VNTQzsASXiM5hQByyiwBHts6XYHXmmyoI2tZ/GebTL4BBfJsM9oPjrNA/HnqKjXUC4JWKIvI+8Bt
iaImRD93R6rIUFmN7q0D0JUIHV0A5yPQHQfLV99r9D5t3O+dkKQK+39EqzeKwdS8NyaGrd+fjMCs
u4+Lce57C0aYk5/UECBQWsBgyQFo+pSe3e69HotC1JVAJPHGk2i+CjhORdcWU8h8JCZccjuVHgP3
kZ8AtwMcKX22oTi8V9enaqHb5PEmQngrWDQQG/TlZdwnn7P4mmQi1Ox+otEeNYajbjY4TQWZSTPe
ikL5Vhvn6ZQp1rEc1yECN76ghYMslGb2g4ZEFhivicbDCZipgdyZupkGTnqof+8YOWonOlVBWDJM
rfgiWTzrZK9YQybnH0aMie4sryQzbxWNeOkTPBCWuphZ90JeYBnbdJ/NJwcQPC2IztSkQT6VOgrz
NUFZ2M6ZQ5hRlWDcT4Q1yLteouXXbmifCo+IEeGFK8RbkwQ9EoPRSOUqSdphSEqROP8LMCGvknbg
p5DDj+6fRtw6+NiT59oWqlTuiT5laPM8p0ng0ke86qWq8W8ngvpPQwW3E8j6SywpsIFe2mHztfr1
1CSzRYC8/4UcUn23tVfElV+lo/NcpVR76JesqeS/6kfsS7QZcPqT2CNIh6eMpVCfQDsJ9HcwX8mG
PsjgBq53vybiW8umW2zOufSliIpQyqmDIfqJJs/IkKVpPrv5xxGDJizT3UEEo6cUj5kNs1G+bB7Z
d4qUIVT4oM55aIN5RXhWAqtG2VYmHSNInSaeD1FlNCdBqGt7hBh0vABZRgi6wQoEwmWkOY2ayZo2
cOgDSwap7X3MXlLtpsDbOgN0wZrkUADHzlkNFnHIj+GjUlSt0tlN3G6L3jOdwiW1so9Q5wP/zEn/
aaKYB6vzt1j1sVO0tEPCz9MBZdEMjLpemYt/LMhtxb9XiQ6/5iCbSl+ztprLiDIA8ifo2aQ+qxFK
BsYSJj/nyeTvQxRbt95HlJz1KWKwxaPVDzzwOtI2+8h/Twe75sIFNkmlc5oMh/ncvDnlX6l1hAHQ
EWXFnixyCw6BwIFzXt+8zBXaT6dHgOlZn9Ac4MeJk9zWoaGIJ/RrHFYDNNqrmncrWnXnPMyLMN+n
IAzS9PEwRD0ZbrejIY/4RynN7Bsuoa2fiO0+WuSZA/EOL7WKsSjQ8RbbqxUUxlnykJ3nyiAkU91+
h34LxTbeFedu+FTOwiNplbGDgHQgAlK+DpkZQZBJQmH+c5krINHm3WKSkJGeBAiLDpkycHh1ADvX
/l4+zQ1Y5IVKJ0CK5tXVxpY7BLKxJda8mC4fBCKFYbt25Q3a6vXBYW9ybTNbBbtJ5E+f2Ru+b5k+
0HxwPpRMS0Y7Eo1r0uxq0S/Aao7NwX2Eh32ggHBvkQjFVP4SrS8v7/NTxO5e0VWfNGfqSIbqBQ0r
sVK7EW5PJChkvmscEFoLOrAoEgx2G14JszmDf4VfimkXOTEZwVOELErCVPZJ85uMQemxZpAG9Qqo
gXIoQvkrgyT4fWmvFsjf+c42Q2AhwDsEuK2PqcGvcVkNmm0Ab7zD/0wj6ucuLAG3bXkCITX/3b67
1twHYznfhVOIMlixQsWW8BfIs7SEy4zdMkP4aUgz7N2rhfaT7+jl3+r2WI9Mu6cCom8aUrAK0e6p
HGZ6CK4UMuISE2t3vhv0snO6nGpVkRmECHeXY7G7+YNB++6XihNZ8txtbwYkLbi6w3LQzUEc2cls
K64KfSeCGYJG618o5Yyjn2bZn+14OilbLZsEw4bZ+LcePxYIh6FenMcrOvUT4PGkDC9VtCbjdIjM
YyUT2haF0kDOLnaJyGQIySqPLwX4Wp0VoaoHEK1lqzx2LGIe9uP7BY0Jij31i5AjQBOVLLc4Jxr9
OzpwwLCPpnXOFUEpLT5BH7vvAnc5rR9V/xn3nJVDwl6908zSA2joMSs2NSDDMUyMMOaO+qOsYyys
Ec/2s8zuEk5gd+ilvJlwZy9O1Ny02yNK0uD1+Iheb7mmd1CsS7+YrptA5N8gIJ9WquOfzUDGtuou
RCwkB2Opgvm0BJJ0dMo8nMsnDyuqXub+nk+Fr+f+7EBscw9KTLELy+OdU6pG8KTSMLeMaA5xOPmH
PS415A9fnAg+i+Szem5r9fdAz+0G40M9Ur8eXHndKGwqb0tPwyiqcNeaLCPF3rKDee9YZoRBMB7R
HfYZZ9uVjiWEjstfRhi4n9HW/YdyHKDi3EwOzAR7oc7Xz7brexBCwLgco4aD1ssjhC4I/vsJbt76
mHKlBSZp02+zk6UCfUcNLq+lzvIOuSFOEQm2Bja8ZzscHkqOuIJNRocU+DBWbnFJnicUxkTu5pM0
rUF5P5/fGhXyrsqUbeIVSgm0guQnhIxvSQZLIfP8BBw13//OTkJ6U2pB5ipHIZpbs4US4ZK8UjC+
2UCNsLWWW7IYZ7UPezvZGJA+ReCQexWP+JQwOQDYHnJN4FanfhrZz535zsYos0omu5Afz54AQtyx
CeldcrPLrx+DAaXERqUWu3SfinQj/t5A4NTTnzwP9PNxxyN/d2ztVikRgREvpn8zaKj85+POP2YB
4689pJPXdT8PP6wZXp2RA53zykXFBPi07NbSaghMO/vEZt9E0YyO3TZuOwlbmg6/aazXc+xd7c1z
b8HXTCH4X7+NWwAOYlEobNxdTftmHZZh2eyMqFSNO8fZuSGxUjXY+DU1d1iSCHPmYBHgf7e5USB5
spwcwaB7MrOvoiSJfmuhvRscCEBLu210ebGJkkdT91QyFI0tbZeOQW9YPe5il3XPG07712cqpnnt
dl+oOEV7Ppfkva3In2WRnPwW23vtUFejgnhXLpsVWQ9JakyPYcfwNvX3tLOCwTs1t5tf03Rblwzy
lOvq7TMiNEJafPMOLy8m9eoVq70BzxEwRtVFDipY5d2S4IY+73Pg4VxdjkCpMRI5zX+8vjhqD7jx
TaicTLAXRyQ+ny/K/H2RNGFS/zaRj+CuGPCYSRg83z9pUheuLCovsHEgQodEQiEpbfGfYQqPhdKD
GokZo+jI9nwObCR5weqTXCynVkHmulP2NeTOx+q5nb8nMmLay4J6JhtsS5gKz//XsHG0KJxMgnEi
eAFMNEL1tnZ5TEb6W2XoTsOjJVlwyHDvbkXD7PMK79G9kEnMQk5lqnljiED9WZpHJvBBCWnP3YgU
9kCRauKy6xsMdfbZBgrVNvTITH0V9ceXdvuBLiRXiC//bTllU4ixsN4arEhwumjaTthWuLll6alM
JpQZFWE7hruzZMxq4ZjViJfFj4iAgngrBjEB2gUBzIoEzFe6n9I44C7D0uPl/GTGGw2el5cWPU0K
qgCeTpzY0Cgd/7/uH3o3WO8bj4tT/K+Ibar+6CkETIEk58K/fiIsGRbLYgNXlrpxVlvggRdpObBO
NeujHui49FPR8w7nhUw2jdTVBCrCPNAbpvDA7oBLj3Ry3GMP18Yn5SsdJIMHucwtc37KCPHN+4zB
QUYxCXP3fafts34eiVjM/X6iBIWIWjiRSMrncb2U0lxG2vbZMLAqWBEIV7RcgVktsCWtX9JuttNy
ZszCyEl8EQyXCwqfN2JeUZ8z6YsxPWkJ2VhtHU95z0O52xio/15va9OnPEj88fiCvxWgcxzekf9L
4SJbuEshZduXjjhutKyazID15m6oZxSLA8PZb2Ua0bqUKbHIkxHZy45Hwm6izg60XmptpvZstiPo
0filXyxghqq54dpVTa4SVLVA/umYg2lSkT3z0JNY/d/i5PRwxbJ7cTHcH/YHg99wyBT4TspHBPZA
08qmwgmj6fbq4J6cjMB3MkoDudNxs+v5Tb7JlTWCGrIxEElRqUV8RpZbbjkuQF+KIFvpwIpf9Oac
ArRi+BgOzi4ZNFp27J0qg5BvhEE89gRTSKfoCY2zvLshIRJrRXL+XCP8xyt0zwA466XkJUpY/m65
zHzQ04H6SN5+ne/s67qzgkpeXJrgVxLVT9L6nB7ot0J0wmq0Y6DOBSy0irp487OzYr54zKE0ObXR
AlV1x4s1JuRIcdw2izpGifO6y0h7C12QDRIuhdBjhdakDkhYBvgL8aozMecAEmIUfhNE43zCFXrP
7f0ppvV4J4w4AFQtEg9nr+3Rz1fTF7Odk1uFN6Yu741Fj6vzRHkU0cx8TP7PoHxYrkHiZ+30KnNE
A7gOpXbu9lhhg5wWBm36rqNhiYHxEIn8T6EQzuMinB4Tn7fETwkCIgGtWYrzT7TCKzvCRxX6JgD8
pb4gXTbjTuxptaKm9hQvtout9Z2Gx7025a8eblSkoJ3QxTcgvCHu5wBPEjTLOU+9EGWsAtHBBImq
nkp4BPDWc8Ohvy2O1vCznj2+7zjwVR1pH245OW6WgT0P8ss6z8cuUTuVMHvgoTPXwDd1vHJv8Ojp
hY3tb9/ay2jnuVh7sL5lBg4Uc1ACKSdk7KKPKh701592WH/lOK3BtHdjYur0VhdEuS1EzLh2u8/R
OqDdKmhgVv0u2g2DaKN0ucvFpddBfRQ41tdHgUTlxp7IHrGKdq+1qN5RDEmBGfL/P87eCbGIX+Tx
7itmKB66XbOAQzH/3Y14yuoiJavUQq56FGd1zjP34aFSAw7fBN8TN2GtYXJAiZTD8K8zci9GNaH3
qIje8h3gHOGODm+6yMw/yZNVKGnv/+5t2ngih/mjzLPXBBuQzTj+JPu7jO1J3ZBngyKNTazFzz5J
7M7hZEH4LuQEVWwCcoqhdHGVwQNZwXNEFSNXVZNV6dEw9aYvGHxrLcfm2HV+0IO+LC16cI8A5RJn
ZH5CK1BI88S0vJ0BrGgO/vfviVP6nH900og8VUZc9Xdbw1ykpYEgm2bgRCTfAXjWCX1L+5k75ivf
U0HTfsNBWIp52nodKYoAcwAT6KRMikaKvNQjNVNJunH13XZD7AiCWEHlIi/MKjL0uUevPjLjT9o0
fGdFCAQTWXRnLILTuUh07MjNMUekZLIqv7woM/ib/77zu3jlrbnKjHysU9dkzQN9ZRNZucF9j0i2
zN0JjrEdHIutsliHzDrf+0Rb/GmqMMHaTkqO/PdF2dAPuP7McHnqVFNW3STgapV9JenFFkiw3/us
LNGLx3flVJXZ2yHGUaDp5oZvzK5i8FgEcT+4KnvF20oZ3qAN/gjq3o2KosAuTplu9N/HGw6+7082
R8rTDdMrMVUk2te7rqgLMN3Whp7P1N9c09+TLJcsb5x+Tx6s0p9buYz7yT4U/K3gAIH++37xNUPE
ziQ6uGWJaawWw/gtimjSpHnOhvw1CLc6njYcBnHRKB9Icy3vvX1xy3cbX0tfb66eDYJKVkH+i07p
dIG55clGzPGTDI/TJZAIKJTYI6UH+HeaqOs8kHVU9awBJJMm97dabzx8J8GJTkQ6CyM7Q5vaXLQJ
AlQ7QWILFi1Jwb149cQh4kN7Kn59wWTiFpHVvv7RxXgGxrvrJUTGfk4+8Pb2olbgeRIn+uxaCZ26
NKVWI5orugN4CgTdj+GnG6M4XL97OFS2p8nhFpa96wBDNCYL3ivsbk+TX+ClSwhbVqMJkaJjp4dc
ez4s9DDPhMfDpMM7XKVmIlv9WUZGVPPsxfjMiveIFuKs6iwq05WQumxWuabUkZ8y9y+qlGQH9r1F
3k96lPFUYhL5s/I3praz/3g6VN4/NsSuWTbY3WEiQi4eZuCvHV2PCAWuNBG/6Nqn0KIgwA9SIgga
eeAMh7XZSQIxv/4ngiUCEJI4SyQLdOPgo2v+21aTi+bEa9tTsqEIjdmudMMu9671LQyd4CGi+rMR
ZbwzHE/CpuaxA8oswSG/iDcmEgkIESIBibTqHGlBMkn9UulMIZqn6JWKkgT8AvZX63UlnVOOpyt4
SInlP2UfP0BTHrV/Kt4P3255GQ1CYfN8o0vvMN5EhYwj148qWTY4pkdOol14S9ihkVrx/G3Hhu9R
UEgKMAKwos8gTsU7rCLU83TRtFbe4dRVutDz2vs80ll7FcCOScHRnXiW/SJfltiv8gytyTmTrmzI
UqO3Nr1pjOPWEakkR+LsWAvxLtup2f34nAz6mXaIaHl66v6EP7jUYcaeoePnRlJZHdjfbUh8WcOB
9CkwgVMYzT3HBJwAg/AVLhM4cQcAxd9xgbgioUHMJ/+D2KRecn3B+kZnAOT2C4A5i8q7iZyWj6A/
jbjJ0xp1MmZhSwj9gyV1wnfrKiqhwqde+BWDkBxxGO9QZpulZA6ruXrfuPTRZECbnARWJEYHYJdv
rQQeBxXgzYPshRIi89ascFrpL49CL4MT1YanQzu60948a2UrUrHTk3O0AFjju6tgkMRsIb4xFkJl
lhooXZwRj8YfO7WDvEsyl3m9noDKKvbVM9wA8NgMKAALWo3B1YpJ7vbDc7w7Nq291K+aKaEKNWP1
nCIjxSiuCktlVhlNfJ1+RJe7Gg3lSyhK3RM8oCQ4WAjTRb2yCJzJotctclrm90dJFd7/4JLzkkj0
byz14KwyWSOuD9cN8wOlNqfoeDLnUVJ44uIzk0DyU909QzUxwSYArRwgdhGWgfb5YLPneHbutfZT
wy/obDr5TdxN5fy+4taiGMJNPGkZ7PvgByWys+USIsIi+OU1sktUHqBw9Vk3QEpfXUGH9QjuWqjL
/UgL+faw1pyk9nWHeS86unDO4tqXB26FfKw8T8/mmCJkaL0iKc5W+oU/HI6X4g9fO0eMChoIQFcf
yGRwuqoDgwyWVQ9WQrelcgO3xo7YstdQ4VMbPrfhFo6YzNQP6c7ZoCZWfBEFHEmwUhhnE0jnyzTc
75jVI49g7f7wBoo6enx5olY66rNOrMAN9r7FTZRWrsbzRFRxINA2wExNAh0cGjeRZm7vLXdtY4EC
Gx9rU96zIAx7Uq2dS29iq0AxHprADesz/2/uM5jgZX9XDViVoxC125LCGT7SDFGGcSEWnAcK6OXQ
8EIhc1lgPXGx9fPrnJFf1pc6W6kvFU+I/E8EsOgestlzi1wpTD/v7fgdchek/YAhkddFRNQuBk50
uNO57Kss0abHxYjOLmTyJ2qMbEtgLeV+CEDYYnMu3pndU48d8v5dUl+XVVpC+mpTMqUmLEbv44pk
Qer2rRPxnUSQjp/96VW6+Q4A8aX0UVWTDOhKg3kkTc0X8vCtIqjHmSX0JYmboP4O5MLAixHglAyE
FcLP4usE2mggMyx6vzsmWMxYw/+88Ojba1B2qeX/uCcGxs9qhd+0AXHJF79olAI2FszyD6XFmdR/
NF8YztEZdzSR1bvUxpsF3GLl1IIsfUMulcIAB/fkL1V50ulcoXmR7kzYcQHpLixaXJgKp0caaDj2
jHqswR+AgdjmAhNfC7buxaPCB29/BQDfP7mrrIrret5UiVq7G7Pz2IfuP64x+n/Qmilf1vbevv/A
az4CbY9Zndx5VZ6kD1hc+5cdnvBW2W2uC1C6Ao5CU1bCkEG2GTnkTXSf9hY3GgRArsqmDf3l/lo9
6GxvqaRAd7Ks4JaM8TFSBoJ40wmmundSOp54Ip6jBxheHdmG+yVfRuspBbDR/8tR8LIe5QTzd9fM
aJOrY5juhBtpVo1Cg8X+hNHE52YLsWc7vYxy5BZw/wcMLpHtkhTHd0Q7WmtMjBGyOZE/vlibA8eH
Hoecl8cnzFZfmwPHdHYcYyzyb7d3g27EMQQxPkzs+T2NEwi5mqSDxCMh/HQ9269xPoiHmL3J1OR8
+W6W0R+pVr4GWtltFHuFof1N7JOUOHxRJkZBkWD2/hcWAKjf9t0BwghRR5F7Q+4490lr42mt2wt/
h/bz59KPvGndzWP8cfA+HjyXgU2KwlZZJKgn0Yk2ciuBpiBp/Llr9T6Iy969yxbk+f0+kgZU+gib
Iv31cg9mJ+hU7fxZWlZAuD6hXEyA3hylYDEeuR8xeQRMIRZqFtaXay9DYF9Fwtv9XJRXTsoOrqS5
Q0yRVHQdvQdwCZeTVHsJ9FgS2DAe7t53caLSQuvylI2PZ70wJJcSJpi/ukz3j3oimbxTUi94im1A
C51dSGUBYL9PKBki9Ps2UKeFRt/d/5o6T3nRXTVYQzQ8kiL8P+36Yovz3hLvdyD7Hy/WKCBiPerZ
Bl95tO4pxdLA/Lx6QCtqBw8ZziLP/1sTyDxhAkKz1deSb0ghnaz6yX3OOhU5p9sGH8G5ggee46YN
kqLm1ucKNAQODTHG+w2qYCq1YduclZoSZ38WBrG5eMrydLW2V8SR5QBE7d3jfwuMcYiEbZ4qkIm6
lrrQuSXe0z2BiITtInsH28m+fQpS/Aq/ji4n+XkU3DykuiYE+bI61I6jgchBg7cTW8GhylychRE+
xtu4S+S6628zTv1+SB+lWbcu1AGPJm8aJqGD1VrRD1S8ECFa5iTYP8N2hPmWsjwUz257ZitbP2ZB
HlTskiIYOf05+hn+VSP68gvTI3rld5RRsP+5BC0EFjfPVDvnjc/xl2BJ2V0c5P/IsdnKiN9lSqjW
fNCxCpAbupFzMytZT7TIVQv3lntDjZ0IU8yYuyaa5agvxZG1Pn6y5FncvjjfjTwlvI5Em6+/mfni
OAe3f1z9dlPvSZxJw7OM1MSWCxL8q4c0A7nOybEjlKCackg77Y4/M6oKhnwieLNed39FWRYEragd
zWn+mc7ptbq3xOrIfqaYK5sHwUCkX7zWUA8QojXnOgDATROA4rtSqhYX5ALzFvo5m0rKvYf9iFIo
+HcU15Hr1+CM0inJYSq0lt481X3TLwORWRKNyDK8g+ZxKiWfOJgRJ819K3RnIy8LVjbTmJDbVZ6n
Kd5LoTVKUluebbiJnajWb1DGMWEGPMDQmQvyHEt+XHlWpKlHD4PvKSVnNdlTqmqE9MSjvAomMo8R
j8GwsEBqhcE78vRNI30fKY6f6jGGn5UgP4hPe8Q71ffG9wnzM28VhEvDVbY79eE2bSRfc/PAnHHV
65oYtQBdfsseeFTL2I2o/D+SSDwqCwRgZB3tmqBkz15CstpVllhWK0n5+nZPZOT3D5TfEVjGEDbQ
q+oPlVLXAgQjbaVG2olXq212svVICQFaHUcQ/LI/iIPuxrHdF3Pice8qQ6sE8ImHNJHOYjD5m73l
vOgkZ0KECtkXbqChpJO8+HbgyTrEOt8A3juMOLfPWS1XLGGp+LcU7rScKk5chpx83SJzPyKSm43P
u5RSzYgCsARuenAB+NkiFtzQ+0vCcEMMz0Ej1UTAwN5CzHUzqEMBWwAAMsFJpjz24JU67aoRolwe
kkJUIeJ7EwPONpJ4C9FWAojtZ/BX+jYH5JPuu6r8UJ8F2jszl6eK5xb7fmb7CUa57tDB202r9z2U
yPdQcxZmGmSvOVePZv+7MEIe+K2u0jcKZrkLPaIoWQHN51rSVWdD0n6PCXbCSGO7EAMFDUJ8i2kP
BvpVInHhsx12FsqTuU3fbMUjAL8ZLma1l5PLXhYOF4GI/a+gvwvlBJdW3ey8F3zb42r0SoNqWIhR
w8qhb4sSX9ncwyNg8r+aWGaMEm44bmKOj3+W5iBDLfNn1xw/uyU2SsPKxRpwvgXPWdze+eCbKgF0
HKOvCSw7Ae6O83p3/QZngfXLWgV34wwmTPohfL11AQASWihzuxJpWiUQ/CrkyYPXcm3VFrp9F3jC
pmCnZgS1CtMrhihp4iJieTUdtvi5Ou4qzhVZHew7Bp292Hkaef+dTZ1n4QDPF1KojzQT6OKnmHRZ
7HRL5H4qEO+RkYm279v0HqQ2GH18GYQLtFQdm0QYfXOdhXAX33vMhs/M32eb9DjVlNx/vRetiFZl
e8gB24H0p9m7Do2qiGjUWJHfFgkqb9kJQCuCwQLkBuQvoIjlhE9qZtxNtXmJZo3DZS/WY3Zw+k8D
vRWSnor21fkTrBY4UBuPPZ/LXVINKMQ+spKUNz2hjAj2ojc+cczHY/HLABmz7SeN2Z1q175Hhqx8
BJ9vXcGSddGeuVFrTrwyp9y7Vp0jTptTuocy9RH+Yr7PYoLosM4yIEjr79LUJYVgBQD1X/adLENK
fF5os70hr9nr6FAlksPtfW/tvUdF5e+6urPiNduRItlh+ai602x/bGiqpVyo57hclKQiKjKVBFLI
m8jIn8p3jkKpse1ppQPD8uX1zQ3CCwOVNX3S2XroxXgHjZc4AHt0cpLduRbPxIWP2cEtHV9XfVht
nOK1hpjQ26tqXQKXOv3Jz3uZt7RHDv2VR3RqraodOK2o3PxPYpCFox7Z8g16OfBb3upBeFxWDUPH
OYflA3kZ0/e7+5bgHlFzaYu1yuDLACYt8tg5l9VgbNXOMzX9N9TDnbD08NJSNj953FdfXv3XHJy4
LS02O8OdRoUOdiG9UU0fh7KhVzShbXC9Mvigh7lcfEeL2jsJBwOllsJkkGOBdK/Lw5GnQXbs9xT4
Fcw2cDgU/w8wsbLdtI4S17urGfT8sExZzjVRpDliQBrfBINCRLzl+vNmMah1EXAShKEk/nYDZfjo
H6s1A9A7Rodl8snYocDdtywlyW2dR9tFCwwaYMBA/RB4tdP7aIg6LeOxPCq6NuoVyjO3blgNCVE7
MvnJ6OtWTKIdpNePqWt6tyEqMm6Jy/1OR3hdS3HRK6YJpRbH0KKytWKz//UgeT9AOhlTdNSm6cQM
OZK/ERc1l/hyzjuq6uBk0uiNvfAODA1maRXsf8O8nhSQBYRMOoAfHHukY8qPe4xoPpnyjuKdxrdF
2dw1y12oJXhb+rZHDSguzIIM9R3A7WEFgXichAXR8AbL9MrZyzZwAbKeHEtaoxdb/yTY5ODlzsIs
YPSLULaoY7lVqCb5IZKWgC2SjoNV0MDJafiXrQL1+GDW2dZ9zueIttKdwfAfFMhnDWWG9Tb3MfGs
9i0P2EGxfiHqENypL53C2rP30CZlVTNYGCKOW1k2kN9al13NiUXNus9CqHjsLaRJNV2cV7QyaGsG
IDuzBHWKYeqGnuAtOgh3FxQrdxXhXm1lbyoUfTVm/tO9uoj8yo+5JF/0eN9csu4lu4Eo2hgh/R/b
B/tTfZJfNMkHRcy1K2z5KQAjKNAV0rG+Wh3eM+S9mR9cmJtF918cihxmVxFN+j1D3Y4RRpCNojOA
imERS0y618YraTy6xRCDq0g/mgzWXW3aeARcNOcQN6SPyRmhA3LMgSeXwHEDunXleSGS42U+mBm7
sAMUOfiC9e8asi090z3oBPDAEbEl8JI47a+I3zjdrdhiK6+ltEx/dRvH5HU6bFWR64vwQfNXEyLK
0+o91m9cf14mjKe1zbyMNmsJ3dxkG6ZW4gI6oEYJKPVLA0depeXiqnwP5hphLjc2Ga30DTjjbnAY
MB2iimFqk/gfOae/yYGY0iN2Q6JAmoYwPw0exYwhHnRBpjXihM9UgH2IxjOPb4Rc3mVP3/pUEtpl
RFl8GPbW38y/k5A4b2gIjGAHlpcFySWcWOu6Ib3ZsLyZLTIwCSjX8mZd23oE3uUb/zTU5FXGG8fX
/BI4aIKSQDyLqWQ9us1WC8o5hrt6yjgbHyF18w6pHiZm3w/ZgGNycqFK6v3KHDsdZtMXqfJl3V+y
aE1g7LdcqCJLj7rD/S+Vf8hvPKjCXQe2WHKFdpeq02+2WTAj7UAlkYhMq4cQL3e3GMoUCTungH72
Tp8CLlInUUgqiWSohY+4HNL2N1Q461JWljiuQrEFTeqlLA376r2GAglN8C+4rQGUduG7EdpYx6x0
WQ4UhroyWfIA63bWOFq/zuJE03KVXuNajMFOGe6Gcc9jZ1rUZWc9GeSaZylz1DfoIZv37xfbNisI
HINLkaj2prM7rgP5rJdbU6fGScrmA4NnfeA/yRykn8hxjOiCxHqo/vj+FpjX+/smIFG6ckBRZ3Ep
CYl5FeMbTNMTig2Gmga4iLwgQ6Mk7Pajk9xxzNyYgaGtUYMpgXyjdCzHXRSf2FBQetqpqDAnzfHJ
OOfjeq4QwEzunmAG4KkXYvBv0cAIiKnJwIJpsa3HewWPzvNDdBpbNEhkvAWkeJnddtOzPExmMYkr
u75nn/g6FCCIdsZGQ4KW7tGYJ+knDTmfqxSdl8pSGpkTq29kSisjxOOS5kGu8hsKOYauIO9o9F2v
BR+KYMqv1WsDYkmGD8IO1yKUIXjT6mbOJHuIOfo/VANkOdBtVzHtDGkbVKHvPOvnU0d9X7t4gYiX
wgg/vntN9Ac/0MBKHlTIXkcyxs8u8Ge5jk4ePWpF7cSDSjW0GTVAbLwbfkuL62Tm6qiXnZ5m4prw
/zjmahke9S4BDuydGq/2voSbfsX3UxO28aSEQEwG2tkc/786lJ8wmCVYkCUCi7meAqiyutZw1OzJ
TZj7SdepoZsgmbz260rJF0IiVOVQijxuNPuds82pUwED5E9/oMMo5MffjqAZ/75s2Hnoi6HMgCcW
ZQZBwOT5Cjoyz/iOWaZ1sysVC/AgBJF0crtlMisEObNUyjUQwBUJ56s1OLr/JYOce6ozEAqXp3zv
Z/lufIZDMW0GsG88ht2wRr605FwwUCm6reDl3MZcmiUzQAfoqcbQ0OX2Nt4ocPKCy5/sCDdphC7q
BYwK9InC8QIdI0b1LqrE3RWRtS1rRmRkNmEEEvymaFvUXnHBHWVNqmXevLYfqyTWNMMKThh5LGrR
y3HBUZV1YNixCOsEIegPQUhcDN/CFmmy0n/6fTd+hOFxaeQYzTtx+N/EZg1ayfhoWGbaOOlYhvWy
76zG3dCHk9pjwmxK5COlhnviINpTSq+cB+X6nDzhcZA6rFeVO2z9hdW+gqpCph8DOEnsZrcbKjnn
c0q84H9Hf5PpijVPoH+qHaPJbS8WzmjyI3Rhil/IM0L5zL6HvEL5vNCXovUv5xnOnd1IdpRjVcsd
SoKjjYM4KFFFFipI0QFoKL1yg3TqSGG0QmYP1odsDIor6jd6iYSEpC72znBd7eDGWD37cNy2pYHe
nnV08oduj+EOs+mTCCEvVvz1hXNr/P8wAzGsJToaJFL5jObLS9t1dgTa1XarOUoF88P9cIX8i3ch
GhTV7cG0f+U4BDCwtOewp2NrmVkvWzooykSk8WwQ/WhB3a/XVyE1FVFYCUo9gNWyWYrZwtBQURKC
hnLGLA29wFGbANLbaZgR8YBMFcTMwL8z1GNIkMW8y7esZrRuczj1xhS6kmV7S+rBuRVt3cKx6eM0
0cDOmQJI0XS/b/iy9Lw/C7Jx1ky+1Qva1zy+RduRNwHsz5IrPZK3rgwyB3yqxxduxNXQm8NH6bwV
2QNuGt2PCg+zjkSaGZ5RYwPd+URy6Iicx1SKAmpbd0GDKrMxbADuJKtxXdP3kdxBbn5BEFEIoMU6
fzoy1jVdG0ILHLPw73L8PYiUT8V4lp/8Apq3m5g41gjhTKIAe41kY6GTpHywtM/5/jxZAvk8sB13
dSK9NmWk2X53PmqhN9PRZXrLcDZzKghdwYZe+lR12aDx3nZMK3qbEwTtSbfYc+UGP2OieRNnWheJ
C67HXajAiueBXFyBRXYq/ewVQJKOrfdc8zmQZOJ1tHT6ztduFoNhsJfKhm4+CXE20AEzeLO0MQn9
J21zYEIySVfenS0xJ8ctYbcZKTVj6YvtWaaxPHL5yKR4h68GBleawu1De0Cy8ndRKTb3xUSEOiy0
FEGUEUOipcil327wrN4VjAse9QV6P052kSA0yGMbV7ABcXbO56TSirnq4ZAuj3oScIZl9fRTZPWC
QhvvzwIBSuYVXls+wHPZU1H6BWt5mr3HHh3bRWjOC5o4eNWKnMbemWcRHzmNba3R+azelPiHT9nK
27EoWUo2AppW+rSCEykTcUOWeYtBlwnOsYgmnjmmT8+RCWg5me5E9Bu5CV9gDKtMV8QGbWGNGBZz
fFCRXgkAH0IxoRtwyTBxY5raNeK+hRyTkxsc6RBst4bTczK48bLuAETTWO2aKCYTNbfbIqKqzWOV
WfNYtK3XMsn4fswWB+hhshiy9xlO7rGM2iXQ4ciR6weLKecNMRNR7qAunKBXFwJKb7ibj/m3AYmw
eglv3rxbDp84uw7voHdhTtrT913NPxVcvyhLycOVC+/0yauIwzeXweUgSI5AralVxWLv6yIZHenX
K1Uyoa1lWM3hz/Eb8rPFZsNWAdBn+3y1IvwjpHlINqr7WxzmdPrB+Y8O70iyABVV+8GYdaiw0KhY
/wyfPRQBA+F0HWlyD3jc9a4PKdjwwjEdYxKy5yYCKX9YnJkOTzcZIsuuPQdgGcWwlb40fmTzO3bl
xMyavAKY4xSOaPNRsq8LZRSN8M6uItnkxa9kI1Kmb5CnFMS2XfUc4mcqxQsRF7Vqjh02mxg3GwpK
C4SyKPoqlWvlnxMNSUM/UCjFBVjLwdPnjo0HWPQd4b3sRIC/IaS8jLa9T/P+4wxxIKHJenkEl8ln
2iX9wjISfbVpx+SxKq3ubwWlMyHRcRdUs3nlBnnkgnW+QsRA8O4o1WnBkexwcpkKaGQaYBXqXkcB
cqF0rjs1/hL4c9Pc7cytV6mYj+t1wCdyD22+Xqc16xSbK7I5xz4dSkoYhehDoM3I8ZWckCimd8HX
I+ELXPYUo8POfJD3kMV1jfnPqn43CcNn1bk3UTJKNq7/O+9zM2vZv0FekGD9XmYDyff3k6tAA6YA
JT/5u5oDT89cNNL+XG5Pt/6eRJq/1azXgyjbx+DquO8hS2S6jvhAmtkxG7VDh+nszH25WoH/0uI8
ufg9EcZvaiLSgmAQilpVbdh3nwjtrTLcWPRmkRmICuNJgxg74DeBc73sBneL7t8sh6YRh3ldxIFP
hWSjDlGq7he+BlMNKkXtvvatxzyNajc7pRoTyHneWhYvTUP/Y48Dsk5GalSlbNp7pQiIyjKqIWv3
QgjwdsAaERgYYMcI3uB4bKNfqd+f/SEnhzXnAW0ulgKgG2crsSVWHV+3+xHx00T1Qmm8/ePlc8qj
8yjy5e3wDA2R77IbztPlNKOJOjFnTFrOhMlcGRrbc9p9aH8LrGJBiuF9LdhatPWl+aA8nJM5nub2
NrlgU3BW6gY3Dro8Is4+k7M8IuxB5EzrzTd4+OQZop7FCvTG4GmiwXSIWIJLJvwC9TgMKCBc+5O/
yfT38/F3n3aBxJjh0NIQd8XdVM6ALUfeq7QJXbKeGP3R8PcT6RVNJnMDROldV5xZVvPI041Wj6qs
tUPvyxS0XeZEBkTSjnkjZYDS9PYzNmxWXeyuhOG2dBMXhqksx4ILmeYqoQNY1NK+1SrLZ5DTfaQo
AckLFJDiIiBgR+fEC/rVe7E0l+joVmQYrJXolECypgzG4nX41+dJbK3OTAKnRlNsQlVZrOYlc4rV
UpMK6Rl0gJes/qblR59O8jA5P05Rl9zSpW+eQHWx89SVg/4fcawdZdLQRZBnD46qIr00dSZeuIbK
s/JefLUty47clYck1G/EJIqWRiNDarToM0DE1OQUFTPC/+NfzoKzzszFQ0a+S/iImxT8iKrM+3f9
gwOzNijo0XhQT3LPrCP0YVYYPC+B21Yg+TEUJEfe0V/wFTjLsdBRKZLHbOKNVKkkqJfAy+JIvDqX
0RSznHzhfQEQ6pqqSlJGTU9Oyx3GtYzgN2q9L2YaFTZIY5jS6v8qFwG2wBeh2TNmkS5zW1NWtHPB
dfbliP1tCimeCo2xN4JWdCP0npYzG3burlmF0c417qhrgPQRkR6M6ksKBmTqH8HPHAqfMIeiHrae
lXXTQ5L/je8zZC2WJ/vHTEYtFffYXsApDpguiSftQXJXjpAgr3PWNMci2bNVZmXt2XTjr4nmyvft
YT3LZDNAaZs8oJZgWezzDClhx6oNw61Dv+dHyDSpi0IsvleSLrTn97m05KrIn+OKut29UAQHuPdS
5TmNiill1mn4QA5l3Ak/Y2iDEjLXA55oykUvXonpGm1VtOdxIN0Ol6/z39Dy1h1Rk8Aq8MiYynkh
UhcJUe6ngX7IU/51DiLtCKM949P3IRe/re7Lco8AUlknc+x5NZzDlxFKm5aOSg5JILS+LSUeESR6
r4rPB0sx5Qo5/FLJ2UzKuj5qYRuB+X5Bea3K3CQLF9ouTmopH9IYUkbOif0j2kDed9tIVpB6SG9F
YIqYYrjNRx2d+DI0AwST9PBAmfB6TagFvc7Coe4tNdW1HBIon//dv7z9kpmnwLOk5+bGlQKgUTfW
4K2/Y0xeTijsdnhLR/VT6GkcHwfrFTa6TaClYbrXr8sPbXhK+M0OtRs7PmkSJty9xUMvh8FRRAHy
Wj+hSD1D6ZbPpwLxlRNWXfUtQdM2+uno8q/d67fQE4CWxsvKl72a3Jk+wlPKCfOQ5IR2fYzy944z
icHXH0hxy8tTfd2yDDPRc3bcegi5AmXN3jPGZZD3sf4DSGGsX8QKx6NOIaNO2CNl1lQEmtHHrEez
pEiMIfCe0LyBiVyviQM+ywSzIyPcpJKw8fzeMb6mJ/1GJn+iKLCie4nptNZnuQmrBr6A+Qy4XERh
4DEyYVoDyWZ73qemur0qc7wYWXyVkFWYe4dpNRXXFslCa7lRk26la47ahByCH0zvbEMjhNHYIHHY
eLP4WFYert8CDD7kwo+kXbAgcRPuHZlEsdD9gQ7D39ancMw+8E74+1g8lmmqn/W3jTpSMyPkeZBE
zEiJgdA9AqsJ947avic0UJ7Z7JZf8EFKrotZbY3OlnKMX4rKFIPbRvu5nwkqExiQ8s0YJwccrWQ0
RaE6FlcFuKubokfz82kK19NAMOQfRipCsY9vfGmJAoHQir3KoTWaVx6l1RZS4Hns9UzXAWTtu9QW
96ntYI97cNUBKFKoLrqiRHXpYaXPCrb8ESQpdYjagOBN/jFM79d/MvmMvbpbt+oMvNnc7vpeOxE1
eOMV04KaIbx+GgqyuRfxy0Q3V1phOy1E4xcKncPA/Ypn3m9RwOXBWxrRjCmo1ziR0r+lgCo2fsV2
VIuWVrHy5aJWBiV6kw98W9vxQDP209FKS2DskCQBZuzaeXNb7P3O8uQp+j+8E71ED2Bz3FEgS4DP
8E4mL+rmkN69oyjDk62tvBxWh5Nci3iQt4a8n26c9rp8oq0TXJbQUWp801pWPHKecXzdyVNIwz6k
WvT/e4/uTL/gjtOw3hjbb3K/27n8xfhQQSOKVTCuQ+P0/pauc9c2cSSCm7lp1Nw1zDJonnXCEFmm
5NBU95JSVLoATp4QENu2tlDCYxUQlFOy4B8Th0hrQ2f5juf8UxhjZywdPAfBwBXGoeFnWl/xOAWU
SojpOkmithKUo7uk5fwfT0wdMXz9ZDMImzAJfAukrF58ewkbDRyBGnWJPs80ivqvrEhvrERqTGXu
2bgYdAEfj4v/O9GOdG3QEq8HC2XiQqFMRHlOCZkdNFl6PSXSnhm+132AKarvDIQPSl4Nj35ntZHA
BLcGLTKzQeHGS3KXFUGOH37epocDFQO5F+isBf8a2ZoBTTSk4Hw9LKwgcqG86ElaxT6Z4+Es+r2B
aHTWXAu3PgSuOZj1UZfbMLURNCz+kbrn4JOemUGbkdA5h2K2h1yCWFLxtoDIcMKxVB7aSsEvxpxo
pQau2ZZ0kS5sgAEUAKhf7a2toz1TQkpkdNFgIPHQ6DDfmcRtJIT+Y3OnKtg5FRmGxV4YU591ESBG
FcmUu5PpdYQAc6ZEXB2mVFqBUGi2A+Yzh17t32T/xiHGjit6KBthsmmG7SidsiHX5nH8t5AUq2w8
w0NA0ieg8qot3Vup2M0cietjFdkVNdI76fVzbQD3yngozYm+Q6yMMN8dH8nUbxOV6oSoqHh+XeMu
+XjYjqwsqIWUr8qx++xf92IxWQTHF5skbHFi/oDUbRDUbsTROCTHyZHVIA/9rhSICPkkWXQzNc/B
hxyYKdIXQd0x4qaw05cx2nhCnTbd2D8VmyKm9eGkemOcdm7pivt3imXKd1BltmQ7BqmzBQa2y3t7
3p8hTB/+5h0ywi7w/G/G48f4fus146DvMqNI+SVX8WZjUIzMY/9W13G7rdzmaoKWJWe6gnhE+X8I
Prhihk+jfpwjCZgjiPHWaWsZqeP15OHf7U/YmXOZN1m58KnO42vaNk6QWkdYOet3c8b7a2Syusx2
ickng29tiNdFfgNeUQrDgf0GbHyF1PexwQHUAIXo4RxN/EnFdVKsRHrKMBEBJv4y3hEZ97tlqK/W
oQA4w2vKC0Trwhl+NkvyTJ4W191AZ9SPCQHxBcGVYOVQ3RB56TISqPJZMrDT4zmyxcIWvalRfitX
jHUiVky4OfSJEOJ6run7hCWthfg2PMahLHBDNREZZZKTZy340DpBF8zzs5MOYE/KFCa1lp6ipXGC
HOKheqtCt/iqSEl/95++wWU1n4pBVsXOvW2T9JZXiWqr8sNcpcqD2Zl6+6/kqX9UeUN2hf04C/Hd
Rwdf4ujIptpMEVWeFsClvWTovkvnjkugd+r6nf1jPl0yJwAZdFeXzcl2yFi4jW+XmiqWkGZEPorg
o+s7v+jBHcJb8F8aQYj3yOJY5ZUYXt/FQ8bfSUe6FeBvcGw7lg135+nDYyXwpAxcWLU4W8tAmjf3
qB0TkRiOT9xYPwlCV0EdduoUQU08FDdd35heLX28vhbrQUOOwH5tIljlxuDL3wr4iSIyHpq9Ns/B
r5H7Bm/Or1+VJGQ8ySOHpavfUM818Ao9emvb9bH9a5RCVbG05vLOctzfAVuXDd5irsMGIn75A13a
Z6RJ8T9GemnZNL0BtWYYNJcKmOx3Qe4gBGRZ3zdhJ/2eELyarx8VOo/N1B1qCn0ytsSG2mqnVyb4
cpwVhdHsz1gjkBPjIiOOhgt486rNYux/pEtlqN+z0YbMGs1mnyIvuAezjPom/C5w9xFFU+w71wuR
UcBM5OCbyrG9O6NLd9ZZZ0MwStEiWdmDVTk58ZKFDUAExYCl4N3Q3TaaJADkF6JXjEbIeUlsL7ZJ
YoTfm3UXo4M4XP2R3DzBQxu6LTVBaOT4KiHNRQbxCFfFqTs6MC2jZcHFRqxh1NBCniE7MW6IChsZ
Ftll2mJfZJdgDQzIrk7ZYCAxgQYGlMsc8v08OGjkVhP1aiueTwdpgLqUm5CkGCp9Y4s5EjXOapjF
c5KnTxrjzC79BZX5gW1/pIy0AvtAVqArv8uteVfffUeVBqoagBO5gV8uAgKNo3ZVWfb34DyW0r72
rLZ6tmIfbK8UHgW2Fqh9Z2wXVsF69ds9T1yZoI9woh8alGF3VgOmrVXjX+C2KtjxAJRK54xtLF3q
bS5yjZpr6Iyx2N93KDicjKezABedWN62ZlGJYiqxBXQNokosqD1nTzrI7iKiSkXgu/ntGTYiNgwC
UyBcD08yYjJDmFHwzITVE34wxqUDwzby/zQalIJ/9+Gx5FA0TRWerQFv14fhr85L3RIB2KhH68qk
/teXsdtULC0VZhjjRatJbbT3AHwlyHRS9lklKMGp6XG4P/TmgPkKDVdPalQNa84cnv8oSmmejt/l
sTS5S1SJF2M6xurDy7JftVQfiI0yTr6QHr46qH4DjAyNCTdEk7vEOc3GjKmp/wpoqlZnPSoRahOl
R8xmdNb2gL9cweRwFThK32YtmtLv4hGZGtonQYK6prSovqpjDnkGXQvMVoTutFk8ixwv95QaurmM
gfghZNNe+Bsz7RuNLWGJepc53WLSMDMc4vvTUve2tLzXJOPCnj6Sk2Zg8JUgfHC6+qlBDUwh1J8r
9S7qEGp8rvGIS4vLUhT7fwhu5QoduHXNhLsu3aj36IU0mV8d3ivsAzVGqJiGuxMfkpeJklwgyyJ0
a33JKXL5toH2SDdujxZ6/hpeIML3hrqucoC1YUIOI6Q/UhWJeoDjV3xcTAMeV8zNbuPLeYxv7RH/
TmXBh+tA4NHGeGYh0WW2VDyL36yV0hD318uOGIcgrVDYDTuyARVDxT0Pgs/eja2ADh6FKJXjXTyg
wjhDPCzrp+dvWd4kg+uW0duXMSljlwdIOiY4EqLkAAK0974KDO288D3QQ2FvbbqDIm3ZVm4uIXay
+EsIDE1RykXfY6j5IkPmODLKFqkpHHwqCuXC/kVHWxjKuLnSb23FQAz6yeWa+qZ9kXnX3ZyrnpAV
lWC/g4Uh3z8MwlG8HqWmpzTIACmFo8BIWR8T4sflNilJ3SBLL8LC5qhpyz5h/C8TBNlSVFXE8smq
/KotgE6GSXca2WlNUn1bnNeInaz9bnyZX8ZzCtBwQsieqVL3w9EjzC5xx5MGnmrrPMG9Fm4bwwgr
z1H0E528sexNTFPrO31CZCYYjUGK8rm//PBREf62b61bNMS2urEeKx0xParq37U9+db2PJcvY+M3
Vo5lBmcelRTiDas6g4BaQeFafQkoJc8FShCoieQXiJXMvpZwbbE7bmqyO/BhlpF5yAHyGyAnZlGL
stdT4dYO6wXoMqTwB3yFaao3Cp6DGTyRHZMQ2TS7tSZTFL9/sM2pnjOMZ53zR7Vr5iRLjNXu7Dqm
qGACp86sOhCBLLH/N337uWQWyMDm5ZCF/iFZPiWNi34gZSoEuTrZ8VvyvDitjZKi/sJQ3/ioOLal
GWSYS24uElLU7jsEZIRzkT5SGwWHcBVti6pQNONiXVFhppeCaoKJhsZEr/hLD0UMJKVH6d5S63R9
lIj67860Y8Yqu0a9ujX/AGeTwQE4CIw5oDzat/Hul9kRT81wwvacWHDMoSLDQMu5cbQ+moPfcJg4
N6XihCo2EqBV0r0rMcsR98zqlVPqbVplsvyqoN7zdkT15ggf8Q9NaXE2nLuzI46mHdtC6eOGIUUV
SAW2NqAohWlixgvVVMtTpljclgyE/LwNirFiTRGXWFxIWWPZhnEL9pZ/Ctur9zhcEDN9KaFKNake
b6irragZbhenqiu6nsaFD3H19cGPE55vFuFAnw/cWcxjDcU/Wx9RqR7uTluXkOI6h87U4Yv/Qp2m
Uh5tmxjNQAC/iMBt8e+uogD8B/+Raz9nj10kGdgtOJ+BS6uiB9fecNEAsfnnQ8NRHSWoPiUltC2g
vYjmy7IEkLWIk7FY6brKakzma0xPKw4fC7jiHSKDc9PRNPX+GKYm0YYkzAaaCjd9fsZSc47zZCyr
Ku/mkwV3Pn5PxDPBHV/9Q3KwXM7EzbuHipq8w0fEemyotR9KCWvOsQji+GQwxopYWIduOK8yznrm
V/xic5b5k1luaTY7ElQ08dlvB/5iKTJyzrHNYr72oo7tUbVewHoWTaR/b2yAWHwtPqHu7utnVDfq
eC7eJuJG4yAysYVYv9cOcSLAIPt/W4Sd0TrCuzHvIFoNNA9pqLNnR8cBs2ROX0fvv07zVjC9X+Fn
tHIVNfdCapWUKLLtBZRbLHfmfI+oCPdd1COqec+hWw2qRgKFPjGv8FVtpMLP9bplgnXKeetyynss
397vgqGfKBxtQAZvCsnjvabDZNIn3+1wxCE8syyKkkbTuizZLVdxS0zDr59nF04qV2Ps7IMrdcbK
71HI9tlMrHICfLG/LJY3F+mxnjtrfHAcup9udz00BEwWMS7keVzoHFR5YKt6GJ7a/Oeys/5IdSS/
Nd9BjpRWk9reZ/+zLMGWe65YfLZZ0kQbIO5/61kkdEvLc4dnAsouuW12IANllMrbAAGiNaSHVEwv
7jrbBqlcYw0ycFaRASlDNlbpoF2z7jZnR2QCXerCp0PtJ7436hienwaMpZVdF44xG6IeuzRjVoQ1
2/9Kq4xmYgerghE8vMWVw0Esb1SmOR4v5k/Vk25UoNT9JIMXZ30VH4I3h0kxrF3yq1G8ao0vIB0S
Hwz2AkRCeqnCHiP7L1UBASnJxMzfEnx6Jv6AFP7bYdnYAKydWd8eU5L4oKT7NVGapIwhGfSo1KD2
+4KUwGpj9AuAPNqa856dnM3nfzS8ZA4sbdqv8TrxXk8hOnco8hBxo65cwb7S626Rx1PVFk/s236d
LUWPemSVcN56LoCZtbHtzH2cc3Fzj5hD8zS+FimQDgs8XV5WI04CzXMiQucs1Y5ef+2r2oaqHIRP
O0z42cUtiOaEAZelsow3Raq4jv2ggZA2MJ/u2P6qv8JOrfa6YODMsHFQgjcvudpg2HNtq/mKabo3
Ia8tYYxPGHWHHFVUaXN3IVHIL6wJYhl2XEPQHaEXPl9aRguMcdji37xs1Imf3G3boBsoVpKWUh7H
GNLbfQVtCPraHyZ97QuvS6GyEJL0uwHrQ0m9QXm1ZR4vz91i9hH8Pg9+hhBbqzMFOPS2SsOb6OYI
QDzYmdsT5mf3tDN6sktTvLBftlJ7teYkUfnxwN2yezrj6upCz9UHBKrFA9MGzSWHIzFIBtqmOpOR
lYfULH0DgjsXSvLuOfHgqLRB1YjScDz7UUrcCQogWQgzSHt+DtzUmETAhd6alZPpSANtBgMRojcf
UUoWVs3ojYP2kuGh8NXD7Wvl/7f1aOUYjMncx4kmEKnCMPNPHwIUyAuR9AOUqy82WyId06ZAf6gw
0jw7ceWor5OO9DUW/e0I57h9xSN5Vcto3UAvHi79lO1RFdY2zbkDpJkSroABZturZus18AMbwMT4
2dvrBfwvXYylBw6imMt0vJu8bZ5z8JTZcq//A0fkFhZ2X4tQWIorii9Ug6j+BpXE+mHgnWo6XROZ
ctnOlvh0wWV+7OWrusSt8N3Z2nXFf0G3kHCCEEt8TvEBPr+tK61wkT93PF0fznkP+C9Q+9l/vChZ
rmVZN5ATulOZ6ySA//R5a7L+ubhHNJzMEPBFjQ6g6o13ERsbNCIqrD4IVuQZuuz8CRm7LOYDxsl/
t29cxgC7/sOO8ScNU0k2x5fq1PZB3LcoYktWrJlhXa6OF4dd7DRFRY29fgWzr3Eh2NBMoumlJZLo
DLHa54heUfOVNkdFQ+1eDFuotvKs/HkAPPbtoAopJSF22NqC8AnM2toBfiIKLwQ2Z6A9yczhiaX8
Ky2BIyhQ67dUesn5Hk5a3IWmelxBrWEV4kFSTSmrTqUJ5sT9wc4LCOfM8TdVpZD1cpM4bSiz/U/p
sPgX/FxZFvc+9TkMni8/g1jw/nOfMgckn/LNkUSk3lIFYBM39xWzXdYb1WR3MDBArstUvnkry6z7
9ByPWpX9CQIfLFl1JCEA4P94alQZF1gpk2TeJB7JolDUF1j9QXAtNt54/bPgGXyzqbKjpZTLROFk
vLsFqHnnwgrsOfeRoVGlouWCgGHT6XAEgfVdiY8elJF57L1vCXQualJQA8M7Fa8V28TY7tFqqD0L
3H7MwX/jOfkBeDIhnpO4iWXUxGA7fmeuTICQPEK9c2rU0huf9LB7MW1JnqA6F1P1rezcdWgMZnSj
m9lqV9JA2H7wcxlrB8HcwxJg+SvD4Ilbe+JHhIM/7K59M2N8LEaFj8BijPAH5SvMBJ6UuU5NHMwZ
oqoeuAuTuO6d2dCE7tw4pkq9YdDYux4TW7QgECV+mTlx2tMeopKb3ENqpy1PhZGnTeUNChzTxNV/
FpJrgkaZvI2JWjin0no2rNwtofhSpwzu2lZxmUVndPtqQzUcb8YpF1/nKIa8cGBxPHTEOU1z+k1P
pb/PKaFxNvFwUV/4/T9GBUj0iMzxeFTdZQ+mTewj5w2sHtcyjSwIAJztUXF4c5vEcqtESIcKPmuF
R1sbRErp2ac0332n3qhsqAZd8kyHHxu6w+aR+GFM4rFc6TjpVWahlOR1HqzBzcf7DaVpsSOdm3C0
Fhx+Uf+r4FPkdUj2Q0MXgbTnAkfQ/h2/gPAP+a18K8IiTBd9J2mrMFfZFe9oM0cNHOuDp6w5F8B6
ygmP5990LcVYHOoCh9NOxCgSpLX+Y86unPSU9ORe2OBsjX6/HbHtxUEbo2iux0oPd26bPQDNspvh
qOg8tVsQS5lBZqizTIAZDofwC1svPYXJySy3XWIxxpI/myOZb+gsOmsaC4ddCVdraDlSCA9LPkBb
hi0ja6CJRqy6FLmq3oQKdjxJMdq4kkf8fRlqfLqDcFUelqPZKIWg0xfi/sLTGPSO83uU9ZrOeWen
RZR8oTIvBRb7O5knWDQIxlWeWepfD1kf+p/5wy4Vg1u/f8gv8+zFYkSeVRqZkSAlSDO6k/FrgTe5
CnsGwN16QNy9Yi8S1qFGpiX6qRmo3vvzf+8j59K/kVcZZ/yVibVk368PsKSsfJ99KPt4TNnsXY1b
FHsaRTWry6hkfm9V9fBrqLFq1P5wcsXWYJBPMqUu0LQr7/bf3qZ+V2wtJMNV0UCbQZRS0F43geef
XFb9Bw7dC8aflUP66GIA9AMIXE5UQApOrT1vcECI3wLqryL7n46DmABxjv7C4+UWwEA76WHJDBjI
i0k7nB4cfHNDvWjFUE9cTt0xlcYYfKsASHoUy85NG72tXn07Pd4YTSP3iyWuVxA8jEL/lg5YN09l
M7FdtMxOpkCEfyoe1L80MXVXdZeZqJyu5VW4Hsjvv9dEmSBoGr4V8AEGbFVc1Qrdk+29yizJ9Kli
mASxrfd3KSjhDheuM2Gf1lZfKw19Jj08cydpVpPrnUx80UiruZ2Ud5mLc/IMNNRu9cdK40qjO8mo
Y47maoVkq0/DAPfnmMhQSLQFdaPSxRz7AO/wPNIhm0rKaUYiQP+Hs+Ogc6qG1O5ozd0ymr6xyyJm
N2CwvOdy6nfJXvQRqsgTirk+cTNQVLxpbnDxxc8fos3sxN4AsXRaRsHiqDUJaXhvvumDKxvYnrUP
3kZMCjHtAhXNqyhumaioSXaamA6c7LDBR6ZDGhy8cGz4F3QWlc6cUFP+EoLBh8lMZqSOBiotpuCU
qsnNyozSeyqKLTUzfJ8yQ182ye3ijY4Wlbdgr/KdIyQhEvKd4KdFWQdTDJAU6OHrvSKyYVWDKPiR
+FVy5oSyISryxaVOoBpg0T2BpLUWvgh47JiHXk3sXNWxU9DWvywrxF2PxjnYr7RVY9g0JBSjAIKY
KsG7jcppX6/NzYi595cX8aD+JOQjSQo0g84xBxbW5qeLB3/i/Ejam3PiSi5VD6W1Nb77q9SZQPtN
smKBaX456EXOXsafedtjp42tlQ3nEx5SJj+nvFMXhHZ6WYGysBWzfUVmKQUKfnDnL5/LE2qJIe0h
tq2RoDrlz3LJ/PE1UHrBSHo37lJWeOKDso87eNcO3YGiZin0Astz1WP0/GeYJrvIUg73oVtlxgsT
7P+pIlrgjcVRCwT1xPoZDeKEcQ5KQx52DpRIL55Hu9izr31GUk4GVXyeVlznvZa1pKPzPAUDeHIK
v+WU0eAxNQYv0EEeGMzu+FjF4jSjHQuopEJKGGDfg3KJaQrSbhioeiLsPyYEfdeELkaYs1epsKR+
70DTvF39U+/Go9+O0ZFikfG2ZEtm7puRJ6FzmUnkJbRboz1a6f0qKeFfTxvoCzSiFCo8yt+sFiwM
LeF7bJksdbhscQ+BdJ0O5P9OjdqokAAA/YmMyhJTRprdGQUubnwMHXvLvIVJuJxOX15OCFKC6l72
2m3AdGNLoXlLO6kTEf4d/VVze54p0lHv55ET9+3LiYJnYfkC3oXKhpMrwlaUtNI6DMJo6E1R6dUF
2C6V/k+f7Y1ZFnVv16W+ZERxsEAOVbsaRaiWX2UPVS7IU2fBKIEWhlLyUcDAsub3l6T2U+KlQe3F
iMtNVsWgkz7QRZe8PXag6CyuExwL8DC2GHZ6LM5+e4UViu60PjlqdybubIfjt46gI2gVH0EXm/ew
d/EZsbMJ9bty3828i7HEZUJL9bN2urgQBYmTRNs46BAotKKjgrYWmnftCrBprdcowaRe6q6W1y7E
Tm/YDgt0liakmwwUPUbSJ8XbTOnw69r2GkHRXqwhk/qySFyfsNkbI7bAkqCBk8l31BUYmvKvDOmD
k9uUta9A1BkwxaDrqhB97YG3WcmfqVk1UI5uYpeJWuWUxl9VdUpyLqGQOP6Rv8Hu4WsEs24udjY9
toCw2bZ6A9YtQusnROOQBBvkR12aTQb6MHCviGBi3RQxM7SMnvvoWZIZ6RILnOWMkhho79HOb6wA
M/RAzedpJ5Tjycd54YKztRuhGK9nO2pKuL0isy6FZhYmqnDnAXq+yNJtYHa9SEKrsP0978XzoToT
Z3Wf/pBg5G7xKXZ90y/rHZOuxShTh1xFcB8hcHhofispFxYnCkfoDTDde+JIvCypELs3AeojVvbm
yVoFZZEGBhpDC+rDAfhC7iBSmR72O1t9Fr7Y9uKLZQNp/Dm2tL3zajNBEKpczZPZlZAcefAUlnUK
8aroXuKkRhzNUXjWJHcvMm1wuBpX46O0fnjrjSkru+HgHoPbCon4TbgTnyLbMO3RfM0++YjiVZdn
GN94Vsl6YsS33Hu5jxkIKsfXMtfYMXp9sduT7nUvvbIuW6Q1z2YRgw8L304aem8rJrH6UTfCOpzw
upzHNg8HCGLN6ighSOEgefYmGBq3GIkCqYagip3HMa2MlkuU+gqv+wn35eCcasosuFAHajKVwINW
tGifexOXcbO6rDD/oGNBGOnuVs2x6tP0LzefmUkCi2wZsyOKhtWHAkzpCqeyxkL8pwbiYbde8YAI
HlIQ++NqfuIxlUdR/557r/cAiLGLeMFGAfYhtbbXUVi+OUHpkE8Yu5DnjrX/BiRADqy1ZxYR/Vhu
YF3krb+ykCJ3ua0B2pYiLRPaqs3r++3M45cqO1UOtOc6XMX31tXl3+Hm3SDtbCUID7AWoqJSf9ax
02IpakrPqurWL8sjednBpDQfWKpMEHkDZKnin1DffcA1mtGB1QyZ/rjnaGhpMyHHgFeUCiQXzJ/C
vQxclC/IwTNOxYLQq/l71KM1mou8tkLkAkYwZU6p8Bhei9dnDNTfNnDuNrOF881b1em1/1gVIqxg
dVFiT7l41r5D2p0EUoek2FRbdimPjgh1xYOlczeImXKla5VAP+qLBQ/HKDnx7/+s2JqXKjA3BiC9
mGAuAx0jD2lpWigzGMJiK+gTOqxsLC5CO4bA/v88jzyTRQ33wiMXdcag62DNTwIpvAkvLJKlPWsh
6mYJ/49yPYXoNQij70HKL3lvgstyAg2/8v4f+zoM6R7BzAKDJoLcdwAJhB92Dnq8yyQHkJK5H1ZI
63xGOA0LI5rcmkH13CLoQXizpXCd3gOdPbn5HYjwg8XDu6cyFJsut3hoCERngg8byzPwDQA7tNAY
mNBEh3hZgd1uO6lvMgmUIJGpNmFMS77j8FxKsJky8xKr2w7qA+CAG/9m9kiIqlo8vbBesUXBv5ab
uVmtFHpuT9rLrH214CTE0OrZ9lTmACypC7XEnXDZ7sdMuvfujvHAmqFmHdKhbDUyht0awlqay9IJ
o+9xrUk2DV1qUSo3f6dshtGoPVDCCZxEmFXjFG+ESycHQ/icVnhZcF3WLYgtVYoNvSBqESsuXkEL
/xULS9C6i0vJphwCOUFKfM6+d9FgD9vOpdL17HxjyRj5tZSXgdiQpZ/KBMJy4qUtuUEI7200AbWm
AO8QUx+hNS4vfctq9K6b1Z9zpoYre0u+Hic1yTwhN+/TbChXVSgXSaSg82/RK2lX3m1tFsbldfeL
F//Vvgyjs24pyHZg0cbAZTFtf8C6dSjSCdw8d2x+xjSna30TAulv2V1aZ/xZiPlQRBUnMT2gPbOF
s54Ko83pWE2uugsRN6CEe4MmKZkA2wKz521Q8MOOQ6okvujTm/0j/NYVKGnJ/2H4Jf0WcQJf14nU
QXPP4Yx2cRm6lEMOyiIlPnV0rskDNek2JGRvf7oTVow6eL1UIKaA583Car3j+eJVw8UAtznHF4j2
/YFuG9MzmbwwpCVojAdrtaiciIwwIq6kzfXey9DRFh5a+yqOqg5H36n4yXtg/e8xIK4MHLWUpmZO
Mtk2NE9tOW+uCMipSiFjwS0KUaiFkf72I4Wy9kHyizgahS6iiap1h4fp6TNR28vUS0oTDeteno1m
YeHjoV8Ox2OAd67r5mWTO/J+gJyP0x0p7PxdzPMLaZvZXcJ6W6/AQuDgpkjRQUhhj04yrtRtwB4i
vvUL0E05rxlmcBv/IQ/nPJfkV2GDRJr/9c3Qjdn5SWa0fEo8RNV13FeELSiixvsyBFysCo7/n9px
aWRwZcmKH938CYTfeYwNEkI0M3DniRiQFzh8Ry/MWa0NpQAscV6uJ2X8svDL8fTfjsYjWxW/yVYK
LRwmbHOjvrwNjsyQ2brKekRUT5zu/n6KBME4RHgggRT3rXbTpJSAQDSdy9QdwjXxJYqr9i6Jb/sd
KLsMiX+JP32LbjzdWrFpTkYMley4BTHlcEvS0kcFkrl27RF7LoiVzyc06E8umGk7UI4kt+0XioRl
Q95HqQT5VSa9LQnppQcsrK4SpUga7nC8EJO8qXxWKusKuTmUVMnMkWpIDHhECr22wFSLSYzrdpbK
vUu7Oh9Q3bw40jwlo3yq7q9gUY2uJK5e28r8THPBKGBn8SDOv9CJDETX+59T3DCQd+x0fsqYvs1e
k/b2a9faeq1OXGojU/JAV+/FPgNAnY1kThrWSnboE+/fRjmOCfXaisEDGLfeEiRBS5WS3StTT2A+
sa4j2M3MXqEwYPelWTSVnIrPNuNOehJ+529GmNlQwKl7IYHKbjSS9kL/rHCaZ+5WXKREPr4+HIdE
CoMBYTta9qBLoqOYyKTY/4nKo5HipFiWCo6nAG399KgEGBC/A5cXGMSMwPWlINin61joe+H5yNyB
CxX46YiJK6qjquo4PrY68IJiPxS+GJvlZE2h1+BzzWOeqpSpPvztNbwTLy0+FIS9KLtG1X43e4/f
XQ5abaU4L7Gob4ysLZN9f94WT0yNUs5LQFS9cY73tdKiFVpUTqOWJsLQDAYRS8dgAQlNtjiHWDMZ
kEiwlYAD++8VmE5bxfeEE2KSl7wOILinBmP7fSF2vr/QoMR6tqRyv4jS4xKy5Utt5oEWZI0gHJN7
1jNJbdK5QA2k8VsIvQkmCbqb02mt6WZIhObjvIPlfCBZU+u1Ihq49AbVPLa9R41r1KWwjDhnfRZY
mVSwxBvyWxc93t5iPudoTFPnH9U27x8uJVvdtbITnyYhvEapZD8T42GVa+GsAdGcZYaVNAsaZezY
+amebvZ4wO7L0X7DpzR5XJx4dAWAJWZ9fXkAmI6/l2VN7a8wJDP40AueOBKQbv/E4Y1TLKQivDZ7
2iej+UylywSGc13rQDhwsniyRFVl4lblACPDQKYR6GIeFkLTfaBR9cx6wnFTckuheRzwUHeVUv2v
UNowgZUTXa1wrAX4qk5uoTiBMgrjKBskHkhHmYlY4APXsHj0V6setHIBo0cpNeVv2AtIs5sF8bAp
LwJ0vDqk0cwSWdQiIrmN1y6TXZrRGVin9uNQe/kTh2XDxLO0e6LBaNjWO2EeM3RCMkh0MEkOQOyb
Hb1viJfcMMSQumhRXr20DeO/TvYYoiqnrGTpRkvQ+EbTD/jNNdmOqtFZbwHd779jQx22r77G3a0a
H4UCmVp1/cwgo44Mf+bdmep4Q7BlPqN0d6jCzUPTqgzDAaNDexdfxkYZ6CN1WbpRLeQFLsQ6FyDB
qNm6Fs7mSqiLz80xuhHgkyJSY7DFTyPWM4Fo3f7mODG7K+01eLBh1eQONB3CXS0qAgN+e3oL0O0G
eCpXz/AB01SyTLb9xPCqVUIzzsHqt73ugzpSax40OgptIp1eP8aZNgUY4PBcmfMTCN0FI5VplzLi
KB5vhphsnEzCHj35ocrrlY0d3vR/b7a5sjaLO3GZtWqTe2nZlbsxZGX5VkLqjBjiBaalq5SmVoUE
v4kC6m21/Ty5pHct8BsTzpCBJMMGpm8/Y6K3Yhxwm7ispN+hePNK/9uu9pRIi5z3J4ecYkz4nJ9v
oFWSVhDVa2sqA1Jbdkol0dNHFYKvuHQgEvzyLdrQ1j8tsVPT/0sgeqW1eVzAwWtCV7M4Fu3LGvkC
u5Ti3P/qN/SX0R1BVD7wH0AFWcgYa2igpfRDDNsB8G/NwHBHw5IW22tpGGxXrM6x7arKxrchQIxh
cAnTo4YI17BIPSjpXPwX4IfWoDUEBw2+wwhIncsfy20N6Kl4H/uMgLFLBQbe9V7XsCOF5iJqg0Ha
SpZRmdROUSxQAL8MbEoAztMxffQ3oJk3eCXujLoCD0F6yCoL9yL5c52uubGyaOuLmFE7qvsw/zju
S0rzlRMgJtvnr5gtnknZ4zRZ01SF32N/9uAojETYCLRHL9fvLG1bErQ+U1DM/z3nW8fW9t0GnWMh
Bdwfxud0UakU85MM7o+CQCT/BAEeLPZ0VUyS0fo6qSowvVAooOJHyv72xHxoqvZ3AST9uKLf7RXG
TcLMA9XVp8KK+gSKtMPYGXfYzo21dPURE4viW5I8ENg6rBTauzTbBtBpxe4SXWBUf8o9YLqrlLl7
2AdZak5B6QJQGqzuE2chFIrP1gSNly6ScPaoMahXfwl4ik+sUvYPfZ0POXHfQwSGw0IC0TsCr34m
6axJOXSkLA3g0VhLkhRfdtYfCiz/8Emo0q5HP+LZGx7ePXtMA69wzOAGrSUcy9JH+yviCRzGUR8R
3WJgSOkN7rUzZfLRmisewCgiILtkKeDvaBSXJn9282NfTTuA8TlseLXPXVMp6vvoT5S1rD1CRQXi
p641Wyi89lBakHqFZCeHEOIH35AWo0mihCRT+dI7uuJ59OFPDU4In3daE8K66W5dv+pzYoh5yJZg
BB+3efbkOx9ok+2ljPuskc6OUkaJbpHyRn2hDIuKqAuteaSiCkIlK0oOBAPaRiBkPHhn5WEucb21
+rKxqyQdDjOhKPqorzJBxFhDqI1YWC72IX+EX/q2amztYm8TOtU/8GAiiEK94WUXiJjETLOhsG/+
L69O41lawuhtYjUIeFqJVE+tJTs2UgTJV88oDkK1aWcsPsUB0NPogVIrJ0cZR0JG04HJmdlY3yZS
8BO8a7A3+uDG2czV+J7C0L7c2yJw41lI9j1qIMd/GP/9Gvxb98ShN+6mdJU7Dadr0OezoILmY7Ia
/5hxGb2K7ffmGD3VnGR0nU1/036qEunK9fMj6gn8hLauJK4SA785XZyWTBJknxineP5gEO7Diqkd
ETCOd4ZZIF8CifRj6iKcvz3WDgIBRMLwN6HoThPxWeCFkANPyvWmIiDh9NYcTxMszIKGYv+8l77i
HwD53se++sQj1FMe52J+nvr7MAoaW1rMxChnzdlxBiH7SsD57iF3lox4JEH1xUNx7JBwQ9HzNh9d
1f2LIej4smzv74MAy1dnBLCUyODf86X3QK+SuPqPupJ9AwSixrKgIOhQ2JmIItdEJJ6HzXZ74Viv
Q0EaYOvyeOE43bI3gz+rAYnShvk6Jbgvy/5PZDhWi0+jFGuN8tATHtb1Cem1bd56hLkgPdZD2u++
yCCJoYp7ehEjimtkTrzx8LKMNYa6s8+9lDwIoUmCUXF/z0SD7ZSnT7Pg1+Z3KXMvq3Q0LvZng5VL
COoWdV9zZWgesQum2bmWIYbrnYql7coLZ2xWmkIrztzly75TTSxUSb5H3tPQdS7XOK053HZ/ZA5y
Pxol5sGNKltRfKiPGrtngjA1A3b3SKZEcSmHGIRk/Uj0I+19iAqHR0G/nEklRcQTROZCjsBrhwEr
t7NuGEGWoCYzkaIH5hli6nI7jmHUhAYVkev8rvUwGsYKh52SpjVjPzDXhk84Zo7TV/W/jvgN6pMB
I0hFFQREU1HJIRZKP3iCrs1ZBCYVsuzWv2mGcWZ3W3q3uvX5NQCIrv0WshLJofPVd+eNrNWxYum4
1VCq12gGdINj/3JSe/6Hh3lT5s2Z3EWo/1pcGL0IIMemjwiUbSwNAdU/Y7sIRF7ixXJAMeye+rLz
rBXZ3w8akC/W+PxVtMYrCeSz/EAiFsngU6FT1NfiFPV1ITiKKBI5jKGX2CFzBulve/LMwAOq7dz/
oYp4KtN2/KRO2pAU3y1hkvy8+b3qL7cVasS8qy1dlXybWj+m93xGCd7S4ZcKtQhr4bGnqgEE0hra
hpnazHpHvvID6zCO7OhBVeRameHZSAZst+m7x280oBjKrk4Dx+D42jQSLod30nNccY7Puuz3kbP3
zHv0GrA97wXhIK6xFxtiLiIAbPwoloe421h4RE6+HRB7DzWDGOLvY9/WoZ9QZVO5cMrzxwezc9/1
J96iZbFA0dThFtdRzkejz2VcE6yNX0R3XW6fEDaTJaccnqvQrapksvj9skpLvL3JAcYohIdGyfg+
c0sdM/qFb5/h884Y/YrnnnSTCodMcGS4Srq+bow9AjbrW5NxBcTaRf+hUhtxbsiaj3YsLAD+LiJB
TX5ju/A2bleBSVYArcYgIUdSitJ0L5kxmJGeJwfsdBS//oeS9MYT4tqydH9TmJajcH6mZA6oN897
Eq6P+FAjqKlIKDIa7toLF8I/r4Di0x0S6bUurwlI1RCd3Yz0lQhvRPkNy3hmMeSW9uvGxLHohhsZ
sYJ/79QSEy7Zn/2g/kVmilhPSJ9xOTSKfJCMEDOhdO7PgAP3uZqG8bQTN7AA57sZdfTMmqqYDBH+
3GtAcapOSwnL2TuhcSYOcfGcBNvCXiR6cqGoeokPNandRQLpx8ow6dazSOiL2wPd/LFCoN3AnM5P
12AH9cax0iVrQysM7O48hvACKddGlPhPJ84SB8dUpJ2UY4bUca3kIaqBvQbJGR3YkmLyl4zDQfpL
FZi0QmFkoMYI9UqUiIiwWwHM5XUPp+66u3JT5uhLCRIJ0kWJIO8qEHJsT76gRJBh6ubJ9TadRucs
h//kdru93KIH/5WesSTZPXg8ZnEYVrjc7GHEIaEus1TzE7Q2BI5eL88fMLC9pPYAc4gPcKGyQvIt
cJB1UbnEbSIZnnX93ldfpMY6znqxLtDOh6MRM2nGRR1UoijooIZcAfTIv6Kf1GvFypg7lSKcK9a5
GqTOeX18rzwPzSNG+xgMVcVebTYqGbg+jtFQ4gUkd3wKW9EJWY/rZz7YRgvlFn+4wTXqd4Zrkwln
kKri4BDFhKC/BF4+ryx2qORkGx6i47IE6hOsKqq0KtYx0adlPvrJDCjr0RttjPtbjRdsmu3d+muS
u6e1Ld1stJ00160AhQamgBoCYLeXS1CjNF98a4wcbPs57ySzsxR6kAI4jSDsiZpNG0EO0+n4CoW7
OB1SqkIK7ASb+A5K/wM4FahgZ1sDgX5JlEZQgHPmoPSm+rIchWNjeN967nOy3ewqYurxdC8Vqegl
+7OA4pj5aIPNJ84GOvaVmOhp4aS5Wz1WK5u0Rd8L4IpoIsTTOZ11Bmc/4g+Yh/qF33vcYYUZWJVc
V1YRyxhTLMw1ydKmrUiTZKeGvCOVffqhWwABtRxPlvvd30tBGJas01VXNIrDaoYahr91TIul/9py
f2tWsNP2dj9P9W/X0dGwFNOQbHDMsfuSyPryM7xaJgY0olExep8eo8pjsVbrTVM+V9RURurfprEX
Oyf1tLb+0X0DlBzsLiR2tFBiWzA1U3McsA+ZfaRqN6oOiosznwZI3J6YCip5xT8l7FBGbtQm1f5q
JieNP4LSBoaC2GeMqelr2cJSP/+pa3sqFQjC6P0mEJ3BEksIH7wP//phJVb4my/qEkHKMBZ28QQT
nAcxlf78SVtYWzC8ubdT1QUottzTcltg/hMa7KUAoi7ZWkDnZoiilT6C0Mrc2ItGCyF3Bnt4iWiA
pzG4LdhKxJ4d/QY7i+y0mKlBGWNCJMA2+brTq6Eczu8R2O7rxWM4MzObUmzkoA17P2uIfXS/TXSR
IdUtiAvz6m0BXOK9hz/lgIp7Qj00gbF+xZGAIxGFHR1vJkx12O9SLF8AWX6wERJXzPXgzZNMuvHJ
Fy1wQ0/9E1wgTVI5+Vive1FWQaaBAArfqsxP2Q9asXVoyKlhAW2U6T4h35yCkzjCs8RGK9ndJpoR
zyuOqsRUdvau03UvCmFlxUPutKN9vjF1buqspJleDPw1IKx/Yw9SG9v8h6lHI27BxI/y3tm6EjGz
owQ6ux8ci/k9Ra1cubAxRohb3au7dEjsnq0zTILT5+z+L0ggMd6QLoMczJ77L+cnbh9NVqgEDMbP
GlXY6GJET49YXqoq9PHy0FGIcMspxWwejYgmmMgx0r76rwFZwF/XKyvplHpUicUhsPCc9XMTIrbF
GD2D/+q3Q4rcaXsl49cpue9bHPdP3202/4vs7tS8FbYEHwg8HDRhDvz0nPqUlcBULis5EtR2jCbT
mjoqOroghBVQUHMikMGm04YyDG314+Q8s4afs5PYIVe+CHZLK5K3h8r2Xqb/H5obkOJVlZaWI0FY
1Tlh6GWMXDQzVOX7amhjwWBBSVa2d/hbtNjbIT4iPOra/yyKy8b9PJ+4KKRtY9nS44HDEan6Fzs0
5SrNTW9vd+9FDW6P8SKfy2EJwckaKBN+knzr5DN28zFxz5VLRnhkLm+ab8kcSUwSDaMvokBIY+ge
nlQLJxGl54oKlpabW9jv7PJmjZgee0cZJ1ne1xLaTo30AGI3Uq8BuoJn3Nk4q6/a/Oak1AmVtFjm
2VMX3TLNIsDaYAoRxDoKw5upC1MWxAZq30onQhqR+qJqrNdAnSUPXgoT0e7+LKWFGFFg0CSmXdYq
V/s1T2DFUXs/Veo6WYMu8MI2FApcz6X23X+7ejUy8N+GFK6aO9PX8vZoQBPwc4jb9ICO0aikt1sv
64/YcKsvRFC83bewPHSCtUsqJLi8h41fPj9SN0tj4OxYnjFodml0bkegvCF+4zPat/GfaXBgfN4t
bNP3r6L037gh2U6NfvqEbrVcJlbuahyoFsWcdqkuexXA1+bQnLxd+Bbsof3YaO4/K3w/Jr+3+UYV
4P69YprjE2ZZD3L4jZlO9cGkvzQiMJt6tZTjLB2hJ5JbjpUFzwzBbUeYVhz7jc8LzKqi1EhFBUVQ
PZViV77Jv/D678iPS+BtHaDoGOywSo5U6nsH9WfFT2tNJ32mnclP+chm3povbZ2GsUp42aHpCoSH
vk71vU1n1RX8z0aEaMyPKdzQ1wRN5WK3cR+eFAoaiDzeto9qi2MZ/AkixX9ouucjV61/Uty8Rvn/
Ejp0SJ+DAccxkre0O74+UJ9X9U1huujyRHDsVkuF+BHhj32/6iqjhdz9hrOJFdrEspwh2fL+mHNC
fJTnF0IYqF4G6a2+pCtbQfQqJQPjdMoaWB4luDZXP2hTWHVl4AouvqGwp6Z+XBhiMZzvHs+2EmNl
Q07xLwwDq20hLltgpy4QDEl6qcPT6I5xQV4s8lY2qZ3bgTaw1KpAXu3S9Vwv12bE5NUwNq/9r3WG
ZGWD71npqY+cXO5N+grTLUcpNO5bqCXVtIj5Xg18nGPm5p8O0mVCFl+2T/FFQ9++9cnsbnaxt83d
qjzhOGkJj7NSult3O+7y7Oqs9sYDklTG5jXGPC0cfOuYAfOc8M6j0t/V2VOqpcc8d8m7NTQfiemL
9H1L5c6Q72G0etuA3Wdz0hZSSP5RDRLuEG7XhCy4jJjCT1cGusI4unWsgJl2GZzT1CP43BpwxoFh
l0voG0HfC0jGF2RemqP4YLoDZvNAZ5ZHEFr7hiixF+CHxNoCu9bSFoqU1LtiWSO/2StHHsn5TAyu
a3gjnr0s32zRebqOAyqvetS7ck/yjyVX+iEgwnHTJsjvpr3xo1CW3DyWXA6BxmEf1uHaNtxrf0vY
TovqNXfpKzE1rVZvWs6/IsSxvIYLd/jKEf6p36bT8JwgMcZFSO64Mweq/DV7qr9e4f/nR2VflPN5
iNZDk31Q2zKBenwWM84Z0aIZuI/6SOoHv9zJLikHm4eZfp3qNJSo7B7EA9d8YchaLvmt4IQQK9Fz
R9TwL7g9ovXTgCVdMDKSR6cui+LbdDiYg0sZJ9Bt1zefIoZDwJZBJBVQrgKyVCafdcKSs6cG2UOO
/Gdu+SiVUW5JP9N+hqGYf2t2kfeI8oadtGatx1teBTYQsDsZDgvYocjDhMhnRzqCWAK2n9Yv/E8F
qMet8Xn+4yWEQr4bPtrSpPjjU6rjHOP0Uymqmw0KTntReK2AyyAcx85rIFZVYMKR/BdOwsA4YDEg
dgUILMA12EoCeBmS2yP63vV7bl30fk6wdV6hdVmm4BqKuLNRtpMtCu8rrWDUFKBc3TgT/FOwLbJY
YFepBKS4LJ6XVkWK0PJ+UY8olVI1F/mD1Mx8GwKkSCUNQLm+iJgl92otFrfuZSXiq/yEc/ehBn2J
Dr8U8/+F1KEvsEziV3FaD1Puf/wtVkI400emByC4m4xKRJD9ZhmQ1dX3sb5zP2Z7QFfK3siiiK2z
R+pV2bsaPA7bX1ekwodXFGnO2FxEc/UNf8tLAMqMnBqFCKM/NnfPtxIu/HgxPBNTn8qgw3egr7QP
LpbBfH0JZaVFVDaxNPPPX8cN+lbk3KIwhR6yMfqgA2BYWKiya1lIkagjrP6Q6/xlpkIgXUl25pJu
d1/QAgz+n83b25JV57+MAPsyIzWVAJRuO/uKUHbNBixCZeh3TeXmbV6jl1XDQbXhTJwn9B2sHAVQ
wXtZD8UMImgE6CWtIY+gyUZcAnvqVNHCsc5rAoO7+TDqpdTXLOefhPYAU+wRFmMkvZXAHZuMjksl
peiflA6UMX7Qp+MC/F3ZXVux6Dq6Ac73RtgKfHjT3rbgt8B9ZRFbpftQC3a/WYJ3QsKlYo4Q1uAN
slIfM5okgWss2JR4EesPk1pmzQ+ADbQiWZfmErTDULsRtq+RTPkHpEuCxzLSV/lURdYh2JAS7Peg
Pz063f3OqEx0zlbTVl/gbn8mKueLAytTJZsqCotvL30d2Z2Rwjycl04xuptaymrJ5EgTWT2eDWA3
7FsI0bU4Li6M1QfmCdIxXrlcX+lY0oLd6NU9ai2Pv9Gi80mfEAKZ4gExD37KCe20D7GbQNWRl19X
udkteHkTqG/74QaoxoY+6vKOVPD6xABbQA3Pzwic+kPsmjn++llHGSTCckNEVp1Vf+9b3Kf93/c8
QbArvlb2In3qcJAd0SolU9OAOPQv1OEHNDyte7gDw/+ILDXXgCD5tySePThbt4bcUhbAjXo23GyK
kNH74KDjm6T4N2yjfYFkvZd1gbt7yJXDhjT+T1HtGb5c09WwFqBEzTn2tPrgBmaaybpP3BqJnX8z
ADD0DA29ddUyPR85LaMh/Uw5MaBZRPijDNFRT2x8lPAw5U+43uiJGBSTg6mfxZchH3g+R8wULY2c
kMb9YxILoS2YUGZYPAAAIFZrBYBERXwVipwGUBXyTStzKi4lYuLTIcvmjR5FHWQkMSqO7pt36a8D
NAt4/TZt7umaw3BKyfaILg5EXMoEIk8u8mbKN8BEUkbh6LJfYwdj4VN2Lka++L+7vdlKVJoixofg
wwRWIU6ZU69sNR1IZjRQVSxU32eTHP39Hy3lOqxcouWSayKa906my5+7lYvBGvMosm/FFX0WyNd3
WACTllzuFJl2Wt6IVspFxkOwmE5ArsKnbP7YG0cBRr2ONYTHI8OGlgIqhFG+6w1saqkx0ObdDkI2
4Bkw2R4R0A0T7yZe6S/yC0tbVrkdmYsJ+5pDddcXxr0NJYZx2AODnHUavH13/XMt2ZX/jkG5tOAe
XUPvcFOi79cJ6vdQZQdqTTx+WmDDZ5IG89WHxX/y1gtELJCHCupmua/pRyhfzqgL/K1INu2+LWXG
m6jgT4MGkfBaBRWJrx3u4ORbrt6jYKyPzY3lzTVvA0jyiq9jV9I+Q79rqYBCFwPq54Mm37yyTIYi
3dtb2EXVAH8K92TOKsks5Pq89yWYL7WTeIk7JAkuwZwoODgVG/1RMXzFnv1H/pLSdqKFMBI3BBL1
xDO28eZwIHo3hEdPA61ORxjUnp4paXEWzR233d+yQpyY1y8Wo/MOLf0VS0YUa11P/E7lqrSohbSO
cK0UNfk4Aq4FBHPg88ASZEP6AZOcLyf71yxYNUS4ml/8nl44cN2JCipteebzxjiw00AvdEd1YZBF
6Di/B68MOhflQw3LoS3qzS0Q8IRLqy6OfIiUrrIni5/ioTVuZqTcvtTRowzz0+7sB3xuGCeblL2u
nxpQ/RNRdpxIAGARo1WT9+jv4iZT+Af9oKu/6U7OfXqZNj5WDL6VFyd9P/22+inGBQVveg+TOpJ0
jKRa+g166zkhsUoxI6dYXYBEb/xTopETbHQh40si
`protect end_protected

