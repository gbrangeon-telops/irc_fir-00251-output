

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iaGK4Vux1Zzm9gBS3KKNmBXNdPq+lSqE3Nnx40zW9JpQDS5U0+JlSB5O0czPvIZs1e6N9M3JonU6
/VRFISTQHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hnTIGD4PF052NtQspkoD0qYNWsnDfk/EZli95x6g3PoDiWDo2i9hfthnklZPOTwcwwB/on/PGVLy
LOGgor+yT4ZX8UGtoSmScYDFDjshoGWHhtXrHczoGSF01e42zFHCzF3p+Kqif4EYEFLVI0b3qWfo
JoBwVA5mSGa7z6eKZ08=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jM4x3jcOa6ByCa1VWDPoU4L7JC2eupLAavYhTE4GTMYrnvE7xP73g8zjlwq1G8Zy1ODZ+0DDopVA
JY2gdvefh3SJisXvlbuH55643svFB8C9ZXe+EMovXErk8XGGsVfWZZ9248m2dlrUXREntbWGdORb
Fvho+MXYXuv0DV2DKImT+u2TQDacpvX5e8ltSYsMmjYxEdkZrVMF9C544bgDvuCE9PfD8XjA3SZW
m5oOMSMtDQabvtrFCxaEG4NyuxA648giN43WXdidnKPUkuB/HxDMEcw9NxHOVNuLeVs7mrwTNW8a
Y8nkGhyssdB7pA+UlWrXAfs2U9Wpi6SjK7D2dg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l1zDcM4+iGcttYyoR8HHgtSyP4Fiyy45WEsaODDzemrDXcJaURYpyLa2UgO2HmqSNgBK4XdlSO3S
QC2s2wdlVLq0nr6twxtavd0Mc90p3l2akMlkawzSfWC3lR7JsZexWZNEb6frZfXhesr8/8i8wphW
9oH5nUnhDJDdlXi2xk0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pHbCg0c3yWoABGhh+X5xmKdWu54K0QNaj8yiI7dbYcl0s74Nnt3O7DJj12bDcjZRfdRoiT43bXo4
30QPK3Jr7E41USUv0QfI981OyCHaIYD9DzkFx/42CQBEOSHNBrRTW/rge+4hugPE8z0ogrEZGdei
kB3oPw27BqROJcBQEhzDTOz6PP5L7SaiUGBsXkKo2TeQ1sLfd6VNm52eUhSewTFcPcdSylZU9gjA
/KlsPUnl2PskRWTiOzVvvy7q14ROz/8yTOqbBslSCNrDfBQA/bwCsE4HN784FAGU2BIu6GH0W9gV
ySlMw5kMiPDazI4NmLxMcJvTd4Vi8xnRt0T8Dg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5728)
`protect data_block
u+Mfz3LOMdGNqAzo5Fjqslv0FtsJvj04qFhU+TgTkxclkoFMzbtaJ86JrpbBMPhqV0qnilhEV7TL
2h0LHAn1YV2u/LoPn9SIEt3P0Jsr3n6okz5lPHMiFfta/k1GsBg4lC05gU8w+SzjrpZ1Rm69eu1H
+xfL2JUXmaUvD03WAf8GYuT97oUBD3+6+oL3LeSNboWKoEwII1IKqN6JiTROvEU1RP0LilpAZ9Zw
y04qyhakgN8D2mS3Qhgr02jM6thXmoal+OJpQxVGH1j7sihdtjsN3AP3oBpmWwQidjdu25JiOuYa
7vF0NGQj+u77PkeqQ8QJ1JPAix6C57+MQV5uEgBDHYqHb+FYky0KrZRKutou4hELqpHxI6SZwnSO
tC+Fd8EFFF/965uwkTtbckVq/mkEf59C3Y+01NgxtqsYC9tfJijFXngGZ9O2U71w9qwjwq7iQsZt
LWNQclxkC9L3VNetpT3CESBMBxZYzVsn7XTbOY56qcvR2RyzE+oXnU8WOkfMzitpDeCsVB5FZvc5
TeVjVN5v9g2ldma3wrFkDTaQ8RlxQyJU+pyPsdRFWyARtQJLU2hHdO3o+kKFaLfaJyJPTz7yeqMI
IrxT48RGmVh7IlEbtQiqjv5TpJOi2GOJ0Fo5Uqxn/+L8t9X3dun6lay09MaqOeOpe4yWUv/oQqtV
IvVU3w7GuuIIArKa1FLqhWJIZDHiEOsKzcxN8Zni6TPWqoG9vXdQv53hEN/kKv/IroDpsCu9AjQX
yWQ9YM6gZHsNfe4yVh4mmeyvdARWR8X8+oGoqwxiA3IeoyN+2ta9vSvLfGI5u3VkMzXqlncespQi
dKkD3yfcSjvrt2w2Gbjzm7onhdly8VoEotTGEw/wBxI5sSr53pWMttWNknV+zPNXp1O7ZrETsRWI
6TBmQ72tBYKGgCTeC3nlxMe0a1IxjJ3SO8rfhl3HwlIp8Caih3zfXC59Xc6jaQGgP4/uI13NXzyc
7eIi9eXAdO6rAGEREEQe/hN4KGnj2sWJC0pIMFeZ+hE5qiYoijQVUYajgVHBWXQnn7mkC8+uTjWv
eKEKioO2M4vNSRqb+crNFn9ToiBgP4abGo/ZUIMX20tiL6ETXhYQY2nSMC5zEaJiNVwiCGfYJFL7
Xea+8Bx74qOMi9dTdsvWJ+W/8wqvWYsgiVD5KCLSNjgWIlMtKOcVSE8uNoHA8pBYY+DW4pA8wovR
9qt7i+3qAmXm4tYfZyqy14/aqjnv5wu2KZlu7wbkoh+zqrmce1/7CE4Su6sV2v2d0ax1HNJymmgi
RwlHCsY0tK+go2qKp2qPJb5f/aXvYkJaYOx9bjztgU6cDrY87jHL+L1evg9abTnLFv+UHrnhSe2k
/Vdgg2gr1XgfgqAyNFxOwR+PsNjny9aegA0gRiBaZ9OjsQdvLd1pQg2nrCFq2leIOeB1YER+eixE
lKBEfhPijDX9Zq73AxH6/Xyzh/tVOheV+Z5Mp1NECTxbJsrVctTeHcXCPdLmKrgUfe336i6CinY9
kKJC9HucPrR68sIoGTF7kGXfq5O9QJxQbBpCdsjVt7iZTFfEXLBgOtnodQv5fr6dqjkCJzcXC1Q4
Cm1MtVzryMXCD4hsX/+Y70NK+9njyX4lR/oyX42paygY2hAvUoPqZHF6PEi2A56QS9xjOI7ejIIC
1odQccGIsAHNskRyP8pIDS8fxuTiWzk/G2Os2lYWJtn+Rpp3I9r8CXJ63Wt8jKD6rFtNJw/5cCw0
jqtyTVOeKn0qrhu8mU9+csjCi4NlZKCIYt6bIlKrm5p7/Y0TI5/JtfINGMNveG0pE+xbcv61HiZC
ZGxf6nAUaLvNcUBMQLoH5/Crdkcb9kk8gzYNCCqdNmd05dtg7F5AQCbWTztrlhGPvftjS/5f6YQA
vyloy+H2F0sONvCL1+dzlpaIQLxOCTI+aFkM5LCHIGCtu5khK3vLE54A4Wd62Sm8J2Jk1+B/179o
B7YXVijueuS4Qt6hpZZ72eHsOoFRmNbDyHRB6fWi4PBEO8sOcWEKaOZvKCWg3tsKt+HsHxr0gi/G
cQOdRJc1jMP6gRdt4erQcvg2xab6Kj6ZSKVIqmRYCDfD0eEqyx1dDE6BpI2HK586T8p6+ONijOyX
7HkPmkAQWyrVNQFT8whKd9y5fzcWdxx3kNNozmolAGmPHr9fijxz/wXuwh4mzarECiPq848EEqHo
0yNGUKxCci1cAEW2+CiZNM8LmzOYbBKOBar/XCWtMa3kNNcT+zGbKGRP/TjJofqfXf9VNbrTW46v
DrbygSOWWizfgeYxjhjoRAhhL8tdCGrkHF9So/fBzfDY4vSZZdTNQR6qWtdtd6vN1fazyR0jDZSu
2RHtemLn4j8nK5ggGmhEow6AKaLMLfp45iAoF11lk1BCQljcnZYd7BDqu9UgTYKZttTsygjLSs1q
wPZJw8Xdk3D0XScvOHkDZO1RzBNVel4z8B72eQS+K6v6QHXgERDhSEq6HIlZIWsG1QzRBJUt37+i
AUDQgVqrCsnAYpnrRp2iZdHFuUlRswKbSvLfUhohshUzY0kZnuHjagTRFaMjQGPlB4bbRLBCpFbt
RB7Urp3oRoQbsCvuM9gR/06zwrst33aeP2P5MOxjuHlYZdtarcoURMG349sb/EDAa5YgVprXnSsu
PO3Mxaf/i25mdZtUDcokYhLtZ0zH6sLmxBr89cL3jhJ9ZXUWIuJ+LC+xeytQYzrAR5hTO7Xp1ZLk
cv3enAN5YPwPQ9PvhglbTvRveLjSEA9x2ukd/F3FYAVIlFTj8fgLemiKOs/BfH123NSKneatqreG
pEnuk/+bjtgVF+/dD4MIAI7Mh6c03xHkG7vWMl2y3U4hZDNQruaueba+B4syoU2hiFIFFkzxBgJA
3Fp2V4b9/q/prWon+qRu8/NaXyvEGMfSm4bx3c+0zVSZK+ZA45yhz0GqBqXdj0jwNwwqNQSLZDsL
SBuwWy6MF4HhcBy5h7Z+Htfk00APWW1MvcD1wAFqTw3CFwccaxcI7nlxAVzAHNztzdkn0kh6kvio
a7rUrGGc4kLaItub3QtZg235sQPWJKbziJCHkzzzxnL1i1RMYu2Gdc0FyqFuIv2vmtFPF71TP/Jg
HIsj57xhNb6eoXYv6rMVH2xe1P6GatzFTcFQGXur1T9rhEeBatbMoh9Er939aWQGRXOZNe2Y10mv
NR1S03bAS/02Pjy29TRbo5NYFgvLhXTrDn2IFNgEsYzgqx9nJd+DooxiV0wHlfcZMZlpy33mAO2X
KPHvb+sc4caZHbJqWnDuLs5aOU1l3lkJ5StNX/KXJ0qvqBQrREmdkIKVG/5EaD6r2YUHlqzOemc3
94MIG9qyJ2xlPupWsD+rtbxo6PNRFSUp86+msxm1TUexwEwm1cUCDKchhATw1hi4Dl3TPME/mPZv
/v+Y9MFPgqjFTEwl3x5sziUys9+fz73I7mq6zxwGaU21VhTZawy3Q4i1quDOEeLMgspvmLINnE00
zFvHF9rOidi++uGrFAQSunEVNCqvUa8wZS7h2v4HV5SWMd6ZV6G8zDDmMUL3FBH3Mu4P0FVfoNzr
8lHHeEb/1V23J6hJlWHYWDarbDwqT1CVNMpvdCbVA/vhxecK6P42kbBLVltLL7E18+dfC6c1HpyR
zSvdgtd0/TMknJqkAiyDnJt9z7QxIXOzrDEu5KOwksjIhAZMyPNc56wiwp6stnJB+Nd9ekfHdTJg
R2MRSDTy2To5qaNLc3tbp1cIGoehvPeO/CMDxf0RpHeqm8tie3hEbVfFIh8c32cwx++rVKaaUJ1+
t0RbCjBs6jBRCCQVHVqbZUaNn76sUp3bs14IAXDzhIWQGubFfjRIM6Etxk7oh7I1kqxpNx2WhsI6
CcW4ZXQlKBk1ePUuZipoLnvZR/6UuJxfNWPo7GefEau3tyYjwTwrAEuV4LF0rzAF0TLrktpsoRzS
WkHE6PaqLyQptof6UWrGtpjs6AJGF+ZLngNgLMduQL2X0uUriqRyIjkBB5jWe04Ql2NbJFU9fr0Y
lpiAHHV0n2DaB+CKABTG8pCzyF38q8jgBXZeC1TE2MgOFq0LCS2Ey+MYKcxwzsBPf8+qhYZmaNVQ
DK8r6UM15HFyEMQ9EofcPUM4xfFGvr+TewzIAnCAkrSYK2b5E6l7lCjxeI6qb+RHsbQRfT3lHlIS
91SK4OhhplJyM1Kxpqt7ghxa6wEyChyRJ5mO2PlixPr4FQToEh/6TzqVDCjzXMInWnYY5Bmm1EjH
Lb1GV837zDVt5NWwpvOGP8zd9bbrJswfQw2auY0e3YPS5mepn6VL5QssjYs5OMYAKKXewyJv9hiX
lse22n86jzAtD70y4HoDCVsQFjpqTExLfREKePa/L2nDIPhdobXCY0RRhjQcvZWM851ny/sTsCBE
+rq5Sn4p7z7LRXdZqaSf+RX9m/hd94sGGMK+XO4IhPO6OqQ7E6yn1MKQh1jFSNOb+bxYoejMW+81
aAzaYJizgBWBpoim+uEousYy/Ts+9hPD7G02wKZzW8ZlY4xAWFksCsHQwAPF0RZagq161enojsxT
vxB2YGaPU6kRbpuNJq7wMifqrQUb1gNtzc02s6UmSWOxiJjfCbvjjWMKE3fYzfH6mZXW2M0jpYrF
mWt9r1/cKWPnN75N/TmSnJ6Oe+HrNAIvjL8CaYku42mcPpGIGbOmstiPcvaHB5t1bJsHW0jOA17J
g68CQ1rH3jg5LD19U4RpyxgZSWI3iIDJP8PaucGgJasJSm2S8si8XR3znSBvXG42JPIhhmWl8Q/X
amV89wYIz6ErjdkJSuyhiW3flzq7RiIro/NN3wgIb60w71wTXHUprTXjASi9ewQXj3PP1D+rUT9B
zt5cwN1Fn9hmUDptJm1M2sDNewxkJF6aZN+Wz6Dz5LcyAq8c5aSK2Oy9IebHD3fzFQ6UXkArC4dO
foNzJImOPXIzz2/V7pTNwb90L+0UHn6C8v0VtkP99fQ3SITupCQoM9Dn294VWaCfpIn7Ey/E68Pw
a4gRoAHCEHbEjdLhodd5eyFABdkDdpdtscIVosO1mgPwc5jOJ14UvOhnH7+MXhmLtP/kucuqEuFX
Nh2Ej2eSvFPuD8NXSCWSqoeRusLvxrSRUKoipAef0TvcEsoHcTGDaeqJVjGNZEvC6oSuZ1kmYRSy
BJodDjE+pEToLYFlNiry32fZp0qnV/yDrkr62A5XXsSPW0DSR3XWqRVxIHoc/HcMjrfYg+Beq0AS
yjotkFlQbnxE6Nzmo5U2wr7V3DM0ftXql2vpfnVjiKhxlM4zxFqv2dgrgVYNA6cun4GvDHIXLu0I
gvMPI88xCBpeD7BUV4kf7tWYKXd1cgUPecxmaEVdZuUtEc60SqSKJuWlBvn8SYXJrdTrzufnkSKh
r7M0lCBGSxISG4VaOGEDlcrpD1XVlNBBjFUjVyc9vxmFlKj48ldUf8pLpVT8Po7n7mOEZVN+B4Bn
PaN44vd1uEDI0Do8GyBHrooLzzDlt91I8e9thRMbdP+ZM2+JVoXJbV7a/GE3QSysgAxDRmLnr4To
MIHWL8N88yF5q6IE4u4npFJlZWqUCbASkbXzlU0Md8lJMv9Q7wi2qVBN0UNJ+g2sqHIxRdPl7RYU
ARVaLblDvKzdvvkCXGWY28cl8GCnkURX6+vz9RRlRSLDhqd8/N5EmR8upQphn2gmdRmfpd/kktLc
7B5Kvhk3GUwiD3d/G7imz8XBnUAZ7GWvfRneCWa4MJFMGeztgFop6TWiu2mRFmeLyeWGl/O0vgIW
pc07zn3F0jkdK2xCZ9CIGmDNS8y6rX2UTfmHqIN5rKzSpiXRgdd+mIcyRrCQwN9ZfMkrteTBEG0l
sxkP0L8pW42Nj1PapZQuyhGwhq6aa0XmM7CTDojoknh/mlAMJe+LCqr/4RkqntR2z0wlVpoOy3NY
p/Xf3x029fYjgLQc3MKgGV8/qjrYEb0N84GsByjoq02bNj/knw4cS7jJMdAKkK8hNREtbFXPfPb6
xxagNeYTLpu+Qq+xvKrkEA3GFB6/WA22uui7E1v+I+lvzFkomqSyewJhYZKrjOUxsrBvoB/Q0b/W
8pmLYAeLrcDwNi/4eJl4Px9vrL7EBKccAFiqeW9qwe3PgrBITLJLj1XJUw+F83plTaSl3OBYL3sP
5J6M7sidx8ungYIPJe7ngvwi1yKTpeSGEq9g18Y9aJKz0eJTi9BTPkchK3e6D22YJIgTeszgMXIc
yRPKuVK4qK/Y00EesjWmrxVYGsrjAIuriReMhFlEibl+ruikIJCu7Z82gUgdw+4TApU1PzhRpZ7+
u9AXaTsCSlxO4SSg7IXrio2iK52+tbBx6I+X+aYXCwKxlA7L3/9JsDMHHQnkgAXhzyKplu0i3L7Z
7hqNewuqOTd/vVMzTBJpbVpAJWYz5MSW0BKYew78/5KzNOHsXz61x768uWFj+bgk1wcssH3bzlSC
lsRky5oRaVb4RwxqTuXn9/VyS4SQ9/Cbmp6e2zRnEJTKFHPiDLmRQiZV4sI6mHysoVAr257O+b8g
P9NlM1jOzHcUorvM2PCWB+FQPyuOnR9AcIdPAC4f1qvIZs5DrjYj8qZxcUjoolIUX0B95giCYmAj
cnNMx4S/g/1FtjorkqCev73qmDtWtlWFkqBRQccl9FBVdbhMl97+X302G5cDBXyb8jonhbzcv83s
ulWQRoXtQtT3n4d3CF7rJQErMs2/5q2Dg4RALxY/RfGT1mfssONQ/9bvJk9hzWBExiFgNrkc9nAn
PuVYjK0nX4tbCNEZMqjwomaX2Oe1ilvUBvLY/eXKpeShTJDUmviNtgfVW8zK7AqmrI/O0BR2VluD
4Ou5uyTeYU1LmE9wtWKEn85mcyVsO8Lh0uJj2rodbbDSv5TIAY2/yHcESVtgB9SPCPM2W4GSljE7
i3MfQb9F054oxPrjsJ4VCTpHYxGEvgYwfGN5Y6EwcxajZ9OmXcnIUVDa7nJUEmCq70VtP9SvlSvx
lwzL7zhfMBVIbjDc+4QkZGtyELnlM76ekZankZXEaj/82RO00YdON0pmNHFDXx6bJSYDK9veVoId
jam8ZhwB0gGUFnO6xiuiy4sQlPOGGBBe9fJefJAtBQj0+IfBM4GcWnrs9USXH1JAXWHCjHhUmvdl
PA3mZsDZBuGY+6IZFc5nuTEvDvmmfJ7EJcNM9ygF3d2D1ZPPWLk3FQh5xNb3H1r2hTFppD5lRdt0
B/9gSxiULiIIq4HiRYAcM1M9waoHZsEnfhR7lRThjmuM8WL3vNpvB2emeNbKU6ABqtdbImcxVawk
woNtokGRS0ImsEI8cJjEV4wdVnfiKftZIP0x9Uk9jOjCnfXUUm19pr0OlaMjR6MnnkEsHoJpubHj
a372YxdZcemwIlC7g6/ir7xgApECNq64FF6titsNSakRe9hxRUQ+HD2ImznVOGsmY3sek6narI0+
Kf9C4WscYShrgXhwiHq32jPm6NXgwpE0OLgBoSPZBYh5YohVyshlVwuX5YIhSkIqQ8Z7yLs44HiK
io0M5xSZz/gYk5eNmh4GkZzCcVmIE2Zay4O2hKHL0bGdu134d1KiYcoi5BPrfD15IzzhsRH4cSuA
utUBhCu0Hzw0xouStmKJ/HxiV3s16RGIgebkkQ==
`protect end_protected

