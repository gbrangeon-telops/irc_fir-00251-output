

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ahdDAHzz440n+Z6SrLNKLMBChQ5FzHxmtmolGyaGzRzZ6AsdM11MYnHQlmkXolfzuQvsH0tiYFpA
bdhL84ynJQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qd5Te5HYUFbAOVCK7Nrwmf+xhp7iHLV1qESGeKRRemMuPlhm9gxKzGI5glBpEm+Bt6GS7xBHPesU
Rh2RxY+9Nst/QoTZG24XGDjT8gulIAFW/37G7vhPLNVOq1gP33zQ0iNDRVgAsbEBqL2aP8fzO3c4
Dl1oSNusYXsdFmxhv/4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0n9Q8CLs0GcRArqoXB7pbLNq/7iI54QAnaQ3YfVTrcoLuaPhMipi/u1YxvxCeQhStE/q36RmAWKU
vuVvb8WRD5dX8Gc/5jIRt4ORXRhrtme6cizBVjYhymzdNTAgbAuH8k+0No3YXlnw3iXuB/bUUXlS
9ThgyMn0i7erFTJ6h/eogbI8EG6TwEBPQ11D5xXxMjzz9Q1WQ4L1w3R2CAYnCrSSlQxqvapc2X6+
HzE5EzvdMpbru1PQrGeGwaFtvlT4dq9BRwJcYQeIth/77QtTOb09uuY2bIUtRjnczrx+97he8zc4
F2HQqnZwdLvPbSwwqlsUdlME2ell5wSO2A8Cdw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fXi1UCgHICyjHcoUzs2uXfr4QL3Zd6fFq0YYnh7DHj/Uz2hpTBP/xGkihvbT84E9/Kgj7lZnbxyU
NW3Mn3WgobnvsYj6dHFEG2LfnPYpGw5nhTQMawWoftBXy0o+AjB6W5RQ99l/hgORyzZ3gEP6q1mQ
SG+9quGTTiRQQEHy3Sg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GxP7neU6pelOGsRYeMpWhq9H64emJJW3ch5ZqO94Ja0S7m2rL3jKbNa/UebfsafxW/Jq07+9ZHQH
nakVk5fs+waKW7fPdCvasFZq3bHVoH2M3uf0FMGIXnsyGlgHQ4qCnawBWxPqrfn3SKY260XmNThN
PHkcyDSRI2OjZKzXzE7AHiKXBnUYqYuy5pZkIRpG5KuuXSL3l68wM2qwWAk4Dy7OFak+VRDwWWle
Ve26y55BBWyX0cVH+A1y9sHRRFBM6x678gQjaKYO8u10cSkLQEatg4BKcHaSLpXozsPkT0ktveBN
etZKKhExPa6BnJyzgqh9xypSTFtCXtbhEF1Eag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22208)
`protect data_block
rbjXPs3nw1oRR77nGKh/BJlKqIeX5zEeG7xV40SXwJgdjvlWukLI9ekqIDIgO0S4hCyxOLt1Jpcq
bOsvug077f3Kx1PQfzGtqtBAPYPOctcx0XmGBK2fmg0ZdSiIoEcSSepF2RpIklBoQBxqex+zGy1a
9u+j3EQuQn40bipfLs4K3zh0iufee5zlGPhrr6zjFmScWNcN4wDu8jBSbiV/OrrbeaEQjgWCkyG8
gjyZx5I5xHGhwB2uChWSyrMlBb6tFly+Rf2nRBsr/ECLai0EQk/UiN2ReUh31koPBzjSZwM3s6T4
tndb+ZhbHsQ24cboyIfmxScxOYA3l++//O3a8cBw4D/vuqqpApg4HweD16coNOkT6QUvmOG0AiQ6
713ctE4wChNtrTgD9beF3Cgc9RbMFPncvEACLtypU5QDEjdSXdmkmVvupokEoBBXluWbDsrVv0Vr
VPAZg76RET0j4ba3uPujQZ/gMMdBFAvqsLwAK5P2na0E3BbnKgx2atO5OoqDB9QX4onxwAyYR7Bu
gzsNmGtcQ/Te7NkINUI8aGJM7VNIG9ETQEaPrXGqtsFDcgzZWL3fi42XaDe9ehL1Llwvk8lYrR3b
MIMoYI7CC1QatWkCmD/9B4d4EGDns4Wrt2scOeM6D8s5z3kmCv6vObgV440nyCIWWVkIgVK8TIyR
1BJPmQeqv/3ggcexdmFULBA0/nN0oQQXZe1VTiYHzpNONNKxmn3q3swtRf4MUfheJ6F/z+U+QK58
lqI9I6BLrhKMTAo6n/hlDU4u6xpF+DU/zkq6S1uNb37zKVP1kTOpajJJfvApD9GWs85dGdHMPAb5
uBQtdPaWB/SD5YQM6UzUv8KtpVpR9mYJtTGb4O71RYpYQdZofsJe266nf0hb1BbVgPiAeoiHZz0j
pYRi6WibZU5yKmbmHz+pk1b0C7exjLQqBJb1oAL2OYqWHdYmCMm9KniPN3/zkwzxgaU+5dFklHCc
/isLvAER4ogHmHckOhucrGaeZ4wk2mDY4vnJQZmpJqybtUS3Tbua1nH0KyqBhE66NyxEvh+9X2B/
uEFmtlgnhyCQKnz2uJ/ueoVWUWjIlrk3herWmC4g3kAVOdfr23B/cqYg8rdsdCmSa5BWKqsDaSbo
kWXdUutWsgOjrSJlfF8KGljTOYWtbcRkBloZuQ4phOPMJvM8+YTdfAZfo2tkvQnAowr39jTaMUQo
M7zZDfUhc65UezSM1wlf8rwmlvgfBRx48wmpKNhW16yrmZxO+UNMRBnT04Vk+/hw33Zhq1mR/6JQ
LiCwt/a8XGHVbccsSOS5sT7TdkMpfx6M+5ZTRg5zKMmMQxNq2Cb7NLobzhea1pxs0mNkiPyB3ExS
sb52X5FQ4RqcR/KsFACb1uWEnwCrXxr87g3GQwBgeM9IAQCGsERe8mJopsPwEJq6FUeLOHEfQxbT
caRZfklKcITDjfg4aQhWLjNpnuxdZtZqtm7gphxpywsiW8R14FCGY/GjHeJGh6qmILo0yFsAjunz
XvA7nC5SNpMdHhPdbp/TrUrOIDjSAbYiNfitPxR8ZYv2wx+3aOf9lfdylAADCTJWpWZaF+Hzw53Z
IOrJfY6SODv0mKp8pEFLddGF1ZqFPCzGMJ3QDdA/mIU3EbOw9+Y+UEyVjUwL4tBu1W3Valw7OyT8
GntoiCUv/Dw5KJ6ljUsjeZuvBr+XPLcIx6ER+3DZTDpdkE0Lx5rJ0EqClp6286gHled88bT0paRL
oziFTaBvPZ7StIkxieXwaA/HwFpdfKipdxQO8NGRJN5eaKAUEr8Nz9KlG9lhe9Sk7LXNLAqE8FiT
N+2obfaKtiQhF6FVyJuOkn6S3kVlWmNyQiXe69HpqFcpIctniMTClnnFfenXA4ZZGdUAPmxCxb6E
T/0uDYuvRSV9XBiSeLz6kbMRvIaJ7eqQ8PCMGeBCiIlVwfq5qMYckB4lSxZQuDxFMjwf732nKmq3
46OTIDLgCK/BvZ68aw/Ygk66b6tELQzWZXtBtIGXrmxwXCJ4Yz028NiZK8x6b1FjcaI2DhHMUb6P
w6m1ryNs1GWBGkhAuZWKUtaGBciYV5hyQD2nc3O56nwZhrZaMUGKqy0RKDsKLIu2/ErBWdIaPna0
JCIuUEGpSWbqK6ACLPh0hBUk0JQ8kcfDlDNDJM5P3sdooeFBcuhyQTARYLAQ8q0fEVBZv6C0/RIr
mMWVbwooACpaK9l+TbOXtEvJObpl7+1CpjTM55bTW/YVnsrdFXsLdaUVdb4HFRmiJzRFb3QNZj5s
Z/vrLTPapOkbk2YzDsCnC2SUEtwQvxo3yB8N+mVPjcg/uZk4VfK85HhohMRrdhSE1Jd6+hXqdVql
3qtQJsml/opd5TKLRb4jsuZA2cC7OLZt3PVGRTldOjsNTSsLnAFj1Z4l7vg/D3s3DVjMZQcapGcU
AKLwTSnb/ZC1grPRqrV72+xlfa6yoE1C0SsFRQwKpAlRlL0F67Kxjo+4WG3FpSxJgwmiOPmZVmp8
h8DkAmXnvkRyvYugANvIo1WnRXP5hD/huK9i0joNGF/Hc72mWNxezbxTa/je03kmVMrd/fHpr1Jd
FFGUidXzYkw6fapU6vlKnmW1hzBx32qSx4OTXuisr8MebMHNmwkRTlyLBChfr1TlDDsWxsnWKDvj
4UOxzu505q60tPNzPA6pKh5PA2GmtlMOQjQ+/84kVRulXKua3yp0T/2pOOOItfmcdKWWhNS9aRPL
0m/vyf+hAeXVaisoFT7tFh+bkzbMaZBcEjzFE1aw0j/+MCC88RRTWAkNdxY/m4Jcv/ifE74MWTes
V5XSzqwi3sEEhChjeItFmKXBvz9dYb5hg6B/vfXiMCMlmu6bJwB+UBWH7lOb/C3rgNcPfIsNjf41
+aLpMjPqUAUX9h3aKE8ukTDF2y/RGXQyuT2DsTuLBytJmxsR+nhOtlTPYG2FX0f2B7/XFL7Omh0q
PX8V4JUFRtVFw3ffQWIR4FnhYqF2PW5GQMILTqDRjTVGF0IxL4gh33PdNaOeUrw3sguWZoiqMHQm
9epkadVnggDeP1UxsHeAGHoluBDdRtrUp6uRKf8pOs7Q3D1MpQUxUMh/iJSrosRHwudiVcz6FB7p
Vi8B0zNExEdeQM/CO0Dr9wD+Tx2Adr+Ni0R9YFPQHmbOYDfzJvp2EpCV2g+K0dadT2VGLKUn2Jgj
7deWsZJNstsKlVy5+Vd5NXAn//h+a9nTstQ/5+TG5umwt6QQ6IZ8W3HOkcFL4qNNEb51/Am604qu
EkUuakITrgwzzLVUwESEQchg/SUoa+DytLYOSXfoqU23OQhr3iGQiNkQIMKFaWSnpg5kT7AtKYrL
IMPmyrb2PLqChs9UP5AjP0Dumhk84ND+Sxadn1xEELpK/eDWWwB7BVpuuz1gKZx3oEUiZTt+hVW+
BG6T0Bdl3SEI/1mdwAGS5gqhPjV+anCkcEyFcpShkEOUcXqZeYODyGYXggAuu2WAvcYsrAfLg3bs
LYwby+LSjMWJ8n9Gh+JLrrsFLPsBHvv9uG9JtOe7p1uE+xyz732rHY2+8fV60w8DPSMgyfLglDtm
AcrW1B/qZKr9VLaHJBMD4e1DYYK13xcF4uMvsMQElFlZ/gBsAkvs6uFqMTD5DL29KpkPFDCoMH6G
OwDjgdOZOz9zTK6Vi3kr1qnv6E1GxdZSP7elWg5oTokuqxIyQzLahcIKdNI905yu1XgAQnQK6Eeo
PAvwCEhvecQS23Wy3RpLHtsBmOB6Ko54k2HH7qrX6VES3TDCj3uBRNvNoU6fhYM01BumUPTyGcdk
IYNfT5ah7/uws9qb7gWG/vAGezG22PWrkUbXOICjW9yiIKcuKtq8334iSH5mluUFB4QgyM3h8lJm
EFICWYV+LZ5BxrEvv+8voEQ2Ie4I/mP8jKExON7Ef23Zb76CBFFTy7dk9VrjEiclAZSzF8ZK/2EJ
6EY053kIzze8fZ7MGq6S2Lma6auCZa+0TUo3biE571AO6Nxv85c+8s4Y0QAMSrfNbooY6Y3jJQg1
RPavJSjEPCwuMDEWKY2aI8KfVppuecRF+LwN5YMzArtQtb8Pxa+cnxvkdYtQ0VED6l0bQ+QMcNkr
D+K4Ss5YwVR49jKa/KYdfBYZxXK4DGHkcmTVXvXyjseSWIYSaYUpaOdDhplI50nhwTXpS3MyHhbh
vd9FZu/G1NbukJuXzohVQbXNi2qKrewNgsks5OUkFZe4cl2BNdwKj4G9rmpqf48tZvun3hTeAD09
S77CDTNXSPdnXw42VVPQoGFJpKgGy6CSnBTxP6OGA2bxbp0yONxn7HW8QO8E9J0PEdkqbL7/M6FK
1ND9MAhCJOxaX8zX+MaVsZF93sa4yhzq0CJi8jbURNJTjhW9ZU2zwpTgUf9rQS4OmY7Hmc0qAwMx
DThsyJbSOviwkWy8u/uQ1npULlm3tfaugSZB8MNeG1yEm5Vjj2OowA6N3BP3TL8BljXDs9KoHM/1
RHopdSSI8dEiIpW2vf0rIGLHmURqum4dA4tGc1r0aU88RV/aDF45CGBPQI7p/e20q/w7Dejw3E21
E8TLlwUkCVKhpEHOniazwXBqstVL55V5yNW5QyKdFLa2o6AAcoxSEIDw2m8Yd9B5QpZkI+fcoHbC
spPsWZxvMKm7mdATnuPVztu4kK6/ddpIS8eQri5UkdbMaSSkl0jfA+VSamUCfJrmyYdCiDRugmJG
2JXLwKXO0tK2kpxBqeviomk+rZaVWJ5VFJ1cXRPISjp1MQ2dU6IAg/CyJoW+OBeG9lf25v1NhVbW
xPraRrxaIub6FvlyTvm+U5D0/deAJU1r5mbsKw41CWkorX/FTADO0YF8+6ygVRy4chpr6dVL2+lk
Z7qq/JiHK4aEo/Mo+oqTbIA+xezzPzchaxvj92s0+xlR23BvOdHMQu86Qcy3cyM8VETkp4lBWdAa
VoGRoNrnVPMHjVT20e/Gi/5g0tmagvImXS1zBSwav/+vcPIcnmm4IR/o/CIENzjf2cRG2eyaNyIH
E1TjG5nVRGdIfS7APHL7dwouvxfdmwoQSFVzJ/noOXJknwUUc1KUwZMmr2UneRf/OGtXahWEtbom
cnvJQghwM9bbEuTnSPzD6bUWIYjsZ2h7qCVixTm6a1bzdVqlNLcvC6dtPPxgtbo4FjtX4pvNvmJH
GukMH3aGWBDT2F6Go4BndG+crvL0a/XjlEXppNTZULX5wV4V7tDh/3EeIwIuJAEQ8lfD+AdP5nI+
ibFK68f+E9e8vDCMXw7So8EsbtcLcZ7krmLBhylp7keEOIx/2q+KbuoxfO66XHYRlEqUaMjhla0B
0h4Bf8CM3MSoz65/ELImnMjA26WW2/oqVE8WC6BWwmga8M99vAL9i6aYbYTh9rhBdRy0ERqTbC2h
tHLRzdnuQxs/8DO/05n/5qPGJJOmkBVsZr6AH395AHySZgmalfKzuQyA3DvMKhafJJrJQb7VVxw0
gq4J6XTJ5YBn38FBwL/q4W4gPtehcSYIeI5N0dwiELrUFAmcdu2oHkpQdPzc9aVez3AmiGsV1JHT
8lK7uibwDotgGW1EvHOw/rP2Yu4AYHt2G6UX44zh9pnYsBc2LK5uxyZQNyAesBUFSjBap1Rnf7Jk
rF1ZHJ+daB4XA2w/qKYe4Fmhlql98RVObcDbRWYCs4zZLo28IOmLoqBsOtQTBPjK3IBz2mQDDbYS
wuL21B4oFrci5MRXmqFtuf9ktrgvRc26KT+yD0X7Ts6io0kexBoOdixF+cXUt01ayQDmtD3KZZR2
PbpyPDgwSz2l47JmtenNVc++94aWyY3sXdDMETcFg6Ua2cQMpBU0I3OUbE10Di4SF1VMofv4b/cf
o3RI3Xd27my0iJF75VEx97dznPJo32Qolt18AukuTK/kL5RsfnqyARPWkFd8bXEEkj8hSOwPf/Wi
GjZX+ZCsV4o9f5OOH/qmrpNUCtgN+AUMMyDAM6qsrd57U7tw32L7KNqmbVoCy8CXSxhJzpEC95mJ
1n9WGSsyQeImpN7CYF5B9UcDfSZmQau8IcGCqHerY11dfDPPXHr6qth3FunXW0AXEKEYvyb74Bw+
mio4o68UHmFTFp3HzecL9cImwjgiwa/RAJnzhM2f75bL/FsA24nQ+ldmk9hvR/E/Cxz45lUn7b3a
6PglW0RoBdCNzQqSE6cZ5LMGt8wtEFbfi8Cquf25ZacvoMS0kF1QZABHmGDSrqUeOo9/iAaYzfQd
K2Bt3TFQwJXDyGcK05JpuXW9BCcoePX1RdUidP8/hzU6JTMSygwfmFJe938Q47sqKVQmlYAiTZZU
nHoPOn+JPFehtKbSZ7U7INOfu/sRuc0f1bxmLUBsBapAVnH9jE1F4qhP2xifoHVfQtlmtn5hmLr5
KLCVkDbqUBOEG9rWYvCIYcZN1fso+WAm+eTjZTOTIugokvPBzzt7j74gKlQp3iIksUHw3Bd/T73e
wuGvbgPX8jQjK+AzsDHtvwBeAXFFfju3ijly95UOmQ4pTTDnhI4unSMpKuT02/qxp7TB95EfPiWl
Qm5c5lVtWVZaFdrTkrkXMHiZ94HO7qgkAdzmE2VQNKQk7dEgRx3r7KUafu7+bA6DFrdAXm1z6UKi
nrGvfbgU0eCGz0AKu70gvtCdq2DjCvC+yrYe6hN/CQmf9u+GUjSz9QGozgS6gTHsqKx16y1G81ZI
Lgbun1PZtbWOZq7F3YjHdZ/s1GxruNl3ox4lr3wyxxk5efLg/DTdr+j1dC5cQpTkIQYpzzPnXbYt
iNC0kDDSQLSWwedkU2IZzVwKJv/W3kE4UBTZhxw+Pva06ljuGCIw42OBXBErqCOCC6WrG8SWBudt
ycqnu6d7t9R2tOpKQTv9GoTPNrNiqlZwu5OBYMNww2JI+ks2DdAEcKUGwHKn/gHGvwyvbYjYtnzq
9LOaPQSp/VRx6B4t3Psjbpg8bS9zqRMFCsGbUL5OQku+f+LIEkNQtBXLJXNMubb34ngxpSuQE5/J
gMXsHBzG49loS1gvWPJtWGBs0e/XBiUytog4agy7ytD1zazsRDI0QOPJPRTG9DExXPHDblstfkbW
mUxoLmzp6dRkiN33zErpe7demHpAqHm/PyY1pktG5FBDXPMhlyuzEofdeqqVhTKjKW6YCHOdoBPl
e5PccdKgmcKAwmcauztwJVWd2HWok3NQ7hFbcbHdwj6rXZsJcprfZHL7dSQO7l1snNmAnYPVJlh+
g5bTlenySfIJ5iRC5avcZRhudCtsdvqsvSwVjips5YoCGSe4zKtX5TZjGaZPOgs4TI12tWoqQzHw
CtOwDNTr8FsaH2qGrMYaYAzbvce1RbS0bQBpGJwcGxxMWyGerAnKCiJxyDQ0EAY0/G4351FOMxiN
JOU9gw3B845uQyUzyV6teAMPqRpN0sSwdQlaU3rSwsyn/gcmMnXAl0JTmup9y30nbBTDG9Pjw81q
LJJe5gBNYyf5qdHyaJ3/yjbBfxHZELNtZltPrP2fCejPHLU1/11g2wCGMX5rP9zMk2bGXiuMpQVK
56H/KA6MQoCNlP6FJojS2hv9QBAwPQrgME3vquS8WHdT8G2bOQv/F6mJmwD4ZdO+GbCSfDiT5j5g
/VHZX8GoDQZg6+SZzDu3jljqt3lPzOja9aEieDUIA3eMXq6qe5BWYWZXP17XHXXCwMWrMcZKPyDF
m1BKaJ9TgxYmhC9OxYr6ONQJaZTck6rDArq5YBLU8TXRQ8lk7d9fP4VnOFvGxuxaFItp6GMrmhQu
n0ATn0gtytTwS/+eMh3n9r1Z4bgtK57yhy5TRF4CZgrrQaXWHEwVEtzc3H54etNZaDsdKq/a4OTY
+mv7oAe6+OSYPZXrE838x0ZHQCJ9g2oa7/QkEY+4YbpBU00JB+UzLf/76D3Je0ncV1hgEqWynl5u
1EYiqbipygsij3hZFQ0PvDtR1OtGFE0NUOayQpUY0CLy10dwoMp0z/6GH5yDrwJ8T4nqBW4fK2e5
AWxh8w7nrI6ndwwTXNzgHki1eXyNc26efcD2PQBFYSZaOMlojRwGAHZqOUGYEM/qq/9PaeX0c4d3
9Qo/pdHPoZcOaDR65v0oqSK/j8b38l+9FPUVDQEemgfslxD50Z1R4Gz/FNmpt37by27y7gEqhte0
RKFWNJOSWTt1rjPlXO1BslZSBaTBy00f2FUomARGc9cT9faajVLlOfVsavl6uMTAmyITDz1Da8HQ
x/pNsE/sNvQYQ8NhtxwditgTf4rUyz1ZcyBITJMMZnAVuPXvI9Mdn3siZC2DkPZV1woPFST4yrtb
0ZMredIFhCrpQXjXcOcdvO4IvygO1M2R/Y175xKyuHgpRzBAMpCF7nD4RaazxSn4ELWMK/3vW4Qd
UwTN69VBeDvTAmtmtxhSAk2l6x9sydiuI7uwG5BHqb1xhR2ODJ9hxNvm/qkOX/yc6l84VKIzumEB
nM9pmg7yvYJs5UsyK2Sr5eBIwC0STTS/Bgjp83hblFmDbCcMfr8SxMeC2fDzIi/CaHU2g6BggF1/
RHNpAdCaFIxm32BH0RL0W1ritqzr/C/muvv+Sdwfyyeze5RNhgdj1uyF3O9ewOwtbfDV+jTE0q/Y
sU5WfJu5+sWyegJSP1J1cMNdiC9vSYdOS8Uo0Gd8IhR7rCNPoFd0FEbgBAV0trSt4h55yCU/sYUY
L7AJZGxursl1r6MoLZayg7t2qnsVC58rZx3+j+/Vfdk6laillK0AG/h70u6Zo0FGSMDkErbNlaUZ
YKEqe/LyknX5diPGcdKHHYfQsis1wqG+GZUzLcTVdhVWCLR+N37NuS/CJI8JOM3CfAr9Cq3hbzYn
wUDHh007EFrfiC7ZCZ76FsDhxd2QYDJmWpI2nuEmVrgUx0AF/oWYFJs+LU53MOdBannXvbXUwU52
6i4W0w4G3JL03+gOhHtWKMRoVFdRrzvb0dSX2chQefm+C8Z3BAEhU4EW8rk6iM1qpvCvO7aS4rRy
zceAfLsQ2qRLLGfmzv4qjGuGKRF1YkQ1KNWxFf4Uqfs6qlT9jvuvEa3SEgumxWfpbndsz/KUpM83
35gBipylQpchkVQ+w7gzasVr/LdlGOnuzfqN2iwG3IVpFF8bXAkol5jAfacBpi/hSf+OhkZLKuaU
NvnVEmTZVNv7qmF+wf9LJ00+MnEy19G5xFei0rnpRq4J5oLPCRIwCknvSLyAMNWPWz2tnEDpXCIM
Plu3qicuRc1qcW2SyUSovYEeTQOyC6uarYJCWiD0hJKnERtFyVbfqKbexnPsfVVALy+VdxpUhf/9
QGqsJvsTucCenWB3ctLlbO603iMYHBp253pEj22yFnLvx2z5J5/lL7iQmL1qXzqrCDVYM9/Q1bUR
l1QeqL20UlYuEVLHJgxs63I+/D1Ju0U/wn6Q/9hlD9tNHQ+gvNPJ3wDrR7iYVNY+iXMog2PSabRV
pGRHwLkKBpQlvxINk9kj89xWoiDd8PDDPYt01NA2YEPR/Ruj1s/iQPr30RFv/RYLo0ZxxdqmhNUz
ynlSohonlTHEywvXdtLzqybHFapzUrlyWYt1s/p9dIBAM+n/5LQUYgt2jkPYoB1rkg7cMAhLji/A
y+FLZrW4vkppBk5Bj/h2unLxVfQU08VMqFnCdFAD3dATBqGrnw9coibbBEMEDejPnqosgiWU0sjy
eSEMnWOZUm7oTHbQ006QK78ZjL+L+Fp53m6kMQ+5er2An7cgVYUjMDlRspE4G64dbCvN3itZ9kit
x4jvSL+/w0qJaTNlj2EMUKtPj6/Ewb2dS5PZ6D2a1MTOrtXoHetGbUUwAlcy2EZtpOsIJJvdIKAf
GyeGbwitvgVyKd6YOmk6B2HoFPB9GRdupV59R63XYRCrSPNGfg4RO6XK0JwIV99HQ44GHk97ILYm
ymtuqAsLbtnQjQmbme33y9rqlsHOAFxBYXfl4sHYEJURHibwau35nLFhq0b4fSdntiB8QRaINhBr
GWOOwvjdi2XDiFfAd9w1tndhDZKIjp3d/fqMNIhdJR+83XzLTg81fvidzCOYhXJQv2BqPvfqgY2b
8jBr17lJUzeUZ6Dl+pw96FNgofnCA4aYBjLwfu2ETptVW/yam00cOgWFueMK0DWXDIp7259nQ7+M
9Jut9o4XF6wxljsRGPdHPfc9cR3cmOyhF3zDjPPRQQ41AEhQf64prnC1eS6eyOVyGHY958GYvwpb
tk279VVWCghKvf5nusJqsyHP1hF1UktnDtOGVvtKPmUFJ+OBatnY2Ak4/DR02nvndUhyV4tqJLUK
NMmvT09/WlnJby6gxzxvQqVwOzdjc6T9vmJ/9YH5lV68zK3o7t1mLXCkVuH9Ai87kmim2n5a0Pix
Czwa4E3Ne+ZX8l+PvhyhSGl5DronuDamWtp88RDOmLHF12PLyFSUHn+YkFfJ77yE+y8KMDakIp2U
yeqCej0hBmdtDps+n37TizWVP4LN+BBRywahzeosFWlS6KdpyMzcL4n0jaKWqf3eyIP1GYEAJi4/
uZJgPRyciAr9+ZLcoDiJAEVuNaec53GVwmzRiOqyJaJK9XjoFNHQq8GK4TPvxVBeaB92fk86dmXY
qgQ4oBBx6RSdYcN1nXmuLymNVfX4DCDKTJ9TRhgnKnp1QT9GMZ0I9zUErJZzgFwWtanXMTj9XI4J
bGGtSxhU+TWUBqOz2O9OpYulzKyVV9cbD/y95BPD5jpyD/o0sE8euuqwJCkwNQlJIm28KPU2Og6Y
nYWyh3Dl0qzcb3Geaoh4MsDTa5TLpYhYHxx+US1D066NlYW86UpXRePIBjes/o9lHTt2mkDF+oYO
tAohdxlf0zy0CwoZDWHFIt35kzwKb+OoVnkkNY1WF5Iy3dp7zfg5ZKil92iFCl5LfLv0Hs+hFvmi
9tvNGZMbhYudjDHu2GogDX3ZWmfJIhl0V1ROR5prn4I8GPKGvN/TD4h7a6RuHlYP6gkmAiBDa7Yu
7MXIwzo14QY5AmptRS8sHj0lD/hSl8VJzqk29ArMkvGSMdANdvbLUIz034qZ17iDZsnlrIpRA9Sy
HUfD1QnovIfYrlJB/CQ2UaV3k427WiOM1wdPBaQtXU3BZiYuC4EMuO0fcdoDKgJO6TzDqRaWDPtP
tR028mJG7FW4Qr6dXL6OJkMnQH/NbLNz2aDWzqQG40OL4i273rsnzCBucWYEpUJpyA6/O6SJ9ERU
3p5EHBP79o7lkfDX1iVMXBZHCXXD38AN4X+yqZTD0qpkThEkJyk3tYgrYQaK3J+9wzl5x45uKpwX
m/e3boFrDxjnhsqPBS2R6ZsIqwAfcjPTSDfKlrt4NkCauqj1NQPUjQAduEA+7Zwa29+KHmffbN43
GsLVVvGogZXYmNpLjkAcUr83TYkDn8sxlWBLfdkx5nEV51WOiXQtSeZnSroZY9QVic9PqkD1MNYL
mEMpRj5tvhwr3RtDXCW2NlmIcy+7QIXnlXllHZtdQ6puNEB0ALBSQ7YjvfUC5mJFHLP3rvJ9t+PZ
COP2WdeukQwtT3JTgI9EcZwg6HsLgYJS9Gct7wVYksKnwloS/gdHiMqHRWelZibHsIIhnbDjbsyn
EJrSpizT+E3GuzTrpkMSUCAq4lfs8Ehk7FrW7fwA+gl7od+IyMCYRFPqgiSxzFbgOj1SVTy+5631
155cdtNTvDpFNilfIBgG0kkn3gczOA5qieaVFOFL8BG3AWXkCJzKtotmH6qO3aLhChpmvuCTPdqi
m8hpaiYn7LCLfPgo/B6m6TeiIWkrRVZfOeFBu5N6Oxejl3r6O4BKgdOlJdQxvx1h+/AVw6AYtj4P
TEOoNS9XhopqNN1FH2jAIa+Vl5U7e2uErNI126ls/qNMW9tVBhMB/Errb+hO+BqNVOdF3JC5Kwxa
/4Qds3R4WETTj4357g90ZTEEZ9OiSrwnB30jn8kRqK2M64hJgGVLwR9JEPzqSURobaAwBBHU+nzn
RXlbiSfLgAwpW+7q8DCRNpoBzgV9tmBrekLZMqXT/t+Ecxfty5yCJugPPrZgbrr851vR8+wrzIS2
3xXsmuhAf7y6g8TQhkUyTkncncPuxMpc2ZxqAy9P2uBPzWC3csf8s4l5P6Zpi517Rf8CCZI4fUI/
N12T3/SqaZQbrgOliPft771oJLJPItnGmc8DJiyUk0tT7RECxLZxdoJ0fsOCz4vUVsvdj9mwkuuY
wduyst5mfYeeB8dycTZH6uHDTvKf+zklZWxWJqFMiGCMIC++fClCwgBfvXAUoMczjJDI21uVe4vb
1WYLVLwiUgTRsVlEaj+zpRczFmXMl43qtL09bwwIxc2R+Nz7TMadgRwezNndB+Qci+e3waS6db5e
sUByc89EzNSxRZn95fbfTMrzJWL4o7KOdce2X2BL5IBFsCH9WZPXclFGHejlOFukLWkvFBCw75w7
45FeyB7UfDh0wt10qtw3eIqK6BK6dmfUKhqI4w+Bu6Vd7Dq2kaW6ROW+bFt4Loj/CbItgbh2OjRI
sbTe6bm21vYTIXgRgLoNXf9u4ZhQqepUVPkSYx+Le16vn38WtsknmP70Eeh6ofdeJUgPmk+VlRJR
BMsDirb0aXzPnGj2SkzSPrDJupLbNoxbPjVEKJErd0dfMWpd/hD/B9bZeBcTtO3tUYT6kDF2UUIg
g4X4MZk+uILarhui1R3776ZvqlFMtVHVMHCXJBOk9e7uriBhIBPEa5pk+osChiFGxvrMrrN8w7oq
UxllGRfH6d4+9mnWR97+1LsCwYjiFB2OICeKB5xY/c0FYZM3apVY2iSeYNKwFBcPaIfAWNevDu6x
a+V4saUqdr+dSpEHBqlZ4YTK/EsEXW/xGqxraZ7EvvB6qoU7HMl/QThRJkgLS+mdUj6ESUpRlqOX
27v5gWLlW6diPMU3pS8ENYKSguQrnPyD5LY5ywwcvitiXPmBLVIvfu7N9gnuS7Era4BCLaj/9SoH
DFsjpavi4MdHr4C/baZD0km7iaiAvZTpDNTRc7H3BMWGOZPBOtLXJSM85DbN7ZDpmv6FhQzjZIhW
OydBtFZR6PNpJcb17u3YYSfd2Nsso75uAUDqbdSjLuWQoUNpQ4fD57ktCErqJ28g3akOozV1TMBx
B7/EPW5FpoVbMzEJGUx1NA27VLALDA2ILFT3/14lolW+JKOHLDOb8v+v5NrAsoba+G3s51/70uvl
nzliWGXy0OJX+Qv9X4T6kRnFomkss0OjYn3RdQA1JffCnB0cMkZqgYfBZ5SKkB4G9Lh/RQued9NV
sjMeNp5P1/Yn/qaMSkb5uR4BMY9u63usd4NQy9SIQJ5G8LFQXdq+mY9/o3iu+R4net9sfQsQtzEs
Bm6NxigjDKbMCXRQuV1vt7gDad3GkkDAbjH9ys6YGJ4ZPxNgNWCSz7lE7JEAQZsdSVcwy2buy9iH
5sili/XhaSC7bxQhAlYlGByRTPzZNgvPx7ut2y4Z4JY8Y6MxwGScKdCisggNnKnnDZa6IZFvCfFb
lIUV6MTovfXPofD+wBdHGL2VolV1LOQ2vCvLC8Gie7fTPh+NSM0mIka69JqKa6qmAcGJX2CA/ZHk
XbpuOk9P+tnm6BSvM19UnMr5ltZDP+VQPhRK+cJggpnMih4qdQROxZ1sZVwdufLEHY2beo78wMJD
aleVt1A6nOuAiJ48eRDuw+jZKhBJsQ4rfyU6ZuywjaBE/0QAtrGGOWbnClO84IzODSR/mlL+Ood2
i6uktOInOflmskn8ybtIMQAMGi1ja8/Xm9JqedcC1vg3O/pIbPMfPUCjZ50LXgCPO8QbWW1L62np
J1f7jxkXwnVTgDZeoRUb5uCLrgx8eVz1hsvNDTg782KnpJqB7KwSTU17vcYNjmh64xKrKm9uyQPl
UdUV4oXYQCoQUBnp79BdpZJRaVX06ZtF0qzOjjOl4udsT3UZ7F6Rq0Lh9jBR6gTntCNAUuM3XuZC
JXCVaU2yJlv+EcPiQ8TRE2K0N/OivFEsGw+iDU9/m83Vz6qqCgAgwe2a8+y7IMMcQuzjxN36PlDW
uIiRGxF/L4Gikr7IV2v+XwuoFFA3l+DHb31RSkld+XwksOftYu9eSsJaRsxdj3I2UPfxrB2wnyrg
T1o+69kUP9UDG9tgk1eu10rgzGRfvdYvw05kEReDZSnHYULOlWspacs5BPui5ElSGwgt7rTINEvS
oL8x7rBc5taFsDDAaOev8lvOPAWlhGlFDkq3QvX1ULz2CAiRy7wcHW1vREEfTeGx7Lr7kuUKJEZT
rBdSqMgfZGShKXIaynGPsTK4nXMdXyBkwxJuP4T9XU+qHmPHxlm0BtpagKVr7Ay2poYiSu9JR48B
kd2055Mn4u3Mpy/b3X8bvCnAJMkwSZKAase9LQpVTTONykpvNFmTScSTQlmh9RPZ3/y0AmjH69nE
qwiVQWeSWshBhhrUXrgPn70eEdsothdSk3DjYGrdYK1HhZAQFjGag0IZUa8/GBFfW6bNuqqJVqqv
ORQylkVaDg9QsfNTHBt4rkox7xIk3h8LKvhD382aeNu1vCYIDmnILQy/pT/tTzyvRmykOpKh6n/k
hfiSW2XByR1iSzCNhT2bH7+OWntpNUuA3nAwHKLkEoOLVwKLA3EZ98HZtvI2W1JUAa5s2eeepgU6
FIlu/QTsRjmsaoaYNVIxjP4ArqAA5rYIrTpkN4JJTP6oNDyIgORDPpKYDdWeF8sGTogj3b+5OdoY
SNRYM7MGXP3nw5ZAz9rHqCKzC0ar8UERYZNRfZ/G0pD9reE+b19EpYLyiTNjlz9pWTGqTopIYdkl
vAOyQYGRkhwXfAgX/ST+7a55bMjUDfYb6vgW5RxMY46O/LvTemNjiuI3doQpqzcMr4TWUmnYlC2t
mfl4iLPGP+W93BRyQqgMV3S5WaF5xwUzsKTblQXnbbJke1PS/Qke5AoUXlcJpBl8dlHKdy1n32/c
613/OS8lylOCtgsIWgIwXc+UUeFSaHMPMUttUo4BND7k7QyeqDkEBofJG1gbbFub3kxrzemZIFIj
DPThTrN1fKdTw4MTvFWIj5FmComoRY5bhWpk3AqfIzDpW7I1sHgTivKYtWHg3kwFIpKaCisudZBQ
lG/NBKkb3bknnkh7NnRDNeH1Jq7yffDk8nyvJur1FXsFD6IjwIp9/0j3aQs+XbFoulmxG+SE1ILe
Q1xsa5JfTKn5V77iUZIE2zjnewoRUG18H6cUfQVIBqhK+2YVB6uAmp/VStoj26dKSJTJEbele8iO
hoyO3Gg23oRzPuz9+8u9cxr682f+oGdSISBH8Rgf5QLRsnAMVyJFzJr6EpwQj0Twu5TEoMlu5AXH
ksFwy06b4v5iITQvVwbjwLn4Kg/lCRXgs7WjPOH25Kd6F4Vs5A1CmmTsl4oLtsT3Xtk7Rhmd0Ec1
g53LrCGDn+crec768yBuV50xB5Zy3M5KUa0eVWfieg4SbLSpjpO5uBkBh3ly8dK8UlP1Es0FSkdf
GmpFTHDncorzQe8M+xbYp1A7vfBO02HAULmjJeUOmQ5e6qLVTRAqXEhaI6vOzddGert/VUiQ4LTU
TiwW44iiwAQ3K9S39xY0MvbusaiDkl0dX98fZwj16YIoFuS9EC8bZp32uS5GUwG26rEa8oEveGfP
5GSSdcmFxLSoF1IXP02wpXUbfcQ9iK3r07LJGCVo2DO5IbVTfKSR6k3YWxg2lq1z9eHh2Ym9pROk
6gCd4yUlxXphZMw0ufiWxVJ7V+e9wHzODNGlsBlBmIzJZFbWBKkhWfG40usTlQUdiaiA0GGegrgj
/6p9m14hesFiaK0ArEfIFvd0DMYMs/VucrfZe2+8HWYcCS6ovUR/ATb89iHSnm9VrBtacKfgefKw
DnX92fAnQpjb/euQ/FdeZP9b4/xg6UxvX+h3QX/dsZJ4soapLNIGHe97ltaLDWUDsrjgWmehS9Jx
nsVdvcRfD99YWwotQcu7MMxj5GK6YqHakboNHnUrhOANsJuDkfmTR+b/elTnDVpYdKR/DBceGshs
MsiHko0DMMQl8ER5NKmK7LE72k9dh3sgQXvsY7VGKaYFPibn8z0BqvuisG79tv1a0CYDeGHr0f/0
aU9JJOROGeXZEBRMwF4oqXrI7sl0uJ02pVEOSUMXR8PVA9gUpNSovHJvF7TaAEaPd0ixMiOkYwTL
Ye6MkQY7bldfKeXga9TX2pX2QVl8DsEBMT3NfROzLcLctID0SUuX+1YncOs7KJYbM/kHJAsYBZoF
d9qCRYPkEzwa2Mu5dUexgeHK3Kfrj4HaO3JrVbONpkj28L9FgAi5ppsyUPngOzGZ/XC9X1mg2jDm
K5R/B7lR1le9tIqKvzi+FUAn/3eFxmrVc6e459tG+aVvpdZlMmuKzrwzYevcfnA6VkJ1cIoxPA7J
b7ECEETfOjGeDvIEAWgOXWeNmWGJbH73iKWPwDOd0jt5Zukp9rcre/rFKMOuOY6et7kbKyPmuss6
fLFbsuUer0Iv9iqtDMF560ubCUCGBJOJ8j//HfHMEsnniorF4LdGOue6OKhtbDvoXaOKl78tdN/D
qxoC5gNUDfCWcp+mGdNaKIR88To6LB4BDVLuVACNsPZkxUJmIaFk6cnv8pNZTVGulbQlXR0qdRzk
BrwshmpAmPn0S/oLxB9F6b5rs1RtiV9pDauxDgLl3REfTcQrFPtKeJUSbBtX5sQ+8JoZ6PJVIfqX
ulSgPgo++3EUdOhL9QitZjzFzNE7k21IMSb1z90Bqzq6gEXFIx/EJbQ5AM6CEf+iDNoHPCP0Yr7+
QTglT/+7DxkIe9mOSq8KTiJ65EfUrfKSL04tR4WKUILx1szAANQhfQLBdDEg1GRR3CFFBEF4Up+Z
k/2F53F4boa1s3j5GYaDrZS9sgZ0VXHA8bp9Fa5k+vevF/EuUUnBUz5jRU1Hf1LI5lmGgi+bJtuA
ZbHHWjmXmKX2A03DG2IldG3pO+JWi5OnPOSFcL05wyTUcwAT5IXipNO4Pc8rtFGiRCjfPY/tGGuV
Yv3cZZmyUzMkskTTZg8nZisn7ek+lHmJ9CCB9vwKJOuuQRrY6tIOA5kZQBJ9cqbveL4hLOQhq6ii
br8JdadS/AI/+VNAgZwFHXoXkRPS235QkzE0acrHOYWZmvBVEeqf8srkwdPXgaySqBldH1SjPBqW
hVWehoau+qR5Wj+cwpzkw7y3JWVISBTH/QfTnzVa6mOaTxiUsdH+zBlgWCG1amv6qYyC+o2JgGeK
mrtZAz3+cEis8vTHltc6oOZsiCcQrxuY+o8uV4T7KBVowwJvdlFSzocOzxB7YyhjWj3OeExox/im
83cruzQOHScuiVHkcM1cLnJi/e/0zDHZVud1XVR0atrgAkObf9zOKDl8pz2h+u8r3fHEpYVeZofK
EO2pC+XsoU2CnJnk+stsgASxJ0G8D63oc61DLP7Ut2Ry0qPZ+2BTpZSN1LoJ70UzJBQk6+Al55AM
W2TcfzGFytpcaXahdW1b5v0N20qrkOy+9TcsF8qXmeZ4EL3eYkmpv7+ylpjy1/2AueA58geEHzZw
kzdulJjqSIiBa4WzqOx8lNeIJcC6FvnSUpyUe4LbEsfmgrgfuVRTpVEIynL3OrZfAClA4PRvGfFZ
ox13iHIM/ghMaqP2HUKJJ2uD+y1MEUT0uCyMnSffgAFcm4rZxFyeRdsNSdjBiuQvA34EV9JYEcz9
KzIbpzU8EV4pLSl61ODB7XRLw/AbZnlAOVxKTqwSa24w8ENU+nMGEmBvj+qVCnGmNO5+NBsXteXp
T7LP/79mMp8JkyW6kgZWeFjrPdA8/sn3WlEOcD4j8gR01rTyhRXGAHMRLq2LJt6nzPKfzdVeZ+Cc
sKMk/xvkmjaOaVBMNJlMdaosYGOHhYUVK8wqHYtvY1yV+aw4WKEBELFSxViCq00rOpswOREq6hAG
pDgexHqsWOt7c3bJw4noL0gbLMjiCWoeWO+w+ZaJg9S5suN59wOr1/vqd6lOBbHPnRvDd2hxPE/3
1AaW1i+FDccDS4tpxEyv9XdgcVAyccERaSKZbLVji3u0msYBdk1Xyg9yLpdnuRLras6c1bxr7/IE
Aqtinls+bmccinSbjH80swj/z68oTVY3xV29hR3oOC7UIsfE2o7ssiXUfVNeb/UQNdtWXoBFIhEN
RO5HbIi/gKhq9s1dAIlUAB2Cevvf1xJ0gUQZMSqQ7rOzMpxF6gJdZrzRmNBi+1EiPQn+mdyolVuZ
zJDE5Cqx1n+ZFSKFqE08jNkGE14K8m325GZ47YuSXiz75ulD9ML1/IpmFZF3xsDoaqz2hFAKJIoj
qPFqx+r3ve7bB905p16a7HoyJlZ0QcMh3Io5f1jMEN3HTLAJAUlM7IBJGDdBe9IZx1ph9/peoST0
QrKMm2H7bKmJLlNenB34Ao7eks9Xl1+S0nEBob76hBPtSC3q5R4YUbigef4qPwymjWWQcFPyvtlS
U3f4sB1Mqmm9AeGUiRIiGCdZ+FIwq3XTJv8mU1PMArox7mHIuSujMls8cCcww+/Vi6/Ep6MkQCBT
HPzpRk7OBsKwtKFb2rIBw1Pk0KWUyAjfEC8n/s4c1U7RJIh/bquV75OOwiMNYcS196t+hYd/2EiH
GIZrWOqZ09BSo04mLKMzfw6/kYVtuKGgFCxhXSWAinL8bMcPEcgHzy9LZJmjxYaeN/X+NS6A5aoP
/igZo1Cd3ZQAaSp5O63Nr5/GFv1N+AE6lK9lTHtPyADSggKxbZhTArPRBbBKVnq4cFxn0FdNc3BZ
biQ6A0j3x64BQKR67roE7NsWS5E+Fv2igS3uiGgdeWhBUmq0fRc2/fqizCsRqfVxIWEXq4vdGkKr
+5mvrAbBelVTdBotudoHAzmAhBG5pN8wkwyAdSthKpBJGXKBOGjFjpMzFqcchKrR8jCZxBy5Ez20
/SkZ67xM0DN+3iB2KoFtTer+GqEjANy3RvtEvJfZx6skd3D1fc6TwXXpW9bj4anaDHv1lg9YLGOJ
UZP99CRQ0S1tD9dmiKeMciTHBoWu5YDamJ13eKFWdKPB/hOae4IFGXshOd4tGxJby7fo9GLdxFe3
sUpZioKZLBjwm9FiqH0bf6E0YKmGIfolAM+l0uqSJAD+zH2zT+Y6qCurSxBUc249QrwHtg4aAi99
7rpPry1JSZWS9JICTDkZE1OwfVMMf7re9xd3wsVGThqMmVHuvhi4Nd8KNL0dgpp7Cu9FLD6Ykmug
jGKmW79080t9b0nm+rrbJ6SOLFgyBmG2wxS4WLdVodZjqmXIo0vW9XMeW3/Xrchrie8ZIFVYdwCf
PyHraZNymkTGQm3MChBFKF8rQUZhnsl91GShMT67ZNTLbiqTSZCPu3O3hzy2Td0DbNiBKWruOT30
Fy9YQ1KHp7NEp8aUv/L3uuIDIyPSWXvaz0s98cMzjyyY+6/Bv1RMP4n9zdP/TjlCiA1hnldWMJcV
3TnenaK8sE8FknKDzTkZqcqYTtJN/ErGRFXfvRtNRMkOQeItaEfydLXPU2hMCUaPUxfRvEsz1pQT
m/bW6lp3V3JEZAhE8+l+c4GMxH1gvZrKP4IchFDqiOXGLq3i+qOo1lkdxQRDu7JzszYqNVFETgnz
iBCtCc4jwiBli1u0ZTu5ipFrSy8kqEF8XYNsvqJEmYQVnU1av65efzq3G2DWJEt4U4qQM80maPQf
mvHlPGHxiDlno24UrBGfGkaI0LRIBNYQyKiGUEIuZgprvP18HUJAYzVddt3dFxAAR8KNmbYoVR6z
hWZxL1PNiTG2nbN25cgLSbA65zGgVBFAxb40Z5fARPuPo4LI+M5U5V0k2NfCyfUVjdVdcCKEb6N1
LR6Zq0jsDLmlLdhFYLhiPQ3oZumLiZZOS8GMgUgXvQAxMvjj08IxUjTAAct5G2GBaDHFhB2gIYOr
brEncMJ0R5OXdjr+u6Aeh4XldVJFkKKAmqDLOYcf3B3QYjGUSrMkGyul0H2n3cfS39r5pckYytmk
ywipgu/qIy1fxdMk38SHSb1UUl2C00xEG4fXH7/u+liCJ9O493iqjS+E5sYPGzPtjLJgfiDRVcZo
Rqfq5zzsJ7D/K4zXjUouambcoqo8hUAOymU75uOvbrvtROFiFgjQWCmUF4cIkW7KGMErDuYFkw/3
Eo652JowogAk8V850jX3QAjFLhov3Ux7cjZvrNsKAZZKNjJGiweFBlIAX86gq5XhLXkN5rV57LRl
ohuth8cTw11/96Bvg3sMAfArpaeotK/BCcQuj0OTN8z9QUIYBGbXlWcbobpKi5U3Y2K6FJTLHPDQ
njbzhQckJtHord+ubKloLgO2LCFttkawCUhJgOlFfOYQ6PyjhecrHuIwjVpEAQMs+jlf+0LKx2Hh
IoqA5I5RkA4zVZp+OjvINnYXFGHPMhLEpeV0TlAEoOiBkVZNENRGA1F2i/6u7yrJJTXd7zRWbFX0
DrJ1DPt97VqS1LzxMplMf1ZQP8POyCX5W7VoAJgR34tB9HT8jqRbDAwM5E2fix6nmwRY9pL392yk
TQ3Kl9XbUhS4BRisaZbQk4m4bXAZBxwDCFcS6KvHLbweNnyKHuunhWqdbpVTEQ1piFqLMTH31Hb+
BNAMXa2wsblUBvy5OEnJX+B3GUPVR98qxvCG+bvV86OlB84UmUiZj1mHHO8Qhf+SxQbBMo6jsPqh
L0YTdRBvkepTLdtKGjXlNheAtWLD4JbfysbF+QFFNQsj5GeRxE+Naspfb5dHuNFSsF4SOwiehX9y
wc0SxQM3pbhrxS7LgIobaPBsGOhAUkDdLVtRUlo0gHhWuGpfZez0FpNfm2bJqge0gONMNMI1M1Pr
0O7EFNw8g6pzL1+cjycEx4aofHpNWuioyzZNyARN5j1/+vheakh7Qr829sXmxct0rerlb7lLbuhv
XBs+2dbqQuYyfCH8QP0ZXapNg/l9p3mRL9Jclcb1Ig/DoF8uNgeqDhVtzVWr531AMP6InhG2icFs
Nk8yJ1IHZEnD7fHHsvOy1U6W7cv81tXWEjJ2D2uMJrZypXQ/9pnthsluqdMSlq8BTySCOsUBVe+t
cJ5H4w/N04csB6W23H0Y//zu/y1eA4RmQcAv9UmUVnFw1doKQv8lV6fAuon6DKE8xQgWmJ3TQwvj
eN/1i07mk/u5mPYlaDSnCD7p2Ip42dIuFk64z3gAhpsD8LrL4EVMAM/LFfimh3nnK9zxCmQ2hqo/
9NZ5FfhaJa9SHHoXuF2dwG/RhtHLaBtEZUa5EffZ1i9yvC+RLwAaYeQsZSB89+6Ej8n2kn5jTCqg
WJyZlrXVZBKc+1IUQwCYlQEK13YRgmOGgEPxAUG0bWTyfqdTMwohsv9L4WCI1teoheYlE8/JQsOn
PvOr6WRiyk5n5EzVkuSXghsGk61T2KutKsyQ2cc8uXwg40v1ilRyC2jxKXIFq5WzI8N0PuBWF8pR
mpLqV98xI7zi7YmAII5TWLqCFR3pclwc+Ky7NUMZyyqQB1LyE7lXLl0y+/w0i8iEK5ZVBk5nv8tk
L9HLl/6NP8qllyPuNU0hNcDnR6ot6+5U/qmHHgwxjkCs7NJHzTFBWv9jtjjCCJSbl96OG1vWzqCL
j36fMw3VKtd3F4tUWQEmahijRIVvJs2W/yDNfEc/kcBv6X2yE7Cvu8IzP77/4JRktCujuuqTuUmu
JxKdXTFNpk5hT8UHbkRf5FxBSL8Knvq3ZNRyh2axszazKu4UXqhfAzZVw3F4siV6g+O0SCqS9s6k
6jLIuhvR46Yx07NwV8p9vv7r1ucZ7z6l4zdDoTRNtBdLq2suYbL/cgQDz9KyDlzfh3RjGzGyHO78
Flvg77Tk8jn/uFiuxo68jkWye1rvhDndw6TMtrcnAl65jawZiCmi1nNTPI92lesKTIP3oYHXihPx
0/qKlgXGzgUNeexOGrFLdOEBeN6IsPlwzxJbN1Lfc5S9fo/tSz9mA8HbiCyxFbhimH+gFyKkqTFM
UFm7Gj1ottIzngdLkbWEiL6ZWpomrYykUgdxXcuHML40yB4yiPF/8lCiGaZmr/WuiH5ILeKMhmiU
Y8Y7xXkPWDtnmHwzv4lghx2CGU5ztMabYTBSjEikDSR8GDkxaIJtZ1reEX7OIsABJZBb2U01Bdm3
WWczSfiptj8KL45p2iCOfYn2tNWQosurPdWxLixY2bQUPK/JDFV/+xN4jc7rHv786iek05Rq7Z4i
T7r0LBbjZLg6MHQRO6HCgDGSBVOZmaxnv9Il52XpfIuvJhPaHbEYbK/nGegBMqqROSAa1cp+gcX7
6wNMR5+0O5FWKwOC8fWohQETTdlWwZAb9/GoWD4DJhy8TFAEBX6prdbppdznCzOJ6mvjHVoB13va
O2c5AcJLXiuOtUPKF+9UtNkVhWLKnf9WdcVmtUaFWIBSyZoLgGyRrt/qQOUOtP45vL9Ppls+wwGb
26Ppqlq5J+MGa2prfjJrsBB6x087C4hHhmXGiVPD8KC4m+4jNCIGM2dZDcm2O+j9pNk205D4hTPt
BO+9sx9eEkkAGn1pJyOo7peW8vSOeMYmEKoTyhIbInKZzu3Kr+WQl9xMM4mH5zbPdSiBgGI1I9kM
BqdWZxE/n3KRCTkSMYw2ESwMuQuTmT9f021Nd7itx08wV7Z3u9I+u/L4v/kIupTR+M+XdTfBhstq
WiN5fyZ86hmfXQOzMDsHWQws3j53cO6eOEtsPv+yDTwtuN9r2D+RQ494RuFI5EdczvbBlMj76FJ6
L0uYs4uwJkbbX9mh1sVvtnSr9XlYhO+HfarNgsM0cIKiUUpuSFRI5iz9NYkd7k+7NcBRtu8KWtDq
epRjjm+8zzY7ioR1Ts4UQRuyEAnU9JGAPltbSpOzx95SiDwkQ2D2L/O3x1MmoBgxjd4vLI6k3Z+w
9jqEAZ2CsCj9iQnETpxh4jUMbjaPrYdulukgTwtWtkpOmPO/RytiZtjrsQ+TfuE951fXjTYil6OD
xyBv3cD/IpvrNFWpXxRuHMiAiSL8+9zpvWPCMRNYFkWo4FubUyWCbBOh7Ny+ne1weqgXPMU/lL5x
jZOfiL03BXWak66uABGjQapGDgn6d7WykPjsB1eSGmmDIXlGlnKkwRzdEIK2KhOyuOd0dG6dFMeB
wFxr3L2IxBgf2fDOTX73vckt05xaNqlw8oxRx5v/AIytX4fKZfqXGnylZ5oVP/WvwjPgWRkBWzAl
/HN2udvDtSQVdrebDA2abrc/iKcrhqhd1xVYZnJwur8kqsORqwXJLyogyZMA6FUGYexlrhdOiiJ8
kp8UTs0FdPnWxj2YFzEiWtAlRuRGscskDSsp18r8zt0j+H98izPjkPuu8mNlE85RsdQLCPwJcgHk
rnxLE4FEn1qKCIFkVdv6z2sRWZpEcYhOD0JzvUW4/coLC9VmXxFn78Ni7YtDD+3beU3XBWlIhwFs
7VZ3BnFOly4nFqj/nwTOZCdsVH9amxahpycdV03VsYlaL0ozlma4LIs/wz4nlGwbmn4gYjg/mZAk
JudU13e3kEzMX9kewMhcFuskz+lb6VE+y6TDgNMbTuTUeLKX1AswY13m4cOc47SJGGlRTQotjYLZ
IBj1OJsl5LmBtOGR8wCvhszZHQvnuisE7l/BueNhQMLseb0lVDPtJWUySQ898rTVAJjqFsEk6ZYY
9ZI3DXjLDedqG/bASIg2wwGbL7wUi9M2fT3R0xzJ81LHHnkHd+NNOx51Gv5kPiRIssdSHA6pENE/
IQlbRkKubqHXMS5cGAiWs4xUtPqnKCHwoDxy2wdBH3uG7ARFx34+sSFgsrdJQrbevQyhvgdlcGqs
Xibu1zUjnmxWTcFh4baOY4eFe1mb4LNjhcARBBsy45khjBFj4PJlQEZzo/AkSjzE/Ex/mYYFbGy6
CeY2Z1nWt7HCo13C9MIwswGFicgkmZ98MYYiRps+GO9B5sCBzwu5vhJSzo7Ism5apr+txKa8YVVx
HHvH1vPMDA7PPlPflHQmeEEISnxZD0tIs+CRW9wExjt48CsT7SXgLyw2BhSE7ytJqjbcXLx5NeG6
wmKKLLNU0lyb+CnqAt6x+kV+eZG+Ts1O0fgEn74oqwLwnaijjfCHwNDjO5bAbAu8IglItb1iDqVQ
E9r3w7pSVlocW1LGxIq01VxPsLP5fv+TmsIQ5WB2KGgEIdKheScfaNKBhcpRMdiKPgIuABXEt7XQ
z1LT+jKOIMM3lfnONOJmdeDxjcGya0/qL9qRIaSgQmCX+pWiS9Y7LDTJBxD6PUN2YgtbmWXydrlc
eZx4qfTni0tYNXyfMF6/ATV8ckEK0+XcPPgQ+PrdxF2o1scsQJpRXR0kHamXY9er0jWqslfL/kwG
8jJxK+GlVxw5xQURn/vwWoE/fy2PAoFT1uIdIzGdT8ZiLbfrkHW8EAFd1NADmckPRRlUWR1AdzHO
ZOTyN26/0ld1KV7k7DqSZpIiY1H7BNiAJbLf7o3ddU2/aDrGbUrnAn6yXkMmYH3rYNnsXDv4yll/
BaQNh1QXgZtHEHUhVGn1JQQIWsiGlYk70rkn8rOHQfV3aGrwqZcZlhhYJkldW+CGOWm9JtuknNFa
OpsGi1JLnN3EhPwcAbN5d4pwihuWR4KM4VXwSYPnjKTrPIVM5aQMgmIOmc6iQZagu16groJeFwi6
HAz4JVy1cqpbtgCdImdkoqNirJ9nhaMKOxd7X5G3tJjuImCKMYwzdCnhV6wRuvxFFz7FrOHl8g5J
WMRvUql9rr4cMzr5B/ycU41bwfQOQeOLV3GBaxOAL/ojP+LA1n6yeSmoIOBA9X5czMv1VgWoT82O
fTj6RbVN2M7hEFQqEGHHOO+9C76z9/R2kHHWgsRaycee99FmlZ9lpkH7g+nvhciCWo8H8v6sZrvP
RvcjRwBSWB7m2BnY35R6tsY+01sf3Gk0oyul6xXEjUBC/PVYYQyrvSAvT8+na2EioxfhCfyF5esb
eXzB0U7dEGVzbaUCaU8GtbYDrd+UIrbpXiUxyZYCATFbQE6a5XAhEzYpqDewVtn8gGdrw+SasSUM
3T8B5fdZb/x3LCMp8GSOu+aVHtA6z0OA1iXxeMO3UCZaPiCfBaugEKSdddEA9PKzMrERVSEU1HJ6
BcPPsaisGTs3AwyBiNH3XiVlo8WiMGE96lqVwwlwM3HLHTr/dT4y3JCVgjj0syxoB14ZdyxR6+s+
FD8BQKxm4cwAuWwJdS+SXYIxUoxvgHQE5UXNDFU5R4ZLbJdJCize4AwjrY7DllriHU49L9xWQZCH
c8o+3S6Rlu7NC2xXTMwOUXNnsoB4JPIZfGmHNUA9nA67diQzoHARLfwhvnqMfns3QdwVSdqvRIg9
UPnehOcUh07S2VI4EFcVWvPMjDq8t6x3N5gkTniz60ow3y92mJyqnIK6GRFAvukb7VmzR92c1/1p
+Vz7qpsXneAD2tnW7N4gMpgRZnVUDQ+uoUDzEn1u3bvnRSyXa0caW5O3+T74ejZvn9y+6nV4BQcj
4Q3wGoVmykUbNM06Hm7JrmkeqNZFswcVd5oHlmoS0jbLSyqeTfTisUefldLkBgPZ9Av44dmPk4Xx
t5igG2HKyqRqEveLZbFPiYIVdIBkcyXwHdsVfeNOsYOSPmL9UtZduGCpqMeqlUbO12p0ZHqzuEsd
F8CD17xNNPWHTxxMIm65bJGiebLGjgHuh0K7SMZh9MRamcmcDwsNg5UCb6GgoLu3c47+ZuzD5ugi
PGb4cN1zWZ00e9i/zTSnut9PzpP1H5A3FkAb2UIyYg/d60JfroMwsG5b0ygfJ8+tGEiAlp1h7Idd
v9WBAk2nJiCQ+uSI8/nRQ1NEwW9nC9Eq6knrQeF6KoRX8iHKGf84gsXhqqfK9FRxWOprpxrlseQm
gLUPbMrP+trWdwJpe3sb7hY6hZIQe7vlMT0sWXg3aF1nzmTkaHTUC/KIXVoCwmPPzfO17WmOch1w
YEmoTit4G149Oh5bljjLdd5RyvH7VVrw9AG/yg9sRvcsvbgcFkAAELf7QJUe5AiZG64QZEOBZoLZ
FGXE554P9DFJqs1Sft6in0keyjbcIyhY9Wx4q8aLZEvzZEhb7CXK9au/kLkbbuK2VEMexLF/LcU6
QjkkLVNMqTSV43NyjAcKFio0ZVlW37kljvMGR3wHr9+krv5d3c53EQIl39O6hT14H2cx4xn5xA0A
KBHFQr6nVy/NLGKnvxmTMPsXZOdt30PEYfrpEBj4lrf+jPYtOeibQmxf3TWWfsLiEqIDdnmmFPH7
WrL/+ijIkavA17RPC2HD+ouOeUo/eR+IpogYgcgO73OvKWGx4Y5ZQjd7gUD/PVTVTlYLmm776gl4
hjaJSqqNBWB76nXrdfAxV41N4h3mS+MSbLYq6LWJJ3AvCP2hgrdlIBf1206q97N1O0iTmai2y/kg
dk8gHDFxrmCzLHgf0/6iVnHYvgXptta2/uQ4ZCAagcWxRih9FdCMHMuALaY4J4+eGJKMdesP4VpP
xNAxe/pjL8X1+hQZnwPXkxNf861ov7S19r9i5XjMGp3yqd5RMxTmR8tQh69rdICWogu1Qj/bSaDx
yUt9mFeHm34w3f6kQk2vHsG4XVmus7AK5U8P6Mo1IKmjlDA8T8iUnPM6amUIcgL9k7z5H3kx8SK1
7aOZb0Unqv/5d8q8ZY5GDZMnQhrQTK8gfbz2P9VdCOBhJBX8a3jYX2Fo60ALA7QvztsTDQsN0Q41
x3FZmn0wW/Pfyo5/vBTFVimvqmnuWvpDiSKFgph7yYut8BanpQOBy7cSLw0bzK5qvogOihaukZue
Qdfoqr3BGO8hi2tiiAfkJFQ7Af5W6uJwH7whRcNSWs0w3Ay4Az1Z1SPdUE6m4IWT5TQESVBXhQLJ
7j2vw63qRDOYWLzh33ZH63N7So6LzD0u1QHeui1blKnhSBIW1aHYMpoWyTFqt6ykWtTjm7OQln9H
W3+y0FRLufboi1j8ejenabS8pKuGVMp9zcCsLqakiiwojlLhgrC84Coh/BMGpg9T0c6pMcgxtKTF
nCvj/Eube04jnTcqi+0POmoeuoA2E2FD7S10NtTDdu+JYdYlij18yTeoivatOUqFhOuOImulN9DA
tK8eToDctBVmwasGDulScVj+R0obvf5opDZGAXyIB8bPbgzMYneLMnwMEqdgpBombwz5WrJ+Nfs+
V0vM6SP0lM3mO7Lxbl8uMNpCAy4cggo9QotE9xTdn7wAsc5ZAtoKmbBaPcS6ur/SKQpfZxsZgzRO
2BgfYK2qKE3nfa2gHdFmhqve2fs3PAyWgO+ddNga+bTNQv5LCWlh7k45epXLk0RK0Qj6ESe8+Rl/
NNSfn3xVhtbWsPpNF7SexiG3DJC+oEDcx7NE/gvUDjWbWffy7LxTyGcv4u3qDMpNGbHEQkiWXH0U
IQhOb85lSxhCcFbJf7S0G0IPjfM9TFvjghhECoQwjZ/sgk9lKB5DgA4skFATg3b5SUTyxvE7heTA
Fv6ootgkrF7N34WPRtNouoOuDEGsTPutZEOUdHhJL3cv2vDtB9VElUqFAdpq897MVs4FaE4VGdKI
CN5m2X2J+fMqcBrv4PQ9vx421dfLHys6IKOHJ3SvuhP0iBjjM3vWbQB4U4JLPLCsse6e4flLxCJs
/stI5Ewm2P6QGtlD1itsyYihF0QYE5obDk+A5rIg/POm8hDuQwZRtC75DpENEzQmhGjtgY56+Bv1
svSEsD/9gab7QtQBLfzheZwOb488GWPC0AX25LGuuwl4VxONn0FHFoVC1Ao+5CCeFgQ6+8O2VLbI
zmXnmxDMrOyeKFHo9xJT4Si0oEukjj7DtQVinbP3mrulwUAh2RWKB9W+uBLxMd5mMb4JXhdSe32M
BdIbZztjd86YS3GteefMNg+Mk/jcVA+Q6EuTdy5Ogl2voBFGktGwU9a//AaGXlN/9MMg/nEshtnc
Oy9Q+TVD9b3ppg1lO18iULYZ4kAsxdpvd0KWxzTCSFwjGyUgYkfUE6ZMFZLKUOSr0f49rUluCWd8
yZDYBXtsOEGfZCmDYuF+cBBeF6FvRx9uCFwbJXiRSAvXl4uvwAOsebvEi7hOV0gri9thFV5+H71V
0Z20Th0a3pQLbU4zZkh0x1do+ftvnVnwnp2JL0hyaVoEWnIBtn08eW7//tyNBA3031kD92tVHklS
aYEo4i0YBf9JR1UFzPdwagxAy56qKjs1RVSKQnsQJMj9qF0Yieuf+xJfGZTw3o3QK1/Jkta9BAAw
Haxpo3cGe8kFIuy2d+Or5C7NoayXfZjYYRzAOetEesXUp58VkFbuMFcY2lsowet3PtZvSKsg5wSR
rqERrIq/HNBaG7g0qVdJf6AJga0VFqXHi5+lQ4H+1hlk/KjuytnL3cVZrLP6qH74aC7m71BW66vl
1n3srCuLXrt87KpjmYCDQxEwRl7EDuglciZrDR3DHgZYrf+jfPNxvNxh9l0DdmYZja1OPJ9EsWjD
iB4EwKuzCxFMwfRrxlltOMThEHM0KLxSuQRKzzJELnWP+/F+wBBt5xzZmatPl45/N2gkbaZxEKt0
IOW7CKB8gkb3fr2B3L5VtuPpVFjNoWBpxTnRRL+N+LPFBZ+U5Vn9PYeF+prhdBYRRa1l1luLCn+1
Z3C67+hFNTZ5ed/OU3TSjPhAE0RO50O+wUlKUxM9KVCTDvkMkjEj60sDNKs+1SdUKJtrpG8IkDva
BZyysEoJVl+/HuxxT6Qc3Dnj3GoDSOjW9Gs6gXMlyic2Q5d63GWaIR4jv17brncJe4RU8eX+JquG
5ngr0oZmDzd5Wleyqm0tHgLK/cxpoH8q6J3s30mZnmyEd+PaEIQgAXZmQZakg82C63JQP19boDzb
ddlxsKxmZO3beYFJl3ng9NIBpGPMJC8Rf6HQHFX9MXGUkKMOEkze5+WejqaafIxMNPLnlIiPL7pm
Eq/D8b3tqIbdj6vaD5LrL68gjbwGZtJi44xRgVfk75QRc29L7CR1iJdEdN764IJ3oaiYTVcmtSBo
ALt/OiWWhk6IA3pkZMdhBQtDkSQFgOHceSDkIE6tA1uCksW7tx1bh6GR/8jeD7q6MfIbOMztFxcq
abmugSOvMRC7s8tlMR0V3Of+UaCXMYg6EC6ebD1raqjxH5tRUHPtRAje8DMmnvYEqRl5mbcJeMLJ
SL8YYkxj5yZlv+b+NVLXufo2Br1iPtDVSYnnDw32as/rhrKejXptreQtPHwrOcQu88Wr1ty9V/gC
p6I6rUeQnEV9YbmVMmlUuop7hu+ouRc40NVjJjE805Ikzi+EpX+T0NPBLpX6bpLQYZIlqBM/dF1q
YNwS6L8R1u4bikQqixyoMY1dZGCAzRDtdJ/AQpFHBCrVqeimGqfmzl4tGVcBYRiOUMzYU+55g6jh
zJPOoAyt0bGAsck+ndUIa0upf40bqp/abfHgVfngJKxndvi7Ifz/taz9zghFj7eMU+orq9RUqja/
KiGT8hhzhljimCJr2LccW3r2vELieQ0ZOpDxUr/n9GIA4/yf7PU2L2LJiiE2LswE1fzxexdYVjqV
anXvn7Os+Hf80L4Mw2Rt87Be/Q9DSnGNihQPG5mh817Nt8VwgDFR+uXVH7ZV0yHWC7cAQhqvpp/3
ofVUSovQF3bVbal8wuVuhCLsLZUhKAE/c2/987S3FrnpM+cVsfGwcHEe8LELTicP76CkJ1Glrepr
UEiqE4ATho9FokumwXBC9KmZYQvenVFJmQdubpOaQ3aWUWo=
`protect end_protected

