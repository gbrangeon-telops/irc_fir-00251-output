

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pabZO1I/O5UlEfYaQEPwd4l9eUai0bqYoMxFZDUmBPXyS95K3GW98Ld97MzJKAXXnSlf1PewGW2v
0RIeWd32HQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MnYS98CLv6GUlLtXXj0MDq/aXJWBamrEeFXZFkhzX7OjMU68I3JzEc2/1UN3CHInfTII6cQBis+f
MSPPkhHYfjWA/UnlZNCfIbUjCA7v4zzzEDOXLdUwHhey61M2PDbtjo4F0M+PSYsHQUE61FCJYZr6
+aBOwyo0CpKkCUVEbxg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qncW/Cwz6DQ02ZtEcvyp5WdAA4sItotGPpP0REUtLyqefQhCtJmFILcg4T0iyRUg7VuYEwIANO5+
QvHNNc39qIJv9lOesalgHBZQgvNRJnIdYWaRfS0GyacwI/2JQRwAkuAQstvDCp4RTc3l8lwP6/ls
9Kgq/wnF0FIDD2zIsqBFYPVau5gOg+E2Yv8daLhsLbgUNkGI+w4/OZjRbQGSUjwZLuzAjcC7dEzW
IiD8iCe2E3P5aTpTA2tXeuvseQy8KOwVCxJQuur+f/bmnE2QrPi5PPQMRcOyc4ok7k5U/64SCKlJ
oITfL/xIL/xwZa26tMPcLgkkx7p0G3RLvL/tVw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Dnf6vaqe/V3pNaiPDsCpL4mEkUhuRTF8jsptuAsYR5QlsF0hNdnCfK2+aKM5H69faCvd5mpbM0GP
Pqz+qhNmOYPHdckgaTUGR5o/7QyV8YKLvzwfyDMqTu2isTv6FP6Q6welH2CNBnmC1/h5T7i+fy/Q
rlaoXYJxfrB3B6n9clU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IMf8iBP4Q72XIQn7cHjsTbT2wNsnwrpqWy35OTpGthg9IgmIl2PQf4/c9imtaZPdkPVpIBywT+vW
p0seCgJeCim8uHSlCA4Yuvzi7NiJqnEZtjEX9xSzaDj4EflUudOJTsvuYMqv/3kxvUgkIK0AS+U7
CWRV3RwJIjyzXaV3SkeD5i2xf0d/bezTocOrvt7wO8hz1n7ziicW5bgdFMZpO18+84bLDi0MzKYQ
Ad5OLz8QJgoCqRTe+B2lLXuByvKd2+XBYArz50J0pDfy4RubYe7FYpZdW50ze6dgBWVP0HOw0tLX
Pt7eQrmsKxnIhjnIQBRBht+Bb5QLkHSbaJnGbg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8352)
`protect data_block
EIOHkG4ptYddnJA1v9lJtVfOLekKTP4I0gEUQsP4cXJT3yeFd7kOCeT/ths91ILk3Uw7U60wj/5C
Fsey9K1Hykc1sVUWxWG+fRy/b1t/0oxselgo790Lqdd4Y0mI56+twnKIcn6wb80U6SwHOP/mM4J2
jfSSEXZ5zUyuAGWvonLOXsT0zy8NepZes/IVu8vZJhq3BaMHMy+SsOLKxXvvUSNlTutzELe58k7y
5QepdDRzB7tvI1za4zJ69aj7dQxX65t9wwFktgpd0ABjbNm9zYHfJa/CcPKeJiZhpP4HbjAQ4v4v
Q+PLK7UXWDTW08f7WlyfDSnR+zwaGvVSKN0QaA7IGVO+IRGq6C908eb/Amn1RndFbI4ejUzdFBB4
MYwMrILwWUdIYzUx7q/i0ClZzUglpOoHtk38UDzH4dBmnX+9fhrqvB+HO2hXSybTcrD9GLGIqyOS
cnpLINEdh0+TZb8sbLn6vmZY077CUBCOoQCPdB5xq4H7J/ifK4cvwztYJcQOzxX4s5R3PK0YBWfT
pzfoQm634ZYR6W7cJWDz9J0llP3WmNQ+oExp6nYw/22xzcM4017qBRsvKEXZwHIgUNE/LBCpl/lR
IW2AR7FYq7TPqzH4IEFNS741DLKf5vPOxtcvQjAx1VFNvFhgJPWr4p1NaQsfEpmeHKd0Z2Jsfyt1
UmHTxpyuTs8BrljqYiFD5YKk8PByYA+h+B/6OBN/pvi/NnbevJlSF8tJaptmvj0KLOjRFHuyeSp4
riNCzm1xl3p1+d4F+5wCPqrZNSGEU8/bOE5hO34+Pnl5e8pyL6apx15UcYqXbWcQFmjOkcnhQcPP
kZOmvtLsVdU8hnF1EcFPOpzE355I+wYNHCOoFWlMas2pJGdqkxVJAMgf1z21vwpAj83Bo9BYRXMg
5WBz+CRPqClb8h08h8GRgSkAv9tE3c73Q9KuDapVvnhBr57+BPwt3k+93ygvFd22/dpkTWvs7IsV
AFf3ZPusNlYbcTjsQbT0GZrKp12VOhMmnkP26/LjzP6kZM96JTDhWHbxfgjX2+TSFJJOkOgiCXHG
2UM77PBTfHURQlJvawoSAB4KLTqk86PHDBM6HyME2UFBEAtLxihvRV2T1JmxbXLEjs2kuBuKuvRM
hlhrXC+bUxwCTe3oTKo1DdY4eZEO83vI8x3AlUx3sYitTJN3lcNfD5cvJGdcleF0oKC3W0fo7H4Q
jqjNNQL6If+b1t9z/+EeTcQ2H/tNMnjJ45q33NAIsHhfWVUOU8Y6Lr1T38Q1XhFDUI8jzeH1EkhC
D9cI9OxXMayZaIdj5bSXiqER41SnOh9mxTRa3iKD1gL3UQkL+w+KqopGFpW413h6/2v8vPIM+DAH
6IY+8DPIdBht/jL8/U/Ig+rpxpTIWimK1ytP+3ahar02eY61wyL0gJ/aRdLjQxX1tMyevvnj71XF
S495wFzmGvsKuqb0G5KTGR0xsuyx5g8G41M+iXD2u4tXETwHY+yCy0yPLV4yjCIhdj6i4bdQ6vHm
RwuoHKwyBxvkn9EMUUbUCH1zImb0VXPSJ6oVmUvYCW4FG6uM6bc6sl6tnmtkp6gHzRYNX6jyu6o3
xmPBJRPuDlsjQZHHF2G4klXNUqCJOTXdSEAK39slxdQJdncQPDyjol9kNar2Hfqyj7pK0/V6w+yW
O9/ulhjsfMZeGhVpxb12nYdp5pqRvQSrQFSHlABdbs6e5BK96oHDtxhCa0DbZjU48NfQynG8HlF6
wuHpXaMw++QHTr8ZYBg0D/ToDJX/dVtjyITB7r1Tg5MnPFv7moh2lGkCTTvHCM5S4PyCaD2P1dVo
/i9XTipJE4+SRWqqPfn37GZ7Z5lzOgQ95ZuMceHEO+NuT+zRAGIbYHRZ+QtVB0L89cltyCo0hAd+
kLa9mA4Wccz2MpnMOqs8aTc9lrkPhYcz8tZCK+qs9Op46gV1Ek7JC6go7HqOfC8bgoyVI0j4zi9W
l9BSPCNC7vDDG5b74a4EelsRMlMBSYcqsJAOlK4XwMzCZQsuZFxH5XWIjUZqABN+rC82zsj+ZEYA
fhdCK6iojxxRrCwB6w5XW4FTRpxrKJZJl0uhmg5g1t2ULLK7GVi3PTSFRKvK+qtA3jZCS72mga/O
/u2AzFAZSDq9E0muinEOcDjsLgU+XCx8K48rPa+QZT19DoAnaeCtVbb30CkM/XFnm2ob9Rre+XGp
0UnCBmrBL+FFTABRHe4hYsVYqcmBuHFJsQCkraXRZifEevEmccrODIkcjZBO7FtzPGA3l663j4YM
kdfWbCH9VCST86ZWIrYatmS0drg7kbNPK/1Bekgrq96Xg76HstgzMtVDTkWBQXUVdcp+B0X5zcUD
khJPL0bv+9rlf7gtoX5B17EWkafm1o3l3JuOeZQbNxxOmr14uBIf5ERv6bHiVovzmH/KXlp2CJLP
K53avpHWsprI27wAENDEC3yxGQ2FGsFjdZvjlab/XMKY5VWlgWgPS4Ag83zx7k6VWcWuS8K/k1aP
jcdSkfhsyJuZqMDW7TO55OczpDuMEHMbouFfTe+mrG4cV2rXpcHVgTx1IuD2LEv07BhefRr3lguM
mToaL1PPkbbJojey5Xk85j3YdJmqOC94knwblkBKcbrAkcLpQXX8g9xUPOnSxqexnOmts5lSsPPB
LP8DQJGayUtAygRN3e/X2a79b4WAY/FuHn++Ig6JJUTsMHHkyLORqnkjV26KCeyIwgu7nr7cuB58
BUqvgUV0zvRcQVYYKZbn775s4mMbOI93rUiys22MurKjmeRy6pnWId5fRo+0XDSsT7zNgo1y27kC
cd1V18qoqGBl5gh6wrbQwY3KlOC6nPFjCgXDf6R2TsMMXt+rVMjtfv2QUt/H2vXKiet3qxy1nSLT
+WmxP0GvML1FztPgz/JPhbZXngXyDEdwqyxG0ndotG+9fDXZcmY/vb45UOK5lSy8v+fANRBLQCq2
OF3+V9ogh4ooMBnO5DLx75dmVCa7UtECOARZ8I07EaWXUElWmqsgr5RXDcV9Dot+jDQphHHgh+Tq
cO9vjJ+qCow1+oJpUXIBXmPJtyU0lF490KPu7LmTcEMoqv41mLd9qhII+iBTXZ3zZjeRUR9p6F9I
bb0AEEmjfhacBB+HIyTbti6YnqW8LXm5HDDnivmzwjITuA3ek4JxMl3ZLYbBsbFbk3GK/J3l77bj
GWmjYpVOlOoyhFSU/G6roLP8aKqGTXm38KPfxlyccZANidMIoRUcHoIDCIeO8snMdAqjqZk/9vsq
lfaQMim7RZ59K1t0KpLNHarA2ymC51VZ6E4jITjmKXG9ptBoyxg0uGQa2bvyXf5WdBaXZJa+mSph
7JJq18DFxMh7b9VTmYX/CSCoRJbqvnkeQr7qIHOAn4HAl1DNsNm4OB1fL16oTAehjtV++8Omr9tp
ym0e7Do00TTtLwcOgZBqXjWC8gKt35T1dcEBgCp/YU73resS8WxlLPQTpL9lCkGqKX/5CzCfVgUK
nenZm19H4IdGPY89E+rlDmPeEhPcuxKg2+2PG6KN9KDDWFyNBkap01bUf/UB04ENwcK7qR+oxKDf
TjgEvKYlUCQIEvUPY0uyJ9p5ceCM9g09r3IqBGUp1vpDqAev0rQNhuqFoz268FV/t/lISOaDEGA8
vZ4NmyqXoJb6m7rxBQOvnzi42giBR5yOltgXLlKtdSkFWsplwj5Ft9vnHlllD5GQ0iWwVauuQhIO
WnMP2W9PydJa1q4qNxwYq/hx+YnZltU2J91PMwVaynj5VS3Jzl+5FNZyyXHvjS4oMS3ne57VbK8n
BiGHo48fL9lBMmhV+fXHOF91aSYf9A7Nifd0XGVOrOAyUk1Vp5kHoCahrX0fQZHUBhwiLe6I+nO3
ydA5U78BJoPfqoOhYWJ4tHNg/eHRApaljrLJkuoaqoFNLfj5PR7145NzsSfv/efVaBFc6eLj56g2
Qtna+WGHUwHtUMRcquIU2AseJdx6AiLKRSi6M2o4aewX0rzXAuaWhtsK54bNT3pO1Kbb2j1iWner
zPbtd6ISdK1dFEiJeYk3xX35ABeNeLUkavRh+SeIdj06kNJuibyB88DqwPCTPMe1OlYkGxk66LK+
of+WFrWakUy8iIv+27dbLqm17XL7RENCKOQZt/YyzV9RdQ4zUk25wqw9O/ypRH+3Z/F7bAyLmMVI
kfk6bcjIS8NcHLbafBa3RlP5KY9PRDKQadUcpqOW/xOuzxQM1BJlYKyRbp0k6ENB4ftR95YeDzrm
P8BO0dIu6igtEy77yHeUQNd98tbvB25SRzQ+HIsCAhWUQ5eHNkReqvqtpyBFcVdH94uV0AaI9KAC
Bzz8ZBix0X9/BAcUOYodln32cFjcdP7Ko8bKAieg6YZwGfdwGz/SN5BLkNGlTsEI7DRufEihgcFF
lW6yDJ4ADSUu6BC2lO3DxdY8xa/8+S8sbNoHXOWSCgyzP96PVCquTX4XbteUY/LMXf4Ib2rqbA87
tt1fNmpo5KWdinRpV1VZ8mT+t6tqgbzBzN7GMqOGli/wS9VJbyZle94IKyDaF87SwixJG7J7Ixzb
5l0tUrWp7yyV95WkkdSJq4uOR3K0rLhm2hicgbTGaCFU2Ni9qkhSpsXmK0ToKwezOP5+ZlEJ1SSy
bOJj9O1mB8g6KVurz8r69DhSu3Yk/Q9LByGkVrDjiDcxCwMQNuK1QyShVA3J8m+scJ74iDRsAggA
/lLzpTlY4KhB3XT0zKsnwCqX+Ip/xVaLH4G8s6LNx/q8m7xp6Rh1SErzMJ1Ktt2E8B8ROpUteRzj
V1jYEkYOm7B7jN1dKhq5h/KkvyoCvPqaXAOBtkVnUc69Jg8hYNsRwvHKqkxQzyBMfz5ZjCB/YSZy
rImpxLvN59cbmx39TWvXUmdztOHiSZUa4Jc/TDw8kNEUOHD3NvdsQXAw6k8M+ng3OQslnWCoUYNB
EANzO0ae4N/ZDzyJaAVdVdnsxhX1va68+bc9zyWIu1vZnYp1TWIeaWk3p0yCz+UzBvVtOx+LT1xa
UUV0leMH95OXpFNVd/uGH2t7gYQIzCzx5W4IF6nS6rib+QOeIENVAI4z3FztkDLx0WbaCisaiEhH
ISLaT9g4snXYPN3UG1TT9xAVDBPmLhc1bJAPqQ82hVIU6S6ygd0V01VK/8BFb5klLOq6LWafP4NP
s32jiVtct3QtgJ3HkV7MGNXXtmUCGk2v1953nOxkwMx0emcKjjrLu0zggHMynkfFJ7FaKwV+ArBl
9dHaRg5qjhiHtKBmdUjZUe/RaqtNMh9bJpT0auNLaIT+9tPDSP6AJ2kO8T+iaGyuS6g3ZT1sCJnq
mAhlhC67m6Ymz5tT7N52wiNvkTmy6x2fV4mdHCdJqP6Y/2u75jTvhFPs+muheYFPQkgyZ+h0gvcQ
eaFUx6Pgzbl1ffUy3g1GeorLz+izTk4QEZo2+ZzMIPw86FzFWctiD9k4yYR8+0dNCdAuZwcDNuAh
xXxRs7qxGWW2C9ABM79JMwHhqZgmKcAu+EFIyVB1n7l0mgNPWRYwp2jCyAJHdpyBhSkg7lqK0r21
xRWwwDi9MYA6C3ku7qUSTVKKw3c4Fl9aUeeUxaQKbyjsnQPgJ/gkZq0nCKbHCAfemSsQglhFH7kD
ameIgQTW5ionIFJ2C8RP91LttqLJ1BTlTwoTdqIdGKfDDK7eZ2q3Zxtp6YBchhEfR5JOPpbDbCkJ
V0Awwh7MNV8/ljJEjMM6vi9EKlcfGyHpJvf5agj6xAcjB3uq29+/Suy0W69EI2GVtpCdjMWXLPu+
dQTzSa1lSgX+9z78khmIEyN9Hp3swVzjdZK+glb9ndv3ZZn2jNo6BrB96NbZOWy7m5Rq8AQ9b+Un
qhov75L7euI/1K2L/gS7mtB+4ITzQS0JGf2sL9yxnPI1GUwGpQasHebwg1WyFdjigp+VfMJFsRn+
OOfdaXEJexUa8DEmTFZ7vTLI/2YQSno98WJr0pkd/lhcLIDPQsACuyrjgWqrQryztx14OeDHQPaj
a/C40HRfXysyIuhyQmmIlZxoIB31oKkz//JW/9taxMXR+nLrr2+vXSI3nuDKMzVG1iMqd6pP2Vqt
1uUPh/XEmILTmtY0OTZIQ6NvXzSPcROpvU0NiC/xWhs5+CwWFuo/7MsQBjzJo1iwAxZtPTbcvjh/
jh44NSAXELajVCoDIOzpa/MDwZuhCS+eNBw0lXtl62ig3LALWFj5d0PTvSAYwn4GeiTr9VcGBq/3
n7EkjeDpnYf13v/ukP55fbm48nT8plu6SkP9CCKq9X2XU8/yQ43yea9ifBwmGoHjbt9OsWg1lPni
QKr785ul/1OfENMWQ/lEc5m9GmORglctLtfEt1Lm384omfXAl4ajrdKeSCJUGBZdBl/mE7N5t/jN
sOj/umnnEDAg8VSj2/xdMGyy6o37DibW9xURqq3nt3f/p3ohWUZWhw0hlo3l/lWL5ed8Czs8PPR4
dwD9WYFGnat+60gb4UmxIQk/q94l6DJ5tqBCP4bt0vzK1FItpTI0JjhCPYWHojauwhlpvXSgd0fW
BOFoAN0EKC27r9pDuUa9hQR53kPfE77buJAbOyi4t6UUozDJDRfQnhrzxezm/87u+b45zChORaas
qlR4tYkkj7WSJ634LoIM4dgLSLLW7YpVM+uaSkMfhKA9TCNKpS8O8DbTJe0zBVHuSmcdzcKVTxb8
2iaaO84UaHFpUrJ7KO/QxN5MDXAyu1o6zrEmNjcYoPOJh+rZxztH72SGLkitI2akHty+oiFrJd7p
Eks2HOU1ZieUikr1DYIVCw+VUB1HR5lPUTRgSO6zIdzIKKQv77IXvu9QY/WNrDSXkUyqwpnEw9YO
Ws0cIwdH6UXcdg3S9S7bVYgNW17SxX5kQbDfPG7U07ajsASaBK0B3aADoqSXxcal06LMUEsQ+NUJ
eIeGXHSDSrHl7h4PZ6IhpKPw63hhROg63A91z8Ci0TPv9MQd0/N9OKL8YVry3ivyE/TGwhT21aas
2ps57K2xoOIZiTNUhJ1D9Mc5xJRkx0KZHdWm2Kxl2Bg/D/ckZlWd3cHbLsByx/LOMF3Vz76iqlkq
th7dbaozv21CaoMROyJBPlidsHArRsSvtwYY0PPWqiqHzARzbaihuj94lePKEdtrs91ZVl1RxegA
McJWlHvo2HVRjtCeO+b+EPljL11emv++o3FF3D6sJ33zOmdBOk+FLUf1SXIE5FljVBwhZUIroK4k
c/OxspPOxlI1fIxzWmuXyc2VYjDe7F17p3igQ0+lRCMzvGPIm5q/VZ39C+3L5h0Re2CjUjB2MQFq
M0zomxZCwgrOPjADP2qYbgpcH4q9Ztjqp3DZn2ntphcfT7MfKvgq0IYw4e3pJbYvrohqlO+qDyr9
31oUK1qI/h0R8/i5qafTN0XAmGBYKzkxu8kRWLabxG78KmByeFmIY/DwmlyvtCLrBX02Wco1DBgY
PGc8LDuMg+oJL0VuNc6DSpqA14MWfzlebb5Wfhz1dIbVYOmJuQpm08yHUyCI39ZvBqKNZOqcYuTZ
RVD+n7NtpnpPkX4Z1GBOvu9gF6ukAUPBj5zGsLil+meiNXkKinCmT96eE8nkvNM9aKRhBQvzDoME
KhvD+1051E3zwQmuxSiIldKTUzg/Urf2OV/9YthkY66bCWR8Yjsofr/wgx0Rya5PVEwZKxL3sYwZ
2cbRIwhxgDxD3bDNk14SmZd3jjbACb39nDecb3oLlHLRCGu8oRI6G2cyKbnf4j4MU6lNwSrPqO6+
ht4fCWMYuOqhNW9GRL8+/oDuwqfhq4WgU3GGgBgxdHb9ogqmIjZIDqbEBS04yVa7YlCRb/8aM2Sx
EqDGGaDeSAxFMt9I/+E7LNl1UZwvuN0KtsfLNWRiFLfzF8yo1ZuAYlzImJCAPr5QZAk9bMVTrQwE
4yoLaBIjxT8EMclqg6alJH8MNHwO0t2L79ECCeZlKqoPPvlnKwwwbfxNt42WdXaqwZcOPW2A+iAe
tJk+vYDjCynCUr/eGlxm64dV3m3/R9P7iJnV0If3KgsxAVdcLoxep1hGC21wZJWCZtiqZSkNbX1Q
hO/RX8bD21pzc55KDXY4yP3BK051zVh4rDVN1bJqdydOyHgYuAM/PBnusqBZrbKsJhWwDepX2yyi
Ff5P2NteoYFyHgWqRtCE/MeJoJdYl6ogYS2g7TD+bB2H5UPGx3wwU4e+5swU440TIOSOay2OvIdr
VP7yAZGtWVt3o+OCDZlpN+KkSqrbnATM9SVcpZ0/1jR/dLhwGi4dz+3xCEkaRlMtZmhc6Qa4WhJY
0ezLPMLTBNE86lEJiyEf4t6Z4vg2aUvFDEGFB5AWbcTXoPBNl/9Cg7gvUw7z0X8XCWgdyJcLcmfz
5N7K3WrKmj6qgyHY3EeMZQcp9wxXnQck7MetYy58bUmek2v6m9RNcaB/Brx9bwZy9Zs5t09CkKqN
QT89AZ78JmLQ0NVKf66QRjaJSP+EgI0vZcXsRvwl2LQ7TB0HtgFSRT199777wCkX26p9zZheFVW8
VeYoleoyMNnQ7K9EpXV0a3/6sq3+1dYz65sz0DcqEcOLonHFufddRRwPAdJvy4CrycY8Xz7WISgh
bFiJEclOpvk0J3LusVUYMd/5saXDe3QE+BjG2h7jJKmwuJnyXbLh+YkrCDPcvshIHDmEFM1SE6Nl
t9HImgpyg4Vn0qujONNiJEI8qUS5pViRU0m6NycClMWhfuXVTEv7/yiGh+B4bVJbKixdGmA2h5b/
vqzVrVbMD/SucWIKKkIGq8hqxRptMfJJ+LvAvjOWtuuK1e5WR3DQqOd9/+hMDadRhAnXGb/8K7Zx
d9SNGni++67U3Tct+TkU0apTj5zgvTT+KDnYsLhrugGjJYcWg7qK39DTHJruXT/8++ENPpSuo8w/
GuIJfNosRvxwamlYf51eLrq40PLNVYStqqVUoIquCwtJUxfh2HADmfgLm1L8lnV1kkoULC6cIogD
WPqFbzlv8quo/Ynp+D2aV0w+e/O9i/cW2TI1d8moi/yJtqRw8A9Tvy/bmoZuiu3BzWgm+cQMSRHT
j+R+cxsflMJcn8fxuangX3RYsvMp7mY0xvfvJPAcT28KZwm4sol4kjzXewIV7YiUAQ7MGCFWy3Fe
h/fycJCryDEEiTCLI6LOfXO7uKHC6J5Eg7lxUqTBBvn6EuiM44qSDz7AngtVlhPeKS3X9ZIcci1u
Sh3/Ro9FipFSuFXifk2jNFVjmm+7YPrJkRDfpkKg0cP4144AlJLrxo3biVAJv2b69GZxkgRec/kr
fvxYcFJCftfhgxOYvQRkgRalJ7jDv6VG8TzNUsHvgx5z8itYsLaCCuMrYlTAqafzs7QlrLhqgA8Q
buYCNkMF9iT3fAeU3xodD1XKAFGDBIgJqblWV6pIbPIYovvZonlMOi3OPJxSfXaG5r23l4e/Cy9K
/srPiTWFXzWFqq2m3TApF6RinrAhMP+pwt1fUGZdDnFV6pYeLefaLrk4N8fvVjawQT7LfosHqowY
bU85kEn9RAb+mYqEhmWg2NTM6np1khl3SkRrnnPp6vfoaPTqCy4gvoqvvjqGZoGWv2IzQUvur6kb
rw6y13T3unxXkPEX4G8b5yNuXcZSPsYTRvuhtc/IpV9NZcT0edbiIeHso44k4d82hJn6yonH85W8
GE7r6w+HnNYvdXqw/kNktBp5w0LLZE/WqLh/AtIBq8rX6Jl/Fs6fKrVuibJF2eSG2fnkjOzb36kf
XMuHEpUaTmACESx7Pt6OClCZJr6NQjiiMxDwT+mMRdBHUbIeDxgseXX6zfDIA4azyOX76bk0Krx2
H94xF+pCULLzJMEJ/EF/e7YOV1O74pe8XEzzYmZtmKG2Ix5qv3vdZ06QCYJqadScsdFME6apm15x
YN71me/BKAt5gxiz0p2SeodUiw9hN9xvhD28vdC3kRHiOq9PgvmZ2EY5ajfn+fxxZUKvM+ctF0Ez
owjOPNfkd7KHmaTGaWMYGdmf8imLodp+7c0rt1xMg0NtYk0qB9nqgG29dF00QSS6uN9733MRWTYM
RfMLSiuywMjKG9cJwNrji0GNV4r3WvD1J1D/+3rw8JywoaCeOtw+7vrDXOX0dFWbH2PbpmIF90Do
fbYwUroL1Q3dt8SgKuxim1qMTo6zIs91v6XluWpKYumAVVMpgndzmxZBG81bKhiTuSmj5OIlFEOk
9GFcvM24UaTqODzK1IKXU3T7JkjQmNhEEvCxgxtIERFnhLtUuIVbb8ofTix3olaX65aekFeha+cP
QyoYqDGQRNIyvJfaARJSIq1KItETwmoUWzE9flV2A4yNW6sBziUWMAoSD+ufWaCSCkMDu6pwJFFt
eYe3t5xwGc25V6kLC9xTHEqKTSQvJhhcdCkvg59JQgF6AwnsFdUyjwtWLTfIjDfcKTB7nMAfzCOJ
Z3aj6xyM1lkGLlwqrcdO6cz22QN98JmNzZPAL7Vt7hbvvaoWFmzGNESyzWXWxDIbzL+BdwVxItTK
DvzzF0Oo1xYmNrdERXm4v4lFkMmDSKixiVjoOGe5tsbWhtKd2vuri7oCYkpsaJusnFa8pE1bkxEj
RY6hAOq7TSnFH6lWzki2aVtdpGnqaWChp/XWK3eJtHoRWwM+lcBv39hEmP4iPbFCx/wgpcH36+T9
xHqNUGZykd88MWl+/NI7WROONnAHg4WKRMZtLmFCML13EojfmAzFx/Hs799K0q84NOVqd3VJIRXi
ZMVfbKbe5V/SVXOk5CZWXxGtI/nDvVTX5ivWYbp8llsFVPhh53YdxIqMvoJJWuLTYQx4oNm6NrGn
OJRbvVTpro3bsTnsAYSetDLVMx+8/2uyRQiga045S7UmvZhhELBaabHf8N3YyCFCY11CnfM+lr0c
7GN1I26j/K4hzn07I18skrGs/v+jrWrK4Ln0HC2ihqBP78IK8zYP9IeFaXCW3euc5KRP3yNm7IYx
jwSoFc3DV3BvzAZ1fyNe6cnz0Bko2vMYx9UAyDCQD7er7J9o51kMjgBsqJdfjYWPO0maBNHUsf6g
nyBEjUMQzr8va4QxY5A9O2AiJ0VHIhHU3rKwxOCdpXlMrMVHShAeYXrObTUi/4htSdUSvE7xpjji
1viX9PAOODokcPNkckBfi8wU/8CJvsFJ66DN9Xow
`protect end_protected

