

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WH/1Hfau3yp/7ANrlzYJ6lp+xOi/gEnoXSHu7RquVCgxmSwM+u6NJ87pS5P1rM1REfM6bC/4VD/K
djLzpKr9YQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K9OQ7UQRJNNsqlJeKiLZja2cTpdn/7D08GuVLJ2Q7YwPyOa9sKS+3g/15LJ/yRa/zU+A98tod3ce
QlWEn4ue+HTvQflEH+MpavwOpNzd9uaRdRTecGrueadi0jZCWhKDECPBSOBftTcItmWjS+iuOrYA
UzNSV6gBgTESSUMmlbA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rfuGizF/z8gCeFD2+mr9MbjRWuTPDiFayAy9W9SH59KTv32ja3WRqyFVDNKefGFWmFgyXwscsdSc
S/STQk2WVtfaxUn47IIZV3HVYpgEROzZ8tdQyrDPMbi2HwmCfaz6YD5xdrfG9Tlx4ToidJJ8M9l4
XJdd32TWh7NYEzLxqVy6SlnR9JfF+0+Nf5C57mxaFcf8i5qJ+wGXhxEFyHFj5aPx81iijRBXdTZB
X7F/NtLKVCgLQvWL22LQZOJhyZVP7Cypy5OtaouwesfLnz7akydXxvJf1kqXrAdSNY4YWjxfZQKZ
dY2m3KiIO6F542kNq0ktevUOXRqWTgZJhPauRA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IUtntTnFOD14laEXhqBklNwiMVlWXctApP9259AAx8PFHjFAnJ8PvitVWk2w4ALBNs1tWO3QG+lc
7ANJMKcNRDw3DKgO31xMYxIed+W9fGmJO2Vhw+W2lfZUNPYCZDcGN5zCsW0hJkR6oPg9+0a7K7Sg
VTgdoWPi0vZlEf9gd0Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NobNPEAvOyayp1TtUWqLiTt1wnKf7VjSBi0esOl6kg2wXxaycO7UdL9j1KzK6yLaXpPqGWArWcdZ
OHZWjNgANQMvd87WyNjFR+DZMXSGqH3lTJ+rUOlsySu0gV6nE+CIBmIaadzXmtjlUXyV/oEoRCZr
rq22ZdRXEi/z57ExJp2QenIf48qX0mmYi5gFLdknqEc/38ewzEWm4uHsakTPzO6DKZ89VmneHDI0
7Rw0KBtgnhcNeggKkHBNrVAExbuEzB7b9xOHs8SicGFL9UTrJpF8NFV5zuKj6z6MHtvPDvJ2GC1W
BJO4/x680qEH+0G3sdhClIkA5Ln0j075tcfv5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73072)
`protect data_block
yU1Cp6t5dxdvoDnK2tlp6gUVS0KnwXtsD9jYNTWrkboG5eTWH3fbfVJpsR9oXLJ59//BquaYQ+EY
ekMzWImBOR/sQJhVqTtEMHUI0ii0ob44/oj9uVXyjyo7DKvOke3obrBqu9NDFG9N3N/vlE29oexT
3yoviJfGxITgeh3o2QAbrsjiYTnh0xwrfmWUlpzfeQB5C63AzCgdYP6bJrfxp76qGSSV03SeQnuW
KoutuWND5chw9if9BS7U/g3QTVsf0LzLXNBVTt1FTib4jbC8cPdsl5lBhO1Vuj+3tYYBqk+OGDSR
5+ekGtRFk1N/p9ao5RP4UzL6bGqeDb138aio4arQMZNRhYdWEmE91jXD1XjAzerBIneI6oFyA2Rb
zVVP1V4PNVliu0kR+Q8z+FbwiNJLxVFhQ2pMeMIBD1mDm96aEq/dLMpIuc31fqr0ZUdLmpmMNkjU
EXUDyvgii8wBBj8ZXoF+I9CVNyTASYLC80CUhVmhM6h2V/x2jp7JPOPkdJ6VZdwErcO21R42Et4g
vtKEnvACuYGkUS+GtnCecHGtSH44cmqQBoqA2pfqUpn+N+tDAG2Ec3eo/vovMDaCp/EWZC9VVLr1
z4Wj+sXjQ4//3dCdP1yLWtwrlUqFCvmdKTFTQ8vw67OcLHwAdda3bM5St/6SdchbRuEnMykF1c3Q
oN4tta8oH0q/efbkx97lKltwv+L/4BKDLL8OR8raZh0vxkVsOKUpjq9TPs26k+xoDcKYsCo+L5oD
u0kObupp7p+eDpxX4KmybJN2uGId6i/JHqqPDBzdIm0FV5mDuDSSs7EVKK5gQeZ61V0+rD+OfQyu
iqvN+tjpqj4xPfSoRL9Vy81YsALTTxv1+O1oJ6Cxw/ua6nK2Cg/qcJMKu0mYzp+DbvqOvAEJADzq
x0+PL8LUntvHon283W8BqhmdU8iOovBMTHnP2on71aumQGRjjRY54Du47YJrP/ptJyQxBfWZXMaU
zn2qQIM871FmEadWgF+ZuBKL+beZkyhJqGQ1TyRJNMBRIp1n0IfAyTqRaX6aCQI7T1cbdb8ZewzX
WuorPAVto3cGt64bSxKhY62SZK6fhx7SC17G1ZVmncsIG4+aINmqVKSxaKb0L7aO3fVsElTpuRLX
rQQOcXJi76IxN7RBG+thGLLflPgPvunyHcGtvhk/XL1zrk2gNEPIC+oqSXtZ7WjUCygDwa7+rpmG
vpJ4sDHw2Kcy1Okp0nFUXP7xdUxGCITsPEP/wLNlKZmBVTQF9A4/TEhdmrEZQfrpzVZ2HIQr1hAu
+kOYXiWu406ZkkBkk2/sDj9DysIO9nE2L8sArxsZ6BDZo/LcaIqQViAyvesKQ7gMLStzujxq6UEo
nAWchALX3i/txMCom+5RILvWJPvLg8Ahfo4dZpQmZTOPDqh7usSRe7mDekS+Rk6pZyu61T7uu3QQ
9PyPeEVsJBuAE/Qo40Fj8jlEGe0Z0N8YxKliknYnnfSYFQ7F6q3VNIOUXHj/XDi1DxzzN7f0r1f4
HclvO2+ZICv+UgBWnjSDnhogr4iON6jFheNo94veXi8K0x+HEhiXlIz1AzgPNKDKCYldjMkAiC94
u+ysqwauqcGQVjrn0MivdgRp+Vsi6SNUAhNQiKD8CWg38F7j2LfXmsm86Mn6qRI/Mg4/5XyzSdJ7
QyyiPRhYQtO3DBaw8HJ+k/bYiXig0dPahMzUKLLbxtfPvaGdJXbce1FRMXQ5P8j+NskJvM1P9mnn
iZ4W6iWg3ABk3tu8wrtQOCV3/r886TPPEpAcSmnItUNHiLWG6kqhGdeasKDtGuk+aAQFqTdHSnog
BZnO9E0Lu4dm0paeOeSTvP0OXahNzHHd6fVq/UDIrWZr35CedFCdr/29XTR/PD5njzkcFqDYL9Ax
mQfXz1uu24FqtPTpN2ILSTywkWotO38+a0L3NBaK1xNewUI6wVtZ0s10W5QNKCGGkFZ+D6fmm63a
2GjwPuB58STFcWhnQkHKJH0PlXDQF0jT0YK2wSwiwNnpbnDoSRSrHaJXzK3t4wOCAYYAAdggkfas
HqaXofaUo3tdx7mtMSugyWatOk3d8DZezXdCC95gORTFfmNx+RyKJrsfvKGoPrYzRtzH56gtdX6W
ciy/bbXXOvY8UeWFJFjD3o/8XFizsNpNuDlz5xl5z3K0hOZ4JWxuKzrfaEtNZloRZyVjIqwCX2Dn
inNBc+UC4ujRIjLPPTka1ECPkBLHPeJRMm1Wanyqh42adQw4tQOBdJAHB0JHeNtWIVSiECVkzuNT
ywVBPv5Ym1Txr3qpgaKErW+9wwRFPonQkxC/WqMU4F28LapAqaukhFr4DxJ5oD0wcQCESTQlJLHX
HV4fCAjePF5Xmoe2FlhpJ+Xzpx9GRng+ojoMcE7QGblmGdQL9ga1Q+Y0saumgAZJ21z+OCt+DErQ
QixWLFf0jyYsEgkJJ9BR3dEi74EGLGI+prgOR8+gMzeUpZ4NMvT/ugwD7ULbkdLQustQWAZufl9R
Il9pMaQb54B8B95llgJwxmbLnvU+VQIuRXA2AcY+Pw7v1ajh5Hy8p/dwNsFrwe1mbkKRmyD7etjz
PCXXgGBXPEe6QpyJc9pG2/72vKE9yZlaxVCaI8c6rRDGZjKBMMH61NYMaXhDA3nMbacLiFfnA26G
rDgIj4GDGmligZIBP7ms0U6fZ57ud7xexQknwI7rAiN1GpGYwuKLAgp0PXzBnpDSDYY5sgnAUSmG
k6P5hCPjXb2z/gHPqH2KpNnsq2IvbttuZPHpZLKWXbvm9ZcPq+L71z+IOFFagFQzTqHTlGbCPUiS
2xNtKPQdK1hOxdgZZyFuU+6oerjTqZRaefeFnUs4ERtN/kvLbL1Cqw6Niqn6DV54Yn0g5D/v8y91
sNYJLAmQb+zV0R9jShsnVn/318TwpttL/1C41XNrVgZRecH95FJ+c5awUIUUJ9ysLi4JJvmep3is
+eQQVN/RTHv1Hkj5ncWpMoRCP12dbw1uaEgW9T0Iz2f2Zbe3rskrn/5Bz1uif/gK7vY4x4hSPJfm
IgzR/Pn136LOVrfFJdkWNB1AUCuN/JmE9KtHR+TU68eOOOAw4T3SUxrVYEjcQvqaHK4LDt1zgafh
/m7gbTPXkO/eH4sFxNlwebIACLltP0BLXcuD5CcFgZ1HR/S2E88uFLViAI+yJDmrc5GFzJkyDELj
MdJHszFMfUe4p1vT5jPfYUgONWOFmDkmwddTqw5myCbe5MzcLIgVjQByP55XUTyTvirkVKWQUPCY
5EY334O9VkJCoqE4uruu/g0FJSQc+d0tuce5inY1L3uaugLpyxCfZlng+GrjL6Z3y4/zCmBCENJy
oDsK9IYm7lWsxoYWCN0mxGXw/CoSy8QrBGXDUSECvR3znTpyEKi4421rrN9vK/AsgXd5NKuKdJlh
IFY60Xai/nDOZHOvy+KuTV5rena0krB8fX+nVPca77uJ7ze3lERt/ZPULql5nVOtnxnOD95qnSVs
XIKqmKhbz9yiRrXZXTx0q0+t0/m5UrDuv3kPkrPVEAvNae6RVlwltRQzNOVhuhFWcambC7rdtUyd
HPTld9pBgJeTUJO6L8Lx7fZ6oxvhNu5Twj79kdhs44xlSf5Jz3bqxRNAVvqlzgplBG20UVABl73n
AsJe5VbqBSOyml3HV7/meTgnJ4iOpV7R1qq98cSwvimhDgld8TZK4X/j9817smy8Ags1a11cnE1f
qaMFX09RhguzlF6kML1Y6fufGxYkBQfka73iskocYSF7AKeCTPC0Q79OHkPec3bSiHih3duZB7Pc
1gUaRLPjSOvxgZHQJq0Gcio3pKQaZQh0emIgLCdwpNKQ15FPS38IIBx9FLTs8Zz1TXU1l7Yu8WI/
Q5WYn4lZgLAAPg0IA5w3jN/uTfrXowaI+IdBA5+YtO29JDEjFkRgbIWn1lyy4SwK2wHU+tseXQOv
9pG1d/lgBEYwmNSBKww9eZgFP34RQchLewBqXkmm80QDjdIIafjmU9alxIXve1qC81DtbWCT41u6
Fm6hwxONwxUbtMjDU6JlfurPyFx+4DWr3qz9+aOQ9cca/bUVdJaTmvvWI5f+l1y9IIopsiO+6i5S
HXrgpHnzE7xhTDo/7AUDJxRBZLID8ncpfikj8iyLndgM78OBOEHI8xN85XOzZI3LzWVnxvoMO6Fq
WoFYN6j2oh86tL2QYBbnIrAw8RmG3+YVdEAWUCNegyf5Pch5FtsFltA7pECuGz+7v8Varogrv9sB
u+qT6G6/7WSjB/Esb6avB0r8v7I502PMyrZEolfRLymH58aCGedDOQReXSKy+8Ek3bbqUaD0rJoh
TPi6VNB+x6yvjGCQTAChtInpVVuruiKeR3xnd+jZQXgdHgERbbTSg4ck8PPFm+62REi9aqkvGRLZ
v7SNoLcJ1yGkVNwgBHNNdlX+dc+BciDGUbgkD4x9i0rbBNDV8Rmwb9Ya1e1N0fu5QxtPT9ZktFSe
neGRhJGrDxm8OZs3McYJdIo3BR12twemkaokXkKoC0xpGdmhd4tc7u1+1o3hiXORNEiYDEMnOfR0
c+96unLRCokKrE+H/4aiYlmD8eoM446YW63OT+t/xbhcM4jukzrDt+oXTT1evPBCUquYx/G65Z7r
4YWKhY1Y9JmGa1DwsgN2g4NsXFkos9JhwSn+M5/QeokWJK6e0j2pH4RdKC/Boe5RCwVGQ1uA7MIY
zcPYBTziuxNjmi9AgJaFYOZfYmv4TeT5cSBVP47+Bs1ejt+kJ5R61wsck7/4kIHrpIS8ORPeB3dn
HxvDnxPmf9dncQqIh5u506M9EeV6mU0GseWMw02CwbU8q4/Us6xjwuC8nYGcnq+nU6ldZXuXysqx
2lOjWdG37XgAODA+wNT8+Cd5Gy1A+fuDUg1d109B4qnC7fCgvXgArdU8G7T7+3CijpZN8wA70m2I
e5YhkyXJfjZMNXUgn0K/7IVwODZon8deZ0MFZPXs3NHxK2GiC3U7IzMO7sOsJJYH923Tfe/5hhFc
oSqWDDcMOqN9zrwB1PrcT1TCEm89BLXxTHTbttcHd1JjV4SG1f9n7vaWBHWFGWNtEXY7+IRHiHDy
IjljPDrVZz4JTBZQwY06rvHbPbj6f8pv0LjIsQn7RXzUgXfGEG4CS3lGNyHEd+SPG7PACRUfJVl1
RWHCzMlgDuvmfI1F29+M+9YmuzbXJxGPsaYBkxk5Y+TsjSZiJht/WiQ76/LUvn5mJeLP571u019i
8WiE4guaYpYsm9agCxliTy6qnB23i9gWvLSkA7rcsl8FbV8HSFwCWi/QoYp8uxTG+Hi4lhlMFrPf
0lZLUw/1TxupvfuRrO8OSoAGuZxiqTSWDeK6PF6D420DBKydaiafUT1rotUmpDoK3JwWJu1XPSpA
sUkrf+wPYUrXyxaW1xAOw+Ou7B4TLyfZS9tB5I8dUJoNQaK0ZXE4KbXDH5zvD2VNunic/3pZnpUC
+kXxUxG5VLycLpXAlZxjb6COeV3swgg4phPMFDrtGYzVyNXRxYrJpu5K/Ady0CtradMftcSxIuc0
VYjavAPGOdcdYQLTkuV243XJ/tXLu+bf4Z40roXPO41b4YMjm2YFxDhkPSv3l49hMkobWEa6N1ob
7n9bMiN7oP7zVHKDZRKp0K0ZwQlICfCVaZJjVkPw9wvV2Kz6ZQf9myh44P1JOc8Tgc1eYC/iYo6Q
HaGXmqaBSYarSZTTpezjg1RgyVSygm0x6ewt9Y8mKkNBY4g5EzBfeluLRGICpSxrRUG+A0630RYf
S5UAS7hBj/eUPOF3IDevCnmk2SdykWups7oakuJrlaKshlhFt2hZ/Lic8ZbKzBjstrtyHJ6IfOla
HVjl+JWRyh0fIA2hFGfnZk6xgctxWDeYmfwkLLG3rxAkqKgccOlSLrzZpGqRTfka/cWGlY8DYD/n
CMC48ws1tEQqD7CgWi+GjlHzN+b5Mzw7g/eun3b3NKhsB903vQjCpFLtBIa718SnGSa9SYP7LB5X
CvPM+7gtOOlEcCtJYxFgHj3S+PwLiAv95mfKwPJzh5rwvqVL1ltLUVovLr7azG1mi0Ap8v2grDZL
120g7OWs5Rt/ZS0N1eii3KABvFLi/gPJA9gpK2UrH2zGZml5BDt5nqCIRWHiUCKJTq1difzVn+U1
5l6QLJ5w0n4wsD4qipW7eKAE6/KtN4hYWbqdPDNU4DhSgBadSPRZumRE945Vf9y1CWbL4+0Kp8nM
uj+GbnKf6ItBgHeUkJCU/bgnw89oG69zBXN6Oe0DTvyXOBTLpNt5QIWSzVPBouJH546iyo2V+2Vd
iGb4mUUj78qPFSCB92R6o+69+B34O/EGdiO23LQQ4cpoTgJmPx7YRd47lBxshHefwX/Bt9OQkru2
/QxBawH+K/1mNfA7siEXk80gyK9RoAhJ7Ay6pF212XFcfQa4mI7WEvn9FHKbiZP49UGi0jrDTL7U
QuSSy/9Vx+qLwbtYv1q85d3yGqSzQW1DP6tkFAP3LuPt778lICbJwT9e6fCpc5tKT5BZaNTwkv2x
nGI808jLTFA5SE8UnHtfwH9GGIZFNYTFUc5jTe6gndSzu9SFumD9WcrhhwQC6/oqX5SSmQ7DyJKT
wSX5Ykz7n3FX2xu10iukLwu0TQGtc1W9h4PHJfFqRlJQNljXk36fEf7dJPiB/EM8MjkIW+P/kViW
EVLad7Y8CvGOkwEg1zPBtu7X5uzGjaE3jRtNC1NXhX0Uw3tB8HC33PD6XqZYudwEc2y6VC8X4FcT
8peFQAiXeZSVbHqifnc+KLzEKTVk+dFhNzJAPLmjGPRNJFUl9xPc1k8tnUgmbfB2vL38tvibL3z6
PpFHWCmRTNwFSww9jikiJka/u3gKioBXMi5HRpU/hy0ElP04eBMK7nSyuWq9aPisbyx6l9jzpYJf
hPNzhIW64cef5bBjMlvRoBo03yV8BJH6TR1ysjjemcmI1Isqzga97p7ZzXgGxcDUocfUbBz/n4gU
nsfZva/DC52QOMBLMZVgpzbDqOziV7uxkzOfVrRULhqkZF3huGt2iuq7itpYp9mZV8vX6F1ufhjA
QI0zZc2OId90Cekv63JtRv8Yn0zz3K4WQ2cLNk9Xe1rzSVMLdiNwI9lCjFFLiGzFJpmYApHsqgKn
An6XwailLyBhHhcTnZCxSn0diwTQQAe1NbmDTQ7Nb/6lYAcYnH3CfzQRoZuH8Fzu4QOpIM8hb+wJ
uMoRlvHb9Nb/c0Nt0kqr/j9P6J8DSMVjsB8IAEyk9/W4uP/mymjBzl1aIkTWplM0m7c/DDyHordc
TZDhVwenP6BcrPb9pEGPvNuiKjOCicHMRgWyc31Qo+EYGcZ7KxAQv+gmm4gDkv+cu83Fu6iy7YfF
QN4w76cd9lmDmDy4QMNI4cVl4wszPMjI3/TX2rnuKnS1bCoLQVTOTI5T27g+pA2q1D7afn8XM7VI
XMSGsgb/VSRQFC1w3a4h+JSUEwuy+myPZogPO7MVAKnUx/M+rWBaMowVDvLhLJciF5lsXE8lQi39
A4F1ESq5pMeQebQDLiYBKhiG8BClvxTvbLXXgG4vwENfhzyeiu/fmLSRLzZ5rH5jSkmUrKG1/hVD
Fz/B8f7FCFxIgWFp41sVEIRfZkymT3Cukc7N6J2kor7sXMKVI6d0pdPDDY4Xa//tZh7gfyfl5y7h
JlICz9Yt1djOP4zvxBQHO+IsB7UcW09GV3plE75DubeBcY6VrWi+YdMDWNvPwsYNtbdAeZBg3RPX
3HszGQM+BLi6xaskB7+mylbhQiTSiONW+u7xwLbkfoLGG1K3/sj5aKYyqCWY6R2vJsdiSNtj+TwC
dCuNBRgDQ7Y6sE43CLiEEePGbvbpuAqOKyQIlhYIUJCb0BWp/2B38gvAb6kFvoCp/x3n2uRjABJO
W+t4GhzrhVvWYRVx8QytSH1F9OBMDmjE7K1sgUQtHEfoYSi/HgrAIJ21nUuyP9M1G1GH5o2vAh+a
RnnNaf/Lhhsw2ZAatYjCajSjc1CBR2wUnnM9ubFPxWrd2XiriEE3aa/cH93hp+f1I3q16gDCBdye
VltQoIgbeq1GCNdyVJNvNoCyEyJmOlwzpIjfhCQ4lillOb8SYGQkFALNhkdbDLP9nV1wIDjNYJFV
tIzwFtU6AbuY972aEXLuhUA0I4kzzria+d/9PBPtaMPqj1k5617tF/cj6aawpUsyGJ5l37zL6wSy
MRbyzqu9FWbPb73UOBfb+oJxuxMtsrNMV4lGkexB2nvNEnEmyMB8nIHWv2zLafmSDSgy6lf8cCTG
dKj8XwHRwG6zX04AGbymdzR97fcPKsgsBEslVyXrijJRQ2sJwU6TptVIiNhRrOXW5nRu0ODn1TD6
7sNtoYTKj33aUu+t+U9m7gD6k2LZnNTayCfuuepuT25IHri8wvxc5fsAhesXSNRQCv7HBBvmOeud
q81R2fZ2t0TdBRYcVtDn+kEfIfpGCcIACgxlR92NazqKx/KlPz4jYbouf7vfIiCDZYKiS6seJ0Ba
MG2fXY3FeR7/rHDuo4/t/US4rXwWhfCIpQeCRYf2rw4Wh4CQm9s9ceauhzJV/mPkbe1banzm10bW
7UvPmKSUavTRtV4y/2Nev3ulewTdomhek8H9yXhWwAESOLz5V19YokPd04SYtZRt27HXTXyHLBYh
aPJTjtu2FICexM9lmLL+9Ci3wtd9t/S7NAsBmyvltrzOJ6sprkCOoCAe37lBSAdK83j6AKo1HHQK
tkxbIAHTOZtImuywELLbliVlPfkfhUQRubSZGM9zDRKYnushb4DvhG1FowXae6QU8HTNeR8l7436
jzf1rxbpZun+tc+Z62N9RPbYJzyHVEraQa9tVy4tNg/VXcSLghVsbj5GT3+dhwjKtQ42aeeLIXX1
cAJes4pdQbjMNhbjVmxY2mU4LjDlVLIK14bQh3tJ9SIJsUDzIrnxOLBdaeM5ltSSFUFPc0o/QEGz
naIE33rVYHC0OxEjwFHIvcTVMv3bFF5bgMQzxxrpcI66qTglU2VubQJH9WQZqY+tenOuBKIl+lwL
jZ16bs8iij+Pe2yA1XaqBlSsQBDoRwP/KrA0PwwRrdtft1SiTwyBIZhtFIFVWgLBhcKX5V0ySf3D
MtefGA11PKnaW6Yx+SzqfwRF494ejNZ3IyjZ40t8TSvDNsRXLjr9AEApGd0gPHV44jF9wEksejhW
/WCVpZsaApqgHzcDMOb642LlnR5i5Zul7O3EtoGu5lbbh7VDFmHsQk/VCXvhoS/oKyw2v2AAKYZi
l9IVANF3agL6Ij4tAxdLsGFp/4H4mTo/JRXf48SJpftLtnZ5ayMyWC8VscX7jNSEhG+omkRh4Xov
Oryblckc12DGCEkeRcEdHQ3DPqO4CAtrAku+vbBuSXXYS+V22QTbdpEz86Yk7zG3sen09TJjUNyE
dYZ1JBkFAooAuRuQizdeGjEh4Kuzdu1+pvaao+jzVfxQslifCiWwiyHyMMRgyI0SXjN6fgxhPIuC
Jk4hPm04fXCNNuulx6MCum4gr5OrJNsEqWVL6rvqHELn/DbbSJ7AIfmLVBUm2JNNn1rCE/b84nk9
hPwOmj6bdem7YFSJNxsGRe53cK7uxG/5QPUxq+oVvYsjnFRwsd3pMy/P75g3qobn06cphk2Hc61S
15sTC7WCYTY/pomXJdFx21Qfl/TC5Xez6SUWOV0noWTm7tzyoXDkHK1P3xl5hAouKhIQMy3hJqi6
S1tycNu/A9xy3HcVQlzVaBSg1xJOq/LIm/vjSkZgWM+F8ItXDTpq9tc4yK4bsuXmNDbjujjol/xj
llln8mv2Jzy3xWAY35RVgrAVZGuvVRjLfy54IjNGHNozQkIj4KSwQHF9cbg9pOF7HlmmxXeCD2FM
MoLOo0ntgpYQwH8PEvRR0MZuHt+VwdhoL7Oj/nruL1tqTXud7QP91KWODFvFgSjTYdJ+cbL4C9x3
NYuAS5srZ5GpaPcVfKG38l1NbFIBOojK47RR5rbAgOFVuQ2VI74NBT7KC5s6wzyYdERWY/Lggc4M
+UXqbhE3oHOtNDx9wtvCdJmlWjOic5AYKo5aZE8QJg4MkIf5ZiwTc0zquj6vrcHe31C9ngfEQ85O
yd9eT8DxP+2ofDZba1qyMYoQuvERdNV4H/xyBNz+N3Cq2T88dCMqdMDD3xjLYLMpgEH4FL6ih+X9
Y6RAWOaqmNst9VRhubg89CF6AOy++ds95MM4B1ecpKowN7RnvnprX8ROBZCJoXNffy6bChc3+SR+
TQdK8Masu5NjcAx5gLEmiNxE3mSzK0tmSNJnic0tDTaJn+N5f/Rm8t3sweThzczucuQWCiNTyWw8
Vq5tOF6jq7I4FPZu6iy/przBygyLFcLoLkvjLburk9fDnpj2cbHNXt+iKOzN2+4LB7KehD/9UXUZ
sRk4vVcsR/+L47MGZXW1P1wWrM/mM7vc5F5xL7yLwo3F000ChpjTbWhXAOsofbmD/zrpDqaXAniK
zDer+o83AgTuVS7wNxEsh3DNQWKhLWf9qsDD96oq9DGIoXS3ItD2vu/7lFh7xSAuZESIE98HiLAc
r8PzdhlY0mnCuSWYY4dPvF8ng6rG9JZjUD8nsXM5HYtcu4Y+G+YFkrHXH2U9JUIysJBls/uvsLBC
ajJj0g0/G8gepwYNiNfbFUE4fgxAe8LJk5ldnCQLVryMjoRtUYUHl6wx+TPI/aPq3JnNjXkIKBTH
gDc7/vxqbs7eo76hB/XXVzfIQLrmk2fweHjyPQRS/u+RZZflp7T7ZJ708vFKf1jHCke0f9fEdW0g
AIHiZdUnVSxw3+6JSS19ISX9WO/TvOfMkug94bn6EQFHyYLO1j5X4PNs8E4qxHfqnVwc4nAt/eX4
1tE+lGBGgRydTJcRzuIUq4qHyvQCWLTIPNydVpg3mwxYdJ4jk/6Sz4ya4KfcQx4fn9z2orgEem8C
8hXRieZdziMIklR7JXTdrde7GBpVCVV7WwIFNWZbfNkMCWLQdWuL1yrd+1J3pF/VD/5xJLQHsxwQ
CCQHghWIrIF6El5OZ8H2dne28stdBforRGzE2OF8jRDDtQPDkla/xDLs18qXcuMrY1r3cXtV5HJf
kg68BziW+CNRxmtqiOBBkEYSnlXlqNr/Q+dbxYFPGd8Ajb8oQR7mfuKUdXhEPRN3AzDy3o+zEMiA
wmrnADE4qqmv5tb0T+7frpJWXFPWbOe3KC4oFSie8G+mX225RHfsDO4BcNNoqjNOVFfMLXKHQ7EC
LlFQg21XWOoEHXud2NdOhzmwGbmzgqOeWgCvAlJ/ZQmbNjNWxtQfY909aXUNMxq6lfE2hc0W50c9
9f/QYcjdrr7Qd0zIfQ+D0+6O/z5uLoyUa7JNYwhmcVNzRdXjbZHzutIxPmpXDlgodehDXdYSIslb
Ze32lCzYsFmnDA0B6VBw5RSOTKTMc5Fa/lkry7XUcRHNsFadLAAc2Y1ZAcyNC34H2OTeHjk1iY2K
+aRM8rDdtiGvmrsQ9IfyDmfp7OEgPGxTVHl8W+IqIR4RzWR8jpS6CM9sIwApiQ3W5B8eK4IGRtSe
CA4kcrcuPZRmQjwtP0WPqbwLoPNQgKLEb6cyzGyDd0mGd3clTKqeKf1wMdnG0QIjh/DODBkXtH9j
AITXbSuRx9h33RJh0qjaPuIaRb1/LVtOqBNfOnHOkfklRshlQXuYPZOLv/B7wAQAV4QqYXCdH3V6
EoVDcS0cDixpwfTbRajJk8XxtJ/Khe09rRP24p15M/thRza1Jvos84ENC+GK2P2vXyiz/lvDCcNC
sjbeqsRGbAnBKwTFP5zt4ZieOq6PZN4Mg8ly3A0V+aWQlB454V62BVxRae4t6zx4xiy5MbqNo62d
b++bAUAtjHSxCq29GzAcWi2tS3u0p90vITPpFj8/QkRCull/dX7zXgr6c6Lx9MwtsMyD4iYdEah8
aVb5eeS3P76ZuUOcvFh4pK7rXw02qkvnJ0s6WlKtKvsAZongAlymVFX7s6OmvWBM88x5F/4peeas
ZzmVS/8tMS9V+CTgVqOV8J4NyA9IBuk7Qroldxlr7R2ZoNKXrGuvsQe80uDmU3y8xPKr4CKOxgv6
4UE4OWv6ya3If+V504vZRBbre69sSeEGpIiHRkUb/u71Q7LixTALOj/yyCc+pwhlbDdNLoHSTPka
CNSYqCYkzfndN5a7hhuo22GBQlVW1MWZAQV2llzpB951bCj2A3OUSYOqgpfDkpp/7eBE1kV/2dV6
eC+kdGe+dvh9JzLLywccwyLeE95xklFVma+xpC5o4X5LQwpjhqcyhkDXmYovBRC6EOpwlK29xVXc
DqSUbyqxza5aRv8ZsY89HyMpRd90ZNZ7j5mFRP2oDCRrMG2H6v66wC6CMe3F7HuLKA7WHZXZ4sWf
duu1bsIW+hJe8cQCNaN2GXu+wBbhl3WgQWN6TltabsPAJEDVwD04qd9TETMP87cOc4Az5ORc2qDW
TsnEm+hykMF6C1MKtcLRFjPLpdrq3/ZQuQcDtGbDyriDXk+U8raXzpTV74sqkBdl/nhIwITRHYQ7
Vnxyza0jtG9G75GW4f+LpbvHhtIskYJ+QgNSP+zeYlPPcCQv/ZiIj8qA0d47xrauBC91HsNOpIMz
Q9U8cyXCNTPBFcN3MtPCDdm80vUdz2BEiMpePyj38R6+007iE1GSUcZhhxg60kPEsjoQum+ZS3Rm
nBhcj0kV1YU5k3CneapsgA728teAPnebDyEESbx1pXn9sGE3o24IeATsgfvbIGOwwbX3SGMT1HDo
2ynEw3g04da55QJfKg72fS8oAdh2bOzn5l9lC0JAIk1xEo6/3lB3eC/SbneYlDUar8bMtix6VdgH
YqtMOOoVMjxjpPDRWbhuHA/4IPNmJMWy4FjECoyDhWHGvoYENlhTkQGL5CseUcEvrMKeE09XskSJ
nNzx/+k2U1CgmX+6tHiBFsCf12aKp3C4CPJn/hnD6NtYVM0AZewhVt/NR/XOXv2F3HU6s2xgs3jz
Uk7o+o5qGF+67RjiusXlvCifXE0XDfZ/mycJvQiKR5piVAFQR5V3u09ZQoGFIfqQ/wXe6Kyy971q
j14kDVu6r0y8hhNFrkm6pgA2jpfRFSWfomZlV2O0vZMlEV4o4+1Ip0hrPrP1T/p2RNYJQIZ1yy7X
wUa1WOY145DVd8cUlxQkHD2B4712f/CEJxiZ+aGiX0qjs3jOOGVyQfYswAEJUV0fbB0sqxITHMJW
RajFMquaX5S/D89FCxR0glubv/GeSM8lE8LRzRJkP3rvIe6ZlMLu6HJCfmIwx1cVBDxxgkN+eeBx
24N4c9TrGq09SMs8u1lHWFfkJGhnFBzyioivKQVRGZ6qV7xqe7Ry88Yab5myM6aRKXd/gu2bqrlJ
hwoUufCsD10DGNch4uo92uiiyrcXbwIc159CnJ4ZnC6TsJai6Exk0PUliVn2XDEhYQi4qWZT+ukp
xKKfOXYkjrpDsfr43xVGpVKwYOu3CexkbrOGLDEPONEPkn3kyOBni9TKqT/jHMxLE8wWoNVhhwg0
7uIAUAGxqNa1CI6w7hgf5dW7KEQ94nwEm98PMwOXBIiljMRgcos7a7zL/402izFw2dVVEGdMyB1u
7nmIaVryBI/a6KlMV5AACa+JAjwvJ642rhEps/HU6dmg5It4Dbx3ODmB4oM1e95Heh0dPg4vcive
v4UxwzU0XIqt6cjlyEUlTd+M32hGGLLlGdfovzGjM1MAKpnQrBHc1cfZLBohE4VZLej83eUCqju/
v3o8xnCKz1GKcY+qnZqPQrs8wtZGYIfIvcJt4+Xue9K+DLIpMABdTOGu9W9k3MlimJH2/Ie4aD/U
9E2MsUhgelfU0qnOlIlqJjoQeB+5JaSiISnTNJ+iuJFrbqoDVm5t6jqnhO0e3NQ0vExX5UgrroZN
JizAEUhhON7N5UnlYTDZPJVaqdauj6n4/i+QyzcEBCtjlVlFcRrUZzB2GazrM8XZ30pJ/m+p67NH
v2clmj+7xBByOD9D+MwpUY93jCZpBDR0TW3UUZWe4Uok9upD1qxpqJW+L0iyqBr0gJbk4GOqj8SJ
NFp7i+uf4XpfqXLq78AZuMaXaKQc6/3lArxsxXaASHLo2zSOyaG+fgg7jnh4xmq5DVbov04ZsP5h
ojbEXRdliR1JNeQS6hHQyBG7m7kfwx9lZT5vbNktP9/0RPILPuEBSw4tx+kunLf1/8e+4vyW8kDU
frW1nbTUQY91X05qtuYmnrffRJriWyBcLPN/462sNLPZeYVsNqeAq23d/I09WFtdiO0Nzr2IXTU7
yZQn1jFUjvOxyqxwtaR8NK/oZibqzBPuiAp2FNVjNT1ZxREjy8Kk7qaJGBTWRQ0HoGnun+SXWgC+
BSbqpombZFw0BKeO50vmHnFWWwlzaS0MusS8BwVn7LcadE2WFnlya9/8mWGeo34juo8Lc9BVliKY
X5VfGMZg17bnAvB1A5SsPNHxc+d3oUp6HylOD9YKsmkilQbBUwpmoJTOPdW4C6yZI7D3uYZ0opS2
2iFWn3kr8h5+xaUWaWbubmzNz0/g9ICIVkjVMzgLrZI9sQsWfL2fE6sgHhfG4D2tR+RugvZDkJGL
kHcjk9x0NIBCOW3Ok894u4YC1VvQ8PxcCL39xb7TGcLrRGNp6hu7N7OamudZgz25vQA7d+GZZOlq
Vej7ZYAyc7fI4w97GtFV2XRUQvdJVlWkbbIUd6KpgBvtD6lzhRwoBOniXAgIooj/19KPkMcKWy59
K9Fwq1QYdMXi476T5CTaUgZv5T10NIsm0HBxtfp5+hK/Yw4jvj0jAJzeufjK1ylhhH9moBD+4/3f
YxgNUn5r/0/1rlpr1knEqTLg2nwnHDXdCJs5tdjRmU0RgNT7rolfPt0CG8zr77WHsWi8XYE1d5rV
8AH8jMbWTVcxgkTHT2XCrj5Lgc81G8uPlIP1mee8a6mWxKri5dux55sbveFaeuCuB9GSqgd6eGcG
wZ22b/nHnDYHx3Ld37F3wr/C7icu3t9ys4xcXIp5zBx0xvsRy0izQptzd7N2tqwJEr1Sfd+i+/ns
N7RXSU/QDxR0WDTgWas11nh7u9RKAW6AM1CZzeLLsSkR/NHl5SKqOSMSJl6iwCCio6MN018W47Ft
JKqH45RSDorTFCDegVTIDqef6cOqwgVSHbeQT4nEgWYXxH75ld1jAvIOd2Xg7HdjchDIpv4O+6k8
RGBvFdZR3V3s9zgi6YK+YJibTPqNOM8Jne2MCcpJDzy5dqQNwy1ivoDWiZnAZ9kbXolBJYqTITv1
+GAOcq4oMKpxLbDSUmd84P2M5E2rweIL5gbyejhbYKCp6FuuAj6y/L0GHJtjv7q3hEfmOaC4rpij
e7LQUOTVnkucEptMjmT9pi9fOE3i7kdn7EF+Fq9JK0h+NfqFrJ7OOVQDb2795RMPbWlZZUwVO4o3
QhLbM9u5mrTxv7ATuxl5ttPcjB26e4S5rbZ9WRq0bjsSbLCRxmHZt6xP8s+pFo/018JrpLCAVRJo
bbuGB5colrCvQN36UzJbA6L+STcUyQmVjiY0SOyA10TzHM1EFqbYuR9TNFU3Y3JcBjF9YrSi5Mta
hcwULRJ50bbI52Xnvk8stxn2XOc2/E/YG/isHfN+ALTGZc67XsLoA/vfagyKtlVX0V+vSDQrQBPU
3gDCNw9fuaxeLtai/U2/k4CWs8H0TYrJ9nNoDtTahXTnjm3JTAUY5oyCpmQejetiCwlS2ZfyGQ3N
Ca+CT2/YIpgtUzBv8btzdJz273uJadEomG99dDi9qFsC10kNVoxSltuz1BVdWcPcWBUZFM2ia4tR
b6gZi0HrvmDNizG24eZ1FJwTuPbjMmZAMoz7T3ruIIZ8gi4tzwxQbAKT+q49wMdUwO4lIZgJp++V
PfQBB4Cm+BxL1eaypnH1n683G9EyCX+Bt1kQhfAIsJ1RgZtBRGEdpxPqGKZDZeEpLxD8W/VmpqnF
3hWfHl1cWts55oHHc4zt17YRsNuHJw9ErSksAipMtyje0RkASBILvjHyLMrxwv2d617e43J4XHUz
IFvQxcm20I26nm1Fo+Dm3DLEUwqCP8uJ914mrGJSvgFU/3ObHtQdsQ87bOQAqcHC0XMfUOpHzjw3
fVIWCs4qE6GKABsCCpTi71/ybNqsRRodtxkzK6YRtStc0c2wtBvAD9bnJCfEdJ9ITHvB4N+TK0J9
CpsboQ6eRsYvx2iHZpwKrWfP7Xnp+K0s4Ga5+WFvwSXTi3vdSLtL83QmonU08750aA47jadjNWV2
znRVHgSKWb73IbKKHHe7/6Y5qif0IVkKeymzkLUGKg22ANoVxzxlN/lcdKSGArLD0pwG7y9LGMQd
vcmEFCx71+XPRgnBYZB6/D/nVlpFU6QaMrHzEnEhYbNgqgdm7hoyjCLGNAtq8mS5zHysx6TMAuVv
v0OizyM+A+EYhzjDLZSDO6/Dj7akPrm8r2TdcZ+FkpSk2KEn8URegiJDcBQCFo3v7tiOg7e0HHqH
B6rnJa745vT/ehChFJaDNgPxJVIG3QM2qCEUusLoKl80Iaw0bbOOKFAW9I/mZwC5+XAuSy5YyuC/
MY+ZNNMZlnuFgL/8Fvl+MX98uMaZ22BmrUVuRj2pNFYHGo8mGsqS6XXiR4q4Dse8KzkwA7J5ZpHm
uaJbxZDG7z/0cyUK+FyrJdfDWh1hZ1VERIMlXQSgGJOtxeW76QCuRS7W+jMp/9DBmBtjB0wzuLau
UW7iaAIS2l9fuypWYu5pUX/Ek1eMl9TfYSbS6ww3r7e22w67F+EUgIK6TMs/39ImTgDR54ETznuX
lEpQush20QsK/TMuySPwHI44/VdvjYNojInUAp2e1wQGRCqUNMRu3xwu14DLEQZQPszf1hAhiU+m
AgvaNmenaFnpzSd140Zgrw6Zh4WHzmjLTJg+vhfUYvUr0pliz/IzlWQWmaUeETIftxdUVvwmnwVe
m+15RpdalviDu+VqclVGoXfdktq8ddybWSOjdmUTSDDnlX/Q45i8hWkALjAoREN9OYE4sHGteLHW
eki0XhiocnDcZPNd9wNviIaK2F98E3aXAM/JwK2NqjKCfpFiE+9Rwfi7VCPuMS4FuRTQvEbP6msi
7Fel5KwiUboE6ZONVj5FxceIbmdZdVxPFbPhoyj80R8mcaAX5YcBhBcmsjk09QEc4XByvzyuJa+u
xCqiPS/m40k7js41CoT29A5X8qqmAAeS7A+8bdqC6TXcTASK8AUGmAkOIRWceO1GT6TrjCHBSklc
PuJXUqvRy8ieprMBrCEkJYTEuwnoRsBPKOwM7xsfs1/jknQL8XJZRsyGlutcsDpX0qX+1a49jyiy
3xB+yYjTmbnGnDJuXBvnrslo7c7egw4vaVRvyf4jXWUUdniejAkZC2XLiEsZ1LVlOaUPbCw6mSRR
85rhB3kTwCkGgogSnU1LnR+mYIxFPo1FhZZ7n7JvMToMCUnaOld5lUd8glB/Q3TwGTBmEzPJ3VEY
Aypyz6Tmxg6frXXiFGDAeHiQBm7V9JbOwLSibGHXT30DIfF7SYnDWFb0SdJENaGTbsU7xiZE0Fmm
je/Jb+j2q5uPzkwfpubmMduIRe7qJV9sdMztBXJOwgUCao8D05ZJ2bW/SA1FgVBfhtO9LcjxFAgj
XvXq3AUMmbjWyzQe/SidprjfDUhAshXW2ls2r2Kx+jmdHDB4+2by6mo5djSuUxstwde0bsPLFlG7
m1Ax/oTrvED3YFLVIJmRDtC+giQF6QP4heJr430q6ogjGY/kwEHWLlaxwjWvgK8ZyvYOmJpV3K1r
0rfIK7ngKx5ro+koYqMppClyeqAf3KBeP/qYYFwkgstuYSl5vKclMHEWPiXaMzmV7f6AYcqA7KF8
szxKjSq3cqCGKNA+H6Ig72YBPT7xUSDhG2NitHzWLAaL1JR/413wzSrpBdP5iXPBAAYtf7uuOXme
KsMf0kgSrUJQthNVpYJALpU1Yu6OFffL8CODqiJvQGzDlFJmX+KuxqQcSqDkkZY1ZRnr2eCirykQ
7PIF4aeZw7DuMuw9/kR3ZfpXrz5DVs5IRgMMZS9+cLu7iFBPk685GsCyPR1CIQQ5+fJGiU6paYB3
vGOBr160N1GKYqS19tonKEBMC2PKP0aZGP1akjieOiL/uNMyaZbNlA3CRE9dCtsrzD5wLtRATHlH
p7ygSC9uBW1N4r+4gH6zhZ8l0XoIr34reoKk4pd+E5N2ACAPDiXxlLm3a3lA2W1d9fGzXl2hJN9/
LZfh2ROHFBgIFTR3lJmueST/nFTKtjUhYfhWaeQELGldCXg8mZW/1sZi2gSWDGtBmPjCSY25s5zM
+2A4QSfSrXvrcDhsn8ti0TN8/cOd97h5ztcOTbiKo9b3qAK9cYU/taXHPahasUWOo1hQ/ic0UDGF
JdxFu4jmiTrxtRXZwdfvfDvy3gXVp/zvP2yDa6OULrIiDaF7ZYldjK62HGvz7GuVY6WGKDXh4wiQ
PsxIV1mH7km9GvWQr5wEUvCAV1PHdpqpZrFP2VklF1CHoO7HcL16Q5a96vIM0Cx/WtJUAXQvOJbS
TaCeCitGqpq6FNOw3AIak0rFqw/01ZlgjX6AHNk5GNscGTbM96DMNCzz5UYDJcNMZCJB7/BcvU+v
WEvJBTooJWxDkDtPi5lg/qOu5uJTIH5dhxOS/5AjG6pgnpCaxgx8X/o4sKhWQHsl9TQfpK0lZUdo
2hTVUUg/ETQw6JqKQrtUCMaHiC7N0+XlowI+7mHxRF2d7tGK+FmrHR/Cc/HPJwbsWa9iqaN4b9ns
pCacqSBo9GiNnS0X2ERw03WbqQL23dFDUH2y/c6x7LJpvJVxVLevgwls5hY5izVf1Cmi15/MMfog
TBJVDZ5XDzXdb4P4ECG5pga6fTvI3XKR8TI059dOiKhwZChjlNCpL0O5oodtVN+5XMPswHNZvtsj
VZR5KmILU/sI/lvJxdqljjQfplylNJ4KYKWqfOcGqz1+LTNRa+zmUtJA0PdH4EPrlB0Btd3wa9Wc
n6tZH+/OgAad+VQj0NQLRbIIgxQNRVar1B1r/WaHbCwNTrlqXXcSy4PLhcGnxSGN9IafD5p0eaH/
YD2uLlHth+kB9flQTqzzXZp4Jbl7mP6XKc76aKxRjMi+VkVc+mfpJvcCUZeQ/2fFezcltkI+t569
WCaTOU80fVfJXtga5oO8alL533C2/PZ6qOSqdp64PFAIodZPsJDlsdoKU1muwHPlwniKc7jPgp9K
6oZd0dEDV3QaIcUcrOsNn9Q8y4FtGdfFAWTKbwmYDnOOHa6ANEv+lbYtD8EgrDh0/P5pzTQgTrxR
V5W24RWWD/B3ZZTYMbDEJg78xzM781jDomw9CyrNzwMx+6Nh7+Kx+eIQPS7suxEYQs1+iPDHpN5a
Yy31kjQ5Z9JLKkiRPwkvd923G1ru3ODCkQwNBipacZz+yFDuPjgcD7kV7MxmdKCvO1MA0tsS8BW9
IaDBP2ohTQfqVCb181ZRJrmZRi1kWpXh/oJiTxZZhash+hZmNAEA4Z8xiMlg+fhhOVUzUtZqHn3f
SXDTMTwkcYi4oVm/jFuWNEeO9sEEnzyx2ivo6Ku5IqanlplR5bSAjIyd6wXtEzmHvm4imIlzYqIx
l/wyiGYaykdKIb0qMDtz18VP5afQ7+cwqKNAEP2bdCwP/RMORHj5wUtESOdUfKrrNgkCff4IE9LF
b+jn0uLd8qVE+viFFhb31ays/vbHsniCFSjlijXUQvPF9iJn47LHRr0Nw2NiD1N3itNm9AIgYZ1W
Suw3CUpQASSx0dbweX7p5mf0Xb7jNPNaaQ3oC4tcgRRpeTh7hPvkaJ/Zi3R8AcbQ/bzjbgCHO0LV
ETPeRZFBwXvzuDoOYqgCxN/eeEuWfChd83oOp6upyOwViAx3tFAEZmoaG8V6a+YvZB08dUjC3abU
y8TlRwW0BFctHLDoW+oTLDH/cLv0mhO9xxfmpMSEhj+Tb/x/CXP4RiDHOKwNh/m0OK6KnwNqG9Rc
VBwrHO22idhwSXS3jbEd6Ezq8vPT9ZJ+48XgPJZ9wHNaRx6DK1Y8lCy7QX5j+BN2yLPR+sw71KX6
PNjUyjjj+w9egTi3D0i0ATUW+LqkbRH1EwcY/9Hr7MHh3wSFvP/zC8h5aXVd99wJwqLdWFmWVmz7
viGMTY2c176yRMN7zSaD9HWmG0+shywbyrA50sxiz+9H2tf/Wps0d/kvS2EBvLt/aOBOrrhb8reE
nx9iv4e0jtEWazjGkOf2x/UTHXOGMdchNe/u6ht7dNrMeqs3DhFhjPpXBvF05PvFaH4519gvMpQr
qy6x/Stmjxcf0SASvdsLtuNrZ4lxpWSocZO/M6Ax0y+T+6E1UhcChNVNReXtxJRwkv0M0dVECUsV
4LYMccBV2KenRYdegeMPzJx0oBKQfvsLfs4i9CGY1yzmFOyZoPvyQlgGwtUSVyzEvUSvs3Jf1tt/
tJM97GNkMdQ1WGdEbGbo1fhkjal9wKbHjg/ECGnAUT/PDdXRJQ+Az02kIF50BUA0LmSCIJwLoF4P
2tCqrE4ye9cDaBnHfhsOi+md4/NoScxUVVZki7LJOu5xy2rlMjt9xfpISrGdQYUN13F4pVdZnISi
p1b+53x3mXmiPNWIpHgwnENW89VPg3GVKJU4/nW10fxa1FrCGVUoK0goVFbFN/LrZO492agbWSg5
Rp9XMY8VK9TWOzOE/9+2iNkQ1oGzYXjKeZhqiLqgfE9LZVJxR8mcIe1lRqz2GyVsATk/HBJTRKRx
YbCK29QMGfrwhmut6BxO2lZfkSPsdBs5wGGVzYooO+nM7uAAyvg9+tzPFpMIZQUnpfVYAfI5EgoO
6uKsL5VGBvPJGyuJ5uXDI/yIJB4o91mgOW8z6nZTdXh38eHnKP0hdS7K3a12DRi8sGXMnZ0+1CQK
Y0eORdV+21aRiB0qVncOQw+yXB8JzEZs846JSlTY0bd3ojYXfJAYtIAQoZfs+W2HR7Ca0fRK3htF
84JxWCCPAYi1nRXAAOZU2bFZrXxJx2yw/9SpFWSwj/tMtdYhYvrhXZArE0d4etXFYAXRkpO2/EBE
4855k/HGDUpS3x6UKjiBarsqYa9tB3OVK+KKyimnRUC/rVtBsK0dgqfMK9ZCNeleYZoxwldk6s1o
ogV6oN3XiBRli13P0Ed+xou8VtLg2pWfwEFuuVIo8WF58Mhm9hvzr22pLf6R2Hiw7XFQA2uYLqxH
aiZ58BYtc0DbLgW1zzBK30dlFG6bCzPfaXr9uhCcG//ZlCSo1/GpwuChIfWcBRMS2PiHgj1RD8FV
SMiLupGvhcFRYh9i5zzmHnJEwgsN4LDj51sryQGhjrvtFE3k7vZ1p0ph4LlinQGX5pNkFy9W0MFt
jzGIZRnZKVrqsX/Wdq9BbyW6S4U58JyeJPQ4HWLyUxm73olZVRVDpI5BPLB6HbCtsJkuQYneCkUj
vgg8rGkGF8Nc5fiTG/v0uNCYxPhGGq6T5pPSpcTTzs4ywtPQaPQDV3vZFK7tBnq0ufGS8jgpyDPz
E4yA8pzjeMeDEHAsQRZ8OkDqBWL5ij5XvR/HR1LxiYA0nIeOVx7TuufawrhCHlnnDzfdkNObLT6/
TzzeImmAXxHe8kUhLDl0D+CYoyQ3whhL2kiN2dCk//A7/m1r3NQpLvl3p+OnD+E4iT8KjENl47gI
rKrmf6BFojCGGPrVWTIA86Q1MQjd+nRdrXhrYRYmvfooT+wvDtDuNR+ROZWXo7z4FEbCJPy6DgAC
wr/C2sZnUosO9TkP0Qi+IBAvplPIYksc0gKA6mJnsFtCMVYukU4i057IkoFBcCuL5yNUv+aB8nzf
PAjPZHXSQtooahW9BIMIEDJ9euWU2yfx20vww8mgsh7IctMcyeA5gRiCZdZ3uYRTh6DoOSPRX6ly
fv4PjP4vCKdz0szRF//0FZ4catZRfklbEUt4cSeHBbP1rV0jRluRO5COwOwSL2E1EAA8BXoTnVSd
R7mmxLSqddhpmY+N1nY8v58MxJNUb6SHBM0z56p635EbAEaxFsFPlb1pJOEmJvMkxdSpomRMch2z
WyAjip3hDjgWkiQGrcKrG44q2XWaxG7mmY8RficfSfyal1PiMn0xNzrT3iWh2C4gHu5rWCYF0kub
KFIPnpFK3TiHlT0gO8mSzMwavf1dlBAU7IlxSQctCaYVoaqG5BzQ6UF8aqlE5wpzeqC5YkYj2orw
rR8N9C/O4wMYuihLqTngMkIXSYoTaXZwa84MWs1nYFZTe2NLKrLABJcCT8DKqQON2EIqRVn1gIRN
tC6PH+uKThXIXF7+2HRediRUcp+rkw69irrZmcE1UFbvn+pEUPvUHXSOeGe3DjuUXba5/V9j0Y5i
EfrcBFuXCEolv7bPC6zubLk8JQFqX4zbOB5EQLsltztY/vHTrYtuz7EEuvSEzai+s7xCu49rkN4h
T1mHyI4UAUJZEmZrkz/oaPki+gaZifkrpFnGVD92k6EzuzB5Ma3MfvMqoTIfBU9ujdpyIysrsSCs
y1e3/qZi6wgmK0m/mm1ZLvb3mK4dSGVp9travYM7scRnZgCefBlh91ZsZTOHluTOacVdWVRB/0G8
nfEZE0oAl+0rVijoUqR1HpapOMIkIHvFlAiNUE7X7P4xqi+z+6sizISeG4/hI33pwI7lZOKPYrWG
LG7t1p0anS4pU9NGNsrOOyA1h1HFuvdNLPI4OFaOs5rpo/k/8caBwbfFUMLPmSJhpg/fBKNqvGHm
uHCJTgiH2FJf7yzutvPejrF0W+2KaBtEcI4rgJBYhewzWisWmH5r4LgUMwoeXWI7ARgfvqI2UwrZ
uWhHa48Vu6R4y36wXukifduK6MXLIE+g9CKGlFctcJRvsDxWvwLXruA4IIeCYifEHperTSRp7mXN
+9sXmQM4suGPw8oVlspGBziQUC7fM4iETHkzovAybfUOZrHmbTVR34YhiJYw2T7aweitROF0uhyh
v/KWlXZj4ZmqHoDw42lKv2lK+t5z5K/BE2+/DRa1tgIgtVc3temErkjotcTYzPFOLVqA7atsKVIH
weoQ4eYwJGGtcUXEGyuTNWBqKQzeQePNFCrfcygkJPpD1pfcdt5HqBbn9bjqM5LUHkhVndG4g7P2
w2coqgI9kYHHt+4o3BOPFvVbr8llU5OtPzEFcHj6Z+o6JtNwqay7L/1Npa1dVlMlGUnjPGRMw4uJ
ZN7tR+9IO/QS6ZvDWLb57Tf2mmEXEodgdiN4X5V++UpHAAMw3ESo8IQIYs06k7Wjag8HvT1uUNKL
S8j0mdzCuvNfHzYpuvZHMzYJMFyFRrL7UxZ9K6sXv/Q5oRKQhr7tQZZRDrM4V3ncYEHQkTCfyxhB
DT5NFC6JkXrqDebJqba/eY3cJ1+irg+r3I9HmNDDg7xJHupQ63q4Rxwtj0j5jgA8FB6Z67fX8ezF
XkxfQqnouR05EzdiHLVn6CsQ7SEt64bMeM72INg85Fldu//WylhKuxVKuyeMl7GiDRDbEOqvU+hL
DaBf7f1gn5u3hwjlcnwELNGa1z8FoYfevMgk32Jr1itJ0BiOCeADQpe4zvMsT3dOJY0Xrx33dtLu
rOujCttHLgP3fLH2DORB4JNr7ASVvZNhNY4VIet37BXGqr1Wtm5zGXxyFhbakk2oeTivplfl6xcW
BEfnpJBiH7gP3PHUJN3vLiM+09Gqlq+CD7jnwAktxqSP/vibJnz11RQg9cu11P8OKWYxFx+36ar0
0DDDPI53TXWy/vodzh1S0mdji1w77rczGxkoZfxJ7Xff9ZwTAgwP8rcFiRSioVbzU4mkuOFTEyC0
S7eP7BeBsM2EwY3hkJ2hOQV0dmrQB5MhvyYkCl8mx0Qq6TOirEN+BBmSnQPvuAh1CPYMY0DErR9Q
vawlhND6ETWvCRS19pLt30KuAFEV6Hdku3YMHtyq2d1V54AuipwfVupc4JFRKQTJ7g/tg05RK5Hk
fepYBzRn+zNprxbJVNx/HFhGjd9fptqqvx0pXER/0S5xKzRJY6BNCZK6riBhQX5J5M9CwJTbV+oS
L9FNaCVCPPKPAadKTj6xcH5SgsTW+ZlutsWypmxyy9whjEWEBVvHixOBHAbNkzBK0izmJCITMilK
HkYYl0TvV2wAUTIZfb53dI0jwcKgGpd3V3IH3R3IGc/uT3UYycApO+43tlpIassZxe9x5neYeRFc
aC70yM/t+bmXZouU86K1tadrtxYsaMofC4HFpAIBIEeD0E4rk7322DUNwxTpOYtqx2boiVGTtAg6
V2QntAT34vB3kWbM+rH3CmX+6R5wuZqkksCskC820IoOCK8abAG8TnlTotZ08anBDIW0TPLDVdc+
xEYpWIfF77++NgUfs6CKOr7XGyQBltZ4paM3ix/5IBcTywUJpIW+/bkYYLTjAEMYIr0aUrtCR5Pg
wbPKPIWtKwPnqB39jIeTCwIRW/LCmkE48OGQuHlvJiF55+hxZMghCTIK2f4/anQe0vkAhNum3tix
pZF8HZRojVa5PRTJcumwYJ0dWQAZwEnl06MS0m3wi1m8sm502mTj3ebos5ixGS60s2acWLAFYY1P
iMyzjkwHb1QD9h2k7rseqcVtYn9l6vNvyt8ncSnVmZ72C0TnnL8vly6OjiXFOBsgimzFQ83Ownlq
+1FBsXF5oBr6dSEd2XIX1/RuHFq3yps7cN73CJTfLOz3eNcXZhmCewPbOxAm5cLvMOz2yFe7BEPa
YpDCeRn/UnCMIQT6eq2JTbYUITXKdbZs0uyOVaBNkctOcQ9FmbH9qhcU9E/En1KI6LP7AovVVdTY
Xh9MSYxplmqgH0Ww57/8/jj7MR3x/QmhtVG2dhahSVk2noswAwte/HF4+avF2wtEPhIwtDz7BA6y
USlMZKagwYYIdMc3cupFFMS9KVS6rH0rcCxVX5E5zI0dl+40ED/Y4QB0od871zAFTCc/hx6hDoEm
szSa33BVP0AMvV8TUPtWl6M7422geQ4YI/aOag3TFIxByazIPJk6/bOnXtQDIQ1FqsTNacju2QvW
Z/6QIloUUkybPUqGqpkHbh1/CcN42Eg1j4Y5vCS6jSgWg49JM8rUq3rJ2DEMVG0Wj05HoEbE7TTo
fDtqU2xkQyoAx0i+pyfQ87B7ENmtwWT2xazfVZ7B1S7tt8ZB36Or38sj3mAVkPq+RlS7ZVuhuppe
NKKOzAzHAIyl2U2tPu/mUB6WUebr34zOlkD7Gjk/0WE9Ye9vJIx8y3BoE8pNV6083vZ0LbZXmruS
fRJSQHuGUc4mOXx8nBeZjfZ+Qs9LdcJDY6IhnACxdLq3K5yjJyq+J9QqAUxS2n4jde7nlFPvwrEU
Yelrg9YhjqcgExozIeh6p3u5DiziEaikISx4K26eCnznyZ0bM7ByV0vBGY0DuIPhGzfBGMRkCWjt
lcUnZRDWy4tAsugHN6/HaVTwgdGUXCgemFjqI0ZsRtIl2Ak21feFzLeBa7gy7RZ5ZzB9l6ixiE9d
gZGdACBoBv1cTvtF0EEUZgKPudwN2lhDORFmkYPTscBzj+5ck+DBULLOs8klXOxGHEhVz3YkH0in
ZV1I5LP0H3KeGS/sUDi2oyIaaIW89FJ3vkRmkkzerFn+23n9P6t1HDAKXbYpn+yCMQfMmM1oQFYZ
vOGmJR1bHdYxXmxPiF2DQgQ/kN9MtmCBvQDVwGXIUIZ+TqXZYrq4nJ0fZA1PR5bwzu+ytogE4xKJ
nr7P9fBb6u/cZ9wvK6lffhH9JSxbagq8BZhI/2pqZt9PXIG+hBaEjC8cfP4i1me9D8mJlvNseQ5l
uU1kl9OXhi6GHP4ZrQiZ5dDr4C4vJXrn7S3Sj/ZxPQMDGvoBdMGlG7A5Ir/qCmJTout8oLApzF9j
t4QN9IW9e5OvgkIKUFYhEvq/8na2nxBfDEmC5dlovuiqXhnmfDfMdGZeA+UFU+vycwao7Y9TSp8R
W/gaAokcwMFY58yJ1xQ17gUo74e/9jqd2K5avenpoCq23cP6qyDMVEVVz7IlQXJ0OIHjtDXAsTf1
pH0hIxrV+sUThW9WeLdvd1QrF0Qy18DDxTpP+qlLSKuMk/PNEYJsWN9ZCnKPk1/GNUyJN5info0U
m75GLeo60jrIhU6cgZhUo9ydZkQ8C9LhqsGJ8GE85TTz3wnH8PepDW1w7IudeYAmarTdTA7PXESq
j7JxXtUU/5sh2J3onS7LCCFFknoLcAjlwd+dJ+QEbfxEScO/UFLkJWfzS/s4KJPv+1L7F+32QGgv
ueQoMcAKOEMytITQXBeYbz612A0hdVh3G7yeI0aO+B+DD8wGkB9CV/jxcFnWlfG5yYjxoGN4FMEs
NUyMYsm1Td3ZCVl/py8dUhu/qvoI2Pgw8pEUn0Peu2UeYE2hAZlUdxaHizSLogY/hRwkJQ49MQqO
aol5V1+isgOTiAEwHBu53DkgchVvjR7WNfPVtV0+1Odiw2m9iYSvrvyx2opnEb/QI7b3IsHjVvLf
UtQyEGS5R8MetuG7Rk4VO29xLsjqVfp1C6ZiFOIto2BDRL77Mzh61aC61a9iTSw4EZ+i4zliCea5
t7xtWuCKUBgaIALixflhtTTX1CmBq0U90KNUCLXGTURVqOZqtY0hwlD3hWlNqnvodOm/oHLGN3bn
PL5KX/IQvQ/Yi16J1Q36DWD1NQ266Gwbv6g860+QA9fX4n9fxf4Ak224/qmhnV6AhOAckaxBgOSy
TYzjGw2STBNG1H/H9Y7UNbWaAyUIeZoZ+gyltJbakPoRcCwdh9Ze8WALZI0xW5H+G+WKAF4JcpVy
cxbtP6QNsQtJlYKHkAZwE87OVMslVp20hqw1J+j3Pw65Pu4uKz9nxj2diGOi4SRnGGBdNNcHr7QG
QSGyGlqttSqm6FJadEC/po1jB7sxzqprq4sScvjSDZ33RwzaMC/iiyIwyAG6VjCOsqvj0deEjvbH
jQTqQDgjpoWHUO19aSdgg50VdmqZVkP29JEcHKbpBWlvHuoHk8zVzDjR5S7CUzU/A6G7L7GyGOPI
H1YT0DcyDHgH7x5B+//NEAM6J4Zc9xNKuA6o3BNPGFP0XHrKUTSJKTHzayBEE7axAVHrg7E30BGc
kjHGk5tGQja4hC2o69S20tj74z7D94KEVEaikT6qxEo6tiStFAXy66RCvhi1nwEU/lPZZbGsjqGN
KBqp0Fj/mG8sOtfCpwfn8KzZI1BUT441zdG3QeJ9m4MlBZr97kpNpbNaJNHxvGE67+urc85BEgP6
XOtDqwP6Ffl7QWKK2vrhDAwLDiY0HtnkOjhdSQzMIMIPk8kQBTyj8TyggBGfRh5LMnzd73PXOfYl
rHMYVzmqLL0iTNFELrlMDsBEEHLyWXJmHYMSReXr3T0T54sELxGXNsmVkVHIUVAne0fCoHxlInzc
OqK88lzOAXYAG+PrbIj44EK3kqeyuXHJJBy/JmuYBDxAlvOpJfY4QF015yt2CQTtMVOlebM3Ruz5
uy2a3cyU9xn8aFM+yAm/9ExcuDNbPUF/qsv131SNQUpujvErH4lA50GMhmI8lbhUjUuZq/2KitDp
IyJL5o8axVdXBViSven7OgyTKNyar0gMTpXFsBz+oTIL5YUaiIzFyfsYfd5UOQcxhVW0k6IcuH8x
RFSI9v8pjUven/2OE4t1AFvn/lZNVZrz7MONKNF3ooZv2Y+Gbv1UFXMzRk4Dmp3kGcd8//loAHTT
CJGUKQIxESaP8Kw9tHqudlDMVMh6DKQdet0eXmPlBUJjIYwVDbc6R1m5jtl3mt4wucxtkNf5XIuH
4TwUwbYnFdSJVsSuRa5L4/T+BSCa6pukvkxJ3nzi2jyNAWtXr+zr+NVYN0QnZzaLQAcd4/2Ke5ZC
99J+9wf2/ErPCezDM8MDT0wJxtaFf57PX1HCQYYNlPCWz5WlxlyN0ULA1bJTnOvRe/FvVmtmK5Ao
B4+dvs1PGqUxhYglVKrgo3VTd7hFlIYL3h4gAnNK3XB2VkvKHAhI018bWj7bpXO7G+dPOduLoKb0
zlYYRlRpyBGgdO4GtFLCsZyLtzCQAPk6q0CIDpnIkzHX5x6t76HVEsE1EQiaCqSF63zdHtrDV9Fc
+ch+B756HoS7SmLLO46LzxGxS4PWctDK5Bij6AN7guERAM85B2cwCdLiZGUkiLv5Ye00xEnYm6yx
z9lJdmpKeDtzwINxTvWmHQbwP7XobDkW9hXK+NMWPXq/aZirZC+mHGlOqN3B5JFvropg2gZ7Gup1
Y7xrTdS8jOin9VH9aRe4rhfhRMPITN+i6aX/ODgDXnv3l/OvyafrLZgaLas90HTfSupv87VIRhHo
+5tarprmA22+XTV49OncjpqKnyId+TeRPF113obb12SYrducS5kJSsQpYaGPPYXVUIFcPDHBq79t
fqLNOlMwIvBMIsVW7hn0zS/sKbHsRGQ4SRvt7uTw+fJ2RUvdnIwpgllvFgEDcdh/qnrNu6N8w5Rw
HL8HkaJsyH5FE7dXIvceqPL1LNX3XSjd+geUslbZ3/guqKhR9D7yc60xa7RMdPuOlD4clVP02mbq
zmNUP+BVGjB/XN6PhUXNr12qw9alTR1EkU4uJQRHOfpe3fWAqjuYFbRlsOZw0PkmMCoVJf4EPacw
HHHmVrgfiElOH/uehihxyNsZj9D7nUIo3tSORmA4h1OTkxMg9ujN6y+yWV8lodKAZZ/8V5SskcVz
Z3wgCRMa3xeQYwco8742r7GAf3RtON9szNcI5EzR/dQCy7HvSQYRAP801JVbMxYXP2XuYPf4u6L4
lBpM6XK1pvZoJOhdpOmxeqcPdcoxCVGiJuKVReuvBz5moHJ5v1Z94V5VtJgkQSResauBfLsOafvJ
rLVv+h0oi8nWMvd6EDoyoT12S9mkgxXAAsuPBT6mcBvBZP+J0wyBDEhdRZWDmm6VYS/Klo/JJQjg
v7Lq0jiTBg/ga2fO5gfzRjrFUX+UAgLwTGSJwPMYhczdfic8tr/0/0CVGYEVabo0eNvW4dd9NgVM
QaRATNfoI9JbBFDDXEkEUVLYkgehVwW/Ox+zo9+95VZmsgFeXmtfqanya+zNQvRLEU8s/9tcvDNE
83gQ5AclaRfmKH7x8PmrP4kfg11fu7VocKlc6LTyWj4Qo64Ki1JBGmEHEjmYDwCmvUSTeFWGTDH5
51pRURlppFpINgf5AzKUd1SdFe+/oRhetBtOF+r5loJZIT5baENAps5FvUsnGkVTHBc6xHImMQm0
1dMtbCk/YBp4UvxdkZYCVcNW3VOibLuLh2hWrmlSOU7/G2FSXZ62r04jc33mrcbmExPlXxnmv0wD
24GmPcgm5XHM+xhUGod22mkPQjI3an6CbLD1B2hDJO48ZKsmooOAq60bUoJMdwDtJZ32J5gwj6yI
DDfivveRqQRvI0MdPxsxVikfEopO+nKYeTLRyoqHjTJGCIviP0ePsDbInkVWVeVGQdUsm3Il3GbF
A+/80dyaG+TivNHZJ4ITPbDqIhvamfikHHKioMq25gELxtM7E4UgdGTQOZkMoHueIyjnSUXa4aON
Vkmo5vmFXq2XgqrS9HhOuYxyr8kGgucJSp/Jk4f+ASUDF1tsGeuSo2UNBIskrvwBioVtEPdUB2Sa
COGdbCvijSSY1eAH4h0wvjLL5fUpBabNunUULQYh8ggokItz+RmuxHTN5dE5iqaATQIqqRmK596x
5UImNreUS0kWWpxqq8qE8Fg6THPVfz2jpfak/BWsjajHs+BAP5TXVN7HXV15kVuC6TdZF2VpW9fz
av/weDzagjCm4TH5mM2OpkJwZm0+dwpdMHYSy6+EyIGrP0/t2hdi+SmBymxZFG2k8GqVzu0f+W0Z
lOJ4THweGnnA6lWaOOhUlqc9dx18K4r3ik5PBuotAkr7mdiRfHoaqojwt90Oig6yC2Fcn6wRVVUK
0Gri27beHEUR5ohxhAQFKWg6OzUZkpeNq54xRcaoIAA0iGftPWdb7neUV7fWpOogOb8aAfsxZpbp
pID9YZ2AxjWiji0AtqMQWI/aD79Ww5TroZGPfKPR0aMda3nTNe3zLNbv4kch8w9IcMRf8SJ6vmDY
tzaRHyOr3c7kUp1kwDQamni2LvJAkeRL4EdVgpFVex5a7BGgn3DTasmcs9qqyGOAM19N/U1+cO5i
GhtEhwFGP1ymBEb/X8VRLVy4F7hwi3ka40Vk43m5R/pDDRS/SFGRYUnqNx2acrk6Zv3T8cPfgr7S
hVxbGeAd/Iz5lD/fq8wAOQiO4rCwQzfRcC/X+pjkUlNaKz0x+8ahys7LY222OvCKXqpqdl4PoDZ9
cu85B48xUNCMtE9HwbDexP5WyfXmGPXCh/JNgnFZPPjgSvvmCfhyoCrjEqx91UEvzgilS5Xo/pnz
QpJcm4nndwPwbQEpZ4IlXrRl/txkxnhnTe3AJW7K2Hf+PTMfDGOTbJqiCHN/XFgnqWYH2B1jAa58
GYahyo0yL0cE0dSZ1tmgXITdI090qvl+gBRaBWa/10wDTiC8HWVyRLHeAy5xpe84maOplXqwlrTm
ivPwipT8+qlaKjLWB8wRVTT+e3AdanMOJrupVYVPnPmjWm5st2HYgv5CaRxVx5nh+H48H8Lf6Oz9
xU8+Hm4llF7F3NABC+Q2TRmNg+1sj3+I4InV8nDvZd2hOvW/UVOlHcqzCZ2OA74Wc0thf1r+pixb
Zrfo24Gqbo4zCSqQaaEsGtb0REsBMpUVfcDtZVQTqnQ8QuHIqp9EbN9LmaBa4i11tRp0Y+o3eWXC
oSgyP8QIiFM+QH1y6ZVA7SqxedRFZOZbyaOoQw6Q2YUz+Jd+L5N12xahivG3S7avDMaTIGlGJ48A
KggH3Px22Ake1i+XUQepIDzvHTx0XJ7+HHGA8zCDzObIVz7JwZDpTcsMGJ/X5Sm+SALeGFMiAVGI
ajTNQnQdAQgcBop15l7WNIgkdIpDOz650fSw/Jhr+IUIHVftVg/phQ9T4yTAN1TR02eOFHiPCfn2
1+HeFRT2ihCUprVB9lgULOFExexNsSvDF9Xpc3VmkSbwo8wvspl4DNMgvBRTcWHTH4FYvNV3CmIo
7bbJEjWwLq5NclEIYlaf7nuZfm6rpkpM65V2H1S/6XZDRpuojHQA/el/SPiKojqHo4v5qpZTsZcK
piV9+Vs0SSR+6RUbHI1Zpk3+HAkbtSAaCq8aFsky0DbMg+qorcmrB+hYPuNg138VBsomn+GH94qH
Gn1n3kEiYqb8D2c9f+EoBqaQpjaMv81wH/Cne8FDgjwYZRyCsQtG4CWjyIv/NmXk7V/SBTSEi0UO
/yvf/2Q9ZPi2ifaqBfe2zCMBusxJPIXd3yjtAHGqIRKdEJ70wTSBX202qlUbaAV6Biy4eOhw/ScC
DyqfN2BvvthLSDZGTunLrPi+toN7WtyQilhdaAO/HWvy7jJTPfGctAoRNeV71QI+Vonprg18KPlp
NwrP4ESBEQoABg/ccK+NjwDUwI6GfASNXKGkxd1Dv1u2rjgJ9e0N1QUfxi/wFT09DeBThM1CbvDu
CGfRQvtnJ2DdvyfkK8wzMjq62p64VPjAbD/2WFWY2+YM9dnZX/uwFYQezy+yxwUYTgEHa/ZAXbkS
x52OcWkDTDveVHqGyH+wGwt37UQeAdqBaOzkzi5qGpQug+9RKk5Ra+ZVB9eooAdLRYOaXA2lpLem
iocO6O0oK46hJOcRhAeNoTr87L2uum6vklK5yW/j4s5d88pKV74F5sAtqKEdCaAIf+bIjYh8PtXB
AruSSLHLBJP72zqifonW7Juf3CbNElFTmLWk3Y5iNGzcmu5IqJq6A/0Rr5rYNSJDSut1z9ucucrY
lKsRffhJAqb6gQRI6+KOkzIFneWME56G2JzzFRxBxA+Pm3mMyn5FUb5SqPlv0qlN5+Q+h8Bh9mZT
ENoi0Gj/hya+qhvtmDNHafnhL+fZEVhyucuQ3faHYDM3iayLeEVThgzqp2/2bs25jhi0v6l3bO6R
4SblRt8CwpgxKOHyui1VtAz1paSLsq0cRoLY+MEp5dmduhXKlUZJvzylxmger6A++fkvseJCSCdm
8dYCZgk88dgZnVE2+onVWQ0jjGvo4080ZNGC27/btXmykY26PtrvjKMaoe0Y7+r7zFANZ1HPfrkY
Qz/pySj7xDx/FN5nDWz7fYyZUF5h0bfxzoqJrzL1BFepIyhuH7BMUqH7WcAzLebeCDZci6K26ELh
h666s1gNId2gxUMMRHMattS1U76eUZ3hagpwa+AxcHv1DLNSe+XWxJXmMs8RiQLG8RgkgylW5yvG
tOHyqfI8yhFRJZXXTh4BF8mHjK/BVY33VNosW0tAJUpayY+9ggHP2qbJjnIgUDhF7KthWC+XT8v3
aAb1WFIUTDIrpi4V5OmjLkdep75nRDOBOHqeFL9bOP30/6KmZFqX8JB1MG8tLB1ApoIBFCM9jTnP
CaSyMbXTQS65TRyi35Syd4nfVeAOxja4r12Sc7YGdt+1j1XVV3ltgznJHp1MkcM8PFaKyx8fPv8C
v2e5jeEtidxpJnL6wodk+bJPuZJPmwKo6/93JAfvVbVdCTd2Gy1KcP86Et1n6Kx3recUdLR3fm4j
g+dXupGeslzI18Qa/xaB0YbVtGYRXbZHZmMxjpVuMLUy4Gtg6u8ZHa5Jq9tnJ1ext1YgCRbcZ/v9
HSdx4fH9OcTKllh9lKh+GHtKsu1tEximuYutthgEMRtyRdkmB9sFY7qRu92k7iFXCAxpLMVa9kpq
Ee6Hhtjl/+wnLGRJIOnjZY8fF46N0kYgIbf4TsZ3muCc3tagfxKuPmow/II6xLNWYoSO0dvV8Kc5
RfOJqXYmIJvY4YbgSQb84HmD4H6xQscnfTMzZiH/XoSlBDgVxkEXDEWHRcVI2KHBNgRiCQ7R3qoS
rhDxsJ+FwjukIisnm+7Kayloi2xxPUPyB6syAvc7LU0ksYbC+wNJDgecmnWuhXyERV5lr4XcLG+A
nOmyclFqegcui1CnazVnyilV0POW2DIKeLBj2ruoDc0THus+jyCrjT+8p77cGYMibmXUle2W7j4F
wDvxvTlLojcMwfjKVAnVZZ5OVLlFH2a7CSy36CApERf7MBSryBuu3Y3mCJbX97+o0feTtx+4ciTM
yR65Xro8GK3ojIsIa1ENFPC8sIXq9YX7nc8ti6HE5C/rM8AT35goc8t15gHvjEXiG9Gim8IJpMcm
WFJd7x6XEvw4P7zIcC0HfXfxb6+WVWgxEfbSEEAeH+sVs4q80ZIfKR0a+D4WyLJsUEYz6pfdSDeD
xmQ1yDSEF2+8ItczLp+i91BDjBnHL3YLNWR8T7iaL+uX11fkgJbSxksAp6SRh6hHAUSBzIDR2w1G
eQvziLCOZ6MW+8urdCX210AxmopQ4SzNFnFlOoLVa6rhBTXSSUzsPzvEmekh1rJZjLij2R1KlsSK
u923ZVnH1BShMmYy7zP9056pXxdBdSOq6yjYVoFl3zb4Xed11wTrWx9uNTLosJhxdzClfgXBVB/l
oSFy94V6zxLuwfnB/HNtCo8Yk7aXpG8zUb2Jaojg6z30cmgS2OhKzGV3VUd3t5AS488J5FkOtukm
P8O+fXkErFjMbyoSOfJTClFdf1R4yi+4jIyzirdOwWNHfsqDomAW49fvAafXsDeE2lCJy2xvS8ER
KISFnW5T9znAJvGzQ6hCc4vKntViaUEnBV/wx/tgCAufLxzooF2JFwFGsSZAEcwq1DgDcd9M1ZPE
IyT2XEDmcEUg+rq9pKFuRQlXdwCuHCy4OUDenUjQEIRaP9/rz0Mk0Z6xTys2y6uUhLckYFUTDE6f
uS5qBfWn8TLP+vt+m2XFNA5BG5kew55LEnVg/4ZSm/RPUpk0Dmy+3ehd5D6epecd1P41YYWFerrS
UZN1OFIFFzKyBVb2CbiHI1zETYcxWSxuoTWUmOtv/d8JI9bVTVvPIQdlqHow7QNYlcOn0bOIDDC9
37RCeeSXKrX1MeeMPmwL8sgXhKXO2ngG51PbBuI93cJfJcrcAKyE/wDj6yYwo2zI1owrZmQsC26N
paD+h79wg7FFL6F+rMcXsv/zCkUHWI7mj+LrP4rI/+YJwK5mUBIrDB2mNshwtTrnyCCk5rFxrdoT
kgrOQrgjnVVqGhrCgMvbi7EPCcVtEB2HFucpKG33gQzcb8OV7pt/I4hzpu878GFghLmBwl1o/M9V
lq5GsFTpLR8RuTuFE4enMMrHs3X5H6b09MnH+mOmwehofSgSdHabJy6JJ3+HcWcwR/ssgN22qsQv
A3uxknlKqGZNNsOraSTBuU/M1Zkk2xILdMXH5NLGlNvzsxZYNg+hLPVOJKidxvtkoiB0ItkSeLh8
HeugtuR0OWaQNwFGSj/7BRs4YJE92dfCjEsLKOLAiqqT1IexZMeLySYKeHMUDhPOIDCsfqsUluzj
0dFdGLnfgpeImTO3WbS/sbFQhLFADw6W6Vc647GDxJPg7B7ZR35evqnlbZi16evKFKm4Vwi0HodQ
ruPbCAdnOHIP6Hl4TaFqyY/MwrsJ28JKxZafGdKK4BO4RIo226mtgIn7yuVYYl4ZBYYx+RZ6W/qg
HcBi1b9eMydVzy8Hj+lqgyXEBUXOA+PCt6fq2XJMtLfiscp28yVp/BUwb2BrHbZRXr+sgVgQ9BIX
OJWv7TrCnuE64TbW4dNraI1jhLKnlnKkDyTzi+Wqb6aV2ixryJAzGB/icggO44uvlRbZareZSiNX
YZhW/qC6VcA76yyUlleessbfpD4drlI4cZbftRZWhkzPi2YiITWPKdYkzy7fNPTdGgaPjQuo6yr/
mpaznFIb6jQnX9IwC7q8fX0PEVVwZkGyl9U1qWHnFQcvaTTDmutXQD/XESinMQ0liL6+iPPA+yRa
Utt0ol9rV3/7Ofnc/2rjkH0LNNR+8NTlPo5sGPVkHGKNHVxwZdQhPqYHfoMfHeIYqy+9ylVz7Jrb
styAR4ZcvHK75GuH8q+rSVqNHCkMF3nuBcc4hR/yIf6mmELCbPb6DvTEmHP/KH3plnebzdfvM6NH
ka2jUkwzfrdtUQpDNRdibyiPHAq1SLYbuCFjv0oRFopIuVkn6YRUHn9Y1nirKXtLFEf4IrkSA0eA
BIEuvzQa+4y6bYjPG6qBa2ZoOQFfv7gUCBEByJ/W/aKYuYKNj7/K6Oj7MU/oVKZXwAEVjGg2HxHO
CHfCiQjXn2XYyJI2Lujhb+0Gw1AT9ex8C7e6rIySrUSN4SR9URqPgg3LPnYUnGc0pwnP+/lGpcoX
huNfv6YZqcgIQPXsmYoobAPjN+rUuMkZ7coyyPWdKMCoydVqaEbvmkOl1VKTmQcXe29jwN80BcQr
J3Cw/BtknA2JtBYaiE6Rb0/FN9V8N6s58duRbu5lVpAnTOvXjfmPr1JykuJgAc3kgz+atE6DLICa
hISTmFv7AFW/DwDjKsWiI2Zg4SZeMfkikm6hn+/bgSUSgj+667XmCR6CykIGoZSNb2hWDJsKf/Su
XKGKWePThkQ+IJcGTIOt2ivylhoiCQ0Ld36IhMKgpfQ0gOwEuLQ0UY0MqHwytQpaMc21hhfNmWFS
KWNKc+ra05dIXqu1usVp+CV0JRyBEkSWiVSh+hr72v5LJFBSUdhAsymJAf2om9ibwtjAKCvvrZ8z
EWQ0EXh9ZLWRdDqo0w6BKkhWCrHH230Y+OO2LFHEc30DZIXB+ckRDjmBCtQOncJcMT3mUOhpg2bC
yOVme6XYAqCwrUzZNAbbSrvcPDQGn9ukXwzIDxMS0YF54xLDr35VG9qUH0bC6FNN3/kOlkFLd1Ys
T61rt7ilbg/Rl8GugGerr1DSVMcNTNOE3nhe2575QlUfzXAE6rGu15xXh35LfDWrSVcFQIEKDNjV
tb4EfnQ9hHsxFMd6bki24Ui0rNAOOLM4asZKR9eCx5c+0BC24bvENJX01MyYo6Nc7CABYAIyoALh
SXRhLtb8LrpDCLmwn7X6AsKoN+UuFCr3j5F9sUIROpiSpYLZSoiDRDw8myuQ9veXYHC9C482bTPo
gnxSi0YSGifeu/alfe5CawKrm3Ax+AcZOrYO5l0ylH2DVJufWwykjJirsgVW4MQGv2LcZd8btelF
47r7GTllSa6KNV8Z2ie4iLIyl+PcFr26s4eX2oYhl4Y67a2kFRySGpmL2Ghs4EG3CCc5cx7cF1h3
RvwPpUUDqJqor3oS6m3DMOZJHeRAw8m5F88OKhc59HQQoafWPGqIMMoggOOPaGEt4QXid7o1U9mV
8UPkO4F2vn9W2ImYAEZx5GcXvM/xVnCp4LKJ/+HjKuerxg6wiw0yzTvursHKSXTFoZ0dT8UTJm7F
ZsLPuVUERIlEtblNMYt/Z3WhSslOIsJOJis8XnFJj+EC8ON+R1qDc/78u+isUqr5EfCib/Avv3+w
dRG97DZMfUFYBHKSrTyTOuR+IAHnRKRkCt2lwS0b1LzVihHbBgEKt4RYR/vBmE+58sBXyr+B7lJ9
CWlQUD64rkQuB1sDzqfPcfJtxpj6aX+YSJjBoR6zDPuKfTxibpBQllDAB9bBXIBIRDEhGw63rZrQ
Q+2jl5YTywWeXxleCRhDjQdKLadC203WfIYcP9Q40z6YeYvwoyRWNJXbQtXZdVyUeKaJWDXvySrY
qnF2Ahxk44LrRi3huw2j/tqO+Z7dAYNTGsslSM3dtlpLzqWTrVSMhW6P82yp7JlQRK00Rh+mZvMM
gLg7/aYsYCA1IcvldQeoS3t+ZM+eVJfeHkWwRvek8BjamP4mQQpJCzFrMICRju57JThgRjXFuEIz
kODGO7gM5fIqfU+hDkvPGfGN+In6JhkiSYnv6Zb5bB8SSUBx2qCsNEJegavZW/B4Ci5FvTQpN5r7
Zpv9RQvztk6J6FmRVh041+dbJs62LtguExkMRxj1SX1ndVkhPWRR1Bx35lKnJ2sZ69H+HU7EGOWD
co+IP3OfBZaUkdQtlsb5mTrqv8aOWSoK8Dkcihiuvo4NCl2152LUNDS8jbjjn6IcwJFKLJAdChsG
l1uSo+tCb0cc92QZu9FW4uXBwgfK4dBOUrMGpSVL7hQyzO0kRE2XqitiklGgQ30qJTvuMwej/4qD
l+Vz2kfIGfMfLB8bCAh8MbyKIAJvbkOBee7yvWV0Pw7TsG9P4Yq+cIiqVq68BvZ/H2MinVTZYWyV
J3pU2cq0OKRsE6Tbc26yhfK0VsFnA+9W4aeANinDWSq+GpvVq1GgIaj+5vH8fbuIzysPLJpDzIJ5
mDPIdp0kl/ZA53d+PByxy0Fm7ddvxFFqCEZmRE3xfpU3EmjN/01ApjFcDEET/BA+6x9wo6kTLTsD
v1+tcHW0ZUvPNNvubG509cUZW3axAWKSi/grUMR1NLMnaPomjAbtR5M6UFhF8/RVN2RDJiGK9n9i
k+jpS5uQGFV+h+88icAnuAeEtpQf0NxL1dL/HKyAwFgGf+HQLqVVNLELOuTmdAR8T1UbxYcvVzk6
0AgDsrFnVnB2igHz20/N6CzCZd3WQ+W1Gi//7y9fZDMld5HbZK512LSz8v6XRGGGBzD3QtG9nz4u
5w4IgV1e1LWejJKz0z04TEofBnArar2XW+LelJPDOoyB0QK6JTo1TO3ol6Kz0Weo3zRH8cnu2W5n
toO3qJ+V8le5bBhlJqySOUgSms2N+t+pnuYsJ2oXp7a0VkpW/b7wHE00AjGb9QlxGhqtEDlloV2J
tNCDyO2UxHRwyd9PsiWEWM9AP6G9pQZQu4H/vJLdnWzWdGt+4nfk/Ioj9o0NFGnyty0gYET4Hj6C
BMfFu6umQ40pOCZf1Vm6TJOThdZkfykIcHvs8k+RJ01j+kwMjfF0vcoXrT/vxiXjcUUF2C7YTf8J
NHFHZXHf+hl5gVs3/er5n7mz78LldmL/ToeMlQG6Z4N5cjRw2w20cZOJQNiYSiqUgZtdm6wTutoa
Qh1Si31/XUK5tZKa2fmJcVliryL7SMGqKB8Sr77HKL/K53iguMUd1Z6RtgNy07YtH9edhJnMyg5f
mmbfI2UPtq8KIXmJX0NEmh4JsPjnZmGHhsYGczgse+adZr0bcgz+BkfgbHGUp0NZ9FOPJvkEXMtK
59UcWdtuHgKTsQMRMRlNbJHNAbuNo7IA5IQaQsJ+mZ/jihM5Ua8x/fSRHSZn0jEpDewMQ34FEQbk
TcB8co3HPqIJ3K4q2AkpB9bPrUHRLbw+Bo5z9VcbvVoUPixB4xA4evi2gXAz3njQ4qtTmz6CaUs6
VRhvJRFwHeP/uDkutn1hUkyhSdcOT0sg6Xf/cmvBGhV5VgfpbJ4LcJ/htgF5k9nIy4MImhtkdjLi
80ixlsbiLq1OfZBH+iVvZyQFTYK6LtU4KImRSdMPBCUEDUTeTVsWkzVlfAqJgJY2h8OW4ylaPBov
upYY98BoJjbWeRAzWF0ZmhLXvotht8k5GDc+Jol2nDWI2HcroUax85fwd949TRzMw6pThvZQXZ5k
ve4x2GPv/Q0RCBRQd4IJJM8qG2yLZLFy0gOxVCkoSemmtISxRLJnd7jD16ZQYnJw7+8tJac4/OSF
B6TEmjsi9O9V4qHwb+aBkGnDNEIVDGOh5Kjf0VUfiqSODY5sy9CSh95mlmrx/vfKQqLJKPrl9e/B
56ABFdIW7bskrfJnriN4cbwJdNIKWg6HinvIx1tYHURHM9GO794zFHIK2V4ETkPm9oQSVSWT/2kg
1h8gUEGxcoSQFvFPVk+PPTJPABIi+ZUTnm0wYmVSuU31FVf8DtUzbCr0fV/4anZs/Wsn2Vbm+3oU
L5fELA0Xdii+57vdm/HyUMYV4L0D3t2ajF28G/uQTRZ+NTg71aykFaUG/8VFTU6OS9LbN2KNvOD0
+JQquXcOYYgJREmANnNH/P6uzJXtYhbQjbm4SC0YtyTZ6sVoU5fDk18LXLwqMMA0TvaDUwYrwtSt
iGqaqnPrA6/6bwNPr1/Vg73a7Dt2Tx4EsPFQi369w7mXJXoK3J3d3LVDMTM7RkIb4CRkj4QvftaT
D69rE0iH6/anQft3o4GQQPuarvgUeE6RujC7lVwpzaiKQPcd1vMOzNOg/Et5uW9DlNuPBkLe9j0M
dOeFrUYfEjK3BwkV9xi+ZtTTHjbdpY7v9+m9eZ8J79M+1n7caA8buVlU8J03KAQ+COnDVV5HUe+9
Sh/4POVpN3xfGeUcUoldADFhL3I3m7wydp5r79/iXQPVVa8x2Hy+YThLo4a98qWt/+L6OHBLFO6k
4TP0H99VSPrnmXno3pLCtlBAGJAd5cuHNJeJ2Z35rJjtYjojKb+Sli9XJGQJqOb0GdpGHfF43AlV
nD696PnJULmucGL4umsHBz/vDzQJ3t2nEMQqYU2czfFtgDZ3vnsLEEuGGZgI8L9Mb0S/Yl4XC3U5
/TJXCMUJ52QTb2sNH1LEP1jtO6H4U7PbrJyK/QKH40Crz/qQQINtMJE/Z8xza8yytbzlK0wxq1sp
rM4KXr1dkOrMUmwz4lHLRbQn8b/nlw5xS7GiGDdegIAhVxs5hiU5dimQGvLFLuYLNP6WhrQZ5vU2
ODxCKXTGRzvxsI2buKyF3kPqYkCpX7TIN7STNN5771fTw3wOUIS4GqUFsUc5GEsei6Kyqyrj+TFi
9+Ni0UkTKn84Q9bs7pfuya2gFNBVlE7CcDS6USCmGGaCbz2s6KI5e81p1XOjXj709orA2JAeIoQy
TZxnLpbYUvmIAz6eorZaCK00HhPl9wxEzNF949X+eLF9iv5ZJ3b4KhAiu/hv2AVwWYwQbMe1FRUC
0+rK4779xmanR2jSuU3dNbeRo6TBqdccbwDkEuNsieBzeH5BFwC31Xh70ve6ArW5h5Ch72HAVALm
h87IkuxrqPszIu9De6AA4LO+1Yx6+qEQINjWpcWBZVEmJ94eVnE+AwwW80nhnkwclj2wMEpT+7Bt
30JjLnRJD6rp24ZzknJzYET6qNyJ1ay+SGB2zbfG8dkSDnyHJg/UMwVKZiNves198H+5Bb46XTW4
dOquIUdj9BlD0zMzDiEum2Wbtg8g9pFD3O8QmRPOVxkEea0o3VV5b0gGhUq9DZ8u4XMfrzUuAU9u
GbmRye9cz8IVt5POEoA/dvf9vXKPVbqmfBxjRKe5KxDFh1k6rNgiH7mRutp1KbBfZR2T35FDBocW
3S1aMUgULB6Ie4qkNvOvIy8RBKuzY3tO2Q69HdlgEa+GUAatumWFOSoqLrZlJkDRDEIwywrcN8uX
jkF4JJTP4LKyhfkDegUJURQVuHVBv8krI4gROuRgEHY9EzXra+lISq816UdGUqic6DOEK0/e42Ug
v+HJn5GQO1LGKOBbk/+8dsC0dqHAwccDu0HkOKF4swnV6IASEvcMGLDtYcGzFPAeayHLqpXGgpE1
JQgERpCuOgi/Nrb9fGsvzHe4sSMsU3mmdhk2ScYZRE9m/pIupagJXXqFrgRg+7DAzGHwFSHVTdTy
EK1PgHqwYXfc7RYFuXGVc/LAOrLP/Lp7cfkE97gOzf4pnHR954FrObH3Vy90gD4cSWtesk5Ufihh
wLaVVvDKxFXVZwKW8Nn2saVBRthqNQtkcBcUgm0WOxb3PjOelxl+k/BOpOLlwNMZvjRPlel5aTbo
6FQJHRqO9elA16LXfQv7AEdkE9p3W4G0ez+OROOne1R4xFMGsGLeAQdHPONpPcXGQfM35gE9EklK
xokiSTsuccAsYcJuZk4U/CxYtsd3E5ZWweyfzW/ORw/DHyGI8kfJ5CuMC9j1AWNhXqOcA7HhGOto
DyJkVLkFhq8wiKSLveGRN610f56ldYoVpmNtuTmsYKJuyBYuJqv9zi17VEWKHDYc5RpktHSB7GEw
x2CwrUWGSY+ASEYN4O2R3IqqJkJbSnt6gohenKvLRAeGxPBO1luCQY9NN0aEBNFtZHRGtIGcU2TI
qpbzIqB6PaIcPYaidOE1vg+zL4kM42JpDK6C9ByH0xMdgTtm9WIQqSfcmuodNDL5qQAtl2GsTfH3
gPMhuasjf9ncmNJ2htSNNRj6mfvIi1dJB5sqANKnPmW8yIwP4INoqbdTNVX9tTnySIM+EDdtiykg
70XRqmvUqOHQWQoYNUlWCEdMeupEcqhJQDQ0/2Pmgce01BhMk5wsMVyFNnvBjkW+F/OC9+QT5MGn
FVPz5iD6ZduuEQOwJoedg1B9PEt4o6KvWXHZtRoajoF/MpRB057kYFeztRskGGJkERNlWD0L4Z9C
twW5A0cQ96Emin+NfXRRmWVBgWBaGLywII99xTDArl6KAVnV5ov9ks9izFDDdL4FqGlrNV5pQQJz
DPToNd0ndXfQS8+lYYWcMXZnpd7Qf0W8FXVf8tiDemdJJOlRadIq/EpMI2UUCYdN7s3b5z4pak9X
tJNOv0fIZn2BVJu5bJTdOwjTXNTTNl3tuA0aWC0/+IxM04gufPadIwV6+VDmXPHhSeSFGyX7JqjK
9/8Bwm000DVhL1WMUTdBnpLSuXct6yHwjHDOBTQsU4uVLAC0Bg/Uj0Vg/uIotpsSvrA0fkv4PaRo
wXeKnhmGIyZW4r1lsN1sOXAP5t92FhYWOrnUOlrzSu6nAbB2bzJyiHIotCR+gA7YmyXmZ+0Grp3l
GsKPnbRaJEyl20lBKHz3ffPzwrEQ0Q/OOi2K/2jIAGtpUUsw31pDMAxUOMAwV5oisgvp4Nf38tQn
b6LILMTq0UNqDkQ5NJ8oXwoFMYx3PjMyNU6bCCCn6I7PTky8pLBRaR0dLNF2hQgWsyeeg/n8a5WN
Bw/YpwoV/yHcScVxImMPGtKxABGo7kiN4TTZ5Z9DomDVRcOaB9F48NQa2lSm7S4Z3v6eevNRr/Hz
ABrgDx69UyunOZLpVaJuJ0gEebmidHP7A4a42X9ddTHgfIqWJWeHYkKFogs/zKKFkds+LA8VYU6K
mJLZJeEiXokj1WnMBcnzJfpA6+/nR40RJCfOgXuRqMLu8Oy7NoS39ufLr9heH2sbwc617TJjyieZ
4ZcvrDWNY1KO1NHesiiDukfZRzslDMC9ESrTTfbbbT3QyuyD3LcR453JGO06sp68PgtPA9OGI33/
48FnL0DQB2+zo1mJyVyWiAUK+bTF9xIB+ySb6BzVVBJR4TZClzqXf3wwcMq3bgmUMJwfzCIglnvb
QLAy/heZle9tIn4IebrzMnaG9/U9EwPRkGLqwUzeYhZZxCJUAISK+qO4xZTS4u/HJV3UOYA5j3Q/
CuDJ/6PwYFSiJVGn6bA4Y3kSKMGkGlmcvGYSucKJu6sA4iY/lrPwsD8RuKZ4JO3cJ7yxhIDVgvse
N6peZ8jFDwi8dRHNWyRRLTJEtoLXyy8egEuMaPZcp4EwA7nH3DrzWnZJuoDZUd//BfhMhipqztx+
aQm+/ytuj9w7VSdVY7xnTVDjETWHCZTMkOHjwUHT5Fv4jmt1gubZdyZzN+Vk+JOldltqv6FLKo0A
bVXNqAmGTef69Q8PR2Xrdof1rQxxcsocuXLnia5MAOnOJS/trbEnUxXj/7WL7jHLxFk2/p+oDTZh
W6RLid8KtgixcS41d0vy1AEiDmVrrNaOE1SwI9uh79WPMHDH0IgXLFRg1kS77np3yzSq3H/4phQT
aVa+yYS51KXK8oZEu5DJK2VkK5e8IvOO+t+52XlNc1o69/GIVY3GHQK1XuDrMqkTJGR5lyiqNjJR
wd4cAMd/KnBqvOY9Z/vUXaY6kLAadoR4P+tiidaUeE00h61FvRmF7ErQ7y6kDFnsrrSEuhZNil21
ESUC3OiAWzxnxUxUE5nIPZo7aZ0nonQWH3KqcyLOzIoZ9rH+gdV52kRmj8cXm6ylqA6/MlyEqxrV
qWFEKOaX74xQ14euf+McdE9RnPrakWXLMvA0qQXn5Ux45wj4d6baGZH3RsDrOJRh3y7P241BKnaQ
76Oae+BOyjRm1f5QEyxViXLGCD+y3a6+eHEIq90sBQIX0e3mTTypAdgRfgwuhmK0I61eQDcCAJPT
TiNBRARhZAMy7VgbeSOeYUYrKbcMwBuqnuY81yVb7847gecNZnDH9zTvhgWnFjRkJO0LTmwY7mOg
9qujWE1akz5+y/1X7r0Zkj66Z3mJj4fvtY1Ks1+TN4KE/R6JvZ/+v1pyWzUJdxv77/FORetaEe1h
gFBhmEAVYaNXYzT0dnM7g4lnLLH/hKFhyRCqq0oi8mc6Y8YkPWUppJ2cqjxkAm894N7SpKiSlrsq
M/OxZgqFyOKth+/vmRc2SphejE9PCm9DEQUYzlgzF+ncrY3NYAlhfxukvgu/Je8Gomgu8pAYX78Y
b61cJpafokvu9wiTl7qs/gqZd4Jm7W2GvUn6bhOVS9z+AUsqdr5Lj861mKnyWTxn2o353CZb5muN
EWqY0azaNxmXmEjnFbzHFUtqw10mOLF++GPoVn9vYpFFPFBhr8fKQQVD/d5JZz8kcrogdU0/1fyq
bCKzUYVaWSD7zrtkK2zGJTM4+r8Cu+XfY85GBdwNv/FjyPdvYYr0y/qbdrPSPLNkplRZ2c5/HXbK
X0Ud52buubrB2PrVITtmLKle0PbURw11BYNTlbdE/ME8b24KaWkVl8yzcqbXwyj5x2gD+ZvYREpm
qnYUyyeB8+5/UNh8fP4N8Dpaow8ujCgw9vmBcEI5b59QGxFNBxyqkQrHkEyOyQCNHRs0Ikn4x+0c
f30vxvNBwEbdUu+xdjaEZ2mRwTHg4ZbcHYnNRw77P2Co6TiHcCaBC2ygX+nyaGB3Lweu0W/4e6eq
9dkUK+g0YOSyEeIW4+FryThxE2UM1nY7YRCGfs7efukEBddnRVQstDZx3IcpVJFBL2ZNf+3NzBcF
Wo2OOHanbSqz3Q2K/94M9TYArd0hqlnrsGBM8cDoiJMJTBKTlgdY5IIorPFUxBd97gQtqqR0zubh
GqSaMUh5fsM9Dik9mcE0dxjuZq+ziZxHL3mT3cY2M6KhVTyjRY1kh3o/bn4oJ0aARoQGUiU56rtv
o8JQu/O810xgFWQLg7hr7q6rdBxstds+70B+hK4yWYCfHEZ+OaaNlD+o14dTRafujAusIQvsNk4Z
QPMzx55NFkQRAzC+IOOI6slhI4g6DNzlSh1OORdfApl7Jn//BIclqXbZZ7hFErM4anSwBTlhdszk
1qYq82XZg9F5LQAk9gLHbi/SjuRTTrjgTM7KDUCqZpg8UhBdqS9/aNXxHuznWtAzKtgnATO2HUSS
l9sgtR5rH58sBNwYjFO6Xe0AkdliMF8CfzeVL6hsFqzZfRDTvtfSUzhH3fsduoR5kFjlbgYDTPyZ
WiyfluolatfQcjEnvKHnfauEw+fsCVmvsceaOJM78w/fji0OSzcWhHXyqfdaOP/zeO5QHIZaOCLW
BkmsgRy/mYDqJCSxKC/zFsewE9lgCzKgMh4psQ4wkhMgUysGgGjRIQpMUjs9Iah/xs29fGBH4afB
8O0ICiyjRktkehkqRHa8TyXKQoSf1yvBI4rHkNXdCp2Z08XrVgJIGU9WZKc6g9r1ZKFqsm8wgwxC
A5noYTxG6xi0mmmGK/wBvV0zQVrTygxbQkU6AbGgq+6sss1Ly+eeelE/uLCyIudYzqJ4GS4Byp5F
F0Boe5j5vnOmZBwP408bpa8+Mq+7LoUpHVaL1T7LDNYcfrOwh4mKeLoF6IDPRKEy1GpMiSTlGTkw
bFODr1nVPOoxG9kWsIfj04MPTmQbg4+AFHbEZOqBIHFEfK3jsxF6bVPzMDC0aH+OopBS9lgwvYq7
i53cZ08PoDRcF5zlzjClbGKBbX7V8B20f99P7muMN4mW1IiFgoWv6lMRGdg3vdSCPADiNCuT4T2D
AITq9sJN2m7Ri0TA1yeLQQez0xcwZx20bvjq3QHXmbflajKjEtKfrF2CJDLCuADQ+7fAtl1HjcS4
Z3uX/eBA3vCwYGVxbgyAF5zE0L1wjXNyMwCBM6lwtL+UunLqa9KHTCr7Zowz8n/NLaTcrlQdiKfv
hKhEaOLFs8HB03xSMKLHPXEecVtuBU/Kl3JuhR88OdHZj+N70FJKCKQVPaH6YrRanas6aQRN73CK
M7frn3Z1kdXhqJVVLObV/+8HlNrq0H83+bUgu08WKpcoOHMoSCwBIrgEsIihSjLm+6HRau/oPJx5
VPj14NpUeCMIVGibJgOb1jQ/hZxxU58Gfs99F+fAWOsy3xzzmUMUsP5EASFHqdSO73NVF1pKxt9H
SeXrO5OXzc5n0abhOHpOwrFmiZ5ZcyKJ/NavTafITBh9NNlq3zFlZD2KLZRIk6o+uEmKFjd0Ljq1
ZdYHGYdjNqrmfYROYWw/hrRyr/e37dg8nrQgI4JIlTN523oxY/wO5fZX2hjtyvg3hlPVVNJzbByl
AWjXu6dFYkmtIRq1DJwTtR1lWd8upgNWApomYLd1u2XpJOfZmVmnnVV14sCzcd7KHwxfZrNsQ0y7
s6c7iKBLr6qPaKwD8fOd0fKqOA6u12/mar7Vucg87Imvxmp9p/FznI3JmkRqQupsdVMXMpD6Fblb
xEguL5/dhQGVnXKYA25buC6vVukTl/HI98KmqqyPYrrEfvmoGib8fSRpsaYSXxKn8YALnAJcxXi7
2SqrGiklo0jlJtLD0rShwcnrVOXkJfsU6+0L+xtFs/2PvnllRfn6rp74Dwe6ybGrSD0u3XWCqpFh
HHVJ4ahJgosiQYvAwhWtRk/gsIDdS+lAu4UxPAZTlTK1ByRzEnqR1u2ASecBYCBBphwk6yN4YDG6
3Gw2gCRmPjnfg1a/kIV4HRsWfRCnEri/+NgFkujzCvmJQ1v8ThqeUrIs/f9j6Bwrg4BTvPyVRJ9V
S9PGZI2rxt652QQSTnGjTVqG3msEz9C8t8GXIJlIbudQqiy+yTlotGnpG2te0k8QReYQnNmodcws
bHMNgwy/4GuH2CTv2zbSuDkBgQXc7HpLwqTPNwyiq2HUlEI8pBeN6w/ENezOkCGAJrr+k8gDhVnJ
1ahDVYJfDXwPkQKayMefOO0Lsw/d6N8zroi2HPmect7NlklwkOmtISQzTnfLXuTZiK075DYoBbu4
yEETQpJUZJejME9A/tc005rwFKZagSRPzHnj2A1rN17axniYweu98NzsWQv807ovpvPj9H4Lzsic
4JBjr1IUxPWdPWjUkGsTGKTA9MDLJj51Qp3p7XExoB3iXo0VroUP/yEQpkisBqztTQSjWtIWCMJE
M1jmaDiYDeT1dxc+PPbPCmkTMM4GBvcl028tctekeHXDSToa5/wDyXB57MSKOVaq0mnJ3bmXaCKx
Q97fuAG0KG9LQrDq5m9dqnlZK6YgZ25I9Iu+CKbFBdNOm3Wx2ahR9aauKNhKByQXbExVWxKUXFEB
SGuRPp2c9sqhTBc92Bn+gxO5wngHTYSzq8uGD0WsObLpXO7mILvx5UGNcWKNx3xMyyFbJmkfShCs
HkgUsZvKwznt0ZhZLoXW4mbJWxLdRTZ6i/TXkn/o9BWahxSNxAD6eO+8bd3pc0s6BOy12TkAbOaK
Mx8N4dI+g0DcmY9GAPCxilqr/5wdPWIMAQdfWU1VO95gPNYqjL6YvoWNVnHSTc8W6H9Q5BACWDIk
hEBcMxEqrrYKLClAgvpexp9ZSNn228baEAB6WRgp5EPxdLG712aqfQhCZHmgUFfgl0sAePui3y01
V50y8mfsNsahFByRhDdxW5CkA7zvOvyH3rz+1wnVnEO9YcDLQ6qYNLwNNVenBRtoj77zYXBMZ6jL
GN+4kpAQhFxM3p2YzNOoPgghrJHTntjn8U1FmUQJdVqtjf5i4vo7WjRRLHViLXyUiXj+0WMxzR3A
pcjTqgmEkPm6OBxKmyxxQVMm4tZoSxeB0Lj+snipN2OYz+m/p96jsbzpqd49Fyiq8d/HoTllnzH2
sZSrjRhLoAY8pDpFhng9dD9ms49FlJWZwScPdr6Jqh5p5XgSqOLKn1UqXUeBKrYAHQyvoTeDIMcB
M26cYiLwCrZSlKMu6U8ZMyBXKrU1KylvIjFIcmlo+EYXF6d8qmkkc10ZcDqE8dZLQQjF1gBTDD50
rQFrH+GA1Gh5cH1Zl5lOBzhI76YaEdCRPX7J7rd5J44QBFtG9AFfvDj4qSojZH6jTTE8+PNFJyih
/XtEHb7Pw+M45kjQeN3YNiT4qcqzqOnZoWgyJ8wKbls0KQwK6VxMUBcruRRSQoquu+hsw5Cka3GI
JQ7pxc2FsZEIChKXzfaiB/HJyKelK9FK15JUOHYY2CxqXa4xyMgn3zCkzB4xUViktYGl0KayToQ8
gaOcCFSG0nKTCvlL/ag/upXc/KeiNenPmnSzrCkVvHxhg24mTspMdiheTnU01LXastkEF2yBYJa7
nDSTDEgJfEp8imgZ9pkdJk6Vk9/LxnXGJvMH1WXeibYYSlKWtxgQsVpYQsBFp4+NMi0MFdJJYwRQ
J3i4w6ZF7I9QyiqUgCHpHTwDETqL8a36BegPh50C0WnZ97XFaC5ls4kZg7fOLsjrvMuRbEuZFME9
rMf+if/mjMSL10Uzhzb3AZUp+G7dcCsNz4cECZxH30Vg0XorqSnlf6eaAoK8c0q1iSq9iZld4AM1
SuRI68BxPYbfSFPor6Ib7C+QeVpTklfRsjmxO5ln1KhmDh9bGBVo74gPxvLzwmS8nNdG+sxQ88cW
w7J1KRLS2fviPvG2rOIdJKr74guhAd6nfHn2BnYT5xcWX3xwP2Axmk7HvSozlG9YWMVovk3g5wJk
kP/novO5ISh9tGxYXCNnEOYzcIoCJO9jBKe60jBAJVA2DX57x7VWAnE+VcHthiKnzt5+5Uh07uf5
+r4wHjdJbewxlhiu9huGaJ3RHnHqhAXAQgSyC9laqrUo2hgrW7gUXyBTIP012l3zBRgVpayBgh+G
hyB5IH8iuwWaF+hJPIAi0BrwWjEb5ESBiKtedNLBAxGADTWHV7JgSKg3yhB57z7qOSlvRa6X//80
Oj13/8cdPpuF8HiivTCGtJdhtweF7xvdRidUQ31rWDG2RiZxFv3Jn0x4W6en6MIJlev2n2Owr4XQ
CNqPm/z1MZa/Nh1uaXJYE0p+7J38Cpgngze8M85rMXtapWszDhMlJFyCGH6IGx/K+27uvVxUCgUz
0geBZ1zzckBHheZ75uFTNNYuLP8lhAOVIp+qZ4XYbpXLv29l7/tuxZZIiqbY54gAcPbqDzk26sfw
nNv68b/YfDz0sWdsrEWp5hNHdtziOu0/W6vO3MpZ9tMaSl82fs+xlzSsYYOLGq+JBwg2XwsTvaum
Y7oK3am5x13LrmptDunvCAwZ7XAEzDCS8K938Lu9S/upPOYP7IFohDwAOTcE1Z0kxXwW3qmh1dxN
S1LYoesdo/LbY/aTjZZX1lehbIjxI1/YHwytjN3xfIWaEA5wYOG/xdh4rSG/CZxzO/PAbJQYQPUy
aj/zvbxjEBy8BAMBo8MVO18gV3WEHkIr5CnV//skln0Z/I+dTjGM/WkHi8V1iQ4lcWx2N5EBsh70
WUN/OzAH7DIi/g2miHvEfrJLyJWvulxNgn97ewSgx3C78UHozGscBVczvwz1jkoXJ3X0fjaIfamt
/J2lOEC0vgQgeCkrq5vygC+Chkm54m/aenJO3gulBdvhwX5jDS4XZfO6KeRPKOVU+ZaG/tbMRGkj
sOOr1ayTL+mdHCjgzdK/geZDlXG8qQEFzMWgmkvJLK7OteKbwn4OcY4/em3nOcnawqg94AfbbfXX
vgfEKD3tjob6lKkZ6lwZTh+J3sFcY+j8FaDdp8CK6xOc46ZgSlaAJSbkkljxb5uYZIovWQnY7nud
st7OyEzvKP1IW9FxtOfAAG72p8FP+5Io/Vp3MuU6dXPYeIPG2zCmbVtXeMYSZm+xLXO8HLxU7H58
pY25RI497uOCGgFW3SHZL5/G64cpTWyI6gyCUt6M9GJo3/kOiQmjnO3+A5XPaqlHLQHZ41cG083q
KlK9yjnXmQT1uavx795Hy2tZQrpwB3PtmY1dC6JKOsT6E9mNZ8xi/jATQkvTrOi18dXo7sMamTDS
5vA1Jv9xrsqq1EZ0D3QGEM98VnBj1zSy52RRyeugu2f3mBhaNB2FCRLh7AVVIT3Dk5eLSrIXyDXV
i8HHjxLyhiru5bNeybLDUsyEhgjNWvKAmLL7xYCOY6etiLbAU2/HIB6BYTDe4c56H92k6vORUYIQ
qww7A89X1YdgWa6zxNYa3u2Kqbp7NsZlNu86ywVCE9UkzdHcGgd70KKzqGKK4C30vD5Bf/1j+8Ub
xHe7wQI/YroKaY5PpIRAHgjAO5XWQs/whe4sScwVeqIhw0Ma6A6GK2TjtzVx783W26SWe50iVLsJ
2wAUwju0/YrVRhmoBbUp5+OJVHTXJezRMec+4Tgo7FmOTDTQWLQeJhPHSxv93tkqaclSecdNdJ9l
ZqvOImMylAatt7KvO6+8Gghgr00wLuhkHZ7ttB3P/E4wrC4bPgzRNmvMuSdCmL13efCPDCvV9YxZ
Mc3MKqA2G0R+qpzxQi89gkfBtlToqwiY/fxNhbEj8DG1nPleWf58fl/4us2MUVKlggB57N+k4lGJ
xjfn23Gjli7rKYy2IsnHpG8mR9OJuCJSCMyMnU9CVtsk3tXOOqzpM0KrM/NWVQiVzaAKyBA4693S
oBNGwyycMurjhsYbNiIw6aT61N0ft6yZjOIxQa7h/1G01rOBuZQSdGUqcxMqbkhrTgGaTNKlZQwV
XzArM/GBD29m8h4x+QZDEjdiPcibZYISvA5SW7dMPH1UmCcO/SLxKoi3tc+zqjZEchHk/meODINw
PP+7eSYTjFdndzlEvPJ0gcnGxzbGYW6IMyXK0aagTECEFbUS8dc7m+IZeXsGJ75orQGHxHevcdAT
HICnkXowCep1w4qve/AnjF0oHXWd3zOK+YVKe+ANAKUvi6zuAe1dbP6svr964FE003zY/4aO0m2U
ABWXnrdTSnL54ZlZapJgzfH+K/PO9gsTZ21UWF682mnUwk0Lua5Mtsg3U721XAbVUz61p5fTEnvZ
+L/tpUPE1nd/3XAZUsd9E5kBhTRLtvgHCfIYGRAo9jMtpfAAr+yCApl11wpj6TjT/DsHYvrBif0J
rOGcOjL6EpBaZc5AERhGp45YYUjmCWw45bmNC2g7oi/JhJD4gK0YVzUlgmcD3zpF6yumJ8HJWcJd
hsOUh4Rg2vcp1PiL9hgs8W2GX6mAVMd6dCEOtYTzExWYaKuy4fhrt0JHlUmUAc3jMnlylDKTQ6PC
Bp+DlKlVhZFkbfSL87vvo5Lp7cOEA5Ax3S7DGXjurmB+HXVHl0PV5y1Pdp+lKmeGU9fe464a1FsW
Ij0P61nJi5vG4Uu47ztSYQQf2pJUq6WAZCAiLCK2t48hziw7p+oT0Vy+hQTBx4N2YYXy9RbHvSAM
LefnfXgsvnhwkNsEZgdEjR9EzNkWZGDdvAXJK216lZxvG8kGhr4thTCKlBgP29F2DH6NzA4/72oe
hnnFO6ZpkF0NYBFJivu1X9GEVTR4beCsirqufjYN5cQnbepXV7yxom/OmeDG6apP8rT7o0WQT2Zc
rOtSpglFivJTZmSBErvVfsnOcshewAUZqOvyBlB+cZD7It23aUXxfdh0um/pN6eEedSs5LfZe0Ll
RKJXprHOa4i6CTeI/MPe65DAW6Q8rYJ1qYhQoR8FsNwPpHZYz/i6PtuGm2g0Fbg3kNDXYlRP/l3C
KY5oxwQzJ06pimPZLcGlV9KioTSnY8VqDFtWx+NFdnbdu/x2Tblpp1UZdeXSbbvii75mCw1jHof8
mylW3HTfWy80Kmhi7LzsPW0//BW+vYZoHo50WVfL0olF180Zee4YscYXzpvQIamE52OhfKr/G3qv
ISuLNCQqd70DN7Op46mFeITfQBTl4s1H1WlHrkNuKeBID+c9LapDZbCenwUA77Nn83nayhVQ+HpQ
L+ikHexwiaIa3z9L0rPB+shfffL912ZYzQltIuIfacdPBSyNxLth0oBuMGUYo8y+ECvP4qnjovFy
YDjmlIBVHzcbDJVmOGiF/tHBaPrk3xUnwixe4jTogrDMiNxMDsP/RAgycpNb7XwkOu33s27h7Z7f
JAA3l/b9R3pxpzHkwHTfawrXdR4+O6ssfBiD/HvwtXYAeDAeNIOKZMVdy8hYwP3lfQ5Da+ko/Zt3
rWX43fA9auwCz6KLq45dPvknmaCHZJf28K6aqauXPr5WcbGHrhG5KeLbJxffwokQ6d/rfo8+UQ+G
j4fnEG79FktIN/oJu3/U7/rSynERj+rv95YQkOFfTVflJuecw1RnLQ3TiGCnMOOq7TcHHoC802YD
DLnDAuIPGV0ApcqO9fPEO4r7TF38Nq7P94QPMplzC7Kc0VoRJ8Mhqd/ty463fY4+gZTL7cYxW/QO
Efj+QdkOun60SpR6sgUkDda/JSOmhcCXwr83kcMBBB1XC/enHeca/27/rZTzBUCjFL3g84cIN9Z1
fgUHu7HJFc3jNZ2/pfAnoJ4SXwEokhyUqZqU0LMBRYlKL8kVgUa4xylFDDs7HP7450lcuh7MG+h7
Wohv2nWJY1rHF4QN2gsN5R4wlMUDp2aHKFfNHrFUG2ZQ6NtKPTqA9zvfSK7UNELNPj4gThgN1ZJp
yrqtGJaiRYX+E0AbtsSD6CjOI2dheRO62SASL3CRxnSlZyZr6VgbubamgXsicVxYt6TRThugcFlA
qSY87spPbrc/py60u8VsDZx/SmpIro/cLBhDmL8GVUS8br565pHBsl+3Rt4/egaqc4I1bC8d6Bkv
L9ifp/av1aZbcHO8QZIMDn7RqobtB8lFYw6QPYG+OIxXVU61O5ZKM4OYT4GBG6CCgoJVGny5rinB
jYRlr9WPVkKX4HUC9e/6Ex/DUrha196MSpK9Jz7surEIpYdLDEu80EGeuk5cv52H5cIV3edoEYda
I2xW6p6FnG6GliYBGNNo+8V5TR5c70mEWMLR71hyk5zeBWmyg27c/GojeeFApN0S29ulviqGyXhB
no8DvSirO30ji7dSNJWSg2onRtRzQr3wk0H7kB5/Rjd+ibrxWx1CEM/+H4OD1IGgn2OdmYASDxoM
onCZ+W27rjBKwkZaAkLIZnEcw8SkHK4h9ZswQ4J1n9rdOCBqOYH0JT1FGu8A5ALh8KH6zom210Db
XnYM1p+HbJ4zJSS/GtiJCnJ0ATebaA+Qtl+JhYJeehcA2cmGyeqZAg00dKtbflw2CBDgJsiPMgmT
sUoT/5i3Z+UiOknjHeAy1wJ6rRNvObhD4U9h0qaJnpRq0zfRspxJQEYxQdw1S536zCc83JYMrK78
y8EWgD8Kf4fmEwTwcCRbmhjb3Lp3183GUy8O9Exszehfg75nmg8VqnAfu1mpMDZrwk0OxJwvGJsx
gi9g2FPUYReg9Th0O4yqVU1wmKqEKU3gt95wXrx+Re2oi+7wX/35qjoHCVBa/vtKxLFNRkpc21b5
Ab+QPBGMnyQGzIkScpT9Exfst3BHQFVjbhxs4pVGPOzomBq8KFjIPSQPJklyV+sDpjF/c6NFy8S0
mROXxcEp92aBtFTZGRYB09ghoA3WWNz/tabLIQvaHUIs2HrB6wiOpeOl6ocEK/a/T/Y6gR/WrVZ5
+8pnukhQhntgmAgaoNZnVwd6eQXF6S1iclauTUkM42yONzwQA6galOLRx1Hrlncz8zT13T4lhvtK
WlbuNgc5RIVpi/qJl9HSHHe8nAOC96k1iXZs2b1DRw4RBpZl4NmNasQpwZHlUYVJGeH+MdyPhpak
nnM/Ec5LnPja58XDl19eM960ejsUE3TSx00iMpnHTAuCfzZ0nr8qlYGkgz7ykGgDOYIzHVWDMsC1
ogxkBsWKLjFkCp9gCWUam0lllIdCocfYprxZWWS2KU314M47VSQrSOTHDSHdm+BGtQM82t1xhKI8
/tKwto5D01A8R1FGc28BxJizJLPpWdQnGDGmg+aBxlVL4JH+xAi7R2CsWXjrgQAuRTd4DGnAMRU+
pWi1xm6fmU6fIsCoQJcs5v7Ko/LEgGkOIQb2MA3R5JFq7k6OuIdo8mTx6nuZdAYZP5cwTVGs/WmB
PX1KSLKJovET4bfja07Xs+xzK0U7KJuz460cKdJqFhw9/ks6xT8bv6lcnOcpGJK1BbPH6KIuLL7g
hyTQ1jqYa1e5KVAwIFSOaBldv5+cOfXbBaVIusPG+hTANkM3IhZ92aNf6TM2BvNSkcHnA+Ak0AOm
2eIjS4WINrkLv/WaHzl1T4cRoOIKxIcKv0M3GVcTRUmtGmgn+FoSG7Fp2GwTDplS61kdGC1S4tfW
mTYKdvTemT23RfVW53QYmOjSBe5UImAfWFkZFKaTukIW1R4S44/MZ2FYh/NErt38aj87PB9NS8cU
OSD0cUO7bKTljtsHZb2Ww7fqq9lUnNHBGxY61VzzBoKdFzQze4JOIhoCcwf10dmsRQt4dK/qBWiy
9j3eO4Q/hGF4f0iSAXNH3PmmldZNq1bxl6plEo7M2aDS41ewiT02pKa37SHBG0E5T9VBFmSyFyCr
r1hsU5OwqLZS8DWKF4AjaZP+tlSpm5LsjeGGPCjYo7eBf7/3Qc8+BZF2ioUKF+oeKEOghss7sIcl
b+lM0gWZfwz16RIqZJ44f4GjKI0YgLWR/tEJ2eR+3Sa5DOWNj4051Y0KQfp0IF38zkPoDqlIyiKn
MOqMGLDw3VNFqi2DgMmomIsVtiOo4FHQjg5IB5KLRTJCQCoKiWdK7q9TRp4/n6BSTkvFll4EeL+2
6A7EYZVzH55XJTNlEqEPdvfHfs2QhZp+DjxdnWl8dHFlaNs5mRnRJ5Xle5HINsyT0dG2Tvd1h7T3
rYrzggNQD5gyTRFQJ/Px/M+dKYm8zK7UTII1Mnqw8AxQfzcOMjBb/4Jz3Eag2oqnlXyvS/WlLsJW
8ZH4MeStel8Kv40yQQbv9NCeT371C5vTErOfUSx0f29ILAeQta5SFZthF/QnKFznSFFaImgegDUY
iQTErt6YrEP1IYzsX7gEXeZrgbAa9odwOP2simQPi3g7jtOI0HHtqAiv5TMGvLPfEtENeAY0p149
4FzmylpdPpFCFYwv9RwAyo8DCS+kB12cLwA6/sGqvJE2pbVmDmDXP3rcX0y/A9rucwMEDXNWiQWW
rQdrSH0Rez3R+BS+VcrTSWTqwgRHRvXllYfRXmTcwiux3dvv0zuQdBUptEGYzdH41auownc2KfHT
5R0n9VS3YgjA1Hm5FEBFZz8c0xMdHQaDTVNAs2oCy8B1qeQRyEqiokYScqpYUOIVv8D8QSXIMXxP
Mpr999oT00RE3dkNHS8knt7lhGBjtylnRSJOW9Fz7ZYFt07Ahqkj30bhF/pbo/z/8yippbOkqLlA
VQhxaCoVGjrsfyhfO9dniRN9pM+zWowOYTzjn7m/SWtmb8TnhneuwJTHyNc1H+1B1x60zoDe9fFU
43OQOK2zKrOg8L5K1jdDRBVuc5AbTVE4CGb7ya1IEhkRNk6MSh/BhQQDP1oSODCcIV+W0hGF+kFd
rVzGZDNOjorWHfRyQcWOEISkAhIZ6gsMRc2TdawoYQSDd8sdu+8llRwwgNrxTFal79WcTM1XTOG1
YDtsZPPvrmTQ9yEdE1xwENyTvlFUMnIpOglXnjgFYuQCBeHTqWZy31HuVMPe0G+qP9tqG4I8khrM
YWFe7N79+980ydrdTC5AZgenjPAL5dw2UH38/yyfVpc2zuSKkjqkzblCgCxQ4tlleJ5FLywrqyAw
hca+DMRlzhhjy1SS/bKmFgKZFxapcMqOK+gYv5dWd3+BvYu7hXg+EDqQyzyiBBjfA7/wUIYS3SAt
DXjl4RS8mSP8olSxIFiM81akdUzNDZ2WLcotJsYqcyzXCXEKkSJlVCuAXCMGoPjyQYaflHk838/P
ufsEkH32hYmoOYxISED5YXo3Eop6JDJHTtzIfJ1Z91W0UTtCi22+nNckREHmx97V/QAGF8hEgAO3
VZ0/g0tc9KQV8NgVKCzMpnNpAXTe2+6hg/yWd7uofWMjZvIDWrsQhl5FKxZsBuVsK6JI/AFVSM8n
2WYKCZDtXY+siSg66+BOEf/qmVvACDHNIQCQNl6JDNi08eu8DEUrSHLf0p2E8jiEDNIZ8RHz05Wz
nFIQvH59wfmLNo3LrLOOHq0RzacXh0sjbuA0lcDi8Puh6yIwsei1iX71kY5wMUr+XOCZEwvE1y5B
rXRAlL51AR0WWLH1G9yb8wFsny1X2VKGN2IQis9KBddRQtJDRjVnLNpdqozH1fUkzuVY3aFF2H/P
JJn49HYQXk2Rea2oMK+LDRGPPzMshzESO4aNAsqo0CS/pYjFM1nikhv58rRa6pnKw1IJSn3Yt5V8
pJIwn4oSPf1L7DtY00iwAW2d0xo/G85yMazFpaYvvxdAmaMbdC5NHZ1NguyDX3wKUOI9drsBZ7DF
ehEALZkttY1IFV+8p0wqO3mF57celYIgsXS5q9NTS1DurVQ3iQACHYTWns/WPDfE4sZTBIqk8nJf
XRmLhfq2JU9JlbMngQYz2fVJAQVVA6R9aCjbBXB/5Rg5mGUc/EYpj40XRVlQT+lgd3ja8FdhZpd3
Miu5QHf0gulFp+/ymZGB+2763/lGA07ltJPHc3nw6ZaypgSjcYMGq+sJeHnfbeHZCTeU1Mr4bvgm
Hmn/Gk2tIM5tA0fC7ilzUgDcxiSiDaokdTg2AxcpE42jXaGDRlP96L2cxoTRWr6j1IFZPTkvcZ10
vgIpLAmEMQcK0jcGviUrQRoHfLtX7Oirl7xV5Mclkj00DvtHywrQZyIlJruCEebHGlkBArt3dQNi
LDb/0i+X02+MF+73A88ly6SLRkOuPvJIqchi4ReDsvqTcIwqrCRWWfPk0d3GZe5Si2tR7/BlSWTZ
PrhG/sdRYmn8DgcQ7qUI7EFtEcj7NbfsGWBLTQdd0i+J/NaVqpS39rtEzXj2PG/D0X005E87SqnK
34Yjl83gmPicxLUZL0SF96Fm5kTsPPoeuw44eVJW83UblemZfGNO8hya1yI9oYpQ5ZaDJS3DvG5N
Cgk0JF4CgvATisHAjnTiNqdq10Su6bxTDOqLu8olXruTMv7lbzUUiQq4zKyTeHEsEE+a75dLA7/S
JSGdee6Nu4HN0yICW0jR3KECeOoEAB+D2/W2Xw+TIWk9BUFFWkJX2AVRNyeK5kgnAt8MfLN6OcO7
xHf7ZtaBMPbzmUsEpcClO3K2cqG7typdOb/OxKHe0A71gV3VZMjft7383aGXx4EWLTUf4Xb3Ug7g
aG3AhDKqMXdgz1Ldd3VONAYfhJ0OrOXjWxno9xEjtdZw/kzgvgwCfGTto5GTcp11Vz3xx4LFzGgf
Pn1anpvuwQqSVyXX5mQmWi5lsK9YE87Qriwlkpkc9lL6dxT7GTgqBEfNdZcKhk2MaMJuOEgggyyP
v2cQbqxKQ0v/xuhGmKCVHp3v4gvrzilh0Ts0SADVcljJx1RnT4FvdXClZ82WzTY6yXlBP+gaeC1o
ZMENkxGx1k5yaE+spj5QJvLQc0fuIbR1VCdkOHJDplh51tX8ymW/+6SbKIWGQ31JtClmDon4HyL/
fvpjoeOHKxqN9a/ebWHoi3hdXI302zKaUANLtSxs84799rnFmU+1mVFW2qHSKsOSBhdE56/paDeU
gCvHt2IsgbGeRrdHN88Oh83rgqOXpiTz2iZUhcfaZggpgFvIThiucCZ6GBDs3vkz/qLJ0RVBF508
e89EEperhsDTFb8rBAqHZbcusnd8srxZ860SM+HmDx+dNvW5O/mLuf3WmU4pfhpHDZYEGtWjXALp
GguKBuHs79790BLjUvqn3r+lJRdJbTSVQK1AQduOTXWKn2I2v7JF/k/Ir7TcIoSfgmINdwJxmsRl
Vf1YYGPitDHq+ZovChA60EI0yUQniumtwqS13gApDzgNdxm1vvjKyfldi8AiV7oPx8FqVdDObdR7
apTGWUrsjTVE7INwx+JHUFk6XkGdRt3VlPsxyYpXSPzB97bzhn3erwmtunAKm6XYbyHorF22sRw/
HRNgxmho02cOLI4kDrAwMI+lHLr4oh2qwXlnG7FeQv36J1CQBQ6bDZozdFqmj63z9yD3gJCKrA4P
A4uVxMO9IEEao+hy/rxPa0frRFbRIBG9bfySNQ69QH6PfdjtuzdQpRBpnPjC7MCy5al12nHjb0x5
nbBOkpZD/p5t64E+KaQenu8QedV2Uib3Kc7LCpZsfV5S8yu7/NgVPiW/GsflAe8pHw6GuJqnV8yv
qLLYEb+6SZmUXdINSO+gNi2PEK81iweVo6+rlyORS56lbevrb6rpILSkSWXSil6y7jppG/dPsjkb
/dNYsK4tzTeOpUM/8FSqEewbOYBLRmnxUu175L0UuWTQvyc+e+MATqay0X9+sgbLxJSliHUcoMyz
1aDhIfbDN1Et5+n27TOi9TIJHgFgocSBVslFhPtdre/EwnuJfSxuvUqEQ3d69qKQyHlgcanI6mvw
WEhapLU3FVwjmFeaY9Wm9MC+REdvd5K8U+A7neq+H2+wz/PQ60uAVrewBXl32puptLL9Z7PI94HL
1wMrzzCZEa9/JM83iSDBWYErsHLTLVsmnia7GAZxRwqWdwtygcEWkC1304IO+NwoV4yNc6nQImPw
zxq+Awvfs6ZTYGFAJOndXUEfdGPCbcYS2vLKqNMn52HY7IeUn+HWGA96hNPjqfiolVNp2/8+r6Sh
hHFEtGO46OtTOvKi746H/0WEsO6Srzx6OlGxJL/eFZvpS8CxTp/1dpJrZHcbWEG8Czvk50HDPOzD
9ssAXMJTe4EhKnX6w5vZv7A3AVg8bqlfEoIO5QKNbizyloKXF7eGaU+UfLdrEoWnActnXz9+uSE4
+MlMrGs7OzA5o6BCvxGCumuuWk4f054cfpIhnSIQpiD8m4aAnwaZTer1HZoHT5YlcOMNXsNVsx1g
wpIZHOO5jRIAdzMUBVItdDEJxOVdrtMXAmI7xiVd3kmsuF6ltXIiRsK6igVQ/d+aa+vKD3nyoq0O
11ecggnvNf3+AbXdTfnGfgtFHZrlkyDQYlrYlCZHluc7cMCBSPn9SkSvb51IVfWZtwU7EQ7T2FpL
Pa8zEY3KeeMvkjClMgmrNlJYVn4Qsx/dEtr9jfgo9e/ssW0ZWVxYrNgV8XQZOxTzm+kYgI2RI9P3
C5mW6bOG6UsYf/ta5573yq1EAFePmn8rYol29JgW6bWIb5Ofyp3Rm3fBXqN0xMiRHzM1as4rpEH3
Ha9VaqVnMCBsBQHCb2KDj9bYc4cv97u6MzPWq9ZsGOEU1xf+2EqHLxOyNJn8Lg260CDW8pG/TNap
YHN+UO5s1X2A85AraL17Nph3Iau3xq6xGJsm+KmBUicLoeJyK1KNxj5PpLkcOZaB18ulYfsUwEV1
xV9F4CEvkS8xKReu5D36JU2wRP4zeswcxBZF4r5vnhf7JksKYZjA8PZaabEZHv6F6id7wbLiS8Ub
Ng17gTU2qJ1Mm1tHlw1rKtHj2i3sZJhXd2oO+n0kV7KHdyohWXgWW9DDdFXEVyQxwq0JLsokST7s
LVx8TUrNkp3APouxXD2BskAIajn1DU4d6UNhXpdOe55aLqnMH6cxyC7FicoJyTDNXrYSLwlEkgQP
IK5b4FYDob+5abEqsJg9gcQ2+7Bu4zP3Z1ZwzYHEZ8XTJOtHpI85VbSpf/ZXoOrPhHU89WXrkl/f
tmkQMexKZo24pWVQ2lmOaqQWYECFrP2vUp8J3fPGuSk9+aeUkQrQczCdMRqcFLmlpX6VtI5w/j5q
CvnmwD2+iKxGdNdSHVpuPL+WFkIuvNZfHSAgRmNmKSdHTuVyivGYNQGbgF1OD8CRntZRNTEHHP1p
pTAoJhNRAd1s9QiMzS5dPzXaabmJgQscB40HQM1lIydNGLdTuBRNv1rIjm5f9iHRh3oSYXdbKt5g
KkDhN3VQlj0nk1GVN53OPfUueZyimi0UNH2jwTbVxUDqUO7AeY81jiDEjOrx/Djb+WB7b1bg/dah
U5ctSQgXs5gRtwKVByMGZDifmEGEojeKXxLfAuMwjrq5taa19hO7R3ro7aGnSVdpme7ITIEjOU4w
d+y/TWqWnaktPd1xDPjqW5bH7INpSwMi/QPWRUz4DIXXwQ0kUmVcFKlRUffR6YTYEpa1WMzNHSSN
n+iPSnZgR+TWKYV0IWCADT6LTbntJgecRiTZSe7nVX42xKJu9dYpmGwjldoY4aQVQK880+CukvUG
XKjfQ1dvxVBGa0Ewif4x7ow+Kn2vVsoHn9MvN2mJClU72faj+zfYJNJfie4GyIRhl3Yl2VJ3fenb
Gx0ovXhBZA0jpNjSBUn2iUo9XvcHJ9T1dP0YNa+TWqgtkDc2m/pt2k73CnZQileEC0ut4W1NukLu
Z6knrgUIuP9Q0CZQyzbnY/whgtQ8GgwJ60TUpmDv0vSfGX63ZxpgSkxb1yJwI2BbYTLF+6ziQ8xE
ChYIlWFO3JG5ptqacRLu9dbvwf9O5tn7kZ0CXe1gTs04W6JtU9cglx7PotaQNd/csrTQMdzcjq2y
k9fRFmbrKcOjGlEoPAcPc1sgxZ5fNi6XXTwrz/5DV59njCbQ3QDYqyf2o29pLI3WWSST4L/0nzDz
UXZhKDFK0aK05YFLcdPRA2I1lp6vLUnE8MuwBANJw9jpt400UWr6TnW4s/L5ucPHAC+f5VhxvPZ7
0O0IwCdcTWvAhfusMUL3vZxE0CJnCvr6ejb/TpXZRNPdDP5vjeWAgTAGRYNFjZofllOBFkwNx3De
NandsJpV6tjw5ZHj5RLrMdFdhRn9w7usY7pTCMLPRW0aztkPuDpdI6s2Ny5sEEbqi5/n2+zaFftl
ZDFEu02x+ziA0XDoeLrxmZ7wt0h4pQ6c57SDtsvH4vxh0KgnLx7tCmSHJ45vmm28RIsaAjsqS/yb
zLQPkMmvBRxMA3zVZQShumqj41djE7nCmQ6f/klNHcPLngMN1rBYlXvAn/hyhkfAD2PSu94LxIJ4
2YQ61Kh7C/bg/6NB69QaOn3WMeUTY4B8NvV+7ab6KFIbcGyvDbyaD03+jv+RUIyZCjloc8Fi/qed
h0NLj0ytzfVYekrLjOVa/j9W1KiU3VI0bZAoN3PHWrYuw08gUYI/2IQp9CDnYOMwKemo0LfTRcOf
5b0CdBQGP/pGyZpai5yVsBY+qLIETsKvGotiR/GA9JUPBoYQrE/Za9RSk51WAvW0aWpDuRLHzkQ/
114zpZOwCAwtlRi3IeYC06I5lBQkGysWXG2XZ/67VRmZRsyDt6YH/YFoQa+mfDi7wSbtlsYb5K++
o6Oos3T6kP8wIPwlkGhfqhlWse9xT05oA8LBbFg+fDgPqFDpmuYppZDH7MZfiulyQ4RW9KsZYlp5
ge/8NgNeeN1QiFOQshXnYjTb1vVMf7ab7qdeoJBpzmmgi2J5rApIPbIany9sQnApuzAlLe5g2TrT
fF3H3iIvFRvRLykWr23/5HeDMc8pqHC/epSsy61TSK2myhjwO/9rcpu1ukAQDrWqSLviZM68CCLM
buC/HpVchbHyN6GNm0eUnHO7M89/ePK5RwyqP0NlRySxiRuxRK3s7jf4Eehn/LE0UP/awQoIq/lG
BS+m8EjDBlpArZRbrgHu0xg1NcfbjZDuNxbDlSojvokWGzdTQFb17oTPMl+p/157p0Jwa2jeusRi
DCdDDhsda2ApY6BukpIjE7ezbNlGQjv5rQTxV8sSqDdwQV+IrpsSVHYtQdXeUQyF3tEOuA+sCTE+
S36ZN2PBaPZ3ej3hbTzQGduX4RToadCkAM5EG6SSPK6KPX6tv0+OIkSDgClbAboVLiXPBK6E+Dg3
e7nmFOMhzmT7UvRbe9XhiVYcVOpgsUuSigmJFeTuyhRyh8JABTu0/RYiQl/PuPigapBAKR44ZTtv
+/VI8KRGCAoLx4f6SOSMt7kSOPD4qy0uk6Zgl7l8FEPamHjt4gq9Q/1JMZbPc2mYjueLC8a+bFi7
FXUcfEEYDut4ida1tXoxA436cgLdCQVwDWyftF5jF06WdLGIQmvSWZCyoKU+dKSXg/Snimo0I5xE
aHg5YZDyIzVg0IlC8UXE53S5a7f1Z4P/lwQcKBn5vraWI+aSFAADTalcZvcfY9UjaFcNjZJV4vuI
QCJW2emHtTtATGsf5sSbdP1GQkpY8TC2Brg6BXcETKOKzklXtvPN+R7zHKm+QQnJIpm385QfCzNS
cVhj87XASiwAleTieyekCT166pdn0n7M7rYMnuoVpolumg/F0ZjvCaKFSbyHC4+S+Yb5nczojF++
xm9nmDq5HDFkVaqpWwqDGXYhkPKveEKZdV1Y0kxNzfDG9LWQB3purz2HBLxVuD2+LSdcowHi73oW
megb7cJubP/YQnvF8nx/kshvL3glEStReVg4+uvSL0AE69UHs+H03Bq/wHt3d5Be6gc2y/oPLcFw
nc0jvOqrQQOoaagCP/ncdpoqmBLh+4GE3lNzyh5QADJYlHrCjpez5B+E6I9toedFq1ix3CmICJwL
6XE/HHsqjS1LdUivO99WRzbnJ4yjY6VF4fhdFI8Rlk5czNXG87HB45ltcAFeN1RbqRumRWgr4bGM
ZFf01HbIrGijm+Zncd+BgxIQjZumZHhIYHjTHWqe3ySpANN/v7Os6S3vp8gFmESZtEiylD/2QyMI
R2Mivz85Vjpw6RwNuOnmzeaIhvu5tTdhd2/mohXPPpzp8OR9TCCO4fsTXlUKmnOhVS1KnXrX5B6t
OqD4rCT4YoEMWXt4H0i7gsFq7mX2L0faY772HcfthAu2Ug4ywLSBDdyCUN38gXEs3bnIm99B4pxD
JftcTOZc+YKSOKNC0CioZbXExLfaDaYKF+dKJFbfl0p5v0ikYtPFKvURpMu0qnY/rA3B03r6PIeD
qey2QI88d0lgcATyLypg/TQxjagbsGP3XQIK1nXAipuqmctLC+erQ0qpV+VHStgLAYJUQaQF7cfe
JjBkqZ/gSmaOxLue0mb3V07kR+X2NAtwmINFKTx3jcKEjVzbmRu92Q28yxrMfufpj8dwtA6kopNq
56PL//+kZxo0BHSOiFzisrtLuvtjEwpL8xzE1ztfyJ0bLHshyZAufSAGtvIBlIeXHrXUiemmLjQT
GCDJbSinJVkWONi6GZRhwvMpxg7mLVoZo+va5Bf1RIs9RlR9qgjH07tCJzNvvM2Z6maOyVl+1exQ
bi9oDeOUUSi+8sbAENznxt/BY6u8Tkir4zU0cbTd4ZZqK916TUgYN7e6EM9JrD7yLzht8jdRce9u
D0I7NYn9wTFvRiZY8VrtuND6eBNNy9RCdKaOLYQpn+FmTw+aX96KsLQWdSs3EoxPFzFqEX/63Frm
5a3v2EuiXYI9WEknt1ycCdWZ/OhoEs+d07rHy7HqqSR7SNs5w1ePPMdsUHzaEUkzmMmm3YxKLWr/
5hkcxBaKoVRFzXNHKtuTyh0BhD2kzPDGcgSPs95O+iba8j0ID4IEACHphHNQls3cUN/BpOdWtZdP
tbZwWdKRDdEZ8RNkIgPgrFbMj1nnhR31CuMsCR8SG48wTTT6g/oMwfpfK23KwBe75I1T5yUbKjXn
l4A3sfpZX4WPG0rPEwfLMWZrSn7p9UGdqW9mabJ3F1lKu8tkblH2x+TZxO6qSNPRdGmTRtdM9rN7
dHliSSyLGCm0x3guILhCS0StD75bymNnoOsjb+2vvoCaowjbydpdUsjxNK/e4eGMWzYCLX16FWph
1M4zMKU9bF0Bja9MerbRvPPoclhBeZMA/AL3vta8erQfb+2j6ypVj7Sp5Ir9oNJvwflQ6myaR0M6
mdL3JZHtVAOgSQ0fIIEw0Chk3doT7ukAjf1Zx/wJ4Kp2UymSZ1npZXp407yn+8js1lrb2lKvlIiL
Q5nODxqR6MDeTnyyTiX7MLV4Dehw8lIabzWHukCk7TJ9OsAXd6nma0J1SIZfj1OPKJ3bBqgv/1xI
lw1Xtk3I1FAMkCwddxa5J+4+svLsKetsDcqn7hcBvuU490mygYO+U6CEn/zMK71wL5kehiubcPre
c0N52ZSpmaFxoeK9Jfh4KZmRfuvGJNBn88KiAO9pbYYWpQqX/jAA621hr9UB9zcpzivuY/rdvCFZ
uxhC3UO1V2GAI1BE/CnCveegLWEiV5lp3uaoqoRy+q6V4QvvXgahqqaFfggUQyHg3BJ6wk2MdPJH
uS+ioIqPaP1DCxi9GrdF1ptrE+9a8L5br4uUJxvWhu0pfH2gHuPPgYEzdJKaWv0C33GRBL41lzgb
RECyBMcaLR8KXEdBcSz6p2PSFi5IJiewodBpVE+Uy/g3TJGVXBFlkvwEleUpuk1uh3eWvwv9oC4s
5TS9Wubul/Wt4oJGIYjpnb9syu5Gma5YQicl9VLAkEx3pOTCYBr/t02sviGAM604sbSsOOZ4bdKv
5nJpq2UDt56KK5QiEZYRChSBei0GWbhGyYLTsB/PK66zajK5mjhChMwAUkujmNq7JMQdbpmyhNTl
pVA/2hmRupeXbOeW8IebVcLu4AmB9GeZljYOnxBnEMgYb0Jp5vqjWzoUyvU8psyeVD0kaXQfWLjN
GQM2jgG3eUhN8gnmS58naxWSTvz9q6eSRzwuXf12sH6uS5/7wsgLr+RvTP6+IPEIoluZy36uzHRC
IYrDfzq+vpVfHboNHlYl6ksaECNvP9WOdvL5VGlsqYL1d644GMwyOPGM7DjFdP4WPZfeRAPo7/8m
rW0Xkd7s439Fu6sJdWiMrFuS1zLAMXC3J5DW3JrN+yNflE+sFuBtZ6wb11xeo0H/0hYRwN+HpwkM
4CMzoOz6DX+jgBQ7XZ3OND51j7HQMHN07a6lbYa+c1si21LjJJrJZn61JI6AMlgXW+YPNHZVfyio
3YWpVFDdI41l7Tx7TrD3rGCtiG6C2/dMqFoL71EsXhAgNAYqYg4o5BmIu0U6J3I77pFDIdizRHA+
cU1Jp19Lnc+Esgj/DM/y93IWiXULMiyIPXINGbnwxR/k+8mY18e1fFqKYTQIrnyT2SFStfMTzQOE
2lIeYmL7k5c4d+bHd6LL1K8h74C8wvTYqZxlrEbjZR/g+PvKPikXMRAdLBkI0ztPH0H5aw7jqGTd
2aX5XunxROw8As2a+8setYQ6hvQ3lmFoBvNCpXMPdZtri0HyUNJu0K4IvRWbdd4/20p70PrR4BBX
/zU6kx0h2+MZRZPmEREVBkVo8pwj5xilXGx3D1ssYia1KFr152dwW99Qgq5eukhimW7AMmSw6j8S
+DsAJ8s5+8Hd+vB0UACi89TzRQSnTvUGsQpchOoMAAEUIySi2Aaxmhu7QHDdiOQowcb3hKZ+jR5G
78WB5zyv4/UCHmcGV17sUqNDmB0pWDc3A4Jf6snT8WsPo7MNEFgZEwu6u5iOeaqPUnO9CTn8uc6C
1rkyRmMYI4JuiLGuT10k/Srnk28bffe/h2Mtc4qSig4jAmnu+3pYDSPnWGFkT2pqXOKZMY9JsG8/
/nFKQyh/Y5xa4mrm2DmC2p7X8ltd0Oy8M1nTOKXWq+nCanEMGOaH7k4m2hQNVqTExXclsiUvhvJt
anGonogL9onOrNSWZdqsUwUdi1i9kdAXLPydqij1JHMxhsSGnBppQpp6cyrdD8m7Ne5ov9aZ1FQn
iVi77Nshf+HDJ8v22RIaJq21+8UGMEqdwDVfJ/HPmSfq6c7H6F8McrrWnX/sLuCXpyoT5mgPYair
AmvbqafOmjvMmqJKklF6PFo0Kzp7xPO5RFm1OW3AMYcyhvPey/vrzQD+/2P8VGF1j2UGVWwoA8JG
f96Yn+pJThQPx8XKumIZtpIjQmOUNoa0THDxMqfNiUFZ36ZauJq3GyVLm4CRy0nkobZxEgTwGLMZ
Stqn1YuKvy0ROhKDdnW2EIQbr1RG5n7o3Vl/8RRZajaJwDKjT4Awkbd9Zm6LIBaq2/li1E+CzwDd
UtFp5LrVvRYLXBj2MofmZ2lCPwmm1YNvBu/XERI453/hOArnJA0iM0BiHJQc6MkzpEWox+wwAC+o
94R98ZrfKqLFQ9Eyb8HrKy+9qiEd9LIl+AWJsOwi7PpnjNnZQYbSNnNHAsfUG00AgCFSPZVAZ3Cf
sLQibnIPykioQ0UD7H22zQ7PR56yO5Y9RPULAGDCie4n5pUMb2jn2pUJmCnbs73orFj2g+r59vAW
lb5wI5p6Rxa+zbeggLtah6niFnv2g7wTM4++cCfE/+hrqtA9+OV7AdT/pJXX9XQQ+BoDD1zPMaG2
UzD3QcisTH35h41Ux3FYT5KvBlZi5faO0a63fPQZvpEc/L4IAX17NPZCj4S2apBULAsugBJp/zce
XoCdHPO208x4Rvxl3YcyW5ugncHXbjRpLJ1emD3Ytovt+tRABBgzGzvCmjZWofrpJlWRXSDdhndJ
GfjaUFQEsetbUxCRM4E7SduqntwRBsDlFxCaOc/uhC93ZKiloDG5KrCKstf2YAbWzTT1zjmhw7F2
BgNzSt7VDO26Wb1JcnTUKx+bNaLBOrpkn9jZiev+YP/3oMUfwaS4Z6zmysP9EPSk5/H0yrRPcYrp
3J9aBIGBxWNpZCjcht3fsdvkJVr4TY2jpzgsjAvY9wsBEiHeJGd+TZ1Y7qeQVmLXe89LqMxPqFDB
5ZyxDf9sdernNnCZnDm3xZGjmLv7eg4y2Pf7Z7lXVadKIIloFm/F6ACgYe13JJz6zumvrBtjkXVX
G5D7q3l36kJITJ5BvHNjVpsARQEHdeCEuMPrD0r59Js+UXOOtPfMdjVDWoDPF+whiFP+XyOweDdx
4B/MV414+dg3KGRdCRayKopoRx8FjEt49Lvf0kI+m38B0krNjTeNhB7zxHNpwL5U7ooMjEpP9auZ
5P6cLW7o3JvRvIaBRl7uojRFCqSfBzNPoYfI1jlEU6u6QbfQrky1oKcaBOEU0Pj0n3FQLgCFS9Vx
lDXBfs7B9TWi0wEte0ENzyhWfxACLEQWHDOC3NYBrRo6ovmIVUFMApt3CyskSQWSJAGLGjFVh87d
PdSwxDnMMv0pVRFWw/GUR0FR0plpVPeQQUd+HXiTlZcCS5zjAWvd5b8Xj0kSLrvlSRJlmnOpLjxN
W7Whw/faobvB3X1f6M7iyduar7fe2g3kR5P3t78vZeqmNORXbZmS9FfOkdIDwYgPx9HimFYVu25T
FAenW2TNVemt39Yf3PA7nKx+Qwn84Bz8Evk6pfBnHSp1oDZ4tnbyeWYtJGf5lAAOFmg2jQN6RVSk
sMZPGNU6HMgGiqqbjlOd5h94TgRgNAm0ocvIQYojHqQrcSqf35wXoTL0aT+hqeW1P6VX5jZlhCpE
/lxxjI7hnD9W0lHRUL83VP7cxHQMXvxiJtgJIkZyzie4jGOrl9g0A//4k8bS7B5c/MWP59ke3Wt4
PutaMF7jFDvFir45tzXS1lJ+Wc5MD61r+/3odYJChYr0gJ5OTUI4sCoJWJ/+ACRDb1wBKDdo4Ro0
zYdrTRM3QO6ERoCSv6uJRVYmjbh409dXRiDOp4rimCiF9wsV9n/4oNQ0R5o7dA+HJs8OjTlNtS09
QEoy8Az3JEP3QViN6JvG0qXwVF0zv5NpmV7o2pm9W/NZnANedDKqGeMYrMNSB1d0o/QijPAeri/P
LZ2OrnDWlIH9HS1yMqDx1gLYDuiZMRrGR0XpgjShwX+Y4lvyH5hZnX3s4v5M/+AONoZEpsnDrpa6
oXG8qMBLfknCVgX1dUZC8PgzQbbh+BFUFe+RWk4UbfFw27ZXHH1ABiL0FxIMDlGFhmgHiPKKPyEy
NGeIOuKeG66J4dCsqpKBB0lk7kuRkV5hMsbGzuV0hEUOKmhTSoycTcfRillUnQtKQ89yJGCLoI6w
ECE9abJgUTiTlwNsSV4l9361dJl0XHb3ngpLTJi5cr2oylcExGp/C07yzGE/HZmmGHpbijQf0Pci
7MkMurr4IC+D+Ts3GfECY1e7CAoeSz0HP6bTrOEWBvaCVREIRVgM62J+ImsTShNzomcMZWMpeHOl
L8t1/f0OVdJ2A4OLoH7xC7xdKef4EgktbG80xt8XL1MQOkBX+Ln5PcKEx68fqcDj8XPnNhcXb+kk
pzE9XEMmi8KkG9zBIG8uzr8rijmV13gNjEc3Ck3vZwaxzRaC8A/aRisc2bzSalkZRQtOqW627Mga
cRjMQZE8T7iGDsqZE315nYGyHwoBLZSGB2qushdRH4Tw1fIMJ5pcV+EKgDWtOxjRANVAtXn3eiKw
TGna/7da1sqX8ymEcytELHHtairHPLyjooxZgARdMJ8BIoo7qeQE/vHOpCeiZEPjg9FzVYv0xKSB
q+Jh7U+nqYI6IsRVl/rA28sgID6UlvhxW963Twank2KZ9JXAj3XUWFX+nvNzbGQwkxVoKRioEdRn
BMMwqCpckaqBep802aepBgju4zSWesWAIfpFg+2IvKLCGyAMM0QdkvewcmeFED20i6NMs03lSIjN
tsQP7k/w2CmRrMoZHfwIwQPlIOnpvXOnSHI+unweWbwElKcMswwxU+EFFuY8MHY0m/gYlhC+K6mr
Zq+i0pf2sLpP/bahK+cNRIOw6YsGUz7SKF822Fp67AKHdUCay3KnGs8br9OyqBykxwS6G8ro9OIA
9TBmHkEPWnW0vVNFhSm6iPrXRP20hpqgzBObLJqqYmxmytOHxjma0NlL79VM5JCJMcQAE+y7v1F4
bWClM6aghJq0akp8OinzQ7ZT4nHMwanL+jVifukSKHEe3+dTGyRAI3fqiCPP02Xl8A1urUXuoHmN
X5jXCN1I3Z3Ks0bCXWlVZYgAS2QA9zu+2tdCMcUU4IKzAhNe6jv4S3gJg5swmqDOFJbQ5e4RGLG7
G03MaUNL2sG24CIaodCgITTmEs1K6x+FyCscd5j9fd90z4/rTgwJHypPjhK24alBJn8iBQa5sLCz
HUTyx54SJC0IX2Q8hGreqD0uxKjJ01s1jlulUMRYzUucL9Vqt7lsU9tEfShpBTmAOc/b1BCjnxPR
EdiZ9ARdFnQShvFOZ5miLnyNCKARJn0qmf1lK83EyY4or9O33to0oP8Yj69SzqpwaBPdy77ThQ38
/8wCUw15oTcy2t3YRVfEzSHztAHLFsVyp8m0eSxjvURjI1CgUuCHxMRhSWei5A4Al4ahsoQoB4SD
/WjNntcOAADFg78zwc7cwn9T75Vy6GM2KloAjvf8TXyUIMjHN1WLZQoF8/CJK+7xbng0xMcVA80c
miEeZloBuHmO2NcDT7VeXENighSNkqJ+FNbkUViFDwvlAQIovtJBxlizy73+V7/zMtlhQ+CGFPDn
Nx/w1aFlfxofNrR/+4lwHoe4Gi52w/O5FAzxBRaizkf7yjozjO3umSSbT9dVJfUqTv2sol6ezpeB
JfSam7YsE2skAxKid96Oc8IDJetW4a0f+7qcj2dy9vN4mGQZkZ6wCy8qoJuMEtB587gUY03n1D0S
J1J1eMHUKpDYqB9XYnHEuvASVEiCWHvnVOdMXAGUdbuvhIcl3tkcR7p9JsqyMjL/vTame6OguzlS
X8rxi1toSexLoR2scXiykGYXYFUvQxfxwBCjZbqSs/0PyOf5lggzWfM5KAJtBnqfHpfi2O8aVxF+
w2f/KdhNOThOdQ1BU7y9WtGOKK6RYCjoROfDoVUrLBs3qb8aPmbTCsw2W0vQMksh+vQICrscoex7
DSMvNX57Skn23roC4TPNi3AW8gWjAMOxLp+ksjqnl77i9LfQmNKRMgMK8Je1MEIBYAmtYI/iaJFz
b+fizsc/6rdtWrj3t8eio374pq+4uf1igvjrY3WOzkUpaS8UY3FkyUcNOuD9I5XGqxGgARZW33EP
sJKbT22v9f1BfA/VUzcoKbjfeqLYnWXe3YxBvh8IcFg19y4PfTaSz1hhWbvQy9Vv2KxibOQhJmqu
1wUNbgJpOHTIcs2Z2G1c1JmYB3mlijJWHY7YAsiAA6uE8voeE1VReaZMY8/AHZsL3XDWsqe/XYOR
TKQooBhCgU/rqVO95ix/MKSgFCSRGQxuerapGVsQU9EqlUw1Qb24Q/0mbqluHRMj6Y4N7cbPps0I
CACBCpRhs2gA/tGoWc01z3I3AOcdQqGfIE08O/CvLIgKjQCVHimjXEPJJNjObK5EatJEACRGfCNV
WeHW5Z4nPYzmz525qMsLKS+4nX5f1ID9ONpCeM59jKgNOfCun3HBPcjSyKG0SbCcbrprc5NCBzx2
2p1X6PshOktkyumftG+BGxPFC4KI9ciDS5rAG8S3LoutVHFqJcbdoxG8dpHoZ0BJwof2qx0gzV/T
ZA1yjCIc/KU3Qj2+dClId/MHPDXWxQrxJmtGVPnHKqI4Db9TU0jlzAZ+UjuN+kfVF7SS3q7m2MLE
rt1W8xb4zIt37DHOqhzrEHYPsRNKV9sUUuVBT7wacYTnQuC7GTA9r3RRN1ONP4b2NsHOx8RHrKl7
QsglSgKiKLsZvZKeaQK49XSYAC0Xc0L9fIl2sF0smG/BMjxPBy2FnauBeK1VtbBEo1yqSuk1DWlT
aBka4S/As9AImFwgg7B1jubUnS+Eiw6rDQA/vOGwJK6eGz2l91ijUG5uIvFoEhAIezNQwm1jbgfv
6kmL8sYtkws2+OcKFhbPIlPp+jA9zCc2MQmKDTlFYewJ4VSBefrJjiwZAWeyiK0thrFdfSZaUy1F
/MNSjcQzk6P8zczU5vAYqpfe6E3ECC/qQMabDBoGSuse2S0ciL1jxL3cvNpIFBEkgd8c3ptVs5Yo
oWzcChW4PUz2KCtQXq+qNn0ffzUltPASLTOCuAY5jEC/cZ9e8jxJJqVc0Y0hHnqD2/chS99XFUw2
yRIYOV7rwCetFRGUZc/BUweEELfnFaF0Fk1ngqhhuKysWiD4I1e8ZNj5Z8XVvz4ChPCzPAQC1+7y
rlE8wpR3b/+yTEo3Dn+9uXjP/OnNpwojFTPMB+BBHjMkq/4dMEQLviNgA0+jp8ybbGs8BZoh62pG
iT/+n+79Jm+/yYwSMIcDX65mJ+FtAag7B2W6pcuKkbWC+yCnXkH3/+BGU5s/QWpvdETdMYjVH08G
x3haoz0qTTUbLdqzii8OuZjGfL087POr2I7LWth3PwRR15KPTlwDNxIVfuS1zc7E7Utx8OvWHBgd
cV4yYYPJ6OxfUFMezxWt3p8a2wHtyCcBYyBgTltvsdmWdG0/Dxk42eIzyZxH1n6x2YLC7Bjcy2f0
3dGgaKwwWd1bfG5WbQESHzHTZaxjZaT2EN/K4iBd+4X7jgVASVM4IYhy1m3fqtPIAVoTrDtZ9Cj2
OlIFV7Ku51FOlN6/6Vbtkghkr8BaMHfM4/CYT77GTgbvJyeMkwwGIFrPFaXFn1bq1A8HyhrKXpU1
PR2YLs85ZoZi/8sZuf6IDx0ooV8K61El/fESqtfSpUoBEmXYsIlZidPnKj8rvoQr3XQwSv9cQkze
IliE0ZNLP5ctNIELtY16IoILID2UPCHT9nHNfvr3OUEB1Eu+V6+zfsHA5ul2APGISI9zu4jQwnYD
PNiKzkYHLnN6A1g5GGr87LukrqdkunZ1f24NRZMEoh/lwJoZXtzEZE7/VCHVaoOoj1RAnAlKDFcM
U3k5luGhJ8xUCrGxGaQHTuXzBXnk4TWuXrhcFoOeAzFl+Cq2tW9wDe/aHsKWK9DGQVs2c7iA/oou
TFbUqxPuMli/ftbtcgXkNpHHA2hgxC3ee5B1ilpRLP/oq3hdZHmFE+sx4wxCVMPVE2LtusDNYeYm
aQ1VvWR2JI10KRa8HELrQkvKgoEcFL4HA2TIq1hUCMtLHzVe5Ur5kWMqXGv+PWru1Rfq4HoEvvz5
hD9DKvwDg7IH0phGPb2eAy5VihaU22Pbl03wNxanYhrNhVARJVjEgZUw4Enqla3pi2U2/3ga+HE2
gCgtUP1uqG2J4dNnAFBG9weJ6HwM4ozk7TPQsZuXjd+MmBpl6btXhX5ymik6cM68A0WVWWQxSvhg
zdaLmH06Z347PsftgMr1HQtT7GuBYXI7vqVo5qhAjQolgk8aBuB5sGTln17FiUqRTGI8FYB7pe57
IVQ6iFFiXitqGirwccZYgxq7WGN+G+QqROz7P+lSOtwo+l9n0XFQgzXVG7MhWSgbjtgD7aDIDrCs
O5vEvNKHfwYLWk65Cut7mWIDhd7FYtuRTBvpzrjJBP5siAT15itbzKME/UwHEPDHNhHQ3ehd05Tx
hJX1f7DQ552oKi6qefLR+emOpWewLHzhjDcnSCDsL5iEA7CVlijmnd1+kkm+FR2fb/7f2kbhMPkg
m3aN26yRsnuBD1W744yoq3zk+u2Ug4YBJDn/vgAmlgdGNP/MdqhLn+rbJHg9sM3Ws+bj/aM8OK4t
Q3ZSMvQYIxEHPGwXs5AAnGfOLC0AGDF3B/9vyCGOtsx4oIIPb7+k6DoYcUCSrNc2U1EzxGMjSfXI
KVrxOMbekoEOEfhKFWQe8J8r+q7c5+JVtv3r4xabUDb4K1vt+9z3q6fv1jGiXvHnYKD3NcQx06Nj
aZhlMtLlS6OKKL2r4p9tRRGfSYJBwewMG5WW5uvFD7HCIGzkQYIXUwE29pdjFaAQAe8OCeQAMCpQ
H909ATSvmqei+vvMrcMBWXSAq9UK/aFF33RT13lOPfSdpHCHn/41u/vP1/qeuAMaF5tcz9VMgDLm
1l3ZPwIyLX4XXRjZaz9SAOpjHkUIJG5qithFtyyvNSNhhWLohiTMR4WLsMfA0YTkcMg4Bg6vZ8VY
diU63eX7GXIzrl0vjxU4A5R6gPOuvEb/KhcO7MPKnniylYGX6v8fVeS4sURHJVUYVjHtek7fMwhF
hRmXVtppIjyPPTLt/idq1SUUEyKWWbLcFb+SPV4tDbQFohVQh8C61O+z1DFvXvy1goVDc29RO6sl
1072XumOfYC2ACQVtdmsaGj1K878of/OcVZDaxi35mmQ3grwgczpyA8Y3V0kjYX2Cq9dZoeqBZF8
oBKcsnaieJJa1El/j/LJhdK/SAM7ypfzlO/cc/3BO+hagC171G11x/3jT0GFVT1wHsL2gcSChSWl
0rGWeOK4b/bvx7pHy9e2QcVrhE29Bqc2ttyoPV1JBYGZOxddx8vkIEymNgUWrZmUCXjYIuUZSPJ1
01ltK25HnB3dAM15D+7KSwHHIl1ut18RxUlWymQCn3ZPcy7dCaFiOcDHfKYP3si6hsOx7SHEAusc
+Zfgl983nUd9uDa1IgnaKT94q3f/xIWCmn/MqG31BaSStwJxfAjVK/WZffPuI0GMFkU+kwPHQ2wh
dhv5Utj1N3tw4rv4/HRbxS0D8y8BdIPhKI3fbg2DNSEwYFX3hiFLEacYlSMTTANLLUCMnrk9UNAm
u5Rd5ZfCVV0IRPEP6hicSOYGNWVZeYR+Krxzqq5b5Y9vXS7JiZL8nyz5sWQVBI3TqoM1bW5RD79l
TRZCyTjVmv0AJK59KOL9EgnQcKX2ExgkY4lvSsZ0oyz0An71ARtLvYNSH4A7BRDczgGwvHTitO2J
I89oQCQchOQXMz/TMEZezBdsdawTBimEpDh88F1d/lxw9G5IZQQ57kNeWixDHreycePKCwRxRuor
dq3sD27q89/lGWj73BFV/6Wdn5ga5cl8la55/JTGTamBy/bAS66PY46HZQYzATdcR4OwtcjPA+1n
bmETxHwyqZCaQcIoYtsCK9879oFNFnft1i2L7pg/p/FCetNdkDuwIg9D0e8b3cBFMstuw+VliQGY
kyK4JstQk6Q1ENIc98v7/TBzRe2zrj1YxemwcarJL/aQcykVZDLwhNqP9ftrdgLrX4tWXh6q1iWG
gVACYbcEQqMIQ/HvmIbfsB3zSaaZ+oq9+Nl8+COjH+maO9EL8q2I/Zdc/l3YWPE/CDeQZXLT7IJ3
gvSSiBxdJcYDCpfnNlzhqEhc26YjR3ug6ZddcYp4rD/bVuZIodjU1fHQZmrO7eOIxvrQZAfLFwdm
lfgmZCMEgrfjxijbTOAf25zVzQNjjuPRm9ce52xp5cEN5zrbXL11CTMa8pliYEXL1p+rxcgYWK4a
S+AoQO+OMR0O1hqauoDp68BZCnkOnC7ewmdGCdInAq6eTJoXnW7F540vMxRbxNMK0+s5EiYuYWlJ
0ElTh6Oq9rrQozD/ssQWB1Ia6vcFalQ1nPFIV4Gmspq5p+MWZO5ecZqn9ji8kdDVDryjHvWmuw8c
YAZhX5zxYkZE/K5wczYnELsGnlOV0z3RyJvHDPbeQVqNsEm0f92GTYsOgEozCqghQEyzceDOt7Bn
4qnS8dTtCDLvQXoe2e5BkWVc/39cRb71CtCSQMYDAZ1VRweZ+LgsNbZ+bL8NtVKgvS3Ixy35NESd
SchMigp3L8V42T3JIzW6SMofvLypzSakHlWmLNxvTXD5XvGI22a5yGRrLhHBmUR7zWj1fIL8Im8D
CwFMtsQ24VGwy623vCPp+32hFmOfLblWSO+T4HH5XTeHf4J5ELhT27q/r8+1o1UU1oFIhnnBx4Oh
XyQcbgt143yZlyya6mXiKk4VLSVYxpvk3rm/7egSYBiWzwGafkST2F/otxXVxh4eB+Q8hjvcRUG+
kkid3gJShgPs7Cb/+FbdX2w+uDz5JfDQ+M5F9OImyWHxWV9oWufnCLoXXgXlgrQvn69k+6hgDms0
mMNJd0JvCq7Y+OAd/JOuPh3LtU95AYfdo4r5Yq0o7tOx671J6457rRb1jXvNomMrDJ7k3p1BTiVR
48GDfBirrCcXyf9g3SnNYzszZGoN+O9R7YWVXDTnJyOzoVHMkHlcs9pCzyGSZWv9XT+zkK4JOwcq
GvnV4+aT1pgkybi0udz7xz4rs2WCUe66fvJ8Mxr+KfngRKthPnHjk4GTb0brTG+sxLv7pL+KPc73
z2pKemW6eG2BvLH3k5B4eH++K9RoqkUfRAlYQDUEtNbKGxrFOsieZVX+x2pvPqorIzQijyeLZApY
UlNeOYs7GMF2Psusfxp1nGrzK0q+iNHh3ksPyoQzsobB7/1nRb+TbbRsZ2Eyoph5OS4hd7lf+S/V
2A/ikRY9RPcJKj+Ar8Xcrw7oS2IJx4nxVRRjPvNlvValIC6jiO1FB0Hl4kHXl3P0dIjtS3cWdyY4
wiHMfBOAR6nJE3m7jnmBgAsXuMT5ZPvbOmrhe7NzSUuaaHVWi4oG94NPkynRozL2y1VFKlswNK2l
xTHe56Xq7HZ6eSF9mY6M5Cs1EQmcgudPmF73nh8M1fFur2DeHRJszct0VKM0u+4HJRMAr+jBusoT
K0kTr3JHuMccb8clAJezMUv4OkKVsniGNTuGuYIdHStQ8qR2EuFNkj9FxOvyqmhJ4ae80g72Jmkt
BFPEA9snRHhYLGdJI121keepO0C5O6ZBrp/+O/YAogum3W2yBJp0xNDuc9tQxKSAGf+U3Olkjm84
K8zH/pZFDyOGhUFKuvxZyDg/jtz6iwHYWE5+AtjKKpECpuJPnUvUpWjiSh6vC1mo6rPMTfqC4tre
PCcmkvAjkMxk4GMvLIBbkv546Yuctq8j1/4xolIdyjxkPRQX1Fg6uqvVmBsyNj953zDr3VWEHobi
FQL6jF8aedr4c0r6vG8BRLYT2Sr1sgk6Zzb1NnbsqUSG1r4HYw16VUUQC+gI77hTFPoIElrmByog
InssKxso6K6FbyCDdNyzjkTkczzgha4QrTYi3Bv2WVdmLRA3ZLGEBcgVVjLWzQPevIAu/cNrYNMC
cgkanXHfc3JzrzmpTo88G/YOBVjZjEysQnFRWrHan1iUPVn1yWagSfDl8jDPMnvdmr9i7jXal8EC
YsLBMZryM0bN6cDgV0srqDEhuQhDCt/po/40OGXGhHGAR9EWWEfrm1woJN65N8oRXl+sRksdE5BE
ZkblF8UqlttGkHPkPwTA935ZlyxK2Uiz5vB83PqcdIGQHZrbQCdlE9VAaoS8jXSBBW4/ynAtxQDu
nNVLx5bPZcb1+VqNp5yz9NXpjdk3BUkxTqrrDegbCasS8ImclapDSE0uKau9TsmIQghwZWLqGaY/
+lTkxvaccp6ZQ1ur1QMCj+URqH/6EpnehidM/7bgANN6szQSLPCAfRX2Xh7E0NagyeQ9bBWAIiQP
C9xEAvA66/CqHmVIDxnnrrZybQWIsO9CjwuO5iLPIIt9opm9+OF1FCMRRsMIAkax8trm6jGH3NTj
ne3b2V61XJI7Zy6EhlWhAMpFUMtrrzPUGxXWK47vKDaXfHR1awX9bFUO4orKAM8DYKm7WvDzAKV4
sI0TJ7B/dwXUxzJCHDI6By3DskKWwP/sb+yWd9vwFGiw26BfuYDml0pK49Eq66WETYX93RE5FvN4
bh0jpe86wIP0fUREaN2B7tTFiu6Vzuhb1Otih5Jo6vNeIQbx1EUmTiz/GNOxVA9pz0jKYGczxQgT
ORqJh1ziCHiBz3GVfmUOAP2eDJfvtaGjxekuGvF6AgimCyFmY5MxVIe7vvx31HQIszu+jKKdX8eQ
vGtwHdtdmUeypMdQ2BgRfdpbuWqceQ9IAG2MRZXZxok26aZKt04Ji36xZLBdpkDQ85cEo45CDt9Y
lbMjtrSr2G5JMo5uX4BKQl8Z0Sw1VEVetssUPbBG2KO0QdN2DsOOr12RMA4VPaTxfz+r2VfJ/Guh
UQ7huSCdYF7soxX+KPGoyZj9X3JJwfPnpolzT5XjFmIKp9uykcOImBfVmY0YQV+W7OCExkc/cJII
30Ym5Udisg/Mu+slzS4+FHqt3KYFQc/wML1GaCPLDsLmYthWiCb/jHVeRL8QnaOfsdYlY8k78mVh
80k6ePIOaRRCBzzwyYPFjVCPBQqFH1YTfoFiVreeNSt/gi8RAYXYxkECotqP7R/VCxY0KcEy7aVz
iZrsqJLHZEs2DICuikbK1OGLtd97Ppe4KODFXhtjhNA9l25nxg9ppFlv+OOpPBQJZOCoWQf5cR/o
9/lrznnhQap1NOowg1ssaaSJFND5P1OjQD8sefN4oyvSFo8drMNna/BtDWIG5hlQH0KgIy8ONOlc
enbMB+EIXFabi9HBWhd/GfAXetJZfIkI22eM4P8mTKkhi4pQdCB4HrR8yMO4xjDE6zmVK/hNrpse
vnaRkYl2Nsc98DBlpzUHoWOcvwiQ5WSs7fy5wcUeIGUeQD1Ys6Z5b6dsmYLHbxganBC6x4CLkZbk
G0Et1lbweTVF/XnK6WH84K5NDZqVi6JmZIQCBHq9tEog3iSChqh1YsLXv2rWoMuIjdqcYxONruW0
mqJ56ow717wk3OsBFRDCyyAIHBjwi930jXfXjQqKE9XwrDSAMzSAv8e9WiYh2UWwRuG+I/TOVV1+
ZRV7PCOYjCQT1aZIhHxN6KDqKnR/48rpyWtIvZWmXQDXQQrP5F6xcEWvziqFxJJfTpj88ZC3i4Fg
pyPnubGNsInkNY0MuQyLS/F6bFCRiruBe8S3ceyoHdyia+JTbdOWxHHNYL3nsffPpGsOXQoJJcyk
jSoaYSNrZy90FeK8RiBXaTgEudTOtRJfRM38ADYDrvnDinB+FKj/yhpcGb5+O5fdTdVdFFLpB721
Eikrpkm7F6Zaj2PHxPFiPh7lhSXAPao/9U02NnWOlVPHFVa86Ux/ocHlvIECDFPwq5LAanr7/Ti7
PjKSregnBo1aePHZu9cDQ5eCFuqNEC2SUO5k3SpNQVFzVXb/oyCXv3zGh2J8DApypBSD8l1qevVO
/iDJmObUlpc+Ub9UTHK8T0UlIqoF+zgCSRiZnLxAp8jgMDR84JW8hBtk1d78fO/QW2E+3ka3E6Vz
D+n7ayaUP+ckfhFnnkWEc6lv87CO72V8VJvrk0cn3ODPzhUOatezHMaP2qti9avyQg5KlGYs/gOq
q2CGGAJqlollbwa5bQBCo7pefgd4n+WTxHDaj1iICslkkrzKq+qbpWq0aBKex/3ng0bIZuUwy1Py
sg4fRDMSCncmc9tofNETkO7B87GgFDAFhiGMV5EIpbBK+KwjenjKFkBXSMwke0cMJPia2xGuVTUG
fGfY0+9UjEJ27Ir+iUNmDZmuiNcQaD3SOrV/xy5ZnglaHCyHG2nLw3Ff+V6J1mZpFjfVh2nwHMV4
bjELwGKylALwHPd6TdAjqAoxlLo+/CovoJ+htcahtqM7OJm5BybStMwr6soIyVaSZHWhjxJWxUau
isTL/hoojxNL//u2Xz/KccRKnS6JkeIzuVfdvCOIMaPQ/WKO61++y8LQ9l0wxGnlEkT8TH+4tQfm
euiBV+3enJU/SK35cmLCmZSLwMVkBFoHVot+zvG4gUK20WQyHF39rJMpjnN9cV99jMQXmj4bij4U
V1zm+9A10WqAhSq2P9V6mPaYYhgfK9PS3iOJ0WP9av+fliff5Zc9S6pRC8UG5XMoMlb+pRdO7DVG
VZJbEHczNqvBln4KMMsA8MKl68mboXB/WaKe1geHFt6zAFg6ipc8RAEuImAjaVV4eaQH1RV+ZqLj
jaKJqSDuGlB6uFRplIo85uGtkLAe/GVtuO6DVxDv4mTSNoLZD1HKlzI6Pay4ct10qthFrx9LENG5
+OlZmeIbJmzkqdYKvwmLXwHPIk7To1WYes/JxOClM5h4IAT78OoYjJ68zlRWrPnzu0dW15IgUkwQ
eQGXcBpxbr+rwnKGvLIS8yg2JQl0qrETWNVU8vurcEg2pycyadwxUlsmAUexxiZQ7bCgMxNCOy/M
ZsIQ3ahLoLYzLFJEgwykBKJrijBNBnRGo9a5XCmy52vuI2TITVMWKlSQdRWcjPsWuBViy/YSDGxU
mCNphyCvF3UYuTrF8xTPOJaV58TPulvwN1v99+pJyj4dNKUz+D4I6EaPfZDy/8uGjMs5nQVWHcgV
nm8Uu4ZlQZ9GghMtfBReohLcPVn924ZSXus4w8yWqeAw5TG3XdPYEDVY+VVwUbyRvg4JxAhoYUeo
QmTcBY+fuDQ7X/UNXmcrGPWbVX2YMlRImyJr48lUBrZW1+LX0+ytfqSvo8/1qDmd0YD/E3P/Jp+O
WNvZ61Z7qRz5T7V1MPZJadkqaAVRLwdn1mRHPyvDle7J/e8LLITYbrS+nsXoVMD2yp2rh5gA8lMR
05t0ZpQrQZPFgVxOZaN8ki0xXKhKIV8pqs5RQxAjHmTIMKyeLS1gTeXR86bqrJnzx6jLxRTYvZnL
bvob71RUVKNP5S/oMJVi641R4psGmA+IgEbNR+UFFSZBi2OWj5Qcby6uc/grsos19CWdf4G/MpBs
kYckn9wXUKH0oYZCdOJqmshBtqXIDrTPZNog+18zJESpNOeM1PZ7xXTWpa5MU06f12LPsAeALFpy
58Kl0lQaBuFt0mTHlygJ4nRNRCVUcAZSkG0DOwOezPmwfStz5fnP7Qq8uDOwZugsWl2sw4W5Tnqj
2QXuFK7ANjFU+aZ71CbqcV/HkpMSU0iguwKDllXCEjHxpmfUotNcClB/swwKiQMkEpXdWsjquMQT
irn2baqc10gGGcmDzy+Ab7qulqUUxvWwxGMjJ1dmmKZnbknl4aama+iCM6ZqmYhYYrQXHRqGy8eF
Qlu41OBIpLLD6SM/oC0yu7PpBk07qxTCXSAbt/6FBJFRCApzUMgSVY6SNdDNbYjSP41hsnocKrP0
TtY7q9TfQoSJT2PIowEqYGFBQYx0LuHWfwpXv6V5/LcIWeWG8aQQ2Zi6tOJTEaIDp+cx8XWQedg+
rfCj9LnaVJWnCQdLjDDCSFGyjRKw+j5VF6CBDu+Ok7T2F2OqMKjnqT1yRNj1d5sdb7xjgpAwW79A
Y8SQk5sM6kWP0chf46PqIwuIPGRNavQCz6Svy/RizcmwD+JtYqf4L6mOpamtgBEzAdA5AtreQx4s
4WKiaf6LbjyXXUqzZnjvygCzoQDIpPXDnSYatfRud9v2SH8nEPA+Y45eq0qqljd5bseSgwYWaxAo
knOgp7sfgXpPldQXDLHUdcLY/QSHRJ5z2KJTOawgRMIgr/a97hGYeFokBdeMQ9/uon+t/ix9fhy2
VjwAqPuocGzWvOBQZCbHpAOi1mc+MyHOKip+47qpYJMpXVMnpuukDTspohT4iv1SzsjayDZwWzyp
L8950Hn6DlBSp9Z8xmKI2O+fT9DOszeZd7qozKvXpLDcI13Ts2qK1JEKjAbi/JMX2KdyZ+1vhASx
VrI13szMdQJEIWwvk66VMTZasoO/jsVawfY0LGPHei4YtJZWJaJVDzX2HBpwb61hzJymnEGcKueb
Ys9ADjqk+TdATzBvfIZbN/caW4ogoANZ+YU5TEKoAo5tMlJCgURjujTT+XxILcK8hB+KZ4km7/Ed
T70khS+D2A+/kBxbg4w6OV6e3Suv+JgBJk8tGavPT/rdL9M7jf5cZheK8AOW0f97IMnL6zBYsAWx
R0i71Rjx9QsiBbTeMQZDc5l6+qUauZ+h1rPHXaqDILuECqsQ2yxjYOX7suQsRYYqppJ8XSz2HdT7
tkzRelzmt+zU7OP+SxYHXA+09PLKolpBLw81BlrO3yku0vNf/Aevib8MyDDaYkdd/6DO1h/gXgUG
8PaVRPnnXo7ipUB1knfrwwxAqzIvaZmllAcI4Dl+suZzuq0Sms743nomXKtNXQTpDF5WFUduY0LD
Z8USzFBLqCrWJeQie8D94ntl+AlYhVWxwRvw5cTsSpxf4m2PHGmox8Odk8M9/exzRrSmVXWcB22z
pKgsXlxFOJn2XT94rH2kDTGEoYFseEorrPxfaOska7KMm8LhZp12OfOjt2izFda51iq6Ry6oZ1es
iB6Z4FZKTSvjXIK5oszQMgcMH5S05yutfK8GLhi8z/wggHp8DVEILD9A1mlrHZqQec8LgZ12X9lD
DGnOOtJ6pzKUe21nAAILFbnSLBVotfc8pwvn2hBZQblPL83TSJEH6Bpb9oNs2zkRs9NBO7qbplrn
ZX0xuEK0Y3pJmDNBXN7if6FKV7dP0NRrldY8rsUbGfBZrELMlMODz5iboyE1hz79b+Q2hK0+OvRe
1h0NkpK1R4Uq0vP/TPIXHPNE1+K13Xikb1onMh/8uVqZbnJyc0fKcPdLUiSfoiTzjeGCw2B9uyX+
cB36+PGRtQ8bKsdGFOdVvViDN2hmRiSFvDUZ7ip9/7b+IBEcF3OjXZX/KX7H3SNYbV8tZnD8kk0z
kIADkcLU49n2wyMhVEWuKo9AiCyTaDCOoE5bxRUlaqPfswO3YrnrTANg/GpBeJdeZZB5qyXXSc+w
MKut6OJBkZtLMNhjpb3CAXDsKYu+6NoNOAT4odkjTtM2QZ00FaE6zk/nUqf8wfZrZogtRoE2h6A2
SBIPxpexHzE4Py9olyHdO4aHyRDJu0BU9D5b39YszJjKaYuH3MxCFwJh7umMRVebGXd98++qW7Ku
29/LXSskFeIc3vUxeMer9wyL59Y0Bvha4cjo5ymJq7IPHnUaTsRnYGsvZhXWjior64erIDJWh+/Q
UWr5ZZfPZv/43YEbZdzge+sYq2QDUqpBV7GjnzWxltCSuMFXT553lQHSR4Kk/x/KuNy6t5Ed7xYw
TLsFULSjkk1L9OeZpdYP46BE6INHyrA/M2pqj7/FYw7M7K9QBEdLd8D2/blog20ihMoj7dEZVxYY
4PsCoxmixN6I/KPu2+vBclf4LcwlSwdIv93oUICQMR8AktQn623n5fK9fX4U1+rmFsA/XIkNSGLe
mihvoPfAhijTFlhMsPPlWWmpZHL6UIR8auCariVOse5MeyqkeH7XdwJwSNREptbMAWNtGKMkIs72
I2RCSucBMtnlx9FwSfCuQeTpPb79JGB0GuO6B+puX2OPAQMxhPSpM6W1c3enS+ul5axXiSLucB25
pJePdRbxqaaVkhrqIa5TtUAXKhWFNpxgSal2jE02h+D6TviMjlFqGuSwLGrqA4qZr6tF2dS+dKUJ
G/pE9l8l4SlShTietoZ/m2TettZg4adFmxv2Z/AhM3dkrWDbj4Ofpren+ZkT/UzcXGirVqw/ZgJP
54VglwZCYHO7B7iNpEO04QkIykgPCqZn5+NiSutiGKgJFm2l2gHtKCOdar06jdKwsYPAsdj3uynn
vFTSPtnphFwHnJcuOwCcgUa51/S7bm2yRstTo0usp0yXl59J3700mEJ7D3i0ncjkIi0O22sZVzTe
xAkbnZloPBf6DEXroMzHqGIhqlo9UKG8q0e5HbKjJgnuySGYbJqgI46BkUM8Dzo1bRCLV1vQf8PJ
K57Inkyn0SKPp4ngmqG3dBnrsuXKdimIHvmk1DF5JkS8efAjFRlKjKfkU1++CCGSfJ6FqmU9mXz4
tIHOwwNBwAgqkKKMErG0RL3wuyp/ab++mJRaWRoB3bF5+1iTp8HwjR+yQfMOoAlG0BEL7hCVIeGN
Q/1HnLsUOzOfulVwXxU53g7EqbTtDysmJDu315Xwh0++UJGmEJhWAxuXeILc7kn9yZ0n011g7FRd
fQ+a4bkxq03ZHLYyI2y3n5iNXrDrKsHjqUfiLTHU0VYAg/OoReorxbsxCKbuJceci4sTz7KQmkBt
VZI4xdm0vdnpBAmdQLov6Gmv/6Z+/wABjmCqx5Fo5zJL1HQ1sFd+IV3boGaN5k/xXzT9w0EGDdwE
DZz7D2UsNnKzmRRq9rPrLSbK13WMkwJTdlABqA/j6zFgfikBt5RoGOigYOM1kYPE+0WJedplAiXc
Nuh9gNOx+qhPzx2HAXhC+d0XTJt6RMk5TRKCWX+SJ5TtSGNG0Zp8OUO73GHMYooPtAaZZF8HNVRT
7xDr5KINvZ44ArZk8gaOAi7xfdgOO6lV2rh11gtC591BeHpFEfj6KQU5tJ/P1Lnf3uBfpOD5Zizg
YxwXerevIEpE6JU9s1VdvZ1KGjXpM0EL9cKqHqFwZAK4bpqvpWW00GMD+AmpUzBeS+fEe0bhpvIT
VBuGIiNyzrmsN++cVx8h8V9O8OM2DOGDXR9Cqi/1ubvinCVxflMYRCGlT07JC2yJTycGm9C0W1zO
9CLU3oPzXu8KlRYmLWMZJ6d4l3kA0/JQCxH7GbORMnZtYzKZVbu9zK6eISMJo97T3sUu4pFlOSZ6
2ZwuULNmawtdmP0ZbW7fPosXYkURRlH7JZ+xAQfPOMjRIosuzY4YNmnGzrShgbuu2r1umDo6AgnJ
glFB/fYt1H79sYwPP79NkoaIBsKAd657YTRoLZ0VGMzzr1BEz9E+mNH3W6+ofQDMd7BMLjQQMzcZ
wr61Xjx2bO7rMRMXLm25/HJH8Wahrjzpb+6KRxq6X2GUSYskDzAmm3y9hN7PTU8XLgh61C1iTMgm
Y7FT25xaGH2OpTAsziZMaRi9WchPuKnIWg5OvsNpQQWxScWjUyXjbwtunD0whn454krrDB1dQjk5
cGWhLuumfwdtvxrWyNm8gb8/s+mX3mgKjWFQAnA8dbYlgM+suNRr1GNRDgYsbS7Ckws4NuSY8VdL
4ETSusmspyIDfr4L2EMKIc+yqN2j9rVEVgCldS+Zir19VnPQF5dxw9P5w5F/8kBnL7SvonV/ofZ8
HH+014RJG/HU2F0w5kMUcLFgWTOgUe8oZ4CATruFechP8emATDKsMLWNmo2Tk1pxZ3SJXMX3wO63
vNGBH4B5tkhq9WARHlHySjpeoVaDlgnViAawfv+59wI536e4DNHKsRHJwhOO3HywsfcCekhHGzjn
SPqvSv9mRvjpQXo+WY22FEeGXxx3ANqbblj47hc7pediFjR99YbQrta6eKpHpgx/gaEE0OlZGMSy
EkZxayeD3jA9/QUQNPQWmqFIOR5/NjBBKKazQtZZAdg+kjP6ztlnBJGNi1h4EWgxK5cL0fpmvilL
7/jfCOBwEb/oh/O3mrqJWMqBiyi0i7pH5rFUcQPGRUtiRVKI8dCvnwsIZHQl6rphhk89a0y8IiGU
XPM16xAaheAyxHM2HG68O3EcXNlg2PPBnTbpuey0AdizJPQ4vgW1H+Uk0A8ecijrtUoh39Zvmhw+
6QMuLtQzweLms4jzb/LvSF+N6ONz2WjmTgZ2GkFWAl6SBm458WUrLh2UDHMuc1RG/DpLRM2wRv/4
P8e0HUPVX7ykpyVPMKROMCuDX5TQ1oobrRSDUGOMSpe3DZH7FtkaYsP+fTgTCXVfFs7UaqECJ72o
x5wz9o8JoTwUaNJ5aQAkX34ZoJ6Vyv3EskMjQeQV1UfRK2Qyg5HPNdUawr941Zx5BUYuvzCaJmMr
i+T9H7UQIOVYKlBsHvLm/c5gq0hQM1vftX5YY6ntbM75BF6n7DKvap1o0zE5n4z72xU7JaubxMpB
JBLl22ANESuDduRIAl8efKbeCDyWC7h/weTwc8H2bWGnM9RyAbQqz3s6bLgH7hWv2P5B2siq3Ttk
H8dNH/rDmBwMle3TxQ8PAQXdwlxCKFnVqVqyOxTM3+PcRnkrdVwYVFQBz8YkDa4eFRF0Y7FSvena
Kjgrcq+RNS1ggOIkhDkv6bHMX1HSCYfRrnGh43Y6MPMxPDJBUC1Lj8xegbjT3KZzC5mnqEvpnXY+
l/6Twrjwc0HFuHcNMGHOXIkQVq1tFQpzInA30zIorZV+V/ts31Y6Qi3z9RvQB/S7bS9AvfoRALOO
Qk3fjUR498J2HRZFKTJe+d7MRTo+sXMWH7D0LOQuj5xBYHvJu37fnucqmp0ZvcSSmYW85ODLkR8P
MSeW8F8vEE/56u4tBPUPgcV8J+/3k/Ao3UGc/rulVd3ckHYfOi7r0T1COI86I/+jCso5X265L15k
NKCumSrCJeKawXuPibYExKL2IKpN1yod1f0rnvAB1BXC2TN5Ezsust+st+31OAFdbroUXgz5LV/4
kt1cXVcKSxBTgu5XEGP3KVwVl8/DvZ7xo0GdyoxCE2UOt5sbGF/DDmWnE8IK3+PSByZcHkcyJ71v
u284Hd3HStb51sxj4KnQoMhuvDuXaLev0k4ARC67cQezS+5U9Z8AFA2BQMEXf9YBsCPsPUt/w4yZ
MS7h4IwrggLfvNxX1Fy78PaJ15arGTNRrHGf+qMkMdLVqVwukq7CHKziyshHPXAgXGdwNKFpGNuV
n/8npXtPsl4qfKEN2YQ42ExlA1GjaE4vM3qA1zPCQ5TqEmbeG5p4RYWHAxqZDyQwNXiiQlTaqncA
VJqm2OWjEm0/EJDBKs5F+7aAf847iAUi8zQP2QXEUtH+5D2RJxu28YdsIiNyR9DLMk8Qrjtsgael
EhfhgTtOERw/pUy5lRZ00kq6rREWGg9F+s+FehrL4kQafzuGdTa75ZkmYzyDMGcoM1h5Gk4VrnVi
dLjgqfl5w5MDXx2q5zH+YR7qXoQggED9PDCkrqmF3wn1tKbYp9sET+mQVpGqeWhxusYpyqkLWgh7
WQz5Qf1g782OcSEuN1WZuUbVaOjHx8+EKQyi8JsQLOzXRsF6zmHW+6lvSC63kiqQLqZQGawS9aPf
U2ezQRYePCtzghbGhyprjgm0cYVj5vjwe0ceZ2P+cP+tubOoK2EfYvIFMYsct4jZ1Jrw6ym4Fnq3
mNskWTaUPjLHI1nSeiYJY8BKIrpk8yH8Vv6SF/Kl6FALKaOS4wKYO+Ae/pgAMvWQfWbmU9SsdS1c
Pmvp09qrjHMw2jQU21iaKmlzsGP4CgIzRTTirpEkFNKSr4U1VFuBkvceXOAj2wWlUCH5B3/flKJ6
5AKZONTCpUcwPf43awTHrC+GJDSRpOnBWzsoRq5TaRW8yL37nhjK/LoMymKfWmipq4S3HBLLNfs+
idxsGbPZ6cPUXFXp0XxmQu1+2ZBTNOvvF693V86oO4jAfFs3ixkI88juO1KXNOXclCdHrPErPtIJ
/fDEpCCbbgugFbHIp7Bowld1KqcdPSN4FNyD9sAUDD1ppXt+qeq/oFzMRBsuit/6c2tk+CC6tCx1
3Lpi1ZIBBs7GQqSrblnkVK5KP559qH+Fwl7djgvUqqUBFjP7U59FqaKmR398Lv3NNo++HiPqKfy6
+hpuIV1A/MRe/T/7hWsWz7iYtBNPF487RIb1+dMEzb3LOOa4lKqWA15BTkEmbXMJi80cblzWvOVv
cQNF4z6jR2V96gqXjizW5pB67Wnwi+sGPcDQ7oHhCJUqJrUt0ZRfh7HP/TabKN9gQIw7I5Z5wD3s
ZSCAoqr5+z46dNXSbm1QDV6hYRqhQZg/VqKWmV7NNKC0hTRtdi054rDsrZkdbjo516okWLRQJD08
kdm9H+KMUiqwm+hwZqAR9lkQg99BuArDR4lOZLbi12f3FC5N8tTlHdqD+1x4qnVZv9e+ko1dB+M1
Kk5ogwSaatF14/655ZTlcaPEZ1nf6Q5z5JnpIEMTO+C19lFu2zJ6ifLB2qXr4WH+kmx3ggCxSdmp
dSQMNOb18Z1gsvXjjPyiyP9NpU0s8wMja+rXls5kCQf6fywUi3EUeaiiC5zx71bX1OUg0k1lCY1q
eQW+um4PEPQ5Pijz74GQ5htzBSMX3iQ2fa/qb1jQCo0U/92IVd21UJc/gqE04vHHjinqteNYLeJl
W+YZMhCPGNEKC/+RTeV/oC69WSl/B7rpW7awAPLemA25J8Pd8+rgRRjR7ZzeepSDHoG912L8s2eI
w8elweoGvGB1VAdPmqm3uIioZmvEd9GyoFIRpt3ZZI0zS6sm8J05jdjD0qTtXG5FIry2gNQqdx+T
jByOgGe/17haSQnm5TEEsq/1OtjTu5V1i389IIbq36nK0R0x/giWwrAzkGdicK/oz9dcRtZoD7TH
SQXegE8QWN43KdVMyZMc9aEX4nEW0vo7SP4kPT0eG3OgiqSiLjCNTko3W3JMKVsEWoS1krlpE7wU
BQQD+KviNKsW/BHBD6YCQ4DA3n1z87BxNutYBWLguVcv8vSxM8VOFLrfV3rAYiMDB3rKJc2IRAg7
tMk9psaX8cCC7LoKpGdf0SMCcqYOWF1Kt0sx4HJCfIsneJtViZfvimoFjC+5URmLYl7hS+62Cklj
VNbm+JVwpfGcKSx9rJMepUHpM+jJjaF1BdY1NQn4qIMiOzy0nxW5hUWPPeJ0nV8jqf36sO/XBGa7
/fyoPKFSFwEOSW/ke3b49las2F24Y3iZQcq6Tjyv7fAVB0IUXDqq3IP4V6EHoGwH8VIvRX84JKEX
L2lugd5Ck1n1GM6LIOeLlezu3TiFEgQYrbOxiucQUhxVjpfnPc7xiAnyjvAv589ZoYoLIQzyts7E
IrzYbpVgcnh2+LbHDcYCIVnkNQv4G/KPgWWuXq1maKjJH5aVguiqEVa7DATYJiBDNPEB6pXHQIrY
Ck2paj3qFYvuGmpDEzI4tsJEkqzHRIVYJsaBwFd8mZCvNsffKjZ4bQFxcozjYrr4dMByVK391cZl
SJd5OakvGMG4PV3Pt+/5CFzwAtqUYE4ZmVVt/7t0Doz2pPjSL9xbWdAOzn+wXadfFEy0xJX9+Iyk
/9k1Xf32c7ymxuv6Y+Ak9cd+11JLzlP7XtRJCpGMFyXVYxFKw5jgSkRG9Qq4kslCklCBGj7liMcr
B7NyvIGGaLmlvPkyTdsDS01jAwEwUY5MkfoJtN/CaCkvd9ImP1OP0e6BnDqG06OXe4QMIKysUmZ2
Un2fumw0Vpg7vteqYV4GOi4UyxiLhxhD/FZht/C0mnaWbfiNeZQWPgOimNqz+tFFDJF3j0NKIgPg
s+TY3+SIABay+PaFnzEqE+5ju4ePOkUIAvNztcL/Vm0Q4JoxNyZTY8wqtNHgyXm8HnIu5YkD7y25
CNR8xZ4LetdFVV1MWdlJci+nASdF+r8VKFvrewhFN2XB3G5JOotdpdedPn80tPiygwm0KBQuNJXv
UJI1FP+N7R6YFhjTvIj5DJ+KJCLQvwRC6f/v8uU4HxgkzVo4ilo60y9yrqOh93UZF0M6zqJ/8OlV
dHJFAzUjgy3anOaWc+jYNNIN9D50Vko0IqHMZHJQMwxYRwcnKsSavG/gAm/oHMAFCTEoRH5jiz1Y
UbsCgtJJHPWaZZL3BJ3Nm9jz4h8VsnufAfljzvbpFnZM+f/w3pGHyGkXAPqR7OQiZQN2IkDDG2SF
p8IsZlHfg6gCjF4s++pvDgoFLQ6kiJkjQSuev+iHPqcYbrU8PzVlQHfTSwGoe8A7MwSqQy7P7UTB
u8HIOj1+k9vRva0nv37ZZjzflnGQNXLDDWISaK64kZ0xEjGmvOrep2ypKodIEc5XwC4nqkOiftBp
LUn61ubljpQM5Sb/huPZU3z17TjBoCsIJUW5QdOM7MACvIB/BfOieHUsQSMcjKZiUwtXbcYf87sn
Oqgk3gybIvP5W0NeiL9jJczwucpFfJmALTTVG6rizp5djgvlDOn8y1RxyV1DxArMddFXiNRdJ8EB
wQdHVburBAxEZ1fVqQDmhTu4GUx9RP6apNdSrWuvluvsux84Nv3K+gFJiDyaeTmzGi/lYtZaVRWM
JqETPv6INHnTsVZHCtDbk2p3sU/QGGCPTl/DUo2cXgCCcY6W9BHG25pBq3dY+swZT8u/7vz6/vwE
tcJVDAAkZL6QgkhnG93b+WW7z28T5wH9GDFCfdqeZkVS2whU71WnBMTtlGBUSm0BwmcmwNlG2gLS
gc5ovPE1IS8K6CyEdeiYRuumlcsw+51ttZVGDSp9CZ4OGUTTi/LKAnt5fqkwhGQgWlS2jfZbcCao
j5cU0awuX0SC0PWhrNpxHQV/XE1J0SVnsbF7HuCjqjgoX6GcOc3lmh63rB33SYJUqvhz5BbDidIb
GNd2u0XyUH9UgFjdReOxIQwiqB/bWKUxq4opGe7JDlkyA4gscHMLFle5TRF5csla4dh7VRstO2Rf
7NbfsvZC4oXlZjap68KqAqjEk9ZxqGeH1SLEtzmNXwZ5V2aF6jvRcgn1DLtMI7mSz+BBo5JsE15Y
hEVsFJ2UeqdDwilFSz7LDOpxXXTFhQMU3Lq3ZEnzgcsMdCniZLFoAzHOmH+znKB2fAUYU4N4QpxH
g0ghcjC1UVDGaMrJV4RYXdypOGiZvLhDqB7p9RpeB5PIUjWcbUJVa2rQBxdBv844kmR4dhjDf5ZD
PCUspp8w5JQQOcW45YkIdc5TZe1+KFm+HV4qBD7Aw1vcXITwthXW1TpwAOVR+5iFp0E7wew6xgq/
++y3fVnnFFTN1AfZ9SrGcp8XIUsgNjF01iwgI1sZETW3j2goXisadP1SrZXweNDahvjzSLgZol0r
MIXuugjA3S+8ohQmoA///RGJ3Qgd9r6ZJqCi2vUMoH7jSOXfdvGY+aVpHYofg5WQaEHg5hyWGFZG
X761mobf0yGapucgLj6na+WkjNv8RnRcpFyR8l/xWZA/QQnQ9nAn55sXHjk5JKftXFwBAtiu6Bjy
g8NKG3Mj+1hCXuNvdg05rs98O6W6vz06DeddotPfkaGQtJhUUjoXEMgA8dysEeUUT8Ajq976FmTJ
HZ1Pmsw62VetqZRbS1DkEJybVMIc3QH+OaagTGDfiLSvbZ5NljJKrcNqGVZUR1oWT2dd3Lt0Bvt8
HD8yc03wyF22QWbNMuUhgfVD5VFQ8yMbqy0u770fUgkvqulTNRDzczY8Qr+DqF/hbyvHTLyQVnc8
DSBEUBljornvtaFxSH9TheM+GBUWFN2JB3GqwC1UwtrtSFRNqhpgaS+eUxYVOQhxaBBzhAypvXap
5QTQYySu4Qmlv15nbfaqUW/Yoa3ba0LdWqIAGGKNqSSYrQJ5GO9QulweHzBz7vtTs8Ak9qIM6Wfj
Ayrvpz13enkb6vqRWfGV2MmQOPwdwXjbx66ixEmoQ6bSe8e1KdHK5e61cHnYJki7AmSzHgxO44ru
r5k8hF7DtZb2x+pokmRUv0VB7xHEDnVnpNCPZ9vXWvDtRMi5YaPc1I2vzxfK6lA/A8mMb8FXw28F
ie6JPMvO0mcBivm98++IWAxpzkNf9jbfNvnGgl74w9TsZiD6AxdOavqzs6af2MgRoXAk0s+VJkBL
PmMMV+Ph6z+qRJJV07Yqo0/COfEDlbfbTy0kF8sWg/RSLYTmZ2g8PlvHqfP2yOZQj552p1UTSJV/
eC2pew1RQ6v1CxXVDgYDpnPpLeYG8zraz2Nr9lCK88BIz07npWZfu2VTDwRvlObAXKB/x4vD/kSm
7SPV8s08uUOxN9mw9PzsfbIDOy5Bxl9LV6zqE+Xcjt22zKS18WWWy7/2XlPfcrNjLUVad/hpFTFy
BCd9c4773WEfQMP1ie+whTWB6jPRvLWvoK56vq6ShomS78C6nYrTicF2zfKjTmQM8FR0M03A/zj2
8XwDg8iIo5idCWbYB5XlQIbioM7bfF+o2iA5nD8qEVE2a6kgbiQhAvhU0CA1c3CDHoPfPQWII5NN
Vf3h2yKzH39ST7LJccHLQM9ZNmvkseavyoXmve1iiArw3eyIPcUSF9OxNT0pVsqFkBOg50i10drO
FtTbtdE/5FN/ewSJyVelFpm6ra/ZZlRNDftEw5O1CBDlwGx7RbTUCTJqgSWbAwHJQ7phIbKMQB8k
B/XK1oYB2AUqHePDCf/TjU5qxuKY+a7wUdRjCchEPOuBoOyNgqEkaNIPeDtX9yPnGPd7KbKmIEvk
Up15ssS1JnOi9X7Y5I8YrQDrRhzCLenPUXDnJznSdqG6AjSB4sn0xYMekAuh0aMyZJwwV6lJ7Cm4
YJX+T6kPBiUcl6Ec6DrIjhDCyCO3Ekt0G9k227ALylMVUMOXok+CIs3mt+hdyWSsk/oE3tvZS4Ua
t/OPm22dsr7Md/fuTvEFzZf8jBtY6yMnrVWM/9umOYbztKQ3ZvL9xG5PkcbRmXhLa1XBBVaLYxD6
aDIFsyQpTR+E8tQhqXpMt5yKcQ7j8vjJUmH8B1+trGDW3RZWpEB7PjPpjEKRgBnb/5i3jQTYLfIl
L81CcJIVuXV9mxoyp8H8Cq7tY9IovCQJQRI4t2S2Q1AhCUhaGtIM3waKjB6N9F292Cf+yDbb3fQS
BtqSe9Va1iJtScNARctaPhKqp6jptFB0aggNaYl/rZ9XiSRN/JB7ebRKaD+GXNHECRMZJprn5RXD
25JFZpgUpoRH+281ksg3cx84qZRdv2y2OXxW/YDnJiD0kEt4Bwjy9WLOfJiPP0CFiUSRbz/rwZw+
PUPlMy3/O6GhH7jO2W0sBbIhm7o3Q1o2vs/Usu+d/xDGhaGf1vChkEjMajdTaODt5zlvXamFKuyu
SY8FTEnfCzXVxlmUdyHlSSh9Po1S5zayFx9FGfZbH1TCHvURJiuUIDA0RhDjBHtlaZZz66xSkC7x
wuPFaXTbRcZXJu5HBYhp3DEKTeAnPWOQFPbPFUHBKct71jhECEPOVsleTB6uS3pJrTKr4la8hODA
v6as2ApeklEMY1oLEkjDBC6Yff/9eJRGhTIVvcOZNZqA8IfA08U41e3ySnaf/w5wvskB1ogbm4Nf
UxOL6BrSaQ9x4N8ouV7PjM9OChdL5jTjlE9eLMvrHqCf/uz30JzPibw6Dt+VautHU2bI74dzb5Bs
ogexPrT+H4v1IGFrBOADGFhvm1CqNIzlkukJTzhux2IxtYt9AI1oqPJGTetRS9/CfBYB0UiGRRlw
q3tucTpvoW0bab6p7YcyEa8x4yKv+dyfyPxo6VkAl37rQ0qNljLBM8gC2E7UOPm0/Nkca+/oHSz+
QFGtaM2IAClyHCX/IWYd6vFzwlbFrgKHSZLn1CcgbzuhPhZn5ETJDY2SaLtTtevof2hm0DQSXnI/
EHquZAvBQwXrSJ/aGAAhKppr05JqtgML8U+ROyL3fP7A9EaJgYd2ya9YfiHUCTSA4mI+s5zWt3Gg
Di2d/h1qrkaV7rMANSUhTgEgy2ErCHdn6Mc+sVpwOm7IP7DogdOFqZksv7RLdphB//J4xxDTJ2B9
/E2xFAN6LRaP2tZGryzEiGmpFJqIXwUQi7Kepi2AKAgj9MyiVawANNriB0Vrk72q6zqJjp3/+NJw
nJ3lxEyLgydoIbgqojOe1A4fcc1HLHSSN8S+VfS8055PfeWnhqBf2rRrpbCb88KD6sHsuL07sANB
Fk7s/LIlhQM9ziWvS6APnDagoImbBx3sQ4g7qi6pi03YlcP9qfodHqutTIij+9QzDblOK4Oq6vaB
jl7KIBZtDDgp4ksgvoIjQGs1k7rgsM6slAqLxTxcavxfiIEY4LQRjOSo+/mlC5c9PpVmIlyHo5BH
yebw5Pjr/jm/UbRjm1af65qWW5ManMwtibRPogDM8EkrP9sqbV7X5D8jcZZHI0OKu30EqbYL2o3T
yvZ+N8XUnx8KhteLX9nZFd/t2Wd7Pj9ZEnQzvx7nmlGQhhlrlxeJsqftTFUVPHoqg3eDGa4mJWt7
TEYaZfpzbwIqS7qXZQ8ClBl0m4Nm1xPEzOcA4olQyQj/CKXclQo1s4DIVGFXz7seXrB4HXJ5jNZj
cTPVsQ0GI//VDcRxcD2w4kYAiuNberSvPWdBDCN2tGGaswHPcP2FQUHW4HadAtoj0qbQXifHF4ug
sbf2e1/LumSLKS0MdKrgmDgx3qK04i1Um8Z6grJRgQmAEP/qtheRsofZoohuEanejY9kuPRsGUFP
t94P4T1L5qlK7SrBLEezFUKm3V6Ha7/h7cmjz4hygMxi0wkfuHKu8ZLDw2mywF/em5sbnB/1c23f
SRYcMoXq8l6g58IlTTVY1EktNSoeoB7iMiuAJxdee5vHM1AQcAOFNCS9Glx7tVPNemTE2YZIe99Q
GU3MOWjmnGYCjTaxRqIA4KjmXXY5iZr7P0D771XmzCc+jVbW2UByxFqPq7ptwW11CXdU2hPag3Mi
/JuDZ+4Q20p1W1Nq+AIoeXSjdqeIz3R/wQOfC/cpMX7kMLwXSWY8oOjAOAo2eyfSi+PCVKLlso6w
g/hW3wlMhA/mNJ6Sh4NB4S9sZ9TM3aNZkXxS66RAiTBcYIaWPYTj/aRPsd4A/08YstA0LfwimQOU
p/vesYsST2nrVOmqp/jLRM1TqW6fNiFVe3VMDG0XRg11eIoxL3f0G2bkA8QKulTWJaiG4o9FWvuf
bbNAOVYNgRQpO+/jDQeWwQMy6S9JaR5kx5IGIwIGmzgwu1NrtJJoB9+AZOR9bodydfGWo6n8JDql
y8GftFUaWl/dX7RJdSMqiAysc6SxJ4aYWcaeup1np4lTuEdPFrhttUncGar/Aa3ZR1b1MweBDP5I
wkh3GG/mXOFcvkBQvjGVEf3ZYfgNYfGCJa5EgcYL4IQBF5wiwyowkqEHLmfc038p0G1chpLOsf2Z
MXWaRpsXh09t7qlLIQjIq2ANY/wskVgTE7xjhl7XK9OhSN27HaLUv6R2v3JWi3pOne5fZuAZja7/
x0M2AaFpDfxw01LGVmqa8LKLAMD6VTtaWVcoZA7WF29wLIdQsGzx9jdV9LBFgXsvy/E9eHCEspVT
3rX6P//h7DkVkKjgBUdPqFrvxQ9mXauzftytlj9SZmvb/Q2j5Ck/zwFmgG6YNvbc9x9c7G6kIVU6
xPFg5B2ZYk5bh9aGaLRTpZmVT+fRAm5ABice2gg3+URNVr/xr2OiA6Hc9lUkA8MQKFIoupoT0FwX
48R2dL6KCYsG71JY5Caa3FX/9TfJzpaLtbpMqX/0IC8w/ekCKN6M0zjr9dCMEz9cZwpgM31FWGCQ
60c8Od/LdSSCFzD47uCfI6t+i7DjS8PqbTmAoZuMOEkl6vw27xKLEsHB0Z5CQkFFdFqdEFKAaAm/
Keh4stjsCPM5dszNHAbrdY87VMX3rKpxv6LJXGe3QyV6bCTMYmSs1+txqol7r5ZyZ3ZDVUK8vEnO
ifRfdZYesE3mPaDZPhNCgCJaNZAYNAO4Gqrdvh7XWKI1qqsFyHF2y3qPeF/uo5rwWiGeTwnG8xCP
7unjnDh3iV8yLMoPulUOWS5rUt8XPdz+4f9+e5AIKoc4LqAs2H8y2D8EgVrSWTwDrl9etLE/NYFj
gWIlzYawaqjNpTsYYoqDsqqmIo1CSfo93irNCwPeqZGaYyYspigWBRuCrQas7S/GVBS3fWTKDjWv
GV7Y0ewSEoGmCM3dEg0ERRE3qFeVaKHh9CGE3gpefxFa9Q/6nyeRu5caz328RShvEHn8uLThwqxB
F3Hzd10sXRAlOpi1YuRQyN22jmcOrXmQmdAObaP0VyAo4RFd1jF0DLpvZf5JBogBg+ozoxxvuoav
QlIq5VVkb4mpKChl8YhxuD7uk8W4akV5ROVWldWHt7Vzdt+UERC+hXicbQnkOIVlhz3XsxQrolFc
tqvYZV5/g2Y2LF3GDnxVH8Ef2UkwH4gSclTYhpvr+Njn/zP+RZxbt84vUREws9oOPvLugkEufmdJ
CwsjSP04EDsRwfTtKajJiHTAGHy9h+ieKoeNDG9ZZGg1F6pnim3urLH845EJv+jc0DgmJjjsUfCf
DgKAEP0w1uVHLjPKqfbA5TwhlDP7rGjTUwVezD9pPsk4kul8ZoDSgi5ZTDy8aMHIEsBmd+Nx+DtT
CLdA1c3U7gAsjiWmuT+hIpYa8KcTPzkmeCF7U6zVyiEOb4UJ99Ddbs+nbMcqhT6z1CELNKudcT5e
6xUltRMIwMI+ru1axNkrjHRX7YTyEU+xVno/fJiyW6eSpbLNmEkDtVytRBLRPBelc1ctGG9mfYu8
A6wF2zTlK6OrF3Fe9ud2TJbguDLRy5wlKVAtv7NoIryIu43xur3CEameEh+iKiRWjU2Yza2jHzQn
rj/x+4u5GnMlbfXDspITU39ak+SsqxqUedENIWymgSh0CLYHwoEQT9SObow3Xr0BaQaT2TmSLo+c
WXsypa5A1QlRDpqNGext2MXsEpRXvf81pRM7NWOJUaEeaiuxUNFGGiQJYA50i9ogykG/0vQnBgLw
bqxXEhAgQoxGmJkLT3h8G0nBqTc6ZHzzqJwKcHiST6uoxaqeGI7ZqvHKqEVId9a4862ZUPW/zJ6E
VNcCw1bgyzGe+jpifmY6yTM0qQ8mcHR0gXQwujLSa2u/AalFoOhdGWOJTfQnka/LvlTngGIcL/HT
RGNsrn8SaSSjEFCHj6yXSEkUR7J5/vIZhGG8xtz54yG8o3AWTcbE03alpneqGODzsKMyUloSeGAa
d4Eva+OyKvSqOfjZSexygPoYIS8jfKWkRhF0cZgbomyzUi6sLbW1B5LNga+hRRhBtbFRQINhWxXS
qEoyVx/AXl/7i7XjqWmTkGwdpUifg/xaNA+hLqE06ZBM0Mirk5skvhY6hXKaXDap1LwA46oI94ac
VaOXSmiHn2xqh7iaVb3vZw8iSoJG92RtuQ3JWi9g1XAR7QWkIYEoVcGS5xGpk3CWXwM+3yFLV0hP
FQ+XPULWidDtBXh4ggSF61KbhUg5g9qwZ9fYr+vSFE8rpObO2imOHwK9yJw74SLGx1MrJKn1jd6p
bkuPh4jLH0SqEjL5CCL0JoLCfJek4SoQ5F2EpS7G22it3VNf22hg2upRRfCjM69NcVLdJRGzUFsP
sN8F8DfIKn+6ycw+hjWUocmjSuBZLEGsz4RWZOM+Z4G6PY4IeNSx0vTCihPu5rvW2PDoJdK9Uk9m
hl/v1weDBjuxu4L2mRNxpENhrqCVLCBUdsjHzGKVha0nLrA4B3luUdyB9rIINGGKE+ZSget31RbX
vBIfmcMRD7EagYZunH6CCpS1z9ZCVODSlI9cVewZc4Gp1ryu71hPCsAxCrjcbAGesaBdcFp1gVOB
0z1e1UX7rcslDf455ZrMPX3IgBwKznJWoIGzjb8LJ2WmRclo9EfHGUpR1V2GqxWFcyvOY09yHPB6
1qO8sGuYGlBT6VnbRwTgrRk/YZVvAefqKmM1Y7VbVPijBKoQdfWbk/nPTT5q46qrwKsv8xuUaTGG
NhwV8KvlDPiTFu363bSbZxPL/1qntJDGwfjIf8cr7oC0gbBudzpYI2SDGQym6GuadtNaisI9UQww
Mj9pFjKE6fhxKfk9RnNT9ZAvru6w/E3buMcV2Tgog8bvmUjEtEIVVCikJr3AqAC+//QBAXee4lgU
Ds0V6YcCYzxrCFvQXPaPieLov8dpFMRfl61WRQy1ceLuJDE7cTfW4Xf5SSuFPuirXJoHVi6r8R6q
qJCxCdVtWlc88ScG5HdtZwGoaSitUL64mcl6uqpsNgfOdGBTuM+wXkt2KaRNn+iSg5ywUc1UvWsm
bDrAnG/MypZZJEi7lhi3fJYvvgZkhruFuOj006npxY966Blv3WO4WmdVDdKQ2ZNKGnAyPBTWofQ+
WiFKZ4TE1aXqYh2i+MwbxUUzX51q/wL7hxIOWDzes+WFbw+9JIWaj2nQqm9hHexiudyLgcM+V7ck
auj44re1OoyTbdqvru95kiX4zSSe2hbwg40nzcZwd9Ow3jEMQKRKe/6qvPXlnts9KS+AJR7fp6Gj
+EwP1UB4WIuCSslhnC3IWaF7J7YHbiYyyCDdQw4fXSOrTkdlwjhYNMkUQt5sD+bk+uVj2GGiZnrx
BgCfalo8AKiTAH8FGL5T1uWp7VkhYkyGiWoh2jcZEn1oayJHCexluwev1y99vMo/iWIUFw6jFLQM
QDupl7843wv/xW6FNtdSUWGQu4/7raxotntFudjd6kSvevQSHL0fwo8YpAZJTqmGJcvl/AV+tOl0
l8JjzdbgIjJ0xRP3FUKzYpGyZPIyblP/Mwpl9G8lc1ub2e9HqbpaShUGEtrswbppXc79am2UTQcP
wO8lSfYfCDFf80DPWF9SP4JmJhAiB/GpCVUs4WrKlrPkaLUJEVfV30Ot3B76LTEa8HwRnrt7Qw6U
THRXOmup028w9gh6P1pGV/V6bjIfsdUhnmoSDNPvhsxbSjNLa1GCMuxjzSb21dCIsqTcnqcwpwPG
pyDcU4H+bxFbaurV/ORS7dWWnTKCEyM3c2ecStJuDD9ujmLPxHG5IlvWuT5W5hOPjxYf9oGkD1cF
ccidZBm9vQSpj3R41pfRX8CKDuG3S7602sl1U8NNDpOUru+wVVdTcIa60Gg9sNIItPuYIHlDVsoQ
evYXIN12+WeGlrAoDElu9JsQEaUHT2kh/8bQj6yYYYX7DiMQg9Vr3Ap25tIGjl5jNBWkqWaQBLWe
9xlDeA5qsOEmSOSR4inlrdWH8bBYcnbvKrc5srGoNa4ayYLuxa4eGPvbwLmgGYCuywVIPVNZnxWb
QWi0DYjUSXZROAkUhU9rPu+1zlnRuANjoIK4qRfmNxMYGgMvVie0iLAgVdpfNBzTyNy/o9kqrCIs
nn5B2HvLJ3dUVx+jxLNtJJWf7bRrfyTze1FicOcl74mAOCAy3uwGmQZlui4mnuf3sPYthow9YQC1
oz+DE+OnoSRjs1176NIaxFhhsYCdo/mt5HoCJL6FjFYoCYv1FegkNEx9Ixy6q5zyaIdUjeLlAE1J
8LS557ROizOyhgfBDSy79U5G7RM+gHpOffttHwRo7h1rngzdFSNDPKiZN+PYyk1AqMSFBVlTfbCM
b6KLkeORKDw5SuslITO1a4TfvkLG1kg9B6biQt23yXgQe3up09R2waZLptwcu69yc8D40Pn+7hEY
unCy/z8y7S0Jyz4pMJsbZTGEackAaLsusgyWo1BNkvfNG9gylsnGQilRgiX/2/uw+JlSYNWua/pF
GDQVXvJdxWF4gYItettreeshB1BksMYE+GBE6PmVnst05k185wBB5W/4moX3hKXPTM03j/xYWJok
9Fe4bgEe0dymB7XmY9CeQ3gX2PJ/ztyevHE0gqfGq9QJnrhPvcCO76S5EuoYT/XY8fi0/eBnEdSn
J22+p4AP99573HApha4L+RDLeEg6eYySf7oBfUWUC1QvH4Tqpuo0E31CpQdcT+TgTEF8ThCDWIY1
ZpvzDy6Y0rY6OrMUp+V/2GE1sRnzzUv76+dgewL+GpVhiPoZZhYJiyRurjF/MNA8k7hqLVnLkvtJ
jV3NoksXlQx482YTPrInHDDtGGv1a/6StjsXimmvAdE886hCVjegtcM7B7Zx+C5lAWw8b1fM1X5B
b2veUd6GuS0nuUOE2t1iv8xcXE0JRYUr4N06+73oDha09f7JI1c4whmMZ/oBiodTObQxUHwpk1zq
0xgxWlLoMddrCjugL+yFxCsQltoNXC8Jmdwch7/HoM5AmqBSPUjI1omQuO6qjpbBy1j56n7u7whC
CAUNWtwyE5RdMpyMkvsR2g1L97yqc07lA16iA768n3PLCdvZ/a+9uvHjb0FPzdRH/xHG1/jPUJfY
4liY+A9s11YFo63T50UnNfhL2dbDenRljz8CCGe3z9UKaDORi18Nj9dxEZmrNpgv5tvlILlmvGfg
84F68+FtFhS3vlEVMJvP3HsIURaa07f3OE9I9A7qArSnoektHy2NsuuQB0hhR8ccEGImSmc0I6IX
IJbpRSGLvn3BT/YXFcC2VsWgW+yzrwbknWLj1sE2XU3DrQGpDaMRC0AqaN0LC49PxBpdzk3Q775K
WJ5sHbTKpia8AZvqAfOhlGdP3FFdI/10boV8EuSvGYkFv+89XYnLHlBP+FqWPNjN1PbTbLNEnIKg
2l+KzCFlcZ0S40SB56HnpsFWSX+vnxO74UPEA4EAhTVJBO+h0Ro/tRzZYLVuy29xSMKQqlkhHoXY
C5/uFbeSNFyF8v6SYu8/5HVk8x2RG0ccXkdF/KaQf6F82WpY072vE3zySKVj0iY3M+TOuktzGmjA
xjcN1oMRn0Mf+BCMzh6UvXeySqt79UgmC00F1ksuU65dee4uaU5Ll+3FFCZ0a1j6eLwwFWFs6QA1
lYJUS4qmgxYkqXdF90FeZjd3K6kBMTKqtImW/witlmK7L8vkt0y4Po92oe/BccEPAGb00Lk3Zw==
`protect end_protected

