

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JEmZWuLCZazscYOT+xp8tQcgcJoo9xw+tt17VTk0Ee/cpOS713F8lYXKKz7qKA5t3FpvNSj+LwOT
FOkmwv2alA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IW+w81BdrtEdSrXT08IyeN9itdwHkCyvXK5q8xF0K0oVKDwJZ55f8rUD3UDvvDXIcAjvU+645JL4
ch4hQtC7Y2FokqIuMtHZi7cNrCDQXzP1bGPJjMCZbuYkodHhhDFZq0vnJHG5npJwjfiUcFOs/BD6
321VxRY2LE90m/fkP5w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mn15icVDdA3CjzJnkJvEX3d4TytP/AnBNj79QG+E3lCes2UF2pZhqISOBY2uufaQ44Iz0NeMSC9n
+tRGbjECz4+Qnwa3jPWzed02j/IF9RX7XCNKwHKcmJw/yHIa2jnhfXGycV+rW2BTSaOcvd71AX8c
xlCKhnyKdiYayGwfRy3hMXLuu2cdwaKnu/UJ1yLUb2SMopRlt3x1/DS/ujprioIUaznXnUPKvPI+
tY5o7OvS4nta5AxgAsVoz+HHq/K+cZ5D10lOXIDOatM1ESgBnEMFZa0ND/EVV3+YXn7orwuIkC9e
CVEV4WCQjR+/QOWg525B6zV97OAe2sVt80NsNA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3K+sUBRgBhLO7z4XKbbFj5Dm9dnCnLXJtz9DyutJQ/EYt7E+7VQGJ2l3bkkVJ8bn/YxKZD+Rqqzl
gzUxIUqSuvPPGmd3z16szdtLqj5YRAEZVXdNbeQ6P/rYfI4kn/0Qw+0hS8K2lRo5EQLrCely7fSf
ojGqs698Kv3dVxOM2uU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EHFOd5L9tY2zUSTwaEQFpNSik2aT5WpldK4px9GxR5cWZzjNzosBm4ckg29GsE3hW7YJVXJwn2ft
qvaRBZQhqD+DF8s0vynZ8IngOkOgp968BazD+XmnNms7D3n8pwwWq1DBwFf103zHNgk183z41Fww
ghnhfPrVLnkJtKMArkX+0VsxpoDgdODsv3fsT7CkMz19ja8WwHPQXCAKUD3p2rptjKIU1LKJfHEW
xgEccgVmdaHJ8o7kwvdgJQxZnf2Fl62jKVF8AJCrqXWKtvakZCxpEqbYNpoJ6R3Ns/YvtWdsZkRH
TW3+uPSDGYDVS3Az7zcuFIC462DOhpyBpwOGGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31872)
`protect data_block
panKA0bv3PlK6mDYG9B+EASQUJy/RS1iKZHJbzMofOlYe/PwPQbwSBNB2wMldslZpLUnOOqlp2Y8
YgCSMdHE0tqePoTJP9EE4AgPlpK9mQfoUPwFK896Wbdhg6MqBYzJErzTc0zqrqpeQuSn0mK+X1Pg
vJTYpugK944CAw6Xyx14DVSsiEvtW5WJsiH+CMY7uCvpb3ykG7TmqSNKXPadNcC74lKbh8RriVHG
y/vT6CgP4FHaba6qkL93yEnkq32nGBscMZNKDehNiO74dUDx12hCM4B16m8wzrm3NovncddQGLB9
Pm9y01JFWLSOMI6ZW7OOfuaAf2rwak/FT2CgJlyiaPzCraqRji8QTcuSL24RToYW+Ita1povpLV+
lPgWJgmyyJ8L9Hv8rFS6QrVrdHF24CsykQkDyTLjYwy6Gm6CxpD2lFObNWjGxYBcr1ArrZAqLQgY
tw5HvWQJ2cwCAFzdL9AUYEUVRlYqbkXnABbnCx0lyjXUKhSZPTvXv0QK//0uizsA0Pdb0rATgNsp
9gbIS9Vs+umqoOJAXsXhRLI1iHvOsZSjmBbXUgzOJ+/z1UkZNkMPtOIlY3GrDwTUapB4cBfU+4ef
r/qoDR9ecCRVVGc66Kc8jpjNfL98Jm0s2yw9ylzUqiB+N0lBAgcZjYNUJ2w3Y5+TpULH3V9/Mu1Z
wLkRKuIMoGAPnNFR5yidvCI0dMXORD/GONwwPl6yQF0LHFHdMJ4iPnJCExLFfms8E5dW0KN8PLcW
YrhtW/ljdLpLxORui7ZHJzDzAMUleXtCaFc5tdI7s+0AiVR929CUcrIVt9sZ7zEC9SpU3q2JbCGq
RxV1bUleTXMlk1eTgHdrfkk+WbOdxtT4rxJXXAuAFEKSPbH+xMh1ji+mBxDEYzvhlfzM89GioVEj
7WMP56JUdOLUcdfiUn7kESYY1VtP/U2EdMTW0Y5vzKES5ya8qwOPz2Kaiq3u+C0ypHlST8NqVgao
TQp/MchRpWl46nE8GTBTKLY8+kxVMFEiTqxbFKLToKtKYjQ3uu66e9c3A/ntrdiOfyjPnrRcEPdn
iZDvRtP2VNRfwP/BZkcxLp+pgJAS/2qoR+axDJ6e53dPPAuHAyL4PnmI5nwc0rGlZ1jLUTCN4vBO
2fzjYHUAPB73DLMjLk+iIwefO7bF1OA5uqj7Nou8aZO4INxXXwNnHcW95Raz0TlgwRtNzEvq+tbj
Rc3oYacWp4ukE4C1T3FCX8n3jXV6SArFsttQX+8HUA6EgBFxPSoIMNOuNOYGmDnJLaZF6JJSH1Bu
vScRwP6aBwlNSnipwQrOPzOqzhYt/Fef+GtSXD0dOtrHsdRGBgrg+Ot9O2OG3iX3xQOJMSMiLjld
sDneSvFFFczoHhpfaa6y67fePGy75p63eBOWviUx87CNU5Gxu36dLZ1/GCC60z5wWqGye1Wd1r5x
/KE4S0wytclD1Ty6R2mr519Bnlz9I9IkYwxYotlwXnmi/quWSsDotUsefgFhMhB1JBk24A8l/uan
5YfUL/KMmbRN1Qm0479O4H1OAsWG6eDXFO/BHNxrhf1nW6ZZqeqaRJSL1332Tun+3hjrMleV8UX2
HOe/IZZBjSpyD3Ac2vA3FkXXTQ3M7s+B0Cqyl+vQMWDjL8kaHnQT4jIUeyhH4yoIGcB18gqpp8u4
aPtTOFC53p9yu2bnC2H1DSSdAkVRS6939qFcmJiZPRKkeVlIWgy7NL17QvSdjYQeHS/MD8k2A61k
YPS1GyB9Np2PJuU1glSA//mQgs2k3IT4DKvcQF/ExOmeKuXsRdCp96J2inpMSJpxElh/qVi5mAfB
u0U/W9QRWxhn0vcaeRMIt9WvrkcUQJU9nXWC5QOjAhQSkXxKYoIMfctLY3kfTfLN1mEDo2PMIX52
q9VQfIAbv/VCYaaX7tMzwzaSYOvZwv+RsHW5Q1jvhCX9Mi46SP9/LOMUDsHFuwgUaHiFNN0IioiU
uwmSeXDHl8U3FDUvBkL6CUs6nRCnklqZWwv5H4v3kMsd+QOzXjBonV1xfVrhtut2OlbTofBimEmX
dGy3DSKzCeuBpfIJtTHb3pf0xdktXIxgH9uC6iECi/ImGTGRCYJb7NOgz3BrM41CKUFuqkmAtj1W
UWgBuITHfyeSt+m/4tVJc3ZFsTTvbahgMezqVsES3zRMImMPLwnzbTDgIe7xey3ye1tTLercFR+q
c6xoqVM6gnaEfDgAfooPOM7KWgUYSaYgajJYAI0yCjBitv5lvL3IKS6eeWdc1PGa8hAaEQftJLiS
CZ5WykWJ+hv0lRyK+AFOm0WoU2xPG//vJFZbRgHQKojg87P67nKMtZY99xTRzPfJUyh0lwQrAZ1t
9Yx6GqRJRqWo32dcxyUbzBQ+QiEB7hIEwYGBqDTN9LJ6+RXgydzemEd/PlhLiFTjca1IerauJ34q
GdnXwe9xjyRuiiswRhfXx52GGesKV87zVt79WKIQBPCKVEBOm9YUKNGTbb9sSrgQDZ02e+dL/cHn
HsPxXsfgQ7JYSiAwR6xBkJqNzwi1d61yV9sh3U2mdjqyMALOKuC930ShQqri3IBRHNleLCFKWjOE
D3VIsAx9hwGh67/Af3sIV0BLGRxSc/M2vmehM7Ac9t/+7SoS4bKemxVfTevQU6rVlJgbBh9WmIfy
QR/NffHSJ0cdYXzZMzu+XvTDUEmRaMxQUBQg7cutElGc+fgkMJ3VJJTOrCZBJvTxdL2F3JuCPtOR
SLHtavqBrKMS3eNps5Erk+qcxUCV9vgt3SKzKVKNzFCuaf8BXHPzWAHBpHUBjnc9QblxXcW5bKN9
MB1oMQkvxL+bo/b5Cx9eDUjyCc/Q0lv0Iq/CbPCPCZooSscvF/GqA6RIXn2UOu6I5e22C9JLcRkO
tX2Kps4uaijT4MQ1Gab0/awJL2taQUpNFOeTaTEHi+2mOcxfM5z/7uk7OYkc6CbkTkwHuSo0MUxc
Dwxy1hGkv9+6Yj0asfo9VNpZaxdoTECAb1YZ7U76+AsY6AeI02NS+IrX/xJJBLPFJCbrFYoYYA0U
YFjkJJiHYyBc8gFwlNZvDZFMSa64TfgG7HbrJm195RhXu72tKK+Vl+ohq6F3ITDL2hzQuiVrxb1s
tca+EMESHYj7dlxgZl9vp0fLW2t/DQQKg3ZxsjtpSJpfqfiRu49adcvpuoFfdiNngZuw2eYMTpja
Hqt4il+nopBTq+GBiwwK/KOvlUE6UUpd95R4A6BtmLHqma+SzBNypTi6XQ89l9f8/08F03dFLjuB
xkUSfo+QIVoKu/3CqRwBfp02Og3k81Pg7HzV7UyhT4eR1iTUvC2LI5QZusoNs0Pg+whTZG0oTJVh
wLDyAef5ePf9fq5KtKGeD0SNSd/dE4KSONb3SN7VlLVs2ESu9RIperDYsvB19JfPeXwQlv8v7V5G
rbM8NeLMvbW9HBO66EbxGXtHQTP7xCeQyf8BDRzNEO+bPGozfYuphQt0GbbjT/Y8U5YS1yTPO/aX
q6sxYUskBn9V8x6NTfqzZodGVT5Mz/VwlLhsVWriqjUWHUQjcnptfeVU/bi293VI0t/NW+jynyx7
gRThdttjGwMmTndcTTwvYnSlJtaspYXQiiTvZPzLkh7PVP+js3FGXwyK7WIgr880Q3rFSkHaf5I5
5EtWKSRlLMkgtT4Sx7uAVICjP6m9TB3nghkKRRDZ+12yd2YWtDHnJwXyJsi0puGg2cItUQLXsiVg
IcXKSEf3VRXfit0U8Gn01smulM4XlH53MwbjCVirBN1GEgBGr4+lEY8cE0sPhputUfeAjBJzhcgP
9vUrU3unzGYi33IOxAh2qHvX5bU+mP8AfvIZmZ+d/3LyAPNV+8fjup0F5BJ0mtdF/rILP6m2XAz1
7EunKrcaP/xLq/WDjyyG9DLBHhaescplbfVkgFSc6+s/CWZdTUSTX8oI4d3v09jTTkdU7id3D8ZW
5xtP1Yh64IAzOpwYPNpddpymBAA1oG+DMzlDkNDEdZUPMbFooS7TM+cgxwOoyecvlBlDenADusWs
WpLaQoVEeLLNcs14qQ6nxF29HYkIZGqslNFBcjRKeoD+X/5Y5czeFWcwjzRrpuBNo9RT3xb5YRJG
85Tu6JURudfdxetIC2bjb9HPwI5h+DBIVpjoFgSJjLsRhVeni6r/jkk6uGlRWaVx9TlcpvCcotxq
2UmrilMzYUue6mHz1M1APqpngFYCHNBzAttrQmqlgSiJNAD2Srf3EOb+HHLE7U/LwAGJp1mOsLrO
cqL2IrsWAEcsV+7Izg5braIXyHX11KgfYGVcbPI4mAGxr5pThhoIDKSxMjl6gCzjbIVXpabVvQNs
P3aq8OjaWyecaTKlEgB7dMWjrZWxNIE9SeVTCSXsnPw7uCLOvCjmVJuR/f5yLY9xhwkDYX/VGR1L
bFYGXXnmc0DoliaDLs380pOOhcwseoNkbLZ12phZIJiC/5deuGzCdVEuFsody+PlPjOI2ua+EQzB
Pq7hGvd6bnqmn5jWvbzK7Lg4NIwdL5FDMygcDv/uWnJTGQ0rp8EIG90WHVs8L56En5evBGHCXtz5
utf0dyIH6AOU0PL4D115vk0JOCvfwzxnx5OM6/FVEIRO7iyct6GEHwqLM4P8XjWN3M96P1KGLfy+
BmbMu1NQd+sjiDwHOyLfZm5bPrLEoTT41Iz4zYuhgKnUfPGNXTi0RlDR5xa3/v32h3mICpnjxJ0M
HV+X4oZhP9EZI7RJNN+rGdKwnPTTmVYhZjEcCZhzqGDa7IlMKGtSMQVZ9cAYpe7Gvt4jaTIgf1gv
D62KlSMuJNzgHyjbad1AzpDvi7w6dM+TvwyNqm3ahlxGGKaWhNAVcpvZ6zj2PLwTRVsfYc4hcXQd
Ech1TC7rfPiM9GPmZt6vkaX6Vqe//gh4L+UOKG4ZrFZcWszPzegQIa6eD2GusHhTEzWAn7f/KoaF
5UBMCsHYtvstn/jvz+c5f6uUQpsL0D9O4E/YTNvrUrZOZ+Gpn544FfpvV8a29PGQh2CEa5b9Y07e
e3dkiNaZIbNf8HTZv5D+uYgxDZH0eJxIoyGoCEPlwR1PAZQLf35qpRxDZWlDXRlfoYyLozIwvGtK
Kxa+mVceBZ3Vl7Atsgdx6TVTojPjKonBFy8qHgLdNQbCdNnGf2y/vIyiq+q2CFz6XdFseYZTA3Xd
fvgJiy/DXRSprIIm5nAiJMq3oMvQDXTH6g9VKVlGGDtbvhP7EGyvc8c+o2UKOZSRtDhBi06M4MIQ
Q7KrczdWKAGif0HZfDR6DjF0aTAByGmxFh+J2LGaWQ0JatCZyDqTKYWQvDi7Wei/IprOb5EIJPOf
asUuGLZNnxNrD+eZx5yqbxCkefoSWZzpE6hDGh4w3tizl/NHXd3DTVvpfUkHtaik0ACjE+bpxFQd
ZxEiXNmUGdy2YgAtbNsgmS0Q4aiyzUdK6A4mF/fodE41yI56bO50YMduMbV22cJUAXeDOy/0sBMp
6HgQHFcjsiLrZnAI+F1LYkwBPz9eAig2JousvgCeRwOZdtsye28uNSndU+x12Gd5v/j/8gzp+9fu
csXvDMl/CpWCJ2MoxYKgX/t7aHhqNOTzf4cGmYkaLjvmikj+Iz22is557nPmgEqgCMGobSpZWAFP
THN2GPMGROuPxFRQtwJEc/Aj73Bfsr/AtuzAwk3URXqLHcLVmFkAVhp7ROw/qjxR3/WvE/ccusCF
aatdjiuYeyYbQ9P654tLqchl8yZPsaiIg55Nyk88U5B8cxLO8FZXVslmAR7uJM8vKo7gpPFR9qbM
ioi2gWYHswVpK0KdKChUC11Dn9x6GxoAm+UYENR5V4NPA8pVYCcCkCy6qNYMs7B2KePtrF4Tqqij
Laqza/6DoJQ9RdEInXgN16G/lLV8QaSo+9Mk0E8EzKssboR+muhMM1rcl2RQIyv7QuMtOc+ErfbC
EHTo2+4jnnvsuR9lT/DzBFJDyxeXUaL6RsvvuyLwVh0/pjuNqyqwbQf5TiVzPKdXhUlTASYOYHhj
9dlqphqpukv+jQFdJb6ZcLRTorblvx4EDQ5Ysq46LrdPYDmVeMHt4etijsYnKYbj82lOUMZ7I5dj
S34uKwfsLEpfg9Rwiky/YX0x0WAOmUeeBRfUYVXCUfIdxz9ezf/KClech3Q52Md2wFngLwXBHvId
nhgEMg/uuFWIG3O6g0eMUzj1N07OXYNcb8HFyc4MbPa+UtVrjOn+23JU5ee8sNmVfCq8kkdnBM+C
/EZAyAokrEeH9i5yTL3reIWCngQW4JN+bhJgybuYZN2DM0xU0cQJSqYesFVyjTCqebHwuP8ojDn2
nzicQ0kJZ2Z/5ZQ6aJcFQ15lXVYtMrC2Fr7/akaaedoiSzKLxe9j1obn4PW3Z86CyN7KzbL4ZP0T
aadSjYRU0P9FXYGHtnv2aRdSnLiLcQus0LJm9eBMDvd4lc7l87FKZvXBMX2tHOHUq7r3c28w5yQS
aRQbzNToK/mL6Usr8ntf+NizlXpCd++Lrm562Ra1mtcd8peK4ZM0N2Lqs68iEyCRQJLoWETsfn+q
17nV7MXqS+S6XiO/oieEjPeBTl3va+2kInOtAt1nD26A71Am4asRK/uKairINfzVQk4FKAf+sdDx
jkRKJCRe57BW8Oh0byDKNuc5TcAAeAZrGA8I/OStTdUeU3knqAamjaPsjAQoj3DtLzF2zoGKt1A/
+UX1kj3QCOfFS2V/AyeDXVN5lMzJcugdB2w3G/Uy4jchr8zIg46EBrhdnjqHpm+qXBfCKn0TCQ0x
ud7jOoB4G2J07CWP0o/uW82bFaBLAWtDx5TzbAsV7uyJ2C9KRpIuiYRN1/p0p58G4DnrfMtTDqlL
k/IXpkB+kjUfgoKJLaMMvlNT4e107y56OUpX5j5Yg2fqm62QKvc6Q+eTW7WGSWrcv5qmLwHLOM8W
3k7XVOg681FXEPy0USRP3n1vAfdZ1ftCqAplqb14Csmjviqn1ZGkwwXQyQ55zAPPaj/A5eFP3mlJ
9D4orMp3yiNO5N+0CkrQIGKo/nOFeiLBTqoIuSLiDWigFHOTOaEr4XfHImbLrTHF75NFxerwCELg
ztNeJ+KPiHdQJ8XdMtxYDIsgs1YLLKa0AnxWwhlnQGE1q863kxNzqtTXo29DDgpt5c5nTHgxMojM
DYUEMbPTrAwk231jEYk+lrq+ZmKAHhUVYZT4JhffyO5LaJVo/EiIi9a/uDmV6ZmzXv7tma/vz6GN
nhvShUcPg1FE7xL4z91HJEt9rDHPy5OowN50aXWu60a3zJkIAEHUWbo9Flk/TMe59oL1cEzzcBox
/0Uq6IKhIUfXlnegXJoHyop/JEKVjF40KQXRDCoHOiv9KiJ28zKx+CDWxp8kOjHNyEY6uCWAcVI0
eCrW+O7LrzubbrOCFFIeCNknsg6CQ9VzYqtksb5CzymHlutOMbXNSxSJ/BqZMMRx5+p5TAo0DBJr
8iwqEi6V0tZ8DHdapoSA1ms28lFl3FfQTNAMu2Wp54NdUSgJIbxeq/3NTsFPMiCf9j0mG1Rqe2T7
asxmBbrFiQ9LYO+CR85murN6oNuNEgOX92hjZHYHfLtHx7QyshLha2iz1ICmU3Zb5m9NEMOnxjzn
gnrFMa4U0pOgUGb373j9I4EZdppmB7NSSAP6spzj996lbx3vtB3LxrbnLimYC2pHUbc0vu9WVM3p
RYfEuyYMarVLKiltFpk38ks2t4JlgsvRo+iz4OaoPln3zu2G7orwodjmu3wf3fQCNmAfQffLfqbA
f1k7qqWNefv0yFsNbLkoxIM9k4mBnu8EKLsl2/NGq8u259nuCLaDU7soO52lvbeZosKoGYpbX+2E
MoaW/2/EatCkrJSUHgIGfnEbq5yR7Xvf22/ZT8l2n9EUE2HEpbwLx4eTKRaKD6UEd4M04T5wFsNX
+24k9v7rWCA/o0T1sLB8w3nByJGbr6dPXpMQLhOotn4fwRVwBghlbB9M6XZa1MXz1QWuR9Td8iFI
hB0iWi1HCnALlMOU7Mznekf7RWDotctxPmNRq6z3kkWpkeR1h/Qofj10By4sDISmZrAyHaNIh0EE
bQAmeErVQ+loUNTDMH2KZjfKvfw9E8NKqS0eEyvbX7+kz7Fe30qsBtkm1nzXarriPGUGcBDls9Zo
WhxEBM7K/iLvKrtPIw7ZcRZkNYe/1E0sO9/Z0pvzXso1WYkrI9p1BuShn1isPr/YY0CIY5BKDZo5
bNjxRpxivtKwt2wd6fuicg9psN9K7c9iOHzuMjUalBaIcKGIpVjhyErZ/QYvmMPip56ffZtRLSwV
DjwlM6wSJ0dkx2HPBhj9dXtLGYidk266CigOJ8khfH9WKt06V1InSsklj1IGuEyn0BTAJSodJttU
MDx45CLMFS/YiKDI33ifVNqi5X5jcz9PYvksS5ryWERppre74wUDzEy0LAEovvKf1ugK6VO+z4NY
o9VjxOXL8WBNexUcHwYpDGJazufq6ogkVPCNPXuW/v/d1Ay914H6nwU33gNC25Bh1DNMajLINMfu
Bo1Nuxqrc32p8D350jcTr+R8FwBNHswcJn7n5gZnL8jsGegRDsQF7hsVzDiH9i2eLr8bNj6Xz/Wu
+xNGiymHeLTyU+fInvlFFVNAKvGNOkOMcX4d1+Z6bGe8IwPWhjZNLmJPok93f/G08r93DkRCFZZa
4Ty6riSkGosu7KxcVftJE2qFA6+ABFxfu/e3TJMLAuYUihaCC03S7LN/ChGBKk5y1M+F5XgS/BKO
mFP3bmR2WiE4v3ps9+EXugWpogt9boo/aLj0kKzazCVw4AN9qcXwV/DdJeSiM/Wyils2MW8BlHZm
xIa48irAj2K1NocwZhqKo7UPg/zssMbgt6ebiwNuUCpldK0kZsZ77t9VTrOQoQjay+AwMMO2WAiG
8i/Shu/FkQbCCyns2xgDKyqL1Y7r1v195QRJ+IBZxSXaERlnmiKSsJYeVlCr+9MGKfuUPuKSy+u+
aHAS3XTP1rzCRqBPDrLwMk8t8Zy+jF7I1KEcs9HK3OCDlEaFnuk6Jo3R+vbPKmIx36j5+HaTPt6K
iwSZfNESFVEbm4PFjR/CAwCv999zkwsFf6XSvYldysNIz0HPPz8zqjAj6t52Kso9UCUnR+G21GMQ
dcy1gGdFbrQA1FE8yhN15YDBEctU27bIQCJPAQ1JkHSoIebXqE6DMRwTGB9ac+cjmgY90DkWZWCB
VusA30hIYb7kGJbyZKZqD5qWjk67DqOC35QtIsPWeuYmjpHe+zMFiEGjhd2SXuI2BB7jc0u+8MTD
TVFf53Pk/P8xNs34Yy+S34kDGqCpn0uyfNi/3e7blnqlTiRgj/sCHxbPyUO+agGUtMih2ZMry0V1
TTzJX3Ff+H357hxVlrs6sZaWY0Z6f1kYaxhSzrB0IP0FeUn+oII2ymUel+ON7/Jdt5LfwScY/EV8
k9A4Br+l85+h8K2M1Bg/TbY3Gm7Hum3dJJa4nbI07HlBH2jqXDUNUVOmzyGk8w4FTRFdqG2LNaJe
D1iFY6cKypdrNRdsZsYXAkTGmHvtLq+pyXFb/HCMQQVJ1PKXlXkJRXb1AJMXbZd9VD6wF1lGhvuS
6y4ncrlLWz9Ku5Kxd2TrFIqWHhFvVGPiWVUcZ48C/T4Ldezimr3S1WyVW0YaLapoA1AL4KyAEFB7
4m1wDczG7lQR1K5LEUF1AqhOf2yu9U7z0U+sOYRgVtHKnArkXjqr9TNgWfThbAk0epxdzxGhh4Kk
Wa2aVS/3ac7GQb6doQrKZ67Gir430BrF0uoCdOxSqmEcDxPCLMMrmlnBY201aUaxD7bCAfv9gcet
LhpmWeS2BiyozgPRJNuSq6JBHcE7qmKh/amgw+5lXD6K4izgaCSlp+pm3V/KQbAvbGbbewfZc/4M
+hu8Kl1XCwtKFEk8wsAAxlDmso0eh/XlTOJ4uU/TkLdAkZjlOz5LD4pNHLJvz8jjaSmYDpSXfvpn
ourR8TLaWePxA1Mkg4aun16Zr60Hm67LBExDC/7R4jQp3rPyUH226hysMUMmmncf7YX4ZHB//Mwq
HVO+MyQJT3WeOymi6vQaQFwgQQF3LqUWBkL4NHIf8iO0+2e+jz5/UA3NaNa/0L+vP56vYwx4NpNl
Cfx0a3O9MCpooNe8lyBJI5V06COJSnD9rYi5ScUBqKSb7q4EkgwCc3Jo2ezNdZyYLPD3xf6JxNN9
qnaXGD+p6jw5c1n5rx8giRR2G1MHeQcc3EDG89zeBompP1u29MkSqHDXscFdFPqEANI/nqX740Hl
DCk7FoV7AxtOyYip0kzgLf+1M+l6LvCKwNJW4T+cLCs32EeT7yCzhfoMIVMPuQwtjX7ptBkdtJJv
PJKHvs0Xrh1Wx1jThIu6MxtElSctp3WgDIIHLYy2HxxjcjZPc4WANp71v2XA1L7tIAlxFn8Qg7ks
/ZUHHs3TeLk9HDqev2wFNeYmKTqTnzTezVsK+OGKunszBKB29SCv22YiaIwSmy5pXB7hZj+SA0/E
yIXCk++wY2kiUN6HlGiFI7wiJFr/kkUhUzhPPEArMn+uIEQr7vppPLt6rp7KPYme84ht4h6AEPsq
6/opZcOgtOKFFVNcRjgddN9ESQ5VSSWespo90bYmHnnb0yvG9em/hXtH3Bdzej59p7nCKmM/8Uu9
kTp3c/PYcsvKpj/CwdrLjJhn01d1WhSayA/1YDGcOoY6/FGvx7jOFm9RBNQ5CPa+gSK8K4gzRdmJ
jWuMGcRayyrdpfuOnkJ79YhZOPGXb+fJp6dVmiQht8nBmRd7zYpCU5T5zaqcf2FyTXV13Tb6SBsu
4sQISvqFJsDoI8vq+FWESSIyGkTVJLQ4caKIoVuJ40WNCDq/za6E0RWoFwjWQ4ZC0wHJ+qCdKqIQ
T2QkcVbM2Qg5VSKr+CoJXnB30EtZt+ZATK2j5oZbQ9BuaE956AQijHVWiNDGEUQUz5t2v9A0l0Wf
Uwnn4KE8rWVtqmAJAgIHj9Jjw4AfPphSkBMZ03GOml7nkgGGgylGZhDWPVVCqD7L0zWmCXZTkLsq
NVTffRsLU2F7yfPjSOIzZbR3+0bVOgq6Cob3hg86LPKvVCHjO0s0bCVoGAVp15qt/9sQ/3moWuIy
iwEpp0lOByJkymlxPcV9pV9jicJ+jSMwdV5pg8DfVJpTvar1XC40jx8p8kMDXPBEQHqqW8zxXMHO
aoMIQCkykrRkDAqunt+gycqcMBgi6W5rwa8TgpCdmuKk7dU+TSXpO15/IiNNiYbLRuO5vE0iam5p
z9AoI+hgaHLbx3mcbbmJ/cMifAkjNuYFzyjH+hXhnJNY7fCEuH7sIk8+dsboG7471xWXsxDzjVzm
7bFqUlQu5FVtfuaoSZDeql5MD9OHwl6KnM4QYUIRwA22+LQdSnk/oCC5MAUutbRuLB0bC2S5cw8O
NgqsTYgPRsg8nBniM8PUYwe3Ij/iwoCO5U2rvjzqgilxBm2xUAWXsOJbn+KJQ6u8kuQ8U1RAIbxQ
C5GZ5A0IG7VropVWLbLqKXAYGuc0aP3wmvr4OkI1+EsTsXMEY06Br1i2l8dl3p+9E+qUeiA1O66+
CEGEVxppY2wpe+yesV1uzOYTfOM6sCa5lo1oYZygpBgu1XReoEKOCjnBosTqipFggw5hY6cc4Pqq
H+Di9IGzwoAUZJsOOjt5Tl1dRKxz8DHMUdfMSScDsz5pcU6NzFm0a21D1E4YealRLt/sDa6fNRZZ
6FAd2iUDCiqLt3x0QW86LyQo3twOziqOcvfQgabBLTJkt5+4Ea6snMUmK7mi+fWGvR0NrqTq+vwK
sbdBLhqwTdrc8anMqXohf+YFmHpxoJrIBY3t/RBH/0aJRH0pr1hmAKNbHMP0McNf9ee8O9WqzOsq
Su/FBr0S0sfG7kaKsD1WIQ3MZIvDU9UZBRkylIGAO+Hseumbgx90DoEmvAzsKL3SuLGpEE+UJE0P
d2C26sBWBposv8j53aM+006vEaX279YMZ/c7jWMX02GUZF6OxuMBiAw7AUPgTiz0v+mlDa8wf8UA
7e32tPhMsSJnkBcft8kRufMk2sFcm5e8lYPZLZd4WI5MJeHZwB3pTgVjHv+3Kq/B5gEfObOqxQur
RIEandpmRjgZ0cLCdY0y9xHjujL1S66+uWkMB6VAQUw/EAHKCqBG1O5iFhMyUL7pkYBj4RBMCa0d
qzTSzlE5h2OUVLEPwBi7JYlA0F2KNm1NYXuABXWqv7UtLvfBmefzHr6VOlX9fZdqIjbuc6yuuB6z
pFyMfuHZHXvwXLiQjeMu9DoZx5AZs+LAML4Dv6D6p776ixMaD7Y5x4wrjIGTNb9L37/cUIlk9HHl
qcWgxpUGb7VzsGqHJTZakMHsUY9r/Q+GerJ+WtuhUaUrUvHRnvXlKGwPkuMIE7qbn3de48kSs9WD
0YzN9QGzCodlnJrOKudszFDxyoEODTPgQgMO/IpMUQMHZosG6W1PipcW0EWekxG623Q+Ti1CSOFy
rwYiqruqa2KzoISGzAcD0q2vYlYyyTF9vbrFa32p95jjwIVGkEgo/3YKNkRcOmcP12SvQIvYIunq
pkZpWerqFGu63R1amFw1bVIUdfLM4bf1c2T6WB/UvKMlBiV2FQQqUKSCuOa0k3z6QkJ7xJ9aCKuo
tHTC0rDWefKUp9n899lhoiVZfnmg6VkqDloCv72gLxjh/6J9m3a5XwoqWPIhPAoahEx+c5I8ORFw
lZd5/R2uP/EaYwGl/7qY8MA+3FuSB7YzZAieMoB1AmbFg/BYEUOdpHmS1eYNyRwlR45mQoSuBx6f
XQi1I/B2dF1btrBeO+hfF3xLP18TH60cOeCPuI9lSFWHNYw5zT7M3w+bKe/PikE4nrd/b8M2F4D+
B+bZk15Ulo4k9DM8KBhBglz8QvSNQ2cARvTQpOyyyBzJhjOdMb6SX/Ct50r/b6XHZrvEuHoz2hPW
vUUPTAcrBbcX6rWdVDXHEMM6GZH9VOR2w4ReSLQ717On9S936XmVwyjyZGrCZOJw2K/baF16JNi8
yQL2YIxWZ/3ggjsabXFE0f2eAeiBJDDjXnsHBwvJsSxlIVs5uqvF7rUy6gywjw4U1mdF224xm3AC
dag8fccGzs9VmBYYzspnfUM/fq/ftJzsPV4tC4uq26mL1l62Bbc1HJUXy0JwzmU3KVNMx4TkHUHK
XgO3Xp6dzhZdmB0OOIVEUtaIrLUsGyxo4fzurcbNYtD1sjlMfzgwLw7kNIH9a5oGz87wc8+9vGF5
7QTPnCF+SXaC8MoUOo8ke45BR0U+5oaeX/d377KQTWM/4xmtK76RUJKYs/d9E+ion4q2y1t7Elcj
T3UfFr5eaD/dcm2WS5t0M6b2rRDwct6qHKst9LO2zG3SHXRJydzhlD+XfgkQpf1PfGSkhSCEwxiA
uj3nTWjN9OQxUGN510/AL4Qcq3dmpzRw0266HwQ2lBkOBoxfkXBDf3T0hpsYaQO3Gi8tE5xJXU88
rEvvTi9k2tsaj4Ynfc65KngepYOrovjm/PP6wE8F2oafIhgZPA40gc1JBiUETt8PqKxo0PxbOyf5
FPz/98PowZ9LJGMIoSD7N/or14i9/9NSaHKK0LWVANP2JVIT7gym2zmG1+LvF7beCqmKzM3fAsLH
o9FgIpCJYEFHnzXf7RnoYrQjJmREKI1277Tx3r13iLIimSnVHZyRmbNj8Qdq7oUbgvjzssG7NyXk
oi5600LYNCPe7bpysJcv/RS8Hpu7BDLNMUK2Gf8W0BvATA9yImFMJNBATxzdDeALOzlyiIh+UII3
8pUDU+wmdlIqOkYZaxrp8gnLmBwtcgGl7CsnPPtmV6yyj2xKBcci2RvUA9/hNVFNovGOvVnKqjt3
CV/4i/q1WcNroEK7pVXSJCyLoEmZ4Ztthw1fdWhw0TlthREUuUF2FDqB0NgT3mpg4Ssb9G633O39
B6Cas961LlB/W1bI3w+hc00kFRNemGcvwwQKvD0x6kincFrT8CJKCVL/+hJ5oCSIdTBwaPgZf+K2
MEqeJcZAI4gSGrSx3/2PWSIhk5wgccDnORaqXFF1tdOE1BuIwzikBEbgsTJnyRGia4c+KrgzYr4K
j/QAjDCwrYFMyCIek8+4yBrAs7DllkiumzVCozBzvjrQNIfoEGIUskLjeyaSFnMuArI0QS/7Un22
+jtESysIlgPw14MJt3J+gKgvR3dn4ooHg5NPG4KZVxpqexGz25NN1+yuVP+5tc+FuTtbVN5O/MZm
Pmw0fMqluHAcqyjwNtD1MWmJhV8RncU+aeBYLQFlGBFjp/RI55p1yuKblBntUelsQq6ckbgiEqYr
giX23ChAgEHuD17Qst3mtpwQ6ZVngMcdosZ5tGNiJHvT385os4q4EDzMaQblnmp6J0n11l8fXtyX
avcsmgEnZCyVC1JsI0CHL/sOrO0q4MpL9E3snTzYbidmRcfUowdZRJRDANN4a6a4BCuk93KtjCKD
/E/vXjaegLuAOK3XzDnJxB/PZagoogrYLsRz+ducMdqOR9d77IB9mmnHpPkT9K+xdSIRwJQ9taqV
gnViqfYgIEOEGjbPeUQ1/Pn0Gl1do9SsxMduE+BnNRMy+g/2lifYafHYjMk06EJQdZpyen4AKyR1
SiOALoYi1SU82hImODDk7uxtO7dSVs0qGgYoVAZ5ClOkbYado4SdLepgjcjHCZ5yZLy2SfxKyN3d
ri3rKOd43JYOINExCt9cP3YqlAqLMrkRUXhwpbQqz0+yzKUeBr6QRug18yonJke2rQAqHvnzKFC6
fe/7Xo2V8Hcs/lli7tP0P0xrJmRXZXDJW/2rktZqrfDlB1sOVaMjB32QkMYPO0W60qelkoJUBwSl
7FCD6TY4nG6XaVWtOHr+e71KACwZgR4eqIIQ34aDs52CNOjSw6CyNjWktMD7iVQBxOXU2LKCWAEe
0nY2wMs9HXJOxOJ6v/+gZja//KtwCu5g2cT3G3+sEeNpmqTvQ7LsQg5KgaCmiiD9KPwUO6g1ebkB
Fc8k3z/ge1MJ0HacMhmEqgiGZpiEExxqGX1jV0Zr+jne+TSs0IAuhYLk3Wutf70UN72/XKjqBBOb
AyehjfUk304tJkbxVSRQNL+u1/ufVuz40Brxiw1jJXBaUFcDvwUwUF87aNUW1hN8FNcP13uMt5gL
0AjfyGaU8xQ/elFP0QRACAeJxQt+TaxM76xqp8PTKA+hnhpvJkuBuLUOCg/6r3jJYJB8QkWrmu7s
0pN/w4AcVBtIJS+O4MytPHusjOXCcJXRaCIlfuuZM8L+0jNsrBh77Cv/zLaIDPxTNwuCjpwEGyP5
qa100mfuc7JOWbrfwJ3rwjDR/cONkzxNY2fcjQqHaEAU68wZzWPmxRkGUPM49j6Oy+Xiyy3KRDXI
fSIJwEEMXnVwHfxUiyFFMNxgWZMLSWGeoPzPNNekp8655rUcQEC0U5EhjyBwYTR79nYhsyEIURak
oHO4ra+iPZC9Sa0pqs9upAxlxBk0Rsn+bT6+aR5SHGt/QYj26rCRSR6omQNnxPKUfyZLxVvXzESk
KhzGQfLwF+K7ZSJcrihV0W4P/iPVHIxM1nnMa8SIKZHlmVRwiJ59VzH+/u1vnaUxq83LzVcRvHpr
sirVtQ5nG9hNLPD62uUBQStEgfsfKd5jbSv1T86zBjAfcCtWQ9W3PIGx0IacAxoWTqlEGqSWnba/
WV6odk8d9N9YNojmPFRkD5WP6xp/LmGgqDRnxbWvnSY/7kMIoOzhRAU98kZLC0GJ8ZuEJHFAVriu
cjfi3i0y9Asqe7RcTCtq5vY4VsBnd2xit5sfV3RdUprnvKx9Lr4QZjlJnIfk1CGQ9b2whpL33yyW
QcwT4hhDkt1gRPYmgZljUXI77y4TIi61zFx9aDeypMIbujEbAHXDg1pCOfXP4p32ncmA5mEtkawp
6qtDs2vNoug7OpRMKhi4lrB1eBJa2pkh5Pt22fnhvjFBkswo/swjNRRiGnycqTImdDJZhKwnxpDy
1Fk4kResv+BDk0TKpXuMr+5ox3cw0ewlQJ0Qvb6BpiUNFg2jvyEjtdYk8nGijR5RdDC+EkfR3w+h
0EuoTYv5T7t2J4lpAhoWWRIVadNfAghXIeL19VbeyMk3qTtgSkZJ+p/Zgh3omN8CdPWVWli/Dna6
uh29Cr6/zMJaaUohheQDZHZBgTNIN+nqIvewuPQbHb1uAngXGr5ukvf/UpflmcrAD3Qt0poZcI05
X5I5GMXjCSvJOZBk3UKe7Ld1VcnC+z8B9WdravO+F/lgw5dGxkq+8FTDiuTGr0j9u8AM8NJoKlm5
Ua3tawLblEasuOLnHmvEvDj3RtgsofLHLzlPv40HTHYAMljgrGMxtcZ/mrFGC33ZjLr7FWOjeahq
9td4+T0kpuBnOrN3mol4jywSwtaVvxCFRrxPFf8F05M/JuHPRXy+CmRaEVmmaIF0YAn06dgtSr3s
lTenGs/GdN9SHL8bY3tiwV5pFmn+izv/2j93TLtREOk4b9MlJDk5N4dgnGMVOf3wVtlTptuynAq/
qjV82vP7ga1xA6tb/pzYOK7zq7E2TfEhvVMbaVqH6y8QHQ4x3ggN2YpvQ2BaWlajqbYctk+R66M4
x3utL+LdPeNzrg4LRzhwtOCY3TxDllbIQMBDdodU0ixst2OrH9EFFniKgwAnI3BMlEKif4cFnZHv
PjKZZAOq+M4OlQrZ2zeJpjJ3TgfKP3xXbjFfP1hEhAL2rOiXwFKYK0BoV3Oje3+e/MrEiVZE6lX2
pSumSA49cimEev3PinnqaWOvaXhb8FGsq9lf9CHIFYjkOmJ2ygiaYSaG99XVly3MDHa/JkgjGgW0
6plw/rsZeY/rhHFIsTjWkXjm3ZL9KmzX/eJQUdJ1P47iP0e5Qfo6uDacmKlEGGLvWH6slpwB7BaH
OYYjhefTemwHVXEus3GOc1T23LouPKKIGSvnTzGJI1uQVq45/HzJxdRxAZ1wAhT0SfAHpDGiN8uI
7Z1ur/o1ttGaU8ylD2W7nOR1VXLgKYYHl9NvALXec27VmA2c3K70SSBYSpERYP5fM3RxTq95AS9S
rGhNFPXupyW/LJ/Rm3afG3+Itk7gUORiIUHctYlqjs5xPIYZ4/OelYidnIe67EJ5wPbbRkVqtCxa
Mgir6CCPLd2cANyvPuAE2BtmIJAF/5ee1OaGMKCbqaRhVrQZM3kNsoio2/m5OJkLyOVzPoKlIWIv
sHTvNuSHe+oSm/X+y3QzP+9fNXcw33srzvDtgXJlQ2UAAdNJrlSzSmDJeJ0+GUAGhmBhSl0ptGQj
bWEfVsyfv+ABMfIzU5ICPkTwXTekiSXSaPqoN/cbBFKUbqf9Zxmp17kBDjDBOIe+EtrqylXTZWYI
DHHbLW/eI7Jj/JBbQ4vmG53uKlfoMzbp6FPz4liBwPmCdVu0R1swF0KxIOh9c5FSSQuFsfBevJNa
dJjth0zzi1rdZtqLdkMk6Jc2oqzYVvbrVRsMXtj4C+S7NR8Rz2c0y9r3mw9XQx7I7JtVyRiX2MbJ
5lPr9Rhf3ZrhEj4kd46RXAT8eArhe7eXL4d7d7UxdN1kcUCHub/Ttgc7jq6PAOmmxaDH/k2Vvb+h
cnHwdUlzeu+yppWf6dQmd0+InIeoVnzKaDPSRwuV8+9EV6kw9kg/kZFp5TlvipEJuN/+rIP/uOll
/sHkJulaJ3SA/tFPsGXlQ0CxQK6RccljiYkiLzA1qiCeJ2jT0izJi1AAUAdQaoJ8S/TxcfomolE8
oozCKb5F0FOOZigWIqbewwpAZHaii+Ie+k9M3qnSwnoriPWKFs6JVzQDH9Dul5qrxUWcMt0kVI2z
EU4jpZjOJGnhPBCdLk4hS1wgqhzokxjFboQpNlMmaS0PDR/bR01GWHSRId+BqLMjKNYiNwPeg5Aq
3K849wHNv8Y3u732QHEXSKpknml1B2pNapqt2dPH9B8IXtSKwXgOfONL6REbHHaDLXfzgq5/9hmJ
F8C6ZBQUro2T/qIkNqbufJHw9ebPyslXfp2hF5rWlJZTe0PoBBAjZ1cpWyzNAwKmLJRyusx7bgLW
kNEio0UVO9+B6w0d/E6xl0HU5EHoZo19Uy2d9/MIKyb2N0EYtyXTWG+MWnNNR8ERsPLD7xKpC1A3
5Idkvq3//q4J51fEGa7aqN7FUM2tZlmTS82erFPt+HsxE4JvEIEL0yD+/g7muwhKkAFpfM2iGazs
tikDXgwuIVrxvIwaOIb9o2O9o1wkthE5TGe4Z8Osm1C/xbXhc5BR6iqWUj/63PINsPvPFE92/tAe
neApcS4G0ZyAo5Oyfv8cR882IpLN7OZvq9OmwX59eXhDMwtazde64zxJb/CkQnX6aayZqJruFuCn
6v8JUOnIbHtqrbuoaOoYV8rj+Xhu/p1tN29z1FW5hKIWjmQksIwDra12QM3c4i5zRmdJMM5o/eFj
z0nfoDMS0fUKcJPee+nuqnGJOZjXJG0TGe3pCQxj5SA9vf4KhOw3F/RYO9xAK0W/MfkJdgEszyD6
8F5RTdh42yc9JjeI2qTSDO4fHr9aI3iey05rDlfTul3tVAvGebi1c/BMTd4909bHGX72NazYUU80
Tt1by+dMqKzP8hZaazdAylZUJR+4nJSnWTk9C6y/xRUaDUDc9StU+D2bo6M5cjJMKsNjnJOW0c6M
WQBqX8LgMgitsBC3L0fjYWcVOrAx8BzSxwtLXEcRU1bygVjYM/yQhrBrVIKRdJruUQgSwPz46USl
ShX5MRQZA2LD6o2Zsywa35JYx7JIyAanVpHYiaoMd6shPPoIZL6b5fMK2O76eIIjMaNsWqdAZ6hk
Su9v8//UWIhxYpFJ2Q7ujblKixnBHCLWi+5G+nWhD99UcAAh/A6qzGkj392yX4RL4r94xg+8xcUC
jyWsR4IFOJPnaH5rCejDWAEWg5KVqZTDaLxhXhPLaCG9sohFaE6Eexip7J20Tq9Ws+o6O4hJALI1
GTIx7YwixCQFSQTLkDvM2dI3Z63KQQs9e7nSPCfsZdU6+mtA9NcIO/OyRFLey9Knk7bQF2qt6mnG
iJg4WNaC9huDNWyJR98bh7v0t8LllPvuaH/NO/whhu0DYbUKT342v/WKx2sxbZ92ITgCRebYvftf
FpIJE89ePNQn4VVHW0+b/U8r8O5K4rgiQbGad3yAIC2O+C80HzRZA3iNDJ5haksDHbvvZ5nA88pN
laEKZjQsKbkS7gGGgDjXrhJmx9wvYjGGgpvjCVhMeqaWgPFXOBlNmFWe/aN0Zav2213P8TkLGimP
12eOCn7QnnzWB3DHwacCCwlKUmmV6hEsuAXG2mCohVSEcMxzECEn0E6yBEXHtK2owM0brm2AklcF
VRNjMNy15rQtNRYilRq7TA2cQ+8Zpum1xOf8WxARgPf9BG/jKftm5XeXBT+fvboC8DSuFIfcFoUx
XKKHeqHdUu8BGfoVeb/0LxJcqbZwlGm0Vm2S5K0VXsTEw1jMqgUQum5j5rtgaeJGTAWmzCisoIh+
F4XyNFPc9SUIC0IBPn3n1qnQfyRDFlHR+PZSYuuZZ8HjVizrQuBg/IOU+ODQldSdX8Gl7b+teuh1
+JK5Gk7Hzu5qVrevCUJefSnTVsCqB9CWQxIdlYXTXTHnuGldO1bnWZmwmk/TPVErtTJ5ZPsEE3lu
idRnx7HigqhC4VUabpRYJqx/jAcOJzB8iSF1b3bid+Rn/fjikifNXAoOI0B5yi6P19svqHyU9ytO
6vutgrzQuOSWCLzHXQqJ/ze0ddkx6n1M4UXluNtTTrzMLCbbhGNmxfhOk8jVGrqY1/2gC7qUdXSG
zp94mZZM/H7MPn7sxSEK+YYWADGQC26+b8cTDyeGumeZ/wd8XueyD2hA4ucg1WtmeEnoFeRaEi26
BDCrK1PCNsSAuqpRBLMqP//LQlnQy4iucNATU3kvFIe2NCu/+01l+XEDQYA3n9RNIywx/q/Q6UWH
qwCVhRYztn4qY5V5BlteMMu8X01PLR8sOtEQaqd8XovZK+xk1DJqb9Vw3QSM8ZVYFh0qtYDQpD7k
/XKTXLFawi+G/a4J5u6/i1qQ93SBZ+bfIej2wARWTXY2epuYs7NuquLOd+dnLVxTCwJykRDAAQya
lA9Qydrh/JX8wvUjRFeV3bcdN0QML41Pjo4T/Av8WlkV8yBgJLaDCTGvpzzWQZNCSVkqbd+Vaz7r
erbYyv85Y7hUpFXW7YclXs90heZuILt0NDtFc0CPS9TldyEqsmJwneoZt5RIqCNJO4eN2+vPK6lH
v+wyZjuN8Lodvf5rYKVCnzIfDo+Uoflpgr/lmYsfHwMeJla8eEoA0yWlqcY9URr6N23kiZUbIUAZ
EKkrUXu2sLw8XJu+YMtKoPTKXmPprM0UQySD/6JGgjdQ9divXquWfFS+WESvzgpXLf3eWBbsO7Ja
N7RPcjD9xgkOj6GsgKr/TMSR3D30WAOWy6SgVrJCqh0nNbnyOvc0pmfCzD2th623Vbdy5xVeJs2R
zMWdrv66Jt0NKowQc1xBi0yvTR96q8I8qEQw4a+cFpPugme1w+/OhSfIB4h1XlPCsfUu4CXwJzch
wzR0IlfyZkXw6AQkvHnvQF1ZghkqzjtL0+cl3H/rCAHUNJAqmIUX0ZaGH8pVBffEveuPcT4jVp33
vtctZqaX1Hz+pO+onj8zMgmGz8d50R2turXZl/KMbrKLhMhV2tIZt52j4q4UG9OHslLOhpHxpjmw
UThZ7oRislwnEWx6PWPt2PB2YbTgEgxNdB5dVlh6V4tem664Sa6EjTJ2T20Sc/xxFiZxTNHKVIaU
kPbDrUd2YFtD8xMcIfsp9/OoBT3IEEwX2RZDXXE3inkKNElJq2YcR2zOl8dV4JE800JNciJPv0YZ
C5axra03chRAy/IqYx7acA8yMsB0EzuKVip53uJ6rnW81lDlVOhM7WEGsJ3TCyr5EcA5kslswG68
5MnruUYu0rb4GUpW5d7nWcKhZ5f+cfcc1lIIbI+rrz7cOsRJ8K6ymx4fBznAfdnc76fzcQqlOWUM
X2JvMOY79XxH81B1yhAbfkj0GxjHMtjPf37k7YyM6RWclpadyPggoB0i5yMIYT5THG7Eh2PhaG2F
1QRt11jIomWcsha6uQPsnAPJCUfLHX871GXfWXPKPMpynWYn44jpke3fttF1OEGTPyEwMjy+EhDB
yLbb5YOcI59QhneKcmWZJzA+h1Vw++4ROAIWq8LSc+7W1nDHb1yMpUwWy0gOMzmrZ6G2ZKfSBHsF
xbESyEKUIT9It+pPxJuuJ5kx0SmSrktunLzor4vfNfjp01cR/IY1hLdwvo2xMxzt0aANWyOu767Y
2c1KL2OS2T41ZfaJ6gllkIxvaeyenpJWCnrgKWxTK1xjPRHXXgJE7jZ27snJObfcVUkB2ISfTLyA
HKwHUdPm0Gm9iJ1/nB+EnNgsDrqeog1c7X7RXHsvwgFIyut4+bWTXDLslOJJndmijva3DPXJtQSb
aztT6rYw4sTRQA1bHVRDmjwyymPMOlTCN3JP6Zx5MuwC8rE+LoAM2ly6PYhIhbUgFiMGM/ILGeCu
LLHaLPc/kCXQY53031cEy9DqM3+sZRZMxu0uO4L7TYsMWGR2HClvq5nD8c7eSbhzAlDBzkBKRKuY
NyFgC0lOkANxfrbNb1/o0itIhQI2joq75l4woTyuHNUaIhsb1k3+aYUzqHJmD9UkZk3C5aafOlvn
i7rUuPBijDhw7wCQ4UMxdJLOJ4gu6F+sHU6zOu43y+Q5cyCGnwbj4dRzsPSmLMJUyAGxjmc1WjpM
PWeq3WTvgoObq21xrY7j1Gq6axvn+lNddj0o2lBqmHI+HL6kyfUCDnqRTGjrqzuv9Hp4RcB2UHet
PUKjfrFsZ97yL/J3i8Q3yPaNnAU1MZa5U+XdNHjN+ZY3iSKQkBCoWletq9bLA8SOIXwup1xIbqAO
qYAqGppaAjGQg9qtexNzCLG3klWUb5R0ZUYsHKp3EFxpoQ3GLRcIbKoKKbKInkoILNTBTXnVjuPu
Jo+e7PAHhsTg5m28KwA6tahKiFYLvWxb8UhSjvjwvYE1OefQoMiIiHUjP1jHWAekdFVlWCrVt1QP
8NXuGKBMJflQuIeq4IIhbqIYfeKOUDfRN4XJhS/ZRDbKVUgwnCj01LzE7OuysGjDMgJPvbSpNDnb
born1Fl1pUyDJDAtjwa1fQNRTkaWBDSK57SaV4xeAFS9H2FIW2t2JQVr2kghSQtKz5RXMvEBfB0B
EB44zNYyRANx94snF+YBQEMXUbXbU/xJpC/KKfJSwsutlbca6rSM0SmraEwKKs57o6bvJ/8vg1+e
4FXO4pUc0LMGapvpUSDU3vZylPIBOWpjfyFsNv9fKacPHEpZoqdgvJ9Jb2B7bnBiKT0j/yCRRkRP
Y+o19qDFPXQUisg2smFPJtAnA5j3sAvYUdXjPnwshTxjZ8t/DP9HTdvn5qtT1KM81qPtzCVkl3Qt
hWg7WTu06mD/olX26V7zEWnbUv2QelHmskkbpwBbbrnLxRA92MZnMW5XchHXsJsYUX9VvaKPsO4T
ZDLpHLG+wCO1mkk/OiY0ADYq72K5whAlR3ZXoIu+490zICzR301JJcRlG/xaWWU8UW3+9eldQolN
HXKcjdi+kPtcoBlpHgSA2oE0NzHb0wp6fcfTR3X4C73lKIfJwVrJxP9yuthfhTPRuV8ZNunrQ2Xz
tkAfSbuR1Q5U3oVCoIBjSah5fV9YRhLczTvRJnaducx90hA+YSuf+SOTp6XqyaM88Pw0Do1Mn/EN
e94PnFqaTo14+DPMKN0rJdAgTktA54sBYrkZQoDLRvE1YQVex9K7whjKZ0KmuEWwdzCBPUlkEkl7
q8kPWmsip/H2sGW0T+iQsKEEoGmqm4ilo93CwEZ6vTPxizMHch5ijJON0sdlBmt15ArJHLHPCYj1
O50S8s+0GU8vN+Yt5SikDjahGlETAkYw6zNEH0AlxvdBsagdm4bJIPWKJzsVw4pTG3aLt6pepmi5
ak8aQHH9F0RMCbmwmW8uEILL0Niv75D/Hj0rMg+zXw2XU2iMC+WCUgthYWdGU1uAFEg7OuA4LXfY
1Rb76Tx9eyuEfyNHkvlVrDeibHDW+N7AS7Fl7BW5GpRJURkQC8RX0cKE2z0/V8/mjLuT2P2xnGIN
U0ObXXcoDAPKytidTEg/i8EE1Fq/H5JdzqJ3cKFl1JoQdbNNXTiTMTM6gvvGCnsSfBeK5vlth9ki
5OEXqjNPDkeMaqBGtIUBFc4ue+8z6BuFyQCb4ugvVLMH1/n6Jy6JvYQDY9xWx6YyuXb0Nqfskdo4
1Kr5vQcZoAHmraj/o8f/P4yCF1z1m8IDmZSdJWQV9oxZVIuF/tXsEsSQrewItEY5oUWD9Z+Llnva
vp9cXnpmPsgH7Lh96/rvZ87/0oTwX83ce/bhXuTNgFynPEBRda8z7Dsb97sA7luz9Rc18ZWqY6mg
2AxWloYVIeFyryk86pIXNZ3uRVDNxT2SV1JE6uW3/x4Y8LI70MZk1rK6LelElfIQoNc0I5ukCicb
U8IKO9iOa56+caz0amY5U/EWnTTd5uqrYT2CnVyCsL7JUdhy50mbd43q807BDAis6XS0MZ3uXbex
0IzT3sdepft7ko7xZyK1VmalaG2/7lfuze3JQUTAHx1HLRG1hR/LonFSzCvKp5SiD6NlF+tKsZyN
OT60Slpe6J6Z6vH45MQZ5UO3cjXDxP4zPier261WsCzZwsw+Z3Tn9x2OfnE1+nkOwehPflaOOMG9
DV+2H6EPwAf83gC8biQlQG33ay7VAno4Cct8yOkhzNhnCjqDRSI2FseG1J9KZio9H6ha2ivfJBy8
wAobJKCfYbvN/Pd93XgO6NQxKi0bvVwY9RtKKh+6FBWqcRH9SNzsmv2mdW8RbEkhn14t6PWM25+y
hy4YcrixULQFW3ntmb9LkVIe1epZKJBiiahz2StMOd81WMsHoHNKghOeZmxHIO4a5iGJ/ql+/VGQ
tFaDmqtjgDBNszHlpD716K8s68+VrHG84wa7NdZ+e1MT68fZU8FZnpZ7zxf4ilzbiSMkW/WNAJlA
d1DUv6B0XkRTj7KvCbFL5kp4op+rK0uM1A2ikCVUwmXwKx6hKa4h/H/hAq3I9Spq034C/LbG++xG
LxGBicD9yn4iigOrSHEHs3WRnyACv96IOHBRX4nxYwblHBU9MQPdWZOVA+NadqoKZvWh17WhOBMi
0PZiOgTGlEbOY6FBd7R293xvWZ/JoZFcKlIim5bzee6NLuNLl4oOyn4eiAmOsJq3eIn7xxv1Cefn
OHNIG5ypHoTt5ozZx+1R9nMpjCqf8qq2ufZHD0UPke7Mgna1e1gV78fUIqNT+tlqBfwZk8s6Tp1V
QGNQjQ1ZnFUQQ61Gd0V+78EH1MCqSZG0W9LiR06R6NnrJDBbENaqmWn79SzNra23UDAy8CmVLWzo
RbILGkK4CfFPD/7bV+zHg/QCc4UozC1wyrF4uZyXr+WO83flZU9GEtoAbrq+qor/ppKan2GUV4ix
W6zM7gGxIOuER7LgkHvy8OgQbvpLpbDJWqiEYPyrbcIpXAQq72lguFnyD4MYO+/Cr9iDnrJ5avis
CFjU+18JCN7DZtWJIi/6LOdZP/Atk1hM6ZfDoYhzWvvCH4J1bx6gMja2DdNhxnAlWCf9co/YESYj
M4WWS9DgrBQjOxfL2pGmHZ6/1w5NFrUJW+vk2Nf48qzR3pXB/zvNf5p5tGyZNF1/NAEsf1HJxkEO
VKHFnFHpkyXGRw/LMXvf6OqsSc3GIB3omBkygUUj6eZYByWDpv/FvejHNemWPkrUTNaA/AQvgZbR
GWJ4PBvADuHFOjHlFIKinYUX/IOURpQuYRk3s0X+g483DA9H0lzLmyZA7wY9+qNpzf/240CYuhJN
SKJfSh++AqmY70fD+SIL4YyZs/hZoB3unnMzD65RkGbwWvB4E0q8aEplf0Dhd7NCSGNLRHOyqY3U
+xV8MIWpFCSicoeiXzuvw2Z4YSmp7b2QjEtfODif6EeTbmmozhxSFqYQLC8jqWkeP0vEMz2fTAye
4STVbpq73dxLNci+BDO8rlR2rokHOswChLWl+SGNYjPofK92fuQ+ETsjY381V2E4bjt6IPzDQJqm
lU0UJyTZez/HsJltfKakevXv1HTPGzkp0RjazXEXm3uQHSN95UHRwoln0tgGbxp56EblAu6WLKVy
NFwq6YusAPd1yvIAtKekz1cX10FfT4Kj8adAUab4aaeB63WSq5n4nWEU9NJhyrqidqc2vfauV9VQ
1XZpt6KokFRhwk1wHg37aEjvw/Laz48LpYHSzI2NugkDPLrYY4No5IAI0HEbCQaaBQKvtMeJUaLv
4pIdGPkKzwI1JN3lOJC+EgbQVq1esVw89h8gY2iEJXlLt0LZlemLye+mf0j0nOr0+LcwtXcnnPuU
PW9rH4JG2ljsPMn9krgcUiKiVponN9sDKzJ6riKJRVo9hlwGtlPUfG5aiAYWeSWDerWyxWBeJLVK
ALCjvWgALgSmIr3B57ukDhw2NogMryAJHFgj5+EgYCcLV0nd8lnGOLIGnSG+xVY+p/m3DXyViEYe
c+EB0DfrS8hSjIETciS1jErjbeJc8xsZjZ0vW1DL/KGtCr5OmfH1LHp5HUzClDojIwyM2VmbdXww
QOlHjD6UNclu/E737WVjgj1l37MtC8Kpwgciq39oOLQ37/kPm7QYlZNFoJVwqMJEzUaBgfy2HfQ/
GpBpgqniWXZu43RoqNls8uhfmMFeNNyUFvIWodVgMzKZdI/GpVm+YV0Q9h6fvZ8ivuHcaejoXun9
cKzq/gEG7x6ufapL+EEW+cgWmkh0LXQqFF5cWEqmeaaLkjk7uzfF6aFCDFArNNDb5cjurzvggWIL
HS+9BsJBKbkoKKiBYAj7XnARgw56hUelqNHPl1t5ysO1Wleg2mkn5uJb/Tf4F7IxpuZKbdYD1+iB
oy4OgGqUlu+PTTRO2zkPb1/TSt0XntMZs4BXmeOnoP0KcIBORdlOJnHfn2FmhPny7T7L1dzyBEbq
2VU8RIU6XOQOHzr+qR3KUKmJFNBb5+LLgz+iNiYEPehT0QVN85+bEBOrGcdgw9Gf+vgnYx4boATI
hoUmAQzccROvyf5aEVjk2t5c9wn7HAs1n9w+BUvGenFD8Xtq8Yfj0MtT1NL3jK6c70TG03vakyrt
L9pfGYlh9t6G09h4gsyQUoUUuRpvF2Z2DrHNdqs2JqXzvpiWo4F3J9ylWnNEeYupbTRNG4Xlds1b
mFnyURTZJAtBNmp3xQXjyXvlNOiG6NwYaNgaOh38avgOhBvR50msRpb1L4JuZvaGRNKCNKoVuLqv
Ks8VO8Y+wWidkD23abAYruvqu49L//xLwuxZoLO7+tag3LJGIcBe1yK+Oh33gA4PbTjt0NSXO4M4
IS0+grf6GUGv5dSPH+RekJ2Vf3LClmth6YlZjIrryyqBy92nfdnCxFn2AIpHYLjv6qzImh5g4Rwa
ah4ZQ7fR2sL+EkifLfplEyv7uEmd633UyXpDBPhmUvjnhyqLZFKWD+T73O4Q+GcLETbA9c7R6QRT
WrG4Nm0x7+kIqeTETjBdBqxsOJ4LCbC85yohIorIr2HRiOOoSKlOohe7SR0fVMSICkNK6XoBTbpU
fkO7+R0ikoSpXDDvN9JlqSybRO6kGNaGDtRRRXrXmLaNC7bx56WwrvU5Ibt+X1UXVNTyKhd1BFjX
kQ5dWxf+kC0QpAKd3bw4s+CK6mkG4qf2Ylt4v6sAmlMM+xQHKfOMEFUABwS90N750RPlau4iVEBV
S+eXrIiaHvcf3jmeJNWAojdgEK0Bt78oB9/aAI9q+zbc2r+fOzPVjqa9WGJnICqON0dSn+u+anz4
vIfMyDBxVx6rVj7q3YWqu0upasTtrZVb42f0c6jMYHnA1izOKKCjzxF7nAzBg3FE6MczqYjF6mOF
hACrs1osEiU4iYOA13KVFG/0+gM5e/RqX9TxhwP0+g6W1/MMDDZTuUq+twNrNqgUk/1zAF3gD7Cr
NmqhZ5nOxJZVWnLC86hk5o5mf3oqZPz30+hoSppeLRS8H16/RCZVYqPUWTxsWFBomUPiqoyvH97z
hV4vs2Tlk3rLxs/pfz+aaMvB1984+f6AswsnX1nPC3rvSM18vX+PrS2ZeN6awk11EoVWIN9tsoRQ
EYhPKwU9z9wIFmCCJs9c612iYR9wHhAysd87z0e8cCSc68P1oARkWYmBUexQAa5LhMaYFIGa0gWg
4EQvKhOIbyEntAsC5NyjSQQlNy3dMh9Dfl1cet05vtX5HCOPg8Ckz4Joo0qbcNWqKTE+qCufdnha
7yYlzsrUxsQSKsRZnOcB+4pJzL1MZq0aA0cpjKCB28O21OIHcnkYP5FzXm3nkun9mLngUeZHFasP
+tfC27l79jnt+QoI0dzMQNBG6ZobxIV1MUZsel6i3B70YRfvThfwM8IQIFmiqBIZvc3PhPUy5RMK
LLSg+wGuP7Nl6vLy0gK8LOGAfv9GRbnEII9Uk+LZ4P6H0bCIE9Xjone0eqRbz5cYzk5xn+mnZuaN
xCvm197OnqnJ6jEwicG7dp9UjYcF2C/PYVyW3Xk3M1nmtOPScX9aLu2iBMy+KTTMmoIHNaReZPaJ
VW9GaeYB/Q7eEXnuAlDDyE6fv9QBocR6sz/Dm6YdDuPeUGTxeu3VcaoRN0bQ3HAhiNLU7HAKsOaJ
pvIony+LvJ6WS0bBBkiCIp5Vym92ldxsK3EGMD7nfyeWm63D5kpfWkEnV8tA17fmr7UpfmwzuMiD
7lMsi5xfvMvJr244Z3NMN9HrJorXH/6WdnUgYA63gZRyzhYvH1i7nWaRaxztBtK+yrzCHsKKsdKB
o6QxSOjAt171UXOXUq2+b3Rt6acGL7bEpOl/AZVdtz3chzlGlD/OWsu8DGbsqPoBQUUJNcSuclUr
GWjXsAfllbhdOOYPovj864Fp+et5tCW/ZFVNi5NkAItksJAr3X94kKwWf7z2k3Wab0DJeOTpF+qN
i7Aj0nEBc+83p8wzE0y8hbQvsz+iTeemh5rceRYSaBI5dm7ErQHSPesS8im2GJrAUxX/81tmrwnx
0EQlgtNvU1+gzp7mxlOFXFrKSiMfzP/a2A4TtStjYoy0yjLQ2ukOmqCzCWumlgOFAqSm5RMjRSyW
wcl9Bv0m6sUlS8sbJ6Txo9DVxn7VAVWGWCboLtUXDs21EVIkR5/opXnntgHqbWoo2Zo7gt0UwHy2
JEMjS79tV5mhBsIW4LMEFdlfAGdomDOac3y1d/n2KrMeUHMHae9jE7bWaK6EHxE5MBJLRDo5BLgA
RXsglNbuLyckce61cBnXmrxNSZJEu73TEj8+t+A2NlpaI5W19d5aX4YpcLQnIwip3+iDSqIL+JRW
ErxuILTp81/F5ji/6LCdCRjH2TI34RskHJPMJID/2YVgxO0MtosbjFrJ9ceaW7Zkg16eTf1S7L0s
+vXf0iz5RQU3Em3Ekar+VekCUtcvay3PzSgoWhA0JJMgGjI7dLoc6tlkTV4JJFkwDSgqJpyJOezd
SPBE62Wza5Y7h0I2us3c1T6Fam9o0a9DvRAQ0ZXuwkwGpZ7b5zxDRf7T1Tk02KCxx3xZpN7EE46b
lOUqfCNPDmFElJpCN11rh9J+ViVnZ+tQjSoXCCl6/My8/fIiO9BIYp5cxUSvXwLA9LfTybgVV1RO
8Iqy42KdahsllfvNuGLlPrzIuQGhzqVcEFu/Ahv+vIlEG+LiUzxmKVUMhh6zVKll/Bh8zmUwFrui
SKUnEEizVuKL0c2plyu1p25REJ9Mi+nD3SY5Pz4Kzou/6QYTFqCQU9V4Ic2L8GGutrU6P7O+jUq7
rj8wd/PxfAJlc4J1f2TYfGKg8AOkVv5ZGTpdpqMx/S5aNk8KxKYYcKkIzo50ck6VhzLCEUH5zm+4
I7dsAA3dIcNVNFxCAM5loSx7XU5TrAZP6ezSbOnSHBy3D4u319Mm1og4dINCwkItAt0wjYxU5OQH
pW4u5CnbiSENtNkvTQnZDREWHksHPgH5NJLoYKCv/6dpZTNl13p/YPoN59M+pY6J00LlgzX76rTb
sVyR0PfG2SejIPtQ4IceIT9QHOgGPalDGiYSE0ijF3/q/BokL0now73lIwwK3J6q0XmO5rBXtiP8
28obpzZ8aRNkIE2m0oqDi70P7GQ2PBK+LuP4V/Kt629Zq5VvF7EbXRbInWppWtf2MuN5bZcJPy8x
z2MzAyTx38sPIAohrJkDUmHm+JmHvVLmZ5RzrmO42fNVva2tG0l3s70lmml1W2wZJm0rbn1+p1uo
JAAGCSbUtKP7GCJGOfvbnhGuWp0rPPMTtInZULr1YAyIQAm9uruYdRnQ5XyCBhK8GYO9wp5azbND
9kBpgdiXpkZl2UGWkv12mNuwDrZ327x9AoCeRoWuvW2RPmUotEzMChPxKFDV8dSoORsWqYuTGyss
j6zTVFdzc8Vz7JZ/3TGgSQKLDEFGuaWZDOeK1WcIsznSwBVimglWl73Vpkrkhe8+/h/cSbK49dV8
fIoAgUxc1zvGlo0pA84v36w9xixfSjlPK2D5Jz3paFsbfTZvjnL1Q/8ypYBs19VNCXMmFk7Ql+IO
ygUZgS6XEC0VUN1nkS1eCCK6c3D50pCWBdh+NwaI1o7slX0Ha8JJlB5/shBiX642HIWtxKHYco5Z
VRGhP0YWO3ow65XxqEs2OqH3O4ocvUfrAgdQlNAI89GaAJ+j6QpEsSh9CSLmw/wO7Gew5AuQUZ3l
qrqLszQ3qRl+qz36Py2GOBU1mW7uZ8cO33FVU2mSiIuB0L0nMaVOmeEMyMp16vH6/E4VwG/8TxVk
cW6PET2BDxac5J6Adfxn/QIQUlIjPGugT+s4YshitrHRofZst9C728VgjZhuKnIpilwrwUoQeLPk
qqrcq+OJbYJiD+181myn+1Pkx/v/L55QUwWONYqNWXgtOUF2FNhxzbgbfnUvfc9xYV1l0QlEjK+8
/98AFoHz6lPCpSh+foCDJRT2zaSsemUP4ZGpHMMUTvgWC8WIjtTuEl51JriT1OfOxC7bOb+d+Pnf
UuSLofMvHZ29TDbw4rfNShqbLsWs7E380PDpHPzrek5nRHtRLThCIj5puwkmA2ppPYNQTIw20Fx3
Eo4ft0kaA6dVjSQjZs30KX5erWST9qa1CJVJh4L6gU1/xgx3qPia3zA3RMoLIIbt2CXTGNVKRMV2
XH3MfMxi223ZMYo/Xf5W4CcROQfKNfh3e0QwyPJkc72s52BbihlnSR5qcIWR8zwN8Tbpns1uBMz6
gInD1PZZ0Dlqrq3VjvLYtdz/5XbzxH+f7aPmKRnpCQL4i3FYOiQPMe8gRMHs02rCPNR2lQiS1uX2
jOA51CeH8S8IXh/7XBC/f6UyjW/Ps/XYLnhMsUtwyD0obD4NiMD26d4ibLI1XHN+TMVAEo38fcsb
xcp1VWXIAeS/IbLi2mgQzepiD7Bo7bxCG51LEvSu9D5qiZD8TXY9CWF6W2El4VJs8BhO+BRuniyn
3+nW4vATU6XJ2ufY1Tew7wEJxHDyVTgPt0N05RG/bE61pJccXomuNawWphYQs47iDs/c7HNTLCX7
x9tEnSdrwPZb2YTljQZhKgQRKgYEaAH0V+DB+wvMOU1MsmHzxlktcE/Q/FSlwuDrlcfKF2BOW3Om
zZb06RJfGl1s8xDFAKDDCaqqEMYIsSw5oNeNZzOPMp0ie07w+HhxHbi6BtJ9uFuAB0z03308yDVw
wydj6Cs1irStfvVqBsVHbfhIiVBEQ0v1JEhMeX5zNJEqIluDWqQfJ8Qu+MT0JYCZorLSurWNqtwZ
l0UiF/wOCd+W7xoMV6UQKKwjjkkvBGrrCRi31YLm/GcDMwp8M6v8lg38d77+wrCPtTMy81ob0hJi
R92en1IoQMXbOB8wXlXbPE52xnLVBc5WpFbECsDZUoiv639VomuQ4j8xih7O8oWdFEU+sDlx8e8T
/06luY7lxwT4P8ekHCrjgniCWeQDaoet3Jk/rtsrteuNGFSfP9NQ0aIEczjh9Dkp+9h/JwGf6UZu
sPtDTx02LYUxy6iawVklzASLloT6E2NuluyleHCVGJpjIBldfnckwsd0r6Z8o301rNvoHjeFPPgu
NijYkgPmLB679Ay4hy36GOU9ok3LZLRpdEJ4aCH2YXF+tMg1FbFsQjazN+RISP370vM/Yj5sLV3O
8Q9iITmosBq8v3YX8tlzfypvh8y5zqY4eH+qMT2T4eluDHEyiGPhNBiz9yf49MaaJlwCX/sLaB8v
7qfSZnDontHoqozrs3I4WIkfezY3Vn2AR2+PNADwcWME4KvcJtrPyjm/mqGmh4Hswq9C4vxKLYsn
L0VsNXn9LP8NLbJK6AhwtrYsDbj3P+iXP/OPrqzmc/3iFfHC9Kyr/R3fMG0LDkZ/7XoASEvCM77d
AVJ/DB6nqjvEVeoPzGu7bCS0eW8Z9RrUXcWjqL4+8ho4Hrr8PSeghvTDQlsIncxZR4PG7g7ax82f
BmJpgvn50Hqs4QND7sRZKbbWolO1AUpfxJvVOqsOJm/yC9DTfWq3k3qZmHhhh/aOSMQ/ycJxRSRI
xsacloUagqmr3D2Q+FRZz50YcG9vFj/Oc5AB8wP26hpimyL+h8H/ofu2/O6DeEMuBOzXPVT3Uc+G
uxEfP9fLHWoQsx18M9SxJaUBRAX63GGpm09r+ryoXJXVBbgRWQjVG4mnuIkaqyxEkUs1h0uLkol7
xoTCzaN8t++Zp9NFKYxfUvz8VdFdvx/xqG+GsTGnBRzdeuan6nrPdaCHO1Z8Cl2DEPo5AzqHCKW3
Gcdf4qizDsdC2kIrB1rMBHD7HuHtslZ+On4Tutn2TfNtnwU5wiKUJz/xIK9soQF9nXMvyb2oY0g3
IYMiEEv92pD5N8TSRKYwvWqfuAwyBc0dotWlT5ihLNBypLRAIEWFkrOlcG1Hu4+rpJl90e2ZpOIp
YTxXZ19zxZ8M+3TotQoEHTQA/TnOycCEP6AvoUB2q7aREmmqzKWKGG2zJ49mvbbb9KgEiwE35M2n
mSjNgEwh9nUUT58iE3ZuvFK5iCWi8M3QWcJk3+LWRp5OyZw/ui644/lf4SR0KZUvgdnxI2c3LlNX
+aVL7hGBSAA0zpANNYsslauWJvPGYNol07UNS01bVsHf2Wkbtb7KrcP3Zu8hYu7LItWw7hppTHti
Tb16VDz260IjSwCVnxLGRNSSjmYu4Y/iKxkz+tZ1OIaTPRYCtQhsd233K3RCMXXdMH36c6NdpoUF
s/8F7c+llZNef0aYi5+70g10tyvmzLqEOpitU79uG1ewnxEWYhrJ/j+64/hs+YVmoLoUp4IUNK6V
8ZR6Zvh30KubC6A116cqwDJhKUG2lLcUQiKJgWOvkGvMa9UhaXM72owM3JfzqjcNkjk+XMbMeujg
Li6lmEqdF9CmvyygF3XCIBc3yfBZdfUXMnz/WsE8uZ7/1lLeP8rJ7AWFG+OjCtYAgQZfi0WLPu+U
aFxBKA7OZs5a8oWnBhOqLDM+aCyHZvpvy0B6MDGdFoFnWC5xXWgmRh/rykzmktcObZxGkl9VuVEO
tqheOuxr2Yf0fkoVdECRDKnE4B2lkulKtSld9k4CzmwiGRxAgWNDH4lEtxMS/NZKaScR6JtzLITa
nihWmypnLngwyEfcVdzsqhKIiLT9wjP9bSXTHJ6qniqUaJJVGDa3Dl8hqGWm1eIeUdviVUV/9nTo
HnSOpgOtnFeGMcVETSd+Y8mpIvBD9YUnmZsQUzWCNnoHxpLZUOPoooG70uqkqC0sH5l3YQMQXAZ6
QA5VDIyGOtJUeqfOF53vJ07ugmRLNgiYYl+jH4a5QffxIZpjQg2xC/RT+ERguiTb1sZGczEF/7Tw
xtTdLLyKAYSWZb7CSHNrYrg90ZfXAqubPRMWtHh3H0CfPrC+DntKG/DCuz41CyJ/kn3tcqN1IQ2P
ifN8FzaHtv7NBaVn1roQUDvSP5nfTBoWXQFbyERnQegVm8TYg3frUYHyMo/F9NvnHjQ4XBtZ9M/Y
vRfjYNfIrI0IwU8zU2cbqS+kl3QgZgRerQgVAa1RAiIQfPO5Ym0pV1vcvh7dg0f3F6t9telyvkZ5
u8WtLdYyU4mRyJNkr+48FkaZCpv5Bk5MSb4CK+8cd7qyMiPxw7HpDDn0BaZEeKysM8SJt23sIcAq
PHcNfV4IKWjDdnaYFqDZI80Ym9gzTu7B5cxpR3gc6sSXHK/ZHYer3DQFdtTBTHq9zWDnLERQMOZ9
xxUslZLwHuz9skBHWrVrjSwzTMdXBCkkDsLI/9u5314xiX6OU9os/tGHsJRCuQsEmQMEkf2j//mS
yFE66Px7irDdKV0aCD6tASRP7MpWl2oArZ2Zkkl2MQWpVGDW6rC7q7sKcoqvUvNfuSJJVWgBPA3o
f07ICKyad6MZHyQA0TdZINq5Ht64qMnnsSrpCAgalXe+YtUXVuNuejSD2uTQAp+SPC8xFLn/gEt8
vsennKOfQxZ5SQVlIQbpJx3F7EJjjlwZDRBoTObzFgwpazhDFo44DTEiepP9TsHKGfwdYL/v0IkN
Tfj2j67nwnFF5pFeoAF7gAv8QmIWsUMrp/uQtNPM1w+TO/3Yh5/VwLVJTMb5KcA59uCxSAVL25DZ
h0Md3xFRkgiPKC51HN4vYYuqpxPydElTOXAuw22RyOYHU4mnB/o8QF/R7LhjHUCz+lTabtfVybXy
+bBmLsecc7OYYT9ml2kAoMqze2dab0ljtVXSAWCvjQLEEGyUKpwSwuBvYtVASzzLFF+PivobOWoY
SWWDhU4cVVBAWB6xzJFR9wrSCzf8zzEPCcmW4GnhzMpTrD1zgALE3EQc7OijXbKMuGAxQTvg/Slo
qDy7Hi90SidxLpKwB8zkXYQbPh3rnIK+Uagkq6FeVUOAUb4JJpgQm7gL9I3e34j5fadmo/sfQPT+
yBW5lDHjcRFDsnpslq5pcmHZ1dPCOPtc/EfBy3oPUBKIlyZ6QXKnXUU82mnT8oAm6YB39gTkPczy
jeoOh9ZvHtca3P2kyD7ocscx20Bhp5rTqFvuvTioT8vCduDX32tlW39g3D72NRmBY0/+ZGo8qfA8
1iKkmL+QHrYNkuKuPxMPFVoV0VQvcmG+r9B7z8IJ29pGZRnXUyz82x6J1Ek87ytm1Q8uW+z9B0s8
0PwbmkdoXzjMvupUV8wBQ1Um7Pa2pkWTzATcYgoAh96fjdaHjM6mhH1NDKYOTVb2wtZ3HYMv41dh
v7tIZ1WDzg34OrvS0426gsbqqW232oTAmAQ5j9i42ZN/fd9ur3O+pmFjT53+a+7mWkzeG959mKND
DJPJMXZONqQDTt53km/+Is1vhDKayCY5tDLq0pIoMM/Ji67I92hKS/p1lnkAj/GEoLzbf+KvrqXF
1ew194FMuIYMLYyOMm2ork2VbHoDWgGeGYH4a/q4idrzVbNKN90eqSpXK2vtER+ycWxk8FBffHw5
Aj9o3BOY661VDSRSSNChDuNQHOU+3sP31xD2Urvk7OjcO7pqdyKvOgwLqtaGeOXSP2YDuirgWHEY
IduQ09WZf4lqlfVN2pXzjXJBtWMdTtoz5U4PEOnwq0vC8BXRdDQQhcmmrueCP2iUibq1WvkhnIkw
q4zrHLmTBJBSmw6I45onrI2hRC+X2zC/xVWhJPz6Ly+yVu9r+s+T1G+SrW1tzWrcT+Li1jdkZrhs
XE/HRks+tegmv12WCh+Lxl4BRB9FgieflZj+M/OyVDDhw/gYc+YRWSrQqEGU38ImswlGU2C15XCI
fLcxT4k+U4W+kcwKE/lY2tyzCR5XagbIHF04daCdZakGZGPkmAcakgq7JUsu7rPW+m8nwQ4LfiOX
wLsasg01B2PI/n9uXAi4o43Qb+DbAVffGfBwGA1scOb9Uy9ZAmJ13GobWur8N/Zo7r+UEOWUpBZi
VJUaGd5GEU/aFIuUVZD4j1AFIHbIWNQBGzsOp/cqTifx5ohtwEQEjtopV275mdFHghHsXDFzQH83
yVIqbPopcuen697YV8s9sN4ptcWzbnER/f3kB2CMQ21MhX9TKwjkLuz5H4qkxWG4aI5Mt6YPzPV0
K+OxDV17nhvj4gveYnbgrs6m5fv9tGvpsWgggGbMwsm5DJKsi99jYvXaSENrLbzz8wRaahiN1I7J
25gvRTCHCgIgqFYWMQsG/nIgi3HtRj5u15uUKcYuohT8DLCu85TUyA6S+2qIWcn/vQhV170KrFAz
tp0hw8QgTHbD8suL63PIm8TpFwYugCKUQwqtOwmFXocBQKkv5HEMY4NTAIEpw3ZZO+bcb2NR9EY8
43YEFNAHDFQ/vEcwdFM6cGr6mPrcK/TjeUaYVf+v1CL6uPr9t1wzIZGEgiRIhbKyrALEoWj/neJU
RlJJxq/zrsIh51DCS/9hydpow6O5gX7JpbyRs/jMTqXFiCuFRONLrwJZ6g5gYYO6Mg/up0cOPO9h
j12/aX1TYSbEqp3xGUAKI25xeSierSYu8WTbGe6r24t4akbPLpleI00kgTJd9UqAmq/f7VZc+1q1
DRHDdRo9LlNOJz+wjrqxJogI40td3UUlA3eaGZdh2WpPDhKz0X4nVZCXmQZc7382TRDiEq6OD2wm
aEaMX9eYeLX8ZDx5sYjNR6mMFQlMgzmPC8kQ3gXbhQaIkSLv/7Kek3kssHPaTUSiafxdKMEhE8JH
yHOjL0NEWK6/3PxdpABPI/r5a4QwLoT4lkILTwArIIRxTPALF1GWLkawQoCn8Ubo6RVCpkEr0poE
RvuhaiaogF501thrZmdV+9NEI+CCFYUaVw/q1AyLD8r4mvxFNvU8uVo0z3afzGrSicsoEMCfhsN2
Gxc1ZZxqWsJ3DZoEfCQlaLlt0+QNX0c2OH/QYnEq8hvc6APuJYxjknSD94T95VwdWwXT+OFnNjPV
4tKmMKQqpWk8uDeANVnIg6UDAWPK7zdMucC1ORySt3QqgZwcGhzeTAxpkk8EFfHSEW6AAb8R74vF
MpKD+8FvbSDjyY09pV44zuMHUGuIxf5pGjmz885tERuRQqZraxpqtlO0tMH2p7Tc+1j807aMyOJG
DizrttWj85hjYJ/j99Qfks6Z/gFo3Rt3i9U+7tJkRUGOM/V7bxY92nUti/6SFKqc768K+wBsfP8s
BouyB2ePs1ffjgNaT07bxvSNgUPHFU3JN1RhTtzowyxQmW6aJHdDQwbCCmkUtkubWfv2edqKZFiY
pqlKGj0Kvn6ZyJLulSJoPR6WBExWkFMawbmYBwecazs8UbxyZj1R6F/vkif//yOtuTpEdQLmk9BE
AqluDuF3azBMk3xj67a85LQUDdy/FEDm+solYgyUISiNkkTRNCxtH76V2XMkl0ulNtERsYFUPJut
ebBHDBvTK8Kqo79eM747fOsCit5LIWeDUgUaGFKLQ80ZG0vxqNMEtWAeqRkwpLPxxU5ukBoPDbec
aKxLPbh10B2BXQJArnaIRsfWv95gS8c6bh3gurn0efgW77HW1AIxND9fBLyP0vhd5BmE5+wkuu4G
bNsx4oWtf0RVgguRD7twprRgnDtX7YbIqc1bLt5XW8BR/atATVcOAFrXkNHvzwXQg+V6HtwVlt2G
HeHSggwN1RdiQ/NXlsgd3QlBHaTu2pWIJpp2ZmR2JCIeyELXWv2Stg41+9YZXPN+V//o7YM4eKXg
oTLcJ9e5lMtU4ftqxY4pbuQaDxsYR6EHkMlWx6a6rXGy4/sxOxQuLtoa93jqEA3jC+EXiUHtfU4+
VIazdNjxSGNn+MbARzCDBl4/azRXSK2eWaoonyII/dsoVhVhvwA6mxEcVpLsHxqqfylDYci9PMXV
jc/+lAIEW17Zpjixy7tmOifc5eF+Zt2uQ+0utGGxoqBpbRRiZqFhPMUBXBpkMqcmKQh+0cqQA05h
PStncJWi21nOGkkfbECs3AxjdnAtWjL0X9yprimBok4Qdmd9mMzbbjZJb6UCMxGahLYUuApECa04
XYGq2hqA7L8K8uqLUwP4RKbaDOpCu1MYEeda8X4/OspdSqaHrjVtzPh4vvjbpuDCnbG1dzTq8ssN
sVEmLWrKMhcly4kzpH7WtpcBleT6WGkkcK/0P20mynZIrdjepinNMM3OKGoS68AAfrq9t5WvzeOs
1/0MgagNO4RdOKPObLpKlCLIPAdmhj4DF3ngdMw/PLlxpXp9r82D38XEBpEhx55yl3TiECKMaRRO
LNwXLMtL3Ic0mKxU5pBYLIZEepM8fJjzxtGk5OzPg6jRbHWy+R/xY3bwGU0J9I80THsggJDLkmMQ
+M3N49qHXhyFiqngD7aJw6752rBUp4EdQ4x87IfK+/FgvMlIOiOY/CoH8nPJIrdO95PqI4p6FEI0
z+SMZBXIB4ifOdeilIpZpNIXp1/Uwj2DqF44fq+n9P62ckJ6e+x9l2EaanogdNojUl6jxy2XaS8E
cZHvX9QV9kEh/ISPplO/1Vrf8cGoSAbYuz9/BkExduTFIrQLPR9TE+a3cKqYzjWTdXgX4dHg1sUd
/stYc552B+mJztiqdZsSgcFb/ZGsc3ztR0Lbj7kRZNKH6R4PzyV56By/fwGEjMUXiZFGuYN4SPx6
C93ROV4wVnTRHxuxr80uCtci9Q4YQy1305a4B6a/5u1p0VpONy2x5bSVV8XM5jQzpBRtf5q4ji8j
V/SiLgYkkdWjSdCLCtf/lOu5O+tyOBF01cFcJtSkKp9yvyVGkDPXSPU7pCkK5aLhZVFW6f0ztfOR
Dw9SEhZ3598MEozg/VX1EPZ9rF4zqLIPtktVauFIOj+gMo+Tp0DzOp+HP3FRCVYZAuX3Uq0Xv7Hw
3YbEw8g1kR1Tp0PaiEoK4vYPGgAnhqvoiknvuVgAK366CAjiTOqBVWQvPQHHVcsl1nN+rJYvPXBY
pVZqK7Xx65UnUVScC0JoK950NQeaJGg520D8AkzeuP27NrUCfXzTde8YNAqHMOLRCgO/qYzJMTuF
GEhg42n53zCoCn+gKEh0cGY/bVOreDVqm71LPPoZYRfPKzpuRTl8orNSTbvcB8BnrF2wkDNzKpyA
2wKUlqf2R/DaZknrBrEAur/XM7gxm/WBRWqfkhWyub+X7PY21ZkjjvypHKGBRv6OdsL+tl7ZCJ4S
9B1NJHUYJp7Aa8Kp2WbPUpjGCwS+Porgy6wbwRbIrIP/RKvhlyEKNDQqYYLXX3CJ0xa0c+Ljcu4u
rDOzCdCguvl0plo+/qRytoM1XEsasJnudsrkFXE9o5u/PxHAffLYfUA4xpbVOUCSRMsRKX1v7p2w
USnOqipIYByBUNTB+DS7D3zLJNAZRmgTbwtPEaRiqcrWCK2s7AoBZm0vPHaQdY1El6y/qedFNfCL
fVaqzyIZ2U+BlAPOWYE7brH1maOz7OkrCupW0iPCr22vwbK2LyiVt6rJWxwCRWoBl36SmQsR39pz
1jVTfwsOYo26HWVEyWjMRyAQW86Rt1K06Ajkzd7Ph8M8tNPMHhrTbzN+ahTMMgP5qtT4CLbkqnJJ
P4g0ih8/iWUILTHEIPHGvztycw/WrqaXEvRo6DxPXkB9VG7yMRfpRo1UmhZUtQeQ3QRte4D3r+6e
o5kmmg6kaVdIfKZtDd0+Yh4NMnajeIh0Ix7YMi2M5jv40JgeCEwGHNlAOwgEQcpeXh6oTe1JL5TH
FQtc5ujltFn53xGqBWSHuXuYjP3KijUciXN6Bhkm7XhB8xPlDAgdEEgDkxlj0zmO/1S2LUR8s32L
u2ZRMRrYkrCJjhiSvka11W49rVniMf19Pcjk5cwhDba/rs6RPxNa5t1Yj6nplv0AzG2Gs08nSPaa
Nyz2it6BkmyZ/XK5iM1iEjUTGMZ9Vev5SoxxH9Cm3ydGnQWcw53OUdQIMs3lwmnLdQiLEPXRFODb
Cr9tLSqkKutiAsNiKMxBMkOx3VBMakZ3R6i23Ujqy0ji71GjGYqaHO39YfYdON36ij6+3XT2z8pt
2vGJ9hemBeWHeSpeKMFEm1GbWcZ01TdxdAVdW4NWAXDm1d9ta5u5+6xRK2/dMXnXvdeTF0HQdSSD
8qXV6dZmqjXxDQbrWFu8VSgeLjrLR84/K0FOb65UVMy0B9lK2vKUDyQWEgwkgBkHJx0sn23GxyLI
LSEG14oxQFcnWEO+ZMze7brQ8mkuI819B64RtdGEvAjwxDt5eUwILC4LtPCskA38f99WKwWwIMQF
A/0NF5iLNYkk/s0QFVZmI36oUnVP8sKW03azT17iQdEtJ9NDfWIM2I4Oa2msFBBymb5g1vbQ7L7l
+if3JXmQdJjZv6oIpuOmmZUSvhCE1F/Yx0ydtMA/1EiDYsQ7OPW/X5uLB4V6xw0UhN5BEeU0kgAc
Wb040cDemErCykY/nE2oj1sERJwTPtXF2XLcgw2uQkQDxpsmeLY7soA/31b9BVkGbDHeazN+nlLA
rspOsUHWYUqWVSdBgMo4MDZTo8vwUYW7PazSmjH6GIxSC5htMc8JqCd39Z7krPXey75fMohonCkO
YKd2qv4xm1V6do6J9U2UILDhWpRziCdxXa8Eq32HLIe0S4Z+CqI7cqdtP6Q5zBhPzHC4XDSG5TGC
fItwTu/Pxb9/CYT3Q2anJFODJp+T+Z/PYpjyximv97Dqmehv730hGPHsk4rJoQ7Q2pQq3uxBIbAY
RkbQNG89jhh+tvjtHuq5mM4TyyJHnQRfWVMeKbXkJCjh5w561tyBuDlzK/CsEOJ5V/egaJP6Ffem
eRKHy8bTkYPrjkNaGDHXP88FunpES7dVtOtdoOVRi1F2vIEqwsrdX3l1et7GBup+4yKaZfgviP6u
ef1P4yHeSE/iar5km2OlPRgMxJPWX84JaHLW+aNxDKjqkSL79xvO6DGzJvqVPO2dwL/0G1UbDKV4
3KZTJs3R6cwhpXQY34Zy5BxL0zXxEAHxXR/srbSrTW73KEqiT5KYrN8122j1O8ehBmHVK3bLmzbQ
Ggmk6ejCeLf1TF7zpsPd3XrDT0oCLbBbb2r2VlhLnZlMHwmQuSbRM4oNH+lgPayGsceJ+ou57IV4
7ShmOwSfytGfwSYgTRN5EfC3O4lx2BS6A0+e6KZNhyDkVefntsI3gISUcm/GkZhf9utc1EV6m/XF
85sW55pBeaw/aIFSDqWGvGXL/rFme4HhnO8rajsNtGOKE7tLHFzxHIaEOzalAdX/LJ6m6xys1NQO
63KCpl9+oNTjdEEMp1Sd1VM+ct/Ft8UU12EQAMB3063ro/lT6ctC31uk8V9BsYO1WIolal618h4V
Gzq/6fMN39UHlp8yNYH0o0UgBfCR0u9MCfnAYMB238b6oIP2uZkcUjyINliAbo3r0/z1uRZO5OqA
YtaYc//Jr+6ZEgNw93YvrO877LBNVmqk/oEsS1mrw7LKcaAqtWpiA+xhUAHNdRtWPXK2oSDkrOi/
07BoMME3iqr5EHb4DWr/hEGk9yWpEMrlQUohXIXIAKCvktTvdh4TuWApY6bOcV/ZdeFRPRS3elqJ
L4RFJNkcxk9Y6fvxiPxpfLkdoCW2EI3KCNOau9szgP2gRX4qWvkt5Oz8vw6r/Um4kFtdlHlciSn/
cL/I+vFiKGUBGC8eT1aO7g3v0T27rg0ZOCBOpwlSnei0rGAQ6BwR07oOaCE1+SDLyD+dXjlzf/V5
t8zRUUjSqBhAjYtlANJlSyUErooJ/pp855SwNBc5pHXV1fAkOBVSadmHjXRDXsGYQNjecophq9FH
/X1slnyN/BhAGuZxQ16C8F17zss8oBGgiB0BaWSYt1FIiaVGJbfKYvncSxFGkEPC3piEd32VCQPL
JqM2MyKU7T1OagAynkOrGE/Tx3ZDL8NgMUsfNjXHtAv2AlSMSGrwZMvbp+9w/wAjtf3/uM5fNNJH
Ea6sgxvXQ2yB7MPXNeu7ULl3EJCTqUyqzkuRn6RJeS2Swxx85/V9bM08x4Fi4PMY3UF/0DZhoKmV
4aI16zyMnEtwmBBXLxeHFSRTZjKN1PYm/WYut3ZLj3/j+umJIEc/54fm5eRysS6eFAnA/R1LgGhD
8tlMo8S6CtI1Z7f8weRaOe4ZEpeDMFEO0bAWU6o3huepfwIy3kybkCCE4443LVNfBuxB0msdEoo1
47AKIzrPNYP1ySM5irvRe00rb9+cOtKXdtVgoEx/WntSaB+aq6bulzYFtkoFAOEsGykUNrFnek9n
kf7Rp4ivYIPw1I6VmhMgKj/u4xIlFeIgLO8WwvUu2dJboqwiNAhuRGDBH3sP1ESNuKXlmsWn+ThG
tXjKy5+ot5okWoPpFrZHzy93YzyMIU4BopyI7hLW7A/+0EQnLo8HyQLMop7YBHxhzpKIqgglJNbv
jo8JcGqsTaujl83bfROFnrGTE3vI7ebOuI/0Tv9k6pZFwbwn+N3t4op9Ms0QLPsOIetVD73AQZH/
LmHVUvCBIBIiW3k3WI69X5yaRtVxxcjR/8vlwafIoofRX33DSiPPBPS/QNRo6UPafXVkeAoB8gRN
nqhCA9SvSeGoX6ixFX6DTuksC0tgT3+sETw7wf+tvpRbfHQ8qiY+17phG5puXfqZk1bnWRwclbg0
s5hnWjUp7mfcPjR8EQkEOwyLoFGKtaGPm0BGpQog69DOW7cFX7DZnYDbpdXlrCC8MupOtRx4rbxt
/AUP0HUNH2CT/zMr2Hgqs7ynDZ9oAi4s4tPWbnz71wS+zbwcA2UQm6+3IBtjr/VfWb3FcgK5ik19
9YEIJMTPKLgNnvIouwPesjB+OoMdjkf5E3G9qZ4T58i24J3qMaVydPfh/NMCNeLOo9kzwcbYBQGM
T8tiEW4zvq95ZrFdr1oQEklab6vnKWHzHbQ05Mu6NMirnn4yDKLnGwB2a377RFlwSMRsVTXnCHCy
bzhI2nFvyngevvviM2CpV+pXCd3IgXfNH4UQDmiQNwrEMkb36hxfYM/yVbmTRS3JKSTcJXGiFLfl
Ua4wiHTvxOLWHMhEMZsH0N5i6hKoACbAWKAKsyTDFG4YWQR2Ldz9BHJeSGUjCKBg1nZ4qp5tZo/5
JdwHzHJl2l2uc8dkmYzcyZxCsl2WOO/jFys25uhf8Nq1bosC+QlkGhQm2FFdGgQ8WHk6cJEEB6YO
du6km3DjT1gpxbOX3hhdo0rCMrqDu5ACLA7ME6GvJexlUYd9xoDQGdff1eEFpwsv2Wx4Y9vtRWK4
+kW9Tzz7vjBemTyEmZQyXmNM8MgiQjMwFqlkkyP3rTCExBU0zGhsxMDmvXuw9Tk7ecid0bZgCy+8
WyHrcyYJtbLBAKVQCBg44ZCtMGQdWQQ98VYHpHGVZ5mbZ+qTOJlLQsf2gS6Z0f/DSy7VnlraM7yL
eLY3TGvKErhyptWvrsZGFdLl0jxIdkw0Lcm7DOK2xRGDUE6lomADPdgg+fDYJQbXU0Wy9HytVmOa
RJMhfaVR8fhEyUDFbra6sbt/n5YcYcjFTEzD5fpsznYCB1GrZg8YR6mnTpsQ9+RtWFMVRGC9kv1H
YRWRrkMlQsYsl+QgZAg+Hlwd/E8qA/me713dY4DS9G2z2dVQxzCwuzhsMvmidJoDntTwMa8rpYZO
Ddw5m+2FnLIb
`protect end_protected

