

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YqipQWc4JFBZb16rc2dodhguFDkilKhXXsYOnDVSNRAjtkaR6AZEesZX9P31kdm98GkKMNT69IgM
oU3B8PoxIg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Th08Wi4CTujjzYeFPRrbrk96/H9lqJHT1fOXWDhDkZaqyMx5/LmUZnPHzc9Mi1qiTcgVKZeTpkDd
lm04xNkvaFBlZ5KAxEqjMNmhtMTNyj98wbYe1WGtUEppm4URdSaGhgzD2gvskrJEfU0HoVjNKsYv
Y8g1ek6gYioQSqVo4Vk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3ST6h9XhpdCHj0//nno4AUPlABBr9tQ0cisrrim6ayZf3P6t8TzMqSxgV/q0TD5pBIm//qvgm7Bo
W2S1EUuvf2WqWkW7p/E9CPizeTTEZkAYHckCfZTDk/HTJdolSIFeCHjfZiRizq3RlOIw44CUEMSg
PXhJE4sbT53L+d0eIaNmJBJnZPN29vIw8LbE7t+Y1oivoLSh1BhWy3+lZNV30PrceJFjB3Ylx53O
r9RULlN7k4FVXKoCkEg9NcpjWNJAX4azHw+uuE/ZZmEDfyzXMbaQPIzErM+LylAQ/PYfvIwSeBK1
4Z1Yudv71r62qTHPKAu2JCMEmzvKCe8RAmGoeg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iNgef8JJ0zz53Cg6UsIY3rdr+PhJG3ZSgPvV55cmHG2d6Sfxzk8LG8+nTrPNPEPV7qefhOfs2qwO
LV1XGy8/zcDatxxl7RZSBTwjwXvbpgbJIb3oKBLjSbNQOSIIh7oK15z/NbQ04jpEoFW8I8unz0Dr
X8lH8UO/ss4o3sjSRmY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gdQRq0TszGQ1sYR2djmFoWhyazt+0Tw2kvNbiTEjaM08h64rXWx+KrfH4Ux19p4jnBVjDnfhSE44
xN7ehFd8XzCnm6T9eZgkCDf8dP3IGf2Nl73ZHXLjDsXHqpK6BXZEG/Ko8+LkLz9nw7Snn2cWezi5
seVqFQ9T1Cl73kL7otmtLUuX7sR7LkwbgtAzFivUF8Ml8V/izjdNdzsqpzxjHY9vo/n9JWZSxDHg
dF+BgQSeU0ooY6vwulhfUyi8hYLdbvSFz9Xlr9vUXABI71kCIOeJMQA6BrcWbYjoGqM7KNL6TTGp
K4Gc5G7xM4ucj70Vz377eDl1W3KXvVQRmQSA0w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6928)
`protect data_block
VCg0yA4+NLyg3guwjQZDvLmALZJmwwhDwmgK0DsIm2lFrDWaBcempNaOGzZwMp30BWbgyLFVZkFY
Y8Nup4ZIegeVohHZJZDpDXyLEUCf8tl/9q5uRlo+O0A2jnbF9GCBDxqNTi4P8gTeQeN5kxsJRnp7
beerrRUN+ow7MV63b6YmK0DAHGnrt0ggRQIPkqJoappLYLz6H7cLdK4VCW+bw9X5GpqGOJA/9Kb3
vY2870lHvtpwY9ICNCnEp6MDAPP5hSCaaHxkb7I/kQbRhBYea8o0kGOXG08Kuxe65oOftAjhtluN
MsOuI9be+AGGuQP3c35I31VRJCGKIC3Vde58IQfg10HEc4IbocR0VzWiaoidC6p3HTeKkjWyY6IJ
2XcWAaP7HV/aYLhba00PlAwJ6736kYJ4PJS4uT/jWD0v+aw8Uciw18M/UbsFnAzoZBh2UIFKiGrq
DoxGTjGGzRfxFNtCfG0Ynfo/yGcWHDHf4c3Yj3Tcs0xN+T4iqU5UrfR20MeYCGHbCdgLv1CjQ2tz
BVYib6b81nSl+Je5i83ZD8u+lF51pCToNdzlFEJvRDspXFTw6ae5cQG5k2CIfB/ALjVIXCwH+Jxd
ScO/4OPHkFlMMXA1iAB5fneYBh6D6VLWO8KWkvpv9f5AlF31/wblEq0YT953TV8m1ERq2oZNE+bi
emk9za5voPROmZQ954bTkxiEFS2U2NLHAaskyuBobf2gW3ZhMSof/I+vARsE34AJVTzlBjRIjRt1
4Eacsh2XVacY3DzExaglvAYAFaCaWSfwvt5hLVlg8MHA33WyoSTQmilKFsbqL17aLApMOqLlkG3A
B4zuhaTP8IMdcjRjBLI2EGqTQZfm84Oqees30MmWcTtfj2b9JU7onn4HcjzRB99LXfo+7ur9Gcqf
hbSiN6ZNYxGioc02kVe0WTGoAiMVn9bvhbDFR6iDmvYcYJT0r37SwJdDJmJ36Wem02PYUi46WtvK
DTBbUA8+z3ht4QnsbY2aByzLHq+qdCbJB1T3J3iGzk23XEOp9qs2Q05VAqSu5HU/U/zy9pOSiKWW
6aXeosdJy5pXMSszZfV9UqWuzjWAEeLM7PPujXh8p67LDo4m+YRflQ1CudBMkrr0VZN15s1WAUGt
KoBkxQYscf5oPlDtG1HXFkfGjs3+2Tcx43AMkcQ/bYOuaMHzaHJgIaAP8t9SDgcKgZJJbeQ53eXC
foZyEP/wPgJUPxnbeiOLvnARskXZetubS8e3xcc1cm35tm2yIk5whRO0+rjyQXqiLrY90tSn2hdk
SmlC3C86EE4xkFPzRm+VeAHE8amteQ65TJ51IJaBq3Gnkpjp92VxmiWsHnhId/xrg0br+XLXsQty
0bBE+iBO/F+9OtcJ1cyw5snKAY76Ntv0KsZCZsg8pFact5Hm6l9SI3U1mxzT4cYvTCiz8SnKMAUE
Gfqzp4NTZ9jD4Bzd0bxg4S44CqcuRzBi+h+eAIRPs5ztHSmWD37sclK6+7+8cPYqYa0/VJTsse/E
0ICLYaFLyoGyhTe1CAppAo8EMUNcV14mdrSgJ8IskokQhIx8OqVwy5Y1bPhZ/pt1Jt3RVYMKa6ib
+IJu43pljPC6t82tVz0knxGNThDPQA9n9aHYa4VFw3POIhHONLb3wjZbVTR+wUMm7w94KTGlyIfd
2V+gH8FQTCA8QwHqa3scXc0EAXfZ493vZWVPQf1PKIys27NQeDjUyyIQriPL2F0QtlUWlNgcYfkC
qyE1jm4bOQTvJKpmetYGz9Y7IkMyE2eMC4jeB60tfU1uRasSIbgqKV4TiExDxlVFSg9C5aOgrSnw
CSQuWBEfLs1nEdQZnuwqFemEbdnUzBsjUjS8PGPCUgrzt5VjJyBmECJx3z9KYGgDOhbFm9a1d24j
a6K8Yq6SAJTSEspNqB40lbyTlN/xU7dzneM+IdmEIDDjsDUyt5a8PSxkOZygqscOO3+rt2Aut62V
bggp+BsHvRIH8FgVR71CPY0a05Y3rq16pOOReJJAiF9947DwzmSL2LyR/4MMs6Qf3iB0x5iOYD+O
V9XSzZzMUsAK4WQ31hYVgZFImyZcwV3H/nH6PiIQv+rfxE5K5rS4Mgpew92XF9EqJjLNKXd+e0Xg
CNAC6nWcWyyJ/UhW8LUhHRlwpcPw0enlLN07oEkOTrsGBn2w2lIgfWUPf/88wzSQdS1St0F+EujO
HIErqzYxoA083pM5N2pr9LtaMjckGPwjPwv4lL2qj8hAWt7m8Zv14gvXxXaCjXoL9/3id2LGdRac
sOi+oHDYdSNlBCu1g+E+iNYgUTrrmMl1rKxBCLM1wUmOjsTIV766NJLinS3ujcL7hVfCqdGLvn4O
0hxTcQWd7F1t5GiZhBmFF5CJGttPnaEZ1Tm7Pp7AEZywKTCosmKDjANLWn4lyOLSmWafDR2WSYXJ
yiC34K6bPV8xhMRR+2fwuiFcD69hmSGDMkVYEkeb+Ylj2qJzPlHSpx+ExLDO6Wut0Wh8MJXxXFyE
NlMzPC2d/z3MF/wTlb6FAan3azs28oLiwBqkrCIlLq6C1ZDhSh/slS8FZLq3gYsA9pPPaneFu6Jn
pG/8lHZal0f8lVXlB7l1UnGw2So843Ndm6KBOoVttO4w+xnMFNKnlxwQ2Qz0wTKPmOBJQ8ISC+fy
k4zVlKSDIxEIj3GGyd5IS6X+8KsS6Pt+St8aP2OyHx2mohUXXw448qz58dSPmhfXNWjCyQ/E7ag3
iJptJO7kJunPbx2lDn3hCTCPzmFtW8D0OZKMDgV+o8kLYEkfNkVuEbWHm1fKrtPe6iSM9mt38RuF
gp0JkImjeCLMhF45HYFPUmBw6RM9k+DnkCuJHaj+fjRrunwKokmJy90UV9Nw2fn5kiVVxzeQoJBV
GTUQp769kWiNL3W5EntvBMVs8sCqSsH61g1aOpv4vtrmeepGlW9STxk5xFbJJ74pT5ALIAV4s1Pf
wWf0VVKRYZnx7PC2nEJohRg1+Rt9OHkbZnCh6T6vPIin65Z80WU0vJoggzD9m+wMkcZzmO3xqYor
qhkShMP4WpGHk8Lu3pN07jDfHU1dB0666HvRgZ/E1puI9ozajUL9CJHSCSN25SusEYBAif7iGjFI
EMV1eCxkz3VRc9ecYjCArOTJLVOg5XUi/7S1Y99G0q+AxUM/Z4lnQaACMCprwWKyFa7kKM99x4VB
KaAt/kgjHzko2T7ds2xY0EuiC2D7E/+fHmi5LFjBXVADycvZUNNUNhh9NJOFT+AZpJyaDZVWFldL
sqqXOh5KXrUHAiFpPjjhYZFC4oCZxoWKt20LYznm9UFzMlikvxIFmyv/uyAM4PepT6//NDB5YA6a
iJE2XtMSFL88qhPgGeF+8Cv9fnKXGhsZkuGooj1nQ49jMRNdDRgaLnSSpkXe66RYt472BiGnoi51
iTcDBFNc7OXvvY7lxKDUPSPHNTBDSyMJrR4SzfoiazQOiAL7OQBWHEPm3tzYsxaF8mjEyzjWQ0Ge
Eb3xblLhP+maFkI8NpPs+lDvydSR8n1uxcZLX0CtPpIaszrakC9KUHOj1HRKXMkTtj4R4HAHtSV4
3ymtkHRFAk8VBvJJ4K32uADGB5O/kNK11+bk1UGEIrdLPs4ivhSBAUQW25hA9WGcXStgBccXBzTm
swg1O0dZhtS1+YsovSh3mqzNUk0TCE5Oka2Kwtvrn2YDfRx/qQN7EqhQTNuyDQiLo35zdC4XFFQt
rlFpDfW5PxDdTwNaX5uF2Dg3u7BoSz43HEyCMMyBDYAaEXLBNZQPZftZu8giGkDdeJMRlRx7KzSL
qVR9S1cGXgclUug80t+KG0tzDPLVCQLFbgqcvCcYGja68vjvQ4cDIfWxyqhlUq/iI3bR8Ljr6pxP
VegOqzn3+D3tzMDZ9f4FXWBeCk/z26sw7bKrLztt8tamHl8MafQRztBpDkHwYXsef1zUzXG9r+Io
tdZ/Ca1+IBrvEPcrvteeeXuSdsy/2zSMFUrW9I0872IbUDzAw60X8CiLQa40fAeBGbJ6/zra8JyA
3ksNRBAipYs+YhkAJblbG+KmsR3FEtFbQxHX33JeWghblB9fCn4EeFaOv8LIswXmK/2mH4zBGdYJ
cwLR1WgQm4ElIKLWKv7H4lebiMQIqJ1GsDSUfdYGWyRlnPLLmDY86/QZNUxy46ZuJRMcbkzubJe0
BEUKEmMzlvQCAacaRb3KCEPC5IcsVWpIy22YilTyfs6MoSC7pO8a+odUg8t+iKE0CsR7nPSl9kkd
xlXDzh13Cu/+DFanTpoOrRAK71WXYlOcOc4CFnyNOvTbCBvBdukUQq9XrrQYNlFG1dj8ji4UCJkW
CzJ2pPaa+hMbw1wAbthIQ2QZGG2qjdaKxXfHnu4yHVWkIZvw75VJx79kbM18UVp5QjVtNNy4SD1V
BV7VWk+L2TwaDMG7Im648SamPC4mOaNWLJZsH0wXM6wcewmzd1hbL6sEipH8HtvYIqskCNXNANxY
2fi7MNDxt++QCRxFHTvbkeD/7nfSbmzoBt6iBUs00jRpldlpaS4flMFz5BAf5w5Hzb3f1HvCIsPi
vGx3Wxa3XjgsNfa3gB3yZW6kQiQCivsWfe/soKyB6Q6o9zpQPv03ceCkPl6iPA/y826DBEciC0DE
UeRZ5TkbV/vi4ArqX3v9jpPY94JFBYNIEaUog7hvEKMtsITbktW+uAJsANQQQhTEd++ngoq7tumL
KUbft+g/7nMoHDQwWXN5qpvPcQJP0QfvndposzERQHkVeYx1+Cot9lYVdJ1R1GcgpfIRQn5SiJxU
84pMfzuL6xSsYY63yiwnOfjVJ/RvnFWZgf7aCG130RyouwuZP/e6LPphkhrQlwdbXUYS0/cmE+aU
h21whBcyz+7E8UEeBxv0WVStcSH1Bc5MpFyIpHe+FGvL69msqCeb6Tgks5HYy/cyGzu9LKqcxpAq
HS4Meg9p+i5rPTmRJu74RAw4FG9eSwzjEWO5fIG/U8ooM4jwV83ohBVI2S9VDN/1VRYGcPdmIxrW
bEgS7UWL/Alulj4c26RtTt4j05BlS9vFlpHGHPZLAnUjnIFnzq5f+EB2uAlcJ1Jom/HqHm/w0yi8
7dw50f4yMl6g62zI1CIkUXalWV4OXJkcnYpBcX712pzhU6n7zVS0hP2GyZ5wmWhNwSo5shn/xedK
YTtxDmw6cuYCcaf2LfITvlvn6HHSsHOFS0cgwbW1AlPvhlG+4z/1gcSH1Sdw03A1erNO9pyTRnUo
otnCUeS1oqSN+YW2YMf8YMVM/vs6ER2/nSqAouSYwLXqLZ2UHKigdR4ZvFB89XLCwN1VA8191Vqd
hwBBdgTefinDGFHqXdlBwqHQRXgtEyrt1iOG/g/Iwjg4UonWJZuMYUFEzfCfbNMo4vVGgyNn4h1q
D2jPT1VSmVNw21F8l2makDES8/GeipX1ainFmkmZFZfgPVURiwAS+ZalxdxtPLFt+FxfOWApIF0t
QItyVmEdGXUsWH17pirfd+U+k2r3TfQ8SAmFYuD6CBnQd96XqpJpAa8Hrd2xUVmcT7ntuWerKanW
PdwGU8UnV7dHEpKEdY4puEVB/XZB4gsNBG94sQocP+wMyVzzJTGhq/1CSyH5Te9UBVHvkSsnWOOI
/RKvd/IsOJa2OYfudzmZ+Y58a6bLuLf064T/nFJyVbXC+YBllaUR7F8o2JzRYrTbybkIpHB81z1V
XXXhZURfGng8B7pVdZyZdNoWMjtdECQBtQtnr0dhLzQ+C1MbF+OuLNFT37BgAFH7LJ6bsVdqEp8b
7EplG4lj/r44BAh0Zw9YOZB0b1nxyB37LLZ6d9X4Q46lXAT+A2J6h3gZxrye+/YW7C3HD7wSSZXJ
w10XFZ1UfLTVyYzUOuKHqDizK+3NTPhI/Bfd79/xNDL0HUZXIWmi9DZ3wX036qiKrvRD+7B6LHU2
9CQrvowtB2mb5fLGOgkXNF0Lw7ZMaDKgxGURwkyhuRDOftQBVRXNzMcLgvfX5MkpjT0SpIC6cOjZ
slj0/FuLqYRmvnxnnIn4lRqRg/t20P9qtQQ8xh8VgYb4hTJpnUJJhS1+Wg8ZRC3oRYQ5Bpe+TCKJ
Hd4At/PVpBUch4rldxAmhtXZJl3A11uATxpitK2Ol4MP9bkgYgX7EYRus0VyCq33k+JGDI3q7Cf3
etC3Qy4k+FyO8pH+FU+pE7CUEyzZ7hANPHyxHT3v1lhcQxHuN4VhSh3c7HSrQf7METfwpTjoe4Ue
9L0O34Czvb2vwvuAVZyiL6MPXt6DBCGjqwMHPkS0/yurOx26akh8Ma7mNTtwzg7r8gr55CNS6TsU
Tlncjp5yRjNDUoZv7zFjc9tEcw+N/xLp3kXhrePGUZvmC1iu63KvpCi29KOOoQ/SEWp1N9zFY+43
zbvjL7hDBOWQM/GHLknwo/3zEshNZvXwMUi3oRIy57OBSnfq6CzJQeHXrWOoG/32Iz2mIVVgIbrM
ZA/q60Ly4iPBlMyCLz4VjuMtal0ON//xCEAkFT4XOfznIgi6RjIwR+oBNg0zlX/7KfOL1Enl2/pa
acTZmepoIZ9xDjnTne3UTiDVHx01BQi8PUbko18Y4F1wQZPVur5vvxLRg1DmoJmbB1Q73xbItp1Z
WhlanGENGMBJPgPuPBh3jDpWlqEjEFE6Kf+TZHx6Xi49g/qleLkaajK0264NIfAHa33O+EWhiBf+
9mxskKAb7iLBuMQWg+x+Jfs9A3/bcRR5Z94sdTuS/v7l/JJOBE8I94Y9MiXgUES25CrMW7wZmOfe
XWtlIEc//NowiaEquldV117R3Sk+9iP+JxlZFkTHVC1a34czvg+4N/RPlLGAxPlqv0vSgRBlAcpM
SnXttniSwJJ+Htc7oQ1v6eCmwEo29m+xs7RT6jivCH/FOyuBba4CEMANLfXlB7lgfqNstSuiXulP
W6uxDPqQvOEKutsYi96UTaJ1vol6BPa7O7M+SPOJX48zPkEAd7vTO5m5pF4JJx0ao0bGYrdSjL2b
00yZlFN6bNNI8epKrb6QLFxyxwfHSZ15MiXcUuvCrFsaxIoDMTamk+0WnDm3+7rpBPwUqjWlb1Vx
aAI2JcZ09YxEXErQPPckPZVypp3LwYOzh6G4lIHf2NncUrpbgVwonul+7LpZcO4fb19oHEl6hYL/
g58jvnLoWu5MBNcSSrjXokqpO014EeP6Fj8LrmNrY91Be16Z4TqflVeo+65rqIRZ3MpgOzbjkn+h
TngUrLD7/PujPpIXHNfM04d+VwUHCu6kwrhxoSLV5AvEPe0+goTQWa8hddEEnM0VAH4U7ger686t
jvJh+kwvmqVWW5cppFo+nY8gdPlm5dIrNk161vA8ra1kTiutOeHktv2QAF21bCiK9GLcbnur/a9k
KDv+4vb5DQlue4KZZv/tX/c7ev5gBa2Upj4PODnuU+p7D3OPl5RPWA8nIv8TU1ibVM9h/9yXgFSJ
CyaCP4tCraCA8wHx4eQz61rG5Ny1s4VQMhPg317vA17H9i5Ucsvw4blZUnz8WdvWCJsVYOuZ/qPS
pCi6AeFJNAjwGP68iTRqV8ZGvgzHCbo0r304alNX4f4ZWGU2Xgq7wrlfEX+AIiIkqHpBKofEM3dE
lUeOpMOWiIYbOUlYjclcw+FIy5Y2gFgpsfltSDaw7JGX40RxK2/0kilb8H3OdApCeO7GfUr/fMdL
Huab1n0gLPLFD6Fi18FNo6rdcgf5E7vba2IiSDyRiTzffde3PQAtiYy69juDjux/abezlgnOeJkC
Wm2gQC/3IloTMN8+ef0XzhZCizWxNmAp8UTF+rvh0UJbDwVWaI+4yyt6p1G/OYbXr9YXXNpQ72nW
uVUDge6bPVtgbOJZ0tnNCCi721ljEe4JRs9hZVgpMAMaO2b95CZfwgSptkFXSBeksZx//0+8XFrz
gSJjmOLSZ4CW09UWmuxPVxGW/qv2dh2Spqrs7LHjB6jLXLX5XwaXik1xALya4FguzXnBT6toCMDI
CzWB979iNvqdBa+mkv4CMZDTAvWNWdZ+ixEork7Wl3R7OQhHkLDQWqrSOIGOgGqxU95zBTGgvDLV
4ejBzPzI7QunF+oqjT7GhkYupdmdiNTTEIbQgLWrdPp7O4fiD46vcd3PpemruTLIqr29fEFM7D80
4O6y8pFQCORBLYzC9aoZ72k0KPG53Rm68l4Ph5TUIFHvIDTFbBwN9Syb+5Khc89Dr6Vem8TXgUmf
tS57gRmfL0EL84yEcTq+rmVI0x8NGYLH9WjPa1PoMaJpXZyMUoELgdxij4bXmtF26eDFxkUjAZy2
iMaOeV4e7xQz6A3L4jFLVbZgCvZ/PVtWASfpR2/nR/8tAvud6bMoHNYGhyazIjiF6iAbBE1Ad2Xs
6mpBXPNlktj8tpfqFvbPDzc/gvQ/bJPiCxTdtlDLqAarHatmpOvGLliTXZooeLR8M6GrtgbTc94W
NZ83T6h+bIof6ojJzIqxh/IwCaozQE5e+Z3upqp5zNh790xcNsQ/XnMPReE312ABYtuhFX5VzFgI
tcx7dA1ifffwAG6fOlm0Hk/Lqsdwr+c1IYZ0Blo1UscWnfJ5CZj1HE05pv9UywRLFy2Nq84yE3zU
KPAx8Z6J34KW7DXbx6cfdnUvREg9le5f/tcVSmaR1ksxKlD57PL1jdZrauj+tb6oU+KdFB580Ui6
od5huZNCFlGpkzptiAOJaaXfUSyghJ6GmvYVboLczqIrkQV4fnsWs8TQP/MydP/uIwA2cqEv8ocB
B6wiDlptNbrkLK1DIWseTkr/oNvuXzmo9EbUqR8wJfeD/momctNfMVufdHNy1Xh7vMvjwS870yX9
FuMYiCiat3DBl0smxDzQ+qPX5hpgRFx/DUGtn5DK8E/UdL3JUpynniEFocY2X+flMq1AEQE1QoUi
EEuMrKNtj+VHxrVQtoMLHWuLZOFHMpb3wTeKgA092NJ4CYFoLqUKBxtoYnVXG+qTjnXHQdclW8Hz
DBR2krzS6mBYbgMVYzczv1M/OtsTQvSNdN0ZIEdJpj+5ZSZBStPmuBs6SrCoRPixPKnlGa0+edYr
P+NGLZuBXDgrMJX4vpyx5z+WXVLrOOnsuGeOBG9xQIEw5ZYMSeIn5sWjq1tLDusfTxB0L+j1VVP0
KIoT7iqbkccry6oUITfIDtpqdWtj2KpWzp7nB3AU7mf5MRW2wlzJhoA0q+AS0+cPpJsr/3/uJy30
lDjYrRsA13htsHQw6ZZ3XbblBiLeA/Zgqi8PNfVz2g==
`protect end_protected

