

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pTeL3lbzyXpg3zBlG8xXBsi5mPcSaOx7zOxONTRBSW321/dGdDH2TpaC43BqFdYZqpUNj4ng67vZ
qArBG995Sg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I0+MKhxg9FScVNavGFQn2xkzaE4/JyCe16C1b5v3ObJwo9nXDzI72pLgwgIfWMASSmFXtaAAw0ml
3uLnAPMYr1dgB/uJGeAtmT326qa5BMsAV4vQ1Yunxch6eAaFBVMMeEWawv99YiJK9jkH7yDAOpb6
smI54SxBdohXuGVE7bs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bDMpPv/P03hJ26zOMeRntjG40FHNolyY3dG2sIAWSb+A/C9vMJYUZduiM8NsMGgn92oqltQI8itf
kfh0mxfLeub+eu7+DutH/IonvZFuvU5PDOu5gXDe5IZcX7PKYSeWlg23QrTg/K5l+bblhZE0trh8
gSCxX9Y5M/tKkk3Ah7QmsxFm+D2iD3pm82WCrtLPh7JqPCGwGw7ZkIH+rqgZe/fQHahkffxj0VdF
wp7Pe3wFKtUoiMTg7uNHWsoKi6g7a0GVmS4unE3L9HQtqDdu8p186XHZQqxkv2iNX9KutOONjQNy
x1JPQknSlGZ+dd8WmzTlL9rwhQHGdMhFcdrMGQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CqlfcKpSPaBiicqGT47t9PnrRSQ8njMbqaZWYqvnT67KXQ7fxmLQJl9EXGvFoMEq5tU8J3rLbBm4
9pWLf80+KgxXgS9WPEn1zRTKt1wiye9VOUHfewp3QYM+B5lPR0EENtCdssVC8DxPUBy9Aythtbty
2YxNBkGFMjMRSnj+A14=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jiVIVHHI1er6oSZsM5uji5FpVlbZFUX1C20PfTXKPYBzpAjDWZhROWc8xFgszwvy5guzSmUMWOgw
XoJ7z9N2ElsO0s1NH9ojznzy4rNB66tyJa27TZfjI9UYZ/9rfTzXHnlr6WpUX3IChRrS6x5LI1mY
orERQz81jyLKT8cB3O8KkjO3g1Ks65ZIeY+E+7T5cJHzOHJQcoiTTtwLajrQktJS0RpyUJr3VZHu
CSADq9QNuiNkf73BoFHvperz6rZhWbdV5MnpWKfmllMNlSqFwzZuWbMdZs7ZNbssXYmUZlJVjM52
JpTXdo1N5lXyKjXVvDlv7kCHkBmnfQZM3rMXlw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17184)
`protect data_block
N4YoebCEFqSFp8iBXjEkaH9E8F9PHdAmC5xt2PhL9VDb5y7yr5l1LAfVD5gLOaePswXESJdTEMhC
79yfFIrBFVILT76lB61h2nhBdzCB4+QG883HVIugC9UnfdxRJWPVLKCUS6lx1zwuO6VbtZGyqW7l
/XPmmbFiupP3fC66eoF3SBqPS1aUP8ByuoUvPqXBWBHf+Vl/02v9Pi1HDppxeqJkAxDGD8aBB3/B
sjv8WpgnpaDTJ7FEZb4w1pR5uazcEZhpOw4FFX/u2SXA3FoVXdEEWsC6tTBubw1Hbc9RDk1Z/lb7
ShejICHal5Cc+TSVsHwsURV1vMeBBHHXjhQupIIe7GUXz0xKxZBynCFg7eJzLnUrX0OBGHG+v9Cw
asUl9uveS94XRW5u53h2W1fx7ef7fbLWnc+ftRe1KAbRmLWRFDj7fOTInTXcvvkZuE1z0tkIZvB/
D2hevKxRPUW5kaoG00B4G7V6HV6haz+M1n4KHSLLI9VMR/RN3KCtPaNNLLzT/yxsJVqkZRBu3exD
Ef7iOE/7bKg+qIp/sgkEQqJ4T36MK9Jn5bF8hgEdvvvKhQ8t6H62mNmg/8cufvWiV5AVGI043zsb
YX2CZ9cAV902JsCFvUulZMR+eaiicBwXmGRQpgA5rq7b+r2zowiYYVhiXSUKBsiffVK55VDGYrlX
5sI0PKMEwQa6V5SLY8BTk4Q4FMd3qF4CHChLx3olhbG38jjLIXkNT9xNsKZdjryEkMhzLmS4EgwM
gBqP//OQngmoxuHBSAXEJIKXEfwsM1I+RniP0I4gkTQnw0a+21dUxYF/ujSyF7soW9I3NUz3UiqV
zJB+cCtXUv9H3woAs4FoEkTZ5eotUjt1XuAT0IBBxxCBBGXDqZ8ghu6XzKmhWLI5VvDySFDSdIgn
ZDbRBirkcuYDSW+Wv0XJmqnevvTMPmaYVYwucZs65QI6jVsGZsKGSn+DhFsyctvnpxGrm4uxcMC8
4dzNz37p2HZScsSCDdcL1rhMivVCSOIoTbFtboT8Ppanw3/dYsiehO1F950zOXwY054NrbLOWScQ
gvgp3k6YkNjAySnVQIVcyy/QRr8HrzRbDUWodWCx+Y+2Z5d8vRUAUeMr4LuM6W72BCWmPFC9cLdS
YYvaK89kMEdBmf/lfqVmUJ4NCLB2mYy6M6ryieT2LWYn2aJzGC14YYejRmKidzbFUnCmWcL0vKON
pNbfLNHj51hgCDVX2g235MgUxorqfjX3qDFNJn1R7J/hfCD6wXe5Hk62QbYH53BvByyja6G8RkK9
uQ9WZBcJ1ZKSofI8btfPbnAOswOpmPgo8MO+lM8G8gTojE6xyUXxLsnJADSoLAUlIT5I5z1jztPh
STXU6FTitO5QEY1UaOpQ0Vnt7onFG+kujQ14soDn5fF7EmBQJJ3bBccQQ2vzHrBdxlv3zbCvtLs2
VDZ5UzQM6ZgUVey0D+qJ0bsCp2B6r0jXbjLZq9YBdYvKybGErBAhBCs9zfZO1Aiv24SYj5bTGXgn
huQ+4iWyPEoRQ9Ut030l+d8r0TmxjdMB4DJd8aB+Hcx2RWXk+fJJWW+6Xk499bOqSC7ck9wM0Vo4
9SO1kLe5mmvTLW+7b20LTMmoQggw1rsM3kwcb22TvqgM9FY+Mq8W559vbkTdxXQ/wi57+hLpCGvp
o+lx8OsefhY/UZas1O6i4ZskAgYRGR2/KKyOJfgCCbx6Y6odC1qAkAg8O6snhxHaFXz3tTWp033w
ngXbRMcoD+ASQqhHlqNkhQKZm7JKyuHT17mKwKmCK+XYLKM4LUWvqzQk3sjSmGOIKd1HxODbZnIl
c1oJcJa09/jweYhWUSl9Yqso3QnkbAxGuhLw0brMAdA2W30bRZ1ai0w1L3apiyOr8H2ydUjCYYqn
T7ayoF3s/3V1pn58Ig7Yn8tT+F1RCMJBRQ2AlKtpfurU8q9pJ4AIwTwNsEdrMXLpvXoFzTkmOd5x
XIbRDg7rItETbbWVoqXqWWnlppL1StVUqKKHEAvleoIx9qo6gKcVOmyuSkdQvbANawU2Pa+cxaMk
qtZcXJFtEgEvxkY9iusBaytWjGVKZot6UykQKbzwJ5rliY89mKQLlj/d8palviTyTrxPfEeupNWb
Iq054Fw4Vv4u2IoXEb3L8Dm13l0A07VW7Gip9S5SNufGype/wLlb9kKXOGuKHS+yP2WE4LwygW/B
myjT6jRy1OMDddPUbx9Oqfq43N2ZnyEVVvGUTy6y7OeEOtiwgOuTj3Xg4k02byOEUlffyNFu0aTU
CdxBAW8Pvs8A/Liw4eoL1IoU98EIQpKOSpX3ZRWnpXC0t3W1EYpdumIeuiNBrSR25OTlKc+ZVRZB
7k+Urr8+7A6PXX4GQy5Datp1wK+zGSX2le6Db0b5YRmFJUTtWFKkL7FG7T+NzXq0YuI3zEnDcqn4
uU6TyxhlxU1sTAj7wxW/Dp1+SO1zC9QHNYxkW+LaPsGkBDWJcJ3jq8knild8BcDXJwVpHQS/rhgn
s47WZtC3Cf2JlSsAH3szFqc0spKAXUDz7+MjoR9haJajY7ygBj2tm1qFV/Rz02EgDewXZ5YkVdA2
OuQYIfyd7kbE50JdLq7aTgA6tpvc/vU/3uYCGzE1awQiQqVzClM7o8RF3CB/31l8BjxDNNOsmoyF
p5+HUFYQBTiQOdcgGRG4UNB/XKaFx8e6vSBrViq0hXsDG6lQWZ8doaWv3wShbHT9S+Vd/mFxKOBM
cEwj5FzW98ysmFb9CuZ7PSFAlicJP9qS/fIgzVbrGtmSsCEOqOz6ndj9Vqw8utMTLhXl/uB7QKvu
UaDLabGVsg3oaYgawAjkuOYXXti1eKJGiMj6Pu3rQS5toGl6yMlG3J3aSBXIBOO3tw/iXRADqxi5
G0PX525I8BhXfDKs9dhGrXiGyzaqjMJ4JiLzFXHY9vajhvr9I4IaaMZ019s8wwwO1MhHs3Arlm1w
kNrDsQCnumUj308MO08E0yhgVvpIOKBs1JeFAVb1Rm3q1aHcfNO4KWnyEsjdI7bGCk2qWticpYQf
mdjiu6G8mbR7qOwHiHroEYSR2H8i9I3CCCeP0/Es6uVj6ObEfTD6QWu7Lofu6NXI4MLcwTS4O6no
tV62I0mIf9czH5P9eojELXQ/glKUBdbeFhXkFM3pkWrEUsDkeIn8oWXsTrDui/6+6VIzc4s50zf0
yy4YZjFCwxMhO8uMS/plpajGM9/SA5y1rsEsAJBh/2vbKVktKBPOOc++nYaPa+6aucSyZxgIuEyU
joCLUY7AN+uHo09youJsiOibxgbvr1Cv6o2hC5rf0By76aabqB/f4Wa0xqXzb4r+tG+0xeE20K6K
pvLS3gIjYv1bjrckCqClwbEOjhLR3c9mH066xDeSoSRRSKyNxoYdmbgruMAaIjMjunRAVNt5uyVH
vGzYMYyOSgqaUMddFvY+TP45LYhXahiKRacnbnR3wEfNlDItmeFMVP5hyr8X1GKnuVASo0LlzPh6
rS3b6AmipZgxKo4dhqTuWatV85AYXEYYO3mCQ+Bg5GVbNB6N2pKv1aQeZOwrHlObfJ7NXecnSp2t
1dezbefhbgYPTKnqEm1gBPILx3RTSui7d6M55THXN70DdHTplZTISSC/wDtnbzv0P/zHc88BPWR2
kTX+ChFFAcTW2jP4HFKSYTZdBWq7aXbZ5qqTIGI7uYAAwpc1uvUKN39aOGB1yhFSTaW4SD6+6JnS
jG3VlOTVRHAhgBd1LnlBsTlRKcV0Hco7YMNC/gshCBoE8jnPtInF0+kM2L2/81OdlSj2XYkeSG+D
cF7WkNUQkFuBXEaBPenhK8amkd2MfsZvff0OZMvClmb60+VTjrIIS0osb4ebyexEHHxXzHa4bcNu
d4PPxwnqI691ysItrQjbkolaTsUZrLKK1mOmerADhu0oSnKPltkd7sCfD6ot891Fout+KPI3/e8R
OBGnnbV/Glt31KqfIKMy4j/vHq6HeaY2fj+XeziR7RMeaeNf4cUDSKH2qsUExAJil6IRmvmltAP/
SBCc2FFj6eMtvmSG2mdom1nl4qk6ui7v81GSNhDtuLSYaAItiwX6DHHTejgMv2QpyelPS7yg9ttL
wV6KBbGc9NFJNtGJlpgFT0aVaLiRRq8PbSnAONs06EBGoi2Ds2IGzYi2okAuL0kRAbh/uvyiQoIc
wbUsIwuGCdX51kvHH+tLG691a83RO/mWUakzL+CMXwUvZCibcjudiDHRsBUI/plTg+HPvz+n/V1A
1JFfnCvPinWEfqTpOCr/ECDIGzGJ1LZeDtaqfrv40+KezOlUPmjErM6IGV8bRm0lsYNOGH42T3oY
FbOGwUHgYfxo/+Q7gYux66RtEHl4hz5DwZWe9fg1Kd/cnI5pE4w64/1aLc/yyfwPbKMTdFfuYlOv
H3CUww1IVzarZaG2KRPGNPLNMdM0lBZILQ7CmbeipXUqIUJHGe2uqwgQol3U1n7NwR3+uxOruA1G
j6PdYZ3MxBaUIlqhZhJO+1IA9neJAStfUnWpZrkpgwRxVLRdpz9pQPn8svMcxpvnLDW9iF9yyL/c
FatmhjD5KI3Vs/inR54iuhNTdXwa1LM/KtPfSlU7jH89nRXMwnsPY6Nz7IG0RwbiQvSF0DSTwU2w
PGvVbHr8l+AjtVmiqMK3gX9oAZZQdt8ap43w/Z0PyLnHL8kgvq+7dBP6Rwadc7un0nvO41r0AjOW
nd0linx7/BUq75Gcuo6LIdXH5+14Tc+G8mRlvEeXiQT1gV2aXp9wZj9icj3dw95Jons0DwDTh60d
fmyqg9kZBpFA3uJCmjawPhrAv3xrojIhvCWKbeB34mA6SQmRwDn6WiqjqityjTaQCMLuJRTWR58a
iJtSDSAQAmZXsHVHeHgxx+8U6ySc0QsuFPBNEurhxsT6H6/00r065xsnutKmpTuJ34YBAuRzLG2x
ws0DIF5bv1tAFYeQCoKp5b+8leqWxVGxucF9j4qTkozp4y645pHM375jRn8F+y3MdZFmESzzD7zr
8gEexubuVeUnhrU5YDgkQ1QBBYVm/ZFGfE3xofaYR3g3Pe1IW5j7k2xrYs7gNzTqftO6f7PHX2BL
1RfXi6V9A4aEFlQRuS+l9X28wqG0KLazZwG8/It4izeKobwVeU+4eau6CDvcaNC+jiwTeZ6npxgm
i3GxAIkeAPynDNmTvBZPrSum0ShXv3DMTd1LjwPBltG/i5mBCaauA9EfEBG4IidETKwCVJ1PCsBa
9SghMCO/kkslqY2iCkRENuDEpJZj4qpRjdudUn0RPVNyN2SloRlnS2hkVegF4R1qxWLQKcuaCGRK
4grNeMFdqAUYlnsUfkxg7LzZm6A2pAahYMu6hcKjyFZLDd+B8kP+h01Q4xmjpxpggYrVRia/xjJY
ffCjQ250V9644knJnsyr4nPWvYPRM+CR5kVN8RocFHRLTXhgzEoGHsBZf8up3Nicj8hgZ023UcYY
gc5nwPoYYOkplCmkPlq4hKTH8JCVsftRdi9bOa8F70gqxIWJ3VKrDjqZFL5UuCEd5/2Vi8SQFeJv
veXDnnJwlsybX4wLkZYDtUW4b8VMJNU/PlzFlAiYdXuJFwCRni4GJfFZKjmPRp6XVUdzEFC6OWu4
0LPmD6UUETCJBuN+IEI1Yd8Rp2wHkYCrg/maqfaevqDjwhcB03OM6zuqFCDAHkMY12h/wTrAqSLk
cl5IEICjvmNfV+5/i459lxwRnVcw83dntqxWC8LztrowzzsxCZXvF7comiqE3uuKOWEyVbKQ0nWE
YOjJvp4DI8dWlIpVo0zqJ5N38r9hBMxuhGHG6HNeeH1/lAm+AMKlrZ+Snns92B0izhFiPqtl9T4X
95c4Qvjg0K9tMITXa/acA8nMYnPhFegl4xhvo1fTAS6HdVwgQC6yzkBTyqTaaczfBcZ9Np8ef5gA
6swWlMHaId4S/F3IvCKSHm64504Un2ldyQsbps4pMdwljQ+WlhPe2Z0mQyeJ4VK75NutRO7TtB+d
p6ubkzR1tsjIFdX3qMUr/jxlHAzY3euw6ljUxfUOympa3YYKZkGLJU+Af2HQBBXoqxjTCR3h6VLy
BloXopHDSJtCLR0lZQ+rWl+vSIuC46IZXwU1oaZhw5LsfXeGYoDXG7qx/ejgcg2bXTbxXU26STHQ
P/XtW53LXT56YJ6y0ZCwrYCv5zlQKkd7T1ro4a8RdjRcKV0Ui2syeKgPXzu2Je8T++v+PQX9juzS
I2UAE9Uw3FFm7t8vXNHmard5V+zY3/+mKkx5iJ8P3gH+IvBdw+uyBgSk0GBePQUcBYBosE/9I/xh
Cey5OpAUBHTDDvR2aPtpwRckrqU5bQebvybse43BX+iaj2yRFQNA9XImNtW9cnqcb25LJz80bOoJ
ZjxmgJFa0mbktSI01/VImahWPB23u1ZAHUedKA04r/2BJXdf72OT2EXAjR404z77fbgCyQRZUEDV
uCMNcoUASK3153OWipz4CTyl1LBYtEW+Tf5oAwHzItSP9WolAJu6/Pz7kzb71mMNCkBDi/GnxocK
fwGeiYgThGYeRECsQVlA3w4dQLGQD3YQZjiTYJNEwICCrBUxuDw6ZZNJtUWVjslftY62fSVn7QxH
UV6alM9qTXtzrGHCkwvz1D6G3ZmHPBsgGBDFdc0GpBBx0f007uNzb+Q3l0P1xX59pMZtMsjuzcr5
rlbLxk3Wcd3CRnC+zvY7N0O1RFbqskOx27kyzumzjvA3oYC9OulmAQ7q6WFN8qkOZDyV9kQm6VtI
eX/uZyRiyLmoGclJ91jvuObTlGIJsoVtWY1BJZEW1F0lOLHNe1FTSLk7xTCMs3sIVJVPEPvBDGBR
hKsbKoibOjkd6v+AnXWkhC/hEX0BMyysEBGR/gicz9yBTxQlrSchg77E/foFGLuhVf8SHGDzq4tN
xayHiuD65Hz1gm92LBFXMkIEVMzmBCKf5nUNRCn3zqvpr8PZKQ49d4dPcIh27F7cpZQlHpbAOy/e
JZVz0KmMdzBHawhPCyFYegecRExWBjO5ZxBF8gMk4nFquYMhYBx7coxSkMhF3KDL+OKA30ef9b8j
fwZz/O7SyJXq6MLvFLesiwBOfG+J19HjUkg++MJAtALZUPH9GCe+ww7p+TZDwlTvgPwuZyCcs83R
N37ZdeYR37iN563TtwMr+T7skNvBjgPQeqjDrrtycyUK0xrZeNGGpirpCImF5qv9Jrnak3s/jaPk
GWjoh10Koe4XalCN10XWxkAjWoHEeMoGfkOXqcjJueCNzNpnN1pfAQUL4UQieDBWT4kDPQT0o81H
zVrawqDuDo/UaQLeGCm59lmRPnz8YMFMD4wVHS+ZFQdZAhJC+STNX6rnxPChqBCXJsfiqul7BcDV
ujjJGv82SFFJmi7ncuPgOTwJY7zKY3BioJf8/9kJwf9lP5jiWtlhzrlap55bfmlEHfpLi0wWuXln
+csbkrzz5JDwZZZFWNTSGhMVY0fcCXu/GqKC23XquFgqJQkFj2KPv1mAudEG9Ia5Aab/tyxKrau6
NVdhxB8KjsifP8pCfMUesp2bk+tv01qkYt0+d+w9zzpE49vdnuPMb6nIrw2SfsQu+l7lgqTQLFCB
19T4YqIxiXtumIgW18Wbjg1p2CX041jDNBvlgtPHjl2nssYHVWhyux50BwYEhXeUukGT0eWk9hxp
GUwPeRsZIxlnLhr3Ud/vnxvofDEhfCsJNxj33C0LgTOVyQczmop5DbGsYjQhE6/PEa1oAxz3YMrk
+p8VQ6ovDjx6U4AvGMwLYOKexnxm0+BP7W55Tsj1PF+WYCCngwaMQpldP4/WLqBPFp/Q6pessWzZ
5w+lsjkUdT0srZB/vOGJAjGRG+yPO07M0AdZr2kHn6tP3XVAotlhwYg9ZA/J7Q/90uGIKiN+6aaR
8DYD15aW523RsZ1Wwr9qF1fB8a0z5Rgs4TkZW8L/DM/evgljosLgLuy2eaz8aPghiH/UIKxEVnj2
zNaVx6dj3wsJ+KkpTo4Q4qvtrgp2YUJ4pOdQOGy83ckG4CPi75Brr3WLYlIOhaDzJXMKTRx4CvIR
EhizngA+K6e7QoU21MjY3olphJbXgoghHXoTwjDM5h/5q0k29jfuq267RtJGYyTGlgNxkmCAb9zd
rl6Ae0GNXZbRIBmyVXRHpNcFNEm9mesDffP0TZZ4xjWvHSwV9WuJqWWRg/V1tmOj2G6Kxn0yM3HN
2zBlhyLVfLpsLmkMGanyz4C/Id8wYgXJth8xVlFw+cU46bDQgdJu6qXe9dOnOXAra1FzWTS+b5eL
AYkM5n2VnWFCQc7O3C6ZlB1ZV7mjrZDUwNNtOt/O/xYqiqb046QJzsZAmaNLCT7F9DZe5mOQcqzj
klB7wxnWXmSB0mzOeHBB9T5Sd+s4eXDuvCcwQwEJr+9usYdiWZZke5OZuSkHa2PyHyWffjeBwEJY
RPd1iX6mhNHX3BI5QI42Fj2wTZ6YJh60oPE0xm56FDDUmrKXkjSG+9WdDcvbRhINaA7Lvflbk9+J
8D53w1n4nbQQrT5VMqyXZXShcBvYCK9k9ClwbJcjwahs/B1qBzY4ft6/5z3RESGL9NiVaTyawSda
xg8aYHwKB75xLI29AvGlCm+gCerY2Ls/zZcoqOKZs3U+bL2lD/dBSMtgRuVQRzMZ/mOrrIHoAcKL
Iipvn3R+R49JwFDDyaqRkO9OWUf8vHwW9peFXtRQZt1uhnS++Il92OKoPYfZg771Aqo7NBecD+Wg
fHO8mZph1fOhhCWrwt2jFw5TAvrZZBelXYV9ZjpH6hhVfyeYA5iod86K1lTYlewnMtXqmbODnll/
tTDCp/Fa4jotHl65THP8Ul2FDo7g3/cCIP6nzfG22x4c5DWq6431yqtcPs32vylCzE8+0xUf4EMz
csZtsKRQb5gZaC/O6t/VVsXpDaWoNO5FkZHtaSQYaimPkHq4KWr48F89ki+d7o8Nasq159KJmcKN
LCPH4O0IZg5KuwZNlF+mTBnBru1Zff1GMS98TFDmpoBvueqTHBEhp/+swDRZRm5bBHlGnoiVNOR/
7/TJLjDAtpSLxmYVRJ2OziBZ76Qi55pb9KPLgjKa/FmYKoRfTyqNa6OGh7iNjnkhBQpO3R8jhtzf
uq7xhuK1QMPqcvFe/G3C+af7dXCxJQNqKNNswj75LjHuf4noiIOeuUNNdKG1O6fL04Qyqq8RgnUK
5ozzbCQJzkSy1ZS4DJuiI6Cjz2J2SYwtUeaCjkicxaPLF+bhT46RRPRZ5KCi6bdMesdewJ9N32BM
wdUZ2SPo0lOdnUIk5oP2NcZpEYIprdQdA26pHx0uRw3+NxGpy7Wf5TR6SRJIsn3WqRIvK/QosVsN
cI8NqDQT1xJ5IQ52V+eeYbXsAmkYQtssQbRrwu5ksfWs0rxYWtmDLMT9BPj1H7P2SxOTV118XRKA
O6kSGg2z/pdox2zatn0oy7yeox1iQShq7LuyHiVxydx6P1epofh4yKVhUxqSvzBm2aMnIrxprjEs
gVQd7eYtl1Y4bsfTCtXK6ME3xCM8L2JP4PDvpMrXlLnc5RVdSfwZuNcwnEf9WTf6ARsFWVMbZ6RW
tWamrkPqwB4CoqEqBXigHaSZ2NJEdbCyvqkGg7KrhFBbanskSCRhdJjx96g5DywCPnjErORVpZ7F
CVs+QE2/BjmIg3Wf9WrUGdWNwMtPdTqIodqnAwJVtDGRh57Q6jvH/W4Qg2IPE63BaIRvH3IslmHO
ed8WEtqIs+fn622UHAPJDSIgT4W9xbicmG3OYOYZgpxCKtRvBQ7dLoQvQJWjALOIL8pGZkJrJbkO
5rgjFxj4W1agx+f8qHIDYIs5ycVncngFStBsR1oQbuDZkgN8ZHAZU4aNOHbij/5cYZv/pE2Ve0pj
z7Uoe+992CDZ0EmJukKWDpV4DoDk+tjkDyge5XLcBQRBGmGgbVYvuwihiZ9Bem2TJfSy0rWO3hZT
iyepmKax4RZ0ir0dLii4T9i1wrUM6V/WxX30Fk0VbOFzIqNf+ryLXI2nTZfvXSX6rNnmYLGrGAb5
GxqvOaie/BANqVcGFH+IThp+A/82euNF/d2jOJK3cv3a1Zh9Ta1zvAE8QjTHn/X3ELtHAX1q7Rl6
WpBBijflgppbgFj+IoGaCGrA/Bl+FvJmWeQrqifVEFR3o5Da7xYVmR2DkoyzFlqtUu6Iy6DZJWf+
NYNA+sQVU9NfyCI8V8LRyK2nFc8qL1tGgF9Qpd8EJ/lbtDG7B/Admk0SFqDLoCW2XMru+kV9k8Ii
Iq0LvZ6nRyZTWmXYO9KaTFBCYb4aqLZODlPA4DrjRidZENHFchfyGPWImCJeSNUkc0nI8Dk/AOPw
PGIdw46zw7fZ36eBsS0Q3lIPYT8Evfs3mPfzWq57WD8qSewP06LHTl6EWeDqZuIU0+k3C1LgdJ1x
9heL+27gUVVYH/hNeQcl3m0buKtYMhIiniGliNiIhfdo+BK3lryXiWN8i6cCH6rp/iDF1b9lh/Vq
AcUT2EKVstkYdFz+KzamtcVPQUMkqe4g3q3gctB0hLH2z6gCjP3gzlQut+ePbYPdnB7WpgSIDbvZ
JL12MxNjnltuvYRlIeaSka2SiMZMi9t1OaZiLfOCCpZ6LM3fp3UxUa/EXIje8AfSUy1Hkvi4DeWK
qNlBxt31T5yTGlmz5RkANIZvaLldJ9UQxtRequsZGf/YF0VdTlGXx12tF9NTLz8d4vb1PJbJf53M
or5/QFGcf+YL0Q5eWrSsvQsOskCcvbgOT122RALoQAyHtd0JEnvXWtWkxv4PDHX5HaTb4L3wpQEB
8uZ0pRECfHh41/7Euu3s5qubBqE4pvee75WUjLfiWyzGyNWKHlapWVlqGj/HmmwuhZZKxR6GWzGB
YO2RIw8Jnrd3nacC7R3F6EriNOV3a6HoTmxvJZ4HvdJahiY/JoV1bc7/D30M1BZDEt4E5314o+vp
PYtC2GJW+rkJO03dr4OJ1QuUw0kJcWLlag3DnQEVBAhq9RK5nMwbFnolctZS/GvIDhHDbTF2kAwq
z5yLrdkbfLVzK/BV1uFDkWmz6zWti0SDd4BvLBbzcIj46Q62V5kjIm1Vyw4EcGeuX6aaxOPKPr5w
Rd0jdgFM3kalbm0+FvGc28u7lJMNZAOw4shK5tGxINwchVVklFWAh+vmA4keBIdEJrvYruwbPLrd
D2NXabSE2zNeX1OTRvwFPZ7ihbEtMXQ6iyiDgS/Hafvl/gH+aQa68vLXu09IGBSY0E54a3cr/grd
7MmTwWwWiOBVM13Isz4fAKVa/J/LadHFl2dgIot88uqok+SiunVrpH7XWgJI6AK8EUF9f/HjG+iX
CT1nTmP8fF74TRQrcqNgGxkFlYq95dWgVZndgaWlaRUeaT2LPr7H+1ZB7D3ZX3YKi+4Caav31+VT
3maql6YlZbbugRMoKvx3Fx1psn1ZFa2EnhX9nip9cw557FrlXRHft4XUqZObZBYZTz7WSB/6A+qh
C7qoudEz7Yk7YFkoULd1JaMSNqDLgJUMfanCMdq1A7TwdjYJ+7HsPmZvg0YgY6l/QnJvjaxb8d/p
qNNktJ8b3U9Hf6D3nDLgC5nNkyqDKNGSe043EUNoaLpgMLoJU7Lq0zh8K552n6blkofGzNR8Jhyr
M2FYT/87T1HGiZ9MmN6ZvID34Kpy2TFX8xU4hVuQw2D2RjIrJ3DpJg2NFyxvsCZ7+wIKV0IYQSVV
M0rEQQRBUi6PWpsAY0ETx3Gcz64DR8zIKmaMihWu4EddOEr0V8omvyLvrccCP2jRqJ3CXacxCxez
k3rySv8Owfel4K+9C3UK672ciBgnuHOApARNOCsB8pm5+p+JE5U2r6svcDBoQoKfW/aYpB44rur9
jStcNePryskyXJj6WlGmCG7xFauXIKelDUxeWcsKedOhE8gQYwkvBJpN7x910vTh517ySlsjQwuP
Dr8eJCSnHK1+J/dHSCuC/lfOXC3CnFk6i/NVjivyHI5xlUcJx1jRezYIriS8m4Yh6oN+Bbyj76na
oQchR/OONce8tAWEAb71ocRW6RmAZeJNAWqRZ0uuj6EBwUy681w6f1Y/dcNjGjqapOon3oJCu8Vq
gKWBbXk8tcbuNdj2G1CczCC7Sg81QzBhuu5a06WUvt5vynUyvtAtJ41aLpmCm7JHuj+uK/d99Edb
s955QeKf/Hf06G4Oy62O8NiO+giKiMBPMpCSdTCg0KdHWPTdQj3BzEdb1VxlZe4U0H7wtttIywa+
FHzozaZ0RteQ69v0KELse9YtJalU/VcNLMuxXm2IYVKOuU/O8ZZSaTBD64pu5o2LphM5GVja+HS1
E1CgFhvIggQiskGC+AgTDBJ/ylbIguBfD0c75nJZ4fNnMfqL6inxi4L3ktaZvE2IJUQozy1R1Iaf
0iGcQ+yWqtRXDQV7Re5Jwzmn5yl6UdtlR1v7KNM4ajIvLt6C09T2V0HaS7/uARv4bA6YMqDj689N
pn0Yqzw77eVSZmg8sOuWPP2Qgk0R5vXY/TRsXXSz7OxtlGamFnXmDs8GETiz1sBHxY3sqOeStSey
ASlAxX6Xr2Im522ZwXFuRsd8qB2UrwYl0bhDKNfkhyLPLkts7+qMD+9YGn5AJS8eF9S/P9yv5pgO
r3xXJ7M4t14KcijoKhE7Iaua3kUb7Uu0y1LU+TbRIOvYPfkKOBSFkm/rhi36eSQ+zpgwWIgpGx5J
CggYOP3qmHtbnlMwpHo0L0HoV2IW95ZBTGRj+v7bGbYJErFCKvcFlO6KDWDjff8DbGNbJeCJL84G
P5u+aKRQmTqzOGnpBt5p3pGdO8o9qF70KkBrbSwZdM6NiOuaoZVFFfmH35U7xWh59cKnIKf9d48P
zA7tHYeTXDCuYiMWpCjQaBZLinnEhhqZCO/ote/jVlQnIyXQp8Eqf0v/Mhw6csAxwsrQrGMzr1Dk
BAJVXhDjqIKrJgXeR1XzDlK/gRBhfhk1n61rDx+9b3ZG6oZZ1jNl+6fKDnMF8DLrOU++w9La0O+T
9bdxEAyV08V442Rs/decD8bX4Z4EiFZRV34q/gn/bobPJp+fxGj5kELujRG7UmP7hnDauk13SEnu
MLhxqw48Qg9Fxkv+iVCalxer8TAjlm963acqCm5D6oGHDuX+ZPPiAU8KLzY0tiATIo3YvvXF9iIq
3p6N9WgTqeVjNoRyhsZjxYlkwELQaFv/S39Qhw2FtUWfBQmj9mO+bM10ApWyioo9zQrmtxa6kEkj
f+aqA9JA65KoT6pOoCDuvh1+zMNagstg3ivNoImUR0BSvpxRE+fivhtjImeRlleu9sTDUf65sevv
qqeQdSUIO/L8dY7U4LjA0iK/lWmiRnHVJpspEnvcOGDG4IwofYYqxQwVqzJqX/D6l5bQiE0b5031
RCEbaFuDdf6lQzbijGnyrFyVSkar5pptrBrfvcLQLVkQOkfbuN5SG5TSndJ8QN1RN34bjwfWf+is
64kUGm8Tmi14E0MNx+a4vzK1zGE04Mwdey+cTb64L6A00wdQ9N1B1C3uJZ1P6CQ87k/I5Fl4y5C8
pV/NMlyU8fPKSca4MPW65ImXOGz8UdcDJWJ8bPmScHBywk2Qib58qbssE2ok+CZOxBhsNNQfIUkB
U1i/4MMSm4NN30t0kAL1d/lM+1RsI0UulcHgJNK4Ge4agQ9GmWzLf9nvLTVVzzvMqwbpWlXflgi+
zfXJK8l+tOapeau7ttZkRbSU/SincRvWfpGXO+zAzaddH3UqUlg/WdEZhSa0RdscFRm+vaj3yA0b
N+QE2bKEvWWVOGIylJSdvOjJiDwG484fNG9AbpLaSmtF6I4YUMOTk9W7UpJ6nWy89u02Hz+9tXg8
VlAlRxSYkYmwMPkidciqjTRPY+pD/TwyGryYovpFpJ8hP3XcBcphG+sHhpKHWBRP8/RZnt4guxO5
8eu0qKHc2PyPrvoGuIDK7Zl4nWJzu/B8AST0rehJlZAjnjgBBj84i/ZrKr9ZOMcYzSkc05O16xz8
RREdcZ4THPiAwmhKVVZFcmFyS7AVD92znFUXpl8nd7jfTSKEQrVHOti8p6sOmviiBWtq3SOmu/q3
r9tPSAQAXmPon7WUXQTzI0ghY/Rul3xo6E1HOrmuVWlhtbXYiLii9U2Il6W3fsChuTB7F1itrfj0
AZyzdhPpGLnSi7EGYLYGiuM6ErFCerRkFCDZu5wRrBzugyilnYRIaOYC9XPSq1oAHZUI9eVi8zeC
KvAkUbB/9fPPoC+HLI9J8oQf/bMV+7qJgFRwoUCbEYUmJLT9qbZOSxiCZtLTtNhDM+8AoDOVCmbj
hqBW/szOG2VaCmc7CmG0Ifgwh6bExCkph8WzquJbcYC3q1+hnlOF0242K3OlElgQTvk9yXfH9Lrf
F3xG4fCdJMuw0dbKJTbY4yrgkf4ew4FrvIhGPT+t8MoMO3L3QFttGkbTXKkQ3BJbOXm+SCSCDK9Z
y3wxlGWBHucRPAfKxQt4vzJmWV2m/N5ISlK5grky+Wi3ES2eYc/W8z7YUC+RqdywjfG2lF3lvn/v
vr5b3eDtNLTZBzjmNF3gmNEyFW6Y8LVfun5j5Ix2W8HxOP3/RXpjzmOC2mQMVXsg4V14gp0ZLNT7
2pTS88hgomawU1WyOE3u/vGApPq0LXIR73QGG15RtnQyoYJt/FQomwCd7PLiT4e/HIo2wU7vcevB
7sR+jTt1Dl3jsAjZLrIb140+HDKOlDok+59Yw722nyo61RzTi/6kknffhOUoKzocn3RM89Yz1nFJ
LBXOW1U+c1nCnEf+CuUzawCubGLz+5SvEVbRCzq32EzTJNa1z89gVa9a7ZJG7QpBG2RYf9/h/EY+
Lm9vXHBOPIcuq+9Nv/B6E+ENto5w69iMW0rcouUixOnm5O9VVlxIFs++oDRyD3kNtb4EBuoqPBi1
6KCxKibkc7k7D6jF1vvP1Su5RYgZC+AWtPhMpFbHjDcoLhJM/MqngWzAfaYcVVVSL4vMObTW55UQ
896NrHboKWiM2SbBTRbZaphaH7V0SMSnYUyCmYOiFq0BceBAgaYVPbT3BYEfod+ewSZW0sPkjxUw
e5XE//MBzKUaCQvxPzDdKklBClGVQ25WLt1frtj34VMEUtiwIsj7bYbKFR8mr59Cm5hSL6px3njc
+tAZNryh9xMBcu/P9/D9aSfv0Lyvp5nxyR1vPn111QyoZxjvB0Bqp69ba19sE33vuJu1LUokjPfO
dlNaJ5hQiYObcNolGz50i9L4G58fKbAnKo/PfK41OiZ4Z6OnrvrTDjjcxIJ3foFv5ujK/oP36ua5
vVCC5YY79q925ofHnKbvkarzKYv59sKNuDbkdUWaupxh2UEOdcps1riViwS4UDm2bvbClAUKnDxG
DSepTlSpGD46of0dFG0zRi5naK4Vd7L7ryx7v/L3GiCFenwwFpd7gCtyAsgf3ULY7QUPT0hsBwwl
ms9AOdzQQy7QMastBMqBi5x9MBkPZWd74fymBdnHW7hcClJqsNGg9Fckx/dwtBpPXYWpjSmlSC0c
EfeSWIyyRX4RyaUoNAcfYTshQQmgYNLfeWUNAqksLZc1b8cuQtXyQsn6PSKon5izVyqrzNHZ2q3s
dq4HmhIeH1MyjaqIF8JSvoCwI5x65QtrBMAG2L3AqIJyAeY/caUV/LI/l0WkdgeXkL5yFHKitXNR
j1n7llF1QeeePLRJLviuwCo1xMvJB8egLz+JTBO2uEZ5VumgvixEfn9BL6DeG+d4gxgmMjs/Z6qm
PTsyBOPkHM+byrClzbygR7Etd9pFwlhg7E//lDxeVFpiK6dZz2oal3wGRsKHvMTNLPAb9sj09zJd
U5mv7MnTuOmKc+cqSH5RldUw9qB3wLXojK1PfbdNhtmSfGvXLbNHCpSQR+8763FA+xjJzB00HRPo
PxkcHl7/yPDM99BVn8czV61bUaldiMBUHqgj7cGWOPVDF9gRX4ZKEGxyrHqZ9OJaUEjf1ukNx0E2
0/psnH85YUZFMLGq5mEoynRKQVYDjkIG2xl+W8iHBlNFpcAijnQJ4yBCdch/XUxlbz+RKBqI4fsJ
ru0q3j9FzhHb8WOA70Kl8YdSFP1kpqsXWVp5JQlQ/MwkBVsVGXRZIqSHyIbmALO04rdyDAAq4bMb
vLH2Tk65YCzZvMNfifAmj4R7hQ1pc6zKd4xB7eMxYu/8Z8S7zVlolQ/Iac/MPbkc0OKjA71hzKlF
Nh52hocdOew0kTmNCeYPFLlTzYB4DrXnXwlsR4cM1+EOPdyyw2zcOMgheiprYkvOGEWpqL1MtWfO
jUk2hWbXNpLxlGc/f7esSMKjrdcml4LDS+u/KHhSn4RTVHHnCYD+OpJMqcHftM848JVuxXkSX6AO
UZinnARckP6lNxyaL8tr58zzFyx7jLf6J8FEXSlIm/m62W5KhjEg49ilVPSAZ5hlA8tPvbWCzA5F
x+vJ2dNSfpmxj6UIJ6YfQwxlXixAWwH2NHwLJ7qqA+03qN0tVqQYe2vDFXAKUVKGN5bYst/IAcTy
NPRR4ievAcHx/k/2Sc3tVq9Zfau2OONFJLgvAozS9FWHbpOKpR76Mb7JOCp/ZCcTJSCP/TwPuinM
JIHrSiDzYIqPDiXxfeBxKpO4fo2IA53CgAHSR1Ndjk7KUtRdtDROfWjjeaX0EbmPdNczkXXc+w4Q
egvzjyVj7PYYsTD00/mfT38FZ4MrVRMu13heYsfymjLddYphMufyWch7/mBskxo7fsn4DU69UKtN
I9Xn814WjNE8beG7l6l2rByZ2G4A18nMRUknhmNiyuTi16lQBcreDMl4geoXuliQTMPXMhvlruOg
k2QaK91LFLK7d0G7FEgMECfChU8kTolzMDsYqMnwIAbUoruj87QIC/R1Tkl7k1VsnTusNz8Yfrsy
aCSsdj5LVs75o4EwLzJB7IGfGESshiZ1t8U9qvf3CidYCIHMxVCdT2kJgKAwAaInRcJRsL55VSvD
Z+q+m/BeZR31u1wOF+aIxXWyMObeqESWl5M6r7jy0AvoFJGdsX6SOSUk2HXpV1jEYLEQkfYah0pd
U+wwkpjVkH9QC6Au/UGACtWh4Mz+sumn1Z4Wp03HuTbhjc7D9yoywIz9V0IjjVwJi2wcwk+f+wvz
NnJ9J5px7BdIe70QZ7ZUtTULuPz1tgI9DTkiFYHkvd8SBxRKAv7+nXFrSmRNPlv5Qblog3IM60z+
R7Mx1xT91ZcD1394fGmjs2Cmqd57hZMgV2QZK4yS2HCYlJ/q/WNYAdwR/SHK/wEZwFMratXuQSIG
0yTgUu29V99P93/MSDSS5K7BC9R0BBGdxWzq3kA90MHWWtbd8K4lYvUopBjAyynPX9goPa7NFPJh
g+ihpId4Z5S5tH3jeuNcyxEO5bkSYEaNLHsujJEbln/tj0aROLmuXGF8Uh6Mbr1TgJdl2iNMsavf
BPqE4NMMBp/sFHKGyMiKUJVb9xxzoUA1gWd7H2ZO4viR5ivIxiOmOyXz7jL5OUocf9EOeaqw/gy6
xuDGhzc++AX4xA5EdLVsqEDTzLCQ74ozyoXHH7AnkjkGvCXg6+zuvt86d0+qog93BgBd9X1D81uk
dq8VnmF8EafXvsQrbkk9ks2QYguQXN3v/ZsNUAVfg9kTihzvQlPmuEzPaxzEq02Lw/q1a8Jo7737
uV3tIMO1RlsC38C6BfXnYu7r2bc6Q8e0In5665dTMInz8C/NLlAphqD7RL0X0oSmz9MxXuOXs+xB
ZGGzkLUHSZCtYu5E6y5Q9I9AZFxm485mmsoOFBD7wcLTBKjwZXcGFUUW7SMedMmNouXBlYII2wV5
G7AF9dKw9EmqTh4d1oqwiiFb3Cx32QBqqrRxVuDQ4qM0ECeNH9lwPqRc23ZQ5ti+AT6+x+UAHLKw
WgfeEEP01U82FZ/aqiD73BI3JWtcNgjO3Z4PR6tiMvD4sO6/Zky5rYdH5UxGrKnBUkuselcAzJ+A
KIuqYLRsS2mY2f1An0IgmLC47yxTQu1B2GVrbVfxm6C5HEAWlG1OhVcYiEctJQrO5BVIHyvEZ2hc
QgGplZnQkP4Id07ymBJfubgao1ZICKxHlt2jLHJjBubHgwV1g4JJC+GjLIEKdWP2ARbPSIJgfjLi
DcBVuGALH4bU9dHiv2ROZqNLdTiMaz2YrBmDeD26t/8Ok1Uj3xOoHG+ua/xyxPNv0Tqj6zFKD5fq
KR8qmuclnDfuDF5bmHL39qWim/2iY2OVGtjx01VVwr556jiGC1G5XIylEFHicLMSWwNrmoAwSRs4
HqpLjmvGWp6HAeQmDO/S9QMQA3Z6pCwgtwEQoJN7XGCCFgSxgZoikKqZpw7HzvK3cHu5GOAffwNf
P111GVLFBocu3pj7Urh8gJ64IUnsUF36rYLIhGd8bgcGOP0ASzLiOM8ewUGk+EMsw19FQxO0rO8k
rDL7cXTC2HTeBRJR4C70HXtX00GcCisoFRwBv1kMvtu6Xdvf36ui5crwX0qa1/tmlMnx5C7rN1Sy
dyAYN51m7nBjeFXJPvN6GnxKO/ZlmoNnnTiksNq9a7gk40Ltln9pNMCHFMlddcE8lFgOKN5rcC5A
Uu7zBrJVpn0kZCRf8+Yb0LFi2eLIrBBWNmJPlXMcqZ9+xxXUKw/Hn5wMgZUd2mF18OT6aoT2esaw
vskZeTR7OXG5AbDH+GUd+EOifMowby8aKCou7gbuotvuhndwdqzLM8LbFN2N/y1kFDdxIY6T92QZ
0JcKQcElYDBMMp7tjSy76iksbasHXO38tkhJbO47qBRMunsLRNudnqnOdcoiPFdAaM+uGViJHiIp
xxw7ngtu3Mi6jBLx6z8TxRx0/U9nC1heDZpdSZMSrOS5eg3pmvGrWJ62KS/eQKieSV+cPezIppgc
UKZC9L0tVuDy9PQJtFcZCAnOw/mJsjFrUG11vJueWPP/DKphYHL1YZmGMzAGfHHQQ82fTp3tVwmn
edvTvwKC0sVBHSd7sEV8O4+CdAq6OqfLX5xh2n5wcWD4NkUNGY9Wu9kJPIsGdAkdeQw3PQ8eTY70
oaEPSToFNJ49gereeoOJ7YYVzHUmGik/E5GeEMsVZSy/jjDWfEH1vymIxZnFqfp9GA7Y0N3BJ3P+
SwRbvC5KaqPth9NoZl7+IRy3D0I97aAl2Fvu0/8YgJx30TkNRuQA3nGqM0tWooixvQJzjpfYhql6
rIVlvg1SQ6mIoZ7fMAOq4YZjRxRn9dB3Ne24Is+vqM5Wi/G4R4fS1+I5vI4rKTPnM7y0hY81szCc
VnzmFQZVFlGZriCS0AL5akbEj0VW1LzWxPXymvDO241Wp4gpN7oY5zF2frkbesi9QQJPb/LD6obD
QVCex8ua6XETm/ABCHqHa8E/Id6/8/UDaxdOnRRFkODlTHfjrS4qSDCtKivim9nz6galZKjw7pwl
btV9Urff49VJ1ubnFDJlmorZhYveCl1+B73Obdp+w0r+3J6jqw5t+KFrl0kCsGLAC1Te4fVTfA3J
tKahEo2veIRM/M19jzQ2adsGfcxiOUDejSrlTEzgcnv+evAiXJ994G0SRXQBpcPGunu20o3hRGqj
IuhqiA//cKJb1A9C7PfCe9+vx5EZ3LqI5s9WNTjNP+XY54DNuG8b0KdeEd8pyo/tHhUGUau/UB8B
wolz5w3fDxpeBZgYvpWWw2lebhDEwDtwGXVPWlsHuadIU70npujD7uQBW6DbDE8ufJka09u25SY7
wT/e2tjV/993X7Y0CJ+yO3xCjre9fxw8fGCYcnWv8VEltKCiDGf5xXu2MyC+mCc+nyG2QONXGKvu
t2UAM8Ds2Knl/jDnJGdfUahO7av8fOpNtLHjtWUWjBN6ZBbN/NDuOu/OKJTWIwgZJITuTQKZ7DQK
Y4iOQ5WTIlNo0mJ06xKESDwuKJA6HiPbspPoxC/o7vKfvgzGWZxKyJ/p94tbMm0BSCkyZEgKhign
2svA5lh9biebRiRWQAsdGLn0APsz/YQVrpVNVifchcgjy+bR3KGwYZV2QtNZWExENNeNnXzx6d+f
NhAD6eQ8peP3FBUkKbrS7qtWv6k49FoRglJJ7fnyfhVmjl+ziRpmJQKgmGucXz2O/LObKim4MVYP
04TKCGQ3hK416mHFg+OVTXmGAVvKI7iA4XuHizpqpEEnpLdj1tRMD97Du7bxg9u2AFH69AtRtcF4
QAbo5A0y7SQYzNwmqPM9AsmeGh0xQrDclC0I1cZPhEP7LhNq3rb1R0FsEm4u8APeBLqLYeAVrtZN
zSDus7XVu6FT0HS+xDWWQPVwUxezZDCfkcUIX8zZxNFS82z5q9gDCJ0aVMZ0hINXelrpkBi0sj7K
i4W1P5nm9kv4DsRGRhMkI1NCTlbWMRpoPIhwrcY8ZsEu4aBg+Z1VjVRPO7pernZUSZuFotC45R1j
h/uaQR762c/N7wNcb+CTAfhDrkdEUFKEhcMYXFDgDoPW+KdCOkgfu/T5O4xCGV7XEd8K1bBxSyK2
aAqinl7JFtzK8eGc+Nf1os4BorPBPss6zNJ3V3xTGJgiYYMhlQPIM15GLoX1xfjkF8Mzm2DQG0UJ
pAI+s7HLVTMp73Z+ub3e79Ka6ny0HEa2urbbBLd6Ja+se0rhhLmhwOpqCa2f9Pt8p25mW9N0no4r
+Qlzj3e+QxdSeirEeSqRgk/be0yLO/xtciDArCyxSj7ZIH9tg9fHUVb3MFICwRoUK0i0JWOwW8md
TCWQRg+IDEVSIv/FOkh32r3HRrQqyPNa+CeqoreVq8EK9rhzUarpgPg/XZu2fxm/nFf3cDWmrF5+
8hTMHyFdrsQWzEtVTwe84Sm8Haj8Fcb5et9FrnvCkoITBsq9rOHjr4sqYNLRq3jGbI+MuRfk10oA
Xc8Jt07YMaAQZZpM/XEJD3qsXgJtiQCSBCXnwlywZaqHh26ZEjV8uO9txdLTWMrrrAn6lSDr0W7+
7Yvt9VMoktrJRn/onacTQMVYcPmKpHOHEbVR2isHPTIj4RSMpnN8BE/1irvvPdX1+Re71l/rS/nh
zs3FoSGJSNHxdY2dlpZsnL3oc1zYHuWgnLptK4GFVw+idLzx9wpwfRBZET42gIAs+/OlrDslziWx
j1ObH2RxgeZg2AeV4SZEjLwNAG/FsKUqW6L1HOzmtWmkVFEYrwBeJTfukUCfgxgOpWdF9Wzor0QO
nSObEV0RAEiAFEqrFiIxlMj+/Nmdfo4zxovzPWMNz2QYOaJdiAttY7R49e9mi5/yOxGcn5YDjk7b
8xJteKaNUxRjzLxcRmE7SNQeR2tSgVtXWFITMmbVzRH3yDb2lVazcWvNf3jfjFSdPHWIjafECR8P
/4JfunG6izPAtfnWspx7SpUHC9X28d8cYFUVIhc5HW9gpNAxNBHAJJxmtcmeLAyUBvigZ5aEulfG
YtHZ0G3/J8SKhtR664GB0mtufgt5dkvoU7GvSlhkmpknTRuaSuMp5XeypaP5dVFc+RvjOJqaRqwB
kujnv4E/h4HVPHLygiVgwsCyu369oTvN2Sn8oWrRiDraxaZJZlxdzpNeuaUGLu9Xi+iDfOo15LTG
pnVBiYtkuNiYON9gPDDdjnWrxOO5fmISIzB1xxizclciNRQtTfHeYixGOqxc8CKlTKgu/0SqC0Vv
YfoIrlMJVJzEpR+x3Ua9A74UMnEmJtnoPCogAlkhCI0NdeuDBCW7PQrnt0ML8VAls9tXeH0ZfUZ0
ub/GbAM7FvSO8hRbfoxceOFBZr8etna4n7qSkQs9i2bb84lNcexx8gNKPHd2px2UnqUjTdW/JUMD
jDFuQK8QW8KT5RvK1anwSMdUJG4N0/2Skq0hS2lqCTCd1i2hec4/YqdovE+xvAsQLZtqptLNSrXJ
KfuAzVq4GBUniSTscGIsBhLylIpLinLirp/ep78wmpi65m66+Ya2OxMC8CpMd2P2DLA9ePpFHzxU
i/kQ3X5cJ2F2rTYNjS8XtM+OmivllKS8610G9LEEm3rPprrAj8YUnIiYc/p1STnQiz/2aWe9ceyZ
ZnKt0v/3ft4DjFiVnM6I5gk//QF+GEUxKnn1v7JkqT13NgYgvpgwsQmrqU0oxOrBWzEOUetHYE5o
yh/vNbzvrYu2nkyVuicwA1Zq6tVCoZrAdMvrV+R3jh0X8sX13WqiYXMzNQI9wJcmO46QpvhVfz+M
3QFeGqt8JXFffiFXNFnZ/rKQLJTbxQuIPO7AFIyJ3x6jNP0FVFGv7/Eim2y4BLQ3Ou1dsvyheHkR
j3fN8RLW9QFgvQCmMORlB6bPUSyjsbq9aZcHB0yObs5yAr/JIhPV8fVuxLU9eVHKhx37LB3ARjCa
tu9FdHZ/1e2Wl8ZQIjJRrCUlVgEX1MuMJjXVLZZVXdKhyb+kMJlTzld4579YRIIxB3lgGDM2gJDe
k5YhHxo/1Sq0EvkGcqQKyhcRd242OOCUINBTlsialFlzZK7IvYr1FrU17hebrcIADh3G8Lgm+7pL
saSJBydUoiTiL9tQC85NPoiVPluhOBs4MR7tZAt0+HOD9GG/msJ8d6ksbYdeGMrzreAGp19uWYQS
tdCXXUCNoT5QQpERZiJrsKJJFqmA3Nt6r4n70c3/kSuXOG3Kt3IEjypXsTmhVn2thuTInqBDlSGA
Eja5DnbNMPfcpNZTjWUr6L6qis5IXKzElBHq3rr6tbYV47B9ie9OOOYbt1DCGfnXN5ZqIuzUYHsT
Z2GUYQs3Jt+TcKzzjTESXYHrDJKCxN2ZgMCn4NrzxE4y8MVFTLcK37VUZ9fJyIqhR8UkuBU7T2VU
56Q3kVqk7MC8N44u9YgTzTXJxYFsuiEFBAIbA9MHOLrrshYoZxqJYxydufOIYqUgVFN0uTipNtq7
1hs4XG/2780TYcOU3If68RrHhc7GzUkMhnPIlJ05lghU9jqVPmYKVG0s8+JSOSAsjZPCTBvZvcVT
2uGxI4ff8SIQA5nyzAajIykt1+5+NrGwQcyg
`protect end_protected

