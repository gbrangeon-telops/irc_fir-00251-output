

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RZm5UrZFV7JOtGxR4Pzih7NQYLp7LmPE59R/6o+hZN+ZT+nCA+l5YH+/j+E+cmHHWo6IUrn/ULaG
ZkaGINks7Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MRNQzUt4f7a/v9KMrin25EUCYvWi/twJzLlDdceTmDN2GCvOURSU7hHpsmsqqCb1xCeaV7xbvs0c
MXpZkAPeQc5Coi1irNf+9eKbc5uIh03B/PevhS9S+La97Aj9rjHplzcZDEBFN6fiyAdKvJgOrOyz
87nOO0u5LoaEOeyC6ao=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L17wVQWzSUChaUkUbjAqDK1dFxRQ9orAmYas8htY5fjqeIDtBkS/PldQL1EGRGrFVbxZVbStDyiq
iWMlaMSfJiAW0codwFWqGkqnH6YMctbqpTZdQPbprA8qa73Xmy9S5tgWXo6y3vZys5HBTFHxXMXj
HSJZBGLfj5+GGMkAkDYYBZrgDs/jxx605zYzRg+wKonRxjx8C7c4r2cekqFXXjEfMC6t47HLGKZO
Wp8oqSV+SdxjNfsxTeAcFxqhiABG1hbduxwcNIQO/0mgU7awDWqjimqvnE1+KO7vQU/MVpl+J+Y9
bwvxkUUMkYnqQG/HGWvvQ7Zp0u8+rRyDh2dzOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yJG5RZbV6QsAW4khC+YjJnbI2jNRxPOtee58pTXfgJVvj12BYVsRuhi1xiVJgak8Vy8V0UJ43Wc3
ydXie//gOHZIACOddgGz8WdlyWauaZ9sd1K4GlV+vX4K5HkoOyunq5QSLYwU2X/ZYYkTAGg7My6m
h1UvByaO98o6pNd+n1w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QjcZeibYm0SAHW7YliT2StC14hkmhpmI1+m8klXbQfAK/yXQ8NfNnDZicIHqHpAbgVQzoGSkcmXa
qhjmF7JhXI4I11rujpUqz61fAf/3PeUiYimqp9l0xnePLlrRBeItzqfetftMnQ8hBAuI+sARuLin
j4+kHDvo2V/A6kndknmKA6lyd7gI8Mgzy1xgvua2Bfq25TZ30r76kaSXXo5N6hFVjtfwPGqnYepq
02yTg3lN97x/f3REjUh0T05iK9mOISMgvqQkxFwl6hBnLhp8WW0zJBjFvAguLZDf4CMBuYBnnmGQ
axcOzl5DWDcYTgPm/DTciq3eoilijus/JUHuFA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8000)
`protect data_block
P/MuG5TF+uMCQPWBY2ojmPhhgQf0tCRflbFlymFzJe78xBqI63s72y52wIpVV8oVK5oBPZuw4Kip
0JPpVYYugpRtWvF+h3zX1PaTU2kUcfXQSR9ndoy5Wb4jqhMO54GRPankB4INHhy5pNnRa/TEqeZj
rkcolwh4kBTzQNel5VigRbWS46d0G1FIikCFefHur9YaBIh2wQOdwt14ejc8YMfjJx12oYiCcQiV
b5GQ65GQrZr06L49F8z6V44lPvKNVbUjGf1xnO8Hgdf6R/9EstR6bbLmZZcWcENsTM+QdPBSaFGr
BBUEuuVTHB1nS3/E7vDtibjBlKn8SIDv9Asg0hSD8Wjf0SGPNKn4pOTBvWzYB8mJwzCEgOCUKwEw
R8Zq6fgRsrcYfFm8EoZpxVvclK3S71lKUj99T5/rx+892mFekkfnx31aeA42LHAuUJYBS+IwPKDI
4/K6OzVjBIxHz/QTpVQbWvm7Pw4Wl3FH/xNk43Wbs7KNbB7TJI2Xa+vh88Rdth0mz4dgYlhJXx0B
XRDBvXnpUkDiTR9hoHi2JOJYQpkbSIAtyr/P0rBkdXf9VCEfnhyfMj33N8tALO7v4YvMspC/3YWY
DUAzFbv0+mJiTIpHAnuz1xyFL05PSmCoMcml+WxlTdTc97/w3efM/80P5bUm7hAtEi+WED00U1H9
Lj5rE02O28+MagsNo7hTaPkTqpWf1A38ZMflYtQtb7DF+7/capSBwdYviihKuk+get9Dtj7jmxDy
GSuqekZDjWYH6yuQv5tbXMAy54HxrhXIEwH00GB+BRcqk+D7fROaL9Q8sDeV8+/QenTkkNw8iKK4
M0SIcbJISnXcZQtyWS1A0Y+J3VXeFzj+Q+De96HjiiK5EUD+EZkHYqtY9XLHo6x7XScL71E1bQz2
H18e5IPW4Y3V37CDa5LcHmzb37mI1FCJl8+z1aRPb3pH+ONaAFc74IvopF34BYu+2TGMEjyaRl/B
aOfML+OugckmgSNBuAslzHqB6LDHikJRgigHqOqzowCbMiG85TfEar8/MVpT8IxfmX8yq+mJWHOB
OEttCPW4ecgaKXtFGvYjiOziMaVYC7wZDdJTJgWC7nyAQHjYe+dRfCPNXzbM2Vh00eDSnIzjEoA0
+gmXIy2Dc1pH+e9HRfLcQ03AY1ByZNmFg/wbORHKUha095Ks2YdN1WnhfdJ/ucu/uI6oHnMbQy9P
1XNLpHywglTxTGNP4pfshUzNPjk+IUrXA79ppwHEnP4wVu8jRIKveno9ShXk7eY6b12TDWD4/8wx
0LlxDhjm4C6V553iiJuxWjTyWSNZjn65MmyyfYxSK7NgMMHhOmpCMnULdWbsIoA+w9Aea34d/Gko
KBGfx+aBbVA0q10em9YShbBE0NgVwedRPaJH1ivJVkWVq0b530uyS/gcD5eFuOwW+fuLDBVB7Oj1
KHdrqHjHV/0GjzFBIxbANS0OToAAeZ5rjMceP93t1BPRVnge1s++nXyizLFRJBdCwvLGhulMFwqh
WpPhVmj34aWk+DInNdJcvLQ5qgarry39Z0jQyUbxfqgrSsmNcfe/1Em7NmTVvQzWdV69Nro4YVab
VfinodN6RkkcPXmQz94N8qFxFSYEYBnQz9GWcNmqoMfkoTRXgpMf6svZxsUpCtihkLLl9lyirGDB
dxB2feyyOagtyuEqi1enVkIi67vxH1SskJie3nX3PaLaYlLv6y+URQKfFuKPGm4Qljp+63SrjDS6
IJ+koZq13EVycE9xrak+tNUK+gsMMBtFnYtCKOgXcZMCZpKF93v9gE/L2oFt6FsDTlGYMxssFW5T
GlPMvem3CSzIkC38oUYnhqfl5TmRhpdV91dkceobh2OfHfjmITzNJ8nsBFNjhlSmSkOthUFj45vL
bFRqN8Bxpw/TK+oVyYjqQYZRarCSixq2BUQvfQfgY35eXIIpXb5uXFnkSdnL6ke0ncjLWLBS7KbM
o1UCfXYpg565JXa5hLOARHQPR7Tw1QE+VRIVLf5bzlfAxgOL7EZO6joNMVsYvIN6a5Of8Wm7/tuI
WM5TKZ9uSFsVHnmeW74ZCYPZTEIIY651fApXj8PfCKIU3vP6uMVzanDj5mFYyRSM3Q+c2uVP0SKx
LGUJA6cSE1lcIk5WRHWlypFwQSUW9jrd82f1qUeMG0Cya8mIXjMw1dNA/ZjanYckdRdBKMncHUtG
mlSNJJXL8CPIX9HIG/we77dZon+mPnc/jbhaSA2ltMvUVN8R2C4mHriuL6zwIr1naI0jmemdLqTO
V0A2VHg9S8GekCquUq7rgLp2c3MqhXSyPpVE3WpE7D4ijuw8XHmBIMyJxRAG+j5rrB3tnyMV6dPI
T3BesXgqtkQGpVJWEf1MixI5JGyde0Zis3LOkkh5p8USFG/RPjaFnElVD+8WaCLOAjog/6N1mqJ/
ncyGGJmEo1HDp3qUoItXskV+j+ASwlwFiDe4KWTtlul4Jww0Xd4gCU7UdmshNFowm8LbBzCCXRC2
bkQC/gUJ6V50/d7DURvehg5GaAYsW1UNzRSrqxnAurKvsmSTdPbN/CAr56U/qgHNTCLvowwJBvbI
yiUx3xwqq02DuJtM9W9Ra2mps6oZ0EBvequcRM7/MdzdGMYyIFwZ/j1wYzM9FlIAkQIzStqa3omB
yADVzVTHbmJhYVZbEjYtXBUwZ7CjY0EB/ADayiL0xSqlbo46B4sNsT+dgCv6CsvCzal47wFCNh9n
1+yAYCbw/6q1ktcAJ/53Nl57CzY7s/aJdxcPFMdpNP5pDn6PAutZOsA/sCtF7Zj36wXIHPwB+4Lq
m/bU4BBZlrIn2dPvzplMZt0mZSthDXoOMqw+Za2NMn4Uzb9KyBsPnRObOAxi0LC+/u2waxfmIhjr
H0GdgDN7g3RUdN4lNezhvd65K59HpA1j1E4PFe8qV+SnJ0WCDf0iK6ck0plx9cYyLLewaXyMzi+C
IIOjDa8X8M8nvwBdkfsw2jgQQaDxgZdpGuhAcdCd/Oms+LfckwfWkK6IDvR0njgS4a7j1VnAjJ8w
i2FkmSxkud4azxyzOiMMOz5fSuxLL4DrrRxmCGi27FBsrmEKMAcnx+stCd7+wR5Fw+qEvtUY67E6
b/HawJ1pCVS4x98BwxOWecDlBtZ92NCxoOdV97aFrRrDS8ct7cKBMu1AyOC4lCrurXbRotFd1CXB
6YUXxRj8df/c+zBmxqBMiZowGQdmDMM7NIQb4zFfOzMacTQohWkgc5EbwLmquUSeo8wdm4bzAgkQ
9+eeXtS70Thb8Jals5yZZ2TUaBdN/IF4o/tX//YAbzyHhNW3q1ywTJUcIdd7fJewd6x0RTibhFYU
5ZuxqEOWDsD0Q64Ttp6DJOzln2oXb33piobWCO4lbzrD6x3PDdG4mCoFDBupf6/gdxAvToX3VmKc
Rj2xbe0QQeqUsY/x67Z1vk8tuA78ltft2p159yXnQTfr4aLxKXs7vZyRHciuZbhNs5xQifMhg9Bq
GxVN/Q0c6bZDnoDCmL9t3XKz9Cecjw9kjvnAX4ajdZtuVmoOhPy9aIaczuNT8geScZxnxNtIUDFx
vlkl3pVUrnUlnJfwm5OUE3oAnsGROapKrdB+hh7mA8WMfRoRDUfO+HTDFT3uaHwd/V4IBYK+x2nv
VaJU8zzlTkdtIBurCit6yHCMFzFZQInsBexJIKjVSxGjQ4VZm42IZ+4+Yumg4W/JXZE8fo5jh/bE
96QYozV/hPhInVnWzaZm6JXTlrcpbfUQpj07k5fLx99FKfi7iO46XKnxM6zZasSXT7jVBrgM92Iv
6Zz9LJdB6bAxD30zk4LkvLzSYW0sz2h6YmegLTvqb6Am6LOZuluke7VGMKh1kQNSp1x018iZuy+d
Bo6tnYLt6zr0u26DhofnqPUPAPW6Cs3lsX9Zi73ugFTfixuaD1fYShGck6wBPXtRkH0UEU7vx+3O
lMv+b/vrRe6NcM8zm43LBefvDpSNPr9BRYy2qEoSd5TuCTKyriCElGEXuxG9Q4o/jmV0FhlZtszL
Z9MCtnXbe7ZhjONYEAMPp9vI1Fbo5ukxNHcTkLHQMb6J0fur6oam/HYBOiLH2ef+1kJEmZXuwHBo
LLI1nBFwwwBtsiHB/siTYS9Dy20t0tuKB1Z2ZpFordcMGT47Yo2vb1Z6KF2pocanG1nJ8ckjI4xP
6kcyPU3LvTi+DAfe+EYkB4at8+kA3WIkUtTpB5MjiOb3gXTFrmpnj8DbcxjJ+lQwgSBDdECUoECY
RWbvDNepYt4q1s/KZxFoLTBTN4TRHO4qXc52rciDTh2LLOrFHm2jm/crEo5o0OO3NOa7S8+v+2IB
W1APzBir3hE3hwBRaJv6Xn+qn+Ph2k81RDnyyefRvJrMy+s9E5Sw+v6fziLkNU81G06/OiJXEjGC
fPGQUKg9s6bV+evoa3O08/QGgvZM+74ElsoOeQwX6w9ANjJ2dTfAhdxADXYFuMUy4wYP5qXdsXR2
onj/ZN16jxYa2FrPg+ZltqbL9jvkpNDBoUJKySCMAknWXqTanIw+kpfHgPOPJCz2ZBP866U7nGZk
WwRg+YfXTl0NjMsn+XwK4mIkN1EOhv1TrXauePR/X79lmo80eU8h9IXVbHKSs0gtERZFBaz+zned
FEiAZA7vJeokeBOlZ1HFqH+jPn4tMh256CWCAxqHhifTBI7TV+J2RF9TrLelxD8kDxOhpfPYqD1y
wQDBn3Jj6JvET3IhPNMZYOd9paoYWEjQQfA3Z8lznXCCcSNdd9bGiRD/8l0rOksLWeG7G+N6y6vf
6jG1dkPZ0q/foTstnBYOUcZp56UTFj331Mxz0SCETyeaFrv1GWpYh5uDfIUJqPzvhCspjQ2Sg/JC
zaElWnhaKQKkVbZGiJv4L8ldxX2ny/qL0QbFUEIgxivfJRDtbiNcEnhd+JEIldJhUaimCOzE8Bzi
EtAs5j79IB9NkDLXZ7Ty+vx8m0DRcEP3fEfbYjWTS2/miVoj0PIb66z07Y7oyxTWoMMjC96a2cWP
vgTw1f5N4fExtqN3bgyWyBuCegvBJ+jxFULWVJs5vvUaqDT1BuXUWY+362Av27Kuks89HL13fAvz
pdRdKoJnyGSOQqpR3kvMSjcd8+Xm236rHJpU2EYeyyKT9Ye5Gcs0iAynB/BDVuwsPMmmnmGJoOwD
VdAuMjf7JoFsxob5R8kz0YXSTw2rCZ4/lUydkNw8rIUcQClVl0EVk9R1qE6gPjXrw0DZ+0k6tFf/
dZxPVNLTHzv9uHqT7751EPzwilAjThvWHQ5kAFVofSvOc5m/oUao0H24I3P5DnsnB8bIF9rlC5GL
aBlFrdCJW5s4EhTipIpK6REgnxgrWdWNbmuZ4X+Jt4DOkQki2dxYAlJodNBmMIBZjVKQIVcqR0fV
1/Ouxmr+VqDim3Pznejq52fAZ9c//8x9Hz+MIyZk28V1hMh7wdgbZO5RZdOOHwPWUAFHb/WVZkfC
Jq1dwmlAVaZt+mb3d+FZn65pPZFm7H5XJSyHN/Rej69LmoPCK2p9b9DYVaZH5hMIikNuDAdRWMFJ
b44D1Tnpk9RpdNlfq/J/ipL/YLtmJRmqVE9Cz/v5sCI0KJblfVqhJCOkRohPI13uujELbC3Ugswr
1GMmftg/OafhtPd23MIH/it2JIIHUT8llq8aysiJnfIGEtBTWbn7/BGz1Vmg3F1kks7HuUweQL8M
Mvd8KEUuZ/6aS2A7lMSqJfM82e4N+r5DzbIfL0UGif+vAjRfa4RY+/9nIbqGvMKvQ3SGDdbXTxlp
HzzF+BT0UaPMGFBPKXk+GrxN2iRZnH4tgnOHn5cca22pJXW7hSYCA2w0Y4QJCVzmg3/dBUiQMCRr
a7jrQy/eygHEUf4HRKV/CrU9MlH41I0JnaDF5OFWgxFHi3fgAZM9BABGmm2T3Z3drbFdliuJ8w7C
G6zZ8ukrYA4aOUD895bYlgALbu25gUp4Ig/w0c/vjwZgK51yImQxmRDDi2OcobjX7yaPouInD2FO
2u+eyMiyDjlfhLT1NVupgh+R3nZZuu5Ti1FhAuz99ZgnIB7OIg25iRO3twkpc6zUQOPdmeWufgvg
zbYSEwdt0l6SG4NCF5jcHtqtA+esoIhHXkKaPB1bMB/9KgiDACJA/k5YWN5FgDmbiyq9lhRZYeKl
NeoyMq6gjs8ctFqCo8umQiDE6E67S981SAhIZH9jzE/+AfV8I98ZTWDDjm0MGHZIO46jF34zK5mS
1edK2vMKu8X2EP2scPG5YbYwLFA/t71u+09a/1Z55L7GjSik4ghOcmtwvO2vIbuJwogrXh4tJDqP
rWEOC9OEVHr6GRHjUu+K1siuAdBpgURu/HsR8ymV1hbUtXnIq/b8PwtaZQuat4H74E+iZVYOyjhk
/y8jbag7qjWgrh3o3kthZt43mfIR68Su6JRX5dcDVMmqFzlRkxYNQ0xOOqF/8jnEQ0YAuKgQcCp7
mMXTp/spxGjYsD+Qdxb5Lk5UMg6+7fA/g90/8z1puh0x/qGJM8Sq7H5nJM1UhXAJsWJWI/BxP0ku
R+bGjMQ/TTl4tdeQN71KMzuj4IWQYMcxdepEjYleQ3GncagXXhti6Iid7FaviZzZfsLIrz/jnn0B
eKYhcxgZBLoL3F1iFGZsKPpgAFPSRGdUTZT0l80wzwiWIem1iWWS7EvK3/9lLugs0JxFu03tmG+4
FKMsQDETnuTIsHDEBDZiBkRGJcgPKmcIIIkLXa8u+HV7s7QWDgt0ojMMota4zoFoGSzQ19H/7swN
1E4FGR5jJCTq18q5RnkzgoCmYXInzb7IMYtyqb+aOdSQ/2QQvQ78tdFp50+25QdS9lQm5frfnYVf
OG57ipjeBOZIgjMSvIevU2WAo1FDxXKELjU+Fyb9JY2lKfHabspVGreJ6Kc9srDDn1ftxUwa4EVo
ZYxSwKkpV2eXt0Fh65kIA3A1Q3hBwZ+qCQ0ENQGcah+TjLTDaGt8y2r3DFuj32Rw95G8XBpeRrJ8
hVxWBLoljiP3yBHs8J7wnuqQ8PAc5AcLqNc5iWfWZEClYNXH3mFMAgg1begNFwfGLgaroAUSU4VT
nunTqTh2cciEPng+2RDrd0DASHwjYFixehVQt7rGlybh/s1RrU9Em4vh1oCjOJsEBuB8MZqMCt8u
UWmrFIBR4e70p7Ykq+QgrKunGnm0ZIb4On2i34quow0+J8rhocIVGHzxj6+Ljw1eqOwKeFnMBWT4
lH1LMMLrKKIiaF/L+deg1OqVFNRHJEgMSqTkhUr5bYu8znfOr4CXVGLMRRfLuAr2Hg1v+bgkmS/z
Ylgv0hwWgVGCXzm6K1j1oT5bBNJHyBLfLDO+ibE2OrpY3oG8jUUMm4NoJHhYIrkaPgPBEg6qpSa+
uKhsci6VZw/7hwgubLDc/QNTAnzT8jJDuAn5q1N2VnOIwp778GXpbPKakOm031qfzL2IyAon6SAS
1CphO/v/umT9IHiXgFOYA4ZXHBOAbigWtFuguD7Lc9YixytE0qKSF6QA3mTuGVbSSR1HT9hY00H6
nKf0jnIuXKT07X510Y7qhtHZh+NuPDiQhBS22jEC0+Cjh/4acmhN6Fuho7HqsSLzcdqltZjylqO5
GNv4Vuo7jF6zEb3Ce8OJh3dB1O7Yf2fHaSS1CpK/W/F7tpsaje2Dwm5qPQxjZDWFpiyWFrfLlFRA
tuCKGEFwYLV2hmqa0ys4fyXZNPtmHLV/3zjvJwvTNY9k0jyCzuwjaR+6zRoyCSK/LZEkOZxdBQxx
bs2JOZIW3leBgogJ1ItAq502BOzleBegYBmnvfV5zS4bIfDTaA5E3Ph340bEh5r/EBBUK0R1mkVi
gnD66K1cbWQgn5RnusYZbGgJwU4U2JYmk0cp9kYn05EuuHoV6+J+ReuWymUnJmEJvOtKNzR0LH0v
SzOG0gJodRuRToyKfxFWZ8c2qRelpcSgULgrWqYm0rknnaSeVNvgtIfQqVsXTK6v1pnrVlyUZwzw
xLV+YzrlGimw7vjJsHerNV6ga/unjvMRqVQ23YFODb0YA88GKqyhDTk3/jEzdmDocWFYf4KFR4My
1PJzU1e2v60DmaybR81yLy2RKfh5RvJKcUAJZE773WaCSibrNNwIvt1KkweSRCHUpOscGYvNz2A4
NSDAtE3n63estJqFQvFIUTOP8f4N8MM/UBZm7ERjkMTLADm+MSOH0dDF/0MQMNdy16WVP0CusCEF
nES+7WFzh/r2BpSOAKVUsJHrpAtPcC2UOjexiypyQ+U7Wjy5tzRFS36JLB9nKvoH4sHMSA9aDgKs
5hO3lWWtBgDkoTXedb64smBD/oroj2WANgSBxQazmStB4yBfA8g0SG9Ifxbfv4FONGQJpPvOZhq4
A17013Rgr2w8EnMw4cqdkW33fSSA3TrZ5ZgBRbeMrg339+3t45ISgI7f64xHR8uOVyY4MjTqixmo
c0yi1K5PaSQCA7kNJj2qjwrd3CxDdvoPSoVMW1EmHLxNk4qy6Ofu/o4CvledMWdkgGap9JEbhR/g
3CS7dF8szZXYnN1r4jgCNMGFfViR29YUhmXuIashH06uiNYsq306rOxLEyPl64p0+BG7Uid/rSnk
hz+aevwgH0zMMZUGXS4aky9ZdD1SFKXXmxmSQk2NRRXaWVad+O2mZ1gGh3XtO0ajmKcFlsywVqrt
sJgj/UOch0zomKps7ohcQmMTOguGoT1Qdc5zEx3ZLt95sI69R+Aw1eWu4wLD9/156g9vPa4DRDZ3
6T/oooIrVtza10IL6sGDiBwJLfMXlsz1CwLz/IbNowpG/e0VW2It8/ysWIgKItOnzIhVH+mVu3MX
bHLlIc5cpeEFa6n2+HkAyFbmxeaUzulPfAQJq8Hrsf1OOJBx+eOEmMtWur80t+ZEcuWD48bkEjUg
oBJ9SEYUeRho/6CyqHgKWI3T6Pi7A+NQkGQzz/dJvhV60d5MMFsPi6JsbgrxL5YcWAvH5je2bI18
a7YOBVxChvV0CoEsVJqFikCvfOpMikqI7aTQJVLYUjN30NaY7yFqFiomxV1OTCODuHjF2XssRnWc
8AFtCRjl30q2Xk5W5oMAV8OWO5hDpQbhu0ixMQscb1uyFIWxTdGaG8TQuwuZdNvDL5i2OJHyXzFc
I/3IfVJy/uRHRbL1KBMCI8mktITyHzg3oEWAw8BFieoqG3uOjBNWpo3fT8kDhzdlNUwzs1fWmS+C
HupL/5Vdxzy7ZoU4cKPe9UuECFUMiPo9Yi6mVYAcOCvE8z/PaGHG3PL311DSa4ArzXzUacUbWK4M
VcTspAPbbXX+ddIxzXm3GgZHiLgvl2rpuZ2GLD/xda+Sw4w11Pex+9r/UItEKhRMZhiNSmFpj2W0
MeMsKYJ20Xw/rqTg1Soh9si3U76rFyU9oiGCH4MkepBJekP7ZabJmiTnWx86XG726fZ44ivZkZGm
CRXo8F153WqzgnyfgCYS9b/uiL0CZvHHhVqvtFey6c9Hv740iRKXHh7mtAjIO2KJCwF6WiAyAXyX
IdDH0+Ka10YAIK6pMg+qi8WKwdJC5ojpPCWcjZvXKRCp4MkHOY1+e5K6geAmv3KTJjQU1LNkyNQQ
iU8B/Qd0brp5Y1FA+66AjYq3m2ANtxyds41PSY8OX2Gk44283S5h910XCr7qw5c2TcL3cRZA+Iq5
OgYhA6CNNkorOb9IK9srHHqbUZJBJRPd6Fo2PMuqJkUNNaRc3+Oj8MRDo52uPxmZ6/cCcKFhSpqt
O1PBMTVO+ofUtGxGVVfZVg7vrG3EiDUfnaAnmDgEWS/4QJI/Ig1sUXKFBIlEUGhpgld5WiQJleSN
hG4cK+pnUXAn+J99WtK1ZH+SG/ZNLGrJB03SWJqSGJM6iotBN/AuD8IJY2GTl7cC7zqY4B7yWPsK
JakjcBRpHCGgQhBzb2TdXrmYQHe0HZ/V7dzcUcqaLDKQHVmItQMGMgpUKcRfh/WUhNmCScOv7gGc
fRkB/lQvaX1cnibMWeV0ko00SWQErm65EaKBPCBV92aIauRsAJZ/C8FVJgIqeBLtk3EBfjULXZpi
ymZVRkPXObu51egz2QA0yOwXahAS5tgZ5PcbkQZHFyh/qZptidxKLto0an03e4dVr0EgcOSV17/h
Weu/MgeNd2GL4tugyYay+bQZdGNjDcsdsDOHG9nTsKIMcYO33SbvRLYekglJ9M6+deTuDvcgl+gO
2SBW2tHu/1e0Fd2SlP4ExeB0l0DlEygMx7/rGAcD4/Fysxvh0VfvZhHy88JEF2ntoVJ9EGE/4fNt
XvVOdQKhQStUAiEuT3ZRBqLX7ZeKrdecvKh6A06dGnW3Zf+3B57s75joiqd55Srk2fpy4CGu9p2i
xY/QPvFVLTPVdHFnqKCyviWrq34hlSYs20i8ypcxBPu94CaqppuQA0EKN6Czz69aIVQtFIgXNQrs
AFpZ7zVyNQYkd7XFeR3RQQd5dX9A4P7uSzGVKH6fcOYI9Xre4E5iR6alP+F63dRjMfaKorSIR85n
Wvr2f7MYLd8V06U0ptG+DR1b4ZQYXRy7UIld0N1ppt9ucwu96vsFP1E4LsV0+WQOBylddhQHySmY
dmuSoTeZ7jXxq96G0WHtEq9Awr4oVZCRlKTqLi2JaZ2On4RlGemRik/m0UDxaBW+HkIW29pW1uw3
pq0wN9hw+pSu428OepRBMYvCxyQ=
`protect end_protected

