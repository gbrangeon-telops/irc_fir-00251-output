

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VQBfeXA4hP5orKlsy+AFFAe2QBxKheQVMjP9iwMw/NM3O4tSdVMF5nSpUCi2zqd6Xl/0+S5YrDyH
MbW21sN7bw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NYnVtYYKs1fo/NxKyeagmW8datCnZRNIFQJ52Ut8vKAvoM6z9G59Louyi6BpOXJlK7hkOA0EyUcq
xnrhn5QTbG+/jjVXTRQq5boOLx13BVtwMvklEuJLJaUCJSI1mkPVMU1Tw6P0C7fzMTIVY1MXBSgF
huHBAAQ6j+Ca7SHEJMc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UdRiCUwOSibQJYHOoWlsqKR136XIPiU7//1vC9LO+s6bwL8gocVodj06NRrITDP0xKYK2ZTek7T4
6OlwV+xWr4k2Xf/sx0trTcVrHoE3bps3QkJHk441qMX8BKjF5fCXU+yOMX1xkQlvuWSD8+NvN82l
uzCDbBA0KjOv/IsJg1WHwqG44dahfC4qa2RHQtygQ4MsVR/PxcN8lnUdpguLi+YyGmh9q+fLgQBq
cNHly9YC9ZC1urY1hg8yqWcJm8AuonE47dIMtl55BTxzCygZ9uoRy68FfVsLU7NHg3O2kl94A2uq
uulT+/Y74MIANEyVFkVes/FR1hhgCPd7uNhwkQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tQM9oFLCOLGigsR+dGte9FyrpKbOg0a2HEe24uc9a4zzPMiWT4Zq+VUMyysv3hVDjsM6Rhdx2y1P
MMtJydYUSv3+V7JQyYwaG874Tc20f583mvfsydp9rtOQQwZoTUUdaw84/pibQ9geh55pxtJYjyzk
ltK5Hf2dDqQ0W2qoU2o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D9jeI9qTFJwFpVSxwOhVsb671/UONJ+BqwlU4oe+K/dJiOTSOoWnMaaYQ9Sgy96AbPfvmkY1YYgF
jNHbjBYJx/eNgXJH2lhqUlU4xX7po7K9tZYQraj2oMsohZUwz/eLwj91c7VL5ZRmCXaHh3hDU0yM
tta+u+KG7UfDjSpBDQDdNd7gt/bWHfns3Zj0BeTNOQ2o2kTzIQxImWuXKku154pI5L0sF72lK31n
Ls7v+PzriYFrSA6JTTtqAnDF5uCY0O6Lpa8FB2AoeQSutIiakkT+T39fToTawon3SeQIsthaDWDT
WAem4lxQFA8q64KvDBTwguerI8Z6/8BM0gLy/A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20752)
`protect data_block
RknCXp2BxTRBwf8Q+oesz/gFqgP9fZBZVtScBSE6ZtwKqW52Jv97V0tIMQ43ZI3CrG2MdazJ5yD+
CPpZq/7T4w725HIojvfez8Q0JENiY/lKAX7BzCymeJA345SJunVUzbaIcw/vb4ZXkpfGEBzZ3c4D
DGehVElUxD8DdOFxUdAj7Vudwkkg7UPzynNOQ9sQiA2D/I4P5YF2sQBpyhUIaEysSZPfNQbQrDG9
bffvAAIs3IARxleG8VcLJtp7K1g+vQZ5gpFqZ6Ved48dXckE8sanokJPmA3ULoVwDupsFLf1AMNO
5Nw9T3uhIUxkvEb6aNSwMaRhpE6PxdqhCMNAkSuPomCxxA4/1woU8IgkoDFr5q/dLl+0xw0z1B4A
9n/XK7OlWpgLsLre2i6PGUtremAYWxF+APInWO5I4kvk/pBohTL2egQuu/HiZTdkSLLg1IwJGtec
w/Zyw3vDpWX87EcisTOf46m7CEWUBrx52Pcl0oHvlkWXvusX1IXCbZ+GIylTrqBOkglCoHjvWgee
8WoOiKVe+oMt9uDdmFEJkmBdJ2e0LTU9SiHLAQbLuuhubVp1UDeYTMP2K+0/tLFwHT/wFpTpkqgD
wqUNbf3ScHFDIazRH9H0jbeQk67PVPilNdYZkQ6Tbk0/V1RYE0dOYWggufVJIDTZSvCr/+IH1WHB
+OUMNTkyjRtcRBpDdbTANHfqCKY0Dg/dDmEhoux9vg8K5tbs2Cy7pFv18rML9G0NKCjvlHSS83Mf
SGiXXwkG2CSFyBU1OeemnzwWTt4HOu98gohuanKOK2tKtZ/q4r9sB9xpQj1WV9PqN+jiWdbZ1F1/
XFJXK+aRL9XlKm/H1v7L80rrpJ03KazRhBkTK93KzxO47v75v04ufc+Pok8swI/nU7d/SciUHPIo
2pWpnG88uU44moHOl1opfWQb8FXrCOn4ff3wEcE5a99peNQMbq0lsNa2CKrkOryAH7ibIb5mVBKk
oU0EFOYD9Q5r3NKP7c7ngaB65Fk7fD+7CM5gt19OYTX3lKsvnzWWZNIxlfJpwQPTOnpM70B5ZTJO
auhr6R+/WDv1pzGFDiUoKQ2sKiLx5iX874Zaxh188XNmK/GHjmxiYR820Kqqfmb6ClpWszLXkirv
RZ+/aqhGdhkDIYQGl5kiT0smYFsJHaDMlaESeEnRshw3gfShCxO7GxAf/x4krUJdxNwDJ+kwcuSf
zbSNK7fZMgGSm/MaWPR0+7Imq/cATk5d3pl3c3MkWQfeqOJtXZqa7aq/qMRbmANwQ2QGOnIuwcFG
PxBVlnYocI1EQJ6x6woDlPCqGLFTH2UhiIG2n3kZCRJox+TYgV+cTV1Zg9JVyFVy6NOwMrQvBFNW
vxU2m3p8KyIX9ikLBC1oy1PhBRSo91sJTuQy0bitd8o8oozUpugTLeAeEEJHUkj0EtuIbPKFspa9
5Xw6tY8BrF2O1u1dwVshOUb7H6rM1B3665J7e0MCB04YAoOwGCyatuxKvxr7xGQvjaCUmdU1d9/D
Aq7SwTr6zucxP5N4Ju1hzM5mp31NXmnp5iioGGDuwDBWUnEAh/PAyuiTTcg+KcaMyLrOdE1dycsU
R+R2wKIRKQ6e+2GCONI1iBlzDf7zuTZ7bJPu9nihyNkTwU3x9m8zwfCqw6iOu5fGzfxSIvR4q+f9
zu1wLjwluXvp6mUtJXUiDDpfjp1XFF9lIyTBbvHvSffV/QFije55gE2Z76B7kkFuomIyiT9yZKeD
l2PEFzBFtSwPHsrK93Kto2DBBIcWZ7UikKF0C2IMkstw9DSo2Hbb3P5U9FaezLtak1axBsf0XT/r
4Yj02YFVXCPZS1Qs3cBMpkMKJXR1so8smeSq1u0o3ObXDgdx9N1CP8b8eORIDlD96e8/RMmtBDzf
5kHriUATbHAJcwySq/4WaFmwJMmJScZRUdRMUQOfhpVpyaVcBadzyKwkMVX1Xxg16Aq0RFMzFFzg
ArWzuFm2JCAFWXFMpjnzCnJ6iaC0GQhu4OUubYGDRxlXIYfOci0fgvCnnJToqYZeB2hUs7GQErpG
Gto28pLK6iwPGV/HYWIA4mwIYHzmzdb86BfhuPsWmQcKCEor7ehvpZIGY9E/aK8eI+VZJIQFAoVE
ZmeSSRUC/BzbR3UL2345k2KMVSgPe/Z1hQQ6f++4iW0A4GN5jmsB3w7HnZtmHcgzZFPhUtsNwap1
BlNfye9c02kwTrkj6aNvox+8boht9WDy5+6Iks4/zsxrPsgQvvjvNW/hR8vqWgzqg7ySdMcrNX/Q
Pb5RpVQ5Vn7E9WtmtMUg9d939rtz3Or2sbh/zkPwice0TUoQwZSK6xMpVnT4UEAZW4UV4lA9+QUB
8qEFBQ+T2rrNm6gkh1CWOahMVMPldWOkLvcOy9ZSBadYevAO/+nKwWJ9Kyf0KvobFn0iIzFynZz6
usncKbXa5gpi8LNNq1AEAu7lP/wkusru+SqUmSzLKoA98bdD0WzTIDgENah7794N/kAslVIBrXU3
Wpib+RHUcpfBs4i6m7JJhzh6mKldX2vS3CZieWj/szxCXq9ABXQPIWZUR0tKB/tWQbWgUTVBRSBx
oqXOnj3k+X8xanZhe2724avinBfEW7ziw4DiTUYNn/8a8VEs4TpN/FoCjbXC9mBzTswHhnj9U2s7
PhSiefRs6KMXws+BxM95DcoHocOYfMeDwJfFmIDluIwnnIWDCq3ADczZhyjBIozEzXj+ca6SPUx8
OFjBMPROQKTYBH88Yj/+6314RCyF0nMoPUQ0CaP+0m+//dpmXz52NbAEQrmuyzpAk7Fk+QLhOqzv
v9F1OK5d8VZxLwOVKUtVHga00lYIIi5CdJIa+e82TMNSqOmRyY5RovZL8yeB0hOmKYsnobeUhpxa
i6mpBsbXSGX+VZ95Jwml8HlRyj2AoTfIeG7Znx30Om692zrAsMgoDBJs23e5Hu5WEe8pxijgMKWd
UTM7gZWFbkPI4y4AlrB6z55TfVYo7sSar69JbiZ1g8kdsqk7xebAXtYr3XDNvijICAvPuAwX87l/
6hwg4mT9ztfYsRTB7VCa39yaLV/3RbcL0mhJhBCfXWxWAczJ4/0A4ny9pnPk/dzQ8FwuAJZaqb6/
ddAtvYyeqKOuuRfsTjpRdG5WBZFMbHGP99XH/UVBulYRxB6C05alolVfTngp2qalXWJdvVQIBO7F
nHmHmZojHRqrV6s0i8cWu5x/7OuDe+fH2pmwrL08jaYgBDCj4vhyc6Te8MoX6/XQZJKqRCoNB3Af
EYJ7lrYPGg6RnNycoswiutn4CDcQCL9obUGAbJu82QGE8NskX37D6V8IcnsCfMDcLZdAA6U0k72g
ygw6cS6LLPl9BFU4mvLs0HglktMHLnx1QeGhVhvPanE4j4pJEzCYhHdDv0b9uJlDa6XQwNceB0hH
fTlfYXrhd8TlJ3jQl+KpztqcflXLIWDsTwWFJYPr8fGjd7hqFWXf81ziA21+bK9dgRheFEVETp1g
sztSkl9IrfVU5Hoeo0UTGFPYsWmlGoX/LtthyXa718goHh4Lpzznl/W64bRfD0dibB3K1oiFlQEs
FX4bssAEnk9fE7jQFnGwnuzrZnbVpNqb1cSKrCAhUC3OSiILqf9GXPOQRMMig8hIZDF+2vI/4RKd
EX0J3Ej26GESzMt9MjTGjPqlrPZ3y4d2WeIwmmuJHFHx09Xu4xubTEDiUtWGNKR4zBkpMecIDyUH
8e8uiBgAPltnLaj1LR16dFWUFrqBZLKylIUFMt/ZQ6yzggcIjERN9KJ3tV0U+UCShMkDBaghvAXk
IX4hKN/b1brs3l74bf+Y8GlmxzuG+vGdQ0JgnGQlfiWVJoAiKfUzPzwV19/YkfJgWYW4ROqx4D9Z
/O1aDhlTQwUkrw13TTtc0ZyV5X4TyhC1i4Sfdb6gd/DRpIvH08cCHrsnoAjCYJqFJVfLTn81EuNV
FhobVj0K4Q1Y4Xyayk80JR+jLdOC30pYp72ckLs0DoX545TPf0CvSB8Dhe0CcM0GpXjVtPSDqLBI
0ntZR0xG+GyufHILz5O7TKLCZb+oRq0VewKqatA7AAY99oDCPbY9Kx6MpSYQUyaH05GXVrjaVa+D
hGhEsOCF4/ffMi8sg2mFRKyYqlcZp2QMjeHpd9NlOgT3k+lnSQRuNhkv//QAnnwJ2PUJwktibuIt
atV4EU2mex8IfbSzomkN9BlTQNu6kP5b0K8Vgc0lIcjaDNuY+UvsQsJ9TNFO7RbCzGHQXPz5+Vt0
AsPZ1CCnXUoOBiHHZAPrmS32eG20RFoL/qtq2je4CflkynzzX+Bs5FgPiq63s7MUjCfEvn/OfZ7Q
rV3n8ceP3j779hAofNNuw7Z636INxfmEkjZa1nwWYXtk72EdnmjcTsdqKln1ZtjP+HGGaaub1ZcO
dQ/FmZnkTNidMUlCy/BlFH/PT/q/+tR2ggJYJ/DtMlgks2lOFZTrCQi3r3gFC8hY02hvn04E1LmS
sbUoqcLXj8LQweQDoUbfK30SW9NpklNho1vswepJdImPPif29sFeLbZOkwE5UINbrocsY151ZTBG
9cBpuVRK5p2A25ZB0CIKpuXgZrXbIg3icgv7XuVKhgfrALx7bU3F6xuPpN4Xs9Wu50JUuSmrbtaL
IyNBztlImun2Ladt63Wf8M1FEi0bqa9vIlhaN2QeuhzgiknCeg6i/jsJL4X2wgxHv8xgETQThPcG
6MXoeVMt3Lw8UZYtm1SdbU1WJ1nNgtSHXOlrYioWMRav47DsDEWWho+kIbJerL6mr7hrEKzaQT+1
bpZacA624nS0aa7pGHWMxWeRui306fIfFpMUImz20VnLoc7bK08lyU8cEtWWux8eQZtc+CPpvq1I
ie3FN3X/is+Z9vatIA5ZB/jtL86YME4TsHFTVDG9TeCCmpMQ/wOUv5c4hs7NyixWblXypW1EKdma
pYvRWBWtLJ9QH6/h9yaJpMshqhEd7ZfD+r2clzcQ+gvcrnF+IIcU02xILF5wxIKgZCsf0EmULSQz
fhSfp/AmPEHHdZx3O8G21yMaruicGjdd/2apDyYImAydasm8gxs9yokYldu5tj2Av+LZfufCWtJQ
PmV3KrnppffIKK3tN8FeHypwlu8G9Xs+8KGC+gGQA/l6iLDRyd6DQOdW5XyggEWzoTEwsMNeX7Ig
3gO9dC+3OXRuxWOA3dtzSCazHReN1Q3yztPgvTkB/6jN47Tj5fdFtX1vZ+bUw7vm6YIXy5Tx2b9l
PVOmihJpJW8mL8ZwiNj4SA1UDcYYWt9e7wUWd2jdzdFhC7bt3j3w/gFN03Xy1UimOaiFwTV8sKYL
RkAp43KHVGl6ELE5JUX4Bkw4KSBkcTWsfyeWvKuNZ4g2Wk3Mj9EoPQUx6KRnKoWnX1m/M2wjX6Av
SY3/pvUa3PMCKVSc0gIYlGbO2CDa+3e4YNnHcB4e7DJS10EWjw97EohnXjrOP0R5HEte4qO39xKj
PePmCVcnsh1BUzP923sjIv4WVnO84xlo9uTMVGyrrU0Ptoh6Z1rJrmmYklLn8DNFJUDMfOyuUHqm
Bn5DXyNfWBZ+TYHPP8uIFycwCodKgngz7HcNHo4NJTI8eV1xltbG+aUWpyykk2Qeix4llbGfwjC1
JFuB7T3M3bVfNzByFbIeyTHfZPHwWUDLN18vuZosoKZNEguhHA5mF6u0g3m9HLsQ8G7UFfQ8AggA
EoCY00KLgHz1SfWbOciWqHNmxyLuSA98qSBh/X5W1PVUskEZnLIrKBnK1jP7jmbnToQqsuaO/XUZ
KKCspIO/1EmVWZN2M/fSKc7RTafINbEU2qEBLgvG92xTR6LPZDVTO3XqVZ5XcgqTwr8WeF3hkJB6
s9q/6UY/evKMUDTEG4RdK6LtZVuTpofWp52ig9i+sHfSIlKNKHK+ji51UWIwnSwJteAUluxegkBy
zsp+HJ/TeUGxy3G4ZDTQqxU/nG9stVV2fNbI9MyZiz4L9j38st1MqrJegz2MLFtaJAwAYDcl+544
KqqaRK6iR5jszLVuc7idKRz1mLQnCdxLUgbDqaCZ2XdU8Blkgs88apXqdSPlyse5DDDBvKzJ1Dsk
84TysEOY1ZpCacOwPHWu6rntx1zcbVgmnJxnochdzGcmPL4Zjui9FYKliOjfHUbu+VrilvC0BVf6
BboA3vnRtb6Ulf8R+GJbWApmPpKl08MxT5rMrEjWSbIwWSRtHw1iotT47kpSm1nVr6XaZDp6vxNI
CETykxem1Y8Ya2cc7N6t1hgM1P8bb3ohxn/+u8SPymW7VIh0ciGV1cMEEHfzQKw0Aih6riNYsVYQ
FE6e0EUKJB6IfQ5o+l8WpGSzyQlRUwiavrg1XgOAmW4Mr9Ucaao4gz102tEopgDdFwzYrjKVOpaP
KJnnc6QN5Z17+WZNd17SLXViIY8N2KRyZCkgdUBHTUyngxv+zcFzxUt6eMuz4AX1O9zBP8ggcPIT
5tQpdbVKSb6hcJCpBg8RYrHmM8JjzomJExutbDUys0AeB95vQXbadsOOJmIRK+v6Z+hF17dLnhmg
dWlURauiIFaQN3fsxyIP2SNEkmQGj/C7SyRl5MSrm80UQyMlcfDOI9VhHoO2cYDqfgDN14Djd0R9
C1WMFyMhiWMaFtKQ/wees/D1Zk2SpZbjofcNHVJkytd8h2180TzFuwSSkTFhxF8B+vh7hwcJy73r
oEQxGCrukXz0IgW+AIPI2FNbFHUX4fvQmfiulfnWF88cKWiS/ldWhhNl4OjnaF1hXHcVqY5EmqFt
5n7JzueXjHc68rv/ljMSeahr/odXiJCZ7w03We17jB6sOw6IHb8pi65ulLUviX7t8s3UXqRIcv9j
/WujFW8eIJjmyb3Aiv31w9LnsNojV7OkygxRyEtkVg04MWIViHjCJDC/oXZ+tOVMIBUXitWGUiq7
v0lCbU4lrrjkfAoPbZIk6+8cifxtERrJNQ+c+IosIzSlKTR/r03z/N1S8+bCvMB8QD+rZi73buvB
Og66gicyVDR9SRf33EoMtUpLILW8OHZkaNbOqgaSzPxUIEfR+0D11s9DOYuyuLlD8KmTVRsIxWKY
fmTIFE5acrclNBEcKc6thZLbF0rPRGeyhU//KFaSI0Aeko5x0JMy2XETcd15GG7mWjxAEADyNXL5
P2x9lDantxjX/kRKBZS0HAkRtlOAm7IgezypE46TKESHf/u1h/EaEntAxZkQzifD4aVQSB6KiPTk
wNOblJYI9i9U2gI/snkkxSn/ZhzHZcunoyAPEGwD9tXGaR7c+WmzehOZJqJLCACgAyY0Nj0TRrtV
sjoTFUMLiYN2Kdn7fcnlbY0CjINiFncC6hd8LU9N3derku2qeivqHBbSTi0K54H5ek/7OB7Jf/CZ
saL4dpALpA/7BFHIeygx6Ln1BeeqEaOzwJwlpqo/1tSoa/WqzLFHumXQQSupDeDzS/PQQ+lCgdNU
j/QxodIPiBinl7VngbJPq9zp3fBhdvs7qQNu7lalRsDarnAxfHkYP3f3yCbDSPoF7R3Jb8O231F6
u4/qJ41oBAsPQJvwdTlAHdzzATuTRAcZWA4GLyoM26RLyazKQQRZumRbe3EYDWo55d1vDKd81t/X
ikWT+nJmXBYuU4aLc2OwZbSJDgM/Iodjqzb3zCgRslPcT7rJUxkwCBdlfAoPm0kGojSaVr7UITDg
YVPMNCU0YobQuuGfztwWevJWX3wGOr+8x7XFhCzVqVsNzMgkcVe+iIxKtejQX58SxMya2hbtTNOH
z2rbQVAl/iwFaFAYJV8Tc9NGA21yO0WmTGwX2r62rgPkVgbjHsQ5c+S0HBgSSoPAP95Ir33+D5JK
DkViVOxUYhH+Fz4jTXKL3528n8rQ9IhRgsC0/CgHP/OO4gejXNwfZfF/hD/nhfpBObL9T3tj7BRo
etc17SHYByoN9a+1heCfF99ln5hNwl/M+8GHk1EraBQhooxgYt/tkTXFRE9quqbVsmvOWIuob0PD
DWrr9BndexJMzquJxpu3k4SlC9D5nwwFLiNbuw7PMuAwGPk6de8a3hDV/WkLB3FNx51+4Nl7ozZX
gfPVFFDV1XpLJeYjk2RLV/7QYQDFqrCY8nY3jlDbOIwHCTzL23eebtK1zJQUtjPxloWXfCtft+A+
Gfkr2RvfY4Rk65F9JPBpAxianx0s7OH6t5QyO9mfDD5yjO5pcO6hckO/FNFryFyoC7KHNmrsaR5C
hVhsd/1T7+8zRUhwqWyW7vZ10t+3eGDOU5jtp6MhQa0BxK81ZvDqqJtla58ZHSlEpnVIpL2yoT4l
5B1HO3N7tgfftZR3+U5q1jn4alVQcnWVWjMZN+OZFc9utLCv6OomMWObnTjM9dUrnKMHw4akzqWT
9rW9638NYYGjCUWvW6gLl8kVXwHp+d9GN0OoAU4dsODN24QXDqHwOK1/OD4nPzkFqub4JaJcCanf
+4DRjbpvWWXbhYZSG2Z8i9jodQ1NHR8zHZlV5PfEu9RciGBmMHV2TSvAw7M2/RdomD9g18LHGPsc
wI8yuhbSMt3hlmDF6ntyZRenT0LVjvJ+cfkUq433sPycG08YdLoysflnmVGmb4vXqNYyI2OQPHgG
L2sW5sSYflTYs3yALCP1JSwxYEeBvYuMajV3FNY8rako30MP9mm/RGneulGRfvYDXcedVXwvc2K0
6K0n2lcg/PH6NOhjebQBnhsbo7CXF8JBau41YOeY0+SfFOqZ8kPhyWZzMq3om6/p1PU5IldXeECq
ZrBCpGxcmT9OEsL/rBx3yPYf5/1fqjOMO/2jYLr/9kBSR2ta0CmltKT36JBNAIcb/+RzAYMLKypR
RVKGDbNyoKisfzMSZz43IspsmcGzayYU9FU3ZBK/UcAxkPVAgIPUMCQXlR7dKb5ZlMN+/HQ4Uapq
WuzH+9SbOJ6uT28EE/c0Glzi0HUHS8//dw1DfrLD9m7sc9G+V5Yr+AgVcJJsNf4JLQhWVopszymM
6i56qpcKk/WzRMpOh1L1J8pz7S//k1z3s0n+aU7j4wLuLnx8CMWvFBqTJzpAHlp+IY00+WkfurVD
O1pDuXW64ZW79ovzelAwdtRMttiaTtuJTLWpDpds3UlaYEcOstYPMotktzDafG6FKF0eRX1ww4jM
I5r4c7GfIJZThMPIda2fq77sZRKmHvV5hJIA0iAAaT1Vnl/J0fItbehly5RVMhKtJmuBGEfKgrsM
dhwO6VnMdWXNmjLgGXruLzgHwBHnP2B7xN+K6N/ok/o4hquIWZTet3+iuttOijsV5gcQseUUT4FV
C+WegRkUnMljTk4j7BVkFyAMb2BAbvu2nkf28XzrJmcU10KGMv9ULKAtpy33TnGcRiUbv62TKTIs
GertQUXfod0IwBv+NiO91PLG4iDSKkM4Y6sskZrt+3/WzBtLvkwWmdW9n53uS/p83xMLuEW0HxMQ
tmoe/EWJUKRd4tF8eE3yx94M62dlksJ3RK5i2qieMsIkImMEORvE5Oi1jPaEqjespuG17tlV4AGO
3lM9ptfglzS8p8fAVh+yF0F7i0+80Z3D7wgUV0Eyt7YhQNHEevl5Qpdk1IYHeGm6tpFHTrOZWrss
vUrAP7lcG0tsyO2xFrpNS0J0tWBovTQJgCwXH1rBKd+vIEysDTtFEIbZCQspPexvFzEIV1MuviS8
vUHPlmTtAzN/siUwzoytp23rqqUtmik6LowPl5p/8kkWY/+//6qNPZnSj1Mtk7toVdCPA3/IJa0M
aaYgr4O2EouDBdv9Vsac9d6sRkZQB599j13wEq+oP36svp32kr1+bqp2h2NAcYvLOW/CPa2wJa8H
iaqwfQ/vm6DbdngY+IAmuE3fKa7AL9pqiJoqEa0vOsMzJi8nN+X5AHOZ2uCZhP/ab8wm060xWGcJ
S9/f1SZ2oYokRvfXAq/7wAFhPZDw2K+AmP/n5F5U2/NRUn4J/zgBWC9MzxpsQrktX/1H8h2WKkgC
OcdcQrzNJj6LYdQbsSVOlz9mKfZpCL07M4GhQsHny6ZgyPC1AymcMZ7VkdVmIVsjrK0ZtQnOn5Vy
oCpE/6u4YMeJ/CfnHOkRLR1V/8VImPGQZpQVszsn2xtI8/xNacMY6sr7bcOwahroOpKLetAAHGQw
2aG98PG0VgQxGX/L3+yDRcGstPSckkWmL9zjec1Rc23Ff2U0OpeVK8LuFtSRiStdeASuCaE+jqIh
4ifm8V2R6HFkZqqRuVPMsvM42p5DPNUoPXXeDXNx7zTraQgO0gbxA+kWxhgyh4d+5kqTtAHFwDs2
S3a+1xCXIboto/EiH/1mZDzqocm20p8qX3l9n6fRFPcb/OXFWRv53hM/POfNKB4DLuuapLw+KuV/
8RSpfC/SYI8Bek5Z67ymous8BI1R7gBMtN6Val471GIlJuPWE61i9QFjgEMKwC95W4z70Pckhb6Z
wY2bj4w92jfuod5CjJ+FNt6d3cocRYgAhry0Roo1ZqZTPOokU8FrDB8Q0QqZ8OEokMcIT/SiDIAd
4hEIK8WdEgZty/lGjJ1ZQV1N6trKoYsAxYU/oyZyRgy99QZu2Xnw+G2hS9zn5i/6j3oAB0DZLXQL
05tLfSbKDrtyidHmF6pHelm4m5Y9ohCdE2pB7C0OwUM53JlMYAEA4DYpDjfb8YbBpsiybjCMhg4z
kMYNVUbJVKielqn8YGpKAJN+CYj7svetxyBazp70b2f38VaY6yj9lZvkOi9kLQ3P+6t694w7Quro
7y6VtgQHYAi8iuHvPSZHeY8nuonE57yc6zc+n+DcAMu8ZfQ3/eDBDPsPGLo1RGN4fifP0GzvEjz+
foEFMxA+0K5vgLib7kKcnDUjVSwVQRWMAGChoVpL35cbXrN/A7ovL1eB8hWYwHqw7cHu/+/aK0Xz
ymTC7q8AusHiYiyV6TaZ1k1PwHO0SeG0RRzsyvDBQZn2UPtKFFLK05Z6JI4BPnMayY2pWWTAHhk5
/9MqGgS3lGT8H4fpXDXSib0o+bMfRnjKNXx3eLf7AcyBann+CzlI/jedOmNMX5/n2KaR0a+UatTY
0QTnKOxrZUUGbr43KmZ/R5apIzSe6PpJg5Hiv823FIS55h4KCIqXeV031FWWSdhcgpMxQXbr7KWL
IuY4L76XNlNXOXEMgGhu0vcegxGueCR8ok3wGVwGLM6PMSx3dyyJW/BE9RpkqsGWPPaz6w1F9cv1
XixUbE9B+9uYFXO5nK8VLqRt7IXcWW63m8xJ/A/+rlX5oN4PMhNbOHKeaxvFZgCiAOPS/BmfBhBa
60PigZIyCLYwFPXKZREm0OKrR6aQ7uR2t03OueZgQWoNHRKEJzdkmmnKWajEfVP7Ta4eG6Ox6MQy
54XEaCmy6UP3z5nP+KfRMNnovxjfH0nXQBk9b7X/11LfZ+mjCHVoUJmFCX9JeDzk/4hbf7m+0ZTa
yqLIrrWAzDkKD4yErpo+nfE7Zlo2AS3XxkarlRBn2Q+19nrctRy5VadyR4KLPGSIkpYx1VYvkJe8
LCS1ErKd1CsnG8Klan2wmzsium9xy3MHjVMaWToIVi/UZvTpENLqb4iuqsawAsSBrSAPmFJemYCT
w5XOevVSj+b3dJSW9j8WlgD6N9gZnRCFtyO7DltExKdpN7kxeFM9oC07xohZoK2t5T9/75lBww8N
EphMuGzkBSrmGr9/s8n1Rt8TduS5IrICwIor23jK2GkVl1VmXADDk5Jy5SeLh/1MyafxJG971QM3
CMMF7uDGzhMuQRtRUkmo3vtgR3uzNIwEwpq/tfwJ+mpSws8RwxQpcY8oxy+uL7VyJcTfVxujY85l
QIZ0jAwmHBoBpO9lgPjRA0xA1Sat7/hczXUwZyD2bomIZvFmiOXpzOiwD5AkkW4GK0g1jrPfau9k
cCnFdTcQlwB/6/Nh5HA7T7NEnq29lSm90eNC9PRgYBEjPX1b2NynxoLIPkoSe4EYJUJlbhxM0MNL
N/+ApeiIvzl0rmilkq73zC/Dfyfsr8Fxm2/saDTmxizZ3PfdLc7n/0xBy+aWbD3QUGvOke+e1Af9
IkioxPcqrW/BFvjsW0TGv1+OwAB5B7pLmxNvi0STXk+07ZOj46i0WL2IbGVYhAn/jdyrpQfaLBjI
6VkoedPwe1fQ/PjMxHeMu8Zo2oHnNqKy7umF8wg1z10X3QZU5ka2WImu3fUjMZQn5LRo91NVVFEE
bM5d2vxLFld36H5MpGiG/SUfjsjJW3/J0bthUhBerA2e4ZVwHtdTgOJ/UwhBEVSgLkI778XmHt+i
2FAVNLVIG4M9K9HCkj/NcjXZhLQ7gL2BZVp5aVFZi7RlecEpxypgQugE4Zsy4wZ3LJI95mcq8M8y
GARaEGwt+/S5XeAtEjT8XCI5REVew9fLP95N1wOUA7ah6aDmuH3njRusH5aMvy3/m6Cb7hAGzsvX
buAl1izeVj3YIDXc0nMxl2TZ4/DPFbqCdLU6IoL0ejydpQgtzFZbEeH9fLqJ+ceAYVUxLdf8gLQy
On9yuy6kBzBSxU4eXF6Z1n+nMvfMXgal+Mr/Ost8li3LtA9ug3lIc9nSa4GmynTkwCQSwBKeE0Gn
umTxXdu3GlFeFtZlgahQu0tHURNawXVXJtrZTm0fc/+ro9INikdoH/NBNOSmxzlOSYiCMUr0oIIx
3feXfqnzk6BJ/a1xidXdGMnlPEaHl1yMsUKJjUttNMp9Rmjnu8Oso+gm9mbZvBQsxjMMiPgxODdo
pbn8RCfkwH8bgvaqlY/tCFiLsJhKdVR7fBP77xyqAlcF+nRvJhnd2+CekDEkMtfS1z+7CRcu01JU
vVZW5uIEEzQDovctGm7MGgWAE5AdG1K84Xhu7n7zEhktgraNgMs7M26ONoNXUOOE5IkE4ayp9EA/
dAe6IGyfA9U5oTcWNNkMqWH5fKEAOqBvBCeesgVIlUW9F9y53ckm9UJBnewQodH3LHbY7n5JX0yO
toL13tawJbB63IRPpVGgq7h02S+QqKJKDuawp3eBPH47znpmxkzjoDe4p0qn9/Yg8sqOyT1W2PWe
4tgwqq7gbrQDxe83TnDW7w8oZaXJJFqiKjpGtOUKy35cKH8aWPXeNHgLZuuIpId0DEUw2SKxP2MW
FgAPa61gqUWPSs9InxhgUkgXO1fsZXRKnCXPArDz/TWl+C4odniyqjdSdNBDY0ztvlha/F/co+WE
bViPC2qq/H5PQjs40WCF+tn9QltPE89dgrZNBQJb6bFumajKpP47hkINP4L/uRh+xiU9X5KV63s+
0Y0pM+xj07JdKv4yWZgbucGwnH9lqnmZuyNnfVDmCD5WiSZyieHUlrThsPNqvIrBnDtm+BOpFhm7
NWhr0EyUrA+o5H5XKUxdjSgZC55kvRC1YMlz0rJGtig0m7ssEua2B6Fk8ypwYyDntdKZ7qhEZ1Oc
A2F7PMsxkEe+A9rblSsZ8zJ+OStXQNAv2UoQ0HGvJcxQ1tDaNIgYWbzNQDetcMwA89zCnvS1VVyU
Foj5obDRThhPyJHPGbClzUAOaoXUVq9muxjqJCp5SkSMjWsdmNS5EWGNXLTQffs0KM5ORvizPnk2
X9rGhCCYxYqtwG8HTo8BuN9ZmNixv5UlyzGtJoTD1830wsLoeQFmkqJ2Vq9fzMG09Ni/x9g4by8i
ZLe9jPRUirP5wlcaYsSdC3Ee/5FwTo45z/Qo0EsSaTR4GcoEwchDNua6vC0JXSu4ZDOmb0utHmBq
NsGuDrxXSy5CVCD4dLJDAo4vh3IonxOCi2l5sshpGKZLfDYenVDMWZwWA0iGPbSB3i4R13tkEggi
31qnPiXgn8z3QgQt+wrnkB+DdFZU0v6jMdVIpsIIz2XnhBFlZppKXTFONUhYt2+WgGgBqcg1qV/9
TvUpDnCa11UmuIuESCLVbdXuD+UCWrssuAcIKl0mKV7caEttyKPQL2mRN/B1VoBp51MuT+bddFp8
Xr5vI/xxvNS9OE9QXfSzqpBkrEg2JO68DqoyDk2pfZ2sKRfgA8wLusldmKmt2Mc9fIxRESmcCND+
yUqYb4W4Qhq0Lg0/KaHjcxoUygXkLa7xcrOIDoPPl4uFJ0zQsUpNpm08zxa/+8KmG0bD20aQGE1i
IVpBAmhjnjk5FW1+s7nDw+DZy2NDV1a05NEoUjLrwVoPRJZQdI2jKEcT9FHCZqw9XBoMZFQSVKxp
mS2XP9hlnkN1Iu57np8vCYb7dmEzjoZkehi4PmgQ1iHd0a8wNqLw+DSGdtiw6jQLKRVBAUJxwSm+
JLU/Nd2Aa5AZh9bE5Lc8RW7Fhb63FeSMp+17k3v12voIQ1HfxncJyQZpDCAvSDVE4DQgYIs8xhu2
/bz3HmLbRUdc4s7Wqb/zF+PX58lW7HLwysbo6aLLo9gESUOs4o7P34YnVUBUpRdCBSREpD5t0d5I
p//7PO75Ajurk5TWKhGHd9rfdQ0h8vvdm/cEivfNQpLUeLN8vc8uvEMKdM434a1exTLtJfaWuDfF
2Zhqhl63Le6AA6Pq922Vm8QgBM2/WG2YWe9aPs836v2eg3kDwsAMjhXbGn3ZVZcYSSzJPwqLf14J
L5I5ia4yY+Ob4bSCfTFTretAe6v9mcg2NXbXrqdxIPrh1Ncw/KAN0ht+lQ9/V8oJBmc7znbDcuZt
QXN2EN1yTa2Xf6wS/XstT9oAsoX1Q656mIGyEDUHEcu64DUU9VVYcQQjeKLIj92Pw7Mxg991csUA
DgBZ635TBsxPRH0TpCVG12aXi1Tq2VPFREsuht3TWcBCQAKZLDUjA1EtZpEFekodSU+AJ3nrAzVp
O5I9OKK8t24mLcemzeGDLyidgZ9nuhgYmoWpD9k4Dud1Gk6VddYlZtJQ9RopT7203ocMjbTcYCNP
/tcY83I+qWk0Vs8f35FmWTPN2xVimCvoIL0uzthqJvh4EaW0qOxFp15HzmRKGBTL+YZp46XoPAtO
6uE0qSS4zn5NB9BG0JmOXQEZPtGF0vpTpwJ2Un2dmvn0DcYYj+27r2PgOoLdqTQT3kljMlbZJAqy
A+X8VkDYkJBjCsibGcqkgB1sq1yio6tkMNAgr1mdK2nxZ9XNd+So7Umd2p2v2RBpDKX12cBpiZ6s
ERvhEejT7CiKPvLjDjL2Bm8gyM8V0n0V3rSzHArMgYQKXpq4VbxkvHQolICN2697jyKCeWd8IeBr
w408JF+Jo+10vGu58PVtREqZcKoZwC01sJh9GT+QxJzt1snr0QgfGAS6k0PTpvX7blxm7Py12+A4
OYpORm77z4k00hYJg5itwt+UuSt6o+HSx8KLXcFqgQJvX+39vvNRfgn47mHIFjOPGOcICYat3N3V
FxgClQuw2rKPnzyed33AM2bodeS8ES/qfPZYvb5TBvpUe2KisvV/Vaa5i0UuQJjTJrHEOKxdytwL
55j7CGwil5FXUNuMF8Qhy2hI++Ph9Iut2HEXJe58SbVadm22e1PcwzTr5/rrrEzXuZ3Q+0HUh+GW
bob8vbX2Ob6y3SXm4ke2A6QJVylMe8n8rZI9VVdnJcV1JRbojt5xE1SRLAw6jpaVo//ViHA6wZBw
qvzwSoYepAHpUyTCmPCMJeLUekNbbhtGvi2WeK0IwjWePTu9EHs//y1NwrkZBRXfEN/OPYa1yI0q
DyEo6bxEZQImKBYXfFGydEqpcYY6L7tDUnvCtty6cCIgetLa0DMmxx0CSXQkpBSO/3z2ZW1Txs3o
f1fPBWwGatYIzKxIuSfjeSBGNILOf6yvNj1IsQPb8efrwuXfBfh1c7qbApnI0vYtcS5Cw/+Ry2nR
fHgLz4HwZ7H9iez/xrhKeG7yN8FJ+eACvVORQei3/J0uRJPy4nyDTQLjGiFPeMpXqEv9fuiTf3zd
Ioh4LJF9V92avR2ja+s3mDypBjuAJVbr2iHWoCZ1TkL9yIHfW7YvaFCGdqkYbDqxaXS/l4g8rMxG
7zBAx6H3nVScqqido3Czugc6xvYDFq6FIQskIKoU/iu1lrv9ctq9sdOvtBOBTuKFBUIzYZrF9zJN
uiXrlWXJf9YlSuNE9OOyGz2tVCH4gpsLAlY4AhgSAEWmTeKM4VxVT+5wU3zqPz1QjEchfgWG4x6D
i3cvgc2E4iUJZJlrQE1XyrKEZMNgeoNiGWq4jqzrqX/mLi5Cu0MrVc0UsQ0WZi3qa4rWaddukdcu
jeXMrOtQCrXlN2AjoSLGVRRmms54oD+Le04EAr/7tAycH90XfFUbxnBfWcWkPhcJiFrEi3YUNOde
51vRTL5i4BzmbykRLDTRiWDQvWwBUPJsmJy7xeQXRPpaBDGaF9ZnpAy5lDHXb/IfahJzZNasTMIz
q8p0Mf929971S85XzRcIdtbZz37K+2MKARjnqfpdLzdzuat44f1090cICrCupD21ybfuJ3sjIqTX
Njr/MOx2BkwNsuYlOuwlqXLZl64c+lGFd/R2HlS0x7NjynSWGMr9AGDQVixinNt1PviB3e2d2rCX
6STr9qqw+b/hO9IWRlEVGo9/Ix4iVO7zR+eZDSEj/cs2JtZ9LwFoixEwarS8f/H7PU0ZgYhchfzh
0UOoI02UTNMYSvxDL/4LltqhpRmxcULHj7V6OIUePHhu23NauWREEUbCidHlRORRWyAf6xOXaDi2
coTQHXTIJLGN48lw8Ig2xzJx+8i5qyJQsNgc9m6fnScpHi8bAVhHUldpZc0+kfr9w1M4mkwjJb4z
a+5jJCrIOoLSnlrJThr+VdCfI7y7eFrH5qHUYeOi45w11ojOqAcdMqnCpnW6nfzGj48DHNt3s4CU
gsKI7uoWkCdMAuw5+09nnmLjw3/CXfWnFi2rq0MNZ6BTK8z11Nk0Ia6O87EfnfwgWuHAN8qU+nMq
KJXX3w2n4f8nUv3z5JLhafChzh5YiBAhlP3TutZQ3Wd2eK+kVyIf8hMNLRcHSf/j1T6BXxX1sAbO
cQrKL02CsKLdueuj5sYurJvzvvSV8aP9N03GbQjugOT7JFs73LwYmVtIqYj4viwPdptzOLM81w57
vJjdUIVvdKQyJFeQ7HhMO0JFaEmQjHUtn1UEkyBJ5w7DFs4+7iJ6mL8Zn1ZILDBYC1i9TVm7r8en
a6GZfFpP3C70GvAeZHE40qLtZ7tJLUm7wKqyQ0+tHBA05ApdYvm4H89Z4fOeh4LMk1VUF87tPC9n
t+DvALXO3sdeVA9VKasMx+mw4m2v2jXH//0M2lEtzmyRI9Aw5G+Jql+jULItwwUh7Ddh2TV8YHqY
q+VFsO5lru9pjxWo8ZGa/ROuXgBD0imwSk59KtWCTIG2WK432i3Bi5U1YLHd/6tnDFryCyNzpNxD
lH8cqLwo0LvRKn+iDYI2VAico1rd80SFhvIQo6CUv0BquqMSLCjoQNe7gCj4QSiCB50tujrWuQyU
oj4Tw6i/v+LI/xcj4r5w25FzeQYuEVAdIgABt+2JBsBOm2MxH+jLmucOF0y/JStXiKeQfjVWGX8J
DdcM86CS+PNHUaQt9zOYmN4AAfW8kRYFOyFN7KwtiLkVVYq/Q3S4YXJfw3z+q3sV+kT1jso8+7hx
JvBJL90yfRq2snnknsdkRlHl3Rfw08DfTqWpG7VGIMdc0iESM4WtoeW13F+dxfgjy4MWGK+DsiY7
cbSGR1w3z2/L5sHsOc54KZ2yuKO3U76zSOHb+zP2BBg5hUEpALwVmXmLw5pbPBpdmMvI/Y6i/OZI
as+i9JaCTY0xOrzHrlko2EyAfRH8dUhaW1lLsATC7YCL8IxSvf7/sTLOYUsOL/E1yG+TgxklWuSi
Dhdiu07Qq6x9z41VzHl5H/eVF+hVmWHkx5G5VjGzEPv5Y5zmCQsILxFGJHdENv+/5mEasAud0ros
phFg0sdZsfVSIdLX11ncAK9Tx7YeYEzYYE3k3LhG8FAVV8exaMmjxkGLKsuJVIVxKY8XXzDWXkUa
lIpaCRXPs4xjMpCX3E8vPJQtxaNu8aKIdEiE0YtXEmVudi0XgDYmGrQbBHTV0WAW1Aa9p0LHIV7j
tu9xM6iKyxY4jd1MLxa4aO1Q72p1HvJvSMDz0L5/l/jMOJd0bKV9acufxpWfuYgD9e/4qPIZ9UxM
sL1cJ+gqkWVxIuQcqvgh29iwtfRfJssBVrecrB6VWLhUABRiDEe+KmTEeDeVjlLYUmwbszYrkDUf
b+jAfIs8OVx/MpQL7b007ssJQ5vtGuBfyYPbbaAEfhOAPZJ+EVbdl4z0n4cR/DqEKg3cQOh4fW96
cBAFqi8EMsebIZW9VZI65T2TrkkMv4hzuOmEmWwLT+lDLUJM5wpI6DBLtPdGriZD/MC0Bp30itGa
57l/8a8bOOli7eOfLgzeITiyUBOQbfDwOFYeF9ybZLGlHo5Y8712liOgHNEMe9oOn+IrnzItUp1M
eWH1UTJKXuoaP2sNHX01Z6A/3/MZOmu5nQ5iKPQnXpdf89hDP6spK1ou01btUZdPNGffE3p5HeXr
TPraJkryy9m0xQQMxDr+aOcBIcnRV4kGZaT+P9wgxBeaaEQkL2CSEjiPPyBMhnBXL7itDXYL3cgY
t1xxW7ttBTFdicWEjUfEJ1sKWOf9N4Vt1IGErOV5rUvf2V+M7iFjRqGHgNwJEcqsMPdTXjl4/hF1
WQBpPEorCaVjcoHLTvlvL91pTL+1lVIPJVvl0zM0d2lXAyUE5ZMleS+MaRVZjF0mto7ptASyLT3R
Hxg0qR7n9JxKFjBp21CtLRBf8BiwxhKBaVr0ymjDKx+gL/DsLMKwvKdK3BSNPEBhLfVsr/aEmZYP
rzaeR0V6a4t1LTs+GCWZsrMmvLGDiwfalqivTnTfg8/kyEgumHqUkyHcktwQEswvnNx8ZM53FKbL
QEPTb6a2Th5gytQDb3ka0prsOo3Tt3dsjJ/Phv2qYRAx8Ea0RNUZPA8rRZmV4ZddVTjc92j/3eMT
Yq3HAqFk8lErlL2r2gZxkAFZABj7ioN7xVK39MG/V1xnaPCStksVLqg9YcAah8mT1utuo4Kxu0mJ
sLLzwch0Z406B91Vw8sPHcW8kaVS3PHVmQsJQKbrBYVIQVcuGyhWZTol7/mcoVi6GfTaVMZF27Mg
TihEKw61Da2tVkuNnLonLpMbib9vM+zWLLcNgXQTFYLxFfXe4J0uysDaVOZHP7UrktjpMM36DnUG
WXNLMgN4auEn9o0RNwSofSTBd0M1/5iynVqZPxHbEsOFVRupM1zb0zH6qMaG6beJ0ib2TknySezB
z+abojuOm88uX4pCBAvoVIA7xQZzOCeNbgF1aXngy54kIcyaEx1Moi5Kdat8T1Jd7Wdlm6IvkonE
sfvCW9YvdC7USHXbd1K3+8nnDdG51J33AS0M3LnlLsM13kPs4nj89zU0ap4f4HT8r/4nsQA6LKI6
PLwAz1WnLKSqFM9hxTpXNH+PS6c8YAkBl1Kg3moXoYRdBdOas7UxYRXsCILnYxS1LeVO4JZf0LSA
uRr3l4J2C5djkkCMzZcqKPCB92ZjT7R8f9dLRbdKVSYXRL9XSPL4CqCjN11xGBgck6ByelBJTwuY
t7c7F1h5ziBmdtmYc9uNqaq5kcVW+8HbmXWQCMbLON75BiyFuK2sk7LkKtoWxdYlqwx59Sq5qOuF
O4L2/Upxt9hDWR/8f+hjy59ewSOlO083XMluukxItT7fjXKAnbzrJVXm3fBYo42PT1kI0z+Fz1AA
6Gw8bytROMPPGlDQ93FaGnT1GWJ/dbNLoPTi7lbfYGGs4js2KDkWEbegZNgCeXiAQzuGsLSNrs4O
7VOoRmjsE77T6orCKr3AmZdxiawW6YMOOxwh6ShikJ16r2PiGNLDPaeRvdYQRM+gP9QK1NRYPJxE
NQ8h+9zMs1duXAgublrahq0CnGqaVC8yWWP8SK/RT79Aa1sQopEI+TSK9WBToRWAwWc6D3+OBFxr
Zx10p689i4CwbG67/cV+XZygiTGpvbbq/BLclEq8WFAx/tvUxPJj4G9qUJSZEXa2w5Nr4/6haVGM
8xbrLSZiwceBG9CgR0S0ytj1nuh4fBuDcL9vnsx3aZqmImx/yd2/xg0UN4XRFq8X43qXRJM47sRi
bK26rRMosPmICFVoWfA0P1IZDQxOjGo08lvUVbdSFAF90a3Z4JRRAmAnl+47aZ85Tt2/BhSTaSI3
vSlDHhTqENcpz4j6EATp+P5jDx5zuA2Dx/1VkSVZgCmzUTnNBYJ9UKEOgpTsUDuWpOtQTopuq+BZ
a8E5Pz4BI82c+EamtTN1t+Bd13ta2J9n+WWAWSgFN65b3Qy9sH5GBmAlLN8YwQEaLu7tzdCkX/h9
d7XpKzgO8tirMhZG+8rA1qyVbZRC5l6PvscAa5yevDf7BIYd4zR38Ne5diNyVhlDHcyz7pYa52HS
H+XMHRdht0dYvovsE95QF7ZRWnDt99v27SLMdDM5lFZEU5LBILl+rCc9ac879GlsJaq68/omqx8s
3eoIi1/IgcoQx785NHWCQekSiiq2DHN5Y5ayggYRwB9R1oKF2ZUrMZPLWiksJscMNY08/BOxK95k
jbgmPSIvC+ErlYgXN2bsfh9/HTtZW6mlO8AmX/23kGIAjG05JVb3ZrV+kbXucLDewb3gM/M0Tp7b
fwMXu+KvaeT785hb1+za1Z1PQvhN84qZDMEScSerELdSmG0SyaD5pu9yasa2kPsSfQumQ2RznGhK
56pneS3R5ukasVGG66ARbPNmZ3uNSQEYaXlmNwf81lWRX+kW3e/hWH6hld9ar/AQxrpx6+cy24Vh
Gg3UYuuRWMmfNzpeCzGpsCMZxmwKv7j25iLBOFeVBO4yFiEHaTtKsXLGi9DjiIj6MNv2kp7BRn0h
o3QMQPgh/BBHYnbNwBfuHJIwtYdvp+nYjENhIPpoWQRRkXZsfTzlINou5b+CsTwrzBY/C1y+Ex+i
cvroaoe/NulNj3+bKWoyh11qDaiTtyHcTef7BXazRjHYLiCpPS0r79zrhZZqH4L39wUdnjD8EXgm
Ggiq/G6/q3qkoT06NahgJ3LMEYhnzuAfUrgq9mkjiGwcufevCGfQzzQiE5LPDEG3Ibafrv9bawPx
hjGHSMVxaSseEvsFDxyGh8rKGkmzDuzUAE9iQoZCUBqp5pY0Dw78TpO6PlK+qfdV1KSVS4XHybbS
DECsQVRWGvT20Fhg90VvJtMNgV6JHUkxMKb59Saf/k0Bd2lAGCD3amJc3UXVREFlJotFSPuFShap
d4z/s4LplIOS8RFt2ICD/yeChWpvYekscyWLxKTsTagt6H8hwx3i9egWon4smqbCIcjRDMILWbAr
ACUGee9GO2p/DFdSNOU7dJ5lpLCJoCA3rwAuVa174emjN9sQ8V1NrttsHYHs+IiCY4V19RJDGus+
Rm26vOJtHm3T4ubtMc47yMcLh8UpaYZ0IqsyXh9QgFzEGp/LkWUY2JY9lgmA62Q1zLbreqCfCWtE
B6XleIra5Ly4Q093jsVUaJpdsxkxx0qiwKv9SFNXRx8o3pSdOLHQ+lhXf0F0qvRc48tcwavtBwgI
j6vTE/sZ7v513BZHmrNZHz2+m2eC4Wvr0vWDkT9qvMVZSlUzYHg/1HMM/Ca0tZ5a7cJicvwz5HNa
1eyI49jttyCnWuhDS+d7QuLXSnzn8/zCccW7VJUEJRQ1DiU5B5pLgaMW7Wt5pqWMQp+9pphR1AnV
ShS8/Xj05tVR6aQQv8byFukYRFkIusIjXCXEAXF1IAWYPNcuCO8KNLEvGYFkwD8ed3Dq9txwCNL0
Zzt4QpTOo/RPUycNnumoq72glAlVeVmKfyu3CdcpXBgbGNS3HPI8n5U5ie/9r8zAHQjzRhgSG89d
E0AG01SIQiqlqMgnR39t8wNjNuq13bqVPh6AXCMoKniAGYgF0BrhCBxgRNg8w71SfttCp9TZaIve
eSPwZ3Y73HLOCCY1Gg46y+E/ofeEQvpTJsVVCKAcBo5+ieo2ahDhtpj8XUZhOccKIURL/+O+Ht5h
lBM30ecV+Kbi0rZWLaGSjwolDdBCZNYzTS17w5ttZjbV8e9EWHnqkuOwTYM38QTG2KemXAo9n2Wg
VB/0P/E5HvLv5Od/b/EV9U8FyWn/w0C0sNY/0t/zl1ah1POrQx9meYI+QDBTGUqit9TPFpL6k2dF
7TXC48Zo8YLtp6gbo52rf0L8xSDLY4uMuCAZTvidVKB81OLfBbwDd9aHzcsso1Rpj1uLEz+qIYP+
TSAAjOg9iTp2cYr6+CYOJtEkaOFQNPA7J++lLRmIDYES8vCCAnBpnKYXqCpig1MZS/KLq/MbZoHc
91Ypt4UxTM/giH475u2E6TvaletNSTVYdK2Q8Qqmiv0uLs7At0o6w75FxriaiAMUUkNY8Uoo5g4p
p2b4GMXXzDW+6KIjOJ/G1TcvkuDWgASteftjzX110zfUr4AShMWVZWfKho3/tyH7Wcc42BGlo0qR
rmxfdInOcM7c5vrK3AdUAx5zTe4II3xRRf7HRFMo4tM8F9VUr50XXWsmhBjNsIkFehKVJ/jsYZGE
SdE2OoBewo8AzjFzPQ6jxCtup0zOyGQzC/GXHO5/Y3vqP0r8cxdF0HvjTAmk8K9VufILT2Y7y+TC
hbkuVNOf1i0fWhZ8st6O2W+/Z8e6U97psoTFp6B15+/eiN+xK721NGnR+H7AvbfnzOzLfalQ+NgK
LDMNgYVh5ZIcmE+YYbN66tCNzOEWDunXK0DJ29R70rQ6FHdI1trcvdpaoR2g/ZJZCqm20C2RvcVk
SJ7IY6SoYNW8E5dmBx6dRMgyXlbnYMbAY9xflmTX0Rdz/KzOF+Uj9CJSFdEX5BiDRwX/SE+IBawD
QpQZvgrqEXoiov2twKchbnDtFyAYBZ0SgF4XuXcO7cK290JCOTTAqPOr9gbYR3gpSsA0tP1/fqnH
ibPGZ3jJ81oukujYtM2S+NKiMu8TTGs9oZx0zz25Q0vQOnOLhar/aYU/yr6l+z58who/Pp4RmY0H
WE36JVkNneD1q/fwW7bk4p86vq4WZXu/t7ZMpxkheumzFXUbh4VMySct1QSAOzd5Y9WRCrrqiGIC
5vbW/ctBFrcAJgMUdm/GjA67dkCPGKOEzj1938lkgQiijlCI8Pkgr2vAbLRIama543A7I/pZoahr
eW1wI0YGgvkClMopo/YTbNbqCDCgWVcZqd1Cz752YHAMzQj6liLav//tPSDUdIWpPW9sqGwN43Lc
fqbbykny5BhMUfSpevYD8y+sRdgGzAs//S1xltjaDJ9y6FTjZxy0j/i7Twn2zVAoz6n01zhS7o/C
8AoKRm0eJ4SmN8NS8zntsP0QW6837D7QlZ0K45XEMS9jSXbPw7y9LhY0v7C1EvZJEwUVjw50zEw4
zf8ZtE5pZu5loBKRp/AOShmREEXSTVf7JTB6Dhbf5KYKdQd9QLrMqopOr6A62RHbBLtvd/KnFY5p
GB8T3LgSQxJuZLnUwZt7ONC3lyb40OdEfI+Cqo25m9+nygl2PJQ3zlAosO29sbaXk8dMd2FF7UY5
wsnRVedUNzSBsZb3wVy+21rWQ/gDXelH26Hkt6bd1aV/L//KNFdmjtfWLUvoYw7m6W5+b73NQzal
Al7p7jR+fBWn11raJYqhdkG6jf7/iAmqQxTsKPlY4hxAalMPaL5fphNTXYqoxq1/cBoClOkkGNcP
74ZE5y6d0EuLIyYkKg+aMshEuZlX4TO4xOMK6V7IubFmKN3pqrDUSoMB0MMHDvRnEJ0LuFJ0dIbu
xmZ/NZJynF1AGsVeVl1f43Nc/OULm4S04Z5t234vNf5mMSLtBlVIY5fvIFBPhklD8FappMvY+Kx3
hJfZaRrERo1NE6RAEkb45yWUP6mQYzYlgB38mIosSTvlG2WfJ0HKFoCprOrUn9Ovt3JjUnpGG0RI
pubYrz699WYLauJ+WxMtaiLvEFdsEy46j+YNnMqjI92Bs9bGIfw7F9A4KZDb75y83LAfrj9in3qA
ZaTwnfwNAM9PuVrPhXPkeEH48s236f0iA8OEKveJrh8Ki0qal4ZYwQ8XDfof2NDHBBnJ6jw3iU/F
JYzwyx07orJ82uLeiNewuvQVHlSzi2Jqk2UoJhIp4BitNTZbgBdm1QodTru9Gmo8l44SAmmMgFua
2M2DhfrP9rlaHoNOaBaOB017t5+5SZDf7pMaIi4osfBhzc9GMmWdJ7ReIgUuBic6sA66etYif41I
mPqHxehuoBlcLL/PbbThjjG6fl2UVbNQjr3ANnSOYdP9Cf88lNN/IDTtT+rvcrCfTIQt1vV9MyN4
l7vPmLBcXIWNW7IFOjJv1qI4ESggo/KSJd7tzP/nd5q1uSpOnh1giJyFSyP9w3EcgvJm3kVOGBJv
1JOGhcsn0P/tsNvlZo8JdAPaLIMr0L2hHBCGXwVUBIpKbv2LtMC+vBVL4FVvWtsAAvkmOi3HbOgR
yyM92dm2WO0tKTAb5GvJsWSEMyCUHvNc/0OvXSnuSJylk+Wi9IuEB6o7M47U98nYJbFn5WhXpmqI
WUPczoKFuWQTQGhYdQILvyrdJzmApb0C4I5etIZL3RgNehOeXSuIZ1ueYErnVE5k9uSQatZ247U5
h2IXFdf3tJmZiuCOQcULyZBE2rAARWID6zzKeCFDF1nVK8OdVAKKlz0nMk61u/pMMBJHO8y4acFF
5uT0J84gNVLhElxpqu315xdJv9sGA4nHgAidai9OJKU6HnByu0fwfIeDgOu9Of6jfcSt3ttgJTiT
jyX9dykuvr4WXMWvEHsqmYb1pRVuUdv8OrRw2W+V3h5t1OEZTIGTPcZgU5TaJ60IqlkhSsZTzHdC
gmcQKbe0aQomVyBlyj2eamHciZV3SrPTuYGd+rRiS7jS4kT+pov4XZ13wTlzzZAH+ARvQSJgH6Me
SlW0CITlvKbWJ8ulED2SvQhJFZrG41ZO1u7Bd6T98tHrMcnaFtXO5mWE8B5jMHAppUBuWIQUCdmh
EiIFUOqao7AYMtGQ5PnN85BsK5hKmZ4+F/Yg7frVQgmDNh5g+V8THe3n1L5PgrqfJkVpBaiJu8Di
KdB89prqYxETd4o1poXwqU8YPj+TRFLiDfBeaHZxENJD9OeT41wFoJMM4l6qcZJnuIapdmYyvq5u
bsbMgCyVXzGTytZFk6NPKdncB+ohrTWKUEkquvn0T/gcinIM0DSjy2+j2peVdP2danorNuk/tKnB
p+KvYsVaByCT3noMOE3YLRTD3KY8NMXW6Cs2ln/eXT0gmk27NEKgq4/qVoSEXBrAM7GvF3ox6WQ0
Lz2WF93TTKkVomkW2F7RemlfdYG5pgJ61LwXmveGV86pjGiC9M11J+Tt4EKBE2vt3+tDLcI6ChZE
sWbuVM1oyEj8yxY0UIP5JK4n9haQPMesPfmOZQXOL5nwygUnAXdHt6V0rMuJOVU57E4i2e4mqkMS
qOu+uD8N4l3b8sbtOWCctifFrmhYSNJ8cF5+2ISDq5YgjhTa0m2bopv+4pmK/4lO63oXkioCHPWh
kzIqRLmIwkmb+uDPKPHlFkT2blRqg2YVmY4Ak/8fEZm2zm1BFhNGbKDbBNa8LHibfTpp1SvrufVJ
wDYHH6idh3Y35BBckhsPwW7IvFjYY+eobrevGuzIPEeeAEeYv1yi85Sqn0PX/CxJEl4kN8+/Fz+A
M0AfYsVsqUKmk7HuhXZJXZ0oQ0Z/LcJuOPSSXMJCIcOxKSJAntdaqLlwv/Bk113mWmgrlgF9mKFL
sfyeYFhUL8ZsaaJRO7vpKtDpoVOvvNurplmsF2QIExh73jjEJlFa6cL9/FQALmOSb4E/ll1p7z7S
ruQfvQlAWu/DbIZbfx767kM/tfl7L9L0NX95fc/qHotFM0qHqdioBM7OgILO/TKZjpI1tyLrKQCo
WUFSfic23tP0U7/hlVuNxSonLZe4SVwAzPfhI9YBPnB8q9iBW5kqaE1LW/KxhB/jEUhDbd5nOaIz
7gY0nZdaM+SaLXxLkexF0+DTeASTB/aojj2aoUy4rceL3k+4n/xdPPzspMz5MRqlaW9KFKC2oJQ9
MVgY8gACMw5hMtYM7H/Ta6kxEPAHGtylwHTY8U0bhaFaqrcvalRyBs6gUHhFznH5lEc/Ob0i+d3W
FuaNe1jkw60EAr/1Ge6GBERhY1pwsxs0TtMJaxQNGkLwrtMU2RCkeACwoNJRY0kZgz/gLIZw/UIi
8EbewmdPaIRZKdRiVjzj1Q+hZNpcxwVUCjK3NayiEJ2hqQjHAzZd+CaDqj2Zi4oEc9ZeMMBMmpww
fZltmlAt1poAjg4S+MdBjyNMvVxPc2qlRX/1+azRuywrOHkvBfnv6ojgk2G69uCH/v4jqxqZY9B4
YlASplYI4ixQAH6oTJ6mUtieutEubGi1bJNkRfEnYciwxu0BVERX0YfmRZDh4T3VQDJlGawY0byC
Lw7rXSpRdEabE6wmAe4LrzTTqTKlxBWBxrvo3UpM1Ffaegegpi7NgRCtJUXSr5k0RWqU70l/c1rt
dJBNl8ZlGzPbUUWNjunhTPU0zBdZ4ri/jX687bxCwYcuUBXuLGeF/aEEFRcBZ26E5dj/7ZSj8Dg6
SxqqL8o/59IbYX65VqmfnYBr6VPc5KMb8QXEFoq2PBy9jB0KxP4IYwM/MP7MgHXwF7JCN/rAWelu
ZVS8C3tNLg03tN269JoMgkABZhdSIuOOUZTYM+1jRbYQz/HgIwysHqvawD9PysE8LPb/8mlPJdV/
ch+CxSiWsaa34LfiZvSf444yuHK3RAmr14F2ILjmazn1i9Y4sBuXBjVi83p4RA5A1p58LnfIp1oB
iYDP9hXRfV7tDn89j6ngxZF1juWFarxs4w2bDnyMESREeYhYIvUlTs1L7oAv6fgatyQ51aem6ddi
tQiGWA9jiSJTtt4TjZV2ZUfzQILowdoOL+/ERjbraFrZ7Cy4s6UwLagpJPF/Ml4q4Cq95F23Mml5
AVY0NtJoVLv+MDK8QDnrTV8luc5uNXQ/heCykpsY0Xumwzl/Kvs4W8ah9xspW+9Sib0aZembeDnp
ChxktdJSib2rxLZauphB7m5/VPRt8Rp2H0hC9WPfXpso5MiBcJnLybUQqnU+2V0f9N2gXcZcVlLo
4ng9aQQA8YU9ODhooZvEUX0KDTZqPuQtWfkvHDeGBLV6qYyDl9+3DwEOGmCF0ON0oaHBd532prc9
8OFQM6V30htr2BPdzV3QV7OrNq5N2ODSGMcD7lPzCv3xo8rAB/J3Jgh/zJ3AcVHJQC8Z/SqkydYm
cMtjF9Aw2QrjTiMGVIbKabWk5iD+TRHQFr3wiwVT4q1bDUvdh2cb4Eq1o1VUv1K7IWiHJDSfqyXZ
pVXU9W0x9JuXl28R2fjnoMJrV8Y8LQh+71TwS9+/bL2v3C7gAe1N2HcJ8jwu+9pCXc/eeh6tDKj7
lc3nENj0AirMNIV41xBcxlEwC/BoCMondVcaM5PNPxrmH8PR0P2nauw8JKckmjwFR9Uz+mc4sVJ+
G6pPQ0zGqLgprGsN6t/bvsUwzi+flMJr1gzjoavPSviaJwFMUNOqpgwednqgwYbUSYpXP0CJ4Ixm
fQu7Ajikzsv9XodQXB/fWXEuQu+TXBZwT3DlpQaHqs60y3uhjNPxTJxuSMt3+cxFrNpPrwFrDqD8
JVhcjfwV3a6Mn2TWBvWFP8SkunwqwzBcs97YWK60aieHYUVfvzIlVTI65DtChCwJq2gfmNwHW0QL
qex1db5cHU36wA4OYYf2FgdUwtaD8aph9iuge1FsoLaahgN5vZKimKV7l9K7y4oFKl73NLg3RtNN
rZ5bPA==
`protect end_protected

