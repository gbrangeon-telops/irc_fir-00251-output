

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YqipQWc4JFBZb16rc2dodhguFDkilKhXXsYOnDVSNRAjtkaR6AZEesZX9P31kdm98GkKMNT69IgM
oU3B8PoxIg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Th08Wi4CTujjzYeFPRrbrk96/H9lqJHT1fOXWDhDkZaqyMx5/LmUZnPHzc9Mi1qiTcgVKZeTpkDd
lm04xNkvaFBlZ5KAxEqjMNmhtMTNyj98wbYe1WGtUEppm4URdSaGhgzD2gvskrJEfU0HoVjNKsYv
Y8g1ek6gYioQSqVo4Vk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3ST6h9XhpdCHj0//nno4AUPlABBr9tQ0cisrrim6ayZf3P6t8TzMqSxgV/q0TD5pBIm//qvgm7Bo
W2S1EUuvf2WqWkW7p/E9CPizeTTEZkAYHckCfZTDk/HTJdolSIFeCHjfZiRizq3RlOIw44CUEMSg
PXhJE4sbT53L+d0eIaNmJBJnZPN29vIw8LbE7t+Y1oivoLSh1BhWy3+lZNV30PrceJFjB3Ylx53O
r9RULlN7k4FVXKoCkEg9NcpjWNJAX4azHw+uuE/ZZmEDfyzXMbaQPIzErM+LylAQ/PYfvIwSeBK1
4Z1Yudv71r62qTHPKAu2JCMEmzvKCe8RAmGoeg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iNgef8JJ0zz53Cg6UsIY3rdr+PhJG3ZSgPvV55cmHG2d6Sfxzk8LG8+nTrPNPEPV7qefhOfs2qwO
LV1XGy8/zcDatxxl7RZSBTwjwXvbpgbJIb3oKBLjSbNQOSIIh7oK15z/NbQ04jpEoFW8I8unz0Dr
X8lH8UO/ss4o3sjSRmY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gdQRq0TszGQ1sYR2djmFoWhyazt+0Tw2kvNbiTEjaM08h64rXWx+KrfH4Ux19p4jnBVjDnfhSE44
xN7ehFd8XzCnm6T9eZgkCDf8dP3IGf2Nl73ZHXLjDsXHqpK6BXZEG/Ko8+LkLz9nw7Snn2cWezi5
seVqFQ9T1Cl73kL7otmtLUuX7sR7LkwbgtAzFivUF8Ml8V/izjdNdzsqpzxjHY9vo/n9JWZSxDHg
dF+BgQSeU0ooY6vwulhfUyi8hYLdbvSFz9Xlr9vUXABI71kCIOeJMQA6BrcWbYjoGqM7KNL6TTGp
K4Gc5G7xM4ucj70Vz377eDl1W3KXvVQRmQSA0w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6928)
`protect data_block
wgy1MJnDEVt282kEapjtmeOr3CapRJSquI+320AA2PFxsstf4B3Zpc0mKKIv/s9hltF4V9KlAM+b
J7IA5bDuh5KGfzBTLkXxotSSHH7NvSJjUTv4KE911I+9bafetS8MEzKEeX3m9HMGjVAcT+5zxDvT
FBUR27mcrqOnEjWnWRpUfpKu9rAZcp/mkPTq9IpNyeGagf3cTiL6pHPXGFcRe4uFZG/yEhVbQb8m
8Ngo0ITW8L7b3NqqADkQzKG4mx4wE1xtYXzN+u5sagunOk4tzVS+z3eQOfE1xX3FZVhLD0O+a4Bf
BAksIL7DF2FeqrAxbOBUO62nzC+oOH2vsaPfHr8Gto8yviuwTMpGOYtl0GyhX+Z8J2isFpwkoZbm
oQYsxJcAfZ3RMsUGZ8aPCN0JbypOScyqBITeXwISQm7UzDcqmEkQRJbVDo0o3k6MNsrZmez/rYE6
uKNPUuJ0Ice4vojru/0ztuavU2ZvquXO6CVPTTeZlZzY3YxMYWBTJmtiWhvacdvKurfWcXsUoBZi
zMHsVlOlKNtpsuzdETy09mgx/l6j945QwF8tOONzjhghAT13ZnWGZgJ3I0cUJagsx1ZfAO2FXiDl
LURCVGF5Ajq0CziKHg/SXZ2KKsdeb+brYI/rtjjnObjL3h4p0UwpM/sl/brG8GsJY5pMrKr+2tpG
3MHITkDDuq2P4fHcPDS19rZB8wT9Du7MJ1mVEawjA8fdbbMOM86u2hCgGfXVlEjFa9/DoTglIgIu
U2dq+WkY3YMBwR76W/nchSLKPBTayJ673LaISGIC0B7d8JkXwj5cIcUkrpVcO8DWbfwHbcu1oZk/
vqCbrokoPowKdl58uvRKMz64Zn0u2ySQMJ20+nskEHpT5VMoLInvdE7YiEpzQ0TzukRIcfc53vlo
KFD6c8dyEcUfRfC1Pufcz3rDGU9Rm1YOUbaIF6D6aG2Q95qsuN+F5DqE8/54IebktMhzB/I6uo6U
6a2JrJxem3dNGrnOR9f4PQtxBKRedsMdZQ9NVOZZ7jQkiyJz7+DtqY6XO7+sFlysWpkZf8Iktxzt
+nP2Mh4CqSd/nPDa05q32yqAXFMwFbYLoVDlyO7CK/3LG+SGtgkUsF4pRaumO0t4R/6aby8Fhl7A
c8WZUB8OnfwucG1cKu+dnv9MWfRHzIvzUcwhI/KT0qH/BBeM+k4+8qJf8Qj8e4FptapzdBDpPXRO
nUXA+JXt7R1M+PC+cMHShbxx4rMiduPYVueZOKOIro/RZlEFeKszhSwf4aj5YIaH4c5lN+YQMIOh
ks6JkVnjxw4SdxB5z/fzBfYjKNYhNZM7BGxCDKtlHRrXZhKs8PfRKSiBeGDTOIwvaHtu0+7StewI
6ZWBVQVsP7eiziHfEVzLv/MEYvFx5YyczJcL3zVYma+lEu9+hwpKNcZfPq4Ix2hVYYBylJFLRKmt
+6opT+Ebb+x76JR+cUM1J2fD2ecv6MtTKyEjluMeeV75zNVztiAxELbi9/2x6OtqDQ0KrCU0h4E+
5368upnVmUU29tlTmj8Ja2y3IP6EashVAAftVGNU2WoBM3yMSGBYIJ6OuxQS4iKYiI1AJ1SMkK3l
Gz3Pail3pV9qTiPNm7C/9b3S0BHBZkqDnfj/NhQCgVhrH+JwdVEdAJDZ+wnQ47BsqVW4uZLWx+X6
/IkI7h0IA3CluEdZoXaQ2bXpnTkYAGPxGSwD+4L0ec/b5Zk7Zp8XZSIuqaLqKjFvvk5bwDeTi7Wg
D2nOHpyOg8cgIBJNrxsvub8ZSFQgxd0WgHDiAFGTIR680uJXDAyKkaztt+PeLhdfqrLOgBrOhcb7
BKIkOe+R/Aui8F23uf4/FpZGVgrU8cOKUH6GbS0yrJvVK213YZUctFgIBBaTBJWiKgwvC69PgUjo
zG++95gvugN9kTo9uG2bFaQ5oXXsRmPP3WPX1KgYcnbK5ebhhJx/Vi17CmBUuAowgSI53F+LWpju
NNcp1XjWWvUuR9VSy//5/6DEMDLsZ8hMJ7cxpQgpPbIff7KvvAi42Mh7TxPqbEuFbdzLFI2nFUPD
IB8m1ZYuiKSg/jGA7ACi/U3rmkYhAWIic9NA7CFqo0aVwQUnouKVRDCnGvznoBtpIc6Goha8mao0
IdybMpVO6oH2d885RPnyUbhxTWnxz3LSwvN7EdiqeauVn9lTHWBYmSi5SYRSh0O2Fgoniuae+Zww
O2f2XZhgy4E0FH3nOhUAPUMj+OtZpGylQoynPuwarWFXLCVZpyUrpukefNb39fhxXIYLwSCEOGtq
qkpqubhlXrFsSHF1stMjNCx4iLRNCunyWT8sGxTDX4TfbABcu8g6uWT9Wdc/A8e4ihMYaV4+CXIn
STegwCCCuJEZO/aItV8wRNJfVhMV2q0Z2Cc/avLVcq/P6KWu5cn52u3qD+4ZIPevjpojVByDk9uH
Irvfx55k8NHGUBXtUpCN3omQ4FhZt41iEwFt2LT/wsI7lPoQhXaPExVaSpXVCar8DbJdtGR+QI7c
dm8oPbWYTR9Tpsj2GKnWjJYTOjyNbo5Ckc+PSVuqf2CGYY977PU1HQBvIPE4+wPK2fyH0lmR5zlq
ucdwTK83S+NaR6SX5JWTMXlfQUsL6aQhwEpN3bSuIaczy/1JtlWY2ttoJtXbgkVAcu9FzD++h4Kp
thkUmbbBx2j2KrEwl6o2orXMXNNOCBSI4NsQOfqj1kDQWFDSqjluY5xTn/F9Psar6KRNorrSX/kk
uYo0knTJ9fJHuP52wPluEoFJq0jrQf08pB927XPKCIyTp2DIlla/ltlTjgWP4qunFHVTGE/bdgLX
uaWIe7JvNuFW224/j1P9XQrHPUWCQaAPRzxCmZL+eTnIJr6KDsNh0arSQyEMfVs/xn7I7KwsBD4N
cd++paPL7t2TrPZrQwK+Mge9pNj4Y2eTh/feAZRA28KcLz073Dou50amRbi2t23OMRXT6AYExgje
nq0B5gOlkVEz7slil5qqBoCCU+5ddAwieChk402lWEmGSFRsGmEwsBh2PNccYPLj+Xq/hpxRR4l7
Qz2kMtQPDcMgu4M9XJqvIXCBM2q3Wob7UDXvLJtww3P23Pw8iA68KEDwhj8N51DT+r0B0iT9giHL
bQN0YGqJ+7Xuku0nd1FIuWC2KNwlQKU2C+ztSStVHlWfS/133EF5n97TvhL6C8ebOSf9mKcyHoPV
dNVn0RfjUMGMtrHp04pmyMP/0XuAP8r3mtz9jw4lqesVsJPGNnYiUaHSqX6t9pD/vjcNJc9yc5PY
/FQ1uqfSpaUU30kpeQTN4UpANSobBJXQBDMG9AFYWuMX9yGc3Hj4rYdv/MhblYRvIRmHqyXj6xzg
6ceLMhTcNSx0DGAttd5fK355RA/zzzefbMdoZZZA/DIVqpEXRwFp1jhHKzr3EAAhaA5Gt8bq3FrM
SVNR1pym15w1dRpFj0Xqojlz9uQwckxJgApY3Yxaa/60Tr7ApmxarPSz4gCkvCg+HB2wYwhq5eWm
XvlMa6Ccdz5gY302Rdsvvcu8YsvMH2GIyR21VH8ia0Os6syUWePTX/TdryCPwEJ8GY6XTqDAPN2b
h6WL3u7E8F4/j8L5LrlzoBaCURpNApbonPyQ8iJSRGjDQsEaDWLac1ArWaQZAcLrSUgxKgZ8YU3P
+3ZVa3kzR4fhxoNtWtdDy+HYTvHyhoXiYOmy2e4V3JZU2lC0BdUv9CLQuY2w8yOviyj2LAVQA46Z
qUU2gq45xjke981/NgJe8pS0d/91/HOIrDkKesWwBUpc35PtMz0liJQ8PfFyhoRDzhK6xwnligo+
QPE90NzVqluT+Coiq2QbVJmyRocVdQQLXV8FIv2uX+JgOZxFZawHzIynUHFMoVMhkY+xbOm2+jK5
mgfVY7wVqWeOmtm2VWZEW2GWtEO9yF0/sz6mTEBC3c2zNsQQ64S0SMTToeUD1oPPlNa5fuwDNIfy
QXtYNHL/SUtmQsSxNRVSIyxOoZJnh/l5AKJrm3W0aPj54P3L9pxzm5zYZNU0rgFECf9blkFH6X4w
x9dFyP4MPSnAn0eR5WFQmuz+AZX/E38XTLwP/ffN4ZP3lxiQB/kxRApf/LGOgkTJDs1C4BMNE5WZ
y7cjEX4yufakza0IA5nayLfjblOkWLgnTJ2GTctTM85JEzQ+wSOVoPm8wxM49DLmNCiIVgYjhtZm
PPSD/G/KWuqEr8b5Gekj5GOGrDYmNp2go6QXZKqzm6uPGnxWMX/h/8+prnj5kmfzQ9qxrycDkAjI
NPIB5js0BnkEVtU2e2tHx1Q/D7sUrgbiIC0h1IrH3nQQ6Oxy94MqZpB+d6E3dzuyX2li8jsCT3ES
M4XhhatbH8Qow5aHvlg3CseQynLIXlP2T77CAGQ1IfNc/Zla2hYJU1Cqq1wNzrF2hWiWnJs4J6fr
ZYjQ1Eavg9WI6yagqTqmNRW3V8Jbcuz7171fDeIwn5mogT8/iGDT5Ps/kdFZgsSD4XLt0rKqnlM3
Nx33RbKnnySi6eBRTUuJmCvav84w7orB0xnC02H8cA160x9Xr5bNJr9bjPLs6t8aCUlqxjihXKTe
gWh93rg8hxYjVNr8ZyYgodL3lFWl0t5aDeioSlxJ0ohqT2SdtRVYpyXIp92zCIwYc75FGg0pXve6
DtC18jevk7IF9VwVyHDHf8qDl1lepnozXXiMtbIB+tWkgGAfQVx+ndPLmafO+6lHc8yw6zC71SS2
K5JYcy8qbwuRu8+EcVdnLYPE+25VAZxYu8ClAb3vf4A9txViJKvYooZaZHLT0XIJa+n16h2TRJ20
JFMb2Wrm5AU0GgvHS3vpUp/SUKGtlhlnKdEOoW7HAFqymXCCiYsvpwpKKrGrnD6yV87BjlNRK0ck
8WWY54nwid822ToPpZB3UISWW4tOxS7dJSbU6Pgkue+xjzX5JGtSRVwfj8sg0sWiO4vyLb9y0lmQ
9rub5uHchKLTHiQqUWIbg6nu0TSjEJgxMxk8jJamcoYgrHAvDefwO3IzrgrytcCNJkj8IcV18/Wd
luI0+zTV5MhNkX0YL4gDUHUmJlJsrxjf4cyHou7fl8XNhXeJi+Pvy0kN3HEXVO8SNh6N+qcDL2PS
tvEB84ES6gNLrhF73CX9dnWFEK+9sqT25AKJH/1LfsWaRtFQUlR/oTzGBbL/V7KCaQemQ1zQHjqd
yYBMMPQnvhK3EOnULep+7GkxeUcFIVI1xVXISYu/y7HZHubHYTgFyKgBm41Pi7vf1aGXwcT0lXQv
HBfZMaSzUf/vnEpfnGFAI4HG69wv0/xR8k8v5Rg1HOZgAVK/n8XUAryzT6tFZgpwp++SULnTFQ/p
hnWbEql1S8isgpacjnl9EZY2jiop2bziV2A/qzIsGyamy0pzjuD0mzotC4AIBJfC/23wbV8QGIKw
2FJ1s2zUDuEU1z/t9CWpkq/xujeEr8caKe0ikGzldS1SX5gez/xWbOG5DPsE+EdbrOg8aIHc7GWX
hvDgWPHt+zqcGadduhT0zZL4TTkxO6Fplk71cOXU7Z6xOej8ynMGFnbtVpzPMSh6piEOEDWOWYCE
vjvojvyXXzPx2qedaCckXg6RJaLe+N4CDlpny9vNdlAst+oTs0WdhV6NMvSmALsFqOzeP10WcWzI
3tyvLbCdvmpQxyT3D0BHpPro0bEBwa0qG272hWGmiokTnIS8hjO/GR0enDu0PbZKR+g6ASyM0iFb
4YED45vC9N0FoM9QfV8kdAHZauy8btgSDOoTarjsdF14DJ4mmCBBjyelnjf6UUjD+X5O6CzNe/RJ
WHq1VE/II+0FW7FBnoOzQ+39bX8GaK6kFA56lr1/sjFQAAhIWxma8ScZhfnZ9zU5g6+gct7+x+pA
tUvPLApDFbUQ1nWy1kby+pixTw/BgfEJodd+ixMeqvJOD6XBRBKHak0mEEHHROEs+eFqCilJJK6w
4n2TA7XtFTk0MKGtxIj+JGa7esayJl+q83Aa5c8vpZNnZkJS/5/MyTJDlrhTb2Fxp9oqrA2jgYTi
xFSpg8w7GRAba5b/NWLqKvFkseaS7ddFrxsZ+6cCtmfJZpJhYy0KOSBGupdr0gdxN+q80PXIzYgZ
GGlMEWlcOwHSj8gsddtkEXHye1N7hgVRyuod+wAqyykaJQIbl/RqtSIG/zxLotgNL69z3prW03wd
of00cPOKOrZqxO4eJ2KUkT14xhQexUE3ABN0wH284p0tiZN9rtsao+AISkh5YEj63hhiORT+WGvU
cKOr4zGl5NulK+wOgSr1ouEVMZuGsGEiE2/qrC/Mb+e7kkAXN+iLBR42eI2IfoNmnZvDt9Wa4+SC
IdszkEirFx3ChsZdmbKfANsCAy+YKweZlsEbSeSUafkEdRt55MZuzJhr1+6vArNZPXF2oRELP5s0
gvRGcopIppxW2sVHGGmnDbRfbm/y3z1TbcthjCXoccyM0P7GsBkNs+lObD2I4E5+vIm4TJ+IpOkH
LqN03Kmms89gElP9Y8415eZb4AdalSA6evZSCDVLzXfJ0QCdViinVrn6cVEPaxHEuesnnuIOBmzp
EUJ+LQ4dveicOqQ9qhP8EuZ/tXiBYSVeGJuY5Qs3VGRtdhk59y/tA7F8dOI4o1RoJgZJXYA4fp8i
kjql7D4SLu/4zL+pSnFV3QX7CgRcHZlfT7byCDnB9+VGUQsyJ1vlZRP/P5VvhNJihENHZPqkZTIk
REiJvZH8B75hAC7y5MTCu1RZed99/i+98/leIBodm9m1dNNqaq/CoBaFjZPUAMlP2rawFq/n157W
Md3lfkf6SaErZY5gStzJBvLU3qAdZxg5rYzkBwj7DlCSofMkbphN7bPCaC7rz8KtR6irxehM73rg
z7RUY+OWRXJRq6xAKxJcfqZFTbBERYBqkN13eZ6M5BUVX9K/d77ya58gOXSpu+iQBbB53QE1fBCQ
C1MSH5p2GGOpRdFJb5nFAX+i88JFGpFaPpJrrKM0glWM7A879oyLgjrAFmqzb4DOHqhcVZqK/vIq
dfQ8wH82y9T/1b3C5193hTbKnbgIBaEu+QoabWQwJQXr/FTqXklpzTuZ3HiX2j+C0xjrynSYK6pC
AoNx61YcuqLItIQ1H8qQdKV2Zo4DL6CmLi9bvukfr4q8j5224SKeJeaydQhat5gi4c0fA8lUIX3M
PUYMxhKygTc/t8bT43vzFCzJ6DuKVzOsh5F/2p6q/R6fASvc6qWbyWU9M8Ns7ZO/UQSkseVPzPr5
wJ4hRIyqzHzR8L6yHVzgJEuzezBO4vPeni1TSzbQlcR/2PbkM6daw2ZZqW009/RBjG3PcdPEpeES
0vegedexoOD94Io7AL1b4P/+lpy/7UHYGST0r7nJPzd96VmJIqRmpPP8u11hanh80BhkFlrW2HtO
MuUGfB+u7KIxJ48lFGUcHZ/V/x7jZYYPsr7MrJjDhLRHFAkIlSqpKmk8yfDJ+qEgM2prKPAgsS+I
SjDuiblzUHFV97JVnYD/cjt1R/YIWiFnOF7GrHXYJJQMGJEeaZ21pEZM50sqJ8t157eXwtdSijc4
ODN8XTVzEsYZ2I8HrNQJpX9iWskbHn903wn+96aJdgAeUEEAQN6NmpN5RJ1BIX+XsR4xjBphoL/i
xK7b08JpaavRwPnJAKfgvaaFKprvLo9RxJ0r8tcGkr86MxFkZGAkpvr4moCUBjY/8y+shXroONCv
Urib6yhkmZrsice3aKQJDAJAv3EuBd0MBqXoLoi47whuKJkVCHwQRVKXiRGIx8psoDCAo9mIvurQ
TxCbKTDV3ZMIO030SjQDzcajyEwbZ1iILRH+uj2cAQFn5e/aodEBWfZwWxK0MQK1lhWSlFdKt6EI
tPTPe+wK5U5D42Tw8H2a0gBzu9rmyZar6mZ+zl+4ZFFRE/E6+qjuvCGdS4/cn/Oy4xhfN5BW27jD
bXtfCyd66u2VL54DsC/IJPCfdrcVZB82sAlqdK78saqK1XyRXu4eXCeK65DzMPr1ZSEyKg3KYKZn
WUVufWz9Fj2vPv9I4N3YTEPxVepctOxPW8qRZ7usR1Xx5JdmngaGwDey5/C6fHOu0jbHXqZCAxTJ
ssg6H634VvKWVz8IMDOQYscaKx027zBn+ou8ZzhN83MlRctfX4zQP8+c25KlvmZN70TkfOXQrHUC
BffOmkw711fZE3Om9CM0QPojio36vF/08MXxRfI75mYKPUAFfl1sDvrNtEyD/Z21sY/yWJ7aSM1o
18mwh1zPAwPrqI/HUz809kLIGUB0eH5XqCxhgIi6uCtpfJbKV7dpr4GNSdMUECOb6hvVrbDpgAx4
K9znYFzy3/bGwu/LOI6MEcnK80Z0E1I29VdXZRkdCO9R4c5QPtkx6VE6PJBPDabi5whv/87l9iOz
Bsb85oYaUirgAbiExeh1PG3n3wjkYTsDYL0P8t3zMNqewV25iLKoUov7gOUq0i/kS/wzRqZLr+sf
NgKALcTipJCc4cVoXMQTDqggUWovffTOHjAAKI8z2eeqXHDYDNH6wcfayiWNPUpwbDhYKmwGEb7s
B/ArzeZgY/jx+HVvmAcZ5IW+f7mqu2X+gbPREBFCasWPGzblyhDhOvWfD96DUYJ1CGWK09bfTmj8
VlvPty562+pazWsPEvmgrTzfIAsPaT6tXDXRRoQbcQLLbBKHsRU5SqFxWUlnAnulODdWMckW5H6S
/gvfqrSiKTgyVcNGionKWMj7PBkTeuKoTbJLWz8V+V/DdHZn13rdoVCkTW4emKmUHgRk08ys7KPg
mItL3YRZ+s/1KApgWxGp/ZhRraFrB4O7F2iTuecsSYO0i/Fvs5q3M5vzwkgSvPg+jmN8MDGddIqr
v+YMWpERMTOAe6rr1/WlaUlkFS64au2JQuwEbScklKMtg813bJNrIXnGHIOEOnxsbexATs4Eg/Q9
DBYT1GFDHncCa8hMPd68uU+6WIIUhG5KpiqzHHEX3YuOikjcJdP5RD3gxsIlBjdtg2pmqJzjtsfq
8gWxrXLirfnv/nXaRCRSY8lgypSelQ2zSDmrVTxhsm/ViqeuanAJyaqydBVxEQ/ScmxYFaWUITZb
S3WKsjNXsl8+nmfAMWsmbHuuFvW5ABr4rTfZHBKjJLN6ONbJ0VSZUtL/gZ/tV4a2vAjOhS3+aIFg
uJKnCjsXW1lSZ98IwVYSflcMEH2Dxk06491vLIOhjzzejjpfw0ILG8Cxf/7/6AytNSsWIPQpLToX
SAkSfzD0yOMETd1Tc8y8TG2Pz76t372J0dT5MvWOOw==
`protect end_protected

