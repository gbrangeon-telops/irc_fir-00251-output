

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gqDFw5NFAM6CTSTQpb6ewV0dkTDze+wC3QoGAxwxbjcNW9/DsOht+2F009+7g6jE2OnhGLtqTq+c
HspFg2GBAA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OROCzcjj1wgCYlIqlabkGZopoXwccuhDPoDiFwbBlsbzl7flKX8tC5m+07o0XejIs9tQT70vCTz8
eor9UB573WqZyEwu6nS7RfReZTn9rXIEfFTmb5LNQYR53WQufFJWXVGGzbi12Azu0TUMNBykYjra
GCJvYkOLjulS+N02/QU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y306+4wGPVAAsHa7Tcr0Z+Y/dNy6G34dYeGbx7ATqkdiT3xoZwFMriTbyxCB/BNDpEEpWtR2x6B5
1geIXl7xRsYW2a/OzYZ1VgC14cIMMrlyvjd+Q0oeBhNwIf7zzOU0YeLe10Ln0VhNNlM9hG1yxJpm
PklN0o7dbe4z3qSMhzdrqG9CNO1AfE0zEYRDe4xK7ci9EcGBPeIBnjhSSGUwaUeKV6BzeVeTBH5k
pFfAdDfvgi3P1VwvurSSAL/VyrhWR7M2OhP7fekXRqEU99K00pFciI0NAEcJPUl8pbYtjc86ccu3
OmuQ0fZKcUeaRlPX6glqeiiehMLm/EPWzCdMgg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gSn/ibMO73s4UyV+DQBAOvPjnov0A3ONpbzDn5S1gDHbJc8laliw/uAOvABs0KKAN8Q7GKr5UYxh
qWYO6FhJPBG8V6RCU+sAaoeSnleJb/buC83HgJws4chUKE1EbA08UnkA2E57wCSfAlSkdEQl5xrl
E4NsCY7zrBmnjMH1Xu4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lI1FhNfWvnI088CMtuEIyHMeXPGNhtlppeaUXaQvRzrpC6F1bRvO696fznybaYq7K8VPJB0YyXVb
8oCJzTtV2jMI6KoF+McAzbvubpz0ru0XOCjjvcTsZJ3kGxHGUlKh6xdlB0Gez6kASJJe4GeTuEaI
VZNg+Q6ea8OLPKgQf7VICmBv1vM4svyVLDI/pSGiGOmfSMrfWDP60zo6tHpkaDS7uHEj2WN7lXT+
Q8c1SGnQvLeKyHV/kGG66fpNSvILAslBR0l5Xt1/csaBtahK2IV70dxaZkLZ2c3pylf+SxXTt7v2
CzVvxEgWwmwKjiuhBgmVM6qeL7+tokO6P+FlQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 41056)
`protect data_block
0r37bjYl1D+c0WVLN+70ysUoSCk+E1ePlOIU17qqrO1fq09FafAzMhKQLIKqIoZ8mYjxIwBZuUwH
9nHLr7Gz9QURkCyP0erQO37fxYjrZhsDQZ7N5WUe8ml3xC56YQLPbOly25WVSVO42oMBhS5++S4V
IwnoYIg3Wyg8lDa4kAlQzxZr8kwMT1GYw5WZLXROGbzE0SP328RbjmSKVpa/RJAyUsu2e6vWRms0
9tOV6vlSZhRH/4n4GAdqWxp4JYUQ9gG8UxVAU9Xh6jqsB5xqmhL7iRY+097W97Kmz7it1MPgqert
wWNnW2TT5b7GacToCZOIIXbpcKHbGFcfjeTiTSzjO3MhY+7kwnp6c+e711gE+hwMZP5MuwnU2Fmb
0iboREucgm2997SN/zuYUeiFL09Y2FFgckj+QNPE94I6KEro0I0cQZpEdnwaHI7NKyVME6ouwSw1
3tGbMRePFzgjzPpQkZY+p/YD53ZFiq55F2Ahpsm1L0mffAf2PyEOFqLbebCMTlRd/OXa5S7r+sa+
EY7AmCwFUK/W0Od6+BVWLIZwVTI2dJuNUD/HFioXORgU0NHuW5Yg+0zdgTOWAsHNL5DJRIQYTIjp
T/D8dS2CyEUM2Gj72VY/zJ56JM/G5oRLNVGBwgCp6jEQerKuVO6nNLIL47vVPZZpz8OOsCK3dzUQ
nkIcmJNK8lC2+7QzFSKrg856IXfsciMVfaLEyBg7dVITCkhjwUsugwmpblpDfABXbcDIIN1Xa5wM
iyMtE+Psjc9iK58Gci6HPrE73pBNOWi60PWkiLyFtE3RrsYPg9PTTj/JHyn4jvoRRbc6/sXnWSWc
T6u895J5n5YTS3BoR70usWO1Dfad2Qb16cq2h3EdLrADcjjbXnTewhtJbxfOEzwKd4f3vwNnQdJW
H17JRLEspNBYZrYOT9Sae7YgN2ukekoBTMJo6pTMPHYqrPUb66GN9N4xIJzf4ytqu8Ms6UwXhvSB
7d2TwLQGfAkndit8fM8gxJGH7WYcRpkI8FRXUdAPr2vIKGWALIQkEghs+hSEnfpQXlCycFqVnXIN
aOcjvXRX52eU3vgz7sEAg/RG0DnjJb8W1QNno5G62n208Y+7UBEXURoXazIJGrXX9kHgzyiglXgv
dFVrAQ9yOLqPHQDlP0WhpTJkldZcQ3Hdq+i9tUlbyQ1s17EzPE4K8YEpvOKtJw5THeYbd5WhX3Tl
9WKrQZ+2iTjMObBd0ibhnqIl06qbBBICEaehCuGG4MY3PzjVhV4kMzBigdRbnafD+jKrCV8z+vn3
ndSIBPfBnrSdK3TLl895O/b0C6ph1r/DPEKWr1RDzc7XW60Z+ljqgL5CBS0kAa4Nz8hSuoa+jzHp
C5nx2zNQbkm7Wp+AOeVr3RPeeJJ3YiRQhDaVEb5uw8a3ml+vXeJXp1ONaJO5+2wHHYQlonHhVjtK
dAsuSha70vRFWrEMjLGWweIZzQ962d0o4E/veW2MumJGbBzKnNL6IzNb84RsUDBz5FIATDEYVnAv
QklXLETIZ675dbIrR0P4aB+7OxHeqbai1QAjzuqmkL3Jt7xTcsVaQ0dWWEu65EVpWTzws2swgKen
WlhniiE0eZrvPgJaOeiEBz0pqbF2+lOovI6bTXBoPDCXKznK9LwE2LYrGFqpWRfNUtjf3dzfWpSM
BvgH1u74I1HnkKsBNmx+1YbN4WjvhBircM7E6EeeG1THz8wvXOq553K/GB6wQY3BRWp8ZbhPTQF4
/OlyeMvTERRtwf9aVNELcAwlwWxePuIVbPKg8uR4nr544WPuaNersc8qIpM3zoJVFudW2fUUnErD
0rQgPNHPVpDKz+xzJmVbLw5Zh6XUDP6z82Yul6GI4qEoi/EI7Ep/7/yppa23Q1VETcPn7Y8vlp6e
S8U0dViU2Tav4kZuw6fnx4lKBE5Wx2p5z2kfW/nh3fMJY6saS11oPPeOQPs8GrOYWbT7FWeEE/hd
N4WVcnmOp5g5uCgRxuVfe9AZvacMp0jM3ETfF9qdYa9q9Fcb3Eik8sHvjPW4eJ+ZSocAfwHsNClN
xLXNBdAtggQZtuYKDzAJ0pHhOhEx17yrZ7kSg3MFdw6/MQPTUd6IU86ueeJfnQh4kDSfMAgAdbIR
bS5f7Oa9BcO87gHyQz/1+QvqLlTPsZVQFe6N+vNChILImXveanIL/pXCSJu/ViLu1dV0pezye+Y+
skGPuxujqARrUaKX/t0Y7oCeRSfbb7WG+vjFqgM3Tk8HOt4Jm2JwoHnC6go1AVHoiEkWvfQHm3Y2
xQSoDEnG9S9VQ7nBqr3pL+bsIat5f9orCH4Yk9cyf3lvJrRFWn0ZnXyKLet7js8sxoRht5UkXwKJ
pNAAZjR++xxl2d7Fom3ttl4+Iu61BJz4tytGHOB+AafQW+UO0JFskq8sItH+EuEKUWXOvtc/PUQQ
rE6UxBxwVjCcOoLUVNewS4DO2lU1vGHTXArq3YkU72ki6NTl7PtZF+W51AX6RCaX+vtBvwoerkD2
8Jg/1i323+TLScQ3M1j/vVliXk8GIzVOqJ1oTj0pqlU82K575wjK9i/U7RMHK4iDSuI9Z5gX7rJR
L4m1Qo5fAxGWxLPSYFG8Q2TKHGv77nMIgRA8ov7bbScJ0E2jaq/d2H0TGZOQIDZMZi3kX/0sNcWH
zROkKORtc/sQmdEVSNF3LYFUc3NRZLNWm00GyvKqX23bjFD+XMRGzgmZvu1ky6jE201TY2e0u8QL
EXlXoSeQTgFvqC9X4eDc//Iw/Qub350A0NRoIIszcKfX/38P5lkeAt1YF9OmOJSlYxK1d5lD/6Vo
WZyve9ztIpKW4tVht8X7ZhYAOVGSn0Teu3L81MEDctBcwx8ruCiawK6PWV5fFLt5FliX/TUjAvqG
F4lS8m9gvwHzu3FaHMGl7SNFmY+ptvpm3mcBGoS93ev8l4ZEeLyCgML1n8HB2nKm0j35cS1mrcrr
v4UJo7eLGc4shSgohw1f9Qkz5TXrBjm9SR8Lz8NR5cAsC5ozMXPd6Z4i2qfDVUN8eaulcVe6oCe7
TzwatXyl2HV0KqC+8pcIM7VaSMWc/Zlbe7yFgHWdpXeBEYoDcCEdKEn75q9Pi/Yb9bW8D343Setw
4d6ZxmFLga32AZjHTAu5r0MyHFxMhkVVCbmiJyzGDieLX7tVmvbcNaLfYybDUCCLt85SwmnFDUEL
3e3rc04/UbVukrWOd6YbuFEeHpKPRJj7G9lwk8ZPwUXdbfLTuQa7VCG0IK4jlsY3Fdh0yKNCXJLx
lRaaRJs2STHZaudMxC6y+gLjYuh457hQl6V15uW6OQnWOwblyJ5sHITLnVHBk5Moq+meCwNU/2tc
7ZDOrPf0+UeRq1glWHUxUk5MyaFtVmO/wT2UqKm5cChr7IUzw7XCfCjF2CBaYO2kSg6ysksV4i++
Fqfv+SfNexL37GNTKMxHa43ebMirrEBaVz3WHbJ9wLr5kW1TbESMEVjMizxVce6L1+kscc4/G+v0
3l94Juxf2zysjTd9VmkNiP1xsML1dBFCMa2NT2n/siMTnFM0bK8zE82ga6bmxuGoCm2rg2rK4k/b
+wFY95/sQuAs/kuxO4OBiqpdWZBUCAQM0flk7TW6Mr8co49eKsexPEcIgPBblN2+3c57QeQWze5T
zFmaw+EK+/4t1pikgFYBtYw6myHt9AeYdl6Ik+meBxQFwDiSZuVgduzQq6JdVEs3El9eJPFyFJMo
mjMCrG40VzWxyRaArzdLVmug2JvyN05ap6+ijPCxusFqQtj3ufHG97S7jTQBQ3UZtkav7zUdu3S2
QfPMKkqEiITrb6s3zwatg7R85tvalbR7v+QdQkJYHZRT1/e7Tr/7ICnPEE8S04fTPrnkW3xos7q0
ImP3PaoMXIiGSmch4I9ehNeJ/FTnurP3btiA+nkQ+lSRUcSkOzlVZH3ktahtCWpyDjKc0v1nFcO1
kWPbHz/oF/JSLkpsk7mB0t8jK83KsWMK5wkdbUE7MSfDseEBEkvguge5bgkrd5ZW6V2/cP41Bu8P
g7Xg9Q/z4H3E9FTsJGsC/H+8N6Bl9h/sw/Yqp8VPFWBacNYigLU7K5+fl6tqnRL4u8vlv7y0PP8U
DcYi2E0VMXzkzUQDn26wry4yjhsIJvcfUZwqdLsTp3JIj4UCz+aWi1a8dG28342pTzVyElqTLbg7
T6Ml2G/dMfN0tOR+/5x2VY45vNhLXI5PvYjCeKTzcPoJr2jMcc773NL0JjvNa58QGxTAnfPNJgOg
GIWdw3Z8YmPeoy3A6VmpgBBVdLVtAuYtWZQGINb+P5jTMHXKfbfHNl/PwxUjAnOBKag1N76vl55Z
WapRhCxPRZ0BmJqv6MXJng8vMrFVjJfpmwBDZCqVJv6gXh4Ye6d5Qwh/VRbqhIyZnGT45JOH5aZV
51N4uWdX34xCChqj26+GZ4DicxoETLvoRwsPPPtKypTPRv/zwgdHAAZTYOO50pzI7Ky/lHKifT4S
0PiRjA3H+FJXYdK892KPIZuRN6B85qfarKZlv5ikbs2aVv6seOm87qKqflNSNweHGiGJ4nfCHfE1
RfTk65pcDQztnXwzZ4nafBohe9bPzS7poagEMmkwPcuY9cT2Ugqp87QoDVfdDjLqS04Vwjtsp0gc
KN/0ls6csmQCumn0MZHeUxsfbQv+YJOrmWAq+wm5F76FBEQXsjleSMtoOAToGynWsPM957cO7gJ4
tx4kcUcJ6KJSERAVGVbyuUCINS6y8m7ufi4rxgGYFmrFnv9NQie7+n9QIwP7rdUpHd78R4FnzSER
zYKGPlZme+gFnleFXCgmfHJUDqgZgEBS92dQZGkswX4JMCBD0Nm677/SOyYa6iHJArbINGY7/EMS
tOf4+RvslPOoYw9D6kVPL5n9IhTVglT3HpQ030pA3WDeF/s2kULu83JWqgqdjwVxPwUNHNsXpwCG
RKDB0ikNCKIIpNkKBzXqyhdRKVywPy0iQG7Vf/lPvB6OFgS8G7Xu76CglgVAVs1OHo2b8d1NBwU4
GZB1iEch7xe1hk/+mJzBGZcXh/YGhhp0QmyJ9ne2lRNtxIqvEgBIygQNQCd5OI1zRnub7iPuqlFA
qzJofAeFYulG551wDhZkASi9f5IkiLxuYWRGBVCJHG2PaaHeFZoH2/fj27DidnaKb0WYvMlynDSY
+HSK2gj0YsPGzmkMPpIlTXVF0uE3FmMmZTfYbjWoa+bNJ3Be8T3Kx7FEYUUe1g++0p7zh+niAwzU
SGh2vTpFj+oJ7uD5mxRwHQ348ENljXydtja5mEL/qiaL35y8ZbCN0MqLDwufe+vk2+sl1OOoxSpk
6q3OG8eGNvElmZCubs2cnTdhb7oct9dmB5a089loWnPKyfV80n8MMzijf9Gcq9B5dldRNvsRdDQu
SA/yV2kLl8Ne7qfAnigCPhkr9kFQP9/I9WJ5nWzpTGWOTWGgrChucK8afQjYTdWdKHtDyewFz8Yc
XU81Tk2S822kJGm12HSVZjdNA9r9Onoi0GLz3PnUc4OhcIK8NKta52X+rIypzJD47pw/8ZU78744
0O+iT3xvVEywzpslx9JHMDpg1KGwfG+xqAB+p6fkMy/b/errKCEahLJEJt+SXVG8M7fPvW4zxznQ
MekAfbL9+un9IpehfuMG8uOPVHopoYqIgB8/5lvW20qrJ1tac0n6njT73LbHC2ScE7vYDoGZKdh/
Zk9di+V4t/zRSluqSoey7awJnptDyN8KGqLgGWcVwHtRCnGYauObTTbSueLpXd4pQLf05MeU43uL
vgJ+gf74ZpaOliwclc5E1wycrwHRVWP0Do9h1gr4MoqGZylZ7q0KoqY4xtqueupoqAr8sVj5iIY3
A5vboSklb9ckv5CO/19IgMSbyhKy5nHh4kzkblWEehfa18sT0jaPtaGnILWTp++zG5GrTzasmYbP
LZ5kO7shlw3702wb/hnQn9avTHcw+V0BuKrGX1qiN1E6w6GR60CrkXHQsQYMwKOxGgRCxE350AEN
CNrwbGozmC9AsCMnZpVs0ZgEYil49qaAdKXZ5NERzw3k7Fw166AjPZP9XvpjbsPESjp14tlEvAbh
X6X47rPqLvjbqGCdaFE2l9QLTPVKs9hLLR6ivZxvckQpjhm/Vnqc+Lg+uardINb3frPTrVwPZgIi
Oc82IHa9oTtsXLT+teFFGE5/DxaO91y1V+0DVoEbMt/4FhRgDr28xf3q4HnrhaGpZ8uKvC7EM5iP
LLfBI1mTsDUlgC/5PIpgg2Qom1rQyTAv7AT4+N6IaXWPQReymZ4Gt66TlHHXHEKva8aWnLfCXvxn
yGwM9GKcVUPXNA1vqpj7NN0BcFP0C+c1yCcyOoMLq3veN5/FyO+XNNfEDDRahcI5lYqIOXpqDBtS
rbe6dXu9ZWsXLYiWlpKyaKw+7mqXo7b+MUHrV/lvsmN1frjuvend26IHEZSuUrRAkysWe/5ZrehL
n0RAK268euoywIui7c+J4GFYP36PnTltkbDBUag4p1WEazWLVFuMUOioA1x2z7qhLC5w1xIYr0Ij
cfOwplxAhxKXRDuPumEJv+f2IBVssMJiyR5iPgt71ycZnvbjcGXgdUc2nazb8AUbuuDN+5fpSQ3i
Tb93raO2kF3mTMfkokUIGco5818oZGXjpDfzoPEUgGCOhn77yGFL6mCfj1yia5okE8jajXrPxOr7
bDMmLoIUNHJ4D5wwgWdgCpDXENF/vDN7dfLeq4nQqeM9Mw0oSZ4DhXmoPZNc/DyYiitQ/O662LN3
yhpdkmAhLyfvldbpYZqlKdLSS3juahGlqx3oQAITX3r0mpKgDtDSMUekqOBWK4lUcf8hPphUfQD3
FbvBsn72eAN0mk2BvUjW4d5sFA2KvZgc7y/qXeZD5HnyK+w+dMnhfuLhqqm5T+cbLiuvhsju49R5
g+bc4sy7xwRiRbmENZA7zfQocTuSTZRGpHPiM/pm+8gs000b0GzEySutfXSuPH5b1gUNfyINEk24
4I4i0vM/HKMcz2N9ItwhSK4HjSLcBAlll9UDleouoOwZuIaDKyjNoOjsGQREdPF+thsrbvGt9ECO
VQ7phwwySiENhrIHFgYoWQT85b7kb+sAxI7LiSDed2UlOKVGbHsUYRgf6kLxY/Knvki832qaJGDd
2Y6KhJOUAg3xDlob854vUD5FTYjpBVSc90pzTIXwnnpUmIrKuLpcncbbunBrmeDOvDE7RimeWW+q
7vR/YSXH5KukUUgP3aW8iRp9jL55mo6DkqsR8Do88gaoZ7zRs5xlcUkakNpDs3p8mgJpq4zAnrhf
+TLG9THsA47DXivdYHpSG7jyImmBVbofiSCz48N7WcJmx7L22KacuXSeq1EpV0B9ozFm8ByJAKaY
CuH4hJXGR7O4yU5wj/2XSqLLnHhyTCGVskstRmIT/OTZK3jdMtOXq6nnOh8TgNYc1QJgAtfyj1c2
fJo409zhnfCurZpjNrElpyZsRH4rHFQt78IrG1WsnyO1jSTaRI7f3b6qrHnmBGal0eXrHeDx3Pyr
5PIL6dBBJndsjZhRss7Rw9uJk+1xYbm09qoRT4zVd56ZlV/LOHUO+gFfRWv2NEidvjwuklOLI6Vj
IT/HjJD3pDy5YfVcg9X6zcCtyMdNEL4deG07nmoZQiXZNy+mNMLvjhmxGVTN0tcZE+zysYkKy01V
D+wbvlCPOgSUxHsE8+6OIwhRy2DOmdhwM8/3AO9D98sgWwFx6chHDlLg8rH55tFlYxDLiRPQ+q0N
7W6TZrxfm5h7FHeiPxexlBs29baqj++JzUulPVqJ6SjU73YjSX76m//0bhrS5u4tXI6DBRX2Iv9g
TtvTcRhnAJ0VMuLjKg4Nm2O8ecgqu+Z9ssNJ1nRPkpNmofxoBzYRHfP9+54DpfkH+IVyzI0ZuIKF
py7ItRrB2dY0yvbP1fpWuSOjCH295L6vnII7rWvvjPheO2cEv6Fk4M0EL2XmkohyADGfMa8qr6Gd
+Hg1fLjSGyzibsXBYRqSB0h5F7d0teQjDf9/xkFPUHoRBu/BXI+ocguC39fjDSjf5Jv4gVTqZSvE
8gNMGoLSjBWeSVT48IlGtNtqaEQsxlz2h10tcsUhUnCKUuFKTBPKGN9LP0GqDoMqvkua87keX5T7
VUrRSXPKBK963MvTR3PkRnuaRqVaAYNRezdws9lh5Od8gOV4Xe3/kaB3pXJQS9R7wBuRGdqI4e7Z
LZQ8gqj2dPONisDfWb8A+dTjuawere1jUKWo3xKP0iTBx2u063lh+LSFx5d/Jl8GxX7G5e/IoqN/
YGTlxGgxFP2/KLYgTo573DJu5tjVUeacbqCGzIBSs9b1fW0y+PvjhHRS0qtQv0lDMoOlZbH53wak
F2HMsAn2dgqrVi9egBubB1x5G/fuS+T23cDidjeyB8rWSIhTjN+kubDvezlCrHP1Zfgau22l/SSk
YsYY2jnlLCGc301GRzGEd9jDfzlledf4+DtjZGQFEm5QAiFKKTBS3prevP7TVv4O/zQpQu1I1WU4
59vYreTCY8m+KY+NmgX0HSlDDCvoYPx7/1Nr0o6pJ9UcZN8gC/eRhUCB9mTzUN6rJ8Nu7uSuWogG
coJ40k5T32k82uCNeCSCZyJ/BkQCZeB63aMjE46mF5VnVBYi9t1cUudwzMuL8sF9x42JH8qFveAZ
JqHjG41NZSsoocbbpgopLei6c8rqd3oUfbyRfR8gvZahq9ruI00NjtSo3qLTQTOf9xXV6XYsmEfu
77ELQYnbgBvWJkGhnXtfUEmdZNWQorE9oMMvgX8aVplDEA7raqb2NHDBEIgpKMHkWVf9rtriSn2p
S+VbCA/7OE/41sEBaSSvnY8xl9+UzGzQeqlbbf42OsVF9PKUZ16moGkMXuEUBULlJgbs5WaBQZsL
Fvnuf9H8ELnGNfaSAF1aKGy5vyYKNk6EtrtEw826Pm+6ATLZIKy0JjnTEpdi0FNi3SeJhBHL8xsy
u7PgfiMOv9i/CCR+K1GmMp9HT4/rwTUmNFffjGpQ3Qf4t7OxGQ4TZdO6LJ5xNVlUoXynigALb2pI
EPB5fp5XYfTqHwEsTNlipZE8mrahbECnMYYwcd4XlaTNBX7xDfRMR6GSpWCOu1wS/+DbhrSOiu8A
Gw1wZAyhQoqf38ma/4qW4kgKVnfyptNjLPPsTOYVoP2mTfumMrewiBNWUDPt2BNk2qY3QDCKwUOj
Pi7KOtVoggrGZ18w3ZhV+WFx2f2SXR1Mm4OooPpjGukl7OhrR83QALgHF+U5cWrh3A8n1sDDbhOH
WnPlm2SopWV3bji9btlAcA3g0c4NME7HqjG7GvyOs5ajpOSvjLdXOzcvZ4rCaee4/plDn7IBITYr
qts2hemTtrzp6WtNbaYd7Ht9S/HO+7Fax3XbhOxNhraspiol9H1D/iyyhSHBHNKUb/AaTQghOvsf
ltqnBU6uruBgkzm1LQkcgnvF2mL7Jf+z+4IYPY7udQFMq7k6Glyt//VlmAPZ79v3PjgcvBJsWd/c
Yjkd//4WkPgdLX/c5tCwW5JIEyOZYYSemBFMHN1YXDD/aOgrKmyeZ0DJXQnH2hVi7O47dlNpmMec
amVFBYBIEQ1xvDY5Zl2WcuJaazSDRpyMmuKkvv2pKDETAraIQH7TIGQqTLz1MYXFnfLQkmHu78ry
oDFLZkJo9R7nlKR/aT5jG6uGEl9mm9Sh/2uJF46YdCCSYYiJghtSklxTjEHfS/NDB3nE3hO5JRyw
AFtWfpZRJc/X63UeCtyMZCSvo1S8Zm04r1j8YPAalzvT/5kroaH2hahhgrILGqSNedJ76XTzchHn
R/EiPS0p1Sk3JRwY25Qvc1OCszm7fxB6mz9X6q/DQMaD41tOhYqsmBhYGjx51bGisnMgP/7vNwdo
tz8yfXSmbKPtqG00WCddwtTjDmpvW48/IeiINgDdidNVvI28d0C4/b4r7nnWY8e3VvYPdHX3+4MR
vdqe4DtcfdGRgVnBu+mNzHbewgaBouj/uz6oY611RsF/2VaB0ipnz8sZsBar8WjjAXcY+a9s63qo
xh23yzJiR4vg9QnkhipMrWBkNfdvsceOwm4FwGfpMXVCqN+nxduKFpm3ELa7Y3Azz9TGC0HP80GV
sNgF/jM2qfWM8eV1/Tofw18djsHWKeebFC1gODzyThzG/Z7DOrAgEl3QxeRWS+68jKuymqFustRv
iOywC/oS+xG1ZpAWSSexghTehaUpNtF6CSTxhVQvRA8JQORnQwg3wXRAXXTWOqllkxNcK2D5fLQp
6F3pMsys0f+1KCGjx+QaGaidsyu+LcLW5Ab1YRJXaRpNldmgIsX5t+8IFIjm+TM4PmyKsF/qwOED
bW8NSllxxd6ire4mwwj5SRbvUPMYgU9JIgajlFgNOcNAZqPlnMm4i9qWiAlfqqz41DKJRUOLLDKD
YZ+gUjQG33GJuOEpS6wGjMqmwKSbLuGPN0uE3e45NoxETYra9/xW7R1dZZugrVUbgYXVcLe8uA/j
onbG/7rfvfK14JElJr/D1qhjpWtMr0IfssMxUJMw1ccy2grhidk5cSqKju52GAK5maGev6gR/CFH
91wRz4fkp/X38ht6+ezgX8Va5TwS/yW0qT3VK4th9XCFtTbpHH0DeUZJgkHGdyscpDSO9n7gdYP9
5q9sSjHvHERMXypdQmEb4nSNAWBJO1oklvUCM076zcg+S98XH9sNLAkThouTw4DK7LnBRYUH/Aq3
WfiDHqddQdyGOHC7PWBzvCrxubnHK/3CUpRVPIVYiXvLhwXWqnPhow8g+mQhvKlPHsSgAnuGRY6O
saHkacGBOulXGJJ60LLZTq4nZpYpAnNf7oEwIzJl/7q0fi1WIZLw6h/+T6rnfjRAO/SCnrnKRa6i
oDblzrNUUQdMQ51kaX6wiqDhJQO7wftiYDy6TBVEtgJDUHwA4r223S5zjW/177l/+fh/T8XILGdu
KTb/9wF9nIG+jtWuwJl62mWe82K199zuZDz6uUasNKwIQ2Zk3dKt/kxly7uAFOPob9XhwrH0caHo
1yHrDAuk0w+7ZnalGo4zYxgTCb+GshlLCl7NreMRWZZPyDa2CYL75Wg2ZnjldIbHBqVa9ULRbD7s
EN9Ol8xGgkf8EciLYF+kVOPPUv7xOBqi6PkziLOKg69rbFhbw/nN9bEQUTczc0tPWbCbOIA6Ap/U
KCY0PhFVd7gw3E2PTk+ljzc9YSmzEBfkeLihXotiBJ/iAXgSbABoT5PBObS4MKoW6eO2/5jZwu/m
xSrSiazs4CFZ9Ms7O3lXQdT7llD4iWsFEUn6UDssrP35vF5AGo2rDOkKavYAJAiWiFJzqEn3QNU6
po+064mUBrzruC1zklVZYvYn3MQL9uqwOrC+eVxNv0uRRhjOpqugq+2WmUhKyJr1oYSDTgdoKA9g
tcR74u1nJNOx92ExU4B/BFgcrKF4Yyi8HDTrPORTGLcWzKT9WUSRpQljwtVh77Io2OL9KrupuOZB
Hvswrnpev1mU6vAvcSAerF+oquEuyVVos7XC5G4MQe4teA/KVUcFBy/kIoKj1lu4hk58rZAo3X7g
kfGl+jlSsrn2fK8tD6TIazj6e+SGxTESHJgM0zSKhIrCmUop4X/bdLT72pMGVEOhqPu/diIh8zoa
/jOwBPLzAmkYo1SWnQdjGSzsxQ9dIBrzKUuy84anBDDF2keXeEclhTCUuAYfL7FlI/KpYaQ3epry
SxzGk3i3Sfb0zCxdXW1EZRdkXYZswXAeUPn/wklodcYIgS0QE6RzJH19rwYpfoUbdh0YJEe/dr83
EH2GkGxelcWOccnyytz2I9qPW/uWv91z2y9SKY8PzR3fsmp1hn9PJE5zQlSc3QDK3vEzfHWa7vnU
qC9M6VXrfHRYTNfFvQ+sRSoxjZugjozTDV7dT1t2w/BIHbgbssp1LTcjmeKQbdKo5UTmvlSWZ/yA
DYMobDQp6BYs8z9W7nQQNNOAUHjmSxmWD6R4Cco3/soiKBbj8jDaB70pZGK2kvouJHf0zhlAiACJ
ip7rz9W7IccTiSMtVRemOxyjkEIc6qlFuwarQoK4YFEPj8HcaafJrF47gbGMydTY30sz9VtatB2Z
VOlSPJppJDv0QvN3G0AKxbHrIiYkS6io/4m80wKZpf7FSU5s1uWu0XLi6r/n/+Rc5KSwT+sfQMU2
McV2walnooour9lOuSy4FlMQrcOAdsvdzHk1q23LZ2Mdjf6Is4DSY+D1WdzTDWLf0F64M0TDxdd2
ZPKyAbuTTD1ieCeLsaXAJfxEgSiYEMls0CffPERb/yC87Z1dByXJfYhoEc/2E4LK/KhOCaEJ64Le
77eeT7QfUPJbHjs5N9v163k5nt4z+dmAUBg7XVlqoGL3geTtm0LODMOZnNZMLqcRozevZ68zLK02
Cj571w3Y/W6T8ilyKKmjaWv7WWRiPK4065yHKTzjsTGx7mw2Oz5g/42/8pxTOXPzxoWyeqK34U7V
63IClBQR5jnGubhLd9Y/o4Wgd4aDW2LJFl001b+Jd/kiAlarEboQvr1PIDdJV5v6fw//l/wHbG7Q
ZWSBsU5p2krvI4XHpIoy8q1n/mLZM8UsI91bjLSDXtcwjHAuSVj21Wx/jCCWfIptHPX8Tpm9d/mH
I7pGwCGT/PcXUgB8lvK77Btp2B27sulJB+jOZ4ePPbY1EFlGXrRq3w9Qt0lcc1j57b9Fo1eBNP+j
UFZlgID4VXVmvgsDEwm0TLvYnaZZ44UyeyDA67d50jdCl5QmvhvzIRr1wfVdK+EsXhOjh+OCMUK9
RgfE1ndtLowtiDLsq+LTOPA+2vxInoxGSRft4Fwbal21N3c40wNfcgv6/CvZV+o4UaEDZKmRnhJ3
ObzyUvPcH1Egbaz2CyW0DHjQzVksyN5Bj7JNZaWIpp2GJd7eMP6VKSIK5qGOmnt8YVZIQQklYuKX
VMEtiBXbTi19K5RN3N2sp+0fP8k8rAMgHnoFRD3bzdAdqUNa/rEsLy8GQdTaY2kbGo/Ho8ESCTcK
ADS/mugnd6L8COvoPz/L9egEj4fpi4pNnRvo5/3JPnvUGOTxzm/8sr5oj07m3Try+kAOlAgIfd+E
iqim8AA+X8Ry+LQFSpHM9b8tqdflT/Jr2gGS0UsatcZ2TPwVeRk6uEnAu/bv3aMsOzS0JyWb/ety
sTh8V6A5/oAin+PdX9QoN6AXE4FIMnUu8YLyDeRMsl2L2dVJica1hFBpaPQJfuyg5VUX0m/+oBDG
iS5TGkCh3p1Tle3IeQzAu1Z7+28yrfgFY9Apmtzhy/z9sDXwEZzkIyZGnExDf+0ttOUBAtSfwiZv
vgVbK2yusgi11aB2EhVJOY98UAYmmAvTFRJnA2AS5UBURig7fOjso0wEBbpk9bGryxqlZheoTKC/
LeQcWghT/I3AptCUZ5XLJZebsk0WT+X0BPHPpY/SflCc/9dwwnnKT3UhmqQ6w95GvrMYyGi2q3v7
pLRCeWqZc5ABfSlUraUHWnNgCcBmewLqiMIVZ3pM0jiH7ted0ETb0/B2oFZxwMrtXmXBWmmSzJF2
As46kqQKEPeuip3hhmgdSD5nhOs7UFBnauxAu0efJ7g09x2hZPfYJAjzYTC2jDt39N+FTCOF2m2L
UPcQ9Ubm1qLLE8rfU0UaPHQeJiLYCV9Z6EPGFlIOza0R5O11nA2E0vZ4o2TrrXU9YqP0dpW/9zwJ
0E2tgYc/3swh4ikhrKFdR3aJRoz+7awuhS5whUsT2raTAYeUkdahlm4+1RUBBQA+4XsLmqOQ+OzN
Z2v51AJjE7/bRQd/lOYyrsXUxVSLx0adfxlj4YlKX7QlvTsG0lZKRa1gQi6oqiLDY8dcxmqEUEJW
PbDekE8N+LhG0vNpupuT3SbO9kbKwsj6uzrNxf31G/ndXcjA5i4a5Cu7wRXyGpEVeDXzuO5QcnPx
Y0HG5cFrSy37cBLBmBhaI3z5SdAyrMNj2RmjkhVGLxg3qVdDSEYiF+xq9zhq4JRE3Vc1G3KDvr/d
i3YHcD+9LFq3f5ioIdvb1j9u8tbhDCeqFcfrEksEXUw+1I4LE9mba+k0Ys04Bwyqtxkkxmjqe01H
0RW3FfnhdDoF4rFNWZAFaM9l9R7sfPXsg9iib1IrjkYMOWHE64EF7IANUzci0Ibsht6dajamQhiv
sKLx5817cpEgoMWyJUHU53/VDnH4NeWPm2ED+AtUUYdlOZrYX+68hsSz9QR4KiUQgmUPr8fh+2Xy
NczutpUoQ0MJOi9N6l2sAy33af/gV75TbUfodeScuobwfEVYF8s6ZbX6rQ7wU/TyeH0Mn7+/nb52
CREGXkBpo07ddYPrDVf86LmWKKnDKRHTv+mYy2+iW3K5qx1gVv7rufSScRttXdpfPlkrVauULeDE
k+0ENJ0Bn6wuGrlXXYz+EQZDge34yHRRxEMwHFRvVvlwLc+TrMWx/LRl7r4ynAtzhO5unDLdeB4t
QvZJxNMYpgdHr07C2OlpI0mtzoU1CMnTZZNROEnfGKTOvdZw62FfB20Lqls1ETA0XB6Z1ArV5hp+
gOGMCubhzaRhqJQtgcXs1rRv1eS5EM9WElLmpvXBDlSQdrzjFfodaO+Z7PeMmF08D5nDm4mIswX1
dL/BCAWLdtoYCfMhNLKv0BTmeHAo7FSMtbsvQd1qNF9SBUB/Hg2P6xZHrNnipzlb+/QrZumnjT03
0sp4GaGXxFvh4KmuuIN4MAiT/TuC7A0aRfqJ3lVVLveLut/cuBdam/6YQNmK7lIBUGGfF8KRUVyf
0RTo7lekaAOvAye+QSGBSZcmpDDvF88JDgGXVjFpi42mGlofPT7HFYuxO6KobN+pOaa5cl81L+8h
RbOBbPoazpUwMYnFcd6onlIDfCqswwDc0UYMdW8c3bMiARLUIDxvkjG1hByBNjsnUCpvWzDEZvNm
np2LsUQx4lHAgfexEwcIX+yfDn0jZoiPu3SD7VFPjMpMgxYdgoARgBdy1Yaq4ATUN8ugq6bNwqbq
Nrh6YPnyZmRgYZa9f6KK++8ybRfOufRmcvPYyoUvGOGS6B0jmEPhvxdxIt6lWpRwyrMdCsRTU5rU
2+CzUiteboK1M/T+Eg/QUrg1fOlzHuVi84aFCLmYw+1VFwaJ12o618MnMzOspwbTlSjK6g3ByOct
EGioIJ2qzDh+nU5q8YU/VsjxEuui68G3UpvhXO46ywST4k14peKR2i+MQgF2VKxq/822a7deDfEh
Q+TRFwGXVOTgnoxv8TJkEkpWInVEVPi9c98eyd90g8QQ0lasbQheXU9hqJpCGhRcatjEHM2J+wAb
PbzWoiYg2j3IH3RtO20yeKE47PzdRV1ZoTSOIOgkpphodPcLQTXDEAGUThHpEmvK4RtRwHDiMt+M
osJJTUY9bmQctxRU/5jtDSyi0pnSa4LsGfbANYjjmFzGTbZx0KzyCW7PbaJbpVZqT6XU8EmbqmHy
FEubdd4HQIEyOZvkerHQMecHGQF7ymqTjsDlMouYZXusCQbRrGVfPvDaU8dcB7Msql//6vUXe/Wr
9Xb5siaPI6TgWLuFJqO29z4HyrsMwn0Fclg4xk3/LSg0bvFBThsLAjmmty2dHFyxeBs880UENlFN
f2beNc+7MiY6Fk7pyQmyEtsDAJE76tC9S/H5c3pS7YX0IUF0gL0v9BXNuOsyvBbtzki3uHEA4tdC
Wy8TfL+mEJ/yBG3qLIflk179vtjjzxRykOA/QPbMrgo81lvqbv6ElpGz+N7Nj1Se9sS0HmkPP/zq
r59kTYCW+xVh1aHdkb6y/3H8SGabEAC8pZV322u5wj8EliHmk3ZyfULXCFOq60BPbsuLIdD5tQGN
toPGtj6+gaYwoOLG54wJ27UCz1cv+yGjVKJTbLTbYQa8JK79Kg6vvYw4Km24z5hPVtjEgNWC1Dx/
byJimE4tkhMLF+ff6S65uziLHaxBJGG4vD0AeSRaJ978JDSVfBiw84sjInuHOmhGHF8KAVIm9fKp
1XKrkvxqdBIJ1AY65nOZyaXrbmh9uvntEbIas6Hy1dGnVM8MLjuMOknvuy7MKX0DkOkwQgrwjvN1
4D+hM4OM3z6SI5MDCmHJ80wP/G9mrPHyNZ5IIgt7l3+1a6GVaJ7UYSz+87FxWSHQD67EOQqMCSk9
zQJT05NbtS2tO3PsXy6wFEwEX/WtV16gyR3K/QdgwZnHY2mGb0eRekBz7iwfm8RCnzjACDf6VgS4
40zgXk2Ntb9W2G59ihhes+36akpm6mlZXPeDRelJhlofotbsfMBzgtqbELhNMz6kHUTTHSGvDW6q
Ug1Mzgt9xG7/MEQQRoe/FyM08foDD28pu0+bm4Wrloo7a3ru1IqjIpP5bwjeAcV3EWdJa6sFL9kI
XtSfowEz9joYsUVLSXGT508FPYfr4ZgDOZCYLDJofLUR4PKRASTnSWjwf4uJJ/LsMhZERBVkaazS
LrxR6smSR0mwWrNHD8Q3MuZRkq0xRcLVXxDjTlfN4qtL6oUIbWuP9BNyvVPI4cyP0XSW2iM6fbFE
IP7jW5KXQd/hP6qx5b3kJWq6aKjbYtsc22QxlAmFRQn4+VD6Xb2dGZU+hpy1TDVntn0GDH/L6u0S
noXBhJhRpFxm+o4AyeHiNS23eRRpdpd+/aLcirIUJ7CUrY76z+AKj7N/9jlDNxlPU1VBMXGu0t5U
3fAW0G2+WiwETvVwSs33jj0qwn66zAFtxrzYdf5WakKIZThG/iuyKqJOSi62iq3BGtzAFZD0b4+t
pMJXhLB1hXtPvrizseKz3CqmVLXWePb3m7PYJ2X2l0ayQxqdB6IPJjtrDkwbJ77zI9EIV7/fAVY4
p6SJHAS8NW1h/SHprlxxQ7ZpOcGfRKlwx20h/QFUb7/hDaBQuev7pniDtiLGeAAD7I41Pca+UZ8s
onuqPDpEqOR1nEIqJNjOOYH4X0UwRKSvGzckSgzL7NkEi09WhmtVdJcFbva3Y5QQpmzxALzDky+3
iSqTHPXQ0q6NMpdRUdESbi4LFJuI6jnPmh5Li4KwZRf5qVHJCRqrebjFJYLWbtOTNLYL8cuPC1/V
jcfQGVL63svv3FbxEpfox55o0dCa+r3mXCwXMcE+/gbkj4FSWfQ8nMmQhLMMqK0Qy2COgeAcEiLc
bxnZqvArzSfysDcsWUsNMz0WU1BDlYd8Om039M8eu/TU2nEaU0prYRuHfbDgt132vygZEn0azm1z
8QEdJ2pHrgUCJwVqsB6sHDCXRWTAO3tJ0sL8FzwysFo3rqVOy0yfvTJ74LSzHhR35kQ12PItkDpJ
B5340pwzDgehPIJobd7XVtfX9szl4geR3UPw1bbgN1EjSkVglzLICuMI2NtuH8XGOsa9zssyMttZ
z2qBuu6f65UeE2XAqjStXdni65ePc77BomEyHptS8e3XiL+w1iYRQ/3KG0tubNkGmgBrpgPIBwjL
KA8wBV4BQlrOJ1V7Do5qtla43UteeUI2VsWtM79DurDSCU/eEOt0lWaqSZpGEvsEBp8lnNpB0955
hSELviO1vViNgWBuvDJzRmGSIyawdaYqiBPW4NBtnqaa259T4P9jFoKOzSNwpD7+eLLsQlcOo8bD
XXqyysQlqnCsSSWxZ3UVAojknNdYMDeIb+U6DG2H9XuIDEHGomNZMcPIfh3ZdkluFGPuSV7nfOHq
IDOk8w3etBCt3qoW/JZw/cRPExYwbBWqHKlD3dkLMvF/Pz3G50wSlZi3Mu0sMPJtmd4LAZpBKv1m
60KqkdCOwdxoYbJ0H9nnuRB+dJSXHA5z7a2Hc7MOivpY3KCNT58Sh0I1Dj92M3KP4aAX5cI9MLE8
L9u69j1yvcbg/T27XxhEYlUeovEQXKWthZQ9s/0Uu9GNsFcDpL2lafeuTZ4WXctXe9Zu/givdSoZ
EDv/5KrtxcgLPT3MQnmBQ74vmTNJIZ1B3KoPs5ItYcEDpO3I6/uRvPTEEkPBFkfpTT3fGsrO+3jR
cvExir122HkvDmlzX06+If7FVW6f4inCMWescvQs3WukHgx+mubxQfLBKcBS+alpwxsvZk65H6bj
22YQwn1zHpaG6YYscN1tU65gLQ/LTo4bZ1NFXvvtUrXJ23wRW3FsZM+i/bq84K4SQcd2K28Wc1uh
eAdANQGqz2x5wkZWlsYH51pAiCMfO2Lghh/MoGjWjzgBcV7cXVFRavP+IYwTI2RqTODvuOrsR2dl
Y5V92M3ei44RGBdOfd7nbkB9/T/2s5CoE/d8MJCq4eWqQGlnN4yHX3YvpRtqZCdtSg3+6sLvZ36f
GhU0rPKLCCbVxeNri5JGdcKq2Jpt68dOTKGHwp5Xtlwmr2+x7gl2Ext9uAu2UMvswpKBSeV8lxA5
Du9egrezePo2WwQ5PWB8QGArU6bExijArMJSuM9Zhgauc6DRv9D+6nuGy152ws+MASs/d7oEA2D9
OK4OCVUh7C07PafQjSXd8UM9h07aN7s/7fHmLRhUgB8GzH6v569it+DY777MQKw59Y1o2MwXhb33
g+EChEL0Daqo4ce1Kf6ssryBigzeBY08DxsoYaC1VDvQQMrOcogM+OYwbMqkqf+o27avpbYb8tNK
YEY/WmULJ/4aMU6/GUaTxZDlvbAmK16F82XdGNHqvBM7VoVfIGpfWhOT2iuQK6AV+pAIaikuAe4n
NmLUTLVt4cPRPCL21Z8FkGiwEAKwAOwrM1NwaXStPgY8JubmO406nvWY7V+GjWI0tAHegBfuyJRE
c/jQge1RHMiBHzYPhy3UdfI2l12GbnMbeqipIe2TNZLDQ+p4LuAfQC2R2c3tSekKO48rbaGNNFIQ
FRBXthMxNdV+cPw4U3LJKKmZSCAFPy8fagNnnAzQgMq6j8XWIoYcBSIk+4DZRKWpynScvIMxT5PW
Is25vV0DxqTGNUtaGd4yezLiVuyRqye8pE+QPLNPGYNM3GX0owV3otS2aCPV9N0d3bs/o0cWzMTa
KR3VqVDYpAprn84V2adFwwT4P3jgLhMo5A0eU5//IwPX2PawpFBibXl8ncDjAx0pUCcretLysI7v
tMEz3r6WOB9H6sqxmqPBb4sfnzhl7+Tqqhk9lDH85vb7lfktG5hNMFfEorgqCdNfC93KK5E5RAKB
5xkpo9lmr84b4KL1WjYmFTWGGdn58A1Sj3K38/i0PxzpMdM1DMB00cg32E4dQEi1FQ29GSFcezkL
IbB4XmQypimuf8NoLZTKMZk88W3WFh3vgMNnClAGQUn/t3kniGz4mnD2W9z103YPuq06TpqxeAbd
dXSGazOErBYf+d3KMC6OvxSXLRhSv/2So+k97iP0Bpr/3q05v5rKTjBC43J01sxNNAy1iX4ORMJk
ylnVX4MsQs1n0YjU54pgKHI084vp8TjpjKiRHHuKo037dgfQrmskNKlqtERSySG1wAubVTwedRL5
+TmNmLtPKNA4koZwiTRuUFXaGnkJlBDCf3DQaJ+AcM5BTCdS4TbBFOvPBVNW13BF8au67O9HM/2d
17hCZuKkE9l/r2K71fAtDsLT+9ZBBO19E/CnZ8gTJY1XnT6L7x7eB7ByZEavYObaC/sybcJiSBAs
BFTUmP4iG0K2m6AviSP89bqTsZjYfenJcUKiQMa3M0odRNFXvNDha41+Irv9i9nVuDFmyO9P4bV3
pwVivJ3TT70fBWW+tDO+54kieYJXj+RNWdFBrdw+g87Um8y0zYeujkv1pduUDq5G58BPm9qqdjot
1eNVwup3JdUU4YRuFFYpJaIEj7sU8mxCD5JShLqWc2Wut9oMx0IhdGLSw/C/BJIw/hSQiXzAgt0c
if7wznZRhsB0Dh87DF3JIWV/gY6+y450lcHRoPO9zhDtcq7xDuVre+JcnXBtEbDUNwXqjHq7SzLd
k0lw1BptZYbO7MVmebTEPu9l8KmeDXBJOnvroUcWxfwEN1ltNU34LpdrgTlL6epyehNk70QlsFmL
OB+2AZEAU6N1rAGpeIrBEkVbglmGshsr17dBenfUUypVKa/kQzUKkVOZLOZP51HBiurrckYKoiF6
a5k8EkmwlmDl1RzbHDTrSLFztG/I5qQHwmYrxo+YRPR7KcWcA12K8fMZMDAxMW0uIoVy89sJbqTe
Owpfd9riNb4vFY+AFdJTppiQSKJ7I/8+GVyc3gQ2asoI7iFSV2N2O0JxrOi+zc9wsXCT2u2gZj1K
x7UPJv+C+lksUSKrupTadM7goY98Uu+KWocBlj4KRyfsmgf+qFyTM4tZ6jRpg7swq9W1c9IRma4b
VLr/tuwjPOu13KYpD48Nt/jCjkoc7KPYpJ544lQYi38/PKpjq0GdwFT4xOLA1KZ5VA+fazdrAGt1
p41CyStoi1iuOtGAnDu2ZpWc01NSOeXs1hK+KflROk68J7sG0lzJPDDRd3heHRWCXcmVKHz1FsFs
pD6JvnkHJ2eCwdxnd/EaY/W+BJ8ZWWLgm6DLco9nXjLHQNFT+0gSUSze07qDNXsYACRoAvw2RWdH
Tnca/z0IJ2ZyVGNznqpBQqv+byVNGwP/ICbT7rCUqPIzLg6xb2QZgduDn9G4vQN3PIh75leKsIXe
TdWRSC/AqbV3tBOMJRiCZ6WfX+u1fWpu2gTrR+uozxQ1obYUM0TnU/jGtjrvbIhmROryg/mB/E9T
MI0Fx8QX6BqQXChYAmp6gMHc34NrUoBMm0L0PehhfiyRavOWc4RFZbFW9Go7KyNPX+9xZhyoo+eU
m40+RRbfYGkYHUYlpxd2ZyAWqo7PiYKF+AFlKJGhsD0YcawAcTR6mUVECyGrKAh8dthxMarpAnBZ
XNprBod+3hN2yDEcKwggMdooT0CABvsG2B4t25Rx3LtdZAGRUFXPOXRubajw64DoYeuoLkK0iJKJ
RDyhWmX56pmkple/WL3tZ59XWKwvs1LjQHrNg1c2pVBsxixkyJoneHyln9uKCA2V/iET6CR7Tj+S
nwX1w/kSWc3iASEzb2MuZJ902AWwaf8n4YkWFwC5ZH6HDjKVk/myu9YGWpTcZr66elUzn79axnxm
EXu7TC50Sl+YnI4dIDmALTT9Jxsm5H6L9rDkDyB38JNx1wanNBMg6jP20yJINE9I+RUiM2mPGy3M
/cRDgm0PjK+SCJPY2me0Tr8Sk5Qk8gblhX5lq1Sj8YSuc0rBYB6Lt9L3iI7pCGGhn8wFo7WYez96
nyOIZNHLoaH2gv+Hb+O92ML1cTejZ1WUTT8G/bdaAciXTG0u67x7OVhZIUm+84S1Oks1HrsHxaNk
/RKBC7MtRwjhrLpoINAy8mExo+3tJBic0oeD16QikYu/k4KpLQBet3aZJqdVdYjJEeEl/1XydgNV
rAR0AwZqaj3G62DyuG1G1ba5epp2w0JdnvSzn1tUi8CiRtWgzjDkkV6rtECwLe2Xc5BTufkPNZm1
4kEipRaEoYmyXEU+lXuqH35ZCtEXaXk7DevB/GvgpEn9mfvJ32obbUC9Ws+Z0AYsfEpR28CIiGBc
7D6J3HBvDwbf5K/CRGDNwU7Up3CQsJ72QAJIRJv3u8XCgcvYotzDm1s+IcRrZ4HahkKXHq7ziHtK
rX2YoPe2fjT+DXSlTU7+7/p/VqvRkZpq9tNfJI6PSnEdM7E2R9JgGbdHEDnOJmblbuaWkzPJfFya
jJ3z/QWjCNo0+w/RPnpmaia2jd2hnHz+dPNNKs9/pa0h27xBKEXnt0du5qOJvuBYUopkFOpgEOH5
d9dVz5IRHV2br284NC05k+o9aMh+2nHmw+3PD5Y09zHif3oC45qDnJEvQJZHbZE5RJNjTpR/Iy9r
dF1XUuxjADcvmLwGykOI9Sk0vh6SyuzZCgt6NSzGi/poKWL6eSLwqTKnEHr9GsHIyPXsNXvzC0cv
vVfKXBzCpHsRzqgFitV4qz/+FsgkTnSEz4Wke994k0ZPnOn/xRgV3PhiYnjczJReXnYR1KY0Le2l
nZQpvdsnYRFMTfC29xVWvK11pCHIPATz9seObDVPrGUUr5fcTe3XvTCE6o1y6PjIAfBAcr22nepP
oDY7H9QGl1dTnpb/1PuzM30NBvZVdJUSgqdErQZSxstDudCqh9KiJTmxzMzE5h9fHT+7EjV6LWEX
51pj83A6zwWAsu8tAYkjbjBsc4Vac4bJQCCxNKiNsdQOqUxlakH8caN9TlIMKD/isqdLwwlTtgiT
PHxdAr0I83xwhJvDvwatQ/VPMFehprm6eGU2kx3ew7ujGuBs1XRiwgWD/AmJ+C7ZWq+//dfb4mdr
ycvpHxiFZfaHP9UKBeISCKJJrbSthjB4HUBCNzIpQgAkTkSo74DB8/fE17vYrrpb3p+nTfJH+P4d
cH8MNb4F6ooQAbdbYxkyoRYadPulNUOSiKQfp3L9JEnksaWtIquGvAEgZjXh7HzRkn6HDkn5OKFY
M6dmnYhu2fE7cp6+QMFaB50HeU8EupEVv126uZKyj58s/FiXvhN2qh4lizT8Tm+nNKHyC49t4kV6
KSopZofdm77ifIpZdzJ3+FkTCgTVv36R0a7sydMwtCcvldQzY2WyQ+phQ+nyM2ZvF2S1kO5ceO4G
N3Aw1G8nlvo6PRpBAcZ7k44QTbL+1Ng7UxVPt9lEotUWIOlLf93cieB3GgZidsqXa+tE6SKK0+es
Vb1b/a6cackPzNi/5Xi0PzMRy14D1NLeHjXirt0beTx54mPXYpxcpvXtRtsxg1pXsqKEcvrIOitL
JUyWvs6SFIdkmdD5IhsRxv5sONa0UBwOjBFpA6SGOn9+9sHuadK5ycDOMbiwU2vYFiPi9VNpYUXb
EWeh3tSMclQM5m9vxheLB/Ap6PwbGtcgqvo2q0xFEJBWuKHtYobrw5poA2SFE9XIJ2juGoHalG1k
oB/uufg4zIR0aqJxHfq5Lbx+uYyK/7gIMSijdFmtDwKvmzCl4kXXK8p5vAZtCXWQo9WgHRj3xEOI
2dR3pe1TuOUtv45DYeOm5NOaugae5L7fqAaKAwzR/p0zhapo5OrTG28BhaTrBF/GkLDDRP20dvsY
sDJwnqIcZmO5lT1Rbe5eXc7LrCGEdmX8lnlTyGYHe7KXhFB49DcVm6fjac0UprOHYkOpHvl/i7Bz
rQ2+fkHiALKqD61juSukWL9EWDWgrWhzM0RYAhtL0R7B7BnR9agI+y9QPEBGS6Hm1I2MOnTfnM6W
5LX9KNrW6T5FfFtM7vY2semy8znPnFXKt/PzD+ueoHCf1LghygZHIAIAxqU7qui30gKrtFVUVkaa
9qKY/pMmkoHETsosZKDDY8Wp8O2BzDEv5YxmfmcOf5lk7DpBRR3paVGPZn908oKarn/UO0cZ8iQ0
mUdcqawAl7xlR4LKsVWelxyMEEHKSkRXlei/cp2eKYXuImkhsHusgZpFvvaOU5Kqg0X6bcGsas/J
07crB7s7xwLLf+PdeGxp3NYGK8kAfAQaMxYoVmFGK8wve/D/1VJzdeA/F/csaj9hFII7BIGrjXn8
4q+N9Lcr33B+sM2CVPznt+B9diktrwi3JfJ3ZL9dv4lSMtoPA3lMl9KUGGJXtQ/MMtrFP/9xdfbE
pla9a9KlF4VPXPHKEDLZZ5xh99lX2hadYkS9MF1iaGvzIsI3bcp14hzrPM+Snp8m40byJVcqFeEP
4O42qwuJek/K9W2oDQswZPbWs2XLB0CmFitZWt8jxmHzXHjeRD8kqDUszz5i8ySvKy2ywdzKfOu6
NT82kWkYQSihTY7kaxtb2QWpVh8dvN8Pjiv5+HvEkAPEd0CpcAz3FnBAYpx2+3cv0gf5mWcCGQWo
RMMdsI4sUbX9bCCnM6zKis2wIexf/U50bBxC1SpH96JK8MJKiHYTjkd4x4pfS4YMFwRcxMLcpfM3
iYES4/UPvL09vD+8++mQS7CWo3fyGEgPhPIpi5SjpgcdvNmSQ0+wISW2+OmB51tps32HO83jvrQy
WBzG2nBi0oZbM+VGuklsxbY95riwTcig+wi5cNyUpztEB8hq8PfntSNqgysMyrhHQvGb+o4t/W9q
V5UGBTwiCtkfWKvcp1cdwBE6WNLtEUJ6EXyzedY77gviSimlt31ZvT9VnARFfcVB2BTZgRd0puX2
O7RwJsiC/GctofQdcj3AwIW4y2QWY7gNDIDYTCy85CuLvYPudK3pM+pCqhsan8M+z3VdCSbVO5CZ
Pa3lFv93djdVJE7FDtCMa7uS1bOn6jh49+y7kAprkBviHSwsK2QQuj4eMnMYTgYm4KiT1dMIZqOx
2YPcQ57PmVbeBoEph/sHEObWIRB2t7qzv/F8MGBwPw71ldtByi7cyOb5vkbJS9/676PtjM4dpN8N
XMc0N0LaO81ob52bQFMCGR8NjRGVj545tgleO5yK0CgbuXN+Z4UPU27mPNHsJScpjwEGlhZZ6mFh
x1fZsV0scE8eRtjTr3oO2hhuv7Jji117Qg/M/Zh3A0/MzC77oZ/jqizjC/dJt7BoGLo3+G9zhJ0D
byFpdit2CLP/cs/RehAkFdCwibYRe/O/G0vCSq1V24VTu4Y7kdpTvmDNoLNHtqHzOJBH+57XfhTL
KIOcr7pbuiFZEPMRRi/SFZ86Cz2xD19rMZbD/BBwnPkygIIypqXLMbFCb6JhsDeIr1Io8QaA81Dq
lSAunjbA4flPck/rCyHPR/+UIaSljhpsm80ZgslMkFdKXYfUEFz3meBKP963CN+VQNPTiN6ipk2A
HWwVYCiNUSlzTJDOp7K04qw/Ih3WUEe9PoEPbYqGuNjhnATE+CwgQsdwn+4Jahxwe2wKn/6Kx8Sk
Nz955MlKjqG70no9xMMSby19jVjeNtsjz8ios+3K/hJzRQzRxj5uzxiX5ve8ni+QHMWtvnenjASJ
D3Au3t3nSoJL9t6Pa+z+Z7ZszoBZSJy/8MP0AbLobGYNVxE3ptwPLNSAafkCh76NfFx6wA3zD6Ev
epRYXNIQfC3UA5bSUHZT5CUTWf7hroTRtnzEdhwM7ii95SH1U2xrgES8dFpXp8w8QaonCfCFSnkf
9QAgplgggosPl36mq3kIMp2pMOvIh6W4q86bVasOrSlCZhBIZ4R06Zk3DoZ70CkPEEKol/GQ0Hka
d6PaUP0IcRuLND9djCkcScfYa6CQ3Sn65tGzA+b4/6fw8b5aEChgk392vUmslXORUNSvyO8gCRRS
eJCg2Qy8MVmx9Enz1J81NpkeemxXZUL7Lzxg/ZDzbcSxofSlxFIpVTGvstxwH3jhXUjP/g1rQYYw
iwUdcwjY/uqFa/Ft9m4sctunOaz4ead51kP1TGluuaYDG1EslBgKwUYxwjRRa7PcrMtwVNNHHU2t
SejG6izADGnt2Bbi/uWearT7sGCcOCH7Luvr/tOu9nC3IZNwFZdzy+q7ZszWKp5nXMobIY5KCwwQ
QtnbcEk3FyAGUhiqSGHRl/DkxkY372W6E6r1tGDaB/ZZYzXzAc78yAW2FUnFrda4EUed5IWhfZiG
3ZwFND/xG87p9hqJiI4mRl/Ftlsum7KlKFEFSiQi3oumWRMF6GbBuJYobp8tDZf60hvWKDUW15I7
8kpV8RrI5TexC2Qm/S1ZiRCmq9tQv+1PwQXf3IRrSZrcP5v9sShWWWLunqZkkgyT0pNsQE+6GtZ1
FqFohbUKUmX9PkjPAPyAm7V5eEOhGJ84cco/DUVfuS3tvOukU8dSiqHyj0qDgZaqse+Ulf6kM2Rq
3Y3uN2kBm9jTFWk9ujKO37sbCaEV0hjio9MRy0yjVg1TEOYC2AQxzSWQW9N3kY/IdAYvXZv66oV2
qMHOZhF2MS4NqfJr5drANMnITZWJnKoX1CXjx1ll38n6oleJEJNAp2+UIQpAirZ8BNAzcpbAKM9x
IcKXyECPE9B1MAs/NbiISkTpED2xSAp0DZeJKwJc89d+ST7froijYx8+yt6ugUF9jKkdbfWWOLTt
HeBYsn9W+/rJvNlaHPXYPUM5Q/tmZklPcVkV8WBJPeZEn2qJcxj1opg8WxDJAxaspzciXa+RWpK8
Dqeez5hST7my1uVvGsxdKhHT0XK+VY8/udzBbYeAj6m4jXrV6UQPUhjoG37gwuleQiIyOfwQNvem
MygYJk6Kobk5ttmrqQI+UlEQ7ZHCe98Q5NMTIGQAfvXsnsh3XXSfTcmYcyMfxErpIZaQStney4fa
q+QcNRzz+ioOc31cg9LyCqyXmIE7fXChBZtYABpZLUNwUvAFB0vFBaMqArBY2wsJer4vk21GiQGd
JiUV0v7Q232neu7ion9FBVtvVByJe0IFCG/54Dc8aDNObP435NoR2nIMrxRtphUBumIXMfwlxIrZ
OL0leSSHdq/yMRt12iuh+xHtk++pX8HFDXu4CbprUjGsmkiESW7jTk5+8uumNbILgw0qauJT/ev+
LZygBDiif/7yFzc2jrKeOQPXFz9NGhixmyCGjx0jx+AnDo0e3YctWO0qa6Bn0rsIWgtcNawCVqCd
y49/XHyxD3bJLnBCwK2OjjrHxt1F+tYkmzMJ1UDS+79qhMyU+0ljUuW/CotajCWojuKFCxdRCUpD
FWUeJ8LelyotTnftbAPdeK0mGj2T1UOjE98rd0BG5JHOOhNY/GHWMFHX0fboE0qGP0/1F+cC4q2U
ZSV19KNUcmMEPMmA/jhPArJZ5APq3zR2ws5UQuNjPtYkGsqFGah+pmCUrdt+JNQCIgTlGhm5t470
w1KEllxyBRL14P16IBFpmVhbGi5yDoKEz+ws54y/dOo0G2W9cGOUAmhs9oW1SfXQekyXPc27eh/e
BLsBD1N4wLHYHf/2hXtsQrZbtNprEkASZGLCPjbCP9GMCXf8GVhP/Ynu6NTcMdA8Mkr2plCKfgsV
382oBkcfJE0sqBBPmggI0+VbtJST7qQpW2FzTEZSLtu+hwhKUIc2igWBp2jGyCdee41k6wMLm1fn
N8Pq7NjYUxY0tETbEBlh/bZn+8VoC54Fy/Z0dWpeqaSyBEOiXmBOYsN3ZO4eUELegJDC8taUp9RN
sInJunZ6x19jvQza3A1eF9sYwS0DJ9736SY6e25vZYdrWl1XVYSTr6t25RlxtmfL1J7n3qu32P4c
CSISbcZYzMxteXPiqeY4e18KLK4fLFzwFsKfrbJIK8IyOHse1XOeUFXpI1ZxkuHs5aMAxDTBb11C
AvtL2HWVCYAHOvW0hPpuxVXNEMjIxQxUqvcjDBscTCEQ/JFL7bzY12KWUh0fz/0/FDdWzFR+lFpP
rV5H2dA1WHBBVnR1nXKWeuy84TESgOEchPcPr7jqUxMslpqrGgGrdka9c6W6AIF73RBPlyBAnrgS
DINPrDb9CT9Auz1LBI4WE/B8Uuys1ghbVu5SUUWWf/aXt/DPI9+75rNi/Q7kuOvH/NBc/yCbtZGJ
Fa3tNwljTdOkVJwSw1Bu9C6IraKsg0ifkLQSOnAdncT8p6oQGUnVVHvYmAMfGKKV99wEmAfyvCf+
XZRLQBb8MT86QG57WTk4mq7RhddkQAfZY9JS3DHKKI4DTyfBFNnqkfXbmdvTM1m4uhwmndnlTeTI
a8qVLpfg+bSALvq5wMU2/A1jZxncfYl3gcGpPtfS8pItjOYC+v6XFVPotNLnRKMkhM3+My5MY03N
B8Rj0MwPSUhTPFpKInk2AMiiXvrNEFKR+1gTLpQqD0IT601IuGa4fz3m3VgBoAeNUE9O+KRzb/fL
FaUK53n4P2+5LA91fEKqSvet5/1op/T+EFROOkYYfwXwL5/fuR826R27GBhsqwTkbVsIwQX2s/Ch
7t2Ju0NrUwCMcLcwxovedHqbJnQwdDgL1noV9O5wWurZHrk2tGONducPCzWgEnhJFOkn/aGnOxRM
TlktHQcBYEIZT2IhuSIYozx39AEoXyMtxHuHmDHxOILWZGzIfsPc0YLHhWg91FI7/9tUKuZlcg3N
X1hvp80ZtQ3x4FxY5D+pHoo5jf0Om8b5ZqCloapx4nblkDGeNLNphIgPCWVm5wJbMsSZxBFKGJxH
LSwTTry0z/FNdN7X0Iy/jFUpctpX6s7OJJbJh+a++kFMRu7MR7I0BLxj80w6Sw0VWkmvqv4fgLzI
SDN7b8tIpBNDcARF+9XuZ+W3pt6h3yx9yIznV4NfPnAejQk85A1FkkoHfoHoEZQfCVcn8yTm3mQp
U+uWOTs0vQZeh2oqfGq7l2aLZMei/aelpLNRjaYD70nlpGotweddxQ7CnQb8ijVVG8PZOYBTmDvj
fRD2w7qykgwImzJAb9Xrsu85qgSRaA3eUCay2ZFjNiLgIZ6cvwCeEeGy7PIuK/QKy+IcjCq8X7+J
dlIjvFhRiYDeYo41/fDbZHeuIg6sXml8KoXdU5h4RNeqWec3DtPazR0uPOf4SxhykC/sCyfGsgBl
T3lWB8c7N030CwyCT2EPFJ/PQW/HkyMBxroUIQ9FyDz6b+h57YylKkZkPg/qIFMBo776eSHSv4RQ
lmEqoQ98A9era4lvaqw2Qbt+64no9jaxynr0Q+uFbky99IwMThuoH1S25SkFC8UBOFppPpcLMWGq
lXH4V1PxOxosMds77tcxKnt1SNq2JiwdYz/mZpfIv9SP3yHMiYxTXOmRNGSyEYgPB0iN75HdUdwl
GHwqFgkX62K95n/bJFLkdzx/N2NJfm/AxbGt+xaELeEvGlaZtDuSHlv4a8PniYnZGM6pn3yty2Ey
Ev7OdwTlovDul/KjYQENGlWa+qyHLKIWzq/KPDqm7glINnt/77FJLTb3g5mwbj/1W2XQWBIvgHwS
S3qgCNy7s+1TSLg8l7WBam1eoAgMOTkBVOTNiJdtB21vI9WPWFDzRKy7zJqtxR77WjtbFa4rzmxi
Z8BoA3W5rq8J9Am4F5pbRs7puF4qEGxt8ULn/vbj6U+DxA+gvPY89+S7/1zJFUcfQiraNIxJdIBR
NQBrEVv27kGJBucTyvhXVzkZ4uGNgiqjV7NRx6HaIvJUoj3o1/Ek3kaqXM6ichme9PpgLMXF9lQ4
tnwbR6j1pWZjGti8XUrNIAvVTdTBtOr8NLJGCPB/h2DDlcw8KwxZx3dGgaoOEaWLmRO2YABpsIm4
4Yoamtz3oxwCHRyGgRnq2Y+aUiRvQvKzOTz68/n3iGT10yz1+jB9+ledqedU3wWANzDmbmkNhM18
UWu0F/jzhhk9XJN/Fm3VqVdMnBcx7Wm5a0FPeB4ovfpmJkYO1/kVvGqfz1e270pYZAqitHhuBMob
8w2WZ4r8q4zgGHMws7At9ey7Ex3Ywm3KACN1slWxOZzEoeXCdmJkko9rpmm6Tt8+Qk2i/r8I2eXK
2baRRYQLYsFFboTLZdulS8aJZxN1tXTgkAbJX6gJtkXWZ6VmjccozSjhQRq30IHHHxAuSwJ5h8Kf
AWvOWXVVY7mr2LxMMLCwiqvq5CVvcYptffOXj5zr2rpJbCu7BKTChp3CS7WBfEkY2jLg3QEa2XXE
HzgiC6YnzN1KcjmEo9zlB/4eqMCrVyjZlmw/0rYNKs3/7EpnFLbX6o53sYg65QJBj1l5+lTICVHr
O5T4GuFsULG2fTiX5mWPM/vuU7CloSAMXRZP+T/PRxOID0IbNBPa0yWTAWHP3NKxnoX9ERXaLvrp
gtDTrbs9a5qUsCpL6+OforBZomdpoBqtAApr+W/LclZnffrYk6DGKxTV2oyNUH1ZHCvsPZe5fAvl
ootAUsKI+aSnaKjBiE8C2lwXgAciNycBPoOy43Kb2cfhTZIZ2YU+xJtmtfHtgbTtU20eUn6YUgDC
Mapg4Q54qZDfDnLp5wHEKUQ1snjrxY2sliEm2nV8ehXyGvylOWkKlKbcStKmnclnqxkdvsUAEgGw
Cd6gbY21mCPlW4mj2RR0Fjy6sHiDe4LTYj1yDjIL0mjULGid0wKyGaeBRRBS1gASLwGhlQODBib1
amjbW6Fcepd+kYH0n7xOGV5hl42e4phUwyO25TWQ30kZJ96TrJgh1jMnmKITZke8k6PexhqXuc71
AoWcj6Jxt20AYkojL/Z4pCucod6rl/juvl8MCjQnBwJPx/Or37l3h0IiIXG1ygKtP7PDwbYyzrnP
ZS2pFleBbxS/OOv1AYCZNAAL7Fq8qE5kTQ3+sAENdU781qg/WnrUEZ32CCkkDY1xOy8wLHLVb9oN
bItFJZfwPeIa43Wa6FMSwH6G1tCCspMGfYwgFggxSrJBubGQ7Hh0vbgpk88XDKS0f4urjAiF2DoQ
WMD9hFAb+2kmPQWPTh1WFaj8+m8BqVfD7OdKxXUpyfyFj9C2bZv90dwefsVFhMGh8Yyj4sDBFQz7
6zaG7QinIWel1NHrJsHHO00B94+BQ8ohsizLFrbtZWUeG7GFl7VodpGBq55StJz9Y+s2c0kfJjpH
jNtfWYu7+o/7MQLSINrM926Q3Q/WDIJJR1eGjQl5PaUK/WwnE8Y8tZsPGKqZUVn52bFC6Vl1xgDJ
6RfLlNKUSqOdP6KiGd1wnjGsHWKXIWBZiFskWQLyBIMmjJv288J1mzHeJXbvUueQtOwXzspBzJmF
/h4eAVaj8MHcK/JRQeiL6DTlXovzFqSwcoueJbsP+4rvGx9t3akl3oIaq4I8ue41mFHOjG1Z+ikJ
qtLbLVuLlWdNKlU/YQoOyQrJ1Z1FcHWPbegIbdX+ry4dFptg64B9/Ap/we6Tq2X78YKchyhucDoX
XJTXhYhwvJQTaW+Mfz4FsEl0yTcxrMQoWZ5semcN1MuRUrgVSz8Xfj8m8Gp+6paRuosULqvgGHvC
ZdXfcOv+CXhxvkvb1jFVr7uR4FIva/G/yJuaU1SqxOLOQ8ShfJ4cBMa+bHMbhtEWryh3IQaBz+pm
4tkFmRMf5KWlSK3G0n6Bu6W5ZPY+SiMqVC5U0JjY0JTc10XRNJ7ZUgdG1nQNEymgaUvBtbvN183t
IuubzCYSadz8gD3q+84zseUHWHKpQb7TyA1yVBEcIwL4xhqZZRuCaq5z+o4ftQm3VfzGSGRTw/Rq
lNOJ2ZM3szTH/wby7KlDAN+6+XYYqcym9js3WvayVawv+LnZ29o5fVhsBSIBLr78wF7/yU/7yKvo
3QA9PrT+zz/Vk0DzfWkBkXIcZtke4etJwwGAMvvIOwcBFxmxtqzwGlFjuVZQmTUyIer8DDdspAVY
d1rU9JqkKvpanIZSaWzPMgfHoaEbAFa9S9YRZqDVrONMgXbTMdFkdNtNRfZnwx2m+K1R5Ejwrr7w
6e0qz5sqOTgaphtkRKyOuYrxbl0sMeCJlh6F1q8upQAwJaGtdKMFdYs03T4colD5tuVdCDkik67y
m42kqBIIUsCvRNVvdmeh7xZnXGoma/NnjQVuRXlHXJbpKBiMx/gWfmRswzgc3+v+B+3vgarNsaci
KN/XGiTPAfpPx6P/RDjTJM0rPaDePvYoy6qIXzg4XZ1EFNiRd8Zg7IpSrBAKwTU5ezWjff8ZHCYi
mE0seTvUcDwddGPIEYi5YK/PYxRm44I9JY8Nn6O5kWMojwUk+jZuTqioELsdLcQzzdKRqECnXTfN
uSzsjNB8lppLyzZAoEIWnIAMPWwTQ8kaY8pg1K3PVjw5IlAKuQijHVQtiiqAM3eUhaRI2SJrQzqH
i8ptPxzAZlZzntAIQpEgfpZd+0feQyc4Qt7zpr0bPoojsZmVvehn448/zJb9kSLU4oeYURgcoQAU
WlFq0sHgDRSO9As25T4hO0mKcyJmIaus+Pl9TkrrROIIaF2K3QHBlI29MbRv4mhkWVKzUltOrb2Q
/z5N/5ymv9QR1KIZ//V/FdcVCBuy7PVEAxz3VFFfnuGqgnrqEfCNiGa+yfKsMbf2rNyIUMmVrOwO
QCS5T/vNF5KKViP3sVlliUdoviVnY5kJfFUrvJZiCKtOg8GP94seJ9K9RSBUh2YwNSbg5qunORfC
IcUf9Ve7cedvTSWG/Jhj8q+MMr3aouwe4/XVxGr7BOIcrElHBEN1JOh7c16f1yKdjItnNk+QBx4f
5HpV9lGWY3N2nkVteyumlRZD0oNFPBqVCK5C8yJoNFeSULUqrvo9wqir2bpabBd5UH1jeqB0W3NJ
MV366XhrluLfGoougN+XnETtwfLBdMvfFoZJ5ktoWt9QVE1ccg5OKFjYdI6GkaS3VumYJAbk7HwN
U7JYlAmpVHoM/DUDG0Pq978XOUFPVsaVQTAqS+B1D8yzxImaNfDkOdMozDbDrWceuH64pNBVRVFc
WVTRYDdmSMIdqRnvXMlINtT8S0SKxLy+7MvrjPJX9C4ldpeB41gEwi5qdaCeIiE88PsJ8Oj+OOYw
jr+t28PxgWw04vXHQzMJFZAwsJWYGxGawvOBh/CYYF4ZVwx88zzbn25Na8KirRlytScm9lcI13Is
4DgjajlFZioDeztBdBa/ox5wUKAhguFS9MLH7rFO4mhG33dxnjTcch3lLdqF9Nt3KZZpGrTG2s7J
x86rQSBY3XhT2IXWe1niTAmCKY/m4dd9JfwJHxwvH40hsYcdj+MlfYSK9Kg33QZtB6eMfbDXsyfs
LMSsk278ML7mW5NtrKsTTgfY2sWQv2/DPLNYX/lHK7+ncHN4ZAVWqlhIGBBRP1pGinZk5REB6Rhy
F72PX8CXnK31etEdoiJZPyYeU8sjFnczF2P40rI8vZj5csm1OFlmS9n/04s4YzHQdjdBQBOzc2hT
6JUctuqw7C2T6z0PoCNgVwO0UxQnezM5pNqmnbHHxv9Ve+LMVXhp7ptbav4/6vdSIn8j6AlUA0Jp
zH++CfMFfJlqMswrCCUCuz3/BGC5Czjx5Xs+iiknhlNZGaiEnzQQjxELR98J3e07hoVg6EI6UzIp
3Fl8KUgIalCVbeBq5n7HMUXrD+DqHSS/27K20V92ZiA0B7L8a0MkswXvqj4odWQWWbfvc2UELHXg
MldXpETK1zTsmCVcGnI18nCrURtqfVbN91w2r+w369nxBdE/X9pRAdGq9HR5VmkWQzQmG01iUVvq
eFo9kznAhZ1NpMvrwiKdLxt5+Dh4kdzswtXH5ooP8D3Jz1tVAamIcZdb6JD/TWbQ5HYVyj038eUO
8hh+1pshFRRdLo+FjS9AxMkDxBcLc9bpU1YnA0IC80uVmmT0P2mWjKXIj7gXvMQ9A6LWj+Ts7J7v
GoJLifaEH1sZUSJqBZHaI8+MlP6p6WD07WA8RcBdrd/4aOkvHZIXYTLC/Kfqivy/AaUlEN+KKvGN
P+qLnN7F74pcQrxZGbmffrqnuKjP7gePQVefZIQJCNpT7y3YBmvBOfsU8WZMs4M1DihIjcihwjig
8RYpi1hpU9yG10SfLqicfC7A+JZD2wG6gNt+/+X9PSCMl8KB1kbbtvOLaSZsRVb+rhScSigBtoZr
xeYtEGNXJRDJZZxF8Qo2uNjGxtSdGi1dA7bl71UWsNKQLLRegJTexOYd1Yxq90dEPhHII1iW1zpL
f3cpz3WJvaVvkkvBYg/a2QZvLWYBQlqtCVIWgUFROkHnvmW8VUaTdObcTRdPx4ehbfGHDfxxBGqK
NKgTth2uVm2Jpi8oU4iDfJb+4pHkMijlor/4q9sylzpEMI7A+9aPNN6glrEMnevI9toRtnoWSRtf
09kwUUaI5SeIzOUzQU0+GOl0CUa7Yj5VkXyHc82bOpf7xHR5NB63wDHFaXL3gvW0Gf/WKLglvTg1
Kk3Ki+QiBWsb2drtqBXx25Nag51GbErkG8YzMq6wVrxqyvRizusNwF647lp+MuisuoDuphT8vNwE
+LOWF93H9oq3IWHc+cN6opmGVOP7fxxrmWD7SsuCqUClxAO4K1K6K2YTm6GWhX9W/r8Mt7H5/qr5
5noQRELkYrSHlGIAnzXpDk0UAvZsj2Lv6zrmQeR/9/+Be3b+Bt934DWh+t4NQ5lTmBFc8M4LjlbV
hPO1dR3yDZ/lVMG4Z6sh3/iG6g7/lFupBTMUfj9xZ5Hkv4BIy5cpurcGAktQg2An3zLsPW33tELt
Y91G/8AMMq8yLj/QHZAAxinwk5M+IkPm918g71nLsS4iYoYYrzKWO7PC+tY2k2TGHOLni4cqYcu7
fXoALMEbDg5zozi9lWsKt4PGJfQR2sLJ5/MoBs4ygwoDB4DDXwlRCmnrXl6h927amhzPjhwsxmeY
FugU9z7QohPkAwGj5kXvBw29SbgGOo5o2g4MNkK5Yt5twzgaz0Vu/VSatSrhduq9pJy+GXZxcxKc
y1kdseek15Pyq2z7QNePX+1g9zSR8tm1rSbIMSflK5eYxrZRGxd2Dei3dit/WChcDr8HE1+oNhaz
FjsM92XJjvJXmC0GCn+zNjoxBnqco1YAwRT/0yNEFXflwHUowacydjdm7+OLZuHaZn95o630uSOi
uvWkX5z33u/hmRvz3YpP1/zM5C0oJO6BxGflsk+Ibf/WbCjB0mwOSuBRwmviToM7DJPe46SRNdmn
HaehZg0R0XLEXYXv80Hm+H+2gr3RIrx33JKDulBmqAbR18wQy7NXKwUl4MjKor5KyWWTD54afgRE
Fu53DH/a8/4lWins75eM3YGJvzEV1NMPkmS7fH6232dDe0Kpn+Ngl+FP5RX9BMyj/B/OKBAWLvvX
MwByCoaIve0pSpfJW1Y9XNAo40Ke466lDwya3c/lMRP+7uBTQeQgweuYlbXE1qYUlrPeXZ5QUuZs
iQIXnaMfFS8BYLYz01+ALvUFAcOz/LGCqy8FKxTFodb1cORC/dkbtgOp8Hf6/qHne5DfQmmBve5T
MUBwJwyt/wuktfkKMXIWfKAT2s2Vl/Jc177Jkl2C9Qsg/z66LXaLStDCDF2nHTkQgAkZmRSOUXRi
14+9FKWt9hUyac36jTMi53AjQOzjptBQ77HJ7uOh1ORD9rVcuqL3dVrrzKsxkxI2PfzZayDnorbP
NnA5kL5BeBSuyLDH8VFFdH1HaYFuOZ0mLVDLzhijcr9VvyXLjV1aHEaTuCn//w/nVS8aHhfjWZxV
CpRYaXmyUoMYDQsmDy10mrT00IkB9PCZ5jnvQI6dprON88uOg5c9Ym1JtBF/ZkVJfzmkopWzrGoC
WnVv2BuKpeMKR0ODHQywODjd4JzyewgfvHEpaX7UPqNUUucJXT8PXyBw4QsmCDmA0jLygUoGmhC8
qHG3AkHInJ1st1iyzYTjpn8nYl/Z1clGOkUwngUtY/ez8Q4d84v7hmYwfmjw2SeW/7Mi6D8bXTZC
t6J516DVV1mJqvDkfWT8j0S7L9Xxrl6SX2tDPBIHhf5DuVzY+z3o9fmv/HrsO1yXKzslDjXrOJ4m
pakVXk6NZyJ3BEjgxUTrUPgo2AKL/BdBsD+SSH3IipTMtsCoPK7zXCwqVg0PEE9rGpSskHJkpb3Z
DrxUE3+qlPFVvUwL8M7xQ9hkhNq/rDHfN0L3q1arj5N/N8W3V7l+Kabb5q+1g3XSV36cp19EhsSD
nJ78Gr2BNoYOc/VfQmjTzI2tq9Ive8ZO/8ImwjmnQCo//fHgiSbZoas9v2c39n7xwV3CLAXoe3GP
Ag86h22/X96AKoYW/aTQfBj9Q3g3k1dHYQZTDMBEWN/azlVP94+AiXFiY3ZLTCFMXEoPeJlvamew
l8AEd/JyM+remDt7UlhoJqUR2w/X3OnzspeI5XZLmZv/zOr0GStQMh00+226EEvs/cYXovZ9MF6Y
kc59jVQ/cIMN342xjCyQUfcCjrpieYYkAf5WQ+bxZH356B9IocTONn5nboo/Am91SZX3MoHncaUB
NnW8KE036yPvnwSxiX+sl/yNSKXd3EbTESBJgxUM8YmPuHL5ajVDFjixitfNt75eX5+Lg8Wn7VQp
Q4iEVRjLGrvGYIJL+fp82CLrsAKoy439jPA83ybI9qR2QPVylmf9AZ0ngXCeOmCNg7q3JeaKO8y/
qG68jbYRI4mhieRwJuNzCgLrs3ncYwvyy+cIdGTQBchQnXnZSjetGtgd4KCJ5SughL/YrMo7VhAh
VZtWVeKWlF3WCWmdoijEETvlqlFYmlHbK+j01bQPDol5NO2pIh9ryKmS3VU7/8LoBa0MLHZdbeEI
7TfWG0h888GM7X9+NKp00TEs0LpbdNf1tPjs3JD3sgouicqwHRe6ngp4SQOkUKrE2YApb2pvqXH3
EeiwPgUAnenAdP7FR/eGDxDaaNClOgGvs/yamnXcb+w7gAQKUy0C4jwEZlD+q1ssPJjUgxIef/9+
Gv8QUK6HtxPYNzMj/dsLpFDic6g2BB4C846mvPvoyfu53kyC50TUD9MoRGFVUnhQSyN8jh2fnLQh
Q8zlxS0FsmCZl52GVOeaT4yC3TU7J+Sh5VkXsTw43vwyGw/DMCfHHiKwT7jRFcTECjy/9r7t/Z9s
GztYjKdv2oDgBPFo9xDTWxJ/IeqamJaOOumbe4V0LkQvpjeUIV9Nx/HtGgQuAhWDBbFYAGz4M/I0
QrXbdRcLjyIHEi0kELjqUfM5vdukO/x1cHtiDprIzuTe7pWUk/MJVPIbRP9miaxK/a/nlRKr8Zly
fFFWQf2+ZE/8ZvzhC3e2EaykGM1klwo3ZG2xmGDjAP/WeNW+IdKs/x+96DCg9KxFPhw8zAgPwp5S
USI+WpF+Z8TidjgOKdF/55g3fYMWHsHtNo/jpeMuNdOgzFpMycU5QtXRvRFlcSLyboRn8Rji+W3k
k4HSfnDOpNUr71NeFdVwKDMSEr7IgWxz19qL7ejBGDRyVQLu9acgLqyk73XNXSeMSCaLZcXKwpJM
oY3ns4Gn0fT5M+To6gNQYr8LOtEPU4VaSLjdWdMF9dWi0/qNyFg9J51PfErwaKsaT/nnZZ4ipk3Y
MCB9PlN22JItCh6olcT2iKGjyZ0IWeUvXrzeWJiMphPnehf26+M3lFSztVrNCIsIgAIY9XI7hJlE
TYmAsNJNho6HSYIcMNHFXbl/oNWiZ+uZO9bx3li2CLPigdtEMIsr8tOOQgBpzFUUtTgFwFMLjTEu
glSHAKIRj5/65peLbzGYnqKe0JrjFm/+Rtj1hnRfZnwCFKLK56mX+xDOF2m3XloebFo7TRCm8a3a
mXDA7AyKl6BlW0TXYZr0vmiqmCJBrqEB3rN9tHAG27okl0COgFmAuGNNFGWKIEMDbp30pBj1A16u
n1TRi3naAKMl+u6hrWRrO7+DqvTRySI6HdJWN2JRdxM+wdqhq+QCiI12qchTRg7cqzZ1QBwntCwQ
QVNhyCi4qYDHbf6ty5d2c43lhZoKSqtCaWoafkiDc/A6mWwjr2dvNQFuqjVpAicCV8P/4s36NnU+
H0Wb0a+ocL/GxD94s/cv0NZ3RtW4ccIw5x6lzH7Zgt9OvRI1wgXDxaaylaQeyFv0WRjzl2tp6cRu
DrNcBhhP2rPDJFo3Sg+G50cX3SwUq0qqJkf/W4R+54o5eKTpLbDV6cw0XgUONj/m9avZ0TLiOBuy
61YQTP8fWCOihaTVai+kDalYr5Qa/7pS1jTU1lxxSI2sIKEvSVCLxBzMiDn3G+CMsAvE2XjWTXiZ
wJ/nAQNEpD3+KenfBWHjGGC6Vk9aYxRx+f8UMhTPqdr+PU5aAquhN8k9s0WXL4Q5bc/68HK/G28s
umShS9uZliTUCsFQ04NsqKksoNw1fClVawA0kvrcTvZFFXOiL9ji5RsJ2I7wi/l3DV7asnzrBjla
Psx+blq0CXAR6uhoAtGZ7748r3mOtvSiukU91RhHQ15f0OkZrafrWick0cy62Xbxcrefz+I57FCg
unfoFoEUF1WEjq67+x963kS5mW7Npr7b/Opnyt/j0yk12/l0PelXrQw9C9XNGPOpJ32wUQJSsNq/
fITbL5cgnGRkPXu7dlqXOGynrhV5n7Ftj9oWtN5qsHE2IxQbhra3IMzfmA0fEFb1hiLbIwJC/FLT
CEsGkoLplddImnYkQVkCRIYULrWoWy7tiPIwDnZNcedk1a1Q5b+cffEKXXQ8WTHSoLCE/zV+7uDB
845L/Cy48z3jaVA6lzuOIcqvyPY9eMcuWHrCLEjLxoGnoQg+yTSYxF1+sC7KxD6EQ/5x7dJ5NMlR
vrklsOmrEbJ0FzY3GL6MXi/2m0dUtIKLYFXaKR2gJ1z3QOjGMH0IU5TiuU/FsbUp3UA1B/P1Au4+
AIU/GVSbQIKrdYSHJDoQuGsqB5tPdZQnc7M85l0gIidAJlYay5hPUywF1IxfAhlKt7/1F2hT97EU
QVL1XEI/c8agELSCOnnhTAa05ScYKgHpUdFX0ee6GsGJ4ytz7lezzpiXqL0uqSZk9ACdoDr1GU9b
3oUD9zdSKDX9o4GzHiNGVsxUgynALvmDAFbu6T7fsxWMgzCzZbqXAFN4cttf1KIa3O1kiKC4I5Ux
pEBZ2TG0YXmcX8F7lWdCdklR9+MHZjAcLk/NBzx9Zl+Xj+EayusHmfuy7e7V6k8Auv4MKSBtB+sk
/f9jiD7FrUniUtHP4HAvYOkyxpjnDVAeKvcO5LX+jwENqVcougPWGovtJE/GAfPYzkM0kGpKIUFe
scVLn/H9iAkcwi7sLPnBUMhHX7P0bMgFRgr4XQ3exRhZny8X7KtTqW0Uk7Aa7svDRn5ljg1aulZz
FvTekGvBQM780oTf2zYzK9U6cgpLqJcZsoOMdwVESy2uu8e7/zxtVOyl2JlGN4nfHkvjUdSkfK3F
IWoAzMiJTMlZovy3GTReuyPAYmBc28Qp2K6g2DTQbW8zVVnWguHsOieWQHKxvQRi0u/AuF0fzMov
fnYJr/oQhXqiGMIzrfMC0Rh5Ch1TgNdLxJdYZpmhlv2gDbaxhEqMdY4fiDT4lbQYGFjvh/XuRs/c
Cyq5dGf8ZkuWwxcsCTFJW+lEoJjmk+XYMH2cx35gF6MlQ2LWc8GJu2zoyTRK/OsiYF5R+q8kqALu
mdPtngrRSppPgWQbWdFwvedg9NZtF6N9+lPmCQiPpX8XoAw5RnipboZXmjkQ7TG+YAIX/Tjf48eA
/SL+L+iUkbBrTxHM5gmnIwtgGFzHn/FVzSzo1n5kTCAtOc58dFQKufdMyiFO53EemhlTYUzHXJEa
42QYJi0VLYKpy7KV2YFJ5v6/eNicmeS7e54IXXFXYvZNoSIjCTTlpy/0GmolJ2uCHtyq2zb5EjJn
8ww5V3NFA6zv9hqQZTqJ2f8xcSrruAB1vp4ClABeGKBvfBZ3MT7NRMDWlyadIli1TwvibTk7GLX7
nYqIRmB8MqAne8LngtC6nZ7AMeqGahP3AYrmsv/9AeJqtNgl9vaGA1whbI4VsIRJo0UNyPc6I5T0
kxvv2HlxRGgXi2Ijfi1vsqUM8wev4GfeXWJwFhU4nvIndSlH28QkMunek0/1hEt02e5cFu/yQLBV
bgNFQq1Qr16FthPhut4m99sL/DcsNRHX0fn7xy6e73PbT/FNkgQMNUJilQWLlW0x1IIqxZb2AjhO
VNFOaFRQLL0Zf2lDB8w+xghXGPzjDH990n4W/od0TV6eu5Pxf5wC5J+rhzndmxpqyXr3N1MU+Kwe
cyS2ITE26VVTWMk8mhsV8Ayyzbt2TnBomeHLuD2h8V9kV/eJQJjZR9f5kJv6sUQNJHVaHAe2l3vj
XDU5u1SBarxbsul6d/Ow8Mmzz7A/2/EBZIBg618Qt5FSRNDQtjY25ITNGiG8+bo4DSUVXfEHDD7J
vfDU1Ws7zzKceTBgwFo3BCTN0vW4lonC7RQNNiJ9oSOXBN5pjQI5fz0N5qQTmIZZxSi7K6C185gF
YmlUtoyxvENm0neziZHCR4rHPP291gN1sX/NaIwxMlI0UOr4DFgiID+7UAtucwNbqJX6T4Qailx3
S5P3TPzCqd6mYzT8piVdBGaD76U+Lxhf1JKuzdjH5vpPUyO9+BsE0EwFDFK4P7VY4nP3lIAlJp4i
6VK0bVtlNgZCBtycOUWX78buNo29IEqznDukI8f78IQI5rbokhdhWzkwUyav8qBW743t0l9ZxWmU
j0SJrqKabj/hU5ubFV1VYkSwS1rztRP6BLdlCxQ0lW+NCMul9BvIPgCRejBP6NtVprXffrby9pJe
HPw9kCjUEEK0ywEEtsZKLgp3rVmysfg9g1VWqFgNQNY27jMl6wzZlyYysKAVu+YohDwRc4OJhdLZ
PG8VHylheS/sDj43lYj5sI7tT2GyIKV68MiK6JM/yUhnNDB0E0bfFXmK6CuXyieU1ZqdRAQGZp78
FOyQBODuawdBcwS4gnnKb46IhoVsbF3HEFPW51RrsaItw904lJCjFObu4z0IFkZC6ApuOoKFpRLV
riGfXIGcFEGxlYyXrOS7AlejRyYlwV+Iu7L3u4p6OUKnFFIVB355ATKjaaKUpj6oZqUoMuZyss4i
uK3yAWN8LLtvY/hmcc5xKqpnO1fdhuFxgXO9NXwWef2pr4wYy5mpe2l8cbpx4Qb6BW3eu9ZadNlQ
gly7t8jCtuK9p5YUEoa0laq2PoR59i+mG3B9VY7mrfPTVUxG6We90XAvNccMv0FOQebUk8B4FE65
dGBWzZ5uH3IZDstQcgFOglijWO+2MTsKZzjYXLNMH3w3BQfmYepb7CxN+HvzeJoaJ9R/HpOESjka
XMNhJMior0+O/wKWz31hb/kiWrMSXaJ8YmfsM8zamYybLwIyAKutNZKjxRB2ZgMuzl+05OZQPaf4
Zul9Ld5MkWMj745gLdbFh9CbyUZqMh+oAykSsFYJsVdfS60aNt5XFwr6oHQz8el0awnmpH6HLwvY
bIyJ1bp6YxLAsT5aBb/S9eqFJSpJjL8naEm4D1zjUqJkNr5bYGK8OxtZyPmFjfBvnY8JyrbSMvcY
4y8tCXyGv+7+WN868Kh22iagF1c9kWa1+CqxfOlzS6HVdxZqPE9H/zwZdYYjpwKpz+0Yx1PzO5ON
eD0pK4amDNgGwdN92WA63C0pZU3GLs9gZK6b+zFT8BeSQsUShNvuRDj7lfcg33pVUjaqiabnrqEl
7EL1jAMPYexraJPx+kW61Hp+e72+0MmNpJxQRrDhQag35MIOb1mxqIj8PDcb+ohGe+fbpLkxXLpH
hacKnGia7Ge9YWcgBEjbGt/4wDBjZKDSRPse7+OwrRRow89swrfecwvjALujU7qvcvAessMrmz82
v0WObYtwgGK4+btKRCbICtwNJFTFuUQdZ69cMa8GNnSmS7ZOvblhOJG04sbplGodJwNJkkdVQhR+
p9oJ3x3v7C1/G9P3yLtKHbpvslEMQss8ChcAhTMUQy4RInABhXnGyQ4YBBYFYM6omn54lcE5+RVt
YcVewlGAEzw6vlUFFUYSDSCkFCFm4T0ZKw6G+V70eDJgO0NQmkvJ9728GtNHYayHFHXyUmEEet0L
mKc7rrj4fp5YVT/fgkIJjVRo9Kdd2QaiJ8DfZeeUSKn+7u2invHehDuo5dSPB6ly5jMiAFuADW01
nyTOKnX3ipnm6c9w7VOUaOz20K6HLXSjCJcIYE/AosldosELx3dW88CwIdl4wzWa6XR/Ft9ZaIZQ
jfkdsvf2qQWjUhF1hrKe3jLwAx+yFUZoZVa4yiS2QGa5GCPvIm1KsIv819h3sDd/5KPkaOKjGxzN
iV/MCFVJUIT1G2lL8kayvMCYfyQLr6eViUziMqMp0rdaQzESopWq3iw5KztyimjweQkjqAlIyv5d
qcPXctwOIGo4xw4W6vUNaYsI3gY6hXumaKYqI/dnMo9FxpzPmE2CdSYKQYeqT/l3tI0+i8wp9qKe
Y7gmWsr+ggHUuZKhf5Q9tIAtDtAdUb8vRQkt69NepuxBJOUCmKzSurbtXri6HBn3pE2F2wMja7ay
qdXPaesUioZpnVa9yhK/KVTTg/Kv8DielAutXvzIPuWu0nUuWajT7sYHx3jTMRhey6zJotJ8D1Dn
4To6zHoMuXACy/0NiKOH5fmLbMWDvbtrOMzsiwFg2yGJ7aQ4+cxwI6jx84YHizXlsdu4Dx/CM7pG
np1Rgb+Gd9A0CZRGjIuabLwJd9ZNzh6VYoHfktrkw0RQiE3jQG/jD4XdcqGuAAXtErs/YWwyudCK
KKid6vyrVbwf/BQA0E3YgRWH/QGbv0s09e5eAUqVO1BFSnZWajkRxh5ENBaXLDsn6ftdRCW/SN+3
6KV4AdPud9PKO8JBicra1MEH0gRARi0EAYg4Bfykf+BZ0hFE/wXUBX1fJfngjZ/8bUnSLBeVm4GL
eDAzwtZrUmHHg6pYVBtgZ5ATpu77Oqit8xPnZJR0voEd24Zl/tDMmi1c62gwU8M5y4YmpZ6T7zto
3/QaIH+CD+l6gggAE3fl9u5orWM7/mRfVtskW6bWM31jCNSBk4OjR/bZu4yKCUSJkwgBx3cAc1Lm
CQUAh9V9qFr0DtH9cKAZdzaBTB6LnRBsJej6NjVXPCnplEhRKAWDSRnyV+9rQ/CANWwGCcfGd7dD
iDUSnxoEzzwE+LPBw2RuEvX13SN0cSA0/M4Y/fcfJDEBERnjONN/46206CWetTg39jYUvh3RO+x+
wzz3Sr1BubRlToIme644VVGWo6SSuxrkwwnsyfECdoOUBZLByk1maH6O1c7TuX1tFoqukHq+R2o3
rWXsQJNvGIURZQrWe0Y+RhAE70LNH/nIC4rmkX9pcKtWEzYgm2Z9lmj8IZM6X7VxK5+K8QRdfOEC
YVDTaCSUhx8lR6+2H/YOvPLJBKjLvfInW9S181aHTgf/Wz4BTlLJWreMoHkWtGCwNEoIMSx7gLNf
A0s3UKos6NOQEit8cdLXHR3oy/RYRtDD8EacpdK0dK5emWjpnvpPR8TeG9XL1cBzpMkPVHAPUHDD
R+Fo7G9hKV+rAWEzhcBxBp7+7b8cTK38Q8qwBNVnT0Ac73EFXgYi0t0YWJ5NKchse1R+g4EKFztY
b4ZEmq+kN85DUbgD8fV5nBKP1ltnvwFOMwT0UlOg3vsgv4VrHHiZJRyrdRzoj6Bm8JntqTIQWWpW
LiJrOKOG2y44/IbEI1dnau8gd9UXpofDzDdrinYilMTZ9ExfwnM3ezn0yJGL93kFRk3G1mgKj9VW
oyJ5S5r2tLJKs/k43licO8DgV6NuVP3ujzYP6CTYap2+L13DNeNZ01/0lpAg1D7ny2YchwwKEr9N
t/F1+ZHRQspbqvYynRdz8+pPpK4YI0/xc/4bNiz5XImB/CSUM5PABjjN4s2sP4PIW58NtNnBrIbR
DDKC9ZgsxSCAWnNFOskA4w2U+84eZOXOFM9vTra+3TmLD2kOoq5WHCV+meDQrrpkywoeZipV3s+s
EQtZzwGHCb3EUuhHaGirl6SOKKckcttslNozmhdMJoNF7aRPpVZvO6giAq173mN2Wl0FXWThMZPl
qgj1gigD/umoNBo8y2zlSEV7aHXOfYL+vfiW/9i+V0UFmlUYDtRQHg8q5GVeID7T93MKLUZC8iSF
LAYhgTJjz5FgLN3kuQb9Rjf3vw274kTu9PgSGfR6nA8+NSDIo/Yy5TP3H4KVKqE+5ZEuw49UnUGt
jbC6lZBMsvrpcVBIzBelQc8MsEqc+m3G5aEvBdqh8YvBgL0xnQywPzTNHlsL7NcYB7LD/6BKwW88
rO1+i7R/aWSsE92/rwhd+XWbhul9O9ZQEntjQULxOl+5nHBzGcaJkqzDLXiVm0cj+IgSHqJw7Iyx
rYKXkp+szrps/pxz3qRcE+sRrUzwUGLVK1EN5v9c8UGVcESzJidyybmJw6DhooJhQcm7gwpl27JI
naM2U7aAPEagx5su7doVGMgarz6FAb+q8s4AiS9X4QqNiQSCay85bLaHuzHHX155tibaIsDVllmj
UcpjmcvfjIpULr8Ei4OGqKsLPeNSaz46cI+2teHcBRbQDNrjK4e7u516JPStwmFqQHVQ/fdiEiY4
F3P9YHpd/IslJuJV1e1EoIAuIXYhNl9xpoaNF0bymHEt2QZ8CRZNGbgw8jCGYR/0o6GuYKrMXeNm
VIeHVSMoSL3fj8tj2LVQ0z1BeKtQaluQfddI0wa6pfaDfTCzjZIhJImLpLQihechWclcrO9UngmA
XQujNwUfslwuYAiEp4T2Qskgf+Q/vHjOxqjz7AM9JNVSgHEl2K4WGSAR9h77szlBeHT+MWCEoKdR
3AO5VM+WSsAtzxEyoG8E6NRgys7CH87xc80mKyLk7pvEaedC2GVfW3plP0FqD9/YgbIYEAWL4Pgf
4rbw9LmxxMB1znygBNlGuiH2xaG9eDXYgzXYpZMcGVy8jB3YSSERx2lJp2Kaa8U7voigfEWtDAyV
GaiCXCtePU9jqSr9Vz+CYedFBZGDlF+5Z1VMne12iYBmf0Q8t6p3hC+AV1w5TXy+wP4NmM3Agumq
wRpdiCLCxe+Cr4LvhRZEvSj8XjL14bGEB3n4zR1DUbOTxxZra18tByTwsahVy3oarBo/chzi3Qk2
WTJJkU4sPGq5HkUv93oV7eP+nZvEzVt0uRRLhfUSZgyFU+aopqHrvZY1hykVMLoquXkMa+6Hxo30
vgG5tFkCDoUABGNP27+X1CsFyHLIyit9mVhGZgi/WKVx4w51TfQ6mjVN5EWkVK3paKzbHzQlii9f
5F+ir6ItMIU9X1kNI5YvLumAXL8jqvfc4m4vgOzTJqtuHi2mDbIDt48DgU93/aak4GhERdWyYsnh
55C3fobgeEW6TanjmdGJVNbN9vwBDfft1CP06z4wvGpLHWrVSQXZ3ZOgmJiqBZWTGIJ8x1I0XmQo
ELaFJadEm8YNYc/3ZDZIBZUH2aUIaNcezySRz7oTHdUKlNPVP0mhMfdzY+gN4C1VIC6qEwDWXZSv
my5dENMNrK2Jv87N9vRGpV2z4vcbMhIag205CsO2dBuZ5cTwMuW46MUT9LYK2CVxtJW73l5G9pZW
ip20vabpeGcdL22mhM8KCbV4sCyXFeLKPk7oSmlIVWJKjLIJNwE8LnyV3dvDIrm1wqi9RaVgDBmf
J1Qlv9UqxaqDjtNoEeXf26DfUaecfWpr8lYskX9qL8sY6KgijYPSzZ6GsNVwdY9/hBhePDfr2uwr
oY3vqXBpUtKpG66d8xTxJli5/xxxq8fUAj0g5i1bQaeg+TQdyM1VaBc48TY4T3MOb3HWMGZ29qFV
o9gtsZmtxcAD4UEdSeodp5RWAf5qwKtIiGjqil0qrtkAvthf1u09VVRJ2DVgQgpXOhJWF6ZeZQcl
s8IelBLk3lks5gN7mmWjl1L87dPOtCtEvvPh6/yKDVyP+IarBMgrACSWaSuh3cYGV5aNy2cPTQ3j
CNiNatU5H8SeqK0pll1eUbK7MT4cysJN8FUuUpWrDvYYqaSSRu08821hQoluk6mJ+o3nxRE9mu4o
MyQJU8iw6sut4r+mA4OoWDAfzvLhtEkh4Gbq7QyJlW/sJ7lYy3PVCH6JVPlgMXz2o/B+Wyaml1SM
GX++vSuUd3pfdXXoun8cCOSPPW6IarcdYT6VsIzKKeMYXKT46VGWoj4i0OEeTgeMqwF3YPK/TJig
DycrQbI4oYnFH2JIFPc4Bf/OkMkWdUqGan+Z6VLj1HMt+hDh7+7rBS7ZT9GmIazI4BKRnQEr7Iqy
LbM+/mPkrNeAsCaXx6LeCkVpOgdqCBS5pZTqket9B7JoTivkMJ8XSoFBPg9j+AEak5jySKUxzmB2
D9HkSiqb6ClBcPUa9gPRsNFXVySmSmoF2vandRxE5/1cGgoeLkl94lIc+6trM2IUd30sjIpEF6cW
lSkCXtpwpTVH2lRtybhSVUe0wc1oY31jgnZsfQAwGNc7oELFMdo6Dqdev3en/z6dQ43fNY852d9a
zZ9DcB5yVt4A6bPrrYRiFCUOp0Enw9DPN8SAOBCuas4uUMQFZAsQ0pAUlmpb82MBPLDNxyUENey5
P2vyEaFbfd/XiZzxVtuvkVauOAWl0cesYZh3GYo52RIDuOMkwo4dfhjV/umyqcutjTIuhLiVXkZP
NZ+Zk/5KdePJwUl94d2Dl1dLgBYzGZ1hAYDaVB9YYNgg1WGeU8NWd/ZrBcQmTj/ybGprRmVnK6dc
jHCP3a2QNn0gnB1/0XasWXl4I3tqb5bpjvsomQBOTi2EApH5v8daefoO4uOScewgr/UAQowKTP06
nfJYulPFt2YBP7qAB6aZ2xghbICkFE0a3eX2togr2BjkzXJseH+kYNQTVdJMaurANYdBIL9fkVdU
Zwm8d3xaIG3PBX4W77VW8rJOr3nBXeGp87Ak9NXbQMeSpRzzm2LRBJJ/IyYHI0aVNVTp9RjkX4dZ
0H+LTMth/x8BpwluqtJrS3I8bpxq4bQtgxE7VXm2nsqaLlVAODqICCgcLg40mxDsmqIkrBsoVSQu
gf84hb9/XYBDxNEEPvyHprdYiKRmaZe1BxeF1F6EVG5Fb4gWYMrwMT0DBGYtC2EdS6uIOhllPhqG
Rx2JEZ4+1LCvQDWqLjFBvMsU3ayeoMVg7jSJM37itfHvXZa8HpG/Vsu2kBc7Wrnx69F+/2x0j036
VRI+B8ahzvYP6i7FV33bWWccFWJcTL4eNGQPZuhYzJjYOFAfIW9NkNWWVQKt/nU/Pp6JoSp2hq02
ITkOBEogryxUdlqgNw2uWyQK6wUhLOHoqtA8Ygs4+cF5hDkPKRWlcDetw/OntCUc1AOVdN1DaVXL
xEs+FHD9OMnxGEmi+ZG6hPsrkbzYCCeI8vsKCL6xcSO1AYat4dX7+9DRPjm/8Si6i/jG1TY/fiLj
vv2mEQpe9rHnLNQ6hx5T/BHkJ+zbdHZTvZqfHT9JuZQvYZN44ls0NxmxcJQk+PMB0V98xNzwQhvz
GQoDRApT22vYgCwQBSyhVMHIXFp+jkpC2Ota5uRX/cf94GdlC5Giq92IbltBG7X3FE+WfstuhC6V
+y0XVpj4DmvMdq0IUiLCVHBTmfy9vGcRnLkgBL0qhScbvnQ7BhRGjJTDcMxFnmfCQHPIUBXQU24C
d711bXgbREzgmmoOtyw2KF0SNreKk5BUnbv195jxe8dNXfPq8j8vXXlVk1Xdu2UT5CTaxrcZhnaL
4V1zmK6+eYo/Xpe2lodpqxYRcVa7WK5brRgA94O8hgaDXwKD8AzuTynONHYnewjLJ4NFuiyByg9N
RYwo1vWhoFO5Nh1avlhaOKae6Fr3qQuWOsVA+cpDJ7Xbj0npamf71mfSTu+Vr1riPHjLK6jkVfkV
SOYa8V5z9Ml1t7QB87g/TwpmbIP76xQUIBtz7WTorzg5L5cDDj3uZYsGF8RneCs6bymbNnyBhf4F
fa4gS2VeRqqN3bonkASyWwxZ6pJ4jp36x2/Nsj66jMzKQq287NH8NTB7ZTT/s8/lvizyU0wzKHKY
NyU1A46HIp9fybDBi7AZYtTavg/DJhqOnf6rQpa49JGkZIEFZqRkUutnnyrCoymSV2X2ilBvqZcp
oQ7mnLP5WE4ENlxRVXryyo5TUbnbarICcaQZltpMlNQvLzyPyEk3cQEP5o2rf9W6dVpndTOjun+L
VODdBwRcfXlm5mUfBtP5glGbVY47acU1FQdwsecZWaGOm+OZHPiiqwG9iLNpnx/z+4eTJX1oAUVZ
XU7LQR1l/cUe5d06xYGfEb4EhQfit61DB96Bm1RYosQYWHadsOCdaiZ/E87oLZTEidr46QxvDnMg
Kfr1mLEkkNIGNqIqzyyYfIBOE+xATaWFkIUg34HzMvRae8DTUaOsuQnjXxuKG9zLGf29cgfyLRx0
aPfOJFtocGB/MlQgRE3JZGakCONCUdNFGw91lET56LZG5qQMlJQ+HJwE7mRfD4yNcGJRT56koWoq
J3RfINaB8V2pjuwIhXanqpWV1VkD6yEYem4ebtA2HzKcVy8BMAd2QkBsRzynPuRvDA5Y0HtKOajj
/8/NlM5HvC+RfMRLFgN/jjjyMNdMPepXA89asa2SJ5CK8PRpLff6MeKUQLV9UjSTx4ww/7/jgpsF
6YqtkJgVT5xLfU20n1JawhBrq97nvbokqVXIH/r6Y70eMs2PGerlyI4nc1iFXF3u96tSDvESEUoM
94jC68tVrX0Vdb+0kgih5MFIUeWM++pISHUB8lx5TQoSB4Wn2OVb5sKIYLaB1EfXm/L+bXlvSNg1
bRcBRgEyQCunZzEoaspielcsnX92sKLVNdkPb9E2p2sgNox01JzTTHXqJkJrxSrkxxa5HvwRhnBf
FMvWwRRU0biqOxFHrGXaoyxrpVogB7uY3P6p5h/h+nTYpLJ44WRGrMrnCxLYnTBpDPkkza/KgFV8
eh4PYlCdGnVpJGh6XxdT/pFVCwKkjSNDaegq5bje8XoxoVaQuBnRqwOQ4z/SbO2Z2pyxx13quegt
h6R5UM4jXiUvYd7XLiWEpXBSUhazj4r5i8eW1XEmDxJh29fxg4TJfS1shTyPtXB/1mqSDf9kjdqe
l/LVsAdB75mGKv+WLO01v99INNXFV36/c4CtDstaoazC2kxlhQLErjT3h+3IgfUBqdfJYzF8+QzH
itAT45IF9amKPfCzVQBaitxwdqUELZRwgQNYiC/u4t2PaxX32mO5L7iKMeKk4RbUGe5ihE/00DRl
WngPnAFgZABSYrUiDYlZL1c6hoA0C4RsbLBohAPw2dKzx1vyWXZnpuANoImeetyaEwpDpfPK3Hfl
Tawja+q2JfhMjKzVH9gMFiFoAw7v3qIq0THESjZ67P30IjOMDAnIpxPm+NdFHOc0mKW5HMstbmGv
upuU+o1AdMgDu8/eoBbKdYnmfZW7B0VUBGxmu0ZClwJVgJpJvS+TAx8yF7zXPW9Nsd/Y0E9dGqi5
W6XN8PoARYdE69d3aqnMKQNEsWAk5zY+tTXzQTPgk/pFz2xdu824I7yWDwlAHpSLDthsiB8WVKlt
13A+2NQqcTcXJP84UI09lHooYEgrPeXphIynZpyGwXo0Yw+ieRO2uJ/xB6jx8DKcdwRhBJFN7PcD
xGXeOPRG8+9geKkF7Kb34+C9M6nUb0x5YCh3tGXxrIGcVyM7dJFe/ZFUOmy+qaWbf0C/KBoivF0O
p8w4L36s4CnCth5fMy/ZJEkz5QfrKOGOw2lT6uAMgqse53Ii0/s63VSSE9tZS4z9dSIJQiMdrm6U
hAX1EgxI4pEeEIz4Ci//Ixyrz8fvV/f5uNITECxyP3MKg+t35l+QkXBx0ExuB/wCtJU1C07rveuQ
WZomz7WVEd9PrUl9UYY2T2Y0E5jCcag1nZnCdYb0CyTlQaRXhxraUqU4sTqyRQunmu/tKSM/8g0l
fyS296rYw22fypmJe1YLoYxHvMQwoXiiPlXO9dxwoR+sB00j6Jq+cB7X0W0uquiffDFAldfKhpFG
HQELSOXxLj+hS/3mCXHCxYY/mloGKlDmPlnEN/81OczO3cxHJwynYJfGXPw18qwXPghOqAWbUqDv
2zZfPkOXb1NsyCuskJ8mvzAGVl4aUn9m0gD0LJmDYbL4xVT6uVkkQB4Bz1rk9fXtZXfCqO29SSsE
PP2p8bwk8pzYjppC49Qc8aAZ7+zqWCGSX8BReawLnxSnT8gEfR1K8iU5W1iBSNCQ7IwQu1suMx+F
SGW2cHP4xF5e1LLH5SXBhGDp9uZ57uzkRZMWH74qUoWLPZ7mZnFN+TXO1KOANDeQz0y6tXI5r/2Y
yDq32oKDvQdkqrVZK+GI6eZgiDoQ+/By1zX1N5TfwZVo2GQDnRVJoP6ROrPoAZkdHAjDVW4o1tPv
Irg0sS3iIbDgJTYideTsei84DsFJK50aGXj7q4NxToYaofCsxWTPxGvuI4MIH2rzRO4Q5zei4Wcl
+tEAxs3ablopnILPGPqmIIC/P0ovS4ywjvvuobreQELNyk4SNk2r6F7zGjpA6uRpXARn98Ay4oyw
SKSrP1p5WazRNS2bIUIQbVLbCDEeFzpXaGSdNcu+tPq8nUmkoq+XWfbLlx8mJOY/goFZn+Si9BBy
cpvKS0rhLiFwx+sM1/QEPrPdPYHneYS0BJFna7wI0+JVrG/UNQcEbYQJcyBHFb6y+y1CrxCQt+27
rzg1h/SrlC5nQAVnHTtqzSXLo+p3WGtM5VQ/kczrUjoV2RHn20yNJTaSHsCC5RisKRzyP8tLC9Wv
7uNjhFDCUnZp7CRq0Re8qG/rwa52js7xVCiTvSUqLuKxaza6oIyn725Nrv2F1Tyx0M5JNNZ8bWgN
qRwNcvnvmafMUTRt98/dB6NU08y0CsOpGnA2AdwnTjQdunxPa0b1ApmQVc61lqvwYIKQsPMN9cwK
PhdJ5meobUfPk3+cQKWDCvZivThvTpNQ9l3uexR7o3+99PdI/VSgTIHSqeJ58AdO8kJ3gvLP6Wc0
yD+XEPKk5KwkRCQ42o9jErtotKY+qmam2PWiYJVfR1M/huiwQEwKrG1W9qCeNWF1CoEMMFeniQs4
mbS0/yOKpzad4uT0B3yMW+mOHrJrNaiBzFLARSw6/5fFDCNnfjYi97RfBcGc4y82SyLcYhL5lkeE
qmDNVFLoBUj1GCpHE/Qm1BuSvE1vvDNMggKud6URX7pEnpwUZvxoP16H5SFxA6INoZY/0TaEvKjR
h+QqKRUFB/1wSL9QknQiIWEJKLRJt0wUXjvwMmMuWT99spJqh/X/aR7f+7Q8aHGNg77GM1Jdfvam
3e+iawpR7mPPdzBFewzlAR+Yw7Ii/iOUz0OCJ6dYLXtGF5i5/u/07Qy9oWZAYFnm3NBBmTB7SILQ
eeiisU+36PpIsvX6WwQpyNe+HpN3Y/0RIeKg5Gj//yf084a9Grdc9r81btze4USM8lw4fl1IzqeY
4ZX3MryHiaoK5NyMVTipUx8e2t3BtsdGxH3W9xxEhIHUTcQ/+ztIeMvCwv6ZeZSmcc6Dm0NiwiZd
V6CyY3MfWLVodKCht/fAHk5PUICMqj/qtuTd1M0/qcTh42UdmpbH8v4IJeAolSZ8p2OfWQAoM+ng
p/GSSw3CUjFKAPoyB3QuhdJbrN7HM6x604NEw6XbTGJu9bpJ5LoL/7xD+Y/IoM3JdLMb0e7fVFXu
MVtvbzeR5L0XNWMlQqOPVXWRaO5+nPKyCtc+PdqZ5mDFwL7nXDXsQJ6N2fdESDLH40zHYfEwtLul
QePAmAnpAJRe5vmew2Dim8jB2sBpQRyNNlWgzfFzzhZe9Z2hLtJ32xtedJgf2kEDyQmhZJPo+hyO
5Mz/70eyNNuik8k1oTp4XcSBBZ/IBRQcXHyiQ4j4ZSKPTN4nwzUahLo9fYW3Ds87H/RJcco4bOSg
hNhpafZeAL/XByk6ZYgeTRXlsLhUs4z3lDXKwKhkQQOym/rdD9zgYCf8TOutjAvIja7iF8ZuNjEd
1ObX7pbhCkYBK0iBABB0WqFYdIK3oqkLDOTJd47krgYwyt2m3AQ+ph6j8PFZmrBwoFi53H9l2CYj
LmikqFBNEXrHk+7BGRmALI1eaiqAN/v4ok/uzD3UcSP/UrHghJF4XB6Uzq0e2YV9m0Pz+GO+f0y8
Lm0GmTXouuh1gYqpISZedWyXmBNwvk2tSIHqetwYtAnUC8tcm/g5jp41Dgx++yrQZFhUyw/sGRWN
YxQsyScYNNz1jUyEjjkWrFc1TL6h4YlUuAr+3VCTb19i9WyEAXJiP9L+HsDsxXJg4z0hLkqzlgDx
AsibRUtnFgq0WlZLFfbZmsof6S0WegLKe93UOwjKJYgS4JD+Oq+NiiRzYeSuWi7OvgJglriN5h0r
bF3NvnGSQQSdOTBcgTJai7lVS53Vji6T9sD733edUvpzzbAIlbNP0OvdGSLJc6EscoY5QxrN3FiZ
++cEzT6WT4aXqu/gWvAeREA4l6+arxB1TdYykOp9huf6Udq/xa8fH7yaBca4q76jxH2ZMFLgcneZ
GAaCaq7hCOm8DpFSaOAnIGIoTFsYVckbyTlpoJn0/Ncn5dnFxfHFG3Si6XPfucAgfA5loOLFjQ/0
LC+BMXfU39bFtSSupNmT1R+MOBKB7/bAjf6P7eYYjf5K7xJbEKVMXWi+6nJy3X8N/y30Ci5JnpPZ
Rff/4f7CTi42huWUs6UZ8oobSUw/VXpU0rpzHgAWlUghzaEbknxhvGiKExq6Jq5ghtX8JeuzD2Nb
/QzSy3oZrIJXrGtU1jLe7madYlerxQmIdyI07YX+qNwWZ32CLEEPAhsOf8en9NgsljfBcOiM27yx
rk32mC9RtVRRQAxq0M4YrPNQIKc/hxDHQWYUGrt40cGVsoWfjrKvZ3LGopvFyE2Dc58rXpJNFOgy
yAlq1knBus/4jHqjI3wGmqvUC5TW5P02vLc9mLBDMw+256e4L7TtXesZ37EENiH9l3yUQZV0SfvU
3s2VGoiScCHZl1WhD3exRHkPMYPUkEZMaU8Z2hXwbEBZqlFTCX7B/hjbQD7rXuonKbDu65qb0YwI
v1ykdO8hR8bordu1r2oyxRaEj4oiQvNZkHPczZm6ujH5wEpTDDDwXYQHZMTR61sf2zxZ3rLAV1YC
8+PZMEKF+dgk1wKVc2OXlFC3llqzK072osjmn1DnFl7ylyc6BDpCFcXtDSS5VBJ/4aHDuUL841yl
caw23tGLeSbRfmM9fh793bugwsgTgx+0XSsWLiV7HD/pys04a943hgLC+PjAVeSeUWa5fAzDFTom
kW8w2gDbQkmR33NSUXxnqViuM3mKFx6HHbdI3ocTcfSMDYsqJRMhq1oAduWJ2VcpxbfMQwXtoaBG
ml2lnBYKLawhiEYgdIjMkT7mwL3nRJ8kPAGHO+g6KqCuxMc/LPXc6T/aN+EZTV486+Xidmh+trm2
soQQpgLy1enOSnqmNJVFyzEotQE3YI1CsI+XSPF4z07SzryTWTbbzk1MWrdDwN24dlD4x4cdb3az
BRUhxVsyVVwP4iuQVfNwPaMhEDpOAm5oeGBi2s3sM34kZXgeL76uDKPZ5uChxye/O2ZUUGLb5khZ
VC41hdnmIkm85bmO0f3DnvUpwcSOYcRxRfpf1FlZYyOesTvxMk6bP6YdUVEmZEBtm+fkSmn+gR/f
TZe51riuiTH8IJMzsdyW7lwoKgGFRS1CRbGKCsrRFWTth9zDvZmiN+bunGWKK2mOqJhwFJ79QLlt
Bl/41UNMgtnl0Tlw6owwn1hzUakDzm3I4kQxcNGDMY1YgOuBsYsbJCaH0baWnEO3o5MpmWxsQ/YJ
mAh584lnTjkZijYqMsWfEdgrlBeumdNQqzBh9WdEn02vcC3BiE0xgzvdOie/Q4FknSObEK4J47RC
Y/UaF1SHR8jmOf94eRb5kAeM3FkdZgLsqeKllduK5Q/Blv46JsPGVAGjr3iPpsGzDokYRHexUeGb
1UwIjz9AyI//CuWrrC6/1NTcQZjgjMBN7Kab4g5WNwNsigPa/QZjwevx6rE7wBFKXSNIx0jLpemP
y7dwViV+CEztFrVbwGkzHTme68qsDSqTopNkDA8Nj0DXJZYiJX+jHQ/CkHweiuDTW/rWVjW2QEmw
gbIyUfa4X9S+9GHEUdY8npU0eRdCZm+ioKTZ0YrG62qpauHJraWloN8bDzyCYUyesjIhzblTOe3z
LKEYOpfdVHheHlrKFWmARijXMEogS1vYyVOBiDPKHqA0vFdtcw6oteeZAb4iFIMXgM8wy7lk2Cov
ADGjny1ib/0PG30ZSBHi3d72Lj+8XHBRZFOAGx2pGMFU+7+aI1eTUx0mP1xxXwy1GSuNLPHkxZHR
cQbai4uzyJmiKhqejTQj0cTVRxlUV4KRiBdsqIlAT3VuxTjagrfctvrOq+/YR87HJOubt20OzWzD
Dcqh/2lMpyfBaJiQP6aj+umtMmHnv/OHNABucpwYzlzsrA333S0oUcU4e3aH4RM0VbNB7orOeODY
IVV4eXPPzDEQ0Z64v0FAezNHR2P8itxvsIisktT8MPRU6pgH0rahjHbnaxa+2V2YImksheIAaiCY
0GBFm1jvpt/RWlnZb3/GHsWV53Wih+evo36GyJQlMeKYGKTF5SvUT/hj0E4GwMNijSn1YQvegPtK
YRazwO4n2grT4BfK/x0xtl6e7MKML8ZT3Xa/gZPNK+tz2hM7BhBN5+zB8FCdgI+fhyKVjz2uEW5J
y7FOYwLierkG2dWn14twNoq+nELFPHy57+DEQQJLeYjRkz0KGmg+HilEpKSdfnYsz88RsNv2ynPh
o5vLUyxpH/YsEUue+kftSC0KmHrVc/lt96pheAyWU1RVQOBTKyTQf0lmDm9xbPcld0NzqZcmY7BH
bd/o+lTmqca+yVL8gkXj7FPpoM3As+CmIK1ZpQsn43zCMQlVuGApKNLpjvbQJqiXYKRSwKUBWI73
Rgpv6kE5zCDxpeTplJmyUtVguUOiZaPKTD80NP0j+E8KvMhqexwNr2BkjYnkPpwevmN4W2Iy3r9X
sPMb6EybrTTn+BkdPNf21ZtwrwTRRiXtX7IX1BCPDia5NenEytimBK0EJxFm5WBXeI6dZAG9rfsa
KTSUzXlvEF9Hc9re/tSphEV13GZxfItTZjCbPYTQUjeCnOir5sG0gH/4I496QTuwg+SRxaXAMtKe
xeYYW0FvsQEmE6qX4fhkVxHM+R+2Tl5lFv0LH8bCNh4W/IdeVCMD+UwdRMsymwP97JAfOErpt3Mc
QL5dIC0eGLtCNp5CU4A/EyF1LalWVDfqT419vynTRl/lu5hnCCOYR7Dd9y8HtoA6w6xANfRNtStu
3/aYOrOJqGD9P1l63qZSEe0cVNwDCTJLssez5sBiR3978Dk0eIraZcz6u24KC4bYX6+cewfTbqqY
KoMw3STki9yqDFZ4rcrUV+9DH7nsu/vRG1/35C6YTaRrc9vPtssU2djCT9ALHgKm8QqyMzuBNjUw
J6Iu7vAHG41REmR4PNUDLKGWe8OgbEgeEMPyVDNANpvidzQ+OrktMKC3EDnlAKlbOiK91B3E9gcp
wK1LdtP6ntMDXQkyeBva+VQ1HyEaKwXI7Na8MRGfq2JW1u7XKI7XoDshi852gjRHKF9wbRADcTUf
mvfg0CpmgDKs+k7m9kxTaHoZVHikYzrNYMH0hbprw6aXI0W3CEVVVaW/oH7SdFhIVoIyVFX5Dgfh
8EkA1tkqNkDBopYqLQKRqw==
`protect end_protected

