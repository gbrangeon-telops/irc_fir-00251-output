

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Cqo+FjfIOIw/0Kghh877RN5JtWmUPj/KfIaTRt94dXWp8zshF20HfBCWrK0/KjFcQ6xaC5bYfJZ4
kTgDE7VoLA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P76DAxdsqqBm7Dhm+Xv4UBWtxeM3n7VV0uwUkGrQnJyruFJEvMXWtTIk68wS1svCurmxJblglPTM
AUuHl8lZTHelg/xsbfqIjFFpkYurRbfQPaEBBncWEUkGXitk2MsCEJd1XKoy7X9zf5gkivM+Dtc/
HmQtcrnx7yMmBEFf0wU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TS87/wLvg3wp8BEZbJFwjKct5crsKQKmGgle2kFCdS51Fi9lA3booRtYf7PKimLYtiDNKzFnNmDB
yS/M5Wwp3OXdwvzTqi7m8nPDGJzv9CPlgJYl97xwwfb/xlITgLx+mE3FLNjQYh1k2fW/YeWIYcJ6
dHaLGRiPpSzATplaiEnfWr4z9y5Zgw529sAAgbJqopXb1oauD9xMSn+2U51TKQlk6QzJOyaBGs0Z
cYN8i3mMrSJtz9+1CorRnx9v0S2lY1WHtTTmGGV3GXP4WDMI7lTnhoLYTdqSlyv31x9qhFidZzgn
WXAPS6oNxDavoZXEycPxfYnQwSx2gi0tzG/NZw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NpAOviX6Xvaq+L0foSrleTOrW/NGnS56aJ5rqqn2Dmt6YUNEPYGn9LoXqfbnr2nu7OxEo+FueCzR
GTO3m2J9405e67h9qARcSi/hF0VUlC6bqx3PVbV+Lg35W+tGaz80NE2OUHws+A7UXDQk1Cp7m/EC
XxMS909JUlXKjJHNQPk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P7klUwNMTreRZK7TaA1WE7CMMEOTtEjomJfZ7pHl1XNp0UR69ZqgBrqFP7D39H55daou+YH1hnHn
RPI1HarNWCxtLMV4hOqf8NjoCFBgrnnB0U1fZ2Lr4Pjyi28WQhnjcgxXDHuFaQlXuyVOq9XUsvMJ
ssrZQdiUjtMyy3njm+Pnbmk63891Ob2bUkQGGCsGTzQYYho8qCUxVS8K3X2BjFQusmuscPspGR3O
NvboEcmhCLzlJh3n01BooLiI/MFAc4YbNKfLIovvQV4EihZ5noxjjP5wWP91DT3v8RKOECGo+vl0
XfgG1PKzgtiiXSw82pyP+WwelLF2xj1qh8+H/w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13728)
`protect data_block
M00yemv74riSztBDYXiMCZQ7l+BGb8BjVPIsHclBDbJiPGYxW8lXTCRh3mR4tksLo+gX+4MNT/KQ
PjMItErmGnBfi91HJ1xuBTqwTm1936P7Q2isfirqmK9LxK8/sy4KUgmTBQqklsn+rN0uhOm/KoDD
JMMII492mtuSB00EFXNOE0++RFqasHlR/b8l19l63gwsnPeyGgJcrOiCg+b68v8XsvFA5qyQ4uhZ
On1XJ5L594tE1VzOufMQmv3E3l78oQ/ed/uWoteMBBfsfJAPRTC20GnPstYREu5qAK0yjqtjxAuD
mIWyKoqgBGSN71/MDBafHbzEtpyYIDPVzJWevRfUGd2r0HSgPm7/OcP0AjzVRYugBhAGFOsYuLgd
6aKCblIMfr6nW4lvZt7NdOJVOLBvE+TlaIlg0L1vaYOGlIbda6QX+FsBx4tsS+6OC5eU0xe2szYc
Yj1whMdQwdkaXPx5SoCVpEGUy9V/LxQuXD1doSlpJ5SEVVoCsGm3NcYudYOGXQ9ptJcInREm8/uI
dfhkiXcN1XHjlwM1aRrbuzlK8RIdfWp8Xc32vuXz0eWsf2th9bNUGGaHZHBCOS00TAaPkjYOoYit
gJezjiidtzRYFFJgqrrFmuA2UdSgkono5DBYrUhmS8SyVT9hSEGVYshniPBr2jD8k7B5vLglaKhu
LNekny9IL5+PkZlWq8q5/2kkRhBSFndX96cmIK+XPFagYivnqZg3oRlOForFUDaoLL/I6XLtshBv
0ugF9E8jaqMB9jSaxrs9c0tqbJGTJ/k4Z3C0XQxRlxDU4HUFqlVqCwbMDxSmgNwy+yXzJDDXkLs5
ekqEH9WMk1ffnqSx22ddp8qN+iscfgDtnjdsabS8k8di9KPPAuzMCHa80rm5wDb6malqWWwEW+pE
usktdXdPIftJqH8kVH21P8rxYKLCTlQSHVzRQKdOfA+9yGO7br/w6v3MXSwmX+5JTA3wfTOYMevv
BN1OJn2l9Cn0icMgvEzNkfH6KuPqtSUeI0fZ7diEsmDQCftHZquYZLKZO3xJRRMpk9gNJpO79/rr
jg1ne/0DhFsO+o+Ew3EZstImPEVkdO7Baqr9I39m7iVvtsBKdv3M32vbz0zJYqC19jdu7Lb7f88n
3CC9RgMGMKSKvcQCiNvvP4Lq+NU59PZlKQDVqL8Jzy1IJquxUbWaRtsjyBR3aLXd/MDprXa6c6Iw
AhWi4fhqSOHqILR1pIq+sDqbwEfzp3Vgx00RhkyV47a6z0nXi/6Qw+JjlqJU+LA1tTQ+Eg8Ncghw
e7hft7ppIHwpGQDVJi/rh7Jqb5+8Chm3BWZ2V4fLnJGsti6aZoCeN420jyMPYXWommZ02W2n34wm
s1o4NOl4Qf4W6/pUCGAyyDuG/urFgMhg+A2byt2oL3JYHpso4m3guASCeR8Rwvp4msLSEl7ElF8+
6cMuQI6w1/LztV6qw7M3M7jbOFSqr/OT88Z9+tW965GJDlg8po3EVsYKkxnPbsAfVIiCE7oGIVc/
qy/UcxZcq5IxcafxXEJMXOO22D5e+BzjYYu+yP9iNg+nc7wQYm+B6Mre6NQR6S5/ZiuzEueRmVle
F+PNGeDd7FB6+MrWddsZeOBGj1podY73gfXFJokvRdsPiJrZ9P1IVMivJYscfTpMQ2/MSPzKQXvf
mtigClcioml+vmvEvoa4fcoLSdky5uNtk5DTuvRVdjnyRGWAQp/kpk6XsKeH5wYo/4FwYV0I+plw
U/ZG1ygETbEgMa10kP+mI5jEKlrXfBoACSgtlXqfO5mNX8m5ErSMhdn3T2+URojaNlyiETybzwxg
N82VMUbEZvwf/DsB9I+wOU/dFjFycquiAsymMksorfkTvXZwgPak4V5Ya74sqwxWMVDDZeWVTx8q
HpElErurb5puGHc/kBgsgeyrNvklrrYc7kXZzqED3hgroSRuapjp3YACvmFbAfhXtcrAimgb2Bl7
G6FvhE4ZuWUWa6VjMhMkyY27wKBJeJbQSghp2AaFEgYPlFUcbFrmDraV483yhr82BDTejOQgolKg
6b1nm4mZB7tZY8GEyE/vxAy5ScSC3LMwiDP8D2m8kDrILv0wdJH0fSysb7MD2KUCch2xfRGr+o8T
WBn9d9HfClSfwfSo3iYo/gzlZGChjivYa71laDmD3hxLign2S3V6NwMGc7jAv09vTeY7uY+j1JYw
sG7TdXViyI4FBKI1rN18Sae5yX6foplIEKDcn8kDpDV/s6CyI4iIuYDyLrPfCnKMS4U48UdzppIA
FcEDuX7P5LS8aAlQAWPFB2P5n2FEVdlFbZ9qEENEjFd1sf0RIDWc6uMi5pKSrqL/lqMBJO6zQbSQ
n9Tp0ix6zLcPSm21hR4nl3ZIJnZ5xLynynyzRC0bzIZMw2PlRxKQzTH6Y13UXXDlkRpzkqva7wb2
J5+qwJgc+kHUhEefJa8hKo/mu1WLJbcnIh8ZKSuTVDn1RAsR5vTxjBG0JhsC1eA/NoFPjwFMNSdv
zitAfA7qyd2vQ8vtNxKDVrhWdt/+jPpp6b3xqwRidm+OunIAs+pV04v4UhnpPutdS61p2ackVRoP
74g/tP4gpNhsBfldnW7YQQStRu2U63K1vcU+T/p3AV19t4oHVgWj754t8xC4h/kWXdPNTVyuHKPa
8fJ3bs88YaYx21VGM6Wg6Ez/t7uHm6eGx1PqnzcJCbhwZpzkfCXC+DU37y2hznnOOCXuj0yO7nz6
4FLwxu4YYsnkMVQMFsXXqXCd5odLnNsGJExDNepEWxpFGK753b3W018mHcTxQBY1zKPGq7vYVgK7
WHsj4FvzRP9PD4AMWl62TqxKOa+QKc+oaJMBIPyKYbOlCR4PipcjuGUwuxq7nY/d97VSTe7UE/1W
F8KpVnb+aSl0feAEta/XU2kubiXi+k1yn1bUoF2+CT80Bm6sY5+ICUOrL5cnKZHWa9m0DLbohRIS
57tsY4O04lgpBBisWYpcYzBgVycvl11BYWFAza/Ttu7UUAOIoZHm8BV+9k/2o+/6/oxpgYOnZ+Wp
AdX21GGM2LVxKWn60vLcXieT+s6R/DFHj990m9c9kwBpiXDXLjscmM9Px/raTgRvPGMeiGZebMNc
yQpEGzaSevxaH/yQm/cIilOdf1rUj8unsDNKvzDX8X1l62fiE98Ry5CGLK/ju/zea1Foz0jPgn9j
98vNWfY+qx2gtayiROjZMfaibXbZvZPpsgKyAJIrGKyK/B00fRxWZ38rjZ2bv42sLSZ5MJdgfwOD
N1API4cQOBB6VKYqfsReNNJoWjwWMGw9VDLVga6+zq4y9EtQ/yx6/vwPGJ3k7Oew2RUPKQf6y4WJ
oz9imyy3VuH8HK1NfIG77UmIh5b+YiwAEGjspTyLoo++1PGcj5rMDX7LB1O3V8kCGKWSFyx+gvel
Rdk4vchpBGeWYivJ2mkOn/OHHSkJsTzyP1iLpkGref1iEL3aJxkzdKK+v58bC44KxICotykBCxhl
BQy6VhszmimSw/DtTUsKRzWjQy6smxu0aa+CWukKdIg63HZyeyuK+q41993nr3O1pcZBgjQzk+xf
erh0sbjJYbuuLEDMbuxRkGMqUX3h9uceNyGG6IDlGLbvTPMVT0o7hMrpmG/POmmeiit8yvFI/5jr
paRKGrHPin/aAcctfL493ExI7/IUrOCl7oRZLWmoZkxuhFnezTt9fAZui3HZD3N2XsQH8WIzJ4Gq
ILtet3/1LFqz63l9cSJ7dHnmrplISx9LYfKHQVPwsQux+u36dObpQYa+1drM58ThR8mKSI4ghetE
vzVp4tnywU36qaUz4th8bIKNB7RjdzH/HZSIl56KJJHUavjOp02Zbcmx82mVwiVghq2tt4qVR42U
Wv3fpwlG8kQqaZtioocPrq8xQFu0ABvvpiP6WS06d9GepKEPeAw/xJ6X1D+1V8W98VJFZCDgrlRx
A3Dq7VPL7RkwZsqBwsieqLBAXmipMjzqQmS1ZX1vs9wWc3azn4um3t0VddumoDGXMPIXkVFQdnos
+HVsMbD0gON9RcBRsc3phn8Dgjn0lI6LVebu/uVO/nXMYtfHjW+UeXdBPVe7Ml76Ksr4KARCmisz
IwvXiYpZ8+byiIRHMPJXTjLoXbUdtQOTm79vFrZwefbyltr3jU8KRy0eANi6L4YqEiw6gwsYB0zR
l6vfq8ilSvwCjl7Wv5OlksSg+weHZ49dQOCYFoqG6fa+8SyxtYw27MpADFiIfg9tnM0xinjafe+0
+4grQOiKemnLL/1Pgo1/1pVw+3FiF415qLKURaQTwaws+NIDL/pO4RVaDcrrblQNTIluLlqy4jRZ
APpBLZ9K5oeETW6pm2kLBDBOcICEQm/HDak7lw4l76+i+ly6qJwyHotdSPInvicYKFZx2Bc4xudG
JzBOaOXTkUWlBsj9MMz4XhaphWX5MWorlY6P09s7YIz57b3VUpDAQtHT83nGFe15FNkItZGS68Wx
tpPj0dRJYFuzBslrNvw/FNp7/DSTvYipBZLlOsUwK3pY/KM591xw7hO1Jt1h3Z/NdPZmjZ4EnN4N
Q2HjFNUsk3ZWIQy0OqWcuM4tdJx0ZVHJFVF4WAtLoW8qMiJt0unbbbiEhcKfldQ8k3AiGOHD4kUF
QNe4epkbdBNh9GjG4ihItfqKOPqAzdt6xf1LxwAMu+CBA6uPF3CZ5UDlFwtEJ+2F3bFDur+dkmf0
QWlLV68IEW7Lbihz8RqsxMv0sVJUHnyxscppIlU/PfVS5NCFGniGOqFcqG8r6D7obO1DvK5QAClO
+Mr0ZDlWZxSNQZkRUow21MMIXzaIXEsgouBLttciOnjW/OkFFauP+9TMFfeNgLVdhhPQitmjTIoM
I2BrA4TXyA6HiQO+8x3gw0eq2plIfCuUW0C6Mc7U2y3NE0RkkBHLUzBEtrqbKlDl4M/wh2CPTwWr
4T9dVRPoNjj5gW95ORqD7T++Mo/KnY7CWztC8uKXasPs6nVxy2NvnPGTWNFaO/AmE6hQ+KwIS/lZ
tHKQleQi4xVOGyalwWlyprX3SWiY4nvChfbZOeS7cRPmKGMFoqk/pzp3Yl8zuOPFvuFgZj2UUR3m
o5emZ7IBLFz4tKgQ8xxxicHZPdrdCLFKBONnF2k0xXdSsIIDwcf0L/saxRwf9rszknI9r+SpPqfZ
PSXlVlrap4Csp2OAOR9dX4Wrk/ZvPy3DBF78XZZigtXU97JXRvDs4W+uj1MV9xAPG2Hib2heDJf5
VwS3cWIarok6yJdPqkHc5AyAyNqVO1S1Ip579KLnbbAGIniOYo+7IYGmb8r9Y3DW7X4sla0tnj0c
VUR7MihEKkS8c5XL7ArggbrN4yExTXA6TQfBKp/RbYb6vrNJO9CWJeGu5Z9Nrpgb6FcBfZhq+15b
XFLTVHqHRSzwiJCESkmBb+RdLPJdMUNF2YrvTy7+XA7jHpQI8FHXzzHzYslPp4qNLb5xxDyQRU5o
zTj7UT18X41XgQtyDl2h35q6lOaVRCqU+0MAm03J8bUZhkLAWPm2ebcv7opNPEuLEItz9Y7xeuy4
smtp3ixeKd+VlATQLP1aXHbYqeGP9btnFPzUmeePUTbJtXyy/2AdRWsz+QdPSsSK9GPKbYEEpWq4
gzZ8fbIxqy8rjJp8WqRob6OeMz5/6IRnoVf3k5qX+1NsopAoIJ4Erkxung99qTOIi+9re9X9+sJu
ftR2JwW1DVmbjVpHxrRQz6SafsagF+FvY+nbd3lLwBOP74bLvoiItwCvg3A69KJigtHweLy1udOw
x9yx7r9wXmlvkpyscqrCMrvbeBNE5GGjjjaMRWDYVVrLBSGttUkVK5tQCmcIXalV7YuZF9pd0ue2
6oj1R33tA5aKwz9JlLDMBuuTKC9/Nj3TR4NESuAzL4VK3VNVrrmTKkU7uxi51DQ4uwiW9H2FgWCB
Ad0iLCOBxXbbewfxnGDXpl2lwpptLJYztxjf99yhukpb7wuyjYlKV0rmTla0v7eBDgPP95CKpb6H
MoEwW6D8uS1XCTAU4tEXA6r6L0+xvpJEhdzRSodn8WrqVajTwIxae/zCR6qZDByBwLQ/lSy5r6C7
VCdTYgJdp8A8CzjJfofmUpmT7iaAflOB5oMelwmuFGXYIVnPZRFUgz6TAm9jMXt1l24OumEhaofo
hu4iuPCjl8O+xhr0YnZe7xZC8S7z899d6R2IIQeiSpbX6XLtMFDhleyZqYJR8m7wIfokEivSTKqW
agDaogrkJwzihjuB2BS7MY1Tz+aYTbpErrQyl5JxmzxNwrpSP7UGUhGJGRzakioEGgZdMGjmDutc
X1g+vDtTvyHb7oAPRtrXFXu4s3IAgfjyDnMHnrwWbCdsW+Uy4Vxz8UR1Bo7IYcI+JJrO5b7PnzYX
G+00Ezv/o814PLgekn5vvQUzeDvhQ5DA6iuUAjAcRfA/TP6wATYDI81wsLcgSglx8N30dR3Y7BN2
uB9I6d431xsAJmKg7CtipULAlZ0g4f2zlrJxEW22ncrtNtZTPrUSHPetPJ2qDdG7EA3BPQNLsQFU
oeGK9xaXiMiof1jwwJDRKwlOcM/zbTJOBlMuIZ78mPdLrp2zXUeUNuQcWWlCm8gs/N6apB3vI7o9
g8Z9tOI3p1UjCeYiqsgl4NVAd9/lXPJWsKypqKagx6DiUQKX+cqloOd5RyfW5aj+wqAxeIrjTzww
ns0yALJTpe9nUmifE3PXvn1Ck4IhoE1Vbcj8ZGdLX1V1mmrKTHVRJcMdT4JZ6eQJhpUUE79p/IOz
KQXu4DFXsMRYZtZBteHaDcAM2kR2at+maC5fG7z0eWd9Gfca22ZeA/YyUNglPfpVxNTiHqNgVJEc
mA5qLj3z16Xt07HHBqlwTKP84j/8HSBcQ7tMh8Y4ycBYoDMrhxCwhKcs+pHKn5CDzHi1s57IkI2O
WTstQ3GoMMBAi45e5FpugfTtWdReyO3t3/hvvOBHvTl24sVi7E98Yr0JkmMhanRqukH8kw+Ln91T
LBkP4g54gyp6jHgXKhshxYRLdOvFVNhZQIg36+bPeK9Tb/g9QH8Ezyy/vxRQK/L4SRxJdFlYI0HM
s4X4BFBkhayd/2Ybkrwm1gVTSfOk4JE8LhCOdid9viS/b27ideAZ6V86hjXYtnkjpL7rSigOVSrB
QpMQePKSCw12+rT6NvzMOnMcTpfJ+U1DP9oce2wIQJvbLh4K7GJq9xxF/pUU1fdjAzQCnwRqwTJy
mSgLhhTqZVgb+rj0TL2kDGbl9NuTDsBA87uiYAZpnyeTD9Lf8j4DxI377G51ud4gD1EzNnMXGmyL
7YA8EQNuG80pRW7gKtxOlkf1U+ryyqad4xfUZI9G94Rvfw2SKoSoZFmCJd/5ffWW2iE/57E2wkJR
ESSsOmm3cQ/SWycmUX32ePCu3WtZYL9z+zTc/s7LMEg97mcl8F8MEtKk5/6GLYMXU5OMzZtGDTVy
l2HsArvxwJPNKpwPH3oBLslvwVJYufVwXPjCEDUvi4noFNdxgUXaYFhXdO377RUZmeH/sc/FRBpR
6kwjVhzaKLZKkj9b6y6JvlWiKmmQNgxcwqC9VpgpWeCk2R/PgaeCRUt+INT9dgR8Me2MxdffFmZ0
OhDUTfSXiF+SZjwT7JTdNrpaRN3yTeRZlPNI38929v4AFUnRT4cGM2zFMwL3+0Waattz+cKO78+f
ByGIIm2AkAbmD3tcQFYlOOKsnttB6Pkc/iVPWYdExWuDKZ2myGrkXHJtSB+g/1hqGtwZ4KulLevT
q8L8vtlgleU9bvV3/aoQ9MW5gt/jiVfaGPYRHdVKhRYDKm7Yv3dlWyHSBpXLrMG+pkUGtKOA0OiE
OxyPsrff8ruhrTj7bstD/Xtka4QzSN4dC05SMgd/geTg+ellWZjgws8XuUf1bxXVZlcXWfVjflq8
rEEb3BPMrveyf/6wE9w7RmUDdsTyFoNkPJWk/bWbMiVeL8/N2nGfZMTI/LrhgtNXacF9XdpGdq/A
F7qYEMz/4eZ2J1+lOeXzy4g+/Qb9lKjwLCQ5je2Hq37NH84aO3YxQ2PNgZslvei6pCF5nRL6zbrw
07qBhFUJpFsAMl/8zIIPQZlvzrcUCdEkhAE5L28xXPSKSzcz7xDOEMpPkkn7OMGHUln5fhQrxvg/
zh0iiTd1Lo/Gq0YuiTs2ELjPrHY91nvOxf3sHrEjWiag5AfGfUVsXTApD0piBunbrOtGZuiDp7s2
0n5HTLuDK25RC5WZ9kMPZ7VISHT2FjaH54cAkGbAjHKbAGsdn34FpyGWwE1OLh4LRNHoR8l0wslb
LGsw3nq+EjmP9eXPz0/FZnxlQECEVm1Lt5Ho9A4Vys3tBJlW47boNYvYhzQQpYFxgWdtn1diO3Rm
PuvUDrRR+ez5ip+etNitGi6nVg9b9XOAiFqC+qNnwPjiV8Xg0zWvrpQOly03n8jlHaJJ/kSvFXNn
RtE2VhQOHS4b3JFmvWCGJRy8sHZz6UAZVJEyb+etSWMIiM7+IFkufsA85yzIeKJEpmnyR4TIWqsP
OHuyhuXgbDRgn+Rr244WamjxnLNNfEvJ/fZ2Ea64aY+UrNNkpWv6ur+VbWNRybnJnaCaeFwU9qSU
h7lE69bVkC79wZa/QmxoHtOFH/Xkacm2DsQ2XCgAdf73CMG6OG1hSgFx3uzsHp248d2D+bw/ucu2
HtW+2T3Uu04SepSeMVR+h6hrkS3LQ9d5aQV+W6elTtmedwj5Ypc9mpE/f+vGwk8ARZQAsf/yxjHr
Y30+RhpBCiEp0ftTEF3B3rbhpT4FuMQblJHupDBbN6CCqPcU0Xxma0eGWZr6SYv9qOnpDspW4SxW
DyDTynKZBSd8WTJS+haNeWwo3TG1uuKIuC1l7fk5aC6DWci6L4o09hy7NxroxK+PYwwGLnqO1ACM
6otmZr5DoXhVkXNCb75FS82CzHpRXgsjR9E0pzfFu+0ZTMoWKcUIU777kVQxWqtIgPvz00s8QsSO
e9aZ6OJ64U9dHClvhcs5MDUnZy9f+u9bGQUDa9OUChe16QipQs0sbcLJOFoa2pVceyJXWweh+HZE
dHOmJwbOfqXf8i//IcltXvsABrDbfM4/8x43OHtfuZ24Bo9xbmaZ76QsZWJVlJo94cwSt9Zj02ST
xLaI6cXb03v5Z39JGENfhqVBJC5vgV4gMR8isb+gtBRKbS9c83PCPme6wST0d4fPLgUgMjxfTJKY
EEbvuNaZTLecbQq40D0NAtoSuqD4gKEv5XYjPJVMdZjiafxqoJwCSjUh6WQTfVcErcOxgqL2mz04
qS0DlfEVivvlLY86PYCIlA4cNwMJVIriRdvI0W7F0mVLgCr+RTTuWNEyUKUkJ5vyaOPL1mufGY7p
pKCQF+guVdXBBh0JrX+eN5cMA6Z9Jc27iZ4Mgh9DLycyE3waFVCjtzsi3ZA5Dp/AWiqCzlI1E2rA
98gZTgAFHeq7gTAaDlvBWwkxcaaSTA4x5yqJvhnbR2LyQ97eMnITk5oBacubuAa4PeCtYvpwjUjS
kk+rVglCYdoi+3YJEl26nkYyKDI2QbPp4oVWnD6cERVhdaSi0E6n4ajPfRk11V1TY8LvqQOM/WIm
dhqhUfPwkkoCBN3TFewrYQ/UZR/6hMqkCzL4UuYPK7lfHaGHIZZv8/I82BvlWfrguF86BTnc6iHT
3TaMh6JEmQwJ2hDaxusbvu7Q4FzD425rWzkYRxr8323U2t8Ft2SoXf2v8ovjFzxrVa+Csr3XHsfM
YoofWB3M3z7HaX3PH6hDLs4fOBq5tF9VGmCdpdZs96LewBjcpp8lsK9qFCQHE+FoFHxNJlANl2Yl
4sEllKbg3N6Hy/5cTLA+w5QkbTQPeJ/lgmHvUb/4XysLSURTHCETjFJTonnHSCvAOaZ5gMxthdeA
2atZD8hx+l8M97kywjkielayTQBnUhtQuWkbgiyZeaS15WhNJiwUCyyZ6JH/IG4E69eeLet6u6sp
p9SnGW5VCJF3qWXp3aY5mFXcuXERB6r5G9SNZkd3Q1Z49noFP9QS1L8G7Q0HS1TgLBfIpWUAFdSM
RUXl6vtuo67ibzwz6buoI7MSBBpEZRcyzH7KYsNKUKxT5dwTze4nUooudMnYE95yp3FbY8vb1IAA
VcmjvNWiYVy4BhMRcdRhLzGO5Q2JmySphPqiiNqGb42RpyuZ2pISDP7yRELdfy6amC1F/FgUngMV
pENr1aXHrgZPKE9Np9xfpv4I0xPx36tvjFysXRU2SuCAVaaBuBCz8/RMnuUTYWrpT2qzH4ky9S+f
SpDFpFXMfpZEqj+WbW+44vWTry8VGUIxV5XoJvj+Jgfmw/BHALU6SJRWbfXVX0Wg/Iq4V34IhlzJ
fKwtGzvRs1zuWf9HJv56Ia7l7xuWJyXzlRJNPSMMiUHSP8oXCH0STp2Z7ifwwk6LsQm97hwk4TTy
hU0TlBe/qJkI7nNJkeQMee2ywjK36Dvzl7yPnYi8fuhysT6io35vUDidOAbakswze2Uo0ff0olge
VLdtaao5JefStjsYEuHmyKKSaxCeUNtigbiHwbRldsTJo81LAnlI8vrgQrSptjZLQ4frCzm6sjTa
J2tis+Umg+FjUxiujlgxhaFutt2PHSQAMtOIqowjAMRnCcD5Zj16a3voYWO15SBHjX4LhuFVdMx5
RdLZhe3MtbeNRXRukxv3yu2rN7p1DkTkNPi0CFhnlws69ZkHSL+hOUCGr0U+N/fOjRYclCgHVI0W
jPAdWdy+zHrStcXnzYOZGUd9XjIwEI9pwu0rZNSWWF92spq9cnev6m7OcSFwzzRg8sps4FJdA474
LzIdABjbFlD0hRVjMCnYne4BX42APjeep8y9cSJpqoZXGw5nJKXLFEDTviAPoNEB+k5p2FPxOGQT
cUwH4kI8FfuHyQ9kzPDUF7XxDUfWMrF6rlUF746nMzX83VEhIToifbb8U4upn3SAp9IaE5FbZKcM
NM9gXmcmxdjWqOEdX1mW/Ajc6NtJD34mu+ptugk/m77s5+rHyua+kMEI7TayBd1yMg5lgZqOSYux
dW85j3hGt8v4fGmGl+340xGRwIyRq0BRrt4ty4XPkXv+VSNF/I+iqZAHjEVSiCRHp//65S1Ictzf
BvdUTteLnuOj0pQN2bMIjuLqBQG8rc6CxqM/nq8H7iXJoLgp/0tS5/0bwM6601467iXvGbTCjN/g
Uj7d9q1hRRzlUvtwUbvXhv8nJ4XHiM58KMmaPWT8kW+oLFgKY/VZdD7/rOVNr5ppPda3Cus7pycl
DnGwsBWjnUQhCzhpD/hy+sHZPMjfFuVl/rA5AYko9W76QRBwITSF0I1JcjpgUKsCHsVWY5/TCLan
YBrrRjWi8f/d/GhNn1aOHKxfIvi95AwwyZJe88G6JKxLW3Qy2I/RBOcLxwIDNwxsscw65ZdtntSY
PgC2Dv4x+uuBEZksMovs0Pko4uR2WZ7atksPziSxSj+WLKwEmEDPBSUo3j6a4wnVzzFMUZnHHNFD
S2d/FWPDSYtFL6/rYtlc25qD+pSd//3X+oa1IaJZcbzgsLAWNTeISOaSRx6lEnPoYyHik4PvNZJL
650ZE3u0vGPIKPw1As4PwX9ZinXEpm4N/LU8KKQlfHHCBSBru//K1mOvC1wnTF+XnAA9onmOJwrq
uma8Vz2I5ZYQESr8QYe7qRKP7TV/SjtUiaMYMtttainMMr2u3f4BmPiVMJ2WmZyMkmSXujH/BG01
Hd5Ru6ZzJOFEiHtv0Y5n1UE33yZ0Z8sxmkSLo8CSASGCsu1OgBHPpsiu/SJGz9gqf/mWjU4PnezA
z3nO/O2MPDUlhLQhUhWths/6Jip4ObRqA8aOlGXv2njN/mQe1pigD7K3SDCTz8iZ6VZsQG+pgrbZ
Q4cPhm+67SRUEDcHxEaoAPD3F/vgdI5g1xAy/csVw+ph0XYy+p7uJocEMN0BTNUT5o3E75hCE2zZ
dZR/k4hv4rG7X335GfOqLJNeD+XWl1W5VUbuuV0y48ixB89wXk5EXmo90ilAUyU/5Hi5Oof2ZOW/
oDSJymF5tfyEJOlpjbacvpU1/xqx9T1QdcrYYKgY17wRaqcytCR5xPLfFG3NCUZtkwZ1Kw2jI+6N
vm2ZdGXqJx7QTLbwnJJAXb2SHkOVw3I5SMVtXIZ3Ash5NeqriK3OqWFgZ9s/zyzZIAqKecBsEo5P
il/YrrJLHbLYzb1NWgizQ4VfxWiKZmNoPKhx4rbQzuYzk355PH4eEpxRyvR3P33P1Wg6M1ir37hz
WJpOT62TRWadftWRFC5iCQp9azUjc6nRV5kWwXNXfQo7UXhqc2uY52S4UIXbZlKAKcTQg1dHwSYr
7HZhGAAK92HlDCQ2vg3w5EarLANlgjHANBAgNC5appznG/tGc5cSJyY9jdGmn+Jy9QGaIFDUaeLj
Kt4Sg3UVPmHJqTBg/V54pP69FoSqgfWSRUdN6oFet4r+N3E9FxLDvMcsP3t9Q2oATCTVTqtecMod
IAqBYCgdLqrkMGLDDl/O6Vx/LkEZyzQCAM+q59NueDD5UgYKtBZcB/1esGcTs32tvS/b6p1W2jFg
29hryk/J13/Kmp5i1CVIGA+WVV3oIa41e5eDg8y41phOV7CAZV+ja3nya3omLop7tSrZGVxAZfOF
Bnn3sVEzOiGh+gbHfGUsJhnfM5nvOqBVYYo7LMPGGRMXFPkdhXAw0a4GZCf3s5b8ecyKzfvzlhkA
+Dg9f+0vSMbF/kQDaGYhABaHCJiusLVqOs4Gkm3VEGV1H8BMufRHTZdYX1O7aNUKhG9+mRl2V8pa
Yb73/fJmy3uLVG2/d0dPEF3owfODEzF+pN73GS1d0m1rvYEFDabBK/71UnWjJJ2upszDRIn6UjKI
gbRFMSD2tEZLMyLMUjQYOkT6Xkv960AbzhFBTNW7KMFre00B4swJtBSwwwFAtgYgWim/2CBwWoER
XsS9wo/9TWQXKIcIE6sHJuU88r693LyWNsPeF+fJdvM+pSPlmWHlsb/i3c8CEvYw2G14l2bLNhVv
LRWKE1jWLLD3od7+UFph3ib1xArbwtDe+8D56TCtHBWTPfzerdoSo+qzmMZQxgxdJaem+egBuJpZ
RXfzYOH5KbUkzNi5B3WMWSeZadVzp6MedwKAP90cZViX2oVGtY7aobgLbzpJQg2a0MkFH1KsWPqV
8c61wfJoF7+tjzzasgMebeA8v94uOJ9P7iUIfPygrT1jTpQyJKpM7qrD45kkxjjnYcCmkzzIE1O3
oA16s6gwBmvCUejf6gWV/55C3Q/D3GlGFxJMR7KihGEhkdP8+fM4d+mKOXtIl/i4csZ0MqKAPkEJ
UFsVV331+IVR/fZz3epSs/xdBGGVsQtmaTkN6XAYk5Ke+uScjObQWGrfwjQd3Y3x7gArOoUeSXm9
Ci7i0Q++wyr4C5+ZjVmdvqZoq12DXlRco5IboXk8/Y/IeTGhNtdX8nGOErDlmZqFJIaQG5QvodUv
S+AfF4Xs3pgnXHm1TkA3ZW0YL03gOM9fCcCCHcpH9EvUboCBVj0shahARtinNkgkoT++GLXMzpH/
dWZXUsZDjywVOT5Y0TDLhlSdVjpMueGF0Bp2YQLN3zNiSEWX1ypP/uEmmUFjovWGBXmSDx0xgPGA
5QJOqb7FjxOVWobaEP3VI5EEhFRYaOxsarkHvofd2nbmc5mbTQtiZ7QCGLwaQsFjlRtvt0A+NsHI
/bQrRZrjpOQUwSr7VeyBTCyDDNh0Omj9rFaE2ZQZABtQb4m+qeFhZAWi3JMHZjfHJbIcyo8wgier
J+LDSgELAYM5T5HYPUfpeZOTvuRGL6uAOOLvmCp9a+KaF68Am2MM8qt/JUqHUaurMdrhXXEk3BJe
oUs51BanbrKpn3M1abbvvqwumUJ+6XR+Jdixa7yVh4QwLkbWl5e1iw3eyUH6Yd2U0d8uPniMYW+t
brRVX4cxb0QrmDLBn6OQpGT0US9D2f0Ug/u3G6OmkGGp737qixfGLWljl2DjaSXiYl7UAI6hmX1A
r1MMdnCmTZVyQkuELYkd0dLYNDJsexhLRS7CdgyLW1VT34z3NctjeDhJHWzUXtvNybRMhAml/vjK
eYopw/YPJpQhBQFDyL9cBf+UJP/AiBbF49mlyozwpVL4po5+fqOF1vvO2aH6p6J+OYKVRkAz3Ner
/U95Q6K3eD9fZQZpl8ZiFqqLUbFAW+BDV9zMy3NwXxRktP1KDGGx8G1W8X/zuIGz0OLcJczOSULH
IS59lPPam9CupulfNdd1b4bv489pNS31NNktcVCnRf6ZNI8G6KJKF2z73n3BiH8GEO5Z1/DjmbRi
RGxUsSvmy+rJgoM+GMUHIMNKoV76o6hbuL312uOTn8K4eW2SevEAWhQJXKNRZ4kmfIGWsL7OV+Ak
Y/kKc+rF0M6h/fKFica8ocpkyDfYzjr/9exIJIn/l5yHOZ2CSdAlpqBu6USjRTFaMDPZ41PIGeFp
GomC7MpglgEw+rrLJTKCbgd/JRdgWpTyaO/8Yc0y+vODwrf4yvovEQcaoEoRDyr930Q3ZM9fUh9d
Y8GWeT7h5j90X5xcltEtNxubC39fu//IqO9KPybPdlZSPf2YB5wv6ACqbKcuGlZl85bA9IydORxq
7meBd+YCwimggey36EzIvxKErnDa0GlX7oJ8JBbtrJIaJnSJRN6U0w85jatxl64Vjm90aP1PE74G
bi1FwzuAVLneJN0DFswvGojWqk/UN7HGaLIujNkkhBHSF9BN2ZrW1AVvd0Dj4dPicfBIuUp+hQi2
kqiy7EJnC4OyJKbxvd7R3e277PO+bavv7aWSyZt7smasc8QXUwxp/FC4HWQsXt/dx+CDlmVgiByD
+Oda4kD5ChEDNUb5xTT1ZOQgMDUdzrGoIxdF1RkgFwy7B67IHlisqBJetdRQUmPdvoL55ZmtLgV1
dOqWanfiq1qeJQ2ZhjsqxRRq4s6NjXeW+04qrJCT3IglX3AsUOrfWG/a/5rzYkfrXAYkbiqW5vG9
ZK4vZ7ZRFhT5I7658fQIVU2Z9v2HEQc7WeQx8u+yaeMEhqRumjnbANnH6W36FffdvPCX06canrpm
YwOI3DSFRDagHw6CzS9I9t+L5q7kzcKnbB1CpZuSCzoPBq86shutR/QHb4dUELKRBHcgWPFhbZk1
yD6ibNXHRM+WYX4NnnJo+9xbFD/kA5HxT+vEJ03HcK3uIfa1sUsE4w0PCb9gz1qzE84I7mNWRqML
JYNqLB2dOdes3qpGXEm5KXVZhjHAq5wSHLPtuynR8PB/bKOwCsQ3QgbyYfTWhckqZNgWAsi5VuIh
IhdlA70t2c2zVXUP8q91Mn8ngh3uhp4lkK9pTIaukBJfGiH9hLoVwCYeHZPwDUVS+7MQ/+0UATME
2DE3oiteLhVn3DkKJDong1n/vyKxvBZeTKEAMTYScOTNQaAcTlIfUITtd07Ql6HZS2lwZpNbGOQ4
fcpomZ3/MqKUxDELkKm6/DlKw227vV+lKh/IU1k60nPvxbh2Mv68fDMEvKoz2xP9IVclc3WXN85q
f9v0j3V5FXHBYM5NArdUqAEa8g/c1G+vYcePzNvc9jRvNpmk4f1Vz91ZAgigoB7ctU+8SCyqVO8E
yGFXVQGmTn/PA5Elxs16fPcLWJXWxG7HZX5PJff2gQr9AVV5x/Q2rOymuhaNlKP9qKl9qI7tgtlM
H4U3+TCe8RjIrdw1RBdDYQFfWcy1OgNZ1qtwB43JlPwV24YZ09uBWj2qbDHQlH52MFhltY+LioLP
5nv9ZCv8eZXGyFeTrFyOhqM2QHTzoM29pZC5zuY4w8F07ctAtIqk9lZOyBzK99IXSIOcjFTVpOor
jkZxsTB+v+Ozp1U7ynuWJS+d0GJ/+G9ZjSENxZvWb/OfAVbxYryFzNB2B3dvPj1RWK46bGXBAdiB
80r+isLZSUxZzIwHsIOd6fHYdB2bSkTJeQsXUqVhagH+0rGfbfekok8Dx8w+vPH+vI23M177zuFc
Q0dJ1yvOktVgz+T1WDf5OB/7MFlzON5f/prEe8bV9xudoxA+cdCxK9UcBZ60mde4ocFi/BtL8PbZ
JfzpDLWF2vzniCA3lmU8cH7GOFvWzRziuAMX5V6poBSLfi7D/VvCcvlv1cp4ureyN6/lKo/EOZVV
B4MbxwsM3uU0ysdZvPobRclrtyLYiAU6oQ80y+VhB40m/a3PK31NauF6HoTP1j/6hkwpj+H0Ynxf
5JfCf8gPcaRztUKCdVCYNylgeI4MPKLh4kCFBsVUjaORwRvss1MK+0L3twZpQ0OUFSxgoW6JPhXn
LyFQwZ1FTXcvdlq5v84P4bmeXWiZC/uT0p3uZZP2WAMmrsfo9X3owXZhfAE6eyWU1KErk20Rs6N2
urcP//8ibbssRGT+UAjzDQ5SSO70bNVE43tVPCgFmnTm/nbbR73jEP3ReJUqHrn2elOpo6YtPBnT
yUR39Whr/aqBNSXsxxquhF5zKkaazaSyO1RC3ATPylXFJpfDGFNZZDN/87fLLiUfSLD1pjwympSS
NBbeyr1OGN9PHupDbiA3O+MGgFLCkH2XwEjstfttIA4ZGMrJObdEvrgJC627zU+VzZN1bskHbMde
QvynUDXV/gUj2eCqKJHZJdYYfXiSmy6PAVbW9w3cYgWKdTnCld8VwD7DOGoe483o/8soy8MxCzo1
GUYBZOAUS4JOek4mOZQgZZgqWQaLBFXqz60dC0BS5DZdPsIYBJmHjiICAQFv2N72QuBGfaAU0jop
dBM8cVCv37lf/sLduUf48af5WivHllFYIpD//wsrCkETts9Q6/IeLFuSjLSXukjyacM3rEnP6bzu
WAZ3PR6QasWovc3KJMzwdUalXE3fb1M42IhqsDlSvoX3BH5zTj44hEiQzwvDKV4d/pRZpZVrvEcO
EBeS//lTVPZIBrVVwjJYipMhtDpR4tfG/GHEXmQEuPwRI4VHNttUJnYoqEZwxSqIXf3FDovECTSI
HD4wqtwgkWTiRBFBR+Yo6sgH0+G92h4NwEvpMJhRAXqL0/8T0sVJLLG0Amz4trhm6S8nOxO+5tyn
TgEY9Vz+D65lcO4teFD+bso7z5eyKMq4iosmTiPuMHJWiTr45otyacwN4mBpBASEE1QOiP2gzLn3
q4D0X2S8ImCWejq5vp2Vu1rQauRKeK+SZ1rKuX42ui4kFyQejfSUTaf34jAQ0+C/pSUczoY8N8WR
1amz6MiYSYZsjg4glHwVA9RXQu6TNiIl8PEv3ugbF6H9/HLDkRk6XDPTH3QB9P7Y9E56ezZ18CwU
Z7YC7zxux8GVtFPrn8H1FaBrxHU+rBbl3v6MbCgHycbU4k5zfkOS2TgzgA9QUWDXdIHIOD2jis6P
fiMcYlqEaRD32PNj+2scd1M1taUiD0A5206oyxyCu3SalxF71Lw6oAzY73mhF11BTcQYnEWnY10R
PzybQ21YUg4DR2IX4J0ofItUux2C8nompyD4DTuKyfhSwiTdQ09bDGnhYTYLVS41dnAnMzjZKz90
dqwsL/G77qV1fRg8RlCJt3rOtuRcknY4U3q/+CeOOhHEvoZccWy5YY6UM9PT9+MFc38sfts431/P
60HrHYGm1nra3k40QWFJEVv56jpzIKfxuBCIh52648Fb+YObugcQun1jINWRCTKHRBCe0u6N1DRi
wXWSyZvb+csDHvAwcptTAY0/0ekqqVo2KTlR1uivmfEg5JgPH5bNMvIo6S9QlL1GARBfYkAQ5GDN
IVcEdNaStnHSRme49+lTIFsMw382P5GM6Acq38t5WTVHJvI6WLZjsuX3L54sGoL9C+EnqClwNhdN
H+9UvX8bYhAg3wOABuu3EmqDM0mONlL99aqtBiyodI+zOPO8pC3F+3j1F89FLEaQOhrRd4QZUshg
DSsK+VKSg7juOksgj9cIXoi/bBeAtlA8CbtFRnIDxavab31hXXZkryVWCwVQHv1bJXmT0ONc44HP
91UUD5SkvCraX3bmsYNUtS3vqiA5YNnmgU8NEKAt0vOGvSyQtb+dSq27v1ZgjOhzdLr2W+ajBF+Q
6Yj7dqjTxN7JFL+kkxYF7idle5MCjbztVCjCH0epRzbFYmBqqBVkWhL/YSAARTcTiIpd3d4eJ0at
qA8oiLNyuhvYQz7uhneVFo+g4nzMoMsvHT8dHWjSCm3nvtcpOA8qiK+IB6inNCUCtwY4uU+NM9BW
LMgQ7CtzpxMd+mJSC0hXdeGV+OoIcGnA3Vl3h7HUqfuZpKp5I/GyguRZJ4fbjXE/5rHmyw6LMKLB
ZITRFCyPr3TwFvvSKzGpy90s6m4Cd7qWPjeUEJl4D89DR9tACHETHBRm5h6rH/he
`protect end_protected

