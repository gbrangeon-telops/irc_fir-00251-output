

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DYkUg37UnVRJ+X5v5iFDmCWObMw/mUCrJuxa/Cr9wGl4FgcJi6OQesLI1M+aH7+emQJssoNWrh+N
iL9trwbpEg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Vb74X6mc2H0e6MLiEAhBKZ84QSTgHhg3aAfwLeb5H8AGScZ7UqNDKDmI5IhuJ/LPpdHQCtOent5+
I1p5tELHTH0LzN6BILTKGZBdaGJ2AKKoofyljqaR51srCF/ZJLUOrn1XUZMkdlutYXGikghh+zK5
6+/HFEYyz6zhpfFGpAE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DUY8u9eRLqeXCDG4E2/8OtDIacK06AysbSio1XfMMKnofNQFNkb8eAjngrn4u/YZ6G16ZNMG7YoY
jk2Rx2Q3M5GrNkHLNcW1r1FM93KBIPYna3s3UsOdPXI8u/gdrTwtTwv/xpFT5pO5KUummozg1ol2
CfVK4phP0ptL6RF00qSF6IA3NotRdVSf39i8Abyti2fNqAeVQtQbe8y1/1WV9RrHHqEjarv5sqIY
6GslwJ8wdJjPL0QS11gBEh6rDpndqUhWIIFTUrFMd1tEU2WzUCNSxtbBPYlWfpU8e4/l9e5xSsF6
weW3wzZvwjgR473vdWcupdpbpXFjQjfOA39+/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
p0GGQgjzPW+6PIUsMdZXTQnjW6BUopNyvt7ApHmGMwjrt0lKkYFdeq6NnHPNeKi9xrrloGAO2Tha
FhPoK1WSUQvFoRR4uKVUk0OywXYhciTgYL90XL5T7z6pvP+T2xdoDnAiUPoqzH/Ubhhi84EoGyo2
+zIDCCcTvvnznOBjfpk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m1/kaqW4ETEcDTOeEJMS5yQHRelnhe+7sXgpcKiP6lTf8NZHj87LtgfMx1Oh7TGMtL3OsgLwXKl5
B/MVSSTPV7z0P/OvFd/MWYJqIMAVI0yV4hJ8dwWC7KK/kawdL1h0Q4iS0dxjn9/392LJCmqkJJmj
TEThXH1uoH4tMKV7xRRg0/MNNOk8hPErcV0Sx7ZxMFsvJk/PuOEi0wzy6daa+A+gop4M475HPjAb
iPZ63o2focv37v9R+NETZc+LyDzZAZPFDxIiHCnZlRMpU+rYc4lLu+Wj7afASerzvuIcVvlJO0R8
MuDtSunchT2Nxfc8io8WUTVsWpkmP/zQb3BvSQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18992)
`protect data_block
926oHxKI33I/EzLP0SDoPj1eAJQvOBlQ92tvGF7AFnDg/DMyOirZdeaXInS06M6lvoRUDdeXcuvK
JcoVVIEjHjhS/VC5PnyYyqCgjG0w9ocnvNlTPvawy2O/bCTqx1pToxaXP7il0dY7sVJ+1KNCfXn1
x1erDO+4BHStuwBUMgy7xUAuPUCi3md9nxRHMWuXyEJLWjWZtjxyxomqqTfkk7gp9OLFdKGs5jH4
laPNfR4D6IqeDx2vcXdQNXeHBU2ox/s26zB/Z54mctxVZk3VnLdR0I2QVFql0NoAKl99rvy9xTBL
73FxXCJwTz6htMuHJOICsPwu6JU2SOMJfbxfb1q9K0jVWjCA+hSxh2kx5dnppkP3n+Ln7nj/o8Sh
VqjCmEk89dUrB+WwAFmyISG51xSnNqM4KFSTzoqniVkanPFE1YAMNUDLEISmRzq9ENKWeG/s/FW8
x3lIlRyGc1c7OA+/h95AjXJkRtB57vYj06vnGivz3Wc3n5/umiZRdR3kytjVdvDbh8hLaZbTSxei
eoEF6mwj7RzPkkjjsRECA5c4qxmc4WOZUbuviVy8Ci0jRBcaS7jRxdaVWsBcLinLAJA1a5h2gdN+
YarsGqsDjuEoyUwDKYU0d/V7osIk9bcta88f+6vv8gY10o9wZyuTfsHrzmH29WCY3+ma91VGDLVE
lwLGBbOBMo3qvKKX4rNbA9niXDWMfW2UhNevhhIOg2mchLM4Ohs5/7QZ15xVEcKz3mKXFV4se7cE
FzNyTaxQ6S4AugFmE/jmpvMW9oKUIrJyZfTRAqkIjt4NAFF9wuLpz6z/SPu2YZ0Uai4nP6/FK+0u
wRxVqX6nzbqW5/Ptf57WKAEQv9PBHu3e2aa3k8k5UEC5QwphrZgRGD3o76BwG2yasRroOErg31Uu
TdDvy5Ail9+IFZ+8KxTjQNSxAoa6b8+Zw80nzfqzM9+a8wuxExUr3MI0sNZE6AiMjS0LEmhmCYsw
XdN0OQSTrIcdpKFNfcxh2nMrOoeQoTRB/hPlDbAaWMlznlgh4Bu/YfI2/jhDU4vSCeosPMtTDftP
7PzC6UZx67L0/VV64Rux0YFq30fNmeu/oTat3Ts4Vk+bWedVmPzm/wKk/NqGKgC1Oj8c1gXYXI+W
600uhXbqBNkd37ySdXmpL1BspfTDgdrcqDyxHK86hLaQ/cVcJMyVZ5xWWOeirvilOjRaQ8EUSePX
wV6uaEqZ9jOwg13O1bGxOt8wSaBmuRtH2lS8qm6AYEkppEd+m+HMTjL/hfSNyQeugHNTzfboPX7M
4dCY1WCvgggwIGIRnzFsAMoRPF3N5S/3jXnUkQvR35ukklzTb4yWx9qexjafw0S4oh31sXq/uSoc
2dW5m6thJVexXHETWq52GpdDyxt/5vpQt2tac4LPhMYaRj+ahmhx2W+0r3B0KByeFHp3abtain/V
TVKdElajVmE8otJv9ye/mBHqu+DnvQOrnRtzphZZ36bqwKgX503jdOHT6k0MG3vdXzm6NKJNZnEf
ozXRRrA0TXhsqXhfyklPYuHNsMknxmHkfeS1y/ubvn8g82vc/kjwadFDAjhmUGtHZoi9oXduxf7E
+rrkQrWViasoTLeYV82+YYEnLtGgY/iCJZXp+oVnt03pe4T24ZmBuDJ7OaXMSwF5foRGFSxYFVO9
ni49YvKn4TDpu8s79bkpP8FIm6vx0Be23H9yVWnWkDbwv2cHubYYHLGGrN6LH/DtAtOaos16P/NT
/no77LAomXvkR4rejd0IXj9ni4+oUNdk7++CIz9su3bSkiOe4Sg9A27RW210dbkJqO0xm7wI+/sK
Jk/FFYMFdK5UBhD7LdBRirwM3HlluwjufceOLyHaJJO7VMrM7D6RVy6cCkjNr7kDBmAaUouZqyYT
k4nhcLUQblZxFjNhCVBovrr8FM2UBSTz4MT9Lo++OSMKGWS9M9qFA8VcaA9kPlyS9libbH79jSP0
iDablqU9LL9CtMwWmFURn9W3SIOUxRSsKjI8Z5/WyAlIIDfYAHOB7voNKyma9C03jk1lyDoNHCy5
tFgu9YO4Ov5HJHzu/FzXxFM+jxPbluu3+ZhDxquuQOyyHZMoi14ZsO8saUypOM6rjYcUGo4IkyFo
etedcuqXYl+zdoD1tDnBQbRNXg3Hbx+bgED+i0didPj/lS8vJQHoYjlxqiimsbq6n7IhgH8GzPCn
jzdF/rAVN5Y0ZPYqu8RrQSwy/N4cbok1qA05WP1NVxfaOl2vFJXkiX7QrG5zuCCVl+W6iTSntGpZ
2EQ9ovzSkZIGBSv5DTMp8UbxuFN4g52aUcRIwEEtPjDfaXLR8CugStyWKrA3DqCbk+crf5MtQsJ7
8lBaVvHLTOYcSdRIMEvhN1EZV8NKTPGWs9ycSGp5SI7kV6AD+uAGfLM/kuDJvQyNKSVv6Mv4cqtk
JLFSnfLcoYNkHIIkl/u51FAL3c8U1oOAPbAO4X2h/DN6gOyEBUyHW94QgBTR7mTfGCfnGpbqne7m
A35IjIMDMCCQTUGv4jBIcUtPvL0yvaGA5oHkJfxxQNDO8vm5H8lJZAXFwadZXBSTP8uepSNUXH1S
D9TecgkoDvDMf/iL4mxuA1ip2FwoOvi+7Nl2F+DYrhQocFa6vmWylh72HigbI3Y0692Ok9Xacv3w
eS7mgufmGreU66nulnUewnazbWwhIA55BZrPdRGln3N2Iyf/AlgpdQBV1MqS31LWB3yE0+7MpDaX
RgIlWqVV0aKOVMHLf0dRiOezUl9JD1lXlVjr8H0vKeAd7AKa2a1Chu618u0nnPbAX4vacFnAhjlD
Ak+cWNkT66vGalsSQuEz7rluEOmTboQFMQv+3aAf3gsp6L3WwT5BBnVWiREEHbxSNCdJFJgXgODl
so5a/rRi/Qo9WdtXBvb1oZtw0OjSx2TWFgjg79WWRI5WY8ud+yFBMQlf2ySf+1BvEnYngnaix8Ln
QaA5lppQDd7/MwxK3r0K6/QKm9/P+34QpmiBmKSuxkqBvLx+j9pUCFQEEHOc/j8c3ToPrzEUGYqt
j744ihdi7O1rGwEBeN2wC727c55SnZblY1Oc1wtHA+UUPLQxQIzqbCzFdTqVOrVONeh5hWAuzAaw
QoxFQdeCmkJ/6BA0eR4j7ZegsjOPWl5ik5eT5eyd+y70JN3BkhW4++PUfuJuw73XnuZobuhxuWHP
TVK4agQhY56OQwvI/19zouxL0Rk2GqxXRhfhr+PUsS44+LB0zKA7LAmgpu6Jn7N+NlTJd4dn9L0r
KcOywc2tEss+oPg0qwnT32gN70vGbHP5+Yi/2hBsnsT7d2BEL/lLkukMryEErJOP9ziApg+QICyh
aXdVpNpDdI5kyJ8citytkere/yJRWG/Nccvbqcsd5WRyHQ6nDNDT52AIMWJfMRc5vGqse7S/PXvE
Z7ZqKhZR/oxrsqB3Lq4h39Rwm0+MZ879xBqDuRKvbqq2nr+72aP/Ei+35xLtESu2mNoHIABbuf/1
Tu2JGtEdvjoTfySgn+8j5fX2KJlH5c9T+uFa4SUoFMKUYeHLb5Hgr34m5faahrjrqC/k3sfwzmNq
Rs91FY68+m9Q6M9g3Q5biIVJE/xcztp+di3IxoNC0YnlHft7RnxFxqrAtO/+TbA71avDD9VFBzct
w1B75xOAtb0Z4vP/xVYkW27bBuKDwhUmUECNF6lpbBCJYE+Mtg7zzjk3W3TuteADZCcpHlaxUQh2
cFsZHOHlXaML4oNkHdl9CTz+SwNH2339gosDVTJv1skwoqt6WzhI16nMCWH3lv2cQuSRlh1GRlxr
UkzN/5P3n+cKw42SvSQ53ODhec8gH2uEaKAq/4DvaDCtWOaq7VLwGBlQURMA2EYoiNViHfU4v2Ee
y2KGYTjWI5z6OL/tgytk2eBIle6WmMIJoETLWJcOIy9VkJqGPJylKWcrpTLGNF1I671TtIh2EDiq
AbdvIsTMudgiGvmr06HqpNcHDQFfLfitpmdRf7ErVQToHKbcntZy9Mv+aMkuko2264mhfSB0cypw
CyZTN7jvv018NbEg7Vp3L/sFuC/hMu3RdvdgMHV0rMMTiXXZhMDI2aK6WhHu4HD7aOT7w2cgYuI4
krxL8dZbfJmyNz0/clTNSg2gP4p1sj5z+PR6Kl+7s96UA3xrf1AmOB7YsiEvBKRXdqIXI+q//MCe
moM3vHXWH1rdFfr8rSdtt8FlzUWhEW7c9iHq2csJgmb6JetmHM4GRpu7Wn9kPH5rUkFAiPJKv5uP
5XH+mlUNU6Tyk9yA11Bh+wX8ll+cPbJUTaRgQ3zYrsa9mnXBsXKl9w2pdd0R9ty15+bKkn8FJZQ6
FyonWb5o8bDfyMXh8wovIpYM3pXJDXZfMqziXWuAnt/PNeOx2RJowB0SLPSFfTiZsS/uDNBvIyQp
3LLB08XZuVtN8J8ZDwFa5SPGYWJTIFuSb8n6r/FLuJd02HUFhM0SSwtawJ4kL86CV1DvXrNTCX5p
T/drFMxVdzr34LzV1LmqTrAFLcEFOad0GiOYOPcyuCjcZotUzrk2GaiTzm4RuehPMAztran2eg7v
QjoU02zCs0vKHl0zwu/pg95wGTvEUEM5SppV1OszmtnSVdL0Ri0kK8etbLYki5ZEf/ucQ7ZUXx5I
jh7kC0zKH8jQwc/ukCmvOjTBh7/dawKba+gciQhWEcTgFCgMRE1sFQ+KFdnr2OsuywL4LasE+2yr
0sFTi7pBGwM0o1IAXIq8zP62TXhPpywviwBdrPfUkYhTvOWVzUGjWF5a9KzRzrmvMMdzjlOiCLCa
QfAtUXEOUkm/oouNxEL/nAxYxVPWUft9lsGyfKyNvTlj+yhwlbWpGEbghurHLguABZeszpC+LmSi
jwITSqMV3n/R6I668SBTutj7MOL/lGk4LCG4Uu1o9TJw2Hap9D9vtzL+QUDXudkxOj+ariN9QY2G
TKLVpjG8UcW8s8BWjRzMpF/0Tty+QOO+nQJGzAhJ9l9ni0jGHv0bAdM1VTWXleRpT/1bwK0i84p3
mF+PIkyO9REJCW8k80bNpoTU8M/tAi+Obu7/Qqz1k6wXSRkBkwrUg432c0sxC4z82N8NtXGe4kU3
nP1Woxfw8Dw8WiwPWDzq6+2V3MyQmmHe1mTODepV8ZDGydY93pwByO7bK/wXG/Cfl0/FqSNL6+5L
F5sBhjkDgjQ/2SJ07WgqMr6MuSt+H1ymksI9fiML4vQcHhcPeJI/KmaOuz+NgT25D6yL9aKbPrgl
UcEGtQuR+38WX45FzbKrFb6YYZcPp420Io2CsYdS6mQw1udcVPqiP4vBakU2ZZ7eGSJbkk+9qTZG
xPvn7O2ld8iih6gPaJWVwLIB8/7f8ON70fQHzmsNO1AotQmyX7dKHSRfLFV4e5t36V/SCHYT0hUJ
T5vjEo//qkwLY+XTe0+LVL4hjXbDBsz1T8nFbrsT2WpvKqNRDqkpCN/+wsB03sBmKMa8PCsCt0vM
IDo9uUq877cbFmxxrR3Qjiq+zandpSQvO2uGTGgE12s2YJf5+d7Eb5BXnwn6afb3bZgd34Q1Qfq0
Y44WP6mOo18JmRroq+153mWlNp9qoPVe43qjoRnspSDGT5xAxv0rmkZLZPkBFvaxagS6AlLkihTV
4MgVtXaMtu7LSrgBcdtXoa1R8maXV/gYIKWJjtOm/o54wzv0f3PmvXu9YKoh0ExiG9cVPagZwzKP
rfeUZ6cDygaZC7VrLaE93GiCdkRwm9gOMFB4UglGpuQdDCGjmUk5ET29jzIQtVyhvjuxBwBKcMI2
Y5TCo2NXiqe2PViDWdwliMjEitgg+JU9wQ6iplkBDUg0bORB+/jtiWLSRnGbQx8Pj//5XgM5OMPV
gi9vooa8OSQmUcbhGqGUmeXoyhB3JO3cU1s8rCs6OMa0DJLUWRn79gRZbBxuXuaQy1DX49mrci3H
8zGfuvJnfTOoZvFgGVklfLtrHVnCe5vsIoggAta8jJ6A3tavJL4u0GapGPXBmNdK4/AiOp0idiJd
fibsAoNe83+8bEamwNxTMOjsQFXm0Dm55GTyJgxmFdBQZO13niBA0KGLF8naq/ISc0+ngzSI7lAV
CtjsFYrbAXWtUVkBGSXHiZ537FZze3CL++ZCi/Jg20MfhxoZaSwMnkuslrT5oRJvYogh36Mz9qmH
9C3xNI8NUr1kEx/ySlVUp35v+EcwERet6C5gw7hV3u/a3rIy9PPnlE7NmsQiVNFEG4RfnNUyhmEW
hZmNfM66GtnkeHJ7/DWnBVA+4NWAg9UQLTCiVoagLjoltaCuNEYalzwsJpClg+lZK4ShM5UcAxeG
l46QA7oR2B+rEE1XOO8Fy2+m4g2ilzctFkho5jftn6KAsU49MJX4dOUShSSHyhF0YFeK+7+HACKE
5NZcYSDyIzbAeRK2OaYD+JBLG67K1CcrwPsqpeUTP3WUOhzg+U5mMxOhnFsIZERCGSrqruqcUOaV
JKBnDrTX2+9jx+Ch5WlMsJtXwcomUBRgw526ehcAfZJGU8TK9WqSGXIUsaTs7c5C+w+k+u8Y/mlD
3JBFqk733jMwjCtppaJa95N5n7bXqe9edhr/XAh7b92NlJPszC34iUQPnSIslVdD6iXbrLLg0VI8
u22LmdI51anR9/0PNQr/y+UI3GdRcRQN6BZ22lPqvSADtmwKVYzq8zclMUduJGp00pDo2V3NgORA
ELZZ2HHnK/AfVBQnfumGw9JNr511/xyxTnVPALYbXLuzoUEKR7UEMisHQgyPu3l8ZH+syMez6so4
Br1TXNILXHL5x8kOe1GB++KtNZ9ZRwQgq5/fb1e5rTvspjDWEO/mwVHQrFYKJb8gNcq8pGsVrEB9
PIKTCBBK8fcTKWyY5vbC8qiuVsxkbYJfaZs+O1mlsFPxbdozhE7tEiDT0NCBsAaul1nrLpuQ3Jj4
lj883ZI+R09vrM2I+RkMEsqXFyihRBb02tdteiK853qMKMfph7V4yJnD9DYi+aaAul22f9v6asUk
XmyC82KfRK+7qsWSbXbDyMbgh/BM+4Ue4W4WPn5RRFQ9EDWsm3SgFuCUk8CnPmUIFXDop8Y4DW1s
jrh4BMDewWHq6RoORZH7wvD0RqP0rGCntU3T/F7ec3VxbFpKDJO/NKPqtCWL+/ZF2UhFXlnjNPcI
XtL1H3vNuNQ01DVAmKTpb+fD9JD2ybqXRs9us5kHUJd+4yTOkC118Yh0jho8UC/dQBT2Wo01J0yr
DhEZRDZiBUiIge/+fD8D1LjEfKD+aXaMt3kROO4hFc1iPGLYopJHSHIZ2epYmWWKMKKs9ptwHLMQ
/4caq/9O1vtrm6nXQKxMEzEUK5dOjvcs03EZDBwr2u57RTmp3ffH9XP0xStyqN0EropX+SzrgILB
tCWTEYUMCYn6MNPzRqqdWvh5NXBoz9OyVFaCI7ARNX9W/+4aV4VWeRRQtGK3JkutKWnGXqpzT6Kn
ORt/0EoJHTU4hwxoqJGMUWQEzQznbD3SN+8oHdSbnotxKNuSoHcTxNj9wU7vwgwvdqjmmy09HHQF
8cif3wHX5kmJY2+ZRjEEhoNSAfh6176/teGNDoG/kTxQX5eThqb3nELszrRT6lu/WrIT1ive7CHX
EEULjbxhkOFiozNT2kZ1KZ9EIdqcEEsnJ2AVOZgwxaAimrsgHHH9du0tnytgOZ8y5QeEYKCUWi6p
YZXd/JtJLYw03kLAkX1P+9RcE0uvNibNTDrbZA+3vE+JygOwS59YX/m7vPAshXSV2jBrW4AS1tnz
dyHTueiud7eVGDxXDP8bGPR0xNkHq2j2hpHPP1or/JKj/nAE7gIJYPC+0BSSD6kydXOz1u8tzp5y
9FXg+y+45T/fJ5yKq7P3+rUL+4j3RA3tq1W4mjUMcVsEpuSuXOvEu570n1tQmYiKvst4IbhxMO+d
RoYBQ4g7y3PSkSX5Fi0zwq8OHR92LFlWzLBMjmJn+bbLgTaPEo/f1iblbTwVZJ/9B6Ufs82afMk7
Ruvbu/JPQk3zD0I1ocXi4q7oVi2EDUeGh0gaHD0qONBKGN8jgv7tGOWzKybvxKEI6lPiOLC/1dxt
NZr5MZS7EwOa0/28q88/XKAVyTIvhlbqcS9SLnsLFBykKpdsrPt7vStnzeAO1MKn8bt78L45kQsx
4xDoYQuxLqvubZHH6I50MICSrYmSuCtO2fNeO/VsveEIBIzN97aaRB70QNYjAE5YGRCIk9jN1ZFS
3Y/1BUW1hrwtrE4AiByEYJ16jzGmyIY6J/leC9G9wK/lH6cXlsuMZRGIuBS3mL6NQAo7efDkQiVi
LcX4wTN5sU81EsbGBH6DdeQnT3rwfRgx/pWmrYNkJEMarVEhYLqgkaY895cw4NxfxbnvIGEMR2Xg
9oAMrN1HwXuey79ErIwfSGsBayVU8HuvcmSst0Neumvu2wtoEETAlpoLYeIrUKQkXNM+b6ke6R0u
iS0NuFGh1l4dSq6qZaO+TCLz0yxk48qZ77dhQNLr4KkQvLBEUQdRx5dcolMWXHJi3ITepDEadCom
AQC8+eF+0G/B9/bN6X5Xt6AmEU1t1gF+Tfpg3Nhg+UVKF1pXECZl0E3qrXvwejSOHiZX/D7zUJHO
QCSudOUuJvsuX9Q/pwbiz9QIFfLi6HAtB1JGITthKL0ObCZE3xFhewwwYgl/9J4tDfahhHR3W6DI
aFOwn9BFUP2xbFJIa2OGQIq+/8tpu6fayxXdz3lSXEeILKlQOFfZX0IwwdUz2ZeoB2EysEq0DYap
mGGL0lI/kxkeoZzybv++JvKkx5kP5JeL7BZXqHbpp5l+SI7Br1lI4WAgqHnNoDum2g1UYw7p7BEF
K48rMrue+ygpVh3oz3dTgQIdpnwjJp9+NKI5wRaqxpS3FTIJhAkV5CLlUfvMofeUIknmX9M20GAR
1I9c+3j2JGs3+3JKG1Ko0/AiskFSr/wGn6EkiR1r6LToTofgR97xKiqjBMiP42v+4z7kqlEeNyHC
ZbkBmpeHFUAKrfyJ4BWH5BTW1eM9FuGRG3bWxgdxEMfH5xIEmprhvSVZ9bMJItr7BsnZShz056QT
za73ZCz409hdPM493kVbDA/Lh0XTwmDfXScC7NaJOdWGU4RoxcDuEmED49y+3RW/Ur8GEW3k+z86
BMa0nB3K9DBQYCXoNh1b68dWKSCweNUqi+ebsqvZ4gzK7AH9/uGf5PCiHklJVnAFj+GO8v4TTjUq
V9wvuMNiQGcp4bQdrfYmvUEA2dbkMu/UmYAojnSnJAHJGQlnk3a94zks/9iJuSFwBZ8SzBVXVgga
iCF1eVlV5B+qCqStlEqgxRR7bpqNV8/7TYD9AgyT5K3c2H0XRVNVMnpZBqUI8plZlHtOtG64KB1u
kiRpxgu3IF9H2ZSKIBoL5KcUx/Zv0rMp3WNbEhRexp8INg+jYHrQzAmRXteiGdC3DGtUeBlNySUo
2/aXS7ZLi2TqppXA/GulV2oZnKiBf64aLYikGvu0wWsLqt8wTIcgY75nmhA/DgaRH+/XpCOnLMLc
jpBL6VPEg3RydaGqEI0u0C5y1hVINWzAInB8u4bai542em5SnR1f6s3UXxHoCG9iyydCUFYOPHZZ
91wRTt9oox3AuyCQMh0K8z19KpA/7B8IXFR4VZJh9Ff5scWsijUpSprS2TyvnAXUCmi4rIFQnbkF
8KACEd5xnTDIqV4ptDu/N/hkPzFW8UI0bnMr4WdE3+82OwvxwhnQJVOzdTAu6ZKUrzhyL0GGnAEY
zkV3jYk4lbkQwFWi8uiUR6IRZOZQ59LZyLoFxc31k/9AoFpe66JhS6MpgIyT3syTjCWDnEi8dnvG
e/R+GkdbnqxRCmjk8spH51o3yzBlfzWxuhezwZDc6zoEEsY4oiv4YZQaGNFTL5KEhKBOTFtwyMhT
3kdfqaclzMapGVpbHsYNRIrbzQbUAniJuY7HgC9B/bv9lFY703ETo1AehxYyY34k20EDlwXCx5BN
5OcLJ9UkSEnB4ba2sqdcrZ/0ygG+Chd5A2uvgttbb5CelIgcIHRsLm/Y1Z3HhDSqip49W8W5loRi
C3zC5BhiPdbPIXWONfrJq++yPSQHGpgLakl7Qdfx/aTGjPXwKssvHkWjVmRwV4W96GZE3SUQ0lqu
1cdOeMJ/70pl6hD5NoXJ1MEcZZcodU8aPkA19LeTzzSrsoidbYxi0eyPdBOhd8ituO8DHaQGMgzG
nz0z1CF/div+lbofW2YCMwdhSkiOthQfQ2eHRhMeGTVk1yvx18OJlr/K3SSmjTAK6HPHrnPhFpMn
dXcCtBam0M9B5e+sHtlB+pjHbIS9Pa/3A8wveixHey9Aimv8RFSyRVGRP1jZTm7Ct4M538dBG9O8
ydibkMkUCnXG6ieILxTLkkVD3w1pjlIOL3ZNWSk6jvEny8opqpxl091UfibzUv4TkVnl7xJdR7/u
CO9KFoB/MyJopLk8FhgEJDowriLr53JEKGGjNl8dixVOdsjmyrO5XazaPdJf19PRIuJBxOB0Cbtt
VSsEbrE3l1nOEVvVBXQ1OuCW8ggOyidT92L2y5Nd6KHumSNfUy+/1mMolPWNfaP9ZwApsFOb4xCG
eNRbFvjDUTSLp6wO3yP0yFufci0SfSioDrFZkMchTfA9jnAdtuzakaItLxb4w8Zcpx41aEWPKt+x
FFviRc//8dhjTVBBDrdCOpu+TNut9hV8QZBWJYhY+rSKMady+hGjIlGi+vURbSukdPMbk1N+zSBJ
1rK7J2bSToD6ZThUxzzjcMHEq+FRzMBHKZk5VM9Xkuto7bbKvfMrVH2rWZASCGbdk8J9FGGHFv0S
sNHOa1EfVq5v6Fq0p5kmRQRbKTXTpwihyWDBepSWgHaJe1hhJs9kLZ5v2Lg4ZKoDACkwlf4PujGE
JnM3YMXmeGwCUi/7+wHqnrXYiDlzJEXGITVws3VjN3bbSlbapjBWYWOa8mzRv/NVtAQfQsMZL0p0
Slk+5U4mCgCcApUuS3ke+MCYbYcS+1y+rMx7djGI9Q0GPw8ypcpYuTwkBC2CXzRjTnjiKYI4Tnf6
LereZvIOQHq4hQqR+Eg531SMiYQfj5uS1j+o/Jv4UF/UOoJTrmQ90G7Ndq7J49eQBaNW/LJMCaPs
x9OnWUUz7mSB77DY05HkwGxgUb/rBCVO1XhBZ3WSPs5p9VNxgGxX8pyvj11vK7y1mou2PDsm0xiJ
Mbc3ConNVFd9/eCvbaAn46nsBJIfI8jgIf0mIQzYCyATXncsUukTzHB4aUPWmA3WgFv4wZZdIpR8
PSyYuse1JwGILXcCroyVv6Pqyv4x00N0Hr2LbNp2ZyHtgIjWEZHpl8P4hV+qyZf/kxAFQ0/kbioH
KXLu+HZTJkoYTh/b8O9ykt75tkAuEPy58LQGuzzl0qOyHSPve+pBlwUSN5fQXIK80D280gjX2e2i
fytly1jfBK7VVVwb4WpmLGFV1ThXecuqzzHxWizf23FTPRIC4BXafcscndmViuLG6CoQOjZK8GW4
SBpzhpr5GoAw21lKYxLCAI30EvFDQGOHCuK6g9/Mz5+8mjqch4QIzLpR1ifOiRkiMwOXC+ylkdpk
9pLc30tm8tPla8uO86wJCXtizJsr0RTNJmHngu1F/chHDpbh8kuT58FayTOblHR8zPwKAHEbwNNv
ytRJwVypBM+/k8lhDe+aBtgm58WeA3DWQ2DUEyYTczP9oP30USro9mJlZI72K6290325Ki+jtKRm
1WKf1D1z2NHVR4CSewfc0tbqPSMp9zuRK0DI6gVpuMo9yo2eXXxcc8tJBg8lKxfnIaa7AK7DjV0r
RU/t8vU8gYiRK8ZTBavCosYS08H99jhMT5jg+0YJ5RVKiJB0vWNYhw8/WFUPOhYU68eM3oKHRglH
IODd8rBWxLQ6jTcGGKrN5B4/WaKP5qfdegyzvJtN+lwJw4hLIXPDS+Tu+/KDWUqFMyTbU75jehHm
z9r47O/Rv/X937YW7aTbkEXRqHQ7QjX7nSVPD6UOWv+b8tdaPEVIb1YtAEU7VJL+MEUS09j96AOZ
xAX73M/g0+51OyXRx9bivwrAYuTFiRb+J0Jg0DYidKu6W9Cd62R4tWYZbOWQ/IEvp/3KmQiHACXT
a3n69SyXI5ivkL7OntQ2vU3g80fwVwJbGwDm2InArYW7sVP1erU5nJZGolx6yGCajmHnAU20x45g
j5D1CNHw4D0NRhKuKlXuc/8yCc1tjEd0tQGUgh/2EWMVvExNA54GRgeYv984uuGWiDs9aP/yuyjL
PsK8tKtdXmigia8p1KGM4QQ+d5wecgvraOfFgOp1IQib+Vg5oPYcHEzybA6siPqsFDeDl4SrzND0
0/lvFbXpTe7yjLAzlQI5Nm9qzDB7ltQepQrAMUTt/+/Ac+0Tt3iyeZKWE5zsUgUfI0lEW+MPbdm/
fZ2hhoPxMg7gfVaPnm7tq0I3bjKKUSsjcqREpk+LG+1JcPVYW6rMSDCoyhYj8nWIT7zFDzDmEtt1
YNTcPqUEeRtRsZ9LUD77jGbTek/UaJrOGQO09/08PpEb6T0HCsfnSM+puhR3ejylB/qXmfaV4Fxg
vyYbBSNc7D3ECoIUma4zO4xlvRZ8SwVcn1Op0jvZb69u+yXjBTi5cl9UkoT7gmWuwpyhBohIRG2V
WfCW2ShoTrR8yThPEotsYXdzhYDGSNTf45pptAj6WF9QGAcSNsFNDVBBoYP7miVrzfyDS4kXED6G
TTP9etl4ApyVkNznwwiy3t+FKdq2nI5glGAmG4WbSlwm26j3910lfiJ0+nPUHsoyZD6ZETs0hKWe
3lpbxkT88J8N3YJLkZqa7/dZuO/a0Ivp3iH5f/9WiGodepmCqo6QQ5fquEPDycB4spzhEHxfZ0AA
dxnsGMJD4g+6eWQNG7almVfkBsIt823b2SKARzwYklpIGoui2b0GqjKe9qsdhSj0uiCnkHOCzOYC
Mv0tVLX3BvY7c95wuHEY4wcvo2S3fEUvKXAH9Y6zTbZTp3gE5zFZt4R8jS8HXybKgR4TTrt7azHh
GSRJYOh8CF2W2U+qtF9MzkLoiRIKn01Qf37YJ9L9yQYgJ8mc5LFuhhcfOCKQjFXdi0VXnZt2eOE4
sELJ9qYIDO/AQgWQgTXEnkHrP2CYYKLPdLGJDbvHOYudCSA4DTbRUluC6xnW/IlXengOTA+vyYdD
IPQlgF++Yi9f/0pL+y1CcIc3eoxGESbEn4mT60VxyvyeB4akjl2dbC5CrsHJ+FH+x1FboJfz3dKF
ekcyU5oxTdwfeigA0oOzMjxd6cNy418K+sVb7+vuUWO2Xd43qFf7GSCDns+y+X6bL9dafuM6el/9
rjOFVf961D/RfENeljZT4yBet3gpwiNImQ7zWbGTMuqI7acchgGcfuzf+aM/GpLjNCFuQUYunNGU
npjOQBG83BvpLfOMdnKVRH0q7dhqbIMqzntCm8UnOKklodyJDLMXq8jZ6ecwyGNgQ3WCC0Es6WbO
+bQyaqEjYdSh4DRwRNkkcLbpAnHTovwOfCeghNjL02BnhHTAquWM69zjyKKrmhTNAw84TShHgWR5
vwyLKSgPCGYDarhCuvyloCBeAYgquLSEF1VZTad4lUWL00IYV6463LFNtqISWrSOSwnMdEKBgicS
ly+kjlN8mlBdgbNf5ecDrRz9c34DsosLlNW4nQi2mMPXO0GRJSE4zLi8OkMpj9JdC/WtZTUfl8qg
V7s8pUqmPme7Vvnac1kWGzooNSI+58r/4LWmw93uhns8UHOb3nLql2ok1Eg8lu5Xr2t2/Xa5ku3n
tUBZujkq5ARkpyjyjQ0e7VwSQjq0u0Y/pRJyIdq7bUCU2uvJz3hfz1X8dg6uykbe25FcrS3OvsK8
/GiHiN+k5zEN5mXX8+AqDtEF3CfsHDiDoZpMdkPeekAvoNsd5KQDzPJd8LaRA2BUSVa2K7ZDsGMs
hrKVJ5KXzFmYgDGJF97BKhvB8t6LEgAFl/lU///H5hTtKWdee8s1NGVPZbqW5KSYtL0k1VU8OdcY
/6NSrG7tx3k5sHaYHkquuXuTJ0zo8NyNXlIFgygF+FkcVubc1Uafm78JDbRYEIOE7X9SwYnYosN7
Yd1+MSIqga8zU6VvBCyugfiCFcVzqoiFoc4EUiBQzCgoI666kE1Jkxh/5znUH6aDg0y/Y7ZGGDz4
FU09ErCeKc276xx2ZML/6DhfkBa3PTFi14UBtaPt5eDZAdhSFsgBrmolBuHbFnCu7KcrV4lBk6g1
1nMYHGeCSx//Drf1DmIczk53h+zHf2AqpmxZYmGQzAV2FV87GUWDwcZkzYtVAPmwyQTtGTV9rj79
+3r4hnNQlfH6XvcqKilHDp+T+/s8Peh4tYM2qOHFjFhJfOU/c9TvXs6yCNWARj3tBFa8vmNlMPQ+
CRwvKAssE7X3alGyAV2L5sJ3do/DB5ODiD84bjqP+h2zJhna82oHQqRzwzbbCeVQmyskm8X2Q/vI
d0Ujydq8oKjaiC91JDBk5cK6i4654A5B6og2lpeMgq4kVy4cIcVNYPZBAora+40Vz4WgRw0keu7T
PczosB0IYtmAThjnR5bP6OChnO2R9LHA6W9KkgtzMhLFBK/3TSKEnrrqoP9RstF9sSYKU7EMKw+o
2deMMustUOPEo7yzDq3rkORKrwt1OaPA3p2wLgkmKDOFYYIRvNfPALK2BO3p+P+6VrVPwOWA9RFd
I58sF8e4+bLX5DJwdfwy92lyEK175/r/kiiMgHCZG8yzmTZaCVWGM3WIC7WaR/7o4bTahGYA+EmG
2Uqjr5VbVXMa7Vrl5SxczvpmUkobJ6g8CenPRNjDh5STWEhU5uf3ceBMQ1ySjgHDzDhQPaIycLYW
+8mQFwKjQI0LQTKhYoAR/fDHCMmokN1mq8OeFzXVVKxUbD2+u8/dVmbBD9yeA6OBYVErxOe2DX32
JjKc4gkVPNdpY3NSH/78zJ9VEGldSQF8rqyS7RdEcCMxML7jdl2hXTnvN7Q55DIOOqHXooYbzoK4
wRyJmHVR0C9E7l9jR3FZB4WIOSTG02EL/C2gZF0WquDspZzckUoqqdTpyxH0EbauIYtc9VEfDcid
cMUeLdtfxqVV074DaSOHUyxnZUoPcSlsQFMtzhHiP0l4uvEtcj66oB5y5MzVyS79YsToShqpRsCm
0aUjOxGDWy6uwApT5PbKfOIulWa839BNu2H4TioXakyarXzgZy+6nLwUJurv9R3EUsskMkZBZp7t
Ubipn0QFfbaUYshYaPdmInCHwqogogu1NJAanIA/OTkBw+nh+LoHQfmWjfKjkOlHwXTPFeqW2fPA
p4U57m6esQgKXzsicXzmG7Mkx1LPSiOFNLrBsnwNX4gSqOkNhq15Hay5HCpzytnxbYZn6GYsIpgV
2EC1yaGEEBHXXoo9qQCtC87gwRgYFExo+VEreHYWcWEGtdhMBH4dYJBlE3RP2F0b/1K9yTDcNUlH
789/mnON2m1fEg3mkIo6jmE/dvuHeM5x8jwWUpOK19zaGpxOO2g/4qlrp6LVZmHyHdMJHDmbhsQJ
14rNlluNIPjj5xKZkrJQhVdRDlPoLSJPCeYiEv4CPulRD7lB74FPyxO+JtN7MvbF//hs/6a3NCMe
52TjFH2UmnnpvNclxWq+6dXycBtASXbJ2EAuSPOhGM2tt0jyprmU/zEfZydpXIQzEF9xGCsbgz1l
EPNLSqRn6rSAXaKbbWD5BDaS6ftVhRuyrpJfRzmtxlkibl8XxEcQfTW2HW1/3008/TJPGSu17ICj
scUA+wIxatFo7s/ZpuBYsrw3xCKweQzYXH8+4urtttxZiHBfHWcCB9Zmd2ThEwIgIwi80yrIxSmB
LLkUCRzK7P4xdPc990dzRxJteV139dbh8FC68h4ID+q5264hOQQ7II5ar76oHfgeS81Ix27qhcbr
39wLn37AZwObMuAnnjDx8kLsGuAl7j+TNqq29e/xUfa2aHJ3gEDLqH5DMeJHCzSD2gOBrK08tB4U
RQjZgmjE2JRqEz1mfateKVG7PymGjWYha+ykTKUpkJGbuMZNJBYCwKb6RB/uvSYQllIT9mGn3Co4
EyQK70QwrZJQzpJbgWZN5CPiheGwxDvG7W4bgit6g6KH5EPb+K4nyi7jx6xMJahZd2v3hbgo2p48
J7acj/cWxyRBVazy9fyIuWfiIBCMY8fKE5Qpnin2YeUoR9fIZ6GBxpTarnwcg4jeRDClY4XUeqXl
c+Q1T91/Znzke0Bjb+m6dCLWA0hXCEYzFMTf1DU8ohUmkIrbRALm2nQdliQjrrqvDSZAtKVJ9kUW
V8iLiD9erts5FnWnGas2OKHI5z+in9izajHr32x1j6O223CB0yUgif/8PXjgvQXKIi74UJ/tZAsc
iH37QSeAnMGTrCwDnF7HUupIvvaYF3oWzy96ROl4ymeucOwGkmNOJP5F0pNxkKSBzp+LYGclyRcp
MjfEX8Oq7fQgYWAE7cc9le2PqfhI8n/g1X8gchtcihRjng41DlrtkeY0VnGGeWjkhyhWR8q/YASW
HaHUP2sWZq2u6yDC3kqx+2t2G6ogcj0RAplePoYCoSm+YoiOIj2b4iHU7Gh2GBIZUd8/+zt1O/C/
iUTDky93zGiBTgAPouJw5Cbx7QlXLsAENv19THhsRSeIv/LQH/TL60CRlgVcH7J7RfAeQx5b9ATc
VDrtDNN4P59uobERJx/HdlbyB7do1FjTB2Bb1rF7nF+aOA6fuD4SZhK323DN2TlaDgnlMhcLLZCS
stSiGZcsDj/7txtBm3jMCFCh5nBe3qXDbM2cDYrr0cvtLxHlnNEs4FPcPGmocLNeuwLl7k4N4W7T
/shcdeV6GeglN7rfC2qS7TJAH+ALtxIpRqxHEeYmd/Y5SsuKG4FmbsbyVJvizq39heoH0Av/eSLM
7XMQWwIKw/5tjMOruDJ2eTVVHjviqFINxo9+zWe5RzMX1YqpEBVE9vskmWrELxgFytWddhctPac2
q2EKvyzkibj2xYio7Dz5AfMJ3Fpwp1o29f2JpAddtzxzcJWM2sVz0F7PR94a2iSa9b8HiifAl0g3
ycvbc5jVVVEb9Wavx5yKcEgUM7Gxv1XrKsVLQZpkZ0NBCZeq/W6yypEjjCdEAVzGaYUSLqnE7FKA
MN9ldRUQkMo7CfZ9y58WqYtnGeejI5xPIX/vUKmMtPSKpkYfEJzhlhJ4YnKp+9dnvoz9NGJBIyhC
k2xghMxSW2vbZr1G9ilfSEoy8ec+3huo7MGtcwJaSWhaw7VuVKpcOix4iHDeMVAsyusoAtW7cR7K
ayqPPZ9FdQSOYOA3gArnKbP6edWaMxHvdDo07CnLADLeB+gQXjxFjcHFTh5kLV+43uXJ2IsEXqva
33ThAzNX8iWfiDuJSjxkkXQ9fC03pe1FNU6K06c40pAPep6ZtPTOTnDQOggWmvG/HlwQTHJVLdz3
HhcopxEc5uBxVlJNZ7JcPhDTPMm9u0t8PGJJ4QRGTF8htlptEI1UNMnWemQJHV8Wv5ZiITuved35
BqIjtbMZixiDu8qP+xnuHq9FAqNUPX00X8tV+SxVb0p1YlH5obNnjJyzLdXl1PzGgxQznU+UD53Z
d6osBKLF/n0fLnmWrm+WUc38a2fdjDnCNW/ImqUe/qrZJltJ6Sad4eLH7vg8aQ/r0FnS1vKzKRXR
0jQbrbeVDLEMt0eoD7ppx/nfVxgXnP5RL9jpcxaRJ8q8WFD0aivNZyMH0ea8F8ygHuckG+thgdDW
D7pqX7nzf8D6JTIFlkqjZGyQ90HII+c6Gh8TUoGVbBAyGEin/lxpyTr1ydYRO2W+Aoq16zatFGhz
CFxeLY1Nn/WVsS6ISEtWVKwHa66MylNaSGYhqWYTHpV4kQs4VI01DrKI5iJzbutx+bOvbOmhDnah
LA7MC/U8M9Q78vEQ8/xLtQykThw0yze3H24sgt5oY5OiRoo9FkX+yy5JK80jTZDXP3tz832befNl
8PQH3RISctPwTrchFt8rAU8XKW/Ijl0AZuIkMw2Nf2jIkloKxkDMppWf5wkjA2LtC55qMhhLgbSd
HvmsSAxQ+BiDdVUlvU2lRZ8AAh4ff80TFikFjU+kl5xAxLhXDz1+pFI4B9mL46VPdk54ASuXd1yj
d6RDaNn66yTHI8sRhDnbaRbHQb/WjxFQTz2sABiwdtF4cx3cjMqM97qBsibvjbRlfP5ZU+82DCvc
NVC37k/awmzQtHvxVwIcYHqy4ggWvXqN5TFwz+eImF/K5ax9DsmKlBhWQo5pzrcIRXP7QBCnScr6
LPekxe/cBwgcXIvW6PMX55rfRFU5tE1kwpiCTOssNB66ZVSBRvhDfd6JNzdMKPAPhgJpxJA3NZci
4fzTDoTlzva/XRJqG2mV03DJbw7Y7OO78IbJ6bv0oCTD7XhhXfIXPDcDpWqr92OkSRSzMDPoV2GC
pnBNBS92XvNBg4ba5LjztJ6tJpyt1GoXF8WDmDL+7X/AYQjrLTvq7BW8+PHoCDR8FmJlKKK22l8X
gBIPJLNrBNXuIPX7Bv000APSxDSp8ugkoS96uqd7J057m+XYQM3vGXX8zDALNSWVNIOpKMA2/spG
QxEs53LfqeLHAIchiYSmF3CsQ74QZTC6wTZmTFfucQTYsu0faVRpVYEDI36UQeGYu7O3pMARgma7
r86nSThragFZnhteB31y4wSo/aB22Ms4EpsaoC6meFXmri+XtEU2xIwmaUhdIX/BYl2lZ4u//RBo
aWJbcjhISxgg1FztN2zfb9HeMmkr+i9DATV+d/+RLjnsCY6C2uU6YydkcNndvnwqBLok31VZi40M
XI4pQTSYFbFwVVIS4kl7NtUi9GvG6KcV0hu4i8k87A4qDp34OcOSkr1Vcx0i8GKNHwym0aHGg1Dp
9QKF6L8POj0PH0v4iuX2KOgIWBBHB0OLtsS7u4MB76VhREPBPYiDIZ8GvqwSlX7wX2tpFMheQt1A
VKsE+wzxMbfevijl5//oEZGEOVF/cpK7LFed50bPX46XXZxZIe1+Le4bsn6wPwB/T6U3YcwY6MtC
4EcO+2eqhjsSVqdyaefv1Uz8eHq2fbbRtSOqi4W1AMm7StgmSjILBIb3loBfmP2/dR5w6N8vFwc1
qCHGclV0qE6Oznh5enX4FypI4IOHXe5CZan/sMSXUIkVGJA/qgK6ky8rai9gYqFd0pRONAKgeIpd
3eTk9TsIfn5RA06g3VOojn3zeeLWr/HlS+LTIzJrOx0JlyX8upMWyaDixz/OpsXkhHzxV3D9LFCB
Mjd+ZEzJEhHpQRq4vn75JQ/9P6KFrU9rF5YhyDVye4+IfPC/dHaxV8haOviy1QDrYn8MOfyOGH1B
TtxSFQqiKPxd0XFZuBAy05GBpDJmCfld2wm28MPhEKLlY6MmFaYGqB04iM0SLxELykZ5HbhUPIXW
vdxn6GeYSZSZg0ld8rSUavct9VDLhBAPsX93wKxTTYUiQzLApFG1MRpDcFFneczIgMXqnVZuVY3O
zVjxpiqHCnhpMt+iRuLsu/KOd1l1y/3IyA2Up6GRUT910WvtUbilx0HQE1rbJufqitH4Y2jnU0xy
G4VDhw20EKgW4oG+eJ/KWj6PTFMbiXvEGRkUY5nbH62JS5xoJcHxGrkpKmbC03xQ+aw9aq9cBLjk
1DVpZeJNXcVsVxmbRwD2ntFIAUwviC1gd1nc1rhl//u1IhtiQt4sIUsYLqfqX8l1nxmkSZpj80lE
eG6okfiCzEv/Hi/f9ZOFfQClti7/ZJE4P3BT+8kf/L4Jyuwv7E+zYTh1uyO9Xd2CkNvFk63Pe8J9
uR8wrZzM5jnXABJ7tgQjdHRf1AZrtYVJLNruRhhhYAlL9gyQg075xK7B04ta4ohjYqgHPNQYYCLa
fvnjtt8m+745DkXRPn0uNLVFN5BH405hvBv9QhRj6g2wOLDfOAX9FU4+CU2nQmxeVGeE11hOYCcA
EjAPpzrwAxN6wn7cWMyaAy1Ae3wLtdxcfA8f7TeFEtXZu+GLvDyNq/64wHLoqhCNiLw5loY2JEN3
TD3ClnyaeJ/eFAaG41WC0oyPPQZkLo91oYwRmV2RVZ5bvxe2bXqaP0O3J9Ed+C04tZKu0A237qT4
EvQN7ZhPJ92yZ1rP7RfNxpcYkD1sO7M3wfnVRdKWXMVqfjYoFkCuncP92lHLqsOdk/ncjvDifDWe
6K952WaxACGPGC81nafr4jZjUJyU7gddWVPQnQEoptxTfl9KLn1W8dJUUM5dr9kZw5n16CXfgVJC
QeWQAODw/gIPjx0pUrD+1uYY8+3AMobxvfJwC53Zr1WuTEAb77TMwQD/MfgRfZCHoekrWq3fOQ36
LE8hNYl7CNJF3ufRqvgnumpzujuIMaHwWIhjHAt1gwBG4+Zk6wO9W61+2GnOit6YZMb3PTaCSLZ3
UKrCueepk5F+bz8UY1xty7UseyM46gMkmzA06ZGY5vPWE0R6XGsaU+Cr7n5E0UQeeVrLkCXGZzDa
x8LHDu2C5DwsYgoKIx7UH/GC9ARXN9//bCxNa2C6IvzuE/A59xtFmHkoA1yUK0qprINt0epOYEmX
ocNIvwPc5UgNfKjTIueQvp17xAo7o/cb1JhX9iCxS9E9QtgDFRJfGzCP7LptUgdzQcTACjiwR2AE
WCr98YLbPGGw8g1qMQVEbH4Agn8UuigV7hmWWF10+EWQlYyrp7UMuNr7920w93J558CsNe+UBTxc
50XdPiBX8zwCvhBOuQ+1pu8mLXkk6B/BcXwVjlQG1FfJcft5ZcsH6UviDYbYOOtE7rnejsuo+iPe
NcYHqCV1M0oqt4VLdvGMk1GjgINeR2/r+jEk2nl/6tic+bHIZd5zhu6WF3XMkcfun3ljTvtxacDK
kBnMyFzRhVJ8NVJV2864vzpAys5GFsW+K/YBLTVjL9CecE7TbHChfggn3BmjQKlijvVfEHx8IgUS
bCorVTxCEh3Av95uc3uUc3QLuDACqdavdCBTg8LjQA6IZ+ox6mQs5X8OtJXmES6cJUVOPYHmH7Io
2xk5JUDpEIJV/h+H8pjDi/TzThJZmsApBxYOfCOyG9xi4bpUsDLRVAM1lSwOHhcuoh+vA2Mjmzcu
1J2FAQwA8vCeu9jkV6eQFVYXqXfYr7SuvMLes4hV9Pq21w3me26Iu94pioBP3/kCFQHGgb9ibDmg
TTL3SGUv8oPqQ3mraL5MIbtaoGMBI5myk4yVOF5FSI24NQ5F8DsFQaPlJ0PC7KARaH5UROlNsgqc
x0uOx/QJsMLryUVXlym9RzYIDQnB0BRrXGz5R21e6NfEGmG828Rt7xIpzHGmf9lueqyhBKmfveJl
dIRaXIni7j0cfceRsVJS3zTCq8LhgUwgoBFtx7FtnDj5ubJU7XYK9c7bt6VyrYEjwMxpnClG0Nwu
FJuPjf7d7jt4rvITSN7aTAURv+AplCVNsLHwS+44EE750OY8gD3VCg2IqoE/y1xiOlSc9Gfsb9g6
mRwh8+zIlwQpP/pwuqNPNhJZf7yehepf0YZteqDVpnNVDOIcAs16swuwHGRcGhhAI9vg4CDXYIC2
CwOV7HT/CJjQ24p+zwRfF2+KeqLF/jgbAMKPnt9yCFSDTX9vMsvsXeT03pr1CdfEMxK17LUd2mzt
S8oR6BTwXM1Lx70FOzXf0zOlrzG/MPtY3OqLjstHcUYXkjYTOYtaJG+G8OTXoV/lamMMNg3YQ0BU
47o1ecj35JTKWhnkecz01R/9rwdj1nbvXl3eJ62Qhg/eKliLEGaiK/gBmQNQh5aQ9QroTbBb1cye
E46CJZ4apTxkLlK4tfYc6B3RVugdz0cl4G/LuyZA0eDwyhQeffOKokr4x+fRc2i2SUXXLrhTOld7
78OcLN/P+++qLxGK3b1XnXovTgkaaxPTXDKHyD8oloFvn8DIXhdt6pj8xhjX6iKSxy6hVedroowJ
j3BLkQ3Db08o5KKW/5BfOkeppWbH2AotZCk0Ol/BzLn27p4LiSZemXt4aToXzJB2I7ja9gqiTGPX
7IDjpcVHJnV0m7aHm1CLXjnpKDHLfwj2YcjnEl15U5+HnYAUJVC7NhAKVx+T7e+0v+NIkxvX64gV
I6yZoLauxSYaPjQ7C2u3QdY7/VZSwD2t14iV/7TvN6Zs2cAz1nDdjfqdiJFE3aLE9g5uku6JoqgV
ss1i7ueQ4UisRxVBX5NuKLwW/Otp+e994B9QRamP8tLo3nVTlf00TzLifdYY0Twl2nPV4J1gs6FH
ZGbOKsiSsr32jkQEzl97QimqB6lkF6L+OLRCXQq8nKXxtaqrEwKw6ubzhsLjVAmZG+jcP9agDG69
Vaz4BzibLZw2wFahAQ3OvFik4sYdPdWOmmmyCRK+sziyGOTD5LPvGfOYZs89wJZ6njVQnoiNmyHl
WKWQIz01VCQTD+qvqH5ImZNlOX6+0FNvebt2pGbCPW7OniIPQYoSEG25nWzvo51jkSvOUJwg8sY9
CpDokjWwXHyX+MXZOHVE3AHUtPF/QlwEF8yJh1Gbrgix1WKX3fLemXNZPWseA0ClO3r56fJo6Lxb
SWsFfYCXvUV4Ii1zqkcnxFcmZq6CEbSLvzpLWsxpnpGDOCS869vRgyfc+o4DfzIaF+b24qHdRXKJ
VT2I6TEcD+CwFC+4VfJY153PWeaHL9HvGHTCotfVWYWvQiP+d0Ad51Or4b19MuxVoSyoxyYf/lsc
eCHEcUPwXE4QMcvBCkeB+Lox5sxf/5uYhv58/PWA+2FhmpWckSoOAiEWIA6gg53Ej4t8uUk+i+GX
GCYgWL1WinfSqJ0TIRLvTqToK7lPq2eg6tAHTdGR2EvAWBpj0/T8HwdhwLoan6IOZC6u1mIMR/ha
MUuSyGKx/Hv0bZtMFmp3D21sxadgnz120AhqZsEQiIjJnSAed0soLzzmqkEa7ddc91ZE/wFZf1Yr
o9hPQOJzOL4o3YqmMfLhUrXkMBD1+AdULmzMqx9syrQHSz682AJAWveY2P+raWJuR8VixGr47DLC
HnkfONRpvGTqR5AWX/P/Oh9ep+3Id+6+Z53TlBnIXjmB6L7ihmMpimpY4kiiKvB9n0E0/9M7RqaR
UG3fVmR6L+g8B+cwdCYgxm+srSucJuuLiVbZHpsbKc5TKwhp/7ftbMwXUav/aCaVcwM3lIRD2nI0
YY2Eqx6gJ1BJxpRdPXRH7FsJqhhmidv4KOxgP270YU9CDpEnmMPvOXq8hC+AdSbkyT55vFB/GoNo
IqVTWIn/rjczGZPLp2KlkKgdS3jIg9+Ph8jeeWo0ErNZ6PoZd6n6TNk1Hgp/2snz04a1Ho7F0Jps
WyxNXkzmDfqi/BQAqHNz1lrwZHySbhkavbxUZgKxx+TqoHNwp9i2LHTyBpUPb1nf+bNmwT3KxhnT
12Sc6yqEbyr/DxSGJHcNznOdWTpjWEmnOXeEEI5d1z69WmqJ6sf/KAiHNkvHwLJWuY5o9tIkRiy+
hQ7g9+9AkZJ+khRjuftaxO1eiWEiaWOGjWxZixeijTbVxZGYpcueOAptXyJWCKOEQxp4CZjP/BBR
QimtGP05Tm9KwDmBv/gbx0262ecwOEXc7Gu8DRL79ghZXzIgD6qmW8JuespMvrzbCpTnXMdWcArd
6VuuSg3RfEHmp0iE7dHhcT4w1B8tGvbeAxcI1AQY6Anzes8MmdsbRVKU7aAn1lE170v0gnx7y91q
fp5mZRDGU3FpyprunW5XTwiLQzfheUP9EzcR268Ash9LYOWWzc2YtzAADcRMuQB47xFHbsFN8QBZ
mv7x8/MSSg+i5nuq9OPcAj67IOJ4CLrrWlRp91/ivVbQGhuspXNRALD28vLJm19//xScuymQETOI
CGb4GkBVLakKui8KyqJc7HzZEWhbW4a2J31xi0xBcPdsdJsS9cUmQHHydnrj1pxCVtg+WeX4afWD
HesMjIGCptKrhwfbuB8n1msOGZz6rJHJLfRkFH6Df6eaWvOZFZrGdgoG/Vgu7B1hqslzI9h9DQBQ
v3wxOMf8YDWR880CfzNUNMK0aQdztmB5tanG+qpwK7LBqXtKBAJmZMmlTgJyqRY0gP+VGNVLJZdg
Ky2HfmKo52kdTkdIYn0XxG2lcisyOYzUvkkJowDTka1X5vIX5NKde0ydhDl5cInNu3E4CnjoHoex
gGwUGBPf36PZhbjnNkB+c/jxg06LQofB6AovEHygm97kAO08It8o+tuwS340MmlPuU34kG9xxLsV
ZWIsI3jqxoHXRzpG5XIJPyHEfYWKGJgX5xrOukLtvQl9PVujrdXsuBqvjp9IQBzVz42H4NgdZsJS
5aE7stmf5z67KoV6O4Bnf/bTn7b4G8xFJGFEq0+Oye+WsivrCCReCAdXJpuZsnGXZupo5pgAoiO8
xNP1iaLj0FAT94WO8FfP1rebQkPfY832Sya1zGTnXNXCCAdmlWnzrrO7Meegh9V8xkF5S6OsSS/Y
83DEOh6X3nkN+xLCe2+ON12hmpSB6z0vlzjXO5cdGqpToCcRazAOJ0TMewzuScNtbXcFOo/MAP1P
TPDbew0qTuz4aJG1o+9I/FZjAkO3QYlKKwQSnnRDn5W2A0Qp6jJbn/QVaYq5vnvH6ymn19aialUz
Ir+bLgrebvJ+kVtUohw6S7pQ/lsdvezPNMIFtzgslZEUjPokGEtDNjWOtpKJt5a/qGpNvus3xK5l
bfAabKoUmk/SePYD6UmJm7Mw/iqUx0bjjR76oUxK0erNSvOsUVSfMTwenE4onX82+XmXf5B1nZSn
jBCiPwV+AbrpogNZflGgsM7vJJlg7vDV73tdGHQ0/TNt4iSGzq8dz35H6Q3r991aUOJSO7S0TWfr
TRmHoXCh1bjrFVjiCogtumAqnYmv97SQGIXyEZ+D/+StWF+1VZxqiw1eGs5F39J/gitb8RJ0Vr8r
d26tigB83cOAUTiZSkkmZaRvkv/I+h75gRVxUuPnnpTrvGm/3uJRWp3iKRLEXrEz0+eiaB/xye8x
SwE0tT+y+HHz/Widv3Y+MJQQJhKnBiunKAWJG4RZYxvh7iLrQUJgreMRVSRh/MZk9mAV3nW3guqI
4bcL93e/MlzegW8V22mHlnHumuZ/AhBgikMudeVAhcEse4AXy1CQ+3fBW8C+ZZr0OMveMOVMMHBg
KQ43+esQqvxcIlBADztXy2JoAnE87wX6jJ2htPwC1MO3Boa0udb14TzeLvn4mUEz0VPLVDPWBQfB
IgJ5HcsQjkvwT8xF31gHKz9Ph8wmhzbtJ+NTPwKklPaI0IeoYmyInE6YCJJj0caR8fXfQLvj7fdo
l768R1PdRgUppOUnggwVf2veZmtxFiAWmJhUjZDaugBGGdIjBLvJyQ9pUnljev/Kf+IiweYdzcok
Ejdudjxt+SFeS8g=
`protect end_protected

