

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bdlZLEAewQqpv1o7OoBr4R377V8Hk5Fd8+q/Az6G9nxroFaOnD3V9+lWQZaiTQ+UR8tYlBixiDT3
2rrbvlUYqg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PNj5XhRRPylbuLUnq16m36512+Iu+tuxUNOB5vui/U9Vyxliy5LDYUjGyTrkosJ5RLmSfgYfmdaq
x3GXyG6MVOiZo15XiDmGz5Xa3WMM3TuUhfpzNItvR+cjVJcfSX1Vpo9/m4Gf2HbgWDY8/uge9Yz+
pdDWTg9IqOS1f9m0bhc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tfy6e9ewB1av8IAVBQg5F0wJVpezM47U5T38niEmKqoHE2EAQIsVtLXdGuC0EVCv8iR27vcg17Oa
mBfBXWB60tzPu8Q6DSJi1RmV8OgW+NgUvCiTMpLKqqsw6FnhMEK3lQVXfOtnfyh9msybPw9byzXC
dambJMmCpKtH2TBazWP4yb5ww1Nsz/1jL5i1zPiiJqwiUek+yJBHinlLsKOdmxiEOjEIxiuXMNyg
LMJzb839xkVhlMYTWXZYlSQVwwm/sLGnZ2Znntlf9sYBoE6D2vYri/PUGcfI5TqvvhrwG3MMHoTN
rPYZvU5TTqkZ0UHzprP9ZbAAvBMMlhHGjyKLgw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
enscaK3Um9KpWwQm1hA2XwO16XJLOAeYZ3URNnasJSAORmdXiuv1QgNvxstTqRmJdf6aiVcX+SBW
QAS4XOQmaHblVVCTrTFxq+i8/M/uWIiPlKdwfgcbq6W9GDVZEH2g71B4sNE7sbY88daOW+dsFMn8
evKdCCrOhrfApxD2w7E=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qn8TdDpu0TmAhfXr6OjdWoz6rfyBW7fFZKyqPOjjqWteCvm3OM0JlharuS1oWtO6vCpto2FAzG/S
BlRFnD+qM3W558gotDG5xKLXH54U8vJ9P7HSKDrDRZfcvgzYnDlLOZYqIhF3QcOp7QlIfdgIFJFF
P1RDJ8d43uSYKR66QV0gPXuT19+tneyhi0YpcaupqD9/Z/vQdGHiorXfqzI+zmAX5/7dF89mvr3v
Pvp32AibqOZJekU7QCnp4VkIAFQi2sNR2R1SirejbeSwa+gfCdYZC/MT0OFTfQjM0uxBSK/I4IyT
gWZgfuPijqASxDrsrURmKezc4hgCDujIExBWaQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21952)
`protect data_block
llnDAmN3bKLhgsWzXK9ldDdHEucPtfdzvQ+IeQs2pP0c1IFTQG43FJTRifX5NC8YSff/HEhS6RB9
G8iKbLuMw/y+CzDxOxVqz4048h5om23nBdE2FgLmL5ZC7XziZYZXBDpc2R/vCFVD8Ktbi+vv8+Np
x0COHDW/bx5TjIUzqdcapGN/91xfmbUc5XXXx+kseGK19ZLUBrczlUBlCEuVylYAmrUS+TpwJ27/
5a9uWYNc4798uUKwybi8w9Lv08xJ2AQkm2nf1TVPoQYAiLfK5W0wgCz5qUQymdjQDpkfxUpYZPIx
Ca4VOY1d3IlMN0l/sqj4hDAyPg8L2yOzLuAMWeEPOGeiJo4t0vFUDZZ/V5Lb4QSFdtXjPn0hxyI9
c5YSrCEbVyUOhLc2IBePxpgEAlqYAM5yJOPBJszLpMRrXXXBB1yTfJYVosV1qYlYsIyPvqAR0lSf
+9v19aSJfSfBb5yOVZMyjQ5GW6u8Wtf/nxt+6KCxNEpKAR0cBE7ua046JFmFcTeGUlxihzP0u4d0
UzkWW4D72L0o0jpgBF0p1/TDlPegFZ0vQEIs+uzrXcjKl/ua8H8aCtQpXolPV2ru5/KSSMMzFYUG
YZu/lVgXN/IpWry755UzuuI54B1NDsL9CbI7JTQjFlS75/yXvH5+lxKSj78wvH2E4J7DPrDc2DX3
I031WvqDY9a/xH1Ho+qa7PPaCcsBOPrAst9ce4KzwtyD2KvL7Nuu9F2j3w47V0g/m34QHW3I98Sw
Ve4d47gKc7fdC57UCsZwE7QK6rYhlEvJld7Az3XmfM9okY65BOPkaECRzY0036xgIOKgDIJtVTPI
N9Nhp6+CfwfU1/M+0zp8PsDrc2XAM1yLSggqRHLKzajHPVG4ubGFUfq6JIE5zyOxYnA+dPjZRWTc
X8s7LPEJD1ybhsR52bK0hDSHePYlqwHiy7A8z3leoFpiTqvTjI6HRazJjjg7jINIAE7oWWMF9feC
jtnfO848dUB8/RzFl5e0BMr7gK5J/2EBlE7Ee+s9e2y0H3hRXR50kkNHtQJ7XhGKTDuROHiQu3vN
nZnE9jFhVGPRsYO47CPBpbSa3y+ZJb1DsmeuiqlQWFip12cb3gVRecnaN3cApxJO0Q4VFLEfBiZn
XX/bppTXYapNMbMxlPNV+gNF6LcI6xlnedTP8V7QlH0gF3ln6NQL/YB69L3Z9XxkOeOAhdsYOYyn
+7p7+my3eDBlNLQzx5ceEdPyZDtG2PCkGYCYtfy0ZLywOrBHsWCG/zwXq7ghNeDT+tNrWeuBIio5
w0GsVsTZHuKF19eg5Lf7j4lM99E5nWJfPdlcEUq1APhGnFsjEsudaNwEjUB0Hhrhw3xJ0fVJgV6d
B9Y/RP5CTTtSQ1j7s2wiruDWmgts31ZQc3iQkVJVsD0ClwME9t/aHP7Pm7cL/bDZEm3c2dOqGpyc
yoVFMSh4kllsud7PWXoS+UKW3CVpIwMFssGqk31pVWjr5s6gxei4KqrE1ii/6stKkm+2TkKp5IvL
a4EBRJahARhzhtKnrEqEslOZ3qZe2XZx5YH6YUOKoDxangW/cNqspLss7/Ia6/BDGZKSXGYfYxyJ
T/anA2EXFSgpMCDv+nI4tWgW1HPO6576Guy7Px/ueSe1HmPIczgAXUz5mjc67oMnCzg6iaSLEXCR
wWUej90L8WsxN7R+ZrVN6iR6LKamWXr+kC5H6mK1U+P9MR8PptKQTAdqynjfRZhQRJBot4st4Z8w
E6eriPORVTbNPPDzFqbj2BOhjce5uw8DmkZe17U36AFHnTGnRQwGEFNAqaek+YvIaQ6NKGquEUUw
6LAE649I2E4oVl8TIoyZ//AeI6TxZju1ywGcETs5RW2jBeIBxU2TC0ZuJZEKZ99e3mijmfvv50hk
9vu1kERuGy/EX3wueTaUYHvFuRHFlCg0eoTKVbvQf4zgRxuMh0dsIeqcAKLUQ5g9Caw8ybJL8hgB
UbvycZyGjJSYCWK4WlgZmF0E9vBoId1IWnYk/YWdRo0gAe8V7+7J48uyvJzYadZ5sIaOSA70J1PB
2BWjyLFSBSBtG9JbakgG6FUb+tRuuM39LNcaRyvYuR0BQMmfecCuyapg+mOP6DwGpCBLerDxx0UO
apbtt9IzelhLVqgg5PtTlC2ZXLoOotUOPo/S1lODPug9cD48ZPB3GRC8NnvWKRBQMpQaXDUWGXtb
Tte0Pn7XH8QAgC0sevvfjt2p29ZUNns0EXyKdlokc9Uqbig2H1DkJXEoZCbmBmQpbDFNtLI4hzs/
k4VOMkxPnLag+Zvt2FsPP74M+3KQd79BoBm71saF02LEbTJOWMihS9Dc79DBV/VW8ilANjuXfitk
zDVS/s+v8p4Trlb2ihofVMI1Brn8kBUFmSL4I3kPN5ZSOHgDo/AoNYcwr8hrL2dr8Amw7EtLFblx
/o8YIuKlQC6SDeAYRh0rgJLQju7sKsXsUhtJRpW9N16MGVpqZ60lxFLOfTtA1HJNYfBuTBH0NN0o
KLMeaOSZnO9yaH919yF+YWuD5Jd75Thx+RJnqpBu5HJdlxdO8rrnqTkmBJ2qWiE5MpFfixKYT1Eq
ypB/jJTZRXEqQYvUd3cjA5GH2i/o79k/ctg6nv6K62xyPZNH1tEiB/Iuueqbwz0cuzGwRk2XNb/Y
0UqwUU/LP4h989sdC8i8gvDSeR2qCeE4ygv9ekUigebVh3Vg001dWvDX/YXbMN1u+9xoGlf+q9PI
lWxHkAXgZ6RuoklQafJHDqWucYWGjqn559VFRoCUlvh3OEG5cjSkx0nY7WJELdlfJno5Akx7Wb6f
vMVttOcl/w8DpI2e9w68wpWlkXKGJQPeIdvkpbKbg84+zHKIH3ozYWcFmyEf5kDgiq7TojC6/BcG
OmOmczh6PLrHs9q/tEGIO/qSWOPbRzvDlBwwWIsMmeLFDtqIJNlKoEguaZXhC2TWmMsqL27SwoC7
YFC5N3LHIZWgxfYR8la2062pnt6HzNDfGFfGtM6DiYbt2jdE1mRDcHOOZ7o2aPWwiv6E5SArIhDR
63afGacB73t0JMZQOTPtndSQ0CLkc0YJFu//kbQIGqSvzugVXNdsaZfbamWppj0P/fuWFnVipWze
JT0YElZrktGs8c4g7JNTUVQhl1UpxzWcdvZl52NDCl0M6dxdhXVnpUt2hESXowjJYSzEKUH6Q6UL
y4ROgwCH/QIO3mdayuSTJ4K8jJY9/tqZhNW07685v81yvGs/Ed9Ic54/YU32t7JTd8/5wFxx8Hr3
EgXQLqgHsHqJJs+/ejF6xWsrAOW+JTaGBd34UmPV4fVigY3+ZVPyU4PFxEq8ABMq4sCw4Zo6Z4HG
vZCtPXRx4ekXjQxDd1gNX/QLdcoGbMdY89LNGpot8+B8/u9pLIyYu1hQFe8xOJ6sY+MCR/YH8F7r
3UiCTopdlZuRDUm36t37L0gd5fqkJJzLgRtCGVGvVanRM2PvCpaRz7u3tRYfWPpc0W/xLpV9AYhh
i+ceMCcw1s3mUzT/u3JlBcZzg9AYXKJsqHymEZvfWjhbyDOMog5AuOnu8mWUbQij/+Ns9opSxg4i
yyEnMgnqPXdrS8VIQIs5PT96rFHKxfnyCVtqgB60nYIaaAXKGe+nL7xjubmIDH6fT0+WE+JI8TOG
XDlCv7MCv8GBdJtyrVJhpS96j0hdCTs/JfAUpp2NoBTEBbRLKZHvqjbGIjCQXaDNxNag5jt4bF5P
Ou3FV6oNFr58+3xwzKLShicxaOGSlb9WPUYTzgLn0vAe0Y36WB6FK7EDVMZNKcduUV33lwrx7YEi
SQCP19PVEXufFY2LWHLh3L0k++dghaBbHcb/wdo0vNIh32HyzZ7+VgQKAhXO6buhlGNDfFohUzlN
GOeE1L9rOM+ojtfdy08JPFlKTQwGXEiDueaImqG6pslYhaSMFgw56b8wNdTMtDOBuDYpILLIk2tb
MgSMIVcaBf33aYLVMjlOpEnSRtfD/2nkmYA1EgCbV+S69UnK51x4h5/O+ONAKyv8wJVsO24KQ0x+
wA9ifoVhK8c2Kxq5pMI/FS1zmspk115gHsDRzthO0RO+BUtgMZKxV+PzWedR5EvGhcu6fSjfeiJc
mp8fleizB8La+VdcQmY/JaJziCUsQZ10uReLHLFTy5epNflRlFO9jt3d8+4tVj/UwfkTqhko9QXD
mV5ZQraTjsc5UvBAxpbLO86mWkR3KBchPvtKlgmjakyiP4ajjIN26I6dZcFuaunesjVCB6ny3EhJ
bzw1W8rX2ax6+olOA1GjvVXPttsig+IFr1rbhTdEnXJGWodb0Y8r6Jpi3qW7nTNd/5bokQhytgcu
Gz+Vk1T0sIygH5o04bDyD5Pm3RYQeMZ7d1xaEKVnVc0ive0ftbEz/3Atee1Lz4WImop6GjvIXTeF
EhSMXufRhHWOX5ghHunvCyiz6D3UV/E5W5YF/t9og05P1vQmeypAUSA36FfZ/9gv9ZUniX13Rczz
LXjbx0c3jb0Ea6bD7JiHmrGnPMC5zpEUTvIuvxHa+j99yMHXD/R9JIgr9DlTus0YnACY2+ZxUz9T
2KwAe7us4UIwKpmijre5pwH8c/Nt+smdIcCbN2niHfhHIKxDD6cjO7KON75EKHUDsjDtk39eRLeE
awvDfVWxC69R6qVNbiWFfGVy8xkFz/sIlOo28It8S3i68ZCqUC+NscJnzC2VI/Fv2sW+fo80/+cJ
rWrq3BIAiIotrDOWzMVDEyCjLiQuJLrhrTRFx1reHn7kcF4vNHAXCdJrtTI3j6Ux6JUNZRUEEGVp
DNZ1xvFB09v8yrQuXpTAx+XZxJHk8fPOqia8IBAnL+uAyE9e1wD5DZ4iL3Z5QSPRPS9vRKoUtsJA
M57AwgNRT5YuDlizBSyme60sp6FmSM9xWi5B6G+uF8yeV/hr9sPwwHS7aGql+4YUQkcq3RMKP0mz
9o0d9tYJSDz3YO+Ny2mEN2nUbHTGM0Rs9C3eBVZJJwnBaD/82/btBSNm/qlbjjXAtKMGj9D3xrn9
UyWEQ/Mh1Af5TbU5fL8U8TEFlyA3LhIXqSSVsTKpRmdr8nS1JHcIAduyUJ3f3mDiZI3KDjj6xYx8
edfcrGN3f7vf1PdpC0yVohrUtGufxghMI754jZ3pTdhoq8PF1ZS5bvLtvmu16oZ4lOCZSoPzQMJE
YpyNCLdC3QK0rLw2H7FGLwQDVY6zC7fj6B/vSgEhJlFu9wFZqp5TEEdOfk8PqvbmuxOXKOfnN/9I
EYu+c9qAWXS/vUJ1BNEnNbHRYYZ55mzL2FbxwGDTJ3qC3MINO7XMSZ0kmrou8OmCz7iSUeGtsKG2
ninwaMoOs7QAsmRDzmwWVjIAOBvXUDMkqpa9p/HR6NVK/jsbCuulyMLJEhASr30hj/alxndnevmL
j0nWXyS7BZbRjis58PwYvNoVy+71VKybxNQrWuR38lHrnZXsURSJrVNbRFAfwokiQ7OycMziTjRi
8mpzS2JBZFQuse8z4APtx03S0C080/QLBxg6a6UBgHxJlcCim8T9849wbI25uiwG4ta9nZTjImuy
GrTkcqaqyYuCHLOvhTSjbBxv09hgJB3bE6yBFDCD98MsmzxcJyRwkQnTisPhYVAfJvyfmoyQFZ5c
bQCTjSNO2N205Eu2m7oF/gsN3Bepfm0uFk5k+hZfv8PteyhdtztgcyXAi7PfbPSFHIdsT1Yy4j73
drl/fg414Kvk4BQ0m8WNywDD7+eNsvMfnb5Ub9B9v/dO94EWwfk5xj+vHsS6mXoHiYVm6XW4LAOt
6ij3ueUen9vg8LmyxOk6fzAKZ/LgAA2liTna6lmicLPr9hwRzy6Dcl9GGaAC6Fo6AEYGUeQqwj1t
eshTqd7De6JxcGo5z6rrpyhAlk7CK/9SEBxwC2hE53gsnpCZatPk7skiKERNdRjswYRMgeAmghCE
1q372Z2xwySyCbd50014hjzCUKxDg2y8hKrvCRVMEWyK5xXN51xLIbWlQHEkIEx1seOclAvXK9Rm
G3RYsmhnTENYodhAu2fAVHdFPPLQXlCH1TU4qUh5Kjpa+eYYE3CtCQCMuYxIqYP5ESp7515PrV5w
N2bHUD7DgPgOkEwo6d+jaa44u1nSqKijNULzdAXsIebvkVAZhdFfOeDSbWQrIvVtUVZRjGdyuwLE
z3KKyOBmkNNFvs/By7TuSYHW4yyAgWznHr+0MA+fNCWDmFE+HSgxtKIcjXyGLhTq8L0xnEi1WkfV
TYbrEOMSF6zn2X/T5Sh+Nx1Dkdi/gBea6Xlkie4y8bjWjEgl6dmQwuX1hXoTYojrmvDlh37lHExY
NlZIIK8+p6jI10LIyp1/LLmVHR1ttS7d05EYBs2kejQ61n0BG85PECv4UJv5orr7zoQmTMTMMwfA
l8XQtGJB2rkIisurtlLKHv8Tf4UtNugw86xBAIVGlMjn+8V4DSgYMkwhyliYGKoTeSU3oygMSQPJ
gJp2LwNSTEcIWWfXaLJ38n3pdRp5Ysmtbt4qH+BF+/2EVzwLJg6ob17UtRxlJggD8vMKK65xamQH
8tLGsA4bJf9H5Cv0YI1xHzw9/DrVBZB4XahOVV7YO23y/oHLEof5JYQaJQ4A/PhKQTiBoPTNL/mn
xPIG42UUZZV4SmLClL3++53zq/WQjAc/C7rhStVkzSMoG86VFWzZ48+QtLXVjsRV9cnJx0BnHC/H
3pTuMQbWV/FNtlGky14rkU6onqW/0yHKWYzbsktgpHFw4hXze0BcF6NAFBAMmzyZFFmMTz9q8rIO
aE22yhmSLw9ek76Rvol04+iGm45sMGH6YSxuHjN2SFNQjRyb9htPh3w+47Jz4HqxnpY4QZiVSVEY
gKuQ9v7SNbgWrWbLrD2R+/MPNFye3Bio5DR1xR1B5YfbinmD0qNFkc+YBw2AA8nr3+/CkCXZZ21Q
4NTsiyQPgXaE5ZHRJjqTIV7CMufB0O0ACxRmQBbdDr1UoJoA2gou0mY8jJzPazrj3zucKJySjJNf
az2OnnD0l+JV+7eC4D+AJjMew7zKi/7gUTp1GNUmCLXUjZne2GQ/u4XchDiywwXFtbrmmwbmmQei
IS5gL7adrUZVoV9Ykr+cHRMrlRLyauBAqXZ1NyfHd9+B5AZ/MpEPq6OsZCuaRMU6G2IPyKZoJFaV
VBJTwGA3pWbuzLCfN2JAEgiiZvk68bLhWUb64Kx5yqYaXCHJKP8AuUdvKJzbywByU6/4hw6Bf88z
6Dn5wf6qFm+TrDFkGOtze3avUKeD/iD/pBELomC1P+KzBhtWDPApOQ69EHRuuPfoAY7uiE38fUYD
OujWwGZg2FbnV/0ElV/F2xHiolEEdoA77m+hipq1Jh4uDOiTMp13dM41n+o1uyRZvRk+uoYYAQRu
xNNra6T9dQfJb3Q1JfSFmvdg9WR3khtsyIofuPFeOFdHEQ4SLBwYZAwpwZ9LJ/3tG2FNDdP0cwnp
egTkqBHawNZv5larLCmB+J99MfQvmfPdIpYqgr68zjuU1KTZ8307r4RQVGroM1Jg5b/aWjIEF9rJ
HaHZhgQaRovPvn0+xoFE7bQv8REkmftDbuLwroiHxrO4dGnfCLvZ1gkWW8ODQmKOCMDS9TSvYO/g
NEpea1Y3ZCkaqGn40R2x+Kvrr/3LU2vRyLAl+8W0/FT26PGYuunS163p9hyqO8vp+37XK+ZGkLac
xhku8tCDHAtQaVsYtR8k7t5pWBhk+/3Ld7cQBvXxsFh0qzqNEp231GY2vw7+sF4s2jkc5QHccblM
++iFIpo4bmzQHfUAs193zY2blKk2j7x5Kipwhe07xtxcDmmT+yLzcYU/ihts1s6WazP/9M0KFOwP
F0XiA4d//eFQVWR7CBfGTR5T/BA+V6diwM0D+6M/vJ5HJltqv6Guvc2R1ZSHGtXEQ3fHYdw2ZjxG
FxkFlckxI1P2q9/JAIfmjLCxNmk8qIuYAooWqzYRBEjWSIWSsDsznaTt932Z/2MLYD32kIywUX9p
pbwG1fe0T6gOfjg0P24XvdutGFVvtPClI12Fx8D5EBVnrMPfNXe09I0zmydEFPlBjGOEizCBzHlJ
FyrC4a/1GPuPOePA96Vc+eWL4X1ITBC3M7IFwCZpCG1u08bnsqV5z3NQs4MvnI9nfggPUF2/SOHt
pYegW5qjh1mR+Y8V++DiXHQGWpZ4qeZNLdhRISl4Osrv1qfFYIV1ERTt7ptfZwLouFeNgXGqI7+O
VQWV40Z8VLaCm44o/Q3xdccTaDqEJbwKvLXymcmFH91ax4NOXDxLWkHsvTjXYPs1Q1hYrSB78yU/
Ec41xbYq18ljkqoPCCe/gQlRTINRoG4RKr0H2K+oZ18FMyLzj/qqA2D7zCgq36d2QUeo+1uOmiGH
WJTK0dwV9dSIMo5JVet9COZ/GEdNfZgLBrciHjOdnsRs6PfQjTUSXKGOnlR6Gw46A6HIixztG7SU
8f57G33Fj86etpvxbT+c6pgyBkpbT+O8KhrfNggE2ySLLHiNZnHYf7lEunVSSZuYVQuh1qYtOYAz
B+zft8vvrRXCISi8TVb6voEQOG6HnEPBqNuF+1xZTghgWz+bhBlZ8RMFOKINhnaQNSonxJYsyfVB
LDeiCkIVWsZjcAeBDVsPXv0x70af04ynCRhawx9m7n4M2EXzGjVGLZn1CCJhPdUxS9UaGSwn28Px
w7+Sre9w3DsZSkue6GiJWuXGPmLWM+nsEoMNTOdsRxyfQaS1BugDIju65EQ/ZJ6qfIFyD+Cc3FGJ
2ErVwJO/uLsRBxwA2O5RT04DeRnsbOmi8BoeAWE6W6E0Pvhrjd1+p9OyIpKld6/XdaTmj4sZaan3
WxJUWw+cmU6ywo4NzKdGIGR+IpP00Rdi/EXeO0pCAGgTvsTpJMDJaOuBpSoQe6zIZEOMjkFrFmLH
iHOBmC9n+csmJtcwZONtPC2HDHNzQT/MJf4wt+yGupDXbgn6VjZyJorWDKmDU2e0kS1VapI89Mns
w8Wn/fq40rTw2bPlR5AOhkQjHkU2Eo1OeaddwTpC1wLnMfh8fRAEzxUuCOBCaD7eC8q3PJvCLO9R
e0sG6ia3QyuRNU6RvBwWD6te2kPy2AkiVQI5axZqXQp/nCZosZj133oXRjqDexM7WODSJRLoj0LP
7aGM/qIqSgwDxrOUaroKPciR3II57nFAI3pp7P0bv889Zp0UHF1Xf95fZxiVmjAbykv0caE/b4er
te1EyHPUvJ2vZS9w2JxiiHoLLpV+ID+GMVyi1WxOk5xht76p+r6AEJk06YJ/sda5Zq069FZa7m5A
iXg0/mRneeAI3MopAQ4sqBciKLvUVRGPcDZTkk0MnTcYWSer2KoxuxUdWwJIe8OAO7ga5VHGlgrK
iLFBxikwfwjhUie7eOFrr1Ed7rbku5vF2pOlJ+l147Ogh/kaYKfK2xjhSFakbisBx7PhPuLiCq8F
9H8cYcWFfKCIXeu145Q9jZ37fXPjn2Dah3HIAzW+7u3tLPtfBju9O+6bONyvtW6WAngjDvew9XiG
DCkL3fwUYER2oe+qmNB006hJnTyjs1U61QnMRaF5EyKetTzy9/GSfSKIRgwgPFxQyVOFbhgRT6vS
1D3ONvAASpgt7l1maDUqxrLY2p4LN1cGQxJuTn1/Z90DYpsFo1hmJpbvzhOklGzF7F62QNjuPFrp
a9m5mAaqbBGTg5Xrcv86GokStH3/LEYhio2r5lkJINBYidrsO+lgQr0OCvYD47nj4YgNhNwSMh+4
o1lI0TAhZ2eXnsdwfz0xwyRDV8W3GrOP8VYCkkn2wmwQJ4u91NfeU6uvIP0xdLAlHlabxDigGx0B
vnhVzgFeAobZvQAJbf8mxu15XDQj02vIHJSwOTcOBYGhRnh1s+CRppbUpPyKcHcEb59C+h9ZuOI+
2M8H9rc+h3VttP0Rnpd98Cje+U219Pd6ytI84okiZmK520fLEKMbCuDSUF4lU68Q3XzMBRMWB5vK
2HO3iGGsv2sQK6YlnQeMSaUr148liZ4acOcO+eQhzezg2JV1xkJRRPKiw2BEaLEbSsrNxjgl6an1
fAWyV4KC8HokXHcTgInnkQjyBsxsO97OlhsuAwiryMVC+j8wUxyXtjvsnJhRb7K08jGwhG1c1xo0
QLPd2Fs74hWbi3M8AWPhiGFnPyObhwOKbPuEtc80nVrUZnIcwCEZCNxGXSS74ya8+APJp7KyLKhI
wl+i11n+Vw77lzT8yJebLNoBlVgL9FDPS/KaW37COl1Vmy5pD4mFf0uKt1Hallqk+ten+NB0pXiQ
e+K6DJif5KjgRG9SWf5n156oYcHXIhyyHRhTTRth/1CDwWs3nTSTXFR0y5i9jiu2FaKPEwv4xkoQ
sPxxWUmc7scoWunAQ5nDGwxtkq9SiUC8FeuEYNoooue38GUyvc72mG63AAUoM6HQYCOzKcZm0POZ
7F6qeJqbvQf1T+Icn5DD6wFvpiXOWL9DeZ5zlk91ffXDeCwkp6vNf8sXM4JjhIztTMMe+IhVm2Lf
sQ4ElLTGLVZ0Vx8UNBKThsJ4azKgfKKld+ROvhw8xM125A4DlYV0GDcWo/Sz+3p+tdtxTE8hkIDU
HOvVLRU2JAl3b1zLxCQWw71qTgeNhdt0wYoRf1Ugc070RMut+6WtUC6g4P1coUm0YEziC8GmanRd
U6fb8YngoIAZSiipJ13Vn5YFetot87uu2OtkSlJInFQm2jShZcmKUGAGjQe+8BFY6Lbdilkehn5K
jNyl+3VEI0HW6luAqNSH8o4k5VNxFElW7/WpM0WKb5PDeLV7F9fY2FaUVA4rAxAe6gqVy6KTXNGZ
YvDUxJ98MnEkraV5XLehlxBFbQ8Q68oezCoa9pmM+xDCHY8E8t2Ig4HwAV3XWQs/VKXbkxhUAH+y
ZdM/xNNPwM2b5QyB0r1olAqdpfau8dtO5YTPaPvwaJPcf0sWdZW2vn8cmFwp2xzUN5JUAeeCujkk
YC7VUfn/lZLLkOxv9iKfVPnOZmKc9Bcy9J/PDt5jPj8MRRr9AX3FqAmy6IBZ7cxiYnae9qxgurS+
UZllxw7cFKr+9+GEyLuaHY4wbFJKYN/24MY2C0Bj98i/88tg6KzL120D1Tdp4YnycXKnCBbwMXy7
K09N/ZVjDgmkcO0r9KW+4w3+UQxD7I0RCX5qXj5zkvxmTeB6/OlQnX1ZOBoeLi95qI5LSpjodL4U
+iPQwzWMqMyoR16enz67GXEPfccxSP2AW0WTmoVOTF2mvzkEKHjPTmELRpFgRLwDNNZuDS0i3omP
PA3AQwxB4qOzcbHicuMk/JcOpg/r4fHXQsgRi1UDF2peKPFTBTgkyP7xTKHoxq7LiKAJo9Iwku3n
Y+jMcd2mMHteXxfWiBH52nCE2EXw3SGIVOE/d7zLBP27TA8/ClAW3PUwJNur03gNC+kbAxSUQ20b
871aTEy7UUM6H1XLzXMakb1518BcDY9Qm0JENukWD1/rIhh7H3rrlkBL6kuSQYpNPj5jDtA8mtND
75NiO9nzrxlTsO9ILiIL3k5wPGsxDOK9WalZKGqNz8aRqjJfn2m2CkBEJ93I9xevQSTNs7uc3Brg
ntYcqtdSomPFPkk9RkebMp5tzYC4wRcZBPrpyl54GhJXPuUy3pPG47J1mxF5T04/4vQI3O0EwbjE
m8wmBiRog64QvTm3CJZ7KbmM/pGKydZjVuJ+h6DZcUkd2cdxIhPvBrKwNGLlQ8xHPpQEN4afXo0g
Kg4qoXKVQNTlam+LdGGckURllRVysPZTpxBTYqnePLrub/eiF5k4Jq2FPHkJ4ET3EsMO+myxNpGZ
90L0DFA8bV2FLAQgZtM9xB2ghRdM1Xsyz9svYtQVFcYGDtmMs0Gwl44SOdzUfB/DRmozZ+W4fWME
Iwg94xJb5l91M26G2msYNSmbGkkpbGRxKDrC3N+8wszuQ1kzEN0xhJaD9uWRO8hhKLjeIHhmTcST
O8/GhKPjCtazVOCXEx6TEU8bGcT8AhBCKjaPxPqTXoLGzoeRVCzGDLLFXkqNpItQAB/fbpJR4WYC
Y+iVIuTqPoyJE38PPq+axdy5/IvSFOQx0zUAWPM/ExCkCVUvYxqsXYudk99jOXV6A0vwZPNbmC+f
UYPTtk7nHzEOL0chObsZ/pg+c6ISm9gIwwd6DDRRTaoBCcnaRJ+VcXj2qqEemAHGSEO4X5LKwane
VtrcYntp2nXA5yRcWvSjxjYyU300NFIdtQO2m0y0wQ9o0nWN2vPx1HbOsbc88WfOmYzTQrHckKcQ
RRaMpeTqXxvRpxRsxJrEumDqEOyYW0n0IhU07bWIqaqxdChX5+a8BQ5lr1qlWLSsA5wMRS1fGrAr
OXBkPYw0Xy96gdqa7ai09KTKLuR+wJNUHOaVoj10Zx2D/VKbbZrRS3WK1QOV/OwggcF/oCd1ibLP
UYrk0ZKutERGMYQCB41WjgFHp8EAAfRuTvxN98w8Ryt5FejtNeO74PUAWaJhtx0zijhlo4aWK8/5
vOvSn5Q+aXKkoEaPDX3+bXiM3ZJdXjwKc8SB6zadz4NmVO0zPHWfADWqBYJpdPH/ATr+6PMQjSM8
lRGVhf2JXOYks1rapdkBgNLFxn4nO15+8AywrzyPZCGwNZDs5gfAXeYUmtwwz4ZuIQIThx5hKgtV
Sr6erKRy7kPeJOE32CSwPShptYLlE1L72osunXnJ1gCqlNMRCk7eHnqe/RshQsejAOzcY/vIG179
bKf4p/R1ImW11EkrRFMpxnwfA01x+bosyxNA8h4fJf3TeAboZDy5B0RH88RYsCT2z+LMM2Zbc09n
13p3arDesNpLEm3EmsH8FA5zNJGlEKkPUlPWtRMZWeY3iOQxmiaoWVxDGs7MoUcPV2Xvp+OyNcKW
Z/srU/anvoGM8gEkZASuLJ/gftX3z00ghFV+R3BXYkqVLnaVuhDYcRhLI2lfqxguHyyrk2xEMFf0
qNglPHnk3ev93ujBIMeFa2T8CL1C5DIoeJt9ijl6zB0TcrNIkLtqCloW7LQO93QGYucuvafGVJZ5
BQG/VX4KRnhXoQRBVv+WHJMg/8GZhdPHcWenFJ+i2yzGv4DsAZ/YBGMt4zCcVWAapYqkMTSY9FAN
NmCJYek30f4xPA3zox/TT3FWGo98cjGnoAJWPimaQvt51qapCr1z82ZHlQsueFJY+FjsGfShkqTq
UY+NIxklgUJUvOra2eKQKZVA3VLpnUKhsEhjAm3Zzh3XiUeXU8v+dFbzSuXhA0i4W908zL+kP+AR
gkoMZFk00fkY9lCYbTL22bK11vQ+/QYSHkpKx0jwFEBfp3A3vaSRWeg4i4czvX73u62gasAm1JB0
tnMVK4q3mXBpT+CSg+TboZnaqdYL6sTHgnqk+9j7/UYYY700jgYWF8SZjvPZe4bGj8NTs64YMfl+
j4eq22V09tUr0WtnJblKH0vpQV4ios8eKazddXFQ9TeZiXBz1z/6lXyrS0SPnIArCBle8tawjT7c
mD1OMhuVC6BpQiyY8PKJCRgtBL5MgXvsFG/EaFS+UHIRXRabafOzrdkd5GoiLbarE1Lmk8Y8i16z
kAR8CMmP6wiWXNux9mMWX8CaQoASeiNImg8oDZh0SzAsWi+LmNPatFNZLoA2OPL5mcxRybpPKcEe
6tzo13YUKyCNgxTLsznewD5CT3sJ+8i3RobiA6eDuJNIzWvjd+0JP/xE1BCw9RzF0jOdFDCxrwic
/j3QnYPA/MTVDMdozpCyVVo28SDskxZar2+XrI7MOlTBfW42R1lz+w6Jj3UMZyfNHOQKpujfeoRP
PoVPFpDeIyvIYxu9iHJd6wZMkbIT5MNAXyei70UCY9iK6jpcKVnvbhuZMGffZD0Rfz2cbWsG55/8
XoyHnIBVT0Klk/aMoQHc4o0RnrZgT90ka4HTwv9e9dkJAVnwmuTlmrxfO2Itq5qETcGs2eZ7ptI/
o3MKhGOusyRKm8cnnddIg0lYUJgtgwbaIe6JPbYcCn7sj1H8b0MAzZS7tjxL/ekP9KhSLCa3gu8z
JP10inUTwrr5sqh5xfMS5RyPl/sG33rRwVLQtYlNLljWKQ0w1w1t5Ocv4meNyo2ielNY8X3Ll6xK
fXXW2veT1Rd5gGJ7HHXVfDV5pkozkrfULRHkU8yeBwDy0axOzu5FnY/vcIo65RZbwrEuWHjHpG0j
RInBhUCFQOvHyVcFUTkhwVBA8qSazVx5L3jLNEWVUSvVK7rs8/KPSjEtnLtgEgtKZH4Cxcu5+eA9
bAreEhXbkYZ+lpE1UKHSg5xJiubhnDtg1B/NE8q1U3J5FlmJvAHu94Wto1Xog/iME3s6gJ1bOz1s
FnZxH689Z96xs/IbUSgC1UxvqL6edJmE1rytwsKQULRxEvZPoirA5zQGXsAs4FZRSmc7PvuAm4sT
WiJTuHNpPALD0lnz1pREgOLnzbmDTrKmMVfKW5uebNzwe5KUHDbONPjtTjH0fKTGKo8Zh7OThvqA
d8hFSwN6X7zXF5px3xmLm9b2THSMQYDByqgwYnO4NzHR+c+QmOX1DBCoqYZO489ZY5GOEj2CkCw4
SqThdFnN/R3ZYiKgs80R/kmCk388E9cNQ2XGniiS06OgTiR8JxunrFQDU2Walai8Afc/ic7SU4G1
D3ml/JzVn+7cxA6nKD3yktP95W61BQaIRE/tIceLAte00CV2nZTHqs9SfuHShdxLwiffes+CJlEG
m/dzmglLya/NO1T6qXDv6iy3rcSQ9RP7oblkAWHBYHRp4E4/t+yVge+e+Q5rqrtmKVPikoDAgOSi
BX1BsQMHAPF/EyBAfKFUlZT6quP/siKoOKnIbxt++2UgLUKNpwZJf9BjFjCMkKA8JiX6ywInBMN3
6pTK7Im4Fy5jRzEdo40vMOQoQR2+cp8cO9mLlVRYhFyUmTmilK3N5TVQEWQbFfDgTTSie3n3CCQF
L7PcUwkzUEdc+2AP/dX6Sb4zYvmbwUxZFk8p34iL/+QxDhSZzS/sUUy081BbAQp2g/mm9v9wigNA
2bTTvICOwMQrWWYwmoMV0JFnCPY3qpZsDE82m0aAs7QA9IxLCdvh+RW162qG/fBFdvWE/VFq9B3Y
tlqVV00Tq89UDekLLtvNy0Gwc6piUxhbc8r+5WY6ZMvRgaGItRGHwrUfRqUaQ1cmFN0e/mvG34D1
QprKo2OwWZi7coLFw0MjM0aH2y4eDVmQjWrYfhdLrx5GkuO+srwvniCSKdCFb/ME4ASjmBQmtgqs
SEsyHGsm5DPjXRi2aToRcrl7i3JHEcUKjgv7vCSUlZZE68TiwcQi6OY518P3yv+R5PMb1zERdzNN
5eIy7xJmOWQ8GVihZbB2kViDd9SiyFFWc3gsV3Xwe1cpeAiXroWiSjFUD4WAUz3zwmpCxpMtIuJ+
qaeyKu1YyMlj3B150waRHYUhEYlcS4Py4JK4G4XtMAIA3TnEDMtRKHnp/kf7R5Km8mrJBVTZedw1
CZeJNZgCklR1riAVGjYLh8fKXX66wGNKvNzVFTQi36kevyOPToqsDSPIp6Kyl7xwX5zAbDuHs4Id
3c4Lv5tcIHR24ZaKpGSNW6LSxH2ocfVLaroJp+0Rbe085FG4/sRQYYD3bmDZDNJplZeUkT2J9Shq
rjHKCKSNyZtZ5AAUYFZQpVnySTwWwDB3BcLcvELdS033ogpS/iHSyjrRBsVsma8oJzJCicfE+2i2
hl/TiZTA//Y1Bsac7pNoHeSFvSBLUGm8aYUXfM2mXRPUGIHn4ha2XKFbGnkgDqNK4LbGiSQ30OKf
8CyLb6WhjVYtQQy04akl2FctR53tHACxm4DCpPbqEDUps7aikmVwPlOjIguPgkpRQvw9QvgoIkMH
L0BcKBkczhKxdNJtJ0n7BgO9bEo6SpS71GMJM0uq4ODWRjbc64oW7wO0OUm61NSK1XYTjfVBU5NP
RIdDUHJsQ3ee9e/CGBbvVKlZGQDP+5w/FA0yTaCQ92OfOgVK4KhPR8lUOGtibl4NrCP6UTubeOXb
pDWXK0KOGp1jcjOF2FOBdpLvXQDcNHuVUBCb+OIPi0AVMPm8ps7HuYIdgGJql381iWyrXaVUsg1n
QlbxVEYoD30xVnmWAcuHwA0yopKBaA/6lJ8mTQWEQODZHvSBbWcBTrB7rS86eunswBSs3y4rCG/F
zMYytRSweXfIiXZflftmMU6kBTR0SpASDcUX4NnO4Pf2LxE5CLZgqXwiftZXq+aC2FWsOPg8uLSw
Vbon2FxSWfq46cQGa9h9NYmWzZOHIyg5OdGbZ9Hwm7AyA/waklgiexDwZdSfKPfFKKVq2XA+Dm3P
n1Kdjdcu3c4bumBuFzGB++FH3A8iGyJbbN8Bds3aw6taCt9VNB1JXiKqAuITO0yjgRu7pEhzwGgb
mTbm0PlyoxCRR+w5OnwoFaDOtGYN4v3o9oQ7kfC9JtJGDSScimHXrB939YUvh2FYOeNz/jIq5YH9
zakS49Z1QVBJiNqg/l1klAMdRlFnHZ/7+aCAf45lD++pbhEyzk47aqEGzPBgvCmW9ADaZkIu1gkE
4jrUV/n6qTleLaUfriZntoWhPbTemIrQH6ynJn+tTxGlNYK3le38J3PYiPYwpmVDOHTG+ztwMabt
uFTmFtjNc+UwYMlhs5k/vNgOkERh6+dgyXKPbh9OjkWUwLhPBN1wCPz6wt+bn0Wxd/Zxzr6uDUtA
cnoRBHl9GqOApkNK+dCKV4J5Iu3QwlGrnOsaKKJVb7PXmHP3vIFhDSbCtqPU0D9djEA/ZyXLWMAW
fJCRJ1KIuKsUBBEcFxYxxHenplF0UjgSJ7XYwE+OCcxRd2W+ZYQrhAv7v/7Snwg5BZ+yXAh4eAux
cONeQVxYls0cruPuk0lhXxboU3W8DSIR/WxluZ4pkaybXTcjQ1UgXdJHSNUZ42xt91hz6iV6HgbR
U156O8vhDm5xPtiS+4IOSY2MzCuP3ZofHlh6dcMLJ2buA5JIcXpWxfPd/Jd6fxElZN3uvbN7WpqZ
5amf27GpXDXoPrFA243P5/3MbM7LDTjBPfe9k5yvOvEnME+6kPCA184fEmEzeMndc4Xunxs+vLqZ
ojES/rCpx+Chq0smFZ4IfwRTDf6QYl/gNjMKGzE/Y6mykwQj+JqeSg1KLWs6Bc03e0QMQhwJGlI0
0OiNMH54wlJn/7tH+ZJasC51vpuKupy5yw4xc+Ef8aoKaoLSCr+lLX61F/umJ1MZakvMtrPGVzGy
EAcOcMz2aiwhuamccDNafoAJLiGKyCpb1fXrQQvm+vOeuOviwmNKzqtG1Srvi6D3hoDZdGTkmP3n
Sy2tRrpV+rJVnZGYp/5JZqn6AYWpB/UlVvG5ohcnjDMzWrt2llDu4KHLMN5SZLGeMe5/jHgd3E7q
ef8LRC4pi8ioUbqV1Uxj+PKRBppjAfsLLfIWfYgkpKZy0heQg7CshAoV2m+Hz8PS+sf3KPeycztB
9/xFipAllAsz3bvxCGYnykoGUfmY48BWE1IMocwp5DaA95Eg2AO3x/HnfW4dxaRZl4qHlO1frLwp
pcvT7IPn6r0zXcMHXnQKdtYJolw8tX/eUS1z60IcfJc7aP7gjZeyuLfQ5WPlg9izUd9p+hFEeYoC
XwtYofTsB7TISvU4ko1lsMKIimpb/GLhfbUJyVA9gTmJf1Qqx9PfjOpJ3HTErYXPqpWkJVLVgEe9
khPt3OcN80Q4u0bBTlAnCw5igUvv6HyNXQ8BEEeLoheTD7Rr4pob4tcwZKKvajopcoHlADoEtsUS
mrtki67qhU4S9T3PEUN+Kxl5vYjNP2hMZWinztKulM/emdaiFuzUaKHmlnTnNBqy0VaGKide4/hb
cgs+xJkc4AlaREaXU/hKk5YS/jUJKZYjWUfMHFLaayzCnVru8cAicVFAzbHJBgjpiLsmwCW7WKGL
QY9vFZRPaSqjHbr5qY6jvQ0zSYRSqTfgDTML1IJ6hGeSO7PxS4/fRCdughNwrAT8n/BfRUuMGx4G
HDCwg1dd8Hy/kc9L+KHZp9EFU7Hk2zE6iQomcaFZf6+ebVZvf7gzGEZIyYKjhKH1+7+gq405y2hp
m85y2yeS/1Xo/PESqn0BODKl/Ywr3585jO1lv5TGMQ6nUXPvOlLu6H7fL3tDG+d+5IaUMA+8uA4c
6j4fvtjQHcyUMxC6t27MBVVNaUVtNjGcilhYJIwxvrXD/lDcQiUowpvNmS2iYMm7h7UUAB+jaakH
OdniIoQC1/QMP1LaErqot2G746YQhYbydhvx2jVlkMeV+ZLFHCU0JYJVmmODgp+rT8Adz4IBbc8i
EUVepyho8n82S9lAn//Uj4OpFdW/zh4wdAoIrmxIqc6epKIEuRG24WSYeCC9SZuhRDEYAs7OFhzs
mUQb+VfVQSXXCN5FVsLrYncwEnJwOAeUQzFhzMyx0B91NcD4ym2inFo+LLB3dTcZ38e6yxspuGeq
eI7FKMaBZDOxSgUEHF1Gh3mQ3CvQIjjwHNIwQ3Ihx2sGddan1abrq8L8whRP6+Zsb5eEWXh1gLCV
yQByFhqdQNJNfY9ND8gDbNCv91tSDUIh9EXJ7yz92m8GE8b17WqmuX2UXoqxoG7QCv1n1UFB44ug
MHdNkSHS/2eP9K/2koMaKYuSXBsvPyYcP615KS6U/vGXcir6II//sFR+ZE9z435704sDpebDSN92
V/cYLpTVMFo41iFNP0CIf3yJBPNoepUF6tgOERhreWSVhzUF114tBvdSvUfE2QzNFUG21HffE6wR
ENjDcywS4EF4X9makTOH+72GlERevJdbeCLq7K6yKByxQjkHjyrWHr6UWDJun/5a/1xuakMGIgbR
Ox5ZFsqtNLGq7JbUYeBhTLhzbXzzbIWTSGj4In8/ZlN7EbXXmi8HkqTlBozNve02oM6flGFi6Bbo
E6ruHxkk3QJmD5Sytr3c0YFy0yGiKRcuj5WeQ02pjStKwvNawBMK4J8nROfK50sm+mCAPTXGTzXO
2c9dZG2kCPDAeY64cKl5h0RrPzJosdhHhgT3iW3W2JZvHdTbqLZLLDpvtexslQWAKW2Ho+4MPXoX
sloU2T5neSNGz7SvKSWPMB/ez8AWO2Cr04LtvcXw84GDRr7Im9NsI/BZDvKsbfqmJZ18CnVbez+V
4qSrnIVxEbyvlSuMV8OsevAHgkMmkDIEdPjqv3jKcd3Y0NQ6hF4wzv+n+UrKKvfrxDt0VfzwL/qd
CN1FMKHHALdh3i6GcS71FGtS1IpsZBsYul4NUn7j8b5Ic2nRxOVwqu0Q/COMOGMqJrjPZmtSOAB8
6xm6NH7IlqPZRs4VWkY57LTjI+1u/HieH//N92wh0HQPFoZDu92uWw5z7o+jtrl0lCueRu2iIGlE
W9ff1KsxuWR8Ls6R2MM3nSP1kkQovxB0muZJ7ipieNaD/KVvy/+Eloe8ydts+HCdQV6aXYgg1jr7
h+t63pEM+7ncw5JilSaJ/04hTuZ3Vr1t58TeFehjGoIUfze5DvsNxEW/1hZoRBI9ryAv37xWiQXe
gNi8cM9jCBgXitxFS8RCYOHPpaNDSx4fuozrP5iSf136GGYczveLBEqUe7CkOE2RaeKM8vBB9LCP
Tn2S0gTbDhPRDVHWCQLInuUgEZarsdCJ8MCgAKXuq53jznHn/jD3yDRPzzGsx5alsT0Dd+gG5+Xw
9bu1c0OrAA0w24zc+gyhe77DgG8o9J/h1o4lngH40cb75BkEwWKhOEJ0ifouP3hD9i3UVTrTfV2u
Y7xxWTUeEXp/x7f1heJuQakpT/tu4KqmOMjnMiwrbdQjLy8paEKCEB3fRqL9uGvTs3jU49O2Wd9V
N1SEuLA5CneQzTpWFE35OPVDnhW684CnTTddcp7mzlaoGlZRLUSw30Sqi6n3xgtzlfeuTl3xr2IG
Exd/XmIxbDNPlQ92TyA6aCUu7EoBuvrZxxEDyL6DBm12La0YRfCkqVMpfNC8efkwAcBRDbK9j66b
0mUSh5GhImqX3TABNj6fXf4uRSCWUGFSVBrjHdzoVfjZklZlBMr9CmCDy0Io9JJ+sNJqG6pneS28
S4SA4DWgKekLWoRrIVEaRHehXzKiTQOxYAB33lPioGjDpIZetNutqqr4/qFMGlxWNq4rlmV6U6ym
VYJxP3vVfgmcWCVg0qBEKhAP5yTX4YDGVLGA3qZ1ZhUs9SZUAzp5fSKz4qHMbraK87Ue59NWUsno
wiCDD3Xo8EBOh7RLT/bRSLr6nILgP1rTicg4ryEt9eKK4qrrSozR0a3rbHlGg6zboUnWI7rkdFOL
3ZFLKdJfLVkFR/4w1M+aey0Kene//qhhFl1tEysitmrCBRFyA0pAdQQmRk2dpysMAznVRq4nJHCj
rnocEfonuOAQmPFn4rINuX6EWUMvEdpQB4QHJSEK5Wnje7UqHXuasAytWlp/hW6o4lJAGZeM70ae
86sqzenANKho7c0bhRh+h7ZXDo8IUpd193PjAvTV9rUF22R74gF+U5XMgSo5aJsQD3jGhiv8Jt2s
dfT1v5h0CRHUQRcdv4SbSYVG+MO9mJahMG3A12n4re8mPIlBDF62eLCubrFBVD7gqbDmJu3y+0Ea
agQQ9GSvFQE4HfJ80LL/5MhUSlhp1Ku1QinbScmoiI5Vu6j2Xo6Lmlu6GCj/ihv5GvrTN9J05BBE
nPMcnigIGDBGeOdqhpsR0eunKTMFF50dEpO6//5X7bOdGX4zAad40bcqNHXcLfDbASoSaPWQxLil
C0u95eDs8s15tN1ZlxcJ3gteqCS47jIXG/ZE78idK730bX+1IYZ0DocC8M9kyQKOUTDH+KltTYdR
EUplq7mn7Ag/IuWoAZDFxuJjc3JXxbtuy7+3FsGDFPk4xoNCBECiSPrOpwiGaxwSXrzL4mcPrB/i
n40ae2Ex7rk5nLROvBIjzFF1nkebQhO8e+3hKTsJ4zg2QJcGPyljY8HD1Ju8xtzpzT2ppL/JOcwF
VUmRoifcJ6vWJH2tB33OWePWL7tYv8G6MpYBvL0O7ztaE8/ajJ6xE++5ytgYu0NchuH2mQU05WEr
fpccK79toRFZSykg4/1D6YRquXFwp7WJH0p/jEXBIGv3pfiMq7Ml3thqm6TA3FKM5s03VYtgGeQF
VKQJoBZ6SE1s5DQIcNOZKoJa0dzm5rVI1WJfc6m8uR30yzTenJTqbsUgW5Uy8SY3g9QaFhfWCmb2
FwwMBSbWDQ2lbdgFd8uvdwJpQY3hBQGTcQQoSWh62ib4Uy8uiitdkco7RuiLu4kzNW7OuLYmQuAM
nEtb8JWfECU8k4fGmKbwE51Ouy7md1ljXeLLVuZFkyiyZAGXwLImltZt7bZlyS2O2ShEfROpBPB/
SYrfnt2UcxYOLlIZREHNQZLllX+2bBih2Q4JtBflHFjsz07u9ITLYjwZoTobFsaTUkHHnV2qqSMR
aCIk0WbfBuN0qBf6moEp+FEQZYAW7svzZqZI/p0Zf20zIRGqSxAIIR8smoj9c4RzZD1Ax8GruhBv
HLXpqidgGUAQZPRLogg/Avg9hY09cjIsHiNM5+bBTu9ioMVB4aPDQUaPPezRHqSt43nbQ4KpLJG/
ZQOe0j7M3qFm/3hvQfYrjLrxv57GPF6KNwFaX7NaF4w8//nLV9OImnR/Zt/tqDIo4XPyBWPyIjPp
2vdcvwjCSW40pP3tZgypp7bPK/eaLtcVPcRsFeN1DJEwcn08Bk7KMGU25ytF2abJRxySyTv4m6aJ
xXw22nmzrfujF5TpywLloppZfyu0GbzzrWX3n7jLSN8l7sFluTV0LBaumE+I15fq/139N4HpN4Ow
SALXgV8I266VB04hsBp7d+9xPQGpjjMjlX0KNobMvBOdd3gx1Jgp4SliBjr3MzC4mJcxbvMWA+1B
/xwM+t6ko4DyIdjbj7CeJLdFyfcmN3JvZtU6XHDLcF3jtEqpqSwDMz17JXw0Qq6Pkx8fIs6S5Qj3
BtieNvL7JQdPsljkofm5T30rq9R0uBi0sXoFVItFbJEC06alSsbBvV3X3ZM3JoMUs5LMjzCTtsmR
YLvB9L1psdR0RRp9X4mgX7+gcpc5+l6Ax3Fn3MV6KxqEz8gO3QaikgzT7jJDqnreZuBr49ElEBVR
uiV/pr5ZJqcX7496ExwoxhDOqOW4yeA7QyFavQJYvLWGXnUMonVgCLnpOw0TeNRMrdW9hg8rxnmd
soUWTDXL9WFPof4LY3DKLqXT+v6/HIbYpVkIsmrhSNPZFt6j3dUasiPiRih/zwsa0Xitp1syrLkW
T+ZTsAzlY0dOn34v1TNldYV8xnE+GYdgAIxwgeBBWrWxwmokGr2k/4AtsGAdOV2x/wit9YKuJhYx
eH9LRb3QlRqKBgvMfkeqaLaV88/eo+/XWdP9OLZRbGdFwR4NQI5j/5Ce6vp9lkUP52VBXELZ5Vvi
I9PNO2mspCSy2Yl7+xked5YxC0ndVW/W2JCtCJzpe1XYk5H8NsWo+pKEjI90HvlnbF8TXFL39oXV
hQ4+EwnHxw7ubmiHIy8WT+RbXglC9RKayjMkwOEjeoTnjzbNrvSZHiSPttlhnoLaAl7LYyyI9o26
YoUIEH8kAJJ/hxiwnJpq501VvQuQIq/XTecq6s+FDPfxQCXFGn9KX3UlEqkdBX2uJollh7X+hRbS
niMts/EKEhNTVQdO64TmnUyCCx895LLfCEib3/HuAsd4lW/eFWaqmgnYVhv+Wxt2eEwxUDptWIP9
RpcyqGEmbeg72yT12XTZKaPQ/L89x9BKpQdvG1Q1kYJBKWQk08woTOKZKDsbwJL3E8GgakThfXmO
6FystBvU0oETd3pVoeFfeV+Qjy+J+2olnbWWUKkUi2jdVUETUfUP1ckbcP5Mkt+xo8cOBuMWB3Zk
2SYiRRwtznO0ugx6NJtY4y2qHBDoii66+08FxrUIlkZtKO7tDfU9OULbho6codnEojV6eMmoAQyX
Fn2/rDJqRBj1EGhVy5KbL01ojLlwL40R2X57dVdq42Z4/mq5D7CPj3akBUCOqu9HzbxzNr9ZLbiQ
w32n6bJoJBE6DOs+ZIobrA2hJK82BoWThM/eK0yv30HXKBbcJTQefYmooCBRoIIF4kMSmW4aSXBH
+iGE4VqWmWGtqM1gg/h3y6OTFkyN/dxmrcVqn2IxqPkn9t3/Z7+T1vn9BXwhKCDwH1U5FJd1s2i8
prVNzbRGLHnWxjwv3QpNVMazqqspAtukVANLsRED0Wf0i2InFlJbfyDw1M3tVe9Ab3xOWcIE2UOQ
0GJwEVDgx1GClemv19lDbPjeLb336f6pxQax2YCMce/yshtS0Agql4+napLyLvxBLclF27GDufa7
jN17JbxVeGWvsMcyXaClZip9YqpLFZaa+G9TUrFYBtKfb36p8Dl/k9UG2VgNmkjoRbjfMXLT4lSi
N7k1EGK2XO9gDkyOTioJ8Mo+SDxreOJDZrinWq3yPXqmDJO7TgcJEWuNnsC47dIreamXcbU3zZZK
ZTwYhCXAnqs7Mq1GWXXpiSr4yfRQtqQyEDrs7/e15wz5PScg30kSst4awxVdtM9R3RmoQziJ8zri
6g1DoBrw2XLQRq6zJ23vF+jzEBNOlBT9YlbFG7GH+1iJpqlcn/5iFaGdz31Lhbdw+3WQrKj3uvGY
G3TeqZypcqDnzrGln0Rnt3JxqHT2wJtfDbNDpCgQv4CjEm7vuIe2/Jyakm/Iu2RO5Oy56YOQr3GB
XDBqlmrDlqI7ptqrKpBi3WiPtc8aGDoKDRKtSDzdXSzDp2he7K+RAI5NI0mVni9HlaQTTiJZdnPg
uAgBZneTZq8+AT+tgoIu8scIuOolzOlWCklqnAuokyzqmK06Bc/6i4KrW7P+M77qgB8+0bA0sy8U
XFBL5f1wStMGpffsk56jgh0IZR4lJlkOED9lsSLC1AbbDqpQeGYTJqJvnW1pwk0uvgz9zGRR4pbV
FZ8Tq+20HybDCCxWInk3pi0ykZVaP1lUQMles6EpbIqaT+hZYJjFH6Hp4pR4qubIYcmB6gMc6n4P
SSB8wMugyJrjqtpAtpFTASpwDGjjREB454QwmYb+0A3oQWHA2JZtATBsckwCCvOrdFNSP/JqSce2
1/3RXJGh3vGCLCzDwWVTLAzToQ45hG7IHDELpc81GLyD67TJcGPwBJ7eLdlvLKxZdpyPwUiYCidz
kcfTZUR6iLW+o0dSa8m6j0VT4U9GkTaWPld4FaztTzEU6ZLM7q2QBNHihD6YHKwYAR7ooeJs/tbE
huNoB564D2F1Hbbv9vyCBSKUb7dXd3X5jNKL2HO/WVn6cwB66O+dC12qsLg4cW6KW3EyWWI0KEaq
HEfPwB7lBX0QxD/LYrBiBkS5rSs2+4a2DE1OVYaERLR3kwW4D60zzN4Je7Pw1l/Pkku+WVIRD5wD
W7ksz5hgqyVe3H3LAf0jh4lAB40PCmvIDY5mU1PlRqFvg029Xys5ikuyZAuLnS8rfOum2O0TLEdl
k4hCVn0+qKFTOo9MUsHfQ37QlJjfOdRpToycU2+bEDck75jHqRvXGxiv1l+blSBHGRn+Lk6TNNEP
n93LB3/N6i5LJ+6r9O4oq6c2Xa8Q1KfdJorhgF4SLwTw7Fsc4L2vJfq3A74DGcm8brI0GukYoOYi
N1kPSzll76+/r2sqjqyMcMPK/P5QsN1mUed27xdtNHQUAMcO7kOpc3SV56bWtt9TeGyyAh1/mLgW
W9+eiJ1eHTK21addUWL5nJMrW+/z3N6FPANOmsX4k1ubwGnqO/HoTDOSRugH/8Jm1iHk5uOQKmxo
sD4VKtEA7TvUBIyAoEKtjK3W1WCsS+Q5DwTixs2rzxqlz62wheip23tJsvqPt+ila02pgswXbo7Z
jjzqtPEfVyzJfOBDKZq0ooZTJrVb4JUTE++AvQ9V2vCyD46zRFxHqkY3wsvMaTbVgOk4W5dZPInY
odQ1z6/ogmS9Z02GYDQmxOV18Ol0grSZwPGx69qIiV/Z2H+50GZ5fJBE7OG7/1xNi0triDmg92so
GvxUCVaOwH0EtU3Aq/CtfyAgCGghJ9AUiktz+PR9p5WDaGMz3bA5iMFz57Usj4LVCSstqJ1XGl9b
cHMoohy2txPoc7n+B3Eu800ON7vcNmRCgAgn8a9SfYNHgyHl0YIOtHg4LXYBxf1IJOqa91qrwLVN
Hai5PbaXlDcg59VzHMCdliZVNQdMJXcbxmM+0kFxc/2A3293RQt+M0IPD5ehdrXt5Wlm6MQm/cSc
PYULOtVb/IfwyWQhO+5eSrcye1DFrtb3jsEGRyHC6da+FxAmd2fzMSTqNa2zLMfCt+VzYk1S6eQg
+x9EkQOFYJyU7LIqckrSKLGgVBKRNvcPtOtrZStVVJpFqx6s9VCVn4o02zCbaJTx3MjSK0w41h0x
XRXrGydTThXcv9ToX6RGYLUkq1twyoaa5WRixX/SKse0l5fVOqyoT/aLKPVgdkTXOQ9syfhqABc+
vwoRcWgJsvsztrCAmy7hQZsoy9HcRQdQhFfY4qwInXhra3okwNV4CDUHCb9VJp5Va0GGnwb4N6U/
wM0tDolkmZAgJvqry688ib+9xYp8P5WE8FgIoZUKgU+CFWLYWL2uXLah/DYlnRwXyAq7Yvtb6v9o
RmIYzMB3L6tW8X2/OSVPdeaM84G09qwMDVP9TT3snDow4XYbzHFSYgQ1mhWE4xL5mh4QLf/v69bq
vSh+jiqWm8tm/R0UyYWslPXiHJiOmF+lbEOpkoKwNBfNS6YKDkGu0pEE5EVww3YEJ3dx8OCtV5ml
pzhDVdiNH/9/QJ5cjRyr4kDruMKdj2QnXTEqlWpJypmnb/H4OEAwODx4V3+6Vy3Ijkze1lVA4cJv
8y5tEBmTXMgn+4Q0naOFufdNVZCEc60f3iTu7H5VkGSstBuVxE2/i90UGptXGeU4Whlwz0mgAOXq
QrpG1k4hSW1ytoUmM0glV4mT7QazANoMg5ufDWtxVQnxndZMZLxqjLokt4K3feygYbT8AQ8Gi4lt
Wtx10pBv8yiwf6ctcMgwmmRPayu34hU04/vG2fMjbtKcDp8q7vpLDRtDQmBJTCNOVpy7O0T4xAI7
e/ZeUmtMrxOiHL5435T5Yf2k2N4XKbamqslaglSIntxhS34PoyYTNAMcOCvn9xWjkmzHuQGk7i4M
Hk0WcKUzraCUr7PEj33G8UKacrWH8iT9wUQtJXgNaJ2CH2yGD9AMlJsSkhM3RUu9AIP+rt+lUSNQ
HxsV9OOwI/8CaQHDla8ANlluNp2evDZVrg2Z0rOd0ZZcz+45UQq+26iV6Da7+WrYs25YdOlyZvI/
ZfqiDGU40v584SdVn8H9yWOfcON5nrcAvjkdaX+hnkTuB/kGhtJLahKdTePXFSEgXeypTgNtsfDT
rrdIaBnt2BblrZKteFqGWVIXEMEpMoth8UNyjwhuvqI7cmwndYswJqaxfxrLg2Y4ssz1Us52Yq88
NTB0rKnHdxEdvIO2Plr75wOnwOf2WtJyuRu0c+jOUgEd7GCozcnoS9LQpBwttn/BuPNgLCX30arf
NoksrE5FAIEG9jV2COBsVFfaDshjbk3leM/CRiQbEaJS/Zuwg/Ytd7xO7A5zLkYaQa8wAZ50rMmP
U4kyDyIwMqmZq1d7lABQswsfwvcXUJwXHk5zk4df8olWyN2a+YhcJQnRXinTC29lllxaqtOifdIU
ZcCPPCS3Q5OTMykUBoTUIUxTJc9Sx6wW/QfNQMtGGe+TM6M/+sMnGFA3yT9SpduYLAXjmHyYP3PC
cfYr9+PHY7EyFbvn/zOzQcLEXT85H0qLVRw7fn5O7TcP5GbaWdHFRFilFcJorfpNYKk0g0lAVsMU
cJ/mIKVmXt4TWWz2wIbELAmmAOsYLlph6FT77XVeb+1jli043pLFKd7ax1XVhGYMa7RQwalK7XfN
8LkaA1wUu4I41+IS+XH3ONVkS0RYr/Xb4E2Bn59ShI3WBxmvWrOoFJTjRmMyFO0BPfxYcmh/M7CF
008FUyFX4SAqQ3nxUwiUoDfjDSBjvTje4PthsRjjOuhS9srZvciXuOFdnnLmeUDRlLTFCg8JVqmU
JjGzH82j8zNfu1iPcR7c+SswghI8DkE1LfJEbat9qi1ltEoprXAuZfTeeIyY+0+zs9yZYVZX9A6h
PXZ56XaakxiObEShAvDDuPym89cBNS/Uwk9l/pBfwVel7xN4NLf5FyPgSNrCPOO69auptVfy2tJm
KMlCq1EtqTyXPwn285Zvc7OP/H25zBsmhYg51QMwxcq7R99+/l+uMLIGTzanCrGD2LK8sUDnoTBZ
5EEHoPuDAttEgUsubw6ba/rbUgqcgo1JN9/3TRMyj9iDWidpg9lbYtxstIt8aCd3+qUQNyvOORSb
izY1Yyn4bgbkvvs7HLAhfC055wu5GfkNL2dyeJ0vDopUSjlVJ+CMcFizhUQrR7KIDfD5Hmk+eTB4
tNAlM9CVsuFy5al0m1EdxYVeUstC2OET0/iKMr5JJL+C799LVukpiWg7io2zeTkazkiigpGJmuYn
M22GuX1aEzTDgZyVrtTcqmHAwugRA8jvxOSW7WN0vmM1oddRYG1SKw4Udt0iYFy45Assy0P+djcR
0jBPgK46fPrcb9JrGkGUHpHDHNwyqobM7Qp0fUK3peBQ3UewnECNGDniaWBMwlbDWrMGdItmA9lV
q0q8uLrkouhxWUYX1Ew/obRTqFtE7aXy0HOeslO3eY0MbQ0l4ZRDt+LRWOKRg93AatIa6OZR8L8w
wpYvRTbvAxA58Cs2E4nhCzx+CuGmDwMg4V+GbQPHF32cqu9hKyWcXz2UiaLrBfal0sSKpOqmmK5K
zmeEJv2RYwnCNvytu+uyeHePsmthuj9Jrs267W4w065M9OBgk5CoH46fFLiPwDLZX550UOJqm3FQ
zfYsLxvzWX/E2Iclb0pbwQqPr2PpZzVI7oUARj6fyr5sAFMQ3+IyNk8y9vllM65QlYIVYchDO9k5
2kC43ehbg1+iFH8PlkDkxZnrqG8iFxAqk7p4ahkmTN0XuBh3dCapuFSRgjBPDHap9WSbTieJjCzI
eB8yarjfo4sHaTRitip068dG6H4hkcS5O5ei3Yun5Gkqlj7w/0r1hyGgpf/meIZRo8oQB91YUZCD
ApzpYxFNRmcnvAJ3kzizSRI6YWRfq/9dDBZ/XGsAi5LazRXWoeWf4TpF2jTALdYBHK9E3Z43HZIU
69RTOLQbWYuEPNL7yx/B2cLb9zuBB7iJ64fS7GPLvFoc+znIcGNW2SK0lwUJGhDKyjIbv5iYZqbd
dBw07yinTXFButzXFGSVAdzFoT7l9LFO95S+XRxlO7uNBp835vt3pqVTEuA5hxcx7WlTYekBNLgZ
3e7lOyKd2zsQIe9k1VnaBYcyfrJsH/02zOch77kX16mDZ4grLeHsCyzj6L9n9wFtlkzvAAHQ6TLp
OGnL9XktF1yDzP0GMsT2SjowOTzSkcmVJA3OEEnJjk31Ow/8kPVDO1z4tdExK2e8JAJG476X07Ih
1B7SuciPB4iJeEkPrKt+doKJm3jKkG3eN8MhEfraDGxmBIlv1oJh8LWA4dt5nlHmSEyNccTi3prH
qiR47H9v//8HXWx2Vye5sxHpPoScjUR/Oq+hm+XNa6LX5+sfwWzSK2faPG5J8cXh6YTzIjGLK2fM
24h67zivLgp+nLKjhMep1yhzSxSIsy9mloGluiekg4k/DiMpARYpdKQE13sBD6DAZ9xn4PydOnHW
NTUW+DNZw6g8kGE3i/81EhjGlScAjGUwqe21sIOHaoWgq9wED7E30IDQ1tl8YT5sfTf1N4HxN/6Y
YQTidrwcemrNZ0yB7LSsPJ11JXhreEaJVm/3Oy0W6sIdlmLfr4qFGo1GsWoJ+LytRdHic1W5EdJ6
anohVp4GNsVfsRfdJxXoq1CBX4bzzXigXRuo+KjqiyB3QSCPZY2fl8P/NtKjoAet/QuVr+XjRWvj
fSGaJgFSQaHWCdqQjUmB/8fJYA/7PIzEG2fUthqFMCpPmdHAkHHO+YfJYtRbUZh4m62Oe63BR0LB
x+iKjxim7lebVWbdD78mSKN6ASDYCpvv1avjdyKA+g+Gk8tlCaKEJPQs68bbFia1xpt4jBZsHBXi
MJDdlvfsg3BOiVFzdBBKGGs6zW5OZXvWV/fDw4u7/El/oGvIu1dHekikJluQTQBJHvaafDFqrp8u
xEa2pxE+p5FVcvyasLR8K1TWswqIjoa345V2nAQfZHzHuhvjbjIUzxRMn4wpnI85EZcnrYLq5k/s
ay1K+78KKmfv0K1+qmLhO54wtuROrz4EHGP4D+3kTgK0wC+f4LuyWzvc1SYn8IqxmT4XS2wjCKc/
mMhs1JEZ4A==
`protect end_protected

