

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qYvaWTl2dVn1UYauUm5HneGLdmTNfKYL2CALcG7YBWzuKWoXlk0Id+l1oLffyjtPstUkcnB5XMcQ
6NZs7JK9Og==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QYtaB7bKNbwxVddRWt78CWZ0keZknIQG6IQKSIZ5COH+hNdpgy+tCPVsEHq4IVZzTG1P1o7hP4Vk
F8E4xV3B+P4d4XumR2TMQt1O3p//18K5GFLVc+tXegTNm7nDlHWB2EseJW3Comce24tPY9JdBxY3
PqZ0pdNcJu1q3elLkyk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dcPEPRyvFmW4PpA4iDmUUiTH0W6w8Tp3x24VnlLzTcuDsG/S9IG3GcyE78eNrT/x0pAgwHhrMrSY
yZo9WE5CUIc2230lFJdjwqsu1GfylgdJvImjNnSRTPzlw78/vxcWd8GQIKrHyFhACpS0FlCWX80u
ir6wyey6yythPFMR7YL9alngEab5jqlcDLLq05xFb5xa60ZtUm6H8H/kSZM2WCTQ/2EYo9aRaoyP
YNJgznw4M4JlCmjNGCsEEMbnrUH5XC2MOkUpPSJ6HpAPhZTjHtmrQy0MjGpBzDrrGJZmxlIzL7x1
7fFFHCW51Ue16QvPlxZlJr0kCC3nTtDv9f7xsw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zhiiGh6iqBtYa8uvzkWpAts7vZ/x1/EV8yeLKnAXP52susoGuPOfmWMYojIG7BJlvNdJsqMcu4aO
YgpCERsfm5E2WNcFxUppU1uIOa+cnCBSZ6N5aebRGghJrQL1tUzWpRnQ2slMJ8Q+gRbsoc3N0qtc
A+A1dAH+z+hdTGoZBRY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lbE1QAVb48OwhlUCQuKav8khO5ghQAvoWa4EGI1wknY/PAoHSz/mN+mHHLZytFcumXquM7gAj5vW
FkPYXzAy7xSUZBC0WEUc0yo4Xa33jDRDxY7cxGlzHmyb1RsXl0duhVMcX5rDmM/+KiXLbAmtS7n6
pXv5Z5tj4x3AoNn90rxrYgdqN+pxQ1GZhPZPFZggV3JHWj2LJUr0U/7aGlgZSQCcdWV2V8ktlt4l
b9BA5BfHfgn1UuvjTl44uqXII+j7cWg72Zy7D/yYZ92M5Y7nPBoBrEiv0PrxnHLMrIv8+jN76TPm
TMiyhLNg8NAb1xNexvBsDmGJWQnxf5cukp8uDw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60368)
`protect data_block
a3kZZIyYP0rO6FMST7FqMFfVLc939MXq0/TPA7qcyf4F6wYZcR+SFgRYAEqOXqQMrgKMIIUCQwNy
O+fHya0Pc4N5/WoYBMeIARQWWNkUi+ew7DjGFe/CWW8JwhGCdwopGUTTh4dOyq4N9JBYTGnD2nO4
VAoBAbpg7oGL7NOAR3xAA1GRZO+dJa0mUImyVnfpxSq+ft6qP2aSNglpm/jyU0JomaguyXj+ajGQ
yxKyTsEhasWR7de2pfWssQtQOmIdDEnqekdX/lhmufMZy+buncLJF7WIjMqai1DwV6LzXK8dCD28
xeLbQb4j0Has8NWYnRk5JRg+8HTZ4k1QBW/WgPQcVXJn1qa/vMsf+/GlHYSnwPCVsfU3HJ3YHtPY
JHVFK79yHDUKCpkvOH0ZZ+YfQpUy2xx1VOFfftT+OwvP0h7uaBsbYMt8ySFFTdKpw5s08NMXrIOV
1FTNa9M7re6zyBpgK8yVJeQb8iXxfPDUzX4QhRk0TWPgxXrVuvD117OsylYyIOYMw/uQfoQsWmoC
KRdP4gLCF6d8oY+mmOl+LwsotE556ybrklSIl3FurneWY4gjyvKadZ1UQv/ytpCBdKpT8vAASXPY
bEt0XXQvgTQH1lFmLjAOC9h0Z2kAWFSki1VQJud6aQLVCNCCmUV1dermZxYHfbxMR2xCJw4PG4vk
gIgxJPgDkeIH+ZBXrc7q9U8wkyZckqRpHQj40Yq6gjIb6/riYiMzvzx4nrhMXcbg6mCXpVLXvoaF
Md+6R6+hV7jjvmNFx09p4zeACY62ghO5r+ea0AtX1U+XGhqVhbe9nTJadiNmMYCo8kDjO37e4wVb
VPzv9s3Uu2HnNekz/jDAkQCsl3oyEPaNxstRAu243jg1yF3OVqf3Vuh3aCdo2wAoHLI4j6aZH+DR
Y9zPwOhr4GOsg7T9aRHYTP0d6RscVgT4RZJRwEsLhfcGrLi/1I7lp400PXQFsUoYIRC9YXefCXHE
4aqV1ltSNlpT2NnC6ScWWgwT+bnp/yfhx5ImpLF0THHfOAuBmMRjhV7EL7vbD7duR0QoHpt8V2HB
5Hm81aCP6cDFhmydlGWVvtkWYSFeiQLM5WuUxX9L6eszu5XhWs/7bS9Pqhp53zVv8gUn40Z2kbI3
pQzfzM2e086ov9DfT819zBQAvIi5jgm7u8XW5ImBl247ws88YuIpOhpOSZWxviV5cQMDeafGDSr0
CxdscYx72nbJ7Y+1nBXr0QHKwFF2TLgt0zbPHtFoJ6PDjIPhJnjCseZMp5Sd7RKVLIUHRUpLEL+I
Qs/EKVUZzgzdPhQOYyvj8stu1oooW5CTw9xTavX0kByuXBx8JILbIitugaZdOw/ntVdWf7JjkjHw
jmSnzdUp4ZLpml7KTjp7ya2gEuzNJo3aFd6olmVrKOb8kpeOmw7JAeFQ2Fs+GWcHc/5oNn5IkJ1Q
P8b7K9ukza0MRxO0dM8fv9vpI8fLzmjV1xn8XJxuHcGSPiGb6F6WpJBR84ug0a/jaupTfJB3OPKV
culwheIFvez8aABfXqF8H69oPTgDEnwClCsS72ugyzV2O7x0n5n/Z4xByHwiDuAowSGTLSGL8gKG
fcn+fkkskbB0bsHOTIO43a0pV3UYPtcoFqfrKPCoX3C5zFOe7eR8FjedTJwb4fTdxQetvJXKkz3K
AWfUpuQI1t9P6zPitHzLW1FVor0euG7K+EtLoR9OzilZ2ppOuEJgVXWiyOf2cs+KxAgVZqdHCtOz
tWD0BIZAm6RWQKTE5zW6Gi39FqLC5BP2jGHp7T1WXame5pZNdXFQ/tjrUppG2JKvoj7PnzBHhsqd
lfDOZ2ddi9Xt/7mDeSC/bbLzO5Hz5g3tjzs5r+BhaCOpZ6BoZ+vBGShiNuq2sqCOL5Zh8ZjcyVpE
5qJjxtNl+ChJn0CXP7CT2gXtx7PxUU3EEXo8CP8P0oxApS5Iok5qjAGuKN7bj+JkPAxBlgzcp1Fm
khpn+C+iSlGLx8EpNHL4iC4R6l9jMotb/8NZE7kd2DWHr5lHKWtxeeBnCRCZ3PECfxgRJYYNMFJH
ogX83kXKPR2badJLN0HnlH/up1Kz6bkOyJEnJ+m11Ulc0/JIDTQHLP9hl2wIcq+rylNqHDwdzF/Y
QZXtI6QeKGIfnuf8dZukZMewp+VfDZkzd/CN9JI1fbct1O7ou/nPlqkBujzg4Uj41uVFVsWqjiVJ
574NivJxKzPE+BDTyq3r1Y36D/zCqK0JOaFgwEzLgHuynIEuTm0ypFPR79v3KPw/aEDmWZb4C3Cr
3p7kK2u7HduZ3U7OdlwDPToaeQaoHXQLvYoHy2UU7rz89bxtsmMaIfMDvbQYhjr3R0R4V/gJ5o2e
KJIUyV1DJUULQcsA0yLuuv30u8LWMjEIsKzhaFGxpWnNOiJR73w/inKg4YdxPkI6pByiOoKTqFjM
dYwjoZKwwFxTvPwL1FzRgRNX8uwg+AYNu8LAWE3d4fWOCbs3+ctRPU1qtgBW9PGlvvM+YG694TMx
7rfSQ2gUHPTFdpBFL2HeIQQjaPXIlmZ59ld87c53HgT+jzAg9AeaRlnjO9Ngb7H0BOCWRJxixsef
MLHSSVLRLbcL8BFn+spTLyJM1AgJ9D2P3C1dKO/NrNWRq/K4zOpkn4i/xYhElBXDUZLLEg0VQm8M
7npGdfiewFQsWAAK2rIXoOMfP5wTEp19+Q1g3vDZ2+od1Lbmucb4RLU87GxOxAThrBwgUbefMFmr
gv/C32zJmkxf7UXNmV9CjShNjYTzV1b9UZbvRBSzVTcPYf8GqrEaNxjDc8NmJCjI0B1HnwZMQpbb
JXjpq06MAttNEW+EOHElPj2CgKCZt6LOCu9WToWVqPHosOMIJlUOO9Muc5NNXC0Q3umNnSbbxQ8Y
iFavb//4kouL8hfGw02VM7NIfrq6GUEid/W7sMRJCoC6c23P8smDXPCVhOv5vCsDvZ8t3BCRv40k
p3eejPmkhNQqd6Pr1b3ycyNbAJ5/nXcxgRxoAxtU4320cmrLjaUa/nP65YUj8eNjCVCt8CoCCbsj
UzxaTgfY/13BN7GyPSSKgsjLTpZ1xLH88g9XFS4aTXM84GqH/KGxARAxtEiQsLD88ChHKeqPdKZG
vaKMBaKeijHKkSYUBcrLOg6SQ+Gygy8oxF6RkW/BZh0ngYwsSt0fnuoFJ5oCyGDCyb6QGgTkmp/D
FxdDaa7/sT6My75/gLLUZPRZZ/ZvUM+VeD7Tq0aNGB2UZyqEWxfGo0W5A7HFptfrsJWyo1LnDoqC
IXsRvdeWkjymGowaabb5bxZBsgyFjn7SDztzXy8i5PNnB9vVrJ+HuIvg/o+c/w5d5ErTfKJc/8Kw
1WJN0fbIgpIvsT5arOJMlRo4APYL49BPvPNnzmDYRQ1zw37qrZdOMl1JeP9A1WWSnNQdoyXwsNea
/TOC+FqFski1mYp9DRjV52uHEfre1qVMwilNyitqJBszUXtlG76Pw00s61OvFDP3D6s3O8wSb8tX
3mwdzeIwfkEUvlNCb/tez7E5h04xkpekPk741eVfDIFW1K4k86mLLnFgwO2PI2B2dQUorIrgTWTO
HUOv2lEc9JzURJIXy0Cx8OUao+AzW5hcwU013T8lSXPlA+71J6Jg5ZWVEXvC2QOyKQv/abK+LzFo
Q+GYIYWPmJS1J/sX6YqYr0kFO2Qn1BoRGr0OZ9V4U2XjqayxHwWwGLddKEcd7UgRjuZEKrcZ1GJ8
rYUx00PvIC8bZgKjSTSGFcYxSvo1leTBXN975Jp5xTO0YDJXeR8IGGG0tnCzRqDPKxFmwkn+7iHi
diNUQCMljEk3HxITxKOrpo5XtZH/T8Kpu4twShAVZtjjPfNLZB4plHDCo6/rTYfIs5pokRhStvNH
G+Vka+aRhxqPWCXmzFTP6TkMVSkOk0ED8pIqUDmxMKvV26q7rdPxp38A20E9xFD76H5EznLKCFQA
eSp1CaSDPwSh2LYzocKzyFI3WNaw3XfLyzrh6D5DE2DzmZvZjiJADKQooB0T7fjTEJjqj+pFPU55
CBngIOwnp7+B0qPHDdx3n8w/PwrR3JT3yYx57OMitF5OKz3jOZNUtLiTJEdH/t+uzMBqpNHwiZpY
zG3G4rV8c5YJ0XgTqq+4bmiYx4djRXLaBi29/7CyqPF028AL3gMV0IPgKq7+GiRPwoihgDQACrWo
cj5Fv1/FZoRc6BzTjHJOgtLWK8SzcbHGbwnw/Yn8D5hILfpQ6nNp78s4wF7NbdYXeN/s71IMsDWM
Lw9kYJA5Gjn7BD5CeeVZQYUN19hciRkeDKrSreM2kTphrzkE/+vY4mJwy04cxyn5tcS/Rossncn8
tMSwPiofaqVVdJkFbTP/vnhBddBM+io3PrgaxS+JzI29C2VD9Nc39BsSCoqnwcIxd9jkgjDp9pA9
pQCDF37g1uS9C5rmg52K+dRfXDtak8BKbIKUx/hScPXRbSprqjgNGgMLfpL2i7PRl8t9Vw1XXVc3
7wROQL/qbOjdFw/Vzk83Ni3Oh0TfmV3tS4cfqLp88tCaepxRvwp714uvvGGXRsh2yjImqvMplL7N
lFRvO54NA32PllqpG5ZdyM04+QC0SjqG5Cc2Owim45pEp0kYi/riBED1pE9f5IOYRA4VAS98ylKR
iHdNDdtmJjQIeLllC1qis/t+CntYElb8Hd4j5XjGjzy7TEDJiaCWzaB38wIyvyuCTe9R9YyATHZq
I9QYFri737MZjwhzoEJgOKElHqU+8jSaF6qGRw8HtIu4ZI4az5ki4EAk9y1cYIBtsj/oHbz5orPw
Vme6ii1xzoUXJHa9XYYpquFcpPgPpXU9yZQdLi9X8UIT9Gu5rr43vj9DwrmBZ6xCppZja7s2Ce31
yHTbaiwrmSj241By/5h9/znEp8lx6pMdTXCmaxfpXKdH5qyGbA4EsWJmC7AMU7x7ivR2ahDpfORn
H8WmhTmqD+/0kksoWn5sdpHFPEzH4Di3vGcsdEaEoOUVm0kHnlIaiz5KzlZfzIFzJTh3VPQlAsdm
KXy3hCgoSYzNPyPSuHpC6ykeDUErtI0KT673ggHGswEPgAoh1L3XVHmPOcvc04NaN/vagfWefses
RB2s0ZBbGB3ES09COozFXLrcXMxgrAXvxvI4aoVTy9soGPHrmPHXtMFnki4iDAxV90aHP1/j54Fk
d/C+tt/ozkVBtQGDciSjdnRciNzMKtYAB8jqJN/NDPxhreui9GT9Hf7iHRBTAqkEUsFnYC9i2vYD
ZVt1NGt1LfGx9U9ucDb21XFYC6jAj7IzfbTXfsFkfj/n2y5oiE/DHUdniBx11++ni6/GQURNcMTr
jX8Ew2m/gU0HIr8qLtTVJjDPAVhbzj+zDeZWdqbjpKo4S5zbROy62pkt1UGGBMuq0kpNrrgLsm/w
h1Ov0k9b92eQ0AMUjTdu6tPqQLTTIfMEcpWGT+x+OVNEhcRdmjWTk9kLhpX3Faqqpsi2WnUHGVc3
YSfzw9d4W8sB333NO0q2irosPwVj+RHOAyMT7yy4D4ud2j+8UreKARsbkso98LPMCdZE/rWxzjg5
4HyP+hEDzAg9uc2I7Fe9qi2jWEx2guuxWJXGT2SrWn0MoJbWi/tvWuZJ2nvWlMMpu9SU1xQQ0YKZ
S8zbeaVURNZmO9K9kd03Cd9nYUSpVuvwKIXLOKmCQDYFKD4hhUxF5/hjSxvp+TaxSm31Vce0mVLZ
YVkqsR84zjXQ8HrBslKQdTLVDcAO1MB7WV2GrBB5euGyyqFXSliBSOGiHz+vV+28FfdCGtS2RkfL
yvd3V4WhZ7YPYguzBa7+regv+h0GywsNYG48uCAbMfVSHBNSC+J3BLaaXpwRRFloxx43EJy6P6GU
gbGx8EfyI8JB7WncZCaCnzZjhB0DQp74bdOZ+Fk41HabH9gm5wyhYXwTnH8OTBVp7n60aBYfIpMG
9EgQyl2DGTVoHBMNt60t+sbp61yHrz6t56lEVdhRfnHZFmE3r8IABuMK3OmO/sYzTZBKQOC8EUpG
7EO6/4K4s+lNa0OF8EM0/FM976B7A6DaV8t7sWdZBBWki2HYFwTgNVuVfJxLuqaLTq3vxUaMTtYc
TdOY5pYN9Pw6YkBFNOy4z18rDcX2Ydh/9/1E4/Tzh3mWDasREMXS8GISjiElDCq9s/1PMqosnw9A
YgSHwGigjRFEFEbd7kSER113XWCb1SFV9w03Ct4OlAYJ2BarNUSw7SPIHfp172vq2jrVLlgPwr7M
EMHnM94FnAVnyvalp+vGhaon1jFPJwaaQB8ie7CDanyi1QchdrUx36esEeD0wZE8Ty7ggB6elYZk
qbwOFq3PXELuxdRfrpEtIYzpT24PAlsmFwG+YoWfMKp0UjfBlGOoemNkZhMJ1UW2fjJGvwQceQH9
maOjjBlE5VWBMQHYUjG3Wn3r1+sUoV+416FOakkVoBSPQFpmUK1qgVOobX/0JmJWYhROjyYSrMuG
MK8nEaWUx12TssMKP12VDOVi4U1LoosGv208TrBxEGU6B2sSZ40jy+2/pfe+ZezcOCU5njVOJYPc
6uQmzryUpVfX9QUzVsoWHrZ28xvVVclNpYl7hiX18Lr0ltw0dMyhbBhdMe2T6mgXSP5rl8NSsqGx
Zuyb8sOTd7wahbfvPkFs3LR7CX/REUGx4XTU7BFx6x81WAtIVYdqPYR4N6Ll+wsBlHcg1tGRMmBx
PXqhduYUG9lJtDMZo2QHFyGiW8NINKbp8QNQad5Eaq8/WrHEBgYFew+NIkjsHv+PHEwmfmgX7csY
bK7BVrqIQJSluQa+T85hwTtJoO9/7XUd06HHhNP/NyZxnwx1WznJjH+JuqSJ9/IZUxfgLgf3JM5Z
N7ICz4z6blKOOpABePspoSFzsu55Fsgkq3TR50KX3IBlL3oTgQbOc94IeXScoC/S3Geo+8To7KHH
CfKb6SEkW77iuY0ikxVngug1OvMb65zE5QpUDJP0rRnV4vkU0hRvCm+qjgp63TllnOoenn10Xi/A
6bec9J9tMk10RaItTrmiL+UgnEPYBQetzrhD30cULkg9HbLkbE7kK5/tSQm3uRA8LRqXFlBVN3sw
Kz5uGQANy/aZqzj+HIikRtECw6UOWNXsS8Hs6/67q2OXpusVyeCdv1ejIM2fc1fP8RVj8ZdlPICP
VhLto7SmOerPaVl43dwUeMTEwf7VsZhRIVfDeM8WlKrVA2ywk7A/AI9mMX9gwafLgo94f+VCON+q
SxJtBibqmqUBhPKWPFl0qV19/oKevV8q/hSHoC+lwW5dwIHc98wDA1ID79r/Qxg9oQo7iXDcTw0w
MwlsAdIvq0Blnw4Zv2yBiJVknEhoLbngIOV8dXKAQa9Hqs8L2lsK7w5gGkKxbtjpFo5mrzqtkFTd
s65C0mwcXGB2fjtPVrD2oC70ucD3tWf/XAupWB5bT5BgrKTx4Ush0Bfhfz5V3XC/eZYeQZCtP7Ds
I6lfa7N5Y7DMzMtqiYfWIKNMH4RCmTpSMplMp5Lmwnamg+tYm5b4GxChqqdKbrtdcfaXCwE0K9Sj
sNq1bXMD730DqQOvqmqGOaenALVe+M8gdxGEcGS2hDNdlBp//pnITNGLDi27umXrEI0D5j2uJCXT
f75Qs2llCzcnW6Kzrj3Wos9n0jJZJ2ew+qB1eIUKrbVwzkJq5If7BhfaWjqzbu2hI0SbYhFGC+Xa
FzBgWGwpPOu1a1OVMfJbemzR/Zg10xUP57ZNG/HZrWt2WVTbLeSLY3FRaxApQU3Q8qn0mDPVApaT
mcmbtZSKUWwZSXAVyPr8j0wk+BGEj79mtwe+y3/CeJfI50OB1qaAUZc/rBFvCeCtl474NmKYPtPP
ahXGb3X1/cNWysTDnBAwpghnd6/U2zTjcjP2/zu+y/RCDa4fTXx/8Y08r38FhiYPdREzPZdp7h8n
iR2MII9nfSK6BmCKfodeBHSJO+GnEMJmjzhZ5bzmW7t0G/kNkyKuY5IRFizm7GRtkaA0JekDDBOk
7o+5UcSqKT2nnkDf8xcRX+J3frOEgipG9S8tlSJJgpsWH+78/4676YbRYdk5tOo/ctDELX5YKYWh
Rymkmx3p7I8QoqRhhlsS47sD1MpXjmitnripmp+lO2Zb3qSZfHVVOJpgNjV5EXor3k1Z6n1Nk96A
ELmVCLbYKky1eHhDVGOba2QJ57Wbgap3tN48krjO1Hdm6Yjffi0ws74n5zKjfaik7E7Su8Umay5x
iIQ4+YYe/0VLDrpyfiHXw2hRDxoUg/zCKD0MUPobpBusciQoALFxhA1fhT3xPnWVP3wZlHHdRr1M
v1aKLkeGIUHxDZAxCf37HHqCgdaCxayF/bE9X1fpDYhA4pSdP0/SSupNcPKHjupcrlOQsa0It6ku
gc8hPdUSDzhc3xqEwFGL3gERy1I1kYf7XQCSzdC6N0eA9BYKZEOJ0kqdx+kBOuzOFmDgQ+7RuOHp
lsm8ukBiof+PJOhH2HesiCbYyWmjoiM3G0Xz8CKbG5hA6t4Vih4z8iHwCkvukLZPJpkagTPIbTfd
T1ziCYEXxOX3hDbr4Q3Y2mJe1YuXNLI6WYV1aiyP9wlFnMhl0BMLmy7CwfTK/HMijaFWFzl7kmMm
1qkE7qw2TSW8hNAEqqFpjuxARwgA57fHuNLJ66I3JFIn9J1usGif2fpCqdBTXsQx8QJD+xxfnQJs
nZbgoD8/iab/OJniDSVU+W6IfhCixV8hUSq3r/bqRveu6/WB/LdJzpP0e7FIc8aTFuBTPbX2RDH1
OFCa0utyZTEJ0l2MJMGfnBCCVUjt3yJ0bO45l/eXcg47DsqQIKIcqGfrGxrQHaSGyhp+Axe2svpY
h92aBPzD3tQmhQd0dJWw5tiJafeNC1RXElnpft2bYCzqq7zHFzuk0Uj8TfdSClmSUXOzTgSciLM0
0ciAtWdXBiF1yVPBuOQq+nPseQkEdDAzf8InJelApwLrs7DMNpYNkflDXFSnQ+gD3uqVsJjtQ82J
DkTvds+u4tGYFfownjWx7Ngl4lvqRcYy0OrenwvKz2tahN5Zts52vmMLwIBmH8H27m0ATNkoTnRr
Uq6f/nrs+wBw6kP2xzS9pFW8rB3ABNYKjdglp48hXd17qnZ7PadioHT3yJme/5kOxQS4CGfMDfsU
kxg5sELDeSEaZwIZoMs2mpNk2YNiS7LceiT0xw4pcTKYbbG3nXSip1fAtad3S56eWCn597qvb+9F
SSEzaZ/RojHBqNbNJX/PrqpAFBHnOiIqCuDqrf/WylWpO5w9d7gwlsP0jvY1vIJwN48mUcwPpIaN
KMkNG74Fp3n3XIgAufrFLO1IU5jN1jpVWBaCmlINqRMdB8owfCJMNZk22S+5GMgHUEaNkklkylKD
iqjUejlZR0y8Um6QFHnWWln8Em5+3meMzsbwCtDJSaharo7FWdj6ZrQR89K5slb2Tl7sf4ob8oj2
Fc+pjF5Q09qqH4ENi8O8YI/GkQIu/DKqrA0S8gtMl0PgJ5vrk4BjFBNF6Mwlf5cwjz6SvKaoAuWn
lwN7awJkHdu3XYSPfNiDHfyw1Xpnt8DajsXk43qYbCpyOecajWyAx5hOXdsGLsu3VijCqAw9XM6E
vFGCalhmQ/xxQX+Taw70he0Y9KVaRrz8eylRUNCVdiWhyTgL6cEVYL1d9OygCZsrO1sYRItdtM1k
HJfIio1+U6PsOtXvq90WIx6zb7mr1Z07sOw+TeEGGm34Vo3ia5LsI0+2V8YGQjnYmuN/xrSRXu5U
tcS0kZMr1qk/cZN5EbOlpUlTCzvppVaZpYhJ/ZYTiXG9vE9BDSTmxkkEUqyK3AsluKdAacGQ1XzJ
dFAoABcMt+AJpFSfD9mGjv5nBeFMXjiHEGYGrYzY/3tLnQkf9om4isgt2KB/AGsot2stDoTOF0aG
14dVTJu+FOWI4k28G9k7c6JDVW2Ll2WyKY6O6cHCFq7RfOjLQjh9H5XT2leYq8hovRiskIjJQljP
Ni0/adM0L34IeCNwI+EzB9TRtAhF2M7WsfHFVCbk4T3lA/GsEsk555PBnW7ShREs7pibf+8CA4m/
luJimFap2YkBfk0jF7z4wYKArM+OIAZQNqc9Dzpeqsyk60OslGainnT1XkvAqfombHNoayBMwMk8
88+Rdm0CDOsMu0K10rFQ1i9T2UM+/k+9UAdP53QwjwhuxsQOEDGrDhF4Q4nFxQEtG+xVhEXf+KRq
xtCHSGkXaGvtsK4Nc3ZQCMAgvnWki83KcgqLIg201FihdfO1Aw6XfI4HBlHMuFPvYQO8LZ2uD0Gg
yT9KEi/aSkGWHxLUqdpJbcFKVvJHSvO+KtvBDbAq5Oe5JpMmF9ofTNqbynCsWo5nF1X+lkWCz/65
qEw4zNpm0d34u9C4JKzDJ4Blq44aOp3BGsqXzj0YMaIrXEsBjHCtx2uWhl2+R3qnUpkZ1gsKRRWG
Kz/r+bSSMz3v/F0e1IOg4IfgNLb5kfEgdEkilmM13wPa2jeTsmgez6AW7Mgmab++3Pmp8s5AL73B
rabyWWuiPFH7GvK2sqghx2Nnd2iJUH/eXUg/UJzUKPkJctcUkfmQCTW41bQiQPniY7IN13fH53IX
akSnF789J3cKSJ0XZtFZhn3ZUbI/IflTXSvvCS9330oIZmobxivsPL5bI8BCviRQmOy+Ky/dyfov
9//yIeUVDyf4AzgvGM7gDBfJLo+CsLwrajGtyfLYRwlg8zXlVPC3ebSGF7aYPWwAEX4PKp7QU4vQ
HY4qxW0UY9TIJbilbYD9UL2K62p0qKu5tbEnTyujmhjN00PMqLARe2zoPQyiyWoCU4vY4QqsOP/N
5wH5kANFC7pUjIsxAn82Fgx1WbgiYIR7OJM5Z2qFblUCideCt+exB0NtCNC3xAnDaaxSyUcuKWus
dzRIio2qvxDcLp1v3hAgj9Vtqb9DFWUGSetdmSqDcedu5HokpWBj3bOuAcrpTPJtSJ9PPdAphBMs
FsbvrqqJfC/bZJCchXFxhHdF21whtr2xAc9cU+MjGAtShvETtApLmdCR1hyfdd5+KkOA5sZctvrR
aky8gfqTIzwMI1GCz2tzEmPEqOELwp6cO7R3vfSQGuM5SOr08jDwks+yyblc1pI+ekbA0wN78UDR
oerJuvHjyyB8EtEJFgtSXzlEfSB+Squ1ewjF/au1TQppmQJHHR5ujPkVi8+eK6hl8ET9VZFl7dFd
/NQKAFgHbzK0zQ+ZJglHfjYUqXSl+Xb/1ITIQkSwdfz/WE6E+wA3gUso97A/QN7tpFZmoqRQ6sPe
Zr2gupOvp8ioRXucVyYo4ebsFpfL/WFRCeFYYwyGNiCSiDi0L05lrcKT/3RY8IhHIjBCDpB7xBcf
ft95RuOOtxkVcI4ur92H/VtF0zJnvDjmL2WD+pCuZ8rWBAwFMkZRXu8gJVTxwaO+tm8GMoxj95aU
CsXRmQ3274990zOGZvRkK4A1sd0hJHv18WXax8ewOUapaEx66S+UdmUuLk7h46ejBS7mjIEfnJd4
XRjawa/+JSlSeUvxLbHfeHxhYY5EgSClm5UocYWbsmOLtpf64YrzQ1NOWXGMtD8ZnIzMEIS69cdA
EsHgIONoyl1BAkPA2zmkF+Afr0afRz/kYjLlwvw6SpvhK6F301rsTI00Tu/pLBbiRF6Pkohe/el3
/LVU2JW3MBNHSvUGt+xw22E9yWu3czM2xPgJg3+bEnDKvQH6k3Br7UD4B3hKN4zBNdEZDGenK++j
iWIkyRpGx7n/VKr1DmF36mVEH33eyZk7pW2ZXidBo0rP5hSlPcjnosVs5y8YsXd/Ik4OKGpMvYss
VkCXNaBue/c261EV5FQugyjMmtRZjDx81/OFy2Qev2TSHeNcgqdOWK9uzF90XMD/+oMKWkgeiMN4
ionW5NcM7NHm9Pu2aT/sYZv/2hUz4MO8hEJrCsv5+teiAwA5TARieGpu7rw27jFCKsUzAANm9DYM
6puxinR6TWe6ubrKv2cpNTMYcpoIi6NYTXhuq9UXv61VZpbmpqSrYakevuO5m6RviWqD8DLHrHcH
INHlklicbkERYzJLzSQRDReL29LDpRWEewjDBPEPrEPhQnBIlk/WCqCpODmLPoz769IyXdQeap5f
lm1eZX4DUqa6VSuJ+SIjSoscmDY5c/iz/IuRoIKlu+92kF3bD7PelwtO+GkPs9r2JsA+xD1Wi0Eh
Cs4TEEZnzmHrt8TdxHQjHjnY0kH8Igyu4gGH1R3o43o+hWyVKBbF5QJXFDPpeQTDfeJLJngBNoux
iWxvY6MlfBazaltcjT0xlRah/Gfr2AL9VCI2FBWyQKGSVEaSK7qn4Cmxx4RbWBR2hU1KbonvIGxm
O1P7EXUtOnz9O4+66PrICczzRmWb9RwvJa91Z/TAPd/sNl0qE90dRq6Xv5+xQ+iIjS/IyP5RklCq
oIeinSLfl1EBgat3B6+yO17W5TwtxEfOwtRzRFPt4DkPOPefLa8YP7y9liAZm3A6qNZKhlX0wsec
ucod5InwWdunqg4y14UEvqoCy+AI2OBcedqTU/aJlm4fFr8XkQUzdRuTH6pKiIkXMMAWuEanlTWo
OIPsCr9oNB7ucZYwikAJmWybwsGZ9YPMAyPH0XmJCSY/qcf/gho5qQaGTAj0EmQ12sPePaNCDTnJ
HnVKroShgjc+rjBZ57NtqqucUGFcprqQQ+QrFY9zLM+rDiY8unEYElruRk/HVmBk69T6DUZJM8Ug
fyLCvivJwlGu/wcwAWs3GBRXBjzYlVBt82PWym/6AuZcIC2n3U+Nk5qE2nOLICejaWT86k3e75au
ElKuLo0lNNcMb5atiKO2msNKb4Om+9PTqHJdoNqraBUXCNnuGu35DsYZhgIOFSjto5yXu2MxG4Dx
ETSV0SVvdNrDhwFTogPHmq5DXWCQfIPltrhHsd3ulfIbecfnoC6WT9C8NVZY5RJoABtLj9sL2YR6
gUMANYgtcRNJuh3bv3oVY90FH6W0ghwoa5TIy4LM26NSmWvaF3lYi02Ys4TprId2LNcNA/+wpTtX
OfmxXXqlL5IS1LrfhqEDhLy+NyG0qozCNVrBMdY5GKjgLJUlheWlNWmDfjghgS2XgI2xQl9WPqha
NLAVKSyuUpsuaQEdvmYFMuhIRrok3DxjuYFp+ov5NOfpMDp+Tq/IVjBOOQpjF3or9DzDMpnINm8l
8zd2XKCfqPMiiV1MoNnSWd0BMq5F6mOerlTnc/OtXYMtjtTdSFtmCR/NolUq03j4jzqacPY7oRZ7
feYZWI+tpMxrza0qzXRdCvJZWYjz/Q/3VpfGzFJKqBNvduEAM2U70UIRH3BOQfo3EHLxJaqBj7y3
Fd6wDD11A18guBFGOy6o6DeJr5MoeOWJHzIo6w09hyQNx+bRbWcGzuZQvHTeOfmIiS5rqNnwREc4
mgqwIXBb6uyuLs3I01q8qcjsTi7ag4Sk4PnHTknErcI/yhFw+1QFywmdEqaGDV3lodEh5+dbZz+F
LelshpNHSfp8db3bFYCE0isr1CAMmk4GkUQvZdzpnxGNDZONsTzy9ZEz0pKo+1AMKvE5jHuTKmAI
mN1UjIBmvB0bYhzlwJp5ii2V/DC4lUVHPCa9fZFtV6q5IXf6GDCY7ZgUEtBQSHviuhw6XPpaSFm7
dVMVfUS3M6b4Ew6CbeS+N0qy9lFgr2QRGWn0RYihGKTuycjBfJ7qHU9rCoE5fkNWVUvydrBP86pq
/VMDxK794c219K/S2yOEPSMbUiR8ySiUDYcKiOg5Q8JbtXeOYQJi08lQ4ZJLbZZMDg7de2E393zn
8XCilzcBu4IlO1WIFN2RFxKSN1MXHyXgjjcDsfWwiio6DrXm0+8C0J/nDd1jdKAVmSNLc2xLawMS
3cewaEJmxHNsvfD9yRQ6wx118Gm8+e5PpbeCWkDUP/teHw1sjBqzO9wZuS3pZoA9nZUi+nhgz8Ew
UL9p2/TELD2wI2o7HspAtuNkmFZBq/Ye/0GXPBkp619vMlrpYGYA36YP6hwXbiCl+/4Wd0DPBU+D
DNkj09MVX/WA61gNkB4nosJp6T3FR3En2FA15VTzhZ97G+G9T6u0T1zGWx2gYEKS22AaiIACFbfg
oCZVvjbIcvM7uduH12kV56htQo5VbrUrOafwoyA19Bl1fuNg4hGzCD+67j/MTZNUp2DGHejsGsyO
LIU2nYQtWZ6R0UWvSEzqkjsiw9sob15CQpDUNaaVihI7Bd9oXnMosxQKJJFAr1c5adURH5PRn//v
pgxPKx8yZebZgIlZbInozRjKgN+RcwaWJcOnusqH8taOrdCkX7NsyFfu6f2lmhncW12UKNIX9xtz
CH5xBPpNOo4MWDEE+caLdRdK9n1vNdF/Stn40+ZLpiHH/7RzQPo3L1SfAUgQcZhHDfQeKW8dcUm7
0ctAE+0A2VADJB5WoqAuy5jEuZn5+pR0xkXnELuJdFTEJMieiQLeBhuiAeqyXCC0KSslhgWvKbjP
/2wbrP+p8AsJIcbO9NI5w+WUilUTFb9wh09XcXcPLmWUJUiZ21YAjJq99VRjCeqtNl31nIyWVf/P
OYmGq90EGCi7cRBnkJ4f1DpTOKYIwhGLl60ZIDa0nwfQobRwdHHkTazyBsTw5Pry1rLtZVjfl8QJ
5taQrxNubQeWlI8yqtmBTnOkJDK1PfZ+HiQe3UzV7kUF5bnmvNXfkftYleeEvp/c9YBTNb4fmug7
9U7gpX5y0FDawMZBS4ksmvr+Lw6giJA8FEwTdEDQJGI0G0fhRPkdJP25AvF8uMOfL5stE5JlvGwN
hlkR4EMdeU3PnjTrAAwsWDM9UAvJfdJKxSZv8/wM+n5zEUB+t5BTxKoYjQS+UBaaA/Awckq3VgD7
yf5B28kLkMkAHJc61r3TEv/MvL5PfcQcYP5Bu8A41hFS6n7huA9VuInRFN/CX95Jn/8eWmSZmKeO
gVO3FI+T5BkqEhHvNrSSXa2+4/V3T+X9+Gs+rsH+I3DZK8Br8vpvT34Bjecn1m/uzWu9HL1zjSkF
deTMtA6s2XftWMgBsV4H5lIEmX+YNfR2R/n4B/y90ZbLR62VVaGHViuOGlhRbn5LN4KsmeY4ngLI
X8Obb/MLuFPV/Fc0l6EeXY8TJHKuQxhf5IhEeM6VTFKof7I2hCkx3yPQZ3Ig1/3cIuTkdzD+SkET
a9/nmYluMB0DVBU2/rR1/AI/6hGoXyslu9PXBiLf/66kEaZDx5v01K3owqJyzHggsiu/QSEqjFmd
R1B0mkiW6KsfGVFKBW8H0+T6kDOYaSkqM4gD+aUG7sQBd+VT/8Eev5e+V5Ww/w0WW3GZ3BALnKnU
Se9O6kN0EBWtlk2fANjfOiefSCHDQv8p7lxwCcEC4Gn5N1yrOU3trBeH7N0dGijqKtmr+HFvIEqh
9RjyhtwZjohcwYztcoizUL5vjlVJzTc1HV4GARgtT+uCXlCwWFrnHcfdFHIiW+rRq61R8G59eXUD
C6WKLR1F20FiplCwfqoaTq8ec/Fu8ETj6KRSd59Vc3IIbQP9TMqoCQ8E0BVVtTd+q+3qOEyhtBDP
wSEunORLrgF+yuOaKfDckKpRRys0/gtAN1py9WZ0BxjIzoLLuLYtOUT227E9LH4osOnH/D4rNGOo
Cg1FInIxPgB9v9qdlKvWmWNSd6+sNaPJfjUDN2Yc2ZH60BJ2zJ4ePI1qADdVcg6lizqZl7a6V6c4
4QxBOGscLBEY/yTni2tM7rA86BsEkwKVnr5ywSoKIZMro/x3y7P+MHuvxYorEnQuRRRrzLmVoK6a
yAeld4TeFDsEqZMm8ubmr13c8t41o7WTNe8fBLDB4KZ7mybEvVhcnDAq6BHy6hslcFEpOA0/UHGb
vtC91as/u0WAKGVS90h2ZV0gcUAF82NIeu964la+6YYl+KUIvDR53+DkdUqMyaIgJ2CYAEuM17eq
ec6aACf4nVWelWv9ROK41FeapqhP+ZFyO0oFz2QonEhYA+Ie7MjEfhWPNeBQI14aMl6Xqzf9BXZ/
oFb/kk0pDbZjwNbxbdey1b3F4K46eZTENUWeaSaqFFPd98L2uugUofyZJPEy7p4NFPvN/dJ/m3id
vjjsF4LMf4Tbb9L04KbMELmOvfuTB0wnUBz9pcpDQUxCXs7YhBu18wa5fQoJwgJdthbtHJrU9sKx
XcmMORqoaYJ52zgAH//ugA97qe0OqbEs4mlEdKsTjwCI973TE/7lbT96WxIxwODqJz7QnosSb3el
NtDlaHsf1pbP7bjoKcHXCuXn4RTYymMay+n+xFyy/Waf2uphdMeZadNFF2io5NbxzM2xdRI/Fv9b
hTcO+anZm76RhFPFFLkPSbt8jlvcUsOJf5LYY5vvoowjgdSiYbs7aP7WQHMqEg/eDia0+C9Wrdas
MCvWluxJC6PhMdhI/3ymYnWJMuj/f/BynL6zaqrk1x0vGZ5fLH7QS32Mo3YeY8SZS72prtcultZF
6BFcRLCVpTmBmHu9aFuVHEPiNzSnQHqv0RnHgLGoEnSAZHI0o+eQVKbnPidJ/63leYVdubYunNmn
dupEbIp2lQjL7XcngGrpWQCuhYB6EGxiRSflCRXD0sS5ofJvd9h5lGlDBHDVUHIwh0vnfeQQKSxS
/r6N+tLTSB0jiAPjfhiAHPKwxRAs47Q5j/1c9h+JEJIMhdjfrfSAzYAe6kQt/vu9QEV+McE0VV78
ufyThKeZvKJJzVyvxPhw9lMTXQBuam7uE+5XZinrp59SbvCZ9tDh/0ElIR5kyinFEZT8l7xrQH0H
rc3KDClsYNvKAd3PV0msAKPH/PZY3HUi/R7DnGW5QTordoAS0aDHNUqBm5KkRXVJc3iXz7LcdU6I
X/xglLZcFoyFSP7ftJNch13R3734I+avv2uE5D1ucQ07DkJP7VVUTaF7S4td39H7Ur3ZjHRPnzCp
Bc2FS1/ZZQa4QOVgRIpLYnJaJsiNylaiqf1rd1WVB2IgPyAOOCEkKGJRQtbBLHrcqiPfraM6vr4r
kbNl3QTHHR07vEo5JG3g70MY6SOtmgCI69HyRSXuPc6BKA0qAxJ1Dup+dB+faNwOEWFU4kR9iacZ
b72Tm2eXYBRseCm4JnIryURQCZ2S9vq5Xi89Hl6I5gRU5KA6sUj9vYkNZrpGO29ygP0/xW2Y8ju0
bVbUbsm5ItLX4tgJUKduhIMNpkBBiztvbPf2omBrCOwKU2qKNRtSBc0RO0dIjUQgPyfwc3s5DcHa
aR2o1UZGFWBuBGuFNu6m65yaAOVPohiHQ/OH1s/aN4NJ1vf6FEbpYVZl+amj4ntD8MuPshBBr0U1
9T6rHod9R77N7b/40FwHIbq9kl60UdYD1dX9RT1pWtMxOImvm9EVCw/TY1RtTvnP9gScszUvsWpl
XG4wpicSZlrGNAo8g/WIyYe3GSbJV/43ap06z75KJ31ZOxeuCr+h6PvaNeDphSaf+DS1p94eE8zG
CHhfLOk07O+0UNm+VX5mdXN0DL+VAjrMoTMjzMoFGv0WhvzbtkvsBn6bRb4bK09t6hgvcD3fXgaL
iDlNWpwWmNMO5onctjcR2OeVpldZnENN0geJkpGQZDiCyBiyOP1qgBRBe6G/6467B5smr0k9epcN
lgZW8u+jkFXC43TAJm8vuonftVzl2Kp3Niu7eQ+377ETDo21KrH4NDEQ5oSf7kzxKMAjsNre0su8
N9ncADC+yL317/wHqOfdw1A+rojoBDuCDg/kMmbvUFyFu8w4d0Lv1lsiJLKmUMEyBG3a3P++ndPF
2FLWJUkxg3pMPCOm2edzYTcj2MjNzzBhTUIDli8pXbk+tlQBt5yVpaq9A4tDhrTgJkxOjLGSbWWA
qtajCGI0K01XYe2kwXfuU2+SK+Y2LWtc6knK4pHxtlqWUZ61kmC+d30NUynRm12wqqNU7MXwK9ma
XRdGR/gLk61+So7CmdBlhr19m4xsvOjeIsUZUENncx9ARy07O7ZXjKPHY7aWVPq9ke0NKHBcR+sA
tn5oXtxvVMFZVW2oOvmvwDluqygyvisgJY/iaXssLNWyRTi+6r2wTabgMmQqsylSyLj9SvzPqvLW
Cy1yiqixBRUdqMrQynCH460kjW0b/RjIeury0YNPEcxRwJQEgW8TQ1QSkKhP+HnmaTUrvos8OW9D
pg798c7nzeXd6Psv1+vnYDr3nEiyTIClFP9aA1MPzjoOiyAzt/XrCGkyR7gYtFYrywdqx+M8p//+
UJYvgQBiggt6W/ABuNd0EMsEp4A5XbBGdYk5iXF37xhLeQ4y4QV8OgJFp+YSO2LyIs605kzuotKF
JB29r1E9besA1Kptz5bwYLouQKmv72f3gO+fTqshiV/1i84WqnyEUaN/uGIaEPpWo95/6G8swSMQ
2uD3O1Md/7a61/sw674PBG9jJ1MOr6X0XNTCVIYEfCa89XQLktB9f8HRaJPFpY0f9vQnHbKV9eCi
7FYvMQOsGQTU7HSlRFaiBKfPlzStr3JN2N9tEBK7gnhkOwsdTAJXfqyU7WSjfOn/CkJygGP87CFz
wqLj0bgpJJ6gfFMjL87Iyya81eaBG2gwh7PAyRVt5RbV28qcBQnPKzYTJ9AmMk1u6rX1vBANrcoF
9mdDI8QwXXgSk9ej0ps3ECc9Y5IOQ0wRi7S+d4r7Epay/XYttUZgABIFz+6X1Ouh1vjUTJdFarwu
MowCQ5RMSuFm2i1yyteNXI2ypy6B/Yz5At/mTDaUeLAiEgC+e13lnIOFDe5/VA2ZVXaQDwEUFUHe
Y6o4OdOltUDv+ugPb6mEGxjGy79D6UpVFk9kZfuczG6oUi7al4J/69NTxninkZz7NFBKHwTR+Hoo
FfSzlZ+1s/tECHGyR/mGF8ZpeHC3ARzPcD0DBqCMJLsMpmZBA2Xt9kN8UmlSGJXTYqZO56ioPdoD
qoTowFBVw6p6mIY76sdVrCzDEw1dmlCPU6zf772sPphlylyCNC895Cck0KnWuCi+mKOKvc4xqDCd
b6uetPGxS75YcDWIZGtsQP6Hni1/cX/bbsW0Ty8bgyDyJPwYr4j7r/a5ivWx7T1vNTYejH3yXSyh
RYHZ2QcjuXPuXFqDiC6XgzD747KluTwBGDaRJUkff3rTVlTB1Bl3NDdPCs+CRuY9aVQnNIfOJAoj
ls8ZW6m6oMLMs9YoLlm7dl8xMSzm1IVodWgE57vL24qY3lSqh/enIjeagTMFLLlU+a+ZzoXA1b+n
272iPFzYFeuo1wFyTpU1FBjtGrhQ26MK0mbspdz8hMu0V4R0emN7CcWqQI3rqGnKcKqCln5vleDc
aRN1+lhbFCNRonbUG/dTTt8Wyk9WwZTPKYoY/QuRgc085hqECs9yiLIVCLXPtLEJ7FUYEfQya2AB
j9Qtcc0V7EM4ERQVgehmWINbZkYjRMqVOASi+WcFtqt2KHTmNB0uDikc7e/C+SnGuXaKQUv42s1g
2X8QMFtaXgVGh6ul5h9SOd0nHJ52FaIs9ma9QFvmWMRFXgAYjTpwKHaZYEQC1eajJM4Eb8GH+vJh
d1EvrI9WhTkNk0YIBH9AcDbFzr0/yt6oBS918krxjTRdFyzVMX879zsoy4WkbEfvDIISmNEGowb+
J1XNYIDYe66PYB/fxT5pjImS35luq2DOIyp938yuiOYV5bbz51WVaxxiXuyx0+iY1gNV/mKjzkq1
Uoi0slS7YYn5LlBH6evU1jjcHnWDFWXEhchETIM24srnnp8wQsHfnyZ1ioe+sjA0yOqXjlx1HQ2e
+peDkMxrdyf866JW8miWrfGgn/78XQ+3a3523xtrtAvoEAN8+PyKFU5bZ8Dy6vUMncCYIWvHWpeO
E2bRCWMfUpRu4N6mFOY2uax2GVDzQErW/maKd1v4zZSs2UriU9sdODkzPGW+s7WsnJ4R156nRm4N
p0kqWFp0D7CugMaBZMbZD32I1vrPxRuHyPADkdJXqi94l70IBHsP4bW7qAk+9NTk+asLBPtK9fXr
SZKkxV2OWYfxu1TrCYb29SqI5RfPfaBuLqBI+wD1eobovZKiIXEg57RLd8rYmJgxe5VxHEctelH+
lKtHsqNVtZLry+p25yZ/7at8PNIf6VdtjgGsG0CN/PqJoBy8Hc7bohvP+3WwIw4IqkJocZ+SE8qE
OpmOI9F4JebwKqZy0GcSR2/PGJ4bwgiFpEorov1HKcKvLGyEagm/2y7s07XJQvZSywsOVx1rPi5j
5JZbrBa89WwzdY3k8pSNabMvA+VzS/Qg2oCPIhG3dhR8q0vxIW2OLTJZAr2yIur3TX+QZXhL+2Qp
wS0f0xHJ2G4Q9dqf3acmDqxa5gro8NLq8YFwTlL3+CbUkB06YNBVOw4kttBUOrM/EM9xhFuWPz7A
yexCENAl/3XUXTQBi3ec1vj7fPLzvzD1rRxBjFfY7hlmfC6edmIMqIadgSGeIQbw8Ng3/pX06Rqy
7xUQmZ5d741Rq+Q00SNQJWPqk+vVkMvkUqXu9UpFWZ6SsXn/GOBIzxXROoe2szHVGwRs5ZM4hcbn
2yOKu89SX7e65HQ2tJzzSvqKjai7TbOdUrbHx3gM24qsGdB9l7iySY8HgDgBkHtuupWMgZyMrjLI
yc7NGBreBBxTGoGAXaCS5kpzxVI2ldAgwbaSvuEU2+gl1UB9hezl8Qt3GsZOJkleg0sn9mUJAA5X
yICB8uI3eE+brmbUABMqONXqO/Tg8JVp58aiyxKnIjtdv4v22hQf9/PtJIPJzbx2c2fzgIVNLZ66
z2zFfjj+F/HiyRl202+yZ06yw/b8RB3QNEAFB8Dktc1R1JLGuEG/+dDyP5etu/O+5nv4n3GrrfCE
bXmLK/z9cdu7B2ilE7SFWQvsu64s2IU1qpLXO8l1n+2rqg+aMWiUwkdb6uKiK5EEA4m9uWKXxnAf
XGlgM4w3qkvY2FZvunfd1iPjgSJBRHW9daKU8XXt8rkiCn2HGBOQsu1Cf0zWytwlFdqB3DLIILB8
82zopBRqb1L3Y91o39xD3af4z24yehRVSSNAodZA8QnWeyXO0t8kAKp0JcESIZErnKgnlha5U6CP
YyBl48d7laNRmcT6TwLTFsNt8hKTQ6jCYa2U5IQ8W9e1KC8l9ygmacCNwTkC2Rtpq/DkzPrE01yT
DWuEdCrkZhIdonRWNusn7JgZKHViHJxFMUnqkEvSKjsHXqd+pYuWbyv6ojGH8Ve8OO7GmhPtlgsC
5qeqy5cJXlepHVZRw+he1eM17WEZMMn3Xt1Vm4Nw9Vi0+Y6SqQY9fr5QXMjQ65pmSIL6luRGWEsd
NGU8YSAQhA39BCVajPhAK3LeVU7n3JTRMIHGC+luJpmEG4FVIhW0UXyzZmf09r/mCNdwcagUH7P1
tQMcwpBbzEzyILe4NI9vNTwX41ddFL/Wyns4zYuOm/fFgjdr8BCBQk6dC+/PXVU3tSi0XXP0u71i
Es/kyM5x4abU4QL/z6rLmwDTEKNJkr8rKOzJoCeD7NHQj+lokGEVMeT3oCMRRHt0eCVZS16k1oo5
WMc5IXN93p2uWvthaz76+ZbLXjZVxVm72Ffdemtxt8ntLAhFaa2KxOrbVp3b0eus7cuPpN0jzsde
K5CUJ6fvLeuihbgPwUTKDKo2H3WKMmGgV7+bHj9A7ZNXnhPtk7BZdzSN1dOnsW63+K5apT65iO/B
gn+wK1WE78QJMrKQzvUR9pXsexSDzN1UhwYpYRPhzSw5sRyra9WnVEGf1r9nxR/HJOCgkLlrBMN5
V2mU8wZONb6o3f6/xKlOK1LOyij963PEBcQyYhY8FKcOfEWF8QkBvUz6N7nk1ftbE6/iWE7t9GMX
dip+DThBTE6ZDwZyPv4LfQ5xI2dx7mvrMEmXHm5jZOMob2YtMh5Ojueac+PBpIv4VsFCoQpE6O3c
/1LrxJIvwHV/2UjIRT5z45tWWDdAmQmSEh0c2Fw4bJaJrA0X3HMpfJvOigunmWeYWSlnZt7csUbT
M3xyFg+0P5kM0dZ+lEDjXRT4V2EQ+cjgcA0REZG85+1pmV2EzxT29hs8opLZKzKgl3ZYqOPcz1jP
n4XvssnzZ7Mqp9vM/9j6F8CBv4FtYASyQLbcHWvYBpHSNQQUNkb0m9JRMBzffyRvuRJ3AuA/OGZs
NzQHlLihLTFOHLAzEkUztg6g/wmDz85bD+57tjZhI2To/XWeAbI+CMQORWcmJdGV38vCwV8BATJ4
xwlVoysSG9Z0Q+SFAqgHHgLsCrEz+Rgkr+bn93lPI2D5ih2LxCCi+BNcWPkcpr/ng0FMsBFvVp99
Cns5qB4twQtDW9b+oryeZWsRkY0uawo4ziR15rrJ3R0cA0tqq2LV+8/3ehfqJHI9cHmXeXySoXKn
khHp/fNaphvMtUIQKIsXpp4xHHo4a02lD+h2qbmQUwFMhYHmeCt3Z76bP8iN9BgfJcPOXcw3sgGh
hlE8eJHs4dpaJvzo0KymrYlSEyjakPzY1cMhBldLpyqo8p2yshXEto1A7dzJfEPQBklrsNR66Rg4
EH9QWZmRZiZo3uEj/YXAJMVcXAGcCGk59DNyNPZQf2tRqSjGRDB4b+Pym1UGFpAq66uTQCBF4e/s
M/GDsHSKExfvifB/D6AqG9Ze9Peg7XfkWGobIKWouQIHcEuD7P78DVMwHv89NcRlwEtbd7ppzN3n
4+rlBHfKMEizRKkRP8s/soM1i3UcEmbkkglW/iVcBqRZlmxI5L7xeG86d4mlUpB39DM0i+/D53+Y
wFw7wh+u4MSz6S4MR1Yx+snHzTDsyf+S2wbdmT+1Ur7sjKsl1FZ3dJJAwz021VbHfOS0R1g24xUm
1vl6z6shCzmo2pIJ5N96Z46FljmxRXRjUeWlZxMRO/iyCtfourTQd4AFEufVOC89skQJJXlEJF5+
2JXsWMXRfRRf/mSMNtuZ9Qg3fOWdM28ptduz/XF+MsM7AlJdaMPUF+pI0zyRpxVpHryTBam58nJC
zJl2jxt1DBKl3R+X83dXQe4FIXGfMZgSbvtxPsU2aHIEAHPxi8UcFPqz/kSA1dPPyuk7mACs8u+Y
gUxIjQ+SZBGoFZDTdVbWACm0zxs/MI8Nah/zs5QT9MQjkATEN9/lmo4hk1n2yr5NEUBVXWsoRdiu
2Jgk1yUEqEIVpki11dbFdFHaZU4PO5oawI2aZeQ9z6B7LKdJq6QRBK27sjMb5/Hi1zXQPuLVmw1x
hYbgKYCeJwweDixRQ48tQTb7OdZnKqXkfWCZzZEGhq8am8Qg/3igGn5H7Io7Ngli0BiJSTrvVCew
qR1mzpw6yhVSe/2v1IfyARwyaFNBbk4VsHAsn9W8C2PspEdzC7Zs0nMmIe44db98WzgY0RAlZ+2j
CYsDLQ/Yxw7hOpArUdoZ41VQf6lrls7OMJFSiG6VNyARv0GSlrcJJuB/gdssq9T+1I7fNwLkVc5X
SuDBfoyer4nFt7j5CkOZXYEbXBjLMYiVTokSaGgs1nYd+t/6n/htCnxLXu99ZSAtYu56bC67uv80
GKU+aXO0HCrJjQBGvronbPYrcaZrbC/5LqSbxsHELl1jbPbDLX31CC0fz+12Oqzpdubd0ORChkaJ
I6Ld1byBnOYAZja/4U2KuDwMz6IN1q/AP9vb/6yEF8BJ3osV8Jzjj4e9N8ov2f5itAuQbDujm/yH
rk3zxNMT+N0x4UauQFsSW2RAs5WTQBPi+j2B8XQAEMNHDZuo1MqqZg6vOa0mN7vz1N16O1bv/9rB
qc+audNtLAXcKfVW9Ws7KAU8qeS2wWZS8VquOaTDEZSHHkqFM+pSaBRFSGHIQ4D7Rk/dYdkIacTy
xyFMZ0TKnbhI2LSOsBQ1a2WoB0X93PBCnOlNTg34RJL1XWAqIm3tjsh46/04+TGuuHJhdwRdvKKE
clC/yymlYP7vzxviVyWfzBkW8OoVO7FpffVP7NcHpxM7iufffXBaVTelyka/uAncfUWEV4BkYz8j
KOOsFReesnoEpFHvKTR4Xn3+PIXlUP6nsMp6o5FZp3s1nH+4iDetXgu0C7i5nsvtNXQOf0NZfHDA
gTSJ4AnlNUi4iPf567LC7nOrxuQBZXpA0CQj3SwvHsONAmmVPSB2fhecM3qcB6uhaLOP6oLQLRxp
m5YkUVwCvu/JXEFwqewPu8CEY/A6rA2SwT+KHWtyyXEhJk8QPToihFIaH36HDXLJRCvWwtMU2AnT
ZKt5jywelpc4oN2NOcNmsCvHvbLvL3Fq7KerIXYCQO74DpXl5YPSyByFFz1wdPlIs+6Pnh5LOeT1
sKhlPfO2QxfjcW5Ty5KjjZYdDDF72ab9Jq5deHS+vXm8WP4/Uj2Nmk0cQCTDgl/skrhfKYnS8TNg
O5XVAvSunLzoFgCf+zCaZbCeShuvrsznI9QN/GEBaalBwgbBFXoHUvRCCenmz0yYrjRw9qNVZZSE
JjT8tdOFo55JazY09zklU7qj2XX4J8q8EZPF8ZuB3PJjpTojjeok3xKlu8aCcSt+WGuIgWBVbQjX
V77ukk3V0ex2XK0Mj3lM6WfwqiN4GXdQyc/7rJ9/hSHEEJLt6vUAkV0/2KHDvUf8XgiPNuPGXOko
LUdFLepgWuqjQNH/TytKr+nsTSOUcv/T+/1LF/xDUhScimSXxK7tvQQfVKJfwNKgZioNnw5uFrQj
Gm264Ymy+v/EEIC6a4ByZ+Dp1M9wxs+Srw1JWL+UOTjDWie4q2bq1NO5Ny5Q+vytLtUXtburj+i9
N9OahwA7pT9L1spJA4EsRliAWGLMBIcUzAbZhM/cfpE9O9kgw+cGBRvMrZhCSQMa3fz6Q0wZRf/t
Q0rsfZZkU6m8BtHFAUsNqn/4mFpeSimlUvXoegOIeREXAZDkSVRVNxnmtk6zq0vjbfJanRxBIKp2
9C2Sgoz2PaT69Nbzr51fcpVwMR9JYNuzg+j0VJApWREoq/PyXXnBr0ia5yAcRR9MwUnYv+VIrXYu
6PYojhWAx5icBnhXNB6LS+Bp0RyChYnmTy2Y4nDck8LMaEmsydoAKKzf0jI0P8eZdt9j2dRPipjK
R2WbUQwJyOTvR5H2SurFdaOmqMGVpjgNj6dOqaCrSJwMnkbXgax0SEmISbRMFqa5yYgTiGT/n39e
OY57BVOHQglDSXhis2o9fYIPCrIRNzwpaTgpO7TFVclPGTJKwxU8jt4YbfCK/Qj2vsIjFBLY+UXL
JFNHjHjMG5V8JHVKePIwDTCJ53jAxeBRRpDKbWEKKZEjige/t6kxm5E3QZjZuujo3bovPxYR5Q5a
t8rYYAK0CE4vaD8T7LJrpHDT2O4oV5fymOt2avIAsFK662IjGBNWDnupPT10mYVbdiyIOEsww3TR
JFNinh7F5j1WF0quPv0m905mSZfq1M1qIli4+WV2bAq4/T6NwgI8P6gwhJ+rqeljGenkd1GxW+S5
i/8hh4nSO439WFM7iZwSxHngA3E3UMDZ3bQzQA+BlJtv2Wotbc8Qg09KvcImiURKxm6D+vtU8Ded
ui7xE65YP1XwDN+zB4fZG9yyiVVMLIZvrsAf+KWbMcbw1bHKNkP+i/y0Ju4z0Kd9giKkJz8xfGcR
0WKqSvVIxVUlpHKEslUCjt/Mm/DCBfljBSE24Q7uvHqeXHvp8KRxBEqT8FVrxaIsf3l9RusujMLH
mEuo+2WKH5X8u1MgADDb8OJ1CQUtl2J1ZvLKcetDYMuB5/UcPsLi27VzTv4uC/KJzG6k58jBhMz6
MNFRjpPPhkhufw6T2S6m/btRKZezlqhIoPrQEf5manOpsOlXwzMAqk5RDHfvIHr8UqxvNK8HMTnW
RW40j/t559geEhGrf7GIOujDyEmeaZFWAwhF2iC5J2ThfR05mHujF/oVlbXuhwazhGbqsNC4GGjD
tM1PXP4frRvfd0Dzxtt/X5frQKQsOB6JE9/ta4mS07m7quuAPHb2+aZhJbPrF105E0ciOXi06V6T
f6tWbfKOLP4KiZ4tyAffWPgbwosoona4ITnH62ZZk6bmlDG5KNeqotbHS1+Juyb4aFuLYLWkrGVc
2x6casJx4nmbItyJ4cy1ct90qDtuGAc2hsApTsdS/L7nQXduJoi8ZNE+Xz2CooNtcxdg6TntOZ+G
zfZLeYolh/H4zc+puNMugvqJ6tawhrIHe2Mbo+gSIPRGNCCJ82eM6ajJIosjHFdJ0LsPbwOAL1ah
K5iYTsu4InG+sP4n1//GZ9s4iZRm7q1dR+wP7R3RiWNurnN9tBFRjWIltlO8S/ev5aGnvTDj45BL
MDjcutwzqUWr//mgsunG5TixYT8fdKkjHpM20QU1ifHdZpPrev+NyUBxTarYOFfHs2rEPPvJo0U6
o355pDsAYVOYCT8+o7ATjk5/wKUOan5Mk4FyvgJYYvIy6f2kXuQR81mSi3JU92wJPC+GgX3G5YhU
EtktrOT6FO4hyWcwGSKY1HHbSwMRu7W4A6pHv4Zl2uCU9z3dGHz034yUFD3egmIQ7fFJVSKhcEvq
1R8A5dloTKvTS4oor29jPn/gC/6A5bZZu9Q3dVbOMgztK4pmsBllapbaRdFfIlmvLhlrWWc6lD9M
ZAPCwB4FixDgh47lWLsj3zeW835fsu8S0W3vYEQ34yRtYNCzzvhG375rIRebep1X8hgaP8BC1sXz
Sq4gZGrCxZhoyDrvm0eJTQBbmFYuNVFdMObGRpmhAiGPMNntBo0MxNWsgMmIJxpuBkiuQE3X9tiF
B7nN0DSaufD86mS0A9nfyACENNeUMWsJFoK+vcoe0CxLMzqlzhoyp3NsdEzMFsdzHVtYfi2aFwGL
CgJElytsRB93xXDIf9uzo8JjxbRx/RLVlNU02LiyQjP8MrJ0v247+CtMfrn+G5SBq8lTsVUcwR/z
c3RwGdPbR5WedT1ScQmN9nOROFbk/731Vh4TNKzhbA4lFp8XMOE95byQ4x+Pr7QmNSmyOTzpYN2l
cZ4z7qQ9weXpzgQNMY3HNESp0IFez23G/bCFMfFh86m2YIEJ2+rQWQ5HiiPakVg9uYD9RHke1GFD
Pv7/k1q/a9zTNzI+dIFrfyrFK9q4DwYDxT/QkoKAKyMNua1GLx1EYl2S83KgAL2HR8mDiGVPVmx6
uDzI4lW7vUPIVz8ZIDz9DlEehwEp1Yv8F2zUgEuJeWXoswrTwvdYz++lk9scVRuBQd+nctVQLYsQ
e327Dhfs6neFUOx2R1jk7tyy5r2n5RY8K3q+M/6oPstZVPWLlPZ6fVJgRwC1zXG0XV/dF2ik/3j2
osw+o6w0Pr7qHVB9rDFK/ivQNdVXeyngeC5apjHZr/DtrQ/1zm6XZ/Wu2BPYKinCsl1P6zfXjkn6
JJdDIJ9nz7x1bdjsQMY290q2ZifKBn/IMg7LhzgBv8KMfNTB0douHzl7gMxgxmKEU7yX3kIvfEz7
3rqsHtcB2D7OdJH2JW9XzDWpa/8+KXB74rNfzH6+y7L4wcG3EFroczwBy/z8bvruEx73147i7tKv
ERSwWyRHqAR6b/p714PBwpONGGugtYfXd6KJhGun40Ps1U0Qa8vQOARUE0arWByT8qRA41hKin9v
AIlomizWfE0/hxvyzMgaSkn2iMELOpTTxYNV844c+r3g9u+0m0olvlVEcbeWBAodCpBLXTDtFK8J
DQUfOn4r6uITjczSzaX1eX98uWvzHBC8ImHVOMu5/Dg8skPwppeiECW9d4XE1rezm1q8aEmVv0RO
kUa+y9M2uni2C4QPLmGL/Ck/1UAUkkrNDSumVHbAppJ+4CjHMNcVoyple1VeNesnfXXWN7TLuYQE
CVbMriK+su+XY7GcED1Y3Xa8+6tC1ufD63sMBoZi05mtrtFhNucZJq+uLS+EgREB+dr1jevpkJzo
3TI7rhp0DPK1z+7kHisyGN7kCQGa0bIBiozTTuZBCJ2U+jPQFrxH4LBI+LYzqH5olPG4ElVyevc/
W1x6Qvrdk2XFqhjb73lqiOJvdr2hm8SA7U1cbMz2FJaJ9vgATFDDa2cag9u6zTiXYceSrH12Xy9E
rzca8uBRAHE5l/O9XdlhPuvu0gdt+1wtv43DCs6YSt9lxbeC5Qr5MndIYxU7aQ456fUrpXZF8Bwy
wPzGF6dG0DYld/xQJjRmbj6XbSqPwpT4FmeG3ji3ljiopGRw2/f9cbE2mgEzWAXFiH7YxxdlNrLg
UYWNMShc0jfWZTIXJb+sHmpA6VV56K+kEPpJJWPjfKYJ8tZYys0iNMIk7t3tpSVAE4Btipt0wg1K
pBmNkR9MfFRUbLG1PrNWYhE4LuN64GSPqE1+2lZ5c4z+Tc6JX54AVZ/DkQjtJVA3cjP5JHo8qijx
KZ/ePGGJM0yc48jFYbIj/T2JtUafyZyFzXwcCaALpTCNgmZoGj186OXpirvjAn0VAp7kI+AV1DZw
/fwQWCeR/yBeuQ/2DmPgfYZbXPlALcWT4FfhnYibNq1FsDYML7f3HdQmZhb3KHjyoAIhEFmVWkLB
coTJ2T7MDeS+v99ay8+K4Bv4eJrZybNRCvHx1sZba+ebjEodnM+iCd8VTllhvcpCI+zLMOkcA2fd
5CXJlkQ2nCoMzfzZrbKsFYrFcQtLZgkYXySGlrXF3pJrgGV+FjAwoaRXaA4NRVSld/PqffPosbJw
6qIOc0yRI9C9LxaYmxmQlXJp8SHBxfRW+UUsGr4ggMMG/xjN3SSivCdnE5jpAKVXQzwdWqIk2hMQ
18EAxBXUwzRqTRKB5V81TTKv/MrJyNVkp7EE6cErAr1zqC4FFVKm9DzbXPoW5ms5sEZAArNokac+
7sLav0HY6YFIXP51oXPPfEhJG4+QWJEaMeURASfvawfZoQJ0Yxc6ZVUHtigFMuG6FiD3NAjWjbFz
ixVikTWUu7oIooFYOhR8TXAbO8CQ18WxqCULAylKA5VY3dc33n2kxJrdsAfWLK4enJc7NmBmNLCF
O5P3R23FG2Rwy4Ouu4zZS2wIJ3kdk7IU5LS58AvdewmIxJLbJI4o+5HRb+g/jI6Byzm4WNEj18He
M+96OTzq61wSf3GrYfwZyOOa500IrG4dEGBE7PaK38fTf++xA+82KQN+LqnhYuqZRMqGvd5MOFZ9
xxXcv3Snu+D/QDFlGWd64r/MhwR/c6YInoDyuhy41juzepF0g6+8UiiAmJcjCeK97QvQnhG/3w7K
hlmWhYWjvu9ONpdURSi4j1yd+a7svUEoBHffPjtSHODPP1SzsYtIMuOCOuQZZz0SemcExEbQ5/MX
LjQEkAetiTNiInH/89WJzNffP91XSOsBxhgEI0+5nDqTdwt6CkXr5vkimN3rs+RBUzMajBB+l7+p
0Nk8cJa/IL8D/vD9QhNgPYmE+IyAKT4LyyavMjZ3w8m4iQmbMG976J8JH9MGr4yl2sScpUdOBlkr
GUA3BmAoTazNzpAG7F7U+T+OOb9e5BG621WNc2PgnVoDOnZLpq1vYxkjZrRCABfiZLi1/GC5Car/
OZpdpPGJaicXk3iPjZo7/wbYf/bgRqhGBSIueimJxCDHVyiHWWO3QUc/5fp+toaFqMwC34Q7XgLn
2Q3g4dBk8U9pt537j41a6Xw0APyTWL+/YYS7nJLSx0IopDu5vtN4JxJeRGdg5e8uqusYwgr34512
k/dQlGHwSQJ7eczrD+eqbfz4vWc5I+fz5agUUqFXtRsIn2ZdiMv/N/MdrVVTglPSY+i7cZBGkMfa
+bBxorvTLDWqGx8jj8CUy/qQ5Y7woFOl9KoK7u7A399tEDmtR2szbmIjB6XPafKDZSEzUz0bsL61
8krNbQ0ZwDVAym1ZgX4zgpsMQL9wSysqPLNy3RqRJJDgsGInud9j81XSTYc99eRTy0NsgKWsgSVv
8jBUf5UkXw299EAslKBeLAwyRRZmaa59cOSfMb8gTnXPsCbH/lSGDJKVVtzrbNERyBXEX4QlZDAH
LjVbS31EjpjfLzKWTf6E86ntZ14cJ9zYr6c1QJn3iaJqrzFxnjtchXUgM26PirUoQs3zuP3+4RnD
93Ym/Q0vwop5eJ7d/9DhhyseTg+xv2s0rDPeOAK/BUIe7B8n9Gp24FKkzWauRC9TEe4JWZ88f30v
2irsGT9gqkt0DPw7eRUG9RbCM/RdYOxal7JMFjCacAAheCPkAQ4+pGRmnR84pYqynShBxcrenSOG
X60OMy/PMLTsLb22Anps6+rz5xmZ8oqQrWtgyl2buGFQV9QRifXj3GFWheOJYydRH8CSqeu7J+Hm
zyMRttfRM7o7YtmJivZXgM5CF8xHk91BHVybZaJ9YU+92F2wpZ1t7BZw9sbCM/izUsLQqKKgmZ+q
1gt3VbwxVEyWLxViU6b1gmLCwubIar4u1T4v2o3F2yKmuglE8s9P4b3/0wbCoasy5pqDLEug6kXJ
aBfQWj09syk2ZJFZQdzm+iwcarrHJCxG6g329tn4YrvRvQZi1YzIJuY2J3SAvBhDun2BN07QlrzO
cL42NkXc4oWK3YKNXrTUVdQAEl8USy5KrgxD7WJz6nezcoRcH/5tAHC4TyMhXm+b9PstaF6LOM4E
lurlSwVTQttViVkPWgJMf3zXsXJuqG7N7zWx3dg/otcV9/mYtNDmoX49NZUiAgD2mWWTosbUNbE+
ruHVRfsXNFhUL2oROpF0/23Du2XfHahQANnmIKZ7ycZlV53OsVVUO77jEVlmqclGI9fZps8oYMOq
PODI4+sn2IFYSGUq8BqG7f8vBMpU+tfFsl5x8OnEd5CI2+hXSU7tz/4gmuzjN8SBM5TLPbqdusgf
FJyzYlQlFiHn0o9ArmskV1CJ5L2bfxnoBmAft/Ms5QUjBaCKnIPmXJZwlYK9hoZ5FysOMvTkXCUD
WQdePXx99BGmbs7F3ex6a5yCeWVVesL4xELdsepxAT/OEoy9dS9p+Ia4FRlN/eRTvgKKghvKvIHp
kZTH+kPTzyzF3qr17yZ6a27eroQ/pxD8gpZm8c/Nvc25AHPnJE6iopuQSLbizpz1GWbjJuH4Wnn+
emzH1p31FPw9nqW+HewLmKJPgXh/+qvQlnWkAdMz4yIxY7u3dB1juP9D2dDbu2XSTqnAVvhrgcUc
x1kE9c7AACk0EgSpWvxMxBYBSKeIZWyCZN76fl7wKZjtiFGscufB8L6tWj+JAD3vqd61RA21X1u9
cPCAE3hkeRiCQgQmD7MqqeSMuEqAqIA6X4OUcKquhRbEyOA05h15jn5CZmHlgek/6drk/I4Au+BY
9K4QmTys7w2p+JzNzs0O0TH4Ms2aGJEd9BDfVpoutPtikpnJoWAv8WMWEBj/REgfLgGmIkUx18D8
x+kp/lES7nWggD0FfFMkJybDNaukp8aJ2Y2txzosiUt3cJEh8JnLc49epb4jSGdMWlcbGdJQtt30
dr+53HFPJsiRonypgKoOkTrQ864/yAHvqhmEwRMl2hqGUdVh8/WL5NIGzoPjIjo7GSASStjGlVJk
K2ys0jEvm5xji9Kajo5T9ZSCiZ2wyyecDbsb695k7/sopg6sQvfqX9u7RTlINr1grq6EgpEgGTiE
v88l6MCBFPCGgJlOo3IGoRBqYDPpGgRiev2SI6ebl0VmR47oYCvU0iLQxPc2RLbafnaBItSOGu49
+803bAqYx/fE251M4fsUf26mDHZgeLMD+eaKb3iMNpnTCe52SdUzOuXlkuUpWFhPlKDlVV1uVTBH
P7UucN407CfKBEO9KTv8DgAXnHlWgEFy9DdnjuMZQeIoXcjUfTnWU0evtS2Ix6mFuPX4XfOJZNUd
dOItDt9zRtaeEGhG8r3AgkmFXYjTYukLMwLUPJksO78nU+xJLc2eldr8wZ0KbLaLSf8Bk0WV5OUw
nL4UlBxozfPYa3AcMY5yBpT612auKL9bRtuoNtekC7j7q/HbPgOs+OfI2/IxkKBv5kbkz1ktqU5r
uonCAP1/oFWpQy9WOYFew0+FbC6N2O9eiurpeov2XGWMiDE6+eMyf/TJ/z0zkRint+J+SVWlkJSa
ADmBsiqQFj1X2Es0qQCw49v4rRR7N6V+gK8D6lkKf6UDMHu4ha8e3I7jf1VSqugVakF8jBdlCPlm
tAHCnVa+OdupQcOZ6YeWW2WpjuNok0yM3MTJ2sQ6iD9HzsDWIgVROiy4mbQCxI6B0KSQRLXrWtJA
fN2qg6zfbHy4SYa/yLctBOlRhKB63CfIy/fVAtqhw9DwgWZmUJ5wlFkmd9+3WmnGY2RY0xev89Pw
HD7LeIQZaxKKCrgMmEHyb9afBsjBudq2xGU4z7RWrBrfDG4o/SB30yrgFaLa+MKgqZ71yUOAfz+7
/eQ2NL+SRt5dWcGTP0rqUSCGPD9QnDm5BC4wfYGKTJ8F/+PU42Q3/479VrR2CZr4qxR42ws4+snB
Fi19t9Iwq3kyPMJNer65z+vNu1CFZ5DsiLu6e8z0nX1GgxbKUK6dylNgWQATJI0i2ACw0lL7f9n3
iTWdyB2tL7eIpPNdQnfE+rUUx4+qR5OhzoUwADZhtN/WOVdD40TcArMAVNKhgwcs0O6yPm2Hcxpq
KZYNGyPfuYP/JhtVcGQH8qK9YqzLRg5QsaTK4uKGtOTlMLqDeDhO/2OUWCn2Ww8E86f4nS6LFszk
wYQsEFX2/xhx113U0d3MozXoQWUfbIjMVZuESSVVZFfp/fYFcEE7c6uxk9IV7WS1z0M7OzqMyqHK
crtTdRZ18tGvyFXt1I3h7zi1fwkpiXFivcZogSmIlfUZRBvdwY8m+a3n+vLnT0ecgrpL9CgBi4VB
XNXuuRxffKPMTPi6oowsDV2vfI4MnAvubroVVceVD2BxpB/CSzgAMXt7KWqGmevJG3Or6BTHnx1a
OcEpI9V1BogXPtxN0gevyzF5AyvGGkvFZ3XZZzW2YdwE94G9/rys53WEbBocZDx6VoaHY8EBQw2Y
FSF5iCT9i8YmxmUj5tn+EuRkQasHOX+1Km53xsFen2ZR3kyrCsMJmWZiYKANM9qtixd/2z1hyIuZ
qhQUbFW4cCB5IHeI/hptLSzLHRPPqL81SMg4h19p7TPQzS8nlePhPSdtTY0poUN1LVpGkOKpza4k
pozhUYwTDlq2k7QzTVS9L3a30VaFTzSbr+/BxjjCb4CHYqQJ+V9BDWJBp/p/hDBJ0dMo9oNAWxNp
NrqW0c25yHmKnad7h29VDangQdZnO/A68hAb244pQjyWzmIT31ZzRtYPRUCvtU2vP2xQkrzENt6B
mHmwfAvqinp01I2VRHg49ZMasEA+T+2I+AHuGVZskemRS6OnXuj5LA5sWRKzortwtVPJ4NWSnDe2
cBq1Mb+Mj8+CrWRZydEAMpKNVxOl8FFAL5o7Gt8vGAWsNXd2wFkOXrqd95PpGZoOuTVk/L+ozr8c
dE+CyFTtBTP1n5UsnnR6x1+B4UA7XKB1VR0KQrCKetgFqMsf8YeRZviORiw2PSMghR4lUMz8Myq0
IsgJyG2z/KojHkQuJ3T/lPRkejpuc65Eay2aUbG5t5ockPN31LRS5v453LUimR5KpYux/OSL85cz
MlcgxkO2k/hEII9v/QUYHzGmbXz06Co75Xt+qZSf/7cUlhHKFok1OamrRzgZ5HxB/aApocK6+xnU
EPqo+rGGP8VwN5XrGuqigglpwgA4hbsntoZ8RFgy8jJin/bhXsfDHPyomGWKVTmcWP19TSCHqe1r
NhWHenhzDGTGMFJi3UWixGJiJWfpc9R5npKm/7bu3tyY3/l5NZvQEN9jmP9kpGwwXOveino+/C1e
VoKMmLEh45HXun01QvLmxtpRYP4yOH/N+5YA18SpoYy+agYYXSbEggPzzNx7P0d+OWE8DQfWI2Oj
1FUz7q5UZ3nvYMCU5ieeBeta/QPyNvbhVYCsQ1xoEHXkX2XpIJm3q23qxf/FTUwfez9cEAiqgs3y
/cEowjxZammGfB9vIQYdGpZ3+0JVG6OYUwwNVRTx+A1Pt3dWj+JgN97c/mM3376Wp+56XJSoa6Vn
wlQWR826zO1XLhr8/vp92vAxqRKdwuCwUe64UALlzGuwP0IzX3WponP/Ly5F1hNJ/WG0vHP7sd7M
Hh76Jn2F0cRWTqaLG+Dn6d88rVMjn9jN/nQmtKeuleLQKTivEL1QJaYIu5mpLSeXgjxs+RnbxaAf
jNcUXr44c1zoPWjZ7r++492UzINWPdZV+TdAnVudM+5rh4tG7+Z+7qQbKa6Wmsqlp7dkIq8/xCzz
/Rvi+mCPBq2cdzQsHFXUYmFHKeAXFg30h6JdTetkHF+vJkWhUEp7tzGJKfi6SospgeAOQza1WOQZ
njaugy8vkXCzjpyZKmxXMLE4QBrmqmPijgPK4aetQO3tv4v8aWXbD2Wm0PA7oSqnFtvsmcX3mMlr
ddK7IxPgEdQKfaXkl5SkkaAC+N1pWq2Y0dGVbmIH9DD2dSQwZekskLj8ie8aCtePEZBk1gEwMl5N
6S7UYajM4nf9BzmvRgYz82KDVcJ5syJirIrA94BKOdMAIGirAEhYOCcTB9/F3LtZ0mp04ahnnsMv
jZSfoOzEN/MLGwLBev/5Jh985AtmU9fAoN937a0wo/ezW/sH0W7Ieg7zACcSgziYostMVQ57tEA8
CdjH8h4QgW7GwxS1rVy7cTApyHnQHKnWX2jlVgVD5Ylt2Hikh9K4jYGfprSTDoHdfuHTa2uNSsJP
Y9lwY0ZGhZ0q1X1ULsSlyTMNzn7/Sq1zmodej6RJVXZ5q1VSBnBi2UnCfftWPM0GB+dOj0KD+h3H
Vu4m6CIJKWfVDf1JZxysle8midGlgCp0W5p5gBWqxzXUvqOpsIKn61L6knFqq51TeEFVOOSEWPp3
XBud9mLkAyhTkWhHckx8Hn2hPP4ANq9s7fI2HU2s/aYRSIr0t+wtZPaYoXRueK1oBM/G7gjNG42V
4wgEGLXibleCcDLiuHvWXEaLDw9FLbBeaxzEn8hfyHVRvw04MxA16rRotW8N7ofAwkJfjdv1q7kB
oTEp21jeNusIGGGZh3KYhjXNGVdjNp6AVXR/lagfzO6M30XDKknJuh2T4pyJUqw2e4TH3djsC/QP
sHkYBvIm2ugxjjMSZzJ5+/vdj//Jc77Kunok5lL8+ZRHWe3ochEfcWcp4MgFtYJczhHuhAFkOkUA
qhtdgxhJTPxPFFILNUuwSzz8p5pPYBXnzG8ee+MU57U+MxghcvtmyWRAPPjiPgOlfrlF+K+1rYO0
wIVDKiKMsKV89JyXzBxVl8WeEoyHc36Lf2NKeZDKxTx8ioFKNw4oCxIglwmNJ1/bYJ60Y2iZlAHH
GHAmxRal2k1CMv99nKX4G7HTkEskm1YY5L3NSoMReXeNYS028gI294g42bhxuMyM+IThF4+1uQvg
vAIStllMaOwVceTI+0wRK5xPDL7hPX+GALhU/5tPKTRO1R7MXPXQAQjM0FfWZ63mSYz6+5ly3SCl
Jj8jwKZXVVCdb2YmKZom8zqWTHDhjwNcLgSe0zG3dASKqFTKK2fRF1/c6y/CZjc7aU8gOeslpuG0
gbRdlCBBRDgfp/LKVAMmfDoXrTYBD1NDEC+sUQvBR52tk9RgDcNVmhkYV09mDFdEWmLoWRSGY13k
+4f3r5Oifc6MwC7ioGEe9Se6iSTVAlRDhycKqM1izSGK+VN2VrNjn86wzFQ6BxohuSiPUx7irsBL
/y17wLnqd5rL+8FpzwG8WbXOUbpej52QKqjy8ctGsNmLkqWZ51GkHVXDz684+HPnhBW+5m1peROZ
6JxCzYgHBURQUQFX1OoYZBUjAmPKFv7PlBMVxRX8gABYDE8Zqe7PqN2NcxU4NZIxKQ46VIxjTmf5
+ywKi0jVcNnc9ioMkxxGTHk48EfibtohYlsGEg18mO8UKcgDOrzbZICx9/ZN993IYvAcnc112368
oadIKMQRJd56OQWP6A18eFfyOouizccTgHYwh3jNRFw3kcmsat24O1i/P0q804LtBD5WZrUrSlOK
eKyFbViKLFVK2K/QP0eNGsCpu9KWbQ9Neri5Rb5m3IDQlMFnyKeY4bEiUd8CtoiV9picyUOl48eJ
rgRBdzhVyRxYttslgxMPHYmAWUM34XDbQ18DP2QDij3ely+LGvdS6N7tmpzYxFxKDjQaz9cEO8bA
nndBwWPZx5JhJOo1KROR4AdnIyMDe/Uzcv28vxpSr7jNwBoEB6chM2SqTrWJjn+r0UutbLLGbXae
Ay6rtkRRqppEAOeoV/IiUhOuna7OfBcSUzQatzBMuUXcZlGWgNXZ1Fmqo1M16MHrL/mnZSw7d3U3
4YvweCrsCcVfSR3tTLQegDm+bacvSLjRox00zxnFHXWB7bJX7aEfZ1neEv6LUKYOfvARzOfOmjxM
DzwW4nZz2ZzOQpBOk3AP0GBsYckAouQkfU2VOMGRa6lSmMVKZfal38aTY92cAE4QJAbyxfhwWjaR
9+DoBu3NyCtziWNgLevvMhJ3qUIiku52vsSS/3N3n63UYUw0t5sHzRnJ0+zmr0q7yE0Bnpggohcf
1fILycNRVX7QT1Pwh7HJLisfaefZ5Gw7nCza4pA64/HcGiu+e0OfY6OsJXT+g8UVoz72ZszWeLF/
Pi+X0wSMQHIp0yR33koHmGt3L6BakLpP5J0tgS8PyuOU92kashGR2zXbxwqiCifG0Z4Ypp03c6RP
pRzafwc4Znosz3uAaWqpINE0i0fF+iu9e8O5rAbK57n3OM1rNy1v7AQkHAUhDqAdpNnBhoa0PiJU
fjZXPyV27P8EEvIe3zgU0hYi2osUi90+Bdaq4TFcgLf90k9AW3gMfkzpv1KKvWYqwAkhNo5m0TS5
l7bPm66UYo8ggpYIfhmJUNj7tnh8LijnYKuRVzSBkxKknMTvNph5VC5yMVj7ARVb1NFht2R1f0Hp
RSAKftXPOD0K7q1U+r4c2l7pBJ400sgglonsGUU7Wx8XvnjYJB3RjbVKbKTjryhNcfJ2ZDq6sgeH
LTqE0g6oiES6mIm2+Nvjj6CrdJ3eckKBLQMeKPJPTsfqi89OT5FSRpsA62g5Lz+biyblLtMtoT4O
HJ6C2PKzz25NNTcMFwLJVg/n4m05QMK8+q+FkD9FmaxA4AjJ3fAfUELHbzLagXOBO56w1jII5w3E
HKmB0iBgvi1Qw11UrJPfIF5qKninSFghL6gFl5rkpDBZjCMYJ126fDVhOzXHrk3NESI1sSaj0mz4
rAvWP7hFK4nwO6UVyqugJF7bz3ei+7Y8pKwKFiUVUNA5ikdEuR/aDyJkqW/slUXTNYj308Ux2eJY
g0up6pM0Rd4u0zpAD/oa7XnLy2htiM6dzVkHgkVSIVFDwtZ1jPrOPvsE5x62t0reXryRCJ0lq92x
JZ9dKxzfPxje799oflqaRpEQ0K2IS5r85du2HvkvCAi8UV8vzYbBgJxL5bzwIN5SlrHjuifRytRH
YOgB0GK6xM+dBmKpz2jL8tc7XmjbEDQjJXovrGC2oeURgYNcYZT3CnjBcPinUw8HPP/hfMhHMHDW
RasQiqQRQYUGb/DaxJzzMhzvv644p26w0wjYbRkJqUsxo2+NgiPdsdHAgQcjPFZ1YOL6OONetnYT
Pu+/cslywCTVS2KAny3F5Nd5LE6zMKMNAsoi6QhlAWhTr8Mhpc8XDm9CGlIs8nNFypq3o8DhREfW
EANfVDv2AsDZXv65OMAZgnvNaeo4Cat3DFthKoLk+C05Oqpw4oZyGaJDX05nRFFxu+c7CAMSmP5m
85gFd7eiPmM4iMcGeZR0AtsdvlS3ZqJ1WMKP80A2c37w4ZA3NRxcNWQwB3VNglz0VQVhnjXa4kQ2
fMCr7e3CPJ5TdkCkwV2512DDx4jObQMSWxuFd4MEAiNt0bRM80J3r4C41PL9w2rF4PzbcqCUj4Gl
4XqPAMk09trPg9TIb09fWpM2cOPvSnKFtu+ipRVOYUI6u/MsH+tlR9Mcp3v1XkHj+ead9Rha6iAb
HiiJARZgNi0fM3lgmM0S1xvpTt0naRjpeolEbbdHE5UTKdMI0Ol4r6x4yeU43UMdoU9XrxyOzNro
uiKEVTRxOVsBLRNH0NpaLffChw5vT9N15zC+t8PiXFrlRuA1FUin6JvCC2MhbGZ7NacZOtpZQmRP
mqMv8WqVdLyxr3/Z/KEFWWo1JeP/q/xkapH5VGJBsZQMvDbbCGUciNMj/nnovKu69k4e/oy94rAR
St5QOqodsaePt1rkI1TKd6pqiAly/+DPLHDX9qZ3RTwTLXqcEewIgkgc4uBMPhPy+JqdF5I5OtiW
Qei9G28XzArEzF/pN/93VAvrfOpLJd1cpeFHuiI7iDFrTa0zxkyfVTivUuFV+ThzexAm/7WfnMI/
oMnXzp3i664XqHOk/v/AF96zt4X30VTvofmAFWITY30DKaKgbS83zBAUmtKNiCiMwOGK+E28nnO7
1BRFKiJFhPVOxpP+oZL9u5bS+XrZeZhDdj8XBt77LmljGIsZZEMT44rbVva85s7BAWDe3w4wH/SR
ftL/+yS1LeUMAaze0miQO46PejLE8V3xe6qXeXekdvzPui5oORz7T4IDV7AW7VaRsrNi4RQMEIME
RVr2MUbdUYONgAfMl7yOjz9wGy3LK4diXQDsdTpI48SeBHWO+TFR8jZvkWMycr/O1wx1ZfxSiNvL
v+iB7/z1/RNXFdJr7ZMTQdCuAFyPkwRylw/tnmiVnOaXnAnG3NK7tSS+dwbX4WRpccGrt/D/XkK4
F0BAxrQgadd4Gx52yBs8n/GwjP0erG5oo37HtfN8xcWkxStWX7Sx55jv/5rBEaN60RBpc+u4KUEm
aZDR4Ub1rXvq1WaWWh/IY9pKi0XwLMIsl6cYjEjO8cmRimiSEcqj8/Z7QXC0zkeenlBePCoKI5pZ
1rLxyc1UcT4qqv0PSudKraqchN0OCAA+5FdQbrH0VAWDN4ue3r+cfEtntZXbSRbkQ3Ew6UgrzOcZ
ais4JGTo1vboWEgysTTto9zukpcOUfKzokfzIuMRzY/YGU6AN08yl543BwPI08FwRu98sqdwmTYu
QIPQY8IpyITS+N0sKRmatbdAszdId2hECTJwkSW0eLQ6iNVeUFrVkHeknGIeU9vjA0kDEL1piB6H
3ZpzpYhfaSoN3ZJ3Cc9wV2QA4vO0Pk8QdizEQzUW3xzuugy1esmYfW3RuaH1JEjJQYdKXufNoFjI
IitsCG9N1DRuOf+7Fo5FpR/UKCWJwK/aSBZWgsZ8kB1vDTcOPwbDjJ+OrLgmJRa6MTESKi04cX0C
hdGdt3rph/vL09up2o6SS8/RzJ2H8afvxzg0kyKE7IK2uDVMG/+WYk5Hlg5x9Cot/+/BierSQCAZ
dwDe0Pq4rcDuqbxS0yRGnmgu0qjIHEQNG1opnX3oN1hRvtbYK2zwHBq+3TYYmRfBKdZd9EIQXK/Q
Xy8uvxRrHvGuYcJdZSJ60x9PPjLfqj+d9yURUEK6amiJjpWlaNp54zBSPOCIHKvCn5lJeXedEzQp
WR49kAabINBhjmbCz4Xk03A76NEZfjKIZupQ0Smd5lEvPZq0gxoUSKpXELWs2JALl004JiFhkAau
rWseoaD6J/wHw9z6rGVYVmQKDcVHBSk2XX8OVvncIuybrRCkMGpXSPE6JnXTSMcaJac4NB9MpWFq
+Bs9nfScow3X9Aups3S1s9liOthfSDZRW9XFH/y2zCuOwqTS8Ctffo1kwX+G+oWWZ4RdMDTrrzxV
Wsa347IbiDUJRQDVFrZF4eNeE+YNNbB20qu8b2icvSpqJAnHE4/5KJSlKhZe0J0sV/3fKSM6ln+s
IdUFgLPR65eV9vqekbWNPhh0rNe5KIpJ5XeRVeADZXuoOOjZPAaHjmSGiS33zABxIv1ineBsf/LU
wNOgBLIEehlueQKEsQpBrpJumhxSzBQRD03KhP/7DKGYNZFhEDrsvwemO9aKkVyt3G0OIa+I9ndm
qxIvIffKluFLha5DQLIi+h9UZ8q6N3RbUPJSvOEqmkhgVoc/yPbw2WE7gpedYxsfL5ytfsVx/7In
/HUA7e5xs76fKnsFvyfAeo8gbh/Vyahl2CK5XLvTQbW2JAmj6t14HSP30Fedenr6+D4t4KfVHRXc
PFbmyMugHcMKMp/mKLq0AgKC+l7fry6zZ7F60+mE64P6eAh7y91js272q61NUKL4xakAwC3lZgpy
AWqgjLWNpoAYiWu2NvHr4UbOJC3joWJfj70p06pR/Dn1zPglCkZKzQwuoQWFxCPkbkxy8NZw0Evx
B7fMtvZsBeJASVHqq+/PfJgOQR33IL2mUwxqyDWrThkag8v0mPDTew7o1VBLgVQ0DR/IIS1Nf42B
b7S3KcKj4iV4OrLVOQwFsoWHS9Eqn5XjHMfoP0bF4cnORVU3UuNygv1QyRJwyjr3cC+43rLrcF+9
mMQvWAWaUe0zfKH0hnZmtb+nhydvUk68Mfki1tCv7HzJCynvWZdSlgWueqRym0AFCta20wVGxohY
ok5wGrJLwwhY8bHDVHkTwsYo/Fvu8Zdh+yViznhWUPrx7oVgQRSePzR0Bnv9Oxa7LzzcCsH5t6XC
fOrVHMDSLzerD9HEh+nBDf/j0g511M5g6ZNeeaHroLpcNuKp4hm6mute1tMB4Wny1taGJO8qzo+p
W87WSALZC6WQ8Hs4ZgtExl0RXkKqLeviiZPAyO5YZy1//2CbADqqPhLVtRhWe+wkouqVbY7W4rni
oD+nXecacJO1VuNjHZ9coKLQongNzIF4Js+tEMUkp70i0Jc1bSd+4/WA2QjvXUv10/a9+Jvai4Dy
Ga8Od8cAeGa8kTdHyAsHBOlfoOzqZAidErN+NK/iXkcGjcwVFwc98LPrkaG2dYXx2Q4m2H0Hyhuo
i0heAjtW3+XlKuM6otDtiP5ne3c/0OpdND2iaJx1E5qwCGZUiRf4rMWNIoDV3OMo7loY2kWdfdR7
Xd2OV8MObbv0JeOcZ0Iejsss27WixwOMnInbFGEPvi+p0c1n4uKJDIOC70M7PAEAX2GmPbOubURX
C2VWEfhfteGbPzN3TraMRa83Sq5l6TX0a9qM4/O26zSE7eD6le/uzJGv5HC9msDrTGXWCbYMzJ/Y
SKc/zGr5+jZiNIgSBRt9Vl/qc3vWEcAkeWgnrNtEZsfBtriP76+pnBjeLJ2Dog0OCJyN9W8LEQW7
gSAay2eHQDkAFwW+F2/Ge3Edb7Z2ApLe556KoPv4T63y4FC9Yr7bV0odGAM6hkP86lPEVHEou1Ix
bs1jhSjjUZVFQrTP4DkIJRSnPl+0W/41J8i/aickASWeawabKEbl3xYAKWtncfKkDbfZVmt+uKk9
eHnOsVtnfOqJEybq8Qb9Au2nTzivzQhflfo6Ty0neGaiHGNYS28wu+vDSQDzDV4jLjBKnbarxDfw
xTWg/g1ngUoE4zdC8JSVY02w38xpkSogFLqLB+KMGHI+4NVUalQRHf3V4buIec46uLoShI2v5y0o
RsQ3U53DAves79DNFZf5kDHxmvJBM1920VYHxuLk0YWm5HfPwqaLv+JyHhSWh3ehRImxKaj4r7NY
VqNH1wEoA1bchxwdmgnAoCl4CKA7HyiZ37W2wc4X+ayM5urZ6bXcE/ZZ6aq5nreSckFhKT84NHu7
uJob0EHcFPn+q872YLYn9nZI6hif1QByKL1VvSwLIbHCloma4n+gA37M6To8e1KNamBAB4DV7lQd
ho7rMg1xO/Hgi3j9UnZM5OisMmU95I4PcALZR/2ByvcclGHXj3EbjxpWZry4WSczuh+3oHn3W7l0
kYZvhOB0c60Q1ZV3Menl+QUYMi0w/wGVk+oJBhrEy1jl4dK4zPZUY0bXAQIC+pJr0pbMYEVgJlAl
LjNrxxFpwwlYUZTjpulwn8I4bU1nednPldWhhvW+MaVR4Nizh5EK3zq2k2Ns7ObTLvRyUTwper+w
gng3SJvfTEiBNkeZtQ8mDjK5uRSO4JPKcJRnfOUWQPLTG6Yb78ynsVHv54mo0G/e93LVVHVh9PDC
/2EirivIe0nsjTtvb/IJDizwXkM77HEqhVNHYV+9T/r9WQM5sqL+A5MigNeakWZrfg4gKcM1clNm
wxaUBowzGauQxB89w2+tpLRhL/VsKI4PCWe/quHNB5YGlQMflBMpavVj+uVtuD9LFUwNY08RCfIq
gUKv9BHsZi7uChjzkFYVhdE2lZ6j1vjDQMyuFmseAcc6DmM3ac0P4lwi4+LoBQrJgEdppeF7g378
1U0Rj0WjegJ8bSfJjGDez7pUIFJykoNZ6qc//v02IElUrWjQVPE5PgL/RB01RGMeFZgX3lwMTf42
lNUio4N2g1sSMs8q0p1FHjsOOVk0nRK6qnEW9E4zPsfOYvoSr6PeuwT8IE6Jlj6gUbxklZ8trKSW
jkDqEh2gyVBTfmTxDiLeDlY37bfvtNVgZUlPsELghhc3wWuzYT2NXinT8ETj3tjQDTGDtlD+SluT
5UKmNZINDkbQpGUnO5yJcSP1jwe7tXeRl0ts0E+0II1fsnkfMyq8qWXs2E5b8iBArBNaQEZXa4lG
iuQg+f0nlkAjwFNxD7AmXgCpvgMEIgMlOhv8d9fQ0rHzME7m4AFtyED9y3SzuwbQFhfhUZa81R7g
PZT/dUxYiF3J5bRsTDUuLRdBIND4TJH+ZDEgmLwJBcV2IQkmrq3gLoF2saD8ArFLfZTZGsApO8uZ
WiF65U8r/WkhaFRs51BEzwEcW/K/05vJJZ9AvTOutVib088WzQFAGbNn4YsggZO4UTke6YAZG7dr
jUrjucmf7rF2LYg8GIo6/hpp4Rh5qIcgcJSLNWARVn7FqQaIHc2gCPbazlcSsUATk87XyGQm5QFp
xxkliTPbwRQgDLCERbfUNLX370ygcNN0V7tSCO2ZOITtbimgE0nBhDhXA/DR0xB6swctpVo/L8y6
vLzG7DdjCPYcPI2k9FRvTfhDKlW0gOkiptNJZ5xFvq6Aw7Gs2HUPpw6vlEskmvawPNKz4qRwwa7Z
CT07DeaiXYzZs/sRtZnOx9zbpHjY+Hy8z4w3vAUnXTq3vbY02LdZ23R+iNn7NdxLWkAl6a3SidnJ
g0NlunOCaPZiASWEY3KJ324TJiXSss7MV9QMRUYzo7YNltGvNq2rKMtdxh4PcG+GAdDbQFoNIno7
MFGmuxs9O5Jdfm3H2TJsnwCEz8oijB5lZPTPdbkIC9IgkeFyysCPu2wxhGIEEewUEL5A4uTKJC/Z
D49gD1Av3zZFALnjMzT7RZROVAPc1tFuzalVzBGG1yvFf9LR+41tpBaYcQSsWSkSffC6va5VUsY3
YOvlbzkNokU2SfF7FO8eWYgrwWoRRN/rb2biltmH0Fc8uEiyoZo2axT2u4aOowOZEY6rP7Zy0ld4
WlAqWh3Wy2URq5PtSTjTDpk13Yd3IF2nX5mdo1H3vNtHbRsOcwrWlVk8kYot/vLAtoHgxDNp3H1A
3HMgMQgwiVVUbVSEgMTScrglNxfem7235fim0fmD6yM4KzRgssHOp7xMsx6mZCC6fkYsoGZABZcW
d9JEFhKjsJiQ+ntdBBMPcQHpBvgJ+yGZFUWghr6DRdQZIsBDsU3yrZEI4Vm3PaoNsD5BWJwMO30C
ollZeg4A7ZpdGltmZd7L6CkjgxC4HP3z6KGwz4JLR8zkitGHMPEXhJySMBzc9hJ05GBWwNTe1/8E
4RDVcQHCyDOmbUJ5SLtbz6pALU1sSj1qaHAZEFT1oFN8wBppfZJBHv8Thl6JpGKcd/rdg/O0h54U
V1lNtDlmSb6N/S8oZMJI70HSgIGF4obw0ILCSA3MjVxe+UqYm5ms+PBxnZ7f5zpsxnQw/8j+ssvB
HyDxt4IwgF/DOodRqCJh9cHRsa/UKBcVFqIzZ70lruaem9zeBxp+0el00FelRjOcp4Q2WjzjGnd6
RPHzFmvE6ZqmJdFmwazod9sz0GV1gWXLWHQr+Yrw4qc0nvFbX8f+xkGurxdM/Z/iCf+puVBUuf8h
AHtfIvxOdwgkIBTNsSvnKY98sIjjdJyELNyLOD+gGZuTQFvljFU0dIWnSfzYLJHfvLoPOKplHb63
6N2Gzdkx936YPYJ6fJirJoT8AaESnWucoxzY8bD9vxaV68Fq1qTZ8yiNFv2+AS8VC2eDuDarf+dZ
DIIuXIEHDWsvK7SLczkUF5GYtQ3YrTPAgETi+wGksvw2nbtqKgHQHGd5P1+NGBQIUOxoBZYjSq77
zD8UjXI5pMKThH8ubMza/+Wq8K02S6i6L9Y7b4IE1ks+AnFagfRJI5iFUox8xzpc1J4L9jd0Zd9r
Wpn/nzW1ugWgbhcYimpeaIjS+xcjj4XL+gcz5ky/g7xZdVEg0Z+4ftGfrECcBS+SM06s6mRfPYAU
qhsLIdLjohrr1gcCldRaIJLmNwewsHuTKAIFta2xleF/jRSPip2JPHN0bYVvOofeyqeeP/LsOAbF
1SCLCata51hrgORgfUrlDobjJqb3JDp7+OVELCwpGsWphxbVxL1fWeel54DdGXLtESRJKtfkqjR0
KxIMRim1h8xKsQHf0RvbOA7asoheLl4llXKMHSydrktmsWeafqx/CmELENz52/XQv/ntWisr4I63
p+dnoLAl+5H+mLu0ndCCz7hJpCqrbZZIMNRM0C2o4gYa3wtmUn+KKOe4DvI1N9oBdi853feLIP6W
20O20dRH/QGB906wqxBwkDLzCpeT7kDn6/NR8PQ7kPugNY/nttF7jRix0dKvp/OJql094hULQ3DL
OZYhoeErvQ1Xe8EEEr6BvCRkkWPrqY82J3+pHbHLT797bZ2nUzeJZ1mYidLU/4zUSw5vpP5fMnqv
Hzxvo6hF414AypGtBLeu8ZFUBHckOkulTf20/tIwSzqk0qxC3eCJRcDmBhe9XFLJUcYIE9426K7F
pWiqSk6nARKgEhWmboB8bsiccwrqmGFyRqoTLatpJuJSJm0vxB8x+n0x9GRyRbH27tf4tFkrMPpQ
buNcm3oUJHWNZHqosSB9AEV4rynzRruqH1PmtZvuCu57PcaxUku6ZdbZwkQch5+pr9RakMd5S/2H
3csXFD1Msd/PYNQ7MeR0U0bRBlv8LjSBBQcpZbzoxGk0hQePF9vDyZL0lGmZtF6R9HzgiNgg+Qw7
97JCJ/xeYEXegu3TM1yx4VIsmDIDErM1vhMciGZewcY4Mco0fNf1XRbkd2Z46/V2/VqzpI0RpAVj
kptsG/Zgm8pZsLewNHGba2SwvMBsZfjlu1ux6CSbXcqJ3tcSGCAWnP0NdS7j9GKLXrSfcll2agB2
mFJh9iO+qA44HIhKiUtJkH5eGtkkSyK+rdcuGGfI38aW1jQPymRv3MP9v7LtHXelPrcOrDPehTBS
gKH/RKVu7WaYi/r7tMYNzPqXTOXrJT2vcsd87XDvqDp9F7nEmLpod+SxuOGetiRU70vjoI9bSgmG
S8KlJnx68WZVEopWv0XxvYVrjB6Xmbw0z/UqM3RqfHbgXnGiF/0sm4CUMj+oCRNi/fbqVQ1DvBfl
jj1yfUQKarJP7OJRMMbXwWJNJaS2+TNsuhfW76hdhjJSskCy/Tt3Tt6bCBsHI3nvkH/UWyqrwwhd
OkC0csctduHU+nhz6zYLLwVT67cz5w8FGWN5R0yNn4QmvZR8nnSz7iXJR/1xWuJgNILAXPVOrXQd
RfqBtbZeFoRJigrTZTtvyiSRQz0Im3HYwKKqjbvuiHun/sHFmFHZvy5qdF1G0qUBNH5pknxzP5hM
apFeszl7UZbYwtwQXJjG8MiBmjyinMw3icqKZp1I1o9IFFyZyuhTDMFSTHYQ/zA3rjqc6Ii9gWSf
yVWzq5Gu3+8XDTHZP25vV/pgFkggvEi2qtb2cLFNAM+UgrpjMMuVga9QZU5T1Mmu74ZGdkKzbZoC
+B4UTJDPbYHKoJfqTphVoWbL4wdibAL6/5C1dSiMqHMUQyzI0QL7sf36BD4dZFSnWXGneDYkiVCc
mOk3iM60YHgHnEtXSbmFUWjIyNAfbp+Av2rR8nNgt2qa3XhSxxqFHpApzOMitwVqb+VlmJcWYJ4i
zk97Hv19yw0ZDbOPB52X4Ftk1oRKHw65npQ7uPC/vuqNhMpKReVPuHZ3j6w5AMCr9upQXxa/4WA1
W/uwRd64qdc9VGBCpej8SY1mzkrHn33CagvBIPFn545gG9YHS9D12MCa9BlJH9SabdjfqSfKBauz
fcpNAEDlT3txBKZzV4gHFaWsRWsecJyST9rbCOuJGZ9nh0U0hkMvzPiKz4m4jMWVDjf8zAcYtF/t
lNvGtBsz9RvLrzA6s6PyHf8ljFrTM47m7atP0hNMDgKb0fQ80dNGyyZVETWiMPMpVczn9JrKLV5x
Fb3PicIIv3DrsarJmZSHhlS5wxqz+1tunmJzsyRyxncAtzAsdjVzTK3xkh2RZkdCOuqUzEDUlt1j
GMWWGYedqE9DZZVay0nS418DLl/bl05uDN6ffo+EbBwY9xtLVgmI9DVhagZwTCpNje8fTM+F3ure
RDISV/tckqJ/HGSWk4K14/hStJ4FedI/ncq8kH24SSW0hpd0dacqIi5k/gwb8oWgl9NVZj0nexfX
j9piWwHmGN/GZVEZ3H021VzfhL8xlKp9PidvOqAWaX94Iq2QHDfs8ugyejFzbY44waY9fUmGjTW1
IUSYR3vq3w8oTzY5akad/JrOQyU6/F0y7VAUvxR3py43IpPdHezAQCBxsMQWI5EHYJEtvwFw24Kh
hEXu0cudzezgQ7/JAWQSnh1xQmKhNxTrDenwM0Naq3zV/QMdizVeQpNC0WbtGGiJL+0c1wQY/0j2
mDGAkZF3ViPCIDYj+5pwF200DaXMJjf9om+9vbFHUvxhu9oapAIQ04vl4xoE9sRBoH8DQFOB0LF9
26IBHJuadBnkpwaz4H1s0UxfXhL6qalvh77Y2r0DSWs8UlW123PPmRDJRA2JYxqmkO8YMHNAi8vs
dgww6kgED6F4574TADz6yW12trah/I7QUJUIEzbMioRJHBPdUIUSgiAxL0oNDBbGY7Ud+rNW1Ji4
6ptywBqE4yPhIvHrA0/Aj1AuRgdXbD7l6QB99TICJpbpic9K1Tnz1Z58rB/SFLCyVxVyF01RXdDe
qtvraMCkgmzTqZk4mglHijpj/KJu5bBQu6tUdT+LxVqkhfsP0AyfLjlk/VDYvjoPMcCmEa7ikZdy
Y2IUVfNro8GieMilpcGebrWtuVldKVE2SnPzftAZZwuUAY1BxobVtfmWFoPJ5y2R+7DSOcbIMvIE
WdAx6Jb9fbeYp7cN5Vj68/mGM0g6YEMGagv2Iwg7+FN6NAoBsRaPMMpuRZPfd1jsh3x+sZk5W9tF
4i6soTiSyEdfbVpWPtJeyaBbxhCtyrBvkgoAMJhy5kTpeW/RIoffa86/nuJFrLOZWhzE5QosJc5C
YXDBeTvgUgGPUth601xjdOLQjXsPIQKRCbuV86Zr8Qiqv1yPYU0hCcrBuTYYYWIPvD+WcHtS904K
MoaMfGr42NBc1+7wQC3DJPBxORXIg4cCW+Hjz7EVWAXkGBXquNvXByB+o7AXezfIkp+Ey+ejlLHQ
rS4LwE2+ZMt4vF8a44+tcWnWTiBgIlmwSuJGWPYfWNcj8p62BXlS8F5/GMmuefznbh4fdCWF5Tlg
EKsiKji/7vdTVd+U0L8McDSHfyIrZlPPonE+KF8NreF7ZjnBhHwny0B1PaHA6d8xNS0Ieqn6fTIK
LY5K493RI3H2jiPc+XqquPk8GuqbDx5o46C6l1dlIAlEBO/DDAaEeTqWIY80jAEWT/fqDz+XjaNt
Q7oreE0Vr3hNld/RlA1B/LC/K5BHoDlN8k/xWXqMbAoy0k4A0Q21ASda9YcDt4u5nKuNSvNejL3d
BCGEhjhEPp9JGuFc721uS0PIWYZ9xgzNWp6OWOdHgwTgpIIyvFXyPlJKwrWK+124djFYQhD4KU2c
gEaWTTZtQTdHckDF1oNdrXx/XzHYIhrPY2diw5+kPPV7biFBc0qVo1HYC/IGJ9QTSNr/7l5YcFaR
35ntW2h7Vut8qMQD26QWHGYpuNXyOX0axdgktxO3PJ0+x1wCWAhWCqhfrvJX75MDFFd2/D7gzCpg
Yu27OQCHxYNP4bjEga09jipVca+AIJq1VYeVMXtIvNIfyOSEda1CUoWPlFuAuIjjL3ZipoDkMs56
pbiIImSGOF+88Z+GSh0F7yBdZi2SnpxRKNULUvc7InY0Mv/1BMdRx1IO4+i/f8wkvrSq5BaWPCca
wTFi3oG7fgdUlHiTjgHzkmP9CZNnF2Inp1tvGPK+kNrmOC8eENyY/vW83jGM3N08FiY9Le7KKzhq
CTRsq0gcPLrEluLmKoCCyN3jpkAGoAGvs9nv3FzsO/Zf1V2rpCEDlAbykgre+rasLYMU/mu++wNZ
DxxHmKw6gjvIRTPvz9a+G9fZEi8Zqyo+bas3Z/RmrRBXySAZHJQ8A36a6bRhP5FPUjuB5xLVG6dY
Zvi/1a+mLYPSsGACNPiwzhfd7qoeXB/Fb6DRBFCmcmviWoGRHNZ9zGcynaSQ7GKgkdawoLeLLxZd
tI5Zkf3iZInwRKme5Cf+STaVPrgpg9GUSvy20HHL27WYbCJ7UrJMfl1GAkBYyxkPA4ncQZLTJmRY
UTCOXx08xfPuFBLjwU2Wch/QFtHyMQK/2qCnwcgFtU6LqKBu/cYiub9ybPxD9VnnkPdV5mWbq3/J
9Un28KtVmnPchWXuElvKadbZDX4RtUFLnH5d2Up2lO1IOFdFFsdZIK0rGWz09t9x9yiApeYX7iyg
VlRK8iAl34j1c/lrNLH3WRtJkMl4ELgQ165sN6b3p5k9ECj0d6uVk1uymibmg71X86qpYGl5rjcS
gf8vLbfjmphWgmn+m/jSL6gRHy33mqs/uoKMLGOkp3JTg+sRiew6SZ6iytM5CR6+05+p2GC6XEKt
46rp/yLOWNaRtAYh7MrwEf9ljKNAAthRfOvLSsjli6SfZQA19S3qIV860Owzsq0eaB+tgwSxloo/
+MHvwn1GSt9ctkdDFzxIZmGkRMcDs0o4hCVXciZZ/JwKlHzYCs21W2ZDT2PGqvLRBbFaSFRraW5A
pgZ1sP4kQZr3ImCGJ7ydos0uENVFxAEsbHl/2xITWJ4saSs0SsloOiaLqi8J7/NqTyK8tGyPyWbr
c6FusFn5jMcPQ+7oljlh8PJefHHCi3rRGdlgo418vHrDod+f8cZUYz9XaNwyT+rskxoIVHgRrWW3
LaY7wG76OWGxQvz38pFBPZ9nnAnm/jhuMHjzCFY/mQEYFI+j3QKt870q0NLDEVtzl+DSFeptoscU
RPT0xVn/kHqqbiMeVXJ1cV/KSMyCAxZhfPnPvjjMmJgp6fa1WPzDvY3oHit1QI1zPE0gAC9sBv9X
IKB9fI2+8bm2RKSo58G2DflYQEJQjVO0N3sS90hG8KZ3QwvLUUgznmJGo9D9SF4FLWkaznexS3hE
TLH6weqYYQZNCRnPHt80fJGazT6ZCDPYS9s30TmFJVUmxCPNH3iuPiyn/iVqr+in19EgvNF3pm2u
gPUTLRk4ERqKs6ZlCEGkoGMn6dK1pRPA/lK++iUWHiFoshEyHoybpvWOP302o2Kn3OHkhXtkP44W
zrayyQkMGXYSlLmVVVTxjqJdAzQYr/Fl+HDK+RpSwQD7KmRA6kql3P5+1Iwy0au530Uo2qAY1U5g
2jLe9nf1nsD1DVmUKDFer9S7O5EIRDT9vf0ep6QBHXJ+uRzFDvj7iz/CJ3fh9/4IJ4CL+9twqg/X
QihuAeFpG86iSUl+JvCqLVjHZYTKnH5ah23bUqiMkXemIuxa/PkklRmM161RPOBigY9XLSLlBGFj
PcF+dFtpqVR1DksKJJ4kxP7+qRsTLFj5jJRmsXrC5KP+5ZjmilaRv64vEPDIadyOEWXVxi4hOixP
63hL1L5d1YX5vrVriiavJ1Pp2B18YVoeqlpD6D+gwYDFanwsi7D5I69u+KnXyxxYF783jK58mChr
5Tu06domPgZ+Pk9Ux5gzCOXzYC0JAzX1DPZAq++FU/a7xhBKy27j4AuX3UzRJLz+sXyOuIJY0luW
PMB+sezIS/rvGuq1zSvtfc/K+edDGRZfp/hN5uZj9cyuPnXAQ9w2qegSE5QcStWxr6P/OUjxCiPG
eTWdslTVgeU62WtzI3qDxLXKz3bd/TtwVChIJG/8eKhfbpXM0W2CmjzjnnOF+gXIfFE/R8/O+dgX
FIZOGYsdr1hFhXzcA4JIchxoYvuUa7QjkVZxlsqZanfD9nJG+UCyZfZUcLtpQfACDnGzJyd7H3oT
Vj6d+eeK533xJPIzFv3EgCiQCX/bEaqu5/C5XsoGJZnZafpwTzjzKolzBPPGmWOfbA2tFWBDgsqq
v3FQUArGLr8DRuKttmBbmhWD2MGlfCoGyYlKg53CwcfRAYq5RjIsGbpT3y1iBUwoCCC8RPtWRWPJ
tdy+mnWgJlgwUSGmZojX+EJBtZFTXoseMk/xWAR7vX0P8zBDwshlsczcFcOAK7GmKlhRCD/maK1F
w44xUeR8EQsKATZXIbjVT3dJadRRK52DkMDbFW/JwmJVsyVPIpuD3xGuDEGz8mbuGCDfD/Oa+cm6
H8jV6+1Z3vsgnhBxUTMw9piDTPckxYzCRU1ei308jCQy89flAyyTUYNQXkBxxpMaFATZCZdWXr7h
sHzJKYbRhmFJ2CLt6upri0IiLOwu8WkVTOxbHNyAlZVrTfkK/UgPCaT2JSESv8KMJlRG+McSUPb3
U9vsef1FvpvblIVcbv4IJjCZSS0XWZIwZj0Rmznzl3vnuTkPphBJNXfC2sG81T2S219LgGd3+O0Z
XptbxXuhwOCfXzZVkb+oZ2QKHgonrICGC5EHTWlGIBe+XoMla1BMNCWPlF1RJ51r4DawcvDSNw00
f3zuaycXPxKukAvFfusEk05IDVQURP+kp4zClhFx62pztjpYPMZ1//yihobTNyjEnujp/uGl8RUs
axPU8rhBjd2HEqGDx3cMF0fKmoARKxqqwRxo2Wc4c1ZlLZ8pW1urKnJWDS9vlSWrCy8ZVa9Un9QQ
bRLhHhzNuMWTTNcJQxliHW3IQ9kRO1rn7NTRA11SO20LewHRlJRgJ2DLG7ca5vcwGJmtcEXEPikR
jkNxSnqq8REFFrnh2ZAdmYF/ZAbL9X09tUrELUcaYvpFLIDJ/Lkuq8BR2wAaj3zCsAmETIcycch+
XZUJmJsOBBa9Syk+ir8g1XeDOwOiSaYzXCIzc7uANyjQzY1qDU1TrlyPH9XCJoK+5TMuAn7RiaVW
lGnydqfRBXU7iOnKs/FFy0j6AmJdNQ/0aM+QJlZgcxCM48d2TE3WRwJljF+Uc4LmaBtIK4oY9/u/
RD4Ay1C68zYOY5H2/7BtXEdKvzoxg+q7h6uvYUS2gpfnk+Jvtmb5fpnW2YKP3iGbqAR8ANPF+o2Z
10Fo7Q41xPV/KfkR2gTU+VMINrPyb0Lst8LpjI+qgSPv9viT3JS7EAMEWIBVfoHj9PJiDQAWu5ua
70oYJe/YqfMF2Rv2NfTJxghDGFYV3AQYX26up1g17qK9yj5D4jRIB3gIisvDv9LjzFZU7sKsjbrF
MSyzV44ZMI7aBMFVqUALSsTKSwla1CBHYgXgArA7soKRvZ8Es5Ah5f0FxulTXrXDzybud8EbA9Ug
6BdVUkRqaO0iyyHXmmlfR4SVfx6b/WutG535pwBHuY+oC8S1+tSLqDeQtZ0GS/WwFz0UjeUMOs3p
KpaIJWOOaVByTz98jpLqLpZjX0VrAb9Cbz7C34XdbRgtIEtabah9eyBlemHAL8a/25aSPLeCkLWU
9EwqFkS9YTcJlMzNnjr5WZBzMe8GrWbRFNKnnTS2VWkURtFrY/btsFrVrXIY2ebdD0En7zrRS0bx
hTiqRESp9cHMEQOZPD4/9MTVFAfPHGmsCrKZyTu5Co9X1zbIYAcO78kMe+tcgSUgNnyxugicEtuK
gsqTeCrN0rUb3EiKA4Ba2UGHiIz+0pdpBmolFRl8LQhUJAcLZxPMSAAV66E2OLOxzP1YJ2A/GvpH
NjJ13GujT9Y9VwbBgZqGd0cQiorn/MsvMe+dEoiqVd/OpF//uiRQephJfwSCgcjqU9SC8C1bXqDx
9RcVma/cvChNKT9PnXl5YNj9BVFiHRcliBAfQGXNqI08bQDo/B1/2xf6lUAT18bBT9y/ZqymYBgO
3w2220th+AbwyaG9dgjDUygKTtRcaMlSXDLzfBkrrV3OslYtYIaQoDgkVAdiWgbWDT7WEuB/iGhv
W2CXIizDQG+t1ZvqDvbeV0AZvLCQKMpiBJmVKoyasP9LrplzgvtvSFn1zq3puuXLsuHH3bW3p9zD
ajnlpFRobtqdg0oJqnw3EDg/uix4rINelUTCQAvrijnxc2eAcjL1ZkKL/p7va0lVqd9WL8TA9zq9
jhaFFrJ2I+vCjxRisRWEba5H2J7wxTIG8L6tehI+KYGmK71FLZrbNWNbYWXy4TWLl0So39qWOf8N
oNnRonw35YQpgLMwP4ezUauvMbwphGYzKqgDTL/FwsSmVeivAs9+F2okgVKwtv3sRTnc4A8tjDw4
RAOVTg1RPKqYvoUDclipiga5yVxDRvZ4w7g1GaRIkG3KQjEJvRmexJ1/+jwlipTyzF96BQCFcH1C
5r8WVV4U92ypArLTORUUs8VftCLHILiPyLPtu4HBaQzoXV6vGO1WD61A9bJp1VvOn6+MTWnBd/+v
/mVmYu8EUvuvK4UZ5cokEb9MhWgLt7de8f7NIqXnpSyiaQpfNtXG9nv4Ri2gsSESPpmw3Nonqsi2
v2hRAbxe5v5Z+VKwh2LaF3z/EYaMY4gnMI0DSpvyuU4Cd5hHomUL5FI2hrIN1/upxSIL0hT+ArFS
E0/bEvU3FVLk1yxx388j9bDQ6f7CaTstGOeUg1jsHSZle3BTQeL768745vvZ+XV3H0XlZL2vLV41
4LMF/G3D2Gh2Ss+wIZXvMC7DMaEVwaoOkxUzipvFxYGUM2zbXj4sQ0N7nH4RWtZnV7NFJ0dfaRiN
lvSIa2I9Vq0GhdT3vMgZRDnPrDKCIzRO6BMEnOPeY2jeh8rZnF+kHXOr6d6pHleiHFGi6JkiiHHa
TrEUpIC6Mow1Y/vUw1O7Anp7utEXFeZQ7DhHrlm8M50X+gqC4svUcBCT+dNX6p95MLmuai5+pVDZ
b2Jexaers3hh1sF/sTcnzJNupSDLN3m1S78OeKQZoHjOF8Nsfwe0rvTqxLXuv7LoyJB4Z9USOu8f
Pzdg2WJEvEtqMSUf7IPkzLp44KX6DCvI1WFGE4HCclaSAp2/3Ub0HbUK3wp2TFgxN5TfeumDKf2h
d795dQMrAq/ht5lUqZGG3pNjA3oJSPY6v2bFE12RPRE873xoW2s+iBp07z34GKKT8OcfJ/21ibqQ
vw926uLExNmPLX3+iCP9cI0cebM5rW4NygntBFAhmknO5vFsHfqc27UKd3u9tlYtWdF5ftVvrhIv
b8rBjZViArpiy0D+YHGdv5VLP4tIa0kxx5sIhS+X3DGDxuoRZaYD+IyZoOMJRv5C+GJWfxDDiKFe
6l2ZAZq2/90schQeJhhImzH4Nw948O1pIowPccp3m5EGevD7QHw/SJwMHwFsn8+wyfgAg87u/Dom
eTOSHsDOf/V18IuoYZR6WlZF+qdudfGKgIr5uBr5LaDhKvmbqGq3gMP4fk1ReddrXdhO1U+vaVou
ck2P3q0ZBDUj64klCzrjjv9e147ozxjK4VWWeqxmGg1Vld1emdMAM2KCC3xMN9Fk2qFnKh18Qn0n
VaetgzqimSrdivM+3UjAFiZAM++gf9w54lRks/Rx2dX57XdORxqeOKm36S80cJdNiybbw1tePrfY
0OJDxF32MGGq85Fd15Y8iP6+2q/ksE59h1UaW46lWO0b+SZViBAclrh7fkwzv3o7grn4NZJy5yEF
K1irQOm/7pMJotqT5SSQHzu9IF4l9PauoCKy06eN2iWKkc40WIquTrToeJsYSfK2yZkb8gpfF/cb
jY9jKOMnh4jTeOtDSh1V++XY+l9JMd8bqd4r6zHz4ucelBKhy+Y4ky/xG5Pkia/iDw2gW0FfoS1Q
DBmnqS9SRBNSg6N6Oe3/3FXbkPtQdRh1w8gqsZTD8uGR/PqNmQZwcDBYO/5KdxMc3qzwZJ7NaTEY
syOY2HGPduHmcqr2lKHYR2IvhdhdO6C+H9+iK4SxYRwwvJrsODI6FoKlsQudL770O+xF+MJi7nG/
ICWWoMEVFHGiUMcy/5vzdNEiDhYUUzV+aLbHAKrjgHILjALQ9rTLhuPj+80jXPddd6DBUdiCVyjK
OZFgfyxDudMKNkb7yxoolftYUyDsYc1p4hABF8pe2vxwTpOav0iuhBAhGHt6Ulv656tmnZs1boRF
9zWq4DlVBvYOHXNq/tifzXGVPPX16GFG0S4XUFDT2RdbNe8kHUPVjDreFgpcB3uE303pMxNWKQMX
zlOgzZPuB4pO8/kshp0p1gRTjb/9l5YntqSAK/T4zZAFBMeIZ+Z+kXl6iww+rRrgqpq8+fI9qo/X
03NOLgIzsOJCvKu0+5IEeWYFZzvf/4cC2aBSuEiU710/VmPJbPu8m7g5g8y9LUYdgChk87hPriTx
ZQ659tTuRTTu9GdzQGpEzcYOoIup7bv0dTZtcQxa71LX3mTeW5FEqdZAFrBl94LQtu3h646yd2TI
YLelvlG7o92zMU1uFJe2V/pmLcJ1o9pcy4LkTyDCJ/+MKJyHzYSBwOBJTjRYdtbtp4JR1JHzG7nQ
eQQ9TcplVxBTJTkmkjSliXqGkKLUU7RfBAJEQpTaJrKeDBBpBVQSzSzsupRHCvC645YgKQjhn1t0
ZZKN/hnJ9dOXmWyh5tQCnFkE1+mEryH1oqZ7JVdkxwLAY2icP3eRe2S9rnj6Kt30k+1wW8gXBKbN
1SEvPyvN/lxli/yXJj4udFKn1lcItz2egsL+MqhVsEvIfJFYtPzEEQoE1zCTlp1oC8CUQA78T/Zz
l06t7qci/N+9FgnGtgw0MRrNnMf23IJYdzcnaPJgYh0vca47GVyJmgNxDfu5WwcisSCdflVA9DSL
C+Gu+vMituaKxbBB3BCA2v1gN+AmCb+Gyvf34X04y6tUZDyIl7NlUkA976OMLu6P3ZSePQJ/2BXc
q2wf2Adk89Bs0nQX29Zafl7OXYmY4inAiORoIYisI3CuukrynVaK94FJatslpUJDn7GmveIKI29E
xGDSo71o06haUAQmGrBrw5AIqniLxMQjh3EJbRmeWrTgFQYP3Ha2FKij99eQN68QRjaiIXeCu/MG
mxMOHoJQvPPLCBPcHFB9Yn8batn/cANdMw7YtRteKBJHyCO7a+6grnQ2ZheMaU6PXGxeBUFOmYNz
7mjSWP8l2cY1NTih2BPYsQ+Iu3uy3a9wC4bnbgD8NLxq0W4du/HAjEwSb2Xzh+hsKF71152lctB+
W+ypn6bNU01JmOhmkUECKbJe03F9gOZVhAYWpiMnLApMjPARfEZ/Q8Zi3Rq5A89poc0AGVfRkMV9
4fONaJfyZpKgLLeKeJssDHXvvEAnCvki1o7QQgaMpkh3s6pecve/ZUbbY5PojQC2n5Rt7nLP9wux
9MaZrKktLdbkSYMZtF6udyEoq4iEj7/+lfGh1BrAS1Y5+0nvv1V+ZZOgrQMOYCXwesYJAAH3Xwut
cOeAEPG/p2jmnFFYT4aUScH2GAWr89uf2ElbpXSO+p7zKM7UF8tuCbJet4Ax0hQFfZ/gPPuppGeF
dY4KqrJD61PrXSqDSPx+ECL/U8NXThPo34p3R6y1NoHqtg3/NNhTn5CCa1/1ABtVQOhARg9cChIh
Jrsj4NAPeWSr2FhRezEOH7LvBGmrKQfaXE8i0a9rxWHaQmaaTt/z4TNQ1oklRpiyj+Juf4o/tSZF
ad6sUah18UJsmbasfd1vhO3BbR40FFdt+nGRSfljXga2XVHoB6e+ph8ZKVlMh4IUuDr0RGmJnty4
qGyg0LB2juF00d9dxPIOhS0BggKdpox9+SC+Dj+vOuBT5l0kcbnk+swpvRPRnUoNKN/d3qvKT8p2
VVU0Ti7jYF/DSxCap2MbuRWZoG5zK2cZK3NIWXrpmvZQaSbwlwH0ZDOkpbclLz7ZoZZOrh1ssjlZ
zauPhz1EJWjix0NYEORt/B43amodz882GDKG6eXDZUfF0R1cUhTIN8r/GhscxAK85FHe1fuJTKMC
xdJHvDd+2dvPhqmir62w5XplBpx4doa4BEAE2q8kWl5pN5eAAavXArEFJo6pabjQIysFY0kIBYbn
yghTNN2irR1086sMDtmkC8QFBcNzz78gXqMGlnRUE2Ix+IpHG7d6+I/WHAE70/SXA9VFG9ovrve8
FV5nmz6MeJXMglxnop82zeTrfjQnpU6TSILslqlNfi6K8cmFPl5X4o5MHsasApFxRKVlej92pE3h
Z9MOyLVwOz5bYxMt6TlkNR5PV0LfsJuXD79PYGF1dOHwlJU5zpTHJus+h1i4/RfP6qQm9L4sPmYK
5P2aTe/uGQ8nznUYSQZbNj1dPqky4cvoQ0tymRQZjwz8A89nYmRCDvbR/35REh0/VcBCuSJZS9w5
B49jGjyP2IvxlBdEpocQBeesfxfM83Rucr3fPU7AMymBPOlwZPii3ZiJ8qxyszoEhG4L+R1dFKij
uuxeLWD8xPPEN/+PLud2HwF4bvZ9QtuQJmlT+3hKxYPwpDJ5tR0DG0/tQ9vyjbaaaOtOfDcSfPI/
BWrQWpgn/N9nu2//n6iySrgwHcONws56exS4zOVEDFfV/nVQMj/2RTCBEz+kPw/J2SnWGtNf019F
sxNY6zY3YO5cDyE5Fiksiv7r6zxdlQrCmLdrmPjTqQsSObh6n3pEMXUgwbuH66972bkDvIjRt012
1XpA8l5AxL6uv135UFt5GD5EM//6fMlUz4wydAohme32rNUGHcmiMGx6Zk/XvZQ/5T4IeZcwBte7
d/SzQB7gljzFMd8Et3KibAf1Vgiew23XJQ51vzwxFuk8OH0MTu0d+vys0tGkI4kjvoE02verxgsg
Q+4fB3dbHeTXZUwEv0l2bIPWt+8Skqym7hvsI7ndVLfRSAMzf6CMNdXx7/rNZ+JRuGUXHUJfecT7
41YJHY7rBTL0QvE0yHzdPbaRcU4ZlR7edqDXYn+hXg194HRGzABjF91TI7hJXvjl6Bj1U2Je1b0P
BILDvuWowoW8STLDf1KFAXMKToNKjJDV+Xdp+urzkiaZPJ46I2gNSUYMB4mc7k/T6BmM4h9y4LU3
d4jD/PCKEH20OaZ4t5mRelbvHTN/pOQIa/k6iuYBHwlGqYGkj8DMs3ASRXkAiQ864loXWei5LcXz
dsUkFPiB/OazNrjm6CVgO51yRwAENGb52f4ezz22cOmAUUSwz5NSAlJnrpkUiUXHx7fTRhDra7vq
b4XRkHWuFZ4x4HqV9dTZaigSut8t3UDqBdoL6ILQM1koqDbV+1Aubk37HL9kgBN/I6Sw5zSKTZGh
+KDTPGkGe0ibOJ40ezh2jHFaRcPwgkF8ES/DgW+RDRYvHNdwvZNb0Qyajy+Oor2TvikfsTwNuW1p
0uEeAHnvGdKk6WzQu2U4HvBkFxZLTOgWBUOVxeDXPCLHcDvBcO4ehEfsJuFWaXBfLRgi4MPH78DE
Pg9TFRkCE653/WqW6MIsAI8BVPp/wlC8fWhe3Y4z2AkYzjLDR2owbHgF/+YhGLaSq58RFFFQq7dE
UA3lLk/Du3vfaEJDZlti6wbjRxrVVr6irCTWzCQNM4pt0ceD3eMoIwZsSQM4JpBzMnhDkTcwX/6f
RP3tGqV5QpD0kYHw7MuvIqUb1BoBeRhq44axSkZ24mZPqx8jYHmhEMshqOSUZ+k5YDBiVigfa8/u
VIMnA91GxMYnfQPSKoBCB3bZunh9Ln7xd1czOgQVqTAS0WbEd7PKwkOpLqSrjdIRmW02mkk3JBeb
XeV3pK8JW3F73DRx709Y2G401rPTz7sWj2mBUI68jpjtf2UxoFka/5K+0qDkII2zvbPSzlNs16WB
q0I9ma3xIPfVJenqdUNsG1aitT1fhPOnKjInGPTrzY1w/17VDPPCIlHINCWzu7+AEUgalN5pCxtH
hAhne68gBMmZgQ1vmd2pIX4DJbYuioHqkOSbz7CMJcG/ZXn5YVGJMj8C1445rdeKsQ7gpuN3GEw+
cP7M9ePV/XBKH9uQy/d2Jz6jx5jkiteMsvLED57jCvXLnD03uTFc64DYotkrX+nCIrCvZ2XeTte2
t0pdmH0I8qfW1iKVo/Pp8U5PVRD/aWh3tgrAPAuUV46/ZbK7kkCVVV6dwcCPtegeZ8gzzPCs7RT5
uTlre4TpVoHDMoEN0z87i8qUIZwQQ5LmFd33zG4tTI5D3CsP7bZbXUWhKZXoaaRMd7GmjS05XLmo
2JN9G5o4Z8sUjqdmmATRfh2XiRhA4MqIzrw5uZ8lrIuuYOgKjiF6QvZQXUEKAy2iFc8cDPUUvzOV
5RV2cwDtL/6aQRc9kwKsmWK9VyeV83/sU0I0tS0xV2XqvomMm2kAL+gT7/2V02/S1E9Bd5Faxvqt
6B04NCzz2vLsNxJ/Ka11uMcbWZv3F6J4KAfQ7n1SbvodBXA+1kPLERXt9xtaZAy6j9FKNRMeQl85
OemFCkK5rWaOGgjKpo7iiiYVHX1PdwEAqVjr4yUEYRwuRpcGcfgJuY4lplWiA6W0BEMZJrKciQxT
yMxqk7ImQz+rWuMnywDsOsjnOzA1IFuzmOVkSVAfxEZML/KAG4fafI2J6hUzuni/0mz+m/5Z++C7
2NVjpagBCQkEVHePkAOEjnPieLO5LKxaDaKRz1bKMEZWkTpRis839Cdgsq5kUtlSulxE6Z8HXDgb
JHn0Uog6zeCZh7HaqkuG6GaYhMcPUtJPF+qeLayFnAjOj/E4Uw4PzRBavIkg0t8/xxKiyPbQNTGy
Ec6WWgKBfX2fn21eQFN6ZKY16nt6yE8O85+jryJQocgEj3LCdA6W9q75B75Q7usFS4CBoyv11Ms6
mqUS8R7fgKchlSTI5DxSsRGOgwQnY90JbmLTtJum/9Vd8TAbu7mls0VTRqfRm18RyZaWyw+tSbF/
8hLYQfa7BQQ6IKkOIunUhqOFm8b7IASjWdZKbs7nVhhtRJdh3EpUp17/H1kXeDds1RbwHJm34Z8C
i7RQq4ELCe34Ae+UCV+73hi5KQ8udgRBBYz2/cgGie40SCYmWK5qAB6o3FXw0Aeq7cFu0u1cZ20s
sWlnVvfJ4CVqGQ+3qu8OIfgpY5ZqzHge9l/ROoN+669tlA/I/adPQpIpxXE6e4rwLr5v4kx3JuWd
FSJGpRCp2g5hHZvXczYGhoDiXYvLgh/u50j5ajC3oJRhZWCumGQhYWli7cTORnIAguyU8i9QQKlc
LjjBaIGuz7nUEpDnGZkILm5K+HQHRUtFby5+9JJRlfqTxMnB6/tdr3MSC4akv5tUL4mU+CU9A4J7
ZuDttFKHR9abQiPV0dCzk9Eoto19ZyHxHOGEBibLqrgGZ1uJ40LzgxCCCMpcAHinmddKqRqUgqJu
SyA8lJqr2Jm6TQ6muoXBD0aJQ/PZKnKmN6W7q3dMwVcDUQUf6FZghx29AbIrWLV71R5/zgJF5Gbd
LTH2GjU0THDzvrkmeCTlprTcSngEJ9NBB+HhnZSU2DzrUZFuxksBaVWYsqaI+7Iz6UhL5vTo1VWx
MGbkAFa7uLGrFvbz7DlgZrnHxRiJwXMhQbngbK89PgtgTK4vM0Kouhth2eY4GFE/YaX35dJ3BIQO
6pCGJUKheyos8b7n++VsO76Q6ud2KpPBYZ51gdF4UFGD7iJ4MTmdVAwu7w3fm8Fc8DX5wvpR3jF9
HrGUiL7CUw2b7938zB0MdPshTjh5VSWESN1gBspfhMAc458DCz+8KmapbVJ61JegOfaZmdWkQexi
kT1G7CXa/U8KW7AZx5+CEy+V8yp2a1mZChEZzN3S2WdpGwpq2b+DBVlOSf7Nzgg0i9GeRa30zigh
/B8DQEVw9QO/7Omt7w5MoPpxizm1yUmT7+aNCALlyQIffWi2jKFJACucec1OT7vLgPYip2ZzuiIw
oOex8w425BHCFVQtm2GAPJ+Q21kweej//Db1m9wNQgsaDGAlmBnq4mdJVW2BostD9FcbbOIkuyQq
/9deM8R5fiUphfkBwdbPBgHA51BaEFzlJdDeF5T28gg1vcMnuuvNr8jBeBdlAvYMKL2CyQChPGNe
mN+OBXO0b1RZVZeYFX97szZEckMebMNjVwHLTjNa6sr+BqnSRaxojDjK9x2YKNj9NdDBWuPQR5YM
+PIlJ29YHiDVBo5xigI5P3KM4N2b+daMZfD59+59hJyG+Rl8VpovgO+p1NbdK8IiCLZwhgtrega6
895wLXoGllgGstCpxNtuegTFyIkjnwBQFIVQvXs5It7a/M5BBhsotj0JV9af/vC3vnr+SqTkk8tz
3IkMahFYNeR012l3sxA4JJ87o78KmDi16WCBXYyo1hzHyrL2MJjlEjiyWZEietQIOpVq7z0UNgKf
RWLXKim++OnK/tI9mNC1zXMs6uZ40dGQcChtNeSlFb/Uarh2DJWr8ziZeR7C3iIPY2EdrK71dmP/
a7wRiBx2DuWMlrPIZEGELh3qbH6TLzOypiL4CdxMYohvvISsuZ15g95OO4m51as8tNB0Ne39o/Gf
BK9auU7q3TXUDHKS/5SUg62Dewr7Uhcmo4ko3G7pV474Ev+0pLnJ6Pe2YZwbG6fMg+H2rh4KU0Kd
5MlZbv+VtaYv5AqRGQR8sJLBdNIaEM/uxefiv4AVHnZfmHK6pRFYFo10AhMOCP2P+wgPsPrDeftA
t4QV28hEfG90eSWo0yBojbxIOyw30eP9mVylCgDjUpELhBLyboRPBTjJ4udeAeyB/hneyWO7n60a
ojmJey8QmzG9tgaL998SHnmuMipLC/SwG3L6bOVBoSM1sgIBRjpnfuurmQew7wfjvp+IZeAtOC5m
lSXDkBR4v4ueyEBEfWhXDDVo/K1zT8DWhGxnRLXi46FP0vIfCPEF0rGjrdPawLll4SewW05vTqzs
feHhttuHYGMmqZ9s9xwIFfUgRaaRgB7DR0ZMydXXfeqSjjy5G//a326RpcBtKI7mJFc7EGM5h0DB
iPYVZQXxEcQkKnWmQL2UTWLykjwy6nVYXbR5Z8zjiLq9GJKjFsSvMUK5HHnbqEE9Fz85s7tNwtJr
P0ty56wzc5Hgey9IDnkLufy7mp1cW5V0OrfOjSE9zfEufPJMDFdPst0toZi6EtGwrS6JTNBgHbSK
g1oCCudFanMFoIXij11cVA70OQsF89maBzlIKgmY2z1xGo7NH9gGWzwK9ndjalHyVZA1lWYCLkqC
4/0nMLKwHHri9YvR6Xnp1861u1Xz89diCqhefv/NeaEoSij+4pNc2xqUp+wwMQnsIzT8XmsIddPn
4E0xvhcO6kjLAzOaRLxQOcsntF3IMf06CGM5aJ1legukJuwplfz3pQVJs4yCJCJKJFBb9WGmt3bW
os2gjZJJ8N8NPGt1d2HcxshCHMFwZV2cw8EGDQCwHkK5GxCg2WDHo7x8zkGUIBp1tmiNDiIpEgrB
hWfu6eIdMRcAGkOPbTD97bLKR4SxxkHIlDSHkDPZ6RWYenBZKVdTn11pFLRUvffgMYCTQOTI/NlA
DfCbZmeSnA52RwrN9U2tjRCvjvVVyNR+yMyZOJSqgQEcJK6gIyn9xCz8JwpIYJOe2Z8ScBaGUfa5
yslwPqTBhm0yCxeakT75rWsCJVVCTy2Poxy++bMJxRVYy3LxIt6ajS9IsPIDoBNBjGQDwAlCODcn
UI52lo8Ll9UkJGVHGU2uSh4NLM4lZAKitdfQSjpYkFTCm2mK3zSwEQsVx6v4iKHxY2T3F8eatMN+
4k54lV2bGCldt32QcgSkhXh3UpqW11IA/jLVyJjbr21QuCp3MENpz/aX5/EPvDoorlGinvmDJR+v
lCUeI63jNLavBF+ORDe6qDBDQNV3KTgwxSBDDuSTyt899bqJLZiZfShgiNTO/M8loNoL/U9LgLIC
2UKLeytEZoQrsyYshJFK1QFmkODbjt2hreZbuk4MxSlkTMxm8d0nJeNbmcvZvCoqpcCk28LH9tuZ
6CrFcEr56x/A+CwvkYMs+IqWGZiHRSnEL3bSuHYbU3lRS5a9t950eWdhkydiqmG+nY+ohbBWkqjV
d8xgOVUPyUkKr3cP4S6Wqshu6eX4vitBKAMVNOZXJwEzV/T/T1/XqlETTChZIG65tlzKQu8YJWVv
ADpIaSKtk2LIczEkFkcbqbERL5TzmOEWqLXS5pGAeTWWOkjwWrmOm1I2u0d8c9yI/DboUuxAMPhi
BcAl3WhdNeYQYGxNgz+8QjUM6KYZK3GHxRWPDH13LPC41n/GXg1NVyJ6Bt08cL25zw8nSRMf85B/
R44JjL3BjdcdGOD0A1a/Rp+KF1kFiGtLzLDdnWpx2aiTL3itsd+coLAFrBJTp0ZKpdyn00bsm/ps
RyDk0uuZ71OolXnF4SpGMAJhQQs6aD9MXgxMPbUhI2b/Ph19P1ALxMPWfnHSW1RD/NHKv6V97Qdg
2sDnnNoy0OWsMa5fexjydIVHL9MqBkVl9ZAn7kPjceDOUpo57mtu5qnIV0L0+heaJj7n8rvqaW0M
bSJXqv3m1yuvJIurm3BVfZi4H01O8ibSrwsZhAck+FLspRBhyhhz1xrq4b77670/w/V91jz5uyO+
WwA15hc212ZBvcH+bPpX5ui+ejhddZXP91zET+DG8+ifghCvhXdj7JGNWkIXb/peiAFetkPW9Md4
cIjPP5mFO3ULB42/jEiX5V3onjF3BsscgEpNEUFH3TKqbKYP+5s5IVwrHzJ7FzbkogmuNtv+hP6A
nN4ySSBVPWxD8SO6UK+D+nMJTO5yZMBLeRGqFLr8BKsqRnfU9qED1KHzoMWhkXXeGojH6jimCxIc
fXlnF1dMrd61QxgBjBWR5L5RsFINTAJ0/KjdZJPOYtUQtrVdzDzywlIju4QZ+71cIPlgkd8ZNxhM
ZMPFxAV+U/OSzWKZ2c2Tk7U2wKiyiS75ZbxV2EJetB7s/Xy37lkylWgN//Wl65mu715fUifETdTS
KYPg3gwvbdpnldGNCsCUBtepUEarY1IIEFEM1ulhOWWucFJFO0gVOjSZHpHRbTIwim/i4N2EQqLS
EpnO2hJ5fX7RB16UqrA+udK+jwyHYKxKZfjF9jFR5JFvuxg92oRY9lVVlC0PQ6ySx43VQ+C1aSuh
muFdurYjvV9cezTUr7d8hyipNMuUCSk5Wo0NX2kwt/sGxhWU9UYmjtTz5pH4umuEHZ7A5QUngtwN
rKGiuy8goHiWT9tGTy66hnQiZLbP2brCxS1c54jCbirgO7ymJpn8IYAAuA5ppPKcTB5m8Ssygij+
LKvBTtSEWImB6nOGEpQyeq2ta3DdJKZ2y++r1Efx0HB5S3TQHk3DIFEZ/WlQ0biQin9JCiMlX8XC
iabxk7E3lnsWEH3890uwK3EiWNjaNeAGnQrsefyM31vcsQpe8vTxYY3G7ISE8wREz/jR1YM4WWyJ
yv7TlSNrjY5T8A2lLt0gKB1QiRZz/jr1TRarZ6Bxlw38RjscstECoKJ/3e2y83lEXNWmTvJqQ9ta
l+AntGgcRxX2kl0SO/9c6MCgaQdO8tcdv3AiI0hYxuHYIn+qm1xC30DcBn93qnkaHF2VMQ48gC29
O2rEdUOwxtZhJAYVK/98nB9ImWmBSmEuSmPIs/9cTR2TqATU1DhDX9EQerK+NhktRDfluZTDQ8sF
xtqcQDipYIWqMfodDjO5ttFicPiQdgHcY1eumrgfZOFmCNm4ISC7IuhDKe85E9KtZyBd9baXZvt+
EhfjLbZKF3YQz6uMnph5+A2HEa3/FdvHgpTDl793swK6Fq0X4g8NqX9fV50XWePIuFW9KY+4zogx
ir/sL/vJPrllLdeGuqZ82kb0bfsUhYucpAi3oxuH1RBem0T0T35BDjSOMorhp17S+OwlyVmGiToD
Aq1kEKrQDQL9VGRXJokdqS/PjMc46jnA5w6RAceHJ22qTBwKlKVQ2xJagHWdJUa4W5HQty1yWubL
gQnB+Z1Mp4GfI8qqDAi2tg0K5+vZfj6MZHDQEGNXTCJlXMuZlN3lZuv9PbcsxIN3vfj+McveHag0
YZdktKElp34wxdOrJ7MVB378tgv9FGyc2B6x4FSoyejJmgh8TYHXcxe8yqZhyDaXUHf0ghZSoSCc
DGZnd6t8aRrplSaFtPAhJw6jAqOoBWjUxEJ9KGIVrHnrWp7be7Zzd72ID+9dW1iDx1l39QgwFMpW
VPCdu9qIBrfELz+J/8A22nhXs5uPsK5HMXdxVoi9MuI4VSr6vmV3J4RnpYCGRtEwRmb/0f8WE6K5
JuCg6zRc4hC0NTI1ws3VUWt/97udFESXjmRt28EsD8uQwjisgmQwnugED9Em4HfLXa0NRfW160Fh
scggW8zZt/BrpfKFEPEAyaYUD7cX37dJuidYRDRJQw0ARcsmsOBN2QVS89pgKpEgLLPriOY+aIla
Jb7Im2RskrGcjUUsPafLrJ01GWzv8AS43EPIEbT5OSJcUPZPIqsE0WX/fRgx7vIV4F67Nr88HT5z
ai50iZUbqbSF8BevLH8U2kzawdorBOrBlhHWGgJmKGiK7hmEKRd7QJKRqcafX06DiyEcG5FC6yLu
7crcwcNtK/rRBIxG3+mi7DsBOmPeG5CPOxBMIdzHAIkmTnOjcX2UmwTb+6A6im5HLxBg4UapDP6j
OVQHWHBby9tr1qeK8gRd+oCNgcXrRxT7MBE6XGh7bh6YNFxNK0p07hBj1S71tK2RST82SeZeJPPD
OBJvsbkhSDmkxBaFta5oLTU/BJwN9LB4EtaJ4LsQBkyfWAJgmrXLarOAZy/u34KWbrNa2Hkp+QKW
ropxnoyUP/G8KmmWpjz/NOduTy9YQ/WGyFq9bIiVgWJIsFcKZJrp5ezOiIBM6DlHwtkPvaYpdpy5
NBSeS2GDwX+cEFzqk/g3ZUlayY9r3tQvT6Wnz92SV7a+lCGOXS8izEQ4DM4SY2o4KFBqC4uRmApP
fj+3YQh8anJ9mNfykwOoYRU8k8DWduDdttBkj78yJvBG4YRJynJ9G3rZTFov8XcJMu3yIjI1J3UI
9J8reetr3GuI8+y7s7ROZ1GVJHX23d0mx5sVLFT0jJUZs/fc9afW3c/Fi3+nisna9iMXr6p7bSiY
7vzcnuEQujAyQFD2rP9qW2Lig6APGFWfyq3pbsBk/7Ed7WsC8hM/eKLi0zpQCeiLDCkodoZEQ5Ew
3/3BPGy4wWn/Esi3JBFCx9Z0klYZLn1JDgSPuE/9WEWRjc8qtos3Z20bqRD3Mdf5br3/URwOPvb5
D0bW0c5Tx0UO6hITxHa5D/BBThv3oF4Amx0g38+dvbVi/iP47GntDbUbkqDij15N/bVGJQe94FKf
jtuqqBs786fWhlyfXuh2/m3+iodeClApz7mEkAQUII8F1LE8tOUerzh/k616xFjdrhhbG6XzxdKE
b5txpmcPW1DBvw0uaevQ9vuoXimkTKbNismsDn++iB23dQ1xRgIpu7/aAy/ctOoE6+gMmUpTuSBO
RE3RddxDlFz8yQ4RFEulZak8eGmd9gvBpMd+Z/J1uLm47E24iGSwCd7qr4GHrMdxsO76RLLKZyBv
rmBzz+SyNoRE7X+bhXsUfx/+QBd0EHpAlieH3fg/dUeMJo84eYSQfAmGIVMs2E7vjvz6mwHn7JQw
c3a7OIC90enZBxB+6dbKfPJuunEe8C844VL2u0udtN1d4pUpAMl7maYDfYegVkz5jZTCaLZJsRuK
S6y8gFAGSBkbnxL/SxmOQ6CRPSRM6K8MIQJNLJ3fqSermM1jLw1WWMmI9Q4dzbyZntJbzBeu8dFL
cS5PX8myO2GfAjOmXd+hnaafhepW+qmRtJV4Rblek/PTw/Wx9zxFI3og9vo+zggPLBdAUXpMGFJF
lpZ0GPBWPX1cN4J97kxIBrpesgYv63fL1YsVWMLikZfmO43BkGG7PqXyCX/81OPdBEJloBD4JHat
LVD7w/2WHMEC4CSdFf44KuYsUFI8+vq053C4WmdbX+H5SGJ6kWlZMN5njNpyl8CfNJKjcKo8AWBQ
gvQANojhK7Cmby2t/0bp3zOvCpXvDqIjy9ZXV+5r+N4CAaWbe6thql2kh9dkBev0nn3tvkoidVIn
a1/uO/uMohUdTZLJ1dcAi6/feBuR5eKMHRmBQ/5L/LyhGCAZSJgCza+dpHsnD2ramh0ZC2u//7IM
SC6txfwWYIfPvopaNuvna+H+jeK/0Nye3Uc41Pe0a0No1qBZHwr1ogIqA5s5vCnrgwqgbYQTRaC9
V/X/jiCVrVlaabvlWIzcT6p0Zl2qB9+ILLIh2vQf0fXLUvKPdtNO4FWzkRr4VGPYLrx+reQMdCuD
jSlrE275UVJNaU6I1LK7ecTYCX7G5HlbrlS0gc5Y22AMUoeVtVf6L5zzWIcllHd4Cc2FQQIz/nW/
hjwSX8TclEvjL8ZpQWCfTOko6BHugkbz3qKbrFH5cq/AV4DFbgygaxbu8eXht8ta9Fuo4sfFEpY1
oKVx7gVen96jTallpge7RVF9M04Utp/lT/9bMceImvIZbt+/TobS/hOC09cUkSM8xXojOgo/BizR
PMIIwTVuGZqiBRMuBDoErjP9SO4NBSrlezFDn6Q61MrtRB6UGfNQsXKeTLvu+2d5RTEesMXKgh9r
MYejE9EUljsMOKdKEcw9y1F4n+YS2jVOB2bu33SSmNgje/cEkcZzjwkMGm9lE3TT4DWCtDNb0zS5
MDgOO7y7rYiFPw3VEgrPiCHNs9nVqiev4e18MTmigmGuuw8RfchsSfzSh3g90D/sPb0mxmJUjnV9
JEB97Fg6sSQHUia9J/M/j7sKQqXoatV/t/7WzXpKTXzIRs0PhgSBC3XIr2l6zD2p5phD7j4J+fmK
338Gx0OFP/tg3yG028es6fUfzQ3Qx2xXUFGnnUGuk1hqJG8CGpISftvIoTdlzsYc6zERrlkaSZS8
KE0B+K+5zG8oqoGfgSxbVat/to/XwPpPFhlVOHMV+dr2NkL8hfjkpg+vsY5bn6B4MpG4Zjt3j9eu
zr4nr2VFoxYX8evkTDcUmEa9u5kIWrG5ppESEWLcaFl6sx6+uxj+PRbKv9RDhFc6VzVjOugRoDJo
U7lvzaIBO2ToV/SB9sZomOd5BKehtwhkNRAl9qL9zM4lnmehFLg1QsDBiye1Lc7FnSF+UJKctHMw
X1YM1V0u2h4MGKITss9E31mWB32SUmSbAUcflOZZeagI6fm8NWmCzJPT1TaECTEq3PEFadyGuPvN
UOV/GeNqMFhokkXeHTEOc3n8lafQS3C9+no33oXuo5xxr4k35Eyf04lKswuMexBqViqOOQSf5qFD
LyfkV0vrHDUfjqT4Udu6opbWhr38ia4i7jtXqHuYYouHe23e7VjLt8gyAhCCkX8MoeBVAMruWY53
AHbf7/VOjknz5/tkQnS5LlEeYnzNS95aAIVX5rkwzoSEcR6uWBUwBkePIEmibeyb9E+c/YcbwnXO
SqEoInagn2Uk9SAWCJViulxZ42eUWVr37TIOWBpLEv7gMMF0XRAn5eJCCpUtCqTu9XNxvPg81KYv
/UN5mKLpeumMsRGqXNjezdi9lGtMfqrOBV6m/Zb/jWN8EYhLFHB84DS5JJQgJcz2QDLd1yMAEiDC
EUt9HiUwBsbrO/PVCHlMSd94mVuvd8qss/wA8H1xsglbyqZOXRLdrOAY37LIDH+jS+Mnb49ry2FJ
IQ9GET5eH4KZSrvfGHz8gydQipWHkNDrX32AY4R6PzEPOALpnYteRiJ0bk3+Tzl0MR0hmoTYwCFe
9muvsk0/7qK+dH730ZjwKmNksAlpc930sgEMeeAT137Ca5DuyCzXVprbult2EhT/AhhUivVnSdbo
LLUOB85aBUOWTD5cLCPApG2I8shwmIUz4jCQ7TbL90aRdqb1+oqU5PkKvp0CDkSvfziE6iZQNpQp
NjrZ0L+LjxybRPqrpdr4eWEHKWiKRITu6YKX8fNzxBEq0XMpdxa82blmpGlkRmfppDdeQqwioFTC
RmgOMUGMZO+8dq94Ipq8m661/Cv8ZUd1ayut/Bb9p0S41PTkxllj6Ww0RVdSdOjHnEdzkY4p1qZn
JsqCBFUAPnOlBUyrFCiHbaVy5W+6pCBl/15SbxkZQ/MSQhBB1j4nQGRRm4AXthlKcUMcZ9sZKOuh
iEKiSDiiB3rdMwsfCfaBvCXvM3da19FcC3GdO2GEzPM5nt3jrJ9TVI3J4KkfqSBNzVbQ0B/OBwg+
znk8JMPxNKpqMmxVFRXqkOcUs9g38H99F6jnMuiXr4K+mgWL84XHoRtEPx2FetYyALejXVlrWWVj
svj2N1UwSew2w5Pf3hGLou+4weSL2+D6h9U9LzaG8vwJH7sS7xpGbOAhCNFx9BqWsxk5nxBpWdsD
vvGxSGm+4Fj9FwgNEI9O70m+33bURwikcp0sxlUagjrCRdo80+RMvwwK52A+BJgcrVz5k9Lyaeym
wbO2BZmqm4dZsnVbx3K8Az8EbqSxv6+wPAwpztoFU18rfuF6YJ1pF5ttOmWInLPiqdMRlPclncF1
FUQy1FQ18Nct08vjXHuCbtr3cY+V15ocj8NTcJ1eb1KRSrzOsqovzbXpozAij/Bo6aFJtRqIuoiE
2zAq37CBmH6A9W+QL7JOeb6dLnAWGmIgt/v4QaGVk/8nv/hSzsDLU4I45CQG3BAcbgjiHOV6YCw9
l7C46141Wsp3e/EJhgrvtnq4FhbNphZYA0m2TYQ/WY097xPiaHtTvGZm7CxTnIzMpKjbMf1em6cC
/e1VIdBcb9dkAXJnnIkCJ+1VUAWb3tkifKTqkHKraDDWGJr72y+LxMWBGC+ZVk60nCv/o6O+hNWa
uJK34X3vGjmh+Puz2CUGoL+tm8gaUMQG10cF06wMaM9AneL4XdYntV8Tkf/SRr0swawOEW9gBQ05
DPz4KkXx8DxtbkvL5atIz2n/6hbWmx2L2Z2EFjUDfEQDXWec2bgmo4fFs6hELUPWdGuLyLL2eeZr
RyRRb/W4usEQPxpIfVAlz+RZ/aAalh4VFDuPYOvzHChsYdX/O5uOHJqc5XoeE9PLX36ox+yHACsA
KXrCTiTldICKd0uJPLBXa61GidddaCmQ+uTsyn8D5qJqYUdfDG+944Z5J+Pt47J0dIHOoZhumXw5
K6HCC4WwlvCUSIs5WljyaaFzZs7mTSb+ZaheVFFKSoFRFsdD8J6GFx9jnUJuJdZ3VhLHQpmsvMbP
P5XIGxVF+ca2L+OSwRaC99O0irZewWZ/wCIqdEct1O02AybymtOD5al/myffJqUoPHPUL5nFapbL
ZMv5fs8MNitJx16qhpzNrxwzwZ1fRuezl5rMQPEPuLu7CaFT5KGWaonRZqibP+GypfllUPm0/H0s
3xqnuRmsCjOe/nLBmF32ApF5jG2W3DSswjkbk107nqrFzuGVKlJexqDs3LoDZF19pduJXuE8YGc7
8Vjx5TWFob/ouzn62auW3pv7OHouejF1Y1QcNOOfZyodjxyTjag4li30cN4ED21HdhmITC7rKSDq
M9cN24XDUH/aRFNnbEvsLvC/fAOyBHwdWTLrJgbKkGLBqKHcdAq7whKF2C0Bt6yj2Ng6d4fWJNAr
MKz5K6NBqJFLcdhLpMXHV7LtCN36nCvBfWtz9yJXizE9Tj2fmHdA07suUzr2zzgPvZrjqdGsCRbb
0ZIq4DV7omC7k5EUceiATVQ3jF5wPOQeXpdCBJGHGOdDy1tMkQYfx9oVqqdr+bLOMpkQBYYAV01G
RgeRLBvC6ac7oDkg0B17hBp5tJHQ2Ms1nR9yQ2yNHa6TnyeXjpQDINjnqVRmuOynt77QFkNCDPlG
cJ+fhONXa0oHihMu4s3Iv3s5wfnnWhasXLWkbKSd1O4NPjZZkkSz+btczEOgXKl2azh8n9uiX3XI
XbOxsyqw83Pm+41iZxg39cnBhKD2Cdn6B+kIwEVt8G6TCEbJv1n2JRVrerRO31x2OKCakSGGx5M1
EcNtFJ33CL2P8i3NFL5gi9c6MAsXFW/9+Qa1l8SCKAUROwfVwPgMT3WmEEvvBHw/cRrvGWHF/59+
kT1axNf7cg7tt4Z++yz/DiWy/Ql7C5n6KuRNUkGL2H+fLqhrNRTQmR8wcwT0FhcaCU9l8MYvndbr
o7gTI1a1QpWVEdD6ZCE3UyythLjQWYddRjsLL36QXMXNdhQQnz/jKjfKyp6PPjmhMr4GYcPG9PgE
h3V3nQnIip5PDu3Iy4CyL5kiXgKCCQUOzVr6m1MwNcclrp/fYS9v+a+g2Zb1q3/6eQ/X6jqulIzy
DhIeJ5W2yCSAqF5VPgmXbyFYEev3VuAY2br9FGlQEEqGSzLS9UOOjD4wx3go5RvsL920jVGoZPQ0
liSGvoX+2CUQsAXKziXYhBsTVAZWJC5Nhg9swruds/QtzBP9MU7/OYVXcGSxQY2R1ZKMqDPnuh0N
2/bya9TZNRQpEmpmXNM0QRCeQ+pkPow6CQq9l+LgBioZN1EkB01Uzu7cxAS99yjKxHV8hqB2y3cV
KPM6spsbIosQNF6NrhPr5p229lJvs2NWxx9Qo3KT5dKn5tYtz3vzK5yWkAnskkXFqZeHQNs/n6cZ
qBTsPSilRAJDCS9UnDHLD2nAV/YxIMQb7vmVdPC+vtVwsSVDAGNTWMZq/TBJR3AggP905XerPqgM
l8yKQoreuIwb+cFrPWAn7lo2RENrUpvZenWc2U4BA1r6Kyt5e47U8FgeB2EttSHE/goHfDzFsfBu
5TQSKGsZ1A2S+4rWmC/Zm6Qs35yIy1CyjggavjQncf+41p+lmWfmbbm5cnWki5MquYm1gKcBATxO
deFSjmQP2u5x5V5dKVKWt6DEQUXGo7p72g22tKVnueDGucWWnvdRFdUQkSGl8g/dNOVjx2FqfNfH
5jEowplE+mUeFrKfa36M8gnSt1TaPVXVX0SD6LF/C3lEvPHDLLiOEExQx5Fw73JKPZVa95YoBzjy
MylDspnc2Fet3uKsNv+o3gcgl8hx2qC57bCZRuAoJzqUSQ28c8KAk0RWALtj7/DqM+SUFb5Ri2MC
wlM/6p6rg2K3IDicup1nsJGBXBxGEUEGvHD7DHOvCUqiVHTkSYxQSgQSfaoJ7l4pssWIFZXWosyU
h94JXtu84gE8AHCiXG1ZR3Qag/UcyHT16Zcmx11kz0CvxbPTwcndw7lwqnp9mqKwW6xdPMfmw9Pu
IQDXxZsu5n9gcUf2qmTLTtgK/oyxFNfwgDol029DQ1fJbOKgrAy4040L2rK1W7m9qbWeqM63Ye8B
Tajp3yeQdHhxJz0/rn+dC5XJk6xHtsIrpNpSFY623OO2SU6oENwCPUdGBA9yrt12fEJctGQRQuQh
9ITE/BF0yXCAi/Z8V0FkM+w2uNcE1MCUfKQzB86806CYBVq74pPr6De960pW3CEfQ817+GtoAY4b
4GuaAqmRApQjh1SWCNQTm4o2oYaQD9bZL93w71FpRz5dIObOiyn1ySj+jbN33M3h9i1Tez/2LPEo
OnJ2xCa4g6x9LEvv1m7QOx6P1d9rI/DOsu9rFc4wlKy+IEphRhbLpzJUzRiHdjyxCWYv8/ZVytiv
P00zi0jGqpt1kF3vaD/dxMNr2sL70RyO1VFIDlohzjCDGsmFOGFAG1u0yOOYRw9GYZCcchm76RRB
/JdsTYZSs68zc7YTQCgobWdUwfl/nb13L0oMLFB8A51ufgplLurkzEz6/qpuuZSekQhEwVdxCl3H
DYB3bhbiXCjSv8+rJdBV21OuniDUJP/sd1+k4dXTviF6HKyHDPSg1u/bzFqGk0V80JMhfE3GBO1V
YVgBPnWzglWtdeVBPK2UwLwBeATpow+SwBH3U6VjVR2wnqAMWn5AGU4ezHjYDCNQk4fFurSgufos
Pd1xYgcPwoHpCBmvBMSSWIa5M/W4oEGcyo0HMOxsNjTa4G6CvEOjh00amTAObgaAeckVjmRdzNLH
jR+VmC8w4TzwA0JVySOC1DZlX1u+k2WlnyYSz0CwD+hgYDDwksWk+l6UaMrctR8mJ2w6ps3xhzjA
jNqmwzYXL0lU5ougD0QzGlzER6razlQZDbEoHH9qQV2UaVyMJ0bdXvAnPV8JCx6dqIcKMa9xw5ey
hskBDrLNvrmocrCfsL3s94iK9rfsyg1RB2paJ1/GV1nq8jU4oKZ0aH61Io4UGP9QNzDBzjIuhNWt
1ibBYY0GnV7cma4h7JTn7UTHAw/dVgOfYxyEnJx72m4zClRCdD3xKTWxZSik9am4Mzuhf4Xid6uE
u75XEK3GDM4WETcAxaVOriQwFI1g1zqCFjvpm6LhbUljqP9Mie7Ggd1QcdOYKNViJI7QL+ZSQlTu
6/PGlZiliuo8pmquch4TNlxnWAXVtbWWu6wnkihmMOVgYNAwwabg18eUtm7ah6nRRo6RUbp9dOBP
lwPy+lBvXe3N/zV64e75Ku/zjNJmvk3VCKW/V/5MWG/4oKhAl6n24fYgQb8HapEFHnfAXWrelop8
sylj/QRcAppjDEVsMMr+evAKtzNWgBvfkSFcI+qsefcdxzs+5h7aYOkp10eQtfAgkpqUB5GrxOJt
DItqBPoDo/04uEIgtR+ZVsc4Pr7JNms7YFI7K2z9iRt/FokRfsiRrPAEOEtlLLZhV+U2eL5pq3r9
o5jNaeNxoYHFF8cCHOC9YoGLmDRc3bpcQ9FK08sv/y4z+NNqrQg/W5RH4sezFTlJU9F1l+ZM8oo8
nHw+ExmP2oKxB0412QLmKOdLUscBBVsn+16IyD4Zx06KaATszx9+hS7eQQi7LeHa+/WTqM5zO/43
AsUMjpXY8716K/QHi/EDx98fW3gnj89JGj34P2Hlngn4gqv8CumRDCI+XSOp0iT8pVCVRmOqfvM5
VIOKd5HdDetXSMxIIRN9tp3vkq2+eSZSDkigKfkbjaUoOOJoCvkg3542xq4/V6fj1ClG1mZLfKU/
aoi1WFe5+BC/EzXWltyD1mkKLpL54VvEMexIwsOfUn2jZNO44sOb1IMzdivp78lpQPPNvwgMx7Zl
oJC/tQanPt1KaIAPFB4andIPPK6YfGWG3IM269IlR+Eb9qPneHWhxKZHCZ9sGXOqNoN0ldCx+MPa
Vp41BS43bZhUMoV+jmzImUZS1PrrEUYOe7okBVzQQcfxMQS9ZGxrLGnSiFMXdSQ5fO3KmZfLUGH8
RypIMnaWsfPqgP8pKkCrjobxAaXEvD6H9LruNPOYGk/n5p9SYjFXXaOzzkOTybXSdLuXW19E0ffF
PcI4PpI/nHATsXlmTEkDB8M1nIuFjowJQwkJqC0ZD9/9F5aq4ogREPoyPNbUh11W68rzBB4C13UR
YEtFNzuhkJYNjG6zsWDZ/cH8xPgcADleyhJJwJvY0yPcALt7mHC4JP3CDp7v7QCb0eA64vS2GBlh
U7ffiEN+64RCTe9qJeAr/3URdd9CZKxSjQ1/AcnGz2u8GwXLyTHi3cNjhb+pjPdbWR7OEg52u4Bo
Um2BZjZzAwzOFgrRelDUr05IBIqtemXAFwKvtQcfXx4wdSTXt7JUZPoo630W35sKk6ldgqQ8FtF/
4jQBZv78Hvyzx/Q0s967zXoUIWKAU6WrbcoPoJgJOVdPwwh1d9nPttgx106e+THxiG5AdCpwK0l+
enl2Ai0Eb2kCt/DpHLIUdafd5X34WGS8e3zhOLqXu0KqQFCTZAU3NzqZlLy5dh25PCLgfmUP9SQX
3Gx792gLC1GdpYRCw7ME5lSsl+ouNsxQFwBzxTFu4zudNNCKysXADfl7MWvWhK86NbTOcfhPIQ95
5h3TNrSJFk2Yedxuwsux3rVjkyPh3vGwPA1CpWYFLoPHS9wfn4j2XgHIPYekp5GaRnJ4LRJAqUmb
1hSSdaiMvlOWhqqZtO02o8ZEZ80p/ZJiBaCI9hXQc0NL/Jp97wey/2iBWz6wM9IYmK297F4hjPS2
JSLq3xMRPPPsMgFy/R+1MmA3dtXfh6Cx2EcTIExMz/JFKiWa8tdUI0MaeQnFn8oUO7FuI9nHDydT
Nez22uxM/CT92MWRnDleZFlDWm3vVllodlwA//MM6n0Grt9ARuAspoz45kVTQH6T/94Xog0EGBvH
DT4i+mEikXDbTCU6nYVGEVrAtOs7d4sbl1+cOSUsTMKAA4+tH88GxBI6+u3h8HsFkdsHQehUmcc2
uCLPXbUezi7+DH7pCTr9pptxxaqX9FgTMJVkf311uxRPXrJyWqp3LfAQOk8Zmvnl5sfyg6Op94pV
gOezhBqoHcPoCcjzF9j9Eay8CD6YGr0TuySmeqLjw9mPfWs5e7GCiUbOwFHnt8Mr00w3Ay5d9JW2
oM4qIjcMDQ3X2c7YOykCIJ9hFlUz+F3zYs0vnXt00DV3Aijp6/JvJRbmvs5bqgKIftt0X8vzv8ce
yFlNQgCBHZuh3Iw2qymCXyVyw82XIavBQHv4v/K3la7ktnzRer2MLsPuPQ/eiN5JcLIhTTcCWXgy
84zbP+qDRbbsSYSYtAvrDUZAlzSuKF2GInfm52j/hQvqt+ynaVUyWinSiCDU7ClMs8fCQyupUImS
2ZaDm+UCP7ykVHTqmIjGlAkAkFamaHpcsNx9t2x/VGTFdbdl3WtQkIs6mCg/JR0e/1DnAwbsRsoy
6jx7Mvt1rT+uuqgvZyGw7kIP/tbThAN2EnSQgJCFGP+TSG3WpnE+xQ4Pe1Jr1prQgK4S0LX8TQpP
OErcKIYTomcFFW80KrrAc3xoon/C7Jv529RR/IXl6W/F7cvI4ONxURu0dWtn1JFYzr6CXOFpq2jp
QQ2/dBur6rKW4kahpREbBGqRkRZMTuciGxjW0JCbNFr1MHr/48f+1MkW/YdgMB01ihXx+gRx2BN1
6V2j6Z4m710innnLABbelsrppVhYaWs4X5m/J+3YItsWuNwwJ6uiB9O4LfHme5Hd/vhK2/6ctzIJ
qBJIVtmW+67vqNNvj6jhRgc5YpfiZBCukdkMzBWkpS6THiYfU8Eidj1A2Ieqy6f4rtV9cB+VRtIU
d2wGNGt+L8lz8wZXnU1uKW8bxJcLaKQkyuNJYYALUssFABaFmYWM0U4hyUAjcsT0OR+dVd0CuegH
/0S+9hbvZTiB8W2RzaeulLHgefo+ITdaZ0aFbsN/UKQ6cXLtg7LEFsH8MsVp2+luAwABG0LUJv4U
pm6yrdMPoXUAjnLNFZJly+EXN66XliqTkj4ZROtjNdTnt52btKcPPX3G/O7fiYe1Xa7exZouWk9G
Ncg8rDVQMKCnG+/0eCdt8nLJlN95N4BvnU/mnNlut06GxjLyp5kio/dk+sgynGPATL8IR7BBjpiU
X6kgVUTUaQxB419t4xl/Z+EguT40bkIHrqtIRuKgNe54rlt6+cuUPXNtrILqPRs3Wc4B2hqG1Tgi
5DlXhXdst8p8soSqlqf6C2WYwrUk71+FiZ/vCysYvVekQIAS3WjFebnXIy7EeXPJQdw9biy0r9Xe
8t6EA/7IWOvQdX11KBRV1XKI2o6e/nWQz/NZjqXBPe1c+vbdji3Fu0wKLfUQaXkXRrV79jQsOBm9
KOXE4ZQsrtr9Ov/f5E1SgN+C33TfUhJtiMhr9X7g/GMDZwGydmlGRZRpkJsW8hV7f6D6loVdWl8n
lK4xudN/glr6zuus5941bwXj4eYINqXxZKBCNCjmCSUwmEy5K0ThckHS6gkG1XW/hZ78CP2csbVV
AZxrVoxELWI9L8tNIRdvdpoFWscBM0mTO9y+ufVm0go0PTdhwHWtKja1YeGkphmmy8/Fa+6kn2a3
ebd3ArA8OumYn0YVtXXekfI6P9mKrTWP7OsFo/Eh32cY1BhzedNQI4v5n7OZVmropIFK2SitiKpV
vYVwF/sv4VX1bftRN4cdebvvLXUmZVYguEmHWwnLLJQvrRh1LWgYBP+Bxqtst5tP6yKxum8//0JR
n6mx86rcleCj34+4uoHrndmu5rMlSKpjl89D5OE/Qh5jkY7X6X3ZfUrihisrpTOV09z7eNFTe+6s
QhzOuOddq0px1K7tEu2OdRSlA63NMQFH9+B/ZicjB4CI5+aRhauVv4xrlzz0XEbpB+tvpzE7cQHy
HVhd2OOjexEk7X+JU7CBAyLqYOKLBcJiTHU3PVbdb29DGhwQXPy2Wvbmopt+oE8drbhJyznGr2Ex
6e9OU4gkLijWDOzGcagY6JlyVaoW0J06cbJlkJ6Ixg9ezb0R/DCxutc5s9xxFuOHyfRfpma2uQAL
RhPWBUDiiLQuRn5cyQq4VwYnEJCXvCfro/dLoo2TZFjy76PBiDcS0fo2L+GMfXS322nbgOMCUvTM
CHWmOwSwVcg3kELzGJm2TdMRvp1KzM8FjmF/hA4v76JpYfp3nTtJVuOMU4OmYE5TBhDiPD73e7it
USPmzRWoTsJqSss6n5qmoBvTB61W/HCrGOZcnyIcvKx+nJXEkCvUMAcvahiJ64C1j/53716YBRcJ
1SqfD1kcc7tEzgQTaTG8mSui0imfkXJ4CxgoU3HZIVGh7wGI7azhpbr9N3EGEddQJUUIGKwZum6W
anaW1H4k/2qODiWUvjhciY5bGDMJzk0CyOIninJluOpuJZeTfIVTjTetFiluwV432rstB/2LG3gz
ksJl7PA8vNteoX4SM3u1a4XZqUeFfjk8cbohWsLmZLAOp11Dit76Nb4DPJOwtkumUbXrfwpGtbsr
ASkd8ABNiwv2HGHnhlleFxaOJ7bxsYU2WB3rodT0dL+YvArbh4Gme5TA5z8ufJEa06wUXFF/2Zyg
nF6fZ30WvYJ4sXBLdvEb18O+1SUAYYgF8IStRTc38s6qlc5OYSx3LH1REdSPwY4g3j4cf29W4Sea
XD/kh0p1TDtQOd4MZwkyCP6A0A/9haQq6haiJRYYFFXYVCZHa7c/05B3ZwdeS3kUTLLKp6vHYMSB
iV4pZgazWtqFuFw+PKP0h5N28+NkQ5dmhSfl0XRdACxNHbX6/wOX6EInhb9YUsYKsbTYZezZKFZa
SMPkDxaNT1rWJjsNP21cCgvYcE33JL2da1Ch6m/YhLSWEiIfgd1dMEM0nolrgMyY+noQk5+NBo4y
duLLPo/RRHrbvmdHlHeSQn7E4QgYi8qkz1SEpnXlf8JdPcIC2hJZrh1uMbIprLdcwrCJvouYiMsc
wxHN2pJvHnyufY6qttSUnAL2IQcAehKLQJtCCLtVTOaG7gBjuuCkuknlZEPEIOvV23iFfl9RQ5SK
ZQEsLf7QLCWUKV49/qsXD3D1ANgweh/0XzMZ2iJdHfMMqBQr5uFs/D3BoeRk/+oCWDpDA6h3EcVt
Za8Kj8R28gLEEy9nak4/h7CXm8mWGon47M0pVp4ohhRlZB6k1lRC9BXeUTEySDl9KrczH6AmQrqt
6dfvU7uYRQvfW0K0LP9Uq7xk8e6nffVaeWDLVMikKbsH5l+M2PMJQFYfEp2WaAhsUbdueEHq+4kD
KX7rlmRpaLI7LFXq7P/znP7hjSBejcl0mLfepwHTu4bvP0IgsxdVJT/WEFBdkj3C8JjtpZXRIZSb
sirdDySCxjGsxX0L9/VPlzisvTCB22wf/TP8cuP5z/6V6vUlSpO3mA/1kyF4QWApiHHKqxThtINN
Ao9QtzcRe+KW1hVNTxiYXqK/JRZwIGWQVKOUMAjrf1AUp2MCDSISnK2NBiit1RhbUo6tw6sP2G6L
SlotgDLKwz2TrQSyDRZ2JgBSl3k9x02+weoj3FHFTRfFsjsEPdHo4mGay/Ij+b6xgm8JXNWOmiSq
C/9cYH1TBzzW9odGbBEvhczT+GVjppcAkv3WwLdyVf9n9QqC4ctJdGS47nmKyi5pJbK408BiPEG/
lyL/bxry/iAlJrG6jigxd0zbT6IJ4GbVFB/1L8hEpSvRz7Yz8WsCQnGmoBytymRyjbnZadKsO2d1
m4obp9pLD59THDPKVuT3cvmHpPDCoQq61TnCQgJ2LY+iKvCbzYRDBBCcWilCLINP4nMsXqqlF5D5
UDRlzIitfrbS3joxTD64GQeYB4Z4DLQRVrFb8pJhz79zRwL8RF7UszsP/ujhzCESjie1xqMjZABZ
S4YoJwtdYRO9lW/sNfzD8taU8NHJQn57C1VRXUzQt80PBp5g98vx7+GJK8BUy+iDhTLGPJhh07Q+
lsyNlOt9fh0knzKzF3OxEI8C0AaaMco6kT8ZVBbv5DJSXDAYFrnJWZvaT5UQ+mL59DMuu+HvCSdu
QanAYL0GyLEgJ0Ym4mFnva6Udz7SbaGVtxlO6FTChPEg4o+gzR+axmCh4/4qlocTzmlKHq+9CINZ
Gi8476kBFrKpCVnUdEbAELtxY1r0u+m5dpwtv6s1BGwh9OSrjjC9pBaJoCTd8/M8WmuR+TvunfJK
zXEcDvSqH33qHsMbbUce4L3w4SoG4S6LbXEiQPimknDJpSv86vcoDxGcNFEzxiSnImE3eansXeK3
m2uU6luYwlo2QPXqcj0u295fYLuuiV8kQxwbzFEQNKTVUGejOXABThZGAomy2KUKHOfqkaBP8oTv
v6tBPSW9f8ESLi6t+rf+kxtPSrWMjMH+WAqdjv9JT6u3ig37vWl0vxfyQiYKS7QY8nVokDmGtsRd
f79SfPwJ88ut5nFcgvLaBcUdUDyDDQ4MmiKxYiWSQqV9CdOhzT9NU/dgQj1FR4OXmqfQFSGvL4QO
5OBzzpFGCE7sBALj4jecgcHvbjrEsE/QDxommOjtGGjktxFzqP/v9ZMVACf51/wp53+PTpHi2OTH
IO16++1RTsWi/uUkGA/5SiNgMdQAqrAb5YaGfYkpwUZOBaHG5J0KEpvwTbhyzOzTMHYVDDhRM3RS
TZ7kRXU9tz51vAevGgTFp13K2d7nzq46qn68b+CXCAhUNEcMCUkLxyJfxxhRuv9LZ7VVlWshzRNd
MwAGd16HiWQ/5RbhoHHmbn4nH0Yv63DT7jh0zNXni3p2UCa9sLgufJfXZvNR4o12MetB1dJV12sN
gh9vJwZx960KBrKxKoNN4jFXfvO1bgxcwbgrOmRZX/rQCsVgltxDMWFHMbVX4+Qvgn6Y1mF9VTtf
qhzC2c1gYJadSy7cUpvNa3RX8RcgHHNGEdhgYBw6uxBmv5R+YjLaWCUqyB1xDNru+2T+IIdsntAN
5v94Niro9AAMU4xppdmkQUqCmKx+DQk+RuI/dzWAsUeGEGHHNXdHp0rB1Ws/lnmA2z2N0dB6gFsp
2KcdRI47KcOna8a+TwQH9CjFLlGD4XkHSAk+s5baapLfvffqzEbuwHdiHD8uM/abYaLhpNdbeepX
ZVBjTKy7Fz78JiWd7UIEBH/g09GtF1iYb/2sz0wqH/RQvbMOaUy9zll0pA0mI98OuEa9U0qkDLTM
viTLYk4S0mX6f8Gymjjyp7KgI0YbYfhKlkCSHwRiuJutmjKtIxcVqXjOt5zr1tCR+nzlcg++cLP7
71+oWhvK/OM5FxoDHxgM+vTmLVDFV56pvRJA+zToPsmoPJrNO5OlFH2TVy/bK8IBGypi+rSKu0Be
ScHRZNbVc1Y0oXctQaBOl8fJI69xD3HYtT/e+DOa6q9//4sw84ocsDJLEgg5jENr1NQb0C92kAQV
889mEbFzDRAIyZJTwnWgoV9R6AI/X357WWtclwwK9BJSaKxdYI+mmuYHAHr1ZN0Ve7JLEz9thgXe
3jS19rmcjiOfsdwQ8OupcRUhh1rTdBLnvKtOAWs3CewfpNbZarBWK3NHnWlexgyACBHOvoHh9+TB
iIzREMA7/F+QwmmeJe1eN9faQQIsoDRk8bB40xEBgRSFVqxCbVfqRbi/XzzXA2dxH5WICjNQXZho
zWnLlE3wqM3pRSG2ZozNb6ykRdeeSHDsBHgXNMn4NNjLtodEWdjJXUQxzY6BSuo24Ro5NS5w9sIs
amKW2UTbi2zjcc7duJ7U3XJknL9xfQATMB+SLibRlT0FfrZ2g55DB/Cabg4GGlV0PovTeiLuZD/l
DvrR6QEjnfwRvJ6ZsxNh+sDg0Kq1zaiVjRRiz4NW3W8EQaYNP7wIdx/lA4UCmUfuG63vaaqpMdGN
bKRGF+LLxgR5uUeNqkTVFtanPrV4ZQWupZo9K5H4a1gCQyINcVvn1nWF8KAOtWTiQjwmPwniAfeE
tu/MeUTuDcfSxLOa9N29oIMDl9w37onzOdGFFrMwDYCMfBXzZyh9J256TRLb2AUFJzMuxufNGCoW
B5+pW7TScXJ/R3eU0tU3zZzXuEi9AEK+yjvT9nHe9Gic30Sn8wgubNgElI1eG5atOdbcf7dDZZaq
TfLHKpaqERGFNha3veF+2tVcz4bg5Bu3YrcR5Z3HWchP9r0XFEsDEoVem8PQRYdqVnYLucYGDOLB
MhUsO3nD+Wwzx+2IWAF/JzTzC2t4DIb7YGAog1B4/Of/az1dCtvaFodS4SuGNee2THAT6eXZ08RG
v3Afap8Ils/zQhniEG/YEzVF/EuzM2I8F5z4OBqFXddFk1YKDRN5rXyeesJ5gnTetfk29kdJSbHU
TCUnH+FCtdmoX9qZoAiWr6KtwOYYYuy4l+0bAoABUgvFrjxygMF2tZVkkLM8wmn7voiEo7xu/tFS
uATcenc=
`protect end_protected

