

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jAc2elpDF3eoKND1/3jp/zR+PqlylbAiYUxqPEeJkonmmMj0p4wWQxczZkP8HQmv7tuBnI5hb1Re
XvZ7MbtjgQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NcCSQniKJvfmu7+yh3FyGy0Ym5XaJUypJ6Y0uQPsa1akcjYi0ta/33mMsV5QsYvu+JmAYVNroROq
Kz/qydAoj148DuSUxGpr/Dh6K6KFEJQ68T8sjkHECM7M9i1ksK/n3u+J02M+jecJiy0HOyxQBNjN
TYNC60RH/oHr8eLrkFk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bUAhd9meaxo49J9KB0t7maJQYPBZ/miilGsGpP50LlxHKsJESMzras37N6FY41fj0BrwI2d8gwNc
EAnUne+xYMqJWaUJpkx5tkU3/Cq7YHGk19i4FrTEgtDQCfuJmvvnxIjd1KLqJ+tz2Gc83+JpCcen
LoaQjHQoa/X/vrkqv+GBi5yvXYw3CmPRVPihw2cyPAHh/aKqVK9U2rN3QsJFh6K1GPjF0J0zEoGU
HwvENWUy5CJqY+RhFtoI4cFMx4zvZ9LvGAYIaSHNcjGEuPxJtjqEiRDoZaxAPs4fPiQgVWKDuDze
FLb5NkzGHVW3Pw1VKV9puYBInovkYfTC4nb12g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yj/twyTkVkmohkM4L+pOFWHFJL5INTv01+xvkfId4SWEcQdYpyZZSWwRohyHdzU487emKgHzTSTy
GFDvnAvaZMJxmURlvGRprcX/FxMbqrYJ/QXjtyclneLv8hDwZCLiXegIMxugiwW4gYlZjMaOoPQJ
gs8ya5IBC3x9kMPV5rU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tu3CqLR7y72d6lMu0BtbwhwW0WER0YZdVAODwj27MZbWzMWHxGpAy3KeDW2xQMQiri7N5lQ02ec0
GWpokUjyJkcJKOv6cAVA0bMYymP9zM81k2IaifDaYhtB5Ah8VbDj/ArIWXDmp920Nuuu8ntuPKBS
17ifrJikBEgCPNkkESl85/+YxK58m3UimCI0iHmw3WvHkIj/sAUsakbfIOXt9rbFyqcIak6vi6kx
Gi83B53duhddmOvXqbhgzW3SRCCdyG0CtC/tlZjBXsJNv2kpjQBMBZf4BiACBpRjP60jLswfeEZE
bWRI3cRILGIwfm5V+sLTGxa0jiUVbd3TzGM7gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14464)
`protect data_block
pEvtwXSAjhTfzua6aHbKrYpqIBWF2gEAszBMj5icoOwwRqNzOCv7h5eUpDJwQ8R3cyBPKnaslTeE
oG2ea7iILJVHunCGYhrxO++VWVH/TdHQbPpAGt7p5HljNk58QM9zFlGYXPSHcJw7BFHxp7TnXAV8
buqTQS0vpvlaa+JKlbDh8CAl49BV051as2K5O1CV+g42FC7P0HMM0QuDpxVa0VxCr72UvHhE0yiQ
W0EKgSnTPmeDjfXTsYnOCL4ixRi3x/VXWtVQLyD8MHHdSzeQ5cWWc96k+IaoWIyeGKDMN2MZluWx
b2KAXL87OQ3Zi3JJ+2t+pq4jSlkodij5Wfok6ZMAuwWIPkV346OtrISUIIbAPz4gATkRx5aiQB3g
BI2Py+L9Wv/wPBMpaR8+51iox/77occXKpqdKbL2ws4IdSap7KC/3xzdMnVXX7h1oUsEprCpAup9
4kpKl6U7+BtRDp43wHywxH4QZh1ecAZGi6CPoSic+gvhZ9BOfm1cZokVnOXA0CoXRgfLRQwth8fK
64vtLD+E+nzDRlyeMH1GosPZ+LVx5Nzdt/8QsIaWXPbCuQOjAsNpdTTqUM7INbaYfgKbXZQ+3wpf
L6XxwhkNGSShBM1Z09pfLXXdFM6MdMH3KeDNOT8zRSq5dgRIDNQiv8I+/cFiPEk15XbPB9BtxYHG
4sAemGTwstdYqt0TkE5IMvLrT0TgyrgFsnKMV0SZiiIzDd69Bzcfrp+c7FhxY+zcxYiOJaXho9F/
JjTIEukCAK1bQjdhP0/nBgc8fru5ELJSWPb9O+mZnB6K9yro5VpehRz7NzfRk9k7EZeRGizt12Ow
u8sAGrdAFEXbB4V4EaRh+CsGXKIGLPbkpNXHqVgaCPqqEFAFJrKJS08DoN+44bVogo8mt+WxylKT
vWfC7c/HKyWdswcZ/s+ey6H4ICRfI9HhW3YpCr1sP8LQI5LyPStlgrqU2IzlsQ1y3g+/+wz7k7WX
4mNjFarAiK7QISkSLaV4Q2MBfjr6O7oS5k+zzC+lIvaDkp4PccJ7lxIE+nBqKwk9apNZr20NZO0H
5spObZT5Mvth6tzsNXeeAGj8Nm0AhqVMvBv8LS/CtrPJMkY1bowNbn6F34iqUxVPu6DemrFaN5vJ
iL2ICxOUgyy0hV3qjgsAJfOSrm73OfHluq6UBiZCCPUKymxL1wkC8moQwqTMPxObG+SzGa39c3pY
GvErrZ74N9lo1VB680drGmpJNYLtkPlmb6IFZMSI2BKCqwT1ogFPnslPwNWZyK/xJQMqi7ShAvXv
3aAyzEgUNZ2pgVCrHSrS1HlJUneYdmnHeJQUNxqlQbCNie9J/hTmqTYKWomTK+tA2WqzbAzy0zUZ
mAKRXcoYaV3nRKNJMrYB07p1de4Yl0wL8OnUuQRhVIM9S196w+t0Gs8ApejaSw45VKzy6PrU9w/C
y3T5kZpLhIIOP6AK3NgASOXSNCR5jHhGplxYMLL2Hoz9D/BGExfjtWSqIPiXnuEaTPU/FIdmoupx
bI0ArOBzv22d+9NsHEVjAfTL4v3TR8XTZS9/9VepYoNVbH87cJFxZlj38Ens3+tiBQ8S6mT6KN/L
0Pfvrc6ra9+oLR0CbjTgjaP2e/2zV57nZBv5YDY532Q7ufvpTpxAjPhtrehderknsl+PcSIDr8rJ
OByAu88Wq5q7k6ycaDGLsD4bdhqYkbdtPu6VUSxDVsmVXx42kM8Gn3FMSODDXlvl9zAssphJPcJq
p4j6ASSYzj1B1CGsFep9BJ0n13ynuluFNjBPrIWMsRO0sXcGAtrGLY71rQul+K78gT1lQNsJf4mK
PY8CgEikrWimVUEr4HT2NUHz03tT9OP1lfKzPBc0Sm6xincAYV2Dno1/CHysz2SaIaSU8RCMRkzG
8Y1pP04yNI+4mvYo5jUs1LIrSX7u9hl1LX17QAtVuqiaT1juNFfGvAhC/p3J9kz+8kLuHKJcFo2X
+MJvIgqSpr1XeSrMLX8PLwzpVf0L6K2/M/7gpe7XmzXkBP2EWi2n/9wpzPBd2ryF/mqDvwprmbqt
YhYEBMrCJ3OTQWw0odDTF3CrBSn3GfEhYBk6iUKUbivE234MNm+l0iBOhYdcqneOh78zkGuKJzy7
cb1FqWUAWzE74fmEqEP8YHF1nnwdI0AOoQHk5tTETHqE4ojCYsP74E0lSqXeVd8G3oQ+UtPVSsf/
sQFjl9MsZtHdPclKtDRiadW88x2W/IAfHgKE6sZfhdqK7aJfzMJAVS4lwtvstPzSeJJt/NFRcilX
hyTdCVizZf57r1MDl7cMK+L+/2RmZaNGqV0B5visIhZUOCcjuBQ3+stOTND7yF8x5GvdwWDZsZEQ
nkzZK/ygP0T6BtsW1MouAvxJRfLGnYBKRD4RXa8q5LweFUhSM23DCqQK9ucKbmfnZbJy7/rxsflm
MgNNswdDKh+G35iN8oW/TAhrMmovnVrN3Nbbvuul+C24hO1P8XYJyAN8DhSsUJ8A+Aoq8sFL2HAs
wH6hbEE9lgCeieM28zBXpFzgtbpS4I2RRKWoeDWl7IOfMOW2yUHqLufk4+SZWjkkyF04mwpDafIE
8eT+Cl9NW2e7e01ttCZM6LCNJJ6KqOC8nymZownXqeZTGxMTAiJpar9tBbQNOHne8jNaa2XtHvAx
bphDsKzNaDUzYM29WkUZMfd9bxON01JUajD5sJfDr1X2eqbIZPPNmirNaOlWt8VRnA/+9/gYG5or
2DJpeVoFCXu8Nn5eCkiY8e0y+KFbdyvjsoX1cKgEMY9jat+nYsBk/dcuWM5yymgmvig9miuhmA51
RFEIa01D12aHeDZAUgKMpDbgyusO0ATPaDtY6G74LlhJ3yMXq3RxHaK8+qgeONgsJvpGvDIYabfu
BNhb0WXuMHJkB4hwa21DgJj1Yyhi/BGJD68wNKWCzCqnOEHJIMa6wQjZQe4MfJQ6yOoAHcyi1XxD
gCB9WzscJ1kBkfDjimkPd5JWw4pxjC9sA26n4zMdAZlsTVONlTlKMT8up/u3ft31/OEjyzBdFvqY
zLN40mEEgJX+b0ZybuE0VzuZUYmVizuxfo8osp6RmQ2oCa2bK7gDh7xceh6Ue/6flcjNf/6z+Mi9
ANMIU3bPlurXzQikRmLXA3AEXfHeYpCiGt7BvGkjseU/VnTnr6qntPmI5grjL4Th95xCuWfsWAKB
402WJhZUOM0dHmKI82qvGUn26Fp9hDMsm6tD/8+j0YDEQkbws5LbxjecflwVmBvw2B+JxLNBLMeO
1O80VRaX3tHlRDLdUUhS/byqYiClYPcrEPO5RhTVZGb1axJjxCH5N7eocHgLkyH9U3ZI2KzUqKOq
uR1IB/G0zOOINWFxx2YES08CfVlTdHkrE7wQeuWRlsHjTm/3Go24py1uc9dyUyISul4U+E1rZG9R
+6lt6ZIZattX+GVqlFIvYyy2Ofu8T1zA+vUhA4BooI5dynk+Isl9n8SCkts6siMkLECuzAxBTW6v
OXgkF7NLFyzG2hHonpNruNyMhqj+I54h0dOgVJz3i5cPpdkwbsIS/4nsGHHTTMwkjZIEf+DtxBOz
DH9CoPBG9Nlk0yWu4GUXpbH1t9MUL1ygZZYNE2b7lFpgYhpJq7r+FxO79fIkANBlAwiDr85TMbBL
+cR2DhiFu+0hVqv0cZl8gSoqgd+QqIuAcUVK8WLlDbjyUSB8F9ac3ilacl7jreGI/s+36cTncMJI
FEy8EuMx0QbrX3gJArBuz8O3otoNy6EJ9O3qk6JLfY3rjKRKdUACVjznucPuppNYBu3Eta2SFXw5
z3LmUu3Nizn/GzCeCLVhzVHp4oaTlG4RCRcoofNYxhFGXcawUh0Jw0GoFUj8JLbCYrauF0r9knOK
6HG2+3PMZl7dLoWbrabpsikLZwEEK1A26Mlxo9xKtMQmS1A+UbLGPkBLDK3fl/UIpyA2tvSmuI54
jhX5obrkxY5WeR6CAvyfxuzaVfmWSMYDW2hXFdeOiGBHdr2t6YzaUBmkPXqe62wCtCfPnhvqtlHD
dTtxfWafIXoiD9MTFuWHqN/LCeLlLiVroZFBzaZmBEWv5lC8dj+CjVIp8O0wkpKC14rQOdvsDO9L
VmkeJ9fS/tVRQjKGjCfwl8hbwf0SwPL8TjZJARlNmtXGQeL8SYpo9OWT7Fy8uOTfIhW319G+lqhI
oGdnfW28/iUVKrkrMXGJbOSSKlIXDObmOpxerYMUhZQydj6oTH8+1apfJOdnt9HlaefEsz2M5OQg
a/uvrxTaSQBAMBAnEVMR+ZDxb/rmwo77+7I4GmjoG8mDjEn/lGJMy4D+pB8l80BGhB2c4Hp0ljrU
yOjocIElBWdstEzkyjHUuWt6zbSt2IExSEjltc+fveGdrZBSi8lJ5w47XNajt60nEJGRwt2GM07J
OLUeV6pkp5BeeXRS8PH5km6hHnwcMqicOug8h4ckYVw+f5a98T7wg40WZOSCg6RxINhT4nBOSx2Q
aOUAY4ed/R9KvPhMKDXr4k0yhvMqWypsneGZT5SYYKqZF9aOAyD0zONWpZtT6cWuYZg01VWnzCkI
eOWK8JgUh5jdgk3kIKjSJptZDngrt+5FPhanxUpZXpsChmGXXhDoZv+i0nhtdJNsXyR8JSKT1x6k
sBvoBMbtDGTg4Uimq50F3OrU+8Ji+te5dMC8iiIWmQXQXs9hk7JQj/MexWe5D6kft+AIzL1bimGh
PEOcUBFwRsUIRWgjWE6qyE1sbf2tk9vS/GWMgfMQKP+y9nBOjg9eZjn9lcUMzW5I4h07BMu2DmlF
9sxfHOUS1b6QBu4x3YDDirOwrUh+bks2tPCkKClOcppyRC6bObWIR00AIk5jXPzlG25Fvsj9/s3S
FuGtZdtoQBX+9pG5AocaxuMuV+AmFpCFfvFRsbZnO3KmNOTYAP/34RubKa35BhqmCjlmTOW7//bE
gEH2a2kYRSAiwsV5rVr+QerAl9wZeAdimxzwO5WSo6UL85be+SZc+6tQiN+iyn+g/v61rSfl8IoA
vVidMuU85dNwupB35P+h9rmmlr6wNa+TbRi+UfOSMcoio3GygON4IfCYPrVLzUChU2k/956x7U+0
gkB+aKhL2kiHAWkdel8ElHcrbQ8SpE/NdDnPEozx3zhQV48xGUMUrV7X3RC9mFs7xetrawBdi70A
bvZ4bUpp8FhUZwBlXzMoz+cIFeYHFPNDAPkYbxco/Fv37t2wjquy5AvDhOJzN/w2tX+F35Uumf52
gfE/RbWkxUAFJj1V43kzmQFD31Llp+AQp7LUgxnQFfaOg1iSkAi1/QzMdaMLy38EXPTmdvuu/joo
NDEidmWxGT7Q2HeRbjJPQ+zi+1E1RXi26n2eSaIWHYlwH1rSd48ZZjdsgrPVPR8PWftp4V0Fg0Et
Wh3NfhIzXG/T5Ve6MNQjuZ3zye8OzHuAiAdI/Nnugs8+2F2uY3t/0PV+WiFvOE2nJATiCyN6WfiA
Muk4fXgQuP68Gl5KxknN2dgee/jD2wjnjU/kUd1wUs9t81hxdyuEkQAC+3zxJJNVkDXaj4p3N1z7
QHofYu9RlkEXh80L7QYoRmi6hGGvYzxMn/OaGC6cM2bER+OAxTgQs392lNkfT2/3BMUQiAjwPl/4
DCoE2dUP3N9AR6prPn+DfruDY1+13E9Sn3pUxsK7GI/617Ka/2YpQqZXG3iqIjIXqDVbNjw80Vbb
vyRnO+v6f/XXrBrHRvVP/C+OvbFi/UtsWlKkKeMWztUg5TyqVUwBVImiuvNilWjC/8WlwcEaXm/K
IZO/a/IEd4L7J3+SeQkpgHg92gxqTsUQjwVm5OP73G4sbDe2imJn3Tg8elB5jqq/4Ve+Lud73h7r
PXfHOK0gKQwrI4CbJEYv7UIpcwI3CmOpkV+5hZhyskJjr4YloFTPqcYBsBVr6HNJx1KIwUsRpzdv
0LDEhu1ULf2AMaEOZs8W+CN+3xqsL2Yp9kHZ6oQnaGmWrE9/8dGng3AKoLt/Kalk0BSwlG+VYPvg
xZsVzAhu4dOh7Jf41FklzA1cRBuwAcX/+RnfTypIsIUspAvzQnll/rhA7IH4N+qAanGmOH7anmw1
IecXGiMobbJgT5ntpaUDxUtzTT0hBUrvGoadoMsprJNq1DUhkc+2AaK5H11a5XRsnJmWHs6Unifp
8sBcojDHSfFKwwfSNALq5nNFFqUGphZJQA8PiMqWvAId+KYODhjRiIodUvY4c9n/esQpKZHEvcvU
+KFBmn/ugN6f9CjK00HReZiW3ZMzmc2qSkiQ6DFJZgqYJpaxmodxWYMU3h5hVRyFwNNy2rNOI7Uw
kqn2onD8Wo4yuNc5Bawrylwhlr6FSeMv08qboAlnx1g1th4gO0xY2IH6dEXC2pw7x1J1HmXuBSvo
ESP6s4bkOYIwV8sV1HJReL1a1daNBKExaAiroryw2AC+acy9zY0a8thH4J35JSah90FXsdQ4sXyO
X4OIMQiU9gsNXQiJo3hCFm6W6oEcgbjdPIbdhibOClmdKi8k2ydLQbZGyMIHUpftPnRHw8KCHgD7
o7hUbRO76WlZYqZgTesXQ2UP69QPFqXOxO/UIyB4x4jIH38zUKpX5CsuLdB2dwpxNKY9I+cXI+xO
lk0nBGScCkod4CVpNArr9Q8ef8roVjXANLZzioQqR8Ff0MgCQIWbNKlAOUcnKlk7UQsy1HsW6pHa
US6tCLoOMwBMyxuWCy2mPS3VsNUUK+qKpa8jZgbHEYHMHLIHyDKAAtCZE4sHZaHNHrkbYMopA7Wo
EfJgTVJex3+eapzQBsIXBRZzcuEWYk14nw+nBy9qXWnkTrExXqrE4YuCfLx4Vr9ouiRTPjlcifoj
bdkvjlWFXGzdkzajNfdZgsLeHBsq0qX4Ge8F0aSK8bZCCexy6urx0qwStSct3DJncc0fRcYZQhyV
UZUIqv0EnyLWUkIUg1RRVd+4U6b9BZHrynipGlZXxO55TnkNVg2IHLg4AbL4fGxYdXNgl21a9vOi
Kk/gkZewz8MxSBR9EC864xOzDz7CQyc1Wuu0o08GXemUkWZ5/vi5lgj4qOkBxuXoKrR88b9rEeYy
iCZATb8eh6azHDhs5pyL1bYAC7d1uXZhS66Jx1rOnqJuw+i7ez+s6q2Cjw0HKvZYFUix8WX5zJQf
CMfEoc1zwlvA+Ffl9qejO7/OZ8tQdD3ul90j68CqgQO0omiLo0un/s9lfd18OwyXdbi8JB39UfoJ
Mq1splqwEw2mwukSC3ncKN7dCrbfK5FIKa1HG/WC/Mcu5l6RIvImqib8fkC2TjarKvFZvdlYx6Vs
UWg+ZHJErQ4u6jRGcSVmhmNqhq9XRbEDxk/0aXp7Bg9kp5EUk8pJ1f4OwoSWpXIwkWqMot39iEF0
JSudKN+6bxdDtpVOQou4xPcovyvDOPL1Sw4VlEVLc8wULS7m72VdGtdkYOv5SZvigtVC5rjnpdZD
9Or5sXTiO7dkvNfgE9UsJjInH4n2S/ei6fPt0YyvzKo4yn5qIZsfbjut05eipzj8TKkCCMPtwyHy
asKR0ncGUMLz9sByz4ttrA4VPBAIOnvRMaM7PCDBC8XBQbY/TACrn48zYgNfBBN4vAnsRwCzLxgr
UKVETs2HDI7Ry8mJKsjv+lqG6K8T8bAN0T60sKgyVOSqtjDfhvrYjuMMOWMZYO+fdmLsFqFHmnSy
NjOsv/N16loCOLpSUGeIOmtSoDykrkW0hM6qpebGyvF1rj5ZTwEmFGq686NLpdLvud/l10FeVkq5
4TW67ldoqNMdMNfm2cqCjdu9bgFVV2LhhBCYsDnlItn2PoX2R8m/oTcvop72bX78rvC4ohWTA5hj
oEzFCIFMeH6GJG8ZaE8dIHSRrYbydSfvc6X1tfrxvoNFKnSf65vU3PqO1hjD67BwYomo06gmA8RI
/P36jhw+YAmfPExIELXiAlI23ehMJzxAhZRiatjFqgBC5hV+CBq0vTndSpOBFrK2HR6qfc0HucQB
7Nk5bEu+yDBCBXmQwtGWK7SsZJhiG8V2QeugMqgBYiOaXyJWUqIHODzlvuH0PHwSJGtI+uLkDDWZ
/nZaJB0kswFFdpzZL3v60WFDw84TBCfpQh/2tIkaamlK1NuSqkr/bsPiKf4l9N4iRF+pu1UDVyzC
YmzCNQLesPS5cXFSgbPc5cO5/bSO7O/1mRd4WWFGybn4Yyw1HhLVf1QSk+T5P9jk59BbkJ7Do7td
UZIUBu+xNGP8eCKDKhU96ebKGK2Ob646vSAdh2oNi0P+FPbfobAh2Sv4YDP0Rf2D2VX2SF89c+V1
eXBmK5QtsZUCsFUljbuXKEHUnQGX+1gAQkoMwhidKXMAV9acS0rxi3ke/QZKpam7MeTZ6LKA7fjq
I+4+d8tG8NBp7Z8SMsRIdu5gmeeogx7y9aQzvlJoiHXYQKmDcN4NHP3vMuCBrWzZcZ8d4O99Ott5
Jl7TGXZmFi89fyvPUVqNQeDBowa8ozw+r1XVct1TCE/oszGHLA2iotBJWj5rrMTfmGLrXl2begVF
BMQlarQpvHBfOC1QsZ2L1nSU2ddmjWBVK3z6pUtNyxlhka0GZldD38nUmTps7VXoAOqc+K78i+tc
ELh9UO7qoqhjl9OvLlfrrY6mppu3nPRi60TqjoVbMIcy0aOH+jhoVAoevy3wkBiPTvm7cTMUwpla
T/HbGgcQrbyr2Al9pr9tkIE5xxp3HJXeS7QbdSkVWtieN5mwDqVvDl3GXltnu1cOqvE43E7IbNYq
uoR0vSVsF5ACgWLBlvQ3mt9dsB0yuxMHTwDzjACA2rNFepVh3kyUsG5uotV7IiKwDndOhoYHDXfE
EPybP6TNE4VaXNJmFOwAo7im/1KdGLPKddhHkaJ1+D77IHWx8WpilDQQBNiRkCvyhje4yLKj4+z4
U3HjQH2clsdS3AMjxI6sKVmbgUGsg/V22NZ0jV/kUGXtHCAOyZIE3i9k5NVyPOWJvlbD3G7jh8bH
b9uvQxZowNUjrBzTSTtxEIqjY8OinkFxbrBsKR4OmW3KF91+bKQ7p2doP9DNBVB2Svv5wBMrIG0D
Hb0COzw4yGZwz47d/Km3h6fn0H9w1ikmaNDFNBIOUjGPpe0z5BHuJ/c07qTo/Tq1y3jBxu0p1QPT
yb8U0TcmANVkTyjorP2RKKcpY66PKLN7rwHKb9TW/YB7ZqFiIHUHbxP/TsWV3aNfQs2kpm/lSiAX
0ZPnpbu9BZ5NpzpNnq4Hv63yvCbL4oMh+6hBJF3Z5JG5JmTHu+S+ViK/x5vTJlgEkoYcKq+CvKo/
13oGnX8uLhZQgLHK7SVyUgQhPeLOVuK785GM0WzXgFe7zXCZGYElTbRC2vwpI6ZuxIC+rZmRmU47
eUKNhFGPysoXCf3DWaxQCv+TUYO3tuxsLdvkh3a6fFrjPgM6sOp0cUh6T7jFUlzO9IGem2MlvY25
lcu2YZqw0jYC/szTdWoP/7T/LP1uhuFbXC0vspbHZlzB03ZuK0HPsBMQcEXXkpiZRsJuRU1F7Cgq
9QAVx4oZreTCLupY/qiw2QftocqWzVZbFM4fy3nPMdaXpryipJllzbwaP861/oguN8aJf5ZA0PTn
wG2KmTdZxjXtwuaN2LVYVxdYxgVu7LEyWxd7IDYamS1iP+w69eXuQFHEjsVeFqjvNug6L2+IZSTM
8z6wNXiK6AiiApTSEf+FwJexaDhR2A25X3m+iAJPnAGKpu1G/6I2YPkFlG+sOP86Jx7tVFDzbTfB
3qIEBsjHCetMm1W1A2WCE8WnIj31YkTW4h4QMbV9uddP3XRSuFSBUjjepDI0SYnOvCVbsIrB9bqV
buAyvLreZUP1bJHsXUY6ulkFBxFnY5c5F1dD0hgNDl6dH0sic6fKJwKAmBoJ7c0wgKOJDS7wR0zw
DHJpJugAIHZeDBZrxwj57U+fZliE7rAuXi6p5o5/Wy3kFXtfY6CEV3EAoupeEBeAy4UnjuipWQBO
dde/W0TYRWJsvjjVHDL4PXC2DTg9aGljpHO3I8qHk5Oi7LAOLg2TgwDqhCdGKpvO4yoChb5WGgsm
eRTwtkKrslc07Q+NVY3gRc1729vBKRJoHX6qLn5bfV8fiOZxX9XhEhVGYL2RMX+i2rsoldXqG8rK
ecNZH2wSSbK1cJMxUnFG4vSZlcsAVlQL5vKMCKSo9kjlLnb6L/pmu8t3RYet/C7ApakNtoPiYpCZ
8bTYu2bS2prOxsYIAxYFWo8g7yu1Bn45FPlHxPL+X5CqkCyqoaw2uOZRYdAVmr3u4DAOHs3xuSti
GrIdVm7LaJNT8ltE7oBZhW6qG0NVJSGSNAm5fJW9umu08MFdw8WE4kqsRMdHnrkheSgpMO4iHNra
WQtcQvfy0jqV0657cO5zKRJLa/5yzF22cC0njOfFafpdyUnGhozLmGwsq2A9b8tBNqCE7WFx+1Nc
qj6lrlQxT1SRyXFaRsCRpQFGn8L/2qg6dL6yhigAABSPutEzEimZVdRruaLK8YLz5FAWvGHu3C/x
TznXj4vdn3b34Sa9mB8eg7jyvruqWJ4bSllw8dZZy0XYsrQgpT6p85jBhLlzrKJyto0amT0MgF4g
VzkkK3Nk3Wr1bUcUBnT4bJ69Ewcv3q0DPZyJvWFMQdSW9tnyDuoLGFvlkR6kBvqkCid4tEf4oCpk
J+kKVXyiykdizwk1ieZb7K3FKINGWXPz5FlJhWywjff1nv69MLxlqbK3FL2YkBPL5uUjepSzFOr1
xrnAf3Ih6BERgVbYI+x19kAF2ZegF5SUzwWDgej9ub4qJcx2onkTzfl+kQqYEobuSzxl+GdJyfOl
ouOZKqMPvTR8m5uLySQQL3T6qKNdvwLDB7RWuUrycVsvpedTLhtAuxTO8+uNc2PE58eYR8TI3VXi
TQ4uIeh0W55/PAzQOjG1V8vonYknf1rO+QNXT8MeoWqt/rBm0QIhdo4wHYwQXCBOyiC2qAd3ALkh
JrVtNWjlLX2gEnLbdNUA4XkpitKqMK4R9U8RPRvYlLFD4k+cwX05l4kRKwSBGUqQOr6Y1qsup8Ev
Lk+zxfCGA6rSJs7TCXij8F4xj+uLkCBOgzXApqWwz0BXUoqmoCmOSJcBR3EBxEMqU7ZriNwAsI6c
8Z16GbWxu1MSPDGSJhJBxv75zNZzELl7M0NJWbAx77mAzjhQVeD6EEVBX7kBMtXoPojO7MkTksei
lJmiaNVSWbbKp9+3L8J02XASIfm4cvHtvqmhVzZYu12o4eIaaTpqIl/kPdNchY94baOPlYIWzL9x
MpWQ5Kza3G0OcdvkqLUw3GmuS/w/xHtOnmqL9xsQE6M9bqHRiBzH+du9YqAjDL6gTqdQewsnky/3
iP+t3KYM7/TFraCH0hJ6VzsUN3d0kU2pFBKeD94aEeQPUbPb+hwncsDhcnlTIv0TzGaeZ0mQr6Ci
CIZg7ZkYSO6uafgUaTH+tGXO4XD102oE9gBZilsp1VfRi1Xss6h8ek64A8AyP02O4gGw92a11jwA
UAzfqFUD4ea4HIkZYAZTKlc8zyDXFew/EIJ60150ZTS6vrXU/OsFefA9xKcYRF685iybgm2qxwL4
Q1lIKZpjR2f+fz9HzWj57o5tabJFZOiA/14UZHp20QymKrWWzXK4FotzgOjVdXQGid3c7eECx5uj
bMAEZUpCpFeEOCC6DjkifxOJgjl24Zp/4qR/yfA8/O9vymAHXGBTy6kwanAdH8yY8t/imix2YUvu
ipdap+4UYXrdWc70gD+DAIsFUC95MWg9DhFqz+7IMFq95GsyhenaZlAAGN5adNimPy4oFrpUfs+x
hjpqSH0/V/64qr5Kh8tL1LxILZ0sMwgGM7jFd2p/TAlH46QVsd3rYZtGh3BMZjnj0kuj6Ln1lvcA
96Vo5j3AeTSVbMjAtmgv9ss8mAO7UiwpZebaqgHN7Xw8jcXIJJ2xuHPHV6YTP87dJSFbuIjnmJL5
P8O9il0doQCBgYEDFIq4qniuAcAjXRVSssANlEkC9uOi1/lNqkx5x52pIHKwME292f9QcLPFs1QU
wXV5oSC2QxeZf3rNVnZJEzTm9PHsRlyHd7RXwCm6eTGqwFTxY6LsWbjVl+qhLwa8SHLYPqvzKr1+
wqrBwrTjCq8P61LO798rDqP9yAW6LUZGc0tTa5jcb1CTNCEUtt+wmj2slPVEpHyK/D/ZvM3q8coz
KPVNQBdjX9QCmCtdMjdWpwJIESfISB0zFx4x8hnq6FLq8ngB3c7KG5TjQIBrlJPzM23QRaKD03kM
8AhO6KnNj1CMdHDU7zdDpYkYkQjUnmeNTeOrbpXw+QqgtomB+WQFft5HrM3rZ2hvoag8R15GXFYQ
mZT0LX2Y0tf3BJ3GNPdAKfocN8+PYBLoBhKng2Iyj/iYjDdW84rSaV0Bz2QfTLZHoR3AzRRv3aGt
4JPPy4+lL8xgNqP8hJEV+quTf0bN/cNVkU9sFBSCwBD2i/IT+afmqKf5ol5uDvPZxmSwrhFncHpX
Tbfd9NpB3vNpvpXMPN4WIKQndeys8Pigjkwg/Ame4iVJ6ai/c4OdNGKh/1cQ0TFZEV+EeYmsz9QJ
pvMC7sqHNAeExm+7Hvg9Hb7Lxf0QxZCtsusKind7de3g+bEcFF+h9HTW0vOLDop4BAa8Vu8rjj7G
e2EUyneMMZJLtCh/G+iVYxNzudBvmFKFLOboMXv7ExMSHI2gIeo2WjofAW1yiC1oySzswe6g8pGl
7MjSmmNPz9E6iKRQfikhMngt30Z6OyYhY7FwVbwMaowTp0utZMwNuegIxbrNl0gv239ha644Mvl6
v/34WlOqFKQZpJ1/jFtL76nsPP3CJiQWRPTclJyDUV0rlgnTWHMpNhKA5UVRZt46902Pwv28GFap
20GXSsm913A6aMuxyLgLg8woyJRtp+y+WcJ2uFVSd5jS5QHcvQGOYGKBzMvApWmpXaJ1Lh4gqWmu
RBPoKwlnKdkxtQH7V1H96/+fHfLRnOiJaNQ4I6bb6p2PI5C30/9cQMWTTg2pcIc8+at+ByhdZ/2/
IpEXqyoTGEuawlS7BN1soSsr1rUkgHSR3cc13wARqzzGr4M+S54ezDyMBOSn0ShoDi+ivlrkZ2TZ
nIHSrAkQVWlXtSj8Ndu4zkmWShvtwgjOR2/h/3qBfbm0//X/nDCt0MlGDbQtZyJNzM3a8pwRbhsQ
OsMV8ucEHUrHBwNXwJE9lW/utVPhWjYvqVJZrUk6+Hs3VXHOE8j0vSxJhXRPTKYYip8EM3PoWIR8
A47aM7T2mFT/b4DL/dcXmSZycT531SIbZARNZSf97K3eMV+g8Ar54RQ+UaU4TrfZuFgznj0LaVFk
mCauExLuKryYSnDfZV4/ko3lvVrw2eGQIBshQeyYoUoVQY7TYcoKHNup58W3js5t2XOQq1J2EyjL
p8aNmiqNz+3K/95eSBXuSlfIRCOkRz++JQJgpfqCr8i4j+cY45hh3GGDvK45ROTl5wcql882Ytkb
rvEaNAoYCbeXgEo4M6MiS+7uGVNOT9Ba7prNm7KjQ60KrtZ1H/oRjarVWWS9pv2j1donaTklf7UP
IrMm77A2BJ1ShHC1P2NuUyX56B+lKypff5m6BYR/9euMa0Z+WUfGScxWhZhp6qMXoFzbMK0ESwaR
V3D1F6GfJnaIos8QA838E/pPuaEe9lMrupmDD275R6s8sXNOuA7vSsMnPtkeetbsqPDpb0pohV4J
xcjA7se+PSlc8Tz89F/8htTFmd1tZ1neX5Jcwzhp11pMwtaS1gmWA0/ACBSC04Srwc59Hk2diZh+
OKUeX3l9mR9QtCAM1iqDSw7UldY9xkT8xlWLLuiNkq8+hbXzn7fzNlVNFYfHMgsIBAEEjoz/shbO
PiXCwAfK+ev8qBj/I4QItZbEA1ZZFrKGLSgdI5TDBvKUvhIUM6thGQXFwq9qCyRRSN1M3G2dU3pb
s47lpO9LcE7G+vDMFpkeGB6r+rieTQnH2TmNxq44ST6D09QcmCxjm1wyHQY+ErZBHxB6tJRieC5K
jaDpq+BcpC1hCamDGvCVlRIMFd4k9yK0q9C4gaBoz9NKA/0+u2udU+29Fg15NDfRoyMrddH39LoB
RHnPxeh+KCnrArgfcRH2BNrg77DXm9y0XaRQZ4mhP+sX0z1HajQRu/63eO3ENqFa01cPOORiX8Hz
Hbm+2MLDV5fd3d/LLQhy0HDyzhpBckAZN8gwuU/CESMSnWAwFCWrkbYQyO2vImSZT7omJ9cO5grv
RFV7tukFDplkKxkfKQ2KdDUH03DVa0f8v9ggiWblmPOscdyb//BRwPzn0MLIxkkI2YtSlG+hILmV
p4gmO4YzOi9P6KpzTmSlZbxOYHnvoqKGyBH9+wr1rCGeAi4ceb5nhDh7pVj8bBfDty1LNDjiWLrC
lRrWfebx+zBJ11s6Owcxk51LCdursi4T+2h1hH96J/KY+0z1Oy7Yb+Q3BpGh99by1suw3+RTXdMi
ngsUIDaV0HtTmbSWKqMl/N+Bv/i+1GNuxiM/QjcXemoBofqTDgTumJZpI7TipKiDLz3sveim00aZ
oK3C42nZZHHL1Lqkxu0XmT4iFY0GNAN/h+1+v4IqMLH7nuPqUDG3dbE+EriIeCBOLqUFmrM5QG9O
5XE1McA+Bise0iXLREO0SauspfTD8OKJzhEao/r341ixIMeeJcfGNkIq02v5DKXU7/SDdk371+B+
+H5D4zvyb/H5o4lKRVN9RxF9uZt+uZb4ePiDt9HcQfeQ7HyGawoH8hsAJSKkGT8l7arnST01VA8r
fQdGjM29JKV+IypiZHl5VI4zopceLZWYQhgOQdQErg18OMEuMGL2TSdk72cDvJjMkhY1BHYlXG8T
q69lZnqYGrSqanKYOj9RdApekFTmFiBnHjiIhY2XQsoPHUUqE05CcpxtCnaIVeU4372N2x5D5fJb
wmW8D/0F5fXhAvdUHjsJfBPg13EJ7t16PmF4NxtX7BHREk8mrCf43Okzmu5c2i6+bsO2cCxRZWOF
LK9yWEVeAx4NZixcXmC86I7ydUofX4h73U4QwRN5EKQREwd/dM7xvFM1X3Mbex0jwb54Pw+LyxWR
5fVV8SBRTtl+Wp5CPjK/gBip16far1j5tVPyrYkGXcw+6xMa2P3bNbHkSXGR7G9lmy+2PDy8REbw
fah+am3BS7rY51j+3eBFiBqWHEErTmh/HKRbDR9513MadxDewBvkwHlIln4YCkR7EhP3BzhHarLb
yYNICTvpluB3eot5xcx0FcSkWeAcuY6dXDlStvyPMc5zZ8py6EJw32k5dRFHyMpZotmb5yuO4gwt
bXZmIxIwMCmkHg+WbDhQZ2MAuGZ8lW2cBEepvKTonBoVmGwWgYhCT1sEB8zUawW/VKulA71VjtEC
tvi778AvkaprQXCf6qV0/MOY/wYQU+sbDKK6l6HqbRNtpZKN1IWsex4+XuGdXN3kvrCkhBIi/1t1
B3dy/X91PDncQ1T2nOSVD2yLaTfZYZnJWqau+OV3xCyDPZXB6j3pW2ZJlG33GzscXq95CJZyWGLL
OCoUEWj5YUlTzZBWoQXv+BEhEByoQxB/G1mOm1Bwu94vuxa7bJ/Oe5/oco9EyvpG33EHZp7gi7dd
Q6vX6VA4Egk9GHyiqM638+REU1sBYH+2X1kGkqxj4mnT4sP8abJOpCa1alHL2ALifQKJZ7gDGtib
KQuKZEuoe8x3ck+d20435j3I4hoBuQ2fO6NaGhmzB7Jx5td75VIF5QD+rwteTF7Tb24NfuwD3qHH
W2ciuJp0jlpigHQdscp/o4qT4kyK666Ewv1BrCbQSgzKad3O2bxu7/rTfhAHEolANn1NpKr3pUBQ
HcNDiFC+rbTcPIWY1B55BJjNo/hSbSfvoPeS1zn8oOm7lhPy3JOvX5oZtk2gSilXyx8Mzth2oS9S
vniSRVtgLs0f1HYajOqjvmofsRwyOTUlW8J1GoNZs+K7dFxcVCZOl7SB0dA4FMUlTHfD/6CDOMht
cpYwBT1qGQCiLGW+6nOD0CKtpRzncB8CZA+jUdXpGLMAcPqQWfxOmKLazlRWFlMlSxoDNmXZ2sOp
a0gXCN16ZeLj/G/wXW6NxOESE46Rdn3vPbLXrI7hBBM6NELDQKkmUtgFKMa7HmMw2f/5AUKL/1rR
uDoQwS0EXwPkHRP0aBYtk0QFoiAe5sI8CJSVPcPruWZcoU1ULf1dMMDw4o5j0AlrPqSz0wQhBxvH
TsSy4bUX4DzR5uBlIxTwPQ/gCYZI8PUFy0JSNQKTzseHhKSJaNU4ue9Zn/f0+nTsSY8JAoxMSdIM
JOKc29yCVeaCiC+8yn4m7Fkrail9g5JW6oBkTHs4giM1yTVx2R8F7a572SgDH9qLYTwf/Qtnvqi3
AtsHQzSlVO+rqTzDuaqIowteWINax/j7smCPsztabSp8NQHk/lxUxQ7cPUiJUmghTGHV0k5J4Qu3
qwcVap4bGDpOc/1q8f5yz7xa5OuCcj6GZOhorLPdeaQneuwHzOiMklh3doWTtTwm0ihelTSPL+AH
FLDF7fNjqg7mzmTS2qcuo+Iuv0ZnM3qQ1HiawhoFinId+I5wUKvaOlAQGnUprVh74jEyMqlJyZCV
fBtbcJ/HjT0BJW0ZIO8SQcnVPF8xlhuY9vvZTKQsmoMTCNO1FvTf0irTgEYLKFNN/G4qaHTkmwb9
XVI5GnZEFUVJe2O2zANZUmTBRV5N66o6JAl9RuTdHmDmC548vIU5Ttefwk2KNUJZj9YoQ4y/GeLp
clDfXv16TAGLsFiS6YI/cKfSQzwK5x/kX58TJ7LCh9Rnts3a7n1046kXeGi2gGGZqfll0iYK+rsl
327QCKDmnyobSNscydzTyRXfBqsjMXpr15fAU7XFifZBz7tV/07lJkqqX9QuttaEWC500HnZ5X9S
+5mXyLAe640k3cxDfdo0mqojnTlIB6Ic0PvNWQPyfxgwGoaq/iL7aUiW9Rz8qhxhQ8xMGnbumVqQ
kgi3+fu2ezGz1Tj083tA4I1czqPqXoF1J8gRmsj3cKldqvxiVOLQINob894tPY+0tsKZWdxQa9BR
6b+N5S9EF7kYzQcH7Ij3iBtWxdX3vmIDxPlaqtPXe8bjZeiqaaepvsAXFIrFjWNPRDQ7nVlUQCn0
4NJITSlNWHvRTRWGRjn/9M2WeXhiYjPFYGirRUf9iLuMWGsrpWWQx8Mc5jByvHLqTrt30Kp1iw+/
QqtnT4ncURxLO+0PuK6KD4C+AJpRnZ8RsJxHTHH/EbhSgwc6609yk7+xcwsJSaFf/XA5s/z6LaQR
XtR4vpG8j/7ojHiHinGB03mMTcwmq8RqthMnHuioCe78FxTIxLJYxH1AoLzeowXKNjIyvNDYUP4V
WeS78Z0K7Psjs1gUMlWhTP0x0vjSYlfuNElO6gbugVUOFAq20iobU38c7Q3hQijJjg4YZ1p48L6b
n2HrHIPDNyhyKZVlGJUX53xqu7BCbLvDCsUpCAXtAXOlFx8JPmLhnF0oliJrfj5N+fMVXcPlSvgD
Mhgl8LYDMWf9saZdp3sqfa5ahXk/vbF73ggBauBcc43xJbpzLqsS6oy3xt1hH5vnWLfFxam9C95K
ifV1Ea+JRiNDyOhmR4LTrQSOVjg9Tox3Lszrc69dhDzWyqB7S31hP+u1I7OVVgozK4cBvM4D8Smm
iinJIxn0vWhxRjp1fu8oWWFPuT/I64DYyvZ0qbUT3hZ9Hojzpj4E4dRKNBk4DWniObVJ4SObAHW0
SesOWgVqjzbNH7yw29L86a/M8A1A8jsB/TjLEKj1mIhxIQo2cpEp9gXs1DGrazZhkI7cBEsQFCLd
TCBcDfR00XoM/9IrGWQfSFtpZJZGXf7yL5+Uz5NyJrgI9IrM3KWsmhzz51r9tcnjhRLVke5oFCtO
T7levxmYdjzx2I1XMuNz8lIZ/0Xx7P0gftNjdMHEoITzhxGP7MVoNYIf/UTEfT2KpfVj/VZmHkqt
5NRTKBIIyxWF2frpus/OTceiobFBH4Wa/5wriKOi9EGPehvTaOAV/UXXmnUjkFeqqoScgmyugCV+
jgeBEJaYScg3CgclhLN77P8JHEZb5RbeqrX0ORbDrJMxHd9K5mWN1jHqkOwwpl6nNDcGhAkT9NN3
XtO0wXSFOXdLaXzfwVnP4BCV/xnfJQRhjwHUvPaKpx+dTqeEqI3kNgejDlb6RQWu3UGPak3hTx7G
PdEqHmfjRxwlOTuFB2hTYzeD5W9sOOyPDZe4h9pFmsWOkmvk4jzOHo8UFQCDeRjMuzP+0P0GM1X+
K6NnsoJjJ5LJqsB07U6qDPRO09GtBpay0dQ4XSaCiZOzCNrHyi6MuckZ+wX8yRrMQ5wszfW/WG8g
e3DbyEnR6+hPV3jAdz/zB8WeGLRSLfVfX6Mv7d0VQhWZX1PiQByT+O3xY/cPLIx+lfgGr50/MHwV
t4z9j/5IeldWYuduMxwvIx0ce8KVHG0kRF9tJ1M3UedrYAUcTW14qQ9LdJNzJFf8Y9B45U1Hwum9
KfMMEvTPwiqUgshQxb+ixzUgHyARLTw/5SP9uWgFPKrMqATAwB2nQY5qD1m05HLpg6unZXFQikuJ
nLNVdhj8KmksBKyk6i+Qg0BGgMYmJevicM3JnjFI7e6pddUFB+BbNwy8EsfvkrzKHrup+TiUd/5x
5gfWSttDTxQcyGMsgwr/woHAMHg08BL8O659h8Jaoq0pU4UC+os9XLDF8eUigLPwkhlzd9Y0LBda
YxZNraw2cFaT3S4XBjQ99OtlxcAFAyWztpq9WdfiQaIAWDwqkvGqyxPAiQOC60JUqfvHJAVVa3f2
dbnSKK39Nh1s2dF9rQTGWFHOHuHXDDRRxKW4Ub2ozmJF3XynKkDrfWGg6qwi0UDqYhHZnecMxiWN
cBj4eBSO4kHWMpwiMNbnTj9pmAPLOkH91wxyOe9WWPHDz93/cyF5LFTHqsLIJWLTi14pZHdJuFF8
MqkImz534XysK3b5XACgGEk+UrIesHYQf1r27rohnlpyzRqY45cdJ7F9u7f3o0/Rp0IEZDkfQd9t
BYMCS+WRvdoTnHVAG1mLwk3sg03NpO3RSWdoqmo5xo9ZDeb6ZCJNeeWFwZ9WMB+gGDEX18PHHxfk
6u10RvYn3Zafr85PcBc6M6OOxySzGEKj0fZ1JBfaoldmayPMNB8eWVMjDCYK3lJ3m3cWU2+mAdE2
r1erAnRLqxLsXVCma3ufXQPlTqJeoBL3Y+qi31MlvMGCSoL+ZgLRT57Z/7WpPvnijiESt7pPePpe
oGfN2kAMinsC1leSRKzDOg9QXGLpLlDCfUQjMjvKGhAh4ZbpMkhj2Meq+Q==
`protect end_protected

