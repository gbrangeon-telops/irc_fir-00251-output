

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IoOiz+BDpEiCAzehQDaKkNxXycZX6DxCheIbVmZVnOeE8xp7Q+9Cdt/GYV8eq/1L+MpdyADA71Q+
diEx2Z9pJg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lwiDFOkaG5HcqeigSQ6a9WNJOSnncyPnebjhd+6IKLZk0I0Ny6LWNpdm2fV6AG4pFcvx58T5yWEl
Q+/SeuKD0HNAWdTl0b2fE07zxr+edW2hoGXyef1M8toS5SeJjbmVYB+jYYVGpq6G4uNelAjC+U6H
qvBM4HmLQCceNGUHSWE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UFVaQj8UYHzOV/s9ci9b6/M58BwxIhqPdXQ4yEijf72oAEn9ivW6AsDsNzmhpHIiBklSohpBNUDU
0Mva3SAcsX3+9Czy1ShJ5GBV/GrTCNonRWGYRXu6d9ADAsYZRaJCV+2s1kEifAqI6MJhteonJeVq
EumiTmv57LCQxMW5bGdt9ducpN0oI1Oavkx+FYROiHKMHPR5ux/CzqaZUlRJQvJOcmbQcmUZt3v1
KBK5x+Z9B/aBdtf5Z1OOegRTMkPGAdkXGlAX/Ax9OEiQYDv905iua1b8cAJu7PD39JX00W/YP189
CxrWyFNefwoc+rk+siGiD7Jjf0ooGeZDZmjyjg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HK3O5vzCNER9g8js4SKz6W+Zie9dlDlDlxGQF2WrvDyya1unL5bBpCJy1w0Xm1cUo/y5lNUI/ADI
uYqE7JGFvbSauhLZj4HImoydapRAa/ZLL9nSRfszIVrPI8v6qGNzlAIC3uzmQS48iAygYUrq9YT1
qPItKzIRjW+YafjsvhM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
haBqrpdC8sHCosML+5AEE8iaTVrDueP49m0Xd+C16lJUg1YPcQ6EHNHA456bk66+nGBPSp3B+PjS
04UE5wn9q/J8cGL4YbVE/GY5wVAtR6WtFplMeOXISx0KcrI3qk/KzRrP9Ji6/ivM1RBF/A3FJtrF
qq4E0RTyXYa205RDSyJAQ9RjkwZRwEtkcJ6VY2sYCysbDHMzh/lD130AUg9VBNSdV8LSRVpcwCzZ
sRog7YjwhxC0jQK02UyUpzfW4/xJ7RqEZDh6icr8dQvRuVfwm4y9IzcnYLipDLpn1iVw+wPGS0v6
ZJj/N7hNXBnHUH6mTiT5qnqc1qaRllFBLOzRgA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8144)
`protect data_block
9dnhrtwz827SEPUiVasr8EerE4CbugI+EiwAjvDeYTNZ5Uegt8eoLHd3pDJtDy2/Jbl9+mioEbbT
KMrnVyA2H7m2iqYVJ3eNH/htupEdK7GlhaZT+9Jn8txeg2xcBnnGjHS14L1JjpHvcpX8spMnKd67
oaYn3cNGyf2jzM82P96sA3So5i5nd4YZCcBF1/SpLeuLlIA3q87DMe1s8crTxh0FUn595a5/H23Z
VHmjJG3QnV7HamTepx/Jj5H6LmrRLg6DjmjxazGoaJJY8dy0NwoAMD/NDQ7UkVQ/3yo8M/YAgkZF
OU0z5Uc3iTX2zzNVHtw0P4+FSUww2zuolQthYAznUDQkK+5p0JLVKVSq1BJCqkZXUFpnxPdNwOy0
HIznCjckpUo3MRe8w1tkRz9eIl3kgxjicShRm3G0FJJxm042i3Io9cyQL3czisswyK0WWl0L1cBB
iJHsKW6bDBeBKSualM5LFhmX29/2Gp/Mmu5dgoIt4k53uquN1U2JcKVY/MLQQ4+FdwlBpTWz7SuF
CnETkEc7EnSfiJX/diUqtCQeqYVpJV1nq3xAjCw7ZdOd1UUoVB7gvebOjHHeuzQo0qko99LZDtlf
4kwqfulVxkMxg2wrKpqiZTPPy6SRO++xcv3j7vnOpDVm/FTV5XdNgNveul9/3u0qmxUFoU3MDPF3
lWwNlx3WWSP0hlJz87eQrURZ0r1TT3X+9aZbUttF0tf7qtWLJRAyUR0j3i89y7SOkiQ0dpQKxZzV
a2VyJaEsdvXs3Y58JYwIFOLDvt9hU5X1m3KCx39+y0a1CYVkno73Wjf2ttaYp+bkGLTk40EZPI1J
yhjzhVZZk6vcdPzPq5gkX//2FDCO4ccTlqWo1gyTSMf4enQd/n8mqasV5u7c3avO80WB94VPYPKE
lxptgdlEkB8Wj68ZEIZO/t+jUnn9+0i6uHhe0rYY5xDxY0X/PTxsJ3orGUnWCSrgZK6ZuPHzXNtn
RwNZk4Jxrc90S4hHNzaoIkSYmXNiQ0q3y89fTgtWZZIdP6iKcAdGbr0XlDDxCSNDEc74ca5HThBv
BgZFjVSAfn68IKzYuoLZkphRyJ+Pan0k5yIPT55YtVY3yaA0Zu9I4P/PhpjOc7Q0fp9kzpBnmT0n
OYLwbJVCkWOcy5q+bJobqoZ0iqfzyuEQoFQU7o/Wu+uionmStjFJI83UjIhak/MZKgYYO8gijji8
2hzENakp+nBoZMfs58CxtfbzUtaU0uHKuAN8L3TPM1CQblMT5DaZpDs6qSiaCmBMgWvQ6y0XvlXb
9W1F+qogjb+anHrPdze4Xb0kWf1qd3ZQL76x3NsdFTJCccBh10kjgzo/oL2DGvqMIo+LEonZtrJx
D2NL2ngLSXW2rEK6YQ33oQLF2z6p5w4xdAc2u6ZCQXXaR8WBNSMZU0egAItPfzAjN7MBVkU3NAzq
5AnrORXyRew13k+241GNEpM6wBX2+wcEJ761UzC/1AJ6FfKYRiWI0UC38NdE7+HCv991Hs5Rr1OV
v5Vxlm/XjYMCD79cWBsz+ecUgaq8+U4JqzCcGHLbIBLHifbVibi/LPVnZroIixHZPLTaklYaFhig
lKdz2fLNAEwy4BzqcEBjTaxyotwSDkjN8BcXJC7YXnRXKTrWg64IlJbBVBTPtpDE4wkAaweMAS8r
+tsMuEM5PJM2Dvw7k3aRy+e7neIkOi62q6rhVdp2mGuE0+Kari1FuhfjvFPw4M17PgqyDh632OYg
Bfn18mSPVBKA0FL1MPbdC20TrAA6Pf/3iEWJlx/OX7joHeB5/575jG+PvKCQDxU7H1+RuRJicdTr
2jejG7TjsruqOD1vSFAtSTk/MI9sfB/IQJDQO/7wlQ4CdYaPs4di8KBXRsJ3fz12dmZdg/HS92ms
dIEHC8ylk2Bs/fRv+sfYLBLOPDQ1VCjsgJDD2skLso1hKKsO7JpM38+9hc1kRoiAEErWlKCC8M5z
fW9QE7tb+j/PIkhkVUh1VGQjqIzS8okSc5Xi6uyjEKDHySHdNH5IplAgZpY/7DUJGOxySTyidrz9
OSgbm5leEVXGrlE/0ilFo48E7dXyDqboG/vUZADc2JpoXjhZWmOuv62md8UZtj7P71frt4/qO0dp
G4ntdXSSlsOp9KceMe6hNhJzv6ePRvfx4gMW5tZxjahGrvuJaQK6/qK3//O93UY/sukxpS80IJyo
gTRxCbRZ3CACPhSvNXNCPiZEpcw/9eWuBeQ14IkmK37pKVt6sPk6pfFG4y0mOxYkb7+9NrE6xgRm
5TJnGBVpydqOG+ETBjsMcHyTJfTyKU6LyUnV0qaJKJQphurcQFwvV8qdQSmyXTQNf7HGf2DyCRlF
Qz6rISvQkWFGXM2Bh7YFRS04xm+OGOP8EknCSO9SKAGJUvVVffdPWIHA5NZLOBRNPPQf9eZh2I//
sOa/OzGfbf/3Jo1ESlo5WTQF+9KWUP6KXNjZZsBE2gx+M0EIvOc5E9qv/fOk4HtCkn3AV5ePQe3S
gLtNSgDLLoULS4d90PjeMe2D2HBzwQbtJ6RWIwNc/kf818ET0kmGaORVa6MxA6Ur1gkJvneh6piw
3wL8oaV8zDOinkHFdiUYruKRI/KQIxpu7G373Jv3ApylUdo3kcfKQJVIaEZTHRPYqxF0md7iPSHi
sNBXEk9iOpduPFCTk9iRNQjIC8xd8PH2rW7E645/biZFW0tYTUwEsNKvQpgxeQKXEqMbeinuP54s
n6mu6Hp9IMiZ7Zg/npA+lhulDSKXpO5cMwKjcja9cT9VHalUqhJucIhDrFzoh008a4XedERpzWBA
WmtL+e6yIwkeaGNFdstMHpxUIgcAYleJu1WX2kFb+gcPWf5fhqd9NIQOsLxdMAePj8kPfk9I2qbE
WzKlagZ2KOBf8T3Ve9Lukn91Y0lVvsanwfZIPh/dr4cs7U5RWjirtdyJhkIi3Gaf2b4I4Xup77qr
glx8woR/lkCdd9hcUUOB96nYj9GncqPfI6rEd0C7QBjTZBKYSMsRd1FTUlT80sTNIbOh4unOZrV4
8FYyD/XpDYblAZGghKGpOWGKB4YDQIE+UGew1+AKoXCA71MNu/x5YJ3KgyhWd2cRbzi6kaytaRSI
LQBvs3QgBDklkkCjkh+AodTf2Dv4RghtDQd4YVpqu5EclqVrVS6GhqJt4M/+1SSl54gQ9wS5AHmF
S3gRXEP/ktu5ImJwUHE28bfsjk7is83DEu2lY+BF8ZzyU0o3Ts8ZeAoW1+R8m6h9wo2Tsj8zfdh/
1R/1yMos3mCgIG94rp99rtuiYq7bxDH7zPDhm2TquylJUKDULEWUp/La5yQz5KDEO4I9O82SwSkU
jpebiJoRfKVKub6v/0Mfxqs+09TQ8zw1rU3dMNfdnmW7AI4zilI90BouTi+5iZh1FLnI3P2mQiTd
bxJGawuRpMfubPYInShR8VaBOGDTd69XTRcxNZT7HeBlbHmsv5DTCGPAyxmPnoM7Ra6SwR3CsE0n
+LjHxUwfWh1Sx0yZh+n+mawMKOYpWug3+kk0/TH5vhI7sukkZUiFUCsYg08LhptOR4Lt44atKOXT
DqrMegKsb5qoX3cKbgswskx8zSY3JaXYI3/jVHMwY/Ct7x6qBcVTKFAgOrXVBjeLmx72LG+24l5M
O4AdpKL3Ck5336RxXZQd6xsShk/hMSXJOcOBuIi9wORjOHuvwdARFnJj0CtwF27oGyc8gsQHFg9h
jHgG0oHuk73eD6897IAfc5WI552JXgMwabkefSmpzT0DDPmYY39pFOgWP+lxUAA2rEHw/O8FoiNb
Qr9bSN+WQXJsc+tsI1K7cOTUXaJjiV2zxzEWWKJNWx0hPyaKSuXwPTCJnV/cqf9C0PZ93vg62hLc
d97Q9d64yJgOQpvhrgzo113nb49r/7/KxQRGyL3nYqZx3v5tgkXPUhS8ztyFNRpYtpc5+Op1gV+s
sHb83BRqZDQzlMZzpXyW0EOBj/NfCz7iCgzCVjgl5WK6Yp/WsM7fPlkpJdPpjqvLfz6zHAhLOiJ6
YJmzVSlv7edpOWr8mUVvHlba1gYE5sZWb/QlPFnYZLqA5zQWag7aU3RKghJ+p2S+Q3JdTYgPGrSf
SyysJPzBm0mkArB3yy4Vpwp/GW/B4R/uwUvCnm979HA5e69c5db4IB2eOZB4PU3cvBHOLwF2Rnyo
rfpEfVermYH1f7W5h93GkVAOUfBNgjVT9j4CxAJDzqXsRjoBDpTmgv8+lSa3MiTOI5dZx6VJab3A
75fhFpWGXYrkdq2ylkladBD99EuDfhydw2bamjfK1JDGEd6PcGWTSk1h3UtLa+bNSTRXvxkafUSC
9/tGlPzNzW32LxnApO6iVG99uRY28dXc8EdGZSNEEpJU7QuGUSkCu/R0lQIWowsRdO7Lsl5shLlH
FlQG04gYcFHKvfld7fXjYM3fs/yIMYqUEOkQZgDhN5k/uEUAGDx7vs6IvPftBmV2ue/ewsIosbQE
ZsH6i4D2zDrgztPu1+Y5xbgm54vabvMn3HmRKkLU/jJ5EJbnGR4NfHL4IXp/2AEIrCXZIUPHheuk
/wE+MrhBk2OWymBFX1JzDfjqkY43tOvhWUvg6GsCuJKO3Dtjo7oIT7YKFo5HXarhqOuX0xdkpsIH
9L7rtT/rOVwITWguT0praM3hsdFq/hsf2GnoseXlBw4HdnGlKxHIhzYhu968vLLQEdH3uzIxBbcr
bE9Zg5VzD14IWwcFarug7v3JIIn3PDJPgw1UzQL81GgwC4Pv1p/L2E+JnKz9iCZ4gFgeU4pMXPy1
dZHrpLomSDPCOekpIpxqNLNuGrg7b+/RWUU4NSCkCIDiwCDkbULajOpWHGhCYW95wl7E5aNpA4Lv
KJo8QOt//AKnD+LbLLh3d2B+pB0oq1MjA+c9bV7PpHPnNJY9ugvQGayGalBN4iP250VdNMjnfQvh
sm0mlgGIjtV/3+flTv3X+lhVIe7TkKtP5iRtDz/AwWxDvlfn9H+H8LpyvEwERnSjSIk/kDaUt6H/
MXtWAEJ2eVvPGRrjEb3748Tt7yOAJfEfBp/rqBLESSobqcEOdiIo3UOeAxc4jtT+ixsfo/UtCoUa
Y3SRfHSqf4M9fOjhwk2wm2Ma/v1f9kyremEsCgpyhcGSWm68zjrZimqO7PhyGeTUnjNgFDLWgGDJ
hWcE0EXiViU5AFAtnuYoUoDjNOP234lthgfoUbzhyC2c5jjRhhnNjMuwLgzOQ0BswYJtLA53VU8b
mAL5ZALjWTCADP6rYGSWXHj+bQHyapKw99HNRo5DwSrvkuLS/YsDyGuyIxjpsQHDdnaAQX2CSwEU
aF769Ba/ksE3vWPFHLWvuF8LfxLGzLKdxs5UcrpyI8yPEM0XlKzgeGtTnJD3C6YWJIkz0sq9lD+O
K13Yl9dMlZPjuzzjRJYrRNwKxer+xQf/szZ9IxqgQRoesnpWVoitV/VmYUPhzaxZ5XoCwTA+MIoq
B9rULq/exNsUqc1kf0imO0R2MuWyaVrZdZZM+tLd7oGvRt4z3+yIHhZJiPN8ZarDlrzHrLQ4dVgP
lP8fpA32P2xIB5N4BC2gc+vd4jmFjkMku22SEI3YVsZ4xofgvksFdf4qOJZSfXj1Mqr6Ch8OJSN4
0VF5UXbVKzR0slodAk+Uw/Jsdx0nj4kdu9BxTmR7lCtbIYEN+KrnSak4QRjpIeG3t0mV501+SgNF
ycu7w+99+ippjmRi0F549NkIh68X3bPBdWGiWvsgnWBAmZFYzI2PnZzIFr8zmlksWkoSVYTjlHDf
rDIfG30zDWFrPOqkZT4ClYMBViuPxIAwxC0P0sP8hSj/ax+omW193yiELf8rHyEHmNUZCShbmg0I
Esaeyd9gDPTy9lPUPXeX7cPnKPvEjLGwLS7GUFchOjpaNiHoc+xMgw7Hk3Ze0sjQF4HyjBPN7VdX
2KaFnTFzUjZNCSNuBlIZobeScZhKRqbUBG0FlN+5V8E4rZtUoRldkOPFkrPQgPuC4R0NYI3rR06+
H9Q39kyCrUqeHEOvdjM+50C3y9SGanlGXp7J/o0oabDZUptYKplI0y2OVE+bOqt3qyOb2BQ2JG74
VBCAgowzdPar7L6gs4jXu6abv8u2FcysYUZBa/IhXSZMXPNVrWNkjVgCTG1JiyzJNaEcJPTmXoG3
h672awsym+XEySL5pp/hbtu3FQE+0+PRyqEPhZlMJGEg98rqPmmWBL0/SJu/PvgHhOOkO3xbI2UH
x+rMyx5AsuXqLdEUFPc/1NPiEHabTO2iiD+WIaR16YXHktH+ec2GRBu8KJp0Zzcl8mlrF4BjtozB
rETUAOeoztsLQpJlzC1ZVWi4APAVHpNx9w1AXQj18QL0uWHf6WDdYf9jX7FaqtpRDqo4mKWGRGyQ
sMPR+V55+Un+FO9c90FCH7Zfm049jWRCG0lUaDGwzm9Cl84LzMOLyCTUrrzzRrtDtGUP3auzCdBE
6nlc73OoouDUR2XjDxT8uXQneURHFJAnE965e8WqvYud6iUYGWMylzFg/LjbrdotzQYs06TcPm29
M83KR058DiyX3cKyXfjI1KpKp01lxGNPXvjphbvDsE/wX+A73fsSq+hx7FRCW/zvFBW9dI4Ify11
W4lEYSc+oR5w4h2lEZ0lA3nNsulDNlcHl22D0FzGM8W0RUVzxWpW+3kqTJO1FgANztcHehgr0qEw
GOZMUgqFuJ6ZP3ggD6sX4ItKSlf+Ng6VVE8IrufyC0FSXcNPnrf0/Ro4RkX3q1oFS7qQrqcI4bFE
6sMl3oa8fiYkEPPrFSkLTDQCZBmT1C6DsEpBICNwbAejyVVrcj0rRxW6agCWa1MwCzZ5Zz8R/IG8
TEFhHVJuDwN7w32+NHNfV6b+uOOLCNKQ6NhAFm6RJpiKQO8/rX4Ye/nH76SZNFXiOdk6C/PHjShu
ZKJSEsfGARiLijAK3y7zkJy/ZrBLYaziUlYoJGOvoawu+yULs7hf3zr0OrUSVvvg8ggMrx9JhphW
NxXg9IJoT+MezS7S2UW7YelADar4swlF8TuwVJSWyVibWWrr0kyBfYLSVsfDaHpMJRtXEDswgs+p
BP2dOXLE2QygChPLK4MNCC1fuRR5I5WBlYtSDRHJRNNoZGwbPAntuXnuoZ4ar9M6HZHD9CZ5kdCn
ZzQ41dKAzTfhnk53gaeQE0zKLTRT+krPIt2s7t+J/BUxa57NI9wqvXwUF2xXwJnFUcp0p1WNgdFp
Q1YH6Z1K9JaafsFjt610eXlB3QOokO0WpOZ9MZ0uec2rU8Cwps73rxnrXlzPvJ2TxOVkgSxsUxnD
Qvvz15Vt8P95+V1H5SvJRhcQlg77y+atH63d+DLqajMTKvOAufOMU2uxjSgjtYkkU47+ItPbNQji
mgxCB9ygQlORGk6C3jxaPQemcnn55YcRGOAIyGBi4kRCBcMYCrureCt47q+tKBZIdhfm056u6Dqr
FkiixwZSHM1Z25KT6cHn5zHl6T9HaFox4VQfQIJI982Sunbp2kcoKpGXvbxuKiGYdiQx8OkepCto
DRco1hlTGQrdIvL9Rvbi7/HkNpgCqExDrb6jwGS+Es/m7Ye0EpRE2I8dmCkr59pZE6Drkmh24la/
GyKH2x2NfsL2jIbmgIEuH09ZXSHuoNSfIt5Lh/Bk127f3WwblHq/QH/rugiPIRt2yGZDBz6S+xdn
szWtjK9fwR8SeVVDt7JILCQS2Enrdj0sgSe0AxRfOXpZ1b2T+DenzL0bTq/uEgLegZNyJcpeZB7J
7w43DlVu3hjkqXAT76ih2OsTpdgZiyGRnx5M8As9l1n3c/RiOhtaMytm21TLXD3yMdNRm+idI4zx
opAKbc0m4ymZZ+YZr0QsfMd7OIZSohyHSfu7ABaxYptCRWFj7XzC8KCUXSDVg5DvX8tMs6YmNn44
EcccEfkp36IgGtur0tpdFnKzYB4lpTsLSJ7YZ57jxR5LpJk7OLTSpPgBM0xVuBIK/RstFkojxVgv
ZdRhsZuOEkkQe2Thri6c2Uoh263e4H9ixKcWtCh2WQPM/7H2xei0mWyLKTftoM3ttyoUuxn0PQOZ
79wa0DGjwFbsYY08qopxFH7uaz3mIuiCJHhBuvlcD+TE/1X/oqBHK2bkdT7tH2yVvywMnMH6U/ee
oS5EaubVrvquQij5vnswtH4wHoAQx3Dp23fa8Z4khlZeyWvdFO2vwdjBj3W6q8gfrW/eplQZVZZ4
EqpkQTcvRJ1ezi8tKilwNXNz95xNrl1nv5NV+JWC9LaoO0lBLnBnW1eo9nv6fJXLshG6MbL5mAo6
UgZWEaDm8A5c44ph75MomdoPXpx0cMJTcn6jOuXfs3aEMnuo/RigElzpl7kgL3QLz7ePdy5RFCp2
aSNQXqBSqQKL5t7QocpQwoaAiOGxrYB+N4lW1kG2qq6UXu6BeVc0fBzDt8W35dI9E2KYSaQM7uE6
rMjn5wG0+MJWUuFicxvEpn7gISHFxThNfXcMemOy2HxDYssrvKEjOFnKE2LOJaL9qklP5tjB95Ty
5wcWS4G2wVgXJx38OdbOR0IuVtyNxvWg5qj29mStXMAAZqT5/jaIklSzH7cFFOeaK/E9LZsG6lcf
WXJZyxvzI41hYmHGcIRAO0V1HN4CGt23aEyiizQJXnUjX+6SSKg5cFadX9quXQn6GBW3rL3wBF+V
73n46pH7w16jOPN48t2bmRzWDjhRcNLIjrimzgFgtSshaGgTPLH4+H18UkgtSS+lmiCi/+m4x7ve
OUe0X7WMrMk1jQ3Rcj/3mnJwxtj5CP97/Nd3R569RjgMNw72gkDXC/9MvjKkJHj6QDVnB51ESWVg
uMOCP2GW+csbmYA3kAbM7dHuuOG/02G0tBlOglXtVvMmn4CPAXUYP/LnXLDscqzVO1guFaHCmPJg
YdGiSnE4EUM3Rk1SwmeQv4BSa+jHZAKZCElBn04Be0l3j4ePIEePMGULPXQGYvftavR2Kc/OrctA
5aHwzu9m+Hcrh2Z8oRp6k7//m3UbVDVtVITVSIpWE3KzGgmKldg454jYHLs01iYpRoT7G6iyrPbd
OHULA1r3TRbCsrFp1Tav/sP8YaOOHpX5IzXWkyV8M+U6QM3YLvYDN2cAmxE5mNxvBzHMPGYtzjtM
2xeWUkmqARdlA+CZMWh7yaJNYyiKFe6SWpq0RZZEiwi0Nu/QipLWc2jM2d1/QGcU3vOUk1BRSnS4
PuxF2wn5n2BHgIzE9YEbNGJbG8JQqv/dGiDfm1YjNe0LHrdI0sYkbocpWu2VcYKMPLxSLtXJ2NrR
IDO9CsWYJVjBtmVtvEhwIy4MWofMCVAb6Qe8Ok60v9WhWajQoW9jNLWZu7KBG4BzCVSQs9csHwHs
t9H5sWk6KROSpyDJLFfgO96fihAymFzxAfexCtXyO5XrVHtTW3ZsbRuvMCwpj2Z9KQ0ABO1wIUch
DqPDHKfcHF7fZ4h3Esym2l/lvyD5wsmK+xJSYmvsXglo6rwn/gjkFPgIxRyTac1D0PPw0o/+9eS9
hK0vGKhV5zY6I5+hsp1o8LXgw9NNTXbgOoDtIMBrh4uaSHe2KBP9nN6MosQTNzO7IarIYIxpUM0I
y9fTVOFxlzJScyXiFI9BjDJ4xm839d9vnVJNTxfQzpF7PFABi5yaw1XbOqLNJWNLVZ/QOLyFwJEc
G/5yQ7CD4harZXn1OiGxl6a3K7XeAbyqpaSsAsemeiI6AgZO9dbaui8uW4/DsH1yXnrTYK2W5Hgj
5+wy9zSO1I761sM5PACd6sSoHq5tQmKWweayPEYb36N6MDQdIzoIyJMV8SmYhAobET7//EleklhY
sE8b1tBKFGBm4OKwodkeCUHSjLHoo25fjKS1WWbbgBlkxekjuhsB3xHxPiLNsRqt0Scd6xK9DgAH
fkbpBe//TJB4G08WnZji2BFTNXU+5aulBNeyOk4hL5QeROEsqB4/CVLJONW7uKqadAlTQLOPc37n
vJJOTrXEMa65wm6hV2aBsgABsBhgGL5YgumEIIlX9BEHC08qC0MzFlEM5gUeJFJdfnRry4j86L76
sPix9QLi+QZSDSAvWb4wbOUDKXh/+aRzDr7JdJASmwz/632pAs2/LWxQtC81WJ5LJEyC6i6iO42I
Tm2yAW9H9r4jtHXEskSGv+XSRS+HYBNyCz7W89jCJKHsCkHi5XAzUGF+4tyfvv8P9MkudosF3c47
aCdGNAHCyXZDzKMUrQ5lWf9uNUr0mBUGMO/v7lQRipLIGTcJD5L8YlBjDaJm4PF3fcnoZ6CWT3Uy
GpyT4Hc9a/vuXbs3Tg0WO/yjvlEB34Un/UnDbMIelWT9XWAGBlfqWx0OVrxznxZzDymxT9xfKtt2
jTguw09yBiRM9DtGnlpMLAqYT57wwnu2aOmscjdSLdpA48Z80dTl81pFaPz8WV/yV3BAqiQqjtLr
jV5QiulyYdChve175SAjHxCBgu4T7cstVz6Cvs3GoPThqtf83arjgFECOBQGxbaP2ZebtuEuzICr
ndTg7a0MPkzqa2WT9y202FBd5P4sDRs6rosTYIpdky1qn8zgk7j6oQnIUDKy25AX7I6cRLkAKJ4B
rfq/KNF6mmglPqqnZoOd6g+jEA2f5evnglMWCHuVilnUjjTo3EYEhEZ2X/SMhxon+06xCYasgeeZ
Ih4gm/ah9gl2jDLiMkrJDSRhl3RgX8844RFRTfXDH9xQi19TYpyqGL+aZ+7M6XqQI+SEjg566/As
iRhirN1mQx31vTymzHYdeoVkwajOBqznEo6JUVfzbpdmi2Kh1JSzbieFPDQfxhNW6KmgYjubk63I
6+enVfpZ7703wr93SLbm152HBtuWpNsPCD9J8znw7Ps2wL5CA87DyVFtEbSiUZFJ6XU=
`protect end_protected

