

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JEmZWuLCZazscYOT+xp8tQcgcJoo9xw+tt17VTk0Ee/cpOS713F8lYXKKz7qKA5t3FpvNSj+LwOT
FOkmwv2alA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IW+w81BdrtEdSrXT08IyeN9itdwHkCyvXK5q8xF0K0oVKDwJZ55f8rUD3UDvvDXIcAjvU+645JL4
ch4hQtC7Y2FokqIuMtHZi7cNrCDQXzP1bGPJjMCZbuYkodHhhDFZq0vnJHG5npJwjfiUcFOs/BD6
321VxRY2LE90m/fkP5w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mn15icVDdA3CjzJnkJvEX3d4TytP/AnBNj79QG+E3lCes2UF2pZhqISOBY2uufaQ44Iz0NeMSC9n
+tRGbjECz4+Qnwa3jPWzed02j/IF9RX7XCNKwHKcmJw/yHIa2jnhfXGycV+rW2BTSaOcvd71AX8c
xlCKhnyKdiYayGwfRy3hMXLuu2cdwaKnu/UJ1yLUb2SMopRlt3x1/DS/ujprioIUaznXnUPKvPI+
tY5o7OvS4nta5AxgAsVoz+HHq/K+cZ5D10lOXIDOatM1ESgBnEMFZa0ND/EVV3+YXn7orwuIkC9e
CVEV4WCQjR+/QOWg525B6zV97OAe2sVt80NsNA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3K+sUBRgBhLO7z4XKbbFj5Dm9dnCnLXJtz9DyutJQ/EYt7E+7VQGJ2l3bkkVJ8bn/YxKZD+Rqqzl
gzUxIUqSuvPPGmd3z16szdtLqj5YRAEZVXdNbeQ6P/rYfI4kn/0Qw+0hS8K2lRo5EQLrCely7fSf
ojGqs698Kv3dVxOM2uU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EHFOd5L9tY2zUSTwaEQFpNSik2aT5WpldK4px9GxR5cWZzjNzosBm4ckg29GsE3hW7YJVXJwn2ft
qvaRBZQhqD+DF8s0vynZ8IngOkOgp968BazD+XmnNms7D3n8pwwWq1DBwFf103zHNgk183z41Fww
ghnhfPrVLnkJtKMArkX+0VsxpoDgdODsv3fsT7CkMz19ja8WwHPQXCAKUD3p2rptjKIU1LKJfHEW
xgEccgVmdaHJ8o7kwvdgJQxZnf2Fl62jKVF8AJCrqXWKtvakZCxpEqbYNpoJ6R3Ns/YvtWdsZkRH
TW3+uPSDGYDVS3Az7zcuFIC462DOhpyBpwOGGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31872)
`protect data_block
sgz2gACFRtf+gLHVSjQfW4nSc7JTFe4JUv5RPHcYlPyDU01eNugzuBfmWI3CJCY/9DccW52zQrZL
SUXgfgcTspSBCoZK8s/nA5ej+N77NrD1yt+tjec/YVCekMyg5CGyoBH+f+luqvHk7HOMbS2DAZ85
j5EQX/Yfv8MoEOp3cc5ti2MIQgkL7tYXjdU8mph2O6VQQvRdAXWbbiAaVCMt4abLCQmI4ush8QEW
7ND8ResrDhd8zpnylcTRJsnkqrOJE1PT0oWzpbX0/EMWUlOAdcsMPIZ8Y36obo4AfjPQDl0FSb0y
dr+9QDGzRZkMdJp9L8otLKaCbqHz9zM5QehoIEhuY8U98o/pcD4XpB/HSHGy7BW4kKhU88i+8JTv
xFXrGwwzYckbUXZdHhkIDcAP5et6LoRhaDqX+GEhRPMrgZb/bUFmOq5Of50HGBT10XIw0olDwnIe
BzAKl/ZGAOFYeqiInLFYpCawoBQmHCdjzt/G7xjgGJxJ1mJCwnKDaUdPA/H859HkaOkmzEVWsksR
l04ViBLoSqTll2qZNgmwKtCuWEVGi37JfdOaa0/+n8JH2f8vUrCwwimlYAVmXCMVgyKSMJANJP3u
6OOVxh4CnsRk/MKZl09mNb+IIzZMog2jtsAsjZMu7lRWLkZk2OEK6s2lDNM1EU2iZAKDjCNE5YIo
MuNaFzc4bYX2cz0YClaunNfU79RpvBiqHXqHA9JDvN0qVSzVv1NqzuZyZBk+aIkVhm9gbSkhxjXz
MimG0kebBop0HN49xlBVhDGmtsfWUGOkkC6IIHIUr9pCuiw9WdjDd5JVFOEj7ANzDGIbJIAyzdvz
FGt9dTm6DROB4rIPZEzhWSkmBkT+2MU8O85ajouSZLrPcqK6Ixm76j+C8vpYrdZDSjNqSmkGwn/h
dgCavj6Y6ThnMSmZGLBPjKFMNfXdbD/amYOGgpZSN7YStrVhgGly16BTBL0KvYQ8EaOG9GnQeb25
SAp2PBgvlcxV5oBtqIPOIQVVB183d4u5JPVo4KeM3iA7jg08oW7wJGc3b3NULJGNfxwKPo5VVtbD
mUCQ7PKq7z6zlr3KO9mWJT3PhSIhtjhRjUv/N0ZdYk9OI+ZuKW8GqXqA1YHUVF6M/Fa1q+gBktKz
64t9c0stE0VUroiJNpjezqShkcrdCtSpvyZMk3DzKYoFMAol2Fx1Ci9qHKkZui56PPVA/seOZzIU
hSnbgVqIUIVYbZtg1EF9SH1zpxCrb50e2R03VoX7bBXKnyNbMmNgQ2nq407a4C7esdg58luTAljV
934KoEpTFxTORwtTRaNqvdGCCU+Uy6hySArVNd38t5JqgOMHx6i3D19qKCjEQxfVyGjdCwHOUEbx
1anN+Dd1RjSVZ51lSagtnH5mt4Qe1PKv/NTYOKnN7MebaWVCHLuFn+PmM3ApgjmqG9UOrBH6BJ6/
s59hl/vtWfMjKUKJwBAmCrgCciJBrsGuKSDb+aVCSU0Suk/3jNRpptizkOy3to3U5tSNJko11IEG
0vOHRkcJD+v/kER9fHuVUbjO0Z7kxZOBDsuZoPJWo2xjwo6Cv5lun+Nq9cmyxna3wj3yMxKBZpEg
DKKc9viSPu2knZSXvav9hQTewDT7xQhI//P/TN7aqD0SgpjbIBUxowVlE1j3GhBrQbm4rOsos+8w
EVNCmyOZpTdbr0FBliaS/fD35mpjZoNCb1wq9YQy3ua93K82DSLZ8XlH3lx0yvARh9eSC3eK8isO
nH6uuKnhQbiDVoCKOvRAIMKhHGJWXXJ6/hbDD/zlcFbs3fvtkLGE1+LIvKWBLVOP/Lz/TYC6V/YP
a1kTIGEyjCdWKrCCVRptIofDF43A7BLgrXnrCS473ZkEuyGYabCEU9nIr5Fl5mItMI7xKCzXd0HP
OMPwdryF1gfK27m27jXfxt3fqd1EpkPZ0UZkXBvOjKNqPk6fX0ZvqTeOvn1qz5U/Vu0dzcDXw4h6
X5cYTaMj5Sc4R0TtC3kasCXdYiismmZj2eispyhuTf/VvVjmUqvz18bh2arIwA9iiAeyMOru5q+/
RCS8mMXGMPnQfddA4MQytM+vRHJmXr30SsIA7eHLTtJyWLqxS76jk6KiQkoTn1rNgRMn8LLIo9fr
GFDPGFQPm20cz2Zc8eZJ8DcO96A5SIVnMIJHUfNGgsds6Kk1OWcoqsruPbTviJIfbk1otIUS1YMt
BQhOqxxLNU6qSLoeJhhaRENlW7TA472kc2Qo204ZaJFz33GO6IpweIMSo+Wgc05s1AZgmjaahuCE
I1vSm8AGO7bFvC5flxCm3pQMTkdoB31M2xrhAK6gxsz4m3o4ggiNZve+BM/qxvyFkwDe+ZMjrkzR
RicJG6mI/de6OCbSnMvZd/djPkNo7SeyBz8EiGa7jG1iZgAulhrim0Ytl+E1AlzHmG1TLrp2OZNC
nEqYIZyriB9dBWkKr/hiT2iKvlZ03pvBl28gOFrj7vT4I5yY4Z53ppeMPCaU287wYt0HH0aVvzjP
CIG5WzdWmWpkdxofE15pzlqLCjJ9CBlbyUJ7QBsP5eyaJUPJYmk3jw04nkt8Xhw1PkQN6k4lnlx1
71ljsikKXYwvjW8DhqsIs90qxqN3mQa+wX1hKOBM+JpRZn/2eW0N51JI2DEW9XmWUBLPgpou/hTC
7G8QwkXYrQQM2UFr7AH1cafPIIL3kI2otE8TApDV6fQKUyYxITuJuzwthcssyRhfip19o3Arp4E7
U83UW+l/fd5l6f18Ec51Ji9T4F7fypEub35UlINZp1TW9BqTPg0MXQw4MaRxjUEjQn+ICJd6593Q
LHXLNcbKB/wsQ6rExIWM0lsxf0WgDwV6fM3X9/dTsTf430RkP2FMqaddjhXBGVdKqWKHelV0svf3
Jb2wkGC7WknOd52nk1uEYE9/T5LLsaYWDxN+wForx2EfvoHqBaYURbbv490VRjeXdmBWbrGuoMOs
Lnwc0YYZF/C5nUOClc41QW0tZ0u2Ri4i2ctVHUMeM7z1JbmfrcaW7dJKQUc+b9D3KZ8skxNHoYwE
8pIWi9Qo+q28ZvkyDHSZjXYw+GXei9vVitnwfhQRVzWOB8izudJ7Fa/6E6opUdAkGQM/iicqJ0mK
1uW/8eQ0OY5R2VD16Zed6P2HvyYBzDHHiCayrajnkTnjG9YthlTpdaDtra8zZV940CK8UzXpv6xQ
UwOm0luKTIX3bNhCm/jew2eHiNHTrsskjHrwdKInaHUC3hnZUoiUtIb4QT4Pk6OPQCXZjUeFKwQj
t8Kq2arIAihxtlIFFPNv5XqDGi9HNtrlrPezzd7/RcQCmLj0i+oCuRveQJffnmVoa+HEOMMEjOC3
yfUToKxAwK2/Mjh2PPxsZS4IBA+zaL/KUIunKM6e2lHwIsybasLkxYwF46KdTEoW9lot5/PF0bV9
eTksjAxJEud6ZC14mjfkExztYFRp3CHTQE+RDvldEFtSemw3OQ+BfEtN5k3v19TJv/zGr4X4XT7g
bXRS7Dz6OO9grGwiN2mKvT4wiy/PdbwNMQXMmfKj00MbdRbX43cHh0P5h+CfJbi7jwJhLkG+sh4/
VxmUYb9tOjZhDpFU3oNHnXtqv+HaIqoyTsiR2XF3igGbkIm8C1aHpY613/j/Hj6X1oxKy7oQHUXV
XXS8otgyR6e39CRXwDs96aVYx9WMNFZ+pW1jp2zLWXbJmCCPO1qlBxLrJHL/OJpo4rxwj6mgIJUd
mK+MFfc2V8hPKWpbyspsVd8EoyoPK6byr93BcXxLSrxb+iiBoCstkai2w2VKZuaAhHBHA3+eSHlY
fHfnZ89k5IW9v5NzGmuLeSJIxs680q607tgaIfZrbofbZE0xluq3MFHcGlvuXPEn4LQOFUZa7XSw
8y/PTVk1i4FXMbiiMmTdOFxOiaKquu54ZeUCmq+MQiaxZvYY01HW8/54SZuNI/nk0dk7GeN1Oo+z
etzAfIkwRPnuwrUGW1Hj3j1P2yGl2lrDvQL0BCD22uM8bC7tYYa9C6Y+3jfMm6mUBMKidUqgqSQV
C5pXJjo24PAJmjkfR7MzRKxLpYmrUy/GrR8+C9TNnlospGvk8acltIOGtCfdtAvWAL5Cc/Ph2mL4
956CUClaQKneQ362iTTtTVBELq5cPdz+h+ZQaRsdxqXYO4ubETLFJEh+/0sMlbsiUyw6c5xx1R2w
fC5nVofFTACsHB9LU5aeEK9ZGOqE+hfvN2+unq2dBU9tsfNcVr7cAxUpR5RSkyKjr+5vvH90bEHu
l1BiUB8LAGsSfMPDIpr8DY1M+Qrfi5IKrYJ1qlIjOChsyAQzuTY+MhdMbWICb66WdTQZdCUrgt50
iQKts5S/5GFSUmUi5RpVWQ9kBed9IOkgnrK1RZw4J0U9LgJ3Pn0EamK4BMbHu4gd1BwmrUF+vt/K
j64Kym7dHlBZapaWFZdVPuMGgN9S0dqQPp5wFnfRhvw6ii2pbvuBDM1sL1fUtbie5Xu8X9ELhLjk
ENmhC4JLNmXuTPuEEA0dLSkGp4mv3Vc5P0vClPq20gDmtEnJ3RjE4o5vn2koEhQ08JYh5wD5ImQJ
e4eHOdFfj7zKVFVFAXCN28AjdiFZbxSUmTyrl3Xz4P4PaF3VbtN2i4pk6Xhmn8O5tUm08OlTBdg3
o7L0NkF/EmPfzn4jDJPhGzk4MslPpEKhdPThGRltdWwLfs6acUbNaap1TfGpfV5sLyk912WFWEQt
e/NBkPP1ZTEGK/Jf7rqpJxV1pdLDnc+WVOrIUgLeZL+lPW/qPU3bZB/NWYr0PI61tYNUrrgXNkal
t0IoCUhGLHwVXxKDrjjqXa5pcPOwfkawNzYDyPazRQrnZ6o9F66hDFbQvGpoa66HizGaNJouul8M
bvoIxq8gkbfk+xndTdh7YnYa1x9feI5QoMGg+jUb0wajeNazlgGe4rehwhTwgwVB1AMm9WOaDd5s
pw4FSUTSQxvtq2dvuaGJqzz1+4OmuaZ0viNNoDWLKZvivHit/SIVB+wG8Lc/uYLZwfdnEqDMqolQ
9jh9kH116B2hALyAiq4IniQEeMjC2YYPIfVJWlYmAoOwCTQ1/ho4NkwQ81ZAmG//VVpsSEcc85/p
Mv3jPKw5rvc0svwvbnVOiZUS2becDd4rsK5XXDP5cIzNRC+YZ4kCdLf9YtVp4CcojPyCFMQPGUoF
BBWO8d5egelt4rgZbVHw+Mqqx3gr9tKtYP/jc2JTJAuUbRHyAZV3RWitvcVUHIsUqXwmblkZfe6X
YwMLzmq8T3xOi4ROKkGIDlLE3zUD83N9+jXCsHTx2uV+cv5jaNofHUUxQZFvlX9terjslO2qEQ7K
JXQQbaj+BCF/km+V7jOOJ/DRpwaPJGFQZw/vn9KMQ1WLd926D3pjnAbrfMHwQAMdMLyDrC0q7Pqd
UIYdjXxU0zuQhgjtc2JdhTEV+eUk+zi1fh0IkvN0f5hT95Fw0Ir9Il11Oa1TLEoBxjZntJiDYXIi
39hd0DFH/JzO6PjOhK8y5MGuscobAOIJASG1EyjwgPTqhNhaTc2TCwnqllnIhmC8jPxF3djunzi+
4Z8y+vQlTDWCflYf4jF1fMx2cYyiOVDAo4gmSDmTAMHqxSOj7bJ1GhqP1CBKnxZPikA2z/lu403i
G8isnqAg2bvrPlGMk+ACRpMl6T4QcZyFRR4LdnCmprlEVQX5Vh7tGXoWak2rhxjzNgm9Py54mFOx
TLiu41j1nPJES5M6Jyw2pPIuCiD+Hsxp5/gPV2pyxTk6Y2iYNsKqV5mM3cUb6V7rkURMPPtUfc5d
3edV0ykOWYA6QfKztT6aD/N8xy9dCvMVZmPuGq5KuON1ggGyT35EOtwrAT+uA90vdeGoNtetESBc
2kFCt6UmzplSuBvsOUbsOG9M04B0DhBFmWuSNunNbHOLQArhHAs5QL6GC0/g/RexEwqblJ28OnHD
tq/schoxharXE1g52bvOlR/679eOFT1CFC5ts0HH5uq8bokJNxSrV4Ro689G4cJU67e2q5UeDuZo
7+qX7UDYylJL6wI3GZJOuOhTOrWoCHTrQ7BKaZWV4H0jUpMUW9JQdgtve1/2wsaIG6IdeozNhD8h
FNmRgZoDp5WMegaEgfex4zfS5ksjg9iG5cj6+XM8XL2aZYaSSlS5awe1ZuVls4t2rGhNBGm8f6sv
t0NRPn2QndIF9R9pPMzoBI+GSrcdj/4yLS2S+liQlECJs1rXb4IRj43HGz9RYu1ZMqEKIQw6BlkX
snXfCWMMzZJqr+BIPmShXMUeAgeumYTe7D9SMGU0XynyvWB/uHWZJxtp2W04VIFVgV2FEuKIrdpv
fEnjdJIr0q4R59qudL0oIP+fOMjnp1i7sQjmGuYAmEJEvKwOO7KWRrOVw1pnTLEUsR1RWsiryj6a
6ZWGQaIsmKzyhORYybuZOyn2Mj1rLrMXs5OweY1SdK0w+HDOmQBdWE2oEUzAHqpcPpw0tzh+tQ4y
3st5J9OiAhshAi2KXEads6TfF4j6Lz3dmeP/MvPVWYSvc6EaNXFoLZmeHuNkAJhJgFbGSKjPS8zR
So4nLzVnbDtLZAaiEFMaQKz+/9/dmDqbzufZpfFRNb4/TJYIH3FO0dnqHyob8lBoHFOFoCnOY/EZ
lXmmGGUCnbkn/R9/J7m8lOawnJM36uq7mYMF770E2pgF7DgDbUwZonIlhUuBAoezMjXUzqIBOMyl
xC0TdOJmIyRWDrS+EfrV/vYwn/Ap/kDh+dUS19fT81o8hXAK3LpyKpIoaA6Dkex3PnsCVQEN2Sbt
Oa3PzIuvhPoVbjiZCMXlYmXwkHTcuDNzry4zN6HucD2KRUeStAYhFFHDWLfj9tINRfmCRvJ1oxD/
smKcxWYKErwFSc1vruMu49BLq9PTmyO7SBFK0XexsMv+zBmVujYmxJoJwricxUK2J7Qk53h0OXRs
lx/V5kg0um9VCLONjrDeZBQCMQbyz7XOHVQF5TUIhWQAV89NTwarqDBKLFUQSngj6ZP9Vvi6+vrc
mYeMjT31uLheWklH6pEgXiHIdqq0ezJ9DilOK5pWnBRZ4i1Natz+Dk7uYhOAuss1wZaLlQh5obsR
+kfucNcIdJdgVkWvaWkl7bDwNrU6nyQpoN3Wf/z2LjqClastC8cZK+5Oh5gszheMbQMjc7V1Tyez
SnaqXt/lmLm0slwL4+WAiSQyn6GAxMXRO70OS1LImlDJplvqz38Ywh2uFYs81ZDrDK+5xTkdR7Yk
9H85nRHN2MfIGkH/y+scio06MkgqzbZCpr76BH537kYRtCbyHKbWfogGx2wNjniVyYidFmI5S6kp
n2ZCk8149vXpevNTMbi0R/hkoIls9oSA9cHLrW1zr3iiIboEZe71BWCrGZsEF9iSc+0Tm5iymQAt
JADLFcYd7YLiCCqbHQM0xVq/vTid1Ibmm9gEdipxcLffchvxsTM44F036qPzbJsb0VnphLlP2tpE
IQYgea5CKi/Uwfge/UIR8DKoEVUzYJ6Ma3LNwKUAtHxhQMgZsqcHeI7otT/8P7Q2A/au3YJMMpCq
ZyMT0CZqzirfI3DVxB3h7/5qhwtasW3jcPFwlVrhRkK2W9EIZ5Div7BE0VlWsM4nVhDJ6qj/fQXL
+XTNKjyQxOH266KHwtVaZaFv/wsMtT1FQI1oPkn15HaSWMiWz5nuMUEwpATB9sptJozqdjBFsWoO
hetUvY7d2qxXGRE0X7TqgamnoJzi7dgIEhlSnX1V1FZXptv8xwKcqQGeXDE84ShP3St4+NMbEXgc
Q5T39TDARqoV4D/e4z73xyZJikOFklwfUVIG+N9g2Hug+p7S+6dNkk+RG6cVEZUCc2Lch9tl7zV7
Iq9Bp+ElpDUhTepOc9RY9hiD67/57yMM8Y23lXBXhH/59799+LFgakxhRWIDQVtWg6DtSr+Av4p7
7bVg2sxZGDfh/wlQXzLgh3/mVxXWkycNOiR93P0yeb9u3HKUjvZxRR+Gl9WcgQqliQWEkC67V9Ps
Hc7XhO9rIQ3DqwpWlBSk/JWOykByXzIiY8XUhKt10RxKbN/K09Tx0WTNA2aVsuHFHxygEHy4ipPi
tor2F0lbnOzA3M6lR8NdkT8HRYQjhcR/DpUvmORpmoNUOVvLSW+TBY6kojk0zjbJE4Ol38UlpYJu
SuHJnEnbGczlHEtqq3EjL+96THjGgJnGmQzdURZnLVFnXRil/x0wfHdfQojucFZb2IJRvTllpjA7
vtPUlSOrxZPwgLc9b98TDAgoplRawtJsgs3FbBOwc1GaKPCsuLxTx2StqzuOMPLxYAxbEWmJ2pNj
GnHpan5v7FzPh9m+eBDVlrdUqcKbAmRgPZjGkKCY4T/47GbEh6978EBs/xSwr/PZV/GJF3FYUz+I
dytOFWzI3qCh0x9336sVN86+fHUMu/ytO77e1+O0dkLbAff1qVO1WnFzeeU7Rd46M7uneHrS6ybb
eqNX9NMkITqjMCdRoVEfo7OfQCZIUOXzt0Sz0oRiq176Gp5j4RqmTE39SQAA6AMqld9J0+vS0Iri
dwTVeunhNe5ICqb0PyHAN4FXRfr3Bgnkz+npkKrcY2ZsYu5ykJMWhjoA/sZCMl1sEYViJZ1GFM0j
swxcajvURwb5+/BedgZLstQD0r1wsaSKtFTepBg3jUoaGZjiGDRQYlDann9reYaOT9RNZN5XXsjl
BB44nuksN918XB/N0iORMIP2ffdvbzbnmCodtF7onNZvp5mRKwewnKkMfmxbqwLEtiANa4pRw2c8
lrENuaXen9Skz9Cy+rmsS7yMcjaa/IKs2DbsEdGtmSl3vxyFdrfmc5ovV4YLoCusmVND4JQj2BtR
vgWRr2ZuyXSkfdgjTX6IXnTeywJ5s8g5hcbb35UZw7OcpgqAaPHIbdfb4YVrqSmhly4N51bttJRI
tnuChG8V2cVa87W6z8POZvZryVU9xow4K46c1FoetYQQcjJj4nyN2j7eIgBdoXpdkZvpdh8mw/3W
ca7jvrreekmXHzoC6g31qeHq1aM3dyUA1RPaFPe1oTVhB6C8Ah1CG1AR4D88vyIdLsc06QmHHh/5
j+bzlr5APyX+SxGlqnE7+yLT+BRLDB7g1RwT2cbQr2WPWhALfKmIXciXBITCDIhkB3/bLzR66kvV
F63iEkRz9Z4rKlQu0qRg33TxnUp9WPNtsvFWztllW2fpP+5JFcAdd3DjmvcTUKLMzXnwJvY8hhzJ
7BTFBKJtfHGTQMTqfR2yf9IOjOlueNj26PCE8GYUfZj2L4xwSeo76PmHryezpJqPNC+4Dj+xwn27
o/rUPtleqytB5DCx+sz0Bb5mCvCJWKRrQXpypE3c3euVGG+WrHSDacnfdntBT0RZ7Sk177UIYRqY
AkH8cSbSW63EGoPJMI9h9DEGJCdvblhKBixfVcdln/a15cLSig+eYqQjM0CgrrN+5TSl9zS6P1Nj
od+z9clqy6BL6na2S5qaOxulV1YzDcZ2wxoyV6tl4MriqTfJBmtWCVDYz2GyCLJOGzmV0pKih7Sm
tTTzIjrB6MuD3Y9XhKuCV+johjUE7gxp9T5uZee4Ns7F3IX8O0sxyICs4c0AT+kFCypy3AkhwPY+
7YG4mWaPbFt+nIDdJqiIpNQzNfYiP4oLtHT1QvP/DQRlat93/jgvcfL8JScgzWiQGEeifAeP4LUw
oD47H6S6Y5cgjYynpHYJ1LkG76DNwzxcDGiR/p7Mrhkopd+g9D+dV/IQ8s3HBKiIjZ8bjoE0FlaA
ttBn0OeffrlTndlf/Gy6Ds6R2z60OVSAtQGUdahlfuYArI6okbyq85tbVaqjm8U97Gneuk+ZhA56
jZH93rSQ8iVh3Fur0tSOyUC+OvjDjPEBwKwU1DobjEH8MWkb/1hG6hiwZB/AGPqXCQAZWzakCOoO
dgBKGDFMPhYmONy4Eu9NMOs6UGhOWnEZE27uthrn6AXxdzGJv+orXsLYPId2p8TMh8gABSy8BI9M
fxu23S+msf2okYjCdbbQK7oGwLVUHZY9B9Y2Vov9lfGGIw5hllVCwluJC6hiJyc1z+j5DrPVWoh7
FRhqubEBDlTymgyql+WJkPh0gt2YKBpRSW6pXf7EX3JVPVxBK1q0c9gihEnO7wQ2qov0yHm81Qw4
FK5mx4Gbf/nVwa5DSxt8Hhv16ZWeFRlAWznNjKWBXHVgGQTSHvfA3s9a2YducbZQ2LexnLTiLm6G
Afxju3HPhr47Wzr6/zTJ5Ne9xS1VCWbwCozwSXxL6yuX/dA2GbUYtYlBRZRyTVUuN9C2eh2y9rm8
R2TxuB8h6Bhxz8H4YkkesKA1V/FLi8hIsmR07rCF/XsPZepQcwgGp9QpNSTphP52KTUSlaUdnK/M
/RDzxCzseQMvg1rNBqTFtKtEBgooMMTzjX+fk9EKLeOfWUXyOHuKivDBSth6av6CkxzAxt6k3mx+
Ly1FOs3Ey8k2ggjs5HSfiO66IixgNa15XP64q9qnZMd+zuJ7fDzouFmxZpBiLGwxhMIdFmtzpOr9
LzerhzMdAZlDLqQwihz6Q1hbl9yP5nUvG2A2wRZhg2yLpOwcvMW+9+N9iFOUNHURFc52aaVX86FE
8jyyPKdEbf0mcwpDulANo2jGt+XL0yTQ6AnWEg5/yL72ZfV+7Tf2TMQQkU6EKUjhceW6RhaE51Mu
HgNYcFt2oo/MPc+gPLWMCrzEO6GoBU70iy9d/h4b/faK5/Gm+2iWqsliZdqaJGUQ5QOSOEvHlm8J
/BgXe+vLoebtkbLDgVwQYBfT4qglg0lpH8AOxEHh/Un/49o7bl7GPeqhRzfHWLe2HULubJRZjNjr
xHadaiT6Za2wdAqbWLpO+CE4+w2voKT8jRQ62bXAyfy9VIt7ulsGsRKqI9l68/sA2NAB+pyxeF+m
bcjVs8YMF1LS7AqXT1LgrK3EEHKsNdJksAM0iHgD8PjrMU01r7R1kMVQ/FLD57xJ5TYTpPqbs8gQ
1bKyDZVKCNL0hVNlXPHSkrkn33e9TODFSriygf/ijpKpS7Rv92ZaND0tHpJFfp3QnCLBYw4iivqC
lVWF0zJmVhi9vtEsQwANvpS0sknAVYe3a5kxd0e48wsk7Vv9LOcmZ1MmAuaw3Tih2F6CEdiMLZ2h
X8kxfHu02DFjiBhgHS74pe64JEgtaI0kzhr1aJS/vfwcpV4JdnxjQ6A0MEHDDr6wCMuOkgTzDITQ
5ekoD2VTpmnSwNzsGwQGVmJpvXBNGJ9uBly6FB9YpFbeH2+mDnLfXZsGm6JGwUo/m3+y4h6b52cS
eHd55dxVZ0JwfIG0qlNvO8arZ1G4qFUmNpMP1uRdoJq7R6REWYqy+vZ3H/RUT64ylO15umL2jw5e
RKMbTpdcgxT+wM3xUi9PW/EmfkYRZ/pItm7iXX3RrRapBycmYyIBVM57jT9h+IqrcYt+mQDzTJIt
3BA03pf0H4ArwqJKqNurvO/ko2Pcrz8WkWirdFLNGwPlfp4kqddjxf2kfRQDvuX0Z+UZOrzrEP0b
pmQtnhBGi3OyFFO1YtL3sBKJVCyWtZVXDwNmVK3c6xn0kIGogOWjtebcQaghKI800mnBHYaD+Cna
ygjB/auaBdd+HsX9qKubpD2obWB9MdYApnlEQNPTT6wcg5JxOLTizI3ph8+LdRvwVxYiRmiCGKAQ
9DRhnSEuG0+A4CYJerv5aFUvC9tmWjpjuChuKlQAPyoJWKkjmIDQUKYd25IiKR2bLj9S6HXkgry2
dzmHLBFiyiuD+rUAvgID/0lSSfDhnZpJh0OVruEQnpuU5jTPqiltBI9ZXe4AAkLrVW5NS7viUUV/
dCr1HUkfypjhYt/91Zg1zzByx2RpF/i02VrndXS8Ws6MHcMGills0MAB0hKN83V9raJ5cKbAcCG0
Tt5s7IabPMFNdwX/u7y0y6mf3V0XR8QZyf/80a/5A7SqlaqQ3/gqFjIzINvuEeniGUHZSl7BFPk6
Cz/gJ9knDppyING1yH5HHDiKyNABZ7QA+3xLfm6FY3LseDLkNxlbcDPZB/QGGwJ1tKv2A5dlKX1f
SCUW365ozKQKdA2CUsXNOZTg6VpEIBmYk5il/rEPv0+pUkMVZCyA7bRJGG5mLHmdXBIQMfuCKhcR
G+z2bN2iedd3MXNR55mrYGgTSJPYJ/p6dN4pmhoI2NtKVSv19XmLiITimaI3IDTyMMk4npzrx6ws
XIbOsWz/hyBq8BJwzZZ9RnWJJNxJlSaIdtYyaJ6D2Ww0Be8eB9zfJ3v38L3sZuti8Ntt52HcXlck
I3oSD+LMfW8YVBFBL3y2/uA7JbeyCf93Qu4vVqFpGkYvBRK0x0Xsaj+/SS72DROpXRXoH/cCJhn5
TjZmK9dlaRu9O1eFz8VVSxJNsKHoylj+zmyF9yQ4AItqq35RckZ4gSATbN3FhMMRYt6yk9nSrqQ0
ztKukPX5H77cye8glMoWfqMspFeEGg328F+QamH9lLSXDe+1PbB/FH6EIW46faRK1Zc30bBjQJOa
GsrNt8HBOZcMGL2IRMYoyfu0jUoSxavNq6FD3VgpYhK/PyGs4e1gITi5AUUUK4sEaoCjI1QPvCL+
OJYZ6Le0oAxJ3erDu3VRjeFh7m9mcvu/MBEL0S9uv+Z1/7ln6uxLpF8GVM/GsYK6XEYsNDtl/Soq
6HOqgArRhQ7U5woSYrsOUzSQeqmn+1okNXhuzP70Prk81oMoarfTg3+pArl2+ge+39QF4ppxs4bI
6EEuuMM+uy+vVDVFL+LAoX4LL5iXCKzHj0FDhxKLM7SYSYfmRMyX3BhvL6wSoTwmJaBdJckUx96R
QErrcFKHPsECWrszPGGVU4qypzNo1kPYoOp8dn+4Tt0nRiysxvkJCQoqgfDnUHHngIVjNN1mJGIW
4tJ6kLGP6AuhOYsfQ9ui0zx5tuAATAVXzdT//BEsx4Y/+INxEeQV9UL7qzysJs+qAncLEUvDay3Z
XGUMn7yUOhQP3DmuQOWVkaFztymnr91f0KOTtrx5QvnxdTnTWUyykMSrXv6J/k5qdKvu9VMJCv4a
RQb7EF2JVdtnylIFj3y5Z5lNQjq3D+9fSIvqYgDHbU3zcWfr7G4+APPPckbhctOpc1QFs9Is18VL
J/Y3sgNtmsBS85RezadBiUCei4CzDlYgPJZ9ICM48+jg6TUr1MReZiBd55iErtMS39rl4oxmTont
RFWDQNPZoQJgZt6jbsoxgwo3CZ7Hvg0ac8hSUr/bpcqHjft/L88ucgehXWzwV5Y8uFO7dwmKQTMU
wtGyjLsfbyjv7DDCTuv6zm/Zxq9xbdUfJpKTzaSfvyNWQg4UW0NC52+U0Rr6CC7iwvWsEPU/DVGV
9QC2Afm9JW9rxOBXn7D/9vxulw9KgyAQAkBco78jpRAZTlJfNvhluXs5Kk3BUjV+EEj9/otag2tI
5WgnOFYVbFeCdKfFAGi0qhmirmZeao2UN7wX5DZs+/bg15x3fwYiOjcp6pNE3u5gQBeaySgFdaZ6
/FrM9bpfmrTnsAg68aG1lulH17S7neAx/+59KdW/iX/D/VobhsKCVteBY8LGJiXekLa82QitMXpd
01c7vgw5SaC1lNdVA7/0SiucRhbrx8122G5mkOSa38u8ds4LtXXBAVIjLxACTfmK9bdmF78Zpx0d
OZ/E0/P4yXsqsCAej9F9NlDnbvJrGGzd3zzAymlwWeLNINnRXtBbRwjnLaIxSdfmZbKCcCVf2pWr
QyCFVI04uyZPNwLX9aplX1OMGmwrIs8QlonSzivUHrcZzA5UCMXtI/mhL5h/L4iGjyY9IAYPDGFF
a/v4Uw4Gz2RWIrbqA4Gj31XhPSPHg1+7m1R+SA/RBtzLAa0Tez/2d3hFvkWZ+fn5Qo5oZwxMKV7S
P5R7QqjT03AoHwQ9CVxmDKFON/Er8dSuHTaC1IbxELSRrzaK5GP34j+q1hl7aXFRJhGSpGDmddEE
AcgfKXwpCkXerw3HEafqVBOZjqDQsXSP2aD7swhexuWGJyLhw+2ufDyohqahDQ9b3f+ORVFaONfc
rwfphMyuxXhiOPh5PTTlBmwQowO8a74Jpa6eGNJwV2DZFO/gLJG5PyNnEoOWyAk1A5eE4Ti42L6Q
b+2uQJCxdEi6CqG4tU6K3+y9e6+RpggCD9JdNFxx5anorVgfTjDHALzdQwSFsZS++fcH4Rb6dz6i
h19ilZecMiTzyEH1FjmHX3OMhwrSv4VdlcKCCplMgNDuqc17/5p0/vFCNxJybi+PxxyxffFwtITw
j7cVjGKGjU07enIxPLzvefPtZf5apAaWJCiWjT3410uTRuCnqf/83lOajybYquVC9+KVI4+4Bu8K
BCHGnM8ctRaoThGeyWGebcYtcXUbJvROh25P6KoYbAUU3e8PPkaKJG6Xn7xXducFXdWVrCE+WjX8
ZIccuCSkO4k2kxNuz/9/hgCwQliiASiuDdyuctRMR0qBTwvtDjFr5i7fpZ6ekxvuW5r5BdZRfmM7
7pFddiOSC6ovW18HgPPk66JgOjvvSVJbcoZiCrUKtA+YtbmgoNt+OWosQ7u6Cf8mm5ai5sdej/IA
rHiUkzJ4+ND9nLqzYgC0swy44Dl2ZOhRMXIxmacbZOAGFE4EpNq5hozn+6wW8u8uANkYFOcgXdxE
tecY5/Dg6AZabkTIOiGIAVRZP9kLWqdJNprpTW4FwoEXVDjBDTOcJuwa1dm4rAHOq2RoYGENRMbp
ddV6bLjLuJRPvbfbdOb69l7dJ9etCMaET0y39Fm6lSKeZKpYJhfg4vhMJiiwbcESMOJpX/fKUOqz
/JMx9IJXKbrMzQNRpjXD0hPaHhGUh2bETXHuprU5nVOkadMoQbccjc28nUEhNsFNGiqwPve8GJb9
Esu0GagCEfI7iz0ex2Hl1UBZ3BaFfatxkzOrdX2enyDyI9EuCh+2VTqa+2SnAhPOMDYH1JqK/Sen
1dEyl+FKgvA/UCHOQIjsLH+cDeNQZ7DGF38YT/rvYvmcMF12jTL1ht/9bWDfNNBwHGUMjHyvqFCd
MvZyw57e17Iu6OjgfcqnC0Yzl870giK1kxxGwcpxi8kwsztQSEHuY+E3MYGX+xqPOYaQygMxiVD5
RziIy5ogD+t8wN+qFNdB/iKArqvaAYRpLxoIgD7ZnXfQG9gqZDBkfj08VammF+muEUXAdAhcRoRE
gP+inz3kFrozl/2gwO6TiNAqz4ypiWjhxYDNcNu4VpmK4PN//gobX9oQCiTVM3fS7q/TW7/rRtRZ
DlZjv0wiS4byHv0EtEYV2+9zwu9QtpXmGYRuQkeCuhFCSfIxT/hR2PMMuBNNi2GKqJe3sIqsVEC+
Q80t84mCa8Y/cK8wtud87x7sE3KnsbKiqdrpn3E5COpoPcAap7Mms2CgiyUc5ewxukA0q7QiIoTh
ungxa5544eV799WBuIJt26kwP8A7TeqR97L5LcObhgUcE397ny2hgYgmte7D+2JHKEqpoDwKUIxu
6DGqeP2uGm8nQAnnw3WWQUxMjQIRaSHcDH4VtZQ3J/G0MTynxb37o1GxfCgOuM0Ca7CVhqUyrhRI
Z67t9CUFGpsRx2GgtMHReBGF3qdvAAZMDsEXzGPdf5ae6BMCdcK8s2U1F7qREyzVi41SXH+7k1kT
bShIIUvghOuAFcmv7pKr70j2bTqTI0fY1ZZN8lLssZXPyMb/0e5BXtt78s0LdRlqjD7EiRZTJIKg
8mpyJl2vXXraJMK4zjAcpxpy8VvCBTPY9LiDq5uI3eLRnXHY7w4HTb/5wdHinrcpkapSt0geujNj
/waCnw8LldhdAkVLxaApP/OY20Y5iZDiwixf2vJ0+RLONl27CyrSNDyg9S1Iogdy1O2xGQeAMT49
rmesaEI8PKw43UIGzKUAPDEZ1T5apNUDAxEROnCMytB0UMRhTJGOlGqDO/rUr6Jgbvb/k7B2YpqJ
JCD29DXtA69A2rfqVu8sBDf2oUWA+tGgmqkbbXIrAt0+WqQtc9iLYXrtWDQY2rwV00fyby0zw7L7
fLFLV3hVyEGGW/STXHwv5W6BAEXbLtf+5u3LxKvBf5GMh9lhaHg9grT3fiYXLbBJ0QakmXhIeoD5
zT+RTSwGJYZNxY2jrM/7oCZithgUXFlLyPZ6tvSVz78V9mnKtNw1iUMg/at5djQhZRZ7G6Sh8lJ1
2/A6LC9wRmM20URjlbWsn1Z/j5KcS66YGwpbr3ISYqZv6JHhKxXcpDQ267Ip6X2zYQNZV4drm2F9
U2XCJ3v36rYlQ9VU13sgBML1Dt13UUcVIASw7oWByQPSWAVZEaB4Rs04WXBkHl29XaGHTQuiuIl0
Oxy2lUJ/7ZsfLsBLPeiKaS2uR5DkC6IhjqwjqlHL3i4Oq4cGQ886I6EcsyJiVrwZxy0+/kVGAs4M
0Mna77Dk53DpKGpLGnb4R48kntOQJQXtg+2lUHY+WsOIR7WV81siugEkuDBAao90QKjGgrekh/Rx
cGDqDFfTQRrcahdAnpTjeVFxnxgokvICChNOJjGh/5j9pg5wklUzwq4w5x8CRXOI6RMqP8envVCd
tqM2Z0NE5oKAKBXm/7Cn+v2scoyaPybweuVcyCHBeijtuN4Pknb5Ut3v13SB6kFKr4g1uGTLil45
VCDeYrMQ9RWwkBz63i8bESZAFzEW8cUzbltukUo2poD6QBopVESag51szk5N98VSUtcKwkNQ8d8j
zzj/df+v92q9moEQ3Qf1q2lpMoslXoCNLMK/mw6BMfKvpDC3kMsZE1TDUEld/DlL0iMxaY76zALv
fepufXZ135nC7h01iGeKhKsgtBDF7RQ7Gq2GjMve6c449pK0FNilG8rTGMUqrFQIEgDM62AqvG8k
+1tvK32+XnbqFj3b1svsPcEhm/d+SbkIToHgQNE7P0D7yKbK0kEUNpUGuQSlLETiHFp1bKUfhp9v
1KDawD/AByhxMX/SWpn5qBFcaGAPNmXeO21FZv6n2DRGs+7G/fIO3+EKnmUuq+l++rPwJoiy5UUK
1SXV3JpdplwYWhLyqF2NWbKnWiTzoV05v9GnWEwZc7K/vsDUGCK3Ciy8W0e7bpJ0nJn0Oi5Vmebc
UhyVAfbEbiEh58OELanjFn1JOQ/3NR1O+qkEfdy9Bxw+wP+dRcgiY0RO2kttls2rWI0CnwuYeaMV
z28hxYsL0IqNErLkJweWlax+Osm/wdySjzeE0mLiVzglAoakF1aKHFpzXwSBshHuSjIc+kOT+KN+
j6je3nbj/stV/hvXiKular8YOkO26asGOQsdtDVlJGnUa9IBzRf5rGPdSXTdiQ8ir6AWGMFCtW95
J3uSBarsmraiIfDdOI/xBFVsE4ABZhTS6YWfdIe1tdp5F5M9BvKLEd5VkbJ95xCdhEROXVkbpJLW
5wcVbl1/NH6+uOsieVZwx+zeMyVmmWI2lAg3H2wQWSP5oJvfKSkVoRF0gy+guOMM1zMmua4xIKmg
6ADZZSceZRlIVu64Q9qjp/Ab3UWl3Q9zE9guemHMLc6z1bcFn7pEmV26hi1t9DWpSDhXzWQitlYt
VqdEDYFlTyvM0/t1E5RZtrDHFox+R6iFDwtAFj0nG7idA3aWvN3Fij66S/pKyJ/lIv96ziVYPtVK
b2N9iJ/Z01rxPUhWSChLMZcg5D+/DSf9hN12967CFKGuME1wKa1fJDxpd2JLdjV3jRfjkKQNnPGX
FzfMMobv66BcROq3bpILTBcgJenly31Jgkf094LGH36soOOXRb2KHBjZNxU4sk+x7QF/RadhJEmw
X7iK/B+G3H54yqasQbTIjtR43Kf3SoTJrTpwu0Yr0rH5PQY7WH/BDz6njN38xcIDECTnhrDfOyJY
f8HATxzy92cKx2ndLErrx61xQ7TsnA097fuS1zS4XYYMMPj6tNjsVnbypiPpbPGHDoVj5lxgGn3S
9NN3RVpxThR8CNalLDvIOMG31t6N4W7XcTqXPqoVwK+96HXBg2JBGw3NhjYXQXVnbZOEgRfLqATQ
Tk3D8O2UAAuWiUul2qdD6nYqSU1q4rs47dVuIUYo3w/IX7VNQaFpC5mWbJdLHkn201M4lCtJkkBH
3LlD5KJgkhWUuAscDbDnAsq6PvLTnN2RmFYqBxPVnwnvEf2B66YcXOp9EUsN21eDR7nIulKoLuAb
cneZ27zNuCGHgSL8j737CrP3XYlHeH3Bd2gLdfS/IcxUnyO5ddGKp2bAtX/ockhl/yLkcXRXeIGA
9rJmgkr3XwMmMoljKfvuTIWRJAdKsqvFp6cJ/ULXVQXMyXb/gz/WCviXxDbBSmz3zdYG6UVP53QH
IoWnVMvrh8eRLWQRC5U0lNadHtaQ+CxKWeHAY8+c1TzzpLGr9PBlzDgpELDFHgLlrZ+WPXoZswil
/enbDvDsmkJtMjA+WvNeSijGwMGcdVYoh3aJUcAd58igz43HBKqKMVFrLzXvKMAlWoDoH2RP3Qfx
bR4CCI5EYzkgq6hrYaRNO87IyPorTSmPaDg8QkSlH3tEAsHanhsMvDsaK+xZr1pIvCJRql4yS/Bl
E/4YCLsgod+TKbeYJhy/dIMyfGDQP0hh/5sxaMup5AMfIOUySR1QG63ophYrVh3yzT9njn50f7N8
rx2beZNNgP2dMgCZznEE7Kn5BffsOpN3F4LLDFlPf7Uyn2CBwDb/33h7zHSh3mGlBq3+dpddU68P
YeLF6Esl9InH13lN/mct9lgOfgK8tYfNF8ewUGFa3k7u+Te0BII6j2nrYSiV+AZKORCG1q9+wJDY
JgtHnKFsEEj9ly3v4QElvo0WxnLY5mTQKtDEso28A3hQka+IduqRC6DXYaKkO9dzwZ30rGN3ub9S
u8IY7Rh3FsRlA/Ve4LDnvk3zh2aWYRdliNkjNPFVNpqHBb17K4E7KZhUj+mB6UjYfu3IvZ+zVk4k
wT9uKWiqo6YPGQkozw4h6Vn5lD552RDdBdbwQ36Uqqzb/bPxw8QtNoeVsFN75yn4Q99FYO3q1MiE
fQNlPZMiX2umiET5RhQlHgbWMZoHPzzltAOFug5zX0P516ajE9ynrJ98gHOFvEE2MpG3IJYu1V3j
/jlsdpcLnVk7mAOVFcEC3B3Jt8spi0148LcTAcD/4MMSljvkkc0EndKY8fsBtfvkQyTwBThw9Sps
aJn8ZEOBBOjJKgFeenMx+ieaZGKkv+zdfYCbkgYWM++A7j84RaFQLL4zoV9t7F1gzrPywCNDVwm9
LKqyKzIBukmwZG5C+2yfsI1bPHEIZxTb1nKIWjiTfcCrQQssVDKcXt/LdzBMJ/C1rRJ8aiUwizjd
qq8BlNqAVWdgTAbd0D0LAibRzyxsWZA9PDLw1ZbDk70Q7T/wMCgPY5Z/JdqEHOaIo9iJnPXa9PKB
cLUGz8KuqkoTBwpg6mzgxRxxNweWl27eT6QtRVhM02mVjGIvGyQo2SdNWWjjOx+8B54lE7fo2XC+
7Z1jlTeSanLos61HkxyOAj4R+GxFAucap6jkP5wH1ok3hwHupgBpyDGR3Th81rhHk9iv0WBhcA9q
x3ht53gGq62BXKbtCD1QXljqftph9uagnHQQ75zWSM0FReIxeTDcTkY/veKh2OCrPn03gmT0r+NS
tlSYHnPTrPU2V7HfDzP+MEpj7SmNJqqq7fN6jvj/T2xDQvy1BLPLcflWKSJ5riGKsqZ0p7OWZVXQ
lVBn+7imgFKGOsCBSQiF72gcvLFDOJFTosWp6+g3GN2G5NjlfuF3596iQwylZKX30r3AcbscX3o0
qEfnCa/i3v1dwNJWeZt+Ql01qqg6WV/uCEEXoUmeYAK4Sb1++X9PKK2WSMq2ZK9CACK7a31+oyCU
riDDeiSUsvPUGvvbGj6lpqJAEseyUPLdKj2QpPLRY3zPX4ga9aqvvXZ/1fccdB/+ZtNNnEcCmn7S
5OB/nRmgn416kyXhP8005KK7JT+/m18qnxWPLBMpyYbhxW1R07ZBWkXgqVkuzYKRkXveLVvzVr8E
YYedrmaSzl+9nsvyqOoLt8JGrhKUio3QDc0aNyh8HTgER6VxZzclVIgZeFMQbrmw4p8EQ52ptwiH
DZ97nFa2ZzdbD+uVcEY/OFoWyNeLFZxUy9/PrDjYvWDKE7p1LxYQ9VUNI5/jFpKye/LbQhKRNTp0
p6MkIUTv5MJBBR+jkc8oTLxI0j0MZBH43hhh2jp0UM9P7a+Rl9CG9M5A5Jb1nmB0AzoXSchdSsbW
n++izAW8r169ekXZ7/SsUohnWlJR23WLGqLSb3Nzq+z0xSsgPzqiSXLvS2Uxi78o0wN81wPTRD+4
2KC3mfwJwYeSMUCZauZ7G2jN5vllcUAjQk6H2cIBKIeMxTmCbqsLMIwWMt9K9wOzaPaG7ukF7R58
ArqNi39nDUb73A9yxmw43OJClZNUhQgJlvQu8ML3eIdi5XyXkPe/o+g22B4R/REy5rsmDUbgoQvc
JurBnVThCaOYMLxeWIP9rXiKFVVxgBwWSCpLhbgXM2NzZDbi+7jS28mY/mm36IyOhjc/Rv48/ur9
1n/M2Dn9N2GPO3m5hy8kp+3DydixsHYdWWOpBm9rUr50Q18lTZ6TIojpBBU+9TLUP3Cz9bNHfXrY
VdE33z+sJD2SgX6tfNLRyucgDvoYF0+bdnbCtjx5GTFdCTs+jMnuiyNLaMGEbHdPTGGA4Baf/0dT
2tFPztxBimrhN+McRrhkzl2um/LL6ygkJIx76HmoeyQUl9sF+D9oWbnWMVTZk651mTQO62oLbRPu
Y6VshpCjwaENGIKXbHKh0/A7m73BEOv4+vM9oTIMqM2+NZLAORkf/5yMQhSxCtKAUwL5XcwMz5Jz
iJ9yPq8QQbSL6Soshj077ii/Q/qpzNNshBEb0+aBVaz2ujZ2Y4fJw+4WFgcNfTc1ni7PZFW5wx2T
4mGzNNXh6ieV4yZE6YEtEYjAQ5b+11JBBvACdqMt5Inr5J/maj1Cbj3xS4KoTtoPk//WLRb+rO9U
Iemw1s1Y2y3aESrxNWdy/DSNMKl5jO2vR5rbvQJEGtgQ0rMbwXBpVlPUL+1fsRpydEiTk4DHtX/I
faT7y3Q9QIyLjin+E+Gz/pJdVrCFShi6/Up0qwPchwy1WksFtgFhOOsP0tuqeakU7/d/1MNv84Cq
UH0xm25G4zpgln6tHcc238Xv8BCODx1TZXpDH8dyklgjqpLQmcUSKkgtksHyK4X0I/m2MXL41BN0
oP5FgU9JMhMDRb+s9OkBg0jX85uY2xq8/VEdbCH6td1gr0f9g2/DOSFIqRzLVovLo/Da0a3iOLzV
9YBxINuJCBYvtS8FI9lThsfDjZ0JcKuUrX0I1t1pG4Rjq+66esZX3VZpWRkt7ZBNKGUnMNJkm94f
adgUeqpSmiw732OUTZUkT/sYsn/eCiVL6wGFsSRYvLi/thDUBMvnX0oUg3Z2MCOYMybmhGjaFOYn
ZNQE5+Y35Inmec68fyjqcCi2PAXw+G/Qwx1XB5K0cncbWlunVxHOL+hue8rQ4T8ycE+zPXqjUJMJ
8xhWFmI4Cu4rZT2HSKikyEbdLxYuvKpMvYL3ZJfM1Bhsj6Nx8yJyc/hdFIASh8RswZxSmvK/dU6i
OXiD+gdgiW2baFz2eLRIUOILEI/fmBfed3bJNvotAH6v34hHhshI2NkQcSHrZ69DC99Qf7uVvB3o
2a+LsuAFEw3j9uHDWYgOvuiwOCFYHkQe7U1/bPFVT5Xgi9AXa9TRhX8Vzqa8u3pU/sJ0YLUx+8sC
32eqzKDXKwp0C6hjDOzB3AbVj7Q7NoOHCzCaNSlC8RClkLX15tYwh3AfBFPLpb7xksFxc8WIc1eR
21Gu74eyscLjK1Mq9QpXCsIquGUfqHYNVRXJUcpCBy0XrJ0DjyuLkYu/9VhUDFm9K1GZgD+e+etY
nKqb5g02LhEXm7aeN9WqqjoO3hhv4V44n2ihKjRwvgqO7zgTgbvCRvMkJDsM5WpW9K3qWzO5JroB
UsXhQ59TtX0MS/k1jB+3XYgT8qJ5uwQAjzZqWuIkhJrDeKdhbc4bcxTywA6rK9mIT6MHm33HeGB4
PSlmwAAfn9pzTHIUJWxb7aUPWzOMQxSnZnDIdT2rPq7NxhoC3a3WFKRkj+Zh3AV4fdS+33AoZigP
0jtUm4E4gvu1DhL46dG/6SfJdQYX3sOC/UB4NYzZRZzwJDMZnr8MuCsva7hmp6uuzjRzlGTJF5J5
kbSODGtT1PIzoXMPlX6TYpXu/rRoMtqJyO6Bk0bRhEzK5qkhZU0z5tt2lta+sCrkJbs0T10Ixfb5
Y1Ynfd4V3BlIjYO5ZY8F0X9b00vyD4uz3aDcyrl31H78nSOV3gmPmP5v5efC9EZNdlGdXjB09QYk
Cv2i2+sXzivsdhn/o0w6qA/TL7dsyKx4Fu/1sxbhoXVfJMNc9IRIxI77ms8c3fQu3OlMerd2MmD8
JBJ0r3ESD/vgWYmFhomfpOr+thFf70+T+kUTq1J8punNMB+y0jAXMVREWcvgBSsGIhzvy9lsl219
m9ShY9JDyiGEs4z1N2PPTOa+FcY9HBUbFiCydJ9v4pn9hFnB+djpQiDH+3ktTK/KIZcAyxV+WtSj
QPblxc0fBsKwiSAhDtdYlD6/o8ApIxSPY19682ajWtBGI53YlcqancZnhaFiISpmM/MFV83j0++a
FFSaedgGNb2mWR1mAJ4zrihWDgnozLTJzNIkx8BWMAUZV5XC8Wo18k6ZRdP8RMO20OTn4XUFGy0E
Mxu8BPbji7iUqMOOG1W/vB/l/t9MaphXtw2CISvlOqKabw0J+OAHXkeDTtHJATVVNzon7RC9Doit
axvzxx9upKACG1JDM+X+yy0ZC1VkmFuHJy9NZlgJCK9AJZn1XO2VIEUioVtMo+49oaRADaS4TCuU
ruC/72l/zoxaJFdVrRqJikMRZe0S+bHVbCxQOcJy4Is4gQp7jZGroFLUGYAblHtY2xQgak7LyxYR
hxVQnphZnm/DFQJDSENpk+QCdZtIgR6FZT4lo4W90ge5+aXB7DVzwTi2PJMdyOrNsNMUolNCaKjJ
HfrAjvHe7Ba3S5bs/RSPIVuByXso4QG8rAfJMrsv/xcHlru6jC80aMUo244GVEvs9gJTGWNO7uPs
5mhC07zoYh+dIfNNDZyJAjpMDeEaPtP08I3zjmRQmKDR0saWWZ0J+VThaSVuFO3SmiraDjOAJW6L
ajj3fQdUmGaSfqgHu4VxQxj/WC2n4h09CUQhiOoFfqE4PC+M3wF7zewu20XNnAX8mXHOLPiC+8lb
IMZITUGP+fOnbOm+tWiFNg6+MyYIU/qhpSoE41LWpWL35ivw9dXEbNz7E5iAKAIDEbe2cUiHdjOn
tjlPVg1jRC8Zn3abaVLv98ycNHFhAU04wWCLA9xFpDm1rOjVlNTOKgI4CMZi11USUdDIpURZId1T
875ratvZvp3oh2Po3ypeeKAyq6L1T1uHXxDdqvV9p9gkFTgsbXFxxZhOfO7DQm/jrq85hkVkclnx
RQv/feLQSEcn9k4TSLP9+U1g7HSzJCxccWnSrOqsVkVldIw6AZ9AfGz2m5U3lRij3mMzmkAV/z2m
pTbHVkOShaS76ffxTdWJGwvzsINmC0Npzie6wOQ8WZ1dfSwq1YW7yXzsweGkqfc7PZhd8wthyHWS
RUSXYM1/KWH7HX+0+EQZh8SaMKDKZZSQT7y/tICtqUIeJPLhcvQRHaY9eho+sYmlzYUclu+y1Bzh
Z4dV8h0CqL6sr8qGAfgH0PEbE6/sdu6G5hz6KwYqC1dqHlqIoRRpHwvc/XJp1X+IpTjzORBKuibX
yJCETN7a0qLNgssLnvsHFYN+Dzv/VWRPTwDeXZPfGojaETm0vOOGx4HGamLqPmDjkjfXA14/U1sD
CdoFHCpVLxoPXeedyylGv/ydUh7PsUjOD3VvDiiH5pCS5njSgZYdcUdm9QJK2MMQVsRGTGHdYNig
tBdN18syr/c9v4LiNjh9RxcYIxc0YD11P+16a2Ht6lhGR9KzXiCMmd+8AOPMwT3oudl8OhrC4U4/
zS5fiZD0hTSTfkL9ugS1zDyFs4D7a+svdbGWN6e+NQpTiKN+hU54gOJ65fdfjarFqKwLkLn8uMix
bHNhaagcHXVaHLhiDJqmlplNmcQK9lTO1PzLqmFiK9hDDLqI8zs/ZKsb5uct2+Rm8vu2sZyEKHHB
pcH6x06pVx8tc4sZZ4qfipi9uCpuhbGIz2wG7iru4HZAmxEwirxUnVCff6Mn/ltU2MBr6Rp8Sc1B
oEvyolKAHhYJLpUAz7mCEHkyHZ6sgymtB3Y6qnspL89/UmMc17rkPGc4hvlVxzLOagR1jbR/GIty
fZBVMzRZYZ33b4tAIT4f4G04sj3JrwV++VsBZDkGgMwajswJqJOVRhVZVF5jIVUpliKn9xXhqjnE
svN3y9Kz8wlUge7W8Tf/Rgh+2/2QC2UGg9E+T5tyvWOXtsuLPE1dEnyVDDregIUGdavmUuMhBXQW
K6QLfLrpP4Prmv0wALVSL60zDZpAyc1ToO52ZgqeLvFPHSpEExf60nEyC9cd8ujMc7WNMJj9NYbR
kHZ6lLJXvjZ7E0bzf0T2inBts2+jFYsmd+qylipWUOzOJdxRyNj2u50mnj0PxqQVC4QHiAFD3IGm
UqgQr9kWVJC2q5L7NH3sODVB1ZY/3/pjeGemaV6Py4IdgRElijnCorwLVsOu+ssnDKNwl5DNmssI
JZkb6BYmVqemPPMGGw/RlFNGmY8Cg474jwWaLCzkXHH+uibJh2RwUKGB9/N9HLrag1C7t4AQ37Da
5lc0f/QnmE30DYzM5vqr7HZsPTNsrIWZP0rDgPNr/VX3qr51dmd9WJQ+FpJVhAlSTOXBQj5LuM1w
w2mT+eAqFW9kgGCRc9M3/SRZUZDFeppRRo7i6kfmDbfhLf5ybmniQ25USsHTyNit8v9F1ZfMueAR
dCivEPgNjFwdBtE0WQjChmQMUh25ZNYRBKxWwp/iieEREBGk8V8LRAuF9SPNkUWmFV95AriRoofW
nignj7extAOuC1V2XgvxPnrQxFjxSeA6UCsWA/E5aS3excP8+djW8BT5sTSYnwmJ9roOCslrnTls
nPA6gDGIJXvkIl8YBRb/Buf+64s8hh0YECgyrL0s0X6rF7n/Yt5ZFuYaxnIHVc5/c/YNwwurcp8I
bkAU14nUVl4ls4hkH+vvF33QaOG8qjP1QIQpMx3yzwTWkIN9+RUfIXi/uGdAuqXglKda2oxBcfEo
Zex+8asKpkGcWWm6axT0hxeDh8eEam1D6X8PI2qzKugPxYnpWdApj7vKBPKjijD/qtZ5w7kb8/aK
DVOuKodAB0Ad7PFU75hBBAUUFEEBLrpCeF7i1x8+ahHFg4AvVpp3zoqrXgLoqqXQTw1uwWaQLBwE
hAbLVeaplV2yRuGntNV42XVy3UTP6OE6gRx7vZa3dXqMteP/A4PsJCnmSJcqsIPnJi1giUg3r01Q
l7zItzfrjwyGo+CtEfmVSuTft00tIU+RkOXuC7H2EhC0aza749L3HpMclHysa6NnRfKx9zn+F1vK
9QkFHcc43QEqkasVXicTlQbGUOFxn9E0I+nAQsX4jCJJqFt2OPn0Cpy+A2E0YqmYtIWltHhvwPQm
II6Ctvnx5nQeIduy82yx5VF2fHaftijaRM8PJ9SMMQLP0VQP0rjBnOsCJlner/pyNfgsDg43bmAR
4w+6VNididYHgxzEEoB7cLtMdOlEUb/7wmuJndxHM1FG+c0vUn0HduJLa7OywMCoZf9jef8MBN8z
/cPm3ezi/DnJkz+F0P+zfSLd7ey+xFokcpOClHuT0X7soADzvcjmazRSklNOPdMdmeS/Qp6zQFLS
V8yQLR809evPIsOmbcGAJp6aGmA572Y8H79O+TTnS+UXRiituJywGaCu38RhPYFcZJjhex1KyVi6
Lfv6CCVQTmtxlUnGkpzMiHvaOFCw24fFwzp+TOgq5flXuJxmO+Xy1Cn9c3iXijvhTrxDRFC3GGmQ
CmRvjVKHKVco5LIOCQMt/PqWnPvySR8rwy+cj2Os4cFw4M2tOWRpKN90+ePDXdzyK+2NlvzdxCXD
LnwEMFZJTM5F8AZJt4G0JuLJuKMudclBugYNUovVy9YpvArPnp7B+0166eKhdk5jAEIyFB0Mv1Uu
lgdhpPlQpoGWUXt1U8FTUZ+nWnZdY2SjhuToxGtdSaXDceSV+VGA53i8zOgY88F2w/OsyJXI6bG6
ZfJz/ZZgqyCWslE57TW014aJBMpULjmOKdDqFdvhJxpNatOHS/BsM4fjyp42McBuwMlx2MLg5KC5
0DworfV4VKhAP5fD2kCT3aeppbcqyebP81Lgd7kZ3B+ht7BUzB2QN+ZX22ZG5Vn9rMc0uNYvxHW6
aGIR8SR4NQLBeiJmPr95S4m+K8QzSOgNzxmh+mUDa6XMgTJfkgLhqp2I44KgoKoGeJSUIC2Idg5x
hY8ANGt4zm0b1bE3AeFHlbGbuhnU307pp2pGMbYxIdhzMJ8u6cHGnui+5rOOjNZwtgcL8BqlvSN2
YJreKmiIbD6Rl9tKRMVn2Pyu9ghm8n9cdQYXmbQP7gHeObUzXX3s7YJ+yWI+bsgnNvDS9oR0xrUJ
hxRH+XQpustFBvI3rbY8WgDYX8lCJkhYr/C/T/GLQOrCoDBSRvAzsL4JKpQsi02UALybpwQTYx4c
4t9i2m62fGEGpgdy4+jyN92bZw2wwcoTJAwNv3T43Lec08UaPHY+CPR09T6EKEUvTjdptETL3FA4
6cJOHPPec4muXSxQhdFqKdxiCsPfuf3LGilaMIxLPH9vtmdkprotzviP0JkeCdPOQiJKJeqWdI63
9WqG8a4LqrngBQQY7lVqkP494FNMKNqxoBbt5p87bDQR9tXDExaNjMkc1lKzIgPJE0ooGospz8Iv
vHle8knbjhnj/Shotruw94pblOwybM0QSGzn1Cxz1ZQHj9pTlifz/oeoqWfjJN0s/Xla2QDmKHmj
0AdvWEcANtB8EfEWdfggYLXV/1p3QVnraSDXTOTj3SazjEysp0eSyghheMdfStjhTZkCPEBxkerY
rytsL6nR7Fx97x1bT7SDhDMUuLG0PXqcbQ0p7wUDKcvWKfy8fvl42uv5JLTa98+MVHxKVWdM7dEs
fB1lmFSjMOlSJSxW+UiRxuYnh0Jt36bONumUbIknUQOLUnAlrLnVtx0L/ZQJGcVH8TYEIXT+e3aH
6/oVQc9EM7ZERuJckc1OAZHzc3zvtmhOqYixCTLEOLDZxGUuUcAbUoXT0lW+SM+qiWA+JaUfktDL
Z0Vq2zkFd+boNpRvCFap/rkhKSP1jBVezEdD4a3qV/JkXSzkPBA50SJmvqSgfcNs0jLpapgtpdlh
ngZz2ATplIaQJdVfIihBZb3BQeXhD2k1s99NjFJYDnR9lcHjavyYQEcx7Maznf3BVNKINK0v8umv
FEhXDxzAFAfEz5lDsSwU2mJ/Jp7QHsVye4PRMmTCWm32gJOf8SKbSxIFJHZLgQEWLbyeXf6jCefg
MwUAGLCa3SExg1tAH1IjDtKk2Ulwdknkg5wrKLu/VaQJ2UkNwg/bsgCKFSPXNS7WIig1Lz9svOwr
kTMIzcj53bs+PyDkotc+0enXHk94clz38oBVnKS7VkjAOwIg0nJmIsf63F7fXniOMO3tb1q1UKf9
Fv6Z3SAzCqzn32uR9RqplCV6YsCRWPN4cx47RPmv8pTK2nwIr7dbMYICWNlBkl5uVj0XmsCq+sDk
53c+IEED/uFQo4aE7UgHHMqeR2ffa8OMGlzJYxCiqbfAtO0dnOqa17/be14NrEzUB+Nj48bUvv8G
lwDBT0JJh0DMOgNlFBOx2mU1uECVrD6LEBz8wdcunpIJpMl6z1H7uzt0t2+t1yKoCAXZKnLAXBVg
IptOpAztofAQzfRtmWNgVgfh+vzVGVj9tXimb9G6wvdXfHRzAD0r57mP3+iHtzUb9QCgIKNkNMCq
MjIjmRElIkKew3KJ3z382YmgseyvI6YRmKU8IPzLLLW3E41tt6tjfObNa+4Zx0S8nV4SFe8V8uo4
0Epx3F7HrUJmmyYBWG/Rl8xWEVaJzpu1zAD/0hJMdJEsBp1rnNaGdMIleCB/IRBmcROKMZw0MqT4
W215+XPd0tK4kWh3jejJfMzQrwJI+jrtNHFSuxhvws3HMeT43Wig81TnlMD/+xx6hM1Yh/hUSL1o
oZLZ4p8iqhc2DHBY8DqD7n9NlLVgVOETKCkwJ9f+V8MmsCN/h+6C24OimRU1AK8ow/4mjdOHtPQV
kXdZtP9rBWfhUndwbAhrY76pDqV3tLnYljftylCuoYt6xDHIydpLZoT+BakIgz9ndbjjzOfBt0KN
M26Ca0UbuTI1K8qf7MCMWJ5tLoK4IW6uEHWU/v8jNLXIHXJvM4SQAZXf6t+8naNvf1wZvom5EscZ
gkHOrRAMuMgkbhO/gdjKSKFfecxaE52t5R7m34bb7bdG6LF/dTK3JaZXL1/giVdhQJU/CNYqBpJ6
LGRBLTxvQOrIVE06O81eJp5GBRj/kFv9Hk4Aeqahr6qO65ck5HFkot8k5Zdsb3IjYg5Is5ndIrkD
M2NkA3O2er7ANnqOXbo0+kwDoc7pRE+8BeTFVGhrHnPaXKyBaMK7j2qTJJNn358l3ITwP1WxIzLt
vWJ3HeCkStUjS6K42bI7EdNV2JeqMFT9yqyI80f8zBg3M64oQ5O1DNPzXQ+znDsUQEc61N3alU1N
OFWsbkJ9R072W9EagrFg9t35tVzDpN9L/TLJ30hhTa55dvyXIt9NX34GP0bmO2AV5oltmD5/y66f
dZnxp9Wyb3W6lDjOTj5pSLpG30P5JAlkQ4sCvQieD1Ph8iD0PE95IKIp7o0iocMx+HUI1mpvQODI
WGa947DvggSQRQ9yGDNf0eqFQGSCCi7112XaZ+c+Doj986sdgR9fKKwTZEyxRNpB7B9Dw2Iwkv2g
I6w6NTatBygkehaoAl7L/YPm/IaI0BSq7DwSPQIA4tC/xwg2nEQahA4UnUh5s0KiG+67UU43DQ+Y
vN3v8hq7wZ+CZCBivenIky/gtmQQ5WWa109k+9JeAaESP4gHG16Q9w3+tDcmLnSTyI710gUr5Xhh
do4ZhwD11H957FHRGvABlCL203JXFsXbhrgA7F1s/JQv5aVLHUPUHVjaYST+NZn/FX2k1hXFz65O
Ug180gBy0g0Ke+LivuC1++V2gr4jescuR6Oc2PbFeEOmYH+K3tImqx6zAse23OvZDzts8m/s2W+v
uH/GQF6Qdo97uKeWEPY7qaHB0SWXjgeUHJDaeyYDSLJrHK13ewb8lITLaKHsWmPeAPjmONmtLom5
G7OvDDgqzmBdbQkwhoMk0p3qm9vyQ3i4prisr54d0ISvVS2/eXJO/uLVuTLLSVC5Xd0U9go46toS
txTS1u2DdE/xFV9nj75XyuVpqxleJfnbvfw+PE+ENmpZxdL8TNHfDkoMRqUj7cHFG/G5cKRbr5Gp
rOg1qpQnQSA7qvULeUzyYKUFGSsIKBEAFektnQn80LtTY/hw8U18rP7O6yFp9NaQYmGwBEl+GF/G
1pWE+wCnmfXdKoSWT0j7MXgFAq9hi24bpT2AuEWSCCD3rzMejwtTYAEJ45H3U8Pn4402XJWLGeGt
cUNeXBzR6RBMj8u7y9HXjug8PM5HVgBXbBYBOAqWbRwiXf0Z+T6ujQvWs9TEo0WMjdwzL+BO9grk
5pQCKIfFPTAGk+Nq5z6WsFAjguxI+FseOoDHXjKXA/Y3GdFs+zJA47WxjJvRGxeIK7P6euuNVoB7
TK9OgAlgZ8cH41cPDCvn09wry2Ch5BZfoLGL84UluUu9RL1QPprCNj0OSvNzQpYcfmWpdSoZwllN
94a7yKPtPbvSUd7QjgfqpNz99It/NEJ9cX+klbKTRTR9UfVcLEiPXj73pxNrMiB5FtrppVe6Zd85
3VqRnRgFSujBfiZzEwUs5MB87YOYa6VqX+H10YyfR7y+DaVWJW2VqmfbpaiAKeB7yWI2HFohCkMc
XZl6AadzcMalVEr4UZQuUmbQDnuLe0mUt0LCw3+X6Dhkl+8SX5mMyZx8u+u7qspdJDeZk9z58ZZU
wlJe3nwNrmAP+lv7q7Qw9oVu5vKha8uFQs8E3Q6OdiUmR2b19USVubJm65knqsGaY7zYhVYKFlaI
a7PDNIvn/S6vQUN7tvRbGnF1MBdFmNO7ar2fUxRGgd5BL3D9UzUJiPmnI4pKriA+X/jc8JirzXRv
+zYTMhIk/bMQjJ+8i+TuLVYR8vaQeb/c60by1GEg/QjU+iNvIcmzXyXgAFOSJ3uHOiXBlPVptCSx
KUW2QzpsnWYBN6gVXsJ+ECxUw5u/PwSC3AXeA1XRqtfyPVz94j88yLVkHIZYZLE6xjO5HT8xTcHG
16BsG9XPmVTOjSciGtyZy2qtJhupDIJAokU6AyIzyRVCXpDXiwdK/coxU7fH6QSI/Es4hP6bixD0
/JmCH+5EFIqdbjPYh7h6UeENi0mo+w/hdNvIPWjfNF2Rf4o/3XW/tL5zWybScuPokBkZji2SSmnu
WSwS21GBZnNfBzaR18MPD4ZsAuVwBP9q42sZkQovfhWLtByiki5XJxK0r3WRy/OkwMln5pxKJhGh
RofmNbWORwzgfslnQzFROlaVRne1o9Apgx4d5SFymqZR9UbmkhYLPhjaFSkRLP4elB9xJK7InVbD
rXUXksPzaVac0XoyCRZzEKuvGs505+BIvk2aIw+ypq2WZV5aEbF4gGeyVg/gRzgjfg9zCL/iPz0+
kGY5MQFEfXjjv5wEAPeKmFt3tE5Bli6LXqO3ghcEiFykblwhM4/comz6ml0eagxGxABDq9BVHfPQ
x5VR8u1lqqhPrJMgPcPgOF7+KpkEG9SfDbU4PKHVf5NDkywFd4T6OQ62aBXhI2fnz0sVfZNLyt2n
PFFdOoM+x5oawgCdPx1J07/Uw4rvIZwXPRzONAdfyIAP1FIROxSc05166gfLfJBw0r3r1GHtQsHU
T9izM6wHSAjsq2gW9F+9FMltvsNEZ8hOdDVkgwoNaPPcU/xPPyE2wV5qa3x9cUJbvlASn1nDJXbH
VTXHqz2BAkASDt2Tm2cpD1J9rE6dCCcXkbBhS/yICvb8H+KRdOA6Cpc9HWPSLU2Lcc5aaoaFLlBo
S1yGN1lRueh1tfhUuMSYww4UYne4BhfRBTGeR0RiVha4l3GMLnlmcqcdayQSvSELQiHspIpSnz+k
ruRjucPpO+Q5j8E4dg5DoanluNAe0XbNbQL1AbMPsOtnAOn6glegP1fyb3xupC6cQZjQ11KfZy/y
PZW2aDgkjQDs2G0gl+KZR//cjxowmSXAtx5xOybgkR4LEk2RclW1N9+V+6Vjwf6KvZz4aiQKfIbq
ckOVSnhUsiG/ll2wjeriwi6lrqooWAJGauhXrLGgpadgzHBaY4pkdH5rcZE+zMGQKg4cX2W5rKI+
nELSjy/UL9n3Jynj1ZbuIQBFqhCC0yPipl8gW57wrJA7LVNfLRh3Op+5PvC9K+Osy1HwiwjHtP2E
AkntbPOyrisLdL0BWGxPM6vKfd3Wu6GPBTxMv7/DCMVtrNXJI2DlqJjz11E44CbRP9aAxl2rnaIV
/L7vtVt5waGdAGNSaLogMhEkt31fLErKRcBautixSqF2CfKF2bWqZzM+Vw5+bIgZQ5yEn2c4bxgW
P+LS55OpqdcwXsisRPOFr4ShMhsjO3+Jsd1aoYQUqGQmrstLbOAAgOWIjuprLt/jaYfRLTYyZtOh
ADXJxoCE6boOZYG2DkV/Ox37PwPi2zayU6/d1mrRzLSzzNgZkemxDhZCDRzRg7Ek3ZdAWdq+SnvW
XppWCja6+4nSIytrDPfqC0dNi3/WvceznHnkL7y9dSTl+q+gbZ3wxaR/R233DkUd0R/LWimpIw0D
ksdfZksxcQZwMBcLQrfhoewLFIEXMzLzcWtskUiooVDXQKpyaNfIPYwqEmC8yuYnTqam36mWLaPi
2c1+7AEixPjts+aO0JR4+0XZIW4uUeyaOPvEiQHkT1cN+2QasKRPzxCy2rO6DNX4Y668BXOlE3C7
VqyDHwklbDxzUpgKhSVHuriOE+UOsh1ys9ZX9e0LjfOrPZrayFeLZeq6PXcFsdRvxc8dKiUZBccp
ii6E1OhxLOhXbFornDRt2NbPwGtwVVQvFWYamYpNstuoitQW2OERZbnx0xf74tSHbFL1tNagmEPE
BFezbOubBoK1KWm8yLKVzzxyYrxK3DFfAES5Qz1lyck9Q5820aRNLvKA8nlBucmniqVyVlyp3BLN
p+QX7XBTQyX7XeQpFOuaRabtehK5Ifj6a3IDiv/p2VnitDOlfEKVeKBWdOmt9HnDV6NaL8K4Xm8q
B7wmH6U98NocZDN/lnozTt9xz/41wfsSQJ9rm1zyyNd3R2KN73MmrbUDWIvUwPJh0L9OGEVQjIqZ
MBe+IoJjvlNEz/pSn5J665cUH2EMdLuOMPU+9kE7dlvnIXC25fulmkuDRL7ICfGnGxmUE0Z/t1eL
XvYJJC4I2dXpQPAOCMzB9FpkqtvZ+N0aTvvhc6Lt+848FH+x5IOUXgS6ZIpOBqrsCec+TV82VcJx
5Y5Ia58pXOMkAiU5zeNuEjxfSG9CieSyj7JgOOETCHgEfqMdmjyELOSgQhlrJLNJOnQKi/vpXkGE
tFhaUp41+JRhzrd+NFsFZ2e7xNHdEjxZhDXXZXbgkaJr0fTM6H7SfD9QJPnAiOsgC+Bb3MYrFIcw
T48XtQSMkMqHqL2yBr+1qnobLOrmkHkoqPTb3QDVr2XPlAyoDAUFus4tGv3d94uV19PmJWp0YZqH
SAnJfBlm70lDFBDKVzwXZdKX2se7t8TG+RfaE0Zxg4SS2GqaqgXS3a33KtDihiwE4ytQIxjA9dKM
lZUaTZ1LpHFlRwDuYQ1Ib8ryFfKCWjHSuj8OGD9CouCN+IUnhg2PcRfVn3Miv24/cmtotQS7irOL
0blUeDfunuxSVjQoN+Gg/JYi3qSWD4DOC4bp1Lb/+qz0HkE1TVUvPYAgXArgYbhzBVKMTnDxb3Df
FuSIY8TdnAh5Fhkx0Ol6kmGPaBRIGE+CA/R3xV/C8J26uZspoNXjkZZZtsHr2kfvgcUps4eS+3TB
4wDs7+r0u+GBlVbmBgJnktdF8dikSeOsv/UOfRpcMm/l28aS8Qf1y3MNOgoiyU3yQSlRQnFVxxFm
EhBj1YzrzEemFfncOoEzfDg85z4G6+RPlrhQq+ZifImhH52v9q3qRrJ5W8D2017RSc4GfE5JoabQ
E/VjLILjr5giWFW6rRrrKviobwgS3Q3d50E5HNb0UNIMjBz1wZ8OaSMo2Aor/bQS+1sbxft82OF4
h06HbPNb5o9DB6+KaSwkFCZk++qC0nlvB0TzBvmrTmnPX43246vwoIanmQ9iFUZmfGo8W89xVgKg
p8e9amBGlyLF4w0d00g4IB3oH5jnqSZ6sxh/qopxAbVxLVCUphGJasuf49OvLl0Hjt5Mu7ooFce/
UGWp0CBESZolxMYVaX9DGN8tdsjO2KQIJRt/vfLJPuRVa66eEbfsa31E0lJbAwzYm/dtfSbWR6Z/
VAc+svtsFlTtUKA8292fyyfz1PMVgxetFuky2jGZFxZ7I1WT7rM+8aCPNgo7uWuyR3DYVqTyANXH
aqgZjvwaab2p6Fyb6MB/fCk3/4DB+f4unwcBhro85CF5qFhQ5dMp+8yw0SJt6Gf9ZdjVPBjlwUoZ
iYDMdF1nJoZVfYhHsG1hqyIlAzWv5iPsbXET2+lA9YYvTHaDJt37fJLiKFd/q9fy+naf4dOexO3u
MOJk9Lfqj/gR5XOBfNqzK4XZ+z2hwOtO2VcGmj71gLeCED+1B/oakb7ZYkk5qrK0Wa5fplfm1Bs4
ta9M9ccsR+kIOzeLsJA/QuabVFFHRR1H33wOSakBQVrNC0A2kyaft1KzSa8Oad6P0kSl5E0tj0CG
vc3Un7BpTr420iX3BDn/HilLV29d9Ca1gQH/FFLZ22nO/y2WIF6SiXLdlfF4Gd8VZPMOagNQlGQq
W6c0NTx9/qx/IlqVMz5zBq2wrhqVu+4NScUX01heOhW5KaS1IG6JrqrFzyXVRUY4j5nTT6OeMUOw
hZU5MHS5KbrGM5PXE0EVHimOahLCYjr4+IoMLH/Fh4fnWj3EKt7WB/bnsfNT+Sn8RrpibEOSn7ML
2LBuIA9nJHUCcqCTZLuCcor7YOjoDR/arSHoYm//28pTQFBAklAAXFVvMN4AIvqv3BiJy82wyJZn
bg8qFph62mBRSq6K2bJBJLZsMRQFkUGFlPQburNpbK7VgQgNqD/S+zx/cwAYkyqyJYSlJ/mmEoN0
+fb0xOCxzSX6NYt4j1hCBs5IQOWvAGaBRNl3o9HuQ0fpfXgZkfOb8Hz74UXHTBUo0seuG4MwJlbl
V89YOuGjf11JFKz1Hgg06GToeb2g6vuzqR9AZl56L1YhwN8EB4nLPVK/PqOMIIqjdA0eKSh3mCjv
BZc/0cj9rxuBib26JzYfU5o0CDrK0e/3U1RNFnL7/2iTLv693flNLjPi+LmlvWUvMqe4HoNRkdxt
aKj16vikNwiepi457dL6ubFf1b7kGgDVi0xCGsV8P9elleoAo5Yyf/Y38oyGUVV1+u6xAoaa2XoY
FhxQxOYlhNjn9SKYz0x4IuDCUUROlLus3gL2Vl9JdMAq6Q+PzJTKh3QBnDToo2vderuSpDX81Rke
vjqi7jXDYgr4SABZoiElyKViCFCTxu1l6EI0WSLZrCkkHDTRoO+yKtryZqd/CgLA+S3IQ5vtmJ7y
2bQzMGWZptRqbvjNC9Mmt/wqascbUntKSbJKNdJ/pGLguBkb0SBztlRUArrU16l+EOHon72H1Aat
ds5xACefpZbDlvrpKNFSrsS4qk1Tvxip2YVXrvrNS4J4GYPDms5/THX+H7z3zJVk/098sPzdX3PF
uGJi7fj8i1h9jPem7rzXIf4Hyn26k6rzbVXrmdeOHjO6KwDCzB7IqhjbZeWiahAwiWdXQJPls8Xw
Au3GyQFV67Oz1BfHvFZsZtkaj2IwdGmXuMUkWLjNOI11fMxgeMFg98bH3r7MfwR4J0vIE7tKtgHW
C81wxTMVf12ihoQDfEswJ4f15RtgyX9bwHqi39AbupQJ0Gh22vFcdd3dAsSSpeY4kSY7MbX+Mk5v
r+su7Wla6Tf5xxUY4jbZrM6X5XTxPsQSDFtZcQv0AA03wAxP1wX4b5ra2H4nbeo1168l5QOqEjMv
s2vkcsXa/t3iLjFN4Llx3ovSJFO8+MOgie6Zjyc7P0zP7lnG4gg0gpItOKv6GKKZimjAkc9Iy5oD
T0eQ9X7mwqU/4aDY1MoPS5vmOgAk/3/Ezlubkw9uRyxQPSB/npDVl2uzbaw5QNBfiHBRIRqjh2ab
N10FlemuJH4VnVLA7TzaCHb+FsS/BDgwspIZYft87IT17JI8funKpZcQBfc+FxpWrBhNg//HOpXW
aiBCJi09/CXRnGAz1bCkxCWGqCA+YgcD5zUzUlKKVcErOo6EAeYUNjMNEzuPGHP/StyAGyOcl+uU
B7182webeFE+9igbRnBGRM8QlxuDNxI1S/Z7zJIT4iOwOD8uOh4QEDpZaOxsLIlDXFV4rCpTnvfU
okPQkR5ewEp3se4dBRX/R04UehftnQxWM9Vd4k49jgFjgsqTpvdxNN5tssn7uAnPNGGGi0MjYpnB
b6zBePRChcPdVEoNpzQqKyBGt4yt8nIjBbMQhEYy+SFvZWffRe3eOg34StS+opwYXW7ogbkR+3ZV
e4S8W2jvzGueu5mwq8I2c6mOvmfJZEjrAzp642VhXq//2nfA6MwE8GIae9iXMV9ZJGZGnf/E01Xy
nhLjc5isDRZ+DPgKa63Z6NZmUx8znpN2M35r5+tZsE+A7O63uE9GUqoJEcdO4Gn5gu6nx3Je6LQe
AKbZE0EcupCQi83zfRO0FdeKDI3qVA67Run3hUQX7D2Wa9B7M90tx56UFm5ZXsgKX8aPCHlsgZxg
PR+CQL/XaY3Zy3xYmZ6VBT7KCr+bsSBC+z1VRUe9XAczs4nbGucpmR/ag6N8V6MHTProv7aM8/12
MmQnlVjG+qhHLo9uLqscJQgKn+jBDbRY2meYl/7UxZeIsmzqmH+IA/2miBWi6TPfKGps5PnNYa/8
KJM+l54DRiCu8n9wG1WB+gWj+z4Zns9Xn/Fqot8T2HX/YD0SvBdTmAdO210ijTdFg1XtjQIexBcR
CtoZlWfNlNj0QcxTcEFPp486nsOAo9YNuhiTlNL+vUs1tdmDpcvNVQEjOwnVkqWnoymdoiZlb9Xu
j+aGH0LgLaa1CU66vgHAgfeyhwfuK8H7wC8AuZcFC7Dye+xPWu0J8f179T7MKxlNuN31b+8ilYY5
1N1gR72ODKFBkww62Q/dAPFLuwwiUvM0kqSA8ixao+ntloW3EnReIXqBEbGLWbgD+SWeauMOn2/J
Y00nfnggKPfwwa+O6iT5La6jhKn/eC3o2gYhrcJ+6a1521N3k3bCWYi34kycVBtLRfIP6MqxcBAY
ypqRXboRm4hjkpwApIQcvS6zGAyoSIYa7Qt2bwoIJzY4DS53aBd9STZW+l+VDbtePQUZBwIy5v8/
KNb8W6trv20VDL07XaU43blN0owcnEZRCSAtMEm23FLDTK5LKlsSl3IZrOSvPbTfcU6yUACD5cH1
06TVHu+eKmkk8L83+A6Hrgerue0Z9wCcXanqwvdvcJhjZlCyTjoqjOfesHdr8Gr8X1LmHhEI64LX
V7YO+Md3v38rCXYKbLjM+rhHmKUyQCODdu5qd5Ft5me2u9UfOLYS7Nu/0Zk7xCQc1npoJNqj6A7s
qUA0W0r1b2xsgxg7/YWSLdgCZNi2apC0AUbij3mrPY3GrOfspFlUL6Jwj0uVpLQEK68dCZQ+mOo3
Py7kvKp0fihrs8zRfgsWuvD34RDmx0XmxCOy724/acX+m1x24KkAUiXsnUSZA5nILQrK6pgVn9RZ
ETNez1iQYdM/XeWBXjx8GWxWFYVZKDrJmwle71bigzRAMoiqUh5K6FYSyyazBc2N405WDXCU1fxm
RfW4HYVHg0P8HWAsFgpYOX9va58U/GHYz3RLaaMH1SGT3n+zCoiv7kQA805gD0NI2sp4Urtj+C/c
4TlOK0ytVXqOAIxUykKrdIQ8z96UiOtyoxdHiPcOJz3v2iKJW43xw3rvjDXbmxu2ogtMsmvcBr0k
TYxQnhTdlD5pX1kUzH8uKzVl8pS+49tiXN6RVAmDBek2agMuzXHFrNlpBl8IBwfk5CzATsAIcIIP
FU/z0V5r4iZxJpN81f6v0jRLCX7dP8HvehL6V5vUBKj8UFDFyl6CBP1H9IhnXo58Skc0EcAw+yp7
tQ6gWK5R0T+g6LeTvdiBGw7K4n885CYfhZa+TRB8o7nlD9Gr6R1l+D/wYhnxqIMzU6uBXjSEJn+r
umpjwMJWpxxYDnjs6p8z0af1B4nnoCV+64C3CVrqQuG2SgppgYYTORjfJsuP96Ae7u0e36ceVe8y
kXmWhQ1cKUMvHzHvLsXrTfySW6FPydrA7QJEm8NoyJsisArN0texfoO1zdARyNOQIhX3971jPUGu
2cMzcjRsKxstKHrx40gUTPuLLZSZ6ZVXX6g1rB1d+IUC4OpKYc+sgb2rT2ssMh9zfQkUuQHc7HQz
8UzSWNiCFDh9Z800UbHgNXKMyMo8p28CoOlJkKHXPng8GQ9gmBcg53sAx6zdk5WPkHT5JkktoYzN
2Rw+qWxBvwEfydwZmAc1EUHbVDssvQU5JwZ0I1dUPu3fXd1UPu3/N6E5cgFY1iCw8OHsvxDcCfjQ
pDgULoEhCKFZmJfRmvq9RverVKNKlPePiBSNlnjrSm9dRCZ1g6DDV/0tlETC511qEbLTZnyXkJjg
BFPc3iDF7OeDxvlMsB8SyEXOAhI5T4N2FOK4rY4EC0uX1af4HcXXZu7Ch0sKnx8bD9S1WNCNLA15
3RY2hotxE9MlaNXIZ18tQ0ScmRTyzHv4G9dKp4tzgUwN2cCXeFSe/t87YMf3lSOzgFoxN3bdqhbi
wafcY8YLssFye1SCJjdCkNLDSiJZvPGjK2xnZTeCu3mmAxsCZDNHhUVJ4MEAMIXIBscBUehdukXn
h9tPP/lwTMsikj7XNM2nr4dILrksid5EsvwyaSUyyRGxb0ohIbQE0BpeqBP++VKmo6Iqazv+GTZY
Qa8g2R7dDYvDF2qP4dEssLNSJoeuvziclzelhPYrh6EmcJTnfa+ey+WnfduCxcvtj3foqEGn/DhG
RGpo9q3kPcprr4wykftlU52giZWSEeYaKGYSc5tDcVrQJkFLlFjP9EMVDKq4wKFPI4XIAHeNv1Jm
OCDQr/SNkujfirKHLidqTw4S30DoTpLbpbP1k9BQGJLNHq+E4bUA7zxYXESlB10QbVb17JChjeKa
nm3lqB/pxaVgRsV/+Lqqb0f+6pukQtqPVlYXY9Fk6E76Kk5HDvflUe7jBClILiZ6MrOnK+YSXC4z
PVHuQdakauVY64bkEeulyEonu/WYgheqiTW9Oz7U7Y35ZEIecerCkIE+ssobLY4GgKaIUZicxXLg
nvruGlo6XMlHbGyuKIu0jRGaqzj3W8kHxdhrkfE1M/rFPCuQG7k1K0NAmhxsZoVyWEvuQyOTVLSr
TwLkRC6WLWoIbSaeckwJX/T5QN2pbrrnDEPCBrjRSiIkDFN2EcU2hfYTaqrz2WVljcSfuG4hcMsl
TO2BS2NW5NH2Oq1hvbUmOXYnkaTgzt9TI9K1s31tfKCbQo9NjFd3KLNI/UR/6hcvB8chzd/45W+C
caKC+Plk83UiVtmUTQ9XaqXfq7afPcZy8ut04kG85i26R8nCs7thYfcCXFruv059ycPpHFSMH2gu
x4/aRCXAyndIXGtXIH6qLLTPmyqmmpDDsgYv8khddfH69bY1HByKNHuUQR5BkoHi0qC5dNNxT71r
q9+SGODUFvgXk17diaskCRnmOr1AbMBhhITfIpCwbhbyrExmPexH1H0pX4/G6/mSDci8L/eZJDYx
rUs90sbgcCrwFHQI5azTVwuZKk9QSckOImZR2aqw2cHQEZGmoU4EZ4IKWQbrJGksXcqljEKfaiJx
C1ebj3ARL4PjwsTHZuz6Dk+jcLIb3b31a0WjCiY7VV0xNT/im3bUokod7kh2PvH4hfkdqDWcAc75
HbJYz8I4CDQ6i4/feCsx3EPcUswH0DWHOXsbuR+ZwWdYpWGAmxWDUUNA/Ht9baZLVjM/NFwvxppE
Lh5da9Gd5AjRVuwIQNFwIsdm3mqVfECeWv8owOhOB+XPBV8Zo/yYJPTNQqtCj8JN7Tu95pCyMMbA
PFzpYYTvLdzG5Ga/7gJoxnDGj4JgGLobfSwBbUmatAZRzx7FR7zci2TMiLWjpAGcVxczS5sLmasd
XMNbgE2YdgwHVrZkZ3vPBFTbthxGa5IUsFBiBfAOiIfI54fB4eGVRw3PquTVB5tY1piqQhzmbTe/
AIL50ijOrcDVTaC76UoDUq98BDfXwPs/co6myPWOaGHJUQscS9gwpBKkkRXHW0AFv6MK5FXcoJDR
I1XWzWG9zyazrsqb3bUlLcQYdNCKSNex7apj5gWUn5P5Cq3N3ROvU9Blzw8pd6U65iv05yeYsQwt
UZFecH9mrN/kqu928p7eLf/iOFqifXwO78c2RMcSlT7UNL3EEQctPbgRUprFElztr2vYMA5qQktR
8Ko5h0ejQihPJg8b2Q0+Bx0vXJSBdFQm+m86W3F7nV5s7Jrode0uXAGaF76Vruf8zKoIiYdz4VuT
Xt93dkRjZndrOoyFow+dd0sDU+8qJjHI9aG5MRtrybXaHtbd90n1VYnPJEKgY5yK0OmnPRtFN7uo
rVkMOdjx2Euj7FlrP/yyzEsh/ETP/XAHB6POu9mYL8TKs2Dedc3J4xi6duDc6NwdKPdWyOv3WnrL
ltMT7lp70asT45lNM8rH5ZnPvCc/bY+aI2ALtJzVypNx02CDUkV7EXu3W1vBNRsXmWEFv5DP7MFG
vSrn87pZvT3g4iVg/YEZOgFmiB7cgWNpV1CpdqJaG1VmBkTrNJoUst+5H6FlPUddAqDyt9myyhuM
AxMFtnarvJp3KHYk1eFAumKQ3dSe75rt3C/4FUc4XWtSxBhuWufNZk1lqLTyeXj+jXvU30s3oYsx
fQGOeV6se0XInKezDmW5zi6iXKpTNfg9OHM0nqVAAbw+/tTU5pCvTK28TSt8SevQfiQzkkHciw5c
Zknd6gIx/KCDt4uD8KXzkge4cxfKfxmK8TpVEBFNRhxeQ9T7Nes9U5XKjwbGnaQXOeenZ5p/FwQs
o8LqvGXPK4VY46BkuDDM0sR44jGDW5xr9yoRMS8UBWYU8uCfZxmD6bXlo08CkxG9c7L0SpxTIH/J
qWjaLQaXic1ZKNvE/z7r9sgUfCQauHPqpWcVavwhQvBen71WF4dL3odltCvWn0esUuV4zJADsDEe
r3vsVOTHJhfaiHrPQgOAd3aYKmxmH6CBt7HHPLiXBzDlbgQJrROot+VXOL7Zn03B9rHs9PlNfo2I
nm9VIXbuecM8anABERCg1N17Kzwpxlab/lYCpBhgzaC4QTFhuwcip+7WJHRnOVS4RxkriRJh9SM2
hvKF7H+NBTYInW+KHmgqcM91XP/llHIyNlfcCM8JFvYsSJoIs6i9VQpalNgnMF/b+6iuXiKdWgCj
nVZkVUGSP26XIks74+ki25s3m1zIoLGfgJcYu35eDZGvERlyxxsVZG23+N4aciNDfeeOcY6qXKpT
Y158M4afsIzJbXOa5CbcqYyZlotdF1ffsxY6AMgoybyO6kOftidNq5uGNHr+ZKv+BcINQyhle615
UXH0VxoEx/wM9NQ6s/sfVdDZfBC1OR/XY9lIjGq24VHieXpNDJZgSYsIUUxs6wucMlg3hvcxCYrp
sKVfPNxOFjf2U7mHszuO1fZOKmLWwOBUAd4swlHkESXSlL5bs2MuqIvmVg6Y+7VTiFRNx76wVNoJ
xIhnPdWGUsuFVt2WXCThy10h1cm0Lxg2LeXcKBjyu3UXWzyvExXf3f5Q46Q13cEJ6NKfI3Otc7nA
P7FIyqNwSWxKuyGHDuLZ2NFva/srg2+6w4xYLMAAYtpYZzsOnfmhAJyxoyyYkFQl0scXGLhocxkB
2cAhilGBQAbA1npuqkjoFpX/u/BkzTOq7M38PkdpHjlxiJEW0DBhF62rvlPA+fHHQr1wti9Di6F0
7H+2UvmtcTlGNXQC4A/PWN4nRpH5/aosigZ5wdO3KR36J/f6Z8kRe54WLwKNtHpMwnWXx0HlX+f7
xpTolIOA9TyN6qgmBHS69iQ1ptVrct2dy1gOV+H/vjPMeUj/aGz+Bs7xEny9wZBTku4wdrbI1/DP
UsqP9/TZUuBWw+G4RZbESsahA23zumJMiFBuz85n2JCeyTFTb8xYhReUzmYQSqZibnlbFSKxKNvw
6hQiaCfIeCw6Us7KtOtHShqzFF0eIqcCDJv3UxBdAVCXMhDTrMJHXVK83Uhm4AA18lmh+ru8b/SP
MCPv31VVVcYhWuNGqqPgdDI60zVTFqOxzNGensMkpxkv1rjlBcpoK9S6xoTWpNpMaVI2Z9ef6c+d
quC/Tnb2xcB28pd5AjyPdCOzRGeGSE75b4KmkWlt1S2GBTNXB6NJ/XjXVZNJM1tbbu1gKYqsgRpb
RLGH3D4jLt246y1CI0CfhoYejCwjN9YPxcrOkf70bZacy2DGBco8dVlc5Y5jPltDkx5UgHXm3pOD
SHyY5TatPb/A4YI/FKAVNPpUGcouIsUU3L99BooF3p+LKdHoCG75yl3MTjitZUvGbbM5nKoxMnts
Sz9AI1KpPPC1MVhlCaaoThZUZ6cPZgJEFHcGtCIp6eJNiRg+NJ0KVOecFTfGgmBkk8KbvvRnf5kL
bTmceIDQ+4HNGpLiQZ/ac1H5qzREahsbcjC/qYhstnLpm5em3ur8v6Rm5mJthKINseA4S+FasQ4t
D1nghLcdLqGfzFFNJxkbY0eRg4Tex0xpI7Nf1U6q1VRBOGYRuB1QQSi4FapjzqB9DtgGN6rfyI8J
hEK22HH608E9QN8cUo3LK0WFl1jEVaxZKTykwRLPGkpJPb3Olh7mD1Ydk431NsmWKrqVHnxpu0IO
2cfK30r9uA0J4GZE2M0Ekl9eEKjwqnRrczGrhnWQUWIX2LjIT9aRDY1VMbU8iQDy8pAH6hIWGlXa
BxO+HQVDN2TqujbAxt6P6nSu7fwAB1fUAM59YNMGB9FllPFCQ22Jsvyu+ZhPnGTYDx51HWFWL4Rq
JUhFmTHvA1mLsIWf6PKWSc4YM6syT4hhMpMlcwu3WhFgHjAfNFYhTFQDWVv2hYJxKonpK5MRSQZf
6Qbt749yjh4mKJ1VzsIl1YzZgX2LMK7Jf5tH9fMioZOzz8wVPA4zKGHWKOyOzpc+10QpHyS6UACc
DYFok5ey8088dxIN0mwbR1HItID4DNlW5gTP7vAYoujx9yEmPKuxpGnEFF7R4M+c7epYYtd3vTQ2
xL8sl7PBZKPq
`protect end_protected

