

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hB1MkDF7gDUjtp9+r0pYANUYTDYvtQO1sWNXspOA3ppM8SYB929/qlOMzanhENZQcOQ3aiyEm3Wb
ozapXP+k8w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nob9JCRq6vcsk9H9VmyBE86hdNvS8BGq2p8Ka7dLN2J7EaHNc5IAaDkHipJixlCbGOjVeeUZyKme
HUzNgZTvjzVoRv6O00gQMvGJEhPJ3XxSJAOF+OM+ukp/m/tTtC3aiC1VdkFrdu6+fpapkZIb8cKo
kmCmWqIF3vlM9zcrSOg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qx+ritZx2pDvnekLOZeaFDvpDAtmg/hs096HU3U8xSeFyrj9v1CUwvI97hgO9fhp5hx7CLb4dRhp
iabDmveFs8T2afhIu9MmAO0ZqxUS0SV94sOYT5DwWoTjy8BTwRuP8Xrs/EEWKwKuWJp/Wjv7M9k+
wpkev7gSf92vj7uOWX6J6ECKwgIRjUGLc/NIrHrXqaq0yVd8j9fP6cvhVKR06OMq6U/6hMqO3Mwi
SQI1xdCXs2NXbTiCZKqVDbSBBvTJTo2cH6JXLB+E/g9NyF0e+z7oxCuyReCUVFJ21DVUfLxU3OhZ
gXG23tcqWGm/l3ZWHVqrETjEni8mwIO1yFoO4g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IXrSnaP8yioZkxR461AE2w19esRr4/fF4dA2RHFQL4fY5TpvMbkL+7RQBJ9eOLT5OFH1DsXcS+My
6KW+sTOsl2ndsfe3ttRCDI7Oeo8joeNZ8xJuwUGdOxtV0ae9PUAaVjkgDttLOomzNLph4uCXW202
bI3eFzZlGpn1iGIKiFQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iqW10+NxHcU1vbwMjaJKEOrgcrSi68eS0/IgZB3xPrIkkojO6+T2kz9ISwjr3CN6PcPo+hXCdZn3
Q3TnU/fMPFYF96Bkmhtr7AtYZE8GinVZHXJyKmm5x7dcsR8FyNv3nSOE/XYU/dyZhfnBj9H8LA1H
EJZm8T3/SQk6AB6tpXwh7kVAfE+bMsPCp98Fijzd/ynv1FX6O6GWv4CZpIVUKm7Fr8lIGCex7lCq
foNktfSIPTqF27RC3UxvVuy2VPf0Ck+rGl7pVu7l375TxqfmSlC5QxbXyTQ1NByeHr2LVJZwC+Xp
5uMCktl5vyr3uh4gEJyZSJlJ7E+uSrhstePVYg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37424)
`protect data_block
DhUqpdhWzQ9IZEqxhRV71ut8karxzeU4gbje4V6/L1ojKKXDMBqlGLd8VbWU+bKk5X5FfV1Ap7f8
+d1ClLSWKQkNZG0p+UwJg7ygOpq7JCha3aHipLQZY/B8BbMNZ/4vHRQ438zN5QzGvmQIJ+V5lopO
klXSuJuaRVFE59Fi29B9ZdYkRKzZR3lUm+8+hOxW1tJxZ01o2XoO8QmP5gJ6KUgzudVBVj7foLPn
aD/I/t8p6yaSY3ld0aVsypl9pDgGgmEsBa6PD9LxgwRwgQT6+2KM3NC4kYfPoPab5f9kXOKr1qnw
ZucYmu2OH2j7j+bidOYu3FRCd04+18zpvRMneGf3XyapdExrv4oKVh4769PhXoXgfrT/3Lwq0z0X
8psGz+0sWEw1wv3lMLRyvEglhJ6Nl2L2Yn0fD885TNBMKH92sR/nmLlEOZMdxn/MgXL9eY1eLuB5
HU+/oflvImFJXCy8Qo3BhNJHoced8vX7u8wZZoGIPk5iurZpje11MTi4UNXhZQIweZcBzHLjhC81
Br4FYbDjJUnVgYP0Kqc2YZgjLDKQC1JzHJAJKUEFrrB82k3/ZP6gP6jdbgtlyUacggjxPYc+wmvB
eU905gYOpnkj0jjUY6XFVDIp6Oj5IL4TnP8QJijwZqiOY3uQ6xD302LO30MarSuLFih7Fzk3vDdL
2YxNcJ5ayM4zZBsluawWqj12WfziObnK0vuWKL8EDNvJdExFN+7lwdpykpAN3+aE2kefjm0T2P0t
dx4zE+mPa95hiDW3HdbvdGE8RlAUHqNMrgHzjgmCgVVRQyRmrJv5foP3ofUMNB4MifX446g55yBi
tJUGjv+5rJrZvKKIr0dcCBnbvFwi77/IiSwT5kyDMKJipQPFG/2PNVqJ8tF9LZ3waahvMCPZAp7c
CH1sypWE+i9zh9DQpS0nAUpD1jib1wPvnPJiTaDIuZIrXumbHx5yd9H1dW8jiACY66akbnFNl2Kl
k97PL7OLU0OsnWZXvG1A4AZpCgRLka4JMjzZwxCwiRVCGgjDaeM8jI6nL9kE3HoydRkbCdb/gfBd
bsnOl08Qr0jccRzmYcBWoIn8uR0atkmy4AWhJdSVfrQL1uLe/WTzhnFcvt5/N4vamHoMRf1nwpqv
63AuNOhgDzcJ0VvJDi3rDxT+2jB3IycLJ4ew16XoK5QJLVmzxvv2/tLbg7WYtXkfUivNsdtpxkJn
vmMutDjuqzETZiP+Ecax6OxigIE6mqGC8wclgIJeF0FQtozbxA95RNF1uoImL3M9fv4twx+WDh9s
4GBa4bx1+UXXkhwuPn+HLINws8Z/owFbC00zD53gxiwNVgXXfXKANNHzB/IHTMBBDHCATxAhzXiB
6xkiEujLePYPv6uWBJ/1sBLY0LlNNHYduGg6IABNv3USu2w+uwbocJTvS6fFPQ50f5+yklS4tEyQ
35EtvSI+0gublsOJ5r9B1Y38nSj+9/TtKLCpiTlEMzU6Pr7t0HVMPYx9o+lwawcHn9PaXfQMo+kX
b08j7QH/eMBE/gL6uuEmW2IPsUZSEfK2DZI1/kwPnDM8xkNMqglFeEygCNvf3YcPtV9lLvDmo8y2
hWE0g04woziXtaMg/AouagFtyEXM2+Bc1P8cazW5SoWhRVPhmf7clMP3dli+DKFUvIFRLbxP23HU
fT3HOOAlwu6DzdwO3qq+FPpYN2pyNWejU6v3BPIayty6lMOHSt4nnLwUjVGS/EXd+Fz7z7SBF8jD
wVJVne2vgoqYIGu13KIyGCuX75fcQurL1mMdW2PvO0rzZkd8gAL79uLv7ytwdDsVXp8PzFbBWi3T
P6lQs13Eu0Xj0qIaXXIE/SAUbgGye7D4aXmIMEW36kxlHTghXD59b6U9PPrcghmW3UbwSYJms0P9
DFCsuYEsZxxcdQS52amQK+kmXu/AVu5brQ+YLFovsk2TTMgrdzrAHzqs5S4A4TRwmsowzCMF1bP0
rvJBbSQWkUQvIVM+bqADA68Vfrvzqm0i+0uroAtGC2DyN+qXfeLXs9erNLAkU/vZaT4n6ThMEU/m
sP95irjGjrPBl8IVH6YDihBwRKnV14ZfLTdgvFVwhBIDVzGr7o2xerI0rFqUMltaBJYBhHUOzryh
jmPj8DDcSbnJ1AFzoqd1oyqgXcNbtVETL5rPBFtwn/l83Ja1npLhoWC+dfGptD8ZwR8s5pG2bFsk
VEu9B0vuQgA7kFRiK7b8Hj0XjF3QnqbYb8o4b9RI+nRrQSSiSVZyqxL0kAqvegCynvHz/oRvjXAO
vbw9zN6UTm6RQuPaVRqj6y9ENib1D8twSkvQr9BxlhfwB8f+ZQwQwL+WY+CBzTiQwJ4daLeDh2YL
E+QmUMiHPgP2ywxtcGgLmoIb8Nqpeakes+2fKJguQb6G9DDKtjEu2yx34N9aZl7DYavKlE5VL4aH
WG/QeNk6VvcgS+C17id8V7KHA1Zw7BjYze7Hj0nbWQ3McGt4sS0V5E+4QVEpmV1fa2wGlkOOAJx2
CKGQqByhvrJz/H4GXUKWMJ+zYNlfxi0qclNEn7skU/sLkWWepa3QXzZzJsz+LC32P/xSWK81txwy
eOQEEwMpgKH1/PUcJeTlmttYCS94LS9M1f7Tl7jvQ9K14/kmpiZzBY1Al4X83fb+cZi37M7pbSpE
BaIexLLZvlw5Krawu9PazwL7UuFkaEFPsMbChAMFvJAeH64G9O9ErN8//UtQRE9tA0GvfQOeRYSs
eSx3kXEP/g3PFurcGqcpYt6WsQyLsFo/UcMVCzfJH68ahRl5TvGbqshWDYPR/ptUnWTXZjlkWHba
3GUSlM5Ck+dUUr93eRAGYS/ck3QcW/bY/FRMQqaZ0BS7+n7a4uErXo+KSDfU8spbn84BqeaJA4kT
Z5aJ1D55aLiTsuVXZZr+EWBl4+WARNDsWNp0AhUcGXVPCnaaWTM2oDGeQKBJ/yYhkf3u7i4i7Dvd
wclGj1BFYKsWzb33W87QkWV5PTh5wz5B5aTD9IkbXtnoqE+CBGMLMck9CDJArSdJZqIJB7fgjv+Q
VeK/NFyzh6bhU3MKun3BtlcOcctjFLSgoiEdzNMk63jGY82n8+epBak8oHjuwYP+IpG3Pa/zDOp0
GeWf/gpV41sj0+hrkxgH9f7aJgltkxpzh6d/L6DXClbTiPYk8Wqdf1QLaV5FJYOAVQv4hvv6vTJr
FEQV8rqxwiCFJBmFfHKVzHSg48mxsbMsXoN3w9W1rxVOOpRXTT2+HUNoK0Y7iV2CQ21HI5tU9iXy
7orN03bbGwIV546UdIRj67Ani1DQZ3vGTQCn2+qRriXQU+ZeTafCSklNKw99S6dpBaUdtBurYNhb
tQOBQSsORQJP72uvcSohUff+cb+afbYhbm5ifw7bvoWo7D4LL5qmQLRwTzEK5V9J0uk9Hh/3eSBl
HXkGmWEIZMRTDNsfN0HM5oU7H7GtXZ+Xk6IOZDYvdQd7BCwVm7RKeFl0/qufjmuDwDWIjwyZYG1E
4hRRhxsIXKKWvOYZTb9kzUG7UfN8C/Iwu71i/aY74MwoNBd0DK2z5uK2JEOmArGNsrammBeTB1sq
YGLHWh5xMImTdz4W79tE3VnzCS5Ws3Y7h8m04hI+KO+eBC+UHD6YrdrD7DkdzFbmVS4tfFUnFfZT
sbpMg6IhdHB9Em+63D25LB/ZOXHbWRjyW8QgoXfCd5xYtQraKZH5BZShdli85BEKhctncUhU2gcE
LT93P26hp5ntFKSeQAiHcQ9f4LQ8dP09RycwuPCWMdZ6YWp60ggkVTQjR3ijSpzc0ALF6kcaE/ps
Rj3KGV3mWppkvRKENfU23FRdPRUNbGGWSpAffpBJqDTD8uHEFVjoxLKIRBotZSJgiEMalzMe5fLg
EgQuX+ErNaoJ+WPXZwoHScnY8ImVyarVOU1OkdPlxtUFtnXqkBwGCx2gdlbBY54i/gyRUt7+sP5z
VGq9dXrUQveYFlWQHDOyaiDy6CAw6yOCzuWDgGyNQmWwN7ZcUiHb9d8E3/CklowhyGRfD8umHT9F
Jy0x+PuM1MRIdTwQA535v8UcRxbtco8qsIO1vsrVsMBYknsnoVf6gfYInBb+u4Y5fRaXSYaH88RY
FAYAqlLoEjR4OHh73uLxZqeAlGKkXoBIR7ZQGpnflcNuxMrUpWXztfvIKbpmZp9MkqeKw1jMFulC
HWjahTxbti1ZgEt2VVK7CkuW5EJ4DXxB3qNkx06UezsGuvkBRgqSu8sr/QCNrfHHXOtJfsHBxU45
jOL8DV7J+z94X0WznkdzUSdzHWm36X6E43D7+u4CrS5er5JFAy0HWIC+1Rx5+FqlOPCn6GlyHCLG
j09OLY5CNhBxhbFl/BOX95z6waLbabiuybtNiMRUMe0Gx90dgBaBwO9muGHDGFoQ7ab7tghRZxee
JxtzWY/lUQojgl0PPrkwflEBvX571piPUpD+x/Jasg6p1wzOkMN5l8QrVJ1Rnykxb/rs961tRA/1
F6CPidsCx55imLi8sNvy0wxG/6/ycmfocsF7J31bSJiGxIkIP6FTJYIdbCuCTgSWsbA200xlK8J4
22iqzdR4SpdcKfFP0OpTJlGWsYt5C/rqzDPfmQvLTYs/CLDAtJnF8I8SOo7hsUGu7jino6Ud31QS
KaXSENFKPz7SVVt2qHQcI2EbnIj6ww7pYRi9U+0u5GKZ4YEOl5TaDq2ysDn5OpAcn1A3Iw76by4+
yYLDc9AFTR13bVZtpNvXJQwWYKFc2Cjp/XAzMUGAJ+qQZWhuibbQeEQRYBGPdmwqYdZlusx2VKr1
0JsHUdbjvJVbOSEx3UV7V8jG+g1V9DUb4Ikpzlpvn3y8C+RvlrKLKqEffXB2Op0HaNrWdC5Vgng6
AwVv/ylVBOq7RP34Ov3IZhZCBU1kApP2Jp+ht3whmyvj4s4T6/QG6movik1kPcwSSDRnU7MxKBrK
NFGXmdT4iykRze0sqcct2Uzm71da/ZUsJwujL4p49Huw8KlS2QoEZJZvOOsMbpTu9Q5i09fywMcW
9eMtgc+xxd6mPV+b8zsc95VkaZ6HKi75NJLQYCqTAHCLZX5H08Ix0yt1jPCYOKwIadCv374u+gFi
pBp3GkAv7PZks5gwKos9ri/pMyt/EqmG+enauafvVgvdEy78FA8fQ7mj8fWY8AyaVWU7fncp64IE
GjzI/yW/9kItmMSZv6EnhEBL6cMNRWs/6vaE5swmvCJdNm0hAoc28gFmNTTNTrbM8zucnN0cV/b3
UoTOyrsGXTZAusAwHjTf6KQjFPFUvqbBp2Dzevi2lK8bjcl4JQPlj1NAsPkbj1vMJ4dXocpXi4XP
zwnDCNMpjJRWv+Z/K3HBRJZ8xF6QzDI7raLO3ePRXsLQPM40cwk/Sn/CteugOy0u4MofhF+gom+L
jIrSkkgUWa5ZYWKnSW7EapgynD4Td6VChGAM0HRgtbkP2n3gX7LW2NL912qfgTCbpbn9TQLujzo3
Z5vnAS4lAeGM6zHIM7Sc2yLM669LhJ2/M2mU066bAGa/VTj0J42rV2yDjvMawRISk191jsXl8UEw
JUnquebdtfnTli9/7635Vujm9fqfb0XCDYy7ZNu9A5XJoP51yXbW0vVzoZavILSe1YBw3aq2ggZU
NT3b0aWWO3HIEezxBFBx7HJdDjTHfOcJet2hG3VMBzPLe+itkpFa0pZ5b4f6uKWapttTGXjjeSrC
fLZOhwvYMD8HjcGYplWVF553pGjGu9XAlwe8skDNj+bLwOVvKvM7EBmBJ3zMwM6BDmQKkD1CM+g9
2MZsSLXFsjX4a3uqEB6AwW215Ly4PKb/np/gvNSyRi+n2L4YWlPN2aIfkM13p33MdmXIFV3iUDvs
q7y5T28Z1wbWdmFgnm0YWZx+Epcc9u1Rh+6XINIjD1J69fnP3YD8DTnUFZLwXtb+XB75V1Q/RB/l
L86AC2GQcussB1cpr8ZYRt9zX8Zn5YhvgJyBj6pxGyRkSa+SuJqcA2933zwNNYJY041JUUX5pY56
3enfSLmNrLeVDvn7m33QGMQAcc1bYZ+/r2JPOssGRbIk3KJCNe/tz3RPbtgANtgrRkw0bufj5Guj
ayvA97Z+pONvee7vbXS2AfGcO9lzGuEgB4uXX8aK/QwNmKTKXNjJ9dv/cOPiJ3a6qa54dBBNo0hZ
jxOfYWyxhmc2Mh5AY2NZBMwCeO9tRlvJyc19XfoEvrlC57eVuS0Zo/r6XTWcAl5rd4eqH44CyL/P
/uVB5Lv4+ofTqLdvBD4DZArD3gpOlBdyoq9J9Ylc/lLxECGFfav5HGTnq43vZ/f/0MPQspOFQWpV
A2QG10TDkpUvnzOopHo+PhJH7zRHUHzkkgg+EJxl5h0j8SSvbsstnNrzJLqEKwcXIOV+7uiOrlTT
pZ3Om+B0KR6SB55b3V+1h7J7pZW9mdkpfT0NKQd80pBEEqfMax8396BszGORw+y7/ELZFn0PQTj8
3HyM0Fbq8DX27qC+cPdji9ZC/zqS+zT5EUbAXbOJBOm7ZXR2nihnuz4oU4wmLpEz3UMN1+l0MAme
ChvhERmGIgfqnrGvLGpWISYs7JOpGr/JCXBgtc3+4g6gXhmjCkzLhNJuCajXjIpjfMKW4sHIt3j3
4GjPtIP5msqmX7988z1QKfIJF7pxYFZCKnao6ldhmUPn/GqzY/ejOm2nhRa5ReEPaelQhtEXHfZ9
v9+gyASjzt7KW8fXE7K9G3Tp0I2z6IfB5VbOF7RXBivg1YHlBrbX9LV3zawv2XT1hlsmaeKzc24o
PMRjMaUz2mRgF8OmDg08oddipkLPs2G/6EZ40zn7qnr32HJHykuBoG2/JKJnLBF5OVjI4dlwAstu
B8BX98M0gdmz0/qnONOU1ivTlXWgW4qU+FnwUEXL++yKlzr+S5UrYZV3LUvzbXf+/lplL/qKAZOc
3CWo6NP9tKt+G3XHK/PW/3R3UtANGAileH0pIqAFLG5UGEW3ZChsbo15NXFm+SyWJL5IYBcSCttm
zwLOSIc2TD07nrfTgaYayPnx2JZXSY8Ps+44vYm2zL0BoSCREPT2EETHaNU9MjLalCCXIbFZyadK
XHq4es2FdmGThT8Jydm7zZUWrlHeeDJhSUd8AavafjSCG7QZOvAtFTba7SO8XkNbn1syuzxToCcq
B0c0xRNswtJoukXYCBSGXfexiaRpHlB7zJOiLMHA/huxtRhoz+4fb1hxheCsqDnrSPgv4vVsh+Y+
QouCLmjFIe7jJ7X9z6zl44diV6hyaJEg07SrPHcyPcVTRbAAKwDICKdTAWGc3wwG0RuDEPVfn0ce
yj41VBMHMLOOZNcz6TZprb8217wRmmXBjFOAujSvXPhlRurPtwnZMryNDryZWDTWlMgH5UK6hBst
MkRSNcZUKR5o6vw8EJ30S7MUM/O1yJl1AHnY75hEmdy5TTq7iF7U6VvTjalTCE/nZVovtKSELF+S
uUMIYRa/uc0YOd8QFERbSkcmOZOtFJ+KxhIr5QzuNXqf+5rTFJBjLtycfl2fk8MtO8VC7PwWBg8u
T+r69a2GVmSbqUvUjyBE+r3oXIL7U35knmDEj4QAY2Scuapir4gq/YVm5JVGRVIMh/s1zXFtVcyu
euIOf+0dxQDqYza8LlvElUYOp6iOdgDBP8e6IKaXilFGKBFQ4ik/jtrNTYN8scsUl7UMBNuS8nDu
d1aho8HXH0RGbiXAOyeRi+nI+kEfhQxWLpRWY+KPLa2Xz2GxexPQXfGAKuAWR9Q+WEemezNqG3/y
XchA5euPRhH4djwa7Dp7WKL715C8MZ+iO4R/HGUNN2RB8if3x1yOrJXXpECfVumsvKySUVO2GKQx
8EIRqFmS3xat6JtK0jKApZgwK4DxX2cKNLOx58HItVQY7UqZoP55I05RwoxpmOB2RjG+NlnRJnC2
0yzt9rzLCRiBjUlVwrBavkQKUaOPoTetF6RYg5gBnOcsTFR8nWLBqJDO0RWpc7u0g+7mGeCMeCiw
70cMfo8hZ70XmQlmNVolChNEkgycE8RxHOfHQDPdzi8JXGRlwHT243zN6hW8kHVao4CS9GJiwbAM
8XwmLitqQYHpUBmdGQ7pHtf6RegYs3dWWO7ZAtjzYB221ffMA+3SWQsAgX/45CzZOoloXc0Nm2x0
UbTCBPu2iuc2AfPgw7+4ULft7Wve9IayEMPMJw1v9q9QdfYV88+Ib9whVFi6yopjehAhIcG8zInM
oBO9PTyDhlA38Qj+6rih5f19PPDA+fNH0cKC6TAy/v9JpyPgwvcLm5XGH2CbwvpbVLwaOZnZp1WC
m1OWD4uMyEC0yL1ii57KuDZIQapASiY8/+NvxsKC22/UMJwPIODcXMlToQnEyhQypsJFCEr/zJ7D
nwqaXuPFE6VpiFLBu5hJyUQFZJKbyBAeaxAA1ixLXu9aAWIXzv2QKA11nG10Tk5bctbgWl+mDrNV
1cajnoHeQrjevtYqSUhV0dc4mBcTMOraghVCiVAmk3Nh8BZEJA8b0l9QFxPa6L2FAQ/R01cPw95i
MYbn4BLq2EetBHazUrASzJKhsQ5d+RO7C8wEtv1m2M8RZ2rKfXk4gxuxp9tYfsIn7R7kBj4+MLYw
IzxEtqu/cLtxQkPABz+BCyAsscqO7edcKzRsy2WwBc3DCJiqaF2nzkwfRvDQa1PNcb7O+JPNu69C
J4Zisuy53M9cXujnMroJ7gez3OMyRBdkS/EbftG87z+eHO1V0UrSAg2wRvb36xqpfgHu/ho9yH5d
ow3Ult7dR4XqNNsNnHuVpOy6f/6KIbr+27X9xboCf/9SAvv6N8dZX5VdNID9nUoUT49cmJs20NbL
GwCpwSKNQTABdSjxDOnuK01evw2M82JLfd/tllPlQ9GeZJ0QGXG29qC6b87FW/9jkBNlfm+MzW6n
762eQHrk+Aajh/tF59WLzK2IVHD/Da1E2xqIdlEUB4hr2RFFKx0iqfHQpHcD1TjKZCt2jnmRhX18
e1lj65ypD8AWThBH5noT59+IC7vaV5hww2mSiC0tkz9ZayuNrU4kRCdCIGQM9PgrAeEsSttV82g5
wytyQm4LbD50B6RCaax1YgwJXuCTl1KfyRWgAfDQ7s2HuJKrSyB+n42602b3pLsc/CnYzwqOqC9N
tOfKUTxdBfpAMu7Y0HO+s1++hyBvE2i78/4z4kVvFqhyvVutn2EhXc14ykgz4Qa9c1D42/1McI3G
g4LLgnSF31LU9igOT+obSZ7yrb5mLHxqzuLywfZDZPK20W3nWaq7s8r3BW8Ao74AzM3UW6rhw/Z8
heH5Mszz8XjUEaQRMx5w+m+hfP4Rwi6TtlOf3oapeWmBmwo7DWjYQEcFTJ+yWCTVnGcLY/5YWLlV
5YGKT4fubWNst/KKxWRjhCQ7zK+55q7tTT0dUvDGdEgP1HKHmMrfYxA5hs7/HVjkkdWy04P2iUZj
v6NFJZH/FfOLFrL9qDb7fuNEEq9MmGPd/pPfK/MUCGIStC0nzbf0IAvq8eg6bD0Hp82m2aqorQaK
4MU+wdO2jbXidF1tOk/3L8D+tplcdUsW4nMlRs5fT7Kv6AfnBOngzWPTlj2Kx06PnJ0w+sbukRXb
M7QbLz0g/F3vxXRm6roVWgXpyKAZQw19/QVBzhWXYe7vzvdPGXbJvXQVrcPsDY5L+inY6SVWaLP+
3jwNzFe4WmaupCBiguR11iS1a97EDIDf4uujQweALL3K6LAOnN8uEFaidkskxAJUHdYcc+a70stx
zSCC5af9wDSKUNOXW5jJguul52vT31JK+ybbvE80+9Wt2vExNukoOeg0uZY6PE182Ts9vEPUre2a
QUSBLGq9EtkLjigUQi/QGjaz/TgeC93JkU1wj3szUPeo/7kh3/wzCi6GJ8W9dqZQui8xoGmholHu
4kAOpcm2SLFmDCxZXhzfiG6wpWhhT+Nqlh4/lW8LbRDaIdpQLmtftZuqyuf1L2b2nrDRoVcgU0nk
/lQtyfTE3DSjFbCFRWeuD4n1heOHfk4OEjHG8hOefTZuZKvMtCzhoHIGOE7gvFtfUClvlCb6QeDg
f2HDIk51v/5bXM32B+h1MsZxV+ZblIryHwGYtKrUH9bcUCGEeKXxat6dPKwN9J+dSXSAksiEgQri
faDjEnrrgxHAlnk2edLAip5qNAvQ/tex5tg6oR0wB1KmneE54sgrep5cAPcdiKV/rPwqlJU86A/p
dWVL0QMXSTgzATiy/oV04gFjgQW/tsyCjy6fARnMxR8ALce8kUalQivovEBoHcdcx0Ch7lPuyccj
jI81uQrQBrE/62tvmsW3W8S5AF21xv55Z/bzog+xN/XitxAt1F8fs27YQrCLZkkI+r0IpPHAQdl8
gwrbbYdJNs2IkNXmZVGfgBufxFU6ORWsnt5q9/ePChNU9hcd5xs/lb84BPSvG2bKR2466BRPjtTR
i1WV8KUFjAEjQTMqZIUrRKrZQDWemGB+pxafWajx2vtfQT7kJcGHKx5bYPV7QRlmpcSbwZiHHzf4
gi/nYGjUnHEEM3L3QKJWDJJwB/MBLAq9CEsfm7zKkkgdQqLvj+jdaYOxcO5mrCicdmZQHsNg+iHP
mM7bS3+8KGsbSLgpAYVO174EMxX8mLI+XykFFbOuznn5WBuKGzKBcfaISXZeu6TrrnQKdH456+h9
Ava15s/9MI9zfO079WMNg7kEPm4BtITlP9MtRcd570ovT0I9bJm2rEZocZ49bBfZhP2eDQ7v7iIs
3CiiAmS93ke2Urt8aNw0Ks4Twr1YIn/lOSqs0PKt3sTqE7zIylW8S1NnBrIgV/x5zzn+xrHNrW/u
+a4ewEWFNHoR7x6Qhc2yDDvkrKScQqMaYjlfnSmoiNi/SuG9Vp1K9NIHNZoC2v+uUc8DTHj0XuJr
xInHB7/MOuUuK0VXvc49iQThDYDbAsZyzbM/WJNvyT/o7xLc7yikkyljYJb28uYhkYN6jAMgFICx
3WQXJwGKSY4tYWAroGn7XdnJkWkSDDUwsdCRMxfMOj3oZ/SUQMZTuXSWMK6saFxRDGldKtzy4BQc
EBhFv49RHKGL8Nzmbsm34+M70R6smANJ4eVcckWdtKvYduumnFrqMHsl1kNRE0sz9XgODqOupNAr
uc4y5fms/2S3q53e8kEB7a3ARSDyuZMo3lPlMwVqQpBSP5HD2y1NKlTKD6nLti2a0BOXkSfWuHUS
uvY9/28kEeB6MDEqC5THfyQPabPWJgH+tZEH9jD91DbR4FJaIYW8c0y+D7I+jPEWlSgKin81IMMl
s2O+pi+9x4DCKxUObm06LNWaX8lk5v7UuYDwMugN2QNggjKLZI7kj9sW0mJbdc41O2/ezG33zN/J
XEwp2UKjc1ClQ3AbrpDqcAF2mq7kun2l6L5infJpQ7ENedEMSchcovJGhFnsqGC74M6l5rL77jRj
TvHFA4NMA6r6x4qd33Ge8DE9ekGxEpT2jg+Zpo6FzkoyjfoKkWonQQ3a2sPez17V+4jxeae2nJ++
t7l3hPo3axW+4NOAr5RZ1drtN3MRoZMoignbhsm39pGUJQJOFPCXcyo1x73Hq/UNHMVBi3644Ccq
lysLTsqPSs+y6HOIEcaQJprA4h/Cyvsi2SDY9vbgpdNMKRluSLyblClYL/q8NyJtM5nLxeNa7aU5
HrrDQ9Oo0Yul2oSfxj2o7YyEFiG4giVxS4mERz3YiyQfLAKnVzoAUSbJCoc4AtMFjWHYgCa+3va1
vMKFgbwZ7h6YMLGttb7e6q9tKHkHh/1z33zveirLKYSsnW/36bppYmxbhcSrPQYWQcDfu5em/o/L
ykZCqKRMF2gx0yDXXQwgBxONJdyBRZ3iP3lioL0i/gYGqX8rKtjXu/ggU4k445s/DeQgJb48wsil
eD6et1vSUnFRZRHU5q4D2nlilAyGwjmB4BYSF4nmiO1HYcm1AOHvJkR2AuJ/3kuzBYVyoASZTsud
JLQnup24a0KHj0G5kja/UxnAk5KLRwAHcJffXer7yh4piT0GZsZzSFu+Ug6SZSE/dXxvL31UgK6L
nUetdXS3wYN/k6If7g2lKGXpPkztKe9Y0JsxOLSh2UYKcCTFpaUyAT6yGZqS5YHmKjjZJHcmllOl
OAMYiBR+b0q1TLolkeFY59L3VIZybq3XZPFqQ6ZqTVTKMLeZ40ZZ0UMsTfDHWpZy9LqlQRrEEq7E
OG1xTFw76NYKPLPa6pqtothIEEfikhK6+Quy2C6067/NAkn16Twgehv9U+rmZDY2SvGc6we543MZ
A4ubsHPXyEtUhdTrWELs0SGFSbRenTkhkCcMLc2hEbOo5sufe1/1Of8h9D02EyO0AoSVqev3HEbc
Nulp929BascbVDW46bBg1FkwDRbosbzfpzSmY+HKBhe8eNBNJcQv5pqD/hvmNFU1Ptm+HNLnotgh
d4WNDHmOb2OJTEI6mRXUsfTBg6Ihs/S6cO2R+mui8TI3wv/TzlphfbRpPoOWHYQ8LCBt0wloxZeR
S5HSF0+oBqLXlhX1LppBClgm6Y3jZvsyABp22bD0m5lpRT0cP17QCjW0/bRJV6nsAKKfzfikRDZ4
zvLPDAYL4/RKpvnhLw2efu3Bp1KH57Xmx5MM8fwmR8LolRQOiGW1UHd0zps6c0Zi3XaCMs39mXH0
kiIQ8bJeCHo4VvBWowfhH2QNp9Tbx4XTTIiP5EWWqOAjXTzooJULWaZrH/VHE+K8omHYfZa8xYuM
8G36YWTFNsUTMu44niP/CwG9+YPtso4HwKG6R1hUoVzibbJWq+VHEROxoQhgXrhbzO/k7kn70pfL
YMa3fPDiOCKDyxotpFIKjDzYmwhNz5yv63u4sNjPjhKkHb6qVFpzuQ2JRWSgDfGcOt9a/cnI7oHc
wy1E1tr91XiyJOp4+jZfqeSlY0vPBgAnselFh562Zh/Qjq3pkrK0QqEX8yTWVodz9IC/OyFbF70Z
xUdHKMbO3G8sRGoVfON1h/rNz0MdM+Nq5mET3NsFviOZr57BSddya9tZ9EhRERJ75Jc8NmT++Fq3
Z7dYTlpLfHycuoxE/1mQzrTMy/S59SK3qGTaZ5xaBMQ+PbhQb/j/USsprHujdbVO88OavFS/Jkmd
kLQv7xb6Blwq98N/qX0iWpHWHzYAp1YV81762t3jU29NcF1z71U2bdDOyy0CX8An8SVPHg/u8E3z
OboBJ5EpRQ2+1xIrvfjGZ+M73NNbuL46c5INg1A5eO9w8jJI9fU6pEeMKHZaxhv1dBAkoh8Dh7k8
rDO4T6cScRc0ux51OLTXOKsqDAmFOKRrPCMJJMSslUe1jHG4DPjix2+J/bA2hc25Zye4pVFJH0BI
hPxGA6Un4KYutxVT5x2foF6wOtdTmUdoY4d3F0xVLLaC23n1yS1MVLY4UadVDY7kw/G+2X7vo7XW
J2MRUtp/DxA4V/qlxJiHlTByRbCSzlVQGSkAnu87TWi55ua4He4P3M7hAGejDkqpod9AGf4+N6WA
1wRTY2+//ZYN5Ped7EJ04mhtaX4Bg9HLL4Oc6MH6u0FqbWEh6VlpCpFI9KNKWVt+ffDISwtqYEPk
snvHxSv+bYW7ua34zbRZFg+E+nsfsMHHKI2VicBJb/PaClf9uL5706JiIM7exltT4TmxJcnOaCSn
rBN4tcZw15it9wZLsqypHP52PUPFmqe5lxoD2yLC49DSB95pBEyAhIqIRB9IqLbI9fz/z7COBzzX
gIFuRNF4hBbKTFOTdMahH8NJXejBIf7o9x5zOt80Fqezo687EObMUiCRJomd1bjEYY1oSLvKlYPK
+PrYetnuarfi+hVcqc9wf2XM7bP3SGS5EK+E7E9tM/gdJUVckVYK287FdXZSy+ZfcjNsaMTBTYkB
zqTcMX775soC/fdmk8jkTXAB1Od08fY1ZYcHulQf14tjDVAhAObA/GqMy0Hsy3dfkz6v3zTlATdq
XOW9HyazzVHw2SGVgN+PXLloqBwclAwMKKuqasg2dJhBr7FyyhUJZ6BndqphCuEV1erZoC5GvS/X
CplLn7sWX8vPvwGCuhd5BJpoKjInm+57CoADgaJ6hu26irC4Q6WjPh1wdoGKthGra/fklnnYOeJj
uBx6dP/DCvf6y45N7Hz9FkrxgE7DSFK+DzmvueDv2ONGxdZO7PiQ6KChYNUnAnZF3CCH6h16WD36
De+hT4TilZhbyDsbLL8wFMUywjZiQ3GAfl+c6Fil8F95yPhAKSJFHyWHM0qd9JYBocAqbVVGyP5M
IrgjzSmTg4Y76IENEsCYaJTlqOsy4ZYyEyNMryfVpYNa2SwglxBczbgyw7XK1QbmjRpJBVrX/pnc
k8uOM+Qwdo+kljbZaEnPjhv11Ydqe0oq7tTU45xxBix6ixyHN9raGe2CHmv18wBKbXmOUbqDbito
UhP9PV8d/fot+NvLdvdREsZqNgE32QazNanfmR6ii67P35qPcXnRLbUZu//qR0/uI1Dc18AjgJPe
CdGiZAPqjEwec/eJ1tckMX/4qNNBMsoi4PcH+Py//sdWZIR/vElEJ/WgEM4QlF06gdh3Z/1J7jJo
GHosIls8/kB0/lCPpSE82pkGLjI4i4e+ci2IVL5/z6zZ/oj1a0hlFb2Md7z3QAL4yWr+ZFItn6or
GbnZ5b6zDMEiMuxTRQ4aNMLcxNpTcpeh/pjBVTAkDi4ziZ/G2PjI8UrZOT1qYrhGHzfW1Hg2CRWb
Z6UN2ZIa2XRuYkhWBNQhOuA31ufJmDhzPy5u6J2JVRxbMFgKTxCaNVHk4+0C8TEH3+7Ob870ffQ0
s2E1EtLLi8hL40VS+872qt5pYMVmEpoI2id22LzoIgRf1XOZkLyvGILdcL6J5UoXx6MnUzQ14lGk
PKyN5mBrriZoGVfinvr3nGnynnzMhq3uNEazEGKnaAAQRJJNRt9StIo2BJgAQTQ6YGLh1E/lmAZR
FThnK6CbuvoOVszQvoYyQV+wc7bW2BafBwJeInE3rjTjvZxUxlYYnzMWJgpG3PKbWVV7nIET0s2c
abEAVCjg7yZz5exXIaGcWGFnoDsqA1abhiyxfY/AEQ2q9wGAa5//9XoTTOHyyVgCSCVywzCWp2RN
SHea/Cc4lDPRdgwI1BhN7/TWGcSx2dtsDNvXUNrTft140LUVgI0pwhnVhhcHBsF5G1Lv4Br8MT9L
o7TkSCkfTLPHZ8DZfbT7M5gfUhCDAtt1nOwwcIqy/U030LOv5g0QDkvfNrFd2NwOtVnn9ccZr2XJ
TJDnVwcvXfk8+PVLb6qiA3mG1DdkMNpMFhIrJXRUm8cxuWxrfe9HBDhyxHjnwbjxdnvT+cGR0x0l
k77sBN/PsrVW0yolYrdYa4rK4kF5zu2CSb6I9LM+3Zo1xB/39boq+mXd5VZGwo9MyteWF0JS64XE
FOO6T7dt6wYgEl0ZemBepkUwp6W1SoFhM/VUzOEbphDhbhBJ5EL6VxxAUhOoF9ASvnAxlQLmijAY
774yDlrPyNSI4jatCEP7MqrnUKQtSQ4wsKpzkBW0MMuWpzc29KDhmVOA2xIIKss94aoCNWQzTZ5g
42iDIfNaKAU173JUc0bchVZbViuDKe5g7fTvsqoHERJI+YCiaF2gUjg0kKsV0sOrzK4PgD7ahRxy
kFxlpPZyjn4eYQC7QO8keO3PvA5CFCaF9jfw9AAoXaYFGhaQBnh5hG4AAsLivgrsso/P8AlS82Pm
jOeQBXw8Ti2WJoH/eb7r88jf8eKFRdouVr96w4yWocMGMc3S57OiRhrSwDA3aaKLJHLm4FhW+5y9
5pZB6vF2noADh5KKzdxDddlzXUSH5fRv9Bdo0AdzxLiRQIBWFSuS5RnumQ/i17EGrvlIPxX+1rH8
LiEYQQc4OUk9Tz8R4cAVMcbOqlsrD+9Y0bdxKP4zT8ItNgIOPRNHi1OuNcF5b0hSqRxuGZ/lMCB5
9rr+Zada9J1LWMQwauUFGnXHYLCHuHuqonfkQdLglAmvxzYKESX79MKlOh7Q6nkJt8ENtNpS3LDu
+cyJ5tctFMa1XcEtgXDCUk7OLPb3C4veHs8JlTUusXd4lm5YuGEGTNrqRwryZwHE8P4QywC3+hPY
Y4BaXurt4NuaUDS8qPKSKBcRxOPZ8reBHVVgsJdViotNcaq8cfwqFBElP+/PGoIFIYM29p/8m2X0
Yh7qr/5HAw/wd0ItF09ususIYFRQEJHIId0uocfFEsDWoYM4HxIUgjCauMfy8s/iaxpXV9j0jX0n
peSwNBMLQKHf2HlDgUHBazwZSfjhF67XKRrZcCV/1dlDqmJsUmpJNja4hQLAaHL5ylJ0Aw6UAmEU
2VM6pIkZswurzDYAgamqlcIgiFokGGw7dQXyJGL/NZNQgQUzEFE9ULn4XR0ElARxRWfyza7ALJAq
524zq00BBm5MUkeZOmrNek9y4x+fvhNZuTmvPcSHawG1Fzoe21x8jtMB9ojj/RMOtKJ/2TzFUUvN
TVsgZEvw/MBg00e1fJyr/Q48AbtmDX2ihze3HxbgCs6XOzAqnTHhPKOsiiGT1WXrpEIM/jhoqmSC
PlqlqnqaoFNwtJ+etF+dRHVQLlV7L7+u1nkOzLjFEF4SfRvYkbACLRwEl+MV+3/PzI7oSZ7DCvUo
Eq6pT/qXJCY75VZRbudZwF/J5XMOg2mug5TQc5vGgJazkhs+fKP2W4WY2f2+bNyrHyVBCDQ29Sve
F9NLOmv8XCmV4Kq9MRX3nrSvKpMMWAp3cuo77chJo6lZi1phqDAJpmSa362mKYeFxhL62XeQSXt5
mJFNSbsDAf/vrtr+lPLaCYl9XZXegasqeM4L9fYQp3tjNcxY4NY3ymwTfPec/J9sCAifc8uTyabq
wPJ+Au1pfyS2r0Z2TWYtq5BgkLaEflAKUU1zU8dYGEmjQrq+Aop+GV0oWG7M3OYflChS52SuXN51
IwXfdJWoqatsmVaev7glQdlqguan+0U9vKIFpRFSFovwIRWqafcHeBCKS3L3sUUH19B9RtN4WJWO
YQtVtuqbrshXWZ/ovo3htm1sXWCBOLPGWOUN8xuJfddF1tLMLIPu23N84RhUyG5HI/8VmnNOw5tR
rkw4TuYmq0JikrbAXWaXoDe+Luzm2R+zN5zP8su3u55emykEygbcsOhR7sOEMpkuVDBk5CPOsWwD
idOf2NGnD82WQyDa1ZiSfeS7m2zHe3UtxCRDjrgMKD3pcs7l/3E6Lr0F9Uf5LVwGlcKEpTkSwvnv
Nk1DH8Ca/aEnvpMPSBxKKEKcBRiQP3o0zW5Rx8EaXN7+3CeVTlaxrwnHMam21QofB1XC5w0CiW+T
eoQ+tI7nD426871tFlxAJTdsZhZay1iAWzUhibxWHnZHj9lvQCyURYqc+pzihazPVoaYWT+CJNAi
Ii+tFlJxMvMFsjJtz9fwnGxcBvy6L5F790X0DH6v4rFB5MX9pz4PmFsiKnClBwirGaDqU89Ooh9b
ruP3Wu+woWZNLRgPjM9Jy8ArT5B01PDD3026AFJktmY17ZrLdkY7itHYb4tHssPVQoDjE8X4JyIl
JgvA4p9yBxz/xchi6HI+nnS0Ss8EAdt2HFa8tQJLJmvFTx0hHetWB7mFLTeLt+iPrOEOWxaJcTO1
TRMmUoTJv641PC/JGkh9wRbozmTxAXZB4cMwlzqAwWAb6nZVhSs3FfEy/r3+xHQSPHZfDR3omm2/
9SsfAj4KuO+R4fy0sY4/4vByzHhC+XM2YscQuW/hYOT5B3Wa4sa0goCpHveghDXwv8VMPFlNHIz0
GwxglqY3G3RkHcSTqafqjOldcCv4nRdtQhMY/7fZCwMPV/t/UAS7zn4/ZehoCpHBdWsJ+4qy/XVf
0yHMPpLOk9NHRPjhsTt21ouPeHyPn11ETb3azjztFSnTGKj2lzZ0eFnze1BXETUyQB7TKb09yVB1
a8NEB/y5vTj9q72//OgpCo79/KVfzqLnKXKDZMZF25CkQ3i1/f4kZMjnk5yeu7Kku838K3EbfsNc
r2wQllqp2rxdL60R88uia49JzEuKnuM4K2VMGEROUBVRhKghGa7PEMgbIROaOyFPmJp3pYJt6tY7
9tpiVtL2wO61F+Jc03ITU+lb3ckp8e/oUAl0Qb9QOqwf6Y5tWT2Z8/C1SJ8QW0GZ4opzTUP5gdpJ
oGzhupgTSI+JRrm1LRhGqGsJfWiGRS074qjhBBihg5+ZOHkWRPQdpP28afyF6DWE1HaxBrUt0GPl
Hp48dgblTzkJIrHIKUGzA17DYff00PPQm/dA4+0gQPFmq2utLAeOe7vtYMUreNKLFml5rEd5vR2n
dtPNDmv3q9/NPZKUQ5tLw+jUoIMG6gbrVDJ3+xK+R2KD+ABCLIF8U5aRi920stPlVMG05K7BG9u/
eOCkXWlGbdrCso/aD40RMqAA3A0+V23MC3pqWhzGv5woqRfcNMALsMYpAO1jv0xRPyE2HddxaWEM
HH86R2AlsRvwWunh7XugT4n/BMbYzdwoIC99bVjYC9MH8BxPZkR9vsXGOmcOYZUDPxPFe7CONB0T
WSUoKuOMTkNrm4bYintHjfzAWs7PnKQdv8ZXGlXu/rhd7NZA7zKepmvx4uVn9jYMpr5LUkWHhn66
enAQBcrXU//mzliGqUy+Y0Jlw4v0Rvq30TfooGQDKYf2AzcQAczK6+XenWBCvvTJbc2UGNHUMrod
o+tzzClFO1q9xncAez5Q+fpXUEG5RhvG46cD8qCSaeQe8xXNDWfyMQOOPoVmTL0s3CTk6CaGTOx7
bHosbBLdE3GF9C0IIdN0TM4/kivRVwc4gg8F1Sc+ASEHXbWBmR907eKcy99nkPNaod9ntPmvWUPh
WNw0SPJJ6aNW0sLC1yam9MftrLT3pKJ00jhRT7XB6GfLu1E1iHebgk27eFMKo+ArngHVzumbtAZh
yXiA3kCRObAn8jrjhi9JrriFLKi0kThYT5AgtHWgdU69T1cMEFLSBTLhbN2Vu1lLu+sCsA4yidT2
MhzfWFayUQITLFj58NJNZRyLBAC2kLT1GZM96aA3ITue8xUywKltOpXvGHFHdNe6BMFko7FUmuAu
knmig8BvZO6hpio86v6noOWZr9zQESpoCB8CYYUlDwcIaNZQD0SkBUAR229VRaB1t+q8lNfOblVe
/sRdeXgnjWYcEPVCgF/h/ooP3gZydpZFmHVoh6KL7RA7b/01jrJO/UtUTVSsIWqAk4aCh6qaiJ/8
MEzYWwTgaZpGuoJhmpYfxde11OKuMIR906F0OaSP2a0/HYVwyuYCwuMY9Tm7EpOjkGwmEb9dv2A3
h8G0cmeiELlGW3x+T1W2y9XjZ73XGcr/aDgex7Q+xVYwcknWUKEO/dKQvDosT4peQ7TJNtJ7OF14
XJ1t1EMmOy1xwBQDJX3dup2n/vX1oUbd4pvWODzfSRLcwB8sjN5cAp0oa9dwlYAu1FgvhA8Y1p1/
2bbXdwcEGU7DSsV0Po9rdMe/kerN8rp3funx9b2OpF8zLy8HvX5msAfjTbGAYCS+6kX6QOVbJ760
BUXYwpATx8INa66qeejQnHVr+Z219Tcu5d05BP/28Q1PFLLTQklTQb8bVG012xE9HDTzubHDTDp6
2tJy9d3qVPlvNgdJrOWZrDsp1550zwjOLukJ4bhYEGTvGJ3eWARjX72MsIWm1oC5o4H/HbrvkpiX
Zs2vrh2+PE2sr9GTlCE/z86XAUVl8J+pvOoQLkzVxrSRUSyVf1T9m4WcYnSbWa4E00JTBb94I990
lb54DIq0GmGX1pz0I47Yt5kQhy/Qt4xr5kFJ6FQ6orFv58AMxaeYyCOyrn0gH+gJ12f9KVk+2USr
bzVH3NoOtPmz9roGFzLjyWURkiLuETrxC8uG3Fx4CU3JeWL8dPV09ayUvU7TF5yMnQlilnM7Gq20
rr7okNlOeg2nHrogHxOwu+22j7+KioLH6YpZlcyZZI2nX0SMYSk5qD7OxVcNGNYtrGwFNLPUg1An
WUggrDWrRBzsP4z9mW84INClg3qgDdDwRSkPeVPCyeIzy5frI13F7iGNeWp28gnQnqmi89bptYcc
xrYFdqsTMOSPJl8Dj/k+WtWy1t//hgb8tSfBmXpDQkIuM/vhnRfTlE8XbnwBXfCQSIrbBa9QNYuw
vpkA3TcbH+PsGoX4BEDv2RzPmuGKTDuB92LOH11ZBNRuf9q5sr6XXteYfT+MXbOFFY37o3e+Fu5n
R0qUkHNgHw+yw/Vq06Ub19OemssOpJaobr9ObvjW8Ou7t6Z7pvkgdjxVj8KTNCnBwfeILlrDzj9t
329crZTUt2CDwiCdlAyreRueieXAAeWcYTMdlvA3ITCKEKJIohyUF/JXtBPPO8Ma0Lmi5g2iR5iP
nih8xWjIMkX+GLpQsOFX/zgBstm1SCbe8H37fVeSWcMnwdjJ0kdloAp8a+MdJ2qwyPx7Nc1vQkmD
fW3PQOteDZmV3Ti/5iX9OcMBt4ZpRkeRcb9e86dD/UQ2pUyZcUSLh+BNHV526xwrk7Wr2In+duud
tMdmNzo2OgttGSkvku2NsjdJy4JivsSLN3YKZOGzHcnlFMWXfuH42rShuBuXr6vYWaEiES/xG1AN
rOBFcxb581NbiYfWSmMK3x6B61N/5/u1t2FoMTReRC4EEOT7LnuE1CbjHjsz4TE17mbrB4HqVWO3
inp9qG+6fMhd91xBFyin85cklyjbQxLuwft4yCVj3m03PvnQ7n5E4pTGIj0NvQOJGVM6u6W6UYco
HOGv4melWIFxAUiTb2LU/fCxPEZXxitHMmBl0SXJD8dHBMluE0kSp82wES9J4q8xrj4fJj6tpFWR
WYZDmX73BwnP5byog8+l0qbgw58DKU4p1Qa9pVOuLwWbOi3duGu9AvonSRzuXz6p0LPrCrGNDPfK
j//HxX01w/zSQg10aqadb5lxk/i91clYRfoQm9jW/VEuB5885n+v/vy7sZLUaLD9XOTqhvhJa/tw
TsFFD0cYM/C7znHAJx6X//ZOhoDv47n/VsEyDMKDZ8+zMiVYwFOvFg5l0JiSzZN6nkMKkWcR9bqr
rvXlWiAJ8gBXtCTMJ8joBy2cFXY1A4RC6dfWNPCnlT98IYIi4wDBpfVkQ4z4S5hg4gENVwOhf646
DEbXEBmLgy/+ZSIj+lzCkDMnCTEVT1q2MHVCYvWMAxrH3dmB3y/aZrGNtlU9SoMcPEv7BmS9FeW+
LoS/jBtKzxirJ0CfatiXca2zebZ7fCBpfT5dfEOuuepUpSIadZ0aVv8CxESRvgkd/QuBZpACSwFh
FT0i/2k+4LcluHiopUZzwmNvBM03E8LaZJfEGGMnTiak4slgebJhtdfoLlUSx0GraeEroG6ShHu7
VC/oyJKPaV2bspBHAddIJO5gOjRhWvgF9vzWSxcdt8L6ZKuLbck1UYOb7i0wUK+7vvmNs6aJ4MuX
2Xu/E7WKBFppW8OZG95HszTOzta6RzvSKbViE6ewi86GYRjFvLOU7hNaPkMekXgC0azMjq4kpIpd
HKihNbYI84e5jre1P2uXV66eVaAh/4LGJPXJ7bciMCbGnjgSm6WgNPWrhv4W8Icjz7E1VUSGgfXz
uGTz4h2LUKvKnepU1mGan3h5pEvPb+Jgx7wvpc3LaTPbmbYA2KEqbs/JzP0rlHVyKZsMDWkH1v49
5IsKR8fYYRZmj+tf9WbvHgEmuSaZHFCFpn7h5DFAZRR5Q4p1zZTuzdusWeNeUzUONy4jsPAPGx7N
3lhSpNiOIKMe/KHcTR9YxeFb6Ey7zC1zyiqzgHkCHStj8CaS4QaAnYR6sxzypAdG9LONpo4MjCEN
dKurOguZakf6Fcxxt3gFiz8kfvVPhHrR/Cb/NRQiirR4Oy2ml0TiBr2b1r7uxag5ccO2vdWopAmv
SvPtZBI01KYkQXgFkCl3HLBoPd3dbtMhJkQkYS1TVo4MvjGCyiK/nKyJSldhDR3pOMOOOkqo4+n3
3agYAnKZPKwFcy4rCtR3KPxW8c/YFbgc/EfHdcGimdCgUmfbjLrQmCQYoaqSf1gMha7eJFeiTq+/
jYxB/d++8nleLoXjsU12A1A/1gDOcgB2zwx7NHbNudc0mFCaNCxgS9PBCgl1Ujrhw8fyeGqMOrBa
tOwnKtSo+v0uwHrjabL1MpYaLtaR11Sil7peDQaTjR/8gw+0h5LPRu5A9mIOWj/wgXInwncej+9V
+vZ1UIoBL43QjiA0Evcic4hcSARpcLgOLb0IrUW6fRbfX0txzdbVLrWboLfmEe9CD11VIuN/Kr7g
PVNq9O876D5v+eiGp8DTpddMWxHvTttxnIln5V7BoGuZVs+yTwmXqY0p2c7A4kVtlgAmyuxGDCmj
heBE2FNvC3JfkpHdELj1N/b4k/dNG0feYIeOWvMjTitx8zTiNL8rntOLR3NpZczAmAjFirpH9ekY
eLP4JG7wMB6WYjHGgDP6HfJRYdpUOSu50caBNrTvMkDarVF9OVKZtJ8dkABBYk8GyZ79wlqSy0kh
Re2JSKyP3HMlxtV+WMw1fTC5z2fiPhjy9hNoPGtnXSWit4lTDt34SXCs6/7jZi16/IXMvoZrOPLO
0EApvXr0TPGf7I1yPvSx6olJPW+70Q5/D/ZASQmngi88Cd3FXejn6IdtJRt5Ar3JRUy2B6yXN6a1
KG0Bu858qNZAKlCuoEsZxXduLld6gm1GRSjfYrGGpSIR4JxGlPRLOuJ9hDYTe+jTuOMTkHs+w1Of
bVx3EyVvYKC8SMp/wjeY7Skl/SRq436B4XYKC1ErA61LSTPwyglfxfwd2ivVwb3hHiuyUA2awfF7
JdtwqJcvLBBS/akBgXKNzOa53foPN/ejnyMXowt6yFkCH0eSI/MGsAwNQRHfF8F792t1WwgVZtqY
nWLlfavha9cqAv0xeTM2DmAOJ51fmaKvh8doQYpHjdo7AZJKfjgyr6oO7hQrpAuAOXD+F2PoCYgf
N/biH2/rLS7WtLERp6ti1r70ZDRQHyNJOrw29Bo4wfm1qF/d2O0EphUg1BtneFYxrSU73cX7yWMg
OU/SjgLX2l7XfcPNzhTi8wt4txDEVvwyP9HjK77cx2Pmu2OkMmr8uPUVx+Ptzv8qQyVf4SdxrWUE
jxZpMh5Ih2baXmfrfpxXA6QqDdaqa5gZB9+FddXRP7mHneKwkFUmqF3y7CsvQdSHDQ9NqGRVpMXr
3IE6a0QC4kdEvhotQMDImRso7XC5GnrMBrHB9QQ4arGi77hRXk+VElWh9aYCXY6hyVpJmQfHxBnK
HwSqlH0F67RIBh0xha2nftvyNsyX+MGyEPyuFj3g53E/w8PI+9qwoSMfPaf4ywD57cT5U1Tk8YHb
6h0WXxn7w/cllm84tFeLYIge4wF8Y44UkkgSXOnoJq0JU/3EE3l7jnL7maOirx86sV8F4fPrPG/C
xEFd/pOVPZyFxlG+/ZCi+Z82//VvfQkRnj4zMJs6Da3gBNpiTlMpCUqnmyqeY7xIQWb+eL7NKE8q
nuvTA/7QY86vCQE4K++XkYS/f611RKTUW5AcN9sgjWnJY/+9D/SLgEsp++VZzmzAQgcMVerncNMQ
ozWE3ca3NfZZPHUcj7i/AbAKrS3NlgtraBOnY4DI2hJs6lD+CDIkqRH25FLcd42yk5dU5qx5XDno
1xXxcf1N9cb5TRZUMi5Y+EZUAIP+BT6OnzW7gud7aYteUmcPfXnR66JpUnYYDv9zXbhQwWukeYMk
pp/Sc8Fp/c/3C81tDyOlFyfyChMGReVBPmU2TBc3TNsDO9014Llr82Dgy+QHFK5xvKca/Cha9Toi
5iPNGsujaL0w82yoNZqAL+ugYa3GO5M9JqI5oOjcBhIh3vQIJehmExr6oQ04aYkjpH959IU/UL65
xKK3ISO4iyWO2Ak3li/hy8yqGQ8b+tdRm3IOdPLMb0mGqPj6wtsnhXkgi7rVx+dKhRZXhU0TK/yw
9jKcwQITTSvEPc/k6qZflJkL+P32gDdmrj3zFJOAKB1JASufMBz42PqO/8EIJYXvD1B38r/t/wFa
CMHCpMhp90JTtGEHmBPZGpJbkpzMxsLPSP02p1rzKftzgmKie7BD3iwx+WJIlE3djgtf9RWyfzNn
sff9oUm0jtPPxSj0M9TblmrAZ+3eGWVD1/pb2W9qwruAzOkjvEqgHJYDD2Kk0XVPWXiKuAPjIVQr
eYP/qYnsfjjr2ZOwcn/RBsuI6IRFcIjflIBDfs73zB2uLJW96XAXCfSmfTzWa10WWMomRH4yCnP7
MDrIng82v5Fbb7QW59zq+aIVbTJMzxEodPlIYuQ8rFD+uxkJGqLCDA29XgdH8xNrrnPQpKrAbfDQ
t87FyG+1q1QLVdGEiNtMdHjsRaTFxuvBgikGn7Dl7quzoy/sQWUQglZoUorJf9Tq4ZqfMeJAYFn/
yEp8TOutJzl3WDW61kY48c1gq9EtIcaF53fWrLq1CkyQMJMrcR3+PJVrGOC4DhVqcCZkIp8SP98V
DHjEBicnAJZaynGf4rPFz5Zh2f2OFQwjovE3nyvWPd3fGgFG1xFGFAGFKl3AhHarLB8LoE8zD7mK
DWqlEJtAcrmvpRglP0HH+LurVMJUZJxdRtQ9qgwCe4d263v1k7RO4KFMPFbyL+XFNhdtqHGcF7R3
v1bqt7YwF6PEchZ8SZ9Y/9EeVCv0sum7N2vjkXoIFZ+yAcQNfRp1MR7Hw5V+yVqeKnsOCzPXktHd
RJZK0PBmd7pHBRRnNx16VOBXlPNeMq1Oo8WOPHOZl/LI8a/rbkKHm8aWN364SovUfk9CcC3bHDca
5fL6SGzG+tjiyj7e1K+g+uyBcp0C8lxTucyEWJUToQg1bjc+ruWZyTLPl0FM7NA7TOHLddjdFlGP
tjksaAnTVciixeuz8RpEDFuLBK6idQzNgWPFH0SxYrvuNE+nZAtkXVQsOcdAmZHAsNgjuJSPF8Hs
vlygg7Zq65t6RFkcwWBygTQKn65p5IRkwcLadSQORk91x3OPpFI/UJ9aheAbOIsTv2k650YSMWPd
MP3GrBGquIWPQq5NeNcY6K5Mp8waQ74jHxgaSY15UvAvzIfsl7n9quYYg/Ekl8UarDVH9uEf9luS
sTKK6S5m4cwmHRO/pSiAZjfXWtR+a+5dSEhr4NmVgc5ncZM4YaUoxLpGj7AkG1mMmlI+x95V9F2G
OQ/En1CkJ8/0BGQIY41lR4I+aHr0NzYrrlY82/1zHz1NPNmKd5nj5eL/5feX/rrSQ0ehV/40eXtB
NH17HGJKviB0wSCmkNoyh4uZvNqlvo3V6/lgoU5gqtD3wY7nUfJkL9mT1rc1Alk5TdEWiJ7P9mvV
3g4nZYlx5mcpMBAY0bbXL4bl3cNejhZinrTLoQ3yKd0NILDavvIcl3/jBToqSWTXAiNcQbrgLoKN
M9xtgN1Q5jWx2R8vIc3jTeW4/mHF0ZqGqAvZhQgttWZquHk510ilfTIFNSnqfkl+UfRt1DnIfDzz
14eL4jmj+AELYpK3RTvO84gHZx9OFVF/Z+k0LWSffxsN6c0Z4aqrkVL03qf6yUarZ2K1yhCAXV+A
JQtQaZKKUcnukBlF+TKBsfN1ilEojcwfOnkEhCxWTGALE7PEJqohyq2I0sWeoOdUNsVN0eJocvM5
g02OKC+iVPYhEjBlyXnJzEZtqlRvYBhQE6QQmle7FJY2dNtrf/5yBukiguc4DO4aIxNgKZGnhAkA
BvDEWM4omTGit3ZZFp+hMUJPWmiD2d8SJOphSfQcAWZedPKfwNl9Poax3dOXWBnlZK9viZ7Msu0A
tBAC1PK37G4NZCUHNV5A9tY0rNLJ8w6BlG/KciIAYACOnGDikuY2hpSmL2T6gweq/RLoXiXhn8J1
hMQvq/JFVYLOp8tRsSHdpotACksLmkzO1+4HpfprYFr72Gx/vScho/OgI3PbkaW4hj1PcYYUCaug
Cn/r0DMsdAEbwPKnknJcwdFWUZ2i7hJdm0ALquRVOF1hHGxiirtnrhb5410CvZMweEFbDurH7Zjt
Qkeba1am0IAFtXvt1xjcH1+ogvjEH7OUEck4e0Lz7ffeWHrD7fSUTu4C/KcMbS55rsnKF8mz9SU9
y+7lmM7EH6RAvSxp/EpLw+XCo3uIsp4GhhKCCEGpy91TlXtxYjpqmfv0Ts00/KMd/LRuJRxLLbfl
5i4fxEcdvYIfmKMvvVcxCsr1gwmIl1sUA2UM84Le0H3hXfCAumHGB8uRzBTj2aPph//GHUNyAh7z
FHp/VXsHssZEAXnIbJmkl9B6yAkH30CxivYMI3yL/wXWYrkGlnHXZ4LGiz9tO8G1MeYT+0rx+j0l
6MssFQyMwrqZKWGLqDUuzCD6QijSS21nmSFzD7XvNI1EwUzeSPAOjKBYcw+fSlet8J+Wmz3koK9d
JiQYv4+WSfc2DNnhVrgfOI1wiUtvRxR4HVzaewUPRoaptRRt0x8/V19gDpW68TDp8FFsgVixsE4N
NGWvo80fXIvC+BUiofr31onZP5HdrHfpA1WWnXPvC9TTAOM2VFo3EmGl4YDrVJkbEow7Vg3tvNTe
PAX1iFsgDZGvlkLdDo3/9EmloGL+OhfPJqY0KIr++JS+A3G6ooB0i9wtbJckVfgwqLwC4w6IEanl
VuH5HMhw3EMqdXnY+RIGm1FouNfyvuFgrGMk8WsCJ/2NeNQyj3u1XPdM8O0F9teWlG7zwYqsES6k
BoH75owECwWysgB94MXaVAbqKG4loh7KPIoATRv1bvMk/ycOAt0SgKyBhNvS7ce/zzHBCa7pF0JB
M7GY/7nSQYNQhph7kK+T6HDQ4Y01IijeUvubTti5HATdOW8E8SsDym9wri3xpyvvAju1b1Sqh1Pj
PB/y24Bbv6MtWIVYyDRZbfQEKe859XlC9x1ps/MqGtCwebBRmI5F/pQtLEKlSaJA9CgdEMohHyOt
ZoEkz8ruI5egdWPqaGfj2/yBfzp3yBZwiJoTb/AStotadHIcXT2wmbgZCR+fWDcOttR7UpLk2nnu
2H4tWJdTIazwjBXBStBoZWdOWs0qcMVrxVU0DJOTRWSoCW8s+NVLyHDiUmOjLK8E7MlLc7QvwfJI
8bRNm3qllfjYkVnygeIWPedrOYZGi1QqIezEn4A689XvHLM9MzN8ZiSqbdAoOyQN/VW3RQB9CYcy
6ZkCiE0gg9dXMxg+KEk7A+QGON+xrH1XDIaoOz51cn2zel/tjHKtN8ml48NQzqRfoPN32I/c0hLw
nWXe1Vq97GjAI9VaJUvE6NFtwRBmD3fd0MA6XPHmb0uf9fS5NF53cs6tKqEhjM60h5JGzwyO6HCr
/tnTDM/0FXudEeISbzGmeGsGRWpSJ/+pjiQBZFZOla1iU93djyT76RSWz2Ve/4ReQc/1910ABYOJ
0V2gU/qN4IZPMDyUD3oYnnR61tyDDw4nJ1EnGWJ1A1Skqp6Uhy5uc/Yyu7r1J3vf11Fx42XOCss3
AkzbYjNm5K/XRLGzaMFmBUkUmimCxNyzmUOsVV7GfwAghlfL+tfLyuyaQZruqJAP5gQhqC9SrDnE
/BPJ4qcBBWJ1iAwquI6+rsxHQguAqFnW/bWFocGjxCVCJMDyEjY2RGYycSflayUoDkMS+j/Noar1
JFVIUtI4zSZ3aMXW9PpUI7LRKqfOFJcl+jIv8Ko7YTcCuLr5bk4NuP6sohmLr0j7kxdbS1FiTaH3
aC/JXh1Q10k448WzF7b+Vb4Pzj1HPJwM/Vvg2unvj3ENnPe4cge6wUfsVj+csTvs7EWh37rzn7rT
1UV2YAn06CSrTfhxlx2fCJ8KcBHbQHW6nnsHL+AQ2GZbxcANndkE/ih6zDl42OIGM+kQeqESL/1h
FVloIjc0E7BdWo2JifKWImgj+aTij3kEIsJ8eTVwl+N7cRsgd4WmsEnwEtM52IkslsijFHu6ZFSI
pQRiKyd1xOWo96BeHf4vuAwEi5CIg9r5a+28/ZbN3Cfhj8TJ9HTb6Aow7+Vr67wKIG7fiaOtnCE2
YFBWK3n3UEFPOKa+UGV0rU4KV7sfkrSlqB1vuU8JiOuKhc6J84k/akUdMECuxel/rgAKTPpizJcj
V7ZRER8Y1dTcGwPYk7G5Gx71cNMWO1rYEbRtbQhgR54XMK6aqWty3cPnMp51q8WWvntAcUIrCji9
cg/5qSUFVCmNtd2Ogrbr0FseVHD7vl8Z+QXTeOZkl7TSI09y/MF7EZjonqFauV1XIvXLOGVOnJIL
EI9Glf124oYM2yIQOYu5Sok0TMl+pmRskBuY0BzGxzXxwwAaLvtBMtTueb+QDl/7bVS+FI/i0rg6
06MVR4TbevLYitmrg3JaAkKYk7cAFs78uRXv6rJ81BhBQJ56UvFUulraGb31ntRHdzrczrpCNIoS
5fxBrMp599ZPUKfx0q5EbiIGdB7+0VGCm58Yy34+EX1dihoWPYucwuGZKYtqxGzSx5ip+Sa3l1/J
LO2uWP/ZpDWgWWKdhlivJz/wnsHmNXxgRGLqQEpPaLUKgq2ijBJNJRJ9dTJb9jEhNnezfvg1qwyo
ALGi9gr8eTckkZ0Mpo/XQUtEaHnoF+XwJVQGXorqv0x5b3X9BrDkty/wuScp7HFtI/mYe+eGKQTG
cvPFoRSjoiMlBetV16xRkKeKq35XOGchsQQMgHhN/eqkCixVaCmFNQeg8WM/CZTDWx8sHhaVMjB+
TNgZpOPBVqnR0sHxBIY934AJOI5ksjuodYO9T9NnyXbgWdbNDyqZosEUWh3NdIXuMRc3pvrAUqV+
8IsubgKveswnxOoY2X76Wmx+GMlTKMlBe5e5fL44cTTKezWHGqOvwEcRMsPrhlikqR+zLiMQtvmB
YB+yKp888vkf/ad+lKmMS5URg37y5s8Its7zvKPVwctmxBowsZzsmnzq1rhwG9HFildFzyrvOt+K
lT0LJ2JzsUEWfET/g1rf1K+aCr2Kza9exkrwaGBKdTfx/FSg6pHDlYqmI+0SgonobCAw/M5ZhBPV
AvRBLimCDyyhmLVQbusuqvAqx1kdrxtB+6c8ONTD/X14e65ZiS4i6Ra5qmd6cSrKnr3JpR2HI8TI
Wd6uZBCvI+l8ZlT80RiCXgY6GnTxNPrwJPiiNxKwfGKi6WWIRC5WLm0UfVkqt/kNNU1EU4fc+SS8
Ps0xzZm3+2m+SKwGnxG39KJlCO01v8F/Wk4xAq66TmmF813HqGdVL9DwdFkioezRc+GbJAtO91Mo
cvmtBFE200ejO4ElzaZyv7QkXPTZWwDlfkJ0Fwh3ACRbTLAkp26AxNdbsllksK/5KVBi2o4SMu9J
Yxrow1XDs4Db4opDwmrJrLp5okrwopxoVoBLQ32TkIsQpPP8K0T0JvAA7dPAmFyldGLbGEfUuxM1
vhW/TB8HkIU6uJkCVwbA/I8LsybFc4WJ8NpuY6k2ltrUPyFJMQfetuENXRdHT+UisM4c+zxwOe80
oYqdPeGFaqb77kSBFvLsRT9O62uTrJUxmnZa5TRKcmP6LtbBkUHw4XTiLueQjqPoS6b+CRJIAEZx
6u/u18bDlvAIRU9zU0wQi5S+SeutgT2MkaeK6MFP4yjMbowYKSHpRH+oGlaZjSFLc/oPLelcZzZc
GXy1fhuG8td2VVr6qr2fjeXxOczuqfTUlDxNuxgOHlzvRANGNzTdFOxVIm1xT+goTDhpT63Aj1fD
bQT+WfJF9MmtWrX4TbqlWwV73NsSfv3GMQIT49EacRZIZmzWKyvQiK9hNVf6pHFOot74eMahmjKR
PrxVJqMJqzif8ZJY6lrT8f/inu+zdKj3f5akGAYv8lyKDwqGclKMMaXS0cKfZgHDghMfkT2WR/Xe
mR4OfaJvULkgtE1PWj70zfHKxaUZbmv7LLrc+IBcMc56Ghx9mwopvPGij5Q0V5VF+F6kup81TZh5
irPQI5Hz1JcYreDUNLF1y/T/NCo2aLWwUx+ApzhxXJvZKQ/cbBeucCjN0DvFaG0Qnvaa4eR4B9io
ZhwX8bWZaAbO1pcO3jVhaNaB1c/UmuQZOUUOqKVOHyvVxBwCMAPZJr3qjIHp8Vyn4YSJps5bkPPO
EUtV5XR/XabjJD+MTL/o3KTsEPwx4SeeKE/1xn1s7jZImczIqFkpjq+J7ruN8DCSqBYWCj+4aBvA
oRIl7kqhWcWpV7SIlYYgkKlqdZZ+Upwc19VGf5y4Ao7/VSbLA65F+waCZV4U3NmG1UsYguzRqGIV
lQoDk75T/owfLogcuO4y+BFVOKp3CNmU4mP/CVmvEhaMA/5UvBvvGiqF3HN1+MSRPfhy+X8Dh4sq
qQlUOskzsSfcUTrr18kiwayLA41b2PVZEUvgo+ZoDU6RSjZ4myKYO38JodR9byQRTbGkk4f/w7/F
seFpCd9a9/3hReExXzmkI0OaYwAugVt5t9Can9YRAjTKBdkCOurgavEdjxUZToaJEuXz+Rw9Cd7P
p+9A8kbVVzH7dYdwF+62vPfCVBY5nYUUNjPHby56A0SvPuBHo2BTOTv/7Xstm9hbnJqKjcusqowT
RfXECSvKSxrwBEw/7ncHLlK4qAf4w6AQUUirpcI5qZhjUj9+uaK6kuH8/Nt3HzC0vpeecuGmLd9B
JAYWbRVq6cnjceH5WDwee1ZsmpzOyg8OAOVYNQ+SSH/B5G2veOM1qMMY5PcViWChXuKNEws7EQUA
sgkeO/xsdiNzqSAynMXOaFyF1VzouT+A8f73YwRaWEUpXSmu+rZBr12tE+ja7ZZNhLEEy1cWNvW+
B0Wut7Jt4zVj9QOEB//dxO/zUdyCvlKf5l0PeMV83Z0IW8UvGBe7ulirQaacyPh1ZhbrKUSpk7ly
0XeLv8b60/+EdQu2y035bqRuyBG8VrzI5cSmh0oF2qn3Oc1+9GMCk8YbGnL1oJ4nboXeiWU1Kqze
Lrcnl1DmUXyC7h5jVVD8SiVzl7n6joo1M/bUQC/BKt4PCv1WNc6LeOKcTiyUDKSxLpdvVdsA+mAb
stwxhxuW0YQXyvhQ+vMGgu5vwZ/RTX1aPRDcgpThHZRDJ+J2QOL7+tFGK1dKaBLb8uYqPwr3rEHe
PEuP2e8KLk8D2gAFPSQA5Zxwo6kO5sgHVZPr+jTDZNg5C05fFihM+9sViIYc6SeFov3q5hALbpGA
wUanB64sQ1r5LsrIuHKZBXnK4NTGmgC8HV8iW2KaEGwoQbQkjxC5Pgb4zpleNbSD8Lf+zIwTHhsS
ieNfHehekkt8gCFQAnAWy/DXhQPTmG5xzhPHUsOFjk5nxsb68wgAhUTgDPNw8qK8M7IEdEHX8yTr
3mny3PBHnzYnXHsxM3iD73Qhp1JhmAI4SB3mh7T0kx19kKMmAX3Tyjww+p4GbAnLMSL9+XAmfSq3
dHy7gToghf09O0ysnbaaQL7VGNzprSq0+ktZGGHR8UYoI0oJgIWU3DhcFM+gVX223Lg4kWitmv4M
UvGTVqW9gTYtLMbdS/kPNOq3hbNOH/O8HKHYDRkCLnGy3UixXorgvSglNM3zOn1IlVvWG96jGi2C
R6XrRAfX/2BSIUFeF6sUgDhXB008KptWYtEVNXLGmq7HmPwp82OdJruFZcvhtdRzKjg9aKjCjN8b
4YQ6s/iU+RFRmduY+TmFGIwLE+GZSAn6xmKNfJoIKMacy5viEmBcL+mnQVk6Nho5eY/gyM+SMkKf
/EidozwzEKUznbOlajD98WfUnW36xXGLmewaqE1PDXHCEK8O5LUx/sn62tKPvdCnKCsq0H6nPiBx
iCXm67cMQMUx7/FM30dypmHtMD5tM3ksyoq6eSzKQvs9dPCL0Ujj24aQzf2fwUlnJOiG1whYo+VV
u6A0BGVeO+HWSa2BfC8j8XKDtfRyDLZFO15JBmL8Cx1MA48p2ViPByYAAQYkn/a901Chs3h7b3Sd
YmRSV491zuYsM4xuOH0Twt0Qb6oJhmHGuMGlXcKKPBSpDp3sTVJN6btm26cVxNK8/7JdJK2osjhm
qM2i1E1XgbXKhI0JkorbWxj+LPKj9YOp4eb2reAULBcbdpsMW8bMIUer9su64Y96UK/0E7DTTv5Z
+R7bJ11vKyhcqFL0V/T7j2yTQy5/Kc3ri1levwUv67srgoauK3n3fGDh3GTvU1Wd6x0rcTtzejPO
pkjI2r68uiQJxnxRd4ucTkLFNPojzVHxMW52NksjynRpRrq6iFprYRyXD3yHRp2VgbX1VaEiMsxz
Y3GPcXrRD+Yx5edP0bnuVAIjRHB0tNkcCrJrYHmq9HsmBa88GwooyKRpUfCFG0b8DCeBjdt6A3BZ
uMgcqhuaOBvSuUva3K/VCCM5UAQ99sErrtcVqB91Fu9y14O2oSsjppstixI5pwwIgWJql/po/JAT
meBTFsUFWcIaJWqicSFqImnDJPRvBfLQCutPWrGkdDMYEXr0fZn82I6vJYHAJ0ALpjYaund+kNrs
3yBwoOGKF/B0+dNv8BVHFxWffLpRYMItJfW5dxf5O4Iy1r1Oks7XPaPpGFiyec2E4xpgpkPFPZE0
Io1DDD1msXs/1gQklGiX+K2JQtBqvMnytYmsjoq0ol0mDxngV2U3bxI1hAsAGIsY8QE2KS6V/Zea
k+tN70whebv9w4mksQh6Nnl/G4ZZUT5aJMu6I3D3OgxWVtWPtEgu2NZaNm1c3kWwkLCDGSndITQv
lUn0r8WXvFCbV+HCOBmqAmPdfUsLRgi5L8s7I8LhHfW9af3WeieIUYPQUefpAl+wEyXjuK9WTJcZ
d90FVBV8KNrAhGuZ9N0JrjFt81umxKHwxHzcj9OSBooQT1LTOySO7qP0FgwCaS2LC8wDxh5zZuZ3
Cq1WXrjamAwfn27+0nlVmmYdkYqRB4HJrUNPS4tnUlhQWMuYaWRXNKKxVXADT128AvrXYhZ1zGgd
X4TuvwRTWVQ0/Eta/KyvrgWPPQuBJUes1CoEgPXvaMV7YLKUqpOTwclYgKiTwkzyKq/MjMZ+Vmnr
ONJZXgLYeRIMQYRfJr9rMjhNAw4+IpOdcGLOP34HmLvTIyaPjYCk98sB3/bohzGSZJg12Zv+0wv+
dTohSTmUUocC8eCprI+ug2oPbuPsBEOJdCCVGss8jP9J0vgK1nGtkX75b93CAaNTZgWJ8DehJG9/
xejRXLPkjwlDu1G4jxqiwBe27kZvXh91N8F5HdPi1muI0VczCXSm3OQ85vsfURV6i/8OPe57A1I4
98QudKiV5S4PMhNZnwVdOWJ1c4jtSvcZD2CdO2hs4JEDd/JIMT/IGzHJ7Ro9ePTJUuvB/hPdu70d
iBi6ezNadaIGTxPAApilOAbFJO+V1VASdXjV5oPA7PXkbVA6/ut8/UnCqrGVXwtX7U66Yce8vs/c
F6JO/JNDFj5UTxjYXMY2NNxF7m+sxkeC/xRLPtHhxeu0ep1UCLJsbbHVP2W+AUrxU4LiB/HKs1tD
i+loTHvLvohBU677g7bSEcM38pWcamK/UIcT1VKtVmTLoBKGBR+QPTiq57zTZfyLX71xIXy8plyv
9wt92orlnEe66t02E/wSHRhPVnrP1o1xS44AgujzgwKemBEgF+AWZPmObcavAsHouVGTX9eil2dD
wz+6kZ9eX1cEj6Qhz9Akv6Q421YSzxkEnSBSwijZ83BU8e8B4khwk412tyqKsnQyVKj8q3k5zNCb
d0qSmlyMG5Ew5aN16FhVy/vRwU2C5LMdoNwu341VNtT9xQMKHyxm1lZtGxgjKdxEJtHL9EcKShb1
qXgxu3BP2oGsYyRZYjEgqD6fvJxjODjgrsOIv3sp2a8darIOOeXq7ITbSS8Pk0vKqjDjjnNOmUKD
dacqzREi8MncbCqKxFfL8SK0lt4FVasKgxjUA1iKC/zmiPdXG6m8ipAGKFwV3sa19VRH4Sj75Xm7
antPjH18Q8jQkKhoDdgjtXbA9rx6ZUUnBoBQkaJEWXf668hpd0l5MamAtK70024FMYZqQ8j2Ftyb
QI9ayMJiZFl+6LmTY896CHfQkFbe4b5Az+KAJub5mLX9hqT+5NPWA+3JlrdIXUPIZbaeVPuRsAMS
8reQ1kNQZwmUt0A2/wg+VsCGRIuQaFe3AjqgTuTnBbuiMSUTTOTksXkOok14pzmuifMiKb3xRyag
LU/aqAbvdxwW67QgDInm2EsEq2eCTCjhl+pOtnYpw6N+QHIbzoEfX/qYqco1Wtz1KVI7BHNajx01
KsIkC3bcPfFWebA+B+iPVP5lEFJ2zLmPjSe3afkZw3fb+Jyw2i7dE3IhghUpUKbZczlcOAbeVLkr
8aZa0Kc37/mDy18rc6tP5Dh+8IiamkXc+OIbq80O6Tt82/7rxX81wORJYdl10QLrA4PVTS5SJqGH
Xmu9WiXzMlk28rPcRYEkiYu7rM3+arBL3oDcJxuwwVc85hEV6J4V+ffA2S9r6u9axJrZzmtWM4FP
+G1NyQVTwMgt8UA0BgHk7RrLVRw4ussVleJvewehbUCNPvc5fti3quxJ8DAsbffClo6ZiifVFi+R
ifVQVcx82V/z+GozVPIFFJkVf23kDqTAr+wBOlF4Cn87HyW1g7weAKIIfbIWLjeKMqq9BeTNjPgi
ou6GYZlZhZaH8mdmzztW88LdzUa8nHXdTv2GyqXUtkMxXHg1OrQURqRBQfMY5twlG4hgD7SsVqo6
tnZZ7SBkr7UivHwaXb2nYiAvDVATBAcaquliCjWTM4+mWnycATZhC0hVHIM0EWIwBKgTvbfkX+lm
Wal7f6jIFnHPPBrOIeWgZMGY23si7Q0chI+taqA27gl4+L3I41MCqjFHrUewKR4Vg8fgtMi+JARs
v3pRNw9NOsnowVxnEkniRLtokaVhk1wC0B1XSOTM0wwDEdaGmnFw5Gx2wje4slyuDw93ZTk09c8z
TVgeSk2iOPqnZFOdOY+pxW2KcA0bAm0t21C5b6dFiZlsrkR+rAbUPg69w2nHkvzx1cM4sdGbdji3
hBKRRcP1L/k+3TFYMFCJFQGHEwukNcHZUUb0EN8s6a+t1XDo4TIv0vsCHlHNS6S0l2D1mIB0tGH9
FrKJrKE4nh6Z+s8b7A8cDubVleNLEdFRSspUUyp6hLglyzue1aCYlbF6zd3aTuXQxSf7FuvdjTjx
Gj8sKfEBaLoJdzoGcMVNsTGK/2654OwEoKqX9E/ZYNVM3OUsnWOoJSE7f3/saYVljOLm+lo2qHrl
64whHYHEU08bGwqKPUcagOoupx5hyH4w59m+pSfUa5tA3sGS8XenJO+QVS0q+qXblD/UtDFilWLV
MqnbwTRXXGGf0C6c00qZBMOkz/chWAbdAormaCauWKTD0s2T9UXobELSAa/nJ3nbnBwS/3YvT7N4
0d3Mq7zEeo2rCCaZiv655uz71DlqXTGW+e2j6CluiuWRJ4VkQXpHYkMhPuo4NOctOyAxg5AFY3Cx
VUtkYTevBEfxjlqPmVGxG8gvzXd/5QElNMiDEC3COC6pGq8/sBR0uMZLypJIYGR1Ihqhe7CiwOi1
U3D93Yk/1HdNEN1coL0sz+W4khDn2NkA8MgPZ8zU8Mud7qWr6IjTD+FQNUVxO03wRk6kmvzvbQ6n
qBpW3ssFNAyumpONj55DNKy+SlOwRzZgt8dKGUJ7iV2WeMdP9oiyCwLdzlu2+sn27ySyiDG2ltGQ
DNnX12UQo0TW6Tr9Q9nRw9kmWHaz6qyesehAh1xm7vLkjwtfWa6QaS+e/phVxrXQZkkTj1WEa+uK
Re9G2DVHZRPpD98L/AY2QslFTbv9GcojxfyWx7uJV1O+zDufojrJOnLQQg9Hyg8Calo0tLwmJm4s
2WO21ygLXqFyTdCz0rBQy+BJDCXp0jGJSKR+G0znMz9zh3oensXbUDfn9Sq4Oa1aiDSodUVd9B0V
ekynbqUq61N1ara6HlmI82Ds/GMvEjHflXaaJdArttYEShR1gfxaTJbgnqNO4C5gEdxpk10m1XhL
ZBfqIWbSYVsg6xpuoRKFdWBxDhdSL5q/vLMXi6AQS61rWuD+5V3pD1jG0TY4hM2FMjGSL4uq2/DE
K3Ut+7FOb/+DGsMrw7rHx/eBqMqxx04AeqaRppO3H3Fm7WsqlihILlVyiBuDjvhIizAgmLFaMXc1
vRwheymqcNtPav1cgM6y4xSwpX3gIDlFxVFi26S8isxkn0qJLL/SoxpozSvS7vWb0UVTtRGf7oqU
s+jrHGp61meIBneclNAMYzZV5TGrg9tSlwlgX/J6ArUW3EjoFDC2A6Pd783rR1NnBM161TY8Wj4W
h1my6C4RoVeJFJhQ+cc0MCJTQ1QfsX6x1FQmxmfGJGKoZMpDZCg8skWJTGiNJdVv89Ox+j7PLKOF
Q70vHKbuKBzBPaQovuNl0jk+wlUYtURULNXyIBi9JHqAPl0hBqbDAlEqDs+AkcLTJavjjxW0Wtq5
TnTNKKUQFxlpTZBro6YG2DdQjEyesG8T7awqKK3PHDGHXv7/7eYcpSzyWfOzOPSBb32Ad8j7Sf/g
s5DSy85EVnqP7Gaz54OSA5VBXNQ8pq40FoOSw5AfzSMnn7nIqtnLsjo+osC1t4usWrd2xor0H0/W
jyWWt/VhnXJkYB+Jun9hYhORjN6TnmQyLyS4jAwh7WLX46KoL5SFV0dtAfUkf+YX4TLgR/lzgnZl
EotvffCDdaPb66aUVZLHpjxWlUpvbmoho7wg+qSCSxTPrBmAbPcmgwGmQe9fqY0EUT/bDPE+8Sng
ljhE7srwnciNvvZ93AJERWwB7e0yfFX1LkLVtXyNP0q89pKUNSDCkmMfAe8Qssf5A6VrXUennKt5
h3j8D/uBMQRfRLnvg/KSh/rtErs6WlCn1bJ1TdQm48jf3+fAUYyOPade63JihSY3C9YbekMWYNb/
BAAF2cri7UnBux2Kp9aQbA3CwQCkKvj1Xc95U3CmaTb+YBMzl26Z+0M+pAjt4XmqyEpbyhcxVgtg
0zEjE+KFnifsa9k5ckj686To+Blv3awkXr+/F8AC+5+1ALJAWuK5Xjea/zXlyw8FHF8qgDj251q0
JKLqK9HT/x2ulUDp9/6d6cPZ92PJBpMAUAmpHj1pKwFQhT9Zb9FuL4Xfy2wKI/EoSMbMQqtSlFqw
11dQeanSvmYSTs3QCQsRhWT/3sknoMgMIRq7fiuZsZ/biJnUAc1h+krLw9PmVrAeRhYCAWPxmCHz
iXVO7RF3MeL7GORQ1zEFST/CViIQrMZA+iup6wop4Qovdy9xL5n0Mssz2xt8CMOZVLpuGVrA1qbE
QrR+woe9uqFQ1uHc7ghNNrhpzLWZFJWY4QUrxlHo+k7q196dMD0mZfU51evI2rP/3D1/RLVKotiQ
VnLo8q7DM/xBGgmcQg/UVP4HJhkpuvG4TNWl6jnOgK+5Vfp56TsU2cGnhxEoUn72uSEmM4AJy13n
w4xXW30pHA6H8srzbc11jKjQ37a8wRVJUGYrDKBwgMz0UN7MWHdrnesMiKu4F/IueiKmBLP4v0XA
xiVz8ZsQSvTuMmYewPErUrYksxz1zQxwEJp1EMLUmPb+HCLfypFZV+52pqMEHIElz2s8h9NJNE9T
3UceR84iMg1xl080C/pgOpdaTflfEQKkVyCX8FsccyAC3n5iRhB0aWo6mO6q/SMM639p1AGzmkLb
shAde2mJeONyW+xpdgPU/Hyb+KWZcLF7KbCkNTsfLgEpbq8UBAlRHyn9Phtn4Uyngtd62cQ+y7ZY
P/82UIObXKH54aI3MNfuF+THuvOXfKhZR/i4o7+vkFyJtzstpXfuE2eZYSvSxbvhsH93eSNsdFg2
KJBIHxeCzQZW1KQWpZGVlZa+S25quW381IMcNvrCZlAtbDQyogL8waVWS1nfNy2BRdhjqdTpXQFQ
5M+NpwVQzuSFwS/xLzk8CJQfJZjWI+p+VeNltfV3jqixH0x9abcdPnYF91OcI7CGIpd+T0XdmiO7
6y+Ogl1ly1UAcOnCCoPPnZ8W9UJTf7qnNLr2otaz3ypc4hOSlp/OCIgSCFpAX5Et+ETwuXPY9eom
wSiTrPtd57e+3tc2LPAvrWj8CThljE4dC1EeZnc/nItHWm2zInMRHtU7DUeAVbXdsRjv8GV/RhK7
3ozCUJVItxNmLMxd2j/SKdiiPkM90z3XWnRJoXroDep5s5S2qZqTul3cLRr0RpWanVbnq6bJvxV7
HqTFDqA4iveM3n4J6eQAzXtp6Ri268N+k2QlGaBiBVs8+qTPp//zSGhevCa1UoLhI5mQbta94TMS
2DryckWrWQ6Lqj9W3uQE6EnehOCaUt7xZsz+RlJ52S8oZLrJnBepbMN7NJVDKNlusLvO/ObHvdFK
o4uuqJkkHTmaDvemikyDOCbfsv7Ulc4dRv5Iu++xQqc/W/SQfoGRzrbT/IGY9iPsvXbmeKEa00qd
enA4yOCafFMRiwZjdGIJwPjq7RuqeNga6PvbZwr7Kc3ELOlmI0mQ1vQygGsGPSC5NMMhYJJ0t4JF
BfAkNkY6KfX+QTYmpivCEUTRuGWJTtFmA7ilLr6kbvT+8fP/MgXpjG2gnX2j3ojAEu45vlwlqnho
uupPdID4mhh4rt+V7zXSKN9ArvbMjtNSaCeLVWtifdf1upLv5cLG8yJBvZbDtNXPETuJukxEzvSI
KILaUfZIvvSyRL5yinmZFZ9FHOCYBTaT/UeorC3n9GE//3Q0xS5pPJaXeOl9wOY1buSMfluubsdZ
61DXnHW7nXcPGc94tKzvdMLJfgghralOeDguIegEUbghuOUp7plL6VdOFCfxj7yU+w0CfPgHh6jj
bfDKZ71Ab94/vAd/P5jGqXQ3pvMjFuS41wLHPNkuAE01dOgehIFS7iJKPxz7UIk9LtGEfvkmMGH8
KkbjPpDOzb+rpTOLNhHLcWpBBh/3Nogwdpk9L1ExgR8oGLH3EduUuqt9Fur7ihpGcFJULZuzj79c
r9uGtqBMYEL1IPzTtIyEnmYaEEH/yeAnlWToxrlLaUa10T0z3tJYIqGc8MS7lM8RBFeVDJhdPuW+
zSq9FjxPhjTEkToRGHKoKjZl6DNgGwY85ywtIKtuzx0Kam0jyEw5KMKakLrEa9T2ZcLomHSM7OgP
X0qY+8cFB7JRntYrYbkWSxuMEstqZfzockdBjvomWWllBfcpbFSLcl5u6KCPiEOQvo+6ToFGruI5
9qEeqshODzaI2CiSCAj6DSm8hA1n0BEv/vVHKiTdeN0NK1c0d9+M7eLFim7WEFbUJstFPW3kBFPn
5hDJVQxTsrE6RJiq4jQPnicFSKwjywEAmX7jdTVMlQ1YHMA7mNy2qyaD8Fovx5V9g2SCFD3Nd1sv
/7YqqQUfPiMUGVGv1PRMr2Ipek+4wISgs3BMHemkia9YI2M4WfRBaFJfH54zSHnBr4DOJHt4ZCXt
R8pkqSPkVHBvLmA5AysCxE3LixhD0JMtv2aALawaW+Tljydj80PLhL87ERoqJdR/11rXPPsSad7R
3O9VBuCsU7SmZe0RIcDNfDUtdfRDCtdIk0CCJfzgcLvHK27MZyXrHlE+g8WFC9TFrpjYZrTYbNqR
5GhZmRl42WjPfjVyCXlFzhhjZ3HC3pYAwJOPVvS3LptoeqIAPlQi53HXQfwjQEzwy+403gv6qZoq
lgGhH1XtbO5JBQm9rxX4isTD0KX5MgA05EErkwv9xpH820EhKlH/zGTCC5ohe9aOebt8+Qr11p0j
Q84wUmJ6v4hKOG7PxpQ8tJEe2qrSXE4Pkzzq9hLhyct23kJ1p1XTOA39u/p0pkAsH2BPmQGZqaW1
Zwa5SWvpLt5m3lSVOCdu8mb+oY0beHxwxH/5fXRl6Ou1fqpHhw590RxrzQ9SxX7m4J1vp5IIdbWa
Ir6lRC6OozH2BXFaNYgsdWA7oQw+98c3I87khzXgPAmnqdtr0JU4ODcsg44SgELVF2oTI9VkH3hN
GelODmwj+cZoquMhyJr3k50TUebxaxzqMAUMwFM1jjOHHuf2eVbrdPpT8xgs5Cg6gzlHbLTu+WTs
bM4brdA8Er2iEPYoMFFSSTywrGIzi/lkzxAT36XadARTyV+oRDZEoWoYTXgiijSrwArjyITq7SBe
CUf+AwOSJ0AisTXfG0gEkpIYQvDUjWdQaYMj6lFXUn0B2nWFE4qAmv9WZwptzZ67HgQfblU4Qcev
AFnnsPEC/4pz++ccwmG+zxPC4axqO8H2N5qpysmRu+uACo+W1j6f2o3NOWfeX44+/Fukg0dVB/kc
+pHeHILMwrvLtVyMZzmVjz/KJXP5QzznCm306tcQCtJb82gOcJLe0X4F6X5jnPPVJpEuIp1nQWex
MZF54q0sAyL9fjhf8eaQyUxNqikCKEp2JvEanW4jL0wS9WH4pWTc5+KXcjDKIUCgOCSvD+9Xtmna
K9AvPpppBsLR8ibNFjHoAoLjSxSMz5ojMscSRUKFpObDFRQN7kkrIu/KLvZRvCOFr5kvIP9ygPGb
PXiLZzzrqksNqAQPudVAYsufg/CL3+/bTtoMMEC3PF363Gdn6yaEFAxVeAUR9BNITbcsC4bjm+6g
Lk3xyHD+M1yFKIB8jrkMa9hYq6ZX6gYoc5Y4jEMoFm8eZE5bARbU/LHJCcyw0QG3f+4/IE8ev/BH
GhZr1bO6eeDE97eZOapUAV3iEx9O6E7quzExWsXRZuNc+yS25wosg6GJyXNl74cpT+SkscSmJimj
xOq3lt85RJXrL+Qp7HnbAzfjBxBlFYuVjiPDtocAaWipbzxYaL930WYd3PRwwo9aYOYw59bYRHvG
UsdTcb3ZvCWXIgQLV8xvMtYOXIL6iTN7wmYEng5vkYC9PcUnmd+Jg29E5ve9mvmzxpnTSxlJI5JK
jBB9ivbVvdnUhspk2aIoYi++v3AWbAX1aLax6cfDSYoaS6jQoUVOnaYW46MHPI95IQqZPIT5JUf0
EjgJ9HdRLbq4ELoyvOXeRxJVsxGE6/eZSh3S1i3UEUsZWbPc4Q1q2ALuZterMLJMDyZJFXhm/WSA
3hxPvAaDm5Z9I+V/fo5rSvwnxjU6SQdWYBhIGxOdbnl8/qVNIY80GnZ+R1+n9PD9wR4vfMZhr8Cf
OWumtAiP2CQ0QNa4xLiLF7MabdticwSmJ5CV/f4QDnGRMh9WUmX3uBvitxeoQTo0gdRsqtVRV1gM
XsgDtxK3PzbId+3Zgn02dRyvUUYLFknasNSSOhkPF744DZQ78YQqlLffnJE4zYN5nQ33EdaF7WC2
qBBuMg01b+/uJ2RmiyokMDRgYw9HsoPUETdA1qMwKMzGrA9mjdAJgUf4tGPwKq7Ck9bWgG389cjJ
wt3vicWpneukHtCBrhtXm0sh/Ou5aYv7Lt96ft+9rdNFnJmEVFNZOfOUPrnxkY+YXqqqCP1tjYxg
He9XB/Dxz1j9O8hTvsOzZsiKP6i0VRDM5K/fixfr+lEhe8hcN+GG/wrJUsxmdHyuVZ+6rYflCIqJ
U7WbsWpgkpDN5lLeSvWsKb6X3TT+karLv2Bt9BgONyAvqe3/Sb3mWEJylOkpoz5jMGLO6jdNm56w
5BhNjMp8Er2IazYPMHgxWwM/SRynY6xZXTSUDemfBxT9Z+GXYkDSattHWQuoHPc2tDkUGs5GWNxs
fDCBUvV049hLnkVPYEA2ZCzMBxYZS4lndg10V+m8f1oPmaOGY0XsGqaEzepTVGpR2qpQ3zGoorqq
ktS/OldeAjUEN4Cv49cBrxnA8APzouqgBWdYSAZV614l/t0i2pvIce72bpZm3uSd2KuirZtuV9ao
5ir2EjalYuxhTPXEkMMvWETvd3Qku4eKgHRL0zHJ5vFVedpRFcUMxShlCpkjjJTPuRvsICtVPky3
IabqL0+tBTHwTalIuKcqDMFqftv3bJe82U7irc6Xgljs9DydPaVgupGr9vkZdJzq8US6kdCqJUmj
8bNIErlheA/Oqs+h4p8Sa5eex/bjgwilWaGD5TVNdg8IdsBhDNo/fC4WnetQpWCH4DEPsWBxfY6F
2NJyI02zZ6FmV9+b2n5HfY21Vx9IDAgpixcBcwLXWch2Xf6s/OWMYGjG3totLfmAX/bdp0W+b0b6
onfkcbQv4JTqdhOSgYguPjb8s+KN3HGzKGpbnlVLYMszjSfTOT+dM8fY4p5b8T10xOEyLNZTg+2W
ilql0n48CE60A3qmHvuJ/ZF0a/eZGLSIJepBrUBozxeyyPz+KVxDVGDE7tnNIYPtMQF7/Pc/mCUO
9y27axqj9h5Qu4kNwAHcXM2XFqFAxH/TTCUvKGkxs78RpF9FK9c744wfygeTBXVwVph/iVq9ZaPL
dY5ipuznjWqjchjeXwk0+zwuuCtCvKZlBYRZek/Nz33SFo4Fy8gI5w0vVeWHImA9tzk2U99AdF9g
K6QfnOYFvJdnA2Co9dbe7/lno4RFl8yEbOfc8S5mffTyQRXAkd2JvFxztsmGxZRfolqZRguMC25l
Lrq+RTN8/H17ma2rPSm08rfee2YY5LCAa+61oAIQqNHck0tz26wA61UST4741Ie+/tFtkYfipPht
JqSUpgUINRi+lLQqpQZmrteESiJVRrTPylLFZPulRG3zWVQAsX5mqrbGowHsAaek+NhdMRfaGaY+
3eFBDvzrdfFe40ORITABYumGS2ukNz/Vt8ahnYK3063yWFHCBrMNuxFU+cF/QZF8IOW+3ZaKoB3z
bRhl7DorEdL2SgROpZaidfXkXCWWICF7f2xB0TEXFiI6rLkHMwXFLBzq+7hKZCE5uFit9M6YZVrx
OAm1kFinqJ+NGXQrkivGqR1JNvnhhCrxuIMDzhPt+ynPmDchQj2mLrPNxeb66i4ylmBwqw9E8V7J
zN+WbB0m9lh00pvbu1JxaHiBAjy5t3Z0DP8q5XCxueITDo8L9Hb+mjJHrk+5hcu2F3xVwnejheZX
PrS7iXJ2KKwNwn8UxvFKGROuV2+q3I8Mqr1L2f31hGyVFyMNzC9IaofKP2unbJ7Mrpo0BnvTo0eE
a1ua51j9eydFzmA7+GJpj/LGqZEUhpv4xjczLqL6Nrirt46YNqL2g6VQGRJbSL4WgBUhcqU7BNQl
FZJ+oKR45w5pbFEl2x7oOZvAnxr/EGKCPK5ra3Rt0D+6rDzBLst5dhUetqIafMYVNKa31pM7ZtLP
YjcFMYLmM+91AONlI4i3kPgxtBmbkgID/K6Ulk6tUNbj4xB2WNrxssmBDWdvvetAzLlFEEcAvB1Q
gMt+MLi09yR91+9GlsZBTaBNgJpzVEL0Tr8wN7M9GIGlgV80qosvypkdqkjcVOBj0S3bby4QXHNl
hEcjobiHvvIveFTJOwnE2ijNgMmkSktH2dj5ohp82H6BrSHPZlVnJbrdRVJABSgWHWh7T135hgue
djMXg2duNxiAC23v/s6QNADIL+w4I+fHJLuH3WoFntE3154exjTUDMqwxVO6OPpVZX3vbsqdMZZi
v09w4uVaK50Cdi3IpPlRTBkoAIDabottLScfgdv7VnOAfGR08UaJ396IUhfISK3HNPicA9BBdC+W
9p7u+W9hDjLe16Q3e3X/hM2ppxliOwzBWmpCGZWaBvb9vu0gOuI1WUYEgPjJH54BAo81yho4XeY5
IT1J1CBZjvjiJzf5Mn+SL7KgrDlWinhIeBp2BUIrfgduE8RPJH+OVn9KpiQNjVAubA/E+aACKf7Z
9gw0xRWUZZos/82LQVthe37Ny/47KBTjNPA07MjZp6WUTfIUl7DcL8qTDOc9cHvDXSgmPiouKBbm
RSQnC3mUBbhV/Na2ZW0iiXUbOXXYVJy9NZXuS8M+Gloz9J/0fjnKHFXupRrEGArdS0mhlXcW3A/J
6yjQ1WmEHjbNiDmlx6hIBUcYhLAtYAjf4K2ePAoT/2xp79BEZ68ZlHVm8Cc7F25new85rNZujmvT
sG0TmhF78Ms6Zqi++8bNSRlfqzVdFQfUdo9eg3UxUIiLr9qKNRztmAZnIMrV1DsJzQ40MHer8H91
sktpe9os0yUDE7r/IrWW1MBD61WAIMsANZyhdiICl8R4LvMcuEr1/+LneexBoGrRgNVEe3A36tXd
4zQshOPHPlx8fzenlkTQ5aEhNSmx1628Il4yqk3DdJE5u0BROw+wQSt2gQzUourkIuwcIlbVCS/t
nWAySdusTVl1WLkUK4oiPW+xZ5nijGrdgJagKLTwth7x4lY7x/cT0+Gw5PLd8h9Uir0LwyQ/f0QT
lOee6x8/QurrINjEeBIp/g1LUf3gTNdcpP22YUiXeq5BXEmV3NvSYutRvOvkE58yfqP/BpZaYOFo
8XRpvtvm3NA+U7YAmFVzETrTuEa3px3hszDSHqtGFSKEvp/nF2Oi0nKOajEMT4vcQxep24gseU9F
b6w3bCy2Hz2QxljDs15JhORwXzagkDqWFQFJX5ZiT1KhW1BSLfV9HumEELi+0jwmcmZaMYUJKzPj
imp4R9zXmbXUbXrZuknSeWk1yK76IU3uhno8mNysH0K98EPTYfBef1vavth+bYlzwF1kzaI6SAkc
t0EAb0rLvMcS2EuB+VjgB3fIy6NzLXIVWy5wYWEaEgLJeKW+6G/JpoT03w7ct0IwGCfIPxm0sw7A
Ar6Z1Ixk2yZaPvO65UW+a6GMGHd9UDSRX49NKvdc1HU4A1dPcEqXxdw3C0KzYi953+halpMlGQTn
+p5lgd+400kKEhpI58Ltg/8RXf4OszAdUu4E2kgisa+imLsTZ7S31V4c2+NRDAjGm5VOupSiRTyS
SxkVFLgatchpS1WugLCz/hSt5UJluDGz4amHU3h3s92mk4lgECsVyHwGfz0/WE/MtZw8G2SrAmJB
Y/Wr+xh48dQ25JFOcnbXiviy5g3KhdvUUnwJW9zN7I6YZNUSImHDFhrjFSTNy4jTGaBZOonX+rKi
8dwKauSAUeEa9KZy5ZzCYztpLsSt3sXYZVw8I7P1zz3pKOcGeeV10E2x7BFKmDRJ4GQNMynJymLJ
kzjdK1fUqD6C3A7dVQncMua85hNmxN8cIc0j1k/Ph3SAt/NuDzxetycUIbc8b0967b5fQDXpWKIs
yAPfGGSe56GnBF1mumWoXHqMveeg6MZ3Y4HEm1Do5b5fIEdHBtFpCHluyYeTMzAzlg0N9i8/qylS
jSM6vs/73+RJilMY2C8jZpc56Jij+yDT6IHYFjhyTnmq/F85tHEe2TeHqx/3MMZQuwmyw/ngOEgE
MiQkQgrNrv11Lo+r4GCmTZaXHu1aM3aVgjuoqS85p+YFDBrGRrbMM2guoAZs9qQBoRZNcgMTey8+
vcmMjpvkzFkuovaJoPVvuV5VCqHAkcuUvg/qzCELJMpYaz0QBSHGNJ9GYZUx2lyKE/watMLiS3fV
86JCb6FToQXv9IsqAA06x+EudR0h+Ckvq1zreauXMkETpoL5eQt99sNOtH/LrO+vkW5TmwqdRIBZ
JdloM50rjxKtlf+DZGYyeoDFocnbjLtViY8F+7uxfXqQFwUHMm9Fo3KOTGncmq30DoRVnuCs1ZHW
OC2QE8d1Myl0N7Q6Nh1/89kbeLYS9Lyo8OIhfYaRD09PAKP4EdNqzMAK/q/32ooy6mKWwWgDEViE
MydDNQ0srBN1UQiZmjoegpVpV85yLI2xB8vRU4WkVdv8Duc6PUEHIKLXc3F9RL1chcHPOw+h0Cti
0f2aaVQWlPqD9x5FOLcB9ibKtzCgk791PsDyPdju3lSrRgHp2/lRQV6JOGrs6a31k6eaGheSCP+7
kDX6T131MehhunbHgH2jtlLJXdW7cu/FwkPe3iau1hy5U9GnMd5X/khrKHi0Ss7m1AEHaPFJgD6Q
8R8ATILbOZcwaBfxtIY92bZjw5pdiehwudwDyyWd/CXsoHphyq3De/WymCeHZe7kqMGUHjUfOfkA
u8gWDVnqVG+atZLA8LSLdX8e2lf8solp0SOmJgPITcFiaOTdopWm9c3//lPSM/KBqMstVKjC2pdr
4r8pcnq28BcWBUy4bm3TEcamZVmw4pid7j4XO4vygtpT1JOLuE6awMKKo13lEZZLZhQm2drPr6Du
FHQIdEqqdVABPp3lw3DZdk5XJEyl2GOnk39j6yRpj7nuJolIuOzanL172iHMC7g+x8yh/XhGQgQz
U1CJV9/L4Ap8RGUYkVpnh9tk9elVPHGWG9qm/Nb0IRTLDmBUC9yaWuzCDgpuRBTSgfGFFKjA4YIw
JHvmRkGZ+1ZOFCnAa6CLGU15A6VORzs8MzvcyCwrZpvo6Ndem7jCe0DHhazEC6Wq9O739JtUUqF3
KqH5mNvBjANimQSzBprYMBnNfVlz6XihLSaz8vCrvhulrRFfop2r+zFkfNSxTDmiFBpHpLsSIzgC
UNuGlzEL2oGtbcRRfXGYOzCB9Zav+sU/gLZa+SQNdBOU+YCxqlx0Rf+pnvCEgaRIH9n3/3b4v1Gx
N0x9N5aGmedFSR+doTZDrPbLi6ltlNU9rMpci5636w2PyYmfeKQPaQx29gjfazpkCl8Gwp+K4zQZ
oV2xUDHcFqNJgXuwzz8rtkSMJ9IkwueBYo8ia2x/8mhJT1oykAL9KVhWMMiRp3knP8QorWxnzPZm
FJG2K/iRGdr1Ji2WW41okSXIJNZ1/iyry+CxxnJj7Wl6fZihWZ47G/iIXbXQMYUZuud+/hKT2Puj
Eh8a2UTAD815hMPoarEZNdTkzdkKqnTsN4cD07STg2VvfZKeQLJbo33aGk9MWEEw5Tmwf5gHxF2q
G/MBpc/oHV+a61UNy6N1zHrSOg4XD8xsZ258J+aGM7kRf7qabL7V2Mm1nIAv+rYQKsLk+vsKfyZQ
uA3jm+aYif5iDBJg9A6LuZo7EMX6wICanvgxcz/zL6d9KHC5mathur91cZ1ULR5MvaeKEc8JW7Jn
JdTWVUYWxARO10FxwOQ+pdSLK3lhsE/4Sp33zWETqEkFMWDmBzOlEY6CH2O3cyK2WgDr4NbpAYXL
oeU6ep9w1EBfjxWSyAPwWcrC8TKeOUYOC+QOzy2nI+nrd/V6Wh39BAhVSUKeJpW7LLJAgLsdPrNt
Fp4fVrAPBKmQQd9+5mkblCkOPI3NLFWY0nBGJQ/3QJop++121NZkE+vUKGv9OBtovqOEDzXh354e
D40wcQG5Sez88EyOV2qLL9LxcEMFcyAF6uCopp+b5SuM4t+8Y6iFgj355F6dHYXlHVfFIR4NZkT/
xTjcIq4wr9iXoViuCKu/3uhlsQ/QdvBa8kbt1U5muFQ1vk1s4qVpVjI6yBDuzfwPMJmx7yHIZt8+
wumx6P6XlIe+gWORIGUUJwer1+gWhI7wvJPveva6YXzMRGtnCJD21eW4UJy+WalvUw7y4gY7A/vj
HjtfvExv5Y6uHagvKbOcqlWymQTw+f2E+EiLSyYjSxGFw+HHbUatJsKaIkeHtSgHBV94qd4mAb7Q
8D7CnJh7mvCMccbbghIRxTWA+rjQG5vF9O0g+/O18O7gO8s5Tx7fn1zG0huXB9EGm2bu7xV1PZEi
FMyUpQcERNHCT/9VZKmy4tLAXkaBvhv5T44bG+3kvjbxcf/6Mv5ZPD7MMCvCRy8cyjvN/RU2T5TW
2s/Ak9me9YsmJwgh80Sto0uEwPQo4HWbXuB0E7fpCH1YKNmLz1g+7HxT3dw2OwkdQPXAl0xzdA81
1xeNpsgB2TpUNFXH/VNUptYOuOcI9TpearMHBCBbpT4EHW5pqGyX1Oa0B5XgfVcqrkmZVpMt1wzc
B2LHDprvh+SxgdtVrpoRUhuo0JI61Z7DwDmvimff+Dgj7ilvr+ta3c6I8itUWqbvm8k5qKUTo+XH
UM78GmuUnSEWWs/qIuL5wNyifWnGZZbt7HwRHmjGau8n3tWSqH5JaqNwQKc6L0OkWmmLftLigPRK
oR07Okyi52bwIFxECdyHtJIn1bRzQlu2M86gJi1ATnQ35/xQu6xsyoYgNvo4Lfd2RLDUxn/bZO+X
+aRFUOPVmlKBOL/L0Gr+HBZjzt/P+t1kpyV5jnCd1jdMwXiZUFnUK60795Wqvt/OPf5zakogA1Hv
xHeo0yxkn6b8Avytuy2LO0nSLD48xTySzJXPAya+mC869tG5LZrqpB9o0DLnGqMWq+PcOi1yxDhx
VAIQ+ySloLzg6V1L4a/ZBYL7SprVVTN2w0TB5RT7QDKd6aXhut05tpYRJ5i1c/YQeLZ4bHw7Oyt8
lkob39utA67O9Y2JQqVv0QbZCkJWTnHPxOephk6loB9W6Y9GpjcZ4i22+Y4n0HFKHSRbNyZtfBqY
+4Nm4lNn+7Fl270IPEIRyqBTFfxj+tdtEMvbc9w2UpbIGmBvcJLSxzX4fqDnxeCnFjbsS0doDnhg
61bhM8VzSV3pxZOv8nOvE9DMYSSZUjy3HSBncTt6PTEXO5ivXaJNyzHcQp/HC2TKTvI5M0U/brwh
J1lHbcChwRU1LifEDAMZoXn2yssczBuUGLyjTqld4NW2TAs4l9dKz1B6jXAEbBHDC/J9hKsLnGBO
Tfeo09J+MrFTteyjEWbt/tneUKm2cZrmH4XHdX3N9yUTvlbO1iVatGT3IUje0x/PGeQpo80DD7j6
KCHSQCJrmySZSucewBWmEAoyCAITaZopubDxcbFj/CN+jB1P8wSGM2OucZ6ZX17RioKIpLmZjXJV
FoQDCQ+IR5iZu9eTjU2nG3AVeM8bdS4cSShP/bUW+VDd6T1jTOYKl+zvof5yf+8gI04nkoUx3Zy0
9nK0FCvkj92gHZuM/vnrVwjEu3UvMMWmOGUKHEVkbd3Gvaul3UpXQXhPDMu4wAmM2QxEG2ncEWb7
9lJJIDfT1sdCQgW596E/8RiPGfFqiDXQedvHfMmnFaIdLzHaaCA7p5psne0jTPKI4uPKdOaTPN5h
woeUnH5yjJ57hMLvxhGzGIk+ssoDqaWVenoutCwRW/AoUSwcDDQm1yrsmXe2u9DcOYTtrbD3PSCR
JyV28TJ+QXnT1eWpx1VZt6uq/IviwAqzowY6JvYEdU09lWyeF5+QmiuMSDpHAp1YDG7HnQDxpIXc
kn3AelNWyMk4zBi2y2Td39HDBpGJ7hSIalidAEWpNmK/tUhEL8GSzfyEJAZ5PA3dew0wpkrtRgHJ
eXnjHlFL+ulJxTnf6bK0vQFXrXFXA6jzsfCclr65IEU7zzJiE++NiBuXQQ4CIP+RC49hy0mU5EPv
0Y+ctZIMSmdXkO/47EkZYyuZdMOnXlq/ycSNHshQagvirRkQu/V4ZxrQfcGSVI8v/RzEwYhpMrTv
SZG2Yyv5XdsrgJNImd7VjhqdqMIgI4TyjL+PFybpkibBw4jryouO6MZkYa2JENSvyrJR9VNj2psk
63JlZhUHpDm5kecZ2Xnx0UXgaIhmVfZ7oMZJtT5Cxzbm9NhBCUF49Lvq6Md2KN8UyC6wkoyJHKYs
tkaAvKo2K3uiDmyhIv/1GoxfPqPfESwArwNHeiuSgX656ov/JObByIX6f0/BvVxTUX+/gYvlxP1Q
r1XKui1tcKSY0SxVJkiptvVSfK3OGKTcB7lUoyy5+/b0SN7c88XGHJqHC6Bsd/GTcFh0rGrnCBr/
idxPxdMfMH5s/LVHR+BY6F2ROdf75mzyxKm1v0pAcmw2LMbk6tmYSNLBqA0J24DPr83vMNoTyp+y
2FrI/o/3fmyR4nJA2zXFoMPSOZ1sZCvJhTiRTuuIS2GHDWHSu+yaE6YOPWyOXedI3cVi2A8Ti4nJ
Gbyn0/p/eaeJANnIZw5f7DH78xYBG4oUwk0vNVcYl3oQEcISeUfHXhkqLmdvwJp2xw5nmYd7xHco
qqBj6Bfy3S08al6DyItOwQE/9uaDUtHHs4+3teRngJM4ju3tEcmwT+h8A59P2YRE3YXXJCjtHwlA
05UJy6LIhv2mMxx4Ku/X7LEOOYdcyb5VO9VDHFmcYjbRX+9YKCQslUqvwWoqm7anHIJxIed+DpSY
tNSKIpUGOqeE9uOONs9KFEw5nIDzKrcah3rI6tEdnuVKck4hIeaPuTBukTXv8Y2YBnxF6dXqqqgK
2pA4IQpCawwxTjuNUbEbLzrlty9cXJ6+8tKDvtQ03WoeTs2Rv7t2wxNCrkR+E5mKlTmikCHOykQE
4b17EF7HukAKYgTQlK+heTwS8FafUNQGw1asMSGwwr0=
`protect end_protected

