

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YqipQWc4JFBZb16rc2dodhguFDkilKhXXsYOnDVSNRAjtkaR6AZEesZX9P31kdm98GkKMNT69IgM
oU3B8PoxIg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Th08Wi4CTujjzYeFPRrbrk96/H9lqJHT1fOXWDhDkZaqyMx5/LmUZnPHzc9Mi1qiTcgVKZeTpkDd
lm04xNkvaFBlZ5KAxEqjMNmhtMTNyj98wbYe1WGtUEppm4URdSaGhgzD2gvskrJEfU0HoVjNKsYv
Y8g1ek6gYioQSqVo4Vk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3ST6h9XhpdCHj0//nno4AUPlABBr9tQ0cisrrim6ayZf3P6t8TzMqSxgV/q0TD5pBIm//qvgm7Bo
W2S1EUuvf2WqWkW7p/E9CPizeTTEZkAYHckCfZTDk/HTJdolSIFeCHjfZiRizq3RlOIw44CUEMSg
PXhJE4sbT53L+d0eIaNmJBJnZPN29vIw8LbE7t+Y1oivoLSh1BhWy3+lZNV30PrceJFjB3Ylx53O
r9RULlN7k4FVXKoCkEg9NcpjWNJAX4azHw+uuE/ZZmEDfyzXMbaQPIzErM+LylAQ/PYfvIwSeBK1
4Z1Yudv71r62qTHPKAu2JCMEmzvKCe8RAmGoeg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iNgef8JJ0zz53Cg6UsIY3rdr+PhJG3ZSgPvV55cmHG2d6Sfxzk8LG8+nTrPNPEPV7qefhOfs2qwO
LV1XGy8/zcDatxxl7RZSBTwjwXvbpgbJIb3oKBLjSbNQOSIIh7oK15z/NbQ04jpEoFW8I8unz0Dr
X8lH8UO/ss4o3sjSRmY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gdQRq0TszGQ1sYR2djmFoWhyazt+0Tw2kvNbiTEjaM08h64rXWx+KrfH4Ux19p4jnBVjDnfhSE44
xN7ehFd8XzCnm6T9eZgkCDf8dP3IGf2Nl73ZHXLjDsXHqpK6BXZEG/Ko8+LkLz9nw7Snn2cWezi5
seVqFQ9T1Cl73kL7otmtLUuX7sR7LkwbgtAzFivUF8Ml8V/izjdNdzsqpzxjHY9vo/n9JWZSxDHg
dF+BgQSeU0ooY6vwulhfUyi8hYLdbvSFz9Xlr9vUXABI71kCIOeJMQA6BrcWbYjoGqM7KNL6TTGp
K4Gc5G7xM4ucj70Vz377eDl1W3KXvVQRmQSA0w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6928)
`protect data_block
9cN5LHJyxcWfFkjRN6skvmr3EXEzWNaV5xX31ijt2exvjtbILr9DsXoGiLeRPopLMCoxRHRbIVYU
tlp3NDYOiqJUHEw2b+oADGQy5mFB8qCmvTYVRP0mfzHmY/+oiPGKjatKswSQp56vUOmNZgaC35kq
V4eAzcQXS5cIv3wyuBu4NQAEwMzp+eMUnz+PGK1co6f0DQApeXOx9NUpTU2Sva50Xe9lV/zKYBPV
EhOf+Pxq9uzsm9UuN4Vqx+s3SaJe+Z6UdRo/1gj7dcKUlzdL+gvp0KyhGzSB1UC/XGkj3FYROwMs
LsRcJuRRTPf6ImK//uEHWUYMMNhh53tN4niQsq56dXYWWKzrgaMsESegah+mNWOGOg7MVDCDpb18
uIUe87lg1PxSgBd7J92nsRUzohh+L8Mwo2IM+vOwShNAd+AKNWiRN9rMS9zIkJ4oM2knyak/pjuZ
ss1Gk0BdQjpPbEzRCDTt+HP8aN4YrtllEuQGUiGn/EEamut5BgrEDIxci1NGF3wjeX2QaZX7u15W
N5EyZyfVZudICl8ZJCWlJ28iVEmvb0j17B4D3SuxQgDb0HG4K624VnSwgCcZtzSjsOboBtxfyBFQ
zR5tJEuMjWtl6yoT+8OaSh/eUG+dklFp/I5anLoc1Geb5NNuMDumkPFg08U4sNzupRzzU4bxXgn+
t8AdpXWXYaQkH7lpJUfSmY34xPAHplvMQt1a9e4IZE0NU6kDdmlHvJ1dzpMe1BJPt/NIB4/2bj8u
Qa7Ja5x4lrDHmpBBqWZMGYa2j2bpMtQTheapuMa3cJmx9angkkovKErKrRILz7SGjKjYSzL2pkFw
e+Gsc9PXhjmWUFSdtAu88s6fIBUvpQB8ajydmfR3Y7b0jVla35nP7cJPBQwD8tS0MoZonu/WQy17
uo5u5sm3BNTCKx9rOdHYjb98uVd8dRvW1cca5Ln6TQMcrNiczi9xrBd/5gdars/tv2s8T8DO95XQ
FMcrU5qO6ToRuMqSFIUgQxX5i+q0EBMdrpMhCLTuOpHs73o0zgRB8YwOYZubb19DtPnO9p5fuu6J
VXZg479/CKweNVtock/RLn/on113XQ6GzNMnwNYSHwsHKDHQbEotwWMSf6jb5Oo6XBOocU36ZxaE
B//YMfdU3izY/bD7U9CH6ZdHj69GJLSD70jA9i8rT6531++5GfKnn4boIKhrp4cvlWaBZyjrS5Pn
m32IwgGt8TKNprz9kIZ7JMxNdAvHX9O3ZX7jnZqLPxctarRrCMA74J9wrJQMlFuBtJODGkOcBFsq
dhlyYPpVCW0NGlpw3+HoKHKDRwh13acsRyH+oIkEIR72TwQaI1acdW3qT87gRBTPCHvfGkKiUrsc
PSnGTjd60ey8g4S+uYLZz1eQ1VAfIcUq9V1texrKzRRXV4evtkhRh61x9d2xn2KLxKukWbNl+i2Q
/hZOyrSbmKIkdO3c4CD6lAkdB5J3ngw5QItA250s27XLoTqgiHCLyHnvCP+SVnhL3lpEjztC4VoM
0tXP8ZCXbe7hYhZOvgHUd2NQFmuJf1hnND9diXUld2pZxWlHDlvd+5UxPS/26TMChG38O1jhUj5Y
wG1BhpDtMOo3OYv5AxhOS0lo6jct0ANpPsn9i/dHX79XAi1Nb4/XU+oxnaX/2+PZMQ0BOhRo2HoT
TItPLS75FKIsqSEiEi1edr9EhrikBd7So1kOtucK14Rxzaq66aeKdaPFqZaDKBoBmm2t9xGbFp7N
KorINp6ddG39epdQRjSTmV6ZyUEAjXD2UtgS9Td5hA88BRBP2A2B0BjyCb7jo7xgDChi/n23fauM
YMCqzH5y1XVEKGeMD5L2zevP/2vWOL/xIrN9Npgq4eWV0Lni8fFsib+E3mApB/ZkFKB2RpMQf/fw
twjBtzSrI8FgLFYh36+t/igheRaKrrYmwn13VDCDZ+fm6sXS/nX1eQXG56VjCPX9u0DZpdw6XmKm
ZPIsHeyVcPIdxsmwggN+izBx6UVKidWnMj5gNeJWOgPXS95uyQjJbdE5N7dAe0GaieufnhfNH+DO
2xJt9rn1iOnd8FXRPYitv+Br9umzkm4iT16wPQtlElGxh4hGYJ9pEbFuAZ5Jq3HPOtKOpNBAfWmU
47I3NcHJVfXCP7mTGiQof4bcxENGBY0f+mG6anOzvzPLkL1BadzVhl+TuW6lVxdRbtuyvTv8kw+K
ptDTpew5qdDpW9PNnbWV0oEiWQxRUyPJ/X5Xs5udpgmYhWh63fO/B2+YtjjI+hpNUW16WRdW6dDI
oxud1pKEanVlxTcwljrfFpFtgevL5X74FChQ/Ch5TU6xQ/vq8F4YY9r4igcyObf//KpA4Q3suSi7
esvImU8X2jZnLgOdxyVROy55zHwzPvd4IsXnQmeLWUeAHmNxJrB72fWK9mNUlWvOi9H+A3ZHMZyN
Y0hN5LLt4Zpq/MEXzDkhO/8WVxs2WARmRP9pQJHGCVSmS+kkVia8l4rrsxvEXC6IvsE1eDRh5buz
LKN5+gQAb7SQRm2w4savKQ2pWFM/AIWdV7mOR9932H+KatxvI/nqDiHUlm/IxsfYA9XCZ2bUQ4kj
rClVMY9sTSoJYCw9G/rInKgXZewBt78kNy55sMbTEk/4iBkr53p+KTYIamDvubOcGCMipHi0UXz3
sqxJMHfhoqkRrsSiaki3y6XxTwGn/47EnSZ/6BhdlL8/uDVOLoH+6pEqCBDtYyfGPD+ji3lMWDuV
Gqjah8zKerjHaYGpciBqs8Ss+Z75RK8RPjtkLiZ4h3nrdT/+bT7lDKmU8NykqtSHkYeZFW76d056
fTsLo7H/7op1ZnbzWjtJzPzzS6rxRiFe6DLRDHUSjwQ5CiaJ3K/SI4GRlKGaj/+hsLM4dnnxOabD
p6Z/CyCGvqPdRi1LMDvQrzLotSSKB16Y5PKv1prBiDcjiB66xfsemaaoHNQqkefL9AlP0Kxz10k2
TbIygOGt5M2nY12kGmLnDCksQlg/p6lPjjS+vj1/ZbjQRTbioTvIgMT4xWwSn4oZHIoeTtL0JkRJ
5rq8uN7TOFN1QeTl8l3mSc9gmC72Dtkb+9IAbfmOMEFt8Mv0g8WxFigYASRmqj4HNO+PixUYcOvU
mnEn71I5blD4H6pq64cISUdiSkeJo5Ev2W+PE0hc4nV3j1NebBi9Yo445oGfErRzPm43uNmiSkGU
I5hGrc8qzOIaS/4nCIOANCCAzUcxNSST+vUKmC+QXqjocV0is8Rlw6Gs3X4yNh4ainHdBUYG3EWL
zple+ARKKjT/evduHhpccPX7R6IClMWIjA8DGAeUhbmqXN+L3wzEj68yA2upjM1WTwh05Xt7NqQ7
c5VKCT5eaXr+6ajTJKl9E5vsh4F5Fe96JEOAcjUMEZ34qRApq1setiTaxfkSZg1poJkEGlo2FGLw
Y8nCZpZjnpOdRzFR2Cj6XSeeqPcMR/Km78h24J6vDLpBlLboNGthPA8woziBz2ldFzRGqSQY1+7B
7SBTaYcx0sOCwcT1OlAH1+ipESa73zWeiAuc3ncmuzcS6qnW/ZWy/dUOlgF4bGWzSuljAJ8Q3ZWY
An4q/0oaEmie9iZSMFLc2ethxaqRP9yJ3NNr5XDUKNZPShh+GsODet30odW9TmoUaPa6IrZ9AQw+
FVOX+xRNG70TNDmE0Mrqj26X8pHaBH6z1YN5QAX9h/cb+qEI8tzFdAYIWArQ8Yjnk1ljp9tsGEvr
SpC+aAO3omybA8jOpNLpX1ItCdctzExwWWrJZCNHpxVC9oibowdhWNEN1Qr4ZZL59faDOTQVutTh
am5eO67F+CaPFH31hKBOkF+Kbhk+93bEQTJVjDkk/sy4jQkKkyT7OMVQWCcOYgotnwWkpNR0iVQI
PkgbojHDihxmeqqUOthUypCufZ2RnIbtpffjk+aZifgzXJRbAVLFGYOUyInlgAx581rCV5Ec3JAP
O/N4qz+76dxqtczg7qL8TTOtHFcHCR+gvaPyKSnojzsiGQetD492E9E/x4bvwc99zqn/Xv+r1Tmy
JsuIOaMAecGYMY3Spy8DYkovxC+o5sJ1MxMRPWN+TlI2J4K6YyRTq/0RMjwZFA8qGoQd3JYshljb
ECIAW86Bj145c3MuVIeAy4SYt1E7+3U+0C51k+svdWYZYJ8293uwrgqp30DfFTwpCZ2cssqbWHEl
8l1b3lknc9a5oOcDo2EIYWzPO/amza8UUKR1RkzTwGB1DUZ4en3FqoJ6FO0g8ph0Kd9+MVP5i1/x
W4u44Yoy+8Cs32a/WhQepySoo/NS9EmhB+dE+S1/3cnU4oLuwfXFTIBKs5APjHC8Hm+T0PV6n0e7
0T87IxBEXTBENctGKeGalvR8v/OsywnGQVwNSJna+KPMDNVekptHlDFq7fTc/3o0jOfGzHrqq+aI
MgTfKapaQE3cjg9YMJfy7yHluOxEOhNzb8Ye7ZohkJ9uhJbjDCu05GxpwuoibARBRHFlRj4MEVNG
lUIjH7IWlDnN/nyVmHchiOSrwM6R+QTxXJ90aNgjcH/6QLydxkR49NJupwVOr8m/uJDR4biF7d2l
bekKvAoJmhtch9cF4baoY9VcyoHF1JF4IK68+SBJArCsaFEKo6qXOdtGixBFUlLOaZ9sSmnoXmeo
9fBB0DKm1EYQTKkwoFCm1vDlJ/F8fWyWTqnJGbKKmAGd0s8oudyaF9kODgXYrrG6l9fC5tqN+tcz
43hU8rNgqdE8HntQ+Okb0SEB36f5A59E9mxqgpB7k8feVQcgxU0Y684EFbTSB05Tnq54dBdPz8Qp
mA49fWCrv6So/RYE6qpm8kFP5whmzK5laOh62gFVz4hnaGoM/r5M0qVV61H66tyZF0+Iy7b/N24Q
0soyJeBonGT6tgJjNpEHsGPQfBwqoPUFwEjBxx+dwMAS7FFPf/caJspWr/f/8ZjBP+xq/N747xyn
1130bqOmwgPWR5rPnN95YAgW0ToatStVVH8AOe+gYhzVlYPMSfdxpDLr4pQ7/T0yvZ6ojOP7cDnF
NLM5yvdloqFbWNBiUMIAFtyvzMAL5AOJj3BGMDm92ig0DWBX73fvlgVOMQUW6y/5WFPfiMKXC6P8
6M7mIpvDLTswuKiG6MKOqLr/lYjwdxznu6QkWQIQUFjN+wjB3s5XekeuzGuojFqy8lZlJkfER+oU
tdlayDLiQ4cjxJmcBdp8daMcWzHrBrKP8o3HoL8bBn9cwqTJHgIbE4yXvSgPlzdq88MEWrRJkeIM
DU2M4ccGCmb9FpBiNUKKP6Ir8SmpeZZyo4nXLDuwMDZLW42YNhzfHqGbbpEp/+0v+6eSCpyEJ3OF
c+LZe3cdSUkLE4+tT88CBXbVK7PX5Gb4hXPOX0mgckf0h21xvXdy9U7XwAZDwM0aP1T6NysP691M
BIswdA/L6lRY+SVSvBWYmVvTuZufFjUhMx1DEY7123m/Z1wq/c4c1jjrl7+sp1T2mrA98UdVIpPD
J6875DKntYds6dk7fmmX+BRUJwBgrn2nKATAUmcX/y5XvLdMzCIhHxR7jwrbsZK/4alZLRawVQdy
WDd2VnHQ7NnGUITPQZLD5TxWv+48IrX6/LJ+5a+pVM0ughjRjbLCd4VXgQEj+npiRtsMz4BbBCie
WwObwwg5xw8TLyMuQXMeV8A2CW8zh2lNQoYXHlaAEaM9bH5acWETSsY3lAvwtPXbefLLTP195tmv
ZY1yiHe+Ra9rfkErMoXEqgnx5qHHGgveI38U0e4Gp4QVITG4j1Y397bH6HbGl2LOXgJ5Vg/HR7oH
bAcFQmaRhjgyRd3KMixfea7gdzUiz/MX9c672Uv3SEA4QcHX2qNyzv7kkZNHCOop4knujGUPnQGh
0YU2wSJI+prX4b2iYwGDhp6/MKEPqTjPRE1e66Q45ib8V2ihcS4vIsQfXaQ0e/xVAe6/OyHqsqz7
P5M7RjTQILzovwyvWD/7ZETXD+5FdhoZb/K5pirTzzjseoQvm5HNSCDOoUwnryFJkdENnQdYg/F+
KkFNirrjmBcV6kr3/s/HyGYQIDlBmWnyewCN9ELF0N7AHvn0dIfU4BbVRNoLkS739x4jpqvoxWqm
FjTwsV6P7wuS4WZMpcqfvRjhPC5h5WqWkH0ncYTJ75I9F4ytEFRHe9mRhcu3kcCiPKueLAiK5jdA
cuVME4YeeAm+eetijv+OI6mSBRzCW0oiqgQWPqrDIIkWkwvPN/fB5IFRiOAQU8e5qEL5uKcd57Wj
H86ZOx+Gzqjz6GxUdG2CtI/1OCXBQs67r4FCZv5ywMKrGB9KhDRAjkm91aXLvC1xHfDk2+whhU8H
WztGQGVhSGdnQauO3ZpZz6vBzAP1h5TuDgKRVOVJpTzyycb+N4KK7GgGXzbDQUKfWWOsDCI2KjxP
tXBQKsHRkDXpiYxTecgnOZClf9UZgOmRqIJ4dMI8tmwtwMhTEWnTSM2p4o6UTtJMMM8McvylW1rS
DWn6d9MMlqxKggQ5RGwJaN/l5VLXEX2+eOp9pxgPy6LQ7400REjme1K4kbfjtnkHqcPt1VpbGY6k
6OFJotYkhE6WMinMUtebSS88xsm9b136n+gDG469c1v0jOtPSKtC+mgU7Zh7OD/j62b+vklIzov3
wXofu8IYxObJKT9mv75TSiA3vwCqdVbyD4ZbEiw+BGGdt7HSRbTTlMZMrcp6WPh+gfMrzKcVQjir
bF0EjA3HFpmr+qViqeVSiqn5XW7xm5Cx58VD3P0Kzk+sEC0tOXRC6bW/wsM3jMTD8I4GzMN534kP
8830dysOWSnnl1O7yhGcqHzWc+GXq9MvGDLCOiGXvHSTZ+ny2rnHPJ8p9EmFphoJ38f+dBmdd8pf
ZbqAy30EbvYoBoZOdfhdwd1rYm77yyY8/8g9kWXbbeEdnnI7EEJtHRd1n9QbYYjuKNX2BSiBjvK8
3iDgoyyOLISu/eJNHpiLTF0np/2hdV39MG0spOTMqe8w6Q0kzDrbxbn/yWovWjiI538flwYuho8U
+mxaUfotgsia1qft2mcGHNLPy+N/fFAEgG2nSARMnbzPt2UcqM3x1g2kdQQlXqqylqFLao/z19Nc
8eijl41fEFLXoQfj1yKPyjkxUAXbUJJOyaRt4L1Ffek7p1ZTfZHnutX8iZO+IYPulwuo++7U6VR1
rmactcjdRwPyAVgzpCTbBvIFQCKQSWjRKnpkL/5dz/kinab8sllzbiJmz7v/5lOz67+BM0Bn9h+s
NA70mlwo4jIldD/nMFXzK9bW22hUScuw54yN6+Lh9S+uVRqzrgMzZkmzJQagT57JUt0ob5ADRmWD
pGxy1HvJbXn/V7VeJfD52ZMXV9Yb0q1GHz4Lc9SPkKI8bnOBq8xAfABc439LgmiKFTZWPI6tGm9D
FTXNPkCBDWPmT5QteBtJJ/rEMuTesJ5pAoOl0WRBEPY0jDkN6n+xeP6kW9cruaSWKkEdmjOQco+i
J7e+3Ex1b4VyQjWFDVJMXNfgOaDrr8e6aBEuF9PKKB3RtEWCjKrsCnubIsC3MMM5sPMs2uj4NIpk
GnK0g2gyMEvVk6BCOIuL0/uE5XjB9u4Hb/pcEatzhVYQjVo2hXeRhCQdDxiUjNQxQ7AL8VTTzQIA
EN+iN8hEaWoOO9nyAN0RT0AXeuzKko09HdMlhtExNykuyZ5mdugPaM/I0WjwbdETCv1WeCkVECBk
pfNtxVaLdYYhAYV+FRkuP0codjQEguC5ckkPS0Y++tUmumAtYrlSrNo5NWiQ7YkbuHuQbB3esaJU
FyjnxWWZQNFaBz3vZ+xXXBYjjkTyzmycNEulw7J4VFVwNazyB3Tf12mF6AN/CpZvLML73Qordh4R
CAkm0QP3ktEVrhx0EDL9ZsPUdf99e13mG0OrS8ew5WMS+x3s07YhpBygWMVhPWMyuzE3/AyPCMYm
c5n3v2/MvPNej1yEFRhbuz9WlcCzQjeJr8nsE2jCIZ7s4tRDFHTF+b79rctPySCjVjyM66iBit9s
Ilgk6Z0T+h119XRvy2vqFX+yEdPYscGWtcZLOVWgTWdX/qXqi6CnDEzvZ9WQYeGA4Cfz6kp+wAXg
1sKESJvFneJZabAzANQKL2dGNHOhDgX42bgqAbndqXozjQz02EcZadwXNEoj/qY70gIy7AE1vMdS
Qr+ORi5eNqQgxKv5WW+5mvcwhJge1WJQcR1o75ocvh39A6TT6/A4+35tT7SpZDPE8Rtpt3+rN+5A
uz686IM2Uq2PSM3UHNe0r0c8Ht7f63Le/gCSquS1YQ/zww9sFkaYSjdTYNl8z1jGbybWAoSh+DZ+
Jk9DWluwJ2aBddf5YZ+yb7aNmQN7R02+anYmFwdBRRm8xZnwELyfGkUk+QeFl4YjMm72U1RnMesn
QUqZwa9tZK1bu86JDLzjUJWoBLAwOjoDopGA7lLNb5RrT6pc80Rs+6L2qh5VVhg91QvkXb7FOV10
enKF+gCTEniLD7e2n0ShqQwlb78wBkcN27QDxheKSKCfQLdmH0xRhdQjVGDPOg0u02YkifijFxYp
jPfLVJFbBOwON3SwZaBs9LOkG1qAu67yzXjJK7O1LPTbPLqwNPkhMVcfNsgtOo7tai+8cZLO41Ce
HS8RJecrrAOq/3EZdaTsvADAqcRg5WtSHOHPeFEmx+L8Dm9H9zX/z06v3LDwgj70gLXjLtkPF3Gb
PQ+fsVXT0wW0H3NfASz6wyNasbKce3EL3XvlN1i74evW/2jv3L2KRRVPAJkOhYzGV1hHxxxS0N1F
io+e+I2xN/9/4KvqyPxu5Y8uXDB2ECxK/1svHo1ANmJn1sVy6VMlE35jQk3QF/ZuAOBH54W+LuJ3
Mklaysgnk7Iv4dsUHZp/h3s2vlLCMqYOjGymFxYBBNlNmGK8oyTdSA0FWT3kWXfWW+ocA/nDxoDR
Y76yCczPWzILfnXe7D/AgByuIwRhaIRQ5sg/7jhDQqtd7AmFp+PNDa91QvUCTgfIpWY09zfpGwnr
/pwNgfjOpXtAS8tjQEeQq2hqR/I+47zL0vZ2Yy0MZKefFgvQxzfdwK65f2n/byXabucH3c7NeH7B
tWO5f+6SYx18i0T7fYCQgHZpq+nMwGgxpsDPFbXF3ZtTuU+x/c9nWTP/nd1KPxdibz4E6T6EldLa
4h+kxb9XCsR+HPJYvEleQowgSr09F+M9StB5cz9aChoZt+L9mjHLtU0SYPXzV7uhj4Uk0usIDaur
sO4u0dCOZp/jBaZurk9pC4u34s3Kad2AOtBqQPRE2w==
`protect end_protected

