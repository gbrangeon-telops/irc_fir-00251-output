

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XHCjR0nUvMBgM1clzO9mSr8YEx9qhDtoXdaphp+J1JlsC9lSFtsV1/eTy/jaNsyBimTHmHB4CLra
VqfCr1I3uA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ebEJK3bmI2t+WsBGbhWIt2XB+F+QW56z7Xo7/vGiNjxPbaq48cjkY2KIIwhppzuYFDUdRDxp9Iva
RlWujqNPGUrxJ1F5Pa0zN6dEMkhKPrWWxZpAFto5e5cB6DM88tJus2O1hLy9PRfKWKn8u2fBqIhs
zvXwIEX3Rz7kU3GI+Wg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oZLpbXnbPC0EfiuqzOyPqmT4FdlvB20VtdO3P1fZux3uAWynrmGeEUk81RKG8dIjeHdSPnugG+6c
jKeGIJZZbH6MRScqnz2QBuupQkeYWE+dCLOq6/P5LV7F5481QZZ3bx28u0vHGlRYhLiMW8KnJ8Xs
JLZ2IP5YULE4cFTCCV3WAM+IdulnwSP3p8oyM0uQffeAJkOTKR9dl0lslKFBplzuTZ7EnXSmYYXA
x4iYEfwbmUZvdla6dJXCCjtKnKqL5vI4L1nHOaep2f0bW/K78py/TJVV+vsvE7+Fi81aNwDFBE3d
V+IzN5VNKD8wM+OpLL9AD+xsAbJ5JCLz2sqFWg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YaruXmtmo/2yQOaZLp6UQc/TTak5F2uchK3/c4SsORqNnQQMwFmjpORZM2++MrgqzkHH5KHH+0SE
PP+ha/JFKIuufLvaAIVDYgMKSDFaxIIvD/8aIAhw7TgTE10+TXTruuPFiw9U65VaBnD/nSEGkP+6
2M+aqBTG/2UNkEELi0I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SWJkuOmi8gVneMbAS0rfK4gI+24fr/0jQv+b5sUWbuvKyCco423EdTDwW7ROH+M/MaGP2QTzNz1B
sh1p0mypy290KKaGmvaZfJU7NOmSNGAsA7Eq3zQGPHDW45/4GXnri5xLLNnybO7r0Ndv34V/fxH0
f64f4NRroCys3EmRDJeCh0D+WDA98E/EHP+OtfmYOGeO+CDzxS2m3FIcGKs7pkeR5dgt+S6srqxz
96yb5/UwV2cpnC9ULYZHZVQa9WYc/XM+Dk71YUYpaEFd7osc9zT0azChQq+XAkJsqukhufRg3dQK
YVPZotO8blEly5GYlPFGnRW13eEh9DRYsb0pSQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13296)
`protect data_block
C/tAWEoeVgZfDeAl7TODgWX9ppodeT5fMBvL8hQOacTGPsXAjiOZgxRGlWzksmlb7jr284jkcafU
xoVOoyItDev8UsokBh2RnlMgE1vR2OQd7mYEeWocKP49HZJHJo7L9vBfs0nnWnPo5a4ibx9Y9caq
Jqf0/VYLj2k3q8Rlx0RQfG7GHeyUsjQ+8bNXzhKDwbbmUkNgDFVnK1tFlyWI4JpC+XZ2CcR5jVjY
T9RX1OgBMzON0bRpkADy+aic+tL6Moa1LAuiiBMf+6kH9nuHD5RSYdG15KuCzpLXVTmDFffN6lwM
MI4ejMLmJ75CJvJLPJnYob8+WiCTTt2mCEq+OZJ8hCO2PQyMjYG8a28kZtdpiSCcErvj2IU3RtZB
+W888E2xdHX+tofQ4NGgNyxImzdS7jz3uiZIOW3yCk37TIXqmyYF1JX7389cChOF34MuiMjiSc9N
TcMpqaUWevtNO5GYfkCOOEq0p0leuO/BVSWWy/HwlyyWBBojcFUqRuGkOTahHbLZrK0sKZ8WDGP/
7PJItTAwtgChofboLIV39u2wYsFapBPHcYel75U7e0GjsP0jpqQYQzuGjmZY+HxU14RZTYRspG2g
gT7C09cB80IxD1kqppbza9Ht8hm+Drf9s/efOIGUSa5VDp6bOvNqxNFLYr/HGvSQQwMwxzTLu0uY
oRh2z0SHmRYYn7bMRQJoJi/VfE0jCNmNvZDS2anLtend8F+CnJvyjGsaJLw3mjAA2MrIZxv7UNWP
0c7WKqCGdT4owXSINW1JgHJHO1PsyKm/S2OI9IyDqY28SiUpAz0yrlGCRkjU2c7s6wOhT65pDH+A
YZYsjsOuP1DtUhP6loUqzjFm7uVRQpIuK2pGQbGV5ZI+xyh08pu/hAjxnbrvuMGE0NEyCHrsG0fY
QVjLKZYOfzcO0blHb2hkM3MieRh++EjyHF6qfQpS3eObL5/eBMfVbxy8WXcA+0taSmCK4STHtaeA
amb8vm9PlFe+D9kH7uzEjTxhlw7PlqISLHUgxwi07YV4jPGvg3aqu48gTGBOBYWMJ3AnNmQHywRn
9sd7BJJPWwogNdaK6A7Hb/iCpyzUaGxv2BGS42e77RcczV3SoXfwAR13irg004IxVcQooMxLPZrc
I5PrhGAbn2kMAYr4BDNJRokmuVKiahzkJDGj+X//kDZbtdEGNg6plsXVNEHAr0+pVZFuK9lufnyG
r9mcvl6DP6rlj/X0TieRukMKHnvqFw8yE8hbE3kVKYR6W6I6udYAuzBdCLjzDAjas50/Ja7SVcOA
gOldpT0pOPzcKfoHCIKT1E+X9wG06Zq/DO5jsS8ttAcNL80W7Z03nq+8qrTprBaYK1G3mtoEmdIw
oRHBPEqfL1HnA7xIalijmKoIlUe/rel7AK35RNWoRUh+ZyHq9XfJZTGy/1o+jm/PSjDdFA/M0HeG
wTGNqx/0uHWXDr7kXCYk3RWR6axB/l3PxPqVMd/69XHlKjlgZCeG2B78iAUv88wIedvUHkPZrPuw
GJ0xLGnBWj/9zgcCfLxol9Gk/9IHO0OuS64wAtVgWu+f4Swj7LrlCMUV3BFq4Iz86QsoykdLKRyu
SOWQoB6lsbAr/VuFRRugtGgbiE4hLS34B6/Ml1rrYt8Xc/z9u4P5Tnq6wa+yNAa85PKQzmrNkqiU
Y8ilqoiyMRrTpUwsWTqgyAVDTysaPUFqZhT1MwVO3/l1EOx512wWJU4JXFQNTl81Fj3R6mV2ORGk
fJu3f+kpQizlBXiiB2Z5GmJC9831fKS5Iw+N0LW9xK7AtadCdgObyGRrUFIkmsJ60yXhF5AQ9R6+
eQtgn9CbjEEsm4yqnRx9u+OYoY0Z5NRtUtTxZO7cDmBoejJQKmlPdeXgXKHKXJYAF2g9cZ0q9fX0
2lqTrifPitH2EqaETGnCwIKPeojJdbZ0cTBAuPnNPV8KvaotCXwRkXW7mBCODzR1C5LHlqCpwZfd
IxkyitjMq4yjFQO2HZpHpcGGez3/awmqWKtGwzl7bLct6W8kvv73fo+unq5xY2XbCKIIENAI9XDs
9lNzgrLymRVlhFIiV4dI8v7amHvlOOyUwnCahrLsi7XMxFatS6RtCzOEPDHu4Tlh6fP5I5NsOabo
WNwIxnpb9OeguG+xy+10JWIOR+Lpyq8V5Vkqg+D6tRPXWHlzIO4okufrLSMu01kHwtaM7o073Z6+
ZsgubtRpJABe1ht8eBvVapN3+OAhsd4dVBRFirmbkOVHmO3xvbuG7RpA60iW0R2NESm4gax1XcNU
LcmWH9SPAv3ca59IxeUOj9V5VVqlHA7TlH15TIXDpQ9pTMqINL3D0wUSXCg+1vfVYJGA5QiB5p9U
pT1SYS1wVhaX25WZQSD60GWmBqcdk6Cg1KbLAsbgjQLYlK7bUKbXniSe4wqLe9bdJcqqgMpW1JGz
vfn019yJVJHEVPvNbPCdahNiqaYyw2OPBSZw10Y7OTm3y0HNGj8kpgo7T+1NsAIbwzvvECyDWYki
FvdBSC9VqrmBkt391UcVUh9TK95JMzfmjeSjw8t7qSDpRvd+xSNP/iVIo+cjRZMD1qDpi6cMyrby
8FiofPRtza1qMaduBEVSrlMhK52Wo47xcjNFGBEgPlpzdXhYVKarhiJzalPoU2+U+xQwZ2gs280x
l77PP3Ig3WLhwoSMV1LRtFfijgPJx4CgDArrDfn/eKf+5y/1HfBMW3a/DH/c38YLRO2TPxsZB88u
NBJdARIgT45ddDofuDvMLJrG8PzFb1zM9HFTDWH3EcHajQwrRuITHleCEKrVzjaFpkFpVvEHxCT8
y9Rt7HB2UOMliMroy0XfItWUDmymkTN37jJyzA6iF8TeEZDrJ79QfuhWI/l/Y0nd0dMNrxDsIABg
pViBJeCxeVHicNG5ygNA7VyU4Jwmj9SqcnsGBOGRfKKnoGRI1pp5z7lTQuroH49+9OjgVT1j/K3C
HgtDjwxCzvQ+tKT5BiOOBaQtFMFYMs6wE5CJEc69EHgDB4krbiYKnY6gborH3gTYPSUMZmtTUnMy
SrIrk86t3sFhEvdLaqu5gwjyDHUMFGbJ9vFdE3VKezSMFcwZgVKCKeQAXUcNnfBbnDicSNHvMWZV
4p9ppHLJb+cnOx3h0fwIS/gc2u/XZHfLfT8cQUl6eXPHIJ5aA4addWROMf6flD3dOo0BxaCrfgkE
VYSJwoDVEZoV/9/zfBLQvhVN/jz4VWD/5dIyF5nDNv1YnzZKzT0DbRyRhtk3HZwngS2tmAe358I+
a+e95iZ562QGiutdlBb3rwsq0aSl4Hbmxc+Tk8ijwGFE/a5TFDvfg+0/X7icCIlR9LHaiL/Kq6Qr
rC0BUcOpGrFyYDJU/fDEogtet2Z2/Zz9xgmmCLOJ941i5zCwnq3607u74FQBSFytjr7lJttHqyVh
KyueE/1LoL5JM9YF0Itl40f8bUg3J0FqXdym+wMLI93yWu1ks5f/RiFL3ClQIlhwQO7oY1FxyB1S
xaDW6PmF5LLoHUw2Tz1t4Wk8RoItPoZvj5Jv7Oldsy0HzJJfsRLyy/BKh0ktlYkoGV2XnwD+BcqX
5rgZvda9S4yULKzDO+E7luYq8dPzLCXiiy6p5x0ptUcmj334qXqjFRFMxjD1DZ0qxnZ49ichhcBg
4l7v2F/bC/zUpeWZeaIPv6eSChl5vzBKNuU3C2mWTZnAiwNQV3Hg2cti/7w5GE1uz1FPYf2Le/Lt
sDlwvuVxLH+WHNxuafJTYDfC5Sw/poIOKKJfmklD1lxxTRxizLKWtFrYsOBUlbN60GFmHrJu2lNS
j5T535bGPgyVaVufbt82CISw+ZCYyT6TBh6bzlzz5oBltfMAzNyABsx+BH8vVp2uQuBCtLUwnmkn
S0b0cnyF/oAQG2uNPCXBiKyjSWNllLDTF7bmf4qKGsIA4z7O9tz/qZBNJngO7JxzV5lp4vsokWBi
cmEIrTXgGHVoiD76aFgE4y1SjpIhAOqAkKXkHNpywY8bq3igFktm3yzWjM1I45/xomTP80YcdPhx
YpHYE628sffNEwYLaGGIEBxKO4J38N6gg2innDGsNCkGzX220XoGyGOYnkv7DQWtMvkG68qjWeyQ
jeAhHJAHSPWUwabIiY5XZVi7uqlYx4tGfdgVksPQHoTUZjPJu255jBdgfwlLYCZ2ZdUaOlWdgeYV
MFW7FqLB0pa861g/+kYkcw7/o8Mr/7VKOfsV4SFEUJMvvfPHJItveaAz1J5oGHInuwA67XnjhTGp
cG0+/7N0WU1GfC7YG9pYiqWrksE+yQTdTrVZWqSen8TlbiawTtmVuMUE4lWXu72DUBREjwV8xUyk
+ieoulM7HehXK27fQFc2fEZQmStkhgKdr2JTd5uLhFPexpMqSxZ3xLS1Kfq1TALTMgNXwg6y8GVa
hi8D8905ANNB844FCa7+nI0WS4jTPut4Yb3KKNTAxQ0enmCpjHF1A0sye8qw3FZJlXiPXsbUX/fL
bbNau7b9jAGzCC+7m+nlCrGxh9pCeyNaDWdKzhVD6f3spdMpSVB3dU5O94HXf/CWmu+cZnikcSyS
IcQVs/x5tZsjwenDRuxFV8N1iuzcDUStxj/+HDkqRnxass0CrR+RQvV+Fvb6zb1Fk7nfQ/3EIKhX
EN8TmsMs5Rr/XnPsZOn/ahF7D+WovNgAfdNLtTxKIfUMGegkGP4e5ybonGcgiJVntHjRdnFTWZos
JNKGdsvRuhKUM49yxHxuo5PJl+lRhs2DWVk99SLLZ06ojUtk3ZB6Me1fF7YkPMuAHcN7N1arBSnH
s5qz1GWAi/rUKFD0BzwsJk1eORIZtBuUoeQdJxj7eN86NLjVU86VsryFHhxpEcc/p+8r2dzyhGn6
smCqqTCMMsp6rxP14O9LzvRf54o0UGzthOPaNcjJohbFRSwxCRMpQBGlxRT52ghs69hx8OD/HF1G
ebyz9zpWt6x0RkkUb2kxaS1BfOc2rsRLA4jDVQ62vEZvaWF07r8eKa8Vj4tZN8hVskdR4xEwhI07
Uq/hNPAkLHwLIchUQsWrROPttqGR2BpWbfamvqKqgc1h7bNSk+tuLKJ0ZNRNsH+Wp3Kcj/v5+D7w
HN3YZYBcIPAmn3aKOTcwUrZi03qz5b5bReQAw73XA/fdMGNYMSuhkZe3R4Dl5KliIewgSSPByx/7
a0F/HoR6ovr5zq3oQ68c9fOGeu9tjZkbnogLMnrbqemT9lNFTmBRSQrO8TKI94W9O0TH5ihHCxNv
Gnh6cthO+pFtpZHGBBU2MWkqDFN88uVs50FRnQyO5UlWSHz4QzoyiXfcjmTZ/bZq5bSZBWqEGaj4
xP8BQZsE+xAxfUq1HDPSXntatm6O/x2a/HtRTkGwwE4TJrTPIhyhhoIrxkCyp6gpZ4ZfU/8pQRgb
NZfMv+Xe9EiAF3kSifDX+AqBgI5zCSsROuCviPjooXxXofykmy5Ne8OwPTOEZn0i0gTsPxihS7Cs
Mci2ZTYPJOWxW3CFdf+cpQiRdUkDeogV9+pmllPuw7T1j5gjlWYTHia2uktniNCTaCkARqXStZC6
wDbLRFyC9SykF/jkEAMIkCGkypdgZaH7vjyuOJ3exiR2i7zfZ7aPfvDD8G8q0V4UtAvPEtZ/unPF
p+wDMAbn7ge9AI8ufmFiey8sQ/kQY1hbFnG88oDG9laAtqh218g3V6fGO7fgmzexTE6E9kUwJLp1
PKu7pAWeaik+78ghrzj2z43fZMeIUrkNHcjjtWMgOUYPEFDXfRNVLOTVbnq4lAwgPkE+oy5P6wob
t7Bp8AWoINz6jJJU7BWZ7yo9hFD81ClpyJ7CtA9xzfuKecGyHbU9FHdKlFhuPIlRUj2odYFsHiOm
WcW92RBcAV0nyVwQXxKpyhOwNVYumQEitdUVIcfnkq4+jCTfFrbOhTyc1FpS9Czo4RzCeaPXUpAP
yLQcmQH961gPkekqo4BRK9q7dRX0B9e4eiMF63iSorLJttm/o0SlLlt9E1d5qG7YdaQVMLYaQQgf
nMnZapp6UcxgZ4db7EJcIkn4jbFNLRQMLdpvENStAsw6IT+94Sn2wlr/HKEeirK7ny7sMRenh1Ix
Amg+jaZ2EpoAtljp+FShMrGnEijFpfezd25PUtfB9p08OUhnYZagPsxBI7z9I3TGlHvwoPWCSKox
mw+li41vJIDqqBD2nBM0Zfkjg5X0s3OOEwgVTNTHkGRN9Bpqcydeq4B3TnRNIaiUTVNFASDDX+gg
xkFha0JEpRYdY/F/7Mv3nTyjTA3geCX4iH9wrjgaPT9d6B3URTcL9u+FiDs9mNqR1M7TNX5qH4To
Myi2HBMnlN9R9U+62wOU3IMOZkof2A0b/DytkYOKD5+IcVLatJLsIsyoIWeAgXdY89ySANAy9qrg
ksLjJ9Ql562olTQcLpIeGo00+8zE4Zf2XG0WkvNLw1yLHcq52cf69Y4pwkO84pgePAELrTuJJUxa
3N5vgTFOT3Bg0h4oPL1CKK1Om9YiFqNUAdRLfc/mQLeMem62hPgAMBPWssKp0lNKkjog1Acca9J5
Hb8JQW/BxhAX3XEW//x9PGxUGUdS28POfES4sJDAMNX/uO0NWv4liV9Jho+XKTNRj4EAlQAABEa3
WoltpSWIL+CXhB54hH9qOq0mO+6DfSA4r9+nyY1Z14kJ/xI4+3uZazAB4jyCZFrCdzczjRy53kxJ
rIQlLtqdoXBNh2UDhnEh+pFnp8WxR/PlIYFr4yQJ3PqpJbXjkuDqMvEUCB8fhg3b7M2UWuXxK/R1
/d8vYUa4JwyqXLLHr3p5LTA5F5sbc4+VTLU0/unJzPkpGCEI3ycyLoMrRM4dZaKlpBQV2tEGZu61
l5pH2glB/slLO2mMGytVr44NOh/S42/EPX3E079+qZFhoKduEbTN2/znr5rzdDn+6vdCvJjldYp1
SyvPLgp2tPBESe6UBzJUHI6YUUmgsSabnpPmofO1FV55B4xEq8gc38/y/6kIiW3jmeb4B57TxGGR
85nDtTTOml5Mo2aQCM7m6e83jif4RL+bWkrDKL0iPWWDs66cMprejwAs9DnZN57B5kwObAvTtYaB
AG5DeN/vCmVJlb4GwNUlKHes/8a+nYRoe+QxBkkAccRqEozwSThm+w/p7FADRAdQ3yxgDHw4BHfd
psnXHKPaQFvN7hyNoxB9OcDSkOOarS6+ULPG9zYMaQQWJaxlkk/7gSXPwLR1SE2Q0erjQ7y3AaWY
SBh3YZ/JwNWrdk0aUGObuQmDFll777WeILchyjfW5M41AUW9TL39tm9sOcqBh9SfrR09wVGoamJD
Hxi3AZS8j5k1ROdfYwwFjq4QfQrLbup362JXuxK4wk7AsEFd8fvnx1Q8x22JQ59e1w2+p8NyHady
KkN3Jsbh0wen9t9M/za+56QvAv2PkeSteooVGNS5AUHXB81kv0Xe6feGHYWyWjTjMCGuZuu7RK4g
CQ/nQn3uzd/kW15S2UDOvkKA8cCsNfiZz2lQG+jLeVPCaRuBGEKnjKySoFZBOoQNaK8jufTLkMnT
+0BtwJRnswJgZTQjlQczkF5WERYd10cG3WELHbDm6GjC0Ftp26E78PlHYCEkKQNpa00cDiVuZyXz
FKBsWWpmG4KKDJciF4oGqK3B6LDVlKEBTBtODbFMfRJXuFjXrIXUjEW/45dsyq8JbaI2+s7fWETv
gj9252CtGa+s38NwSijyLJdVVJerIGAwYpuIClmrYx+r01TuadOkjEHNz3kFbh/pUs4WZdnLlUtG
SyD5kLyRvBCqfnUx56bTaOsSamMBaMBCer+BmRdYoJlmIeEmm/SRfwPr8Kz15u8wqB2S3kJjkib5
r73V2Cl5mZuH9+h3BM04p2x/uE/siD+pH+mQVPgBM2zYLjz3Fk+t1rOfjxggadIkWC1hu0GPZQ8/
fbwM1qFh0N5YLHxuWQe2J36nXJvH/kwjVGMi/QR2cGMno57XNO/VQWzEaKCNvuPbOhTeqr49TFsC
pzS35JZNqIU32Z02k1Yazn4NLOBDcv7yN15348x5zWWXINbkoznD5jv+KmJMSGP7gsp/drMu3fa2
VM95VCytQ/9ENe54P+QW23fQG7ZdLMLGJaryBnPEQzLKQMj2cBK+4T3MANANz/sCE/mCxu9WsuYD
wlVpfLQG+QHjXg3doTeoU8z08ck2bACIKqjAoZor34vKznLYKwqjTagXBvJEvJ3xCmFd4M6uGok0
C2hR7/xzbpdaBwmvFcBVkn5IBL2DAUayRraD8RG4gotW2twrXcLbhrrr3HvjGxE43UrXLGEufVQs
/FoBaBwxhFvXiq4CA7Ix9S+/BsM3rie5Hc5ZQERt+btbK6xzx1sSDxTWRm7b7rKlhpN3qkz2zeCF
yzd2T3Vl0d904c6yf9Tg3bA/U4w+2w38gMjTj62AAm3O7f7ZWnq74ZzLYm3AEOn4/Sa07xIU+730
qmrm8Q9dWLU9k9O2xMqdSW2j3oq/YaOtTqz5YwOwFH88dcvRCuWtfFk7TY5keVlam6LBvs5BTgMl
oe71K9Gd2RIRfTftCtGVQW17t/iQFGttoMuc/hGoqfDAguEythwNdg5lZNxprrT55Kg2kEGJtzbM
Vxm6MBzkaAhAUFtx6UTiov9QS8/EhK1linCmVYIMV+ZpGQ77EdgJRjPmINPV3wI+xCPwpcXXqJZa
DYyVisAqvHGTGhhz0ZhmhdGKrpKei5lZaIWJ++M4HPuQ3ZvO8u5g/H+O4Q7vumAZrCP0LsNSON97
+gR9t8wGPdID16q4SFTqupFhO6aHVckB+n28Ge0yxOo12x7OpMe02yd2GyGvPUALd6sswr6uaUSa
Xb0v8h9EGGazUXHq7Bn/fnK8XlqNPMAAE6isdryB9+6XsBYY0zibDY5EMy7jYYSditx3Ri3aNpQG
H7NdILE7VE78pSIx5RrXm5FCRPvOlfNhO0mG9CZov9reYWHyomi81kcQSF42omtVfxEXgNH5XBZ5
P+AjqcqIvMe66BO7FzA2QE0XXVttBWIlzvqJMkbMJ3daerYoIV5HkI0lRTvN9Vdfd8agY/ki1UqF
vH2VH5A7ONYWcNEcbCsbgT7mzRL5vZErqay3HLL1i1FXcGEDkUG0p9JVA3sBka6pqv8uLcaF7ODG
U/jiS7Doo/2UUVqC5ZKM1qKRISTc9orGjtFcSIkjUxgdGLJ9vcuoLaQk53blFaPt95URSmOL+7J+
AK+v1W+Af2If4wRR12NEIXwfyA7MgpMVDQLCruymGpHmHO5KG+UDmOCsB9XHKqAdnUM2qOS1p0VC
eFSmlF9egK/Yw9FvmIeJWKP7s70G7YdRx1if0r1NSg5DxYH1D+rqFi8yno3uoSQFlH2YScNcLS5h
vn8blPegWKxEk1nf5vp8XPRu+bBnEHPvz3kn1zisI2h03zRBAWNUQp15uuLnQPcKzf35aa11QmFF
vNqdmPGAfrdIsFSy4Rc65oPPvPO0HnLPE+gV4oT0sIfslZ/J1+M5swe/APblyfF/nbzGjpwyfGyR
kkNLQp3i3UiXytB5rGOyznsvOp13Gk5s1zAPB8K5/C58jutW8CrEwEhjuN26tWB5fXrYiVUk5XqH
Tvh4unaJ7WrPDk4sbKw8WgUktuu1C+L3Zquc62VpyHbL3/jS7WncWHwPZdfIaDHc3pz/1CQ5oG6N
rm1up8G4WA2K/1eBqKAL0IYc7DkvEpfb7gdhuaGmJ4tpbzs4akFg/DvESTid0P/PvpAoOUyK1jwz
/IYNKukrQXHvSjmYh5HNYqJc4dOcvhcNdbKB56dtFJlsk/y5mB0iOu02CjguJWt4xkcoHG7Eg9/i
hKm+GqO5g+tGiZT5/8RR0pZyeuBRY6dx+tkf4xAbynnykkInvs3GS05/OKktrmlHRyP0pfmL+xHj
6AipUQfgJ0KHPoMZHP9gBwba5qAuC5/ZfAszhm+Ct1veyHclKQYHeXCev5a5JR7Wj8GM/MZw6pce
f60wWiWWb255iu4rMXcIhptd5Rf4GHdHScyJ78VPCIBBYz+tda179nNCB5L+DHgF86OKtafkPV8I
PNytpn+6q900HVlG7g+8YkrKdbvo//hzOtNB2cvsItybjtHw9BlkBCirjDtZmNpRysF6KfyZ6RVw
YaK57scpt8bYNB/jADgL9DNPdLt3GUz6FZzmn6f6GNnjJivUlL3HHHIQz4UjUMLSovrIx6Cb4D4u
vQk8Bv7HQghjrTBp6UzORegFiJrHmuPGxAlDmwFEk0iSQaWwUH7T+cMkqZmBDr/0aEUOUh0UaJAm
xPTFRR8oZvyqw3hf24NcQz79Up0kJm2U67DiR2hcM+hxk2Ou6BrufwicWMgzBj6xXgHrFajkDkFJ
qbPI/QJ6hPTVVSzH8ar0J2N5U1VuxLdFcSCYlNMe1KOAcHSHO8vSqWYp80gURwIpd+wo/eBSmxvK
6WouIKwMt1S6CoQpdAEza5s5lbO/eGfB778GFVTWTY0Ag4K3zUaROX8a/VznlrhIwM7VC7tjdVSk
Cy9xbRR0MWyBT1ylTqs0kvL+XOP7EfyrIc3O2o7sj8KSMa8/FW6EtQIOtPGkZ47osr+NU2a46oLr
On2gkiE+4x++KoHLF5A7HzsVC4ZM3tenonCnE3ERdH51+AtGy64eusSBxqmftWGO/oc+QUPwLkpo
qwOPzNBxcGbkUWNi5ltLkjmuvC1rFVFmSZbrocS9xKdGL5e732cbGYR457qrJ03RH3r+b/IboMZe
u0AacbZg2HPzssbaTRR0LJV1mQ7BtwPNcts4NwhqI/VteW/Y1Iig0D7fTK6lsm5zO4PS98HgQWJP
ATs1qViwASzjfpd2AVwkM0qbd+7Op+i1OM89lfCgx/oOseMqSbzHQLEg/GJBWoaXc74FWF2BYB3r
+eu6VQg3yU4n90vT8dmwZPfJNb4EqmKTmME/kq98zHFDMibjRkC5DbdRYMj/sh1Lv4oCNEEJQfQZ
EOCtv3nguCGK+sbxIDYBeMR+wrxA9v8390LLRoym/niBeO1Dd0WWoG1YF/dO/7NWsKcS0w6dKQHn
qAiAu42TlFt+K+MyGQQcVaM33mt1paJbnBQ709a89NXmCn3s6ymrQYsFuXn6APlfj3OKDzDqZfBF
cPVBpsYCgNEm93W9TE/kDrwNn7l1lecbYnU827Pr9XDAirk6PMVNNvY3Is6p/dUcm5NyGTX6cGO2
KBC6tjWNMFlH/5puBApCMRTk+qjBbF2MN74itf63eSDLYxeb59pg+6zWZn9pr+U2HB6RY2eooblz
5XpGBopkeITViQEzNFfD96PBi2CZ3WqB25Dp+f32y8A/EUkmh4ikLgJD+TxZMJXxSITZ8qchNL8/
sbG2AVQ82igeSat4p1GzrDW83hbzDUbJF3/mkiCnB7DZEFDJYT++jyGfi/wossz8dmKerMuIhFvI
zTEaFhv6rjI/iKpqUX4in8sidgSDv/DAOCaEU0JMldC6LpVwn+rh8DGiOtGvjCcbXBhFK+2YgV5i
XVa96JYRL5UKyqyGxlzNIVAWno7G3PeMUi72ghsj5gYvBui2gLY39H9+xjDx3gCMrP0LygF6YrAE
KM6MjNC/KWHuMCO3p9TIa06fGFw/MIf4C25SBOZVWt4DVSxglUoSyJltstP693pG5BN8k4h4Mgao
ZuiRwGQ682ypC4ADnHegWPJ+h8ylfqYiN5VooDSO4ZWlslZhDaB9CBOOhsMwJRd07BBZAIfM4AYu
rP3neUcOaFQ4i2Mzm9TAv8Gm9clrJGirVSPaOchzPL0hhBEZzpSmZKrsDrpuNxavowAe6BDzFYuj
BYdMj1eU1DFkWHOeE5aT83LMB4UJHDPPyJ8F65/fl0WkVTCWNpy5m179sNXdqm0OlMLupTtccz/n
5M8ntbzPAAn7NIBkwUlPT8HSDjAutunikXUHHErvAfLdhl8zMPYKM9yB40JTTetRvShP+VEfj6wK
ZVEEUZC3O3fEoZ82tz7EzH7NkPjSZgVeImBNic39D8AwkPP2Agw8Uxnr1mvPSf1c52wS4oz/Pj3X
SzLf7khdyHoCBVW+rav99pO+asecb87wPiufPAubYb48csU0ewt66i17pYl9QyB0FlRA8+rq+IcY
MNhK9tBjQLUddrWUTq6hvW9Ax6BnZ9ScQIvFq2rmff+SG+jzuhGOC1Kbc2WwEzRtYwaDFNABg6aI
KyJOVMkklTy6VXM/uV+5+kN4H26+SgDaTHd2obd7onth0sUqepoiji6FLmNBlSNxOXqEsZvB7tUz
9kNqIHBekoHjt7bite4uY13yH+Un+C6bBi76F+6206VpiqMUZILckb2vn8LJzWVk+tr2uwyN1W4a
eUfWmJKrrpXgRFCXwCw10wN99R0TcLSnslE4J1G2E/WKKfo8Xf8V/FoPw1tcxBER4/UYszi35Byw
5F8EKocuWY8NtOSgxtM1SoOXTtMBFfU7G5zL2mxYUr+um9cnsfXsykSPm/0DimWU/b9RM6H3Cs4p
4elqd+Sn3JIrSheBoC1FSNX44USjcVKTBEBspYZHG7IaLDR9WnB73DU8pxHvgjWJ7bZUdGWO6jLI
dOYWk0wUkU22Rp0YHBETmWwZkKtYrizdlhOq8kcEk1/CLD+Dm99J4VjRgNCLJmT2j68nPswCMw79
QeTWMA9siPyqPDQsOS00cUTO8tHmkBoGVvBzvuuaMUDSwT0UmNhy3oPoNTROGqm1S+69mODihA5Q
dpzsxiQ+HPOUW5n55N1wfXnNG3f4//PH5TxqqFozyE5/bZ8JjLjaoYP/4/gewJ5LhbIRtlFH/A3w
c7eDbmOdF7cow1qd14rHwFv/dOKErYFy4TmRxHnWMkupbNiP1aT2tw5dRNUxdxLCrOa2Lmn4Jl+1
rl1ja/PK/HkKIbko189OXjoU8wr7fvMpDvOlBcq5jocK4mKbNNIXbx1eBXD17l9plX+0txHYywna
kyCu5MgLlIlFPXia46JcyeT3fZNuhTMLz/mZN+B+n1TkbpYlmHkalAwI4FE+2mXisGAaryho7o+C
ca6lf4Qj3NOeY99o+4IdyrPntxt2muyFqhh0LFRbbwCV0clRo5IANsj7xmHhIzCcn15zeajM9ZCS
XBhYVdVQMWscyhM5QrcGee/pUkw950IviSn00tJGqMCYB6u5cpx3LIRG2hbJcSXswYhP0O/fExz3
TmLNnL3EAtj2UAbpGlEQx3kq9IH+38qcc73rgzfivSTQZWGo3U3ADgGRF7hx3flmLn8ubKN4TM9u
470dlNOTuWsYtPQdyn1flfqUkgfWSNMyZ47PI7pN4OEmub/DyhOtZaLoSUsi3JhYh/u1iTIn56cS
x3925Azc7kevmoILUs8TUTh626Z31eoztNF90Aato9h9KXKOFQpCIGFb+uWDybst1fieoOCVQoWK
8Lhk3C7B1z9Fk6caUIhHY7sV7FqjU3bj0C4X0wwf0LsiAjV26kvKQ6NRN+utsmKSAXL6zbT3X2Ji
FebN5wvgT4hYtBfFcTuL6D6yoR0zyz9Pbj+zYncUGuSyLYddLJgO7lRDt0V7GtTJTgGBBw+Lxb7K
yT9+yTGlI0H8cBkOu0itrRYGd5oTF4aODUAgC0f2nxPCQC88r9kxhdw7SpgZEYgeGz4Ru2YBYw8u
+1ZsksF3qutzZgW/YI+6j+UQ9tepa7XJQF/ohNwdfBkQCx04EnhQNjLzPc///DNygjONSVh45I9r
vNVkU6k9AipvpMpbYFaDVysJpEv+fxE9RiHtpFsl3hzV9/IklfusNBMyXmotTRRE83yQvD633mW+
ycFwTalgXUI291QxR+YWu6n8kBkWkpCELBhiTZjJN++SxGtGyrxt477gDn40OAsNI8j+VJJIS43G
qNtUe3bAK0mK67/g4hsH1IlJeXVRu0V+Yr2BaHt8z4Lq9c90nVmb68arNHJA9EaZNdl8plRhWLsH
k9nFBzElMJpIZD2zvQqL9AZPJqcpOIZ4Uz0/+rR2F8v5YgjpgiWFrdGFshUVvaUmriGGXjKOGbh+
N1RGpfVWu8c0h2lEbWPMYU0JTlR5qfp5kNm8+ls0/Wn85WTqY1w09dp8BWbErAnIpIrhDoS0FukS
T5qDOpSuYgtYruvoG/NzYjFxD05B+3Yl4tLzjsEGuXchQv/OqXFl90twqKQcHr+ntjYfcYCiqtWr
i1qX3ao7hMX7CLn2e3z0xe/MSf55l9aweGC4BfZ6NN45ongqp8P8/coTN6rKDGvwk6fZ2ovSqtYA
gtIRznQGYQRp61E3V3rnvF6rU3bRmCm8O1nG1Dv1jx3NL1zxddw0i4R3HnBFxFhcrdc0KRiLCg8U
iFVUPWRlOgn+pi3Hbzi+241jTJaeCOEDR4PV/uG5uZHY37Lp8KbZvrtJzY4hUnzl7Hm8ihmQKEVv
nCMIoEAwDTqTHg/HDxiWHeVghAbRYByPFYPaBYqmMo8PhMCZIYbvmumSSKRLyJSrYzrIrSDuHI9V
I1soQ5WzDnBGd4CJfxtTF+B1eVJh+qDBatilKjPv6gP0plQoE32TLeiWVHVNUYeKDrdAxeFhpcm5
SqJelpmaliYydrsX5j6Pv+ATodUfUFOO2042jnGpVNkvP4Z5aVouuBsC6QO5JSFS97A6UjNPY7LE
OeNtrMN7b802oPnzUK29ZuKJFnlXwvPtvNquSI7Y28+Q1mTZnnaJWQlwuYy8wy5rVJqEqzIEyOZH
6v2yWBKaghsbfhZFgte9nJ1GcBxYVLL8TJXlCeM07K8Cxhxj4SdxtYnat+XxBfxT3Bpo8L3+ZTG3
gMrmdhp9ystIa4KfNNcPytCLhQhO3/iFQsqw9SQjgbLnqmFrAI9sjjBemdPIaq/V/mxbAIwVypob
gkS0n3R6KEUvTGdo4l/X8fBTeNOG+ve8qbAD35wJU4RzgIcf2+xSV3dsNAkmk4wZfmQVIImq8VCf
iHBRnJItt1PZjivpY9JQgRnWOcOKGm39ducNSXPlrvsI30l8JRoWT4nBuFwitGLkQa4rrdFjsUu1
+wWxbz1xwPKAPVGCBW36jKLe5cbluZ+sDUv5F+Z3ootRBlLOOyvV+5UrZK/GjSlQQC9nksIhJ2iG
PTAnDSrq9roo29N01TXMt4Zm6qjnvgs3v+Jm3YB6u5KClUESbb9hwMItoYTxWgLU0mrTuzcuJh2y
CxHji4JW0uIQ/++msc9Jd3v60oMze9+MReVCPMViGfSCGe6kLmlQZoEbopEsOSnvFZhITqYFoesV
+2bMQvztvKofWe5QY5hHVFgqOmFhf1UGGSKAmwE6ZXc1dKdrarpPgznl0O6jg3G0eyzkSODapSnF
HWMrSG+0Z2gmIfB0XqKPLezCOc/XkqSDbdN+m902hcY8a0frBZbiOAXkC0UvHHFnRMBqTAuWr9kI
9iaBxcZGN+bnE/70B/s+oA9wDm9GsSPAxwaK3KrUVBwnDUXSbpUTAcXjM9Yu/XqlBIXrdPLCgo+x
5EOww8sDq6fysIjUUbK5MXd7F0AwVJ3ZbUrcXnGzqC9qA5c0xAC18bPeC6ONy7hnZTaTJAhqdyL1
Gjr5WTrX+HVQv/bfq3oRxZhssB6/qljpX3zxqh/Bt+OpEtljiWzGk6vpUZR+EzQ5CWWJIVsLRABX
A4DK6HDgdBpSyhpY742DjbTLXTC+De07xL7rJjcgABBBQKItHLeaSWYM33ebJW8CkmiJvHmRgRfy
A39ZrDEn764dZE8rxqXK2wfGab3+cEGosiBzfAxtL511EBOvLKmFMH9DYqk0M+29Lv6eDseRIedq
yfbMdDD286yTSp3ziM3hHZ4fXOFW1FvnHcbm4MXV6EpSFP4mR0mjF0s/aG3DY9w/K59Poy9+2U4t
yomBvUPH0uVWnpN57trGH02k7563qgZ5rmrxcSxQ1wnPC4LqktDL0dSPwcyp8ocSaXbMR/ajM43s
51aHRMZAQp7M5OrK5dGAYlc/2PAPLsmwKgH3PYXiZNVLto13IhUfxdD/aAksaHQDOmuZ/uOEkyju
3Hf+gx53Qoe9IN6nwlbfwi2iwciqzCufLv9s/zSOwS69W927+31N9Ec5K1iEFUXiuNq6j2dong2w
vPPeCfyYpIYapWzPN0WuiBArpeRyMt9NjCcUV7gzyR19ylVPYMcgQp0cfvH4aOH5CENal6MvbvqK
y8xg+eZ3Sd8N9gyzOadvqHs63ADizYDfEXqaworcMPqaqYuo33yf2I8ljxz7tWAgJUMccwvAQXzD
5ZtMT+PrWhH4bewyOIrY3Q3w1FRh8rtcaDtthTKmWC+/Rhv7jW8HHIPIHlaPBc0SVr4W3p1e49oQ
4dvLKO3ZH9iVte+yF8aAuKkuSV2mPIW2aEACStFLknTExb1tRMiXH1QlkK1fSYEKcK7TQqfE50iB
xqNYPh3K5cHebxXJ2tp4KlZKmO5wMhs3evVZj63doMUgJFpsLJL2zk1Wl+/PQrNu7DIFqkYWUdQG
kxOHRjgDgfDiKv9nUraR/2tIFQ7osseHXbMmDjdtK8NIF7dTarc66Oy7uOKf34Nyx7sezd2nT5Ht
IAvLl7/xI4NLJkwOog1yflbK70Q8A8sB+1NTSKMftruh7dFtT6OUwOlyzG35PsqfLmeJl7stdOEh
kqTiGYxUeSBxcJutOcowo0v0lY3+ColL9uqgCv804sHRxTSO9z175cAcGBTN6sOiF3l623mAAjM3
Z76iLDZQv7zOLoVlJGdYFsJFLdHAOfbVFuzZbrXTxeP4TFnySle3eKw8sZUP1+YCFR4y7xvfbBrE
5KPzNg2yK+S61Ke7VJDYbac9G9YlwrUBQAFVJxbAeLw5mkHs4kiOgMmeGiFdfiZsuLLT100UE8Xu
1lsXUg+SadlRTekF/B3vskUh0OEGewWOVOW7+QXv8gn/vB9ygAKmiiTicRy3XJhojLonecHv3O7d
mgQ/QzirBVsmrvAz/R0hMlicD3AOh3GG+MtkxcvYVMqGSnuvKWtHcvKXizVrZn8lnWaLFHJY4/8b
fvyf0PxMSJ9ukg5c5f3gjsqSlJeptgrkrdzOFo68wtceOwd3mPLOopxAx1SM4/0V/PEWxNbSUYxE
gifs3uj2JxEQ21nDpuxjxem3wmHhQviAFf+kAH1QyNeJFNw7eHdHuTPqj5yWQ1/gI4BnG6kuTScQ
DozipaRifrfLxzu02DhN9+MGmKzPEGtYuypsa7tAmUbnLeTsnIsIeFFW9IdLzm9B4zdsUQuJiw1t
j+8nZ8UapQ1cm9/MjkWHGK3r3+1MSX3AjfQfZZ04a+cZ6pKPWkFCSdf5GBkgUpygGK6X3SVGpikW
asULBmC9M4MVo6GBboL1pZ2w2rfR7rVWzzwGNIxazxJsirfOCEQXD8s7xlJ+6WJm6oXoOr7pr10R
zF7dotZWxScA5CXdWaqz8bgEoyOa9BlWnlPggFZsmsVaSrOKdvWz1rCpOxyDRsnuzqvpWnC+Hyw8
OcNnf4ZtSGhxgCXGvlksFsfom3grokxyI+oxmvrjercrYQAc+WjbJuI42uJeP9NUKBrnEJXUYUmx
nTJwgJrhJRxmV0Sz9hCM0vIQNuogwunmnA8B25jlbbHcAFu08p0jfCsqVyNxL67q28wkm7nV786+
z9wCuwTdYMRp4fwVq27msfzzYALwjr02Yd+WJs1Wn48/2W6esA+nYnQaOsCi4QnOatqGlusRMk9g
cn/T145fIc2CIUeBo6gw9mTHK1AaspLX2wIyR18ft1YLLxmMZGecVEp1D1FMWLGghTgxENMB8F86
x52P/fpGNUWZ/nmdgkW3
`protect end_protected

