

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SQUyeNX8cyskpzvvW2T3ssUGj6xZX5vHX5fJU9Ms0M+rWpNjMO6za6Zgr1K2FMwHi+buwP0Gw29j
IKEYpdzZOw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hoBaDPgZL0nmY18FE8yzpnxIEfx7SKisNM4FVo3Ao91EGtVywU0Wb7yA1enrW6Xd+oLWYcrMdoDX
JTxy8JdlM3o+jyjU7UKGIkB+vX642Q6fBAuo3SZKPKM/RE7lQknQIOi2Y5V60nbw/AM6mvYDKdTS
wiPRLcQIZpvU4dn9GkQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o9OFQKQt0GaB68TjFqZyGwbFj1TRgCs2FzlOtaWTgxoDRMFT9IEssmRwHo9pwJ5Tn3OigUlzbBbd
XTy7vthduMEKESguEgGeFDAlZPJdvm6/cpwtG3omF99Y9vBxA2K/3YI0+jDh2eyUvsHMcDbQ/C2p
zFKW1hcipARgm3A9Ys4mkgzXMVKYnvnQiSsmezjrXPsPy8jbFYPXFd6vFSGi/ZwrKMMLLNZt/Boe
k/Pl01HBEt/KNoY9VFx6N+e2ufES+vAz0H+DJSGPch6YdjmhkZUj2llujVX2dT6EzXeB2X9+1Sar
qYaNJFQdqXN7nDqoQMCiwqUZBJaHNrPJdzAMcw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gMFEdGC+ckR/NJmX/aszkYoB651qUCnYvXxq63Zrpc98jREIyboMJaogrhiyZ1kntx31alD51ug4
ZAed1vud+wZB4IN9oJ1STjbhb+Zj5u4I029j7Gy2lllPl+1O8Em+DnBFlaNak9VTW5oxld5AFJs/
EstFEKIMT8MSbegVIEQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I2MWBDnGcReW7SMjRXdvt63Rjoo/gu+NQcstRp+eRPxV1cdY3BaChhCXefqNXs4HwrSwjy6eXoRH
K9pkdKW/MmeSQuCCGBXm3SZnri7VuXOoNwZoR7yYcuzRHYCe4OVzWrXYc7CJVdShI1TzYNVzTc69
N+748OjVGLm080Ri6+7tnRVNASpwPZfo8iBz5hClukZRieQCUQgdHIAZx2RjUyVQaoW7cJ/urtOZ
zr2GA2iDsweYcuo/xtEmVehzY9Jjyk+XsH/W+/8SFJEIN/wAiWoW84/gDLItkUU21xaixyhQCl/Y
sHoICo/iHc8aTOV1SPHo9yWYmV0UZ8KJqveuUA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`protect data_block
3ovu3sl7IlRCwU2siriigmCYN5r02MX3DM7IdgLXdyAgpQU+6DzHr4JYOVe/ML9raoNj30rqNgkj
8D6964c4W/JnLJzI9hXFp8rKh99h5LQR0CCWrDbx1Rs9VyCVSVGYABnwnCcqgiuOLZmKo5KjjoxF
U+mErazXZKOEhGPG8P2+opIWq4pApWhA9t3mi2n4T8jTZQs9keqlMHXgjgQGw4+BIiH5FQH9sQWc
PEcaYH4/Ytx413BRP9V3UYV/InmmckGVh7ak3/zHbvdqsWB5uive08tbOH8VWeneIK9lATvTB8Vg
1ybkS/KwlX5WZ3sYWW0XhBtF3AuuiZ0nMyJr7+8m80wtOo7MtVlOq+wWHvCQ+ebi3vLmoM8NVDB6
LT4JYCUxOtCPARZkC6gS9lNfQTf9pT2+PNfiL1Gned8ChKj7LJ9wWEKT5wgrSGlX07ko1FUWvVEE
7ijm45tx1JUQvze7FIYVdXwa4Oh5G9zv0M/x/Co1nUTrg8uuXy0pyb4EQwj7MxFb5CJ01jjAtIaK
K4D6pKSvTTM9LTOZQ5TIPWMLNGyOFJHxjYEwk5OMfFbebp3dSwPurYk0lm6yAdNqmP8CS/8mR0pc
gt6ZrkiNWo2lVl2WbU/8d568adFWNmn4/HieXVtGnrE4xOtIqjfpUso4RBiD+ypiBcE5IxdOitpt
WKzhsCxTKnb+0Pnoj7GPYYZDIHGeAvEaYf2xuzD80tY768n/zGkoncH7/aLG7kNbE6dHR1waY+es
orvQ4BR/g0OC/KmSbrJa0D99Ty9+AnCO2xyiEmu5W3SWRK7JiP1rc2I+G89b4DV3qzyMJylN3IqZ
E4zCvQJjp8aS/omIofO47tK7wDoOTwGCzxxbLmhPV6nRyv036yiEpn75Ej2kYKFy6xXznl+wlvXV
SRRJYDem0E6hJONIvqZ2TEBr+8WPulJOTkUcEhwpuRvjyv/02XqpdeFex9lZpO6IGDwa+Wew5s4s
kKKuDwt4s8LzKjppKReWHiQ0qckRL1mtZSR3lzkPzFU4MLXfqiremMlzN0l9LvdG4js4Mk7y5Ign
iBJIhlk0FI6EMsEDjHIGFJ9H2mm64V14X4tnwkTXfkO540ZUWnzb1OdllLnNFAsf76Zo/go6ivpX
mG1+7IAJcc+eYwuRKptlp+dYEGqeLvDoY3kXPEiIHQOBlXrYrNz2EBhtGsZMAwUkgtdyFfipAS9M
vV5Dc3Zxvv8r0vnCIi6M3fkckK3AUAj84eUq3u2FRMS9AuGoEN0am3Il98AX0o/cFAHEmPYPgoEg
K5vdc3YbIC7HZ1pQMwsRORL0sXqhAZXir0GsbKMXaB+xBBvXAMmYXNmqe/WHCLPyi7WCD0kiy6R/
jPOToTtOK3Gu3FmHHMfmNo7CXPRgLrFI5VUSP3908iMEi+GEhvbOAhe9wyBMmXAOkNo27l4AALp1
Frw2f3eNHgFuaL99Ke10zd8TfxafCbF4aUDkmllbR/i+CZEbJmyRRb8NX58s6tQgbSK97zBh1PDQ
ymZodgOtJxTnqgCeXZAUxCHwlv5R9rcoQcx/vH7K0mKhoBaU2dbXMQxGxVnSbP25ilYdPIeiQcxM
jfpnpwlXRIudGvkNqXIX2PYU4y9ngAlhpZbj+BdU/2s2CbRyFaTEAp7AFnEAhMD18g0BK480OZvz
niTHnHlxZvneN8BkR2vn2i4RILewr+GLXrEVMCZ5YX7hKDDpZ2XGt2yvIT05fDX6YxSADl4HEXTf
ge649bABPe0FjQKRBk/k7fPODENlJEIxCd9uFJCASwEiAO4CoujN5JSwvCIy9xeOxlEVZOSFF8rK
KgqFGcpOUnogLeaJ9fg3yS9I67EyThoT8NoRwWz0ppqoA4mdnYo7RNc53ob6WJPsv2yFCYQKsx8y
uug+OUtYLVdlRBYSb17n/H0p97XtUDMCc1wJ/8i/IXIJkZa6mfgFSWXtPMgKFr2AHDNGbuEW4V6j
Dnsk92ecoOcH5rIOZafiV0QEd8muEWO1Zgq8gw6v0STiIlji0IKeM8KH8V81cWcG/H5jAAjmRQRN
xW9bE4qy+eZeveLJVw095BxWPNhnV28dD73Aod5vBsqnxSEGGOg45X9ag0mEpdsc3pM62e1niSz4
v/f+8Iq5lZenBNXjR5sPODaAHdDr8NHLgPX6GwZq2kBh7ifPWcW50SapwFuAiTm396mrcQuzqmIQ
MVCm9Fv/yMX8VL/L+u67ME2qTwWsNoQX8WedCjG2qEgxJgNhhiw6LsSmREkGVBWKNuAmbur+Hqg0
IhXqYlBlXDw/dJafm1Y3ODJ2Z9oTv6jQPP5eM1GvxfSnfwTyjG1c0iBiJacglL/woWooOcoUz9h3
IUHaGJE0suAl/k3+wuNv2HqKFDG7ASng7+YXqGRR0oQzxX1Ae/d/EL6g6Woa1X27DFjBca1/Z0SH
jr+bJgPFjxV0dSiHrA5wJ4nT7a4xXFc+M8K97Irp75Z2zveJRpZy1F2T47Q53ux7nn9LnB5NOYD7
ZNX0bmvoViAGGn7LsU+vz6E5cFeqgWI0FTbjjtymQdRNL9Bu2xPJuwMGiXFAL19svuLCLpwOaBwn
VStAg7gnVqOYEia4Bvl6/UbHqG0/V4GdXRRVXsT1xHbYxtEL0ICsVgF05AaTSokE10ioQOP3x1YG
Cn0cZ4zzLL3uSIOXvjl81Q9dc6Ye/jUjDbZOvY4DcWONMaUoMqvquQuERvPAGQQXUOD9ullJz0oo
qW9lO/9MvFOLy7aPCQ+/IicD3BbBDu0URUa4GiauPP+0Qpy9Yb4jYtwmFq7DNDD55rLGnlE4tKvY
6VnwKgyYsA2ioEZQaY+laUcSRTGccvbA4Y0ai6znBkRqiCShXJWJxfBUc3YhPJFJGRVVNoWUwzvs
NbQ4YNIg0+YK1dmhsO7+oVeuXdjqnZGJeUQYercD6gLy9xd4mHWg/+sqmmCjXAZaXU8cp+5PkO2S
/7Ux1AQ6XSnYDCzfeG4QrPY9UZULW4X3WeuoZKt46haI0qn884+tbM/LGMRJfGwZmI94g5wvEUW1
AFJTycjeWSzga4DYLwUJiipr70MXzczVjbUGuekyJ7fiik0+q9rr4z+xpNTlJFz/yrULlcGPXp+7
i4mkh5hPf328WNlWcdFpQuv98IOwxNtXPunoR40lEHZcTD2HHU9FF/1JEVnx0Yj30v/6MlyyQIfB
zvEzbEvw+YYXs+4KeyCfAIMrS3y+x827p7gwcwUP5VB/TYEMtukGTspcQTc0VLpYaJd6g3JoFt++
5gU4vOjjI+n262XhaG2iK6qNFbvTMHDeCzicHOvmk9tuGdKom8Z0oizjnajJDg3Rif88+dHwf7Mq
85TmN7hv8rKwn5lhO0B02BYhZsBe/Stg1YUDEmijME91xrfskGm76R2FhHFdTbL+gK8k/vJ2EOjk
LL5fvmCLNXc8+bQX2sHDPu4dS17kFTh+QGaqxu30+qsZZHdjAXto45ilSvZGowuJBCOieBhuJ9BT
YoYE2P8PpDzBHOKXWvylRYqbTIBYBvQe99RAlrXF84/5arls1dKMfOjjQhis2PkKIcnn3aj6S5ZQ
NP0nEK2wJOQVvnXEjuVFbATfGG6BNCtNIPXdW5gKmb9IRwh3/NSAcYOazo8roGNgrE/Z+Vfr6Y91
nH8I+L9wyWzimpgTv7ztSP+//1YoComnyjDcUX1Vurv/uJtY8UPuXeHn6yMgJyF9BbwyV8GicWmz
3AP4HbAJD3GjEQLNVG9wPBqAL5zPxb2XezNOfSNYTfS0KtR56wbM181KeLc4fxvywQiA1tyFe0vP
NU6bkvYbi5ZoE7zaCKotjnMTMcAFeiVc07jy0lHBMh1lk4Qw4D/1mxoB/IhSOuTq8kAf+paIdKsz
A+IMOk5IBotpCSUUMvn6zq5DSqvuZyqTqAmlUrojtpL/bcuYu3qGhUsBol1v5cr4bBs1jt/h6sKr
cGVMlkCkrurOxi0JigpD/MaFMHV4fo6ubngAXSc/hRa/CVff3y6WtUBD0L1zRAT3xG3DOCgH+4K8
ENm12FQOIxfB9hMQ2BqnSt7pKerb0oiT4RDRJxPQccO9tvlZDTzceKHo81yLjBQUcEPK2xNaPWvn
cMHl1913NAM5aXdp69QCTY/i0zCLiQ4H0DMxMnnK0++NvkgB5bUDEVe0uera5GEaeOmKrn1zGgdC
deZeOUgxmDRIzxY3LSJRdLdV5Rzn2Cnu/lgC5sAKxyuzq4r4u0WpPDJhMN4uuQ94+0GsGsFBnQQm
sILagRUihFhjqf4q05CKpXZqKGDOzHFVT9ej7o0cQznMrMNjwtrOZg7ctwaaMt2UNKLJ9ewmnkYC
8QH2hPOFVVYITWpyUejhkYs2A5uYf+YkZXLCIwJA/QIIEMKcjWRyq/IjdEj7qnPgIHUTWU5fEswP
A0woKAXKOhn5MDcFbl6ZJO7zuGiqdf3IPp6iwW2Y4bA2rnTqvml+S4MBGdh4/qhAttSEegsrHCSH
om9A8AOgGiR1MS1+ET2cuzItEpHTGSxv1GppE8kdKnsE/pmUby9a7V3kf08bwJHgvHLsGV9hcY/x
I6drY0FHhFbTM5+3NsvvZGyrKRVYxgt32PjkBPNOr+E7qXKqBzjrh8F1SX2GtM33U/LtAwqgRJkO
bEVc3G8WpScuG7JUuPR4kAS/AITnHYJVXeZkgAIo+AV5pyARksr71dKEVKuOdZwNc42NHeohZlv7
dAwZNZ0QGIVDnadl7EhNolRxVGbmKHLWjNPVKAwBgVrX3lL9FbFl9Q/EHVUbHMnIYa3Gi+G3v0Fy
z2fURzinCtmWhkDADKt/pDhm1UW01KdjTwIJf+r9jCcg2rTHuNCr7qSyCdvYmzGZB9ghros2VyLH
M5WbrsTzm3eXum5szVAnWs3J00XGy2NXFX6E2iEiR6KlMfqcexV717EjFRrGjC2lPkDXrLnpAg3d
Th61XPvsscSi/yMmVjB5/liX7AF9rgpxE572OrD68hUz7RiSvVSIbsw42wrICxKBdzgyAPpd37PF
aGRxgu2578tLxNW4u9j9DerswgXLI/5dbPmFvhgK0vkfQtP7QL5y/h95mB/YdNlAu6lPipkq9WFc
ouhTfuSY4DLwW4TBwNxjxuIORsOWuExSNTnBORM2i2GDsn8wAOTH1uwrgQL2QlWSKmpBjMKye6cf
kvSB/j3z0OyLQW5Zl1VIh60aDlS8bYOGRErrYW5FaaSCXOu8XILzY7pjKi6oeLZ9r0r+cPueJ1JR
jyuLygYSdHvr525wNnpajh/GoD01HuGRm11PzQFUX/vSDJC6Y/BczOmDsbp85oIuuMenfPkh8xYE
Mfh/PPgdBiJWKq7G0VrRf7h4VpoeR+kTCqYLL5JSoA6fsHofdM1dm4nemPGeGwO/W04vjIHs0ryF
Nvai32EwcCqctKLvhf41FqQjh0gcviR3lcf3QcBQ8p/RY7uWF2O21Uh6+jIOT+rIEjtcXXR6b9eH
n+/eOJlBeHoneFEhpBb7CmTiJwLDhBQxuCnEBrAdSD1/wh+n+Bb0+iRZI5em+LuBaIu9obC2Wn+a
M0EXOxqZBazelGN9n+Dbwx3LDk3NUE5PWljBJ8DzwEmW2yMD1/8LVNuDh687xQNpX8lVmhqLMg7B
1wAlEjnsNrhyv5j954Qovg9qQXCRbhcdOhHxIk46d/+tdh3Jvl+G7CGhgCJeiF0Nyzmnn6vAjgVF
/n1E016dh2EKjIxybgCqVcukFZCdOApP/stpODgN3BsDVXP4xJcHG47O6vIqrn7b1b+Sk43Hh4NR
0qzc0vpmiFv19dvEB7ZvkVudY1ilIr/Jdd5dainBxm2kkL1+qrAxRr7t7eXwDedY/jaDUUYIzQqc
Z+DmH72CY94ECSnFyrm1nQu4XnGCljmUdmmC3kIbkO8pexMPb83pfzzQd0t+YAMWjVKZm+fhPdaN
+BhUwr9FTKY8tUrv3eMGdXv7z9nWoxaXUNjzqrGi6nUGFQOoREFYV1abhkZTmDdC8WW80zkcZAFh
DVHVRz43dk3Y35P646vgPwB9YdyAbG1BHooTrGeWEEUpXMiWxjKwk3iKeWi92p1xqAqe6zYbUNaM
0mkMyHIT++Nthhatmf5q9vDTDVAK35jmNjhm0TSNv8qL54/DDpGIgg9FyZdqkZxVGtMTcIfBlVYa
gK1yIswOh4UunbxJVSppC4osBVvXMH1USJRrv5HljHpeV59lP2if5H0iEigHr3qeRbHi1iUJUzKY
sdIivTyhdwvUCwNg+5CifEDEb06+Rx5tT0R4uUDHHVXgZe0MlQKv+j0fJwtiRHz3rbqshliP8XN3
20yWaXAzd/F6PydhViHQkl4zVDQHrTpbnRG2FPe53ssU0zjffxW2LNwjr/5DtPeAR3a/IjlmqwmF
UgOdQJkz3wks7QTNjolx56VwqMEl3mdSISQthyLaQlbsAWVoo1+WxZT9P5qfeU8wnehe2zr5Nro9
h3RKZ6CzgyaucVSKuYe0CFmB1zlJWZIi77fR+dmBx7sCsn2IaWNy4V+dyum+PA/zPCN2B05hzaIB
SLrr19z+V1Hd4f571uvLh2okyRNi2VFzAhpqE8UmPdYmsHiJUYBFnwvUByINAwus6wJuEup8OU/b
zZe1k2khfXKhDB6A06ou+U90/ktajbf0zFM38RXMDw0904IqmqWtkMAXKk8+Pd6NxQ6j/gYugybs
uzMFegIh4e5CAV/RLApsQnVbz4LaASu0yzi7cAWXSh68uFvRHuD7Jeno1PhHlb0yo/jzrAEwDXxE
GzzMyYf3FYbsiF12CSr06/gsJ7w9SV+PFYXluoGiIA8d156rcN2lmpnDwZ6X0dMqX5vtUbzmNULa
xfAFPlneDhT+9L+rwc6xpqYACC94lzMy+hnlCMWOlfVd2D5iPJG4Tg7gWYISe2VlsPSGGqE3w1aM
yCAi3p36uz5FtJNB541oeyshMLbxjGNl1tr3FSPK+jR9WoY1L1fWwWgcRsWrXOqQUSgm797YI+pa
RGZLnQdUzOI6Xa/prJQjZe5q5zwd6WwQKVL9uGAHkaDTKJmN+pSQOSFjRr+6O0pXCOoEVNIeG1V5
PRRvrc6TM8kJkSBSGZGPUZQpFUspn9V4slXZ7PzQGIkT4cPEvyvd8JQXi7P4ri37KYvDWS0JF6Zc
4jp8u1JNa/WLFLxs7JOJb6bWylbV46TglcceATPTxvuJMhRRLd8MyS+YDg9S6DQUWasxvfENBZWV
MNFeG8HXmdgIrTXXx5CR8LuharjGdIUv+kkX9pvItoAuGv3YiBTeB5QMsufpBeeV5LdX0wlFHFml
GpJuuIxiPPZaYMFe+xdYjfEY9IQtUyUqyPcywQjbvzy+X6HgrjAsAvNfFYEcKy/fKUyEsOaFsApH
q2HgXTI2SJl5IF3DsfeiW+f83x+FzEeVhF11ZBsrQjack6DcwYhKlmHku7NJ15XbuD/QG7AplKmT
lDM4VdqQBxnrmbJf1pAZxteZHUYdbrxTpmNKPe9MSBPQhuu1qS3bYX7KDYG4cSEAHj+qzINMJEm4
1V2rv4SS+9SSbFtLps3iKm1t3msiaf7FEiFbKUalaQJwuX2HgkYkjWEYfVFm1B4ZlzbhbUEkdQ/d
MHytUJtp75XgCz6t6YUblfhkQVxVy3vthDXw/ZnY/HMwx/2SaH26Y8aWXGHRiG8bxsWiWqN4tINq
wQGSdZqTtnI0dtJJj8ar6WXFS8lvoa5wZbrqEBPAf8r7LumPvi/NSxLHizBp/9M4A+50DLCc8PW6
EcP5xT5UxZPE3anXn7RkAkToV82AnDZcKTcpt/tANZ8rW8flLLovMcLl6VnVcLNLxbFc5EhgFmio
Mf70kwocD+3HelbdWPIP7jKU+SsP0unKoK4yYi1lIAhWEgrCaELs7pM6jYryWI9QQf50Jx71QWXj
/Hj+XS1nC4NP0y3DZuXiN9cC6cO0WbFu1ppO9qIPFHnJKg8evfg1HsVotLSoplgsZq0ob/6xI8Tc
Y74rPxVDMRM7jnjT6+o0YVGjHRqkjkzqe4i11NKHbiPH5whB68CnmpHNhIPZX9iTr3lFTjRf18i6
tJ1DJxc0m2pjfi/BZPjeYH+HM3r6PJxinmsc1mSCk9CNASYJKt/z/bXQWNZmraPxLzpCGp4E24Y9
aCcEVEYmdCRHX7h51qHfxsmcibBUvfiiIsFhOwAURF7czAIJFtXwuQQ3wTUp18iZR3dR31crXBtA
VbayZXPZ9HRazBL442mmLwti3/qKkP8IApOOjRpYvtEPpK6kJ/3x5/uiFvRVcCgJjaA70nlpZl5V
yZAjbSgJmJpsoxRG349tq0Ia/SETSjvH6M1E1LwarxrG0WVo8zMDvLfGfi9/MH+3307KsQdXVHP5
eDSx0J2Bzd5pfureQtmfh6QMboQwUWjTXIFZwnrXaow39A==
`protect end_protected

