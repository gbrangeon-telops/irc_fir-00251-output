

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VQBfeXA4hP5orKlsy+AFFAe2QBxKheQVMjP9iwMw/NM3O4tSdVMF5nSpUCi2zqd6Xl/0+S5YrDyH
MbW21sN7bw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NYnVtYYKs1fo/NxKyeagmW8datCnZRNIFQJ52Ut8vKAvoM6z9G59Louyi6BpOXJlK7hkOA0EyUcq
xnrhn5QTbG+/jjVXTRQq5boOLx13BVtwMvklEuJLJaUCJSI1mkPVMU1Tw6P0C7fzMTIVY1MXBSgF
huHBAAQ6j+Ca7SHEJMc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UdRiCUwOSibQJYHOoWlsqKR136XIPiU7//1vC9LO+s6bwL8gocVodj06NRrITDP0xKYK2ZTek7T4
6OlwV+xWr4k2Xf/sx0trTcVrHoE3bps3QkJHk441qMX8BKjF5fCXU+yOMX1xkQlvuWSD8+NvN82l
uzCDbBA0KjOv/IsJg1WHwqG44dahfC4qa2RHQtygQ4MsVR/PxcN8lnUdpguLi+YyGmh9q+fLgQBq
cNHly9YC9ZC1urY1hg8yqWcJm8AuonE47dIMtl55BTxzCygZ9uoRy68FfVsLU7NHg3O2kl94A2uq
uulT+/Y74MIANEyVFkVes/FR1hhgCPd7uNhwkQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tQM9oFLCOLGigsR+dGte9FyrpKbOg0a2HEe24uc9a4zzPMiWT4Zq+VUMyysv3hVDjsM6Rhdx2y1P
MMtJydYUSv3+V7JQyYwaG874Tc20f583mvfsydp9rtOQQwZoTUUdaw84/pibQ9geh55pxtJYjyzk
ltK5Hf2dDqQ0W2qoU2o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D9jeI9qTFJwFpVSxwOhVsb671/UONJ+BqwlU4oe+K/dJiOTSOoWnMaaYQ9Sgy96AbPfvmkY1YYgF
jNHbjBYJx/eNgXJH2lhqUlU4xX7po7K9tZYQraj2oMsohZUwz/eLwj91c7VL5ZRmCXaHh3hDU0yM
tta+u+KG7UfDjSpBDQDdNd7gt/bWHfns3Zj0BeTNOQ2o2kTzIQxImWuXKku154pI5L0sF72lK31n
Ls7v+PzriYFrSA6JTTtqAnDF5uCY0O6Lpa8FB2AoeQSutIiakkT+T39fToTawon3SeQIsthaDWDT
WAem4lxQFA8q64KvDBTwguerI8Z6/8BM0gLy/A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20752)
`protect data_block
oQ1nuFqT2ZlA7HPdeJg2ncgj47Gt189PXmRQXaEbMFkJwRxFSFJpoimR5QGfVmBdr9pnRQmjjlm8
tW8fUOoloOk4h1fLrENp24PHAocHpbwyfa+YgDxDMIxzS6O0+OT9moVoAnGZFWHINFBzIl97sjyI
dKKmfseBA/Hvcgk0/hM49fxWJ3yMuHWMneAGMQJef6Kf/p5vizBZUEqwxe6ysaReyFHWNPW9sOjM
2QQmyQCrq7bqlIEyd04Y0IN6LrtKAiMeCp5VJ8owR/iWGsyr6+bZRDcAHKcrnuRAgkThuaArHfB0
eeOrM3Rip6oiP3xqtx6RcU5DTKtFYk80MzfPFQhcWsBG9iI87UPSrT4+VzLKBZwATUMb08rAx9PX
QBA/rkpeStGYz0Pd+RLHMorys8WxQP8DNkU8Ng4UMHfFw6Lh8y1lb9xc3WEmGKAtDodGpvlkI/eo
BYvD+8KQjWYS7bj7deqbf4LxP8Z4ToRyivvR22UFTFVs0365i9HcDYg+HGhN7IWNaz0g2ae5ISci
BhPamHWZPBpjEHbzM3GYuExHh42K9gW1flC2Hp+r0GkuRah02Yw6TLtBxiQzW7+tNvIABv2sWMg+
2XXckL3Set1yPHnEfqaG9ngowpjheLYszOKSoxgtH6pC6t+VLC+OPZYWQ8C2013u31yHRNvu8Lya
A/zjiZFw68e5f4SqnR5rASq8qV71bK4ESEJbm+/N/G5uk32Rl5quAZ83mIm/GcEoZAujRVXpga4t
N5gMdGRxQxJenTkPs82e/Arj0B7NI0bAxwjYovln+l5Ad9IRPrSUH9Ab3NcBTiIOIAmcV/Wp3XLy
ABjqeEwuyo1jp09d7cZEDjXXzeeEqtzIpJy50AvPeH3WD6cYXprm3KtByOeRGnhlAngo+A6CuSF+
SvYzB/SCUcHPL9mnR3rl0O25Xi1ZgoW09q2xWiFxMnMvjZJS0himAfIEBIqplm8nrQBBl0sQrUMA
HsHLU9XPWzmyiKEV6jX8yV1oGo9CIQNoPuwLUhKSNPLP9zP2EfMOeV7y+NX+bNOgQd2O+C103gmK
GzF8j2RvG0KGWOkluyrpm1Dje3VayF5ngCLmZeXm6UwEd+8lSN05n6y5JlqZC5Mwy8Kv2mrzfW8R
6sxM0dtCrd7QWhfpDEOmPlhIYXMNU/FpyBYUibM7sMzo0h7E2jzOwe90ad7b1Nk/MynZasmH1s5P
jOtDOfYn3JZxhks2TRTVRkB72JOwBzgY5mrfCBIHuUuvnf2k5PI2N/6JC7W9oBddtZYK2ilfyUV2
uzqfbB9SySymA1S7zjqjiWJIDMkAWCs9XSJiY1BunLuBzTlnuf9UJZaOnbNqARotklShrAGTIJsz
wUIAXcVYLUqgxPoIkhs8ctZavxcaBGLHCFdfBDDsjma7kmJ4hrmDvStWwG/OV/1pGUJ6AYjus7Kd
tYipQcMDZRuOb+SH2EaasoSjxr6uc920OTWcH9AoA44E1xO1EE8hO3abY8+eleF4Bv+oFRM1QQhI
zRa52AvV5RzV9mrctvCSB5XUAonyWLq95WuhNZ6hpjURTM1KDY7mlnQA206o5/SGPa+9nHWi62ZS
3eXvLYcyurAWt+RlGJjlel1exEAizQJL5GJ+WqJ3WmqEtXCdXULh8MeF8Vtf04kYy5/9WUodiOwN
xvPesX7drhMVoEqBzdTVP+WCBIoyl3h+4HbmIfyc8qrLG3d/b1BRC034JkgbDxjJ/yyHo5KJKxWH
8QRW4YwYpz/nVJ6sj2kRxI98RuA1dGPLENMIgsTsAjsHmTF6J1Nl8EjDnhtyh1lKos/UABKaB4SU
VGV+74hErEJhNATBbnumDMvkin3Gcc3GNSc+bhAV2hVw+eFDIgRXJQ3NuHBjPdxRkj27M/xzwjfR
OM3ho7SLjF+HV96H4Cfglm2fxZFIXxzM7BvjXwmDuFdEMP8epI9zXtbD7IxIQLg+bae7wK5WAABr
ygYcJ5ZMNihXo9JVciXABvRnASvU9oXKGY43Su97I0WtpV02RTDi0XFQxNkGo/ZIe8zIaHw7fJJ1
w2MmV6m4B6GZ93bmfpQW2tLZKf6JJP0HfZppzap9OqkudD8018pfgk9Q5+G4wtiXHJbHgSu6aEa/
J3En3rynNbBRSXbw6QF+R+rGmYgR8n30y5CXXBvGKwo2Xc8AACMZLbM1DKrGVseYdyv6NIpuFNh0
/dAhSC6v235abee4sfx0HHNFdgTeQkZURhI7PYdNUtFUcx0BDfW8LqeYeCYIZt1s1odg42g0UFdt
mTIm/LWuwkGhyQlzsWHGSIQFKhoTZauZ13muOL9MIrZAZsDlYvHGS/mtbdYBokXJSuSYzAcXttqS
I9DI8hobJdOXfnzoH7lQOkXqUJSKzasQ6HsR9tW6s32+DdSwFyjIjM6chlhP4gyIgIM+WV6obn/4
W9gSRxmE5Q3OgNOSwuOA6aUClol1g6Pvb+bSZkUwlIprKf88XPx8kYmOQjhL9tKD1gpPjuH+NycK
8f4IFbSJB24Xn0dYab8MuPrCN4e6xe4S8rxyG0UMgwu3qNSc1IuHIuAUveAONliQ+YhYkCA/CKHn
srqQnGn5glyWxcsEaWZo2pBOzViVC7GmmzCGcrB7eelHH4jQ4GKhilJ4vMIkhomSYnwl8dNn5s2+
Whk1aqibYx4CgbyuEqTptknG0LYyqesJGOmXTQiiQ3zRzVq7G4OYk6r4BemWXWorxNxO8UmWaglF
TY5JSELgnOJFYtTYNaDjeiABPvnzNtQ29IVSc9v9qm+Jd4b4ClSkCuMcBXUd0vVjvBp4ReErQx27
FAgJ7/C8UK7Si5iWVdDXRF2fefuSkIib3UuqLt3/wfIKIUcEqQDlcymh24ed8CG6SvH9A8T1veyV
5Q2AW1xAVIYOo0C3Z/MVd2Bm34uvtcBaCPp7s0LIauMA6Vb9aSomyeOtEUPjeLEgKLE/DYVz7q18
OgJkzOSuoOKp1Qe9WmRPIAfkN1Jj1LyTFK9gb4MMAZ9SYNqOPzK/WvOQ/PeTAoo/xoBLNGWr2wzi
cUAKb28yRZ0do62WXJsGE3pSiCyjLauCuqEMOtEEVx37WCU3uejrso2Gu+09jYAASsMbeYECpn9I
86OvJdRYpQK4vi4TdgVGpgFLuxZzVxSHhBIPhnEKxNPuZl5JFhLiZSYaVVcKfXZq4O+d4Ma6xxPz
H3jL/fNTemrTce1fhstFU02SznBBkY26qO9oH+h+XxvE1bL1+4cKVv1Px0ypicyjNi8M5sR52UYe
BWXO5MfnxzuW5ijZxC6KzmpBSj8bcDcZzWRPDjQgaZdSIeUYICbkXvmgxyrV89V3u/OMhcaMB0aa
mjpL9fAyBWz0gNll1k3jdMLYIe8OD/ti7j/VsnMzltkYZbM7dXRqw2KuUnqOuZmg0eAdnIh1KAib
sk1NHA4k1mZmWgADA/wB5PN6oqFMNtg5a1QcP2xuWCi2VFtG7jwNWmDxwdpf1Jt204I6T8FycrN7
HKwPFH1+gXsfyBr1Kp0fu3yTgbQC2rSOJMTneDrYI557JOJlsPxIIKishaiMvkZIhcftkgDQ33wE
LoDuarE7sK2v5xj3xE0RBAXzp0UDNqYRhAfw6GHXDF6LcUIRpvEenTzbVXxuLGDemrCRYiCa1Lm/
BOeVI0AZ+24nD5ByEzXr54NKYU2huia6rNzZvelkEC7Y6NQ/mZac/m9DBMac0l/sT7GllCHvCkH+
ncd6cLZPwvj8+kfrKumvnCvzd0PAcjwP9nmDWvuvV4kE4GJX9miVq39VR92Uld63J2wq10u+02y0
tBLgi8/1mfjEpK4Nz9TgMBPk1Ly0tTAjBNU+bfnHGixErr4aGegY5VcpC9MXaexD6GX3eZMRg99U
/aWKZy8g4Si3HIFd1y0g9jvmy02LgAPTE7m8zwvyNNSNSfJGJE26lSZXDAvlyJsuCBTQElnh6AK8
uAybdJBOFFHuOXw7C1U/k2t1H11cnos/BKz5N95dhNoSo/ModApFoZZZFPlsOrxP142ZwOcuMQRT
iBlMF+3N57aAaPZQOW3CVyrz9cp8nf/uHPaqvS51rXk3GTWv4Icd2kb6YhNeQpJAEek+lirgaF7B
O2Syoo0QGAxJ+edsw7VWoBxY6n1bHnl7CLdwVwWnX2s0hV8FezwjNcri6cXMWsNaEA7MjT3SuA6N
IeHXHJnEuiQ8u+76+14T9Mm1i75ej9FpVGlIW+1lh+AiXWTBmO1NupIkZGga+QRFOVDYslkHschZ
xUjByAfqoXMvkODwjjbqSaDxzQfQbTze2OhFkBS00w4wdJDHybKln5gfb8l4AvFUrMX+eNzF+SUQ
P9hypYt5qXAfG6ABapgQ4x+sKAJZMkiBrqkqQRjmTwxFfurXjrBDDchMAz0+NblRpQ7Ho+LvSdhs
XRgUPUjTSDv1rTX99tvukU/WrhWrloF/5Cbft1od4lrM+9MbnyT9i9ulyTI8hgP1EsWyTKNZabhQ
CXN6F10tUk7vtVlB6P5bpZx9ozIIS16N94T/BeZrUI01OgP5qY0SYakhDpxsuBpC1U+E7vbvT3UH
zrjLAjrYdViJviq7PzMb69SCzsup7lIhCqVBfTKWTkdb30ul2Qs4+ljzeTa6gdUeyr32LJ59jZFa
xlY6tLVRMGnU2Ecy3AF6tDPdY5XlvibTBCmN6YiU11PoY+HX3NjgssOcQpbN4PpWhLz9ykLIQqyp
Fy0jpv9oe2pSpce1ARoSSTSM+nxCV3li+FkS0ZnZB1tIHfwq1Ceke41HgnFd7E3LQRS8/MlD31rR
KIXnvARdmtX1yFTv+k89VsnqSu3panELe/gcxJkzmMDIPMq55g+QcdtfLdzQM8e/K7JjTDbbJZCB
cOaEcl/toToO3/zrYJI+M+6A36iZnWtV0E2x7sfuLkBQl2N1wXVr/+f1EPPPuEM9bzFFB2BA4VQa
6Xo9B8GWvdgt29vtKZYAJuohJupvn8qUqKTVJZPgU6fkKBxu4Nr8/ure/lkA3C4FjvMWxiD0o/K0
Fpy80QGNGOemx6r3nsPS2PuBxiZ2Q6iiECYazkFpHoLm5CX/E+1VObQD+QbG1BrLSjmOpraH6qxw
yxtCm5mGZQegXMlleT2CvQBs6hbTy6wBrq5swi4Yf/IPwrphSDG2Luj2dhDBv6L/N7ddxrmv3dSR
7WqgYcnL2fRyVLspBDB9JLBs8M2V8D9l6+DmgQoZkWRaluL4HrdxTvN8hH8lWluSAWpSKdhWzJOX
NQ3XbY3Fpqz97cI/C8B+C6B3ES8BBKuD7GqWwpvTP69XtGRxNd4ahgIWZV5PnERt+Ge6R46PnHv8
SRJTNkB2YoKgf0XtNfGk9aSpRsJ7BHZ1zueaoBtZPxs4eW6bl43/otIquTILXFlH4t3FXuw7sDM6
YrVBDTdZI2P+x2eYTsFRPtYLGRmdb8ACLnrc/AgoTRSceBEPbQBxVrqyxQ23jMTXuuBOKoKFwal3
z2ZvDXk4XCr0UxkRMoVZVbLYQxTwls02LWQy1YX9Qmeigt/Xuu4/XqwuYWs3ThEIFmheVvRURuOZ
G6iDwPiKRQnSRxbINH697wZGMy14hMzxPoel2VToWxZC79t23msSBFb/HxLLtmjkRTk45T92QK0x
DNYjQyZhMkCllUB7KPRraO7STnWmuWB3+FJkk3jE/dOHzIWazuUKU8j0y71luACRbNGfVkUakfDi
wxiXCtSiYnKFzMpJ+3bwalVnnuJnR2n6qaCOtCEQSIVvSd5im5Yo7MUSOlZ+88TcjHPhAaUcOxvG
7tg8GdEnJhXSHJhjZqYpTxkYu1HfWxPxtcrr1MUvgc+n6rIqYmBev5vTxYYDbqfPO5gsG6zZcyVI
+javcGTsLZSDSElAnyGA5gc05DVrOcj3GoYCDcFhtE0qqZFBUkYvu5NmXlOp5PyrJLXiF+f7ecwz
XKncj8JA2KQTXJMj1O0nu8jk6D5hCZMpV4ns3m0DO09Lp7ZzC+T/SW6UFtW6VnRyR1GJptYoGlQI
N4VlYcHIBGvhWIwN+kjz7Jh/Owp59mLvIHisgVEmnJYvcF+hlBLDJhHet1wRlAqAWoB1jSy7nW8X
VZzMAG0PHRGfwyIHj4OIuBstJ1tb9kI+rSmntAV6ktIjm9YftfgKG3XczkUaB21rdO4pQ/Qw8s7T
ypJY5JKWfxKdOhgCFBi4fRr0u0k6Zi6hmfRCh+T5/tYfqpBbsMk83aO481/wQMoQSS+SOJe22GuR
ot4RKsKK4OnAbHelksfh8blmPs/fshte6etPCOZdjMC66uBFr9AYKogePs0ju/tyYM5WyqNOgFgt
1tk71ZBcZ4hdUV9Kya+y33LqmbgdwKxIKtdpTOH5fud7Jr/17HxQDQwN3g1vG5mfLUF5yT3+b28Z
cfeVowTW5mFZmerBvyfcKIRnRoumN2am0RwlTlkFv77+zrKq2UymAz4CG+89D9nJuqcrcCHTmB2+
K0YJW7nyjYg4bE7o4o7y23iPcAGK0nZSZDL2PgTDXGouwVnF7KMr/PBhRY1SKUkacuFS3KFHeqDs
2/crAyFUFqKZSCg9Or6txpKcTFDEjI+A2eJFrWpAuyFmfRI1nsH+M13cwIiLYV2XcXLVtXhxhX9O
oBfydywAjgZxlxbNRfIi747syXWUyS/f8jwD6B8HYRfDose2BKymrs2GzlQ6o5jl4wpz6zkQrDNK
RX2TPfVRkyinBtJ19fetnC0aoi1BgzbHUaBam8dhfbBqtAr9Yg7bv7ieTP4xRyAuam27Zw5zDpu3
1JXbIMM4LTsqWbbUAjrCeWRwnMfU2UKIEPVzija1JHV9Y5BKpYE4fdlaU+GKlvEU/2mIVn/Tb4Z4
Vhvla+mLUEimRayt9wPBAlEYEwcNfcvmkSHvSfoywB3vkdGNghQlL+Re7LhZwM9zKs71jKqqaTo/
1XjTno2pFmThJv+2ndIXhBVJ5PDak+9lzAWOwLNOxzxXp93yJc9T7yXUX0Rr/Rnt5cvyF0+QMjQ2
St1v97YNAC/M9oxoKrUAoZR36rWAikb+mbyqS8aqW/HFgi8ifMLi55vKS42GZF18wjnzv9H8xThJ
m0VOcYADkco640OUTfcFfl2An3eJ6zrGJ34c/llmppReS32DhtTIKyHW9/xMD7WVHMPgLGh2YpMf
+giZtTm65MJvqeJzWDTl+joOmFHTCS97XEs2kimQscNCbGGypa9biCo3l57WtvZWPry508BpQ0Ub
fi8/nfkw+erzRlOdhswiTo51e8s8n04DPbIYdCapuBTPzlv7I6YHXqb4jlIk10ipX/ivQ0jG3yLI
oo60CjVFScCwcXjfMc4aWfM/03qeyFV3JcP3CM1pEC5VzBz1a5lhKauIFEW2KLYABG2AvngIaUDa
DxNoB5DlFgO8Bq82AutU8Lot/SndRHkffeLgG8y249HSaLGpkRk8e5wc46Y6POpdZPyP0Cbys56Q
54qWI8yHUlJMlJMSOwjdmG1//4YUKz5AghfcRmvb7kEW8/ME5V9jvOCQ3UNwJSRn3x1TLRH0SSIn
1u1fI2S5S2T7P/EU7n+ZPT21XHYh4rTzEvZvbox5azyGWqsHwDF7zkN8L/j3sEtUKvdzzsTgQuxF
UvHRObc8Tj8BYvwSHofkQD/DrwhUui4W2PvR6khJqiSqVEAFkSuuFOts3qKyopR5FBZQ8QtJke8q
e6T5g9HqsfNoFaTEX6uu6q1kGA4vydhL1hYieD4ARQUx67l5twhVo6idUdh74Gx3X0b1OiOq9ohj
F20DrcZom7dsqHp4TexI/WdxAik8Xjo5jfqJDGuGlwXhPfKJQl3qoXmsVNgqGVsNgHxf5ULNkpso
WM/bjoN8aptr3ycRgNFzP1iec1otM05QLNm46JaMMXPhtVIRIV8SovNqKJqkYCLiUdZ86pr0AODB
ZN8o0B5ryHQLe6kEap//x+zn+wF+fftDevcN6ZoS65A1exklsa6LgNNI0P3KOY8+zu4SCbTkS3cf
InhFWS0/kv4L49WGNGc0vuo+RdSEqowIGWNpH/gGh5HHPqG3XbZkVkX3oCOGFmNgpkoXqJ+v0Ili
Op2JgME3gCEiSkMhAGk1bOmMzh5Rg6oaoWkDa2V+DhV1aaZULwnlklW25acQP4L3IzFpKh2V6nKu
B2nyGZ6TggFiYR8kVcIisnXaEjo9W+kqR7LB2TCViVAvgEajQKpWbSmEiQB6VgCq6teYsE2pCb2N
FR57YkfdlyDTvjWcbozh3ik3FWViZC1OPow9hsmtQ+IjrGbiz0pq0ntP1qQWVFJAYGEeJ+2lLspb
vUeqVRVLas4yT701Sh4YGinKjcdqtyfb3PdW2eQGeM5VppfPuKhNjW9sE03tFaoSXCBoTdw9W1yE
wUXXaETbOOhMLgLX4MxtnbLlabdoYvSADVdVKIiPCY8QKZ2wt3BWGe2DHfmYhSt4ufF/bXalJKX1
SxzQ9R5bvAnhEHTl5FkzXiARPUX2E/tAP4xZKqpkVss95Y60zDTK9X1ck3MSLfT9p0PgPhUCRAY4
TBT1VgIJ9AqT5eDq82m5BfK4LY4/28NZqujsbGTw2kM9htsQgq0yzUCuWfpOpC4UtMFaa4vug9Zg
f7Em6jnGBWCVvWwAAPBjNUKAgDpnADtdd951jW19ibMdtSKXM54CkqLb3523OPKgfGGPgr87/5jZ
UuO4c5spXMrOlI/0u6PBrBh6hWGT+oDSn15sHZvsdOQYuW3+CuqhUp5hapdmHFsPe/4qFRHll6Gt
SdBWHuKNcJeuTX6KmAzlthR10O3X9CqQ8ASg/XBb3Sellzp7GKw7vadUBQ1qME99UO431sc512Xl
t1AUrr9KTbviJ67e3LvROhaP+Mt9h1Af3JMApdSYVdyUlcss2Dw8TyiOGXbcmO8QzdqWwr4L0bNM
Fa/itj3c1YTV+PRGvB1zEB0831K6wXCmIwWDA5AVtY3Jb5PHFVW00G0NRwWUdi9lewqHgzQ0F6Al
bVqi2u/Av9nmn+DgfId6/YwNq033aN/X7S++knXkZ3zfeZCun50XvVIt5P9wZ75xxE79IEYPjt0K
hLZ0dnWd++QNzd3lHMPIx5Xy6RawpaDcoY3KHrgWJ/nVCHEgJ5L4VVc1osxuspJ7OJf82NmlSnUP
nVMSy6PjUg8ex2nJO1yLdDxVeAPwv+YUfM3TKkR8oq7FKEreDwLXlYfFN/PoWWUeu3ECV0Bz7bFM
k6NpHpqplFvlClTzo5NEHp4gfZcDZ/irXp++utawV2LCwMpMmnFmoEwoMnJxKbbLw8T7w3xdbfHt
Q2xeY4E9mP+vTw1pDUQuvnHnmDnc3zdfBC+I5KmxD+UBJTcXvZw8krsBnkLY6AjX388AcNzv5Wbu
dpkFZRqkEu9afA0p9SdUTBBbSkgYojjwpk3ABoVo4Yn+S7QlnIycZzieESy+BXvCkk/R1nexIbzX
ietT75Gxr6JqEZR/jWEObL/tS4SK3Mv++V7W5qb9t3G0X4TnqIzMNlQvM1k9rHmiXTKinRDHyJtv
KygdZz0+z1L9OKoIFnbXrwNiTO9g4QgKOQvnmuiUrhU3qEnsZVH9kO/YuY1RP7nzGkzOx9QDBwBM
C90KiofbNHagukRPsZDg3T7UBDxa3XSHoE9Y/yAOscGLWD/t5+N1KNvwNtrORp7H/D49499FbfA4
eaLE5FaQDd+feh7IajZLNbwExOpHd/67FdZRXFC1HBafOeqm3a6Nb7DTNsEzosFXKB6gEGK5pZlg
8IZEaJ6GfxETJUj0TDuNFmEFLluvw6IBCC9wg4q9GXF+aMzaETA4jNyNwizj1tHxvdUq6iRblrhv
r5z6W9ucsJRHtTYvbsNc+fMFt5D5q9jjYTzoshsAZCXKaDIaXPBArWPCkLYpUl3E5IuGq2Uhxxjt
HowP8SzIOT5t6Zp8LlFNkuFzcADDcL8/00I0VVjaBebROy36JZ/6a2gPKYqU8iqteszqC6ZXiuhm
Xwp8nOtAPyv9TG/eou0D34xvGwwOCOdkJOWLpKSW282J9qe/bBuNzMtRI9mhYf05powEp8u+1INE
ekIdhBWgBWb3HC9MFgEUQoSTmcPFeQAkvK0WanAlAhNENOwVXFgbxKnDPG2RaQQbhAnm6w8AHkxY
iUqWfOgWg6CGEy9aEximaSTU1tM+oZUgKyl/9TGKB3xR8fRiBuPHb8auvNwsZcDP7fuApojgFkm1
lbFKDMkH5xFMqzNfxxQkM4Xy8l0V7gzrMarJV5M5hEsY9AtFR85/VAx9zBkYDhZwbMjV1Im1krTN
BcPbXAA4DlWdfHzDKZ2EGRZk2GS1C1Foseuz2hizcA84Z/gAkIMAsI3YyfRxx8sgwXvoC+a2gumH
XuMCYZb1VdJXZ+6l/u+rxz9Nxcq8FWiT52HphudC56vXusJSdcQ7Lc1TWFYRWvaWW8Il2t63ut/q
vVKB04hwJ+1KwPvUo9+xTYjwhKODkYxTeKuEBC0Z0hdPaa0SHltXMTjf9PFzHMDSoLhYoTIv90nD
6vFlest7a/XQQRSUMiNqi6cd1eDxi8oR3WVw4taSegA40vXkbud71/ahzwKElVi+G76/qeo/GVXV
w/mkxt7i6l1HWKETBlCsvzSE4YAkGU80giu5MG7XlIClGQF7KA6gQOUFFhW26nBxMCFxKlRcQOYP
MZzxngyB0fzCKIwMYNZGhBZ1boCiA3zm8nPST98AhBnR5bJPgH72V3flA42j3q1YlRj8/KfN3psq
4tpW7S0jllyf1plyZREVN3bJwR/9hCijPa7Q88bQ8XDLldGPUj5MaJup4W+j5//6qBbKzaCIn6+0
DzW2OCPjIE9t2UhOLbK/IciW1vSx7E8iWxKOEIattLxWvLtQuhBnw3TlDBcvTK0TviaONjE3qq6D
B89lcBGRQ0Kd7RzTuFpA0b0diSjJYWVyfbSUMdHar8TcrlwXQaVgnpkNs1EM4/BXOsvmsLIY2Jsa
ZjTEVb+pAQ+wn1NmSMiWJTnNzEJeNV9meksU+FSfdmeY+TIzdnyi1Yrgk1GGPlv8K5j58dkUjS4T
fz0BTIsxIo69bCoeKk+R+fhq8/jT3J1TXl21rEjh9qWr6lc1gboYgkjHGy/VTesNjFtfeuAoL6Y9
jvI68Gqsg+EH+ApDFpQUAUCqDyBmb24LBIr3loSujZ+DKrW8Q81nQLizEoLdmMpTCnhwwBC1w2Ge
3ZZXgHYjVyzfb36dvMuZPRDlrv7G1VqS0Pr/PBbQfk3kC5WRg2NyNSwY0FtrGnzTJlSNaSzFpHQb
EurzT3JBHj0UWMSVrrmvbEPGQr+Km7RllB/Kjg3RUpCoZ2jBz6IsmC8tZtZ5gcs1GtX1ExDMj0zf
do3SzALbfh9RF9GBviQPGR47Yj3jK7LLjbZnfjSFzPVBTcD8Jumxl2gri2ZjB/VzRDSasmR014NK
QYSKS61MsX1lXZHJsCQ11Q+tapZhNN8ntuLdD2bILedxGil74DakakH5UMLJxUaMLQQy94tfwybX
TT4M8gnNbJi/EMnMr1WKSHLR0IbB0b6/l3b7ygSoS6mtGTt1Z9KLYv/VOtT8X0JA1IOPLAyttvdO
zRjTAA8c877KER2gZrevSnQjiDHjK9Yk9OIEoI2iWM1i4Y8G4RaTp1jfJwU3G+fYTD7NzMjTyIET
CCHITlKVKxwggZehHdj6qGZhKoaUJ84PhThNVfX9C9TRuh1TC/jiIiUB8c8SVQZpNipMfS/3AyAX
i9m6G19R+izFdxpn6XuqHByLTQRKIEGoKeRBeDj2e3yMDKG9ZC5derjOA+IGTaFzL5nWw4iZ6C2O
XE5aJMeL/inWheeXFbaH+XcBWdG1SymRdK+exHLhBDxWO78YAq8k0B8Ys+RH/jRwf+8SSQo1BmkP
EqSkeCUtiKWmbIF6rxLLJqGT3mccCMFuwHQMR5zdZ6yLV3hlmVR1Cs2pBA5sUPgxfZFt0TJGxLV5
+vfxLZI3ZgzbMN+JpNYx3+/QCuQXLIuPb4acLA67DX881ahOZpsXq7ug0pRwDYVUYrynnpuOQCG0
dbkqs7ywNhGk1J6ksue8Si4BnTSykkYt+mnr3VLv0HYt7CdbCDVMik2LiUcAFVCIK90zYdO6de2/
2PwUs94ZsLvUOmcLlBzlWtXuWlWNqIB07AG6v5aR8ygEL6CYL4GbZTLL6RhG5OMo+TQYdZZ2avCG
U8Fpj8m8KarIAU+BLiJ67wwROrlQlxt340VKCxyjqAxWn8b7MJvFRnEtxfYPAUcFEoOf5s6Pg2yo
jLAYEZTqaJsIC1wdwIYzmURipMBujgcBTnSHlsOaOsHDyzi4I+6/cJ8hr67h/aph9O+sjcGJRPVR
MT20RZBZpRselKBfn2msv4AwBWdffRNgpZsJiaiTA4yYkMY3PrYLCHPsh4sgvU0JBVYhNdPDQQUW
Bfj3uVw2J0vJkE7RzT0QbpZdOGMqmmvi9nasIkLkXjGI76+5hSBuVHWAzMU1Cj4xe+mBL5Qbqlqe
UcKZoFkkxTJiv4WHLgZWkCxyJP3GqEwN29HDNi9dOBZb8SWiuj0HgslF+x8MdHg4hMmo27cuT7Gk
zxzR/mZVcdmb4HExmh5XUWQdod1OIbvrauxvrp62IBrCBX7XXYL5ou9wAawOBrTVDCsEibc66i4+
Au4cGIXwQUhki7fItZ/YLSkvWZ++LziIyhuEsdJrOkZM6MIWgsRbSFtJFnF3fMgRAaWwF0jYgJFR
jPT6XMjm+QjN6q3s9syrOwucgS8pDaeWmnNe1VZrofRPogBThTN0GFQDMF6rgGn/mcwTSt7PfFAQ
WBm4N7b6UtygL85GZgOYnF4voKUihNFkX9vepGgfhztT1ayur74kalWNIeaZ4vZ5nZXXQPJrMYXS
eib8ygPHDzXOI6Y0LQimKzdBeUKIja3LpON0yM7JKrFD5mqhN/RytaXobNlfwz6A+O6Nh3sKmgw7
ZGu2jPEJhbVeq9VUwYeT7K4zvffhn+NzSC02fW9JTtS4tAizX3CJ+hZkpvWZWpUHWPSrPFsAqtiQ
OBw5H1Y2skkk18UvfyYvU47+FRRtUfL2afePx4aZs0oBLyl8uwrAKsYlvaqUWzqgP6d/bdeSSReQ
bsSatkZU3M2WdlPDie3tD/ontMmxiGzW2DAvdVHcARBJZ1C4SBaNWV3UQTjRkjo8LNp78bazR3Kx
6u7iMsD2JuhsXBeXnhpNSY1hEmhrzHIoqJmrZMQ5vbjW1K16UV7kRkstTa/z96lJzvXKc2rWEsCe
2zQlcpovUYRMEhwoQYJc7ITWnvT1eoyRfVuw5YTiOZFKwrvlAXHshO/jvyZJXit9bkjOCa+I3F0H
QfHAEq45L1ThzvzXrU1VMws0Y080PZ08c6YnqLE0y9dn0BuxDwUa9sjpbciGWiwGNMra/clqqGEr
dEUhLptfJe/mDypocwXG67hpjppzn0nc9mQAp3gyb6RiQQSCV56mEAqDGCrqitERl9/xC8ooCtd8
I+e1FsVV7638I8Cu3tsmlkT9g97TjBxWwO1yUiTN/XBEgQvLHJcWo/u9yPvyp4xBsHVccxLY3d66
3ygPiUHwxLMG2+9g56gA6Io8rwcGwbHqUbzrx3SKhkUuOY+KtvdIMZuinTSPvPA90RPyMLJBy98B
Zhn/+xJ6MyZWF5Nt5DlcMSlOYNk7FtszOoQvFsAGYE6x2Cj9rKehZd1YIvPJxI2oUvltH14zjU71
32GIfrg5fLSw3Zs+15Tnu7/km/vDx3R0HF84cS2zWaKFcFojbpIOi2qkXXxxmt8PKddmU4sH5In9
lysLVEr021Do6XTr6RLmIo749tIUfRKZRsVEXwf8DDvYGcNyv4OxE3IVM+1GU5rCwQUUPl0GyLWs
OGZ/pvWLGJnba+3tq23e3zDSBEIdq2EgiImCVC9H2Nyy4xRc0RRCBOTcV+iSSSIR4IO7wgsVXYP6
n0vzswugGpXjkRvxHf7A5FRa/3xojz2lIfHf7h8b3XbnK1/jH2VcDvFXznV15q/Yc9/XizHFTQZU
8HodXxlVAQXoZOyw8SuZPk3xLOm5Oxwb9DYsirQ3dLCO6Lq2knHxTEwiVHCsWefx2IXCfYiBc3gC
UXuUG6KWBQGg23GUDC1ucOpkLCeUkPNjc+E/ntjAxkzWiSPCuUGa8H0PSlzdAxNtDBIYtHvtnNex
vOut/YpY2gXaOeaEygC4Y/W1lRPH+6F93Tw5p3Mvk0XmDlSUjr3EQTUbL5UbzWKZmeHCxAVdoHRp
8cNEH7F2qy7j6VSBd7GjBExr/CpOioPCoPwQvKEuI7HMyTUy01l0Ssgg5i4rpTtEOtoecjQdKdk4
6ywoVmw03IWd4AejBsi6JI9Efufdtb2Gyc1NDVmu7FFrYOVsrR25meu1QMds9Sa9g6mzUWdQovBo
CtprH6ewH80u4A2q1SPOe5eCz6Dcllbv/V8pqFQvL5Ix37SRYjCd04DTqCun5+AVRy0wp+cQiGpT
QT3CDQjyqZzhbH5LyP2AJy1JfEq9nDnMaDASx7XMn85pR5anxB870bLMbxAyvOE6y9olPXBsIcHG
u4KbPgWx5LxnedD/xRgvQaFEmMW2dsXcZMWwVJsEG/eaG80s4VpIh5c1ZKHBgkfzWyzKW5jgWSCi
QbUPvQdMYygDSyTKkQi8KPzsJ/9CxWoLb2fAoFPW1eXO8kDQwTn3Eds5BW1hAEPizw2yrShQWD1x
Gyma7552Fu182KkQcwhLDqskc8mQo5aXLZ+ORQ61Hxys9PQ/as6Cw4cXvItSIbdYib50nmel4DSp
F3U+DVgR3NIFgQAjvYrDj82sc41yTV9sz7sxq6j3W+VGvzlLKNiENozmDJLjQ86XGyJDHSzSZ3ki
8A8q6fj/khnoaSx0yrBPeX/0jeOoUiuDvOhD40JfX/qoB7zdWKBRLxAs3tiyiQvrbnstmKiWLsgL
lgRpApIg7U6B67mJJ3JIiShHKcHXiOfxu/L2i9hmNT1D3+JRic/3lsr/I6xNBLmubb7VhCuRS1+S
luGz1gBdobONMvPSAwuU2W61SjIT46UUwHKr2UYLqghLFL0XAYGM4uLqDAUEdfh2LJrUUDUd6cA8
8W0XtmEJcN+S4A7XG6295nh6gdZUYkyqMytszpAxaqmT9RxspnNDFSX3evv+nnS4hwujQrHBIGKR
/jYEhcZSEMfOWlKNWTWfrSEJcempAomzV/oG6X3Hqxt2dpeihez4SKNvKp4b3b66BVmyhDZGA7n+
aypgR4lXOsae4sUHd+38sl+A9r26YubK/3GDgFUBbPMhR0XDC+vYnnoQTnnhnLx1BDsg1+6H7mrc
znKC/GB+awG3BHoIku4p2L2C75y55eeolS6cbkTgMjK/JdSN9OyEYYDlzo8f6Fd9WOPhDZAJduQZ
e0b2qYTxbffTl/bdBzeNSHXehZwZ3LekqZ+dGoHZaEyWHvGAbqVDZPOPFzQ82al2B/4bCRYTJBAm
BPEhF/aJtk9Ai2s94iVoMqlnxioq2z0KjCEMIuuByPB9AL2LIq0tdGxn4H6zLuEDSGEEuNPgEPQk
3KUS9uwVJNsBry7cfpVOkLLF+xkccrt9CYEDmUkp4crUGdHJ2mLBMrTSJGprehXq737ovxkjrhTv
WIqePNaGJbqJXcwAjYuD/sLcxySef4Lq11GFrwofIlALc7cMDslBf4PF3zSxj/6qUcjQPOdFCjwt
0Jrm+DcYprxoGr9CHvXqelEhavV5cWMnDiS8UT51zM0HEywA1YrkAkTgoWm6HnFc2dg4G8ExvWFi
SaYskTmhd45sDXwanjFjvknElPOAQ2i3yCqDFXQMulrdLoWBb6t+q+bUv+s9G1sLP4R1+Z1oA9td
D8Wo7MEExDLOKsslyarYpYdBr0YLNwmcNRq0+OqYaS+hJyZA4zIKWFQNzR/wI1s6GCm3RdNZxW3/
X+s5lvgWGeGl4lcioiJQ9WEfIIuEFeoejrH+sbRdHwcg3V11GuaTQWPN1isf3MuVOk0wmcAGGukR
xh6Me+5ANKx00AWRmvY5m7s/e8DYm9z+2jTf8/lZMuee8Xp4BBja+WKeLl32DLsHLHbeAZJ52OVu
5MruVfe+YQIc8SDbtx8FNMTbnMou+75yzyqOqf11tAKw2oUvDdweNi0w1oVDVGBL3cP/zgQNHTek
eFK77KHXs1fjGT3iMBRyBwHPNRT4b+7A6F5dUTshewLM5vcOU6kvHwRk+2tyFyypwG1APb0Zvwai
mKGKfpOOj7DP2Jfu3akvyj1/IypNSIqT4YhhI7US3x/FeNVGNGfeK1+pu0C1u8pnH5xzckblUPyZ
6uzs9T0atPDuh22GKGh+XYn6XwTX4bzna1Zf0jaqLLlru0u6v+9EAMUTzenRN/mf9S7ZgbbEVd1Z
JtVM1CvxJ8G0KRrAVNxEhM389tIpo+q8htgYE5i9S9y3sQkJX/wGVO4Bs7CxQ+kMTw7VV34m4Pze
xnMswri6vLUaDGkP9mycprLQFnTbTkmI3XU2UYzK3zDeYh/tzVCH377XGOFW7dX0IJD7ODZbDeaW
FwFG8sKBi+QfV9k6DxGpf4w7LFtd9j4prB66ur3vTdUl4tYmPHBKsaW/sDhXkfrVWUvN+HqcPepF
yPmtHNCGjEF3eSczVmbc0+r+WUhuRdV7BMZBm0ru4m36qf500qiaUIMrFiX/VVlyoFCVRLyqoHIH
WAG0r58wIoPF5Zoq/hkFu/xa/cyDGdkVrv1y+R5ecq2lezWQphrOddxEpdyVJ5fiklb963B1WCJU
OI1a25nacDvBA0agQ8roal1nqneiid6LFx8VH31evhqXM2Fl+QkN3uFx3seufLuR2dn9BFip9i63
wcydqwocE0nGhk15D0hgiOilgNt9iwUuPFoed+i45Fo6yDdc5ZUQ5yxuyKF0+GscywW2X/vH4/Sp
xYnyki0NJqYfyOpYq1rK1ID3CNn2PJ8i8p8Ci8sNs24v+RU6xwqVIiQOTxr/B2SbYC4WUtpNi199
XHlHfbJ26ziiL10trVNlGbpWbXJTvyG+EbBknOClFgofG8LxOD1CI3/nlQ5F+0DxJdXkmI+OWL+v
gNooI+wdEAi1LHL/6kVoDcKpfxcAtrFcjyLMzOOj55R8a56JqOb27ym7P1u9JIQH6aH074aQbZvc
hHjYROuZ+p8ZjOd8jCQidjKv0wkUG5SXH0b1ygAWT+klelCSyP6sznspQgOXZpWJsNTBu13fiXSL
WDABvi8CSphU9sugDgd0/QbXjYHW5pl+CD1MeGLTN1npL8JtxAUtR0FzzTmoFUsA/I8GQfuKneCx
sgE9fZb74hrOKqXPyt7h1dDKzc67wiai2bVBBH1/pf2NXtbydjRLawKaF2pYUnMksJ9n7Nxt6sEs
tgd5ERgHbHDvWVgl2iU3ZooGc9PL91idKH+ulMYfxee1KrZC2IhQ7RDqllgOjfXEeQSLlp8rtQJV
IWgrTloTgnu3s6fEq8jb++bU8ZpkaME7gyY0gy6I/zAiJOJh8p7gti5qSmHKaMmu5XawNjnTHB4h
CHVt3S/2avNbJ/IEtfK9m/KhLM+0oGj+ybi6XVLxp5MSyOSeMuLhIhtLo+AZOoCt3f8D5WVg7lpb
tJhKdczUjGsfZ6Wh/p+lOTeMkrtxyVGaU1khbfZNk8ZLP9LbB2QP+163p3B4hlCrbXcLOPcCRHzy
xMfwwnptbiwPWun/e4aLtK4o+hlix1oIU9u9ywjNM0ChlcManmPSxxatQZnrfkoJU8opObeSfQNB
oEWA3pQTqVFxeOOHEtt3Z6h5m2ZX4cgSDzx+5XY7BD63maJK9TWo6XJD9y1pQxCiT9B8yKRs8MPr
lSr3JIaZYEvif46JHpGUAJvtNiUWUAH/ImAURlY3Eq6GM+D4hlORW77w7TP7bE6icRdf2SOiQ/Hb
MTCBxaZN+GjEr+jmwXuES3zDY9LE39dDwH5uisVZV29L7sF5aGQJYz2NaD4ajHUPMjHqxd7oiPFO
i1D1RmrTe+/fwtgpKlq8qk/w5YhMXQEyIDlXd1VIjYSs1fYQ5hgo1T+IPP3UMxfehHpz0Sx1dPVB
Prm/JZK5piwl9zOYQDn51ZvQmhWzMwVI+bsUKLV7xc0ouRGbl0KjP08QXRhaa0OsnegBPB23XQ/I
f/mCgw9HWnhgNWieyAGWuoZN9QUXaYvxIs015pgOdJrDhMU7aOKIFzSRZfr7uG7PNZUyosf+qyXj
XwPxfVrp0pAlKEeAZegHNwNKy2DYQQWBFHLhiZ+vVIOclu+CexRSEJejbEtf9/bSyA2xfQqLh4Sh
R5IYxfCyE9tTgAIAQ2iF7ICAqRE3Bh/i04mTTHlCR2UYmyCKynAY9t2fV2uOMGqQ+UDAL4o6Tzee
rciXElZNaDDTipWLkL/6wMHzGM7D/olqnlH8png9WUeCMsLz3BS8WLsh3wgpjO0IuSyJJdN5xUGA
yimdwse4ipCucOHM/rx7WaG4P+J79pZ8NBXUccx6EPPMaGJYwS572QdG0DBUPjT7CFhrkaCtIEf4
wT4t4dIanHCjNA/npjfPBS0R9wY8ehvqPxbvCRD20O6VUTq5AXL55NeM1x8mfTKV1ReKhmKfFuB8
OFXe5SHeAuWneLx8pFJRLD2iTQjpwjzM93P5mVobAMl4k6fEasiGAB6/0meML9Uk0+aGZA7ukpA4
fnJBsoYGoAXEl3owPpMUMmjs2kVJhDP70/kLMZgXEMs1cRAg1GIUteOvUVo6jwRafwdkgUqzCkY4
P12wvYVL/U1od06K+Sia5v5/6jrfRA+rpf12PEco5CJgciu3Q4VC/LvuQGazmW0TlJw2dXeiAIH3
wyHH6KUnUJhkGLCyhDsIWrNkv7sbelK6d7uWKtVY8KGYUPQ2oZApCFZGeSKjb4Fn75xTEuRElSTY
uMW/9GIglQQILENAjJQ20UVjEJfIybOfVfWvC4FknCMK/HlA6pM/5sXEod7McIvuGETeosMsCFpF
sWaCKMwRajzdGXsGNFBMcWHpevEwnuhDxr+L+BGppCkKA7eAfWf7hzMr7UeLwd9NoHtkqWXUKrQN
lQIH5ziJnmdQ7N63v5iYHu9W8+az42KQL26KY1l1xzsMB5Pol/bWUYxEYqwho8eGpUiBi6LNutfo
TyK0dYxZsOJ5kJu7pYzEcMANnXZqYZKzjhziaijHxyHrKL3uC5TyY4JviDfmXH410v2zJYWh+iHL
aAKTn9EuUVGSaN+tMC5zvVHtzN3F9C7e1d/6HEOqQH9+Yw5lg1UCx9GdVQ96Hi48hx/GUQ6ZGESI
R5F5t4BzdNKUq/KUPvvZG1Z7LkDRmDTc4K36cMmcWRnDYAXh0YTtTvgvxI+S2CrAZQCvCuZC74Ha
RF3idnrtebDAuLxFvqiKdmzA/800Nhso4jWciHEokIbOv8u8quChyOATLlMm0xI+EMWMe/9ik7sY
wEMNSohHpR6Clm1dT/T3g5tQp7eDwRKd5a+5g1xER8gHJq7M7eVjmdIuJF9TGphZRWVpT+lxPcbm
3J9qqOdOvG1mp4VDSM6iuJ4CMDPRLMfkSCv/uLkEyLOKmGJ+NUVazcaIjN1lUqQokKuiYJtgOZCo
S63KRNzqZBac430cAyr4xkqsZ0s6QlPeysAcf5WJlsQ0PDcd0heMNjyyrdshLJtU/PJ5fc7RgplC
3p3aM7lAjOCuNjvS05zsgH7PB2soGSWo4bauhydYhMNnN9EdquIgus5fXHa58UQbHF+WIy4yyLnY
gH4+f4Gf6clG2TTGoAeaVw5yd5bWRZZ9h2v3ZQ6SkUVNlPokDXzqYZoZl1aQoo6o3Aq6OciV0STt
h1XDPtku+6SE/AUApcJFH/f8mo/tuzme0c7lKSUKV94QN2WvrTAGsonngkk7o/hL3ODXyTTKVTci
csgQnNgxy9PvnEqdxIR5LbEMKmMo4MeFYlCmeyjdEmssIBlVPPGevg6NqkXqecwnDogN9V9+cxqu
oNb1qtd6kb1tK4bZU3dJoxvVpm+/lVyHtJZ6vy3lP90qSl8+oVLp3zA4e8hgBKGvAg1c81LogSrU
27VNkNk5Ee6I09XVdlaDt+KSta99KZWXCYi1MszKU4gAQ60fv+Pl9o1RrHAIUW4yf0OI0/ArJ3bJ
0f6qLqOtVcXSzvJq0iwEtRZDhSPGZ8YX+vZERFOb5HSLdcNXp4SB0Ya38dAGRBHS1BzoCJbAQLc3
AT2S9k15YBWKG6FhBDOngoi2zS8L/AeV6X89ewDJUHJ+sRk33Oo6o4ZhnkUB/LzxUhCz22488hL7
XPv2yAVlF/NKiTzFOqb2h9XVNX3T9iiu9N2vULIPPg9FM8m1iKOQ0BHPc/T9Twml2BfJ/7UAd2Ob
ZYwaGQJuuflQaipZiLdhHj96KERD/I28ZtbXPqujlTLIJrc8tQUNWrZbQrbHhFohOhc16ghIkvgb
ZGOHSb0G2N5YvfGsdZl4FTnBKTA49ojg/fwvlC/GGz7wnwDrLRfzZuvE7FDYqyrVDmaKbnhsmc/9
ZWhHeg9EcH4pTgGbcvB8TCxaji6F5JzrdxZVOQcgwWxg8K8dlV6HmPEsmvPR1U8GcEA3XudwnyA8
4pqMN/iO6Yi4vJyLuJ0/liEP8t29yeD9hZDfYkE/kF0i7ZVm4kS6mLAssy9uAyqyADq0WamyAUNt
eAzHwdQTwm14jRNLHNUMaANUIVzKDLBCGsxz+G54KQtIexf0T+d2SucnE9i6JGvWK0lRaYajoIin
U1yu5FZQBS+PwySOgENqqvMKsaoDmZklF0DOmJZ+mP0/zQthuKDpmPfx8WxzG4cNbMHu2J7gAvMj
2l3n19I8k44H2q4CaZh/PXRkFWLCvo8iMEzr+C+/89dnQN84YsGW3Ff3CiH2/9vH5jNRT+ZJ5K1b
S551LWo+Fneg13naVy3f0LY+DPMQvmfTS4Y33PfjG0E2Ixumpux4tj6K0Tt2sunaLkUZhoRi0bk1
0RQiQ/zbN4KDq9umsMUQywCCSxOPzU7RAIYZR5y9JACoxq7daE7a0cMDcHcWgckZQYso+4FjRPvE
Ggpllao/Pxz2o2eNECBkFYbkKBXMHPDyKSipAgp8Dsq5cmEpEhX5YbvW9zPeIzZgooOMx0vgT5Zg
rSxkjq0KJm6lpclDzOwOrE9lul7MmqPRz1hKfUmhb74SaX3dlN5gxtFfY9C7btx8UT/j/YOAtqog
vu29kxjzJOhJV5Fld6+1XapRwFeEHVMzU6Ck9NevSwvT9+s+3nFs6BZTUWVymJnqfjSb8F6xL/44
VTdUZmr9+kJdW4qm9TcvqBBNviwUD+I9xLjxZofhFpI7ryJKi7Gj/71onY0hIrPkLjt+jJuF7oOo
Fdf4JdQS7r4EQh5Z9giG8Wu58clsfqh+UEoU+ZoL1KZMKMz/xsk63zXFwjQSr9JVFa8tuwJBFJz1
nfQgxoMerdPujjGNBV5esfXDY3QANzccpFlNHvKzM08jvYNdWjh9LzPdYSRSLYoAEtQBYhHNX9lK
nNB6tWnPn6SGO586aRXMDtJt9Y/HrxcNdUNLO6TfYTShIC4OiPuQV+Tb5wX7FR27OUMaz79c37AW
+Lez1S5teI6Y13N8SakxIrJBn2F4NIuwSu0ZDgmklygC4gnh/Wc+QPHSt3bBHj4Oo4wzIJtOILH1
4NIQ7Evuy5I+Vm3n9Y3MVw+H+tHfpl0Wn3h1uM2aYciqzlaSPKnkwcyLd/T/H6GPeaDpFM2oV/GC
6jPznw+hyzjQAKFmdAg9FqJHmbfISfaV/vQAexXd75OjaM//jyIQ5V8dklgRgZswuaYJzNvQOc3D
n/L0K6Jyi+8rDTnGY+gpRRL5Nu5NgdKbkm0YU3imSOfdEW9k8J7dEeFwc8HDXPpKi/5zOjjW6S5K
kujTZrR7vg+cZHi49ZjTL/jCmrOIA+0nTqC0LQcR7gJ7T6zUtYt8jTPvFjATd4q9ywIjlO0LAv99
kbYI8pjj9kDDYgBkMZXjXYcyEIcTNk/ccgHsjp8Hd95S+421p691yGXVFdQhPmcDrozWsZ92vjlt
lDTHyIOhnYVK/70iC0/hJE+EPnYKpe972NI6lg7pSLj4/AlWMtkjjx0JRlH+NHJrxf9pnmOfCjg/
EqClrEae3+LAPzCaqkqgwW0KjRObUKU6ng4OfnR7Y+ic2qzDVzj9/rWGILe7wnHRu+cUUc5Zmt4i
a/tTUz0z92Ky7tb899/E6SV0ArKJvn/B6iXma5MtUtHkiiv95qdmK/XKmgYgYsIh8nm7GxVaJz2q
OJurUc5ybuhzBw0o1atAlpMRqnzJKebYH4XroH201K1UbIKmgMobsDbNfnzPxO8WWELdw/Pi2u3n
TbTtxjerHdBESKf15cyNZ1Y8CaN/I1euxDY10kMSD9EHo/4F9VoUTBJ4V+/G3sQMFofXMcmCKVoz
I7z1WuR4WHZwDP01SV9mO9moqcnxeEsFSSP75zC5CjILLVzcgZrY0ExB+ni0wHNus711SG4yRiCa
keOP+a7WPeYGA2/+bV+mwWQ58hO9A6V2gI+v921J8GGBXxu5KVhvdgB1I7NYSyGqHE54cgQ7SqZc
ua5pHrZ8LbL6Z5gB9v/JBFXHWPhSxSFQqkiZuBrFIxli+Pb+TvLrSK8svNgFSnK2zrCv8bd6FKlz
qceuHAK7esXyRe0YZ6S/dou/efc05h9oGBYXmmmkX3i0P11zG8EAFsMWz7pTb8c+FxTLxGtJtsBT
N7kaFaKv4SbHMm6qpgKDzxwrNEg+uVYfzFTgKiUucjdaotFOFgzGiRUcRIg0ICEogP8Su3vweT8/
+8CwsLPWm/Q4Udb29Ogw/r1KBOVY7Q2LgKv/Wuq/3x/f1NicHIFzdGmgyDcmj88zWF5SVjoOSIs7
TDoKfEW89FRaxmoS25/K+zZPpdyl2Es7dbDpDgXpAFs92FnYJBzqVhQR7J8p8PrO9gNhtxktBhFi
5MqnAZiM4v18ZV4zXZ9y3idQkLBUS0TQqxh7wTRXJnh6VrnJ/7TscbC69X9ws8z3yPE6Et5H8XsI
7wkX3oUJGCEI68ezTchFsTP4gdT9EPfnbt/xHhOGPs9anbwZ4mdQt/4UrNPbCTYe00wikAkle4gi
3zWoAChfsxyBg5p0W4WdpPR4okpP1aOOM2SMoBRg73FiT02ZDH/TK3573IIRSmpxWnHmGhDk6Y5l
1zI+AoXyzgjkc3rJqTy3xSvipNvl4zojoBVQjplKCsBd+5f/PJp85pWjlaUA6r3NGVdRbHab+Aa8
vLGxGsbN71pljs72IqgyZ1oI7t1p6Zne+LUd4y2WDWwyYDyexBoLN94hgS2P49+ZO8ev8wGWrOb+
N0FafmSqZjHb17BJaZ1Nbe1r0zrfd0ARFyLkhzcCSn+CO+0dpQnGGxE16rTZ8yHJj73BnqbSKdmU
tnCxd19UC1Sv2YeMaJpx5IAB/mWsL5UrnL1sy6vrc+HoyCGdW4U3mnq9nNVAYrY/8x1r2EQJxsE/
U2tiTObaED91gtztIOivY0MxFmj2yvnfKYvBe+0d1inLuL2qS8sTIb3vXBUPoxmeYRT5a0aY+ine
xjLiQr+o1ileYc9xCTgamynkSP8PTgn+2Fw7OLoP1rbahUNYOCE0zGVpSWD198FqZKfjmj83Cq0T
LKqdDDRI4v7NMcNvnLOz16VDY8R/sSRosw0WT8QGFkVtYmZCrKStFj5md/w4Vo+BQMt0KwyU+FsJ
ovZGPvC4x2AcMT8OPHWwmKoIxVAI/P2dbdfVMBusnKerBPWwcEKx6zWW98ukYSd98u+m3cMyhq68
y2QP65Eyth2fWs3+JGJKhMoWU5TQUV5RrED3UDRfxLh333WLgtaW6GU9PscgM1SIqIa++rHHOMlM
90lMP2aEfrtkNFi3qlUA6cdjf/jDX3++63VLRmwTxjAujVGZaUtvGaazgEEu+ibRCG76Tg93dXmq
Wm9FEswisBIboDnRa/Jsgz94J/qvcK+YJzxqma/+zl2ri1PXx21YKUs7uSgOMav/y7EdAGQi5qtl
0yMD9bYfSANDU4G9qXxcftLdUnwkYPZ+4e0tdujzdwwWIKNQUV06mSUuaJoB9lAeBhAeEUNgfWrg
4JWaKHRLSDthXmwEBDdmj0VZbh94WcAym5qobog3HkfC3YP7pIJT1UY7axo2/yEZqAkeSmPdGddD
lJnIrBR2TjhMlKmRpwsK6Ukn3nPdrqtrtHDRtPmk/SCbumC4oP7AvAXNNJkptxQQfoGBw47vytvD
05P95zEzuHwhL0TzZUgaBRojtAh6USW9qAOcidVnnilQ8X10jAIrhaXzfLD08W0/UabaMT93D6/U
UPxy2BKRLuwn5ZKloGb4mtWZ8Im3+h+nD2XWEKvK+MUFasVIJtaupm8JNOh4krjtaqVJAlitIEVm
Vcs4z5aYtGLGIOliMqKRgL0saPlpqKLjxF9PWJgNP2inXrZsHetKbRAFgusMdVwZKMaxU/ui5RpF
9+CPkTHt4Qoa9X4FLrhwIiGy7S1kVKOMRlQd1Sr8SIiSy7qzjIPf+ErDw2ke6qDOuBY3p6GbmBh+
2+AFsnrVzGtFrOGJTXVXEIGtQdg2rSaiaz6OgAP8AfPjpeCq737dEk9pz1Wt/Zz3OLr34oUup+B9
TY9XeOt7Wt6d2BtrxkjbL3pNKOI2fbWTdHldOSAQ9PXxhOtldB4jbFjudbVb6MDWxCOnoVfsO7rK
awty8DXUM9Z3UNY9pzwB1PlQGQhofXLwNhYh/ZYiu10J7NSC4SRFrC7OG7BXKKcblZKiiY6P1cTz
TleB0T3DZGFwueZ/AN2yroYlVM87HpBlBidf3T16U+Tv4BtJ4hdG5bn0mNPkC3Rbpm1aociEzGvj
D02dV/zoTA1PL55YC8+jr+QKVwhzW6sUjyf3mUccgVJyfeOlVx2fsCd/cZHEijHNq6J4s97rDbEE
D2tE2FwcaEK4fepP9JBQsOK31GjaJ5ej3zOWZ6ved5kxpYq9LgoOjx2KO5b8LuhWQ9TnU/wMrOOU
EfMyid3eQdbGPzNIx3o309crdXY+DHd4aUuUBepziAOL023T3rp8wtnd81i3j5RT1ZDktDqIJyt2
NIVrSSL9nEgjD32auU3LzkOnaAGNn1U7dq4GwONCRN3Yw3Bdn7i1kgD9X/iZOK2T+jDtpbznAeeU
l1/OOoedJbelZlslpN1nzU/V8vEmzAio98sofMLeR4iLNumJ1GoGxhoUk1C8KXl80jdzWEYcUWZQ
/PKXulhNOJl8BXdG96hHhKXxKAtz7XgIwyQJ3gDPvUsf4N/4iLjAcPmTkdiWmPtKno8DB5hpvE4c
J1cv1EFBz+wabcgVLiQMUkNQMLoQUKLgW5dLL/FWI3olLRK7q8sluvcHNCN/bY5XP0QSvBdKztNB
/4GFa8QCBnLtrmt4B9e2QBiTCtRBwRjukLvc502XA+WHuTUYJsRKbyJLv6H0Ws0PP53cxdqxXOml
MdVOXQvAK7NXeVLWlXrvI5nAAxWEtw0p5OuAZ9fqAtRYNCYdnXWjDCWX0D+/Xvd89iQH4xVnT6cZ
cf6R6ZLQHEB16wX91UYfMtjK1cMT0MJQ1ze9R+razT4LFY8n1YlkhRtXoBIRB0APay6MahBilLmS
HPY5NZn91Grkcg9c/A3EnR4P51bIZ7fGwRYZqxI39rjd3Wwsv01Xsjvng1Lk6T+hsWwPdgOfflZc
bDwnMZ+1I1V26Plq012EKa+GmVgRbqrZv32CR8umv6lNHYdQeMRhoWk3kcLXTlCDKVgxr3b9wb6+
46FBaMdv8+QG3KJVOIrT6ND+D7uiv8St4T/ga1OVT8I8hdExlePCPoPfT/S4o15BKCrEhr9QgGat
bPiPNQ8CN+Cp4857u2n4pzkVHihe0lTkx2evKVaQZ+JuAig7pbZZNI0ja/iSyryrDWsdXeVHCA/q
LtFQk3EMe7WcBzPjNqoRNcg55Rh6Kk7O/sLwSL0+njhXw6AMGPOheRC3OH7Ep0kUt1V6GUYMzmFQ
9B6uQB/gfeuQcZaGCgdROSuLoWLG0S4jmV0+nTbGgIUyFZ8q/nd+jhBa5vTyCnsP8Y+jbYMEduJU
aDeMaJoqTbAzlfa5AraXHHl8BJHzswU34aK65sp7Sn7VjGV33cdVTe+pa9UFC9dNXjwV1RJesZSN
//hi3u1KSN+kZf7V7h2Q+RJe13dO8Sx6tnGjeBEn0w749LUtDJk72QQz5pmEQagPZrkrk2F3/GWU
bX946YUl1dYD+M4N2Ioxt9s0lrdiDV1Hnqea7OiGMBrefkO37EjF2Llwu23Z26O+3jyKqlpL0GkF
7PZdEX53YeDxRt2Bzb+nQm9ol+lwiC2HLT3h0phNtXTsgl2p6wx/0zPYF8FGg0d2ulJOKS1rDKz8
Qg07qxeFkPNOa6RQSPOA6vXGniQkdPxRQvCthzcdWDcLpec1Wm3Bfq1yPmL7M67DKdO3cSQ436gs
qvKgfqUAVRuIkTLx03kSYYPInhOVFb/gR2JcjMqKAInqxKkE8njbf/9nLCp8WNSqAZUgFDBdQHAG
k+YoA/PDADVqH3/baZ3rU8hSedpogR2Tf8pJkqbphJah1yGmHH/NmRE0pUuXDs3fTR+Lzmt8L7Ju
no8sb09/VaHnXt2qx+WCascMoXFFzpYmdRvgmrqRVcaCh/G+ydvbnTIFE/8eCxb17P59RAqf69Y+
ue+LrLZoaNa7FrDPRtLNWrWcjl+xdlftbsRVasQKh3AWVg/AslwlOw2elAdlk66qhYxABhWFjvw6
A96FdeIvdWgZzvtOdxJ6UHKa2z3O1jaXLNYiW6mUtnGHiCsPU+6oJYGUYcN3Gfx47Hjv248xiQzl
IbBQw5xcM1bTeh39SIafzR/BQe4nE0hTDjsgDcJKCYInuTVx/0EcdFXTOXlxW/kAt0z+IsuVYghm
H6GipvEEU53BJHVDmHBZZAA0TyqpgvaLolGVQbkz2eKkwBqDS2qZT86k6PfzdSIKCYpblnX39jhq
fob3uN3+Y247bVFV/lGqz2I9gVilL4k+Qe4rTFLd+ksTEFtMNQpOxF5mNWWe/8/JAt+FidlsnQrU
Z+LTNYzOtilWoIUB7f9LhwRUqNGZDD0qGJVwhU+IphE/Y4xgRJjx477Ym40Dyunsf101kMFSKQzC
gtVRWgDPFxVXLZEe1uSxdK3esTx/HohrxxfoCOvH7BVoVDzuqN9HZuXHLCKThptlr3jKgJ3FAeNq
eeMWljS2+r4W9i/jVg2x8R602YWZlha2SM8HfFMykVqy4Rqw+AN46it/Qj2s7sqX2TLyfRgk8DYy
TeiDa+reaD4ofWddsIDwfS0DlJkA3ZhwJERnKivYdlSPv18S0vpg3G7SJw/fiYyhanxt86hdRNY6
MbeOgIRrmrdGAY9OWnAFNJe4/l/+y6UPS4UbSPFLHGt4e5mvV8+YX48Zx6BNcMHq5Mteetv2m9gJ
bPNj2Eqay7dPNifp04wc4xOEIhnW270vc4IZW0To0MK2YR5vZ1DMNrnF7nxamHTuw+9CG7thIP2P
v0Acu72O1ScT1loANQH7H1497o+z7mNN+MK73iOMgGe4iF9i6o5pN2LjKyv2XvP5qsk4EF6ZBivJ
8SZ2H1g1qkD+uoerZwT//kQD8i9X2VERwEyeBPzElshvkUMvC9xNfRi0FOQbb0AElH6ic2QbzeUo
0eAW5Z9Uez7MhuBuyVj2Y0+sBmO2ngdW62ChufzOWFHt723wTrF7i7aiA+HS+1E4m4OxlhGUlP+X
iOs+Tg==
`protect end_protected

