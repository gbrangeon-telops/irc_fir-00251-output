

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZF7Gp+JQYN4x6Hvjz/p/glt8+Yhfw+y+NSJwSgFAT75FGfBEoCi9gxGC1aPKEYH1nKSH9HDVBmjN
jVYDQh69UA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bCrwACZO6VlyUjDp7F6NflPANkTfGVm4hgH/4AFvgK6LtR4U73r1HOWXfaKa3y3uaefm3opyWNhK
nV2TI2PpMLr9LswzFSOsgRzHCqR+XBS+8LwZ+lBVN3PhbED4ykAJBbHjWQapS4mEVXs8Bors5GDK
A5lW6VBcepABjdMHcOc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sWMXC7ertaTFiCso7MQnbVyuVSvzDQRw1zbA8jCBUoJcGFv+Da5uM/ZInIx2vKnorpctjF+RfQ/I
vLvHJ4hFA7ai3KLDBa+osiqXeR3vvyAO0dNGGmO7GQ1dYRUzzSKKrGTJhKWqDfnAsYaLroy6U3UI
uNSRIQtxv1ciGPzcMfrykPy27NH2CEGiCobfxP5HXDyrOVBqWAZuLaPzQRv0D8Ie2O70SiCDKawR
vbedGBup6qqgOpbOuoCX/zcbW+qJ2FxQY5Zrju+0WyLSf0XnZd4src68n6rXZlziL4eo4Q6lUGQv
gUEyqpp9Wiyw0QLmYTxtAKnwwMsfY/jCo5ZFSQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d4cZTzaonF13oHTIDZgb2oXxuKQXQmTrHOYXqYqbAU6BYAx+7y9fxq+NNlLqPYeukSU316ZJ2R63
uH6wrMfXFW1V94ov6Pl2EeLSPre3P4xtwdLCKbJrudZD4i07Cl6ICwNSN//h6MJD/kwUIU4k7zeP
ni9WJs+GmLVsVx0bOck=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W5Ic6b6KWpsR2htHXte3+6CjlmHZcuEa6WOajuu7k286E/JIlKxSU0tNrXH7rL8k7QTBc55tiAC2
sT6Jtn2FOqn9b4N96SwTUIbdNrh5Ew/7EjwCsd26VOwpEgD86kAwm7rEEtRCtStJR4p0yrbCQjf+
9+YuvQ3Ab1Y5fgtY5ijqZPgs+knlZZFAxm+NI7o8f97lEMTpHDonVgfj/KtK8xhV46JSrDB2FPhp
PMezRFDPcrnrGio0JnUe1oPbSneaSJZPAFIoGiaaxfjjDJIOa0DMtbVjecaL42P3+sAmOk0R5Mfk
8MlmwedAmXWwr0D9NdqrNJ68Zt9aVa7CXXiS/Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7632)
`protect data_block
q2MZJtwK12a29q8CykqPcnx8tw1FEvDCgxQZfOiu6TJmbGCM69NsAmIzLY/0eeDCd2kyDictHKx7
e1nc09Ztnjzc8apc74K0hJzA1QH14gOOV4QFHHbJ9Whn5nYgpeM+wPuzGIo0O+xsgas21ZpPm/1D
aly/9KeSrRD9bLX9oLR1OWNrNq8YSIr2GOmtQBy/Pd86ZGNCQzTf1+KU6pJXih0Qjc3pItig1FIJ
6H2M0l02Htp8WUOSM9wQH3XRGuaHEoGGkVh8opAP0fSrkZoVQlOQhJQ3/+PgvlXrYYiWryRPGShm
4ygOdNp8+2iW9h3j0Qx3N4h3vMmE8YyBkfua5JqqhBJ1OEvdrhHJTYtbXDvqQkUIGKipZ/24X7/d
U78RSNYvbqEaqKgKPl+TL/wz3MWtqxzQeOpl3x5nNNNVzJAUiFmzs6yATSgbCFZM3yL07g7zBuX8
2fCvYm07Qt+jsitQ/48iTOQLh/Rdbe+Xj6lXVZgu56fZtuk98tMthFeS26Ivw/uBNT++B3Mw4+4V
ild66Kma50pkZfh6HIdaneUuqXRi1kfXyQZinlbTRffWD3hJr543KlFWkTva8vnKLmq/DNrDZ5Mo
NN5WaZGL4g1hILupD/k3TDukHfp6bbfdBTSe3lMmYbC7vB/u3RdAueVzK3ZC8S7RW/Uj+PmvuPeh
6GR8BsMCjK79JPmllSVjEpyffsIIwBkSsUKDOSjQvdSXKaYdCh60dZi80glAEwdl7I1Ew4y1F0IU
hhwCpt1IF1BAN9ldNPtzaLyALHpyeFwo2a7oNs5hGM8aqqhyRWtDRq0G6a299gLvC38n7ah+bqji
AyIci29bjnIaFLY+BnNOVyKsRCo8yc/8MC5f6ov7GC2aZylaSxJWJsVbf3BVx9jOl/fXv9Pif2BM
XTEKvfamcXVr2RCIfWtFFDrmQawyRvM9+1mDhisn3HEU1YZgL8o5hvstJ6YVYTYCq3NMjWCCclx7
J3bj5cJkxPpOTRsjWASsOSBv1m1neeyM7emajFGDtI6NQd3azYKYka3oEmCH/WQ0e3tp6BA4pMmP
YJd7No4qMPxzaTooPf2Evjw55vi5fzoXuPyz/jD/WZBtHu9AwrrTkfRMeK6AUEyo/Ml1PTXwYpL+
//ZMtqylfZWFtwSch132PZMooC9N+1T22/UvJfLVklLdDHHSIR/2whkHCPWYK4VJTGiNiy0ZWiMG
Nnj80g9cOcgMaakRYS8YKxTIlYvtyGsIWzjS4s9y40RLsTL80mzLUpUGrOBArPSgiI/TMkO1SnPp
/Zx20WDDRWKC9pmEpJX7gtPGe79Y8hOmXzwbibUohlBOYUDQeYoF/h4upTNsBXraqabwLArzx4v5
2bzZR51A7YmgkCBvMmGd9bpvr9TYLj3eTHDLL1z3GPx6V0z8f6iOE5Nru4UG62skMQhSmNXkWl1X
+DOauI5G+rIiHngsSvESrhbbNTzZPi8iODan8qrWe46HpUls0MjIGJoKm5LfV+u8udaV3hEzASIr
n01oR3lD3YcnzacfCMyMaKAHMl2tjd87hZSZhwQCDYDlbGlAgxjK8SlkjVgnOtej9Srdn65eXomG
jiXN36Q8dqw2cAlEna/HdyHjC3wc8hcr+LJbW3Tehvee2gE78B8RxcChmnyAel293AV1qwOe++Hu
Dc1xr8cSzcX4lScJg1w+tu/jJahptOT6bepzMVicVH5MMrh7Y3vcApmPbVb3n+wikEnzXeQewD7g
6R8lLEIm9DAZ/A5il5Fx6bebzZO6diPUIU3w77Xav968AI7HuF42jxe5fNnuQEQ2IZ+j+uIZigEC
noO5BLO/+mlukdsU/P3gvxgG1Uq+HCkX9AAkmRemc5NYhKK1G1AzzYebRWrTWMm4w2dYaIHRhsrG
6JZdSME1dTizqeY2AX+YoUAhKzNDNeIEB+3Tw1adxvsDKG3osZHdD3wySSRR0yoqXNnXo8e90Mch
xnYyrHZYaCPy65X7NB0BgQQtU5FP/bG8jERBwFscAxQ+iO8P4sizVHEhj9No290IVJWXGWkI1rya
+DjyB+4JgsuayuhjHUyzmBtt2ahoqZvaIxozDvaFVq72GTEhEYY5RQxoNldzYFi5E7Ra1kSlLiTD
Dl87orvbMUt0jHaQodjsMHFcRfCGW2hvSbPO5sd4fTl2l3dAWc2A05eLrAclLWz56Uy8oIgu4Ihg
ZtyKYt/H45p6GBDsNsWt0VhczuPFcTOzhoo9XeLpXb4QG82IuffO6hWKAhygTmWkw8YeuZ5kPrqR
VV5QTs8xG43hms7ZN1xES1z+g3QUlcXjykzJvBnrghMSbqcgmBYy9g06XjMO4/6E5HzOawrK3Bz+
v+zFwePQvbLXa+Jh11HMIH3i2tReU/dzbG7V538jbH189z22ZtwwsYLYNZS3EglZovlQeTG7emoG
9jUt5k8cluUZYkr7rfegoq/0B/fkUg/TJ4R0e4Q2DWpcmMxAK44ByEa0zKnssbmfRNt4sdWrH+vt
1ksVZvs4s1dUYr7fAHTagBysOTMxd0tYNEevm2vnlhM/4v4rCARt+hUtHcyklwwYkQf1IhmtC3EE
As/5/eBPqlqC9NscB2jn1mndXQ0Ah4DbD7crJcex2KEOw9fA7DVk3YQ6plxgajnEHe7Z9GVMHDc+
Mojpo5u9JFWFuSY8JIhvbBsyq+hhnclK2I7Np7af/PHc0a1DFYK5QCXnuOeN9OWL/sIf0G41mdEH
pKQQf3rcVOx5PMkAYPjUR8qQZZCg0SVwAkd7FAzZm5yy5RzLg7muh8FgFnbshG5qEH4HxcmDcFeC
FqCC/LLpayaVFhuN5GaGYyymrnQAakdiDGO3YkHN9H79UKIXpon4VKzxoynvWg9mlPGuAVE5qnri
d7hQEaDwWmwLfqSi9xZgmWdYof2BiOwuliOHG4a5UtZNhUvfaXEam0bLP771obUHc3I7sOIdMQbT
RLw1zXBB30IWb0iKf/S/pbfS+O1/tAVY8/6YkoR7gaxur3sil+2E34nNhGjAjcDtfPKZL8IcNeIW
oILPL1L8eh8gIM/BdW3e2KMI3tNZkKvVyfbjLX/7Ll6gt7OOu2VXOwyR72KolMq3wmZAxw8bR8HG
GDOGsTWprINix1obin3fyaCyIFWkgbrIOogkX2BSdfk4tCSxRDillP9UmCcy9AGoyHHNUb1jOk+R
hNNRLQPb6w1K/Y/I7KxP+rg8CgHAB+3z029WsAQ80z4/0wPiCoexBl5+nA3gfHsuYoDLIbX6ORLn
H3rdoa240s66HZbn7VwTsOpeZwj0dwTdIa9FGSkEGL5aCdSCHq/v54ZJlmeP8N+aMjYjusHRtYk5
fic539CPdPVRUrpK0N7yw1HXbe5YZY0yGtlI0Ki84lJzjFErZ4unciL49fn63xTSsAyDCRv0aFZT
pu6tZjq3FSzsTA7VQv1cQGHIiqumbrTzPVXp0NWqBQqQP0Pr/tiTlbu0WjFHCCNywKsWkB+fNeUp
zpnrh1CfiZ3ICsST/z5EBpnpTe/VCQxPWpCoo5GTeZlSRo0u5CTW15iOKYbPiyAAQQV+X3IC0P8U
j4xsPFTodtyoyMKYsIt6lam9Didt53vetytcyog91kbDSmquuuDIZbVSOMghm0L2ElztOX/G9fU5
dx1VoudwdFB2rNdFaOOCgaeo6EKMV+L+JmxF0aw/ultk3Z2kfu6iGQIQPWn1fhg9SEcK6WNf1Qtp
lItR8c6hGzzHw4xot7g+9QMFE761zPt6iHF/ddoiuJ9p2OhD4tRnvL/2RL5sYDI/Jl6bHW8pANNb
yklrTdv6t+36AYo324rRcSKkW8GTA48LQbXuVGSXL+IR+ap+e1rPz8r20GTz7PKp8ZPD8i9kgRFV
5OiWxt3LNhENd1bjaLoXxCZNjkkB857TBh/p28flk380J/MXuAN/9sqe2Hv5hLlgKa3i4vB8GHb6
BtBAAWnXNsQdPQOUABunSnWgqNc4+vdmTT1ibo8J9iMLDum4u5HlLs71mlSBOUY6zYD9jymzEtCt
yOz40QROHiyz4xyjoftU9zXcUUQTr81m7VsSmVvMsbhtKfTu+iPC3JoluLoYV/TEqfu6kJtMIxzQ
g4zre9332L/3sJGjFlRG0/8N3A12KrdMKZRsvscO2U8MS23KyoOM9nvBG8QcpQXZkpAxxE2Zc+9f
ob/Yw2ZtX8wVfvdQ258E/y/BvjwNDdg23FxaYtysSoE/ijm8tLPYEghjOPn8rKwuF0Qsc7655Wyv
SbzDMWu/FgryuZ3967SZsFciA5OC28fLLEIig5vMSAM6qgji8vwqmPCFUNEG29RyXrtZEoHahVPm
/TlqnX4+QDskGX5non/3OT+VqVh1F7G/pW0ExTpV61oM8QBbllEMz54ma4CT2Y1MndLiUxpCTd5N
tsbNbEa0x6JIhBUO9P61HcRSY9DYbRC1ietXCyF8ethZyh9fKPiwkC708CQO5DoTXu1MUFO71FhP
P7nyMBkdlRq28yH+UqH3wlobRMrIsg5qEeNnNTRj+oeVC6ubqTeZMEODmM3yQXrQy+LOhaufg5Dq
oIS12I8MogSI87Gs/zas+ZtaDM7rYwoy1MtzmBltkiy0xBoyvX9CVRdzB6W+5ynREG2pjE6Y99PW
0L/b0rSndQT9RqsEee7CVNr2MS11lgO83f2p66VJC+3uScShFlUegn8rHLgwHAuVpRioescfN1xd
QASNoLuACr9tcnjlJlEvQHzASQMJz6cLFeJF8B74NS+y51RuetCJD1g3E3M9DgCOzZRFdlfp97bd
FWtcE0Gt6BfRCd/dF1WlvMegHACYPX+slDEpIvdS7k3taec+TKhssi9YKi4OYOgI7dBvGUkMCnVb
B13KzeIXTcpl/E0bQR3dEnbhJDm++t2oHeZ+q2mE4+mURpOhaPxTxWWUzmtcbi6OhdU2l7qbwhMT
ZzBLf42stlBXTput26XLm+OdhVxBcLeFwd6+mxYHIt7vRTZe48g7vKV2Rz8IcDH9ria2w6fYjZlk
J/gwqIWS0bBE9NGVQqXJPnhGjvhta7IG52EkMzx60p21z8lAHvCLgCA/J9ZNitDb/fcmiCHu3y7l
s/+wSJq3vOGDnvPHTEwRZ6VHE0195y3+p9e2yeuSMnXbvrGYnXLsiliI0JABsziCB/BAMdMq0Eaq
IcGgp9qFGhRWkBMtHcQl9yZhTxe3bTXu2C0GGH23s7grwC7HX+oPsWzz3nYFhGDQnH/INqc1K7va
xGeoANtUZ4B/HIc9smrf2uZXBFV2Etqs1EOc+ho3jale2mIWfJrO+CS2jFulxpaTjCdf6CJX6AgN
7Xez3qRodFIZgSYrAQIpYkc58Ys4bxctLgGF0BLFW8gyZi45WdOvupPUdEeSy7JL5nfDf08p0rgh
wJzwwK9pdfEVts8Z079OxYiESW4ezcTIgIooYrM9UsuNJl2QgyfnhsnTESwLaRlAthmvQp3c0utZ
Ew/9GSe/Gh7Bt7qYwbk9hVT2QvxPJeonrQrJ11oXzrIU56qR8jsG1eIxV2HXMS7xiw3myGRvsP7p
pvo9yAX9HSdtt/RpL1nGXwVGq6/OPKKAdkL/66cP5KRP9zIGMDwkFANcm+HQFmAXF/o9+YqQkPn1
Quh+PUSP4n3ZbiZ7wy82e+WNDyVDrCLZoXn5/jQ8zcLW5wMVuP5Ns99SP7syEDDAPIxe7k7XCnYx
Krdx5j+zmocQCkDePTU+XEkxpl4RYA2ondAnLvRC6P1TcCaRAtArk/mTwyNCHC8OC55hm4wzIb/5
1YSHm6qCKA7JspaJrWppZ7L+Ioz9dyOILDpJIMlo8O5qGEGZKnLiJEcqCOp3J4ueEWdFdki/qAyy
mJFgfHqtyThHekVL6G2XGKr2ILzDwQ/hQl7DIUg9s4QaRhGAILp4FpOVy8ySI/U9ZlQ8v0WZNQYE
R41WSg+PRKQRh6DkaXGF8A7eb3cb5dxXjYGTa5bZEMBsCJnwBy0D3dCiMzEbVJ7FYMJdha+3H7Wj
N/6EnUGXN83rw8tTzRSw0vPWmwXp68SbfdcAG3RXgRmTMN3ikXKBbANQQjxvqma2SKU9SxF6n4xi
6tshk9yVJwRRIx4yaO7PF+rN4FlfogOFlEDwKGVOb/htaaYMHOUXYmNlLCH0VGlx0J+u+rGCyLee
iHiPHkESw24bI2v5iUA4vNmfjJFIykbM2ZHIRX79s/zc2C+gJNSN82UziF01fWdWuzdTYmmM0hc3
BbFhN+z+aE1wosdSdMOd2ljcxWm3AUmIy0CTJlJEMSjhL/EG33aeCzdK1TeQYoSJmLRdZwJoN3/+
Wec/vH08cu0v1wRck3NzPNx2SPWO2FBvlxjCseHMm+nXkylnGekEIzEtH0XJQZDp8NpIY2wm9MLO
INp6SFm0tjUMgsuU5Rdt8QgaeorTGTdXbiAKRYBhjHjqzfUeoA0nhLVwokjVE3n34aYmYNVFnsEa
NhGL64eGzBVsIGmXQQiTkY6OxasW1Pro7qh1ad+FtjdEZeV98J1j/uvoj1DH8u5XiqlW+iREWCBS
ZpEfZg1oS+JeWK5VPE8O0Q7tx9dmTUgz/LwFN2RwpVRx1nv+HOI/Z4o4LUA7JAYPXFyhtpzQVnQq
FG/28pH0iERP+kX5vUq0EjADeqlLTFJhH0Oq+JlXUesgWBgp80S18DF4UsZQDQCTii/m4HBlBAWV
ZBjGAJjhBqufGDnanoh8gvo6xvVYjj4Vd27Fuom+Csb4bplkJFyyxeUgDx8r5HoHe3Vm8tMTLsI2
MPI7wNYKVgnl7u894SITD3YrCrvC85AXPkUHCySDMVDKfxj9EtFheBnF+I2dLrD3bBSJR0ss6167
TT0Bb4UsXeCMMbLLwVOfspWA7i/ECKCVpL4b1/gbjOf+Q/FPj8OumNxwAGLYJ+mKelKe4WwGocOh
/mm+UrHv5p9frxpsJRS3meamHM0WJrGVqckMmk8dZ0RhLFLhpmpenfTt6rXTK1Jm5GDQYnAd8j5P
thtKh+OPReh8+rVvoreaYLHRd54oDeYc5y0AChp4I9MU6EiSa64JKIE5XoAeUZ9kYFnvB29k55oh
Z4wqqkgmxYi7Dix/Dqvi51tFu3SIvV9P595zdPqiaJvZHqXD90E6NihTS/iNWeMVBTSszll02W5G
usKc4IpAxZJStQ+ZtFR1/9Fd6704JaNSHwAnB1c60v/mBZoE0NzTZK1pXT3QWufuBuFNlqxoXuRR
36HqKiK+ygULaoxX5aU6j+vZ0U0TtHEZVALK2uHSw4OGFiq6shTJYBnZO64SiCV8dap7muSh2YaN
ITEy9cbZU5QEBgJj4pPk8TgnIG8BeGXe/bEmDS26NdOfIrByxKtX6j/2n/ioOvMBgsV35vsTx8ib
tjDobwwAWHPlZ7Ab5s2YnKreP75OU5aLSOc7BKeKf7mHQQ3fcdRSOtiXaBSEZpTLfFty/3p942vX
35mKvYp9pWTDAD4eXfeaIEbpF0dlh2wCRNK86dBlpo/Qj2Ppisn+2NptTdSM/8ts9JgnMEr3JTRx
YI2g1QjNHw91hZ9X48cYoECAcCi53DxtitE69ONJYo2uUwAQkI8oNbQaFWtnU4T1xa5btj7GZADy
aCbcvkJE6ui6iY6D4CKa4R+4TPUFSNaR8rGWu/mVoXxS3B9MNLxo2khwNaBhvPKhXcnFoUvyxsDa
0u11afbpzzX5lt4T84FYMLf1prt7x6+vDGPis4uDufdsoum+weBsqCa8LmWje60tN2CYCpJimbPg
eBmFVT+LLxOG5IynOBhZcLXneP7+eEidnZa4C6lSpP+qfMIVocisMGPmub/dcZ/S0phOdJfgwcKP
qVk5aQ++6AylB2bY9RqocTCt8Swd/UxbCMd7v4ufYxUBiAJFYKYhWP/QjW7mkSv8yoUeRQEY7aV9
jMou7aJ7ogaqcRAcj4NUorowc/KIr+bF47az37wXechpgpW9PdOyXUUIrWBuO36r30Q5Q7HSGW4f
nGZcc1LgDZ6hUnUjycSTPef6MEGtWxfZ6LeGVqFMx13QPJgVA1qL+nUO2V61rj7iFbv16jRy+lI7
xZLXcrNwmLwM+O0DnYs9t1MLQdICKNZ1JNHRXZPhqQj1Gpr9jgtq7l0FfJXa+q8jz7XLt7QosD4w
ybOIv0tJWbkly2NX4Gf0Wy9rcOPhMmpZtGSLOIOPkZ+U1pKdHORWFgWmf0BwgczEdr+SS31l/GqZ
kWGT40cyofVGJX1srg+GVx5A9S0VUetBdVY7qsb5c18CrZwRpIXQyXZiFrnEtRUWsN8qdDiT/kEa
iVNb3tV8U/FN4qowlBteo1ZNKvNk7zYPb/gozjRLZCBEzOwMcSAHe4rQ4so3qk7CYkTGJjmAjQow
XzGfa1YffXTzgjrv5c6DlDIkz/dk9MgIOkHD9DJxjSafXsYrWbYrlo6RQGk2DwJGPc/UZWhBfSm5
9xRGI0uO0Jtxyn49tqie6jXnOmWkuHAKnWvgzaPHU1u/grTKSfxLqsCWY8vnziqYFdaz/JoP2PrU
kH/H99xSSS+GvyHv2kY3tonZX9l3a6GWhifQ4ctqBqcsdoFFfB5pyFR4uvlyb22x107Naup/77Pm
jOF8fNhz89sR0dMvtnPybja1Cr5IQjhWD11rYMRsFtbkWFT4YeEz9PmwZ2kyCh3vblieuD8C73aM
QZEjj+tM+mXnVC+IRmuIDlnd8QA0aqJr6PjxXVBXtkMsycpfj7QZ9RduDrVSRiS16Oxc6WnlrAKJ
fp3HnqtIPrM33XprZF3iG657pROWnsFqg6OLufuypcJGy8GvHjy4Nm3yNiZYhHL7O6Pcww0hI/o9
Kf3YmvdSPcJxc0zIkA4ebSeWov7khsGRaVvi4hvC3xsTUXVlqOY8wwe6xfiJ5RBTA3bcrKLQrOdL
zkHBkIQmouukwQAYcR2ywvhnFdk0iNuQN0RRQKJCXbb14uoKiEkutookXIPyy4sMdKAfvFs1/nAY
1r90OS4HYVQeztGpsaE9El0lnnWQypjsCEcU46iwlpmdOrDjAyZ2DyGy1jdyHS4BmSL3HqbIClvF
15F48NXUwWIzIVlChFbj6QUrhScGspewEWTjI2RmvfYS8jHEmbqHhK3EPCoha0MA9L2MH8USmJLG
a0xxdjO3S+9ivfWXScinCCC4SvQ0cBxZF3xZiG+vzzjxQOIMd1xUhKSP4rCPdzvJDOFdMnH4Z/BR
jgFc9A6Fom3vBeUpQu3Tmf7/QVeG9N2yRHHVbOcsPRyN4Sdx8ThvCzwvINFOCt/LSb0qNya67Twh
POo+RXg/8DMhc9OfezLer75aBjPUXqoM0M4StCb8l4BPPXYMNiL1XBUS4BdDfKlEhdGWmP8yw96o
UTgkYeZwf+PLmp73QcdoVbiIybQBZvgJ4ywyir9aIDgSCq2pkpT553rT+CNJCDX+xL9yts6jxZEm
FEPG7HLjwnh9fhSJb/QcsqgkpXP14wYfqrbXdZ5qlUo27SlhzKZVZTd0mwEwq4/sROc7Ded+wVhu
axxgwvxRKkny56zDZGGC6EEk+dbMHCIRmuJKdPrgS7hSLvyuKAtb6sJZ6NX3BuCy5UGstfAcSBTW
CeYajb3BMIQNS/YOZsSPcZEtQAdUe3Mf3/ntZ6T2zZsOcgRNFvZ4pV6KbivtY9jZYzIwKIe9QM74
nhUvyv4gJa0iWHArUcsDe3kik8GUP+aLxQt7P2Vj9MqaFugmoi778SvjvO1t6hZMA59HBUfOty0K
ZGfzDSN/qE2q2ZkAqyKfWaufq1ZktPB3Bizjy9BVHQHgtT8Ta5yRD7Thfiwo7cWdKXrgrCpXy6Y9
FivULZcp5+pc7TM9r2kY4h1kM6PgK2QqFrQUo+F/gvzWxFXXRKy6x3Yeu1MA34fJRquZGPw5bU/O
h4qnH3toe+5SeyvizrJ4C/4o/F30BUNzK4lxTBjM5OYK4lXVicNIXGG9Tk6vtGg12rO33MZx3eQo
hmmF20Yj4ov73CUjppUT9G/L2703bs2E/m5ekeA320CwGVHTcOoJS+z37HtxvNYJkx7p3Bhx9iHF
BaI6KhMU9vPK3FVZp1SYjkBQHDSdDY1IJTv5UQ4N2regon8lFJb4MAcMJeu3NpAr79j1/M1lQ97E
BoZ54JJPQBp1hREouSixa4DIf0VeTqZk9RJtm9WFczxal+Bpo4zctdHEGo1z7IHcGL0a
`protect end_protected

