

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qm+ahCoXbtCT96FlU7osNjp8Kf3rDAFQ8vMBTpaKgTo3EvHN1CM/XiHNcIsmMQ17hbL+pWxo5SQe
TeNJ1GZN0w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KB+ek3mkpx3N+ihSLNljgKYzWfCbUQKXGho6dSjrHEWrzL9W93J5UQjcPdLkP/4r8XQ5AjiJVm8G
O0+WgdiO6dbDdWggVe0UZIQ5qp9jotaT15XQQVVkD2rcK5wquost1xsRm7MTsEsCbzkhqKPM6ASZ
mpW7GzuYQ2vDPmY/r9U=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5IFnCgXf/KjXBNbWCJPfF+u/Xe3PWCvLt3/lqQEWvv6nS2jJ8qz3O+bSiUUxyt/rlAZZm5DvQ41j
Vn2wE7il4mdux1L3DFueP8Ob6UEbh6yobetr8hrEOpbRcnmnH7rXtvR+yuK3psDEpqbW7d8GyDcy
T6jGK5xIsUceYrUwudt7lxYx4bLnzP6q2c6uLhkxaoLJTWJGh28se0dzlAMX/BnMMfjK0HDKD6kp
1VwH2Gj4iT7DvyBkDmISaH7LPSlLhe+ZmQMkilflhi03bS9w9ABaqs6v4fufe3/pEUeBrvl3gRH/
oCU4QtUwSf8qfFsWdX+C6Nn7mzOb0WSGIH22+A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BAf2bWZTeSaPIqnT3j5aNO9C6t5/rcfC+/QtvmxOirWtcQ57aHowXlt817D+9PTxe4qEx5CjzmUg
9oMYSESB8IK4XXnHzrwWEKN1a7YOhI72J3KxmNssnP6jdEMx0znih/oPMXJaAdPPRUXzSczvXVqf
S7AhrmorMi/7B7tc1xI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dVk9aS2pcwcb0BrWR4Sm4FSW8QQWqHH7xHbqUaQTDLyPydXvHmrmxiDqUJWu8AAmbDSnHtBnMo/b
vhz6TIedlqcgp9o49Jh0CEli94frA6kGx65vbdl7q0c/R9+UB+XDf9B8tq4xwdSd4Twx0zVa9WGD
lmNliqJyvFk+OMbS2OJJyBNqK6eZPVzKMFkUG0UJu6TERfYV2nuxVMsugR94X7JoKx+W2jEprOdB
UQVXsqhudTLpaKEQiNqzDCaBK0P3FekkJJMtZNaV6veO7wX6Us6tTDs6pxGysSo4e6tLocXysaO7
1blW1S7foypb+e5LTkDXsQjIPmjtBTMz3Y2yyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47328)
`protect data_block
3JLodXqFtE4FcDdenMKgObelwMa/SYz8fTmyRsodimGhbTeY2jZvbnaLbJqm5YW9MbfRwPIJLDaI
oipkBMYBhKa4nasuqZZ8jfZnWaSl43t9WNLwmP4HYjlWFU0y8c6sNhL3yV5eyH1reKMM+jFgRDgn
Uj0Od18VWNC/hDyVvbsnkfveuuh/sRbSJPaZ98eynSofS6LKhK9ySJElA0CeKh71T/VvkMFFJhk6
Qm25e/Q2c695YXIL40OHS7Ie0TfpB0QhlA+vgWNlElaAwq2tGYc+q0VdcKYHH7B+SR0bG+s0hSHC
7VXGEuid2zqRY8z1PVjZPxdYVIyy5dqaHJHX2nYaHeLNwihcXslJAO9muySp56DAEf/kCTrjoI56
Q9C3Do4mdb0SfEp4t4Mfmv4QuROxm+hht6l+MeMP+xnNOBKruZ/W6bcwAmhxusMl029mlFAYoT00
LGzkUGnx6r7/w/MKlRHGcem1uvYA3EIIo6KarFu2hMTbKGc7R0QXitNj4bDlxK3pBhNqPpQwCxRi
/yH3nOYSYGaZKHDlr+lBO3OSmHbZv2Y/tWpcPX/UufSWII3yQCS46md22J9nEL0zIkSjPUYB3oNk
PPluAxwBNrgbaiKoin8ljcMBxMmgIT3CnZSXZrcM/FTk1S8NdAa04TpugaM+gelImrf3hK0r9mfR
0sp+qxzNO+Ae0Hjvn+Hm3oNpha7XhEEp+Cy1QGgmdx/hEZFYSjKS+YywLl+pUL9FfcMT4yICe54S
tHpjajXc5fuxhioO2DhMxgTvVlMjKR+earyKdaCrUUpeuxCQJJpaeiBSfOiokFHgIDs5XC4rz/bq
Dy0xQqLayU2V94GDvJU7BI7JAUmqlx4o0XB5vmF8MGy1t5TkrbmntmmbBsnG02OwEHCvGFVpPNdp
KWvtb1iTSHwMNhqMWl/wTzn9cyvJdIMGK+6RzgYevw+GGkiRN63gVo8qd3hkEsYCSTpIBfve9V4w
sEVj5u3XtODH/2NR3avFCSJougVJdyH+dAMoEMpeU119xxus5n1lKz9FbaNc0xi9uAP6EURRXPKc
KNHP3idZ1eyxh38OIN7VOjimP0Yv9ERu1VqP8PEv2cx0c8puDsG/0duXUTx32+dkIbE9j76Dia7j
IZmNIbRGFn0F5mlW92+j2EYCbaoC3QDbO8o0LHMAtuQFjHSgdcq/ghfTo1MS4lbUTyn/qwLjMD8u
EdkYc2AB7AcMsmvdoJA8JFiVYuiNDxJJvykWqfkqiGJbuYmuQZGLtg9Khjbx8Iev3A9IfEbkjz1y
OA4/lRRPWV/ujOh27PPQtNqWv7ElCh1FLmJrhvk1Mfx+U6kQLyNwHrBMS4FFHyjc8b4rQWRIx9Mm
Umzba5D/h6avh/bss2DoW0qbulSSLViup/duc6cOempEss/tdO5xmefHJiEGJgDNW4FsoFZjfLPV
Yo8RHYgf7GA/f5fYunF57K2hXdfSmRUCF/Swpu+B9NDOiLxddemhOpW/k1oAj//Sr+PkEHIgw1Eu
Wb7Ae7In92gfwva87ZgVFODUlLwQYKsiQ4ukePgzGVoiGlSEcVeGabQRz2+OqRJNEkUfqkkK0yrb
8yUcCMHPGbIcEDVsmp5WbSLJc40KPqrR2yCUXf5f2h1y7ZRh66/P/gjfiyszAkEEZh6hHu7jL76D
tHwjCKh+UGyEafVPCo//OjLvjtgwaTCcvItsQZ0t2AtoTODMw6xnUVEIMszJaU9yzT6ZAf3oSsP5
Jl7uqjgBtbE9R7Gn1Dcc5nhYuvlfRuiRigi+OBWqMttoshE2kb/Mg2/BqxFdChZky4G0GqC9LbZk
SbNIPZ/qqSkApfISbLM3I/yJgxuVWO6GIOE6MjqMELMAhcKXRHZvwMc8rCSHhYU8GCxSiyqd0EXS
qlfHACgaml0gHkjJERE6zW6FRWVEalLBEuP3m+tGMsm+u5NNHhDG8syDu7LYDzgn+lOUL2NJx6tY
gpt/Obud5JHLnFrYInAWGY1GT/4xayNPkHcJuVlecyz+1VsieqJVBP1c0kWinMnX2g26uo31JPP7
tzI7zps/S0H/vmmUFFG/R0EcyQOO1GGCo6QLLfbHU6ATH27c4aLB/5QnKX/gSGHE6WsTfqb/eoKx
QcAEny329+H+wrnCPbd88QQTl+In0rvQ2Ob+Gtb0ckzmxhAVUELjfTkc+IT5Yk5XTEDDkLfg70jy
nOV4tRckhEO3H9t6QoKOKjv52U+p6FffepqYVHdgv2sLYLcBFxOaIFDBjD0fK7KdTITLeqsrAgND
K/xOVtzk8dLxlCiE+wB/BD2LcZuI0TS1EIa7QBxPwWetlJuyCXdPej6k4BDIRAiFyptIBGiVMBZ7
IN05wZRjOaz2QF1IcJhpoPptPgKsXbnHp9IRTS2FpgchAvllIvL8wu/DCfVPA21nmALvdZxmw2gm
6vsop1PiqYB+SsbiqyUqsiz+hvoY8e8C57ZUFK9wb+Sr1tYmXUucAjQmvybs/P/sqN4MGtKKSQxX
1aLXMkCXwUNQeNqyLqYbqGPCCl1Cyt5WszqOpHKYDW+DhcGMV0M/3jd4V3PzyVAM5wEUcOZ9KXjM
6QB4q9v5BI/tJbXRCVtuUu14SC7pOFqJYvLUdIHyLFMmr+qZJ763QPei4vtbWjqMjX+oQl1CyhEX
Hbra4Q1SIDnFPL1yJ0xSbWeR+CWNtlIBzhqKdl7ioEHWV7FHpbwb/9xyXZTJvU6qSdd4WAwfifn2
GJYeY47P6XQGIRzekyMaANmbXefqgk15dgUklsYax7Bu1+HOP7lbk7WBq/G9/KadKNVsJoMO4Wxp
qmSHqScfI1iy8KtwslbQZ6S19IjoxJbEJ2/9SQnbX3t9iATDgxUqMJEaqo3v2hQzhAs3gbfqSpSi
qHKrb+OfTepnztlySwajj0joMgTIjnC0C3v77+tF1rXpsc/atmctf/1qrknTWmNhv0aqJ62A2djk
eSL2ELe+JVSIB43E5k/jeAVziszv5t7hiT9zxENgPc9O822EctVVWHk0xKGXnv/GT5ATDmxseFOq
0at9ExHUS4pjxr/IFbQ97HcoPWzK5jM1FBFgkMp+yGUhkY+u+mah224gHP+SQFwOBdu0beBZTTCh
D9kxAgFcEP02iASvuyuV03bFdMG+u1pg0xEAqihpuErxCzYSVa8SSXhNPzGoETtQDpjKdkFFuRCx
XrkLuoYFT7CAkqRWMSSQ4kniAHIfLUCFMxL8EXa05wcFNDc5eSyDR+8mXcCWUAZ1rSz4t9aw+iYJ
MogJHwzLvDaQgMMONIhj7u+DNliLnk/5bF36pztyuPDX/6Vd03TLCN6KhNMAJReKc/P1dRe9nZss
b5aVMkgRhOG4rCyT9jbyLxSGRBrXoTTZmGdjNs2veBpD+O7oT/KITZMEvsi9/z1TwsOhqAs6iq6u
tBGI00PJ8XHBXc0BerOwQEJlBZkro0VBYpjvnNnt89OrhJKG+eD3P4uBPdGdODwih011exgoQvSx
VwaU4mPmpveIF/l4UOxFrUzWulUh5Oz+t1IJSL7aNOROSX79ATrwa5vSJFu7MU0STclOnu1nz2yv
2Jn8pm/KtjCRZSGSRwhOvXpkDXz9d8ovDUTDZBVQEm1VL26sNUbw9m8nqYT2oD1uW4c3DFJJyW7V
rmRgHL4jrSjWejrvFnbTM8r568fR1F+0BNfYpYNnHeH/46mIQjkegK87hDy6kXAJdGXHTi1qVm86
6H/n4VOgyW9d3gzEeX+ZIsm+qJjA3GUDK4ARUs0AswMJRuwjbAvXjB2VQWL+5fQuAys8tBGPGbaV
zsdkI1NhVMwQdKBMdrFXucoA6HaSXCQe66iGIjV9K+aXhjTnm6PnVu291LDpZN+aoUue0jreW1Td
4MhvoTqSwGVtQm2o/46wM0M/Bg8L1WFmDPBWzyCDt+mATrurnuL0p8SIsooLQMpTkAyUkQE5DsDF
q5OA1ImCy/iia2Jjg6gMQMbvhmI14cae7/Hjwnn9lizseaXrAD3Q5YlRw/8rRtgfzeliP81603yz
MmwAFma1/25xKFgrtoxLEVFa0iTnwIBCfhxJTU9OxiFCP9I6In8JLKlrF5Oy/izNEEZsPiUXspQB
RBf3O11982YM28LxFr8GrPD9JxJdy2cgskO2W8N9UmVkUS+lzBDDoAjS2nDJFjLFLGolOyu3nLqx
k4gDctamdQpvAxZIb4Fn+7V9ijrQR1DAV4eyGCdYxF+l2t1/2yQtqDmKx7LSygXuadg7D0hHQbt7
zKrb7RCHR65uoBXN6Byu0o7xU21dIK6SxDd4aDRsRY1uVarKkE5PUNpGhXQYV/LDyiQIL+U9M5E8
twPEg/QR146cnWPzCuLAZpiSQx/QiW56mXLCwXraUxZZRyeL/BOPk3plnuGQNBCaBcl9pQTqZZKN
wrjHeD5A8awEy5LQIHeZm2XFOvNauhfaTUvnQMGHwPBjGd6TWAvZnzDwOKB0xW8bCCWjb8RetEhg
vOTOAgBHWDnZywSKvMQxgFPs3gn69jN1Uwl0/g8RZcK9eBOAGnTTopG0ovn98Aj0VnamMGUcITTk
kBtazPpH7Gw6NA4GCHNTXr5Ti5Lfmsgqg8zPqWVSlMN4sno7eSGWfl3BJEQegytsTrL0VJ1Rp67/
4yAwctn1/b0kbYLRXQRIFka8U7czBkF6d5H0cgIEQTCKpdKRnLF/VvqJU9JNO0lrQ5oK+NmsFrJ4
0NiG2mLbiuhefvnBzxP7sqvAk5rHFEnKCcYp54mQnPBtSXCBpH7A+5cpBuQRaJ3Iy/zIondzvSZ5
PUHTekEKeMo8c+BqzvnBO068gMinJ5UQ4QAu2Ic3/QFEbb6KTWLa6gOZxShF08+hlgYG437Pey+b
shxHpgPhgNLCS+uxrKPrHoNucCGDQ2bjmp8/OYrAc4ZdpNr6K5cSJ/AVIyoiS3IN8+MlO7mswJL0
PlXuC3nyJ9ENv6HX386bio+79H/UI/nOsDB/CV710/4TBYCKTgDKEmjbX7gnoRPA4zBJEZbLmj/s
VL7U27oITYyB0bA9rboT0Jbc3SoakAemlzDc+qn/zhYIsISyLg2M25jdjS/CNbT/rOAkzF/+zxYn
LqpCh/boubr0yVGG1wQyep6fF49tsPJfiDzfIk4V3hbvX7L/jdtXCWOPVMowgbFtnbTQYsU/+Zy0
2oYD5RWzsTNTlT75M5X/q1DFWxI/o3Q++ThiCveW3BejIdDId446xz4ZrbCWqLH6jwIi3zIB5jF3
e5PyBwitVLGSfSbZbHG4m3N0IxHgj/Ai73yBYJX7bS20UQ2SBeUPibNxOgS/r2/7iPQ4UOuZT5x+
Z9yewxMQ3TzKuo78QSRXtr9VWd6NUdESF7e72i9LV5cs+EHQpf/XEgTYl+T4QJp2dkvVDvddDxuc
1LHIThlMJPc/WMdOdL1KvoDo2F3+/zkTLpxVSzQzLULbs4Ls3TKq6EpLTfZyOwnP2Mt+mctdIFt/
HZqy+DzFoSTuykVqNp/ts9A3F1BtWHNp68kF6PEV9Wn6KX61clmNfEsIUUWcaR1uXUBHgSpHK/9O
yvbqCXieFKGqkJUt4bcL+T7ML9FFPWJHahMsSVR7BxBqnFc4KhyaMf4y37FitOekOVgNB3P72LPu
FKcR9BSGrM8xTwCqqJp+8u3Kx9RcuHPMt4NGBdnGpBSUlO78Mdprleq5+BAt5+XyKqlCjOB/+Tb3
+IDDh9/wHxEXJvLhi6V7l/ruyVGFAe0PV3hbwCXzm2K7rICm4Bc3t7a7B7KhPTGDgs46hF7ersw2
W3EguxmAsJKzIwkCjShNoNUCxK6+rg7yfU3BMrTOoyXPkexcolBqfFJY/ecU8pxqxTonZprYElAA
Y5OzXkI0LuXd0kFChe/AS4sVIOgZhXlWTdvlmXuZAta1dfqCoUmRojR+2WBpznDj0wph2rlLgsP9
dQHEnXLz65AP8vriUr5DM0pHQ/xVor/nDIZzN/ZHLPeiWHodisbVwKPfYCmuawdO+Hyp78OSHT7D
bAVvRm/V+mEtJATCvnIEUnIL6lk6S7Vl3oTrnDpE6yRper8ldEd04ZX9uJf2/wT2Fd0nDGFLXsZi
VK2mawys7d1YgkIouH/zHIKNFY/z20VeJZ+auTRpf4YZx+0B8ZaonKgoWmtnPr+fY4IvhJa7CTv5
CIbIlZgkHJ5yuNceKpLe6y8qZ6o2MRTXyVWzPQ0mwu8rP2A+L3nebEaqCN42Oj5ZVDBa6G1taw3U
tlaymBfvmqRfUYzW1QLYyXq7ZXMFTN6n7JbcJaqGYnycNUS0Q6i4f5FeBqYX0a67lwQMz2PGCXHx
5vgzz0mw3m4BSeEbjFCtkdWP2m5EIicNNOjm6WFhlle5yu0qA+yLCD57aPMj9oonEozoBSiKow7N
QrU2IjQwszDDqwXQgGQBZzeY+GzZZOc1B++ixE67xZMGmEZzUFlB215sALjWvW6T7iGvolC1DF/F
a6IDkd3Ef1UYmb88cA5b6nZgQx3LPoptYd5WByw2gJhPOSKljOMZekBTAVm25JLZ5FUZMk3IUY5B
lrBvmTq+uMcQen0VM1Pavbx0nS61LeHoXZ5d2KmtwEHu/us5doqnWEJ4fHwG3neFReIvXoMdHrMP
5+YfrIOEcsNAjdtAY/VpV6RwMbbCkhT06HSYMhk0hPnl1nS4L+2lSQ/fCHB6IPPjQi+8tfi72Pyl
djB2XFjX8/foYjGsO5FOXFUIzbdMVdvua8mdbwNV6roM5NZ3G51rP0+Fwq7/5AhSlzR7kNd76kKI
GozPaUyByQkfieBgjrFlVL4tRdeQt5eBPiv9VE2PWJPB/y0UiQzJiFBzzPyciA6hXD6l10mcnWed
2v5IogZ+S4gWkOtkwxmCytthqN6wIm8CVxw0JzV/ADUSnJXRsuGqUSdyqMJTcl6eDHF/vIyEF+Iw
KRllNlDar4nKqpNPsyRs6CadE5Q+ukJlnIXzhpoJ7MTolBChtei6j8QqonskjF7WDLhDxA8Ks/yM
yMn6iCyVvzvu4a488m6IpE8u5tD8peDfQYCi6shMlIS4lapbp8Hu9zh5ScSAJaeDsV0b13rR9iMe
fegdQlPG1StoU+I1Y/ZVH8UeZIzhc+PQV/jJt65rYK8T5tbV96Q+ks3da7rb4aX47a5l+hyjHKYw
sWNsSMgEXZhIY8O0/Gss7UsR+mCYgM8Yx04UL/rEX/NHmTT6b0gcNeqh7YbjcG+PUCSG3b/tsr/e
PgI+kyrsKdo8ceqcbt6U/ttsxsT/PWNtd5XL+TC1VLUpiMymoJ44dbrPLFHW4PK4Lba94BeO4eBQ
42JsTFQcMYk8KueRotr8Um1rwUKnSOrL7WzBT83QDeJh6QZFGlSZbNXZci5vb7KDKceoziDJiusM
36J+SZ6NF/+s4BgnmHxGUt0Cx044G8l+cb/ynca+omVX8X/pR/TUgXOG/liMj1Pf5MYOBdsjQbYK
QB/0bWtVAiFCokE12KBURZNkL5W2pWMlF1geoRg6cTrWISE69Jf1h/81L+kPPiTb0PZkW6cPc7Jq
jSSoXqE6tSX2ViUghTzhDPPy8qXIw4drsgWxB1IAieuCNsBPzJM/boMcZoLx/lX3864gD6RPLyS3
ZT6wLAyvxk1Z1U1KJj1eNpuNDKJgAJYrQiNb8B87fmiEgStgHjEGBFBgkJmelZIvTfAqhJpnUXvM
tfxcM0z0MSnksjmfLhykbsZK7Z6tDpC2fNUUBQ0Ojt8NE4vQpAh3SM3pXBSzC3AGGuxew4VzxVbM
lJgl7mJCYOrDnqvvuOvMMqG90/euHsl6IjMz4u845TZvz0YJWfrwVQhdMhY+huenCq9x36mlthwa
J0MTwOG/3ZY9OyImtxYHlkLGv3P6sLCSE9UKAaQMMpoWGl/t48loZ0e9az5Rp7FEp/6fvC9S0bzw
kiicHA18DsXYpxR0Ssfe2PzTD1gWnGv+7T9YQ6m+gv1q4Y0GOLn12pLH+6oxuJym3XAcfudVmSVq
bCI5p1FVocL/m7IAkpaPU9B8UR9qThFy4jr8c/lhSfCXtJSmzcVarGCKynHR8qZF8YIQ5Wy4vrPG
JYK1VU9G0cPT6jtQbRflq3OmrhrEtTd1wl0r6jhHDHtNLpKit+YEGinJ3J+3+dIihlIcz+fSfe6J
9HjYcVxSIrxXJ5xMbws7I/soWsh59x0LB1kV1gbeyE4+NTg+0h3lyL38k148OlnZXtxx33DO3FJI
zZGT3LIcRwmhXTA6kTAZK+crh6IfjavCPVCIGOauPQwshyhTjtBKz4zhYUY5nJjYeaFg/mmeHjZi
tn3iPiOX2+L7UdFvkvSRFR4gsuEgFiJ6kZX6F/6OOxFrbpXS/nGKhezPtwju2BH7zxyY9IrFk5Qj
NYNSc2K/pRsp7BejSj2OHC5ux1VGNk2rO+dcpHG0QC5GWWXR0DouwhYxjSlI9NvWB6EhBMDz5JrU
zo23zK8YZ837okyHUOZ5v3BHILDBelBYfmkyQ1JB/wA2iwmFM/AV3ZZ0EhqtpjsnkkAm2xHvG6VJ
RqY4RmpL0124ijDWxha4yk7ZeQXgLAaNk3b1+zhfxHNPzhnpuc4ScSitr8rRKpPhfvcQFFxLay9O
6Wap8LnNrDTQaQwlhy8wqz6KACp4sJZw5yNfTn7EV1WqkhbCDsnl+uEPiysjyywSgXMRLraceF0O
1QoRrXMbtuZXKRS2p9EwCn3/fYB9ahD9DQ1KhsrH6i7xomTCVbeTNuBwwO3IMySGK5jWOp2HpSzU
GZ2MuM4yYBysH1HjSfiyQeEAxJh5Ha55kLxN8c2SfkDFLfEAowc2eW8w5JxHHaiaOLwqjk8ayTFV
RaecebuZRXrzCubXY9E0R7F24mSnm0Do92ec1UZ9nBtcqGddyFAEdqjXM7nr6dW/Xs2Iky6Rug6X
IaaNKXodMyTi8IW54OX3UYTJ2GaP2B6UjfzdpBj1Vllt5MhmekIwl9hrtpAGCeCp9D0gMnKvidsE
75vXH2LrDWR2D1MHBRV/UUKGCDEqkI3+4bi2NW2+vigbBrITVJdoQECgkAx6UHjaky2rbfInaFwb
BFA1bkfHu3Q+bo1KtRlEJIhV7gVp//8UczE6KF9kWISwAMi5pwGTAtE4VJxo9HiLNFIxWS7UAxwJ
tD2oLrzkz1t3suSDCqbLrTBQnKLzJ7V6SjuhgifkY2lLBMY3gmTNs3ZjfXaM/btrQoQIoOZp1sV6
YL6ZTJA1LBv3K1ptNIFPCwG5KMERF3zv0lmaa3KrYUS146VLWlrY7AtUAFf2F6lBgSZMQ4yLX97O
sRjqZozgg4JL2ML0v+JdMze4gxY21enhM9noTDEAvx6kAAE3f4A73K4IXdEenhcnzjXdVsxYlRta
FYkhMQHhlwcSbLlCaBS8bPpSpepZixquVF1mtrw38gWzvYFvjx1CQo62Pc+F/vBnTLI3DKfRTveR
U2i8v3Q49JBE3VBzBPtNADbqxrf++kOWfd93cIcb4IzmFZBkQeudeqcrZgG5C5Q9aD56zqr9xpqu
H3WR9hc0RHg48g7YaUcp/C15EKs+i2rM7GjJkyOG368SEf44qhCWxdUaDmOSV15KIiwNz1n/Vhg+
hIwLE8n5dMwCh6aCoUQD1fvsTUG2YH2DESHb1OfhCoJz6+tv5SC9OUWLd725WC2Wd3Qv3tt7E/gz
vhBY5Ybt4PLvbKlxZyeWKevqfe+9tjDmiUicJJ1lI5OtS7rXVqYScpCgsLAo2ogOc+wEdeKt+Hj2
NJJj28nGAApM+QXtCUbmUpUhk91705IktxgD9XbO5MWxr9VAIFx+A0bMtmrc2uKlZHGMewKUerdb
69ed5z5hQksWazUO7JwGcm0dZEpsHdFo1jCOr05iA3u45yyziYJ+X6WfMiaA+adNXk+Vcwv9aGz8
zBJTVJSgiU0eAEGiuq9hmNPPL2+uhe9j+C9IzGJ4RoOOsEvQLvwBMDDhWRHjqBA95pl3/yXs66AS
BE+sTgO8ZOzKzKhsb2rUt+b85X/m1Wt1lGSJwKEMUOBU1cbzEiMWrgHFYD33p+ZWpG/E6wN4CsGl
TzKF9bvkSf1Zt6SiYfuxJJ28PWRwHmMVQ1K87WsUf5VGgD1VhUaF7xSTWVfKdlVzGVYBy7B2iWVO
Ds/pbYXLOLWpK20AT4Xp1Z8XEHqsBQzzrM4ANvs8KI7ODH4+4hDis4bsioL0oROUVnkDk7ViPYRh
0rfqGmdhEwKUwthYKV0Yjm7puoF0iC14sShkbefO/ho6obsW1Vkf6hdA3PxrXbHnBCujrsnK0m8P
33gXeEd1t+QiDV/UigUfm5Hh18urc9XVuaswLFqOdbj5WMfEZNbr56G5ctiqFoAvhUh4bvRrtuGz
0+eL5nlNboGrEOu6MD5F2oNd+HztOA8VxTWzBdsbefn+dVUeAcZKL5KYThjRIM4ccbBTBt4Hj10E
5W115p+5gCZAbSYpQW6+ow8xQWD3HmEMpm7KgNYAJGU8mZxgICpi9Je/dO7F98i4Tue0BUE9TtcH
bjO8jjDlnxcwz7ZxE7qw3HTljtcC4JC/8cvUf/07/JmXg3ayFlbb8SSJVWJKZrEXPcNyw50/I6o5
M4bmrdAha1+ST8X9VzduyuDY3tXO/x0Xl86bHH/B1diZ5BZhFL2d5tzdpcia62Q3KTgRgeUtK+Aj
i/d6ejm+H4t/y8oCXHdPGs654LiEgapEy0r8PENxSSMOZB6jLgoQr6E4BHrkEu6cS75m9rcE2dwt
pykMcgCygw0y+ZEV9aB8b1uMsJ8VEcMOef8PTMYQ2L1YyTPlJeMXUo1ovImqEfKYYBABhkEgE4NR
LvLrcytw4f4+Q/La30MpfO8QeIaql87EVkiaBWMTP477lfO17ze06MSuv2LqNaNzUKAcRNJ4ojp+
I+WRLd62HY4W2s24pVfsi5I5q1Bracm1hWfgxkAN+D4lB6A8QrP3Ccp6uf9VVAzzJpzrO+GwRN0B
l913/HyQiZky7pa4Jeb5xNRf2LoNj+4ZagJ3q7xSg63d5Ds7/lGRdAiRacOHqf5GtTECXtI6WurC
cbXlN6taDcgosWgltSxO4LxAFHijU7PRZeNehwEnjM/bghHVj81Q1HImYN70VmrFV/2+YbhfHEf1
lxA019NBvDOd+BzSdU4vWf9nwuY8Y6IdhUn3uGCz15rbvbimn5nWdG3Mf0DiJCL6ZTxnLHQt+RMY
U5qFAT492kg727d4PNXkSzDLKbc8HV46OY2HExYgS/qrQQPBAoZkIFm+u/g0XsCBFmjhQIyPUQD4
WOYE1l3R3zi81xZkIJH6oulPZG2vp5LCQomEim6J1hN2U9Jnl5i4U3klocRCU/JpAO/fnUoKzOPZ
xy1wURlS4Jl0L8eEfBU/fwo3NgrHPQLLDsrKqGXbXl5w4JM44kK568xXJvZHVMb/LQTOq96zj+Ku
Vrs/ZGZf+1Xwkh0gXWf68UswgZxC11TcYbbim5feMPvLzhSD3NBEmYoBZmo9lvKattj6Re//xUtL
GVPK8ag4I4ZFol9XsZ99Ne6+abRI43CR0cY++LzF7lm7TNhA3jv6opV5T2q2YuCXMJ5iBgJM2oGR
Ui5AbVvvchALNSp5NmD0xlpibaV3or+G13Akn6NFzB4k1jJ1DuigVG1jqarSgV8yd5jaWa6gkKbR
PKMyB5n/tl6MI0gm3NWsNCGipcaLI3ltFpFUSHiTuy8gp/NqS5zodXd3uEJOknzpFon74FerYLTs
A90exf0C/jEtVNDfIl0wDQt3KW3F0CpHYzr+kZVtE7dzMfYPohf1dpdwgM/xLqojL3m/4c68m0CF
Mumz0prBolvOxiB8jXXcjTSP5N+xL8dkjWVz8UIi9KK6DDHapIgboigYzcj1/ezq1zGYyjYcBXjS
VdWtHqV28OMFqOdwfx6JrPDAKXCrTOuLRgtvEbaPl42cwd1ko/3vTzwhLpCfjFw4ffJydUXN2IP1
Lo0Vx2OB2+NCOynTjhMj0z7n/abwp0OLLApy03sVuP4oaRpibbPksgi8Oxl519f63aUYxcHaJwPd
i3zxRh5NGosaUi3dQ+fKNJ2hu51RV5szLx7w+rcl7KMBRyOPQBUEY9zkB/4rwrPDpyhW/PBbbVZu
YFN5vdal1XdfkmxenQ37NTruLwPfyMiK+BhXXKQccAZ8Guzg+kBJukXiSQeMUbTX53aV2KOxRhy2
yAM9ZlZbeaf4dnlgGaHcnLkMUtvODc6M2mPpkjGdzSW8gsIRuqjPALogTPwxAT/bUtXCplu70EdO
LfzJp+G7OMujNDmR5Gj5l/z+CCbv0vRTk6WU1rIK9MUW3uCLZdp8VIDoNVNp2EJw8xgPEqqSv24r
Gkj4nt16G0cHTYu4l4A6HupPGVNWu3dkCJ1XOoW3pwKEvZwOq/td+tuD9wwe5kCI410QBj3gNNce
UtGDj2bAATL0resovd6a5QKZg0SB1ZgnB6XLbnz02VL+LxHKr8IrhRHbfJmcgx2X1nejebD/N+pf
ljGAOOfjToiM1fy1C1bzsGNwd5rw17GhLxZDaD4VkJs0RUpfOLGde7bXmAyNnXqQ18fJ3dUIRZrW
MqlQLGfP770nxcRhyrVoT50ZYE//bMUke9pxH6CNWjvmWrk2DQR5FJ35b1W5gwYRWO1YQxV1N9WI
JUJczLkZMgDxOI+yfCf8Mv5miI/4b8anlWLyxbtS/NnUolUEPWCG+J5I1yNCQB8EnaCoz8sXpC6Y
N9qfhR1O7gaMHn4HU4axXH5OBN7s03zLkFuGxetDMwjj2CXP1yVcfrWLUNdD5srfZ+V0xhN3NuHZ
ohCXYziVTM4BwdD631lZXtYsFwc/ROR04nQRVcDuBLZ+99VTQUooaGxgOxDZftik2/BsrjjhadKE
RS45x2M5kemUPb1Lej8rSVklpaTKEFaJ9Di6oDLBWP8zg0BGuU90cvB0130RfrZAW+p1YZyvPg2b
Vh+2UcE9cCIJ8V8ID3uiAwg9YIVvHVBmQ4GSwVzHEK9zMtRDD6VfTTQuZhFtoE3JNNlXjsGWll2K
a4zzTSmuKq3bRd8ctwRMvwf3lQGTmmiN0cIU4eSfpRst/Ro/2sBvgiQ2MFybTngDBuiA6cn7UsiV
ip8QLwFNRSCdp29bznNT/abyfNyCZs2pMxgS0tICYhj99U/OeWibXxyFGVhRabVb2VtVUQoe7vzU
ySjBcwQkLZOJKeAbqbLDHrXjTwpOQ8LoY+Pj2PkV32YfAMeA+A4OVBHnZIZFYjmT+52tKqhKVykM
d/wfJ18PvieanqEQ+KL3GwK1lM1O9L3NmfnmIFnwpiBmG5EcsMUoUfMc5dQlV5FU2jKzit0Fh2+3
xo3pDWRpeNXz5CJlZR2hsoyZg2Vm2CskrpzN7PK9XLBbWhi+Yck0Ja6GppD4KOfzMmt5I0rILmhY
6YHVjLKZ2dA5ofsxdKy9lTfCXtCcvDph2OJPPG8giYP9a0wpBeS9n8IumNrLWGHV0B7S8wY3t/cU
0C5ufKN4lB2aV3TRD+KzcjSBdX9vmYhtU2MMEDiLzpVF/i9EtzcqDjR9qfeoJOT1HpEdpzvcCZEz
udQBQrAXawN0fr90ujI4T0UDh9fzm3nio21q96h0kU9nakIPMTEOQc1hfQcZuyVKaHaodyuDAi3B
/6d6w70tFb3nABqxC8+WWGcKB5pN6SKfES7f7thZn/Nqtm8M8i6iVCdZ5XqP3NPsJNQCcjJgFJRS
ZZafu+DmQnUMSBuxuk59wZWucASu6H1Og/1k5I/JgnEcwBhYhV4iUrLzAxAZRII2DbmcvO0iEWoM
RlP8gxY4jmMrl9w1E+x2t23mhphyYJn6eOG7gUKEub4W1NJ9hLGflpnWM/hMrjvkw+l6eYCO0j5I
H67aEYt+TE5UDZ2V4LQ/Uv9Mqri4a7E5vz1JFMufGMyeb9L58NC5gGWIIo1GRn/+/qR4r9exOF7o
u8EWN5mrI8GnHnnhQy179SxFiMZIQ+vyXfJNI6adRdJOoeaEDZzYkiLysSMDzLyoUJGJSIKjvsRO
x4Wn4NttjKhuZAhJJZvT89dDdYczfw+ImbdBYdQxnIEC7YSEXClTV8oSogSGYjM99Si+41J/Uafs
kIAspZ/3NhuoMypORW7+Olxb8uzeBti7rbVpquAdS9noGx9ufjtemfkaWBD+Cfm7X4aHPzF9rSUb
iJ/dMq8Uk24GchomGuvNl2KXQKb3Z1Rkvy6vfDvpMAPbtQmZnAN3Ue6Fypc0yqNR4fr/vzCaVzbU
/cX4swBXL5K0Dxoc7lpqKGzVit+bU+NOKJxEhl5FG6WpsvYWfk62i4ucVn4m3DSydrLViXWHKPEs
0Q8zwGIfcj+mIOSZFxZZBgVb1t0oweFxl20goYs6MHNMzM72X9GU5wVwB7EyK1oPJYysH1U1vQgz
rocJ3QU6TzdX7O5yTlTRuHWfwkmsjPRH3gADocKoof1CCcgv/ZevE389fNnkD3+M5uFp8iULQfiW
/yUS674pu+xULa1riSlHOMgFDK5GYq6qQxdH9ey5yHwK5IU0r9/e0xqFcgUSYduuRnSj79Af9wS1
GGbb0ifNsw9N4K9gdyTd1ChZidshI9M6a55FT5vfyxInkFS26wG09ddx+x0bSikNLJP0cAY80t0L
2vA2MB/G6FrPitap4rZhlUcBs69SWSJpBI5gzr/0vqI/i6gJtdYpiU7jWtnOO4hTBpDB+SGmCfT7
nXzjx3CTdAwStKgJiQ2Zk/RV7S8gddtSUN8acsZpwW6PXDipoRIgkB5EKACkLsQ4/83cQ/ojzV7o
mDFME8jK0LUNbZVVzYIMOxMat10llwbTMixuZrvBksVVtwmUYEsO+QgqtLT+TSpSfo21VugfugaC
oc7QukEW7YqYMhk6mrd/dsKnIFOEmXBieghR8Z9uelrtcHVfH2xqKebtoBizrJ9r9hbv1vn3pzfV
Je6ZSE8pW6WmXZFMxZLv7xnqIderl44uTAJq0PvWfPEqsMjNHajKQojqm/sqGFmK4v6yr4tMtFpM
e/yUPgEjBOo/7rO28AYcqAX094QwyGYj6okGkn94PZ/qhNhCpQHa4cGCJpdEGgfZVdVzMt7aOuWx
WuMeFbQc0GeEg/pUDanpt8Snt//HzVVK2hiLvP5HIx/uto1hUysbq7VsyyJNgXj40NN/7hOxP215
RJy2F7qQoOTdsvSPBT0/gRr/MB/beLoBILMqq/yeUFXJ3p3zuKFEJpx/lrK2ledGMzzifLzz1Hab
fHdenig/hvViBvzkFV1vZ96oeLHHC5FGiU91V3YlIm+00ELlnDFG/fJ1LZzliqjCDt0jp6LxWSzE
4Fk3QO5+n7NOWi14sh6TrKXHWln1s0DqYvoFDTSMs0YqYPv+xgq2TnNDNfdGs1LWeNRPO/qijZ1v
W5O9cGtIBF25f7nNXd1YvjqC4koU5XBadqR7ZeZUl1Q7ebkkCFKHqY/MIHyq846vQpnj0ZmV0Cx1
SrPGLCl4sDaMRD50rAWaDL57mpuT4b8eikDUEU0dSy0Uv0c73ftTvYq5u6k4S6KpE3WU3pnGiE0a
O7OhZ3P9T8yov1Se4pf+LnXkO4ko5stJ+dZAXImat/ZSneUvlLaHqjRB8h58DJOSGv8wisiGe55N
AoAyds37CWGCq5v1MB/Kd5kBU29IMVf6C710iNYY3ZVjAdVgPKxklwj49+DbdjexEg1JF/nQDzMc
ScDV4wOt4wk2EE8WCXlzioomr/88vPl+jt3pOhVU8TK1KBwGJ7qIyxjT8CNQ9SfYOfEI/T82mGAW
bAT7AQrjVGOyrCo3vDGUrF3cL9XFswBJ3fkhA8/KDlDc00nbnryhGM812Yf/5b2lcDlXVyvsSAdQ
SkyKoMTZ3HxCtClkyYiCcQ67nCk3J6TBqf1KftHzkXH8k0k957DvXylL+mqEe9dA37eU8kf+nmoP
yXGkMhfbJaEMfbXyUFGzyRlDFvJjlCS2Rbw8qlREuOs7SeW7A0K7MlnUr3LsvlCfmz0bzLSxFyZC
YBGvqWGWCEuEdUMeKqilJHqIVgVSPcJulJDatRt+2tdWa7slKdS+GYCgKmdD1BmmaLyGapBbSjW9
7Q3gxDJZPuC4+2/AIzLdmS7bYC3TKq4G1Q59h3qiISsvfCqLiMoKK6zGngKRP2Tte0hrRfCVmKDO
KBnDGIXiNL3Pmlw949gkQuSXWrvycMMrchpP0PpKHL0dvpbBT36qqLyjPc+7JmEzMi7CytqrAV9X
bRDrvbrmSb510vhwhANIXldmNshzzPwXlq9/5mG+kVBQFfho798bio3ecrEWfEloOTT7nKk89O2c
hMlQHN7koXAzBzHDqZBJ5HRVKKJRcE08Pe7hT3A1z1GNs3WA5pAUh1CVBn0BTUdck7y+c3I4LuPz
YtjnqgSLEmzWCqMGS+7qagqDnnrQG/0CIuLAFjghukbTLht+VZqOVdaGVsBlyXi9K6Ole7Gg3wCH
Ba1Bdw14WArxhJSIT3JpB3Gz4ihbrdkTgBocMYlgfFGkFejvlJ4sevB+LFiACn2UXrFHYilPU/bi
2JfgttSgDx1z5iIcL46tVJaOGhEdhHTOwL8H0Sh16MMXDjYp5oue9/C2d7c0XzsxzMMT/L7rxL6O
GfPsWuEUggeT4eQa1JOUL5CDMob3IdxyYWizI1MRZgtQ7eMyVB9PYAHDiqMlnquq/FaVxsVUmZL3
xLgOQY7iMttBEAOpiYdjgGhNW+tkuc+4o+l8fVqvPZ4mKgG6Z46DscwW3bv2D8t4iUcIkfQrOeq2
sCc4euFERrxLALfxJpGi3Yy8ey0o/oFR3WgJSNenTcKTfvSZPXIbApBb0kkqjCOoFOZdTi5UZ+94
C2PWk0Eu9jVfBrD4ShCUiENdZ6DjNCENfrwarzNuNujelzK4BR2kfgAiahe110QlBRrEv/Gvy9eK
XJsKyaFWus1M6VXal74qvc8PX/f/02+Q5mVyU+9G2f9jJpZjT1fJf75StBVUdKLi8xPF24P01NWv
vMr84oYjCLzkCDMdlNVg3qtz0SoVr/93vt95p1OJtZohSROXcmIEQzqdEbHM8Bek7mefi9ZgslvM
tOe5wnLy8RYWYm0aa1aSdTVYz9SHfQreeErRqf/syvt/OhqKQ2wtTNKbydtD38xau6RJG6I81Cmd
4hotaQVSRlKwUyNDfgm5Iy60WOcfccIgM16ZO14Ic5IT+Fsn+WyEjj62UxfLkLqkynjSQdi/UFPp
Rmrf14NG2pCA0OGJF7JxYchpJLmG7/MQvEZcWCoN4UxF8CxIWVz+Fp+LUO+8oyee98nDKAb+1HUt
39ssJ6N9wPfGEnNsMbv40gWj3ushKxMbCtiXPqwi6waNtJ6cwh/nShevlmjCn4nWlJjJgNOS//xa
vBvKbOzlcibHRNHg6f2H8nOEVHde8YZNSicbScfmvjGErSk1+RMgO67q/kfa6Y+yIjWG89/did6j
cuUedhvxySSjxJzOIDitgSCdMBR8siFxO8IDIxyB0hcGFzpMF4kdxOiWdAVhf8CD7/XqFKz2yHZb
tgdnV1HZeiCupBfVFQTCqojNYt8RHHmtPqMLGoiPRj+IaD2bmnc0mGX7xvB8TUuch0wG4SDjatOy
7HAhI0xgJKE0zdMPXZ8UroL1WtXu1XpZRjmoiBeLCm4ASu3YUbr5kAf26oH2SBLiy8sshvRLF/ni
xu+MiktzRVJ3LGqrccAgIbkkOEQrBX7Vpljhnefw39wZ5oX1w2Ev8BtuTQoGmtFUmVOuDebG2r0j
qwG2F6sHm4KQOXnk7er/t8MHRJ7maKZLVCdq3pWeOW08YQintkRjOeXsfZNFMABqyYS+e2mtqQjJ
2FDeugjr/1EZaYnalludbKA5rJz5T3oSWPEB/BeP3GQmboz9gSFRiDGxqIx+Hdjosh/rV03QH0kZ
fcMZKx52jP6yvISsZctXBTLr2vtlx3C51yxZDmFceBmGkATy9Z1qZdh4A3UXzZGmJYZRfYPbJ2HD
Md57neCIz+ICFrMFC3jC5OYJy/q1xZEESGdrwCzkdhrShuQhGawoCcW+q967pJw+tAP6Dezzn50j
Fh1PZhZmLUjNVynW7prSmfzTnmb74VKeWusNaopImjmd3QbsF2k3FB+DR7LFSuYXo9wGgC4/jBgd
mLKKRJPvFo1/GyHiU9gF63d4IJDPSSa/Z6mWmLMWZCGIYg2ON/ZwPlAy8O4CTfn5vum5NyAygNgo
SmL40aSneuifyge4iPmgBNVr8nzj6dJDOx9Dv2dCgfPvUQ7L0ARGQ8Ts3H2K1FarZvyxVnTBB5bN
nNzWGoQK0lLW2xvciSP8aspDa5UvPbq7LXDWyxJLBEllmNWw9sZAYRL4JtaooQEi3pxIXGqmkrCD
exoOqjXrNKwG38AAd6QwW3EisEPoR8dkGZjNNnMHPYUC5Ym7m71g8yZ2XmuKncpjML1kwSxTHAen
ubsO5PmSt+uABR9dDMX4ioImmhuHYq3E5ASdyF5qaeVnQ+WpJRndby+XkQTEANI9PZk1OCf/EATA
j8u85Z3Gra75bL4tx+PJLEhmwlKxwbz8yvlaYlfjxtpO14eqLs8GXTiBSStnGbUG88JB09jACKGG
iwRYg1K2jXPo3weoAFCGyQuCw2fovF6RzygUblDeBLmjqhGS/8tCjvoQSrdrTyCK5SDGj+FeEVOv
Kfd9j658qRJiySETcPZYgd7CgaSWqqwI+Jg9F7uHYEgNvfsviiTmzfuSNL3hnn0aDVvVp4TDGIj+
YHigJV0dXYw28ohMZaFoDVI8aVDy5nvvJR0Ff8JQqXetXaa1w7u8qBORu3d+nD3ZWEXmuiRzBo1+
YVKJFwm9ZN7799AuWzYS8iEnzYeFvwXbeb/7TmSUqUZ5hrWvIU6LWv+1qDBmbcRrdSsGgXOyxXF7
EjUFl4P1QsTQXZN+UGRca6mL4Pf+50ZyCmfSNNvB63hNtC7lNuMNMYhH4wFGcG+tFM4zatZDTkmN
JnXbtUlyYP5wQG2NUtRPLoDSrQmg3442Cp3CBZ2AK9V7x8/J0IJkoMrZ5HshuKzM9oKOdUqDPTFQ
ovf8R5c0fE9POKlye8Chsk07yIYAqMJuN5KImUo/ff8yqFN8W7bRryjEMxb2LLwtdjrDvhC56lTf
nQ2lYllCF9l9+1HSVFk22ozrIcOK+Kbpjnu9XmqASkh33kLEJ8DlU6EXBYCsYIU1WjPvO+AREcVy
Ry/zkRSP4Pp7iIwvyB2FIcaN1hznXZPwVw0LUaJoz+Qo4TpOmQo0z8Tzjd5sffJscB6B630+wVwr
fyjWaFOVk4YGlyplMLMwPW/vUWRN03AcVXMRDW3swFQ+jJeG+p16JT/JI+a27rWdHNPAkG6qXEi5
jUgo/kvIJoqaMDJ7Q36KCjDu9QyTnIFvJzDIzeUIbvozN3MkJ7syNASqVPisYlHDGM3QqUFOxluV
WpD2POSIA4Dg/0zXcRtca3Hu0MENUrpYShzLYjLZSZaW9GjPh5q5XiHJ6YciezZrAC9sZMumdGMj
DfvLBmoOl4yci2Rjqb2qTZttdK4R5r/fWII6+xruBh7LYzQOqTixaunda2nPvnI0P3lcfqt5qhAS
n6TLGg5Z10j7OH2fsYN3/we0Bf3qs5xJ9U2Iz7Paia657RJM1Cu59zLiTv7+WswKgGNoALpP2dyx
VdIj4p434ZrFkiJFH4LO1mvfFRLZdSXVwvEBYCcvWsQTF5oHlIQzcAAQGKVywB2W+xX2IUOSJ01W
oTtAL6YU70fkD1lIFOx2dVNQBLHUvpdAHqq7PRROw9jQm4IPGGk4rHeu3C3Ic2ZFCTR8yVCRM24f
wEH7vbfUg3nM5EQbMmws3T9hCgOifLgTDz+APG2Ov8eZgt363NiiEUSkUyU+z7NM1nlHPz75K4of
wxl1Gs2+gMUJ6AL7Q4hv6fbnupP9a3/vsJzlutrdx4IcCF5C752TpC8aeArWthmqyjlz2L06lIbX
jRGCRAPXYSCUfeNVx1pLfsQrxNVvMffFPSbVsD5QGSxEC8YuiEGB7lJEN92eUtnD0hZCxH+cYxkt
eXEyRpdIHjNPd61roWkYX9UtBRViMjCW2/ixbnl2x2IFBPPAct5qRm8u8eLbNwDBv4SRoD0THcI/
am3tHohA1VqMzsJikDR/lUxnSuUBh9OOK5jwVDWkKS6HzJh3QN+cbI/2SbUi2rykOdqKAoauYVRQ
k8OcJFClq/+wDj5jxcQLgYn7iHC1TVJVTdrqUqIoxHapSSHMp2ukniaWisTfqLEr5Y5Q0Akncvqo
0mNqjFpfXED3HFV8si+2lwftH7LxN9uvx3iNaEOh72c9Y93HkeTKkID59g5oYzOhS7aN8OqKa5zk
0eaeSSQ+CeLv1ucC0Pg9mxIqTAbf4LuSQtDZE8sOFcjQCeMM0BiLOBFhV0sUJN93jChDvF6gbDFt
4XoxhM4dWodji/M9//u1W+uYuQiPuv4rKOxMWGbaWiE8PPUqxKNcgwEEEr/q9obpApdoxuuJW6dA
+7gCwy52dvGaI5UsXedLyvrg17UB5qGnQ77IsnG1kA+93h5oYXe+dhQIIuE1W9mu+dmiPQGAz079
deM8a21emOTQ5who8IBO/jBYR5tRWADfMqrMx6Gb7HPEAfxAHyBwN6sLm4AU+23sw4ZhK50y8VLN
vhcJEPx4jLPrKMuTAXpDD4O+UujR6EAapgVwY3DZ6ZOuLKkvjCoxdxTeb47K4E+RD1eJhCVpnVAM
yUo+qKRL8C3rr/79dU6SBIdVVJg51o8/eCC0lZdJSeutK6BYjXonm9kvkR/gVUP12/VScvNeIY9t
a/vaaDVCWHsz5xaEA5SHOoGupSYhSGHyCxvkT/PwQI56Q4BNcsQvjvmp5d0Kp8P3NqbYpY0UhpFS
EDcq8OoM+ZOHuARNWM2fbZaPm0KCHfMj/qpoZkmG+OR53V4zLDfVmQDKn6Qt+rgGYL5X3YQHck7j
D085dx7x62dDzZwX8lejjlqe42ZMxjwptM2EA4tGZvJ+/+s4GHDUmeTwO21GSgsesfYkX+3rg8Oi
Au/c2eCLuz1Bx3a/qPyr6PqGnwjavNOPqxD7BrfCneEtE8Jq0dUgQfofUNkgDEhZUu+2/NZwb/Kb
EoNSPPqTLnB3LzkgzknvhCRjwPdmLjJaXLJ0ky041Qxx+nBTFWHJ0uDe5m7lYGpf1Ma1wqErjyKp
0bnyp21lZeaaNzRqyP6vRJsVEGPB5M8l5uUu3ltcebnEtj5Sm7XLdAOxrKGkQL3C7ytH/ymjznFE
cp9iv8UTcY4ZqMh4jfPIcmJ59fDRY0VWnTXsIe0maINyhNugg4B1D0aC+3nclv4evDkA4h176Kcr
Fj68SbULP4AwfSm/xZMl1jp0xGt1bqt/LVygQ5I96OwNsB6J7KMRau0kX6W/Io40AMsBoUikyFG3
D4x1HvSN/t0qjukY9DmZa/IOwKb02jPnYZfO8O/yXZedymCUILsV16L8BoExBOo8Ck9ZipnuKAz9
r5lNuaoruWzL1ls3aoSxR8iy0qcZg3beyfmMKwCU5+1oCC58J+662yWS8PAw0zD5mZZ1/I12A2fu
6OdfPVqezA5LsK4GGIUtevLWpMxtGF9W0y9/1mYuzcyXGZWS25zqY9IBq99pwxZsjUpMvJYXUCOv
3zMucMixehVClE8GSxkVE55rkkQqG7EN+rQ8By+B0uyutYxw67B94O4zTlLOR/h8Q+p+HEiAsB8I
ehf38DVnZE0sp+kuEza6e2SC/LZHb+MhCAxJpmfZ1gH3InR4tZHxR3j2fD49RwCuT2sN0mv71ovM
PXmXKoKKVHbuk8pDBgoyXB1r9ax0IAYWVa7L2C6YIWXo4WkFsR6TiJIiP6gfx3/L0TFDMMrLKYmq
9YN78hdimXRGe2Xri8ImjIItkpP04x/y3lQyyUg5eYfX5qkvW3Eoteyds+BMgTVcBW3Rer/LWl2f
td4OXor36kR3gma2EgfiF3bZUp0loRhUZFiumE4Xtjm26mPCUxerWVOVNJiDR9aR+AVz1tM37dKb
g+JD404/R0jTjaxewFGhtH8mUKbny4TNnZWF2t+XciEoAvmBdqOvShx8blUWIKM4iKJKBmz8YLPR
5DDK+G16P/Y7L8FQVRbpVOzXJRoQgfY/CDiRrSluFwxKclNox5jHbvusrAgSdRBEK6C2xf9J2ODF
ibE73j8nM/5LRORMpVjSK9Y9gF+4ai2YNGWCdZNYOlvqd0vec86hVtmsEYqJPhUqHPkaQ8UidBOn
wtlXkLMtrbknuXMDiDz/e4WkALoR+Tx7XkDAEHj6TWZS4eqXf1QnDErgqrP0vsm9W3ZDQriJ3QVQ
WIn845Kd0wmXmxtP9AzSMYUOb2x5+gIN0sXCM3vAKNE+FnGqExUHURCbzbUMWp3I+HVm5EwiRfBd
CsOC2QUae5k81PuifSXnaOlr6FMBpd7mgZfsr6YRlqmuhqtKwvMl2fb+cu0ZI1NLsWPxwWTSYZT4
cLejXunnANdmzh/vXM4FUxuhZKb3KKC0BE5vK1tOyUQ92tPEAFNekB5d4O4dpLqFC9LTMYMtq1HP
HnFhM50nKksx8N2yJH5sCEzo6455zk1ZYZQGh9Ax+8PG4YMVxY4seH29V3immsCTU5WgRUGDyYIB
CTnPo5oqALZkfyMIe8xMz0hO00xn9DwdUXDYMUAuzYwFqaHUPI4egaPTXzrY1Goz520tk/9nzcMZ
Q9bCmfqkQtpq8pyteJzQxhXxfJeVFQwrXZo4LC3p2VB/gajAVWfpdJpWqlSAz6GG8sI5lPIMN0bm
Asz7/nxLqvueXbzfDs+hFxBBgYPtenIpqlY4YdnMp+vM4WoD9MnAs2TtRTHyBA7eTC9LFnpVnUq6
9RcuifHRuItMbdSX0v3jOg6SFlH3iU6gX7sA8bsnq7acRqjdBoMDxQcJP5anEawcl7KgdGbxsJcx
GdyRA8E1dfml1z2gstQBh2qP8WaVp0kJ5bRt0IzwZiYmnp9x7zNwBladgia2Pyvd4cem2D816cIb
XrhIglBir2ffvisuQ5RQAfdJayz0veQKyATAjqSFYbPRTSkY/EWKKWsrCCmkTGHy5YRiDHqcgi/b
Cxfrd9uw/4sLqG2aMHwSy3YHVHmkpRE15CL3RTT1+TbNnzZqFbOCDPAZZBge68YWJ+BaQ77fe6tC
t+jw3AZx9tLXwJiL6fuXOpsTD4OjRZJhDQmcQqUz+urWg5l9S78fCpSkBLkN7o7l/gXvW8LPdU1T
xcpVJA7OoAFzqBWbA5BzEtWNQypX+Az+NpwVTyrKHz4culAyWyfGggwOBjRHuA6fbZuwxsTbbN0V
ilzZDZ4hkPtQCiKyDWmKS4NPUVKJ402VnyT3scxvdFPSOZiHojLr9qoPaavdqPWb8DZGoHD+xBH5
Ud5HwQ5WXaBzprrAP7oNT+CCEMYbIbSSPRbllBw80IyFuY6a8hTJwfkslJKNsjy/HDhq30BS7asj
ahvPlklteoGU93Xfl5tzQvFRNAmyEItfTgopBsvfoZonMbyTpPR+tiGxyo8cYQIdNDcLfypTmHAM
xM5mBcuQOgLLZXUw6qi8fNTrvhtcVn8GUkKm2yIgQ8zZ2JFu+f0q3UjN2eMLBsgja0PTOYeaCB/G
FAGb8Lt7ag/EBeSAR3DWlbBMI+4ZmLR0Dyu27cL7jHhqMQryG/QWOGV0n70JvBKP9QQ3ZiJh+Zbw
svZdjrsAakeD91WM++L5clHEoqN2NFf8qNxLKCox3WK7zZ0RwMx9Z00MMY5oXdmDgXoi4X9gQsM7
bWAqMIbGzqrJyvKGRzizdXVpMJg2tAwMFRA5V8PVh+x630DbLcsuqP1+2+CrLBp6o6rfFbdHOkMw
Fsw8engeyIAUL7Gn+tZ51KT2itrvoGkqYbgoCIkNnlM1ggjdaY08cnZiki+BlN2vqOCFFHzrFppp
rDJqjxrHYa40dHlBSLUNX4Egp8ndzB0866K2eQpO/KaHCtqNvhatGMKqF9EdqENo8Z//lg4vSGSt
gMtA5rDIj9BLlaVEUrbj2i4CltCJmOpJ11P7BVupsjwmFjPbqDbM/RbvwahCe1wuv37q7KdbiAnp
gVs7he7hPtPD1gHrjyCd0z01EhIogr0NvPYjE7ez0EaZqunOxQYOkWxYvppbm8Xy0hUNx6cgFCbP
MYXQ2lrAAzwfWrippCrmPXefvy7RK2dJQ3lZksiQ0nm6IqgeODRn+sIuBglSPidKDPyxyr89sARZ
sYuptuh7/btpQOa2HWK0e3ixN6jpmBRVbW2cWz3Bgjnm8+H/rwY1xmcVwZYXzG6Oh6DU54ZBX42y
MgAqRZn95o/4nO7ztb9ntbHM2qGIqE68/XJNKmu+/YFaPgil8g99mRGbUG2UZ2CBGDvQwolLPHFi
zp6ewgde9d3Y47EL2ulgL6G+SYxgjtwB+L2iBpRJA417D9GI5kHCWIO2CR/pHeZzm3Mxjjl91WOt
BlTKNcNi/bBUAas97WGT0pe91ESYoG8jlkLA7YEa5oVKN5/HKOJ/2o0//R3z9e51+d4TT65gAeKd
TnAykyMWebf5Gn5ApgGYJBufaTgyJQrtpCC3SOVsAgwwSI53PV+2vOGEMKwtcLQuPZHd9kY8vCLL
AQgtc4SZ3PpR+0Jv+877m9LuJY15NgYeyrgofpF50g7MrmgflaIjhZlPSSN77eWaRcPDbultgSyD
iUvXAf8d42+qQdBdQaL3HCkUmp1pe9wfMy2urQZrrVv3rtaVRvaAy8hXDZTi9NMvMIwqmMD5Im0e
Zwb5Eg6HG07CtMxpsd7hpDpfvdHlQpgCcQRU1zDpCZOYSNTxkJXpushZmQY+p1FhnSo0kWRG7GsS
xM5V6gOTJO2PdUvecUxsvFk+MnBGK7mwv7p4M2ANpXy81j7q3EBP5TLDYweo77wV06y+7PNuiApk
L2Dv9b8OcRSRhIOtObHV0LOCEAwqaXcNI81oCg/ZxcmJ5hEujdHGQsugf2J7tROBh5Xn30Kluzhf
6lGCbcVT4H/2mpNR2nDSVkfjDvl6X1YEP6ZcJGIDGbGPra8HGEW0/g5q2aTNhH0ZtzGco53BTgoB
MRUnd0tP+/LL36uaNS0ax5xH6hoD7YgJMJOAphtnSPEekAXPzZgp/c7Wy88L7eoeOBpeJx45MzAv
jdgApZX4Ki7zSUiWo4G5JAPp6hGbN6Ddn2iuLf+Pg+FQP8dy/jHES/ZFEe1b+fvbpQ+PS4dp85xw
oGPOoay6LtLXaa5aNjg4umewjy4IwF62RNY5kkTyV2nz6+lKqaOWrD2QgEuvvedLvndeAFPuRtJk
7I+AtIWe8M8Q6NPCqE1FyaTNPhpByODRwq7WupWKkcYl4kCuDMMhK4C9ZpQUO2B5gdRZtvY8SmCL
L/t7jAS/JdHpg+6rVCwznDtgZaJInKc4CwWJpjeIZsoG0IrRWY95p+hVMynQTxi3aoKf+neHIWKn
jbTCuDcKLgE/GBL8SOtrIPbwAWSFkT6z1DdXgf4mxxql4w8GRB5uHJ9+j3RlCVUAPCTzUo1KI/ao
KACmgzN6XIcD+4ELUWR7bDAfyM2FWjzdm7jtYqZOqZEHh50MNTL2vBSLgkPGjvn4woLAdK7aqCG1
4UVigveliXkt7lzywV8jdqiIyypIEOora6+99Iyo1ggSFu0BvVP5NI8w+RgdTg4TtxK4t2643zPw
6RmD179sPielSniqYLa5ozSwJu7bfBZ5K8um5ct/K/4Mv0L5DQ0WHu270R9y6YAwEyJPDfzEaa7W
Ti6aKmRuvBdbBvC4HEobVv0MASpaQfjw+/Ftsw2Nzra47HeTp8POQ2iZd+NdtF5TtQk+fxy/bZe0
/OWa2RFfy8DgJIXHnm1o0ua+4wWyHLnlmutXVI+ltQjuyRHdJuxm1c9G7PC8QqdMUkA+80rEnh/y
HyS4QRRmnlXHe/z7KDIJ2VsvjNoP243mFjZXuaV7tnNeZBBgzJKkmVHC9mohk09m67/m2MS5cDHB
ER4a2NxAwBtZaMNIvcJyTRFOMje9DkRESmHbXDieu2wSciPM+Y4rs7v78iK1PmwFuFUUE4ig8sBe
6f3mwrTLCkrKmns7vOCknW7b2o9PwLNaof7lj0xjqeLkpru73WEoFILpjTXy/jM/DVaJ8r88WUuS
RE9qgfLLYFFKYA4TobuUyIICbKFLnAVwJYWH3/zOgxKJI0Vl3Ro1SDLIu7mtqhWXmT/RTRGLNWCt
HgqW8JiAKafpb4Y3LOl5t7MI7tKgL4B43/hI9EsjsJn+hPB1lR9PE6M3moE6MMKVe8GyFB45hwwQ
RxhXq6r9Vaf6LV+pcvfqC47IUCOO5obgOT6x41ieolgLYcDQ/eEDHOYJHPB3rv2rGk87Gmm1ckMV
rssZPT+ZoaXzVVdMnEVckMY8ni0z3pJ1FMR4ou7h9SuqUygepOHznGf+eFlGSM4Fry2OJgoURgT4
eovsdodp6xoEx0VA92Fq3QeAGBBDoVDFj0CFdbML6QJqsTVwRH1BF/Wy+LwWbeOUp3dzlihAn2Lh
SyfAL1wnAsYLFnaHkX+R/N5nPuy7rnAYoi3M3eA9Q/WoulXPxuD+wsZHgk7ZPOCGhbJwhIwx+kUM
bDNW1ztsFx+4HOo2yZePyP41Rz94Fa2cc7RtKv9XgGLusLHZbOM1MyuVTWrlELgUIo2syzjPOfki
Su3TnngdfexpfxQxtYgH4KrG54/MEIhN6W0MRomgpqF+zoHeT96phpxHx9QyKBh/q3e2otXwJdPF
d0nC509XAi35kw+6gxr4hhTRopiqb3+A71SFupKFqePfyex9NGnhBSLZDM1RsSQuYZvTFl5XMYFc
cdBLQqlGpOc86SebFXiwu4THHbrvNZjm4hZ5JfR4zbI7OwQpad1s7UVWTEB+54kvBPZFnOoPyTl4
eD0EtIPY+h9miMjjfU8pXcnoMy3TSD2LTd8VUsGR0pQfoL04hFNqIyivrwZFA4JaCggzpxQybx9I
5Avom4z8UYwFbclmJibIS5LffZuj05rWc4yROh4w8QnZFaqvGmtyWKfj+83GA0j6b+CGpyNXkDE4
x4hmsuCkFI11LYAex91WFaCkAsaoWjZ3oYtf6iWsDplyAOUXqktXtXnHa5EHy6u3WgWmBbRCDcK2
izV8MbQt15c18s6vGRfiqpOJw0NNcyW9e60/BmpuKSO1Po52FHcLcCRlo7Xfdjrvx7QOHQPn0F1x
SYJwNX4e41TWjL3I7scDDYHrbCMabAMSqlV7GH5+sFkziGsqMbjvD0T8RVeDYZF21rriMYC7wymp
ouh7DSmv8+Nr+AahQAJcEvg1brUJ8Puj90ljf1bhznYwm7eURK2C+NtlI1mKA/iWtpDlVWzL2KmZ
bmnCutaTYNbThJPbB+8cTUjjE5OhLLvjOTFTPm8swkE6e7qnzK5Kigg0s/tddFWjdlCbaNRgC5SU
5MMpvQ2oHm5g1voIW20AIbCV6PyFnedJNU9ElO+WUnXTTOU1mjFlLml6N34P28Zo18wcPEsy4mkr
9+iUkwSxeOakXnycyxdsm2PKvYff3qMz8GIEw4VUiWKrm17smZfBokRx4vgHMPXtwcq19RBFLIvZ
i55vJ2VMRpgsqz1DeP0A2AXnRi+/muHA598a21f56jStqP/mrFn4SzqymzFtWOalkQQmgWfcRcdW
2PHiq09DlhZ4cq86V5xQU1snJ8gJv0OatPssb4Vf7gNoGCn6VABM3P+6rp5w61cdeMT3xcdUzJ0k
z+YJ5FzNl1eadaQC+DlSYaSuZTHVLKpCKKvXRI7u+T25jJkxfoRt5HnZj3e8+3QjusY7qgIyc3C+
0E5HMw9AJWi1o2+I2QqWu0ZEARZCJV7Sf3LD+Un8ZRnO06WSS0S/51FF7EB00smzuCAFMEj91Sox
AAIygGqNEyMZ70x5eGfR+XBegb/tbXhO2c6wvEWR+ypnJ69iPfb5nSsFzwAT++o/W+R6Is7l3G6S
Ahsi6lX8Q+yqC9rC/UUgqlpW2N31rfFJ7N6O84K5iWVRAJZ+te34ItucQwD0X8nwhPtfWRbmMrQy
aRZj+zP7LNAKl7mzo2/+dUpyd/S2QlAZ4kfGWmk9N9mZ80K1LDYAiB6kzKCTGIdn05msJ+mgkvjR
5WBkiTZR0LDTiVZgCYDyEfbgiIepz6SclVhX5xQt1I06Serz+O7DAG1BA85SjxhVBlzfQhwK3M4y
u4fmXQcsqa07rel6tG3dXj5HL+f2mZiz3Lzq8rhBMIKVvd34FSpFAtnHM0KZP+qbs7z5WjrnA8AF
WtaZF/vtO9S0lHl7sG1k1xsBJeFmhTuV+H9qBwnWTeUgt5x7EmvTQMx/p2SNJCJGrWibe1x+o9B+
60thHi2+ME7Ff4ecEXd+wBFHg4U/DpNbERbGQi0MmxbN6MsxkiVt6PalX4tc6FcYj5uzVSq9aDFg
MRGwDm8avSx+AG0UXgy2QVm+R4n8j1lzFHEX3Uzn3tzMtq66676qi4zDoxz2MC53TnyFwY13ZkDP
Mr32+Iodxaq1Rn943nq23WrZJdwtjNdRzgIipPafENPKQZ2f1Z+FvCcSc3tSlxsumR/dozJDsc0R
unJpJC+8MqNjrPSIghol4MeqetO1JCoAd7b6C5Vxm2dvK2jK2+jigXk3Hz317L/Ff5gFsL6iocmd
V4ycRV+SWgjSsF96InPDg9FPUhPt62RvIipu/3dYfuvybciJPm5q8lMg2X7H71eKdbtEStCU/B6b
+Tsk4/mSQYKxhx4I3tMuD+jiG0uzUfxM6izfp2u1aLJk91LIoBDA1rrEfOkRNBAN9y3x/hgjDrbI
Gzg4rirlIjhotoUCLMWjr3FUOIkUsC/SYXRW2SiYmAfzvvH5yirZpBKMkb2xxS6K6Psc2hnpKt9v
jbrjqNRMhBRDSPLrg+5moWGHkkajIu0iqyaX4dKKlRNbKqt5mniPsLjaP2PFHkYH85MkWaYGSX6P
JQ7JzEuui9YNqZkEET9b+LRa6MJGMVw/lri2+YYqnEQR2Owb59nXLnapCXvxwGGDP5yBGGrKnzK8
kWlBiT9vkbxLlb5rpig1ZZUpVoAkHbpqmkU4X3Aw138n4B9J0a0PTSHmtmdgzkGN0eoBT1Fh9y8b
QgEfce3YmaJnqv42WcOPxqrcBFt1SPUsCdHwa3xmDOI1FrXZQIveZKcVhBccGKN4OOgJHWv0fHwf
M8Be/RegNd37Ws7qyDbMBI+wAYr6oE4M7q9OpLyNWjbr/egv9jmFCLhR+N6nUpGOzd1DbR88ZrYp
/knjlBXKtmqCcd3Z8N4KpnfS0d61WnDE1Xw+32HmUKYuanRfZiTPUaL9fVBXNogY2FNgl0rYmPCm
C1Nvj/odzjBDKgHa/5QOKIQeVU5o1BPLFkJOqf5/C+LsQ+dqz+12zJxpCmnlBFiGUUxbyv7rqEIv
BpU85jfvjwZ2+WK0smwJSy6IsxKo4HKpaaj8oHwnUGouRIIdOANh7lw/3J8j8JsNAYRET98NQrIO
6YVO0KgC/XJfqzK0OpzdKslqilijIhV9nndrsksgBnXODQctRi74m2519gbuccytFlM+vv0I9eXW
75xo/VmW7R+XZX0ZKwqwvDc9PbkMZbq5ACXqiWvnboLt1kM4q09JomKUgPN0s+DOc4ZRWgLN/O8v
+9+1UVrkKfLjP37c6Pp9lkdwYqgQHGGU+BuLAT0mH0F6+vyrUC2sBZaiN4LOXMeeZSVlKjpHFRwp
1OxjgDxRbTAgjKGeHsX+tO1oFPje80v9Jr+kaurJLj/5CmUJSqoK8cWvoKkXNwLRYrYpJqOf752w
SrKFurV0JoDTi+egeRXEtljiPn84C+xzdgeZS3pu1gM0QghlweQwFA3w4zXYnLENo+x52WII1S5b
Nfqn7tFG1yrleV/6U3/sZq6xS0hSOrHDf0gMELCM5s7ZaI5v31LfRHFOPMSno5dBC4f43k3O/6V8
QCMNYaVJyMI8YnhoU3wMF1R1EOc0AXEX2oc+xBGWd14xXSirdpwzjqKNV4OzJFK+bvKCqU9wjL8x
l/8E59OeBcoRA2fF2/X0M9+DUZntPdIVlCbZSydMKInnCcrdjzBDplcBleS9S6fhgaiIopQDEPYU
f1u96hTHot61l9HnTWtbkwfAaY8T90Z0z8nEHKlmnTdwoOftSB+aoJXPrRxMFam6TEeiKEePQklm
i4RWvBO4U82gxQCtBraFANcUEQTiPKu7lFRb9pv3lraLhRWidqEgAGDa7E9tIpnWung5uMmKGGqH
xNAS92lSO8yVNkU1vhS+yCaRyrEnwt+pNurLqPokTX2IN7G3AewmH02PPYcncZvF6jRsuvyI7umP
WaqSzqPBCj5Z7ziLtPI04camdkzlVvTYOcxhjER3cl7+goGRqyemePQGE2YX0FCCaf2RqdPcBuOh
+PuSWx0X2/P94PTefS/H3DTNn1FvrDY17o6qFHaUwZYvOTaS2Rttg32cqFBNPNVMnlZmZmKRurYV
xyEEE7K2/SbJDV+wAaXkJ/POzBDPMSYftrJB2k/5UPeAXIw1PNcC2t/MRKmR2AnheU1IRUIFUNy1
AFTVxosqBSPvIwyMJYj9SaLEuB5gSaMCnxa/FNU/xODalO3PxOk7RHt+qBGmZDSb7WpRROPqH3xf
U+w7wXzG8ctOIDpAAPyPGVyLyKkEh+/cMLf64m+gnOcgocYnHT3ZVRFZuCYPYz/ZE7P3mhFsKxL9
piRHBZVCgxfOSlDJBPEDjwlqSfQkFxgZ9722rCUGWI3DgFq1EWD9g+BnxkPdTCqMpzg9o+3bckId
kfRL67HgQ2s9M9QFm56gNlAc9OI/gxAPsp5FWu4xCqMkngb6E5oCcyd5Wt2eC0FW7dP7Ff55H+/5
QcRyNEcrghoHxcE9tc+GBjulDHVvjumnAieogPU2PI+mc3JfrvXFbYm1tWZ8/Ujyct3DNNQe76Y/
Q3G5ke72jJ/hsn/upKD2B6gpB37awoIsdv7QYmevKDhcU4md0eHav1G+VxJHOsO3fUKvOP2tH6cM
+wQdOI/n5cGZaMh9q7fuy3/0xMYXX0ErD7mJu1askKsUzrpTIKIw6OGGaPANOHA19OGYyrwtmGpY
M0Bcb53H0QUHkdlugdbcZyoBIOloB17iF4tAbjK1GB6Y9R9fHiqQVR08RNr0DBlEqcI6p9EOYlrH
7rUcbpCVwviNOKHBsXTRiIcmqrPTa4ZogUJ/qRqW4nbGRGJr5ThE0HFhbmV45oe1bYomxyJuSfU2
2I1qLD2++VQeP+3K2nvx87vm2qbU+5g8lbxgH3WtPdspoWdqqYqQc60OjVmGFn8MxNAsAvKWwVUL
UuwmnVo38a5bWSe/e3oiDy7VRps1DDHimIhBF8YEfftxAtEjrIArHVq5+xQlKm409/D5VZEsivW3
R3m7HweSHjg1wGCJHTiT/rVlt15jZE8Nyv3kY8a1t8D4HRDg3g9o/OBfHWMSf5aMWCaeRtUNxqhz
XBQCz/fGG/5HKjhVVgIn7DMPV949pbnPLr8lBm+dvjNBjfBNx4BnGIOQVwqac491cVJ7IGQ9NOou
JJkVMxIhI6cxIELQubK5kth9M490BNvTbdSOtWQKwoy6nf1QQHGtfZ4xQjuPP9147MREwj5lcfmJ
hEwNZqbJNE0bdzc0LMHI+voJcZkipCx495NtrpTCKelN90fIm/ztTqmZaI3FT69++FsUPmx0rkLm
WvmbiWRwDyxf/7mnT5hLrm6jiEJvJ67cFD4zL2hywm1O1txL3OGCY0atei3EZryslrY9N+f5QIRO
2iTPB+mOgwuDZGP3H1UrRFGCW2+8WT//JQAFs/XL5TlAxh+guM0KdmsmjpnwsTP2hMvR1MC/vEsV
QD+wY43Gy4KxUr0f6jl7WNIR1SeXcURb+OLhT67LZNxkT7mrknOpbj7dmSOYzz0TB5iYmTBa3Z9v
KuXdt8u7eU3hK/GOTFOo11tiaK28fsadrFY5nhDIFQZn5U2wgw+BwIi1+LVdGJfrd6QuhXhfjLbT
RZ3l8RBfeo2v1Is9FkfeMbJVDnfeQjdGB0S7yA/ziAM0a1t9lX7HoQrKCYGtXlno9HsDuRF+TR2o
ABukahI//ciDkueCE/AywI/iQ+zZGaBKTMmWMxYOcr8g3WTK5+Xw92Nk9KX9iYOW9Km5R7k/27+l
Qaz5rHdnJcBCWV2T0bGDZlV8X+K2mBVBR2+D+CCG46YrJUXUuyTDPqVatf5jYxyadiL7gmOI376C
a6mZGCmhN5ZjMsb4LhjCZ8gK3RYmWenqcjUBOxIxOoCXm1gQdGdKQw470oZkobtHSB0MZpDynMZt
+cZ6M6MjTp/TVNoXSHUe8XzPg72N1/ffrVr8QUaCaVT69lJ76kaLYMtQJYP8XyqlhPU4V8VnQOA/
3nhc6pORDfQF7sosiWvAL+A4GjqxDf19+EU8/D62x05sPmDyBTaQpWJtzWskSG4B16rDJ/DBy6nH
cmxcdkh6oTeY4+wyItu81BUsTaqmxJQySGTB0TR86KEWK0lRvW8pC30owsAjDivlp+scTduLQQ9N
+Im7xGjQVr7cBz/1Sse+qBmruBqPa2M2cplN4V04fdX2k38BFgjxmYtWneyejlb/DAkG4OjAV/wN
eTO1CzhjO5ykuPJIljA85AhykqxXN8x44cVOipPJBa6TzqbApliZLQsJ6e6S8vYYMbFk+0CqlOZv
MLienSS3ZJuuCDfAygVf0Q2d86m8V6u/PspzdVjwnMC21VzhnupK/oiwaUyln3F8LrV+WTbouMaB
cgfq846yEYhBofK4TFqzxL6/3ROYMSoPO0WdNapJvRNGVgDU6QOxmKTqYi844xsnG41oSIOZbAV4
27jNAvukfnwmIs/cYVyOX1oNsDxSJRhDDwAOLl67pjeKlPUUFx3si09RRY1a8DveNjjVoZa58EI+
fzdCPQe6Xy7T12BZjsd3WXIBqEpWgoXKaulpndEUALQdU53GypcuzXioOQg/eZMx93wO2YnPkmU+
KuadK/BsUC6tRWLkON6wL+k3iHPg3uRyfV4YL6DdRfZCbBavZoNKUcSXxiIQllyRUqcay2U46w1y
KoLFw7ljsRo0ff6jKkFkYm+VU7woBj3/+XwmJkMLayjVteM1sWkW+MzmTeUY7G30eZy98PJTBS0B
pd27oqNGphpIuV9bx7V8qxUCBiJVUYyQs2JfmCo7dMRD020jPFbU2BiewWJ1/iAyWGrie1SiMhBT
C0rI8IX0N89Ux0cI9RYhRaNdR05NSO1ZueAVwaLuvbFh6r/pKgsccRLaZuK/+8gDtVZZBRsQsS0q
ow1GnOB+lE5biUOWFxVRQzV9RBDgH/J725Y8DDM6vkg0Y7yRWAHv9M19evcjMe1C9I243raEZfRM
iyMVkR8Taufo3ZIGrUQelyTz2MlafuZuiBaY4jyWjncoFDXbeo6qYl7oEbD/vsKtQc9qGHuw/WLn
xq/v5kXbSS0nLQ7yLQUc4LHE24tgBBXRS9X2L+4+BSwwgUd7wJBsJmnH3IlMx+G2ozPp90/Riw9p
2u8HyxPXL38/1nZF/6mLDjWbrf4HQ1vhb3JPwrCzvMMhs6hPJJ1o5jx7p95TYNs3oXlJrDwBVeFf
42tbGd6F7/EvOd71BJa+kSqiyrlNzbdWaOucsBp6kF1YMnrGgxHXTDMjI77A00SuI0lD1shLBhXc
8sKYbpsNEaPZPnGBMzLrvVbEWwDYnuqwAi1NCBVmqDhGhnD3AzOyFC/lyzxd4v5n1MRfZ3pN3Nmy
2PnchBrP4qL2M3leXqlWaGVI0vO+9vlwoadCfT4noH3A5i17Djhc715CoC2keb2Ow7YQWmMs0iDx
mU6YH2wjJXOTLxwTHrKu48j7MKHUMDWVSVhejVu0g63gvyRhALTX38p80EUN8/+tGW+SmMcdYQAG
1xY3wLt5gcF7CUib3pYSsNnldGhDgK3HpYp+1fAerZJVbiuKNyewe7IRATtjg+Sfii9PeouoUAal
eEKa1guY9/d34L4RbY6ka0BNsnZXdRWsxwxUKgAdVtAUOj0VXNh1us5FmgFo4lWltVCYDQnNFYWx
qlXYvH3FY1udl4ym7L3L0OLy6trCY6FbeJeF/74jJQb+crt67No7K2ec3gnoHIHbufrUF/vxQ0+8
1Bpuv8rRaAfe7r6rVzTRo3a8BwRTDK/UfavjIxMNGPK8orTRpi54IVmfLCJlFc40dPNvFDrxOz90
NdC0Bmb7apEuHd/KLFxnzsC68OKH5D70eIWspdSS2a2WfkuAlvZnQTmgPeJ2v6P6jP9MrI16lT+k
2WC9fbPYiCpQOkPUXvfNWXfMjfMr90dfJCZ2GaLydGRYXeQWKYUURED7ndaIorA/Q8Qy59ozNfQr
YNvqnZpKsfxSA4dqoznAqvwjk1nxGAEnG7iiXi+oKQFZQJRfa9fsBqbWjbPEhUcF+rnM9oOF3fhR
IX9RW1XvcB1kB2TRbu9kdyjbeSXUWv+Z57v7aHMioTokbPW24dwTJR6guFh0+d1uLZh1QhY9LXMn
AYNlaxiqyzb0+hZTODNwCaTamI2MznJYZHo8RilBi4jIbwLh8hX8Cn7bpvDCtha0QNi0tgabCw/2
8ZneBhV6OWEjtANE3maiyPW1ShpqC5GOZcyQ+W3KkowC9YZFqJfIBM/sVvjbAI+3Y9G7lNvopnZI
Na0Ze/EkfWh+Exiy5/pkXVh2u+yzhBC6PRnTxl2xXwCy2uLVL5+Kzl2apoLZ0OmKGTrzbf9w35V7
JZFIrHHrf2Z6D9ZqrxXcT41EUP5q2EvlFQvapxTGmA3WPWkixX/IcpNjfCk1w5ofx71vr95edkLj
HRlOrMmvr6Ny53Itxk8M2qgwXXdzfpaVSheD5ysvI9QIs7Baovcfa9R5w+5gQh8ZRjBTh4Orrl64
QTDiHqIc4htD1IITpPMCFemmgCGKFKZo58vCNMYWXtWu34ZN+5GLs76Ld2b/3H/NMv/kGsyMJNSb
aafBIBV5/QuyUr7VWrUKKW5hEDdl1ky2EZsVMMy9puJgT742yVd29yDQZiXi9ReopTfRKo9Fiyr0
C8eEbBFbS7jY99FLBmY3qOQA9nYLHE1aBjry7vq11DzHAb9cRNvxBVm5x1QCFm2xECOWxjPAkYfI
ZuCE0SAahFvjKsiLWxGJgRJSac9pl/vUT46+h1+AMAXYv7h2FNoqX3utQu8bcs3GLVPOhot0DBV0
NXmUrXLprvvRpKHEzirOLvNvBcTuFzdCY7l3KHZZI4MnvukwdI3ccQqeNsCGOBTEyXSR5+/bbgJy
pv8liazNj3aPy18y90wKveqdXd6MaDv++e6fm7Ebjbbz99h3cyYckCFsKpOn5+uo7gzx6CkduAFl
QWZg69k+vdouUIkrD7qYLqnV6PQkQDbV6ntsPKAFkEhseC4xj/DAkdNieYjMxno/ZF3lVWUrzqlA
cwnTc1uSqbI7rahk7mYRIALyzGm6vf+XZcz2JcDDHZToESKUYXdFGl6FmlBOIB3Eeeverk/VKr6G
r5d9P1i2FI013+7cIIHO2+SrMvyN/ltRBAQYhwnEY5f6ZglRe4fAqLdn2ILot3gFLYF9vMI/qhzQ
WSthxLOgWuGgZpxlsZknaHG46Z/6SjyoK01cpGX0ZreX5Z6Ck+YaoZnz9fCURysGRDe5yVcDPLQG
RNJ+/qNvC+F2gFJlED+40aBIiILtPOkBOApYtLFpsJQrSTmkoIDfa6p1yonghSNm1MlmPXzdNKpR
VIsYrDQ1yBWoiwCHq0thl0BEMZFrZ5uRpneHh5K0SjF2/OuS6M2BxByI5kLMRkgAauTB4tVhJ+po
ywX3HsbNZZRA463rn+Xau5JrvDAn9yMHsJvQOoAKa4ZWQ+mspKtsFXnnPLbBlEQM83wcBINFHtnR
DmnZQnADiXnagKTRD5ClOTtwzp4ByoPNoRe6ctibLAr/pTA1RmYe/sCEosThJop+2SGhOzyehIdQ
cNAVVTEHXKmMcrKaRv54bspUYYuj5eXk5qTB0FpPHWSJE9BvWB/S7JP2jgnix/IVCr5SrG0HwTBz
irRC+i0vt1YaHubH6MV3imj219uR8P75e7LYKawpm6CpiCEVapklHh3hXFSldkMwTMvLs+4rrotD
zFMX8oOPDyz+C/m6PkHP2AxbaW6FcxscYzzMnj2nVtviCzhteBljI44ZnH68j1NFk3xk+q+Jfrud
OH3J6x8R/mrI1PC3BlF67NDBMDPrZ+pHmVEoJS4mKfGEqwLs9s2EYiLUQR0AVT/NTm0GBrO7fGl9
4GadJfNLFvxolj8Chke9QLmZcFGyFENQ5VMclus/qNKd+7wwzLKJB0Vp7tkCIVaiMuKw9qAkwkaB
c8PVdaxjpZGi/QZ8nnGXQ36St8PQEWkuuhOUwHKclCbVQ3IUY5MoUc0ZOC20GdRfzQJFpCQl1OM7
cNFBwlOG2g9okUh2hrQK9zAe+0Zviji0E829w1GDRaBw3pna75GpX2jvUnsMCZsfjRvfGo28bI2K
LbSx85LpXyz0apo8e+KmJ2mzwBAhqKoeP7wkJ496ZLHWpXsjVYVpBatvfW33NLs6qPvHAXSBrfiS
Fd7vSFd8xu4/Jea+ej/SeXWFNBDu8TT1rb+Wi3HLBuz/z0iMhcYsH4SFWnmhccayFUbIt5fIi5QK
5xjevrsu+FcfXz8PnZv6nQrTSwz5ENERCjlqDrOuJx+3cFViepeXag6CPzA9esyXPpZjvjTyaGf4
gYv1v5j+mcymlO1ym0XHjAu0ypPnhWPTJBTDktUIlLL8Mw81Uicm0/b4e3Z4zUd+CR/s3KUNTxGK
M/WHFW3CyTbltfuxh7g8uuM14ZyOQQrfY2ThNh1fNzj3GypvjONguK45/QVmfpy9zRxFFmbVDzDz
WjuNn/EJmOK3l03WuL2aOEzlA9WtD4FJZIWpMX4PVDt30upa1ZbJAaCH2tg+Gj1+3w/Ae5I6+U6p
7Thmlt6ppHpNQkC+e3Ogryuglf4EWrMaEXTukQ5FqbY4s4pFKi0wrS8CK1U/qM6xUgzqzkt7whk0
fUqd+BRIH4YEY5H4X53zha7CNUT/MtVy92kN9FUMHmp7qI8KNpa/x0y79IdtUGvnGUC7OgUR1vrS
1eXZxktZV9eZ6bDR512da1jD/oyAJ217RMm5o4lS215TBMFhwE9s9cjHJ4rCAyZsY7LTupO5mxMf
tuVUipxx/MkDcESxHaW+lyTJEVK78TMg6uXaQct3TbMFD8IVBQsH0y68yaILJba28Gn5bu09NmN/
4T8qpebjAMbe3zgJRz75M1OoSnYMG+0r4oySDU4snRUuGJjZ5cvD2Mh+4gUcx2nmbml0TMxtSib4
oZ8nCQoRSIvz0ompxSz+XH2tHLzH+xoYg8tm56b13EZaiRachrk8WX72HLSUEvzI+NCRK+s1hNKg
DzFqVR71f1JNuCkDPVh6afAeyTTplK1GJOAV+Ghz0fbpQ1mjzkZRnGn6ysLD8sqng8/qKsge4nrT
J/eKh8yBJKCYxmE08niZ1C9/ETdIazAcfQqsbyb3UGvFHnzuOGmpvoCP3XF2wNxGpscCeiXMTQEU
2vu39nS7lNGErTYVIUQ3EMPThUdhPph53WLWsFTyUORHnQ+dMpBKHt9Aa++VAFs2/WG4Ds2TFaA2
xlVEKtZIRhDHuVYRlKUOVAOhNUAHOJO5aR+6mNNyV0Q0P7C8Ndz5y4plY4vfIMGzIcVjQCmJ6Vt2
E3UWkyrYuK0IzPWkcWUCxFIPH35OMjcPFhAR4tOrROkXjrXEqdo4QxTJBUkD+ZNnQwttJFJStzlD
aHOOjawTHYkfW7ySkPG9Uih9m8pO7bmpbf7A71wViYj81H9YCUzHKvkCt24bF4Gta64OXBUF626J
rOVadgOTSxO49eHt1rCl6KhAELUjFH+MdMf9DbUXcpX9icpwFhKfSq/KdSFrhdZWYUcRv3WOQ/jP
WrJFz7Ve6VKwhcRjE8yVYYsUVXukOU4g6/cAiUbZ0xcUp9whPEazSlVR3b+e3w/jELSFVUea0m96
1GUk+FyJYiL3FKDY6Muh4A8tEji08WG0iY3BVSIlJbZPronRQFwwYFBmQY2rP5tJWJdwrkgiJEW3
n4VBIWBzNyJaLM0hp4mQGhdXG/Aabpc06QmA4bIiOlMTzT7LCW0bQgo9yjSSyShY6iadQoYSevFy
o1L7W5FqmPXgfUYqH3faYZmoNlB6o+oSiKxPJO2fJoTxCTaKX2Gf2K0X1qDuVXHEGESa3ngR9jVY
DMXuEC1FnzIEyFYMLqo+nGdf3p/PGrkBGwJIrO5kpOpEsrxHeB7IK83cK7eq8ZW7cMqNFOTmi57D
JFoZpK9sbq5Pg5ieUlmn9BZPtrNW+J9v5rao22oM2IiptxJPGKYDnde8WYYmKhVnnrUDJMXjQVGA
fTQeJzq6NpFs7e0LBFbSXUiyZJbp1HS1lREh7WOUaIyYoZb2wO44t58UQOy1fOmz8KwZfM/McwjP
xzFeYSauam7jUBX0XJl2QUto9EEE+eFKWgH+1vNfzRolILAykHnqmLI5PMb+tVq87ULeCAXPiXSU
0HLbIGhqbbSeF/5O6ni+I4KodOMoJNajMDrPUUF09vfAkLmM8PhBmo6uQf+u7mO/CkeDX6ecUb1R
YrBkVRRgPUmuBte0mcXoEG57z3IAbjK5qDC+GPeMqpaFGqQTdfBNh7m95M92uhVXOJes7W0MXUFq
83kSq2pbL/yOVZrxDPzAIcwrEnGsRz5XIQv/yCQWnOTRdJy2cCtH77X/bnO7LqbB4CSQ1iEovP3O
E2uzn7jmGe092+wb/emcX7ul6sH0RjCtW5Mp3G7ewbd6h8w1E3BYFm56+D0Q25bcjJhEpbP0EYNm
ktyI6R6kKSHpju7W8qgWH7MuDxRkyJEWX2V7o0qQ1uQzU/EmZmHySx0ubYZAbe97+8k9ABpzidRX
7J9zAMzFnxcrm1MjjiEI3AwcqtXNN55IDB5VDIPnoYkaioGJ37Tc/Pbf6QWPlyVKvzmyiFncAqwL
/YZnruWUWb++RbaJGAuUXtXgxf+TUblJZSP7SdRUuJHf1y1+Znwg65Y2FgKpUjvEToqmKnMqW/tL
6wG0pxdcVsCkdWk7A+65zigqSdg12hU1zx8/3kyT7o1+wUAR37miJTgIiQZ1EqnNEdtiTrCiQrjh
QpbZwDI25nBLKvs3u5V6cSVdGHTC1Mp5mjigPebJ8skIslRq3ji7jA5QW7yhtjHkY+Y1/4ACc8zu
RycYC3BRibqpHBdsBow2DDjeFYrCM/DdTdSCHxWCLKooJU6WrHwgMSyqirPs55lZ9FXzyVXY2uqY
A2iVmlJGkSCV0WPQM6SVdNm6rXbyh9L4GJ+Oqa86b98Tjzp8fjPT8tUEUmGv8XsQDlUzDJope7x2
KXgzMHx6M3aQAKgYYgMlQey1u8nDhwAhllAo2xhSnsiRFTm0d36WybgSbEsSCWqV5gMdYSfS+/3D
QFlHTyKEAtUuCGQRo1j2/uh3fSIQa62wEzYD5bHltGUUPSL3fku3Mm8JDXKfO1xgqO6RatptYfSA
Tj12jtmGGb85xTPWXR4pPjP42vHi/77PJl4eiwzTVzmbrROIhQOR/YUmvmeYKJQE6DENOwCxVpj6
CnYQltI0atVlawhySuXT3k+eLt7VAN8MSbnEqsBF5orInerkC2HDXWrHq0TROfX32D6EasTgTyOb
hpKJKP6EBImMDEhsTb90gXFKEoSwLXKvhBm7AM0h+12Tng4o5/iMyIB86TboRaKE8UmIsFGL+cZ9
oLlFbmJMTwN/uDabHwHQDNgpkDVK2ztQU+LBqbsLlCiubub1vT5f8RRqB3PMrGuKljB+w5DlgfUG
z14tbncSv7EeKlBFDCLphW3/T4jWTltrAUVnVv0jcVyKHHhYOE0j5deD0M8m/+PdNr3/P7PmnLYh
GXWLxkjfLEfYtdHjETImJj2QWLFgjEhU1hO/cJl9nYhNiuTjmnYf8OOEm39a78OZpF0gIw/7wYP4
PIGmfOmxnMoXm2yNfqTwbjPLZyj//RkFan4wEq3XWRSzOOF29mM1ZQhAjJSjI/QSjWZulpZYWxw+
3zIj6xCoRhtPEhwFZlaeB4pCi3ZXfoZLAsup7BrwgFsjzYjsQT64mk4IwINcTz6HjCUaQaCBO+tJ
iiXybpm4YfJ26f9/aVpAXlRhXBr6KE6hz5eDKn6yIKclMflcq3emAAlclMAAvUkYeWV/yBF7j9BI
KRjqMxjBFGfMIpkJBxBKIR/XPKG5T33RtnvWijA4iY+vQJ9jueGchhPwJbnY/okUypXZ/EZqOl+U
OzummpI8VLf4aO8154YMgKX9xghToaxcyZeY5avn1o1WCchO7AY+EbXUkmjHNaGkSleh5DV1Xjm/
k4oLzYKZ99icBvdcQCIC2WpcyBaeR9LBNnlE9i6xM3LthuVdkJX71Tz1oY7HdiAxnNuJWCgwRE4O
ST0Xe+tpFPr4G9tNlzT4KiDkXtWPD+fFOzRwEgqQbLltNlIKUf2ByVf+zMy7vcdOYHqt8f5t8gT9
ph/VSpMB8sKLQbjbYW8mhDdf1BxfqgMreAf5tqLId4HiGKj83koaXoRjDjubkxPKYDTfJ9JTryBA
yC4+zeZfTESuweyyGvON5zEI9GODTzxLlEKqz6rD1RPLd7z1NjyK/nUy7JFgZ37efQAG4ZZfPgAJ
DJ5YhF3bTp8byDl8/tOILaXF7OOee2GuBNwdRuyfx8kpa+eTQ6egB5KQf0zezwYK2Sov1ghvx/oa
3nu9RVe9gxbxLYpRUyWaVf1KeUYTRUJJH83DD4qCJaijl6CR75xbRcGnCm7i0oPqWX6yesiGjL4c
b3dt4OLLpCqVpvNLSygToP5f+iQpV30lniOS7Zcfh9M6soHFXp0ZsFutA3hQYSASnWjNbzafPfz0
fAWRpw4XoDkTHk0EQ9QVjEZ35nAmEGW5rSfYSy1J9xTl+VdNt0wiUYKZDmQnYekP81dtWuSn3Squ
ZXHOOEECJYnz3v7KC2YIJNxA6hJgGnZh7IZx233CQllKeoB5RuQxjaY3Wb/rAGzT+4ID8XrlEbsT
+Ohbo5K9fca9g4Gcoq+LqFd4xPFwvkyI0QRESkOKM9ioqKRiPSBGrywsvEsnH+0G8QLlFvdCoRV6
d2OOBeJzOp2UF1NpL1EWjMOUNshk7KO/jbg3FhunVehhlSNtlXS0Ko2C/jqFhTh1XOgdRojFQlfK
IpH/EyWn7a+s8XyimDBIhFaUgCOwz3wuR+o5KgwisbjHfufwBuSQCKBORtLRsvE0qB0WgRclBnqA
0bFUOBaxnLtMBE5B1TG9FsnOSDzFppWoHEF3kpuDkTgAEWbmr9FKH+MLRIG2EUQj9urC+xY0s3Zv
C2qjeXLjWBCUXWu1CYCN0vGyyct9qr7FosAoaasGsCpCiqqlVvd6QK2YnWapBiFSJfV6uyK+hlKh
R+bKPIM4++Tjr90XY32IMQJyIobrLMu0JCQz6lzk7d6fUw3jvcrIvNHs5OmPAoPS46Tp2v4hyZB1
3GFDuRjlOLzgjmyA9TbohgbmL6SJG+/W5Xf889D8vX0eFZXBS1dCDMjQlG5SXftNnYgQzrPENepr
FKvwTR2hpEXjuHITysi65M0/MJIeK2Q57iKwSs8M9YPMcoGxnQ2185kdh6MaU/BhXyMT8oed/6Dn
7bezBNday2niwZDbbU411sVd/NjcCNo9/llHM5eEV0LWUL0/80ExBMKUrmZ6V3203eI/sAb1rUuG
injP4b6TD8i2GX9XZN/PpbDfhUxkqqXXSC4XcpHC7FPEdQsVYpfGF+UAFaKLVJZD5Lz2d0WUgRFW
EP1Sr8SSJ0oMEmYYkXaw7uOrjcQQW2cNxx6N7FwmN7bz2/sxsw77tG2b4TfXcWD4AHVh3GfVFxyj
uqZ2HcvaOm5svWpjiDPoeD3iZkDOqxmoE91BXfeJjY3enJ24rdxB2yj5w0Gfjon54gujM2Ha8wgT
AZgtP4c+Q8U8Nywh4cK1PJmbgxlApCoNOC/rB5BnBvIg3SgmlvH55cPx4fKX0vZHMBSSnmu10487
991tttHJ8ppO4xkVsSQ427zTs2NhCz1h3gnFTlWwu+/6fIFQ+cfdiShX7i8EBU61y68YLC/AU1sI
L6WLjJrV8MSFrvnZQhnkTJb7SXCbCiJFoScNGRpa0GCSaWpXZ6yDt16CyVPQ2wHTrtaYADpWI/uk
CGBi/j+l9ugywIZwwqECWZ6fUkkAu7HGRJNHuZE9x2FAZG48iJRfG6Cg/ypxEELY2dA4fmVqmkUL
CC0uzBcHZYl98jJjKq9TbmzD3mfKTFddhqQiM69tvoF8ssejVSX8jkho7wckCmKUdaR+TY41skHB
+aEfkU343JAD21BOQeJkt770m7EKhmk0DRbIB5CQ9cwHu4jYXNUI+d3//cb7uDu/DxYorBTZPSRs
G4HRvVMtiPZmAx367MiLq4ONKmV5mU8Bb4JmKM1Hyb79phFR5CINoWNvFL7cC02NmU4exTLqlk/J
TFxRt5q3uasDh/sKs7ldjMKkyhl81msafa+/4rUzBzt0GDbIiidiAv3Nh6kAHB5mjtKTXIFfq0Lo
ICrsgufZeU2pEiywbEBMEEruKgVid7WbUWHmbzZqKnsCegRuYk183oWSb4/uqHCp4VpsQcvCXxn5
4HIQH+YCrZHKXwJ5ZSHSIXs6gmKLdqtGyl+pCQQfDOWoe5R99ANQhNGGIzr2s/UyHUKNw8NJ8KEQ
x6XXAV5S3vBJGC8lRjghn4nRnwwfWXfm02tEN1ymrhjka1eGKPOcGH0NMW+d8cGsxnNGVFUOwnho
lGhdA0fl+RJpBlUVYRSgGBXJlhwlFmOKykOEk7prt8wqk6M6PbpEtm8q1Lo80uuL2oMNW8iFPK+4
1nue8LwQ3/Sh1AyJnLuBKgm/hEY2qQY5499TcwF3EKh+EgEFQ76YYH7athGwp3hrRVcwMXAumtWY
VHWSgHD6Mhrw+utBl+aX9+uY3Zuf7ojI4Zd3IFUTLRP1H6Pymw7AtQMZ7kU70u43FhXRrAT1LR4U
ttZV/0u+bVXl6bZh2GNhR4d7IFQEvxSZQFMfURSUiB1peInBe01WScSVOvuVTFetN9n+sHn7ZzyF
+mEVY4EKtWJkbzxfkQU9Pqr0EoqrLoL7oQ4fx58WE6xVlB3DgnNOSg5QSVZpRE17rZS+Akbj7aYa
xfW9CRIHlxrZSoZdua8auDZRJwhLNy+oK/KFVFumclgEGNHjQW5Zq2q8v3tw1kK4RdYYFR3pwtRZ
lu460R6TAX4WSoZ4CTFmEoIHwcIodRyl3WHt84Irbdr5rcm9HDmyPv+6gYI/SjxZBmLe5jgr870k
08UZzvqI+AYELnNuRSm3khvrp4Vhc+onKZYwqS3HwAYWo5HDLGFQ0l3RQxZ72+1WUrjkQ/g69IB8
FszH9aWC4w8KRpUhzd8G2e6AEY8TuM0hhsRXgkdRs3XrrJYIsaEHM7/xd6RSJ6mlGgVvAsUULdJe
ArL05qY0cUdwB235m/0JEHMMhlIbJgi4QHxX8I7SSa205UOipKcQrym5INqgYCp9JUqj2NmFEdgZ
QfOv/jOXgzgIyC0yptDI25PxN485DNpqzZMTIOYJmvKJKK0gp4WQok7fC+jC35+o4X9wjt3ZLfsm
I+eMZt+y++X9rHag5rKu3oBoyQbZv+BRNbVBLtQcUNsQoUeIhs6TVchTTrTJzqDJfYmzhobmw996
S5usX2R9bP6Z84sOJWNzZrOsYO7m2p/9EixyXcBEaqb+m4/kEHFpNCZv1IMz6/iHsG0KARkU9AbB
xId2vra9YW7hmNB0uypCTj+JMS9IAZvQ+5qgroeFYz3IuqJ2VcDB5yXstVWpH8c70XmNe2FQ2loM
eAbZ1tEKHo7CegCk3gwfiEbgYIt+npjezpj7bHudLq1udiNZbFAtSEzPcelKAIfYG6fxe5VGwWvz
kgYzdFqsvKEW0CZHSmjXveaJcCgUckG+BYIpjMk3pmGcq20j7/ZC7DRsBR2Lhf/2gOzn5sPUgXDB
PzEYduZir2LAc+b+cWPdMuUk25MRgrmPJAvu7/9/6d9K7gxNVd7mL0/BD2fZnKnE6z9iSHLBj0wp
n7Iafuc0pb2/+Weghn9wsrcFVLeVv2wKAnG/8IEqhdYThBkVP6jZop5wUqa5XOFTWXGA6OKiyRZH
SfrXoQj0V5ux79gczBgDxY/WYhW3PRCxiyDgntKDTo11vIYHL8Yopeqg1+UkAj3rgzn97isDFLO1
+YKsWVEpXhxjHUE0rNIIwMQB6YFMMOVcXQeuteuxqsi4tjuBz9W7sOVcfXk0P/L8FMluynRnbQsD
8DSuJkiCPJbPt3xG3aQCDPMoABNkt5XJQU9hz9CX3QudFu55kud4zWv+9p4uW4CWcErHU+fBTVIE
SRNDQKmm95y/OlNWxC6VhL7eQVg9tobxxaxDgmfagz/wgGHBedNJLhq9LtPBs53LCTY3a3cFWLuP
mEkM/TIxp8sEpDkge8bHgzgEbLU+g+FjAZslNRrrI4+l6uOHudEY0cUHurXhDImGcr+NXlkLNlNT
RyKncVBMe/QjAjiQaYlsDk2avpWiN70ovepz5Wx64bDv0wNGVi/Uyoetgr8crVGxkz28WVeNfLNi
lLq1cE6mkecd6n4wsli2KzjUWIsR6Okc8AoB+a2c05SRdxnv20XWdQqiTA/7EmXjpBGk1vCeVKV5
SFeJgQwfz6hT928WRLIws7S3nieK6RHFa/BpV0sgd8mfLP7VI2YPucl+LPV24ROXgQ5hw8X/C+c6
sb/hBBaj50M7E/dYtuNTJv6osJe6hZSIHsIFsbUp2xCzoPp7FE2VWEyMCvecmkq5aj4HOJkS2fQz
VyrNdoDlHz8xAM3ZE+Fjw4WZd0gVyMeUNmKEnToE6V/EAmlEEyYSWNBZU/zw/f7J/4KYf8WWa7wg
le3RoFJKW7ixiohmh7mNOC7gyrhG6InRFj9wcZSrpTrCsQLbZ08eBLm0GqodsPwmMpUVZjKXKcit
Nd8Fsla94RZ/lh3UX+VXeP8JWkvyr524n4yFby04B7D/OP39YojtaAQywa85tq4W6iFMrw7Y7RRZ
ct9KPMYbLzyAYSEY1rE1u6uoyKQuFT6NKYSKBEj9C5ANr1KN9JIdLcFJoWlZ0xxCobwKdoeWzsu1
aTcKBMO+cp2JnMq4muYHI8b8iuPMnMmkenvJ0upWtDj+7b3Iz9g3JK6vog0opQqkEp73B0AuCkU8
pho3yqcb7KhCfHowMFuxzCMHJ0Q6pJ9Jf8fJtdHbHc0OE2O7uHZGeMIkppRxFeKjTZKTUWSR9Gqh
pP3FI8Up0s5YYJVIbGNFVK6ZRFWpdL+tP0h1BWHY0yRQjuS3+019EDMLJ9T25NBOaJf13dFT/dFN
/U9eKzqJznUWjWsfkpKMCUw/1lCjWrhoVYHl8so1HUSfVch/LK+emaO9BiaI5CblaH3N/hwZAaio
XgWJfEJAfmcUvk7rCuNytwFJpvNgGTqg++A2x4Nu4nc+oEil2jnPKCHEnJoXE82yYq0b0+okIWhb
b165iOwHTAiWI9ILtvI0yd5ur7HsGH6YwR/D8fM1iy8sisQuYGgw/DaQXf33vxyVfMO+Am43wS78
cwmZhctOpFqBxHpXFlbNWXNgZh93I8rU/Nc0azMaRTAHnqrtqaZ9LZksmK/nJT+1RMFAQTj8KukF
ORUgQuEZG4yDG3/1LnA1bx/8WPxwJFCVKJNn5mN8ohAKe6PNUxo86U3m8S3YK9LYMqPueK4UIDFL
ZpCGY7Q4QxMenJ2jd45dx71EWrZp5VaAm8uKMT67PYtAZDrcDzXf64MrIXzkvrjEMhcMVR5HiPu+
b8yJZlOm4bLtb6SE+1D7Skotq0y9e8Z04MayV15dZBDfYHcuuYIc6fEwKAp3ehdrRCu/Zhw6roMZ
+CSQSgxUmPBE+WYf1aqMdWn+lGQldb5rXniwFhZdpCBHN55yN77Aq0VJ9KwT+KEHNWaX8ooT4JEI
7btfqX5dV5/sj3GCUVeYJ3iiZx4n6La325dQvOY5rimjVeRXMBXSfhys3NOL1Y5w5K34M5MIkpZL
oXqVfEcczHxbWCd3nPGsdNgAWSRt14WeIBFSUAHCx2wNZcqTBM379eITzdUacFt6BCMEK1XkR4wV
2BArB2fLZdMxryARX+iweQsdumHx0pTrUR96LoZ9amvSFH4oY1saJ2QjrxW3AF3UlHTMQRYwOcRA
b+m3cksFHTKgD7BgbDwG3Rwbu0V1IkOeRmol37t4CWrnb89v23uYTglwIcUz0FZ+dEqtLpECppjy
wS5EF+VQZ9D3iAPVBvpHMQaghcfuZp9Pv6eK9khGbPG2Q0yljh8oKnmGse5ptzRbypBL0z8ZAr8P
zgmWB4Tn18MKclR5nA3bZY9eWVOm0eYVCBbYqH522f14wG2OOQoIUHaGUZ2kdypycyFqk5eHjHzZ
nOLP6risom5tT7kms4U01Y+57JYQxzy3AyDHF7c5nm/wVRbKcY7Je6I69+At6nsh4jck2CKiDzb+
FmcqJoIVaT4R/SBrryVRjOORo8SQkkXOWV86JLielc81L4HrtJmGBq7UJipE+jwGyWau9BmY477a
tY8XY9OALlD9TK4k8ii7DUHTsVpYPDZzoqwZEVmIw5ofdlEgsUV83e4AnU++WMKsYS4iAlf874xg
IOtSYZAh52LF370300pjJFtzx3Ir6NTuLsdNwJ+1Dzg68A4GeXDATVMxJprNU8cCDBROB6Ctq6DL
hLSrmrmq9rClDiAx2a2/GmoLJaNEGA0sW29ZM716i3Xv4EufpfdUWYr1Km95UpwDB+pf0SUxf+Mi
62GEwNrZuNiEIrFM9q/oWsfCfWCs4RcKSsjvtUTDdJ9GoffVqUFvtLgg2b5NgvXhQR77ZXPgPhcR
wrs/OjSN17G3oahh42OkkISmXGRwWpAEzd3e3DtJgCw+jYLwXA/5aeG6OkDWMDuJQQkCdshZM5IO
Lx+Jv72eL/ru1B+pI0Eplyg3g8iN6i0HUltI+diFPNgsP0jZMy2FAUIZAQOEtwUzI6ldledGxSbV
ROvwAU8dGRM0+ULnISW3PqzIVsuTDwjjDm9iiqFgEALX0GbwD7+Xm3o+7jwulDOxIwIZN6KqPSat
upDvYsoitBhqZATVAzZc2s7gSaxpVYmEfWk2jOP4rgPP0PE7K7NaC0hN5WdQj8oij43JtYcM1aNk
hXJyA6j3jmwwaHlTOa67jwCHelSRB9sXkEE46IlCTjgz4pH4nAe/q8MN4IEDWCMM9HVjY5IGYuaa
jfNyX9rYLeVqs2cCGLBihf3xN64cpxmGyD21wLztJDeKEUfbI4IQbiPhMz9KkhRnILEiO36IjyV6
gteiF9mmQ4cvFbwVNk2Hlw957Ejpr4PBnfe5f4gxyvcu8824dtqtENd21JZlTKQxI311jF5NUwO2
yqGq8sl0SI4JQySZB9c6qBWSn27PVuVShnYTxUwZkIEWvpQztaP5zm0nSDIXXMhVmCPeFQtBQaIZ
e1q0SqkjdP1iCv4QZSUXsZi4upsC+kk2qjklb4qWHSCGk3AdqQGNzNIlQAJRt4eoWN2ZaWGgCIdU
4vdziNn9T8ABFw+Delbze6ZwB+QEpt5TLfvcIRKlaHbny/aFx8Sa6X3V9isL+1mV4hTNSkDIZRJ6
ECqUZd9BIinqSjekcBAD59GB8k4vM5wxZCOzfRo1tOCa6WUZI2u2DK8g2aR2PWgbXZeHAT2eNXHW
YVcVVzmhP8a/o7z2W6QN/mJOmUpp4QftJ18SLFzdipV9f0NmDPEl0dsXHewNliriNNB3Jbu97USJ
3w/3kW2qi5Q9HWPiFECLfpl0kxr1lO97/96gLSIuziIBCr+dgiN8Tq5w4+GHxWcTGRTgfDaAPfau
qVO580FPja2lvgtldjpQmbOoqc7SOMJnB2qLkbLgVNmhtGnrKl7oW2q+xz/3KupGGfBORNDyOGc7
sIb09CqN6wBjuCjlyF9bT42Qexfflz2pC8DT2RV/CS4aJafMnOf5uTsVQulGq7wcxCFAH4DbajGR
HepVcMceDzOBvErrXm/Vs+TNkDKvoA9W8oqE+nhyxz7HY6awPC6RzJZwcxLjWLHEXPwnGfiUWzSD
h6iBhcd59wzUpIouiQWL0SXH5+CYnZQo7doql1uD6QUjPsSfn94EIMZLQEra9v0us0rRRhB/GhT9
5/lAvF+URac8En9eQVhuEqNuUFdwr4mi+d+ogUVNWwujaEIOsexG+yWWCIWmwcusl5BS1B9UapaR
ZTe8o5qzhpUqsVYB7GKYqYWQr7CLd04rTnTuDXk3Sszw0g7YUop4cmO7VdvcC5ADlY2kqZv6+GYd
8/oXhJZIN6JnDRJ5vZBBo2i4AKR07YD2xjDn3M2Mzmo6aJlot7+Cq1mK+gfoCWIcQnG3B1/2xyDY
zYPX7fUuGbSrRZGukCE+DND9SbdxnZimemlPMZq+ml9llAjqJeJZR6Wm9ANAaBjrAordJ7ZJhDy2
SSybPOQrnTD15ni4/j+OWsZ+PUF8osy5u/i7MTRu9hFwVuGm49bgeXn0A+/CeAAB2f23H3xLxGad
ox+Gszo+ihLG19SLfO2cYnOdBlYJW9ImbMTpMKGNyZfFZXTW3EwAl4v4lfRvh+3utyKErydNerlj
NVk+1T7c0kLvVrVU2+dbH/m1DCRPfOQm2IcaAFCdPIXhvFgTSZGuScxCunF5f5T7LidLaVmsmCkM
EIgvq/8jEIJRnKHLMeFrz/dP0J9wkIp5gHjUspSRCrHXgAekXyd+yFJcOF10ktrI71evtTMrOs/c
XSCsGGnBXKl0qK+69S1Kn60DviMrv5Lek66rImMWdpLrYASJWfiPtDblqCoAnDn8syFXW1snD2Jx
Wv2Gj7K1HpcI+y99csVZ2LPB5Xr68UIXb1jmSxnGhuGgSj83zQqF5oR3wwOJE6FX13MjKCzhzE0Y
LJpufKNiri/WZiqmDQHY+TiWquHtbM1WPUkh64AyRsC8ISe6GzGWAyvpLWcEBdx5xoQpodMgI1Pj
i7EaqgiZdVyXtIeS4fxBE5p8ZHeBljFWRxsApvL/6g1yTp86VRy00snqfji0eHydUmVevVKNJ7ng
UIWU4AqPGaGCbNaothN/hSK8nmxbL6pjD2VxLhyc3bp5V4GQFI1S9uGlMfUNkwZlJx5xs//HnE4R
aT4HuHdIDnDixeKHC4f95VLtQs7ZHNC4B0HHhPplUGtFJw3sPl21cnLZPHmjzBSUbYnS/2RFu466
KDLgyGbIK/L2H+JTTAx2sK1h6BS0oToGQk3b57IsTTMi+5GZVfE36qCXuECayQFrOOnqvviTRb1U
ZhqMHVQ/LKMH3prU3vw3r+RwJTgcvMP14exBRuMr4m/O/t7Awqr5y1hDyr5zviC54Ep9ARkOtxbX
Vr8Wt0D4O9uxhcGwZcIa7IAJLEY7o3L7cd+qwWVJUtuxaW1qYaGRDl3dSw0fVAVdFHt07+3qGsMW
ZaIDhD5eQ6bEqYixiC/YioD5QG9IbCLP7C5ele7Yekj+SPZ2MaNOyHNIxpv3mHYc8ruIZ5be8lsn
CO5ZRPsthP4H9m2ht0EiXhqz41ZhgPz0Qx7g7FOjNu8eDAcO5gnRJDOkZ8im4yVI043ZM8Ipv+f3
Q7pdfFqMefGKeNDiAalGi5cyN751nX/ZK3qM6uJsYZ56sT4F3y5SN0bU/h41fzau3BXMm6IGWOsE
GFA8PleR4AaNlNIvFen8G18b2UHnH48FtQLL8X/BP3+Zg+H1dfl9AKnT4kA2FOZ44nDXagxUyjjR
HBM1YiPafSDy8XVqEvZ/GXrnd1wIf82/zLXGWVBJUQJZPAyZAxWlXEj8l45PltLNlJo0EL2SJrDM
2VetwDgS+9smBHn93PppEnQ405UHv5aXY7iU+0MLVkCachR93dp6bdroZBRHYlGNnzUZDGIp/oUb
IHX4kJD5uZlIhafyMTjcxbWETxURXet3MUx93zVSIUtURC6eQWfokyaVwPDha3iyACvm04y8K1uK
RASIEhxLOL5WDWzk3W74cxXqhthP6v7E/BB3tL9VknCxKfgj71sJJg3YCSHHgrN5a/96OYH3pPFS
wEthl0fHDCXZQbc3+12o/5gNhg/xYUkw9yjNw9r4GGyYmWpzCNNcs3tTqamGWPQ54Mt7n5r0nE4t
opGL4GVy+vMVfvs9IkL+Lz7CUf/xpYIoauIuwaUoCcg/abvBNN5br2GpYxpk0VKG6dWhQduLvPKM
RkdybMr0tKf8ISqVupi+tL3rarnN6Wl0MvbU1qBTekFPY+6o5wXGC/Er/PBcmadH2NRvAIDu+Gsk
xaqZ4NNUdfZiRV87/II4OE4BoN70UACRHABK9uqxxG01M43Cf/S9ize5wRiy0m3lEXzKkq9QGJWF
9Wbk82tOPOpBcXUagxeuIRyUb4oAI52ybzdESvo5fRTXLaW8sB5/0uw5v5lmZ9Dz3WZYpdutlWki
vuJ5FF7eYDHqgG/L87MvKSQASfKDLzm7ByCFyJfqYJqhsVkCEEwDGa6k44cS3byKckuuBuCryvM2
vPv0f8DGBOgXupoCY52tVntWV0aOuKTrhUln0T03B8BZsPntPB6WDkZxO/DiAkdfFyCdMt2Ake9f
hBcVP7pLiWeRymqiFhMelwU3TAolbW8OBYJ69hSEM9uvTUebj6PkfueZQDR+3uXADxrNoFwXkwig
XqcwDNnlNznICESC73QuJPb7wNYozvS/x7DmFdnA/03+SxtHoIX1S9jt5sVIBxc5iDz7RrFbIeBO
WKn6cvu2r+QfH1qippvDQWM9v3aMxlVH62UE22SPQnBUcgGZTEiOt9lA8iTa+vw/QKDphs81nhzd
ObyBxiWyQeo3OjyJaX7NtyOHq6SZGRm9ONXOiOkY6ADsi7WzA8O6XMomgSPJBy3C0HFYfIwDm4nG
v4rwKCUXv52cwmcPozrO8cqZMHKh/Tkgzsbm4SFOdqjmz1PCtHpmtxoIx7e8BFoOSKhPTFcpWBS9
1p/dT9tF616S9Sb2I1Y4vrIDECWDif/y3RLtMQUuPOoDscljwMnhEpacNkdLb+nvyYi2APSkiL5Q
Gk3RuMiMXi+oBz+llOcjqI8K+4s7w+Sm94h5xkIHlNT6AXyIQjkk0MJg1u1FBx+rZ+jYqqVF+073
fPUD4ei0xgbwFuMvnGPRS4068c55UxoWCX8AskXrp12b6IiMGIHe3BL2c+n9yKN6XFSlgNLgV1ko
tWOw/IaaEBauX01MOHuA53nMzE59eK/UK2goXprruPL75GWQSgXSaqVb57tAW9QkSvhJvjD3cpb7
0+1xobf4dmxlQU+Ki1DHyhcKbkvwSzItQfEKisj/o+Ydinx34orEJQkw0pJNMjPXEGDp85kNdoIU
KhsozezZOZYP9a4tV4KvFa2kfojoZ40sfDAwOyXDI+eQiL9hjT8BJ5bEY44uLCHItB3JLIOhW8O6
RydKd9JBL127K1V4gD5qiSe3SVPusMKdiJJ/EWrO8ZMhLO89AVXn3QnwMS73GAjWVlvpUj2ecrbx
RBUhTOpWjVkN2O2N5YT2Fx4rBSP2YCecn6qBuT6cJwtvojsySwpQWXIfNVxKRwRg0GaEdg0woj/r
nDKwW78GjNOOdKl6QSMuPC4L6JGFWPmVPBjRxbWWv7oYBkymQ0Jchpf+JMZMrmMz0l31lubRwHEi
TGgTUSvaFC5Zm0VxWp51FFdCYZIEhkeuvD5C50Z/mC+pyVEiU7HteTRu2ITKhcW0aCuLheSLjEGN
VVXJxlHhze3+AtZKA1nR86g92wkOP25VFxPFxCnGx27J6t1o/ITMc9vsHNmrJcR2deEgG8qGg9n1
8tjbIoOJqHQNb8trDL8LTuTubc/4EA7fpWU7nBa3WySwf5AO/eoPi1jMTVvc4AkDueYFsOpW33L7
H4OX6kty+S2UDOHdGKHZgrL+0983T3h5n7MT4Ub8z93+NmgqHdp+egtWqC0fBJbkMiARhkSXp5lk
OElage0ucqmmSI6A6BgSv3nkoTPYiQTq/Qt7+GIQLHkpVWmRqqpCzU6O122QaOsmIr9Vksfz1Ic0
iILZx/7e1f+ArtaY65UZCNm8EhhWcPoefg87A9QT2q+tKBkA6zUPR71re6WYq1rxOpwyh5rBvqbA
/mSAaVoJLOorzmu/5euwA2LGYMOvxxN8uhkm+Nazp6u7DUz5NY6CiggWnkpcJICcF32u6tGV+1V0
vf48tn8Ij0lQ4y/A0eKRT0sMPvWWSYNxGrQGDUH5ginlBIV8hL2SzElg75CGfusu91YpXLIAfVov
AxOUawXeozQnw1+6JVGs+wyKW+EDJSY2oEQM4kznX0Eqq+vHKvFVXY8j5f4FM4GPEga8jmNse8Qe
d0uVQhK/LgwxyJDhdNAZaz+94VBPALwflSgb2hfHREeCXSnJWgPZex5UjeIrBkDxh8qzl3rAPUU2
dWjUHSI9mKHNXbKaeHBuGsnY7qajiOq1gH51wagWcae/1tPrc839BOh/sWUVXxavmrOMcK3lyNLL
fPiJUxKaHo5nD/v/OB60agOcmsrF7tLWSWx4UVkxkSxcQbvP3bjFy1ehtF/LPJkb2RJ+02twDxV/
Hg25m3cf/LVeD/RnCOlXtyTpIwB1Ax6pz/wZLnWWgmpRzwAG9w86srvOmsbG2X67mCr05Y5vzhDx
dqkBCC8jGTQDCr/SeViorAL/nsotjBmu+qVx+s6mWj7NjvqdEgy2SCCeu3MpuXJuPv8kAJ+CBpG9
okZjYnO9Z00CeZNDoaOoPCu4od8BKR0G4R1lGN3G4rtawAR3IsOY7Ruf5rnzP5Jbj7UxwipP5EXF
nHwSAj5GlB816BX6j01jOHYY3sYd79OHNMw7vsjjgqKttdaaxOZ87MJM+Ya7Y/EMo7V82xENWcwG
yQnsUaltob3gcIkm82hB40dWPtOtHFyRL9cbM/1pBPZmU8kKL0ahsHw64kF4HzUaO/DeGGQL+B5P
WtMNcpOuNIW7KEbTlNISLoOFnsln/0mpSsptYdsEdHDxQmEdGfJ6wb+xzCHQrPfV8YfZwSOB0RNv
gPYMogalC4EDrPXl+TF5ITCVdgK0xZ6hCEkRMNRYUWulOiuVfN+02ap8S7Cv0/zlzmQ6DI6JF2iC
WNrbdpY18sWZjhnzJrHwPFM0XY57Tj3HxYZ4TgtdiDoP3FBMQDhtAtzT81Rul+vS/sQBt6h6JYWY
ev7UlyCQGQA5xmiWYH24hjoW9vyaEMhc1T9sqQ+oTtCGY8MquHeC9RkGT60NT2sqh6ceRg0QydOB
jJ1x82hMPTESXHspTyiB/FrBHC+oPdg2VIdWMBPudTnFnQGP2/Y88VXy/VebeCB6qflERb0nLFEf
7gongHugaSBhqIv3HjwWab42r52fkU2MwYYugX2T39ug0YF3k6zUr7l/jx19LSBKGXgB8TctJ6wR
3+WVMeg+4BO+oCOZ7453bFdT72kSf32MwcjNkBrWHXmgDwFYnVpFYPu172Dn0GbJJW5p92QAi5Rj
NSwZv/R/KFDqLBr0iRYlwVPPQcKydchmrsh+WZ3a++gtVVFUMxZ8mDp/5RaF8iqY9QeH8pWGj5jt
3T3if6g4WLg3zli8V8WcJ4Q15M5HbOepYul9GwSuUVV/jxgu3GxymN3SdcvSa9t2pGCjHL582P74
hZbKVKJT9j3lTf7Vbk5tQJuGC1DNjSIUtmlP21JbfW4e+H6jFHuiK2HTPPzcBKYBDjii+lUtDRLh
h/8huJ2Pkf8xtOfnaF6zYn1X+cQb2vz3rbUayMPli/wjRLYldAYRTbd0yFPB3J20sZaWT9bNgH5o
94sXoIS+bR4MZXNAccd7sDA8mgCGohxsOqrgIz5/womSJMKpWb5s4TW5UJAGzwsYDyiedfy3vCBH
3zNxwfID+dFxkLd+Rsw/cR87ndc6RKc+BodEC/0UU5sFWZ0C2HWXQmcSrILDQw7o+5r1iF8vFhJd
m2a6pfxv14RilNgB6FBePhwiG5BLh79YKksUchbb+Hpu8G460y0FeOaYdjOzAF4aXhxWu+gusQ9l
7cdnJUut00AgfB3iXhyhFtJIocqnnottp5Jr82IZaItz3pg0z7dUgq/wj0W4gADaPSkySAkXOanf
w/xz8P9N4my+U6xuXYY1L/gn1l5fOsTdAHU53awEIF+3agjAoTodgNp5FQnBo8WWOYu21ea+vXb2
sR0DTxGa+pxppkg4ExY/yI8IGh4YuW+07n+K0xuaonkm2O08sfHaEyFUNjXNYA0JnNP+Nn3a+epw
VsoqjSzxwgUSXqHHTyCepmkcetR6I506725D/WOmHvnX6LG8MVpe0/xcLwzuFow/onHGGzHkb1CZ
w0ccosnyPyJrfviyiEtSwjdfhjxsyptaJtXA9d01R5a56PQrykloz3IcVsFFmA082Nrvn9GZAOoX
fekzo4h/8+u1LwVBHNkL2bmHXf0pdtT0Y5pbk+J6qymUbRSUbS30+8WwtxGjvgUmZ0CznLwjp5im
emfjdG822oIkajoT9+ANoib4BoVfw/wwlbTfRnls3a0yOcf650X1rOrL7WQfPRe3XV6AVMF5uhoi
B4/XLfMdKLagsAZRzLIzjbIOi1vuhpVN1ujngC5qcCxd7Q4gipCUf64MRih9dXsPn7QJHE5yNgcX
ip3AsNmbS/S84yukh/aCPniPJdo4+mf6Ha1VOwVND50ks1UO5WBc8krujjZrMxkAzkiiMjpyMEvx
Dz7zyW/L7SmRfPeiQGKQDVlijIa4/+vuTM7W5IAwPPxyIcM3fdjFAAy/3C36CZM16S8mqfB1LGPj
hAEJ+3lY6FRyXWZCC85Z2aDs0fBCh7y7W/yp4wfRGwVHxTgY+fCOCE6R8l5B0hq5xYu1BBgtfESf
LFeDj9Nu1i21eL1sgySZvtZvdNUjLiFci8EigKtf2QPz/qmget2ceSHnnPaOrcwGPHY0DN1dPjfs
5jCZuQMvKsFwnOXqJvWEEn4sXn1nckoIsXFc5ziokActre6gXTa326PFZz0gx0MPJGJE2yvc9M71
PLyWv1BurHxjDg0kzJAzSDfx+pVdTgalVHHfjIjV92tbHMUoHkuUuc8mGFt024+QWHBZnEs+IxtF
O3nDXxDGyXgbzDwwOdqu5/Ago9fQil21WO3PExIJZ9GVU4TB3gseSfTJZ/g7x49zPGMPLf98Eemr
2FoHOxww2Q6bmGs7RfGpsRqmnrYiOKDHRzJVhjWeBgYmT6jbbBb2/dBhhhD7LYA7ORkubX+3VSYO
QtEm+0nAgLkE2VpslUdJYBxk7+q4Sa26Vj/Izq5cDAeAau6e05hbqMm6ztxv4MRyukuccy7YXF63
wQI3gORlsOlIVtxoTKnsGW1YIhZYefXkNmJfe6kAQ5c4PqPKGVuzz0KQ/o+ZkJFSXzURkDWi4oXo
mknFYuwh/L0Oo0qwFNp1wumx2sLvIH9ivSS//s8C48TfNBa8O/lpA+LIS1GzqBFWVV4Ldz6PuMLZ
Z1p92/dw1iRHJJYOdhhpzaFJjtcSWExEWZIGhbWwpcIH1r5lsFSAY9ARd3itj5V7qopG3/lxS5zL
7a4XG2RajQ5llQ1i0fg/tKDtVQF392NGkY94tQXcZkPwDHqV/gR21kNYss414CAYA7m767Z2eWz6
PwUeXwI9Fw5JdqLJVLRP2nudzGYmdugJZTr4cKiAzz/yH0QaDohCxDnlMDcclpAx8qngM0S6eN2a
FVJ6rX+EYUvJUV3yiHBD6OeOuX3cToLCB7EFhHAp0k10gG4vMgZ6r2B9VNPy5lJKbxvuJr+G7Tv2
Bnh9cczCL79ACi26RWLunwBYvg3XGISk5un1kjuCGb6R92FfMsWzjV91f49jGb8XJOiaaV0riuoq
6aC5nEc0XO5qjnC6qMzFw342IXctCba0C64m1ZBCMiixETuOkdYAuLp9fl2gWmoUfPLKEIEL75Tk
V+FQ1QUTrJgWi4ec9N2qY5vMqSmsp+23lsnFmj6oN0Rpgh0tZ/N8gKiPHsk9gKEdBpHrOAjsf8Yp
CjGbIldzt1f4YMXVJ1KOCq+vIHHojeE2gSSZOvn9R3/eyqkahlLIeEORH/6vv7A3PH3mEwj5km2H
PFTRz+8LaK8Gp9aEDQ7YKCV3uP8SOlYSpun9yq99wiUQdt0joV4Xky9mbqIgzASilkk6d2U/V37x
MSQkmwSrDecBKyD2Gq2kqeoR6YswiAOvdf+7+FK22SZ64rYVJ/sb3oNlSv5dcr8FPN6P0QxwkbI7
Mmo817F6Tsy18zqxTD6ouOpmK47M5c9O9+L5bnQOL1s4zKq/m3myHicBsgfIkM7Llkd084oZVrGc
XFsR56+Zm84Is1hEyqGQ6ibikFXaNDQn+XVr11c3Rr2uymqq5JkLoKhM/ZjETrX8uUt1qh8yvo47
yVRCEl+EH3UV+1T1ETwJqMu/2uEpGqGoZx2APm6K5xvc5g11u6qi1CP2dMI1/gU7jXorgw+cFoaC
oYdb1G74yWMnuO/nzz9je2DFQw1EQs7+dlLTln+YYBnDiMmBB+kg9O/PYcN1OQc+FPhLgjIfgZNd
dTTJ7P2XzmS5ZC3RncKSI96T3/EMWCPcWw61I6JfM/5WguxwuqT6RJfmKVE1dOcUX+LYKj/YE/FA
1apkIk9joRsZ5ZmRfyH8d4csKyGdr0k/3/b7wr2shQd0SrZihDbhk8lYUINm45l+j6h0i26EDlmU
tf+McRY85mv6toyx4xToz/3Ey8usuYuBhDDwI0ldLVnQGfND3YJyKuy2s+Eet26GL9DR9gdWZjUM
4UY7joT3S1bZRnRyIGG02wOGQq8Yck7dREo8Sq4K9XbnyR4Ad/97V1GH4tNnHwOZgB8UJam6CDRz
s49clxRUgUoObiVD+uZf/v/NHZc++ggeggEq8lxlYHQEdDOerTPEnpLKg6Oais6K1WF7CoPRlgPi
WTKfC7XpDBd3rxiD/Wq7kVMwIH0xX43XzNSitX8b1PV6sQNdN6ZPnjx+Cu43RO7Xgji+PjgILJV1
zqVGVgPP1VIapJlBMzehI/IsYcjIkI/DD6IfSI+GZkxJF9nUS4cB/6UPpct/aAqMaQCLp0dD6eqt
GvMdAE2To/Q7nKEeiIhSYOUnyZl5SkbjOoHykv6/7LesqhZGcp18WZS+SF2mBELS68nYW+Np3/2m
jrnP8yZn2jyHeOdspq78HdelTMzq45cJw9KsUQdfinnaO/5Tea71ay5U2rRtf+ftcIOLeK6xLQRL
bRaKv9KdL3KaSuKanws704J1G8FQJnRuC9YzaCwqlb4rnY8eeE1y4XhdIF7BqGMNwfsoSPaAN07k
zVpT93WLrg2lv8IOwDKERSSISkred/4qlh6lXevrRn0hVHHOpS861ffhhfL0C/sLVV/JwyTUrK1S
TQZR6bD73apq3dETJcNGK4JEWSsx7optfgWJIZLNyg0fhO3hZVyibOEK3rOMqNVLhH1HQ6GNRZKK
eEXBuiqyJTw4eq28P/VO2uQ3XG1njBUpVOeRui7sJibss0hxu5dPzyCD7VLOetMla3p3cJ+gkglS
GglHdc5/hsO7+mN4h7dyROcGjmqe0m33sUGLhoqs+1h0ql+3WbvWMC10NDB7yLU4gqiSWAJiqptA
VxpCn+PFSmHWxtMXe+K7HoLukIG8gUe4GYFd5KJPIoEUDVeFLOzLqHd3QVRmn+/HuHiAM6cXtS2n
Ds5pkVDu8wuotljsMXPqAA/eoFsU1wXA2A2Fhy68hS9LcjQ3MivVKhLv/tF+5ct2h66uILc94ZW/
6CP1NAutKLzShr+G2NNFSELES0O79kZilE3qoRYrnqJ3xFsa60Z3bouM+3bGoXjVhnABOcnDCYxT
n9RuVHZzURYGuhaoAZV6tfUvV1Q/X+rfY1PR5pr7DHtgsMdIU+7EzLbhXD79ZsbcwHPiT3wDkdSj
FFBNQDL49B+Hk1LQc7qTnc5XoeI/A2WIidulv2lzoQ+AmYv+nQI4d2unfu5DVrLoXFQmnjA2IFFA
0sfvtUXDNXHkV6h24s79TDugGWKveauIY6o7FLF/3BnqYW1UMriUps45sxxwrsmXFYjCSKuLV5Fm
YDzXMSqJAwduPYB+RLOFdO+pH/kXthkDejxkP0hYcQWXyjtbLWBuRxAerFq02jGG4qNa/N0uudWO
pcJaCQWL3OtN3fQZ8vk7EuGDdTJRyAXWFNo2MDN4javcvZTnGYbuTdfi2CdtbQZAQykEwC0+S6//
4zaj2JUISCAarxoqgua0D8lQW5Ftin7Cz/Ljcu3KfJxpkQAOinh/2QswPHVS5tlgHH47K4S++jr3
M9mQ8Uwdm3xM1VFXrEQWvXsoqrr5bL9dCGG6i0w0TDeHKRPJqXIRhjmXXYH4eQHN5K4hT21eEuRH
58gU6MbImN18D/xGxpcI3DP3j+OSmYfoHsuU9xTl/pF4JUjEGMC4roz+iATrbjvEIl6/7/c4YpBL
BcrlQKzrb4sp8LRvq8tvCztoSJuZK9UrJXQ0Phkpbfyr9D7XVPcTxJciBktqS67l/0gVtfRojWCt
QhFJp62r19vvO2kw2+qHbr1kLbAUzjx2Gr2AYwE4c3kEw35Myd48jO4YQg4PrnyHE78wjZ4xggwz
crqpOxj4U9b9sgsFuHB/oBrTEKzjpIZWFLLXMV8NJNTA1jJpPC6e3CEBRwXIAFDgXy+qSVPLdjPF
CoTAoS+v/O2HcgwsMKx212kWxRQRIiLu+33QkkEfrsckqBVBrKViHMEaB7U1bkxhysP5M4YyOk1O
OVbzu3ow6qDSr7hcEI70Oatr+yEIdzR0pjb4t5n9IM2Yt4Z9TGw7Bd2j6jAUvQ0DRVdtCibsly6g
OZkG5iUaGe11M2Y2VaE0W+9JsQsm8RmAZh3eyX/zOpNawPurpiQRDtgYs3j5EbET/DA8StREwABv
vQq20qI9sifzcgOMcWEG+XQVgzRQOzKPRoy/Oj3oM8jbi7oi2R5nZI/bBpnEWfltqYTg2kznpzrd
TNrjW+6MNQWkrGsOV/ByXXH7EO0lvcNG7ENKvq9+/PCuGKKVdfeS6HGKl7vFqL/zbQacWc1SFVLt
cNtIAx1bpPnzIJUkj0J9lLaGb90P4k1GdFb3qrINPWxYA8FF1g66nyibvmpOnlYVabv8hZH382E+
r+70DloyINTrx9QR4HwmaqRyN66rKqtzaeZhhIzmc7pyLe/lkVm/kprJpRsWd3SF9bLd+5Rgp/yX
cn1KSwOwrG07w2pEQkcEX5meIcqJQQy9PYVxSLhdPJ8U7MfxwuKbIQ+HlGAmRvCyUwqDWbrpAPbl
rHr06YI4JJk5ciJo05v84AfFNsV3X8sfquUVKWPlzoud0gukatXalarLYwXBAx+SMbaZkAM5mT37
SsM7C0Ab6q4zflrVk5mCO8WaUnJ1BfMUDpg74Swky+/gmJppvtKmFeXxLMn2G1fy9oomOy1iAo5R
0znFU8ZcPOVAskb8mc4Etr5rwiCGCA8fpZ/ATR0bt/PQ9weLzrzvktxEMxepIHS6zm5EnWZff7OL
O4OiXVhG7e08j3ei/iFerwcR9JalIZ/UDNZgoIO28EoJzTTZNdFPOCE0GziuBS+7jc46CqetOrZl
GKKelZ8T14kxI793cJbNZDT0Lfx3EPBsPFn9R5vVQG/jJsRunNDfZrlgSS2gJxWjJDQv13Bubro9
5N++5E+BRUP/tSmAgtk7usKlOVffZvH3CxQcuqRQ/zE2oFmpLnXiAhH8+Jlwd7bUQqXQUHXJvHKO
KoBk5YRwEiUnLBkaLGe6QF7NROlG1pC9BBjV6ijnOC4ZdaVaEwmrBQH2392k6PZtuCQVaH6aMJC1
glVxyvtGouOjOUZNuzCRaxc034hswwG1isAaKZAo+TYGUgB3NtfXaCGLbOR6s89x9LJ2jlWg6UkV
E0nbT86CV8ZrLYzbNTSuQ0ckALyCPvBJKrQV1GBhtG0kQ+0TI6/JsQk6/qxRSjw43bKvmLGb0HBE
c6FfDiGEAvh8UkJGbvfyJb9lJ6e/AAXDcdl7bF3v3TCWDplZR0D8kA9EQ11myg4m5oCzQzgYwrz6
IvcTzlpVojRzkY8mcZry54txyzLuqZNzsH/ziAFwI2cb2p8AAfijVYo1XV6YOZHG8mJK6ZFzyPrZ
GAq73XEYqUCoe93TSDEbDrxfHSp8t2NNeqg/vq97RLsWA3eUGDdIr3op+lO2B+W/afHhuddtFdPp
S88Czw0Gi3msVmeEqoPCsP0OwcmtnwCXr3jEM3nfuBSg+ilAtrJ9m8M4o1Q4O2BmKnLoKU6nR1KM
Pp68AM7oMJQ9OJKaYEOxnQCuD6orozxHXm8X4gGbKAtH1+pP24Ln0RoXnnY47bPZCbT8EAKqoo8q
rk9IsKtD9BOa61nG0yWmCRhfJTW19NwLCnl3beEwp9L9uPZJ2DJoUdCH2DsYSm4Sude9oyOVuXs3
nWxGBR4y+RIdsyAJT8mvbG3GT3zmo+Wp3vwAu3Qly/30vKxijaaISdCIi+vEz0ZHLQKtw8lEOyfO
FtwMWeYCYqk4ZPR9JCSymIf/qY7H+X6lGkQBzZoWOa9f17xRwzvPLopdsLBVm71LiaH6eYu5xcw5
dffcpm/HtA7WYh390Ay+36pac7/Ad+dk5CVJ7OZEgM9voWCSlhtX4O98K1kVVtAgY4uSPo9J0+d0
dzhcWZIPphf6B2AGAy1Qg0wBw3O/gYwnaIMcC+Xh47jRTTPcf8pJa+yB1sIWhFTTi20mW3nBDu+k
8VQcUoShCn16jm29uCQog+oizO8lfrc8q1HQOePZgH1kLWmKbfyOeg3zk0lYbFOm87RuDbnFvLpb
JZ78ppePpPrmOGaogDzvZgW6Qp3EiRok/7D/ekwuDCezYu8Jjd2jvFFFqG1FPPPxrl9f9u0F/LWt
ILswQvhBY2UZ3OmgLyZnflrqtCJi/31BqulALTrkhcbyVSpltFUQcdVtDKoDEqmaEnoIhzSstALC
2sDSuqg9RrGjrgyC0Vph9B7EhU/xTtUD0pEke7nk79+fFlXiCcaSWawJRKzfGq1H2Q9MD9mU5Ejz
7ktR4vLfd5HdoJGVd1jWKjbTWTVm+iKg1kx9tW2bG8RmpB+lXLaYfXyF51gJoEXWcUj+NsWMeV/V
YDDZqoaR2KhcbS+JYTcIg+8M5YXlzOm95Kw2rZDsGGNRpr6XPcuTp/Nk0OKiCcjZqbHdnROtlB9F
suGKPyuXoE3Dqb2BCpD3kzbOroDpUMTxtGKe5+n9EA53GC6+929iMuDdIMIvmajWMUeK8bjJH3Zn
QCk2xI9AmLISy4wNZOJ0ei+owgsdLF1ajFkgo5aJmyCTEctgYDrowsolL+hLjJEoGFEQHcqGFP/l
eyRa8A2p1cx4GRO94SVkRw+Hk+3cio3n+Lnm+lY4MwVfGhLuzXFwbb/6rUh4jXHHGTNR1xcMG4tm
/UHw/Alz6sStlhPd0h50ZtZT4v1tJknbgMRNLEDdy3EIlPEJ3rY7geovE4/f66YYoj6RqKSo4ATb
i/bupJpxwlknvGyR2rFJh7K8+Iygz2KX9Pl1CdxQU+3IIF37YVjRSdwrtZJ34BsdnKY9Fhfoyxpz
ZE16Rpwpv0FB5pa9/o2Mb4524c7QW698U10vH5kyBPv8+/BxONYLMUh5aQZy8ZQWs6m1IM6ajkHA
/N+SGZX80WcL07+zjF5bCZ/yYPIdGpb4VDjqAErNOCEzuzITgPGTFb5d83pd1XkYrS3KiEGEK2PM
hP95YGAzbw7VIeeBETCdDGJ5HpVxymDdKaq8m1JwnE3a2QWFdisHFK/ZSrYqc3bpK2NqZidbcMCe
OXaf/86hzYlXL8V0WNOPyS29mNXUGk2toc5sc3uofGODYv1NMunS12uetuhmttTJCuZGe+9m2G4i
esw7ksvthVi4rbun+oAs8hcBqT5XHE22U9yPuN7MelUAqOecAEp0ZalsT2A6giR4Fn52d0G5fE/9
HfjJkUfz2uINo3yRG/SfKezgPxU5nauZzsHC5NPa7YKLpWLcnT9kVNeuM8dlCTeQD4U0nrsJ0b6q
DNVbNvMpT88pRFGZcZg8y+ZDaDYFOF9Oq/3zi4NSFpjPsGZaj8z/xhqeqhZVnkWxXatNS/u3fxBT
suuEmzDwVdzPXXeiRGgqLNBGwkeEAyPvyRdIr7IMc9bqx8xJOALFvGWA6WK0j+iPm7xpxC2x6boU
+DM1lys43Bsv59zIwZmyMyjSEfxAjuKkivNQfqk6DueUojmSUX/BVeKNaFrbSkKzJrV6U/czMkRo
MAT+sJg0iowyN0vKQ8YG87MPRmqcw7RePz8ZMaFjj0qqBhxsZZDRjAmqpexf9nRtY04a7AuL9qbD
0hYxa+JeY/OwNNmFz4RVkOynbKfNaRKQ9PBwp3CgcbVgQpN+kZKrRTXiRyBL4s+++khkpuKOxCtk
U9+72hokpiDXxm8aTQKQoU3i5uQeX0Sb3uvlN2Q1Hn6boZLEKDvu7jUvlDLEqeK6DDTsHt09ZG7B
kmE2xLinhNA59W8f48yafLG++pHILQYUwvhxlctWrIGYabX9gypvxI9UpD/uSDDVdffCk7vUuWP9
GM0Od6FOfbu0dK7dbceGMYW72CGXZO/+F8oMhCUlQoA4wBeigH59V58fZVWJubkDssKd5HfWR0WZ
/y2EvtZgJ2ALAnRsEO3k29DCL1CveKX9Kk4hQldFnFy0QuQ/3bkp542Dz5cFVwvLeM3p+tEt6csj
+8qBPkBCymbY37Y6CObkd0xHD8Bg42AvB0syShJbVJXUgCoIbEKDUsZX6LWPu6ts+sZvHT8Y3X67
zMwtsabnP59wln+/dsxkNGTHNycftZT6O+F593z57HQtR+oE5IUEZJWrcMiQpj7buNp18+/TMxeU
T/tN0mRhri2QExtJaX3CtZ1Kwgqr3LP3jS6AM5Jbq3gY98UgGwz0BwNgkKTLNIFxWI3ki3T9vc3i
1VtnkKfCNhFPw/xxmUxDIzJzNPEc3TKjr/6JxpuaW5KrIfaRrYOJsTwMxugahynrOpVQdtfuxRCW
UuHGSeUgCJflVcbLkUrDDOQp1Y/9qhefs/RZCJqayz5qSiURDszHViPgN/AtwejAceBmifMhTGvI
ZuUMQVZYMkbewuY+XoIolx1T79elHb32tkbgRnX546Ne18mMy5OQx8KOBTsh6qjZk+O+M7OQRW+F
l9RSHN4JUPuyfHKXA6KCtpHJ
`protect end_protected

