

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
esuuckrrKLBFMMgSrVud2ZnB0pvEqrOMx6GkXz4dnPp4yshTD6+Y2glVVVlxat4oj6oLNAI0JrQK
DY/z82hivg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d/1Syr0Yfz0kK4aSXCIN7lq+kUu10RASco8trwm0ImfJURxtGkX5KSPC9Owus8m9ZNLVa+4W1mNi
DPA1z5v28araMT+WQkx+2smTTBb95QnM1r7IY8WLJwhz/4br130YtPfh6ALhwuPZLGS7lh5+ZNqa
WUkp+2aPy+o7nP5Neek=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EghETPBi398ucn66loN/344Jtlwrx7OhFAMdZLO3Gvsf81gd+y/lO92JbZIwpE5sZICUxsNH54dw
q7y/XtZVcW81UXDzCet7Fnd81N7WGIqo0pJecDfSTWB8jEEqdLB/p9QS5cVBozkWw9ZXd157NWH2
fYI6wtb4DiMK+3xbswRz9tjt4QpCCW6pl02xp3h0AjoDyHQfQiHlsbTSjlklPmKa/t4Bvl+J2OsC
lbC5D/MuvEAoTUQ7SK30lNJDTITWXb0RGcdN8tf/1AbxeMFGNs+DvhkJcoBe11Q4yCS9vXGZYmJD
ooCuGIJ149GuhA9Ebc3S+zqtQIqgB+Ip/rSAVg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XB7G1kS71wIOs+JCFd2Cvu1TIPgCW+AVgVRokt3aIVEjyzOaNQpUv0JxfFRbYs7j+wNszYGSy/VO
ucUpEKb3V/Eh6Je+1SiQK8VPkEGyi6kMKodRtbbO1t51Edv2l3Df96scmfDCuwUmCLxAYCnMI34o
GJA4Te4oMZLzNzksU0M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mYbz74Wd6t4yNkXqEEqIyqTMYr1gDkxJuJW5Rg5GXWUomZKn1t4qMArQDnPwJx4y9XZOu6/MtCnL
fPfEaeJGNkk3xubUfcA48NrBjUlfoqpqaC5sVaDR10h1kTeB38B7pV1iwRz53qngpcQ/++tRqM1Q
t9nxWednDhGT13iznArEKq20RLCcpL20e+RRoIbTe3wwmYnDWI+ysKyhOx1k2FPgh9jb+4RZZgn7
7PDivXP/gbNxEf8PXBmODTX7OG6mMJYh9DN9gjuP32wcsw58ZKTKhK7ryO26lHYq65/5CZ6bVTRf
+77RaLVhpZ+Bo23bR+0rH2ulVAt4vAhPt51hRA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26704)
`protect data_block
7FY0nOhRGAcdWC11HHcHCgXWGu+5GKQpSAV1Owo3eSkisWfvQWfEHhXnJKKitdbaxt0God/Dtn/2
bPaPpnnBEjYtiPK4zeK4j87/qFHHOic3b407A7tZKC2BASMWTomMsJNCWSYPu08hQ+t/RYGX5f37
aUvUjGbF+gWuA/C5YfK8oGHhHJS+IDwg9FstZuZcZDRwnhh8eTPAyGTeiNvKaLdBqrUapHcKxlOg
Or1/3JlvYnzmmnjHvpmuXmqio1sa/EIvrNuhCyYSLKnyNfbpzem7zgmd565W/0pLeM8mglsOoYch
TIgXw1qUww53yTZvBAcBdAylsQMgyCS5kG0TN3kYE5VrA++YQO8xm2Li+/HoqpYXMtU8CgnQzPU+
4+BJVUyWbjoitSgCFK3lhTou3PkWYFspNHHOWB1LSoMvhFabrJehmepqIMTtKgfy2YIbobbdyBEo
DIZWAFDN1gTdeElMJJZ0jermH8AKaqpxzPXyTXOKEpd4qc5zbS9ykyi3FnWYkzj1P9ZmtyT0+M8Y
+z2QbfWKfSG4wxZrG1UKzWDsQbcMe98zrF8imnAcXDgbyx4Gcxlej/W0BsxfzuxrEFejQaT9THEM
8PpzOx5ca3r2CBg3fcQAJfxMMlR78PaapS1aV5ZnzmPnuHcYF8ZACINW9sbQCHs6c95ZyNM6WF57
00hxDNYLP6iOTQoOjQgxzbQM1iNRfmiGL24rSGkL8g5SsrUNmmwZWtFlq7M2/so/MIwoXokgmfhW
yH/Poobs/MBXv4X55iT/vsSxoQzA4YabbvGRUx+f1JjXqLER/v0x2rftOrrqxrJJ2RK9uTSPPa0v
F11jmybArgCKa4ms1871QzfiKC2YTSe5EFrU0e0lx/qwS0G5VH0Sqsxj5STyfYiOQ+K8ONYdhVnd
3Tz1HwmazrPHg8TMt6AQcaOYN3TONN/noqo4faCwYpj3lrLdLi9uufKGmjeP8rAl7YBrZJaTQ4wz
W0BAA5CxXlOjoDNctkzVst4iPwNeL0JMGkQoWaK0Y3hx2V0lUdiVHXKHq5WCSevmh0ntMCiS32bk
NGw1Z4dAF80w+EDkTphlWPOact2DxrFQfl+p9pHcVEJIfpLAtdcVyCuiX/y+UWzqm0Eyk1Qkl4wO
GN8VyiKXG3Y98efdvc5sQlAk3367QvgEhmSMy0/zVmCZ5gbrlYf7UNb8WOtPQ8xiENPvxeZMqD/P
CiukLc8wtltz6LbIpzawEtrUorAs/fKIeVtZVb3cSdLhF6JxPgRg1jQo5mUgdzpy1ATieowmOlK2
GaAetbP4ddKAirZDpMZUB/Kza3wO4Df5ABg5LOZEEfyhMlJg067kbytgE1RfyFu+lgJbImWHPesd
nFtKJpiAHxCtcSBhRkA9zyXGMl2Bv56Ju/OHKREjuasWCeI30+A4rf7Uf6p77NDCdOESod3A9nn0
DPqbG61BR3ffTEil3aguNIY+Ui5Bs/KnAg/lNLt5cMtjy3iekm1rKKZOx4cyBN5iN+YxIhmjrn35
gte7lcjLBVrMH0/Wc0i4yvpfj04Was6wlraiu9iOCv+mq42HL9cobUgC4bEUyM7NnfkC1oL4y+4x
yIkD0IAUUpiv7iI8QUQklE9Nqzz4FZad4iutu56evPESHGS2MaHoWeZRKCNWvC9HH2V8LM2BBvjJ
McDJ/Q689hCQ/2xWDRaUEUGQac7JAAgZBCrg3SYtulczRmsOwG3NHJTwQFhSVfQpRh2bVmwL1kYQ
BsGA8mRK4otdxo59adeAZvcKMiDDgX92jOanKiT0S2aGmbHfq1KzFbczpugkuwp8r9mICbP61ayk
8fnl4fW10kN7LdSgm1IPshGQHMFM1nfZ5GouoUm71LZ91nRq/CXp1yxo46qpD6467jSPDxHv3tjt
vooq+V98loW8732zSQLfRY6YUyqB/Y3oKYQ/7Urq3BeG40RXd5xkVcEDyCkhtyG/O7HfbIpu/n/F
sLHgJX7Egoofhf2Fw3IoPp/IRjVh7CtGeOBsZKB7OPfO8N4w7PkZYlpXBgTc0FTXpCvHwNP1x+dC
0rq6+0bB6HViuiODqUW6MG3MNKlXLqJXKNqsverVVuQEZMBlwqrlEFTRC5Gkwh0GK9KEV8xnkVVK
0FEhpmY3ZxICqJQM7Hmi680AjBYERGd4nsvtwMz4l7s07eH5X/wciB6JL0U6UGeR65HCzvraf3js
Z/hJmOJroYPgjRs81CEDAmX6o2nQQn1yrQPpi6I0rQubqRWPyOtmqd2T9iBo8M7LEuD2qctH0WDi
QIBcFl7T34vbxM/ZqS1GkDMUuiUhOmk0OK+gisVpgOCH6sD52EUYnMU7os0VWpac8l8RtESjAaru
MqjW26mi/L1nZ+i7aJucR5r3S406ATiuUm35YkeeyReKtE4DzwLglACl8mfBtDJH+5BiriuFfquF
ULXvAaVrNRskYKrYvLR0Suvx49t/eLryVM8nG2H+YxODd8LiWdGZRRBok5VFjX6nBCzGhLzc0X0v
z6F9TnecxcRz55MZp2uNQXsjh0AIED+V0tk7avNZL4J9VHqhAdbXxQklUpkkOVJOK+aHTdX5HWLy
OvXGn6NW//IeF+hxqvjup8kP74dI5OpWycpdxcJVyzmOnvQTLcc66l8BshbdhbCa3K/ZaUr405PY
+VUug6Ji73eT8mJKQ525b+27apTCCdbCoF10uJNe4pkw3L+abADLCBP/3iL7xyABh2U8YYNGHYVR
B0imz4Fy8BbK8V3E8XyYshKSjt3iqPXnt8CidPKGQ2bXst5mBdDFKTnmkNWWeDDEWo5h5MSo5S/F
N7bZ2X03GNNRcGFK2dsc5PXce15lD+ZWEjfFbxmxGxp0HMna4+L98YoVqs51tlj4qEWvEApgjV8b
cNrStkkqitI/p8ptzp8WJfyheTIXWZfmZhnFTVhc0agQFO1B9iuk1FzJqv9pmExj6eP588p5Gjb0
E717XwU+0FteHUPQp6umkjIQqFP+tJPNqRCgwOKI/jY8o5ThDZHeKRBpIaVcWBgcgUpjSZ8hHe0p
2hQkWvO/tPhdyy1Y1QLicCsC5t78uXQ4tpkHviSIa2hIZb/YqxKcAQVoGlzQ5ZMxLTOULPCR1ImQ
fBAKEQMWTCqAaP8FaU9g/BgFBSIb6WYNcpN96U4CeVi835IlFnA5sHzeNF8tEgu69gIzFBMmAVFj
gD8bEuiGK67G1y6vD1QebPVy0SYqowApsNBhJ2vfKbZM8S/NmQ8E5koq1RokaS46G9vXWv/sLyo4
eMkVyUOtVc/qYGCtoSmqw3casPoRNlaQkx/rPQ+i3JH5n9Dmv3qGQBo7kWVAlylnXP4/j5Yb48sM
HoK34XOylm5oawVCuDLEaLNH0kae48jaBI7VUXFwCAC5rqzyjvI/fiNLtcAlWv4A+AN9UBLVbwWy
AyurIBfAn2Z9hkk6QaRfFH5rKfJNO4g8S2wL/rYjRef41uU0yEZc04me77a7VN5qXFGkQ8EoWAgF
x0WwTJkV5ubLxWu5vmlDhY/vQB7M6o0XxqYygnlzRoUcjyM5+o6yBnwWoFjaAHfFJfMvz6jaxNUD
kzk/M2P6jdFUC0D/AyCZi1xqpw1NHuwD+AF7CdamTNsWLjbwhUYSQo5bFIvYnE0EjhpSkW4c3Q9f
nLDBGegD+6QtWun5dEgH71386tQfbE9phgYWL37jlKbckGmUdVSF2PC0QuIzMTDEiEjtLGjZvFAN
NhihwtqfxzV+Xup9uh1+y8YtQBFp4+AZx6CWLHkQ+Rr059STdcWS7ObLisZTfAvQ7pteTRuQ8JpR
nft1IOpo+jCbYz7Lzvz3iTXiUDIV6lMC50SXavV4X4a2ukQ8is56U1pEnYiXw04GBmhy7R1VAo5I
aNu3i5kINJIIUmIsa5qYLXXI/QNJnhrfvQwpbwudnq2e55OgLa2dSNZv1mg/UYopPzXOOVzMPA/R
z8Mw2sTWwbNEN7QNoohfcVCJU72+vROIKBjXlInfUYjaj7i1TJSqE/pPy2ihljvnR9yZtYD8sp8Z
9wNxfstS+p+26xEsNo0oZV8i4+RDG/MXPEDTbY4FyV4ypsIK2C2TYDwsZjZwO27Ckmwx0gM9p5oZ
z3cS/ZOWXs6If9eTL5G/GynUCKCItlbLyAgXxAGaaIA8BeZLglAhsovOiIl2glBGFLJjCsG5zW6J
GKWRR7yKzqbqYtlPSjj3986fk8q7PORuDZCZXWsPvocx7Hy9m08Y2POtmimDePKmxIN8asTup6fi
RxjEIU0vS1zJ99pSPQ7H2vugsqDRLaM9792XjPGXptokYdTBBrXCLCUDnKSN0W2I+8fxOhd3boF1
Bdd9VEd/isaS4JLPfck9uuchCVKQpYYpmhCfO8LuQBD4reGNazSMdskXehmE6R3LZX9gfqibbDzf
OOKlr10XTJdugCbZkqeNwYPB6m9A6Zs+NPyNyl1umoqM3h5hXUjQbnAPB4yc3o8OHZUBLA2ePRp7
y3Tm2FS1KBmkHX5kdaFUnnZ26FJICAnCt6H87V6v7ucKCRbEm7GUk0B587EK8fiVkOJJKgoJDwKW
hNtdesqdiPvdHppgOC2i1e+GHpsRM7B8HpjjKwV6Epj758O4eT9nUl7DFUT1ApNepirM2vH+BXBX
OBMRjm3bDRYz6ETpz0oM4hxvqnnrI3WTgGXhXQwhgw/8MRieVCLkeAYcYYheSRJFCYWt008HNZwY
K85Om1AinjNlQ937DJvuebcHcFg1gpSYFu5y5+3QSpqc5ypzSwNaRF/ZAZi948LzV2VztTWmsqV9
6SvRGW24rk/kXUHPOfnoOp5THotgMXXAuPyPSGC5QIIzho89JqMp4X0wdbRnajon6SRxwtJHu5Db
ywvq4VryQkXOJjZEMlCvoR5Ry65CuaiIzGiYZ8evnPnozGSF+NcqKPHmKxOJjjcumSFkiobA+r/d
NRIMOhFqin5+EEuTwqLUg4TZG6SACU92TJAQgEderfWy2MBUtW3I2fJCctrTnNB3G5Nh/eWUPRng
BJreWMEvITJnnvXZatXHwk9XMuRGb6P9z7CsRyvi0IP+k9dDonT3LQKKiwpKL5YoWcJTe6vrlvrs
NkWxzHxZVb6G6uBoS8EHh8fokf2IkQdVeHeJGbEcp0N6TjAnAmw548tsqgR+uhbjXwLSjUPbu6Fw
CuxR05f7TRz8c9oveYgrD3oPH2sNR+DkEy1hte8iBNC+DHh1RrWJrR8t1BBxJO0YjxTvbaa6EgKr
SuTv3aj/Z0rfZQzc0WbI300GjGXC+owuDvT/un1ul41cnbh9D5LsjAWuc6wmblOsJuKcRcxYKgWh
NyAbnTqnlOJEEzbpTExTJZlwHagrk/0FB4JncVkRdvXPkCRtPveiDdbYAPyDH3vPebl32LMd2ZG+
dGHx10aEfk+7r1/wyPBQi3WRXYrTRYvRSTXh0tkazkGNere1olqinspYxvA51Q1T2HxeldoDL1G3
asfJutktfjegA8rpw+n3gJpDw+Spbe9gZKUJqapsQKaE8Z4mLW7hWqay0CkIZz4i0fKWlPYcQEcw
lZPG7/MK34pRFYaozyhVn0C5OLPWpUtwckdxqgImoy6WG76RABBmI4tUPeyj2gsiB5E0MQKHn0NY
pRWQjpkU45zYAnQmqH01LkQxSln+imGMwkkQU6tg1c+AIKrRH9bp2ZwAPqXeCxDV165i/XbVQjW6
HovQYq6Rfet1tqPhGy0gR+HnrIrDFwuAYbDsKOYjQqHpF/y3TB6zj4BIyN+qP06SPZMADhM1ZZi+
w2GAkMczTFmFm9U4m/9LrxjS9ABTM3cGlHAa3avGkAsH+jsHohbAZxcyoR1ygvf0fXKmMriXZ5gp
JD92KC7SHvBG03f6QzwvBBza9rodwWndTjB62EKruf67a6kD/hLomZeEgRCySmwZurmKtvlpEERf
7xdXcXGY/fSp/BhR2Z4d6sp0r03+LDrnz3H8SWGXmWsCm65sfFU5XSsJqiMVEhkNlWcNrjFhRMFC
Snn65mUwSH7KiLBPcGQYCHp0gV/86aCMSgJw9zLojk5fKFZ/c11JO20bd0+RCg0t2XwG9osJ/Hlq
NVckJV7/FfHyQdpbzltlomKZ+s7Bc1yko2dRYEphzrSCswERpQIQ9d6Hk32GpeYuBwz/qbQW1XG2
FPr2czSLzBL+wcL2TQlWxz294neFJZLdQJNlfK/D7Nd7Xb97mHcg8eEenBREPjgr4LaiL1IJbz7q
G1PNikGxzWdid7qtlaqunNYA7vQ3pPL0+rU5XdRBM2wmcl+3Gbk9qUpH63wRhFJos6yDHK9YXJGQ
tpwLDfsoJJYsO3SVCRX9YGe3sltu+RBlxZH3rDiF38Sk/Bi7djnTJJJtYC/ht0fgDJaGDPzVbQRI
JC2XyVh8vx85sxebIUdi/q4XOn5Ws5PV22qWCo00TFfLWsdZGlG7vKN29QdIR6xQb38pba0ax73i
V+fIQc/MBDLftXhYKwkqGWKeqVbORaaMUhRCA7h8W53CFFramkaCWDTaZ23xc1D4/4xZqMFp31Gq
9g6xXiAkpSgA/6B4fq42z/e3GdSdh9/SJiiGiK3b2t6fbVBbkIa2PAbnRmM6Ze4shh4Ww/roIYH9
e4VTHGl37CEBpVfvP+uwLaEE5jbFMGBAaLIQiXhW//rrzro6t5VzIhZ9nVXxXbLrbxRHno57gA2u
EdZ15AR/4j8Ze3tUan+CafyxRROW4pcaJ+Kewovk5219ciDXnx+Pct52tqpqjQnwZBDr1tazScLJ
YOlqpOPQiuSpVd0B5YPMjkQ8zJy4wHBoqvf6Pkqex36n1kgM6s2BJf4lRdDMb4oNiDJqbZz0618l
1CXfRLzqREwP2EimzJkRJQrJ3TAj8F5K8gD+KbEgsxx5PMl7ZIAjWAlbP1mdgGAwp5GjVNyKUeq6
VnmeWTKjkfl9t0HvRx2Z4r4mWlDFGXXvi89P1Ee5NMspcL3YDohcQumDbQneOOiCxS83+sw0+1X2
3anJ0NHOUn3ot+k14VR7jpIpyZ+3CfYVwB7WHvcCdiUXsiwLFrY3Af3tIMy0aASNhgeqofQQfRx4
FZICvKlxx8GHupQScJr1Ta33HUG3ehGk6fGnBPrlqRTci6+jeGYRAeJ4Vxp3d9Us5qYF24nRqzVv
DM3p6u3X5EAK26PvGcBxMscuC4RXHErdg0TbMzBQfJKmS8OjHhY3cGJmCCZ4mdWMzEZBy0Gm/wi9
KF5qgE9Ap2PoH6swbo/OEEl4E4FGs340s1+OyOANrZBi4B6K9GYxYgIIvbtpyBF/cCeN31G5zPKb
YDvXNLtfv4GSUods9cQJYI31pi4ug5XuZJBBPTHLMRy19VXaVaWoOX8O88QmrjTJJZ/s3Dk5685q
2xW4Pe8kIM/jZw8vZyOF3m7p/0JRz1+seZk9IUG6gMNpqN8025dNeNhDRX8g+sNF8u50dJ5ZBpGF
bLRS091Sq9ZTkF28qFV59IcSqj+QLamZNZWu7HpKhrZtdJPtMRZXktutkv11jfdwa7DgzLnnSSTB
VA/9ZJFhSRwu3Cbh7PvoUC4+lQm+oQ8SQ8DU6JJa7M5Q3bW5s7qY6ldFxhrvKM4Klim08XeMKJX9
i0WsIgGPdB7CbK8ZFrSeNFdvH+vA+5Twgqq5LF4tndTDBG6M0k1o22M2UA5ET2U4oGSD9QaFXpx6
oYRyvv6IvUqd95n2zpYPVZqBmEf+2zizK4RdWTu0UzOA+/MmmSugUwn3YQNJ0fSk7FwBXLHC61a0
RQvQRyjWHhPLG9aej4da2WbR0CMoyEWv1jhYiptQ8Xr3sTZ1UZ8STZ25wJDL4BfBqr8F2wRy4xjw
h9goWabzlNHAeiRxWRd1mpyOUMMPYJMxRMzh48RpoX5ycK+UaAeUho+4tgkMOcg0Un3NDZdkzcKN
JNQBVUzsUgxu9+PQIwCOAlxBRnHefbQOy7PuDvj+hqUQmYfFyVDWDSQ36qkGAbmCpqAVSVhZJfUr
ZRyztnXmXiPSmQ7PRLJnkFWyjHXJZ9X06jDO9gNop1e4HeRO7B2oLp8bYwo1ae1XSGYL0+5lq/Bq
3yVKtmiTTp3LRaZui58kcLOxQk6j51nMYU6gLPiins24sBwtgqN6jHd5L8th4TqGB7fcA/KrM5oY
PBrwKWAEnYMxQ+dipo2ZvOS3L5OPCqnbpeHNbGc4SOavTPlQ2xdEJBhTeh6pTrgnxQLkW5pWgUag
GycNaBTfNS76ndHXmYkT8tc52XthRB2zB8R8FW3Hz6JiFxLACslgpdAAl+rbd6gvYghNK5/C9yqs
W/C6ZGI7MAhU6dzLNd8ORkBojK9/DbB8E5PEMuzb7YVEl8giOyrV6TKYRJ7zs48wly4QuISseKNb
ZlXDrwgEMpwtPGNTpTXbuxvXYC1WRpqi0hj1/c77JefU73DCxisT46Y7N9rMcUpTO7p69I1cGeST
kUQQSrg+zV6seHzJKTMNeLPV+hGV+0IKbmW+swYSekF5SYTpTaFFEa5aChTGKNwpeK38gKsazzOl
/pn3GUFuRY2G6SBf+72TvmbOJwbyKsGcN3ZbqyfgVHVkOelvKt3APoqKdtIEPIhdHRHR+ZSBpigI
lRQ2PBEC5FoQ0t7jpscs8WxNOW9cgiM95IeJT5TQVKKHl4wFvFfBaQCetdAESpIQlgIwjhzbzmlP
YxnkOAQmfKaUNk6G6ZMmJ/EnUrgnuzu/saXkfhpoioahOuxgHkGH9LVN/SZVMAL/+VrPswEaB0Ma
4bQtO/C7pqLxsIJjMvRzxmp0F27aU7fAKC++5VRApH0Ue2frE8emKC+0IDqjb6DYsDW9iiwDSETj
JBro+6nHWBtHd4+LmkNOkMDerkZO8Ise7JtJPNtldZg59h5yQKCBIOCPhSKGUNG9ovqzkgxNq1Mw
5sW48Lyww/3DCOCmm5oVcDR1+Nf0E9BD8bmpicWrGSAEDdorv9PkjL1mNySWZUoxxFEf2Aury8iF
9pWOrRrWmvvuMaIuBS6C0GoDt2W3b7EOeBZa+nvaSJyphXhGfri7o65iZ5NBK7Wq+E6hlDHCuvqt
vVJUQtOvEYZ5wiaask+8M4U9Zk2d6/UM+pEAv9wVGr5YLQA/ABL7n4TyVduSrZekex0Xq0UWzm2L
FCU5ePas/5kC3ynE0H0T/sA2xXU0yFuqG0vfH+NXrWRc2KXGjuu403pdw0Kj5nBE37rZ8g/m5Oyn
qK5U+L1riKppkk5iDyiplQ4t1JZ6QaNT+84Mzem6fldg6lNEDzy9XtjTOA4qNGO1wJydy7IRJ5dj
2nPkKHd65lePpOrq1Y/570CcR48gfRCEAszdIsYOPj6k+pYfD0WaiQ494gnesRbU60+MTMm3Wx0+
h8HrxZ2CxAFr+I5wmxNEYUT82V16lAXQempXnJ1zJ9Tg+CPv3nyzG8mJZWTFAkiSsPhdsiN1oBcz
5Fg5TTNcBw6h3wr4JPTrfFDtzIEKNgwJ/rv2yLASGEiKaEyIItZ0+d/9ZcNPQjhNL1ZK8IlnPv0m
4YQzYTux4GDc5zgaWWzKhOBhYiK/WwYQRK0UUe3CptrlBKN9eJuSxJc5xQ4rnV9xs8ZwviPlhWyu
YnwDRWmxgVITGKuHEUal5wx//g2tzYIc6PiCJHZ3A3rB3Y94f7iw39u6xFO7g/sIaZELA1mH0fUN
ZLG3jpcSJJ7qAgVX+VmKkkAKFSUOBeFp2VF/aSkvAuNXRIrEOy0/vsn1KlUSENo4CHcWdLpead5L
H2GOoV8fTSdoep2pZHZKB5QIzci2PXyJTv4xvTXY6gEfV/O7iDPxzibMOkMQmUCkkjfDgy+NPdMa
65ZCWh49accDfKTsS2peWRCO65ZlqpZkEuihQWQv+e6L9AooxwuATo1XZPCr8e1N5jMaRhF7JjFY
m2sckOZPms9Z2qK0eq2ZH16fBaHp6rzgSynZnx728RG4mUzL69DMS1gL+6J9yaYbPIHTEczE890m
uLffNGOw7DNKh0u4LV5g7Sr1CfzmUZpFnVs8BK4kc3zucWAW+4LTH0d7kiEPrgXa4ka8Kfordi32
uh3UN8CvFn3HfK3bIZCEjJnnrDlsZ6s1iFLVFk7zX834OaxFnza0eC+Z0pvBI6rrRyQM/bTbwR5k
s6JbRQk1RYz91BYesndV/6Z5DJvaDsiwZNLrSPCNbV1r6PvIhC461pIGo0on6ekNzit9N1WKjGjM
kavMGAzaOdevBC8agIPbEvhIs9We8fyyo8psKVdgSJsEGxpUsudoZrdTDr7FIfb6Of3heI4q/RZq
2LD7w0wDBd2Vk7B2nKx9B+t52IeLWpX72LzGFXd4IlAShPYd5VJDfwejlpRqXutevpypvck+Zuno
GuQkQSJCbZeQ72buAnsGGE420NpT+3EHE04aYA/cfhGCFKrY003FLyzWGBKSY+cP7yphKndfpivm
A/J9niVQa324IiKCIqjqKmPj44BrgjezwRpeB0d8MAd217VozmDDu73kx5kNADhHFQy4pl9P9WFr
8AA/jWfMLl2I0oQMgN1lmbh6H6qQ0W7YyYwEvw1Y+OhVDbyVG/mpnWcgdSnpkHYjEb/r/GyhexQI
X8yzYlPjbl831GT2PcKpb9FB1RjKNhBu2qxtymJN4K5bk4NM/5+24p8sqSQtckBmSOceOSMFnaxz
Vfyt/crq0YhKLnevt9aS+gsE4vVaHqzWAYH0Lbjja3TmN0eJM2a3o/BEcdUHN8/dIgWNAhB/JpXY
F1VWXe1TSxeLqgPVKOd6epdOKbVTGj6Kgc0eIgWstv2ogw3rGVDTxLitnZgZNGX98w3wbRgrgdhv
3gsCrdhCWMd3l0BGjwmkCx5v3aGKajPdiyvHTBOgtFX8HVV/dr+NFPMu99AkeCak21IQ+mL79Wsa
EGkpMKk7LZA8DYAhmLmKZPF20IZk+AoJk1/JHgy/w9L506v9gPFtnkkj2iRQLJeJaNaIpRHfOr7s
2EW1bCmtIxyJoogOc8QA8lPRyW7ZKLWwvCFp2ikRI8I0cw2k8eKhpbI+iqTP6nu3vDx3q+puGZx3
92NjRzBBuqH0+JdbmjrUAECWAp335oG24iq5Xwie0iOVcXK4hjbiitt+qITQqhWjM7R2vDtj8KDc
YaTHiStel8l+Oj8Lh2gDGSHCypRKguHEALHaQ/ouJaLoeV13i0irnPZx2E/wKmcus9vFSvejgkIU
Tx0b+NMEYwBiCYsb3XkloA6VHgxh7urO/vMcxtQu2DmutLuHcDVw5nSi9QQFKVdWQPtByzSXxKcV
nyhLeTATrXmKrYsF74DZbCgRLti1omMYzNPbTOw4iGxxqIdDthcCzu0BNjfiG13Sr1cRC2sEzvz0
I0SvlIDN4i64Q7OfmwNYS6//3atVTmgvJcDaxxxsh0IXa+Izgjvnx2imtMbHod5z2DNAuGw0xog6
/BqEq9dPL57OkuCqqoUd16Gl6R5DfBXtY6NYzytzcd3hSPabLRZOo+jjaykxa+s1oe4++LfBDfqa
oSJrAd0+Paj5JuAKBEEjGJfChAlpFJ1TmOkL98pUsy17gwpxE0cBWbZYw/IwS4g5rzrV9cMLdBsU
l9yhNiTd+F0AHWd+FvoG62NVJEFpA+lKrDoG+7CGK5fV3He3y8Dp11JH+18sm3jIOeT4VZ433FmG
XvmsoYUfm31oxWhP6i4Mr2XWSPRJ9Uo8Or6J+S5rJBcIu/vvwZGSQT7ftRqO5p+kYAw37m1kIaoD
6GK6fG5jcUpELBdmTYj/ZCIZ7nU1dUiE93EC9NXAfJgywVy3rJG2SFjYy41QmIE9CSqtT3BEsSJD
4NDTeG3KGc4NsOuhSQq6wRSO/x4naSh7t4N4EwLa0ps5QgbXUiwvBTSBLGUof8MtdkdMPGqJtwOn
nZWy+Epcb1AdiOj3fv77KHDEqqWiX5tBlFIHrc0j9JZMnWKK3WRdNxsBjufK1xgkwtFxDsbGucQW
BgwvXWUQfro3GBpKQQona836QdnaKG/ioXkzPyLUq3PTxDSNb9TEm1QBEDuI7Ji+ur3IhHOpR/6G
Kj17PWzxZNd3aDzFjl9vnpDJnyWoRu0Ij3JovritaQutbBr18LkNU1FqAbdzJkJMPYRe24LoFBII
Cnzf8TuBhYXvNAAXHAtAGhV3OzZgpwCTCf0BrQxTqw9Jcb/ZWdZXVJmU4YdNA0YlBlpyGHsDzC4I
irGUV3nVD/0FsqdQCqut35bWofmv9oUrPRMFli++Ib7JEBuzSxn7xCmljTAIwVm6M0Gayu3VFdq5
aoP9ITQ7Tyyb306CSdPzdOG+rd3H2AFzikvTD6ZDRquNtBcXEo4Mz3Z2qoePEsEPZM4lGSYGA8Fk
HCqMMx/FJdRjJPZl4EydlZOdJiMyLE/8/EUTJT/BOskD5T3P3xILOutgX8XAwqRiJUUi+Lm+Fmgb
tcA0NM9l8Jv7rBLEUnt2j1+Lsa888IcFQmdKvLlSN+V2VnMWdLTQKRyz5VJt7bSiEb4N2oCrJAbW
Ej/9uc4EdzU9vFGimBE43m0GtlKH1PqEpped4R9gt4oNWSBGwt72WjXOpCBvG8bq/hqzRxlgW4yE
rr6znpwgoJuTQUxNrQb/C7DE+qUKj9C0sUH0hcyF+sFybP5EeEpLfyDp8tfAbuuzR8kN58RHsboY
QFDp57z0H7Vmy14HP7m9+TQ5Y5IlO3ljf5vRWxVveYm333vPpD7MuwdXNJ0yQQaHJQzrjClMBG5s
V0nsEMkLdRurmBXKBEiriRoQSY+kPoZDOEOx2QfAxkoEFgcdkAv+3Tkg9giShduLzRdqzEe/7QzJ
vCr6hkjhThuF+mczrIwlsbYSOlURoJ3nSUjoB7o+8nQ38VIKIYQUTQ8yTPuZXw8RCc475FIuer5t
7ns/SsedLVYFRhgA2MNU9lV6Ow4p1I8uKQzGcSsuYDYQ6iIgbi+GOlVrGs9Z8WwKZ5zo2rjk9j9W
e6p/h4rkc/zaELLFANyyqrLcxksKP4VJTAPwRhCHXquP0VIM8Do9zRjxzxbl6vCWg9+tMSGk1dGy
Ig9i01NonUIqmUNXkFKUeXM5G7mpDVE8BXyh6OyWuTDTr1NppjhmWGHOjR/5DQJkKIFH+TcDUpXf
NYEx5r0LGjans0kQ68PqqhMXbjhLXXOWYywH7lmpPGyfETv+3L5FH5KtpAKC+3m1Suhd9aQ8Sz77
I/PeGK67zWZcfs88JSOign/ZvjC39kgpPYmpTyBMX1LACpYL6/ZZPbSSZ4QpiZIJr4pFRyYvK1pY
JBewBUU2a017R2cXhUjnY/WqTxbuUIVbhR+F83ukUmWwoxAdHKZ1WMwYrDV/eqVkHj+VjCw+H2qx
J7/wjhpoXxtpkZifGmoIbtU95qKia0CrmE32LkVU8AknJAEiZj+RgDjEIjfDsAGPqE9aqpjVMLif
ROj2PkLVH5Pu6J1BaAUzXIlIhOGBskAbWvsDWT6lMJNAS/rmEKYTKDeVNspXuEVKg4MBfaUC3ydr
k6gAAWUafUfXU0yFgIbiJEP7Mk8hzQKecu7dkjvfEJELfiUK5VpVQwyJa4oz3MWH5yr3unKAJ7Op
ILKvg40AQYBWXgvAbr+MgBZNlThauH8xePzUAQwqnaao8r0t0gzlbD+GVP+IQcD8zxqyyF2uPJeo
t7alFCO8k6dPPj1tOuHfW0KkS9HFeOrsJsmu12xnDApOk5NbjgNibVyyquQ/6ugg6zCq3Ehr8lnT
EkTvB9GXoG8GneBo/+M+i4ffk1g9hzVnz6MH6HDmNNXh5M0QNtuagvbwfr1ELYCrQKTAlSumhvcp
EXcY1PQCuYQ5BBGAI+EoiySQz5qwk8eDLF6TkvivTOP9YqLq6cZ5KI76L+r66JEfnOYqASwIBtx1
qCFWhBLGDVLpIhpHso4NdG6B+i2cwMYqz7g6OeLtWAiEYUQpNZUP2C3gzELMK3DBruFzCnjfKOiS
K2YAKEMfROyML4n81a6m+RLeDd8/tc+WAIC3vaTFTbCCdRfHVdHGCH1bzJR1PTz7p6QZPeImMD31
GhiY6079ujd5Q1xcwRvA8DMXuBNHq8X6QoxJmpeDsWhwN6C1z9twOOAqagIqECTvqHDHQChuVoiG
LtsOWBWe+MzVcqoKHzlQpK1AVntFMYFuqOcTrUvrIynGggYEQn/5JmgsfaYfLg7yYgf5EIcrkYgU
DsnrFZIQ+e0pHVWkh/BkwAQnUuHyotQYYR8AWQ3T9S+46MG37TheV2djVs14yxaCpSIxc5c08ifb
0t4g6Q1PoYbS8XVP/h1vtWJc4Sjqm1X0w+SitUELYBDLJk0Xph9Ow4j9S6WxgGPvEMsAF7mrQcOp
N+kPEM0600MAtauBeg/78QhpKQ/GQhhbCxogz79KdAy43x1Yulx2ARnp/KmiA+PvTZ8TH9Ze4GYr
/Qnsa5GmgD6dlilrjbhC7ckZ97FAtR/jbOiIhtYmZVPTBy8A26yEpaeMsBe1GkGRIUXXakR4rWPh
elbUTPl1Apvx+fFNcSw3FV4a8vnL5Oci63OQ1v1CdBe60QlGfv0opE9JiQ+Zd1La8u6IROOW2Zxr
AmX92Ghigh5x13vw7I/4wrFEEIDNO8WBonBHyd2lQxor5F4lcoU/ytIvi09aBKsXW3xDZOrrwPyo
h+6gX/2TMVznrjR7e6doerAsIJNFT+k2mrHkBpQKKPAQ3oxs5tRCpO+lSyl6hJ4a9A3B7Fn/BkGe
NJvYiAZQ3wjgWRWfVYU2moarVtH5kTna9beRjzdNZraWd28tE5+YAsr8qGAPOzYz0ItohxEoka5h
My2KInlUUAOoendzmfTVeVYr7XXbbHDRgztxkE5AJBpn6nHBzehLVx15Czhm94yN/e9UaAvi+apA
0vxRK2JVbotVWYx/wFQRFWN6bX70ZgRzhntTXTSCvOV8YFqHQ+ildXb85UgnPceH0fmtjYeF4uCt
o78+fcJQNRYkMh8rBuh3HHg0hrLlhUJUH+1B2e95NS4dKDWCacfaZz0g11xQ1iDegW37lHSatArE
bU6l+UpDlSC7NKt0UJB/GOBjUlbO8PrkM8V5k2NHm3CPFle9i7Sxv2atBtK9bLgmtgUotFzW1ijY
ekcOSaVxZbaK50fMjZLTU5xQsASn6zRdDIbr/qWRgeorDxaGtO2/L9gl9RBHjmJJLM/JP67ElrMy
Yye0TObgjk/801TTPV72dvmYGRmdx4QApX1itXQkYzcXqc4bCgrkMOyg8qzhIHWNRuRk/R9f+S81
EyH6E6FimPUb+wqBu1++vVOnGgJJKsMieG7ksQwp6VUb8khzNorRys1qIP1JzV0e9e1WWSLQF55z
eJJKHDauyr1tDemsQYwyjU1vS6GiHw8sz44sTcjpxnvPwGLfmyJYK47TR0hv2YZ85wMu/zfyJh+n
pPFCGi7LDC2bAXtI7l9q35z2GMBWvxi064jeMXnn+OVV9TrSf9RDNZ3bUit+cufO7AmuScU3kEPU
CVTXRY+7bnYEJMme1kvijlm/awchhwubU2CneSoht8Rhx4km2nxogo22e228zxcTdPi5Lh8g+Faj
0Wr+4rrGKd0JbBbq4U6z5hn1Q88EnE4mke3Z2IzyWZFHnjBt/HrTUltZ0Az5xGfNnVOuHVUAPUVC
hSV71p0+3CpqaOjOwM67b+aXv8MjfLrvchwg75ggYViVqLJ2ogppvNfKs4OZZ9Y+UDd+feoHf7Rf
R460TblwwGBjTZRe5XzYDePZmt21nrhBZxRKiFKB0HFr6JZ6yAQs4uVY8TR01Bpg9SYz7wsc6r6Z
07SzdOUhZJzlTnIiNzUhyD7LQ2Y2FjHD9bkobLNNKYRfoZZB/hi7OLlNagYzBWhP26P4MyneeuYN
7eROhiNjYSUEUuZHUXQ5apFcrctoKnIKPBRpHr9DVdeNM1eKFloLu2enSA9aimnz64Xw1wuJP6yL
mKTQ7cK8qjoccq04rppZCtyyOHuHfFM5QEOmWWaIceyo4uSjYpX5t8f6FT4BVZSnHsy7eW+H/1eN
TE5nfkG9L5eDQW5Gyzx3Xjrm8BsDY0JPBx8qrOGU8q0Mz4T2f2t1HHqlkZx1LIkseXKOqLOK7Tlm
9YULDnZ3D1z4L760Kzs8iINW/LMSVDrV4McpUwe2dX1o+DkI5Lh7r6EPMQEIGSC8iyOkOXEjaMi1
yam1YPhuHuCFhsSiOW52jcVJv6GuuA0C4drMvFlgM0pz3I+Vn+jZSLFn8QX7nxW5jBi5OPdE+Zu1
c5usbBj5rSYRmAgxDVL/VQkx+WNw21/PhoI6iOrRGAZrxt6H1qEipg0KrgoYGyUg4k3KBb9Ry3OC
qPGkBtwZ+s7ljHk9O1P7WKXMQ8JWDmDPBfpjTJUj16AgBbrrc3OrsHSTUO08xYYh4lD2DqSZCbDd
pwKBdC51EhZGbwxEC5l65HsulbZgyDhk76MnyIkbL9TG9annwUNCe8OjASF7uSS7svfH5LzKttIq
+/ruPlO2AQYM6/OdZxpmPdMbZAujuAXy1j4iE8nPewKjUdIPF6weL3lOWUuulpVVA66jZJfu4apz
ni65nDtOkCPUVasUbwEJyFl1e0qSZQ8cGD+RTVEXCLeWWx1XPP8+BOAT10qplp4TAKoCLL27m+AX
di83KuDAjpET01/GVPb8c3I96jmMq0br3Ae15O4ZFURbEe50kMY6ARbiBNGqUBaUidsCy4AtbnEX
MNQMtT+U37CsLtoVqYmEVdi4g5VD3x4oPvYQxGLHqX25qD0pwpNqR+p3C86DXjPWK1slcQOtygbK
msSoLm0hwR17zpDozkz37qjj9bugykFeWu98QigHwLPEWb7Hlnwejnj+vLBhLOhz/8TJqp6kpraw
P8oY/lLsMh+JNaIXuqf3nB7R0YkyeO5a4M3FeaL9IBSn4I9Z4ySDUtwkHFf7gZ77QPKDcmeR+VQn
T1ObdJJl9IjYeptcRCv6WhI+WoMNtjdyWNA9Mr+ZeA42q869aBDQScyJYKwVAvMBQyYW7BecGgTf
AOqCdiN0p6khtt0DoOvJ8yvUpHGZDEg8/+PtitzgakycRDkgrKkow0kpKhWF8CTiJmIKUjQjZ/2F
3jt7NMjP7fxqc1iGSU/5miE7l8csF5fz3H8HegrMD9x0jQW5hTXN0RGlb/1fQbsHmGSH0g1qTyqp
E4a/qUGcsnoZs3ZHEYHTMaOtDpwNsSC/m3sZvnGARPx1HYXEFaHvl8FgR1Z2eh3hPqg7+ZALc2M9
AQ4Bp51HKQO7K5BggCtbd3YhQqHllE1Om4yYC/x0e4obF7kgRVJ4A5H32eJMg45p9GZmpPX8nOm6
3yoW2kZkOxJvgnBa/zxjrWhFrJ+/5sdL/g2fvAhdsnGOfd81iJG2LPzM1IXnKz+xTqASpQYEqqyN
kadt09xJouf1oiGO9VA6t03XG850ntlxBHZW6iP1+cyUL2suTQYg7ggyyVc3PpmvII4ry32z0HyH
NM8gbQIbCopwc9Pqdz9fYP4C6Q+b9RDcSl+8pEFjw//bS48KUiJTgusAUPiTVvBROzEdutsiwXLQ
PmtFsR3yrgh5dghkUcDmZwOGOKl/fJeYO15gcvSy+lMEyC+4/0Dq5s7rO6PHXE+iis0SEoOINxEu
rYlBNXw6Nrv9V2vtdAUr5kHEZNnoR8qtUY6Pi+jknXEODJM4ZYr+cmOaptFNeYr/LomwQ/FE53bF
JrOzHjVYH4tk47uG/Ci5JDfETcL8/ahWN++g9vySaIs5LGk26KbPcZhw6jRirtyiZCk1zavmizEI
e3nVri/IptxEsjphq9p2/dzDL6vQ7EjCLfk5Axh8adr5lYSnIQAjP6qjFAVv1O/zsOPPTVusnXyd
OU/Ehc25+Y4PFILUyASPcs83kOjTszRIeLKBFkRghob4QhOnPsKjYdQrJ1gH9g17eamJL1mUXE0L
u9bTIqkBMzOUC1ZjeBpcPRkPYlWW1zzJWUvN50mbG6D0WUqy2mWjR7xpQXghBhnRPw9COzrR+kHt
sA8dgBzSX5BFmF4dfENM8FezT7FoIXFR2fS3FikieDrrwwTaJcSd+FEWrwEdScx1ZRdG+yiu4sTP
siU3QDaxcIbWtwD7Eobd23U76XL/gI1gs1oqa1k1uZrD9jq8E0Nh8xUnWmM29D67Mhs7cmj8U8ai
FRVjU6IrB2hoeV/HOQ2Snl9tHVQ+LdXTtmxZq4cxuYwksnOT9BKpqLmstLG7yhN0lJDeI9zLlVgn
4tuHwEU4Ithdh0J5s69t1GSLAlLi6qoGF1KkoinDJnV2w1ONMRlSFPgCvETpxwiSEaAVgwA5n/eJ
P8O3vM4Ua4isAOtqrFtrz7wV9isIAMK4v5dkhXrBSigmYj2C+U81PHymePY44yfzzQNG+RTjxbJD
EzpSO6CbLT1pWb2vX7NpLnMSOJVHCpf/8/6NKWBELofj8xgdzDd3xV65meYEgUZ6Co9nGt6lNxQL
Uiqtn+HA6IpxUujJC/vKty0R+fiGZ0HOY2dGu39dfbkAqSRBpWeY4Qf/Bq3jdmiti1ZBg9kBeSnl
04FXx2VuqOMKPnqxF4jQb+cxmZWE9HtTHlk9A7QbIS1YgRU5+2RRq91pFYdEeRp5CjvH9cjYJ4hK
4JId2rHjmrF/bwAyszXk8IRLoMX6717TbrPjJWtYLeXWItZT8eHji1UazP9oL/mcQAZsKFYi9gpw
J8wiwDZu3PxVHtvXsvjCXUThFLDScriDP7/+UVqncVuwUxPSAZ8WR99wzUVXaAN/fic0waNr23nJ
U95a4gYjp0NTSmtTIG5+Ts4L+Mu3io2romAISo2xqa8BkJK54yoLGDqTLbDCkLjm+HQvIR2T25dd
ByWYtdgXmhGoTrQO2AdoXqBzh8Tb+w/XO+xbOt7IwmTFjnBtUk3nVR272AwaN2BLWOpq3Swyhc0Y
xupbwOVpbV7wB7fqukmLOFk+RBmw2C9BmWqFnJQnJV14UArkaBzYgZkXZECd2z0fFRib/b+2CeeP
PqNLdgqyD+oIwkvPx4VQize6bAZVIgJI4I3Z7vQVYTZ92DjZTASZbx4KdusWWBYG7cEFuVLhuY6E
tdvhqfOeZsOsW1Znhate4HFlSLhcho+cugDYJ0FVluA45Kbp2WtV+qCmCAows0Q7WHD/cH56BOA2
h62W+Y3gvVIEHRD2ZlYqlT7+otzmjwdUckdeehJZxV6J6eYZD1eFIsi03rOnFSHJHT7C2F0DoquW
53YO3xJuSIKrREZD/abbbO0pXVUgRNa0VilkIEBQqkaZ0Pmyb/VHzE+ik2ZUwhOeLNZeIyWaMAqB
w7lExZeKaVM5HdLQNbUc/QKwPGuq8HRUUvQR9NamrxzkTVb12u2XyIp8Oq/370VTl2+4p5cXAF8t
+mH06g6s0t5dOZpnxTmVI6SOvNN2kb/R5AyGr8U4+wpc7fxVO+/6JzQJrkazgxyjrxV46TzNCTlU
F3gQ9E9NFGq20JZDeZ10QSPrmhti2OjrtjAJZBa113M/1Gc5USTJqmUWTc/2qLUkO8+DyVq/afiG
HGF5PRENLmthSEkebCtrY1fQD0fRWGWkLnR8hYHxrcrxom70JRqfjaWk6DUhmua4MhgJr/9jkI9a
XjqvqVpgbq9wM/kdmfXnhXnTg0cBm33tkoTPnDJB1LFCJR/xYUXsvW0ljTYoQjFqgbYBD6JvEVg2
UMv/uEPlKpXAIbcMDDipT8cMzZ6dyGMSMQdLm26jwRdAIleqICpuo4lZKbzgv3Ho2Vn6CSTde+kk
/8X+RQVdHNbthd4UwmposqKtCkRkZtcbYAtikBl0tb+FuCExZO8Tq//G8xJaXeiHEEcCttnw8VOD
9HlJL8+t8pqtwjIydNncdcnJ7W7D2QacQ/l/+gcTY9YYY4qz9/YM6NcabCYjEufw+9XDP3vs9dRA
Y2U5/s1VK3t8nr8nkNuc+cp7BwkWy8YDoMFvO8To2NCqXrL5AZx9vBDGBhqqP3c1qxlgaX/Ro1WW
N/cYe28WraHSFlNeCzksTwJA+i93nBcaquLf/ojMesIFvOurztJHwaPNKWOC4lyDv87FY5nrsqcS
VHGi59m+sm08HGtoaQZmda7JD95uVIRqs4ZJDDh9Xc9Vt9MGGLtrvrL+27sQAAcu17t6q7NmlRRE
9dDUlzdanGSyADaftjkp19ye9zjuAQKgFPI6qZIolws06lV+TV/p5jUFleJSzFeAmQG1RB3W5eDK
7t6NP3D2sKUkCTgKc3/sfABEkpA2lzO56vLpTUNJ92to2siu2akPfysd4Wg0zwbutNmxt+jQOkNa
Acu8McjHdLuztV2WSm3ZRTW/A2+D0JUL8shmnzdYX0Ol3rG7yAohvYMEG5s3fXxEj/e78FwJB0nZ
E4gMxzPy1dFQC8nd4J63v/nJ4LLGQRwTxjIn8I/a8ILvHz+Umsx25ka5k8+iphGRfKxdKrW1s2RX
fQEmirFvemsO9+Po+R0bTzI0iLwA5Ovtq/xberIqef2RhUXIfm60SRKw7AD6q4KEuapDcJXa2p33
2LSeSCXoyJQtOqPni1nGp8VH9O6GyN18Z/L16osMwCfsOyltJbPXlYapftxdM6eOzWBSPgmSWnZv
URctqS1eg6LCzv0mCTYAzYYgESdyuxSW4JLbh9pG63GCW2coScLFU8z7PwmNrVOpeBaj95DClIaq
j2r85zA/lHuMdQ7xer6iQhrwK8kFuqO+66hvmsKhiVofOGX0W8XKGJSOdqYXVAlsauNoJVWNzpRu
yHsrK5el6z+BftRZNB9DTSU5j4aiz59UWb9l6OJ0+3Nznr1k30VrQNzyQF+DL6RsxfwFB7B/6SOM
OG03XHX2o3qggPJzLiKiBq0a4IgbspRuUpa/MGOXABXKvVB1gMChDmjN5pJNWQGeg1KH+EKzNaQ3
2AF9ER6QU63UClUN8mWvh4WjwDIPnOxqVMSv5AANLuL+XQSirN8ZMN9GPtfZ60iqYUJ7ghfzcZ6E
5wSgVTf9oCcyOcMXwqTIp2BZfZwG1vzC1FVAnVSAUIndIEvl4dra2A75VvO9x1fI1Ia5Ei2vwOK0
8X4qdrLF8qBlzdz33fG6trb8bmo+3nX148GXsCfG/lsNwCMdFTPd7kh5o7A0zrSqN5E99yLGw+vv
479X99eH4l8O5OWxqEBZGF7qEIDC1Kh/hIw+eDAEYmaWfpmuA+/E8JKbaEzPfkyEtvJCOeADHhrL
Vd57d2maqX4jbHIBo6TRvFYQEHQ6EnKeEZW34KTArHjTGeziwkemT+Pn9GkZhmvonWjfHhZd3/AF
F45NPqWy0UhN4p7FI5naEWcVJnIr4HW9a+w9g5zNLyy5aSvKLZntfdp5lFKN5sh6bgaTLLaeTC5z
sTbmGVanyd0guH0oPEFKUDVbNm3oZeuPGxzNNt1LIyI+zAM8/B/5PmjiGIJj2ou/vC1GDH+R99OC
qWHcD6NA+rHDNu5cQjI2x+4urG2COAaenG33WDce3tKw2RZg7GMhoUxmyALikskgsUw6kIljEM06
pkWAYbdDXbbh28fxPiwQ10gsgTy4be2PLjAVHUwnpThvNIIe17/7F1/5SlCaYcQ+KLdcDGmmhyqT
MY0XwbfQcu1N6hWrrRTUsOI4Nsfn60x+BbZwG0zpi/3V8wsjLS1b+gUrzQTVCz66ov9HAEifb7zA
nbSeifxifqQ7shCVXDohl7fH7rM/hQ85EfSI2cq8UKusoZ8dyswAEmow6CCDxXMNf7Yqw+N0KbsB
vfOOubWoy1GszbtZElDj7LqJvRy7djiksacrtF1NQoETR7QXgSSG9qN/TPwrnlMp2Ujrc95IJ4WF
VPHHtHrwRzgV+oxSX6O0Fift93rp4UKlO5rYW4d846YbK9E+IONg1yV0/YmBKa21UWl06EpoB0cz
W7lMU8aWHGkr5n/jZz9EJI2G81YkH16eZ07e+tW6HgsWI6hs/agTlnf3kSV8R1J9CCd3qwYtkIka
xxTBjNlMAEyM8bq28nI0qSXYQMvR9c19BQjb7VtVM1nmwpYP8rRjpbNrk8sCjyNe2ooXXnfG8dtk
7FVYNMdPcNF0KZttJy9GPcBVSz6EfDTf8106CJ/WgNv+RDAWxgji2KtQt76F+nT4P8fkrccK7f9D
FYFY1L90EyM51CEO2z3yL6s/fk1TGgg/u3Wtp5U0Zn9gupgEQgk2OUjMnQ28nmjUNEhIs5XEhN3I
mnnZhXsPHAamQ6mezAoH8BiU9avRfeZ8UdsX2f6lcnaPaN6v4OULrn7uLSo2BYXd2bYiAd+SmFN7
tQ8MzqwBW9GtUktS1t/AVh+6BrDo2Rlb0nPkbSczXbxRXZXTzF3ZZWgBXNWL9x9QNDwYiSQGRR6f
yuuKIqGF8uIR/PhNixJAXhxwsNIdnR4JGC7Zxwn1gly2+0Cq2FjrQiotAYVoWh/FYf4ktZgzRuLk
33IyRDSSYxONJ3E98QjgHK4AtFIxRROgVhIFV+BOL4zxyTBsrc1ZLtgCCJOJmi2GhmJ4HtcCxNMJ
IEkhlBFcTDY1+NuXkRGJuo6K4Bc9WkH4uS1ArYpyMG/rP7LH3edJclSv7xK4IqQCpLw+XMo8DFon
peTgsOyP26AS5bHvXgh8/1bvDFCCOi5riIQHd+YP680fTiBQiZiyB8uRhNVES8NAVBxHojueAvtE
otNxCdVZs9nOtphzTeqAOZhZ6SUqPlx025OmpA1aJ/yJIzavi0DHGtYiLWy6fd3Rp7lDAi9QcrhT
x9WAwwrhhFabeeJhZMH9B4sMsIMesZ5oZlgwfHgHM7KDMLaAganpFZX4q0J2/N5OZBepv4BbyKln
nJBZevuhQEwVBpq5XYqRX1D8+KSZRKzp++Nl10q9BgmyMsO88+C4iVUuvPXYKFltBcWzk559NF/0
+YxdJWeYtsnNZxGO+mAybC1jstY7ykcAFnSwkEA8xv5VWA0ZvZyvQzeIdWhKEoUHqXXSiWoBFoLH
pcgMlPHWDmspANm2I86Wo5JtKnwOOC9vwX465kuCz+JQ+eLDcA9SXK/BF0xlB40dyVo+toLA7cUv
ChEoEGGisrrVS8+nyRpifjkTl7b0sC4CYHiRMgsT8iwKkpWBdGsBqQlgSwrRZSxoCI+0CAa8/Q2j
NDpWrYAS1R4UtKB3wQgcwiGZgg17y9wCQXDbbjtQdGgqX+45Hr2R704sZFPROblJw/gf7sLELIX6
k3UIBytNd0YZDsHqWxdlkenHcgUoYTP6MKZ+6Y3fFfe3KyteW6azEFtfZ+F3RjtCw5gbCdOM7Ntl
5HBr1ylhdGtY0j2IShxXTRFZXYKjx3goYrOyBEA1mh028xkar2H1fmJXHldI6Ctgq1RNHyYN8gY4
wsjp6Dee3qmt9ECZnHwLuEq2gxUYAMrgySuE4KelvImxwNiWoLdxCEvJA9iMmBzv6XdsXK0W08ei
tW4x1vtE6wwAsYgW6RDU1b8Qz3uagnWUGsU1orSQBun+MKJkT7AG5sfCpHtbAwSU5Z8JT6sNFDEP
nCBQASrID05CvOgwmxQ2m1I/GXGMAuS8wV6S4eEi8APfbTKo2KUE1459+k18NqXmQ9iNytGaZnUQ
Om3PcC/LJDsMcwLh3mKzf5qtnVLNSoUYqd7Qt8KX5wHatr7vV1yiTEZILuizFQsMQEYMCpa0SUJe
KvSveakmSrlNW/+8yQ77Dw4jH5wKgT055IWQuP7hsN9tCYHs+DWL7BGPCWw8Po/bP7Fs1Hw0JGs+
vt3ISb4qaj/kj8Kzs7Fmj9kTDKWZ0OkGw0Q85idnq6BYOVgG3vXja6EEqigdCjq6zHFmJYVQyGfI
6I/WNTwyyzXv8deBPQiZXVd80ixbCAS03urNu0uD/+oH4etO2tR1AYTS9zE9bDu3+y2Ff+XTWCHv
RhOzexU5JUVwjgJJtElizkd7SVuBIVnRNBVzlDNj3XnsR36n9HHv2QjEHq6bmiIGSegslOErJ2aL
zON32cAmKHrEWmVcx4cRHIf6+q7SfiMhN1PUz27Qshses/781rHx6GJx0Wp2ErCkCx/nAEeKV1I5
76XhYm1vrZ4jYKsF3McHnVMTOJBGob/krJdY5sBFEHbjWJb7py95oQfLERCwxP+4CkdS8w83G4mS
GlyXfCDyTnXZeVV78u402CDmk3WLl7Q+1Idd+mkJrQFMBq/HxNMnKamNu2oIDiH2IqG+LFnGE0Q4
LjCeBVOVeSnxD9SDogjF8bmE+/Kp6AFwx4It5JvN/kJuSlrc7c4VmM+eyo/HXTYxu2y/QHWolIBz
qY7rOuq/lQNfKiM/Xmtjst2e4Uwn6CG2Fsejol7HKMEB3H9aQfbIuhtsvSxpoQBw2rmv2o3v5ZoP
0Lh3B2eB575coGDJkOZNKCwxvz/PWMmn85lNk1CateGP4LnD/pqmPQqvfcOgjp7k3PoIJmyxBluC
jn8W3GA2tlBFSWaXZB9P0InaHTF17nlqpI3lRShVAN0W7+czIHQSOXtbxQt5hO41lfWeQVBwSlvq
02V5BtKup+UfdVILc+stqZr8SA+BKqH5epli1xvhhTN4YoMH9Bd3qSwZEBIXJeqfQCFlI5AIHaeM
AT7ojipQC4pV40T8ojvbG+Cz9JJBOFzwQR6Ng9p2DqVKCZXWLTBRZyOipQ5xxPxPsVU3qPz0ZkOf
/1BZqApr5oZmemGeYk3HSaOHgBEL7Am0yN8HoizpatSnbtcU407OP19IB0cvGmDUCqGqShVKdBbm
TLw6uaPBQdPMzfdikzjQBiBMOCN/x1nX2K7vgaQDoN0NOHNYzAErkaHZ3F/pGFM6HVByrlAKr3/S
TtfT6a4d+YDFAvAC88dD89zGXrqAle/fkVxWh25gt1PAxSfZLWOnyohkiaXD3kHv73tE/AOsL3D8
9WhVvxInI1I4HYluFG2xuM18iaCMrrIHjcRuheRS4w14//EqD1xjozDJaJ8O4UycxAy4HQzLp7T1
ViBhG1vxaZl7bFbo0ZFd2niFbXqM7rwnlL1MFQ8w/U8ho7unzJI3UqDMO5v6S9hvUz+Ps00ZUYgK
uJZHC/5OMFtf0bQAhrL/6irLDjw32WgrMKsMI4V3ZWGYKmarsc+9mf3vrXQcFEF/MWjkQJJ3gore
a8c6XE4bUKPNX/wT9Jao1TDI/GUozPFSp2DXeQbVONBs7s8CTZxIgTAOBBfGVir/DNX3bYVKZpqR
k18HGn/8RRuUOG2etKvXFNsgjqGg6wkF1YTzb7RsVGDeC1hVLVjc3fTiD6EOx67uJuKyKFkYYTLd
SAVvlO1B56NKFT3OTyYNndvOzjD3Jbr83i81sM6KUI+ZryPzLWcQCIvlc7mhnbWV/obKy88HX7Qa
WHkpvLwP0cEAMwQH7seZbjcsDAGQf17seO2GlgGOkxy/+hTiDy/nEupsTFk1Xvsbx17sRrw4vh4v
TCWgRPzLf6mzBasOnBlZYHLV/zUU6FZ7Ju9jmgiO++csv58vJjicFH7LmWHS9x51L6OrECnLWP09
WyZ+PsysdRbuvLOstxa2EB4h1z6aCKfVe6kKPZnw9i7/XYisqs/D18tW/7xbA68qyY1cT8TaKQFt
gS1AoKC8BDXOfltfGHDvbySP7hcvVb+xTVLs4IcDEze4vn7WU0NQuTL60k/GAj//cLoSvgxUyOm+
U23u3V6tTmf4U4ilFGQgwX75EYf/F8o9C4+5b4ofIbe2hJGA7nSrR6gi6sYO+9hMmwWwV4JFUL2W
A/6Bj76X5SVf60MIrqVF5JcHcVwYOyJbu1Q/w7z/vX+41A1u6x5aSew3yKUR7tQ+FkoRRlIdOdhj
Cw8r6iYJOKNpojO7/oBjkJxmbmP3BVk883Ge4sis9Ii0FwewbAlm4wfYqgqbg9TUHrVhFwNOWFPt
lrONjQ9j76e3rEe1e/LBA1R6+shp+OZI3NpjTjJMOHgsuEr2UOP40XOngcg8ADF5bcwKtipQ+b7M
AdNDf1UJo4AJOY1XwDIonwS5xgIGKxf9DeGJZqM60zaSvu0RqPOI5/cE6PXLldof0JLnX3wqrcWR
anC/X4q4m3608LXJmlUN+0EssTu4bGpKsgWmGS2R6V4IrrhqHVfBE2pNbKeraqHeQ58SWJ7FWCDd
6mFEKy3vwCoaG/yqxSQCX1glcN+lCbnryV80GbSR6qzNx01cLDzILXI6TpJoNjYoThWTH8HNMU62
EWHg0wnB5+vwpeY30ABwB2vnUPbM7iMObpmuA0r6wdcM56+uT+c84jvyHuQmz2g58ms99321W0EC
eBLLxQDnBpsVXGHczMiBFr6K83TXnmtukeXYrEvCbECFbw/RMFf+iH4isQ/enw8MKPuMq4+X6vMV
ccV3eosBu58X3TkZ8y9ixUdFMYgQ6VjAIYGAyiDYS+5myq3hf7G8jsQ0sL/TuIp8CXokYUnhI72A
WgT3TmNAuDK6rN/E1JTNWSJ43Mofb2EhoXjb4ogshLv0gkyvWovsTqR0g3Ht5WpYYdPPnfk8EKHA
Vz7VKkZPnht1qW1F+mQ4PMZ5AieTK3Op4opZtsoY9+8Hd8TLf0e/IBU/0Uc+u1KuSSaWAMpZh1H8
EPvOwksGoltrMmWVonMQ1ATTJ/hrHVIRVHi3h3Q8Z3nm4A7ez2LmT4/YLkYsM27Bgn7Wy8cE7Dcw
kZ81Xft+3EcOqpCDPURQt+c2eSgguQO0FT4Ef9r/Me2pG7wYpdz6EkBw+l4Zth8pNLW8mL3/RlOa
Zg3QHgFUNBbnPdQMeXXs9oi6EhJJOIcYVI0JqyiVkUzW4UINCGCKdoILxliyHJOVeKSL2T7DXG5b
RdkN2979rroz1mOpcdV3uDYgwGyoyJd63l/A+mlc4XBu183xmRrNi3G74Q/LpNl1MeCSR1f9T22q
PP1bzFhYcWh/mhAis3HH9jdp06MQ/mmc5VUpz5GGBF6C8scnjTyGSBcA+aPiMLMI3bAj5ApCJR4c
zOA4I0iEjT5DpwMBvIt/m8o4i8J0N/fFyPAmvWC+OySFv6r7L8PVtgS5x4Aoq9UWfZLI1LfvXK7h
lhpjYHwWgWrfu6ZGNpw3uQEassH47B7VGsc/0MpAHgHKEHw8Wv/yg0KL5blfGi1XVn1vgMHZguOs
ncZD+hd9C9dM2LYUt7dBBKLV7w408S8kT5kwlfZyqa06YRVbbtGbKzVOdMEeW09i6gxGHSwfzlzF
Qyx2rDy+iqmwjKBpxERqQFjX/SI6fj8f/KrSI3JHbC8z0J3jiwMSKiLflqiYB+jPsyx9Q6cqg6ha
3TDffV+GSd5EyyXZH1DsEBq3zCXfiITLirsABj+Wgsz/QstzH5YWkPX1LBOn+tOk2zukDRns4987
rFkibRmyVmDhBUL5/cFNns/KBk/nBpO6kP22NtShF2mFoQKuB0/tbvs1pNCv7J6MZM1RBg13EvJV
/hOJOUTIYBWg/elYp1t1MicJuOvp/96WJy0VVJQ4eSiQkUt6rSVcfXEnhW8pOkEhqtV03VjwvbjM
LY07rVGH094b44SAVjW6bX5P2M7h7uQKb9WxBJNW3oX54bsW4x0bNg0PMsbQ/OieVBPd3oVlx1V7
KUHWLBzesh2AsgqxdN2N8yh5gGdUnD+Xh3kPi9WASpiRwzZ9iuD2FOCrw9J1rkBFvFY3n9gb94Tr
T9MNze4HimrZ+FE5i7w9bFENJH/hqLf77sjGY0SOPnGVnZ+ag/l88emkmKxIJS7WxMInWTQvT+0p
uc3+5XYTgyuTCkwTzp8LQbpmQzmR0FgDA53MWDm3+ZqmEu2Gwyf+tTgXkX61YQHqKdfElVN9bKrc
Ghf2vqaqWsX1k3c32tqavN8gS1Ukk/VbNfbuSkrozCRftIh2zsExGJJr0zRuJ0gztbWCaqkU3XLR
z0i5/NJkAhmsNfF2kG0wHK8Dak671DzlmIiIXaW4CxDL7MFMfT3VaCRnotVxsNV9e6Jx6MJ8QDvG
fZIsYjPX3VfU+HOHmuhTLtYXFJIWN3PSHuq3+WKTwZ/AeKA4MjFGtXeTpJs5YaKiFP1DO6YlKi+9
VXUomvfpFkLuuPVL2wqjEtJ28bLffjzBiMKs7sX29B0VFVvIYvx7NHO+a1GnHwPEOfjGfK/9a1dY
X/7g9g/xHdkU4HuvQRAm7J0X+j+MiOxI+oo+2MIox2vAoYapUrCzAM7FLh8BbXFkvypqNNXg+kN1
Q7t2+muITNwbmhhGZZ6e9CLmUOLhNIaLK65e2ClelpgZuf2Wp9dlcQulZrKENM2V9HEFocuIyiAx
ExeVEJx6DFaHzKvoetgNsSliePS5rvcNgQ4iXzGp+fxmoosTLbGwVis0AD13zGtEI3j6RhDMNhrG
XzqmN+cT59VK/JR4lQk++tHdOIBOIru/81HWbpIV50Q9LV/ufyH6/MrbmYA0Zn8niPAwpbEjEtiW
bJHw5c23SDMWUPZQ3wbvdoV2JUN2JlAhi/G5WZIC4PrUGfiBvHRe0YPYZ4nR9rey+9AZhTYFyELV
GWwfxJua01XxgGjyP9sHn8YANr1MXtbxqjlAHms8SA52YWoIdQ4tH+/gUutzYpirlwMG/GvHDN/K
Eu0rhWW9t74AutETEezNC/ighk64jlgDN4MFokdfkAVOqm4Ub4YBY+9U2JRbykm+taYLDiES57jn
BR4nIf/OkQX+0gVXgrM0w/j9r9ZGBWb3sreutE8kGyv0YlvqmmzPM44nWyrqLt22Wpel4FPbYBuJ
/247WIh94WdOJr2tT3Q4IjXRM+SesXVjhqB276YybD1ymCfR/u1fDfcbbTTPsjMA9wpcTp9P1vrM
9muae9TjFF4S31hZWQxXnURyioAA5RCaM2qxgK6PiZEOzxzbAq9BJAbT5/NYCVoDa/ylmhnqORfJ
KFMcQVYHZ8ZrZyTf75Al6eoeq7e4zQa6Kth1j8tobCcrgGZIb4UXkrxlbkMfxcPPJhCMnClw/yX2
K33zF/bP6jyvoQbAeK4Jj5jugRhA4/KxG754V+4UE8oRAv3VT/TFWdX6SqOjtiDEARqxNa4motvT
NT2AjqdsbAe0QRpF/IsufGT74IHPhzbAXewzYx2Pp7YiZ/6gltBIyQPD0gm+zzbOyigVOJxD7rwp
Bk7Rz1j2+KM+mM90oMG1zyxBwRhRPC6yonl2rhsDkv1qHBKKaDI6W1J0bhKBUxss6jYOUFYNEd4k
NBT74XHHdtKZ6AG7q9LqLl2qnMXM6pf+1LM4omL6OBdTN0McLHYVsz35BdCoXDmoNMS6ci8s9+lB
DcaJLol3B6vWSWEPDShlQa2eY18IQD3ymo9FPwWRbA+ci2bpYGwRE3WVtOaGgqaWUAy3/T3Dq1Yk
6MQevhGbxTm4Zl4eWMo8hfnRZX8BzKhaHuqw3KCFRhDPNm1OgXVPHgUQLujK0llc/qXQXeri3Q3M
+HShAMQn0YMrd2LtgJjSAhXi10xa7Ni/Bw6KmPeMZv6ci0jBv0v0/s0ZazfZRABUGtXiSMUfKJ8c
dvss5pMAoo7a7rmjzRmtCAW8knk33MD3bdngRDL6BsWsYN1ir7MDZ9f7ju3+S3muJQexlAldCZyd
MPBJJJcJqvRrxVkXQtf2jAFAWxKKclpspcq0fwpyZZBcZl9ZxuNQXJX8QeSmEmcRNMBvIzxOwqb0
8gSw0RnMevPg8CL2NLKnkMW9tyyC0FUj8z+M0NGcZim8x+saRr+5E+w3SvoqFRfelYhm0LUXWBhr
TEDOTO+h2ClEK0MfLNVyE1D9rUEYzy4hlEXW9lO4qs1nqtbjrZxrHE7ayNY3oo2oq0Wjw2jEJbrt
HL/lIJpVZcuAz2/JpxpRUe5T7KmMqHHa8kgBfZ28MgCi7a/SweyQ+P7qRV2hd+NHQARFF2yy+SYk
83QM3ENO3E8PRmsXI8/KSVozkirRRwt4yBcsrt0vZSsUJrrXQRZ9axgITHx2T3ikp/jsCr4OAkrD
vtbt8fDElkSrz9VAYeK45xZfw2Haq88+SoTvGwTJPQzdvv674spK6gRRlD9dPZloU482sFqUirTc
TzSpXALkD2+dPVcyR0Pl5sy4TUDiaUjUQgq29aG1DJVY97gpuyO7Vl/mctV/RZyb49DzI0eJHSSn
ccRCoTVTVfNoZV/2W7wXb3FzO9Apf6naX4b03HDeB2mDFAbRCUrAXjdmK8Tz0pVMnD1ipGIdDwKN
kCln0r0+vVKAfJKtNbHpkz4/SuzsxVxPcJokkBXfCe2rKp+5vCaQJNM8bPaZyS1uQ829+chAh9sk
2ynGYmiWjsKhdpqmTL0JB96MQVipHrC8IFc64iynl8i0Za/efyx58duJrl63SB1mBA2nkJSHOpMr
hqCuE4SchkedjODZL4TBxtzxNmnC8GBp1umkeKJ00rzBgyhhE4sNlt5KVHmo2Kmb5sH0wALDrE6d
tNG9NYWyIzIwDfLPeuW5yiRDyEs0ueJcBNXqB8IcKi00Og/kcGZnEEpaGTLbnItgCRQUaDeI9j3P
s7fJ92HL/ehxFPVqqyzp9i/sLhd3mR/ofZQzPu84H0H5qI1wu1efKffLRPkKpJzn/G8v1RAvq9kX
/zwEiu/8siYGG2mm6O8bt+V3BxqMatteaZPvD6WZb4WDulwXZw7YZL3+T4tywXwcgGsu1O9Semcb
IRTjhKdDSAQ6PDfVk7nO41N45q0oCRigykALPM4ViR0WEvMmM89sOMUUbs90S25S+JimyOEmKwrT
hcxSrHYQbK59rVCE/z8OvgR7CytCGAcsFweYedVLf4Mt+H66bpo90GPzTjZ+ZqE+80/RtkSwtFwZ
m+CZG1iAGC+uVrgL5bne4TY3NouYRJj6a9VjdygZ6yuMvHYB99Id2MKZSFYlKU+p1IO5dRl1SBSj
oM7G/ULcKH2p5SXf3d0mqQRlgeExV3VGeNP6QGr3FRPlmRbyHty2RwayCZKeZd+iaxpnV5qEJ5Nq
wu8If3xlr0JeuymlWQ/AmeGSfA16etga1WWW+IA4qkGqfoTKHBZYpOUU0L7jDwE/RhZQ5VcX6KcY
2ig9Vmqo2c+2clHsDWFOUTh+OwaYxSQanjhuFw6ctTrIdpVBw5lCpS6e4ui7F+vvcKsc0qFu3ugq
BHdBdOKiQueAqwa8S28sFOSrRaA/e6hPUqqbocG2ueXuIyEkOFr6ejWRqVNcDtEqximF2H72U+ad
Cz8vi8wSr74qVQLaMWSiysGs0dBG183RoKgcPrw7iwjTWGRnSN34RG+DHP2N53rs6714QLg4xBhk
875hC4RX6AIW/jU2zsejiMwbXZbZxNNnIkys32erHwubT7yVvAk10xKatpGWnzdKTjoyo1Jmr0CL
bkAMXVqa7ZmIxjPQEPM8PmAIyTOmmKCf6QYyb/D4lZmeAmOuquywfQFKI7pskUKz7wc3tLV8d1Dv
JI6qIYNOBTgAluBKrRjoDLNJ1DEAXGHK+8Mgpu4c+zYtELJyzHZ4ZIKgtNrqh4XEX8c2LoIo/cw1
86HJvCw/o3JzXZJenHisSRMHw4TEgK3qqohenip2o8Q1Lme0MzQ13Q6VfAFxF9ZSRD1tSFQmYlut
cwp9OpRFUD25zqSwxbgFvYwLHmG2uthksq6tjuw0HwcCilzZeiKT60OFl299DUgIHn6mXJrJ+WxH
atu91Neu/MtBmiyppShUqv2+Ks5L4LoRBISNJku3sb5JxHOFGeX5KQico/wwcgK3pGu2znCefor3
j5UyeJXGnXv4Vcnlhx6g6iwY1M/UBckppNzNW9VpP9o9Kv+uo+LLedeTBw4Rep5hfcDm8PL7q1Ck
8zvBJMP2X+ht2PIefX9A8gpAeRiglKYT1WjEDJ3xJqTcBnY7+6RYqMjaujsslFTXt0CiVlAIaRlh
mHdqB3ds4mLYOBquipegEeeQ3FSVd92zEUCsRMuCsbYkYtdoqtJaH5x7KXvZxzQNtti9ko2kFAA3
U2ZTcTieVva01CTjI9z9ch7//VzDZGz3Y4sFxIudg7STv1hx6Wv6oVSOu72Qu2ZlDjr1R6jpU0Fy
AvQlsdj8hLubZa761RH28KQrR6XsBLtuul6iR/nDwt3Le6Ht4hx7olGCY5B+6UreVIFZKXS8Era4
xkv66lWu0+woLMmKfoDr/np3hxqoyxMLCBxcP8lUgRBhtkJ9Y0Rllbihs+1NllnLnyQNCPQi27Nl
dP64Q5lhOiOkzFmIhHCm1c9GwCyObSK/Q9RMb87ymvE0EtXdMtGPTCrssdnb63FhvDG+Fi6ikOLd
vn3x8bNj8CveZ/LVVK6yhquEDaK2+jbyVP2ILIjRAB1ttPzpMtG+vw2D1G1OZ0NeoEZwjJdEzM4z
N7y4DElcUf4UJ9bCVBtenBh4mSg/oeUO5OG3HI3nnL2vIRdJgxdJHkHdDp9RfeZUaFljgP37yuPM
inLIEC58MeuZ83GLW2G5p9U81TVizMQuhwYn6HU4SAuTyyYq74lWGSenZUoDsKNNScFw1dkGbYlm
fzsjnnXaT8UAsc2rGPzqv6b7zccS6oFV+WBTlOrT5NE+YybFPm+WLcDDXYLcxl/lSfIzBwKXX3pN
TdmzpDZXd1oP0T4DRtr/DG8wltoq5gJRMj9mpeeyW3myLkTFGZsjWwdt8BunmDZY9g+FPUmkdEgi
4kb2k5piYZjVnQ4XoZ219jk9VrF6JRthr9Kda5dJYRUGu9aLqmYvNeKHgZIGVguKMbUgvexcMJZr
gLGEIg+8yBm6ckhbOsrBHMIDkUMUjrZsBp9WYQ/r2sBecV1diXJriWnH9uNohWSqWSHRBZa0Sibv
IL49WgpLlDi+RFQ842UePoAjjuNwkyH8kqKy+Z8Lo2ZHTEjXaw/I1WyDFXvou52D+w146GHp2U1j
YQN55fUHhCIIMjQR2KrN/Yn23io43Id6cjkmaJCsfbwq6ov8bW+KolC9oY6pUSn1ANv1hHzjZuEc
K0lUyGYDl5LO2EZj/h02geXf0UMonDAzN5isvidYPwm04OCmnYy8Rw09KOO4FVvAa9bHic9qxr33
n5TkAWfIG9zhgWiNNhwPP8+J/q0GNFvzV3cxHI27HG8UwHvXWjd3B1sppkHBYDCbaMoCkfqqpKCl
HMqx53CenaGrVICCMl5fN67PlxPlKruwNqpU6fWhZery508db9AxjPh02gbKSANMGvca/n9qt7Oq
DIyK+cFzpa72uEK38Gwi2WN7mT6R59qEEe3ZEXKlmA6ALyR4UpGWjyp51GwDZiumJ+IAZQ+VjjLD
XGqNffHsIqSbXH90u9juwQUTQMcbqaQPKSGU0fQgdBYrP3hN5ceJaKnQhZPUacQ/hyF6yCCfDF8y
QM/yLFVoDASc8MU6l6XsFfFZsRX+Dzvc6FObklUigvicWu5YrY0W4hrtVpyLKdCl0TgWU07tEGEb
fFl8NCq7b/u56QhaeuYO1cTk7A/2NJVI/7SBvNWRZN7ZkXKtsCKu2NEJ4wVUGV+wWvNsSzEaTlBn
G7Ac48mF5RzQ3I8JuTxyhzY652s93InX6kkvjFaq+pX/m3wam6DJ8sbf9lxI+d1gK0rob1E55XnM
L1pWgtL/zxSkuGvVjDcDsab7b36ZwlJYudB5BPSoTS8EBl3joM1aqSFTr5Z4I0mh+u6xVkbUfLoF
UEpXkeqTspV5WHF3P7j5ttF/aRfLTFjwWe74wAYKhxlgAVkV0JReLxpFAl1ujRPvKCKa2bypzWpJ
XXRdeGsDMvJCzQPVOdEPWtas0BsIX3D1SnMXaF3QVgEU3N2Ky6anQR7eDYXG4kntLMXyXsi9xzB4
dD82YfRvJmtXYqsLpLswxpI+oHwbKls1OjOvXCeSL+pFaEDrgDDsz5rtHvLCUzK6N6uY5SG57VKO
gxodUD2pKuFdD9H87qMG/t7L1tjymQkt5VhqIDAEjsOMBT4xgHE4kWcJqBUH6Jmhqs8fQucD+Ury
n7kpy7Ljm+L4Il03txZXWWIZ7LHiFlkAY7ZDFZmMO0p7Eno0fwZsO0WdC/eXcojmp+KPnkU0ERS3
3csQoNADMyC3Kxp4olM1ei8v1am97ZM7+0zCJqOap5NFFmb8xqii9h42HR/V4q+K/u3KHO/lzJ4c
7aMgz8mRyf0W8S8TEgJPa0RaNFZABI3aqwFYjxzy1spv+tWBBdpat/MWJpVdgVPfClYRHKOOgbP0
sR/CGT2fVllUJeeAKievkbBWzOGmKeuvGm6JOP39VWNe05tO5FUZINTHddOXAhh19+hT/uwhd0FU
JdhCMbsRk9O4JCC4459cAsb2eRTC1omJ6jT64PTBDa225P9GJqppxU0+rdN+vu90VgmFLcMGOM06
hGuevafeebjit1KWNRjxGDh1QwdgUluf49KmykbGbYm3MkyCm+qzLdOvdPC4J3vSGXzQZX18tXY+
RHdVrEPrXbvOn3VwwYUOy0wfPnbO+d//hHjbSKZjjhvNEoJhxjDJpT0tiiOwAGC4PVrMKCbJ4Grd
r/WMttf55zmI/fObLTOE6R+MixMD95xE9/hOfwaaACGZTtmTcdqVh1oLq+ddTTmMfGknsBrv33pZ
zX7Es7OWSr1+VohSuVv3Ytslrq4M4Go3XjukDmUxVDUq2T8yn/rGNrTcnihrmSVurQfQ03iJXJCU
xBumkYR34T7uivxBflIDz59xk1ecrf2Rcq3aqNputgyhxswB4JoFf/F+xM694pXuw37cSnHVqX49
rjPCwzsVIF8X420JhxjpAnP4Rcz0ZfonZNooZKeEKJaxxdcuR/TBCXaUwD5nSqHNNd454sQ6srRd
Gdj/lt4Gv+ZqR8pYgDX9Jwv/r/Cv7YC+zYwMYZma75A/15Ocr2U6DWSVyDiLkuJRCBCczClcAx6D
4lfRS2Ucmvcg1pvC0+/aGGS5ZPCyDcvA78EAe2aXYhZlOoiQutiJx7b3Qeq2IVhIrdTkwo+qLfTN
xgFYlyODp4ByeW2aF3hUZ1L3q285u5QWB1DDOuPmAlaLt+WM+bS4EoP9+VLJWYHPAS39j6Iw6LqD
3YpEehH/7IbkHqDi4kueAXP6vNelyJqf2RxdHzHMyIz+Gz7Lii0xEzd3Y0Zkk9d7HTGnXan2kMvE
sCjbr7JFwDmW/sMADBWXNidHAEHqSuKxA/ezzGo75D5KmS0F0kYdrp6I1YzH1wCELqUPnBytezMp
PELfUVcdlNzTIFdy0Zxa31FQzDCF/u2cp5bJwgoWuXQ94KGX0wXsZ/VXfqfnjrZd5RKvPWHm01I9
+jdMUPIBQz3ATJ+f0ml0vzFYkZqoHO7UhrxJ/PXLQsZcAGCMMiObLANiXB9sHWTvBkKKofEpCe9h
J9rFU6keEHcE435aGpRYa58ymwdVs/U1Lj3ELEAV0y5QwiBsafE1tp5ga9+nL7eUySsGXCLHOydR
gAUzR/a4hcx5hQIIQ01Vi7RahUJQoXKcLNWuMRcbCFnzNayeAH7JBJyqM8T6N2XtFfTpa8y6r+0F
SggvyqID6Cm1nHempKrh/K0NAqyTCg37fUzGsv+OpwpciiN1nowHrSNRn7/93JNQ/SXtVtA3d2v7
zbUlgO6W1PN2FTJ3A0JU22OGVvuxJGUcgSswKyS2jfeCgnMJQ3zaJbcSnAH1FBo/UUAvzw5u+fIA
bbz55Fu5fyFBKDBNFH9RpUiRHDlq/bJ2jfEzbfnWi8jVlD4Y5GVAou7lYG5ysQCA+lalUqRhhauh
bLxU7X/AQ3wy+Fvi2YWT0kA9eQUId9MP19O592S8DThqBcqntRa/P2pGu0G2yORknjxw9r11mPAZ
OG8K6ST0vvQCVnwlD2vOTtxyvSeAdnKSAK0TDA==
`protect end_protected

