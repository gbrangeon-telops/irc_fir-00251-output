

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PFFltKdLY0A82yxFqahMaWdN+zxj5kThYAcsDyz3A2vhpKKQpGJvV8/AkpYYPyltKlIzJB6Md9uF
AN2ca05J0g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
obdm7XtHPDQGZMrK3kNZKnRt8ypfk4aZ9VtSDpnSwNdbgwrFg4uylDkc4YjBW8BFR32vEdXmCKFe
3L1bSMhXRkPXZ88hMJlBty0IcmSYNatn3RV9VG9yYtXM73zMkJ4NIx7KoDtvOCnGQpHNAJTknAv6
BNEUXajqHzh/vB/QNBQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nx2eU410BtrBCSzpvDl9pNpIplyp0nHGgzB9LvwnXgdhN5HNF/YNjnH8WXRfWZhIT380E9zFeNz1
cIYhUxogcuyFP2sgar0PDv645GG14wyLd7prd/d1E3Ur29iNukQkz59OjXTEIN/U9Gy3hPt+oLVA
TwpP0P8RgeQqCkJY93IlvPGfZ/yeDQHrxDZUMFMxHHI51HM/LG6Y5RjcVEJMkX5GTsC4gSd5fEHc
DWDREOSmqmG5Gmciy22xZEiB1SI044vcLqlJadcUhINRbAw0576LfZrf0pjCGq0s1+nEKeJm9MeA
baA5VHd6hhXLwLD9jRkKDvFp76mdZ8cpvFpcXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
my8iGpxybuJuMik3+8MRqWVv3aAmCE4oY3Ij0YIUQTpme5jJv8e5DOlNoLmgXWhUlepBCUyZ1Ysj
JGlFKQ8MBs9R5aa1TLi8cCVfI579Nm4AO6VpackDfb6c5/BXCbiBb8XeC9Q6z0hKyH6xYDDC0Z7w
m1jdROr8ONcmGBJr57g=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pEGUMbCVqav8XqUNf0y2o1L56804gb2pssAnfqbrEzVo5CXZ9MmyISfyPG7HY7huXkJ9tWIeWtYt
bUG1XTbOUAj3uDqhigkZ4KnTE/68izmD5rgLlGDQ1sI7w5GLUgtjCBINeZsiQZ8IbdNK2b2sCu2x
1k1tcyPPvRv3myvuFaOhmiYYyCNc8F9T3cW6mq34yHrMb8GcN1rGLFkL16mdIcoRSSN9znhYYcLe
21llq9uuuR5MD7mOGEYx4bKUQGVdPOHLC411Ms5bCd0IbhTC0qWispRkmO0D1uXT6TguY5Z6gKTw
vMvXdJYpwStmSqzikX3kYI1zljpfWHQ7HMzzTQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 66352)
`protect data_block
Tp6/UrZQbmeYSyRKvaQYlcae9BotFy9FlHUFCCqO/6TKBEMspe9cNKATk+Ni1SA5BkbJkRJ/lHxi
BBTq4tqdVGY+rTmti/4xO5dJFGtaKxeDga3dDlvok0FxrKLnbSP9aMHLEs+B1gcfCkbn2RAWhdPS
nkPRpp/SA+6eQJETJptKWpRUhXecf5SRC3r69Xhez9fAoQlGpDkVcabzIFu0Iyj2jo4xNMX4G0ze
qrnQnEkSQVGP1z45bljRRF7m4CDKqq2Ml3R0V0/N1Gs39ksV32MCpaqyorPt4EmTm8tzOxTp3h6e
uKJxppjckhGfFjujPYvl8PPu7pdVDW9XBT3HjPih7KUZdZxpI3f44ZPn6zxQCwQ8gwZU0igmjBtY
TEr8atj1QQ6r/9cqNtIcB/L5X8VceJpwvq8kUsDJQsnu+qzVE5nCTB5rAIvnVItCiOSMgWbjxX6D
HO+017XS6v3SQ56ple4PenkYZo2fCUSy7saNL0lnGDvfRiKCVEmznWpc4VuelLS4GUeVu61tXAoO
P+WFU3G2zPUEqpvx0h4+F9HaTTgso66WHMJi+l4FZueOe7Wl7gdCmIOZ9mFkPU1P1pnidQIuhBrc
h77CnbZwrGAmOGkArdBraXPQScojYwvXWOYu4KaQ2ZSc13qXvEZYhfXJvCd4FV3ermutxEnqMvr7
eWYCpU1HpnapfTZ4FRf7b4q1YhGuUmhe6KEMWkt9lcgtSHeQgAL3ik3dJSUzkbJZVWRcck8REawn
jpTdu+nFUzha3RFD8MQekkbddfNQGc0d54OIgCyZsdF3svQdqDtXugHyhvk8eqCztkHo2vwCOQmv
FNJWZjH2JckJc1umV01WPi29XL7A6/nuyf6RSSnabf5tMeg0Xgg9hv2GJtRapYExPsFv8/nZcxkU
oou8P+lRMaXZcyd5KA49e4rKwIrsmRoBOhcUMfDAMiMs2otM2w0Uw2+eepnGPLIi/rTvkHQRO1Vk
GUF55NLZC0DNC7A0qdPOnUdTMo0bdS+BiZgWrLqRVRA1GML1lRC62V7HvdMQjUBXt/a2VaCwccoC
5JIUZEKBxvl+HxfQClRbgZLZz329N0H6Ca93Hin8M/vyD0iUDzcvay0PUhjbTzQ/ioC78vie011O
rvpnNXQkdtYQewE6EoEtJ7gPXhgMLejIrmmev5EcmZ0F9BVPQnWqKz0Sq4ypqn/+XhmANYMthjAR
z6NK8bdmbBmoNG22UGQYbBxyqxpw0fay5t8nDWcO5yeIqYua1bZUUx554aA/MVrGRJ9YQ779yokj
Wv8CH+YZX8nBkBN8/WCWDCf56C4t/LyXuBGs+h4n5dFQdW9GHo6lsSoxbIR3kH8foVq2H1LxgO3I
dmyYFXvzd5BKMDwOhleVETNqYe55qyvq6ZVTJdeWgQClHcc6ZUdwRm3vLNZ9ya60CgwLr3ADxuAI
zOZAxMHOMv9uuPqtW2U233TbxX34tTTlDOt4KypNTDfXyrajQjf4pFyUIWRHTiEuvWAygO5lqReA
N4UdhiIrsaS4fOTk2pYDY30Jbf2/p5kZerttDwAybW0MqX7DS6L0dmwiS4h3VF7Uw3PZr6CZ8zTn
vM2cCh3PoZ8WutD033aDd4hIsZUt9459EP2/XMRyahlYNOCV0P7jsQvxGGGlyr0M0c1ep4d4QoXr
+Fw4OoQ18wMrQ3u7zAUU/BxyWpWxTiTmRXw3CPYMrVSlM8lhsxjeGI4FSzlCR+8NxlPVJsrOoG55
Qk+7Vs8tiOQJ+xOmdqwCTvnZsf1q8t/3xPYUtPZZsmr39GAAFbz1rmlL16FA/129HGLG+knKS+9P
8l52t9mLV2xMiLz+wDObo2xVhyJX2z0CpsP7wZo42LpOGcKF9I8wdPSOooKF5KqXTokQcca59umn
vRD2y44yq0mBGURpDE4uUBmsGh8hmkUoPX3uOXOjT5vL3heFTsI8mHDOkt9J71hSc+gpkdF9sYj3
rtcDBE0uLZ9maXjs6Qh6vTuFFvviUBB22nSgdg1nWtduyLUxvStz4tHCbmBjbFfY4jpCJ/MVy59t
M05ccoaEBY+cyjSL7gVuqKQQjEBwanhmIkQ7ws2EN7ytAbqDjPcwAoUverVNjr8Eqb7mAYsPSKGv
XxWdwzM6dyiHVTHvY/pl8gwj9xZ71YOHEIIQFowGYSwAYfc6ZmEhAF8QaMh9UrUoQdjjMK+EMjkp
PxIas3tOMR0s/9EYF92DbPOn8f8+ayhiBV6t9oXqO5Q7A3Lw3mT/8rZBPlk3UpUXWR0Ixa4qvwuH
NndL0uSucBuo5U+z8adizT8kxtRzxbBMVKbMvzfh8zapsk0kfp8/eGnRN+KD4YCZAufOgyRyIjOi
CYllQ9Z/LBvvN9pDP5xOFPLGovNiLBd6Mwg/uTEO43/kxTWGCsQxh9f1Al4D33SzV+pl0g6cKNcs
faYkbkXF//hlrk5RypflUBFcjyYIQYkseLMj22FBUa4EblrQIRIDca4N0thApkw4Ykbq4a7PC/u8
Z/F9UtoCauSuEaYMqwr0txqdFFGzFLGIX9EMH1B2I1nJsqbzTLnKbzNa4MqpFl+ge+k3tYh/wX9U
gptNpdUbodM6PqH39PLT14UdNFzHearTzAp3LUy6sYmnnj1e/JxN+vKSARZJzb3Zm09iN+pkVXOq
zKNMRm2JfM7JKRq1r5hNxUcr7InDmNdKlO/I6MdfpY3MWcmGe6ANquxZCKJEqKawi9i/G5Bk6x2e
TcUdh4V60XVcD7FrFGjif8mTK8xjrzMGKMX4xrGIB1eZZBtem5MNnwB3vyJI/NDOP4QRtUBSMDul
sm9QTgQ5yiqB09UlpBEsmnBIY+po1+MYILuhTbHmqoePC3IcEAsP5Q3VaJIzdOmJXWjz+1pqAhn0
wVFMggv7h1iGA+NvENViGg/ugUf4ykHuvKoE4laWpWRy45hjZNs1AvUgsUzElrU2s9duqN6JU3rt
wg+XU9+WUUvEhd3d2yEv0g20WFo2uF6BBXzsfWLIxHQ4chgD6lAMyeTCK6+M0fUu/RtKsCc8Jbul
AYcpV68q0+FkJvo/57eFuyGePfFzz5KTcUgg5R4EqHSld3f57e3VvWVLxZuicq48QcNZDdsFfxvH
03oxYKPXXHgCCpreedf7MQZVHXiFv9zhqGulHmp+cFzJm9aBOgGMaF2sItB/oiyECvGXdrqbhGk9
YvGRd0hODTBeGGmZ/Kr7F7fiodsU5XhfJJfM3oOY6JsLEucrOtBHHbrkRQbJsJ0mxoqCDPPKCPuG
7B9UDXG1DBdMgISFeJdvE1D+Kk/llSHghWe8JDfcNX0r5QvUl1tbRc+2YNEhyaJJb37WO3hV6BcN
n6HTo1QN1jg7NautGu5WU6qgYzMQSZo+DpqMsrp2aqVty2knyJLFC1m3eZtZry7tCHT5I/K+Pp39
QfFvxsMmQQRZeixT2A1Rs9uSuM+FyGP0yvUjq5lSIrd5ypGDwZCIwSAC0Rq8MwC8/Q+0uX/mTVOX
0vbqFEmA48srVjl/k7z/RVUF/VXIHVWmSpR91nyU+uPnnI7Y6u3dyGGL3axeXGdaUkVlRpU3Ov5U
8HhteJwiVWPWR9T9yh0UsyG1UVQlK1q9/3Me8ANMQJuO15S6HjU+EWcWQup4PHePGh5ngECNsSzK
JDDIAeBjiOVeRaczLaDbZtvbd9JiDHCseLOPu+no3/8Y6hargYgPENRUKqYoL5UM22q83q4mVERh
l1Fe1bS93DPJz3Dgy8HM+GuTm9BmAWGR6L6ZMCVjU7r5M2hy7RVgmi4PnRjRDTpkmlbKAV+b65Ds
6I+wHc2uVeZbCRsnaKJByOKXDmW0ZMf2G1sm4ZgOZf27RouLd/an3oTdIbwurRbzn4pSjOSWzUHK
LciBvVPLWQ4QoReclEmhu0sg2O2Vse3E9ezRqLjZAbmObMnjtI91ywm3DACeKFkGoxWe6zhJ7H/K
iaSH183BhCJPsxOtPQBjyAvzup8VP4VEhMV2+nF/Fhw4Xgvh9zVlbsUn+vjuwyL8yYhibcWGFdOo
wBOV6NBUe5KvVkualyVOEJQnt8Dcwt6UK9GV74qdtVc0p5yQ1PtAhK0oZikH7sYlGVh0iBQhwTBG
z+xcvLmoXb2uXgxR9vZFfFBig9XChqDAQuW58rK+jjrliLXxyFrlNoE7HpuMIlC5D2QZxrUpB+Gg
HepCJzgDwKfbJflYvHQ2/LMnpnTTyqkfFtmmH5Ci/QLgkV3Gd58y8USBvxgkcEFv8g+SDMZt4f4J
LNKcYj+kg8bIymcD9ZwuGzMXSPoePiZoohx9PUTwPFihfd7GWGjzYy6EusXayI0XnKFWuIAZDdp5
KM7rlL+4F9GlHsADtsjpNwuxMlaJLA65oD+2sdAb1cL3XFaZDgnk5NpCf0qVrdtlWk8k5k5CJB7A
sVfEGrk16sm7ha1bHXGQUmuJ78LNsczMjYaNijE4mt6gGTOfcXz3kFHEfurzjx3XUB6GD/e2Fu0D
8MP6L+PLloVIfxrU+rOo23Pabyd4phAEpRbNS409hx9TWg2+zESrPED9h0+jLGoAYNnXCBcAe7RB
KGoxmTJxesFqbD2hHBggQkF159tJFtrJEBCaTlkxxa0x8kiE8IRWsy1X4SwikTbSDf0qzrp3ML2j
QWgnmgl1BCoZe7doUNSYNl6JgNplr2NjHw1y1hdMUb3zaTPKx7pGNB3HCvf4aAfM6OaZ7dHylfFp
g8NOYlq9NUyckbzYU4WPZqFlHm/I+1JmBfRIzJPbjUB13N57aj04Xbg1qzt+jUSfdmUR+oiz4Rjr
ezR9liocQISgFmkv4nlV6XJ0u3hZFatuWjv63wwyRZJPpfzKbhE1dPlLrOWy2+1jl+p6KXF+q83p
/RJKSrErGfrkF/jhIiC+xLKeeZR1GD/n3ymVE2tabPRttyhD8m5U22ca6uVi4YJET7sJYzgF/94H
pcWIyarkgeM3zWPoxZrWhunC7GxtaxV87wGF2BH9S2F1zCCoeYG2YUfOhtPnZpWU+4nlRa/HORh/
HVZbqcIjeqX7jxkNRJkI00XjIxcbCQRj3EYr44ObjyJzuiUrtxYVQ7Rzk1UA8CvbJTv/TSIHiD4x
prxcAGtJ0SJDO6iQmoOSc+iW9faZ2PHlQX8NhzctYmITvfYxhJ4101ty8j68D4IDhPFD/J3H72h0
EhL4M+m4qmubphJlWK/We9hkq6l+E6gW/OeMFreHHcqPtw4Ov6C+wwHlwZCM7410FYCfUsbUJ3yD
yNQ33vNkHeanoQpvGZSFmW9sU0OVNRlKns7sF6fqLmzDthcvqx94JRgy6eSUXDAb4TEbrE/JsLVX
uj9C/2PqJ6JHwx9oWZICJMenr549diVtF2sUbRz+UL1oxOWOHZdb1EbStgaS+VdC7n0fa5gmwZcW
a5cG8j78K3NDi9UEIwnQDFnrQzhXwh+ExkgyWsXQniIEtIcyD0sS0hybquD+Uqnc9f1YwtiZi9BB
UT85PVqDL8HrYknWHz0N+LurJ7ZRl8DoilrDfxkgqkuw0ty9vDzqmUQ7goXpJ6R9gxjsoyXTTxjx
6E7L2BE1uJ4uUDH93AeF/yAIcaQt4txlVjYMA2l30NSEiITlBZuxf5cqCGl6R+LS93PNhGLia93n
8RStHPH58oK0Hd98hmT+Im28oNE6ioNicJ094QnVuVijEau2qVsrCS/69v5qYsk9HtScCzzFQbmS
Zx8LkBo9VC3csMYFNaBH/0mdzM9ukdC5VuhcTRfnxSc4mRmzPorLDR3+V1aSgFDN97MDJId9S05t
vRXuBnIBVJ67ANWxGw3Dly+wMIkVbOv6Usg2TZ0jEOVbOUdNlfXcwbBmYim+du+lmsHV8rHuXvML
+Qqldr7jbeKUb++Md48nBO21Zba6LPzPZaDHDgd6Vne24KjY0FOhFgzoGcYerYzzCPBEGwZ+r0FY
aHnT9P4Cv9w1KUWF9eJJux3y/QRynbZ3suXu1ZNB9MfHzuyN2tfCzp1jkLr45v8IpQmHWn5oAlU+
8JD//bvnAtU3+gwGRNIA911uLv2ToMHAP1sGi4rCut1WmdqCa6e1iBTnAlog4OIXurfSCpiWSpOT
0JV2vcYCkIOLIzdlMZkhuhgJfwqMlHJNTTMTax9uF3Qmqtyebzd3slZhzwDiNCXufqGjdqYS/w8P
afD+BEOB722LqCEn7ITT5TytMk/ubHh5zyzlVwW0nzVc9bda+NQ0+aM6dpgP/+9NCvN7YS+tSgD2
WiI4IIUKAthUtQHogqKDj5jwQYsa9+KSFaQIbWcNz81fjPFBwoncsBxnMh51C2R88ILNq7N1Xi8r
986EVl4pA3rvn4ATw+uLC0aTODyVrbZwUcFG7/bRKI9UN+QclBEcZ8QKZaxRDV8xa1hRm9C3E+J2
ClnJx0vsOEVTKnF2ODpOogcfDdKUgHgpMeYncuhMll4N7+fiptw3FkAp8PNgbHnH1xoZ+qR0Jgms
OogeOzQ13FpyEWXhvFg68ai29HURKeSG403ABxVdeiOn8AAns9mVSbJiWh2VbyNyOSWm8cHC5sEP
7tydvcrjbi1YSWPSqRmYXhqYLhh+Y5mAWPWXID6mgTcakYFnuXQFKQ2XncwijzorCAIGeQRx9fbE
DD30CIpIwg86ei9l5RVl0AaZl+3xIls9L1rvpjFbVhmroSxNPn2bNA/H65OlOySEcTgDWbtfOpPY
isqSbbT5wVmAVYu96Gw9stFXbXrJiXm3VqqxWndcZj2FQJOCvwySPSMVgnjLzfm3wxt+OXRtFIpd
D+e6zxbr1QozkcW3yFDndzC+1cFB5ON+vzlSo6ruoNzoHOSaLA7/IjV9JgWE5BvVLyo94GJxPM6r
mEdB4U9ig+p7dAByvrSuLXu8zIm7xse/bHXcZsYlHYacl6YYuSwoJS7DaS8ScLbMkxs60zJdjfVs
aunTlfNV8n7Pjon/ZzAADTht1Yx8RNt0H+YTaX4+8DyCxZ9XGZ19mhjA+qfS0gAL8cJdVO4dDYeb
/0j4Yx03bewA25XiZPevXM0vuL6C8WeKi3fR0GSNquXw/4YqEpp30ieZX+DECkXZFXuecQcenR8S
zkeWF8ZF5ptSdTj5DsW6qt36HWekBNjWNkkqwFB9fjKPn64TdsTeoCpNeQihz3/Yr6dggWxlffeu
ZPa80i5RXMObQ4MEAK425ieVoeg208KjI6U0w6qRX3TfWIDfZl1LfJ5rlVqxCKi9EzCvbxMdMP4r
rN3RQdoqGdFQmDHbICwtaivPcVjSZ+hgXepaTTPEt3CBxlNC4WJdhH0M+wg+RatB3ySAl9/lGxeX
zLELasWYfBWilUT/YnlwJK3Pek1WfuuVhTFIY3yfX0aI1ZtE9qcbgoM7MXMiwyiJDPeDL1Sj90Fo
4ivgNmU7SY8zNK1EhmvTFMFN56uDb10HjMD9y0UjMCmXsawaPNv0o4Bk5qO4JSCnmrWmVOBY1Ufq
NRCS6FD3l2LVGVkU+RodWg2PhNixFbUqh5d1IfF5lMSPQC8mSg5p65sixe0yyyl/D0uDbDsrS04Z
HzV7nX8FCXVN/3coMtoieXBamcV3EdrBFxuUnXN4jaLQlkpyKyGXz9SYGiX/L9RDmRuF3QmdFr1q
7kbSV0U6XEGUIqktVqMcoWAEhCAuxIwDU9gD1h9rBR4uF+nu7nnjvOVwG87fh0nt47S+PXYLybfn
vvurugYHYT9GqXFxihlDVRHpwR7Bxj+SvHcUBqslFkAlBkSO8uXmTqxFXyYtUx4b5oW9KAOhQeRi
1MmKV/LOdNFgUPLTjhT7Bx9NqLvrWWcRa1q0RVNaS5rwG6ZaMIjLwWdR47M6nC66jBu6ufQkLZHh
tn+lR7OwujpaeU04px6q86ORbwj/vk//UJ5z7Of4QqfwbTMtDsnkqjyr1ygi15bcc2tO9GxUBH3T
sSNpvBZm8i3TXuUpWSCbkWZ5xhlGB1G+mFLchW7OM9qBwSz2FV0nZoTrQBuD21EDa8diqH6C83OR
VPTV+mjLpPXo2oUT2tCq51d1HZfdwjc03Q0mqtM6w9NRCkKt1cyz6mRPw4pR+0BC58An/0hD319H
nfBL4dBn2X9tee6v0Ia1ngBkv2X2DOQtkCkAubHP8hUgKYYW7lXN9pjtohhhmoOZl/uPvKfYLpSx
Q/t1oSgXO8T0B4r3V8FcgDjJufCRIJiNhN31XE3FlvWvp3iaWNDBDx2Np4jH6VG4l4JsyAe3DZH7
w89LZUp07cboHtAJ3qOLIzYnMAh87KcYx2OtSlpIBm0ig+Q8relaeu6hpfCIwTMoa+YIKktq9Ca+
GGJlKo65l1I6ZukV/CAWC4sJTUIDC1YdIvyoMWcTWEd0B3qc82n8yFXQJySPCmXzSPZXWN1jH7t6
F9V3wahZq9QDUFR+pM9odvdRKSqZJ7oqdE8ymWmNy8Rt+dlai9SXSCyISyw6Hv8txFf7QkpBtUxe
nMJeYVXfmKrIu6P4BsQifx+00KnRlHZf18yco8n6yeJF8WoQHHtwqjjGPbAyAwwRn1FAe/u0axnR
EKrIT4YbdvMAkxRqTRdUpmkPVyoVw6zskvRXfGIcwx63aTCeN5wH8cLJ9wdXQh6BXYC0LAB6ZxxO
URpn4C9HKjMzeclRIdFLiLlp8UnbMZ9sjGUVb5z/FSLgCuZteA3uQyxd0hDxf3P+u1KHSrfxoKIr
xVAhCwF6zKNmu4i/vBlEiccVuV59lbed2par9ukEMTW7jrgaBL623sBa55TjoqoBsJ7kVTZr8org
1gpl6DHUB5wt0E+MlmWAffYRjbAg/0mKmZ5RA1TVhHnrZ08H1LKTKeTKD9MovMJLsZC/S26hEY2c
NBKSFlMab9hsS49WifKj6+/WOFaAKoe7sYT/3y0Xiibq+We+KoovE6Bp/5GvXJG3XlZd0rxtSjUb
3m/MxikRReIHszrCDsw0W4S1Tv9ZdnE44Oa4qZYJuOkUefjZ5uI6xhqMnpOonz+mM4StUpbQFxjn
wGwNJD1wtq36+32jl4agMjYx4su3YGi1ODTZs48WWETJAYgw7yLzxmePtHbFhvcxjlUTbraInngG
0uRFBbMh7u7K5DUP0lf7kC9d7g1F21HvAeve0jpi6/s/33Kl/JzXylX0llISG1acJ9JJA7TcUjbM
4hTgnNPSwJLQKn27sRYFZ75DXyGQc2q41MKwz4knj6bBzOW5qqWjAqguhyTOrHmmPQhGnclgsFIx
lMQpiHU00PSStbmzYJTqhzKaPCPZvkRbEsTpyr/oumrOh+MsAMxzOhHJnoCXUjTGSt7Iybv34ixG
Qn6kobqOm1lb0OoNrLmZDL783JDwZ/x0FOoRhNrrmCpsPC/zHChh2FodGdlMNTWGV3LBlyrs6kGL
6q/Z09ATbAWGvLtQ2qdAte3bKomoUl1BdT7Pq+BQAhgbOMhiAvdKE0WZx6G61v5J2xYKfb/L7KxM
7nDguidT6hrMl3i4RT8rPQ6pgs2nCGnM7ew4RuWshZNXGwhb+ZpSjjBnkhsXh/kdEL1wxqWbR6BN
0hD8r6xYUnMZIyHQWzWAuyHaLJ4khFMObS63OTOEfh+qlLeGH1FuWM+Os2i0PHEezMWxFKOPa0wv
ZHEqCbObdU9F+DnK/JP31NV7qIp4vZzbtBEjpRyPjbw5K374vc+7j/FJiStdW6F5zb4ftFie98FE
xt1+9FS7WSkPIOKV/qQ4tcTuMpyQ4v6AUnWYU6wg27gsHWVYJsSX6ytMdQS8vtN8WOJRh2jAA620
Za4w7vwDslJ4r3cAeF+EetIBbvXbWJ9JJWokediMzxuRF+Or/8M81dHAFmtw8xU2+nTWhbhmefd8
Ji/e1THG4CWLwIolTlB9/iRB13ol8VG6hv0ZcxCWKwAyeOl9mGOI3MNIHuT0ti6npTYFipIni/w+
MUxLw1GtJI01iCfdhFdF9H7fLSluCFyoWiUmzGL4B1Mn/l6pPXzPB5pMBfpw5xhMHvi5NsrwXkUw
uQ3gmZ/yENMSEfC4p4BYMIRQElBYboVPQbl4EsxTEjNxaAG0OpeeB9csW2izW1+pYkqmzJAOXk04
+MJSqlunxLjNezKhafQI65wu+uWRnRph8Kf5r2i6hvfQBQV1G6SJSKJnPn20qT1eThtHomtuo0Gj
iaE/c9gHLx6U2o7U/kl75Hq8WonDLJI143/WGgWJJOQ+hlx/C2yi8bJqMc7ApMsh3ShATxyoIftN
to3iamdmS8y2xZDyxOJcUYYGvTATrB/khgyZY7kVt21OLa+cqBVHDJKV7Bql3uw3ve061ybM94qg
gY/A34jmXEtLDxCpecaVoMhZvw4PQ0IHD2k5cc/9P1hzG4UJ+799h0tjz937y9JCDa//8JHuZL8g
BAWOZTJMQ3A3lGnxL8AtcGrbunwOj70ouUakb4KXnTeip/NPK6BEUSP9Msmc/cbmNitv89nWTTHg
ymR7YlFy7E/rGf9P/VOFbccVtqdSUDUETQUrWvW7bF/zZcUV0eJDaapqaS+KemgRhSdkTgtLI3Sj
EAPGxD9maUdI2loSwFwDNHhP7VTxqRDAd3fT+iPrK+tScFMHzTYlSVpY/1roZoBplOS1uDhzlgc5
FjT0WJVbqYN7gNzHk7nlz2Yq0Y5w4dG5WfydpGOaiE2rnIZvVlt/FWVvzVm8YqQKUbRACO7eo0iT
uu5aCTEVmTp4dmqN8IEni7S+vXxZmudQPJBA8iLEDD4tryYGQaeWJA0DOtgjwc/oHYwMif/lAE5O
tLl8/WdhCICi5VoLtQwFmLX4a+RasW4EKpt0BqKq8EK9IVyU/QhzgKkZE3HiD4RilH+LH8P4uRoY
eYPBUsYzmNg+wMf28Que6zRW5fMaDOaYNtt9bpExImtpWOJYhMQHC6rWsQZMcLp2Q8CJYzpESUrg
HtklzgkeNLRvr1yfN3iFNr5NPgPKOouBczQu64GPULj7NTfx3j49JWjD6PYbzZNw3h1xASOv8as9
IBsrKCbZi+pv3JKVEg6RuJP3zB4DmIaoqmD2XKNLHcA8w/XSayyKQ+EPmM6z2XJc6CI2oA34H5zJ
urj3zKSEmLBGZQOIgjOjfUdslJ0o1UePq00gJOXNrAmMK9SkJy7xOwR2C2eJ035IVvUIw+Vm34BL
7qvj8+2hofAAcDMRwhnGo2PvD6IiXyFL4XnG9CH/7RPVmZM7gg+ndNQiUxfYdq5Ebk3gRiB6YULr
vFez96scbM0oJKmSct6KBMsqS7MvfQhAMG+1p1BYpMHNteUUU3N8YnpKeZWSOjV/JTamKQtQj2SP
UnADyAq7vPKpH/w/QOOfa3h30ZrKBbxZLNgpf7v9m0n7xN7iqV/MM6A+bDAD9X5ZgywMS6hNWber
KryjMr7ZTcfrHssqqbWCbTzvd757dlVuwwAUNmwr51BYzSoTf7f5jOzY9E3CbMeRcSSfWLHyin3Q
5npTeLrR24jb0KdG2MD5giitro2Efbl4D3JurNLJdl4xBeqCCTAUo4+AlBUUKYCw/M2yA57gaM0j
/jRMxnVao9V/2aZWfa+HxxW+nG2sdZ/UtITdfiCnGu+X3VpA+1KsrNu4I1hIxW7pPq294BiHX6+C
zOX+hJCNGjGEHzcFW7hZq54OUiL4Jf01vu9wtuF8+Z6K7FL8VuDQLxbwIhUC2ZZp32gLfGyBEN/s
eVkLWVA0n0t+/SBPrYjVztDO91IpgTNRIfwvawdcfkTCulObNmDI/7Br3oE2PUs/LEG1VJ4ayu3A
IISgU1J7U7chJ7FSEaOmFiGDGCEn5rjFYu5RMRqNvixrQUiLwueVap0j+dUmk2WLCT8SV7znYU5E
brj2xrLoELgEvaVxNx4NsBXzVnH3V8V+TvlpIWZCBMCQem8sr/43tGk7SkixAY035yUiCEoCSbd8
P2lncR4pGbhg1hR/DY/u3Q0ums2PwGH4oSZf0ssEMJUtzvOWX/Npdm/G/DDfY7bgYCuccqhgMTap
azt4CoYw81+Sfsv5lRi9kWGs40VPp9W0ZoL9I986e4AVkWrfzH3DKVd2eRvNPgXd6L2hfMyIwOdg
T0oId5bub7kO7cx1myxs5XwfXRqlNQkHy685ZX316tgOACYc/aCXRpUmD1MGY5P/pQSxlr/9mxu6
nmcZjnA2K0PhauiJCxuKv88UzsDnYqBO7FrLQ4YTnPmnTqNKjbUM12MTS5aCnoiQDWKxUUEQYfTK
GQJhH44toJTi4k5RTB5xMaXVvHjdiu+lYKQ5yXTMjRC+DkbyAAuhBQUA4OkcnwH0HejFfVYtWM5A
Lkxci650tAJ2/8xHmRdNYRb10lG0v6sf3QIH0JztDreeb/2NhguVFCIOu9AhmSF0+tHyhxQ8jTHA
WpBbzl7vsTH3xuJ41YqVnW69pxocxY2qdqHyNjuLz9Zi3p/sBsNhynMZeW9rsL01kNCFQMU8fn0J
R9rVWSuSHR3iDDuvStuhS0NeRifPffHvqlaj7TDJBeC6jE3VP/bF/mgsNh8UVEYM6X+LCNQtvL/4
EdMMMx2QzLmED85R0Cmz/niQZ4Gg/DI/NYddOrWtzLzF3PRFXYSkNk0fokh0xSbAJRHhYbz0uAQP
+Z97AaZNqmprHo0cIK/RFmjOYJHdaAAfvn1JRiUfbG55CNpHo5cm9aHL9MTj/j4cXjv03LdN56BR
BHGEf/cahhqOQeCP8UB9BOriMCBF5Y0KzJ5Xk0cAmv2fSNYmnI7gcxDMaa9rTTMRzqk3lg40pd6p
j0CIcebkIxHmQ0s4YdnN+CoQZIbxib2/ZXIfRrkj6h7/a8YRXzWja8JgMjs4GXGWFBLLCToFi0hj
FPc2n6fKU8/AaKh/gLmOxW4T5XcWeF4iqlr280gYM6AcDqwQueLdCMCVJGVyFjSfl/iJqK4k9xCR
GRQuWek6FfR234cn3QcGpfnTKathQw0/14taiNNKjBvKDHBE6HyVGMMZtxPqzTHXBrARaweBLXjo
SMhSLa0h0qBn0e204M21BGkMpR1CWk0KhMrGgLAtKg9OkbG+cN5rmm3IK+zerDj85eBhunqgZYNE
OwQCtS3i7KV3nKOiQSpyKYyUjzOQYUTy+BtQHPQsS4H1hcqhhNKgW/d35BeaLMDY9+hHVN1eRonc
uOvQ4WO/cg5FL3dvLiE9VKhdbVmnR9ODXV+opTCA8ajntasE6VyvAD5l+dowaI4wYW6YZ+AoDQxw
Bhn1fL9vjP1Ye8yP+bt628g4HwmbEfx1fZe0RR/jsRB3fukzimg19tuOB32lyTJ1VNo4y4/aE4rU
7eEABmxmuVty4gVVcbZQLaM2GEcsbSLKMswaMJtHB6PpkWYvD2o3ieIotOwT2ZVFoobeKoLQNrlp
w7Hk+979nMOz/N3ovQ34mMfw62MaajmNEPxmK6px/K8Hgg1SGzccAfT6xc8Rq9S0WhV2a3nA1F1E
Y5pyt9fGa7bXPPAdYNgRrQI1b/Vst7MpW1bOIuijX1jw/MTdTUE73uvLjSURHPuu8ES8ja+7ezH8
S1p2AdB1Y7eK3KM4Vk1+aFbjipJxj6w4rHr4Lrxdi5r1B978Y5uWPmJ8skUJ5x1xjI3e6ZfF0kXX
O+UkPAOq2ntaFtzPtr1nLiiQ+FhBF0zu9wF64GHmO52e8Bco0wPJWpEZVdhSMiZf/WE7SJ1sAggd
Yy5Y8AuEFkc8F4OR7aPJpBLvSQzA2Zy/zhVXjtcfJjteBCFxOq37v1z4bdEU1r2N6zKHptC/ciq5
5SlWmbbzYiLYqrv2lQSte52V5Um1VtG/1y3UP8ecg/35tPPxe31vKMX3RngEwO3+FTvzA9R+C6iK
k3dTZzVaBRM9cJfDZrrevpeObO9d/xmfd01bMY8O1LEpFmoQFXqHfxRz95gKVDP/CV+dQUGveysE
dL8Q7Fj9FCy1B61QT0thvuhZ8+B9XdecU1HZvMD4+O1iC00H6Yc6cwie2Z3K0it3Qab8m5oz386s
2OAhK4lI4043qzGKMM5BY1soEBZDRi5sXx1ChmqbBvGdWhHJKIebYpHBBnLW5Cddf6u4zSv8Q9YN
CKjxJ6bjDg0WGtEzRnfEGdmxHuiEUsPh1gzyjU1slPzyqdYdqGT/O9r1CnQ2b7SML12wA29kb5ht
0qX7lsOn1DIw405/KyXvlxKMmYJEyqPdSPNF+4eDN8yE1bTeGNpaBzUTwb7QpmWM395udrjS1VJO
AHVzlfJbYG/LX4gteNNwJi/N0SDoPFZAg0TkSS7UCc9X5bRWmdRfyyQNKp4nDjI0/vajIi88uqAX
ZaRGVQkEWdFs049Q6aYDaV594t83YlcDHQ8e5q+nzhB79jYd4ySImmWYYlRF2sulvtQgGtrau92V
+oQ22EZAvsk9YdcFbblF4oC1SkH0F1Kv7LaQMnUKMZkae0AwbDwVU0nU4LJ/VRSXgDPui1udkQ39
kepsFBJ/797Uil8mYOXR6VuoDX15bzgsjwLBeaaeQd9uX3fRFg/ZaqAC3Erf0cT9hxY5DyG4sHdc
/lhw4SAJU4ui+Y/Kt6i0XlgLtB6VHDgc7xnK1O+LSrL+LH5YN/MQJqslWgC8iR+ng0G/szxg4PYH
lcQBW+NFtj7tWVQjEUe0b73jqpRiA/rHAogt1GdxypMNRzuFCjHLGHB9h6oNsb5qLyd33VaExuUY
a8kbgwv/GOATt3VCPNu6oIEA5KInrExCe4Jz4PwqCjsatLg6yN8AgDRhRseb3MECTvS3B2VQoZGo
NDeww+wjj4mtFxQXBTLKyETcxqlYjFkbRm8yYD+tLy0eyGglR09ecpZNf3vurZBCeiAdLh6/wmuO
tYVKjSh7RHDeex/rYBAbx/DTNfpGnqkQfqBvpCk/9CgKvmplgo1hBKu08q7Y11S5v/OyYibqAc37
LZw7IMGgNKFcPoC5KG73NcEg0tPYLGERG0tdq4nuYMXAn0xYRlvw/7+cOrGQiHKRcfdadyFdIjot
aXyNw7/RqetegJEFdhm1v27g3KqvqbQWaSqIiuTKgXWWMTFIsLtPXCC7C4TRyIgEwMkHyW5rWl3r
zTbOV0K/HlKdbt7s1vO7SbvsLswfA+t70fmSvrf9chLlOlIxdedQdyqB3OapHGwdywzeybd12h8/
+SDHJF6aq49gkbTUPH8hzVkKTSHv6+X5ezKAI0oy+DSqSIlameeINxNn+Gn8eGN0v/UC2x5tAxEt
FtDMO+If9gZokyX0XgJpCN0rGDfwdSHW1mgIyWUpfLnUHETiDSVueV3xYHqM9xpWg1PuVMGoCz7y
51288UteIW02HAcxOdJScwW/feZZOuweSbrPa0IniQq0ha90wpsk/e3aq138SUAjGkyk3Q5QiBKR
TENnXqAPc8mSEqO5mJXBzI0RE9GyjVzxGKi5ue2smdeR6rjHrFxEXg/a5z8lT5+U9HY+WFkvIyjM
jg6ULA9KOA5uN0BIe3d+FdEWt/LVJYlA3PKN1W61ggA3zlk110WzwRvZbUTcpLWXGZkWtbCSrNf/
02Z1L0KVuz/L1ldT5rRw4VrE6+MGCbiTI5qOOYWMbwFK4sYJ1v9eG1HL0mEooITbtP2qRteYxSH2
+zxJk+SKqzy+pBzNWx1bqg6FwGH7V1Cpg5ldJqYQSifc8NjOtXC3s1RZJbqeTI2qurN/dmvCqP9Q
7zQ+k9NPOzTD6tX/vs3XFUZmuPDpN5Juei877Pv5+G16XeRNbXhUsz5cgXrjtukl8kqu40NNNC4V
mWd+W1YWUeg8DitrEclnvibnFSgyl/Bmn184LHoSFMQnFLq7j2dP8tj4z6upz2dyzI4vRqZgYjH+
kQgiA98yiE8ea9YrCGrPOuPZL/kQw0Y/suULbgF/jrOuzci4dGu8cHQL+8ueaO7bcKpAekoaUW9H
WlVYj0+qnql5sETbA3HjabXiXrYbMyLy8dQX+eprKRmSsdX7UH/z5wolu9qVBD/CCO/CktskwH45
TlvaZSVFOP7FFjqghXam8T0OAjaLf7PDhv/bIYXDlWddyUHhmZO0ifjT9ngo+KCmQmfbOj3sy514
+CNUG/AfeuMqw+N/PHlhgkBnGkAF8MBhE8xl1T7kPjX4z1QVdruGHqnfwqbwPRbM6sBI53ePoda1
akwyfppBrGMxtznZAvT0VauF55Vaqlr3AItnfmTuEj/TLzfVQHiBnOCZ/ls8e7Pt8oN5c+lbfoiP
LbKDMqRwgmaHWhSQJUUcvrhD16y2eG6gHWBvGhc/O1px+I9Lx0+wbgk9n2YTpk6n2mFu7IQXaJ8C
v/8nFUWcElokjOAoPyCaYzUrHnjn1USqJNM/2izddX0WwdroWAsDdko049iT9lafAvI9hxsYbSIg
MMEZ1HOV70xQiuk3whvVxrGE1rYu/dLxTZ+ULCCjmRYIXvaADgXzvVphUwR0tHjjZVXuLhEuHSkw
Loo7yOkD4OBrGa6qQwcpgBRItfXdkvrxVBbaTPnXyDychlere0xe4pBG+bZJ7zHgS5k+GhJK/3MO
Cd1Wm4ZhSX1zjubVEwNxFMQ58hH+X9e5v9DvNVwX6d4XXK4rjDw4l3hC+A+63dwo81x94+52cXMf
6p4JPYhAuoHeOwchq8JJ2TUH3k9X9+oE+vdot47fHci22B4m8+DrAN7bWUvBXKhZrJBnDe7mA0xf
smCU74kMUiZ/y26lD+WbxfvIlmPKbYF5Zm5Z0jYlXpjweTxamJuX2zQXje3SZoKPlQvqP4i0Jeqh
tTxWsevek4Le2kCZEo2A2z7bxLesx3zpAnBksy4YBsbF+U8j2YsXMV5Wo6R32J0w2XCw/8hz5vrW
sP4CNV9LnQhQXHNC4b4PXV/OIF0mq6IfqFtdslzIShoBX2N79N90Q1dOjlBE8+RBOGI18tMDFbtN
/QJA9wqNGd4g0DHsyd5vb37E4bOBF7GIAcR2j0VDglblQD6kch0ss8CtPGmVuvujsWtVTQ38SZpe
deUp/PkE7hFVmoNUfn85LlzgeTVP1MMM2moYP5Tbb/JyMi4AT70I0WBFB37v97yr/gwgc6+fGTNm
bsFFKcHvUbTpMd0hV8isjO9a+GvuC1yTLpmgwlM3zKRd78ikVx4dgp2Br2e4U7/fFGh3YrbAAZ8z
hz8sv1l7Yt+iLdhZ8zQ49YZyZokAo1h8aBDSDdQ7mGbjx3XiZJDXQCdKzjE0hpuBd5Pv+gGxvpGT
IM+o1LwYt25qiA5mXua8hGf2xZZgQYeYebc87Gz4gFEU7dTkbBAfrHO+hVoRDBfWrNogG/9cPQUA
8PNulaNxeGFAzp9bbK6NBjQXhdSo8SuYcGSQm2aT53YKSAOmy3FdVx6SGAJR5IIW7rfEKzwHZwm8
5tAVmtWfMUVefo9rCktQFkzSbc47AvqsNrtcecdzEfJRDD6rxDTW3OD2TQBMTT/uhLSty36AwPmH
v8n8I+KPGl1t1B7n947AU2UdoDwpa0eiMr4mS1S2/eMi+8Hd1CEiAEZw3Lqn7dFvytfmGQJQVjQi
5D6Rctwxs9U8jWpjS+IdUcDKRsJw1jRdVunHnTtwi92Yzh4gxnfwFW+IRqn7b7LqHzKLHxjfIJwQ
8BdEJxDEQRODhyJpLPFSaWvmUTE/WSkqpyRFaglHdLZqMHqfdWahLIeKgA/ToHo5Z3Ooz4ggBA1A
MTAPdDCkVknzEiSrMEpto/NQkv1tkQe0tRDeq0ZUoMH6j1c2gpafeBnWWDZMNs1ZPIVApFGTvZiJ
OsiAyLwLUHG4VSoJeu1iDPN9kiSogK1OfOR3jhS7HiHr5WvwGRx/0sb//ha/TMgAMzrMQQ3zOu+a
UB5URJG8EiKQGOBc0H6uQ0DtO4xzdedxNTJg4RxYcRYuD7iLgBf9wMlWdM+JJttpOneyW+eMo0se
mCA+Ve0jgoQ3XOuZ8yLkzPZK4DX7A4tFgd0PuBSIbCwBJtu+7FgK8hTxYfYTd8Sd5nahwCYKkZgr
qRezYM3snnzaDbiDdlLOxw7s8/eAgWfkex04VE6SqyM9l36L076QiRJS+CkF9QuBENgBfyygjHq1
q3MymDc5G3Q9NAgmOyXAb+xrnYODWI6f4jkk8yHpOJF4E7PNomyGhaqNAxc5Fi+nDdpONbFgIwQG
VpM7G1ao/YTIyOCHC6D7iynpG1aboC/ov66kqiD7MI24JaaF8R8h8Wm5PkdNCCiOUl57h8psVUCq
vgCoc/IGJa/JHhnbc8PpTFkIjXFiQulLIR2tBHhJmouOWmr9aPXN17DuWxZgnyAwpfu68M+JvhXp
mndBgsj56OKXjCCn2TnunOwYmydf7Dw9IIcByDsiN91s1Dgy2+/MALsIGKwkUEUtB0WIRiObMFFr
ftQeLlBLzANH2srQoK7aB7qgEUQiIaRF+hb2wZM7+u+FF7NjTNJ0Sd/BE1SxUIWGGeY5MNawqJ8l
5zQWOM56X0UQMDd6/3fGelBM1JHTqUODZ+fRNgtoUZBHTJ76fp1Qm4aN3vt9QRRWKqIxXOx+K2i0
bptx4DRCwr7jKQYarztnRTEQss4q677YTzZlTcnBcCFRQM5ek2mBKD0VoMxZ7XuhxwzAANV+LjbP
Bi7aAOGQxg84uMg0SsWtY2BKpvP1FY8r/g4E66gEhTjvZzTfVCbshYLpS3v95vrcSSRaPI2eShON
G4uLDE6qScz9lA10KNURtJ36iwcr1joMsU+HQeOlmebOtzXojyJLK3VQ2fKbH5jKu2s9duqn+veE
Aqjc0TXn2PNBBlrbIdt4gpZ9M8u88qpuGNtYYjhVkqsoOQhEeASQQaLwNAlSY3vclO+BtoHWcOjF
ml0Z/RguWpIIg8j/xpPh/+br1wmHYmettGwm0mgpD8t+FAHvDnExK458lgRfJ69pQBkUjig0VJA6
pfARPoVOgFMHkcHeJVIxPG7f5j8Wiv8ldVbhUQ33SuI+lrN65yx68M7YmGsxxSMo3S6HMk0deM7D
Y/SGM8np4if5dmTtmlrwf7Q7zMa9wbpM5cLAOK/XnK5/R+oUGSwEpExZ8k9lEgIxqiKU6yTFJyeK
zCcYCt3v0HaHQAqSvBiZFud0C1weZ690H/kA09V/vKL3n5bcy5bikgUZVnxx0ELUaco3p2sTIKlH
HMnZxG6m4mVS80N3IEdXC3FA5HNl+K70pf6m7WPyTB98xvimorz6Z6mpuDxmnKGwER3Abx5gsBMJ
FeRM5PboIvjLxCtuSnJbApyqwcTw7LVZzlyh+6VCX4fFh4VXnsw0Be3E+shL2FmoTuzgfv8R2OHD
TNDH2okdG2zQo37GANLNqz5NuqgKr8B3VtL48GefLU+j3rv2cu5GEmMYjZIUUsPDHRqXDDQJxST3
5zV/lUPUksYEgk0aI/qyMu7o0D6aQrkusZO5SqOkV5CgIKpCOaw8hnWGo7HHkGqBgEG2NazY5kaO
/AbJDDZ8P83ZTVfhWKvz4SbOqJkeG99EE0hzmDrgJPsHidMRoSHCYyRX8ApvHIXURkXToj8xP2Uu
0rrvrJ1O64VmAAYzp1+SlyvhBBmCgAY6A68wNUVbq2V7fo4PpEhrozVKkawzJxNAX/RjQgbvhR1K
QL4Tne/qudm172umHKNjHVBfpJbWjg+SB1s/2cichnOfA9+SfsurcytM9GBghq7pEWEPPWqBxv6X
3YC9Aj71Q6+hQPW3vqYpSUyZ6e5hWbOHm94XjUKe//GjfwrzPOEjFaevzb9NrONrkcihf7HRcczd
6burf8Kl/IBI0mbRvQcgNcxidje96Kts3uN16i9eE5H/zKeFNR6/sFJC6qK9NCEpm/PcDoiiR0wC
Ros2Udw04hlt66rzWvHCiCUzET/YehCJLYLgBFhB51+J5qNKhe5fMLl7iKRE75s+yVRxVMZlbDbw
Zd0uy+9FXXhjxlijSHgt/hGaZ36zcQsck4zij5yDe0OhXJy67RkAU7pDdPjVYPSBhRHsO2gGqXFD
/oZP0+jy0J8nVSryFdq79H7/kr7TJ+5Bdz3o5T3rKYuW0mDNo8WLLwX5IRzYxRTXv9rO9leeMx9i
fOVv5Z6CQAqdLdcL+gsiMz2M/at+1uDIgGxnD+xVcjbI+7a7d9vtLGae0/9W5YZoukt9WScBb3YZ
jf7ab95jfm2nT6QGghAgBXfUrYPljrZR6ert8BTaZ44qDnkarLZJFIMf/WmtuzcPd1fVJdNK5cin
dahxcoSL6qeEDWYZkIuqShK8ZW8PuSPaV4WDRV26jMfdp/TTFA09T6SR2lSsCVftqUfk9R/u0/hQ
xbjv2wdh6Oh9Aq2wvUAnmpoUMgYjNHUcJPCrKQAV+2IQBKEpamSL4MdFUCGyMyOM8hhKe1yvWhOW
doe7hF5XO2vjAksWvqu79lKZwXD7BFT53pEFCXZQo9cAAMcrgmDdTF1QsVzkJYfKk15YjjLUnFrg
NXAqCyNN3gBbbKNU46Gn5bTMJOVW7wP189xv4x5UK6zf9Ri7aGBISu+G7YMPrqecZrtka1xV/uFo
Bu9+wrcQQ0v5dVk//ZSDeXSOKpe2HIeLnQlft795SQXLNusrVuNZotd0bryZ6fcodsjj+nJbaJje
rwl90eTRhQ1mbgxz3mBQZWrAN/7DfAHMMomglY4ymsDWIUrorobmujsk3ye7INRvT3XgqHfu5JEd
338J7/97yh7cI64J8rULUIzeZEuC+YDvPqkar60NSrYZn4mJjvVeJ7natwnSt4KIZScGMcRpNY0f
L8EiOO9myN5qoHql04vI9z81atFE7wNZZJgT41lhZYsE9as3NIgtWnZqR1YHJ9AWdgzvwbKT11Mj
u4SQ37/ZOz9ckB4SC1pMdgFBRkZH+2eU7xooGUUcMy4IzQ2oINRKS9gNIXHKF9wVBTfBNZpUJc4w
9qQ2/4BkO8yCAX8A3NXBWN21eVFPygsnAZ+cGx1H5mrwk7QC65S78f2RXgj+QokVJIctHBTD0/Ar
UBW4KQEoLFd+LRR51NesDD0JSfJEiaR1R9s27ovUo3/Nm2z5R0ASBuuT078Com19SKTLGTBcb73h
w8bPZGMaKvoUUxHQcqMhkT+cptrOwB2Wjx+d4GJMWw/u0j3KNPbC9lMzz99Npbjh63q51YI7w1CX
rjI34qiWJJBdmLc7i5+3oGwlU5ZuEDP186c6lywA/qJzfn2M5eL2OcDFZFtkN5BrszvaBN80fNuv
x2CT7LoWbWlBbfsvL29ojJhw0T/clF0AxUl1KlORC+wVF8OFqFv90dqCVKWoL75Q4w+g3Vi0Un30
xHK5STKfqLNNb6oAo61DIN7X/QbEmTlQbGkPQMBu0JZcRH73/FoBSswWf5khRRwuyb+NCxtnDzgq
hC/uR+bqTQ6MJmo+P4fspNn9uF33ijEOAAAFKWsInb7nfDzhI9NJ22tlUHZT92FDgn2B/dJqSzOA
6YeIC7HHQBOSIgs4tQ6ncbCe5/tulquBmF421gGvH+m2g4GWUX1U54E1d1iV+dtCX1A7aD19mYeG
A1eMci9DNVjZdnznqRmVm9eM2hBmWsxzRYu5U47ngUpaT87lhvASTyi4a0MUqxnaGQu6NdGdHK6a
LKi8UIv2+RtskXzBqu1YnHRE7Gpx0vMhLIMnbkMg4PLNsGPdTKwzoZknsSxaR9J9Dlt+FnLCihbl
4y3QUgyfy9mefdscMqkI+6j9yMlKmWjNWWloCnmhSBmWW5yHD62as9GPjKi17krJlxv/u16dcjMt
TzZ/3wDLkNbZWdL04Dm1OnUYZT3TzWOk8FEzHiuXz/aiavm7vpPARPozELy+FBm7K51S5Y3mHxsb
X/ij0jAbEhQ+jV9ScGCZFRY9OU+ehAsoTes4G7vNDTRXR5vp0DaOkauYpn8QwrkD1XhsToJZFp+0
rtBl3AkZCVuJCvM5KRj+zJRVigMd/R1IKJtO5ix4Die8VGbNfYuwFuN3xTWJ6cwRTa0qZ10KtBUq
GAHmpU+VLblBaFQfiHN7Le+o+yOWSGqILqdf+t7EaY0rXKFz4AsihXiMBuOWc37uxojN1n9E+7YM
0318XaBROPnsTl6NrJoXy37f+eRyn1LiG0VJG0+7WaNJINYzlTrNYjbXONl80a22l4ATgwcTy5Ih
2dJHBjwnx7Nhe8yFmXp7s5pApnmA7+hmS548jXX0R1Gian4WQXMK/AHsvYyz2uslVHJcbaLCjvx7
Ciq4dGd4WdixVgJjqZBmOnmVqWphUv1UmiTuzCVYdxLlBNOO+Xpwq1jyd2sMtbIZsCYmwUfkQ6p/
Rn/BMCAFEMAHgWGXnSJLwd7Y+zwQ31hBXBeK0q6dN8D2rmVvuKYzxLcN50XmLuaRYy1XaSjINQ/q
wlUVOiMsCDNWK77ZmANbH57skHdU0XC3nXKHMOgp0UDo5uvA437TpLdr9CqDNftLFyveGBd0Y6C1
s5/mbpEh6EnGJrVDuPdNQmgAMqIOSpTiCRG0MvQKIfrcDMepvN5EtZBXO0t7f2oTLXShVLcTDdN9
KC4wS6m9oDfnTl3T+2aHZZD6WfLzP1CTc9GJJwJQwqBcFj2Jf92/z+5pP5EalYriwYLNdOQCR800
V/Qc+vD5iAqCYP15OnLb44m0xB6owmSS7ulpYyBDfgKTpYbA2SFBcHI8QP2bwnZMSe4l0HmLlGHM
VPwwtm9mzrgMT8voBoSBMSbjcWBlR6teJDEmRKsAGehrYEnUPz/PK0AYoFnh+tf4ImJi0yw7kIV+
qLzVxVrouvpQdkyUyiDVUDOKMDjFktnlEcq6rZ8tBxpIZcOD8CH/1JqqLshdKr83Wclp7FNeB7AM
GY6nHXzrkSue8LAnDoWvXwSYKT6imjXt0OPLNOcUj+5nyehTwMewKf5rfCzXtMrxBytaihyq5DFB
DnCTD1A2I5QB2PFExPg+9E7G2Z3LIXkuAVkGn9Txv8ZAVnUEOiPL+YMyhW/hZNG9fzcjYBmzbHud
v0hoWzt/AlPSpi5C+tpF7OsIWlitoPRT78NSfsYzn/D0eimkMY3IU4uJLOmO4VgCX75a8F0sZgZX
jzBvUa39zUE0uuZ+5n34asmkNZwWlHsplSbUMwKS/Zt9LqciE5SIZO4YAYwR308WAzSN5eWtlb1t
47+ymny89H1vNyj0sLeIqPDwO+7qU0d9fHcgCo8M7XSn0t+noryaDhYVCt5LCaIp94dfIxk7zaUA
q91ONWCiYMVIRtdMfKneCneuSbZSEva2zwVFqZYMRoS57alid59Miu9eINueSrgekHeHN9WceFjn
g5Ponf4iV66AtX3zBOmNd3ooWE5xoWVtC6Uywl3T7ohhItj9LLZdDEdpT/CZ/itZDxi39aeB/ROD
YpXOuLzzJjI6hmNz563Wxhwp8dzac3oqneV0fbEi8kPzw90RZmfuoCvaHN+PHTiCptTEmwuVx27V
HsiA+RnDe0AHNdKHzK4o8edWiAWa1UHLF2sJU2ovzAaaRaN4aLE7iFtBE0opxu/quoWLzotujDVa
QxzGId9nWhJiGYUInah/R9vH7aUtsEfLqz5Llhd3syOLPXY4PdHbwat0HEl9DpOpMAWHe3/E9oth
7LNPnaDK48g558oi1wmqRymxiD8lzv2veMXmlL33zqyPgOYgLrL1kD08WD79FFvFDc8IL4cPpi74
KApK2mWlzoZ098RR5MXIyU2EGii6FgIkjZc7XNvMW7se89wwE5+07HTCO9lB2wX1y5R6POuGfT8i
hTGTy+Td9tdMLnvtzx7MX9nC2NiYyP6sORg7DTeIkl39hWOKwy0pNr7HvTYa4kQewp/GMGg5dySz
34plGcCaJsYXB6WTZOg8US9CS94WwXmBFHclcqAPpcNO33iVrY00DPKmludkxU65IUQRJ4sETOG4
Q72YpOEr3obewLYXN/uagv/4yvXGXrS8IT8+6O43sf1SNPyDw62UG08g8RuNiQlQEF59348uku+1
VXaB6bZI2DYGboOmGRE7ajhu2jzrYxtYKI8T6s8FTYlA/X6Xa58OFs38uYqPfWpCKTZOYGv5+ZXz
Xpr7ucPIOu/7d23yGr2GrMSbqYlGpkz4YpiwdmCtx7WkddnG+a8EFWhBJjmfq6zD0zfnwFURrFB5
nCgZGJ6F4CRKxmVDw2Alt1dLR1oT+sF4BnmM9CX7zENCGfRVeY5jqx2f1i/DIdPlivXLY7DRkS5A
Q69wnJajG4JZeLaF5WCZ9K75XIY37An6MISqmYYiletzZwPI+H6XauPYtZKB8bEI4BNeZJ8T8rYY
zic/dl2Yt5Tg7m6O3zkEpMD6DHc3Fn+EkajXkUG5OEZgwH05Yvi9uU/3Ax124v9/d+sGtkY2c6Wg
eWF6q6lSEyYOmy4nIznX6fY+JA7fA3YLyRNAsEHcFzbVDNfOMrDKnHCMBEGLVG3h4sA7fJ8voMF7
nN/nFhi/aKNf91kzX88GIpRRzfe1LG9SlJSokRmckz7/tpp6xMO6DbHbu7VDE17b+3G+y9tsu6SC
gs//GcBHFyCrjWcEj869Z9YzTuz2wwz8mV/SIRTLLj+WtBlpGS9UBvCIKLuJsL0dAQv+KG4gqPNx
AYGWBwaOR9z4reCQkeKhPG59L41/FIksuE/tWCYJp5P+Pqy0VizOlQ+WvfPjUnmF0QFq2o/CjbyW
DU9SF0HphaxHn/uGWAnvFY4aLUShgzaYr7Xb08YRTfOPmuHv4E6SiCueiK0YOHC3D9FU5e5RlTib
+8rlSeVhzJTaFyim+alfp+YlRaFqxGS0lgNqjaLi+qL312VisV09Huf4gXN0XmzGHnUAd7P9xYGC
pTTDLz+rFE70hA8V/NTOY4aFotLNLHUVYCA6gk02C+cknGdJVaiOfCXzWAC66dz56EKj2JUMMkSi
XYIiQGwxeXxRvEAuLXqkY1sZgBzMxvIK2Ox3bR3IWoD/7Wz8idrBH7dI3Q0luJKhlBlO+WaurpdV
WK2wIuvY0XPufwMvC/NSkf8T9eC5n+2xe8xlcZBsrFUR80qr7XthiHRB6Gd5B1R6ALtJ1j8Uogk2
Mecz2Pebc7qXyYAmyGNwstdHPD033ItP5J/U3GJQNGN5xYub6dMHc5vqbDS9ZbRC2UXAZl7EabPJ
6w9hM5FG0y0jDF4LYNmS57lpm5ErZ5442/Y4XLv37vjDSVkRNC2uUUW+4vMXAIHA0Ou0xLVTOu9Z
Fd4nE0FS1r+Hefm87jbvoGKooJMv3pZ+MZo17+bzhHAb6oydmr6J/kJjtLstFChEpuytPE338vA+
zJLCe6pKyjyfAF0UUHqSQKSbO8IQSI9ufPV2aESJ56nBRjXRRuuSbKJBeVswMvA4ckZleC/zhP3u
+uJIiPMWV+EU2+UWavzu0NOvi+3WnDvwy5qdpn5yBpzh2LY1mZ4ODNXkLhGLYv3YlUJpx5tpDM2M
gs/aZ3KWVQNjkoyWHgbl/zvXoddv2A41fRsbSw+Sqn4ui2qSsr2LUayzmteT6TNMrjDjpygruxMz
Bmv0AnkqhK7WA+LCUFkoIhOFmemKJaHLZ2bw97Rs9KNX+acAYXL6r8JCh7Xze393yY6Zvp6dI2D1
H46/43242aNpTQZ3p2e+XnpHRGYcxe3NXM98vpbqWpWFvMCW0oC9h8i96mYFYi7K9qI72hdD1Gkw
/U4u9iIfGvvSQ/4a7mmJQF/wHqOhK03ic/VzmfRSOjyeN4xSBEgJxaHU9Bxhgp6jqrrLVME4My7E
4TC1MfWrnGxVoEy3ZFN75PfORE3gs/K8RTFkhRfEzppVHNrGDh4+tpb36Im6zys+HPN1A9gg4AyV
BzmimiNQGjxmgpVuCxTHKKPxHZCRiOGeySs6dkQ8hQKtwEmXG5u62orJ6gluRjrOkZ4VQGwWcbEb
Sywros03qb9CZoGcfXb64ryLY0AdQdJwwSHitIxRJ8p/s8YphMJm2CgX3CEFo2t7jpRw2mZfyIXa
p3BkWNKYeL0Kc3fz5ScqEydZQtFcU/HwV+NUqwmQA0b3TFHHchYIw0YjLTJiOOX0ORLLnl4IPbfD
WFURz4yqqTAAQVU4Efz7T0eFddqhV8Q06TlLC0yHLaCNjDo1Dqlj7E8rOz4wKoBD/1YPykGwwLbr
5I91ot83ixsv4VbvQysPI6ZCILLqTnbiuGCCrORi1ABoKr1d+fQcewISQx4ojAVtp9RwwvpYW5f0
WeAr6rB9sowaHQFrxkJX1XMCQJeuyjlZ/AT1Ge1Tvm/K+BO+GKhRDVWtxQvGYJGDCBpoKl0goNKJ
JKF2eGeMF/j5lPV7yCRJ5w6ABgZuoRz+bIXiCh8+mbA6F2u5npnPKIQ1ubtz1mBj2Sb7WcTa4Y0L
TosFyzfYlyIIPs4AozReT8RApxlZTZAq9TaxeY/lGaJYnVUPwwA2yo/jfwvPayPnfw2xsAgDJYkS
ayDnut2pngmQnJSUXxeFxCOm6+eMOsiDUldp4Pc7WIlDsZ6Lc5jK6BvQlqxP+pA69F7Le2+65kbA
coit7X7PVlCODE5TsjnwMKh4/cpdLoO6F3nf+8o9Q/F4nW6uaKA1SA+QjZSLHqD169oHMCYpCqUa
8re+tDcVQ8KJEDcpQke4cdD7AIcA2RwV4WJD6ET6GuVP5WwDwfKSxVbz0oWYHtEKAc64fKeeuORR
Zl4kDM0hjd4MG737SOryfFYvcqCco1FdJoOWiOe8pQvHtkXjf7YlQwCQgwYSTR0kujV0n9Hau61P
I6RMx/K4N+uDvdjVmuCqjy5+gUh7u75p/K9WEemoxk6O7AXMssaPrxjhh0JjFVyVEj2VwGk2AVnW
K++nT4W7NUXiYmXyhncNBA6A2YRUwCvAF5KZdoKkXhh847cf+f9WGq6V3j1WOeJHsoSrGKmv1xjq
NYnegf9SSsWSK05I07hUN8P5ifrpbiZORbOlts5NP5QCVtlYk2gDGNsLAc+J/kqmO6KGNHIZ+qXH
1us8e3FmKDNjtUq/ThZQU/zeTFO/xqC1T2eN/mze1YMY4aZv7gkxRpncAZ3a0jN4ZK7h9orfm/Gl
EqvVRsEE7fHgPNdPo29eaC+MbI86LBLcZs2eYNpdTnd11FOzVJG/6ZdQXFrT4fvecOB2vCfgbhma
p7EANzUMXSPjjStVN0BIkBG3sjU9kMafOC7Dp/E3gXDi5VREgHTgCPclX9SsmE6iYTSkFKnvxwmC
b98UyxKaBQIaxC14OLdx9aYpj+V+6JFiX+4PSL25c071Nqr00dSnxHm60N30B/GQdskSX3kYPRG3
s7haUwpSfjCj3w70JrYdJb1iBRyO25Hfs9nOxPY+LzaZNGwX5brOlu6A7mGn8wb+08CFCFKAK0aF
fuNo9xYKDHEpYiuOzAiGlBMNUSKJnttkXT9TmVncQ9PfhGgoO/CX1agcmxJrJyO0weSjUPe8YtsC
xMdlGewMeh6hkOT9JPtbaaHypdPvvXk/213GnwJZiWSOBX+mWaqHlHSUoAcNgIUiMP5Ic4pd62DX
ZF+fnscrPWIEAwaJ5VzlSk7DCaQ6p1zhJR32VgG5WcJPOG4sRMIk8jD2zUZ16ViyAztSxkVm2eYA
7FJ7jtlRGun1VUH5HgLzZ7wzBvOczYtpeR2tEWWm8i+6XMtcxVZo/KU3fT0XcDhLNUF1Q9J67tE0
d9WS6Au8jpoW1XWeJBozddZq0w0RwbDmcMXmTXWYJaRr+6TNBxAosR7cq/j7WvWBgmQZPWnrNgWK
dNOIyQB4lZmMQ1YaFtcCtfQ4ZFCL0kPfg3RropRmfqsHcOg1Z0Sgwv/gSDUc1GAQs0zwm0AE6TWU
MnP2uA1Gh7J5KCh2vlgpsTQiqm0zsVX9uTIy4bN8I/FUc3Fkn7wqXPDONYKBgxE78Pph4JGlFG4G
g+Wpz+QiJaMYQC/phGI6LPnzR6A7qfwBXYhJUG/1QhEbV6pcQp5+4rrC+Jjz/LKBmKScARLe+CUO
m0tl6xgellE3PmiGmI7FjdSvVBIZ7GHl4R0yOb19AU7CDMK9AfOb5w/14zHShQl8UGZF72jBfabz
dv3EXbnS0/E6P9Xcol7OMAOWiU1zqzGIOv1XOWltA+dWJNldN90z2v6y4ydwrHpCNLgbpecYlk4o
qghSYiU67uGTvOiDjknD6HujiSvtqEwukP/JVvYYyjNidgvGgzi1rAQpJholGXoZwHYk4Mh+Ixw2
YzlFaRb1ipVBwlzVBybiJpxo2uApRn5JcBOiGBWIWEHFlDPfeJza7dhjy0MjOdGQOGG0NjRAeCqV
UCIbDlylEqQgGgRcBpuQkHTfDqlTJ/wHJctmZt7bOdpmfDgsvFnrtHzpSZZKHib6Ma8yq7QMIlGX
UHSERvIlQD3ABxqpnxQ/2ZQgZ2nUcvn9FfqZGRhBp1X4ETL26sEaMaM6ehyW3Q212R3LDyK8URqa
8n3I7PYxwTICLPEDtPdH/geEc9wKii/jRnVI5VbNT8SAecWNQoQSH+ThSIJZLz0+sIBLr/QH5pwP
vQXMYDU65S6osj+xtQSXofT7680ISzadxYzouuMhcJpqWI7oWuDSrVZOiC2G0AoaodUh2rS2P3RP
fA7hOz3iCeo0vXFlgiMGDnWohgiskcCh5lHKEvhO5rlfPehQVp4vTy94VyRTh8yCEENRQBKPySK3
D0iHTZ8tZtVhAcPBAjy5SM/OsOVOk7F+ogE6jboDj8Hg61T1xNUt5Fy2w3fQie80oN6M/CC/xnHK
LLXy+NqpJVEq6vC/rXDGfuBwTzYSs+mwtNDMkrph/jjk6a9MfukfGobgGrya4d9tPAzH+r5Y4Qzc
XmJqBrbmdj0upi8qevIkvP1I2bo21oEnhwyBT7LoyGIqZmc1GL4QTIW/0wIMO7SYaOIpRWVB4uz8
fJYOobVP27hxhv/ihzG4/5Zw+os/HNTAF3aFSchd1fd2ZpzE2oM+6goekKjPoKINu4Gyc8LmzyJP
5jsm58zt2lQFSELTDSV7i3e7860yG79R7eoAQ3C15CiFoN0pj/3o8rCqkac7pGeoXSQDeFIN7Eml
JtTH3BlDOm3nUUpr45rW9nvr0/B56obNft3vbhQNWNpT1w7wzphbC2dOWd7Hgwn+z7t1vKxShRXC
d9k3wHkgpP4FzTT1YYq7KvkcywFy67MCvMYZ8gPPY5AjyXlyueCmlUlTjhBPGA9cMIZsbgTO7cEN
ei+1JLz4yyOiC2+oer3giFJsn39H8iKNWKuvI+/qHEGqpeGQnqR1B1+AfnoYKJqyxQyCe6GsmYTW
Sbah6048s/SbDAqSBN/sU7kvVb4bTaiuWceK5H5Oct8zlUT6xcY6UdMhkF6tWOJdRLUvd4tbB4Bx
xZDeRLzYn4tUlRkYciZgAPYisTU8Ig2TFppwkaviQQTH/nX3O/O2dPIXidbnoTx7zrkf2guEeTGd
kpC8fUAnQe8FxPMQ68AFuYfQTq67fAX3EtuHGHMs4mFe4VYe7Re9S6SCJQDuzePyiod4ALltsgwO
OMIvJEmT8hH65qwKXWgQHWIhZDbKMyG8ycj/eYBRqGcpiWMp2cEGgagYrHmFIMAUQ+xC1L3pzuBx
MrMhSeXNmCJ+Ne5KcUVDZpAvBfdqJMS2R8CbndY/0LeHGCHkEL/nOOUDKCnWEYhhTBoMlbQydtA6
CItquDsKSo4vm+nWnZnPDzDtywCl+c9DH53DoH29kU7v/MKvKF8ZFEcTuJuDkU9tK+yYJkp2X5kc
/xg9UwfVrlbBTpQiP4G2vyLyl3AAbDKieVzgzu3c0gKpuq+rvlG4a/V7KYJTaFeKq4I8w4B/u1zR
Dc7ueTIKB0zcXXBDqkkis9hQiJblIe+/f+9em87rlKn74e6L6sjCSUgiaeq/7qlQ5QWSNxptGEKn
X0g5WE+PN4SSaaBZhGZxNNaS2ChNNRabJBrl8nm/5Y2IEl4fxj0cr6wapLHqHEsM+FVeFmyn8q2r
v6GvU/UFcOKUrs67Imm35T/qEGX9Y5Ke1cSZNy9/xA7CshScpFjblp/P8srr3VOcG0Eq4ef4lzb/
wf76hx+jow+2idfvXuPt5F0j1fgHSzlIbXY7uRjFno1KhttziZLUBpWbM1reFDwX8yuxvtekqT6k
rdY1E4BZj46Gp+WcxKzOP1G1p4p25JGp1NugS0xNV5yR5FAHXnLtZOLwleyNfx72ALkEvBRjTpb6
YZhsjRwB8QcrXlPyrsGKbHG0m77Pxf4SaCAUuhtLhiRqpyMy5y/jnwHGrGs3tPKaL+8JDJpX8zaj
nrlmC1/4sIAQD22yOlIjObY5FhzmiQeotoLtXT143NbE7Ncuej6vu9uwhus5sr5mF1NvJG05QSFf
WuDrtr5Ce59UnRANFxrpz+Z4/QaNXrAupci6QAl35qQC4lnT5DmYFlDmKZFLFOGA5jSVagJLgJ2c
wLl9gIDpaEqCt6FGKGef/gjbSRcbRQsIKElRt6V+rLep6vCURVn2MY0rAuU+aq58t1xbdyPpdKqr
NzMjgc15CNRQRR5x9HDuIl1Z22W8uNOOxGC+aBMArlQN0hb/gBUXv8oE1xgwWbDYaYNptYjdKXsE
sfi09skWIOUMQn9Syu/Kk05KXihooPYB6jIugqQ9s80MgQ1XCqu466TvX0cpSm09uRjZ/RQ7Urr+
WPIp+EI8FozBuimT+zORKFzzjBqioRoAJko3qnQGWDQnzGwPArlU79o2g1eg6sLQCjo+SdvZZnTc
VF3WnPgpqaHgTRubnucwXVC/dkI3HY9HAPmrW9wQlJEcP65JMt2DTSqb4m3+VRA8vgn+9wz6EyRO
W/uZ/XdblBHzu4HdESLwuF6vJR+jxPRNJP9crNEnI3BOKyxCQw4vqDcFfFVQxlnSvTigLBPTn9eZ
EGFXWjoae0LJer/a4HIbL1uYAMuiUcZmQdD73GLSa8m+c5JE1mv48AYCncB+wMpLjT/kELJbe8Ct
iJ3YdrKHh317y+X2jLw1eJXDwf9NlA6Nw1nyc+jBhDSl7byyIiSxoLXBHX1p+p0vxqpaWtHEYyDL
Oz/lIEW5jx2GLOwIEm5Q4YFIEjhCbkijg3GE41WUfSCbZ/DlCan6mFM/SzKbF3Oeh3GhOWTMup2y
dy8zUUlwNMWsAPW8CWxwcBKHXW7uPp8I99JKtnTsBdgjbcx3+rJowXeS1X2SKNZe4sBV5saqtirT
T//t7P2eC4ToE7MX3D187edbufHBREfo4LcI5VEmkvMxxcxFtTxmlui0FbqLsrXIaDeTT/vezIJX
3ZI/s30jh9Lv5BVIbSFLoTJr+NCIbEh4bpcEmt2Uw+lLDkhxBac86FTa25u6N1lyAmqhhFVYe3x4
pZqHONa3dtzypaObBGAz+7eUQfX3ZjLVFVyCkn27OtcXv5ZyGX7KZujJa3icNqRSX8ERyN5aY+PU
YsbkaRDi7j9kGi2G6Spo8k06NiHdspsGWYHW+PqfjIltpnjikXEg43dzgDMrfrAkn+Mqp5HQb8v2
S+xzrQDYbb3VGhUdhvXZGsQTZbWS5scTNMQpM2nYMegBLknSictvlx/B8h53TmaCQZsL/uxfVl39
FPqpa7CkzT19qoBO2bUWYJ0XR+4ZPHTz23Z9tFy/fcBkwTmtFNwX3u/YBTkfDrSyhpjPEoZ0mjfJ
9AAWEDe10ZpLDcx2/J9u0AoFANRm649CbcZHtTMAZHPIAI5RkKF4pWsy3gpir3C68koPgfqK13MP
Jx/uvoJS72rykKR3UxOu1EN3L02HZ5xDS0JCcMYMbYgmY/3H14DMm3Ss8f6VujoJ8YUCAgNCh9vM
AX+h4dr+Rw+9txtt/ia5CwlSzN3DlwiIeCF5FbQE1fH1C+tKbJFi1gSa5IR20bBF/4MHBdGUxWSn
SIfWnTJQ6Yc41rtQfs4z2t2NzYTe805yZRChiIfZg+MmHkV+JmL90KYQmTaHrA7Yo2BrHxcEjWMn
ZKc8/OWQXs8PlZNmZHP++7LqZv6DD4Tqma6r6yh1EDPSwJRHAtZsCsQVa2G9ZfsknLM0Rzdt0WhQ
w1dRMN3uX55q6BBxlPo4VJr5EhGhn6argEWCK7997sLyIURfEyRVgyxN5Jsy/9cCGOj/cZKnSwr6
jbV+FFbxlUzT3OdvQYlKThZwGQ4i6KVl06C+hdWxEiWMUZoAWHbk3AIIqSLnjU81s7D0B7epWJMn
yBoANxpR3msOdt6XdT6QC2JS1r2ygG7pTPy+cHUoDTkF3KtPaLgZYPbV+/VV2HgE+lZKxNWFq1Tf
n7zCNORg7pnMdGBHCEFiCrngv5xHi7DZMPZzVUBZ0hZhf2IdNc99dntJPu5g1Cw3qZdfmSPKfzlZ
CTjueO36hL3AGXjz86BgS+cqNFniVVvr63dj4x3WrG42deN3PTPFYs6WoNepbHFx6Gc5umKD2EAY
Mp41wQT421Y9lYyDLzYv2dRkki+2SW7YhhJ2vEjLmXjzSYRVxRv61PON1Us/G/G1dXlz5GFv/WuY
9D2h5MHzrE+Et7Kes1cmaYwLwfmK9ObNKWs0S9YdnAGl/5kaJEwZsFO7WSb5xc2+0xgUuGjhQema
bCleuXmh9J2cWRHamzCaDl0LgyKvX4rEnw/er8DzJnJ/Np0qd2Zr74rYC85sLFegxVqvR0J16Hgt
Py5hILTo3c2mpCQk5uAhg6ja1ysUOIyfsDH2/IPzjqPsTzApHaZwj+hVKKvdGZF6IOtRhIS20xQL
Ir/75DlhGOylDkmhg9LC22O55sRmuCEt8FMTLWddDwoROQxXLoWhShJLLw4+6lEsNbWEFTvnsJHz
S0J1NlKTk3IpEir9SV8r5rvRadYSa7MPZvB03dyBAweNyirKGoCcQEBKWg49nAyMPKfOIPqFKNbj
Wjw8mZHgo5hVopedL0sHhc6enN8lp1dSgBMupfrh11R68Mze5mHrWenBzafnjXGJuJKqkxsv765+
eqqfrDQzzOJqXA/1coIyx76rhsweVKIz/4XBIzYsDh8sLeD+YqBVFVFB1uXnw1jWztiECa+Pohjd
x1xanfI8+DjnD76nGi2qeeNEQVijxZm59ove9I1uk3w4Az2zN4b57GPSRH59phad8oMdd4g4UenR
boVZ2I9+nx3cuy+fL9gt7HhJYDjfoZyBesFKzAadFgJH7rmNQK3K+wJsJZ/sI+EPzOEaX45ShivC
0cezkCEgXkX/InVGkgykuptT+eRuGQkSTLXAMaufscox0OYCQVkLEF7M+RGPQAFWuw/+uQQI0sdP
GTkvL9sYA2awqc3gBokOiAzHPLRPuZPNEh6WPvhCM+uEYDLp6p8cD3z4ynek5ye1FoThUSzugeD7
utbKGjSv/+bNtNdiioQEcjb7XB568fv2Gvjg5XloZqKhxp5XFZr98QUG8KjoKfBX0jsLNuKFj0+f
8Q9UXKEzkeI9TREnBpsOAkcvAyC5ItTc/9XJ+5/QwKKCEj52HS2M/B1mTm4LjyPHxefotvh2TvZ+
r1BC4Ie6b1h0mVoW0JSD9lR6vKVkLGoc0/c6sYJrQ3eoRbIsBFmbq+ipJCrLwAjxxvZxRu3jF4Lq
zhiIqyOpcLfeYSjLfkfWiVYuUS9v/maSwSlrCv/voaPPOeqc0IeJYEZDmRi7XvyPlY8jSKzQyFQ6
Qt2XTyYdIdXHJ0jz9s7YhSO6CeyoDQxop5lSNQ57IJYmdeBfGvPNhdSaLnhhsLW5ihMEMbE412qz
BDKMvQsmLiXs8c7XN4I9y7mv6NA1GR5HGSNGHSxYZbFiNDCDHFOeIKifJDX8jl+jtPEzME2lzSyA
HI0FZFj4ur58Ykb2cQhE4ztj/xd4+YQSKxctEckSJJfAOd9/ZIbWriHG7aUgaXkkXQntyTrF03WG
LlBm9ibIL+3la1j443eHMBwKXKtBTDDLaBDxHbZ/nJGJFdA5Pl9hfxyPttRLrtQibJ24uFKmZ6ET
L7HKk85TRfJQqwNDFbmxnMYXN2l4kJrb0eH2AoXx55N5CvPHp6w2sIff5/Sp5UjDC8cGOGX0lWE+
xNOS9Yiqbki416ePzb/xw/wQqC0W2hWJmgYBugNYuOhflu0s/Le3igelZrzWDcgSrZQ6Ifneytwf
971i4faaGyQ5ylhYtxqwKeoolm5xLSVs5j5HvraSP3Q18iNtQb0CjImAFXoOQs95i/CIAebX6wxV
OqfYsuEGue8CHkQRMjQHwVhKdESYgQuee0j3o+bOb3Mn88P5Ilv9+2Bo+nYzmBBW/PeIgbe3TIYY
ZkdFKlpwPpwqoHZ2LGonDUsnNjw+62CTxp748PtrNeQLA508/VkyPEl0Ne4iICXn7mgUzRLkrL/g
x92Buf8OdyzLJGjycpJXQ0X6oFT8QEmRqke8UrdlZ8rEy4BlrPiS9NFz1v/xR+XYJ/LAbI0nMInU
SoVxlX+PBmlLAV4VLFkcoFS432PXBjUrR+bKzJwdBYm0cSR+BoFmkQIM1bvLQCo/qzPRj94cshxk
FzTbYGqO2FaabkA0o8lWbkdH6sZuOpwFJlZoCk8qxnYTxK7qgIt9VynR5IM/mzCfNSL+pizA7qUl
b3I/lnFjQksSp3AmaIPLYxgC220R9r+YOtoFFN14JNd8f6ogMYBMoDrheyfVe+ttmeHHww904B4v
+8tiz9KcC/Jf/vwsBCwsA0lwDWuse9F1yISSlcLhvMkGXX3syKK61F/gXhjA7jn2m+LHxduD7xSS
1caroEISP/6/b9qovW8FJfQQfw6w49O7t+Wsod9PXJBHDH1+XILP9zB5wvrkOYMvEkKcuqUlq+N1
YOPCy9XdOV7+6EtTl5XpQceQpaprrls0Op09YNOPP2lb3rmLJFhzXzQW17z51GY5eBtneLdXTjBp
CJgNjIaroh1S/0so15WJGsO6TqAK3xHUemZag3V92jp6uStXAeA/C/OPdKCUnAfuaXHqRUNrIwY2
TvLPYEzLVHaMxQmmvWRfa/GosfJQRw2JdBVk0m8yKHZG6I65SezlW1ziVuXsWVw3bICG61OCfk7x
5zTqgFJK+dxrzxJo6v3n42knBhMEATVsdDqHtJgKgakNkSX47n+obi9n9SO/eu3pgKnCJZpVqORU
5lKsQRGwPAm3Qk3D2vtbNDjpfg4dsc2bCJUw8UCQUxgPh2B2fupD2GvfiEeW/G8XnR2Dw+VjvNnh
gCxLUd4UsHCtJH57ZXfmAyAYmrHbmL1aqvIuwKxzLERu+6ZaWxa8eQfIRsWs95hMNmxlnaOFJZe2
v8WK12Ghw/UPPMsPLlQD7dsWye4v5UrzlX5Q10BLsP8+uqbeefy0tm8UXStu/DeGh3WkHCfVi+eX
yyvUbHX3uqPYeQELZ2JRDYGCcDQCX3k3u/3a5+jmZXs3MQbPmpaELfkecNEvlmlgjqZQBFARI5Tp
ea092cNnVCoii+nZjLn4DP6xZ+Jm346ls4wMcUicugMz/rTNfYAMlOWT/vwSW1+ODShgb9ElwhXc
LfwDq7GOUSGqHbMqTMcK08URb8y5MlPR2bQkX77RL+DNXD8fkJ/n5oJ0EKL8MIZDwu4UJr2tsljQ
8H2ESkWpQTa60usA6H3dtrdr34MG6zEEziP3O3Z2GPpo+qSDs2x+MOGEq9/3p0J/PXDIboRg1Kjj
smQB5QDed3P1kXnjlQVn+EImEcpnVhBrgul2+swNeRYmmGvlkuxKPYMJVdlZ2z/9hblOp6m+ksNF
xStoW3H6UbugsOBms5cp4/27b/XKXUNU4SnKc9mt1MgTQp0QVSjNVNgZ8E6EHSpD8j+7vCi0gU6D
rr7L+BZTsjl1uUx6mNLanDuAiFNqDV5A3UTvZyC6vjavO9HRRmBrBTWxpWO7v0KXGHsxpJQZbU2r
OBLkYYLEZp84oCk2o4hfKIMcCUqiehoofkifAfm4P+EwfEw6dmqS1d80PHhTXwqb9kDZ+Q+WozQC
R5HiejZ6YicSRsLjefrRnlbcTW+Wx3pCHleeNbK6K2vueAxa4N7nvlCw23eY6jtRKaiR8KFXmdrL
9mxNaazREoePdvuo7UJl4JksEqjGBXOhjf1JXtgo+BQ8rZvfPbr++ugstUvanXjWOFhMSzRyKSkv
xA4YE2FRcZoGAUwit+beeC433F4MkFJ5eHKuOnQKO3JnpuOoFwEGdyyqQ3gRmASCat+zwJL5IvDN
0yULuOAiVdHa+oAvApvpuHPefCajr2EUUOYWx83oz1yXCTKwuCBWjGjthxtp2Ci3XRj1u60HYu6/
Gv+K7L2JHqJ+m+hH2Jx9UKozIAay0tcgMfEVGhC78QoqoG1PYGoWQ/VqZbS5kKFBfWXPlhcq2KTJ
ZSjojsGHPSwXFKOlJUKMQhs/X2bYTw4Wzo9CF9t71cBPLhdpjLoRmIEUNn7amExTT6w9FFwvjhri
fUfMX4Igetm+Zuzlu7plOhmt6N97Lo0avfVFkKrIo+shhK3mdokeKEwYMXQzUHIR4nwysUo7+Rpg
HT7M97ljX+6T1qNtb7KpR1HCSxuOkeqz0E+RF/mO02y9/3yxdG63Q4xHQU9Jh1O2r0vQI/St8zNr
HVzuZmBa0zc6K5CXgNkyGFpwEiP4QeKBhnJr/NmxbrOHtkQvMl3n4EtGeAfcf2RVljduutqNu8xu
Qr53C2B1ubvY0Zxgu+jTMShbntdJ43KdypSo0wzMAd4Pk5OhZfQe4u5Ltac4xQaquCXqeY9LEh0U
ViEc8AReP2xm9pE3ou2gQFEw4cf5fv8YXl0rLNpsUcsK+i2Ma3q6mFcZRFEb9jj4u3F0UdWk5cvD
d0J5fMEgfNTyRcVeArFo1SJTA0J5MgLzjV4y8cvvzxtCPxqqH6IlZlWYFChBSLHQnogyakcMO7Yq
d/9cU/dHtEpFqHiZ7fnVvstSJwwy3O3FJTmNdVoriyzWz6fV7e0f+w0lcpx1dkxXo+SSsPzyWyZN
kLDCX+gCH4ypN20dt7PjGNPEjzb2iwzsohpRrF7/dAUTyXTwv1Qm8jLwkEKWKvZ7jl6BemSO47Y2
Oi2PsLShKMtSabGW3ln2MoXMQdQfnSzsuiN47R0qm0Nvzjf54bBIhWXO/Gh0+U64kcv3HexaRF3y
0vYY8jttEK2nQ6fs5H53RkE9ky7f51kNPvOJyDK+mKdlsVKPMUhnEIxwL952ilekC85gpQNXowDv
gdyVzOM7AsTGcDUOighh2DVxrjMIqwsX39F6kP0SQ3+xNt+ozfBN1InavKlmwskwnk06nXYDfncu
Q0idjRQViA0SWG9kccde4f+4SxrehrO2kqooKekPNarB8gHqyrSN8Y4GQK+KySWJemfqlh4Sq0Jx
sm8MZIvykSqVYpDYF8fe3nz+WmcdKv5mY6bfjaVDI90RT57KWSE6YXfnX3D4t3gcPVVkA3TCXLwm
h3ZPtnzLYlP0oh7+FhaoJNx7mD1pZpyWEdMP5scJk1yvrr9eNFvxa+g/RIMuyypK9jStv9IQqXLx
f/XwLoa1E7oyEePdeCIjhEHuyQHzpmv3cjoOgf4lN497ILFRcCcW70q6QaoRyDjQ3aS4r8RhTn3d
gljuiAEv36S7LKjPcyjG20JuIzV8UuK3orbTDqSGmTL8Vv1F+q12+U1QAFrmzmwrj1IIffDIxk7s
QefrsZGxze3PJekcDbN310B+Se0Y1sYfhcbNLG9FwBAel1UBal9LA6zGnmGvutck/hq5omRhp+Qe
Qt29YwMN/yqrNifa6sbjMzVSnmXAuKfLGGF6uy5wc3ql4o2HHSQpKp6aNijb3SsIkjATGh3RGIpu
mfSmBpVe+hlPb0+B5CIrsTZaTG1wE4L/a3+JQHhMEaPJx/1ZWPhUQ5YvqX990CQHL8Riu+sGqBq1
SaY672wvx8HniZiXqN5FEfmQLxqomodLlDRopCgdLXtEOyWqZLG1Nz+1MwNkA9lfRitZLNJRkp8v
DBUWFDEU3gafgtzKBAkvYTyiPz8eeUnfNcmvyRtuj9kFg3hyP7TmFFlqg6AGc0hDEMZ5GcDhiq8+
jUEdUPoDpniapC6eHMkZNOoULxULPthz53K7kqdwznZl/mw6gHyE2fiacjBDM1MwCweOo5NmSb0k
FSIvZSjPxwthgu2cnLcHXQZCS8gijTcmymhuZbJVeDJ0+OvMO/fpGuvbx+XLR5KFHdG30hAWGMwk
yKLwNLpdRPA6P16h2M8EnCSLCx5mtRjniRP2AJWNfYed9y8yyhE9NFPHQ7GU2XB2u8UVdjc9A5mH
y4u5uRPI8YJrOxc/rhNLTA8z13ABpVstFNCLZ9fofQc2RxW7m9NKJQBksbc9cJeLFXL58RPsDr5F
xvNlVwb9SvbDgqxWzw4Ti36CbNUKq/o9NOH1m9gst3ieQwgGfM4bLd3PhfMDnmeryc3scwwbizzn
9s7rIO43EGvFmU4G/cSKA8jOssZ8acgvqzhVDEZyXTNUaZlgX0muO8V5sQ7vWiGr0LXElO3CpKVx
vyGlPJp2kkn4Al2M/cB1lERwAe5hzdaEKy1VppeK2firNv7/RJviCNGHJBfbC+eIdMp0pOp3qryF
oG/1e3+qYXq3IAnyo9OkPyHAC2S4Wgk4jfhJBOzdV7C2wtO1wujmLdOUrpm00HU7wVfmpYvPrjHs
Z4W9arlWFfwM3bBr11BlShtvoIapRgzVQEZSG4J1RLRc5/MHNYKDRCjFfOFVbSqs94JEQXwwCV2Z
Ry9E4i/+nhcdXaAbfwiqeMZRQB2dtFt/xpkUKVufcWEj5WpTackTuj3XKYZcyxLTOQMc7/XuSrVD
ZPEUupp6IbymZVNhDhHWtSAUsMbJnNSrUGskAhkJDN83OJyvtZmwQhEEyW+wglQYJCncXEPXlZgI
IRijAphMxxvE9WDz2KtwmFCRhCcBY6KtcQtCc7Gt7et41nwRGe9awx99ADtiuPMQuyK7OFCR70M3
HY9MNumFS0E/iuE+nwQar9YhQMCFqMQcshn9T9j+YYTnaP2EvacjrM51c1i8RlbQ9ATu5SOuOByV
0jbzELiRbYQ9l84ODJxNwwJ/1eQrv7lNYfw+fLkKMLTD7Yb3wtrszAeSbAFsfh+szJk91Yuz6QPb
z/RS5b6QtCMI77/hzu9qdLYg6CARjFYVxN3fEbuNDiOUYxt0DvyD3HCngurvRorX6jlRx/g0xOUP
o3+A6qHlcgWNLYq0CcLaEd5nirK0YeM5UxPbanKdHAVVaxj3rOvePzalTYPSgEaqF5xlVt1pmsQc
Kt6DF1J/Ub7m/A4GRGGUnKvLDHMWMJgzCSw/SirCq7iEsAYPXkFBWpN26G1mcdOV312oVrwh0BZC
HUj/Xcwl073eTS/SfpZpCAZCdWrwST/48x5NwrMJI1m8pBPsCtVIqZ2NAyuxUeFICpsR0wDOyCt6
KCE5Kz3UgMPQrmjQ58hwHUhI0mnhSR5bN4ecuSE3gb2fOpUva31MGDmZIjukaehz3OJ2fmAcPETx
k5DehSaS+NSIBUfHI/DmSWGGTZrMvV9GcpAkl8o5nRrQXx+zuZn+bYjtv5eUiCROvvg1YoA9SOZR
WbQG4Pr152umiizMXu2qg4I6IxT9iTVo7hadKEjLDBpB0SD49qC2gzG6aj/Slxe8/2mRQ9bd13zE
owYHcEZ4/i+4HTe9iybvkOE8h/5alDslYL9WqPSyUDMjkv9OGAeNbA3TjQONwqAAHnYMpZo8nFDy
QeaC0MmdDcaGIv1Qe8bCCgsaKfVQ6YUSjeMS1cBuuteMssPAwgDTji5WZqw8V8aQ5QxunGxCWV8H
eOuTwY3IeqkL/m4Rtl+FpiVDyOi2/U7Du9FuPIF4WHeA38yhmIAtNKx9AEBcI3lJ9MYYUB79c6nn
/o0TwWyCm/aK/LbGF//xI3NnaKLVlqe8p5KCqQAJab3LLQj2Nv1M3sdGY9N/56Vtg6SYiYq4rEzd
mizEF1Zgrw4OeZXkP4QCLw7bIIqiPygwopafv2dlQ2NgUED0fJ/KewfMjht3TtfUCyoQNZts67zN
J3yVell87T7/6tipgi7+CVEznHD+bkuqC59euHfuTdug/LzEzznj/Yf7UBXPXTvdimEnTOvFj3j9
d4C3O6N0lBI/fkj0WKnG8tZpamn7Z9RDTwzaWPrf5wzRdVu7X/4QuXVYMwTAivze8fkEqjTViXtV
IaGc1BuwGQM4awp7F54bFIh1d0nDlhXiCEk6k2idgfJ6gCZqci5EpYOVkb6Mmcw/N1uoh6O98AP0
guohcsSOGYKYTNeNryzxod+/7R/O1njeyHtHgfZQ8xIXD4K3HocJmBuM60iltFQF6RrtchsY8fWL
IY1qYPOOwR72sae5AR7xr1jKv4opc1nvNoEG4e90J5teNL9DC6ECEKpyB7xTlErzViLpqbqIYLej
c1Xw5W5XnEQOZq+/+gmA+J1jyMZ3pzg6Y+fS6Vjt6JPPWju17Mn0Bxe+TLHIMwt1jRESsMkPA1Ou
5djjqyZiG0TDLMXse4SLuTbymSKQt4GZbgomqFZnuVnyC8VD3cF5vXyO8+lsYBkNVDCyQpl4bisq
Hlyq/yhS3g++0zAWco+IodpVbkhf6tHsspQzsbuUoPMtL8Iqle8FSFxx2a04bNjBnGv6ARduoQrV
4HNVcSZEmtoFs+3R+ZpqgsxEg0lgpZttoEJz1Q2OYOsB8K4fAOnPiaUu2pAUgRyKUoV7RJ4LAJK1
G41630jOS47ir+9ZZIbTyu1jM2eu26AvY4SbRiAq340MwIJQ8JOmeB2JgXn13HyxsVN0+rzTuxj0
+tEahe6aDNlmqF3DcVDMLJviGdl6dYbzhqxsoEHQ6WxOaDUWHz7rTONZRfl7p480Doi3T9UW5FX+
yqUFqt+qVvvcmb5laRV3FyA0++0lFTtNXcS6F4ejvswji9yiCS5SYWgc29cv2hhUg/bRjEitLX2j
omqKdvg5lPmUzg38gz0MAzpsxD2qs175aE7/vSulvRFnd5VFkTOHfDoLnIvNR381cr8S3cp/tLhw
a6yaAluatKYJ56/r2nA3xtNj+p7yk0NXY0bG91DuCfVw0Yh7P15gPIOmr3vP9jdnz29HfcySAbY5
+HVEi9j2eUHcrJgm9OwLA5g7CXBf90n6ihHrmrTeTUAb2PJyczYemFzyOAJiusDOjwM3DNTlMA3l
lyW/NaamgNBGsMw+47HzLZgS6I7MP7LkCTq+C1vdXefoNyIjPV0EIzfDL3wdc2NffXpFkzgy9KDu
2UBEFMsU2s9wYXP7z+9hTpQ2iGzcSO/eMejVzHvCZTVeN1EWCVtUdE7fnQV/rTuw9Rd9Ta00S0Af
Co8bJKydrVXGSW+6Gx6+r05gaeb2DbSiKRbYjwJBpzMkUivYnuDdCLDnJgfb7wiaiN+c3L0MIWIB
VdWhlTpYo2wy5vODtc6xRqganAxD+V9JTuY0dUMK2DltNN8XVpPQmrz8p2edSYLSy2b8Tkah18ry
rOy64lRfY1DS+2CG2IMpkWg7ddEZ6RUoydWogpcvPF1rKpdis+nX1M57Iea6v78hZb1Nrx8sen7U
Np8Zo34c9UezT195FqsaIlcTakatmtl2S/JkqLFcDXxLDZhFQdG2+E1S25bIo6KF4JE8FPIjzxHG
hWjR7MnPHFrzh6tKiYQrm11IhKDq9jH0iJn+m4bE7wnzrAGw8CskKVz/q5eSLzX2rqJAbyPfBycf
U8KM8IezuJY6IsmhnFxLLI13UD/dSeWfPXT11y8YyF7vfWgb06N4r6NU6SWssE2UJFIjQFR68FN8
VpIar60L/jFr35DnZ2YfvrydfqntpxFth/NmGL3J/iXkgzf5yQgv/QkmoUUDj6vADBCV2bnoaD4l
ki3YTSyaourN4gtmiYd/ogyNtybBZzOhNLZX/O/eWHkj3Svs2nBHqN3rknmgQP3TgXwVugSJTzZh
ScOfzvpubxclyMEDFEe6wZa5CmHV3sBg3719fuxwZIWMe6QgNxUtocEHENwGxUlnAEDvPYxjDoIX
zVT84I6BgpppIb0rt8PW9KrF3CXYITEzau+PyAwgVIJesmKqBIhQuFOixZOAstkfO2BgLdnyHrMp
ArWTp59YZxcPkPP6lwUACeIGy0wuTR2OBBbO884xAamcJJUMB/NmJwomfy3GFOI3S+4sNb0/gYuX
5+Ef6UsBfoU49B9W0zTqBCCx2MWSkrXVax3EBIuUJ9Xe3syCRcLG2cJElG88r6QE9OVzcmvjqTuC
8mvJiaTuqFeEIbg0TCqv4s97hLnSlfXqQ38dbw0ZNppjYAo8cT8U85sZLvQGkkIGkrmPI2AxObnU
8OyQZCbgFKTtjX6WlMoL/IJnseVadu6zPJWMxFaT8tu9L+QeEcrcCL2AylmUoDN+3OCM1BcNEYew
fJdutdys/nKmyJAuYXeDKNLdn5uo4OA2RYwNDG0+V/Zw2ole5qKcwWYyutwOp8xa+BAmSCtRQAmW
yvVjeQ9DIzUfkBLbvlYhCFf8kq8OLFgzASHR+vcB42WsvbIs7HVLWEWq2DOACMwBrC5CcBMLRl80
RJ2PKEHXb1awGJVdfjmzFHAmifPMkBVlzK78ZSIOY/1F3/YabHnuI8XcVunG6n2Gj4tIcu331aII
iq9scnl0eRWChWW+Qmg1O5r5T3WQ/2ZWNirt0bIcBwQP5AhuBy8bzzcB2zttz99fAYOzC5JujUTe
purGwDi/FRwfyHhmyw2DjKUvUsY/3hLtgRCFgKu0DRKZivdmUH4FocYwTgKctA21EFXzyJ75YsMr
jeno1g5CWYxBm014FM4EkgR/MxURHjUCmzMeK2eT59K32Sh67nQEBnGLoctLfkAvFmNX7lLwmK7D
R77wBAB5avw3q4lgoYUsRqihNYpHaYlAKTOwUYTd0VWZM4FSgKsJztcC9/hG2HvFemXkj2/KRjgJ
MpnXK5lft9YWdEQ+kCNvhZ+R68G+iIbEVF23eddBkXfIHRn9Eb6TYXkfc8GVRD30jP91gi5jwVSe
04cpMS+cuhVwbLr+aaRYgiM4d3lpcbuVmn5ji38LSMRB9xY7bILADcFpXoN6qQBiLuEsAO3rlRg9
obyN0EDS5a78gcldAZfUVT/B5iGKh3HQUuo/wwPK5bSkyUdbCNEQtpvSS/79GthGFoQBeqHHSNM3
oLmENLqXeLRNz0n9hUMHez+zb3HWJU8d0oBjSqSxXGDp4LYIfzPQ8HdtLbJTyl+kAddxjdZ32wap
N7mma3kKWImrFVmMkWjYoNix57iuUBnbz5yzjSl5eUuk7vYM17V7LTM+mQD0VgTJyhz2FkChzyJH
ru2LQ+EN9thE3M7RXdUTKwueeP6MXtZbICujNjERFZAmuv/gxWCi5+I4ysLmGbH9sUYHdCGuvGUw
M4omS9lLLb/HhZxpL/pdhqjR0RDJI99fAZfXrDOBdqF8+aayk0EumIYh/e8BYrpIPVMAuSdkZmTt
S3wJpubtf8FhiGp2IE3BclS22sx9BGGo8drgjuE/kvPLrZUSgUgYKtKydgbZNkq6J4dO4SVN86uH
2C7ou3EP9grzZPWQqlHrN0TI8ZcWTLnqEBoiAsPZdScUzwLlD1Lf+IGorsHw1jR/mb+UTMlEVUwN
tFWJKAJhVVQezWLn+DbnDfTGnWUBrBkLEkERtCtWDcW1CYviXD4mqpNm8LTvudm/TcRcS4Tc86Kv
08yT7jpznYOzCfpO5Vrh0bq7rYCi8h4sazBab+OS11mD9/oSU4SOlmGIlu+JY5QdkQlA/c4YXbBO
eYoHhffB0GYA/NkIBUNfEmBS94cleLfYjTjvRGcK1ln9ABhSKm3SyCjYWcdlP/wJl2ziKvtVGXhM
o4wUYz7/QPQN/h6AVIO1Q8HAhjRp3fF2svb/kz/L0JQk801wkt2e2iiLDV13MJ6YsR81bvhrIcZP
BCa36cSMrYT0bkORrSog5aZVP9sPG3tyyDP2PZ5X1vnFb45lw0xJ/oRw7rUO41jjOxiZt5UC5IYQ
xe3GN+M2pg/SjzssA/9Sfu/eplkqf/Jnaru+cOEXVHB9HCwDnojJzGAwbW5eTBnAhGiAfpV/L+m/
PnXbJCKrbjBXRjZxurRYkXMpovCCuCz+wXoYJxpcEJnw7QyP1BJCtXjkSQQ8uwdi2wi5GlNyfgSR
QLsaAiiAEo+Bnl4KfvZAO2AWIq0B98mUqX5G39darIOF0Rbvh18SisdqqG8r0EQgUPXXmUyKbBI9
cE0Zx+n1/1jOWOIc9NbfhZ+MjX7xUjP2Mpb544mQCECLNlvqvmxo6lLvKJiSK7eQigwepkSfZQ2q
oHSUNbIrloAiC3BjIyNGBjCvKyQgNIeH8l1P+jsqngGPdvR7yvUUFTn0WXsZif6w+Ci89DrHIrF5
+jNv1Z7J9DYLsD+GkCMJ/oLM+1AA8bBMawIlPKSMFc4DSkHG+gyOR5E9TVVB+vt3gRa29rbGx2zG
78KZQH5Ra9vOe4KncT22lGPWGoQN9WM08PAe7CLEURowJGxyjjXiacwp4wBjs6QADIGvDo/s1+Wt
eqd4H2wFJDgYMr9rIjl4Dcgv1n1APF1+D6dXxXn8GO0x5wte0rE5u4Dy2GN5cAuDU/NihHhQ8U+c
kQfDxGJTc5eWdLCMUVbz3qnF5ZfIEfJ2S/qqAWNTZDSKC0r0NgRYiLCWkgPIHSndCW3ZZpb57hwO
7ZJcjpGHr6zYeAH0vXsZL3DuiBhPTjFnNXQdl/xPGw0xDMvKR6s8DNcjLI2Y+ljA8XswHJdV+p0n
Cx2Riv8xVGIxoC5VcM5dsi6G+VOEeVIAle9m/an8OyjHrevpFyW0yDDa4Syirc8w77GO2oKhvDHT
bxOLdIqMPbrjxbPDEnFusfhz2Q4xQDVENgbiwwi1pYOAlFphp0wFwqoT6epC+roaqKiekeiS4cbf
bjnFW7uEe+Ftdy4MK9k2ay58iqliwUUx/HkLzd6dw6Kv/Tv3Jz06BefJxi1F58nFjXCIZltqZkW3
YrmPwsA/PlhAa2/naStZbXVExcGWEBl9H8xehGND5vPHNpQXe9/Cs1SUUFloamPjJlUYnpS5+IbW
UoNCpk/XxNRUPlVY3BHkt9Tod6afjiqYVelhk2RAAI+r5VJipbD7Xq3eof4DiCHrpBK+VqunhAf1
kW2OcWOWk9rJ60JQt69H/sgjfGLBdaYisSAH1z17kWH18OknJWPin1w5fX1IC8QX+UXlLx/G18xC
sTxkAcxT8MtsQYgueTtDCz1CaVO0pM8+8y6okuID+wpU9EypeUgs7Miq5m/voYqHc/BgUgcu3hCl
uwzZNLT3AhxDCx3RAN45hGW4kea/YNrmG4y56cL7QEqVMW5QNht7xyyFmrzWJMj9K9hPNsbXGdfX
+41cSl5xKMXLocxj0ezYbM8zoR2bfafgvErWzctt0MV2wkk2erRdBEzvYfwnze8Nvpr+y1++4TFk
dOQvt3UwzsCa+F5NTCAdyAYphP1hw2ChPvaIzanfEuNCxsXOwbPtVmJPz68yJ/PaA9/rRJ9/TfUw
DxnNNWi7mYI6zX7Cva2MuFm/Czes7bo1X+MNEpVLWgs7bZ60dS487SrfoRHTc54jP9kc3JWGjYC2
ArI9wsMG1+O62isVDm/q1SGIpLngpeGX6mfIDex8qS+kDPw+/clcAbilt70U1CccZzKrMoDhtbzL
+m6P5u/fuMVkdRwlz4i+T5WYY+yeolsWSmSWTJU7CfjQ8Z9PGWw6/sYxXVdpgJPJ/vlujPOz6dFs
xYEYM0GalSPRCa9cVj7SdO0ZnhZQ4lkSVE+TKGNgs68tmdFOFLfvY2LX7JmKFIMGtD9fP2CmMmn3
Eu2g4lugmuI5w/o+P2mMupNB7H/CjjFhr5Jj7cUxW4ggYgRlGiBu1MV2Zd3aW/ziu0Y24oyzIRiw
MwK0a2aFj4Aij5a6y3OcV3GzvNDk+t+CEoUc2SbWyUp+e8+9gbKTQHIwN6I6QgtPXqYHYcwClIOq
VYsHjwIlbXeUv4KCGIdNDcMRpoEapIDpBCf1H+jeseXuXdP2KT4/2PiMdOKRjhtlpRlNk47a7vu6
vtX2kSDiQEsgcS2qVCVy3tXUrRXYYGpl0z10JnSaaMZrrJ+JJ/yn6YJCJIP0u3ZToopyXGJaPDd/
k0nrXSMuzLdc1K0M8cOkWb3SzC98TPFpkMNhk8geK77d/FOinqQImeVgqBb7kuYFI3VGP8fGJGaB
tmZWvj8z+7emhZM9iycLgu7BpuC8XwAatYI14FuPKC5tpYKO4rWZRRMhfVKfIg0Dd5mJL9DxCzqn
FN41q6YPQraetNcpmLeG5JLVzEVg8lfpVECiEfvzppo9DEokeKaWm01pa7062UgUE3v2Vqcs2v0A
DvcY3KzV7jy3vyE4DdWmZa1G3oLyqdps3RxroIkKWXV2ooG9T5Ha0JaBFeCz8grW9lWz4jFUZnWS
ePSnRWBb1v9Soa2njYaF3FGH9S5a737ascMrOzzUHKYoB0cHYqVfg4bxGqEVdm1aEUqQtuXW8LWV
lWgYMtTxxTHlRyL0zoHeH/CsZM5dz1uruexodG9QTBmU3CbR3KnXj79xWCIEgtaoGWyFN0+qFsEF
b3uGGsyn8EAmcjFuRYaqCAS8Z4YkoqyhuEFZ2vIfaTJNG33sa5NojHkmjEFTwf4lLf2Vdc6iTHuh
jIMqR/LxMwTTcMnHTfTJJwJreOTG2GMvnY/cJFqFygBCb6C1uIS6Rp3cWeIcDbNbJ7ioxLv7edMV
5t1jFyRF0uJ+mwADYHRTYr9ikhMjNzkEJPISR0xk+4jaHX3L+h5ubO347q/XJS/vmIbf/Pk41VPP
1sWvJqq9ondv/8hUHxMrQEgmT5eFn/aaau17+4laLvoNRwwvz3lRW40PqCIscXDyxO0XAbJuhC98
b+4ZNCihHo9LDiS3ndh0RXPQ+i/vTfu6rrIeWAmGxz91kKJUBNddE4JJXFJh+v8vwJARVh9Wq4+q
VUPysFTOT25DbRBAttq0hZtXAgL0XmJd5bm37F/ZPp1/+4AbiCyNAsYpwoXznD385dUKuRrg98l3
IK2C7lztFYJHB06xZ7lVHX7rpEysC98rqHptGKjsx6fepxQ1kfG/nPEI4VrjfTCeeYVy7jaCAsi6
mQaQt6/l/Nl8Tx2L++L7pp/6zSTHYJVBq9gbiNBMddwX6zSw8B2tOksksb3I52KycmakMfElRhCC
/s8YA2zzy9QmmTCWFX2hp/YNizqlmmr3mcdtd9a3KvMy3HRzxMbSYXZG2UeVDCtb5I/tvOnzs61E
K319ah9Q3OCge0qbkd/SEyaDPqrczqHPFZPsJFY6Qlrxuz7FfP6wEkll6rAsBYcFuO1pTjNjEXRH
wJwA1cZntF1bY+RF4vywtmhEz5di2nS+KB51UGQDCk3OdGeduc2xY7bPmG1wusdgDgCbwHorko4a
82Z6+jUXnf3UJ32bUczTS6B3WjfZmIa3yrsnxnTxqxRgLFf1Mk0ATjv8RHiOovGUWo54w/clrGrr
N0TBQom8dNKBSkvSP2c994ga85bNNpuQUiGKgELyTciPV26u3XiXtbZrHzWSE/NVR3kA+ij9Z8Gs
GizXekEE2vYB/yc55bOA8CrU/IIS+/cJO318cctrI7zJQC0wbOw9r/Kqj7GjALAQ8+90roSrV/NB
4ru2C/7kCc0lv0W3Ue4JfqWuyxBzrFdFa+ecvdKERXEajd0IDKySEU9+BdwMgWdoJslrL61S1KCU
QNostLNyi+/8JpFN8RRPf6uFYv4gT3EFzJL6+tAUW+xtykQ5iMTiIVGb22YZ81W+lFOPYk0R/ly/
SxXmfrYINxHUevSBTRsxK14WfEhbKyTdlVSVA8dAW2sJIb/Rliff/dgdey9wxCyfR79Anl8jliLH
T/l6VPMS7533A1xc113egIMAghdcRg4OZLPVUFkcbBpaLhlt0doj7/LhpTOvHcwuvRtW++s9Vdjx
CWAU9SHes0ZE2LnPTS5Q4ndH6rOujk5DxXDAQLyCvyuIsifo8GaSHq9i/lRMItcKhzNbN8O504od
ahovb8YLfagz0eSOl34+17t6n2Ya4UjPVDY1tg2zQ7oO+72KzMo4ZXJnH/psl9WO0MjnH8Q/dyN+
r7UJftsXWDkeVzHqwCy+TckuSYLCSqUoVPiRu/ZAQ9rynvyWwn7vRxGakJdCTO/lOegXyVw/Lks5
NFJtH2qYXkPzhhoREutOCMwg/hql1p1G01ODtQcdqRRQcyX8qqBGN11FqrXoBiNGfIdlpVfYDD5l
j2QEDi9NhsEYIx7g1V0IKE1vpjRiD9Ezhpm1LcnM1lm0jOjLY1ThWg7d+6SQoo9ECN1PdceZTOHm
cuL3BydkZ1PW1bLv0Lu6jy5DtYwuTG1W7lEbO2dhH+r20XbiuDCx+YyljGu+i5xp7bwLZJ9JZH4Z
FgERO5vQFc/Nj8fRXkAg6B6xNGzhr4zEPS+tNqryKkmjVv3gNHGB7MPKDvTJSYNoKTKeDZlFdKnt
3Oj17mqhrHMymD6knl6KaxT+MSYZCZEhjhdvsrC10lVCzbf/BEZgoBuQUEiyplYduiXC11CkRf2V
nJ3eMd2MmWrhzmQMQVgNNZ9g3l0WrbIznK/pl89SLVtSjkIc/Qfi0O53vco8hmZfx0aSxGLCziZG
hRwVy5wopfoM/Z7SzhzgvYZpeCI9TeqbbIPPlARjCqNYS9+Hj5zVWXoteFGW2IUEn0kzTHS0layx
ltzGfJ/uKYUT8ODddVmRAnp6hYeqE6hbgY4387W5iVu7oFlV4l0bfsVS55fxO2FUqRqbLt9s3PMj
Kk0Loh+dtaCXJhRoIfZKuqS8DKIUhj8EhdohcgQPovCAvvBkwaOwKt022QcymTRpCY+Xx2MPY3FT
BsJne93dJm7LAhZGRMAoDNmgQsqmGitYUxpI/BMG9KKkBrKTQMJsCq73d/1E0DjIj6BPTZNO9frm
0fGqDLaf6YJ3nbIZu+HT3dHRVOlwkCux6TiFDpvazJESBHVryttmuvRkKYT8yF+gyK8Pv7rvL+Za
qO4KEfrrDENSg53jDapgSFTdEi0GDhFLCvuaS7HqHNvlagAlYcTWlNAAqgrpSPUVOYagZE2K0DoT
AHMxqQF0i0UWWgQN4/p9KEixfzufCWpVHwHPnCwERt5Z3Ad8ZnE9izL5HeqcHA76vzgNnWZP948W
TxkCrYXfC8D61cuUD8GQDDVTbOe5spNDn9M9GVxrD/1QUewcNZD4WepYHh20ZlN3mWU9mSr9a9Al
JsDPszTD6sUC9aFeNAHwj8EWkJ4pnqTh9d/F726UyTAvV+jox9boygIQTNaTx0eJCEKJ2RMDgK35
xsa6JR+6rGEQXDqtnJ1FzcAwGPK514KhEAfyjcCxJYkeK6DArGCszlL4109kPuSRalYD/+Z9QGUk
R42FvW8kZvU3PcbZOsAGn3vuX4D446cyDm/syc1AzkMyn2/NSQ+ct+TtvpcoX5qvN80ZttptRRs2
g3vG98+gjOd1uxTNNdMV1uOMPSVzejuBb5mZTe/hMDkkBAAIWfvy9n9ndDBruaIHQXMoV8mT5TBJ
fxa0Zky0AcjJ/u7wJwMxhQFIO7t6R2csvNBjzsidH05ywT64PEMpH0ORbxLwpEbDXP9i8Sfmldq0
OZk9dVJkKTVqk1lTR4TZBtx06pIWPOg7GM1o2dauop4vTCoxH1VkzZwzvO0IQC4IyJXxZSxb4p8Z
Lv2/ceBzjA9n/rNBvP5+HiyiVZtKpK9ZeuhXBF5htfVHYKoJCMMPE1XTgZTaZkepNdDVTyoVRLpg
D6CL3FTP4VHvG2bdW70NCpNZUY5FDmwfp7L2L416foz//X+mDq1KvsciqSQeLXJJEYBakJ9Uznba
EVUdMnfJ4Ul8gBxHvvQbuV6ZrkKRSpulMyQlf59GINwIVetqse06IWS1IEyeL7rUHlScbyxNG2+l
Dl7tgg9d10LB5E2C/r5Da6XZ6nhPUGbbfO5CVjaulstP6C50nGjiYMcIi+e3D4dZ/6aC4T4J5jDQ
LDV77clkuwRD3xQab0IEmaqDRLDv91/xr4LB5MOYL4x5JQVtCKeOrmANamDxMXHLy9/6KqjVhI3G
bFtZ2wV2lDDkaI58EDa2urh+/obJzKH8BRrYe1YCzSrciU6FABjrafeI3mH1PX4DYqFY9hGpHbDs
Kcm/nswzdK6vOBfgj3L6C8O1w9EcCLvvkB8l3JnRs3GHvHjAqeF1wenOZg+G5wfLJJr9CS2aHAtu
A54XH85WC6GKS4lGF1k5A9XvjI50KOPVN+c3mOQjDdtFoucIbpD1WZZ4TdGcuTKiDFVqMi1OMO75
zVr3HuscsIL4tzz977yWnBLfLm79xx9WZY2OfnvBoVlsxCptdGHDC8JYjuLjOO4HMcQC1jWSy2x9
a/HAJn1Ci4dF/bYWfTmoVwX07K09QcuyKSMc4lJaY2pjPGwAVJWvwqzWhvRgBQ2tTM6ZVQ/kXa36
7ASSCfnsOWGUN0tuPA71S5fe3/nhWJ+ZKYyDVWr3Ivoa5eTbC0T4S26chgveYfEcZJ8lZmmY7bVN
JZU0owHxNDVHfxNCLhNWC9SdCJqg97IKaAwCcaGv4PBVlpwcDx0l+QNroEAk7cfVJZOmXLxMDpEB
rh7o80MALXXmCaQeUmoXt+NqV1FQbsw5Ati7JsHsdsOLJoFnuqLRp5VwzRjACrFkgBcbg3+YpSBB
cR7UyWwP+jBFDEalsUwXioaYtd7pfR40y7lBmSErWfPtQN9r/QG8g/TehnH3lrw393hSK4IfOawa
ibILwhI3Et1jDeQZ9ACIhB4trOfqq9XKo3ecPxrWcudsMqKfnKA7MtKwk0PXj23pQujHZt4+LpRc
jKQOmq1/cCaNg5tcC77D0wBQ7ZGxIhVvq0LQ0xTQlxqDIa4m3VnJsUvIpRNhFwW8THpIDZ1An7jO
rqbKhV4pAZvKnu776HQVwQ4JyIdBlLHM4o4DjjAXptLpfOnE6Hci4HOKjveUqRyC0B0oGSxjInAf
U/7MX6+cxNX09OeC/oCxuxX1KgL9w5NTVb3qX9UWxEY0uDbTVtbdp123XdwhAwLXfBB3IY1hsUpM
CyYX4iaJdVLR2g1Fzig7qtZM79uwzobjqCCrXILYqnjAZb53GAY5oygjAQny4leTd8ZtP3SrElic
cBEcC2b7549RZf7RJsgnsuypceRDcV0K98eXo5tRL+0+joz87Js2giU1TV+hAmy4G94WNS3DeCQ+
tZwn5J3CELdfmFwtW/+BWIInh5crwFRwRZ/WrrVHJySFzBF0wpmgLSIBmLNeO2ZUzrIJx9Drre3h
VQwlzhW3La3saashcW59Av5N1BduJQTkvd4XqGrUCvp6yg18NGX0NBBoOuPIlkaW28H+8iE8rxtO
b4vrDLcTfSV6aboEtLnSkjlyIm6P74v2q/8P83QbhDYRx3koiQyXCIeWBTwY1eWhOk5r05CwCWae
lxLq9iODt8CvjzZEpELgllcLS62HJOrkdvAm9LvuauQuVoACi67ks1JpPx7rLvUL7seX7i214xvL
9UG6WcMoRWZez1iLzmTsDhtbMLSiNPkX37rUk+IiqbFzU/53BeizkPAeLfwoz6/EP3OlpPPYqZwX
ney/C4loO21sU0z3kJdgQAWB3YAhoK8uado0+31Dkxkl1HQnMR3b+DFHscKpcX98PQm7JovU+Vye
sexq6yPPq3iXgEFbEioFVTkKm6liJkWOy/Ni6jiRYjkJ0aq2Nc25tKSqt8k5fLU1nkE+nVdSQXhu
n5y9JvWwIQ8rzmxWUy7Qwdvqn3L62Ue3Gi+EqergUbuMWKwXpHhypErnvd7BK+3/ySrTWa2r+ADo
9JkXlZ34XutkS6LyXO+ta/FHEZFvauYZxcayQfd1dz08JiJMuwVzPetVSL+jBF0cecnZOBQ4sRQF
W37D2KHABi8l5SB3vRLCuR7WYcU7LG1SUn/9O2U+kmheAJCCzQ/zx4ddlqR2xLWZMe6vZe2OWdrk
8lTusesaYDnyFZeSqu1z1u+SPJJPK9H2xL09/zGtmJDpeUpfDQSR5lT9zPQrwXkhX3U8oPPHSJ8r
5KFSj06MNUbo2k15xSaEOLHAplio2TF8jE6ftF3dKNwnhR1Ul8+1SKGh6akrbMUaC1T35E1DScXB
HZkUpCQ+i22LFguWIhlyyNYTPIVqylzGWHHilPAGEAXkGpJeUEC85pIziyTatmDwweTXYEahR4du
5IXjQchklGB34Kyn2q6mH+saJlnZPHekhf5eQd0jeV7BolfiRHHa5HX0a4V7Q/45bmqO29x2bK+U
3eO5d6NJCZxVQkOBaGtqGYMUf3GA9lMQzF3bOH8APW/hgU1a+vQFujEM7ZbkfA2X5zLEljUHYcGj
+morMCKtlHSwPO23XvBYhgfWxKtaTxzB+pjMpdZin0YHE7JAep5r1rweq63a9eAoGX/z15pk2xXg
xjjBML5csrefJqbFDojkBY6j6HGj4akOUH+q7vJFfYYHthlnXG6SkbXJdaa7SOgi5Qr5jGtouZ+v
2wzC/SejyQS97ed6J86wfI8eocklA+2lRUnroiO+PcmbNjxU9CDorsnipMZeuS9KXvXg4rl87GSu
wl/wzO7neCW+zUpfez23ppNOjQS0v+acEUJfVPIKwWILGr1RQHPi1ifxHhiDwfvsD2nG+5AjBoWc
VxiNXFSlMbb8m2wphggDd8858DDmwnRHhyXOxNiDNGy0UTAQ1bGoPwKOTTngwbqkwu0JUxMRQVeS
Xjc6TZVe/Yg5ygKC4Diw6W7p1bthnVg41nioo3S82msrC/5dxbTk0Gfmu07XjTz+eDgKmm7P2w/t
IoHpDOM0jxi1q+qUs/ILWDDYclwkwvaEBSFH0nJEzximK9PwJfbcbiabcTodzghkftbWIdg8ykiT
dViOEFBWd/8+evsUzUUX2AMYKk0xvnjDynpDZVCJ7GUBtQXaPyYxeeMBx4MuYA9H7c5EsHoj0lqe
e1AnW8SOIZ/Z60ia72ipudLMpJSInh/K920sFAmVI7sGr7vmH9bgXM2281PV1if4ARLpFwSZWlWr
pN38wDLfdMnwRi7U0ub7sz2MderATBnV49VYaT5i2c0ybJWGxH3Ojvpy36lFSmeiCcvLNaWd+zet
J+719FbHNYNtH6sFZp3ogmshNYxWfjejrwBZ2GOC1EfotXM1JfGvpPwy9TIc9QR9y6UQ1tVy+KKS
6JbXz3POC6LIJT70/+1P11cffREl6wUvYaKMXl4Lz38ZqYB759/oPdKmWr9d5GF5csN+ZDO+c/H1
6GKo59/JsyX/8RLlojhY5POtMp4MVVNzFX/j/bmmlVqgAuQTDRN++tq1i+RMNkrh0npyq1F4hzXH
XjyKuTqQ5BAERzQZN1EBqY0E4F/6qhBygAfpzj5TyCmkxHaO2AlLa1DbODTqL5ZswTodK2zXHXHs
jPHc/+5UGbRri2YCX1pOg7fKZ0zjOppIDJrN929ntrRGaY7rGMzLzWB0ballmXSl2UKi23CykMX5
Hb7XVc4Da0Gfhn9+WaulwNCqg9ofvkpraep5ORhLqZ0IBYgyPXrDXvcZAPa00jpzPyNLaH0tZmsa
dByYDpaQfmtgWkzLY6UU6eOUTiMf6bunV4zUDjTKPi6IaSXnSwQPsFSM+JDvGbwZlPaLfLB5B/cw
MdncCORG/gfmXobL/3QfK5plje5s8/M7fR6Y8xXQGge2e5WqcfABwLfo667aBniv1wy9pH9AcbS3
kydSBZ8UVVFhKnRDNxwgCt7aXj7iaIUCXa8WUT7WBJTOyUag3gXQM2s+3g3tKnr5TuRivbg7WwUs
iHlWMCwXX8Nn6QDMZRNNnMcNWLjFhysH4WbuThrKqQuVOthNb+QyspgOuc25eD+4c9xCB6Hy7Y79
Hebu1JsxoRUHrWG+2z6MrAkHce8LwKp8WFv7r/mY+PMeP8i78M2/1e8pEAKPfKXqaQMpAVPGVrRx
ZVhEqN/Cb2pcaqEaBjLj8RuKUi4uqLa1E2H/92mOSQ0ualTIvjAvnHTv1ej64Te2tLWdtq2aa+SI
KXioSkQympy2/qUT/C7l+27sHjfKZ0mOBQqsQG4vkaxTnqNBKpVI4qFvqBtQW5r8Hqfgi8wpTxu6
R3D4moCDS+VHBUaOU9cXvafM4DoO2PqSsDXConDIg7mTA/sKZms6zCsn0wqaD1W197xscZriUzRR
JjwfFowDe8gLPd76LIEdKUrV+YUO2Y4hA4003PSSSSTFcn33tBup//EOabHWXXJNid9ka05DhFQT
YdtUDTPhVN5MVQFw1NWDY6veHFAKLIMtHhluo9SCKeCEBPaxQXjGAlYimOsG7DpOUZIbnu4cUn7A
HIMjdfn/CbmfgGtA1M029SoEsvKAT7Lm1ikOBPcNiANJNrLKIlQy/hilazZ7mPj21U7PX1hRFN3A
OhEoSGo+28tTxSF9aQpxG1soA/raubYmVdskrxmENxZ4cEW4Zw8koMLgF8DG82iuUp1eWxK4dXrD
uMgvbUzcFzSU7mPN1zT2dgN96zDAS1vQMi7VlEelsCj56/SZiOj59x4tpuvV2efzNwD+rQgCr1lU
PryFFNpNHJLTsu0n7xKm9Hhfx9JAGWaiDcuf/YGFp7lnLLo8mR2xqMYI0IVO29ILK1zbaZzCqqVa
kX8wpseScp9Up54o/dQyQZ68JJHQ9x7Rq7iKV10R45ZnYW2AI3UtfNGTQ1f2QYPRaz/Ui9NBrnvC
Ky9ZgB9hw9zmWTWKc303g0B76SQDwDc1RoEykuHobeanygzQEsJNTB4m64210FZJK9oEnwptQgZE
ABt6ag7tddfHCWptaJtg+pY2hKBn0i+b348gciGsFddEXRffyqEtFF/4C3aF5aZFLSlD6l8/Girt
LF9ylRd5TYXgmltlGh694Lima2JC3kJuyjmmt4BDT/g/mtqynwQ2C7+b5WGW2k633CGYkUgSYUXU
FeUf/pjFY96m7sa4I6XvXmyQ3i/Az4dQoMcye+a8lMOBqzUdQnycSCqoM+zMSUYzfXmRLqBaBXs+
bxdElEzY61aBx9cEZm5L+nd9ZxY/BQFW07n55BoWpLDoIqU8YH1yqPahlp29l91Bj0a2QDzBLuRE
/TPiRFk9ZUZjjJi8ZOQqnvomdGFPE1w/XlgC6EPiLD16GxbJTWLK4HHApZdV+qRZ29vn8H+xxW9C
zaW/7DmaifQOMN6etwocK1Yydv9PgCR7kNmwHqktwuhXJaDAfh5uAaztxGQ2WksoonSHhJdkv6UM
8mUNyRo7hylkgwwRbD6zzBUwFwcUholX3oq8RPq2mbo/fzeApdWUAaUo2BULlbjH6S8ESOXc5p5S
L/BKklq50CecPso3lVNCHqIiyalP2PECaG5l4c3hffeMb46sm7UwxjqmTm4U8deIUT/poqe8H+6Y
CbQs3GpIFv3HugDf5tSdnt5MWzzxfjrGAjFdH55ucwEaQM4+sALmv/6JeVGXQe15Q3181wNchPwS
4choj76jPKzeQiUEIojFUwefrN4OCwNMTulgHOrhpWJZJ4/DjlCBLrIOqrNDMZiYYhbZiThRw6RB
GSugzW74q0zOOVqB7MBVCyhVuwe6cTunYgn05+XETi5KuhY2U2MI9qY603dX+1PutiU55o0YtpZp
K8gG1KO7Zt9SjT/t6XIXNiA26q8BxdMz7AxBJj0pLNhBruG3cm3QX1HjKlwZ3YH3dYEyaocznZxp
OG0jWIbxr7zwwCGTV8vdkZorj9YsCWIOs6w7KX9/+9WTlHjkrxIPFygXYElTA56ITMX252YWFosd
F9SqHYvzvcdIg8ftjra0jBC0XAS9KtMTa+W/g2PDCfjb3w7bYW2Mtp4RnAJ0OBQ5WDcOTCjokdY9
vCnKyi4x1wMfJxVrsCkIrIzXRl6EUz1O+jJQwGYx8HfbRJCao1UPPKoegtKgxo2dgjImUQyRxuA5
oBpmTw6Inhdb6JUYyH+4DRT1r9Z7qcx+eEDowKHTNfcDhrvGlx+zPh2pEQ+hB1AygD2Y9o5HhTDd
UkN+jJbGM743SkzBOlLo35qKDslckg2sQ59mjabrEASo49adWPpn+u6d9n5+Vh1hMg347x2SHtlf
n0DAoA/vB7+0lt3Ast3AgkyJWlgyPozIiTKAcsm+W7Enb0IuhK+GM0yXtzugM7VpSIyCOfoOSyBa
J1SVqSW/cOXihqXMvSl/xcLefYvMKRMRoGwTirvHw6ua5/sdCD90NOz2yjFrlK4rtzWROmwqrLUe
jaPpyhICQty2lxZZqEsFvIJn/42UIwxMpx6G1JyY/vcRtsufMCSq7fzYBSSo3HTA3dwaR8OB6YPi
LoGDG94Uisob6JQDzwO9nTVSa75UhiT3CZ/+2zIsQbUneyeVLz+QWK7rts2B6jgqcC05qwmI+/6w
E4WpLii/+6gxcVaM0gcyt/p02+pkCUlBH54oQZV5blmLl0l7RhvoJKFxNpb9hPGxUKvTD3iNc5V+
ypF/hduCO6O/Fcf5TRoj646BvjdVJbjugsE78DSC31O5NGxlV8a+SNgtOJgIYx3uzoZJnUT/RGax
Ax56VLgqsoEEAycp4aw0u0gExvrekCY/hYURLnB51lWcQDPMZICezqMgZSz+5NB0607l1gCRIPyp
FVDlvXV5cCC844lHIEQ8P1lPoptexDKXOs2yWHOeXuPPLZ49i0Ro7WEiG6TCvOzhQl84xMrOem7k
6V4wYnQGD4KwgbQdikzy9JpncorN8zqZGR0Zy0IgtQCOXFT62f7T7lBcNboTgnfuGt10s9a0XU3i
1p7467YGrkzNfK/zJXWaO4iqzN0S/5JcUw/ggoy63Gyt1jkhLCqQ3/0Hx2peohHzJuAlzb1VreAB
sTUj2Yj/kWx/Gr+rCyKLAs10c7DpExQBSqr/KbSa0z7tqaob3fiRgy55wslyhTPYeX/R1jj30lMi
Ald5NgfoGOTVz5qpXbO1Npj0FPajq1jXEFbOnWhoIgZqLXwd/a13YoboaSELG0xMARPQMVrddo6o
sCzd2ye5ZGmWa7j9YHBW08uu9LsvFEEUVOPOapjcWhlHAOQ2azFc2tuNhl69ztMPYVqRe8qnMse+
5PaBTKLNfp/LYkPU0/yOQg2BivYnKG5VS605oJSIWeisoi9QodXvdcWAKz72CvfPwTKeZifFu8ue
Cjcrxf76DpGoEl42nxiQAJgd8bSGw1FSu8ylwbOow5CXalBWmvhuV0JIkY30qEO1PycQV2esp/1k
/v3bx4Fe7yMDjWxW6n5NIVAWUxYCO/ZF2w6x2vPJ04IKeU21eZnxeW2WVbiuzBi8DE1aWjfWBllC
XGcKtxEoKFpY6MGhpN6UxF+hv6T09Am83BI/AmTCFsQuyM8nLgK2ijEpX+e2yr6/nCHNBbXPv/wc
1+deyiscIDf+UALDEoZ81KGCVgW6ud8GaJp5Sskj2FvrAVXYEUx+/omBh2F4um69B8lG1wibxhSc
BGLhCdDPNGdpMRPlMSvBPN0RjPne2OEfQl4fTFAO63KsQvogDv3W1hP67q2Ga7PpcvZc/vxTppG8
PslPQkzZUpuC4AXRoT+krdV9nAAV6gJIeNATRN8/YrF7eyiAX1kmBEmXBFO2gBNnjLnAsR9i2XjR
/300UH9wmuAc/lPDIkuQ/cQ/KcaynLzqayapMRMdd08mE/Oe2HUTH4fsHoojkbsqHCSvaUK7hldJ
RVrhsIsrt2AYFOtuDl+Bxhwp2oAc6ZEV9ixMN5vBbWfEU9XSnOpkyQhIakHHyZzqvzqU/cXg/nGz
Vn/lYgpMtU1CtIbaTStvMaN6qluL6IQjl/uGeZCWvUARt7wtbvCz0AeFvLIzs0kn1yzWJJvNWRGs
ZyJLZNR6Rien4uV3fceLzrZ7y27hj9rYdTUzmnI7eT7IIiqKGepiEzl4sF9DwC/8r1RVf3Feat8F
fVrGUhqsDCOVxUyYhkwojItRPn3F3k7+uPbe9EhdXbshBJkWE6KIOLjxqy51EeuYMNLJ9DJlWbka
m+2GO8StpfJ5ziJ5qhXOEKdanBF6P2wQq0XvlEYWL0ukTLchaHm6YWNK6MjE70mn7f5DITPWUBZ7
aNo6KZCysapQIgUBiyQ2vXBgSQ4zvZ/AucnQSdb3qaEZsm2KcU2b57zhHq/+bv65SsdlEW5S1st4
Rb3o0/6C3tkbRltjRl8jqTHlJLLXUqtqUMMWGqhVWpKu92cChGiulLnU+JCKX/6WMepbzjAqDUNP
4iZgIhUiuvNpEO29OfciBOFTlra/au49nWTWwscNL0Tj6IY5gUE8VIy7vK7ES4g/PXHUr97oZbaq
TBT0LPd4i7bG/2tCmdBi3OmFJgCJ7XXkkCOUKl74+aJYPe1LpNXPtnZX8mPg+ZbdVAsomr+Swlv0
EB6cdk3uTwTqz6SqY/KE6T87pDb2f5BjwSu7GqbPWvfI/R5upX3SEisNHxf6wEXASRV1f4Gauwl2
uPiBQccLn3BmNCc0M94ROvS4NBwaYB75bWVsMStrVvdaof+lE9q8gCNS7ZNTdGnk5OSGGVRxAw9s
AkIaF+ObbVAVO2Zr5CpW4HQlOf/nJSZgQdhupfJ6wNOU2s925/K2Mc0rsujbWfvbJO1Bgxw/8Kan
c2NIz1HJe4qrZDOJyrKyqPA/QwR4grPMT5sPrvLSqqPhSKevsg++VTTFl4g9Rhacg2u5ALA9hZHH
X6JoZKHxZs81osh+sZ/nLV3TslY0dj5d2iZwj7OE8yGleHyFi7/jz+DVxEnLodk9A2Q4Xuym7CUp
v8n6vtGvslUgFrO3W00bZa4WqwUwV9UgfiMuvfFNJs2WYFoBcXbU+0vrcwQ5BbM1gTSoR+1oI1Dp
ddbLeSy8dgpC7F3oKIxUnJh4RLyopeJjP8ogMyxHoNq8L2pIx7bwov7086rI+nQdLDRuusRlnXOv
rzV+cBbSmDdNVP8/8FvQEeYxge7P8pAkAwy2tl1mHher0mYT95KWlJ6eO6OUtzosMp17imEKDlv2
4Bla/2fLC9PN+aXTlI5CSgXXnAPTjEETG0D81vQpRS7Y3szS12E+frMgZ8utePnARVdNAbGqBxNU
v2D1xUZ9wGupZra3rB/IIMIpHPhHGyobsO169NUcEwRKOriRVcmRmkvXAsEvp3XPOt9vkWIwLclW
fVc7GAfesWNrZX9sU+e687OCMyBpj0zBuIVAv6JPSzP3YqwVCqrlQeMGC62FE2hHDO/XWanp/rc3
qM0xilawMrmQRpS2IrzIwfFE2SPTMBjdpog1S9hg8UWaUSYnUzUlKuLX1iKOhRYg9sTv3MI1yXDP
240++zS5zkJ24WNMiq6bycw/oSsoQEvJKuP55ap57mpnBY23LjUVSidnPqPMx2eiHcSc1R1vXPij
OQ2kP/86tgE/9gXf6y6+ZEySZyEY4l261FjdZGwupyRBnpQUlyC4Qu2y/dMMVaDyXnn+qrlWU7g0
xdvdMjzyAAo/XsAVlq/YNVr20tZGfNe9cDJ4tR8jLTpgfd49C3XuXRHoyDf0p0DdPpqBxxBbKqTB
1+X6YmXE1E2RnxdJk59SMY/acqamYjac9e8BuszG5S+ODMQcJWEWL75MaVQGP8a/kkJ1qcorYsHU
5DHczpfVwAvA7bc0aFBPyWkPsftLElAsXqrNkKy5nknWzfVXCIhBiiZB5NzTTTcwNqHO5PFx4vp0
8B4Fd+WZag8FMqBgWBcR1TrefJvY8JdA/jmQYeHyi1gYCSp6z6SZ10XXnaYgF/A0RYmVlB7zYuJX
23swX9zspKgFGNqHWg3e7Sj3KZOAaKQ4W0qKlm99SUse4W2FcULs4RHhb9zlMiC95rwdy22c3xIF
as1Gpzt9GXKd/MMVXqDtAxed2c28D1deRkPSF0iQgRSOk6WcMhORKncE9s0JBq6cxeoNuhf/K6Rs
e8fAtyVhyuGvgn7d07sWR4P1VPE7P/+O6kAdkDljbFdMTISnNH0qCY1N06crmwa5hBfLmKFeLMeB
HzFVKJOX9wXaccxRq6iwRf68lC9aixudmUHOJQeUVhAX7ezv4ehFsA7/zExJ4nf+Vc1Ty698BVQo
6JbByP2DJH+ukT5hyQD99yoqP6Li4Twvq2cm44g/gzJ4mV8ub4ytxdjEs0CE1a49ckzm2ZgBGHhR
9AcXHXcCNg3QH+YGNemMUc0rLPw1yJhu7OVo1wecEXFU1XgnEtJcjYdwWcWIe/FWfeJ2ZqTWs/a7
mUvOdd2l5F0yQPidJve52IEZB28RSqvtW7snvi7Lq7Imlm+EtLopOzXC7SvIQqBDfU9AGGJL90rt
W8O8MSx95OnVZYkBIrVnlQdNQC1P93NnZ4pu5eqOMZjh+zEU+vRQsmymrwsrJvZ6DCNVgpjE+FrO
w0kVBK1k4VYQYTrpY1vLerGb9WbCa7L2Rma7rfS/CZ5TmvIWzQevn2Jt817ib1ucWEt3SDgrnplI
b3Z5wM8UyWrOW8xc+GuEXmVuT2bHppjR+80zwBxcLcMTiEKQ1CvC729YrPPUQm0t4C1RKIcIH8WC
NQhnTWYTRGAxnOZHBHaZbpHZjZIFwlTT/2mb81d1pOmKajVirfIrzGRREunJyn5LwKlSycA7I1Et
1fv64s23q9c0Om2gMjdnB8QasW3wSInUlcw+0KbxjxuH8E9PleYiIkJH8lTCOTnPe1Ga8qiXCIRr
a4TZ6EJ0/RqqVZkZ1W+ZiF9c4LxkTBvYAswFeh9Ni3K0/dZcYog9tlUeRu95wl8+M/soCjfZYJR9
l1m/2HF3vGNrRuw2TxfXlOZxfKHWdSKyvZmrahiPBGFTAbrSI25qnfPN4hz5M398VKz00KsofKwF
M2p+caUbuL8SLvKRjH384LcUasQP+Bdts9cow0g65dNPzBwSvhd8ZPTll//jIqI0lFJFqf/kHMSq
HL5upq/3NsWsFavARJHP0wCxG2rCOfcuAAhhoQYUEyEuzru7OPfenD3sxja8ZN5Ipns2X3boA36P
Lnt/uzJUwhM3Zuzj2giqRCeFHRz4Mf4A+2wQ/b6VdRspCTUAdF1f0Kv4QKRpzIfDFj3U4rcXV5qE
IQpWITJ3LJF1EPG4k6gpSWumm8fw9jCbAKC/WZTIzAOjTbYzepX2AjbpAXGU2ymD0mJIAxA2Xvqv
c1AYIuBd0kzWTD7iGJFbMbUdx/3C3F23Xfxu0WwQBrZxXXRic/O8ohR+lzYHvCWmAwVXFd4l6lPf
AwyIde2vsNpqEDHaeD72RvRi/CQolA6PaBYKDuX1T1kcZN9YmY9Z8al1lBZBhMOloQ6NV1PIoA05
k1KM450Io3XjxAD9qE1uZHq7n9c1gsbFG72Rr4eNbbBuDcDcuZWLMTgOWA7eysZBRX+4y+RoaWZI
mcgJLiicMt0ljfqZ4Eu0qHgm0V36RPXw54yAJWaAs8aLJkXhKQ3QdIpIONx7ywESJBBQ3SsgHOwx
3c/SB39YTd9iScHPDnb6woh9yBXHbxJmKi7bhjahH0gkq8AqltgUii85zY518p8wX6dJcBmyenJU
PeD7pKV8fe/AVDjJMs92bRC7hsC1cVxSoZmOj3fmiZ0ARQIYGKxDTKjHP0F4/pjtuPt7zD/DQ/5Q
H1jstfVDFkXu0TRbr3yRiQZM6Z7fYD6qOS6YnRjNCHL5YLFcaKy6aKI8yaYWjtQ3sPVVBF3ZKdOg
sUksbiEa639Dj8TJaOXcMRTX8TNKm89QLruachs4EGjfFCtOmWk1VvNSPdo0uE3Ql+yxxtG4EumH
1jywId8OUMgoXBYfemMs/EWwdsAyXVWX1Oxa7zTRGt9K0k2XJCmKtQ5SfMWpgQnO6KLE0+IevGOs
WHdbJVJY/XCmhy/fij9xf3fulvUF7CQR+nq+bJyD8s0c5spPAYyOaePAl/CUA/+E9h7HgQc3Q/CY
/pBpsVPkcFsI3skeLh71VZz8uTb0Js944HSOj9mAyaOj9ysou616CP0Eyw7XXechj8dSenxzHq7I
jRysHHOXreBrC3yEx10tZxO59NZ3fTMj5wb7g0wEaQmYUbRcE6yzzsa1HsDgpL50S+QYXZ6nqgmX
leNfeeejMq7NVI0z1ZTJoSNq5xJi5oAdpxIDSr4jF5TC5uOfbn8yFq1c2N9JSCLVYKO5fHZwzyRj
+wcPxHlMHhsP12Aq76eA7zoz4MLPt0iVnDMoWvYIb2OYMe2IwGW3kabMJaPAGsQvU7HU/J17M6/T
WPFdsOm36/bouIb/Hd4TVN5peaD476/loUTaI5YOf3LlLGAesUKvxukbvsmh9DjoU+/31im8fkPu
SGTmvy0CTeXq7MlxA2DtbihXMx+pK5qDZOoar8eUPpYqkHRYZVYOkuGoL5h9WQ+xSdhhwkTSbOFI
3fa3p2ZypnDIw/mU/uHElANPgehdmGSzp2XeOOxBynbLBgwh1GzqQxAMW+ib4A7jaITlzi61ADPI
EoV2uAo5TKBSjKo8E2212xR/v0AYiVLbDYz6AKrOxwOiAv0lInFtRoY9hSJLToUI5fK7Z5S1XfiP
KtpdJw57J8LeiIOs3D8NkIiwoIrrsLSvIeEpnASRryJB24gbCkghij3GqqpvRGLROv/50twNmv1c
NuYpTWUJ9mFbNNByzzaLgoYzTwY5lpGtvqOAqAJFth/4p0bvB4BWoZAlkEQCfd/fcB5KVgki83CN
VBpqKxQtP58xb6y11Ob0879g8V1l/Euyq5N0T6lFvREhOmetTqSnp2EJ15fJ54k8EKDSxvQvBf/4
wy6TqY6cNhIQ0/Xl8luObZG5F6QVABs4Ex5eDP8whdMsMMrR2t71r6XEZGhw+ei9Kqt+fUbpYEpL
G5uQHxtC7hjx3Tz2dyXD9D8gqkHrVroRpm7AUs4GGOf8JPZesQsgf3Nw+lI6X/MSKAxFrk8+Y2Bw
QDXYqjJk1DBt3rK9ygkTtZiUL7RQWm8FsagxSVL1i7xYdlsC+b8sYht2Dt788DC9JnkmIp8y8GZ3
jv6YrArIlAU+8pqY3W/8y5ssoLVf/ZZdZUofnqXAI/F2/ZNoM2/Dc9GGiWhLO4jmc3AD/jqfD3JF
kE4xgqmvf5CROkQvEUphS79PfcBSDZzrAB+7ja6ePywZse2vSAkz3pQdwS/z3ifPGb7hPvtEIEV3
2JwWzDh4sw/ZKJniGGxMcKsDwDEWKGOEsWW1l+PS9OckOHpNRfBoEYc1ZRcsmxe25er9TgiBUVRe
OxxY+PkDyJHt6jxaphys9Y7bj8E91jUaqIuVJqPUtu7nN1A+Pv0aUIyaZe9H2I4aTP74IHFzYsCj
obooRo8lYWMVzEtdE1uX5ptKO2o4yL4zZsgsBS4XF+fHqceDASJR7dB8dondfCAIHZ+z/n4qdTG5
MYK480frIi8ty5HpbEb43vC6aMtCXRvr+OwMnhG5yO6joWwfrIc1X62OGeNJYyvL0bD9Swsg80qR
bQ3LmuuRmBL9iOFfODHk8Hae6N3QDK/ExjL+2visC/Lfu/jx6nRkoQyit88H9/NgBDNSV4hOgzXY
h/QHXrXrWc8CrEHyhd3Hb8kZfz6k6G+u/3PSePgatrZ2JA5eLbxJPRrbFgnjUMfydHGRecFPF7oJ
bAc2s5yygLqzbR+UnydTy3Oa571MGRKad9aBnPyXHmTcw4OPQPBT90M9RxwSLWqS3tuzj/ilgWnD
MmNWtnCUZsvEDT7cuEX6rrSUGqAkY+S5UzxBQXR3Q0wKdL4UXOn4RERHKY9s7DtFPF3EQSxIl2WF
LiPgQxiTxWCpUzgy5P5eTmMW+BlJKxzscmh7noMhMM6YhH+iOA6sb5Y8STLY9oP7BTa9AOHSvONa
LM821OpA6mIh4uC3L2ZHieaz/Y6gqw4XuSxiM6RdPYycyDScXhPplsTQRenzO3+IbwxGZ4TFF/HD
5ZNy01IVJzBeIBb167xzDcgwqMUmy2i/x8EwmrdVN5UQf8fbnfBMZjxDLvRaKKS/LQ5LLmovxFZX
PCyaXeOATlOG/bY4vg0gBE0USfQLKsw71ss+5Jg80BcYEjSNehtuatlua3GHHpkdFIUpWJMMPYdS
UPXhYI6rkFGCrGcJ8AEdHbzSyrxYM/fJwLN7YpguoTwfLkJAQ8udEkLMco/lA5nR2HbeXXJkSe6e
5PlhE9wc5fIRdJq7WkC6UyPbO3g2Fiwc5l2wVl8LSMBoIkpJD5fARXIebUe9UDCcUMzj5IhfrT20
jaTzhtNbE6qtGGw+lkdPP+htyrEteT6N79AT97D8ZENyuZGqGCuAWt57+owtOQe5rcKhVKGCL8jK
L2DX2Nei+JsHWjY3gQvuZFzuNO1Y6QytJx4aYxMS85pbfoeI5RJ/GxEHbYBoUQmxRwiBD6WKi0lY
+Y0uhH4eDayf6MBNKm8mXtd39QD/Y3/kjc5AWVF4M+k05rLbTdEljaL/IGY0KGp025MBt1sHj725
BVyFphUNq+I6iQXygNAsETO0ZRhQmzOeVAK8YgXJLe7a78t/ygtPrt1S8AS8mpRfbPSdlSRnVnZm
2MOrhD+S2v1X5W8BapoKXCb1i3hJ9dka3+SEQ7pl8/gQ1qJvrbK1Qh9dGk3Hw35WjnD6D9ryQLXS
BGhy/W2kTZWhlU22uMa/JDTDplZ2FQdaaTTIWqbXIo071qBWnJVjVe1k5UZ6SMq6DDClGnzhLnHS
vaPo8+fpvA3XI5QiWihLPk6wbcIgPTNgYF34qINQpX8oSk/lLwRiQXOXpvWvJ79h+iPHCGAu3c7h
Ou5P+55mGa8vq7EDT5cd5/mvZimffGWw3A7F4oyzUqapIZF+b+vpThRgoszXD6xymUk02L3TQLUP
SA/pgLFrcC+xZaeOxlG8Z+l0IUUcJ+w5vf0Vs+YIPUrrRS9Y3G/iAj73vxO+31uD0o3p/sGIIqWn
vHklqQWY95u4eVVR+Kk8t63H5BaivhPf+daB+1dEaRcrN0CJ0xrleQPb2ZuL/pbOd4xaYe7CQDqA
8pW3aYOed35xlFnc+payJ871W8U2gsIPI+7BzZqqDHRJZfehwuMFccC84klQN1LHbl5fHIsdL45n
Qo24BuxGtcLCwWlxeRiwB7KRxUKrJj74ujVvbcLlPBrMeMIDgWObBd4LXU55uTe+F5QxllnjQHe6
Xlsh/otUkNeYQsD71+1c1djKigWaj3RbrSG0jltLbx//PboE9BMY5xaArowzhKM9Opn1ScAp3NEL
fkhNBuBdYwkkMOMsBdTcmFywvuaNW/y4R07S9PEcxiKqI9q0RleLrbmz5VPU0eArCclSVJCCb8/x
XeFLbDnwZX6vGRnYqfOOnu3xBh6Uqob0bxFAFMc3/ekEZIrgvzR4SDGZD4RJzy6Q0QoYf59iUUbN
R42Y/v5joXiqcswLiKo5XAolzG/hZ68BvjTZvy5PUGpnxtlG4YhoBvT5ejrYusNyhLL4EcL226KD
PFhZh4PGUBbIeCkRaro3aAfMqawe7/um+h9mwSRcUtda2DojWkav7CqnBdNYHLqua4GGf/Hibqa7
Igqe5Th8dK2I+OgVK+mIFslCcGYfBDK57FRPlj7fIaEdfFkxDIr5fs0OtijIsyZT9bKd/mb4UOOP
YNrjyzyNjqbK+PxPApWLg7w2kjxQnX3eQHSD7x6uIXrnXIr3OgzV+QPdjRwRrKRGJMf4WGYPGbCf
+QHwEVpaF6xQ58BSBrvn/xUTP1jSWLfbk4lszLGoJpkEvKJ8VjB2G6xaq2XaURBnAHJONMvWmiwg
0wmdH2Ie56SW9eXNF3PLunh0sg3AqQKrcEZyEE0NlsoVEy8qfBuyTn8TqQFWK1OoSYrmNrpY5w0+
b4WAPSCwfFLnsZGn+E1I59smIDm0ZuMVvJHaDgABX1r2FRwJ9G+7dkwmYRKFgxqos4K0TCPucUOh
zXSwtvTve8V5WKkrlkdfQcvTZBQ9xalVX0ZFRM/CVyEhVBb/k95DbpiEoDRQfSqvY7hNpxQJVmvb
AZndDuVIP2115TU3mmdmyMgeFO/11qm/MbYDVqFovXsOAIK3pR0N8JGIoYvNT4xjlPa3dZHyYZGP
OCq2sxv0ukBK/xbEGrPvrhij6FCiJv9cGAdCWOWJ6GUHFTa9SgDMaYUv4swpZ8/ZFBIyowCsZUdr
Woymp1MjipqSgjotbCy73Ce3w00uG/YI+jpYzv/H5CpvIjx2QkHGNMmhn08RpFtVF2Ns82tcHird
uf4URTtW+C368vni1RCh5QGJ4SkzFOeVMNDTBaOdBmaPpVhzXu5e2Aj96AGo1P/IQ++LGq9DyIe8
bMriNO1Sa4Gcyewu1HnumKjjJd/ki6vHVzedo+/6Mw0ukJ7XNFt5ENPQawqJ6tWrzCVn0zQ3Isob
d29L9JLcZ3bfUxIr7C6cMsRwTBt0WHBloGz21374NK5E8zS1gO2QtHTlQUusEpzHSLM62ueNZqQn
z6Kz6Rc50cILPHa5TIC0RnfmCpVrkAt5dwONvRKOR8hkhs0Tmt5wFUyLMZwUV8X8Ku/OxUmIBmtM
IHkNXiA7NQ6lrgYH1LHkZ9pARMQnmes1Q3JiN0mCtNN98aYdhBAJdtYkoAXCWxmCL/2MhmxSexn+
SDRzcAQBf0nMW4RRsu7gAxoitf8cmLxCO96lyrBcRcXSuLRqShkRfZNHrbGE5UlLogf6Xpj6quVo
YigfeZ8utSQiOLFOpqtNM/O0KhaaI+JkeoixaZDoWLESyWG71rUlOzJs0dDkqDwKnPzoqrjCRb4/
E8lLCKdtyAu7XNu9PBG/fs/qw2XaBlAmNTCM7paWsvz76X2JpooaeTKKj16wCc8NQxVCpbXTs0G/
M7FOde6KO6/IVuN/mRvjurDlSop/wVK9cZRZJTpZlMIVG/6r5OUHn9qfqO//UFpkSeba4xBS7puO
YNa5VEttwxOoN8L2Qs+xMIAzbusdz+Jw9Oo/M4pplekfRrObcGz/XDJYyC1kwBREq84c+plrOWQZ
UtSY1nzQYIWybsAVsDSGaFi/oLai3lQaVAbYm4niQTJppqT7d5z2Fl0Wkswv7/t3CYTp7KYjpYW0
Jr4j8nzndCd92HgtXXYd7oLp8vPhTJD2AWBFLDy9t2r9uhMiCqo6ilLI0ltkhhk1dt4G1P85Y8fN
BsLG51rrkpRnD3Blz9idv3ih90US+61gUiXZ3TL+cXvHs/krlwm1x4uqT4I/1yAHj9Mmu2nEUaOe
AfgVdVF5+I5JA8/iq/VsxHrSvcw7GRd8mEnjI3LFYdxIdd+dcbD4TFP5UToPB3byhpWac6gbfDvW
NNj9k98FfRVnURBWa0PuiECwdbO/EWnxzxJ7V7znAWWvj1HaWccyeiUlzIhWt2AbntInieke0ISe
KUslUolIGtvmtSAlrE9xfgQbeLWtzWrEyMGK5SnXeRrlruD4BG2dypMeOa+Kf97mcrlgRmyt4JNX
3xCTJKecDvaIqXT6CzUX1okgHgbMNkjpNR7MbH0QnZ5WeKonX9mGejiQaWvhxkdV0/BM7T+6TK2R
H3UrauXimUAH/fJl0KzH1CjBKZK1U7fXl44hPsrrA4UtpWGvxZBvVBHdIW4vu5awggnIQmIDLsfp
wKZHCw6xkeSPBNAyNglLguW47q+Zg2R/BKGu6mvNHP9pmKYhwVJf3CkNwp/yY0ibP6ZuV8Zw+poQ
/YhamjK5lVagaifGo1RX9rhnG32/IG0QbkOEY1HoV29fwrvit1NUdFMU5JxOrtNCSJOUC0VY2mzv
I+PGKlf8+n81TbxFKTDhkqjFKVphNxDXzA55DObb08WErba9bH38wwYOcxZHVTvxhM/P5ZQqM+0l
Gkv8m0zmLQqjVMOVI0Q+IBPl7w5TD7KAAc20q85NhChVcnT6T8wHXrrBe1xQVuLi6ZyoB56KBhXg
oks1nHWeRPyXihq9Tc2P4X8ikBMKhsOLuXnKUTawWQpoimJrSyORugNXDfDAFiqn4lLdweFFMNgU
eqrhcA9mzpnyo11sh/kSwvXsOERshiUCtXUv2YpJ0ZbcYC1BJYwcal4wSIybO17Zo2pvoEdK7huX
Pqt/IBinvOa807+XYzYc4KBwZqtjdSid8G7v1lJDPH5k/Pu2O3D+S/Koq6oYZHY2Q5c222hvV8e9
YI0gUjwXIzKA5FRUZ0dAFx8P0lxY33BYvD7LAxabZZz6jIjFyPzhCUTSQCPShdLtyjihToLcx+dP
15R94gmlWGPG7yepmlzQwT3iU2HnflXv0Gn0zTyN4V5EW1Aj8hzkfmS8uv8gawXYrlh9tAtl4FKJ
r4XD2lJkmAUZ8PUTgXw+Rj9m4Q1wAxSPgKUAWX5Sm+B2XjX2e0s31S/qnH25EfCa2eHOZVQwEJS+
UW25q8y7Q4EeqzOZQyiOhFJ5R0cFQzu4q6oRDODnhS45ED4siKHVDdwj6Av/V/g7sfd77zupSxQS
+7dpFvXzL2v7s42/y9FFrElOeNiP0AI73FgHGeV4OhtnJa/ycwF8tY8xeev44qT8REN+xXyJgCjV
heyf3MTgP+i+G02hwfZa+2YX78iaLfIuO0BHR//UoknzitenIEm64UDXsvZyS4pZv/wWylCs0QNT
7wEIOTHlCQq7ZlCaebKyTVylkA2H+Ymi0RJ7sklIHR6EodpNMxZ9hSJgA2+AlmDdO2JTjZBXM6c2
iYsaXUB8xD5NkSBdkNdy/UbIGfiGsygzt8nasPzxbTRF4dz1XeWjbah2ACA6EN5S1G4GU5ODTGV8
ScZZ/c9PivTLF6yoWtbZIwN84a02FnDy9BMuRHTNrjJlk8OFGabAScTQ2bQ1cx1OeEXTOiS63oi6
wZuTWM2uijuFn8Q/vrj3ww6jRU/+2QsIDp4T0m/of9XM/O7JLcVCFSnlnJYxFP8ADatdo9yV71No
sl1NqP8znBXoSLgddq0uCG5ds0AD52lrV3579O2UwwOOTJKW0DO6TPte62a0e//AJ8RV0lZ2IktX
fp/oIzdNsqc7fEbWm1GoQTpNgHuZQp0kPsKHpeSu9vtT+aEUKRAh4Xa9n+zAJdQTF9lOICquBi6o
JWxFIn9FF7+PCDLoav1r8yaZB0BnXu7Epo0RGDiqS4yCiADUfJzmi8BicogB09MUyoSOxKvp/8Mb
CSfuIGNHMeRcvV5dxDf8ZEewfVQi2L/PVkZynWAx6T1PS2G0SJTNOy6YNh4+wShkyl/XH6WoCv17
u9V8R6PnTzwoyeA/r8THIuVHs6AGg82oYkpzSvz722Aibe18gyYm9kZGWhv3ZXfJTWBFoc55x1y6
SU+ufczQphxGTk9Cid9WfmK85IsFhczgdUYzOdpL8GnXZmllf+xTjZPxi7LuOqZiDN2v67Tn9wY3
X+C/iaIdhq3CrvlpEjICHL5gbIFoy4J57EBojbLZjrcThndfvJ58p+mWs5P4dPwIVPkhc6wKbil1
/Oq2QMLSt7DJVy/4qes4kUt0KjN6WfT+Cll0LlNoH6x4LH5XwKL42gPrD5OZOmVfItcCIiz9ivNl
pwBfc3qm3VhlxvmlmGlYBQDVHVAzq9NnqP0kFkdei/R5PoHSdVTEakWjgxqsng45KPkE0SEpvTW3
16XiA0MeVwMzNpigCP8OCGAabBrU6Q26hPG9THHG7K9XF+/FHrXgt+687uXucTHyDNztf/0+KbFp
buIPnrOG4eFIr1lSUxGcC/0+kacyuf0R0dmjco833lwCge4w/ROr9F1+OPoFKaVOUa+JMywY0wZI
i9hxYOnUe/Lgco9tQPvhZCEfm4r2ITYGuUPVhpxeXIcu22uAm4FlAUw1+n7jBN/i7EXBt05viFFA
JSImgYlJYfgZUFaE5lYJfQsOEhXD6G9m86fr27uQRhG9SfiY5WwqWN7G9Nji/R0xxBo29riEbzkq
HH/pb6mqyRYbVd8Q74SQnYqRK5lMa130Q4XOsPRA+U8Hy8+odWnDb0T0Fsul6ti42XbcEg7S7VF+
vry48hvEaL9DiLq7dGCvPRYPZ9v3a/LjJL5WYG9ySPc/UgeXv9HMbC77e6hqugbaNfLOYHyW3Jl1
6jn4OBl3y9ZPlQGDxq4KumFU/izHqLkVR11bM5bJ3eQO/gpdroOmpYivenSCYnR2XdBRUhz7SqTT
mzibTQzNKJgACOoKuZmypRrZwHbpm3GHU+kWnpLv10Cj0yW449tPfgVWe0iYmhqUyN/WXdg1fRZx
BoLsnogOrxiRm567Zktbmzn0rtBEW1aN75jYbGmlqBuahsdLI8F5XYtiJE3uNmeKRZylZkyZLZcS
hG9lzWANoyNYSPL0vqEFZRlR93yf1MoPVlmYFFTwFvl5EvJp71dQcUfWs+5NnQJrxtC0QR0C2udh
BzZ9IozW+8kL/WWOvUcwfrsnWWorWk7TM+FT7HD5i6v2FxMCwX+oarmT8S4IswVdiO1mCpEnDR1U
wTrM4oF+3Mikh7YrDh4/lXI2ufQmVANK9FpRCztIM7BwY5FPxxOtzFqLVQLsulEffp1ZY0dRVevZ
oRreoTf+/dt2AOuHnC0iqwdyYGIs996QgvLseLxtmzb9GUckoNX/ut3VzZosFh2BLcVWTF00ts5o
8TgKs67ilTnwyv8qtXiUBE2N34a/sEdR6bOWDO57GcPMK4G9w8N9D5yihknYuFSX/dmu4XItfPjE
/BxG45+e50shZa+eZHAO9e99igbzo0vCyVgzLvSt2nBPKLEC5AXCAXOiw8+L/CU11XBd6YBykPAJ
XCb3SWi8VVO2NTJdsIrvJOLHsocco+FJD4sB0I82ZSzHrFHAIITjIFonlEse56SM2+VNaipv5dyx
LvpcgSvyYkVF9D+6munSTPaRdTtD972XcScLXXXMOyeJohfkgu9q6ir8mawSNPLQN915+fYbvgy3
dbJ9MpR1zD8KUxkscU0yxMoAJEo9gciCb/VGeRM+Lold5crSAcNv05/oeCifUXCWLTpmDSrKfj7N
mSvYpa3KohulEOqX3P1wzkasWkNBVjzVPWGVsW94MMMdGovxKBx8Vi9CbySLJ09qozc8ZpWHZCdY
zqoU/rM1/VhDDuJzTdeVkRNVTzoJN9J95lrwE+fuow1+T0zGQ55o8keBuZXjxvaz8n9BArmgws7A
B0kRKPfMdcg3G42BjoXCJKNsE3PGZScfrvVKgGiRftqh1eDuomMkZS38qUEeOSDG1sbQi7B2pHGA
I8UzTL1G1zn6M65LfiuQQOIpc1Ez1e6ub0nSPqAHOX8iOi18oLOGFsbMCqTtezqut0QCIbebwCdv
b5Q2CmWqjXEUSzPvRgX6OXOB0zRu1GTAzPlO7q9nv8sHZjwtOibdjbHAh3Iu03297/rWbmxHa5ww
qHBrMcmtFKF/c1965eTn6c1zaju2vHeSUMr1dHG6lyY3QCZiJEsQgrjoC+HkyZ3XHA0wwKMbnexh
ZdUVAaxayMqoA/dsjiKWs1Y1XoSUL9PrhxuTIkyoVq+hc2SHINk/6p6AWq2GM+1sfsmznZK8Y1iZ
DGClo4nTf3u+5+oehKJ0Oo5M0yedvMszlfULI/uW2gk8EasFlAqtDwj9XQjIbprB+Ua4JFiaRx3j
ckk/oWIDfUS4ggBNHV0nctbGoVCbaTxZFPReT7Jc2ZVvHH/muXRMMEhkFNhDySXxEXnjFS/zqIAq
bZLJVNGXL8AQ7BMRLopQatJgHVT+j/RxKlhU4rrkxXsS2fvsFDxVfKdQSfbDzcmOhzpJSBkHPeen
uiTXPbORPdY++zvNRo+GLvc0OdN7QyKXX0L/OAlsPqiTqElJJzIt7Qm+8ndgMhFeONKETBfc3AAc
otvpdkVe7fplnGW7OKeFPzu/AM78Gy1vannIYF4ruolTD8VCj0I29CH/xGoDb4r/BrcqoFxfWs5A
2pjAhPDFyMXZ1XC6X2uSSDxhAYO0xL9wXYiFh+b4weezZUxnyjrW0ECMJTXoceqKYYlPqY/tAfD1
s1t5aHrl8MkHXTVqPOPaVNmbVPnBFgy6UAqVE4epf3Ts4sE4/9BhEQKm8a1FmH8z9s+IQWyCfemz
WAsI4FBU3n8Dx4fy4kLam3SQD08NB+VhChoAWWKGf/EDgmR4qzK2iYpCqwfKB65YkHC96NA66TLi
V3q2rhrJGz46EmQB2WGjUXvlhMP1jjPv012DmLG9agYEEGmWiaK+4MKRwCJSsSfTykkyEF/NzeRx
RaYGljOao1HIm4eLQYqY0DEmMsDNqr3noApWlaOVCdyRTwkF86vusx74JFS2PbGI+ta4HQNDdNb5
coAHrAyZsXPHFxzAjwgsLCkD2PXZNH1UINAZiji8uIUsAiWxLQoPyvbFQQy2e+2TE68R369G6v8R
jC+JcVeiBsJRAykXq4aeegUi4BoHP9/eZpOlH6yGsC12uKBbfXKzwbOCjzUoWyUPj1yyrHws4LNs
pBGa3mj0zauEAi/RLYfovCcwGLVr3zdD7DqdK0El8Uiu3ZHiHKIzpiRJza+fBEKT46hWfMQoLVE7
wjee8ttFjBLpP4OGz8LBGhNqugDzuZn1NTl6tfF9A/ZObYE8C7hAjTG1DtWdtVBaIk+TRwww5tNK
iKqLwx6XLUH3MvKV8lSCvDZajpuobDzjruHH3iBKjGn5tbO2o38Yob2UmiK13nVgbF59izJzuyml
aiRHH3s98kKDk28RBwTA5ih+t61lZV5+iRZnmpdcJogXDJGNsCuB0JzXMDsJ364uGWXr4D17uh7A
oPe9qzUQTS1FiMnyF6Nzw6s1GH5+BfiNDkaHsltSoXhxCsyzYW7r5TaC1FrMTXAELJYokiQuGCMM
zvtMY/OR4z5lvyartnYLS4WWEyVPjtRrMlwHDtU7EfPvEiB1RPMxK/bAeD0YyA6dew8r8puNie1m
cBQPdPeOf897LGk/5/+EYDibwa5sZlT9oPr7B0/WGk93gFU10AZ/qzY9TG0rWKjqhs8DCKFS5HrX
NePJCitdfhgoGb8UzHS888Y7fzNfvdE88bj/xgYjnwS38d6mfPX1Z2zC0Y1/Siz+3vJSY4HJuRcq
S776lzT8Yg2mpUWtR7fCCpcNyR/iJJQ7l5c+W6U0ULMMlRhBzSpE7DuUNBXCL1lA5gDud00tqFlX
VMPR2fhZZCtTiZpF5TGryvWX0i3dwey/8cRZC1aKi9AExukN8itGZtRuprU5VHuyuytx5aTnnkVu
FDfPK9mzJlEP0zWva2HDqowLXbZbO4SCPUXMezT8TJytZKMDK3SyPlLsWKwCLbq92N36PnKflXlp
gf/krJPSn9xcs38xRWi+HpkFUxI9GfNZTyuUFOC0zhf4oouZ48vNau8CW8SqO7ubwPGt004RWmow
ZpRghVn14nYXE735ONFoDJ03QrqIi98sb7EBCef12AmKKmcuo3mrVmcSYo0ayLA5deeoAjNr53n4
U2MGCVHfOM/Hk0hnh6nwdBNXrrawDbSJknH9fYju3CjoFD/FzTDeI1+a0Wf4QakpyqhtYAAgbFze
OGWu/vx8Dw44O2GUjWrG4Ovq6sXePEzuMBxNdj4oHvvSqUtrcU1FVX0y/XOSXyTAzI68nk2dvVkt
zHe1ZemcbupQPKhzpsdXNNI2P3sxuLjM+Xlxa6f5fYlTPyafNz7LeDW15xq4sDNP+Ij+KifSPIGj
5ltAqH64TTCj36G2TlKsFahIrlQ69QNPmsjChoaQ/wTkwDXPfKxtRG2EX7ZaRdYlDol3Bc4FgnUC
IgPb9Z/wEoHkyBWUnqbN4XZR/mmA/ydm2fog3YzoZ6SV8r1YSlLWCajqqL1OQwnOaU9YOYzGk4b0
2BlQAFAFrNVBOA6GehYc/1s1iEaMCEBuap+G0efbrpYmY18u4r4JAoaKqYZmn7lSmbhjHc9iOnBw
1Z1on9GkIL8gYB0JTnJkF/2IwKLEb6wuT8AzJlzPGyv5BY0rloZ43oCN5kpxBHf61xS3NK0gc0nS
K4gY8mnob99ys4phoAWMu7aNd/BMPnvfN9MHnDvbcclTNZ+SYXLG/ZAs8McQZvgO+QUhiFAcMn8B
Guksa8fbB449hfXV31CDlFMxCGOyJn8uOXQENtKqTcEtk1pq7N/Q97AKJP/8uQ+enZt84B+93K5o
+y80HetBkDlccalAH+x1/mSCJdJ7A7yuT/6K9o8RKc3MSz1eYveHrgJshWjIbeZH9BLzSgFpg7tv
jmNJSgY/j4tD6NBcXfQ4mf9oIJ0Aer4Fe41DUVfGfJ0ZlStDiexCCDfHcrArPxWkC2/KfVyOvuug
Zg0PvX27qDz3HRMvRarBYz0jfdnlbLR1YZTziSHyBj9SNRClwT3leMQTaXbfDvmdYflnTHxp4xP7
dtiLcJCUmtF4hMgj+fUOAkmE4dsvnj9lTxu0YKdqR8cuHbhAglITwBP3pAUwuJvVL/LeYkoUF5cy
sVAxdKg1A+w4n3j/gFevW+0NuDkyYUM2sOsn3HFDzzWlTGgFaHvbIZIg9whTWXXQdzY5VAwJT6hl
7OFVPEWrGAJiSHP5c4VouzxrU9hRfvRes9UCjj7l2HvixfPMr60/JHUrhT8ARYDGZyRa+lpywYKg
V4igrtLJ3EB0jUq/YNyPohU4mlOQ2syuwDFNfIePHuSKwoA51txjpNy4W4UznhA4UIZ5msCTLnGo
h6pJq9mhgjgbmApP5ZARbz+ED4PgqYsw6kteqDhaIabKVwPl8PSLArRkYD1gZWaoPHzuhDjytOgW
uMh1prbQ9pgOYhVhXbn4GRFbEZnPR4bkt5dc3OyJiNxaxVck1gVvQvrhVlShzzVNScIk8P30pNpy
UCnWaagWUMpIU55p0bLyw+hJ2NnX81NQe1gTUG3yvg0srOf1KqrOsUs/7ac+fj1ejKf893qZ2nig
HlrTdPSXVbsMBFOY5ju2va0thVfO8JUASyET7rtqDnBZT7oa9QVGefXAXuTTFyI/RI/TWNWRNSv2
YaJ2sq9bsEB42E3wYugsVj+3AfmpjnDnR4Q6anvGawSkHL0tE83NwuQFgQIMKwv/+6Z+OppXjdyh
g6er0UyqimNCVSc18UjO+20rcOBRWNBMWtrI9WrudCVjLppURb/BBzUI5CK4ahwOncca0LOX1bJR
eUzSzERhfQYxjWd8r1VDwkRLveDZfxH9G27I/ljA7K8lr3dv8+mVTfsmD4jfpFwnw9m1IRBKeq5y
UlLfRC1MhodZg4pMkhnwj8ckbFlYnmL9Fot6HXf0R2pc/NCrSnGTSN6xNYbEzJzuVCmIkgv67cHt
yCd4BbxejBi/oAm4HdzWcP8pH5KIinQqyEOhn/5Lsn8Kh/yvQ9PXkRoMd3f+IlzYE8+c9TqdNc70
54xAPIH44Ls3l5FhahbbSWGuHHMKZqqpiiWsmVRZrlnSzgi05gyMHY0WyC+3hD//6Ge/2Mz7/M8a
ywyX7x8p6tGYtLik9xhQ60OW3aIs+FBW9QLn+tJWcx5MfIH3N3XPe4+JGsz66XSJ52rtHUFUAS/6
cYtYx/6oCn96B2z28xoU09Y0DnrVLasia5nHxQ4cq9cc6ocmBka4UevsXtWlidiB/ruDuoyPkVJI
XGn+vKEv/QOtyfD2JnmvuRrnBhFT+n1EBdRI+8TxAaWWRqyNNnEqxV8zYk2YLJSrT4LO2ygPjD7W
YkZLC5CIJJN4rCTfZvNl6CkZdqdX7hZH3mcXeG5vqwrLl0RiLaNTWsYWgaFymHPHWRAoxNJsukTC
CJd6GfL6zUtgeb9gEHRjIhBw83EuUizYeODv/t1pP2iDIlWkMhkiH/NpgaTdZ2SxI9RiwM5L1ZbU
3YprabOt1p79fTSMTUGCTqDAbe8BjZAnerQ6P4pqleeoq0YFTfzyivIE/4hudotEbOaH50EYP1TL
uwao9eYNsuhd3zv7Mqk5vCmsrWrX6fMDpVfE7bSX0QstWH0vQTV3wiK048MbWFY7k4r+80/k3Qh5
fotCG9Fgh5sWkkcpc/A1C9pJ8RmB7M0HyskFU5VU2FULyuNDlitjfi4kE8ictRjD9TjVERKlWoWU
1W5sQgbc2dCYXOnNP72cIHK/BOG1rK6JMFHPDgDHDORQcZz/4ldANQxxzpmK1onKiYCHrJhTxbm5
OGBVviw/6EPUOdlp9PytLfCvbVd81T6DUHBFH5qZnwqdiYjgd6+E1QlHN1MJmOe0de5uZPwCk15y
9qyXScqh/l6vnm0TDVZc7A1LHLjRfrlFA0+W8iKrazZZbtQ/1AO+wT/6qq2vFT4jK+Go+Ypp9ETO
RzLs8lHUZwpptHmpdlSl9qnz2OzrQyeHg7IZOmvud7AAU/oUF9Dh1ipdBCw2QW1TuRDbYX5jR163
lQxiqtzTULde2xqDKyfBTUCLRJmkS4izTJMoK9qvZJutwb1ZaWOgTdtZduE8IBN6iAqHP6rdlemJ
w85VzfWsKVbgFKw8SCHdtUYHVJIgddi4dbm83z0HIGRODfbLKWz+cGZb2+779QGQA/7jHxBbmgps
kGY0L+bBEWuQPoONwQvj0OljcpbzMKuqt3GMXmAzeswk79V4lO8Bysrm9yo2S2sp3s70XE0I8qLD
mQFmwYNjbK3dJZ1s2W0YJQEliNVg4K7UNmOywsJtdQK5CBXU3eZSP05NxykccVdt4PAi5tPsABlV
bQLv1AuFQazMScIFgT4Md/RWGNudaHJUp3vI7wzWhHlAqauiZg6Quy7AHxa6dJym7/MVCeZyJNLu
G/mk2Ykbmg8kY96CVaYBsmIxTc2owcrmY45kavlVrcoI8clapBK0TyjSRzNJusmvd7QcV5RJrGr9
GhXJ+syZwpSRp0EyaENfLD935BXga9lEAXgD1lLW6lGPSIg+AtGE4prsxVw5Ui6/NNo/29fq8xra
UJ8Eltoyj06KiQDcoy+9rDC5KNSaVkOF5noYKNeotT6hy5IfeBZ40oo9mF1nONfSYvQorbSGWJRU
D2dOTkMJfANQNhuEHgPt3uEOFf3r0eXSiUFXnhuNwIfPYENp6LWZxHx2ugp443SL9gQgr6iirD/e
VFSYC/HYVpX0XpYSYuC76cxhNs9degWwF5HdciZtJxShkI7iCfHLubSdQf9PnDM1wC+SqICm2epk
7nMGnkRewk5ZBpqCLJg4oQ+yTjQAau42WFBKfKouaTLLqvD3PNs+Cap4wPy2gB8E0PXR+RP6Vq9a
PzYI+W0OysdUoWyeSbTmFR/NckLhc92D7e5I9Cv4MxQxJH1jOxQVXhqwOrPcMQ9Ys3tdddug6uIJ
Q93deB1sGopUyQ3jCVgJOa5vWj2EK15HeMmjRtDMRb7HJ8Q+PAK6y10dAhSq9xsDsO6iy5lRZEVE
33LJXBLEaYEZ08Wzbhd2ZzhG7EK+z0e4JK2YSJfQD/qF4v1R0CEsiQwMsELzF1nMMC1WazCNXC5u
xL3+snMKoPN6EUQVvp1lIMoctIDtfJXvhjK4XERVeSL8W5DCVyxfWZItwQTT04JHMHmr4xW3bjpg
wxUXSQbMGlhmX6AsP22y1/BNwZqpUXyYNRF/rDfJHwgrQU4P6aRU5vZzFcyP+UcWTSjM9UVIrMiv
BeSHX6SaJVxzkE3jFdgZWI7uA338FZ3ZMjPO3ekzi1HRepX0lv7tf1lGEX+BZOcJmsQqDsv+pC8D
VGCCnYbEgDBCoqxs4HI85TwEdnMl9EegbNgIG0amKyBjOZbIYRClMRzCnOoJwRPRxo09IrSPHjzo
8JKl/Y/VVr66jvLZcMEfbeNWIkRR0v1GEBKcJLcHGv/LbWkC2vKge5k2gShFlQp0nhbu/qATHCxU
ND8dPJJlOccjDbr4mX/9E3NqfZ+1m/xGCQVIBKKpmjtxU3OK6+AehW3yEt8TAZQboDed3wn1x+EI
kT0RcCL/csIbftVYbfE+8qkiUjQS6azr6nK6P+dBHbPQcqK3SlwwYTJ+z3du/Go5Ox/PmOAmDvpt
DrmW2dCHcGWCrKMivZtmsPQPxY57J8ihdRzgcCGcP5zjOxmlR8jjo/5iOBX9HW5ywGZzWNF8XQrY
4k5ObHmAtFtm0J0n/J0x1WzqY9+P7N7yYNwQxPNlwnGlKZCJUqY8JeEi7wCCznqnAclXir0w3e8g
m/ZnEJ9AV9oU6KYOwZJYGtQY29tEEz7lulTDSbEE3ylTi1tIbGgMi9Qc2xcZ002ZzSzIc+o6gxk+
pafHIdib2sDNlUVzrWBXBjtiryD/ZtACgr10JuvPpsySCWzULckJj6jWDl3knOfEyqmSgKB1pkkl
tdAKtSgVBxro0VgaSDpV6frYQf9gi3WWEGpUXNUVYgUwNvfrxSvezk/SalELn0yUbhOr1+etHvaZ
ZHPi/VLyQEnUNbvsjoMsA0wD1Iwwz4h12aI1TdytqnR+iznK7kcVDZyCD51/nTmySFdwdzkrr/eW
6YINjEH8jT4gBhClYnmsJiIrQgZSrquKJPOW3ngrIlYXw4lfaObEbqkmELQRewI738XGUFhnS0dE
fp/JKlpkcJsReUsA0qBkr+FroqZ+VvgDqwFIbwrgid1snSo+XgyVi8xExNbDbepmkugSE1bmjqiI
mfMLQ8ReKXbwiDXLypxza0K/d5wOpXZqmRjp//BmP9zqR0iHaBeSpUZ88Z8q+o+V99thpib7mslG
Qxdqk+kZMe8brx/86iuiUMErPR4jJCDxT147d/rQL4iHCCe0g7Huh8Ouyt3uu2k3y55TiR4n20yU
bVr6/H1n1acrOjWfQcaPvGznhYbPfX30tO94vO5sln8UD/EZGinC+U2Kn+AaHHWqPeYawft2W6pR
MtPeQfaXvz6lGrc2He80JBa5xui0nwNLSx/aRiKzND5yd1NaU2W0hzaK2GU/JUPhQjNowrTEoB+s
0At59zrOP5pk6szm+8X5t3PmsFlvCxAMKRAtaku+TLhw6M8W7cZ/1dDqKVJEo9Qc2M0j8Tg5tOHL
KCvLGeaBoTJr26cMSmtFPspEvkkzKuQ2ASYjP79D8sGBwZzWtvlplecb4/p+iW76GT9qObb/ROff
14sKHg2pXrj9bEXpXDZZ2f/v77nECXPoHLZZ8/Nh7fZ4XxwgeaWiOciH1bmvQFPTmnDrTUTf6TKB
fTai3jCdvvqt6Cu+9tLgiKEPDAfpS3oplfuXha98jbIekd3on5QA/suxWkaYcagR5A+8CanRqaEq
vIcDtPQRAKPyEWOStrcyxKgQbCst7CoceFXm8TEtMqk8Gv+qnnf7X3FrLKei/MzqbfQW1HfLRs8f
0ZKv1euLt0Dj88eLkukqnD7xnFxkhRoFc15cx7J4MFenx8eZo4b7DTHw7bk6Uepw96+YHMYuAcBn
vp02R2PiSqrScHajiGrpSZJuAOJMadI5mu7CVxa7NPOxI+THrBem7aXQmjlC6y/pJaVrE+xI77Ko
k7LYxhRHCoUYrpD732O0OW4G44Ldb83h+/jKow/uZONLhO9/SkLyBttMB6o7Okq1yr8OZV9UBBX4
nZU3NB13fa+J1MayntjXItc23jlJFU+AfZMQ8y3PQIV+E72gu4CVnAIuvo1VL1YmU3/QyDZwYx1x
O4zFBzJBObKE9RWPU3ePd0cX2sgoErDA/qg7dHlk0C/vZP5GagM/GIn34iu/U5qwXUNyEcqMtllb
kuxXXrRVaiuZQJcu7VVbriAqr3YEZXq6jk+ieXNNHRl5l+MXEIHJf6T8rejeRM96jLrka9jWjKHd
eZ5ydk7bDtFYC9NoJ1k5Zw5cfZ3JHM/fDoqpikdQy3hcYAfP0NG9P5MheN19HFhp916bk+L2vXLi
G03giSLtZ5Itgpgmz60Sn1eeWybOIz+aCwcxHS6wZgQ2jXbqancr6pLbg8aUAp87x+FypRO2eIO+
1J2fPKMd/P3SRstNjgg9l0fZBRRIV6MsJaQTTlqGptjAn7ygsLhj30CawLgf4xktgWkpe6Mh9w+o
ttz1hYmntvdzc7EX6RK815Zmowje3tMNovb3wJSjQ+gxz7TsrUL6Qo56/zs7LZNF8XHqjGMXYhqP
wjYsJt2ed/Fp6wbohc0D4XubCv7bq1DJCEE2WQO+jR1R1uYxQ5xQ6TjMoYCnivMGI2ZfjRdfIcmU
R55pehmQnQe88JiYhijq1D1a6K4qvERBzrEpis1ChvEIzOvd+Jo7QWKewy9uuaPiFhB4DQsRkg7N
Wfn62agViSs+Ds6WYpKjpSArzEQHiqr2SpeLg0O+t28pxYEtoBmbkHI3pjeLk7AX4iRInxLOX5LK
1aVqR83mBjNjOVZow9HUByPckKpdLiXiau47RO3zo55WwEFaCIhUDhP090unWyBM8qq32accgA7Q
TWKxF/xOZN3HUAV1OrgqnKHCFhsOQx5zATTBpnp8mwLajlvCxgLk5ISyOku3o/f3lHwCKg0FQeo4
x1eFAOO+ABmfQCDKoOiBcKtA1UJ2VWO8zNQsyn5+WR15R4I5j0+SlB0UFPkuJMVjQkGYoS78Xk+A
HOFDu8OS6WBHz4XF5BnA9/vyAMMaluBM9CsxRx/ojk3zQGjChqqI+6KLG/QsbPcNml4J9FhCXTDp
hXMr3uGiJpB4YyPwYJin+jofoXzifCb8evPz+pHqTPZmJMK5BOVLq9fzwReEc4XKGMu+bc3qb9dx
ZxzvLGkVLL3gD3Md4Gd1hsj/EZ+8hY7mrrlFWA8JPHMf1flD7FFXMCVNerUphtwACYdLusyrhw4d
3e7hm++5Iw8CzwU/2GPcKibXskvp69BMem6gePIIMwxGsOjQUiVf3CdKyy0/eSDDGsdNcPIkBN1J
QR7ea41nfqwriz/SxIvBxOU06iCMhf6LOe2NZP9hKVDJU8PSVVn+R02cAeyXr1qWnL25lParZFyV
bDoR94IkMeADfH/lI8+zRTUCGKri5gLg/SNnBefujhCm20QpcUEjNW92EUqBf9atBBnwaCDK3DDz
MGeQQ/qNOTCLMeuk7+Gu6iZuZbHGUuvKKpw0M16XnZGHDMTc2O7sHz46wDC91HhBLQ/af3mi7E/E
B26M3rzmwSJpiJnn710WjaMhGu87ta3a8bsTUv//MnM91UiTtP/qhUDMv29JKJqHd5TYJbfeWx6K
Rmh1aDMcnwmvps6ZF8SlzOgZ1dxlADTi2+KfMhDPwV/D0198qtNSw/kHdcaSKK4h2cDWMKYOCFYi
AdenC32gxHpTUdY2zh/Y88pi+Xo4vlixZH3IOHcnwZK42e3wpKGSBf2M4oIihlwF72hz44jN19G0
drCpKZHCnpBN/ZJq6xr1VFdqA/NzXdgnBhRbmo1f4K3dPzI6z/1ckHH67gdzYEEWRiE5Oom2f5f4
4smKQqdvrtbNgdqkjCMLO38dC3P9nok3dEpSHu5dWdI6PZx2gL1zSUznkqNEoqSmMS7sac4e141n
dIdrv3qjY/HKvh2bvcOclfsJYwZxIOJp8bysXhIT6bfFknFbMev7PKOgTRc2CsjeNvn7UuZzbH6f
oyBqrvP+QQ2OzoYZFkpHJKQ5JLrBYUeKxe9/xTmw0qbr+31fEZryEXdTYU9gduvaFgHFBUmq1WWO
DAuBrv18MAY5G0znMbfw0ZRD2koEPollecbzGzzZ6C2dWSoZDv3+VeFPE4qqhDucq+wrMCm3bCsH
Yz1onmeE3JarEZdW1R3JT+7+bQECZRPjt9XkdhMjKN24h5fQLQV9QmYet1NKNmmdjQebFaU1HXY5
fQadeylAr/72QqibR5daIGxYMFgkT+/JCwTn57x+ZnABKRjKs+ep5jaHjZ0NkjP353rNgUVEqJxu
T8I4EC8IJ4UoV8NzMrzOBigno+3lQs397WLOxwP9i60RwW76+q3IP2ziLe5ZrQYMV6iEK0xEvU34
rHVHvmDdZIqvfc0y6XKKYMZPRSh0N1sXANPG+WMIdYLZ8yZADxS5mgGxq2q79UsDcKovVfbfiIG2
QNX70bkLXLwiwbRb5fCSPRC/tePkzIg3IJUos8+0tsuVrWjSmvHOxnrBLkW9QmUi1/bJdGNRjcMC
7K5CK7NnQdN6ADPpeF85AZ2oMShTCEo/DxnUzyUzyeFe0xj4FRoG9bZ9+qR6di5LhJUN2qWu+gsp
gnmw9neNQTvX2VjohSsTTJpwVUBYrLGr1IMBYSxOueIanTzOsXKLC3c1AdeAy8yMFIJNNarrP1BF
VWgrVMJQIiVgVyznSedQW3imJLu6s1olZ0dcSZoyioJvdJp64bFHcj2o5G0HhySQ8BZPH7zjiqyS
3jAEeYBqkaFxu9IWw9e1dwlpyA4DjhSkxYh8sV+oxrbykAqX9avnBllIHU8MZPgGARW20eedF0LE
r+D54iorh8BCbAOvJTVuFNGxvPry9hBJL6WxHi1ShfonIz5sc1fOP3xc4kO7gSVPyG7G7BtKi8qV
HGJ66p7SJ0XN6zU+GafSswziJpPUISPmvEjTzhNCzqZHpWpjvwIqIG/py7SNVay0kkhfwONWSNd6
Yy30tzs9RkroLN0RRXeURToqtfDTo4JlCJTibRJsGn5EdKvpRe2oZZAuJwo9Ybes+UHuSadUJop7
0V5MqTN4v6F5ZZFtLFkfmf4Wrsv+bo+PXnU4sf6xAzDu7mxT6VgspJTvxdIjsHLMr+s8qKTI5C7t
rwvFEl1O++XE1Zygs4z9nxvJ/oNCFLJmnOGvdrOzTPjE7E8xZnrqOr9Rymgliak9Nc//yj4LPGeH
I382mixrzFxSZ3vr1gEDsagXO0auzLVk+GLJrHb6+4Pth/MTBp9XQXYIu/kbWqtioWu5/hUWDFfz
7x0/WtpPBrKF3pvOs5desbz28rjnJjODpT5lehnXDrJnTr01vrHmnd/q3WF/83+1dci0bUJEW7Qh
AWsKKaAkAzXZA+pdnIS6BdXxpPYhx/a+kfiFHI/UbuOdL/6/8t48cIJQobF8sTgGg1JcLVZs/LbG
06fXXENFvfjWARPUkVMWopJuYkDFeiHUUJrj5Snc3571jy5535vSHq+FmL0IQJF4ROZr5WtPPCkc
9CBnuM8SdtCOLyWKGgsLLhNoLWkQcYOnihhPEsorKzGW+fgOTXwjiNpw7IMF8wpT4/d6e4cYdM8c
hWbYYD6FMs19Uf8pKkE1TL1EYooE3E087bo+/GNqeH/VJY7ruIjvpneb+GXTNEkhvC0DnI9q4ngC
6ssGKs92MEMr3nSoeSAfdubOQUzkpDhz/g+279rS6P/qzGZFGwsvfU4/9Wqw7KLmpBOamHOfOGAy
oz5KdC4ob/Ww0P714d3mu1m9KKYKMdPnViHdQspRfa4TdLMwhtKVZ8q08UYcFEvCHNcQFtaTdy0f
RGcCivOOvgBI2xbr/oj+MIiJ+0j1kwm916B5KsgOCaEH3aB3ppTgexnm8Zg//etXNHjRntdElGDW
muP8Xx4QMRSMR7tqXYtpvQ15NStVhJLS/zTLus/TSKCGobwwqAQ4JKry/OcJ2SUiikomMT4gnwYT
PKAnzYH/owiNM17vDistvbgPg6bFqJcDI7jYwnrqd0Uv3NESbPdW1+5IMqczxJ7x0/NpP3HBmI+n
O1VB7fHUZzkvUwy15Q08858syjryDtRfqPZbgeTg8q0YN8hIC+9FX2gV9/eIE4GFmfvWbq22btev
hkaiJwFp1epnIYXtagJXYqDZA9YetK9g67warJogWX2G6VL++u0nY9tbX98zIj/quahrAQpWxzFu
TM8REY8Q8NgiNB2K8hcYANAGPldm8+9LAtBL7TPUnivy3qNsQ3JuCyqeOKFtXOcBfr30U0vQEFPv
orKUPBN7hpZ42oS8olV7RYT8qaABaF+/BwsPycfBMt61/0fKMTXy+7H7/SRIcG2o+lsvcVVkiK+Q
D9VOBOxAiiV5tnpcyAdPNxjmNJggFyOFHZtjumvGUYkeV85fWt3AdmkpyknkgGkB8e2hNOSGxtZI
9fVBxqZG9u1q+XjKbM8J5ZnlRhWmcp+qOecxCG8sxLRjbPknoeBDoiI1d0xfgxxs3p3YA8liQ0KR
BU3KOpehKviuv3gRDq9H6rdJtfF/svpGOnHvkvbKgn3O9a/vw2jFjOykRRsVlOTbQ2+qchxfq+Vl
X8DHEjXcx/WTIarGZ80/bGuDkAJ5h/Er2RGSCOXa8pxYsB8NuTCoIyb1OYAI/VFmyboV4JLnYGaB
HzGigy6V8Q/MLc/x4gh9m+uqOVzDd9s27FTJNUnm8nwMJbATAsBlodQCRVms3Ui602jeBYHI7uYH
elWA2ALk9hkzvmR1BcXUWqP/r3tnsiVZvIvT4YMKqKxzwqE/cEqCEPmT9E+nCms3fAd/RxMCOz9s
kJl+6xMWV5BRVSBUDWS2C6SjMW90YcVmZ+uvmzAbaqGeuiQjm7MdR2TMnsBLCMtd5XmvdVIjWLJK
Zk8O6wYMLb+DLAevACfQqdKrIveXEnIdN7GYAHyd2qX2NyoWCu5nVgi+Duv81gbBwHhe7REGc8wb
JVQWPIrH7jwsaisetysjzv1tc2BRQSnZ9yl4V1fPvpcYM3DEFy/oRy8tZKIvFL7kw5zrhL7YyW8E
/oSFUyfTu7o0/XpvyOScy0hBLfPibvFGUjWohPzOIWonSDqqyN9BpbpUHb94kKvndwdpCLzcid/x
Emk62J+nQx21oymg5HbqsbS1o/Lcy5iLJn0c3imzcOcF5UZb4XtwHrYRXFfyE+QqSJGFW8wJV3l7
nojvSoMplGIOUTF/bUCKA3+k1Di91glOBcpSftKzrh92MBUotyO8HdaDLbmxX+GuRXhQqb8BCc0d
wOZfWLOOXd2js5qhLbekzilYPZULoJzwwph+VaxgEOiOt5wWs8uDYICa/BrLp+pXB9VQ6XRJpIUM
KZxZpyBEMT1NF3oFKLWOyvix6VKYieKJpFmTGzJwqPrjWkIFEBlqu5LXFgGrDLghB53G8a4R7X+A
Vobv2Y7Nzn889yfCc8uXToUrNRa7JQkWIB4RdaYsW5ddaKM5gUzLOBTUP0E3wIq8soT+pkf6Tjjp
G4+z3Ls1qB5SZL778Trk+8PAkxlSgf5ZrYe0/ap0dOzcNJkaiQK9BMRT4hoQuc7CgTMoFyzHiGlI
KVH9T98MSL6ZV8gKMkZcKmmq7uN8Vap5fMwNoQlBr+hfR6Qe9CU6svyIVKf9ZAKcIOpm6+Tr7CaV
Kh6r/YCEAqZ4CVQF9sQV3FTDQi/YsdGnVXJGL43L1zHtNZIN8/ooLb0cM746oHjcJcjgMEfCJfvR
bWsnwAk6dtakT0oU85ZhA8wYebNFBggwba8rkaN8ehDtufx47wedS+pzOvZBld6EqE+phjSXwKSY
rKiv9+j6RZjnUAhItEKsDeUMKCtG0DKPMEINCqk/+pOaJJtk0c/NNoQz/o4hcdmMpbWHOVAyttIm
Nq1WYRF0JyLq0CvZaHU14vFm/6b5uqU+XFUa/b4zJuH14ZoYirYdwuGymT3YJtq4RagrSzkOdgFa
EpdrSW9RXAyvl06ckj8Ber65+X1x7q9ZtC9ThmeANAMrtAkuXsqoObCtcaScIdONDg266VuSWwth
whrg+MyEdlhqWa5f+QAiPV3Ypwo8aycvfeoqq0eTCirQAUFgPx8Nd8HZRll68UjKdOdFMjdMSygE
ePOH7rz7/BN+OWFuuLThoaK8qxVvCgET/UYune6Lk7XquD6AKH4pvmCWQ8z12xPrRkioIxj+OIqd
aaOfc+s2Apk212CZ+GqMgBfnLP1RaReMPjY6W7l7OOnMUlmum4+9359Pz06tiQfkLXyPtiC1qYCM
zZqYy2flQHK2Ipr17JdYqY98mFN+h1usbbWnlAhLVJn0HvkuDdVH71kNqAl0po89CuTWVrleyUAA
SoNLhC6TbGskubcyTHC9bjyHy+zA2OYAPdRWfOdEIrHRjS1QsQbdn82weVr6noCpXOLSWky+4Qx4
0YszptJT4+9l/p4wzul4TnneTBVvAaklTceJ8t0L4hv0nJi2gYicSAwAaPfiA8ZUHqyB9YzjxYoC
woasRNvze13tQJC+FAvV1Oo1yx09zIU/v//lVWjHJ+14dwMS0ScmI+I8uqomXnsyRn2biGDqYVLW
mrUemYHbNtYiY4bM8eLhVLRKDJfAToltsAHuokU6jr9BNXU1RGl6uWPiW7mh6kxk1PxIDG7DDpNL
XwnEemo7ZfCb/TMVskjkrKhg+jsSjS2xHK6UpnJws7Fa7sHbMrsW5lFi2FuqSMwMAKRbRA8tQeUg
dhtVwA0BsZNJCU2ETjjhYZuI7vs14AIFrLicuCUhLfJ5g+TFQiVInHiBFfe/Smf8FogcTEPkFunX
N+JWPn8kr2jI8cMMU4I173ok3pHb8LvIerkVcUflQm5t/4lCS9d3q+TTHdt0hHZqzv5aD1wqN+gl
D3ROVIiiK4+v8u+xS6kAoxrIATLV0xz/0wun/d0LgXTh8pZHHmsrUH1FF6LXwDcCNgNBLxRnYuSn
3Xo78mpSu9sH7XDqPhka9kBVUZZrfyfsJtXD0e/se+0NTqgt5PvdlgPFHgokE2/0xUWG+FWk/1tO
1u4EdFD9YgvkGjRvXDXdcGwIInoT0GUDgtiwZYrJMzxN7yZmfKthnw/7mkq+fBfVv4egMYxwzXk/
IiaJUtYuHouQw4yEMgSEOJweF2o4B8Fi42idBfEUU4eKkktrohePOlLPyV79hm6oMOFy9ZizXQrb
nqaoTjmnFl/quD9TkNeylVsg4xYdXRqdgoiaBrEzGGaNk8Zw7yWUQdi8Q7VeOMXAHpcLK9GoelKu
7zMKDvWRtSbuwo3Q6zo6HI7Az/BYvcBTHXe4jHtlO4uf5E8lwtYjqCl6nSF4e+P6JHGUzvuz+UA0
50B4yQF4JC7AZz7l4XSFlhaZJYkkothmZRLWCVCusmUJfyt+Dww1xzPizBozwYbklCkPcLJ/b8ju
UqhnyOoWAa40SHgH/O7qsHkKvYKQoemFMEie6tyiqYXhlPuT1WnClp7NXF4HcggaKnLxIffYr9Zf
/vv7KIOql2taGcrjBgVGYrnXad7d3W7ib3vhsY0KwMHrhVQCoBW0obW4OV//aaKZVSK6eOlfsCtl
PSlMW+d9w7IGOh+TptzXJR5SKpHlH8J7Yqk6KxfMaE1p1q9wWLaR9dYT5GzcJaZ7uxgsez6zSwWQ
7MAwMtm9vnTjhepqz9/ZXWklobsyLuw35urqUxKnsvwguegF2+kv8d4XPhYk6F0Hl61r8tmOOCE5
vbc+NWKiWyp5usTkJ0jMJWOEAP+TC7iSHIpPuEBJzs8UC7vRxkDLRf27pZkgmrC65nTCVhbomihd
a6hK7jEhCmeQYkZBuJSH6FYqdhbXpD8blAhnDSZii0FE6vDByzZxoFCvbL7EZ9yoWcPfPyb8cwwA
qXbwPF7/5sKVTzpDDxmCuURjt7uAwwYAMDhc1oWu1tsK/VzBjBuv1mbdGWAJA0JguUrJ8sbZrU8L
oDOFPgCQ4tfcgXrM9dBkcXy4eHGd3qBKmBQ483tE3qmPq9A2JPXYnDZ9zSJz3ANsDl9bwWUsq8Mv
HigXviXbtXd+IpThPeEBQmxVvILe3TTdLvPuq822uY1N2nKE15qixY2MJsqhVm/phYCuUrPcgCqV
mrescmoZr8qs/STVkMsWatVAfuVphs0uvQoTZZaco2puxXhQU/PXdl8jUjpyc0V/lzehs9CRq1gf
ZUifV27wDET+0qYXDheBDy24+DGjw+STf02tFG/NM8WunGwQCqgYdEYe6ECBY5bQl4Um0tBDJek7
BMlx501rD7CUnzdJHV5D5+1ovyO6Nel1eYS9m5MHjLN80sKsp+FzyiiUtjwXwFAfb/U7tIIhZ1Kh
zRrBGWuyDwWF5d1TeigG65wZc5kB5Ym3EOYJEeRvDi0FmjrHgwLmV9fH0kC74C5H/CzhaUMlTp6n
5g9ZCSIOihYvppiTq04bWIdHoMtjJFclxLLL9nqtj/DeUSIOUeViHJcw9y3BiPEX/Hf8Vuh5Uizb
FkrmjTQqn3ev9EYpmv0h4is9cta5itoNfNkSGyBLmturXXfZlg/0e6mnd99CXIVLfi5Zuu4cZP5y
uNnkajwvg6gNPei+p2uK5HGn1rqifBWAGWZMOVKq7kY5jsRyIyrSVWa7tq4IohoTN8HBvoxxI2Fl
NrXdPOFqwnJE8XFmn8FZpplY3vn0hmDTM6cWElSQuJDjvB007sSlUHohHZzSXRaKxjUntkYTn/hT
HdndRqWYCMLWsLNxD8RWr+ZMuY7AV79RAoOyLW0ocOMaTukjI+WsWXB7qyVLPYMhYL1iXI6ed/RO
ddbvZSDGmL50gmu1prP59vj6h1aBxPFrnOJXKceXg+w4KOYVoGLlrtJy4xijmMZDNcROta7YvIy+
P19xx29UR6/cObdJ0HJ3eR4+54vrSTc+hTCCV0oM1+WZv1/Kjmv9V3or1dMBg49b7ZeWz92EnJii
nRTijHSvyk/GxXnBzfucGq83m6AStNsLU/QJgwL3wGYB6dVl+qG5W8dctfMoh6jGAjVv8KtVY7ow
I6iVcPAuSwKa+FPvo4PcZnv6Z9tldAN3m8WrtSqyfNToaHnzqzwl3IViaHhglM8Lp16iu/GSk0NF
coEs+Q8Wc1yjEqxbrLwvLgeJ7Jjt5J8mSQUfw6ag5oAEdg4w5uR/iLnUDj2HNjTSO8+tHNKxtfK5
OEv/bSxAZ37i3kLbqhLn2+1hoxg5YoHFBQgGpu4ocic/oFODNMAZZpzpYVGtnx1Q0Wnz6JH+Q6TM
TnysvP8bqhklc3hqLIkxEOUtluyAkaJK9djzGbblSCIfgPfhEOfNpn4goidKBW3pN3uE0u+nZsUz
wOGYex2kGPyrmrS1YNI+1mC2QReF1k0FhyvjPvsvd5b9FpczP8GKXDK+Aps0vjRQbqjbftDGrVzh
NhVZJa5r4SmGiXy9ah2yaLeajfyUUyYJGD+5KwMNoCUXc++6QjwcP7l/ixO3W9ry7EGt/P5Wszsq
eA8IWYDa6TquKMB5/aGHARG9Fh/2JIKW+7u8lb4hgyaHrYIaWQyYC6shTuo62f7cRtbzQwuc5nmr
h0kbTmvRUScErzzZVKh3RH9bhzbMGR+YrsurC8vv0KE2TQCVyGVXueN0dRo7tiObocmjTCfvpFcG
HAEmLw==
`protect end_protected

