

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hB1MkDF7gDUjtp9+r0pYANUYTDYvtQO1sWNXspOA3ppM8SYB929/qlOMzanhENZQcOQ3aiyEm3Wb
ozapXP+k8w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nob9JCRq6vcsk9H9VmyBE86hdNvS8BGq2p8Ka7dLN2J7EaHNc5IAaDkHipJixlCbGOjVeeUZyKme
HUzNgZTvjzVoRv6O00gQMvGJEhPJ3XxSJAOF+OM+ukp/m/tTtC3aiC1VdkFrdu6+fpapkZIb8cKo
kmCmWqIF3vlM9zcrSOg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qx+ritZx2pDvnekLOZeaFDvpDAtmg/hs096HU3U8xSeFyrj9v1CUwvI97hgO9fhp5hx7CLb4dRhp
iabDmveFs8T2afhIu9MmAO0ZqxUS0SV94sOYT5DwWoTjy8BTwRuP8Xrs/EEWKwKuWJp/Wjv7M9k+
wpkev7gSf92vj7uOWX6J6ECKwgIRjUGLc/NIrHrXqaq0yVd8j9fP6cvhVKR06OMq6U/6hMqO3Mwi
SQI1xdCXs2NXbTiCZKqVDbSBBvTJTo2cH6JXLB+E/g9NyF0e+z7oxCuyReCUVFJ21DVUfLxU3OhZ
gXG23tcqWGm/l3ZWHVqrETjEni8mwIO1yFoO4g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IXrSnaP8yioZkxR461AE2w19esRr4/fF4dA2RHFQL4fY5TpvMbkL+7RQBJ9eOLT5OFH1DsXcS+My
6KW+sTOsl2ndsfe3ttRCDI7Oeo8joeNZ8xJuwUGdOxtV0ae9PUAaVjkgDttLOomzNLph4uCXW202
bI3eFzZlGpn1iGIKiFQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iqW10+NxHcU1vbwMjaJKEOrgcrSi68eS0/IgZB3xPrIkkojO6+T2kz9ISwjr3CN6PcPo+hXCdZn3
Q3TnU/fMPFYF96Bkmhtr7AtYZE8GinVZHXJyKmm5x7dcsR8FyNv3nSOE/XYU/dyZhfnBj9H8LA1H
EJZm8T3/SQk6AB6tpXwh7kVAfE+bMsPCp98Fijzd/ynv1FX6O6GWv4CZpIVUKm7Fr8lIGCex7lCq
foNktfSIPTqF27RC3UxvVuy2VPf0Ck+rGl7pVu7l375TxqfmSlC5QxbXyTQ1NByeHr2LVJZwC+Xp
5uMCktl5vyr3uh4gEJyZSJlJ7E+uSrhstePVYg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37424)
`protect data_block
s7NslC60miDvpeLiAVueCXd1QAw9XZubItL2HDRe6VT26sYnayWcFWEmWSh+pGUCivF4Ey/ZrRDG
jvCoIX6j4MY1d+d5NOeXfvwg+kwgkL/+OXVumgUgWbImoPl6GqE4JkgG6Pk2gULnIN5iSf7SylDW
GM/57YXjF/0vDIzbJwgVWpY1rNE9xvAtA1hW1N7sTEnCLeNDV+xh8xdzeQP3+VakLAg9mu70HMC+
d0HhiA6OL1kTCqAbm4uK5T5j+G0nzRHw7Bop6pxgEmtFe8HSwgcgln6pR2REFeM6Gvh6ACq/IRSY
EWvkx0kZ/LjFfCm2ne3dLQNWkkDGbnxUxBXgv7+5lLrY1Whwg/3FrXeXZgW8zzL+a4BJ4FoOKPbg
nGGm7jl7yr+P6whsBZ++qauFoqa0Cqi/TQPqt8uQjaXwS6cpjsy+webHKCIMiDkp0zoxGaBYlJEd
rTwOO2G7bqGTVqYMDGT8lyv20NUwSYZ5RpovaNLIcbsNZPzVh9sim+8VqBHpJi1tD6deqknC3xZP
nPrSuYVsXJGvFXf9Hna02Dzu9qSaWXo0jH5W07ExsNCJcyxq8KEGf133oJrgWXufGyVFGWBD4ATv
p0yEXow7nOMCCQVFyUZKU492Dvf+tsGCF6tAiWehxOM1MHQe2Jh/7MSAyfnSsxFv8FnHK3u3ujvs
9qB7bEltQ+4U2ZjLz6YUnzdU7ffII2Gt502IPpblk+KoFx/ktv5A+JsTmW+U/fBaG6kW1QXbg/19
MBHB+2Rplchn4uy0u9x0Fy4hTUvc+qHhTH0sNbTqio2cs0XSKFswhEcaYwW/kmJGNXrfJ3z948e4
yJd7MuiqkVoHvKuFa8d+UNSZ8HLXMrSq14nVDIvp5OktUjs/mirDnjWecvNhE4Z0qE00oNyU4o7d
J5+o3JMMddG8J2oSJMBEkaw/NECp4KwhoQpKXHDVH+OoIwOsx/1dckyCHw3bfEZWOzG7c7HYFuef
AjMmSfIodtD+e+iq9VIIKI3yEogmqLgv/gweunjYXRSvYdclPpgk24UplequCe/pU55FljoLAq4m
S4maE0UrdT82BvsU68tTQFPuZcLKrjwERdcR3iU4sE0HBL3pJ1Fkuvrj34WvGPq8fWVp/jIzJ5hg
YHZGs7evoZ62XN1NAiYOkd7Ul3J1t1vkH7cdeveQiGq7FeNNXACEIUsTgs2YszsvHlmN8YRm7FWE
pKmy9q9D4aKDowPfX9rQU0y3+Lt2Dl7sNpBieWVN/5Cq92VjtqbgzsnBHd7MeAv757iBUI9LLLep
DgVA5+UkIFF4yeWPeqxhrK0doNrcTIG2rmTVOnHmS8MA78ngCRPs+8T7StvdzRmfjDCYdPq61gww
mwzKJ2XiZLJQulkHcEubAPwRNRYAvftnHTatnSuWrebDe5nAWV1eX8TC12S5S5Wzcftqq16Lh0QE
g704gGbR1JFc9SDKUMLDcPKioKLFRqpnm373d9tGgMBUA4Kn/5DptGO/nGk/kytmDpYA0Ve45G4C
JB9Iz0meKl/8PhTMVRBo2nkqs+GIDDEu1dWxuinbUaT1rqIZ6LKJ9eCtfw+JD6vE2ZSD5zwQ/WLw
eA/DnUKTE6pXbYk0NwgAR6QtcYb1F1DQClChiXomXxWx656ueJ2CJi3/KngmADKfPTirmnAXjPYq
pFqAzlftn64Nn0E7hb/8gI77gNT3769DP3ObCOqgBNCaPoGyX2mT43cYx4oXk4mjEi/+/A5f+8Gp
Jfp6VByNvl5lKiiUkfdmUsNrCSwURI8s0dh0lr7GeasJWDCSPv8GoYboLhD0C9ipDYzpAf2dnbN2
/lyez0/ZH5h1v/5noBx6jGD0AnBXSGXmJ3BaPQcFNsjEeaRb44Rgv6O+C0+UidxlfEUJP0Us+7HL
KOCIZAd3CvciIj4tKEgH4ZUy73mqgLAKqcboDLDdNPJPGY58Cjoq1FCrQUjDuZpLGuJzalwT29V8
tmRcZ3Ox+2+dIXFoD5s+ITRiYFtmeyiGITxIJRQMBvIWh3yf6Ns9NUV5ZfXXu8QMG/vCCMGqWSEf
mFqvq6BUvwbrQ/Jts9lSjT1xtWTXEVpqfy+vNug++CYR9tParxhgA2JtF5avQCFNAlOj/0OiUOnY
O4zwm3n4Rvc+nVxYdP+zGgCGwOABvuc4tg9J9lPWNjXagerC33AyWhqZSptwA2Io5j4H/G9w54ae
6abbcR85SYRQqIMkcSQePm1cMJUaCYmC9jNwSq0HPvIUieTw5R28mdbLLpLuSzylwoITxsHLdv8t
fQEcjHWSp4upa0sY5PvEeOpMMUDORt7rbhl/GqSAWAOFZGgzwGatl6juXYmCCwcTCnYQZM1NYASG
5vrPLUTFtRKKJ06VElL+AUFKZVyxBgzLzDJOeVtoPjr4tqtc5k9ENO9bHiVbxIfJFN3j/G3QZxDl
SXfW8GQzEdcXfd1Om5XLkiFlHpqae45rXgH1BI2TmNJpsMiB1QB/XNBmSck7reR5VN60ZgLC2uJ2
U8zQcCqeAOXU3YD1w80I4B7ysy8m7l9ws1yYwMe0uj5c0HmPH8zcyuvrb02Kwyrs9kC/hOxgsE0a
EIaXq2baa5IDoRYeFbeYS61K61vkikYbXELHvI//Uk1WRoKiL5f/m5bFnYx90Uj77T1bWLeiUdhX
3TSMJ+XKbmb3cEmfQ9kE6Pe2F8dCltZCx7qO5W78H4OAwffI66B/7lLHKb1CKB2JL4CYHrMXDPfn
ps4LDK2ltobKV9gFa/OlW2NIJVjeufeG0sCuteK29xPgXK3TBk15lYE5GhdTv/LcSEhS7V/2ikd+
3RP/tJ3Bh9/CeqQtMrx4u7cNdbN36R7jdbzU0OdCEEwSfo4k+A679Pj7ghbIAer3YjS48Ke3QQkD
roy0ilpjvJcQMAurlhBeGcN38LEpVM/p5Gc7ywIoYgrhrfmOTK9GOSqDgmJRl9oFntp/c9Rgii2X
jrhRtY9Yb3+RPqYi8r12F02fddI2TT+VTs8C5f1HLGt/vK8/FNrhmOy+GnUynjzuIYpu8WmW8vtD
vVTZX+znm7mVHbvR/FFmLllarS+ZOT7kBipbbVU3OqXKA91Za1puEFcg5hWkwzJRznfLqGbsTfDN
EYsQza4b1LpWb+vIBpqDjdb2gyCq+uNL7IUGSQoMOmodc9Zv5j9axlr6m1g1VXv3MO3rHPEHH2tF
GikAkmQxH57M9sJ2ObrKxmaTBeF+I+nswmFxjnrFwOM6jR7s0VUurAk4kQoSxRhB2mb5cvENMZHk
tPV9Sic0LT+vZbr+0NLXhfXhJqiZ96A3Pi0xyJdfUcvyJtdQ9khAgnTFM/xxa9PGh9tYVfnSRUBT
t++AioYE2sPAJq+WAY0NwXM4oLwhk/ZoBBAZrGm16QtYaM9aDvwA+rMgCgjx6hOvirTSEG+z14Ua
sX+qkW1diqlZfL++eIGBdoyhU0K+RCXOMkDBJJacTIHnaE6x2xVkenT25D/yCP4jDbMmg5mdTb94
l5du8xlEF/JuxD2VHz59XZX070r5vMm4rpJ3tPhck33IfzefHp3K9ExHqKGVcd0pBs5FMQuJk8jr
MvaaZe9FiahHQX+C/otEA56/Nm3EEteGlSoDw2JeXFoUEOdPkeHWYo/FdFkwe7akt6rHB3lPE5XQ
c62SrGVV8fRX5F0RJpJ/18YrGgZ9kc5N2pld2JQlQVGV6Rc2grtQUm7S3viOomnnCUxucBj9bZL5
+tcX01tqoA3Rln6Tn2xWThEckWlfStDONpJSJ5EncXa58w6xeS8L0TGpJF43AuiySeC9u8wFShj1
wPZj/rlERVq1gfzQZ7F+CwlA8tk1XkFMH+SWBq7NJGyK+9GkJ9Je1V3qznRH3ArMrAzxf7CINw/C
+i8Pi0tLKN6HHK+V084oB++J7WWYrqTryz8TS75n6z1le4Ji4hF4thwZIv5GcXWP9MvlP2B0/MoJ
QY7HGVSU/737fp/TPrmU4ZBSY3DF3/aXAGeAStAvY4cg2FHDPkVigQhw6jr3sfrITjzMkEVYRCCD
UoCzKcORXf7p1LGxeZbhtLN4ysW/NiEafscbeVQ6NnELjmYUBImrlDPxKVb+mk+/6dB+umsJimz9
kuYapD8VKhLc1hlI7hi+Vf2Tdbwdvmme0p9NvK+xjDDzyXsJB2mnWPvIerpGE8FyeQMcaIPgvQiz
fUmmt4Z6gXBCYMX4s66udfH5AeFZtcNy7uWVvV7gsyJxLV1FZeFdkwtOCBD287aKQkQnmYqG9Kzd
+1V5Fx+A3w4eCIyZcW8S3LQR3ECbsLDacrh3vS5ImRvXfkR2V8aJyh2Bj7h33ZEBL9cyQCKSL58x
fANiPr6k3TUr40XX5EEZ1WE742AA49DRDoOMvjpZRqtxBAVPbvJCk0Vs6EHDL7WqH0ZTzY643APs
qa9K6mDXfpvix5J7t2aCNfJXyDLluhXw7ANIVfHJmvLfwWRAVv4E0Wq252/HcEQKIHEHRLnHC+WR
jjJZTlKCaOFu6V2NcirEjXFdfdBLBKYwjqeE+ZAOLd/VPs5PEtLqJR7h7zG2707iYkaXjT8gPeHL
kD7WfQv1nHn0uOaK9oMbTwATU8TCS5vLrKj9cVpSk8Waqc7CQhzpNZpn/E5HH6nDkrDpGpZBL2tV
GbF7q/geIUGTIVoDVK6uiFQuy8Kyhb62/cLxT9gIX4s4HYl2ACE6HEuQXqfOXrIeC1aBZm32Cp73
uQEi6+4kAgTg/R7mgDDbBL5b6dgK+0GJ3+vtMS0pfGtOD0WpYf7RGouLNC3+m7+HNSyB5kRgKr0O
LL1/TP2OcrWUTpkCoszQhqYpm2jAFNSpqeUFyYD5S6Tfza1yVfVCzvaKLhYwowxlwiqG102tQ5Bz
H5tkdNYDXjk/mVrifxq9jUHdPPCrj7RGUK/zYxoXs4OxEwHdVEyLfG/sH4CKXtGw6RQikvU5GBHx
1UrjA66BLSOoQxroUEJMvz5hgx0MSNBnd4o6f4pJfGCw/O9VIx+UiUFLnIfrBzbD8cC5ziSlV5Jl
c7OTfwtZzQE+B3IpfbV4eTGpUpzBMkwFkrux4ZJPBHAC5iTXWC8LzvIdqzHH+GpU+3qD96Yc+9CK
Eb54pyYyqwzaXfQVD86BzavRTEUBfRkXfkszxjoBJaphxoiwWVCKy2PClnBnW5f9CotlI2GxIpal
Js6d6Hk9u5fuoyRouCKez27LpNfQaqblsdeVg24MC5ihDEMRcdPnCNzmR1sKHR3+PJOMh4uJWvMA
bEPwIHUjjSzEucLsM2uZiOdKfVQt2hgTZdfpkxPgm4H0c36do72ATkutf8x4AiBVr1PKn6gdGuK9
KXqYfn5ydYPbjc0oUCSWgBfIl1tGbbfNgk4YuWWl4jiYZrv+EkOTBCO11HdrDvaqdbyBZbvNEneb
FMoTUWYhlL8+Jx3BIIyREDdkHF1ax8TrWd/ECR7xBbtI58jl1Wkn1SnSE0/kyZwalFCDRohtXv8x
nxFpBj4uPpOJWkDBy2t2hRBaki0ptGnk2G/YjnRHmAGylMo1aLn3zzVIQPvixJ15deXB15khD8XX
ZNo1z7tthiy6H1oFrxP5r3NZHBulhQbZQ6vLcoOX4rilASX/NRuu9pSOP2Yl8mBGe0tH+3lbAyHc
/WhgtWvo5zru6xY1oPEhox7QGpt8+Te7rfCcPNoq6+zn6vly4PQDu64FxbbUhwtRLKJNGg/xYigR
VqnnvN3hr6rcPkNWOJMHcevmOTW/NUwhJ7U9oobJYPhwHD9f75tsc1WHSDeRbg6fMo06qfzGH2PU
xv4U9yppz8bgofRFMJMpaHWt2OZbHbCqwtu7WpDCql+xt2aYoQV9pjTApLK+rsJvtpIwOkhCWWVt
7ZRgGHh2hiGnYml61YLv4AHu+SVZwCyqNR8e71waSEiKmlDZYAR54OvxICLpgXp9OAj2gBdKvPmQ
XsUzhOxli2PC7xnUb567G5y2GL4dZx3O53DQUMc1EMO+3GigeXmKZlIOf1PeXoqDq/h8WW/Y8Dwi
IDCRS7SBql9u8C5LXJZqVGQ3nZhDP/DyrkRez9hhhMoJL/PjQwiSuGPBB9nn0jvkj0BuZjKAmaHv
oxSlkHhprs6fhAjlWuDWJIOTqxi9z6KTXwU/ml47+BUkQFx+N5zDwU8LV3gMxvU0kYiI/vrodi47
y84GXTGmx/jYbO5I53O0UqhCHSPashAVfOrMiuBLeG/pmQoCi39YbeUn6eT42mKG/BzIxdytYUcj
x0cqOTZ76TgL7z/389h9rJQMjox3Rh2tGRp7rDukZbPivaDMTZkP3RSXaxd2Y3D0m/xdIgqHseyI
doX1tnh1E9EiM+DzI+xNlvAj8kP9Z1vFghklh81D8fdls/nH3pY7EareqF5p6GCkp00mIL1NirPk
rBbvZpi1svrYEtTGntAJxxypgP+rpJzPXwYogwmyV4shoTuq2BELdR886J/b5yrqfHgR/cgDi2fs
hE3EhYfm5AczUr4uXfG4RLpcfx6YU92CaIStjt25g0IcILJYf5cZRhl3fwrHNVWExFZChaS1DoEt
w3KankXYj8wd1XVCXrRMSjNYsyMOlt4FqpIKUGoMtm8+7Xh9ev8+2tFzLm89YRDJnKwExhoW/VIs
JTSKkBBxzGst3g/Rjofmdcfxqj0C2FITCfl3fhLhAObHwqcaK3HVOOsHqMauoSZ3BPq3yuEIaX03
sO7FKDxN1akPODiqBerZE2JqxCSB1vFaDdJovNforXaVl/3f6OWyz3vl7uRqC1Zs7V/qglNNqicf
7EQnQW+VeX6XKPt0aowPuFp7qK2BeyOaNSfoTYb0E5AEvkHacVcjuGKhj+QrfMHAaSs+YIEeSw60
0fL1TSUHKx9Ho0zLcui1zwIuKs/Tfv3ZI7xTMGfPMzwhGayes5Kzuo8mqanBiT02menDK1lVmkzh
CxJwW6F6HClBOKdx8qyJIsa6/fzdjsUdQ5E0pcJx6P3KjKBfOntoTKwoNCvNGzxVw9CavbyhenGe
7dWrsSZ6hRtoCSXnt4j7M/thW8Pjb25OyoTfy4hN7baUcFiQDb3MZQ3H0ZewnScZJ9sSc2D/VgAI
evGvhHrkMqRghW4y8A6ppo2u/o6/HFSOWLDE8JIjta84ZHAl8WB/rzPe87929r4pXx8Fc/nP//7W
9WAnq314qSRU6rJMj1L9A/4X1z32ufK8L4xCpw0ZrmVq7ew0AjQVcduyBUzlwbUw3smFpjSr9BUT
c+FzGiKsych9gJahQpFIgzTZySbCAHXyG2v0gRZILEWSLsQIH+iUJWuUJA6Ns43BBU/MPohl59JI
fCGN2/fGCuosgM7BqqZ4kQJX0rCxnoUvyJvgljnsK3ANP52u+WgGWnX4XWUxP5B8x+SJkkNbFOLm
tTXSJiEsbO39do60fC6pVWdH5OZ7SoRkSl00BXiCnVL/f4sk7sW9kggprlyTq0x3AgRjpmCUrqEN
LReCF3Oi4vA0I6zv3ncLaCWxc6ADfSKYeoyspsWKqLOfnYoSasR3KvEzQ/YUapftZJvAK5iqtRtO
Zaz5ZxqvfwmfUme+bBnS8dk3W5DNoINfxggXM88akKdut61qLabQPxruetcF3a1g+jbbcMme+eRq
miWfFQR3P0IP72C1cQxCGr2iZLx3WN/6t29l6Yd8r05fcDGMpFssAsApFq9gTKL+9PkeTRmt2hxu
vy75fYL7/8dr998QoCvXskzl9loFfzFYAQUEolGcD1tNmENNoKkNrur+rGp16xn/S96IssyLej9K
FoVR80TV7h+MTeKP7TlzqP38Fw/9/eP9EQw9zgDd2n1hDDXoMPoB3BepGnq5u2L1wK3OkiTOoeHo
Xv8GkrnBHEh3749LnE4yS29p5XoJ5hfmrNWAdgzlE++6HcllSw8GVrCIkWcv8/AXUxTpi82yf4xo
SME9rcI5lJVnkIEqpLNDiEyKP33wLGYukS5SFOi7/8FTdA0g20GAVkreKmd2RY78rII2xdOQAHht
bGJs3PebjL2ijYV2KTwceQ7qzHy58eXYFtXfxC7e2Zg61WOpIVcBWwtxMDQSE+suromBgpOJAVaz
f1hTqSJhI/QSGHdLrXt7XJ+q/uX69nU7Q+sNMXM9syZvlnA+aNJ2Ytd12g6rgQDFknLtFM1Abt8H
CCMjIUvPxvKV8YtMvWY9S5cww1+iZslQ34t1eDpC6RjWTxlCIqswLQSv0B4VfQ/XlhZy4wfWp6se
40NIccXZEIPk+vx6pFIZukOH2YRZy6swEhzJHO5ej6JTCvsP6NDgSQr6dctykNUg0xs0m3tXozwe
9AkCB25nCUZ1OjMEL5X2BsHAfbzRcOpCGrQIPbDRn2snDMobjAhb45y/roOht7E3KftDtfog73Fp
Z+uez/PsqwPMp5yGCjxOyV6b6Cf876Wxq/LNyYU6EvXOvz2PShhRQixRO5LB0pICuDl4+JhZB3gI
xeXV0p3qcV4nciyj3+JhEb6Y2+tYkluCRMEGsfhZ684n1IfWLVecAPiRB4WMOqYpsJOgCNNlpxo0
Oc+Xs7Y79DOCrn3bn41WmvVUeOOQuNuBRYH6E29V27J4CpxQD57WeS6SFNMwhNv1KvT169BrpSdO
/WFs9MdNUYnK5xsynginKASF39h+LRE6nAztOt1MThh70ZLLMwxPkxNsX1xscvFFLmUzwjk1H81X
fa9iW+S/hB/PosR45mQ3LzFvNmemxowSc1tVAX3xQ60ghu/xD3IUq4dnLl8VotQ1ejFJ1iYTEjW8
y8LeuNRUChM9LBT/Wg0HENbf6i220/edHsW70yePeL5KsRVfAkc017/siB+DIDLzdEQ+WTzQ3v+A
W/sWoian1aVH6arBDGqBCw0p4KIixO3DSE990+55hKOen28NFOZ5zeYMvXg1a5XH9rptu0cCS+Cv
sywotPx5+sk2zzCFVfCHhDIfu15Ndqg16c1Zpj+W9W69aYDITdYVpKt2UM702TX3k2iaL0GUdnRt
OrZw52tKsMSeE5HSiP4qIlVcrqNokCZPgHs5puA9XBVAdki1cJiZwYsodht/nfigPz5+0UgrU6qW
C1smsyk7rsVEdmmS+2hRl+jAjiogOyl++JRDlXndWZl5arPGdNkO27XCaocdfH3dJ8Mp6/5+8IdX
fExYrHF/FDbp9FQFp0JEQQ2P67PDvYSZSx7BkT5CkyW3U9ML7kqPB1n+S2yUqX2uuWGs9hirsEcC
4YVYotbXaaB8qTw8Q4bTxp6mRzjtw0uZeQOifYE+0yVlQLxVBdHdOeusMtgdDtFfxR/BEwNDcpT4
uxzgyne/YzzMbA6TYU6WnV34IG7KS/bmPitDrmf3+83K9r8Go8hsBk/r0/PE81sXMCbkOK27sLyC
IoVQczZtS5jGoYj2/Fb1Z5/phOuJYik6t8/n8MPQSS2l98Sk251ehvIxRc62KsML0jVhJVu+4Vrk
ObKnfe2c5GNQIijbClCUY/vZD9piDB2CHeztIeXSUn30ErXeQ7cNRqe72i2628hcWtV09PtwZrR/
5DLc3ka6H+KUqzeByoJxIVcRG8q76lXytvXScWp6Qvl5b9JAL6hJwV0SBO2wZe9fxuHeoDFndOVq
raXRxXLdMU8KFmYAJ7R1NSolTwE27/QBpl+eMCaHmBBFwaA2Y5w5dqdejxCjqqZqYEDgdOCsIXjD
BQKsAoYUnWLbOWRucot+tSG3/rAePu4SC1AXg+P4hR/NK2gl862gU86Tc7r8QA0lkYqrMfXQsdcq
gp7IuZi5B/u9xnC+plGyFrUzpTOg22ObksvGtHAWPat0wljhFrgHgWFWsqv/Gf0V7Au4Ka5LfiIQ
8eqtTdVyV+3H8JvimkHseKoBSORkA9MFS35XRl5DXYCFe7eVZTufS8KkPgQCFsf0TjkfFui2bBN0
0cMq07IABy8GDSyDG0fgrZW8gda1mWWDgfdEg05A0AZ8Uwa+l5qD/r9a3ximY+Z4yE2OlTMnerFk
K3DIZ3jhb+xcjGoVuAFE5zsTvARXjxawXdSCTpwFjrEV7dBk4V0k7lWQ08acHt+AjtlrlcLbCBgZ
hsQEjUF1sXWHUbgknM6A/GDMOgL8JVix0zA/cF8wn43p+zv7lNxwxhjuJhbBN939n18pzHbf6/0g
XN8n2PtdBdPcNSW3mFOXPMu8CVI9bwTxvuWNEoSKeyoH2gEkXKOZ9yCuDl2xEAuzr+JxkI6pLoiO
MXTITVP9rPPjsCXgUvXaCYxkdZ+yYIhxrqGxFYVVbbCfc3NBZvDGHb68Hl727A+hbcfWmM6R/GVX
brM9GLKk2jYWbjKbtozZae2ACcuuA47xbD+rcMlMDGCBSBrE6Li81rmpxD7XZP/pz4WtzlTdRZmO
GAndYACBEQ7RRg2qubI9450gJliM5mbUckS+ys5n2MQQBqqVbKqxTv0H4bBvPgvPBllOhzt+2Pys
94Kl5oQpanWSi20IS87hiAeVZxcWvYkrlEBQjFqOaTqbEbJiIwAAuq8fZLtOUsZHWFg1vUBWZR6M
YXBkbdzNkP4Fl4fu/FCumyrK00uEZcd2iVP+1kz0vlwUEaCb3pfjCXRMNX5oNuWzryfJrIvhn/tZ
fc27hrz5+U1QDNBNIBxVVe9UZ+VW0NAsl+AHyKhZChHD0j4ptSSEKx25IM6ZRk3spt6+rTxiwoo6
xaH7hoOE7EIi/iYD4JOTE1qlK3LQklkwx1T9w63aqmN2THr78XKqQqBWwiPuZQB3OPBXDkOcyrQG
hQyhaRnZYsk/Z8ELhmeKMV9KMeq3T5GADEdCUHPFJUXnhzwD1TazVJqYPms8XuPaFYUEyzWx/evc
ZP8mngKGuO6GF760RBu3qA9M1jQw6RSOMA8SvSkdCdInE23bsd3HFqYvYdkbMSDy5csMdcVDK9wv
rVxqOFe/42itHvOTMicw7ou8SKJC9Obbifc5GjVfGiPlk7hlgm1IKo1jafy0NImvcM2wXtnmADNK
rX3DwpX4FA1YOnaY3mshsTelnGdovSRjAMVaD95mU6KYaulA0Q3r/n98i8+TBVgJru17EM9UDc+P
uNrm43tlgEr5PEBTQvHtjjKCS6EtrNw0bYlG1oIu8vpZyLl7gMQnV1xZNLNXijVgaPDxciuUAiSF
wizDbSKbm+kYomI/gjnTtx4j4JgXX8n6bPofoHeYoIHse212tEBmCpZVHV0FvqTBOk/QnpegaM3X
cYnEGD60QSPvpiRuOxXtN8XU8vWJh59aSlU8YPbLiE+E7ib23bqgpwApk/mM1iltOgefy1pucMR1
1wtT1DLUT5VVFZAbqNPd8J3HqA5ftNkuT8uHCnv5mlBcpJqTNPSoqP32vppWbF4ZFA9lRNydVanA
HuMyuK2QbYGvgnkdgEBFRQAdxI1M1sWnbQFOAzEOrNt34Ge9kH13P6GTKye4/aIULMosMIysRDgd
xSbIu+diDAfd2Lc5KM2aIkUH4BaIi48s+ymQaZrOkA2dVXmdCNtkd431fo/Gzygtz11JNbvL6eIX
XnPAbar87vU2m/aYUGwoR5su8jbwft8rd6vre+6ceJLjVdV5aFAcDaNEDSoMTtz8SnzK3r8LiVPL
B6BeDIazyIffcgqPPw8C6RL+IPACNDcTWj/44+8/whiKqooXd18x2L1vOj6Q4ilIPtsEp+E8j4/T
B7U5nZmLdG9pSTBf6/L4M8f37qQCK05JkAClUTqm4ilecVrgwIALuiUr5guu2hPNXgg3/nvTbe5g
mlqZWHOdlL+vfjxwB1pu1AKFXFcTUFT8a9D9yDpbuQ+TD+iRQdjLS3RBrAjLP6gZgJqNSpeN0n02
ULuIb7li9cYsMAX95RCW4ErRkUVcNLteD8+cXvBBEqoUuhs+CTBLhHtYw6bRQQEp+/JMGxIPZ1R8
WuzExHF5SSzzSdJvJ09g4nNUdAtu/a+gRwv2/O4Bj13Tk9zYErD+Fq5dXi6CljA+7IxVWHE1U+KH
89lIDNjJ++OE/zNFTO+RtIEFJkMCHjBkNfirkgLL5FlyDVe6Yu+OUnEQ3tlCCZI0CzgeaUMAPnCA
fD+Y8Pr3uKVwIGaHPNfnwrreftkB3xTOCEk4Ke6VPtVgeFHymhE9M8uUg/aqDBFpjHltdGSs9xuK
ZTjo2ej/FWW7w6CrSorwdzgHkEak6eV9GPW3LgfUoH9LErpF0PwY4/ahs2DKGnGIZHhVH8WL8bBD
YYXfrBOcDLY7iCnbdXmt7MTqVqlXeZHZEa1/FIfnt0NaVN5/4CjW9usokB/Ml0tUsERmLBIxwUen
Zu6Uc26TAJYUKJkSt+a6+qz2rJDpW6THhWMPkUmnNHn14jGfkeNz+CgQeHy5ZZczjFgKbtjlkXCO
gwnJYdb6SYVwsodpsoRhk9/9M0nc72/XAlbL+R3OnhHk1xdgrgp50G3NeALJEbZP+HaZ/9B13mRP
7ryUGjZvZn8rgt/MbzkOP8Vjyw2r5FzYbYLm42zOgMrGyGV8ltwPVxzluRDnr6/HgjeZu+zfLufm
xY+lwCD+wF3/JggkElYbVDWyddwo68eki/mVcOAMb5PT0dYLo9pb8BjbeUusceB3HAxzdZxA7Z06
LhWEeG6/QgIFphGkB4SYfrybqW+Y5ICero6SXWWZm3nc8mwnm41pdQr75YyO4BWfewj4OaxWaR0s
JrT2EQXjIKHsz5A+oipl3cpkkKmdV5O/xNcxDlGKl+r0dVXovIaengU7PacIrZzvUizXdmNAFQjb
LqYv42+4dVGwJn48fOD1I802041Vuyq+wP/TrpZRgB/iSKtQXwousV/qQX4PL+TIwTqPHWch2V5Z
gUZaUnCM0BDycuXDjqg+ADetO35ttK5ekvMaGvgdGGkLvMz68wBTJdtxxae/My4y3Df4JdTXRR67
NrdMsP5TtAzGxWxoUsPcByMiMAxmnfYAPKX2vdQ/yu6d8ueZkm0aYCynC1+7sQea2BJOQc+QgB0N
KxHAt22LtjVjcWsLV5Eul+tJsaQQAZSxUZFNYT3ty7ytYSsMjzfkVXpuDqZg8HEY8AFZjm95spFU
vWXalJDKnCUb2+Bz3Zli3N5qafITKEHiF2ES5MR2bYeHTAn9as+ZkFB+0gxpJMXnmsl9/H06Jcoj
6+b2dNYHtX+TqGLjNGCEWsVKoNM5p9FY1jU8dnza7WfU6oV6Gy2jy59O09y9aQAavHkSJ/qLPGfK
kN6uh8HFmCGWPkioOLV59ka41Uub8NVRBg/kvojMsRCpBKnJ2jLlEHeeJqhd8UkOAxl2GLqKGl9p
w4XlyGTKpk2sYyJq1dsxVryr1Q+BCfhQH1edxYoxfeLzfA+pRU3lpyvAPU7CJZMDzLsu5wghOkCQ
Iz1NeN4fN3EC3ZjJmOh5bJGCZ8dDGvu9nXvoG+tI00ffS47CP7nlpmIC7yNhxQHnWKZilQoKsLIK
JZCKADrZAxY3JccgryIoussN/rmlNBKSqbGrhlh2vQD6Y0WdZZtw1ElD1Czz3S4U5gHqw73JElyT
ewluBIoYi6V6p8ilOoBFtbVPNmSQA2RTckXCxacpP99lCJtRWZldtGph3zjHEvdnycNT4hKu/57B
TSKRhJXud9oprJn4aHJgS+NQuEjBewvwSos08F5q84TUPwghyqH3rYMo13oRHIcTc6q5OShqVkBC
zhFvtGFUR8brQIqxIWBCOUQbTH16y1T/vNIk3vKfhvL0iAe7qOMwgWvdGDwoTrVM4Ee2Sz2r4HmQ
n2Eh6Y1FuI3v4wxZhlS/O/3pQSZRaEWPtSw2Zu4CgOIwaOCmUsmS8owaO+W00TTnOhM5d+h7Em1/
rHcd0hTFBfeCjV/u8vltA/52TLF8TZscINc43AqON80f+8UCi0+3S6YYOAdT70TOzAggchLS1AyC
6uOaFNmgISBsu9GlTICumQJz1OgrQHoztMIp5Qi+Isr9Ce/bDuoTqN+3U5ea+qyP0fcFBDNdTM4E
ZDXn8xVip5Op3H8KAfXD1Aw5QhIjvhc4HUb7Zz5wdXePbqodStFZcKKKLXFpQyQ1hQI2RqqWd/nv
ufhAruifyNWzTfbZWCJg0hE38FrhIssXsaMPrUt5+5Bfs/7yJGkhm1XdaEwEu2hlyoyHiB+VbJud
ULuw6YSFhlbDY42MTOZNoTI+WF6Ul2AzsNKwNeZUKEFLLb25fAhVUrCYZyMj3f7PJdeH3OnDR16e
sp1jKxpn/3zm9OrmLU5fIgbuITFzNdYZJj6bqR1y2iU7FFlTH2ayUBdiKm61nfsPD7DX9RzZWqf1
UkCEWsRreawAifwHssPrj7b7mdQHMvZs/+clNOeSeEROoUbaKZIRSts3JyNlb8YTE7BT9MeQhPyx
Uk2j2t9X0ZBVwUcgqbU+UpxeKZNeDpBGnLbVIBVAMm152L8Adcc/wgglFhSO7hzwXW7Qhom9a1E3
mI0iH36HzUivcYBqrr8m4VMBiMaT/Q6OBKWkpDOfBrZ78bePgE7g5Pr/XKVw3FiWkmjDKrN/JN4i
9jCX6F9WkblGtMKJeZdu5OlqC/rPEsyvT7yRrLB2j3doLcN7YP9+l2WZPjp6Tbi2J59Wj7BARY/d
W9AorjN8d6n6sRtwX6CX7UNG5TOFRMacaAP3Z+qAtaIuTNzgEwc6GgmCKvvBn3ijjy2uGHYmbId0
OeAhtpVUtvK6UdLsvE7mcY7keZNtP732Mjqt1M7EbMc5p6b84Tyhwbwdt3a6UirRhIOUQ8Td6BXd
HjGSc3Le8JN14idFyVQKf4toqqs/V32NxCrQ4bTfQIechEw0WughbyzssTuWeDf34scCCqr9a4pa
BxUqg5AlUEW5bnTinsUbHryou4X/1Gw6+bJG+E3/BBg3xSr/2D9+wcxpwjHsTHpAG+kCB9OvePAI
bxsdizVQGwbwCMGSRhdOWrzTlAfyK4mCi/Fkl6kn55QaJnLURDcaw0rPvZCTwenv5yGT0j9bs5tU
jacCK0cbGmMu02x8RhLpyhwtjCZxF2aXlESm1lDT4jxfbfjCCeeNlvSSecMykcm67P4qsou8Ost5
5ZJevncNSi5C5PH/hts5GHrulLisJWHrK7PrqQ4xQgvcxt3XGOMpxB2Pfb9qK287Duyv5xTjtTuu
FGV4UQ45enPqzljDSv4j+VQirZQd6pYLz1uIg5TdQQATQKCr51ms8XwY+KBILa4u1OqvRIh2TOFr
qfXMarobTITkswBUgQnqd8PonW2RWfmsQK3LqXD10Hq3Frif/EkkKSCk1sq6aXySMlKDgQaAzUZl
F0j4lgG0O6aSQbDkQHU87EcWBc45VkUp0J5AfPFLKozVYzRrZgdgRhsHKYP3Srw0pXAvr3hOncsn
+jlaTa8MzyH5mKunhMU9aZI7qW+f1Gw5ZKq5cStCMeUM5j29E0VAcisJwjsn1+3vamYCJa/1Dt2F
nKhqgKQvRswYPGN1wWJFuDR9NZy0CFDd+A15Nn5EyGdco8nVrWg2oM/ZTdLf2qUaY3YXvMgB726h
I4DnjIuPOybiuEzFynh50R8L+a/q/6Yi+lKjkgoSpPRezuGicdf1XdEKD3pNROjqTN7srIimhqJ7
C5XFKGdqX3HUD2IlE8uBJXuKe7hSLI6ms+0iBVoOaztQI3SGWCmRC2C/0G1XltN+k/sSnXh5sf+r
bMjNRrzS4JJeRckiCZ77txwczAVjj2w4AZduccfeN0+G3zjUIXnH4AFO+z0Z37gL2xWpYw32G8lX
mP2vK2D1dvifiuPRtVvNuTwXGwIhh2eYTFzXoXhRGGSq08+SdQONEuTpSr/IAAxHJiKYvWQB7Eq9
YAMf3zV4FrihdMHxOMwnvrK8htaHZEEwAqfDYwzjuQu7fIxqLLz83hXGIE+JaCG2IMHMTAWq05Fd
bGrx3zG00ZxF3G1+zcBpgkH1ketHTPbmK1k/LuruzothnWu0i7hKnL2xTTeGNoC9hTD9WVQWy3bv
AO49DcxbgIkAqCnuNaDZ2HgOeeYEpx5Lbs53xCO90e5J1+acLmPaJ1V4bow1KiqNSrgIEB+y5bEp
queWuCI+YhfhMrvdiQYUJi0IEcfitHPepcme0Vc7WaaijFkigJTYmJuRmqFjd49x9B1Z67aHVxIF
4WKbXjfO0Pyq9WVH3nmBtqKgFDEnKtxcc7zvQgALzN+zLIuBRPpF7whtaXbTt9/U4drm7anCFPXb
GbYhZPmKH5ZMBu8ioeVEALpp5CdxBM6v8EeS1L3DkxVLjcUwTnA+EimhAdVfNLG5My3bwZN7BD8g
ga+a87NRaxZ8mdXj8lF66bGMMXyqWfWywYbOxuVKsp8odbpdrFjDxuonS3j3Mb0MNGfSZThag3IQ
wO/2eFAB8YKf+s0Y9B14oOJJsgDYYEhu7Jti75iaaLXKKPOu7hBcAYcLoAl2MHKdCWjye8fVqubH
Uy0BrfESk6Iw/DVh+vvh86l9tAgSZBvF/x6gK0letE7vb0HQzfLHrm3LHuvI8L2t5FGr9InaHHrS
cu0eauVmc8FMBfu5caNQor6eppPOQWzTvxM8s3tCM9Noj+bl76O/6uI29z0brAM8hK72DDKFigZ5
YqHeHfFnUxsH1JXyJJzVzs1G3Uxu4gfZuMKy6plYkRSGBFNcAmOnaYiADRfo8BFAdHs2wdhkAux1
YJfD101dvo5kSByD8u33jjIoFH7S97nnPrE6yjO0eQOI69r1OohXgEyHK/bPOL85utAmDk7+Wsrn
f2AMK6Kq7FeHut5TQiJHuT0mnYBWKgc9cUllesZJmbWpN0BQvdZR/QUe7xx5B0+oHNyF2yPyLSSa
fBYTrtkM8N8NXIjoaMNhZHT4ZMP7/FpjNjzgWOlj+3CYZn16/19o89bIAHGcnetX7yzqiXDyXcIO
ll05pIvCEslTea0gaWv+Hgh91TRAch4nHjOoTUSucGw2pOuPmF2nq7XbvcWwR4KlpBhmN9T1a2tP
eP4pK72WH4RDwuDIZSwVFLSVaB2pgyv+ZQssLMHA3WkR5DrXuZEnbP93OoxkAm2+hD0RY32WEkDY
CL6IuBIl/I29IVyna0kwhSDeIuBM5II++85Bi7qn998J92r/ykUtFViXv8Ju7r1OO6Htr+ioo9lu
vWj1fVYQ9283bHUxTIEKyGZHhBTwerNDSgs0bbV7z/5RWk1ZgmWKngUJhH0uak1INACpzvynHPe7
a2TjC34nI1u9oQbi/CCh/fr5SuTm/tQCOp7poAJtwTHD6Gky89oAWstuDPWtr+HCagiuQy6Tddda
8vZrPMHFukPCViEiVSM2Qdot2yQTnl038LZPeXc3UQeI4kach+y7QThGuy76b1FOdBP7xqEJ5X+J
rEsO2qvjpNkE3avy+98kQXv/711sUYoliJI7m4zXd3jWM/nU0tWn3sdhc1TCEIJPxvjak8J/WOGX
GxX5DZUt35oOwkM3N8lFwFacTP5hpccOAnRcy91Y/wqMKMfr1oWvVssbrT0xgIFun/h+4nOTOk7o
hGwRPaPBs6KhLL73tMVRP1YeWwCJ9suCfSKCp3cUj7nvcbwQVu6bYZzHgoOOBszWAJtcdnHhvT7p
EsaZPDUzq2FOZJa5udXV08zzq4cqsOgGw/T9mfHb0qYqAJyq8tueAu58Zkbm/6Y7FPnPyR0u6ph5
Rfza2ELs2a/LpTL0bA+WpktSEoT9zjybXvI3SdzfTUKsNqF933kSGlmBzf0eeSr8m2G1wKoRO2zF
B7Qv8a/ab5BVeIx+ga2CZg6n+TDYbmmhEyNde0F//X0pkz6zTTFhqMXE/g+9zkpaONEpfTsctTMm
DjwbABOqm3lzA09R3X8ykNtUVdxFfPAiZli9DcMVT+cU3xOXKaQDYXexsy/Ik1hrYgNa0rMvJB8Y
QrTPnQrrsaPJbSslulnO2zIkAIwwIfWbmDqxEFdz0rWEVnjFPqmwnDp4wIcZWmBU6fd/BeWilGiw
2+NQeGlCemXeNoyOzcgu4Yte/rg4KeuT1T1KSg/MbcH5BcmrCKbu1KumbFWiaXscqmqWdNJxY48m
B9F0Y/fbFkGFN+apOUJLQmsMAWomSkemVdkzWTKpIl2KERTB8ZT3NXLWz373fFT3fT+7JQY0xC3+
D94GAkiLt3Fy36hueuOKFb4yVBMi8DntyQgadXAMOF2bOu1PgDnCSEdplAp+ffCUlCldR1QmFS6K
v32/TDpOC3/BeuTvyXkb3Wi05LJFN9OkPeaGFqb61mK7ZDYCM97Mbcbsd4uRvbVw40lZmQ2cQlfo
meGhejLV9kS1BVyEb8nz92kAUBRayb3nsv+jppk6DOP2URyA579dN5cWzEr2rVBfKVqBYWD4IXH+
yE0sO3RXag2Ha4dSpnYNWqZ/VtxwyNG5K2zMbZdR7aQa0E2PgfLxx4NZMNRRa4fcOIBsCppjgOVw
ub92Ie14YLmSvKAiOO3vuskr6DsgrrqF4ElODVz31tY7tRS7K4iteDmDh2j217C5Wi/AJWwcn/1t
LdGsWtA74MTEfPhqsWGegu6VI7eaFjmzEk4667bzTiLMhq9dvUC79DCIZ6V6sIX/o2Lj6EENual1
ek0/13K8JI0MXRHyJxjJJXYySvVJI2XHBbXsxVSERIvDTB00UNEr/kF3I7Mu4c+ENOEVwFosfdSj
9ekiR5cdiGjslrTbET9QCGRLCVaXvopzicEcQSUDVLPwN2cYo6xjSBL9H/PgbVUjIAaK6nh+/9Ol
9Bwk+o1Ur4VU5eTx6bAXGEjNUsT4e3aepCUB/l+KQfgMIxxz8hNyLj12zoeDii+1YiVqoNXxyTU9
t3PnCX/OidxhBd1NrPIc9D5iYGnDCdODhWPYG3yYYx7DvsWkvTm5JcFDG90k5n6qktpcGVILG10/
Dt14rAULz8O7veyoIBm7QrJb3brdaLAw7Y6EWHQ/ZvlkyecL3NhJ/wZmSMEzYrihii36pSqL+GMd
q+qvRsk1zEdeKBUGXtSdMBX71lc4RhzXMF/OsABYuvqDpVz0hX0s9UXbXlIiTvGzOaHzEsLNxLvV
Y9OUV6mAVQJSnxPAjS2Wpcxza1P6JszzAnYlmQ8Y4a1K49JyCZ9su28EKsSSqTi4oiFjDKzK2Nf7
KUu2/Z3Z4+kJ+rmRWF4JX5fuPzHf7a/NMueXhrHZNof+xZTwJGuZNM9tNbUQTGE+/LX9V2eof58Q
SwxE3attvglaphyu7dbKP8cJxegDNlvSmJ8LBF4yOSe0r8bwfkNVFdIHV6cjT6ig3ol6gabRBLZQ
qLNsQLIg82Z1w2xChu4UotNHY0ewz7x8jOVaxhEt+zDk106tdhHPogxznUEo20TMLv5Stx4M/f+s
KoyTSuzKMixFZdy71xNGz5p5VgJiKlEFj0fJaS0kGII0sgqDPURe5+4kiC1ZDqtrpBr+3NxEHmbr
wCQH1qbV/rHW6kLTO3zLH5eM/3kPWVp7T6jMWpMamzi649ajGMKaHO2rt6IlErSwTICHP3Y0t21+
e+B1wVucBy1OzF0H+PdIzEmqPWZLBltGNyJaxCDSma+H+rFqcepCshy1EhoX7pvA8YmDwAlWLUdo
ELY5gZjnYbGKtE49cLQ2TqDQ215GRDkpOX1ZM/DvrLGxjv0xZeSFDXzRTtlOjg0aRBl/EjK6iFlC
gsC2C5xZPjAkl3B3vJKWnc4O5kb8KGbHGL2Fyi9oOq++YvJw14hkc8of63kJFakXisaVFDVUBiGB
mDdTOSA6r3XE2gDrGWcNNQzQz+Al1A2/dKfcKn3LdHcDCYwTOZ/lDCrBBaObLjEl0L6SkbaEl1EG
WfmPfr0hxsyN8ivFueMQFycN4vqs1xWzw7Za+OZvGd7YMf6dy4d6oXETZJJXsM8NIq/lcwW0jRqb
ypaM5M5dMqKJsjCLIz3cOfoLZ4ER2cgtal7XSjB6W1Ds1bEupv1CTLy9EAtbnIlXRa16Hrn/rYB1
5kOa4/xEYW0USXJpvNiwzp0qtcjdE6ulNSY+yDWkVeqwsvklF2K3G7zCEdqkQErcd3dlB/Ps9oKA
vplQo0tfHA3XwivykVn1WEwfLCOveop9iJ7cBXvthIbiEVikpsH/1o5cKaap/xVk3GJnF7+WLxP6
CKOtGfBK+nfYI6oNgU3g28tFGueEHED+hpR3r5q5F3pTiBP0XB+Hjclj7s3i3nHrQ5FxMfJRoau9
duB8hLivnJ/CrDL9Nc0OtMEr098/65jrRhvSjNNx17FwdeBJYVaShp32UHoQKgh9ds0eGjIkm73s
157BQ+gXXfQN8jjcowzg/EqN8bo7YjgGgJEcsNantOe8sM9DnAhPDg3clvdzQnVnmL34hI1ynkzm
pK5nraiA713aoKxNIK2uh8Vbmtg0Qx8l3ZTwouN14sAQb8ffLWLryfP2FRx/tb2Rd/c2g8uRO6Ug
MnQXzRB8YP4ExAsOpH+5g/ClneJkt8zZhRGu6fgRfQuBMTQV++Yb4J2rY/mjsdYfZBkr8j+3orCj
ohpN0u1PQvv8p8Pp46gXadiZH5DMH6LngkOmzO8hF4St0rZEA8Sy6nsWgvR/0f14ELxnEuyBzmDD
suUHSpQGy3ONrs9dwDa100jXM165fBK5AgU8YuuA5cJLLMGsXuaj3Q4WqsVe5G5CB8fQd1nOtxEJ
qe49x2c0WvOERcEEbUgH+jJioLy/962jkDo3hs1ZpZVr7WGeLjMCN6T3UmmwCGFhZfELUIGd/Dvm
+4Uvi/JpDJaeyT16XvSm73jZwCeyLNz583OwyCJ5fSxKHGRmRmpvitd37BYNXnydR8LWR8NyFlWh
nZuWFCSWXReMGvQ6uJLmvAYrMYwgOIX1SGRpuCx9zcXV42br/1dtw1/I11/yL9oonjS2NdHvUPeQ
2Lxtrotg+yh2cOI5JrJGkViManMGFpX4n53NUP45HfUNlPY2JlgXT2QrMiny/BmrwW48UQlj/lio
//h+dsNUD4mqNfbTKK9XfwSppbr+jDMOx8et3/fJ5TCOYLZSUtJgICKBhFY+0K7eJMHvint+dPD7
2e8lYmLjluCw8LjTrWNW3h2npPCm3V6lvtkFhJcGjNFgVPLGTRSAVbsFvlNVSJf4EsjCuqk7FwhP
WzrYGKMeCOaWP6vbs3TpfJxEd4XgRMkusJmPM32IKdwj0THEIwmbMPJZRDPjFxKXKZMsChy4v72w
BGi9xDCcHqs32oqH/w5sp4muXhC5xT9/wHvlIAuQwV6hYmNRbyJsCjT8J7ojIugzabdGtsWZ6Sfi
L0gEaJh3pTf/0LMeZ1ulhCRUnwyob091akGxKR5iYHm2DbYQ+AvAZvnl9t8JzpzZJkgps3tqZkZX
reaUMPf6IOvY11YJ5CL+efiIaMvlmJmgCbyNHWFq9OnYvUrjPcvFVsrLNmirNgvmbx9tEk/jqjjK
on96G0FDQivwIYtqRCw0Vk/80F3thYKaJeqFuVm0X/6ctNcM+ajMmgxelO754QYLHUiD7bwEQ3nF
ZPQRd0aG/L33cqc8BluoCYqfXsTyqCGpO9YctCaBxwdkPSoRxY9M0/xA4xNGkpnki0TTjjjzxcV0
TtpqF+EVnK9bMn7U7iJSGp52A4X3ZVxKH91pNq1HjLl+YH0hHuFLDzfUYg3JUkuL0qb37P/WSUPE
utPtFULYuOjixBowCP9Kb6goiYWsDlgJXE96SoAUzoB5wrlOmiFVpn0EE53OwLN1N7/aB2LgE8PB
pBfazseAsZpVdHH1cgCgPhUcvEhAycSezmJr5RtvKCfN3vcXjVzdsYYABEMwmCgwfpFN4IzJCXPv
Q6i9V5PQ88lo1wqGzkUci6VF/EAtV/VNzkP3Vf9/fC3E3vWe9ZQaA4xhNJB82tHWEgL8oz105ncm
eiZdmkLGcB8BrBBNtnacNKMDBaBihec1wUC7aIgv1Jn8/kRJemP0toLtEj8rIGaLKSKaMU+Vh9tG
4gQrF0V2cu92teJbxypjUY618kkKrAmnkm6L1Y7Xi7v6VFR3KWPZ7tcq0sKZEiQpjfGz/aoSxnB4
5Q/4b7r5y4wFDf2eN2mOeAUo0WMId6mNlL2vJ89vypArrT/v8LnGd38ef3bFiVG/5nSJ1iRzPZ7A
KCXQOFWqTUK1rRAYKeDRTW8OaUUxS/GTvmIOO1zp9Mig6au9q2wxQGzylnQnNtKjogyj58rR+YMF
gmau3Mz+06O30JgC9MPpxZSRNRPDF8pP0Gt0ZaagKzEn/ivEbonVGp7cz0N2j2U3NLcu073JDalQ
xmqoQdZ5U+305UTbPWmsWQlrd1bJSIy8Yhb8jy9rCmWRg6qwIEkRadPhZLS3agAS7f3U4E8zQE0n
ZeYSCSX0eVXDZWG70TbCxlCwS9jrbBkoazQSf5dGjksFK48N622f9LW3+SfZVDj0b5kif1eSB5a0
MPLnE0bBjZCTjREJ67Up0N3udgMS/DGZrx8mzb1TRxIFSWpzkg52Mb5GNVgHzWcc6zsAvjC46vxe
t4yd76C13GOxV9XlO5UR96BlyZgyqioHhfwEbS4ZRqLqgkDBLimlPSjpaaqAynpj/BrVWRihhAFO
Ck31HeFDtnRwFythMS7D0czKLpY5cwFS6Z+FymbLYGh8zcyQSNUvPr/fA0RxYrPmMPu0SrqWG9md
sRlU4Ceoag6/xbknnWjjfy8v7I7YRyWKL4zqh/0cY+3RNgDq2QIOsxiZZ7yfUchgWN5aipLUG5Vu
AVbXEYsZ9qPsLwdDRtG968zVwDWA96hgBlFaZqfMWaT28Q+fM10a6DXBJowO8WVC2mLO9G81d0JL
t3k6v/QSbplWd2eGkM7CiIEHuUZhkijqPckPoIZs5DU9iXxT54x5fBuLihp/WVwB4I+xzujqrh8T
kVmseKGJePxnTpuFfUYYydyB72i/YWXx02hOTAp/50KKMa/HqVSWOBSYDTgsHjU/WFndblrNIBFQ
Q/rHJtsqkGSMbZ9elpvR1y1IUqBDznbvjPbt6Gn+zkIOVKRUueR0tmpqQKVfuNN3MMIW5gY3G7R5
1qmpr9Knuk0shbHg/hhK2eUIOWytOeYkbgxvphe6rXD7JXq1vddaAlmN8cXcs4oRpam/DniLBqKN
dAo1u/Ir0wi5U0rDvaSuxcuga29Hp8X+0OMsTlb/b+gQ8DedDJUPp43fv9tiTfeVx3kk8hBRdJ8G
2U9W/lN5GlvyHYGa8sz7V1rkviKRW6ST2rFyxR5U16fbtKS6bCWXEXjlWMBTpV4vHZWjnnls5qD9
HC1jbPxXzSe8zNyWsx0e/urgc2guVDLkufv+RZjELDh4OsMQ/r5fu3feJar2m/XVFHMXus9M977s
cmmu98JE6RrPcQ75zkt19ORae2FjpnKu6b1fGBrvn4homZByny+WzlGRNs4S13DRTX4w167cML6w
NPMACU9Y77+szuXHRMC4GEasovfE6sv7/fNxRho7YQftutWpPZbuKQQ2kDglNZNlcBjzgdaIJNtA
l8rA5F2Hr2s9MfyZtflj22kttomdV2EUPI30DgwqS4Rr3mjKBwA9+35cuTnAYP/dPV/0UMxpRolU
LfNflJ9hdrokRTcu0YdvrsBC5nHq9v7AsXPjkBvhSH/WZdjxffy+zuLtBKL6/RCHkCzA5ugz/rTD
CI08e+SQCWQIIW+5V0szRNOncXJbQuDXIT4kIb+Eexge2Bh29re+OFQcHAiSRWm3KOeDonCFseZ1
3/cisGhmlsEnxnYMKNTsyzs1NDk49U5vSvPHW9w42gmetjVUTIPoC43xtLezUdPY63Y8JYBsno+3
mgu6h/8F1e2gHCHQSQEI4h0zbHkscAjSWZIBGmLY9KyTfIgNgoPf88zw8Ehc3w0kyrRxwLu6IR4+
u2aKobMsdxeHuOWaHqZNQpqiRfu3OCtu3fV3V0466HGeFYYHfapH73xf15cxQ/fWKASlZ5nNpidY
Vw9ebfyepPrHo0wyiGLpwktV9PTNo4ha/KUXNP7YthD2B4CM37Xs6i2hKi9M/ofpsoYUOwvsVEwk
mNpdKhQYXjzXtCi35JOpfoYOjfNA5+nw4jzNHcvLFaf6u4/w2ISTEsE1WT65keherK2Qf7HSAJ6V
85Awkkum+MrCKrfLynmXxCyUHGIJfnOvR62BSHWmxjOldDhhbyAZ2JwJSWK5cPQDZuEcBBGJlFls
bavDco23knlcgxH/qRYFnBSfKOFMhcZk2aaP8WOFrJh/BC+Lw3A47Pn/tC9JYZuUHVKRe71/nI+T
wyevUnjl0D8EqzH2dTnM+4SI8lOkIVi4xdZjIVcVovSFFjLsWmmZ07ffz5iTMG0LIkWpN+JM0fEY
NFuoFw1cNsbxBg6TfzrXneSnwYQFLVZ+lpvZsCCfGQXw1BB0CPVKHVI/gCA2TU0Xa3eDqvAqs3SY
r3tm+5fxCd4HyWEnqhEXjiY7sQSK9OqXzzGqs0gtRhpdSnwq+/DjYq64/KoVWyfmUclq1Fko6uq0
kXoBWWbUFi8caRnbIbQ4e7Yyw5RASghEB9fiOyBz373WCkfsmPRFwxewL+KvNFz3L1Xi4Kvk9t21
g9BFAO1hjtTbsV1/hU09E8CBDjBNqDwVhf9VlVxlLWWHdNdYiAvwlMEf1NhiuqsjiqYJDjC45hZ4
+ud8IxbB0TDSEuCppfsoPu9upTM/F0DajOHcMpJpJbhr5Ucl9pmN1IuyEO6ya327dQeL7OHf11GC
b2q10n445eHYuuk0U6JvAVeR/REuiDz7UGFXQt/MFoS85Xmy91hkAhyN7i+X/Ez/PZEmBztP6Ogy
S4omAcQwo3ljVdKzdah7n8xmNkzVRrAVr/hUSxqjzZ+Zt+MkYkoUE98U35WO16NOmph8OsmA8QqM
e979+/P6Ww0d+0ZfPh2NEI2Ht49HPTw5Bz6OnDuhwDyMYfI4uWYnyW/MPko/MXLmpzNR+uNkHx13
/G0+AmpVZETuFoADyzsY4doHVVHNfn1xSPNMOBV1rsJkfWNYonqYQhjUw4MIBMtTWkb+U7U1/gTF
ox06rWUhzLrzI9M7M5vdntabjvQY/dek3O7oQqavEjaUaQFCmK8UIJolYzJAUiyEYlF7z0i5ixLS
oC6fOqjhrqjzBaew/FVc+obHCpmc9xRheZnIlW9x5me5fnDMsNarx4KA15eBKqDEi0RqRRWD3MhM
gxAfTR81Q9MoQvjlBiYhHjeF2klCV+NX+2J64A1ceBpgqffS93VyIapYL2iTKZ3/eGnEe8p5wCDK
wFIHLH2JrVYBzUUwSOkZDOEq1TeSoiG3jXpCXZmSH7+Z2e67tkzPlZjLWcKNbhg5B3ob5Hl64qUm
UIjgDPY5xnvH2idAnIp+poBSzRjur3DJpExLb6s5ulIQmTTTS+LVPq9qMrfnYOZ0725jGdCahcpy
eS5UW+be+N5Vqu4HCxAPXH9PSwD5Y8fzyl5fBK2iPZx+f5KrXG/0yGEe+Ti/PtevplPcUdDoLGQb
/ECC9Qf7Uo1J3eoGLH1M7Ciimzoxs57gIfTrAczem97gFcZ5rPe6g7XSMGFatDBusYeWahyXVvwn
OYT1a5U6LF0pHZPsvrUv2tJrDZaWcHsjhxn0+IfJEWA9A1EDw+1hK8WhpKOW7LA91Owvr8756Er7
yc4SIl7rA0NYv1svvH/DEhp/8zfKdO3RPvzLq/RyxWpmmcBxjKQKrH/454QVvaJZ2qdiwDyPjoZv
2ZvcWkwfdXidmB9kmCMnJTdgzVf125SHU0mnX873FruXpfhl+c5dc9UKObGMwqBiPYNmBvGczwIh
iluIqfnND94DjVHe/FuELC6hR1HqXKZwbmY3J7n8Y0d7LT/vatsGFSCtp0vMA5SN0+ftGw9Bqj01
0YDWMcUZPHv9Q89pBAoALwu3yx7PCKBU6/lqyw8Ikc03VCXtBqCIkIjvAT3vkx5tOSfRZzorNAFh
LlwiM9cXu6iZPriVvQ2sKTnixx8UeKfKxMBOdo8/3suanjRU01SuBTaweLPEU6ihR2eM0om8XLSu
QwGa41zfqAJmE9Cq1mX7W+y9KAX7B1PY4n/UG2jvUwjsWn+qNue9OmrWmdkoXN/LWB9V1Z/EaZko
6VBNkjuwHo+9QywJGQ6OpFkt9LoDP2MQD5lAt7ir5GHUXZ+84qC7QuyT4kRiLdym0RUbE4pNG94P
GHMrySVpT8X1mQBmlW5pKH/XA8CA42aEMubjnw63DoymM5DKlfC34LvUmdWNofmg1z1YSf0oOUp/
hUFmr5HsDC3bKzshIrBhPFDVs6vMaQZyKMtHcIKy86C4vCCytkT9WAQXuPVTLNbjSDNpmHIg9Q8e
lsUtm1F+bg7vWnL299dJGlZAnTSGzcAmYbnDYJNEhXP2Vuy/q+NNzsvmO0GAzX+fvax99Rip3zvB
YtSvYT7cYWYzGzFyrYiyfkqdM1zZVlw9aXSd3By+BLRm+oQWbE1cfh+YM6QC6MuhLr9nqcdf7wDZ
66KYLblBcOpplMQ5cQa5kIWVgTtMOo5mgm+V5m9Bj93sCvNCQ3OxndPCwNjachm3LnwNWjc9sxQz
fuKllXWLyxBXQRqli4Yg+vKSYP3RboZ8AefzyCh33FB1M+4OiLewTqFcmO8rdAeVuVF1kJ6Edwcj
+Cz5pXyI+750+likQ9k95g3aOtDD+1irZhvw9IA+elx4A70ozXHPEs1+m7PzOBwutPpQm649Rls+
xQZNhfk879CMbFeWBt8932nRi5qGcy995KeJVDqRka4pQKebyKDk8DTeAce7qGez8zmzeOVKScI6
cH3Sc3SUo5VhPinPWTg9P8RVSnF/aON8iOIZI8QnlESwxrj4t9utCWbz/cLWQB2OEEKvHq6RhOCe
hfKF7s8MaE450622AI65F6yvdIeMWk4V76HuMoSJq5fSeNoVX9CFWvwM91UxOLbrJAAZqqCcEUpm
s4uX2dHNcG5/uRGlKFJhAuZWyqrSMDDIsQ9ifn0ziGQnquMTm74PX8ZAwDC7UEFhCPmCQx2wvOF2
qh5ApVFWPAuGI89uxngli1fUyMg1ckl4SgCas0XwIb3LDDznmAPOPqNXXIo5pvK3yWjjFqJJz2Ly
YxIBUTmhKCc4TWkbsTvGebeotVvhFOGjld9GJ2NJO+kuJP2kBcAF18m901ErhywTaJ0bcJa78URA
LXmOA8bb5c+/9+0Mjjv4ty6N1LWH7C2wbbZr7LzSw3M0p0zjeY/iihH3laNZfpenN61XOvP1Kv97
mHQn/p20iCQBdAfy1nGPyH30cuF18jh5tM2W21VycF0KmTcx8sCcd8n/x8V21Ht8hocYE5KvTE4k
bkjXg/JduCB7/8KNiOfbXYhJC1+MFDIZbfThGDdUOGbxsGs0op0ktIjJXHyvruBOeN/IgQw/Izfb
HH2+XhUBlYgIWnNF+xP89yXq6w4EzgBGTx36RY6lDT/HY+G5Q0RZKdsHjj/1v10jq57NSQemQcO/
Ff4YHB7cXurTQoGYTPacIXiyj8X9/SARUmJcx8qJew8W9onUlAsvedo3ScSJKzVPloEhwrW4Q2rg
2sQPG816QGfI9Lp+xW+OQnITedgnNOsyxIaoYV1M/5tzJaf5qDJDdN8b3OgdP7VNayIeswUTL1jW
GZzvwiCPhWW9mZQ710yU08LzzJrZf8QdlPUCWzijfVrwQCKBHawB1js24F5c4aByaa+zcYqM2VLN
cF+f2pMcxKCymAdptvaD5i4+VlBXg3xHt1eUGLVRMhtmu/Kb1n0qCNZ4r+biwKQNwlfsN8iAOt1t
IyCn69h9MDPPzQ4J2+qLmPfgNnrbth9DcYa9jeXNhObyRFX16x2hWa/Vb1nV0A5VeIQHRb3q4+er
8hNPaLJNtNm4softk1sgV51NAVtT+j9uJkv9H5GZgBcP9RNAwFrdhh3J+nRXT/R1EGXpLOPSNjcd
RxTOl0UvH+Brll1r5FuOjdgueOXwbeUMVQH/LnejLmy54U9//MBewbdL2q7BEjJOq2fi63YrMIOM
2B6NV7QBnmcewDJl8XhY+enAKburaHsGuYrRbFWnbFfNqQfZcOBxESI7sQV0+IKxVUAgakJPCLPT
QMrXuiQHjs/D5j9dtv7Rvfqjp3oMHpVSbwB8hmg+YnsPAy4OqFJpRLXDF0jQnEXTdoeMcHA74rra
at2IuefZbK+zOXctHzeQyRdlXxgrxOSgdiqdbq9XZKlo+tW1+LOgI1sv9u1ijW9LG6XE27XV7ek+
KuYpIGx3bd4n9EEA3uPQegkZ/dpcjdD/aeuwmjPzL6EF34834cp/EziiNr4EixqyYv03s6kj4LFe
6PCnewpYBqRdNQjgMI4rEjo0QeaO4YdMPoo+dWqEd5EEsLDzBX5d9qWKkH8aoT8ZY8KzKMzE6JPZ
iSzVU4+ezmHauFEngmX7L2yys/2kdizcrfLSg2O7yXMJuN0de46LtyTQPN57goHvXbR8KSm/xjo7
6hLmD7UE4QPegsU89Ogr0mY9I2OiJ5n14zLKIzm4njgbtn4yh/6/EiYBUvqHo+uwnkX43zlMuwir
CajMiTpP5Dqn2GDX5CMb1Bevi20fjA7CVYnPX3MCOdfsEMTF9OLXfpk9WeNsllS6z0gH0rpw5j8F
pgdUWTCWL6ZaYuQpV+GXhUAVcct8S+h4fGW28wv0pSu1ckvfcW/MTy/8vDwrghVCVUREUqe1BnOY
6ei/vPA0eANGO0Uus+j5DVJV/XLp6JRRFoEbpPCVe1cT6bz52fkhEOc6/qNV7Juz652v6lXyd25T
IYvHba1N8A50iPwqDU0UGTAMZd95Psp5Ip0gQMdbppewZFD/VlqhV21yCt1ST0X4XOHJktsUknoP
3LO7T4tsoyvwP4l1X3ami22FEyOpZ6VYX4r7JQcpUhjER2dhVuEvO+qG+vxyoeSU0CxDNhG0PuWA
F8L+NhG0FRU34Ro4llZyaIbzaVHXI0DvL4rhgCkF+NcJ8RtKTiUJ6uCn6f39wWwCGqHWZQgiYD/3
NV3ME90Bi9TIHHIAktDM9BoV/3jtwgl1+8aNYjW/wBlisXyM/yztdAE09X9fwd9N9zwyoeJ/znX2
+1Ty4eBBc57Z3+KsAk9rJ5L2bzCVUtLzrRH6OltQ0J9+QuRETWBgwGQCi9e14OFSmUEE1FsLqKYB
bWfUatcPf3KZuo9FG+UsPb27DWcFNM7lXtS4s5gX8bHJMs+2J2bGoPPkFfeHAo7L3vRdFLZDNX34
aMKocBB5cTUb56PVNTRKwb61Y31oP5GcnxyOHr8mRQ7UINpQXzwu9CMJkHFkBaaiT40po/H2cPI0
5NsoiDotntSlI0C2palJhd9Bp2HBzHgJ/5zuUnHZuKAKpeU4ryKMJsGcYb+5OnWJNwfTcm8y5TOm
NUhbuCekDDgyPg68Nr4rszpu/680PzdBflShghIwbDn5MsSUYwoutb0V5dDjfZmT4KR5KYgjFW8x
mcqNI9BJyvUDcCKUr6TQKxN2T/SFrENhe8nyiNrZzO5y3+FQygbUGGgeeenYSpr8AUPWmo0pvGwm
jzWHsDm/FqtUBm9NILSJRV9KIoNOvA8ocHMsz51nNh2HC15iw0IvlZ8cGj+zCIyTm9i+TA0ajrjd
SHQmUI2QVGPLmSErDG6HSx0+eWB8NZZl2itA/Y5m+yJT4BQEI1mlvv+lu9bbheKjLjaCJvlnXB8T
VXNdv6TdHXB8lVgRbF2qH9FmTMfVmz/TUp3Ht8aGX2kqCWPpXQWsUeQmT27zcGsMi6/qUoogz0i1
EbSrb0Cm76fcDgMNBomMbKTjd0Kj4uBvSCS8Q9qxUhAWBnyK9kG3w2haSCYw3NUeDBb+nQdVrEtT
TGA9w5L0CQmvLtqec3crLkJZfzzZJKyz1ieE/ODyizZRlJVZS1Oy9Sjkr5ONu4GBboFmpMrtla7f
Vnk+tyoxaFZQBmWyvfMNP2C+7tqZtpEAXhCzXyO4kCrMMGS1tJNFu74/30uTp/6y9pN1MMN7M1aT
BVMrwjl49QY/OlJXw1Ure+iJSzLMU1ybH4T+6jSgIrF4hzSfkRWwl2+1RgSaEEwBFNGUY8FUAHPc
ZAsHVTzE+22KbEVPwxq013LOgv6Mvx6lhN44Uvlh2Xkbq0QnEoMaGp5z3COVHMbCt8E9lYoeD+y6
5NzdbTXhbbOIinT/rB8f4boMkk0jEYOU087dPvn+t2mDFOYYS5DkTXRRCZxuEnM1ISDusfgw+VE7
iKZlYksqtu+xOTfzNmz8Vdau95ok4af4Ld6Tc7CVQ1grXcPwvlCEO03wZN+Lzmbd+SnKQqUkQqWi
2ZZ3myioy17IAOlVk0l2Kc9bAZXTnMjkKBz676ZrmtCciCWLCaScXiupycTRlhckTjIIgnWleD/g
Vj8wgh/mueWNejYOlyXpU0Vf0FoyR7faJ5RZEGb75X9ZadSV84WI1YiEgfIM+L2dwCJ02s29Q2k5
seu2w957yad5+NdQPrrN44XBgF/yhJWuMficJ8icfZ5Ks7VLb+xLECUwXGC8nWa1SLLDj67DzK5W
BT6zMrySwWnzYJib1fBGuHoVWGnvSZhTsoV1B5T3kCLG6/Qss2PAKSD8YjgDqbKfEF+56q4E5Ou7
34f/ue9y+Fijlg47M+h5pb87dwA2AV5l/LH+2lm85lyzqFQU5ukxaEbLLZge7BJeCEqxwlZpN3LL
X3Lt1NwAPDhWbEA056YlyLKQ/XkX6OMJg8CfmLZF/YIoKyXgEZkH5ejKnSwcsgS5/It/+vgk0Qes
SQwbT27/Fem2r9PPWPRBmwzlFEbjrH8iWshhQnCDn352YCDd77rnEe1PGSh3nKliWX6lFbtjZuPg
OeapCvmSc/x3GZyJuBYkdfvU5JB+LoUcppKHhVUNmel+vII3ZRcPRZMDZjSgh3O7yraq3J968Qae
nQBdJ96nDiJ5YNRpL1mO9ZAR78ba9zuap3wSlLbiSIDaGV82pYMIJOT4GbXKnwIkgaIBbhicMBI+
lgK5zoK2B82QwTHcDHebRm9hakDbbVfZ21UVnui9yyKnAl0v51GtHcxS94AM0ZZZA9Ob7BlssZ9/
A2cb7lSIfEUBLprT8uYcYhQzVcERaGIyPN0StkRYOf0UtleedBUwGeMsYTLaveFqoZGqEGXhBNC4
bTXPlf5YccrTjKH3RicmPzZ/UL66RmsUD4Vjz7nD9kM/B2e2chb+w/36RZvZiq/UoAd+4rXd1J2P
zbKuFEptE5EKss3N1raAI0zBD0KXKvotBavqdOwxkppe4U3VQsylhZbUObQlXRC+jaJOa/PE3yv6
kSGAFNnOxEydbWzOfZtTik/pw2TD8uPok4ltJo6Q8LoGBe52S5k1NrEy2UJiRQWxsv/QF82T1Y0r
EEVrWa+FEcR/x2QMFnu4R3xl1I5zAGE3J9QAz0Nj4SIFQsv1Yn4vuBa+r3TmjBEeOPskXAAcLZfH
QZx5lK5pP+r7BwgfSBrzixp5v8BiI6haP0a/Z1owzZasDj0UrEGPohh9ZjZViag4pz7JtMuBs9k8
NAZhp8N9pzpw2gf18Spj8nulsUawSItRe7qZ3wUqsrvW5pBfSmEsGA6z7FKUG475DYagSTejCLv+
dyfwD8MSxvZB9Dvs0jULbX/mddHIdT+NAhqHKx1kp6v53/BV5xt2fLkzbWFYnsyDDLIYAgj97XBD
43IIYx9/6nTB0FJXrFFkwLL56u+5+moxbW0afc8Jyqu3HnYqQ6XkTHcwaX8YNkL0pjHZvWgZ7KiT
wxVj/yNJFHPcJRh/d7KmWxtDtPq6+6fy29WKkwlbl9Fugthtw3dOTTGaGSiPxdyZHmJWMpJnFi6p
lcMscgw3/36CXftZAhZQi3wzXF4JQsSJUQudw3GMS+cgOdm9/qJPqZlbcaalxbaSm2V0z1asuAU5
sLZCxSQxHcg8AM89K3hEZ5QVmkSV1ul1Lf4AM5z2UQD/fmlNC1505+0ENIhCm+2kf3J9L7zF0SdJ
eqQix27xpHy+VQv+5qm9+djg+05jtyXuEC/stM0uTi40Cz7P/0oR98MEZzxqEdIITHfgXJQyQvdu
XfQfxwszbGtrcFiiIjSQHAc33nuYavc0UygM1sqkLKRZL9gc3Z63ylM3TgvX9mdwSrmvrPF/VN0M
CzxjOkNXChnYOtHEkIEOKJ+/BMBFlzFhAjzWqb0+9ATpmU9TBKqwLFVdqsq0v2wGgFYJvTDbIF1q
npkNKrDplspo7EJF9ZxhhAa38abHj5nT9VuQ0K3RO5/rWosj7BOQr76Ygye9w1xWbGum/8VTQelJ
QXmOKb58+4M2B6BqkUGekqHZRV6GkUcMHAixT8/rQ0xzYoN2hZmQKdz6kvKBWTCTcTuDVYh+OhIS
LTVbb8V4muuISIuZLV3sa83jG9+a5vpYLE2hTQd5vuOpoIxmfaf+Zuv0MKLVFMtvIssmqfMJhS7X
BlUEE37SAGs/kAuswcSaANkFVBOgzaujwRI/LQHePD1p8CsDVNT13XIIfe4MIH51Ra2VgU68iikC
gJUoPQD8E+rX4ebUni+FBPT7Kn25z3ytdqTCc2xyby5pYSXKl26ZlU64zA6eGSc7+0rdShwSoRrx
Br4wuV/FYr2VDc0fB/bvtcWgBIHS6gpfTp3CSEpixdjRPK0bjn6qQ8z/eJMwdGwSnalTfAyzh/xM
zh65JliI2V6Y6eK92GeW2dYA5liWx4t8IGNzzvW8qj2GyMnek8zpPs7QkVjursoZquMuJg1woXgJ
p/rV4P6TBMFs1RZGpNRlM18TGMjrhua54MZ1pZyM5PlKXre6ujhDRGnFn0Fs23d+zABENuhZY/OY
nr2IKmnnt/XMq4crcEDZD0kA3CZ6VDZmSCkgnnzS1M0VVRRxncIWSHJnMz66rjq9VSe51WP4Ti+z
84oJ3PjgfJ7qvo0C4XV4G1x+g9tOw3CerSY9lz0HYVY6zPRARmsx8PMu1H4hWNSn9YRhgWLJLVkq
1igDhH7CJzHYxINpGQVdiiIK16qf42IDNq0B3/h/Wkt4GyCIhal/8nuJhSmUF4YMKAHGEgYGSrcy
JPJi/8SDGU3CbtU+9gS8r7izot9JgwX3/E1v+/EZdpQK+LtqpEE3+X7poHeBgDAjrXZjaCr5rkXP
30VzfDMqzvG088Obz4HgsagRc4TeP9uPaRK0jALzQcydIHLD5P9SQAy1ltWjzX7ERjqEzRMS/xKe
ZP93gMw3cJOdWr6bX5lCtK5UIgVmEX6ES6e1qO9mYXHkF2B0Opw4OKW/4n2xoT6saugyOtyETmdc
sohTpie/TOCEYF5EoBZaXUom7U4N66dQnnBoEDorNOvJsNEVTcoEmfcfeIXPRFrU77FHKrCWmUHY
9Ai4ZsMHaAlWoxE2YY8hKrkXIEsGUhw2tvCYfgVhurTlLMWPs5c208y+r6PTCb97OdxSyM5VGL+e
J8mVeyePVkw+Uj+Xk67dnMvQEc3b7dd7AgMJpel8oKCaVKA5DXdPmO/0JUsd0/8MrcNr8zWbHh58
vDyzA5G2Wg4qfsrEOsMHR5pdxT+Wg38yRkeQ2sQRzNsrQwzR+l+UdWN3Hi6J+ugmxK8rnZFnRC2C
LajPGwnxh6cOV3ApLAUNfX92NPaWr+TciA5WnyOavqUycRkKWGiGOOWf1BJJfLcERw+Z27eGF1fQ
qqIukaVCGpr4ghBP+FZyevwlUcwNMisfdz6kD6XBYcdsAlKmgvW+c39/qzFTWpfMO1EQ4l/VILTn
QPcdwYCCJdW3g/T/6wETdPNO5NDuqIgdFVEgIRVUjk25b3Rc/ynzS4IlX1f/veIQaW4Sp05LrRLt
wOjDzVA9pdT/gTcuivFdx1QbtyG23Mi7YR6zfNaYaQilLFFcfUbaPHmz3ICwGD8xNOskhwjb026V
TlAi1jb7+vwj4Tj4Rw6OljY2L9fBZLRjxqy/TAG3yrI+dYULkAxmBjwS9/5HIgO5dbSQmJaQpqcR
v92Rhksw1EfIa3FYnjIsGzMhZh70yPXqoClE2mF1IktU+eveWXf5TGcdnv8AIOcE84dLZQ3+tTtR
CXyHAJnCW2ko6Q3bsqszOweZ6gQU1r9amOWCV7suustWit3GkTErz9B8JNdJDqNgzP46vsXSrDHT
62yxEli3/eX/C3ncL+ZrnnXycPYEs78eJm8oJLtaRFXkXox9zvoPU6GCcRcWrD+K/19wXNwAOkk9
M8vCWsDtTC4snn0Z8yXUEBK1lwzpZ0qyZ2u+mzm9rl2SEOEhoaD30jSbTBTRYzaw3Ke+LuMH5e0/
DyCxSx5q0qqrET+NLnWZOqA11b88UjSrd2v0FpNo7VdLgyhumlEq8LqVyPKnNp8iZlWdHkbDV0IE
HRAFszpa6jZh+S4QzNBczUMMAs3ANGPIXKshd7yS+8yHAV0KOf9IpQpznb3FopXHCN4usCkPSL1T
lvaTVLa49qByWr+3y3tn/hCpF/xUZHsPAQHWfOPu2eMAiiV4yvzfAgScuToTD0W2MZ01kyixvIT6
WQQZpztOyBfObhA4PoYP+4CKQeyrysHiQTC4u94GZ1vrSLtLvWXqhadZl/LEWApFHwRyYccblTAa
q73o4xOeR9/HdFzG4YajaI727ANRUlYC5hKpGiYR+nvHqChOgYusRYvPBatrlUHjF/YZydbkZi+m
BMCi3Xku0K+TPf+IPky1FxZeGZf9uJhCs4GTPZ8WYly/sip/PjQoSGX7BY84zOZsSCgBePC1Yt/Y
p0Q7l1LAVtqr7KihK8O3QVek6LTKjMrulOowirTnETukHGhl4QvusGnv4JnLH+o9eQLWPWUlYxLm
hiNwMnOfAkF0Nuns+3QdvdrBRyOf85ZoTWeZ1Jd69vAyBouWC9XYK3j3Ypt2NG8rdRR6GfLx/L4J
om+TRnk5ndhQ9+00AvPrcghKQyv7WFQFTztE1C2c7Uviqlc21lw4VVB1FrjikEC77s5y64iwC7T6
RNE4ZRuK1LKrveGfmJYkKYX3Ky0XQ2EHigI4+58BB4TKq2tcaK9wmAbHaP4Tb/UQB3Y00OWxnXze
C6dBGEsciE0mDr+b2gNEzHrqkis//xwGGJn+ml8I0eyn5Bi/yEp4OGsPpxw/K+QqDtDZVMVxrwLw
gx7hsryC0KsULbNUOFGp7iYk1uvF5VPGuayyov7hzbYmaQT6UjH+WJR2s/gPDdnO/mU5a/S/9pW0
4qkDJyC1cYxHj3olGGYv/jeXDs//Jg1s11htCXasZwX48nFf4M4LRxrTo4TQWGDVCt87ym9Tjss6
OPhJDkwQyK7D+RUWvZRGBtEuIUjc9qdWnJXnJRqzQCP5qaZ61l8eBkgGyfboZZvRyvPFJYOCphI3
0TNXMcQ55H1G70HGKezNxAom2n4SSPvKlry+jXdxx6/isZ71xXUXxaXd8InW71JoOuTiImvWOZSK
GU2PO/QPT3wtdXSPOb6boh3jbgQrfAgc88ez5QY1g6RAE0STqYTuPS0xRIyEwlrgK0xyNmCcdHA1
of8Qx2S/WAm76Xf+Fdi3dAsZfmHe6LOYUHPR7QBXUmEXMXm+WHhmQdhFTXyGNDRAIu7LlArRGXTb
sp+sUJlWcwAuNFUcJBNSnWy91VU7cSQqc+jYO7rX42Xyt9TVp7yq0QhOncHr+q2Ln8gopQFNEaGv
oG+j7hL5jDZ7MHgbwP8d+Ujy5/UXGvoiOii86UmdvYw3voa4ZGyswbV4Zf2ejrOys2T5JXFtFcIz
DCCXSpMpqoTADRHMeMBF1rAOxPt1utrx76dWmlAvbYyNw9GKdtP6NblUQzS3/+cq6O15aSoFYZlY
kxVBtZ306sXuwtB0i2NJQ6wU6CHHdm0/RfLnYM57pFeulxFbhej38hheBaYpPOoBot9BkmgqQmK+
c3hxW9SN5FzocNfUHFVhXPf1nUeSc5Tj5xy3Jf+zYC75pyHpnqUofPRQUkf5Dn/lJ6TQctn4xNDa
cD8EOUx0Ka5rRSqxCG866PNn5f7FLXwk99SdfPzZDCBMcjTRMHKFAARqb26ICAmtUs0WvgRuxae3
5ymT5AZMcaTySfs5Z4f2gpBqSKqtkJRibE3/vvzLxDtDo62Mw5w9vfpcS8Jn4CklzgTepyB3XkSf
fFQok9QY83PZoeHNETuA3V+fkizaBHLwPrFf9GabwdGZsh5Muk0qOeie9S6aCTTAOibU8vD2Vddi
W/GfVKKtIhUaojr/VYN+kphS6oEb34YG1E+Hx9Nu3d6DoGfar2X4LstxtQTycxfKplpVyHfD9nUr
KaB1GRzO5FkWc6YSlOHRulZ1nYhCO3LLQIFGTP5E2obHPLm9xQi/KERyhKwal4Br0TEDesAcj9FO
/RXi76dmxehuR3bZnuIBLmDYKj5/feh18DTyglTUPH2MqZt8+43uaXRd8bZCBqwslz5vKTDkBlpN
Q2yZ2AjN53wmo4aOnzHUej8w/I+Q5XECxjQ2eu0scqwU6p4cCPVRKf4PuEEZOmtyctU6VNeStRYd
HQzSTjxsjIMcNnLQEeA7RKLu8ucM0kRxIPmAQPEKvD2DOstnnCahf87g/E5DrvpPso3YmExsmu+C
iz56Eeq549teYfF1YlShPKiu3GPgA2ZQTnnlYG/u/XXq2uBsHwiZ0HhnlkHN6qNaqse5I38rCxpz
w2m9YsA3Hv+joODHtdfhQhZZSbBPMWVPzurO8LNIa4PsMbVz+nz2Dwr91Uq/8s7E1cDr2mO5CaIa
YfjrY24SXXHG3ZqEsar7oYNMcDofEAnreexzND5gq6dyML7GoNZhFUvfQUCtCDej8s3qhdmZQrOp
rw9oghNHiJcV5iXyDeN9dC8i3Kd5ddiLwJTOmjF8BI2QbY3KBAwWSUFq6kO7gvMG4G5AxLsPNlf7
UvPeISkhnPkd9uVhMj9y7kw4X/gPQd/n/K83DR0tlOdyclcmaNoJlLAYKYSZbaMN1J6jwHK6eroE
kBdH2gSbphne49N5i9aVgRQAoWxHjBWEu8UknVDzz6o2okb8WngFZLYryUS1VsSko5TSvxuvjvSg
KMYtJJZuSKm6VAIONmiQJKjtVgLQSKdBeVbBJ+qqMaajyFsF0ZdRjaAUg4cPpEbf7ss97XijNxr4
Ir9BiWRlwXAwH/n40Hh8iUEZshDHsogDZPrRaZ3Bcy5DpvpCNIpOGSQW8nErnEdjwT7umW7oC/Lp
TsVxdWnhoaLDaSbPMvSOjY0DmXxmdDjiiL9cmWYLeXTS67Ghfp/hlwOHubnNhav5btxHfZZ/aHpH
gtMHFlIpopwYJpMm9ftLkd8WsKrGiU4hEfAWsrBMPQnMI8WlHaPKhwWsuFOoSU82qBC0jdr3kCZU
7KkTNbqlKFJYSCaEPNN7dczryBKsSJdsi6qI41PcE0zKkYkfcvC5xW7rtBPyrq11rXEY74txBTjf
EvpQucj25iBjbKfc0W9SK0X+xoX6Xrrr0naMywI8epL01IS0GJL+ALGkevFIG1H/k3Qbu8VxFZFj
2t6OTZqupIHU1pE3TfWbXBhmGUrZGb/A9aHS3IjoEMX0d48crbgw9+eaISPWluB28g8j6AMigqnI
L887S8zOu49LugfvBZdyXKmTgQGtg+ixmDcI7KY/XZY2ZpoqNNq/qo7T2PUKPrP5zr7U49bTb49Y
tihAaLYPCNO9BfBrg77e10Q0hpEouAfLA5kDcQNVcYstBxR7lA9/qC/BLHrXwxzWZTHFeiimJF2c
LqBOeGS2BUWLzrLrjQaT3HrfbDyfunHgulv+woxvVFbtThi8OurjzSHDhJY1NXRU7BV55iZPaCb2
/3nkhjav9c37KefiK8dUg0RqKTLeDhFtn8esFMIthnI8uSa6NYcUQ7iBRit3NbaiCLZHMKCZYYcE
bc7TXZJqpJNYAjVwnInnl4zPfFW8C2B5lvtS0tnIZVtzQvbiofK8h+B/n8PQmh7+m654j48P/0rM
ZIEbPS3VLuVKRK6j+W2WyumpzGVXigqJQaZ43pz16LiuB4u2aXa/XowKH5Wx01X9E/k1cVLDPTyZ
ri2oqxB83B/fU3k8onfh/YeQgYYgqRXLhZtIEPJ/ASkUaSRXEiWkKknBsQCnu2u6P7sVa2jrtgXj
QS6mvyGes+iYuXFZs/PTfoqRpk38ZeyxGjmfeLAXT+n7kXtyw328uyNIDFIOLQZSZdGA2TlxTq2g
wK49aMwBZ2oG5KpTH5GbB/ucq9FvVs+3PrFoNBGZ3W3Up/ViAqWRo8FDlh295mQvy+ejoqEElsU4
7LTiEUwoP47q9/Q3y/ERfu0790J1waBeB5wduOf8n+MLK4I2Et1i2P2YNeDLzCa3XACemDZuEc55
sw7iX5m6YWniM+jicEfNvN1cEMqqigFPYh06pTLPnjzi80RZXULNDuXz05KpOb4iaPRGSVTgEEX2
FoGFZrADmNb8GFDIujCsw4ZH1ixx/hcIVfyVfDbWlqcK9pjP3rIQSAizmypdfjHSUNtOKJjkvIFR
ITKsIyOwCKzDALlkclzpmfAw0PLgDrNUptt6X3eNqqDYZVyCy4cYvOelklk6kLkwKrsInCG4RIve
YKTNlU9fi3w77bBkCNCBth1aifqLRHtlgcYH7DicRhOAqAd0VXyQL1VPbSGVAM44zuvK8Kl3w4E+
MsrmI9HQUBahVHxXvDSiicWBN48H0cqpZ6CBc8piVwbWp5Pzv+sDilOBbZFwHG7XoeOEo8W3+ser
GLp+9Kzydw67u3679uFmmPiUuv33fZ0zDzRwf9yIfcGBJlmXhqv5RUk3oHL0TsgTwzC04t+X977O
W10WRc0DHJo1YU+4K/e6F49sYChyfp9wK2tWcM9EtLm95ahZtyXXwmDfbFmKHBh4JS+6tvzFcTUc
gSnPzEByx6YTDu1Xg7WPCGEDM6lscvl++lkuNiU5a1YjmXMPLn17Sz20ykv/iaaoXLxTh8nJx/jK
xxvXgsy88u2tCpqVw+uvwstykZG/fhx0UjfNh8E/FKP0aiw/RjRokTdpLVuzVAwiFpVX2pvbd5Lc
oln2V3iM4BWDc7uaMAtOW6Z6jfvE0QEo2BcSp94Frr5+7bGg8An6GroVmiZW+LalJsB7ZbYkuN85
2yDubU6gQHra4CZNqEeQuoNh1bFJy/+CgDTbg0cpJAkAd8K3BZH9U81M23ePd2mPGcp9YpwLHYZ5
8qWDQPi7pdZ4RBhhjGezZl88efSAClhe7EK8SsPLizm5jX3UaKaP4DFhr+JGbOzorb7qj3Skz+2q
d+k8OPx8dq4d7zNqNbPuDb27uSJt9Sbsg1wbinM5hXP+TK8gVpaO+7Qf8rOo/gYc57vbpKy1Msgb
HyDeqJJJOggvxVHFukSnFamZenlA6PzcNzKBvLGwW3nD/MLLaFDnJojM8DFO/++juM2bndXvGcHe
C9jqArkUrsZ4kzEPVLEbqH6p7BcrekxP0WV8R7ESEESKqEQCyIAJ3VKmSWuJS3XiWmE4m3FCGOCm
uifrXTX8h7Esn1QtwJQ7vN2MrBIhFsK7Z0nANxGHqpLOLmgsrxfw+OdCnuUhfQXIc4Vi1KHP5Ox+
XW07zQhIW7SFgZWQ76xHoHdSvj0IZLRs3klgWjGa8LnSbMpaRv1c9XE5u43Op2Gq4OnMyYsSWMB/
91lO3oKA5RDugfvENI8jXYXLHX0/zWH/L/+jL6JhGWv8HX/IcC8Spngk5ZVndueLW7hmcjEW0Vl2
ZPnGyCx+d25axOnq9e+uxSJNVEvavk5LzHBGBDmaMNQWvwOVV+j4AEk7H3kHzbvWCMuPiHTndSym
jHCqw1NBTZN0Ud+3IiGf+wT0zYZU9dawTulBTI7cErdtFEdx8fV+rOb5ZUsN99+3b9HQ1YoUPtvC
eiL6LUsR951kcUUrx8UnGx9l5+svkDPUzYiHs1oKnLm2Uwzd4Fq2G9pak3kR/Cj4Quxy0mlaiwuR
UVVioNPFA7uGTIwWnnOsPakbyW44/Su8Oe40KW3ufqZqEXKkYle1gsGLCwr+67Mhey71MkRq3Lcv
tanOQxDgxCGFOsCz6oFalU+X9/ctf7qXaRf6g1RZUm8BsiIXADncSbm2aR0YBoIqYQGus40IZQYH
i0juu5syjjCBN4WN3MARHQJZFN3sf2WNHIiP3WoFh5dgH3RSBUPbIp+cOixUITlwUwlggJrN4/6D
VU5Xo2N7XuI3p3gu3ntOJ946qEEnpl0ucwSComH10431AXRPjqP/qIa1/bIOg46C2yJWk0FyPdVB
M4AvZpra4SYStsjb/KRH+mk3pUgUUOUbF7JM1wYzdb7F1BslRJlBuDLb2snNuiyTROGbU+oPH/g1
yif52Ua1gpSQOFc8UsUIh9dnQ1Iwg7iNJ/mcs9Ex4oIKLme4C8Dlca0OZFoalMhlHwZe4OWdVMdI
5qzSGKyv1NQD3hu0NZ/hxzzMYTUgHpwcGE9Mw8Ej5JvyNowNfWBqYR3lRbGLINtuqG4lKGm0FDpo
4ymtQQ+wo+Lo7+0MQpaoAsgyAD4DZtfT3g0r5Kh0Wx8zBwjyI7ePV9igy8B+JJAarL/srvxqRW2R
Y6QqoaBeUSaRi869oK330+E9OHaCcqWPXgIzPNkp9GtiQRxu2SHpJ2W0LetavsoN1aZK9L1LH/V3
RvINXdDFN2pIKTXTt7Xe/Uh/i6+sOks6fxLsHX5KyEmjPLVHtRz0MDOKlolA5PYf0up2CKdO78sz
m1dHMCFTmARarx3KGUKTo9ihSG4tcZZdE4Ouyy3R66LliD4ea9G1VhqYIKEpZZPVYtXCUOpOxw9g
qaD2FspyxtWyZvAdXivU0MwTMSSzFewmibYWpCE5Q/sW2Xwt/I4nZFGg0PS1goxwb3vBu3Y57Bqe
AeWptfkgnXFCqhar23ZVJ3jqseCMbyA9OnuzARq7NBZ3fzfX0M6DprfTF3b9HbD8KIA2X3u4mpwi
Ffya+2g3ojW9NgfMLDDHOsUPkxGbUknPnUefjdw6LIveDLZXWz6JbT0bhcjT2MZmO3Uytu8581TQ
PDaQGFJAXviU/l+jv5rDHKPtfxcQqK8lkaSiQiF/DEpJBdt+OcJniPeQvhlTbj++JEyhNz0qJWDX
jwBqVOY4JOmSi9NmEHUsnw5hdaWDtlcjgul1+v9hLBKrvRHoQe1sDdZFKMu+NY91LHr0bAa2x04q
Wd/p+/g9NJw8S1IpeZ+U79ug/1//qI7YGolYEJtlSKfn2GftcxGVUtrRBLyo6ZLGrLit9LX8SJZK
8D0BW9VoCqVw1nrGa2VqwbZNYz6wr+6Z90jnCgF0q3bP+qzIYS+PK449yDEAS13dhT7ep8zC6phM
KnxKNeKDbabO3C9IJv+sSZ1IhHM+iQdjEhukofcJdNZy8Z1LS9PgTsuFZSEOCv+edeRue9SJ64Qd
j5219ZhSlac0ogbtZhR8+03CrPmYIbi4L5fktYgvTKDVm65FMuAVxPeBhxFHh77VpUzhG5+nIE4+
MKwi4GvInRehwYqzI+N44CL0TPlVxL5+5WzFf/JyIp32nG6dBWYkHFeQoYn+xnnifkw7FTH+O4ge
WtYohiKDByecFgUUwtTT7VJXTg2KyfJWK4zFTx/b8VHHLnvgyYv/ZUypP1nbj/RK2yWJZ81GZyUE
Xxdbsv8IoVH3aqQcBFoI3MnlSoEiqwjCWEayLjlIAx63sOYn0tNv8Lo8F2ORTIPMtVom0IGYTvq7
whh6XrCTCtgeMhXamYXJQhtyt79jffPNsPmLe67jpX5a2MFchPgBRSNF07zNDMosu13ka60MBRUg
qqudomhvDOjPHxTEf9jbBD8ermuYIp6CYcFCt2XRz7MgVf6XcoTKcOVit0NwYaR1uALMKrPQFWQx
xiilRU6r3nILp41QqHTTZn7701ttgcCFK690f17Whe93QOX/FQxEoIllACYInTwU+HzOk5NJVIAm
oD7zt639YtY6ZXvXhVwBpvWSAS7a4UFRAkZLx6voV3fpMYAFpuu0DsyCdJPzpbRU1blNbGYugNfQ
dCFhZGslVDnryP5iPKDCpcSWJQPWlesjLV3YtxtAfuyzkDDOoTRc2bOkvBtCDKkhATtaBt3wRC6G
XfyfEsYEee+omjwhK+TxL7WYhlvhroeANtjD0g7+WmNFfLdQc9pBmEtxP2EKcNipibIBbcNNVsO/
cC9OlU2QddZVF3Dmhl8VigomD8kpmkxhu9puO5H+H4YwOGis7PyF+liDS+AYKMxfK836a+Z7y4TJ
Gz5SIrt5GFQqVRmNPxRof2UQs2hgLNBuAyEQ78TcqvpJatVWEghcIhqWxJYnzvGs3VnDGvO4IOps
7q93HZAmllodUdooMcVX1R9SpOOjAH9NFOpFU882zBd0n2Uy+xCOFzaVl3ggxrMJCQAw79xSk1Y9
JxMy2rol1ICkz295O3s3YgRvLCEpM4nonK8sxQLSFZjsKAt+Aathrrr6bprDoZs/BRV3Dj5EIERf
q0AwNrezM9VIVSsOKUnyZofE0vv9BCF+NYo0Mwh3osWAlbgHYnsqiNL0k9Hh6tIWBY7yLDBLSvW1
sVmkMPhrj/1KGWmBtCiqP0V2yoRRTJDlxUD5GVFtbRil1GsUTVmG40kQ9ZFHOmyMikyGCPz0FoDO
66vPT9AbVmbXuIgjR7NPb13zkmj3DnOzznslWxv1mxTLfYFibJ1REfpOK4lDzH7zpugZy9fFEflB
jc7RsAFOkhJJ4UJK5NYTKk9Ze+jtshXXUKflEF1x1Xu02/JaokrZuVnZK6UzclelWPHbcVmXSvVQ
UEdBYjm6Gm99Q9gKJ0y5Z1b20ZZ9A/MoytLEumwqML4iTEZhf73CaDrYCrIkJGZ8Qnq9hhbqYdAy
SaICQfl0Z99Di1s6z4ApVL8hpmZZHgHle7p+l4wDCaTExOEcgjU/iHRYA6VXgp0l2xnLbsW8h9dR
FcROodKUIUYhrxI/m+56GMashc0masvmPSSXWZuqYtwndHSu3H8r1I5q0IZsu4l+FjLMFm6TP8ei
dIDvNXwUtBFYBGT2Au4OGI8sw+q+CZ3R64xJf0MwNbqv8TGTm+HObmwqkRaiy6LUtxBBz9cKnRYL
/24aWyS62HP6N4XSOkk5FLSEnGWdcfPn3KDNpWDC/DWAvZ8TaCBi2Pi5RW1YMG4KhH9Lu2Y0wHPA
U3NcxAjDBf7qmKGXiFnJnOIRwIs3wmn/e81r/ZNjuu/GjYkEkzzrWf3CBzrEp+hdXW6DR6pRp0xC
87rF0L9Z6Ff0ObTSNwoavibx+EoV3vA/2ARVcNG+7RY8PdPdlCOkgIVixRr/fq4lAGiQWXv+9Onr
X+37nkPiRHkvxtl0kyiwiKxz+9z8BwaqT1+7qYHnSf2tNboMgO2XSxY4rcqK/Mc2HkcDWZ93s6pz
0PaQQboFEec5z2WezusU2bXvoVAdSDBUqY2oZ8aO4LyKaQYTr5HEJFgOITB/FbeLuk7e/sI5hv24
JpB0cItiOdQ1Ryd1t2OP+RlhI1titISL8ZNmShdqerIpRaIfowpnrDq/GwhbHFv856VL6w0s2ZVr
i07ZyKaA3sz2bZE6HTTfJNvG5j2+wHU4qaghnsrhPkqR/w3xya2Hh/2+cjRIVnnFzUUmI55Uf+uT
ASKbkET4vWa2do7Fj3zbf55oJT6TIRQrSdw7LBwPL8TF8E57/zlrNKm1aN/RT1y4fbFA7UMfemGa
GumppK8CfDcYoZ9YmryOjZoTBWSK6/tvhO0UHxhAdk9Tkki08OSmx5FSta2n3aqDpJ+355Ufp2ON
7UpYsQr5q1qaj48iYZLapEUIkCIIFYjnxy4793y9CwTRKqarIdDL2pHyTeVdWEvjofwWR6rhc6CB
MDh03IKHAhWZWcAMQ08o16cZ7zG+XYymP/zIjqKY61mMbfEU2nYhqI6fOjIS4ifsPxEno438ZJYP
nBw5TQ+sIW43WW/HzkRPW6SKvPU+Wb/yVJdeXOClSTgAa5sSYPY7NRMxfLvxOqYW46HM19NLclg8
c4CMKO20lsC68dA9YP/I4foeqWGhFOtMtFxkiLAq/OMKvuG2z8Woav4VVPeVYWcja9CTQe9SQgWw
xQFDVqYhKOB3L8lwlpEaArH0HJxkGH+G/ZUfxqUMz1gO7ISQzAhh/HIE7WmmpNxIAp04dzqmQ5bz
nSOQXCeSKoC/QgKFvPqOGgwgUTXy8yggy8DAJ/dOEQzNmn1w5mYHN0B6gF++RKB5JXPnBEdqJWt0
L606IpNa9fiNjXsK2GA8iqNZP5GHl3mdEN4VcFEVxfLPpNw1wyR2gnaosREJ0u3B1saz3QXqi+2M
P0DPdiNTBauaXuioQzupAbSEbeVDR9DHwj1jUTsJrymI21tfFvLxmT8PcZ5GFO60bpJaNAKa9khy
gkgbD7RNgXb69UNwqoF31rToUQOqmN12UyalidhZcuHI0XlfXPUsEbKlWzsfnlTGU3gyGz5LdMc2
E+YjMl4PhGEXv9Pr68UUpdZhltAVdZJMw02tk3aHd8xM/V+amTFb5lYrQTyZphebrk3xiy7d+0CR
SxEWM15PDyLLwVfmp0kkLadnp+GWkScCrdnsza/Rb2Q3sh1t7Qqw/68Wdje0ZmYnCqriBk/Iyki2
1XRyKgvsqGMSboMAvgsH7/2F+hl9qC1CkXKObRCziF9wMML6ObYtr6Z6W5j7/j22x7kfgjHfD2TV
lGHAakH4ZYTlU/W0/YpDq31bv5xmUvBryLjyD6Mq9/yXS92xSxX8ccaNHwW4j1uIuK/qklcw1uJU
0axHZe7g51RxkjqpQCSD2AydA1uTdQOWFRwE2v5QhdJB1h28jHnW5uspyEzEnyc79iGXJuLR4M4e
H8AonE1TYYJAnCdSqVFfIrH1hq5XW1ZoBIPqwziK3aye+xCz/sbPLpUfbrPul3HJ38Fj17Uwbisn
CH+bXdXRLxExrAgKj4jprIg5R2DqTZzyr5MgE93+lkuOmE3fhRtuSR6zfyP60MDa221byp8bn8ys
J9KkK4QjtJS9oSiXPhzADto6lix3TtOOQWPUkjdBCzQcHdmnz1KSW15BWn7Tj4k8MsyaE9eoMjqK
Xizq2Az6AluUiXBaUkqbXJ2YICkI6zjymRiNV4D0YJaEILqEXoi/WoGfsKCWqwPzeFeSlqr4AC1h
UVY4oJbYY0Htc511x/PpF50MUTulv+sQHoBbg5hZnv9dNz/zQkzE9k3m+uGeH3iDI6ER0d08irLK
qUvSIV3QyKBJsh10PMtTJl0PmW5qFzLEAJS3a4ye73eClne94PUvWD/DDHS+Ba7dt09aWFwQcjhZ
x8ytzRUcOzZVo2TOjIrKtrEAMpzg/gw7h3dofH0qDLlqdSIcPI8gQ6qPxfz4mJ5kG21obVxL0T9b
aES7UzqAUqU8zsNWIFUaAuVcXlEig8eKTm+U9HniIKTuCgc7pK9IQmzHph331ORgvu+APkk4kDn3
l5pUk/AlawUCg0PUucgxskSlpRjw8Dmum3Gc7mD9iLUtzL92yfpAL8mLVQtu6YD1gK+t4PJ+aCMh
kDnm3dmL35w3+i+egP8LwVLmct8lZhGDJeOj0jkBSScvkckggZcmZKJ6dn1DnbNbVLLEjrzIaswr
yCT56OhC7OTml2R0z2LYpA0oGPCc7QjoYAKekTRIfKitESgGZnUuL0aFHHN3g60s7qPbrqwrbEXa
rXCQ5JBezPD6PiwQyjo420nrRyHas9JDKjsxgXJbtKwVVxVGGyRWQMotcVM3/ZPcp0I5Kx+eZMld
X2J4pZWZBiEGs+JymM2UoeI//AAoVRpajsxqeQl1ReC8upxccpPFD6BnLzG/qQtNqm9XQH/xkO4h
8x/vzJQocS3mGLZhssR1sWj5n2Ow1Y8sMbGT0REyBoAUno/YZC1wG3BnkVU4QZ+mDaOvgvMS83SV
K+UBsm8bqT0xbPrJG86YvAkY68AwCPnn3vhg1Lm9exLg5SyfUOI6Tmb4s0Z4fQCY0oZ4+Ab6QQIp
i1sKvh4mhxk3ZaX0CQYt7fcnvOiTxSMHwNEgLuN+wfgEDYAicO1wdTozqIEaqhgb1BFAcUNTTGlJ
FLMfg3PxnvbdFfx/rTlJ06EnfXDr+4YYyy3tuk6oD4RMClmqQr6mwoWOlGBlny9hcKE5IGYPRT2W
SQ9CJdiYCBhTSCkU4ARw8MFA+wZ+dRtcYXZUuTwEwWDKBejDVFmHJGnkKjUZeOfIvDRPGJ8YqPtq
dkJqd8kwzw5JWu+2U5Ow8/7suawNgR4d4G0lVFGNy7h00NuKSW1CGR8NxZTzVwVLJTlN8XcABfib
2fQuzk4YIKWR/pzEzh7XwPEOUffg+qCILwOwKcpYTnJZ9HA2hSSj0GuXNWre6vLktnmTH1jS6/dU
xy8OOXK4g0XBHGvI3ioyYWJ56c3ka5Cpx9nlysYqjwjErRLErQrcL6L55WGE/0Lp4hAoNB1Xlezi
ZSKriPbdfQhk5pIIFn2PfBjevNnTGbHa+HoKaw3r2LxaRm64P7VLfD94BhocGPiLPNTAhMkxYd60
tWe6RC0m3aiNguMgz4/ru1cEMWmkjkv/OWbbGsY+POjzFmnQyKYxAkV17jq5mFZv/8ZX0hYgocMY
ESDjoKvmZY5vh40U6qhuC85iGxaVVLzEyU/ZUvR4tIU5R6oTqzsDsnkU/yPxGX69DmLLJq/obopk
vPEa58pFWEMmz3peeoyOckru0KVOOD2m+edx84fAaPQp81EmRYDEyLoyDKDn48BKCVqzvxjffxHM
XqRZNi8Sg2nQPiIAMAntimhbTkDmeiXkDxJ3tH0iM/Vl4jYfx2JTVLsEoyYwfrdR2k9a3E0+okpm
tXr1aB5HJAx4rIa0Jcym6azh834Ldsya/b/qeV0FSI+yxwmX//Hv19UEdpMNEoL7aA2iCnOz7QWS
yR6OJ+7esTkePMVUNt6N/JD0zbkOyi29i1SdVTQ6qfhi3COOtfTfOkVAz5lLh+/2Qx9tie6AFJtF
EEN4t+lvx1TimIxg20pbqNouSbvRTfSRulHUxVfzZEKJMTrApn3/CEqr+j7jikrvgmuAcmTvHeGQ
9Lu0/+WiuxDdDVVOxABufCzholkHrJWbMEVcgUyatAz8wUADcC/sSLfcTs/6fgBfeSuB/CeT/oZA
cQ01fw9MLy225ElsdIaxIyW2mTFA8ttdtuFUYHCKTfm1VVVkIvVqpLyqyi02LxONE+WJCSBOeFDp
MvNMvzSb8Uzc4t23SfTPPn8UMs8DLBNvOjVUULOSS4/755AiVp25qcn9ZPBLzPMpKXHVZaeD7PGD
OwrEqZsoWL/7QV6FJRFZMuccPMmYR0wUbFFnu6IyGPaDzSAINow96l1qRqSMicYMuXuZjKdW7qzT
uBa8Ey0+1fSJ5BleKXVxaIOwOHCBbBE47lLqZYSB9iDk+LBD1PmrGtz9SNPKQU9RjilJmOJ/0DLH
Mfdq5aMKu5xuhyhErYZQKW+snX3S9dYqyRLWJPIxjNdPu47vBRUYUBmBIJyuz6jdAB0L90AaZjHq
dRtJYw2nB3UpyLpwrEI5kMCXTpMdvMwEnIzAsy8Py33trzUsAxZX3yETGeBf2oyg0n+Eg0Jd34QZ
NZ3Lr9C8BuVz1iaX3t9x3qhuggqc3OI+2gIo3ar8wU0mCMsPcJv+BM9gAHgnqEWlf7h23CbkOu0q
cBjKmaJMdAi1RCYzpLBvQfCJOK6jI11LHJ3EIKEo8pN4F7MLd1M0UzzYOPg81lXtOlF4sztUyBTW
XXFU45NGiQC3rVkh+kRqVKimmVNnGtN0RruH5oEX2i21rGB+mx9sHSOQ+wCurBUFQDBwWFHhLaHe
VilAVFTUrTsyJd6DWV/eXvy3/Mi9z1qO0wsZbKatPYGm/se+SxVBzN+CdMi09LSc12+AoX67Gty/
e5guJmS0NSPwh9ADr0OWvQVKXO2FFvq9P/0uEGgVgcWf1TBZPReitpK1H5+2474xoxdyLQITultW
88DrxiRgTcsdroRPwvTLZkYjDozWsn/ug/QikeAOz/j+R6sXB/l3jjQamamIARa0NvxxC7Bk63aP
tuKVKwEx6lArGpvsh1aNfN4/c4kKXhF/FVdfpY6crx4ATMMRz5uuowJHNfR7DDlnlH1IxqHg8SXb
RyvxNNtDyvpTUQPJeUyWjSMg3PQpT+7hUwA9Vu/4aTtJmYLewVO4QPkLxfb/djZofjlIuEZp0jHT
9AIKaWU2avWVbJlkGt/nYjK3JK9fOodLWYAHAMTmPJwzMp80eAcrbv01ZZlEdc/uAY83guBjK75J
6XRElYBCddqQIXbxDVnsDdem5B6R4s89tEXRCWH6v7aFTMkfvOfhE5dg/0uYAlugfxwSGzRzxWBC
1mvkXCX6lcTvLq8TCzaxwk8Te7weBR7zR12zjA8f0h5e5aX2meH1SR2Oc7z54nqwvXvTqSXiU+33
QEiGt9clUr0BYYsJTqiBnpYNrDN1p24F6cyPNSjQFOzvY4fimN6RrINqsEqMSM8ArapLhbNPazRq
S8iBUA6U+TQf3dVUdcNLHDpiatY3flfDyKnTGnrbVF9Wo/9JBlXrO4DWVG1XzWJp8zgqqtw86m1k
W4G3H9sCVLkMkZTe1tqpGgqVfb3uwLmohEXKW7HSDtZApu1TM95sWVbodSMUHI1nrcRut+iie073
pL/fLlYltiGcZU9SfU4Y4HqIftOf760iauqXO5zqR38t8VYP3U8kuIozQCzayH5Lplb8r1fieI9p
dL7syeLT3sGXQdMCdKhmZIYbo41zkfp8oBXnKqD1PtaKHV5lEzxb1fHovRTXy0nWAxSS0ULSvZv8
xMSe0wACmnc1nZQq4aEqqFOWUwc2vAUgBgRKylVIgpXvZkejFnqYJ9COaQsRotF2PxaE1r3b4IDl
zhywf2tFVLsLmvdevPgxiL9wVtnJLlsQzmDQdFM2+86X2B3fK1Ux+XRjpKeZAIoZfrnMywwF0W+4
ed3VWq4ZYT0qnIubqnVp9Ay0EIBYrufylxY6JfcqsRYV9Bx21vIVS50xJI8PmoVOhPJfPFABITBr
Ec6SbXIkflCKp8cfLv8ZWu3odyij5m+iPVosrToCpkKHHZEvfppX5JfFYKInU6DGIkstqPeWifeL
OPCRlCrlJe1kkxpVfY8Jj5EuNksDTQSTHXCU9OjTLg7pfSLHXfPY1u2jPRlKiHuTRWT8pvuf5RjH
G5DmmwbrflK72PZIXi8ihQTE2hRt0hfZW5HlMuVOp/dowzJLzuirtaUpYnmRLkMVf8HaZ+jECQlN
LJQaii1vOZ/AWBKqgq1Syj7DafygO7BfwDrx6Q88djnx4CIjy744TGgSczTTezgbQToUzKDWLG3L
Dylp1mRjgdrjqEb7YAiCQdJgRnaYhYMXataux9XewfubQygQglwh+YylPU0C2wr9DLmqVpwKqafO
Ccup78Q1EULZms4/SJzpwVCeI6TuOJT1W0nDoToOGDuL63B+kl00K1IxYbxYpTBlAP7LQcxoxfAM
afIj0IFWm2mSyEAihlQB4AfXWJPN/yG16ZDd31LhKcFN4golN2dG2vxqrkGdG8IdhfoX5ZChTm7Q
rnrJvBhRtcGoah0StINxAhXIZXCK2uVOyplSQt7mcDeB7zpem+Be8FcaA/5vqcasB9rHbM8ZsU3V
4En+Be9UXxF7jgfZs5HSBHUwkJFHcMxhwTE5QoR6BiVjyEd4y5fjDBe4m6RFAtEM2QEW5bjV4MND
tSILEciJGbMCN3o1rkLvDpRVwqT4qvmbJjhUNxp+Ch0nH0l3PnnrFfuZ7+gFpqendorVxFadwlmP
HySsomiLTEO/K2+AkG3NnoIkD6Im4Lb48SMx4mpZgVi5TLa1TmCivOhPhw+DzldJkm+B5X8D+MuT
ggSi0wqvuylFIozvUssnQvicpfNgGqekfictDVjf6TrKL28PSIYqZ5eprWWrkAOiwVl7MR5J0uyM
NBpQ4J5gZ3RvGy5WSVuuPP8mn0OgrfnlsVplyv+lHcPouf4/qZgPtgDWdbKyn4Biw8UBeaivJcCR
BTVnFhrBYJQEudq6ponxkBPenLkEwjGpp43xrsivsNwIhiGV3jXg7D2exjynXqJr+Dc4OYu0/dKZ
kwEvuFwGyfwXKbClOoDYP5I1Et6oDL/q/X147zuqBzt3Lr5/gBk0wZ84l7Dk4MuZQvs1yMft0Fgl
UT0MwFgsiiUCl8ollHD2UABgL//YcsSqY2CwLG24fwk=
`protect end_protected

