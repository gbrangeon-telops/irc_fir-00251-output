

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jjl8vAn2UJruW+pwbvMAIo6yT6bQgTl9+ZqbT+VaAP/dcMa9HxI5w52bG1uOMJkKjbI3shaTb5QH
+WA4TEmwBA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jY7USlQiP9PR+LALAEYZsrKak9VnF4tfhT9SQb5jLUPXs+eC5ZbIVQkPjdV+4wzhB7b7ai6shnHa
gEu6kUZZsMTRIotEQn7SVZESTAIMCGAU4lDLU7RT30ySc+gN3y2heOoScYVxVF3kYNcbErB9g4iU
iZLVkq3ZU0fP1VLA30w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W97r968B0QPwlTs1emSg8mtee0qHNpQ+/n5wfXS0R66Akqy90VsNXhnqLJjbnGJNqaGSMTKCRNVS
ox1Z0rkuemlJn0dMgZtmRgHM/NeyMTSbsBwVvTSeFdA56k6PzciIIQ1S8150Bxbexnd+b7l/UMK+
JO8+KzzHPEIPqou3srZGn9dog9HSSfTUIqvBgloCeGmDxxwlsFwQ2VsrffuE8mB5Kk9lHG/A3rMw
tbJURgYaS/b69KLL9Kc/urEgbRWHU1HQCQDL4hSKE79WXE68MZJ00kcWMfNfAOR1zytQecSerjXJ
iVVvnEzEtzUejpnuhHCRhS+b62dMTzf5a1Q4Dw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l6IXa1kcvqxcIuqXI9bELoLDvGs5XxFfhbXxOKBitloxuDBS5IYgW7AXksTedGB5rM+6jbAr+PVa
4ykVDtx+9n1RZQ3HKQZNsRywuW0+Fcm/MhmC5isxnEClP56JmzAEyD9l7nmy9JJJI11qQTy86iSs
hkUJMmO3Ph4Kz8ptLn0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gEbAM0PoYz0kTXyuDtZRhRtQJeO0ezbVNuHzWd2Q6Djxe3WZnx453sNsfBBqykQPTu/zHrWi/wfe
VIPTt4c20XjDHHTidMXhf5YGMYpytIjNmzV4g6PhJehJgJTQj+T/bAmaDaXLcqMDTjUNont0w58X
XTjVYtxQgjqcVftNf5PS5GCVpRxSTsKbT4CfmHhBwwsNC5rLtE2tRCpmB6tKw/7xf8VLLD8a23zt
cVvVNX0bw3bWCGFmWZjC/1fhYI19WFrjQO9Y/0zq8T/b6JCoxXV2HE4Z2dJ8uXvV5GV8EStC7VCB
DhBS/R4IfNLPojIIJPxvrbzkKlmuEkhgwflRRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57936)
`protect data_block
KM/3az2YSO1j3vwp4PYLI9/L0KLGhTXLrq4SqzDTpVUl7TPDh15htdrLBKwjNp/bsvIgLN4dMLh1
8fAGDqv608Lixa1cl5vCaAGiDgCve86r5b7inR5RB7hoEiD1VQF+uDaq2agad4tLuhafuFTjQafm
0DYmCC66k++IsnTiXTy5rc9csiKbHUr8p9t8VRcq8xGGxTJOfkdHbxkV8uejKe3aOyB3sdI0umXH
UsguAfQ39t9cw5LTETnKuQLSGGeE68+l8aCl3Fz80oKUSnzrgw973b2v1tc04Yax6rImGSvCdx13
64rRNcQTJepwhBW/+tKOv8SjunlKHxhBq5BPLgAMHBVA7clIMYX+qDUwztqJes131WYcGZ4KGnp3
rnP93dilhMEnc+yhzH4a25fgZI0Nk93dWcXRumgUq1b6YgbWTLT+RyDUEhdOis1Kg+aJltHrtNCW
kyRT27UMaDBFOUT2qPa6JCJzdGRIdaJpzzuQQS0A31w/LN685qeXZ+RAp0ToKas5Zm/2MWQbiqOI
hsqVFwHRWkJMUCIo4D/VWCdyEEop9WlW7Irwgcgf9deYMJ0HeosYnSg+NZbpmofkwJEhybEKrA2z
N0XnfQHxqrRgU5BHzJBkov5NcMmPJRYmg9B6PYNcOTg8gEE5JRmXZbNdemjImourLQnubdxKzHl7
NfXHORPN7ZaW9YUnTMjg9fpIv7K1SwygN7EExfzi9VFe9yTCZMaxdWkhyvUrZX6BFdnTnDQse/HA
HZ4mpn7mAOCAOX+OJMJtnGaZKRgyRkGhLf+r2i1M1yb9O6KSSLiD+naVc5AfRo9049Ncn/kROJJu
SVeODN4+zu/PU8/5Jb2I0wg5BQ5EXkHvqKXLe0mfWrqpNI2IWMMRk3iWbClhsNl9p0B3U0Su7VoQ
mMQxKTRukX2kfz5QWdFZxB8pnbebYdj4YB5SHJ4x5wbP7XnVQHZjYP4ajxUDViXaIXdZvVEU8x/+
NGw7aSwH8mQ3pPS0uc8SkYx+T3JIPnmM1Ng5PlCup9ZcjLVOxWUAAi9C7fhOQP0qSLtU4RJkVdJk
cDRYGqN6yy/dOcXyqE1I+hSa3t+PQ/tvmiA7ZhPabbMaach4AwfxnuILdiK3UgzcxojcL7gXVVOI
0UMgfeGHWTF55ZhrXwjJjCUc5w5/Nsv1kQ+TmiJM4bcbos+TpmAR+QMEgy1Tr2DYl2WVn1/hv3hX
Csn++FoT2TETExkQesAnQL7BR1FIBFvFQ1bzasNLJx8p7F0F4CQHUsDR9sScXNWvNpncD+oX6og+
71gjPX75XMUdo/S6cEwALynStFafj+CyM2hbuBsA1sqV4k8apv8enZrR0X2MA9BQ5mDBtvzSm4eA
oOth6VEe5ZF0Pd9CevWfykzaIYbl6BiwgOL/4Buzz0JVs7twkIgPZIY2o/RYlV8z3buYbMOdcrbs
0HiZvhmOxV3HhUyd+h1SBkZhCBeTaIzjnNjV/lot7qB9toh6Qcpc6/b7yt4TtuBR6MV87N69awmv
d8+6zABIRs0coNPFzqTFyfk2rpQjY4odi6Ok3w2yQ1BfPG/Si+o0IzPHRqcKZw0WpzsUE3Ajqgao
GiABUlyfB8ea7byNi4aKfHYHls8zdgZCcVp6MM6I3RbKx4r9S56jZRQYQtLfest3aGNHOpg6PNzH
xvOTSNXBIVlwg1abcj8TQIzWMoODqQvrKEHFC2TRM0UvAWcG+IRKsN7qTTx6Gc5fk98cICEaSBn3
VFeNWxx6KRieeEPeFLWPN6jwlNxZFcLs6JfESgLNtW3FW9eBuYTxyIJC7kmOTe8FAOvmG5b3l/UV
1bfHOVMdlIb1+4LpRec0Hqnv5MyK8cmSzgoGehaYo90O0XmUTKxXmVxO2uorQTNRRI3aoT+PVTis
b3/jVZqWt4kxb4aOR+7twHq78mGj4q+SBbEBL4FB1MOcGZVUryoWXAxAfwdOB2ba9CIGGtESTXsQ
hzS1Qklx0Ie8D4Im7CKzpX5ym3we88Puu/QdLgz/Y1hEsw//FflSz6HjKsef4mRYv+YIzHP0ON0o
2V+V42gXGyyT/30VebL/E3mTHoleAx+3hy20lS8kgMaylFAAz7zug1CqhpKAqAU7mtFDtro3JeeB
f0ooHJVU8Uw73K9nohMVBmjaoO7A+UjLx2XFZ4nCLatRT5a5U+lJ3Ro1O/U150wT0DfM5jL8nRgA
1p3y+/rDAsrWq3qyqMHOHihm0iw+V/nRfClo2Q2XPYZ8nEoGNDgfiPJ3oBmiLgTP6VFpu5noMGrp
Mrre2r+C07xC6QWUOk9sPjt1WAMifgcyuSCSRgIzWBJsf5uch9+cKo2p9LpIALxTcZ13+fsLUq6G
zA1JcqBHebv/BMVt6dxXgwK6/+vDj9l67WsM31iPFbq0G9wwYG8aTv1IdqZDervqbuvXgUAjHzKa
5Hz1mPZVFwlFRz0O66ZBDqexse9BIGRggOEFZi/ND77c6riMzBwmYKlcHbR9KZwJ4tgo+tiGa0jM
lZ7KykeA8V42mRilg8RqNtsq7+2mz4QJZCajCjQGbnh6S1y4QH0VjmKyXVNjSjW3AKUXogdiEZ9U
x5m6JwLCau+mRQXZdxa0/sb1blAnM6cL3wcz4zVWbzjnbQ7X6/TPlsKeSDju5VuJJRgryG79H3sb
DHaulCuXnTf/vwDE/r2Qywut7V1MhkfBVbtDNFZpLUM7igMhqo/F8v/wwkeoxvnkv1941tIW6yPu
aifKpWbPVteds45H+BKzaiDI2wGomECdNBcMsXFvJ05MidUL4evCMDzkEMv8tsew2QVGBhUDCGO3
ODlwSBA5m1IxljEzpSXHus/Qb42DJNVXpN8FjbNbSBxItIJIfiFzUDylOAwhvelg9woP0Wc4YWUk
LNC9JHLvJjWtP3zSmtVfcYjjW9ktO90P31nW4qbZy1p2Q/RQjobwXc4uTO4vxb1qHlDGkvZ6EWqg
L1dsA4xLkubWnR7Dm4gDzdyWsQ4sgjqOias5iy+88moXVB42KfMGDA/R4UyBR+6gnePIWmeqCCpy
LM6exYMug+I7q7vaZ0lVXWs1jlh/NvaAlPJmIwfYIr6fHPDa21Qssuu/YO5Cs/B0e7YbChQDmFEH
IKrQhordWn7rDYSZ9f4hPc0T4A48kfdirr4sCxynqqUOAYGw+7nibMn8QFPENTwj/OgPaDT9xXJK
BSpdCFx5EOlHA50eac6YWj0F1rpcAEtSnGhqCwL75k5kdUiOuQSyiBDy/xAg/4/P3/l/5+tweg8d
w5A0KkvsKmB5sHa/ZzURB3xyje43QPTuC8TMW3yrvzYFopx9jnL2OB7G2o78Nd3oAouWy+rgKoMg
+lS5OSfYVttGXzCkWRLluvqPVA7SbyFN5jOAL7bILTVZQvmYjI2K+zafjBicpYEZh4qs/DEr8N6o
Np+6v4cEuaHYfnJCr9SkMH+LE2hwVqZYClDN10h77wXKre4vMQZmA92vWKcuBw9h/ukTVmO4vIAt
nbHLveXt/AQgEU4sZsfVeEApV3he4Cmf5CJLLet06cjbigohYCsYgu272xfxDFI0CV/p2rtRaVf2
61GBd8AclZUgwzF841YI4StodJnA9b9n932J8NePtC8yarj2rb7P/972QH6WEsCk3y5SOoJ6IDRF
AlpKx1Wh7ZXkMXDYE6WOvQruIIiJCT/eFsDGmTKeRMwUrOlZKFM9IOff95LCv/Uxy2xrdpz/mDm5
MrCKK7RxgY5SnE9sX4NPAGCyuEqFj3eCs2dVFCBxFsQBvamNhrvDGVopkube4n2VTwdsZUNRrhr8
kdGsV02EbLs+rLB7nic2/g209Ln2l8qm5TfjSqWASblrfp17SHZEbf/fT5SL1i1uf0RMK+QD0dwb
8PxVZlCOncmEF31QG3cXE2q41uZgjvh1fqtDIExCu0TjEQwMOIgyqMWmmZfPglFCelDdAZcy1/x+
SaZxGbEwfZD1fu7VwaRxVCjFZHB9yaqw9xfeTclzg8rWFvxAFxzTJXUbF/19S9rm38EzNa+aptu5
hTDyYUZnUhgcp3vQsMeTMaxPi/HrZBPUMa4qw03VGpfR8Ty3HY+feKJk7LDT8JHYyLNsvU9Zz+BU
o2FnticHYIUc/7vfzEqQZRlFVWevI6+08FUUx11H6crZ2MEuOkR7IuI6cZz8foK0OEfl8bwCbqEN
qiyge1jSxSH4jDrcmxuqo4Eyi4lrtop7UEub9kVPfdEz1CrwJugjyCRTrg3lLeEAdzLeT3P2uSMY
NijI4fUGg373CMuavLg3it7EmWKcyTdOI8iKFv4LTE6gb85bM7K6dgZjnBYK00HJxPQeMgsHtYev
yhfa2vWgpLrsUwIGZ7SLHHOXhYSQ+osMZ7qcxzRb/s1C6gUXznl2YuBpeRf7cAJ6voHlYwASlqoI
S1qz6wQ7YDJcaSy96lnuT1iDRRqRc1MqfLPYIXjUI8EkK/D5TVGzCebV8m7pW0tDZVVtGstgo4PY
yCFE9ChwfIecMstJTCRLujhLYMdG4g32ajq7Gbh78ieAXOeyYNqUiR49UEUFAOrIIbCpBMof1jmR
NJ5UuGNoIACklS543YtESXRbUEz6JlHZpm84bI8nZ4ZfOcXK4KtbeVJxRKBdOUlovVCo2cHkFurT
F1y0mrCGFyo5fay0s6N+jocxonr6zWtBXxamjc/MgT/Q1TQ92k/hOjvixvN9Lb1WpxyL+Rdj0vvs
K1q2kNWofyUxmeIUBOfZmEqROxx6PE3pARfoRxUh1rifVtGzrJRoQBnFA+RS48Jacde+3nMarrYn
f3sqYHpuiEOMyfz7I3n2TVKsj63XLfYaHWiq4hmoYAwWEmBmxk9YVOhxRYV6RVojb4DZUvLq4SWR
55EjZwIy0vjdVbym8xH/WrceA42iNHjYTJlbRuDGRw7EWJFp8jFX6xkFxU9z9ScgPRKn3evsN8jC
nRK5RHUEX2yRY3+iQKq0S2MdP7e6fFbGdSLKxII5/ibD7wO0eY9SwzRAmKAIcGXioIuSpVI2nPee
SAc7wnkuBB3i5hcH0wYRG/6Xw9Qr4kmFVcBOz8EGRWCLp/Z97O1o6tHMyfRe05pmCHd5W9YV1J1I
WtIX9eMXIIbsDvW0xILuvmYNyDNuUfA6rWX9vOo/1he9jwsihRgI37GQHVeLihVtVSwh7QoZJyF5
2f71tNX2WJzGMHByM/a7D8W7kR6+guhw02jo65bgXRGgly6D/GB7cmjpkx8nfIrYIvz6sLi3qJrJ
oDi6L8JahwLPIQ0rEOhH7CiPxN6SchvsXNnZG/Zi3TJja2H0hiH9QAj2VvfLmSCM94GRr/53KVmL
UD6NGLd503aOymYxFwWAOWdlKPtADrZ1RdBbxtF5NxEUYCj5Ix3aqTALVyUrDfS9Bi1+VbgsROm2
Dp6KrzLoIDaMf0gnlBUxezb/sysG+l/sJy4SLdxIft1S0w8xbzh770a9gj7U7k7ClzFyZOtJP1PO
LBHhBoEmm9IO54A8xT5D6kMXI1Ux3qu/L5c8QAnOaaI28n/ojJL3uUwov9RaCyHfxTHc00aysw0p
0yYOL7r6qWnXp1LYHV1vuyeIEl4zOpqaSTR9wTFxQBb+lnlJeS0/0NZKxryJxYFY+51dtaKFfTm+
wKHN5VxaJReb1SeFpsA6LWwpHsM/N66Uey2JdioCnMF32Bs31HCbRnOj0EiniiUJv42E6sgZLbL4
0CcWFG0VzU60/ElurqQPniMfQINzdly5PPW9U3POjjYB32I4STBuZ6wMghY1SFuz1j5U3WqzVdSd
Qi/kiahCiSuhcdsri5sw4oLyZcZa61gCoEKpU3+NgLsL32DFF/8zV0CK6NyX3rVO3MPAXO7ubeqd
4Q+z0CCPEE+yBVYJDNHtZD3NoukDm97BC/6HfwaS9R5DOTiPiLzMmB1ci+txw4DIslbG41uZaRtZ
EAh/tpUTp9zDwCCSC+kVtuWrOVmQ+VG1bknyTsy2u/5OOtUUd49d1QF0T9HL15LaBKpwgp4cTVdx
HYgUJ3/CcKn2hjykY8MQmHrNwqtN3XlnWKgMmuCteHTcd7i9FeT0S7OC3B1slxbzWxvuGVS/ZoAM
EMELddu8m3LoLVRcECq1TKuQBE0D+iBzcrV/uJZNdgpaVWP6DMGYmQJGxTzMdl8T/bviFG7ajtLT
+hB3LSpzcgwwMB74+erQ1u53mco2dAqWDpJYkg6iciO8vdE1d2qd1XC4UomWVmzoc+RCMxn8HQTr
uH0n5ciTdq9i8bl0G/pMWPV6bhS6dCzebANNaIOo/lLiE9Po4H/e6GZaFW/PUqBe64/pToJt7r64
echXpqmottgZdzElVxO/sh8sSOC3t4y9p+T8XxXlC1skV3RCs9dge3AC5iXaSy0c8qyjqIWQydlM
ucQ4xxduWs4L2BmU8i9lLMjryP1KjMoqSOyfQIsk2MHaD4PrBhNVh2jej0L3e1TJ2y1DYqBxL9l2
ot6kwfgXHY1ITDO9Z8Ch8vxwGphtif1xhTFwt2yWtb50/sAusbct5W4REZhMibsm/5gCsCsp3Kt8
hu7rglzp7+QEmV3glw6IrTQbgkyVDlpXzFx7Ro3paxLo5/CcBIUHGQ/IxY1SglT7s+x1i9JsH+OC
MEIad7xs1hO89GPFTgmF9jq2ansbHw6EGjSMSz6vOiuj4QrEd8SUVsDGHmipZ1+YSq7etf1/gJnY
KvSLpp0tk44MD2DNf9Rpi4Yx8z+KGh4P3ZoDTdQSyOq4r7R9Ya1epmn5/QhLReRJ031qpegyj9ZH
s4ChEnNFGBp6vyZmEfK5tk8Ek6el/Gi98gwhOTT9Uy/n6ctY+xSldjBLutUqRn9h8lFo1cINbmln
PgCDqRna8SCB7XyHwKBATqdNOJ9ebsJXyHuyS16RBYKdpVw/uOv1CrYP8hsclEd1JrS35Lj0swpi
2d3S0dHs3epW5Bzmeif+AoVvRFI7pr9oJEkOZl75nPq0l8YIwivI8IN4WgrvzDWOg33ZHWIzu9lv
FmEQkFkRr5xp8D+mH1bSi2+B+osffT0lDXf2zXc4LyOevgtnNiDZmG5P/ZOaROEzhaXNApmypmQt
yMh7wFUSZ/0/MFBMKoj6spxDZ8caBe+yGE6vvgJ/gRqQoezrpik2VPqbNs2EEucOuocDPX6Relcf
M7zz6yBQygMCwZaHhrF02F8uAjZraTIGsOwu46Dk6ce3s3AY2Exsn4NOV1CdYq2E37ELnt/J92aI
3nHmtZQnDTCsxyPZPO+PvU5VbIdj3+PdnAgc59NqHhts+VIFUgtqwLTYUXw3kyqF3Hiin1gjjYN9
zCRs7kA/y/91pY4nW+FwSIT2yP8cq1jD4m7lTmH4Oa4SyCXBSR060IiLCZsuPysJoHGjGl1gfWq3
VQNZDOtFGMIt5MP8tT8MwGoSoY0pz0xCr4bIFJOb4f2sTSTW96P4ABl8J3VbzyHQ2rsVICa2Dml2
P402TIHSijjt2HLXETTZrfSCNEFtCmGYVQW0YK53UxCceLhqI+7JWp5UcEgHvb89SULQqZZ2HDFi
WACxk/7tqkzgVcBE2xO6lMf/2KjYz8zim49FXsanQn4VwevLoPYiZ6IIOvP9JQ3vopr2RA/69BxC
AWXUpDpEGH28Z/IkJHh6HcmzKLFMankKJeI4Shyu9OTZEDCz1INtfZ5zj2SCobbxS1i0k4A67LUa
4ioj0MksOW+OBdgNNs/xXwX03k7BsPgDh3wYMIcwegQdPpV686hZrIaffSoL/xbAyHmh5ieoch8b
y7lX7ggKgQUq9KYnF++tsD+v+7758td+vzb8kLzDIVp2npTz09AwSfsdAygLA9NSeByI1e2KRYl/
nfz1xhhMy/jgdSixbUvGjiGQHwFkDLtG+QCYONvS0QCxP/7gL/CRdn8qI/uHxJRTZBieTGkYpPHC
3oCBODgwcmJrHI5sbYRk3m/ZEeSWFw3qaPaO3bWkasfuuD/kJdr85k0hDueuMVjJkgTLvA2oEtEB
I/KWlQJrt6WcN3Cweim/DcYZaDgxSKu5wyHl6akluyjmiOybRH58y8FijfajXs+dYxYV4hej9LYJ
jFzG7mKyiSXqW+pWICkwOZlyN/KYXagir6D/zVBNXkCYBxYs4qw1TO6VbYgGzGLcmyxsngdW3wRD
pXSXC5g8PVksEPd8FpHfj797GAR0q3j+++TFsdM5Xw5tI0ETc7I9vKl9HKt++tsxoLNVdRj3f0Z+
r41F9eNMVS35vh8OmLwZLH1w4X3VFO/Lr/TSTLqNJzzEBNtw1Hmwm3Vxw1H643aDvJq+dFtNEU3R
c83Yaj+lcKy6eJ2LnhS4ydYfQflEIcjDAkQxZq1mG9AhyQJbzpLi8kMw69wAgfV+htlZl4nBfMq+
LmtI1NjnDgikPL0oZdDOHE+rlybSFsw6HsDFCoag9RDSCKG9eK4Wj7LPHjAgPoZ3y1lWOuca31Qk
KOydzgHDeim1Y7m+sadY67jMIgDq5RO/tKPNsjDRMbhQOlXhXis5eb/s8nEYUzVU0zG0SG3W0teM
vJ5B5XTZ0QEbIFw7mAorsmMNvBoutDJv++Dt6R609bx+YCDRvVD+Ywz4dzyTO8EGO8bTlxCkYz03
6Y4OMxzfQeKulyiNEwpJP16GCSSQ4m2T4+YPZMyi6eCZslNqpW67a5DdYVQrTm4tbUKzie+odR/A
kIOGKaN/lIZpRCbMAc81hZ9Um60ToQWqvL4tyjHmYR6KJRBjOYuGRU9NA/ZcPiZMAef1gcZGFkbe
Qdp9G0MyItGrAPzJKgfkprFCMxAgnf5QdUCSRsG0LegKxGoue2yAnboHfTUv1/G4Vorf2FeMe870
hRiMAB/CwgOQgwZ+G1ihU8To0SJ97GndpWvVezCveOgFfykKmfW2oR6NwrnngwZprEnZ/O0yybKX
s3eD6gQTIOlJsE7bUtiXBN5Gmu8gNIzK/brxbkgz72xgtziP+fg4sBWcHlb0lUAfld94qDIYBORr
OmXcGsZQOeeUU5/kki62qfpH+OgfujqmlMUX2kt9FJ06JKQO8DFNgXQkPemE7YArgLPcB0fHCsVy
/E8oI9FDRfhHzw6PeZtBju7Ph3O0Hgm7clFvweOzKvUmEmujRonszvcr41R/w5rs+3l6NLOxOQvj
lYpaytvBHDN50FYkTCgmFDOGFFsD4UO/MgPmgp/2WHfB9SXKTVcE/wYxiu8IhQ/PLnPRCsHM/D8N
DZToS9lCO5f221DsLwQ0tsx2bzFgflA6KBrh4DNNIKhSEcsMPj0s/XKwnvKi1VW94P7Xc2738oWx
OXNPc6YSue0T+I5jVRqo3h0igpkNfsM8kHoY0m7Qt1JjrLgEE3nKRHypafo+LGHr1gvRuHYxVhdt
jiMc4pWiTBiz+JIv2iI5ES0NCez+hXCXtDKeGrH+EnIeN4aKxKezohD5ZsZ9NtY2rKcGQ9UbHcuU
rtYp+XYsZg2sKLUHMdhwZlCd2TDzlL80CkP2dJRtC4a8sXwshoLvMFcwZRTlYrxmw72AdN/L30Cc
D2g1wHkl5D6OrTrtQ/4bJQXWqtnSJDOxJ4lN6ReApiPxeDW2KS8JotFcEwcag50fcFaUdZbuAQM3
dFle9XZMLxCFljY1mWSp/eQOTNuN145hzyrsb/g44v18dBKh0mf+99bREgRygFvvhhmfGmdjymDl
f6Vhpc91xTa75cVvhZHdUgXLIF3H0kRlciyTi7UCzV7J7UBI9TUQWfsN10LxnPo9/RFXYLsJ+b4E
3pAiiMcP6by8ssOo0jH6KFtkKSFecMkEY8+JgrrJhC9dcY6hxwFL4hKEAd3DK9rRH713oM+SoLoJ
uNAMqlb9U9hZKE7xn/m0rsKSyCCeOpLoIruxHtq+spP0rp1+YH1iho4rDgbO9eXNtTrhzC8pnVZ0
r2dOUQbfMg+apg8/vHfmPL22GwhuZMCCqZZgdYhUW9in4U3N44pzfMXGg9SUuKYf97/VN/jXu/jA
Z6Md6AqKsOWoYbQeUkg+/ZBgGk/JUZWB0gUzTkScb50Rwly2PWINAb5xtxrDesQ2T1PZtwyIzzeD
rrxwPOYP/Q9XYLiU9I21wUKahyWRjXylLNFUPsUkia83PyKYOQGV2SJapTvRrKy8BaRc2BjJe0iB
WazBNhAdZm+9BBDlRF2rRZev+l+/ZW0QcqsFSbmAyj+x8XygPjg49wMw4Z+j/lwtj+iw97zadnvx
o4OsYMw8RBK4O0NE6y+Pyp6/pnmqnV1R8Mf55WtGL3wivvUVSWn75K2G+VzHb1hTZvXi6EDrwu2R
vJ+bBbHxf+cC6WnNwNVLkz8aXuyKa92FPlecrshA8R4j2sw+S/x/hwn+aX9KpziD6goNnA4Ewyk3
IOPrK4zlxQUeEtjGuf/guKUuBHWy8kWlCbolAtH7BffiDcOJ3qvwv+t1KVybAebAHbkWPE0MFKnz
udJ/mj6mxRlndfA1ozpjWlu+XyuYxT1dADpFZ+RjO8vLzlJvf5x1FBKsguPF9XhTgWSAoL67RI3t
Ou+idnAmrNnu9ymFzsfk1GGFPcUv7xYe7w1hT3sEW+DLUkfutMd6G6pEc5stE+XsZEr9UbCQxETk
FHg3lgnBgXb+N9+3dMI++kya4hJQiC8b4rYqWAn2uUoE5L3ACFQwOpwTlduWklCqfzo5+mZBvNrP
mgS7BCfu662poYxESPcWF1gynt9uilJvXEJ+/C35fuPOyToG6XBGzFdW1ZLrse0n1o3RAMD9+pTg
CkNNbNB7jUPXAZTU5PnPLTBry13TjSp5WGcTIw/xlDxiOx2K7bnwUu3eP/YZe35K2xvaqsnzoKhL
hN46TeKzUfs7p0o5yKRkqG0qF3WHCBJkOUxTaSBisI9+i1zExv9s0AQUSnsDMo9I3dvykrm1kMWI
4FDreQuN4daFFj0DCk9W4KNLbIxSS1bbiFJRoaoLa713numXHTks2/CyPrGQSwMr6M4U8nzp9kP/
ajLkzgSJB4DO6MFQGnK68HXiA+JjhTPyF2+YYM+N/Ngm5XB0il1Y1+tckE10SIjek22Q/9HBd8zR
L1blRDz7Ijj2bsLhvvOY8be0ZxSJHtq6K3reHq4Kd5wOU3lknbaUNWNee05xj0lzuQIdXBhleyzU
umw+tc9PS/bnWISNEkc0WmYhZ43URJpVyUA1jJbGKSfhBCUAUG1rBcG4WY7yv9XV1s9Qh+tQ2N5J
8WPsLAv78aGWwI/DkglGcUTevRxN+h1O/rt3KehUxKMNnbozYprLQ+aix2jIp3rPQWd2OnlBk0U+
yVkfBK18qBLMMiDgbe22C1BLvCGe+ubSs+wx9HAuxRINFj7oxLLthz605z4Lilu8mUcwu7X8BVuu
i8zZ0jNthrzREd10nV4kRhtOLoABxM86oFRnRLacLJPLh0Sh9HWo5koC2/+AcfD0gNXv0J5xbuPh
xgzy0GMRH/26xbjmzEbKypEJMA6dCF4MhFVuopKcac2RT8+NDGoTdpj65ansfT+3xfBqK2qyTEvy
s79py+B2nhnvhvUB9izVY15dP8LciRQaxjkWDF4qNZoygrjqzny/cCrxbtIAvGQSpG6xHBvr3ew8
6iTbtjOCjg8jfI3ejw/8sFhyWpu9jGZgF7n3Af/oBsMr2I7NW/C/6ELLhWJj3S6QJGBQHIAj8gXw
HNapTaQjLY8vau0NsVOKRryYEuCBm8XmSz2JI5xHi5UtecQytYasoz1JPnmq1THz4F1Ks43ZSFUI
ASZwroKQJRZpE9hxC42zXywzwnEnURXahh+DMB7zwYMqxVauntfUHXh9jrUQCg0yJ6WCCxwYwITi
nRdAfzh7jVWyzTDwgL2SK8DTR/In8BLa9ak7qE9A6p6Sg55XeD//dkZs7ZmiSldcJOTxApeMl7uf
c3RjgbAj1ivFTR57RXLzSnuUNqEwOM1RcGJWFuE1O84j9vyBiouIoV4j/fGL6qLXP2wkHGamEo5e
dmLA+oDjDejFNyZUGKhqbz6PAhSUXTgzvlUqpZw+BRfIP9/ZOL0tn6rS3fapFXHKKSCFo73LW4Gz
1h8KuzBQoCx4GgVlxJG23C7Z1ydMgxD5VE0qNelRhbY03PZG9beGIFOfkbwUzaYUx4DfCocBs5ZB
BmZmi/Pw5uFUHpUBhLLRgPvBiHE6bdRl1qv7WRf2ydIbGIp36lN3E9a7pYFwBUoXbDm+A7+g4j7B
nZPFEHgzGOH8Obi7gb/oOdKFQQIOTkVkd9gXkosAYUkvSGdDr2iv3pn7W3PXtrqic4nlthA52lKN
euYTJCFoDsVVwFreGEc8TkUxIQlg6U6hWvIm+lU3TCX3lTTK2m/nYwF1nKMYGbvvTxpPjV4VvbN+
IckQW/cwySnSbjq8tntiU35nwxZeA8TKQnqxk4Xk21GP+8ml7dJOXjpH8wa5qpLilVi8E5FGkNWm
Y2zMfoFFOK4mwCpFsvyMqgwOQYSZznYJh+FlTAV0IUSQJ5Y5TdXH9M/cu/qmRQoTlF9TWawJ9P1A
BfDAC00h/TpOTaRJtfAoyaldDGSkSgv5CsduC0/y1gvEYmDYJD5Wfrgcx+23juXn+ul1PGAvP304
vRzF4J+xqi7FWYRg0c2M9M56m6ZYYTebiRJYVwTdhryhxi84jAKX8gN1vmunXRCl/dHXYK2LGhiR
EI6HN+ecsbqZ1K8bKNB4OA8fZ4NEhJ7ghzzFfqzPRHZPk+RrrarhEKq3tSvRDME0MdahcBbl1WuZ
7ff/U5R/7TE5PUWBkB8n43xqKwFMTgbiydGA9odwgLNqYB+sJ7Vf5DKNZRredTqOS/gP4EMwER7v
6k/G1cDEeapF2pLlRdDkvnsMfG29eJ69RA2mPoGRHklRkjAQzRTj3jANvL39kK2JE6ZPc7TiMTIA
3+11UYRmTR8Jiqy02WuOyBR/kKll3/HZWrF7yhLidAIgCyYgXZHerjlU8xzIEQwA4LjFD2kacK/u
e+xEE2Gbi4TamA03e/H7RhkSo7SkRuEw4yY23fQbwHvbxfzlx642GjWZLJQmDobhgNjrpsjjVvjq
0oVaUwZMKCAYnrqAUpHWMy0Bw+4wi6ruLy5Fi2ONptYr7H3oyHCflV2tbRcxmcbqfB0hMA0QSE5M
ZMYLjP7Cn7Q/122IHAtJv0V7F7ImcIsIoFJZiL/1Ji8N/7EokLAml+Ocu5yZ7VlsU8ODKz/Ama2h
jnT1sxZoJ8zY7zuSWwcS+Odr/Eb8RI0OmH6bRSq4NYnZLlzjoaJRPGTkCo9jYDOvzwQGyZomCCsK
3CW4Xevtx+t/3Qkp0UR+mGsDiVPadDmSlY871xN+kmfXmzgMp5zp6lmU17lqfQydHo9xdfsi+ZNT
icEWuXhkoLeM4T6594u8tNDyEn0NI8fTvFG7JLJOE1pade92yu8euEJd2PODkdpkcz91OI1Bor+s
l08t03y11+tPmDcCcpcjwKL0qx/Oj4W/YFBlyjRnjd3wgq5PweiNWYBWWCoW0BwZ5ljDC8qB4u1E
xsSRm4j7056mfDVYV64E+cW6HW8W/KigDU4DcfQUbNOmXf58qbP5Bzj3SI8TrYzaJ9jME5RFTx3m
CLdct7Jg1ABF4nqHYSw10VznI+3xMiiW559QouIQj7tlOZlFmTmDzAVo/rJD+VkdLvkx3SGGih4g
Sxh2NKtZ4rjoYnNpjrqoDd8519Gkil4BPy7+hguer0SIrdss+cgeNsWHuNq4Hz1h/zO6giQoZO8x
2iCF3Rg6RAFaFsc7ywCzH6tcUOP8TuvxY3xbWH+UL2qDDtiOO1P24EcmnLKGShWF9c8/dv9eLAx4
UcAvzStzmJlYmw93xc8r1JQ6Vr6SuiUIX2luon2HQiPSoKtiR/0/sESWaNQ7lYY7rniANhknY1NH
sK6fIV3YSZibH/yDyKiGdd4rkfnHASPnNsaBHmK9gy/SlUwIUa1vA4VKqB8+KfksqKO7iBP8kPZa
rCnuqyG9q1kAVd3Yfl1PCXhGZ/hXQBVMQHOqYEcO8Sn1EP0CoFJZZZLPuvaRWK+wx6evehai4+rI
zgeDo+CBX9FRmDDoIclBALl2ai5R0c0uNhL+ko2/nQLdx8xqIIgtgNXVCTbMlLNS8plNoDirGT6L
p9dGmDmDsSfYx2JBtzbVm7Fr0EFLopZK1JeIY40iNNps+lVDtkXdd8sv5Qn2ZmNbFu9xPFzOalf5
NQIQPdAnUHAGgPMMJJEA2QbQv+4d7DJaBACjO9/tIxTnt05+JOLNXmFboYQU/hVRhLLGkGZeEqWo
s+2ZYZ7ZFvQXqfkYnMWMhCmz92F9uCmjXfqehmmkKN8wryqeRpcIV9r8jcHyMVbjA4e1bhNybhsN
TE92z+vJdXuFSWOGInl8yiOGcDEHNzO6IL36sqIOoznUDbooVCp1SO/cDqYTrDrhzqMHFVZRImVQ
zz22eilEnqJNUnXLZ5A6QMiKl5fzOv3ejnBf+4xnovMSDCluTygoqMqxv/Rzn1FKKuLnsGdO1+N0
DhVGEW+AwgAGleI3g5zqPIAvDVjxatDxzL1yoOTl4YGa6PAiTVlAz512KP5sYfMn7PDTK8QHLs4i
KNSAXzvKcdCBqaDJkREQ1YRjw9Lps0MTzEtFHq2f8ZZmN31MKc6JRpi8kbmg4M/gk9wZLjiwFOCi
QZuY7Zmk4sDleOuhkYRJIHNkHjWTrENEDjQ/+w/YNUWwI9HEvxFxeoWdznqu25pBEUt7QL9Nl77I
Kataq6zaBypz68zXonWvgSzGhQY1VyUksWBaaq+I0A72nlpC99+gvoCWZIo7HGME8wyu52ELO+Ez
jZi4Yy+qJ8LbnkxoFzvupaFcjthwG7vtWlNT/G9VW9JuBkdN8t7lX4Setzs+B8gOqI9vhiUTjjWf
d7H6cceXrG6vdtk37SV2/Us4MHx6caI1rXd509qK54bjHDLj/4nNrEC5zU29S9YI/izgdUWoboTv
CONN1JDEgjRQJ481gMfKsRvJsC14yLVgfKX5rN6wFPXSnB3zTXFuyULT+q9bM9PUct9YmOcoZVg8
fRRoOWgd8lJv5Sm0DNUi1tnD/5QitOi5lq4ATe57urJDiLLOfoVjDQYA5xpgaPLas42BDKNnWtnX
UlmVFw8nuTd4ee8DTbGEYnL9LCMffEBGzEG9cK45F5metU8J1ET4Bl6wsMfSvtzEuyfA/j6X1TlW
oIrzjGElvHZfC5oknva5y+8dvQvru6XyzJimg5iGHlIErDlRVhBCbePwFSpVEA1TactMGJU23wXa
TF+nVu7us630cfPeZgGXkOxmZbrpoWp4WZkofruKXSWNqoxqxguu91gF/lWY4SvkSf3M9pB16wVh
arY1SKNsy9H4sREVzM5cQ1kF8GVKmIYhYnuCjtt+ISUpCre0X2iTVJWPlBc65L2sKxIaBFFXCFcJ
rAgffpMPYdVKX0anewDFakWH9GkMaiD+3tSnbGw2h6+4NVKA2O02mHK+XdBW5ewmsHE/NJ1IOCgk
mwfFJ82PQKknU7COvA2UcejPW0GskDuMs1md+Fl8Gy+g4uFGn+LYUiVgnWz4eo5aLBX6mGCwRWAG
hq5ageJ/7ToLKAyElOEFgdjqGnke0BcrUF/OoEXg05pBED5aEOXZyb80o+Nkxefve4ib4gQB8sX0
dO2NxbhUbUmJx6V80MgTjbMvUBwSMod3RZk7lhDkov6o1q8j2Bru89eCUQjaDWmmfXVJObRmnFI/
ALezlcWT3AyrY6jG2kQ61+4oz4f8GmFeXhJ+VGUtuWQ9VR4rJeUclsjpKsPEowLcQPtiaHIe1Nzm
nXKYo9WPgfPGIx4J7bsNZaDduoKfc1JKRKBNOGpwkxP978+hfk14LpsF3y09jeNv/MjTbovX9QHk
cRgP7MXQYwx6sCQhrdgqQIeR6qxwoza21ZoI3bRiZT6tefUkj+jUQbliOJJoJfg1920iAVdtqbWZ
sZ/BH+pnqK8BULsAAmbv7590e48kddcCzjDtKv3OPJ0Gb6/3P3G5iWZ91JdNF02GI17QOnZGG8/X
aMM0IaOXI5FR0NEhITp/hl1+HQnQNzfk7YAAFovPL2EXx4VlVUgG7Kv5q4vie2k1C2xTRWt5sGsN
lxIyZmaSFrppPVhKImiPpFk5OVo2A7zr3rYx1RdfOkLN8Qw0PYSirxgztSmHEWPRpZo+pz+8/U4L
6Mep/SfhwJViGC8UKdIhUZ0mP2nX3gMFOm/rBZjdg9ohl5ot4Xp/mjmTlpDMH8BS3ib18MdOyA+a
WRV90m5aFOZmnC2HGvuX9KuEjQQO3VLoaE3ChGvP5yabXw198PTJOndiw8uMgq9xWbXVk7dKywoe
EazWaMHprFMhyleR8ijz7Ug9C+cQy29V4EAACcUG6T4ZtnWhZcWxWHGgICVCVTF6ydX9RAfWnL4w
uUTAAp1t8psUduGkuQzEBPG6tFXIaqPcgokUEhIFIN/9sVwYGT+u/UgRKQoDF1iFaSUicwmy1OCI
cRJTtXgzE5J5sZCbtGBhH7+EQTyrbrnyDq9hGRmtdhy8eoDldhUB7wCwWdKKn0lndIe+glheZjoE
y2CYFvpdmXAKqRAXcwSag+9jfmUAyIhHahI9ObI8LvnOaIywmYAm0ia0kgmKnVjo9UpCEsbxehQD
ryiP5N9RrG4Xp+DZ0F3jJBuBonrWPWNfoPQ83YUi3mdpW82cdcVd8T2NcU1y6kQ8flnT/bflAS5/
V9lXxqszWeaGE//TsErlwiBLu9JuxPESLhgSbeT7g96+C3/QRJN6ke0L6LWId/Zis8SHrNBh30id
eJkxnsdN/UfzYK2Psxl3bWw7fqfO20hbxy0mAVi4nOEWUVk2L80r1Hg5Dlz7RYw71ZP/cheij6rx
O+SxytRIzrZY3fmaylq36SB4iNf34YzwZ16YCswOdyV4MsF5axXv31meQgqd+Aq2SSkqYsPIDx1k
oSmUqkSzqyyG3Fjy5CbIkXhh+N3BM3/oI9uKOFWpJXdXOZak/+8hfRShmuBEscNAw6101FWrVF5G
bhq0WfhGGd/f0kh63gkWmApxQx59r/6vm4Rx1t5tP7azlPODXuJ6rmgrhjXm4zy1HBJ7sdivSd7Q
FQ++1naYj/h+fQEfUHGCdFfLvl7W18NWmcRjaMJMZmiIgIfFVu9H+/a95j8EsargAMlsXjIzLIFw
dcLo1XDZF8AjbpFQGf+DuMc5J3+XwAEOBNH/uxNMKPK/Jf/sWxEt5y+da6RPHLRmIVUGolWC85f7
fRqqNc7ON+pTUKlCLaGWrp5F57Md07dpmmZCSITt9CdMiXnUou7W1IpsHiEX13zQH9u/TFY7qWNy
MfbgHmUKfnHOS+jMMcv3Xf4/QKxCaZmcz8UbzqYpg4yKmm5b+t5G4SXRlpUNHEXUsgYg4Y/wa0LA
nWyJQwPCthpJwM6uMa7WeZmCdgwj0NZ+8BJfPzsNbU5g3Hrx8vRoaaSogo52Eif5ZF+dsJVkD+MG
PC9/w2MrgF3Np18tiDvQGpvH+OafpQiM79oRZ9asVWDTZ9l5g3QhSZIB1p99naXT5H26bpGPtBdE
x0YM2RP8bMRZ4yFL5iXdycmI1/ZA085ZI2utDDqvy14hiAnZrzW0eTcSUFAa0LczQOvAZ0ZqlKeZ
cT0c/VhtUrRpJzPO//2iUTX3vTTlqPQZaQJvYY1EFdWOqatDkhBAT2eKEmP5DS9OTtdRlvaskQd9
9Gw/92DyKwDpaWB1QjuL2ISU3HS2/SrUUySlXzN01IP5wrCRHTBp6vbOWndiWI06XQpOSD6AmiAC
rydH9Y61V68PM7LkLR8culZy3L2+HwQvBaneNhfxkPExcPLUorEQzAWfwk+imZMY4/81hW64Nay0
bx0mi+5kcIi1GLcL/1JJRCCk+VP97v860pBWCvUuWhRNmxPzoMWFJDr6cVNhDmJC6e2xPwqwSZh4
byIk7HUEHF8Ssj0F/X4rV2keZxpkg/KkKgd5h9pCYjuSOpTK5K3CLIe2CCdea+up/LMDZJEYIWNH
+kd79Ramap648dB2rOtag3WOL+Sfnw/rzY0OPIKCX9weCZsQBBTLMewGtcbjbzqJDZ5uPzwy52GG
GhiwhJFwkYm+ioCIYB0cX//7UPKD3z2b1ow05/n1DCfitTE2puAy0pj4Z2T7CnyKhIsD7ZVWRnsC
75GiOThw4HYkxakjaGmyH06R/7yvqVCEujO0k0EW8fEuYagJB4ajfkrBeQG4ImNyQUermMvg4OX2
5Wfh9kkvjvdWGYqQGi8A6nJP7IG82bf6wxyRIIweBaVnka4NQzHbtm7cRR48DY3CdwByJwEoq/R/
CHw4GQO2qGNW4PcJGH8IQbuqGlHKqDdiU/gWPqF8dEmV3wDqmAdcCFfRVsXUTxm0MsZom+lGjkUn
XhZg3xDAtgegHIaSp2pQKx265Jkcuxb04k6DjEnEj47D3c2lsLaEedP9kvCF7FIjGDL3ucvyT6AQ
Wf0lcqkjKrC7H7zOb0bU3fxrUjB7L27ljucAp3EExsmV39nMqRmwpGT8ZLw6QRDfMFHfoYFDbmIi
f081RLXIFh/QF7WVhPeLwssJYqXD3Di2JBu9XRlTHVE844Jd2KwqMFL4yEsyn3tr7E9VaHxazO+J
rjeYbYgpKoySgDzGAh/ur9pxUaqMlpSFpRpmcaoip0jNkNYIngwW0EXaoBYyXyehFEdN3WdiTOPj
wNLZhcivB3bWwz7s3gFvPtdZKbhh7GORc/jdOP7e0vLUcDzyHw6N7y7Ve3Nwwm4/OFcF+/E5bcI1
iUozau1HX4vk33cI0AKB2p+Bt0pvyKZ2NvU/KXXTWlzD0px4ut8AcYl8TCwMGfbd8fgwAI5MxGi9
34g0KOUBk4iRDZsQDnBCM91VEoDQMqBeEin5gAF39wuDlrMAZB88MOB99V/d3Y9DAYTQKKeS/ngy
cRMu2bO6r+SdgQ6gtDAQbrumnxmEO7wD8vOPY/V+sqtlKAl1jvq3HnaorcgKu/7TmBpZxUpCLh/K
2ed6GI3EWoA9YCP6HD8Q9ahDwMMHOfLKJ13VtypG5VJCusG5ry706jYt0CLwAVIUGS1uXglCuvny
wh/XCfBI5BgsCvgo0u8ba8IfxfHmJGK5l8jUQkKYV0LGg++p+xpRMszFK1Qzonc3qDNTWwF0rp3x
2fF/+swHwbgu4ql+heXpLXF4sKxBGcNtfKgdBE6E1oxpAgvEm+UYzME/gFikAeDA9TJ5UKfVF+DY
5KXS4OhzuTgBDpuU3f9iP6trE32ub+ItG0gGHRQQi0umGt5tn/guQsgMPXgUajcPlWc9hn7uIywE
WGrxSyDyv8ksTbLBZTfTXTrDgmpAfdPlxJ9NDmrs6L7OGgo9cqXnijuzLrDO/2dqNLRCiBYv44FP
tQ2N8jnF0cZ79abCxNqPjiWPzlaOoL7tZq1ku99Dy55UiO77E/doGxzyGpHedPunHM77TLpMmwxu
5nx7UjpWW9JoWxISlHhxfqX39ouxYA9khIZode9d1dYhdCyJmBUjnfPtmHj3hHr9Z9iyAy2d3Zkn
PIhCjphjFYqo332147SPdbnAfkYeLo64gowpUiha5Rda4/DCjbOUC2oXdozo/oh3u3HfyYIbLhGa
uLQ5SfC9XLfMJnObCwVdkdF2J5BXUEOAddVRVeFB9NuMJRUYERL50icGp3x1zPxe1Sq6uhiJ2jtP
rneAVHQvNiQ+P3Rg4MAUh3FUEbf/XjYWI+euSUlLZ9Fk2KoMltRTQoLnb58k726mVhwEQZA+c+nh
/qNPEGnBqrYzTczc3SguEHW4KIfP42OqSQgmqBVNuZaLJgdAwEkDXaG1K29NBffH6Yy/qFHRveHr
0gR2gisEqj9VOpQxp0oVfsfUplXvevxDelWes2Q3wdk4tuf6nyB4dvKqRr4qUZEPbfIM8cNTHfr/
W9VPyo5Z67JY1txey1eeUrUtfkIznWFCpqpS7u+0P6aYpasipUOnuTw7y6xhWw+c3RnXDvSiqyv6
IfDkI/9n8Hor1a8sCHeT7JK+RZkOgYrcWpBhvYXm0Th2aRnH/5AOHWwfxgR/TKxUauiBEBP2vYN7
YRCNoXM1BYdoj24uClAnVZnM8lhlIyoqWr9QU0va4HXfGvBz3p1iqZeZyKXp0RH/SRakScmvzfmU
yLH46pYdW3UXUnnAoEmqeOojoZA5KaRfWG5Wuh/KKpycbuCK2qKVXDcNd019KuBieSPpj4oJUmNi
KVwW3MI6O5wVltjzRKa7BcCyE6p/IeVukkPctQzvuJCWCBbCd29VkKCHBvrqrYuYdWZo0ObFLy2l
JP71dNiL36JUEAna9iS4jFExBRSafN46nndyJUehq8WjfYFB5vo5xP1y0i2fe0o2n14DQ/UQd8pH
j6rh7TQi5WqajE2x6mbg4aXlAXoX29T/T/5+vKmZ1RBjfeYEEga9eK9aen8vXymgGVQLb07E5yjQ
HZk4VvoP0XWyVWWA8Lkw8rc0t1YtPdYt4ak1GvIRzuOhltRQ2hgOaZmla9cWUGLWtLI4rCwANI88
MDyFj1LrP+WN3p8yXTi7mlN61Lcoc+xAz7sJ5RpSFMFNene4w89wqkAsKUfATICT9eyFCy8VAQl+
om3Ei9qW892QfvrObyqSwJKo3tbhU2ExkDnCHFMSQqsPbouTWVR4US8BLFo2fgS+FCa1OwPG1pYG
Oei8ZH7NyVWAD/isAnNCiqyiN/nepE6FIYhG/zDRY2mugGtyoPLHyhHNTxG2PdA0cvnf1DK5rUWn
ZVpGr0MoxtIESiYkviYiPFEsm7lvOeMDgF5Cbw9Aq9U3PHV8n2YlVMjvNyoaH+SwL5yZCb8seCNv
GuulPoN60o1lAgGh49QSrsSbzkWrsxxGbomkX3Onm1fPvhR0P0pvafk3EotJrVejnYs8VOvi3vcc
R0KFYSCav2ApbykjPPb0RUY+YN4W/AhL2s2daCubaecTka8nXW7B9A1OCoTSt4JI+DsUjozYhaa3
s+8XWXAvZ2XeEhjifMb0C2PpfmK5s2vos+Rg3JqCewbtK3S5zfGpLfpHa5UYfEs1gASbsHUtVUQp
CViuEaytgVlodzlLEEXMB4gkimpJZGPrIAo0Y0Uxtx2BmFdz6oAZjkEmyjKcpFbdzFHQf48sr+SH
l5aaJn6KK80n2YPT2mPGqW1ccL2jTliiR0uuQ4oSUnKpmOkoHObn0eXTAfsAIIvmnnnwiti+EDSl
5B46uAfLHJs6+MpEkkAMOAPIcO3BrDAVRBU7+acYfc07KjthM7C+R8SOhtSR8oxFqFmDuLAxJVlZ
5IKRnYJKbTZxXrBJ/4r+FsHjRb43OAc4SFABbi9ypluSie0aFQtnqLenBg1L/gdguxmbLYL5ETqA
eviWTsn+ZE42leb6PU6Dx4im7WzfIb9wWBENJx70EUM8enErCzw7SrATqW6SkHL9FJECUWdmpWZT
d9n4++smSiq/bMh7axXw2q+6lZZePMWqBesAxf1zSXw0ZY90YJKKK8yZg9JFfUOyDdGMSRfnFAib
NPK4sHdm7c26ohlIbOPrUclEgqjmNoCKwv+NCUeNx4E/xOmeoaLT7IolTigbufEF+wIzNqEVZsSd
1x9rGDJrAr9Ou9m0Y6osivmxxEat6ekJjofORoG7a7JPfyHNogEdYasWByPiQU0G6Tp2fZoeabc0
yUGessVJqZIJT0COOdkaFLwcAJr47hfixb8lFpJL/ha4VdWhMAWN6fmd8DgE3Tx0gVLhLSQ8l33j
ztxFs7bTH5RrOR+FETgz5PAnEUO+Rh1IC27u8rLJryrm3SCqy7IWtBvPPviexaqDc4U4A6lMCBY8
zZIgVp6oyP0Qp0/U3GyAJizgEi6UNwnNl0R3jJZh3fkaRj0bWsuBfhxuZk83hqBlOJG5weDpI6ds
J8HQLpeUI6VQ8i0DDq4VKoVaadV2ukoIfTDBm6fTU2fnF93LC4zeDyNardp6U5Sd2rYNacPLpplp
zO9Znhfidmb92E0D5D66YTK8x8kcMrc4XGPCvI2dxouH0rh6UUtEy4LNpYyvOnph0PYK4bhfZnAT
vIS9RCjST2Cx/Hx5qDmMXaM+vp6TMAPn14Ywk3xQ+qHjC102SO0Xg9TH4qAJ6mxKaLU/mPJJfHai
8/W79xASpUd4irRUEXw+w7bdq8v2mO+8e8RXk5ZVx3m/2w6+jbG5mX517gcN8QfvSf5uAAfn7eun
bCVUN2fCQAgePW710/SfpM7J9iPu80nz6/DsDOCLhC5uC5Dz8r/tSD2va3BOpyp+LU0486Y13KjG
Hm23g3FZhSvw+opyTZluJMGpMUEQB5aGES+6D7mhp8EsL5RbmqRPPT4ArTKtkCHsnZSn3uofPkTP
3h+Bxx9GzYGfJxuVGkrpFEmWAoJBJfRHpJY3r8S2TJjzkrsBvCIaQIcKE6tRHt3dSQ4tIatBKRM+
O70Yy5HqSmXgyz2NOHeQvtvxlVH7GfNRcXtOIj5m5vTTce0zOwHq9Ju/TjzmuAR7Gbx7qnlJuPQI
Hfu/QbIdlyZyZ5I8nIZO2cCJHleuHAEQcpioADa+oifOdmabunED/PNg76QCBNqzbKhmMEC1ViYu
xovNCAZ+pY9xxVHV30ERVaMnftQfa8uy/T/9i7q1O4tVkThizbVRoAiIR6swzfHOuiJRxFNInu5h
RIM+N2gGBOINUqtAATAE6P72BwCwmnR84u2BWnz9aiC0/zgRzQK+IMLs1mWahNHTUuiDGRfRMM50
zrdjgywTCJdaG9yqiGv3+i8S7KEfFqWxCv1IoP42r5K/4Xm2bNV5/PhuZIi455d0brd0fyeeCzeY
mS15VA8gMND4MKhhhOBsONCVtEF6tS1XWeioLZWFMjdX7B6ufG6rPaIZ8Rzo7UsX9RYZfjAOcI/D
IGx2yqRdIibFvx7tmkzxEGosbP7BArXe68fywVGQNLbPU4DGcYIY/XMAmH033QWRBPjZKlwt4mkh
ttFOFYiYpUGiyjydcbWEy9351EnsJWbok5Sc5SZ7OL1K+5OpE+xBCTsP1fVukzBkJIqNvv3Oa78q
DQq+y0SGbyHuFWSYhYCWUkC1FSE2KdyTnTxnixGFouXrQ7qYX1ceYfmOp1ZSLORWljlq0imATDDC
zltbIFU2rgAAV5tN1+AbwxzpWr+2/lRMTcIS3rKgkTwOsVkckBkmbv5TjD0ARDRSHNOg9rGQ1M/g
MRDMYefTUjWdO++5LX2GuMha62uK228NCJJgm4EVcpPGsM7iAFR4Y79pvMQ+fH4uYH8FRM8NFwDB
NMD/KDzeoxDSRXwvZfZGlNIJom8NYdtdnA+BRtiiBiv6TIPas5RrQ3YJdw0ULKM2kCJS+TEkCheJ
DfPx7GKB/EhrUrFHuQ+YcNGsvIM7hB2ySA5LIDk9TjwGK0ak5eVvc/wpHo5EEoNzEpwJwwV5M0Cj
bndmED1/J6vj9DH2IZx2YRLnYRpq+huqe7e/X8vXjbmXFmXl5IM+jKpMxEeQULVmqPqKaxlHlJvb
/D922EtyOJixwZItpkl7B9MZyU2w5ANL6AXXP6vB6hUhwjB2sGrFfmOhkCOuMtC66GLFsJxkfqB1
pfZ+JgotbCPL5RLulUXuhM2pluMO/kyNxVVFR/ircc0YDlnbgQlHe2u76teVGatw1loGAqVcbHc0
Q5PfVYRmCdJgVvlqxH68VAha03KpdizAB13lreWaa71pt67oofCCyw4lqY8p5XTc9VlShOQyRf2F
lBupbOERsN3ArESQK9AsCBsfDNMXDL4GLKPU7E07w0CbqYxpP4dT0/ujkKM5IvK0nDi7xbxRsoCN
C/oJsr7H9Y1lNWhXP7WUro85oBkV6hNDAMVwzzAjG6a7Q/iJ2s1sFZOJjEpalspB28pSpRYrKjn2
vT/oOoj2Gwrq1BBBEy9mbGs2DUxWRa2whg0FYQMnoqJdGtSCU0PIgVTj4fTmr6ixCc2LtkQhS5Ph
RS313ItoCEV1scY2iPkYWojT/2fjznt5Buh0PzAHrh2T6DK7DZYhwXiXK10T7L4h4BMCeGc8Xpzh
9oTua25qyyajGRysyJPdoN9Co349Xgs0FmtcpfsJMmIFBtDNdGK9puOEWlLiJqOj8DC/3EAwNNw1
5DBj6/SXIiwNsrIs+RpOOQQx9YFvdIkKpH99x9I3awqKSvkkDo1LJ5/batZHtFgbToVku8V4hqJL
wNil8NTdQk7upDgIAYI5klAJoP0A9UCeKzoFE4NGJPFXvvH+ejifKUk+DtU1H/FDJXMQvZFig4OB
x4dTpo5k/M7Ktl8dJAWEL8P+CuJ+PhxBk+HKiu6DHPWXYefi64WTvGf+BPr4lKhG6ob2fc714Vf7
0xDZby1j4O16gaC5yM9qxbdejf/vR+QjI8/2axml6rFh8djsFGHpiM4nqn8lvgM+fR16Fs3vw8iL
TD90cmA283VPIw6USnAw9fCBbJ4/VOfFHg0HRowTNWXH+NNy4Rb8Ou1Dvrtf9D6oBGR2uQx3Yl9A
rfk29c211Z2V0WQfQ5nUewpjxaIVZPpjqm469N5l9IVncC1cdJDifz+iE0nJc4cvBKmwdo1liQf0
6A/dulE3tw/I9Wdlcda6RJnhvA33sK7wzX33W2X7k5UdT5NO9Slp1yi5tGoKvPS9Su35FhtR5ydO
02n82qg0H8srnd3xGI8FOU/oJfqry9XpxyM9d8pSFsA3PA4FOQ4g8KOeQ9RwALj0dN1WF6UH6TO8
oxxD58ZF092V7FgHQgnatBnKFt5td/YuKOd7t9IbelU7byN2pOUh5orxTeHM90MgqdS/+IWQ6Ng4
Km/YB2v6Y/dDxxIlVTxC2pOvsnDr8dBxnVQtUXXLS3iAGIe9B7wAlJZKAlUnIfozuRRI660vi0WP
KRBhNS9lB3rJRQ1LEO1ZjWQ2n5BkwcBjvHhoqerX1XUK6gezIi0nhxffmCjMuNyCCzn8JtX1WbG7
SbTkzntbbWj52eXn9FIZ8G+zZ5Ra/BFjZHfjd6GN27wMXWjjwAmAZfyxoQffUH7vSM8Qs7BjQDJK
1RTeG5PCKSp0qbK/sot1alU9iny2fpjCiLCCoH9qXJglnThJq8W9N/6K6CrjpaNQKgqAHhK8SJ7e
ZC3YGx8O9jx2B6WZfguTWszApjII2VUacB3PQEAJCR8mvhClnVZDJJCOdilgrnDq9M/V7GN1KqAx
HAT/X01e/xrERWWGDpWhzwOEBH9Kw/vQbfEF8o68uRXXtEvMKFdTMBGPUR09ShQG1ToTjJLE1v5I
RZjm/TptQR1BSgs8vjCiMSx8bX+Yr/u50OtArO6FWLh7WnR3jQR/fyLsl2b16KmNxJQQlIY6fa+I
2KOT/4E0l8XUB0cdwDUUIgtH8lQeThRZuoMBM5TkN0F1LrV8ohA8nX/o86ecoBXNlozxZv4vdnj6
H939OtcXfx7iWye8T+96GG6i7wsy/7i+xWLRu/DVbymRe2GP2XSg1dK7ZyWtmlyVYwX5b/bQBYIx
KlcWeaB/OHdqJLdSNyad66kxEgbTJPce30egTzQ1hc6apZUdh2qvuT+2XOxDFFhL3RxhEE6ivLjV
UFB7+9w2uKLAQzWEL/WgpaodB24jWyox7+iysuyDKIk6eNVGYVTltOdvCBO2c1GeDCdQiTPhxze0
kAEzEaMRTqKLrFUPeotydV1kgWMHlYEIXBVa2esy5guD3IeEtRsKkKkeauKCDQoaPaMGEhjouLTc
hAuV9GfP7B112o69FkT02REtiKe4MAQ/fNJKSs4MTmsbRXNrA9KcuIhsLAUu7iTadhMHhJ1AwPjs
jWrU5rijLBaB9WspPVR7ZpcwhEl7GdU/R8O24NmbXooiBbHcqYj83kWEgYNZF4e6zjnrzvzpwVAI
NIkCa+7QP0sfDJXWVZ7yreqFxI8T54esx1bPpTfGh+WGrbEIBaf7DHsPVWXVVe0OcU+mQaueSo48
MOQWKEU0gPDBVI/xguhDgt9W4ZLkPA0S1sP6k30Iblr7Ze9lIfTAKuzHCnLhLzYjzs+2EtGmtBjn
z0LkDPYGib4/YeinT6J2rmzCe6l6yZr1tNqWoZsU5koeuACk3ZEDVobidXj6km0yssy3FuZ8vISU
vTEKSidrW8KVr8AmxSIpoUcSA1cC9bVX5GsHav5FXOc75wDwX3qMcZHIypzv8HbkS3oHoV2lNIwW
q36E9CAF/Ac6jD/qKrFFAUEOxlOTMsoNhg9ObDE1q/OsynekG6UF6+mgMkLvoxt973b59IDk3mQ9
5G6ejwHQuJoAzP1wzXJ6MlMRU9xmuzhwphTRfXQoReo7c3PB95I7H+No9i3Xrpd96VX4WKEyvIFb
MVE1Rcptp/5PvNez89o9KUPKzc4hzNzDQ+FgXs5Gfi/bU+NXYWws/m53whmmUgHB9gBv6tEv4jan
nll0dOqW5dr8OklfqnNAdfQaGNPvcj5du2SP2tLq+9PvmWwvwDyu15W0oZib6K5gNTbduur9pp08
ro0sI4eVm6igAgZFkCag0FdSkh0IRh4Eo62ZkWh2bNPmhmo9ra061uRhiKL7zqo3rFkyClbvnRli
Ww71yGI4z5Iy5aZ5F2RtgNmbTek73K6B/Zqdfmgwsywulsu3llvpZJvaft0HINZIrTiGh8gd7aiR
YuBiEQjpH9ZXYR7BuxmeL7lBeXKFEgQBkfAS6LkjiH+n4lk2rcxi6wU1T3Dn1yCaJmcYEOXtjpbD
F7dYYSAuEp20PZNYQ+vXdQwNhXsw2k1PMv/dk7c6CZKWsgoLzC4fY8vGcqqrCczyn7Xg7UJEVMsX
rNi00JfAtCI8EM+BENJUilPRlsgBldw6W+oLnmoPSTUu6O8HJM+AHCYiLLY3lQYXkRselxZ+Dbev
+YewlhrEOPg7u2Wje8gXi1u8LB0RlBiq2nJ83jz+dCfthToLKKA0rVIw7jd248wiGmoUGHdnVwwf
6tB2o5kJYTU7LcgkJuB65vJYSO0TaC7eLw6GscFg/TxJ4oGTo/WNY4+oshuwjF7LDYP4jJ72DVMW
4opfahgrV1xIlMPyPePTwodlWmQi59vcFofgCCT3+PMMWTsZNssCK5ZQnhHbIiBCNcNwgBuDfdFT
dzs/TEWgKD9USkJok2/Ws7mnhc1LPhbX+ABVVRKa78dp/CgxKzKG01YMaMATTm3bqH87Rhcmi7+a
9wPy0fVkMzGYiVlo0YB+iQTQMeVmABw9UxVAO3s7GhWs85TcAX1hQ126htXHjnTh1hHxf1K1w8PP
zL4yTY380CckjAg3x4/3kD89WpY28pAEZB8MEoQZxT3GLisJXWOhOLVA6zp/xFExTMpCBnwf5tuv
PkcZq5OI9yQQRRKvZH4OL7Ev45UtK/g2qMydNIoQTV3UZG1+x3l5xLiVIUXghzj3BNjadE6XSSBb
8Sed4FYk7j9D6RqG1AmD04RcLI440sYVmcMOuVY8f4P0Zhh/OA1uaeJ7xGhUXiRer/lpf9J6oU04
mAR4HANNyGNP8B6WsF7AAbXIo+Oaass32BeoQ/4ovJyXirKY/Lj9fge0ek+/I0ChSdZbPDTGLNtX
raPNB4XhleAeqYVw5iaUxncYLLkP1er76xQfIPZE5g7iIm0Uec4JaU7sRDEXLt4bX3QBYmI43Eml
MgwJBNQMfqF6iM3RF+k0a5crxoBJrB8431f0K5uU54HU1lC7+X5zynr4ROnF/VfH6h477vMp14n2
lxXM1km6pCPWN1EbYCEhnd8bcETnOqOoprpkWjcvFTNAEPG09G0oQplF/KYocY3sepVM5GsUWzaK
Ac4DXCDkQLCyuRwDvcj2K4ArNQyb76KiIt0lZuCC6FyvlGKnU+3rg2zNwl9Ztwh4D3HcLubDMTsE
+iZvSErbKlVtkUcDtthOV5T6jUV5b3L4T2FtRouwICH2dhRwSY2T+VPdyZfDQEYbgGvgZ3o0J3hE
j4RoOsDKOrY8J0bgPsqJ96DBJOjZ/QcP2eBgNCtyyVQN9O28YeBGa10KJNqCfDjs8Lm1VrxSRemB
2ruw8uMMnSeP7GYDNcIL9SrfyU+gjUHJebm0EDfeqoYzrIAZ66nXSY7JhzuSJ1HjrR8ANut4lJXy
8lWY7/0ez6yvweIKq8sCSQF9h7ls7KkyFMxxnaJVgZrNtZfPWUAx1zSDj0lIb0URcb4N2n1WrHPV
vAkD4LW9TrwoAANOzdNFza2VDcrlG1PhOLg9nUIH65MG2SfcNlTcgwK3nie9j7Cg00t2uO0Wd0ZZ
TZ4419Fm5DEq27dwJAMEjoeXF+gMX/omnY2AgE5t349FrDWAFMmRZOMlFctoIbVb5Lsq8wxIlyI4
N+6DEwmqtWuPIKlRxXhvVPUfbkQ3qSSs+vrHfbN4EZh7skfmh4L9pynrOWfSUUwqod3TuuN8Q/9N
azYPIx7cDro+omrJq32/aeQ2wnCvL7gnljJD2ZsnmUvfy81kJhKJ45GY3UjJzERvahpS8+GCkPYd
y3pzh/7Jp6FshFLRUZzlxPr/3MvgBb/aJ48bTh8ba/k1KB2lULEr46Sclj+cSOj0E2P1iXQ2CzXy
aD9LIwF2xuaVRr5NAKwZcTxukAJhFXTs7nXPezkwPz14RchmHOxBxbUx4mkq6x5hCvOvTfRpPY5d
qD3uy02jsHB2x9htAm2h4Hk8TAMyEAmMs+Vc15b19pxhWFrnXRYt4HtTGrsnxrpBbpSZebkUtC9n
Md4fICl1gilkAPUBbkOIOValS1eCWGtJ6zc4Bd3rGyR8QnIl/rNG3owI4qV9m504SCyqpGVw+Sqv
YPgPD5Kk16zt++mwG06krDohf2UdaF/V3/YWJQTJESSqk2Yv4RKfgn6WDupWX24NHm9mfcBpP2cF
d3bv7Irzq3IWm6g/ed6lRidg9umwRzPH3Ffna9rNc/HNFoAU//qMB8YYMYQVl+FRtvTK73e7iWZL
7YYw7CwWIJGKynmfuQ9tDTw9Ld9zc+wUe1ZpPrdruhIJ4vbpFQ39SD1lJHgwF/f7JorCrWinRx9E
5e2T8a0nn3uzj0CcOpPMt+9mdmjHKmv4b/d93DWNhk0TBqyY6LIzWEL6dOz6C2hiJTPmSEUoHcE/
INoNSF7epxPM+5JNNG9JrUlnJmWxdeuAHvLSF9q0UcOHxWjEc1Ui+9YRHKyReH16pR7w7oaP5cWF
AsXljLZJ7J6uMMG5Hu81kC5UjXmH8Mf2nVTxGtC2uaLFk7QqXttJWPYw5EZs8vfawVD0OsmnJemB
PCQoa4hPvXRts9AemtURGYIPqEeC7ElNv3cbJ6yi7m2tbyw98eOdm8fD345L0xdIgbR0y/LEAlPW
UG9jDT3tx8yjcOUW4VqKpQAzBsDY7GejIZ9VrrkBA6U56NpbVybzKfqUqV0r+xV/TchoBt7lFwgU
mnIuW2rsBhZ4jLnFMng15Lkgt3gH2WrGEfrspSGkaV372ocJk7ow2A5nToWzKcp3WTvGSVV+j0Ii
xSxh1o7sI1qOTVBIpRk8yiPjwewYmC1kLZt7GUtgjtDSeuKGgw9TunuV1xOFwuW+HaGfQ9r1x3Em
eCWHe3BYJsCqAZ4i9pX70dk8oR7wSo/6v8WJlv1tZAzvJel3Q5sTqZsp+2YFoMcpKKM+WVixZ5No
D9yHp45v4YSH7y5ZWHZt/TwCndS7FLIiOBgtzhoTuqwr2tWFySCYNYIGRqsd8HT/4kqIQKmeggyu
zbg9+zTSAcwkynDhzv5Euk1o6DTN5GDgk7VMzG6KQaegDkYs8C7xuNw3fszRJinut7yWlPKTVCn4
TyHthxqEji6YEKNl4Mleg0iN55SI3qHNNJvf2GHtoyb0r1bh8e/gk3FzqtCoWswO6eZIbT7hY31O
FxmQgAeG0vnDi1gmxb9KbMEWxwgmDyquvc5w96Ediq0U5qg97WuvO/eThzIyxkh/i0/41R/gr0vb
ImanOM+vsuvfAx3d3oQZw8WJYCCfBex8OJ8URB/R5J/vHkhBuPV4rlFdgZmj1z11+xfGyN6/Q1ZP
F4UWYJ0aSJDseKX/MIIEQ77IAvV6PGzTbkcErZec9zbg0O8ZMK2xu+CujrTuvd68dphdtfH070Jw
bYzZ2eqdBpDXGjLB1YCmGdUXaWYS9x9wjE5q0HgEEeAzp4NU0twEAL57+EAvdGcFySZgg5fwlfK5
aud9VaH1uC8wv7+Jf88iRJbbC5QcZpOPYkAmgonm0k97HgC4ks/LHGLYt/J6ChgFbtwIujHB5Kmg
ECrnK9ffzDtKo1jBz6NDMZQOFDjwbjThDN5poaWy2tK49RYnsxugDaLV+yCOfHispLh7CtqHqGiC
UAFk+yv015rqi0ZM+4Wggqe4kyJzwshYAUuLyGyaLUzgXRuiNDRW/vj3QfsVFTLgd29xcNf/9msn
8NH00qlRJUBo2JwbQEm1kGHtBMRAbFejXodEcMoGE0Ys3XEBM2ZVpPOi6yTZxGcse5w/o7Tgvh0f
gzeCcFL/CTKNGTP0xD18wwbKdouK3TBdmtdZTqough21UDXS271ME/1XtIfEVmFiuc1tmTB8cYhB
IK8HCAN65F1YVpH760FikZ7BRf7vjYGvct8TWTgeCYP87SUI62CnAF5Bl46Y68ZCEtjl4oPWVSi0
Yp/Hhi9mjSObUZL4wNcJ6aSOSiwS11c8eTDvUHDahnmmGKmWw3bVZz7uB3yEbjfvuSD3Mchh+O9b
Nl2b8WAbET85FHjKSUxaaWPNgYR5mARmQknSCwRCASURZDD1L/L+KGnA3NdLGzDgzxHR7H2lieJa
NwtTKNP7Iq8HAAXBkIZbeNUm+XqsCEPkMyj6C5e276Afc2Z5Ex1Teg2PdoxsDqlV/YPPgOXxqbEO
brUbQs74R0x2XApq+XbBHATY9S0SI+bdsm2mW5bZa9O6Kw3ByCItxc4Zj7jTQhdy+aa8gVqpxiHV
yVvLBBMHSEP49qr+YXXkpXzeG3dXTa5Z2CRaYUfVU71Vy36ypwnUXEVsyFDAJYMAJDxFKL4JB6Rq
sbAmHGH1YeWpvjZFIUDs8kvQIkV+1ks+0S2hqYvGzUCZe3gR+She4HkdJ5y30GC49mgDVNCh8DRY
bcPgDtsGxXCaicor7k1/N0APJht7cHnAc6Hu2D03wn1eNWU9+70nitM+7K08+0oZMVNlMLoUrrCP
//CFUUdZmgYhJEN77/HXD7hK9CdfW2Ur2H9Ny28+FTVQUIYDOxy4Z5cA8CPBLJcqpmopW3eeqe0/
m880Z24v1l7IQ+/b3SN0LfQbgRbDiN2aHLApxvywDOxuq4ZXLMpwqLZ+qQiUaqBLr9VxAnhlAbBE
VfftvMi1i2uVOU4qbuYH7aN86Jmxxon5eMFaZeU8vXhNYqJV991ViXbCpEcP2AAcl583hz+KwCF8
5ppYwAY85CkQ80nQgjy5cARoX/sXgXyf0agm/9IVVP0QKP1tHOKd80HWsy1+1BBb15z5HEW3jJ3w
NhcBz99kdIXMrfLq6v3Ynhl5f3i+014pcjcoLkpWb9qg24n9kWPfJzCOlht8B/HoMJlOMcJxmYGp
yLs8Ui2CAEciwZQpA6eSfm2/IORe4/9E4d7UjeO80bLpOcTCHr/yzAHF/M92oJvRbgHbR2F65oqr
nqJ6ocP/C01kCKy1scBGMXti9zp2TVjIYBDzkTORLrRPmeb9UAj9x4lv1uH0RA+n1xUnWCN/H7tO
9MrfqolI3KCxPNd+7Wg8mIlrRhB9ri5/9HA6yAvucWSA4g9IwO5y0104kwA/jPjcirZMZ546u7cp
jHsP29yWcj5LfhC+um4mgfgVUJKmVHFPusPXEzOqY49v4lh4hKWoEgfjQlxOmpsEKwU6v8nT8jA0
cDWMf1rLXAa8kijHEKUW0zF8yf0m35N5wlfvGF7PA1E1o+Ufg3U97UQA90VF2saHuMftwOt4Fpqc
qScLACe1M0/tvAQ7slF0XqiUenZ2OdyW92AVFhLVOmhg4hXRpEs4ZcgZS+YAsMnPeeoNYRZT7JUl
25dLNAs3l22A3Qvw44rvH4XZuSzd8SAEu+uZOF9vCs56KdV/Fu7cbe6vGZnh8rl0vdcQiaY+1aZy
qBZ84avgMlENLXOSu0otOTsQ572mZFdQp89t6DrW7uv0xLfaE8Jc0lublDcUguu1fKc1Cz41k2k7
8eLhMFh1QLWgo7o8RVIH8cVcTA0t3PUvTKODK9bOYW4EsK4dGA7bOAj4MCCnMDR6dniv1Yg+eT+T
UuFs7Ta6XUKDczn5ckouzFFl6FcBOmWa/RcD8keYkQaZHkxwnwbrAj+23faRK7EHp7eXhc2gGMSF
OOQC4lhdFe92XGC4S8/3J9MWVT5KnohrUuKBfR78BoE4jokkp5lCyD3kOvpNnVHZB4VSLedKvjkM
mAAYPyiONs4v8O71wvy388bZ2OcstLVJyJmd/afA6VHeS3RmTvkMgqAFI5KceqJNqD40ijND3TQh
BqyEnDV8nv1O3vaZFnOA4xIRcbVCBw1bOezj8cooDB6gjiNvbAs2P5sofP/lCuJ/FM7HMEMSo7sC
ZBXiDyGVUVLJdhOnhctOu2aCrQ47vS1dI5BqVRepgcK8zKQZMgMeJ9x2WXk/PMi+jAdFo7/tU0ij
3h0Eq80/oahKFK3+Ik30lGvf79tdj+Ziv3hMZQfU+zMgyv+Zjqq3axl4rlsIrFECFcOWVtB5oLry
TSabezYRW9TmxBhOwyRZ+QCBOKDqLcQq/3z548MknC6xQ0Sxl9CvAvEslUcDDFlbcjo1B8/Yiwq/
RiksTkE63h172B8mAVm0H72Wr//OcJKMCz0T3ozrKOmR9ei/dRhmpSKjsnq538JlBhIB63q8bJYs
R3YlaOJ3+tFgjfc9qn6I6VjZ9gTaMwHHVXwdfGRxVGP3Z/xd9Bl4vIMZbD9GUKqbFb6RB4lmgWKI
qm/HNjZa4dU4uhpchi/xyhF68kB0wYXniMVb3a9ayP7cLtH/y9p3S0+gZu0EmCYRtJVGVICmD0R/
WPrxDJsn23ZbG4fP4txMla8qRx/qYJnLnKr7RPa2fEcN7sKZLTI0cBWNseEDGjR0glQK2a+vk7Yc
uybUAT9C7XilQo43IG86++x+xScW74KfN9dMVX/5cdoVp0MV3hCyqWF2TbvwiGOc8+OGm85rj+gT
pHf0YV2o9cFcd9h6svtbu5I9YdARL047zCZFqEtnAAI7tv9/waRjWuDit9MQScfhcl1zbi4A64aO
wXTNTRALim/TtVaJURrqFzJE/sbnngifeFp2VwIwXahSSO4kpMg9+835dCEQRNJQJpLK74p7m1fi
hJIlz9+smyLaGXcyzRk+Uz5zhh3gAC6Zc1PJ6yjQJf5s0OaZu7t+MTF+n0/Faoxm8cjBFDNJzK1z
YtY3TeUk3p960J8BJB3XlyCk37OrTI0CvdLdZOqgwHNJFC1HC3KpjIQsMv5TK9cIaCS3JYFvSkBL
/0+b5oaKZqlfoZQVkYwni4Nl5CqTFl5StjERcdn/HIJu5acbU1Na6b88oMpSHJk1YmbrG8mHSm3q
BTMtTp3hepmj4Rct0c+TPEHiGXnWCXTXUgvucPhzwzJ7c67SFMchkfVrsk+vwBebDEKV/Wsnxmlm
sHTAwqxf7XfzOBgShGFujWNl2XYYpch2EcOItbZLM8gmNM8LhJlSEt/ZnsASnQwaZPM1sPTeIY2j
CKMKzzHl1mf27JfcL6p9ortCgvoJzG+r6rDSaR/0jI6nugcPt6kVqwZ6RHXNCKZsQV00bhVzqUoG
CC8wkoeBQLXsz+YIg8dLYfp6hcn6R6+FXoS7snHORYTRGzLT7BWKkJVRjceJS7R/ynvccqDQ95w8
V+8K+3LGVGu0eXgM2iQ0bEt6GVwbuXgvt22EdSI1I9PfRfQHEj3MBPj3KwygUZdowM3pru5xrsYp
Qm0z5Ss3+brOPKBhkH+aZ4elusLqmubx5Y5rOaKFaMt1pLaeI9F0dPKU6kRNkwgU7DBsBJo9Dx+W
+b9qxsvZt4rFI/5gK9zUCigo6W5TbGWmMyZdDohPk3Yo9X0uQzjNvkSHQmWo+SD2Sq9iELGrzH5N
PTajhzBE50VoIvdy6a5E9XH5IycPZzQBuJaiKwVtcbi8wViXUiYZqjIxeO/uUYvboth9MkZGIWLX
HcRr2xrFX10dtmuqg9uruzEimSN3PW7DP7hmA8RX3d7naN1vf2D1BSAMsc27suuD+hyIIcLbkj5j
/OQNdE4Nr+rWenjyqep0vqz2iUhcvzuKQOhuR/eh5BIo0BVx2kfqTnGZwWSeHcaqaikvcbswI343
TPzyHq0Kncv6hiabVISaYrG1w+tf1nh8n15VZCzxNEbgN+x4OsoUmJQi2l1aWTtmSYQMgE4p9Oco
zuhoTV5/rPaktwsnlUDPak4uqzaHUBImOE/y2krJemB8CWUcSLW554T3qcmoMIJXbnKGSo8Uw6CP
qZDG4wZJHj/VacEZTi0tIXejKlnR9raHYQXgYUSZzKEzCnurT/5wm2Hs/KOBIwkYaozz7cv/8lM0
cAZ0FlN8ZfoCJm+zdzyUqHBH/I3BccHNNQDrdlBGyE6GicSE80aGa17+fJ7fWe5bOko4yA4tx9lO
oF3X4FmMRn7JdtHYmoEK64O/qOxdH/t2ZPZzJ9Ex0OioTYw6EBxngXsTy6AS8X9+MmSXLgAbvPj/
uEYpPcMSU+OHknMZbBv8WGGpYILVyqqEziuSJi+rF2Iv15j7M3SkZ9rCTsVm/TEunZaEcOlyLejc
3OwnueAfxsnCRZwJk5Yke9oTIzbMB0PdEUaGSUVgMsVUouMyABOeUe34KQHWVlD7IGn3MlhYK5Eo
78ZGcx+KurY+ApaxEWFAbBpZOjuqRQnD0i4UmcNXS0W/80IBeRQt1R6okOD5fwLuqUhmHSW+n7Pm
hFBg4pUrQK1yh7FdljFBkAyNZlwltxP8HpfcJgmsmqBuiJQiGKZgNN+wpWjDpHQtIi6YiieYahPw
Rmi5oHjCzQeG6W1todOxcMy7bJn/qq2YZLUkIliotvAB18Yr05vPebqiSoD0yLg4zkZ5ItRaYnbh
Ek4nLTigygiUxujpJoy2wJxu1mU2H4+7Ysxm6gzAcEspbEHZgi4h6bM03xSjxBdQoV9FKwnzKKWj
4L+gerdHcBBFv8zrL3m9fAXN5R9N/D4oPXPLtFungl7ZLCRJIqb/KHiCyWebUjvMZjgepoKETwl7
ojjR4bhzgDfMFafluOcM4J44UoQqIUoDvZ9Vbfh28mU7jeN3rBDqE3j1gQSPOuCx+w9G8d+zrkha
J2Q33LPkI3cN3JZ98hPZUwFV1MpvarGvX6jIdQWH2SL2JY8Jp+95LrQpQW77Lyc41s+tfPoLqrh6
OWqavhkhyLO8NUWT3lDfbaMvv1Ny1YG7kfUtQYU1vsWLSUADOt6ZK3ckN/A/nQDj9zCGRg6b59GF
IG/Xxee1hm+I+QkbXaPUBGXv7JiEGIj6Udydfd0rp8+9oVTKzo7UB9dwG9VUqblE8rZ1KnhxepzP
x5aHpKqzalUa50CcVDtwcyIRCiD/voQnoFl/KX7ix7jGFFlvJFSfe6QABtivDjPkErMmSbqmHE3m
AxHcXyuB7FQJ41IapHW5Z0n71IA0EUWKrDDvFMopQmotFa6ROXvLzVNwEp6T4KqGs+WWZghwWsSd
oknAAfWIPSgcyqdxnH0RjqjGexNTGibK9kS8C4WzQs8T1eB8gWjr1ouJRCHcMjOVJTDqaNMrJ/D4
XMTLTKMA0g0oZzW7zzIpkUfeFx0NivPyX2Q1ty1JdL4vCiW4PZsPOBf1U8f8ObvyHv3EWu3JW7UU
LAGChQ4uKEUyZMLwsiuA5ULuQE4g22a5SVyFresANtfiCSSJlThQDVoFnD6i/fh1kyet32WhPCHn
5PKWW8e2qTA4rb6aCN4010OCoGGGsRHsncvDTMiUwnkxpUQS3g+jkjl2dXsrWW8Brp6dZTZ0OdPs
L8QU+kSx2qPQQqvDL4dBcJPlk+IqOqCeS8gTbtjNndpqPbTVffaxuh2wCfqmLmgjctjHMoinVrHC
FYEKVTeMb5K09N7khFrA7qCtlFau+sCRTcM+VRxk+JqAsi7airsSxXIkCHO5wNpruqia1HqTiOus
x7c7WKmMmklVLZzW/QK37UA/AgxDBIVvqkNTG6YdBKamqaFjmK2LxkOT/FR73kPNnRktew3sNqPi
uNK2CbScmbZQzJIC5OWbDKiw7nM5sONpbaCaXj7wgp1a5KTqfc33ZWLAqkEUIT3vjcSkEBla8t2W
X3KPq7iYUTIeQxiBGiKhoKbGo5nBpSrzCg/C7rNfXrjaqmU4WGroTX9DKJ2FkrzByRGxf5ehne7v
UXvKOmQ5u7dkP88KlWAXGeAe5vAFGDPbG1BISVXBQHnoE0yy/Ge5EbRDAgoryNskge2NzxoA1nyu
dVtQLmVhIjIoYtWII7Y0XwhnpYfKrhxrJ1UxLIRcfYhL7rKgx/zIlNV1oh1mcBawtm/YXk4agT7R
6BO6ReP9D9G5Z26h2wlkSOeKm1StpBb599XLATEIhqx6HU5dG9jL5DUmQpetDuKxi3SV3onbRLVS
eeCpfdZ1d9OmcSn/KOWW7wUEInlvuNWZB8ba2Nj99k3bk1+oMjaqDbK7zKkHj6G7Zv+ZjlN1UFLR
FJpXpXnu03NfdabozEyi/hR11KU7MfrDdfBu7jgRLCz3XgdwxDDLMChokK2P3+SmgO7bOgZIN0jl
t/ecUuvU8DhZckvWkXuIqOQQ95XNmI+J0oXGI+1OMhsg/TQmZIKtfT7xVxWQdiPUgW7puwl6+Y7l
8kbf6f1aNQTtcffcZ7mAl1cKTRjGyEM2YgqBRIAOdqqCAdpL4OrTnvRdZcDXY4euGgIoZMt8HgyC
WOqF74dz9eMrjh5VtkERD+AduVwep/YsTjeTQJl/YDolkd/wK26QTuyZOyYzmNfKatyghvW57NV9
5g2gATl7r6X96DhxmeRYdZw6B+AnENR/Wvk3R/r5xoOVZerGK7wcwtnMh2OFP+VmBukE7vFIW6tB
ggQBpkekwKbGNM3SlXNP5d/T3ZfWpoWghuaGYToxDSFMc4hW+JNoCOx0aH7y6vxdMT61RrdkTbt+
7/bsVFKgJw22nh3kfN6d/vmjjyTicpaE3MylawvyVnaRStEvVfpztQlw2HYpaIRsb6PW5uEFNMep
Z9to85l7ZaONCpMg/nzbsp0ng4lyACzvTllKONHN4tKWPDaa0BkhM8iG6RbrTxpWS5pdOCKcBGL+
7+EUpzr8rP/PSoI0GUhrwsrqHpnGR7PfoetdVp/v1+7BMbvggQYH6OPu8DJLRiO4th/9qACHz+A9
0TfGhNiIDu2gU/gRzoazgVwaC0tBmBhdrhkFE/Bm/iKtrH5IrJ9kE3ORXbJSf+ghzB2rqBV7U7tx
xYKwLkS2/jGfOpuPHtIukmJ8e2PbJvX8nA+R3uvFhkK+qD9N//pcpVFITBoL5cyKza7eYU1IgQ2Z
BgPt7sP5shVHKWQNfiIRcxcX4CNszV3TLt99uN5NwgZIXMN/uooE+JTKYMONOaCjyONqZ1VESOlB
+LikQM4m3Rrw7J6B8eSAaEM9CMqzZvDu2o1pC2qJF+wj4544+UC7g1164PmFkqkDuQL+yEiR0NFh
Itl8IScU/Mi1YSALva+R7CpPLkhmt+4M7ZJt2e3yH9lLvX//kzWASMRAj/6fEKgPqSuu7gI+c9Uq
DWNFFNOod97uabztJ5GjZ/erqEkP9e/p5IV8Wuuu4y1eUotW1+h5VIh4inbO/9059d35wY3aPB8A
pyfXXUsj34pWVkldfzo52h2cR9KD/jD697rptU/7VWIdF3W7dB0iMF+uYTpqkBpDROawWyoD7xGT
EdP5GDPj0JkMnWX1vItygwHBTjGlRXIBNhpeCcMFfnEzLj8IFSYDi7vSqNGd81QOz+dwm2nUcVWf
T+t9QOPGOPSs9WXr1TFGOqbYvonOTURHf6JeTCDZYPkkpr8Ygu6cCrOA1E/PNZN5b1Zenq0cFGj0
aNMmCtTbgoOs7T4PG+ryxv+0fOITQOlmlFcsxy3Q9GvztPVaS+ShQUfH7cXn+ezxJ9T5s9Yp9hZk
WBVbA+ifxrigpGhNqE1C3mEMbvVTRoeA47Xex4n2MErYN6JuVe//sCyb1SL63W/d32B46cTmPUgj
dYslTmzb/ciYQVdP2Zy2ktlpwK5Z8h6wCTMY7s/TOE8N/Pzep9OJUibzbcYLh1O93WUcNy/PKc1b
KPAU0LSSpndz0EJw6yYAizr8fZNIRvivGZLNq4ueJB5d7JyLGzt/JPtGOqJ60KOmGxYAgCTrOK0e
+oAKxFbZKPMXdpDv95k2ywrI1bRVnfrDzKO5wsvWAVFI56ypiT8rmVM3JDM6+3JMxFvKqbt/vTxg
PpERDsFnJp9qiYYnyiLtgJEJ2UEgyL1oMSwkGD1G8YGNO1rt0JF4Rm9Ghtfjag/q+/oYCW11LqIa
OC6DhAGe3Gs4+2RwzcCCDEm3GQqZ4Bbjg/lQqtnat2tc5VYrrJ1Q30PqeLjqaz03ZvbOj3oGXPMG
PqHfjPAK41thfy1PGumqlo33qc2J/pKMh9VMZquCtAhWaro0n1FCg9ybVPO4Ctofo/VokThL3mk+
HBIsnTmGVMNhJL3bZM0E05W0G8VyfEBShFfcHcCqVoJdIKl1Z/ge4fVtm5HIIK4UxkqOQwlpgBFo
j+pSBVVt5S18R8hkU3EERYQCawc/2zcEd4/ThVWd++qDmtYEKb62j8UziZn8+BhKuHva+hQf6KEh
XsJQ723oncsrO4XWRInMaly6CfPeqHzj65aYjidQIY7dc5dzM5YC/sR9qJ2wJLauy/sOk1fx9K/K
KaZiIcGeY5OvoDxogeRCTCu/8JPiN+LX/ZQAzmLEZ/L8FxUd/MMWDPPSo2V5iQlXsfX1EB/XUT1H
sM+XQLAzkh4QPkEg4I9DRM4ETRlnBKLYLMArvdLOCqrMZUrA5eAg03HUGch4rQraj8hTND+jbF3M
VRtMe8M6OP9Ix2ljIMHxtuNWmEf9vUy8fSACLPS3w0rKjRxfEIWxzEftj65wqfO+ijX+GJ/OuRRM
DcvSemxXk25xj2K+TjOT3cjor63Hqquy0um46ucXwBxiv9/bWnp/14s6KKtG9WtIxiVCV1CfxUTD
SbXQjOCERGjCoaUfZxQ+1vEHRLTFm86SQJ7/tnv05NNLSMuWfU6aRGCCQJmTuxxFZREVItjzwOpi
xiZkpzsYeGQehh5v4CrAJvENUIKfqNsN1/ResicbwEiYJhKBJDK+Q8Ou1BOI1myNe+qWZ56+bPd4
9+e7E+ipd5/EBIgE8yNIvdg9/rNGa8WATOoaIci59ziqDODW3ie5wyMDJj2Ujz9ceVsvkIUpC9Bf
bpABxQHB3jFCbCdgY4wcxx8BKPRG4AXyiWP6KHsIz5mtSzej4BvQdw68wpqVXRUmrrmbdFT66dOs
EZC4tvenwm2SNSY2JksfB2okYTwOhO1D3av6n+Un9LXSXpLu5FMPXiCV4R/jExMEpLp5idjycfsx
RwPv4ZO/ORymfWJWtgWsZv8VIDQoUDw/3R99rrh7+3KhSdlH/mJmLY+Kk3byoDVhRvFUnAuclbrL
jSTSktEK1lI5/hnVr1ifbiCCu5k2ky7SO+kZ/rTNTh2BaQbinEEglLv9T84czNCRg+yXAScccuF8
w906F7Esnw0lA6qMmYLcFzu8dZXm6B0fJCTOpFK3bgn0qA5nX354KEfLZbNRW3MdoGoCje/jRWPx
xQaEEMkPESIslk4pov7ovOTyPpYlqcKegb36Qk1F92IBFPkKsWSiHdu63qQ3GPuRHwYF4+9PkhFu
/qBlMTDm2X5KNpLgaLUVjLAuwKh+wK8lmPDXIukWhWVlKai5T3sw+aQAzGQROy9MMtlTPouayoT/
hxcwD+uXfCRCYDBeuXTDFKGwxvPwKIAZcnZd5nZUts/OcFm7Mro8Qf2GM6dtWAyfv58CnI6rfzoz
J6mqJyiWhFIYfzAbPK70/d1A6he/InNw4zCfIXhVA6AwdKwBqZsEGYK9Tx1f4fsE0K2deqMPpHmx
vZrZ0zxQxbCQeNjLatxy+xAaFk2hFDcoZnz6oX8/I8RSDiocSTvKA4eP5Vm0262IDMQAtcN+2b8K
7t9YMS106FPSyT7ci1XaCfogyKBxYpb020L/72CMVusv+smUN+4hxhOuIgr1424X7/3YtJb0cLRm
rIM5JnUzeVtcnpSkKqnU85F1WhvV0Fuu4WeBh0difJy1nNSvh/NT7A2RpbBXLXaLEnTnMvnCTcxF
WFO7PMTyOISNtzTgQy95v3Ja3ARh2u2tVtCmuwHvEqcT4lTyGN/ut40RgTIhCUMa97j1T6W5eWjg
j181kHoS1kZOIEbTDvh1/5hghdbympKZ1fRZLimJxuUCmHf4sY7zJA5Tk6kJ0Hzck7Vksy6BE5Ig
J93UvECt/jlBmf8b/beUbxuruh+5PlOS59eEIG6uezN3qwGWnHnL3eb7jTjiFlUWQ4juj/dI/4dA
Xn7PB4f2ksQ3NyLTozn6UuTEYiSS9iVd8DoxZ9Z+35r9wEWObzI8N5P/5hd68TN51aoqUCzDLX0w
tCsNJiTKLsbnm12xwvT+X0b3IPwkTllNcprFNo1YV48i67jIBKAHDn631QfBNiaR4XExJSyTAPNF
HWoiTvRwIZrVZawI92vhkhPV2Q97XPxvxMmTvvWCyeV1FHRSsFWf7XPRmZNpoEO/Oio+/xj3UTeo
CiszTJ/FM7pqhhTaMDwSHG+JRETkKil4qUCo9CZDNOOAHq5FaAlppvSFfEQidWIgUaSgvslJZPhV
R226Bj+E24Wa+CqJxdniKUvEFeLUdKIBMgzbPxf23JvkpfasAiULmRm7UDuExCrCMzX/g9NvaJbI
b1mmzEq3ZhhC2fCUO00LLheBYkNXEjSkpygFVbba7Z5lDfPhca9S//7kohhuPNZCd1dgvw8njpN5
yNDwP8WozIwm1BNIwb3O4YqrsTBPKwAGI4Dz9nEcmb7F3SH51NxRoi+nby9+C0QKctK8hdIVJJFX
wmzmZfxkkJLIm13wX+I5f+Ro+loJ3rmn2MOn1mae5olEGsvY6E/xBbnBlIpvdaEdcz5YWCFRD7PL
nXLBkhU4Y4MH1Cwx4XciSnqpHv0avmd3xXDwwv51ua3za3pcA12E8MznVzaYP5RsmDOiAceXZ+uo
aWaUaQjcJd96HaxXaFvq32xgI1BAIlZ80yhsT7P002/nAV98tXA3XDlhAUCN+qBRzL0GUgV7vTSz
+T2B8dBpkV4V4ZN6wN73K1ZF7wUPoOXw8G7DBun0J6uyG+oub44pwLEJd7q4D3aIfodaZ6cgHAgy
5qDMZU3ET/2VEnzLq37q0n07tiioDY2Tnbi0fAUYXe2AY8YSKxelnh6FsbiGrr8fQ7ho3ImrExGL
nil6j3GwZNfyTJGB2uaMgU8qnkFkvnk066CQPBMe67bq4UI0j+zkmH1tZW6TGjQxdBaxRHFS+RG6
DxCm2ROKREYqkkujJaORuld0qX3BDUdP08ALQEOogp9bgeMQyRBEpwN0RFlXR7M4HoefzCewhO5L
UFqMSb7v/65M+xZX0F0CHNoWUGK74zYYTy34mVQ4y6wGgb4RgjJ2K1wZ3ZCjPqkuHM1RnI4Ng72T
2j0HKYfBG1A10qu8TD1ozww1hseAV8UpzvS37RV2nEzHojBzupc8Dn+OIYiovSwQMNuLsXqzn0KZ
OdhgQ3IuaVj8qLJ0tPTdps6tMJupXWCWCHVO9w4N3SY/eo1PTv4G1cADd1hvfxYiwf0fJTxVPVnW
fZx3m0WUfAYDRUvsBzbi7M+o79SnjXCWm3p+S3B6f7tHR2wmWrWfLGWG05kxOmJvUMUwm7CvCVSI
+xscEr4/i5nTeLuVoaYehhBEJwU8D9CKnkKnPqPLx+pihRRa7LFQ1wuJWDpOjeCXR0Mt3mjeG4Zi
0z0Y9HZtFeUhSa8NoE83wo4k/3fjBNz6NXujUeE2yyI83Gpl2P8gLezvfK+AUtVsLqdg7aviV7IE
YKlm2Z2TJNwHCMatEe0DZl3NK/t6oCu8CLA+dLCt2JcdTkp8g9aBAvRSlBg0R/hrbRyKADdiCOtd
qaD8RFPnKRJy3QyP2xR/Z9v9vhhB/w4OPKftPv6txFgaGKCY0xXrLIsolnucNJVcUaJUWm6WwdsN
R24TloWMFQDV+s5xo67YNG/I2Gt9bJdH4Uww4F4X9ygji/1Ypbjw6OLZjkk3VjXP5TCvGaCsJwaD
0AUB84iixMU1/jVBtOi+aHrEIylyT/I3UqK/3WGf7rNMw2hqZtyC9XQXw/idXAzdwEvMsHm6pqBM
snB0XLuNXWDLHYs4e/Ooc2PuzphcNJMQz9Ga2u0roycm0f/bMB0hBqk2ey44rpUsY3Eg9aTMc091
ZFQXrhmbxnejLSkUCrCb8MhB9+1BixC0/i19/I1kssgKfAkN9s6seIm0do8poC66MSfQd2YYeRNP
PsoOeDtCleTvMzLRUbh3CANxybRL0SrR30eY34ltKAN3a8DwPH0yfh5lLlNeQQVazerVeoqgUvaV
UDNk7ik7lBJBLQAkqJSDVdC/A0fCVDeQJckHcE06iGn8MuAVmF0pH82OYtHrXpnCObyBqYIzq8yN
WZFSNDU/z7Kvhe0V6z3nZ6484nUnBR+AZ2Yya+qBZbTM+G7QCkHpw8calimx6OsghUljpDGl94ah
NiKIjM9qzLXoVMtZleKSmhtaw07yw8TsmQqXrUmu4GYC5H4mEjwyE5M+Gfz+6zHW6SfoxVJHYIZN
VzPYuN9RQova3dkE7rT8lE6LeQDxnrR4PotEbyei2lf3wXgmgYlneqtDt0h5icxAFOL+2b9xA8Y4
lF+jHIEuxiPYWhbTiVZC7p1ZRASi8N3/4xXAMZh0DiDdMrZLEyMsVywjtzIWQDDkgw4JuuwURpey
SrKnYwegNggGhpe7vALWOe/2IJ2aDYHG19Ypg+n7nhO8QlT8OTDjlrCDSIH+3oS+YTxH994XNHyc
do/f7QVbCmvqVDH0R6AtrjVab7Tj+KWvTB598KiGvj1VgLxvj1KWu+MkGXqViM9YPXo8qp1krUfQ
yFlx1quHj2+lSAhYtd3aImvjSrac51n/4FKX8FFI0NAYIAnw4s9NHalC0Dxak+HxMIjjKS+krUv9
dWk1KzYGjxB610D1XWJpIF9nAFBGSF6aFQtTtzVu+iiI5YQfUomFe63mL9IqWzuAFUDv5CONSHw8
tKUu8z/9dBG3I4cTAnZsWCw1sF9uU3atTckZHEvxdLAFhPPjS9ZDt+Qha0PYbOhoNiKszjZl50id
Hm7qi+iiSmSx+4WZguKHEU844c4GmkQ/zHaYzovkOccEmQS62YcNs4zyGd6n8uI6hWFOSZz+raXI
+N6CphFL3vipswU08N3ULkmYSm+b3FTbVKkW1Yi6FOsvY4w1PIq+UncOADA2kOBlxMm5rH+XP6we
6f5Y0pn5vUOTPhudzHkMrai/06Ii+2AX683us6JWZ/MFMu642hEUugePGrvnJLaQtzSVJMtSqozf
tYh7P6Wkl74Zaz5xrM8d5R1d+uVbKBkIAuuxjpJTD6aKMF1GUHOEVM6FM6+MbizQ3a63z/jW9TRJ
XYemRaSVRC0Ui/nyTv5DZnkbj+S1Qkomzhpu5MfuCP2mfhyWUrpgmCU73cU+MWOdO2fr9fpFIjyi
g5fP5mHxEsQxqB1e3CSCGFtiTxDOjkvJmPyfupVWdtLtzLyclI65SHqURzkRC5tWt7FT1i2087XL
WEGYjf0KYUX0AkWDm9SAEh59k8xucn5dPQ3a3xrUcrO0hNj2PQGzNJIn/HQk16fj3cF2g4xWaMIa
7+j0MzEcg8/atqsXmpWkXuaLMmMoslx/H2bv+aaBVcsvGfD4h6CMj3IIubYPyT7NuRpDAGRQlnJu
FpM8xBG2GOeZOGp6rxmn5OabXjH04rLxNrN30X8TDhOJno07bihZkK3b1T0sT3Ma73307GMrxQhV
o7qeaPTVR7cAOljCfSrPHKjVBLZ9jEUms99hvvgMDSZMYN6bYMfzCcBX8B1alJ+O7xZTdtB2t9Jb
131B3V3p5TzL1dkowXpBvw716J7yj5VfwADG7V2GlmhQgjsRpEqb0QhKXDHyzsRJ0Tzox/hAqXZC
6PftLml4l+7xWY8gmbZkoaz4cMvZ8dpB67gpEy4XYWof1kvw2udb3TcDKyZclIVXIhcJS1rZs/aZ
CQm8/io6kdTQIZiu43ieQSPYzb7LN2jKxjoR3TB1j8kykpjD0VYxhDbCSwsut/Vk3lHTvSvRctjn
fP5lmq+mw+mSqVQfWlJc16iiPbK3V/NIVn80c94Qquq9IrfCY5w+zGFVBbG5rUl07e0D7dxBKORj
kL5NhCl/t7twQZzt80BnST2t2h5iwgcjBR+ML267f8tkPZ4+wGmR/5xKbUt2I90qNkCDZPbqrOIf
g0drAXLYXo1BR34I+u1TVEze59XPCcX+CbVWUAVIux0mdAgPSuMui8Qw5Uiz5x0wVzgDzKZsKEBM
mwk9MwiXNFQn0unlLNrB5b3L+nIWkCff3l8bgwwl7hWMueGE3keU/8wDgTiVDePLBmwYyXw0sYVs
DZWi9HUXUCu+s41cSs/7fFxeNxdxb17Z5EQmtufmDZL4jy1k9r5T7E2ukrP0IEA19bJ06r4LLEE0
PnWum4TMjSVp8YjD4KcwtkH/Y4mD2NDL4n7iDPtaW/fZyqdr1bm0DbEticdjj6L15vs/YsFuWRK7
N/UfeRHkofF5m8s0K0pkog/Cvby8K9Ozi01zXsfCxOeRKE9HiUVFY3JBpZFFFo3CPHXTPawn7Wra
65aG215dq1df62CQmHgLWKJhsVUr0lcZPueK7D3yyeM88UhRi3P99ywM1BGSKNHmYIvJ4rg8A7oY
Be8d2+JUK15l/dOL30JIWPVcvch/ujyIjJy1pVS4XYJCgPrf/zHt13ZhVUNyxrsLvV2YjFgjouT6
hfl2+JJt1dnNq0/DMQOKnkBbKH9JDTp2JSslirVPOpEqNvr3PE3XHOTEqQ0+2eWBzSh64Y8Yn9m8
YWfmJdbZKrqINeJBUgAg5bAbr7pXsXYhHKT1mcvol9/eqpVlYYUIxsOG/0WilXTNB6n8OnSjcx+B
vvLqEVB4Kx9oxqHQheNEaJKP/TzBVSil9S+YVOgp/M/N839olCcqdfAfZok1R3f67WShqMuzOYvF
LrTM3bk+x7TVRwMDLLW8z58zO+m9ZqVGHjpbtLbgkye88wcLfk90LlAaDMwhQj914QZXqTRe7KXH
yI4GLGa99vUqgNmcqe2hziGw9vsxuwIKPKLU/mzZMNmhLUoxNaOzmFgIuA+VOumEkert6rwAUzN4
nXbjrU0sFnqg5/GOjDi289oXZQyMVtRJj2xa5HBaXNNDcUvWb+ToT04PudjU9Z6ALg9UnxcaoK5H
8MOpA5UMfXr/4E2cgXIiqg7dRd7ubYjB+Ayy94MZswI8OrQUix6fNZfwu4acbFchzQif0Ghea1GO
vYUqickzp95mpbXQ0nhcznF/gCUx82KP1QCp+tKzHuNQ1XGw4f2vAZn6r8lkqM85IpK3G5CasM3F
3fJAamECh7FJ+U/1KcYxlUhDvi6ZrCANu78Wm7c7gPDyVUvY3CcZKApfp5ROOmjDpQNMw7JZXKKk
cHS8MjWjcZvd92POcmb6dx2SZnwTRGU61AI/VXNdha5dPB3JgOtoqxp+y2vOuF1dWCIBAtFIQ5hl
aevvis1AOWucUYbOH/a6ktfczbFblXq4sfjdfqJ0DilG6T5rDuIY6DQVW1XcoLt25UYxdiEmDYRK
y+THfdrFJot0vTdaQoRSQj/KDKoJ/vE9Xdu4Lmozm/7yJ9bs8exPYU+Eag744ztFBnDB6veEY9oQ
OpDNEKeFVvB7EbLsvOMM8AG4MDNhpnAfYWV97jK6/Yv11gddcp0T/pz+GSwJCdNsCq3VQGnPYAWt
YmBs7uMmmXAEh2Jmi7AG+UD1I4F3EbDp9nPKQZA7EOS5XqiDcXOcnWpocrQ4AMmbuJNmQX7kz3Zq
N/te9L5Sa+pipHSgpQM5w8av8bmMvZnihqLrCWD+e8GpL3FUI0CIWwUfd1ysVNFchnXUViK1fc6E
4vqrcZw2A/4E7NtB49MiEpcYKcjTmxZD9pTOnII/ZOUkXJnpe3fFxJ+RTOg/lCwaeHHL0fL65Pw/
pmQhFw8LQT75BTC24nh8h5Qz6ukNWfu9wOj9nK1Bdfm1mqqcxWOqNShTbcaNO8/KXrgHAo1+0DIY
WeQrHHtCUagydGAIDDkqk8MyPtWv/FYx9HUV1XffhedjMM3l6vp6TZ0ATk5lNWDR12KnQhsxodGe
otbfK+oPRXIe14FBcpLpuC0ujoQlXcnZnORC+oKijAtyMHrqCafTzizvV+C9UTvqJ39mrcbrdUs5
J0O+rgCjAPlW76PM+CxgyDXcrYzA0nCT075nBYZ5Qk8Fq+XGSF45c1FlLIIFQGi6IK4Dw4WkAvwk
FXHyas6H5rbeTcYRoV1WI8zI8EouNiX6MJRjmdPYuNvS0nNh9uzdX61zs9djjkEZZEIYzfQsAeWG
eZmjNBOSolvoIG2YwFssCGHH8UaZ1FMF6oQtLL8DTmvvwqReDqIJkW5pf2QHC9DXYeaCPs1fOOjr
/FYjg7wIpC7x79lT7elgjFddAqMFvg5qXH8TVjnZ5aW72Y7XOrmr5dJG0O6EJrw6TlLn5QktHySA
NCuykibSRflt8klFvYF/pPpGrWtGdLjlkvyazHG3LHZWytys0YSgvOV/SaWbX3MgigN3ztRj+Tv+
My2qxzogEXj0OsAFRFN8VbhkpTJ9huyNe9mdx05MIHhF4r2XPN1aQopubal9b4QjkqK7SUrKkxDG
kCzNE9XrmXcmgAd9vVabe7qK6+aZj+sZAGwILq64XcayK9RPTgHLmiRF44cMdp5vsU5/dqM0/aUH
8R9uH37SvLHNpcdunT46haghsvk+l/Gpi/btBJ0MU1OqXPP4GFNtWin9P0rElZjmWMIeHrcRuYvS
QGBQ1UW++v9HV/CM5F35BsMhLIEI9RYuenG69p3vFBpSx2tE7DPj/EG6TCt0RlWW/WyXUrhp37tu
HOpaNhGI2dU4EWNoYu6SuSoV9QKK2si0nvBe60x69293042qT0yoQ43G537NR6UrwaML+1E3eadB
1L7lpaMrMYHkGxEl+D6686Zf5DbsK/fkBm/j3aMl8WYnl/T2wIdmIgJVH7dyEkzx/IKAKpDXSHm8
rTFhKVvguz45y/ADq7FzJsgisq2zRdvImgv/38zGgicOKtQZQN1HZK1kM/wZXnFgfuqxlEQ6Re7T
ZJMs4gko4yyk38tIA3VwMLJJ82QgNJsu3lkAIWe75nTwkvcsDuPhgAGWzkEpmbb3ElfXhNZa2HSI
MzzGm1x2g9sqTeXAoUD3nZc3WdHSDeVmN2zHaGDjQ9/yWAPauCYVqJBbI6InIByagUK785OW2JDy
Q4dkNO5aZdqC3OyhU/Y5jBh5xHsf15PUO5Cql7a3dTaUlZ+h2+kFJBk/V0f9sAfFMnGIrqdNNs+H
xEW4RJvjeh51T4pQt0n44T0eGlb5gz0nTPnJVFRWM1oeJmrm4WJPkQiwJG8OD7mzOuTxtuiVEv0W
PjrbtIsQC0L0JQPW6Oc//nyuhgEhtYPIQWA666v7v31AYZg9QVHYVIpmoLu0PFzllrVtsnpyxVnI
YaoE24Vc0KTHjTEIqxN5EwOmcR4ascKetSd8MBERnEIxtkkehy9aGnwta6ZBNgL79AdcrONtTLbd
kYp6YBdoBE2CNTdXaJdvf38wBL/SQXk7Jjq+eXzZrom44/zdCOXTaDN2/PLWKtnQ7R9B9eGVFWxA
ycuN0yhm2SgktxgTXixY5PAZ8wG1HkEO9/Umm75SzxGPP905nzQsOhmrxO7k1lRN+PvV7lJwXSaJ
MpGYdL0vsiMKqjbyT5yPTyL9Soh9XxldQUQj+j9VUKDa2umy62tdhF2/F/29lPkzD2CmfRhnKz2F
V4pRKyiUHdZOXQN5/1y1yrhbpwQ5ov6IYV53hOKhb3UI0ragOwTKUYuoqXcUmxVwVQlbm6KePIUO
T5KHTAqn01WFJdlmQSSUtlaP9wRJRmtuVr27dNw1FziGO73gGWZR9EbFz98FalPV1dkRUit4B9dm
qKIuy0B372kuczYm3RJ3V7JtgXWTDNSvKyoXDJX/h8E2kwAnJJZr9ReTdtCqHYeZ0T/20dmZ1QPr
bt3yCNh2jkIieyLwCs30E2itdQwISQEguN1UZE8HEUBa8rdvCkR90hpRypaaaHBEagx8+/mg2GXc
USnEvNp91MYeQkONwkSK4mie62wb8X1ISOYOINMl7fCn2tvz0xsP64R0rwvlpBcjA3Bp4q0vvvI1
UpSNCS5PHf0rNnoQ7wkMhikHImnsiP2gWI2EuV5MX0nCMGCFl9XDTUbVpGokJE+LkeLAImqoUJLt
VbHyxp1qeAmGXk6CSHzrNkHX2cdLjBM97DhPg9fcy+mBSX2/szwJhw9yZauNyc9P2XAUH5CvClRi
8mGt76n7FvaxPBD+Y2BG1n+kOdIvcpg38Co5upaqBh+3GE71wAaguXwgjWd8pYNtKrW8sSYMJQJk
E6lTN14siE+m3ZRBYxwukUayWvTFt0obpUqbe5sWb8M2uxsjnGLUw9Vk5Qmxls8t9XrlgJ5n/n28
ywA7d3S8tcwqDcSWfr6YP0tp+7m28Se6aGrsnIUgfknJI0EmrY6hIiFUVc03bP8nTPA+0tH/kT2X
x3jkhipqR+5Uen5tF4S6y7T++wixgBGFMIIy+n0LHluqaGHeh5HJaadU/EXbvCtoxbI2n2s0XuFT
3wXyqK14iXLAi9hMm+VFTURXyx3gDvopmJY4lhFIMDRkwfRgiJ0WvxDNhPH3ZtOL8zOgc7eLgvmy
i4BXwkI7Mvj2VvrcfOiw+8bDQqtCBvgAJm700t+CGgggHuCDuzLCB+FB/6M8ob6BnCDRzBFbMuCt
M1qQlRJ9XOmAth5KljPQuODoQJUGtFpUydMU/jmms8GxLptfaIF2vUF8EAQoKbFojatztkKKo1l7
5Pw+VdrqLaxoa8EHyuCHJGovTXgMoymVLIlFRz01BvS6dL2QQYhy6JJoKnVUH8D9BZ0ZsfHQOjuG
Hc+Fm3pZdR4V9zp/FNA5G4A4VwiN5TGuUkyvYna1LKT+sGmX/aVnl7BYuzzba0NzjgwgkFSmAMT5
oeiGsM8DvRk9qs8kxb5zFsB/MkXl24dRoHD0tlgXrpj3MqfhzVEzrIZACuNdcpBGj1ozMZ7HG7KP
MCnuTx/Jwa2/twD9AyIzVCbaYWbqGhxvDxLYomZ2xf2vc2pOsPXqIIHX6njeKYfz7q7hfzRBUWMd
kfaaW30vH7Z8a8sYwtYP2s3ESrtMf0xQ/dp8nBgDHb32qYCfrWZ9JCiuLmWwmPq0WW+lhEmHW24C
6PyKm/rG7o9fBqpOvz4bHuEf+b56OpJU2dxUxco2WYVIEabslvhFRpupP1mh/rcQIRD7N/xHJDce
WprirnvfNesvxoS4HgRDW2UhV8W00kcBkCU3HbPIPsC7h6wLVHERjnkjMxdHxztIXSBHAoDash94
jmdUklt/DXviZRYCnwF72gzgNJm94inUnTZcMy21fy/2HmA2yWHfBZFhBrIYuKbrN0sCYFgThBgj
jTrLOHYWDV/mSNwJ5qxzWKfup9KPxxll++cJfc4bW6lEyQw2wfRkJUNBZzYp7fWoRjfAjT66c+gl
+n4DiYkKqymO0QfPcACGARz7dG5W5L5uFl529ipN0C+nSkRmNH+/DGv14xC6ouB3L5XEE8SsLxoB
P3dckeOGfmyjsJs8C6YDFGV3al9b20NEU3H3r8s/htEJQqCzrNN5uFzwoKZ34iZE1JgHgBNn48R0
UOOe0tsT+CAg96QjJXNZUCkmJwyj/sWwHu/kieLZKCtem28NrbSCGTp70PJvzO91Klq6BnCj1yid
ArJIPhiw1rjWWd5ipu3fNbbcRHazQj/6/3UlHhnuYtV9ZQag9dhNn/Kqx+IQe2c+JKet/ow7+nRI
pGHuhoYT1ojXKZG138KHO30sN8+ofkuLobCbUh9HbGRMbQtx7cF3lxEGDnmzl9+CsajcJ+Rb8N7/
eTLVgVOb42XG0gproTYjUczjPtyoGdjMCvaOSsufGAguKvNTPhiy+4UYQtVoDBhZeCefQ6mxhLfn
2Ijf4YxNWZ8GyriQV1Dx/ZtX02Zr3N4+hXRZeC7wBsdjr7Anp/F9BM6ulTLp4JfQKP4gRNNdtfFO
VRggQkePQF5NrOYslmDwlRFnLJPPa7N+FSgdPBSbRNfAL93KZert6JivGeXZDZA5wIadRtSVamsb
O2xVqwCWSxsNWvLimW5Imk6M4yUfgsHuZo7S1pqjakCoYwnhskdldfzn1sC+pBLjZuJDGuBYROc/
orQ7flmrOE0VEVkfxwMl5wv9X5mDcWnkh2kWXnlunyK/fUBa0qTUUhgYgbi8fuRApQ3HYnnJPgzF
2mFUEWm4XjDv/DXfgtSsvX/qYeI9GwAxLUYmdPhmAO96MKOoups+0SW+zVtSk63ec4lRjFRxSzhA
AJfL3fqc2G7bbgUC6rML6VffpDbs208mhd0x0O9yFF5eOR1O6NgyhxTsnPRxrbjgoEYGdKGIvp16
hKnXDv2ztACOqZipPsIvgYwowMOVhSrd3O16XovTJB96boylhjsa9Bf9qIflohOIOTFs++FupWIr
DfNfp2Zl9fa9OflZNixoUASgl3oiesbjfY8G8GqwTeowrAoUriyK4Q4QMFNMtNzSyV8tUJqRRX8/
j+U0QhmbAqnhYtGuLpA30iuAQM5mpEtJqg9wLaUr+ctFjbhSRXkaSzycGoy4e9O+XcQ6Jyz3+/qh
tI9HdltEZdPGpR/aPhv44XqBaAmFw0S6wKEHjkft5uxX41jHbMb3gsSOgPYHHzvI95SWHMXk8f0p
/b5LjVujrVbEAtjk6e4ZCWJAxoDxDU8Hm4Wh22yl4lzqdniG+6S9SrQfEDoI2rqhodGvEyt3J0sx
dZFhW2VBvMujCnZKasBDct4cUl+gKBFEC2tCNkaOsLu9YCn4uLLsnIb8nTXPJeFkzPGpm4P5Sc+F
Ax/gB5uXxzJuPfYQwk7uAoiCFydFI4GggnIUvRw3qzpTqLDWEwDcJClE+aWh0JkD3+tfwYjaUOPx
053LtRuGHadlX6ZQGAz1RO/lsPgNj7NRGuMPjCusElKPs6/0P/kfOCfsrt/P1bsNoh63vognvPps
aZWdT4GHspUexm5UAkVw/xJynRdScO9+P+PxVsEjM00boz6nwH/nSXowCJ0BJ1Mv7xIxKk8tvjew
uLxzpedOY2ONYae/T+twWKJW3SSxOHtyEyuzkryed8ExIdzG1tizTpf/fR+5V4WwB8KWXYNUAvXP
0VVwhAXGxcshN5hQjDtG9sF76jRQ5WCanZ1/Vf/H4gacTiw3UTD3wp4S4+oAYWWFBTAd3+2y7MP7
MWq2FWJwAm7U+Edd5vm0OoPdghzjBSQVo7lMu+K6I4JUpa954WhllnzPSn3E/frBwT1Wc1vtB2fT
xODt8cY8XEES3HEj/sI9iy4052JZKL12AWfY6ezHetCU1UbNnoCBSMMHQv/jzexz0xRbITaJ2vrV
ZmwH1iCG44wf4MrNXdStwXBkuJKbgLA1c7oh4rnxchj5b1ZWgYkSE6anCBq5WyfoKvE+E7lm8Waz
od1+yuafEqbf0ZDkFrTQPe0ewfiaCs00BJZCVQqGT0lrK5ZLCKRYiX03IOL4RcH8HRN31NQI06CA
BGphw/2APXtYlBtWVbGsvpM3vnhbw58Qb8Ll77sMdOEabUPTjrXkDOZ5WL4aieiG4gyv2ldyFhng
w49SrixSdnr7bReYLApt6Yq75WbB/iQlBqE5XgAXzyGysX6byD3WzHMXNhSWWZskiMl0ate6p3gU
0lRSGS6YbEFMTWRG8D+M2Dke62nifQuTruazzgTaeXac3GteXzEPcvESnL8lyeOEWIeRZTS6mwKS
CO+EqQqrM8jGeW/TBVLSdsRYp9eBSGnsPTLgwBYxcJ4ujyqi9BPGpb4bPNYzQg+QYUMg3AtbMThf
GnDiEnlWf0CvZ2V9iB9T0P5Ip21UZSq7/VBNsCcURjVrED32ol5ooCddHiUDULnM5biJOPenl9uv
zrucNV2LHYpNddtIbQ6T8LFgKAPOKH+pmthS+yXdKF7yqGICoHoOue/af/J6jbPCAjEd86N0ouPe
t+BZEUXB6p+Ysp6/vunWWYDvF/MC5ewcVhlugO4NoSeeIDKJoyJ6niz2r458y6fp5PXK/zKxNxx7
H+4fVkWkIhgTEZ4A2O9f/B8lG+smN4EKSm+Th+Mmp5HA5PsQJrlwchXr98QCDb+YhT4d25ABMRLg
QJr811AkTwdU5v1S9RzsiHEIsx+aht8+qRozrfT9o2Z/j8Iidz/Vl3migqiMgKCOsClDqUY4nz3M
bMXKGR3nnzsgSgrVnc/19z+ZbNmQSKe6kvvll/6897UgjhvfdZPVcFbSAvnyN6AS8pqAj2eH3auv
cN5xbeh4P5xvD2wmOwLB48iE9odoQ/SwiirSovYkYPloRjgOVv4Cu96CeOquYyZ7avj0Ht6TOY2d
qFq/52s6P1O62Fn61/WkzbKmY31cWd6erVX/wUjq0yyBFkJV0vBHRMKFRKYER22GISe59Dsg8kza
cpacclOgRa8pQT2JnL9Av1/txCL8e/oK+5LKtKnACeMkpLjy6HzDmOjUW52BIGbaC5BfQ5yCX40O
lw6rwiC5Yq5mFh7Wgu9J3SAt4o29MT11f06gbiWqj8RC84sZcqY+dtwUrlt0Sgf9UDEO/lkxjGdR
2x2CNiHhg4t0BlbTf9RKwhCqt82pXutx9tVrvIByy1RJuFkXNvKWcFLibGa4TU6CXyY0EaXkQJnC
gwWrETKmPENWwPeInlPUgKx/ngIpKMVN0TsOSkfOxyH6AACJG7SRg7INjvHSShLGuLIswcKywKbx
FIf0nw3CtHDksh8qeUOkXekPOVHmJHTbplPhAT4Qy7K9WcketHxmIowDoQUNK+xcFGbybiTza0NE
Uvp+iYMEOem8IDOpz3cpM2dfGZgbwkJADQ3ZhqKF3uNWcvzRQS/huKBH5Jr4nRTQ5PNALo7ZyCGl
1NmjdrNxtXMHZdN0bFgQF/aDFppT2T1lSdTSaMRvh8FZK/b0vMw5m8cEyCENR00dcLe92L7dwCx7
6FNaf19ibbZiJmTMKY7TNAUybNWzxEUfWnsvFLRowz2vNn2K3Sqxii5NGJEat9/YD5F8Hlv26b9F
rvjovJXqaBwVmFr4b6Ko76myeDufzKBaUnUh/PGNKG69oQCtvja9qlaSlRokYnnlFMxceBMMatzr
uYXNTh6psZYemR+Kxh5g6bLsEYeoUPSAxplkiWnNhDhknQRbCYO226GvFfvuWZWuOmKeVl3vuCmr
XB6IH3RFGEcf88VBnkko2is9b++RgUhlOKDZtKIBon7L+lXw0BTS2hD+VKvtJ4Abget9D4Zje+UK
OyE+hK5NG145Sd4nKKLzoU9ww8C8jV0faTG1JeSU1wKBWNs1yi+ViZmPqNbzdPOIS/RVlHKOpeVH
Ol5PKAepZBt8mKfAQ5GPpXc2AwBOqhUx11ueSoPaJJ/c4swPyuG8TddIIbO23Whmj9e0nm1Qw6pN
ghKBvrJiMBB7eTHqxtlqYzRn/Wm/cfPw8uR9TYIvvEqcyhbIRMmyZhZchEIVxp80khKhXuyIMQkt
b4LOh6Na8QGMOC5MGmqWD3I5au4JbIMFu8pi8Se+uWJ6Nks1oAQ36be1WMlF9zvntL9gYCaf5M0w
klLEk2DSviSG5aTLkmlpv6Uv+6TcSO9jA3PFuXRvkcLOPeOv0+s5tvm1GQeUKC81w44rIYjiM8q5
vNZQsETZVlAMLIiGvSNO8uvWJmFHO8SXpQXsA4JvB3O5sIThDUz7CAVuDjSu+c2Xwu/jhlCzLsgE
EU3A15zJ75D/wcXnfK8asBJYODmUqxEC5X+vTLU62bEEOft9Hu1R9ZYEKlv+Es1acgVa+OUka2Ue
8ZdmEDxCseEORXFSlWdNrexjY2NEA+9XJyT10QFYxgPxwptRYj0ZZ8lfKAVIMr77I67yOCogwdqt
7CguIf4pN3sotiKiZdOdmH2PnRzEOmBX3B5rDFzskebjJZPrzXBLfiO23P7Lm56fTtPOzJbieLaI
Y6IV4q+JKsAJ/32TE8Jk+TAB6K07x1WQfqb+qYj4Vsd3JvwVB7R0l1fUXtQOjqvOSz/YJKwRsmgs
WZdTofaGyKcERkwEs8CiyABBgVu1zoGLks+AeAsxuX9mDMVDWk4z313yiPISiTQUo6++YYvoz4j8
CxlvnJK9486K8Jm4OJdE2t1N7XgXQvs2qclLB6eJs0AfANLGhdAEzmEjkzYE0LEVqgU93JWdGB1q
f9SrdB3kD/17GbvKbZH4zxTGLDO1+BfOWkeaNhVtPdZIyQIwMEAy0jL0jBKUroWmMXWZ/wIM2sKV
QjNaqdjZg0D68Jt+xzML9g3D4YUajD1SDB4y/oTtWMgoh3m2Qdzg+zNUld+3RGbotPJeLPrq1fCK
SjosOnIFOwxxWG+HE3pRpM4EFeTCR92iuepDP7nc0y+/5ZBxRHrv+zdhfG4/+YexALyVeCV0y73i
DHfxw0GTGGwq9Vo5J09v08qVn88vdTcBMqOfWlS0WpnVdf9BhAYPLFIE06bBt8KUvvscaiPP1B7T
ALZgC5ogdKyUb52/1Oi6gi4h6GsFVh2/h74JBsxKezfCRy9C28ClEABU3caBFmQoJbo1Z4p1a0CN
Cg+9moZ+Etm8CMQw3Fbr/ZvEu7E1GPwU/IiciZhh+c5dO+YhPpingUAVIsLF+l3dsE6izLC9HacB
o+s8dGoyoN6dSNc6yYoPocSp4lJXY0sTXDm/ElK17Mu2OpJv1mIIuJej9uZZJzO3S4/I66zhB+Op
aoSkfCiAfBgqjIDuwO0psqf5tm7zTXpiJYUeyws3gfcjNzqygM1/zG6NzRv7GQ2LcWKJw0j8tqSk
/5lO6lExVNM7dNSgEMp1qN75+m6rB2UnSwGh3B56Zd6qgkBfIzwB5uG3sDfEN5WGJUsG05RLk/yX
dAiEl+0pclwRjFRH2TaSGnod1jLxefcF8Ps4sm20z76g+u/bXObE3vnL4NGIOROnabPAoCkYhaeu
NgSR6r8zBjv6u0+2iO45NBM2t2Y/gEWQwgKSv7nJHjmkqbeDNkus4rMJ9xPCVZ5LIWIFuRNHDLkp
4YtPIR0s5yDN2oj6lAk1lEpQ0hJghdW3snSA0iORT3sdk/cRIjbCrCC2lay8DF+mYGdiJzaB3n2I
0DJLnvAJ9t3vkfvWN/O6v7E3R19nxhYqAKo/loQtzMGGtbFRZLvnvI9R+Dxc0xeQyANmQmHhz3ye
JcC1BIkw+DsvrpxcsjA1iIJMMNlvYBq95S2rE8TKhC1o7QWzKFLeM7/psmV53apCXtdRek1jkbkb
ztIoHowrF+KdDFH5PVAjT6K2BEiZgnvMAayjfYn60ACqN13/VlDBChDoeKtTzCuN5Q/BJ48BoURP
w/q2Y6zeCignwzTc35pzxqM27mu9adhcMyj2zdHBBfxo5jV3r6ZIH5Dyj/86XsY6GwnTaUE6da2j
Aey2bPSYkrSNDClJamhYJuSnXFTLJ5ALa40uEVN1OEf8wMfRYIkXq/HPKG11TC4HC0sH4qQ7fd4s
Uqir2Ll7F8uQAiMwWeMMR/sdWfJR/IyMUMRi219r9dUOMwPqUP2BHnJbE71L/zULkzwLIPJeRLMg
IwF5yU3d4iZgwYAOIwciW97QNr56Z5ZGQaKu4804x9HUrCHh7okNOA8D4l+PomA3M8Lop72Y3sTl
EFA6B3XQ0MAuDqBfh1/dq2L1xxn1b8WHmUoEH0MBT1WrAkhUwqtGnwCovBr1F89DGeewEiFhwj7x
9bSrBkkFtz+YjnDgAvGk9WJppJzvbkqE7emyywtmxV8kKgI2L53RoVzvMc459elnvNUT6LHbHnRP
XYDUOynYoeou11dISKattmVsVIy/hZtxwQTXN9LO+ZlbAYwreO/EtVfQWiXT8ub7F1WPf/pB1yvf
a9g9IxV3ElunbDXraegl15w9kMMrswjj1cisYQQ8llROPf3yOSXLxpCpNtrZ8qojKHgr3prwZtQD
kOtIZ8y9lJsxmCV7jzbcIaGbcf0JhqRZOLYzi4XJQ6cnXcTrMrPPUkqGz79ikjJOIcLDXkRDIwID
ycVrUnp10TuiyiZbZb1bQlrV8rAKKDbuSgZ3+i+Tm9vx19IoJhLZyFDqymwzTuTo1/t36jUwbk/L
I+gU0wl17cY87XlpmCYVj+zJiNwFMO91deYEaXSfg3YapkpL7wJBKHNHgGrGgrq6Fwo+ETGYFICB
rzUvejypLU76KlpKe9qIO70W/HhDJhTHiFpHANlL5Ya3SYMmSIxM19y6AryF/vg6bkVChp3mNVuY
Ll8tRFNB0TiVjDNZLqjwEfEHqRzOum64kvxO2J2Zr3xCjPWZUNChK8dYbhKvgg1yD6ZzY996v0Gf
+O+FVfjMo2pl5GZqXU6kOcDcuxv2MkfStHUjWgYnkrVjJBpqo59T/V10Sr69apJpqeZUt0/x9sjQ
fY32Ly6K0+h8C4ZVbWgM1bgAll6zJEEtI9NonW5IuXQjzBVHdQpwD3ZlCZs8lqZxjXPfnb5uK9x1
872g8052azOQc1NbWrDGWI4fexX3qj/IH9eFuVgx/iBh7FGFd57BwXIN/7y2ezpSJbMkaiXEmgfF
Rwx5eS1RnWhZUCg+qnBoMDS5TWGSv1QFFKYY4i/mIG8y8W7GISmwRDbMVU1900z3F93h2r4OxYVy
GhaOW/UGiCqoFVamP282kfokGjB/+Rw6oPz/I3UMK564GyAMmRlSC3PwdLsyJIkzokLpm1k6el6P
jWf4wRrmB7bcLiDRUGcyb0lV4/hkn5Lx2Ew8dvf3zrFVEBhJHTb0mFZSfCy2J3astaPFjQom0CP9
YMyVLbSmvS0DiHpOgdxFnJBP1rB20U15uiNpj7lSzEmMV/7oTvH12+qkflbqNQe4sJJWEG+cKADm
DL9Jl+8fQWPt+QQ58Q6zdHeNCxEi5157+IW15Za70eATNm9/ooFs4HVL9kFPaOjK//appCVXUyUY
58SkgUopJRN7mDW1pRBqGm/Peom6hyD8ZM+hc0JZLKGCHP09U2tIMQO+gBqsRfojuhHTeAHg6xRR
QheMhm6HUSAQF4DG3ZHjN1i+SZv3tWh0Nyp5DzWD3qIHNshLOPIQSOZ18sGapqlnBE3nufD7He4t
uaw5UHAn06nx+C9IS9foH8LRFS6wvMhvZsk0J//ALzLcCvDFV3sqS19PN9YnXd04bpZ+V6WQgAlg
FY4iM4qE6ktfnLkr2me9KxolMM5u7prEgDgq7tzG5Bc9yfhHP5wzbV1NwtiVLauB1auSqS99evx8
+SfGpWjIVWxiyhuuL7p1DcJ4JX8/R7kJdL8i9RdX5ma3wMQe4AJ06HkwPBEEVN9WSAwMkv3UqBS/
gvOj/1wEVwTdy97GEm3lYsV044z1JNWLK1QbCr2m/CKa9m63RH7KZyPt+dKqSg9RVfXHJ7XQd/CT
OBvqAUNkBS02ssQ/J8UcxpzADQM/1OhuSFnhqUaY+zkB9JjOPy9rd6dYzKA/I11/a5ulnDWwORXq
2ml4zYH7iNlvYi4XTiyzWQgXz7Ip7dw30rg3+GIToMTEHCcggdLRnwiQsOXX45NFyxbctaOo23eu
GynZHq51FGo7ddms2yK7JOUw4V5Eg21xiRcNW2gzqm+xl7Rs252JLyjPzLnZS+UtJEo2Bd3gXVPQ
F5cXUUEJG7DrP/xxvHPrSPWAOvdZrIySDYDM8xEaVbW6wo/eAmIz1san2JcRb0QwHoc+3EtIFEQc
8hqGPBikgFI07Tl59nkFj6Q+BkPmdBfe4LB7AVZ7/Xdcs2RRAn+NFYWAS+huRy9bK7I1GSG1roq1
pn0emfsT4vMGM1Xnfn19JtGQfnlT7xsoIuR7+8LlKFN+BWERoZr/GLns9rzgHD0fGX+vnbeMQQT/
jelKDZVm3IHs1wd/uiFgVEWBRcww1I36pwvzuH2xy2sP6XKevmMnKR+jdFZ73/TgOLMV8Gf9d8OV
rkcOpYj3YSi5D3dUCCgbz3aU/D0EVEm31hgwM9kUYUhk0QU0RXCcami5vIoSglVAgHPmnoMwbZ2b
hvkzLMVd0aRG8TW+ewLxF9khM0sksP7PVNvD0tX9gMj+AKbtP4xr1O+y60yB7qYDq0vlQWxbzbIY
kg3szC8c9iK5F/wOM8ibRLMNFc0agUCyRn0bx6zQpm0K+iHJ96zPV8j3LWFXe5DRAw9kL1AqcbPU
Vua5FVG0hN5tZOFTv2MYbNn/zCElK5TK+S0+D+In47E8k14mkRTeQ/TpUyXyaPCdx5HnpHOi1V6n
zDSSDZabhVjCqlkAbNUi9ObIoi9CdwhZhkGGzZUAcQE8Cfx1n/sIH04Z10VFbOrazwouiexxQu5Z
pLGDhPw0s5A+pNhf+yb5BtrfZ/r+P0upiB5LHD1g0V5BFO3ESm2ehc3D5AafKnAky8z5YkX6nGyU
DCtHZJFUIX5nkdtTyqdfJAZKV4n1RHNimdwco4XQVJ9HqXfmuubpdrUUm+QY/7Z8SCopdXez28LW
f4TjltYMy1n4/g4qt8WFRQvPNH+jmYhqEspHubSdfAm7LPy1+CFfUl+TxUwri9Hx7bi/wOpCZFE1
9olPp2fPlhxEWh/w6Af4Zs/gGjpz8l7EQWKs5Pa2pLwjCsfxA1AtT5kMA0yT7294IBjlXTeS7El3
PEOo0FTAkVKCEh6NI6rSkaPbql9QPTXH3/0mFKW/U6fkLD+BzgVx0sFfKlRjTcFmKIL6vbSszeth
quaT3SSvTi/bqeaT1sisW2FdPkov5EVX8mPvMHrs1PFirL7CyC1XWt8qEZqJtjbc42mBEoN9vLqO
EEgAyOEP4XQ3hR4yvJQlTfmAltq0wGICuVt+5E3d+HF3bgdmUNd1v4p80DVvkWShQvh6VY60tLJx
HrwQ2/BrRxJtpmQPM+DrLDt1c0PMzrL2oktitGoT72psUTNbRKzOcr5uzGgVLAUUH3a1SnFB1FNU
zAqi0pqeUI2GUKZ/h1+do8PQkCtFOoFhLxm4bqyLn94KEG6fEipdVgPvHF7I1BpJ1iA9rvMIsq56
obauFeomW2prsBXsncEA5tSPNfLvYWe34t45h66lpmDw0qrntwujHl3/HwPieHKHr84D30lEk6Tk
aanlYtwXlkAUNfhlWZzBLkHZwyxcD4x8qZHyoEmHjn7jqq3WN3l4pKaV3UCdLmc6j7gYOBRMp49c
q8DpBbkbTGAIWajsvzpSIzQV2+xlotkilZdKILB689n1EXfdjKtTOpYJO1scqAIh+CZe0bOKuPLx
nghZ0MQIXN7Tx8lxMZ7VFpCmqDgfCxT1AqyjW5ZC/d35cA8VesviklPS5zKlORTYwY9JKHMOXflY
xWdK01xlG6yBlmMK1FlRvfZ7RyyzDBra58kNHAtfW3FAuPtNj2T67XZgV18MhVJ4+V7kvqXlO9aB
I470nAc/ER0oI4TvKLuSO4q4qQjcNY3v0Qqyv6rk8HcjowIbf3Ap48rh2yITsPpmrrnTbw/7KfFp
q/wFsK2d9Kh2anLnlMLu3OzJXWd7xl+cCnZEDJsl2XVJIIa9Mm5jVx3q0KHljyZJ3nZOZ1hKYl6V
ElYM1+W12I2OHB29b57VHJqsIeoRNvGNt/dEaRXXnjOEjpWU4q5PRpTusw3558cjcIF0VwySP6t8
EbBObO7EfN0eBsY4cyfMN9SFBGO01aEm50S+Gi0Sl7uTG3UBu3hxCJ18W1qQw8fBRjbSLU5ZgRlI
SFD+vod1EXtH2uSGQUnLT1b/Yq9Ig08IM/kcHYIbZaxLwKsRS+O63KqGdoZZyY08u10AoxOMnTxZ
dmjuLiVdkmyDbjCFH3KvIBAXHQSAu6uzkL9CtkleAdR15cozJSj/Xe4uXL/MWCJe1IKaGbbU/WyO
W+ZAGg8CzXYqvkcyXIMwxSsiBZTzHIU2Ej9OXnFQqe0fJChTLxt65XqNQC1Eup2CUbMqmxJ0QoSo
vCPxQ9Tbyen8GEn0uby+SG7ij1X8zzLq4Qve0zYQXR0x4EVb0EBlMtu0wpiYInEz/iU3wjvspboM
qTgSUtWaElWgRh3rQjE9wSFnlJkj4btPKH5au6+l4kpBZJ4avV4roACOUHegJZtTXuH4ENMq1t2H
XVq8XsvAloczPNgBkbZV0+A//41MY/amrhmpqgVMuJyDJoK4bXcorVNDbXjqBw5JaclH75r4+CnJ
hib7rBljJ8Ju3dMVd2iuA1WgJnvdG5OC3fZBixfIs1sUEH5ZxmEkw4vuu0quuHLzQRPrgnEG5vZw
CKLM2HX5SdfiGmM8T7KXiHePOGr8RpDYccaxZ3/TbiXEIr9tYhM/AoS6ATUlWYuvqYCjbEfBnBVq
HaCaQXK0TEk7y5sri7VU1dwf1XSymCp7/pN4nHgcjRjZNueMuhf4RNeQRZVcIHhPZigja9JEotFZ
oeZA0ty2HbXdcQYB2FAHUh0LFNwR4uor3nHnslMccvne8z9MKOQu75EZUJzgK19pUPSPVbx/6tHJ
56r61zmfH0pAvQaZXw2ELGd0qCVEhuByO8ouyUILJIdAAUsibmewRT/RbJ1XZprkNg4UCNNsyVBw
VNAOXW1pir5RIpbxoMqx4Viyh0nPf2IClbhdrkO/CpZ9gfxUsuJheIgbPm+AgoT7c/vnQAz+Fafk
ZfXFtOhkdo1KhhtG776tB2/sQ+BropV5XJbTCEw1DipHxlLgN75IV7rQn6H3watTu1aECsrN+AaL
9pAvnLLADyiT4TuZHOPZMinO4LOlvYzaOhzBO9ZR7n/nVxvXeAPDnwd/QGLBBlfUPGa0+RV4VjbS
S2N/XjOgz72N7hTcr1K+SAnxbArGzg+R0fFmX8f249LjsR4AWHmQBAqfC7038KFS2wLHOnCX0j7g
Kxpt0lLbqb07f7O5rZPSgfM2PVtK3yP/Ib5uOqtw8ySNIfj/LhzUhBHXetIItlGJPffVwuBdjX/u
TxgxdGMgPtjgFsNaiUJzxqOQNT+Rpv+dMQoUEyAWQwIfkaji2yi6eE5LccI5eyE4nBMNQ3WgDo/O
4W53Mqo6II6rCBmJUvG5d+TB/o82oK6lLrr+guVNDRIpUuZ4SQ1jg7roPUfxrlMOrdHMC1xQ2IbR
zzgwR7jTrKMKGUA20uLcaPcMT2Vqb55YASHmmd6mwPoTJ9gYKCozasLAuLoi5sdt76tZ0cDRkRGH
A2MbIqqW7jaQ2IPvnz8608djepbClEo0B6BUt7Cd2QjX7GON9wN7FnBc7kcCQFLav2a3NN9ciGFj
9+ReZUjYJ4f3s0A+FtjC0R8qWYevuWylWoVb5Bp1AEWuXz/iLj7rqYWLeHfQNzGSMJF/H6CG4/1a
NbCucz2vsn4EqUeY6nQu/KQcONw8BrSr2JwIjb0F3E9HjgfETi+zNKp0S7VxLgvZ1v5c4DWG+3I5
hWF5Z1zV2R9L9xn0vWLOKxJ5C60IcFtZUtPXSWQWBjShFdIYLutlyECcWQ2wdgFVlyxfKP+gO3+y
Sr8NcRxLVV9GICtOBECSVQbunN+1JqcKFTWfyTkjF5yfR/eJgiESdLnjYtfMnSrjEGqYN1Wvw3/2
fTbrp+GQ8v+5EbH7YF/23pIcKp31eK3qeDAVg+Pxwxy/BESAbrG/FB86PrU2X+CfXrsOTv+Omlnj
DsNvnc049ImaGXNh93is/gcUIG1sDe7mS8XRVdEKg79mr+F3oA3uOVbWWi/fqmR4uAzqzqhlGkB9
NAi+NPcL8bhEhowuayBHQYhb7A0cS+YMxFbHyqtp4F5Cjl0a/0tJOGi0INPz44gHkO2n7OZNE4I6
c3KV3AKTB2jN7SFD2kAdd3BMIQCQh4x2sUj0eS+BZAj+mCyi7efZnn/FQFH7Uv8H7Br5qOk6WuuB
o4IsIxeXV6Nrcm+HJ36580eKw3/frg2LvaTYCB51+mq6CuUaQ+/jnW2IZeBVjTRTXxZhisu/oIFK
IalBPYOGv8SVAH904k46NneDbVObQ0SGcadOLi6qOHC9yBySK+wdBL/6+bNduuJPXNShHAHJPxCA
mDonLmopncbc9qaj33n36SVw6VfrAlbatialCpMmXG9HDZURGeQn6KC3tEhWR9kF19bxe3rjzMae
qmXLK7HgBgtB6T1G/KmHfsNQAKN61mLoJL90pIHsf4REi2+cGb++HvolpDEmAuyiRnoS58Vy+rj5
XIQ4ZRIVkUbQG46UBVtsccriP7Ku3azGjEEKVUcCIRaMFaJAQSJ0+nmlADEEhmPtmWnBzu2ykA7A
OLp0IhKOtwh5P0oMywFkGZdqwxCvcPrMQxtRS+T+gXszf3wfql/Rr5JgfEWTqjFVr/vHTSeVbspL
DpkfNaRRWy6lWQJZt44aBt9jNzZBI7J3QHHMvfLe4qnrnLoEZGlhhzd68xA61yNXJhwil9lRT+uZ
EG7cTygtzuUax9rw30Vy8ONuEBjaP+oGBlk32BnyNtdXypOt/5J3XPD5ADJXtaNojmGqKG+2qLJj
XscuA+3EQxlN5w5d0W8HMKHfAxnfqKVdst9onAiDl2is1Ivk/6NCq6yMoSPLw1Sc4BJjI+ELz9Dt
IEnlr0yKperro3ePTPFiVH6YdCpp/0sxwwwMFz0Pv6GZpNfnVy9bS7OQX8GPTub4Tqu56bTqNG6j
VtUO+e7lbMT0OVoyKAc/TYcLyDSZv61MWkwXWuHO9InAKRdnfSGHZ/vFkE/fmR/HBLdOKuxM2cdX
xWqfoBWu9mD4MJsNO2NKcWSlepMJcxnUOhZ+6k4XWCBlW8TvqdZDq8Dh8F9YAFL74Zm6E+rF53B/
XCPSPf7iGveiMUad6dY6JqF5GJH6Y0fUz+AaUWdxdzz5sWsSJu5AKW47BE+4yl9LfDGvx151wBe8
KMNvYxeOsajB+IzhLpsj8jowfqcz4L+Z3yF5qbhCNXoH1lB3xVroITcWM/M3YH0/ZbH/OQa264l9
ZSg96q+JJYGAJwyMfytLBv2B83nNMsZz/6luzeHQEmVmjiNNGd9k207xz3uVJZ2Q5pzQOoLrOHp6
w0gcy8M9/WN16K4isOu2J2eOvr17bxbi4jWxyKbOK8D/RWlcPDjpcJBF/0B6MoPchjJ08HZqzKoj
nSDaLLIhCDSyARBnsuP6i7BjMXXP9lyb5oXR4DW1WCJHKpZeU2NlJDFD9EANukVdB4Vo4fYc+Cr2
EioRCVS6i7jPh6247e7hf4eoAUJp6IV8IkCKIPdqFD5//vprDUDNqADtLidj4c2evWyWt3OP8CoM
2UzvVFu/31+DGfaV0O/UAreoeG4qw9+47bwsxPnY69/Bk7WlU4HnAQdv/0n5f5i2g5K4k73SDZVO
/ZSkDI6v5+rkZF+SX5tStnN7T4sodOo7ylmqOu3yLqsv16jBmqFt2mppVbp64CY3lceeWcjlHjW0
GEi4tV8bKsvvXXMWIGVY1g1Kr0ABj6x0MIqxGIZ/GiO+te1ZLRvd47q871XkF4qe4B2vbZ/GTs9B
ttRqV1drI6j3PXXVTDJvMot2lg/7GqpVDs975CIvyZaEMFEl7WHV5eihoTM/DS7TLO5l13weVH6m
MWq/hIFLbeKKr/epR6YPGJjeAwmKlu86tNGJKXZaO9ZRbYBvbuyN24GV6yeQaSopWqUtevTLqRJL
jzOyBuzJ1kVATT0LS4MHwlDOszMYCN66EK2KtQedxO+eYQiYJX4auNVXp9uUc3KsdQEmXw5wuVgT
hMifpj1dNmxCVrvEfq2X72QcBTE3GKs+ZhJ50i2bgcWL2M4wf3WiH/NWFVVw6Byljr8rVBg5//eo
sPZwPVPhWHv3mglO4f5diJag6U9JzCrQ4GWE1KhbYW4weVeCngIrhH3eX6lD8gy6toR9/oMNUuAT
TJmudP5WoVs+hl0YFlbJpADT7FcQtUKmI4Jh6PnJJnQpqhsSaemq7AKp5shdVTOvKgzfcvwnZg7i
twwmsdwCnm/z4Gn7GfdXniL2FbvQ052X/18AWbPzAcc9RwiYuxLtRIled57Rr0XRsg5XPB77/hXs
4RyLoNTxF7ozM5QxIHsDsw3/8jdWcMm/O/BlZcOrBka2BD7Q46ZomdGHAftuNjh0THX1PaGhkTrT
z3/w0csMn21tQ9cwtLYkfKjm8jGQXxq6H775YTrGWp51aYJSkGDpwc1V6hmrI9/sgF5Q2aBSeQbx
b7aVI672cRIe+o17zi4GrzM2zSOfl9aS7eqONL/Q5/STWGeiHmtGGs4ZvJ5WF9uNe43Lwv6pHSji
TYwWWtc3iH0dhakv6eL8jwHMAieEqanx5Ewd5O9+wGMDl3ybRO1nfgeQ1uCQqZessiLtNH01LqpF
yRXI3C01NAPdLsOORXI8BXGroiGDjIE5n4FjtIyLQxqTuPvrsdUmI8UzjWSm6ex9PiEd+AD26m2x
llvSnyJFmsdoRXvDyH75fr9dL2QW0AC32Q3guG+HzS0FPiwAwSU5ryT8dwWxiYJFCuHiBVGMQx1J
5BmqxHhqUTKG5GU0hMW085fLD2pPkSxsZXUNIbp8wrIHwYeB+tNR9ILDAvvMcn4pPWYZ3rOAJXLB
wj9BgxYmXvxfAyuacdL1jHb4nrDmU/a+WlhyHUSSbnbSCTXUzKYVsA3Zf9WGhcOSHWSgtzR3nMdl
rU1zSJypfdruTwkzWLkfuNAlfQY4K/OEVFfPddC4LJ6ZNmqRc59DS1yOHufLb5t1iipAxDFOHoh9
VHXjmZ6lA3blW/y3iAQVADl1j26KFUJRliITpaOvGYmziZFaL0rwib+ybLihD0MkQl7lxf3Rjfvx
CQ8ybxDOARsoelLSSoh1q1y3V9xw3Rx5CBcxN0yPOZdShRjDvQFNzDFElkA3unVivDgmz3PneDMz
tsyg9jAe74y2tNKxunkMI/bIg+6sAJ/Oc2f0TH47wN82EBomR1qhNmOpGi4Ss6u2QrbVeAlVEE6n
iIvClND00fo2WkWv3obxOmb1PTcxXlwBBUxfSVzy4xl/C8uyWMz3NdLQ0BzS0kta6uOj+IYG9LQ3
WGHeupiNnlH6Q1aJd1vojBY9h4W3rVjAA2VJZpvPstOLDbjqFWcgAyOKb5ft+MSNtNzTAAFkz2aC
/44EkOCsN+JGxJEIIGYjSFzel4lFFNnOB/tyHgbcZ257ce5hhIiB39J4eelxXPYmJZH4hiRcF7mo
gCwzF0PEyNtfdLMLJ9IFkNAdSVO/Dba5NEQSNE52D4Q0J0AasKpu46ErKjzp1vuuRk1jfOsLi+BR
Ng7FcQagAXiDoWaWm4b8Iqo/jdOCdk7YLxnoM2hArLEVGvy6hPaq0829aoEYnzltsG6mPccHep1X
L9CiFfyvsW+yvIr/BmdYdQkjQLOGhrFTmcVCmX0EVQ5qFi7DwfNrv2nSroakMaRUvfwZbyTKJ/ec
ZoYCwroTFz12ZUeIx8VX2BrVSGtDl0mI+HxzgRXjlb8ToHP1O1K+rmSQwkIdcWJs4OZhAa232T2Y
qFVP+OgquXQLMbbI0i+wr+xzEFy9OeK1Mrr19cuYCZTohSPlDgfHCoWr3Thlm8GwCX/vXcXc9Bn2
q8i8JcIcs2KrYAwPbBSp/XZstGaAsPkMbIZX0jLaJjwdGDdtMzOiUY+SlSieSI58f0bMVvNhkqyH
v0sZaed3AxPX8LFQBdTyTFdXKOu4VP836dj2/Av96uW6elGyren2NozY4pBBu2tNHk4zVyhV4tWU
qGOE63OsMZ1FZ7e7B4G36a8cvyEDPkyf+N/lGadmJzUkax4hrKprhHwiEK4yPBXubPtcvnneZypQ
4oAFJGNLRbgbRvdM+ENiDkhnannm9WVwu3fDfyEl+LXXSlYhHDcZYSUtaOZsWugJdSMxqaEIE7EW
uE3TrqR4+ce+LoYY7SmF4/IkcI3VMVu7UFOEZcqAXRrYLXkxPFTqiMtnd0vCVE7OM7fFILOnz3t6
4HRqkON+msfteNTP719T5B1ZPE6zZnQ2GVJFiIDsP8WztCmdK4BiYkDVgoDx8SlxFSEzo0L20O1b
qQupC+5RCKKAVOzfkHibSr3+sH0/GrNYD25dq9JNutUPgcPRLCCJY9DONz9OorgA3GMpu4FVK0Lc
4x3o7jRaHANLAE7Xv9YnBBsaSashbfk09mQ/y+4e4CApg93uBK8bYSOrMK43WEHqG9erExMFBonz
0pI5DbcqWlIhBrzs7WHE7BUk7gyj/Cy2rCecP5BVHkEIBO7vDkbUIfixCxdlAWshOJI6bE1R34sP
9cm1bTMgPw8FKvdsSvk8snYUeWGF3O1pyZnBORJ/zE2hTWqnTxdH4sAEoM06gCRFmNpTUgwq2ero
F+vr0s3MowhvLXSnBun40CaFVidWpJXp9kEQPiKFWhCeBmf5MnvqYBexvaJUwgmGZUdW9g3ZqxKV
oHBJiRA2ojO0STbgNx0p+XdW/HEme47ioX2lgHysvuH1ZsJUSywIoWl+qtiRRWpV4C/kiNoqLG/F
kewIjZ9VHV2EWl+dLwpZ7Zz0c/8tfsADZ+w36oVpODBWzho0e4sYicUeM1rpFiPvsY/KxTvfaFRV
i5o4YgVq2Vnc2qFMyCU/Tko97o0FKQf8ULyNNwsNQdkzVygPQ3NNKCfdLgFeL5zwR8uKRzZDOtz7
b5kvBC81Lj64WCZ/WPoeMQt7fsjV4b9zYRBIMHEoWSdtlx74HUXCIX8SBIJR0ACBUa/0dFJpeQlM
XVPzlIoYZuO2mxA10UXve0gc4lxUpB7lXcRZaIK4MBQJ7vGVEhsMkBb1+w97PQlxJhVg/e6B29T0
XQZawa1UdPUaU3LIYI7lQ/jLLo0CbVtTR0GV6YSS+FiEjBx9qu9xzEnG7JTuG+ZEg8hVJSYbskJD
aCKSQZ5SM68OCH0qVDjStlvDomsgCVpbeLcAnye+c9Xv0XBm3KUDYcP3N5Qc/Jq7tSv0SYaSEtrP
WB3EPFAAxtJcX0FihMTzmcUZSN48VhD93h1kUicXtK9omI6qgR+ymkJobVZrjjTDhBfuvU8Q2G71
ToascpVU9p4Qh2ztqddk+xF5g+1UJRKxwi0NOXYH+6lrq8XLjRK4gdvq8bA1eXqPtcdTQjw92Ib6
PKKloCmXw0pvZVPMsOcWd/jLxfCsMSI5M8oHS6euUZwYfsbMqYLxVvtQUvDdkuwlmDDki0ukgb3L
v7dAXOKyVykphP+/nZGXiZwto8Cb72piKsBjEoHcpuXcqQ5NWG290jVqE/j6NOUh3fxVtq4Dok2n
WQnzJhqQXOTSGriLufJBHTnvbA0uRsN5bTEIhHuO5Pk2lb2UxCRoYJmThCne7VsLs+/0hBizeNLw
Fv04Uy8NNeM/DkOwWXxR2GvOEOTclTyqkXnmN/KORVrtuElqFAYtQZEwXE9gRCr+dgZQhKqjk02o
Hh6ugpTI7DKGhMISGSrxC1eNLKBoAFCMdCR2EL5QBElM9zg7yBSaIYpUFHHv/JsRgkaqSFlAl3m2
t5OXqHz2fA5I7i3rOO/OK2t+Y4VSeupIAXTH9cFcH5SJDE1Ay+5dmQp3cVEtCgcf441NfEdsGv5t
HDFWwD8dZBAqS0ESPL4TgWnlq9w/S7OM1ZKR9m28Kq2zBfQiFclSvlcY6yoaOM1RuA3HNHI21vqN
fDLgiQ0xeucjc3wSp1dLqDXQKwj+mRq/9nQqtg5bHk32BWz7mk4NRZksnQ5fZ5TQDwDqWB7Z3Rr0
dhPsvcMMrwc2aHzr8KfWlEGBjOO3N3t+sgs0BXkIKL+oRaGw5A3jLJEGsQo1KHvl6Ch+eFSCMnai
8eezAnRSK3nlUi8PloLKHNe/gzG+zAL8WKs9AlhUWtfqh+dOhnrDbT5B5qBNNTy0q+SPLsX98HY6
4UCuH1sEh35kdSLotizOyjV0fnyImD6NuT4aydQhsZHJHFqWNeVXvSdJwC+cco9ALvyS5Pm4AVfE
b/BsD3W/udQgaByuy8Btr6n4k3c3YxlJ77LZ04GXfGb+kJMd4OFQMGqjnVdHfGfiro7hwYhFLi1z
BgvUQrFBlma0q6By77TIIwR7acv9qPw1ekybsFCVJXhc82eyUHUHfv3cG6n8TvrIzjYy2rYissza
N8tPTnSTSuuVtzvYsLwfIkPNIlKUgKNNPEJNJn56v4Py8v0QGzhilrXhvk3n78dH6zZSL1sowxAk
8MtbRYHTJgajxTxwwOfJ4CtLnoojhYQK5iYMVdqIy1EjC4988hqaLLSSJ8fprvmXOv5Zbu3cMyRe
SS3MXOmc80ssgffW9yyyoOQxvetIbG/5HzWyv9hUOnUStoQGdOYgESK6A3VXj6ZfnfeMCIvfpQoW
wNdxIgZUIxxhqwfXA628IB4g1NedJ5PyFTgbhuV4Md5V1O9F/0+DZKiq/XkyFXp2B2P6DOtQV5Te
/SJQBDQyN2c2EXKMmOsW2NTohdnGz1rNqgI44jJPRvixgPJySQhapOcbZ+Q3eOb8i2mLqLk6uNP2
vSvqMcdyLj9gkwp1RRMwLBynVksUbRHclsSb93n1wZnil4llqFRSLxGg2/wO564cKpSrgnWdIc8i
cX6D+vztCNaGHdw1Tsio5v3IfxjWDFCNP6QaxipxmEas6ZjTaqJK1kn08+RaXJt/bBLnWMUK+bGe
nb9H+2FfGPMQbMYAGnm1waDAsvglED/xVfeDQX1E5rdQaVkilG3Efj1b7avft3eCiI9Ov0BaWC4P
Qjfb5Q+9lshpy5GaiyIh8+ZyNMqZgYBq69RAK9qpedR/qHMrzRWicZp+IqDbCzwnHAwNsrwPmHvs
YLgaWyDna1icZTEwzIa16/yg1FUgOknjX8k+fUq0O0kfDcXYXQQrCdISYvW6X7gvPNmoGgcj1Qjr
k3ct7JFWSKCpCSI3wZl3OGMMnUl9D9tD0gjbBwsC1xzZ9cR3CrgssvF86nG9GbsQwZmcIQyFwjdS
CYn8ekFw82MycuJH/mVJHgtVCBbcpwDjveF9jJ9nGZVT9Oj9FshjHzWiO31bLJxV7RnC4tGP+mQU
wWO/biFBGNqPE0/Xo7bjfgmLmt7woWOBjkhn4xqRDNqiX0jvwwIL0UA6bSnpr4grLy8YbH+5r4rI
qlVCO4ZjAGhEYXpHnP4TpYpymNR2/njPuMHCuo5pGQ+3fsKEe0O1GcCPnYRX6acAJ8oT5jUewj36
U70LGbluCifrZ4Z0IQXn47z49ZNzmp9Uta3i2nKjb2qA/zfd7RZL+X8I7VmzTCR9e9rnAZ6i4iic
89BZvvpHgvWQPRbsJiU+VrQEzzbFtrehFApown9Y69ERbpx5ase8YaiStIAr4t7bwSrCxJPUSK4F
fUfRcmPee54PAQFh6/umhYOkROpwgHMinble8iQR2npGJVIGvtMsdi5mLENeUWgcLcCS7r/H23lG
oBqlzD4cWUD6wQPfPh5sT94YKRSUvUp3J0gHtZSBEyNzb7wE4aZv4yIZZ5uzcqSlzrzyXIlWzotr
kTAUaPV1fgKZEzWzwjTQXSUqAqIrvFMQ5jcSgRi/8ulvvrQg9gkGnKFHP/g5Ww8lG7Kq+mACKyyP
/qAViE3WCYj1aD8lqnSCPoKKLfiJ6Q3XwJkBfcIaPpe9oCJJbX1pF+aZ7tLHl3vV6Pm5U7+SV+o/
r8XQGLuxDggaKAWUHJ9O+t0rGPXGczDZHoLbV6JtFQkRcIu5ctzAlTXDsuaPkeuHQeuNJQe1uWn6
6TEe6NTjJS4qv3OsdW0SL0phE3CYGrW8ptzlIh4etURhC5JChQoNOXgofG9gfwWab37jrFkSh2uW
Kv829BwtzhpnA6wQxbAuHgz89GRTqh/fFvGXRJgo066m4jD86SbRijFtZFdujVqbdmk10XDTL45i
gL+MC3h1SVBbjO9nbyt47vU6yf/NvjmllncxUKrTkT+1nU+09DBL/S98WddZ+mu7Q7gI0tBQaGiE
gtfZ8qj2e7q5LY6TrHFBwIdknDpU19NjkEqdMQowJ6DWYJf4t8LZgFJts7oYOO+cpVjklZIA7m6e
SASMFhmPnS/b9yikyaNxObyvaGhavScqXC1A2mYArmGc3PQeUwvLlz14ZZ6d+cHu7RdQDCsdlH6G
5Bm2hc5So6rEAd8/oLuWhfoRp0c+p2Y/yZtZDKk9msg8mMy3VkWn7JTIL3/J/6yEB6DuFSblhdhU
b2llAqrCk0fRRsqOCVOasJw1xo4mXWXa4yjIpU6AvS2IMuIBOGNZWBgdjCQZEd9UDUWAT5mqXLqV
5yLHqEwSFeUYmC32SbJS9r7GsaifnBZi+qV6aHcqScURRays7yt9zL/rIGAi/nJAUJTvpaa3kwPS
CarI2adKQJefWkeyLlT7sMFTGlgrVp07AGDg/Tn8HCFc62JPpdbdj+PH3FnltNgv8ol9QjmOMBA1
3GsVl0yy39yoLR/TsLSll3giTjoAKfQrLaQj963hTUN9xDZIcPeH1beuwdSHFx089luCsT5gc/s0
qXN0GLdFBOgXnITL1X3ODJGYbDzXjJpdBb7pPPeNc+F5QqhwI41F2e9mL2DuElRhc6XZ1TkiV16y
5rmRP/cy+IoUdKFK7HuLxYg6Tz8vc4Gz/xKYOmVHQLOy6myvhslkTme0EwAZ/SuX4tcqOFjybkiB
JESvFZxdnmUeMBptKiFpptBmTHKBHY8KinrRHhvaZx5l+Xo+XOZ7agU7gATVYI2aPP0ZLLTy/DpN
ebXgZrnYB/Bydhd6nOXpLxr3QOLbI5T78kEqHOqimukdJsQ0Vs2ggbHNmctqBUCuHw9jlATaULJX
k07g2tndV+rdhaQicTc+VU+V7fR7l+XJWXkSMFK/sWvQfOHCR9CdMn9L3rBKaSPVSbYo+EkyAiIl
vr7iF6ntXeJ5ONlHmOLwwmB0tB+nMhlWZMoAeTuv9ow6evjsxcA3Tg7ZxssPtjs4VNbRCVeO8xLW
rNT/qk7CVp8foURBbchWpuITgkUG7SXhjc5I2ZeoBtwh+5lrpdljgC2d+FHOL1PHsnD3yEoZpWW7
tNC5d7WBo9jUOUGOGVrCwojiFVzTt1S+M1XQ0Kg8CTbHcPkjgHDuqGX5vBo5j+4e8L+TCMGt8h6U
dxUyekGI5jAFWRujJiHzgdDbKfCUnSCauNVTzNFKqpP5Q09pfwy0uyTHovDcf6SJZaLgNmxU3rlV
woWiP98g5iYy32n7MFo1LIpcyr7q4XcJ0ehsN0cwoILkNeoe1QB7WX65NHbcOxeSACDaw03zBHaM
tQsvasGDC2xRxWgZHoMm2JZmFrv3+fZhN3uA4Bui4IeuthEBMUg97boojjpcee0IcGPCn6LsQ2Nr
sFL2Ik0xQrpELk4Mv6IwKxDDNTLa3tIenVPZAr4Sn4yOW1Pw6xc4HbGcHeVuOCc8KU/4AHX9EKZt
khjmOwfEneQwprhU+Sn2xtWKxpiUsKEQvA4Wct8HtUup/rvYmT6CcKQ5nqKE/LihTRBfZPge1CBJ
9dcA91FQdXHMHHbRmqObs0pGtdZLDknK9rcfwwtDaRhXWEGG4LQ+PBTL1/2QKC9xg7d32lZ6pMuT
9EtWUS0Dw+MSUSEbl3+9/K7kJJaAgUUMMxpMP07yXxy62LWKgvH9S+dS9eQTOFYSIVkePBAxqPNA
DYW7S2g6LjhQDMql031TCA7DQoV1aX6JwBG4bdPT66yavXimnTzigs4siH2nku05wJ6toZYFKnYM
4GnjzTu+e4jLQNWUkD82+t+uYfY+d64nvysG5NPMuya4eLs7hFbhcartC1PHYDZ+Gc90WDM/JQKt
YKOySIIvoO/JqsbHzsGGq+Z7col51aGyoDIl+lakaa/kjmet/8lFqRD25Bp2yUnqT2FKP5G9SU5p
5VP0MLjwXzHzZiqNik7AGz2kZDXOTfcWi08GNcHiNZsag30iLvqJn8C5a1e9s/9CR+BFzfLgh51Y
C4O4OEaerigHrmReFVTaxl4ao7FfZ9gJ4eoQdavd0e99q/DaImilikpN+yht5VRWhxEH/eN6eFux
GcR9eT3PxxVXc1iU7419b6nZZRUnkzDQi/nIivksdEaU1A1E5JML2RmkEGzXpoUCSLL0p6DbPfch
Mp8bxLcAV4/7sgQXSxwNaovoQ/DfvOVe/RDfPSLz+GZvhKeRmEfwU74WuGDI0ACscpUZBbBxQHJi
a+SKhDqyLslm0jtt1JlORWHhAmZ2DuV5nBDJQ7qgEHx6Xo9EPcM8D3KVHOkHU98Dgg2Hpej2ZP/K
WiCcUFrOrpCyMhUYgADWIwAP/LokcFFUT4/LTE3wHDd7MNs57P6ErAS/JDdKLYIxspiwJV5oFXS7
Yhj7A++4MJpMDQjcgjfotJhvwSmWO3KGB3hIyAN4u2lqS7n1p3LCYF4CU3gnAmN15a/VCJEUT46d
Pw4kIGz5Jieq9BbiuHhSaqnQK5WLI/5hoURBxgVIGJhVxyYWQZ5oxEc+oVH/VQhjMqA9guYtEGCl
B8t7tJOuFJ/bIQlXAOVqrqWJ97rNyoyFaOEhZv+YysF9w30tDHvOjZsAzmECDKz9eiR5HStmGxCH
952TPgnylq/ZRFP+kfqjtfrBlnYJVgY03h/wjzg/gCrL+9EyQQtmOfbce7Q0gm5XxlJ/hXj4EtV0
JlMGl7grfv9cFtMWM7SWrEcIz63vQmTVFoKW6mSlpXXDI2bUQX6r5kiBA7tSiORjlIbVWLOz83gn
sujAply2hgHntF/t2Gi1UggTGke1Cr/8JYGxe5SLpTj6LrVa6vCQn/IA5Lfw+q4dUqF+kdp6KUwN
aZ2oxq/tgMO82x/JiKQkE9IBk+UEIoqehOWLbbN8bkvMIWk66t7sZAy8edGZZH7gaW6QMySrvu95
dkqUfkWxblWWKioqGI5mkwKQUZFLGYpEcYtrl8UG+ebkO3VtWN/e//0vl6HDLqDkd0gDJC9kziaX
HtGtQvFYejaTYeQUKRNPO6PE/2g04aHDCRHMLnrMyRmlil8u8BHxy1WW26b8eFabBw7Ky01UZkJt
9GAl0Mw7tWMAdtstQVUQlnnovlB6qGukXwOYBEyF52B2rkNmVX2+fuJnLNOc5vQ0X9moUVQBHZ8D
MVcAsk3jclTOQRvK3dgnHBtjM2BDmXVOe+Z2+Sp+8ZMVGqUXAErC4up+S3k+9kYpMLMWUfG4RYza
wtR7dazYTeOtSd/cCguc0ovGc9dRYVGWDYbGPy1ta0MLElj7LBI1xpBQYYz2YXQK35jfFBMvRHb/
AkEBF/kubqw4WHgdNX0xa041UjmDocgzzcGsjQq+MaD0CbruHd1tdHGit6WwQ2A71WFKiIqtyIba
nLtGFZDwGvkdYoliNQaxcRE5Js9BkOm5b7Y8KLNzZ1LxpWpCL2cvTnfo0lg6+UaA8anKb1L4i016
PjBhYZ38SZg999/MBARacD98hMZlFzyAIzU5f5fRAZXdQs8+FNlje44NIzZM56Q7fERyIzdKXQqy
hnenNOGijUCteUDdd3ZD2pC47TU4FJNC8mSXwDhljX9KVuiX32BeLvQpVE0AhGeyuqLtzc+z1OU8
oMvRRR+nK64rSki95/j6OSSFHLDO/PCjqvv6n2xcaQ7W4GoeaPHQNz4xcuzyxPtC/GQmM98Wb8Nk
qL4MMH3NQKKGm1OQLXaVq6dniaTk2W9jX4G2RWwj/SocRC+ZB+6kCq23t3kN8k8n6+xRhDBZB3yT
qanHr31PbZuLhz7pIfUK6Xb3Pf++LOtZtLVVtxyNiiwqMuYmKh7cr0/8NIZV4QvN55b9WlAozaBx
EFp/Bo3nLiYnnWhydly/o/JX3X0cZf28m2kXJzAmqtZWx597VvqqnCOYmS+xzQDZ1S8K5ZkKEgb+
XSpWnCEGOD27VgmAfP+BddKXUKWf+G1FYXBs5XXuSgEMgigElw5WaLLn+76Fa9HVuLxyf/55jhwM
ZeX5MxShLRyKP+JdE4hXM9dId3HMyEIFXQH8cN1vsRCCx22lEfFrb1dGUiAkHYWto0BRAEqAr2P1
PzeuCJJJhDcQRYO1p3W8bbaSUlX01DUsWVfMHSrJai94CMQW6vRz/RodAcXwddy7HQlYJ9qWJnS2
Rpk8VGsn/zqyupozCujEV/VJ9w/cjDDJpuL7ixVsdKOr+HU6xzFtSv5xNKO0nAjamJ3QD8kiJqkB
sbj/nP9rxNIHTxnAPhyFhf7voU/DOECrQxdpWjSvAx+QQoH8/J7GUiChtfLb99aCZ+5Mto068MnC
Ygm+shYiZ3UwOhX8VuEDtX9KoWV9L+Yz0DISxi3PPom6AejYSQLI6NxEsL71FTKzNnHg7wLnn3in
DuPuO7EF8s+1/cpxil+tIodSkB+4DVk8jiPqyUVfEf6jUmRVEzCWG6Dw+d23lamM6Igu7LQC22NL
IdGe3cfgjFkvhpAXaNhEfRlpauEHse2sqj8ASjy65PD4lbTNT5W9LZXcWCyA7njZLleJ1Eqyo8rA
Ltxd2UdGv3e9KqC1oKjjHBI2UpUtRunPwgWW0bSwbFDIJ6EmE1Uq5t3l3jIBrFhfzZe3Q0h+VxoQ
gCyiVNOJ510bb0uZe3Z4f9vhP24941aipxCycsaWG5NKqyB3bhpMqXgeLdPkn5r8Z3zdh1zwFi7s
2dQNcjW/mWOP+NnM/BBmwIE4Xr48Gbg1iv+NtUfZigAilUGLrGdjYDXV+fwCdXt0OzJVHmBOstm9
e96Bgf+bAD8VAh0n2WW+EhuCHidNwMrtFabHt4T/EroObxMOtT+n9JvzwZpyuYKI8F1KzYx5CYmc
g6A+HIUCtN5FQJbAplNqWn/YbeuOmqq7AgyO4TfycnnLApGpDW4rDz6vX6gzgzbPTQuUR/mTgE9y
IVXiq8uYwueNnotWlbLSC4/hFQb7jathhgYoebktD3NVbZ74dgAh+4zh39E9p8lfCnH2bOsRWWxi
KyYnMyCmdXkInM8jPN6BMSQqrqXXYyvYeCzy7Npv99jjhCXRAJWLT7IBi9zS2XkFSHf/LYGoSSqM
FqBpUaF3umunlH6wckzq4Y6Oe8UL2vFdR8jXBFbR1ZSm9M90eWnUY641n/SUypf8pKRky/yMTFOw
HuJNpib4ixCic6ySXhUw4OMnTqmrcRaGOfgFT06eiCIu/tbZ0/D08fYxoErKnIpZwjTzVJAy+yoZ
8BCPS1ZZGtMWxMJ3QH5ambj53YgGrXkunqkFe1/ykGvT2eTJLBENKPVmvcE9CnPmDUiV6OWgScTE
oh7ZrqDqlqshQGAXZ0SQhI30LJLhVVM/WwK3gTP8VHyCxlnplIRqf4QibZPbzyYmVjfKgAqd507t
+j2Km57CsVG88YBfI05Q5eRAr/QYhbqIHSi1LxIrIgnvhEWTsNKXjoCU5B7WjtC6QYLuoLylAzLe
gLXbcGISEb6emHCaRDkWmoC6o1jCpxX10d51ky85PrWm/EFs/D4dH1lScKX+x+XTfHM8Xp76QxzI
vAeMdHipiAStv/bIeyk32uUmsqaqK/240pMoZSmpvStsaoih9fvWpVeJ81vCTSVg/l6QqJOQSi4j
exx3oeHQjItPVRjpqGjZ40/wN6y8bCNZJozl/gH9JGEanbGdo27ZGIdQ2Anzo2IVP9CBEi+owiHZ
RZ+T6lR3BnKxp62a/qmi6W2L8LXMIISVBxNo81LpQUiy8t82jOYBrXDZLVHUO79vrQyIOOqUrTjm
e6tZ/7vBeEAzdH4SxzZzpVc1IMP+RmGW18nKZOW9pQO6T8krgqw8KwLnw6RkcPXb8GJF4j56Z+ci
8RUWwE9/mjYkhIyn7sHDY0zvkre05o4xXc+zW7VJhn4wqbe2hqvUSoG/Nd8Tudtx2eCENi/XvuEA
K6PaE74t6UKft3xs7HMv81aAsxwB6awLLLG/+4vrM19LjyM6DSEQ8vtPrBHYBXSyySWArJJ8HPsp
F2opTH5pKnZZBISLUH+QU1/z7Eb9BCjQ4WGdtk7c7xU8yV2vVfU2omgr5899jC2N41+3459owKPd
y9TsDFakFIARYija1qIvW9T+olY08wod5RKzNuSwri4QffFIj9xS3zm2qKSzEGhcjPBCzF5JJcZm
7fcYAreDPPGGtOMtI3X7pXK51uLj/5pC4Awqg3ABunZV6ygPO8yihPDpoIOP3rzV/UXItr0ox/3t
t5sQY3KqI7YxTqNu14BtvCJNxfqJV/g9sGnIUQBswLzpxkLnby7dWAtpkJyTzAUIzU6NtSFi0Zvr
P2UC/I+ACNlWt7ZtVNwlzEaxOjorfn3iRVHp86+1eczwL5a/XOgIELAwE+95Cas6gJ8JzimHRAj1
B8ooURkniWnm/Efw7HYfapyG0Wgk9027Z/W+ST+UZtfXFhcih6QbKv9UbJgDSpy9QJr+XvZaG+tJ
x5ll8Gl8nnzTjt713smcxQ6XXyTKkPdl62IOZurWvbhR3ILt8Gs0VoiSxXZwNRcghiYYsCMUMzid
5x4bPn6EfO+ZTOjC7x2UzgUFUNElvv8h9uQ28V5GE5yzQJl90TGQlHVUAgrrVr/dfOoH/BUNiipP
s0eUjOzUcaVuNKtkkyvIRo3Om9hDsBCTugbhqjy8KGkeivjnEN86Ouxd8lPUJrLCvHfHede8N2Hw
niF4gYBTlKEOdRP4x84TUhsPuMkXK/D0lFWRHG5d8bkzrzryytq5+a2CulZJwd4XIEJ9PvQNQaXw
dAkcBW7dCg5JdXuj8sCAbwbxq0vmvvcPUg7nrm2EXpzVSxgijHpNjUry9+oXuAO6boiY9/TOX6ic
P5Gp4NQXxqy41tgr1A83A3SF/kPlBiyeWDQZsv0UY2x/mUJSeYJGo6cKuIKbpX8YhKXDxPar9WDL
pQ5c3NtP5hvALztb4eWm2rlOjTri3AHhSOsnYpz6Dyavq3+ehS/WIhYJvWOoXhWBFVxKjb6R6CqP
nK+mV/2f23kOTN1dfuDAwiDS28gxYJoUMEcVxk+Fk1bg96Zq6Y3K9jPWQ6x9sOCbUAfS11WJlbn1
q4L8DtSCJEzFzSjoNgzTCGcmTKZRnPUqIwPdCVdRmOQbs9lUjxFIY0m2cC7l4GLTRsiKbsliO5Kn
jnq2r2P2mJuXhdsb9VyJPgAAlOOr4kmXEX0xPW6rbq2TjrXsbreZV9v0f4VhDa2exYu2pKy7KghP
cvbRWO4IRqclpIBDIsUnWTOh6p+L2HQhgXvsALYwnsVD2Lzve2GT/77M5YpICr3eqKX52SXpVKIE
gQiTpwtmwrdVh1Axk84GBb51eOR8VKbnXYzxtrCtojn+K9x5FPJc+FumaSQ0p1BdF0Xw09/q5sLm
CeX/8zUCRD/1hKDchaVV0OE1p0W6KoAe
`protect end_protected

