

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YdpNuWNv5ANxG6sesr+pii9y21Kx+NVDp0WoJ8gKKxKHNSppxy07GkwBsVP2aDgHIw9l2ULLZTNZ
WthaAb5amQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kEIsWLqGmgOl8w9T2kPb2uPP5XenCQ9kpxljFoCEGisg/vUEuVE5EQlDS3+mxviS53p6zH5m8hA5
bszDfKwHD76EbEoDDpJWL09MvEqH4hbAV7G0A9Qe7ZciYDi8os/DYZvhR8zjbLils1MINgQgL32T
+DXtGPXNuzJTAMDKzws=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NxGGOrhc83L0V7+Qmwb6+Gi21+qsbQ+hA/5/9jysqY4QYAqiXfCrWB3N0NrVsGWuuTvZXoFNcxot
Izvlkgh5KOucyz0ezFvnhsYziU+FkvqQYf1g82Syrsz8zvyVWXqii6aXcF/WSMwXtiDjm4MiGpFm
yTcu8CcJgBMXYGVZx6nj+IgO08YgHCC4sfTqmgIgkxkmBrOsiH76g2hPxvXPgVWaBlJF0bS/hLIS
Glmsy0cU+pqQlcfbTEV79W+sXQ5Q3KPQFXj7AhMrHHD9esRm2Isg/tuzcRVk1cq3LsMUN//vGrfM
OKoYOozZxl1/IflxrtIzbjclaBUaFr5bvZYMTQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dIJ+Oh/ID0KokdCrmxnp1QfFJ5QZBtIG4FQx5Pan4DTwhUxDWY/BQobSBBDXzWh1TT07UPg0V7Ui
zobKMfHgBNkMD8/PoD0AIDWLDLeXLvIJje8mGtE07uncec5mJ2eGa/WSy5sFj4M/Vdtk7C/Ab9LC
9qAaWZZ72ZUoEHuysZg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VglxNkzPd+guDL8DGRWVtgWGTdJbzbKKn0hBXJRIK4IuLrtOeezNwjLTIb0FIMSJGqYYwUrPN3z3
TVnjDJDaG+HA47egpMvivRkbnfO2/EAJtU7n0hK18OztWFzW+yXOUsOuQnFS20EGjEAN6HCMCAXS
ralqFAJsvMtY2y3dJNuE6ytT3WYkXmZUpTrJPPJOu2l9mCOnHkBU0dRG7RNYXf1tEMPaZrHSYyvp
XKWW5CTowIM6jJQxDVSVfwprGmWFUVJFtAmp+65D3ADXiHMcwre5cI/ty7nYS3euq41mrkrZyEF4
iH4/gU0xN9mM3aF9hBPzu3xQrdML35ONnUZTzw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13184)
`protect data_block
UAMcGBO7IaQ4xOzxyTEFaWL69LD8gTmFzA+b3J7nh/A+sNy0HiISTgQgzl6D9IO4e7NKNzt1dHw4
CA8F8ykI02nERVUlyLoQZed27KZVH1eGq8H79xOaGvxIV+xrrd8y6PEfWmdnNg3iXR7NV8edY/Yj
VGd3s5IZY1p6WZp2+eLllXZZ5Elvm/aIDVd6BpsKCvcqUaQ4QBnXIj1vLg+Yn8O+xxZJEvQUnxR5
7Enn/ZyNkb7r1gJigy/oNo9vnb75RSLe4eqBZd4Eoy59uKABWRAXByFYdA/7Br8DpTN8msjhJVz9
Jbh0sLdWwjkYYtbB4AFXvMFXvUtR0NTew0QgqCrlRCCPDwJHbD5nh/tF2BDkabQQ6yic/eDug3zl
krnWh2Wp8ZyImt8/pDGI0WUiubjWMPXiIxV+yHoIryTlX8PiPb7Yer4Yuy8IR/P+2IYY681e2eR7
CQisZPcs6YC9P4Lf9HwJhlyHgysA9oMJqvyEfi0GrVAYof4alF76CAOIDXzph2UI+CkIVW9uGP+c
zZVlw+M602y4UhOFbxo5gE6e+cAvH6iCxGnDfukcY/6BJ4sC5XSyzmLe3dbNs7S3HCbensKvAtUB
/5+OBQF71rjgR7oaOY5fqaoarf2CFaLNLKsafJMXhW6MoEBcXpvixqvC5hJWnSR2KrD5OqHaQ3LC
cTkLODKL0nSklH443kVyRiM+wIAI9TEs2J3KVLJMjuHFBc7/M9zsOrswZVF+0gWj3mPCqB9cbw5Q
WT36eZFW8WacxjxomBieDmGLlDywUo1RkdGffkpFu449L+JhAJiw5S+iSWIoGPIMjx/5Av+X6Z7R
9YkEWzjMWf1iLDMZa4eXQCdEHA82s54toHfolt8RTmvy67fLTQbbZUtcvA9XcAHijvy99YxZfVp2
d5/9EdEpaLO/ioRuaL89y9M45qmCRsdR8jPKOuMZE38FBKYMytk74aH7I1GHBh21acWiQxwauDVV
MQ9XKvslU3pgO7BbbFH3thFBV+EIIOpttTQXA9U3xnfBI2udKpeDcHkdFXEiYqFFw8OwqzjLZIgS
xvZ6o9ImE4YU3yDnsVC+TH1ufEbTXyDiav5Ay3u5JV/tWKa/PXGrAoJKuPaqMhfG7Nuj266QkKxG
9fHUkTMSvFuzbBY14tqfetMmXdiD+iH18OZk9qf7gjrB//6gYPmOOjH5/Nt7Gs5BBo4ata0FziKp
D4BpmRZawGpM4Yrgtmo4VHI7KY0vcU9lobK3oMI012rkLKahEi3T5dOACH3hoYYcbftMj0v9blq2
O8YpvD4VHEMxTI7BtzdrVWzL8HO5DulhS0fML6A0hCZjvt41e6blKeJW5wX6zofv7ZAQ9i1Hrbdi
HqIQGFr/kTbVie6fvOQcBM/tzxt+C7YNZh1Bu70gENyJ3H+ntD0AGsiVelDnh4IObRvm1NKGQ029
6fSuRcxUYcPjiO1dl9gJOrApmv7okpZ74kbqo0wEbpuIqMHsT6ojWszn2ui7goRFP0Viwtxi5Y1/
dE3X46XsDw88psIFn3FPbccrEtwUuCtqlCzLjIty3ZcRlCXRLxN4tZAMMalJw3tMy8w5g0reIpAB
RdChJnu3cUsOZdJCKzWJj+8R7+utbK5RE9C4kUxm8MBmZ34RZxNNrTCpvLdg/vyBjMSe20fj0c3+
KT4ddcnnPMhaE+0R+KmSnAhWU5gyu+2mFKXk3d/9z/CxoCyTSB+E8ik/Lb78+Ls5iIbiTXyIz2KY
cJSsynrNcm2jEGVTkPqERtKmCadlcJ/XuZSzHPWQYk8Zg/E6VMXYz6erGSjLgIhApx2p4/eYu0cz
vILJwJyK6JmO15NfsI6KhfDk8Idij+QYDaN1+BF1jcnpLDdAiox1LluriLWqDnIQUCRnG8yC3TEY
4rFzrNMZOZY9mi8FS1xTVx2aRUdXJsX/geFcIx+Mo0pKKxYbBPNcrhhF1HxBYRePYbTnwvrMBl2l
yX4Q7dRJV3NpwZ9OeALOYO7nGXZhiqc9gGWdtrh4kVvooc4j1OAzzyU0wgmv9f6Yi8YOyO6nsq0g
iit6isYJVHMNjyItqmI4I2OU04Rb0bTgqndijIaDd4dCIpYzrr09H7/MPFQ6xu0iOhrsfpe9z2x6
v1A/lfZBupwVLjlfr0yPAAUTUS4hRbqLsAlTzPuo2tqhLSAZUQ3NvJCChp03BLy/e6rwrU+ip5tt
cojBFg+7Hdzvaps+YnwZtUUtQ2HrRoafHXo4FsMwppmxuMfTxVEHMlqLOwHSRq2Yz6zLhHw0OlYm
TBgBZ8vm/JecSCJ1EsmkIAxf/nnZaSUup8ZGj1p4PQjCREwznVnJwqoy66pk35hpvYbjnC/LqFZr
B0fVJXd78V66+yzzctBFDYt7XyKCUYYL1fKoXbxQldNFdDYbuBfdCV4CdJtsd8h3PW4dpOu1ngJJ
38TwGaECn7qAYo32amp/tOuakVi7dZ8cjWJGoxwSsanKe21ff2R2dcmwOR+MpmV5t+/kaiSVSfOY
2gZ57ApbKyuU04t04f28m7nCBITEMMfLJWgkAxXI/+bUGTmVo64b+/iOuTXnOKjMFKbCyYdaUqg/
RtUj/IhGeGlyMkI/e1Px405GRblgqWhpZIYjbv1TlzmTvwrOAR2q1GBZEPdNgFhznSVnxZRm77Ce
LUg+fbk4Tx6RvW3I8drB6yIRubjwDay8ak9rBH/GuDnqUT+I9CFvVsXpN495LbpAvz0YIFLjBF5r
d7ZXxQRZczjHpNoFyaEkY8tnI2mLs6P6Nqeqxw4lrSqFrETQJXuszMHugg7MolRtssn18Lg1LL+Z
F1rnQfmkT51KD56d+5WvsD6CVM1L8zlg6rBCA5PKHnB8omCKHlcjGh6YHEFnc8tMppo5rd8Yo68l
Ml5d/19i/d6OL184c5GNd0YxwoLDgBb/X527l+sGVFo6hNzACNWnNUnHUXoeKBcP6tnRwxpD0bfC
mw5oIEhheZmu8E0o9PPrt05J04nffYJyvzqmmLl/ZshHQav1G0Glb+1PVqS65zJStJKMF/i5Vmw3
ezGWNsvaS383sHDPaiuEtL0J6YNjvHWg0ubGpyAcLinD0xwALK246HLhR6ZwKoQ309YzeM8BDkQV
n6aAz3M94CFR/AIXzLfOCHWMRxGkSOr5ZptXtByK5lwnfl2fWMfjbRc7HlapsT/YkZEahVMoB0IN
/5/jBeAFeDKTFJax0bbuQxjwfVDx4mJ741o9Cg1arPJE0Wb4dwn9tqcKBeoLK6CTKxhoBUJSzp6f
uF5DwGa7DhaCXfdsyi1xWh4yU/xr/Tc4DgwpWHNz/MKNZT+tbWfFXgBNHj9EASpPZaGuRCVpGf45
J0TWL6AIlafMZeDTuaD2XkjJ4hZacg/2lZJCbpzzirXcX6UGXh5gQhDhyfPi3WeK26zKhwg0QfZ/
BEk+OQTx2eSjZI/LU+BZkI7cMbFqVsW1IjYY+9vSQlLKTS73mo0uTGOJYO++TDOaaoh5auhV+mHG
ZFS3UQHq4odvQtxPzbu12wVwZCUDSgF70io+eAticbPfBu+32rn8+JfndOVk+bsLeqLbJ2PncUhc
wdRjRrEXxsMf0ydIx5k+IyHbK6oOOXoht2zaG4c0Gn4adNgD/iW/J+kP97HIJblses3UUTaleN+z
KRv1PNuhjdxAl4C0iM9q1ceVnhoifDtwwiVp5qx4xQ5Mn/rmbj8TWn49wGYXhxZEjq2wMLP3zJvS
v1DRUPw+o1gTrlcxNjNGfF6JQN+MbkGN4ZkYDeZKAAcZfLWfUZHR2QQKo20UgVR/sXEymgJ1eSsf
Bl3jOycmcpiRVYVYy82ZjOy0c7AZ19BYOSyL/weNobQ7TmjglbljVDPQmtAZyBTr/5f6Dc+MXzsE
fhwTE/i8YKJLUN8Us3CT6kvyMDACo4s7ZZVh5K8b0bvdeo2buTWarqOl4mRt6CgJSjfHfe/MVS5Q
1ngnugNHl7Zi9z2wIFk9RamIGFuKKJdFeclpg7/QvajTK2D8K53mREKDyN30pKHsQ7tKbTI5X+bl
ZwcJdfbgTHW2nOlQx1RA/fJNWABER7kX+JaycASHETQkCZIwpWWBt3OMN4CyYpY9V558NCFot/pH
zX8suBgAGj/bAOOa5K2zcKXu0Fklpa7Fck93YnrWzsMdr9WutW+4S9H2uIleKUB4gcA8EAip++tr
YgPNrEJbyNhgQsxR1hLtDEOUSodIUHYFLWSWH2lA2kZsC7y+TUPNEImREhuT2BIY995Uo1bpfRnB
LWbtL2eDOXXlDpzePGzrodyDDTWcbCO2dFq5mdqf9NplLm4Nm4dq9vq+hDhA9lmWAT6PPDfX6WfP
srlJ0T+8/dDj3pcZ4NAUhtAjRPsAwD1nFjIvrO5/WB6IKGw6W9ikby1jRleq1lfKoh4F/BWAqF6X
8wANLBPbP0GakSQCwHgaTO4rmgWxFPIBXmNgp4t3rL4rAExvqiUvSwlzBPoGsMqYmare/lSvF9fN
GdcLUamF/nZHUSH/AeNjJfTuz/bGx0gBHbGyhFfWXydlAwcfoumz7im6BPEAER7nlHXauJTBYwNm
uKNyaeyM1/yf1zgnxQjGsCCvrYMCCbWp0KxfMX+suaWEYLes5uzsMxRPaGNBeqNIJxfBHMpkgovM
IRGIcc4zdxuGK2OWgKlg7Fii1mMO7u5hzL6GGaBpBWWDvXe85Tb0mdTBWaCQZLjBv2+5gxHuw+lU
0MG16IEz40dp5NSi+83iqfrPRmRi1I+ROEIaA7Rzg/KntxLiSpnfRUvXgWHj95xc7rkSF064464p
gDcPvp4hEq5ugyHVpGRvfDlCjwFnmmVQz0tOzopslT83iG0Tl9i5pVyapUNsemB+414b+OLZ1iGP
MZ8F2e+R5jWYea2YMjOwbSmSsW2r03KrmVAaQGSYnEWrry0Z9xaaM1to1F6iLDv/x6d8bxJkmyll
/LCX+dMkHyfz9qa/H8WEesmx+mkTQmAVsE0vvSLYfn3oAXVCqTANSTKchKbz4zl3QIM9fjuCGExS
dRKkCZ0mn66RtsbrfoevGmLlTXVy5Pbmq2QhTOo3+7SMDAX78SlmvkOowQIyN3MczjpC4XpK7HzI
2bI5SSF/I6luUsmKdfzlOKyTlLPCovAPhmMPy8EEF9H5H0tqTpBPHRG8urjD+RRnMab0eap4dj/i
p3OAipfrYoFIX2bQc/t+EiyeczqqIxv4M1u28qtZ74PaAQgxWbrrxf5rMWJjDjVi2G4VOqxMb00J
fFzbc4IOFYTkL8QUruHfvVpCQWyhLF7NxeAap38345W1X63iCNpz1IFDcTlcwok7l82PepIdyPay
sZVBfY6weNdyawaMmuLfqeAktdFOlIASO2DBG1iwYNb2yRX8YEC0PTHPrhzAqgdUjrLotsAmrGsN
9IWCe5KHKlJAXCVvX64YPuIdNZeRB4JEQCbcMpX8MmkTX/PfrUqQ4dD45ECOxHYa+E1MvgMBcbDy
x5CeLAzNXuE93k0UP2jsKN7pJubS6k+Acv4uzsHDnS80Edq+tcla8OjmYAvcKwvOJLZaVsmaOEpM
w+y4jEfluKg99Jq1yjZ3kZ5YKb5wG3G7CrVy8psaRByyQ8YspnsHT6NYDxbeRxgaX+KvTaDHcxcT
QM/pj4lUu86haj1waj9TtpfRlwm/S2ULdp3/kQQc5KxCegACx5P2KF/pyuZejfyEGNC/0y3V15xl
8QIEIH5d8eLZc0vW0sAvwwY4/VUVLsjphTnS82mMh+AD3+8InnM206aIfLqm03XTlU8Ts6YrFblN
Wjy80H2pAkyXEZr3Fk4lf0aXAUmq1EcICheAh20pwOk6Vl+PkM4nPcbPYq7EaMANgK8UmK9AWTSa
UQxKJRvHqgk+ZFmFTUqW7tKIedink6u7bNvjyASUWGaXgM9S+s7kPsVo/0rMWyRKdNb/ZhO56uFT
zT/clrTPxEpUflIfdR1kerntU90ujdon6D1hb9fDIpsptrzREpnRNMd6hK8/bo0ET+MPdWIiVGnF
N5b9cWSE7Uh0uwEelNIxN1EP4M5gqSbIgnfN9JBACJytVTpTujATC6UIwhkk+uLrDPAN0LSZcbSw
0oAkjN3YY804hr7JvyXX/dA+ax3OyMWrDUru0Cs3/8TGPLlmvEhwT/lB0n/S8pgB6uytlbCbGDzt
8KMb7quE7rpGBKkima1nRrK46UJXcVRERu9/QprVrIVknibwWGgh1kJPXpY7J+VRrBLN7miom3fW
Lhj5qD/G0QyzlEUnfCUZ0HxU3zYVPlXaz91Vd6/IszlO5lbPfKKiCn+jHcytDwXN+IVd3AMM8ONA
bciYCJegZVuCHY86C2BbzkNC26UG6Wy0ynqov6Jqk6x4oQuQy0iW/Na1sSm43uwFBbXHv+06oU9T
oI76lKkqT631oKawbe4L9X5aZ/XCcYqfYl4Z56mYK86uYsPCsJGnmkh+2A1IpPZnRqCeq3YfZ4oK
ZQGtqh3Dwo9Y4Qjud9YiE/q1E87t3EwOZDuNEuc9VHVZNqmEDPKLKOqw+zOq/9cmjvdw21XSyJRg
+r7x9853cLURlK2i5k7mFtFWUBUj1hdqopFrmOG1f34geRH2cGDSqnFmyWSHaBL4UemCyGhZHOLf
zh0RQioIXfC2DKjSaUBVKfPWf1b8Ye3aEFViv2fQhYYYjBYwIEDU8oi187DuimbDsl5PN9geYK4e
gXscZLkyOyHdGw21v81u9TvvvIUHJeTpUCJ7NTZlomLROUK37wLujkP/ZwtAf6kKW4CW5FpJyFvL
8X8kj7srOlTZm+TgP9LvbXjRnhnGtz6UOdI4g5kDmdriiuzubtjjsGOWxRALLyFu5yNBlFdXbGuh
idZVToTqP0TzhJxFrxR9lZ5kidTZxJko/wybW2J/+SHT8R25lf9xu0MtYlJRG5ggSkhVtB9DE5cN
wWcVUBzeUIMByQQVwWyOuibQOXEl89QYu3h75Uzn4G8mKeD0yyGDWdTr4LRW7mKUs4OzXnqKi4L5
dCeF4yblSSHulrVtQwskEFbNecyIQTm6Cn1T3gNyIBZfgzVYeevPYrEq5pBuznLmuL4AhF6yqf7D
13km0u2G+0irgtY7xu1/FykP8z4j1Iu7aRm/sIxk5vvhi82FqYyoOG9rrPCehkxbV43FCw5g/m+M
ooCQC4sqzSZX1RNBnybZROWDoozK09ppoOhkQfro0keLgkmA7Z1MTO9SF3QQ5oAGUtHi0z3FkLko
Z2udl3mFYnRPuYUKCgvVpvq8XlpQ/JJEJFMdju2lx/XDeeUf12H3ArR3EJEYONI+iaiP3JXUhClo
VARuKPphKU9UqBvgOPi7O5I03HPjt9zglwhuW81ZntM2XpqJ6aOFS19cD19qzHjZReBh+ZvfPHc4
ihHNgnCWmb+Y0dSPnwx0u+5ldaEMhoXHjFhIR8ANolnNVtysvnv8J65yLXQPJ9dbkqkTUkeOWhuo
ywYVm9yhVk48sg4IIRvidBBLzJLWOzFn7ZX+tGd5P/+nSzN2aIK3OW3lnnf8xQEuzLXf7mwLWSRY
GS69rcfXWlkJ2cHneZgTiLVibnorwknBTMPjNZdwAQOqplov2zO41Uw7zC51s3I4XuJI1fEqB4gA
ByyMbeOLm5JI+HQKMfFIP4lloHahz9xKtlsSPkhtA1z/xUqvQGBsiwTthoGZHl0uQA/ZSfFfN0QZ
dqxsvzcfAgubR5pM3wQLjW4HfotrMxH5DrX0GPyU4BIRrsWSntKxkz6AqoN0eFCTOKYEg7Oirx1G
GdoxK4S+tR3k00kKrYMrpwoNrxSmx0pttReBk9e1/keG+G1IXZmFWwqKPNKSJ8ICIKwpIhbcC1hD
8mx8ZEl4QIW5LGkNkEeIsY1qzPOreyfjJ6ce/89HSWRbVAnXT0kbwz+fvb8AIfvvtMCY3MPlkT5X
dJqK3Vd8L932Za7G2s0eEjGaK71iWT1pTfOIN7WPP+S7z731xZ/V6oNv2CA75gXzsTfyti4Nm9AQ
Gv16NkZQaO2wsd5/0K7auQcucUAcCQd8KyMsoZtX0CTFNEnZDyHWanQSMgLOUOtqc7AY4+xEah3B
qu8xFaaTacE8+P+SP4C55tJ15nKVCSF4w11FWqDIr67WCzOy3b76kMPs8guzwWXMcKV1jZfqMjSh
jIXOVn0Iehqw90X45Yv7a/hXavcCZ+efOj0eyD2sqbN+zExFbLIpR1+29iz++sEgMsH42GN3YBbI
v6Hdkyr4I+AuNXq0VXX82v/J2uf/8lVboQhx37+ZWN2WyZSiXoi0vGlNcKPyD5O7udAQnf+RQbV2
RzGgKDwU9ZZzxLthtGL12QmbTOCc0ndNZ+0wdpNXE32QLE8mDhxMeAa2VT5TWLm/uogU5+zEva60
rS8VekXjBMmw0QxEz39MYU08uSykESzN1VnkWkpTc3Wxs6NslFL7SqmirSArOTQYJGrMdJ1IxIK+
g5D0b1DXfYvP5N5fu+DM53Kx7Ot6ye3M1rrPTpjaD4HGppa0jLzA931pceUh2baSqoSEqRjScp5U
Jsvhj12CHJUSLq+5TDAKGjvab7wPdEKUsXc1MXHgYqtPSB7YfqjVZiPa4qUc01m/c1UtxE67m9Ah
b5JYp3Zuz3CSGNkhm8DNFy+Y0wWZolI3dSDW0p15Gm/FzcFLufjXeFV2SGnp1qrJi+qOodIfUQp4
1D7/wp3HnqdHHtUG2yqhCugt/VQSQnG0Mrx8f9c/nNfI4qEe9YZOK13ibHC4n5OwVZ5XEpd5US9l
1UxJDwGuY5ph25kr9plXkXt/96+gm1TIiUqvgNBNHNzp+bXlgUgVFP2U4Gt9yZbc7J5eoE3SeTeN
ZPxINztJct41sEI1TbK24r+za61BM6XOYAs/vSYTuCok8Jwwp1j7Gstyw1g7GWJKMypi1RhCsGH9
AFsuQ+UKaEdDzi05bKTs0ixtM2t1BnNbYmfmPWIk5hhdkwUdYnhpw+DveSx5rVg4w8Zau2qXDSO0
lQ4HWjfn/FENscXi4gCq80UQMukyQrmZjwDHoDim3TH08O8S1IwVXG67J0tqECextbA6ueMGIxLh
//O5c8HSEQWrPMMLfSP03FYXxGKJQJ8hjX18cwegAEUxvp+s/a4lJaprZi2gMwAHvfX5Y/TNG9yl
mWmq/v18U3ZaMObjOoYfgormzISoeXV5/sZG+PfOGfyOLXwky+n7DVQ1kgnSOEIJN9Pj7Nm8wgBp
nT6XgxgGksLdvjVvE21mDSobo3fzoEAm7tmVWq8AUo7mgfbxj1rrfSk2ctjLsRbwIFKPGx9Zs1Ua
kaf8Ozf29jQbQNNVE8mIXqxMqYFnGkz9TPn8NVwD86hfqIvonXFsbxwJX9ax+WPcJvYh6SMYof3e
aGslrahwEc4doZ2VtdW0pzaxh/Q5F2Qvh7AN6l0zSU5jnd+YrxpNOxSM8hvviFVDrZhS8GB2HSoR
dWrDvp0pyQwObOYeQ2rl8/QPL2PfA9AxtjfqrShy81CK3hpDkAK2ncMvd9OoCZpYT4cPO2N3xDro
5qHj/AO8PN4mBlJxH9A/L3hOIT0sK9MzSbeBkwDhiz7rda9eZV8BQmBQuO5uAOuKQnic8C2UjNUC
CsKbVb945WoIJ0L10COy9pLXRSTPPo1JDZvj55K1TqXSpp4fSCNI05JuHeQ/54+Og8tJ4/1jzxjO
YPtHIhx++uwULvIFXIItLbHIGtc5/wDfLogveMMoK5e2xPtmyFVqo286QdKaci/xOGguXxFme/Op
jO3jdKKPLxtJpY2ZCSYxlqDJu1DhikGqtRzxfu7dmOYV7LEF7R7OIPbYgSrKGKRWgWoQgulAU9v/
YITC9fQZF/Vqgs76PWK1GPyIwpGDugoDA27gbDxKH3Zvs+9quzg52FSXqaygO1hlKcteTp70duBR
cXQqLaahpYyAzsKlfq/54r0+7hWZRsfo11nPxw6+Ka+1nYilPIb1CpwBiUY5awxH1bvxz2P4UZqq
h+NLVTKM0jwkxV+iHhVOdR3QzhuI/0Vh7/79y1h3P88iPgEGZY8haMC9hV1nA+/++MaNwEcC3aqC
8L3BdlJJkKMGeJJKpb++4CdpLUy9fOwRMrDW5s4ZUcp9nsR7WtrdGzEBE0WyEmLH8XLlS570vFO8
UoMBsfMX+H7mSf/XzbvBmLxLAEnh3OHR/wiySeZsmL7+/wLXCTPwiMxuFg+ZZq7XLZ3mZzuGMEoM
nw3AUdm+pcUAZeoGKEagiORo/HBn2NUfBmz09B0q1ehhLQp0AO8VzgiJXSQtRPYfPpAeT1Kuz7Bs
u5SmQrK5p2j5NF9VSlp+6/7PGXVzoJKKFMlaiuIiAfwNMhGiRxoez4FQXMaeamz12OSFYXzCvnqs
1ME//Vp9W3OzAN5A7hBlxF8KigN+0t2N8KEC1AKiLQnjJsHVl2Gg76xpFHP1OGQM1uCp3VUpr7ew
mY1uZmSb4PkqspduLmKQP1l23ZS26gBsLnhUQoNRC1h67a1UEKrd80hecLhAwnUTzxtWn5cyoRxj
QzIuVYyA1tHtNYITnxmBBR+mLdGvQStQhNY2DXoSMZdqlWwcQnoMx2VTF9/wONj2kdjy3upGMSpJ
LPtE8eHbOx0Lc2m5MrA4UEssDr+kCZyMzjVVRGM8zEzJZDSiFfW04cCnWpp7z24qOi17w0FAxTjJ
A23PgdFuPLfd1E6GvEh6Xfspl4uZVbWOnvwXQx6Or02YHvqNzjP6ELgjhjhxRE3ioBlABQ7hxJJa
KZxGEuwOlUUaplAtBwuncrVRBv/0eDR5PobCTCMj1plxRE2zjIKqCH9pZfVEqFX7aCzq7Rq5ZJSn
AN8gLodPCu1LwbyGmqcNcPir7401RpmDs16cjAvQNgff0/G4Vok93PNq8gm4YVm6TbB04OWbEN2b
gk1vG/GDQxShVGIWqTMWp4KLj5K7V18Jg4PxlrqO0nEX6HtffMi0pEhjNfrTaAZfqcY5SWzPnyLF
7YSktJ2oaZzDWzzLKITsbtSbfOSjlh5xYFtbUhMoULkmIS+RvybilE2kGIfzQIgd6oiM4qNmBzGg
4rcYBYqQMYt5gGY47+KpPBQiIOh6u5ppNqE2M2dyhXBXerp5ZiOXCWzaXt3QoaL5ED22z7dKVy5m
R7fAEKiRJthcHZk55EeL1dIFEX91J9MRmLpdS0//hK+2ZB5RWEaQ5YbJ9x30x4TPP8Wisjdu7tB2
NwP9XKAwhuroZoybLD7lhUV3fK0yAJ5+qZBN2ol7/1Qh8m5jm2WUiUw+/pjewJWTuvYsg3eq4Af1
hK6ppzwynAuuk175Vf48FGuWyWIzeVXEv7kIqKPhbG4iC27GwFbQvYqMLjQiLwKp3tRKuphS+p6N
MHHU7A/x/119FntJUSjJb/bX4fH1jdtB5w4qQ6M4Jx7f5IyZ0HI62GLZn5i8mLmEr8hVqgggS+8X
m+WQCphArkoCXjiE/uenBkVnnWI4NQlHVRSGMpl4RuPsEzTMNxFgb2g8MW31yEB9o9czozFjyzJT
2mDGY2l5DP93UGhytf+K9jLYiHJtEh1E/EPwzlR8uQeojSsWSlk+OuejZWmMhLWY6b5GjhUdmofg
JWHOGALH4iDrz0pIFzf9NspNX4G2nTo73CzhtzCgbQQr48ZHk1xVNkBx3PB7AQocy2mEQIVfiBjj
VaX9OjRUGGWVIAxMpx2Mx31vmiTIane/bm3PMh2jLqJOQuOaHzl0jIuBduFGs6Yx+xd6kiRCzMIY
y9YEX9+nm40I8+qBGoNOJR+Z4QTdoYQBeOFIZkI/5ans76jt2BYkEQzuusKpgc5pGSM3LKIQrC82
2q6s4B0T0qpQ0A4YL6R7QTet0Omo/DLiZSR3+urLZ0RG4/g9MSWQEkUOeCULZyAU9ykw5GlleV5Q
h+Q+zuMqKgFbdjqykRxJoWIdHCSQKEp/6Kdz88s8jAS4/Zik50kboHQ5+N8nuNL4YfxZnjah8blv
u9Aut8QGr7LasdPUyyUIyGMVRL7Z/JOFxJ8piv/Ht+vtlhg/5yHHRRzYIjSRdCML20wXgcw1NM2p
LvVhyb7ZXptZbo7b+JD9wWldMG4hUQ3nluKcZJAvADK5XQ6bbMomXJtdN/hYOS9lg5SeQeeWRnrq
DLTgQkk6kQmL6HA9FSjYxd8fYrT6lJmDTkchRrGn/jf1jMASr9z/x4bX2zeWPua2iwLfTJUhxFdE
2xAzrRVcSEYjbNjEMfBca78Vn4F490VLhJQlAfpbssaKO4kc3Gfq7NUIAMmM+sKdrjB6CGErRamc
zFKgt+dbOENTISpYlgpPNzqD5lwVvfGvbTYZCwVxGwriTD2GdCGpkQ0zi/jY89xQYQFo7ujdz0J5
P7IEEvfOpn+h6AY8zMT5DxpJrZmXlvLHZduYf21WUX4iWu3vdV+Z0i0K3ls1/jVJwb20X0iftPmd
gyjINTUq/IScWkL/IxqtwX6tQsXx5QpoIk0vnHHMdGSqLMYNU2YTkRsap1Z4jgU4KY9m+3okYRBB
6uvlfElmkwzg2Rk8Y5VgrGxCbxioQU+0gIMaWC7fyI7JXo323tePal1iykWJ56AIsSvTMYkKr6L4
LzLin+NyMwnre35Eu8BpxfOTCudKtsoEUjoGI56VbVB6XPV+baryOOPf219ga4XrF6MNR+BYIZKY
YtVXRtb8FvFm50eR80h3BUT/styqw+IDtEkKFkjWKrGLnvA+Q6UIbFQJqTcjHt2B4GnL52SLh4uU
G4Y14F9QgPPnrf4EDKdRWixpCEs+27TzfPZWyQXbMxlcxxv/vjURQ4l5Sryz0JIF6fAVhWeXkX+m
OnWXZVDZR+13ueZlEmoGi/IahvtcxcGRPOT/lh2X2QiKJqBlO6/as+zPIhU7PxEafaVFiHA1kNGJ
x7zDkkfZEPnnj2jcyfZvkQZyvj6AEIratMX6xSPK7QrggyHccBHzHCDBvW6XISd23c3jdKvEOU4s
3npTCU2rfNetCGQ6XTpYNp15HDli5Eo0cJg1uhNkZpSEWM6bXJ/2cfwDDMhUBUlXeV8lhbS7/B1F
Li/680ol0T/XlG/IcKcPTCVxhqsupguH2iFs42Zs34LkTDaHs0WWaidR24Yq0tm1vh8MHSuxGGc7
HpWrYo86zsijesAujw5ohc1tLKG1O4lCJmeruUauiAEO/cCf+btOKdvTYzxnqphiCn5QUiqkh21c
uWqnqihd6MhAnCAT/g9KChuc4UMrU/NqKkrOLwNzm06CMZw/qxpfwehY3n7/DOwxxyx+L22I9D82
lXFBOmMYY0eM63gsBHwhMIoPMVhAMBnfQ/PZhLolvXcXsJFWf3suLxbMMSA6e+VLGaM7VgKmrvcS
kN2M/syAaBOp4gp1pBtldBEk/ouen1+khCmK8eKRRmGuuqbWE0FRtrt93NfK9DUwb84vmszjmLhP
BsFJopxDX+kP43A1QmRqa7NLOwM/swBO0yHSPShgmBp9XF1t/JfIEd5W/8NM72OvadOwVZjmBGZ3
ltrlwizJNOHEElMvzwNx/4/0zRRWVtrZzXWY1XQH4Hzsk8l5COqYDs+TnIyiXhSRJVV3ON8UXaiX
kdim1G3kuBzxllC/s4+d282/lOD0QyBsuepKGcni6bd9jpF3MRC0kd68NM2978mhhiK95/Z1rgtt
kSopogmqqg1ZfM7Lall1PxQukBcCw4lD+nAGezSui9zcE8w/jNKuijelKlxztEU8r6CXSmJ7Oigf
ezQ39vC+gEz0MH8NHCBjdvRWAeqXIs0AwVByui6ttSwQFZj9E0P3VkytMWx25kktU2VeJZTLHi0l
G5YmvtX2Xndes9UiaK33WcJT/gr00OE7PHaBSi2BN6zvmxEH9Y59YTiQ+Q051Hi4fB1BzT19iC0+
S1E0YlMeoqo2I1QPFfgh/m52+ymi7CNTvcfv8kiTucvsk6lBWL1eRFAUIl0tPqFLtykn2q9v9/YY
CWZf3kwi1LM7/wx20gO++2HKQqr3/kXR9iUqaQY3E565lj5exgOhOma9TSv6oN+kleV1+DRZT4OR
Ua8bBkW8Ujgz6VfO6PkiYj/0vVrlapPDwFGlsbLjnnhcB7BEDBvelCHXMz6S1F14I4YIxKs+P90x
P5W1b3EpwT+7xYbYHaHAbYKp3jX35rbFvtvVA2t77dd0Z9oeSrTRnHKF53y/8lVq19xwwwNUhTcj
CKQFdfjp4POtj/QBrClzvNQKV6UTnn5y923J+Naov5FauHoOWhDhPLdrvrpUn1X+uJk6d7nO6MmO
0zp7y418hllbmwyFz2lJ/E5T4rT8DrIz3tL9nNRt4ELT+FezfszDTf51vpHRv8cBlweL5aXZXGoP
TXzLaJIipUnflFfRkXg3xX+E54IAOwQDgsJaviCPNbt2cvp7kJ7fKo5v3aH29ZLt2+azU7p+dTNw
3EeNzg5DdKqxSyis1rtOqYDvDcXn475VHcIMAY5mqLzZkmOxmTpBdQEhWAUpZLCkz81XCdWCIkAW
+oJHA8jcr4IU8t+9lPQPA6kefxidW3nugGgeifKpWmA7vPhrWHCf6FwoXfmYYkCPbCy0k9oVsA9V
vN0C15eqUcZemMaG+UwP/j/TENOeHhghaXORCx3Fqp32Aq6R0iOV80Iv9/fJNMCJIxOXFH0bfwzd
vS0ImEUCoqpUi+/aQKcsa18d+Lhs2QvPzr1RbCb+jnhlpTL+onq5zeOGka+AZKd3Snqg4YpDryul
stEfPR4E7ge9AYPOO+gzf6cNyQ11IDB4/ao9Y60Ui2A+wJ5rc+b6eYIqchyagbsiyuIjEon2w2/+
KrKc/wLk8EfnjprGuB923dwMDwr+41G9ydHW7qwoO9cKrIjxy8+2S6U1iu3uvMBFc/GJWXWEouDU
Sk8i1/EpYwGwhifSQGHZOrkJ4/k8lzAT1LsTso5R+O9WuvtNFgiHMvt6UgC5fGBNRWjC9ALDfP81
Mq2nv9jb/wl3jrYDyZdnc9EVyufrDW/DIJ5yT63h+oVALdlh2Lhclskb+PyTbzUnTrcOFmnFVpoO
cBBdJdFdJ2vdfe+ydUK2Tsw8PuvyKScmNaR4w41KzbHKfZlW2WvLFbVgDphbbl13L+3a1JX2TsXn
5Nzsq6TkVK/kHTRs8pXjq2CvWock07LYZcoY/tMc7JWLT73EDfMFQYBUfi2YUSxUn2MfahJyXoEN
iNL0mV8wRsHT0mj2/GE3i2Ujd7zLmzU+vXo7UGd6V5icZa5aKuQXRx/IAZKaGyLmkL/I6CnmLhAO
ocxxEht+HvZhyuYNm2brvXLI2nDyuV0Ui+YTswpbAdlPJ4OA7iGtr78XQlrB9W1OcaipWKsWqUtj
rgh0pBc0jf9lX1i8kI2f/4i6U1jI+voQ3jxz0T5ko5r8qfwQz3N1DMm7N1RY2s/CK4UEeRgx0q/q
169pbmFrh/Om5f4fAWlWfNtdjRc6Wy6sc4wz7EroJ/XoYGl18ubY0gMdVebH5+3NpQJqtxyYeTw0
4q+fl2k5ctvFtRzuF5yrxmXlmLasrX41R+Tky5o8JoyavfaLY25C3GIir+o1pNNoixFiSQrPNsHt
uSM2gLD15vToivFjPtJsoPNuDgszoPYPWfvfJnFOqe1TNFiVa9VKW0efLIWMc9fmJxxsgStkIn7H
ksmQ8QFW9x9Dui+cGAV8We5vumbBhNbfez041r7aveiALpp+WHHfZkGpYNWJbZMAgspYpOrE2zs5
xas/OoMWHzyA36h8fFWJZv/K0HDuxoP0dVkP6CZnfy/J+nffLIi4vpY3DZoxsIE0HQ/zNtByodW7
FtPhPd+Kpa82et6W/UrfzK7pQW9WrjTpYQQi5lZNBHJ//7ApZ+f98aIwUmwKXXAlCDOHxvMidoLI
VMBUGe0p2hSQCd+wufbhIrp5e8buGiGt5O2oWEkfU06X2FAh+nJd7xuX0lIsZWYdzjb5whmG71+s
WhsuqHeXJqoIBIpsOHnlKBpoH5ymSu1/JrqkkIbxlPxXxRVJWou336LRkHxxd6mwXrTasYDj0faP
Hd5VWVG7uOjwwQZqc0evgPqqnKFWfnyj7sSNFoiJgEfNyKdElqSIFpERZ6TYmVdwzA1iaKFbxWVR
4zLiMV8ZArh5Mqvey5rGG/wO4D1r0RDwOGSuqdFmUBqNxyeuzf0KybIphX2ue6yh4qOBInnKyv+5
9/MVxLvt4oIuEUcIamqZu3BlSXpolhdPSe7RUR73gcnKsMyyDmhE0uYjuto5fQne3oJ1lgy3hBWm
0GioPRJnQU5Xl+BCkfxlgT5yTxN7SvycOe9vUr6nqHWemEf4Z7jBy7/WHA0OM/KlOBQTH7Zwmmzp
f9VwXOc4wQWuuFtAMujWX5F7EFMZYYtqU82hkvX9n968PdEOJDDW6c5g9FL1jiktywQ3d0ZHOcUw
5mQckFBrEo5hE7L7ch9li+PhTD1yVtRiEuSRDMBfX7idsxIs4RDPkql8OyT+ZuHDdbR4xakt6Sek
awr5WFTXmxjVkkPDD75pPKJXx5AJvR40dEf7SxwnBwZUm2FgOifszdf0t4BoEaD9x/FLWNqmU4rZ
W4C8E0yQ9XekAIka4E9FBIa71b099FrPWhOr97fOywSMGys0da+wf0t6eRjO+pw2t/+TFjUjYzyr
KYF+pTU8pb6MZPLrOJhCu/mdBiTy8TIURFjlgosO8mCIJiEs+scbcwZVBNOIF9PTweHYkN6RtFtc
FUczmsxTZiYrHPi/XsoItxdqZW+CNWwEoHi4ity4Wq356myMn1s0iQykxd88oPTUzZaJ6OR5vbG3
e/K5cgrxrP1VXQzTxE38iqgA4SCdQ2e6fO2VeJLwQarcaLZPCG5GHmBOfUEAVam1HFTARjvzLEU0
Enyj6+H5N1y4Dh13EbG9npG6MUhiogj726yMVZjiv1wu9Suxa2HHSrmgJ2aYlWFOgm8pezeuW6/k
2VH3G6h2txzKWFuH2Vvu+6BHYBruvKKnz/nK75N3HoNHpccpgHXQI44MbcaV+5QtAbqnPeAfqkyT
glFYI/vUoSlR6upiYsXa/ApRmJKDQcvHe2sSnjRuTqhX8TYAVpwTKLA5SWO1VgstWzg8fOvHtEqt
ReriU54DXByfqkU6o310BwYeMxlnDWVtSUXFWsyZzxbi/xk7QeVzcufV1EtKFb9Qiw3pDoCXu4Wf
6v3GAG64buG13dd1Dt1vqKkIN+R15uqe6GyATsrDOOAG0ysFyOCJ4VcpHDK6Z+OxH+xYNNXRiLq2
FA/uPKrXWcKAAqWl4vUxXp0Kn+/iBsv9UVGJRQPz7aC9uEhl574zCBQsCVa919GxeNChyq9I00M2
G62BYEGp9mQdmn7msfw+j8ecylK9uqPlT+1/73BL6JBOTPZDGwZr137U69G8tMM4CgJcJ1o8Dddi
HFoHadaxODjv3FGM7cKcZiey+JPPXnl1oISgg8P1t8qncQgHZahO5spNBzOjTi3W9DQL2YqcGwyh
wOQz4atvoZtlOreeJ13z56BfJSyqfG2dLEapYhCoyE8Ag0GvttwbRX4/nvCk1kT0kxEBmlDFdO1l
H4zcGQX28//iprnln/fYwFXlG27cdI4pp0Hp8OriXRbRXoQesV9mwooc1xf8CEffmZM99OkdJeP8
Q5RWgCqcwjxp8xf/Pr90VYg=
`protect end_protected

