

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MPaacDM0TWg8wcifAVW4jEGylx4PKrqc4CLboKEk0r6t7KyfUnirQwQAphZDsR83L059CNEzB4wD
M8AKmBfOkw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XUT3zAfEi3anHP5UZ9Q64SRw1RnMtcFX7nJsXqsc+jcNnlmbg5PdhmwV7UaFs/PrWKFdgim7UZCy
o9NtHbXd3iHyUEXXZiWfkC6NC5Dndoi/rfKSxw5AtxtcCSaJ3/cb/i40IG38fEOD0mldCmJ0WOZD
xOW9J2aHwV12uWmmUBs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5hB2z6qFvCHrfde+xOJHAAm9Y4Zd5X0rYu4ngUzTSYyHrr6WAc0PuLxe2Zog3gNAv7DFoV1y/Y4U
F6T4flnTjzAqIUvyAW8+maZzCAeWDi8VgmeKHRbLydt/JWB9Ri7GcOoofnS5/hxq8wRCMMkoHbQF
kNzxfXz2j2QXU8RR6+E7pvqcJkK5H/P2HIhS88SnGwppr+eD2lVT18h0s/QB43BH12kpY1JIkQU4
LOR3Ej9QoPTxmx24xAodMjc6qGME333306vLcWETw7evLQ7fHCoyGS8qVr9xvwEOuA+HtAnx7p26
Z/azE34tKzoImCmpb36r638Bv/NLBk+b7agF9w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n2iw7CqdgxuZ5kdEH+pm9NjU5keAcvOSKkOt8pim3KzIVtdYby3hWhnEsC/F1aUQ3kkgfoeHTv/o
nwfMP+AVXxDoH7hATDu0iX0A8s8avaGhFp6novk5xXzwMVnGP5Rbk3GwwADpRNWqzKN80je+JhyS
o3J4z9hQTmce/KBAfWo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sR/mTVuOveJs41YLuqwkxNe6mc/KV56Pt/6c0cIYmcRhmwLHOU3+/VfoPpEClea5ISswKcgmSmEA
91cZp5XMe9E1MxpJldN5YBxK+3XVJrpKIG8b4LM2yC+ZTp/81AZ6CpAKQXOcZAota3bpWOVB7WQt
kPn3pALJ48nc4gaIOk2j5GO0g6BLITkCLwe8Z4XOzYZAEaEB+5dJ58Q/7AbNKHr5UdGO2UVVG5Oo
7GIt9ETizL/sKscnCI3CshbxwDQPtnh9/CAQY2Ci2Oqc2ptOmylUrV0jpazJ/ulKvyLMe7D7sjb1
BOUUkYAI7NZU4AkYW+pW9jcllm96HEkuSjkTDQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50560)
`protect data_block
Nj0FDku/CvamYY+s6tQvBU9M0pkz7pOXNrKVw5+DVidLcqx0N2xgH6Sff2pAHH4DCVzFv90EL0eK
e4cggT3q4IlAU4jj41sDI9P2v+LpNPz/qnCGNvhw2wfvusquIJ7Z0QWdxhjqFaII4JYrpgESWrPb
xy6oUunBltSF/g3Pl61T+njAv4zrO/MgDWnqnSSEAWJtLWZMs9xjoFyltW4Mt0+WTmUF7X1qPoBB
VTa5NoOkgvv22zdOth5v+5IQYqSdrUAVNnH+PazWRtPtBOj4ZtLM3Rfy1lCXuNVjOFdTv0vbsacK
C2oEVX+X7N2z50mZczOR/GGaHAmYjSDebkiaLLGMad0mdWBsCQfM6oSTpqjO8CeoPxtF90piyMSD
TzbqeqNnw3fclIYjwwrDVcURbmNvvFwElZVgwC/mxoAFhj0LoGkFE2e7c5KjXBSPBaXjigNJ7nWH
Xk5xvMaXBMMVTHrUCz+QRzr9v8wVux8KcfQte/1Ao6SIuD1jrgY/oUe0l1fgpcceeuh8cxhfEykg
v+Aukmg0vy5DBZ87GRcTInse/2SflPybRc3pvKM6YciD2SN4JXyZHuIwhTotwydcs7ifrHSu4Zvd
BWWNgLnBLEaIgUx9fdu0tOjI/uMEKaUgVWGUiHpHzQkUrkvhfV9+E0drPKCB5jfBJy+e+mWdAVVD
/7Ua4pydXJIWzJvZdSRfnHlboj3LNYqZF96QbBRP1wN2kvbNjhn4k28kzv0XoSBmgu3XnGhhrtw4
agAcTukn56NYufzuF16G4NSiCmBzX90ulyxSHawOcdZnfP25007NTSXneBZOb7j+vglI0PjA/juE
bfh2VbUkecUdHv8rtdjlz+YmE2Et1xuzLGDnoIvGTnoP2KJVkm6UVQ7+waAG2f9/QPTi6Ajkaj3v
3ftHJQyjuBxmWpYcZcUKzgYw6BAeNkfjo0s3uAV+1Eb1s7uKaaf365V5Obkl9+Y1vT3141UcfmWw
xUelQ4It2BJYK+KlAskqf8OyYGq4/RXR1RMnqIBTzVD+odUqnD9U+fmcuGWz395nh3VEf+Vj+Y4o
gvxjjMbLNfNPLHAhGm+qrSyMbCUalCJU8LCu3XFE1f9o44aq/3T+K38xZafUC4UNl0/2BLNp7XeJ
gu1ptUwYby+Y4BKJAYWEZEga9gWK/pP32+dCEmQ0tmABRPoc8cNKHIgBXMBQkeonn79+7G0hnvKi
k/YhXn5+8LK9nyUBvCZYmuFoxYn88y9kuZpAPkIFI/dKImoQ9KnSQcmuMQNcwpt+TqbYEra2zbve
uqJmcSct844UqrUs/QJVZOKchHe98Ba9peKhV7H9ehJ++wBdeLsTRUdxtn/880O6MpSRm5IPcuYi
xEXk7TvG6UL1VIGHe12MIP4KMJb/1cVvFBn2XQP7wQfWheMc7EecaJa14UZtLqAoRWBHQeVV0jhm
gvfN0a37SxLaFs01KlAXjVEx4tWKoUpsTQGO5E4ek7gWuaRGDWWvY6JTz1wu6n2aCyxCj1HT7wKR
dqiUpRHTe85x+UPh1qYNP9T8UJaHz+X/jCjaa1euYQhYvQfo6c4jpdS9/UomqwAv2PcL2Up/sTEY
UkyAFqzhXxlVvo84JCyEsnatwLZ4fz4OYnf1Z0ivYuUPxK4qrkA1XdkClhDIdSw3LBeE457jZuoo
v34o+bS/64t+pCMOgvP1P+Fm+Sw/SXn3yct4Ramc3HJWjx71Gh/7FCc14dHrPKekD7HDhrqEswjw
uwhKiEK0xwB62uKZoPnQVMs7i4myOa9r5gyrRkCzupqeenTc3Zso9vtgSD/EB5Z3o4lCXQKIYktg
IeYvOji3vEfh8xVylek58L1WnFM3iEKofwiLfvvDxODzLYM3MR9BlWPABgz4alFjyGZc25+4xTxu
Fc5hhTj2gOUl+mGexTh0muaZTRXbIROAHuddruUi2lAGEKqpoY3JlUJQr+pvXjWaPAiWAeaPSeAf
iyF/b5zzImXcINP0L7AIFxF6ySPaqON5QOXAXFmV1FD9RSBRgdEzxT2qodhJtXAv23ItupB/XwBA
jXSYuJDIfY3vCopOq8ux2Wxuyg8SjIHrNv+p7lbQPUaPHZKvrg72p3s9reX4v0sgPMZF+VflFGBW
S4TbREyJILwnNL3/g8aIiWir2YkwkChy4sJGXXgeKspRbTsa7A+9ptcrhIEyCB4wAf+ea3ZJTV04
7alPA6mFvC0D2j5jXAvVPimewX1eAJHKZEjnKjklKw3vC1DdSCGpOyishwpiB1mW/Lmgn2Z6xn4H
V5MaM3ipNAaKvUlASqj1lGm9XeyLROAu09pxH56hX6tT3HTj6iAhnEHZszV/5Pkscony9UMCO/d0
nanmPSJ1iQ4fNjEVBx44kyl0wYZrgutiV3ReK2sSRE1x1gQ2BG8kKYLp1x8li8SR7UcE8w2aSQVh
29SN1gHsDpg7LS557n5ODHBi4Nw8NQhqm11wpzYZmXIqcC2bCJU6qyuE4ZH0ylwWbpjQxNYE1fIi
8ZJzexaZIpMcZr14PMQjhjj60XA+8SwYB/Oqe6Smjp9ohHNrABhzQMwMfnd5W4+oLuiVw2o6+bYV
lqCpyfiEI2tknQzMOVll/ZGDQHhddhI/PBGfbh4RolSbgKQKVtSHEYSXLsKjgr61jY566YymLQyK
D00CYXO1GKuFG5QPPbLw4KY2EgCzgFJlDFMMSA8zHm88vurSCTdwPmZpwyMBnMo0WtKV8KT4Cray
p8BTQRt3dEVT1VK/7xtDDKsprEuSn7QMu4jnrcvy8KF053T3eY9rW4zyMDQ+GmVGHXmZ7Q7hD9Wv
rDkzi/1TjcN+dsooClMz50fGONDGHOaiCiwM8gCfxSDx1FFCpWzk46O3MeAIPMiz9NYMLoursWo+
2TWIuwK91qTzajt3ghm0sJtVuumyT1dujw9Gm7iudRIlMntyCjXDHF3Oqw0r50ZFsZZMP2eBfh0s
e8IFLxfJY6V5azII3lw/0WkGKXzLNpUz9QHsQhkTOHxn5sDFPOiQth+exi/+n5jpZVfJdwKkz/3u
R6fcMXn/L+u4W9w1RGYwhRY0JTZME9s6og1Ir6d0ItoIsXrc/kiX414EPqBL3aX0Cy1lFDNAfy51
qsouzpHCRmEG81DnEDwAtg+1xtOCZ2JTduuwpmOgjKFGAYxYDpI0uufSD/liVYhB9OvZXEPlkA9n
M/WmJjVBxg8E5fPtpixZP1xJyNzoJ4FJOq5x6h0nYf0SqEMS2VIyIZBmoR+CXI6RPAE+EmzGm31p
0Vlgqm8LdF+oScwKZaUtKwc4IENETPYKgmnxGoQaF9L5MDbL4wr4sK5JMnQE/Ae6m3Vlv2lEBj+t
dMaNNDzceOkkWJoN8qr2PqOWVByjeJgJPrrwM3p+pf+Z7MT7UhJHfhH8jvB+wsKhWPYo8DEziP7I
/QqQVHQFDft6DrZrzIjfNh3al1qlVXhVSSiyxAVmOkwQh4IfSE1F/T59Pg8WQ7IjSxuxyFH/QrXf
Bhe+g6PF+4BOFKZNZxrFyA6rVwhGFVjrK7TB+RoryYOohan+6G49KMeSXvrC3vtsslFmShEoxXHa
YTNbcqUCsMjwknb5nGWmI3FIlvjm978vgta/eNCBKwSmSxHFJbhxHSGWC5tSvoGJAb2XzJ1OR5+B
Ny4PxBZBKWDwZTvFhjHUiUDaHM3H5Eg3zESHJZWpPgXWt73RfDfA8rDLF8fbUAxWH1lZF3HBBa/w
OIm8mrH73Fb+s3AYMjtup2M1Zg7sLd9SS9nfU3NiJLpXJ517jE3Kv6DQQh3rfxDi9k3zcxoh8QLi
LsNZ/0+vNqizWI4mu1Yg0p5/nnzl1PiJK4+jB3lyWuozqkSICh7mwmtIC6ZwsjmKirR6LrusRZA1
wXu+A6wiOkaU19eUhamWI3hcfS5lB2HA1arlcaHX5Fz1skVB9xhxOnsGqvGay5S7vJXwqmdna0Xn
PhjZKSey41uE/ycFITIrB9Vr8ONbp+q2NtTeQAUAATXJTg2ptmoDqeb5qs2/S5O8omO0rnECrSEK
H7GCYkY3ZQ/AL1yDBQKfMKPMHKlYCGCRsy2AEtHyEdZ6TeYsoF+zIL4xTX8eSkDZhGK8er0bD1cC
pPNyvt9CRFbGaJBZLDElpOE+RncXqA+BbyUW1njimfroM36dSsfGDBuH4ZIlPDRPquKwgtH3v3zc
xfDBdI6FNjhN5TKnf+yAQ9dWNb+SwPHH5Tkny/Zo7J1AQm1+fPWbZqk5nocY+lAvt4F+QoihafwJ
Pq7FwbvOZ1QBilicP/X0NppAT06uua0jixkarnCErTXDm6UwkcdshkDMssu+s3WU0Hjlc4ujgBcI
kEB8QfGX/V8ke+p5ZENWn36jeEuFFXzJVX6eLvFwfiH1kP/NIKLERJCeG3GmMY4CBvTI4WvR778w
nI9MipkXNzul4wNeasI4hOT/O7Eq52anwkFoz0YZfmoiLLZUNIhP01PKsF1c84ORqZAH0YvVnrKM
lonVe8coeeGEOo64U4Qel7ldGDl544vLqbE2HZ/V5Op/VvVcvuOXoZLeRZXZChKP6RlbAaNpGL1I
vO1ANXfg7MQCMrNRCuzCIynyH70WS7KEYT0gj77PUhr6/FogA+zGX4Iuoq3E26bct1dPrjX/zDmq
XaTqHI2LiCVH+eVlj4PB5GiYHyS9sRWudsV/2tjTJiOuFHvMIEu78k9VmQmpdQyxfgucLy2mGbUE
n+06aYkjNbJ4EAgw12sfT8vRv3I7I2D1Jqmh572/hfEg88UalDbolSDRLFieQmuwz5JHT1dUO5sh
z6VD8vWNdEW9/6e3Disg1kvhJMlB5fS217nUzNVWmt5RxX4mKCuI8GTmZy3MB1YDObtufTwGHHEm
RDVdJhy3JC9Ldy8kFB3Pbv2astiauiZApCwaS5We9VoGBoAN8T5y/QcNVN56bBTZu6vO6dU8cA8u
A7LQu2DMgxVdQCrq03M9y1/vsMU6BL1LHt45+YzN5EdkOFwEmH3yWjQUo0NWcnofEERQ9p8vM58q
oP+/IriD43NPvUj+rQRF426Fal6PDp+C/OvHWJ2Lb2qZ/IWr64ZV6oXLpKY0B7gZUtxcT8dpQ2Ig
wQx8D1l9LaNqrpGm6GvelbqlzGhESGlkvoM8uPgXd1+JmLrjudWoKpu5TVHZZbLLRD0AuYPQzlSr
3mb0xw9sgTp4jy9UOD3iNDeWXUJhR13ZKjpXsU6ShCpU4Hp8MGg2+CnmbF1/AMfZqzIMlo2szWLm
LEBYDON1cpt1iqPT/ro2uM+0vBZZMjQt2SNdsoJt5JfEWtqCG/a8Va3vrD6SGoX5gM6B2KSLljPc
sjnEj4HeFBthpQ0lBdhkLenTU6IuvFMZ2eByFZ/V7mRQZpBcbEfz6bXOUDxs0QyT8zRVVjmnuEHq
uakGeMHbeZ0kQOIAy6Xer49d8BkpSSfwLNUHWKkJiYOeLuK1SUIjQKA9OZJZ/K3qhd6L+LiiT6ug
5YgZKZtarfyyETQNO/ryw0rH7W8Aj0NXnOk2++wE56QC8Mf30iKqkzukMhLJm0i/gMsmbFxppk+V
3ArbCrU0xbpxzJDo70hX3sSsbQ7sJuxZLHb1dB+4tpd3m5Gbrzsv/oczfFjBIXEKbxlb/opZpiba
3mo7MSMBM3BSgF7BD8FbqTIH0lmNiJUg/nJWfN2Sy6V/XBWAwkf72Sc1hWKwPHSnsVe1MOSfMZfX
cryZ13wpFdNVJgtCCKSi3Xmhl5znv3d2y5Gj8SIaZZ8paPOYJObQ/tQBhr6Mk4nlqaZbDZ4L16f3
CCwSvMYteFL6FylZbx5wIoCFOSmI/UY3X8ab6CxflfJxgkxnTwaNz7iDRg0ZujXcpcK68YhgI0VJ
5YcGonMB9aNxaFA3czJjkcOZ5GXU4oE4HyyXqBIzLroQwnZ6zmE14nfRAvJUuFAZBWtKyituNWK8
ZKZPyD6JL8LlpfqOMd98RZlmyjD3F3henvVf7iFl+abOB6x+5TVDaOF8TLUZoQceHnmX3KuttY8b
8XhFnKf1crchJKR6vHfC+yuSHoO65MiRGDVS7GTODe0h0J/6dalWweWuMdptTlxamUaj2XzO33UW
KRUydwyzhA+H3t1ZMlGpmuZ2VCxVHXbTmhohyW7fEH3uB8kTgRUuk7/USnCQ3cTuQgFiQUYnDebz
33u7DozyjZiCvho0P2m3HtU+FN6bNI4HjCYlqRd53oPVecPrbQXmQl1ReR4/h5Hj2zs5IICyrrHh
Vew50r6TW9ZmnGSdH6gWMBN83TFjDfg98DEX3XN+SDPhezRhW8v4wCS7TMcnAzVnIEfSJBs0BCcz
lPu2tOakiZLw1YYLBrn0DH38zMwCdwjgF0vipymN2/e8ttkrQ6B5LM87sDTidjPergIYOxcaAyph
ZCSFRpDjTjeWxD6NfFgbLwp75Oeg6wlnonfFIRbS1vrRGX/CYYmNuKSrq2U1s00D39iSDpcRw3x3
370D81p9O9ZXVl9u8hy46+Z74ryl1easSpAYtHRVqnOeunyVPgeA9rPtKcPdErC0svj/ypzlsbWo
zNwBE/MT+110Sb0fSG17dEiDyT82LrMVNLhofyDFkjH25PflDNqMVeJMPHOueb56y4bDEgeRyOUX
oWEAuNuNRhMaz4Op/SThXvOg1esdyGrmWy/w7ZQofSS3Qdy9GH+HPdhb3KLI/mEGz6DTVltAG8Zl
ELlgtzkw8/mMy3mzphs5+X8LWm/vgkhAH4TfRBVeNuf4zuebncIoLkJl5i4G9nCieCBD3Uc278aq
paAYlYwEPx2FAUErhiKOz8p4jPhcID95lRrpuSRlCU13o+9yFfHL/rDi2fyDz4BuvxHfU83hHCQa
zTYUKEjwlstnfdDchZGlnqqzQkyQJEl28c4dhsMeFrWaLauWuIEtrzXcZjsuxpB0MzwdkxtjlwlE
eQxezTRaz6VacTQ6aGGFNlWHjP7waXY6+pJlqMLAzUnEwPE7B2sDj3ZIegp3fnjaryctS9oCoQO0
oJ29BJdMMjqt/hF/GQSLNRVyNKtW4h+/zGzTf8sXniHTickoJV5jg7B0Ji5d5WExc0F/iOB/spzN
RHGeuKGSoqjCeOJlfsBiGJ+W28bXlFj/EVq9jMpsyUsvdpFCBeNM/c6fmGLDs+IT85/hCIaxI32B
RkdjSuOfI8UHMjVxnemLPe8HbZFxvTSmRNGW4BdBjCxLn5SOXSGBqC9cbq5WJWPMJSGca87h0N02
ijYeHricboUElUUdgQMfiFXPZtEn8JqnMbL/a3D9mVAN1uv7ILSmlglM1XLpUMvehUdgfNnoD9n8
6va1+qCGgWVLBXHOCeJ/uNuSVQpPrbDO5noxId9oa6iFBLa3mRKu27v6bMUdD74l6xTsLiUVpMRA
VxIuDNuM7yhdNx5+pH/28IvOqwHE59fH7L78dyIVl3og7V98fc4fOieaj7WoqNTNrbUH2TwlDBnl
Q6ZhQ8Bv/muDtwfK946DwRVhTxElq2cs8C4pnvwlwr8EIwRnyIkyrbCaO0ouydtSa4uM6X5tJUqD
9tXwC7SmnLfwZTQuMdfaV0PAqtD3IXADwxxowvoiRLPJIuqae8AHNa4ZGc6LdE7qBE3AVJ5pvIRg
s3tnVkQpLJV/MRgQ4nANXPxx7700CdzJq+nOtPECVljzMl0JG0TCWXTPfqJG5+iBPUDyspIWI8Pt
1229+VUsk3NdhX1Veua+zgo9HXTez2HXoxf3YNFzTDFOz+KvfkQtfyCOJEdWKHlbRZi/N5B3lIG6
uSTcPd1OO68dd9uDGAdsmFFUx9Ls7OqIKA+9TTWoGhRcMrx+SnalLg4zXk67CG157C1PriXfT24w
g5ueW1RRp4GGuVsUXLJzpX2M0wT3NhxYJxWtyA6dB13lKHmLIru0PZgRqdy625cYMRO8Bv5GUTuq
XAHx+3NcTdO/Slaq6gS8uPQkC9nFCXd6x1y7ieyhxrJYQQC/YC9H3Cke/2cFcq51XCy8ucz5xK9J
pBJb5YaXZVlBGrOI8eTPPRf6vdYBYQzX6/NFYdFTkEIhXGhg7wzGOw4RFCBDUO4KNJkJJr5S98ar
7rs2JuTmQIfnvxv+D2QlJALgNIgO1WduPe8CtT2znotX17Vjp/C/ltMxyYEOcwd0uAyD6uCLhXQ2
p6xUkySPXxXUFdW/xoDAiQnvOkOzxosTOJrYLsba+4lOTI6YSjsWBR/VSRPp/pmyXA6scAtylW3a
HGp/n7jTEI4bz59413NY/wkbxdE5uSwpWrDVw2eUVtGDYW04Y1QYtiISIdwbVHJSCHUkPxiYHnZK
5kfbLpAfkme0Es6e1bCS2Ek4TWv/2py/54j+c5QfEevS3U4+YLFMnvlkX1+odw5ljsJ5C4D9DWha
TOzC866U4gTz9ZJxh36ELe0qH7Lwomp6ml0Jow6On5AoT1aGiwIncvh/tdMcGoEbtzWB1/J6bNkD
dlpff69YNx6Hr0J3muZoT1IJR4+NKHvOSHD2N0mKS4mj4CYWM94D8s+MnhrLEwRTQ0w0AtIzsQ49
RKVNl1SyV2qCs95zcnTS/3ROvqE0zQRNVIv3VW12IY1U9j0G0ntEW4DRh+fkkECvdNjie0CRlMia
ZzVzOzYH4UDQ5CVipTkOutA8gw+AdTpRxA7lfjx6L0s1MInFh3qBfBPFg2Dp+5FKMLWz9F7h/mrg
gNjHlraPfBYibRVNE59jYka4XZIooAe76Z/DAsl0l1rhKOQf+PFECtV5YmBrQLafkH3+nx5gi9Zg
VXjshXt+/Z7JoAlJqcsz/LTLmoswFJRagnfz4skxeNTM2HK/3/cfAp7tWL0LgtoKV5Luwe8819TL
2lSB+uTTO72JbzJ83tN31Zb0yEo+ooUuomtErvMZzkj3LaEuhwvqKwBdj7mpO9phoy6MPqlAleOW
1vNx2R/j2WxkqL9flWKbyvNrc6dMcNWrx4RtqarGtXPEx1FjSlh1v0wuGrH78xdUGmns+umVNxtb
SJ/NMH98wDr7KrKC9Rouzlw4Uhfpr9YIzHi6nat9Nlu8vVzPzjx4y+hVrobcbG9sNsqUsnAkk3fm
1c7/QFlUA3ucSwECmW3e2hOR9BljvqQ1GixUuP/QjZDIkPDcKgtiJtCjj1bh+Yza6CDfFk63iy0Z
v1SN62rahA1Lhk+GDw2vQ3F8dp+z0F2IEeSpwTx5BYJqQk/YmPOsHdfgi3B7Ku0JCrMj0xx60so3
vozNmIU9hDzxbfojirayhefOYbS5dG5/1o6TvKIjYPjo/diDH9Up4IBER7VfxDmbvfSyi14HQYpa
txOXjCvEz+R54NoVm9rj9QljTqDb/xdTiGkFseDCskZCcaDPrkhB8XsrYzQCKKv44pX0A+WKUtGD
LZuFmoSGhXppIwg0WnOCD//VbjG7L+nxXdcLqjke0IIA+hkDKf66DI55cTGNvjDFU2jucadDT8hx
LreUy1UYlalkBg4Xw2bxgYxyggVNIfck1rw2V3KPUPGOn5IxvIq03/5vr0Xb9Il6CB0PTH5SMw6j
AY8lCJ34QchkWilLX8zQGdnkBa7xrp1/QFWQ0L/tVAMX92xCfn375cVwby67AcihiNIID8P9wWmo
RNY2XFf3MHEE+2+SwW7odAe5begVXISX10dSNndA+2+MW0YImXNNB02r0Xhn7bUAFQ8qTHXoiLPY
CKkxBPMTwHfijbXJbmsiAcLpZ9gQCK/u78e/cNca35em8s8+c/EeTmzLL9BbA9UUnBRHDWUIllCv
6bw2CcGwviULfBQENiCdObkxEgB2pxcolChh9qbbNKgD3kR6CWh8/l5l3fONvcjqu3JueiJUS4FO
XhHaVsvt8mJoLFtlVIwBDB0hyMzdl68stsM4JzrFQlaSiPFrtaK2TEktBv2FdPILPuwHOanG8vEV
x+lvj72FNeQXhMk9mvR8GHliFUt56ZuNbF+hAHxbVw4Y6nCR7G/Ez1fb2yYIP+q7xXT5ekKZ5pP3
pWps00Lz8Nh/GTW9M1yn2lTZ2IEqI7v6uhGCFFiRweJGbx+a1vaAKWx6SpuxNv2VAX4d1agkASXV
0H4ZIIFWcHVBMg+l9lKtlTtp4lLOFKN/Lca4RXHbg2DiGTg4oT3+8mkVHGaOZ3WqkU9Jx08PdJ+P
nPXTlfSwbb4tUOWM2Uhec+n9WiMZuPl55W8lhji6Mg7ctMkvbKw6sGIuxaqYLoqNkuDAfoKSp7jY
l/ODEh4mLgOiESLgandPJl/ofBoCkMgb3GWV9URZw1QhKSe7JeuUnptI6TOKB4SDKr43Hg8v76rW
w/y/06K/VE2+/f9459IGwmQsAewr5VaxDSHFfpfv1B8EsWhez1Nh00d95WxF6rD8nj6R2+y3OgtN
DN6MpPEhHpV/0YSQ9xOK8cRF16KWiXkADdzJGnrEZK88HpJAtoUk1CKZA/QUIPi1MLS5RzvPbPA0
DXoTLKxxespSjDL7JrUx6+ODbNIH22gWAXpPI1/4k69xBJIN0Ij53RSiQazGasnoA3hGCLJUFgRj
sTvHRSOcQLyhAH4lnHMxf8iO3TsLB1sopt5krgjYNui+Z7xcB5gt6m5nxq1aNxAGVo9ur58WUDil
rXz4L9ba5hUjGL/nOsU8lfdPDvAa9YzXeT9JE+YwVVzO9Uwz07ZJwyYnZhjc+n7puYJArfVEfgwC
QlIMVZ3iOuzZXEiCED+MubfmcihEZpGTdEcnv+hbvTY2wBViswkMXu4u1wOyte++dOoo9H2iNWv2
QhdUIZRtQOMAbmcGthIvVjJaK4FS/XhKF/q5AKlTpH6evsk/aDLvmgHdhY++4naggmmyb4yelm6a
HNgfeY4uOShy+L20D+HW7mgGKk1d079AmnXgizGkXhQKicwfsvhIxV16DUdhVMdjk6jdJj1UFJxA
kFMGmvflPK+gWnPplIxzae36Dwp+GU1dynYXAzbjNM96GoZruzMK0PL9nuiPdQZ5SUMR1fACHRvC
J4Am60/qCqQAaFrxqi3CJispX0MsPbO/QTaNXoa5UqFgaLChTAGqJmZKzz1k8tb9FeRM/vVwfxpL
Jw8AouoSWuSSmelkeo9QDNwH8Tv7kWLDWQWDI8Xyp/+tW1T1eTyBwTmZu5fEwIjj/tt2gveOfXdz
zFFBRwNYXIkfKIk3rVNTKtRdjYpDJQGQGM+4xmbfZG+txtobzD95DE0jxiEA4UdAAYSC9BYLGyc2
tAnk5vFmmusrPPDcb44IWeL+MHn08gae2dCCtncmFLtS1HCfPfJTd3pIB+kaXsfy5EdRSIXl+Ov0
B1Fig5tp2XuP5zfGsmNrtbiVr6iowLaA1AX1dWSLKkhe8zSbngr5Ut8T1ohtN6ELIENtYuDgRUvS
4xWtOxIb9ylVWv8+m2JxovwZ+PhI6IgHrkRYXerwh3VOHxy5HcmdnSNrto4n7XjeLvGnLQp/IQA6
NvT7XgSu98psdNXHtjS3drMIDB3nBFDLIR8jFH38SmSnfTtm1ksQG2MxK6aMCVPAC6SnSh9YdJyP
J4pdag0SAjT08XVFMCe52yLiEcMLpUtOLMwAuwKTwlswdyDIFpVlTNF3mfQoQX6ExAY7qHMLgmL+
Pr8rXyWNixSU9GzLPAS/JplQ0X/8x/5EAyq3FmM8KUUgDMtntr7sFJa3kDtaJ9TKSER43hO9dUZg
+D3T5xUd5tDL5MsCKwC94tPbj6f0597T246igfAONFn1482OT+Ki1lm6PHLFBkF8hNnnY32zifAf
L0X74fLKz1YrxK5m29K6ZH9DHQ17ZI0PAx7zSnCLRbSJkOZHX1o23rNRAPcsKpODeXFVVomiUURd
CnztMk4tfWvc79L+GXC6lyf4TMQHsCzwjLjS7DTud9FB3oJ6fn8W6YXazr6Ys6l62tLhcMEt9d/k
7H9Yc5VaX1ce6bXZG1CS067vzgJCCY+uJN7Izn5yPXPUyQRtiDiYCMJtrkY/hvaty3UDEeFULAVF
Zl38lP3p5CfvqgZ0RYYGLGS+oFOC9PEdqkpGPJf9rXomITYnmQ4D7GfjZgviGx2o2oICUqqU5gzA
Ku86yFnCiNYZ+/sZuUymWj5Xk8zEV6XUvsKHzX0YGE2ZHwybdcTCXoTif0EBRsaCzPFgHfT9/2gR
r0MtREPX4zZpR/MrVCZge1SCBTcRvj6E1XVpxOd3DGDtbdZ/LtM/shgmWPIQHx7g/II1D7t5KUw+
1Eq1VkPxmBw46xZZC0xR894B8vxbRSahNXPRPd7roqkUoPQBySkSwLr+vg6G8LnX6YgkLxVhswG2
+aVPiRw+j11bjzbO6EOBgHy9nlp54yw3CPTuQtl5133wj9t1E78I1+jcQnCKCC3Sf0AEXk3VoZWz
UP7Hmu6+h6pDUaJeLPQDG02kB27rskb2H5170+hTuHZzUfZjtz4NhOv9xsxzT5LduQvKVugtUDtV
SZL6q7ObiPh2RnldjKk+QQwbsHtQ+dTbXJKVxwcvvRUGIn0aJxNowMOZS5S3arwqct0G1dFiOKGW
bqgQX0PHyJTBPz5is7or40fPvJbmdZVvvI0rH99PC8CJpYp+UEqzHObxzqUtczVAkOT2Q0r5t6ez
zBX1uCNLxN0K51huT3l+BF5pdFWaPhjfpGMvkUJLoTJ85s3/nsFloqMC38OAc8kQ7co+HWKcH+qv
7SP+NFxwm++MzGCNg1T4dziDHW4KGY9NyXL/TvA2EbU/mR1KrW5gjeV/jnOInWlsi/66cYeZ77XI
iWzi7CTuBzl4lR3CY8syenWfrqG4mydOY3uThfHcBHvm3SUU/y+caerfBTHKvsP0o0LIjqaMhE4k
SuXJGPKSE7ONLAw35O/tJB57V67djgpshzvdVCaOYcSprGvty9lePjrJ1xp/tgywaZkQ94GWMVvM
Dd4SjI92H3JQkcdmX5yyqkeXUVSkaXifP4vM6A3bBX0GH1nWKoryseblmYUh+i7F68z0SQlRK407
4VTQFVzhTT1EmBHvWbTIYm1tFGFZbGshAI73XDuXW/LEkxV4jGiZ+CrSD7fmWakDYqvgwy5Zs15k
NOyX/P4QnmyVtL030ljt466qOdt9ix5edgvzl+4p1GJnEw9pIcIksudpetA1E+VJh/VT97rvWUrV
iwxsmqmF6FihBaWp0ReeebsfReit22mDQdHWQXm0urIH68ZCfR+lMNYkJGIQdnsr+mgdFmF4lzrY
m7cFjQn11OwjnN7zq5GQ6wl6oxLa66arsxh2mhx5hB5DgzAbdH6QPTAAKcRUxRX+M4rwnVolZSIL
/w4IgRWMz+InV6xh5EDqCn4VNMKGj/oOMRXbcSbvOsyC0HiXS/IRucH9AN55apP0bTvqqn6dkjVI
t1zAE83cRPuQvxYZhRnmEKlSEyff05DEONzAUYv57aratZYDDUNtw/0egb/JN7CFNYeGZ93QZHdj
nVm66IYQEr81A6pPqyTv7xieAG+uGnfd8JbhurbyEPBm+QVGDkNWlG0JR0Ei7d6NLRmHf/CeoThJ
od9k8TrB7bNc6XRH9jE4HEPEreWqK/eG0QSEIGF5oPqx8ONwhzPK1Ye+wdLEAbVqOIW1g+uosR3m
uKFT13S8hxETUJAsN7GC1GtoR00ZNR8T+67CuVkJ69tpD54Z1eyReRKtIpeQ7p9161XtKs3O+r4X
jC+npvyqjkB0FJhz44ssn5AfggzkdY9GnoS5eRxq32K4rORVVai0ZHVA2716KgS7rRyKhudgg5w9
Mo71PfC1hhPexgftH3MYVSAtOsfMEqewAXNVdA8ujQbJwHApk36yRcCaO1QXHZEo7IgOnkdoadLn
OQ5Y/fp6pyvgR3ksgY6UfcU6cJIgGePNqRfv6Wbt9ED25Z25yxg4hGCmXDBtGEZgUTH1U+z3s8WI
6PTG14fTWzmd3parLjkfgJpxlgq+IQ99+BlaK+r6AlnBz4mw/QPzbR1yJT+vxqnFZ3KPZlzqc6MX
VnW1wK/FR1Yk5qQtFG1S5j1/726KttJexMVHzBcIfLQXtN1Mov34Lmn9C691tKc0oG7idECR6tnD
d6B5H8Y9AZqFj2/n5w6z5X693qALKNLOXraefu/8uKH0ONkPy7FIhxclTBw4hcuiUD9Oo72fRFWj
YjxZpKgCZ7xWCmXzlQMT1P6jUSQrBb90ZeNdWdj7dfs6fz3V5KyRxLGNvCIvh2gEYuVGILWOVBn4
dCh+9QNJzUAuwCY+xc4UUhxgJN4E6nkWn2glXH92hlfpOsS3cSes5c32laWOD/GF1OlweNGcwqwd
Sg0Qkjq4wP29BdozwiDiDqyUgYWl7C/mhJFnttxsBhGypQUaLf80moOl4RF2OXnJsaUYS3kteECd
F2hy4H1T9F9FftMnUEcdZwSlI728Sxp/s60eOwth7GG3HtQbJ02BRLH45HXbee33VPBr7JYTFjhW
ztwkMqOauuTBRYCg747FV/4uLA8xs9IAcJpjjECp720CKLU7wGA4eBu+fxECcwYyPz0FZg5tiw5v
xolC4Pj72mWIpCqR1gKhxRtfoYOrAm0J3IEovERxyFgUOCvkGlJ9mab3eT1rrIi8mFKxwWeEZXlH
SkgxJ6H45KSxJTNKmFoRp5OEdhLt2SXUg1K+fHzaxyhR+2R+5XRVqvPEmnQz/pAL/yEkjHY6txjN
bvFq7TJQ1cz6zauvHgrVHWcdsCxoaRC4c1/LBSfI6J3I2l/IvMlZ57g+VVYsB8YbmtIlBqfemwq4
EojfW48DLt/qSd6N1Oxqxd64wwL5FHHlEUkDPdQ0+5uXNqnlFaHVCQ9FdQTEz68KdszhAJG94mKy
knrLCKCbulRDCXrj8H51PLecuDxASoI0Wc05TIZPJYht4bjgfjC+vi1YILFqH0pS7TbzkAEdfoSg
9DZyzVjxz+UKfJ0e8hbZVXHJHrLsSdj5PRBbbtbMo2Vey97YqY6+TQ/YemCHLE9KrG3ymgSA487P
tNCzhVG0ZmJw6GGN1UAwGpMGZRXLF8CF3gt3/uXC+hY1tHckZjZw42wh3Mby7nNA2qlgU0ayhcA4
5J2YwWEy+J0+5VNkJN3m7Va9y/kJToaoArBCRh61t89l9AwZ14j6lxRyyFNXxd8vUBB/p9F68lN0
BRdQ0xvhJRjT2ZbJkADALRvTQUUBJdCRzaGa0HsB1dTla0ofmiFATmmJTUYusjiHCGXduMe1o2xd
7bMHpVZ8YS0qd23TeEOt/GATObFvtOihx1KV7AIXUpRJ//LVreTNG3+P8a/uOXPkoweRSr+02UgX
BXA4AoAOATfNYlZY1A0+eUeYPguhco6hgHvkLhFh8s9rLnrOL2ACxqONiCkBFGFmoU/TK6PiHHdo
AwsA3ANWVBXWv6gpwurSP94igzfD1S3fRFrl8BdcsaRGFvMRSGBxQq9K7yZCY1lMA8yKblE+T8bt
KLz4m+VuKDbNjcrmJPr8ki/nuOzcTcB8o0H5s64Nr/lRcMlHovAi16jrciSo0kRclmgJtRrJRuSg
i+lT4NtWylEET8wUD0sdVBmHtoZdhbYflFyCPmRWRrtqjBqSsIUlAnYtNcdLwNh3QaUJGFnRYTvD
MDR9wCuIPLaJLzAma6BNzgWe6HKxjdrI0L2fLat5CZyXtWeTD7e9ZTXxZwwXDAunY3HrMVIuSO8k
sKdPP/6cYA5Uz85Cyx/lIXtLmCEpLfK9bD89Nka9l9uvTGicIfkigoNWfIujKdN88vR13rNBK3nD
lMINTXFspoPjx2/P/D1srWDA1qxap0q+jLcI+EMdg6VxaIMvA3gzf7laqrFgiO4AcsKGNmaf51DH
V43pUDPNJeOnF2zlIyMhhtGZS6rwX/jMG/8ITq0+djOMBG6pGDKPuXtxMiphMEmGEBz726o7a7m0
yZ3XIxWnzFEZvDWbkeswsruDh221jDkaeEQzyDVfJ5zE8srfdSc5FsPmxnUN1AhzIsCMO4mWefeS
NIFHsYqU3KT2qcGZt66G/3lpdLUWfiNzesfkYMaCr3HR/zXQdZy2wqZLC3qBH1Oo6DzJxkkc/nqm
6Jyf4OoLR12jlV0HULzIe88B5aZg38r7vBIW4n4OC37KXS0Nn689Toe6a+D9ly31084Y1n9RKqYM
V9BDpnM5fTQSAS17CiyY99ajyy0ZqiQLAWBWHISZvI1wsdt5e2837T7CrHMQy4I+rDZfrfy+z5pL
C5ZMX3KbbbBhBDD/6h+ktVDSFgXYRcbysWrg0FaI/f9MGcgCNXREpmgpPUKdxO4Kd9e0YuBCVwzl
qy9lobTlbd3LE0OWCyRD+YNTyr2gzmGNS5Ia8+V/cO0GcJ3E86fuhmF5GhDyZlOfvpxbrOqNeyCj
2+i7qajdSOvYuEFdbp2ZzBqUQOeKl25+BdDSDoYUC3WVOOd8E3W6mFHvOuLoiMbWa7s6ZLwctcnt
Y1p/zRQ5Z6J18wLcKNCqAmBeSF1sY0wtx1fbJuYnYlg/BTKyidMry7eNCLQRFoqCrj6EbvWIiQGg
SFtGioZhPb24rgk2Wq01KWExeJdZPSsuCiXUhTaO8xJPxjNghmijH61qbM7EgHfAhL5cAdfa7qvp
EWHaFPAoWiTarBRu1g2PPWO/Yd7Dhv8laetXAMkfXGjCbvp6uAle4JxQ7dBUm74RJQaaqkIrKGQr
wfhqMwfDQDyaKHVmO9lRWJ/D9Akl5zlwXq3hZUHt8PjSnmm327RvjA8cMf84RMqflJMf9mVqtVRY
V6lMnMdDiAQJeRH57MiC2C+WvWwj05XhYb0NumWMTA847K/RhQJfrc/+1ToFVss5xIlaoDmUlK9h
VoKMzZFlEg0H1sKHhOac5myT2HDor0jspnJDNF9S6rZbw/axUM8UL1LuznC5/7adQZlTatyawmJ+
wjWHfPKgJYP0oo0nDRr4899vukUGvpEY941eD2TKTd25CuTLtdiOjmhu3Zvsm3m1b59FkVP7Vr7I
z/zWu/9mpkwT7xqqETw5YPNTUPIVUu/A5ppnHWb96g07DdW32M6AR4B0+dvdZrkEnYxsGmt8Blto
c049zESkXaLV/tSSVO361u58nBnMtU08TZQ0mtefswx9jiL+D3BGxcH7vZM8m53rMkxBh2s+iWHN
c39pen7jMaCLKTYCdLfEQMOzw/Sw77vJIpBR2LbDJreC1m9kUz1Sa7UMOIMSNg2/XV+ydosInnlB
aph35VhHMPQ7Nw5HqzeW5vUB1FNjZVlgGrKHR4EeyKk7Y3kAEd8rhA5N8y/O0Vy5eFeUnEtsMS0Q
WGyod3dbkps9JjNR8miZWeVSXkZ7EXq7zXYYTvB81n0evdgNxIs0ZXECHSlVZJTCvV3JdsX6T3u2
FVkhYIV0mHLSqQwjpzzNz+IGoju9tu7Pmmq7JoildVlCkB1dpLhst71TK02qmGt8Qjg2kEdBTAm9
RMUPGNfKIcY3/9efNAm5VhZgYNdVkUGWBtjpEGKMEDD+/edde5FrEbvfmqCZt5xJ5e7xZLZQa5PE
if7wEVUyEWWZccUgllhe/+hjKitd618StfL20p9OUNtOCDHi1p9odeKUrviHQRD4sCgHQyIoS/Wz
lzG3TvT5t6noXkDXtgyDO1O01xwCQfqmKSoFF6SQ7NP5xp7Jau9+LX9RFQR1Qtl8Q51Lrx8jtLAn
jH8Qn+9KvSew6FkEA/4WkrlvdOZuFgPgOyUI9OU0Kpf5fsGBHKvh+OQxkYdp+91htfg+1HocRStY
6XTQdBiHSwfO8BCRl/Lf3OnmOGy3IY7lxML+xIWLVm0PBRo1RrTNVE1FrRn30gC3ilixL/tlqXLK
j66C7jTrEpbgQtydhUWWUj4+GKSx+APupqpFVmNP2oFQfeQnWLjgXSNWmgYGUWjYFavObn2VWlty
jT1ueaGQJKK8WtT5ZmR4NUv7iq96Ez4tFgLdHNlazNLC9gIONs6b6MemaPJwsoWCKWL+qaj3iOe3
jvfTpGxfn3AuFLdOih98oMAFJZs3ajKZ9BB03ASRhUVT6tuvxgqLkE1Z34JHAvpr3rDrTlsRLJHG
AJ3y2D20FOLm97fbhJp3Eokzs72h6zLtzh5XnxzoLqciIF8WfCTF2H1m5TQwNg9534o4Tjwtuiwd
fKKdGHt/AY3gTRxksAuTqjP8b6bMf0Ctsr1bc6IQltQC9j8qrK0OsNwTGzRJWzAweeiMnxRaIThr
agXXvjPEawIvHIldlhPhLY2cY60ZDHAtLogqhGW/0rW7fv5iMCeu3RWrZj0ZAFTO2wCxGhbyZ/eT
TcCWmca/Jdrg/SqOanyQsj+YCGyKqDFt1Ry8yDDIa8SoZ00TJUCW5xG6smq2U2BxobTeuVXzFIvP
2Ac7rNcnv2rnFaz32eG6PGq2Is0le+SmZ19TnGQEv0iAMQOldpVgXoX2zP9Lp/Y8o/nVOiwZqAhy
7OCqqlS8LoKbM6y/+F7g1b9wKohRzLaByC3NeFNuUmipz/Qkg7M9RomzSk9yAXD4ecL6wq11U/Hs
RvkqK9bPXMSL/ypupL6/LSwg1eo2lrFSh4eh1IA8bx9+ZHkVQpKtywhyYjgqAhtsBSyohX0EdHQ2
FFK79pLoG0Rn7IHOvaYDk//kW8vqoyTBxHzhmVo7qsCfkR7d3s+C3KeS3PAkcsKElIpWG5VeQ8++
sQgPBqssSX4xBTDhBGbVnIVnKMf3h60iykjGl6S5Atct+gEzcwKtv1PowNlA//RRe8Z2mCYX+fkQ
taQ71DVx+bP8DUlp5ra0J1xw2zdLIP1dIfw6evUvnSfZTkDBsxOkv/mNbAgtiGY5kbLI03SPlpzE
RGjAKvE9OPfHHVd5uZmjh+AJqUqAc93ktoVsFdOsMMe+skb3fjhQdFOsNXHMx7LzbxYoHo7XjeYz
k8iJ4grz/KrelGj5q4iuYhmQ9oaRnxMn7rR2u6a0eJHhZMOLw/KhC6JD5yEKxfNzRiUykBvVLtu+
4ogy3ygHG1niELbKwde9RqOUtAZQ0K8rP9LrPi+G36uzBXv3CHt/YN+1AeOPetweUpd21fB9j6wE
fNnS9Dpaf/zw8UchLn1V4kxsQFsAqmIdjAyX6leqGJDktWMuHlvAC5CrrxS83jjrBIXWVSir8yXV
tLvzkGMhT06aOyM78HFQL179FyU6+RRQJK9yEqmqRnP97THr5IEJ9Ctsu0D6knrk35VXAq1kCx+d
u4vM/gS9fKJbTCqm2qLf4nGj1Akapdk6pfH6qvslEU9UrNkqhcJ6cuZl2hu8rErSFSVIRjGsxnF8
2L7CHBfWzorIbM2lJHs7JjPUFUZxNMJ6Avr0yJ56VgaWRpmXs1wJqmU+nQIm8mXwpaALiRfbVXRC
RAkkSw+ZQHxwpbALy656lbzdYwlW2x5VTS1JNf8nfJMb6/iSM2cZaizt+7chHGBZXgjRXuoPwPV4
OKauWUoZD3aEVIDpZz1W5U7oyckyRjYKi9jWh94CwQZiI4tPmVBgsv+hh7gZzeLH0y9m0iFdNKzP
xZWgl+i8od1Iag96iBh9ajxx7VrgMaleD0NqxcoU1axXBJM7fb21VE3LqVF0cZR2lhf2be4Qr+D0
eYAiviyxnLRkRpv92wiLGozujxKG3EsyWXlrdOYDf+IBaI3ZEgSM5D3KD2VFIz1GOG1M7X+aQT9P
3nXgxNwByobX7+Pbl+JsiUOZyV3RwmwPvfjV6jqxza8cUHsgCGOGW73r9ozHktkYZ3HzP+VkYjMU
HsX0VAFJOu4tBLiBhlAQ2gyHAcVWd/c7UzSHoInSznwcJPy7Xyjw+WZ7cyOjpX626mAJjazt61iT
yS3VNBVNYBLIwnd7VuJ+ntvOIuRC+i2y1FMQ6Vk5jr1uRWBK3HAY319iH8AGDldo2MPtkCv4ZIbh
uB/Of+u4VADeoxn9vXgTV3SM65vST+v1fF1dZM0KCOWc0TE3fHNP9deIBhFrCyY6rUp11DBDmTdE
LdCMcg2QERHiv7uQW6RiwvOBjT8UhveW0kn8jIUCEeTa9UsXR6hnzk7+JOQJhKNG7RlUV46m3D1P
iKgWr+7zF0asPAz4FFEkLGOuSav7qoiYs2dKBWrmKBAh33xeVenhLm5J3R0J5h+dnUAnd2hZuzMi
v3sB9pN+vs6RJLTrGBxnZr0Gg54LvBvV4dO8VoLPZV4ot5Afht14pOVmlq6v+SpBomvYZPXxhNuP
riy2vB2kysRfQKmGTQrAZQtSNbzOJ41/zlqy8tz3zwOHMUo87VjMXhsOK8pPlHtHfdIA5Ubb7J0t
o/6vjrFnjHMuxIx9iGJ44DjAhEBB2Kc4lNcY+XVwrlWwJB/lI8KVaD7MoIn8WVLmN5w3RxEaBGWc
ZE14VaKa2ybG0NKdSgRqQ4LuariA2hZGfw4d3KrFWlX7NX7qGBQTSZIv5kgaEZHPxYwnniTl9svn
u3rFbnRMHezRKdYAewbL2KI91JbToYjPQXTPyCpQIkKQISLx0xTdPsa0YCQhwQBiz4DCd43S03OS
RIegror7PRqZm3vHz4VG5pM+2iOudhKjaO41IJ6S0nk7j9phYkMCLOLILW/m/xgiamqE2CRfNDm2
nxPczP5W0sy76D2epLbQPcbajUYdHqrUrRFK867XwU3KpYpG4TSsEhltqAdI3fJ8giar2knOuuuM
VluTuxacxzv+Moa7bMkyiQzJr2zwxHrsSVhjOpBJ/1nAgLlVduh0ZQ3EPPKUil2IRJ3F0KbgPhDM
CHg5ZqGcykO0sq+Vm+4V2B7d8HX8vsLTTni1SXWfQ1Vz/rqzaPdfc4YHhO89cLzj/YPucBCwgT0O
73ex6HnBLBEy9nA7wF4OhxppFzFgbQwn35tGRMCWqtJV+0GIi452JxbF/HQ0P6lQnIOsbJfXcr8b
pD/c16sdAtEvaFSFYoLHCnySpG1iRxKEWAZddvkhS87Ym0SuZUujT8nY2ITYZThHSLMFwKStrlpl
U+SYI+UKmDcM8smsORnKoOboWmTm31rcGqUU73ypHs2eXWphEO7Ho27fvzOiftWeU0Gj418pgpqB
Wolb+K5D1NhYQV7UWMFPRh+kdvpBpVmD6SP3xA8PYINdImlMBiJQOs9z/yl53XjaWhm56FaMRW1V
LfVszh572/vP4FaTss1cwoJUUPvQjuv2sO1M7Zv6v54vqA7Chn01hf6OGnFhoU9FGjC4nu3hpayH
2K4EVjiCW9RILZxb7i1tuguDbJx/LyN3l30aMizu+FEcRsO35uboLnRZdmnmMa9PLzMB+olMcpO2
3j+Ssx58YuBxgMQYLwkVI/G+nc15EBbvxvQVOZGR5K8fdDsLzICb1g6UNp6dfgOrR/DzzB/yNN6R
ducQETKwT/+kQrJE44ZGMyxK70ltACdINIpeJacc5uJuzyy4sLOftfzHz83pHRgnOiNfdC2AAji6
BmjYo25LY5mtgHhy6QPSTEdXV4Ar5HKEiIeocACk055Jwhh5469HVMOWrnDJzQt6vf1aq7OlwuU+
7W0cn+lDkdx5wAw37BK2BA0jsBNlErYQyCfj86SoxzHAlPLLLrnN26PUOiYHBB565Qj5eneLs3qt
LC88WDTASxYwUyPAO9waObQN6ibcRUbBjBdt6hG4zT50nvrb1QhB+yzOoIqi4+IXx2PJj2z+07cb
eBOwP/622X/vDqc9mHS/3ovy1HUugY47lNobkRBW8NzADS2xoofKxpZbAnHUEs1aVV9972e4E6ey
7z9mihAiVmv1dRvq/nqttJ6oWn8ELo/xaTI5pqB0Z2qS1nrEtq8fzBwVXvfDX74bVShUfjl+8yF6
7lh6JJjTmxEd6+NfrY6SagTvC3/Lv85YFuISKZX8PVhfS4NDMBTxVHuukLeYys/rXtdO+kZ9pYuy
w9nOqflQNB7JtwS2QqJpGtJDBBMe3vxtEqrjLyZBuPXuvrMH9ZkTSL8WnLGPG2yakQBuJjgn8KZt
pb+oHUG5JlTsrCLYuOL0+Jry2fZV7ggjUfuVg7wPuqfsiKnxJvA11FkHu0bajRUcEeRTmUjzbN86
1J5+og300bbaXbthDAAr/ASLVJzeIEVYANd2H/nCBTMqsGZimuJrMTtsD2eGNVllnuV9RMLkORG7
aaLjvf1OeljXMIkJ/4RDMDjIxeJsCdzsXkpifsycX5a04q14x3Zq7g2SB4wqU9yJ1ybhGPSOqVjG
53Nj6VAchPusw1MK+667jM5mDS5Izn7wuaOkpavSMpzVE1S3Behp83GnX5qAjO2UvF1zHJjjyrLf
96jDGjCMcx4vO8w1/+tqza/dIsSWUViXSyqMLji4oj6mk/rrJo9xHIWUEtnVEqO4O1kQZTai+s5a
tdKfsz9RLEhVsQII7L5MWw3CIaKSZvgZyom414ImTXrGskMjsfXdni4LvgZGp6GABtVhH2xD2flD
LC6y1aPJmK2+UZdlmsjbilhD7xRhekp45ztMhEHDwaTOiynsXvMdYoL4RTqyfcXYPOcJclevAP8t
jRXH/fDtSv8aB5kmzf+bgDHIpkW/afZRH+8ll4RoWuw4g508NkmRRXfs2bwqcmJNFcHdtsLOPxur
7hJqRtJ8EbercB+fXG8SH2gjpvtxLzdmTmJbYWQbqalT0MqqEXurx8OANb+zHwVBRRLYEeYE+E2P
SkcUsjCfdM4tD+CmP9vVl8Fhvw/xx+3x2vPxJ0AZN4xyRDkdhJSiuz2mEo+d8UByHyhIJa1/lFQD
UpSU+lMH8pU0jdRmiABB/wgNAiGGoOeNYe8/4u1cVh5rjAi4uexk+wbDHipI+z2OvEngwLGU7gbP
ibzU6i5tr/EvQLbljL+82O1ilEr782QfLnqQjZBDISZztLkZMmQhqXfLsxN7P4noo96MCBPogQfF
dfed2oiSWEkHY/fVsewOnh50Ep6BgHPF1np42I0iLJWN62Ku3MnThDGVxZpVZqWzPcABuIBQgUXy
gszM4ZmqmjjvoOADlS3NFzssY85WcFl9lR6bVDQknn4fgQRnJUi9cZIWh0Yia2f5y1wSJCOfS+UK
I+mdwqLftj5ufaFp99eOv188AQLlCOQDqKYpmZGKm3jgMnQzQfKTui9KOXpWXQTNhTl1TGiuyLZt
lqxYNz3r/wE6BxWGxbtgts0RXCFm/+W3lMT58rQ2vrEcMhsQfIn4IZ0gXlKnIcinLcYdqlg4w0wq
PEWFJJ6nrjsHoMBrUHfT34JC2yhVCt5OfVSYjgo8feEwvsLCklU3VOwG0Jk7YTeVgmQDsC5Vjrn1
jFqhnwqNUhYgo5fELkkWR4KiQ6n3j9SR1+/GOK8u4GG/CjB9tZaLThd237vZz2DlDx7SotJYH4BU
BDHSUVFmqxmjpTFH/GX7Sa31GX5EF0TCwmQwXL4CVPpZMG0KEdEhgvMR4xlrV/l54gxkr2bVhqXu
eAf6OJo8hbOmtD9db32ogNT2CQQxQAn6kN4MpV8CfGjTU7ObKiEZHG3NYLK0Y6r8zMmOxS1U4L/Q
nQGBx275+sqbJpmSawxLhNIFZDlCZ2ZMg8DwjC94Ls/nxhd/RXaJfpE/OMEwxaDCmL4B06mcBJan
PrhVFZDTbO5ghXtt0I6KjS8MET5KUWzQRoEHuO9GHX9zTChoi+PhAj/7C7k7XpXM06BSOaG1yNi+
gp97tQ1E6DMeXJRHa6P9cOTrp3EHndCfvFjAhltzaVP0rnnN8pOmD9SCRylkzXdFAlgONPTd9fKQ
xpapTU+V4dxZ7a5kHiNzdzgF6Zj/V4ntTT75kyZ5sC31aSM0KMYOWH2KQqf3Jr6C78hrQonANla+
2dUtazWj1oE1prcL2UwPbybfO5vto+TZLpLwAcc5hBQryE7wEX/W52jykVdrpYbrrhlE1sQQJ2VY
XBnFELnpJjP5ytpYH1NtJBXUfYDRNHVUgmzC+M8CPM/woc8eOvWjI2auioG7LKri+zVFu0kWaMKR
Bkjk3NKhFM04jryptvvCMkM1O9c2/irzhpdtrhcZBEpqqDVVtoPjP5Djr6Jm3C3dc0q8d+aZ2OZF
EY8bSDFmcn+KmcyQBz+jVan5l+kREOMBpV6/DNv4/QvT2oIqa8ryvrYLFRg8D33Fn1Kn+AMfr+bM
LoIOSF1IeIMzuXec3qGdeJHWkCDx373QiyQnbxveX381tNW3YvLPnbaCJyZuhS2jceI0rbscMJxq
3CfHNq61cykT/o0vYL763N+Y3WE2zNtgkosGcLYySqGuYWrDc+OrETUk7tZI+sYy3Ul9umtxcNwB
eRXIbffN9or/2f6n+cLL2fwhSWtcCA2bShoXyU8soxbn0Ks5ic/Cy65PFytfB2QGRsK1IgJMOvDP
dqNDUZk1lpsnRSI09Hnwduks3VXpF8dgpwyYDbmc9UU46qtjmxw3WFLfXPOGcY4xtdlGGBYuZn6q
oPlcxI24rAoui05jBvdBT89qr29BpCe1vVYXMAKuP7VsGkTcthriICJEkGVl94GKT/LI9zkkerSJ
TTUHQbdzZLu9jrLhpkl+dYrH3y1spDPh5bIbT9GRySnCgil1fot+PUSJVHRZcb4EIEa1bREvx3AQ
gqJsRc28tMctOtH7HwoSbSvE/ovLDOSXLFIaQi5nIp+wMrnU58ZQo32SZyM/2Rwr6KR0x8hl0I4p
rSrsixWc8hkLxfVj9FMgrhdgbM/LRGhoVWtRrs2o1PAgoSk8b6ALlJzcPNJi6mp9w59Hv1DJTIYg
/UV0V19GCNe89KoiY2JlWntl0hWT7R4cuZ5aJZxLHZE5A3PH0XkkBfCoWJFWWYGaTA8+1KxFHyXB
6qvNChbq0n1pJg4WxxAfyQ0ixLHzLxCMLkkgcJ4F7k/zfvfGTmep9O1xVAdp/JD2BWtTvTrON/eI
XMYFP9MrtbBd9cM84sR7pJ16l7OnZ+SinEpv1gMpMM7dwvT4cJo2bmPewr+01x77Ajc3liuy6zGT
8yCQZlduztGl57boz8TFkn7G9fsj7NT9o57RWLA29Ai3y+6hko9QtxvXVSs39pP0UU/TkDy4A/r+
+FrAuRpf5LCrC3g5rhHxRTVmwc34S7BZilz/VSJWCsld/gZU4uxPk3l/YtjELJWVAtIbVJQEL0Rv
q4HSPbYuD38MH6Qw0xMX6wJ0W01LRHOfpWjOcjRz1NwSsqoE/7OjxJCuM1xMVEk62O06CYgFInbZ
hzKuELCFYPAKrNWiR1RseUUr2S8U8MvKNwoZXatvszSSzBqFeXnzLmtR1AIeprZ64GDLal10dqSp
Ailw/yxQUFAw+wzFh6FPL1UKgmXExZKtMPAbM1eJqBJG3/JX3IUVz4Ri4Baxi0Dc4eBhge9G/Z/B
ABzQBQrR5zDdjyN4J6HcILcxtRfuRBhXshz3mZbvMQO3nA7uub9l1CO00IwJr/wBxQMwclTkHLPJ
U10GOlrW6Z1s9/0mQzMzICWBrGvk/xoMDiHcnSPVt49qt73G9nGNb2hOyolRRdRSfFdaTGcCEPYC
SEFn3Jk0gW54MyOMSrt6nObKYVFfU9VjwKV9eRUTKbIJ4w861vMaVFVx2IG8pwxlqB2hEphXwn2Y
s/j0dt5JupIAmVT1yIXcbRWbOZUWPBjVJnAwTJYvDkzTytdP2woAdMMPMcCc/lgBoO0igfcU/5DG
lxQ1i2rf4RKyW6NGLIe9CUKrq6rXpDloxCS0DxGqVLQNLPHW5h6Qjc7V7b2jMnLNHc2x2zPLQWlZ
yQTXBhkzhccdd/HJGGtERY1F6InuX+dSj2zO3TOk5Ql1E73jU5uflwTK4koAJFN70nvW0d73mGUL
Qp+Tq+4NiMbAki71LR2ZBjmgowQgpKNaCm311hH1CVj1R+VGHjYB8o/5e+VkaDw0rQKsn6SzdWXi
CuKko2k7NqlA2z2OlP2Pv08SFdOWA4NZQC5bT4rT3mnzBzL+IjaQhLVm+bJP0AOESJOS+aSr69qT
7iHjX5VaDjSSMqk45N+qEHhS7C3daIou6TTQ8Vq/9GoU7ssghQYdSjh4llrx1/rI3yltN9tvwffr
8JiseZ5+neklFQ0xrvYYK8NsbNWj9nUXn3dOvZfHnwCVtnyMUZOxqmMf+oBs0GlYLEZ9pfoEDpOf
YFIKjv6D4ixhTSt+Mc9gJX4tqaE7rQsnLUB7S8unwe6vYebl9ig39hAuRoYJFPbLNFsny++4gP9d
ZR2mQ8UNSKU/tUJIoZUAgxCBSSTDd5T/50D+kDhItSKWX7H16pDj8w+hB2lmi/jH+/LQ9DEgi7Kr
kBIcebc2ddZD0SFAp2D2+DB7bH7bia3SSpuPZObweAl8NYfDXRlKnDe0bO5sXoa0hafN/OXYhafd
RcbF0lNWZA74x7yOdT5WSooT68QWaXlBI4bCxlK3GsX2VcB1bTUIbMEVDYT3r6RZYNmfEm+d43yI
gitgFwXi/jh1gHDVxT2DLuyoNznJpsqGz1sTEG3D/yHbIIKwTR92DEJF/50W5MKdlLHUEnPrRgn9
SdL3LSg6GhmYFIKXxBRARvfZrHtMY4mWQli47HZupVt8QgHE0TmrWMZBwlWvivX6XQzgXBVaBsHQ
beQvYvpXFp4BK7WISxM7lXMTfGx9ijfuspP2gEI9LSWdBA13dGAqu2sozOpJJMkgj6N1Xc10kluy
STEd6GEMs45iiNoICE3qK4gv/GYsUjThVo+NGitvUgwtFZUB+EBc4GpsbUAsNd44hPJmMYnphN8p
ao9eRDszFZ7tgKZpSYIwJUOhiRBe0uF9h+ntGUwtQzAwRUBR1d3zJAXGKOvtW6PNt/wu8n8SV1X2
zwNzHKA6vUrW6LODsnl3Hou/mzqNkMa6KFgX57Eu/5XEOqUjuITNXSNi21QYBAA0/APRh2zuPzsU
LS/wLeMVWAUKVwdDmru97DSvX1350hBhooxBp2NraDNZykwnC5Mj9Bp7XRSrcfDmfs5y1u2/5GFS
orqp6/qYB6KFEKZLwbiMsGSnSlOQweRc+hoyPzZBeMymBm80JaMDKTQNymLY/vz2avvSi3SZ3x4J
Z85lt3KdfIqdSYWq0ZAZ3llivF4aC20ir0QbYkXSC96oYz/BNvKnjUqZlQnS6atIWgQOBvnGxx+X
dF8tuyLBTbmKhmak/oz6rSD6nX+MAzp/J5IF+IKMMV2PO8rUOnHWGMvPakb345EYit7a4rr+5hdC
Y7v/BxrYOau+mqwYs+wYq1YsWxhZagx41PMQPde+RHf6gqAJ2ru5CHbVXue/kKkMi1Q93qMuNGdu
VcQhU3zpl7B/VRKup9pZ/Cnc5Sl0o/BBzsi1T/BT58arhH+sdxaygUfO7NQsWrItF6oFjx4DE+gh
AaJV4mmr+tNMpdS/AOHt5XG6dyF6FEqIKmSGLvxgp4DFoNTkzNzE3jB8YU+SdGlY5gUF6YJdP1vM
aM1+90Kdrcb6PtL22/SGWrQMtaTFho/qUhhyTgkdn7s8ogXD9LgnfM4kYU8jy09hNRY4akq4vMRy
57kcQh3ZKzhYs9oz4FZ8iPqFH/jpXn+VAaAAu01cO4IW86M/6I/s6FG+v/MV3HIaBI5h3/YE9umd
b0QT6UmW6f92qrh6wwHMCplzfRP1uZ77A0ele8ajzLzIgZxZBqBCE+BvZ4hUNFE5FG9zNNaex5UK
A+s4tCLeFKsjvk+bYemP5pY/ENIpaQ+vD0SuCGiclHanVJPfiMR6qd1V3TMUc1iJxWwWzLLsXg+c
8pxiUE08lGoSy2UXgfw03pgdfeYdNwGX/4rUajXxJ17EsLqA2usxE0ybFER9sIEcKEaaOvMoln7A
rXYo8uzkUV0xBMzCD+g4J9qCu+WbJYPeDE+IOEWKqnvh+QLUqHDRhdKFLYXLLASlFJS+NpiU8ue3
iaU8vo5woPaAel/f7PYY3BH/WO0UuOazxk2nDBaoVD4SGWZgvDY5iFFIDoi/j1WrD722G5qPIIC1
rovUyz3L38FaVPZUY5o7T8RARVHNloPTXOkm1JYcfZa6lq3f+h76h5hL4K+eI5TyzWtJSiLy6R6z
lgKq76j4/NlXlkzSLeW1Md2IOlEHufskwcG50aEz+6+I13nNuQaUCDixhskDJuNwTR26BrStFXc2
fI+980OKOR5NhC0q+7syMRBFg4JfA//gK7Ibv2X/l6ei3xmr2zye6XyR+ascz6M6mXRFZWCv4wRT
VVMOiBCsCRkPmEdjc6yJ2wSNQEwa+voytmHe1EtFwQuMJMHVEcqhyeNSMJl8limdVUty2VVOsstU
j+yM2x82P3jBusmiE7x1qcN0bE8HuDNj9YJNvYI6lnDxJApiVY70HD8JJ3ShFpm2KzYMdKCU/5rc
uM1qnLPiAnvdoGQNtyZq+iHFff652u2wGqqF1RfeZtt7lYZ4ZegceaMe3wIp+nLmtmUDapd2xGAK
Ffy9ZDUG7EVNGyhfiWIRZgMLF8dEN6nas6+x002eBjNw3OaUQEOq5LvtzvcF2DuZew/rzITWxN/C
BE2UZ6l0W+RnE0jm4o9qGmWHTNm6YFautJlitY6QbKJH6JAWl/dEw6MiaY4abOGTTUhiN//YsxYy
k/BXQiVA3RaoYF4Un1V4zrqKgs+h4uYy7BLNSH6VIYJZAqpGVGBXZytIUvPESFZnRmYA1o4TRE50
/1ONmExWE8aNQVrbCH+TnUzdTX+Cuau+FWaiJGEfCgxn+Fbz9RS1FrbmKcHnFKvDZ3+XC51Zbzx9
gOqxnvk4szqq02r4OORtuyk69d/F5nhxFRQbrpl2WAronShwwnuvmkTf27yfwQo7D8zipzUDu6v7
h8tkZ6VbM7/NgLNI0IR0UTQ9V153YHT+plK/FeqLABgb1EUIH4OXKOcX3v2xHK7EGf1ANNLLibln
tqC9dmqTDU56akr9QK0ib/eygTAkoH2uJYHTFiAnJixUKZmXw5EP5FsfG2t0Q3OKeXmtCxpegzYS
zsQoq0jJWo5vnQhE69kTELgomd315XtYbdyQqahKmS3enAYWo8AMuEc5dRJGGLK9Q5dKXg1BOkV8
R/hj09Mu+ie4BWGuoaihM402zIc6X5Jr+eDvO5bbl2pKRyFY0opxCEBRWcujLkX4hrk4vtoW/NqL
osKoFByMtMwTDgXsRaV1W/hFrUco7NgsguIxGPkQ8GhYxSrC2pCjvaF2+aSsFVKeVjg2INBHnOW/
9BCRPGexoma0d+BnTLCWHd5h+2VTDJR4d7vT2FZLhVKfoN05gg9jKiajApQxWHs8wfPdjqgHp8EV
h7sjkYxvLuAecJ9gRbtrpKwFie/EFMS4ebIF29gL7wSQJiHR8vw/BjmcWUAWn9pAj5EW17HtER1d
woQwWqJ4FajR16uxqRpGOP4bHF9lXAuLjaum9OVfC1LXSEglQgi+1zwA7jdn3ISRrsIEk3i4mmYQ
Ztcnc+K8ad6JX9b1GXdXUco/Ftx9k7t6rBh8+M4IGtXnnjYpFmnULftDun3Pf7SrDCeq4wtlaED4
h3qaTm+oM+NPXiQ5jZcP4vhOnXjc+IrvqxdXjtzX6SwqzBCXXwrwqSmzrgVG15xIXiebv9sC9agn
gDbP8l9iak+VerFQk4jdVIiv6TvppWLvYo73G6sqrKkY2CDuZJfFiCVsQOfMDb2qh4gSKuLSuOkJ
CuxIdlRBB0eniIGUEDsw1vigrVnk5VVitAviuMBbBwRjxJ6/vfxrqFI/SA4wIAzvjhvGZ8vwsEsY
EbMzGbBjMVQL6V4LqkY81+HfskqTOrTYN9n1UcjufegbabXyRwTkVBS8zmdDaNeg4BDh85gPrPhs
K/NpEE/Aqj3ptgAhce8tq4Nz1QPWHeZunMTAjc2Goh840bqO/xLezS8nJs3lcWUbujRFzYRVkHRM
zjHzfgass8U4uv97V4LuHUDefirvKm874uU+tTL6dhNfFn77RKPTR1/XJgqFw5lTPqAHSKR2vAZO
qegoPFYr+lPt3qkVgo26TGb2IiDA1xw5ZbdO5x3jpZ8Trhh8weRRhlL7L6D67LVeRCa+hD/b/Shz
jQMsm+Jn3IRNhxMwg/MnwgTOenFby3DwXzfmJY77tmkyZpadWI/HXiSPgTLT8kNvmfrOoD+6cTmE
BTkz9IemSCi+OdffpOJGDFtUJtdM6PMhnRAh60HhatIfi7hOZREh0gTSKQ5ZTQ4KmyXpBy9+R1Kj
n94MoYxr7fU6HKvv7f3IsqdE/6LdaHkFZ3hWmkK39KqPrnNBmLGFM7vANOXbMYJ26km4CSmUpjKy
dRoAj4bcIyEyvN1l/eFcBZELgFeFy/s9V6jVevL3vbyQG8g5XXZQ+ZZU253ub1EZFeENc9uY8yt/
ub20WL4basCwQp7ymUrkKwJJAfre4hhVWZOAuKghrF7ChUcl7O5Zf4Tl+1aW+FbHZFOm06PnmcSI
X4EnDBDoGeWFqV7wVolCH4GpUPipnGQqucVjujqc9sVfBeINh8nL/YoYtxY0VihLDtSUY3weamKE
e3wwDJhI7pTdGAFjy5GIgU+XdOAhk9g3gcIBXVmn7fc+Xe8VMtQuJBQxnKAJLp5VP0OyVwEH/BVU
qNdhNpC8I+1mxyaNK4Nl7mdFl+Vsnu7UXFcc2ytOMvjlkt2UpTLMioJkhaITzdw7UMsWnrQpp5uO
Q2vkZTH4cpfsTWaMTEqYoc4asmYvP2HoWnFLEefEKND/rvxJJ0T2IUIphx50IJMhheO09C/n9kv5
avl8eNBOzl5zeOJf1+UNEiagthlCxmgcqu7WuFw4nI3nF5C2bNQB/xW6eh4WSe5bEx7iRxaMesN9
/CVnYoK7ccLXL7SMowip8RvqN0WZ9Jjjre/HTgdSTYRYu0SWbYJtps80eZAxCu1R2WTvQO+pw5ni
heFpljyGjmZ9xI99XY1fiiZ7yLGonie/3yFz8rj9DdyHz1O9t5A7xocSTsJf+dIpydmwFehB2ei5
TnqV+daxR+yaFhRZwFkE/gBOOoQzmuiaoFvZPb7VZ+zvDOKpcnesayGMfvlsTgazaS4DPzWNrASX
fJl6K62oDom8JJXmTdMCvCukpo9mcCodDMN2/KSN3rraFv6BBui4sJYDJzvSEhjCbPUZ5PxZUS1D
oJakToI/bEQUIZGeXV2+iEpTRYUDcVHVcoLdbMKhI6KlR3OTGGGarUnVsQgfel4ZDOL92HdRNfJl
6FSQFjDVYV6CN8bvCR66n6YAg/6lv7bxI4tLGFWDe1CzjJPWEyYbikFo/f02NRNF/IPlrMbVdmRU
lE3aueWD7oiQ9iZ1m0i+DidfzI2vcSfwZAe6VBe9CsnNLh0KTTRsrX7zoFD/PIu/rMmxL0uh4pCk
g4oEVB52DEHch4LlL1VmUDKoQmlnsjMslYHa7FvBxu+P2dFYh3v7SehJcyatZ1JvKSHzYRnT919o
j/4JsnMQ/pZWZS/Az7OWGTLmL4+hMihstykMmzwpExSPdMqHBVcZ+UkTXwwQjLejR0JQ5GgDHk3j
MS3fzLZcqD8oiEpBK8itAZJo8NeCblGl0R6kChYgV6PNQ97Vl56la3A3I+1/RXy8pMl29AGc+8xV
DIxFvK3kxVv2+8I1gaGxkSILr0g40K8q4bHb1CoY0Ds8cauwt3FfyTCMsEAsRXWAsjDbadkWoUWz
VsbIOlniLkwb6gd4WoDpbJ+JTf75mdM6cjBxCYiipC14c9TBiT24GNJYTzYDB351UZiP1O3QvIau
ORrl3nzbSNjrklGqLkW3yuIlsZt1LbmZ25BjWtezttyn6II1CKruEz6A2aEh75eOXzMPzOBnLaXL
3BirXXcL01HieYTrYYwjhjpBRvzKaq8pIO+XVOh06Zni6FcaWL+jEN8SSaC5p+9ebBCrNR6eAVC3
uUT7AGMfqNMoPmFAzWcq97PXaytSPDn88FEL6AKkzbRza0XXo1Fz4+XV+4ZzR0ccDkkI9i6Btbk8
DdlVD0aH9rGRFDqOplXoMqk+/NrGANkKv4DLk51GantQ50dOAejlWUY51pBwMurmn32gcBBiCfw2
zAQCXQKPqNM7qcZAqEmNUJBwEnDTyRamDG4ZYEhAbWGbK9zpVJoOlxQVqe1Zha6Iju3H/p6O+8nM
g4yaNg42Fwf4dD6dfSCpfQbAiU/wC0zCNoQ6ohaopAUqgFQJ4Z88Uac+gfrkeVKwKvfLN9/zCDPp
sf8bTEpmdAdy4lIjBCAmzk9pHriBlAm+hm3IOkI4gbaB6KDYkyUU7O9ClkKjTzTg9/Vc+Df42+XC
vf9PSCHRazPa6+W7lFDWkcbuH1hqGhzNZ62u1HREhCj/pO7n+/GC1+287oVLLq0ZYzb/QU0NEg/D
yuy4wrVhETVcW+50yz0gRD3PeU+4Ur4Pq6nC7HxRrLKbF6UrAQSX/x/WeorLbpDdpyu5IU6yx0ch
doZciniLGOl1VWD1u8fd49xxRiVcoNg+kBSLjaomphE2tHJqFq79jELAmgQBnU9HdoWBngOpsGXr
/j4T4ei/rttquFGDWyl748K8lN21ByalnV6SdnfQdi6hGacvl375fyReuuPie/kKfd0BSvrNxbEQ
NgNTs9Di7Ewt3P3wDFn3/1weDitfmHI+l3zKvZWhtC24XzwVpCeUs1GBgHMRBkEZnEbulzRowveB
Y2a6ZC6wwrWavq98pcjpPYWOSGV4CZbx+pscmNAZxNki4hJoIcjFSvq1nqnEyDHJ/NBYWdB9ABrx
ruOFHDQQsS4e5YjWyBX13Nxq8xaEx+Ro8UrNqTYXmLF44DaMisO+yt++HK5JRi9z1UHsuVUI++fB
GePVknTXqMb70DRwaqQFJH53dAp3iLwFxPE49nx0noCWvHZd0gOHygMxZbKQP8ZitTCyxVkmzGwd
fGbLszSMFIab90nE946vk5T2Uxp1MtTRbvQW5cxT++AigCDO9R8pU3DIqAesE+DfhQ+qTIkTjbGG
L9PLK2XAhQEe9onlF4K+OXsbc35VA/WtYQHADZ23Rg3JrEr3FPtwfY22tdZRXyuYSjCF2jGNXmGU
6XGC4gy6aBdQhHUIa0J/XbdhwOMKhQnl2I+xDXu+Tu7+J+rb/JL81F5z+N3V4etDmrrUfbgSk0ut
gTiTd+m0SI3CHY5cXg0mRyRClkqCwyV3elM6mIjIIgkLbNeLdcNqSqcQfBAbylm5bOpHyFw96lsa
bgL2CREVAQEHcPF8mNGxPldSnR+wRT/v9WsYdTWjZ6OFaL4+2Ri/DPjgKD9GyuFfz/5wrCsmju2f
TMHJNJXpRlt+hzwC431sa6xFK7d/x3CznTCTB+bX0CqKvsoxUhjkdHeqeca6lSqyGMjYi+k407vn
BtCa+Nn7lnq8OeCp2gghRea70U5AhS3XEz/2H2GGgAHU5fqFVY/Yz3vXTR7sqxUxWbjbfDPKB0NZ
gQ3gZqdmJLrMqUhJhgpFYoOr7PmkxgkGW7TVlEQddiY2DQWG2u6QqP8MGxGm6I/l/y23+EAsNozz
3joJ6oQ9ojVJ453fBwX0IIDKXoMjZk1nqb9n529RvL10PYv66Qs3CKpJaIcKlRSbD+NMo4pyCHao
0lHUa6VY5gE3xUri+Pxjya4WvhP9DQfsOSGNtCFTykWZE8el1c71Guy2Fr+hnnppsG0e8opeokqQ
7CByivy/ij/YWPh0zE/FP+SYJjYVGvgq/C0KR5EvMdgiGlSFcCCxfI5AJcIyy0EQS8RKX6VXVMCf
QNk5gcTDjRQGq+/f7vBzPEBKrzmZoE5VNVjvq4tx+MBhDTXnvp2ciwzcSwEuKH8jskTmqxbdBN3/
7KorOaCc0mYu1ZelQ4u6F7fCbmEmf4Kl/Qw5xi4eqL4RQyIYMUuU8+v0HVd4HSS1wXkosEHG+vkR
BWZ8qTMjA2eWLAnompbWJu3g0FprXYhepr269dZXDXwAtneiSvyY99VvC6cj9E9KduFOqUxnf1TE
DiiEWsVjZf7QlWemkl1O52W2fV5S/4P6CzcFxSIRDG9fzhfJQqp8HBmZEY9VmbyCc9IkhT5V8/w1
UOZwpQHsBDCAQ6OLyyowSBzYqdSl0y662RVPqEPguPnLOR8lAAG+9Y7M18LY0AAH6kFsfPpph0AZ
u3zm8AeTGpd56tKorl50CEX6Rtsw0UASOt6gjOCaSnQoPsDAMBY9t5szsYfw14+kM5oVcAPoiEAt
+Gkls5/EnWJD3Pp5jlDdDArbLaGy6KoGknkc5nAiPWWR76WHQlwAseO8KWQSpzQ/Jcyho3P/UA7P
GBbGF2AisINCRgg6EJYgZtytZM/eqB2nwh/JZlB4DXjgaZYRqTan2/QlL2vuuvUpstgRWlimWnc5
aKtPQ3bt9FTVM3WKFWLTB1vii7QTUrWN9k0p+npTEzxjAfPshaEK3jVxyWgXHHdQMlmXgqme1Gkm
Kgq5/qAU7lOe+a9ZSRxzkwdgxxY86qNOiOtdpLBUsNRt4lXFZwzQghvJPMEQr8F3WraGB0XDKQMi
pBoefEUMAbs/72dmYMcB04lcKwhBT6oa9Ot9CM2FYbg3420TVor6nNxX8zQIuWp2Aa3Ewe7A5JEq
safuPUiL/MggEjGGseMCbdpohReVCGckbiPh3ot9+uVHZHVeJSui2TRcnL/yABOp0quN3ccjgATX
GqmLazOKFWkd6+y7/dVzt4czYfVo93I56L5eKOaUst3HSeuu1bMlz7vskDdnHxLmFJaDo2VpzvKo
dS4oSVOsKopYC5M+vohoXr5fnkWk9Rd2VTSJ30PX3oWSGX8U+bs9AlyrjqGVJpMbGO7Wamqd0CSR
eGlJlaaTwJtV+P+i0Om/0n3EztYCqI7sJ4S1IoAcoUHcmboM57W+CADRFc+0P1/tsfBpEFAvAgVv
91pOxS5bvK0vLstcjsDSmY6le3omT/UcrwLDN2nnLIX+T7pbY2Cv4L93eZZJm6l6SC9BkoyF1SQe
mHLhr2sSt3DWYFQJh3vKrpImNReJpNM0W4R4G8VoJfvPz4njq4rlGjqW7VSIPOTg5cR+d2fNtGwh
sfT4mI8Qb4UlIbT9jhvw+Ac4nEcNPCTLNCzhjlOPXgVd+VyLv7dS8UioLjHDt/+b7ysnfLk1F61U
C6VKEy0ex5VTHpJVk7O9I1uznp4CxRYcKdhzzlRYtvUcI+pWwLndMSobll1GQK05oZsLjqh4Bhjf
EFfKryV7J4oRAe1DZI++EC+T89kPx2xHRM7neA7xOHgF/QZRVbomwrX1yZ9DyT7JQcE0r7s8KAkv
vAqgUaxgbK1XmlSafGWhuQIRYcNzjyceXgDGfQ5XUziehf6+HV+piXfPgXMHees8hkRu/7uhax7R
XBlzU8s2Ve4irB8D0lX2aCNqE6h+/Krgg78Igk5QGLncNcj8EUMDo15b14IwDsE+mWyPdpi9HqRm
tzuDEVZ5e5006OfjW4Ibdrjh63Y4T4On6+DjCfPIEj8cqVGaW7jIxiR0edbdEmA0ogDOdJLP7dJq
lG3GrYXEYNqbJGG2tAazpg04iKyPNVUYkzs2RWPlNShMj2qgobqilRGNTRrh/efd5a5WKs3WHRy4
rhUq8+JpHPT05JGGPU6yVCqMZFbacnOLhUVV77ouswQcoThI8dMbfqSazKehG0LfkjFxpvGytQvn
9ccwD3HPlKTquX07jI2DxcszJedN9eRV7lLoQMmiM7SU0juLi6NwlMDt6a22hWG9THg14A/EywCF
qyjaFu72G/oHJfw2rRAGG2cw2/MR79kThdSNi1iVJdcrKBMMsZdaezsxyjQf3U0JoterdLUjXbaH
JF7RYCs3+4YeuzXfRUypl71wXkB4CasELUoObDmNky1eEWEDbbbcNg7tf92blfh3044aCLf7h2fc
6SZZtqUXcZl1eIGZPWo84O5si5zzuI39mz65lLQwUgS5dj07Wi2A1KhSIA2okwklbOIPf8zAZHu9
6r1NTsp0wsd/6iHw5FfO0L+NTx/23f6pjYn/elPXldNdHus1rxE0gLub4wvFDotZjsf3C3fUB4tG
9uJ/wNQM2l7XSKBh2TueBIRB4oSyVYx4M0SYyKyMhxJuba/hTrfsqmF2eEkHkJ7yuVq9ViyVzdYO
1W05PGCdZ1k2G0MoZNreEjj5BTmTA9qTpjnIbLstWpztK+GH9dVhJVydNrnCF4WFt0nt9JLAMsbw
/xlAorlOHweF6SKg3oh5lmg5Olk/iu+AZmMt/mM6NXSWWR8BUk9sIfDfYH+NcAwce90yKxIK3srd
7+mTlqasyr31/7OxwHMY/6lPr5IZBd992T5omUMTn/Ekwj+XzoPTAGZ5Xwa0BTOwiVnvOSyBDtDq
gJwzdCvXrxY7yJXnQkTohZTBQUSxrScyy9uG4s7/Vnc+Re2N4So2Qu5FQ1wi7Bka7PTwvvaYJT7k
VxoKLMfapZxSrWuboRX7WVFY5f6RldzE9BGRn/MMjcVOBDyQgNrC4mIXhz+1eBRQCHF/Lwitkhh0
ILHhuPFk22VKdpHlvEglh2D3RE+bP6wh16siR2ayebZHEjSLiDse4Vutj6qQKsPGnANy+L6saGnF
ftkBO3mv1KAhxYPkeyuP0nfUpl3jWu31ulLA60bz76brqfseTPusVk83hUVIhaWa2itmvsEhIt8/
prFDtCvBMVcO1F1BuMkxbYryjluVTFK9bHNrwLTbgK4f+COtPNUwE2q8aHchgbHqysXnjHJYp0JR
FXEZaiEDJz/jAlIPdkVbSHJDUbHbleXERm8UpynT7Ox+l6tAb/WBk4O02UZ5sCd69lm1jeLb7Utt
GgMIicvekvw4iIJXquJy1B8ZW2xqhy4PCxfAsFzqVSLbHGrhLcKB2AYSpqOztVgqd/oMq+scGtkq
dNfAx66aZSB+BIftQJen6t2CjL0oA0BwjHR4ZHPJY4hamcTyYFI7LNjan5HYklNd+LHZENoR32LY
obCHRyTNhhiSjeOvNJtgIjLSNC2iHWvHUU6FWmOOGZ0WW++8tuEsKIbM7MMoClSgXf8D2Gk/BfKE
cgRbScQRu2ZMOxnaSKeo4KghKMVEd9O2H3tUkpZ/9bJTBm0IRzlBrb5Msq6xBCwSeNK+C93hMosb
WeR45hodtvJHg/I08lemU5oQi/HsexYebvQ1otDZwMfj9ysrg56K21lztDhujnLFfWJyk+OCImGz
FvP8q4jFlwG/MAKMrxX+ZArmP1msJNdjqj/hdDe0kJ0jbA3srUGwBghM8TaYOsfW5bz0z4cnyfpc
QkWDE4KhWA7fesxysV9HSNUh8ebc7rja3r52lScuUh7BkI7LPrMhMDZkhcEMNrob+xSt/i/J0VcF
EMer44o48RE+VAWM0LlperELtP1fw3wTdHDiLQLtlMlvgXFOtkkUXyqZjtJaQpHdxS/ithBxl8HY
da/BMpCvh3Qob9KW6MVD2/CsA1w5TlmXrdAQizDaExChm0x6lSggdZe0ZTDZfb+L7aLIQcS5WMic
N1npd3t+KBRuQQKHKoiORv3vNoK4q9KoGvCXeK3imQJ0+ra0PpyR7T7Z5IORe9f2hlrEzenhhgNe
AP1y5e/3CawTny3eSDOF2VbOZuAVGOWKYOk83HzTqATQOxUFm0Fk8wLgSntRtYtG0YEg8yCCGrAl
mlNhWc52PFGyA1OMGLdU8bM/kThcTMbJ4kplOwTGe7suC4uLi85os3XRCG62diDPkBAXPKnsnV8m
8Z1WER1CzBlaBWI1S6ER400qhbAD3iWIxKqgjZ+JHU7/ZISrNzUk2wlp1piir0bWsRVuSN3tQA+b
RDZ/l7YjrZsFtn0h8zRpwGen5RlutRpgu2tD+Y6enfiGmjTZOHp61DOfnQFZnqMVo3jxCuo5pEWR
yRPMjUYVD2gjEYWWv2NduvvVplV6NYg2RJJ2IvUUYQkR1bzVEKHCDo0j3SdVPjP9K00XI4o97OVC
VNa9sftcCWDsKZJqvbxYfuQOR2/RsGkDSDFZfAVnKxwsUPpohvUGygIr4H7vR8Ru5DMuPLoxmvfZ
MBBUfkStULKX7zqfuFpdVaZ60w8L9Z46l45sASu9OgNo6dqV90e5K0zBRTr7X4y6QYkSyyL8LPbM
om57pMg80rfNKHquku2mnBTUn6m80cGdqp//jJM/VQ0uFolr6EYA3CXu3Uq2siRbAhpTJPs0kUTZ
QlT/u0twP9KIB5enpzHO8JEatXDAy4KfaAW80X8BHVNt+ZLZSAA3XrKpiSnowKsrU0fWiHxexCxR
5PjVi3fHaSNhDOtQX4z/qbi+LJ+50gjDTUUlP2Nvi3Z9OhaBfTGOCs5i/XgWATlsuzbymectfz9A
87CO2F/DWNhPUhGqsKVp9jLkIWpszN7afeCU26rmPnpAsSLQrmEUVdOdtShZSbEBT5Jl/Npo1AAU
XTXfixnfgXUwL1Y75VWI3zTx3mUedCsQ9yG26uxDabVH/RrLZYVwOuUnJd9Ti7WkmmWwpy1u1G4O
7KxjjpwuyfpJe7O/x0sAg76Kp+MO5AmP84N1KNoCYyFaMe4axRqJ3Dp8vomePqPBVOfG3iImj8ws
i8Jl4MURJHsgT3urpmK7Wr3bm6X/ayF9Dtc5T7/hVC+BtDh8tMquYToteG4Q8gOUbA2UPToPRb5n
t1ZMTHSMBMPfysJEnbRcJuY1JSxvSZVWakG2BsxBfqV/D3HP87E5F0r35LRiHGOjxvPHACgG4jIy
LE7NYgTbBeCXRWqkMVKVGDafoH3Ikte8W7KWEqteqTwcj3L/4y3MotMnYQ2BReX03J8rH1xmLSfK
vpXQNtHST1KvlTJZK4rvI/ZgD+Fn0afZvkIkbmQiBFZBD+8EY5u/QoMGmCH/VfoGlrgDxgAd/6Ha
jZDeNVk+DKjI2i+mTeBqYcJ4H7WR9Vtmmhu5Xq6rcYf/8H6wh3CvBziSWh97JRRukmUWytiz0j45
u7QNypeh85/BdBzUxm38vwbjt4cEsXJlY/V7Fuwntr/0zD5F3iM6ZseZjdIQpA9Htt3gC0NAARE1
7qHo9VsfqkCrEOU8DJQ8sc6VMx0hwtnjS1ku9tuCIAX4ZaXPpjBEWpVg0oEFL7/quC9BRHf8Fgkg
e4bxqmXkXY12eYhsRPI9y70KR8Bj03zOvwDr5aQ8Dnr965LYJGJ5ZqerpQdiEsj4EXLq8fcmxkZ5
o3dnnVIJPktVpqAiC6K5k7THSkfuLqeMd4hNoVLgQQb5gDd/cp6Iz7GnZ6AZ105hR37dRRUrTfhl
tIUW1Q8DYhfMSWWKSp6NUa9DismovgUBlniHrQhHAQGSZNg/NjlUHBg7PDnyYpzkA65rVYVGqdxS
65YVjTvK7o6+uwSphaVM6Fxeck0XQIJ+9d+TNHe5kVu5ui6Asym2vvdaU+wLG8t3OLfJGfLZnwBz
74uIQZIwXwuQNYRBWkOi1GLF7n2drFzK7dKMZO55UN1dIq7cusqvUIlW62phA0375kIcW1hydhyw
WIWHR298HJBLCBVc6YJzOm+UeRhnfGn37Jsoj81b3z+DMzEUnn4TgZJWPIpzORm/z08FBs5BD3zt
lt1bcrYVgV9zAhnGBUmX9SomaezoAw2Xs0AuJBDUfPL1sQ/jqY46WGmFsjFAwf6cOrk2qF9tMwXo
Cd5n50iBmWmOem+ItBEimmIpfVPi/U76+Rwmn55wuCe6PhIoeDcOeU1d6VVeLQ6eddlFmFaPPkQf
3BCqJJK8tJzmOVvADaSBwl8ek9wgDndZpbfFLCFYxSOm0GLn7lrEV6xe4tro3AVgQNYRGODfIzyP
Tj6JjFCgNnYlft3v2YLx+ggqaS7mdD+QocLjx0inDmAVDjhqClRHoQD067OdvQTW0ur3GjX1gHzW
basr2LXzxT4ad7QO971jKPoJKoGpx178M8N6sBTNEw20eQ8RyxGT/5QDYX/enRA+B3Vuvm/LiXZv
DlnucP64cLSn9GQudgT2uL3lDiRt+yQsnVOj7JnINxlUDBSxwzR1wK7W0D7aoDjY5vHLAdaEMvM4
czwOcQmLUr2X1AzzuaiSgE2GUbFIfWhmV0AfcgUUSMoSonuNBKx6T7G9BK/lTelNILpl2mtTE3PR
nKjl7Yb6O9VSLHRhywlbP1DRvaZoBUlxsVoXiwM/UBuetiQp39ojOk/+XhNMXoyBIbxDRnlG4zUT
tmzQZPthKOFebezvxeY7Vwr4H9nb8XDfXq1c8fa6usn3O2ki1tL++UKBDF1T7tK1+7rFIrJ1YROL
s9tE8NW98R+6dWMhsqB7iClCvz4d3fAw643rr1xFuwuvvSjQTbhvHrULrnIcagZHrxDdlS7X+w2a
1RgJDojns+J9mkLce0S0AJsD1kqktPXV7Tch00LLZWWxuTz9uH8lsE38qj54rJUtDkUAHuPiaXZo
p3CuHceId3nP+2U/kIUbGG2bcfQqRB6erHzApNygHOX4utvUkcBiWiAkKOHrvRK8p7VXN4Vc/Xja
9xfRR41eMu9F5wm9zVBVRdUTHBlnliJLpyAiFcuiOT0Bu7UMJLZ2xgDthG0lGiHFhBVMcmYhtesI
YcARQFPnnKPCCY1yclno/R/xTwAATJvZgFcj3TCbhQcggyX6DXjOmCcAuCIiNYRzBIWnGtGVPZDV
gfA/S899KXgG8+nWlIT3OgkFSVSd/MmAAyfs2LyOrEuWXKgj4CK3LySd2fr/N2+oJzuJRIuHXnq9
5ujmOut2sWsjFxGUKtEQBAtvY1P1QgzfcK7Ue8mmR74aNEoEf1L6QhocCViyAx3UBIFJM6ZfxBb3
HpiZZW703HQ+iqqK2RpLoURG/QgYYl+mHlykZpV7O6E+KAkYUzuYNtNxqJEKI9IBGpiHkB6RaHfT
quZpN47QsXJkKDJe+fiLRn+im3e3ecW+EQQt4A7/O7xWhWg4abRHnhRkMFEEKQjf+QgVFplktXxL
uonE5OI5M1+yc375jUyj53tFdsc5AmWwzIJj4w8N6JmWdjiF0kZDqo6o/F3vQ14tHBHVJn2ARigF
vBwuEjHfP6l6UkZ4bf45PP6bijgPCAPl4xbegjgAmd1VTLlN94OeqJiZ7l0XiXGWAqYu62s6dSUE
hxQqKDlbAwN3MLnk/JmsBVr+5mJL4a3ti8uiLjxmyacBY1cuJ+DOyQ9E7mx1c+IxJTEHBHCbDSyA
EbPmV/30J/gepec+kanSlfiluf0nOI7sDbuSDDrfFJnb+pPyFJaT1zkfgI0cwqUvJT0ovGZ0SZHA
XwE5TB13TLHZqq9eu8RFbAGCOAQWuAzRpvuSq1soFkg8RkjFoW/FOEXQd1kVyJUA7a2hECzJtBkf
ImC6IBm4EP7VMYRa6I4pBXA2rx8PSS8lirTASoLXShd1KO84lK2crKAADUpKqCQmFTP/P6r6KTV1
2XX69FpySKXnNWzq+Chwc/hVxGDcoI+sc9DtjF20VHiQUOxpYFZVNnPoQP/B0iyaQ7urK7fDTLmE
pZ/lKDeK346zN+GlQl0xtX31WP0LBt2Je2+Ac5963kpS4THOUcjNUqsLg1NFlEZhbRqLODlSty/+
jCZnazuGbZknjrgQCmZKkHuRPVtF7O61M6EEK1HRWFEC9DU2FK5bcwOsccL/t9mAW++FXkcu/AWi
/bA+9qMyBkSjgvZFmvEWd1j5e+7+iW2f6kcRpBdcLpxCYIdgDw5DEzwf7f1SZVimGvFHAAvKlnYn
rQ/+c7yzieZxP8Jh1xKFd6H69gAloBtJ2bvaIEzx8uoFXL1CRZ0uVPFlkrqQUhwYDKb/dbE6Ggwy
PBhT+yTRFvAVD3KCh91G9P+WEjkfN85HTVjwA3GHh0lplI0PkC/nd+EAQ2380u8sfpo40gI68OGx
PieIsZvOqHXVmFAlj3gQWGsPrnEHLYLmj/BlGEnuKmaTYZq3fluGL8dOvHHHrmx5FVSOoCHmc4rE
Z6UFg/81yvGyrc3zwcbfIGwARXlw4XKqlRKxn/hqeYMUvUyJiAICa9uNSJHw08YzdqfAHy36z3Ns
2nFBbqjGYqnDkw9/vKHg9tfdypdt6QUJ1nTav0/hfAK4XihBgani2EeJjgRUti/Us/PzhriEK9dF
ljdMMTma4XIrqSuMj+w14nqP2YfBrdizkTm74iUA2l4aC+G6I6e3S1jlMlo+R5V/KWQ0WEQ22Uj7
kiaBEvXcPTWjKjWr5rW08rCp+s6Yz1GpJTg8W9j1gIlR6egXDHu4/D+9PSdpOFXMD1Uawoz7x76P
lfaN47wX3tlwD1HGjb81e9/ek4Dfql1UfTqnuDjtECZxhqpOnF+oVWGHhTg0bfnnqUDcf2gFK0qf
NzlmJZKI1XBHAA9scmnXAJZvJMfGAQW0youjOrSYhx2YFMIETqrdNU4rDulksJpG0z8Vpi1SwmaX
fM7z7DDqgoP19ZLIGdksOVZZxjE1f/GbYjxghPlZCiShB0AcUFM8vvNs58vt99KWIQ/i9iKwFmaN
WSNdys78X4NlKsxzh1R4/FYOlkwWfeLFIUBzR/Wk/1Z1DlTPK1vmGhl7QDtRRJi9hdI+YA5AGanB
CuNehHDAj7H3cR+nYQXcHsKOPztZJTRqmK4yFzhSI4VVqTPvg1J2wfDdgviOjaHJOKp7XLGIa8Xm
o8VPEndu/KjXHV239bbM5FIPE9G4Ygc+dYjUEbVn+CMWDBLqU3HQTbc0dcELirRHeVUZl7y1Pv8P
4zl0t1DKbhmA50o6WEw96Xfl3B0H1K48FnvORECjRJF/9MH+ATgRdR03PvWoKvpYQgnhXk/vIltS
IihqP5z3/PEEfKezfzuVFEXIyFwRoxUKgVaL/+OTZqDxqEpSKuz03LPhAg3c1Q/OHJ74rnZBxoGP
sM05mLbHlqProx6fG14ITFjxCjJfmvlI+yFQhi0FvEPFJFZyFWrFgYuaA7TLXDAqFQLv724sjSU6
6+9FpNmfwVb6RrCddb00vs5zWAJEBlcei/c08QO3vwO8lwcDcGP7aV9KD0VeKysFkiVJEwZ8AFGx
ZHGN8Bo566LwmUFgYFbkXpuBfYGcZqh2CjM0eUbOPGZ0oVDXfWgaIc7rwRkIfb95/IZCCZGqIWXf
igA4qZPFHT2/R8gLL+00OpyDv52C41vnQ9O+D6QYnnls5GWILtbdFUbI2qFlQuDsE1SMmJTXWhMY
da7b0kA9T4bVhq8ojoyC8LuyRCxqwO3wshJ4i6LSH5Iv8Pa2bwMQPIk1GoI8NQlo+uU5cKwzFBU7
3CDiSGzhBYgFyqQP/apnMRmVzdp0QL7ipvx0Pc9SQKf4P0BtMPEQ114w8vgLwK0UeqLuqYty2xIc
dMULmIj6WJwHE8ixBqfd00AjscUzfiaM3D+NIaK0q23agIDMFsg/R+5jSZQnccyZd4+mOPyaB3ju
e/vsupaaoEKFG6eZFXjvnTnJiDnB0c82y7yG+J5+3On0WYkEsVrnpbgy/USRqv6tiH1H03Ul56s+
0dXHh2J23eZiA2OIbBuhns2n8u9HZNCYkxNoH9/0GrteyGxf1NhibUHQFJBgtZDsCY/wEyI8drRu
ubqnMsI7upj9q5gKJY7welvZiLLj/7SML+Ajiu8jAd91El0aoay6wvoNBmVa8fMdKCzCiY7yzFoH
3878NrbvocLyc757MFLQV9BQmJDIw6cmnUwWLeP4SJ9dH7SM/jZmhfWFuE7uLEm2nJ+kLYMPvk71
J1I1wNQIu92y75dID8WryZv286oD+wsLlIJRDxIePYvh27cQSLXuyblRv0DKtV8zpT0rubnsuJLQ
8DfvOkzGGWauGRMxLVIRZPWke5tXpWgg3tzTeWscYEcWutjDFWl+E39UfcWU0vZ8XJh7MxJKrqJx
d5v7/PlcM7/QqEUYs7WbY0Z/eial+RANdvVRAsE5hxCSfK6+Xm34Q2BzLUdXU94wRpWUXzg4pc+E
kM1vdRmeY31JQQRiAlk8pQPYBkDvyysOT7Kx/ob6fJ0O29kEazJ8JLlaEnY9SJy49vaTDlVBcaMy
qB1nKDY/R6+PYHoFYFEOGhIdfYkLe63IeOAkqo1OasFsFXlBp8OoUUqMILPCWzFnmk64H34368uu
bSGwH4o6ZdTGciKsF5Y7VMUlVk8+SPgmowrKbx9z8LoQxMVeLnWexOrWEO2J3ylZ9mkDqVxH/lZ8
DH+Ceq1yyXc30S/JPdkVgg+qsgkrjkZVTr1uW8vkhO/67vDezDkUChv7iLg4uiWxwCBlOhg8qWpT
xlS8aTK9sxOh5rm1j/mx9wsjSKF8ry+/kIGz1HHx742I6Egz/IcuFfP4W/K0aECfku5AEKO/oYj+
TVOEBiecw0pmDYLc6NRFMXZpcwNNuufHVpcaBf/SVZbuBDLIQ8+fvwOviKDws/zQ9t19ApUqH5Yn
8VqdpH1yVX6qT+M9kW5S9R+VfEE+16DchfdUEmk2VHuJuq+i7OqvZHQlDVZDFt2cwhb9tMeGxi+r
SZz9NOR+Y5cVSjiK0XJjidkzRitR4hvkx20fdeBhuD0UzJo7KkkOgDPl0xNuPYuPjMOaL9YLz9x/
nwhPBcHU79xZpyMwEpiPF/I0Kz6KQauQoQu8yqLjKY7xzFLEWZ29SPMpkNoG3HHzGPMVMLTyB2Pz
BgPbYTxC5C+vYPnOoAO+bQAzLjRwl6whpvceoA5oCKvSF4j4PXs3dY/OSsT0x17Z7E9hoRkrE6HZ
EdluZDeF0MaeI4Qu2a1YZFaLl/E6cDRpUPKxlGjR8YcAsq+DFCv2/t9g0a+mSHiGLinOpvMx7jLz
IgNe7RjvVGWmEWWflkOeEYsLYrtMTpmNaq98NWtA7cjwD8eGtHiCBkV0GPiRGQ/hFhwrpku8NAWg
+71qMlMcQd5J8okNyeSRqfhPnEltztUZlyf1rI0H1q1hYWMXzZYUpmfF6U6MMGFrhgI7uHt90Jv1
95dbVnErvsdXV+ivEkRfJPrUtH+SygeUfvrrrfeGSM09tfB1cq1QWJXpfAa/6bZo8uCl5do4Pc8B
Vcrh5QA7e3oWNafrWsYsGwI+WDdJCsqMfZId/+BXgvEkb0xDbQOgDbk/DG1VdAHMpK07s09TeqKz
4uDJNL4SXQHyEdKEgWVoo3AwOfxUpLJGiJYvtJAis0w30DccW3nappHWn6LRd2xXMYaY/99sBsXt
gEDzgYFDaWCN4s+Itmdl5gVnVDNWkIErc0GlYz1XJXl07E4zW7JyHT96tz4tdnyujbsUByB+1UBK
kr8zj7JOaAP7kI42gPFjzNPgl86NbAijc89FKpLUxO2j73wSdgCmgfYymMVLB4wJxBEOwcdFnlMB
nNly4znSpgSp5KEnXgpQJGy2KSlad4ySr9GKexpRoXPMtRXqhglmM64Gl2hWnGDrwNkscmJMngcc
YGL2aiTJr5b9XFIRBbCUyGBV0cpqcXSbbcPF0LGyBcN8CMwbtzz07BTjXh9Tq2pC1Z657nqQl2pQ
Ja1p9zuLruM6nB/w/VEOw9m8ZZXqEoAy7WQCT00raqxefpD/sWXxAHwW4ehJB9NHjL3a4bglyYt+
LNwrpWoxfXnHpEH1YISOTwfRzMPOLWfVdOAk4OFVoznyY24PHBTNOOOD+L/tn8bqQS4hz903nvGU
ctdIbqCl/aP1MXn8FPH+gOdfWXfbLS5xcFSeFNlAg4yH2VvFoGJjRx9CpJzLSxVqhQiXdFV0fYvb
FGmetcAcwFLdXKnyHL1UPL5+e46DubDyGEPFEQhxWRj04SFczNeiHkXdld+hOpNqZhgwdfBuADCh
ZdKWYbpavGoLdF7pf/P2J4ExM+03wRERePqIYg9zWphhLWhIw4mS3lbFg3zdb4NLY1PD2dw06J8u
Qr/RvB7UOndNUBUb7J47KwYcL+EFJnZcfjR3UkuTOLGuVuFQCAayNFNBlmr8mfu+gEuOmYEWiY9x
MAeTarOCvbfnyNqdcc3lanHWmwxUyV5Asi2m2/8EMXEptdfks4KLwqUJSnVztU8dlRxRav1c1Zms
uwLVLNnmDgELHO3jduilErbVLrBSRVs4fVM2nS4g2jh+Ll5koIxMsKVoHZlJA7Sg0b0HFCX8VvjO
M+oOBNWhRm9nNU1gODN/FGmCvizGnKg+4Pc3Na/JfWfUcYMWnq2g4mEgMP52V8K0/as0iHQzZrtY
WydH2VeGU6nSoQkyQ5nyuBSoRFLsuRgWqKzfLVtuoClCQY8rv9Hw9aXIcI+KSysxFdBqSoXVdexF
zbPapmaG8Aw2OA4kMg/XYkAk0jrA+9vUIhNS4kZZRs2lS9wa6AEjBBSOHD0cU8RJUM8WrHZT1wE9
iA3bcb8hR2qK0bYeMQO6xNG62w4hQsgQfsE+eAmoQE3uWDPtFaS0gOzKvxedh5FUCWwwUHlnEsLp
/LXd5hLLFHL2sY1h3iPtG9Q8FYnPmO9EOHhmIh2QDA89Xt8pT+jJ+g7H9QYYMYf/wTQEanOA4NI1
eTWRkkXDOoPEB72iIBITuqFpGtiC5W+J613kYLHHN7mySLnnJfC3US8sKaHSsQK7RxRlCIaycgkQ
Nr5ZlAvwtNslVGUfzJIJUT1tSrIKCvd+6o6oWeEj/6dJ/6pR36HPsdXNr9NM0O+pmQC3G8e0ediO
UQ2eB9ssSQbTVVtcH7rw+MAZqMfFEh7xHmcybSdeROibpNbRHoMyAJoBwOFZILXX/MfProTbp585
w1OE8uP++42vvUU3DL+P442rDoBokdvmJIEVH4bQ5bFKW2zvNGCIst4UKU4SEqdqnKybjFFgVvBZ
ktHa9LPoBUx1ENlr5MePxWX9oAxCK89YUXC7etKCjWGH8TTKWlnbKmSIfY8wLZGYMpsYT7cydgD5
Q7UipYLe56f7Krwbv+LazaZ+iqRK4Qu7molGEOz8F4ufcDcA42rP+dJxvDGiNWKw1f0Djfcwr3pv
0QFHD3HgFtQurm1+jHcUZwW1dXdFur6jj9m40vIJD5GxYASLt86WMQLgqpYolWYLgaEb3YojIfn7
V3izzvYv1V2cbsgo4X1Iv5vk5DzaG7qFTKuY3G93alibgh8gV9xIIyCFhZxRSnVgz2+FjUBpKopb
INNr6qE5x6J5nyJNIh65vfnUKQMvNC+DdXQ3pGSGI1Ij4QDRO9lvQshpQ3bdjuYmgmJZOlMN96AO
4gPDCCOe2d04B4NIFUl1DeGAT/M5cyqLreN+uVIhbIpawAfouEtnTXr5okMj7zHH03s/yxAUiH5J
tzj7hwDB6h96i9SDmMqK79ouBAlFll0mETXNL0QRatDngXWSOKId2r+Y3Zb5Et7A1MoHKDh6IRWw
dtkhmboa13/DBI25TDnj3QCV09+8Wjwvx9or27Mrxlfq0kY/Ke7kULQqqYk8HisWXwJ2HF9N12hs
/RtOp1LmPa6DJ0UcmTTcsuJYfXnSfCavbgN/mIaPQ/ICb+WAHFMSJMa+ZVfljj6esf8UnwnKj40o
lZg/r1PsLpNRm0By0nEnRepqsq/TqOlfXPWsLOtgiWeHEPLim7t4rFA2mRL59LOVaEc8KbFETwKR
ZQiz12pHO+0ClkS9aTLaVOgNBjJtk6b7XvQC6qtK9GRewtYD1HmFjEOcHjx3EKLAQsqGaOeJAMnW
Dv3gkviXNwe3oZcOo5Hmb3FEDz8+wvITbh3QIlqcXLh/QcJA57F7RvvwXl/JSIAsf4Peqb/cLpr/
O5TCu0Yul0KQl+VW+dnEMgl8AcxgKtGLmvT5XJKQKMjNoWN5exuqILIThoE2ZK+VPqVCaLoRDDKj
LCWi+3sFVSXEg4wxhNnLJkuYOPMi489dyIGX4WQ3XS6mvlCDIheXBskN2sNrvUwD4zNwnx/yoIx5
SchsnUkZGL4aGhLqe5A9TQf9E7CWiED/BwkZTRcMekgSY4RTPmJ0Hr0q9/upksstwEMmdW9qzGtC
K43kHcF3QUzYGKu4BnH8RlDZt4gQcLfvUJzCue/nSYwRwvlj+rnqqS2DnnnYNIBev5i1Y2+8/GKV
ah0vTqV3dlxkhYRTEpJ8QbKnImM9Q8Faw17NVZkUweGuGwvw05JYon1AeEbpKqFdw3xJbs1D1Afj
1w34tuX/0LapJzxa//zVkBKLNvBBLdE862r4RO5ny5ADJJio1e/RsOnFTBsN4lsXGEnD/UIoEkfB
BAGsWnrh2+TqpmkbmRhdeEg+FVIGJMnc0j9oTS2zgoE9tF7/Qxs/Ghd936KvsXvgRlfiYWMsEjS2
47/F2FPsiu1WB9pq//nbU5LWjmWclgjlUZBVcpIsS0OCXEqCp0H3GgKYRxEA58Qq5eNdS2Tz2Itx
rWXF7KO5fCa8IfALCXqT8un0fpM5peNp4Fh2zv6ve0ZUfxLJna+0/RlKOQYO4SGR+2thoIN01slw
GJw0jXfQc3aZnM+pYLQxa+xKiGMdnwXbwQlsQ7GnBJVda2ZezwYRudEWYv/KEcSO0Au8yX6Xj3HR
TJQtek8tHIj+8/A2GJyh5Qh4CfAAPCsjhNP3B4hpo+8Gn2i0NqnVbirIJ8MsxnjcyJ0oxSkC4/0G
kVBmMyxZ3IUe1C3k9YHg+tRRmM+0xy+1A64I79Bsct8EifbX9FHCdPUFkWkbPcpSYtfXBvsE6UAQ
+yEPFGuOwjPzhDv/x100syAQMkwD2/ZrPIfVxWNMiIUC9MFdvx82XDH9IcAP4Ml5zTaQwFJal22g
Lr8Jqr167LALPuJ4TLCgih1Jn8RYCL6Xae7IAFy2dhvUkhrcxbkM6rzExuAYeUECZuqqrVLiRN1r
GXDuNBw8XKPQI71AY4hnuIArkkdmEd35qucHctZaM1gIv/I06yARpYRhC/53yoxT0LogJyHNPqK8
fEULufEfHa13+2ZfTs8xuL7Ph2LvYg7wWZPzvcI8U+R7D99Hps/spf0XTrg2RB2IwSc84bze2U68
KrCVG81QBjVlg81YvlPYYr/iON7pE2WloKFBHeEquXPrzgLCcHDTxblRFuj9290GuGiP5HSK+Xsu
jzaF6snZykt0vcgnVSabra3ZfQCjs/Dr1zdqnUQ7JtW97gLZC02reRXlPNF00PznIG0iL/GEr1St
xNTlE0I1KFGNbaXqved/6Bj7zEjGErcDyV94QdDtNqtQm1hoq9O/ga3NqrAzlW+mnrZ6HJvRtkAk
HrgWAn5ZbeZPBseb/U3RInv2y3Mk0Zf0g6dNgKEDgzTVz6SMavKHUfXkRTq8yz/Mv+pVmStuH4cx
a1JQcXL1swmpKXIHcm+4Cv++hwFJxYuy8WT340XKNyxU0FSfCmDcGcdq7Wj/L42xmE5DaPDoIn+v
yLtBhGMjtR+o5tCrGN90EkLqytXwlGbOs+RGsxeFeAz1NKMXHF3lIXN2BQSVmFesFf9JCUZz+bLB
XS3GbdPsY2OPtzw1Oj6DkMqEfMAHcPXs1/R3+e89mxQ8xOvrgmepTHzm+i1HHlrTx13ON2rfY+qa
OM97gpvBq03ms9YEJ+eUtjMK1ES+eczchendLIYoQfHLfV3p1VpQ4HD06mRr8PJHLLgFHYh2BwVC
uwjuAzc1lRs7lbdCcb+aVvUG+sdOPSXIuBcpiruy4T3+BPl3EXOZQUpM/3BTMTTeCL5MLNmRuvKC
r0OdcfXCpGYZEyS2e+7Uj1Q2w1hmsBI7TnPf+Jvz++qtB1ASvF6AgscNZFHXnlIUHXiI4Y5kUL4e
4nQYCiHfelafxmZxw6p2kvH9GYHXyGmeWDMBURz8u+U9+b+09QcKfF30uuHmyYBvWIzUGAEJzwvN
hVpYv+jK/fbdpTdQWbvZmLeeXL9/XyxVANePu27tRCUkVUOkReqU2VMvnogL0fTzslBlOH9JIgGy
J3KJBhSrTpFDIfckbbf4QXM3obyr4zGp3E26qYyoja9I7ggmqt9MczwdnKazBueE5VIy6YFzYE33
1eUDI4NG6eOo2Ef3m/Bg7cV1kT38IVrXPZB0I8aujHHxpeBH2f5JwUL/aF5vcCFROcz9PINtdoIz
KSMaz0RILYJraGJQ5JwOFxEsOd3OBDOhAigp/D5mLYenVn8s94ltV6+G8jlsWyyKvrr+HblJ2yS9
gqlRE487kOJLyMKxmopNGuGYUPdAXlCnxKN3KYsVrfhfW27aqHKGbAxS6ZqdCXvjI74IybqfGxvv
Z92QRzeuMCtLUeAHMhm5dol5ryo50f1Nga4vezukG7DczF9Udc2cYhIE0bWB/ZL3c7MqyJ4PZaX0
Et551mp2LN2fcMaVksitTrV912tq0u8AgAEFgU4nBW0BsgKdzEPo0j9OeQ9/1Y6nMG5+Y9UWj78E
Zd3jjBLDTZISmlTsSwWJ+CHoeB9zgMJCZGYmyBeRDjLTBco7h4gMH3tq01l39wcRj3ylstqTBMFU
jHWFVsx/L1LomKSAbeFN+hPiP+JfhbqUbVKVjP+oUW/KzG688ZnzM3ENMk2iAKYsU1q3/1/wIgqX
uckqSRTfX4hekXjJhmKMZEK7L96uXWVENuiX374ifDrFy5wVFo6vh1Hi/RKb5OR8MLjs340fainO
N1vlLIqYROnSiihDQAm3nvM11k8o5NTb6gEToTtcYK6fFfNtGbDubE2Dda4P+ekVsJh/W8KYrLs/
hNbxkQQUxWOGyUUqHX/WydSloFV0UaWvAVd/qO/PG0IWriATJpxwDSZFohL0xdhm91AaiJeDFBDW
0vH9vImPwNviiQ/cbYiATM9r7ugqVax/x87yizE7C/HpVihWTUgKoz0ioQj48A9CQ2wZ2b/yXjDO
SxSbZQczsjUMRfPiV2zKbQNTlJV86qUuY7LC3a2yzAiya63EOxN87e6zXAimp6Ib+nL6S/J1Gks3
SL1hIw4ahBBxtSsaaPKrQNadJT5QERGy1y37SIxDjJyxuG07O+n/unmOWEMn4vBmABq9dxhj+DBf
gzLwPkNya8JU7ZNhAjkYvUqQ5r6PqgF18bphZJBwjE+tz3asCoIuK81y0LhUfEaThLfb/pQiN83c
x7LJ4dZiZzzJQKXn/1b+9hE8R+OlHx08uo1Fbr7kfG/ApJLuy3B0PJNE9e+Q+GC3AhXmby+VlLDr
vH/n4+/2wUOTCpU/8/0HM4WgHzko62vXrvCa6fuROCDN8ygfZwKEOkzcTCb3nxu1YK2f9rwZKT1R
AS4111x9SXcg9/5qCVSNeGdSfFOc8084Gyb9c8xlab6RVrSW/3+tW0w6tRVb56JxssWNMulr/gIP
NOCIUBmdDHVWU2soB4qLrKCbQQj7ZnyvTHLu5VKe4sOl4WzXDmjLFcgdBVwdj4vdjS0lbEsc650H
yEBRz24kAjytxOiflTnL/OH41MqCfHWJYYIcw5OrgVDUPyWGCh/EdHWz6/pb176YZTmGfmBJo8Gm
+D2va08mYrjzqOskHf2U/QlfSZECEefMjEOEZ5W66CWMPe+6mSGSpJc9p6x3osYCXOiqORS3FuXo
ZkOYohXND//tsb6dt9g69MwCJgiQWP+eB5yuC9zwbjDWuhI3bbgX9zj6c0HUnDx365OXi12GADPl
8gG4ZGtOa8QZRJYie3eZRoQJE9wKlbH/4VjHjrRBrtP0dRHAssHFdZQNI6L7azu5at0IQVCbFFzC
g3vokBDFsHiMycCsVUF8I99HfhlWQvC26r1bqNaZcjw2MkaFl8wCdlIChO4Ev5xXQkDKzS92s+ZG
iMvujCGs86u4Lf7UysEuO3fyDHXWcbMe5RfwwlncH+N1RgYCkwehO3qeHGg6hXNtu6T6jiKSX21Q
kESiTL3OmYk5jZxRB4oxwnDNzlRmi62RjxLKu3PNK+146y759nVOHGmAGyemG0w0FPikm1o8ciiy
5c0LuEdgPHMRvBIQ/FpnQ4naCZ1vH8vdnUpgHyaqPyJWZHbbTAw+J7HcR5GyYD6M2ck9jhG+Sdvp
WXxovvC725l84PVsnQoZfTxjQvz6HCD/+XpEVYy0dRC8kex04mUyITH3T9RRMJgjczTp+B4mrdsQ
MjwbHpJMZQfw4CP/OrmrBvBWqUaiAAAXlQz6HYObR6VdR/G7orcU4OnGpHO2y9nvaYi7B/AvCuFT
iXHmbRnMDz+COWlXLBD8kFvXxHngFvtUjqdsobqIf+0yS3yzp9Lskj+2gVqj/grJ+Di/Vf3rAWZr
ZY1LshmdgQirU9Vbj9ASsC+CfvtG3bGZzLQkufk/G0SpaVyaOavxIjsL4MgCaIAqnJUMwMaQQ9/R
FTKuZhCe8N31rvgHx6Fa+54uhrbIKz0lqboVc+zDohtONbBEV2ac9UHnhpjI+b0R3jfRVgzwzUUd
4QsPMyIzTanfEW12RP6/bJ126QK/wqBOq8pHv6OPunzHBmjkBt9mhV9Rm/jXR2QhLbILiLHtrMWf
CEHXwBH0/FWxaIdUAAerb9nJhoC4LFOvWAgMLwdXgwWrmDvdpDH1rCOj2AXbSrUlHfrZR1nipKqm
U6iSpRjvMgw7o/bqjPHKDzotJY8Xcl4bvkuVd9IjAKoq5Hb2eDc23EiA7CBXT47BKOxOQ0SM9GD4
C9EWUM7XrOetr/2huZ4i261/JFphEptoYBVvRZePAJU5t8gaajIp43SegdUy/oWaNfmTmXIegXqy
DdnupMJsa5VafY8SP22YMm/NduCxm9IGSkoufFcQuLXec3VX+7HG39dV5IpQEZzPTkbNuOcpQ/4x
GK1tS5/wnUaWM4bCmadAhXFJVJe7BKOOPFGpHY+JX5sZ+GXcJ38wO/g2dmnVOuTjPtqbVKh7s6P0
lSDUb/2UC4ywMzb95jRBt7CetPdKWrbtxa/oEPPk4uBUaXNiMdWMT+wsdd9n7bSQpqaPwCt5BYdr
bTURHIsr0A+cRhqnAvipbPdvcckU7vvSsL0MWUEapta9MBelgv665wV7wUTwEepPEiDUOdmEiHUm
CBQaC05qEBR5zGFjRh03SsnP+qDc8QWPBKFekHq5bsZ9uiq7qZxE0ZRIKKQS8ens0qTi3ILZ76p/
XLRWFRM2alFty3PRlL27aoGMBiAV5BON4hJPuiCnopA7Q8oM3zRgxodW+vG4S9GYva69fP+QuneM
z/yYzf5mqlA7jhg3R+Ac8u5jG6qsLEfYIhrJLLeK0/ISGLz/bnSinuljiCFXnApP48X6eDcFpFYQ
Xq68kHol9ueNS7eKYG/KyZaxm1q6j/2LTDVEIv9+ct57jQuy+I/ITsCXYLQNXhwU8JDK2EuGtJu5
J/DTbBdH61woHRZ1RkSWNfwHNXG8cz0+YAJ6TFkWLod54QBtQcNo2TQ+QVL9uMKmRNOuSrymxcAV
SfnwmYWOweZJYpphFDyFuAuzlai8LC6WQMbIF91FaaHDBg7RdmuNFsPfkto921YdIFbT9tP8SMeF
SQV6sDzBJKs/0ke0mw2wCT6mUcPK9o+daYhk2UHvrH35M0y4pS6F2azIDD6I2z+ZxQ+VGc9TGBSG
W1XH56BJ7vU67yaN36Oz2/JtM+hCABnDgmOqrvziDcyz2FDjh27Vo9+4Gn+pUtT5bz5L4liAW1Yj
eiKGQ9C4UiVF/77ztg71ijlPFzMavah5ManS1f2eQP1AsaeSNO/02hoFtsKca+rmDvfJFJV0KeYa
nAFi3R9WBenA1VoFblwd3vVA+IIk51R93BjPuIB4yF4ATQojPEz7HIDGgKAjHmkSl7WaDvCTo+nJ
unK6CqJGNEMjOXuFjmsaWmo+vNX2JYvcX3q0l04WQgc0R4NNeKpsshYaCw4tS1NWu9U0T3w7i33G
+Wav0qCxoXB4J1on3oohOsINqYYViMKvBj0ACCCmpHVAWVa3Ys7GiwawjS/9pPhdN2H4WytKw2oR
dETKdKfUrKodMJozoklHayF69rNFNZPN5Z4m64X9q77XGwrITKeqGbr3MAKYNDz6gwdtQx18h43c
XtLvbzAAfXWKiJH3yhoMHMk+Ba6FxuythtYza7JSeEQcTp7puWUOd2B2LcntAfjAI50OrjElCbnA
ehL39Hp9meLyriILlUwHMFPmvygbKBnABjT7k1QV8vQ/Ws6Se6PzG4qi6DRbUg02XrJ+qMfQ4OQT
rug1cEaBMrKZFT/exlUVt0hJYuY2WIzhyaFVTQxU4HUG7bRAM1mT27MHbaCvDggop0OyQa+KrCMq
8IRfDDS6gxcMx4kA7WdAfd+mkLg7RWwwefV3JflBQ/Kqm5KQXGtssK9mGdSiE5e+6ebiEV4Q3UMU
NufYRIZP9y+0khIJytaXQTvxSjYyv07E1lt/9iXK5UebHPlj9oNx83XA+zUBx+reO6NzmfKKFja9
5zxhbT3nBFy1YibRP812HIq4jGKwaXIRy+0jjgfX4qCi7R/fTjI1QM8q4N9+faEsh2bmsBbrffla
ZYqZ/i/daxLoOlArsv+qovwIj1OQ8Chwch45lOnWDPS/yqXrkHsYjzqQFAunfnMjWobTFjQmYTCF
mxnCxfRyE8v6o5EwcZP4VoGZ6HJA3nHHZ4CbdneQUHnrZB9hwk0KCM9yQY0w6RFi4w/j15nxnq5U
5g7ztS2TRVEC2PiNziE4XvHdBMNmR3Ya/dbvKTH8hB7WPMKsD70TkWV/25SMmh8YOwjTT4v3BlyO
iF5NNogBq+14Nlq99j+Qt90sy94v/TxqJ1eUu9SNZtUR5WXEgl89EtIEfEQwOz/4GUiXfNK9Fb/O
+viZnAeR4DwfICUXgfwhk0zPPRWhYQAO95z3tnidVJ2GBfQvLNW0TB35LYcSIUna1U7+JJB6dfUo
sumnQIVfbcwbDWA231koyzQLkdi0Y1nxLo1iA1GFjYDOrxhOHFTr2Hp+HMAAPrPLRI0Mz/XWRIqm
4N+U0x5g2sEvlU/VOb0dQ3EXlWdD8TW0ngWPyM/0hYa6AFEnnqpLrvfN0aOVsuXsvvF9x8VbPAYR
mHiXApt7qO5YATG8pRAowAXXuMsaZbc3aOqtWZZzJYJwqwE4om9E6z1r3GksDF/n4qps3hglu1z/
2gsnN7YeBhn0BshYVmSqN9oSpLjWEIBBiGstFtxhksnMydcqgOxE2q3h3Lgc0Mj0yQhpwNPv1QB4
CJNP29VlA4oQ4qBasNqSbOWOWqYaYG7A7NDYFlvC+46vYjDeT3wGFivkOvdGd9w0pcL5/O97niiV
KzmwYJ87WNhVUARouGTjjQtkALgSQLNhoh7UUKx+KiX2Z+ZMVIx6HtYYgMmSMUUuKOcXgK701UD3
lv0rT+D+O0uGGvz57U3p/aEZJgALbqtfA88JfTcyP7zXr36YFwg9RFA8+3PSatr6YPbaaUPdWJAc
BANJExoLCkE8OPghCkDPFwm+aTilnvLIElp2DYVBygaWOb4gHmSQWz7z4Vi34CzKthC51UGhrgp0
4Cg4mzy5WbafL86stqbD1KNT9UqA+/OCLBSdZflH2Hak6L4/yWQ/j137ak2H9Zyl1Bit5ZdlbM0C
SWprQgbZkvrNHXkO7laWMuAJentck8WxLX+b+/qCBVQQKlXyWUsSc4pXzsxzFjSyw+9fk62SxT6U
XnLlzSA452leFg0ggaSaybIy3d2zosP37QYbgdahc8AODPvlVkZKZu8FkZnWnBvNcIsxKVyBU4v1
fF7usDEmG1juzX7r5PXzlB/2Avx5AwXADIBOh45LqwC9btWgtfiKiKqdd5dGcTNEPDAbH+T8kJCC
prnmSNeCjBY9UaSFN9t8UYBgGmPOp711+UI35GP0VPcUL7mxKY3ybXRsmttCGkJkr9zRUwlsiGzt
9Sb/ck6X6/zb1aPPXhVML90qf8d/hgM/FUgleBbGeDLNlyLhshMAo7yRRhN+0x7IoAl/rRClP9k1
xNSB2pTNdx3DTTe68fxHSVGfaMbB2kjkyWKMPfrMZo1DQcjizvdUgvAxXW9tqWCgKq9fLHe86rSV
Z1IAGkRv5q0/tui+AjW43Nb6M0RluWHfDuV1x/JZcICSqQMCl3ObMF1VjjQPN7RYDOuNSv5dFQaS
AIKMhU5xpe9FOIh0T7Nf0uMiRiMhSxuo8NkA9AEeujwYDCB7R5s5ZgFQTtOr+vTq21MA224o2Tsp
Z5Ew2800NlFNFu2ynEll057BjttdfIOkcbJ5HjwnB8FEk6ZAvJ0vPGBbIpAtCIFW7+YpyhFmz+4P
/tNFmJUa3SviSGumlCq4YjF3LJQ9xC7v635KSZhg61fZlVQXw9iQ0+MvQVf88CCsUoUtg6TrvHFF
ixcwgwvJKjiQNTATVq5N98LwBk1dzVNs5js4OdCD40ikmJD4RTKt5xXmxvYCGpRjjgN/viLzV5/g
6pmSKF7vfoXJx9RGDIz4iLwRyZ4Fa/61PXdhieQfVtQKLAo5YLUfCmybNoo+VyJW0rhaRt7w8XHk
bSl+mdIR/8d2d/xJjF5A1vvQJcmNO+gS7T9Ecpippg/X0a8dfohpCm56ySnrun8wx9MKfGFqJs8i
+opI5GRcfjWuQt/Avuwv9PTGi4aOJUdX/1afUfTZCAqC4jgeniuvrvmMZugET1uwF7HffdUtxBJq
DaXrQELSM/RX8Pj88OYMsoonBi7Xz/3ZJlNvQPfwC+N4Mw4Obqnu+88/8Y/rtmhBvZidgbCkl7Mr
J+WQWZ5hdMak9fIXNtrwFVFG7Sdi+FVAp+vnx8nmJdv1s1apQNbWrporlDP3wpMCfHGZk+TvGMxn
PCh+fRXXOsCdbZP5kWLw/2qaeirluo2/7/JOTNGbvefexFC1s1WwHwckf6+vlhbQ/g8lV3///WLh
IEmirZr3db+Wf184TuOi3vP5uhIBmX38Ex/yzv4c0whZW/6YsrOynyxvBLcDi2lKkdOG0Isy2CST
yfBNCGT+UBSTp2VMdBWAvUH+s1D1JJH2tq+S0EqNGEfT3PbsF3LhQxtpcizuxiWmS87LOEiYd4vQ
CSoA44D8h4pr8zeEfE9Lk1wtlTQd4dA4czr/S7D0RQ7I7bChqDQycfao9V3xvqwjhRJNLzAPMBrl
1wAEtdUy5H5elWZUs8vGVlYnwcs0INUOBAel5DooFxk9XXeGNfk1vv0BH+JgTeEc60OwfLKLeYJ5
Wtx2JyaBCtwNaz8zin0ArpGMh3W7jtSHGqnfgNILdduglHRRNjmAEyWt4U3gOBbXOVQIe/ZcnDql
ptzYkn1s+gCucqnacofsZ9k8jsOo4trPVxemMAK6hiut3e2iwIgLLmK1pR75XqFS1N5bkjBAeU+g
J54NEOAnXVLAaKjBVMWV9GfQEFA2jF5xd/Xxc8k7HCzRffCIG6RW0pxacAvlZr2KBd8wE0kNkaCv
BO7PVrBWGFVTRZ92uiurbVml83YuaxjEHsUw1/9BqSENagxAqK6avP16f/7osSahJQtx5Qdb2VHK
lM2DeeeCR3cr42sPByhaApwR6GUoQR4TUOYi/2pWn/Lj3Jz3dH6Y+ebkBii03hbCaU91u5cNT4Z4
dgevmZKbN3q76763LObFeAEqRSDKv6RmG/5Wx/pYl4INpi0PLgMfIEgIuXquq45S6xApwy5+QOjI
nRd0U8f8zo7VzQNiYm82fht0TcBsqDUNZUz9B7P2/us+DFXJNQhiukJGqfSaNohcHUJy4mrDignF
aP1cUl7ynFxF/4mToEffC/U6LlCwhVbOd5wSxc5PQRxXBTM9l22AeqXtINTteVpqOTwOEbs0nE38
rtDvt5S/8lI99rp1eGsLH3NqpxZdnMIa+Y5wq3kLzoLpLh2fx5ZZB94unnsxxhdopXS9PtNV358v
rHNJrH6J76DtAWpbG45rKEKcrnbuvKVI8ckcn3Qgsdb0DBe8x9fFmzzWn7Upl0yP5UpswE9Nb3lq
tkq6JNUAxj5mKAhYXwOssuNQLH6TFKF3vk4p1zfKLRVu7HZCB1yLWTzxicvKF4wbXSfDxoMchbJe
GgP2uo7HGt/Toy1VUC88VuJ/3gnVfNJZ4dSUKNhvAXC/omFqZjGAEDwWkxYwcAwne7xgJ8bKyIH5
305oqISH9s8NpeAY79dfEomgUSUw5k2Gr+3TTk49AjXpZcqKdWQ2V87xMN8t1aM9busnXat8VSbd
ZWRa6udxFLIFqa8AJ5k4Fl5b1hsUkjCyrqj7+oyAMe/dJXqZgLpon0Q3kpX0LtKf7XBz7yBl+JEG
qadd/x/64cD+OrEG59b39FJhGMwSCFEvSOY9L84NJ3Y1gZOryOZqOa7nka11g0oHk+7W56xxGDQ6
WkNeYVIUq3Dk6WgVU+3RLPFUizO6fcvTOaLq/GfWqOViBCjDGvcstr5LFWqGFjQHbB8AU4t2qwJT
YgAtQTF7+0oN3T1HcSx2T7QzB/Yom8RfhhJvRqk2Fmi5rs5YRbflRTxs4061t+qmOfAZotwynpaS
d0V9mXU/ao2bXT6tVDZlInSn3NWWgbSVOyYLHLOFLGMFELjR8Xrhi7c4jVV7wJsoDSuIht4M/+Sc
EA9PDW59pI3KPm++jrmtpdpTawby6ekg1e7jqLAmEO+YcGGVHH2CUyz43AZmoljo8Ibqc6EYOJDJ
k3nP0o/dwhyQ7kfeSBdVwDHTLu3fKEOcyEDruUbqaNK+P52DMpHV9RgIwsnoXzPBXRCYwRicj39F
jJBlMQb9XgBUsB1RiP0XAsVhnCh3zc60voAv9xLCF3GMav/TnCnrsCIWZEj4SY/m6SGxJV9ciXrV
y9A+LjabCjSKWurdeTZB9CJqQQyLZqTmwj5RNmVtAzB2kmEeUM3Imn5x/77F+BayzPGCLl9WGfGR
dTX2UNkJ3Z/t4ScPD2UTJSA1uoLBF7L2rI2L3ZawPwBEXQmet1ngSA6EA6sl4546kCd+zTPJRTBY
+RCUrrfDsbdsdoTI7NZfoJtgGj3Wpu0T+aT9r5WaCYAKKyrdl8CG9CMZfHSdsPAVBSf9AEZ97lKJ
bo1QIsVUdK1o9ZvBg8JJ3AySRwPcPSB/auWSB0/LU17sNWe7xQaEu0DkCT4K7NmiGIYOTO4DUtL+
rZyoIkKXClo41V6PylWa8VWYPcd+xb/L5W2NuRhfFjTng/zdzeng7ksUZ2C104JCLtodBqIHq19o
ZQA7C0TQzaBiAJfVm4o1weCURtNYxG0USRNA+p4pvBmTl5DxCn29/T/ClnCHV2da9Hm6aHnt4iJq
/Z4OWgWPKzQ8NUDsoQbtWIODfTndoTa/BRVXyfjqH2Wqx38e346IHK7c0E2k7xyGc2V0li7H6sUB
Jnv1MwN0dHLD3CV01gfNbFXleve61h8/RyGZv1vcnuCIE3lueU9Jq/2DAcQBKZ9eYDDCX3srQg6a
Nnwez1z8YQGj1puO/Hppq3/cyVR5LTICUNq1M47VgjMwn+idjAUv3Xrv9j2tbwzHsCZGlaFdEZJV
mjZTGIpTuh7zsCYbKK+WZ4KtoK12YxCScMcW8mgJnP6yqil83mdCM1puftaMkdsuSkmRKcSe+Zao
Q/gK3+VUNQd02CxuS1rPXZWkQzPF4FH5j/1sDHanaxvr/wkQgSnCVoFlqjwDNsvCj9NpDWhT0feg
IX1ADANxu4CinonEnor/NHyBaxQ1uIER8cnYDd/2HDIITLpKGrYJ9CDEjm1/b7tO82gD2N/ViVrk
24IRKKuGR1FdzHEYefYSGoHZyoyBWGS9yXxwyo7/aT9hGVjxbit2rm6iOtHuyBy5/fYqAGrgJ01m
nML2WllDAWMgMtgGqgU7TlTbQO7d/HMtZ01MEInW2Ck3Rc8ahnMdr1c1roJ5jn6aKaDYWimOUX7Q
M8zM5Zs2F0kDGX4zNlznL4++2+GQ833foFszudpTFtPBLjHDkpy6s+N9lviM3z2FG6luetM6erkv
EQu5lmaeK2INof3pFux3BkRoCKcp1VnpmfSpRIp+chM2t3nj+A+Fm0B1FL3egXMIEY1DqDPPuI5r
pUlXd/2LX75ZRnesMo/JhhcsmO+AlteTkAQpU8IASaASshWrQdxZ7BN/+aJ3Zyfg/+oXT2U1ZVvN
DFdougiKuuhJzBB8GtnV+JcRDoAWVw6sLbkTNuNS2sdgAb/yd9yHO7BVYyqoCuf3wLZrmpYOkAEr
drhQKDfahsTxbRBN6s5K2XmdMnJ8UN0+BKtQn5wvbY4RztafcdfDCps5u8IIz7R/qHiChbEHDOeD
yHpAqzS2SybsAqntqn7vjknx3Fxn/ux/fJEY9DB83ZWBoEqA4WJP5LLYjkgQUEdu8LnRI9aF6CeG
6LhwHpN+WegvzbjdlCEVmb2p46R3n0oTUBfuvaZZK754kbopIW2u25QlDZvo0olrOzn/qwOe9sfN
fMsveWf0fKVgGzcu0xPjpNAeAuJ/elCo5IEkRK1KgWKW4fukhJy4a/mUepUsvWa6MW3FHI7slbCd
xhtfjv5LecPbzqMcxrmCK+ZrKcUu/MWiV4mc4WfawVh10iooGb5viEeNSGuErmeot81o4uloTLok
w/fkOg0Talks5Zngt50/4baGekTmp0q4Lbw+XfxpwFQpD3zbNSr5qmV8FoDpH/mdENNgeO3u75wp
SWcX1YUyIHnqMBfWACJz8txT4FQJoW69OR7CMBAI9oJ7zzoT/4ZskYU7ThecNQnJrFrdXizY+AxS
i545iGeGzcySQi+U5RbW4Io4fHKC3qY3Qgi29OlgJHLWBHiDgeAwHwbu8djGL40qmN/9l1y/V6HU
Iy4xHcax4ZNVw8ibV1/eHbIpxQy5uQoempyTNQahhkdotBzo67IngfOygC/OY8kM8Mv4Q/Pzcljf
3ypByI2EL2gPUC5VZws8XqRz5fJHXed0ivDiFij4PjLLNxfeaoA+xicUud17FuO/dcpwFWNTV3fI
GBGEaP9kQBCbXKnl0xXtnMKFmBWwa1gf4vmB40UTJC5kfCdUGPbLs7PShHIy0lqgMi2uAZ8r+nv7
oqpm1sG/Cp+Bjk9ktZvU3yzK6FeHqIwvbT5DGOkdiGB0I4HJ0yvTbD1Xf1HgVzssDyLtCD4SekpR
gGwbPj2gH24oadhr9Em/jJjLD3iZ4H1FgECkNAXrQ0UAPiw5Xkbzibnjyte+xZHnqbzzGnk1fesH
w3VPXiuCz/f2MJHYybSr7INDSEzQaztP15b+Hj0AZMhfwUoINTnxD5ynwGFbYzsD4pu2NN8nPnH/
gzZcs3/9Of4Yo1xhrMQrSS7kGfgqfb+cBVQ0JnogQjMjm2RHJV/sQG1sKIh5YjdpGkIQm45heM8e
ibVbsNvOxThGjx2UE3FlZ/or8cbR39y62F9BC8KBXOcieAiIPLnMM5nylKWUPcBmaVE22UUR+Wui
fL4yizw9h14JzBxxxmWSoI6Zn8SJ0SNw3PGAwuLsL+RXg3S9D50+Qf38uEF7x7+PZBdCsLy2kCnx
+toKPWOp1J1E+OwiybdY1ywiSfLP9Z/ngC3EbmjrwenC9NjEwPgTWW9THtCauveOMtkkbv6HhsZZ
/g4Fx+NeTnMBR8NwdTXxnsBTdLemjx2mrUEnUzfGnWIygcWL1Lrmk3DQFaJQvZMiLCkyWCOt7SEv
lDXegeEc7SgUjyIMH3/d1ZdBvc2rHll5uLfGlcUXRPAsR+BCuRUh9Mj80Wm/X9ioOElX7fZ/WgKH
OwX9Z2qarqfTwlkLY+IO/U5NDAXDC9PgEzGr+4g5vuHX0gR7OvWd2fXdvOm8a2Jlv1HBaKpP/NWp
S6hUav4pu8SYB3KgHihPmO/MzXvxV9s7bl+paFz49B9H5jzOPKN3rh8ZEf0TcxSgLz7qiXbd4MTI
VUvqQkQAqhjtKWQMe0ifwNF8m00V2RPGp7YidiQiwjBv2dzbBBuo0lIa++5vrUGU+U7dpvYXtyDL
YkhyamKZ2EkKTwuwujs86HHLbQy4D5lOgCQvdqkCxIBKfQ0HXvLhGPkePBf49VMinD4RZBEFaxFw
KIOXU4ZCO/75auW7ZbB0ynyPcl4AxIKQICZzZEyulzWdZM1MLJLbrSi7teTXnj4eBxyGXJXk16Pq
1OF8UN6Vl54FSo7cqs7wMIagsWdVDRh2Teuq0v70+UpIvzoZVs+dF2sP3b3FOaa8ugdYN/tcmGuz
RpEi45dsOAqVEJWmg5BRFfHYRMByjOYIalqqpP4ysNtVQTY9LsA7VJpELfoFHBMDBN7mDRnmNr8G
wi6tQiqSkVAjbtlDd+tLKxZZP6ZjAynjJIRe4cqOHhglmSIbUfZlCRzNK9147j7e6P+pnwp7ROM5
1f7rwDeKYcWTpCAxTF5LLSHVsD+ga3QiYAi58Z8P3BysZr8T4SlN14SyDb2EiPs9/MgJsjtlm3Al
9zcD8DdcXkS6Yb2l7bgAQTS0c6+LwO+TQqY61GcTzDrNdVcrCwGf++aQqRJ0RVaWafh3yGKhizJ6
QTgKWpwH0wIfIYJkn23s9PuzjMrfnsWvbiggvx00PfIlWNsRJO6JkfBtTH+xmR0SWEzPWD4KNkr3
g0Tg0fD3mJspPvq7c9EqOerHkTdLZ8/GtGSdbv5XJWrEdP8efvSElD+d7YVWuUDUU/9rWmOR+oGW
Q6Kc+3G5wFU7wk1/guchs0+fnwQtxx3/igC1PZQdbHLq0jP1Ss9Ot4MpjLRwCJqfMn+TnFYgKErK
DdRd1uID1JRkV9bCdjFLi9xznV/0SqNZ55pwFH5uDDCbAmoqYCw6f2X0GEkaaNTbAr2Y1HEgQIPO
1Eokl8mFRXtXziMLKc9zqEuYQUwNbKblY4U5snyVMBEn2MtUxJnvsi3c8X8FUXsUPcHc07eodXQr
rnEkHyhxsjb47hL6EO8ZS2+aKv37TPRr7ohgk8aQFe36EaiLvns0JnOyJEthRXbO4eU6Zvwkaxy0
dHx8InGO1G2ORgxGH+qq0D04XPSYAZRIUOJUhRKEVTJbiemRgCMFn0DL+au5ZyUAVR2cYWzHjwm4
WFKMpbrD1dmCYqvOolrSUIpjkMUCUbkJ2j/CCGbkoo8Dt5WZ8JMj3zrkZ7vfgn6TsZA4ATi5evkc
5ynhOPTXqZNmQ0hCV4xRRC2ZYwJl6LDphfxxGBmDS3Wqj7XSYNeFsGt41CNO3ER6Az7FcFt4SCue
oxWZoCj+5mYhJsxI2Fo1ywJlsNjyRcmZHBf5rgDJvtVo1FcStLln7GoJn2TrT60O/0lphuNCnze+
zx2A+O2yU+zJZE9XOIZ+ZgLN85gRCL/l8+XKTpzeSFNgZtzcLOCFAdQmuPnoaOl7ByYJxlhrDLlr
oCPzaMK8NyUejLgM5az3oAqYoz/R5mm//GzbmZ37ftfb92hsbi+hHn3rJNxnkxIMtjw4VB/iZhYe
3RHiK3C6gvfRD39t/DBuFhV/IZ+US32D1CmqOXd+26zKl7CZVKAw57G0wDbhbxrReZ6hv2MsoFdM
L/Uenz+FtNB803QykV34vmV3oiybBzwI89kBTW9l1c7uZUSDgnpvFLo8Pb4pFS6fw/4H+pkcSfGt
EXREGvyZ/Yc3YWeO7WoW5ijveEEwzgVHgmvfhXKcGtybJ2yKnNR5c4uK3GrqSrK4mas0gjnG2YOp
8R/lYyrMpKX9jP92Bp9yxXIJGXOzXV3vHULCv1NLPh2x6VtbrURIcxMY9lq/aDsjAVkY4HDBQN7J
xNGeVTLayNUk0x6l4QgmCM9iOQ5MT8Rbh8ff+SWbWo1CsynF8smhTyAIcYlAWCBn3gy+7ZhmiZ6j
CneXFeEoeax5GYIxDKJ0S8JmRNQgQKnmIPgQDKZZGef19+SaYfBY9Hp8/eI6+o0fx+08b+A99qM5
pgvMYVNuQ/I6xXnaek9TvTb7cDeszi8NYkU+zrf/3gYqJOZQsT2NXs+BwdG1AG1Jsdnsy1ML3O8y
Zd72UAxLn7ht+KQFiNpY4gOl8h5Pl5iqOBXBTOeT9MYkQB/p7LZKWzEd/HBMq3wA4Iqxlvbq6IkX
FtDTU8y2DhfJSUnEyn1TE4DS3f9OkGxDfFDHuticRt+OTsM859ZFzpEZbJFmJBkH+B2JSnH3LOxF
XyoAknxJKPX3/rCRbFKQ5jvRejJiScSt+o1gzJ7TDEgp5Fr9ExPFOVpLt1pJuFMcyjmjdYuhPv2q
kEjG44MtlIZsSTPFUeLbEhEWoXTZWMFCbhvVwcnrSOwMi+pTmbthZpKSrIpPHxcg0A8KTgttN6w1
XOlEZyHSoqeyJYyKvEhWyE1ytx+PsxLr+pZWL7r/G98jCEPI60W956IfxqRkP3+oG4edGbzNJhGK
jKUQYMd3KzGYIcJ40hKA85FkYG6UWfBbczsU4Z7V4i2Vek9228fIIUEbtehpbdyPxrhz+6FKpffp
h148fQZfF//+UEKyHvW/uDUE0NRL6Hq9MIMxztyko3jCjz91IRD/dTB+SzXXhnGyZNoHlYlZBhAx
Vl5RPwsGOuDCqR/6gMATUC4zyQWY2c9uwEb8GF4CkTPVKSgCAFzVHnANeWet/POm6i9CyL6cvQAG
HYiy3HsUtSqM23flNwWnedrqJ/aFe33Gj7iqqQmVgIz8TaDfdNWIAM+OyATe8cbnLkxDctDZK0cD
tXuyVj+RqlQDbd6OlReS8NfPtqgwjjiGFmWEa/3R72LW5A0+9U1QyGr2GRJpT6a4JMfuJRqbqB6U
HPnp4z84SZOOdEfwXEpTtdWQ9D6ivCsCnB2hnu/M3G4TeCZCXniD/l7xXMnL7V3r/+B4Eu5nFovI
HtAkyyqo/LShNa6BEr2on5bpseWuenq4iucXuDHkkfSRkyNAfmBMxt0/bv+ZrBiK+ReY4AMh1PsC
tqRoItzdJVEDUa5ONv892e6s3MISXXDM3ggtQm3Dw2nqZal9jlNWs2zpp5F/9O7jW6/NMcOOy9nm
1NmP43aYFoSKhBv2ljt6ofgn3aNkOKujdTs3ffOva9xhneEIf8QtjMfM+A2XIy2VQX8quEbxJT7Z
Cl7ON9PEmshsMgqC7CeBmNNrILs/S1ymmgv//OlKYlMRKhonrZorwJWsKWL5kHWk3jydCNHV+J+V
IjJmBrq27+NlMNcKGLVk+pYOh3KgFShR+1TDsW+a6T0c3FMeW/89AGjhAvGZKmC4swNZW029J9QP
w1mWEMeGJTGSSRJkuxQQc49H8IVEk+HlxHPNyBsznIm9XN0+P6O6UhjlhAOPMcELGfy2VmM9VE91
lOYkHYZZszzeIA1M4dgkY3MHQXcgdY5fYnz0dQ2xYb7NCyIC8NhELl0ELAjcrg8jBSjxOHzguUrX
lHTte2++3h/n5zXNKiwpbecv0dUBPTZkGFR0FrYU04gHdA5GllxZdZt/lxkHoPlZc2ajtXJDCf92
FAkuLUjUqAEMPkOI8G3GbmB6YcbVuWrKtim10lkPLyi49tsBqP9KeSQ8VHYl5RjzESZUKRERWuk2
cyoy750RTW5iYvLXduEcojado0+hkB34HIE6hH01CiUoCdKsK4wzvjy6AuqKJXYCiXgE4eMmtROa
7Gr816VRA6p9qaX45CgNGqSLI4I0ejLL2ffoAnF8pcPI6C/JmvLkGF0AjLsP/8pFptDxoGk85b2F
bmUwU1vamNqqEyeARCghBeZqwysCMNir/XZoz4QGlDQGh7Svf9sK6ilzpTjq/QzDOoNqpD/73xyY
xObUNj30nnu7rmGQh7NnQEaNoSLKQ19seO1ZOlF++AGJSh4OudmkNNcriJ5Jys9S4jhk4SyzFK+r
IYvNGIvR2IsjVkKP1rmhbBnXcYyF2SBy4g8H2ww/mvCUR4ZWILQSToyHelxc5R8AbOk3mxgAvw7a
WrEqF5hWIYiXaDPyQ0SXakf8D91/ytHxCW96hMCD53Bl6ZxwGUtm4cebTCeeY4KjXzlFXVueNOmW
S2QbrUYXNNkA9JnXzqletL67CVSa6OpQAnwh61Doly9RcPepvEonaICaOtM9goiSFwLfJX8E12lz
XoRiG+6EtfMWdyV7l0pQDT+/zF6DNM0gWa3gBhsrxjMJtJYpM3MkvCjYsDxx55hWFJqBWZD3hg55
4ktLyx1IWw0ZicNC0oS8sPgY56qqpNszBVCbw7rc0mCFqVCJ0lqOE3mL8+mEdqvGTFqlotMt9jD9
Ii9f/DmL1K/He94HTWFUPDOa1WzYXU5jEop5q3YwvrA2ODhQnlVcOKsShzdPURDDT2yz26ORayiT
+AlMN4jCgMmocTp0wjS7UQF9ZF5Kf1TTTJfkqWwwkIEFGj7k2Bp5zsmbePNW+ziZaHzMtV/aA5wL
9t8Ns8M1GqGDsBpwis8E6/txaWJrO3lFXT44xXHW8zf2Gq5+J5RWlrUhupnN9wsvebs13r+Ccshp
bayAYYwcL1vtiV1xRX0bhdRrsPlPwdstzZTXjV0ehP2Zv+he3YmYjuXlpjj9JFYTN4uWuivuHpQe
q36BPpj9iYkprC4X7Wlq/GdCkyInHr/JZ4jzslxtHDLKUZKQpVC6DUt3Oypk7ZQHkUiY3lBl8Yk2
qcyBs0JwGkHgLDNrBuuRWoDUpNUwIxCIrRJL+9VgWTho7LYGh+TPov7rKdxkBYtbwdwBqByaP8oR
jVSOGahSpFAlNxq36x9IC3lqYAxonBN8HHn+ucnlndtFo9lqrHqxuGAQ1cpmiBKAjPHzOQMYxz7u
lYxFDbR8WqxCozFGKpI6ctxwFrr4nCg1khc+Fk4GARidIqk6O/g6JjVQxQvGnklf88io0ksuRTlV
OuU4MfkusX0LTSQuhYcLwdMECqPErqNwxs5R40muJj2VTp4KUya2JZkLkaikT65m7Aiho+yURaZM
aNu3RdZBNl37X12XJMSVKxkvTz2Iq0/uWepkZUHBOEHV5yCnqGCrkxMiGJEPKFeCWvOAti2gd+Ru
cNKIhaKJ6PB6Ro0SdXqkvfjpLw6zcKd3g9Vq3inqhQQr2oRgIPh0pjfuXljE+DywCB8HFa1wJJGM
TAlXmCrPBZLEgcBRYKWzuvoa7UmlpTOJcytXU8PyXralZ5inRjGDFBo7LsnYNDI6y1k4VR3r7vjc
8AlTiDnkzgvOHA11+dpCeZK8sB0dhxUsxxo83rmyAU9YBlMD8VhQf7+aNAsUf7IMRsVV5CyyJZ9o
mZXzXmlpJt30q/9iCtxRZYwIY1c6pN8KkU3PhzFBht4zgKFXRFHL6cLTyEr/MLMkppH3A/gZJeki
HyLIsjhPKt5D4j4hQBuoBSFGnE7bj78M+boy4UeRHrlRFUDkdbIedagU5kqBwlVBEX2vKKLuHNsR
z+QnrTxd/+c1NezmUtkhCNuzdTPudr2paF/4/om11CuhovqwX/mjteAea1pMSGGifmNgQQcMpHmO
OhN0ECU0cAKXzygC+7IRZyqzNeKTBZpuB4UEzuC9m7xbeurjE0aASWpON2Edv0j2uwVlqYU8Ag6B
CU66RPe0NBtqRA/oNuZpJa0QUhy/XrEqIAbdr3TqmBWhT79UfgYXLEwqcrKnLRkQiqYWgfUzfQtZ
xgieeabEMqs0yiCbC5pXZtT2rSaPgMRq+6oYESm0BFBpLkpWWtGvAMbtMi+PNJe6oPROz6TF7sRm
xiLrHNxhDtdc/+UTeB5Tkcr7fQ3zP7y2qXRC7MfKS1eLONaAlBxq+RMBtHYkyBl+1cbYtcu7CKeG
O/CPBc51r3x6ep/s5WNg8vvIijxoYtEl2IacCHHY8v8EYXp7dqpCn4FiRf9JEeuc06dzCR3cs1oe
n1qI/05FISrR+l/fJdz76CizGDv2pkVAqLWKZFB2HlzqoaGWm2l3B2+3LGfGLpkdPovl/PJFdTJ4
VpXCSbsaYzeuYgh2nQNSZK2a/s1WtrRTwdeIdTpupKPgokefNDE6JptGr4hU+5t9fZ5hCCaEdTWF
8FgkYICdTMVJDdafi9a8SUMhz4D6vPkonNXeJ6weiL0gOTQedg3lzfprWqtJZOK/jK4TBlhv9UxD
qNC5t53GslldCajbb7W9QfzqB9riI6qditOE82qQMtpKWYTa/sTbCyuODRPpc/k7phvTpFtIte1X
BTcm2Y5S+4MjebO3NScn2XwZ0ojbYw922400BS6eFdSv+8QnOO8KDZmZju4UgEKrIDayFiQYfEiL
ng==
`protect end_protected

