

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BwHHaRYHij9TGTVh7NqyF6fPKvSJbz6zXpDQ9T0CSRjM0Tr3I2/EoB+qBgzPRFij4R1VpNLIhF/W
jnZk7ILw5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EoffIvgX5Yh3KSkMHr6Fb+Y16CSwhqKyrZiel9vaFNUa3EtfX9ml680qKyH6k7Lt+GT7JeOZ8tsv
GeWg3Is5mnBMAsR5XkmKmU1Mf0hiU70CtdaVxbMu+l0K5NkyBzps5GWZFbpBi81xyWc3mZBrsdOP
SKFV3jiPDhzIXFusLNI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pC+fmAQpqkr0vqse1A8SFfJnAErWB2cTBoy5W2fu+Qfel2Cgg+f01SLqdiCqUwM3sdVOYKq280lw
0KlccFWeISj6EGy+UhrlckR4KPE0XJ2GFpTDwr6dIxS9OpYPDM1MXlxttLYJRqT3qA2yEzsidST6
0i31grVO6qNsjmpW2d7uByo9M65VEOheITjyvjEpcaFShH/Xo714T1rUj9u+HOahJ+Y/IZt5BXf5
ifgOOsFSC4Urhn+vw7WBdTykWaXAuPqSgZ+BAzkf1tn2a5qwxdC/nJyffVluJZjwqKsS2qOqxdcW
lV8I6VmHkVrsFF7Im+SIdtLtq6ajfsK+Fu41Qg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sjA1wOpImDpYBBRjnwY37zkJTSoQvS3OSqKSHwre5fBAKnkrgUJxozoTE8i2Z5d9g73A+Dh1Khan
8gYd3xbR7Bt78jJM+PFuUbVx7c2wSRcHOAp2KIXVLTpuc4ycdBn19YJhb2UIFhm80kkNGNgavUsF
mOqFyOQQiDU6WY7JVI8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yt106ecWVBUI4xOZZkRHweGkZD2nlI1jRN4H6Fzc3EkfIh+DLe1c/sY05LO26DhXbTC0r7f3V5kn
SKvkly14VHuR+p2mt2PXxY2kZUcL6SEF75Sdud7O3qeyYyxwzbLXhAk8rv8ESHYXdpJzGlAIPVhc
CV3MBlzutogOhAPHHcbRbukDx/ONHomfzueq+JuKHmbmSP3Sji52yPtcq4iLW/WcLghIBdR8EZ6j
UoWFDA94p9C7hEbP1WkZCFdBxukr8LSVfTsZyILoNCYLGaM4SAN+KSvY/r6FcDftOrSTK0VkVrNX
POMgLw4WpJ2xpIx+qCPH347wGbfYnUgOpgfHdQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 39232)
`protect data_block
H69KexgQvCJ7NWpLkRCm0VRgdcKz3s/qMc/ws8ErUQH7U1H2VIxLyZpLj/nW+GB5Q1bsHEZOiPil
w61FIyZKG5JNBlP7BjpWgIWNhC9ob3l9BlFPaPCULnuzSbUIOpPHTivK7PrCFCl5wJN5R2G1LQdN
xvSlvpO0A9B4e4LLDq7fwBeEvhJLiUopr6mPeHVBjr/3p2eY73Lz/O+ekH8/7StgoBzQe0pC7J2S
0jXZSom0b8xjXU5rNCHJ+5RSamXOhc82TN10Jc4QADzpWK0cnMwbzylHXxa7g9CRCC5bMvnpydlf
C3ByYO7wL3CuKB+gpTUIpL5Qj9coNfxDBBKvBBEuM8OXbYMXzbgYVszNQRWQ5xaP7hCh17oeVH6Y
Ocx48VcoBjQxAJbDNdNVsPnxqFkWdPvMeDlyr7HAxlbEeErXTXmgoifYUVKkxNTHq7NqqkmQaXsf
y6kypZc6rHgrWQwBOm8u1Qm6vMqQslzF00lKnDz+0GJwUgiNigDdaZL+QMB1KzavE/35WD53ITdc
Jcpl4NKuZUk8K2/JoPRNAmOhtTmyWTpoWGGhS6NGx9Bl2Gu6FHi1TS7AKKlfAHFLixkuQ8Nk6ohM
ZLbFaLvTw5h3x5HuxydQw1KSB+3/XNcX7A1AAJdfFETIwjgJTjl7ZjzdAiYEdeaH/bgLaVZuzrzv
vfy+oKUcuKw7fzX/aGHmisExpBRKjn5+3HDugsKTrUkBPv64CsU4UIXhocAF90wUFDi1FQB+FB/j
RbBgXpgvkslXAKH0Sj+LdkfXkH4JYiKWpTa5TrUNCit+o1V5ZYWM3VQ3Bst59VhYybxOqWshtHx2
VfOqU8ZRGrLvoOWWp2R0+tjbrkobxXXbBlxHWe06ZyriZKaSNEIrf6aTk8e4VmwkvEaqgDaXLLzH
Maz13mIkRM4BpJzhWC0KqCaf2TWnYF5CAOIFCZ7Z64i+CN/cDBFv3Jv80iv7rSDKeu711oozHs3k
USERV3qjT599xB7TaYeDbSNs64SpD5npE+Pkphdyr5cDTQ3miylXd7lihsk4hQv853QoKd06YL3G
HAskv5kWc2uMIYg7e4dtUfeyI1csxzAEOaIWFFZmgugP7f4qbJCNhOIL1HuxyUH94SB7OZb5/HZ/
bDOLPsBhI2fF4+NEe/OOjIQkWcPcN8iNBtSfZCqhQWAFjmWG7L3Y23zNvF7+VTYRw1XReHiQohwF
gNtpszYh5fkw6vQO1aaFWKQHc2a3qZEYXDNF7YAFrL0g+Ccjq5a+BVEeQRY0fOTig8BIHPZMXs3d
ZO6CFWndxbDZztmUdi0epiKIoYYUThkdz8DJcKSR1tTcalxEIO9izDt7xwFSHMaOlwGViXuTzDi4
cyaxounlZ9SAILoaf+rP4QVdTIiTexoMupGSryv/Orh3SYtP9UZBo9SXU+0MPP1nFSuefwGSImlU
YtEMucT+0GbbbnAicWgQNN8r6gyBuuEYI1N/nq6siexX+pA7ExnsN4WoZZSqbUF4+a1fBg6/MXk3
peXDrmdBOz0hTycq8RIiOufwazsY4IM/TdAPxf18co62lLbWMfxuuk006SZYkyggn0LMiGnNccoE
XH2lkSyJjyhkK9Jt5MxXB92x9iiMh5P3F57ZVJdKq68zpidPkl7XfqkpB12fAj+9nwozQjMd/LEV
UfW97uxPT01Hvz6YhlIkD+hTj8b2KhHAf9x80blt6pTRHwWsSU0esMzgTWYXt/9bpYCosBz22v26
Og7ffUsdqcK5w6eFlfIbk0QS+TEYfD/KfGjveXTUg85f63ncQLr8YtS3RjPbrew10elS3ycuJ6TA
F3jj4LrTb37YX9A+LyzkKwyn6LYk5Wrq0RUHVOgMulcdwz+a8Oi8/JEouIx/4NMLhV0kvfZOEx84
od2byB1TfsdbqoYlFAz13Oz4EZ3lrGHE5IoVkNd5EVYOozVYu7yxlw1zJ9NPiVngpLOigaFhGEjB
ITR32ezsQC2O4KSHHksLGOkI2CEjFPQ0OECySdDzu5cndxGJpyxYYhNgJFCipidcB+KinQZD6Wa7
NUqqLPaS2q7KXxiZPYZHdW3+6YpGaW3dz5YU25jClee3whiG4pO86jJAuTzULcPSuDaIW1Cq7LZi
lCbQzdAOjhe09wWnpFilSA1pMsjx+mHBmQDKEt4UJqj6z4rluTZjeSi9fsnPPuhVdZ9/QBW+snfY
dycBXJ6MBFWET/NWGPMxuT49LaFy/493T+VximL66bfuVip6VUEU7lRatIDT50n9E8BBsH9dcuTC
cmgf1z5JLLCN06BFfQ7fqMkHPdma+/TzUTOXK28qILKSx/6xLVzSTdiOhSUhWCjgTKWD2WpSihJX
x5CX9j1fv/SVCrDUimbOQ9+U0PZ9PECbXRRwXo9E7AGIepQqmNFdiG1aZUpBxlysWDkeDHO/VklS
d1NiFoM+Yo7yDcmSEfNhYJ6ib/ylzjRpf7eoUVLJhHp7Tv8B3pqYyxd5Ydt9Pi+gu2CfpHrgDMmb
G+mdvyD7iyGhtE/69QrZWOS/8dMvOIGj2ECYDUJMQY1+dZVSwdAcn8bWKZdRkeA18U53fqwdxohn
J/+IMb1F+ZFmUBeD3rkxKCdiWYar6Yl0Qb9drhLC91039nI3M+aDiPxIlgupCHgh48Sr0m2HGZBQ
4oG/dkP+axNyvYLo2ACEdXPuV6E6BqiJ4vUgu55ppt/zWSy7kAyu2ZeQFO/pz0IZE3ccwiWjvubC
jDjkNee5GRw6ovlHzA3+eD5ka4+w8KlHZc4OtVKgFloGisb1DyqXE6tlRtOp0hr4XvMjATYAL4i2
BZwb7/cn+dkM/2pc6aE5hWtj/ZfRTXBgjrY4eYT3NoRHfzuIzekZMjEYFOmnHWwiPM2xIWFlxhRd
1Ijofi90jts9AwcIxmjCEBVdSA5iVg/E9Q9ROr4N27EAqhIRAjveTc0hUSHV+fOzkiKxhKHDyVuB
h3ij/15TFhuHkiyw/Cf6HGSYduqLXEnAw2ab6/PcCmZJ9CD45YII1xmzGHdYdJld2vLuyltIuUaR
BsUEvCSDh2h2ICeuU0Awu/AKv2eXr/mUnmuFeGaT6Lbx3XnB1OgFygQIDVTK6Ef20wUcVaiz0hUp
y7idehQW/8+0JVScNhVCgA/YtayMeSis4ZiRSYadcXyvwfI5QYkDn73XdePsLuL18c8p8Qm3Xp0y
SFq2Yuz2bOEeHAxdc4RztdUt9TbSMC79+uqtQ9BJo5DsHzO9JXE/v5/b8XbXxkNKyrAzlauMb7JI
MILmob7pAIyzsfNGFJgwNaDmBFLpeT15P+x+egWMcpoXjlN8OtVWnrBfC9ndnGIStHgctzyFrL1X
82l/DFa2K2lFoiSTQ8rAMj7o+qX/Up4BufLOheMbljP5p8OGKi04jGX6L3Nrfmd3fkUrFI8TMGEH
/kg0w+TTrHEoQIbKDIhAnZRPQ6jCeGOsDRM8PfNmWNWl8hJPiV1rzRHHNmZzF+2GlYqcctzXFI28
a/tDcR1OczOX6h2iXs/aaAUm/gJXMQAGIfnGUCy+RqJV5w4c29G6db1PGI76nMWtlOE01ve6+PpI
sLSxRnV/GA3iLXrAJlJt2TqHIBq+w93eRVsjtha3TCr+jZSceiyFBi9jGZcpiQcUllNbdNSnXB7e
4aDIHXvsbZxisQs68vfehjgrIwdsNjVhwJRtk5MsJcp9blmqcd5mohFTB9n6d+wwJjOfc1gPDB3O
j88OpISC9bdqfQBPlTo5AVi3PXdGaP/ubXSnqKqrR08NYWAs7cLtNgyZnC/0JVWCuXFi2ER5sXC1
hOGAKSLyV4c2i+y/7yutMBT1cQJkXqFkwbzchFR57iMurNL6nrPKV6O/RYtVg6WX4tSGcQ0/4usk
xaDev5j9dVPW90a6PXuUeegQnRw3ZqKDVkrEc3f5qM6rHNOJYLz4CZGB3jxJN+ZsSF7xQie8aIIA
cQoh5X6xbhi5C6L24RwOsvzj5Z72+nstpNGwzESir67hVJZsjk9cm4U/JJom9nwfsR8ruyH2ljq0
BdD0ZA/u88gGw/DWhcsfkayuA5GugvHi7fcM++7Z2qApeamjaFP/o2/Yf/YUaJ8g3hPdXHEExzAz
mSUsvMqXfwftN7IOtnjC8dn8TGay2ydFqtUywiflELi1uGCK8yI199CcSa5vkDqg6qt0ev7xJOJc
FWiKkU/V/Z46uBTxUAE+8mfxrlhcnfEQ3chAnMCJaSSSdOOODkwlMCgQkILBxHQFt0IdPK397RFc
hQmE3I6Q+j1WjGXUhOj+OUm/tNFM65D55uef6FhDXXl2rL1Gj8SJ5jPNuykY3lKJKlC4Pop0HPE8
+UXqOMWzzHMeis8u07NLhstwPwNcV1nExCdWwOyUfXZcd1bxyzT68GzCxOnbARQ7mx/BaDP03hXP
HbYtYmzuYEo1jio/aWj8tB5cqfZFJjUmE2i4hRO/EYvo4KyE8CM5LBHb5TYDrCuzqeEYmeT9y9SD
JQtB5lJpy/o/jhe/pikP8QSMD+fEJhzCp3XlVS1qeKHOeKWAQzu3GtaOAndxNgivnqWwfhS3uJdJ
8ZpnX5FT/Z2JoGNNt2PAmvDjv8Z0zF9sWldfhSYC/1s8/RMTMMkqP2LmsL3vMT6/MOD4tmz9MpTR
bFzbcxQluORcHKGPVyjlapg0+T2X5b2XDmGAl5e1s6/vVcDhwW5TvTzCiWnIotobB124kDythd4z
ArEUvz98JzCQA9QF800psXQ3AQVkmWWbat7oqKsbHN4/FQcmiRVEXKw2vi/ZjlQ8XV8KS9Tq5F0G
+ZDdCCcp9bgVO7cpPo5lPJoBCjSVEWfoMtyhreB1+v/24y+xvBmt4W/3Iu/FO9rHgNFObCHeca/o
N/Rlo+r34w36nCtdhCZV3rsDDwFCj0d6BeDeHYbrtZMa4gPC9Rti5jnCzi0wB1mF5mTQa4u5FCrZ
PNM17hNQc9SG7qBaxSbwhhAVq34BL1+7JIHD20bCXt4FxBhAoPgPpAO4h6hRCayMeBPXU+p6C5VZ
+P/uMgs5GyzU2NY38Cu62HzJeOP5izMtEh9fW7FydkVuwE5Kdhcu6GlVJytXJab0mJIqzMy3h6od
JZ/6u5NxbCPHua2LRMUYgfppWv/SkCdVMKvr5D1tPZzwsNZ6V1jULxnUkhgtQU1HRHi4TMur+JXJ
HzSxewum3aJn/y3Vd2s6kYWz5iKqw/cNWG57qb1ek0EyNUx/M92y27HjAV/JKDYvRbY8CNHKJaDP
+q+I2/7PQc5URy0IaeJM2J0+R5k4aOqzgAwZ1MsnCgNaG5HRfrQok8tLnwOx+THg40Q2DTdRPs8o
wFnggm0sJHjN0Lg9D5EgssAI1iz/wwrzOHKMYFpAXmIY1Cvrz9ZnB9o4tvz8BsOzYreypPWnDLSR
YBlc/5CljztQ55IruEWqEXlLUxaVt1bhADn8W7k3uiGB84UeOBQ7WtH+UZxjMtsDbnod1ktVsQC0
C8ZmHXFIuwk0NMMecYH/PXUNSUctMmEMP87O5KHCeKynNIju5xfemLlwC3Im2YMZ8obwpYIccqVE
l5/DM4lEo+/9VNBPor2y8DbjAjU/nbPzM4El2JBzKnEKV8s4g9OOmXcKiZWGzKOOirNF7BVN6SE2
Cier5oVJ9K1G4iBLyyE9UjEm2dIjK4a/3Jkauf1TAR8LFGIPhtvtsW6NYXDVEocwtSLE+bFcfaeW
tF2Zu6QXWAPmzxZONMRZLPT1OVttYpKnXcwAETR+ojSLI+hBH5/5CbOJgesu9yluc3CSHsEwlc6c
WOEcgOFrqr6SuLsJS6dZ1Khm6sLLom4raC5BtKG252qM2l0x2Sy3AevS+2qWcP82ifITJEmv32Xl
32VYqT6E20FfWYix4vTs11TBJs+ugzseKlS/ILhgOGTkY/pQL/KgvghngMQhL0nq941vAy3IM54b
RkTSgHfzKoC/JcZe5C7K8pdtRaWJgNnjyTG8XOvv63LbAIczanHhNtfVqGtDNVDQIjVsFcO3f/Rd
si/AYDfqR5JOiJhTHYI10UwZ+vZFAFDrnoXG40XTdbQKJ8EMnrY80WniBz+fQeKdwYCAnrqTWQeK
FEdvLFW9qTCjiPocYpnv3Dqwgk/K6P+Mr/rBpGelw+/eIew1eEbzYke+Rzji6+y6L2xYGcMJ1UcX
zhZCCjHKQn+d7L7GqcN5UStLfkhYT/FvdVX4EBU152gfAk1nTcm9e5IwBYGobdUbcwrRZLB96OXq
8xAwuOE48tpqf5V1IYO3OJz6xxYEYXmjOJhxh2liHLmoUgoJP4aJjTaw3uTnqPLgcFMLmnXkCVsc
bnRIjeKVjq9stRiBTyyhCV4bG1FqygXJ0yiN3LIc+fdv4G+2+CxddkIZi71LF54Te9LAtaRkN7V0
3JN3LyfheGWq9CciQKzOZCZBUBKNwXoTvF1nTkaj/doonnysrtol3nJbyQOiZsAsor0SarWeQSjb
VDo7/5t4k7M2v22D4ItsPBdy76yQN0d4g2UKTcASTTFnsv7d/uEvHNC1q2WX+ot9BRA2ifqlN1XN
M60uerCLIm8gzqYaNcAG7o+sk3OWCHPuWdm4wa4dkCsjsjuGfldsBe8tFgwr/jFliiCZr73HjOhH
cPZWMEU7fN3/iWfzf7uMHa0bgXy2rxgAVQVIkTl+rYtQoqa0em6/sNhka2Z7ytheW/qw3gay0CRa
PisSj163si0RjCEszTdYq4bGCluua3A8B5Wp2t8o5BCJiFOM2gqBnvAv0f5ox7mZ6ZLdNeVKCRt6
GyqbaN99WB4V0bf9IEwHoV8TPrqalZ0fGxgr0Izf9qaNZfI8goLn3UFAEpg5grxzeePUo5B1uIOB
Q9tdm8D0XESYCTq92+F/8wEhNdQYINoDT77vSZPoiBiZl47FozvedyKhkIhjgilWMHtHpZ/ChmIP
ruUFOA+3lmMo6s57NJE+YOFacH2BkRFwRgYcO5H+96FXPUlf7oedqUc4YO2Q9DvcCjbmZdoSMtqZ
bHr88fgatL1NrD+3cjzt4fHtkxWlrpwjkgzY/rqniYfMOHE/A1dIukpMt/uUfs4L/vxW2Xxi2a3Y
0zZItV+ZYJ+pKFcFXd6/D54CuGY13i9VDEIkmIhbNOHmKgRqIf4grgg79yU09aYgQvsF/tZSQ3Ug
nGoN+4uCBwVp5heLWA2KKrT/CJrsHnmcrcx7dyrc1Nhsfmx5VaHD51emwmHC7Dns6TmnOf00GXhX
+HbZq65Ro8b5mKZFpKuXsfCenwAi1nufWqeVmGligkqTBY+//IA5F38znY01kE+wivgk2q4Yx4Z7
mXYXWg3/yrQRJ2NY11oumvs4Ur7QIUn2kN7qGtIBEXM8dT2DU6wwUbE5kAGzwLzHoSIHXhxzPogx
yzRUl2ia59DJ4TODh0s0s0vS3UtcAOMuRMKFLAvRLpQxGw030EYBHFlcLNF194wVZk4clIi+9tzD
LCuBNezQm0ip4HLLqp2LbAVX5Shl0dvMaEpXXmyxxgCdPCxlbyPcVFjfIA+LoKv+F/Eue0ZsJX0M
6TOvqNxOKqWxtzq2Tqcpv587omOGWx7br+ZMRYY80eQjQdWyaxUn5ENjQp6mcjbGDt0a0sVMbdOD
8iwiIn4lcgjTKm5jXdtxkO3RpXLC+Q7XafgBpDHIyw1DV5ZgteJnPHmljxVHrG8Pv9BIi68Gdt5U
YyUFOBhGsRgrpo4GyhocqU3MnVUO26/TRqmQTnWAT5xnE2rF1DqpokzCYdgLP7cfD/mJpa/TAuCh
vQeE6BUiJPikCCvpgLDXXEC+GRSnUmnOarhMg+asgCgsP7iaDSs5gW0GyCCsgPgUpeoDSi+UAUZd
vrHTAMsdhFl6lNuT4BxXUGuJ8k1VG0YknLB8rTSBLBdarlXnv8GqUheY2QvYuizMLF62OweNIKBn
3zWXwqLkpqR1PB5BKpvF57EMDYrqKvJaylBdZjyEm/j70WP/E3D5fcBZlOPPTXltvKNIigqu3TaV
xvLgj66Jx0jlZuRwQNvIuSIH+ugHvaMqd97nVnddNO6gYjp1RS/ru7zn+9jOBdNW0ZIWzEe2wkE2
SrKlwEu7PoR0h9SWE3RxvKueHCp3HiD5s2+SBFmrkU1qHJbMn2muQi88tMhtj12VaNOkaSjabe4C
9ZiV+UUmfvZ5BlTtHMiQMshhtCODNAjqImkgq2JW3jfosqM/dL9jxMiOMkE83SB6ZD5SZqFXyuKb
3bnOW+/nCeCcdK8sgx8wi1wZGcfSvLi0JT1xa3R3FIhGb72unE8nmKcdZkTLCuP/xnIn7yYmsGAk
zgnp90Nx7FGbYTeNaaV09rgvxfuI4BE6qXEIau/EeNxI2ty6MKL/Zc8BudJV696Si928JoUy7CqA
yG8ymaX86RYrB6YFb2/dLi5JhpzKJXq+76zNxv7W5lWdSWBkQmOaxK1tDKX/IxzZNPQGmar925Tl
BcvXBVcZEt3V3sOv0LbpLt74xDp+84nmFChwo88QKBzMKGbX6axAHY1WJfOvfHhpqFfNXraDnt0O
a3bYgoip93/zu9C1UXB3GgH6isDA+qrTUhb5R9ZJM2TzArXpaJF3joiPeiU8lgVudfEtuo7FnwnV
B2dzo3v5l6qZ1KHiv0EZYY2XqqcY5iZEFZY6d/AVw1ywYfLgzJsOUMS7obu6AvLtoYc74gNu1JTQ
RdLWB3TVZEv8mJB2nkuLhtdepQM1VAHK0vTDOVW+HTxFQCLE662ccNOnULSjXxk/94hLdtPNKzr0
TzyN/xNEwJ6QkRi4rzYDoAiR4Pt+N6AX5u9oNgi4L78bdXyJGXPp3OhAPAvmf+12fb+wiG0nj8OT
hBjG+zTqDTSoAzLavGcQIsKE2lsqgJfPKyieUhB0NEBepx/Z+UnfOmN606uUTgY7NyRyn6MwK32s
Bml3SmKs2xZgOwiJRVqFdEg92L3e/T8yz8hb51XiKqhiG5hPrnCgFszdGipcq5PmBJJIga/ymRB+
Jn1dKYFXDdkY3lwOpIS5hugIQnQcqyDSzXec8+5iA1/gfQRvvECt1cCx2hOledcIhtcSeTdEa7qP
LBCgn3AQFG3EB7xDzhzhsHB0duz7+G5N3+IFB+kCue+1YxVASJwNszLQKPi+u5/WHzuzd0wQYeyz
0oAsven1K16QSqAqtQp+/o4bf3hW9a3kuugXetv6ja0eQvVNLbXKp391xt4IjxtxhjQ/XqiQJsT5
ekkbxKMPE1MMeUYB54zJ1I1M72q9K9XYOYAWlIZ12zTKRMDh8sFOP88hNDZ+jmR18PTNW7QRQbNh
GKASm78MBLuD6nug8mbrfxposzqGwb8CR1xg3D2vPH6MGRNwzoFWeR2J1zFNWXV3WCiBlmixiMub
oww8U+3EGEbRWTaz7IdBo2FJNgP/Aq8NLdyUO3eJycPbrmTXA9K8JMn7OBvZmfhEfhAJzKAJeFy7
d/hlFIsjegZhrceZPxlPTi7/UMYAbv7PvXonSoOSDRblgYKecYE4/1fuHvbW5q66q1Pph0iEY6P+
on4hT7ObJlDyY1zVSc4W8Lt2IH6FWT0r/MVY76URbkGJ4041+YIdYT4ALc5v8rmizhDmCSqw/bSu
k1nI5I7IXwNAz6D+Cyg4yCg5aHayFRH2d+VMDX2EVN7TZoA3xu90lYGQmvZst/gS3KLKJWPivUrM
zIK4AZNFTDCwoofp8pEDk86VDZow5D8Un6JPqMJRjNv2J9RmQvZI7dss50JMZ2apYiwwWAtVgF0X
uxH98hrULVJVhUJkv/8VGys1qVbqG2nyajMMFEv+Uj13zKuHk+Qer1ixdUca94m+wqv4ZeC7yxal
toi0rJusmTT0qsk8yb9noGPfyIjfBz4lFpy+6p6f79eLM76owaoMWxgvJUk0/IfOrm9EscIrmyeJ
+RDCoMEOzXv91hcc6O6tK4V+dMnUy1yV1B3pAfUqMjmSnGo5PL/axuXyn2uxuKl2RIneeB+c/tg2
WLK5+Uz+g4c12V1BM0zdtvGiDMvQiC+dsdMk6bNgUBR9xtcxEa1S/zqynvPHdosYCkahwdfNKEsf
YDoN+lkpRiRxbxWgV09ELkRZu3PYkDNRp46OKwyvo2BxnDcKIZ7uK5m5PFUUQiDNylynpiFLH6Mo
WhKxrFi/j8J37ZKPAwtPz4iciGREKOV6REAscQVpf8Bil8opv6vBve8as9+xqHybx1GIkM7x7pCA
Gfk5UTUqGYCjcTcSN6C7+AfvhoNQCq/JXRxDVeI8s6cRNbhCXq+rnUSiLh84E0oJBp3iYjzQxKEc
/l2h1pZJtA4GEULeDP2aZDUbiZsUAhhxZzPSXRSzxkAJG5LaN/rnpXiY09lQBVWn9DdKd0mpCGvW
yVg51r5wRsmWKSEHvq16CyhmEEsNf5dPDnz2Gkg4RXs9AnUIOFwdlhRLRAxoqIwh0Y9Xt4GsrHti
oFiAvbJuXCtpqHyh+O+TUGoZ+3lWFZ7SjlYdY2+6Jny2uVm4yDyI73kJGgmwITYFwuLgsHkdhZ05
Nx6wFsnytHoDXQ6qg/SUf0wB749Qujl3Ncv8KUQas3/KxysOlRuE4yrMbACia2Qnmijz9abQErGt
QA11d3bD+in6RJ/+IyEKj3l80IGNuwXGsMPEOg8I21POid3l5QM4B+Kf2c1G/NnJ74dnRrBKDX81
YlAy/xDY0GelZ5yGjKNRETQ8cKJM1tjQishHfBG4JNnr5UWLTU8NuzGLJooK/1VB6TCkwTouKzei
DfR1C8T7EVin2/ViM1VPPAL2p2FT7nfkJEn9NwPsz1WBhfndjJTKYQZcBpSvqJo87BC3tJnV/JLD
blYc1OHf1pnczOboxb1AhMDlJM5S9yV+cdQq+lgxIUJN4v5DRI//wzozxal7aqhgjWBCM/u0kPlY
Ew/57rd2ROpQsmXs/V9J6qnQrOnfJ1i6IDTni5BRVIQLvWGmvWQUH31v+EbZEFnPSyDyhRzTHE0A
bRWLoiWK1uskwypbwbAEExhlbVPif/a8/A+rodrk6e0RAhcdKIddR2bLPsfIfIKdAwEQfNl36ijw
v3rae8fPAiWPyzOHEz56x55M3Va/fuhlfx8veEXmbyJCC+cKd7Y5A71sguxNhYaBGq6jOXxq77yz
Kd48FIkTdOmhf4mUY+DoeLYvCkeo9ou4bkikTJgGTU9gSbcVzqvOLSR6AZ6kBPZsCNrbwW1n+UWq
bxbqt+6FExTQOWfdU73xNDhh1COGQD6FT2bjfc9+F2dyTEkkdmE+kfbkiAAecNvD+BKrSAE9Ga6N
EwiVWZ8Cxeoao/xavfhQrLhb1sahduZEo6fP6qkrCRyJktwlnL3rf61mSRwnSGLvKJHIYLGT4m2b
BDjRp8agWoSiDVc9Qc1Fj3N8sFutAXeTWrKzyVBlUTGALUcAU9cUiZ/SBCYQmPj3XIxl+9QmYcQf
gz5oKUEbAmWDfLDvKfyVmTER3maTHtz6KK/oVeFYMQkXzIKubMCq9TD94CUIe5zykFJOI43DISOG
bgQL5Kul1apsJ7jUtrJeWHIm6EBncKLNXdzIaY37phsTvCUWQsVwpBi7NZGz62PzTDLUtnPBnedl
iL41XOqrEReIzkn7Yb79DhVIe3OFTkv+INRiPLnahimYQxAa38aYgYV5x7+VJyapSKwabNlu0HNG
QWpbmyZd7UqRA9/I42JhgKanPkTMJpJ5AtOYIul2/iz5lrSSuiI0HuKCoKFA86s+LtVxtcuwEm2k
lFAYxWRE5rydh0MuMoaPkWkjYYhLZw1jF8K3EpbWjXQMe9M4EK8S9Bm0myRqKWp9IQ8rtbZIyyb4
ca16O8cTaTolJh73EMQ2Ugs7OYxkZ8kIx8mYZGBykCJx/pcN2EBrs3mLEvs/VViPbO/JO7tM7pPw
FBPLqSEsmE37i5cQyEsYsKg/2r9j14C/kg/RE8DT6Z0E272A93OgmDp6j7h8Kdugrg72MzBfme9q
f1fL9JO7FLYelhb6fNaZfkk8pZPAw13qucA37+Zq/fQYqdQvriGxsUDOrBqZ42Sv/3fRZOWk6V95
IU9F3Ba/ZRTKp3nj3dCA7aDd9tfIT4oUEilp5Kef+/ag0YA426+eU8j+RNSx0/ZosF5HyDORuZRs
cKFeOnWRpmUIbdFn+0gyp2xN/eIAeWwW094u63axVXFfpxmzwcWLQlZzbhXvyEAvyjhsFmEfK92c
q/KaGX9g7eqXyP+UTF6Hv/3cUEP0XwywibUlbcdgrSHECLrhScADb3L6944H+zqmS3D3JsGJPI2Q
Pf9I5K4VdJECtc+yqdbIqK5RaDx9Hxm4y0EvOC5cFuDd6+ETFhOQNMR/tm/zbju2Xh7P9NKscTFX
Ci0UeLGKxEV6Ga1j+yEAbhseSTw/56Tn2ic3sKAr+IFEHOyK8fHXI/RPJgOQ5nSoN9tFUzw4wxoL
In0zpCaFEeO9rZpUtg7qV12eT/lxZ/8Oi2Yv23Isw1WCGjokq/wfNPY6ZFZ9Qz+jHH4+k3QMD9QX
OA2IP+8O/HhEohpLuThfJLj4tLN+E72p+nTZktiYPLnuh3wndvGTUQZVZBVL8yH6cuUSqHUIuZTU
N6CaUOwjkI81Bk6ZQbP1N2PntOMUegJvc+kdxPDIpMj7qOTt1TMb5Pdavi0YEXroqsH/hlMU+bx1
8hWCPfVtpy2j4IJ94Qnfbq+jikGrqB9YVp/d+aXRfi+3ghCJgYF/hdnddxB4taopFbZtpzlcmIO+
CfANtCm/puxJGlQZ+rbR64qOHUalcsUfJS5ln2VD1TyAmILzvx8ueHLHMaGGdVCWTrZNoN9eshYF
a2H2jWAopA67ZhTY6kFrh0kpxjBzVG3K6uaUCWA8dT1ytHtMwERBZ6pqR6Jpu0Y4uY4fyF6D8oaU
CeQ7evKLR6WYJqxbHxLESs98iQXZHSvmJ/TGVKIqZW8X9V2Nvu7EQ2E2yT2/k6WrgcyEybDO1DK4
IxJHkeuauqZF1NSkV3bct0QzDdIPd6DGgxuYWycku+MNZaWWlyR0lnI/0Q6RmYJ49nCHvBabuFBV
daeiqCHl8ZkJcSOQXfPzz77+rJQ1/Lduo+fgc8SBTY1kVk0EUtRDfp7omVo5+ctAPnzlA1FoRkkl
uCylYYTbqBTfTr9xZnsAH67uFDa6HeFyvMUXjuvcBZgH7rqU977CWymrcNBMepjh/0H10q9o8bNS
C2QuFWfcsEX7NT1+0Dr0fYUE7uqIX9ukzMBUkovtDfpJSpKjfLM5IrU8eC2/GvgNQQEpJ1AydcLx
hjTw5iJMY4USj7Oa2cXCQyicKGen3kGoFwcA1k90iLCd9iy7GEA8BRgfMYciXJIoR+A3YTr/6Jf2
KdBRQeQs3TfyNcMYuzIKBXKGZGVKc7eFk8rf5SztFDzel6UqyEwf3WwgTiktvJxrPhUkZS05OtBJ
hwj9XJSb9nQJ6MHoaeqslzgp9q9anlfMh20N9sA5tekWaLyChVcQLJ7w9RW0Bn22dw69RwIN/yXe
9u83F6bLqi8RCP7I28Edbl5ptRRZzPaI+NhGkmrehAZDCvuLrnAoGKe+MsK8YMw2wj4bgy4Jbiyv
VmkQv/xLnDGzPGJWQwambX/xaNcxOFmlMWyW+P9hpUHEbz1CalXkNx1jFPLkySoj04eCOj+I4mU5
esFeHI7JLbyfttqNAEUwm7dQuslgyXWpfgY10yTRpeDsDtzMYA5tnkhofKWSmffM6cM82xUnZBaC
VR6EP0cuVBfHTkBEBKU24EAaFfI3isGPmmVuIhs0FIONsrU+Vv+NFaFmylLRsz2RMzThdKtwfMox
mcktQjUOU2cpOoc8MvKt6zJvLvNNsFB+dSf4QE7goaEYIf3Cvz4RTcU6uRXBn/jP5vc7GdhvtJfL
++9eorC3UsvyoPpO3RtqdCT9qw0ptnBREA4P7b2X4pE9cSh9JFWPgXrlgQAnahJwhHxf25cOQBzZ
yhrBvVp2tL2nJ8vIaX68NwQOmpnAV3+BUjxemW67lTcPK6/WmETad9/ne6dmPtusbnrt3dAv0QsO
6OZR4vM0KLRRbxzXR2Unl9ZleGz2mj6iyr1a4ms2r2qK1Tar9JylnwKJjFRL0zj5gh90TeKsLXjl
QzchFKjSmIJ+yvo8lJTO/1aM5J+nSobqdMC3kGCofZRMV2xdMfvVRuXYLq6dVPV5J0VkL+eJ/bG0
9j4j6vWEz4PCFifzB9XPfyXyAKs3ec4Av7vNcvJODDIVS6HkQrckSQYZK8vp8PIg0hHDbAE8Iasd
d5VRRGFMNyZnkYrm4gD/KdbdOACwj8oXwxR44Bw7rcVOSpZl3bt/I2mlKCJC9Hh+PTCQRNfx+XGT
3sWZ6EBsCJusxCqZigbbpfGMH0StNOfiVLUmZAn9CRt0Uwdav1F5f5Zp4zNovW8+rBSG7dGiJvWh
LuBX6wz57xLXADgZb8zf0ZlLe+j61kIKH8JIf7OWYJ69GgLN6yhIhhgjEo300Fb1J7EngPQruqlQ
mOr9KXEsf5rFPmK3zmyzk5u/QhFaUPOkK3dnjK2tClegFr6yEfMCjGb0e7sOyJR9lAdklVZg8J13
Fgl/XkfJ6lpEEzgvmjO5Yij9Paat0vfwG2UXqGzuag524ddECm62Qjm0Uab+C78LSMxOb5c5dPTI
83/cgGQLz7vXbGQHiRy0l5A3VTNZhx1sYweK2vIPYx2xGD/O34a7wc2Da7lP365iQ9D+zQmiydAQ
DIFogqDmas7iW8R3+mmAbEuKaLA1ALRw13JUSkep/M9udIb54FbVmcNY3gXfKB05pxW7VgKnGSz+
8Uu8+89YKTI9mc0BnUNCmDEEV9qK+5Tvq1JBTCuJhP7vPaEohCwaAwpmIGecqJyP1XLVuci8Z7As
atgfc9dM7IW18WdtvLzbT2Lv2QNdKLty9NmIcjOViwHgJmfFqMXEgxUuAmomCHto6zwVRIAkuNCu
U7rIixXqo7yEl3yLGfJLt9bW/24kIKij7Rm6QLV5Go5veG5vAOTBXaCPOj91rfZRMd2aG6R8B18j
GsXCKsIAG7UWiflzlfUirHpMye81w45dEEKahVUATXr2nfoRZcxw9Y8zzYngzjexh6FUClcHDca4
Ep66TzOJYit6JvA7RHpLa180eDVNOLgbI49PeGCe60IeClZegyQp+KMW25QsGdfP14cpSZa7/vzk
Hf3Nslabk2vGFGzUw6BkGh1Z+M8N9k+FnQFQONm70jb/n9LHLKmRPjms6MVO0QwywBf9MP5akf37
T3uQD4dIqXQdjRoxhgXyX1q5ZJenjHAzH0FidF+pE/odNnJ/QaU/5+f34uJvTeljR9iyfarLBeDO
DWFgS2UIejmWNQt7HI2GbpdJOcTxfZfMjU97gs8XcF0PqrEKfACy08rMUEEkfshm76bm7Oqb9wLF
GI1i/lGnwTCubr7VcgoWCuaFoIkwYqehB8oVY5cK1RXTj6VDUSSz/nIMLypSG149jFO26KVqfNoy
1lzwTqRTxp45rqK9I3kxMegVbqtGtGhIeMgO/q4Sww+ABwbQFR9vt4B6g58l79I0Z0Ejen959nEG
gqXN8i2yTlfLKqg2jXytNkjk8GbQYUAQK99YxEBLcEH2zMTBpaxmWnbsIsQSuEJM/7qH8oxc9xIO
lVWSh9UOQl6UMlEnmigQKcjLIEi96WglUwCqLt6QBvi+4Isk7Fw4gpqgvPkwJRfmhfKitmuWSHvU
hh0rg8wevAPBwQkAJUCGTQ2jpZ336XrjIxMOUw7vF5NjB/Dls+2Vn8y/mhYArl5/6/89A7y8scg3
vUgsqdW4iBIr1Rt7XUP3SGHCuK/YEI9p5x/m9AWfSvjuVnhyMriR1Jy4WdlP3k83AqvQVT6G3uAJ
dlu6bmahQg0RpUVdHyrSC6hW8NNPrYEKDc9UVmrvBnHdn0QALJ8Mqxnjv/JrFbzm6k+DLSz+afMm
WYGhUghtzcv4nyPAiAZ0xo37bXcrxlVd03UpCS68a77JutOexiXNU8KiEA0i7/X+o7vUqS6nb24H
Fte5MuRBT0ElmiJS8SuI1hQOQicSgKBebZ/QTQanP+16Rv2lDkhdl7EOBUTopp887IXj8kw8qQR9
D56RobkRGE3Szvfbg1zXthOqMhlMshLQQlK+SRuH8kEgsQOKlFTPvchqP1OpJwuDg4I1Z1S+ueJc
GOX+6H3QDJpcrYmZHo3H750Ngd6ZSsnY6ivUtB0zX33hWBWeR5WBiwZrH39zGmBxtq4x4USs5Zc1
yMs3d8tuvwx/CTIkitC4ICZhMDPlegnI2GO11Y3gMxaq/QW8G89aEV7ii0uv0q/X9m3mUPNTzPmr
6lrqUHvhdljXkkeje0FQxeuaImCFBP6Btz0WqpTYEzXWcIx23A4qtZ63aHk7UA4B9/aYX5BDUp+n
gVjY8KKoTUAmozrcaMEWPX+bE2ARAb1XTP6EOmsC6tJZFWZOtCWQBL5JiBNK07yYTpLty3QRyiTY
blcseKkQEeGnz+tPMo71T5X/SPnW+pTvjrt4Ip/HxxFET7TQAZGAzt7TelGSXwtX+MEtY+Z1mStc
gONbCRQUPwXykdMJEvufTbaO8S/fCfLkWvG/NIZ4/1Kl4loSq3J4Ze62yRvm6VfW8lDcUZVCZnve
VfIlYvxzoiWlvbQdWBC0mioBJOBnEjDQbW3hSlvYoZbafVpl1v9H1EPCFfdd4mehANcn1q9zLXg1
XdmoXPqF2pk/JXAGO/lUHzBIrnPuvGhnaWGPd8X8PRndDwUgwaGb1po1epR+I7EYui9yoMOrZXtG
aqtVNM7Xq0mjr4ldCLdLam/Xv69Efq93F226lHciria5viN8IZ3u77M4kSYlMrR/taV7HsbOVmI2
Kv7IkRH+PVAx29rhGuxXx/q/rBiywyL0CW/uu/XYl9dcnQLrFGLd2yxL7oYgtesPEYly5MHhYIpu
0FB65oeCqC6C249Uu5EwbMDxgcXmnEirA4QFA+szabwtNBux3Xq1l/xpBGnmTjTaV5dla/Q789MW
+pv3J86sjPJ+X2P3Nx/Zq/sjZlmS2CANg2F6ucFufqBWrMlG0GaOeWLsjRO4VupDNOw4orwS3ecw
hvfy07ppdZsPu6+Qt1zRdFhpCgIUS8MJAt8Pm85fXvHzqRIerggtgpQJTYrYlIUGLOautx0e2TUg
0qozhjcPmpF17TFa91heRNl+x9ogbZYYaBevvVu01XwrGY1KkrgtLElZC4l/jZgn97aLzj8LrkLb
CX8BG/Gy//bNP9Y9JLaPU0jR464WxW7Ys4eO+/gqWq7jVmtX2FDWTtovtp+zWR5eQ69rSs4AN57B
brI7ZmFQzyP3+MWa9ntiuBZWuxmJX4IqXUYrfcIul+VuCQnvgJchy5qw1BefnnfpL0BKB/d87FO5
OcjnKg2H4EPWm1ccxmDwX/BEoR/+6L9EfEs49F86YmwPJTOduar5hP5NgYG7kN9xScDqt2J4wg3m
7QgMZ/R6wDwxqAMfRp6F2wOMxilwBUjI6+oy9y7LXLIoZVfcfpqtyJ4Bq8AYxwNaevjUZNrQtvZp
NqAqhN93I+ycydhmlGxanXdujr/Y8VRbIgKrz5RGPIyvO2i3btUwY+xRb/jSY1hXavLXRo7D+Pk9
jLWX7BJQ8MHea9nuzc8+r8Ki8K9Y1K9GYVyuCTm/m2g2cgp0RoC12KSLdqwTIizmePNI5rNBl9Gj
puZqoGkFw2o+NHr71MaR0FxfTIFaVST8YZNIJdG7j6ZSFGcoGzgY0AHYGI815Akk87RK2kLL/6h7
dbhpX6gIJIc2Zod9bM+t+KqwDZG9N+9RFtrVTOoODDATbQZWvsxG7zqV5Co4FT7n1MOnf23ZyWjb
30wFQZgZNohDA9jIMK2rZUJ4+Ryt23IiiAlgmKJpghkjBq3V+FL11vZ5cgEo2xQPuGfcDj0J/31q
2oV2IQeh89T8fMdH7an/9WRq0dGp0dmOU3r3AW38GIlCbnGXdKaLfTnMUbmyvc5UvnOaqC0/ta+p
3WO9yyGXswlzgZXGLa8g49bl1AGtxBNcxVyjckuUjZnSSPxbvbnbQFu4y9g+K7fvVLm4SQexNS9O
VZh0C02u3/Cxrcxe4a5NcK/H2tPkSa57o5loxn/Qba2YRR5SjAV0y5poCIX0xzrWqLJ6cmfj15Fh
kEEt3b3MKMIyoznEKSsSDNsZ6uglsAM4xq+24J8Iouwwn64LVLIB1bcbgJfLXE2zq7XmcDAlWvvf
+FBUlXi4yHgcmpfF+8OrHe6y/Uw4AzCnByDW5J16ZunJkUG49QsanvNaXomjVKOIv3/9KVpgEKca
mFGt19XUQD6xK8ivZ6nYjtbss796k4pMgLdSjBGHhYBykFd+o22Wm/rO1xV+3yvCNVgao3GKldM2
9xoM8YfRAbikaNcQbYidkrSxQj8OqDY+Eevl59fUDh86Ys5X/anYTU7fFkJus2hh4mIyUZQEaFIs
I/VH1415XOKCNk0V6M3LtZy3Nsert7rYMyVXAkRbvJUrEMzKhjn1w4bGxBVlG24PGpDujMt3NohP
5Sl+u0CMK32eF0qcrK2daIYGJpm6AybsUa54qX6QqNgaF54JSkU6CntGwxSVPUbI4xJ+2CQV/6x4
6NRcZChtWeU52SJkiQ/F0HoJuw8tRgvyqqAh6Lo3HwemeR6J0EyqjZHynI67lXLsOmtQvWUDcwki
mhNkRAIIEfkPpaPHoQFDY4qM3/0G/OMsduL/pOkKVaT332QQVzfoIo0HDp4C8J4PcSVQBjo8Zv7b
7QhzW+Pe6RvftJmFqnEbw7ZLhlnxf+PF3kd4RMxTQdXjRDBT+3as7A+sQn89jp40JJmsD9zdYB2+
dg7bErVoOyNyT9LUWaP1PTK3DbwwKlFt9mTtD22a6Y64LB/3p8FJE3nMSrvnm7H3tqhATjowoqPU
uMKjq2seyOOdwY1vKqXylfCoqfjC8i6ZPupZSZgMgrDGINBx6rMif+oDR/sOqfwyK25HeYRsXggH
Z6ZIJ46LhCsoOpQ0B3J3BI4gPGbPZelKVfo+BhRjbEbmqUWZRXZXxKYROkFkhF9p/4JbrxaXzW/B
V0TUenXqNjw06banSr45Vgu60337mmCTgE8TkfQD+SSFE1G9hnN5pA4B5cPRLDOTcDsXQsm2DB9X
QrOhoxEgtajEAcKbBaQd7X3eZKpOu0PEey8pOyaVTDS4mghpaV5S/jXYkXc6cFIRAvim3pObfGQ1
ID/nUlYgQnMj4ChQ3IptaQlw0q6UyjZzjttwbMBqLXTCHcInirDSlnLzWiBBK+KJxxJ0u2h+5J7x
znHJw/0dcreuhQIXKu0Tm21nA0pSKD4wEyxlfxhzQKOUSga2bHSNLbwoSocKsNNdrzdS994sKpuU
8pC4y7x2fTFDaoFXMQj6xxNMQKXItgV6+BeaC8vDR3XsNmI8C+yWQy0Z+3TyMJ0gQdA0es2rhG+L
Z91dnJtuY8R/fwa4M0Sf5ij/DhBOBhprnrdVRj5ozxPccAmeCJFSA6AxODZjMR4cgNHg6JN/9Zj/
VCKM6EVxZG7BeAT/vr+dD7x9d3a4w0VsmAkWvrY5erzLr9XBPd8kOScRg1Vju/fnuuGg0dPbrvBr
L4/XI0wu4r7ctMJCPrtSxYPS+O6R32bLtp/4c/jY5IPrBxJUdz4swiuTnvnHb/z4CI/JcV9WaFWa
izupFpaggXEctiZ6lzyQ8CmwwYR8rlDT6Sd00ps4qhK2/Mu6cQVcoPbUSJjm7KVhcG+I3h/7Rbpl
HKbpidi/ICtDSk4WNBqILWEo5hFnTZ1B0i0OkQBknIyjVwxExq7J6HtKtF0mZLVQ1m03b2Klz0cc
gnL0SfMvBKKHEuFPIiKgim8Q7OCcJSm5WWh6CYPvqhd4ppUCHB23PoGGUy9IRCfm1l8lmwn2+6JD
i7UjMWQ7pJUmdF7VWWGDwZVrdB07XYRkhB40ygcKuzlvH3bowbWrevBTmBwn8fiydR4W6au+GFC7
FX6QO7gVfJplq8KuiuTClMSn6ig1haT0FpeVAWAIMVqMLHqDGnNl4WQZyl46sLA8YYb7xzHLYIpJ
4Jr2+6+HnEroCDJAp5x7x8A0wgUXZ5YIc8jwjNxwAIuEweCGq58D0NeuK3wiE2abaYHuH5BuueHq
M0/LR/RHC/fM2ayuUFo3uktybpisZh/KgBW2EdZxEn/lsrhbXR66Te1Il3A4fPgECgu1UkRexnVZ
a3raj6QL7VtKF1RLYnTJI55zRsYzu3uKCUzDZDD0Icj3hLfLtEah79J42Z8rh42i5fEibsYE3R6t
yNmCvyeouUe8JxTHGaMt93A1aCS/dQjeMP9bSKuyoj5wg9EGdC3l8AbqIVO+C4MVwTbQrqRD/AdR
KSslhbB0az4oEVt5abwalMCW5vZlb7KM04ENxmtWjo0QTYBoRIWtPfm+bx8QgN4Ih+9EKYcPe7h9
xXRoNAhDaKELL3Qx+Ddb3oNqjKcfaHOAFX94hrU1i2bYj/M6XggrfHKgDm4QTncDFoEEPpI1DL9x
vnlgyqnEZdtZ/dHZsDY1ddqWojh+T6llYmfeYfN40KgNY2IfO2HfCFJMhhCqBFqcbuE+hr/iA3Z5
nnnTzvmOqkql2zbO7xst/P4P0hPugTEpI05ixg7VD//szGu63yRLIGCpTx9BudMKVMpLVo73p78r
PGDStHhrBx2wNPymYAn4S99xdBh7CfBsL0ofYXnzqY4QPq74tAoZGu+47lMyslCRtXwhJ5SIOsYX
vpGzwNRQnKQcI+fFTuUpk1Q7CzV9xvCb/4LnPXjeknf5k4D6FMaWYkwo18RbU+p5l51dCFJzbcwg
2eZWsfEFgfs1uFQJ+ZkAsguR96lbSpOadS9niL35tLeBZcT6DYHWXGRKxt9SdZpxtJWjuxUu3XIS
/wPD/7wDZBuiKKz+10a4fQr4oEzywoMju/FOqlxT2/dwvQmCmyxaoLkHCn4pkW44NcAzymEK7DFG
KqWNtLoyhL74BR2LhaPqPyqqlHtLSaMC2IeKxLk1KHu+T+lVz+m6c8rOajoNYFr1vFfgpFMxwowx
TG0bLkn94G4jmLowpB61TOGWzSAiZUrGqQv+7t8l1UyStrRur6MxTKxNIs4i/1ivDjJXUzdEgi4e
JUOqfwpqs6YGExNES/COMwGiRzZ/hQD0dcAJWQHVemdEZSv9cu+tt3bfe95LeElzc8vzLeV9gfZ+
32V8wARWeZcAA0zEnox3pI/3ZAJX/Y8CDA+KI5ZdWaqFrnf1huXwqw7r9UxgxBspqCcsnPihF216
UcADikrHV+/5vllz36BKlDr5JM6ivdxCxgv623rQeq24vD2LfWXkW0xUV8P98W64zEx436gfTCGX
zKRVh9aSnfzIsTbhFlGd5yROneBVOxMTFMv+gg7AmTgcbOKst0OHlAnBdFPFdo5sQTzkYXI3qrHD
OIUVOZi5O4/D20OorTbjDeJ3scacT7Rg8EFanlLquOyq2iaOnKy14Xht7OXwq3CRSlvfLpqaWBIw
dslTvsaizljK67fSFrmOX0lH7xcNU+2qzTBKdp3PlhejfotesGKDzQU/7mtDbBtd4ajvlCyNs5KO
ztUSQ5St6OLrZAoejTqnxGZ44on10FgRws2Mkuleq13TAwNvTdod1lAhbUUa3HwZnDrbztm+O6yT
mPvHLte9DWuroiRalo6jbvKoYXXn/dNPIuIfNsiD63ieWosQHWzzTtzQsbysMyZrJnl/2t01MqtM
zsfPxYsNSz+sjPsYH2SbsoqqChUQCZ34DOh1awSmO2QjY2Tk0dIi9kGlTbSBX+QLnin4DDurEHtQ
GW3FW5/PWC5kNFNOlhIOiLrEZYsE2Uybe0LUB0qxxWym3EDE2qjZvPLFGHMSHrorcLFJPWTQI7K3
hFb6PR9s+afqnXDJTsW0hoJUwvVVjseMxv/gTrxhPIojz/ZzQBGRJkbrmAp2eo4Hig9dw/9E9TZR
QZKp1/I4Ce+laIuBwKur62J759j2fR66lFvUHlgwWa5iFsBBqQw2QzZ1wvho8lkThbQV2ysSLBHK
8NfU4gu8bSk4bQNRD9Vy55TBu3Z9NtZA/YI6UaD6Wqj8Kf3dcaJvkuf301OTYB0QKeS6OCT3pPkJ
sbqyPG6xODEgz3V2+EFNeB2g9yXn9scwVTbiCKFRqPQcOTTY6P/1wqypiSC7XzBpThNozNVE2ijX
954DhLgA8GCF0Qn74cjc9O5ICtkL5zlzIPPeafR8S50twvqa5R6pUN3kX7/poLIm5hbyeajlApWo
QPgGsC9u8yxOfibDY/gPS3BdfkzgOgQdBvQmpy6MfAslEO4Ac7mWAFKiVBz2e8mp1QBjHML7FAXz
QRnWKdndqFg2cFxTzfR3jlyXarmmxtczuIQmpyKymxquM5Sfqy2QmmWFDt9DrtXdymvaJirHMQ6k
yxm9+UpKGBBIH2sdwQnCd7PoekGEWpVeHp790InLw20kctOsEIEg7pn9wq6KjfTiQ8dlLH2ymetL
2UlJWAE9i7cG7dO0F54t9IqxRgMyLJRquJw4MmCBlhYctATGaAr4BFU8uwllTMzl89ArccAumNSZ
TmL8LCfPGkaIKcVC5puIJErOdyWsl4W+6NVzz/ZOIgA2T6X5w5SgUf52Z7bcEFmnQjjNasADmKtg
JYWTLJXH9j3QWMqiG4rfGIA4CRfNj0S7Mcpn6ricEEADkYHpgmk57bYWu6haUhjQg4wG3ifiuqVh
qObMm6sDn5LeQnhron9FhwVMPX1csnJRLEqwga2+LVsU6gKKba8ivaVuqKDsh80RqINHqfhItHas
gKxbN3SeDd8QfGp3eqCseLFj3lQUMNbFQsgfpwOJGWTnuLY9SbRVP8F2011R/2CCBmKP9voVvlEh
2ILr5JYyaFcE5VNjqqs/iqrwJoGPaOIZrD65YkiJfsWnW1d39SnCf9sjdgoaFLMSCRj/ZQC0PtX5
qqAC6PCx9pPFf0wGhdRRw5YYidEK/9XlmH54WDgd25mU2H3AmpOEMukre81Q3qrXoPVltFtapcTr
CkXxp6EpuEvH1Q9AyqyflZ5R9FmQutYRe+QnlvgZOAosN/RpKXsXK8nMyC2ooJdv9HheX59uvGVQ
HmRaLPhnAPzW8gcaYLGx5bFNw8MFdcGvjND7cFnwnSw2so6X8ipDdvfoLLBnW3RWzDxwF4l1SGm0
M3e8zuFz589fDBDVfq4AsLYfh7AwGqq1hI72zpGTEX0eF2eBmnfJ2ssq45l2uebZtyb48h2fg0kk
df5VcmKig7AN1knMX+kcfdaf3cNIocbxSeHp3y7puSYARiJJh34J54iCAgsVGxvczNU18NmpM7ez
iNVewqebX7QZZ4JtmGL25HTUQhDxFGlZjojMhLsLmLvnoT4HdfQiFYIe7X7reYUPqWUg5Oj2gU2q
7+VArwP+NZrcVvkdZslHCmJUdfDoDowe3q0RF4E3wFzknT0Z9TNeWD4362pP8WyuHi2n1qruauJK
fSgtNV43vQeb72xlFYZcnnEjKe3qg3Hr0BMk8/3mlZc8QUEY1BgKPfV+Qu6aPM8I3qweJMlYvzQm
Ma4dubZrxHUott38Q3kwEafojzR6LLjP0OFFEaUOCJv8x4/i8GPHW0Fpj2+xm0Vs2RPjkW+uOUaL
uIHd+jenMIT4okHqtg2RFmSeDv93kAoslcdX/Co1xv3T1oeLNEDhxJ7POURbLPKh+MaKO60zr1rV
gPmnjTxigI88+AqpwGLMjcK3+EZ0yYx9ilEsywzxKET0jOg91B7FOCyOuwRxIYSUOMNnyuOhpA1B
VgzBZCOr4QCPLe2jzY3ZKi6+XRUXtg3q3ktdiQke2YsGa3rDsG9fy5prRgBxSxt1xUe75phE5i6m
RVkGkqWYDiAF6KmV28t3iDaGb1sTIinsxDBON0ngbmERffv3tt3oxfarGy00IFSiEEfuZcph2c4h
XTddLXyK3KL4QgtyNXKlqcrsH0qqJiCmpThu0JlUkDU8zFwReCgAhCc46HAqsgBgYuPqKKIbk8Ol
Tz4ZXuem7gFLAFZow0bUB9PwZonN0iWi2lp09vNTvojX03SxI4e1MQj/R/bKIPMTVNiaaDUQsycy
z72kuSNcKHD+hsa1dhuErX62Ll0pa9fhfZmetm/fST5oam4G6sQ/reMeVQjSWFVMa3e/e5ubWo0j
H99cFT/kkfwXvHQ59iSCJ6Xfq/63yN+ZhN5ymYTCA2RRTsUZtBTxXZhDMH4tiMvfl6TGpVAazCsn
9z+OLz3LZRImp7a8STRG/pF0ObQVzXYMAb3slJMSictqGLdGYYwDh+XwSsLpplAkR0qvjLMscU0j
kJ6SIlVJX/vQQOiPdMDpMsxs8vqJFrWdvzj2T5iSGRKS03dIogekmDTEr5QXSkVfZDfW4Q44qP9Z
TVx8lQzRfZn8hxYCw6vlKbtu2wGBS8FrByH2rK/5dgrfcu81b3Jgw1QY3WkVNswCIqOBEn/hqASQ
mVeaISzJjbQ2ipVibnWxQFl9AjVyiovsT2grHhXGlzDjFQ1WR3PudRQBGJLokjOHo3TjOzvFQ4/P
RRyLnS2UKa9kt0FoLEwKaeQmLyhi5sG/kFwI1CsQXbJvWXLNKG5Q2Xba6Lv/C+fCTjdFA3y+/QDT
k8y/bVYLJO6UuuztPtuP6WqiQjMlSH1zD9gHYLmxAaMfPGLR/rFKVXLH/lQjc9RfKD+StkCiv6xL
v/zCLdU3jos981ZB9+WMrY1iiFsg8mduSLlovKRQX1+TpCiuPraE5UDJ5TCVzCb533xGFtUQgYxZ
MVSt/fEvjz75fkUFwcbMcul66W8e0CpYNG81BHOp5zEzu6j3TlZHCbTVlk6WPjfGeTg3CRXRApeU
lRbbrs1qF+MOYakduSZwAZKoUPo8H9B3ekUaaig8knBcUzsHrVo+Z/BUtV4nR9uBg/KGuXOWufZm
NWKLpf2yaO+ab/EE/9+MLcU33d+ed1FiT6R0hYnHj/6b7VblUtIBRimRwO6vsdPiqfz7MTTtR1zt
BebrxyYlPFLE8JBajDv9szuo+Esia/XWI8LkjiRXD33aJGpbi7ilBWSq9LlgueRsynOXbIAYofUW
zMojH4RsaXuCJYm5ChBvfvELi42ZZvnTCEV3YMalDL6saBmhiHgxZWsRnI/osct+WkUT7/eSmcMe
N9MNeMcdWlw6wYH/JGV5G5tF/53gxyWo+26twBgfxKOj/YU/NzGuODLNuWOncGEkhlgKtVduUmqI
ixUwD7ymse0B2DKvhy64Y2sUIo7fV7ieKzTKOfJEQz0pbOkYdRWik/ORk6qUTLX6bhgTvnrqc5pc
EBSFrWiu0ybQdoADiTUVtzEO4Mg90SbFirQWABQDICSeN2zYA5GXO7TNCXvGe/Z4ArGnhSH/xxAO
/VUwTPIk2j+oIJQEFsasD6wGUXqECeopOxWXy2kmDgxloipbvRZQOSVQJm2J4wuWEnEI1LZAhHqu
0NDZd1VvfufkKiraA55ORECiMCbWH6nrpnvZbx6H00oieIa6Q2oSkdsbigvKjtcobn4bIDLFZR4e
Wt3as3Ej1Mp+IhipzSwRJsGmvgIHgjn1btN9bQ2i9ZMpYUAk42AN666IVc/OhvkXGVGpAxVCpIS/
5T5GF5Hj3uKQbfsRWF/Lc0nalYZDQ5D8/FQOQiDX+4gIEl49RaKJtjWEq4BiGC2YrNGzNgmBAyLD
Ei3kyNWH5RSREgsbTaze1dnVkWwYgnJmO2yob2fm6mU5MA+5lDr/SgSZS8qH4r7TgUf5cGrWQZ6U
FIxwJ1+tZnHwHX2AgTBvU/GAYNx/TAV9wlnWR3sIuf4MR0cwSs9DQwh/Hx2O4VjnCadW5O+TDYfu
cX8udnPd/T08qLiyNhy0HyYztvvYyYBYzhZ6zq3E6aEF74ok/l8DphVZ6Q0c2weOt7xUktFWcWGq
q4Vr6uMUraSq5Sn7+wm0f6T6724HwtQA26AgR3pvWuu7RR/j6XhNXc9MKo1qQ/VgxB/9AXK/Ul3I
dRe4f9q8vowdhhPzL2PyYJfoOTlIRuZ7mr0W98qU5wSEE4Yvo3HSnc1O8DzqzJkRSlZuvdbGrU35
ZsnCpPhmdjZW0wSs5iU5BpagjxXjj56GfPw4CTIauDoG72Plt3Ca2KD2ney8UGJFErct2t689b/H
lAP+71wy6sJQhKuXs3SKkJ9ox+HxUTZSYz8960phZ5pUefV5GJj+hkpLNiDlnivvhMjW3O2iooVW
YWbGQfOyJar7ybyOze1TcHWPfDeYS3SdQguZ2io3QrV1o9PBBHOUgcyga7aYyyZUj92+sMqRzlA1
MHiPwIvnyDSQ4PvUKDuGCQScZ2QNboxNTVcJD4hxpdA/ENi3LXiRnxTYdrC8HELWrAHv4bJI6GyB
YV+LtjjMvTb2ZNIghgmTHhvWT1AtBrXuTUEHVJpR5Vk93hXpEGFoSXGhnQvqY6/ZXB63DG+Y0Z29
7OkJRX8h5fhNtDxGXs8RCIPPWgmA0l9ze3W49hafqDDHYH32XMB2CsjECsWT6G8MRn5KjckZRMa5
gbNEHq7rw55yRmpFB65Ekw6Z9tyUUcBg1CDFE35HfNKXw/ZUaUY3cSAskmJ766CIq0dYKRODHBSE
Oelu43X6E4TcAndwQHZPgfFOREDgRNQTfU4sxkjhJoBQZn9Hlldm3+a8CXPb6xmAxEjKmBX3A6UT
V2rsaNKj1TZnOmCnfV9vDwHSFnx5mespt/g4PZSn4PysJR0PBC2qUAcY2aYk+ZH65zWmhlnMU+5m
FMcQDSZ8bft4noEe6Z6u5ejADwGVLXJUFnd661W4zUsWrRvpj6shky06/Kb64ICsNBSEA/YHFogQ
B2sqDvVTZFHcFsGNE2TCcVdFXOioyNP+sCPD29LRGglcN2dbcMRqc5EjghSOkJ0ymx5NiDzzf+Ae
yaHlZulfgWHV4PnYh4qab/iJtLn7nmvQgJXQp7PQCkJECCUOpdv8fMJ8G8MLQL/Gwo1/JOOBlilg
wZ8hDN3U/NYEN+MJjXw5px+I2rakqTFTc0ApiTu4PkwXK0zTD6Hr92fDqYEbQq7zxkRnBxaeojqO
oJPtgY45WSmAnNDbeLEL1dXWb8aeP2h+OlABR9OiZGn+Ot4rt41qlxBUwHB1wCMScpc9adIHvx9Y
W+XawCzatbrpQlO+I6E0pzfM6N+XUXFVxBs+QFm5voUs/ecixPD+mOTJtQQC9Tj7XRlQIuP5gkQY
pOIgP+FTcpeTNcJAyXIOr9Mm6qX5Yh3xYnWRkj1d1esnla7q+QzlfoUb2qpa+gOPSoG9zu8yGbvO
78n7QYJbMCVO9NGtHdg3yhHjZ2v4HjsUYpI3zSTtn6btaFyN1+WZWfIa7ShqgpZQc3Je3bPqxzub
logOdJup2eiPVYLlWp3we9zhRJaGE53SFCNq3kySjIhD8Rr7PogGBM4CmTPktHjMcJu5D7DOad43
wM6+M+D81uXSXXLJZWHf4F7e03ucY2s5GOCrIXspCPwCVyrH6D7JvsxLroMFbQz9AJis3FFjVkVi
6WDu4X256uLABzUJ8c+IXxPWKKcVOPjSS/bWmEYQR08tLio/mwHs+UohZMKXZHA52SHbK3v6WzmW
8LWzUqhufBwZ9b3rJW0s93dUGzQqh+S6x+9o1yognbfnCux8YtowXpxGIY/YjCe5ITZhvNdEogGN
GRN4BiIbM2NnyRuP1fE/N/xvHoaIlYqSx1s1li9ukCQXODH5rI4sxtlsnhOtMpwlcAIVgTZd93Yt
ae/UNI4A5OngAU1RFptgJSHYKFWdnr+B7qGCl8LGfuFiY9y8TchD0aa+ugM6NW6n++cAB5JU3w79
qdhOUAomVjBYDvI/gnv2C3Mf7Ke9cf2jajvO48WLp8dIA2af3/SaMFNWMPEt7CjFgxV/nD7uSIle
gnf/E7SLuvJuXw6us6FffsEMAe+cWicJYzpKCBymTQVeKKal8zRsWCTrSD+0kCef+FoQulJ0JR5b
KBj8b5npEpx3YFo1/xoqI/0ahpoaJvux9f5KSAraq8ynm+OOLwOvu2icXGkOZCqbaZnNesbwMzh+
oXwLc09kuXIOm2dHp/VAlkqOZHy3H6VKi6AfvKdQOEA4ADlJc/CScPEFtByhPGeqp/6D+FdNhbxb
9Xi3tZzSu6sdiv07hL6PbnzyBO6VIpQMcfT3rXv03tfzpBgWPUGoMz3XQWv/a42L6FQpanRxD/ak
uFAuO7W7g+XlIZbv8FiJUdzc+VkzzRlnu1HhZzHg2miBNUj/AqvrpWWLWO74CklVRHYCGkmEgPjY
ictPgnk69Dijp6hAeS+lVnhSyJBJr8CkLmAhGk2qQqxL8nxgk7nXVCJcxschC8FNdTzYvDN10PLA
NcBKC8tJ/lqzgwkpBPSC1IqTrrj6snxlEd/P+2lMYGJU5v0gCUmqHBIFVZCnkgegbLoPN75oWAmh
FoSMElF6ICokow9hd+7lKffGD5JSv1K0b0ao0wEtekFUEu/yZhYjIXfIDr4IAymjdfD7wfL3aTUD
bD/s3mZ5S2zXH9a3b5yo17C4K6uqzTIPHTzxOls4lkSbBCxPbSIkgPd+m8GAexl7dBv7hvawQLWf
QxxzwXds+RqgOCEFX7KS414JWdvx+bF5n1K8P8oPEK8W6k6RM1marvET3j3PdUPxS5pBZu5c70qu
PmA4wGHCWjTSZMLVlKnjAKz5H2KWWGl/V3VN2DgO4ZWbS1m9Tw36/iTfdsRsfU+HV505qpad3AzE
lAeJ/EEatBJXqaaDfFq1Y7o1WC7A7QK9BaK1H94xBqlaAOPtCH7ZoNuzBoAsdkJVed+65GOux2Vz
4cxJMHsqmrEn1UqYRMR0SMk/OjV0v+bjatanZiTXIj5NvBmwltV2jbhd3YjFdrOFrgwzxkUO7wTE
KVnQSbpsdGj+LRjFzaP6g1L/RGh8p2S5NRvUA1e5uttDpsmuZ+wqpIrzHhSJc9jiNYevYGJUkZq5
foXhHxvAOv8bhIygFFlMk7hYPBvgMGCWfYpWZpToOIjUqNMSpnZSia6Yp5dwNIGet1kZE9LjDstX
3zIiwfu961CJsO964B+m+wCiDBF9o298KZ7W9qd0Pei62gEe3Q2JJO4Krp/bzY+XhgR0/HneUOSQ
7psX1E6pL/slrxIII2El3MJdQysvgftQqEJG5xR391xK1MmD1IAyR5bSvlPgSQYXgaOOeMTaYxHB
eX9thtVkNoZCGBjPWTNna88CedoaGphn5R15vwdISzjIUlIQ57vbk8jouM2+FxdwonjfeeughqIA
wgYhC+l1+TfQP/kuu6UvM5Wy4+J7vVCAUCGLM0E+Ou7Ji4d04ncGmDlUUhFiJbIdfww+CF6ernOJ
mcIyM2gwCQDdF9+mMb9M/P7+UcAIevwPGhHefGRkLCYEe1NbTFZV9xkMfdBqtint2wV8laCJE2kv
q/+Drw0eoNP66U1QYX4EQWQEDyA1YDcARYtnNhWH+/uw5Qc/ll19O4B9yODt9xuc4jRWIn5BUVsO
tGQWdzkX/IxjPTgwFTJvQ8fmvzWOos7qgHazkOLKB9x4bnUwVO7kFMIj2Ho7fgXGeQm/b5/CzpTy
zeOm8iwlicP+CGs4D5HoYNQqyqTviIf2ekCnq4q7kOm0+gsuZkO/SIMIC7fmK8Y9vR+9EtsMD+rs
qDgyd489vF1EfYGbVKOj9lToGRSeJde2ziJBNSDE0MLs2HSc8joyL03e7L8/M1G2xaYhAHqAF+II
lZIr+veZT+j1nfvhfh7Ux5MFzFNOFDL+wpTvbIfKAvUsz2SRWkGPfdXuVtjhmkcBsXEz9J0+H43k
x8dZmCdjBqTO/giv1NKB5p1nyFF7NLSORF37OSwqFX/9bFFJuqTGQXbsVjnYFxLDvMnignuGVRXa
Sm0tAU/ErID5jto+2j2U6Cuyuaw0gRz/S1zb9Sl+mv/W7u/t9g9UZdPh8lI42AC1/bklybScdUbA
xJJnMhES5wM+tndqsOVWITPyCeoqW/6JQlhjnd36DguQqcmEwozQN0kYcN/1of4Dlrk3/hnNy2PN
O5AeRGc7QboxwR3RNq2Xbc6wTUurSDPQmXHUzHWyDhutSunoaEQeMaDN3u0gBbY+avWNarBlaVEU
Rj8lc7xAgxi/GUR6sq94gZv0d0kxDvRKmR2sGZd4UEdKdcVCANV9p6427EEOQ8s/lZQP0PoLjSco
DlaxQ1biqV50gKKHWbeFu9BHWMHcqh8e0HCnQ5cZbvKALYXqV3jTssa062zPOFkhtUEw7c7NTv4l
JmsQYuHc4CaXJPEU28787REluNi2hNGJH0c4kurQelQ+rkXzhjNrTINlm6gZ2CZcU1qW9U5CkXeh
wbAi5IfKTdd2C0UBcXkjZPQ7uHx1JT+Ob+XDNkMlCEwNZn1uZxDRQd3xd1nnQ6DtaOHif6hAgwKW
+trSclYo2HSI4G48rbkrk8HBLSsC2EGQNKJmH+d8jZHuLg2jXylV8LS+KEa43mvIRwzw1YOvCBI3
upJh2z1ewiRfieWOH9tpwqypxE5ojFYgqYrgSmh6A/UP78DwwNErdBKhtnVxLuXuSB651yjJJHeA
dSKMS+wgfzg+FbtVVUR5WRxkmRZ+UDUQLIG9WlJbYI+hHgnpl0RAt71TbL+iOivU9rTJK+p/8zfC
si5gVewbHIy/GDnN1x6JTXJi8m/Xqp6z0AGMnGygzXZlP/PJXKMnChb+KzS1sOP2Wnm129vZZ/Ro
ToZCY9vwqrSe7Z6i2cKEFEI0ZD3igBRV75YbntXLaJhuDVCczKZ4qOHIy/jt2vj8ueOYV6MwO9T8
GCJ/Blp8gP+AivNTXU6xjq2epRQCsRRuFNBSHIAvqynyjG8dwdRAZpR/Epj6nuBE4XAEuytPmns6
+sp9zKjcxtICT2dcQKKimXnFQ+RpMIb5VyffqP4bCOfU3mwpqeZRQIHULrVuO7mO6Fl4uGdbY4x/
RMI5ePJzzuFALFmvnlrhGXlFn/c8y+rX5SQotWxZGkkrj+CPjI6CF4tBTHy0owW0449JqkdOYC/D
Y3SynP4/lumWFsU6yFD0Ei8bhoMvt0Qxv3L0GqImJOMnZ5mBjJjqgAwS8Qz/ZwSEzSbO2njvUXXV
pqxcUrUNaBp0nVw/ODhcg+JFwK5gs2oM+D0TsT/M8G87cJxmmy7Aq8u1l9EUTdGLMRxImIB49pRh
/Csbn5iLD1Z6TowRjJCL7D+JIWTKw3Vk5xn54vLpmluZg4tvZpqSwpv2GjqojRxqAjmKkvZ8tFSe
EkMlceozkYP5OTjQbcGJFZMrHrQi4WUt39ESnQDyPN26LVOxz8625cVht9vC/EiRs+JeYmj59nzQ
yMHmHpdJhGL5Hl5kDQi50jXoZHYH/qORpPAJDlD93yOsxv9md2WW3sBWl5ujlYwmUnFnT0EpAL7d
U7/a/wXnGCkRpxdWWkgN4OWGizIZkc4mJFjOX6GbaGv20XpEjW6SATZP88wUvQHN7zSpHnDe0SkZ
T6QndlVb+PADBnpVUJRwg2DExzIvwffz/XS5Lm8+pU1GEk+ZA9sz144gh8zXGMwPZGqnUwSAzN+j
f1IjY1Vr59LmdxG+PYDjo8dhrzbrvPDAk5fk0/rBs2oA7onEDwRDRiC1lwZyDlkXcqhzGWl9cdz0
o3+zMtxIm4tR7TJYCq5vZCRQ9Y6oafMApRW5OUxRA8sMF15OLlA9vhfpN4kyuWc/ebsZ33wSsCMe
nYdZz/QbyQ904sOILXAh2hieswyMdO9bhfsO2XLDvaicuYNXYHDEFL2CKauV8wtKz/3znDPXNEhn
irJLSyhGKYWPw4/q62h5Mr4s3L1jA0SC13dzobHwCDU3B9/B6SbljDZpZlJJyxnDKiwv8XojStQs
AAFDIlkmBcnBFkhcVbL1mrhDFemZz+slaL4dYvCb8X9XV8X0cC4/MNG5bu6PX7kkfrbwlC4wLuPv
pvV5noiY1ucphHtMvzSIqZdh19/ziVC2v/83uwNF1K4GT9/MR7wsojnjXxgzlXp14ZBgGHRcbCGQ
RDPM6wcCLGycgYcxiKTdxfvFF51IRh/HwdPoaP1JrQS3ke3SjKnlJSmNh2aCOMbgMEudsYkrmt+M
eSuPxjOuRdI8RhJhhQJv1gV5Ud2v5CWdHF1J7f1q/Emi5NyQ9HDYlOqBYA40EqF5kAq3DVXz2lA6
k6a2NO7VyGyqsjrN+wvJxSDGy679F/rg2m4Tw2aLE/aG1fpX3pV6ybA/6poRB9n/A0OonpFKFB0J
rSjUT+dy3jrM8QrMbGBtl0rgODfRR+TAVBSxuF64Qa26ZwEch5ld/NQCNmLZKgnmHiDzYwPYrvJW
J3Nu+xJ7U+g5lxSjTAX4PPRyDUdiFr1q5Y0u52oQ+CfCMjADjeGyHheGrdcpUJuYVynVKrIg7ofV
MvfNrTrz8b4lVSSOol2Gn7ceMzRXvbJ2XZsnNfggyR/QAc0In1fS2S6r3z7YMO59tmPdQeZ39Ajx
fPMmGvp+9Vx9cee1PW+jN+OKdd/8M0xrXeK3aNCby0QKqnwr9H5TDcFga4MkxG+YAUIW96hwO7X5
eOTx07FTD342Ba71MSPr4ieiULvsiP7S0gHJ6Y38UgCNXGnEgzy56iWBME3ydnc8k9OIcxGMwKXH
y+AhFYdxFe0H11J7t59TaN2O532RyqJe/5qNzsxxJC22E96GCGj87OFQxS52Ek8piQGMOM3rhtnI
jtWmcfZEOtGmkN1dV0+v6oaZuoal01ftJSrIA73wA7lKbqLRlkL78o86RVizLainm3QsLXbHtbaZ
lv+3kgAQ3zt/A6WHtitJSy7QJfdTE7kpKbDh2oClMhfU2Vn52+M/Qbd/4opP/BuI9evvV3ElxnYu
3MzPbiDVQl57BnbobaHYf3XWwD1R/OSkAGo9+t5aPKVhkfzY8GNZgxFh0HyzFOgvyWyLRUSXTSXr
3odFr4GqdAlJS+/z4p0pyGq502XSze6aoPQHFXx5Y+aXAfhWSo66W5Ivs3TkfrYl/WInruUECtn+
yblHVVDD7xEWotJivvRihVeIjlID1lzd2oeko5ttDBzwodyG3OJmB8sjm9evqcRok/FZ5A48QufU
XqxpC+v95NNZf/CmUk0CAX1nSwGA3FMmrA6TKu6xt90yomuTc3dx5xIN4vNEfVfigRyqpSsrBvwr
EQJqM37tt+5gackDOgPIJeaFuGEhgoGusaYu7dibT26ZdX9CzVsdIUZnxy4/KS+CYz7slgjwKP0z
ehY8p3hdik5Q/cWlo5M2yxkHcn62p4VIzVH87/oThYRGn2ypxveD6ATX1+MPkXZLo7lcD4KkEc6y
uw0IkT/siW5oO5eLVHw+CS7NWh7ELU75XM6jQZgklviraDROV8nsak/vbUA6RVoppntvQes96Vms
xR6d70FN4/5cXOHWtvKvxcnJd/MvtoGKSyfxX5u9BVUh91cgs1GYmmTyMeGss+hls5jI3OGCb9uy
hsFynBSkXK8rLgjfX8MTE7jOfJtVEhGZA1UUgOhCLYvyP1DYQ/jmpMo0Mhar24WxgWMTkxfUTTj2
haonEkPKdTEYXt5S0X0Ol8Uz65swfi6AQZikZbK6BFj2eRUsl8pNZJI6Fur3Ov74+pjUUhFtzf6Y
WBuVdRoQMDYM/JhShRu0p7JMWQT0i26z8K2RwbTOTEkhZjEpIBbWWYWfHx0vmzHdMxmK7y1Qitrg
t00xpnJRiCR+TP1R0zudXFWrafMSBIWRYN8+RPRrFlPuL01Aw9cb+aZXd5jz9USz+PTK1QYOg6S3
yZkxOuxgjieCqDz1Or9hmYlzv4AicaC8IvwUJnnNW77JUdJeuItTDG8oxZ10gRxXx9SwCxZ8DVxT
KVar54L+H1/kYKwZfkI/pRcyvqpEM+a3IrNl8K+6bV8FDs3fSojtdheus4FgFshwdeU1eTTAwUIU
7ESiBhcSJ3ncGGRBZ9T8EcMgC09vuyishs3dl0BZXvU6IE2UOaIExgM+0DeCl+i1+mIq/4WcxiId
veznmNUHawjittQIHZ/3iWZyflRg/cyU4K0JKObbwGOPrLLGVhKEF6Hp6tqA5qBTE8aOcZmjnx7c
iZNna+x0zHq6fEKuLtQJzSoO1ss7BaJ2wQt/LjR4PpiltUlIyfBlCcl3sOTs70QmPN0cymBxQ0ec
RmeyltALcsqxXo7eFRip/t2qBuxw8uMeBh6Lk3piI9eylgF6m+G8izodifTW3lQIi2dpX5In4fc4
Wz46z5104JAlABoINaLIdpMwiQCj5utUInzFLlU34n26YoQ0BO/xcVOWXoo9rOflMBQfq/j7VMz6
+fi54R2/kU9m5DFDMz5ikRrUkMygCBcm9fvORtP1ngyytQwrLi4brndPxpn+Nz6mnWGH9y9xD5SS
MFBQP2iWX0qArLTV/9SI/PSuDs0KxWBlCUdq7S/wTs41OvsKhNyXfjRwyh9YhHbUz/CCT8T7xgLZ
X49WENTglc3e8IUxY7VcAGgmApEV+igvRF+ObzXLpbF5+adEwBghMqdWj4YoGmp0hAXMAXqS28J3
3CItR1/sdmYP/oFkU9ZtJBLA/Nm7xXKuCd3mmJjT32ehwtArMoJcHB1s7wFq0FiglGJvNeJMS+zE
abK38+siB7Pp/9cPNCO6wM426XxjrZBCz1DESxC+8/K0zCefoJYQPfI6+P9v8/+wXdhrdb8lADGR
fF+BqoTbYgv8Zxd/dqzwdTcbay6J4HzGJOWqjvpBghSZdIKJ908eii+w4e6dr270TySjy5b1ujMI
2XOpFuoasMklY61zWKqjlTAnMgFOtD7xleWgdpvjY8M7X06PFOUMmWvaXXhtzIWjzpEDd7SZpnhf
Aqest+kHSvzOYm4RoV1xm8zN60NrzK3k4rEaswVBOeK9kawbptj69A3HyjI3/SxSiuo2voFh56Gk
MpqDVIu4Y5rzu8jaSA8uzqbUiLXcD0c1zWPII9vLRu7V/a9VzwYk1mi8Cpl1QeMZISBBC57EGiqA
Em48LWNoLVd6gjlbbsecZbo9EbnTGF1Aht5ZvCY4mWLUouP0+Y/aYV0j/mVUzK17Ve3V3MTHFAkY
uZdMgczrryluKmoAFxT3ND6hyrD1BODCbi0QC6DNUWeR9NgQXc930R8ilYOqnt7tIrYyv+81sxKC
sOpgoYLW2TbMl2HN2rIsdrYcm1bu1RyICgAZcjdna+RpHuwjAwxtEp9oEEyipkCisIfKF8V3o1+t
W7pKm97r58ybKQdk6u7iRZ5mZoGoweg7JizhihQ4+htGTWdQj6Bz/C+YABL8i8zLl9b9mq0yKRgc
FNox+BMcRfmMmC1D+M+5QLFInGo39XQb1NKwighIyMzYpH1lugKETtJPRaLhY/n7dQfrQQ/hCt7R
M0IKqAlFqiSLt1xppSBTHz74Zsq0PsakBLCjD66JqePAiIV8wwrSWhBQb7x9Z29A/AtJEd656H+b
5wNBwgLr2WaOkrxvzaPyDfoRySvt8YuCIY7s30090UOiaMDqdvdWa6Psdvrqz1gOd1cLkH1lJoqL
TacrWxBDMgrbWyOI2zidJpCILF05VDVr7YpiI7ydofpCoGWH7amocFYYG2TkZLpfnRZKS0ZOSjyi
BmtcUMwfgZGf5OcwPQFJje1NnLn8fKHAj2x4k8GvtD+kVFtrOU22zT6ohkFmEw2zzZpkhY+Za8sd
f7jb9q4MI8mQZ+slcNhikNkzxbVdr/0Ixthy+3YZoUfflM6+43wY5IfispDk87QsY/qa6/MKYFLg
IvNhUyVrA1qn5SA2jyyMJG9rnk21EseKkpCQ57fyqQqzYXS81ou2VKXdTWOl9WtzlYr14M4fIKO3
LNP9xSdiuieemkqff4X0y9b5hbftxItfq6Wh1hlalB7/eBb5qYn+Yke/xJTyPITvIppWlCpepcl7
rgbaGIuVz8GA/k3XPSKnZ7leUfhTu9viaN5jHrPlMX9kSYOUftPS8lZaNEuvxjXt1YVjkVtqVDi1
gy884oIc7z+bRk8ZXTU1pZUplGux7NYy+4v0ydKGlUSDKiUsgC92ykmZUwF5H1xYfx2oRSgSQxYC
jpOlYbu6UiFS99HlHt6Ms22LollF8GngOTRH9fcXD9njxjG+6kvLuzAP83iaNgmFZGMWg5ihCchv
eLCjesXC4Dw/MJUalBnC36Ev/DuSFMHNN23+GblxgPQKN1c2kgmWa1nuFe+pZb22zVIn8bU37SOU
iVZTdG8/UN0l/NBXoQqdNEAdZMvjeKkjfqxXZTrABEGBY9cgcyiZ6csCNymaRGYkfhxgRq0VI2+Z
tEVCabCd3b5IHr/JUEVhlbLw7l7y4yTMiIXgZYnK/rzdpST8yIRWfZQy0gX0w1cmmRmA1uF1hOpS
50JdzgpFLa4xlo4MUZtSkYexSyVHmUg2b1qfjvkR/UMge1DIqnjv9tHzp+7HQlGnWqxBM8JBAYQf
kfNuzPPF50mmjeyCyGtu4JSUAiZ7pzDTe7uSKRk0nHY4M3Ic0DMHpPs4uGayLtM2bIBzQ0EUy6Sf
3xcw+Gn0H0i3hNEwOPrX/1LKVoZmYVWlbGIm1kPC60LwDEuSMpeg2wKi6ToraYrWUr7NvtuSaYCl
Mdov/90satiXL9wcxESoYnBrfcDJ57Tv7LJSMqKKBKrdRXCoURUWlU0dGSf2tTGmkAw6yHp2uAGo
2G0PVi3TLvg0U9YKub3YckGe/V1K8BB3xd+Eno1Vdsd+WHp6pR4q6dGUTLyPUnvUYSHHF+AdM3wm
MnvhyMCaRtfJqd7tR1Yfd17kCQwK41vmincMdXZUsRSDnWIVmu4GNabiJog0Smh9EU51AO2Ogf89
LUofzlzfFVcFastPPN/cWYnuZN9YiyK1lklxaSSYH6ZCkgv4GeJ/tLPIS44vOOl89gPSMwRNyRB2
jP79JaMEl+DYujfYiEIabL1e1GOSb+W41Fdv7SPP84Cz0aYVgjokpL3QI5QA6i521SzUUeXzgBOM
J4sfCyB7QngAHjccNSO0vtVq0jqbSTBwvgSdiPsNN7Ym6iJQV4rjkNs5Wsi3hsHeYXQ1p+zYDHxF
gM0V90i1ZvvYlIvf/wwFZgKG6shFKTb4VfNTf/WpZhbyJZgz0Gtb7kWG8OL2JaPbUGtAC7+q9DTa
NGp4d/q6zZOYX5DEV0bdGCUfCKw54hEpUBOqZ0fLJuE85oHAHoi6NlBuZ0Tod+q6HDwo2RpLTmvC
LpcXwr/VcBVl5Nk505gXLo2YHlfOLcxB9JoAXXn5ReT+p7+ykj9I9BbwQYHmaIATTeXY/3QIACKi
R7qx1kKhGcqvVb0hJTjFduqOlUiaKc00WfGfCFtFS4wErsvpq8wWDCCYxbXZTYUMrxjHco4BfM9z
dCkzH13MsCnEq+xkaejzmN3mJxbqHG7CfWelEsPIoGa4JcXsTaKMcHgJydw943hTYy6gvRQne8Vn
6kCNd0tmALLs0ndqQdzgqNgumeivKRi1a5O3rsm0icAXeUmieCUVHYs+pMAsjbiEUPO+hq1eIjK2
GbclrkAW8K32PBhDXrl53yKOZ07Uk0fuTwMIBZ0Gkeq1VunJ/kTDIWZ+r+29JfMgYhSXQ9B4MTvj
OkY1KavGClNKzzjzvmM23hv2dALc73POwQRUqnrMgNH5UCW9+L5WBLQ2SjdNt9Na7wF6IzDasZEl
hPJDttgJHY9hhd0JrtWRsaw+DgPzkBBR2bifP7TXkH07PG0em982bp+XwxW9FDPQE/0N7gozlaU0
oyvOqEAwjsrMBwMOOMiujoNhwb4gbZbjo4yXawyrvb5jx1c5980UuoD2Vv8xgU+9innoHvsE8Etq
HLZ2k6LQ81TsB1AY99YQ6bpF8Pyiam25zgZ7MLEXUGrfDCyzXczzoXFv3hcVMTa5C3zM56H/hgNP
1ROcYXNftdhVFSgUEp+cdraQWH91PW3Ay5J182F16ZIeWOOmItH40nOlTOVjduUGxSVw3tReY8dA
F4Fg3aciMlhA50oef7RzvOYcQJ5vF+RYTQ0Rli5Dnoe+2KaxpgaKSwbiwDcIbYzitNYnSFMUulKF
QMAf2osNWPsvg5fXRJLNGrkVr7+X6qLRLmIh623IKjdoEbEWNKT4J8o9yi19Yaujxk2AN2itjzOv
oLCjzGIKwmRFuf9CU80xD9Fema22VsfKsol97+EfHJf+tPs4x6JVBkp35+VX2Xw6YSubK1djbjBn
8hnnxwtAvi2brcf7LbXzX7aEig76tpMPoQPjKd/cNSKMgGBG+53KeG7DDdAH4qGOLiJy9dThponc
5dl+wDvWMW/EOqzJFReMK4KzPrBp6DBvTuTnzGiMBWGKC3wC8Jhd1n5+fKO+VmiDd2i8KczTO3r3
Oflx1z8nVeYGZEnm1eDoQezENWmn4DUreYHPBfDisuqn5vAktZYkYjzwQouJb+hD6kngSps87yDi
LwWFZiD7OcNaqwRK/5rkipasyE1gEP9nFcPu4134DT0oBgyiMg2bwP/Ex5A5XMAtbbq53T9kJIkg
CJ0HErDdPsaTZaQvcEGFmzkGydQIlyBPqMVC+09huoXMdZvdknIXfqp3/yhWghGVyFftOj5Jewlr
1dIClU2OIwiau7YQVnwjqlPLtVyU1e4r0uk4QXIVbxBIwWMu/FlXUKTtLD32hQ+ZyefYxg3uWNGk
ste3GoPI9TBPwJFxJhtENPRmAJdlvARPMSlziKqvWpV7n5EQXSiORICt3e2meAe0yCFy9vLohmHR
LRf0GEFP36E4DpSfBjdxBSoTZj8n2LH+bMTEiemXdqvtlsNRMsFpb+oRg4BzQWR5iSfiK4P6FEGN
qZW01g2MKoUhpX1aaHv6mJ+mLkHOLA/dPwvVy/jj1s/7B12ZJ23YIVHXVQUEDfoTNQlMJW1vZLFK
E6AfjlafhDrVMJUIOtKvhhhjdKyErxThH/AiSbE+kFVFo4gXvVzmJmPhiUz93MTXs8yyxAaaboWY
sZ2N0QbyNVljIXlj6bqTbEGonUiek+5Nf6BplQ0qra59ongHBwDhYS11bWn1u/My7iM7cqQeEbH5
MKy0bfXrngKcT7XgnK06H/PBQJquA/YGWarXDjtnlygFC/SiIlosPVyDxCza2BcdVpybkQi/Dtz2
6zbaDTYKIk9hEPFfqY9/os1FmNDnrGcjm5Bn5e1HBTN7K7dQyIGCu0loBbbNS3NqrlyvIZPFpTIu
CIgORGT+Rc02yRBoH60JST1yLWxRhWFvDicldFdaC1UdP2QLptTSFg7zK2VTSlFNKQWdi34RYCej
f3IHlKDXX5Kl7KN9qZev1wTYxpZeaEuWhuj+jepFQxAjNY/qDJneSj43D/ZLD78FNRn+K6HKjvwp
DDctHLMyjHPuJRC7Y7wR7ximNlQfbnf7s+a4MpNzrUBpZZS6MRNaCuspOC7G7SiSCOWiVju7gRj7
gqkjKe9gIQEXq489At476hlD9bMcapBbVFcmU5kQ0GF5Dak40CYBHyE9TIXhMtjv36WbxORlbjPv
idBMUJqat3FiD6VvT3ihsT+wXfuK+UOa785XTGCeRrApUVbeHwfuZkZ3Z108hO8ivX+MSdfXKrHt
wkQoK2+0ZfS8mI6etVtXjgPkDKLp/m2eKs8wslh3sWLvcIUQNyCgV1z37Pzh+VtJCM0lDjpKL+v6
6Mgl7DIUh4BYdgYV2FnTW7WfNWQD3Uh9sYoPuiyCXft8TYwnei68btqGC8aeDF7pVWlPNqLvCwf+
O/GwvMuhvYti4ucvBU6ZGv5FKvVm3dfzAjtqPUfh0nOvUEOVmKVxyxmC9TgBzrEHgywWCpQ25QAL
dYBtMWU2a0SlqePTocKQI/xetRk3L4W9hRtGA6g3YMybPHd+vHARprukS4XpVcLyF/SLvU9GGGq5
9/yqJqiVHJBEdrm53wjljjSBof0/SekT0dDZ2jhfBAaoDSnOhM4fcTfAHg1JivPDbclyVlMebX4H
HXXs0XzuTfqJu3gqMSQETvbOs3GlktOISmsh5LYOeoqciw4784jkrYnj7ZgyqE5S+0DxSDzfkoax
+8imalCBivIpyxuj5++xKrbUXetE4rsEI0GCrXkVsP91AbOr4xzz4oAEAcG5qTCgOT0tzRCenX+N
KR7sqySGmaoi4xew+BsB0UR5y83hND1oNCZ3nd1gv7Ke4JSOcSJYf7yiFbrfZ1PrOcdIz81tz79z
Rom1QVFLi86x/fXBgkD8USVWleFWMaCYnNpRrKWdq44UiFrYwmgRX/AF2n+/8C5HqDkxUi39Du01
BkhMjELEJn1nxfcGFNkidXAnKSTMO/lR1PstPvOEvGH5RkELNwetMWZjzgUxxijuEQMmcJDF+nVO
y+Wi6ObbZ1Du5uw5di1kjiB/T6tGJxdCV4hchwkhV5tsCKRGzV70UVnKIfpkfOdSQlU4r1huFYc3
18gxuQ0KCflESQAiOcc6KU69k+zvb08qIa/BvSUKz8HOe3lxUY+hgK4SuAsgJboduk3k6AITY8j9
mR+wYrloAlECiSg7tS8IXgOpBpmFdc16h3h8NY4MIqeYA8GL6+gEZIOTWiqe0AjzOoLjUMabYGZQ
V+oycCGnqrhPjCl3tdQsWaQ6y5OoTgOnEKS9+0BLpF4pY9fwx8vsmtOhjrB9m/isX9XlM2FdmIcp
zQ9Hix2Fxynk71MijooNqsxr4FoV/eFMEBScW6ose8aZRbXI99q8bN1eluaHqlnRZCWCe/WsfNI1
CUldfiotp+uLkgRfCNOcCXu8cS/tk4wCg3LKE6R/tG2afiHLqfvPPyWquCpVZaQNZ9tjYjL0aBv+
gu0ROm2q0vrsLKqbLk2QnMtrcBMB7KE1nWbtqM367nGA1OwfiIF/knZloHh5Zih3dH11Bbz5WJXA
ktLjU3efscxyTOKEjCc3UKRjkjvCbeGd1h+7wv2f7GAAbldQ1F+l4ssqOYxdSRdzzp7h+kM8NYdg
QY9Zxz9eeMvW0xsICmvsBxilW+/G5d2xKOKbo8kBMJcJqlSJsrjYK7W56XGeH4Yd0JUODCXD1Li6
AWyeY9jS2sBJVcAY0QHWM+wSMHVPi8ihmDmCWXomJOC11sTbmVWA2EtIxgzXj4DfoGny4rTt0paI
EnE870nokjdhN6u94WAMnwtpln1awZwMWXEEUy1dn8R8kQqgNQ0VWMh3TiAdk/SZkH/DAtA60yqG
5G2sPoAyNlnJwQfp7Q7olNkIdOaCaWWEDsJMR0jHezmXT7+3NUuqxpELX6J+X9VQTSSzyRXsP6vG
5pTCR0AZ2y3+rczrIAfeEO0kgHGGOD+QsgZK0MOc49x6SNULE5LpHACAk9uzTSnEpzqy8we5SSyw
O8XZH3KGVc9ZojWEpsdxrdaGX7/3SGim/JGnUks0PWljvX9gyivrV0HfEjHnFTc/G9RHEpzBgNar
HSIFh6lq6CwVQRO0byiqQcw6W+uY/twjzhN0CKhnTf66gAwRLeHg70kqXqcirHcwIjIl0PSc+tXp
vJJgFJOX2q87BgqqTwqJO9Q88wJyFymAKDVbQZDzZ0xRgvT7YK4kpxhloJRkxQS9CpHqnUItu5dp
oY1d0jTrcUqzHngneruDIp5r33OjXsWm5enTxfLIe2AJp5ByBOaRFqj0S2nKMOO48wROD9iqZikR
J2FLW2rJ0UIqVE8IPiZSmoC6F27DPE/7+Y3ZwrL9iJBUz/8ISzWuiFkUg0Kfb9/F/2mdjMHrrydc
ha+POfnHXAKlJmN7oUJNFPQpElTmEDi9rLhA0jRPhicUMsGRMDELhtTHPVS6N+eAhLvQv3GskBgs
UjX8IoMBunUvhTucefLDU7XhVGJpIezd5/0wbwH7jmw04skM6b36arDrzuje81yyEAJpFFGC4R+L
Sw7u3/tyxCzpVHN0mdnPUtv57V4kNFoocojd+L1meDxo8pvvZq8NAQoIZcgn0eCfRBY3aYZRqJRO
xYimWkTOMezMxXJ3VPJcZNQZAZu4TdBLGOdExYkiD7lLlVfLNIIqPc8vxogVF2EGBKFfMItFRxow
GwchdMTEyiI8CAnbRuQWKq1Iwzz2QcbF3M5j/BSHOxikUT9hn5xm0Y5P/uMbjpCPu/6sHyg48vrw
MaDJ/I2W3gOoW4BWwM7VvRWVgBuKhGbW5jvilmkPKwV8O4jIqZ25z+rO2NKsz4Ac7CJAFuHS0TLS
tg+2lccMsVxLmCr6wBhoqgmIv0BeHNIJ2kjcO0O9kmJ3uLvnTM0IcleSI38E/28OlSXGwEVtovBk
qnwblNU7NR0RlxDe3OCsld4rnYyCp+r+pJCqdMuSKdU/7Xdyu84cnAUhjw8uoNtk/VybLaGy7jxD
NuDJfAT/qNCoEZNWl2xgJ60LhU+uVMo5qbNzeDpVXCD0HbYbM98DACmnkJAd6L/8kvwh2AMgBM4x
JmomXnAZsSoh+AV4p3Z3Bhr1s9EZJ4wjT6Ewhl+jCo1f+G57goSV7nRK+7FSwOGIqOoF+fhM+1tu
AcBhuuDH/SBzf1rq1abhALPj8/i16MrcQvcdoGqNQgsxSAUHcB0W15bUhFPg2KFYWd05Eg/Sh1y3
oxTMfjyXQAHBKvHA/o9Xsz+cuTdFAMZ6PA7uS9gU4tDedzT4xFUVdmQAthxKz/eZtTpDvJ5u6cgk
TjopaRfOtF2+9LUnd++q8WDzX+NSdU0BCWqKLEYsh0pWYFKFLNi5ZYn0GfoQXiTUVOJ55iujGJRg
gwWdT8pczWkqSrLZgLR0+j5fucwP0Rf0UtDxOX8IGE4Go5JvpP/awuVyJ6H9Y5zXNWq3zI6Xi4na
RrP18oTDGmdF7ol24KLeTxHjQX9BNY9QTwGxsvNlJ0Omtemb15iVYSh4yrsmdCnHZDhimxjbT4AA
pJRZF6EPpqpfft9gMHMwRGtsDgBvNK5sGoXKoEnXK/2zzG0rXLStQgtWfiKHBO6aBa3/HLWRUMIr
Xkj+ooMv5i4F59/rPFVGQzjY12XKMx/OdrXnihW0zKXjVE8RsMSrhkoaPqmiQmZh9HOa5m+6lgQI
JscVWOAEcilJyO1TCXHNlZhO0kxbRFnzLGQO6038LQPQHfSeiNcx37UUpbeaynlqqPNCCztgPyAF
jL0CJP4uOgIuN4BGAqCtDdR5mJWQfJWERsS7Z3iH8YwY0j4YgpbIXPB7kRYVpfr2blp1pifQj3gL
jKDM6nYXRyu06aL7/EUPm0Xb96LMU1uNERM50kLFxmFFxLgrWz2g/Z3TYVjAr8iHhKpWUabliFkY
4LdsuyOQSloJ2jPu9In7/gnCkmiOlgK4FmBVaumWNg9IEK044mROy+z4kDKOP6Fzj/smnTXGm2kn
KqV1hsZVdSmHkgZ4h41V72UYEIGxLNGZKIJA7iEo7jV6+U9rdoV2ZsXFNINJ3cjVqSOyTauGH/Xx
Wx3FHLIDh0HIk4Z+zjqJwGM4QSp9zpoFZTiR7i8N5wql/uTSRsxlo4V+skrUSlhDn8S6N4AhOPF+
Xl7+s/gXZ9Dk4xjdB+nbocRGOTAnBqkIXfIIutPDSUCswqbaxZq2Trjetbt9A0tgaTYUvt5GHFnj
nk00vvy135dlH8eJgP/OxHJ6Wqwsnykj4T0tLn3CvclmOIqtkURk0z6ReE2mJB1ZlvoUiyJ8YO5Q
r7Q3x7dK3irJftLbR4MQjaV9wBiQAiVPHGb9vcwDLBIV2NJvgQHYFoEBtgv5XQVdtbJ5feOp8TnM
5RzmQntbwb3YPajerPh3LCdIp8f2Wdp0o56btI5apL2B19rPfNIYM9ytEVfvw1pTU6hfexMUfuiv
NfAbgkQRBywuFPi6wnTN1OebtH1vWtwzDpjDOqLcgzqOAHOQ3z4i6IF6hYypaMZbPwxwfwDuED3v
DnYEfnr/THrGN+imIEnwLP5dwSaN6TFZkdRdP8wMDRUGzOU1urtTP0NiztEeoZXr8M9S8NKRvjNU
gLt5qT1q/Hditpnjft06QJNOW4peK+Ivc4pkCy/jxhFRhHYEOmgDxQC19bpNXSRz5ZPIo1Uf0nvQ
T5UfiN+Zn1G/cA1plpHDcuyWwQCV8CT2qse0VFyyhMbEekxJIIr1MlmxOarl/k+JiUNSj3kVyk8h
O9YXGZ4UhT4EQ8oSbjAd/CxuPWK/noZWAGuC6VVLeX2rrnE9QE6ElrT+519kj+KapCIsS0qumWZ6
LRRiB/mrfhfUy/u4In/+hSA+E1a0zV1Df+mJofWL5DzhyZlbsnxrLQETV3V89EB9aBZGQxon175I
xTemVw00dEyUtrQLNjs9uA77eM7osXmfi41oYH4OCpH0o/cgRMCOpcgPvIIHFD1+NDHawEjXtjk+
vWmV9x/xWnUuDKVC5TKMrB4PtNzmX88LFvvP3JtbPukVDw0YX4V/MiaWsHB4dYJKmivKX9gWI7VE
2X3rxqxFtJP9oh/4vCB6aAg1P1yMn1TYOTerf67bi6uCbAlwUfrpp4t6RKr7LbMIVANozEyD1+bA
XHgNN3bdvG1JXcmj8ggHnFFakil7bcRP4SnalDlkkFiqSWSxNnuDZXeAwQH+5iO+8ypqQ3kIAFR2
1lflTmheUDsmBUC3u4uSfXuO2CwBD+DeLx5jTNr/fU54jbb+45AEr4CCxZ7l99+bMFCzBT87rZ64
6wlBHryzKPiDRPHW/YmPpSvR42Kw8P/4KU4TKrpxk5ELzzBYsJysSygRakMqUgQwpxIPLl0JLkLV
XY8pD4SXfIucwcsmoNvIB9x8wDB9otBWrrRXFaFpCW3GROx8Ms3fAfyz90Qd2WiNLn555lqXztzZ
uTAvZkT83cT1FLk1+9VKz3GSsBPe0O4t7QNoW+8WgJn49ISUn9Mx4KvnBFbfM6N0aXfrOgDFXs71
0eAq+d9oNlcdHG+jSBXb6sWc2tCtLTsb8REgt0L9JdAEQy6K+s3YtthGP6e4XGmC/FEKHfxMF9HY
o1O+PoaeeSXswjZYiaufbPI4QIdKvW6fhLm1jqRlfA32F0bn36aFtKW02NFB1764dviWDXIdapIO
bqCVMwfDWLAjwy6SqIyOMRJBHzcoK1XferbR9mUS8OW+OVOp3nJZ1Z60KFndxxNRJwmDZEU9uDqO
fl9kSMIQIU5I1Uxl4BvenR2Qgv3nA3xW7XpGuN1GTu3jZbYxk80nU7xLYTldymTQtd6a5XMxIb5S
i0xYV7b1VtjneFZ+GFZbRAT8Tzj2WzocSAaCiyygcgr6CTuQ8H2TPzLtit6f2ZZK6RpcVydo4F2z
WgoXbNONKP4hBOZ9wtmmkP3J5oiYLX6uPenwADOHaMT5sU8FQFAQUp1lxUVur3VCwB0m6G6jsBPk
GqqzyqGc3ADbbxFAlU/Wishm3kA9maDB3eZ7bHioydq4ZPtrl3M0aCuj5oYtlMXa7FmzyFfVx1zF
ks/6jguAIT6gQ0oFtfZRyf1yxo00YbZkrrVer4DE1uq9lacD5dx48+/gF1t727/D+4ObFFXnbnxg
d2/izOb6N7OZiETVpwW3TEumFl7K9vi4/uxc0w0xcOdxmdhRDtXIZm/0oq1GvWZREa2r87yXWHaU
TXBzQUQaw7Oj5a0giZKFPc1XhZd0b7XsnFl1gN+pY8zsaavN1u2XbeZK+IgQxd6Ntaj4+h7NQcc1
094L2MLHSrsT+PIekPUXW2AT7KAI0kfv5Eq31ZTmODXfovZG0CzgUvmascSFuSLBYDi6ujwa/4qO
BWtebZh9t/qEAKeYOvrfletV3VwuIRGQfoNDM9EdjQvP3fv6sCV5Anx+j3Bsuqyysn8vHEzbfi61
4Sq3yoVCWYFHj9u7g2PR1cxYeOjT2cZuehTn5pCq6Me+XcP+LU1Z5SunSfe7UbsiXJK8p1r6tgVK
eyTIi1bM/ekhLzXh/fPM3zJIcdWFTJ7AkXYCIczArYj10E5xwKl6Pe5LXaWI92uU8dp+++e0BuA3
q6J7dR2PMnlF5M8MDjrOCmQWyfNCSUqY6gbeuZlVDFQDBdsJil6cUsTnfXpFvAIHpkKHaYveH2Z5
2/tOYTkDJJpO8vWd/r1UuNhLZDnbirrVPqUieUtVWTZmSLVFS7cGB3Zh96yV9oahGtsgSG0KDkxW
dRCSNhfT8Eej6rdxJPuy8BYcFG5/0BZs6xgWdY9L/VKhmUTe25EaK1hyX5LKm/KG85gkOMYtCfaI
lhhvPgYfclLvNTXMwy44s+Wj2+VKxhVLxHwDwyCUvaA2ie+X++xPm5aS0recaVfEaW04W3BJDI2h
CtJb5L6vwYVMbjvIeEDE/kdtEICV4GQ3bq8xjOCdyAI/ox9z6ct5k1AS3e1MBDQzS8Ze43UDj8Ed
UXlLTUc9vN97nNcUm7/JDSGPdy5VwvOfVlSNSHw5SmXfL/JHZ+b/dr7H8wbWFmWslpPi8BadTS1K
P3Nd0kHb1041dCwvGtcNf+hJsKJKtH/R37tt8yqpLW4TTnHAmKzMpx7VKWqeCcIxFsSPs0t+BACF
f4ryUJ4HQv0ysUktFswNPqCswo/wBJ0FxA4iYZ7c7HISjgxPtJule9D9+cSgmeiFXcoWcZfhw8dN
+7XswT8V/q4RaYk5tXL+7MEXgIw7GAQZ0nqcJzw21g4kxIwxJjb7gXqe6QX5phvTs/VsR9Y/irpX
yKWvsl3b+rhVYPpoNzHGmezNkV1MDn4Yi37sFa7HPDCo+79PWsmvf+JZlNDb4IlnDgKkrgCb1cZS
TE/QumPB7ihazIjLbu7dydv6lxxu2Jl2Klgik5iA+j7PoOk6DuFUrwnl6WGlLN+xDWhpUDhndyXN
iE8WoHnzlrYmVsIu69jqouVwKTIHmgyTEZvYOKv/8Qrvd5hWsMqrkuoLgiWyOUKNz5Ro+AlcIzft
BxLkkqcAqZi3+T7gTYxV+ZneL/hXBccaKgkOx+8CnM7cJUxO5HtVK/PFQ8aphTceWDtJdCDYreXM
rWp+yfQ2ruXo1sBTf11Xm0oKAUXhgWB9eyNi62GfLGujyQGU92umhQwZjRlTEtkxGXdVdf+H3cS5
53VWd2qTbf9YMf+ZRZvfgKO7CumDvY3ymR2WPj+E/43GEneUfTfUkXhMK1Venj7e9aMJak7vFetY
224hGEHoFwGqdwoSwZ7rQY7lV3B1dc1GMBxpBFaMGlez5YWuVIkwfQ337owcW3+mXFBHMSKb/w0Y
DSonUfz/qU/47pzZOIV38kuGiiVHHWMKS2jajTfzLxOIlwi2sOrWOsGJfKKheUtUrnK0xbdCWIPk
g4K3ZlJWDXl2dhggxqs00ZyKMMxT5xoHSHOqio7h48qptzeuQWpOhGj3wJCg4B9vgLkkFLOtdANI
MVIxYNcvSM+7+bMWipYenCAksvUotsMdoZ0M7G4nJodp/NL+aBAXkdg1vkMQxkdlS5v+5iXfHgez
9+uHw4GuZtLf/ooEmYtGpR2o2H9jNlg4ObH9n6qlGsixqVWOW/JoFU+7JCq9IY01eKSnZXQV+cb9
y5uC+zZh4Ng5pZ6YaQDfMEsX9oHsUT/MMHGhYlW6xirvObfhcHoTI9SgaNQqwXyl+eApMv3ZYvEi
0IkgWrz5Vi3ONEDOr8cYzPkNVZicH06Tzp2uwwqR1BnmsaFU5yLixQJ6yOGcVtsbtSQSKD3O6t7F
lE2d+yz9CXicFZM9xh1Y4kuky5S2KpWYRYLSJnWBjn/AXQmgTyFODz51XODGZpWQ3QgQ/NR85p8y
W5iS4+XdJDoqPXK01tnPTgVm3sxW2UvxtJ+rAtkCFRE59pXC9IM9nFT6fJ5LGxmaoCTHI1RNfPfR
B4exhfT3ijZOUJPgcWTE1G7st5bvu/vP+33FEwl+Z8UFkiMVZ1PbhLd0nwXDtm38oV5AErc4Zg5j
RGBw1ZumFzMntPHpsZHyvj63DAWXl0n3LasBPxOvqzVBdkiIxWG4TSmFMasG8s0d1qYZAKjHp/m5
KHmxR9JSrBmcRdin90LA/aD4EKwIPsKlz5N5Rmf0Jc+AJTHvSiYEU0pMzcRnAqzhko4Zo4gFEmLw
OlMcw7XdnbnYb4gSvzfvphr/vAzC6mzdM0QxH6lIHz2ujNfBHf2P+BM5VpOEPyUnOSvUCFJ3UB6l
95IQfLmnV+BdxAF6jnsO3zDa7Vrln3AdvK6fbDoD5xP/b5At65V+frxHHyJc+SZcOCfpF90Iq4jB
aOsyazefw/SKvPHThNGYa46wD5sGjenfHFYlKdXG9wMglDOyOfkMH5DGb5cdSYyRg3Cp6/EcYzEg
77Qrwqb5ppg9MUZ5PaLzEtNY2NajP5U+IMHKGT+hQ2bYvW4tRyjsezRLoCFr6V7NHyhmeS7AbqSK
ApDV9hp64a/H4p6SorRXlN/ApQov/7hNGsVy3fuSPSBIsRG4k0PVT0Ar4y/dNRp/kXtx4VoXsJhY
utNHiHuJtz65Brhriq9Zy57HFP8KjiXxdfN84JvK56ehpEm0WK8aP0f3LqRMeRsdYduHcJ6+slhH
Mc5gHd64SPvxkeEZDJgG/lvxTN6vbOHIGeCAN3XqVIAbUQMBji6U/83fgvN9xys/wH8S4fZBeEVQ
cnrrUw+btVt0RCPoKyC4LKQQIB031LIiCnc5kmb9LIAEH4axY2LVGqr/qcPF069r4pyhAEc8/BVd
1RIf3gi7dFYZCFfAFPuQbCEQW+vVuEOjRPz8FECHqEcPhqMBJNoO+VvMVGvhR1vj07dEVBDl6RVd
y6ufTGnWEsUJQ5bll8GzXe7umUqMOmvNPauezReczfUJu+tytS5mQWWjIJ9XPu4R07HA0lYx8TYq
NhUGgD55LK3QAwPl91vBXoNxcZ2e9DcvoW9wqoRDH9CdVEq9FcXBJoRGoCfserSqLF0CyOcL3/BG
GIrt/9CVMkJ2D7+PRiHHdPyNcGgl3WvCtgDY5JjiBTtrNcGnUIpr3Oss8FO/SwugEZhLkILofwGW
qoXHrSHlPn73TTxBagovsDf4BzqzF0KrJVIRgbeiMDEfhXmNzJKuyhH6vF1LO8hPnitE6U165yI3
uYMyEnZq2AuPmI7H5lBv4lU815zQ4DUSy2/OMw9J91ylqXA82DydVSUju5ELGGAbyKVsbHiotZMf
IWfAVaNUwKy7JbSmYrlJP8mXk70/uvsDVeKArJqRpiQ6yMfQk8CKYl7qJK2QUmixwFtd7zaMT1L3
U/A5QX6dHvuZ6amqyIYu5eNSBefpQQ9seBz8c2blXN44NZ4cHGD6sPRXN5qoSd7zaECfliDL1Q4Q
hxpaptrwYaEDkieKJuZ39KO8NGbYQEsCOXwG2Il0zNtDrAqFyvwN+iv5+Tgn5FSwcUVj8ZF1ItWj
d91ASbPtgpGge8hUm323+Hp1CPRiXTPKnn1awypjNAWZ2n88kip9nFndF+uvXv+kJoPrbJCa2IPv
ZrTWIHP9YdZs8drd1DqUrTTumMdnx7SLUmv4LgNGQBoAIZ4damfIWkztZsVPhSdmD8ckRhStbfkz
FVY3cSsQIOFbiOFSnd5O/9V94mH7U+MKebgQV/zRc04j1lI/JS16pY8KW+tuoIMNyPRCBHVAOOAA
8RcRkBfd3qc9kpr7C8T8R+ae/PgDTPo+h5E4x+1vtYD0L+vVB6FJa/Ccvs1ez70HVbcBIYK8GmVy
kh7Y5WyjSrXeJN9VTLO//XaJqj41+iHgP4vHVMI4sdifBY9ZDSdNSZrnoADSFZLNbZDljAfFG/Br
sr8OvvUp9BvHCKnfnh/6+ZOjt3oVoL1cf0W8QCA+auAOJjQ2rrHDCzi3bKsNiRz88so6MnY7t/f7
7DUOiVFJADtbCNY42NJgtzbQBjwzm9MYhQDjxkinm3hVQG9AzpvwKxvK4fgXVvAvLsFQZf0YOPrB
WqdPqvTQdLDN9kFdEzwhu+DqELhofv7vEKvYNnPvda9HEeQUAqQ1Hd8VgPJpWu0Jduv8T9PdLMym
Si3iTeB5lTcnn9sgQQ41i5Yat0VPOn4Cc5+gSf5T0PF+DeL+PXFmZxSqovMSW94bh/7HWw7HhvpZ
zjJ713rfLEdiTq6o9U3uZFZOOhMMfkKnx9RG9AuEYWiPvgCTLlqO8xqOQzDdJs/uPmb8xsH2MBT+
4HDOmQWh8ORPrd+YEcuNkQ2IdZekei7gZBKLxXOPZj8GVBYsxCr4Y88ZLQeDWLRDJjVN8TyMteOj
izcboP/Dwkdx1qkugNndf6G+MzU4IBnqrR6i60ag7RCzYn0U4FvDQGlFDbfmj5dWFLfk7BAgtXav
Q7IqtHOZWuBscZoloF6HTeqmHYCY9iicYAas+tZTFC7l8WGNy+MFaXn1+flTB5DjDdRRkJjyjues
jnQOgBVfwIOf/Hn3tj98xYbN+j0ajD/mr71Ghrxs4C9cCmSN0SVXTOWSrFthoHZDnFOzInkkOECS
4mzRTLlgHTBGCZKNpZjntrQEg9jmLj5O/PMzFBAHuehal2XEmHtRVFndlC5ipK5NrT4ziyWSlA2R
UL/ln3barlVjthD7tpwTTk/SFQwLaVIqbRtpmTDAbNrjxa+hPxyprOnDGd0Fq/qYypoBGDjioO2+
6yfq8TfSIeqZ9MU4XGtbpLb2WhN89GNPZzvchWeUJyT7okQTBL+/lJPnCX+0GhU28liT+zZHY4H/
jcADqgITQKCg8SVAERgpWCnP+e4LEpvvETeqmLtwoKrpoPiKTFoitgdaNu/UJ966ZZkizMnNTyap
5f3I1N841+nr7R4slG/ECseCip9OPS4n37rFvB+ac9m/djjGy4BX63TRZVwe3h8EDCdjhLzfK+IL
YQ8G8UZuZCQWMuu1MX6HRnKz0dsCNQ1biiVfw9XsC9RoBT1D5unrap4SMbF55/hgP9WYos3G5za/
/v2fm9eDkVCyRg9cPr+cPTKtNDxZ/h2BLHhBEt7ZGwiLpH7tPdM6TxhFdUm2m4/3BX65q4RIkfwg
5sKlERZMiHCDAms/VWHepcuEKoXXvSc39vqeJYPyPtx9RF6EddC2D8z5JPVdntMGQ1QKI1S6dAcD
bVKA3VYZhdt+Aqu9VhqOQkuvOJQZ+va8Zpx5Sa0UNF7fMmj7qCAxCiU1m2VVUD1adocCT8Yw/MMO
LAgiLNdcbRAKtRYx9xuOH6PRPa9bGWnCuXx4wHfoZGIxhjcuKeb/kSByTgMLhdVpqWTswwXhllkB
Ic8dBsRS1cs3bwYVyy7Taa9wQg4tu+xk1HFY69lj+9pKJw/8E3/0I4tnP3QqNlpLZ73AfxWk4tdr
rVpBb8Eie5ye3usjP80XbZZ+hgJj4vKarmFLYiNEI2FAspcVrvSNVOj90KUSe4NNN+TQy7XXD+p3
4InfHEmEpce5FkuX29wpkjqrG3aB+paMnyNvFZG15IE2AERBjktrEkZEB3ah3YKNzkjmz+Ds5Y2i
q9gwRWvgb96x37y5fnDLKKND2xlAnikkMQkEePS/zUmy0IM9GqsrOzFltMfRxWaGgTt1IA6Zx/xP
O9u5piJ91CpHJU8apckz6GJfpbRW5l5xfAwZVLuEfxvmEoFV0JiaC5QUZukUA3IzaPfwcIeYyx8t
mGar86h1eU+5yhJHlfw99rXFqdEJhaTcIFmQKbQfhTgsqly8L3xfVF5CXrjQwTuvUUKQJP9vE+sB
+9QuTDOMM5e+1iNUN9Ot5Y1mq590tvzbjBkzAXLpvFFsEu2ejNi4GmgOYArHVFZ0gbXZ8V4f65YS
KZnm8+dZ3vqw68QU2BhenHBQtnF7pbZzdMDIVS1G6LNR162vYhq97Yu6dlWXBeSBPPnny805EXwc
/Ij5khJuJ1FDVOSNs1ww9wpKENqSbMgoSOWbXOlCh1GOrEmoI8TGH2zlYpgLe3X9hXR2UM91i6lP
gJ1fnz/FJnROCtzI3WCFGS26EOMqDOncVKUv2Gy4jT0wxKma95jsI2MG7ys+LLvqqY4c7onORbbK
MKewCGjlS0KopZs//Cpt4bVdhtWv9guUeLybBCtr534alePfA6C0/oj1htwON7KTZgPmcmsd38b9
qSV02/zF39yciOj2C8r9o/GCQwn+tFOFiwn60Z+m+JjngXJvq9orEiyI/ubiNsRfeIqen5i4XjrU
qEfQQMXzkmKAV3dcliPO/HqTOgg6wkoRwX+mML3IXAC1O7x4xA+amWcs0vBjNQWxZaZZh/E6eSBk
oDHRXxKXiSRNikHT0mI7E/lT39EsvTlC54jOVn6AJBNlKQeFNJ3G/6MpTabiTY33yDkLZy7cjHND
ty04wZw7gWOIWXpFpFgvfWsm/0xogfYYtYzLypsFDYm8HPah5QEhrBBPLgOOhIo3cgV9f4mUbufZ
a7alhnDIqmMnlSerWojVDfL1X42mw0w0tCtHZVMd8O95F9/Q9Q3GiyGgL/TyDHfYuv6rIi66YjKG
c1scJU8rmAWwZgcIYjw8X6tpqlrEwRFrMEpV5B235h5/DxJeT5k4JGnAHzw12WORg5mNPIB2wCbj
IgXTChlA8cOdAK2NmfzmtKK+0qpWK9DCwj6TsoDklIoqdt/wlUossQ0xolJtaSPtkC+kgsRkJzSA
0xxklpEqL57B5lPCXEW2dg==
`protect end_protected

