

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZF7Gp+JQYN4x6Hvjz/p/glt8+Yhfw+y+NSJwSgFAT75FGfBEoCi9gxGC1aPKEYH1nKSH9HDVBmjN
jVYDQh69UA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bCrwACZO6VlyUjDp7F6NflPANkTfGVm4hgH/4AFvgK6LtR4U73r1HOWXfaKa3y3uaefm3opyWNhK
nV2TI2PpMLr9LswzFSOsgRzHCqR+XBS+8LwZ+lBVN3PhbED4ykAJBbHjWQapS4mEVXs8Bors5GDK
A5lW6VBcepABjdMHcOc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sWMXC7ertaTFiCso7MQnbVyuVSvzDQRw1zbA8jCBUoJcGFv+Da5uM/ZInIx2vKnorpctjF+RfQ/I
vLvHJ4hFA7ai3KLDBa+osiqXeR3vvyAO0dNGGmO7GQ1dYRUzzSKKrGTJhKWqDfnAsYaLroy6U3UI
uNSRIQtxv1ciGPzcMfrykPy27NH2CEGiCobfxP5HXDyrOVBqWAZuLaPzQRv0D8Ie2O70SiCDKawR
vbedGBup6qqgOpbOuoCX/zcbW+qJ2FxQY5Zrju+0WyLSf0XnZd4src68n6rXZlziL4eo4Q6lUGQv
gUEyqpp9Wiyw0QLmYTxtAKnwwMsfY/jCo5ZFSQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d4cZTzaonF13oHTIDZgb2oXxuKQXQmTrHOYXqYqbAU6BYAx+7y9fxq+NNlLqPYeukSU316ZJ2R63
uH6wrMfXFW1V94ov6Pl2EeLSPre3P4xtwdLCKbJrudZD4i07Cl6ICwNSN//h6MJD/kwUIU4k7zeP
ni9WJs+GmLVsVx0bOck=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W5Ic6b6KWpsR2htHXte3+6CjlmHZcuEa6WOajuu7k286E/JIlKxSU0tNrXH7rL8k7QTBc55tiAC2
sT6Jtn2FOqn9b4N96SwTUIbdNrh5Ew/7EjwCsd26VOwpEgD86kAwm7rEEtRCtStJR4p0yrbCQjf+
9+YuvQ3Ab1Y5fgtY5ijqZPgs+knlZZFAxm+NI7o8f97lEMTpHDonVgfj/KtK8xhV46JSrDB2FPhp
PMezRFDPcrnrGio0JnUe1oPbSneaSJZPAFIoGiaaxfjjDJIOa0DMtbVjecaL42P3+sAmOk0R5Mfk
8MlmwedAmXWwr0D9NdqrNJ68Zt9aVa7CXXiS/Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7632)
`protect data_block
JJ7UDLdP6VbnIwe+mB5gQuWhChi3mtm/4IQARy5zGFAOy0U+rY8czeoOJs23iHWE5cpAvea20X5x
hOamD+qcm33SCvE5jEeDDogvTHZlStg6lBMHpP+Cf1S10mUyZRxv8CRMNI5CR5eP+kTrLIhB29A8
2EaiN2q7FYxmvU2BWrrSIZ6nbsffwzifkUqGB1wY6aTbe4v3tAe9eKshADkcNavxPrR+Q4hwH/zH
9eoENaaxV8BtzTvNx7DkqTpDn4zz+9qENthYeWfgrVvvme9YrJPS9PBW8EtDLc2APJNCabxXYb1I
aQgYwMODShtIjqGWydwlIjzH6fHhbom2eESKBDDzNuPXVTbyAOkNvy7o5Jhxxj3EgUsNKPf9bUk2
T2yOBKx7Bl1Ex+lMVj546bY6xJ+0xSzcesQcl7dZAPw3JK2Jzfwm71A0GCuxhYVT1kHBJFAvw+y0
YPGoRQqi8s/sWq1t6HCkk1P7rzujIE78kFonftsEr+5ar2nN2I976gjDOk0RdwVbd3M8smuaWkoL
gkfo7fEe70WlYSAYLpHGBwCs5EdEJ7drVzA7BgmJZUTaFUrBS6qdDpQUVz9tRkH4GDPcRJXXfcYL
Izsi4Xs13akqcviJfets00FAol+rxe3U0b4jFu3BkLSlkAvPUamF6Yv5nJIMZg7OvJ6iRf542FL6
IVS0rcNsihipbmoNKScBkT3EMf3KuD/2crO+2liZxg8jfN0CEAQ2MsbJsJHRxqxjeZTgCAI8bj/q
lhKEc4O0sUux2Lcd4U/O3rZFS7BFWkXN+1t8IEkbYtTQdEjneFkz9RsAz/9fL8ixpNx1TpslJHoK
A/gZY2cuQTNIb0JlKlZlQg0b6WulGEL80lP21j4bKUSjah+n/2cykLWgWax/bcgoiHHVlcN6HV//
OnOGoEVLDYV9fZG/G9c5ev8yXyYs3PdcxIXjhvZsBBJiNey6N4oSNsnM+hYuxFGzORD/dqTAl4yT
BNJc81KxHwo1vXT5hInzt4ghnTGDCZF4Qxzer9nLT+qDGnVMg8/uHg1EaPdZxGCpTQNFNGKA4cCj
93iN/15cveaEkaouVXAzl0vYGZD2w0/dA4gulxjJLuT8wn+wYO4U/8ZTdZ9QckaB41f3mJu/rEkz
pZCruF0fCM+1KpMZPOHupl14+mnAoCaLCu3g4Rc1unCAN7IsrIO1fvO431hhxn8NjwtO1Ct867ox
S6s9u9+K5IEdq+3YJuMqCbanjnuoW3u2Y1yLSCH+xQ+novlgWMp0+rcK2X4RrC7NhtU2ZleSg+3b
J1AkRVK9q/sw0bpxeqEYIXrnfgQ9SIa3Z9uGYsdtaSsfFAwci94zOuLKcUfqMSCScI2lGKgG19ZG
VHxiusTXGO1CBHZIBXvSllkW0wivIwEAWplW+iRbwHpXTAPlsQI32LttulQD80Xt+tKZI7uZdjbJ
c8BfhlQhc2gl8w+2EELkEX33qYvhCkSz5wrvTSjTOUMm4VNTMlrFyhuBfHB5WyRMaH6BXIlZtg1t
zDGPD3gHPpPf5aAT/hFK10le3SVg4M/pbVww0KMWj1qvDLzVGTMjOPnpTedfCaxCzczDwl++mGlp
thIrx0JZPnOdtnfnl/DBT8X7+Nb4zJwNnUF7jyN67OtNn6aBkFmXH+BTmVwokXivbxdmm97k8VCv
55xCG7AqMIjrKU2CSHfwAAW5J/gu+lkPDK0/9oLk1HZvvtemkN5vsJyt6jSg1nWc8D9TtDj3pZ/I
Zci4Rq6t+8da47GCkCWFUJcTifUQFojiIE58J46yXC79WUE/kpiiPMcBRIvsCELk5JEdcvE82nJf
1raddiSlNMezsYkuBy/uEnwva83AUVKncFTC5lLRD+AcdmabPPRBfAAq5zfN/hI75VHTCHDFslOh
VVXT84PQ4YdXwqSGV0Jrq0/JxUWEoLXqNX5lsjahsuvx+SWF1xXc1k33584SiITrq5QYfLl9WTiE
kY70r+pM2Zz4UtBOz+VUJlcqpjX6sK7nRlB2O4dSXJo3rnDYB06u4dn9QYiXYqSiHgkLEW27O25K
z7XaY/QJ2z6PoWABGHANC28Rz5SdIOCaymGPuqGwESkeKtMbIA0opWg9Ztcaoz4P0gaol8ZeBmzs
EoEH2LmgiIlH4hWGmzzjls06DsK1OIIA6MfQvtdSrh3GG/XtCScg7W05iR7XrCqj8AfYiAxs7fIW
xQWVld9BFOFRNaPrN+ZB4G9PKGrkrKpZMZadCrKOqZ4efBmY66uWs29hWKjEEf+yreLxtzeD3zdl
Lp1Ra9tYyLTGk6hq0SPDClihEG7Yp/nwifu3N0+uFoiFwbJSEl6e6ZFFZDcOiwFJd+7DNQdLnvCV
W5fpaboiCQUHFJ0soj143Y2r0IhaeN3/pXRkLCWFrRNHLE2EXw0ggOOX+hh/9ldRSDpeAYBRE08m
Zh4jlLDO1nHPhu5N9bY59JAJv6XZfoa1D8eSVD9sh7D3oGsLTrIumArqCG/0Bgo5W1QsNBguPhX/
Jg29GvVI4Ox0Waolt968p/muhelYgqR+mrjOJgIIv4nkqlsgyh3Jvk6Du75+fsk9e2Ke/x2UEVqf
eAIJB7dd/Kbz7zar4np57xSqh3GE42MiFnyTiAMifG8ISTAgV9InY/C9XoMkR2lBHl3O1OCnX4wH
doUhtWG7Ljbzrlqysygd+E0wuJuFnShIupBmQWn/lloaTHxHGkqxcCfxiOkAYnPXgMrp8eHgV17j
CzVRs2SZALDuxhc7buYCMlDisnW8qYfSM6plOFvaZhCwzikCqfk2ni1R9E1jIeYRTYd1UstIHWmC
9BDKLlgkLDh1kqRBZt/aR7iU3zEcMKWVd5oOgmQU9suU6qP/kCWaFv2T9oMBzGgSrd/Jd+UZt6XT
LtcCqZFLzMfGnrOnqXaRv1ZpeVhCFsCnebT2jzqGfx8qdCRTo2wtb8wpqdFqBpveNxdFAKRmpowh
XICkTi9uA54yU1Xy+xSWKRROr+Gbx0fKdE7I1Uqv62+O/NXAj01GE/7kayW930xX0lmd5pZ8iFn7
iHyeWT6WrRnz4z5BHjLdS5lhYNNRUUgp5zWBfMD5lxnGVonFeN0PZHcVKLz8jYBhlB0QtN6FWQy3
sBOhKRmQ3rEGaA/AuYnczN5RBUGVr9jSplOjRUIzk58dW5Ey87G/apLdf75ZRCxPQOPyuYyEsjvC
UE/utyzJF6YCn/qZFThjXzWXN74g2Lt5IGS5HhIJrhg17C2qhy65c2y01btsVDJNHei2cjhyY6GI
IWUZMWADlWLOdHMuuYBl6dmxfSvcYose/fnSGZNUFaLjeF+bK7Sy3QAbCqv/9AQ+GsYxpAWoTkOO
vC/0uncAD4fmfzpSMGmowMzeElbVUEVH9J69jL+p185s351Lbl5ToVOOqtca+MQoL2weCNiXH1n8
mzJM2mJhdLoWsPl5YrCkX1JK6W4BZP5gX5Sec2T8LgSTIOVu+FvX6uYLUSCz64yFp5wAnQUFEjA1
XkDFOePLhp0y5R8vfPW/q48gli1sgGX5BHHN78X2fR4bRPrJh79Wz+Whs8hj3Ia0t1XQGONI/zIH
9Wd2at4q4v9gYdxo7pp2hQtCQGo14LarM3zjzKTJVzMsrGjTJsvoMPMuKrrMJiK0/hCKxx/QhZsf
7NJXaHwYT+0ShmRfl1IDNeSIRAaZDCoYSy/KhJSHiYKxZn5kqMJhSL2S2P0AqYi+gNrZLp3Ipsfv
1hjTjkpWGnopRYooiK4oDaA/kDAvrjoFjmWegWq9ZWNGtbjLoIVVvoIUjkk208q1cJbuNJ1NrdyO
6flSXLBv/NuXp92l/oANFQshzp+DMX+OZjIqGL01VzULtZ0JW4SeLFlWBS0x4pCLJiow9uWGh1iH
HujQLpoT5a0xzk5xHvEbfRj4GtZXVqwlOLkQMDX8A9vsISfQUo2OJZMfMFfKSwZwofvYWqmEEth7
hj17DBpku69DBKEjF6zi8wUZXIUlB5H2YuZhJqMc8GYSojU0MPZn97uoGw0IE+a9FcNAJBWwt6z+
H7Ct02O7TrzGnMsx8W+7Qc9AA4Ypa/bUYxgQ+qvxRNr7zIJn4iBtc81MKQ9JD1toqGvA50UktDbT
AJBFTcVqaclRxO3jEmDgM9zFcIi9hC+9qpdP3yNmlVj4ZzrKY13IhyPK7b4o7cuCGlzhoWE1gMQQ
zxJdCYTlLL8o+1zH3PJRk3sOT77QpgTMxntDXA7URMfp0pvPfSgrWtxi93PL8VaubnabN47FRgzD
TsVu5e9xviAjczeJKhd+JWYHdLvRi4213ZlWA+v9pYYDrY7SVu4uDJbkLAwP0hKqD3hdGuccfLGJ
nJUCco5IuGhszZ3HHVxlTlu+f2Dj9pHJU/6qvnNTOx7w7Ik4qYUmIFobpB/7BYdBOCwizGavR19x
dKGJsOgQZEUeUhSKLPAf9+6xpb7L2fMOWHwmtwn/VsH9nmzuWqpOQ62JdfKL1yArAypj5tw11CoH
rHDVal+BiDNEfEN0zDf5tPes4hVAHSNIXwFJyeMOqqs5IoJuq2taFd8zMggoqaXm1N1hQonnfFu6
tm6De+MhnJry/mdX2hx1qh+eTPl33L7cNoQiTQG7RzuRg4M3+lfzW5rsBT40w9s9sdJjJ7UBfyLD
8jM+dh2YTt5Q3X70JsBF31esqOnM1+wng9l/gGDUdOjFkF81CzD62MJtIgtskwI+1BH7jC+G6D05
30u+Pdz9Q+Z4PF96+dhWpv610oeblFw4WhwUaQ+fk3VtcqBJY7dNk0NxAXxHTkeqD5Clm+roDUMV
CNankZ5Yv0gWidxZBojOFcHYdlIfaO7viKinR+ED0GLthiKE9ifcmjJ7wsIYA7PSSrGLNf3n3Asd
C85/L/LL1vJDibLvVgzrFgiGu/qBo22GFHl7aYIVPz/zQynd4aqvxoRXD/1MzXfmO5etH7PK0RF3
KY17SAHxvrrFAMitbtk6iPR2JKtbTX68JwG9RIzBrlu6sXqCd5i9WPh1F0aDVpe4am0yA8GidYhZ
s+QYVigKV+OSh++bpge+SUvib4UR3Y4U/2CikTEqAFIKjIyJxn2NlC/vhgUH5ztTAXj2npLhbnNh
Hx5ji7T8rT7C+XuD0bfyBw1BGu4oVJVFgAfhIO6V0GPm0FrIHCA7L45bk0QiIvCMrUH02mRsf0G3
8bMWpgRF+CjpIl2Z7pjWuy9yPCfpVha35xEFS/Oor+7l5e0lzsFEvism8C0dv27lzu3qrs9GFmrd
AYrGcT3YskgeDOx0YY6rKdZy2i8qKd5pCwCTRp17rMidi5tjzbOqfPjkgaKTqtAtIPFfPH04xT9Y
YpxprNPT9deZ/SFIl3oj7msxJH6li9wlVdcH1NwDIAPhcTGj9A/b8p7xcEUdMoLBGuko9NujJKYk
H0dm/7JvZQV4u5G1BRVdd6TqEI2dwxATPREfvKc+JzwQbmuEg/Wt1OMgwNjiOe7JGVG7MPyLIWtM
L3WJlmASQ2jfxIgs+NhdBOshX5Xh58yCeWIegZGr7rCDZYeMxpdomYYKwD2/VJaJchXbOxWPwELL
cQVTbbMl9cck/wokbgBLi9ImK/drDU1sWCvwxgHGCRIl93vd7pFlSF2sSAnjsyiquUf20DJ08M9x
zX7t0bZ4X2ucQQ3ARP3/qcE/kW2YGKjVIdEQiKAkLn87SVoKEHVd97gOPk5u7rUFTjeE+3SInE+I
pbCKi97cJXNat66U6XCLiHtJArfB9BCrRVxC9Qrhn9MRRTLxDspRc2Dfc5ORXY9vy0EfWqLHppQ3
ZEc7T7opAw2taq9tm1b1TTNxiSsLb5fQ3mIIHTBcKv1vmWnh3HQ6tbXn2ywwe9AtJnYUlnA1Eic1
pvCDivT+Rjalakd3xBHjbgOTAM+J7FaZIAtbf0q+hKp28ovXZnGNhm6Ky6s7FyTHHVXmuf+f0J6B
IhYFtE1McBNriN7UIQFfSve0DTb+5RonP1nAln84cvECNn9N6+9gvGX6kTGZuS7lS/tgNNRrg/SD
elyVp0DDPDS0cKImwc6R5CwmQqgzunLnZdpn8bSOxtBumNg1lbY4cBtwX2J7kGeI64+EZkbrWMqk
ua6Mb1IHDGJql7ee2eY3l4ysrkaAN5wH24EqNkeP5E6JXoODO1afGNLYBM9LXy+HF2LvAxqchWVC
CLIFzzd6ww7bCCRCDyEhudMNbxtIuPEmpjDR2oT1rlQVHtnQYHMzrf9ZY+nN7IGiXqwM1fMjKyHh
eNhueyRZOHO9dv5+4SLwzcw5A4zeBRP2AchswKCRi/Uds6BZH03nKXfwXXx7hq0Y32XvwwoYq5bq
6g+jsUWmMcvsQ4HAv7HGMEB4kDVgLfpeHq2X9IUUFPC+TGXujceHo70Ik7FO8IeoYA2dpQ5nkDjW
Vm4NO25EcUsykYota4E95PeP8IntXJHKRNb4EEJtTUg8v+Fy+s9/ywdGwKVq1QEOzyzKA6JpHJ6m
KwCHnLy1q5oiMPqUBMmVJPVo/eQPV2LZHzuZLdntdTFRTcCW0Cs/XhX7SBdf30qwb4Jz2jpoV74C
6QLHDQCPQzXo4swbj9DIiw2sRqCFOj5LENXTSA9FflP67B54mER0g2SeRP/cghgVQV4rsq0jNpbR
piDWWGSMPcSmp8775ygLGkZbr8BERMkEUVBvZlQ7pkgv8biy6CkKz26xtrMIq4XssCB/Qiz16eml
m6sSOBYq8v0OquHiWhV2SXtrAtkMuU1/Tm1Z+bc2b8Z8nYNchwJf6oG/Cyk1mJk1yDfFVfwiHII+
wp3+nwpm+JubU2Gq35XwtNDSsLISXC/ESG6AZOajtJjmZcg84OP+vZdi3UYWA8Irg88OYj1bhqCQ
cHgXp2r7lCiysbFty1pxy7HczIXQiyMXgaKYWMMFi5PSxVPQHSPzcmkxkN3kMJm8e2HcpI5ArMsq
5UwmvP4jWVbVuevDM1cIV11N2ohj/7wffeUNb8IcyddsTp6zFxpdVWtJQ9YFwhn60URNvvu7+QkR
I4a1KLQb3D5/dpdt/BPoCHf5Juw1hcrF+nsB3ML1EFnOMHLBRuXlikpaoiljWxXki9ofEHSekyGj
LqgyE9PQjPVmRzbMK9WFTq8VnyyLLWBkZtJn+parbhNkLQhJWLsOsmctOqJATgruYCXcK7GMcIqR
PX6uKo5XG+K2ohhCTbLqQxvn6flGwK6QHI8J/15QWcVv3iyoDWBRg8+7K5SswSQm+9MH1Cm2Oeg/
Gyzi+1UZ+1eBydDeCl886xGUIo6ETA4kyE3ln763gENPUsxmWLqwgcAuJYyc01Jw6T2FPTNuGkMg
H6bXqtYoHKOFyx/J/T/foFtgKxwQ5TL8DMfI7eRLfguyW6PHcSRB31uhvi+fwPrjt7m4X/WD2uv4
y7oKfEVNyLGYP6tZS0ezU/HjuZ1xH1FNuKObFtC/Wl2LFNSNvyncSJBKM4+tStOFWv4jDtkNC5mv
xs/3O47PXgjcBKCPFzBI7e7APK1RTQq8k5K40Q5XgfXR+9bcBGjp+xDwmJ9LmX3R58mNvi02B9AW
+qIH9NLQiOMAykXKRGwgmd7exkFFDSGBZXGewLxVjjYSKMBNv6/5kf35wjmSrFAkKZ8XMt+4grhU
gEy2TRBk7rnfMbgg6XMPl11rwJJZdjHDswxc0KTS95mtmATjHBpXMR+DGQRGQH21sIawinLmh32l
afJJMu/MWyIkK3maBkCu2AWn61g2+sFBL5pdzGtZ4I8DWcbnWG2d1kAoFPKLarZUmGs0Zh1C/vGp
Wsclxn2vEWCuaIr30/8ZXw18AOCuJIMtDWJu/mkRSdhe3hDo1Yq+KZlVPKZ6LAKbQafZzSwLXQPe
PZCUW0uruDkTSKr+DldzNmBWLbNKty9D6v0/iITJMuayl2A+fbPbgG6TpzqWraSXdpEh5dnNbjig
XtsVoz1zdr/nC04a7IL3q/VkNWp8trbAFmDpB08VaAULCXLQNaFVWnXMlmr9u8JVweqi5MI59VKl
YsfAo+BqzIWRg+CMdr/J31fmb06PfSzcmb8K+ls3ZuEeDlOWrU842vaRM/glYFS2sJfkCGvR5G60
fyWkQ4Mm27pBfx2JJtum5oHTkLw17fghLi09+g+jTIauGGOKJEAGmrCHxP18nBLlIFJ/WaB4ujh7
qOMgtAA3bPD8QoHY+DUQzUYQtLc+4zZ3WTVJel/Q0zXWH8DGxRYQA8P+8cnVmGgcy/Dmr33slZAx
Ds2lBMgDEWTPC/rgyuOx3SYfe5tDb+slWcbQ7zS+amPLtyyQ5sgTmnP0ClBfXO4YUIcdLCMAHrZK
ShnUC6vLS9nMttUVd8G45r5iXdy1hwaDykNGULyMVbT5y2ogZni28sd20KLHjRW0kFhfrab92Ibb
qtnTi76q7CtQhcKkrxWiKEwsSwv4E2Ke+dEdcQGKFoohbe7Qbhb6aNnT6ZaLsEW/uTLLaBS/EHPr
fu5JyMo30AHYlAedlVDa+NFNgqwxhVgSp/cE712o6VIpKzbaA74QjLRZS99AASVdmaJm4e24W2Rn
qFui/gpcV1eC30Fsv4RdSzeyPgkgJ9BwFj4qlCEMjOxqpz6NCnFa+GCC5yoAOdFp87zsr3JhuZaw
aCnbOsPDtGiNso+81/kD/YvSdw/uF1EPO0/sQYGC5aJK7G9I8gXqD70acuX+tFxDTuH17dl4fP8V
EUU6yBaWNvO8SRfY/xSHR9U4M0d0B/mULbQXRFpgL64jw/8sENVvE3NthtuQ8wqqGB1cyQwxEgH+
8Qak7iYBcTU0ENfSGxnn500ARxENWXRxGv8Fs98P1LVA8n82GX0oitUEd/cHmmjonDcmsUQlPU/K
QfcoRuoSY7WeDXz1HYoxwGdPtwFUvxRmzPbKwASyVOsODPoDhE3iWSDJOQcyXFIAF6T2TrXqrhS5
zdqMSJnUrZurLCznDw9Pe2x+SH8jhYAbsdbPu41ONSEWzM1KelnOjzqVTl2SG2tb/IHoSH9fjdvi
q3xBTopjLZLtP8tWwOOdxiR5qC3g8ZQuwv4Wy6qCmvBgg9DGR2/dGEm0lEk9B/T4CyOtAUkunp+Y
gcL7AFGEY4P06Ni55fOJaHlzlPWwJz/8ARi4McPOtJi0ZzszMxJlozGqosyp5iwuMByxyyQleFNT
H7ocDf4etk9E+aSJ0T/N2OG3QTJTnTBzFKWOp9/ZeO21zUDWNOpWVT2NVzLICkxqDu2xuvt0FQO+
0rzfUys5p19DZMe0YQ2qi/wWWi7mLvLL7VbkmolBimRtaIUa9sRbzvv655PUQfNr3ii2zB9WnNZJ
JfhqT3Gb4AlT1Gs07TuEL61VKt0ANtkxHsKXBMoXmpH+5HjSMNwo2pFD9tCxyJBL2LxXn/wZPrm6
zfMmrTWGnKWw1Asnk+WvMv3ia16Csl+nF+1C+V8hhB8+EwMUHMpAdIC1L8V3pqJy5YG/3n7a69Fl
jWtcHwyO04ALWI4het9+LKicmTV9tfXtbDIg114bPcEFG2JydzqQDcxHY/O8cCtgGdoPwR2KMZ+v
7qTvlrZYTQHmUSrMz33Rp7UtzHskl0L5djlEi+yl2xle7ELIQr5i/JnLR5qAJ4k6+D9uon9uCQ3z
jqMcDa0Uetz9S8L+PAzsWqDLl5rEWyXKMjt7HVQa3opx0E7l77oSWtLzuzpQQ2lnwE1er8vWxRSw
sEqZ76DG6WrZEqD27YFqo/K+Uc6jC20cHz8AB2A70h8fuFE1UFk8OH3nuz4VTVL2vSrt/pwW/+lT
1JqBQZo/VhcrNJIwzVAn2cn+KaxU4BHPYjXAGOOZq05FnzAL7M7kShYVCCuDMOeE3Uq0hfbFBge7
gsPNRSbgS3+Ar0r69QmPFa3C6LbWRhV036ujWvKxpE7DDk32d8l3KbTKUcm+8ZTIuP4GI3nHWI0Z
DgnBbxJReeG9wd02Lz4S2rTrqv3kfwwd13jmB5yyghSWKQ9mNtZqJP6+s+1zTgYs7qECWiNHg3ZX
Jh1a5L1HK842mq4+tqX3gzWyt3XxkIbcxbVpAG3QlbCRiqw2+ts1Z5Pj39OYAjAXm7muPuC60tjG
VZQvmDlIMUmUkj4uGc5qtvgEtUl/XG6cppUqmFhIZIvbiUXdsXzPb7gT4XQCzRiEL6JgBhNstwpn
oeog82Em5DnIA98DDjN8zN1COfJfpqB14X7G6FHKk0NubsHkf5r5ZylJIpUMMjoK6oJs
`protect end_protected

