

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CJc8rmbxQK7PiD9FE9h/V8z28Q2yjtwOLUGOHj92X0D4bGhAiTKxH6Gs6WbTk3x8dF6WKWHXW0Xd
imaqryWs/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KUGgnJN/sGLwh1pfD6BBRkJkdz3qYXsMmFAG0D8TIT3kvn1DM/WYFdJfNjuI3TZJ+GjJhgQt/TQj
vszszvccproNtKL+iK2kDAI+dODbmK/3dk8pZpjNIY8iqG+SZd4LOHkCbGnDn8J5L1SCb1FbgOpc
lYLzGKyKMfpMp2H5zrU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QPilQnlZ7SkqHJ+uQKxasOWlKPf9SmSQp0r8PPqOPGeQK2aUl+9gzicjiy17/DdQAM7rwf++nyUV
Yi5HrcGStcw9bK+k96zmiNT/NPvXPX5xeKvpNagObga/il62MarkWpibvt8B7D5IQi80Rp8/xMyy
QM6+TtOf7NVahw7dZAUwr3krfROulZTDfEY3oalO/PlnwAGr4Z3udXzac9NTOUWxkjpW4cmTbWcJ
unHhHJbyMO341XtwkTUgKReezgKFOpi+gREeBT80YOKcPQyjGyGuc28HYVmxKisVh5P7BYL5neLX
P5GVK+HA7MCB8DsbsorDqal6rxwDeaIF/kJcyg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZE3LPHWjt8FXIcLXD6pONgldgtzqHVcVbUx4Qj9ztf/3D9DwoYFB/m8dT7Cv2OabvKVMu13QC5lB
rxR5Jhd+fouVouDNKYwIESeS4DEkgnwfSJpsmeVaPW2tqCd21tzGTVfcw3Igam9PcTjnI1q1568h
X1Tcmu9paLkGRwvQeII=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EV5YorhH0risCTPPpyQGO+wsA9egdTVjrRAwQuEDG89jVsb2NsTih5Y+XoLrashGMO3AtQzajDhF
KB2YGM3JfNSzKu3jU5R247s9Goe6ZA8J4KFFzdwq4blriCHlPX0eNqXwJaOF7SeF++njAnDs0TkW
tSOb3VJRRI43LgFv/CHX80X62oIhRm2LIRAjPrPj7KevSjFw7diU9sSURAffWyrhgq3XZsUY6ovy
nAWzeDeWY3xrRDkxjxQAN8xOlyfUxlNsf7am6Prp3DCG9ANkw/MCyfCVBJXBbghP4T6GS/pNjySW
+j4cMtiThQqIcJCHVcAXQA0FAf6PbH456gYJfg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4624)
`protect data_block
9bSwyvHxwgT7yWWx5staR8rXlehJVMNxrlYPtLPs75y2InVio5Cf22tjKMblx3v/WwNr/ggvsL8m
DVBX2RnvTnwIIv+/1IN30j0dBs2yaLuoYXBhJyOTSVsNULEvO1j0/ubSacGQeZu7y1cD4I9Pq5Vp
jc2hrBc/EZ05apOy1n59AJF1UQ1ubvmqUE3C5xeBnZ5uj7S8t/XqGDLsawAhbQb8+ZuW6N6Is+4J
9T8/F+OnROpRYBYsCO77UFlL3HV2tuaj+2Lcpv+yjgTJFHpQQ7LNwwhgcfqdU/8kkMKCBNxmHPeR
5FX011MVmlbUmG6USI5X8LpdxYrWHeQhVipZ8bqpBX5e6hH1Kc3Ke069iggugVAouYIhtJmvAWvA
Z3KXhcTiMoAaxQdXE9RWstijo2Q1V548h/N1CMQYMJskd98HmqStA9/u++QbWHt7tuKHm4aVV2nf
k4Sp7ka5QSkVR2NwJ0MuiHHmySCPR2l3+Lzhxjk+TugpPc76I/e5DezCoKLDqFesA+e007gvM/32
eMIiSbUfEJs6xDzBkzSdEEDVCspL3o0+pjauAFrTHW0lNtTkUP9O14h4X+2FSf40xF3mEFxdtO7R
rQIHF6cG5wHb0eCXHKxGmXtjg5/AS26s0+hOpg1mXUTGzv0nP91omhJW7JwleAK8NFgyck7UJFm4
e9vwJtyzRn6i2RBVlYK6e9QdPgtFTcQDP0c1K5XSVQAT1wVRX8zAzHh0kY6IXw8na4PG2m3VJvSt
cv6TP4DV1k9Y3/RSG7fb2qOmNrlhjJcPvungvfb4n9ovn2/8bIUwtHo0+qaW2EAqpJ13nInGL9WV
6ikqutkvSids/TkVLFLCFURG3C9DORQ5JpOmRN1RKA3vjEJq/UfeW4vYmZ+EXcZDFKvUeqiIgZ4i
+o4anj9osogDXMAFPF45DEgud/MZj4yIirmFJNYfeCk4uTi7/88KYosMNNwpAwaVAp00J3do67Ki
Dd+L2qfMNVneUYs1IySdDvNqiEj7LVsp6UGzNOhT/hk7Y/ajS+/4UFQbEnihNaHp78sIB00uk4NZ
FPUy1xMZ1o4eRE7W1E+d7GFU7Ets84oCGFqbyns7MfdcwtgYLCQlBmU5adpTiXKf1OBSpkYZPt0b
ApbO1jJeqtB54jnH/d6xqrKw2u7UbKX1DxFYGkSkXkS5s+N5uIsRXoDC5VBaqG1hO8MGCKKQ+2/t
GU+Zmqn8lDor9GfFsTe5v9vg3LmjrcOX85ln4H5zvj3ECwAt8bAWNeiJkwcFYM7ulKgJVhqWSzgm
8zlPYCVKQSVoDy80nCEXrxVeExw0KFJdZ02g6wHOsYQSNUY9xFFvgqZxT3gZ2H1z14x9Mk6OJsVU
eAl299VefTvDmRiNYBSrW7DcfwlIwhqp59/fwIllRCUgeY1wA2/lVSzzh2b4uaCY8AZc5Sr7ozC+
Df3zTuRIbgkPosYkhA46sataad4YXej8/t9N1XNknNmkbd+yUfMRIj0LeIIW0eI8DCdh/hWvBNhJ
KoLV4voduAH4Gk3BRVWXWdmePkDo2Jx2JdXfc/RDLRG4W9cUgtn8EdQMa6PnGAFvxO94RH+XaIl9
omoZeUj5PDsCIlXY6GAseEqAYlfmljcOYZt4d8I8COco+mX/jmq5cyJCP5al107dVyeLMC73ag0Z
ZE8hJLEVPMA6B/Mi8O9xuMLq8U/NFERNK68XfVv3/QiSOy9hZXimZNax43tYfq+cgU/D3y+l+Pko
ChiiVj+TtaiUnr3EhoIZwFs7nD4OmhYcVs8+XyGJ5zETYa4pOBlI9WnEu0qfDNBax1jVEoHGgSyr
JmlxJbeFEmIzutX/rArv3yy22DFC9pzKikKUWgnur3oMif1yTJ6bspkoaLgZ/cf150JVbbq3sGaq
C8KEBJCecELwgJEJkpbGeJg7Dhs2yfu4keV1J497QY4tx037DjEmIjJ38iYjZLg3eCF5GjEZQBto
RyOj2YLj0IEzvK9cRxDAe7TBdBFdA/DLZgXScVR6iX/42Ms6dFRaeWIvtTSQHQ0gGp9wbbntuDeo
kVEGXg6w4wxieEh1HMthvTh8U0yJPyiDkjLSM9eZaJhDD3/QRlxbMvuhCFuWQnWERZXqbYaGVZOx
TAHzgjIT3r4djRJGhJegX+A8DJZkvrV25UoFKyHX7T68sgDF8Hjiam4KY1YRXsiCKZmTDGxJiihE
WCABim/gXhYKedeRFxZmVnhOD29FhhqldgIg/44hgksfPDUqEJhPG7P5hv0Y1X8zOlXl8kl+4Z4r
9ib9EpFqp094mswI/0v9eUlP/XqftNrenuL+qRZXMaxiJbgm+roXMT3AhWIlCmyec2Hx8CVdGF7l
77RDZmEpxtMGtWKQIs3vFJy6/U/KTRwVyCHY/SOu/9c0Pb6Mz6j4Aa3RCK8jFbGE+IN50jahdn1L
eRlpQDmfYRhZNAC6ElU3eKcei3G4vAnWoeMnSt8OF9wxO17B9KFi62Y/n3Im9+sQFWXwxRgkMPht
cR9OqsSppPffFhnwMTVoOqiVZ3MjswJN6P3jDbDQbAhrm9cBgypEwSfGL0acWdfklf3QXNKmDO4y
hmwMqRgv6++hqcQwnB/ozq86ebVVRNxWauMEV7inml2sKpeHh3tyQCKldjjgEGH7zWboIo0nGumc
0/gBPieH+uVifXJACdPzJp0DDyL+0wbUb+h5AFoPtky8wrW1nswGgcudir66aWNluiXdwk5ywJde
DER4nSV/a2cD0UcgWGyLjmibxWPtVPCDqWvF0NJS8US3qE8JN0iduV+Who6NpGUThn/BQ/4KYlF0
v8TlmYtIIAimUF1CVBcKAcnjAPenz9KKKVuWUpXMPrQa6Q6XuXd+Hn2STurps8+kC0e7ZKn7YW53
hCs/NAJPMXPaY1EJXun/6GW1sgVOJNduEdUkiYOs9PvNNKnG86od8qJzOavFdhfRWH7lVl4QwnIR
OCs5QVZWOiZx0dPf/zQeNDUyxvLJqtHKF59MBkdnnXN9O+yXKUrpGdv8rq/GtcTOa98qppFRGyJE
knTcD0rFyTWw996RhbhcYY3MTrxkisE42I9DLY1r15fpXTrE+5av6dEae1pdTpE/lql5clYXisT3
qMe0/zyBooBCRoV4IortFqHCjCjX4QDaUCNzYSt4Nkcs4z/TP+bqlYDbL+glllA3t1uIJSbtmNii
HBrzc7xb619R05SoNj8JfUP8ir8R1srpM+Nv1FmGsecmUFAHmI/ea5T8ECKjYGxhJ46ZCvofbGgh
Opx77/LXvDWyJ6wahcq2A42mHlC7MGVqevvYy9isknef3xa7SGkY9vxdj9EDO5S02ZC8js1L2GOY
3Hhr3ZdUe1zRhX0g3Mbnx0OVkuzHLqQflFSbOaAh8KDd6A5TL6yRXrVfj8mfmEeC6bToyRLVkmMF
OO5D1ic5Ro9PIjqAL+mA2pi8pqcyr/4GohFPeo0J5IbxypUHMEwWjCohVa6ukbgmbX9NXHj2bHgj
FjDlv+uU0AfTxw8lIMAJtBbknPfr1J3PL0WjzBrMp/bAKAJGkaEuxXmb52iK2h+AwR8LkRbjtlB1
sUR/QH/Jg+CXK9g5PX7YTW9TpbLO/bs66gHeiQR6kaKR6aOAdF0lvp76fqZcP2f8koBxVB70SyeB
tjMleC1GD6Tq8gFomV7IHFjyQv8JfUGtqWobPK/OSqq64TDSwktAUI2DTF7FAm4c95rrzN+mrBD5
4ZU/8IbNN5gUHa/++iy4OKvvm6ZOmqLDxKU2FDQ2dG8dbSXXFiEe+h4kwMoBp7Cv0u/OQYvTB5IJ
eNSLnwf6Qod++XgNhkUZjTRnOOCfnaYsKYRPy2jm4ooByHvkgavIEew2MqNWomC5qLmVMoS2EezJ
zRtPUDJ5ZKwCt4NA2qCVxbVGMecq6r5swjRmgprJPw5y7nsDdkWabjtkM8wrt3O8KJZKEuDsHU4G
2DRPFT5qmNuoRi0MSeaKnvIYLCtl7eJX3Nd8x53/djK+Qg6uKcVfu48dW/jZKR3ah4mtdhhkmI5u
cFYaNsvIHITxtq95D3KTU8nSwiSePcqXgWnHhx575KqfUFfbJykEOPju8zom3+7cFkF3w77ZgN3e
y4P9G2P5OlPzDCkORthFVFlha8u+btu/7SLvTzKfc1ZS1Tlbi4O1VQtL0B+O6RjVyOTpjVEMxZe2
gzmnO1M2ja6PFopymOGrexIeXffJKYfE4lJz+eK/tRllTN0GQg1jAeITlq9bDDrGFEoQ9hirEGda
g38KHYvDhHer01yx5e3ByvZdl1KGnp36XqZ+Mz3zer3opvUIG4oJXjiBDHojrHzXcUWELxhDx1Si
SEygCcqKhim1ycvEQcuCgMwHwXIAIBie5Z7+CaOPq0s9o1jlh9ujRqGRlrEPubBRU310z/8cUwZq
jPBybLuUhjOUfUvWGv/NuBl4nBlVSKKd5oibwZdc3WNcUnpj+h5mccWY8B+Ahp9gyDmiF3vSDslE
mGHgG4KTwTSgxTYkTKmT7vpyhwTbPAvo6ELLgzTrfl0GWnChGnhz4OckqbxVuE3AGU4W2jAQq6dN
POBDmx8/RjBqeqwMt3KWKpWsHTdmi8PqPrCh/xrlPVsOs2ni20RG5esqM9CDPHQHfbuAs1KE+Hh4
HqBW6w3XAKRmhT1SdkI/inwPTCS/TSYHJUfs2QBhvD7Z8rf8xhq+ZGKnxJh/oZUiguPfuRKHg+q7
aMESQcpCcsMnqQ/mkug9igTdUl4Jx2TjJUG+UkuTH614b1QjvCNnddg/NIRrrxCZ+6njE+nBKkQ8
Wr+7/v1LMSl5h4bD/p4L7IFCKvBDp+l0hmRaaFXtxC6FR4FB3PA4Ts2RgykcVFN4geeud8mAmj+Q
z1yIIj9qUEifpn2NiaICobMXzYTpOS+h9Jn9sGDWdqljcIa6YuYhnkS6HR3QkxNJEIhTGoPIt7EZ
mVZRHw0sxt0OPXN+NVN3P/Pew1UcBiMRnTRFcXvfm0ypx6Qe1MFcEP5FeAYwKZIZ0DIPIA+wFtzo
cWKOq06x9GpQKSe5xivZHTezVk8pJ4NivAEpOTmsv3HDVA6qQo2edPoQE8GwMWrq4INAzht4s2jY
r5/R+IF5yk//8J57TDBUmkK+oqhdEsY5BtR1G0BjM2qr/xeX2u/i0ZQfpbBZw5P9KQaLghD1ZLVU
CBQZX9aFkCVaTf0JsUJBca+Ux/hKvsjFSO/k04UCVoVylFBnZQ3XOguPnaiez5Bo4AU/LhkDHxRl
VcIlyxKjCDuAYzoYzz7n72Oam5Ug1yUfxfcVwoWlpqtbepkSs+HGiiMRrQttbMjJLF5ZEGhK1T0G
BI6tkjA/kVOslMlUgJXuBOhOb7KgOmcpykKEUmCmhB6KwZ+jSfUGGmqV7S9owebCdrIM/uBuZpou
nTlIOVaF67nLiuyeQORfb06VetQrLjBnpbVpVwdI0lz8EBm/TVJiQn4GeixssNny/etHBQdJ8n6P
mrxKTV0qxv7ZITDoVj7Up7rtiHrNEDNz7r0s4MqkMT7uk32yKq73AHYCmhpcZMhjSeZGOkKlWSZt
XbOv0GmLYRXBBKeBLsfLC66lTPspgvrV3kc/0/f2AFveSJJsO+sNZk1g1tj6luoWp7Jwmdk/rDgO
LPxYZCBE01rJd1udmF4Vcr7mnODOKvw6/kzN6ekUnu0oDEh53OwuXfUW+y9C75gGu/aEdRhqrq5T
qvW7GWIZevwaHmh9wCF8DhIFLjmygQKa4T+8ZrqCYUr14tqzSFgnQm1RUsdBdQhc+fluQZ72ybef
aMfkcxA5eeKYJ++U0YqPtbNH1dAh2W0UH+06VnPeGHewmd143XbY63ngdVueW1eZjG97vyZ6i4zT
etV00ZWJUDH3Hc18y1ovsfwYzyodNrnIAISQGO5mPcVkzoC5dJ/FIb2X0u2mhZf9nKS4FXqCJvSn
3ymERB/PfPDUEpEwmkbb6SztdgdW64nHAgORYNm/W1PWyhgdn+bm54Zc92xFu/onewoCSNC04/gI
z90ICjzN0ta2TbUoUTTIKY661CZkGu+3Hs0AVmo1tkW9TnP+dlC0JAgsrt4Hix2c+2+Xr0a3hhmH
4VpoNZiwgNkxlcSRjtrCXYWjDTANYYeX4AjuA0Hg2f5YxVco5izK/Hpirjv7WCY2516D63J5GowH
32hiODReHg==
`protect end_protected

