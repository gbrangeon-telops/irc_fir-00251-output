

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T6wVkTPpNtKFC5HWYRGz1pDJeqROUhDmQQB0XOtYU+hhB43DLNvsfjC5KYqU6Qt1lGAhH0laXWbY
sFGsB/1X/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Bo87Ik/z3ZMfvsxWdQ0fNuP7YOCyp4j/ygqxg4KH1VshQEFmP82QDe0umsG5l9IQ7WJ1x44Z7hUv
b2TxMUXo+JqxKnlgUE5S7j3ulzSH7GuiH1ZZMyENkBX9PvYGPAoxkfBZKwYBwge7dC+ekfgtgSTi
JmblFBaQfl2z3igDjdI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OS69EpuOCXkwKDIJ7c3PBFNFMJbX4CiEZKRiPCWgGoIatev0sXIZ8vRiD53mj0pSkbBqScW3T3bf
nStSylNR1BolV0YoJstQyT1+2pFYhZ1LLXaZugJ/oBE6vqGV5u6J3W5eW2CILy6xHulOJT7cesIj
cRuZgsZzN/xmRcR/wqC0vFpdgeypXB6mda8Kpubf32Dxwqfu3L7BPiBg+o1IuskbZi2Weoc3I0l0
OeBzQzAzru491AqXGKlZ7sf8bs7SXbbzXRpVODRt7n1NjaKD5f39RasUxEkDN/Mf2io8pxFG53sn
wj8Vha0LEKNulGqvG45lCg9sffq+6YoB/PA6pA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0V7+weIw8dZ+BPWec3DOIbteiwGwG6dN9psrs14jYpdIBALSrfKIpNuQOkhxmutTucD037ovCmPT
7tzlCJSh8b8Ydyh2TEeIpJfXn05PGHs6Bho7YXv+uAmzXPPeMsLwL0Zdj9PYL8wHeM9h3s3oFmE0
whlOV2wA/y6g8Y9g2X8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LrKyoRzDm4cxDmM9WZQaVOeA1DZCMC2sBI/JOp2hUeVDZFMUfjL+9ejUV+oaV3PC9kYwU9gS2N4x
T5QckNj/uBm/MDZii4ZX6FRa6E86JES6LqHqCKy4pn+VjDJ9xeobjj2ApHw2GympzRIfTHfg3BzS
Zkqs9Cmo3/2Uv3zdNyaGnk9f0Ojhxe+EEq2njDvi1AWk3nuKPvaX2PFiQqvWXWef/JYb4HJ0Tjlo
v5y52n4XeymzBXqfaj2Y0hccYVFZ6YVhMnGGV06K68vVbtdbUuaSPRKXNa9qJHwvtspPluLhH5Xd
ujRGgNTtTMlfDYr0Fh/3k9HYg9NPc+b+y85sOQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4096)
`protect data_block
jyZQ4jnZkoVYc0HBudGe63mkz0/tztd9OzHzts+gdlbY4/wQbjv3nKB0CX8fNQDXctsrM2tVm4R9
npfjgQTFibfdhrG/AU0ThinFFqzcy/6hcvLbEver2NA+paFzt/rWWnUOGOaBqfkJ/YAjZhSdUx02
enFupPHIgQmCcvVBh5MZKjVvKG+KuRNFLFTtCeQi7rV6q5qjxOh1ED/WAmtiwjJlwvVRZe9vdiVo
qp48i+nNtu5/dpmTcjaHnLTsOK+S466ietTM4KRizlTkLfafdVzDpSi09iWutEGzFvrJfh92L+JF
60O0wBGCI1NHWMBtvhAfbv565X0W6i+i2lijgpBJ0F/mjXwzhgyqwFPHBrKCsdcFXAz/2ubrX211
9tZYzcBJuf3nnZFbL20Caf5uaTkgld13iOCkIRXJ/jsj4+ZZDfRL4OIGCyBi41/hf0wOkRHH7SQV
BIEziRUyjQZ2W3Gl9IXOAz3RFFr42TYMXUjYgEm+9IZ+fWDL4r2AA0coOOYZNy4JZno6z/Ia6HGJ
MkWr09bbnUDaEtWPtbIcSVNzeDlu65CxiUNmg7y5Hql4hBe9ce0H+KCWz0uOfIMGyf+SAS4W7GW1
kL2NsU/lL23sadUUieu/sYBSESRt5a9OfibYNSGL6n+x7lJjqmmS1W47g8fctNuqTghq5cazUpzN
whzixMdfnuVQNLi0dhJFbuOcVjcbq+BnZOIvNjbdk1OGC2nU9buZuY+CltssQiNUKaTu+UNAI0xi
3Hj1ldKkaS9+10/KaI4VrtxY/oqU5tdJHPezRnfSGSTQMMP6qSTd5ok2jJoBLwx9CL10uyAE69Jw
elJcVef+ppL2NxufamGiLhFze5vOHBQgo/r8aKLI/CT49QgKIc9EXP3jfPmurTVFTvWiGj3GMcmc
OkEilUsy3JZ1BO0P1xiDvDi98XO9StAmKylAwnxe5GwEGt8EOOOpx8YAUedcOBVga9F2G25NhiSq
3+UmR6Nuk8V3Z3YlqOl07ZYnCN+WqEkWWCiMn8nvGGCs4oVx2rnOZ9AYw/+Ci7auAHirYpgqfkJO
/NhUD+0Fw8tTyXtn+s84+DbWB+aF8DQIKmSXfWxWM7JKxxj5zRrHpynxYlf9eEyRIJql4QpcvwrK
XRNmdQnVEBCGtgZAS5lIWPaHGZvIOcDMYxZlwUJLswwNi/hDsGNYigvxQt8EB1mOhDi8RZdGNJ8r
agN+yOCFiRzuCa1Mmy0TjxHvOBMTDV3ANfd/QCprv0LvjthFL9lOMoGDSi1GQH6I3f6/pzKQXBPs
vnVuqh5HiY8RajhhuyvXFWFVk7sdNd2POW3PrCwzVcRxwP6LZ8QhHIbJpTLX6vuErcZZsvP6sYyo
3sC9VJSUclosGb1Cmajq1pYhNL5AIx00Q6Cee0J+uf4EQweErFtkft0ClPPiloiEtxOE0tbRLN/T
BvFr3aqXUmXYulghups1+Hb1YLEvPvOSqxcfupDGYi0ZkcT5PEU4m6ieimyC0b2Ur1HwaPX+gr0D
0OgviSps0/Alpvq2p1PYzMZaZLio9dikTyo67SxEFFAXt+mwvigpANFdjFdcj4GppeJFOJsepj26
X4uFWY0zuJzrta7NhOVB7Mc697c6FScWc05HQDKeF57vHUsobqVyxO5wnTNdZNpfydbrLIGoE+st
pMD1hxApOPnnJyIS3vhyVeK0ivEE2gavWzkWnZUPhYMKJ9s+YLkd+eeyuoSQ+skDwQIZUP7+XOhN
4zef78Yv0kEWlpqgWMW8FFkcQkafI3TeFe3wDOKhPz6su+RC6uEU4L1hHywT89DgtF/HyVx4osC9
xpes5YkaBMACmMxui2upBPaXip5HBTNm1z3YREosHSyDVtAboiK4PsfQaS5ijCr/bhI+E5Sw/480
yJogccxhsa2qPl4M0aALjwCdfom0/jY8j4LCSsln9pZFIEi64JZouUIyu+GFjxMLSdNpc8h3Ej5H
xOjF96hxcQDjaDrGJFUeVdPmi4n7MRJx6TaatpNamHbLyhdk4oTOSnwz7oDvJyOQeOlsaUD+Wv4O
TCciA7sLrmR4c1XBySE1S2u9FIsQR70FDFZry++RtMY1zW/JphaWyRVGxYvygrs5OVuitRuGPFwP
PZ8idk0z4bi4T7bc73KxstN4dvbO0D0HndY+FqDFVq9Z5oQO/ckeG/UlNivMGHAB8EWtnscdmlhe
K08nyeC6VpLvGYGZ+5UXWhEd6j7YLMPQFB/mF/LYyx2sbFsqfD+1sOop3go0VZ+KBRPk4SEW+p0e
A84HpKdqAgyum/L2C8ijIV2Kx4qjkcdbrtTV6grnLNvigPxFGBxk/zvVv9zRwSxJqxysNm6u5zqQ
IehXkbmSoD8MBQr/fAKEwvN4LScT2suLqTdocJb/gPkjTrxRWRetR4JmJffPFyyl7FJNbOb76qwc
wiy0ZR/6f/dzxFFsUboFQF8nrMmeO939by14IL9gJcQkWU609VI4c1PobdysVQ5Te35WAiwCnmLb
nVT5K+sjI2avzLIuCNsaQ1H7q+6av/6CG9hF4rOo3cXcmHTf0H+TMXY25hnykzaybYgW3DWZ5qVZ
PrPcc3qH0SNYdVcClI9X0ZHBbeJhD96NiJFrMX3IL8m3tb8nuetFwgXZWdrloZzFayCV21Ap6Bfb
ptsTA55/d35nITt57AHFuWB3R/+SrK3F6oOVpGJS+hpOWSgZjQ5To7HxIACnnQf+5ww5NpgOs/nf
K/Rt82rLhtP2DYucBjqSqHijaNw9ugedV71gruEVbLq5aKnV/fOjAfmLWMpduUhAsgjqR+cuwzw4
MIJoG1LyjYcIFPJNdcJOCDytgdMpBuoRVG0DPo48Hf6rYtvyMy6vvMrEYhdYcO623ukxh9qqlVof
aFSsZK1IYOn1/8fNZM2BdeeZuyyUIjOyhbTjdWW12J8xAI7Hcn6gU7CFdAO8d3tnq2VO1udtL8oo
VrA2XmDwA4QGFxdKizm4ENrvt44g/fzpWR7vaMZUp00VcJQIvgNxVBeRfPNMtPlTK5A/YSn4dXI7
jNzgPAG9TBZOaBQNjpZMt3Kf1RL8F7NRicxSOK5TmzH0v/KE7T1AQ1+R+WsXSiOr9XZ+AcQJ7cmx
oplR3CEx2h9Yx0+Jr4MFdo1sbxZBLVUsHlBG8il8QoggnusEH11ywMiC4qzl5J37crpVXVl4/Nyj
qM2t4KW8KtzFKcrWgBtlIi/OI/x2fehJWq6Wm2bqYNgWid00UTscRlZfbNkgAUxGZZoRxZY460uN
wChICXZ4qtW/+HY+CFbxvEWkhZesR3cSogm9BJKe8snofqqSavkh0XHHuLfzCBesEVBuQDhwYDHc
VFH8qN8EV1zlOGfZzkcW3CbzHm4v5xN+NkS3YxVHQUfCzN2mk/QZDGTGwRziMmwgAkBCjQyxvLgA
EQLvKmybnKuLU82qqEGD7It7Ui1K3dkdtnjLxqvSdy2QP2fZQQ02v17Sk8H0to1HBgNp1Edg+plR
Y6Ph+NS3km128y7ybdY3HLlLSeTwUG8mwArPQfC9n48c4BnrSkBOHj6yuAySxQDZhCq88oCW9RWa
ZJdHoRECsztlDnU8MALPSNgE1z53HriUVPTBtugYmg/OfRHjvN4ydQ6GLBNYKWB5BdK83iix9l+K
Fs/EbYPLNbKR2bKhzq5vLp3uSwxQ/NQwPp10wQsyUa7T42f2vSypdcUHKfudAVBkEOJ38JYFyXuc
52wSQEoM+QaqrJnQm1jvtw+TgGxYPQtMLg7PJmkgzicM7/hs1ol4kX5HerOtQX32FZNEUbBz7fAh
4mWGhIgc3Y9eqa29Sfbfl7jyK8R3CyNWx9M2glLRs9gOy2JykipUoHjHmXzMVKccs4ytAtZoAAEY
l5Xh98KOFcXpJtBOf46VP+bHmuz1QQJlr0LteVJxKlazgG2409Sf88eL9v9PmjBc2w7vphCTH3gL
sGANOualF2Z4oDakCKJXMQ/LY5EbDSIgVKoMkScB8ArkhSw3XtZvOjK7G2bT5OEUNtmjqGMptceK
s/sviWydiyvyOxycGFmB4bBW3yy9qUKuHBpoNrQgDc8Xfc4vAq164pg2F7r6cg2m+zD8t3vBoe6M
fGzWUtMRm7m10sHi1WrvLGlhHdcJUuhdZmofT7vMYKOVf+wZXUr4gHCo0Dw8m+9nw+g1nS88sTP4
FWgk48xqfKmoVuTvS3luf+nisTBeCjo1wrKXaxPAcf7YMOOvUVC4RhH7w4hgg+JiUr+L/SwaHitZ
RGXrQLYySPDlaXEgMNlZrkbspnpfbLxkd/A+Kcofcy5g5q2nYFt7E6RUeb3San2r/BNXeHl9JeZ4
Hhsi8PNPia57uuPbMhMGi3sWp49rO6ULQBbewk60X8+1fR+PEyY/M+cbEzR/lVX8Rh4eNrHolEgp
87WYB0E74BrPTgy/bCSWA4Y8t6bTJVArbWdoRtjDfE4x769kQV1DK2SqA4gxescMM75BEd56XLit
mHdaiGFBLHgi0YJs1qc/FcGVuayN4wCWbt+eu9vIoS7NmM4fo9KbwK7NTxibhE0yl/u8AcEJhbJw
tyLOkcKKR9tsagCg/FElKET/g06FujOzIsV6GGiQKON7xBbM2kBRq+Mhq2A9FCoZmhehK4oHqApO
yQ2eT8e8Z4wxLIspjWq+J7G8MK1wWcZHzHrHm3xbOkYj9HoYdIGrReeF3Z6jMzTNMybnTnIQpP5W
HsEdiM2m0wEPKzRm/zLBfuAsUkgQzKAHWbe1KY2P/iLEyz1kk9FOYo/FHYrpybUUFQRvw9wDt4vu
nAllkK7d+0rR0gsq3VMF6yTmALurkKASmRPfTNHekfSUMk+hcCBRu1NwAecONda5YIbKZXmu0Nt6
Yx4KZsOLovdbtvdM0CVsWXSAfWphi2PcwcIDHGQwZFrTs6wCru4VfHpvmUNbqN4qKQWevgUmJAeZ
OZD6o9CXdtaDzt4vnYkeqvQkJsOl+SMADfSeZ4ROBgn7nbOMwpwf1Qi9UT+C2zTJpFJER1KAVBGj
2iMJEFEM0uGONAGlQzRa6woHC9HpGG2JAsDrsV8WufhQ90G6KrqAQvX1f3bbgQPN5dA0kzvYVKXq
Rpu64SPfa0qQWtN2fEkXb87m/z3z2uai0nId291RFtCdLi2Aozs1d1wTQpR0ZZGRWUj2S5xYc1o1
U1M2Nnf9Twyf8GvbDLY4l1hBw8hNYSL/r9NyNnk5E72Z33i02Fm6liwubisJ9C3VkQNGAo42CT4S
iUwXYPeITYPUs26pGoDvj4wVxWI3S15D8HMhYj23XkL+l5nCcXR1lednGCMcYuhGL3JLMS1CWDB9
eWUvXR91hRsOswY4cqF5bs5P8aC2ylF8av5lDzOtbgMCI/izLQjdrpjRooRFllP+0jqiXdrlO5OC
zcKhTJ79juhNsXATFrPSo6KQEBkFyTjUvDpTedYS9cHEFQm00As73asWjjKVBWgkRg==
`protect end_protected

