

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iEtOB5S3Q/0nxxj3yhZWc1e9CYVNx9kxE38Uvw9Q5GTpbeWA/PaP7MHi1hZ25jWcWTCQq2m6lqXe
j4/ejpW9UA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Xuau91ineWkILAnXNctj7ghjv8v9lVNvmGeO8/qKPRA098IIoEEWbPkQsDw9y8PN0Kc6j93b9RA3
24AkaGw7vS3twv084InDNHpEnlN63djkx5ZcyOiUohe4xecSmu6QA9TFBRDs0Woq2jQD5/qd0oJL
/BaRHEN9wihMkCnRmi4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DukDx60lt5tRoBa9fYOjxQXcMx39PTzSzi3mfBKPNtGRH42SBSoh47iSUDQLozXc9RVtQC3PW07a
TdEl+U9LI0QpSHNQLVojqhahZCfYOg99dtV1mWPojzxtpV99k2zYX2J3PXN/YbIzV8ZxTpLcq1Jp
CAIcrPJ/34KYVzvzXFRsvxEfk+CxS8lIGg/nVz9ZI/SFfi31TG5Gc9nsiydQV6NxDLfMTIZ9geQt
WjMt/ZdcVbixfIDM01Blr6PmvrTG06LX8uxL31TQuw5SZfsZBAh/PoXSzsMleljAYXIhMhdSUOnh
qfkHi0I/YHOxbZGvwoECi6yzPk1O8e4p+mbfJg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfFouWl9C67kV59ngW+xbX0i0eu6h0roaptqFtm5oV4WYkqMJEDqBwmHay9e7sJ9CO+K40RDFIJe
/eeImbz2XS0Q6PwgmMgPAHRoOg4fHkGIAEugmb7hj+mXvk7iQo09CaB7HocKsvGcx4nu5U5a1pLQ
6UjYczksNjCCieDaJQc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RNy6OyrkxjF2nMK7NTVKf+mkYRQZVhnkvdhxFI69h+pJImlNAm3GMG9cNkr/rYPBFr0KpngtSqYa
zub6qdQpsLCoZ7qDFdEc1+wws1xQHHeB7VAyyByyPc8Chu9XZcfd6cEAYC55a9lNvtmKoAjppEfF
hj3OtTTwZQDicoWmteMIzi2n5YcjhwpDSzFHpmKq+NQje013CABovpP0/TVMHv74ZpkyX30HW4tb
0iH2SzLvUD7U/AR0ul2kht6wcMaLE9E6bQipSYn1DEnfUpMfQgGpPJCWjykHayljMFWfI9ucuNXK
1XTo7EI77uCstdWwv1uP3ZSQ8pFNDP7NXG8mpg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9552)
`protect data_block
FDHYNkP2dKjA3jtzFKUinQswmTot1XvNyyqe76gkXa5B+J6fihD/ily2NiYVCbLL+zazUGmIs/kT
poFvuI5iKjjAibWevpQTVqaIUufrV4A4MZavHm6If3+zfcVuNPdFKgVna83dcXVCPQ64euke6gwG
KvnLZkzwmNRuWNWCozk/hb3aQcvJ6fq6Yz2FfGV5DEj4fTZE0w47Q+/JFNDB1qe/WX08zA1AQKEl
DhaNmy8GG6yVn2in/c1WbmxHAKpR5H91P8vTbkvCVv8fOmCSnXNrIj4Ess4lsHlwwn9e3r1iIBQ+
SuD15Z0RAkxBPAtWwJYxRbuQUT6XJwxH/RFhDn2boyb75uE3aBnqTMzZAacbAsodcoFYrQTNUoQT
mYatXv4sDDqzFEhf9qaXb7D5mUps0Ds7btfylxm6EBZ2qhBmfJiHna9k1uK9FO7ePvBqylhqCNu4
6Y+8vlaZJ3UA8ML05lfGAFqPrk9731aToZ6VMIpuVOsyjfkrEvFvAjRLJwzCY5QnKxixMx7y+oYO
ekW5zFAM3yGL4aGyJ1IFabJasczpcHu5R2sZkuZLIL3oTy0WpJF6C2MEUF3Y39jbeVqV9QS3tPRa
6czOJvzjzMFmM1SQys+tWW4uJlaL1iQPj7svkwFI5AqmLNB6avRn+wTq397PUc/FUWZtYrOgJVSf
7qcR7tG7qDzRi/LmQU+wUEz4LHVw64GYZlZZKJXhTGA0yhfK0ubiFSAaL1l3zKlRibXRbaw8BFlh
sjYurnxDJpcfRTcNof47RlzR0/tlozfCeP/ZcHimk1TGhcbt3jHxeQAXxMe/l21iodnLiKdV4Oo1
9UePJBbtxc1SaNyxC6tKMzZCehSLkkqLEaMxxR/EC4WAhgStUryYoFajdfULR0KG+kdd1kb7r++6
eDp0OLPBQ+Xs10v4uDxOvSgxv4A5tBlQx+jcyaCw5E0xbA73DW2ruY4tEX3EswTEUYhCspk0fLrM
xjhoQSmRt6lSwnKJis+4M4XG1GFWqrNcygf4Qbn2uh6i6d4StvE494qaf0hyJ2h90IOsYeZ1akxK
qhDf45o92e1C2qnn8RA/xGh2mUbGpz1mbUVzYwdZFpM+kntOXxOiVBeGsHYZr21rvs1LyinFrx+y
tEc/OTu53HdupQR5//ip856STNNt4yWTuQri5mXAasHPTCSViJgy3EJnJef7FeZvKFyAad2O/MVu
t/a4y2CxaMokr/NxYNmY5MfR63f+R244QJtL8+Ts3Rj0ZXwWVIaR05WEC37R5N8DNz+n9NeFdEUZ
b1NElD4a67QM2H+xM0jLqiTBlF2gKbXfC1fT2+3eIL+I4jM1ELkI4CW8NJRJXSocMI4pMyhWjBIq
jN4TmvltQP5TeobhBhaw0X7RNdewmrfZdjjjQV2PxSk9SPj0H2XCZm6ptd/n0JC3ZKd8/nwvThko
CvMQcl9gJxqN2B1Yh0aPHfDv7IzZ7T4vkr5UNyz6FOlQ2tFnB6ShapGLoo6+wOs/xJn/71cZQAFJ
ICtRS8L0Qb7J+dX7FnUtmA/wzyG45w2x1fV69M9ngbD6b8MFDxBVx1xXv18LgvtzD91x4nleXsv0
kPD9sk+O/RTqFusMzBM/E1J5X6IN7W0nESKvCLY50pOmyfkcaclzAHF+HfQiWPRLirdMXUVLbIi9
qxSxtzYerfNsnVNEdzH9uYfyZubt+HvuI6JFKoqSe4/Fx6w93ZreZzQshpWppTbXaPNKuoJYMTU5
a9pVFSN2Iwmbcn/vCANUPEfLH3/erULS3Zu7rDSDv5PVV5zNAKwZ7RHY5vaM9HhhEZtTsLiueMqd
tpb/t6F5yB86tYbbrbiyrxqRY2eoRJfyhNQ9GknF6DlD30IOW4nbR/osQvHnY67ybJ+Oi8l6z6Fx
AfIOGHbfBSoUwM7sa2jolXANoBimtM0d0AiNpBlDf2x9qfbXcptKvkhtHYtgYM4FM8XEV27LuQe+
C3/SoVvEs6TeWAbIc180nmtwL5qUAXGnCv+8dvMfupHnXwq8s/5XtAQ5sy7UrUEJ8ztSX9LXJAWF
9UF8WlyLYhfIsN2r0aQM0ZC2V+brDeNTmbGcvPXj8Xv5Ndt1NSiubShFMXOeoHu+Cd2MR8CAQGUo
PSQhh3/NXhc+Z+E20z0MlF6G2yfke28KcaE+xM5J0BJ/zNkxNmVGwqjMeBVou6uJjlmK40hXAuBA
CEegIC+sypcayIe+wVASMKNtxy3G2CH70F1KMUgTO+qf7bSqbd2rY/wcEfUgV7G5kI9aQrSInQ+R
75z6pnZoSyXvhbBkDJQXXIBX0ZmbHtzPybUpGDSE3bSEp6/ognawP9NdnzSXBy/dp30NecvuFyO+
RgR1xYE50lXVWM3xRrPEg9OSGgUpAbDh178sC8pT0IFuSLfg8fwAZNBN0EBWvHWk3KEoVprVFHCC
NE8T7GdxQI/DNnOMLvsy2eKDB3DOXtRjD57lNmfJyvUGV1DzXQzflznAnTLp3MAZOMrdUd3IFh9/
l2VTBNxK4/FJeBch5F8U+y0dhh8T3RxFiv4+DMsDnx9S998e89cNkDeEUlm+yF9l1N9/5+oDyh8d
ZIw/7HV0VGH0f8gfiqCxP2rHNEEIK/qGdZs81yfRDU8DPhf6TWTPzhbdCG3abkCGh0awwfhI34FR
SKxPSreC/ci0Dl8qRbokpvg/1LyP2LIBw9BoXNj4TwHljLgaUP7+7p0VNvA9IVFStCZkomlZdttI
r0VbBeh2Hp4KVzFmtwtP2KDXRWCZvfdFjw8beur5J3Id2ufSA9cQ8ZFpvN1xQRTd1YvYw9ph7aA3
ucC/PaMpnCETOP6Vx5l+acedDjdeFex0pOtTQ7MX9880hJ6jVfeHTZlIzsMNU/CQSbTs8qLCzB0o
cLnKiXhx97VwvscrAJb+qsb7AVLaxHYwIfZ6Lc/CBrZHzbpw6TArFYjQpTfbfLjwTvzO1r9rojbz
DBrP7ui9yZ67APu1MTmMWDio+1T924eWVjDLra7rTAltY43rm81EmjK1R5yt6WdA+SezmYMjHC6F
t48GsC6fW+q692bsaevIp+OCCA+N3uScvTe53bNM1aJkrl2Z5oRJrMBFbbWTHHdRwTTO66nzmmZl
k0xM4uXnBJ7Y0kYVvymjhuZjTiCPRLC4qDWl0tzpLvaf5GEndaSrMFHUjlc/iCefDbCGVsPRy8fU
1eTwVmXtnD1eXfvTKkIQNyuCUyj8Y6SNwJvW12jtk6WHlgxXtb+kdu8gqFLu89v0dMoWcx0QcHvy
F11NCw1SxAGP2PbJEskBTSXBM3nzyGJMTPEexRgFz8M7HezIjTFLgrZcq/e3qtR+/hYeZnNtF0ZY
QiOBfTKjVrKhXYCpC3/vM87qtAkU1qe8f+vf5Uwq11FHhaiUJ3teOycKkNbdUdbBf0VqbKGNdD56
mb9NEyGMek3ANJ2Ys2dGbKXOB/0zYZZQOqLItX5PUhwyHgtTlyz7PARNiIr2n+xCM9n7POvXRciL
UzQLyT4kQ2wutxTtvTBcAO7F2ra+loHV0xt3QDhRDrANT0XRxf3++UQAWeIZkZeMBDAtrfxbJLbP
/v+E9yjA55yfajV2iB8XCNsn6d/GfA3GwgE56s7n97h1EIii2evFqylyrQEJSGs3ozhAP/3w4mUu
itC0ijyiN6pOUzrK4MYsed3H6eutbwBHKNguuqAgngWEIn5UF4QSR0zokQAD1RfZh0IFy3CJgsBU
Qo6vk4xvkIWFt+Mu8OxXQRZngYF3EdKOSS1N3bI/k1Ntn53mv+V52qoO59Sv2GWC/nlVS60Yxqwn
mOAmHaXZMf+3awvHflSY+deVR3NXe0B/dams4XcHwpoVabNVjMxJ0cpkoixH2E2KbfOslEc/vX4b
wrBVxjTCNBXjdq03JuVzZtG3xidbATEo/rcJRgHXjLQSGA3EVWmWQIsElGC2Z7a9+kcbxaon4SUN
MKcHc66FqX6a6DHWy959dyfdZ65We5JdFUVrXuow3Fj1kfwVdDC+EXZ4Tqlw01bTtMIYmDxLJTLs
QgR77YzbZkr9JAftUhX5YGdbgcwODXrNzS0AdoQlIPBJqW+udLg7SoPUfOmudzKjIN56XtDAxJT0
U7c3wBc+qEc2yRhxlJr1ahInVF9UvJfv8tOED1SB7B8FVvv3CsVcRuFuwSwSCD/N/eJQ4Qw0U6f3
s6iV/uwY1+GLkqhC191AOIKY55YYCOt2gAXb4RUHb3jMWSjnzv5T4ruIvcjlzlTKbmeBmHLkEhTf
6P8I9xSElqCYFK719WJtio7udR8MNWWnk6JFnQDqMqgEMFX57DyJGY8ccU/Hlbrg5IQEbOj9pTmM
vqvoFHXFd1Ng69c1N4Haq9KLPCIPa2Ti0ucNNf2aS7Hl1RNh3cpq6L/p3nVLfeMcUJDZRbzDouef
bzXZ/02GNWCZzwxiBjXUnfeVQ6uktjkyiue9CNVy641zn+iYhNK9qv9+RCNDXuTeNzyM3MfxayIe
rcw5+mTs/xm9Uv1AU4rmM/+jnWGTfHDQOf1n9EVziWKJPQ4WaqOrvJ1WcLRz4PYEuKWhWRnNKae3
T6MF7rbLzLWl2V4eeD2VQa4X4sEegP5VVQvAhOeQOnjC74rUEiRPbq1cVe2MVfmFjM4H05jAcOZg
I6qxI7uj/gMnm2KrfUAnZPwTdBY1+fxik3sGmeL0TOzR6wRoVrScVBuCByZkdgCaNNYXHpJR3NCZ
W+rP1m2NJ7fLj+enNhrvkNtTulTLa73tmMFWMOQYMk3fCT3RRo5Lk8/yNPV0ktkuZohZofdw6fpw
2q5Uge60Ew7yK3iw08aLiVC5LAUsIfJmaPM4OmNDv1+Y2dxF7mij+QbMOfRo1SHL8q2oDQ5YYVKe
EpDVnpnWzdztraQHCYvOBdqCOdsB04sFaEJ2Y4Y2Fiw5k0P3GEI+/7BgWPh5P89lGp5ScRR8ArmX
oHdNZkaCGxaBMX+PFdeBuHlZedXkX5+HdHqjZmDWQisa+X2jz5uXebM3w5p05p5wtANWU58Lhrdt
edXy6Jg5bHKcTEB0bZuV6T57DPhh7GF2S+0j7SryX3edi3H15F1pyi31IUZ149pyc0QMwVFp2z9Y
/bdr7e4CxHPn4NBjR0pE9oytbQ/y35KHzFlq8XUJ/YxDQR0Lc2QCylaj/QZHqoFG6YMg0+umb7OZ
imSd2mix/kohkMxyB8O/8SVjrnIky55IiC7/jPx047jIdyuzdnJXQoSBi5WRLyetuBtzBH8hHbX0
/BPJOelp9IuZxwXAKC/8KSinZxHMEoXl8zqBX6hIdmEZnEBOrdZBQxaQn2NtpeUAqnGOHZV1vT0S
ybQQd1AniWUFfFzAu53/9XP3GOtjrSV2fxslbFh5fbvyQOX6wVg/4WdXHu6zgPkYXYLalFt/W4Wc
P3g/niCRvUQ+AvEcemDvrdCPq6fiVKwlyXg2Lu2T/UZev9+wgscRtzx7pu9yhXnWOyQsWSXWeXei
MHAkDOnPLNiPP9iFPTrZRvcIOtI8BSL9vZTGnFeYTw83DPl2DBOnSX9+ON7VoCNunFPUynUxkooq
VgYd86i/Qrvwpv8w6dXsLU9r+Qmu+khVDltUriG5Z5bmQienJ+KL4iDmgUwmleUU6FVEPqcj/i0f
NKBrLO5x+oGJFe4WZD5VpZoMBgfmo39lso1jfKNo23oF5+gUx6uWTGh0KIRF4tjD5GPf/MVjGLgb
ljKWRn/KnGjqLI0DywWswCen0tdXSORHSqq9F3LUjT97AeNgIO2/Z/ttthiNj3FUQ/CKi5yr9i9u
WkRH44LL2iK5QWRxW1BkPOoT/WdPVY5nuFwxfw2uqZiK7FSzxYliOD8Eo+EL4OsRf++TV3C7TJFP
SvVzoLJse/4OzfMzxxhN1uppat0XEdHCtMtg0oCRZ2+UGeecn1jDQ6t/+svINnQ8xL1gHEFyLG2P
SldWLCgDS3aGDKYpAsVftwlW+Z/8hK/M7Mf4bwPIvhgq2+sl0QT2STytL44q1fyM8c0n4lG/PWlL
dmygH9oZt5GqafNvUMHcrgrDvYTd63u8kmylHVXI7JsSou+ZbObnPrxA/0dHqu2ZIoIJw5OUXRO+
n7lmTX19G57MtEKQGRN04UNAC8jkNhJoR3XaPCrUXzBrbsUVgmtMwt7VJAefR1vE+s9ai03wNwW6
OLOdLbbl7X9D931pB9+QyEo8FSPdJBCMnEgV9zvBfikNZEe8QL2rTpj0A7YmcNSyDWrvfbcmpD3X
M/Piq4f853xfb/260AXeRyaaAVKvfzYxUEfSQ9GcVgzEhB3GdsXHdCtsvlSEZr8WZT0pAezjdNNr
/JRr7xZDa+le/NFSHY+9KV1pJaChzDKiynwUuGc5VyQ3KzK00Lsso4we7ZUsSzKbSGqOCEdIrl5/
DipfA8vH3+pp08X94t4ppsrNj4hUsu/I+gO8uV8qVWblSu8U/5ORN8/JxUD4VlxSR1mPisa24rsP
jXVfD5WP+E0261FfhiwGjAFF4lDuUZ6dz8ZR+ez/sfe5rnVKgL/t4cG18xWH0FoY3dkCFMChdb2g
MMr7sPC/ANHLUmaQD2Nt76exa6B5awkyakF4mzNpOAobVvd7/u1Zt5WvAidd+ikqgzLz2ON9elAl
KftB2YYbufX83HauF/BXXnacEUFtRioblrU10wNYsL+SOwwEiQrcFnvyHqBDhv5jlsoaBcDjkw2e
dojcJvLLySiQ23PDBQjlDD25e8ia/TnY+F46y/6Pc7I1slt7jKy9kxf2hcjK6c8yPTDVPayRoxrW
WGqHqzQp+Cg/jtSHe1+Ale7ObfosG2Liu3A2Zx2qhVTBnEUaXMaMRljw4e8k8oq4UXQG3i4Q0vCQ
e9MX4OyIRndHUiCpSXVVIx4taUyTpiV0oczdtnEEZFRfCq20FQ4H94SfFosvgFeoRY4SVI5FrQA6
cNV4jkHQUsdQLLHQ55oPRHCJwDvfSPMzRz1yRS90eCQh5pv6AtoOBJNJ/hIODAoPRUQBUVroHbQ0
FqIpZhQDKtnEvirM67vvyJrEVxDx/NRT3ll5YnfZvCX89KLgnsR6v5LPLYgQqFnYryHWoVSBZ0Cv
9pvcefa3nCgz9oJPqUd16ynbwisNu279ISsx4S0DHlIl8Gi8CKS5nwL1gLsdeFwmFleeK68XiYLn
5YgUMVkCORKWYqw5gbRM3c3J3aQV4jQS+I3nBccya57kYWuRDly6BaABdUsd0XEJNGE7D9+QtHW1
7Su4qmzkH3kQlM5nim2IrsV8CrlL73fVZ3S27fZV7BB3bco26FFuKtB0mxWWX0x8TRu+wBih63Xh
cO1gkfGm/fMEYdSdyy5xtK3FfE7TSm7fE2IKsEcwKsdspqIX0iBgXme2Z/yx7w6wqwaZrjQT1wTr
rPwV7Bl0B30JtJNl9cGbrpoLY/LTztH/TckEdCqMJArn5FlZFRuqbjt9Yk9yYNGjOhYcrkNGPH69
e5Gu315XdWFimsJWTrF78HDwwSYa/0DWru1bbPFRG9o//BLoZjCAs4ci7WFoQlQ+7HIuGoOR/6TS
U6eDpHkKBOqdkIExc9Po6jCsq6vfzAVZoxd31L8PgrXoqhjWCdnKlK8g03CgX7HEq64J5XZGQD1q
ltPcPid9421Yv1Mlj/7klCanhniMUrjRED/JMwnlVMC8RoxT3kIzuwncplGyj3YiEyHb096xiXro
GvgzBJSYAGZ4rBBuDhhnVIF00HRkH235t+fEcfeppLWtV7GwQcwM0D8OSSBRP2zwX10njQFHGOLk
baqX6JHGfGwaShHJxHSQwcMTNtbAYqor+DJbNCDakV6IjIS52HXtqzM9t3PqOvOFel6dDASz23Ff
gIlOP+kiQq/yvRPEGazlVkQqsZltUWDNlbWaDXJL8T/NyGyr0RKTOB14gmVf7XTTyLc9nFJrJVuK
fHFYidKr28hmol4m8hzrPzpzkGeTX3b3Kyj2QgDZq6KK9wUkiRZqGCtPGbmVaZ4BjQg5gSHSZD7U
sSFD7V9RfO72Pe71sk/IZwqgLz97Jp+3IsYMfDFPHJogY0Ri+A7CKe7o7w4jmhzKybiVISnYQLA4
Fx0gCLCxIZ9IMlRbVkI/6SklDc1GQU6xCCoxgRiCEfvZRRYzg3XCbR6CInKP2aBCatcYGrdYk6Lm
OFOr13FITSVJNerb6ibPNEs0Td5w1fhlt5SbLGc84tnfQHvwRq1sZ84LhH+YTB+um98DCZFWedfI
Jnej5iMBh7RtXZ3ClUe/NlCeyO53M69YCIKOm49f6NEGY3O2V+4VICs4BIjNr20rJNN11z+ShNl1
8MdLv4aWRq1iGcWb/ToQqVUafc+X9n3qLfIC4oDCbTUqkosYOd5lEZb+2+wO13C3mbwmjLNQbd11
CPmRq9V6gr9BNOBfeDyfpFNmmrawq0a7zy2NAM+aJ2ankaYIRmatoxSvlgZXOsyvLEuVHc2p6UCF
8Dv2VmKyALOq/vbwclDMApEhECfl7gEDFanfIP/2iQEMCqxOdWrrIAEKVQ4Q2MyvsC1C3rx5O+Cd
Q3G5CZulN+RrMcDj7ZxSqbvZStD2GVgp5lMMtnGzOmVgrUpPzyo/lZjSScc4cWnCXrnV6Au6Se9Q
Jz4RTO5/PAlbRprLHxzopRN5JE/E2Yz8GVs3sSTjO60PzsqgSIxQMLsFAkOdavSr7J/IRQL8+mEA
KXTGl/FYI//B3rsswcOF4jZnXkqCCcU/juOko/UnJdqrCbfkCsTJTGpS0Yi1RHO0xNc22/fNzVSM
JGv68ozDaE7BOWfrUVhYW1PeRSxd8as1ndY9BYzSG5kuT/QKTvbuajMR11kWdYC6hruxpf9xMkfM
Vs58lLLdgLoycVy5RkvYga81VxN44ymd8ZlvrP0t8J8kp+5l3qbQj7qNpcZvfG1KGZIjFdFz9aPX
ngqT1FVWvPfMxLiBGjfsWctCn8OHoG6uXyLYF7WtNBPBti9OUJOAo2SdqFeZXZvI4VCPF2tUSVXR
deis7bI0pGeierGD7civXPIvXDK8TH5QREdvi5A2ndIsBcNtdKeY9hEhs7nAsoiEoYss1Vi+VFHk
K/+tMK99pmya54YyrhR38XsJeSG117GrASME0HoIgUdUNpcARN4SHTlcW4uJteff+QS79WCwCGcS
nT7MZTO2v8DpQuDBlEFLEUi8cmG21Ua14cctnxyD967k0C2UWzyhUTikWAa0csYHUxxgLixT7IrG
jsm6hK25vkK2u3gDaDM8YFr4z2CHvJNbOQVcuFm5RL6Lp0UQM+piKxNNK2UdbHX4FR5PK/Hb2j/m
A0NvnQVprdGo6xMhKkpQmzu+POXPpZRAWOxinIHk9Bt5wsolDQTDBs8XiUBvZzeY0aURaRhzIRmu
FaSHaHnQoHHNJgd77Aav4oSyZdghkQuDamDd/7fHmm441p1BO9Lvsn0RuYfjNNbF5CTcj6WjnBah
Rf4OyT7CiGYVpC9esCn0x0Ob09tvahpbXVGauea7PqOT6VvApdvpwAYRw7xqzarpcuHr2eN0/6AN
Mj6zvFia09A9j8pwIpCoCysQ6tMB3ZzWU/8bqMSeLLJDWyvdsm2cGWx0PFVm4XlHNaOcbKV1OrHx
aiQCPEm5C/aH9ukTSUOE7+LqO5YjatALIFjonxsgiPeVMAUhMW0bzWmBd4fJGv2Y+39X9nGMAJNf
rNH8kuptUTG9XMKGVpHRr9mD4p9WHM3RIhU+wwW+V8qwQzMLPToc37XDa//zxhqElKEgq+YiIxiF
+e6fS0LxnVqkYhwDo+7BTilZITecpCP4DOfoe8Lel00o/5LD+fYzukQsjVDRJT3CZxQ1ZwW2Nkj0
4hsYCICZrm2PToH5+pZZGuuFnbKgEfrjUF6fjN34aKU1+cJB81xGmsPRAzXxtee28hpdPZhiTOtR
Ax6XKIZjzU3FNaoNRMacXuhLV4vflE+1PesL4IfrF19HXJVYe24cT04c7QfDvA8XXiPX3AIe+Bbx
Oo2RAgGkhDOdZ35zz8t5OKYmARyVnU57ZEdTy4htdRBWtrjI7Ria5ABspDz87DJmzmL7okuGMxiJ
XKRmObbOKRrbmdiRMCIx2+MRQoTy3B8Gps+NYa+6lyOV6tHkS4axaCdPsUqzfdowoZmXqAvafasF
llJcN4iS1CDqBCe/FbwwmXFyVnQYTWV1Q64vBWrOPQzUGjl2R/qJASrcmiDhYZ1865vNOnDtmUdd
kyoyCuEvShXaZYcsXZtoF3HfSounGlwis9VcpCX90k1+o/zTRr+ReL5mL6NPs4Y9YZ2yuNH0pTl2
YHeW7N4IeOoQtWsP8l9GgypRCitT9Jq/FPUqItCmal8W5NtB8yBogRe3sHe2L1wZhnmjC6sXfgOZ
aT3Q4wVq60/ado4yVwYxpACgDNumvUIxrgtDJzRQX/tqJXm1kd7iZeJssHncBACrD+ZxIYRPzoOD
6mxZuzQumnJAuNct99tylfvS+8X/s2LPvRJDdIQiQBmPSGkZfwJvPiP9knKtTrEsjm5U0OI2tb8C
Pn+VP5Htk7tKntmhPUCZgU1bZ9iVAv6MYEUcjCcTfBDQ9Vbk7oVo4WEEzdx/m8NK30uIXAWPS8LF
dySOXUnI0LrRZ+1p1qVulARlv6gQnDDUeU6+Qy7M9HnX4ue7WCM12Avk6MmE6kPqOmukD1xFMVYz
r1PBvIhZhOqgyM+SxHrgha0SjsOWMgB05/IDPPm3TvE38jyRGp1XRIKJ6CPkO9UBfgCZ41DKFrpj
5XRswRGAZd6T7z+GdYqYr1/JQPMiLZzCSj5UzNZNHbzD1jitGzU7IIoStOTVzhHzF6GVAhHtDakg
bxL2oU9jgGedSL+DNas+q4MFHSpaMdT87TU54z4m+RmZvzoIICggEr3owh8vPRhg8k0a42V3TqUO
g7QtVQwsYOkiOEBi9czXxG1IwH/QFEbI4IdgeB1ZFi7fnXOu2NT9qdHScra7mXnlvWFbiFpscwgb
rp6J2cilR0FylHosD99jy8sQhe5Buvl8EfZdwlm10N6c6WRpKFc0mcJrln53B5mfD4vBdpSsA3Oz
EL0PxF+Da3ACShnD2W+HjEN63eHzylw+aKq8+kiDtKoFJ7B0SpNdgNDARBMBFMjUwIoWYuSBO1PH
NflbuSyvFuPvi3Yg9o/GkMh0ISlQ5lNlsEXammhTuxKribno+tiEuOkkhDyfKHeNbqUusZQEH+qy
go30lCLEckJZXMGu24ahFYUoOJNrqiS/MbQerjjnE2g/UCKL2R3w6AcUEj6Yl8Zn7aWDJ91HVjda
Nu+QMlLlRFCDyyrlMZG2f2mTU1ZDEDRFVu0avhcjw9QcfUnCBC/IzX0tsJa1PIHZSdmjvejeFVn8
Vw2sz6yy/oZvyZVb5600hPUk7aLCez+f+QXiT3slKKN0JRG+OWxeUHqTWxLbmfN2uWOVRxycfbpj
/PKZb/mqK6W8hX0CXazOv2e9nE6h3zTeQSjwohpdJH0Ip1EvWnRlRL1s9Bqx80e7NglEB2k+voO+
X3ELk0o/SuwfMUkxGGStqMwQ682fzB8JQNu9LmbYZou73B3NpNVZhySlX93dCsMafJf/U0SEwCxT
bKoVl7dbzGZopRSrxV757zO7DVoHK/nMI0b2hu+5AHWxT5NTegqAsOxGPqLv5yZwOvXtQobRD8lC
Ta+SQsLth14TpzXFTM+lFG49AjvucsrMOAI4L0eLYRvxDcupAyeDKM5gTUinb8sIWSUeE6lFSNOI
bfs6qeB5PqfeChXHAyUSnYDI2JOav3tYxPowIwnCQ0fjEAVgX4mG5Kcm0GzxCDF5z+3bRYbxNMYH
Glsr/LL391OAtf3ldXFRSVwTNRmIaZAl90bbhFVVueCMH0mMO+cmd6+EtPNY9oWkSfKAImCZ4xgN
y3pUOwou8Ceb3W3SPhKsEC0s9R+QLtXYfo6Mdl2nSGgWaFm7OQm6MQbsu1N4mbwWkJMReWQp3BlM
Jkfi+mUW+SV19n0LKSpVGnsThM+vPjqKCSPDi0mfPzUqBiQAnXmx65Ws0pdrfrbzfmgRrL48ZHAp
Hl08ZY1l/9jDII6sFmt50UepcsbOo9VHNLOiy958gh+q1GHkwSaITy7y5enUIC5FJUMzcEQy2ln9
t8MmHNMxSzvTrNvNRnI3Gp/WT/WkrCbSXV7XFWEt+ID3a9Se2qxlWLOHKReIcuwyZqw7Vib6hEBm
w6RS3KMn3th6JwDYvfLoZXwkVBbyZHeGXf9jfVtkK9qBkBx9OhEoK3ud/iCwpccW0U45X31voW3s
bu3b9Bw1U56rgEzTAjL385CUXnRLn1ZH/j2qkwHxMaxjThOEE/DVo8xJMFCIKfE1Xf2eUXlRRLBK
cnMn2Li2Ao9NmublxphG/n2irWVW/Bju12w0nu3gcBeCqPJuoXW1iKwdgFapOJIaL9PL0akSEVOt
OSntNXxBnUasTboL6D/mOMwPHmBLWL3yLRtThm2DRJTeUgwg/uQ93tkjSPXO6wumcqigHQisI9f6
1e/4GZT8ihMMgFn1SSFQRZaCv/58RELpHwcLhbCRHXQHfmakRXq30Qkhq7zsWY8rosYWQnxFbm4m
a/yHx9zkPDHhuZKxGx8GpShr4sVlDCPtOIOlQO2Y+qZdpltuKIWaitT6YCvc+0lTFqR/5wej+VHh
XWQb8g9UPPaLKMWXgqSTlaED60MP8oadJ5MadB+LYYLtn/u6NAcvbefLmyRO5K1z4/XcmgPbZ4wY
I7gvibbaVadAKrWRr3oBLx+OR4YQ5UcD1WDYlWjLT45B
`protect end_protected

