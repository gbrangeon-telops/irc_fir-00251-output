

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SYUpj6do5sFTflpbsRmqzQKFPQDYrJyRQArefGItBrRpeTStPf4iOexrlL2KuY5Tjxr42gzfz2no
s00d/SuK7w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NR3ykkYMNFMRKu0xHAyt5DYiOktc2YTf1JOlIURJ/ThqHJccRXVvH+Sc3vg9x993epLj5za38fd9
R5dBjv9keX+G5g1u3CtBsdqXK+hNOz/uDIy23yxr7rHw0ImE57TmiDkVMvMwv3eYKhw+6jZKYes/
orVUKkqCIC9qrUn5RTg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HlVxjhtCNCKKX+WIZOv4bglrDneJvrVwpTadJxqH8bLj9DfFux8A76EOB2zOay/g3B51jEHFXs1k
cSPeVifBOPOW+4hnoJ3TimbzQC2WXDZLrgI3HV0zvi2+v+260AsNylQU2ks3dLwbxExBHvawkhdm
qLdLQIFdyzjRMD/G+fo3ZOpvx7tOdM4iBWXd2qur6t8wJth9ryhPu98XGfaQXlmJP7Tzn+0ub08s
DCWHug4G341eF+dWmcugGtWe2Ca08XjibeU1gRioez7LDJacBlMb+me+eJNl34Hg9trbjeo+4u2p
UhjBKGy0TbAWhSuuGKcCtfIFOUbYcwT6t2Yt0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DoI+R7m0zbJxCq9A8c+QbVnIsy2kNMG29/strbjpu4rQhHX3C2LKQKMwC4UXbs35yFBTN82oCtQE
LCzB557xK8srP2DUb2FdCBqlo4nmLOUDlZKHLRnMjMktj2MJoV0ExtbMFAErwe3zZqIBchZgf5Be
0C+OuuK2xw443onEGyA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jkJi3dDxF04M0w5noeJKvbYmN6cGn5suzWOH55jYT8k6r3UxrWZdHPmAWJgyGzXTFa2rcCzw1zFN
8CUT3mqhUaMicnmv3k1IZXtmQp8LLIMHIhFQWUBUexg49lQQHlMizPzJBAEcyMQJQl2JrQBPC4y3
FtPjOGWfsQSXXVoSz8O8MOKUSTmbuzqKeAR7KYOBiW1PqJBZo+vP/teWIw2p1h9/ADBVH7fQiL3s
cyUleDPcPx934u+grxqX5IGh+uK/gO42i4Ms1tDDhMblp6piYQ998xcC3XiMWw8hwmR+KGnfqU8Q
VD22eRbZMxNB+D8sxEO3PnV48eApa0h9wT+rpw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30848)
`protect data_block
N88tAffDVUGtijMHuKEkvGDfxq8Y87ERelIhL4xxU12pNDDXwZhSYrRxW1nDk95AHOyTTFAaj9KX
3E9JIUWCaW+50ZT/QS3u9afySNISuppcZGg1VU96vGFnEFRZoz0Zhnx5jKHUIcJFh70q2NIx/gPd
ZtC571NWPOG7n8/lommGa5818zVFBsZkR7PwTKJ2TVEt5xl8C24oZ5IRxJ7uGfouey3uboYvm542
y3iTDGKY/gs/1fud8BYvhKXhYuNP0Op/+6MvoeIYSKa57LDXj4vIWflDDXPckgWK/9lCrkb7hBS+
hk33s7KdLc/0qyVEzGg/N7cg9R69H5BCL+QEdBsAx0Ta2j4Nhwnxo5mhq8BPvbLQ5uUj7ndnvwMM
ukZ8pfiRqtHeGWsX2FUMhFBM3NVmUe577rbZECa/7xnSVgi22x8VVEdPc+ZISx15h24IOfLb1FHZ
krHxUHh6D9zIfzyIOu8tkqWEWXsgRuogvQHuEgoAetMh+ozDfu5aeAIhhHW3N8vBCkfVrYqiB0mq
CexgZqfxidT61CrOfmSLCZXgUikMXSWTG2d633JAB8dYUnXlNw4gB+o1S3kSFzrdqmxfkUc6YJqr
F9qjUrlbAQy3GLokGKXUoNQY8ZNbXdSIL5vmCOkXOMho0Yn9ot/VGwfH+7TWhjPisddN+Ex0youk
8iU0enNDYazUlrbD98yVTFg4vacWJKZlixU+qQFX969BWSK38xPbFsOFrOCbe4oEkgYx6AdT7Z58
s1xZGMXTDiE0xZpFgYkgk30GTrqEIAgoty5bttITlcfvPJ9mqTCHr0+fzK2FqIjDrKxfg3rJdoOm
zm0Oqt1baw3oIegsndqWzvtq+BXSPiCERCWIV3zW1bDSfNyb7X1svL1DsAPHL7FpWb/axLFjsvCN
lNvUUaQW+WKT6URZw+B9ASyA+1R8GoZUjyIvbv0I//9y1PiNmQ/+/SvodNoEYOYeoC8EFvPC8aQK
/qZx4JeD9vA8GM86YhXEXhKOZ5sBNHDW8DUN7f7LjzN/I1E2uTxGx2VZPrvhXb0B7/OM7J7iS+J1
ayr2rMaE0bD5qxWwvdVxR87oWCJIvv6/43PqtAMUBn1edEOV69bySfcajNgFW6tbCK0XEvWWrzEv
YVgEuT2pfbfmyYhOv0eHDhfbY+rCu9fCBbiCXeuKhAUbrBB2nnDRQUglfeYgQhHIOztOQz6UXknP
uoElg3NMVKujE+ch8llB7iIM5uUBq1/B8idJ4kmNkkcBaF3w0/k/vApmfSEXjvszoLpgKbZ8VezA
5XgS0GOsJUzUm/K8rfueJrlNUsGJZWtgx74wBENhNt87AZPgQbRJRB0uKrxMDURE84VeV6el9MuG
+/KLh/iChD+ytGIUTPUFBYEnvqyCno3yKFcqLcMeFbCVjO6SYa3jsW341bSrdSSbJHNSNdeuCs9p
e7bKAlSoKMUQtaLKMLwtZprP6XwOB+JWGMJYw6hmBIsbMztQqKZaSm8mld+HUkNLveoppxR8SKWo
FSNFVNq1VNsNsxIwUejU5QUf4/hQ1d5DV4h65uuUQ0g8ZcgWqwn7yxt6k8GatEnQzvWC5EhfvGzf
UDnoQ8LxpH+kqCBFFFSjL1uJq+LIKLjINRvvfzFqF+3TAijQAsxSRu/rZR1hSQjs9VZIBI0d0s1R
Owzz48IU5vreDWrIepqZd4rTW8yf0mUE4+q1K0gCNtQwRf3OMor/ZXb1CBvqQoEbpIleMbgKo1R0
GYiWUTLVAapbSozuYDBoD9d5+7sK244k5AU6jQcyFtN4fZN00caT6X1pomoRKfvF8AobNAtpvjF1
je0YFEiRU0d7mIrt7XAf/I66kiFsoqBZz1tYQCmIq+WnBBzXS8zMo1bOrQc5AHGRej8OcAgNGOK2
iEsdlBig3NENz23/+SPX5vbeslERZShPRIXbAI51EYOvK+aOKQ5JeYx4QOx54KY80GnlkCjCtO9O
3kp4gNYWKWLs2T0AfVIOggnSI1x4eDYEN/ighgJlL+96I5Bv8bPWhDfCkAO7QMfnkgvHMwrOGpZD
/gmg/UdGGtQ6TmsXEnGjqlsG063modqcseSrGREYAuM4NZT0LkTBnZ5hfE1diSaxPNkFQgAlUUZF
AEtMg+8yBx7sqREzxReaEh7CeTS3os8gwvyQDbRTdfrMrdDjA6pf4ny3sLEKgvDTxqlGWCXkpg+3
PT/3aDziHtL+Cc2Sf9wmDgA1YhGDgQ5OoJnFF85Z5esVqPRfKYYWDs8bLtcLaq+/yl6NW+83t4yh
pXamdhZQ4mfOD1mmNEDu8fFXTkei8mHYhoWZE7J7bjNai9uiI9NAhxQrlF5EcJSP/FRxYAIVT7UO
dSlvpkEeXofEyAS+I1H8dDiniq1Huwx9tAmkNhU9mrQHZAkMewntnkNlXa5FdUtzzPBqCKDEyE6E
WzO/z1wPB/36TKzwezdA12FtgYxmeDQribhk9+LudzmphiSsvwRi9BefbxVZphiGX7r82O73dq01
FwRx83Op9qaDAN7CGN3UknfqHrke2oSCbmRvOtZKDUt4MdHh9YM2ZsGEffHt9Y4rH4eAMZOd2hlz
mOZxrTLJtlCr3PRwXXhVCWZTOHoYg3eByh3zgtLYjicf/82BHlv9d6d0jgOxm6VIHFvV7Q1Gpo1U
iCLQVBsX68B4uej1SVf9qhRMqP2HCcygrI3DG19YB7UYrzVMjOfGoVoZbAoh76bteYrxsJC+cBUj
0d6fcPaBelYWl/qlf0P6A91M5yDuXxLdEBa1u2S1Hll8N77Q1THDLdzt9TrfVACqZulMn90lVURP
8TCaRhbyQAtm+FH+SIaCjRPzKr+tpNbqKzSbG3efTgRCuT/KW6JRhVQHANqRmz7fwukeZ7ykKOxH
rujvCA6s2jwQlJRzrQIWDnYsKRo7GQ36jDvi2ETfpkj3FcjDiOqfTpRYwd3VTbIR7L0YedjvUE5a
VDK3iUYvj+JSv9r5uqJGF3YgQeEv8koYdG71eDNM953l8awNWh9C/cXwxuYWAiWHoY4iF89CbLM9
rmuh9NQBuF6i72Fj+eet/KrU4bvR4DplOp4476iwMTnDTMYXAnAgPkhtHjIOEu+ricF2/dNYCgQe
iWyhmXTSeVecQ/3WgbCuPSb2oBm7Ee6y5XrfuOOC1TEioVACdq2HrKY2pEFA0WJ48Q7m2JnCEN3Z
5pacEJ5IrTbv45CT7C1hEcl8oa/sfb6XZJEZE5q3sTOLGC4b6u6nTCSnFnTyXSI9uWY3I+AWd1NL
W9r9RLawJPunzMM7rsEyG/sbvisQf+elOxm8Q3b+I7IcLoR9EW92dUWW6gwbh/uMat+nO/CEQTRS
821IW3AiK3nw7QU3XXeO1THgCFKs9VyMx6D891zeNDOX/FAFNA6HsPN67iYdMAWNej/0dA2U26Ye
5qHfwA3C0hXJLiXjhSMuBAAZGsyfFDG0t58qxNqVzLQhhxb3ky1f1mCcIZwIx/nnpUE6RXvqq+2A
zK/xFB9YAY0K3vvoR5yaCy6u8vEA1/Tx8FvU12RwydPtPpg176TBfSgZ1KMdySqYFM67coIidZ/6
AqB3HKHVu4CRjXZhbgO3WHjnNTHGN49orj1B/9lpwj6nMYT6F+gHVxeKRcvVo0oAMUWrLHvbHUgk
nFyKC9nj/z228GIliRLUk+B2RD3+U3VL/OPa8ZeJQMn8cn/s7d1DoyTyCu8ZL8xg2IKX2gQeoa1L
oRovn6fW44y6q479/Etp7SXfw0zDlJMQ/iV0uKwrHvnjTAugdQ4itW9kbCwmZlDlHwEZ8BMUQO23
eU08UvKAfkw8RsYsobX1m6PjmiV7cle9H9mwOBCZfD8PWPKMMR4L//EJyZLbTTcTjDOLyiTRMIGY
Q3XA8XreR41ihLRaM6VqHFPWrAcZRtxJ3EkJQ/T6OWEALjfz5WJ75x1kCYW/kTI6M+iwWVZSuc1N
0PUt0q41u0REZstmOWmvymAr4/bh2n8UH0lVFwvQ0V0vHjPHbs1GKJwtw/6fwky967LpRowcZoY1
+aafShszmykMJfefdu3ld8i82yM6GO1LNucIT150cagDSfgDENLwUjNFm9Xn4JeXsLmLvurF1Df9
SykrBdV8Sq/uo9oaS9jly0QoWxGpGefHQw/yCH4G33kS1FdAhLAYiQXbtlKjeX0CgslwW1FjnLqo
72NPWdHq2qg6OVS4/boBhLQ6ADi56d8qbKohNECRqzcV4b3pzN10O/KEeutgg+naVEg0VCrAQV+q
aanePM/bueV8OxZ7IlOqH+VSw2L+RCe2DDh0LbMYcAqtHZN0TUcUasZD5Cp6/nmcqvmBWuYc5zl7
+S/POotQFa0+bqHy+SepYsk6iXe5qt7hzRu7rmb6PW5cAz12+0tkfeqRIEUkIkLka2RmL+XhPUax
FwSLWy8lc05TtRv1YTJQQS9tcu+1tebKD1xJHHQOzR4Ygxo0BO/RTi1KJYx7Nz8fu7Of8dQw8rWa
/6rak+Cv8bTPJhZL1SaQmC4McvP7ST0l83vUJxXAjMy7/L1EifHiP8IydAaldUBDw/JCQczg9nQN
0WwUH0A3SzfDEcogxEgFTG934UeCq28czQ8DxzMeS366E7QOAZOGBVEJ9E9dF5Z8632eqfXj6/Fa
4Vl4GtqbKuedzq2cOPUwjqYlWvn5yy05yEB1c728P5keoalqnnUpYbZUOxEThl4RyESCYf0xJne5
vpmYKIleOlcuJ7oogUgm2AAkMb8qG9aiX6/K0/xkExcr2pYLvosBp0yMQDgsEsCmXTFAzs8sHp6o
qUClFLS65tkzzpoTLu00IWkZOses2puT9IEgK+3tLjCJcxosOqm3ob0oLHMNEjQORoa5P21Dt7Uw
n58M5v5xJ3P3B9eckuVrrPlY8JDE/06NO5MRTs0wnqXZiT2gTIzmwnC67/v526RxJ24uQ4gqt1SP
yqiSXO3k6dXyhWcuV28P+iVP1sZVBLQiGmCZAKs2upES9DfaO8+g5agutfjSktOkhYstoMGOjvDv
8b8OEMmZEnDjC2fN269iXotZQIms/Ohb5d62OIVOd8JTFH6ZNkGEoTi1XAobSpRp7VZX0koAjW2J
QwfaFbnTITE5lxehHVsrDb4CspJJs1xZ8NEn0D8QiqhtluSrYVOI3Q21zi4YPoKdghNTJpKGLHCr
5f98kiPWZfd34+Vs1fRATBTRnDeTR7uEvzXq1JZOMS4YVYqWeRIUeR6TEPmZxGlGUjycEvv0cy9G
sJwke4gYyrzQKiyndAhkydkR1e/IZMgEtBOrn2v57JlDAEq+2olt7k2er2vrjsSTRbMHuK/z2Elm
y6zbHLkbE7BN1TtYnb7Pb2/stAD+Qu8iLK/lv+07s+RadM9e9VMxNCXvmWI/iXvdLDUgcgB9w5yW
MUJPNSEq+geUVBnnMw9lRk7FDcILKp6xJsVcvxWoaj4xuIfQqfpglSAtNlKGsc/Ow6LL1EzuO8m3
vJWGF7cYOhbnjlyW03sabR/IpZJwmlyeFXiDnsP2eoq5kaXpzKa7Sg815jTq6+uf2Z/6sLOwI3GZ
uOvGU+cqRDZUu9jeE4PccZRnXBzNkwUF0+3RtE7SP+4AVxPFQCxvGDiQ4NgM+bJIBKwJ9R0PcbbK
Kz9PecvFck1MEYqGSQT83Wg67/b+quiYqm89WQnA0EmhMxaPnVRo7NDWSuKEma52xUnIgdUx065Z
dqKKxOMumSV3VxfPv8TQ4iUdKz32kZBWNpYStAV3KYqL72sOukmGm5io8dsBELeaiXs++3NCew9R
Yj8v2BxnhcmehSASAwv8iiRQSFiV0fSXn6lFfoJFrP2RkD3pE/IXIXn5cJC8OH+sYSIjQf7pH9QL
hep1rZ4dECM3kualhCxR8jlKUfCE9UK20qsJyMJdrmM/ijyUiOL9z9l5LVdYTGqoHOsBPaolHQ1R
Vpr3EhzB+1bFHViEQl8kZVFgcO85lHGuYKIIYyRgWAIBCe5/oUk+yb960rtTKnREKN0JkjprX0OZ
OPeziTJBmKatrWJ837KJYLOBn5De7mCN1de7is498VTlwVEukI/yeT3uJBzKuI38sB1PcBUcjcXJ
B8mW83FHJ7vITezFu7/UDtJ6kMWYOU3ATVDF7I5Nyhtz3auOq1pFqMzUVVOUSSO0MX9UJsDvnboI
/Slh+z61uZc9VS/avV9nHN8rinLhrB8cfcMUoQquHVeRjqntBVqh7rFsiqBJwiPax+1BQysDoIGv
7EfA13qtxFQMSj0U9ewKaac+miEotvu5ajNXrYlL1mIL6btDuoyR4/UtXerOgwPgFQM9C72sqgCr
1mQlgGfrnY5o9Bo+PF+Z7sXo69vnCKZF9ViMM0E7WoMsQ7+ZYA6kGFGGD0Y4CkNRFTP+PoLyj+Cb
YX9R2TKdn6IfNXG72qm+7GwlWQkVlJoTlV6p61aL1BH5vVBm7FCywAi7YdAx52L69AXodi4kN9Zv
jaC5dcTvZiMKSkQ0iyFPk+IDUUf6NhqoOwysCCi6+dOohKhEsY1vhzXi2KjCO1y+KotILFUk5BgH
oUYUzFNq1VpjRL3J3mzbULHVr8FpwB7cO4j+v0ou2EzdARUMfwWrq1vLUX1N3xrXbCAKqbLHDch5
uOMODDxy4xxD5RrpJT1XBgQRhdmtWDOvmz+iAiGiUUuiRYl7bKFNcJP2Tvd7NGgPDwqEsymVPgxR
OPq0ITxyhzmafL7YA1IFw/OtyMtCSRmLI8yeOkMMefyzJD4+ndwCvTjCd6Hf/dt6foAqzxKjepI+
ZSuHNWW7dzgezPDXLYelIJYlFJaUkeLVoJzS+/ALqdF4d5GMQCFlH6J5HcLAoRynjhPO6LavJfRd
aDZlCuQSFTH0/3GiXXZ1/Vx4ZCZ0EUmbWWA38osIMZ1s3qtLQ4XTYlocpuVSVsjAuLbw+XX5ESHm
IzN2o6ZhDuWqklEXGLoZw44cUj7la93C0+FpeB1qYsRKLGN1ktXNRG/ACVe+aAyC5Uw1JO0YcHSJ
IvnvkQwxCCuWFIBARztCqVBnTHzudWWMtENf3YNpDzgf040tbxcziMg3VSbJhKZT4QKeIleJvr7w
Gyd9T1gNDZXUZH1CGEPjMq8fAnZcK17/1ZP9UYjnBgFWWTtLt9JqTAUmMsZpNVBD2DcodEjWAmj4
Ul9+6i84yujppEmmjNb+qijc3mHkpYlqLz2mxI7NZCpUN7yRbP4V0yp/QD7+01ApuZvx1dFuwuRg
hVUGG95cc2j7kHEQW2oPnqWDiXxxaB0HdFwL1yKn0YzR9mdhjCBCxWsPSLOfyOLXxHMsg9E4xCzC
+Ik1DfQeN+F0BrD5RKZxAznHH0iDrfCV+zTJgyz+hwiNF+G2+5l1kCKcNwLaioXQrVcgmkJCWCBM
SSQ/82A9Obv0NEsLjrxZXgydQj1K9A2YouZnt0tPAjY4CvhBt278GcDxxHc0unOTOck7Lla2Ov5e
eRM2ZkRIWDd7f2Ovp4ayKr8A1H6hJZWAraP/9wNkao3yV6rQ/GgMgNuQ6i/sV6fs2SrOnSatNFzH
Nnr2HreQzNsBXUFRhvGmOIOt3oCQV67NDtjJq4c1CN0Jx7VFIWBf1mU7CnJ7aqP30DW4i/GPOJh3
IpUKIPwq8WgwUpOMC3ZZBho0XJrzs3qeyB2H4g/H7aYQhZCw8CloGV3XeTffysRE7RZPbi8SAJdP
hMH6pHC1pvp+z1vl9Dwhg0UdfKTDfYckzKrcJ0gIXKLaqWier5zSYgSncUGzkqQ82onmCsb5ib70
3igDFQxIIZN4HJOgkHygvBGn3IWo4aZiRWZtKlyYHDRrJuhzxKY+a0eTv3fwZ+lRIBymj3nFMVHJ
fJTbQw25OlpZglD7xb/+YDyy+Y8sXL00pgt9FcJJuzEHf3nQQ7HIv+SUnlmiWj7JgsTZpqwnMzQQ
PxPWDVEAGl0CBuNm43WGWGIuJa+PMtRYHDIaPh1O8A0EgLngSDTm3fknndNxzgzzoMZHzngTB8kW
++KRSVKOu8pyoqjXvTt5g4+XsFRUk/jOvhTJePsBMZ4dJ2DLU0qydviZDmS+dhI71gDGxjUtlckH
VJ+cdG3DEPzlQn4tEZ3Q4u5T3FOlFm1PNqaWLPrRGLMhMAd3jDb5Vk+xmeiltaDQC4Wi6CajHS8f
PcAOmIrHyLtCL/Die2GSqFZdtpyME/4307HnjGp9LKTKk17RWTN8UUnSZRU4vT3GaCgWaXlk/jb9
mr+M+Zn+9Po+v4I74vdV6scLOmumPrc9MpXGeebype2f3SaETAfSnH+JhwM73XYUAmn+xCE1fbKo
GpxE2X42u5UwJjy8hI7PO8F/SbJn4LWBmFiTgyhHg9u6SxfTJ6T11PIvVpoMtkZMxzkR49+9O8Ug
dQ69BqbrlisvnOp2NLsEvAFpe5iojbpw9GnSNRXGGymZiaahjc92Ki7+fjImI8bezmVefbQ8Y+Ca
NbprgeGRPbSGSBWVcIt4C0JIXGXF88enU33hlJXlOa41WRW/G5eRNhM2Y3gU+i7041KbijbSg/PM
vpkS2kLd8Snx34hB9Dn8UHpznqZ7XYvWGtbyWR89uSJWPCAyZFrGhWt6Z5J5/LOILsG8lgTwNems
Uh5203sSkYkSE9Ixga3tY4lSSnkeIbWFxtME/4+jRQM0R0B/H25U9bQf2TNqd8XJriyX6bF3IK0g
uixp6orr849SSXIHTzfoCsL5jM5nH+vHQuCNVSVYZYsqjVG7PcE2dQSiqqB8n0mfZ+VKO4pAw73m
mX/nQajyHjlY+Q2DEOl9SlGS1D/uptqSo6UVzdAbNMlqC9D3pH5dUG7g/+oHFW/9PlFtgDG6Pi50
FQ6Cu172HkR8bcqYLMIBmmAPRroAng1mUZVtVUj9PZBjW0ZlCDpQUvZIuFcFg5lJ2f3VbD/d5osp
mtAwhgWDcyWsCMBBliAHTPsa4Nh6R8TxyVUxrN80LPKOSj9reJ8yfrAuFZOhtEAbBqETjzBpA48J
/mmqKsvJpdlajuIK/9qMTQ0UlTZEndA0HgRnYQetz9qNbwIPuA5BOpnhMqeF9YdU6rc/cWa/B3PJ
2/hleDR3CGXdXKysdaBCnWJC/tXMYJ/nNqGNzIHHrbJE76TYRxUM/zpD0PQGmP7btVBDoJRjrH70
v0EvMRhneN7ipbgIhZOod2DBC30AHkzQwRY82W3QO4wwGAmyCWkRL5xVjZcQ1ie4xE8NQx5g23V+
B5o663CKVZbb7nYFNMfH9JDiw9TOIUq3p+CP59E8hoG96uS6W8KujnxbX9kvJlKghZsZSIJxtXPW
Kw257XSGr8HbYKW8XHEj8enu8A5ji/DJN01IweHTwKtXLh/p6vu3C7qN9gd7rPrbkgE34/Ndzg3O
az59hYBzCVCBV0UEeuysSS9L1eeuSUXDt5orsTXc56BfrKvqv0AjKnW2w+PvZ32Yi3s2+6EaNx6d
gZK4hPS2eGp5uBap4gm7b0IqJWwfrMR8cKLfNq52OtSBOr8oytM/LoCqm5B/5ydZ7OEiZcVWB4n1
XqZUDUf3omY5TyMQDw6QAqZKafc6+XBBRjhWMYxwA9XLJ5sL3x5jL5MhH76qyvWq4W3dR/7f3L0A
bqMlhoDOw4Jm8vDeDhnBgeyyb6annYEWd0QmJOVDoSoU9u4v40ezWkDRbCLhkYm3aewwAyKdetRg
FHCyZKP2y7+HiZoKDTkF992dYYmUcwl9wCowOl+uYAiryaZa2Y9VqleiUupZGTa3SKPU0VinpuJ1
PsxKYY/qaOhym6aYb3cYfB9vPbJ4GcAdmKqc4SLjwx46inoKWJfKxh+x/0H/Q6L+Ok36azu3kEoq
uKR+Uwukl5JZOrWvdositfFsuWA+ZK3NYoQNja6S9xLT5Dkd7D98XYCbFuEJ3LCGS8/H2phcy7SN
VXXJeG2QynsPtUqT1EOn/8TnUAYOQvywl4iwXzoo8F7yQDWGJ5Q9aErrHRofGiXnzGxzaHbxg4YR
tjrWkS2gWo9zhmBvH2DFkw5jKQ3ZHNEtxo6m1pXfyuE97dzc4bP9c+p+ycWWx3to431UVr81sB2i
eHQMR/SyswnjLb4gHVyN2cKya7bs6E5EEu7e9eALG8uqF8OubnNsgYNzXEtW3s+Xh/tHO/xy8zZv
0wWhPzCwYIp2AuNGsxAaSy/cP2GZRfUwBbsI6b1+V65osKGQ7m1Om9Rjvpb5sXjw3MogJXMlOp+i
F7ct5XConIbUSBEUPrK1aqvwUr6izbKKk9sqlx2L+gsxCjyi8QNNzlD/sS2VWXxeaXpgoFRO8wjJ
Gy048GmF8y0reh+wTh2EKgL+YBQqb7r0LD+pLaRfrFjZydiA3V0AYeHrOMfL/lpBljpo/W21x2dD
xVGxI2X4cHQiI2V25u5Us4y6vcZ8vQdoiU+pEUIab18RqJgaAd0cLsPmhHdiUMtJ8RxwYeRHcFMC
2FwWSNOrs5FPgHITrI6kAVvmJ2G6BKE27YPHOWSFOZuQXpj2/kIZ9qj4eecsfXE3L4OB1MzdTmOQ
xJSuiroJUM3kzwhdhJmOlLFHP+X2K0FyBQvI039MSla2vptizJH5Iz+AO+S805o9CTTdwKBmHhoT
emzxD8+rNkys6H/Fdywz+cUOmIKvPZy2H3noYT4sbSLIvQtI+F0eRVSs5ZAnnmPgd9/2L9rLiPZe
pcmObAzGYK8VFy/mC+jSVrmcJKdtpklu5VseWut+7oupqAs+AoCpQbLw4L4yNUzmbkLOGzS+sIsm
EZvpA9c3uF7YLOflVwBhj0U8iQaVGfKnOxWfG7sqyEVjC8XJINbdnQEjGOi+BPhNhM5IRRPj8hU3
rEeRs68NA0NN1T0aliBtc6bZD+ocC3uinRDc3YsvCXK1Le0EmB0xsz953J1oVEK63atn11oW0sga
oUlR1zCTYX+tNX7MkMwqK/5ckmXJzjgTnqwChndlDt3z86kB5iC/pD0n/f/A16lYAYrCSPw2aNFU
OcS/nmCTwbwIknfa3kWgzBQin3jsQqrxXwgVHYtPlKSOTKJo1PqdHEyztYA0vT4V1uYnqbzBotoV
y251El/0ARDtDvIYSOiSakJmAjasma3SdU11wh+BBbMEnnwKfofM1UsjYrm8kCYkW5dFtf8cxcJg
v1PzQ1vDDabPWayfCERq+vGyaAwFxFoz5FcGoIkIlfKSXhA/hqGLgCnAGMiK8qIuT5+bwmAfl5Qs
9UtZRKyMUhB6hYhky9y9A8S5lGrkpRZlmE4/TteWH6NjbFd5tuUo+gjfh4eGFYlpoon2txBA3OSg
QXFVDYvrp7TwjpNPIpGoReYGtT0uKnVd+wB2+YuNDeOm5fOnWIHP66V5NU+yCIy5oLIqHA8PdW5e
d+4kcyHPmt71lUP4niSQS/fqWkyMPs8njaApkOH68y1gS2NZ/WiHKhKxhf8cJqtOhNwL+65CPuXn
1jS7hysqyJKycTPmy28z+WAeJ+WPK+itujEX+EjbLQbG7Kt1V988M6Zb/ro4cC1PyklStgIjIEtc
VXk3+s9MJIiBaq3mzhsQ2EAbiuikcM9KVqkvyb58wAtjJquQFZxMwkZwQEDcXCpin0pzKjFEWRnO
Sv4l0hEzTSxvdz25KVXkAnNMFLlZ5hi5Cl+Okwv5z44VoHYgE/KjBfwOpkS7XxfoLFsovUy/W4xi
HlsQLS2Kbw08K4Heh8M0F/gVzfbxSYFZ+PKZlpCxN9hnJ8lhC/1frgvI5NWuDxouCHKX789QsX2Q
47bucEMR6XtDLbOLYdNyjt0lgCOAM2qKGkNZKUHt2XjryOkW4DnHoo+FKSs6wS7ApKE49gS2zljx
hlzeAJyV1bwRgWBbXjjbWqLpal/EIuE2gqQLxAxqLZ99kOsUC7aHDLnULzssBozxf18bjT46rdLc
20tKsV1GZK1HwjtKSrbmUtOd0VtFHopEC9lxxjAQ8fa1mzCY3Cijj/VorJAskRy6mKllGPfNmtGq
730Iz8txOWOmZqx3RAY5Iqc6hKrZ2vjdS/RPLgikdH3KMKO0EEumRqyf216yo43DtuAHRcfsJrDZ
lfj0s2vOgNJg2WgmiJ+slWhSKU14qu0/V9L4LShg3TNpJMlcPKZXFvbmjMd31A/BC281tR+g2qKX
RNxn3MLjLwhfHgEmVY2JivfLV95nNvt4uxLjdjii71paFkwFMbvhNXXxpDnY7F4Cb50Bs5aMBYmb
x25MYxG+Me14fcxX1/0YO5lreAQO1oQK+I24jUKqXxgqN+j6kZIxi87Tf3wfOEIYUKKtEIpWm3h4
2FZntlHu579o66o1EovpB7vJBwtQWQuax8i/H+yqyEfs67pah1cUV3VjuiFHTp2Xmpwt7Bc8dFiQ
GabzmzP6R0QzpXIqmyPZlgTaFCq2vR2Oz1Uj3R6nsHKs+SLtDHv2YLtot9qWHAIfAXGpdHi20YWz
xy1Q9qmI5qPd/7GZizIuVyzJ6Dsp/azFw6ZCg3dg5MUA/Uh4l3ieaw99gyK1S9tI+9QhlWF2eKay
6hLrCFDKDGH07viFe5V4n4yZxi6tmBBWn+AyMdNqt5h+0VW98fMgy83pA7ERmpUb+8V5Er2ChPIl
myRV2epIFp4SMcN0xPSLOIHWgx84Cm33hymQPX1QWl/WrMgNqiNZqNQveKeNvhDcmFJan3JHpr5B
wFJT228bGsklvYgBn9RoOXpbRQz38hkHLikU2M9rooNqRI2a7fkviR9hzkvR0hFCnhvdGTvBFKWQ
nGLA3lbKEYVnY4tSUDjtluve6zQIPh6+Wn+rXUMrqb3IZGd4TramcJA52TlVNSu61+xfHVmYpbV9
djZdTiT7vWYzaouy0XRc6xVjL2PD8utGCF7anqLjV6M3J13E3Kk6PknJv9hKuUA5cCzxflVpsyvZ
S4uDXIN0ogzZqls7yCuFNC5o1vt1UJJIKi4V3+8R/mZw1hBkAehuKRjHCy1SUqnFPTbjmagNUh3Q
oYIOsSkOMqEWlPDDV76FqwDh42fcRdlvQFzfsM1OF5MqtFZn2CNQ1/rWYPu/bMjXZPXGrRoIFLJ7
vBGVvE6j56U25YLPm01hhgnlzmaLv5XED4MsaFwDR8qqTlkKzxUGRKWfTU01yU0UgY1ISHwx2nPj
NtBimsUeB1cMAuNdWRmLgiRuv0fanormFXpe8skCjjHvTIf71UIyIhAfIxFOsjA7f9RDZ11R+97s
JLs8RSKqg94wvEgcMwrSTjRHN/OY7QkEgxjZrHhC/lIJnTTB+iP0n9ThBmlZzs4KgkPSg3IT0p5C
7CQnXN7Yw01MGrnkT0UHxT/U5tplk+Q1B542qdofDRUDxCIqbuTLVuE3ee/ZewYG/EpMFd3aQNpY
4zS/iFrAcWF91dpbtrAd6xdNYsqS87+Tk27ujg4qGeB7LPXOWw9Ds67anHb6zWWMeDL9vAUOXZPV
sLloknsJK4nyxghlom+Zz/nCtkHhr+TV92xATEI7t9oOWtjbeV3Hd+woVz0iiIHaw8/kMhKIoHXf
Wt2+0A4VKUQXtY5pBr+3BixhT44Vc44kXKsjgHVX3h1vLE+6KCDd/HifQ/23JQnYhyiFNyvs1y91
iMDcMCGppXeWV9uUumZdbjyJ+G4LO/q1Msju/Vax0IWqqOzEUk58hjF5YLr/gbdJElFGtIfPnIFV
dovMT9EuZUQ8fGSMcDn99FnikA/VfxiSaYeo+ZsKFBmpEUYyNCMsU1/myeK4tFFTzV2CSJH3D6b7
PmMfMj4lnHXabjTJHM4vcHQQCdp+xTK4vj9v8e3b0NfZ/mbY76wlQRZA4jbbuMIfeerMr1oC3KTt
4sgB77Gh2mxFEe1co9SYJ1lGCSQ1oCX4vqh+3k0dKeDw/WIRhnVLuU675K8Pdttty01Zti1xXE1G
6H+zCCDRGMVwQFzvmJPRtpe/YGVZ8GMAbFsDgP2D0W5JfHOJYn+u/W0jx3qG1YRybI6+qIroo+6Q
gr2nJd0q3wFPhk7o5aroKFOo1njJXmeHLjX8Eqpxwh5Cdp85VLrc4A2pqkzEEZmlp3tPndJueLlE
h3dZlGNrgIHsiqJdJnYxEuvfF7YvklXzFNBtqayc5apghpgVE2OYTZeh/RrWzFRLFWR6EquAO+xO
879qAayvaJ/UUYPidDKKb+FiYdRYapuRj7S0v+hD489xTEOKuOjAE75QDHlp126HvY2b2hzMkL0u
k8VzCmH2bBrmWdLOES3CtMj+kpHm/K8H+/eMyLXDGHxuYrek7YQCYKioiD+wuM9VhizEUH3cSqnf
gnb/jsZJ0tWJ91MfZMf6QravqWnRZ0yW7D/gQ3/hPXx6B9gd5FFNFyZDZ0xshsBvtfeZsPS4S2k+
qogs/z4hM0Y8370sXwtZG4WSlQwCUBsAPQ5VQTyG8UIOeipNKoWgUEDL8gCAv7UKYEOz2VCbrBb6
eCaPx/U3JzgSZfq6CAll14w734yC0Yx1Jv9q3jFKbRgyShpeMobAWAL/x+PGy5z2YXuSle1dO26I
uYMtqoXjPHdGQYaHYyNl3tISFkg99pRJK2skUeKHXlThkvl/irgO+26Wy+VWVBNSWH+K1GPhFyIr
LHaSdIAHCGefp/aeEeZKH4PMK4Xhfzva9JwNYireUSluSFmlVNDgJOelw6HAqvE6NUMTaqHDtEhO
hCiX5rnuI43CvhgjcMlcTTmpDvaEczg7k1vLqABwDc0ehc1DKTMaMkyLvzN0kDQ1QPMvzZGdjRUu
NaC4ndFtn+e9KtVLdIcSIFgdXqxCOd/c1FxtbaLehtvw2GsjXzgZDexvUY9ycxGQPBus2unq8+Qv
Wkty4DDjR105cXO4l28IPt05NhvUCAvKjSHBYGA7tZB2QqWRtcWLEMQLeIx/Z76kCSdWffJJdk2W
Cujl5Xd8+TccM6uwz++e6I3BYaTAOvbPL3CnkhOj+Wicu3i8q5hZIlzbD+yiEkw2UvtN/jED5Fi9
vRUWWtVQLsMDwOt0zaRbiDeHVrZgCqnuW7FESC6Gi8K2FfvKEDaOB0eT0Mtcen1QsNYiirRjiHy1
HMKpPzC2Dtr/NI8rJjujEPHHat246PG6+XvEwBrQi/6x7r8UFSqVIdREosExWF7KvpD79ak6BcqY
9CBBU20W+fNcao6eePy391NFA6SjKNOg8oixif0VVbMMhh2z0VvgncUkaWarclQ+qAqBiuAWtbpC
+suYzSDyIIkMGGl9tI6OaVMSKlLQXm9Vcci4EK99fqgzFhEaIxsI47iEmxLLkRMY/58aIRx6QI82
bzKhHfj15bad2V12oUbneicyeG36wFLY4cmRIVRYqwM10cgeKXnerEyAjV+8QNBGZk8xzAvt8Mc6
19gkEUBbey/DMDuENvasGCLQx5PGw2xCkaDEgTK6g9+LNi9r8fklxqes67NuYc6uKOCEgykniEJL
8v3naolFyTFlzRElfd03DyYEF5QlJo0b/GpP8pDu1lcEodjuYcm37RJJ/Bzl2Rn+mx3041bg111Y
4sZFs7XAC7PmeFjUInpegBw4HzYk1E2AVlKONfYcc/dJoZplvDCGiAjdzVrUDkae0Fk1TPXuxwJ5
ZBERgt5nNB8XTfxl3Is63lDth09d57TcYPnGgKDznZoTBvETW9x82SIDHs5P91lMFnn7yvwX0vTi
yi3QH8DYjWPCZni6le7kAJu4VqV+1ByKZhIbSsn9TbYevH3gofxO1+5KOdonaWvtGTYMIFz9fKuK
botw5IOL5bBqu2ZZDFFyr8eWxao06rUfYqwmAnck58T40LmxNiafKfGr2IyOEKmgdEcB1vnx32Np
oedhsqyUaccXYVhcnlbomGOKz70RIsvhBuHvzDp5VaF5JoobIY2Y0wihF+M1M8g269nJYD/7GfgA
obqPRZvK0PMMc8xNZz95J2TFc8PMMVGcakhfPdr+1DabLxznkSiPLM6KdJvTSqH4zRvLfD9jm+jY
MDnqt1JpZW7YQJbMLE8FLNW5U2GeYg6mA2BpB5FkqM5LwKcrolrQa8ecdmVA/a8oFlDmb+r+Whqo
tN0gL5fUDIMNCSyxiuyg5SmTsrPviTazlylvAAqbuZwth5zxCEn1b5/ebSoDOZiYv5nyt4JMnG3o
bKqwtHumg2ayjuY6v4ATyM+MdLbHx42a3G0sevdRNkve8V6xyF5bPPYGPPtHgt9fMyZ2wvWjoV1O
mlWs7rnnSqGnBOjNOHiqKajnR1TF10HBjn3dgsvfBHdF5lapPVSu6SQeXQ1KNx3jp1z86c2UALWX
wu/oFBMTr2liqRBBDQwvtMsHuYm2Sxrxof3CjwnA7+pBS+JHIvCeRi7nsMdfukqCmmGzBd14iqNk
1ncZxIFR7iP7NzVCcIZNeweAeMiaSJdzl40HoU7L8c8VsAOqdlQ6qE2mTGKhf+qMdbb6tEYMag0i
HGtFnyfnZZ2KSMJTwguiF4GJhk0ca6gU8wfWZD00yEOjgw/wDpZkjVi2umzj9HGFQIqq9eZBxG7G
3DYkfb+gI+eyvesMbVfww6UYwwucCSB6bXtqruzs9JwPmMPGofbMeIkhv4MDoL4TUwYuEQrQciRs
24/DhU1R0t15Txbjzimv1rByNBmyEmQL8fdEpvyFYOIXI/xnCtp6qkNfp2i0CV2jDesOv0v+SRka
4XnHYBYZHSsLc9CxTzId2ERtnJ+R02nQGdLtA+PkDxRMGyH/GPsZz4TV0IxfU03dmkTTRPcA51Hu
OFZ7I0nAjpkmN0EJPZij49KYZoKpx8hKke3Q18km8Y1owDmwqBQpuHduKISDqX5fqsLXBHrp0k0m
vBgQg8rKtKSjAf7UjB6SPcrK1UBuK3Do3GqKKNe9hR6Yu5RDt0hn5Wt9b/8m0mrEJICCbllkfHwf
MRuc2vm266O7jzZhnyJtOTyS3/6K/KMQ3KQ63Bzgazo/Q/i9R9Z6QyUSLugwphY9YsSh1imMUn5X
HJo5yzxQWR2uE+KM0SC0p22N6+/+ZV9kGjxjvq9z6zWoGQ3XmUy1SAFGTAro1qqczoV5+93t14yQ
1f2dAcf6YUKipwdXImYFO2o7ySLgW1ClmUERxiTx9ACS4cONjgLb8jMxJgXHeVxvubPJPXGs6H/Q
VXEP4clrBtKxD5wcmwalP8sHMKxdwiniVK9yZJ1BLjNJyOo9NPyA6vJMjvrZ5CRA6E2kaczm6MgK
mxA0nIAykfc1ofKJ0pEsO6Bo0mP5YpiOnObv3uZH/o8zuR1NDgGrvafH7GkgvGhyuL+ZOqs3FELC
5UKgkzbrvrTrcGF3hm26B80tVWIIg3DjlCOWTlVTJVpgOo/Ur3EZOVVYcFDrLzv4eIpmH+1wHaG3
c8tWNmdNlBtpanuQ7VIMUT9HaKQBNHHXvHb15Lix2j9inqXfYfL9bQ46fnYI1aaJv0vcf/RhylEH
lOJM1PUi5AMsI6tZIXu1A4+1sx6vqGKm4fR+7QGZpv9miG/xkxfRKAzIs9dzKNnJ0hB32wzI935R
kaE9NTvfbLHald2GSuqGDnF14+oF7vb4kLvVlUUQ2z5m6PLGK/D/I31ZkPLpcO3URojuBdqplhQi
Qje4GV2UL+usqujkmnYzsEZeTWyG9yiePIIGP+96IU9MNST+VqSEtoPRBBfuYOm0dTcM5WFfmRTt
MFAMg5nvlETx4ReAFAyNfx11Rpps12lzRZ2wmfimTzlmg7PleK2St5Ny/m2s1PbbvRFvnr1XVlHF
3N56XJx5uEpwO/ZBYvW7KdVsGXjmDmfxIbc31v6ffStEPzc8GgUVaeSD0LaWqWtTCNchEklrzJb0
Epgeq6YuHzFAaARx2aKBFwZWmYtC76Zs41savycZ1HUfKmfkOR8leRW31HGlWSplv1n1qqSm/xZX
lOW7cDSF5Ss2H+rCtHmmEu1fmQ+gHcin26RnajQQaoHtjwsqzB6KMjvJtv3r4tTLZEyLDLr2SgrH
V1uWfYpxkZF23RLWe9hNXjHj+COiwxgkCJcgtIEOK9+ZU3eciUnIxeNnCLw5qtvN0lpqh/fWyA6b
6wOe7T6zQqSHJ/0WDkbc7sId/XJ+reRj5vwa6jlq6XBtJlQYNKjUrpDyyOLNgmKk3her2jDwEDZz
9ZGIqTRPqk3DOo1uPTLL15rdz6wi20WI3scU+HYClC0BYHkr7wU9xhk3i62hLOCtFkk5wH2XVKXd
0UIaFerabyJ3mtvgx9cKEtIy765q8qCDmvD75Z0FqmPw0ZS72mUJ0PShUbRd3ElbT4I6zeVmbYax
Fjkv5JHZ3GWKemvbSFIKu5bzv9T2yzUr81F1SDdpzOR37BvXiTivhkiEQHHcgnAXCpnwv4xJ69Aw
JUEES9RMVSaJszkStruTMFGkl8Of2dufOnistGOWNZuvrxov2jjlHjgsebGpdi4x4JPP/gwxSh+8
WOz5ZmmfAIvQRMM1TNk9LC5AaR+WZjSKhaCbmDvT+tdw/SSx6zQTbWYCJr5WTaP1fYndUCOXNji5
91ecIy0dglCeAnPVZU5hwdp++VlPGRG3f7CPEXfmffmhWSRjSRkh9ufRdhT0EZ1deJEUvxtJ55ky
S0HtQWqhtmfXhE6PleZa2Fpb1DlUrgHQNjhmK5zdE3kcTXbKKdTzISpaWPCAX4CY8S6RAZ6D9QS/
EHZz6wPkTaefJRk/aKFnNp5O8F59As0p6cLCbx8Adn3mk/hS/cnnqZXuk6bevdJ5rBf2fGMgBDwN
woFNibRa71nU7PR5ldfg2BeNlDmQ2miniGZauy5gchHQQ0njR1S6PpMM/pv/WFcRhIqVEauiWj3C
c2SBqYfAVvGRtgB7VA5xzHBFANd3yHVa2BNDbNV4YYhrWvsvEV/QNWWFmPggNwoOoMjnVfN1zlZh
xXT8vyEt+kvxr2NSsDIb2AcKkR6ahYprWA0c1eHtRxKGDjO6c1R0nhieTRdRtWEjaRjZfJJ1+5cy
eK/idi4hFddgLw2tpxq8kl8Qc/P6D4e1DNLs5VurQPBupK+/Tep0jP00Skv9NFODgXH44sVs27Is
HhR6kfXv3S1QuC8sijjoIvp1M6YKKBcoJrhmwFM6wE7r2Va03CnCnDFkNZCPlS/8ycFvGylN0LBP
LSMq7eDScOD42DslxHaS5KsbbfXJObnTSjzguK177tJJshC2iZEV0SmIYXf6wVXKuJsj+mHFgBBz
V5eVy+1zBpeS57cp8kVQI2GGN8p97c0uSoKZTge9qQ/RPm6Qy2cmR0l0TOPWb0zmEB+dzUyeJd5C
UrKU5c5YmpjeR1eIWyDo3Xni4zNgSqlOz2lgF8zzyODwW2wNsgOUStBGEmVFyup9YSxlGhMiSzhQ
6OP5USuQPovRLHoo449/aykJGCEcJUEBfKDWUTJNMYB9XCcRx47IIfOV7Jg4pAPvKZ8Ud0l+NOMT
5j0iIzzEs5iQ4dE3E5W+zQwEaBCwFKieEmUO9Upoj4KPuJwPCRYtWnux+m2/xlAxqnKQCq1Bh0th
vhdJoedUP4msVk5T53DHZZUM6eNi8HgaPOp4U/1wZuJxGzvl5yA6VgfBqPaOUULtz4BmpP1MKVOJ
LGfcjoXofOkcoVLV1Rl2+KR8eHRvfnYQRIpgUkCSOEyyzWwpYNNhb38EJDg72woFlI+GfkgfGycp
7qxF6dHhVa5A30UHWvHkYr3s7ZuHj1kMy8JgCbG6KTT/NU0mLFUPd6yhl/1IXY5Zww7PFONH1Ekx
OHHJwegBFOaWjGhyPTy6bv5Mn6fFoBwZW2eQ2GmeR4JZCGaChG+y35p1aAKYD0lHnRsNALkO9myE
Au0y5yfS9SYSnTl6qWVfc996tRgzZtPKj1kF+pnU8mSGRkrsnvpaERNSnYbncfiYmf+XeaQ/IZoX
FTDWeyx+Aw29jp6TKbX/izJRqvxket6KundbSGABxShXnkYSovrwGHPL8XAR+Xg5XSvOTFn2vDMC
okDiWpsJ94wl8cDGcEpBSbRsopBqpNeg/NHZlwAcI9BTrXEaayHpz3GOSUpigbA+lz8IFtXxo/Rn
x+oBJYmgDGCwnYqTtekDA3nDMeQsH5oP3Q1fW56GmG8swDCmdawxXienaUVk8HpptUeAK0ZMejoL
O63/NJfk1QVSoQU1UBnI1a+a6RML8u0foQCuBP3cCp1LOFz3ACA2HVKeobMKIWUNmiINWIT0uHnB
Y2MaYk0ArhiQKfpTSCGGIU1i26F/ZqO6H/3ugHyh6T1zelFCsI4o6qHR82lqNdv9tnYExGCcFOkt
Rdjtuu9RtSKTTYRn0VEk4aTgqp+wunndst8IRlZ7g2MT94q/bd+7ftb90B4FWtn+Vt6iLht3iPyj
IVnA4Hj9ZjU83ISJxJlkogf++lao+yNxXmbBAJdYYZXCIXmaKr9mbh+yg4mBAEkl04GuVH8XmL3A
m2BWGu2r7SASbRUyajzACY+q9OhwfS5Yp4TyV30xfhLGZqUhP4D+61vmmLmSJQCpoGZ3hlyPENpH
ugEIEEpgAv8vYy8K5sqyUKcDxqftGmpmekYJP+vZnwRxEq+ygEIneFbqTRX3by35PI9m3E5ZEEBH
L5ddUz3A2sykbpbL4fOgLXYcANaNvu4AfQTa9XLAsH7DR7rlNDjfRPQ7+kpy1g8zA5J9w5mOQE5B
gmdkTB9VZq7BXQSyaYx5hPoBeRB/tYW5wnN2vc1I6fjTG83BxT1irDoMsrCnqwBJSphbTFWlBgDS
+CSX8rfmWOSYbUiSvxnNaGf0t0x1CwY6FXQizEU0ZTIUpYBw0UQaKxz9Ky24+X/RQT0FUhygKRDN
RMnyDGz1cyZyNTyvL63uSjmqm6Y8xhw3uTU4quuxB8LKoxgkv2ew0c7+sdL9Ss0OUMontDoKxZjs
tuBMvjtNcmLA1+Vf6VCDYfrzqf7VIlpYXw5Eha1YwWBrLj4lYBhRGXaOjN37HNsumxNaHPYHyWVG
mgqNDOkXnp6gUsxdSzAR8jwAU56cwalH5C9tQR0enm8IRY2PGCce/LCXLe6V59aqs9X/Q+lhTlFW
fVuPAfCxPE1CmzQMgAiX2+MhdL9/xoBr3WrPP8PSdTrXEHhNdmJ/Qk2Nmx0rkdmq5Hj3gBGkijPM
zg4RtafN8gehBRd33aSlRSlJjK+vSgh8MZHxaybIDtsm4AT/F2P2r/MD3bvncZYSHj/N4YcYjGzp
GBXXReOOExllvTeGvXM++RsADwP5rNhiWss6/oJHuTNMeCQ5WMRGa+IxqlYTgKTZUuQtueq42lQw
O1lHtHThVxE5Dh3Ak1s7MwJgBB/3y+X668rafThnVFAa3kIs51Ev1d4q7N3fK3iDOT8VjcYbTwnk
kv67kuwDwUMN6jkmnUzAEXubfKNqKPa1x+5zZppxdlK1AAmr1Hjz1PxOTiL3tXAqzAA9h0IlaCsq
T0zPNEh8iFvC3/k7iNTSisBjGeiW4lhCYQF4ktqUBQni/J8U6D6fFipHlgLEaBvF+NFZUd4f+Ow2
gRIf6thQyL9U3qWgfFb1IZ6FkNpBDQEJst4yC7mR6iLXX+f939Atb0kn3U/zBLsRr19wgWkSSuo3
EWpMExlGFV5dVBcQmHwYql2E+nxxW24B44DGn2g2Ll0Hpm7pp3JLm4pPzLo/KBF8d0OSSChonCmO
8ahE9tfYIGFtHFXBuV5S2xNfGBTfWdHNe9WqURqDlwZgJayJU2C/kT2FZsCZzmRBn6TCmcwIHJUs
jCtEyisGQnL45l0R7l/B2QIdHFYnEnfTWsuLqfwTfKVrNPF6EJ2CLKmzypwQn1e6vI+7C49Ofi+P
CBZ9EOSUQ0SvHB6Mc0FPpB127uHuAXlH62kIZNouZzODcEn+jfgcr852raWMuw0j6eW4T2zghNXN
DkkNb9Qu65tABt1NhNwHYkwNKZFMHkdGwa6U/O1pvyK+xcmloTykLBF0U3DV0aUoGEEsrl/cJeoa
Ztc/3utB/PgWnt5uGPJt+C7lafbuW8YM1YJpo1BFCWsvmbVCBlp5gP56vChmEJWq5794mK9onISd
Wi+6HkYKG+BFzEs5q4D0WNr8o6u9OXdeoxytMqH8FAZXUGY2SjIYtEvutnJNyEthLJX6kGUG75XO
cQnnHy2pBYhfd1Sv4R1QTgpceD9abVSWdrNBZqDcPcQUj6FxQixsakefpalLfc373Lbj2EK+px3f
jWCsr0Scue0YI0hOU6+jeVklyIKnj+l9gWt7Ll1G6rd+9c/FQYC2H8W8iEpPkTNRF8oNP1pWSOb0
uiBcKkJ/1wAfCnSrzyl0EY/fjREZUbVU35NHgobw33nFyl9ZH/mi1/+R5kDzmB9DY0WD/t+lNbr7
9kRFw7MiHdgJ4UHb3Fwy5pnWPqpXoQLJJJrxALnLmm/qP188T/lXtnLfn8Nt/8mTMa5ycsaoyjL4
TRs7Jv11Ji34qXGG7i+12mOyhKMCRQ6E1BtLDuBkZ/q9F/5sRG6QvObSyE1xTtQ6XdrHqTerQm6p
Q7vEfd/GtyTPqQ5iFcDN/vcssLKAFoq++C5bsV3rt0xZQ2hnVB+mH7OPg6PuuTX1uWA9RfosHSpO
CrcPgsZooJiVAnYy8OVmCW9CB1myGcygpjyTsh+9n1y61VFSUVZxMG6o7fU/UHhe/ZaTj/eLLGeP
BjU1fcXLCqO1gjiqAP+qlVcLxQT+RZ7LzwR8UDN8gwcPwKMwNhyVqPipArLGwGnsCXawk9BBoO/f
HE3B0tjPQ2JzpQAEkTMnOlLZK3LPVfhQOLG+oHZStYOJ44PBclKsomIGm6y8qRzpjnzO+vjTb89a
tOCqXmCWXT8MC5Z1lv8ekyVz6m5M0ajeOGZ6Ltc3NeNRo7Lbq4h7OxE5A1x1IzcY794kiTaKacTZ
w1PYuWtGerDcoe+4Ibd5P1O51WNXzYDoagJKUz0tqduJiogP66SYN+6wN8kOG9AymjFPTQ9+beQd
figQKRrpa5hp+eeMcX3xm6vvYpB7THuEo7Uk2L3+haXUHF/XynsXkDwrd5Rjj2P/jo7UpX3JfR2D
XK42LuGI5ZjHz85UqC/tgfLIv/ls7n9xSpDAzdpKLAc6qjlvbW7IrNwrcwL91MPZGXqFuMvLOEHV
iYEELhdXYVq5rFszoTAssIcqhsm5d7xDmhCUU1eZ+bX/Mh4w73WYopq1due0HNm/wFYj3Q40ZK6N
bdAB16SCtRctee/Yjc06/lr9Dhr1qDZ+4FBPZNxuYT50YG1VEVyCKCvh4I/zYPqM5VENEbnT6QGk
+sY4W+PC53rvrA+L8dLCPhRPxZVC6a8Jgev5PidfO36eLczbAmRoDR2t451Y1UU7PIC0/c6DwDgC
B1auDkA2JonpnKTFO6okoyCbEBeMiNWIWf1JT+q69i1bzJIbdASVXsK5wJmh1mxvVDqM5xC14EBh
kgCRVL+odWVsYUZqMvAmHLJX3UZcCjSIXK9/9z/MCKT+bZhyp6iorQSLZ3Ap/lsoRPwCJz1EliSQ
bRW9toXanvvHkxZtquiQN7bQjFDMNxjbNXb8wP0emZJcZgiNWdeyAmfVJIvY1uNrfy8QTPOREVds
alELeNSkWfqpLGjKVlwT1LhjnLU+OBuWChP5ChOsJFffW3FwuzYz0BxQWaU73VnFb1xOuWauzqGK
IzZWUst7U1eWKogouCp8r2OU3fnK7YSetbpIMrODLZ2+tI7sBQKIFHwyE33MHcCYCDHDbv+frnVs
GuovOXtON5UTg8/m+i4CHeT/qw38F10NN0vXSc6+TxHBs0sFSmlNIugFjUbs7cqfRdh4OrbZFI7w
SGl8fMMP551LobWquFW7U0QDVebOX7C+pnbA8g1Eue2FQA4Y60OdgkymmyYZpWhcxgrdUzKwlNP1
UBfkyxlsqjcyFWTSE07JjHof0pcOdjYmQkEPt9jLRG0N96TvOA3u6B12M3B/8YfnqNKIUc7kWrJ+
R7lAxrpKTFL1w9VlQ6es0QGpHZW+XkLsz4kSHcBUGCt+Vm8Cnwv2hM76LKRtVqOiSofDHluMQRxI
Ddlz/kex4IMy3q2apfGWFLxd5p8vKrdvKHa2l2oZAwwodJ7M6zb0lhl9XbjHDYv9JsNLhepeYscv
wyBBtLVL/nwg6R8Yat9zmW2HAAbgTTbwAxJO5AQq/z7yM5iCeqBobSrUvk1EBsLkNOYIfLxQzbFk
1kZw6BWvFHQ0O8kDqvBtn9mB5496Y6F481iQDfV5zvAeK9qL3UvvtGhafDJGm8NvzZbt/zRKinxZ
t/vnzDQHIJvh22V5TPclml2WUguEs0ZGv6pPWfCx5WOsuKXPkZZ1wjSvWQCEdzYcX5N6Z5Pvoxed
RDBR5ipiA9pM0yYXzFK0Ph8KK4TKoeXnfZ1vqvnZiiDRun0F/CZaMU7UWJgl5N864nsDjLC5Zu55
J4bwL6plJpymvXBRXfG9YCeryIvLmWCYzw8GsgtdVaLEoAeu7iXB7XxP40HsrEl+dcTDxt7emlFy
97fS/MOmToIzi0W0Y2ZWkcBD6oWHs6AxL0Efh0zWRj1S/zpbNmAoOSoeVh5Uv3XJsTrH6RbrV9xX
XIMNP11+gK1zlXLeThVcNL8myZ+mhxr4aGNBVbahOjgv88wQP836lKi4T/Uh50vGmsaBqKrkayLR
Aif28B5jSC6Ob8ugqGTOpFv/0smE2S0xulEuoMmOVEFd5NVAhrkqxKCFo6erseuv8YZVXqZiGAiV
R22LYKQBaBUrCdu85buw9fUeOIOYygCHtYKfmHlv1OERyvqC5GJNZFDlrheKqhZlbMu+yfQsIYhg
4YBP70FwOI8XV7voHk0bT/ahM2T4MjGW8Htk76M8VDuFpFRCkKeiK4PUjA5VBlzizSOl44lzlfXW
BSBq1/xGOBGCussbQnHzNs/ohM6KLu42T5GnXCkC/cvoAIj6li+D12cicUkom8+g1tkrJ/BMCqVC
4leDKrwNCQplHZFDfQ7Hk1uE54lmZZtxbVeNHoWRZE+RcdNLgh5u3MALR9PMxbQoo3xMioXE9SaR
9fAyrCs/KbgMVW8VDImKOtnePBxiybnirJpgQArqdP2EzKxE/cVvDX0jdDWohg/H6xljAc0XOW31
+boU0aHDhFrIF/juGztQvwoa1iM9DQbREaf5mZ0jWBX5Poan1qWMZZp0unmyCGHWAzG0UxlEz3C9
Uk8EyrjwB8URAe9IFSIWkQpK6v8yEhocLFDZ7uKrzg3uswAw2gUAwbKTnGJh5AFhcps+mcXUgL5K
/kzEjP9fwrJUD6ZpdlRmdG007YfPyL/avLxzDmJdGMdCmSCZU8BfPAnChI5doQKueMra3jYeVnbF
v6pGFIxpM/PBBVlc/8Be8BTu7m3408Eb2isdQG0/7+kFN94z+b7CyobehAXOiVZ8lfU1RGUDIfey
pyikYrEpO5xb1gAoh3SON6Wktc7h9hoIfDWqZCK9hIMm5xWeH2QL3OSZ86PVsEBBPyPkMToVGdJi
oIglF1Sxa9dJoFB+rfNWwCqXLhDykwb9Ep2ps2Af4ZW+JK9NadSiBQnqndKa7++a0W5cXvCVnCjD
ncMe+T4PijKeNqZCu+UPcocA2snzby38WvCRpAwnrB2kXo5HQUOVYGZn6U7pxLN8DYu3wu9Zxbbc
M69hXUrK1/nMCtsLlDsn4jSzncv/Es3lR3Ah1NpluAUv8UECb/tjo1HaeqkcCkO0m5msk+BZT522
er8l7h3e3xjBX1BFdaEZaDzJ5yFt4snNvjj14r09BN7FDlPO20BorY4+E/YwQObax58MwEDL7hk+
NJ7zmck8zUEsv+/uEGRRHX9KFLW7CTxMjwbXpom3x3rWlPwjFXrP9X9e3RP4E7iSZnDOauq/u2Xu
rw8eiJw3+rZFEigA5TNC+jxgxWEGj/d3CcYy18ckvaYKrKtVusPpEyIAa6Na5zhVrHhc/JtdjwBl
4BEEBaUA6NzRXM8+hySVwXoreVdJZpNuzHyPltHo3rNf+fabqeLS0HlnaBGngcPSnxcQsCWlObOu
1lnj/9EXGvId7Y2/DazVSIZL6mTZSp6sKZuCCBFIhgYsUBEuI+pyB+esy8zbxFNK13JKbs9eNLgy
QZVM5M4AsNWigE2y0dY2EJLNfCZDPhtBFKl87Gmu2QjZmB4PSqeF/yY6OiDS1S3eZZ29Exsd2fX0
9G/DHMvxM9hFRyzo/WlgTJYeUvzlg2BrO/Mfbj+IFfM+ExvD4RTNxVqWK4cjrK6pnTgby5QwLbGA
BLOxKRS0veb40bgThAOwg5P6tL/K7XKPcyiQrAb8OojENL8pYyR1SZjs0FljYw6zVUriQlOGmqp9
HkuJUWakyIJFn1BQkzkw/ljjnMgKzUIxKJ9PatW2Y9miJShJFnPMj9Rm+ruZinBxQqgIbJcjeFLp
MSkD6/6Fzbhq7oxCP+7rW6PrPUmXJPmK3yc6fnDjrGMqs/5fu6E8+TDw1A189OyE7GM1Ul1sxW/K
ORruS+USMgO5VuZFck0lrPQMgQg1AngUnYM1+CLFWzc/z4JiQX+KASst4g+BzZFO+v+artYr5Gw6
fUhYpE3+1tiX3kSrMzK9gUf8ufAtvNMmP8LHY093iaZpRoIb53ctGMPA8BI9BLOzr85/tZrzNAZW
0gUpQo+tTyFFhyZgjfasRTYpOCS/vTLy5hehymIyDDMjTr8BxVndcZ/uTEd2C0ZgTDw75mXE/Wfn
q1sYtuZpYhtXLd7QCZRxLwJcDLswe7KZmvnCo4srRDdwcHdJ4X228KBSDOM9hrjURBVc21ATifsC
sSC7jYPZB674VfAe+lEc23fW/Ev/DWHlhSNPkr2JyNG1CEfhKGXFLtpx/qjX6a5pj0j4kmwQpvao
QOla8tZ51+WSU2KecG8mjeZMXzOi3slsAP8go94YRerGLkthSap4Qjl7Ng2jP+MGDjcdFhRHerLL
k539dOByLkbAjZWys8GhgPNYwN7yc630ZEHovzCtm4QVmS6igd64l/Pygu3IY3ONInFbHS6fhU+s
lAqp3CjZ0j8ihgz8wu6oKydpBBeW96QMxkVchm/Fwai5+58oPDW/Wfty7F8KNkdB7AittImq6xIB
UI/4zq79ZWCCV7796gkEOeyA5dJZDwqCNN7HjMliB9hA7ARR77Toec6a9n4u00Q0DtCzcEX29sKL
gahE9iBaPE0m2gj0wWsJi0UKC/5IGIMwFrCFNllYTnxbq5IOVXXNBPhok74bCHIItPyMQS5nfP1D
NhbZe5YPLOoW1f16KPdE6V07KHehEBhdONB7uCwVxUicrZKgh78esXjj8hKmubfh7AHCRSy8pjFY
CDySnGGaqcj12EBGC7apw2NlcX9MJL72CAKMVo+L2BsfKHZWImD77ZgD8pcFoUoZDaJ42gPG2Sks
KteUklpvBikTCAktCnOAzeM3p0zO04v7hUhiRPByCMl2uZKmjpUBsw2W3cJRKl20WZncwHsqqkM9
JVNqpnB5n4XmJzV9zOFRKohGQ8f7va6dsTW9TFXYuFcgS6NCx+DOr61bPRYR7yVgO2owssfaGDAZ
9wAvNtonSZpl0B6dROE33fOQnhVIMZKoTyjIeEq6HPoXQ/FJ0ITCcOSBVXzj1BYkUq4Z/HzS8umF
M5zNjHMmoK45m8eSTREJRM2XB0UrkZuSTjiJs/fBwNWv1zGQHhAvbsrQJ/wPtv0P8QGM2p9BDzuB
eD31ue2TNuzKhtRtxm7t+BmJbhtJsvtCBcOBWZmn6eLx+YjDqRi9hGsza7L1ePyiFShjgMm45yWS
4u7Ap+hjljd+WCLjMpM2bQZmTRv4UmX+Bw9lKmZBu/4Y2vCA7H5JSxieXrl9u1U4dxQPEiM1YcIO
b0zVZyURrVhmtOS63JO0aC+t3tOf5qezYXIGjHTHEtzexqc7rckykNAqFXua866pjnFWMljsv1tA
8D8st8wEsNdXtZY7VHbdnwgV+wXoK9dWyQj+WIPU/RiItQxha7i7ThGGXAvNL1/cFSEGeipUx25K
nMp42UBpFzj2eRgZKCS30BVkwccEiCSfOOEnnzWM0aIPaEjpILEGuKOBpyLXZyTpA0/mswLSMaqH
qvUAVQoStI8zrNTDTpN1kJAtn8PnKxtVMl7/nvMuwRh3mch9G4dTxTVA+GKOsCaqAXovsoXcqyQ1
d7UFko87IpO8c2UW/gZHIeldCaTUsGEeTSCriNvDguzxElkviUqr3OHMhV/gIQ3R/auK+Tqjr5K5
LIuGy2T5b4IeItSHOaX/4nyfEanMB56kE1PGVqB3GLBbNYTFL5aAs42zpYSX11MlQnnVJ4ay/Gf+
2U8LZhEFKzWsKX7eEkc9xm74azCUjwNgkMnXX83MlvkP2mHyO2BkfUxDj0atY6X7s6g+7aUR6/Ge
2JmvlfFNKVRFoZyxmTOLekJEFq+MSAiOBOmrfVtn1p2DcxTRu4XSaGr2rbqOsi1q0n7dR38tW0/W
+Qfti7ycPE+deBMpHakGYZGAfYF502T1mHne6iZ9cdxgaahklcFyWHLtDnvpJdXYKcZpysQyn8wR
hCLjWWslg43ANhcZNiqvm1ePRZ+btaekWkpk6QrYbtpQ5kfIX0L8QRkiOBVdFhGRmLn3YkC/mV0p
JKFqM1Lzx8BxFageweQIUuMhA7uuqdFwflTzJtTsI8VUKL926yRkJd2lb58jNhdtAE0pPuK6e2/p
d/T1vpSjOIF7A+q/lNjuBab19ErRWtSvZYww46QASzKPGBI9K46NJWJglT+5aFXGJrSeOGgdPYdZ
OmJRoWWi/mGXPt6jfOv+NEY+AionHqJ1fn3SAIQ8Dw6U+hhQd4g6XsmacjRZvaH0WVhjIYLnoOjS
aAzRpzXNaIJdnNg92iViaZGI/3sURQPGF5NebS+uyD3JnnfHNRd1lUNiYC9rE+bzaSmGryFlcZtJ
p0nB2RLVS6kDVFIdauSW1Uh32iPk7OUy3UsRFJBz1OKqEYUH/x5fycM4racNz6A1/GUMC/mlPV69
6561j6dvmyQ1NcWZEftW6lpBWs/ZybQdcSd0H6nXbTXtKL89AE216aa7dvIfdqjZHep08scH2hXU
Kd2IaorZaqCzn4zWLx1ufuz1jrRploAGLoavgEqesqY8tU4sHvXoJ8pu6Ek3lufcZzC9thkf3mN2
UEymiflbw9SaZt1glqiWf/PwlclwJG+KLi/2UZemVZ96QdnUfehdDGqicoJXi009goSrMo58e27S
HG/giJmwoeLvi92BO4Bzcj7FbzoIVQvsyHu5lWolYDLeE5XngFAF82VKczsx5JIC2DCpGpYTT68U
gUk1NTSQLv97rDtmhmBmyWuoxeFEN73cz+pSPmb45FVsNu4k58UDp60iTKwozOweB6IqoaHzHDXW
mSkC9kgEQiTQGKUJgyMoqNUUSQDKoDbAiiSG5Wvq11BzU0T3GIXu1yStSMxUfRXCN219zGe/r2Xl
zm5Y35h/khD0DoZ3OkvOALrdG8L4efwEPiRJTuS/2uHGlpXmLf8I2xobjY1oj3UekKX9j8A0mEX9
wxr2RkBi2Q2K4bfRXWRQwV0Vwi78e6GSXbhgD7/3j1dzOIItmrOvotaFmjLZLqLvhRXqmmXJdbX7
WJZBWDCImxrzUq6BglbOYYN+809eOmB2tBzy90yk7VaeZBa9Q9OBFOvO926hqZfafmA98ZWejjpS
21SWTdfmscjnPWB3xt8NWjTj1FUgZGPUaEWB7OttUTOl2dgyKt1GEUTbktw8amJhO9Lrj1pjZkxs
IRIE6i3FhwNdxpUzx4RBLGP9E3c2ucHdgs7zSPG461hAe7iTvs6m5eQ1MsCtwk1FaG9UQvjBzt8S
Jxb6wVx+r0WLx4aemJ7qDwD4sioKVV+1C2H78ZzYsQZNjm/Wi2epGlvkZcWHF+f9ZlbnrHcFS/wD
qYMnfqAq4AMod/+mS++lXlDkEwlZmAKUSRMul8pRSgiTQhERO/DRNFq7RAy3TJE1o42oYVlnJzH/
4ggNS8sm8QujeqRq7Vx9GARlQ0AA6MQLJQo5VX4PYO6W45qoJOK8+OsmCHpXyYOgZETrIZm1r3u1
6VOFPlVOh8roDW/eRNGHb4NslJiPGwUr3Ov2bfw2Bz37GRcRf6ldIfa6kqknQVDSZsU45O7pxqVf
jWCtJVZ+vAsFnm11vMXZWPkLM9SxxWO7ntuLYX4CQNoztMdDC/96Ry9AGHGlsSyIvsBaRzCJe16q
M7cTgi9xr7qg7JNizURlJvbzwZKSd/3ryttySgx/vHndjPBVE5ihU3eUuZ+texN7jpcFK9rNysc/
uuHT2Soj0iqhS0zbP6ts59e7PwTEygjFv+AGyBHQ8SoGz3a1C6t7VEo5yBHPEW56+JYD0HuaxLPY
prD6w80UuwJhryDhOrMotN7lnsL/qoLzyypfsiAlBQrS/asyhLrqrHd2A/4NYyq8rgKZPNlScCWs
Plxbu5ze/ANvkppDmNBc+iK9vMnop8aFaPrm+DZjb28/n3pyLjqIfgS05KmTiK0zCIp/SUrbt6Bq
0dqM1xANtIfZaV2k3amVI3YrTBIf1hWZsAUMZe/NEIoJqObj1908BC8Z1/BNat7qz59w4dygW7hF
3rFDh8rHVmgi7TqDmIqIwPCD62nswDtojNjDJK8ezPw75iDrjXFkrWLb9NgmoR2dYFAnbKsk8XwN
yQ1cCTxCqSfa2gM9vtrpr6j7DovSz2Z68po/LpyJcHGuNU1USzpAyZbL4AuzmJ53uA4Hd80KJktw
mfPJbSukOuV0gjPTFvo1NMcH1RvfwH8fDRyCYiV9O/qpgvDWZVePkmsZMBRrt/JxGk1R4J2skOYv
2LvTRJUTZvT3fAS7RJnMAe1NmhQYa/mwYNG5Ijo09ZDfR+s8N1iuBl5I0qg2ILg4OTnPI5BZ8+mX
09FT1ZtoXic8ZA41DEN4m2yow8Q9eOEjvLSm0ApDAqTr/4kEklcCLdFALVYmFKEf5iz+V4ExaqET
xZCguz/D6IjxE+itRYH4SP9/iZHoPzb0hnV5PCjJQ+vtkdYES8qc5wQeaGhg6vwcpifKqa7Clnyx
PS62Y3WVQDghZnVM0WAID4LEDl4QNz27vBJtxov+qNB6kcr5SAbKggSE2DCxkFSx2C3Xmr7qWFbf
xzSgELtOgQV2wGj393GIN1ax24lOODbx7/4PSrtBqY/lULKUacc2fmTtHQsIePWhu7CfQkrQCjVJ
qacw31qJtDVBSrH65w9GugAAzxCbcW89yVCAZpCdYSTglOYev5DoEn2Y7QJlaHQi9fJJOIHrAA6p
L7Svw7pQMDI6tCqNGH6/tJYBAaDBuLHDuz0oI4qNi3LXcnbYu+IcKY6BSntkSBqSb51Xl31LylQa
fGARgU4RMa53DoCkmLShZ83gdCxSI2Q78ULqQeEPRRJx7c0rbdRTrXqVUQdStTW1BF5Ve82VpMBR
haGaRAHGtLZAPdzpGZQtP0nz1b86vI/lumFKEwhjic0MqYAN8e1CZWU/CCPEBvBDbsohJznlZc/J
1nM05tkLyrvLTn+20C6UX+qiJktArbCfZAU++zwB83zI4H6y8zrNgvAMmrIMCLwh6iU0cahtrNua
qpoae56zR/HOWHzDCNDXJNSW515JBpBrT590C1xoUHwfG0CjvnSy7YKzbvrIepaBoO6ePvHAksrR
gQT2sRYk/c64Ix7zKR8WqIhHb72oGaF6i+ncIBXolJO4zcBHxCBmHoCMGmmSG7ez0oqwB73ecgk8
NAxsGzFnwi/mKiyR3KlfPAg8QVb8ozU8jivgB7OBA43UUk0v5uH0qy77IXiBVbqRQbOHG4JB9crU
doSwBbzEf/sJA7hvaJcoaiiyr4Hp3o7rAEcbHezI1Zygv95+JySyJAPhKazbCc7AiBEmX3Zi+jYh
A7Hw0979JrcCGlWIGGPc8Jd1jLu9FPJPzysMfaSUMVBa7Nh2Bo/U4ZV81qynyWj7VWsnajfYXN28
2o4UJMziI1Wb4Y9T/6LgGEbSnr9NjHMf4ukjT13WDx88dWezcp2DcNPRwRX29vtmN6BsD0UnKK1a
VGRsrY+AE1yBadQITVB7w4F40t9yBbU6qHjzLAfzGmY2Nf+m9o32r9s1Ba5Jja2tUnH0EO6K4cEj
EtjfFZEQfcBISVZY4d6+C7q2patVfT8VEq/yyYUcu2Sgx1aekoq30ieRGvRtvktSq7OckNVVXMVm
bMFdTtkIOC4NadEQYm+PzAhZCVxXL+ppnOrxpGFuQsT5d3ntAbXzMbNQY6ncyj9NDxMo9Xxe/Dwz
FXqtNDL4OWtJ5XHYBzilv9p4bsJMTYQqrfzb02ELGd/96HBEkmLdh7Gr6PBXXKHjR6xEqXfOgv74
AnZuQsV7YC8Vhgu2Qht3xlPdQRa7JhBqOwkNBgmyo7jEiT89go8gAKu6CtamUyEEysCh9JS2wcaQ
OuuKJzJTyPpCbhpdw1kDHo3fV/e8vFUCQmDhYol8aPsUGBQ8517hUHi/9a+D+zzZVRLhSyUma54D
Vev1FAMZvC/rMULG+v127mwvvuPwsvhxolkXFQHcsBCutB8peufzEpwS/cjmvR06nYZzWgk7fG+L
/hwmeZXZMPbxbKcxafq0lBTrgQuO4smM0UMtCxn9CvkFB6rMcYKHDOwAAzM8ap782bjOOJ9B43LG
8gkQv9WExqAoN2XHGtEKdwiG7VcPBc00908cBOFbEM9kro+fFMSl2IUMRV9Syxe0Ir/9PuFswU2w
aoWPhbQgc6LiKwztyJRizddp10g0IWd2q3o2CTPd/PpDxiAHI2Yub7pC0Y93VQ0Cd8F3zWOsLD4y
HP4XS0X7T7Ri1Ur93WUl/8i2ows1gXUXf2NH0MX+PO/A7sQomUil/yhg8qdXg0Jn5MGT+0oc+Wmf
y6kcl4rFAs4rXdsioLkR5gjMR80MNFuI8ZFVjNwl9CIKDgYQWP4YkHEaiJ+/LIeCy9STXFRwDWdz
BUwCOCYm4xYX5azMvm/PEBfarmsFmOz3gdIt/r1v38ocB7WcCwPb/lQElPbkDwxbDDhUYAGJAKtb
s4WLoiSjxFUh6gk7TRkIr+suoOEzkWf/8V038SqhujZRRcVb7xL8akap3t+tCDe9KFJWNaSvRGlt
QTW2qDpO7x8JgZDvlO503gO8ndhRSNhRCMJwgcdAAHaQVyJGFwzbImvSLALzXEyx2yRYjIFnpy4R
k8mzC0wtZzPw0ImZhIx/PzjfHXssKSmyMp4OFzp+GpXN9xAAk2VmfnGkmCDKCK6541/NeYKEYaft
gEI/mjx8uD2t8yIfReH4stEeLKcAkq2+t/cbfvq5Idv7qqQ3NOTSeHvX5ncBiQ0DzUJWWtP+NSAb
4eekw5zknzKXaVy5F7AbZQ2+NfXsN5xhXRZzkSlY13naAh+IbQ7zN6yctEJJYMU8QM6JBycL266A
oJ8nsM5+gr6dzq+HvNH9QFU9OTmYaBpJCyaFucXTC/5dQGiJTaIknvwmZn4yHuUbVxnAh7zqCG1o
T/JkG5nn0dX2dpB2UgMfkzPTXgKYlLsjwzKR8hTADLGQ93NMozSl2020trQai0/gP7DxYpCIks7a
4rqSi1nLJn6N6tFKXxJ3hhHOLHWoQvcqxjQlmxvNCBx1bdaMzp0sKAY+qkn1phY/fgmS74cA+smG
Pd0VmP+0gUlnA/OIZ6pPL3b+ECdT+HcH/QPtlzux7dHX79HAfLCBD/7Jygo16HyubL9ZNLeSwaqd
igOclENpyW7jhFRmCfvGF0AMxCLfemttn11oPNmUkkjCZZ2RaGs9wqq1FvwrO8A7+rS2p26ifU2a
JkdAMHyT4KkQY0a3kk1tC2/nSXHrXN53XbcJnW9eji/jJzZjlZzF0xUyVrjj/WHwsHVJJJlHc3H6
1OwAaYcWhVvBuyVHF9IyD0pmG3GR3Q9nppOW8V1r+PMkTYfoKcILetykZKStAnFCPrg5tPhsWPo2
6YcVa+TPeDLr3YgXjm7zihkPNwr4ghj0DJLZI7V+ASplm78zBkGhabdA3pUbLQatHYztLLUmS701
zH/Lr3rSCGis0D3DkuiWbZABWS6u6ADZ8vNkw7E8SAdJnhBN+GdoY4ezFBsgE+Qh6ZA/8sP9XGAM
SdF7rBn7p9V387eYrOLvpS4B5ylQ38HHk3re4fcjq2+qhnUzOpUBTmoMh69gXkZW20rf6MyIPxi+
gMB7r8dWl2B7ah7MWfwjQ5NiSgKonuBXuqF5mFG7UD96U29m5LRNLhjtpP+gMLcAyduVlsurgA7u
y+laI599h7t3yPuVxjzLcFvf7YBz54rSV3846Ljfet7uU+gbR9k1nSnrrAWXkVWiz/8kW7E2r+5d
171wHbB6WqHXdZgndm43qx83o0uEhJBBU+WWzbcU9QTSwVKaIe39aZmkzpFd3KDoN4qU/64M/DkC
Lhf5xmI1sgG4bo4SPQADwfBqBTtUciFCr7BHSKd8UuRly2wxOCBFpeLQCL4WpyV1DGgBdNts/XI7
onAlPZ+sWsWnLB/4MzIaU8WS5/hoW+x13fPBHzeKocHPa606opmy8BtFXIyil6jpciaUTfaPpWF0
hVNtazNyIoV82cGHD8qsy6YK2g1b54h5yeLVXczfg6s2lJth0pKBQzkAJyw051rRtA5Ylh9M7Zol
0NgrFX6M3hY2si00S2825X/SIVs5p0zhX+lrhD8v+GlBQcG3MFAAMWRHw7emGnM9IX0ukU3ggZEz
wdxEv2cOAOtXJw5Q13CT10/cJ5Oo2PpVvaveUSBBaP2T+mq8mNppX/RuaoJG6GSYOBw5jpKlkYJ9
9uv3ytGO/CODNZxxn9euWYF8tsLowJbr1r8thL07S2p751Kj0N2ghUa/qfMzVvkeayb8JzhgtlpW
KzJVnVrj/l3y9//xtqteDfJoKD9/GbfopOqc8iMk1C+/ZvlI2GEbyvQE+zLRi2zlf7xA09qeS8xL
fk8/sF7CdSeZosBoRts++inclgdIEDqO4WiTeH4LQRSKrETcpPIPUrdtjR4znRzuRxAlgdQLKPHm
wGIADhq+vJB/s5Tr6AOfc++unfjmVzTLK03NVQmkOcukqJYob8PuAlYdECK/1AmOGKQn+eRZ49eu
+Pyh+dCESCax2XbkpY+pB73UI6QySpHRNp1mfWJu+crJ3UaQfzjQvwjRyCHrPSWGVibBcAcsKfa+
dujjv1lIOTvXo/p6+7oxdi2CipKQWStz7aA/wsB1PmCjP3//zL4A3XRfq3Qvhs05Bq2S4LxfUqVi
e9G+dczTfZFklXqJmrZDkVlHESVPGdytR1RhD3cOubQShcsdsyqEeeq6V1VyB9ywVzELgWsrj+uY
k95F3Pioy0b/OHFDFQvQDf28C1AEsZsS8iooL61qntABxoIIiY6C2E99734Clu3BK1Fn6ec2kdRY
42D8p3Wg3mf8zBfB54dX400p4hThE8kv7Uioh0ozXNm2CX6+6QgcoXrOhDqT7RJAXMDVtGzuM8vh
8spD9Eu0eeXP9TS4oYr5WsFy5gBJ8L5TjPBZbzHBajnRy4e5dig2WyuBzXkbs3BcquJpFs8JLIM8
OLKTwTG9+EPVIzxn75ZFlpL+un0JOiufzdwd07FdXIrdqA6HItez8xDK4gT6Pj3sAOsIn3X4di+q
t9OC0tZjIuenzb4WZorAdjt7ni7kdxmBtGlIIGLCM7ftD1KZ/RGolcqKpo1XIy+11v1U+D/OcguW
Ain94ZoCetKv1ovpANJr5JFRwZNgTBe6BDyNuZ4S0Eep1WOtKosIJJoPSBC4pzH8BPXiujJBCaa2
p67qoI1k90wXfPletJQWullH5aasmdtcnkSyU/RsPfvE3j2HbEp2CewdtUOAuOSI0m0cm4pfF8/v
dBXHvwlnbh4WGrsSCBOCQS7hO/fDxuIhgYbpwsMCQbbdlnpqJmg5kNV4667SNDQyRJzTj6V8LkW+
Ik64dpmgLnJXCcueYPbmkwZv7IFEW09fwvsjsPv9uEJePckF43baGZ6hza6gQgaN4/7O6eDRbBVw
kXJy94z+wIdKtRsyvSOPJSHKYyzIgJscD13IcFIcjr4wAOyQHAZ9qZxJzP15nSs32Cu9qT5MIssU
A1EE6vRniXVYejM/fitGql3hCB16FsEntYb/kRTNTtzBsl/bu0s9MUD6t106yne3XArM3jeSwls4
0yR7Bm+ENH+K//WjNs7elqZAzgDBDMuHo+sdsOtxsQkZGnserRKV95GEyDu8WGsWuyiXt0h6mPSO
183nSERgt3pW2/mvyu2f250eMdcs8ZoMBUsxrHb4lzm9CEYI1m1DO7SkGz9OMQeI+mGvwwbB6r21
ocBvuzYiOasOtzmFQxc5pEzlbnPgNdhC/WyGUYJJXZ3VDKaP2s1zwmxSoQxcS0fX5Vhrl81quUo5
re6vk3xdi04UhmAy8FCbm3XWvOlECHwi/oTMCJlyqvXFzObu1eo37Y/w2dW+cWZA54iDGACE34v0
qPexie+X4piS4SjMF6uj8u5PzQVHqLbrbIhAUstB1jCUjpybF4xK4/TAIjg9EVPi6cwV3UZo6rr2
cji6r/qL5j1aaRRESX/YoyLRBl4AB8YKsJanFHGacz45H4VHBQcUp/rDl9u0BqjZD3laHzXgL+6n
rKQMINt0QLtnUYTApgTXbJ892NTV+QZvLQB8HotrYiVsj6na9LRUO3/yTt/krfoJXSJTbTsSUVhF
NWRVdTBh9F6dEoOL8nvTui2CCkw6B9BbFk+OJRlF0JoiEziDAzlxg+xiqoSlgxOBrfbA6UPv9+oE
V3qClkr3UZkQy9FcLXrM3yoJEm+YD9EaIX0ZRmnNC600KLWXvmnmf4JfqlkrP12g9rSVqiBlCNzS
OV2F+UFv15jDoPz58B3Mov3z07TH0Gbq4kF3iVmaFEJ1Y5WUtIhVk/iN0wkE2lOL0WLRq0M3cKvw
b+ZKjD+duLfvfE4TMvnuGJVqSqbT6BISD1ujdt2SDwaeaqATF0LES4Ml5vSj15RiboKVbgLfkJep
ym+4KQw2qTHRgZesFWcBwJ7RA0Cer6KtZ1j+kq6ZZzYrkOf3Tu0aI3HgCHNPC/CRaIVMvLVJb1SU
EdR7lJPtAKyMtLysjTRhz+bZ6IrRPfEzeTVSzUPYTxXdkbOsIgwtObuXVZU+xHzFFO7u1exoF0+G
rLFlQYFAfWgxkMFjfGUriWbvGqao83MW9quB0JQDn7xAxRtYexUbmFfToWOhzTuJoON6M3319Nwh
Ta6mguYEPJVGlI25lTgA87HOlU6KUsL6XasM0UgqPLqnvFNPyOD4P7184/+sgG9ZFKola9mwz5IO
xnTOputhV2+GBCiW89fu9T4ujggBxRJufY3yTkMuH1U+iAjmTNHj1UieOfeDnneeVXzbxZn6eLQQ
SPpJWyl54qXuIJ4dJxB8QolfDgg5CIqydcQKqL/sAb8UrvYblj1TUXGSfW5/LgMkXlIsVPie8d4g
Eld4ET1CN6NdmbHj2Z1DPRy3c5SxhvGpGBLtf9gfdlJH26bkJ2KnJ4sCZqf7HyBf2X518od9QrfO
9wTP7jkc8KyogdECiNrw5fRakk5RrSEpiJOr/gKn3K4/fLm5cav4B9BBwlDULV2QG6S7o/ewRtzm
Co2smGXkx6v3ZXs4MgdyI4FjTlx3NzYU311R22VqGoYfsl9EIAML/cfsWdsyyrssbedxiAhyPGE3
MeK1WyT9LbmEuExBZhPCjLLpAQtEbC2ucu7xuQ5NQl5U+TiXyiQKuvxtoQDUZaINfDbzv1OPv9Lj
eaff+neR9x+hmw69GxsHJaRePoMIaI/xxPyjlziQfWHQGbv1uj2ezYhcF77g7V6RuaVGAHmaGRTG
IHp6+1bmDTBKIbD+3XLvJ7dBhNJnr4aQl/QrYTuoRxEJ+OeRNTJmdpioo8pfJjU421eA0WT+yBjJ
+ChUZDTI1GhINWKBPYEaoT4An5B4PA7d44MeAgm8YzxC9QPDYNngi8SovDdyxfbef0ZJ2km0rg/h
qIAY3qhljr1PWSzT1UOl2/L0/LvwiBKtMJCjrjn/3ZsL3XfvwTuICq+78wRL8/Ob+MmFAwk+sCtD
GIVe9SFDEyWQYlkGXAniOqcbvUnJE2XLNRrlMMo+hVjZ/pb9GRoNLYIY0EUPRiywSO7zL9s40D63
Yn0hkq5LQKCyKNqFYsz5SoAPsNyFW66Pc6yGC/d1FSISjDSj4hgghVvCbNTBhSMSlnxyrU4B3m6Y
Py+03KGfZ7CDkrV9BZfJiSn859RqAT+JO0ABNGtZkO7CspHEGz9XkoPZUrr9i4ZCl4hDmDhbo5fC
p+97BwkRa3PBoYPIGEaOOugrAXawacpR30J7AGRba+LeYB+RhowzMfiP/m4ROfcF8nfA5EXxKMQ4
GnRyH2SGcBUf9j9g4tQlg2xDLzdCTmbWDvnlAzQzdia1PeCWN8FuH6R5HGruzSmWGIOZm55QJkIn
3OhX/feosepNFX4I7rCDe2CvVwxWSU2awftVvieDN5SwwjUfpV+XtrbVmeNljpbq0h6KjqVdAL4R
Y3cof/wbdSPIWfhEh9lkmm/ugJQ6e90zeYMHYdwAxUKr2KKK5x/jAil44PWeR9Bzc8dcAK0GnpD0
2vaeje/lPw0fhRfyTPhwmkpQC92u0kxkcg+IsVRkSsnr2lNTUHS9kYD7kJ85TDaiwhKwjX2mmp0B
BHCCjnVd5dHwhDPIgM7oqRAH+rGQjhAYkChWl30OBLYK6nmzivLw+/rb4vmTSKgSPKvganzm2qTg
SMgIj9bxXhT/CZakUGOXxoThApXjvBHHFRtYreeq+G/9XZnNHYP2sqEJkCkcHJTXa1TXBI+Rdhmn
pDV7qWJwFLGqr/ZspequOn52Lr1XjGkVoxPo/XICNmkagqcay4k2NEcTLAF6BZUdAt6gGSQyqS0j
0xU7QqWBvNg8D9105YFtqqOj6Vfxc6bBH8EEqYPlMeaAqQaQfLfbPjN1CJcxcgLP+BeEc0Yhb/WV
NlUg4EbzrXLMC5AdZ2IZIbBQ9x9tELIxkBEx8rLZIJRoDsfFwh1+WJTci921yOanhFJv41OldFSh
Ggcj0x8z2j3PN8jecxSll3559Vhk8u/SzKg0XocJVCOCxHXKc5EaB8S3I5wAYk7t69MQY6iuV48L
UGJNWelYqJTYkkHDJm5rcu3nD+mUuJWdtf7AXsBt7WTfmBR0imWDz8kCSdT08lY2rBeaHSz8PyHY
iFoqwPRJ6eDl40y7t08qLLKUUj3Hx15HiYz5p6rbL4VFmgNrTFZkF6ZBJpMfRIiBGikBpYfjmCuy
d9xgzLKboZoJDyrgKb7jPsG+JF6bFIz3r20XwCAxG7M0DLuvOhszK/oaWjjA0uhlgoBkbTugoajM
tAqcQLKNqO2L2uNwAr6yLBiBHZuq3iTPs09QkLBVytYxlpUwXU5EEsWiG/eY7BpvjJocgXDdDDzg
dL3AUDlzwEEmKrZcCfahSt92yy5ERiwStp12Yz5BvdqpWv+ErEog87+IfI9Ok/I6MjmHpw5Kfchr
bIXIP5IVdTk6F8k12tJ0Psy0WqYx2q9BosvfWLZwKKmMZbgC/fYiws89HtRZ7nvW3sYAqHO4pebR
8vGMx/+vAUMfb34z7vYNEnXwPLRJhn11K79SPMRN0ic+24fvl5U1217iYwE/hVCDPIQb8Myhor/E
Tu2vAc84ECfC2FkOpilgVQlhrTIuyeXNQtk35FMQTOPLORQBa2vRnDmXw0H58Oj7jvasTx7CcDKs
M/pZu7C6c0DuCmmdzLcV8BLu6FwojwlfUTDZ8L0fAGCpWX2v/zyigR26+F7aDNRIcRkjAaqiPSoR
EUJv23Z0SwYNstFCF6iFmlIMHPn5yJ2xaZCVQ8LeiiZ8CIIu2JeUz7PNiL+LLwqnvpTkpaBlLw/e
L2s+oVsUe4s9ZeehQTIo/29LWnTQ+VSaANZpgouVPVB2d0ZOaBotR2L6PV4wCNEWvTa7LFwCWvXA
wPUL70+GKkzJp6Dq8n1bTj9JWrRvVveg49dZJdMt3ncVPDgsWbRfnAgTybpHnP1uWXB8M1BNPN4I
Kxc6bhAxHjLLAd2nE0Q0/IARmE9pcSJvF3++e6CyQqHnAPBYV+UkEDomWMt9LSpr7/3ZZUkiaXTt
4KX4Vl+WKO/AegUiWRYjkaBDF6aUgFzKMmDyQJ3iCq6LEo7PJALV2z5le0aYXAoLerxv5zzq2NOG
DaH4gN/Ei/N8F/EYOn8PS34hxp7GGyExykXmneaEHN+JuLPtBkex2rBkr0n2thyq4ash15Ebr4f9
8JyflyqgbUxT+yDbjBMFgVQesr5ZHwibYr6PIgwRQM9fdG7o2fXBEFI0bsxF54ScsvpCve1lxcBD
2bDc90BrpdWB7jNI/GoUWYKAHSSnw6hUktfUJ35AE2F1Zt85oBqN9ycOex9WEk+QWBluSc26S+aR
0XLrwFMhQ7XwadNHtgFa/Os3HkUjliWUzsQOB4eegF9lrcIqMoqxXV+kPd5DJHOcXa6szOgFI0d6
NFdxnGfR6L2eP+1eLO9Ti2rwW3C/xteBqu+4/SqoKMcm5rHYEwQ0sRs6XpJt1xRcnvghzJ+n519n
0bfbQ/WDC9MNMKxxNu95X9KGeOsAL5cZ952MG3pAc3wZYSR+BLwbsc/S2qxA6LPp3yNG3uZ9DTLy
j91Z/QGXShLxjhnkd8GNFnN2c1WndXmSNvUWFclJxXTSWsXGA6t9kdUcqv2upGZ9Whlic/WhRPwk
DU6or/Ma8M78tLzFWJEq9YHl4A7nBT8K0H/9+WB1guX7V6uAg8azEcb/3mep+t9khPitUxUMOhBD
nUiPj9+8xs8TQZQp3FuCqAOTME/jZiJ8nCUlqQqIZgWRVVjGkpvqfdOt6m3LGAsn7E9TD863ZJ1c
PspWd1hcUReDGeWFGPYqu2ubuWGZid02m0OI+9KuC9CR1jz/UU1sgb8zxwsj7O0ypInkg9qCaHIm
vBIvbZ4AhTxBbf+6Yt7H+q9pyFQhCmm5ANDD57iqHe2ZoVdA4a2ya++Xg/ecRNpAR4YEwMt91i0n
3baipLOulnNLzs0GPoz4qgOtWsqFy5JUdjMhmn/zr2c4Eo3DS24cP1oTcW/KZUQ796/HQlChuor+
qkdbVvVnifjmmH2sdQXdU5oGyreHYi+VbKv0nZnRcVbOdlKK8Z8O5bGv5XF47hrPGDp3lbJAuw/C
E+DN9AtY9rE3N9KsXYM+4a5PlOio+JhnOTuWWDMVvxUT5mCL/xnlztVQS+QGMfNIYPCEw3hAEQkL
+AF5mnnhUeJ7gEUxDUVI196MtNRA5fQIgA5vSN3I1rnlfuJ1F+jr2PsnUTBoHovbgM40858zN3UX
bOD3Uz9uAsfC2Gc=
`protect end_protected

