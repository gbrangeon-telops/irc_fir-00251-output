

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g2RN5TBir43ECxFrT/y2GRXX5NGDYpjq+n5gxNTYWsuzDCjF5YeYUisYseKLr1ryeyQynd8Epzt1
V06LipLPYg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eJKP4nowQhkS+sdlDJ3aF081jbTFWdzdlOBNNOlq8qkrol2Z2K32WIgnl06Lqx6yc1xJY0X0kmV8
eOkRE5vog2ePPioAy86OAcMONOPoHTqykW2qaaCPwvHqEP73jf7t4R18PaTf0PZeg4kzgW5BQXqF
THWJ0viu+pagUeVYQuI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MDIZ/fTOzwhXm05ObJ3zkVB2FpJAN9o34cB0jHfFprFQZmUeUQ3tZW60svZwBPLmTXGm6NjoSEnE
d1b16jr2OvP7e61sGc1GOIzSD5lAxq6KYGFDCFGlb2HKuXZP87xm86ePu57tT4ld2oGvDNavbknR
LLxhx9ZyBV7SuzGo3PKuxBA2tnF6vIEJkp4n2dqwXnKJw+xgySn5xCMvJuNm4ghYOfBAsNQGJ39j
9OlCVz84SN0I+ZhsnI7KhLpJBWOyFN5hfdsD0RVsTRLOBu1rLKX6200sXAdAwmaB9xg+3o0vilh4
pIPe6hkIVYlfHVKU7Znj0kURPqGkJtm2RI+CaA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RvD4A+WtjqxHYEUrji4gUWEBsLfMuiFWzgBi0pzOF5kWQsF7tHiiAC+dbiIZv5TBKh6/SeRqqj5f
up1ybf94wq9EXJ/d1afld/HRqNac4VRPTUzPBHt4z5dEncFPVDK4ucOaLAd/3B1aieNd9xn+mBS/
wR5gmSxp/s9f+zaVsS0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NS2iEv8S/DLjr8oIhLcaUy30De4W+2t5q2cf287k87h3kSCMEoBnjvcyRcG6CE1IFz2i6ewnJ0mb
4oesPU8Xde+4KmwGSKnw2OpNx1aFtJHy7C5xPLKHuYCmY+9zM9y9RMguGvxUNsPvXEO9G/4BQZtJ
xHf97YW4qiiYtbOsAO8R0m9UHVOYT94pj/6x0Itkq5yeU0YXuubMwNfZ5ZRnrVKNyxQ5Ilm1kGqH
N2bcD8eyFlVJydABBBV388JKwKrfOh5ZHUd8//7U9+6XMFYO4OGZzTYmAvyyO7iRRKEjPElnyW25
UoL5ziiALbB2biJ+eBPz4dgChqDQ9nB8HsYg8A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16672)
`protect data_block
sHFYuHfhqhvQtsgycoymLGPAotICCcoN15iciZSzbqSPCQupCsKokoIf4svmhxl0MllCO5GPDHN6
GlN0XVyv0oFsyyBfuw+RxkpirHzUg1vImGvhGfBJk2UuSObxItLn2WPYwYY/HDz7JqU2Zt8tKnAL
bF4FD4V6IyaryVTht8gRrICv8K1xoEZ8ycE3M+AvtgZnvW97wxHCSvx6Lhv2ZmB0UWelVzVIqkno
K62Y8c3PU2Z7WVPnyexgeV9Qc8ub0vshRdK1g/6Q89dSvKrUOCi6QtsvVyIzyQK1F+bUP0YV8HXz
h5JFOLZqouM6yZpb0nBbREPF/k3giGVnAlz/r2Fs2oOCF/16xqotQhZVeJXhEfQ5Tkx+f454DMe2
YOictlX2536iP5KeUah5JetetQMJG2YniTlYZbFbG//XQG6D98hbuNQsW7rbaymxFjvWFhmzjreM
u/S9o1IZyMhFc0nM7KlIHhlI6mk4KsGp/BPmKS1R8Xp49H+y7VBT+EiA/2tN+bURRYHOHTI0rZF0
HDpI0T0XcpvO695tcoXmZRZ3fxt65kIWpTOB2BMwropTD8cVq4dmMWA2BTqt+c1Oi3FcdBak7o2j
3ZmPQlKhO6/+iXraryduPAfSRz4mvC2ljRmOrlEaAinPGRBnLtM8o2f8eFZCb/x4ZJg0qSfL6CLo
G3TiLf1dKC7PAv9g6FgA6K8igFh+yTX+hbUYtW2othGqt1tQC1Z4jT9Tnf4gXtDQILLd/Z2/O+wz
EXQOkJaloNb0+byANmT63o9Yw9VHcX6Nm81cnuqrEdRmI00QatOW+3xyktegt2+y6FGCBjHY2uTq
hvo5hZ6qZCbjdNhlAwX2Clal0wolzf0UaG9n0S32LIGI8D5EmjqjAZS/jV/mWl65H5zP/yzeU4kV
SfPcSUEX52XOBsvX7rP33s+xk83KdAIl9z3kTXC9yU8Fj0oVBaBTEY02gelLekqKROzONRy+szl5
YycdkBR+m2htVJQwTLTnOAb2zaN2N2OiRHU70BgN0PDtRTbd4yYI50p7OkR/CRAxYs1y0WxdTguP
A55oK7omcW3Mec2h9E2G/WVO8swFru31AUOxITvSQpQY/kx+Nc65YU76RVHEtXhMRaxbLyRA42aY
mfD0vmTFdmZZqRckU6NK5T1upJTTuIS5A6ronNI9mL3hF+bljXS3McZZSY91zKQEylndbuJPMRED
AosBQ+J7xzxbIWPk9O7SRhWZ7ywZQPIRKwbPsMC9w+mR/uV6LycfABza0ultVCCCm2QFDOFwuSHp
Bk+7sDk42//jQvfmzcD5ejgAn6NOK92/52PFjv4hK1GHkdPIrJoaXe3q8vebYyWhvF6Q1DFMwHqX
UBE8QarjolS/n6eVaQ6jQ9UAYU0Xf8zHtKkgLprqfOSWm040BM7/cqhDtbW4U6h9DULnzHXFB7S0
4s6XhN4YlW4b0RVvVyEKO0X8nLzjDfb8ZBQI+Cdi408c/G8F82GOOwRvk4DqAXWiJFJh9prk4ajZ
ASDJZzPwyfOqulMW14AY/YanABt68x/xUHumqIoyi8eIaQYYIlmSSxntTyvtZM2FLEebTkXGFklJ
iIHFCNdZID0LruwsSnZzQxWyYEFLl2Ic/wS3RPGSW1IPBYY48rLzrTb6PNxh/xTX0H0JwcpWXBVZ
Ow8GATwG9pq9rwp/Du1aZ/E63iisJIXWdpC4u45JvRKLDa9a4c+DohSOeEbb9kjI8rdGzij+qhHv
2lqcv/l5Ac2WxVcD5WDyddeRz/CtrA+GMKtTcEuW3sJ0pEivhQDlZTIx48tgjyDVZk0ZWBz940Ar
YuICO+cgOoL2ZD+mstu6ksemZ9mwPWuna40sUDfKlkDhmiJ8qLGVxUYXH72dq4qHraUbCdr8daGH
sXqNcmgSYONCTpX/mYiMsRKsSeO41jBNKddC7Pn66B2kujfUSXARasmgv/uZ/P/Rhfrax9UlbiCy
sUZ8c5i6WlaL2DFH6a09ipdErZI4Y64vN9TAF5YUsiW4fE7b/jvjGm8hxSTMnhqVCvbWKRxZ89ST
heYlod6KZsrJSqT/Nm93rW4iLWuayuiwVkFT9t5Zpkh7paStUsUIUi6ZEobdUGazE7KnaKOGsSBB
2buTLmSVl6Mht/Gz4IZnI0b2EHgagL5j2k2FlAFHaseH+++VfCvxjuZrvvVCWexWBAWR52lvYtp7
LwLzyx+E3uCfVSIzzXVa2f0hGkLXZ7LVV0SJCVv2ekuo7eYzWsRNV0iFiMJeIInEOMCtNqg6u9U7
UVGFD6hFn+IBg86zK8+xW38PspSOtM5cmeaS+ZLpAigR5tCO4GDganXDcbN1nETfJ7Mxgxd0SjCV
qNu8w9i96ghoi85C2v7OWdVOHt5NR1OGpwIwCOpAqyDQ1HdBYIV8+mlcShNQ80Nr1Y1/+MATWIU9
b1zDo2KGHQX4gGnTHT3QNe3b9QFV54qrDlD2pBPn9Zua0mtErhnxKizhwqet0xs7JdxSgmafnnUN
TxBTzkk/hsCC3nZpiMKjCmEPdprorOlAZZkdkB9YeiYk6R/9LJ/jBLjjUizmheq+u3dhxseh8NZW
rVnPtFnZusLulgGfh6W9+yYg7nMLswf3wsFzlaF0wEaXX1hgTC2CMJw1ZGIxgMl5E3a7VXZ5yiY9
bcgpZa+RFCeVBwEAVHtn3xw5qGAreiKr4zKQUCRW9sNUDEniJMYbRojDc4vRwTwyvRgQx2UwBkWU
TeEgKWjQc34Sgdh5aK7JcavnFzx8tbyOGco0RgyjrOq9+BQFnwxcOoCFaETntWAskho0AiPMnn1m
/Eyl4NKJdFWtfXel4r3Yo9PGCps/8x0tBn+7EBkTkMulURH5SrNdWaz6/LY3foesp8VHnQDNKJ4m
uJh73pgadgHUAoxxURCSdYTwwjgGVbFXu6RUjM3l7w+5B6gdaSGHPALsnfJWNXk0e8v0BMYHT0s7
1rayLbJOkhw0tMKentxuUA5JmUVP6Pw0WdqlqVg0TiwBOC8cwmuXfozFyeIcJbOGU9hayhbECiUj
5X/6a8XYGs5a7VgsyMhqL5YyV/yZq5IvqCuhdfUn/LzV7fxxBS2ng00V2ZwbL/XxLQrqC/ROMdHL
peXVEU/lQxeQ+ZAvANn28UMNIsxksVsSCpFBPjSSMB1fvkfTWAzhA3tl+VKvd1oZGIhTZBOoj3lS
OLNvR1BhIfBrrtKf1wM96sQhWPWPKp8mHOcCzkpW2eE/co6itsr4bRvD24RG9kCqGZRDn5ShN6gS
ukJOGPiAxflkko7za7L3qGshvRkk29TJ2q/xPnpOK3S+DnbDVPS8GgdzSE+m6QdWNQsrf9Ub1Oqt
IVK6W/ycwmsW7S7nNJCYzG1SHDwYBskT8hgR8yQsq3bEcLYvJLY7Uij+wQIiPQDezL+gx4Nl5d2w
ikG7DXlmxbX/qbu59nIZyeiErLCS05bWxtQRkSPOmJeJ8ji6NPg/iS5YyBfIz5d8Hy4sOF2PFC1H
rRdWTNRtYJOtmmt24g5lobRDHOO7cNCK50hQBFqvBeOW0f0GRVy1Ny9ivgQkRpkGwkopnBBE8FIG
vlh6KnxNtIzaQdDicWZFaCQLdzqGu6FSGq8IXKWpgnd8WYTKkMRyivbWUh6UQolFw00jvlw4xU8c
e3SacT9yi2QzK/mbL3jv8aBMeh8fVERdMkLFVcBdB6kPDScGCUF+uCfgXQQ3Ou0RJiVDsQ78Oe1T
22+YXgaYycL9wxFHMNMtx5w5J35R1CoqZtPyFkonw6JHtcK3/NhPPwrZUqcvNiC+lR2EjHAGsx/4
qXBDbuqhVmPKwrmNVGTD4zw/rEmh1y+sTDYQz+sgnpxPaDLF40VMMgV6mNz76kftVRSRnSrwkWIj
7w8U9mEhWJEo4LtZPV6x90wnkm89pCB+OeujtVg2TbMBl+WIc2WhnHUkIfxBdsOl1WX3PlbEHFfg
mfoWgp5TCM6pjWf0piRUiJ8u8xoVWaIKPJKj+uw1rBmLTctm1/duk7/s/j5fUg9Z1hPQDWyjEvS4
qQjDzBRQHfMdqETYSPMB4gpvbkOQq/abdhtho6IvIk3OxF69kkHPaHtZTPoDphNGN4aQ8bhawAV8
1C8NEXXvCIQjZpfWxzPvqt3sWi9ImZJqEJnmfzZmHqQ7BKvpQ8tFOq+0us6+gtNj/W7/n93HefPs
Tx1FnRlE1RB+E4AC79CL2xRTwfvkWMq5KPRBWO7OZf0tp6RAchheosE4X0ReGTYqRXMeEe0V+DjK
Hymk83ft7tPyC7vPGixyzVlTSYmZK/ZjAh0rBd96P8QVb++gxxd4b5oDl3LNS1k42qayH29wH5N0
QXUzDBduGKAyRR1zBybqLGSlJxS9pKDaEEEQZvLd3IDTKHXLFf2+8ikvifC1JR7D7nYpf5bTz4MY
tFQ8DyfwPQp+PniUy4C9AzKG1hTnEcCwDQS3bBM23U7FLnXpycZv2wR/2ZyED57ESy9xAQ8ZFCKr
colKk2tLMqomXMlHUrng5TMJW2YIzlEIplYi7RHk1vsJmm4QcqjU4QxJuXEflEoVOn3U6bNgNNs2
gLKn4tSQycI17y+NqiwaZt75FJDmLNzn+g8mhlu/1SrlevI8XugGsp//IZjeDUX3z2nmSjXJ5hiy
wGCmzjszRVfNu7h+uOvmOuG6QPclCgu5YZyKbmcINkAR2ymgL+XJewWGHY5PrMpI6yqHUyqtLNif
1jBIsDEEZOclxVSoRVZU05Xry4dIiIlPZ/YSXGjk31Ro6OMyubUICYZujHZH+oRojTilWwXPehaf
XnLUMxtd9fKumoPXFV9nKD0VdHo3XWDOJ78uJyh5owWusOanp8BDAoy1irKk7FE3cx7NFUlQRrxp
PCYtTvZ13GoBQwnbcyt+2pW29rbD3z94C4Rg2lCnRz3zLvn3oV5d9lSfB8F888SbQlUJXm4EIRlJ
wne8DL2AfyH2S8ogqKAtmfN/MW86MMJiG0NmCF+FqiEbQ53AZWvrr05mumF4Por9sWqt+EIfmnuO
BN/mgqLrUshh4nHIrkT/8mHfM3grspRq4IO7ZY//43aeE0ia9c6ZJU+gTFcm/7JnlLMdus0VKwH4
4PtOs8b8VtiywJo/eewajHu/mzDjwBshnMMlhWQvbc9Q+z1aBfAithqXRiXAAPekSdKpGOqkIJhH
uyc2kwHihZlYBj0PG20aB8ZrWV158fJuEcXWQNmNBHpBB44JgAlSEgU7S4xBCE0K/GlfYXP7omFy
BKLeEDx1s+khp5qDqO9TBEqa3luM04OZxqvi3iymVrs+LrRuCBrplCt2neSDQ5cOHAdlDV3A7qYq
k4EVWcg+GTdvNa/H0Nhi0SWph3+3uEpAqIjL0AlCvlMtwGTviUd2As6CE8ooyV5PRTJGvX/ppyuO
7bcpU0cHMAiYVi9hptbDQSOB7sko5ZG/Yj9kIHPMTzOrGIHT0wPfMK21NMyQLxbUmT3Yp5N+K57i
dNtiWsLLXIKg0hmP27P25Ts0/bHoQe/N0sWQN1GfzBbBs74i/Ut+UsXbPC7MX4xZM2CJca0Q2iiG
8BMc3jeYgzDZHvQO5kv60MgHOjoV5nQm9rv8i+rbPT6sR1TLIur3zbnyHbW84g9cNa0UpmT4eIQG
tHq4ImrnKEIJnZCHN/HW7JXzxQUsK9jZhdDd5ZoNMHGTQHpTDr0B/HjefMhr4CctN0d8+/NL9Uj1
FXBSQQARjBr2HyNL7DnT8tBrnNuLl6FxhxQbGXIc5bjTp26Eg0cbWoQ0ZgDrtBqovgMZi2wuQiIK
noTxLmrLeqphxTziML51zcRDUdvu/DdKtWLaeG9P078TVCBeH+9b66BbqsPAo0ddl+2po9xwm7fS
O/aFk6Kxqu1SDgRxAsU1FLN/9oIhsyJUaReOseAtocpkn3LTYh+IbFZZswzaw+1PvqYvsHSW3xt1
uxEX2vG44aI2d2ApOcS/gxHjpBHbmLp0nQS4l0MdLrbacI91RK6Br8WzS0x0Ti53dp9FjCb/zw/g
N05jPYCLmx+JqnTTN75tD4kQ9CR4C8kbZC/MvDzTBSgoFMzCOE5H8Wtb5CxssKewIKbDoTYSxqjG
BIlO5VAj3Ag1h2q/PehNX9naH223NobQDXmHYRubw76IozBzI7UDIAG9rZyMzJe9FtqF/f5O5eZx
0BR9wUkMSV9KcE2aMuymLaVKx5HMlLtgjGp29L/l52j3p2k0jYaFKGS3QIShmSiXapaeFT6fTRMN
uUCBYG33FGX+xkxgmN/8/ZOiR4ZLZzKpzetNMOJ4zAXmL+YqiMw7LKXPFVXVDAfIX1GAGs7KqsY0
ebhU4mchyW2Lu6/VJRfJqeLPrpGrBWn8iLCFANGd/A6uKuDn9ByApTtPctHM8pqTisJ4Z5OmrnNn
r2NWPhKqD8NCXYi7gjNCdjYPGqSCtY9959UmsaaWf0OAvlDtQN2sbAnpkd3U1OXBKm/L6xsvmkCq
W+gb8333sAonEArnAXZDPpuFKQsI6y3rNlXNPyqSd1Xj9PyWSgRDg1OpogHdozLvLPuZ6+SLpf7p
QfREYJzLZ8t81QQQ8aG7mSlFPVCKSLfHl6BYKZAcM192+IdcY+EjrKAdS416G7xXYziiX00NPSUd
TcwwA/6JAJuoaG3PflB5lWnKu3lTaUYf+Tskt9fX8L/b6HJjBBsXC0Qyi2EaioWt68peL/fT+gHU
/9kGGALn1NpFnBrzviMzjNsDqkj2LkcZwBs/MUsgdTryDjAfM531NBIoOpRgNTSSUGr5zoYJGN29
O4tmBHtKhdf8fliVQ57tyq/ONUgvuJVsPlj6mU1wpMIj7UbnMgSpuaAfOfHpuCGVzFn7R6rtaSxF
Uhf1ekVMJm3VIxqbX/4D8h5y4uqCIWgCTK9WwUHCi4ck+LjxLefZOp4Bin84SL0MOP/MpP2izG9a
c2dE5ChpHqzqxtQIgemPQ+FvpnI0NHTj2ofPyFURZ4bqAMLIADkGWaFIQuWVNVk7xkmnCrI/T5a6
mDcCWgbitEGXZ+HLh07zKG8GjyPDYp63EJ4FhCwc44/bVWQcpNlRaEhgcfQqKhiSiHa1e3w70STz
cUNBKeeRS2crDAIhnqywqe0vOhICpbe1ykti7EiEoR5Y4jMu1EpgA8bNh3Q+tF5sf20u3iM0byH8
cMJucYQa96Z9HOfOHwJUj6XVWitpeD2Xr227slA9bnY99FCuQ+AAGr+74wYUFBBmBgg/e6kUugfZ
y+YNvSmjXfRfAUHjMziio74hjRz8ASpxgxoIBEZvZrCBzjQzxUo/YuCfomLC4OvmCDpfZt9+xJk6
9rzY7Dt2KFwkrbIy8HIjdjgdXV2XV+j29GxFZR098hHuxGCpSSWaO4xIsSJpsw9knQImeyzhKdA9
QlsOIyXrLuJFKQg4oY3KWnttH1ArdYE242Auh997WKK9g2UAAzrkR/at1adq9hGqYhos796iNAyW
fOy//wV4hny/610zc1xxHKPqSFnbxSTpkqVqPC+9gX/o1cFxymHbUKLzmswjV2SzYXKAiQZeHgN2
ycpQ1X+XuUYgX5ymdrKIjgBeeUh4X4j3dkU1qaUsVD1nC3JcUL44KnoqxquvqiCAKFof/6o44lek
gJz7/wniNpo82b9rvKlWsJuGesuo7Go2LeD4DV5ctjgb2s1Mzub5FcFpG+v/v8EKIEQKs8SKv2B0
b5YRDQ2YREfP32nhdiSYmUxVh9FejuAn7p2enNQYZXSeoDjlWgr3pz2ZvyZjuii7IjdBtT4V696x
8g7JqemSwHX6qxpIaHOwRyJB9RuJEG3Blb20D/Gt2srSNpcyWBL09BcKhxg6V5FhBfV/Qrd3YwDe
ldCmNOHVERPYzA1HVfQhwy5Ovw7zZ7YdtzDpzmYEnTbKrrn3W3Cbhz+Ya4dN7s4uz5Qzk4aa+1X+
Sph0q+yw+ayjxUHAVJ11qwwW01rWIggMAnWPp7Z25UoFGBGwJcNLOmS3BbTjnFCYO4QTzhIiNbaE
xNNaCu/7TFJapQ7fYfuZpFkg7JKHLkn9B5RGwyLKxxNwkuJFM040RFdw9m7tWfBsYAuffVIU/Dyg
P8JzGO9xM+QkFlRMWf0VLa42HJ52WqMDjxYNQwKdBU0QG/OXJAd9FJbBxciP3yMbls5c4I9t2f4f
ewTz9bsPm2KUi1DYXD+a2Vyir3H1VLLuZfb7ZTsRW+Mv9bARnYNuiTtkDkI0YZ206zIFR9Cn10xh
oEUdoDsmzVUjNBOPVoX8VlKAM+0qgn7Yi6o/WcylhNXnqjYL/k6CrleAI7s7YFkGpGi1UxXgCPlI
ReNN67vScFnbFGgCoDG8+rYqiNmz2YpXbEvkFHfyYpLhL3bIwtQX0b+ni5K1V9vDFblMMEVsg34a
NXXjIL1tImQxJTjM235GGnpgk9OsC5PmQQV/OmgoVWu5yWNE93qmIlE2LXfDXTFbLKkOlpvGC5Fu
D47htO816wjrgHpEXJwFfQhk4jpxGCtStbTW5h4NBraJxI0c4AiueoWaFOXzdSf4xoI86D1ccHLh
eeHae0T6JdX9FsbqIfWOET6LWNg3uC29laKC3cBU5wpXl7pb/5OnMVDtivxKtMCtQYodk4CKBjLB
2pqIBxjEe5F7/p0y9/FG75kNGFnoYqm3gqZh2DKy39905TavlTzdDGoPgFF8ONJIatImrX1VvbVy
19Khl4cX//CuTkLqZeYIu3eDqrw/jIVNtsinCPnsOr2a+o0q1iW1cjtlyu4lh6n9L72uh3mfaJVF
XtdLWrTbhF3JEUsO1saorOgixTRM/XY1ORG/lNGcY8sOynii4VulVlFB+7CNKYZLnxrwNSOgcZsE
RwvfaN40PVaBT/BrMwnHxFayp9Xrp+H4IdLQBU2UY/ZZFuOhosQaNWsROcK14XZ7xaOz96ydwLxF
1PWaafHr/tR9OSDd9rp5Iy6mRpLf9SpN6+Zt/xoPvja9sgf34fp75trRAln6Nvr8VW3UdHr/LP3+
PszHb+Hh5pKBjIJgGGdWZRs/GjcjRSWt7G05FPj9Lz/SXlGw3KmhNErBgDeoyLT3LbGIHlOB7gTE
9WX8B7Dn4ZyrYdQ6AveM5rxg4/i65eTzxYlGDW8fmRsGYpFXqzUkhG87JcUsQEEOShmabuOLOaGx
NkTSl4n48M+Yg3rL6lt4/Rg5YtjD3BsZz9LhhBrqW2okiLac5Erk2F6nTiImU8pUfdGXH8/zXPaR
hNYEcOyBOcfAp7MsFu4aCWF+w9W3yBF1GP2voWfwCvuNHnPBMsPK09C2eUUSKbwAY237ImreZTQn
JnNWhR8P6Gscp17c19lDwTnls7kTH9O4C3xMh/Vmsl+VWoLAV6tpRooAFrsTN1wAGRKyLMsTrxI8
8nrSDQkZSDvhZx0QwoTuj8X3pcf3egKBDVWH8IkoXZP3d0a7GEbD6Bd6D/iuerA6qO2PLe6Tp2qe
zZYUXA/3S8Q+/TOByJAYVM1gy+W6Rh38ZdQE/pk/D6WevDO46YT2mbztLyb59qV+ZI3ZBpiTl1Id
OwKka3qNQoHU02XeITu6YUq/Y2PIKKVGonGNM7UxTFZRg/l5ifAkCRaB9zFTNTxy0gXSouA8bZuo
MnMGjXI1yVaB2/JgWipp4wp1n3hwiAbbD319mjs/SH17ORoV5LrZJNCZgK4eWpyuNYe/hDgFrY9h
soMuXZpex0lemZI8cqoUaRExvL5PEVI2Oz3Xb7a0D8lLy5cm//EmHa9NI/ZDu7TIfKZwggx+d9he
5ul4I5mvtf0hNPh8aDj4LErfMpUQXNXTzH8ax8d/qKckMi10eGwonq8puVkCwp0k4LCIWMWHq1Pz
JVMDEROruQILZ96dSx4JiTtenn+a76pravhuHRP+LTOLzLPJT+G9Oq7/eB8AWjmix3UapreHM6Gz
K7PMb+OvdIKajtTjViIf/UYvv4eA6dOApYdfQ8+HdOqjXLj9D/hhCTMwKLFOrTPHAkjfhLsgC2Z8
PPDZOKdjF3YutMnb9vu9DOKauKZy5fa6iOxmDPPqJ5QmLdQV70gYr2bfwQw8qogiGcA4aWVXYf7w
splsSLxJmGc0/sD8/Dd0TGELjGjy7VUhD1+OfdNdc5d9qfhVf8QX7kySJbCnejYGNy3fLbHR22X5
RsvAdMYYaHqJDFzm7r6zPgr/1GuAGQiHErGb/j2OA68Ddr9VmQVWI2X87zhen4A/RsnKEmqIuVE8
t5eCWwCRyICljKb+aEXL2CLoGTPvXai66wwVU0ffaVYR2+kK6mK56R7o/oFIwhlFoadmk/LeoGcO
AOzgFdgTh4VIqolYJF3HWrLrxWSjDt63gWOrgobAX1UmFhnJouddRBsjqUk8RLYFuyRfE3Y5OOIJ
9rsADNfR9Fi8gtM4FWjOD//GgfITbMczZZE0lvhSpBBnhWEhe9aWZ28mp2fMaqvY4yYzOaThkFOM
GTmn8+Ej8+7ajiuqZr0SnPhnFIettSrIn4DyBajWlhrEI0e8KL3Xysv/T8j51YLSPl8CNLF9QojK
g6XgLNKs6pbsmcnHbIeqDB7xlvDW/B/jj/GEpJu/f4HCO5xmJ9rL7mO4q7erX04PN/gHQY7xJzKO
tQph13RbR6glyDmy9nT9jGQ8C8dn1z33SpyzHgh3ka/c0PVPdH6gcfUZu11WNbpEj3YmDoeGWIxv
J5sbV3aV3+jrE0v6b8u8TJdUA58xPKzaOPmrL+tSjW3ja4rgQwtjedHouHpa7Zr5qmpNO5wGt5Yd
4zqdHNAq2CAi379iA2u/jRPvQcwqOQdvsMzriwSXRUBpb5pwtmNGgDRcFnLY6bYGE6bepyha3idD
8pLoxGro+9zQFdICqJu8NyrOe/FAz8USr7Oj+6kKzt3Tu6e3Zf9cHrRQtJZHwwX8DHc+GVOsE+B1
5R5GnzrlSBKLe6YeJkFtuBvIKQqmtdt7cEXpZ9W2AR5N+c532t5AABTiyvIwb0XMetUila11I1fd
edkkLEMrbnE7udgEIaE857Cr/yHBNIeoQIcibWi0w70DZC2LnE/qON5jFHJteEoG9x/RO25zQpRm
ZJAiGNkSxGSKUbqLliBg3f1Gpw8ohUZteA7rjIi3CvS9h0xBTYO6xfsQStC1Mx+T5llvc9TWwe0c
GGq8MeOtH1T2KrnfQKhf4ZnbJKTxRRyiKohpODbjc0VoMuSM5z8OgaTdNgA4tvR1myRNvYU1VBmw
zOIgaiL672BwsIJphraGw7n9NPlFEf7IkbPN4qXTAjLKf8bKQMhZbtprZiYcWd/Bi9oNEjchhzuN
L103AqbxOlGAWQByQokcGCM99Af0P1UCPvzuFsnEXJSes11RG825q80C5m8ImJXuIuxeHytXnlGI
K4VBlbx0LSci0CuqeDGjK+AFFZtUR7l3IlD02VFtlrgz9AWvHx0vLIae0HtJQQ+nCMMuERL1Ettn
5KzeWM8KDccbmO4WyJAuUE1WAzc31kLcFLWWCD+g3P4lhxXfT3+TpNKbi/2Gf7idNRnOOlj7RKR8
J5beqWcjqAZPzEmMm9mj8rwzjF36N/prsxGbjlLpTOR4xpKOxuZGvzlWPpyL+VsZ9U1JI4T6JxX6
nWAwHVe5Uj906tyxkoO59DiQkDGZTRPJNXu9sHZl3xRAB4bnNw0vBBMixCLr3qfwTn51l+KZ/LaJ
wNa+z7F45+vL49ZgO/eAGm35+Wbe+45xtvzv4VAWR8Y/sHBI53Cv911wYQtqtB5A5I03wplaLLwh
lDLDpaeIDvUIQwCB+aKNsdzG3jdeEGkJpH+T/JcM96JsURHiqyJgQS2hz8SZRfYovR49to4w23TL
Gm/oSmVjqSdZNuS4QmVq99VFnOzX0Y4pNx+PQc/WhrCepO5rC6wtM2Tqm0lqyep7grVcihHWqrGO
IkZ87WOc0HhSVawl2vrQVQuInEWOTcyjzW4MvZ74U7le1om1SAbpNPIzbu1v7CJRpu/K/fNSqRpY
HwZX29dPKc9TFWdnRlS8pfeybn2uN6e+9A0iixk17qZChe/LXGoAUpGEgeir/gs6oQIjEZFO/Ig3
7TryWs7uqu2On1KLcTC4LIV6bzEHri2axEty5OdP4ghhCyJMPqgQlJTM9CK0WEE6Lbi+LpEjdOiB
1yWz53x2MmijmUsagX7SdAYFaJFQxw9fHZ4fIPF8s9YVZHG72vTm+G1CfrZGCdb7r2bTVpGXrOQz
smztgNjupP4dH1SDhkyl/K9XuwjpCSAklWfS41CXE44v+fuSp88qKZwgI4vtPk6b/lpvYXFNzDeR
YpBcrMKOemXYqsvlKBMkHz7+F4iU23hW0/4I5BuMjjmsFfR+tHBEhCzAdmJthgUS7UhpJ0ew8Z+8
wRuYtn1mVkOQ1Y9Xijn0TQd65UnWiP+SDVy7J8amxJpiz5mTsB08BxmMNTbPGykVJA2lDbRnQcHO
3QMK8e4OzclVe/jrrH1XEW9qMsT9XRRXFGwAbYlKspHBDar80n6JcJgNlNBAgTNdpHAYu/3YexnA
Xsf08t/SEwWZB6g74aR4tBW4s2pDqr0BSvMZ9j75DiUiMggwbR4B21e1hmG+/6H5OVs2kbGa/eAh
jq30pM0l1moO/JFf4BQpjg8NnQNDMzzjfVr9c791t8JtlOVmiSOtNtCX6CtlpS81jbu+L1LGfre8
iwb/lqVq9a/eu8T5jW06tNUSmSn5g8fLaEGOC3QSxJyw7EQAPbSk8YkOI1XuzMZ/5EJJraTjlzGd
Ecie2bNU4kGH7HVpTUGqroh0wojqNsMNwJ0CMdkpOkUMEHJPIOIj6iu2Tv+FMIt+v/G/+DTzQyGB
rcQfPLG+/WLCR99hGuGYUMPpOBObC+2ymAeVtyERaaK5ALPA/ED1G079LFPYGDvbHgEBMc6QsGfv
OCcLwUg/m4sZRGxD+NlFiOmPl261B/0F9bmICwaB+EFNJg2nF8sQE2CD5Q2nPVUHi1DZ7+9KLBQO
0ySwco54Lm8h3w3KMIfgxuFvZ3g+RAGDTcgZUGqWNIFbAxoFX9FnFW+s84XEMt7rNYCJPF+crVxj
ZctgYGkpl5wC4mNv84BvmJZIV3UJ9oBnQMch0e0/y1Kfh5kRw08X+0YSgeYijQ0Xn7YSBmfH0YFP
sY20Sz8ic5Tnaeh7VXQZ2glbmI7MvJwN7Ej5MCSC0P1uid4HSoVIfA6XP7KSgL9bCWqRIrVsHz8q
vEJBJWyAtR4yTGqBdEYl4H5NMwuHBa3ZzRVOYVB4J7DgQl6ryR1RO8fjCivqoEDnbSJE6U5nYpq2
6jntnXW5CNBbKV5JPsowVAre5pgOzxS1uDEm2053OhQjepGO0bisUVbxwhxr25s5uSvdpDOZRlwC
IlbjVHg3WIM9A6/PFg/XLEbDg/Xl45AOsd+fxGqvWxM8s9i1G4fvSg4tHJEJ3BfLctS8dazXULgZ
n3t8IpnbF6LYEKUHLJ4Nn2zMhc7X/qk50Un7ih/P2xF+Sp0DeOMCmasR91MlM/f6H1rp3K2jRxam
KYrgnn/MnJCI8b0ehtpclBgock9hgdv8WX0PXGo12kUt+fAGtt7JxrQHJNL4jFmJs8u0EhCL5RGw
ikftB8wUf8KtcAH1LJMv1b9lxcAYV3p11rqW862F8rkZtaTCG3Ncj+90h8F0QnuGvRodoQA991vs
lHtAschb6lS8gYbggoMs9ZloCgYuv4lvfks+c8pXxI3YB2a/1k1ypuvBMS+Bxvc2ogsy+y2Ff6+6
DaPQXm34sec81LzD4FFqbkRagOqKEapjbg7hvb7+0tBN3x091Ed5c86crqZssX8/+Hm3TeELZkV9
nCYSnV9no480WnQDK9VglGTWbppeoehGyO8TiLyRelWxPTjuTvq/fJYLZbv23Gi+8R++NzddOTG3
RGjN6nO6f0zMDTZCqZ/mX8OR8zIZt0KtwoyGOv7w5xt60tBUkjwdCcDFoM/iNpBaoAbd05Hj/mee
a21ZWK5E2a6FsVNHy/7pGUU+AtlvOSozlK4GaMHcxA/4quuA77PTT1PpDfKLNalKKFqNmWxIxGnA
dF8V2EKNKyvx5drgZW1YzTDQfuLHG4CJeryy8kF7K2v80Z2/WVaQym45GGSsyizdHCkMor1biSyr
Yv0dSmPwmveFqlJJE2SnPctmPr2zySfFys9+Xf+qBllkqmHBnUXzHokzY5G9jblfIEyipmQYD23j
oL8iOZ9An8qcCrJSc+llIJAC0Pe+orDKLuleoWJVihcpcNDNelS/uIrR7wkRJDGbvvjbcggUFqaX
snS3QZG0LyxPTagKCHJg/KTK+090rQF78IM3Ik/M5QGphYJKJcKJ72oIN5XNHH2nFDCkibr6aiGd
KvptSfA/2TmL4g2r1YhCnDQPOYKfSaU2mSoUNBAHP6oVoXnL+CYMH/T6BmDx2mol+eqBX9sWzLHp
JhqXKC5lLD60rjupjfPgdzdDo+x12KTIDInqjHcqECPAGli+S9lPdXX+CmaHGayFBfxeG5GFYIDi
wWFK5smRQ0fTr1hcv0r3OaDl1dn/t0sEFIWFm/G5NEyLJaGDu1kDiyipgbkTXYBap2GtBU1prh7A
qQ9/QybyaaUCk912zvmf7kclN3h0AzHwytdwugHEaxbklmpxe7naLkGh9QrVIgOEgNZ4PYo0x9vT
VtZNF7yfosT32FGCKrJ5oSqi0miHYw1DjRaR1e839uBVpPm6SLJaAQcA5kuXuEJx1W1kPH4lUJz9
u9q0jh5iDRpBDBYGS4MkTFGrwj4vU9g+V7mOyecJ42zTagujjNUzEweWO4ypU/d2qopN0bRwFHM2
udqGWe+5bEcmzZFpqv0/7hWV6iX480+hGgHrVZp4U6piEUCUJEPPyDbpCZvmqarMBLkcu2dFywGM
SCHbo7pGfwXXpqvo/OCDr8wvU0xGNu81UDhPTpl97f4vcvhDleJekAuJKQtvzI6EZ7drL5FBPzgT
s+D4wEFFjkwmq+zCDppkiIIqUY+fAH2LoQKsOj6sTgXevEG4MIrnWFfm+Wi7EZLHP2b7uuIcO0z9
9z05VRBnHtC1wmjRP98dQIO2ZZ0m5nxeFHH88sX3ckOSguHzPuy9qt6eTCAaTNrScN0CuL4S30fc
Gd29FUHvGh5D09IrvpuIuwFtb5RXviNbp0t7dYCot06x3LugZkGPstjZWPZOeWDPlM3pkiKWUcR2
XS+KMhlNQNaui6hy17FRDyNHjBOMi8V25XBLXjuNydiEO0zCZB2+WOjKvhajoIjDFuDTglkQIGYT
GbiuYbgG+hpwA8oz/tocqcH1ygJ4+8q7PJ/ENBcYXlfoKejTaPHqcHG6MIPKKTw4GsShY5iW9+7o
49WjNnqStjYGgilreZW/zf5epDdMS5dG78I6mHkUppNqpW8e6sAEZC3rJMUIQ5npSEa39Q3SRtPo
gdGYhP2eZCS8Z9tZ7nNfP7Up4OmdHtuiiovR7zAELMGGP0za9ByhDN6xlFNrU9wtT9BVp462Sqr1
GpLhvsw+sRjsCbTJnvK4If6Pgy3DN5hpLxTghincMXfxqgIFcyMRBk/hh4lUHlcZK0sZ2Y8V9MCk
MFi/BX4NrbZW76CblwUS2+2Aipsb67GVhqX78eHtTjWfdkt/DfwnFIKHDcqyapgcRY4O+f6VBWa1
CGDg2wxgbc88ZYcqbNast3fV80oafJFryyJ0sdCr1ocenKCTJns7QEtErVl+5WjOE/naQVvKALCF
juW2GYiSvkGNdqu0KWRxIeAvI1346QfBPakkl6KpcUYvQA6+A1YPqKCc/d297RyJLE0breHEled9
m9cxHmcOYhBiEo8BitVZkkg7NE/ZG6iUxYbJa3vZI6iuv+3s57+5L+gC68bVIdSSsDoVgsefkmch
K80tXFKz1SLUPqXfup67PrTPqpScaC4x4+N/Mt0hCr4MXiXK94cF0RgYOO24GMsTTssbB+gNfg6A
EwBSgCnKHxWKXlNLncNAUDkT86bsSV6XDl+Fs3c2ynN0VKOylKhdpy0Ju/6W/gFsegStVyt+j99o
WsPbzgsWP7BsBoUI8CZjWaiWCc494trE8lSgWa9YBKIw+8Qm7wVXZdij/6vZOj5+56T9kfapWvle
U5wfvgr+zd6yr2RpC/kh9qApNlTlQLXLtKK3+mPb9bJ8wkUBZajvwbRXudpTdBDvUC/Mh+KyOgsa
YL3j1ctqObUpY90dUTqtNU+AVO0ejQVNyPwcjYV6a5ICKli8jzNN4HoiEPbhvGS3GFqtaEZBUT1m
81aBk0pmZwziEGsM8NJg3cZACqqZY9eqvUSE16bVZbhETukdm0czwHu+I0FgOmgbt2ZarWVaKDZP
YZMBJxdGRdiYIPffLfKzka37R2h1VXrR4AJL/m8QdZCQq+YikfR1UUvkq65Y/BWbely1G3Hqj9pX
ojuRLAlEJimxX7wCPVheqmeRya/RpAJhunmMWAVUKav9t/wakqgDwJFU6kt7VIjVdlyJvnqTSWhY
BxTNX/4xVSelw7HkxL4HZ9sK7dN+HwTMGvQTamOPgTDkGyqKWHLmZ+4vUw5FdryLoew8XI0Fh+rc
7oWbhZ9PxsyH8xH9X2SyAH1Q6kFwckAvFtSMSL3XgT4l6Ls7lZQxO1pDl6vUwJ5Qdb07Haho585X
YUk4Tr3bwpdhWQJtSwoXtf1cMCD6KX0UXIby+XvTuzEarhM2FchIacfNO5DB2b8r0lATECVO4f6R
cvXinew11AnG0NLJYHrsDGPV24N7NgYAm+Dn1gKiAIiZOFrceEl42AKcHmr276vJstOi+N12qT4g
bPlc09rQbhugdJF419rC0eR54hD3K6G4VIivfWPrKamZ8OZC6pHcwUYgSyhJ0evK4WfYsiY38lt/
8bnz4fJfZ+1yuaqlQ9t48vkQDcEFrwrPQeRRH2JYoddJhlNC+i/PEUljGdx7/UzUPqOKBT7XKb+E
DnKNjEcy+WTV7sP4i3gbuy9DbSMcLSGOkMCBmo5Rg2Wjy0oXQSk+B/LNIsW+MKqU4uoutBXU17SB
/eISqG+N/gcudyL69V1F78FlyH6eQuo0lB+S3YeLbVlSpHfeGtqTPDBCxTn3LgTVfc3Po795D1wx
rVQR/yJreFMvbuze7CYr9X0YU+hnR1SYeiPV2Z/kqa6g0cTNyLx6aQUM8rgc9AAg8fvQtfZP/BBS
ySbXcxxPQ4eBxnVpfolOPhmNSu38ECjUhcMVXvV0rtqjIYuYUoVAZaRiVr9eE+dv+SDcaU5l7fP9
8yMIwP+Yo/VIhTsD7+KDQhCXdYK+UoJBdHO9S1PKDAnN6Ybzrh+5Pi+phMHy28VhIcfYF3E8mPlG
XtrUbtj7TtLzkB3bE74qOLXPBt1t2hvtiwopnhtontktWySMmULIJI/iU22SWn14YURyIKm56cPc
HXqXSAE0WSm74SAqHvi2oFxU+Zf1PB6UQ2pi56vIVwSFFpLVIqvpL4/vdBn6lfSLCFLRJ+B6VihD
K/l1jmQavAvJjQJgjZFQVD3Va5mJsQTtzQhae6hu+YeCEwGnve9fRew/TE2DQZr5MTOjwIWXhQxJ
bScvhQCDzupouDukyl6qlnWqT5VT57539T4X4oi90OmbU6BWw6Z2+hbi8AwTJaZguMUnBxlqHEOo
7e4C9vRACkSFvrqrAs65XyI8vV8+JLbLYqxjEWRAAslq6Vtj+2ciJaBFxceulq0FgQg4u94HGhTZ
SypIGlLFgSM7ltCwoC5CorGkC606HSeGlsrKqLtTrNj9tAR+MgYsb8Z4Q6rB423kvqqg976svBu3
XPvV2m+sQOzdDQsqKdnf+5f+kuCPvfDAhbR2+ybEwul1xPW/st290CkcZLfgXomhzCqGqOc53yOD
hoFKaMuM48Hwys6E4YnRbmZ4z6IXsz1+JEPa/mJfhPm/qA8B6vUSgrh1i9G608/Q/EYYIkaEBfz4
8UOFikr52kpBD7bMplvcVunlb/JvDNUTI45eUQSRIElLsZnHk80ZdCorfndtBaZ51dzA3K3anXoP
5AvbS4do1cTe2uPAPlmsp9lzqXIIAMnSqWhWGY8xA62TTLr60blCghVQZ/pLz2Tu3Sf1rDCmAFH1
qCRFLMt7XzvyhJThuTEz+3O9CU61Y7Si5XfHtp+Hnv7bnqDjE+t482PYqtslR5Dga5Yojr4bAi6u
T/Ak7ziLgG8zJId54ZUE8qb/tt7ReNdwXXNOodpCSy+tso3SW0vpshHDBX0EyVpDGwJPDdS56htD
FDdTYhd7s9QIcYBY1qFkLmnlvMLQmQaLNtRF9EhO9iGp+ET/Zf3y35y8wyzMga835U2gr4Wpr7ns
x1QhbUxdIHY0ceh0YPgv3BDbrkAQj3GG84gJx4aSdP3lPDLoGCdE6/rUdrZYVGcFrlZ7UZcO8SEy
mm8aJlSjk+WnB0jNIaxp/xS1XzcTqOBGXhpZ7zWQqppU2SqNElX3ar2rq44HTjZUgB/FyT2hM7ry
BtbLYkCpwkU+4QnQxI0Q6TbPcIY7s7QFMwbiM/9IRWWxj6LzruC8ZwuxqoJ1PZtPdIciMir9+si+
78U7HfqzVgYZyEm9avaZgzfY/lOer2cYsn+EfjFJnyRqm0qDaV01gKbsj6dH0Cb4VpgJzT2brNYc
Z+++CizUI8ES13TxTibcT4b9pYYAAYrQeZgLlRzPXwLLgb1SVnvxe+OU03WNRaiI4EoniDR2uq/z
RiQ29qFpwtSigjIZMdVy4iTM8Jq9VFLrQD0Rz9TwX4xEyjtewHUvVc6XdAm5bwra+hmulqORQrTd
ScJyWy0Ngur/U50kE62SGOgajl0qx3vDBBzhJa57qqioFQ6uMNFHl3DCgCEKKq7MbWHPC5oorCQ7
34T3E5mUzDoHWv+dF9y4Q1fL3GYAhN3vm655YlxZHVqoJ/l9xHvbY+6YCawby0fkBYoVyRmUjjPz
C5YDluEe3IrIPr99qmWx5pDOI9kf1QaHCPDrolvipnYihnVIDiFKjKXGfuFfajODyAg0phsEzlbJ
EzrIY+UhtRfPBNNro0/AqlGHiCkZdU25CwYGLQJgagJeqjee4K+hOj/UkssWoLzoNrCeCcfJzirD
qtkwILcWycTVk4SCYvlpS0TARnnfSRASECv/P7iQV/uxhunF2bLnhIOsclmATm7ZPm2KsRytfPw8
UxVqXaK8D5nfoETj4sXa8YoYHv1/n0sGAHb4w/rdE327c34/YjUAnKhgxN4XmCUvASkE4FEldoQl
asR2FQj3JAxSO6WAtoNbYbck7U1MVkZfZC6xNOBVhqJPf5dRaD8ZHOTAJFIY5YIBfT7xPfCZa98f
61VmEA3ciELWxuk2qBU+FGIFrr19GUEyEaCYm9pD3HI2tgkhjxN8c6XzIOJw98wWqnUNHcoNXFBH
ISUMpE5IOn57pBeOYoZwzWWOOuETz/gs+qur0Ybnl7JrGYsCAthgwR0f07leMHc7QBo3nR2N96I+
+SKe8caIEi1sWBT9039MGc9CSh0/dyirXJKLii/3VdpdbHJZ2gWeyldXMSvIMNIsJc+KOVlIaNTy
CrhldFm+Mz/yWWD2RpB4sMJn6uu+2WzLMJy1QPytZx6xCgPPMdACUipCuP/FljsPaq0dInz19Jnh
bq8koVz0nICY2UhCOiMv0m7poEMyifCfhtdHKN9HwvZ6Bj+G+0RTQtTsvEYrKmQKZBqh5xbgArWJ
D2cQK6dPGd1u86i9GbA4vW9qAqd6t3RiMEGneiBMZsLGGyiNo1wPo2Fk/uh+93hAYhl0Z0+nSZq7
ymnYZ5dkfPA3DZD+vvRKjsCvmEpTo3hKh9EyMjTdmDKDDGVdoHcBB0uiYC6r31IkOTj13GdD2nnv
PsEcoR+vRtXOQyPAzDd7pG/oN8HXYZOD6YmNtrpli5jViVWv2W+0EDHY/9xcFf7biBPFr9/DH+y5
RE6ZN6zc8X6wU1ii/7E221vPA7iU3m8qgPAFXAooqXtRroFfYKfis/VqEnvNPnfxJ14Qav4WR5Zq
3W8Aqi49oOVn8dg1/zfAEr7PgUuKRK+gd5IRN7BHyvQ83DMaEIRFfiJNpYkIE9j2tgSwvIm2y66b
U/kKUM8uLd/AH4cf0josFsP6eLFeM/cwVfffeDy1ILZX9nXVxhw7yPTek3vOiOkcfEMjnyEM0wEK
aI4II9GNdSZHQI9RClDJ3g5gjTgx7ldRTKq1Lu+Qx75p2lJfE3gCapjQQpStCcYViozbQF5bGfSv
FoOpdMBRb9hUMHoUyRFqtQ7YNRHGYnbR0gvMlMAFNvKG6GcSnt5SBOLnIpMU6jXFlfZk+ZGH5EEW
pYlzbahFS+NwPqFO18eXT/0IBEo01Lgxd5sAnOxKBTmNhq4kBlOlorkLKjYb/aHCcgX9Ov4eHL9d
us2bYC4wj0w3wSvcZZQR1IQdQHksD6+4ycrvfrjlbyfczWp2bNBA7IwDFoJceS0rSd+PBrfyUv1a
yUNmm98NVYqYe+NQdyGaDSTzSQ/yjYPPJGnvNfNS7sUf3JKf2gr2PUQm2uS48R5EoFmJGDIK9TKR
LMuVVew+lVhX3Aj3GOBZiaZ7zYf5iKy9UAXLPgK6FX1m0j7MV4OEFSnvTxAw+JJeLZLQlrw5j0FH
voiZeL38IU1Lp2zrtOei3u5j676RKRSZj5272VSRrasZAcs65Jiav5/8qZbanqORx/d8TBDaLY9r
m88wsTdIYhKmuJZqP43IEM4sG7whkOd3Cu89/qlszTs5K6O9yISJ5N2XwNLbBe0Vd1sm8iduPvPt
uIHtCIJFuq7g6zT2SG/sQPJvfklx6FELxbscWeEkbfCaN4cspN9O5PjLSwlzQ/xekufQvbMEONxo
rwZYuAQKzWZLtph2qS3IicEJMZgrffpQ5YQ0G992JPzzS2nHPtlRG/RZonttuUKxnjjsM01vXQfy
A1jLR22xaIr0FmyAJITmosLveqwguSMiNxrPvkWOLeZsMJJNRPmfh2kWtdut5xb8XSjSE1waIBh6
YF3BGOxBCI5qGQpTEVvh71yxKzV48QTS3qf9UVRRC7LXKKJke4e/ujn8OvC0/DD4aOC4agqp+P2+
ulyO7WU8vYq8uTFDl0CtEdNjxgV5fbx0hSwH9x7yft/PWb+TCul11AA0uUkPmO4O3fvGbobgx4wT
C8K6Hdk/+66OUptPM3yNchnUBbbUhCD/KxT51VnSiynuoAo/n7vyffJ5giF38IKdoBBaPdaKcvdI
/ZZjBlGdeABc5UdRNaU7JzT5sRrSF+gbkfgsAXzxe+KGRumEDjYp5/qROqLh1z6rYCW/f3NohEfG
6fhyyWLD/81PUHha0GaMnSmy18ZswrZ3CwutTP9bdEdxT5PzZKsKVX3br6SGH5erpwA1EH4l/gPW
ZA45nj7DHcZ/ecHKAq52GY4er3843hd/8Ibr3ODrCOobjgLMnUCjYPZnvASBRN8zpmxAPO+gp9q2
4S8KKl7UJgn5HJs+74QVYFbkI0oxePCB5hIcgoVSUq/vOxvneiOGjoFDl0OFP2LjCFd9RWtd+iS+
y/tcwSVdlV5kBQ6VomYj9lK48k8VsomjZACBEkiBHhfpJHo0ylS+hwqQYGpIq5aFrL22VTME9Bwl
gEmU8igZVPSHhgTqiop8MicbM9T0SFDIYk7gzYD+v5ApCWaYE1shNXJNuAfI50Fp8OXdGiBlv8Nd
VoxsdOux90C5bz8l+TUNs7nlw0GtTj5Whb+eawwpkAyTPWs6oH99yV1P+Gwy6EXNZvM+W5MktbBf
WWIpr+GNetkNJwuACqd8b8FUq3YbmrwLpMVTCpGDIQQjCjvfXTq4jvg+uiKeJWZAxPJkXoR2WFCD
zS7jWZJ4AOgPBky6bZm2zfSd8mGfng8XEN1uus/QyXZH6Fbjf30upUsezzKvDWQbEq6ZL+iCGWuJ
OnhQMWyn4C2bobtWclDpfoUl99Jpt25HtkI54iFZBv21cG2JDWugJf2+EO0ZAGFx5aUGJiSq8Ea2
klxUKy4oF0VU07MCm7tBTXQ1NxGR2DINeTTe3aLZKcV3SelFrxFJ+u2GtaBT09+zs31XvZDPiDnT
8kMf0RcwukeRjder+XvrH4q87pqd6vZ667NptH9vwmKDsWzdkRBZLtoXvyKUrjgq5K4frhvo5BoQ
OeSg3qSCSln0mJQzcTpi5udd6Vs6XVLgWWCDTc0G59ahAhTwnuEtO8lAMR/NkpBzLVdOMrrry7BB
+cpNhq8ZkocCAFgV0TVTPQObRj4tZxfoW3q7YjyjcWgnsqEyy+uPzJWxzhVS2OHPjnaJZ3WqpUYA
nAukaMsoAe/1yv/1OOzfm9/K2Qgg6Li0u4MmEA==
`protect end_protected

