

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
L9EbKuxxzV/09pnAb0OGW9DxPQ+o+m/MvX4x5f3JCiR63+KWt2eYB17k+9mGgVY+K1VLxoYz0z6V
YvlDefublw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gJD53XIM6IXGcoGao7b+pChhlJwhGxOuVwSTI1iU+aaEVIG37JelabzUSiGlwgboK2Zv8N9/EzBK
Y9pDSGcMvhlTABOa75VEGmta9QvVzRVMjXtd0b/jrdUkZar600zvkPbB8+QESNshxT7B96klkdIo
XvMdlDR/SEQxmh4Mkpk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uMh613zg14bfl9MaiMXKdALr5q+gvlBiCCfJpnudkmj/VEzNaqE3gABSgWbIJEk6l3XEblsHwoSZ
2eueijgOoGBjZq9eDXqLeir52M0Z4RoybrJFqX7YgYE+2quggoW8XJjUPK7bExWH1Wd6un6XRwZo
+XQ53VUhkTgctFKNHRr7bEqxJa0qk8dm+fTRKVmCc1Tr5X6rd28yRrr4koH3+liBwEPKquwcMKJL
zK5B0g+bSiHJvGXlQQpKzQNF3+4MebcveUUQPOYG2FAjfRJs1t60dgE73q6y3I1DMI/3MguCuvoX
78TA3nOFRYGLkISVFXDX28xYA0EnciH3BlzGiA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2ADp5V47yVkwRII2+UsRY3zvclviExupZdil2h787eVOjYg5odQlZCOMnldkarIbxDBoj52vjMGc
rG04pAKa/Z3oDUnDkDe8ZMmBI29kynugqgc8aGxYPVKp3KD8EvhnicB6/4Tt66g9A8WsjHtxXLuC
0ImlGHU3T8u48JygeUs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s5k0DDcwk1Yhkk6mc4rW2ITc+jBCojX0QPFrzARjmvIjcmc9EJT8pAYSdJK1ykoSIGmT8u4U6vaF
5pchZ1NWV4+0T78Lu7ir0M6lHPYDFRgXZTR6CNdPGqAe+Si56W7NnXEM0Yylf/w4tAQ0u+05yvCg
wK+mPCq/91Em5ZiPcvKOHOdJBSTTkSYC7/n0QNniR1mBmd7+dgsFr5yshClYY/q8HngDDE/aNYfx
P9AT4ECjL+OzARXCnbTA6RjbHEjVx1ewIc83WIXkwbZjUYAzp9rYNjFdx68zjq8U1XW92RXAEXCc
AYKv676uVGq/WAryucxGApaihL/izu2+HGUsYA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30640)
`protect data_block
YJODPbrWKeoMTF9N7yi8Wpo9IkKVryZEWLAXCTzdzXTiLYKo7DImx8QBWoQHZmqV5H6u2ZH6Ta7m
ij0DnTT2xLXCRw3N2k5dzHBZ4ErLeFxw0T/RaDR7Ovzi+qOcfxcogGHEZySZMlEf78HnYMiA2x7W
ekH3K2DWC2ow5+REmLgtOcpP2Ao+1WxXSMMFeo0ADw+zzSXFCk1X6VMOmP/BpXQ35vZ7a5w8JhCj
zyehiIReua+o3Td/iiZeTqdPIaSm7Tn5mw2bwiCBjhc53ZrgVKU+9RUTm8X3oGq6MihuP1c1lTai
CoweJhUWuuEENoNhkJnfz+/PKbLOtYLk2rI70ueaBlToGu9n8zvYhfj2OeUqONPS4ZUG6+bbi1n6
5M4RVDQEQx15Easy9xkrubAB7/Mxgz4U3cEsAT+KE1FPHmYtGhehefTOnk0rAdam0MOkefVEXiPw
jlGwm8A0qwpW9Y+idc5T5OZ+arGguHzNz1bifMgZqipJhb2NJcRoWQJtyQW9jexq5vKzGxSq6ej3
6A1IH0PX8SiBInKSl8SJNtlk/3u+jXDmM68aZ7n6yrLkdmkHIOjILaDQdPoizorL3ZUElknHQ/VE
XkiuzpmLYjPq4CSFXLJ39NFF5K7iY5u3RbhJGPyyKZUcvfpDCtCi0vpOvitcCDjxxECfu3XKC2lo
p0hsixBmbwpMBgiEvZwBElRrwwtZbDUDWyzw65ewMZ1tnAjp3w0Wqg+zqZVgNHBK+2qWH0hFfQzS
bb7Ttp0crkPPw6P9seGytp2FuqDsqW0oCSCkb1FhHprapItLQLxyA6ZXV/tEDSf7F8LT/8G6mvUe
9P72gJk0eNFgXaI8CuwseCMKlfOvW8v4/W/alJp7UEkAXXj0Djh2bd+2p/pqhcNR9AItRiM8mz4Q
YyzY5GTNBiq9knWt9pheqHHqJUk451cSEfw8+5w+HjoystrzTEuKx9I5QfZtfNJIR5BA3W5cw0KX
HdwIXbJPoKpEHQK4d+iYXNn4BSeJZKEBjglmt07eKFO0Ekv6E5RdkV0xoVoGYo20MTW6XLa8JzuM
MXjq9WlYQGZJxaUEm7FDCAJp5Jekw5bOB4yDMGqldA3omM1cAb0nWyJlEWvr59yKMaBEymkjd/fZ
UrGYPksmw8tqK05K61lbYrAtUuBiw4MSrnNgDDxbu/n+5NNJBql3fv20aQydxJji1rbTUfCaieCg
V3fkcVTvZ2zSzNc3ydH2y7MD6kjF+nGk3St64axfwRpNl51jALFjDh8JcslaLoKwoWAgD/B0/p5G
HT8ELwZaCd2u+/sN54QOr1ZilORzZB6RsN4ft3npVx4yUtPCyw752PsrMILK8YnTVsBkvS6WNo3/
k4J3FAWMmpfHETsZQCwxRGCRmQPqHY/ueaVJ9tA/QCBxCVI2mZNiuB5yzVb+ZRvyGlBlPRbMECeA
J1ULC1ccXV4pdU1k2P4eTctbT1zPtkV6IU2ghmYZLDMXEMkYxGgROIPR+PyZSi3D8frCnNXPjWNd
GoDRuGO2W4HhvLrdWHAOTRj3mnkiJgJmCn3qzLvfqssz8qM5+8vEt67gmoejHDuoeUKFC5U+GR2G
HkUj8O7iieibeEinCX2UEdZyTsnPmfXL/n8LVGL3NvZJcpJhtdm+Y22P3WuBPLENUvroe1n+roYs
bH7XbTIj50WLxLCnfFuIE7Uqwvl33gQXH+mJO2L8+F3TZ/NfhfsK1cxDU9l8fOt9ItWURslaWQGy
bpzzdqFFd1pDSzY9cBo68DoS2sbRft6LMtsPZE+rSWq3AB7N4WEyXL/+qIv6jggZ1jgKGDFUzLQm
1+GoAYvKj8QKP0xqWWh5cZGLkZLDjIQIcEVrDtN1lRFsu6C2QEQFQSVz1K0ZBm+mMGlazqIFsZ47
12sDEd4ftj5yFHjXOlKdDHykfRnbq3/nq1/p0eXOW9e8bMAo8gIGuQU1qRRJdlWVJD/FYsQfHHDf
CfLo9nDq/sF7MdOAyPTO5rhf7tLUJalp/q7rTA05RcOzQ9uhNLXIVP9Ws3cJvblNNC/xqiZttshr
QOwbZGOtNqPGfhwVVM+3O/e1k4nJjii8JLe+rUi+b8lBY7ZlSSio4JGdSib8slTnHb50BDvCHD0b
EOozSKdHCkf+Kv+V2haYCnI1IPzFaxR0GW+9kempC5JKj3avpvu+eWCiiwJ2t3luGALmQ7rQ5USa
OKJKMvKdIOUiUSvElHRhgGnc1bfSPOCQJRiYJtZzoMoSkCSm5Zt47QsFdpV7TQBZgfHqxD9hf8Hv
FSjeLKc5FWV/+Ox5VQN8pg4s8TfLatdbGZR2DA3dv8sD/z3jDbnaVfGBLQnhU+z73XNsmeqS0xmR
DeqxmpatGJB3ju83KnIpPudy2j4BIVAhU46xOz+8LV4meiWj9cMzB8DCZh5GEQWdUiHGOebtoiHb
TEL4ezsBVFdnGfYi8ZwnlrNhpdSGWQoQgxSQqdHfdjig27fbYkm4gOVGpq/1TAoiHLd7FJ1dvnRC
34klJQR9e5IlVgTdSnJuJpbIU43PTosAi/K0LAiGLcYv1xp+KkGZBffGsVjMy2l8lUZjwU1RZ4Ft
c1NTkDRbBEtvzdMFDku+fIoajxEYuhAyvQO1W/T3mja3X8fFBKfP6Z5BsZ2iTMvRoIvhcgFzbyv4
HxzLCHjtpibzttA6I2dtwbp/2akw0WoyR5M/A8ILMhu7jcZBpLwASjnsSUdP7JoYhc6rgR5+unuO
93XIq9bRErwNVPOSLN1/LNp/haWUxViwJiRT1A4wPZpV9arWVgduZkpH8tq5epGH428N9TApmwSR
07B0ZwNnOOIDLrZHGDhfTrwcNad4uc4N9ULoYYZWgXaxC80OpWCwpOrnnK+7DU5CZS1nk/RPbCNF
NHJ82JaI/Fl52iyHVX+GYyxt5skYssKlqYMu/fU200Aw6qkDdnOumvvrJxl+BsOgdebgIWvbqR2j
0yZGd0+LUawa8ghxUoWWENOS+dLGlZIA4Vv4S+l1CBotdzDmM0cxZstfVBn8zmRdJ8EkE1LaGW0+
XV9bq5h95eAGTy8VMrsfv5Q6Tq/0TZkekfZ1wMtQC4BY1q6l/k2C6gz1h1Zgso+ERUv9gr6K6yRj
Bb/CpbaS2dCA2XuiZJBHJD2DrL8q1oM+pslwEHQvsFysZNDo01D2bHcsFuGtMAF28+NT8jl+Yv05
bTH+SYLbChSZ/FxUg6zJx6QQgK9pEhdZ9aUJKB9m+oHshdAbqYPBQsLyfH2U+8ehLgHZ1u5pHXxl
8563citjoYjluVkXLdBdP4WES/j7dOQ/+y9QYUmpZf1ndpudf8PWaje1vYTgMTTd8FjH9l5/OnA1
xMB4wVK4U7wbxbt8EEPPvWr16areCE0152J/smoKNrhuKbv67UU3FGtjVrZgGyEkcPsqhf+HDXkV
Y3bP8vh4Y3cje+wFyeP6JpdZ+AMlBJ8OFpMq5ASPle2TFLSD4OUsn/+tv5/+aHjZpFNZNAfqUL0G
pD8vZ44nQeXVbn2kh3p+Bp1fselSODU2knNCk0eod69TroPqlU00Re88goBTUmK1ot8UZ46ER+hM
6NLHDTMyIl1n6piF9z4W+iVTNwXm+WWgQQop0X2+58DXGKMblmrcGitkWiHajtoCM8M6Fxfj7CbE
D51qvlg2OowIGndpUvK7Cm28F4wI0KfNaphPDuriG3HERpY8e9gwlT1Ce09tBlo/PFAy+h+ot5Vv
3MRX+J3pR0sACYHCHK/v9t8/PNwxe9iRvhClYiLky3Q/SkpPVqKY3KLCogZ0xhyAjkhpgwzP/7so
os6ehn6YcploRZbc7klVJ66+d06uwmTvfNhH9HUnC4QyNMIwGddN+MpP7O/DGcT9DnRktxkolp/n
n9KhKi6loAO1C6jdAv5FmyPohj1od+v9Xp2qIxXdlU9/4cuDpcGYgOSmfobjvOvJgsbOBeyMNJ/W
rPB+jufjnCIAnNVnU0tvwt+uQwpG//F2WBv0eR/guHgqxvW1IRSMyzLoUz5zNAIHqIO3em4jIboW
YrGfJMd3Pu+RAjjCZUr8fusT+52kCsdqHJ3++6J/YoP6FElhrYd11N7lP+saVDLVAEqqfpTQ+9Vh
JO/7Zwi8COkQsluCzMfrSLPv9Q+/3bvjsidJfdNn7lOcYcFVwd/hROErhao/ZPzGjT5VcHWIY5Ks
I7xiShQALiWTI2PyW9MOruR8rkEjPXDQsFcsOCIG/6DAhskdOA05n6QXqiMvVoYCi07Kjc8PBwHl
c4GT3TqzUiOjRUQwd73hVwI5a2tbHzXyQwgn5oun68wWs/Abh/8OlPNoASLNJfHB7+Rnv1viRGxn
Vl/fKEah12J+in5lIOElQA/d/ARB9FYno7Wl3D54KnyCyZif6JQPANhBC+KiMLAr2CYiB1Z9BcYK
ZaQOMU4IM3psxwZrCWNANuPzxP5DNnojhUCWtIuLiPGNgmXOfcPsNcQoo+8bKEenQd9b03sw04vb
P983U5uy6rCxOqsp3NLg/8mWU8qIJNNU3T+N05NeaalfZGrEILWLQCC3Quib/WnLUYDNNJuasQDA
eG1oHlhu9N1H3Gv5UEabjx+KtTsF6So2vg+z69baJpXYE+MdO5hZkDo6PJarRgEsj5ZLDmSw79j3
TciMhbWeBdDtHWyxaP4P8/IMzODkzwxL9TX4CLvLcgaIDg/4p+WLPX6yZ9rThRUu5OuDy7OzBxtD
R6DZvX7D5oeeJv5kzsiGtX9CfOewuyvb5SJxhAaMzkoPXOn6VVC4k9l6lZHo3Zl9Paij5NqyGDwQ
za6tRhnwQkVOW0cXLLtSyuPG44vrU4QB/a76jLqTQWFzCmpFsHIVmWFZODpogCD0RLtd7PiH07cy
xqMA0a06EnxmPqtdbyRoSRrJIQGYDsCSjdLwHPptsF17GRvCt4LrqTvQiGBcLY9MW9tFrZipQsIM
JM+gYgg2PEUR2QiY8dzMz9mJhPwB+JNllvcrPcDx62zrMruSSawfoP8NTTxc2tcJrK0Rtsnqx21U
ENGWVTl3MPaBocUNN4G6Qy9MtO8i/ZpVyPQIPjmm3H7Mkw9VnnKfSruX7AA02lCXWS160BuvzKyX
a0VDItSyUlzqvuTl3xCIpe03DUtfDZitXuBPf31w0OKKnvnDsFYa/WGbBU+TTg3IkRAbfnSg6oP9
npIljTbvfibPgSmAzD6RSsLBM0Jr/0tTFQMV2v+42ccoy2FHxZvbCZvJBon3NTNjVHzYfIKH8EX4
3lX+AeoCqrj+p9U6sGhKHGsMBrChqCLOmfnrqkI8chr6FeoTEK9FwAOyJAtZGtwC153avmXPy36J
yYzAhbcl9NnzmZLVXUO+iHgwiewD1x+U9RBgzubeHMwMFQIn7jCpqt5PK+BekSL/itsNRa/Ku66T
Cq9gm97H3CI7ldPKNR/ZLKLetXDdjhp/zhoU//Os9qt4i0v7JTKE624+FsOOSzosimeC6KpGQA7c
IxhVZnPhbKni5s7zI3ejkAidISRaMcfXX9bqnUCmeaVK2PUm0k1xN2Aabl7YSX2d3exsdbpxUWsv
j90QD2Wzqj+nsmWVuc4UFM5qPEXxooonoskhNyabQsOmsj30Jf0IpaSTT01ChmeL7n3QNKt5rVDF
GGRoOr5eAP7NGFiW97HiidZeXlaSO9SUPSpD6UdA9HZCXPzf7h1aqdRmRMmWqEDsQw9wi8U+zqOQ
3Dk7tj/dmETsWaUAMH/01NE4IrzTwfAN058uUj9ZKrihsPc8xpUadJcZ3T3JG6M0Cpbc3o2AHYNi
OptjkiFJMvOyoxAkD2u+9F5DaZTUt3ExtaWsVtGJAM3Z0LOZEGae80XfT840DSINNxC+VbN1e8nQ
TRi0fk44KoP23KiPNGotDRxoozcx7Mip0ypI7SYq2kOR3S6HczUN64Qco8G31bVSJ5emjTW02v14
mTNa8eRb7U2Xl+IOpOOH+TSaScvCm+yXhu1A209GpoNqpe71L5TpOEpWTpOT4/VmTPNTOM+VCSg0
vFkS+0ZQvZHZbqx8YTNFa7IV+WAIoo0XftRHEPvE4AbhKrl9mge/UQtGBo0+RM/sINckl+2QMFGM
NFxJ3qNVyaDjAISXI427jKJllFw1S4XpEfuVmrFand2QRVWmqTRKemP130mWksGW0PKV3xPaBbe8
KY5VsALKGLdjCWReOQWWNpH3F4z6DFoYCLSESLp2eLY0RAymZvda5E+X5jUkzz7V8rGZ2l3aQUdf
DDLetKjQ9LsVRDOHhdExXcSh29coABprNPqMlGz3CvtSGpntrDQO+EhNZU3trlQESopXZr0octgl
Kdh3Lb7r6ofTbfYit8cxFfv7Nb1n5Z/9zNm+DpubIGl6qLoYMSOyevQaa7PG0309sd5S1RyfcILx
MeEYWoJTkKXXyZy1h6TDtUwdJI/HpoJPE2D5jQzs2UJagOBAoHgvzPafzeURSMphMJLbrWd+wl8r
mCx0FfG4oVTJmMeF8lJ6DY7nRTYRleZXS2JQ1YnE+Wr6Muza/p13ku5auKVuXyTxozLf1CxdZ0fV
YPymcsYWSCILQZgG1ppahWCE7JayVMmFGmEsprmkO/Fz26Af17b00VK1leMrR33asAUEYqGfZ6rV
hNJRcb3Mb1Y8zejuSTJI+dH0koGGOr/Js8vXGwFlwnTKLppxXVsfBimniyHHbXu41CMhHraW6oKl
q3mlm1Y8CNqkmzmQz4oLFCeiZKLF1K8z0/eoFjgvhezUaelczNeVqfQUrX6BDmQlz+EmSlEKmBBQ
Q+7hbJB1le3otpaGqYKyhecjvXC2unbuS2h23PXC0Qs+V+tXStYt2uBjkOMsYAL/dJaWt9ldHqgT
I61xInP1lNM3aWSPQZZ1N/J+I2F3Wqkug2mw6npBcX9xXB8tXM2/xsFmHjoscybg60yn9+ciLFuo
QR/HjKouiqLWobzDbFnNDj+tMb8eBoaj3SWbpl3bzabd1y4wYetCUGbFY+vkXZR5onSL3gJmDlWn
jczun3PRAFLRqNplaEJiwGhDJrGr8cSMaNQIgEJfUcb2mYPgqzTl4sSXcvUHoCt0gb/62OWp2iT3
V2Pv/6mZenEHn0zWJu1/O6OYe4jK2js95b9PJQeolhgAAUIjeoMfsnJv6RgqqSKixVo53dOS60ck
0yoPyqQAST0d1fsO0N4tQAGQYPTzcd6imtRlfhh902vzDDcWiuRoLV2Rbw3b1l0cfC6eeaMsPfkD
nDtTs+MyUScVO3e4LmyqwMxL2Ayf4kdF5yS7Xa6RIdMOjj6vbF3H73Aehb/xZp4v01RyqrwxUf+Y
7qCFNGO+KWSTjWUGquS18TXmd4fhocF9fJi58/MaXfNFX594/oB1stalNPzCN2NhFaCvaSbKjIBw
E0MhGpCMPTlKQ9dgIgQVw+j6sr3h5jmt7TpPWBm4UfhKmfLtY++863sRyTry6fcYHPziDBg9ts0W
IkltYWl5YM0Ebfn3ugaM/lnGVY6uUQyMOyo+z4Yys/jnGYjzLOWegwp551HwgPCHogrseiBJoHi4
OCbdKNwHSDlaZnMRMKlM0VmZw5kdCTg8gU+LV8CEAxMSnUQuint7As4ZK33ULcuHaUMiFzz0Jj7w
isysOledyiFlg80wCtgncFWg/+uuhvDCNDz8Z9SbqE35Qceq60OjaWOYP65vzcOyWIcv8hBgP6W1
pw1J83j6T7gMvPNBYWwA/p7+QH8FTVjZSuwVGHVwAl9tQt6XVFCwicHDG6JunmjTXzdd8e9vfqqi
+EKssluwK6/AhiZheLwp94gz+2eBIdktCJNZb8k5duYFffoOfEgqE5LNiMCFxPwApP/0xpvy6o84
2NDtNyKAsrZ+VQWcaS6L2LPTJx0lEe9eVK9/qQopX4H75NQf9hGWHX7lcwMh+qTkrGfi1ozUyQ6O
b1tVwO7x4FKFLK23lTrzijbVXw9xi1Mjy29JU9KnxRee1nC6O9zL5SsT3Q3Hc534bWAND+KLb97w
tjlf9WbWP6hueqR1oOywlB96Nyfoe4rkP6yV+y+GiMsJCafZ8TDQkZdQq1ZeizOfUlvG3k1Om70s
yZPfA6VAa8u3zPmvZkZ9gSkqzjahWm2mkoAPY3/cqNwyfRQ07gmZIZjFbNERPZ5DCNEiudzkfbeb
EKHMpZUyUrZ0GalYYtdfMTYQxsowcjsWCv8pfzASFFt0a/F4pYry+cpexLmjODjdfoK2R4W2Y81v
YP5xdSun/0hZOFrTm6zyKeXkzFIkud7nFjDWUEQm/P5Z+0Rqk8UaY/gnTQX/sj9tCCG2/0zFxBvQ
z2LVIVb3qJFIGxUNih5mM8kR47pL4Tw5uPLGT9QkaF7rP0MYzLdmz8FWKiC5MOf+5IZiqz4zyVsW
E+7fxLDvbYxOm+n3tuILqqmSdIdsPlSCYwtUKpcrpvQrdKswV1YZcfHS3gmgrh9tyCqpiuIoULww
+OpgQoKDT8m5eciCKfH8tSjvdy54rCip/7tjsISknUtQ0VSAs59/7t9CdiJ4bpZ+gScoPuzreL9w
/jC4x9v4A1CYbUUVlhqXKnpTj/fJwpBtGWkccoE1N8x5dX6MUZrVHFYqph6XsHE7E68I+V+l5xiP
+UYCZqMVakdrUOgEivbGu8uaLfDHvvrNgcFZJ8RnTYvoRdDLsRW55ka2Wmw1tl1rCazI8Mqzx9A0
0O5OUk2uqWO+WhRYBtnRzPW0Cl2eDPnHBE/r7MmDqXgXWX8i6G2Pi/zGAnvYv+Osxx3gf4l/M7sS
0S/Uy2Cw4zqDwwIZgEuj2lCd0HHJICmgGjcVYj4a0G0Eb+k60N8lXKDfUQh45JgkWpMTEEPKDzJw
TM99sRehfuPHN3IDfE8hiHg0WJzW/nOCsCkc7r/A01uYpXVPRyIvZYxDgcnti603EiqIOdF4vz2P
MsB5uQCw8FQqwJgsYtsfp8D96GsjVOZ1ZfXqNZRZKXLsRxK+TqBr4hJMMN6yl5hY8zL7trqABDzv
F2t6cT31v6W0V0yPYnELgiDci8n6Nxnds7t/jUDES//PvZc+9byupuXptpwpkhuDu8vJ2QY2J5iK
HOev+Yopyl89+FmJ2GOHV+KWaT8igb4g8+K/0Q8QKbDVJNd/Nzp3jHDPIzrp7mGa/xWAk+nbvAEJ
imuIRrutu0+g8mYGJc5oqXrAv2InzR5LGLpFS9OVJWaPdlXgY9LDX2cDhzoAN4FDGDNMKe+wI913
YjEIT7VgHBABo5eIkv0qA0iJeiRhtM7sco0EQpfiPg4Hhv56LRzNA2MtXhfNUgSj68ouanBL8939
1IEcCkIFoWIICDGGuN78j+OKBTpBiJuR0bGpIvhp/rq3pMzhahZzKXnuIpCPX1Z+o4zadkQ3iDjL
3dcRApIjZ9D7++8hrVyQQzBs96UL+u0G+1IeRlRnlnhqgwSvkRnhZUP7X3wsgd7RaoNMMlLOovU4
c+0KtRCityZ8Hq8jndGjw7xBgG7VOqhstPPufg4yiy+3AE8j6Rd4tVbTmh6Tsbnxcz5GF1YGAnw2
Bmlpd/liiN5ZcE6I9v2Eh02D7iDLwg7tZEALc/8/aH60svJRjZD/R+Tb7Dmd8ZYgVr9lnTQh3J7z
a5hkMLTJMltBHcC+zZVih9LxqU/OP2xqJPmdDIy8OYyr87Yid5uy2JEoKUvIwwW7idcwYW6+D/Jt
NlKoYLprpV+QwF/W5C/SqvhqqjqSo2eeUzaoBRDl6P8JkvkK1LcVCDmGq5nch/yXuAX6dJshLszM
X/GsF7Kq8h/623ocZC5h9LlqbT/sgw+mpg936lBDV4cqhz7DhmHHWHbg4y3JlB9l0anwkSet0yvm
GG2Ich8D3SVjDZ7DaKBe8WFBrzJJgZYjiNYfLSW7281igWE1Vag/RRybSkEYBeLinzEPVLQYRZlE
gBoDu2qM5ELVFPgZUsu8wwBjMX52/gDAOesaeUzRCoIyoJEUIdT/VU2fwL4nfNOkjgVWA4U4A2DW
1P5W+AvcAKVkFzB6VpFEl9MEiVuPhQWpkWMxpjAWmU/mNrKlIuZ4shU942TCnrbwG8IRqTYf2oKb
ZUwhKhrIK7rzHsy/uX6VEXSszaVSsLChuJXFuZ3RROaSX25l0IZKkvK2t5KR0lQjFDZ0gIyA18ww
WxpRY/tkZQbRsXvH8V5XGxt2HHklKhN1VT+u0kXqRbMtmhajMniDNWheltpZD4r/fQzsLQSNbCjn
dcVRr/bz9znZI1hVPh8Y2Cim8rWM78Tz3QuHYd82LEhrJ4CPhdMD1fY9RtOjcgMyQzT7uYD74kRk
NnP92HXHrUzADlScHN4+RC0s8CEHiY+t2/691k5O63Ulg1u1gN3pMXiWRZLLrCXKMtCKCWUR8iUB
IKpe20Y87Ob343McjaOF0C7tEB2iA/YivoNH5tm6liUczb0ZJTwvk+NYkc7b17aMf4YNwqHIgg16
o+oNRuQXZvdSvPUKnRcl3DlkRC5qdLEN1rknj4LrXoMymtDnqLsDw4C+DHz2+6N43W8pc3wPYzDx
qIQEitjw8Z2xqsERVxY2gDINe3rsp0vZrfHrF9LKroxrgmwb9RXblDbjappOdKFXXGTq4NPKHN6X
hjs6kSGRMqKP+EVcCJNmZu5R3TftZ8EXCDdYPxvZ1lT7bJDx1dR+L/R8yzWD3FGFBLikAO86XO1S
NfC99UwIydFRqrFpYxkxr6uOI2V5bFs1rK+C55P90af3je+JrDj8dwk0RkGLQaLDZqi8gbnH7lt0
v+NpKyAnlL/hN3zx68N/Z7QLcDFyi4CCCvHSOx0CBZN5g+VjF54w+HvwIFn2/qLwUFHTU3OUv7aL
xl+rmSfzeZ4mh6tECJ10zIxe3gxfWPbUtUd6+Dl+4CLcsYYetQ3lOSanlgqIvR+EZSA+9VSH0aHI
xOp0GeyBUiLK8TDjxGaz4Xi9iZjQ1VlaWGVHPQZsfbz253irmsYm5XG1YzBL9TjNElJ0MOvCxPfg
831u1RoDFA88WJE06P98kuJWSCavjIixDXELn6FRWfDrpDfjbf7RQcA/xN5hh/Gl9zyqNhJ3AHZe
9PB8kv6x/W2rm7u8/Vn0DJ4PFDB6JYYxb8sgCb99m51FQdlorga1paSrK63Yt6PdFKem/3FZBU/x
LPNk1+2ohH5LLjSPdV2y22TlPQt4VRLJI1Uimje6Lzn3m4jsG7gahA0JY/vt6ERz9YcLm1qJIolQ
E/zggrGX3p4IMxAE55BhBLzzcVlbxB0BfJb9MC1+Xb1xr9CbEksoWOYo72uoyGuUlqwuCIp1QLbo
9TBLhuhyzRF4l5kiUhI/wYnr8hJnstIdqVdUC735JT7Baz5jZf9txFMdZSjDehjJh4ZN3Ftwnw6k
jvblOcGHvEEnN/ithq214Iv4UYP60f5dpm2u76mEJecbiWpX1GFJywlkvLAV/Wy37KfC0Gu3hoSM
HdLIyajYRcJe3rmITKFF8jzN+0yNoObK8K08YtaOe4P5GkBZa7dJMmTPAL54fJerECDKZGeG3vai
fwTyK/qN+uB15b07wv+O9UBFudVAPnNOdR3SvsO+sEWBHoTNeoNAvew6wy9/79CxeLTpzKWEkUVF
QYqbyTBcTSayJhuYAhZmraeiHG4YZOjRKtxC7D4rqGOOxiILvm5AysKwCMzHgMG1nun4SW71FIgx
IjvyI8VCXhPGGNtQmpfEVFNtK5CRaPH/uBNUh0UzpvNIB/1Xs67KDAedtatRAx02yl6zwq3wC44J
hTmEfr0wgWt5iEOaAFId+7a+/B9aO4gf0dgwlXoI6nR6/qYBodqdemLAxM5gcqMhu/lqBVDmKFI+
QE7koirxPgyBaeQLsE5d5kFCb38o8ageilDyUZYHh4rpJqLeJFOLXKNPii6Z6CIEEUeGJrtH32Df
hkhwVMWnY/9MXcVjf9/bQjqoEXJpI+OiMs7awkNcnVBcXY4mD7NTH4sbXOMDOhwkE4gqAg+ulJlp
pXXzVlovmwUV8mIsveDY6d+m9rPuU9tyRfGQcmazGqljn6Z+HXwjyqj9/ieAm54N24jdLhcBzIRy
tme+S4PMEu+JuL5F2jzBKNZ3UY78CyXN5zJS6jJ8GtRyy+c0Lvp+Ju0/+DqQ0miiwrX9wbtW9BLB
AGl0aL/sLczM8FQODHHWmlDi+CEaULupxCODu4hniei4nCMKzk0xIbHHMX/dA5v9dpM8tmvZ6Ea4
Ja0/9aUz/ILqj+CGOHsIHTiFoeWc+rpSCmNXW85zFiKkitxuQg5M+eErywpSXUgSUj1NRIOLBNRV
RP/Nape9WBCcnOfYbB7cX9VzI7QmY6BJgV/vl3xB0cfbHEWr5LKfJAw8RaZpVOlleeWLytYBMAyT
uCg0zCHQpnsb4KBA5d0fuKyo3AFEVP+mKz/J+l4fefGBz9XHqXobTJaFJ3Oi5TLKPGA57TKujM9d
YJbF/E/N20Um3SkyuHqdVqas3VfBrBFFtjLgalVe1zjFsVnIHKrPd9Z4Y3+nGI+2krAeuts2EZYS
a2q71IdKkLxOoepOmYEe+9/maJz+GgRdxJ8bKapmPrmQNJ9bWMY6RRZpdLl0yVQNbO986y65dkYN
4qzsk6S6BN21LuNtywyqR/aMO3FWBe4kQUJpvq0opwh91CQ689O6LWkMPjDUCRfZQErHFJCa5/jf
ItZR1USdazi1Cf4ze3X2h7d2YHfSYHTaFI3waZ0JsiOB7M3MBE3IUqatIjGj/nIl54ENlZqNWLze
gLideDJJ/VJAc89ku6z9GZG2zU7zbTsCGy3Lhq+r7cD4AU5g/LEzT3pE407X+0I7Rwi2yoPzd/3Y
Wyg6W3qt9kvwjQvcWyvpoJacmkp7UeRfrx39nc1LAFz0iZO11Ht4JfUnjoYJJmii2LtSz391EcfM
rsGEOvYhIjX0o9fYrHzQ6Mw4dH9dmxOjot6cO7gzbcQUcBwzVuFvPvo61+ZrNifOIWcRI5Ug6QKV
3LyTtyrReudN6Z+04sJgercP6WrJPtbHxz/MSqvWFi0kMElPQ1MDIb3wdPRw//bEt1jW9e9BKc4Z
wMNtLEIdwyz2jgOKX+ZGAUeWqqnByxCKDU8h4B7K4IBOnR1OS07YyvfAgGYDjmUFvSQuobTF+yFE
Nq35MUYQgBSED5NE4BRv2OxMIq3SCtLaqREmwhhvidFgee22LoHFshLzDTHMphd7CD7ttMOSZXSw
hWHWT4UexJDFzrBmzL72zRxNm4dqkq6QBzoNe/eQ5qOPHcwDo4hwP8ReFePce+OdepgbneXx2Dz9
oxKrJukx5RXu6AuOvT1AsCqJoSquenXfWFn55miuCl/KhmFcNLnvd5aQ+Sc0zLCCQX/m2j6bz50N
eyT3yrZ3XdCA2QJ+CjeNxq0/RAW802CWAG1Ss5ZPjkPrig3Dv3e2xFb/npl3Oi+nMjawyTfSp9HU
Si7XYrBl1letKm34nCXh2CnkcDDkxrNZPAHHfE4vWSv1hhcrf8Jiunulcr7A0KkpwoXJSi/XKt+h
yOj78X2roZjJT+Ex34znOVCUFprGWYMpmiQgNSV2iGakDjWdp4Cd7CR98L7R5qiq5Dp3qD34vuV5
9XyFSe8yFonrvbgLVlSxespYNWwJmsJT7j5eJRSfwbgtuxWVxBnCYQtJj5GQggku33O2XJojXebY
inhNLb4QpT/kXro64Koh3OfZWFS1ok+WpWFFWHVSmmM2tIoZm4RMqyn5JSsTnGZCEKzUAEdsj4AK
hskHgK+UhQB9gvolSjeLe+FkB3VMIHywqAZJqhbBd8w/0LvLacknZ933gEehREqgBZloSC/DBAUs
+Gf6LO43BqE2xhvE+gbIZeOJIpX6730iA16+Lj1erWyg3XXUzHiPHMWds75YUcgBG3zDClfUvH8q
vQ3J7cr8t6qVPxgjYSjt8zyWAgGBlDl7Qpx4zpg5poVtlIPrRRh9871lEQwz7iu/TNOwxPhD7Ais
kFVr0M6qe5zHdbWmnz6vKjqgWtWQWgmq3BqNJtS0WfyElyu8GchX2vUSmdVuYYcKtIi0sGIIIMKa
2MB8NyVcuTd5iUUPv2171TZJrakdMiVxYMZCr467zFJ4MXe61UF8qVEAWi2j6NTTsKAgKN4Ov3Zp
fYA/p0psKoPkJnJeLKRflKbdwfD+aNEByH9VUQobNYDmSW24tJYMVt+Nitt/AJ285boT1m7JCzH6
CuEhsGBcvDXeM+oYJc2vgIpGLRbNw2coOGA5qgwtbd8AR6M17crGhR2riURM1na9O8hKCccM2pBd
9I4yMg2omM/sXBupO50gvI+EN20YNc2wsbT+Jh4il5mAbPUME8GR/9+E1RzM9UfLeePPGhMKDMlJ
dO3zxD3wiO+a82AVZ5ellr/jbU77YCuCnOMEYqjAtrX/XkuUKAW2bZEcHMaroyrVu+ztPB9kjqp1
8ijkkqG/Xmx87rdarRo5zjxb76CWxmE+/PPYS5GkfLghK96OrgUQGmWC25/V97jIgYt/K5fqMfzA
cqcMxbO435SiPXQSamRLu+Isf0jkjrDKBrEAoF/AdFolg1oKzm9fC/lPADUCf80Au8RI1F8M9Odr
tls1nK/eeESi/nhaPS3WDvod0na4Hd5+sTnH+A9ccWdXLTIQqOckaEN0oCNAXqqtZvbCgrFi5eRO
a+w6l60W6wHeEPj+Mq7s4EHKFWWvyH1jA6uyGd6Z7EXNAb0UnxA4IgH6ZA8dwh5ODXsSxCFvnGmk
d1qHmUR3aGxd7HS7yuSfqdvhOnal3YogNHH06ijYaP00imfObZhX/YAbXgLe7eHC/A26vy4bSdLa
miDSd4jSnTBkwSElxuHeBKjX+PngfMBjJodCJynKiXtc7XPik+lYEuRNpX3XjZqDLjH9iRDynA3Y
v08Akwkpr3MNcS9rVFIxgTbsH//8ymEy5LpHUDetAi8Hc6dc+vcsqA+Vm1SpEMEJOgHSTS76PYpE
JWpMTMYvAZm3NRZwx1JkaNfDBwNc0srajrRMD++XxAptsm3v7bFOhLjweGHY+wLZehRzSTr5I9R1
46zD5QFyKhOpEpgIoprrzK4TYmlfYQMvZlo/iwFRAHwa0nV3QRlzR1RNwItH8PnBHwkNZvXMsKwH
bmhKBcpRn2ksCvkNBMH684Ty4UD2L+b/8mVNIjeswndib6oTQOwWACjGnmEfu1u3A5rIvm/eTKFt
rjJCtGyCXhvVXaPy70ukzLD5pQq/fOljD4JHkWu9LtyWLPRVdnPWf1HP0EMaMkn0e1CUihVbFKb2
NNG4p0P5Ew7S70o5+YqsPeX3r3F3rXonrIOjTjI7E3p11/1LHUG39WoBKmvcpLtWSiW/wGm3woTv
ZsNu4iCgHJhakM634jWrsMzVqm930etWh0N1/NXXj/w9kFnkiSJ266G6ys9YqTZAlmeP0Z6+90Ot
EtlVc88AoejdF++ZYgGG4Hr0X7I9/50tX8cL2K0sXB7VYsG1VBdRGiqo+DlJns+e/vb/hZ8pOw/Y
TJcDsFKiOpOSmMEi56tu3NHImgeAXpAISOxheq7xpdRXWENkTiDAcz0M/qYwu+7Whg9rGywA4Ch1
IR3T6zz47loo81Go2ynqeUhg4bF9yOxKBc4/8zp3AJ0x3GEgEWX9a2udxV8r4vMEEqMP8wot0fvu
oB0WWleuzvSmb3PaFmLS5tI8vUXQFpppZjOTEoL4NUv9YB/5dKmCRHNNWWvyl2D5DxvokRAdW7wj
cqYHM2NM/PXc3drthRNsyPI6L9gAVGQ7igGRtsDZyVWK/09rHWnAvd0dQSBJlP0LDGQFCZlBHKOs
t/TKC5zWveNDfqOS2PNxLc9NaBZ6qXhw174Zk0KKSbB6IkE7sVxdNdjLKQI5T4S0gFHjUL/KIcCV
Y3KTZiLy9nxgNMdxSe1AagGVsFrV0uP0AXgCXH2+wDaqO1rGVjN/IdycPQpHtv1ssBx+XskH507s
2UPp8Rnk9VsTOp5MyI+sAsdbxV1x4XpGQQy3vTxAQEi2puUqjFyZU/q7e236tXSi63qtG4+TCDcy
ERLjjp+ZHi2BgB/lGQNRY1lN0uHUrvc7Malb9l5DPTokl5P7bpG6otfE1HmvZhKP4M+VJ/G+g2LA
+bxL7RRpb5kZXLeRq7PgoAENtetg/yELIoqYxgP0z8z8jpjL+UrmNphZP4mk9rqI9TShMUCj+XuE
aJkW0LPwqDumfE8IdVgEjSFCBwCPg8gTsm2dRyQbw62ivdm36P9xUa0MDpxTyw+HDvxJZyhOLCUB
nyyH1RASi+vPnY6VVn7RngjGOBFXci5xJuEHDCBcgddPPOhYMUWl8tOdt2ZdWiKHjr3HxOmpbzCC
TPrWmImJDcQmJKR38nH8Q9dv1ZBq6+Zno/fkqerLWrFqqSI4FUVwQjsJvAPW/HB6nCvpgzSN9t1x
CgHX0FFbdcu353sClOath76WDp/tjQWICMZe+uxdA5MzCOIhkLNkqSLQraymvtQO0u6xyVlFVd5y
s+nSbaLN1W/hCTpPpRy4R+tTOpvc6Fcvlrm7NEUibyHsIcKDNnlsbDFBGcam1djfvW2lQmr8IaTp
A1XxKiFcMH8C6f/BbT82suG9QYKdzCv+h2X5dqjqZOSoTtYolXRWPzrIFLCkE7ff+oMKPoRZ83gD
qmyT6+V21xmR5aqVWj46WRUyMbq9gq0MV1ezQ6gyJ5v0wT2n1zgcKnWzjJX5RcyJnspCTFOzpBE1
d8JFVz0GhsPfR0j75+iAmPg8/2XhYeqwZvd95fmQ73KOCpmgjQVQmSHvxg79TMKJOTmdy5LSShXL
hYOiSeeDN5Y7T858JYQadTQSmCvKvNMvghhPZ5zIq6D8COfOP07TJVQt4yvNP9ShkPt3/YPouEe7
2r9a5C7HRijYFi35+mPLJ26e2YvZawECW++3tOaBYS0coBRJl2Q0Kq0jQLyZ+6tiHsPMnO0gALdq
qW3LekhJUIuS8J3EaYsqpSEOR9BPQb2KsyHAvBRGgnB7JWg2qdUWyi4gK3Ntgz4FMKgvW2LzYyiG
tLbnbpsIkzUbDduAPMkKT0+Wfqx/OMwx6EgNr2xTPMj8WWwFw1diP3++6Lo84YRNIHyU7wSPsey7
1qVw+zpGb2J2rZVEgZQrusXJ6vJZhmnr6DnmGvMFJKxweliXwSVdT5HD7vOoGiWqAmRADp1zBosd
JuMEcyITFTp+kOgyQajGBTgPQU4N9hmlXyiDvTlFD5ge0mc1+Ig1yiaOiXRdVKvUwmdTEjwCebIe
iWbt0Gap6MGISCBlH/dDZTq6k7QkXqKxiAYYfgkhrh1QHs1AOcnbgvMhoLeZFW2cRkbhHCa2qmpe
m8Wn9hjXYY5OgSMCrA8V9bqyIGbY1ScaPr9awn5xw2wpRWgQ8d1iBb+dh7W9TVxAyYNZ78Q8KI7D
1ZoawrkS0ftUPIRBQd++WuiefvMUQyjAtaitb3ZgcUkzD3eU+s6wezSpGc+60hOmoLma5rhtvO7L
nDZ7398MvcLeO6rlUcqUki8GbOZJPoVWpkFe8OgxcGv1szOxqdeWx1DZc+98X1wExjQzYJwD6TSU
Yd4WYKhTFek40lQI+7ySk+zdUqXgVOs9TT3rhsEDaqzSFDYXwW3ezmvX4BWBy2KREo+mLqABw4mb
WqH9DDpqQQQ4h834X/4u5Z6+Dza3ZvHjr1rZVYUkdvWJuOuY6maylql3HJXmVMZtr9PoGaZm8mSz
xD7PU2TCPfaTapiCXNe61O8Cm+SSq9kGo5LDnhGK3GHbcX9gNJUAHGMuPhaIWxFeBBy+FnhRD1Fw
KeQl3fLoGUPP+Nh/RnSYNpO6kzqSrSXHiXxb1hLXf6AwVJrPhF6c0nB/hyDbGch0UMlzboo+P81p
2fsrLAI3A7up2oM4pkCbmgSvKW/X2Z+LdAA/e2vloGMuKS5JnuVekvj4CnVa5cn+M0p2dxyn9bAt
s1/0emecDNdSLi5zfn4XSEyoodMJyO4BpY4de06s272w+0prbPRpRePx7e4c3LF3ZrR4/TnfeNgi
kgpV5wHDeR5+nVDkiRVSgn7UII28BQcbFbbJbvq5zWt1PwTop4gh4am3Z8nPYzcYc9377q/YHErQ
SG0MpKmb3vNPcu3RddEmgFnWZbAEakgEXJ3kvZUk9jLHgARApzFRjy7qoG69ScXLqmw8buiksDzK
yNxFENi1gMSrplyfe6qp3rv8CLZ4jadNcmOtEf4C1ZniQjX3Ax0nP8GbPFQo6m4Kb09J8f48/pd2
1s2i/eTfSPVKE3yPVqpFZfJJpIv3sVp4APIKmK1eckCJFqJVyTu718i7aL69Hiw8RBjawOymkUY/
W0xLjM5/T615+YTXeTVpnLm4XJwYnP0fyJB2OVF7FEnLR9TbEULQnM5Q0frISodHNPvLNqXY4Ywk
33k5tbqsSVwqJ2ApBwxkqN2CW0c1kk2lzZPBS4qVr00/tMJnq2IcxeyALiFKxfqf6QTIS99wRiGm
+UQo1mLygn/D0DTdVnu7lFclnvb7lSWwdSYFYVI//raiuRwvptWWx7Adz1840mZux4bMjnXkYs34
rymSb5c+y44u6vJMV3bEU8eqhypTXQNdG04Myrj5u/TSkVavHOt9NcdJt8sngNW9q602dGeSZdiG
g8rwHhvVear6N+ctJes5h07ONqe04G+jlgCEEyVWX26DXc2GDipsn2eLGhkZZDq+EqeMnWa+ovxK
KigdmPHhFRAcSwB+/dRisjArU+bkCidBsZGrWrw665mPZcO8YJjx4+JHWK11rJznJiRHnd78QjMH
cdoMo5oc0zHa6Yvh8bQGT39MEjExmJBZOTzYC0pZcunXOHpMCD8GUB7ihb8i1rI6s+TiEas9+nz6
nrxghfFfHDt18AMZCj290BaaALhndj3d4f/JL2dKNOZksfqDnn6UnKZWRZxbLUXkR7/Oc3bvFt1F
4wNCCNEE3EfOUSi94J0VmTJ8jPoMP77wsGtO8fTwIZmNRayQC5tv5dUBwOIyhDU4BL0kmFEhcaOR
hUcu7GsUGMOvr/XNBn1VceQKoXqhIhBRCYb5ME947YckkZVhYe2qHjRM8HSK3NRFGuQY6fsrscx3
h8gN6uNKfiZJKaMFm33IlMkhuu+DIshPc8N7jk5NSlGvvRNYKCzF5oTnze24JbnaJfSJqDcKz5vk
8YylkcDGAli2tOCFB6+b27zQ9zBKVuN47lV3aTltb9VKkZ7dA7eycqssRs8gW3DScF43pjrxn/Ej
u0IL1j4DIosSBvKPcZR30HEJq2PMMlSd2IeE84uMKrHJ8wUFJPhYAvLXlNgoDj97obhhDLOfcKA0
8zFsZOH+IGFHiWzbj3JQ2MFwDzmjBC3HD04s7vdwuY3Ps6roVre+CJMGEks7/qiPJTjtYcADBSRk
1om5PGnh2vfNbxbLMdG02cqZoSR2/OkjtcjUs671MA3CYqf0gtzWYNtG7fNTF6hZQ3AKxVhnn4/q
1oPEk3ItAZD5hUmEmaPGEYX8hC20prYeB3gi1yvFERQOrpppeckPYPWdQEumjYSJY0+ULJkhCh/f
ri1XBEsNILws21j0SrV3bL+yMErD5SCmkxNgL4fV/5zvxLyAkGUqPI2k+ZuQBVHl8SCVo/FYbRo+
0UaKzp0HpK151whUHy+JQOYAd3MD+nZ3c3H6bQBfCLpRkzKYmzQd1i3oqAUVo8XOK5C2RiQs0Dgi
Yz9CWh6iVyHXtKMiYPp9KcoHuOwqce3TMLv62+t6arRNjXXdjiIuYG73wn6Z8S0Sf4SJNLBequka
pOYw6C47ZOlmyFRDvADUKnX2xkppoO4TnWLN+nM1qBuscjXJH22x0UqJaSEFIjAigo0IGxmJac83
0nifi9pzmcvcEZsmLNF2n2dcktO/KXwCtPy1YUO59jPSy88EMXk/XaB7DJ6R4k/CWW1NwJykskkK
qWKsYrqCUZ5qCTFQelNtZsWQDbnFu3xUJHJn+mcbT5qW2C682vCRuqOkQn2mT25LZutVRXgaFd7X
JNbnsJjl551sxNYDu929f7F+uMhjsbdaWrKv/6RebXXdvh7GWfXk4KD/Yf2gFXDNaAzhqCZxYnWM
3j8V5QiT2ZfCchfIvM1a+LJG9lNoyoTXtHLvHDcH1u9oknYbPZP0Frm91NfMCH6Jyya1y93TvQF/
7sfzwVTMdrppjw3tA+wNiaW50x7HQxpoKLrZss9K59hBF2MgUQuxxiOqHQghVa/cxlVeoShMr/rb
AbP316nhRaxhXLC72o3rcEzG8nxIKOZLYe6EXNXabKsS73luXvglUIHdRNJCwWV1S/gktjfhC/88
b3tzQiEurp5u3KVXfh8KgH0BnwA2y/kMo9F9Z0id0ggMYuSLy3RIDbNcDhbSd+KAj+E1Es27JdRy
N6GCD4JZLlsY29EgQI7RQslyjjdbKi1BITWugtB58aLWuhD/gQiOlPmJuvZnXom6HQCSTRIRpHFs
uWRnUNX9PKDJQKKjOWJ76CES7vQHAvhYsSj31EWPVf17jP5j1Zp+bcFhhQWrxDUVLq2NvSTyFaYg
NlGBMhjykEdg9a9lTuiD/C+lRb0z7JpyhO1sKMVVUQ9PEL3OeVcgkNAqQxUpL/BBT1dq+EO6SlNj
Thvhr8ceoc7pNg5lzW0xamkzEfU59mfxs8jWOatmqEj5R5re1G+i1o16ybDiBJj0C7oNJAh4iW3Z
kuSrIrJygZIgB9DtDUWdjovy9n1RPgLuGj625neSCmRFD/+PsHnxqmf4R8Op8mNbIfxTNtYRKhTH
MxY9PBe3O96MHgF1MlTZ0lHHOMQ8N1F8yzGL7NzFTXQED5SO2dO3cPZDqO6jQHBUWyLnQ7m/n9gC
pABEqDTG6+92MAOWcKpgWgM0Zqv5r+zwc8aPvNBpH6l3FLLgRfu1PvUCkYJhHG+iFVgCclNhXW12
u6McBLkU2Aw3PyeoUvMMC+apgtkOQ/tHEYex4EoTDYcoS2hYGxFmTagtvyDLi3yA9xL2lQ/ngV4K
fYaLk5ua5oFoL03W7HexTIJtNvQ1D1VCuT5IEWd9QOemLX4VTD20APGDoyWVtliXqWXNz6K4Wo5O
6ncrBcMB+3hGsHEIYhjmiAtdy3sI60mnxw4R3GEjevuYFq9B8JMu7m4+ocdSvXYzP+GV59qpyvpx
bRyDEWylj+VJDPQGh9zReUVgUt8GNBADYsW2tYGbA09/VF6/Hw6Owc/2eaQqtFRSLKJB2F1558ZQ
LwQbb8cZ3//N3HOta2d7/rvceE6jh3aHGpC3+wIrOrk7crbMLox/3reqPurk19E0MRDbv24zbAD4
pWUEGpVormlm3wk7xwdJ88B1GFdmqkvd9vUSUwXUo5i0MvACqPOXiDBS4cgB1h5ozYVz86tl5Z5L
j6cn8WEEmQUFeQCKBcUDE/fsyhBGkhq+1Ub1g+0/TQe401SwS28oUb6ErYnBHu9Gnz3YH9GEZBRR
7LMPAXNYFu4+Wk6l7SXV4vjjJmyvnlLpJR2Kz2bzXyzjv0jej0kcgw2l50QYaUhGtCaQoZkr2Ojs
zLRhlujhBaj/poRcC1ayLFhQHt1ZpQEQNASpbaugp3dfKRKHFv8KaHLcPfIoUgiFvUN3CJGTelw6
esImHptizp65rcEDO21Kv5KjUoxrkCkWUiBffRQYspsNxNHXaUGS9DszlpNLllOuw7HMFK6FQsdw
tXxyhpvloaH30pEnkMwzSvuatO9cW6NZnpftf+pZ9dFet3x3GHaUP0vNqKBhmgWED6fxU3d1tNR1
utIvl3vCsJ3/H5weqfPcII65wAetp9siPWvBswv91Ii8mbnae7izzMYtdMbMzbgaRAxkijHIHBF1
3OOqIqlYOfCkD5rYwyUFQALPGvTbNg13F1pGJ9heIwB4gLfGstJZ5EKSlkCUIekjBbkZGXfUjhtf
zbuqbvqBUvi0asRIWvpTegLkiNVGwXz9PI6ye8AZEcf+zJiErcCPzZPmtYWR75Kp7wTo2guJ3bFQ
AHmXvZ+CylQJjXhBR+XYlcWUT0eaTIizHb901i6XEOMVlcCXTS1PHXcLw3YUQvkEuc/nTHancS9x
liVZOHBGPmL5OoWiMDQUAbbJfMOa0f+y2YBAQ7J95tcS8xSe6xb/WY0L6gMQqQ3DSLFku4pO9A1m
3v6wb818Gs+uG0QOSVnvSEdDOdIGLuN+TkCx1JNa4j8k78i5qkUxBFZr8jMMGtPx5mWS+RhhqV5W
nsKt3khlw30MEnCbyqrwX1CH4tKjJrM4oP4Wj9pnurKC5xN+rh8Y9Q57qIaGD/aKXq/NukqS7cqW
VPVctSsQxfmv46F30UA/7S3seQ8LU/Mkjoe5K+m3QW9+TktCrbmrj+Gu/fCYdo4WBtRBTqySb01+
12vMZVKzHi277KYWT9dqBzsF9BuIkCLYFe4+BbrvdZ0z7f6xm+uULO2umoqmzk9lMJKfA3hRHePL
JAbDhM9QJvk2BqQtEJVu+1dTbDBa0tTNSeQ8rgDreopA5tt5mDrQ1AXbJG16qpVXbaZUYnPD0eaV
hPiWepcDEirSJZ1vAD7OFVmit1ZCmkehvL4ph2+d7wyOihGpONLMn7fHApWksfcxT0D4bcef7CZe
JdmYibgCDSDM5HVJw1u07G8hyVZNAR3mJs98ZGIZOQCDAgHKAbv33mcAcyTTX3sJqhNwqDOZGO9C
v5erJJnM3Y6eUynoc2S7Yq2DSUY2HujmI+uWT7XgqtUXmnZBU6cMk0vOIqb1EOb23s0xHsnLGE2+
Lz42nMyU/nvbdBRG3hiPIsLOhk3214xOa5hwsyhkTCXGQHo/rCVabCqrGONgxn7FZWddtu8JNUpm
HIzQRg/AwFsESJ0rIXZzcUcsCRHxyRpe4F45BI2qjOnXX7flv3JoP2QD5DCqmB7nst0GqF/wzzBM
JSFl9vusFfRcHGIhN1VjzLEdzCsLQ/4Sod4DEJqYo1KW4ALQh1r9z9ABKSN6ItnUJT/HnjcKnTcr
8Hy/wO/eJZ60hsSsPjef9lvxxTkpnv1R0RPs128XxOT2l1O6sinrTw4oVhGHs/JM10ieCSV9Vk1T
f5We9nILHYT4FnAIVBuMzxA2NQiy9V9NFhpBA73PLeULt/3ui9loXBj91Mp+OnxYcSGTP1AcCwYw
H0CSLLCGUNgQ56qMOtexAlx+s7JwnMWZwOcJDTucvTLsd5mCbMYl/3dMIGveQCBycZPEKQJbhtAb
hEJvTdLl5XriyB2Wk2v9qLDj9odAIsyAzTASIlWtLJfHA09cBBSoz3+dMP27gdsH56C0j3U1N7az
HwtnTzLnUqCZn+7FUFF1P5WWIqlgS4MNp6d9wktWIuo8vcBDQmX4kdZX8zDVI6ecpzv0rflNY5p8
ZaHsKzXq08Rk91GsLWue+q9xm+yko+7fnvqy1xazpqF8H+X6O4ixZT2Y3tfd95YFXHSfjIKT2jYJ
HspsQUjpOafYjJGDYaDTaxvvvE6rQZ0MD8Z1Z9FwqTGyJTpew3U/iEGYu1zFB6iJ34a2v6q38GV2
WWA2mj2sA2L1Upz+R7LUfkVNiJn8MSi5l+KOk1SXiRFnJXA3yDyDnbpXWDNFubdn4XRP/ykaZ/jT
MpO8PueHIupr+YfTesoBF3bYYJHKbh+I7fYxIVC3kVodXw14qsnhLNls3HbxWJp78q3XhAPXaynk
uIwULWX50SwdoNSOIuQcrPcuAxUlia8/XjDQIkLaWpN7dRq2NuL2bdV9ONqIU/J+ej5vmXKgrhY4
+WK01iv9tbtJZSDTai1iZgW0fKc0sTC8BcGRn+IuCD08TwLlxqyvpz4qZYSiasD4nY7sGeod3ZjJ
v2GiEA6qb4pX1GTKeYa9NC/oCW8Ctnzp0KrvyPevwJDeP7bfDNJWfMv3iJfBi4RnNQbj2y/xWBBZ
IZ6wJT+IXgpgo+zvoopX84zzMjo8L+jTkQ7jhOFJAEvWYmD1IE6weW+BSToODXzqQS/xSfRxmTLp
LIaFRhDPKyHR48O92NHuhZiCUKkoVNfukYjcFiVUDdSzXYIbPSDc9wR2ib/DJeDy+4pYL1eapItq
UC+Fzmzh3Q54DcVOo7mgTVxrFQXOhE9aMNWgQMDSFcHFikodauug5nYKRcGpt8P/2A1A1q0CBq9c
UI0AZz9zoiwXNgWdTbT9ng7Rtjb6qLc1Sha+xWVhrzrAhbNs5KnGst0VFjeQKn2VDCDYelOJ5m6G
86QwGZ4EnEyaHWHNDxCYvex81E+inQ6/3pScXxuGDBRZVilX9/6N2NtZvfvadC5RP73w8l7AR5Ma
ZalrSYpLqJf5ARKWXO1qOUeI7x6HWD09zR7g2i+VXf/2mXztxF8cE+PCwoAnvfL3STJjdwtpZCgP
KeEXYWYwirb1y0WzayyLv75tFrpyEYNZpSBCUrDwaDE4X6LkKg322e5y7TKirQKe6Ab/+G5SB1uE
EIqxEcY9Px+30ClbDi85BXXa0mQ4xq50d7bPlW8YfVFebmV/dD9mhsCrUqdErV9a5Xbz+uiS52N3
C273yBuyaKoqT2K5q3Y2wY/pL9sR6Riym5nQF1ZdJdoxf8hGQ8OWexK8YgukPaZFemmVps7EIJpH
a8Dn5iUmFRAYVMfCJEBn9i01a4qjuTvh89Xu/vWvi1jJqAd1gDWzqC9F0mgNXtHeQDaP7rwX/zKv
7gRfSvYtO0AVk77CVIRFJIfrguYto8E51qXGr/ZxH25MmG0We3w0U0KoqyxHP/N/+DACH2Li6D7T
BobG/liqzRliDDGytv4VMt9vCsynOQ3XbYfQUBKW/Iv0Ap/+S+oAJzVmHT33QSEB0lEl43fbUeLl
WOg7t+Iet0Sxch9370iz0fj0dIEhgYLReV0DcQs1iFOhvmIa7gdMnJlBjq961UC7j4Qze9m6EWpE
CnzCvZWhGb9+0G0BDf3qXFhX62oI5tsOKLUis0jSnJwJRsod009bH9k3b8XBPgSZDYn4/8fpdRXO
GS5Rzy7EgmPDdkYuyAFaTxG3ItfyxzusGoPRWOOtwcnUCJ+NiYuc8eX6eo7qk3PfOBi6/YStxqKE
ucd+1Ia0WrWgVCMtj/pXY5MqwUgloG9yN1jpeI8mv0EpZW2iisE7+uQR/dznlzxuQz6IY1+dbs5C
Md5eeHOiLDNYQHUrpV4lbBzGZdl0+No5HjljggH8y3o/wk4jN0aAjFSzM8ENJ92Cn7fDW04upt+I
5sd4w2NXf7Jg+NBrplF0jux3Z5Odep1dHwpqweA/qZNz4RGXulhu3nGpEAYnmuZZ+YdO/8yF97tU
8cHNXv2z6xR7XJ3EblnxYDX3+RPUCnT34CpV2ko4inrHUlLZM7IzEgklSDNedSGbgDilyCwTj6hl
bbaYG+JxQLPEfc0RT1MBwqKEohfVpCFNRiHTRspz/J54GCDeG/4rSTdrKHFsDny8ZGLyHZcKdhc/
ljXbMmgoguH6cREfNMKqxOaTsw+FPZmGuXEzfhSg7zVRgr9vNDuNoSrFfs+6vg7Jpwt+oE/fQO3T
aKM2DPlc382LMHkqB+pUOnuApNBbxkROGc1qVq7zir45slunfNypyXwHjzKCSe4YafY9Gc7DLe+E
i30E6aZkgmLB7To7/S9vW9VLPtIbrI0Kt6PTEbnlPHfG6iyaDBpIcSfht88nvJNVwrp24WQy0xVB
v3Am7qd0kpR7QsotyDTOGMCpcoxjQ8juNrA80cg6Ke578STSO5z5yIeCudXiGhVoV0+qAxLaxci/
n0J0KD1wWandAHKfl7+rMxWAD8SHO3WkHzByrHPoiANVDfvMTpB9h3vM2msVq9ALNxALZxUbUmh4
rksXbQSMMEO1Yo6g5W6XoIOf2VO3ZIaVJvyelAhFE2yCtJNnxvoljC3veSG5pRdqzHvUMj1cROdc
nRHkGa7bUFRgu78MjmfMJucSXOanPDw7TBknZuppIPCenLZ35MN97asrPvQpdj2zpaqEQntqyk3I
VVRSPDiToJ2L46a1HwkssAW2eROcrJ+WwV046oVF1962A42KPE43d0fGes+utHuXaeUojgpBQVf7
L6Cd55A3aRe3QFduIBTeqSoovIDuQly/U9fP39EHbzytrqotN3uS2ILc3ib8yXBdVoXekYQMLbII
wXIa5rfskjTVE7eLEiqQ1cKkDv3snOYW7EHTPmXyPZCQ0TjknwfA+W3EuMjHBGeLzbu4Kbu0e9OK
EOg4VQsqKam03ExQHQjD2gf+wPeTvmAeLtskd6HO2G0Q7MuDXVdSf/e58eDXwalHiXrOgwutp3a7
NLqkeCFpjtbqLm3wMQIk3CHXyqnYmIid9jhGlfSpG26HKMMMu/VzhETqk4gijpOxZXYRCD5ZljIi
gLE/zsCYJKQsQa0oDvZPwUexkD61R8TW0u2SM4Q9TeINDffnoKuKOMw3qZF42kNwQBZ5kkdO8Vah
zg/CKrtnfDjflKJCxYnQ25kSt0HDTOueiV8MKXsQujZpa1ru0MNErp+8hXHIYcFy35hIHZXeFYie
OyuBvNOtkqgGhOFAivLgxxQEf5LRe62K5pMVRHEHzOK8q2T106VQP9Tj4hyMYLhNx8gGcM5qYqfN
E56VDGpfexaPFQKsjUAA9yn2GxJvm6D18NunxN/PZzEZGHecEdBGOEl+Flf8LpLUfrRFHUnYmnb1
QHPHWztZJiAYaP/xMXumep+e/kZuLnFSMR++i+5PGpR26/qt6YHM9kqP5GTSOkTnM7qw4GUIPTof
2Ua1OkNIZlPMjRuBW5AoXWV75WmxQKLxjs4jSNuYb21OWoY3QQuLIHdQCSv4JyokOAM+HkkXJ3PN
+3ghA/yCGHUGRVGbNwO+95hMEES3REcOhtM886GlKwKJkwbKf/ufUCMcNfrjtKiIfXpZ08ZpUZ9b
rs2hvl/VYs9GN5JY0Jp+V9+2acb/TX7hpyyxI6zbVzKhAug5iQwpjo6YrKPGw0z/ySAph3Luwklo
PEIBT8r97lA/WVxzZW9pnIpNg5d0EMT803hz79c44L2tf1VSAV9XusHutX67ADbwu7fsjLu5Nivx
o1/BXlGZQ7Qi7RHTkCD/5iP2IHVI6Nj4DtW+ZgBIEy4fdo/6bhc4OfxZnVmc1F+2v80t2WlJh6ni
jj9jg97qJJ+qK0vdPbhJSEyT/c4b9RBhMnd4tZ18vlG4j5wXJfx2FDnQnNQeYizn6B++O/GH5NIc
QIvQu/bToQZXwGyoLPSjEHlyKMFR2Wn2LbzIxRuIuP/oZrsXh/k2Ybs8KcFmQzOVCwgoElPJ3AqM
6cv62cFpFfSBymUBYY4uq1NFLmUsEfRx74g/gwB2BHZ03DM8yCslNBhtHA5EnN7uhUeR5EoIY91S
u1F5YwS+olsiuAzy9gOMKkLaM5Dq7GN4DNrFxu4EUWQ8YVdda8Xu64NbdzZoeOjIauyWbRQqYfUS
8xdE0NmJ3TvwsCKfnF3+Dxe0sHNJ31iK9E9lW6AVQEt0iZTaBWVe6jiJTV68t9m7DJD3vYbQS3R6
aXtCrx7HtxKKD1kBzUkGLwMG3lyncTBA+L3XUbkRzrdDAX3ZVszJBQWZTVJUb9sUaKsy6JT0tYex
JS/9QO6JEA/98gbP5v/oWPWUDoWulj2UIdxJtS9QzyGhVhwR+StmfZlsaPPMjeN4gz78Mi5eP3NC
Y0B7HcNru47SDSmLXFB9T0+rP33g1H9cvPFh4ddSbDlvOTGnvuCmRpdlna1ZVzwLbx/AznhjdrET
IrH2pHLYQiJt3fbPv6ZNh++PF3zJYWmaJAJr/pymHzszmk1GQvn5YuGjB9wPjPmkjAZczfy//ZoD
1WsQJh8w5C3jwlSYGKGKS7iU+Iu9gToAQavN48uZ/AUGw1D5XUkKYxt8kGMtXbfMeVdeVmHQ2ckU
kuMVHJKTK9vsmxmW0Z1ecRg1AB6AV8q1JP45RldhQEWhUrb2sYgbsNNJ8NK/979KDUZLONMBS8Ia
Dp3gXqY3NHWhmr9bssYgLYv0/sGoKOVER17i1ZiTyjszCbC/yKOpDmSc9XJnEXDpG3w6e6mWVntm
CE+VrXT9dv06DL3BXSlySrNly14Hkb0hEDHc7dm5fITqvkCcmUwgMYDw+6LDecvHJEeeekBMdLZJ
bR1egdUqMgJhVOB9zRCcf6/sPVrm63btEtWRz1fz36SHUhNGnPx7gisjDIwELK3VsAo0sEMB9xXs
MmXNbBVjWnxn+a9GHH0XoGVGvf92BH8b4Qq9IS/G9dCVtWGdEQTm9VReZgWRtCpATp1xfPlnR9re
4Ya1DK8Qas0roMaLzlBsvN4zo0vrz78o19qgcrYzoWhbt9kvduarZgDITqIRMSPffXQg0vU5Ifm3
dD7Fm1yA9YHP9ref5yxgan2Y9Eoo5vNhkh4pkvoimTR2uZTlpOwLFPyNqOuuKdqzT+Z1hXMvjAO6
+Tuh1yD3IVW1jw+BDbTlpXrqpz13afQMTavKP1Yej7ffnAqKOrpVeK8T1WtOVfiCbMV1OpV6MJ2i
GWUs2rnWEp8XAfeXWeOYwlEJujymFrvPfCI4PV7r+pjFNGLWfSDXhK12GenBVoy2SOCmU4vvldDZ
CsBZen2zwWDgnPNhlgbZsHeBfJcpv6BtrLTVh6Is1FJFxV4h8jynWFhZ/Fyw1m9kGvx0gbr7i+tB
QO9GsKF4KfGtvQG8DIGhoLMSyCxhsMNAq1PRZKCbwwkPHuWlx0VtEz9yyXBPFhT0MQCCxl6ry9sl
eqCPiu9KoycIyVc1r4Y/a9G9hExeOVoWD61TQFfxf9aTqSyIRVtJ0M4QPquuuITrlftH7N7p79q2
ZJAuQC2s4uOLuwHzrHSvVhOIhAWwAgod3PHqyixZSoswjUlM1OoVUfTZUeg7jpZsXoyDZLe0dSOA
ql9OYFlmbcxizFv90fmA1llpoQQHtjse9GYPJDMGroNJTGseU7zPU5upq7IPWSVwlrxW99kvlxG7
Q7wLClrisPNRsNRtLmzr+pXiLu2xvsjtsXKMX38RgxN7H9Fl5POPUOsUorQtdYvbDHy1C7ACvrTy
GoHBW3ch7Ax6iC4BBFe+mc7qSl4JQnCybn9y9NCSpBUeQ4ySMogbgrpoZ14la7M4/pL3hFkZtoMF
NMvcCaF0oYLxGkfT+a/RW+T5hHXbdiYguoQDShfvB+87u4WF3b4AW/lUCAJmQQZ2VAPuzvcaZWQg
gZwDfvzcySEknxNEox3ZWlmL2DukTSe9MhZFB8pwq1BzPzd/+JUPxa1NS+E5jEeWnbYMke4qbm+H
UQieQbF3lc3jEGZ9OWv/YKchSERLV9iQcIbrQeTKVigTBw0w6NJKvCdvMlgCIxdQHl6/Ncc/GXLH
Yun/99AA23YdmEWUSNQ+DP9yAX79yw5LZcxh1uoPXWPBrQJ//k6W0jvqPK2sS4VTk/wAnRSJC5RR
Fj/Afrjcg0kJSxzIwqOSjsQwsn0yR9kIN8nsQRQks26rPhUut6VVqR9RccU//8fi+vc5yZAaeR4L
32PTL3QUCdHN1xMXHkTE3rgyaQhx1Ew1k54TMaARDbUrJwxx6ejM5ic56vfIdziS8Cft7iRDPXyR
8nbP027iEQV54Xr+C4kQO7fTFX+Jfm8sZrhjIiKTfBuZFg3JRKTA+dDHA12zZt0Z14KM3AOoNYAg
a0aYBIqypwfU+j1oay7RoatCxbfxBwk7/JfR4Oofcb82Ijosgftsx5Vf5IK1fAGgucT+OQTAwhLC
XtLM2Y/TikoO9XtrFDADgY169n6NY+jlupGwgZnVGLmY1ln9pNCKL2DT39swryvq3b1W5E/Ks2yQ
8HyYoSt5yJfTFfgGAquU8QPGDXA6lQrzqId2/y1Qz/l++2zIvfq5gGnJW9oXps+KqxSSOiZjHWAy
JAXjcGdLQ4eoSqi0gcmVDZLZnMhLOsMzDzqa83woSecPSrspmFp2/vSWV2GmJyELN6KNpIiC/4xP
Qss+4A8Jn7Q68TjJIy312vzR3d26H6HIMkZolsbd4eT1G1QaMUknB6kcH8XbaWA+2MwkhMqonyaw
lQHA2uDN6mMMRqcLCeN39juZ6BwMk1Wu8rXmw4fwEZ7TIFPsRDoTK+Sa9Vp7dkYzUOnUS7HRGtWo
/wEcV5rpGdnhxD9Syf91mDWtW8XUM79jGsd8+cO+T50GCA1+bkRDBnuEsX9jUjvmbdVENhulYFIm
wcBM8qdfxYOJIfOvIm9NdJzfTRB/bjPQI8jBBOtGEhrSltoXSR+DLa8ic6mkvaDApNjBZHpye0FL
CJ2LceRe/teRdcpUHE6G0gwMdAPqHTdPXWqsZCHwdcB3vLnQKe1Y+pLLJnFcixUg4dJ8+9bKm7GR
J0KMeFz8UzSd3nLUr4XXz5uu+Eevg2gdUOohh6hzW4sHBkdkw3NwTIck3KiA09ehmK8zoSo/c8TG
Y+DLpW45bcI0CNFEBzyAyk6Pac8dNTN7w2MT32jmtZUd4o7ZZu7aYS5ZCLIWtORa6MX3SxV1OnPA
1LqprYKfMn0/apVw6p1ZYkENMx3/5OJlyj3zubybvqNgJmw3RoHGNI/niaa28bCINg6reOzIzN+o
Q8sIouo+oXgGQVw2+uKUf3r9PjllpS5h5L9boSc5zzhnvyxN4wmyGcxR4Yrxm1kyp1E2ebs2x2Ld
aTTxqUYVCY9mBM7HswHO11qbWaOcHPxEQJrayazUYmGG8QdjE9dg+PuRYa9NaPwKewOSHv4crM9W
FtaqLrr4/E8QV2atFcQ57+6MwkVhz173E/hX0dRPLtJ2LuM7Uory5crX6B0u6dxt3ZUG9EjgAGcO
a9EdlGMSG6WpBWnEiGxvK8V8TypakX3iojwiM1CEfjI8a/WqFWDg+Cicl0sN0Nvfjc5WgR7HnxDu
ZFnoFobwQ4umKz1W2rqwbBUa5AW0s9al/SligUCdQTMJ6mPtrOHUUqLtrJvErZAOOAtxdc2INfom
cJEapZJ0db3wFKAQbXbS0X5Q+7StXv+f7OxWkSmYxJb0CUd3WdeWLBDUzI8RW7suNBxDAjklpTfP
9viqVhTnWKPuFpgsvHowAUbfEIUKsu3h+wAH+KRaccXJv3Pp/Ym15TS6L78sD2WudpK7UzjwaA+0
IuInpH/65TI6t3r/b9mHLVQMOR2QBiThopBEBK+aRaEJtqKOpRksXJXM7k8laRNZibqEB9LdDVix
dfzykNhtNREIb/Y1eh0X7RQezgaz+d0BJwfqz19ZoTmcYHb/x3B5qsnWaWkKNmtW4nU88lcSegIJ
YmSnMSP/BmZ5FMyOQh3zZ8F3+qGLW54FBQSSFA4iSnaxK0gqTegmnB49CdLdc7hXeHzSIpwGpieW
1LEt9oe7+vQ5L3H4VslgGW2Lr+zvJFcxT9LbX+qz4VypFMZYhtw3sEpyBeKF6hM4ixPTX/Ix1V0E
B8k1kfvczsmqZrLdzRtu/NSle84J2s30TMEXm/wy3HobXMf8Il1dSn4t4SKzAtrPClyBtCUFSqtr
O2dbA3zuZ3TXy0llw+m9S0453iexZFqMWvKLLueq84+HY+fVzWQTq9+QnFVhbjg9NPDCmvxbwLhT
+3OZvK6dOuN++idbbdqBXmC952y8byVoBAU3YseBP8Xdqb/6o/q7/iqa9mz2ABcAUPD+UcqlPOj6
iRqrifK5+YnVNKIh0xTCFGPd/SALo/WP/fSQIZGIIwAcX25CxWme12LgKXW+8caDf4jqrl3Ca3dw
Sx6bVPEq+Fhtdwwegm4JEQ2vVwEb6gxo+xdS8cN34SETCq59zinrjJvtrpxlXUCEt5LAerscA/gx
F/Q7NMqTtRdPABH4zOpshL25sPW++2krhJLAtQt0fCjBpxUDKzMIPOP2fhTb8n0x5O/FFZ9Pb8+4
e+JPXbIaSxkb/5LoPH5l39O2UI8OMhGk0GUg1Rz5W48HYSyncM5OxSxz6NC/9wCDQMEkl8/0giGb
6C88Shqhx1LAP/hjzaisOD5Q/Z9rPIBDxY7MPmWQWUGTL5e4i/M8V9UpvvlPKC7DGBZNhFPMFgWU
ZqNg8q/n+bd5FcIUSXn7XR9L/kqNeLwY+B24VcgJE3vgpIyrFhIBZSCQchFpczzvO30uxJHLwZ3v
ZsczLbTtdr2xegWxlJp6vUEBtjEFGx2ZZNRUW8xVCXgOZMyDsPsDfzBU6D491mrLVECa5H/+PCdS
NrD6szMpsizaSjvxajzk26T2fv1Oowszzh2Rj6n/bVW6VPKmEkNf8kaRHq0pXdnGiwAs/4A91eaT
rJyn7uSwwa2+yjV1juJ88Hl54qp61c8RScxYU4NQktrQNxJB9LdpKZmgOC8EoH90W09D76yEZuDc
IRRLE43i8nTv8dyX7kY1ciGP12i+VpKEw6mDDwoVomW31NV0tRQ3kBE6EjP8pRc2ElCo6Qb6lCDl
4wbs0vFE4mDjBL/dEPqkfSEjB9u7JVDs7tD5Kk7kLz+/46+9CreDaIdUOKju/H11q5YlGrlNrB8Q
izFllPHqdzj5PgbT8kEDgtd08ln6kgsPu71EnoQGX5CRn4RsMBJDpjWYgNSWjyXCzKCjDJCfeG0h
SCqRlC/u5McG83jCBmlkTPkrOfxDL9opazQttzm9fZbPCSwDB8EVESGXPhq3a+rIReJmYwsxfJp8
lhA3qu1hc2C4Dkv7EtPZHNmO8sLxq7iYXGuDkrxVCgBcHDUuCXQhaorCuoQyo5JlYHkF9G/oPTeZ
Qqv46g8ui8gFLimeHH/wh6DUXiCgt1vUO5GOwTakIetGh7ub+UumYwPNDqlbPscLNEOYg1AxfkB8
UlTBShwfCCQ7oxgCICM6ox7TILt5QBOK/Unn0kxIvFy/CWEEIyT0FDFafu4QqiF1pL7zHQ6LoHiE
ZF4ex9wxzsqXLOcAYGe4d6zn3hJSaZ6Qd3pYEan6uLcb9APSoGq+mIvvuCnE2LBLoxfcUen5dLuY
OKRLoc1bJbed3RYlFN0hnJVUzQ9Tb7BiDBNO/pk/K4m98E1Gy7xzs9HhDJtcPyWKvdIilGupPcCz
4SEaqxJ1GVFXbtSt8snavGddX23TCDu7ka9V0nVeHtYvk1fw3L4ZyS4rBa1KrLe63Glhrgg820O6
YZKpI//EzQEa1ytSgXEkMuZGcGGYfKkfRXrshqpk6Lt+94zB7IWkUStAZMewIR/nbeXDzdsWStoM
e8Wgxkr8TK9U5c+qVCYK/QzuZwVSZiXcFTtY0RR3+8EX05d4ESK1CAtXeIONncHNWrC5CLGo+b00
T4HCvtJLuA3tW/nGuO2SWZjAXejE3CkL3ubrMDBEanIkL+5/bNUlthmU55h87cHlB/V+tz96Qh5V
o+5QX2FaEJE6c2Srs1g3ZSIs+Ir978/fSr+JXBz8jojHYpv/E3VhIZQATerTzzvcO0C3zOgI0BFC
ZaSLg1fR3urGbLdZN/rc414/ffgJuijRrvkWi093hVE/ybgurmZM+A2fqeJJSFZtd/+Dvf2yAwAA
ZLoZeigxIJtj7AeOsfirVp6/kl5nXvcEa1Y1cLgjUaFEDmHDbOZNmbj5Eb9X1tm8V+eOUicmkAQA
KQhVNTPf/muipL1Sr48P+G+R4Awy81r0vAyDh+rUNzQe+DL6nGmO8dpoK2gKDyLavQfn/jKqbUEb
9B2LCTfTs8mJ5/rEolFO0l2FDemDCNaJiJdvJa3Zar8nmBg3jz6o3aVnzO/AixCI4WkvzNVfgfqC
D66cIkYd+I+0HALHIDF1kMPDPJtRIskzB2+Cvvr8yFw/VbPt0m7iJEvJ/t+RWZTVWeNTP3J+qdHe
UpwPS2mWobPkh4oEUnbm+5HDyoB/P8jdN4K5Q2qKRJYVIiiTIoj7sg1HCIFFiCy99D5bvUYtoV6A
xuY2HCw8o4xnEiA9ucWo5YlEvy6S6mE7Yi6OYRGwLBCC/WoW8/Ks7TVK3inr0MVbe7ejSPksN8mR
zD0u1a6kK0KVcGht9IXFybTef7NQBz6GtmOZrljGO06qiQtRYHD85B69VsJ7RetUpmbn0hX34iO2
v+VDrwe6hIMC6ZJY9fOL+8YYs3gvoGZgWkB3GRI24l8gN+eBaMVRzckSMnqlvExwcI+rRQpsnwwU
UKM7oIXng5MdmrswtpIFZvKPui3NlPXPwCBsKSLbfKJJ2jkGGAjuxE6XH3W0XFrcV6ZuJ7F6YXos
lpFrAXiFDErwYa7l8Kp64V+CPS9bFAKaNLXSdo7SC+K64nLHJjwuBhsqmmKM9HnDdtrPDM9aLGvg
7T9FMW27s3z3EyM7aqQQ9z5yIx5Pl7OJKH/KvQCsPhD7swGPq8R0Sutp84keEM1RDh/+cGfth8yE
tKyK2TaZHqItYoypwVK18+LP+vudOuY4nPiMRHACjG9AwSPJ4h3YanLdOOI41ScTUNRtpjsXSPxF
FKqLxebsVPNJZrM2ZTQVMJWbMo4YLb1mfNrXRjMYyhkjsbI3oenv7iDLhCfAQh1x+Y19MB0/65vZ
sTkMk+wXgy+tIZYKWx1z01s6fKxfSy4Q6dRxxoBbgFZ77eWJcgLgCC5qcN1x9HPO+UXY28V0ljex
USRqVsPH0rXl3sGh6eXk/grLGGMh63JwvNSozPOosiqyKYZ7dAkvBttNzVlsNvnSmY1rdfsZNFh9
ntIJ7xEB6XGBGTaN3Bc5YVwgvLJupB4E3ankJkgryo+ocg23WMvu9qOhdGrMoMpeSxGFWFceL1Ji
A0iDtrXmtgwji7SK14Vwa3eiFoeXMTXAQ33rq0TXIPBWWYDe64tOzj7lYVjA/YzVOiy+P5p2tcS8
VgicFTz9TJtvXS7ec+7RTKj6UEligreSKrSCvwhY2ejfQzLzlwrBPmFLGsCsZ8G960PzxpOn94WD
ez5qRPDZZSBkmuFVpZS2JC5vOrxzYdatiJ9xkD0XTspTV5CLghCcw/XopT+1/4k+VG8Th1pgEGNw
L6dCINQXZ+zpOmjRdsU1FPstaCR82u7RvQKGT8/7LVhxpc92R1dzlDx4Gl9vjZwFJG+w4a7Gbf21
hDIW3NagLIpJiw3h7N0jK8tsfqyQOXmZI1F/ntZzAd+r1TR51gsXtn36BATcOX3kFtxv8Vfy52Z5
8M8KPEJQa9kPHoWst6C6HeMPC6tu+GYM+csL1RlbZzXXtatxQzsaLw4qPwp862SYxlenrRhw+aq1
kNuCWs37KiotU7/npHSfTvufiq78esSCDX8NcyZKaSiUXJ7OAR116llQ8CHhcN3UnFZNL9STzQDc
QkUM2GUMUxqLXOXXhkDEHQKGllMHog+fTMEVAchEADTHur79eN5w4Kg+AJv9473V1W7ePoue73Q7
jStVgryWc7THQVqqAiWcTSnq6xVGz7aNMBvz2bWyUUZCuT6ORnLdfXKf6Q81Vbnf38+vducGM9Xk
/t8vehu6nPdDbPbOD5WjLDNefutEdy6OVO4oTLMcqcrSt/83H+yrCfCr9z5oQQqOv18yXeAOyNrQ
QWGWjTYSOItJCN8OwDE5jrq1QlitDmcF/8Jp9kY7uLhR0zSa3gVll0+z9sMBwcp+bzwtRYWarQTc
+BJOR5/gGQtzvU5rw3uibbCUqCYoUlbbGnONtNEryjz7BwG9lH1T5wVj+pX82cc6lD+8z+SAfQca
uIn7umzqarkWsvDmI2xo5wFZzVCtg9AoF831WstKI1eRfXKWrQcMtBc6Ryg0D1G+G7MA+PDrz1ux
BHa30PKfsKdpjt8s57iubte4/UhDe97pPLn9ZgzbJDr2wBrk6fRyH1hFqI2b3GgEMDmp6ZhJ/MzM
+ZNINtuUFYfEqnsk+RwK8eb6xOMQZeBCNFa2kza7tFlGPTYoAnEykALPz+Xy1JUUI1nvhvHas9/y
EODjOIvihVdZYjUZ6MA9Sb7lPJQNvdAr0ykKvrKnfZxqMUBbR3Fx70jaYWnaKACvmwuVdbdUql40
UZluACzWUU53K+UdTlOMoP3Fi/350AaZhZlQ07aENyrT4hGOgDa7GcPhK0jEvv7k6z5NZZYmNOd4
iLIF7UXV4bAWIx6iIpC3hUG4p4eELxD+AcogWKj4gQv+Yy6bhDIa35h2BYjPmwoZNM+xitSaO9w6
zHuImRogJpb61SP/QxYQebpb+AvgnBbNeSyHsqEhcVMnIklL/qPg0QppUkJ0LVe9fLet3fmCtBii
mgZHX+7EqAqGp5kRCJdP4oWWnXl9jIshKSq5ww+Qd/D0VJia6oSoIujiaDbsDnrUTbc5RMDAuVg/
Rpxs3ay1lQGo0zanML+LLlCkSGd/AsXXTD71HYG+LbBElvgZH1ISCY1LWNDJYyAQimkC0HiG6l0Z
mCh+XIBuXwfPqjRg/behUMzcilCoV9FWx9217AYG6wO7eezOtxQFUMDeIgEMdggmNW2AXxwBtquT
UcEDi0gE+Mh9P/fjn8JXV5INP2S/Ucg7ZYYch+Ye+D7P5b2FkDj6WIyT/CZx7v9z0rqCN6gJDMX5
M1GI++eiCBxbvyiU5d1zFmrpGB9ztFV4F3Zg/hXK1PFTJYZ9blzI+JlBmA0GOkWIN4PvnDxZRZ7A
NrCzwBXFY7xMuCySxjWJDEG51KscKaOxJdao9iblLoc1IOrF9pgdZQ88q2vx55IljBKeS9jO6+Tx
DKZg0iKlPnf2W1JuHpnxkibLzF/a9iqa7DloO7ZgEC4PNnDqSqcW8NHWv8kS5tFpwNmiVqowRnmU
0auvJslSyTqnYuZd+gPtdJ33y70fLpfbZi7J6bK3AAQFdVmDRahUnAZEd2qIyoFl+3CGvDGUfujA
VvegCvjE2nTZjboGiwKDCpk+JezcjoA8Fx58qCBoms0Pp84chD+FMZ1oUYIw7E2mAXvcHaFx/yFM
+GllDMZ15AzGc0G7m/uJPgs6ijxsTs8LsbCLhrABDWU/r7USzfYB5lfE8HDRYacSST0MhTuR4bHc
oLMA4k52+5epSgFj9pi54zwVt/NaYPZjlLkwIxRaW/DBouBBmSSefn/cnlVtscWU9w6iJz+xD1Uk
+bYcsULgmw3EHuD5Fd9YBNSiOijsTXKAucDthSefo4gxOmPx3/qk6J4/svDEL3+2h10NM14oW5sY
Qbo1G50dg5pQcobUYyUvL0u5kAPLvUT16828s/ubamEc6hse7ogV/YuYk0J0DL8DxEECdUL4b94R
j2S6MfBs9KC7MPestj6C9WKkwoXMQLmVPzW5U9zRfrzvR2zOj/35+ydHmdkd/ssSThtcbXVicy2M
QI3C5R5M6LkIsaca8RtsIFLOCEPqVPisjdKdhLYYPXIBdZCfqZxDRp6FslagYYpJ+bArz0o3dW/N
Wab8oICfM4ZtdboPm++AOQuRQaudNaKFMhH440ibgvdPq21cs1hS4Jj1XPEDCo/1IswnxARa5XN6
cy4mW4MU5blwRcLJ7rvjxwNao66dkHbNed+ovCbYb8ZsHo64mXOL/0965pNE4CXbFFDa7rnmRlu7
h4FS+4Ws8DmSXZvXTiYkCQeaZ0UrdG8ykiGA4tzWnIxDGQ0IKvORdk9K63wgyQULfLtweb1D1nf3
mabdql3WbnoLeOzWBBAoeE76UKk5qsHR7SGdf2osMMbM00O5uvndDFyJH7loQpVodF775DH6QQHd
5ilr40Y1qWKXs1hbCUAsYiwZ/SAUpp1KJG/Xu0knOV/ptHhSBSs0uufYJa749VzKLu0up/2AOtZn
428OwmoNpYW8vn1AB+gukL6byOI6hWgfNE1/Zd+vxlGJAmI1V3bTuGZmLxN68bNl1jw/z6M+0DKw
fOHiDSk2yIDRXy54eiBPeRBokYYNDEMdRNPrglgz0ksM9qsNgGPR67mVmDwFNAoRtche/8A1qTF0
uP2xYo8SPIeLjgp7v6DQy5E2ax1ClSOgyRFyTdV+guo5PBvORM/T70YzYUuX9QsmWB6OelS5BiSL
BjnsprHyyST3YVRjFDBeVM742266TuiyM4OGs2KPLJTHnDqnBa2T04Oc6kUSgUCXBIIIwJ1wQIRC
cZp2VJO4EOZgoqNAYu5JmSUWAIoMlXVdCxm6dBW4G6nBoPnZkKLcA57bq0s77mqllG4hYR3HNOso
ulLM0sPf6XLaiMYQh69EYjmoxvNtzxxGobNTgsl1oQKhvrtnYzBXnO6XBXYQTFNsW6P4XA7Q0V3A
H8mqFZMkpRqWMxqcD3RZPBYnkrR+NwveTdjjOLt+hnncB2Gw+Np/y2yJUF1Yr8S2+djv9phf7/oU
+zG2BSUoox2CaVI56ONCdt3zOK1EBBLp6Dg8J9HmbVTe6E5+JIHn3bbsRiNu6s6tYxoiIaj1vU3n
4DUkZ/dwH25R61vYvqH4j9v3i/vhPepHfkFp+Tqi/4tkmEd62BjezouaUm5QXXHhRX011OjzYz/n
xBkta7GcPor/a8Ohh3Fj2rfPuZS5jgmB/kiWmDLklzwjS0OxIpm65QhtWFjxK+0HU1phHXKhbz/q
ZYQqN0c0tXOIPeE4PMATqu0gJ7UTvAuXCDxW/SSbie7LrRcoIjhZGEzyzt9XmJ9uNxsy0L5S/fcb
sbc2Oasc466Yf9NmPeCFCTEMlQ74LCRlHL6lO5vYeazYqq59yMub3Bh+b1WlFSlF/Vl+CdY64VBY
o6O4vXf+O155ZZKRnuVXKO2hBAANd9r2fZpdCJZsh5j5nqXtJu4UDLQRhcL8uKJzT7HgTDpeRBVw
Oo0oO/GazyKE1urcAFrOmRubEGBcLyqB3PnSTvY5iv3Go3lzddC5uVfziAQuv5wQaaFK4DaBfLcr
a4Jpt5aami4p32BW9BmvocUGMGIPj2ph2WeB++jX4xB1vg9Kg5oB/qgBxqVhhSBqXPetbe6lwrYa
tIHpWjHD2xDx2qAG2+3ajC0pkrLsY2Xm/vvLMZO61Rwt3CkhjeCgThruVaiOdmrw6HGEMVFJ4JbZ
+1DNY9Jz0tEIFFR+gL8r/+SDTXpVTgq6SjT+/1m4kRS4u2RRqTGXXVYEf2iJOsYxUEj0tz68Sxks
O6dkDlg0lfujmgV6d3TgCJ88GR4gNrwDln8n0WctpmHHlUjdpx34cvsNofn1M9Rlth6MsyTY3P9h
bv4DPt7Arg2u/VffhoMbOuO8l2e6IyReD7Lpcz5EMFNlF0SANCQbrdS0MzNhhg9lOY2iqag3vpl3
xriDjLheAyLgY6t2BhRFIew30fM54nsuZ5MPXg5RgAC6WwtTR3EJ2QJvLzF1DcLb50VL40GNBty2
elpwZi4rKAEzGf8yTlugXpLLSHpjacUnoLtA/v/Dv3Ibtfo+L1Xd9JTof5XNe2Bwk+ISQ6O+3SeC
Lwv6tee63tk5vknuCYdNuGoh7k0BZHafbgQPdjYD0GeEo50Htb0vUQEjXi9bwoNByJm8Yj30Iral
NncHZB2Rl63VNZ0Mw9C+oyxeZJwjOzEpxghwVlDIIXc6Y6VCXq74eJDyHDst8t6rGcAu0T3vjzTE
yLi3+C6cRAKUuW2Tu5krkstZ2fY7/mUbnJqae6BawEzd+JUd0Dc1f81yDRU5Aw6iOnZkjVZ6agVD
06y8c9WEMXzun4HPdLb9F+qGkzg3yJEcKI0XlMK29xssrQ8LbQhbcaudT1zCuIrVsh5TRSE/rS/M
QCGaczUPPIkMfGxniZrtUFLRLATSIDi251nYOfkTtGfmJZMjwT2U1WKohrQFeuXWQfZV1Tg+09C4
M6LRKG4HiSgBVDvX8uw4y/OcPYQVYAdqTRdqz/0orSI/R4/msxXCjXSK4zI0dzsHorUlFLVDXo40
scvkA6ZJNv62B4n+VWh9WOGM9pdcxAr3VDJDsv6M/H6W45zvraFv3MW8dtE8mGl+s6VWNUxBDiTu
Q+c8sOVpcaPxZlFXf8GcGlZhvJnBGL11bbQs1XzptLlQciCXg6agCLyKqLkAgPisxNkM2Kao2TID
9F8SPiTXFP7qUbHwoCAfh6CI4O/J2KCPqTlCJb4ZwNkjJT3RU1WP5Voj/pyVOP6u1BGKpkBg6F3F
5pC+I5Wgfm+nr5FzN5YExs9TRWsBAsnUIMTsYclha0J4UWJf3ZMED9e5HTw/5Vmb1xtdniapLMto
AZXUwYBDZ3JJwTTwQCxfa/nq1yjntmaGMXoq4a46bZA/UfRdHYfaxuruQjD70sFJyweIR0yb9uQa
iIGLr67N4wNZPQJAz1o7DhwzI0zRBWO7MLAWtlqPjIjtWSYYbkn1B8LdlPKycfRBvb3PDeQ13VG+
2sIbeqTJyhs+VLSyjWPvjHn1NCHCW+vTnXlb6qfpDIaoh/3CaYO4Hapo4o0B1mjExvwu4ypvAuh2
TyDNjlx5wq0LhwgE9mJaDd0BQ50f9YluSMRj0uROyJPgn1FofIJE4Lk3Bt/qTD7D4PAPq/h7WRco
+MgsOAmXU3P/yqHa2PxxusS1rUR3+b7pwDTwP24hAtH8LfqQMe8FcRGc60OCxrnpqnw44dj9Mf1a
IO5ZEhgrgdTlol68/2gwQCI4HCIn/N+PMOfI0fw9/vEZ5WB6ktGcuHRn0OEhpaptwQPtD3oDJk4x
enNNc1rrZkbl0V3fQxURgObeQRQMc0/AI2LeuJb1X8VhTAjoByc1P3PHUDTBgPPrPawz91AGYAuA
N22RMt7an6zeM+TW1ekjXGck0Y39Uj+smmCdLt5LSOqncW8KGNC2BY+xrdZoSw0WeJNry1K7CJS5
hvZZGEQfRzfIo6l053SS6jLxA6cD8XH6u5RxGEzJfOsUKPOyx1++QUAaqTUzV9Ka7vcloJVboX0X
UPa1LXos25ZYQPtWWWSEkV9PlEG9lcSTKkQwIXokfPirrDEprKTf14fQ3qA1ad2h0ZsSA7ohSjhy
b9YFcmO3eiWZbsCSqMWXMumdIQOi54OSyNILx+7Cb+8U8WbJOhnZuqxvfJ45qV+aGj1fXNQIk08h
ssN7hq2JvvB6qenthmtI3AIA0ph7ZBdg5/4cJ2p1T3l9QiBPgsf/CIA+8945lUi/E0vaon8i+plh
rBnx4ew84ZjWa5eLCDHVmylPZvo66P0E6A4yk+mAXyqA7Qo+VX7+zDVpcnSRX5w5yH0F3qn2GFCf
v8k0gJql+Mb3QEqbB18Ctwd1YWHKQc2O/4+Xgkd2Ig==
`protect end_protected

