

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jmxpJaVr346lkZ1a+LoDVE1gRSFGUifNjtRZEnGV0oAexMx3qGrmrMofcjVsktZm1VmWfXDcztXM
2yFG9i0kgw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dOSbcKbKyGmwastHjwhWcvg7mo0iC7nVbxSBuuKDePvzqRHFROAJKKkq6GTW/pekpDi7EYOWgoc3
vu3a7xd2BbB8KPxJrQPbDcHKKLsfi9Qu05pG8kNfZPTmVPdeph29tJwJuOY3Bue31aDGpBx9n97J
il8TNCf+vPPl3qN1O1Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oj1u/InDUMUdQbb5KKzCbe7WKv0Q1mJ0hkD57NzdtON+OYFVa+iXuwhtetuyEkD/RFkOZub0bzay
EGz9mYS8JrDX4uhqviZ/lNeQvlGcy4m3aXFV0BaNm28dZ3yofXU/BObQHMb2AJcvSvAG3+NK2bRe
O1i9rDUCI7L9zpBAsqwfaKowW/ytJpmf9i24R0N1DPpd8Du0b8109OjIyuP0B6/WOaUz59+u6rpk
YBt+RO2we5Eynllzej7EOx457Zs2AfpyYb/scT1J2gg+ITQOiXue3l6rpuOlPDO2s8UVnv9AEDol
dBES1PgrY5H3iIxtkySbQdPn1RgrbUXGoP3Cyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nf7SNu0SV1jFULe1qPx1Us0aK2tBb+6HkavjcQAOW7vm2bkkBw9TTTcBYW2ZVktL2qtI4SdzYqok
Ur+7+BvPVL9Si1NxET/7Dtm+YCiSnZRDjVxRHT/nOJoMkCyfwzbKJ0c94Mhpx/IIVydS9opk1YOK
norD0fiQ9NScYfnzaaY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gGrec2cOqGtm9E1Oi+bdp4JmEjroHrWUud/ZaF+TGsozi+qUj2kRQyVPKMhdue0iIQELWZ+mxYUS
eLZifl90wtAXYuJxD08Z4LzdxHrYp8+GuCF0avDcKZR6UMS6GdOF0ZR2WdDmkxgQdaVnCHNmLABF
3DC4E9wBUl1YKYXSRH2xT5Tm/cD2sgS0Uobvp+lTtO/g/wUBgQClX1AYzm6JvXG56K4a0tlrJqsS
O19bJe8ailtvTRagvfU5lh5iVeppPrENq5fwhz7scUcyvohRe2r5jixGcPz5bVE78eEpH4EwzJTz
GDGFrWw8qJ6s5hJeVjOB9tgbpdnAFcvyrMEGaw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16464)
`protect data_block
mUvoxO8ohq1Bp7/kdwKt0TUa6qvMo+bl0ZUy+Y2/OrAS6nfys7MXUAMsUAcSLmTonfAEHIWu3cub
P8uECyBk7Wrjg07cd6+6otvZmwIdJAnRzp/PV+4dW02NtgW3R9mUmNsxbf3YL/BXudXt7dSRnA3/
ygCgnN5bmM5BW2J/UobZ9yZB84gPyuFj7NTkxQo/XRK3ZdqA6A6EAh0AhgXEhqdPUaF4J7Lpy+ot
7D/K9HvxpWe4/Ekq1V9ZSmRxC1i71xNbWAsnmxnGk0ZStRDcpkF/77+4PuFi9QP9dlrsM05wn9rW
aOl7e0AYgtHBkpwpfuBxbzLQlyW3nKEXOQ+Pg0rD4ZAFBzZmmfrKoZjR1EyLXkLkPvY+I0pW6Na4
tu3horDEVd8EiIrAgd4OHmr2mI3gLQIP6nbrloa0hoAg3LU03bsvfe60i5HgoHcK7K5qht6X0m5n
GJMjmBWLsiE79p+BLZQ8xs8dKhiymORKIbYjXtD/CYo1jXvXG/twe9q5C1Ye18GcWaoZAlu/dMN9
AL7chwPMzjV6Z3RAqfKXITC/QW3dxnHh25r5Fuvc1mrd97lycVuJOFUCdcWhU42g6IMhT3wkFOji
VwGddiPccAhe3hUi6H1BYVYGfEj2V8aGOtw1llHt2zNeS1nBYJL2zgJeOdZwnYus7ljenaKznNh0
TYwVumh71G6k2apLtmc7p+qIdf2HcO/p8LTHp12tvFAGvXijA6MQbXdVFM99bzXNgJJ0phxKUUb+
TvntQMJiX4GNO4oT2wIW9i3UHuZWKBLiKmOjzRBZZvyfrqR2w0M4wVhcxSlOKPdM30vakhEixGu7
dboVEhA1MNkjOEE4Gs+SeDIIlWSgOvMxYgnEEww9VDtrKkezJYOgUcBQDCKD2ui+G17FAXCviLoS
MQxPliVbRUKvLkfOBRUKDLFW3VmXFGv8rUk5TjZzHjgDT/71+4RVuFhXr1vgW2SnxcQDgScvt5DK
I8zDi8KjRBICOP2ghmeSSCypFHoSksC1pCGaPMCyObpl9qe+L6GHs+W7CugqvA8ObbS9+zhxeDgQ
EkUP9uronNTgLN+eiOY7m19VjsRnW93LWMJB1ReGUO0r3qBob0UbKg9B2XgnB1OXlq4rgOZzIOYE
W8eJSJbSWINUJs0mt8qDQTVAN+IusE040kJWmA9n34E2W5hGBMO0kDLvakSfjEHhkBxoeTMXDDIX
FUaTYFkYCWl1yLx7P+fQWWDeyCJBmHEI3qFm7iA5mDxPe+Z/NIdY+pUcxMREKwJ4siw3tAgSqN+C
LsGxzAcV4QOl/7f+t4Kh0boSUC/3XxsOkARu167RmUp0/3j9dI8yXSrGsnptewzJapy0GmM/klFw
uNXJSV2PuTdMaXISGP6aZixhlXgp2MDebJeDXFEtbwDkPXzvunyhl4XjFfkrVUBNFV2ZskToQsdG
1V3XWtqq1AAJDIqOB8ZiAkbWGei32JC2lLprGYudQi3R7Cj1jnnGLRAwEHgWSp7aa5NlkyJwb0i7
n7ufUjFJRu+jEZ7pdNPhSNzxjiklJphqud5T8hRozu1s7bXNmDUYnr7WE6Xwbhc2h6jByt9++bS0
2yIlxsQSEN7YFHDO0MEpJn3+kEQJeAHvX183byd4Ct87rMYkcWJ04B0PNCQuUoDtWZJxZXtZbzZJ
cQRd/F57QBLIAa4cMm/r6Jsr5O6bixkd3YG6uhdwOm7Jgckr9z58W2nHoIhb0m+/sSgmTluY/XPv
+xaLJH4Icn7ILRGK3Ppq5s+IzAe217Jhu/+uIMrHDtoVsfn10a8GveNoY/AMcEJIBF78rGfSaaVP
wYMWEzgJv2xJVNP9b0Pacgd3Ev0DjzdVHqtFmNSguhNMc6AUcyekBboQnNN0LBM69CKKvok8H4PZ
Kju0YcAf4G5StHFW5eltgYpwQw6/55+7ymQHgQDW53mNgvU0FclqPib7ToSF6kVjOGq5eYHV8cE7
aorNutDjkqplnCOp8/8vUYREwjwAKINB6j80krQb7uVaUsPLeZ6W/Nwj8v7J1fR8BFVnWrwyb+CX
Pra4R6FUe26rDahBk9DGnPhUhGdhmYVMeIaJ9k0hYYTqassFW9uhBOVpp4YgJSiX4u7V6dllMB4q
Bcj0Z086aVEitsRcM0axtVs9S7LxVN+J/tQg6eqNRZX1xQZI7igrJakFlsFVg87ID43h6/0ISiAG
FwVvIktvobSaf+qkwgKYW/NfMLGIKvS1HgF9My221b0GMBGjtDi5+F88qlM9kWjWEMahl4mYMoZO
rfkN+19ZKPwpww3gx/af29mXW/CCHE2Uoa1B3ShUaALvLIYvmPr/+09dusz1WDZ4+owGS63sMBiQ
bjPu5mQAcPJ02d88zblJNQZFuw4bN6Gukg2KpEiKMse9Q7zD4wsz7eCnfIolmxr3OyHw4QUn8rxR
oAFsE4UxzKXD2skdPIHBaR7EWjANNiSgmmyqPSO5BrGfJPv/5UcCgcF0WduO5X/dDg1MI1qgfkh0
NDXXxA4vmqbpdzYKRVyx7uRojCnC3KKDKj9vho+Pxz5wohWc9ulK87Rq2fhvyvh7f7C+RvoyMPH5
Hq72pGJWQPUccrzgr5Qy6codM9ssNirXr4RsYJwYAYKQBIY/cn2WyQlELz+/3vsaj7bOY4Ft1hqU
g/2O7CHe25L4Ic1SRtr81n+2S8tDM00UR4ZubE37/7+vAZInZ32MTxk9+YtrIv14uCgbK8IWIY25
Bc+MV6gJwUQyQ8euBaKpAmI9InIrehhTRIt7d93j1R2BmiEiSujhwwDmPDp5vpPvDSUV2m9ZzJQe
5VCp0ifwlGYHqsc2+Xaug+DV5xM2pSLwERkLSLYPWVv/RHEOIcMzkY+b6Vm2jJcI3/5PmSWxqxoE
Wa81VqiG5JBMbYgArWA86lJ6XYxp+SJuHEYwBCPu045LjfuKKMmT1b3gJQvmWDMaTANr+k3U4+yT
iZuOxMkrtZAwRGUGBwD6qi8+EjGJ60iH15v7J7lUQAJu8AnXye+fUGHc2we8ygBtkMTwjoABJKDu
J+mksLUUlf4S+snpDAv+3hNXmTUGlSuCqWTf71Q0QtaZGtNYPSZfmJcswuxnHbl6+TOvua8StRQY
vL4nll93k+y4dFZ/pJxUt6X30nfqrsP0StvKC2w4aSMg9feoxN9a0SYjS/8lw/jLfL+N23voSFe+
x5QF9SUdftn1Mf5GohLsD7DBt9mvOIbCxvfk8+GRK8aAkngol3gvR/0dF/SsZErP81SdhyAU+50C
ERpSuxILEfpmcX8J9GymIGxgcUvFVJbFBPlT1lp9V8mIp7wrxzOqJPV2V8MCDWpDOclaBqaCZtH+
RS+5zopnXWbihO7RvgSA3rakYhaTfLVZrJI66r+kmBA0EFq4TFycSmOMQdRQS80tqm4TWgwrJ1CW
o9pP3t4l+As8C4nXzpXGlpnsHAbfgtebcOZQRhqcUgQokrz7/Y4BIWSwNTrTVUx4/aiPk+F6vqbp
xGGsP4S9bS2UC/a2VjRvLYqHO/V32t2zpB953j7mHfzmsHRgFB3jc1NOGh+cYimYicjA0bocKC4M
ZS+B7uL5sisMh1Ne2satC9uT3Rq2ObvEisDhkc52gpEGTQQbSWfos2RwMyCRTn1CnlpZ3qSp+oOH
9+q8fng9vvP+3l01jqcsmxM32z1IgaHiNN5h2egb5l5oaQYDaaM5ETjfgVVn0uXQClyoJQYrRGd2
XcmRqUFJGGms2A1VqtiQ8TGrJdAApwDoUv/ZhwTpYQI4mtCWZlpiEUBZdyFlm2aLNOiDcGKjRkMb
s7vtKGKZzehL8/FVVUv1ewpXBjhrREnDWMWOdS64KpyGs7vz97U440q0XHF3Rx1cwsQV1pgP5b81
DigOxAd8oRn9b+JlD37yggW5xNt3MxDv5DN/JCqu8kIC42YE6ULppVszY1aw7qx1JOlqIbgc9jN/
UEkbdSswUf+6gTkS3di42zf+TfE31U6KbcN/msKbNYNZWU63Vd1CMk2tr9B5VQdYPDurWa16xVDL
bBR2YTUqP943PPMJk9i4rHvklfgTWKyFeAriK5lhUd8ZVQ2ZefpegALwH61wnkpoUD7FqKn1QEF3
rOjGVrQC/wpRrWuJgiRT/NTGSbCYck30o7Gf+hnqysofn9b95uA+IQb5m19Y5948oHMXiIkHHeX9
bqWdw8xGrBDbp025CVZpBItmvuW3iJXSBnkgbcOr1evLbtGT9caXDOp5pb1wZPFpqBrMGaigDl4y
+jZSBYPpEVNxQMY0Xeb5ZnlZQ0uaPJmIUScDrSDeoxbiHyQ0IVgl4WjMJYmsB1k2U+QL1DpOMw1r
JHOHVZNjx92Zo73QqtkN4E5a6MvL0SYkLsp1lZgsnBs1HRyYX53kxC7Q8r1WqU5BQPZeVEvMLRIl
yEmpKV+YfoagtpcYupV6hqEAei4wRCeeGNnCgp1yl1aXDugVBf9utMyuZ871UYHaL+guNdA9KUcy
b9+JGQD3hoXNGH9m2DRE7GgDE/vC+pMRVEuppJeQ4qc4PNcD5AZE8z8Vhe3rybF3NRhGeMU/jjIf
79RvfwyDz+Ir31BvMHi7yHgy+ZQ5lMINoeyxT6c/tZL9fofokreXM7uxvySdQ4Byy0tQKtqzMwZ8
El4K7GKBSYJ+TAAlXZ5ph47ElmHmPG/d4NLPQ1mvBcOMFg+Qmnz/3+LfCRl3v9LV+aszdDsWS3pk
VVKiMkcOkbFUYobL9B98inMITvwFaGv0lDDkHh0yGBWo15KGNdL1plmg0l5Yuyvhnoyr2bo09oie
yzUJfSGqnAoKTBgTVRjfQH6FxQHkDp95rtfarvVHj95U9UL3jg65B6eXmBBoDXufFsfeVfH+yXYz
aCvj2hI5na4gRDfBlKBNZ5SBgP2iLBin5Ow1OhYz6yqWd3Dj6RvtbZd+W82sq/PDST7rfQRJUNE5
YW82/xgQ0e2ITor4+fh2E3EGoIy0rjokTXWZBvxT5GH95Xjv/1jPCBvmpGHIx6fbazz96KZ7HC2Z
Oohu7Iiv/iwbAAf04tBYVTAulqcDK9iv1fNaZn6rhi3UTYGeBzPDEDsFTwEzfWFqH5jdR7cl2CEF
Y9tQkGy5VIIIis8DWB6j06O2fwSOXY/4X3tOmiEDC3Pr+G0S6e5qeqMI6w9PSwgGlLnCyUkzzy5Z
+UJo0u2YuyRb7pIl8tfzz7xykmYyltdIHyNlIzr8cRSp0pcrvw6FIqnc/wnme0wZrMfB1MKdVi9S
J3KiQGCzLY0+EnNMNw3kclBsnLwMajInxIBBBNT3dc6UOqh17C4zOBJ8Ecq8r0VE9Eh8B8P/lW+2
04TQDR7Zz5FMtUjTLfACPkeATMKS09DvWQX56WCS+rsfcA/p6cfJtC2RPACajekpQLnrhtvvH+kE
Vzab8kPm2UBdV7VNe0zUyoEp9wZ+wYjKSNt2Q7689vzer0zoACJlOual+nyA5xBTCVr7/0Nud+Jc
vuN3jagOXPJLQXFlsBtmcbsclXK0vPND/C51rBNkGnNiZKs/Zjc1WXE9+Gs0Qkd0x2kEjsUaZgjx
vN/nNw5hRw2TIY8RpN962jIKDZUGyhTqC3ElC1bRF6oNLVHkONlH0Cozf238eDJHd3Hyn5BDvD+G
9P83y509iFzZOlfn4NW22vXKO1HrRrdxHVHxIoVFeNHnAnJTpfNYo8MxXfQapV3+OKJa3stouohh
NP3cZMPrGfnsE2nJkvt/wchMgVGLDTvTjpAc11HLP2xyaRrfLmfh8MVkvoJN63KaBosZ/NDOrfnB
eT+ZHNjYEH10cTDh/a7KeNdHN7bniPUrzINIEbNwGGY2p55bZEHiUiV4fZnygI6PCrKO3VM/9Ry9
zc2S757z4XWp8O4ZgrfNGKfMqwlP7ERXYp3lulsq1d7RIDzIRnMSQ1U+tHBusvOv6hFppTObOlPS
7lyAgKpSEa11qOkWe3lh2P3SlLM3d1+Fh/57gI01L4PupK3UBwEGXrL+BI2eNpxcDZGsPvpFYHSs
OiUYGK5qNQwxClJS79PaVmEg+UMuXLCSydZjv7WdjuYsw73TAj0sZcEvluL5KIVwVwWYkUYy2V+S
9uJUU1u0k/G6sxOopuR6CRIKLCjxnHjjl72135Ljs4fcRdNV8NL4YygA8rDb44CN0673wBqxitsL
19sczPL3g6DoloXmb1ccj9lzSSSsrIhbNql07b5nDp9JyC+Io9GPz+wQ/xHRf1PxnhTR29REHUmS
LaM0CzGq69JHlDRkvYfGnKtwcUWo1TRfKJgi5OUVNikCK4K6PQYG+5WY8Yb6Q1c/eWF0vl0u1UnG
NSqetlxUNssW+7WiSO8K+bv4RR1yJXW5+rOj2oDj3rB0BfduAXtJiXg7tP4sgHT1A2Cq78otkMm8
TN5gjJsbNUOvGpWCEwXnp6jQhOMtCrAtb116dV9VxhADep++GXoZ6CsA+8t+FCHMUHziqbRPn8c6
Dxf0PLoqXcOB1bU4YJm58nnlNtMDcThkKFGeqZaT/IjHCkh4iNNqKhjjYCDOYAc+wKQc3aHpE5Mc
dEcC+kWpedkYYE/ZsZQkCDkNiGo0gMajTGSlb3iMZvJhU9IJDAO6UeZOO5xZngBdSzEzPtjUqP+C
XECjhEXXzXsM3+YV77rA79gyv/1E4NbsDlZe5P7AKHKftUEx8G2h250uLwBOKo5sgCJV12ltMpm/
2zgQfCV7XpNzw/NqYFu8BWJLIDxftCxBPoQl0Wu5s8zlwR+FfpgWbxM2GDgrHLkUdVTqnbWMkqnw
Z/OteppLLJ55MCkXHXQdZ93L7DAb1b+PmdGtI/VrRG7Pn/btwR5psyIRUBEdMgeucywLGvHROaZC
gPmt1Ys5bCQrUZe0ZlRYv5ZA9f0iG7U6ymstFkxSBGlwsSm/fdkTZwV9heNmRcGwyJHGZfF4aExl
ouqwlXzjlLYSb9x0uHdXoWeljSOE97G9BAnPl3ndTOZ63rPaklO+sqwGFUHKhmv/ZVHMaMUU/rFt
5c2QxBSykuXORz7R4M/4DXNAtE7avhkPWpOEUoL+uRu+NHEURhXJEjIdnj8Z72MUgLAYdMd4njtq
pLVfsH9XoWiUXX/3P0yySX870QfGHy634l+W3rDT1kDuLqKNf3Y/HcnpVlHCGEQnMDNXKphnJdIA
isKYcKJWIFVd7jnOFEa05lET6eeN0G0sW3Mp/tWb7Xnn0onQGVOea6WB18E9GN3rMn8BZs9e+/YP
TJEa7LOw+PX+EekFKf2b9S+y051ZQNekwUYYTAdr/Xos3BFkJ6vG3N7PJ8qRcekDVKIbLF1Jc5iU
ak+xObFuA7gIXj2944MhVAJ0cJBi/yEscsApSSXLHPXNaZtOjFwOx0vj33gLd6wlTEqE+wHsr94Y
mrTaS4F/d0dydTKB1EdM3xbda4bQK0oPlxqzsdkUDfvLjuU9sYlAne6AGdFtSFqHHOn6lQB2G4K4
Gi3J/fQ9LD265u7kQxAhcVVF3JIoDTTIY3UHCwUgC6aG21ltw7ZLRlxQqrFs/6m5EEfji5HPrZfa
La6agoAw3AEy0LMpgWhCgACJVK0GZBLd8yyJB8qjkSG0HrxJyCJSAMwNc3RsGtwbqrFgUOmBRhse
wBPtliWKd52sCbJV0dZ2HKk4JZxXZxJwgAUU5c82I5xw/rtITUacDN6TSZ1XsQ7unPXDijsARc8B
eMtLsEPjQ1SqIrh1av1RHxbQWMvjs+fecCyTNv3B/XlhC4XqKsK+qVqOuxC0/j2HoU4ukrctl85J
D8LArZ5M8F+YQ5kcrm6vTi1KXDN4aOXOW4ISrqOwfNNHEBiVtmRiE3jOLWvt49sMn4jwQraKPivs
4v2MBP9AD7q0WiOvIPWxPHr8kFZWKQPthxZH8pp/KMX60F1r9lKx3m+BqIwPLUfJ/s8MnGmTue/K
COpvBvmj5I8WWAz5UeMsy3AGESKEFxa2msmP3Jvz3Zln9ezlQnGcTPqv0IiTm+FmvYqQ7JKZ479D
yh77oQYse51FaXngH/o6jt5a2mV4g1Pmn7nAYjrtrEa8quUVknKwntforQvIzLeNinMAl1ApSvRM
GY+qwh9bOaReeBqW5judp/guhtmVrm+UnqDHAxcP1sUyI8XCw4GPybur34dmze5GAv32clkbH77N
aE0gY9d1vlb5/SzF4EHt7t9fz+dNzWD3L9FW4Gr3cduKoyYSJpTxTThdde4j9Z2Vm7zs9SfdCIQN
UNsiyZ20545nWu3UrD7vuRoKax8FiXE3chm4Fzf/h9bf1yNZt0ed4NPd+unrBPiKjYiGJ+kSIBx4
aOrKGQ+5edb4ahNTS0m5EMQyNTQ5CjhNBg1RVnlUatBGKpw+soEmYTW+ErF8kpf+bcaRX+iAvX64
aJSoW5tHMJ5gxBu6M1NqrAWhl7PbqmwMmV4dxvgpzxmB0O42OvxNs4ygI0KO6eMAYDhdFIKl+IQg
LVqSBwIUQl3ASXpz4f9O4oX07L3HQdccCFAkyh/1u505woiV+4Aa2Qdu/kRLSXfzqkBWCZfIJy8W
zhji6eDOoLilzkNfl9gB14Z/kPCNAKYGDsVcnjKws7mgm6b5vFefM4KppUCAG1U0SVGO+TC/X0wq
vBWXDOLF0KWrzvuQu16PEI0eJ7NfL02Ae2Y/XkUYqPSYROIE9B7nKjWUpLF8pywmqen3UfFNETJp
9SZdaNPBXX0louHd2iMgQGOsHmKuVn53C7vq9uHFy97LB2RzyODw/RkeP5G7mFYVXxAu2dP6ADeW
kQyBLiUZ7G0EGxCym4AzYGwHYMDVaTAPD5ZhA1fVYWyyetVswMxxEFrvilXoAVevW4e/LSPAINhp
a/3tEyFYqi1OQYn8GtHcu7WtXoEHBVm5k602IyHJChOHhpP/Qxjiydt4U/mM5o4sdhQDbvXbsA2v
/xiBnFniSdZaoZRmQzVewt7XJEDJ8txm3pdHjpzDS8IaR56PCSRN+rb56QC1cGjtAO0YLBhf0JVs
U/R31cbg99Gjnrtv7eXzEwkjtK/VwXaM1iIu4hM+kjkyZlfjW6LswQC1v6t6WgHQXFocqgdXFJyx
hpdpo6KlU9bkuuR+KxjNl4pNO/ScoNaK71VjhN79JqKNZbx1Kq5q/1x/PRsLgziKKDUmY4Fo4nZ8
CTHekl2CgjelVV4d2azmtNGIlp5Got5HUdm/bNZAuw2UELlj8cNBW2W04ya1LaNrMxYZmBWDI1DR
KQ/x1keH6/1Vq54r/wbJDTOdMRnewzPPhzBE7WkTkk+KCGtaCdx+CFrTEF9eOEY/mceM5Uy8Os5Z
/I8KR9Zd5XIg0Ee3jLBri76uGEaRhB5v8gCJS5d8+4MVCKUPcguSHHJlywf2VY4dvvpHhn3nSPY6
52Utw5Mi54FwhmYJCCSzYDXVGiZwb2ElJB/AQXT8tuzz/8jlEPSsdxEdTK71QGoT9gy8dgDWJrlT
yICSZ8LsHUoSVR9yssC0L0wA2P+NevnEaCh+bprumZ1yvwZLAvZ2knn4xl7yG1ybtpcVNHnspgV3
A/PoolObPbDlo16o3uDGHWd3xmnT7Ed2k3pvDGjnfITnswAFaC0wXSHceQ5IRk2IU+0A+50nqK+n
mtouVY0V8KtS74pvX6W1etjY3hg3+0ABIPvr7gEoshL7loez8GglRfGyBRZrPlyZ3hJ3NbNXa8T5
XvfD9nlbhqvhlEmyX4Lml8OlsrJ8RD1XworHWS7BpnNFY8VcA+UH4n30blfK7WjESdnQt/Th190A
TYsWwx15PRMRyiTM1KVeiSdtoGWUgEDfr9yzExkFBP46T/ir2Zb8XKVFenxajafR2D1wwWumgkEu
fb+fcEMRvnjm+39ROydQ0p83kVj4GsAMsYFoV7KWUg3ocWaxB4ptA5/cgGnVu0gBiUHJ/d9JYToO
rQz9W7znwxulclf2TgdZUupoyr+bkRei0+RAZs05inF3PT7ZY13l5Qqq93ZJG39gHrBPPKgcC43c
3WCbn71Ih5Kc+6lTvOh9PaqbbQz2QJg7YuzwKjp8wptXh8yyFBjv/wK9r2jN0leOFS0C/++l5Wb9
+tloj1OUqYARGkWKwGxWreroQ2XnbYPv5zIvHm0PafgbRaFZc+Y4LQveYZe47PBBFCHOm7dN4j7p
r0WHH1yDs7W97CSghOKsoFS8mEmHu37ATAkqTqgV+OQKs7K7fi2rIIt5HSCAnWyzeZySEgs2JaY6
O399hsC/5AF+K25DdcLdM077cm0lg9hpwNPm5cHltwIVLPYHDE7cCE5AWBwjTV0k5JVgQKoxzliw
kYAH70yenoPNQh0+nJUayp6tZ9qL0OFmy5ZAibRBUnGbg954g4aMSdycEn059zCosdGhWTPZFTah
co0bIANE3/DfeF5l9h8sqmHQQuDjswEu5fkbw9d0hr2B9cWEv90rSOstwZgaOwbucq4xkXaXIMQo
2ikXwhFze2Opc7e8YsQtiUghUC+0Buxf0hKMb6jPQF5t8yhwdMt3yOuq9tHtKmh4FB0NSymwIYXw
UP3jvo/sqjNzCe+QwR5I40ZUAEskVd4A56n82VKgRRQBBNA+RGEyhtb7F9i0uQTrkDN2AFBLfrwq
G9+Ac8CkN3Ax1/ITkFMM+x32QoPgbnOfgWx04SrlX708fQzyR7+rXUO7zTII5+Xb1aVdd3klHmeZ
FP0b7rrHhYBbVf30YdAmg+MspyULQ3ARWYehPXWaxW1MdxTKcqmymJ77qZZcrOOotSHpHmpuYyzP
UfrCkqs34ZuMJaBixwTIBJ7j1JYxRdVKLxfyptnqLhQIbxqtHS2bE0CLjU6QaFc7iSgIOEt0vyT/
zTyKx6XgFPmw3isHzxYMmBwO6IS0tcDmxOJsBPxEQ0FR0nZgyhx3JjvpUVZZX5vXxjyIghrnKnvU
Dj59pIMqBmAcD9EsUZfCcLX0HphlNoZAh6vTPOKPoyrXgRvzy1UOEpLOIdxU3KGmhsfcmtPuC2DR
NhhStOX7cCress3AygFK//Fabx8Be4wmeGgS7LtyYLe9myCJR1KKp/VKRqJ8yIm4RvH1lm3uLIyM
S+cAvoB4C+QwF9x47LRnbq5tSUlq3DkplJ9Xe36/2nU9BLI9Ak5NL+v/K9Jd3sAWWlFaV0ZuGcvx
7CxB5oHdybgqpUhRglOdImMcJvi6MF3fyH/l17cpKrledrxfwz2+J079g5VNZJhaqmiQowtKAdjv
qb7yufDNZ3XX27Bt+VKFffAGVYUBuOT+s8eBkZlLkx9sOHOMY11EL7BdOHMaLSmIcSvBipvQfcIz
hXFpWv6debEE9XT5fbcUfdiY1LL/WendlwSzYVoE022UT05LKt6KuzmLU9Ao093diKvvoWQ3J9x0
eAtNPwddofGgt9Je7sTuhkheEkcYjqMtz0vJ0vQxMZnvXzavJanNSRDlfgJFJRUBeiWAiOgUPden
vZhn13x6+JQtIfUQ2UPcBm2QleFMUxrl3OCzVF+Inek6W+3N33XGoADYH3FtdDd4UcIu0jzau+Bx
UoHUCZShanFcQZ7KPB/KIkR/hBlG7WV8EwCCrVrgXI61IporU5wz9usymL9i+4WT5D6TBymsEo7F
BcD9B162+m1Kk0wy/ISdWQJ1qVyptebGng4EOI4IfWsEorQcwKUIBlLiGuZfYjir6DLWDIdH33/s
heegufGhYHeozEfdwDKtOqA6hpXB7+hFzieqjwzG5i5z2VqTYZYc3DaMQZ67dI2pFIvoQu529w4F
EBOKX0lcR/y3zZHj5JSziZMFZwKBpkXo2h7Mk0edhw1hE29Psa/maetycCNBQjf/JMpBmeZHywrE
h/PuFoVp2sb5+IEz26EcCI9jyzZDeHQKxFSzFNtkETxsMgzEdJr8qYc8uGsvY37rr5eEXsFJo5mA
GdMvhkJnc3njIl/YZIOwQw+6F4y8Rxk7KmDfY4+ptJFDMNCo4uFJSnf6wM9cCkgs847iO2QA5ruI
Xs0koWjxji/x6e5y1RO2KTP6yivawDzndKNBK0EgxYQNbvy312R7jWFZ/Ms2Q4ogwuhNW+6iMjZn
pe1XzVwhQCpiJlTN6dw853XMIXJECqllPZmyyou+IRhlQwmzNKrZg11NRlhVwgwZqK2j9kVpo9/g
8lb1OY5Qt9t0jUiQq4KWecPP35U9tr2N3SASgBXCzlgHa0uk2dlT7KFBRNxB0h09uyclPYGaGdor
wujBqzX5Uw3hUiADibwivxfJPOyZj92E6R1Gv33VWrxSF5BUWDPxWiTiAWYOZylVd8r4x3ElM3cm
gDkBP2cA+Hz9SZiO9t9dKIgaQDnA/Qyd0uklGFKWHwBEMopxu7gNvSif9LyIs7nNr6tR/j6xbKDE
DIKKqQJz564XkyLYmRITpkYLTmm1Er5tG+alFuKCYXY3zHvM0HWoi8tuhhtzaJOZLpXObCW8oPTB
rIZEgembezVdE42fxBvCq3XQVq0Y1vcRDpiph+hy1Xce3H55hymEVph07L1XpKeLh7E76E+shC1Y
uIU7ts7sHeQiGFqaeJW6Qq+hXCS/0p5ndnrXR5ZhAgSjD3N8Ku7dM8j1L7KxYeIMJaCgFj6R7+0O
9za8YouK9tD/GA0j2YpD0EB2ZAmLJwkSeVy3GbswDi41mEnbr/vPvVD2l19nKulrtFXFyLstpllS
M9xM3BInukmeWp9o+Ag/iCv8jWSY1THNrwdxY05PMckVbqpF+1YRVcyW6M9y682gWYT9DgLG0/ZV
/7RskdA0nTinfPgZOWQJRVqDsMk2+61JIrUtaxPqYcMYofi6TB/eFyyciG5x6IHyf+MTI5O615mX
BTqoKIm6/r0hVz5Tuw5jhoRw+1Ys5IbesRoL8tNQrX9nMhweutdhfkJfR1x3fX1oUApPtb6r13Rl
dQ9kPX95dLAuvi0KLOVyBUhY877mlGX1Ue9eB8bASsLrcQFzHDf0TzHyzUFIs3xSrrJRGD40hUi5
ChmhgpZvyLddQkwKRknZc9ut4EKZmUkItrhbSvHKAxowlddQlt3mzjh3zJhT/BTTg0BvIx/QT1D3
PFepWdzm/u7oTmgLhRZioItpOfsJtNGeAvrCKmJm0Ka6nphJuXfjSBZF8rr1fsGzHleMnnlQcjwt
pQ9nyM+pWbLlOTlqZw+pNKv6ARV6xAT7s4LG+BiWd9LYNzpk9jyrmkvXKZNu4vxGhzSiS/c5AVhS
5CzHzpmntr8iq3Ymi4EChRYf6HIPkUQmQzyvbRLfja527jujsoOUaPqHt+NpDpQ+PK9rTwkDkulD
J06+mC3jHtxIf1/ht4IbDXUL3xXu3D+UZ3Xj+j/FAKXtzhigVEGYrJOz9gecHii/IRF7q6fszonO
/Laii6tN+0FQ9NwrLdmuWlTEzH+aVqBOSo7yWh1lR8AKtnoGSQI8ADxP1H1GbQTMFWc0JfoPPC/u
QfMaKnFVB2zql8mjw1qGeX3cbovB3c/41R68XNujvQl7dpZyf4HRz9z58vwhiA9WdIZOGAcJoeik
fUqhVF6rkoOLxuS6IoRHEn5cc5uF8J7sbSxw01PptFjIIsO7kEIapsK2d7KAuXvsjX9M7yPFo6l4
+m+Iaq9HgOjiuyPqy+y6Jx+/WP67wjaByicQwjp7m56lEov5d77/31DZyqi7gVgUMM6akrAb6kO4
lh89qg9igfdTR8ifbpr+wqAjr4014XIu5+eZbl1Mal9nNf8TPYf6ZbQv0T6QJvEmdloQiauy4WXK
NwwzLVQV+jTTnCDa6DJm7BTogFL+XXtuZOElv960Mrv2eUu66ek3Jn+gfebNeqmZsM4oSaQNbdKu
pAUqsrrniVVQs+4BaFx8qffSzYXbmQTAPKY1Zfu6plbnMq78HP4C3ZV9WDDlFg/0w5BvWuMj+YbU
MiZod2a9FACRfRxaD9LNIEAL+XM0hm7bZ8RCWDzfU6l1XHI9zLteniVz/WKrcZijcskqQXKIamnn
hnjcnHFntigTSxmansM+ZM1xZiyVeQoo1dKt+O5b4We73h2EYVU1itOZwwiYJ+aH9zJUiFBHlhpr
6Y4sDDpWUONeCZoppFV7Fet+c7aTrGdo5Fvn/KCjY9SZwHrYURYsgu10f/tiVSmav1b0lA4rUYtC
XZsJglVvPKkvnaGU9szq/b+/CEDjxhcd0BpzElpqbaPcKnV+qYMsHAUsFCgHvaoNCttnmWPiQNQM
llmysG+0CXcpztaCT1pru2gYl9Z/3wCnf5HQx88imQF2wBYH6GSWm/Cuy2BjLkngF+LRQGUqlX97
PKeavwlCzIV4kJdo5HLViciF2XIHMYv3Q30y91Xn3o0gAaXh8DBD1UlGfDKXgztGG7bjOPHngFWN
HZBT0sm8+Gu1sfwVT3jBZ2iiVo+h/ofpRF2UzTuzqQvKxxpWHjom6mYJWfyXT3LsgQRBFFJ0OQBT
aLCG6gFUteEow20vWQJ0aWMu3/MUWlUhQkHufmyuyGscS58FKGKQVeXpdVOM0Mi9sIkhBKmJILcH
K62Hstnc/f5IrJS2G2PjZ+DtpGn1yqqQxglELRUn4JuKM8K47lbafro4wh7XbiXqudZiNu+S7TkS
bIR+mc/4qQ14Xr/gtoiB54CEM7JxZvGW0yl9dWkEmq7tpjaLOps4jvY7SSd/qfhKQtBOZbBkkQIy
kPY30NReOhV9+Vgjy6RIW4RiLPOD2PoN0c6dtK/li52LZe4+13cDJ7bIuNC1J1dlw+xtTIOFh3Su
mpshIvqExQYagZYhPknHq8Haook7m/eHM/0r5OnvkdXwHFuLkbk2eQrq0mKoVk1kHhGqqxRBzenr
8apln+rOEAhQdb1XvmLDNHgkkuMI6XqoXWcF1A2Hca6WRO51QjHqZcA3fDr7CnjLd0c0TT00TKXz
4EMKja0hj399Jw5m4cPID3s50kauWyH2OfcWTGQmw9jVLAVJJ6TZNlq6W35aUFQRfFIg/ORGY9yS
rOFojYESNLbU9cMFr775btrMBccaRCzMKEBwGbNeumalOeyfnzGzFtCXgJkgsPZl8ZN4Q9nHKUcg
nXzJBLcOvy23bTjAzmOpws9AlvGVQvmtIgi1KysyQwzVJdOHQ8Jh9aisfJxJC8VxZxb2SkrADVns
a1eznd28+Tr1yrL0nrSwej3eVq/5JXg3Mp4AFKhSETQ62O4RHOexiMxPj+u3rkYb/NsJQv+W4eQL
J7nT5G/laXs5rhsdZBgY5IN4bn66mMN6Bv9Ktq387doKX2ncR3SmvS3a02nUauCbYDe+2tlJDyFb
YVHq8bochIQpJijhRyAeWTGL4fnf2Xvikh3Zaq1VZDZWhcBayufgE0wziV1htDf5/waDTglRlQn8
/1m0/iNJhBXLUBEN2G6zvq1VzBNT1RoJTFNUcATwwVsj6sTU9LY1qX1QXxBWacsuBQQvkzIQ0606
YAcqFinuIW9jDIqJaNWKGvs3PDFyVpw8hxC46GaQ6bTQYjC1TRaSoc6bxIecqp6eZ1AUv/M0Pa6V
oGvMNIu7ZUNPEJOtRpamrS+vWes7JTAVGxQw2q8qrATEFswxcbEQUPLGbYdHTy0KgrWz/70Z2mRk
Bger/LK9AKvKelBUw4YX5lX15BY0UVUt662AoImVYUVQrJtRgyKTadSd2tyPfoDeNYf+gRoUcFjL
3ajstvbwY2tX/JtYg9r2+xjOwxIpH//OVobguthejqJk1OWRvjNZIZ0vUWc1Kb/FjmJJa8IEmdOT
J79Yi9Rf8WDBaYtpyF/3oVF58Yym9TQLEa3NHgtzlpA3YQbxBZTDCy2ReEG1Fd6VKnFXvusz/JFH
DBDXIdDq8EksBfTuB5JrkwEW5r13GwJNNisAV/pdQldYyVuhHYtFZfpfij8H8oOgY3t9A26UiTpK
QRTj9CfUD3z8Pm4sYenLd7GIIq0NwTMOhy9c206Bjn8qu3kLXRfn+vkEggQqTzP19UX/jX1XVObC
0+z7xO58Qt1Y4bA8P4l7vZolUBK6esB8+PleskcEN1djhQ3OLWc1yzh5pNm77GMiGF0jvMiPV6rV
LVvtY6rQqtMAxZETcMWTZvSgAUm/nmVJj70Ql4rXnHYNIoQGBZ5xi+fk+dGw8DTC5LhkcghuY6x+
Vm8PT/JkbFZKm72SyR7BgP+UjgiT9P+Yz2EmLbsOr1r6213vVgQoXg7DFpcxd0f2L4/J7JO8+IPw
g3f5+RcGZlkvLFc2a2L5egb0mkmoHiTGgRb1/BIY2RKgdV8gNF7JLWATWSUm0tHVuikXhykOsepN
eo5bFN/uRYGxZst520qGjN9q7TNy7GZXVBt5DqPcXTNWthro/cTGdmYm8kmNKyfyAiSVpFEkSIYi
O+dM1C2zRVt1AZh490bMOlS6rlK/eez6WhKZdab8Y/upFEwcGy/nu7B+ILUkwGuPN+gzRicxt6dA
DWZPEuynEmPIPeWtnmKGxrEDuSycAKNK3AwKl7/zJn+rxPavr5BfwT1el28pTId1wOrNZFAfGqar
v3q+IO8EB3YMb1IF5IjNUonlNeOhYXUiTkuMa9ljmgondu8sn+n5W8py8AjaEVsi82iPWZgwDj4C
eUdjHxkzWg9K7fwArZtVefo5CBmCuzhaLN7pdSJ4OTlV3wWb+p3g4hATNacQ+Oo6AAoxWw4G/kHd
oKGQIkN5sraj8HxC+tsYI91Vg3Y9mCVs2NXlnJg4flN+/tTQjpDHwI7ro6dtMvC5hu4XIvCd8/us
ApitUU+TDtX3vXwwebEiYioOitLwMIekbzup8XX3dzge3pN1L7CcnWINeqRidf9Q0IyFIXaxrOBn
FKIyIFQbF9ybgF1dLIufoxgFOKeRiU1ENaPJ1rcZw5h4uU/Vcwa62sGzYH0JaXClM6Ez5EYfiSU3
cc3NB7fd4sGG3vNhKffZYh1WTdG9KL4vKj95sPJ+3uexoEtn3SU/kqv0elPh2/yM0u7u19BnydPj
quYXJ+kCLSIXU/RvcBdhMDDeOLHvcIwhFyFKwY1sJSmNpH015ZhEYMF4ECr9sa/yEZRJh0EviDnj
RljF3ZcX3ZMqmfKDTynIJkvdejAwcgqTwMfeO2VcKdi7n5vuIJlk2qnIKwYFzuG82BAHjd3D2uF/
o3cAmMfUk/JAPK7POdGEM2sA+F6rQI2WOc2VhIZjP0+YtqVudEOutO5YngR1ON/8VAZmV1NJoiOL
Y8C73lWJ6wMww3n6lapzLSSVwvmdjjYpuTqU/j7abj1J6LJtguUtE02D+InrYEaIcxEAUAdyHpPd
Ee2g7zuE/3uIbQ4aHBZPFrtoy3ZqiprEyUQj8Ot0QzEg/Re9rT2jMvtTKMyRfjf4NGgJIpn4HDIY
zDa2pIoum/Byx3rtzeXZAcSUq5rwhRwbo62Y4KX2xePSAXdnQ9SNRN2vL8ZjiA0+SOEOFgkssUHH
XqSvlbdvt9m6atRMs9zKXa+p14aEvp1zSBiSCKFUXHvBo0VLgLBGg3oHPeAjeLEDxgtqP27UawB6
+hryp1amlcZUSuzpztjF3pbzjCneDmtIfSD0uull4hVbov59I3S7rOgxUdlKuG72UNK1iTdLWQaX
MXia5KtCbfbte2l1QIpWRhwxbwUgM3Icb93oU30VyNbrHTLuwpuWCVMWWYCRzWZVTK8wpdZoeYbi
T6YdNfTw5qwC72TuMJgv6xFtoobwPzKDOb3GYsgX+tb+A53O/U0yJwiDIAtq8Jj4va+FVMeLLB3V
jvS/IYOVzgpSYOuoThaxyLDaz/U3qXbAkHBOoA1J52k4GdxVT+dzoktwPAjbbWTtPlii2+z9md35
/hxGUkjVWNUBeQ6UgTXgY7dJPDFZ1sq4YN8AivHxOhCi9nR863TUZytH9jwByF6dLCG2qvD6XugG
LluEn+7ctEH97IsLJmBCuxb1mphIJFaR24jPc5bfpUyp8rqThJ7vWrkK7IVXF3QnStRJ1Baanej8
dk8C7N4qSIGIzxu5WwT5WKlnCP9PQC9P7v/XepgTULLQ1i/JIXRp+2zITuJc40PcBwUK2hQ+xHU7
VLf4ZNyPAZN8jUMxjXYczKmRzvbzFYLo9dtnH1hfRwgOSYUy3RicDANF1CAsKyIQgqcWX/aFX0Kx
7ZSbmOg9EByZAXdkoeVgzpySLlF40SqyN37josdoCqAnJryx9HpoA64ZK5a6TI4rXg+Bj7dH7Fur
vh7+v7e+wR85QV1exJeUWE/FShBpjgNeM5VnU40dGHPYsdLMkYXf/2q5vxJnHb4Shhm0h7VqIepQ
sBhdX1va5LDY1ZikTfGH4fXLRsNuWxGLt7tIAF1JSSRgysBjQH27701qYP2anEjVzB0+XkuWUPqk
8VSR6sVb4GzyNhujYPMgfxbQg1rpMtLlQ9IyfDstKHtHlmOVcWnyI1Qc8T3hKT9ZYmrfXkojhUWt
montymDYivEcamqawec0nCKO9xJIMSnOFXteMlrnrRqEG6sH8mNLF17OND4jxtlEjWA0yczLrirG
jxn1TNxOm4bQXRtqrllcyO3JJtp/BV+i3owzXNgwgxWnQdhpocelA5yhpPR5nHZOJl1tLcECLx5L
KwXyn0O0+QAH0ft1bPAfeZREBDfCrsuE3sfbLJqy9F/FMLfVQgjENM9BG4IGChWyuRli+B5nYyG2
eUQbymtb97cl73TAeqyYbhCZffKMcc90zp9b+vY/GKxQ3L1QeYnUBSiF5qnEY5Rpnc2GWMfzD+9M
n0a52dVjmReqGkQ7fUotv5jErbMvk8TasD/OaeN+5sDyANlia234h0lP2D/BwMDRBCrHEWqPVslU
5/JeJbQfS5CF2W5Yyo8SnssnUxkzd5CT4Yi0CRT5X/URMuj4sP+nCots4SBb7NqYtk5YOVGlKA8r
zoVZN8kUmgunElnHZBnkEhe34kt/QuEtp+ZXNIPn+VmOf7WGqFwg8K5lQ1uO8oC9WCy0Ra3ppbe4
1XcZO54i2Ioldc/u0ZSKuU+6a4dz8aBMmX8xg1MdQGs+UCFDINguRhL3RtZeD1O9QeYELuieaf3M
FmhsGw7lCZub99WkxfhHbFImwm9YKXfCDNJlpZEyW7IH9+TKF/rwbNikwcrRkt+r3K7myrh/NkIU
cfso1k7IqfjD01znH6YVDX4hceFEIxTfPEKF3fKADwe2nE21ODgpGCp78azCrhalZQnIwp9UjAjw
PpQujdw24x1mFsJL4aOETSYYwUnki+9v5+RwXYji4fT/iPuElaySnL8ROsxR5cnnRykVuSMiznXL
DsJVsjYGzEaBeDGh+52qWRf8aitzOpt+Q3gCqfgCv9K9jsgEspvnzjcNCUGi2CiNfZ8kHgBg/Ard
VuH9LtPyq445yzxptSsIlOmxRk5lDYv5Qd19lTUDupDaYczVyFQ4A3jWRWLdxp2XsTFD5BqDmKPM
UwKoFxDENzq2BR9etRG8r2eQs4tvyMRxBSbQOVQ0170sKK3vkGJmhQpB0KoxrjXqbUhHKtPDUuue
23LQGEkKOP75KjpH3ZPglhFitEJHeMEkd9YjvnH8RkItL0cXDsCMBf4PcdnZJUoK3n/sdldqpXej
NtGsyqCQevIkWDjWfDVjqZIqa7XvZEhvl1gRzEwMrgp0KAKOjSxAdUe8/jRkYQ4vYUsD/F2QLVZJ
dBbMgHagn5XYgs+dbXUs7tAeWyUUefSXzgIfoLZPZ+RR3dN1gasu84u60Yw8Mpveqk/iiXbKNfBH
N6LoBWz2rPC+tD1dGHRZu6Q/a9Id/WvxSCIHsez7rnQ5zPTdPhOcp3MAs5LncXu2jB5AnNncBzdt
YKMQA7bFlB23Rw2CNZzs7O4iijEWC2Q2UMKVM8X1N7Z4dWUXExFFr/kDKmWO81JXWAtezd4eBjSe
HEAmH+f7uwN/JDzYUA0dUqJj6sJ2R1qcqsSTtkmtruv1DPSx3Fks00VwdoTCYE4+vSweVXbwNRph
72/tSEIFcDtISdaqCvuGhI4JH+Vwmltk6Ymw7SPnhqwyJ13YdmPTEfGWTurX1ObXRp7UAcxU2Ldo
71J1T02KEQSoP7e0bxRnrtLl70zOABpaSxXaoxHtf6dV5GksQ/24VIHOyGkuCWFaJIFDYrMan6m5
RR2Qel6QiC1mPVrLtzDu9VP2fmITOVQCPoqPBDjkqVV2719WDBLwAo2Mgjf7kVtQM30TZd6Hk+aS
AL6Atn1+eewNIAnpAlhiwcFKAcPpFjKr0crInwQjccieVmn1LR9EIAoGzIn6pBKNBvyGZBBQ9d3D
2Y5mndS2OZEv0yZ68qJgsv29j46WEqObUuw2kwFAMy8rsgWKPFhLlwMAeLafQItkzyt8gykwQtL6
lIsPBNYpD0vdM/TuYrry6/9n3mAZwyRYXgmQ6zKQYbLbENwyRLHyh8WA0PqPUaee6gz1k8wZ26EP
UuCe7A0p3lGXEe1pc/vKvyJuqM5eXKtcdrVqbsobDQ9PnqeiO9E3pvtZ0z9JaLfwLgYcz6ePfAYK
iIkPTCq+FPZ+F8YWY6bycFj6lC4oKqH1YYy8S+NpQ49uA4npH32Gk4YXYVd8Qzzdgc7qME3+jdfH
DEQOw4YhZ8zUep2DMwzhPNCgJIY3N1BcqljBSDeYVUAzgQLYc4BkXMawOplD8R4OqQ5dzvRaDomj
BUjxtTs601H+Q4u+YSgeq614rSvSfN07B9eyxgWxwJdAqlonBhH0/lZqIfqpncnK1GzdjjkDbZDK
ON6GCcQ4gnjow5B0RAIAdP8RLVmgJX0T8XG4myUTJHYrbq0k97uPW385dJicmHs38yBAoYmJYyKh
/ftID8giXTP8dMkHHlHSBLNZRKNPz5mnl6fc0cmU3N2VdhJzM9PqkGkNEoraz5NLIOPN/7Bv25hH
YHGw7E03+f0LodR2zQAbFM5Ihme+JhXr+aul44AVGCb290godJUqiVe1w3cx270m2uIPqjffIrR9
/sANMJyG8R/W303UQGCj5hRihWJzpOf9CujwltaGf1YVGOXIm122ASijEFG210ayFgBSn8JFNLZL
1WWYIGuTkM6hVFL2PZxJH90qZnd1rOBQ56r90yiSNQqUDQ/oMGcVbfLTprcM42lq1ubHQgf5Upeu
5x5OiSdWJ9E5JqE2jeiNc0Q0eM1cL4YHgi0X9oB4fJI5LBt0VvZyDBJC3HzApjNF8oTk0EXpszlS
0W+HakmDZUJSa/3ejG9ooEXi3MBTfXxIlMP4f8C2lStexR903N1f1KTYoWCqvUtFvtJQ4HyobW/G
d4O9KEV5/rpbhcMjzelzJVM6pku1WTy/mwOj68Lic07ffLWjK7zAbdVwieXqtV58aIwlpHKGq/bN
8XNWGN4oKPQ1eIkzJ/QkaSB4yUnEqmynsHJTy08BnxJxShkTH0+fXNn01APrqvXbFV7A+hCqz3/8
sKva0AfOcVWo9mDk8JWaQz5/8WQRK24Bhu0VmGu1PsiPVUA6FOUaQhRx2MMRrFnWObwwsVx6H0il
nPtRy57OeaIZ+RawO4aaASPMGIpka4idzTFBHXwRjuhkU3+MLZ/Jfk+89JB070VpCEYv/MfrFG6G
eDiAOhlWRqKOKzaXdExQBuZ5+rtZ3QQ6Kjuk7VFHmJcYnbtDqkV0GxCeuGc5Mga6SlMeM8vFs0Y3
swzIfm0lcneqriWjqV9lopsqlNHnuSSBz0rm5KpprfTwacJoEbfbGRrSgGftdafqdB03axA9tbAU
4S3XVLvlmZuk4GXocmCX6uDn2Z0MNKq4Ie5ahTBs4exYMlMcmflUNQ0seRyOWgDH5GU6AacUj4xJ
Nax9zCOoqfJGm6P12vNtXwDANj9TNFmpqllcR10sx6PmiRjETkg7tfSEaFimr3nKcEnuq8M+bibf
y4H11RxWjpOn8Uj44BkkV8h4pomdRre9OZTwYfBLvZTfJIlVcEB3fVAApI1/mbawajRP5lVud9i6
ljBPZfA2bq9ldoj0P4qjMlHMFxoPgzoT9w7stw/Lx8nWvdjkH5j2JG75nf3iDeDjpjbJYaXJ/KyT
Jt7xOq58YJU2pcLjKnhmZwTdRAF+xHkYy+neumHgVX/OEOb3kYfnr3zfA2x4ZABf
`protect end_protected

