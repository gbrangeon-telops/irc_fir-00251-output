

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HUpwfbtoJu5ljZH1PD1nirfZUiqEH4rdOJmHG3byOsiHMKK3LegkCLnxPuPlk+MO+z4ctY9AQVS+
qDXnVNabAA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J5amwDwAOhmwY1AI7aPhS8ck8cUzk3ZbW/PSkoxcoFtS5AuFiIpCT9Eh2Lt0JzHUUKx72jQhC4xP
E8DYUPCIo40JuI++9z5fK4HwpQiCOB47OP9CCbDUXkdRdGgF4e6aIOfD40xCprloxnLZWVs0yawE
2eWpDksVPZ7exWV5yp8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kHeSBUaR4Gb9xyNR7/PmBoZ6gckk9p1h7+VOSSxhgJTOkeDKrcZOdIV1GDgFDrDQ7kzRgTiYYdNg
fXk4UhiKwBVyrTjV2sMzg3+WqoUQIK6Jy3j+rnKZ0FHbaJ/B0H/GfbBoAdHe7Ll2JvXvA2JrUnjB
cZCpVeHDgAOSHC+pzlRSIpPSacSQtQcR7XQ/3XaxnZYRC7uHkv276AbG3wIpLBG2zxIX3ZP+ackQ
pH7/JslwJLo+2yMp03WDL60KY4dKN4/3Cbuq0p9ZXqs2Y5D7OEUZNxyvOtt0dnCx89ZP9OSkU6+U
STforoN1MyOGgJ2YZ3QN/z5I0fk2RYpfEM9JsA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lu2s7AKqknRcUE5f3UmM0sxhb8YGklEChkrpjNpqeFmWrHZVTV653SjxOWSucZRxKRWERgvAD5Ge
f+lfXprxLknFOXVThhIZcoGHsP1dAaIYcRFINHuR+NXvmYc17FBsIljnkMKM4grLGNoBCK5BU3oj
+OpUaEAqYZcR3Ny7rME=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZNNygMQdh+aYmFNm+RRdz6IwBodkqsu7V9fE3BGXF5I2MBgRK6iGinaX8yLwnKR/gy2F4SnWUzqm
SM6Hy+mVD8IIS+xm7ukIVwLbM9+0zez0kJn+qWOW6DSjxPXqHRWy3fQI42FtwyVBs6pb7/W8Q9NM
y83XMjmhW9gbYNHIHq5e9D7ao/9WQ1Ytg4YhUY4H4cSzY2tHj3tbIsVO5Swzs3K1mz8KunAK9qzN
WNyQE7ctUOauX1bPhyKN8vZcKzkl7x8jPe9GO6BDBcCZS9DeY3P2LTqajNPbMa7b+rdlszJkVZWF
aXg8+G+Fp5cfd6qUK77FET8A+G+lv6qs6bNgOw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26160)
`protect data_block
LvDmGX/FbOMJdqDzKgNLPIbBjXy0f57CaSpJ6zyR3i4mkwvyBMbpIpufy8/h50Hcx6ZIdGeFLdR8
Jan9SXZqYrk1gcaMgE03anRaxOLGXxPc8K0BGupIU1c/L03sJI9Peae2f42FqvhmW5RNQ31b9LTB
gnnS5NXpGPUdIbsIXpPdtuEWyivqUh6a/J3BEcrJj3svtW0xNkCfZUZx6CY6c7d0GejXxMLs6XqI
PoAR2fT2mNz947tKlIM1kxl0AtDO4wR+zCATRv7bYhIUc0Idjxjr19gXxepJ2BWeIfH5F0pJY+2W
tyfj3eDTUuyzz9AJewOTB1qqhaieKhSjC32tbrariit8/QOThecOSVLAZEAFYPbymLqSk5EBQxSv
bblm8aPGj69tR16N+2eQhAEGyapqu35XOv563O5iO4MOkcurlNDq7cE5t4bPUbfLjq6ZyleSmLP6
QDWoOHdXNLWXR/j9jsfmnQyAO2eHsX7+avtidEUrKWlDX06TrCBvxuAKGZY+qwBPzUwTENFvnIog
765uRiv2QyI7QH+ZkbNTV6BD4PpzwEZGk+d8RV41OWX8QZ+AuG1aHn8K+8tezfAY4eCxpyIsYoRO
7iSG2WlQqO14AXXf9SkpkvV7kiULDpE9JxXYMGeed8vT2CZhxyUkbz3al+dxtbAdjJ91FpdVevCb
8yuoXbsHt7b9vgVnV0i8uA+dxCQ9J+U/NoVjH921v1GpeWmeaTA93BV2ZLnwyq7r+V+DFtzU7zDO
I7MaUOduG1Gp407r9q3YKl5QU5y7MkW7828AqUf4hh5Pw8NBuJjGvCURh9OiJgJO7PI+GmqUY01a
LGGIZlWADwmIkDlvklHEZnhvuEjDlYGaoccAvxoQQZSam4rZIklY0fLoY6ALSfWd4pFSZovKZpDN
hL4L9mrX3esbzquGhrGYd9Y9rwpoR+bI4dhu7oZC+hhxw5eX7DjugtvjsChOCFD+E2vUXND4y/j3
N2yTD+gkzgyZal4K68SL5M0TBK2RHi2bxidIUWP+zknSt4zswOFX2cpmCeZ+OL40EwwmdqQ5S3j4
BbwTCux+PFTkco9elLRW1c9GO1nIsTmck6ZxsheYqDTkfJu2zsu6TvR7qcOZ0MgwZD5AZoajr2/h
qJLPjMIRB7dsnSqgNlUG3LQbE8S+iv5rOE/WEGe7ct63YvsjX98hA54uvDxwk1TkAL3u1NfH+Na2
KDtP+MS0iw7drZIohNu4HSVZWJaqVeoofbJmykgYpkTOpuDGvPM7ByJT+RPilB3YMCCxYPB5k7cE
TeDeVS7kFUSV2rSCkIYuugHj9hVcWFo6dacWWwkXfTjuZVmf36YcUJC5U2y9YFMLBDN+aG12mvxJ
AASGwAHz0BlAoZ30PleHXuzLxySwvq8FO4Bajrv+DAVyG2Tl2SliUULMeY7aHF51y+mJvYMy1CGk
jRNRmTEYghNTZejN3TJAGy02RMR1YodeKElssrIY7sbnkXI8oTb+HcsObWJs/WBQa6xmdIDBLiFa
xdRk6qIFqBhEbmIW7btUE+VDcw6OhRi7k/nH/SJsEo0Lq/1dcXxpFRhetqYtr29eF2ILTKKQLlJ+
1EG3IAY5Bhy3SAd5HTNro1SEgpBHVG+l5/WT9I9sqV/3y0RJGqm/AE8YrfCdikxvoReRSsZh/JZm
GWs5DZGJ1qPUV8U0lG3l0NYjqcs1mER7Moix27M+1ng+yYVxIrKQgzpJDY13AutDf3m6bMIQncJ6
S9Rx6J+cs2KIU8aOtdkm1i8ai5jWYhZqPSye40ZsxKOTW8J3PFAls6JLHtnJ5tcnt33EkPT24T0I
IBLwCXQmRCemYO5RbKoP4BIzNsD7lni7bVP4w7xvbDRGgFumLMR/Ird7P7NO+ib4EBr+ug1L49vV
F2F7WmPBNVC1vz2ZAkscGSCi/9n8e47tPwi9Qx7TFNqdlA8nRmWbwREMxbwp0d8dpUPUQTGRSM2V
g6lomktKHbem2JvGLFbh6chpFw8PsiHCojhz3dQDMqqZbolk6tjHV/pQvVYBTIBHIDoCCCSLU27R
QGyxRwWFA8/tDkGMSF6/SGbkSwnookaaP62RJWKjmKg8Pc+PZ35ErCm6efdzQ7P61PzhVtSp9Ytq
2LpJFOzw0HO40luI2Ycp9tZWUuLRwrgZisjoFZTt1MRWP8FVKn5nXE/Zu/uoaMVU6aTKFxdHOdGC
dRVSXCdqvipzwIo6sVl6Bth1DZIvePHP34ph61OLI7uXp2jfnCtN/zJ+FgkJHvI+KujCXRmuxhcP
l041N56qyPrrCtPrNIi2a67Miz3yBFf7wyY0wOUFKIio1j2pFW1jWIDOPOzOyfkVvUGNOxyko4qj
21CPduUyCmb9sGeCOwVvVwGUYECgi3fUmxvmZu/ZQ/aWQAUpMYNRPT+sVeSAZxjdAmzJsQt265oK
JIS5ldJsrCrAX7Bd+sqZSihrYbWx+OqoNEqVN3D5CJWqaGv3ew8KKFDK1LAwEdw2y7NdgWmwabXU
b/nUWjmz2aJ/f/H63yoL13YqxIRjWbkfJZvJQYxqX8Nl6u3p6G5gZ923Kor78hsvXfwJltJ9XwmN
MqFOQbtDNrJw9XHQy3nv3770Q10o3ledo8bRKF/nTC7YsO3XsVdaPgc+QgDegVFXTC452GNBNVE7
l3kp/RWiwDODpN7TmtBDITzF7KY9J1RhG7prGKGGr5DzapNMO3qTWzF5JIySx3447VXIX0NDd+qR
VisU9XEBqg6mBBcx7ECtPC9cciBX3MXZJl4a6E6a2ZBgWUxfO/z5zAdjnN4gI9YzOEqFO8c6XU/S
pUZFqdgY8KY2Mde9AIvSswKxJdArz6SD+1bVNLRnoejxAtCYeC7GXPvn1Xz5FKAkOJcBdPNirYFu
sNRAHkRE+DtMQLV1TEKrcgIHGCT9y5NubSv9p1VgeyvIbSfm6ZjnhFuPcUTiNkksZT639VheRcxH
CM5lEfKVEgxxkkMO0IckZoFlWQerW3DgvKPSvwPmz3Yv/nAunONTy5Qz9uvNNGatXcssajKBgJAx
8JfNtXp26HW/HPlMjKlDbKEiYk8rmhZ0/EEduxlqh+GtKebf+n06RmkSpKADmlShm/Uk2E/xOAh7
LvGPnzUn8ZdpXXxS0FQBfqaBx9Ds7nd6DW3YBzO/Nu5BszCg7e7BEjGzCgMXBdlZl68ibvEFFo/G
3z+Wj1nKITM1+ny8/c9EHD8IHor7F1AIHj/kjJzCvvQ4ZCWjXEW7scjZ07VZSXqAKjS/GydIo+on
LJszxuBx/fH5U4DrdyI08XE1CRF7U8qb74GPWsOTGEcXV0koePPL9+7G43aqW2/kgLdCzUJgzRSO
fFk912JcwPLMXNnH6vkwnan8uT/4fn3scJ++kPl8Macps3JsptL6dz72oKzL6sxT/PNTpWLFSASd
X9FpnWfruBzM3qzpvGHUOYimxltEahx5RLyQmDHelKoAeyDefShc7RD58P905WsKjM4waBPgdO3u
oDUzuibObAn/iF7R588vbs3vyN8hLksFyCq5dLy2gM8hLHJlayk9X3oNyOUUio71kA57THzLNeqM
foyJQ3tm2Uqt+EkMtwCKWNDl5kR1oWSEJxEhgAbt9ocBocIxV9w2SW3L3Vwq+8GVrvRjU1md0ah0
jqrd9DPX4m6ovU77YCuj6CZhmbv5j2FZqmucHmZm7L0DRCwa24Q+7mS3D+1ulsItLlDQQcpHBnm3
UrBoaakAyFznnkM5lMNvFmjziRlGq4DKhdahAoIELalsOlpfmSKNOoHuLLNls1+BHernUVTT5wRi
QGF0GY0YCAIslEofct/X/xb6AdBrqGqLA5Ax/+VqzP58XNwd71tydi3u38M5kmotH9xdDhDmynoo
6O1BtnIoUR+wJajgZawKJ3kY0FWPUR1YXQk/82xsDRJ01h1/MJv2ZjBmTQz8uFlXbBS5VO/nVfgY
7LpRmOFvO15HKfmf5I7OfyBOJMr5EnH7HAqVeH3g0J0CRbJqdyTf52gSO3jnxZCh8ezNOzCOH/L+
lJ6bcolmQBQUt3XKw1/0MtVZIaPJQZYcp6SScku6mVRbqT9OwQVYfi+5uta7fC1wdk3zQ/yG3g4S
unY64/1N3rYSgN8z7k6C7uLz92oaD0a11Xzg94ksi6bzhj4AQHTj1kVxeAYFERHUQZRXD201Ckwg
sRTImDN5nu/m2iJshORm+8iJNUNk2P9VY5u6sapOPG5FV0BKau0El1wC5Vp/2qCjnAADN7yGgpLZ
lfUNHIXNYoMwKx99ZNquWYNAgBzzJhUbieJEmjTUhxgcGabYB+FizbiFz+OE/oUOJJKXqxTuQYVs
LiDTTktXFsYBiKATwuPo1efnQRxsmC7PMvrEzZ4kHGzuc+zGiNITlQqIHgxd0MEKvqxhbuNYHUtH
EVBj9+QxA8fgiAkmDeoIykh/IrrpmEIfQjfEQTdFtXUjatOlyIivlzT9Vqj19qgiFs1BI9ZAzGQU
LVUExJAqui8qnZNQgHgHWN6YLR8xjSooqCQmkV6SBzb7VFcG51qJCBcJUnbR67TbHV3RCJ38wrIE
jImd7k50yPWWoVvpAOp1EL0nOAQeR4RBevmigcdm+rSzA9ZJpiXXWqCc8SCL0Zd8azBhZEN0Otet
MbUSiOoQRjwnKEiQ2l2lwOgSDi3vuIqFoMqMxcnoYW+MGE8ObIiW9DD0/dzvpL/iT791f9p3gX/h
0Fxn8eSvsGHPSqHlatd7A3ZBCZ/Y2M1AZcoe+C8HkS+4hdQhFA4caOPD26sleq3OWKhbLFI9jI+g
MPgI6WBfGa9xX29BUWZO1kMzbtgiP6IbHwvj9E1oW7p7vknbqRM4gisTlifW8ZuembaBAfZ23Odv
zZwB32OuQoY0WSFoTHfOQUwp1kMFlfCdXNnrUY8DtSPI7+LvLnr38aNkQIkHd0Yz8ckVndkOKM42
8OLVW2UU5oQOryk0sboJJvbgbqRc+tP3WreaQGyKsBaU2F9+A41ya7sALvr1fTnIUKpRGGKKm1iO
/56gi0hP65F1wB+c7FNb0XobyTU20ITIeRWI4cCOUQ3gWRM8LmUoPdxiAIsJUEhdEN/uzCOIunca
Iw7l1JdKgGLoT+WpWa3p/fvsR4mhmA4kwgniA4VAcJSwNWN4pl2iX5sXpZh3Mwx+CiZNbgglpAdn
4eq0O11984VUl+R99gK2ZE9jP8rrir3kxQ5vh2IQ9O376VDD17vJDedw0c0tRYaLMEY+yC49OUJF
fVyZPEBFOAUZSOvWzyqRzqmmzY3cq8kunsdWzp7iyPle4OQNmghqighaiu/fC4h3T9VrUc/w76Iq
xDhXjqm3Wf6RBTRp41YWfBfNKCvt6mv3+5ZlcY8yRW+a3noP2zpXmRw7EcqeYxfzdv3U3qqIdxTm
qoOiNfxEbwvZnkH/OSumIou+faKhIhFceGQKOXhzmYEtPhICOhUjlrdSEXCZvtOpyOOEXeMNUywH
upRfFTr83YxRvf0GiFOJ0nwePvaP74pv5D6WK57BwfDNy67xr3++zsZIl4gp50yLE3BOsTInM+Hs
drsw+Ovx/s1f9JAZJFCeELQlg1T69me/c8ak9b4HhK79fofhziANf/cFybT/4Qu+n2ufzJ+VMNl8
4ZuW/sOBss20boxESq8nz9qns89FG2R8eoH71CWtpzwAJPuN1f/2WL4rmsIUavHbkoajSXIs0kbA
wmzRVGUuYFxdQ5AGbDPhAuPR03zB7zuj1vTAZ1NtrrdwCWJ6P/zupynJh+Gl7zBHb7xaEhO4ReBA
FIwNsEdp9DYCY9moP2oszZckAq1jiLiwWQ8CNvDLklcupz3GMAHMaNnzAntfRGlLnrIZT+woU8/A
3fTaux3bxx603OXrVv+0VPNnRQaW+VMW0mrfbw7Mqzcx5DNVfk8biJVJmyDOr4E1moaLeicIhM9k
DXl7kmAFKXVgoL3aAwZNRK5VJBIWsLFV1hodyCz0HeZ0bOosGUNsfL1au0ovWtNVrgbLBwsDYQFp
NqZn3Afwz0Gndj3fanJRYCCgIf6fneQCi00oBMRQN1JXa4rIdn/VC7fodboZTRoCv9/n224ZtxOu
zEIa8E/O6XcnKH866r2k0zAYLspiCyQjTykSiyDuUlL3c1cNhNzQTu8fe1XBcK4JeMuPQUyR+EkA
GGrWm7iWpQcQoew1ym3rJQS7kqtMB+GnHUv0T1UrLuwCHnIqkMEK63deraQxSfthaKXilHbKxS5m
XYoIsh+4+0wZodFgBFDRyPSOaIgh9NRiZjLrVxS3Afn8tv5CbQTJkzPl+celMugVu/bTPNPTaJfa
DJmMa1jFQNyDlfKzWeM/a0Rf95CgLJu3NxCtP+hVpjr9DUQhtFpmncIAho1XY0RukBDVvB7DD8jE
MSqzGRGAwiU5vWKpFPuZx0sVUhELExKhTWUQzPvqyZzdqTq1HRJfM4tic1uSSvZ6shV3iypFK2DZ
olXGvGhT/LPgBmuMEAWMhkB+JIxj0fMiX9h/i2ewmoyGu5WIF3lok7vpLGww3q12hrdErgDHT9su
1i+SOW/k2gsooC68GxcJ5KVzxfXsTxNevL+MlbH6NpAeHJnhbmvtigMAYRCv/wurYF+RJ78cJ8B9
JbFPlw89rx3T+dZRRqzV9cUf0EOoVxJ/RQ16DyEKuO6hKQCjf2tz6xienGUZ8qsy5w+FhOM6foJV
D6E2N2+e9JSrPjv8JudHB0s2Dk3oym027Ta++bTBenIO9H/x+EyhIaMtCDEomc3qy1N0ALvdCWbU
XdJQxRXUrKtj8CRWx9pysVCPD/Jjv0cbIyuWlOsIAHqyZU9KF7jmr+O5LwFZ8IsOdtL0xaN9QlOZ
ZiklclT8fS2qsKeG9W/nEMgMoiS0bOol2wQh47YZ0wLHz+oMs/+lMlmbOtHow90y2Oocfo5mwljD
dv2QdeXG7iSUIEZ0keKuExY9WeN+VzlkWVeVYR0e72aprOBfq4tnlHl4Auj34yv35vq+FpdCiq+e
13qUym8InzJIiZPoOzfnsQgk8WoSE4PELV3ojYruqDdaHvXi017t8uUAr7kRh+MuUxrWb63fbHcT
AHAChsRSklhUgbkBED1Fd0n7+k+g7xi/7yRNWgnTbABqIGTJyX7WqAy6097WqeeJzBhDKsTXwWPr
9xBsyUTDspODr53CjesbUyp2RAmlwjX/AkOzWpvLYkBJNwL+r4QDLSxzlMueZVjWPcL6cuHlLfD3
nxpR+a/TLKruCamwhqkOA6segi+U9j8fmJmsSeqUQPcmBnmLiQ2sQjVrr21S/2wTLO4ts8H8pKqP
4d2rAA4egmiSs0ccko4qGGzEK07wfRE5FiebnYbO40TlYJQin0wmM/nM1+xPRXm2TBwQoYxlsVQf
EbHJk4WHyrPD0Q3skKvYjs7U2/X9hZSThxArHCaT3rNuO+AJp1pcNBM9qj5T6WreGhDUZEezezZu
U4hsu8ryuv7uctrbluuEHZxkTHEvT6mID7CNKupDZJ19+0wOWyrINIv7otufplfd3PxVulHK+QaH
vwld6l1YZxTh891qwKn6Q5kfM4tbKa4nWDWKLcJpL0jgTG3pU77oMTpi8+L2q2YL5Gp2vVBamrW+
zxsd3/p8v1a0AVatnXMmtrE6Q5MhYsDC1PQs5FLD4Q+JDT6PXn0+IJQoeQH49due5pP8fT4tU0f+
/VWmXIaxYNIcUh5yeGuL6BJXJFj/cqsiWQqD0JxHtmSJyUfqgWe6qAxghTevG/puv+mBaPiAb7bR
6z/KU+PvJZC/uMJG5I8VmAL5KLCp5Juh/d6pKZaOy688m+3tYez6ohVCJCuyd1gZCgph6dr+aqrk
Fzn7Gex2uPAjAeDIf727xryeRzg2OUAdi2wgLi6z94Gphga04yudnYt4ebxD/hT/5z2vkhzkyXSr
b0CIWW2azMocleS8FXp3r0wVDIGyR9r/REplVxJGqlmWhPsUT/oPa5Kh5KnRtZUV7UrxfzRYicc7
h6DaAm+NGsoG02+W9YpTLV7pacd64cq4vKrUQui8wLQkckMGZKOFoe1ZKku9WH4rRhBWkApaSyvG
oeck5orU/ooLJ2CmtIKojcv91H6uMcPGWZQ7PlzexgfnN8RJ3b6JuRytDqXSkhYBJ595YUWOzvfw
GuVvezXFbNtNA1KHri7wDv+23DbXT/mE5qFFZEFlKKpr/TROMnKw36WDwc9G1exG3irXOK316RdD
73CYYjFFIM5RqLLjxTOPF6o3y74V6BLEgCNST+AvLOarAVOVeK/2RKCeHsEN68FT0rjgCM5KizoM
FuH+AnuEBzdSOjQ+ns51A0Mtk3j+so/e1h5KncdldBcYlYtHk1LlJii/+I/Rf3GHjFrXyOHBcRfw
pfbz12JMx+8f91SX/qJUfD/ZfGTq4Q9gmG151Pdh2CxcSfQfvcqq0UFlpU+Adn5EPAqG/qqNu7LL
Nk/kpu/v3kMCT27UrtgX8cbTaQj6Wnm+n6G7RuC8IZQSyAZLJxUrbWYH7kjKA/RDwy8Hjzqg/0yb
55rO2CE+7szgLGGiv/mceClGqo55JBhOIKZw0llCWvmCofl58NTcqueVxB7XO37Y+LF7QTgaXipY
SusceP4LfYZ14xt5OjJQYrXYpzqA1ju0HHv3LT82VLYRGnClcVrZbCy3YqbXlyk5Fen8VfA3O3gw
TRkGLXAqpoWGL8PuR3Y16YB+H16lkdU7SYXG4dwyscJBfuYsNpTD0ITNP+2cTmu0BqEwety4wizz
tz2mapHPuxYmayPoeFUIuGSo0ZmRgPrVm8ro1ehhdd2wbttHE76kgoL03h86FLZDHkVPgl6Wwxdh
0ZP7Wkr7VBam/PFFhHE9kWzPqAd6KRL4xo27zU9ducYlBhO8WM3clRBohjwOqQPdyurfWwYTwIgI
eMJb5jpBPt0vcgojWazvo5ITCSEJZemj4IOpHaG1DST5YCUjOYSIhZLw4dWalpJwCXIo1HHLa4JR
TT20RjDR8+Ge9OR2lvoKmZ1ImFvx7TIgN54VyLMjEZHItCCbVN3VIuxMjmVzaUX4YFOHPeh4GJB6
FOq+YthD+UlXbiCldPVd2m/1M42jHZaYNSYceREQENgVOep5BvdmjP44aNux1Qwifnwt+boOJIna
atmIIMWUWKirM/mpRCIMLBr2OkxWhka9Vopn+6utaeXhSTjCnXurh3z5aaOcKoNYtB4ptybGOKuo
8QC4KK7Ioy4eKDqS9HXw2Mln5QNpEybUT8OuUJFuePrNw+tpduVzTs6CQ2BZLUTI9uvZ7misRGj2
o/9n9Zy1/acJtZX3w95Tw0qAodUP6nbDacvGMDZhJCGAJUNKLBPvTMHfz1vzoeVACbJjA8oR5put
Lt8cm7+feSUyHzPUwFJ7Llvcc7p2FGUGIWmtd9xf8jIdsg8J3fHXt2d4/te4bv8aipfwbCJ2Zod1
46nMN3bEWPy6dEO6zUUsbl3g5XzmeEg0Hm9FxHqzUgkbgVcXGU/Y0qle0JuE1Ne7BSYU1UdeE81H
IFsZGbpslv242jYFcqEMnx/brYW1iIa2bil6Ykgvle+V+s/zO/+W8ap6tOUsd2horxZDeuUEI8nd
PJY4J1WUQPcavktmTkbl9VVAHDkLT0/Cljk3slr2ZfUpxFB7LxEDuBWxbYFdQ1a+oLnezK/tguXn
dIUZoNFQyim2eQqFVSpf6layKeQitsTp0v/A2NjqLsnbLqXXFA4YFPIoe3idQzZuHUKLpLEB3W79
oe1SMHsd4w0fYgQgrnnVK+u6y5YsLgJa0q+xjwLZRJfmO5bodP5mMU7Cb9pWkFPsEpdrRFSRjw++
H+AIO73ks8p3BJDabUCswqlYZaIvMVU+zuBGkFWPOrVEYlGn+QYDrDc+rb9AOvtLJ2aSsoMwnQM2
656xSJraxo/17uosLBxKv1Xel4kE3qDNq9MNZgFNo+n+Fdo/KqfnTE4Byw71CnKJAQGH6x8ierPS
4jCbjUfk3CJKDwIpeKcAhFUkx/WUU0gtUq3tEcC4XmweZJ+fVbX94Smkeg5SdKVcY1MeaFYFvOTy
0b3FiFC/Rn9GAQEa8dZ9ZQor9xmaaGBbhPj0Dpjg4rsq1kIyGBI7oUIxc1YIs8FnhWJS/07lIeRs
YzoQYdaKwPQxfLlKyYlc9HbumHH3tpI28wDj4OmQ45jaHzSej17MJ5vxqvleXUkqkKXL+Cpzep5Q
vm4RGnBY0IjKM4ph6h6k3A9Krcwxp43d3ipjfwf2exr9U5r3VQnTLjjpWUNMUfy1xlswQlCWmg+P
nzEJ6uJ/4uw9fTrQ1ORu4EaoRIT1JkV7ZbvZNv5suBal/n6UuP7Q/H0NDSLAHXPj0Yi2shISGPM5
sk1teFm3jWEOig0qVHn7XDkBoShZf9IiVp2LP4QIlEZhnX0zuHDxQUrc4W8PeOhxmTCzAq/ELenC
K8vcvqih0zRXCnq4k7HO6VRfV5eR0aylbh0peqlhVQH8lh6yxh21Mkw0D0GUK1TxK2BN8xtmTECN
U7FrWvtckobJfHcVaYsvcYL77vfKnhInYvZXRM836SA879Ltx5rqlllZNjCBIh+4ajqpENBmnLpE
dZqvVBUsqe5xHTkcqbsLF4Reu96jhZPxlVOjUhubFi7x1OQQ6xGHppLfbMUwEd8knayBjtXDFpZE
hgadsOH1HxXLCtH2VE15Jlg4/mbeER5EUhzUGF4berx9TeG4ZJeNLixfyAxoF1D6voe91nS5g2mO
yzHAoqnYahGJpLj6FwCGVRqlE+y510R37aDKIGF58c3/yD//6OAszpngf7bARFKpUzSezZmwuAl1
XfTcgHs5niO07jkfDuMj9ad+/OqGfSwJ7CCXDTBsdqPDWdYEJsHFKamH12pE/LbvFktqe1uEBhd6
cCiiKOcRWCKANClE441SOyUeo7DsNWhBCbxTd2Ok7FN+XhcD895EgEat/EsFeaSiZ/HD2PtOIFjP
ssc6Lu1ovAoARzFaaHDkcbKGxuN9K7GVbWAMhspcAmXZKgom2a7InXxnL1fslJO4nIVscX65znfU
XuCgIULV6uc/IEUeiELQyfq2Rpo/41F6W+uzsGJ5mpDWJqXwYvgWopbNrCIDkR1qtCqz0ke4iQIN
nSZ6ZsMX9femWE7y09Ob56Cw7A0IM+vS+QQxX/goJO328m+fKegFD9ohI7nMW+Jq/EfUEIXvcSQ3
YjLxbikuH2Lz/KFIcYT4LRTMhZoVnn4fva1iRMRu6CHZu7kMMeRYhZbG2/FFzsEd9JsWkyRzniMX
RZweKPPqyVK1MLPilhveJcviQ+5ZVdAjdSFMIWWATRJNmUsbxGIMkzOQZoMjzExQz0GLfmqx0pAy
e4jKdrkenp76gbH9vLoOuiaKQSqxTxpA1NN/Q9BHtbJg4N6vvhEB2t7cxOLmPPMvUMaXfOoyJc/Z
jDFZuZtbylPdMqUk2XTYRG/8HfBcIDRxl11JuAcqaqlA4W34bo7lQP78h6CA1CAwwbfvbS7z55ij
Q+ySpA7k79VwMzm7lKHEeqd6kUo6e5fcmxp3VEMmgn+sAyIuuH9xCbnRxfeU7iE3D2mrG1roq9K+
NNbRxu0bbtPjHMyu6TEm8fhh66De/ZiXzjAKDCX7WEOnajQimtIrN4aC8+eiw0J5PsZwWiIvz7to
/32c66LppBhFnw1gd9YWxTBImh4jbzpd/e16tiI0k+NUKd36pCsi/zjKWKGRYIdNvCY58rYsxUko
Rb8czgKFikPEGDnjeAFHoJ6xTGKv78PybR4K4eKcpIpY+LPw5hRDODb3m6leCs4ORTQxGJ+VWZav
IOgqNoDtEE4Njck0pSY09RbA5/wQYtzYx23+VXp8a9/hHP04NnsIuAK81pnlDAA6CGdp/4nEW05Z
m24Tn+CoagEUr02zF6IB73I8Q7iecLil444K1N4SjJMbwbzROoR5f1610qZRJ1LOsTrXZHaV3j6T
taiWPUd/IuLMz1MWuDUSjwbbyKGKxFQWMtzayHT9DSGT7IQNzOgT1rNl+BtzrevdgHUZVAnHh9Ey
aTYVrS2HdRucWc9vXeSezwfZthpK5rjcZ9GhwBVUpaDdK91tGEVQUQIQX6AfXs9FxTExEkfsLl91
RpSHq4FgxyzzjRT7qH2hU4nQBAUxdBc6rlvB5k6CQCjZL0+Wriq249H/y90dzockinCgQ5+3WWtR
CDOi+F6ZZ+jw4IYhXPCUlkuipkYeq9Lee0Q51h2ny+1GIzXi4FCCS7oPpak6RUv11F3oERNbkNrG
o/DErmWvUAWMZvjRtVV33TNF/0vJj9Coujgqq/dbihcRzfVqhLcm3PtVnf8Y9Lgw1aeZ7Df1BwEN
RR7Mi7YznR0vLL21WX6UwWA0g+q3zwYuDcQ6d4LxTD8S0YOKpDnMQmLhQuf5guipBxd0FWjYXv8J
Z+DoH/IA8qC1uS9lN3l4AqVsvIlXCrsNk1uSbCnGvTVt/ifMyQKem0mTy5Lz866Lx/YxFIA48GBN
DH3TEoet9pKKuE7iRQSfkN5QyCeZkwyA52grxDex/MMMZGwtkPcOTlx+Lhi9gClzxCq+WZGg9LZM
JL8B7WmNLfknZkcq1u7IRiRxPQKTjDvKZkuH02Op76FZ4UhT82W6lKOV7ZJmDBFqlrkBzWATEvGY
SXgP/1Ho9AxuX2nmMZSO0OGmGa7BKMxdD6IC7fZpXdjRy4HHkvvdbbX0JfKKPuUE8VTRLi9J6gPF
YanM0j1MaIHCXHG0rZf6PdVbhLPi+HX4U8wy3KFIHfkeJxmPT13WnXdBa9ATbAsiPdKQ226FYNeI
32nCPwoz3DN5irHET7/jfjQxgdlYV0iPO4PYezCCbJRX9P3ccmdP28PzWHyQZzvgNZvEvckkqucK
TXw+DETWQsHYC9QDdoJ15DhqNUE5ndMht7SoD6W8ZUX6wZ7W70nqX0PuVcyRJAVwgjiU2QNFeQZy
sWgWvTtf3wz3jH+GTeed6JGK1xrF7+95n1ejHLi+yoidGGV1aK3LAxmDnTBkumOwixs8gb1hux9J
EQEzarueV1I9HaXAZOXviB9eYEJ+jjfZJQsz4kYE2KYxoHDQnrrE3y/gdihpwbEPsqDcq26Q4kyG
VzenJ4q9i9VLXWjFh0mrKGMzAvSBHulKwNFoe3czv2CCRWXTwU/ZvigDjGPHyz9cz72nGHCGWYTZ
OeDkgJ+ZHJHstm+ZZy0qgPnl/94qnkB32C6I3Rh2lgg0gNApG5VG7Lai3fNajcbAx/e5r3LEz+th
kOcxQCDoKdS2IgWm5E2wm+Dwhiq7LfzrlLeOOefFOxaImEZl+btx8ynN8o5YKAMDwznIeuanz944
82hr3eIOKZuM3Iyitj6nbR9Sgs0nGqUCBUPeWCJZdm2VqPssbWiTWL536RJSY/2hlomz5qP8E2IX
84sf+v8KKUuE1d3KVuRJYO5CKDXTR3YE/MnvQdwRH+1dbcoTsNyIOVC5ZKvDGJawcPfbSbt3FKcl
ry0c3xwVygo5HLV7ZqSl0cYKg+h9TuMirNLlqGfs6h0jnFxE7HkDsHiXuxP6nu3rbqutafGYyVq1
Gku+yfSRGucBOClcEO34xsr+R1x+G6jUNwzsuAW3T41Ybjvg7UhY50eZKMyKVTNACVIDz/gPoA8j
XO3YqrhwjHBJKbluPu5Ux8wlDKQu6ZiCjM9a5jfrn/fT3ojYGu5BdFWDD5M60EuMy5qilxDR2Vyn
vXPzufa04dtpEBzei8PRm6lrCBAlm0+BLzFCoC2+0dt3tAOlLz1u3SSlvSYnHM9w+qw3sgFmCLza
vlTdGiS65dyI9jVrCvvKALycbHD2NtBvB2/8qXP9++u1umSaCmzut+RJEXGY6uThEzqtGJNAZc8l
lr2lUs0qeSf+NXL91QI8fVT0jroXu2ixpkV65criZZQo2zzoAqIh9YHsOLyOSjpykIzVo9VBrVoj
LqrBklE8bBz0DlezAsZFXc5/ZEhEYN6MwnA5DQicJFaxq9BjHPwPwJzheethKzuKFkCW2F4f8a4s
pBDoMqyYiw8LIXo840oolkCOwXZ5T91NS7V3ojNv+eWcnL99cz8rinSLUsYI5a+v21qxOFHzohUZ
qLRWWdD62CPUYvW8vT7GA+kFUYu6WHXj4Udgx8/oiH9sFwHLBajoLnG4EenBoZpw+1p9p+j4GAlx
0PKXTcYdA+/sFo/tcIV+hOTN4rz9AK6JCH3/tREuECaJsX+z53EsHoUPxl2AzTeKNBfFyMBEzjkK
5Umm8WSllYAn/RY7T/kWyTqp+9UgTE7ewpLxjEQGoR05AMvQr2uKHovgv/GodqWuwMVM68se37rQ
PHUymh7BWGMjZWBv6tYvqDNQh4/KEfVSFRpRKx2kduPWamu3NwgNNGNmaBB3mXdx0nNKWdaftebN
y2RsxSV+bZnsCvVUn5AsvhUzT118Xn3DqjsULF7tF/HB68rdR87krry/6QTr6BoHoMe5D07SQZff
gomSmkli9d3GwvzKxOjpVSJ97NmbdfMECrMrCq2D7Bb6dpbUGE/oCy4PxGmax31Cz9VQjgXRdIax
LQC9lVaWwhjftjAjNsNfGsGbL/cRptHdkgIG7FBRuMTgTZaVaUSng4fKQe9+ynen6aBK+JaZ4MMp
123upvqIYA8raFECDgbpQmF7OajI3gHs34AJZVuDf8oKTa4/Z5fqLHqIkoQ8jjvmiG0loNx11eqX
4+mBsr4tF0gF7EvJTxY2xICADLmj6ZNnu4SOh3BOuPnwcaMh5zy3J/4C2g3kUPNAbVYf79qoHbbc
vMgKYSTrKOlpiiqCo+9lqp6jQG7ZtKb1C+JnKAgEhjO+ZJzujSVYf/ncTJ1Cyjf2tt17zxzzS0lW
LdDU+ZJ8elkNn9bwx7MkecZr843F9Marnyy033Nk7IbLqqUk6Clpvjcut3ztpSCk569fpAjOCzrj
NG/hXBKMmhsI2QfcvNrMzUSwn9lYNgCFVHkn3gNeP3oAIi6R69RzA/fY4FEzR+SLBlK7rh0WVoZ6
gETudth9UdWfXmhv89l3rDcplbWvj//hhCMFfrgz+Ghofqu2yWsyDyoEDasrDsVvW3yCACK/QAKo
MWJunDhrgs29ZYeoF8XZQB1IvJlWLo6qo+4MpszR/KHqOpcqO9YmHAoZBKITyrZDcZ+3EBmACid3
vO6+W1kv9a3MSnDRPAhI3bnqYQimKB8FaHKxBx/MH+P7akOjoV7xei9aWUnuvumTJkYENwPe4bpZ
18mx2WQ7MaqCacqOhT5YCQ9VgNoUgZIjn8GZM1VM2b5UgPpYF8W6YGv+hQCnxwPgv/hPscp/gFAt
0au/jnHqkroAcTVBsOD4GKwl3fj+AXoQmB4HgZNy2lMM7VWrjuV8R1bhDXtM57xq4jCcm52fQZQ5
S02otQu+v5iUexhTNze16ZEVaapbUxqWVsqTvcJNZU4L6KwnIUUKNb9MPv/bRZMGFwbQQcp+LZ7b
c9gPkjg7ZouARCNiJczD4LL97axFCYeNdBjwh00sIpfbDED4tdzlx0fsE6C8mFdK0sO6XNiWz1EX
F6XYTZXayQr8JM9t1VwulnJLglrHIkIic5dCAyP+4P0DYtmySp5kl93AMTtTJZaihG/XNPO5t7ch
y213pGfn7It33xnosNy4Xtzldu+BPEwb7WoRsJWkBVVKKh8d+dmnrXWlxqyPmOD8AgptG+6qSoJP
vOvzJLOfFv7adXz99Dvn1v5k42HDqmJTysy3RwAXmZBdAbNnulPXSXuwamoZwQrxLCRk0F8vfn7e
4R8CPsH4n3vvrC9PZ14cW4AQwg8cP/RozqleQK3YAndTuCX8Ji1GKjZuUuFFNOWkMmtLsdOgc71Y
5JQ7tmC9syNtUCQDDZv8S7/hBT8cLbxX5XVj9o1r4A3xkZSLS6qfA8lgAteD1O/24jBoo5qPxXY8
mFvh4wYOPK7iGH6jmz1DmIHfg+teTJGmEwS2PW03Cwllaqod6DOGEmsDViDR+3RETTkcelho1ht6
LU6L+FVLz8HsZNOqEkmnoOw7mm9dPCYxFBfQMoBBXacjqJU397BzVPrwYMP9qGZYjgNuI+zDq2cU
wk1TnCc+RBj1YZL/+QB/lQJYN5NeJ4pPs9nmgsI9w6Dmjd5WhJ8fzej06HKSxPj1puPC/M4uqR5F
v8wuLT9b3nUuSG/p1VV8rF1yNc8QK/mewFQayMsZaJaCmY8LB2Ja9Yu3mUE8GCZrYEBAVMutm2My
w62VCHOqC61g7H/cd/P5J4E9SrSuujYfvvswUmvcb/gDENj9rjl4B8ll4HYMRdGeHSEwyLa4nAgA
sI0waW2m/CxtvduFfkW4zn9zSCnr/4wQjAyHi2KFXtTjGfIGqM7UBxTfMiB3SDszwCAi3hJR3dU/
maGfo2HR0wO6RcqSUhRqieEDqR1peScficQjj4h1pgNJcAgU0e92lnbgcN5PnGJWMv6+M6JhIUVJ
szZyxmYHv0dxv3NSEgt2zLPu59Qev+rodR+15/qjplTtMbMHZPT6iqW4dQ7THNoAPn2mT7yFOE4G
cnM/YThwyPlhxYact0NmdZA0jXN6geXrL2JPSbdIngDR2t18UipKLlcFZEicwAEmS0zo0fnaoGwR
iZ6sXQ0zpDEf/hPLaxvKRGybxp5uErufN/oQRAehxvQKyjLvAg7tXyGlfdpurocsIyaOXuRWvXi3
bsyZ44oqsgHOABaqwNUfBYVfriHNib4tWR/P/AXghV/aj1EavaWwh5GnOY2O5cZe1gd4DI68T6co
2syut9gmmLkMyXUO+ZMqhJAafSQL8wcuQ8YmkNK4XC2gCLkIErc2bb0uhGYmgBvdu2vI+UEBxOMr
9Dr5WQvXwSGXZgr5ZZeg5EGYhZZnestw/bB9IyJWIFrMS+A2R53uUgn2THzTpfdlEKkC9pdWwrel
CG8EE1X+d/o0m3Hnc+r2p2KqHSFzQSSwuUAxuctuo/8kXuO/FdDbEZewjgYfLts1sRnbtziiEejM
f4YtBHJwsJ2rt4QD5RDfafH84Xg2ipgyeiEnNJsoaKsEX/3Evzfaa0R2RyD9RgD6XFPPghUwkV7S
R12OBb+sIU6OF4/iE++hE6M7Yya2MLYIbXyb4KGFgr+f1diFbNZ+eWVeeNlZp9mX/F96R2xUcXqW
vuXd7xUAoJb9x4mGs5AZRgoOGGnPdCJ2bjmhunf98gTYAWb0C8QOkkx/2699ut/Oxftogli2OUXv
92Jio3DehbjKSdMasG+7fiZkBrJ2sO/XzMQHFFG1ImQrGPk+wG4Hz6wYp/ruZDWI3IEt6mbGlLhS
l4sTxHMEiuiBnSGePFMeN0238g8keMKLl7TSyExzM0qfhaKWVL1M2pUG1qOpRYhrkHQej10NsMAC
vPbUe/uSLgi6ZCvFHXcU7G6doI9sAJOOlU/zHME06M0qJm5ambZOKaSL7Q9+ixpwZzrt0MhRpiW+
VZIFJ0fpOR8IOcbM4ihh+c0lycynuBM1qXOXQCyuSxSz8MyIuGLumPj2jwAYo2r7NYd7s6ozOoJR
Fi7oI/JT/3I9Z9EOdjNJV7ho/c+Z+iGgtVb6o4zJdhNl1ZKAlGC3XR/9GxGEIkz/x7EDtPqgWa+M
UQCDvU/S6dbdjnDPCiMuU8lksD9cUTZmjWEUy1CEBmE9PT1TdmS9DqQPuLn1qo65+pLYo6ewv0PJ
t9O3dW/qwe1rZyF1/Bzq6crstRkFfJ+HohrtWQ5tzZhqGH7FUlyZ2cQ/sPGtfWxjojbX+NmU8gRZ
mdOJ0T9EcdwmNF396W7616wesKqSTa4qrrVGRPL2MnZh8YhZ/wHri++PNOc/MOhPP2JBGWgg9iUK
ifrGBE4ucOc2SE3CYuy1CrEABXpcM9jQJGLwMJvo5vceZOo8PysBz1cRoaMkrMMXotT6KM4wnONF
AGbU82Z+HATbimgkrzu+ih7oaVdDGS9uPPV1W/xFHSRYiC3GNu6awbn3CHGhWHSDUlZ17yGkF+p5
Wbi6frtOc91jXPrTScncdkBrF8UUEB7Zm1b1aRpnH66VvC5TRFGNifDV9Zk2/z2l/tjCEao9w+0F
WgM7R6Y0TV4vrtlZmkr4PaWf6etKA/VReJJ0GqIOCN9abVtUD2oWi/DKTnurl2zU5YTxfRWYwtZz
40LJLLpOsyWuQPctDDnLjtCi8UQsvGTM2abZ1sZ9C6HKgPo1HpmKSbHojKERoPJZcwQrYMgW7hKU
UQLD9hbQGoQfl4/uSI7YgxaOr/wF1ES1EMA0d7RlUpJxrw6h7mn+gvQ6aJnL3PCUIHaBjjnLDtXY
0gPVrz+ohPX1QA9CbHok2wUEiXPWscW1qSALL/lC86gr7zXJ41iUi2fgixJcAeyR9cUxuK0rlD6J
BcWSLXkfatdR3CYTXIqCt92JxCXTAhX42LZkEuk9BqRSZO1AD2dR3Gvn3CSDWf7qMfhH4glka4Ao
RaHacBnlY9hnPKYK/hnBedUuuDn7dB5JV3K8Js3eKWXVnKdSXaqHBdx3SJLCXgH/82Jcpu7CkwwV
Qa2V4tOZYEkws2GshTE+Wu51G7eHkr0MulyEEWNgzqNt6LseVP6I+HNFxC6JoGEBnpUdIuS+Ou46
1+9gtMy14lKNTC/Tf7UA+YONHhJxcIuiukBwNt645A6tV06zp0xc5r/QZYmkzgLdmbDKj55G5+fX
uMSmlzsn2CEGCLzdJ14DPYhpn6uQwkuTRa1Ew5sk4AQVh3hn6umuBR8k4e24YOJBnzghVgKzjIYx
IVCTvybCLWqjNrEDzxx0RXHtzGwv8+PMPoZgeXyRUPsZ0VbuRd0WzUNnPSA035tjk7z+L/fDvwwf
Nbdk4v/MnzuNCjUiIf+bPl9nbjLb9NS9SBwNC8JuyHwaP3wY4352o9vxhGeXnJgfFDWgneuiZc3X
/pFPQ3uC/cJMO2/MizjCP96XG3LtRCvu7Wblnv1yRSpPNxFaV02zDoTDt6S1y+jvL4hBtodTj3f8
WHsqTWcAHp3yLlWrbdwCNVrtyX9BAcNUGjbyZfHahOtlQ1ICYZrck+rDl/aI1Ur8Bfe/1SmBhacg
Z0Hy4I+PiJ9wsjEiK9Yz4ooOCR6AlR/Xr7QvpNcCh8RQ73v6ZVpWoekKFPS/Ccc8rbbM7LB407HZ
beADONrMZPeeiHHGgUX92CIh2zb2NXTG6wPIUL8/H6SmDg+H8Q9rhLAaNLYKMd4RgkCLWRO4oAK0
jbr8MdKmOK5K9TWgj6ohfQ+2oplJyRCDShqEzp6V5OlHVJhaeRG6g6IFRlLXF/dV4PVGBH8ypO+9
QRAexNjmy9+8cp0VAIoDdlQGerQ/8dePTJyJI5x+co91tRgR6GD4vNGltolDEfZK1dZ9oP0sOV9O
Ch8jEFTrTjVVSC/JPcFYdoZoSloo1BXXTKaSoDAVmByTu98mefMMVy0fCdXorgM32zVIZXH/SOKD
Wu8quTEo8ulSHbdA/LQ7sC7jmB6aHib1DCJORa58vSOdiwJJ8/ahgnwT7WUcArpq32qsW7dQ05VH
0vhWjKBlHjcgh13HBbSayu3bmdfRURMA5xqzXX23bexJCBdv/apkIQm3+NV6V8LL3HQwzMtiG767
+c7Qvjngn3secYh55coepxTuMSBC5UmT7pAYxxkbWUEZCWt7PEEovVenp0TEcXM0GQCGc1Kn+9bn
L8+CRTXh3xtTmFFWZ671JrsDXGyzrbr8RGLAzAUr5CRGfAFRnVFwCj3ds3TWu9OOMx1l15HGmeBQ
0OLRo5GRkHM50dwvyNAyg0KhFIAkaTmOQaHliv+RwxCoVrc/0/kZcQFkOfzO2nqMxzwkoSNxAZRz
jb/EGHZ/q+Mvh6KGJHFsH7nZJOfHaSxyXSyaWLFhE5lNzhBBQ85duM5modZOvl27lgatDYzhnnQU
BYhVZ5p5JMvcg93ININcpbsy7F0HWE/kG41EaxdCrEDr83TfvYcwqBfGWo/gJNBBEIhVlYhBTQrD
S/Lqldxg84AQMdus9eYYAffRkQe+qBYljtuWEk7pKOg6OlBlNdyhKipeixgtvT3fxnpMuTR+Lwbx
zFs04fV5EKLnCTKSnqjqQp2UHPhF7AMfkvwgA9xeJ5oOoNxF6b2yC/BtXgJi8FcGXGvq7NdJrXgB
cW49/WV4/R/6QO8a9yS4aKJoLUdtzXWUJc50wGigEdi4gb0vuHJXdeVQRcnr7cxvdGcqiyrPH8NO
CofSW7+PIYCFg8FEqNWdG8sdJNVbM/aJ7JghrEHVZoReONqS6n7ZWhauJbDI/JsHshGT9sJcuhqU
p4t+K9XyEiOgOy88BECArEK/CHtd8Q7J18T0t9xmd//uUtPxoblCULK2lw3gxT/429Z43JIJaEkj
sqJG3xLO9OXVsQ6/QdWISnnrTRS7K67pnUXz+U3rHErHYQoM05Gld73siwx2+BmKU8Esu3hb5pZK
ruNy3805SHA3d6tWKfVeuuAaibTOCUFj9PIF/9kMtO9fbZgFKUXehbJF/xWveKKu4ObyjdKQbRh4
kJBW7kKD3m2k88W7Jle7Z8Kok6PN0MS7DcsfagaFchS3HhWtWP88WbkX9ReNB05fvKIbUObWjYTS
e/bXeViwkK/qOiNJf1ozW0lykLipWJfSIazjHCLsI6slyQOgdZr6VXD0AFPCHXPISaHSd7S2Oh3+
Bd1j6Mnl8bzxOaCqKMa78k5+m9m72ODvwnFxkSy/B5mXgqTETk042H5txKiiYTVKiJeSeOFrkO26
/NYAwwhR4mr2mTLPpqNOervsHMrm7LzPHh2N8whks5g73gum+KYCAMIJseNkoSRMh+C92KY8YrVJ
PFIv1/qTAm6AzA4dycPw0ksAy4u8eDNGF+04GldlIghxmtSHi5li6a4raNl/eGm3Rwy7v2bqoefR
fGhPjVKajoUfoPv7iHKfyKK3DXU1nCW9JZE3/motxiOu6/OTTOSpJkntonqADXwb4QtC3KuT0sKZ
jYp7XFNTUAot0QiGVE4YlBsDOPiqV9vdZ5uWmGtVMjMPQ5XPsj1DHQTUR9JXzlzPC8urQtYdvCcN
i/SVgoqBTyyoGiWhoEuqWQrWTp4C6dlW8zfsYpT+DEbMQ/TRUOEABjW+Zx9W/2KdmWuzZJud+XWf
KQUWYz1AAeT6kG7Sc3C6mtXp1GKsuqyftGAwk0gnckgueBeWRw8iIaEZHJ3RqfjgMS7QXWJA/Qlz
cspYQtlYSY7dmDyQS0pTzak2tWGDDPNnkHtS6Bp9SBZtgtGwqZta4tR4evf4PxIfi7sbCFzSzKor
w1gwqacflXh61BW2uVmJMXhMyjJMBY8GZgG1namxqHDcDMw71FcRpEaAzF65BZmZZzXtbXWFXGOS
StWsGTlB4XyLi5IWfYCBLHJ+rc9ZtvwCEyCA0ssBmR9Kh/IAnDkaBnPtn0EI+7oeNc2PwIUeYajx
zuSxN2OECnFyaF60bFgdtawThef5uo39WjueZtG2manFCBS7ETBvwiXudqjz4Rg2cP56HUFfPX4G
zRf2h7VrGsfJT6D7jtagid5A+RsNn/czjeJWC4exDZE6/MsZbQSmXdVsa7TfIDBfj1QPJByq67Fr
7RI93X6Xqbmq2sLjab8yoKCgxKJOUTDWZP8/86tD5kMEZDeqNidsNtrZyyCfd8IlXVbEA8m9dOR7
cuAXyLSCdUkEQvJGvLiXvDr359ZuB5TVJuioQw2n3ts60OB9P/SCkyTgDGrKxbfomE44gp9Ily/h
GD8yF5aAhn/GaGfLxJtxuD3aYlYjWgi8gFYg68cQard04ZcSYiI5o17RM6+AKo1FeAvtcXNH8ZRC
f2IKitqHbM+rbozwd4ta2bVaOgJaFoW5sQpVqO2x9qlcOPqW9JsRHgnCTOMV02SDHHZ+BwKnaP/N
omagmlFNnW8OmGVW9/zTy2CkaU1ngVcVROKfypjv5BgbuSMAbojUyqRxdBiJkGJfRLkNyOXVszv+
PddA9R387Cd9zk0XRv/aaj1u77AuusVbrFLo+dU90rQwXeVG3FGPaoI5MFliFj1s3NFTULXaQwtb
ZQ3yndOMFjAbDTMXxWMjgeoiWRN3JDBfRFe4TNWye/n6ShbNW/3ibsVXmlHeyYcHTZyvL2Nj9gbg
Sppv6G4mno2SUveNQ7AtB7A227g1HI2mEvsf9sUyVgMdf2ImLmT/AA/lolFPTbu+Ai8Tlj4B8dlY
3+1JjHwj9maN8MUDpekPS9kXajPflcdA+DTzgLCs2DMnFaW3hudxI0mBJFDN/baB6PzUs1exUL57
Um3bSlGyE0CKh9RYEyuAfxdp0jJh45r5B4MaXjtQkpJNiOik6vuBzb53ouERrfm3fIwvVtpF7NLW
xp3g3h6rzQAqf1BFecof4IYNQn2ooSzJ/HkyK7K5BGDjyrGd38NtvNsyDbnqWQWW86oNDheZ4kC+
OJpJg6a7FdaMRdo9fD/nbFjcZ2JY0REMweJnqGnE1kKwA+FOLwieEwRbS6DIn0TC5OCgZxtED7M9
OD4TwpvUOXFDV+nsAQYSUOwcerqEgfnvBvjYBs0dxvsmzQDexOHEbbvkUBwN0kpy6GH1bC+VJdiU
wmTXaim4aSX+hvW+dCBlfIstKVm2Wlo7mltJERxhmfWrsDrOK5M1y/pDD4SmD05LlftxW+3QSTCP
HMFmJFZCjD5f+X72Wz4BnaTqKiFzv5OyJa1ZUw+LcXRZWQAHc3+oWwN6HVqID+DvxG7dEQPUtbYu
G4+Di3KEAh8kovvfRQcjL4WK53eT6qq1DV1IhdsT5MXxxIVxqhoSGpt7nj4XEMBLvlCfkPPQzZzo
jL3UwFOe577rnUjL+FPJhawWOOxQT/NjfSwqoGQLybg6eV+G4jdfKKHlx7z7+XSf/oXYwN+XfCQe
sb9m/4D4yN5erRcWQNXObUoXREYgibhxtT5dqd1XjfbAR4+kEeZTGkhKlgh3yGHhkrD6Q6xB0euT
8waxX7gXPSPolovsEZ4I475jXp7t+1gkxqqb/rf+bxDYfgjIdWtqF8AuSL0vvYFCayw+8P9lpoQn
z0BWvTn/3vbj0n3R8Hrk+Zgj22t8HnPldlwjW/1acJEm/Zy6kUjpCiRiFac9R2MVkTL2YGww6GjM
9TdaFyMEWHFReuWKB+VFvvcBzW34cM9Wo+FFCrxAYQsjg2uHF7oXp7+Fim2xXGBiwHE2jklx5WG1
ktH37JnO6sQ8NKpozWw3AJzOiKge9AAj3HAS8uQvX61sGaqBGScUtn3wBVsuV9oi3+5GnJ+JheIV
n+StsTsl4yH1apAbL6STnTgSy7rLSAeomscXkXkj61FWQQJ4NsommhCff/N5N5+xzQb3gsNq+XDL
FNc/jj2DFtA9CK6iLr4mAmmTBDXTzX6Y+vOPrSrBVdCttUDptbbmSWAj04GLYwdzRSH5iKfmC7f0
F4oRalaPf+RGWc6bmVbKuXN9GNywPAjOTrVBeUN+GQm+li5LOtfYZH2DsJzw04W9/5tEUiX2Xi8z
JHThRk5q29uIqP7le00UF4/9bnQ/PHFJZxnppm5KENM68GlNzP8QLEb7vamr31AKoUKJ/tzGHB7e
mah1rJDpAOKhQk6r7sVQunslS5OT4uZDHb+Nvip0ZDttoSzzbvYUwgyyWTIzqdVRgEZUBWGIYZ0k
h9jR7/7xmFQ5y7Oix+nw9iRK4pzgpkFaOqDdyuG2ilqA+4kZEFehm0IHBViHmuMlRO7QdYHqZLVt
zYUcYy4OF1YH5siC31DGB4ycyFAO8BnlQwjmpzjA7iF9xax8MVDskynY3NYOL0hE5Sq05gSrUV/D
qBYzffNqd7TBENFS+ZEpdA70eAXXaZKXNcYUxikOmEFttK/raOxToM1aA/dWvsyE69ajVcJI802g
pC1Zd5ZDlTLa4og7eXWvZXSvlDAjPBegF/qu+kMsbpLU1dEedaCfO9EfBwvz52bGLFTWd0oS4SU1
WTAQKDPZfAGiJDI2ifK20D15P/3xCN7R7Rzzv/copLBpzz4pVDrihNqB+ss3YlD3cKHkGvePSWd8
BEsf38nk6fznCej0Jpi/9GfAA/WnvOuTmHLwQW2+tAmZEjgzGkGLuXvbuf5nOdsQFHi/xE08Dc2z
N4QeHXxHz28p380+qgtlgqBf8QhnVFqzEbOxs0aLzyDWg6TLAOKBBn+3mOeeqYwQUUQLojR27LZI
iK69zGpCFdHHe6DnjbcwnaeRj5axW4+syZwfxOGDXwqL9SRi2Cq43m6d4j9aVU/BLKZyGG7ibmGi
hvYx7xl3BN7wPDAItNccR5yBlBB8Qu9ZXOgVJYAYVBIfc1xJa0umG8hF4PPQNm2Bxkyb73ZR0ovy
9QKj80v/Dvr3vezOeXwBMXIWX7x9t/Y5uw0vyBLopMZHNHiGDOXjkGGZnhud48ea/Ouly4nPm/42
K8epx+qW7WokYtsv3Clh6mF6OTkg8+kgJ9M2DdPGYopSu/t3Hd+r14sOivCxYrrnGM0xpsAlcXES
io5dd6m/C+iVD6QcBAj0fyzkAEkvSkxiwZJ4otOnIQD1X6cOSeTAtCGBzJVK+yli2dyg3FYOz/bu
oxGBB8YBsCGae04DJ1uJdWonU8taNl2nQxG+6ic5/3pbwhtKzPSANvxB1ms3+JQfsyLF/aaJSZaY
4HU/6WnjWE6OSqr5EXRumSKIyW333ugLgUh/bfJGV6qNjSQ2fBFTr6Lp9DNvonz08PaJ0E/jZkdm
VBsiheZWrQFLZKyO0Bg7k8ZqtB7kopkUg0020kanKrQ0nT4+cLWc1FhHq9TfPneqkpZkbxiJwRxb
DkeRY4IDIDt/fwssJ9iDR84iCAwPTVZrDnoIG10f0LSz+8U5X4883Qa+5AaHai0uddiGz6YGAjfk
JAq8xiQFZLB/4X31XuuI0sqevQRx3ON0JL3iBsned2vMav6G1jldWwu2LIarGmAmT0bkmZ0OE7NU
+xDoUw3p8FmGZlnWKzvAm5t4qsh5+/F9SqJQmy2E9w+EuYTiFRpw2Dw9QNGcZeWKCDml6zqVWko5
bwSRZd/cowbGGR6NAy9FI9SRdgx7mNHYVwD8VMfyADKPa+BqsKNGK0Z3G8KGQdhDZHAt184hPEP3
kN2vASow2evX2Q8zFrbZE+xFUpwPvbCx7yJrM23hWKAHUCEj4WUZVUs+eW7O+N6QYXHCc0aYkzLx
bWVLy2popcXn1fC6Pmz8YTx+BlrLFlmeIb0HoqZSDTqJZTeZdusJd40I52bnAEVXiVffkwQlfKOY
NXnuHEbywHK4LJmeTjBp37ZDKY4JmDlP187+ZdCDeOgS40xPt+WkwrzS0Y8SLptsJ8HtzjM7EBsw
2wbwZFP/TdQDZn1rlb1tGTkXmpyamemB2pDc3jl6M57g3ah16Pb1DVqya4m0nibUZc5rPMv7E1F4
3GoaRBE0xT4SrvkMdHgj/mHprEAa40vwDdOzpKt7bfYFI34xNi002C8XEStlL76mVBzY+ooXMxcv
1FF5dSEG0epojRFwp4OPGo0veeHXwGEWpABU1xN97wRGJJL03/CyLxqmVhz5qo9x/VE3Ak9R0Z1Y
p8UDXlIVV6lYJbIXv97XlVOytym4lr3ereDnZGdHwJMojjtm8F1pqPCoxgBjk51kcRU7jh17/q5I
qG22Te8Wtla8CCx4R4Xnl1+gcL8v6n93wXhi4E+R0sK+jigedlPOh+zXLbaOQwb5OgAqXXdRtgye
LiSkHd3LhGPpyirBlmUKJETlQeWrmkxJy40XGX5bEuLBMavXGmokCeqVOTrOxPB1snKWhBlfV9Y1
G1jfU8+SWfl96RkfLl8A22mDN6ZkFNYhGvtn3sn9xP6j/uCB5N28UFSLFdQ7IaewVNk3p0zyj6kb
sHpAbMifIjZBkm9Fxz+TqVDh+fivPICkJdzXPkxSX94si8qrqLrhnGCSYIJ34sbQvvU4dmVUuAuM
G/lBUmWjUwG/ScVU5JGbkVMJYOqv/h2mpPJg8xOmJo4FyK+UFP4l1O9p4AnJU5MU702dmkVGbajU
hZmh2a8G36TCHgDhKCrLB4gN2U6m8IClfT2km49FiTkikPP7kOBOH40ODMQtj5PW11CtETnTAuKM
zqXWdrY9347auN39QZX+rMzmyGCgLi6zgTO1ti7P6PZh8u70foEnJfS01luAjXZhlciptj5l4Hyv
fZd0kSzc+U7V/gFgXEd3Zq0g7eDGk3JpkDjgPGriCeBnxT4vTGupg1yXQSqxSjJnvSF4J19ritSr
N93+3jCcZkX/+xJz+M32QA2H4SpbWrM4LEnzR1J7V+mXIzuJCWxiLI05o24Qxs0Hpkv72vmFYagk
GL7tqZSIhG+tSZmgpsqRvyBhwOMhcSrEfNWFSkhEcW9DiPq3mVbL2Plj0bRAuz5mU96tCYcJ7hYU
iyyimkT+YSyqpHl+p2rMuh/YGRNnxNtyUuRwu/SAWhL52e+a1dPA1wvXULu3Shu781UVgrTX27fv
k2gboUoLT6VUnDvZGkAjq148ackhka8GwYCRO12HjWBLMoK28WqG+UFst5x/nbQNAxEGM8AjmR6o
GbgeirYzzxRZmhrD7F8Dypkrs4k7KSD4FHEvwCIhOUJ+zCVEFssW7UDbVfOIqbrm8qizWHmRs4Xm
Dfbi5/+wOKRCcKSLP41HO7bEEAwY2a0NFBYhJg/YqInzNZtE2OpoMtqZJrVcKKnQz2FUp+aMDimF
hVRNL3Tmpe5EC6B4NjSJuJtSAoRJZbWU4hxeoLNoDrS0CrzIZQMCWikUlWFcuJP5THe13vgLVf7d
Y5+qzqpI7ILkHRB7ibVdWKxaMegs2VfaBF0eubmSX4HsSnsMhdlpIRYQqzcYyWYnke5w7Yu9ykw9
hirelUQ5tCuYmaWUypIDH3oEETa7X9bS+eDzPIWAIvHipFfflg5FbCb3wQkoE3AxifnZI8BhJ/jI
pwfB7lWiJVU2fTbDeqEqoQKgWqZA/CZvfz57IRzG7nXSATJL+8LWxENlKX2m8r764CJIK/AKCEja
CciD9lUHrXpzdtZuvow4OH0aBMv8qKXQ2ueGIRgXBLSXJj+aaQltRmawNDb1sCvkGoxNgc/O9PaI
BDTtmHyW0n1czsYpd+0rwVtxAqYb49Z6Aarl17dFCiuQ0rwvxcQB/aNzsAU53rAEg6Z+AcTVU/au
XwGoI72fUh0jK0rByMKibw3f4u8ypsillKSGzn1Guck30jIQAlQCO45jqUGeI8YBGV5lc6eTGUxN
kvXiMt+s9ICPtg6iU+AgGlF4oLovktjZOq4+dD5qdmDsrcvLKR6HsUO+MR+X7o1NnHs9GQkonAfv
y8Fe6k38xfOH+dKR+FV9YSQ0zrexFJN/qLHjXqkxMO7cKT7z8kgY9mi2rsgKJ2/ud1b0ERtTN2x9
bRl6XGafQ2QpQyICM+0WEJ6kndt/kVeeQ55YMRVLgGMfN6J279miDB0sIZK9gjF8QDVjV8r/p/1u
qQIGrA/ID8fGEfSyhghR5B/ZIDGOCfSu33NfO9GdIkzR2MYuvOM0O1NuHLeUWkX3cpTXBy3dTyOG
DvKT4bZB0B76Ju5bfASd789gOFVp//qcDU9+Qlz9MLNOm5Byimqco0Sjk8LSDxjssMcXQDBuDZtZ
X62zAWq0XyQ3uvImtbcQJaxSpbN6EAZubxkWSXvtUXzfVhrolEOaWhhrvKJAtP0DATbQ2Z64T/lt
9UsjawyQKzV29Yn1tXY+OPT6fFoFvjptA0JemIxBzYSppN1iBtee+XY6HrVlBbz/L9ox+8mvnzj0
snr6HcXpOVUJRTROHVXaW+s1RJipSSmu7JC3jKJN/kI5GrpK0D6LuJACgpyPyYj/WjfQUNijUi++
d2tUJWxc9ONxAVcxW3fTfGwcTjOWrXt80Nmk89E5niKRBlUdjSzm9jpni2B/76Bgp8agJmr0tD/v
wmLy0chRxl7w/CWT11Y68zx38ttc6xmeY1ipJ+ExvuNYWcoI8qiAgNf12LkSfjxuWWy55EUyap+F
HS86exEY8RcpTopFhjRwLFsSxT/hbIGAMwXredCsKaZS8gOMon+Z0DyY7FfrSmpl9AoW/Stw0GbF
WxklET4c4gfUX41EbyAxwJkehPwKn0jriKhbRjU9bXg8MHUA98MbLnxXo8rEoSvzJNNK/3BBHF0Q
/2dehDPBlo1hTBsdC8k32bR47J/4OQjzzXaVqbxECrTc5Nyi4VwX9aT9chz7lHvtsZaNs3HdaimV
zO2AQAFlHvFcFuaEwj4+iViZyxuCpAoCNF4Cx7y4jbdRcdU5rDBBKXv8GRW2iAuLqVsh0y7ySL2y
RgPypDB/k6VsKgrOor7hDtA0tq6w12ma/sZbaTMcXujUwuotqvUI/5XaJInnHG42Rac+lUICBf3N
vyOhVEc9oDu0tqqxy3oR2rk5MoB40gM166Dq5pt22yhx1jFI9iB+7OCTkgE/jiVaSCH3Vk/ijFQu
2WvEYLoCYv/A/lmImnq+ckT2xM8rs4jiJW68NLRr2LHh5ZT1QGibOXtCEtCmQAbLGUQpV8panDPB
oH9aPfAeM/1jw/rgVvr2I2krot/Y5xJQW4dLpC2Bee06WIcNi5nYsAFH3ZuLKtDta+g9sNahipFw
O/UrUgntNiA7V/dDh63K9u2uZUHVXZKy5V2XLA61+Be3FLow2YHG4zDi3CdTvOWw4T7voxRG1hq5
FoPyzZB0hxldUG6c+ErqQrL2/6KVsLv7mrOmBkhzLyOdImJN0Mw9iV5CnuTi0QioSGTPmiu3uSU8
Yspj5SNugnuzraOBl7xeke2leGnaqtw623CTSoLNwmoWEvINt8jMeL2VOg5AI1JZk59afpxk0WnI
hK2srzypkN++ygqEUTWkn1x3nUdPrcoZjLwz0u/3gkdFX3fhdou7VIiJK6w6qAUpyZjY2lqtsww9
pI4i4q7AXLiOmSrqSZ8msoeGnjmGTaLpIM24eyejkDjKPduztgE9xXX0C1hhuCHufxOidmd4jk+F
que2PK2th82e2D6gY0D4Ze9pRfJGKwsIRPl6Z7qwC4Zk94thEup9zLfKcGXy7VtEnuIKUo9/VcqI
I7gOLPaMeOB5DUAHB7vG1uk0IRNLqv9aNS3D5dk1mMscLW/wUlIdS4UIQocC28MeZq4wV4EuKxAt
HySNIK1/MYuFGkHhOMtWGAWi4kaDJjoYO+Zs+CbbqdbjpytbWKWepr7kZyr9tCq2/xLQHfhDXexy
Ix5TNOxaXrXqvQEasjDr1VYvyr4SEwqX/IThU3WRK0bqvxsD/y7M8iEZjG8nMjNJrZXb+3AK9Qt6
KGvJmNgB+igmkiIptActZcEJI71shJ5B+qg7EOCAokl+cnFVdujLoPd4WnGmWlA6ueJZA6umox3j
TagtlP6/MbPlNqGQcx0fxE1fsRf8v2+DLrRUeOEUmy3vgOQfzNG1IN4u78OhYgFvNULQMqG7Dj2s
57Ti3J6ujqW+mXoUMDgJ9mVPUkN+8QQ9r6bd9qIXAVhVpBmz9c3TdsGtiN5Inhy8GhU/PWyxXd4G
UkIyVBxXmfCE7NGzhp3FUjPMGkMURLnbUql+miss2YKcbnpgrBYSRIupx6uz1xafrnXU/oDKKcQX
jLS4YYq7V0SnlwGUfwxjFv0JrnSBdCVxIPcUKPMox6HDWMVyZgccpDLJ8YzxprvKbNGGrm1jXrm4
e7Qba4VHvsvWDsfFg6LSBHWTr8ZuLxEOD6060bhmCY4bynd1VSUzGORIHEZWbjAjv+rxzqb1dMpd
l1id75IX9DH5AaugurRsewFxapUWM4MSQYYfSXZP9sc/uPovnzOcDl4WbOYe8hJVvdK35seR88te
iziriBfktoZuPxQDTBNmKL1aA41Jn4tB+tl1hWwouDUkYGbaaJ9WPiELui7PQYiCxQkJPhZ99TOH
V9KhhGqlsVyq7HOM9HyH0Mq5d+ZUPeejkr1J1A4guFVXBh1OlxlSVmi4t9+VLK0QVLnXO+3FeiV6
jGQ6Wlc7/4nHNiHH6HOaj2lgmmzTt0+E9pScCbxceG1Zvfyi4vBUt3rdDr5X+Uz/8Cbp1RDlqwEa
4EuaPOt3oMlFeAldZgluETiTMGZE1Zku8v42b+TbFnnLTfNQ6lzEQ/X1HMDG1zXruwlCXkTpK/CM
65xBmX6sIPW+ezw66n/xLZW73VgMiby1oviUnNp/kwl3zuckexguA1z9ZfwilzB22TARqyqycfY7
XWyX77IDin5ICIPBiimoNIurbmaiKFX0EtjQEwhaJm67oO88qq/JgDm93d9jOeG73MTRKX9P1lwH
h3kXaKcWNqWiYvrmG983alfqo0UkUZMTV45Oxao+CeP58HtMIEb2r+9DYQY3Dwgq9Ct01ozYSLnk
Yj73u+t4QUD1KWA2vAB+XepoeYESeeDYyCZATU454hV1QEeQ1/TRD54eskrqWf85Ztd/ExD2/m+B
0LguLyiswivHs9uZrS58FWZXFZ18RNtRtbWjTLGQCWSxCw81O/NIbftm+4VIK1TJUdXpVbdmxjGB
NorPSWl+6R3SOrRIW6XMRXSyfZpxDtU4YmDgSNCcrNXLBafwtSlwJr/Xm/EO2XAaahnOYaUhMYlu
i6uNgjajPlGmUQB69Gu+UU12ARV+CeKvug+l9VYFSOVbaiKrTqZLTl27HkhJ8rlNj4X5mEPcOmQg
uQptYW6OHd1JwQ2Tpl9mgJJmZGz2EFZPfp8Afjyn0x5JK4Xo2Xq4kn6bf4Lqnc8ex0cwbR8BqaRQ
KEPg/kCcxOK9CfNqhTlkXMw3G16oxvj1X7GSlvDVS1Pc8sp1VDXpGyq1XO32WCVdUO76l697lfpn
AhCoph8emomagRMeDc7qslk5quejX0MO/8UsQkk0lhJsqV48PNuGF7PmxsLq8KKNYiPGsS7cQb+n
tbkBieIpb8iHZkFoYryIbkm1ErpJOc25S5Rhnnk9sL38NvugzAvMDY5jTm2bn4Y+utX6DXdhSlIH
70MEhISC2J0WaM6kPqwwSBpOzzKmcHLQT1zm4ykElP3Zir4nd49upd/S4mwj9vLtzhVZYUnNs5Lm
FuQB2kKcVowqM6nIubbheg/tUtoU7beMiTrg1TSbYUJcHi8u0oI/dNbc+QRVt7RtFYA5AVq6TGJd
/pafT9rxr6nZADLNi9KX5jHwr1b/VuzH/17k3r5dRMA86h62EDwY1WO/eP6jPUIATrgZi55j4EVY
+0ELfN2H86YDjX2Jb3qodboDCW8muH/42Baix3eS8wuUFnlLBV6uCknFJzn+ofMPllUOIjFU9bTP
kUMa3eF3HrR73x45cw06Y+DvfSXbdAC1MAEBfHooUOnuYLkRrG2Tm3A5Y/QNaZKPYCoR4T7We+AZ
QmFb1lcPzGwapvQo1kR+CXAMf/tqy5lMdZXcvT3lBXhf3hOS8FWg0SuXEa0NGasp0TSMM5uWIGMe
rSnO5fKb6SjsSO0IM1SwFl4YbIiO//vdO7LiCq9c3+GlS+0s91p6m9mrxbuxBgm0NsECnp4x/kIG
IalElP8cFgHtekScWZ8EuMXgFWOQUVNV3MSPjc4LmO60lL1tsUvJWbLTDSDP+MdnBFT3b7Knw18p
iiX3U6fZMS5hGm0Okb8rTXmbImb+oLG4J8j74sU2sXkExUibdBz33CISDCn2VDTamvzi1yceP0LQ
Jt2W8ABJVaoWwrcILJSF4YwgUwDKAbGSvCKkzn1tgGYGEEn1Ii/pp6uDLbxlwRx8qtwVNZZ80v+m
QDee6VlqMyrOzb+H2urunx0xtEPHIrFJZuEciO6geTFqALVfrFjjWfnOJmk7NYZGsaSb4X3b0c3E
CyZU4odl9CmqyEpcc7K1E5Tt83/QWnLbuI2ox2aKA9XiMibWBBStBEc77xGx8QmW0/QcuZRHiMZZ
dDMdfq4bbwcDHTb52oDdyE8UpJAC4BAsF2F1ke5T1f1vp5Q/2byMk1zP96J6KMlMLt8lJ5LTxzCk
GtIxXxXqw0UX/pHVHF8o30W8u03wmc5p/JmJkGBeTGMt3r6N5xW0P5zM7aBiCDRoo+i4sIORgfWg
bJ5ddpSwvDZex8e/8B06cSexqvoUMw/rxXLtB3ybEAn531cI+0N5wW2Gb8PJ23EXNIwhqHbBw6Kj
wruROQNXX2UyLAbNxyGXM3Me+CjZOlShIaAdNXxYCGe98km/CMOZUKEH+TXT9e9aV/8LRWYVAdZe
SMzfUDhO8DVUry96EMOTBg/q/3cNiFj8bEuQputYQo4pgADgQavZbaBRnWF85H9T7WvQJh3nqQdw
S0EdEwufx2d96wWl9uC6k1En/kYYvCWEivWy6jw/LDMut34IlQi1DRLRslXGvaj9W9veJ2drVr0X
mCe1VeYAdY6ClXAsJo/ioGI1VFi90xEtzac/6O333jb6lztSfJ/8THdz4YhbyBHGQrcuZDO+e+fV
pIbPlt0vSsNuK0kYk5PvolwaLmnGoKFPCD5SCV1l9q4tD6igMI0wvmpqUuNJYmDTVVAqZbsnW7oF
zosX+Du55O/FAXlGL0jdV3tae6eVcFBezIf6rqNMdEPkSukNLf+J7jQOBm0Xtol/pX9iT0U2Q0cf
J7Md5AAa71zmrQyyYj0jHtnL6fRgQK4LWVZlKQUEcivhMF6qq1toufn+DnXjWHpyv3v44VupS8Ve
olQmoU2CNMSjvhwiG71uqVnIptZSzMBEcpTX5tVGSRhmJgdj4ZTx0Kb8mttsGixCldyLb6iptGDg
9Ub7UznD5Ae9hfERHssLBYdhk5rwnZJ7PNNj65fUllCzaReSU+ofGKg8dd37iRV5QtZElFuHU2dj
OA8s8c61HkAz1w0/7TOX81m1IZTPocpiWO/am4XvyvL9glpDUO61En6NZG0DlCF02mhW09SCB7Xb
zxNC69/qEWZ4cJEbdHLNdYsauj/NfjRCA36EM0pWMCsTK3L9reoJNJ2FAu5ZDRaRPu/WduixAD8j
cOWRiiK3W6ka1rYK7hwb+E7rMeqcyjc/U+HBC4d9mn1xchtJF9MF6TqNRTgPmF3nD+GrRSJT3E1i
wnWJvbW+RWoDNjtlKQcxSNYb4xCUyVnS1EJ+M58Csv+A5I140c0YB3IziTCg6GP0d8gROrC93W8W
lzgd/Ts3UBDKSVt27c1WwMiwQ2AUXaXgtHmFOcbVs/KLLUXjoHPNN08DSMwMZgfd54JWNt9LOsRw
lrlYF+0KIAlfVoq3dOQ5HvnwV3PfscR8i6LcncWuKIDMMGcd6xvg+Uop7gBqBB0xEbOlBF9szlsQ
7I5iYSDemBNG5a8mTsxlCjxX4o2Y5hR93aXPvFluPGuqrzvWrbbYjPDwvsy3oTFGiIKxQ4rz5bkG
l4KGJU0Bp8uxgfhTqSdzEiI1A96oaPvUcEpeoCL5OQtf8fBi/wnyLGePT7myOceDkqh2VaYrd55s
7VA1m+2usLGLjz+TMwv/2Lria7kO9AGJRrpQ1QGhfiB/AWBmhgr7tV7TW4A9g12dn+Sc53BQuazV
P0tjW085syTr1yTHPyVnowZ/6ewcJd+kycIgUF4jVy5lX31698WHroKzD86mVeMqDNBLTSeTCCS5
AkXXGbFOjWbUJu8yS/zO9jHc6UEdmL3U4Rd1Lb2+Cq1ypbya648gSv7k5Tm2Rw1/heRtWsLfmyo+
J37wP5X43oqRSSvhPq7G4IvktrNuASVBGCZwWi9jgoDzVTedCX4B4NUuCD9pEYoNbjVJxeXAeE2C
SZRw05m2Khe0V/YBi/ZTY7/2nuD1q+yiWdHJS/74C2eDeegQpctSImeE6dsKyVVRWJQczBjSOHkM
QgQunVNJ37kZ8sddVRYVE341moKGu0+aCMwLpOC/xSgWF+UL7Ytk219HaTKyZssUiqmRmgAuJhAU
KcJRLd9WehfYqBFO+Km4xPqFfHOT3Ag7P5YH6gMAW4vPSwAOv2ozEcjhGcIOkdZWUpNvjzekcO9Z
XMgOjcDiITbsWo9yWelFrnVGUvRIwBRgNhJj2zjO4uamNExF6XuvEC0ctss8O6yWT7qSJwFXanG5
szh2UUD1htQwCbIEkp3Fr3IXs1bGt16/0ZLD9VYJRi5/ryc8L3DHO4Y20NPnrhOr/lu/peDRBt6M
G/1crkhuMxlwkTNgrQ+Cljc0m6mLIRJ9bKrIB1sdN0jAV5Wb2bpbaISJv7RdiUv7BrF8HcCfYEOj
GLsTI8Qz+xH3YcCbBBILodBkOD/n0zFTfhY7OMCinqDhdzYToJrzNNea9WdK8KfLGyaHD7YcyjFK
JDZckuywqWtnQmX5oFKqkhmxrsWQC3pJ76Y036d4tLc6INB00Pg7cBPyf+cvlsqhBwmDq67EVT30
b6PAmSUakS+0Ss2M0cdXHHXxQYVfhrPTP5Eo1INhRE9dNsJHpc276VMVndA/EnPSYX6vXbRVvyG9
Kgw8xrh+GJYsd4AXTGy1AButz5PNZiobgC1PtITjObGxq81C7U22QZr6ILNCbwx04wUMuRFloq7S
flTqJTcu2Y3TTepmDz5wdb40VIhh4rZze1EnqwRxDkCFjtZQU1ip6tyi4v+gTusQ3Trcn8jLPL9s
L2JhZ4EWZTZ22QWNfLJarwWB26OQADdkwun4NBYQuI3VP/4bmoBMm+MJ9qR9hQlktoCGEj4x5Ml8
ynZd29GXNe8cUx/itV+ulPeRLZ+FTJTwXnUglT/6NviC0v6XHh9a0oey2TbgGq0Gq8aWsxtxKx6l
mv3bNn65yc/f3MseA4Irm9j6Muzz9AclctOqGsSyuCKZ+ORarcNOi8Mq6/zmb68W8eCG/x8m8ubu
AgzeiTZuLrzbNZFWgcYdeIOrkxkjDCbUgF+iwvIaoeiRRlREI9cT7EbSk+JnmQ3ekj0Py0nTrRyu
hBbIqrn9AHSe777aPKKKZBqg/g8mG312klz8aBR80uqOLeelbbX5PaHPm+FuQaBaXoDOer7voLZp
hDeYB63lskrzBH12D9XEVLbESJuRxIpgpQWsJqkfDS3JsxihhzCGwd7OmqYIZ47G0qJ3OA26
`protect end_protected

