

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
n6SxQ4cZpYT/ILbURpz0n7m3/CtPg7Srwf+5G6B92ASMc93ahDGfXsRmbxfQ4itjqNp4bImRWGHp
TxDOCQa4ZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T+03ThTlMB5LbidY7dBVWlYp0mNjkvlbypoxh4ls7n36ZTLkklcCR9ZkGKPsYI13rJYYLwxb8HQ9
lAxKeG9QmQNzwwKufgYFwBDRimvj8pMxUUa5UvV+Um8vyzZZSQmIWtsYrZE6EEbBovwAJw8AOtaR
U6gMXGczY3zuLvGCvAw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xyeO5Evu10M+3X2Afou0ntsX5ZB/pwkUmxi6MkSVEZEp/q8vhRIBXtucD3zi9CwKskciGYDIN3V0
Echz03lkOALKA28V6TwxpTDjOCcWnPUs+SbNU9hrNos5LOcUeyT/Umkuwxvon+y1+GmmTNBs/HsN
LDp012R0drMTXSZtr1fQtCR1xHLj1REwEGmrPANPbJm5g9t7g3uQ7e+eNRUcylifmDkL5SHkZMiP
o5a6WQY9gEml+rOEV7XkaZKFEUQnZO3nxTVqbYgCz7Fr3B2jvSfBBfXQPG0AKW9Iz7aUGng8TS33
LFSc4gt02mCKBH1NOkwuxP/U3rpVs0fnK6xENA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UaJ6dwyNV7zPNxnKVFOwTBNM7GBgDixNLEFTEeGL4zxIus/wUjUkJRcBksOgUQrjesNLi9rSamfz
a+6oBrRU3NMz/a6LqvgLX0FtqLiIT69wj/tO+121sBluFxMRAbLYxwtNx0oswICZG6ot3kY7wUo8
MIP1BRyvBE7h7gUe8AY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iLkN9pn78C1qipOzfdJflxHJTY8JBXpf4rPYSCaQgqf5yt0IOulURCvwg0EGtXIXYL5OVuC8GGss
Cxal0AVlk6DQJUg5tnhgoani3XqnRusVYV7ivY3j4fNdUj8iyFUm29wArxnau/1wGXLQIbXlD+l5
Ze35HAoJRWjnvYyl2fMDrjYG0QtBEQHUh7moVIQ+kI8DwofjU8zFsu1KHGJsBje+80Fr1j2xEByY
nscMu+13hzF1cQaS+Ce+aroaWDuHJWx1kJ8/T+29qUQ8IgrJDtRVEWayMxcA9x6qrZ8JHoIeOcCa
xCl16mCCnpbqxuPBt6lvzV/n1cAzp3w9LmCffw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 87504)
`protect data_block
GJlZFfXVJOtNbKZB6P6L7k+dZ8NOc5b1pvZvJCWVU4K2amd5DIEmy7hUn0vl5VlxnFNVJ1OkfkO2
jTSwPTkgOdy3CBEZq1n0r4zWB4cn+Jba0YktWJvU3weAxxM+mUipiMWKmqWawTZsrlW5c2k7/icl
LOj4IYNLG7He98+mFYTj6N5YegNWamSZcs1HtuatE4F13SCilMfVv1vDCCO09uHC7YwPtuVIKKU3
embFbHig2Dz4LDglG9yj0aJvH3RBlGK3ib80pPwegtqnpf6FybmZe82Mc2uIhMOEGL+MKbRCuSZy
kZ3B50rW28enDuby67/cRAGPicLud0t3GlXam61t3FK4eg9I76/1z3PPM51fq/vahBZeoULVQJRp
U7p3ng0VCDjmi08yTUA8nai3EgONJkipBHHyO76ajBg1v99KsKUHmYCzEoH8Y2bBU7/TWBXHdB+l
GMVPHte7oVBTXjo42w68TUKYwwOCYmVWKt+AMC7tVTYRk20j/6ido/SZVnpRWnIKz8eD6ZZKUWUk
iTvJixN2Oqkzz07p9+1e/ypRyWPM8RSJFC47532u/9YoK4p3t6rs6/bW85AUv5AT9tle8vkt9ZCI
6KDZpTL1EaTHdgF0Sl7IGNFR7pzIXG8txNUbiZXnv9u1tJvOhVqmpIMX7ygsdJsiM8CAa8dE1fxB
/f9vR/tAbqYFg3r9qitqC9UdxcYzVfeFltxtNV0p7HdgLiUlyDsJSq5lXzo89a7RdKyNf1AM0Oz+
buOl5x7JLUYALO+RntwDrxSncAIoyONAaNI+nBxVnqT7h137kzRAoK2Z80yaJAPIrBOqcU8xtl9A
JjD+QKwHmXHeewqAxU07wbywRcseUl3A4dYU7C+TwVJw+P+n9YX68bxkUhV7htrZbNssc7bptJBG
S8CSj9rRV9pNYKVeUudKJZGiQlyYibWEJwIsXgl42qmkATbYgoCnrbkum+KOgdlOJTj6rU8KeDks
Ej4DT8iZ+LjeeMYbkSu5Ch18cNILru1fKS1yh0Bi7zJJXpnD9aaWATLuYAAkS7uw6D0VTPtIBIXC
JvC2pEIVscgjiZxfjTZORswRRCxv6GIDKy9SqR1aeMI+44yTO4iRjzDtSjJPKo3Gl+hyfFbNxJ+L
MdVtCJnbICNx9libmk6f+EMpy2qDsxv5ZgOHR6TI6qYFzFSF3egE4frcFufkNOBStWoPwoc2YLzD
nQFTVUBhucVgOkefwZ5xfRtYuLK+t6ABnF7ZV0N6STLK9+/xYF+wVnm6vKRtdR6xi+Qsrc3mqSbt
BUsGmPgOHDAcrsMVfWyGCQG3dfgUw52jwU9sDscikOmp5WnSXcGU6xaVLzSz0LJiypDuB9i+hf4T
nOrqNzlVJjFHkL0Gs7yTNleoVnjBDy3UB98CVg+PSh01xVFNQH2gb+j9pANeIHh/lD05ABU09TIj
4T2PFGDauQXLH22qEXYTdip1WmqvQURBSu3GVLioY2uejUZUmWuJBx5KNo2zA0NMci07GwvlzW2y
mSNoDRc+uhKhLlQAePnY2qLKr2NKezAoRX84upzlLw9P/TsgKlxUYqzhCUsib69R/CZ9KqBr2xEj
zuJ7IEUp05fflEPxvfNurMl0wzPzk6DpJk6z3TYWDK2Ueie14/uv3JFwTgJAn4V0/bKXonDvjBoU
lZHgYusT6qp1eX3eaDoKx9xLpMxdY4ro2Bwt/xTa/gmzqQwa1GEgnqWFP4rpceFFivs9qzPLk/uJ
pHnTPKQd1IPM27JE4aQn3zAgeninTNHVdC1fgibw9leySqXVr/UGJODT/F3QrKHlJZnF7cF0nbpH
GJQSzPNsAuaMIXUOBgE5ZiHpEWW8zSrb6SCkwbfsyXgY/e6+wVM874nfXVpEeQylNr3jnO9uEYB1
P05ibWlFmxSjjoXRSZBHWhYENb3U7uno758jnmLwDNeQTjucxdBopN/ejHyIifU8kXoYQ3wTky4d
bw/TwEhgkvt5WYMWq3WXRv3HZp+C4HDamAUAcnGG5SoOyv7LRm13CH6lOomEQ5srd5ratG5W+hTd
dkWtRM4gbQ+smH4XsjV5t8VH+jqcBAKY478y0hvNhlFdnRjeRY/FVe8IxWtnFXWs53oRJ+iRz07i
cRtqQ1Ac4YDJHWqUIbcofC0LOpipd1AI41NFRPIAh8H7pUmEQH/0kEK5JdYpd6yPUI7SFL0FDgkW
8ZdOTiMroghOmunmNCInO4B80+vUyEppaXJA9ilvvPnvhM+pv2kOpJKdYzS0MulE8nh+o/RPn64t
tefhXvFUsqtsUPz5J6VLKg+hDvy51y1NCUt+l7gWVchyRvEMaJ9hsxb3Khhiz+hoGdXJ1K+Di44D
1wAVyOLA0A9sdimlRIO3c5LpT0yX7GVBuuaDIgv4cXYpACUdEc6G4Vj3kKBxnh+c750xq0WE/WuG
QEecpxxMSVKl6JsXStmDx9DAvhPBa92E8WiCHUODG28crErlsh1hwpv5s7e/mOMV1F86p011cODk
THseyZA4PSu1PVhzX/Zgwbyh4iRi5PIyxpv+jDZS1KS8bi7Lv1hEzCigH5tCon4hoDWrc7SdNbhD
zA3p2m1J0zml42n13J6yKwl+uOfRDFL8cm3jxVnuOIgcmlxSMs8otYYZQdhTW+KSMiLwWvKM/Eby
G9PbFZZRwtFBSSVvTbpy0GpsPgEWUHEn3nFKz81WgHTGqEN6s1sBs+p6K86gHCNvENM4teYLp+IP
EPgqYel4ktAn+rmZhVWw3/9vtrr6DuhWA9feO8F9t3GqyLZ4E0fZHEfs5LV06Yq9pwWp+LSibRAI
tt/c1/e581NfgY9v6EgYzLxUVTc7uDNGyizr6KL6hDLD8DSGv37xUQk28WsVa5mP6kJnPZ5yDJuP
w0sQ8bk0J3Y+gGVHF4Hez2tJ1u5Ir+UrRriH7BKx31Pu5bX953SLjK+WVwcE85tdNDJFbmi4GRUg
B2MgAj2kSXvFapOOsNNTtrNVkLNp1YdBg7GlvxkSTd+FkNEe4Wh2VRmDUSM1LjZUJNyXl2tvAs7v
nCBA9W2HNwrrWFebqAR5mlZYpWIWraKg1R7ep7acrdszmvSAONFOUM8TzEiOIrKvjMAdiYJ9gnyf
Rt1BTGJ2Y3Z5rFb3yww/30phn5TQUNvK//tAHg5zgtqt8Uc8pZA2r73RCBq6zBUHWQv792B7jJhG
8asIHUAngmVpqf0lfPTabtEpSqqvHxCdkucLuVIiDrFg89aOJ8k9Uk47eEMWbpN9+XdNwFXf0b9Z
LzCNetVjDG80DdT3h9Bt20j6MeX+CJCfit1sPCFonP4jmXRSA78LXVE6Fo9qwSuOMXWTQPjI5IgA
JU7KSKoVSxyQE/YQIp1z80djdoiIE8JIxCY6ETL6ajayguEk2Mak0yVZsHqXd/zWPq+++kS86Hmi
SV//Z4mWx0nF5BsagB2gIHkYSMY1c8NqjaM+Lw3Zq4wPqrMkvXXlZ97hVoEqNqWFA7jcESMOSEvP
4DDTnKQbrZ4fKc50GZaX9hQCrS+9Lukeim36jJQHX72+gXImvLTW75ymvJuUiXwReU74QLc6+STI
sXzp20WbQeDxG7jO2TTv4bu/1wwdi5VPvvupw89FsWdCLs+Rkgy7cMGu9EguQLLUA1F3/3KYraqM
FRRn9VABsa+wFfys9SBQK062lEktwgZITF5yXtj2iMtxnNoQtTBDXVUV9iv1X8Vd+zdV2TENDmF5
So8egO6U1xARM/dJyZtIyCmpzL/CM398Jz9BYdHHVb6/Np/lTcZn3rKfYRlB2RmWmg6gfCyqF9WW
EWctCrw/8r9mdpurdMKjDImeLPSTlHwtLWvvZRWEgCnGzOwZOsTI4N5VBUoMEwmMHVnhBPB5fKma
nB37zI/NB12bk9P5RdRi97QUq971GxelgnohQAp1SWfwHylZ8YHVLxud8K7vXZtY6vozYPeQKjA7
8agObQWm93FUkcAX3woasjyEd8TUNPT9kHBmI9khVOLJtbOns7arvTVWjRABa8PkDoBcqR+7NcsZ
HdBsgCxLAv85YVXEdHiYtFDlBriQm8l6YpqiGjhs/S/bdi22Zy+xImVZMKYpleRU5vpR9Bu8xQlS
5Ye+im3SGf15ppu48G4g47gcO3MLOoUW3Wv/CntSCtnZcKRSwdfaq16wE1Uei/DuIOcO6G8gtEoh
UWZ6q35KlFWdLw/O+ucyFk9qdnOvXJkqLG11MyyKrEt+BsAo+8m4GD/9t5R+d0RMQjwYMtsaUsTA
JZMeegrgYysgP/Kb5LHKUfKi3v1Akt554l7c0e101WHi3pczbPRyArFI0wXl4MyowJ0FmWFtih9b
NK4Mf1OP6UNgA3CTg3FHreLREgcCqe86Jqvl4ERmui1vQtN2UHzHG3WP+7w1Ec04zj7By9cW02Bq
DBzZMhnlObqH/TiSSvRUSBMNXoisorIEfNBnADiDCUxop0nJa5xDnU6CUWdygJsg5kfzXc8ng6WG
19T2dLf7dGfBkWEAisCUw1S/J8YlYZGdRGtlz6iKXXFn+Z6hg/6BMexiVCWMcfE1IxnZc6tovyxu
5rTNT1cOyeXvTUxbkZueCFhYzTcbyd57d1QqOzuFpYSq3F2IZ8+cVjU6AXZCPmrUyvmlnB76wvLA
fjzvIjhvBs37zqBMoFCT9yaobXLlYE8mol8J2Jp0f+WbqWFWkX2EFSxowJIV0ym639Kt9J/n0+q0
zkc8Bzp2ptQ+HrxnBCQd3n29rHrmJ1QNZEdli7+WDIWHP5Ht1EUefBp0AHZx9eCE9YAii/wTlKc2
I+2s3RoEys/cVYjq1Gg04PZhZfz5oX4aCy65A2lRY0/n2swMKBqqI89vNsHIG/d9LTo9/z92/PBZ
+Pv1ykeQvngeiKuPLif9dfQMuLGI0HzBLW2FE+6TRIEYZ79jinilh+YgvLYjI1a4ukxGx1ch+1XM
1X5Trfah7af78UWabdTuM1yNUzprW89m3I4Mw4hjuqNQR1IwYoiwXw69bTakcz6DhVUFsaBTnvQf
8dXNkywWdekYn7IuHJPunmVRIZI4o973wW4CvCvSXtXJl+180czaxv9QtPnJgJuWOIGjOgAJeSVy
NNYFAw09ooFbF8xCiozTe2Sld0GDmo924JqUf1ceOvQ/fzObcmQzcwrCwQyWaG992Jdm2YMwDNn+
HE+G8h22ZqgqctwidffaU50l6jj1amUTsSJH3CAmbLa1jlqho1W7d2Pv6z8bU2wJ4Tz/BYs+pigy
ua5Y7bkowKN3O+ynsJnJauSOG448Nu9V1X+14nIdihnW53/IupRARUE8Emf5hw6oxJMdp0GHHatL
juvecvSHUi0uSSzMuY1Vk6VhNLOFkWxeBCBW6qPvsQ4WNdj1qyRh+Da4Tx0ihjJDzXybw0q5bbo8
mOOVp5ECzROuTA83ngfZQMPJsfFKuuEYY+lyrOIFHsKMhrsUyuOHltHQcbhw4ASvLVsBt2h8jlE2
yGf9U8PYcmuyFV0pWuxK+0oBs7n4HFz7vmO4AUbaQJ+7mCdtJF2+DUIlMjbPWoyyEWoW2z3udD53
TwTaiI8a6uGsgSV1JvPKTkKpzr2i2U9lwMKS2C87475Ev7Yh31Azy8qO8ntZtzvDG/ivGUJZ93Of
E42mBFJNij2iBR+FNiKSQjIXYjvv18rOjsOG00QbR8lDBowSWQOqE/mS46Gfq7NykNwt9DcQ/kzV
jcLgf4HCiiLq69VY1/pNfW2kh2wNTztdSaiXBDzzAnnDv+sUlorRKsdFFCVLf8xoheHYe1pYAn3C
XapQeSNLr0iHMXJsBmdOCzIMZ9lw+mjuUTcjTQ+NkPW3C6ESErnVL1zv3RCUwchyhBTXYl+Xnf52
qYLgcJQH0vHzYmcuFf5a58lAiNljp6pAUkYxagC8nEFge3gmGg0MhuNj0oQEivAaACdc4Fex4AjW
zMXGsJOURqJUJfHRmCpbKmu0dP3xEAiPMSQq4+4vUGkpwC6l/Zj7FCN+Hh6/bCXmmuph0572hJ2I
O3jXS3BXRn700tcgAFzBmKKmKQRrMT0xTBeu1a7g+depo3a9KbhBbbrdENgCvb5aM/mjPL7PIh63
GP2yYNbYlUu2Rrh9Y6WHdLfuAoVrq1BWn6ciDL90a1hEoR1ekzeknr9hlFVVBcLCEjke/ApNL3Nq
kqhRAX/d3lSlMb2NPYO4/mM5C9zq430exeDKCpFMuikiVkRPCjRN2QJwPmdCgNHiDK8kzwclFhZQ
sty8XK+eOHPoGbLwU5n1QDdN+QLcojFWX1T0a0hANHJl7inzkf0P7SkdwpXCJlEQkcaxo3WdFFAy
JxSRTnKeGdi11E8YkL04wDOb/Wf8+Caq+DqDf/2oWKGbjSQsIELx0OXfLm4aTVca2b5bJSL7XL0a
9oEdWW3GdiMxPCD2TEt6JdZCTct/SShtaMtZCioBbPCOP1O04ON3abdwWRBGK72kV8nuRYJZby/h
QQCsYYLZ2FYsT52eDQ/thJVFUC9quxuCutBEtf9UWbmRJAmEiPJHmESeFf31WUPiT9WOSRIar9Rx
jaJQRJKBF/Vx2bagiTt43Y3frH/916018qkMHM6ACThyLmu7/j9c3FANvdemT2AUo+P4jBMiH0Lk
6LTMfgK36nzNG31xT8X8ezLQ5LBbC63GtAYihjlOwIb6vuCvlWdpWOT1Le1Y2qHeQu7YbQU4xM8E
yOtlf7UG2R9O2B7i8s9BkUq7NlSzkjtEDDO1IkK5iUSx88s10vfRuGm8PAzX3y/An/Jxwx9dmQWr
4rjsUh/yp3zEmnpqqKPdg8Jd4Bnu4JQ5Hn2YSdOZgbW/iwpngfFyL58zuS9gpor1hXwLgcvHj338
SCBlJpECPSmXfVKnoxevEFymQkUDvlVt8t0ZcpjNvm3v0IrTzPZS2lgQJOPOtijhpb25INn0xv9r
9U404FPL/6uGNsxkyTXI3VoW1TXvcQr33XWhPJKgCEqJSat0rKNPt5i088uUioYdmuUHHy3QU7k6
8YlLm0BNE6NtMHUOLlX4/kS7/qmKjWTDTb7CtgxHMavdeEHQjzqg1QA57L7/QS0vZu5HniWujXr2
gqyc2gN+63EnidZagIu/RetzFE/inSrIL2nKWf4R3jtPMDj2ZzDdlXPJK+BKZZyIvbvSUQm+t0BE
w5d7hPdHBC9ZQtuzaEn9S1RDhwRpOaKxzr9OAiHd7XLLuRt1Ytm7oXjN2k4en/XOmbcJhQ9+EQjb
S7XRvs6IoCI69nCZuLYVndSdSOlWbpNnKdvt9hk3KNDvT0FIPEEyzwhbUhL4CU8mBvEWo8Nroa2Z
bcwUAfW47Z/dQQSNs96bzmVSV/hhBf1D3O4F96yUGKP9/pZyKyiqF8/f7CPY3OsKlDmtASku6dLD
BH6/mRWurbBCeCXURtE3XLOonrmH69G2CgsRS5uF+qJchfhPCF1AvTiVjFHUMJyXtSpjAdf4MWQC
8YXUwO3XQRfGEBsk1MM0NeernGNz80MS/z7T1IKJWpIsKSmOtT7yEH7PB/v0Sjh7fW0Rgwsi4Uc9
2BDctQlyH2IvWcpdpKjNFlXE7FbheyiVwfAwR+3Jwv7SQB9Qc1pvsiZu1MA4e0OE9Vc0hkwFeByg
VZATV59IdXAutq4CNXIU75LiLCLLVX0WIILINrwTstFo3I+QwuGBiCQjUqTXf+3iG9W3aORYWvyC
Nqoxpcx9Osjl2UVKh8++gBZKkwvT43gleJesUh9LsnSxBWEmBxSObp6jMH341wblCcJDxPoVxHqf
+pK6fZyoDPEDismjQ0by+jnhfS0NdYmSlc9tlWFNIwD6k2HX8rUk8Zl6QP9f2fZXN0pU4dY3Xo3h
WjUQ4q04/Xunp+Z/ilAoaFEZBlqFI+gth8E6VTOToTyBWZPKHHw0C8OH/IbbnNEG296JRQN2ocK3
khU1ZiojyV+QsEWtSOFczuziBVeKntPE9uPRruvO1Zswed4RKfKiKgRMCum0iOFNEMHsvmkjKFBY
6yRhTORsSXG3fzqerFJ1JiGAiZWbWuYLIElDNYPRpfcDQJJS7LjnRHEdMpWCf8CnC1JTLDib7PH0
9gq8rLPWyiTDzGZVRXfrA9ntg8WQZQNsar1vuoRUgGN7SDYp+LgWShoPeLv6urfHNFXidYN4bPla
Gl/fZYxCHuh0EAVLgslWzWPxMPm2iCj3ha+C1db7yaEc+BGV+799VHqxzUwLnLffVynLb95XPs3B
niSW7ZdlkUZKN0wxRcgwNDRUUXAaHiVEX5Plcsd/q+ySCXhRQgfRca533cS1e2G4R0vAjC+qYlEU
0cy2BkPtZeVgqyfWPLxH71EE5ndcZiy0CiBSY55csL10OuHGb/NNwJ+KZFsRmYr3rE9OU6mJLZUW
qtIxfpB71Xg6dJxTu9MPVC4jsh44ZdKmo70JtdnoqGQIWqHJ71EeO7KtzNfl8aEH7lOPkcKzE1NV
2RRCVJmAdntI4Qfl6nzHFr3uq1dsswkV4+0T62RsKL4077D5YQf6d8Tc27R5VEDtT63wU69Fjayl
5nmya8lK+fXwNobIXh+l8F2WZ+GUAlVnfYVfmpPXS55vsIzkraTdFlAV228TcR40cAVVOCzp1Zv4
YCDLmNsGMgHqaUP6L1PBRZSxfTgtzCfeuSakBkVDwjrkdm9bVsO9lQroYYnKo+V2KxAvWmEF3O8t
JqSDHWPBPNxRoIWskzFixRsFNBvR5kkvphSmcB45TrGwSAAE3hCVmMqEpFx5aC2D8iJ62y6GPtY3
ljdZEmR83hjV029gAElScW5uA//O8/n/yEngeXCqN96+E6EjkECPijKxvmiKq8PlheaS+Tb5YEs9
NcuVBcNw9qmQImEAjAMMN8c6Qyuxl1hWefPP1ptx4TiaXfgjXMMhQ1jdYonUTmAv/uMve8Nvh9FV
UBXHvVok9LsYtDEQpY7SChJKmi3x58rFhckkSyBMNUgjSrXuSHtCNya4uyslO/uMZoJBqB9ER/TO
piakSrYDaq0vhbR41wtrHge8mFV8Bp1gXkm07wRSoCCYxDdocTHdTN7RtQHAFmPvr+abWJsb4ezp
3rMecPPjFwqS1PVFA2KYOhkTMVa2STpoy+gmOFk/mjYe9TZc6gNyk2QGn3a2O1KtNivGH+atUYfZ
M9ZCg1/CBXeSPVg5+X1as9uGvVctm/vvXX2bomPj6TK2le7vdQNH4a7F8wYECWOCAX7vMiC/i/qN
g06x48W/g9eujmmMWBzAyHLVR7Xw0mmY+g0wAS7mM8YhIk0YgBexf/s0hW64tb+Oh0VqsT+4QqbL
Tisv5DfKGhpm+OPmAscd3VfIYP9q++C9HC4WjC0kYO0TvCOzpBjxa5icFKu2KB+6qdhsYIExGt+R
mVCr3rBGdkNlP1zKAr19tcPGcwZBSoTAFtqcgXi7yK5na/sd5CaG/6kLnclVSooHCwuVkD1KVly+
fxsro97CuE35baCTCmHUlsc1rTIA20TuP1EB9k28wAUgTqPwqda8876X3jY9pxXVOanw2C5ja3nM
K/o56PcjMcbUxRy+nObljIi8/yVEM7JxhKCCB5pcaldCulJNgQ3/yvyP9hFl2+DfNnEmXyhUPQ92
fx6RQk0wG2bD6alw8KyvAPcs8HoDAGpPWykezt/2C25UCkrNgJEP73Kch3XJ35Lkw8hywv5Jt7S4
egFxt7B4+Da5oH/qIl6bxXJM9LH6rd/ZaRSl+8id/8Ag5YcSI0OS/g87slF2ddiuhkhcS3+K4hpQ
0nuCTH1maySuRFQHuAvCHThgJ9+stTFNBS713U90h6nxPz/XRZtacqp+1aH86edFyXk7UhZ/hCLY
cccYccXkoUlKeV2gciat4uyKz0bsa+yaxqi4zjmjgW2jrTgmVLYDAd6qqgCGqQ8JRvYClsWevgN9
auOQWjPhqODaHNQbbPOEfAxgDoL1xlfJZ3QcqvlXqN3tIu8KKHXpfGrNQBaD+22TDPopFI3Lz4/f
jQ7ubT6QVl4ci1F1i3TT0B+BuIIS2Tl5myZKgSWgALYMbpHcu8U3AAPCOL2Y0duMYGzsZZRANxV9
fJeHF8iP6/h3yJgQbp7tbe7tz56hZtxxCbdQZe/bD2MEf0MZtCVKmNCR7l9rtJJrhE7VIRyR34Cs
SICHlOsj+9vdnZ9i4aIRNgkZC7Mv6O/oqldA0WgoZ+MslPWj5v5evJfT9Ex+yBTVKAL+63JN7J2I
wqSFZNyC3Uc9WNo7tgg6OsHbcubaWC505sAjLnQt2mt6yhZsfGR8m45pXpV4e/Z8bC0YSIxkZfxA
ogH2jHCrh6TP84unt3u4BhE5cKOFnigW5m2s3WMnivQgbEx0taKyyZ1wC5yMMSj+a0ehrjcDtKAN
V+VfnpY0lFihLzHZGkSm/EiAJBKbWfpys+kUmHpUmXKpgjoE2llu4C865XN9XVWuDU+Uuz5jZzMU
NdzltySXKrTVEQey+PhLt+Xs+ipSwuemjGAV5pZwIJea/E26+qa+bRDv4AOxjD/NhTcbKOMUy/o/
x5XZ8IjWdlS874Adnl0ZNqnkgEsxpXGjzfGwBOfeJC/4Y9SAv7yDqqWoQUxUh1ARUOfvG0Yo5rBl
+axw8sDJ5YKZ2HL7oyyLubQii/IY/T5i10VyQMmHFWEl5Rkm4bcKztTkfDOmgqQvX2N9b/jFHeDw
dNVhKwkjp0jI/tnQs6FHHM8+xSG715VeQWWpK3jP1rz6CQ9Rakw3Ya9QXwAkaZxlSdMRgc84i+M6
VqYzH4QkKqVlzlDTfGwp2OQJPEmC0PajaKMWE5p4ilYdRCXxjfJqrKdLxZ6MUE2Exc4Evhqscjl/
SsCjZi8zKyHz8JxQU1j05mXY++lulA7G+tofX4NsfMEd7shQ5SLZH7C9sm2EGoGOEhIaP5+KenSM
ylSsXw2uDMieb3i/lBE9ywTdZxEJcdl14AZb2+idPCx9Zp94s1s4jtyGEP3sgRzWvMIJBi0xf4yF
ctN5ZdxjBfdup9UH91bCKyHoRBUDXw5MAWLFAgSPKxfK0rXGXAynnQ+tJuXYOSqKAqPxD4BtvGJH
5lOLPeemgY/C5VnQTznE9f+xxej7OCv9ve6q3BVS7KvO/RRDFG3UzROPFqw475XTf9G5EgpYCUwP
JgtvrIcD47BCveA89scjAk0k0K9RKzp2j7uZkHM5YbtzXGdNGh3r0H9+D/QSdm13NAtYo5EeY140
xcpVRC7+pUcdndGKaLejqKbXKfKQ8fkYw/cTbvcqPAfKgjLdkTnwX80rRJ3rZqa+oc+sYUNNg9+y
j0yMU8W2Kr0ruOfRhHjtgmwQEsUIl7CwXVV5i9EediE4jkI9glLLVzNMVauWxQclzj8d3PQ2LdtZ
bRhO4NNul9VtdlpOw2/ojxfmKtBVwurNu9fbBAB7ki3sARHyxVqzOceLmYV31tweUJX0BuO1SGAk
M4Z8TFEEjUZRXRAxvRzeNwtlQXyrjM14amZsode8ObGPqyGtO/lNWjfXUeB7uf7UrE65WXEcvpGS
OaUbOAZXkqp7T2VnXS1XYhpzv060MqdYsTSr5b+mGgwick6BcFyADvmkImQGBSTqNMY5dpk9uNj3
I4caS9puIWrNCpXv5ZSfTtE4qF+Uww3kvthS3G1lciKaLTOj3IAGVh8OJGzf+FbdQVs/BJH3F132
1Z5lxDrpjpfpFzGz4ZWUVeUQE9Aoz8IaJzdYkohar4sySsIrvICjonj20mB5GNo+0ZXCz+Na1JHa
nbsQ7DlgR56OoLNkLsnMWmxLlA/FKB6hPyo/TU4QCfuGyNokLCutmePTVRK6pdJ0350to6srEap3
9tC5DDG2zEsilW1Nv0cXVp9k/ArXsiSiXAhtfiE11tRHk3Vfivbhuzc5md8eVD5szbyjBJblwG08
b8RdqqmuAQjdhTFD/8u0FlK1wv0dxqDbdZ/bS0sFZYPCNtrr1xNrJHK2NWlcYoZiqy3T13yw7Zuh
4/0C20dnmwYspM4G+dqKwlQbn8b9/hsCQrpn9eSITvF/q2az9aTRF51ZS8jA1x9VKSTTljx1f0pp
ssK9FQ0EtLkaA7qF8+FKMTnklKA8TyuQqE8Olh+pvaHfqnDuISSlohQt0gmNxsooxSqYv15CWa/8
PYHv7SieZt8BsTM/atsqyvBhcuHyU3S1IjDLdKYS2OfmQHttpW9t2/Lpcb3g/JffhZc7YINQy0qa
GlHedKoYqlXbS9g13Dvq+lfDxBFDYeUnXrlxjxQgyOK997lV1Tfv5GRapgjk62hBOmNCmHorQaU+
OSXXiou9pCEnkMHVZroN6ElFFbFMzx1q4GmrcBsUn/j5qvI20c2pas78bPgbcouHF7vl3VhbJDDh
Djvao/o+PcoYFq34+5A6NCKtKKg9F/of1mIzwEmuvNyX4eFAeM/2v7l8hk53+dmsh2JvUtWtf/H3
040fdFabByF+jxK8TJRCrTDzjmdWnWbOM+Wzx/5YZT9xmELRZsrt01bwYiXbQpkEOPdlSUqt0XwI
i6xuq40E8R4evA4Y4Vg5tzshhVDXmvw4CnFMvlTlkOOjBhXxF/lptC7p60fAmTDzKJM6c2PLja9m
x5uCtNbLU5tpgwqvjE+8SPiXgHzUEjmeS6PT5ntW35h0NKVohXDoEQUnQ//4evqVh9HxAzqDmbWT
a3cP6vEQQLGPk/17zF3echpu+IZA7TQaKNDnUEtVUZAV/Vgpq+3Cl0A/qrMa67R15C1rtqdyluXt
ygU844+NUYTRrzItSXrJ91sbFwJTWSYoFhHXXznnszFx/RdlI79dmzuQEH40KpG+OkP1KclBE5pa
nbRTw6OhDeTn6My480mRlBVd16YXJviutasazI6GXhcoFIIFy7Yh8RwM7TVXE63AIUMCEDC4gpWN
4XRUtm+s02dBfyVCUmn9YmQyr99I9Ww3G7CEdcDO2D6c1kdsq3m8zkg4hLWakSQ+Hotr0dB5OnFQ
Ix91YbPtzHFRUdpB/KBahiplRLSeqD+Ia7qbtL6KQExXCXkTFUOHVD7WVsKgtr+jblkMuNw6mNfH
lBVjkjPxsbR5nPK3hakhYNMkj0F27yuNtBOYRaQuMYabk8lMIqu8zl1rkNuHz+ur5XX433Wzav4g
k4y5aFoIfYgAXJIjnvT2Vp4oSg0SabvvMMJhyf9TB6v1suzmuw5DDV+4Lyuj+iSUBaDAXEA241w1
zm9i2W8fvkOP1cuCOSRdy5UN1WCr/g/JICf0jPSyxmj94u9k1T7EgUqwCz4F8B+8PxAz5kajPwte
Kd+jm+QIDBGou57C5JgyPRsPf+UvMwYXePiz/eLCH67ueFOYBmvukBnr2UZ/KjzqAShCzoQD3CUT
YF3mB4AUWT9LFTBDP+d5wuWQAGYwcvS6XNiVM9tC7RsLn+tSUxcAq/fevRNv04oBaoKra9KeXC92
hqt8fO2EdEJail/JQC9OLAWau3E6I14qilIeb3mVkk/j3Zwzn3Pov0FP1iblaxYtBzI7gmJhzuOC
fN4T9bDmfOaPyBkSpaPlkw2fYmgbr2+UkdlgQxkVBJgFzxV0JmSJu7BRvBe8MO94tiOu3DTrYayI
kx2pKe3zMRaDHhrVV2yfokMbk9FhdsfAF7CQff8ai8ncQVgjhRXRrDxxjObDTnWq3mCh0AqVJmnS
UeF/EoSb0QVFYIO+OQF62RB78AoD/isa8vMwcCMFSO9rbeXEM8K5RWgI9K412/c5Ud7OugEKNa6v
aSGqe0JcRJ+Rmma0nXzHm2zJ9/hTEhx0ZDQyo6aLAg6lNzSsrXmrsmB+rDVgrtCtbcW+j0YHyeSl
dOCvv3EmjgR+SHqaM3sk77ZLxZvZV/ODkJ/yihJc5DBrfma0X4oS0kqC15qaEuqL7pvOV1FYCW8H
81N8LqS56HqfN/dNsvIjR/wwHMPSEOgzXlVXgpCbzGhikQeh2Kntp5jegCmSKRfZNeBjKEjAOmlD
HzofSwFiEV/exG/nRLE33AjYZILf8ZRUbrUhfgB3oHXiijPYE0bI0nIDJfjzJB9mwaEa8fJxGyJJ
EBxGlLS8DNWHN+20nEmi8I0jHWv6UAqlSE/fL4VQZVY/+n3mgc/ci23tv4atFaFexcONaYsUcfA/
Oojalc7+gmDc3kN8q2z1ZDDZlf7obOimIoz/3u6jl/iY4R/4QWFVc/o5xBwoPBm0Qr9x7vpRSMzw
m8GEOwz8SDMVKaHY4TzcbFBJtfhu28/a4cQ/T+PsLYPALkCumoR1zyBWWSEjJB45UCnJ8yz1fdDz
DUn45ksPVFercTuOeXXcVDhVs2LoPRK7NvKkbT1TQR8HHvLHEfOHul9imCfjfYQznPG/8Prsn8ca
rqw3zsK/dniuoCnb7Xsf1YK1hVs9oyOLqa9Gb1me0cAYvHtfwRAdHrwpDuNYJAHFFifyDvCc9hjT
kLwsGAmFyUnfi+7mng6how6SdVTQyZ/g180bj2mhr8PAmIGtTlg/9UuEYJLr96BmDBrbXQT2bYlu
YSxc1cB+xJXMXlQjm/kkfDoSWetuZ85rIE2UgtOuWsoPrdsBKEGHqV2gKlbfkhlG2Q/ObAhndVrU
dsPEYIGADkfGDwaumvvH2KmrHvTEi6P1wpPLVs7515RGjyuIC1iZyuDwmP5n22L31vvWknJrJnUl
+w/Ml43DXXzRH9cXfwEkjeVhvQNfpGTaXDkewfRbSDOhnri+rgEkGWEGHzkFzPX7dpdSc7uSQaM1
VfVd0fNm7fogK4KBr/bcbbMJHpWqfa8UzRRPKcZIdinBvbwin5u9jf1I7hfCSMXTMOexN9HM0RTs
cmwxatHBAQLLEM/lVS2aK+q93BsoubREsUa3gQvxRa/sY8EZipDLpBksnPYo/1xuBKH1k7tPCJBS
FKLz2pV3IejRCtQKo+15cz77MZylHCnKow4t6tz+lMXplpMN7EdcWTPVma6V902KV9tRnZLgTLQJ
sBO4Xj+/1E09L67b5nbzPnWrgHCciez4OQF/6VLx9hle585x+ny2Z/LADFV8PqcIpXD2BTSa2MJ1
GLBa7Vo++wjXlIKrS2qmql9eySmkjOVpgPfuXlw1q8BXzWx82kA4/ZeZ5NGf3r9kUH7ap4eEP7aT
nAz0uqMRuv2TWAFPJiiJptxT45kgxXQ7N6GGZjFqvaOogRXMpYknWVUxC4+O6zJIxkfvPgXfeX4U
LnXdcXR8UNm3QBz4oyo0IzRVZjKdwakMiM4G96gp5fcg63K53QUfH6U9iidszWmeQgfTY9zLX3OK
n6Y96//Rqo+EC+dNgBwXPgxJ4MvgIdaAoS5tr2Zoqj/rxOzh7foQZksX2vNpUPwEzFjrtstQH6bf
QrDONYwQyUc3OAqPVwiq6+XGLMAi1TGrq8dkrovC6qzMeVR/Vh4IPTPPIH3uUNtBvCftTyfVRDbQ
J9riwgZmwEUEm7Q6bAs5eV+0QJh1yEwT1v9rIG1Q9Oi0te85bda3vHjshv41UzwAxuHLlfp2Ipwt
QA1Ghjpm+PvtLL0nMD+AVISxeggpSQ8k5MOznRJj3Zvq7tALXlbJgOYmnWn5GMoE9zNp2RkYIF+/
uSsbmeAAoysVmm28sJQgB1ewStV0WBFvJW93OdJBM6TYKPcm2W4vmRXJhmIJTfwoNW4MX1nqRXnu
M9VNr/vHSYabEMGkUY1y+986JeLv1Lm5drZPlx3t45LhL2p5DHtdeiWMJ2pyGD19srYFB1kt3r5D
+gQV7htojMk9LDcxtKOBf6gD9lV6aKnWNhAfFXEqip3JD7pyuYPZoYpxk0QgxtWaStwNou4POSBU
lkc4DHla7/NtUsnt3vf644ATd686PHAjdJcAXgeknedtlYn5kG4xNzOYhr3sxFAoMygHDFIRi5ha
1PWf2K4t2yEmeE8WF07CHboG31pQtrBp0ILSgi56RL1q5j7zRJ0igVDbP5dXjO3vLSIfFBtH0SEP
yZZPUqvny6DxSZ6gN04Y7gY/W4DwgCylbSiP6ZMYHMvN+gmdVcfH3GVV8ppkwgQvGCzzl2VIpdvj
DgiE5SSOFxmJrLDlsi9zXnvfT8hP0tAUULhIN8LOgyer9phyS0b0xxz2b4G7EaNJdlsX1X4k5jx5
d31FhAq2htJDVPPIc30fhjbvQYS+Ck+wWOL+0mLSGyVQA1UqzoWzUcWOyMtIrZqREXKBgTx3eEmD
qdCUOo9Uwd8IcRm5594BNxZoQmyG1w/yZICYg1wZE+1RxcFktF/Akx+OdsmKg98OPHnUTZg4/mfg
hIuUg3Vw+GwBPAcXGw58SwFYVreAagVGD2///BJoXzgBtz7BAfM9IX3ihOUhflWuh387TVuSIwTU
38JsGArojed7d4ltmMNwPT/2I96FSJO9HSEWip0fPGSubE610g0IG16RGSHSd2sbvj/stVhfvu0t
0+uxbjNmiDX2+pQ2aPWY8trfOWVlTLOr4AjtOlkNjdoSFvTcdzOhH95MI8X7W3G5irXBxy9O4mh5
iEc4xV6GtyefBKG58nBN59R6uQHxykCtfa8hn7a0a2EdtS/QXvuwjXPLAy6u2FcuuD4Dd1v2KP1h
L6HjXzblYDTIaVdRX6//4bvi+6cDDPNAN12kVJY1uR9MFkX0JijF9v9I8AYzswAwKnXeXfFnVdeK
zieHwFTDmgNnzDQ5Bsrj4x9SOZP7Qm9dduqg6yswYkcnKUBnqiPNetc+YhxIygvb5gW0TcMNfXgH
5mpfHfV+tyNfCm+5vENw267L8PgrsRlu/wQ0nSDnS98AtPa1MsfpmhJ2MkpyrjNPxBUYVhTIEbu1
0m0ddKr9foNDHpBVKGklkXn4vleCSIIlLJCGvcQpp1jhgHaqbjLFHGlyQQvb+VGjU5hw8QBQnJvN
V5WsjdjeJ4/KQFJ12Oo5fXrLE1mCM8I7A4Nu9R/PHRTlnaKKnaGdgWG+uAgqY6jaD40m8LdG0X4u
5eIFvo75XhxNEx2EE3vWtMgJOHrds+EzmR86pDtcY/BYiUZe1S3aRh6zuSZr2kDKz6iqk7EHu/CN
2ZK7rhEtZh1oBYNNWh6dvEVHXWRbNAoWOcbjDChQJWM6JPb3qhDsDPBFEeR1oPElVSHOVW64uCE6
j+dNW00clStQOjWoxraH0X8vdces/4pvEgF3eza7WZ+ESfi8YQDANBrhtnbr1u4bTgPHVpFnyT40
nNlyVdKxRqDjVHpoasYdyxMLbaBFkN7n+JoqOQJLNZ6FBBeRLAau8iujjuHtG1apyARiQ8E+1Tq8
tXewQ99yh1sxkvwEdn/9ISjz17yc0Ucn+kB5hKrFHg7XwlJQAQDuULgjUhIZB+gk75Z5WSMmHreO
E2/jRf+8P2DabKvnMvaOpguDZf5EkdlCmzAv1KHhmya83ZopJhY4P2Iw9ng19DKre8phViTG9KbK
FnzondlfHbv3oXEYHS7eGz4jmeG1dVGbIcHcGrqzx/7u08vhi8SLgh9DmFbU0hC9SqEpAkNhTDND
GIP6Zv/7htFEdrhB6z8nQt5usgwLoJv6mIO+IQkcgRIOrQXf2xcfEsLV2ljugm4XSLyGO2akGmgh
kHwuE8Sjh5si6WHIw7pZybDU/xDU4TQqM4YMUAw9icoeKGMncok+X5ULnbfu+IV748jQg4qizvR2
sphF7bW+U3G+cWDT3FJjF8ApCzeG40ljOGj7HtiuScT+FRaVyIYVFcKT5W6dM8WXOFlOTr5wZ4k1
I7Fh0Gj078i4RPP6sAiKHa9F6YHZI68CLhc4wKCPKaA5FYRZ37ycPyXDqiI9c1SJtM1dS57eoEHJ
5P6AlhlzJPT0g+Cxs4e8Ht/VTzLPIddFrFmius8uvraKLTPraCfr/mQUZVQK6EsAWYfVJsf5I+W1
oyM85yEErg52pt/vyHcUYyscbJokb6zTzvXiboTqR4Atu7PTYKP2kkDLLF9DJFmok5lGzyxeITg2
02lFOdxcBprieadHSqu34u0ig5xB/taHz4RKyBOUvjWFpc80PoUfh/s3JA78Sz2iiPDiVxO68d8s
1bL7o65XmmdMqi93WmdQmsW6mIwzsC9cCjU2ZvS+RzP6dsJjCXkWGCO6Plv75A/Ul3IRbkfPmAsQ
xcr/rhs2fmBhV9Fb+ZO1/oHpiKPOSjehVShv4IdKjwb+w8f+82ieXERVvoKFRa6naJsFdvxwEwCN
GfDib6mSY2lAEcXrRjFagvR027RBG60Z9Jgz7dXNx+Lvltkc9DJhQt3SzJ95sRXQCRKsh//BLCc1
Qe2q92uk62QAGo7xXaxwryr91MFNez7FgLMVJNBZ1UfvHEZtQKAXoTLN3hbdGiSSd2r31s3VBNC5
HOnusDmYXz2UwUKk8XePRluDdlGGluAd1mqQr9mJjgNiT0z++vmmIj7nA2YJbC9MR2T8+X9cBBCd
ir42LwuYu2Vq81fNewPvmamyUJfgFRbrlgLH+7PvKiv7qlvMuffFZL7QqQKLLaXa2KRzqI7ozdj6
ehwJK0VVCEkhZH5q3iqmt3A8+8AEk6JCNTq3qXTk8wrVGPioUL19aYXNbEJ/YINTuc5ThWJJKAga
54XiEbmyD+Bj3OKlPQrOiXX3Sm3ULAF2uXVga9lW8u/gPJwIV1Yv3oV9ScIA3iBdNJbEmIeArumv
oyEQTEyv9fNCGAxRJV+nZfJAM5Kty6ShQs1Dq0oiSL0JO+WzwBa0fQCKQb+XaocVkGZ82nsflihw
v9QDNOdsAF7Pf//NT7b5VFCsU3/VIKZDakpufuImc4YIPhL51ju/qLIKgUMY9+eZSccSou91/9B7
AvJ+8yr5W0YeYtNf6ewEptuu88OawgFje10t+NlIY5exonUlJmAZydmyRMEJYIaj0zZgzu62xy2c
BZDJ2anZ2lIeVWwzFU+ipunVUBlep0J3iCE+aMsM+hM8+Wobe23sQ/oUCmgk4ZeBVfXRtt4ND7iO
8eRikJazKQLBAVf76l7aFZlA2UvP0mFhOD66qw9ukoKW2LVJY2NFMwGZYxQme+2joAQ77Yo51KT0
6/vg14yOQ2NjNUGofy8r3hT0+Ss0zCrcrtmDZZ3BD7Kjw5+yvdJlq/BvBkzLVmzJ2AoEJMSMrCfJ
/mah7qSgB4RYVA0oaV9L/zPkOI1RKlt3cjTYLf+91K0VNzSFGsw1lslPWzPJJPNjhLEwslWdkl/j
LyMY4Q80izy9Hvzs6jFfAyXd/9AeIy/2pLfqriA4/ICb0RI7yRyrxjOvBvfP6mpD2DI5ANjlF14s
wk03F/n/eX7Z2dkTl3NuZ5Y/Ko9UodYT6IaHq6mfGhR6W7+y7/qPRZvr8ciYzfkoTF2YCFmBrmAB
xGxoUKZ7YAPoD8LmcTicIKhZ3tj7RDr1RsD1FTdgs4ELQ9DH3pd0RJiKxAwIndAWWgxVDe3uq9pO
M192HhAPH106aQ0T1H6ipdXHOy8i1gBXp8SEoE4Rj+NFBApWtmWPg83e95FsfbXcUiawsFf7jNcA
mtQdLJ5BeYMubvLa9CJJ2Mgk0b+5jemhoI6Hg8938trLekEpss2JzKaaUbusz6siD3qALrcXrVxl
T8lpLrTbRltnPomDg13XMa4uVtdNXED5q2VDm+2mTRMNe/yMhgiTOmG6Jg7l1Ux7zpmYitRnbQTC
X/fvXCz/MPm53wD4Z+AP3dR2ZgA9zO9R4IWI2YYaRNKxJ0Ca40feI2NJoWm4frtGHbQZ9CfTdDxL
KcaTXoktCJTB49Lm6PJpYUqN4pj08KUCAlu7mfVND5/6hlGUHRm1dBtEYF4tNZGCd6GB9DPnlm6m
xsnTQs9S9D0VmU16yttLD3DujcWaDwjxpUoBl/2Rw58nGny0wLVY1Z3Wjy6y/eQteFd4yZVLxiHV
DvjUkFQVVZVHPq8H+e1D23IqnVIKrWOd4PilAkalwSyumFMIux3+xnlP/jvw4CsUImZMO7/1qUg3
DTr36a73nfFPXNFvBBT2e++BWlvkqreuwhoPIjnFdTttqPxjXcBGh9PjEfXAoDImOVOeidQEQoER
ex7R+o1sEcpq95/FNHhH0woPPB5h9nXc6mQHfg8OBZEPOg6nl92FYzMVxJbQRuT6Ut/JG8I6CG6w
rhEsIskso6iQQ+vx2GCdEASOvqHGOh5HG9KYJtzaWBNgcEyN7CcpjvHY9ZcPxNgQ+FKRodY31pI0
sKxWbbtUl5EYuceog+kjep7LaPVqwo3vuExbBV82oa2/faHoRu82TWb8TJn9TgCXxtOr2XgUY0B3
IjhPFRc4UNHsFDYkuIE2ZoWMQNU6lstjPqRgWxP47QRgBoFqhnukLdDQPUEAhem53IO6vudPW21T
QH/nJXUhmUP3PWX8Lppnd7WyVxcF+6QeGNNucu87TefuDwvPjCZwas4y8zdtm4XXQ4EO9mpMiC54
Wer5gxGI4ZdsxqgDT5uy9XR71zmhpo6k7pzvOwbgJNuvy+XadoBwNeb8K4sWUYOinvbzBbdTHJZt
nrnVVprYw8IwgKjqnf3Ci7qwqA/9EazwXRLl0Zlx665P9pMahthz3nXSkKmvbGcdMAnHNgRD8bMT
jXWOc6WjpsuPGgJK+X+vYk53qehxsp/qFzCgCXiLjHxbD+6cgvfK9lgIIdU0oPrEdMhxnxwy2XGy
NQ2ryQLWGjKDFXgxE6do7pi1XqOH4URPmG3zcYVPgUe9uPVY0ETEOEoHRN/yEBjM+e9Fij3+hPq3
Rya7w/Y0afHwGasQGGM/RbyME8dWflqylhkiaFi/sfI9rlv57C8U2bgVSiGYGRRNngxcT1clGjiC
CKQmxH1aZYy6HurGyggVb3YHiwHr9pEqSf/FW+STPSR9LdTSolZdkquUdIdlpN9sRFvCci8riPjk
fjUwIB5ac6hkIKji/w53CIlA8lLNq9M3+eJuejSMI5l+kYOq0MmDcUKaZo7QB6yaWw1y0/ik9ucn
aEt64Cycc0fU3HjcU2GybwHnRN/KNMDf/3ZZ6vcPiuIY2sTWrqpUh3lPDcCNdzjBBWyqd1qEfHI5
HfeYohBZVygX0PBY3MCn7ftTNWP3YS7htnlV84YE4KZzyzBgxQsan5AAkeRxiW4UxPmu0x9fCu1a
gjfAWj/9KYiyIcuyUA99Mh4GcMnUtW5OLGopszh8wyEnt9hTYIqK4f1q/kr2773CxSk4FPfCdPeb
InTDYKCz9zSYv9z3YFJOkutXA5aHNh0i4iDMwAtNTPUKUL0BSEg+KS4isN4hSAiVLdVlbyjYeeMZ
fKMciktdqgn9NF/2zVseBzz5l+kHOVX53QdPV0wre/2TON0IxaRkz6KnfptLk/Mwuv/IKXWRzFrG
sv+wUyHc8SRWRDZaF/wrGYbPGASYM9IdI0TwBayN56DXACNCLoBOg+Wbx1wb3tabMTDSYN3DiqxB
Q3PoAr4cpwJOW9NC2oQq2bcKEVM9OJMCBHJshZo1U/9oe+tEOEGup/4Sl+8OPxXOfV4XefYmzpG/
VmrxDusDZAlrHySi5XKLkQEnk2SRn9ikiA++T/nlbUXrHby9w867aWQPqtFJhZhE6LmZCiURZQVU
woBsIHBfosYSzD1MUev5rR6VOSpoLqX8NF0TzqYa0I/1Io7HKYv4YG/GNeCl4arbabbOX28bHwY4
wbZFs+aklBqw9tu6bLF3eIhsRCVNPJCRh0N+PVuaeYEf0Hr+On1rm686RpKum1CsWS7Qsgz76d3F
4XH/2w98mnTEXKuYerJhwmbiO6aiE9eVLs6vzE9cciFwcSZm+sa+AhFym1enQr2WCGz8u/mFDDqb
22PtfsocAfgzOhBM40nIRKNFMITo/sUVh0cF9lTr2a2J/BtgkYOQyq6zpsbN4UvgTj0ALT4zKa2z
9KSVb+FEueIAfRqp8/MfsM0NqhMNyuTOjMUFQ25hJnau+38cddilpJfBjyIi7QjumkyurmCBfc+7
S/dJ63UPEd9hGmeAbPhmPkGjqWKalYmz32peu24w9Q++7dngjO+s9DnzqebtPxvcNaXQiGlmaa1h
bXSKtm+2e/0aMNSzjN3VVHnnsgilPY7XCsHymEi8vRB+npEF9ygeTjNSni3mL0jL2Xw6nffTYr9b
B2meH29F0/qK5Z8knoed50FixB/HSZyN7Vki27q7gl4TGuEcxY+9guhvRpe46EyLC4SN/iU22foW
9uHlomrsvBtUS5Wus12ZMvQKmoyGxrn1ySNrzoaWOYbCw3GKGrVuGgnFklGDOvrfLUqBvpfYtPRK
3PI2EbgW9ZtJD1DGUC7qx++Tov395cXjjmnYQFZh/R6/P4cxtBKpvuCnUZzWyAd9S4wCztUj6Uj/
tQS5fBNC3gXp493liNVq5mD5VLRjihw5C0WHOabVAD4MzAAeB4I2N1C4XSHJh3H+8yB6O/iZ5mC0
/a1tB0MADwWGekXe67InWdJWPuUONgj2P01r05bHkhKkYx1DCWLiOSKqN+YYmRWjEdfPNdCaXk/2
aicSNKm1bKv5WZH60d22DtfqiEb7UxfIfN7Fy7k0M2IOS0WUyw/Dbk6DVFHA4f48ClGzmouCSryY
rUISX/f2HG+bVlKcf2WscErABzTI1v1fUkttt9CXU9eZdqIxmyI6s4sYGivwHODkE30K/P8pIoqC
WfvWuAR2xCtYX8tKcBcJhMU0fkOqMVYsS91vlBlK7F9Qx30Vuq+mrDQOd8Q62tE6ZP20DgrnF9oP
1mb3yI2R4irORW6nGCB2OlCmPd79n3346W0qEBUSapO02W9V38o2H7N5D00O/xVxN5ZNu0RmvPDB
a9jmsprn75rt5ngg8VkisuQuMOexMKmwVwWSznxcIJ7pXnO4NrETTa7eqV1BQ62GzHHvDoZE7Zr2
0zn/iZ5kUcGVjr74NYb7ozL8+Zk1QLBPS4jevVNXNZonFA2eXlvKJa5A5qVpcEEIaxnQL32IE64E
8oMdQsJc0h/YmehHOg2tarwLO/uhhExV1uzYBdGfuE7HPJFakgoKdlvXENpnnxUayuF3k1TSTgYl
66bm/PlQTqF2yg461zcJo6PGZMRNfPaZYE7IpbefINiRNZSs5GIxmIL9n4N2/ckakFOq3n8/o0Gu
UAULOpR5PoNKvfs1vSdgtGEPA3AzFL8+ougQuPbLXWdJJfpLLk/Ml6cLot639BYrh3qGVooJQ14n
WPin7xOFAN4lL38oS1CDoKZ/QmPfSTZwsMdOGeR+R+Mf5WX8YEl5h86Qdk5QMuAxITj0ADYU0LMH
mLRzCgT5EM4/Nag/V/Ed5xf5BHXj8xB4+Pyp7n3qi5nsxrxK7/2Ntjyw2GNeYYLG6c7mP1gNJj7C
1Zb1Q8W1d+9i99IPmW/djFVUIgZQRpx1MZ8H90zYB3nPI3CDWSeJECwXpEtuS3vii18HMPvG4BWZ
VXvGy35nMLi6flWklmbQu2crGRUuwDuMnVCmQq0u1UsRJaA+qzdkh/jfVF8TjmKRhSKSp9YztfYZ
Hy/7gEw+Acyk/1zXQWiFLbiJ+t11aN8abTCtssnoA/hwJ14LWen3hEbgZ4P8d0LxsMnhCp5tQa6n
lqheEadtfOtCZatxZpu5PRP1wc7LqdSAB77Djy72mFyyIrJuiGgEwEWOJo8OznoOKqtqxBFkZZn5
CkRjnYprF2j/wQlxIx9tVkj6A0QBQTdsqhcN+7Wb8nPdyPOwjPxzwOPbh1aqZzeY0C6CsCgq+D2B
H5aohPwClnHrnDyKAAsG0d01goEVlM6aVOa1yloOc7fN1wmuekKXvSj/i98ytaBlGxzOJO5Qv/vl
KaqFmgcQY2FmdnYpB1Z2aoZWZ+EJZXe2d1YRkDREttdCrCSUjaHaYDphdWoEYz9o5qQMYUPiPAvP
Z55/x4TrcMWSlAfYpmgAhBmVLN7a7PRNX5RgOkWybY2IuyJ+nZ+QSK1h8AXjhrmC/PzRIs+07P3n
wKxPsbelHf+v1/TNmdLjbHWc0IXkdFPQS+zK4YeQ7VBVfvsVA8bf4mdLn0nzg4hy69DihQypNpDr
RZ/TSAsKLNEof871nJ1eicmnTP7M0TMi2iQBQQf+Vue9Fhzw9Do3IYwUfAHSycR72nJuzLopCSIm
xHHg0tSop/WA67DbzBtaRogqBNy7x0I+ijww9Z3WwRux4qAvTW5rpJ1T5V/0aQAshurighbXcI2y
dJMQxynkxMeKRmNiE9pib5R2LWqVQZvYCZcrsTNs/3pOGgFQlqZWv0857v6tUoZC+txzmCu+5yT9
fDqXGgSDBp+k+EDhYAin0UCWx7VlZ8khA64Y+qz/AX/MN+gUspRoEUb9T9EhBOLf636hwRffCZ9h
Ot87oPEE0sMAT+U2pqgnYUFgP5QXRmnxQnMcYOgz2F7giyowRlYe1HbzQhTA7Kt2Ok9AjRpq02he
s3X/TDtUnb7PpzBjj6xBwBXxhxyYP9ls6mQ5ubQabynApPe6ExlAqbiIUTkkeGsxbS4c+H7X7xRf
ArtBkb5AEk7W5UlqFQYn3Ft6n68qEB+KldQIk5Gw+m9+ClguKGYHeQVGpbSjBO7e0INAWDjVgppm
u9/21Xl3kVVY+4UHIc/uWTIaT+LVh1Tn+2YMj0H+NOg15MsznNAShmlCZtzckGOUJVwpZnHwXCs5
MG+6Z4lGE6tz5VY87r0MomeI5OOXMtrL6C8vR/XT1YQyMrbLqSk+FJGxAg4bknlnNCfUR/t9SAR5
oOxs+k346dpqZLVegBhN7IA8HDKmSrgmAztkQmPlCWu1vCAImi2IDh7WoEHgQiyCF+p2SZFABJLf
vmVpupTb2GUA+kROWW2FspcLn1vltmuRN7fEWO783KOxhRQyi/bM92dILSA0nol1d6pFtPBL6TGH
fpOV1zsypmAFRFZnuRYvRTD0fTRPVTK6d3cbMNZXe0Y0IOwkjcTjRChJwNPxVr4LtuCt1kilWTjI
85a/MUwXLDwlNBcOVQFF+AWG3KhtBbuYTxCE9INNCx+bpgIwoayxQKUrXBGkw9fakmCBISjgi1cD
tls9/9WBlhBQKTp112r9rGdbUyk/zIzzrqXlETp6fzSUvBIbw+czdgRqR633eEbKAmpbYTi5J/bT
GrTw6zzqoauFZ1W0HtAkXPzOjYrfiO4tmqkglZzlhewlS/Z8hXBXwmZOOtb151DYEXAf2orJeOmh
4YmXU6NRPDx47vk/sIThDhyGVeKIapDue0tA8KTfZmF4kwKSbGRAoTanwJquU2Kos5pY0NgKY3gr
0qQjCbKW5GLbWe0INuuade5ieak2RA9mTUQ7XTH6Eowt//kpu8h4ow2JTHaNJD172S76e4FpA2RS
XXJ8UIdhWBs5bNXH6fDkXKoXzc1eUNtweoNctzPqPH0/2B6P8JJN4QDDBCJSL54xGKZbGhVGV1M9
6Njs0aUkkx9gzXhohI4tiTNSf1wbYf8ZQRPuHe9iJqwZsThrhcCM3hO2KJBoDziXZsDECgHgjcdl
8DCJ/TiC81cks+JSxHEjFA7TkfF5O2leiVecy73SFsIBjBVT8RPjiGlWiLxH/Dg6v2/R5YZL8iy5
H5c+q/DxowDKsYWjFhAAjk85C3WRSDCbqazTaM+z33jHIxz0ZiI+81UewCeoGeOx9CCxpUGRKh6U
tdn1nkU6pWN2SB7wF8Lz/0fCi5oXLDvUF8AxAWWuju1OfmRQHKX9sweTRL+ldVqUsy4X42tcInIS
36WD+k+bIksmZVG5vKMpJHmtU6De0GsBf/maISwo5GaddEEwrknikcNaquWI/BV3iV0/R9tsoRBO
spZXAHBto0meingFmrEjZKDY/1obdy/dCl2FntShoxWQ5m26YW8vjHYM22g/1ewMzfjdnyfi9XI2
ZEUBI7egFYbIY+fiM4BbaWnGH1yp5f3CciEpIioNK4VDt5Ok+/O5JezIBZ3Krk+mrZYLuy+1+yNN
Dhtyjg1gKK6FFhqhjKKHRJJkSVx8ezbM+9sHFdRh2wDZQB6qCiLQ1YCWf7+sklnpHIg4ZwJaR1KS
vuskIqGOa1bPDYRRy+MVIXgru/lKZ6Fm1wL7dLlcKk65XAz6h6jALmZhU5vWFJdrjOQeQ5zL+3Av
Zo9CBauOI4tC+2KOPZMTpYkHOwFNQmxjg4eUjjqk3xdqXGeQZiguf/mKO94u+qb+nk3xj0Uie+9/
zfU4dfwssKmrAtM2fvm6V3EbGQ36sIBxcCpW3DuMoA+q2DiFv6rdmU0wc3ZeuIcUpRRZAKZtJZaq
PmypqQ4Bxe5PWrAswBeTINAnP5DA6WPQkApKSvSz+6Eh8yxsQEUc0vq73iJwgGAw7ClHhRH+RG19
GVUE3X54N95MdvFN+UcXFX1yC5BLd4Ad2fRdfhQ3e9ChH5y5bAIObnjVKnTpZu+DIFLkVCdxXrOo
by7VMWPrnVWa/+lR7nUUP1vz+fKrOf7bsmzw/DiFTCvK/tn27jjQKc4vNRdVO/mOLNdztUz6MarC
DViU9vcB2GLb9DPb+qeIXz/RXxau62txns8A5ihwV9pCmQGD52sjUhP9faUL0QfWDb/iVWAJgOkM
hadd5PbYFOMrzP6RnMkG7FiPSNbgPTf1++FBms91ySKRCFkXO3mPtixLVF96ixLNxaTDFjtwPcJq
6cbZUSZHSZw2AO3JpImoODfQVoZ+VlSd9iBE61W4AgefeP0QZcT5AXrkuW6NTZRoEh6TcjV+KAO4
x0XVs0z+jtCM8GStLoLhi1kGOHYHBZq0f5ecSV9VBvWLZ0IewCR/g9dCENNOdq/kn4inbEQD8V3L
kBdcqgJHJAmn4be+R8XOuuWsEXYHEF8wtRMa1GtsUyG0fTgmLVvBQ6/n/lWAlipKx4wr0v6sOeOU
5KxJOeW3X3O6cILluJOLpLD6bh9N6X+jhtsMMCM43cVjeLyVSq67F7eaoBjz3bTSxreHdyj43CQJ
TCV2TjgGCHRwwHpCL5ZfH61tcW7gq1s4QikXbMH9C+f9cstNiOVJAEhFP2Wvmr0A1I+FIcWhDSiq
Of9eg+Y709zPv4AaG0XznJfdVUu0beSBnVziJbq1RDfALhPW/SAisnMKgBlPl3GY+oqR+LFolkU9
JqzZffeNANCyHsEMnponzdiMej6KyuycxnjyP0PubhGb7yH4nGl0y9+5EXmAenTYygYWVcXWsoMC
1HbSrC3ybsKCZoSViSiQdqaoJfX6ILY1579sTS/KHDxI6LzlwDykaMWEZTSCwdj1HCpzHW3ZBZDI
McjaHu71HqYFHGC44NdAz6gBYzmQU2AQVu2YJPtjIIIzmLAAUx9sXHyFwe9MxfEeLV8e4T/ok+76
OqOl6CGUL/e1kGrctyXe6cuYc5ZMtp2zQMxG3MaWwJjn6WTEnKAfSnpo5MATZzq9U94y4+6Rm68Q
ztpFbnrZbeiA1GwsRJ/NxPbYfPa3KCWo3Xxc6TWz1Lv/rHka0HQyI7P9hUI6+YY1jdpE2oVoTK64
kzZ3TKmvxfTu5sAhERSAbKrLGvbGEh+OuKXUKjvrV0obPEI1Dhk8IqUMzQ1Q2pjY//Lg+yomNRcr
9pdH5XJLtUwpEjxTCK6k3F1CeWqTT8XHBmLUVbrHcov4lrHVnMR/jh9PBWUvCi4D5tZdVCGfnTMm
v/a+7EFwpJLHt71BzUx9Aag0fNfaFE7r8ey4c30B0evWeIShps8p2xLZQz7wyPSVMPv0U221AjuL
cr8wXATSkawk3E1Jp/+6bRT3rlPLYMHd2WBJIc3A9p+yqrPLCG9gxqxHcapI1ztFP3g4iAqR/RVu
OQQcJE54IvyfJArJyAw3rbXCZ2XPjH+drbk9ZAnqpxm1dT4WLPe4KVWEyMro/Revvt8+lBvoZz7d
cazrQxkWYnjJrbdXVlPTif/RpRHf9flqOubi+KfFf+10Jc4+nppfdJQsete9INc+w5ADqGrRrIaI
ecP7/8q/U9hiqzNq+BSuHiFX15ZyjZBexXIeJ58bHaAg9RSev+qsrEmkLVDWnfKoSdaXdtCM7kCq
nYOeKZLVRNtg2+FyvMeBrB1eD2HdVp6Oq2EnfMC+n1e0x26QHJWBV7LmO7g4dC9aNlIckYMnrNPL
S/D5lgIAiqz7pS1j99z7O+wfJHLo2YsLt+HQnywEGCUuU40/lIJeP/+nmiZZKxBx1yNnWcJg+Xlh
nUsyBPcavpxUZuQC3lY0cIw07wN1rJCywOgGemPnhgFWn569lJHUU+o8875h1/qf9MTDZPBSbnMR
6KKBaepmKKsZVsFVuq5oN+Tk8b+Ymi5ziWoIduCRZ4vVZE9UgD8u8/L/Qb6Aiq/hexBEO5CiRY28
sQtcZ5xP2ZzkVVgR+xKiwFGCcc2oVPFdTqrX7VxuckQdugAkTqCTejbWZQMfL/gM0gOOcfZwu3ZE
FDcu5X5bw+kLmSblvkgQXcrKyn3JENKAip+GAOsixQHJElV5HKrDO19fniBzjUlD/j169pcUob+a
FC4/XnuNKOIyodH0IhzVqJYIYEltbwCIpcPhliQbf/ztzgiS6vFipxSAzWfzgHs5PBeHGRaAH9oh
KUPQBnQmbq6VGDpxjPQVF0qBbdi4i/GhBnxBc86TMiuBI9kyMu9aL7ijsNwceSbPlSkR0e307Hd9
kKGk4iOSa3BcoMDPmK25lYkFi+S0TRflRiU0uUameoDv4ndfYC4hzJk71tBLL1Y15qnnRhRxB49G
rDfAxIaeR5nQkbALFDDpPG0QoMg3vBY2b/rJzJTvt92h6jrz9I7Z526Y0P80n7o4WNEIy3taO6G9
kOQ8/6ebP/kcWpy04PDWgaRgupv+VfTD7d8vieANjXBcN5thltQi6ViS9RaYLtfoX5OiZO2EqrAW
L/VObfZ+0C0Md19LY5NeVoz6VYwgoB8dUtmZICIqyP/+XhZ6ClV4PSkQzaB0A45e4wya4SWCPrta
3PkotbL2j2kFiLlqgHQEUeUw4L5zwRV05jLAOOLs0h+yvYGwEmcywjSzZtCASr8gmgwfbZqjd9iI
e+LjdSa9tDwee5tzNdaXucW7+dLIM8WVRSuceHmJoSWT0/bI0yu2XDH9vhNND9cvtB/x9LpvaaBL
GFPXTAB2xzY8ACp9HG4EOZVWsftLPslE9KWG2hJQ5kJ5T9VbPgufjW3Vhz1k7LPjjXHj+zl/YFty
t1rQmO+LwHgE2HLXBPL9E7gCL7BgyYVdj41ctog7lrice86gTo7GQH0x1+fwu0X+qvVagQ9SBlFw
tbEFYmqjh+tXiB+zzXd+6ILaIa9eN5RScXzt5i1N3sBGi5FVvKsxn7j3iO1h7wu0C473Ue5q3fIa
sH3kxiDbJHp4rCJk6T8qNJYPvSHs38H/KpYIgdWpRWkCQw8uAi/OidTtwH4AEtXOkCwAnnxCoOzC
D9BdXRoC63qJwROlcz0xQs+8NPYgBYsWENVnAJtKy1lfOsqNsbhHFnzblvSkQXX9MqBbTDY6HzYK
XVrDEChKuz8c/3weSPbCckSR7R+Fyi+qHI7iiQo+CUiaR4TbF0cK2ND2X/NTS/Cc4Vo4ZVIyW7LW
wy0D0MhsnT2toJSlkuAc2IqkPVsHWp4Ro7BYZaN07dDdrYFz3e60vyyEIGMGOKEE5z73UPS/yKrd
hwXO9QflREgoV+yo49t5hdllklok/ePihi16aTTh6QAEFmMhSeXUexmeoekOD01ks9K+vDJvpYMn
n9tgnfV764VYIljPh/30Yc5bi9127IKhxRTR3jc5m61UIKf4er0ACkrobxcztmcUzYEGwUlPiOIp
aWaAIaTrGfwp8/IPVyv+UvEojQpzNGWp4GyblstwnWBNqPDQHryGoTPB1k9B7k7Y6xdLLmUdvf8z
WLXapyFQZNEn367ra2Go96MbS+ql/bayopAoAWhaRteU5/+gLSxSHqVQFgqwZw1PIGbr3NR186JT
Fw9+Tm5puMtRwC1UDMIOCIxaaPCefeJBKbDle7q2u/9f2g82dF9VjtBqstS33sfVyK13YCnTYQp1
IM0LMjz+LB+YF8ydB/Nuoxr+GQ3ZgAWtZSrQ7xsaTs3l8PG0cxUyivwhJHyzOa1z8s5YEve4P8ry
y+/KyLA0TciqKgdthquQw47QnON2TTQkC6hWwHr//zUhCmPsMhLRqz6GzuorfN8BgZQlr3G2lknS
0dalv1dCYtN8hSXzi/VfsY+7nSU1uAaoobueo4NEf600GHt+iFGfxTWTrLGnbHbrni6X3vAbc1bH
WyIuzHNuGIhcfOnf8UVxh7fnjKlGZl78glJYLMClSITtQDj6nfH4CoTOMbPSwcSO0IYJeOUgzl6X
7DtKNnIZW7VxLklbQaTge0iAPcB6+dvOuo/C8/Z6P/6YIbvMXmLUN4O+O1+pAkV9utRDOWAunU2A
Crw7Pd0ctqFIuJUkQTppMINEvWoMplj6qy3TKT7Z1muFJrKS1XwDWycnzak5D7Nf7zTw6noREmsT
J4vmp5EUAIkYHbq76ssygaaaR6jqEBjhfMUiQXVnrsDoxZuFaw45GiZg22RmIUClMt0RORyD9LgB
P2vCS+M8u6OA6LFZbJIOJZbhGKAl7jl3ivCCuHnPywolA0MGi7DoRnc8gzyAPTkruTnYlIKLA6a2
7FqTQD/j1LCGvu0MdmMUw58nznM1bYyMbvM0Cs8ux2Cpc7/Lw6QZZ6ZJxyaaxUx5nv00zQKiTjtB
gS/N16yNcrVVxRkjqwT4h3i5Vb4o8du0QGBseZy4NTlyjsRvqekH4oNVSN6zEqnqLRx681u3QEWs
mG95CsAZIOT6EyC0IQ1Uu8YZwu+Pl1RKb5jU3lDRGtzUle5xaTj5hb7X4nKDqXIW4KP1A6quaE0b
ha0HP7+CnreK6fWuoaX5NGc4WX5fSUCfdYEknMjgOjUuQTZEZ17SQ/Fvuk9yhgLuiUiWspvGPKRz
ryEeMTeeNDCfnJ6VcMYT2mxsoVHEJnWH0WtTwKXU6YcteX2flC9yAe/EW9w2IXUoXJzL+hJjdkoF
3JQH9XkxrcBBfkuFv/RoCajQEeQWS7Lyj/zdJ+14KzQOn8yEjA4Mgp2hPNAR4qPchm5sFrZ7smEc
Dkk7hDWQc6ZPxob8vtksZsTRNu2gqkKSo9TvwIUan5y0LPid+cSC67KfJ6+ZAEUKzDgrUGK9IGDB
MHPIx+xF2zHx3Wu3AnRzYag/z6pj/ldes8en33zeTCZa7HxZA2KvozfW3jJ+LW6jcWWvYK3lktkE
MMtIPN+SYgtNDMHMUY4PYBMoDAXypGrdgRAzcf4AstmXqatex0T5wWAT3e7IJKKGn/JqB62pufGW
SAeEYQa1ImPFM/X/1xVaJvoT6jis9Os9LK8KkvBmRD9fEQg9uW1VJWRYqsF8iQKzEEwSoO/V8pay
PB6mBQNA7V8BJRFwaOz5B9Jn6lQpc1gMnETITaC8gBd/q3ZS3LNNM68fWcRHeBaTjqWvNR1+L8gU
6YLUALDfQWBHhd/vfGwf5twT5Ukmd2cCXvntUVPH9Ir8Uhm54VU7pxZSTARsjQutC0H0YvDMH5zl
8aIaFA75HFpPj/0ho4gxyySB0VuUtEo2Ectj+YAI1bRvRguhSnNL2zKCj7LeZhrqUYn2j9Opc7Ub
KnQBy1nAje3EJTWA3upbYkWiiKz+ohlbyUuXOY6BCX2zDZIUvleyjkmZpM/HRkN85BCpUreirQhg
/sYGqW68jJAj2wGtQVLp3Ozdk7Zi1OoW4RqYvAyESsHdZfTXKFlpoJiDvL7wYbBfz1iStMKW5Ldu
TvsEY23E7HxJJV6opF8heSo6v78LyHjtCwsIogwKu63JuQLdx9MkSslsLfrlu9qGLtiLKwDyFKiI
7KLZyEXbX9VkE0FJupIUHYO5j4BBOIbQqWiHEH7b0qSlYyjCo2yt4altbEvD2SOdT9dSyeNyP5Ca
qvAtJIqezYFYj7C2TcVCir2t34QYZ9Vzyj9ttXct/aWbMSoiXI1j5zT+PRLAdTSGCznd1JZgTTWt
7TCcJHdaIgyODicD+ZfMQNe+IvUqukUlaYWyKINEQHzur8jLSCKNOqSVev+nXgvSsEChebcStKkF
Ke5G1sVYEJ0xW1S1uKIl6Wuv29lWo8MsOoVMiVFkF6NM2yvYo3SAzF8J4WZ2CkXzfFA8zNdJ884i
Re6ppGz/hvoFKBxljDl+Aq5ebPz4vOXV+VNFWDjhg0xvFxIxCbI9ftqgPbSas7RJu1FNwyB9qO4W
rdk0cAmpIcuMsedggZiJ1C6oHUvUPZrxEmtwHKD6r/f/gerTpSLQY56HOFYW3G7yWr3RUrvkGnVp
d7VC530bf1eIN14TFtLZNKNmOriNW5NRNHRxMqQ+AX99Q8Wy1MWxmaqPTMT50r3CXFF0/oN9qbhR
Pf/1zJU9Q5JD7lNrn5J1n9xuuFVKRac2oPQCL3XU/te4TmpepSh+d+6BvjcZmUKq/uqorV4gL+KU
voCI1g6KNJLIFcaPvNeAghmvJ0/j0gfyZCS+oGVeZ3tl1oh4L2I2rQ6nNg8bvTB5Ujkd7VSfYebH
2ec557vMKIzA2H/RHvvSgUpU3Nto7xKo10GCfyAI2j3Pgbt/mivpe15C15ZQtk7dTXJYuDAXlkdc
0OUdw3d1LILvWpUG/ftCHWvjY3frQpX94NIKCwRjEHJAmJ2CrH2mCMtgWmyMKYQCjzJVhkHNUdC8
hj13pr74B5X84LLHVOwKYCWjCP3Up6dADxRVrZhg9YW29TcyU3FfLjU4w8vMCHidkur1rcDxLtiZ
bW375anD47qKZaNkGQkj5aJAppxZZmSows8o4lDB2MAgHrWnBBvqC+V7cFOQP6wWB8o6Bvcchk7Z
4doQP8/5H8SW2Qse36KBUdGo2/UcYdAP/keknhWlmvCPLiMP9LHZ7R2eFskVJrxF5/7OLBQCdJ4Z
FpQvWIKRyG65CpNizLKH0Sz0Bakf4ILPQ9kB8Q5jp2w9BHO5t7R8AjGYu/XBI0v/Irz33Ao64u7O
6nbAlh6PCTortdMjFeVEInF15t5x++7PzstSyX0H3DZRd9MTbEh1Y8H/ZTs0QIzy1R/iCgKQy1ll
HU55xpy9Hp4lzBywUv37zC0To9Po7gLfyiUYT/IhGCM6RTfmXxmMEJz3x/Do73A/2g2GdAtZ7K0D
fwMBgwLABytPv8rXNpTN4RrsFsWjF710JJC4b8aaGKHW4DD8XnQaaJx88bIpeQBimnWhpFFN0Ceq
1O5rj/oYQ/BLXX+Qsz7GkNnZ3KdViU3DVnsgSEjJtUgtg6dyD1lVfZN7ITSriTfOeHYWhNIJD/TF
3jzRR/nk9/S8BK6HAi+3TADKilqYXbB8m07i5cRNlHvC5J47XH0PnO8hb4be30oVf6FRPy8mTf80
WgPnDsAPFsBPBQJ87jLV0uaeDXrJUOdnyfoACQOkFNNy42xVj6zXpGoiZxSoFXqgQh8HcZ4aHAgh
SS5m1wzvlqBy1gqz3ShJIKtO7aKopj/nn9s4sJ+cCTrHNA3J3WKhQO0WEbdW7RRpxtUTUWceRTDI
zLuh7c3QtB+l378Rgv1YNCDKU7OvAcUgp8s20GTdBcMVKSxp1V7vVdLwY9mPocp6Q+TnzkYMsTlh
igndxy2+CJr5mzAkEzHkKY9KKOR4UxaeU06m6Nexai1vgNb0Yie4wA7X/Jn0HTpgnM6BzbDVAz8K
52ikkK1gSvxhD8CIWLAZ7ZpuOqX+JLLQps8LG2djyDz6bN9z5ZgrPMk9uL96FNV0mnsmnrhxO1vq
+3kt2kWFcl2XW3AaKqbfJ7qoSkqUFdw8q2rD9mlyioD9jXnGY12zsRNvW2RZhW351pkU64FzTSeP
xXE9iG/KfWcFTFmWF/Mgfb2gBnwlaS3G2V/+YXT7Cnj2G3wx46K/66wPbzFsIYTCAKKGqYU28jPQ
HAOfaY4UPaBTMoJitYwFH1YkbS1/S/wq7OQntnROfj+gUkdR/JzJDA8vjb5fSFsaKPbGqO9sgJNI
FbXSngYKuCRSp7OD4Rh7YqqRBngG0WcAMe/IR94DxH4upFs5VavcU2pBvjiiLyjy6cJ9mrT8/+Rj
w8290blap1tWhEuECdDD8zkN7oMRWvhHL20pCqQQHyLHPvEx+H9Y8CKtsXCmrCiGxJlUXBK/SrEp
BQSoboq/aUAlmLGGZckrsDDWEo4cicCHohfFLUjTykK0MmxYlMZfi2sDWfIN/Y8/VI9RnHo0A3R1
QoF2Kt946RarH24d/2f4SRhpAE6hWqkp3ZpnEtHwAZx/N+pbUIRDEzXNf9DEl/o9eVifE3XrJVXC
RmZiRhWFU9L8qxZBUGgZapRVifR00eunqk1aQT6BzxDGjdF6HlQD5PqbOF4Wa3DeEBhCTnhjeJBO
Lz+GOWD581klEE8Rxn9Rjpp7Sa90J61154TArvLmldc/IjNSpsAfV5UPVQX+znXwCiRzm82AaEIf
uNU4iKoh7rLMAmtcQHfeVgfdTlXKP8OUE2on2m2Hty5DFNHhZO17w+S+ThNDaI53SBTcI7ir/myp
k/hQCColbLVt6PxOjuSW4OyjrOwg1g3c7W0Vrfqg8ptbaDZQMrh/kia2d8IApBErtvwz8SoTyV2o
SlyjX3XPCByCtlHg0DvZGY3dFyymAFozr+E+xdS5Edv7rr+df3HL5alrKebbKsmLbCBiiMneHY+A
uPYFyGxlTawZY3jpbC6dgPipEOG72XXGTY1FLYiOj9ZmKMDb9MeCy9GERy4yi08CaNi66IRXbQGv
FbnMzp2m975GX693BDz5zUbUAeYayV1vvifriOiyB5ZZMtX5D8ky7CHrN66ddzS6Xqwjwujy9Lf+
zQSoaRHM/wvtTtNPPOdzeIZqQ5dWwTzPyQZ9huVm5jLQSh4jFPoiC3RRKHpIS5BZjuOZnmyfD2pz
6Z/3i2tXDaFTbyuMTkzTtvQDhBSWlvOdbV7J1Sb2lEpJqh5kUxCwfV3U5n5UvDUgH0Bwym30qoQq
/vAVg4lBpulIuti9scZeY6SZbzFozIgEYb2JNC2odVyQt2wMv//ogUS3kkzuJ8erM8XGc1RkpjlB
0HllMlmBUc+1KAp9KbJSweBTA+9pily6TfER//qz/1pt0q+L52H0QRHE191uasqYhSWwfrLcsrDl
dZhY2LW7HIpEfP02HbzXVoq8zuCqD7zscgRL1IBx5jn7xT3JleYYMrrWcPl9CP6S9HDcbmmcZ57X
EiTCIUMrEnCm49GTuiBVxQEPONlgbgKbi3HqJpYA9Ip/u+ymIy6Sv9vHCpeqFMGXHr29YJOG2MNY
om6nNZlcb1Y7XG9HooMtpH7AwSbK3KmGuBYQ4F6ar/9REqHLK7AXQVuxBTMDgmc/fcpmH0HgNqEk
LEtmUiBKTNgIoy+rD11BQzCNVmBHu6G9JlNvv69L9moACRdPCe2fT4ZOUJcdDKEWs37jzADmrOz0
9fOiOB7lXnS+IyJG7NS4HWF0RFPLMvV1iU3OcMkC9Jx1UCv4sgrs1AKb2OF2sMLXkKS3wkmbocK2
soZT6PGrX3AYxUqE2MCZcMeyIrvqpE2OhfkR+ixWOB/fPwdJVFZBHULfomrxw1nUjsgotyFDPyrp
kW0oMlf9W98TahV7zXQdAU2lkoFSasx1RIFAbl7iXWPgVv632kJR5LqKspnHiCgkOGhK7huNOLl+
bjnWdVKxxefKioi2IwsJdFvU2jVSsK0OWiqOLmi5XfSThmJMK4ejF1tl+SKeyKbqRk1T1RWO64o2
X4hLZx/a5/de7oGnIDFfpTX2r5RGtn4iky3868TEU+TLH6bm0Yio0eXTmRr3rgBwKjNHh5usKUIG
FQ9/BiEId8oLp52LwwNBwvhDW1brxiI8/2II/V0MOlF5TM5MJ3XrB5wFgTSEM9xsYnAOriTdemCS
i9RKRzFmq3wTxOwBOTZznkDZwhu9Hug1FGqgo29k90gTVnLKlFb/NldZw24EJJ6xoqIawxBXE7/G
Ll6UNZRGA7LqD9yXGI+d5BUBz1G34dBfjvVwDY/w6HmE1LqAT68bRaKJ3CZf0PylsURlQ6diyCvD
ok9PoYabzxfXsZE6U1mAwzCK3akeeIzSnXoXg+pIwXd/VKMUivm8RSQ0RMlut5YN0jJGFx1YKv8y
veHpVRqaFM/S/UDZTTBOPq4cqG8wsaHQnkJ/mFrYBG9Oy9nOfN9LXDksXq5clPdGDziLwkBUbehO
EbIAfGVJ3MSbDbgCZ3YIyS/EwvVJb81SzEHV7LwMeTcVaJePgxefz0ZUFnt52IbQzN4zIS/w7jjB
RrQdX3vpgifRUrVpdFMm4N4mmnPgBWHmvBHJi8vUx7DMZd7+V1h5tSxbaDDdlyilxFNOwFwLdH8T
hLA7lGEhjoUIP4IDarMxGs6xmL17cy/QOJnRaZTu9atXTIEvnOokU2spsiDPjyC9hEz19RQxpXYh
djqpSmBAEEeLL0N+ST3svVhB8ZveH4Hni7bX7dV81PrKSOZaP1RMyoVBW4/RJaScNtdXbWajoSBx
nLR8DASNN6ojblASP6lsQflWFit04x1bVT5BA6TXTBm7FEmb+hOrLyVQTH+AVD/wAhVTuttj7SDw
zs7Fu7xkSnWECeEnE+AILW8dDN6nZrvAh23l/5vnXJ4wc/vy5UtrgEz+26GOG75aEJj1HCUCPPUL
NesQHskT+A1nYP82roYsRYVQRTu3N4ddIuPdYvpXBOu1A207tsPigu4XdjOdQfBFvx2ejKjIh9v1
aS3jXShb1/LWo7RdDEk9YhHFCVs59gNma1rTJeXRtgL5C83PbPln37xoWlGbbTvqiGgha5JisCW3
O26ffEVMdO0n0uHyfmMAfAcC3CEyWJpYl+6Xnt1ObflyM2n2BISPAMoK/uHMlCJGP8a3erBDXyLO
WoWmvH52nmGbVFM8CxlKOdbuf9gr2aPDuFf7dUh6a6rZNxaYrtJEImj7hnLRNQj5RaCKbR2l3MGC
rkCDQ2s2fGtHpFuLEmB+V2mrTHFP9mSX6iLLrEyIIkEvF98hlJTetEnavfnRXna6sxajPeTGdsXs
IczMC23N0sM+SYCOWxv4PJDVuuSFcHIE/3j0ar8DwdK1/mtK9yN5Dd8j6jpO5JDqDx4RLFpIdCJ6
8aqyZKx7VOB1okTtgExIIwHiPubf1bnIo126Rq0toSaJstT2bha4UBYflW+s/e92xdkGNOliWHVa
j0tdPD25yuPIk1kawPxCWO6p3JsBvYIarSYMNIf3UHEgFki5WfCBNLenwMkJeQOyuFYzYHpiGNEA
kWiVjSwvddNYePqJDqhMEIpge9zYJoN95gumdG3RFeCun+jhXViFoyyE3MgjZnzZTS0EWgHb7aIA
VwPBr5yZgdWPsu4uzQBP8i3GU8bPtuOgPSkVcy/eYPe230XzWDtMB7CxAZDImbAi6orzQgb4FpNp
AL/e7E3jcvtXt8JFmMsoBLovjTNYNlJHG4yfe3hSK6b5vxoQzLIAVuSsoeknkmUMq7Ie02pClpLb
YbWElek5utbS2xE6weXexZ0lZ86TAKdgngMbJ9iu/L213b6yVmg3Gz+m9ShRiitnTVLN05Qew8yL
d3vo/W73I5I0mGBGFiHlCTquF0t8tX/WS3y5bLWVKuzGhwFD75WU/RZRQQMqtGxQilxkKIxWLIrX
f0Sf3TQs2IqhjbNCShT/RRrG93gd/NOAD0sKLyFMqsk6rqbHmg0JrLOGbKWVHeVD7Ur/3HFMKGiE
0nmFgw2SVwyhhn0TBtvl4ylZ2Jg72oNmDLP3mU2x5nlj2QjIDvNsDT5Q8gf9v5SvGQq8BhCMUVB+
LGp34bd+D5SBTwfm4Yd3uJk1EQ7LkCFnVgmhqKo2Ne6sJRAF1WrKVaLy4Fv18djcakYjyE4ODhIy
csQJnVneOVSyQMgP76j3q8Z2Wg2ojQf2Pd+pTlFKf0emlmj/wZsWm1vBOidpY258w1SxZO1Nq/vc
TZyGXjcme650MDKU/DCv0eRdWZOlaS16t0MJ9ykeuE/B4mXvFPY6A+p4lrzb4doA0Oj1CVX8FKkw
s2deyUBu2y70YMG+9fsWaobfMiD8JtZ/7RSHrQen734yfR/xIfyKmNp4mGktW2Dm43MDpdQuiM02
rMXHQ5/OJY4hwx1HcGe/Un8LQ/g/XPSU3LxKkz7urgxqisWY3FV5S4I09amdbO5e/RQbqBAZpXcR
0/gn6xMJbanDeW0SKliwjbyhKIh3hlX8PMhe7nbX48rWYJ7N7ZQzN/rtCud2FE2rZTQYofg7w1vm
ZhF/dXQFGoLWfJWW3mLbaUqpCezSDTU2l2OjeTm62Jt/k7rTdS2yx+6U6JV0Nv57VRwk8N8OJieI
jTPEdsIkvZ0Hi3NMQW92tOREoXjU3sqtzkycet/JrcgmW05cBsRLks5S+W9uY+OPV5145MA0RQbi
CAsWRufiIxcZTD11H59tx6XU3uX3c7LftEOpk1yKqldCLhOG0erUzIP+pvhyPYtf3es4FFjTT7tt
8B2dM5exulvIUWO+NehyRvlTBpFRnCN4xFW1xnBJdStwfj5MY9q1b70gw7PmYseey3db1YQWKDju
fUOxHBYP4+BlGhYGzAOzyZ+y0hVp8KxT97Vqr74A97STyKhoRxUqRAMLzCpoEKX39JiYswJjYBAq
yT9UnaztqFCTYfLseihmcma1wL/euQ6PzEGItcLhtUSQIU6S5nOjYHkCnF9nx7xo4FqSabAuHEwU
dOnwcJ7sRqZj+TlhJNGPDEZv6a/wBaqf4l4OhFv/HvGubYMmoy6G2l1h8B+5QY1uYJcwAeZk82aR
kUAfH8/gtzaSXYdSt94r473boLGGH+z78u7Y6+q8kVBhSosSlM2EYCtEPvLRhg5We2QEjJxCr976
8H0UGAa+uoEMqZI9U2hy2i/sVAz4M6jD2M3Gdh2D4FTPBVkrHEy+gdmooVIn/tw9Qi7a1QCpP9n9
9aIvUNIrnrFVes8rxIlAQdKhVIJXLf1e7Y2Ca8QWdmAgKwcHCL3mwmIKyfXHVXgR6yJCoXfL27R2
7UPoqHju9l3EMreFt4aXS7G7aMqjRVFq4zuSeHMx+ZJWM5SwO8FhXPXELqGpQzl5AiUG9dkwt9N5
BDac1junkrhuRtL90x/iUuax3ws0elWrf8dHVigTOR4Mu6dOOJQ0LyIdwTivaE9tKW2aopj4uNiN
HPjDUYFN/qFq3y1HetVCNKRvXTTZbiUyuAKPPlfNvcgGSyOFr5jrjJUuNIGWmsj+KLEjtrLmWDgY
JmJaTdTqNm/CMVtxIOfHrH/pglfkPweDCh+p80vHDRcsG14n7I5dJxb5wR3jLTFpN/bfNG53ZgNt
DfypHnblJ1RXEHkLMi5rhcvsSzhDX28aK5ypHoYoy5bJb/mYkBm6ZNb+FDruGQegxECgJ1UcdFwl
/agTLCl3g4e3P+rDKAdP3aIcfnI8aeh6Z7OWLHkoxv5K/GFAUji4sNAvcf4o/UcDFrfaKK9O4HBe
KTigQQnOf5ccVa5ko5+GPGVA0hitXYoyNmkaUeVcAzk5725rQrXvinb3n6HgOoNYRno6NBLdUNk1
kLeUAUtd4Hv3q7rVeoDBQyR+SiftocJgD25MkFKSkwg/NtLkAabz6w9cE9ss5xM/dpumeb9TYiia
qEWuaVdy5C1e039FEv4xN1K0SoxU/I9DZIZaqLsUITEmGZQUoPVa5zwG42ud/J6n7sFDqyLeAgcI
9J8+E1yBcjDzyaoH5qgqn4MOolx9ytEV6+rSeRFAZ3Y4a8W7IXYT+HKQkwVriJxj00ULD4NY3PxK
qMTZj+RUylQQ5GA1DKsmPRFmztOEIf/TuTHWRlOLS1hsxir5+6sbl4xwTrILC+CzXqGfJVvkN7Dl
gUhX74TtkNwPb6BQUdO9vxZCb0soztTIUFs8DbVG+dDx228RAp5iJa3cJJmwrZ4JpK11JpYq8Y4E
RD0PXxBnCUQNCZjh33Wz3+dtvBkYzPth5QdnllyaQwF+uP6Pzp1MgSV4gqFmoLVdujguo/FICXLB
5ayKyAZoYOon/FNrtgtUWabcOuW6OdZW3p447oKRWnuBBAWkMKTb8lokQRqUCXur2Iv3PUDshuZR
D94UzLxOa+pJz0+gOrTP5KOVHnthMmZDfOQ/eGaFw3nHQybroKHy/HFv4rbO5N9iHztgvbm0tLf1
MVVXmeSGKlS3ifzEIFtPtVVymDwikQXBVpynyV7rVgBFjuvX34C0cP1RD8Q74imVZ05mpBzViicp
W9LKeUIXC4YUZbVSIUzERhkXyo9O5SOudUAubdvPc+5n3FoJQCiCrxB5S2M7PuVTmIyJzLskvhaP
uNMvlJnxw1MbvByrW7wWbu+ZBhBB4Rm1AqN5aTkLfq5smBA/qljWRlPuKy+B9n6CPjLaQJ4faGsf
Yd1yfHPRz/W51jUwzb9qai9GANmdicFsxMdGIm0zQGiSjYzCoMskGh1t/JEb2rluNm8jnhHMP5qt
KjI1oGZPVsI8FIbpJhZX2KebTumgrD8fP179CI6NUkZHbYuR2VqWeU6pGT/Sk6RitXJQqRx38Tg4
6VD14CgmBoiCbYqtxEMbsrr0yhg0JdD1tY99zgvI7h2Rt5ICv+4nr0DTZj8GEEAQnMBzWvHtIhxR
WzKZuwo0SGKhAtBdj9fc27qjeSUNrJwRZUsoftx/afn2fOLU77yNXWW1v1Gp6VYTCRX0xPQB8y7A
XM9Roe4x+IkxLU4PAabV0ORe0c1TEok/VpwviSE1L3XIx+J8mpsmG1mNpyHCubACla7cv/4AXLpV
h/Nt5fely2wacNmG3nOQ/NfNyKW6BB1JArvapAxaZJ2sEDo3Ca3Zbz1Mfm81++5C8kth06H0aCzj
hMOObA1rAPBK1CS8MBK3WDc1UUldHuvAc8/+vZq9lxEAYWiQAVvbCR5WsS/O9USWbymiwIuQBbCU
ZW+U+wnv6J4qJtSq7XBaVhXCktjkvnYFc6Av5xFLnaUaaohC1oalqHZbOL+VRpaD4rb25RUOSJiP
RyAp1q3uXrm7nzeFI1PjruQhwXu/3UR7EoPq9SY0PMccTZ7sNVSon4l/0BZOj+5DgYbqeRpegY5k
zL9UvEqn5xW3brew9WVeUK3XtaZA9LFUwPBSMIufGj/90mzra9t7wTBwOYznRZIJGX1BunQE6ept
N0PSuKl/xWW858Nt93JAwe4Tlww7FsPPa0yaCRkIFvQ24Fibk+O4FgssikMhBBOt+23GqBcwk+/h
5ir3rfl4MuHVyXfUNa+HCHVvEKTL7t7gjpzOKm0E1fj7svdXWTni1rfkg6fZ6wgTp/cO5lU0bOyr
ZRPDMA5LxKNkQggseC+5dytwAQhFDZBVZQj13jMekJL4vpozAh/N4FxfOXGfl4wWm9vTGgPevNag
iDiY/qTEVT5MCU3ESl2chwLoD/DL4xeu1RGJ/pwHNg65uoJVhuY2yD0tVwqCnRYhdsvNNZug984o
cJbAhZIssefzRfNVxIisAH0X1VHUtZJDE81ialfSlAGiYs3IuJHSimd3vftcKoEGUqOXX+5gR7Nd
XZJWKqzI/p1vduFOU2phsdXLMG2uaVdf56FPjLXssTjp64im/lCIuwDMsTAb4wpA5YKD5S1Tcyai
81xXAfwdH2ohav8JSshKw4VwO0M3Nqn54AH+nDOB37E3jHgVEmf2wBLqFqNWFJ0RjKjnaTVPwv06
RyVY30fpumChs1mVsh5urGQKZbf8YXznA0zVBZHWz7LN8QhRkLVMHCE4ULwxrU4aYdkQz+Qr9wyo
kOuDSNzXFUlCsGDDIhZ6fgyS5zHXGfp99m+qhkqoNNs4K2HJTv4hg6zGUyY1z0uR4DeZ2FEw7ODf
+aVYoZWZGlVsCrpOfTXFPQ8mOSQgLkSffvaxSMnswe6RfW1q8Nt+5fbf5e/CWq8/pQFDt/XXGhkM
lo9pYYPvNieUwLjUo5d5Jfa13NuP1a62yDSE5uURxQspwsOxfdXGBbrAf97vozvpwhOmhGRnENsM
DsWJt/cBQQiY78Xf36cEjzm7RWNoynWLKhLEHDNp8hj0QvWr9YSCHymgSdgl+CIFxnqOApbAnmAl
007/FElSX64h0sq7DGdbnlFuZWOGt4QW068F1ZJ9LWsRpVhonTzfeQwUYd81BdDG2BGORPe/r2Ey
jprJryVSk7yjHiBXzkLNCgf7efQmg7Ob2YXcKUbJwhpqlDxHaTfzcmbuV192eHJ3mbSWYhz6UYaj
App+ciAOefO/LxrPht4G5OkL7NA2hTcHAGAHkK4roO1UTSRW3RS4y0P0RgJonjUQ/3eNipCI82PD
bRrK0/UywiDiv7EOfPVgyOGtkXrTxDaABVTKI5hR5ZGTx81SOKpdXJ3YolWqThk3u+oiNaz64a85
pUXIYMz2/BGobtvgClKxs5iuh995zn3hT6UUoZpQ3a7/p2tMdy7sqaJVZDPkWLXcMonvn8gEpmj7
u/40CRJH0PNQ92Esb38ciX+x/ocbMgHmJWXjWR9W93KqsCzahmujORtofDPeZFBIabCXYpqP5TlN
hLGWRLrB4huleIfTo53D9zHCSIDM/QK6YuyyiQTXRwCmwP6dRHG8w84jeix7orRK7BzIqygr6fDX
rz7i5JCD2r7T5R4MLQOfGGNwcKGIMH/mbciye+lQ16LmQztrgS7JtywGhzDog2ZKKBd8mKQ51IYJ
Xr8SXfSHC78eY9qUxvP3InNrtYfA9NvmuUhFaHseqkPIm1ly3CAHlkELXGRMu6E+Lxs3RjbkQ7wb
mF8kjsk4m/SZMOFIiTK/BWZt2PIvHyBTccZCHq7W3CnX75nDYTkPwZ4IZqGY4wtMcEMm8SCVHYSW
NUqOf6ruUMYfohSB3QNqiBMm1Ivm/zAU+VwXnOYw6yUVe+1FB6WTHpKTr+wBHaj7AbQmt2aKzgoj
3pq4EDGLGF2Sz55B8Jmi0ZNm2O7SxaqpiaILjiJGgDZTeWH7nU5BnmMEyN+JrmqEKX/GLq9W10br
jHAFg8u9xdibBTnGY3xhlQBwWQH0pKgcIKTdf+eniOgLRoCm0UojGMPvY9eeiOqB+rgjxZTSqn7X
AoGZvdM/MyvY75/WyvinvWD6NMVjXFecxVBzniVm3Brj/nWagvUvzD7hpMcRKRGP4Q37pXt+p4j/
k+tLaXoY/hAkhEWkEljc9lnRq00EzPCLMNG8pqxoQhyrTDgbXqolJCigGv3MTKRGh/1sPePse+tz
POUCthFggZmtBQTwczdAbebHLHbgjQ3jBBwz6NwGXhvenPa5+c3p6HJ7f4vXCIvrj5wbsru//GSS
P5By7EODqAOz2TCkbJGke8TWCH8vax+D0UzImbI6/SDJtr5wuiLXtk0R2c4NgD+6x3+O+ahHpmGf
UkLkwZ4Gb3prQKIDWsMy3rd2hMt8qTaioCFxeuzb591M4J7bmFr6e5oXwQSF91QXM68KTQ/66UGD
bT3zvlaqLtt81rhOJpWcTfvfLuFWlOqiQLPYepB8yJ+RlkjhpTT4szuMonYli95dlXUoKMnjF+o4
K2jKMJUkLuyxLWG21UCZjnMfTXtDQPraMU41fiBT1xMOjtLs7yJ47LhH8nNUfvmzfqSU+f838Hbn
JHRRSaEeJiec4V/OW80rL5IfUkjHEF5ijyZW/QiM3AxLwld1HuV3V8lVXY0jDDPrBC0XYXCQZ4e2
IbAA8ebOUjhhwGwmtqWC7hZhAR3nT2tQ8CldmxTRP78Xf8rVJtda+1RIh7g3SOXBuKIfOzVxSTeD
cNRJwci1zfjfvQZkV35Gqlyn34U0OsQjkq5jalJFLxtCDDUqICa3TBJNLPKPLYUfmFpJyF0oqta1
8kYQN6OFUngS5jn4TMhyWUW6lAk4uLyObZ4WHOXsUd/8DCaVdHqYesMAPFqSkyYfIq61AlcSAX/0
wRD2N0TLBV7vzqRUqz3nWhtVazD1vvL7aSHARDDWZli69IjBUax8Hiva3vultyhm0WMI7By7wmDt
yYc3Xj0MCvjXY0x13A8ap5rKD1IfQacvGinBFIhYheRWp3bSV1t0FzSOolFLFAtTJmWO3So5pWSw
N8ZqxTxh7hM/I4hbNX3/W8eNW/SVWfzt2xTGuVqQYwXUbm5OtH8g7+VWI7SrPSK++/znLh0u3EUj
Ax2HyrIWGzMmcAHPLOa9SUcldtnWiph+vYbzuZrRG+jK3P7D2k7UMWl0KgBuA007MC4fk/ylbMEa
jR2V3VwIJnxEyBGWTSBwJ2aqERqNViS3ftdLDhOfummxCDzAozEr3uX1FJr3ETTghzVQZsO9oHMD
Vub8vY+EyXYdhK2y/sGaFETwA+5AajIlr14k/OGhlroYzf1QtlCrWeYkUQadPYRroyR0yHQ2RbQ3
i9dzse+qyiLmkmHaWAu0ajpRzmEczoRX7wEoVJKE2c7yPajYAARbJiYlKGg9sP2MB/+tavGvikEY
WE3eqAz49ZrCopCYBgcv8YlgToCDD+aykv/Iqk11SMOxa9uxAI/DDqDdUvN/w2czcTyRL9dZ+v31
IXdLNDwiyI3etjI9MLCFg737IF9n35Rmr5Lm8SoEC4t6Kb55bEPpL/zAPLh8GNJUAwS0LJKqNKRl
2LneiRMdEMJE2llu8BJKIGRl8zGxgNUAjVKCRXEbaN73siK0bzJw41eag8g6BVwoSWmdvu/vhz1R
4KciZ361KI/u3Q4XiJyADokq60u0xkdWItVQ5ymUbF4trYxRq8C/jIEjcz5cCNB4wKTO1m0KRoU4
bFhfo+ynMBgUlMzcZhHqtXDkd0oMltEWZM/8NV5n4G7svUzby0566SFTlfX4lw6T3qZAwtrlZdPc
gILP7uM+SCYT1vWzEU9dccSW/0cWrOLH2BBXKeDIoXGg+Lfh3YlFRgglt5fxbW/WV4DvyqKYMYCG
oXRjaAyr4k4JAmTLgvympzknXwhDFQtGfvUBWw/Gk3LVNJcAEtk+GE/m0VSAlQ1fs45435fEByk8
vqQjDQWr92zjbVSJ5AL/5MMgARb+23hnwucP1KR/+d8v1WyXQr0umLdRVbOflczFyTSX161JmQPH
oP7A0nnTfy2D3K9YieD6n2ZCGwuFyoCjnm5E4/TDey57yDeKKdfTAJaaBdUb8WbsNEeDfJSDs2cy
jBXX3Loh/9ETaXgrrIT+0THJ8aibr7JR8reh0sSkVbbJeomSTKHwqacSzsKaUazsrF4fccb6+2hG
3KGTj0eBbO0vlH75A7ipBd9Rv/PIdwiLe3YyNq1Or4l6hrCXJFkqzBoUBD1sHoSd0TQBwSDFvqWM
sZD0ZlgnfnSBGP2o8Y3UvaU5AfhACQl6l43jlAwmq5qUL2AKctUYKDw1DACY5/DBWQ1W5gkhMZQ2
9yCqcpYadWUZ2Q7h46sI1Eto9Zqt9qAYrcza0nj0n4V1A/h149WAbNPukoebdMXwQz5RyrLEiE3x
riNMQPSQ8pb6MecvT3CIKFyFCCBPs/+wIkno5TzMrq6VZGA7rs5C5ncbRQPi+gMwsaN3TRkwcdIm
CIU7glNDbSZWt5/sHY+0AeKCivt7JWZYDhcAznuYHcgpwzoFkGsT+VWzZD9x2rfJprrx3K7JyMlw
eCaKq/pdUDBrBTe1S4G8/Rh9vlPl3zX3xqWS6pXXuE6p6MINBQyzf6Xu7zW7/WNuR7bEZt0YmcPO
SMMyA7gEXcGA/NYS8plcFj8nNkFVneNelFiUNbzGM/Mf78o2nksKHZGgqV/0BjkfjweK0UHE1nAg
2l+TEFcXy6IHYL6eq2F/GF8FZhI8D04fPTFWWVnJI/BYh+QrW7rUQEMKPnZmWMGsAObrPrBkwzhY
Hiu/gDakc7DoGhuab02oiiYqsjp41DFKECMzTIxeQuPmpJf9mM1sd6xr+kzTH3gWhVFt3qki7ng0
+ZMCQ3aKdA4N901LSItsfMzcFfEAydb/2SoPJ2KVBDa4l2xCabd0wHCNia+Hzo1RyHi6yeP44GLP
Xky1d38oVvpzOseO3Hldpwv0PoLw/qYCK78DZnK72v5+knzdZnvGpGIx4tqzvGBkns1/JOFfP3yL
P5Jb4O53zUR2TAX+4JB6Tf2PoYD1Hdi3sAcCoB8VsoPURL1CTnwgiMev1ZcagtmQ3L5Yt14YUdaA
zRkVKWAzDvSA2Q17rnpdPh2IiGHC2WgYVtaJIlSjs2DgVVQybIPlQWEQ/yFq4YT0kv21WL6gHOjL
mvE5Brl6XLp9JOXb0nkpQyHmj/zQdQQoUVeJfCZpDt1FKVslnC/84Taz8Bm0WnHVMT+wlSjB6O0j
ewL18FzzNUW5cBF++U5bJ0jwsTgPGLdg9bZEc38/8cBAJ8lyPXBGUScahGz3VwOLapxvLT1cxMHB
C06wcyzmKieAUd7AZPBmcsEtXrIACVXOirSBkwRL0nj6VD8vBHh961Vga1h9ME7JholsM+o9aLLc
FUscwJMAGH/WhHWUIQVFZqlOhoVwMrZaEG9EC4dEtafu0CYa33GDpSJnABeegcWODSOoe11+WrLd
zni71NIv+6lck5lH2FM7R6w7IHGuz/bT+bhY6505E06L+oukrdxfYuSu3Jn1gxRKok9ZyjqhpQJI
p1IocsB2cNG/dHpRpw0Uv01DwvQ4I3l4/lw+4ApEQOsb2IHimEvFLnlNDY5GZdZJ6ng+7r+A0lNP
XYV+0MCIshyQfhWqZCkCUzAnjzTyc9GrE/vD8IcuUHkIiok00e3BAbVPOMrOyfCvBYbNfe1wfoxI
+aQZ3j9l1ExjHywXMyjgJJqu3aUmiHDuOVNsFNN8YSqvwRljCfNsrDCn/qwCxGCWDRFmSQXPJjZF
wt/pm141qNR0Mix9HFuMGdIcvIZQx/HpHrMvcrX2nNygt8UCJ/hMLvimvqNn8oRhhOFKsmQa53vn
uh0nY/H5sEPtzR6tMn4FxcrBMz+51UUybJ97LMVFwDs7mYDmfgpHLimPvZttK2IR3M15ik3zSnCp
CtJZzPVxSnvzjbHsJXOv3CRj6/0Dmw4J+jKkZeH1JbnbmjEIF40/WZkB9LvyXJE1aVWontQTpDuS
ms0tVb+J7CNu8tg9IN3BHB4jedB5vA8myq6ZQlVQbcDCv/K/lbJ80fcqelvnwfTlgcvQul6lVwtk
720Fe+fTrA9itZ0a2mgAVzX/o2AYvw2Wpy8BqeDLYzb4zFU7PSLHS/CRFM31ybaHvdnKMjsjHth2
Dt02FyhNYTN5U08EoiotdvKJdVklmnCFN7iwC4n4QKyYc1IxZS+q6APZxhxClHKFw3233R2s4DSz
2ImY++HUTksEBNSZJtx/ntInIcoNABoXM3zx5cg2nBzIHzEKmlSIGki6eTrPwlymTRZZRIHETb6P
bW8VnFOmLkULnVxKfKWFVPqgA/JsJ0sxh+s9tl47NfIFyuEjVyBb+R36idoQhrIXVJb1K/fKU6Ra
meeM0RTFebkE+fF1t/AQKHz7YiuK2lcaJi6X1eh+yEjv3NTrngN1EAfAoh28puT3u5AI8QTZG+WC
SNkXSd8G6yfy1idY+U7seIJGHSIJLanQxnz2O6eSILYGYWo3InExLGmep7OUoFFIYS/5hatd3FbM
5Z7LsDftu3mHx+asVoU7xRKNiRqzNlt9WWUYl8FkIdPOXboM9mpiqrJoSxf3Gu+eEJQgQcDEtxLt
/Fx+JSkOyq3G2BVBJRD9bNJoQXs4k2j+6IgOfzyL3ekpE5rh0/kWKUdtXSgIbXg23TmCCqKQRRdo
s/xLi+JR7GTYIpA5KRdYs7jVflvvLbYsUUALVsLFUzDuDYJcXB4OjMoezOzvZUmaNAFqwqIosYEF
INYaO/Dx/g9Plzqykc9w3HJuxMR4y38dbtAz6YOIZNEuBocBSnaDANnDctKQupDL2gsQqh9Hntm5
lB9Oyg2g545BJ88bTXidY+n+5u7y0fw1IbiRUNfiFxD/B0PuczYZYrFsGO479yrmdgzSzMbqgxSa
DZTe+cr5tebbNqFuZ8SJlz2m5v2effX3rsu6LqbUODBO1ieKjUpYr06Zxh7OOqjjVyv7Hl18wyVZ
y9bgvGj/7eqgTq51GTKnRSzlbdr7CaP39eS0ZkL+knYT9lGBBwp+v2P+f8g+PMnuf+eZpN3i3RnY
jAY0ImmL4lfUL1takxIHE+aPQIGaTPszegMB8kSoChZ/3x648bVrgJsUKCUhjawRLk8QQETmJPo4
KyMtgkHJOcPUoCElEO3rWoyk0W96u0/fm0saJ+WnGwlFZm44KKA/1qLTvoqRJMixsF0NW6CZym+F
zufQVZLJVkn2JNHHGpJMMEkCJRRFx2JbuzRnWuhdfUe3XApp8UzSc/75tAehj2COZqJsg75/cgxS
r23BN5IvsaCVkZ6xX5NiaHz+x5GaMN2y9Wxn+Axbby+Uvv8O0byDbxtR/2eW00+MMlWCmOUMr1ui
pjg0NgrwqngRWCUkF6LWgRCO2bAOJHL1cFL7mJ1KTUIkWHnO8MNTH+HwuYal+nkEH5bSLC6nM1PQ
M4j4P5zoPAgocfff4dorK0aDpGlFD4kiZbTgom0V1bFL9FvfOxiKo+eV3OrwdbAxdD1dZE3poLhJ
wurG4xaYeCUPGTK8HeRSvuL3ieSvvsf0ISDIBcpoh0FwZ87NnJ7xcBRayO1zCcbYMfITYwED6RuT
N/CHr0jTPDk5KLOWq/p8mweHcvdku/J1u8XD+x+WUDLnJufbDXfTXSfVYjWCinsHeFhWStrSKbtm
SVHiPFpwLV6ioTfGzAms+zI4ueyV6hd9NURHY5cIJ5Z7s0bpC3KglkhWZ3NJqy/Zl/jQpyaIwP+S
fhrOC41FCdO5Z/wunhrwz/JYV++K8usAe0CC4XMbj3rGRRTJD2k3sOJxpo2wWrg3oPLsczdV95c8
W8zn6gD3Ctk3ioGtpZKqFdLZrGl74m06Yy4IqcBHTBqT2ewJ8r5hagLEnIard+nrAotYf7YCGL3j
5FdfqxzraFbR2IQBhtSF9ljr+3YPSGUptt7i0wmD7am0awNZti43pD3ZJnWRQG2FDUCbfBSoGIt1
kQ/CjebXf1FbyCrEAdKB/wf9vhBFu8lNian3FgFiq3BbFrBeImJ5lTyApTXJ/d+SBqksdxl77Tuw
Fw+HsvI3ApoQzs3eV6Y3L+QWryu+5Fd5QaNwabybQcZcCWfHxDFf/JlBW0p1nBLn8d+Be95hzTVi
0JAFLrb6PRKqno2NUo9w7tx4traDEXZcU6CAR8bWHCcVZuKQkcqTPZ3sljq/nQVWXH5/1j3uRGId
dKQ6lsrvDBD8bgTzf8jcKq2zwCsJRIpHyBcUhD3aVoBonPR1z4OjQ/+vewt0jaaSG+uCHDnYFDFz
zykdgqHNGVuXjDMf2qdCWCLM0Ct8CzbIcsJUBEiLqR/QXQYRcNKaKfxs3CxlO68utKimqE3Q6foW
M8yKGC2X44P9okKowy9eilSTS5/0Lfzspu3P4snU5TOuCGuBYi0qar8sxkmHNcu9jjhO5jKKjFT4
42Aj1t7z1wM0Wjg7CUG0yFbIOkgIGi/DVgtKiCJGe+fe1/4pdYhr/TlGGSORf9P1NuPopiZSoidS
JC4ezdPSHDvtSRoNXNDuXRFkYN5PGw5cfCx11fK8YIcBN7VTNgYC9thG+NgXL7KFbpo2kEsZljOf
OFLwj/T5K5vRYtfKyQOIsJ0PXS32cWXJz4vuL8PhTKy1Vx0oFJ9OkFq77CHrczQtf+pI5q2/ldcV
ZKya4K1VfCQKDIEStzXTa0ZHuUc/vnLugT+451HhodC+1UsBVSnWyySWRvzWKeuSNDbemB+rTvL2
Rh52g2zFejOpcNqEdu4QI4lAwJB3XYIDXXs3+0GySE0u439JCpI9u4sxrX0g1xz1EE5yQfV6ZgsN
lCrSxl2Juz1gmf0MU5FDDf4o2SKNcIcT6p2ZcTz9AYgJJMZVtI2AV3iQVTRSp8/tRqPOvKkFuy3c
8jhOduFc4NXGBBAkw1UBpNP61GaGLudn3dSfwpLubRaqXXk0FVwf3tsGdTsiKCnt7DDgvuJGunYn
5BfcZfUk9kMNWvw/sd807eW7Iha0g+G+XNGbnUdV8klJnnS8mgFEMhd0GWQRIjS3EgFAgFDYC3Ls
KyoPzG6pe1xqssLenTPp0ZnVNzvnA//PrTUVvsEXtIp0WiPBm/NK4wg197fi+crFT9NhcWlgNDJ/
dpPChKqCyDk1JRIPu3dffIz+HW4tJhKJJubd0zLyyI/jimAUhmp3E0Zni+N1tlAHxrPc8xCOIjAU
FelCuHNianhJSkELWaS+pp/7Fx3FSBNCA0mEk0i7vLICJAUTY+GH5d8txVzFTP229lpJQ8C6Pliy
OFETDyQraJtgFSn5w1Qp1VUBe7iVp3h0vSt3gWoHuMCcyB/iWTlz+mXh4PVqCgk5iTlDbOdcOPyV
Qdji7Cuc0VJ4DuaAo+HvWs3GjZQWPmb4VzC2OpB/1T/hJU7FGFiGfsK9JS8K2H9uExeKegwjxNET
TSLEoS7wWhQqpXZA8kmW9zjGtdhKqMnBbYXlRC0x+XnDL4rfMXbs7Ush1eS0IGLhdvvHT6XOMeAN
saMbdJB/OxmTTuSn+vhk6YquBRYd8AKJ69zNS2ljlzPakEYZ5oo2MZ8P15SGJxWceVmCvjeAjaZ9
wth2z6PFngBBBcOBGJxqKInE0b1J8kuD8mllVWUlucNIEjM1oCw3ZxJkVYL+KL+0ybLyEDqjbhWC
DrGOF1yyZZBOlJhRXEHXBdrn4HOthZrvu1UuvMG93desrT+8sb643U70zOODrSyLxlKHh3smH+7U
Q0sVJprQWBdJXWMvnMVYvC2NBSRAeR4x2xw98F0dHvPkwc7d4f9GNZoOv5Exep9rWPHjldAQVLgS
u1euVYZBaaBMpX9etsBdZtpgmbAM2pXg35MxtH0KHmVCATePbZKzocvZdWdn9/wjt8tHHIs2hPVp
mVtTztLzm1ZcdvNVF1iUb4OTFijp1E5FYCp5eaCPqCFOGo6sqG4WLUrPzOhwvi5RbnI+1053PH4H
ByYC+85Uz993nm09tM9NWDp09e2a1hwxrH9SG0C+pAaP7k18NBIm6qtadPpN1K8oIz+WFvbm5caz
YdcEevNXRfH1TZVfsQJQkp0UporFJlKKXAFGK+NOGvza4bpBNNiU5cF9RlS08oHqg+PG8M77qbJd
s9yQmjWgt9OqPqkgTMem9l95wIx3ha+mrayHzcHMjcisXjlIKhmCnryKkr2CE63ABkSm9qTcg3Ry
siYZRQrS8Rx86VuW1Uz0AjL03NSdfynM3MpnXSv2GKWvn2GY5lHCMmUvRbm8cEfDi0/u7mbv+ZxZ
20I/XtIkL+8koKqN+OyBJaBVEbGOvzsBBRz3rdJtfNXTg6aSZN1bscHmhxYPVTnCL+uTdohE2Due
7cGAm/3Cp6h/kHjC4H+c2v7YjY6BTyoerek8QxNRXvwiBHX+XTE2MOZ0im7yAPjNKWxfor4MBn4t
hAiAM3gIlQp+2lkXGlXV7rdwhE95AZfNoYQDZeAFS5aTsGW+Gsd48oIOUF22u3OeLEgjN+cTWVIN
0CRXvMu+ZL5JVPt2N5tVDnsSDz5UzCVskq65THJXaLXMav+wDXQRTCWLJ0fuxAGUA2QCErBML9wt
vcJ37QkYb1ZmuGCCJlsIu6nEAgLOBa462jmC1LxoxGGqrXRUkocGOts/uxd9IVncGLOyiW6/mJGt
yE9kWbsEj2+6+SfKORhvsmtq+mjctZtAuXjfsprcxTupIwCCYhOatrbirK32PsDRNqBgx50AW9pB
p1+68fQy8WOmZDfj8GUX93c710u0g852pijFke0pnj4KDFR3m5NCR6cIuQ3AQ/JqrF9geByVbGpN
PRphexeqKo4thwqco7TR648U7p/Q5LJX7vf0j02JZ9Q3TrAFPfpie9YGRmSaDJpvDcuUCfVH7ZZL
J7bi+Iiab02vcKLKz4SfacCrcc9yz+JE/Qj1tC7OVwf0/QKO2d2uhR3LRL0wwulKS58FGvvBKIwz
EPjaXlmV792khXbklvh9pWs4WpI153hRy7E2Ychnmptp4M2Eu7W8b84iv8Ap8RYHPd9V0FLAp4Uy
hs0Ba+1W1D7ox3VSU0+9bwfx5swxRev/+WO6eNaosbyXsUEKTEfFeKmzuGBLlHG9Nw97GHioG6fI
wmZtNgG6FypJH4aIoQKT1qh5OL+u+eMu8tLGLHHDZJy2Y43BvdmrEfwCGK0mcboY/JWhPnPKcOD3
p5FklrYbLQlMobTUxqvW0NsmO1t9cLpLFIOBHAF0HUQE+p7OMR5gUm/lsqWVIfegqm++4dC6u3+h
kiyL8PQSOP2XELEWCThlD1VVRZ9ws0yxXuddyDhOgm+SuAHDhUfmPDEtRKCdnMF2pCiWvIwqrbPU
84YPpfULE+Hyob9RlK6WVZjczEGOttDBlvKzg2+4LgZ6C9+3WsZPtiEnpNAHNf8fOW9+f2MOeR5z
3gtdspGEKiqWqSfGqo6CkS0ykKuesCxe18MnoeFScE3nlErnUsDJRg2zXMbAZACiO4MYoQZZQVTB
kcmB1JtGTwwPaKg9pLgAoXMIjhVc9E0cq4VGhH24U5Ie/QMOEThYmm4PSVS19q5vW/6iVgS2rKgG
xWBd4Zpe/PDdKc/HMp45AY91GiKXpUJmN1yVlJdl+E00t6wrjPBRSUw3VTtFjnxQOAaZsA7z9xbr
FyCYy1lq8LlUnFgYjqlc652GVnQPycM9ttMwTOYbo2B03rNLUPnzAgbs81OTkMq8dB91aDWHHmu1
rguRDRPQB5IvfpKxbHv9ePPew7IAzu5pOQFxT6RouvqHoLUxO84UZD5W1JfB0httNNIz7HiS81Kz
dRM7QcBbXCp5wZSXjEaXbivckQSVSftwiTBAIEHPTVwzeG6A0Qe719u8y1jSfaESKtWr2gdyOR7e
Pp6AfCeaDr4q3UJyh/qcKasxZAhucN5tLbpzgoKKdvlla71yYbDjI+zx8PgpJwYkP3E8qpMrbgHe
vBi5sFM30jCkFsK1wIc0UgPbT25DIE4hflB96NjbKw+iOP+za9WCEQetkHhcNaLgqKnnJkg4nknj
As9lJZ4gye/cKR1r31zdzZJ/lnrundtstxQu0PN0sVzS2OxeVATf710bcZyDyUR23R5//ZmiKw69
TIYZP+dSZBKcwDV0LPeC8EmsNVFOFCIOo7K8n9lTXHH2XjEXaJKRxYWak0vQmp5JsdoYsCc2Cnic
b3gblAIffCIhvvZgxH8NR3dDxzb/T8xI6rXNK+74tgSiRAU5iMegqH9nkyu0h2vJTHqMnnYTOqVq
x2iA5vYx0SBVcorv5KWvpxwvV+ubFMRSnehoUOzzurmSIgTUkBITLOh7sNAwkAu8//brNKjRZXaZ
RXtfFj5nteU0+RgtGGRiPOt+MkIvrkiylvsEmnYbKym0jV4muF6LUz6XN2VSArnOE+ur4t1CYLWs
SIPrObmAL9eyvBhuSPi6EVhb7FBf1hM59eBVr4iMwGB5mDyqjtXgnHJ3I/j6hhIa6Y2EOKjCHCOp
fCUsPxJ7LKUqptuvGVNEKBLoyC9GmsT8n61kQ8K1y5A9eJ2IuRQFjD4pOoko46EMclcD3IjTxXLq
rsoKMq8AfnLk2CcgSP5hSTP8RcALq0mMoxGTEXKqG/75Np1knsbsMv8ygVJuZmN4VYnPrZeknF+q
Uet8BP/2SYFODdP+Yi1n6dGWhiaoY/tyRFi0dqMZsfDNIMp+FNPybl88y1y/yYZOGDPpn5gZYGoC
hiXh2pCa4ywWjDq+0srU+kb2l1z8e+H8Kvekp/9ZgZ3LSqyb2uIKtrd+KwGQakv6b+D89jLMst5y
cPFczv9chiJedGXHd7g0EPa7l1WSXIugaefhy3Qm2Vadkfec8w5d5fBKXx1QGD3hsLifd/i2cg43
kUBXxfme05AJlKSfja3Q3ocd3gr0hT3Vkviuu5RkfwtLzqIYfZe8W6+FtFCCeXar/7LZFn03JIzF
56euSl6kJXQqTGKjPEcMg6mJl1x1//sO3oYfY01eR+FHnBFvGB29PwL08k6A1Q7CBEA+mnGSukOy
Fm8qRq5xQ5sDwOHIrqfbvrEvwpS5w3SFLnqMnHTfqXoIBAvjmbLFrq10w6gWwiwCwTkb/5aNqo2U
Bo0/KQHQmAkL5Bv220FzNySWSX5/6zoaaq/ljBJ6A4XLNKnaFkUczujuxEmpuJV6O/t8KeEGTQ6M
WBcM2yH9v+4DjVQ3JifX5l/BEh0BFFYR4DYGH4jHWniDGsLUXQqB8vAZ3nDvf7MjCxKvCoVRhX9q
RO034OPm8csDazL9o9EOERRYbScKCd+QkXOkeU10PlKMPay04ObYIGjXOhHPrCKJ2wUPRjGVdVEs
fw4D53CFdwuE5jfmL8gr4j4KXMFEVvfrFOz82gg/KZYK0ykyt2L51GrdjehUL5nkzv+qo4Cf2yEy
KZrz58DIANOojL4cjW6CyHXvEmtv2Grpasw0JOSUslStbjnudKR0FG1QL3WsZ6fuwUhL8cdH0O7D
hHbnAkKPfq5CB7+3gLzqR4NOMEsW0tKveQHLmV7Lnz4fpK7a0tvfFLzx+GdoFujKH302pzQS2nGI
X5uc4j8xsGI9DwiLskPUL9FbLKfRt4UokXFYf57VeGzgDZ3VPmq5BiBgBdIfgyUP0/lgRqfjkDHH
riE5cqHU4KgzeurdBloG7Er9r9kM1hYJGaI0TAFDfxRYijei1o20KhFWiIDTQ48RmpDBT0tG7Kkr
L8D2mBwny4bC6S9kIOvyzkJ4CIW+qV2AQAtIEHLgfKSmxZmYOwNMpoMIwK9CtbEiw8BiZshpIz1g
wRVpiNyAS2ZeVEo3TZmufuZxgRPQ++o+dMWiTINXkM3MrmEriyjjAc7B6bN0iv5jCm+lrKo7FJTt
ExVmmP+EOloFfHCt/2dUUYpiGgR5ym5kxdRjL4uku0tGBX6OKKUdu8yEGWMVcayLxlilZINSNNoX
bv0hta+6Fw4yHk/2o8KGEuCxKsVZgNTIBku3BqWF5KK6T3SVsjMdUEEsdkd5hCzL0KgJCHkWxB27
4I6bqUHKBy/f6Ol5wXIXNwfpiinSPmndRcA8uOUvWdMJtPSsoYIU/OswSqRGBc5OIHGxg0F2rG9j
sknlRq58lXcx6WaHr7N0KE6bO5a303M1CclOuYKmdH/jKrecDLHir38aFphzOfCIpc+vJidIBtgv
eUFfN45tw45AtBg9+8CuDuiJksCo2ZDq9+5ce9RjC/nLHMpWB2hze40irj36xqVVzvuAK60kuC1r
2un6jheA0fK0wI5hYDIedn4zE5Nn3aVnueLvM25KqB3tR5qQ2lHidTaPD4SbwWti5NbYvOUOuNq7
KoyYnp8tvH3n1Z6Bhv6YfBtsR1HCAXDLW2svzfzxhTjYAPhPCJi/IEcieGx/rt8IcRGA3lYnk+ut
SwvvXs40h0o7AGUHOHbw1LxzxptESo48r6rASREmQ5iBrt5+dGH82OUca3vK7YC3DRvhtetudntv
FtoLS78tkZnfqIFTAw/9j7Q8YJYqU8Q+NwKAc+MneoqrKVrG+i0V+Z1leqdVLvnJRUmKkxVtMljP
5wMHo0Z9PqYoby0kctfW6K9+n4ArQ8Vzh7vcT1mrjnM1EAX+CLYQDXA02/mlvaUOPrBVA60hM/AB
tWsuEA+PILx6nVJqpY/rnxEq8FTxi8NcAoMc0FiRRkY/oGkmc4c6PFTjU6mCScTFS0i5Fp5qyPau
FyP+HYU0niucLz1mnbwqVR9E2cPAPMpYJtfWeMjlkp9JOSKSG/mNPCsavu3VPLi06KltcFpxRaCX
yZjoA/rj9ZdI0+hN8UKpcuNFCapTLHq9OqopCGw9dIHD7c8V1+/C9jn5BeC9V9TQpu5+kgHpDv3h
P0U0CUAw6nYAAlo9JRKg0wQNtRXmiUt2YUrWMrOq6PzZ5c5RxLJaDz+pVlrlfq4GR4me1yQekM2r
iybH8MBgdVUrxdzHZ10FNYNkQ8UaYHdAxtGAE3kdfeDqMPeMzebI+QNY/55UerHjusF10K/JthIz
D52xjGhbbjFHeThhSplF/z3sbuYcPfKYB9YUCZ9PF/K+xXzYpZLcToOjJsTVyH/qoXbW1oxjK4cF
5aye/wIdZOokzDwCZCR0B9e8uVrMD6XM2kf/3LatG699CdwSOIGAEVTMGdhxn8Y7GSwtXCOAGjxJ
QtKW/T0w4G+xoosGcjVe3rtHrU0+FgUQ5ybdsX2Dedd50sptM3lro0ZmXeIZA2QPD4TNrtVRM6PZ
esgfjLp3oDJxErK0H+7BzNr3uuAqbFWSJroWpjN9g+Pxy5Bl/sUbs96x7XEH9P38gg5X2piNry96
3C7M/cKPwwOcVowuE3K6Yiy90G0MFf3itDUD4htyHaHcqcL5KJ3NHmn4Hy6tGbZWpdRTbgNXmk+s
zkp1RlZ3JDuape5Uwnc6oxQl1evPfdFTdIGedPR5UwLfsC0cpTyJJlJzXuRJdvYDegjvKb3AUZDW
HzqpPavHCaE1yrA17GUqhdiiWn8PXxq6NzmQnKPWndfwVszzZqmHDgoUbGS4tscFxiSFVI07tHws
cfnXF/lQA8UsXO/p/clAegKxoilTWFXVB4cu4sIPQUAJ5RhXKQcZn71vda87SFZcDO8YzPwIyzBV
qp4p21LFizQksP8Bfgk5W6XRP3ILe/LUom9pV+1dXMlEzh/T8NIEG44IYLYWQEx0Zszai8xyRhgo
AJlNUVfLNMfLdlFMH0op53YRZ8G/KCSHpWila//TzPpWxOxhYScfj4h84qkkrHJwKm1Ywh5vXXP7
w/tdJ198nLyQRASxEMz8xlLXAMou+2x77Thra1naRDZCkQJLm2KGFn9kBqIBt7FN6Y4s9qKvdszb
rBGsf+hlBjWhYebZgbm+Y9Qys259wbiqjUAF5bAZId+3S43a0zzR2Fd1hN9RT3Lc5EGfiZ4b4NpZ
6xIDOpFUXmJYLkFLmGEiXrbTxbxYEM46UAGHTQ6kS7o9nUZvUobFpieV4+49PLwGZdPIjnymfkOE
Y9y2e+vGoKHnc/xECRBcvhM5jSVSKRv1wB+i/FOgHLjga7BZZsLGLfX/HupCIQJ6WJNc3VnIj5Qi
oz1CAz/32OSkWsWGys/3YUgNCLAFMNVmbgMKSfA/L06lKjM+un6T20yWGs1F2piXQjBCD8dVk/9b
VOzlaysmRO5mDLeZZwTIz3Ahs8UhVYQg+vud9qjPnRViECAo4+fHkGpT9WA8OuyF93DwGyAP4wHN
A6U/EOKc5EXkKLlkcwpd8jt70zePTEX2O3i6sVDwq6gefEn7R4Z5MnPfL+5wW/UcX3WmHPe2RQZl
LPemHxvtsNUS81prmaiUHfB49UnF8lDA+LJpdvd0xEZoVenTSYWFq2/qgEqf45yVNcLEG8APlkNm
oCnTl5TMUXvunDW01mzvnmjZna9c0/s2x4kr8kOymcjVbFrMdtILLyfoLb6cBgfN4RLDbarvYJJc
wL3vZiRc2o+9kWZs4MLtyXb4rRUC6OK3WBmoQO0zW7NYzcFNjuXFSpLIh4Zx2qhK8O4NocEO04hK
/yPKxCzUUaNXSzlGHcYvCsdP1KZrQeDWCqKT1Ml401hZjgEPuJkb25/fKTWAPovQHV3fvqTIMGSI
HDBF2sKJdpOHyceLKsGq7sGlJdmanvXa86TP0rJ/CGCh6FbQXDCKIh8KZsjmu0x6f+XRgD8yVxh+
BXC2SucUkQCoMy6rDJBB4UF8LVXbOWtYE/90qt36/t1gySVFUon9qfo2FdAqbYY6RyzxrpOsog2G
J1Vtz72mROVUPdjiNjNrz6RwR9g2VwdoowTbo3IcsGD3dJB8TGaypai75l0OmmMQRqzEdJ7pM+Cb
ZL9UMVL/a0dwtWxFS15HLyJpjIAwAeuYpRgMesjHpTOo29aFO5vZM3AJiofDI3w6xetec+fJVOQ6
ipkYei0iFDTv77OjMkuG3N2N1sPIhekQBVONZVQNU1B+rAIeTjgYo2PmPO4Gp/4dTDj+15jfh2Wc
Gh3GL5xa8Un2KPWGtfjgMVwZy6OVUjyJs2KDF575NgC8c33Vw+Gf9LhdPNpIQebQaSCrPmb2iffP
b6IKEeF0iH9hNIlZt7eT1VQrBMuJCHYNgUzrwmc2BlRdciHxfdXUdnWiG5vwbjv6xrNSyIhfu5Ce
YWrfdT4RthimIgHCJX3bWfTR2xFQCq2e54DIp3ziYZivai6pXG0xfa/wf8MbR2l8QGPFgjYsu45b
XPpIVmjC5eatVXXdfBxhPuVGxFyjHsAqPSimemCjlFnWOUSDTHQI4UDc5Q3bT09CWVCATduCSPOI
0sA5GfJ+bf+w6vmsBPohraG/YQeyzBkZzkRfiP16heDoWhhEHaQrEjWmZJ/YyWPULe8TvaoNBl5O
HzbXH3C9lUooHqiVXmOK5hsv4iAkiNGXJdZibrBe5WfmWhUUyNNFXuS2fhxLBNPoEWzuwyVshpKv
0DBB249zNY40T/p6OhnCE6Qqep/idnFWAQfzyXYqpqkCdWuhhaHszrGfe88EwhvuWkCiJ3llGjQR
yenM4UtmSXaMu8uIIi6A+9T7EyK0CCDXtsNckOLfKhIsbbzSF9y/L4BQrInNUDGnKvM9wdlDxhAk
0pMMoGcLsYt2BdbjBNSWUs4p8QyDJyyPsZQIhWGHed6K6/w/gtlw+6y3oktMNofikzubYGfsTi9U
AYj9IIfp6Jq1j35t5sSxnAQQO0DqHM6p6rzeLqb7q1oqcMlGSX82YVx8105p+JI8jsMT10EbBm0u
y0Vj0j8X8fvOTsBgukoPpDjbzJoG5kjUITBDBvnfr6xkTCKb2SvXyL75QlhoWUTBCmt1nQc+s5N6
Qkh4tCv3Gn18rz0XyO9/HSFBDyPkQM/TPlaZBB6aHBepZ4UaOsdkKW7ttak59x0ZsVCYBOc5X0LT
u/K2NsAdwvKtJhVph8otvGToVPXjTbJDjX2H2Et6M32hetcsgmkxb+P+fBx5o042Pl2HEzWDMpOp
fHIw55/fPPAnWcYrkIvVTIdXSz02tdEQsAex5LbNNj6dx1ZPGfQeL/qDqFPUJCiclHTxmsQUQj8E
lfiZq7EiM1fnXnpaeLcjJ94CvnKD7XFgFV0oOyj9uzIkQhpttnsNcOopd2sMKBKx+FZRevI2sczk
6pfQJuw4L2qPab5duamA5T+2ynHNgii1Af02Eu4fYE38jdEdTkwlRYj0HQ+Py4mkYTDLHlWefC6E
1LGQ7ag03pl303qWcmYlsxdHe6GYEMOGKSFKngx33UkpYgamA+bKqkrTQv9kwmjciI0L+VwBiI1S
Co30oV/U6NRloJP24WCsYxZ8LxMTSKuHxe7jogGfoXLnLvmAptidOk5eCzc4PjY/tU3/tijn5wZr
bSoTgjoM98K/5B79+ACi5PZHHMTpY2N/+PUN78BxM0GFKQUHhYBwL/vfLyiVEQdW6J5tq529M6Rx
uptvvElNfYUfTisMALbrwagvEg8hItBLdu+JsoTwMTttoBXsQFOeGVNJFov5h63akmKoB/gJV0S6
MarRUfDwplFPh+0KDfMEzZUEAr2fGgrIAEto7swGNmZ15x0lg3cgKtIS8PP9AvJ4KZNh4LlHKx5v
jNcjjmTTtVi0UOQdqZsEw1ur85qti2avJ/h+FKhRUwxcCkIIIOghcnzvNGezAlzYbFuFueWocRE5
OPfGhP7lQhJvtxvHT9vtQA4g7PznZPoeutJPuZfgzsUs6fek91FRGNuVMaHAis5JTXQ+/TDX+6bC
3bNSsFC/eBk9EUEe6PIS7mQOj1ffQL9d6FL1wbgbKJVyGKTcjoogjVlI8IaWa33atZZHzoXBsn3P
TN1Tl6xX4vd4gaAuzFqZ3CPUIAc/KiP29OuyBKr7JSc3wzvfOlJyi+FD7Vy11uHib3VdabKt+r1Y
WmljioH8krEMP5ZQDxfh/+ZiWkjT4yO/F+KQ761eP/Z8WI8VxK0+uPAg9ugNHuZqLGIEDvVH+2OO
aWXM7ETka9/iY3qL+FIuNBpfdunrF9fHFYj0OVsT7hYrn8U7owSzXzhe/3DCuqBJRsymSc05HIPa
lr20JPnry9/PPH4WKHosTcaSY1Sv+PPN5lyZ5UMP1hkddXmMN2VJhRy/fVF8djFwZ0wGCs50x/3A
xvytJtqax+2dGcqFbkgWIgvjrqupE88CkG+Uuq5iSiYVbVErrt5W6ba9jNEdWoroJPTiHFPW5y3E
1cdLd59x6uPdAbt6w1qwW1IwRykYns8RCEdmQ9gGhsxM+FF/85fl/3vlS0fkjbORh520QFBKjXz6
cQ3kfoUK76rWARUmu0WRcy8RMWPpmWHO+qoWPCMiLDbBmriUwVM6iL9CwTp4UhqyLnMMwt2CRuMf
cIjxWvBaDT2CuFpaJDP4xmqTQceQOTy+b5XR7Dgqsx7JCJaKgHOX2nphxxMcz0JgUUyPc8c4/vuE
3oTpG41bcQHLS+UZywuj5pVB+P2DtXXBSc2Vy3oMpIgJTsGsztjppxN2E8ot2eW7IyumMhRueKmH
FD2xznVnGzc/YQWlrMg7lKWVnMlTsmnmGtdiXuMLPGGjbhAN8x/sH1+/zvTUcDxArShGi7iQR2en
fVZK0T0vNAT3peHMRbt9il8qI6xLJhu2xrpWgTrjFePQKUmP1hVEJFpLfOWWOHtrz0R40SwnS/yS
r/Dj0kf4r0QlgET6HcqjKUbWUKdpQFlRC6JyXLIe00StTsGo7layWVd47ppZD19YkQHbH3VHZm5s
1aTvYe9koMMo8FWbGUBRq3XWL7j+rGnbtMk8RgJb84SU6x9D10Wp0LO4JT1GBKh2Qm79kx76QgZx
v24MT+CmAlFVraUv9X6rImq0l9F59RR7XIl1AAM7cKVEq7eSbesL5sn4lhdfXStHNk1F/IB5yDfO
httCXy3myoXqVS7nOhPHZq3VAExaTMfomxrGzLrliBp5dMOKXzKb8EB+DpXZk/Z7PNI/FGSfS7Vo
LQt1GYYw2gZtS/7DbcipUHnx9r3HVPhVFKNvdYnn5MJND0B0lj5fQb1uxC4Uncqjk05Qq1zd7xRn
EJcMD4pSWQKJTx+35n96Aa6BlPtkKIdh4aKsgdZFNnLZxAMzf3U5lkUNyKS8l5IBqbODiZDMJklK
wUeynQByBN/itVlP9E7uifK2c4x27F4uGP4tz1hzBxrixaUd5XI4wyAeSN/cge1wuvaLpwJFru5j
ldrKyoPC5LnBsEf1wJBLraZRG3D8UVh7oAwIgfBVg8DWl+O5QuLfKnu9GMbUdr98U7NvcACRR6Hf
8CXwEoP5L/m/DM5KG2rFjuNZeqme0tMgxMlFE0arz12vLicfefmgw0PQ2ISxvnl6HNrIbs2OyRtT
WwiM38Q/WB6W/sACs5CSHpEY1hSxUyi3/jywrGQbuQvpH0LXaLHK/gRaxhPhpd7VVF9fL4hF2B1b
1ZQO8AfGa1bjt2hcIUBVLuaaoFkj5LaICLXoLo/qDOdGVksKnEiqeE/6NsCoYAxBi8DNd6Z/Ymt5
jrLDc2Jt9OfJCIi5FEBicRmZbB1c8O9TQJbzwSKBoZMcZkoP8CNvrXR5pdYrCv4uu915ftgAWJDB
x5s5NpweB9AQYylNFHYltqOXBlUxnc3hulI99XQ1crNhsvKqM/n0V0PaaWLEvdgqf0DAUpcE0XQN
u/1pInCQh/e0FEYLNMOiDL7ZZhK3DL/foBhotsEZoSf2aim4PwNC4/tkibbzhDvdmQ2WamLyiy9H
RVorQLMZ2I9xbKVzB04meg79AyaIEe+szn2lbukBKiwALYlyyhFZGY63T1vgSTQCLEnT8wSfravi
0SFji+AXI6reLBacW7t5/gdj4linSmXEQm00B+HLpcFRQ8acLk2VzSdjEyCsXsKouUTg7In5/2pu
MNPkotpifJEMnqW/DyRnEifv39VyqzTA/NF63iCA2QvAmMMdxtt0YLkeq2FJipdGCHelAHPNyHM0
qtmwKyO5Heu73nTvFVLzcqDLAYJ870P3gV+GmfzvG90k3vW1ziJ4b2Y7aPhZRr2r0c5kMKbY5a3i
cYcMW5LLUNuHj/Ni4SHD4QC5YklpmMCz6hpGtbTBhg68cpe23b8pinCVpiqduYyLYGmeVnFOmx2L
0NjL/dSPhNFzbxgDVfpK8Hgfc9OHRK7dm9W7+0ZC5ZStiZalhvooqMjRxMwyzrq2Dp8QeNYPQZ1U
iLaYbOl4IRqSjck4R409PGBkryZXcsvQ2d9KZif9whUSzAjtOpNCMAtg0hxb2XdBoMhU1KwJo5Ay
ZrtM9ne2MgPDYzXJoe0WGTqJCjtZMD6trG+mapMdsAXS7uvR7tc7EC/yMUf+B0K2f7L4fnjbkypV
Y+Qy8wId5Bt9ONAZLRPXRVLA63k262TUUyJAsuE2JfEnzcGGHlDgFVBIdPETXakuLJLrFI3ra6q6
Xms0d1CTFvW9e8jiREusBTXjbjGmCfdpjGOxGWFvaCRZCS2/VkIYFS1JYJv3HPAFdHA+lnJBS+g9
POle1NugLmWo69kS/ZMAWbJPLhglK6hQhyXi+CPLaNz5wzamkg3i/n1jGzvLZeq6BSEjx1+RaNHA
r0qJ8FOplJSlVC4xHf6w0AxGiEuHO5ClCb8xr1jJmPdKSBjKwGdKLThelGkYApq9PBwCAfgULNmi
2feJO3zwq2XtAatakM60JHOb0wOWuhP17ar9j96iEFbpKKjJhoAC/uqRuSjz5vzaHYBceanlSxdm
HR0Sqlb+yyKvqL4xOdurZW4KtE1tynqzugJCmZPGO5gYRlKywOvcJc8uNLRZnY8+EFVnyUi8s/Tk
00r0Txiq0aWMyy+DIQdR/sVyqzSp69eMYplvElYevxl80TDbRoxoDbsW5DPFTDKXxE5hyN+dT/pG
+9JcDTmyHZ9lvIfFn1MVTU4u2tFGUGJk+oxu9bsdc1R9/z56s9HJAJRXVzSb9XzKJB9629bjiLk8
WvRNWBiys1GPnZk83tOtxJcsNoDWDF+emC9WkgBtXQcY4vZvnSnEx2vdQYjnSGoZ1bb+Vd0BIS2D
NdSK/nH5gt6L/EowERA5IHGrRrj8/i8kW898DHYq3OH22eK1tUTYnundP7PJDl6rrRndiTNqNO+u
zSEi817KaUGYgGH8Cs/rZ+RZ8AXhDUVYfWOBGcpbTyhhZoUFNzRyGoaXwNsCUEyH1J5V1cwoErG2
0bWr+ajxFrluJAZa8bXE/PRZGIxz4NGgy9w/qpmHtROOfAmS2oFKbq0+Zhi52EVq/X+K7vsoKjlD
ecpcuxczmqsXnjRNyhKvN/38FbOrDEUJ8mjhQ3YN+UWYRCX9gZrpX6iowb6oicaer9EV+iIkevF7
ttK8njqXncMMrTT+5zOBrYMQzhqf/qLM6CAJuFg6gv2eeyTXF7u1QSIyXNX8YWSg4qOJI6dtnYcr
nMJ6jrEhG6qVdMy5f80OF2Pjg1m/oROUc4yCOFla7lNaAZS4GNpQadZOnyMjNaIQKVtIhhh6xbcz
5MAZQWoIQx3FqjgzsN8V/7/VXkCUOsf3qrbkdW3m2hLkgB1nU/X1wU0rbGcZGaR+GhvCEcUgRvnI
YoJ5nWrnx2o/oV++e2kCEbmv2x2f0duMS7AurZQX97alqUjJh50TEXiIWzc5CO051Vrlp8+pkKwX
UYIUn5KyEW2GBR8Za8m7ts/LYgFirYef8QObAlpCta3Qxov++JztZcjbQb+zJvlCuiUmt80UDouO
0hVBHq8ktwcrkI4wxTgOAq1QRo+mIrZX4RANO6Q9MplGKGi+/9mE0x9I/OUyuz/JEjs5Hvb3KlGh
jHcrWATV1W8IX4n1UVBFx8fifoz7yoKKYcMT6+46vnqvtkxPV7GLiRlrhxzn7vOC+FFusUhxLO/5
ygewnSNMgzqm+KmKYDxwh06wnGo9Rer3Le9fW/00yzAy4bXjbscW/NFA2Y6XxqOdfa/Ah/wEYHYu
IKVATL3Tlwi7Lcm4rU91D51YGmfKySlLfsDu0oC3Z0WxZoe65fiBToa3b/P5NskZepLoeWZVhtVR
6FRCeJwR0vtaFedk/135BbpSuyQPyulYGwJGFF8TJscWhULadQ36n7muepa1Xx7hvbC62dLKXZ4K
8M5C7Uja6MFLsSoGWs38GsQUpkOW2NdvJPTudsNIw+66F52MDnf2w6T2YuvcSg660kB8to9CVwQw
v29joo/BgAU48RhjpudXXXLZjblHnIA6j+hIO0vnE0g+d8yxsMv48VallC8v+ZACtx5zPN1YnMaB
yX6Lj4th0RIStOjWyouIoumJQ1ss+dtPemt9BFy18rwfFTCAsj/4al3EYR6OEGR/3/jmrTzVE1kw
sccPqhhOMxw0/cun+xZ/JFMnCjphsr+fDc+JqbqWWDSaOE8Gx41w1zw0MT4ZwNJ80rUM57DxpnuA
CBpgHzSMzvdwhCKEtb87EIRDnQiUD7khxTHT65zAouIDOtlTP87seUFRvB/ddL4cXmZPQ1yrvHAa
t6qteMXjTZqnpUmTLvzTW7f6ERYIo6FwAO2yvtnrTe3SiMJPsOSRnJnSrnYfAoIkbPPE6LY4kaP3
H19ZX/sX50rMI5lIGOW2pYtw7Qk8hRRNdStMnd6UcWyDZFJBwoqKQFJbO7yo4ff1R8/l5BWDGoWO
MT6AdfbGX18FG9OXBZ8ougdUlLAKNFVD97aRmSkQmdvIJOPq72qmjnwJIYaM5zrAVtz6t2wQThFo
ZW9Rniow0lkU/tJY73Fypc9S3dh36p/GgvMzzgEU1uqSc39V9/BKJtWi7ZGoxXG/NKvgxLgcAt01
74m0eWgpByt0gjva6WRfJbVq9yJpMc0oOY2yTOW68q4cWqnr8R6NUG0Lt5TxSm0rNfG0tELfUGII
tLLgKCWQTwAp58ubIGhbtW3FAv7WlB819CI5oNq+pTVGuZLIJSEn1FVVsN53yP309WoiEIeszwI8
w/H/RLFZpzDnaBTL29Y45OW+AytMUkUw3+39rq2eS5qfxoh2ZHm4l2hgTR80BS3Wc2pAW1FLQKsf
NzK6qfLk+hT6KYoXFsPSl1K/k9imv3SgnJnj1mZ/sl1RZoqZg5TL9EoqpSm6S2aSYE80oOW6Ebw1
Mjb+PcbmJ2JwVENqY9Vsn65NUqsfYidfOUasNHrDu7LSoKi/blbeMIH1U+ydZhJ7oIFtOAZ4svqg
NjttC5YoXbA7dxlpRAnIDFdrkSguTS8iMe530fIm82ZfV7XbN9AChFejTVYbKDWQVBHmtCMK//bf
9ShUbhDXn7V1DrB9zJn65bw1PurM1eL5Oh3Mm3VM7xwCxmWNaTVeSq+aMn5cnl3NIzgxzuDF3av+
IBFFl5PXkrbCfRs31xEkVLDTTgUPArn3+Kwn1yDPNqKaF6KrhCCij6URo1VGqppDOSyocwa/cHPm
oBW8doDB942ND95sfkEChYn5P3wq7XoH2X6sBrA8BV3/suUtdSQ0om4azCv+tYR8mYkXA0v7HDDf
Y03sp5E54ub/FiECWZ5eNf9qACTD6t++L/gFP0c3IdhyyaXJSpqi9J5npuvrd9VmHrwWAOxP2KKK
tS4UWoJwstDBSrOE6TuDjjSschs2vLTg/YqaZl05c0zSdPv7nqEeFYa4xTkfJ3/DK+7aaoLm6oYJ
LRx9HhhFaCGirwTt3hgDhC6mzYb0Fksp2WtvFo0XPfNpw6xyS3VRhTSzXmZyRJfIfLkY+vMHWqKI
F7P2ipkn6sTppDr159g65LDkHdntayWY9POisA/lal8p5t07iG3PjSa7YFZY6LLgR6MFVCs9Y1Cz
ikTp+IUJ4j49StH/MKlANNiU5nQ+BKPW08t6guvOcWOqn5vcsaHhlPVmD/0tOsbeo+rnoR1Lrim+
iYnVwe/zTijs4z/AS4PSS0TtWV3MiOLKCHnzlcLGwGHwPOK9KKqCxCHejImzOmEenYXTFVz2rCtG
G4tVRXTiP9slMctCHOXNNxNIOGcqqo9tjFLZWTssQVxVHhubKOgKrVbC26JzIRBJcuSxnit4URla
I2VqqeZt+3mL4ryWoj/kfU4uTdtw0I0gC4j67Kmcs260Om/sLjbKBT4dhx70zTxnU1MSfiq1qVWd
6tF8J71zyiP/Ssw8FmiIAyYIPUFr8iQ8Md3jG3xKfLfi35XFqiU5o0TNm2kMzb5pQcVnyAKf5zla
I9Va5NI7DEiQ55NcBqPGDYiItBn6Y2TF1qZhVvZ7HuCWYaDU9MDY0P4LLVFczfB6h2tFahWMgcOI
s7goCG03POmMCGaDpfW+2Dn5wB9DF+MGnf/eiH5fRvVMF748QaLkL8jYS4p8ZrX4TqoBPHuyFOZV
qIpJIXSws7ckGupUwwKEMzLAPVgiFcUPF3Zjfj3BAYX5GPWtJFyejd2B8p+uc6v63F8agAA6TIUW
s5/m7G+QuXmyr1FTjtydTV3+1csiMesbpvS1lFte9e05Cm1ZR4Z1J0Jlx4TGPgALPfqkSwcW9j+h
olaLCySpRcW7TMwnwMvwkuGousk+zYu0QPm78eSZICnuGDegMkjSluENkiTsCOP3tHRnZv2y7skc
i22NqV+NeeIhOAH+xMyf7bepwmEVsoK5u8wxJx0JE1uH41quOTQD0uiF3LNCLMXWoGh5r4kCU15B
x3FEUUtBTIGyPIy7+IU8Fx5U0JQKgwdY3JJI1Fo6qvLZi71kEeAbqLMjX7LW/Hd+uhg4pEbbjdON
QQpITIC4cdOCCcEO7GjKMvWY8sO/D5bTcV5b9VY2ypn0afZLHt2NtpAVirjDeBlyIYkAOEE9cZ6W
8sbhQdq8ikmFeI61tGShp2vuZ362IoqUntZbZ2m8kXiZAfVAnkCo+CnKRCi7YOcSTsX2ywJc1+6I
oU45d0ppu/fCOJ1n/rNAa7WyO53buyFKlfGNgcYzlAAdbbY0VfdaojqV6EoOH4C97R4Mkecsf9F6
uXIn3XSOHp/gCPl0xPwctU2Y8bJMm3Bp62U7BAure4RbF6PVy7Kzg4ksRBTMuzfOKE60KQOkrNJw
j/GTP7CE4yovgVxO/6npavuD1OOyzj5hK70Iv5vb4ANZL49A5nXFVBjnun9C1QiviFnSmfXLJL5k
XSbpqUc9Y0DbD2+Zf9dJ4V+5xK9GQrcxHRBPBxwiXETWdfoKh0nAIWYZ9iXg/9L4iIAfnejP1ysd
cPKl3kl0dxIfrUJZxZHLKgNPZW/gazFgCDVAtjwxa6EEzzOQJ2BWKdmOvBFfCn4zRdhO0afXo776
Vva2g4gvqdX+44S0EFpD3MYtNilk+WjtJ2FtYUs4dJY8UXEj0u9QwTOGAUXP7t9LAAm4ROXY4rHE
4r/EukC2Wwong9SgJBA4GPH1JOhLA1tAA3EzlPSUeyHVF+8ZxciHTailcu1SqRofxIssi0gNdTGG
b0tZHEwjqb+j5Nx7TCrcIQJVA4/zKKgor2kYeL6CD5zZZBlR7WLQ6BgA/sW47THOFU3yvS4aP0Jh
NYiZu/2a+WPtiIinOxwEsfd1gnFih2uU4F062Wf1dynabjeqLI2uM4p/lAjrR6tSGK/qGPdVzEWn
bl8Dp7WwxqMb+PpBUF0IL+KJnBaD1mhJtxKMtaKdFktkisusf0Y5ksRDDYqzZVozXkve4z3tJwPr
zUdZUwdumjCMR4Uf48aPNCBhOeXvBo1hI5V5CbuhTI+z/lHu7B6x8Vl9b803xBHfbxyAzUNsU3P6
ggeD0jh0HZTKjhzHO1FMt7Lhvw+2aiNdpBK1XsivbrA138HqiuDgMNuk3o9CHwBX9y+SR9JO+Hdi
iMIa6l2CUImdrRhJE9wTaevTXWJfoRhwpGHZra4mI8oPlJJ/6GZZBNyrId4sRZV9VKuK6XvurdHa
2GmFmmbNTMt6n3dOiRuUzjCK+rODOQ6wh6Rdfvb1cv+g3GsMb5Zdb1oNzWBC8AnzJkbbUFHDxgXS
3ZvS+hyMj7anBCnFZn1rqy2bLGh4m7hWPr23Ik7cVeSaRtEnk5pybe/j/xA1NSW64YsXKt9+LxuY
IfgGJvJUDqCCeWZ388pC0twQejL2+x41IA+14E585TlcpqziPyPdqxyPzen/j3GqE4dlEU2uFXcl
AM5d/Q8HYp//AwJlposUXzXY4ymUP7pYp3o855dtH3z3vYFdWVtoMVxqQ8uKk5lQUc++XQRoaB8c
a+PbZUsf8ZegurRCq6L4/aXyHHOscybb6mN4LxNWKNR3iWeV0lU8DzVOHbNidrQWJhz7R0JZ8P0X
B7Utn84cZgqlCThNgeo1hwVCbiFJULYITKUH7y7PhTkG6kq1Nj0NsFTJQ6j0uimSG6Lj0GQkAL+p
9ttqbFLs2AdOu70gniGwY1Xl6BsGnbglFK8SrSGGFn10XK0G+cb3fDQOwKitlmTO63xJxm9RAeba
QVM1rjddsi4eV9jvB0WjniSWd2YIgeBjLFD6YcM9fGQniH7skzknq+RrE6Hb+GmkMRcEK8V9nuYn
zovAsxtfZ6MmzfKRp6Un6h7nFJswCd0tsrp8AJE8s6WUf0oVmF9V61q5s05k92k2eBiPOmpP6eLE
lwY7qIUuT1d+XipumH7BkdFA9RtidBTMWffG3+qlhpaNnops+4bGG+9th9ID+ydix4EnezPZ4KH2
1qO4C31TNTryLS9b4ZPejKiVjs9k2tWFu6S8LsSWjJpBOSw2SUNUDnZ+Nq+2nurac5no++8fNjIk
rJCSMbfrTBNoPcIuRJhil6LjL+8yJiMxPXT5q4zp16epJr6QLGv6gKdDn7P1ss4V76PH+kBgd7uT
xXwFkJ3QGexJ7/kMVcsmz6s0CgrzJ38iD8gzOmJ1/EHpAdVojms/q6Amlxa6h9vsJHrBoWmfAocO
nWrbrB4uzSe7RzXm5Qi7cwgmdgB1RmRXM8vTTI5nf1NkeqnhIWVe3YWqr5ki1o1Wz53Wb9t7Yf+x
b3YFZ7fYCBx9Ne0n0gkQhH54hMui52FSl1JAWpdcXthxo2mHFCBQxkXfD1bHU/3TvadG5xO5QhpN
g8AJFQdaIAt42GDLOiaHZ3DhA5/Br1kJr9LEEAn3J4c42rPs7GhmWoX391wSzw2+lLCamwJzRmF/
LpZ83zpyASz9LYyGUmhCWH6977Qqdxz5+Cl/OFCns0uXDIFcL2kGbqrg5BKzIOJnzbtUDPh06+z2
ZkqqWBVGT9tdUcN/vkJA7GW1Qt4byU7KHwW2bc3xv5Dbn3vdJJRK2dCQ6ZFgYKoJQqwxhtp7NDDL
2TgctwoiEzi8sjAdmBgzpuslcO0mYZgGOJEKhQ9c0XE6VQpCt/52TtvgbVXcVCvVOstYzK43xUXb
ZqSZIKLOqU0czbfGVedAJzUZK1TWSMlvxZydZTax81vbWk3cf7brZT6xHzZPMVccDfehIcKN1mSy
Vub2AMxnG5X2QlPTybioReMiqLvdk76CzCDQGFbmlqDh6muliUeXezrTn5r8zRuWjTEcgx3pAzhm
r0ebDv/+HrEudJRSDKTMjciz0roltVs3ZUXmvRKjFRDVSua71NlDhoG1PnK2EOoYBGdfbD7Jl7Ax
WTvFnJeKuvJ0/FaH5TuFDcv8mdAEDxer4FsUCjNXP00bmvoiPejGQuv3zNYGKO+0KM9Axi7+uz2F
MG7pVTJ2GIbA0g2KyDjmRhPoKl366kVH2jEZCfKb/WzjneLacuJZg0+fVF1MaIKsswPbEYb27wON
dxoxn9SpPWA5ZL8ts0/JLHOhWd7+mjvHNwW67WEkPozA35/oO2NOSXVZvdelYpWjaF06l2r8SN+y
d2ykYfWp2bAwWbL5HNk7oip1s5hYw2DSQrh1jrweXAMnx15WggIZfYXe0CdkfLdZR//Pjhyr08Dr
cW5rHQjzrt92ZLUWB/2sNaVRyQ61s6Je7ZUOoG9GTUu2K87Ejo71QtW2Xf5TKmWirU9ElQ3PNns+
duJofYF38AjVHXxva1PAkEhul1v1vVvmarUwFap4KufnsWXZ+5lhiC7PR55OvLJZVHcNayb2FmtB
0nTtmnWkvAntc48LMgfx7KnE0qPjQf0X2QHXPYXZbTMAXt5H5p/8BrQuNm0OXh8DjzN56oLVH+do
7EJfgvRuGpsMRRYrEr8n3IfTcFvAq/I4YsX9opdPY8BrvpK1Fz9Qqrl9NkBxshkptLW8YiquJR4U
e8x1PObkN1hXfaD0mIv5izJJufJP+vUqgUaqDgPCqB153Dn7GJtyUF6h/2ouV5e7ymTa6umE1fKx
OgSIJBYsRwYPP+9HUrMjhv+uIX5KGLZSQ3Ok7N1f+1zohoqKJ8YQx3RA7wPPxWsr5ZlGtQa5snSa
8bXM34d/ArC4wjvrHV8wUokpENte7R46CIq5MGXGzTPkVrXjN4BIfzKv0zl0+ICs/HL3EVKuNw1W
w8dLrOTA4qHxTx+dZfpuFponaiBbcBRMCAR19ueu/uZ3YBy5tMhvTOVNyXKxvE8hKGjRFrVl/vBs
x/oT496S7yoz3Ue8Ta5GBvn8DiSEQoQBcb6sNNF66s/0hgzJgaZZXLzSupoDW4rvO3VeHohb9HV1
3VMxLVcFi+TjCMQxbZe9kno44Zbdco1MtImKtoMyPiaNRBEzek3+PmHOdcluRQPvBdVh+PnML/+z
XHhlBOTFI50hD2i6QQZcwSW2e5p6cdDzYxk7qNT35/E6lisL74YEoHJRi99+/8bsHp4IGaU3BTFP
ZNVwfruw0KwCRowswh1AcEO0xqj8pz+SktDA5LkOosF98E71l76+MuW0m7GIuk69iJ1unoN48yzk
bS26rfV/y2I+oQlXUoev40dlwMV0/Fq6Okr/9CB8IOnhYrvjkJGxmnMufS+ZlswGFotPZJs5FAKL
mVCcKsfJqPovACOdRCRORpV6EM75wUIE64o5f+HG7U1l6exNqPG93SIMYcCl7Q6I/HuJXIuVQ0OI
U62478ASqnDZV/2wvs5lU5di+UtYAdi4nWaB1HMRdCXBU6YumGmHMUH4Z53RUEtlcXSRVPyg238R
m0rYg3M8tOoXnPXPWY7bZekSoBRhpLsKH4E7LjqUAFxegAqfggR7B7folCUhz7C+ZagtXLi/xjL3
7pIsNiSPu8Cao8iyuDOtAMAJVEX0m4/dfqTA8NOZxBqe8AaJwxPeyd6VC2BNPpze/C+XK5di6IPf
COcBd/bs6SjkgULR8R6QHs6kDTkqcAQKVFK9DG/Ic6/zTaoNWxWyRVoAfYb/RNSGaJTxK/jAPtQG
9blNBqNI0T8osLhTT28jz7VBtpHF29pjFq/hnrqfQUhi/UGQhGXyjQ3/u/5ok9eW3WRGTYdVA0SQ
WhwLLQzaUDloUm1v6o35jyzics1n1Xm2cd4LD6in8XDT/RmHnJirYCrxo7gBFBOuc4fq6XvMEUHj
JnrLOvWjLQn6gYPI4UjWUwO/5pLFfRRq6Xbwv8KAm7GbCvrqFojsaBWDpv5C343JxqBFuB5otd/k
r7aaGA3hupAGnoQAVKoj/gUTpjDZtK7inUiXtohy/adm+Xd4lLCxDszF5SLXb8lOsJouHVfdqQWS
hOGb1mpa++jUmYHNyyP3JM/jM+C1iDc+c8UzHSFIfIK/qQPFM25U+lmqqCVP3LyiVB0VSSPSevy8
zQrnh0i7Lyi3Zyq08zFE6m6TSPi8UveUCREOGPeYEU1STbiB39yBXz9NSpySWRuiiwR//nrcCVux
k+0/WWvzajtVeWl2aZGAc6UXV3lBgdJqBtcc7Bz8Gq1Q3Zylnm2ef24jlLeRuVqyKiyAgHo/0a30
uEEzGgxVwlHGahA1zsX+sYcFIisErwg7RaeU0K0RewyLrEXGRXQqGbSa0aMOh9jSpd9DhAvqPSJs
CKKcv8mAbQk3vde3IRLfo3Jd0Be9GAlVKI6dB6KviTSZMFyGZfWFc6I14IQz+maxF0UBgEEv/jzh
VeigFWwqBnjdTVuAoN1i9DQASXWs0wHtx2VRBJ51dDXzjcQKubyPALzVPD8BI106mVs17VCO+L6A
l5r+Z/smghYXqdCciP+cUbP2z4QT8HN+d6YsfInKytDUeqExXilDfSwJhtzGrXszs6SKcr/pRDev
mm//2g+WVy+JfvJcK3VLrDisecFviBFc+dHRSqPkSfkOLws6+sj6emzAWtnowJkUoNylTYw7jMw9
T3qppXqok3iCSsHgUPEX81f+uuwHDBb1p3/RNMC53QO5j3wuUiwYj1W+r6+ehRRU4toE+X1ZASqu
uhl7L40OZsdfUk4iBMQkHVDSt/VKxHN+Gp9UwKopPWN6wZpTa8PbF0Rv8SKV3FEUNMfbhsczGN7L
qqMssZZGTtCDbJHetWNDkplvMt7ql9h57OoXstf2QGaf+Un/dK7ikFHc4FiQ3Tcuy8WQ5UDmYTKw
cvZXemUG0MLB++bA0vFUUtD4dobmWm2SP+op7T4AkVzYiim+MPgXYQnaD27/SmasOEMgB7rFUQS5
E2wgUKffeueXUz7LpcKO9h+24Jc7mt83JULcLuxhY43BnBgcjgP/zxl0pXbWY5rfSK4mujqtm3Qn
CKknCcsCgt1a5VjYLZWLTRhPqWGIoF6K0M647m1UeM4EYbRcqibyleie/V/fnTDmmeucHaB4Oawr
EHRsWeDT1bNEF3LOct4X2Dl/HJU9EI9UPZtI+0i1SoQqDHb0oPcYSqGA1LJgBwXbC/Ys3siptbbN
vduH9+sbhCnvvgkQ9Vc72SS7i/Rmm3N8Cj7HQbAOB7RBrv3Zj9viTOwJdIPAPEPRWx2vCBndS9/3
WmAvFj6dw6dqx+FIbYI7rXycx8iRiXt76pEPbhWaqAq4JTmN1qfD3pjNUxw5LSHdH9Cd9ZslyCpH
CTq9i/IF7FXt6krdKNDP4pdCb00iJo6wHW9maT4Dzo78YfuvNI/M4Dt1DNNg7cIall5HzOrj8zBr
WfSeB0SAfD1Uoi7FvaoNrwDUGBECKORGxjMxW5BLHM+K044/MqPukUOa/jtqmKiOguat6Z6GVXhI
PR7o4v4dbmiAoF2QSEa3Z6NCZXhYnBmA8Fd0J/IeAKhx8XCwe8SQkolDP2kVmnXvgvSCp3S13A44
/GXLNGXvV9sSwn0xe1176a2lGvDueGJK/j9gvuP7CYt8zLfuHw4oSSHVQg8SjFexuA/IsriID7Pi
c5si+KE4chqYw8/sqgphDaljD5iZOy42tkzVJs6cVr87lLBjEqj+7Y4B7CewlLuJyceKR1qj7JzA
jd+CNhZDdmsNEyc7ed5yDBBx3NYTgE14MCMTpaOYPLdhwDWV8aktP9Ml4c+rVqO5elhzpOWzU0hD
TnE5PXwymEIGtFhI+8HPzTNGoBwELDDGCQBBvzEBxBsVOdbfxAwmertZV58fpMgS4Zie+XilcN3E
QPYiT2bq4F2xkHCANpHNF6tt6lfUffowXf4qCqHwoCA7jtjt1D5niutQCBMtRB/McW9u3aHogfUi
SoIRDCLzuQgvdAeDsJ5WKYOURWCuimnp8GzZkUNymXVDaz9jfz55AVocJC7vlYYyvPMw8gIom4WP
zhOkYHwlZfx3i6HhlOrv1a3cySI5MdSBA/UuRVXiz5utcLbgp2MoJAYtsqOoa23LN8NIfTtxb2pS
JeKsZItJryGmkSKnKCqTgldeMclGAp3c9SOHl7qbSgzqljLjFn3WoPuLK8MuSQVn9c/GPCwC698J
hp+Yjn58iFrHReF9yeZGeWmf90ahFTKx6R+n+hVqzPcsmhVRVA7+CxcYtVH+o51XQlfFtaImXmpQ
MLKj7YH/xPwUllKZKIGRBahY+dNz+YE2h1BYvnYtxmJsOYhr/zZqEV2urO68FFPfIivQf+AouV2B
2f9R8xHn4P8O83eMXEFASC8wiiQPTy3nstK8pRJyUI9x3ItTE31wQRuEI1cY91MTjKTF1gi8c4uy
Sy7J2kPBmeLMkTeQj0Xqm3P2rFfTG9L/MrvFKfxNzbDlPJXqI37tLuiJH3K3iXGrxeuw3koD4vly
inA6263mcp8ssKdcVQvssDSMxr95Vbn1Uh0aAFs+SWaHlzyBDsPqQVe0LETSKLeWpoXNlfWkmYhj
ishZpkuHIsl39S3B6HXzcfiaAGy2DCXlpOs6LdZVE91jKh9z1MCM9Fw6h+RCMU60KYTL3zWtw5dg
2NcXqGIWBwGBBJ3ErSrJFtPZ8AFBYichhd6Mfxu+xiajNxuOjha3xcCGh7jjDyjypg6ckwLvDnkk
vc9I1p847xWnb+y3pmNbTpImYyqHh19e5zfrQTQUHtz/dtv1jnyQm3xbmJIeJlZUWJ31e0ZxT44T
80p5FwJHr11QbepFEcWDAO0BIXtMnbiJ+FXUIUSrwjhKFMRZxO0mkpolZ7eZEDD3NVlXLEQ5mNqZ
E5MYTFwDU2fTEYGX52auadHqQnhAriBGFY+aZ3oo5HnTII4L82UlZ+shG79xitQ5vP3PdgU0l37h
eipAxIOuH378kkT12z3W4vYnQSUI9Vz41UO6woSo1HzJs7WMoAiA5EXgu+mDBLcft0sLxtwZC0vc
HzIHrO1khgdMVcFiTr/QvvaT8KsaRHEuzRe8nzcJMnQPilE+bfrmYr5GQC3GONDTz+xcxYnOEaFs
qcBaWKOeERp5NeUNYVHOxnTMA0njzT5R+feP7DLYY8SdlIXV0qvMpSs21vXeKm6IrOYqUnyp6lGQ
dt2W1pg1xv4q8wdjgLWbSC4nxnDsfPq3KBY/U5VT2eahTyF5U8XsB+gv+3SWa9xkgQpsKgDW4GX0
orLm6oWPLujveaA483HqT8IbTvBcmlbSIptqslbLV51fP1xHaXsCjo8GQYe/NyOznnjHPfBP5XSk
kfk9qokgUlNJanG0UHSX63zIqNBXBB3IWpOcGV/E6U/o5VxUbKItTEBRdoIL9jBcX6v5RD2bc1RG
2Y0cpjpdo6JxsGsF5W2aATeQEvmR8Y7rUpS77wYCsE0PPOM/x1yyEE3cz8KX8UdJqRUBIpAgl/FG
EiGBrKXdlglie6007mKiN+epa2MB1aToRzIt1DcMgAD9rMHbbYNg80OUQLmCqwmgbwV0WhU8K05U
yN3K6idDEzwrZEwsjp5nTHSPNqgu7nwkeVpEfqC7Y02NVwg+mn2qiL26iwot+yyOYNSvQ4EjY/6F
GElRxzWo/vG29PcpzLej8365D8IVfrHwLUMBc5XMx5aExdbvPrHpDO32oxVcuU0gjvv1kVi9/UZG
twheRk8STOU5plfwg/LC/EGb5MwtnXP3oCdHnou08JWftegSScg47OyQZa0nLZTyGyNL38qvmqG+
rV4p7FSwayyKUj5LuKj2Ikg3HjxWi78Efg+F3cz9DSeVOVABY+d9L0WAqXjNadv6G+tlsVIqUYg4
xnQ5pUozGPLwwMhdEepjEbqJekSql+hk5SEjm+nqIb1kK8MauQbOcV1WrfGqMUxtYHYP6D7dmHJ2
7XKduzcodDeJcfld2M/x39IpMEUlX1Zk9MT7+qQic8vxUX7HIYknv/GzwNF0eti2h2HLOCXi2Sit
QQuf2DjuqPTRNAowz7tpMXzSV7mqJ/olarYYpQXEVOm2ZPAQgl9lR2pkgICmfN2f7Dxe0cMZ/QAz
9N5EW1DawkTsnwhSZyxWYKVm1GROIl6/+XzRf8Xp8mxSfbNACCSwKDXzViQnzo35RvB2t0mZnmdL
sJ6FHi9calmlZj8E1PIUJtEb3liB0ER5vxWEqBpyVMoUt45LIgNCv287CQTsWStHja5leUlXsB6e
xNiJU7tRboEhWfCWj9NVgDOTW5MWE5Xpl5UqYqIkSWRzJcewnV66wulDZlCyKknzBZxOpD4bOI83
s1sWBSKypBNcdjYZU0ELP6lTt1ke8bDGdxed5dtQoVnPMQGHOnFiYkaLsHaMcDo42ihT1aXhELLI
+6zp3goR5PSfVo1wyY5gsJMLpgYrPig/MvDV1lPkPekr60UgM7tK2hR4jlneOeRndwrhFjXX8AR9
Yq7SK+/iPVGy9Dg7KmxOhotX2sHZsJ9Whk4bm44E1jWS7u9x48cXN3Gk/wTQZFgcvL/Vnvgah9VP
HSPoFPdQ9I8i9E29fiCbzt3JYBXHoPBQMzlQLnmXANdZCwBOr2LBfX9DCVGTINw4IvYO9NiwGzeH
Zjn7JGxMlhFC1bgLvtCnYi+ITL5ij6Z8hqyUsJ0a70D3uJ9tpgvwyrwad6cYq0wRgwHoUl7IpHC6
nlR3lW0MCT7gpOw96m0yWnytO/COQSGzoTkUSy5nG0sjZdQ9rQvlzQ4O5/lkNWEcXubwvmhkVwq9
vliD710hFhGuocyaAmAQGJ3bssQQ0+upKqJMwlwTuFBshnfF03qJ5l5GB+LPA3/w176eGnt/RDv+
yDpfq8O6cfPHuZWXYHbUT1Jgvb2NxUKfca7YZmXilhnNuyGTMUYlNFL5VRup/Bnlcy5zbW28w11l
l96+ZjFRHI3W/lTyMkPnjZNke5HQiOw8d9qE/B1G9e/j8FpusCQO9XR9/Hvwv+pyDqJRr4TOcGSo
CCNcRbutNxKvgXLAHV3EAPj14g3YWZUGIjrsGSHk8kPYnOuf3JBu1jwa+WV/tP2QEsiq4vX+LYnE
sVHHl/i/4Lj0ttyqf0iarJeDk1sGmRF9zngnWY42uom72s0mmVtswI17TEZip5tpB7Gte3h0vkCq
8NZUX5cbVIOVm8VErZMdelIUcz6R5SSaVB3CqFhsprCxlU9OfqtcMv89XObOfS/cetqzbmg1AkBP
AjCLFLFIdORbWmk9HPbfjxGBVp/Ng89rwydomDOKqcBkveUWnpyI7AMfaXdCbz9Trcbudztfd0Pk
knefFlKk/2xZT0VzHSplpK+YU78oST75UB/C4GYJIMJc3H49VLnfeZz+QaBVE5Xw+I0aDxQDdxin
iQdWaaRyBt4ljc78n0E2okOpTtMszFJvECbLjeuTKYqQCRz/UroJra/+2twSKSrc8gdS942NcS5t
ZOvsrqrusxp1mtpA1eCm9/DXZtdjKLFa1aLVNkvrRFwRKmwCaKNgr8V1Hxc45pIbZNQXi0RLaVG9
66yByRagCBbRUNZ+1vdAJgZKamh3Freb1nodKlYvhDZTZnuRkzDms21srWWR+2NOZk2/NPlWk1Ab
ax5HcVD6+OACU4fFOk5lBWyiaxiY2qTnq1RSps+gGlV3Goba9gYYImEbyaYZc31c45Ky5JKN9BiK
iPw5xK7iriNoswfzkPa6ipWZBfenlTmMSxdDmDzj++n9M51PHjhHTp8tquPw1p33KdUXy8QWvanr
4o74INKzR9dKJNdanYL9tUgp8GD9Xm2PBMnLbJ3mdijKJ7kfR58C4w758DpFKDaFIM1q5ZLvYRuC
Bs37sL/r766FnxBumw/FJ2/FL0whDZnoIOvfRx7JBub6GtcOVtJULsrGZYERg7+WDRqfdD2BIiZH
ZnSE8fO34upKnq0twkkfETaWU8+C8kpgRdRQuvzbrBUC5MoqDQryIZDkNcmz0q+sjA2d2qKITz9z
A+8i7nWL4uHfPg/2Wk1k3vM1T2sn23yvzNvf2cLgZxsOzu4fPEFerqRVrWFY0792wnLT0+sCBrxk
NlDWiB1i3Yt4dWc/Nxe/KibT6G7CG23bCKXNxk48gvoHb+ezcmoAew1UfPfsStjVG1v2K5hO1kV8
mZK5/BXNFdrACv+zYXJ7Tnq3yQ3ZgvmQrCB0b2xGraTt4NFvELyXaLBjIIYECLGExtZHl576DGPV
P3teYtZ0Ph0JN1dIUmzoheIIUKL3Br5HC9gibWIXkLQc7etU5cuMsL0bOKmLlVX/I6P9pADCAdq2
XEzQVzZtz0LKFq4PnltHPiCBRshPPeDUiBzUH0YeroZt2HgpwArdevGdWc6z9fTblUlq9FexADrM
5cpwU9Ha+zTPUtQYi3XfLc0vI7FmR9bz2RO6RprsxhZigrX/nLTAFxwL1+dzPKdpbsSpjDlk++IQ
q/6chJOiBTr7o8B9k5GnP0V0NDijH7ELZCvoHrDEeq+u+MQLHCNNZI6DhBLV2Y85eMnwLz6p5FDP
ENqzwV22ERGrvvcb3xLcuTgpniLAO+H00PIuIsetHXAirY6r59xF/8mxyQLOTp7ytjXVbYZGEOvr
Efd7tXUqOmkZmlhOr3ue7vH/IedTWL6W1ubfNQAKeBiyUuwXOsan3TVr/1/eqNaYisjVbq7lVxnD
yf/94P0S9d4O6f9CDiC84M8aKqY/fNrsV2DE1X/j5KToAB7Gzj/FoyRjdsa31f33ti9lBEcYMqHe
B4fJOsVm9YTYMTSCZ4BblbP3ilYAl9LeW/5Z727GtCbKLY8tSeOf7iGzu+5b7QHVcObnyBbxhMPG
E0N2XfKRJ5F21W4oOMVw5DjRn0QrlvZzPy/scr7l2y3eaIhKjhidAeIBRmXs0uO/hJyk0EYEjN5Z
aTI6ezx0mNLIlq59L+OJtJdHtCimKgOdbCAoSHBwm2NYdNgpgR5Wb8o1UF0Z10kIXCs4p2nM+PT2
x5HZoTZNdgyyoM5FJ5PzAX05GMnKhcU6Nez/qz6MOaY3GHhx9UYgzKngAX6m3d97mHOVpZHX5Cyi
+6UJcmmq1wQCrt/Y4xm6PNSeH9ANnERzTSabntfT04RTa49WwvexrwY7CRtEtZziiN9TJbIetvbn
my+0x2IYeEZvcF7ckoP/ou7uYAv+t6EEjM1srIHANEn4eET17cYnziMJdnr2K7VaOeWlVjv8XHx3
LiTJ74UZVUhenWg49LPs6tamPSEoVE9I/f/90mEEoJjW/02skHKL9302ont6qrmxlM33vjjoATDQ
GHBL6+i/kSHIBT9+bx9t+8nOiEPwELMFnxxi5NxqZYVmMECY0334DYuiAICKv2Fu1XXGnPsVvs/Y
VIenT8LMTrEz2Sj83VsNkgpUDVpwPm4RMhRzeQmiWQ70xhOq+FUos322+aUd1k2GPBbicrHsmSu4
dWV1NpxEbgzcCT2mV5n136juEXjVn0HFENqcNFdf6kts9OuGsijBKKxQakhGAnxRXCp2H984usma
qCWn53swkdMa/qKihD0qsJiV3Sh5/WfkjCEzlM30wmVxhKYw2EVpSEuL3DUL10nSiOy98/7IcP0n
loDfogBlPriwoCoKKZQo5EsRMKVtwaRrIaM9AOqYsTdEPZv2s8XJr+XewCbltf3rip10srvfBl6Z
V/eUwUr1BwQaGKbZv7dXbDbvtF+EPXjDUe/PL/3nP8TmO3pJ2ySM4fowqNX5m859VDaIfL+IoBvi
UYT171cmNePRubbrThqv+/alMeDvv58f92StCFnZaM0RCxDGyUio07Kea8lQPY+JCaACE6Z9O+8o
78eDU4zLakdrAJAFFCkyS640V/gxk8cemeibwJm9CQDSbTfgKZ2OzpejhHFBjDwd98kp666zVEyO
Kgzd+c+J/La6oqPAwPb5khFs5j5f+UIcpw7XaMBSarrN+68Tp5NgAlRF9kmcHWXlZpR+0gTeYyfg
8vlOkW5wTGN2f5WcYbxpClYPhKT/1Y6fMAjwaiZAdWJH8aPCV9xS8QW4nRR4njdlcjRAXn08LThk
sRdb44mk5bwySAMEhSZezYgEwTy4YmNOuj1FlquVNyQAYLkT8iN1MrZGfywUsdCTZaUEQrpRZeBa
XHr5oRScT2qhY3hri/k7M3iBT2jQHgQbVckOleuIgaZt8bEEj2j6FLPQfewUfKHH1j4iz/uvNC2Y
1468EbOM+IoK0LKFJxKzU8iRq8WhUcVsIOba1rPbxv4HjUwh0HU8nhOiVJUWPh5bPz9zNOg8NjXG
6n3kpPy1QnRP3NmTb3J73iU1SKciQI6YrbUCGEDPjsN8dvnpgPbAd6r61HJOJkzkazOGGD+ejFSE
nvtOzTmjj4gOtcsuBs2XaMk/0XXrcLN7DheuNcciglBUhHpvdStA9sKdgufG9ix0feAiGNQyX/MG
9nGcN7LfmPgM3KzvTQO1NWrqPBdvgCR829zP6loeqIoUMhBsxJMOqM18DNoiDvGxFRxjQKs94mTU
5cLn646GiXnOiZdSkpgq38rx8qCwu39R1ac5m9K0N6lAu+4wskU0elK31LjUsskM3mYOZzjDQScQ
OOzmATVg3ULjHpiw4vALe+RTGZLAHxdCphaquoyuxvGfcGh19tkrpjhYHSOFUZaAU0rc4Pnn9PGv
giylUG3z5zEkU3yAE3vhCvSvITu9PUd54aATB0ADtIA5SahelaIR5MzJp4FYCm3pidHqKGe5W82r
0+2WNxZHPHDckC20b4TJBRkETNQBNiGui6sOpFcyXBP80E7IpnEbGWpCntf3o7KpygKpoXkKgyhG
LwvniW2kySJnx2+ONaESug8OT0y4q033YGkIdUxMN5ToYPYt4PCFhCtn2T39YNh8Ic7d9uChwvWY
5gdMgnjZdj4M2bBQ3UAM3gN2MZLPet1DXy36MIskOOwutFSVyBlUDr9ug5btw4i0PQp+pwAqfb/K
31ppk8tkp7vFiIQM1HD5tEyh1To9CN0G76vNbEP7DiShHRLMxJTKyb7kkYCaRYaPg6+qbQauL1JQ
W2sgUMbZr+y/vV3GQHfkYjDPnoz2uywduy2uDX7knvzn/hKcAJA9BWzthOaYYYeQ+eJgxeFunCr/
lREtIMk2yvbx7bOYKqroCPHSm7lttfXHwXNgXIfTlNO+i2NRycvwU3Lb3ycsTRZlS5mnup1IoQ/7
TefvijXjHPwn3Wet+MN0b3QhEJoYYOOATiIf8zlUb13ULHLSqaBugkBfItHbZlF+vwbOfAAvEZrw
PrblETW//Ga2WQN9BLFkbd0cc22poH0nEUDovdbA8hVciBlucyWJPSjwQaSeSKmmRDNJOhTmeUNz
OzAjC4AqefuU9JsuZq7bkNH+ofg7YzDxMHUXNIZ7oKKXxA+w/4+iu17K7Z9KZi0gJEoXljpeh3b7
8U7vyUnL5zZ5+HW6QvG5OdafYfRYaBNqcE47C+Frjkq4i2Es+D/ovsWs9tPwi12ogoDONKcjoT7g
YsM9FKZ6dRVHQXlyn0GaKnMrcCI3Sz/LF82BLanF8LCTJo8rT5zuNjqIG4jldLizbiGZUdRY/DE9
PwKHeDP/dtKSwCqgBCA1sy/QsAf8af7Vg8kFWMKhU5/X/I1aHpd+eBoCXabSid2Ta1ZjFEEfnMKg
Suo/+x+y2EdZUJ/7NWJTcfOu/DCJssFP7MCn+RUQi1tGkcT+nTSkST1ndlrmFMKxTYk5R1Eu7uzt
mTtn12KzlH+x8JL67beJBOrnKpEHof414aYU+LswncX43cMxuRN3Rw7SyM1iw0yF+fvmLAyB/Hlh
IQuZWB2gja/qjqQl+O/qVFMY4c9SV/t/45A60Tj6Vlyoqgg7PFqhndAD8XkCcTJ0FXskvnia9zVM
gxSCFTAKL1QRhN69gw4SHp0Cmv/lVZ3boUQSKRl+PLm/h+6NynvGMXYQAr2kMIpJ9sdnSf+gmzvi
ptV742cdcUa01Uj6HTEzbODEMLOuv06pGxt0ekeCAHnXY7VMtRGNq7gnkpKxWv6CGjdUYyPjEJyt
bYKU5Nx9b+kWGIS95zR6vDw0UwAtdbZ9rp+oDdaxAVMHTnAyR4DFs63Kvr71InaeUy8ejmMigNdZ
6w7LA2m6UcAV1ln/Eq2/Su+QN39NeCu0dE8QOKcdU+Jz9GQ3AbaFOFMSPGgsY6zpsDGAxuNRgCi1
7P650vx2wwhR5/A0eUB7olORAeVjJd4T4wNmnmoWc5UobDLgqqCifwvLgZibfoo7e5ESTb7VMp9f
Dq+4xgnqOFYxX8hebb1WJqsLL3SpMDzufwuU+EkZ8CS0/EnpAyLJ7Er4ljx8PyEnCkJqdPcrLogc
GTO+QCTkhUuiGLOyqkaGvA2BNyulp3YazTp1pYzw1bVHUCn+nqk8Abi0WCPcHbQ+uPjR0YzXz5kL
BXHSWciSxY3EKjBXe1gJYejsjyyJU2+OGAGIss0hsvLi5sW94MY9RkBjTiVVqQBaIVZz6Wbk0Ir3
FeKKyKBGDOad9pcCw2E0jMCt0lQDNsu3h/yVst6CHcSAtS2asFj12eDY6ReJScEgshf+CqVe0/Xd
Gedl1LAKTKfsj9D9s1yWmHxBKS4raRbFYIFcIPQAsVSs22q8V3QaK3x2va9NBESzVF7wOZVjmeed
wPNV9NhYYFmUwtU9fLDEHFg/LTlqczfZ8vJRmu1knP25YqJRP8CBO1ajRU5jk8U16YX7CaTstsKP
w1BuP1uewzEOMotlGG/hm4Rrdr/OmCw3bh+sTP9LwUcMrNwLiMpVsuBkESYeUjd33k8VwxHBjEXn
+Pf+auhSBiWLpoC9h+ExlmLee5W39AQvo/raVjfp88Pg9iTyXxA4ijsDBL4y6fZVHhXoPPvHs5Ic
5JiaDCqIjhVuidKYy4abTb1pS/57ZU5HcYA+zqcjEWZxzDZYPxP+SLbR0x6KB5f9iRFykR+HK/za
LU+VwnyyvlkY2CWiaW6aQTDkHAu2kXgVQ6cdSSQ8866oCZ7eRHfcXhlSkLAguRgHy/9YEFhRs5VS
uDF6YQalin0A2XjWJtQ+WU2szfGiQkpE+k26X8eD/Lb/7/xp9np+tsXk+b7TXjelRHZQhijWxStE
e3+Yp4woMrt3GC7YtWj/3PsgO8iWFohYWpwZr3JMw2pFEpNn9zBpPbFt3zpQ2KIAKZeenCIxEiVt
+Szfn1Z6mqQQh4goKtp27haG0CMxuAWzjND6XPVbtowqqVG5MtO74RGqeYPskX0X79w04FQ8Y7O/
TQCsXlotggGo2NIVCkLqY+q8OCBqolfsVOvOHZKgdZIBhds1bvNA2z8AoTkBouLvAOprmejiGeP9
xA6vGWrncn40h2favqlporV4HTNFU/YMmiBKTe98Dk/8xgbw8b2DWv/oB/3uLj5Mk3uRJ1E9wRNO
by6EJw1mz4SM0MXZd519qkMD5op0ZrHyecEeb0SMsnpORddsNZxUkYxWUH5uyuJCx/MSCzBUKVOF
ohZX+7qwqRQvgTaAJIvfLpE2gdnkz2/LfMMcQrU1G3KbxYG3qt63oWWu0F8vCYaqIkOXsvrmZIcW
FC+Ar0mMhVlu/o+YYab3zpM2oJBsgTHa/rXrpOjiYtRsXPUCIRwsjE9/XWvQkhfV7HI7gwRC7/Zk
fLUtrtjeudThskQAlUIDau+X7APnwLXpqIsuUEbtgiE/pCQdafm134zrXksZom4oDiYBwJJW49lK
KfE99nDplrny3tVkUzORfGufR3Eq1nFTQsnHbP0FVRwQmaG6fP+pKAmgiqwEZvRQVFEIL8q5X4E0
/r3wUlgqOlSEHRkDIYVAYyBjJ4qL5VcCMTyvB3QeXUzAy6th6KwSXFvtVg6jxYGr8gRXSvevgeWx
E6B8hem3nBM6ATavWXfwDDqGzrZ23YuLdUvpp52AouPc3CM6SYYWRqCSVabZFs+ViWJcPNG7vf9O
rklZ8YE5XS/DGJ3yayQmIe9PBUpMVgA8eckhLlQu8I0BU2N5vppcKu0JFK1h9PGDqlIy1j5ZtTHo
HTUklSUZj+hAWJPpqVeBPLpVpPRIW3L1sfcN/DcRPRJSiOT9/CD82SsY7ZwaEyGEURSmXVLaiIfg
zO6m3UGJHOKbyZGilptuPWnc3dI16KZ1QCYjQ0r++oJ6iJ50A0B8nTEc5zKrCSjcCRLP60NERoYE
pK/sWdehDav9HXg8kwxnHYLklu7jCQG/fs/S3Gv5uP8yw9vcBiWINgzU0ImMEDghZZ0f+ZTDdLvc
yMv8vLaig0MzOKzr387x4xhEDCf4rYdMDlEh3AlOCQ4y9/VX6D+TdQ7GNAUuBqAzBzygxdU121xr
ZwPHPVQWtQ1Mz6j+9sY6TLc/L6jkTANNRDbmbpWJ+6ACupx+YBHHKv5gpS/fUgXm5cGfHpcPSE3T
uX6SSXDsF0dPWb/sFcGKUjGXgf8gM34vS4muQ+Nwfqnj177O9BwShtejFWLbDqd1tIFkS3oL4NTJ
OMHtb3hshsNtRKkv8RZyNzyN/x1adZwP3nCMDhiIffXUjC+ftUMPGnJ38gApuXvRhiZt+lfj1rNs
TkmkxEWkTmZ7myD7g5hlqrfpf4v9MC68CsODwO/2nqJSc6yFKQBGBcZUDY5NvxqZvaa8Zv2R8+bD
/89XRlPZCYSfmCoeedNUOhLUlGZ2/P7kwVCwI8BmBbY6d2rTWtcvYuGotlu0+y6/4lUKBOHwM7RX
JGEd/v1+/bM2XkN9PRBvu2WNplx+/sOoYyUPrdbBILwly9sbDt+2WnmY9I2pZhIBDbPi769hcufZ
8gN922qRBmpjq5KntwaAzQ2cv8/+8cS3WDUVBPhbmyYQ1RVtmLD/5oF7y7AYiRAcLRdKTHOhz1qz
njV9MObxCnB+ourKVTo5ct2gk1DeeRtI7bD0/fzTvBAXnkwnsX9kR1kfN+8cGaxF00bNfX1OWYEV
vaISCQwKHMshBXtk4eBVibBLkNH7AfiWdoc5M4FvX9ZW6CJHivRAgVIAEAbRTGxb192wfJqVIjtc
f+6/hzgcQys9Hkg6Rl8V6fgu91Br4W5dB1NCRYfUiwlrD9yxx/FXoPzcbdjHSHJFKmkSqDP1vZ29
PWjjJ5GNXRrkX4iVAGmutcJT5dcEai74oq1PE5BIT5OToCQvpZQ88fC1SACFPW5Nha1Jj1L57VRP
Lc4jJbNj+OsJOh+WIOrkrVOvws0lzR7KuuKt7uY4auNIznbRieHZkjB03lSF5Ndapon3wEcAV4X1
HEmmyiXWeC0OGa2G9yrGLlnRDpRF8xEVJnrtHQhkKflGvXULwk0iN8W41dj/kXwLCZHCpvTn+3AD
0Tw17oVTe+JTvBb0MlYQUY1stMjpyNGbmsyySWDQhVoXKzv/w/uH9NcaEtbgTlsZ3r+Xxbvu4ziV
PWJr3XKv976PaIlpPViZl0OZ6+N29GtJA9dV/LwSXrN+YxSEi7R1ry6aX943u6Eokny/hffyicXr
jtQ16dklrYQOom+O+iKVPTEZTuCzHEa++bwlJ632upCWfWkpbcxEEAJun8KALVPnPoXLhXayqk7J
Gg1buro7r497nDU1/rwYMwy5qQpgYwhDyiehIDHfg+XGXO9uLlID2QTfuDfhK3/n8armUI6aEjYm
etdbP5BZfiaTQbf62PYFcyHAjPm8xNX9k3ZTTkTjNH/Q7hiB5vVGpYqQ0z+wOsl7YP1loW4v31j8
S5r+FV4LFhuyLhORR+qAjlkZYWiAw+qSHWb3FaCbbkAf5+9bzTRpeOWH6js9fFtcWJnk3uBtcUei
2oSh7lL7E65BKsX34uDsMy5g9ssxxrrJfLbwvH1tHzvRdURjYDf3J7uZByiVYGXASAPak2v+wFjv
Tj3Y7hn5GVuN+GJftX/lAneO1ZPhKRVg7Vh07FoIdlvb52yAyywBFHmvbwlsVDiuzGTi8w/hzdgk
0wtmMztjIdZQ706SlwkzKMEX3dYyrNTb121TFmzrJQn4B2S3K0P9McWPlQnnsQCT1IBjIfbyAPlH
81UJx2wbgHY0w9r4mW4MXDJREjWcxhT3Ld60SXFxlBUla6ZQYiEESVKyRSunZjzWgKq5u7xoGAIt
IObiYVUJLoid8mu1DUvHY8t5vQOUSMHEyJceck5dy1hgb6vkSECGXgPv5iLsG1RRZO4O6jGGiDuK
k0rJMDd4KM0gld1LismPn6+Xajt6JPgYkbTyNzxlfaPz8hVUJ51Bq0e0IcmNzhrvkbytTbyYOar+
OMk+HSWISbZ+p3SWkVTYeA1Iawwv0ELfNnnBizw3ZmEboCD3T1YUknik/M/JyH/DYYgYYM0JrYXn
HoQrRJWqxiNTZpaBGc3BjmcgjjpffgC1AKhVqX05SPKy88VTmfDCw9taIedElOFtKjEKS7TnqcC1
ZlSa4Nmi/0d/L5LnuLEHcmlAV59vxfuL5RDYNQZgEeeUyBSVjq0MmCemnrmAjjVQ0JF3ktFYQrHj
JWA6wQSf2BQOOctSJ/BsyVKlm/tRNf97OopqXNh1kY9vK+zAFACvcSVJFZVQGVKiI1npDjud+f9l
ZV775N17C9D5QRKJxvKdr5UpzilTOYo9kRn14DqV4dDSGZzMYj/VkFBh3kUssYmKFNme7HdDx14M
Rc+rwsDLnZzUt5VJAFLB2hRo956GML4nYijmPzd5j9CtgHHikyL5JldlbmloLcG5BZp8IaQAnlsO
2si1kQ+2zpVPytizQCOGmmHDLO9QrzbfRUID2jXJG6ZqpZTf7WNvo3bv+7GVDhGSGtkRCrIrvN0/
Zr8PqhlwtScZAwHTClzquiSxINnQMLZDBhE5XgpH2ZMC/KGQ9TrteuqmK/dgVi8UY8eGpm24j1iS
b3VHPcnJ/sZbihbzD1b/rzf7yN974i7UxZhQoo7O8nGH92Vw13ybzglBusbgYm1kmkeJs1KFfQn4
QEli6FgN8Wst/SYGwKmAaLpRfifjZQv0tyKYwXLULh5F/6CURRumK0MIPPQxJZ4v+O0tRIY+RHLl
+QyRRzulMIgapqr3hwkGMm9LOqmC/4WzLBPrg8LRBSCzTQYoMrDgGRacQ1D+VI/eLlfqvrsFDwnu
bgYvXrfYnaPb5URv3vSVgmzuF97iXJ01otPVJz9MC37jTGyl/hgRDtlHuL9aa//Ug4rTR0I4g44u
ed6Tx5Jez2hP0/BgSVdXH8SQsj+ZYHv5d5ZP5V+q08RTlwpJqc7N/VKzp+ptF0FOuPuTOqUost/Q
Binx1B/8J2I5OJ+hVzEZ0MV+kvavpV2r6+mlj6DkCv12HiWKbmrHsJxAR1uE1EpzW9g7tnHtWVl4
m3z8tgOTjg+etjn8VkbPRoH9deRorNP6GduLlSwWCrJ272tOj1klXPPNwl6yMA2jS5Ul+w7nwXCw
d+E1vMjOCPfyRdoA4FoqVNY7rDFylX+ffE7wM1oOJlW8JdSbjhmJwG5JDKRztSJ9Gmb2rYWnuxuX
2lCgMh42Ga9Rv1jpHG0DJIuqqLTq47E+1TFAw8zpul9NJwX48jxdjTjTAOXDDjNb6c/ThMbLDwhk
ikeJWuEmbIVfluekh7WLsiHQ2xddDreLYEOuFDoChzJBZ0E96c49M+sIRUcETsgil2J87/xotOzI
u/JB5WXOAWHzCw0u/1W2Q6dZZgi3C3/lMjpv6VZbxb42oyX3oGsqxTQ93xcSwxaRwR4XUt/4iZSS
OLj5mGESdvXCOiOmb57MJ9Ry9pxa/NRpdfFghlE/glnQ20blqeR+yJ4zKXPrSFoswfbKCqgm15U7
iFszGWJu4cNxd9AP1surInnD8OtgLGR0wswh/vCOUFnDtLL/YGjTf7YKUNUSMrG8VWjARF+lxaS4
grvIcEKTjPQ0PdGAxCsc+ipCOzJIT1X6ypDE5PNlD9+G7RxX1vVxYcr86ScaNxKCBrmYlBMUxYDI
y8+smJnj2f9Zf6Ghl4ky7B4sh3lyqr+lVq/olC24CwLpn7RK0Sxed8HJ9Lt5qV2LgJISXXkYJJ4A
eOViYzR26FgnSdCd/aIUeyhxmDZAV33Uu209uTuGo0ElXmqprYYLXMFG+TV3Q9SzMwYM2Ep8uV2K
dA12nOkyjMowWXVtFbnwNdkxfPLZHGoG/1luHpUi5BPFf/o/ZLa6zjICasCbQwSPZtOJoa7eRthd
nx249/TPizagJLLQgnF8v4LA+c2lAWDuLOcOsVUhbpZrJdGrt4Xcr5wwqrpuZszgGGbkVAc+b0W9
cd5weOSJjKN9D4vUTJ1OXUps1oV3i9vLq4eINXaFN1JsyrQ+STBu26/dPAqZt6MxN/STLXekdvDu
UtBfN2gKRB1KqqYLJaEDkuB8SgEXr1zOkh3NpRxIIoVB5XZ75NynuBhjhAtQnXPYHpcU/6qIxW7r
Z+UBh2On0D3LwWeicMsTAnTuTx7VBx4sjmbiJexocflWQotlpNUVFXXcjiU+ewd1j6MPXAS4zE6E
bBTP7h01YbSWZ0bb2trnkTYYWZaDSfsufiUKaREivWTzsQaJA9v/oi1VuMmC0xMxSrnS/U/auh6i
/l7FxypYiWygzEUoXspeoXMQUM8CPdBxJKhZ5n/6EPV7EsOGN3xww1pulEGklzZ9DI9PEv7BtaNo
rlyNc+jQHYcdr/qaCpqOkd9jVl5q8VdW5zj/C/k2rvhzjty1KdCL3sMovcVdv7uKaZWsnxi0suvf
oDUgoOEVr8syXsAiFpjOhaQd+1OH6IVEgO5h1gJquURY+vpRUsABF55tNTolmvH6sz+WC8U9tmDk
Aa7NOP1DaPFJTw4YzbenssyjOdx6vKidYv/ApaPqCi3PHp9hqBu5ASfQCu3nlcDJrgduAZWKTy4P
8QOOa8AA5RHDV7g3wA/4bWoc+pe85j+vBbdaDn8kJQUf2XaWQlSRN+L86GxkJAH4+DJLwlQ0PMxj
1pUpb3XG3QlSMwoVdeE+M2nqImA1eB7lAHe/l81FbCjAt4i7qTdHc/PIa5TCkjcb+LfCC5RnQwL9
igruNMWpUe9/mNTW9EY42OKu5k9/QUWV6mpX5VoYNv7fEsRICGy5kXMPbV1uMKJZBxq5mUgI92w1
8rmYKjIR+tLi6atxzU6ThCc6szeOYlZvX0uvzsibKbY1MXbMQVhEbqb5g46Z4fro1VJRAkIGwQZe
zSxsU6D5+lknMdPuMpngrID/35LCr3wZMYSFj04tsv4TChXcAoHM09tyV8mjvaArkS34ArI3Mir4
Ist1Pq/SE8fCAiJqot1rE5SA0XCX4I1EgZPC2J//5j1nJzb+JgrVrf4pe8WPJNdxs2Acxm+3QVwG
hKSca7Fk7IH1jkMXMiHpIItpJ+gJIgfhc26b3XWrnSIetzE/KtgSFvNVm4TUH1mEoRt5ueNR/5e4
4TqaA+kRV4bkUoSZIubZkbg5ea5a285R2c1Wfxfwe8DjyrsX+2Yk+oQmSKyHVWhNpYBiWKySiJGh
IOaCHemUGvemBi0qLOfIscB/VOLNl8x+MG15Wf5fSZ3VAqwYCmqi3ZYfPxNlBiUhXvhCzjvbePWC
e+aZP5TOYwsNlhiZVGd6Omc+XdzNyVfsVpWMFopSrlg6xWWNknbBRXW31+k+GaNvQWJEtfzUOlcY
1JDbjIhe4ruzLePPfXfC015B9iO16S164bKiKE58gUzzTIl+c5snh1xfamgsb8VfA/gsCWMv61cs
rtoUbp0stlWruR8dxHznaDS1MWw+sLfANDRO3KhtHtHTp7jLAbuc8Fp2iqaKFIzIqvweShquhid3
n9M2ecUAQ27s28YWmX1Qq69JHKo3x2vGhdMvseTzImo06btzEhnUy005B9He0cQ0/Q2+zK9ezwHw
VZ54GLvjM/62Ije3gFYNTD243+zddNeBLEBlM9k1u+KWf9tIdj4Iq6jM6F1KToxKZ1jWEV4JrIik
ZxsEnaRxlvlyhrwbqcYAfdqN89h+W4LLnmAZiE0uIglI4EOjfMKuVnRr0CQDPxLWWzAuu+ck3hCm
iOcNr4ynK7raV31Hn1kL+eYcbhSJoFy9qh/5Own6Qdl8Dws35aijOrZkaZYf1EmOAncsK4lV/5Gf
d0RmXIxad5LC9HnXI07LXdaFa3ltOQJHitnjHK1jzuwEhN3NrpyZOm2NhmsnzBJAMc0dPsc5wQVa
5Z9rvu3+0YAB7c5t/P5/V8bhNPPMauQ9kO3XX6Sju6dOoKqB13aTaO4ImOgLcTAN+IFX4298Bu2O
S3VswEB13Lqb/S4xy/P6FjZ/fVt8+KWY1yTeqTmxkK+NXL+CJBTtSTPOMQkdX5WKX//AeAe/hM/t
yk6kqqyoKfGt1yB7izjiak1tfC0GuEL/+th+J0PLA+JoM7XOmeQo4WmLA9RjTI5NchwgQe0njlt+
6ts9DihGoLonofy5tvfF0Tb4WXK4Zpjv9VAgC77aVpEp0TSNUQbhdK4FuEWU4Ujg7eeM1A3F5sb7
7K82aRDo8Xft6CGCssnKtfLX6Q/kOjuTw/rFS1IXnoH2GnB3ejInAWAR0+0T2lfpb5OPPOQpYqbl
iILBOpAm5O2QC4H2Ds5SNchqrPTpcupto8BlxM5FpoEU4pSQHpaeizE+DXjb7vTCOSZ7w38KObqO
1EJcbxbSpzp3roQ9TNtVSaR+nRpWmvph6IY+5ZW7T5/RWPwyYezO2whij+Y+GmCQnOOFlQyCcwad
FfD3l7F4SgiF4NS/Zbzhlm1bplUWhH+oiXTq91I3aOy399b+B5nyQtIjHTW00Cth4mPVOkgHmcbd
EUDsAy+F8sVrbHjYJOuud3Ene/dQzR/hpYIpBuS+sxLvPk4VTDPYWb195qSuc7eSTwHFTEwKdIkT
Fr7LE4YaMhda5boKlwHDRL10MfvY/lz59fd56M/diMRuxF2KTh4D0Onu/P7exYDNEgcRdnirIwij
XDRrmF2S05CSzRtGgzY1Zof7BPP0l3UfNn/1XD/3lwe9epmFhIh6KBa1IOS1tMVDiI4LnXx5CZdA
BxOlE1tBHYW1oyJmP+e9JbPUAElmFDF+Y9rUbY6v9Gdjq4r6XBWNFyT22O4JnnvoeIppfKTDjip0
Oo/Kjtzt9lvb+iuaidV3ro7ubIOWxXBjgEu7LlFuS2TX2b5sOZlzdKw4lBkPVnNcH8W+LhffoeEz
k2v84neQTlmrtbU92Dl5lUWcb95++9+K8ISGJB4U2t0ahkRD/NqTNwhjeL5hehcA5VTF+3pg1f5f
yFUHSwhlCCwjD5WEzFWzsBlq4mAvlGliicSIKCZGtczYmUEcshzlpM5E6iOviTzIIAMevFtBgbzQ
iBQNkZQ5Btg5CVjlMoUspvKnzSgXlXIHgijg/G5AVZSeK8Eq1ycZpwMMXiiwNJXTU/jaoZv12UmU
XBNsW5TDsrJ0TCMtw6kFbfjmZM9/K01BpD8YIUeqqTasi9B4OTi89gsf8CO5dpBvHohbKGnrYrhw
zsyeNUlFx7SktToYOUqTVW/rcJarCqSJjsepbBf0JWEzj+0B1No+k8PWZMvGZjw/md0ABLe8In8r
awDnUeap1LCOnnGuUx8lTgcXOTUrFgSgMDVfAiNfeCsZZKP64xPfrR9Tdazshbdcw3RXjA8r6SAs
3BFHtfVIP5eMBRqK3vEaxoK+NcKudjA4/xWv9ww8sQjYJTve0B/8mvRJ4+TrpWURfEr96H3HvP49
/sYzlE2QVqxBeFzbNAtq061naMcTGiLtzpW4ow/7Vf6De7NsGwd+FGAAUdosQXy1rW2ZEUuWr/ar
/IyY02roXiW1z8KZYHpCsGtbXV6MKYuvqsdwIjpT8PSRZWt3uvJkydUa6bxIXRYnx2dZo1ZXB7iq
3+HKogIWpjj2YmMLBRp3B7QibWtwcg6EVTCABYjz0spMDQNjHjN2Bf6ZUT2JarCWFKBXlQOXuU8Y
UGQfFACt+PgoBu2brH7RYFbsUueqkncPjGsjvAnFEbha/c6GUDePtk3dR9ISdFnGIZDuhpcXrU8k
WzQCKJzOwrtLS//UyE7zmiKkfykmocKszgKXwH5ZcbaDV5YUiun3Bhw61e2/ZVzjtpVkJUvbhgds
thX8r7TO028DWxDsl40B8IwelIDgw6H6FdVnTJxLnv6WC8MhttBxXsYBMxmdzIKV0aSYGRsJ+wTp
urtlr8CD8AqRLvUjWSl6HdGQHLI0X9xDU46majaKthZi0wzliPdKRhNBnZTGjKlywXDJGk8KsahR
lHRxZZeL0WWGA4C1xuNiNP/oH0tEawZfaZX8kZ6XCYKtj2V+4SbewL6XoGhV0QdCCVE7F7zKXkcm
Ko4pAZZGEomF3S71dfzmyJsnYPiA6uh6Dtfe9fRsUvyh50ZMj+m2Za+naZM42dzUB+rJAQO/8nAn
P03xAjPy4z4USM8Fk1BI5zoxA5Hb5j4hrIpCJeAEyiuPbFj/9MQP5tfE0AF6/LxcrMEdnTUON1Oc
79NO4MY7a/td73LvEQSQU5yfh1uCFQAzvFzC0CTQpb0wNW0XA/xFeNT/TKhi2Jm9PTGNPHHtK9hb
T2piX0gJGJhhvJGCktyXMTQkN7eFs4u9A8zIM4ErQs05ItdRPgs9vp+r7kkZRORC7ssKlbjlizxY
3mkGi2nSOWgkaE/S7FDPHzr/QSmBOo4LNmMObrs2Vnl8gDqDJBFPvFutQuUkjyK+xedk+MIqh3WX
M96N/1wvs7nbRoH4Z18ZRC49QzDjtm7IzXiqNrLZWO+5Xs9yY+D5Wo3lDbWCL5CIzwzsimWBLBNs
ZDtcRQcVXSGbcMrGVKG3JnID8gY+pK58Ok54Qe+e4SVn7Wvohd/CWvSGMl/0gZkFkUrnZcg96OAs
KYWLYDcjl8FKmJN85N0YtB+Onacqc08osG+MnKclxivNBqB5D7VNLwpIp9SRI5LaB49tYI+7KxwR
bl+viZV9OQmRbjKYhsxRRAuTK99sHZi0AaWBwIFiyLo9UMYMDZkEz67NiR1tbuEmPnJapIAQPnMe
s5HoEfbhp9RbecUXNNTb6aqjXwl/IIqpvZDQE0/B098g0STv+0h7sSJDkhATfuumHToC52XzrZW+
ls6WwafGkYBAwZOtlVJkJCTeLSIemPzlapP4h7byYfKatM1YVlQw0f75gJuKR9urvBVG7g/ige+2
HE53xPpetxT4uyrcVwVUANQYPbz9E5Q/7w2Sj+C1injPs45/dmmBGQCh67UyvjC7IAGVm9URrN48
IDsQj5AtXD54HRU/kU5MHrMixDd2aUPG/2gF6ddew4Os49px0mQKyHBtxekM4cceHNW3UugkXDKn
iyD4AmZS1rz/E6vMdq62U9Fb7Zyftzp0J5iIhgZkj6kwde/i65EYoeboVJjKhzZn43B9ZbpG5Q4o
Pwq2XteF6d2izVFByErvLR3MgbUOqj51yCOW6mToXVJv2wiSgFvW7enNWOGqAMBYTBDYbuCXNMw/
pRNo51zVY7ecVYz810MPyEVRQRla+hJDi4gQ+ircrXixOXE+wSX+56OEbsie3tVfD0omgHZZXXwW
H/g3gIMgge5Wg2AEjCjP2iBVwFOEhQu+Ysv7lVJI+PXEDl5rOSRC7EV4i3PtNtvtulqgVFMz/A9t
L5MXEESZNwoqa+nYSeWWlTTOjpoQbvdmDmkY1QqM5WJ0BFsOadvKEC24b3lbUsfF3wTiLN7kZuwf
oKY0wMTnEkaVkZu8Poe9n/NH+UgrWnIPnYybOPpCQl1W4+gEX942o9PhPXelY/cI/ZVGwSR+QYQu
l3ocGrLkAVt9gmZW0B3snKDfeAxpklLtfegaNPpMNOtmrCsnjF/PGnIPXlhOWdu/SvEavyBUcDCG
xc9EBQme095q0GZEo87UdkMthWH810eYJOPDqdbFmW3H6MkrCggAjqVmPwBkZ5XTlWH3ajERw3Qi
/rb2jElkvrB9RZkOs/v6vlQf7NDFN+vykuOP8Z7ruXpUv9YYjlEL4r4vGpqtZP/+9G9f9+cNWZPB
RddY+7KTc9dpHWrREVD0ED9V8IlMCBijlWWX651KJkFtZpWqCe/Z6sKlRUj0T7Hi9Ws+KfirvppE
NSCkyF/zr4e0tXGxMMLwketJHvVtFdE6ukNWWerKhJwP4MLoxr7AvdJYp1tWN/RWvcHcVB85CjDD
o1BtwOxZmjGf019eKNy7xtRKIOyBN/S6lAlX5SPCZ3b87ZhoHNiVFqslsBdE4f/w/TR/n0hviQ4k
8sRpXB65EfesR8nPeAblEKxGwLqHeQ3FOO7nR4McBnFOA8GqYdTplJcd+xq2bTJcxXGLqVdY+5Oc
bfc0Zvju0hEuAwyym+pk01Gt1gWTXBiWcUXUXm4ca2nk3v50XRco+mGX8MF6ezRwdkct2e4aMeSn
zItNmJqcl8mf9oDfBZvfahPqnE1Vh5mZi210g8Jil4H4jgoUv29gjFNKEuEkL8VRNMj9j+ItimRL
kqvIBzUbqGPHcqesijeUPAlv1p9WDFxkwLqAGSV8uxsUnEc/Ox0EoH7z0AxZb7aEwokBLLPgpi8/
OeoTZlT9hgcyfrEVXdGkEkT2W0SSSw1p71o2RnFYcxwDmfOAMOZCnzp3FBHzEi1iE6ctx4TaArxf
ejcPPh9/g0ewpflGaVhrQjhCP9fGBu7lOSVrmwdMX4nf3phhTeg76cBOMzAdqgqPa4L0HtR7/CLY
/CxB2jp8VhzyT3L6pT3PreWJwxdZgpzzjgF1YR687BNBWWyrUg0Kg1bZMikFlE3S2pU8QDnYxyzk
12P3f5vZOxXUTtU0DpD56IzjjPfh8jHCZHYuBWuOwh0HXbFj6s2qRGY6p5jeLp5pboOt3/4qDq31
3ghEAsu7hq8iuX9ddYkkBhExiWOFw4rsmhob9945+fgvuDAdd7sSJSgQ/dwPfbVt+3tQG8YvBLHu
1JEUZ54Y4b2gVyfRKmomP1NwYtir2iV+7xhLMNt5uc0fhWkl50yuknXGosTgTLG8jVDA+Q9ipqRj
c8lOcjJ/7EnQJscEPUmvy6U6bQajiFTk8gn5aeucNJ1AUdhFyx1PH1TsIuTUiW+5fCejlUfFzpwy
qJU8R/5YaLwqnEp/GjkL9vJzARKaoWeWp59YLz8zzuGevZoJFoBz+inGYU/AC23xqPG/bAe4aBdY
ZtrqV+o3CohN71U4ZLSq+ftm6iDXJm/87s4XDfZQp6w2b5CfvO0IAF8lfNMWnVEKF6DnCJp9CAOZ
H76ckXdp4R7kYoE4Wl+novTFfRx3EtIPGtrJD5z4HzGeqX/MrlWfHhHk229TFDI28RH7lhRBbBRr
q4v3e/X+I9tDp+dErx131k5Y6Wd0/lFcbtyl4zPunSL6TiiKsz595lQwpJtDKSkM5bAUuNVx0f5G
/PcgbpHdnq4JsjYlE3XtLzSlkuzZFM1aWUqaCc+K+ylLHsXzMHuBZ3furlKbQYWTHuNJ+3Cuy1Qk
P7L+2ycceT8gUIw8o9rafTXWYrYMA2NBxTs9RhoGYhRjiKjPHaHa+JZR4w8fUOVjq5wKx4JxyTPk
DfJr5hZfN/e/h5EH5coeqzTaiiLhqDVDn28UeuS2ZnBNUD2KMVeXJX9EIoHpAo8WmLp1W3ix0FLu
oQ7QWoqxQB/F9hCs/nG8CbiPcmr5w+ws5B4Pgg09l3iNJldTUG97NgW+E51se3874yw5uMux60dO
6pWF4Dd+Sy8HtFD1kZxqWXnRGEkT+e/lj8T3U8D9NedXuy0339WPTmQbnb2g1irHVigZ1GX7/Lf6
MZgSiGe43YBgv0mgsP6kfDboO7SQ0MMgGHXn92oT3TLCKTSPYSUXRn6kfxJGdH5vuqy1yZFO4FW5
ODsDWMyEjP7rssaf7oXiJRAcnMzd+040xjf226yYqs5nTmPoLAdwUntEPj/O1ZqVv+894+QzBPsQ
V1iolcTDA6Kz3QyKmiVYqizDEWQyChG73Cp1qoH0K3gzK2Bf3gIUWBArbyMzl16gzujFxJA4dkHJ
yNTOyJwoxyDtn200o+2cRXX3mApQ97L/F0t+wVltNsTLvM2Arr9tYg4A8Z/XtjcYr8KK7IIdy1EK
6iq0GmhNEWKa5f+u58rfnF1InBR0sJvkZyIspymIoc8YKPQHmWwdT+jVfeJ0Ur9/UXnzsflvfsCb
4NFmgSw+aHassNARQ24LLFxGfR+PgDPoJUgHoYvL7X9VLRywGgkPH1Lcf+E5V6ctCQXSWfKuj4+P
DV6ACwC+V6hQu6qJnTZB/5JnrKhvp0Ash4YR4Pi1U/go+molRWy5TSMsGJvk+XBJ3Qg+iCXd1e32
BRJZU+exzUf1rPT0Oa0rivNub4PgvW0fdyYCB4yMzpBAlRsZeFEC2hSWq79NjQPCu954KNQdN2zo
jqps7uU6dUMseJaqeKNAQ4dZqIooiMbM+6egRvxc1zhI+jJHl/q0yu5fMbfEYfTobPTk5FOgKfUK
58L5ErrpseuycRbPHJg7p+rUhYQSaSM9fGQByXsd2bDIV5h9fddRS9Vhs4pGYyzy3r6zuS7JcNnv
72rpJjTEwVSQVAzlPhPNHugn0uNBxJGr5Oir7CUeAzKS/hqKSbTaAcMuYsTZMJaeb/tKQBEcO5WF
TpPO3EOA6vLJt07xsmu4pvwWIJr/928l97TDSPISU8CFqnyXrzqgQiB0sqfgPZUoftQkaDFcoHIv
bpAV0wBQQVxHzgG1EkpHUYF86Gr8r2iSspsfdHwCCScAhKmvnkqSMjK3l5DOmREG8JoBrcQwE9N4
qQz+BxJg+5AhH6EIKtzkk+vJ2Mp/UAtG7HwpUlQTU2bPePfMW0cKUVVzZ5m/NONRoyufMdjhAJmw
0dwbGPnozfox5otxNkCOGP2AOAppP3DLI/n88qesFzs4xwjCs6cqjGRSIT/GHRZcsx9DKw7aplX4
wE2lWzZJoTMIwHEfCM5H3ujSO7oFazXCLmhFQ6DtUCmswKIlN292GCkEmaImGntK7ajsHjJxJXfk
OrFL4qLoRHGIVgwj1kU/QixHPnCJq1zoIhByjLtIvHn+yJ6f5iqn4Ob+wrDwUaCxDSc0PfB90RDE
95o/kiEV8aSgmEPM+rs8aighvJhe/XCoIZ0xlPnhPCRc8r6XcyEwJPNI/NW2SpsAGbXG3CfysWLP
t97qcHlA20kJt4AVcIuuDQsNNk7KfQ/SNmmxrQyBMlqzpLMQ8JPBYiNP2VsvZ6MXRg6TpDcOL2XX
B5QKcMgFIcqwaNiFY63/+S1Pc1dkOy1X/KSXdU06Kfdm4IW16FvalPC/NLZiE9i/B8i4fKNTv9i/
uCYx3kcDxnva2ZAh4nNpYz+Vd54LLAXA28jH80RsI+pMmMeeiln/3mbyLJCvDOtvBcj+Nqw2USRg
PXgectPFHE64kToNiGJbyA1pcQfm2qAoq7lWytHxNER1SlwReIh8oFi299STNwc5TSb/JcmZ/CNQ
Bas70/y2u2Lq4TvAsf91LKkyNmGi9X13kzS0tr7PfhPq7r/Ta3V55FuJ2oLAA6vNAaCpCLwfc1ox
b5WYuFA+QRhZazYtqWHk0vFu6wjMRO9xCIXiXbWloRn1YUaZF2hHNhyXAVB252UHjqCw0MBKAqIS
VXLvmlWMcoX3aDTcwlzui7vXYocASBa2LQmjopxUwWrs/jJIdRwZsrnTxOkiOghALvXg8e2aM6kj
BqgUXjHGiiwRboLdjucP+qYCBpTpEYe6Q2M2BS8Y5w+oegkLL9117hp/R8nTRtiCT3F97MS2QgG8
efB6VHRyvX9Nvtua8mxEwkLTLlFgoTAZJV62/4MMibY4LKGflhyvEiNg5/CV0oDGS9HF32k24AhZ
37WN5gnGpz8xG3bLey9rC1ZYfGY8cxSfU2yHGQT56BQP0ZgmGCv1xJc5tojJQDbkJ7GI4J9YpRlR
YNboe54iHO9p9g1MuIUwJ+fUnqTJ6+5O1D2FwaOFcQmP6bumpk9TZnIPnjq3d9WZrbgDLR6nnF6N
i470ZInayTl6KXW+95KAwjOECC1zg/Kx2WT9C3Wai1p4/+j+w3GNkyHd1VbmUJgC/6aQ0uZUnoh7
DOvi47TxX/6sOB+r3mw4xIiH119KeZY5y/d7bcYVnWhvbPeMnJCu7l4oU5LZjevas8eKIbii6vvO
Pj0zwV5MMFCc8+sEHuvNkOaUoh8Sp+XJSGlM6PYc4Lt1Gf6Ttxzbq7HWn25uCX7b+dErfl+4twJQ
/b4zi7R3CTuceq/LEkZPV3rWQuLp4ZAvfFnjqA/zJV9u7+5Hc9+D2RxvXbWjrmz2IPHGIokUnP6Q
013HNksNLGPRXX1YEChyfsRqOaPVhlvjXWZ9CFIezWgsNkkUxc8MDtxDSAKpjPUGQzsiV07s1lZR
KDtX8bedEX469bubckc/M8puEYUN7j36baF7VKqnBWDnZiOYg4iepVr9L1IllkzJAu3QRu5UeY4L
TXktCgB84hZu7847DK4npCuuQrl/7kIgmFDJImGSP2Tl3yFMtptiC3WNsIziKETZBj88zsDP0cVP
jaVFWJ8M7S5WWLy663dz+i4CW66WA3Jw5GY9P4DnBKOIH3ClUeUxfWnuNllJc4h8RJyTrASReEHo
a+7mZtQ76B3PgcEIgwjElkukapGyYGYPZo5oRK6G3zJhQ7rMUkGMg1JKRCeesFHKZMdmJuQDQqdV
PE2QYdWI+ffaE8b9GjajwFINF5OnBf8Zj5a2vtVO/1pIblzJblKW8c0Hm86cuIap/t6a79PIzGmr
6dhPIdPGBukHYANX3I4QNNSJYHyTTuXYc6xdkb+gJh/t6gY84/sTUDelVon4r0wXaZcH8mEPrRGz
GbfjtpZfoImS706Js2pBx0XYd+w6lLabpdjuyASGmohswPwR6c8PQBJRNw+R2w9L3kigiCB+oyAk
N7iO2GsAdF3gmBylM/DKLnxQJrOX0RbTjuXu1Es6jYL/aWjVj0pa9UBfUsuo/TJ3NBr8d2PDzoAt
cdQkljcpqe1Vd41dnj3QyZGMoOlJbkap7V4ftJS/4L6N+r4ij9kNVQk1JDoF9Iw1GETJ1xxIQzCZ
6PraPyLrYCAVOrnfNFMYugzn2tfXn5qLQHq7QAiPwYabKvFWWGEixkIsDCiJiYj7/ffGdv3JT1WU
sQuiDJCb/Nm1OnserH+nS+AZhX2KAqg+TfxYwv9BkQgGR5MAeCdBJOF11lxTSGQAKrD8vZy8UZp7
4R7kLdzVTANzAZeJsgXdEaSvHmbiP+AKgHiqVo46tDzDLxBg1Fnp5ZQtMplwKulxlKgZNPCWHvj1
8g/aMAKU51FGZ2azcg+9SCFdNnpo0BXAgRryClZZrMhrEr2O/TUEzbHdnkl6fyk04+amRxVcmF9t
DElHvTFRj0z8bCqfrH86CiJv0mObYZJMk2AntSo0736qB+xfRvqOKua966S1EfGhhmx1kqDWaJZp
4Nka0SdwzoqvmqkldTf5rwGJyPvCh2St+/wdGDEbhiIMVQPs0sY0bl/3kLkTM86zdPa18Af9jWIj
h9FCqzR5JD6WNcXQRbb1C8/83Wg61d08DNp1YHFw4mmLdA9fq5kwD6wp+fymtUO4/RQukHaIIMdK
jAXYtwmPeQ5xby+v5vEycKH6Pp/1gzaYnoE4/xnl6/254D9gn7WU38mfMb1ljvSfvMalkN2fwm+h
mv8nsABxIrodDVzZOqKaNTmp2fC9uqbVilh2CEI4tTMrTa/rxL6xoFYt+4yfcz7TijGLgh41rFT9
EIlGopkJGWo9ejUrwwr8NmVPygvva8QfoOmpHRXje3A+QnOcgnST4rCKMF6PU3N06Boka6E8IL5N
opzy77iBl+oqK+vJd9M7xUAj7gVTrxSNJxDahlEmOJMB1+A1tnS5MW3vuWrO0MpYu1FxC4vSbw0a
NGopIgrxf9NW5B2HxmdFNV/+mXOsFlDm1TjX/D3+akmg2fjrneJ5qt/heQVXjWem7dyrol2mmnTj
aU61KO8EIhihrLwA2L+bX+QZ2ewMZCfOvXsMdFmacr8VH+SwrhxSYw3yprtPdPjAeKbZG74TOY5P
H+3mSofvDk8YY+1c1pWOvgXq8CTcmDx0aAOjMUB4LbcvqK48zWRvWfrnTLAUsP1fLcAMq7zrRSt2
JTil+lWtdUb7YlKaG+e1FMU7OHu+ww/nHuj9/2VzDAeM/Ye7YL58KhOT8e4vAVAWRc74YW5duImt
32h2C0PenbLJ/aiJHSSyhnuxs9QEr6Fy/bLiQi+mwulXdeuI8D6STBJHHRr67/7yNCNrBuvwvB70
jBzbmaydrfalqKcmmD1kDxwDDDwDELL00VUlz3ea+/LWzjr/bkPZwoszfcyMBAfpt6V7bZbRhHm9
EE4G3FpUbGV9Cg+nMjrojgJlJ28h85BQrJZ42HmtcPw6Xhwo0tPBApLUWUn1Miy/R4fgMf/YzIE8
Rl7khrbuglPjYI4cn7HH+/cnARboO+jHLSEsWv7yPCuxBrYBrUtCkIRJl1Z4Ic9wQRdQj4l5cOda
N6KFaF92jSyadvZ9/HxZg5/2orwTe9zNBO+hLEDiSa3TL2UWQ/Vc9vK0t9q6YUoTfL4pUj6k6uPy
7sD4IkuIm2T1godkfX7xDcDLl1W3u+tH79uqCHBzPdK/CIVj36j5i7mLRFYYyTt0HVTpazUhfu9u
lU2q6ljHuc9t8na1akc6zTcuWoy3yKRfMK3sv+9iMG2uMaTrJVlbw0G57GjdbdKrOA8KNGzNABrG
/CGXR4m6JMG7xCLJY6fa4gtEaniYC9wtkpA85M8uvagNaoAH6xFvLilvME4EMZO7pD+h75mon+AB
hruyl9jPNG9xmBeb6Omjwx8BO3NIcMbaU2/rhHRCQmcq6ibcvULk2yz6ajMmSCPWzid9NBsrbSQV
MecwZMjgE3TxOdzARG3UnMCBlz54NzyfK6jye4a5HY+2fnd9k4dEUn7kSUuemtsVYhzlT6mRFW20
BA1HBkQVOunfwaGbKZS4Jr3FBsBqHIGyEtQ9OuQ7X2pSHm1M45wm2rN0PLt5Cdy3j8bMg0NAETUb
FGGJyhpcQ21P8TOOKYZhS4lsLQfivPOoExBi5RbzbhKJk8aNLxNXUZGIdkhMOW+qp8V9oe4PbZ40
wTYk7t2SWki7lfNSdU6DVM9C8mDrVGby6sSog0JiKTrTuGKAHItKWeuOiv5Gjrd1537bNKwhCqYA
TS1ak+o/rTSoLxXOiWQaL6mBxR7kAkQUZLc+sQ3gtnIDe4l2Wc817jxHieE/U3SZTm0a38BgrzVW
MLfZDdIXnBpYQNK2o5Dawe/7Caw/NM+akuw2k7IB3TKKf31hSQHXBw9O8XZedXxjYrnofEXQpwG/
zQcwTzxT98YyLC3RBf0hTZO365zpxEj/91kqnH9jKmrxsdLb9rtY/xA0UX94D2Oti5ney0M8PLDa
9xGG9lspE0J0+zd2YhZWr4ZyLpNYYBqLOMuaux5h8VXj1tbkclTRtR/joodIpF8N/3mq/2nBSDA/
iEc6nn3l/lgO3VsF4L+bSsiQlrNytmdhQVrMoNK33ohBGHrCF7OAKYLAKYReA7GdTDJZmALRjTNE
mNGeasMUoZ3OAsicUMIHdoTGeVFXiqBP4JNQ3cv6kczy1MIBmX8SgH8CT1n2jV+aBb1kecu1lEIJ
tGxFf8xaOyZwkE3xIgKmrV7nVlcA5UPG7JM89OaOPK6uTd2gJoWkFxqKrIOvn9N2Lp+S/yvaYJiz
UtqJg11b3hiFsFyvdwVomb2BAR8tc6hDqznhXDWku510TRZP8b4wzzrVBQ+rkFtJ6czl/Vq0vq6E
SC03KoVvEiEkgkBdLq+FHOqZY7SSj+rNqxGgVgYSFs2zGHYot+C3tDngjrVOm51ft9+2vpmHgD9k
+oAJlxharJ26HNikjInKkgVlTqmDL8l2afssAEfNa2/i3agXfOfKV0tiblJ8zJTdGnXXJkYw1ESW
3QWBGBZfAE9lfVeFoezMyIqylnIwHxMWoPaOC6n47G9/Jxbc5+YBhubfuO5qDbRGCIPilTybw/7J
h2nMXBLNw9YRnAOyi8cmMAre8NG7S0eCm9KhXWGk3jyAaVgzPUG5X8LsU8v0qmaNIUC76RaZyn5t
T5g2r/Qk8fXKFS0yiCFs1Sf86mj9G/huooal2xazWFOaI25Dy+BSqHnJYU1zZU9v/yjZfw0o5k39
QDa7Jb7pIj4RwH//VYKtWm9ompS4Mh2GKxO20vyEP1So2neT0aVfYnDGhdHTHBPsB7txOa2iUeJ8
y01dnEDpPRTv+rgkNYQQcpZRYLCxHN0FQYQqIJrnbV16yMqHQ4LL/kwspbSHBlQtSTT2vhie+mJf
/uBA3Rc7rO0lAsOXy9XD2K/3Qc9vO7/nQmzGdl58f/O5pHsVrmFPEs441iYT8yuTvE3hXUG+Vg+8
nEii5nn8sAFMLE555cVwSZve3TlnLpV+zOWzXahigHdnzQbufTErZgyoYwv3sjukGWjFTV5OsLoZ
UFw3mnRC0waTK6H0yfssPAQ6NBnmKSRpyqt2hefdGqX6yZjPdu2El7rdA00+skUYtMd3Swhm6CzA
nbyLazSGrUpiNWL803w/hgtzp07UpVjoNLLwKy17g/JfqD5O7pJPBndOiNdfR4L0bbim7jVF5zH2
3ad/hhyBgYT1fFWLB0BRJvZls+fFRLZ5WoqWYngzam12yrOMp/8U1X6a/Uw10dDlnSZuy2TlPreq
loXEgI8PdccmjkabpzX2/RVuwg5FMCYzolw5nTJPO+BxE4xLIvr/SSWuj+IgMq5u0NA1HprPP0Ub
6oVgub5k16SJk8lAHaWKre/bbzeu2kLY8vsRbnCO29cFDMxbLaCKJUlPTNJCISE5+WRYbKcMugie
qKnS2GxrZwHSfBboZ3HGoyIM3nbtugTo8o8JoCz6rTgaOP7+skVzVG3gVyvsK7HcqwChO6Nt4eDw
16fTG9GTDBQDFqJwIGteuvgRSa5R6p0lbyJWN5FCofA0P7GfbCrItVEm45FC6rleKTxnKIXgOUB7
TITWlfCtzbMyQmLDhrLJcBGVHxiqrRtu7Me//Q06DjHaqNGY+cgz5BZQk1x241cAolXwBrIdE8Cl
E9rrU9oSXKQPCAWz90ggHdNcfhEt+CMUtEBeL0CCeOP4sZOTAunRNRopodnW7ixUGbZAWNsmHnWa
eSfO2iWVVJgS6mn5HpbIR6/1Q4qEFH85gU9CLfitAbxi60ST4h+yYg8TNEoMIXvguUsNKDe0atxR
7oiGV8UPeMYrbmzWvG1nlKYWM8Y1bBAvZ8i73Uam7KKcZwZTC4xbvmRvVn5+hwhYG6Tz0BATf44H
uVpdsRzbdid69a58J9avGHZYOLPIszSJ0x2OLuvpNjzuMmPotwfF7e3MqqDcARu5bFlHfphpUXSQ
Y8vr5mBY8Ie/teVv03+OUmn9IXWSjB+QeT7zeX51KpeuVyoxVuSQENB019wt+XtodhXNc1qJHaVi
dpCkp++W2DshC12/e63rFYeBAU7mcmv/YWkEGZQPvVdA0XVLDfzNVE+7TP3JBRKL9wOdLbaiviJd
TId9pJakirwfeyOvOj1wEV0cvpz2gapk3/pF2R3DkPQu/dvbkaSvYUOQ2me0OoPjNKH8kUP9//p2
cNdjjv39a1PR1CfHbvBEmyN/WvSoG4LAvx0q+F7aoKVq5fa8gIMHd+i1FzyIetGHBjM6LgB+HAr9
Cp2NtTv++V3vZKW8hj+dT82Jv1Are4EO3u7h1q3lulBsXZAI4vqg4xHCr9JKymv3lsIS9EVi5+fH
aLQIVOfLgY4r9hVamle7I/fKi2TwK48zsuuEKhOZ9lL9r3nUIFvfj23fc2qcxJzuoPJyXba6sI9M
zQsxBeM29jKJ/3RqWLM+L2mJWSsGqwd/qa6Nf5S5Nk8UMkWPgWPYgeTx6KuAKlLsNgCGg2cM2M9r
ivY6ggfb1Sgr7FGho5HrbsNQfwD9Ucswjzddak+6roQn95UZ4zmW7OfUKl6GJo898DGdIEYaQowc
odmemgXR2x/hPDl+zfS6RHkka8rF1SIsJ8zF3e+L7Omr4mZ7vvDokbaUk1mHu+5Sq4ESGMCVruH9
DYb1OSt1MmYmXH3796MQbwIzZB04RCGPZcmiAZX9RadGJXaUahkGYK6pbjmUnBUHyJHxQuYAzdO7
QfjKrHoA/RecL9rZ5ADwKuh6PexNQL36rsQHKbEHmQLMB6pILxC0QGzpRwzbvB4JqIyary+9TF+u
1iJCtS6bPbhtn91jUxdzlWoS7EN7qL+UQIbhlfbWI1bZq7g9T9BjtAe3PLFwtT2rnZFVGotoh3Ys
Co01OONLHbZIAB0Q1rZiYAyHRv/wCIISObAQnblE4jATYML4CEznwuhUXDOT0TVYWou2+ayDFPTQ
tY6agUw9ZHnAZrpCaLz9ISc8BsK/FXERl0G+0FuUJkdeMTxt/uluOs17hY5+dPHbwk+14uzQxkRC
ofa+xmXDhRdg3Xvb+zNsCHNabU6/baOgYszWjGQm/vV/7p03DbDluAi2rmX1dF1MJ8UCnGeiMiW6
hcLilOFodYM4Ig8I0hvGwIFiX8QRoTWqpmD/MP9XZquDv7JD3PzwVPoker1oXBCB/yGfxcnxRTyt
XIulizv3e+qwruoBnuqPRBzKGdminOUh0pDarSqDsVU/lFH7V1eXZrMnpVA5LPBtuIbg3GJ3a+aU
T93qvR62OJYnL3H8zdP3c7qKdnCXiNKr9/lxaFxoNNb93uERs6g3kaX5Ljcv8+K5DkG1jgptEVfg
hBN7ufIxOcvxWlaaC5fg+L69Acljvpf/82dw5LI6I0QIS3aQBGneE4HM+gOzm/4ued5hANK0TZl3
Pt+rFMliBsCy5dUhqRUUVnJA/2NTQ4UjtnHF3AJqU/RFjXpXD4DN8c01rC5Nss6WT+ovuFc30xPK
yfHDEyYJKCcv+Xxh3GxWxlwUuzuqhskaB4q+CI696Z20uyJL32yDh6/NGFaY+x7XBuwePXqhIL7t
GzR0JL52g21vtR1J2f0m1WF6zCPOnLepo0tTwdVKSo+yXZWXIykvOSSRf7OlCzzRwRIIbs6bdYqS
c+VUj7UAbqdpzTNB14Mxo6JOQmvLHM5/Rk3KwRm2FXNmEPVq0Q5v1M4dcRbVu5DFO2UvXYzqU8N0
L0VPCkOF4fSmsUqk1YgYXNzvQUqziHUJtcjAzin2e3/9Z7GGfz7M0czSeFQcSB4Gv0olGlhnaPDV
r3S1jvtBWNRZIEgKzxqAwlvFa0EdMUT6UEwfn5Bbpql4ss2VlCyxvfORXyN5zpZDhP0E/fIlgPqa
YXUAirDtvqm5aVgY+lM83DlBdwABDOsc84d61YGz9tYRW9sOveikbuMTLlkULiWmpNi9qQN2MRNI
Tm4d04rJXvcUTzrrlaM1kNEihIm8JFPNJqvIEtcYvOBpNvRcgj12w6h1gwbaUhIq0p5o953c8c0u
bXCqo3NSqoiz68gCxtVkvLGvOWeQ9lRMccq+euBJmc0LiFMc4k1nfpKqTxNHBGK7M34UvuxD30cS
9iYUsoFDH+3Af7iVSeKod36CpLm35GkbWC+kMIa4qIUpWl0OGSgLHjEmTjqFdSVKcrUrXEsGIu0y
uHQxCcVniQAdndbRAAla84a75cS1UgUPYmADAF19HgFRR3+knMlzG12jWkVmo0UUIVlGLOflhk7L
t7qFzg3gtXHwyIqH8RhlQJQeigeK5XIrTC/J+eV1XhBxVur+Sj5VxrSFxMEbSVkIY0By7go9iJ/e
6mzFEYnW3Qn2It1kZ4gouuuGgu3sEUvIXsWto+V8wBAfs7i9gR+tRVW+a9PjSgx7V2/3BZt1GJto
lCLsPNn96Or7+HhnrySMEYeiPJKzEujvivHZOKCULfQoWCLg+zklliP8RF1ZvmqM/5YuYa65bzLR
qys8YvDamTbY/p3tEf5MU6IdQwXw1RdQ2lSuRh+JVu/rMsYCfL+l1/m8cdyY2n27Huy+vdnK0A+l
qLXeYjEUCSjmCrL1klcnCzNCoCw1doSkjHsLAZLj8i4R4y46gRwIqTEp2nHYeIL/2H7S6yGa8Os2
Za6I4CikYe0rLkuy1kQncW24zDUpkNs6LFkBm39AnGxYWxHUHbRKhszGv5ylixlS9V7vgDbzs/4Q
tLVtZGdA6ZP0vky69+J8yOiSXC/+8BVhon6Xfdum3CE8ZqJ6/r/O8I/9tmF0+1vdsZZCdYR/+xCE
LSHbE7rO8qOda7kJ5SywZNviskZVw9jWwJMSsh7WxG1EgthAdzyM28BjELtXGrzRXJza9+c0IJq5
Ume2of/6B9BvV+HBAl9s+42wTNtmEszwDRoAA58Ld9g8AFh07VzgMGsF5OWBgd61s+zkg0AIbX7k
EcPj9NRapXNaVoXSkCJAVnCkTX8xpdOW2rX6kjqaa9EnjjVWZ9+ToJBuelkWEZWxjkcBeg4anga6
1w12XlonGWva6STTlou6m+badymYlXtujNxC5LhhegCthiXDsyVPwJjo7si80gfIMd5lVLVHjNUW
JvNB4DZW00hqh2fXayQg6Bw1xh6LbBjkGbJEnO7LXNrP7k4QHL7HQiT5dCExWkG2CzOws5tWGKZT
19+1ZIeJ0+vn4fj/kP9f8GSfSBDJ7N/bIzdg14dLWbQsEqRRZpnsL1cBHUW9pG6SrGqVn9QVzLl7
tI+7D9muuCveK22DuXiupXlSg6hlSqspiYisO8M5yDUbWcmg9/1GKTyPkSG2MOi9Vk9H+w51rB0M
8Znnd33rnre4IyeECiwnYYY07zm4g0D06nqXtrOid+eIa7NQArjmBjPrzXjthZr1b/MIClZ762sG
ZNfyXJRCOuwI+H/N71uohVEbdQD/Zcn3ksnGE5yOBjVrSOP+S3XmqEKdcnt7uq5MWUNi6HdYKm2P
Ibv4/vobw5K5JH7bU1Mu0MbcnfAfHr+r8FZH2x+p8zC4+FLptX3r4ikMxAqGXTXoBr4NYrBhm6ys
jyq3j2l0ymUs34bv4p9mUuz7jjFKujPJbhubf6yB4RpbJNEX6Y29n7WL8/dsa9Lscg4shjZ0ijPn
hzgWml5lxzvrJFzP3m9CZR2HMJV/JwSRSKVl6khI9v0GGTCtoqA/NHLVm7kdgv9r7MZSrQJkFkwP
moQnB/F8QzcjkNiIJq0UdAgQxPRq+KDDnCfH1mVTa9lwXU4UKiQAySCi+SsylOAvABVaZAl+3kl0
bx767rv9mGERfVe0MQ9rsFUqctNLXu7h3LraB85MG8slEYIRCIHk32+gJik/svOS21U6fV8OXJu7
ALybotwInBQaw8VPpSNpdlbizec9YCM7lpyp2afSLs59/Mm99IxX4Er6pPp4CFTKssBLde/gqpvf
DPgon+iqMG0i6CCx9thb3DpkTWopbJ/ANcmHrep6+Hz1DaMtrN07CaCuys0v3xd2rLZRaY5+4Abn
DzyRbkq1DylBpQydZsdwzmqZr9dOvOFNU5g6MrwME4lLDBs6fRh/I4LQLhBslWU9xQSGrqgqRHNi
rjlyW6mD/ZgOr9FwjIckcLfqgHDhOCv0pSF9lB++rH/8BrxLd7qY8EWSmAelrcriJrDbnUQLEg8+
a8yEzYNY+G9H/IZoR+LdjX11uu63Ybgwsb19DTs4oL1q0j+pgnbcbDG6gI+nG9HTbNz/12D9c2sR
MNIJt1+ylN9RPKo21vhbZokWTIMV7h3Vk5aU0f/SQxB0hvZqsIxFajqeBfSGHLraJyHEFtWO+9qH
0rNAUjuA43TVNaK+ZIzEywCUhNKLfqZoD7NXx2Czezoyu6itJkYb528CLfIC0AoVRmGhiHySftZc
CuCQKVeB3WBq6N6+PYWaZanvIxiY7J3YQ93azYUxFwRCjeFK9lJ4a46OHCTOJ0IhUqa12pS57jSF
rKahYRuh2aWm/o2mMv/bZ7PZrk7kkqlQ6wqEtDJOXAY5p6IMY+brxpm678nWIqo+s0GYGVMzEhmv
JdjZI/8+srUgCf8G+l6nOydnr48Khubudk57A0IZQU5S/MZUgY4FOnwPxRRvJ1+VL9f276sfg28m
vAslCJg27+9qPG4fAeS2/8ITyh8UnotegGhhoSgp5CnlC4XBOd69SipJlLwwiqyxua4Q5YXWdMh1
kdo5XPQTl0e1P0aIc3sfJmFHV+/gZdAbDBtgYFRH5p/GiFb1AAzid2JbJUAJM9HQ2bDxF9tOQMQi
EURqngVR4glYJCvuzgDwZ3Tdy+gu7/N5Rv8o+35/NEW0wuyX60OFKPqJHKLedPHSe5ZJWJdu6wU1
I/eOjoify1e55xGV9+y2NA8zwiXjFhYCKh5W7rGteaqDjg2caP9USBGhWNBv0QsbfZOkWCEpyIyP
kOFy/yCBBNmgGaZWE8DYeL6cUg3MVnBs3+seaknBMamgKw8GIUeKFvTeLGhRj3hioLXHVl32mJxl
niFNNmeurLCbotnJCS5WZ7hxSCT5Oygrs6IjVAOSM25ixQuqFld0S9zKcuLowRkWz+5f7ii/6D7W
tU2MelY8X+0Ttf5oWsox9cMJEK42UX/GUTvA+q5sHnY2yYenLMwSR6k0m5a8mWDtx5W3TZZYYHkt
z/DicSVYWhstndO5zvoONXtlvPh/koD3VaIICR/CBBTqUvJfxBDv4OH/F5CWD6lA2/BnasZ/Vmhx
jvinjpBu158Z/5d0BD4ogNf98Lj6A6xeIM/YyRMHhLt0KudUhfqgh1RkUF5I53A6vVY+EoFubKt5
v04MRv9G8XtjIDS1l/m0/utM5BgcmmnZEJq357AFQ5synQ7C+JTYZNa9UboiwVjeAm5vAThwCFBL
MJq7lDD6conGX/EtRdxx7gRJMGNP6nCLTgxLgIvfJZFJhE+sc8lITyKM9iJdJVkVdDoVdkkwd+rf
PzO7CP7m61BgNjCzRMRMDmm8EWoyI3hxUJl6dzpoWCnf/wRb9W297ABWHd2uK6LSJ+u3WSbcjWdA
sba7nu8zoNRbzNAMvpDJGqEUlPL89LzRoxQWRBHQHorEb5eFoTD1BChNssHwKPuMGIfRczV7qs+y
EIGg+QtzRD42XYb9lGL+cyFYJMYKimtXe3FiQaP/qeJU6PgVnPTYDceioCZD28BG+8tGlZ0GCw6E
Xq7TFFxgDtNrdbb9vFwG55JoSDA61WXx2ZgLV6TkIWyK+YLpcN8+i4TwlHke2cacf8wE7dD5MWwm
/mJRiRPt0Aod9oWWJsPTBc0mt+FYbqwHn+u7SsTdCJzzaYf9Pm8PXZIOxdsd1j8kXtwJPIUx9eGN
kfPd9KSZbeaAWZ2WmHFBiomIkwT9Q2BGWbt9mRPJuLR0hTPtb28CCGDu8Nm1a1jvp0T/kAigGzt9
2pw6C/F3I51YZ5bjz4AAMC+dB4ymDCU2cmcbduXiOAGGDjZYeW0Z5CXikcAZH5C0mpuTK3DU0kNE
B7CtAatSnsenoRUrcpfdGZEm4pKwAGuNKwtIuRPdNv54XfxkaRD4Q4XR3xB1dPnrVZ/fZwQeSWyW
8S1p2rzPQ0VTJuoYoJslcpgvxBZkXkWLxgDuYQsa43+Rn+4edMaEkhpVUo/Rh+RgB+Vwmivj0E8c
xU3HyHdmzblTjnKQGXuEEveCTIvSWw3WXz0X524k2FAk+pf+cFkVeOUbLHXRWsQp5AObs9Yg9ljO
JBkFXWcHQ07oaQ/1M5jnv6AG7wzdbW717RMLQo8ErmuSw4J7N70xECDBw1OCHUBLrHiN162EW3f2
Z/3f8yU4qMHa5e2WllU061Ja2GoeGEWuTlmYVN5lqba5DfWtSpfgjn+AloWqpNrDRYK6FWkx3DAq
KwncVr9RpFJ83ZLoQzmF3h8YMmav1rA50ARVta+iUj1J5jwPs4dq6fYkgZ0xIlcTbaVYEoMfCm5z
7mmK1ny0WzKUL2PmuePEDkmSgI/OdsBaZ/ny7ShWlervj4OMk73u1oAHTS2gVmWFVisLuLYPHE+d
7YzdTq9ov42/3SvdQeDXE3GoAJXMOkMpuQIX0u2g2E6bnPCs5RL8BXNzENuuPq1wKWFSr4RkOXXN
UKMkVoXxoQneaS0yIL9qIU+5ru2wtNdQr13yzPVx6GMj51xbW4OAXwU11fABfhglW8kjZFnjkQqA
pca+rZUjyRkgtHJbSxu3C4iiGYJErePi3OIe9X9gtgXpsWQGjJKWZR18HWc+zTipsIbCM3dOtvd2
qRDTVPJa1Rt0e1HsLcRaT4I/bJJcJ3uIhFSOUXyVDuxrmxombU7sBImD6g3hB8IyDvVfYGO7wiJu
HPPMxv2pUNShJPN6T2z1C/57+uaHDsew0rGRi6kfLERku8r75Ua6a4nY3K22Bscs7+Q6AcDRa+ij
IIihYgOBw6LX6WqpYA4Vq5y9nw4aLOSVgq5KPCO4U/J/Kai1f6pXpCCk+vD0uB87saOIoI4uuTPN
BmEQp1WRmXkOVNNCBP2pSKxES09ALvWYtfOGCxGYPaqAyGdNZfWBirnxC5JGF03OOc2eMcrN7NTE
4Y/hM46VUHcFXYzhyf15d4KozYCjawObAISLUvpwOhknu74OVAGmrRYOjtGkpdaxL08U4A4iKK/s
KjsEcmyZ+h0wBt93hPOzrbcRMSsGGWLO1FSq8F7T/ShBzs+81ARKM9MoVCjag1QVOaJxOHOAO/ub
FwbpKbvMww7cSil8CEG+WtVfZDX1ol2BDs46RJpPV+89CyE0nY1oz9cvJmwpwE1IpJ0EOkd0OY+i
Oh3VMdFvndDv7YBSZ2qO78Df5/eeRn4m/vDLe7+dBjVpxMYG8xWbtNKTF5h3RLvDfgBxN1/x4qxK
SFJ73E6D1fSIVXCjcx/wPNkkGF9VyzWSybvmwF5jVAoc3oKCNGlqNExDZTcrin4stBUbXyj/X9Z0
fHoPTv9l0nSSSjM01aoz5c2srwsfX+6icsT9MA8v9n2l2RFwBgC0y79saRGxppmBugdY2pRDTMhd
HZVrFP94Zna/Ie4jTTm9NeoO/Eq5gn/0y+j7x4BhRRJ5zZl2RV2cxZ7BYgrmFBeuUZEw7D71xd2P
S6w7mR1prlc1Gw5xXtWL+Tr4U4xdavP/RSEkrVQsa6PP1FxHJ4Dsojl88bfa2TfaumsP4Ue5cTDO
d0H6lOunE1WD1d5bXmyijuXg67WyCKryU9y9zg4F2QwFgTzdh0crTkXa7rfrrH/fdyK4gG+rAnsz
VNchv+lIFcHKOmnq2yOmOM5FgLshgvb+LdNV4w26qWHeW4uC17KVxVSb3CitxyHMFT7aBt4guHB5
5ijT18V18QQ3SxzsMhf74q4tin/GxaiNR14nXAvdQorXENzJTjHYEsO1KNouO3VnHh7eannhaf0E
yWsSI/39yCplIFlUbksA+l+EYyt0Hd1KRrEoZtWht+yWiiS1+VrMqkv2KTepOeSmKg1TKMWcL0HB
fmvRNpipsYqC9QydIiQ1g4+O8kqWPlRqmBKaMkua2uc4HoYyRJthwqlSzpQ55hqQTssUgjmRnOw6
gKeSjsvU4dkAAj5ng8PV6ab4Zx+M1qNrcWjxWTTl84s/XKbq+aymAkC7GT0AbwEXIsCDyR/NkhYh
D7BXME5JLsSAgertxxOxNqyF4yePX/nDLs3qi709J3dOlKnY2Cz5m2hceg3XBRDgeBch4C4tRpS5
IZhfIa7S+ylM8Kw+MprMFj2M7a6W4XtrfIYeDwCq0gzJOsJzLQ+DFvbI0J5UAg667Fl1DRc6cc+r
vKnPJX0bwLEyW1Dsn0WqqSPWol6Ool8Z4RKnEerJJJ2S4BpTQmJZIAGaa11G9VFSUBKmQU2nhAK9
uMYLfkP/ZbNtGRK7hTOieUscdOYx9Otwa2LW+nRJqdd7s6Mc2k8xoUxxpbdcjNRpXWTiC9/RL3EI
IlzFxE+VJpEPs8cn54jS7/coDLU/hFPaCyxLl4RDRR2Scbr8xjq92/AvUBevluMjOWQlu63e02sh
DqRJRHc3yMe0jkKrEqYWacvLxgxRDu41nJBPRkumuOW+ogDjuP1MK+h3CN+T7Jm3pnWUQRouk2e4
SRAjUmtOCGMd5VXfuzK00LNVycwv2Ejf4jAbT8PULV5P8+5j277hj0vBf1fQNacM64b9xbTXfeYv
uyBLsBq+yN0K8R6YmOmoCgPpD/OiyMn4/QcZYSrtYCR/bStcAlhHUQUcqYdqM46PcGcSa15nmgby
iIsXso5ZoJpD7Wql3qJzABaGyvxNS2U25m5S26M7njmxKFAswnXcvlFU9RzcP3I39jXmMKb/BSAI
cNqjn5S/oMTHzRNoOUtNFptYvXOrWbm1P4QvLsyStdPyneIcRt1NQ9BzDzCR6y9EE7MNe/6BaN8j
do+n7QYwJaYdWmoI0+8VDlwhlj+SeClQHisHjWtXFu9sCuYDMPTeuvEvcszCF0vFof1rqQs/hFbb
4y1BVZRBeioT7y+o/XQ/Q+NfCiwnHfj4AkBudMc5SUfllxUwLCEWeA05iznn1gDp7R3xQYGQaYmc
YC64nJWpb7G0Iq9mnsEDhsqdWpDXKsz7Gw2cxvWRHtkQyGZegLq1EP1CGkXiVligEdtkjhe6RFrC
M/kZUBBmWFlRH93QzBZUOuZU2APUYkJeXT3jtU8lTD/9MgtUqX/QUJ9r1D8Xjr5fSZC6L626BNN+
T7Pcn9wNk+2o+cz0mVPcpBkADbgoa7KU3FyxHeSVWLnYg0ATVzdiW9MAJt/deIAq5AWbTXByJ5pL
Q2uSoyQDOr/NpUo2tIPATXHmSjleP434aTvtlDCWPYOF0qeMhJgP4VI5M6abkDo7LzXaLZ8ZbwM1
uBoWC2Zf1A97LhakkKD1V6xa6kupzdyPq0W9/I3sSMBhsFAvabPHb9O86joVJ20PjcwTOuuFvn3p
gvnx8rErUxdLTOEPS3wK+kx92iG672Kww2QDM2Mvj2A7RisJsxRZSgGI2PDVghjaqlWrBLoQFc6o
+jOMOpg8zOq/JJbLhVtFkJfp6lR4TFrvwiWUzPT7b8mU66r1vzwhoIRumaPxNpXcr6lLw5t9i8z6
/anxluv6kcwPKOqE4V5RTztUrj80vgnnH5Hu/qw/EvXvNB7gfk5cQ+YmWzQ6W133D0Mh9qUScOdT
lcxo0RayV78xs8cUJRHasuDQcjQ2FwH2uJakFTyOPsJ/rdicExoDqE2aX+e8vgaYxa85CaRsEPtj
ndRlgE/Dnd5SmuJBF7t4qP2rW/82Im3YxdxZA0W7biKa3oqP6NMNN/2sNZGcGqxNbvxBXP0gkupf
cj7MYpaho73WTg/KEX7x6ppmMNTpNbT3TkKH9REMXTc3tmU6HoRZDnKM5FgJM4ulkC6WPqGRHd9X
FeL/ct1GteocVs9O1EVq3Ygt64dfALQV9w2gc91UX9/15Ql54RlxQr96l46PTsgmbOJCfYdghkgt
GwmC4oxe8keXN57InLT88yfp5CT1TKWG8eSVVLRIrNGlt+P0el04Mu/iys3+hfFBt64A8gi6x8FN
KICGPCycuXTpnvEiy+phH3/4iMzSczWnd1uQ65rNBEX6ZaX0Zyvj4CdStZk200gyhSUF13hzrJ4s
YgRsW8g47TqYCJXM1bw5b802pFdZxcBOmBwoKXG8FdUbc0sDmgTWHISwDSoIVrdY8sHf0x7TIsy8
pg1qR4nlQD1yrB727yI7PVCSeLSNjpXWRUCfJG14DO+AnLFkzvOpstod0/mWgimapguab2wnD0O9
DFSzc8k5G4mdWz5M7Gf9P/IMqhZAXnqhJPacoh9Zh7UrIgpGVgfj8NzbyVpkxpwv9X8knzkxuM08
xpULibS2yaYAIavAzFvLshnPZj16UHA+4uyGx7jnSDsNXD7J//rs0bkxoY4RXemYTMc20uuHPwj/
lVXHJ4uLUomk3TTaEslQcN8wckvyOkzVOx1++BbfbFZu1gLdBm1QE5ldXVPksXw6/JqjPEIIy5/B
xbwkJ/dmATSw7Juvhj3F5jxMAtELXbecF6Fs0hb/Hz8j5A1XMJ9qfwCUf4nYgO26+bxJJJy+WUTy
QrY2xyyjDfWRUFQxEKkvqTeH9krOMYUh8CMzcx8eiDJLHi4X3qPsWYl2p1UJlqBRXFPxN+yjh6ah
zDmQp5iKf9QBYNszk1pGDJ10ZH6NGV/oE1oY0m5OX2DV2XsjEontSLLGYfZFk58gV1PirCezQuMi
4AbPb2lAxJzBcWTyZJjuX2kjBOxdkoCmD36mrveHOLQyDZCemJy+Q0Y5PHdhc+/OS/3RYYUOEq2I
k6AWgsNaPp2774uCQMjL9tSKe2LP0SiyS7ue+4F73t44JJVGoZIoiXWOZYVUn2Nnk+r1jxb/7765
9yJZwqHNr6ZoFisW3g2mcwrmJQzBSuELA8iIfHStm/EU6a8xb8HX2mWZZIwe0K0pVImKCc4DS5qy
VTYEhx84xQYCAmO0Ba6d9xZOCwyEIHFqrBbtN8J+Fmeq+aN/w3JTZn1bRDvF2RUXP9Z8DWT9AQng
rkLQxaqD00RscWW38SXyHFxary1oBQYhgdnswHb+Kat3X5xpeHmKbDkyMjnll4GxUHMxP78vgVhU
1XZ1tpG8SoiZluCukgFJpR7jSfQdPHhvvSePQEeSLbglm7IXoDfcD+8maEpp1bcBwu+WZSfYiC66
VSMpV16omrZ4pUart1zayfZNQRJDvn3SOX1b0is/0n77+jL6ErEvR+zh+XDr2d0ZnVuHk4tnyEtc
I4VlqYEqu2IFCYwiaIJ7oHNR20qxK44apj6fG2SlDEQOVbtJ8nTwvg6U5x5CVNQRH/Z2nEdvMN2Y
elnyy18lxjxRgL//nz+aTvdYZyFpkEHO9hEP7/laM3gxBpdoiPI4bBMVZ0wNXLUrncuT6PBkwx2G
cM/7Mf8gVaHn/16AWEiZarLe103P86MJL7YU1bfk2L+84aRr3hcsqGKc3PzMMEOxfHF/I3GLn0E5
M6ynlgOR/bObYVFTbV6DH+rJalBULzRkFHUZu3mlYSWPF8EkoabK3pbpz1I3HolKLPPCB3eav/RJ
9Pa2uO3TSqiVU3hzT8lh0S8RrgIKAmnJ5MT8HlNs0FZ1pGXAcg1/3G0YCQNKJ+vI7XL1m7rhn+H7
rFzHu9NWvdbf+1A/s2uT/Tv10LoVpkPguJOVpPbxk2MqwkhXdDnXfT0nFtWBhdP76oL9fXWJcgjU
XbMObC+Eizd+5FVpNRcXVHG1APqSTDKKnMhYyifPO8nuyWOIYW+OFWVXgaf7pmErRMIB7bz6yGyV
XCdmjk+jc49SNn1ycYv5va33eX19TfdzkJbPXo8olmsW8d+IZ4CB8EBBQxU1XQvQtJsbrhTPzJ93
nfrcoJF963e3ZL8n2U+k/o3kBncrXrBuod/K+wBDsiqUQBY/K5lU+C65HWU2vK9mo0BQo0BMrz11
9W28sqG0huGRz68W7khtuU91NgzV44EhJ3qrSZuw663L2vDlVTGXIPx9RMcyyblT60Mxp/DhXfRY
/jRV0+j4NwnZ4LcB2NHjf5JdUkcZW3a7gYAlWOe7J50jGJk/BhOrpr/Jd568YGDzl9Ie8woAV8HU
mlxXNtsNkj4qqaEpSdkBCgE6RuJfFrqXYa7mHkHdfrESurHSDVJL4WSrxge5rj8UXVKDw+7SGG7D
L2K8qPjMgwl22Nl9X9CStcUXfIMeTp1RuQLFytSoCSqFm55pe5T55YyAnEwK6LkK2racwq2I7QW/
2CEUNVNBJvYAC4myuVvITkAaatTC1H9jl6cBudhoz3JENaEjnFJNAu/hIK5VoZ79AmdnflASnn7X
VWApFuJ5pwSq1FFuYzoYkTS1MLLV7AxBtjEvIjMvUmT70oyihgvFhd17K2ujL6IUMB+pWzcg533x
i6koyKb6E7R7vbGQLAEKsfhsF28Qu8ZB6t+4fOHdnRUdRo+euqu1+cpxO3l2+TfM26LsSJBvJU1d
6/CO3YG11Oqfl/UpVEi9VXiGFpdV9Xiy0YPKUZcrTOvtnAxYGPWyfkND809KxAxFi+EiIHcSl4dS
45miOWUnTxe+wHLgCaxucfH20HJ/nl7WwPLqBf6bOpa8x8nGd6G9xgjAh/R0n8qbz6MauCJiSgsb
fVs5JqEjlrst+raxbzVSA2WGuMC7gGupstPi7H14YlEqT+OVUbT3XTegt4E3BwRTNjyyrw+Nxvdf
hwS51mNdUnFy5EoQlJro1xSRI6XbmdzpEY+/IVUhHEi7WNe4dSYh5XmZ+jDIl0HIOuj0iTgwbBWc
wbqk0mshgxJtWijACTaaeQ2SMTdryNDFp2Vz7yKRp9JUsV/2HjTQW35AKrwLgY8WxK2b6z5mABVr
dcQSNg+xy2kIbQVDu1PuFSGANBbRUK3/QKMKN721zF+jaop6GGmwEFFChX5KrerZJVvf8lndnvPO
HYPxFhvN9QyT9a9Y2c/VsMBLxedQcHslcL/LqiBKipCSop89kpm1EHbX89tveazTYPlGYteWG8qT
7/apteCl1NdQq4jeXGHlkxDybutibPUv8aTcLOjHBc/hDF1HJAd+1t43Wy3f1d0zUICNrtNK5M7K
QqTaP5UGHe/kj1kEeigVRr5dVbraFqJhEDj+q6zZoZ4niohnxfDVqWtjBFh3rfrvnOfciX5rgqB4
+aLpRXnGZH2TZJd6Jw+bA7kSMSWOd0magUMHvKposkGx7eGbhFwICMtkpy21oks2pLYvVyJYtuo9
be0RVpdosqs1+KUMiBcbIalg/TDzC05tzYYhZK8XwEQ8ox4n1g/w/hecMo+fdV/qcFUxs3MBZ6+1
33VW7lL7Uri1R1hh85DShzqmZIEa1ycScUoi2i7/g1BN9LRwYn3RPrIZe5jDtxqa/V3VHlXCAWww
KXcO7Djeg+YNo5YVqifAFvuBy+nYaULnDsuDw82dAe69ujHe7CSBjnTikTZA4pu7qliYA1yZVPXS
KuwGc0ZsJbgZOye+TAx3nf7EHoMsvNjEyimbH5Rr0bqVuPsSKaeEsA/Uo6eA4FLGmFTM/F6qqzQY
ym9QzXlLwndjpVC/oFQY1m88uY1ddTVG6Ate1wdbFFjso1cLSCvvQnP+BsidaL2ATTIOyBrQzG4P
bc0ul7qVzqPRR0eOvmy+BjcukOZ4qRKlyFlYURI5dVRtvyx/v3uZPchdT07/VzuF7QF8LrtiAYu8
blMqjKkf2uos7s7BdwuHCe761ZbO/WGcFkfzPH+5L4RDSBsaMXzFSIARhWBq9qGru/xSMooVvE+A
7TT9DhWPHz3sjTMno+zU+T/BgvueZBypb9uV/sRIC3e28MHcRF9j3Ww5Lztwezj2I6UVTNELns0o
nMtN56Cq+Pyihxgn8MWXy7Flqyd9HLnAoRBexNMq4mzTyf7lEjgY2MlbKoYltlcjAhmqgvZLj/2/
lAFcJqCQqBd4nPKiEX6MvhGmlgoY3f0LIN3qD60SJOLTTN7zSu935yhfBxDDhoS2qqi3ZBjMKZi/
By3GnhrmBlNeBzn1PvvNBLtxCmrxb6TZvGiSaZbaetHWv4daZ9ukCrfDLwjZ7lo2HuKc/Mm1Jbf2
NuqHBhvoKGHpnRU5Q5xarInAiPtmrQNxXQOPmjheWnZCB5CNvcx1gRMM56tCuIQ8sHQp8+EcABCH
Kpx8ObjJjoaWqrT/4ZxrsgZEnObO/uAwSvjiDOOC5YcyAGXooVcIMWB3qQJRG1Uzyaeb28d0i6lx
pmyLjdMOBpd1wnQZCQ2RG3gRba/cEv+ioXxF2qqq9AmBHS7v3xQmZd6PpylnuQgwUJ/jolRF73lq
5h5/kJw3J/m43pMNxUM7C4ZRhucsvt89tiKlZ1Ze8cXZeoT+HDFaacDk3Ne469sWs13DRXjM1mFQ
v5UsDwTNqx8J
`protect end_protected

