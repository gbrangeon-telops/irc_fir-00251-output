

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SOOYAbmSVdMSmEhVcX6OANZAlRBhIeIgp+j8aWie5qMiZZfkKWRKGFlDj4dOK2MxGgpLi60kolAl
iwo8CvQQmg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XO8hvx7ayNrMYNs+QowHbS9oiS1GjnY7XWvxUBWvS8S0pBwgguPJgxI5Jawjx75IEBra9z6gur8D
+8bJ3wjB5uOzP0Op4TufbsYZTMy5/IRaR1m1haAiZDNWpnRaJY0iGIl1ZfXnFFB/FNm2d6rg/H7b
+K1wV2KmxNsYmhxGeUs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qrXPktUjITPZaeyYovMGSvjyrwEeWSEPCoXArB49zu0J+taotc50izauZkw4BvtuT10+TUqV3pWu
H2Y4+wBhbI0avNdhBTQ6WysNgxNkl4xSoIMSUDeWLPrThpvXqf5EM2xFWnYEsoSt1fOlTzsbNp4Z
xTF0/8eRzGcTqQK8goNirFS4li1yNxnvMyocM7UB0Hgwd4r1WhVfwqexmsE2F2aKD0WceDfUKvzW
BkaD/pggzoFKe9ZBj4krjm5QO6MJe6tmyETtklCe5Tp5KFVAoUG5SSUacYfOW5JRRQQN1B29KV6+
B/PXOjnEprmrDoW2/GvnZUOJ8iICUgvcDDx9Gw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RfdpJMuL5lneUspdc3THLHWNRfMy7ZKvo7MAlgXNSeMyJ16shj6csIbQx7zWlYY0s5cmQ5qBeuky
S0nRybRR8cWMHwN/9rEo4V+uesao4mJ5GbtqRFTH0pGXUIW0hSA/qLXBAZCtANiThLFmTTovXGQx
QWChhP7QcQZsZBRuEUY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KfAPtRUOpYg8KaNj0Wxd1r4Bcs5Lt64mregrxrObBeYBNNIje2iGcuv2d5+PQzzomKwP4NoGlbzx
CSYz6XLlhFat5X0Kad65Lvso8ilyZLrxVgz/cQQVMyGtqJsflyi+jbqMWdWQzDlLboEzDolIGqLM
T16l7bjdTv+UHoBJFQNNpgCUB8RCwZwGjuOrDkNOQRBxFbXP4ewZBD1TITGRJ+9yag2oeIszJxFS
OnxOibAvqbpn5K7zetHoNiQFD0HLxODP6ACT7OZWy2QVwDRr6smLhIBBF+7E8S7up2WgvZZ778OW
7Swo175PkHbmEfmpa+y5XkNQNOq7GC6XNCURkg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11344)
`protect data_block
6wsUiHnZjyd5Sm809MO4Rye8ZfTpwzqqkQfzG+GnnXoj+XH2/73ucp7R3lQDoVnM0bloqlbhfXEi
5qx/e2nR+Efd56eyDLcrKyutYvOqm5/dw9sbyUb1bjfrKSEop+iL7fFY2jkQqPO0NhrkCq+uxbAL
YAs3X7Prt9EwVTnPUz/Ot372cblXRqKoOAAqP1958kU7Hva0yks1wkH6sCcEW5xlnr/Ft/NEH4lm
XPM2Ach5S9FrQfRZxd+MzktDCy3sXxl2eMlJlJP6VxFJHxVLfK1Ec2gM9RCjDIjz+7lDU30Cv4xI
YshNWsUVQPgdqVdw0bfHArMwIet368zk1m3mli3lkiww7kTK2O5FLjr+iA/0Z12hlncgiJ9g1fnN
CSf8d9YPfCr8XmMkHVnkQaH3EaGur7v2anBfAb0nzlEUV9KEM9pHLt5MtIalLh2G0KozAFH37MD8
sQI9tgRhFi3HwNUEFzw5PylY37C/AqWSapXJVLThBDD0o3oQSbNJdOUhG9wItqngspHGCcXBRpe4
PfPCa8iLfJruvd+gruUhsPvByHsXMiEcFnC2YV6HvGASFpMXh0/T64sXi5uOXDNoWhRQEaTQKQO7
LQF6nogr5p/xT3Em8kTuidkVRPkoqmNjceYYgRTul5s0xR7StXDr0su4yOxVsH0rvDqmcIM4Zo8v
Hcew4agJ1pAKpHGzy34G4z6jXkKXXcPLNHa7l0WzFA13CkFiTJm9C6ufKyikCCs5tzLz8ngmO52V
yQ8dhbZwW59CQHK7SXfw4sT2v0hfzKl5ERw3+unX3WL8ZtZkdH6boWfmYk+aFE36ih9bjwNCi6rQ
OQIWTWcXev4SArgFi00x9QZJxspYGeOFJd+3RR98utVFYY6+u/dIbjNITgWm56mtCt41EB++p4Pu
CHkJRqMfol5NlqqahUBPpMVB5YILr7ElzmZKd97j5Hhl3SErg8U7sTxkgLJ/wEwhcnck4j5rON3C
1zrzaGxe5sEpoza0EhlCB5fm/N9jy40799CyvtLMUi9FiON1vqGEKYoJ7YOT+ecciOsJ3ySe+tQp
PLoOzy1Hv6kQhWqWEPU1NEmnkTAI1N/xm6pvp5rMq3ILDPsz43YBKN9TIeI2JqyJ0if2gmiRzNQj
UCMBHeovXhpgSpZpQ7iAinMBvDd/BBPUm2O4rI0QFUAv5IgpS6SmhVEHsLIzW/m8mp7EqZ6ip8px
sqWTmsSfYzD7Bec4+TKgU8QFNRkZ2Ujy0om8RV8aIGQOUi7+TuJM/BaLy+mQxTqpEN3HLmr0ntqh
4hvglBkTPlQl92OQBRy8mZVxYELZ6q0Uoplvq3+dGUsLIIDQRsOmsXjkEZ5FQnBVdqS/ad6qNNF9
Dc/7BsW0XbFRvkdNr09KapqKPJy8YWw2nkO4SFKYcKIzNhRbKdLjiah9iqJHPeQD3v3ysmoY6Cx2
VmOzKVks7O4BpUQx+2RGirB5ktxYxjXiMmTZkCS/wFaDBkdGUQsi9VSgU7627JNjiylnSv1pQ8St
Y5UQTyqEpYZFqkh3bsTFQ8zOoYcj3CeqbrlRDPJMeNPvxujeWfZ8l0lp5dS4IeEGlir1EzkqICer
ey3vuZNwxMpHNBd+JPm0+VEJb/UNlpOAUfmK3Q//FzclbeWmk/Uuo71ImP5LnUIroN+u7ZVQMS7h
hQKyavvwVXqylHuDiOHMMyDPSGX9hfHi/I7Eq5/gSm6x58pmrVIVI0G89sA48/n7nVmmBWPdPcpC
s+NDZU9DlVIoEzrwyCKn3SLvoghItaT1W2l5O34IROF2udI1R9vEq8X1LpUWbh5xZCEMMARDP7n8
xPSTblaIQS0To4lQSNiA9NuWhRD+m/TpxRoUNk+v1RF9YmzgEPziV3Dh6eYoueUKHbNrBRSovVn7
fe4Rky4DPUos86tlnNgSIRpQ6SfRcqQpwqTP6lnmOAddjaCn3X22GzHYxu3Zbmi2rhCqX48qLLjq
abIiC4HZDjvD+AhUVkG5k6TM9Vl4tkFrIo04NPpuLARb9Z+jf6cXDuKdercUAxjbO4SLKB+822aj
ftxZTyAos0QTEVFFY+l+4gQgX34juMmdEMn7n1uFsnRzb4PB4BeRukttVb8tXmPbBDARyYiev5vK
G44QIsM0KMaqIc8s1d9FVpmOx+7+YlKHu36viCpTvhCjjWDLViPCyzD6KxHKWHqOK+lTUjtgomxZ
EkvPVkiCCnBcM3Vw9oxhwkPnkYR17RRvVRR38V5CRJ6iazzybJH9Ao6c8OqkuYpd7fW7OAbGov5p
Q2llX+1Psk3zKtbwDNXPzDq0EF+kA1Mi8CmootrNKlQMBf/fvZeFWz0Qs6N124+2zKaR8ErrfXly
imFqUL4eAHm2emHqg4VpQl6FuOdQeor6UYBhkr929A/TLZrhp3Ny/APPyRlmv/MQke/5IrTe21W2
/0O0462LXBsmj0uk6a5839RWOzm/Zz+Y1dS9upDmHcM4Y99r4UhYI7c8MxqJvMgcanz99Adxq6EO
LG+aYkraFFT2WZ8upmfH9E4Lzghn1LQUjxAPrX6aiqLNoYwKexRaqAXp3qNY+6ZtPLdTEzUPl7km
I3EqChkLzPnXwdevRFZm3YMib6aqnjKpmdFH3ohiRSbDVIqpQt2QphzVoauOrlUMk+Sp0qukM2Hr
b72haQg2pLgrKJcCo1gsnTtOxGMZZDsR3jOxvBdKl1AjOMd7AfaxnHGko7kVS1t5DaQTsK7Zqlz/
bCHr4b4JSouZIRhAiDeZv3+E9GoIq9NkM37xXX3Llqd2RxRktZSGME8W7+Avs9hPiuULY8IL3hoG
i5qrT23+XcdXI6K6SLikJ5lCDs0ZprlaFN8cJluhPBbCZnAe/JUR7VyRtTYk9YYdGjpG7ni1htEZ
2wMJrshAtRQ8z/bxHWw5FykePFbrl3L0ES6hsZxgGZr3gwRKH9a8NwyFmU1SPDbYS+MbM114YY6O
dZFSW8HRTlVjTY3dJ/XExMfNMcdR/GTZyNsIBiqbwOAGd4FWdTs7DKqoLoqYQcGqlR83MMw0VSwY
NsRxUbA2D4rxeu6mI5mt23DP3QfSSj8Cu7PCtqic/205NznWfg4xkRTpDKCip9uHXfhj/baiGVWA
ccj78iqvDzRNNpQIncbedZm9GzChCA/RR/2UC4w867ZXp+QvoVSaxJsj6USN7z7MYqvYLCmcNg6A
WbFTSuzYVgiUaQMOeF6UjLQC13SdMLSAq2lH6QKN3tbdJzAMjAPlzFux+HLcaRSUC9G3riGMe1lH
7/08WjLkP/Y5vbekPRNQfYIvUmI0+Hrhmvzx2e4yVbZoWzLv+MFB53GcGSEMsC1kQOg8j3yFhIXe
cabjTYEa3CSJdokneoRxAarMx/UxanFJ1jCggyEL3VtkHP72OqqeJODgywWb3u3QK9ZptlrxYMnv
kJSiINWQXVSDKmH+FVPTUWhCMvVNxloxJTHTNaLciZHpimmSQa5h+2jXdm8koLnpF4s+ziJgH+l0
v+besM4V8zuYygY7Q11MCjXU709TTeC+h8bQEHoG0KEKHtOi860FYBkLbdtSTemH3YD3BJeJVa1o
/4ISYzflmCVS/xZUwmUlsvRnFHJk7imGFu7GNku0yLSusH2Bs2sir0pTdJm/WmhpJCiETTOCyytR
e4jXNJ+T5Gu8q9E6pgSj9T6VH65TRzxWHfw7vX5g+qE0tLUhErjb0QQKwoMxFG3urLlBfYCE0pbG
rDnWL4pskv2+h1GevNGep5ZdglhuTUwzgInON4rmkdHyZxoI+OGRAXXuPhqtIE1gEQgvfZZQRUgj
BJlL2ntBtwXYjVgpw97+nfia9eZpTsAVoSNtNr5DdCFdD6D9AqPkapQC3FgCKGUCKnANbmToq93R
TDWt8wBsX1ASX+lOgp5DDYtOpUdyHXDkoUhuTngpoly0UQnYNVO7sKBszcNdng4iaKYDXtuBEw4i
l4Iq9b3LTWZ/04xvUcVXN4RqojbDb/4eNlcR/ILS80agif3mTbLlL5EUxFMr0sOlXaSB3/lKhJ77
XeTJ17hgWgHM/d9ketY/nL/SrLPhQH8VV+RQfEbsIeSS46izlmvErFiak1MLRRrIhKY5G6Le4+Jk
nwM3iBGF0vCIND/w7tiXmHqIZPHoJc/072VFqGFu88g0jqqQ9pOGuLvMENRjgIDiO3cqKUTFCS9X
JDsLqrxtZNwpeK1OdqaQrky1AzmKRIpmBLKTjakbFiai6gQ+plOy+lTTVekjR5MfvP8dm7kXmmwk
2p4WPcSGxS/nbEWhcsm4JLh9z70P09apcn3k0nfSyiKsf4cZZsQOYxlErko0qC9X4v7tHGmy57Rh
cTMn/YbmCNJXkihPbvv2CCNcejKTch60CJ1gsGD1m6AtseLPNPRlAJALva2DR6OdYfeDvn/Hbg8v
KAQ3/ny1DysawZVDcdsHmE293K5J9Y05Nv1j6jhV/YWs822cEs6KGRQC4DBrY1jzcmVqKnCefrsh
ck5eSCLzKTdGyV5uV555S9C/q2YOFbSEr9CrN4xoUKtsm7O4QqDeuSziwSjsqEr2hrsDi6AYJmQ5
6QDXlrprW0CETqG4qv5lRsA93m2Edwmkc+qeHgTSuJfH1X9a437wWkQCQedxRDDeNDrd2CBeumuG
qhiGWGI9Alxww4clLr8DOl0San6UwGS0RgPHcpV/FlNk2ewk6Lgy8iO+RhQF6KR4+p0N+vqflXdI
RHEI/fAXGLfnyU9eQsJa2kD339N61sZIvfZC4vAFEdSORKTTYIH+WfKEeXLS7xLWsKUJMWpMmj/H
oTHwdxL/riDkecppt6P0+JSWJS8ofKfagvf6Gmya12g/1OxAugjYlWbiU5vAuaXQKsPtRGrDIuSI
EZmLAGO0CLSwt398nC0SPzLnZ4x0+BE0MgqEB7HKU4I1dPqbWVRUCXr3JrLobUHmdoCY4yDAw2gG
VzykG9thf//DoxPEjRzSgXVZeScHcje9jLMEKfVTzKO6iJMvjO7Q8Y2ZKh10IHU7+UTFVlnNvH8d
gB+DM6/a0pyPbH6JPboI4xd0mX7mqGylfjACUyiUowfFxBOGThRno2VmB5eogj1JdkSIGSEGdqr5
4VPzkgPZRzE+6jzZctBvv1sZeq4kaVAehwhnQM/iCpL4AZtGgZ+DQnBXUnvnrBtnPpPMSEko/rFE
XJTMg8qsQ/X+c0dkhbYAC0euikoHCx0bWSSiqU2CP0YsTFrPCIBa+q0DOlroMAxBon3idQDkG/Ea
eNUifMp2taVcISMhJNB6kcue8xOI1oUk9jwBzVKp5QMrTUmK+OiB1oF3jjrwu8cKblYVPaAfRyw1
ZASJ1FhBkczAUVWCk0fJwoEnpoIv4owEtXHCt7YmQyK+9mGO+8Mi0yhtReR/QVZbj0sdJ+eLfypc
PFRKkj5utXx2rAM+a/6/jlQsGp8Nis7jLLdSwSEy5YBOBW1yj8u2hIKeVAlG8FXcQjI/p88XF1/T
QPmCtBYVynt7Q0XWoZQVQy961lxiV3MesPnzkIoRJjRdLehOQKbTDlmbd1l1KKXdltW/YJ6kfXfC
szqXzTBptCV9+i8V6t70HTPlqSizHf47bhDiJ+w4JzWUAkjf1VHAOKG8p5j2unLPnwn9ujemIcVC
pzJOIb7B6nEkX0U7jqpBqIz3dcbMDyas+OvCsckoftC+eTRJLgnFO49T9lP7fez0SBT5iISzWrjQ
1WlDsTykMD63ivxaAF0hluQHTOwS8VYZSeaZ49/0Jdwdq1qyty4uas8HDiPI3Xm5Ug7c8EuGyPgE
Z7LDUQC8UkZHuBOlKDTtznNqZ0M5ZeVNsUMzdjBWtQI9qTDG2pcgu+1VETKob4MwhOUQ2Oliem8/
qJm5/TBufao8gGQbUxb8JfrdHvUzgg0tgpk6D+gThTiriischHG4Ct5TsvdBjJvos6164CD2llMg
z9NYFfmdGiKECuWauJfqnNhJfeG3SGrzYaVlm8yGe97t7n7dcUjzoitIG7sV7jRr+IDtAbNioq83
hOblKB56SYL+L26gvt4ZoRG0Wv1K1hhumT41Ltpr9NrQiOIJPXrGfW8HQ3CDGdY4IlulsVaANRt/
PNBsvbUNRl69DP6SPEjYD3dMRke4wnQZAPkrEfbXnXt4a51GRIGtatfQTpEtZ0Z36UGxKe+jWczl
PcIlqklb9modEk5+dGA4lca01Kxa1zv3RWVGJg3m7wLkJs28ew+nBLxKfwwWuUSVCJsJKqvfQShL
TXNM4aoVKqPiFNINVaC2bIJpoKgzngOPtmiZXB80l1QUSGoYtU8t/G4YGOlgl9BRkrkwqooDYvl8
4tEZC++RD5A5XYDjNdTAEe1b/nbVtdOw74J37X9b7wZGvQf6lF93xW69q+xFBMOic/jkixec01bL
wkgvkM8c85BOnanU0UEIvS7WwosVHhxTP3DRusJkNe0ZDFhMCEaTY3aoyTQLT2PCOi5nRkURM1i0
gR7F0JsuHtEaz2+KnYiINSUfDaScglPwAb7stZ2CBH3ajw4iMLj8+a/GZrs83XwxtLa3h3hOUepe
mtva2wdO3cPSqda3vt1mOGk8ZLx2QLNnijG/7PWQFSCaVt5cHS/fHxDjTr70BWqUDNNKOcW47J5I
/21MaraXXxIRBvueCvCy/MEJxlhkWElUCurmfR3RPD81PD6eXDc4yc8DJ5iXml7rlwE1Vv2nBWDE
zkDE0lCJFHeSswz5X3kPCKKNochFZ3csTVim6PZx/gkCeU8AJyGUxhtThcF0iDVW+ihXzP7PIqgI
yN9R9An8Ge1dj8Z2gPeSSBhoOvzognJhlOsQtgKyPZ8Btb/2wfv/wa/Wy+OIWC9f5QJO94kV6nzk
+rNV8JogwuUnHHejbFjOOglm7yBymFTWdklaywu0b8Hyyk6tYhUUVdba1bw9S8xbz8zAWnQW2IyJ
bo8smbvBqYUyzcgsEj6J/tK4yR9Ct8iLiflUHx3jS4ooFJY07zNzxbZ/qFKxS93Jei1UVX4Hs1Fr
XAAo8PkWLsM0FQMlx/twwTYqhk+sUcy9MHnDHfEIA/rJvM5jjgZmCJvwJdc9zCI7/7S/quTmgWnC
KjGkl/G7iy6twvV86JNOzAzF6GexJ+ewxYWTcnMwbsfznLseCtgutEQpirCdagE/AgQQJC5tgg20
AX42d+0IManesMClSrsByRBPbnLwrrlvd7oLE6RmHYXDdGWZUW9QFKD/Ym0XB/qCnO+P2RnuI20/
8SD/cN74GRTjLDVXBO1kjjkgs+iQPnJLQAoRpE521/kOcNIIEe4S9siA6JOVr7nVA73tztgcuEos
MktVEooDyzKenFfsj3mCXWypRbpG84t8182A9N+0xbREFjivdzr2i+VuuMnUOsV9gWWpvOYFMcoh
xUHPJ1vmB4eWAlBRkPot76dWlM+3KJM9asoPiqVq/nOfp09HcQi5A1/yM5eSk5M5IdgB3nPz4XUe
1GWjBIhp2uk4i1ODmHEmOuCAw0RslwF5uaOxwLcefUfblQIfa1uHTKIjYA8ItICZQN3Ou3GeusJz
wbzlE83+6uPIMrok3S9Qd7ShREOaW1ZaDBk5bg5G8rhvMAYICB6JpeJ5Ptxg/89ItJESL1A6+38C
+lM1o+YozhgbLAnbxSv3M3N1RbZ6gwOuzOW2SLsBOo7/UJsT3JBovD/5hJTW5kUM4wibz/LJzhGC
geX4k0NXEl8LAe1OYrcqb3TujufbeVCNvMkXXzXWi8rtjFH3M8rlG18Wi1dqZQoIZgc4ufOtioco
Rl1up2ULjq8kV2WVu4m6JmM05rye5IcoUUGH48BEARfgQaJC7RFpz/DToE52wJ58Z90COyyk4V5A
aQ0AAeTv9kv/1M6suFR1fR9Gsi5UPzkSizIFsiQClAOhqwM1zGej9GWIOK0qIniFJcsxKOPIS4UN
ecq13DautfUnRa/3OW5z6MD6ecLreIHaZcMwgTXSvmnLOzfWO1A5q/hKnlzId7offuQnwk+RKuN2
+QDpkI2m0TTI/bxlIYDHIXQtiskhZEufN7Xm+y6VNRctrvfOQNIQgGbv8KAjIxBR+wxMe5i8AzdP
734Iq6+Oe5cV32YWJNaPTGPJYrJvlIezSrAvKqYgyu/gNzW+luwJNmWY9X31LNKPIW0iO+e6ebtt
z/UPPukKgaI6XvCzJZRIGhiELDlig4BxkIK8x6gP85d9la6GsLZ2RnkXgwfcQS91neGJJoxhKDJn
UDOOzDV7SPr/0nQ5xtLoDbNDina+TrobJQ2iZINWoJBl7q0azos0v3pwWe2y8TPbQi/PPSoB686t
BJYFe5Nj4ACFj/DpvWFojMF61HmAYjgJfpz41lY1moZFAtNKUyUIqruxr+jmwJ8SuK7A+rpvOAM4
FazO4kLrdKoq9uHb2Fn85YJbjCBKrMI5NYW53BydRn8OdCzeTxcPvhmA44qXgyoe4uj0hDQunI2F
/BiNqLYQyQIc2mGpvVQ6oU2jFhsEx/MUQsUfeNxwm2XVcjh3WqK1mjMS3yOa3HC8CVrnaFedykmp
yLLmY9V5qYvhrQH2p3tdmnuKrcymSQ+c4S6Ypl2riqhztww50F5ULXuWagVUNOFdDk3IWiZOyKvE
cTDiSIrOou6eK9nFiSoryDvnqfi3KXbSip9kJ9RUHlmbX3KV/E/9sXjA3hBcQGCBI0QzzOTOTkBH
BIj40emaBBlNNt3XeUczWZhK1kIvDUxx/aOw0KX2NuDT1wC4z27zkeOcyP8fnXy+eMQvnPp2mkY8
UiZYBExPUmxZbJ5dp+kp1d6v2rDW9lfDZHOazIIWX1M3N9E/Bab5njRIGc2FAIYsPJXmk+c4XREK
73QZDdWImToU0VC+Nrcs4OBiijbMlv5RS3rHaRB/M1abiGnbb0wsffy9gNsmmDzYwHz3lbkbwn6p
RCSmF5KMn9lT1CRVBL4T6vJVuuLg0dXPjdSTQlu7auiR+JSZu4fQecNfiTWOkL1AC+ZiaXmmpA0M
8wi5qgCb8qgkjc8hvaMOqWkYniS53B+tyzWX3AevPEFlQnBf1AyTwA5beWUhk3YJW6nbUOGS14fL
LK9WlFAcJlPPSvlxVsaFLTIoHd342M6KGiC54jdF8Bp3BdegsXdOhCI4DvIQikMradqQiDPdWCo3
qR9ICmQbdbTtnZbl1zrGcamCT9qgqRkjbQykNaqxhKblOGzfaXWmoEMOT6Np6m9kmhdeE++hk2b0
R+L6VeBa5qIah1LLu0h7j6EYQIZ1K0YFeCLU9+LouxGx/2CAMlB045omLxP7+ixo535yhAhlQQi8
QqQlJCZ11avMJB8Fsb390ZDWqB30tGtuUbtVZ1TDJ3eU5/UuzFqvhVI8me0DDCYBy8JxTbVDq+AC
bX40aN7vHAk8sd0LIq2kPDjNIzv4jqBY2I4JM7WdhqpAqGI3G71y8UNrkG+707fpcA4NmhZb3oJJ
Da07UAXRTisXyJTcD61VQEnnhjCAs9cvXAPw29/tMe3Gf/H1hS9ayAR2yVkI3PJFmuepUOwPa33Y
/+aU16+MmdIFUTEO5MUqrSAEh4vlG3EMtae7EzrUYxosflslaTduvPJCcvplleQLeDppAAy1saUM
n2cxJdRoAyZvtWx7nVp9SS34u6uJaniCIMOr6zhF9ac+akIqK3I0SCmYT5ZAg2xsxZwdkJ+olnPQ
P0qCBpp+y3NdZbnWBxX7MSZQoR1M3ImhoALgm+HhK5pMV1UEAA9p9p9stsHpkaAWfbulfGmEUyFL
NLSt0DPlBE2Jo1LSGc79iLmm1JgYVJZhG6hj9Sh/ygLPzT0R0E9k1McJwg0uSrTZP/er32QdYKKc
sZS9brn3nzm1ALNO9G+baUO0pqlQX4c5sqn+sgf/zUdrTAXaWPtPVjS+Rx/HHBGBcKNGYqIa4Kxn
iYiKheHOJxSMVx/GCAgI+IyoqbvjBcu3bYIr7Maf9GBdfvfAuh9ngQ1D3n0QWfQ0NYRcMBxg0xzA
rQVAsegRz81hmV0MJBa8xXL9rTHwdtnG44Xyr82JosYS7GCnod7moEytNG35OW4H5WOHLQYDEdMJ
krq/06LJz7LZYf79aepOrxXLmxEzzT61xcJfdpmsvzPAwhD4x7Gg5QEvJtkU7l8piiQSVNt+bYnq
Girj7OcE+fi00LajYzE9kKa+MLBbCUGXharqtvPXmbVoiocgghRju9+MMG/6CaohppIpIZHbA9tE
ECCx0mTomGoAuKKjcwm9sUQjYSrvkGVWpp/sLBBtyP/zIkk1tUSJbM9A+wEOyNzQ7AsAK46fAZ/c
kPmQhgYvxR9FhrQ3FIAowILmoOZn68O4XkNXBI8FFoAiqIW5YatW6y8+E7noEDC8TaFUaTnfDpqS
BxvF81exIS/Pmx42XuBBz7sT6A3Ykv6fEDbCZAY6c3T+qBlDMbkv7ZUmCFICzW63zrTVzgqgIWIZ
dPMUABiQNjHsAry0WKnSVWOwtDMWGtQLYMCltTC9gCRs45ymftffoGEJmlVWlBFU3Ol8nhWJ5ksb
ThKGRU7WdWCn6Yfk17nDuxqpr5Ih0TkyGX/KBvvwL0y0tJOo1pMQPnGWqWYg7SV0WUXXNSq2eXmm
oiyVzzMk6wsV9dxuRwAXbj1O3RBKqAiF+1HA2u0KXbh5hlNcjXgrCVpBvs1L5bFZlBoUnHDgt/WV
6e3zRxBfDiA2DCxGNt8kXKhnY7U5djSrP8ll4Fnxka+XtgFqWmsh0YaCnF1uALHkOcglBD4nDm6U
9NchOOg2a2Ah1yrUTq3yPGJH/KhduQXMa/0or4sl6ZM1XqSlRtpmFvwdIn5D5ctgwCSbHaBsNi1D
d2VzcawvGpB6U1qj427UPSR4IKONEBZewuaF5wKz2ZNKRii9AxeWpGfO2j7vxUlofW5lcarzFMxu
H11nBmuGLWG4WbPdJ+uZH4iaQ4yDcTcnAkBms1NdaO9vT5rJ7ouEZPFBRqqqq1MFKyJA5VZWdCks
jpp4mA5qKKBsxM++GTYV+wIO0IaE7ruHlYsUhpFqOovrWZe+c5MLS4n6n2MD+BBeqSOfzQ+SPbCM
jI3yZON4tQ4FMTK38+oCgyf9cRPtGAAeQE5YMvZbbFjJylfS2bcuV+xOYi61Yh+9YuPP5Y/zuaND
gEMOvfInCcNdDGxhTFhupRqufNHRTUxC15YL+M927ZTYLv8Pcy4XsHitWq4DS/cnsbpWnAoYWkmr
I75JXzHDzVFl97Xclc24hyvAMsJhhD5Y+nff5us1DarkhLMvdhRaDjOUkeU0VS0JkkvQwJe71V4O
rjTBYOT4xGXybOoLIuLZ1dZ+/rSAv4BUTnhX3xojfMCRkW1+SzUkr8s9Z6aNy2iYAuDadXrgfurC
IZ0NlIYv0p3y5JFwF4BxnUwd+w3fZ/Cw3BQ+5zW2yURQ605bd/C9ElaQ7555joNCtznficnK3i3W
cGXHTY7bTeWcjFD9Y3aum9xGS8MNN6DDFJBtdN8bZ0x74u1OYdkFubtEJC7sDIW55LQyTfEHiLLK
AqMPjZMrv6GBAy3Y5Ri0vRtvYKgRSV0DZdeF+HZXSf2EKdjThYWbDRsl/JAm1opzzuJiHrLFAX8A
58hb09OpnPi0SrgE92xvRMWNuowL1xDHVEEDwyjaNe/P96SHgHWPxL5zoIVB5Cz8uiI3gtp2a1xO
sU5CITR2KWLU0j1r1IZYj03XlOrfrC4cR4VS+2epwX/91k06u9ucFTlikmTW81NzKo2XxTVNh7DZ
R1Rl3wYQS12ubiylEB8i7JOZ+Xpl2MvmcbEGypPZvbilo2Mh751BsULYl9NufXa5U2sMzgHn/U5a
gwvI3EWarimuzEP864eKepBr0ZvE+cuAjDE5i97OtKK7cx2v590opAg1L2VULNfa1h0jcBm0yDHN
FyhHyylkfSoQhYVQmuwGENbbZpcsGvYE6ioDimLebByHV6TEXSlnrV+yhKDo+6YMBQWYqInFe0mT
izu0uBdEUD3q+Hh9Xdetr4jdonupdgkTfX/9spqC7MnJrNYZGsVYXyCFY7m+ETkqExVTIbKuyump
vumz/dA/GgdwwgvpBMnOx1CYTd8edQV17sAwm1xwHNxBQomzcg25T5mdEAiBGiQUoo+5IWN+QCPt
oE0Lr3UYjfNm9o13nl8durolScA4VSJimSS0UFjvNG5INyLjbznE50h/c1lsDYKiWfst5s3c74vD
75kK++NX9t8r0Cx2UTvGUXYFpmYBVcgBOuivNG4bkw5Q8sPnGMzrLxIExY+ayvZmIjsLqDl2YrsE
iFbJrdyFiIo4n6boJuRwoy5Dus3k2+3n8NHCeJBUgcKh4tSWbX7Jlk+PbqaMgdDs1760eILFG2nF
fsGpoLdZsTXbGNDCaRjczp29rw4gs+6yy++RQzTWdooZAKl+wx59Q1B9MjwXgcZrmDxZEJstlMM8
cvahjQxw6H5jjor5VFvaa9qXTCFqJ5wdeLa5LgUUbGrQ6KsX1jsu50r/OQ4GrEKQf7gIzmLK7kya
2US8n4m2uJyesKYWdiJde3N2s2A7r8ZwIScbK0Tvs4eKUp2h+Iq3FK65jxFo+OXIzpzDJCI8x61a
ZqNzOtDCXR9XsZnae9WIxvzZFhKjkMmwzJc0boI+2ciszGWMkcjqKxU/dWnYwktxfr5hZC9CQY/f
NDrwagJ4I4LpiCt1qGB9y83Y9yUtQsASojUQ6rvDI9RgUyY5sdaw5OvD34shGbOOPNvdSt0aP9sg
UQdF+L9uZWDsMk9GYp3YFj2ooYUuGz6SF49gcr0bH2tSIephgq4U4KNcqAGacFmTnEMpgZE8/A+9
ehBZjzMn2+1rY2Wu7pDGnb8HXYHUyx5femR0f9owJGe3Ji6UNssMyl1DJrpNOSvbt9jGgorRp3K0
L/ZZGwUw6MYBUyjkRyu+NcJCgw+y/muLdPnJ8UWEZzFzNLr1a7dpUGWB4h/FGWwp0kYGR99NIlWW
EdueZnLuX69T/rdDDKrC6c3r/xVPoMdPerVJBApPgjoAWIc/rOgS6MSEaN0UMEuZPVIi/L3FIu2e
KdEzCMRgur3ls1EjkEhz0JI5dOG2gpbQLAus4GkfTZfJ9AQNx1zFceiRTlPFYlCGo5XFurq3bpe9
DD3Tf7p4lOJHlgNcqgUhZD0nXAKirUo78HdaBYQ5blqxONtOhGHaghvK8fgsDrLC0DUCRgvz/3A0
2eyzV7YqC8nyX6VFzBRHDT0S+bsqf6ZTWqG08r04exiqvR6gNpgOAXqSIVx9TvxOQgIfEzO97CiG
4abALykPecHmQcq1ciz5cp+VctPbfdI1nENNRqbCZ+CUwM39IbJSxcgYJbm0GqewYJMBGd37dnwL
HbkHA/Zcp7ZiuAzofh3HIIeu8+0uGtoDeC1+GVs/tHuPmjIOQNBLy0F3bZ9qVfWxasbbTPllgiRO
eC7yIAthPpv6QPb5559K/Ez3zkM+cCTpzQKEoQED30xsOdgLXw8BJLSEjPKs6ARsDj0RSIbpDKzD
DWebFnVmTyj6hQwdEMM6PBM9GW5L+UE6s3g9QL85TYK6YjkiI86KcKdundwc/sW8B3MwgY8cLXbb
0njtiDhWxyz/75/Yuu7WKwBZi9GORc+jjyTW13YqYo6JtUj83Ho0OnyWV8kiDONc+NL4S28T21q9
amJ9ZUj1EJ06SV5zXqZGfvdP3Jn0Yg3CUKEBDkIdIjGPC26lJ1rPPVsq6Uh97cqnAQI97MnuVarb
o1tpcFGwG73gmH2KhHzJNcq4Li2fG95uem7qRHfWbky2rOP5OEYnAIXX2TK+fV3nXMeuYhJWjVBT
3Xu5a4gZ0ScUSHrwkktXVNeeYWlLL6dIPZIib7ujItUD6nbxbQSDx09/pdtKQQko33qt7hnk/sCM
Soqh0J/U4XwwfCaVEfl1p5UYUhz3tnjgrpomkhXkoo/0wjMj0cI9rWxwOtq48CD+mR/1TkVBn1W9
p34BnK0D+chH93eZhgTaNqeSY1DvJLo6Qi3tvPxES4CGvwQG6APpnXJMEgwBRmLHbwFkUPnrkome
PSwQ67F1IUeH3iqNCqD7Saf4N/rNSkllQlAPNsMeVCUddUug2BObabVeQHiyKB4syEwMgbX8Zlm+
wpnENaOnHb3Kdt/WbyqZ8IFTV2R38PkiV4DkJ9yU1GBFsH8CpaqoW/fHGg9CLePJ7Wx8gWpkqe5w
snFxsVF2JfgY9a/xwqAMdaT+/KDUkAC5gxCP8869bbqCI8M0UODLJufgMBKOLsnKYPfsl5errUM7
046g+KXmR+xeP0ZgLO4WCmFXjgAaRw3qXH0wu5ndK2t2uhL0BwHfP6yelfKf5OLkZmhiu6jpt6wM
y38AKdsFV1Ujy452ig8Ww/wJVwTm0xYcLH3aNVgh5LV742b8f61H1a3Sg5yjBPSS7McWyvOh1WR9
LGd0ea+9DwZ15TQ2bylQg/AThSqtNWgBHRpqyIWPxlLu2IzFwKbzDLVwRDsy/sHJj0gtZu1uoaU2
J0XUShveD/yItQXlV+78onfkd0HYV/pZ6yNhUQTLk5v5pIPEXH9AxYmeMT7M2G7pzT939gXlIExu
6/mkf9GKnZhwkos+ZGA667Asw71S9yc/66gw0LdZAyKG8lxzVHlQYb398woItN6Z17ofYwOKKrAS
Zd2nC0XZaXWo+E7LLwFjIBthc3sw5F+Yj/glX2um66oAuJCgt+MrwmkypM0MtkjKOg4U+qTgdfpa
srcVi6A4mN+d64ECJMDyOAFV3BRBFAFm7YmvkeVkmjJ462YMGOi8frMZDa2Wm7+VE0iZsBWmqPSJ
1UQG0bBlkmETBUAizNgstI3jVXSUVntSWVOOnFq2rLvHXZT8DXjEhnucg3foUHT7B3dK5w2oYYjy
uBil8oTyxdFDNbOpejxx6oESDQie9JUTBlazfk57UimbRq6SjIdNOjm+pKmDhdQ4Bm6WbdWgV/f8
JBNbmaI2IN2VfB9RVly/XLKlOiRcX6/BFNB4kNNyWWEmeIBG5M7XkSEYluWelBpwk2aIec7jcdT4
rlAKCN9Eh8cexlfxEp9g58Lf9RLsrdjY1LSspCi0tWxbX2u7CeVjwleFavK7qhMYwlUReraIyO1w
CSv0amlHMoBhhYYvPcaZ7T24czpPBQJi4tG9rY5bBqL8RZHPze5h6IQvzNCQy7KGOXNK2DsPaJjU
sg==
`protect end_protected

