

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mCyyeqqjg5/0TkdJEsEEwiyDfrhah9gG0fpTMwUWGOKZ3he/dpUva8HsS4xtl5XP9zdNgeOXA7QE
z8wIFX99RA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X35C+3C9De7vC0qODnacg9gsvk+3IzrNpqQYzh787Czr0LrIg4SN4n42C6CPfkCBLDXSXwC/eOXr
yWqN/Hj/SYBmrS5kjeF37AKShalo68kYRaZgUNEiNvBgjtaJt6WRpWYojbh+ogFdK3xIXCNq+Qxl
K0+QDwwSCDU/YMofxGE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n73jcH3HYbuczKsWgG6ox7VZK1YnHzJQ1B4KxEg4B/kZylbLOe/lb0i8/kn+CjmMlUuMK0WQWfed
hITAZaScEDQ3B6jcHH/bNliHMpa5PCxNetq1i73KuqIUSMzdaxGWTSuFoXR94e0GNel9SANUqOYF
vTOS9qeLaefJfWuMi23yYpmliTIg3f3fAbSdeAfef4vuNm+0XcFw60RpJQs3nrsFq9KW/GfqXw4u
TZNQUQbt6cL25X91FZ9ygQq3zmgha+CzhVMH2888hx1Tg3YKoHcpCHNpnuDfIIlbv8c/WTDMb67v
IK74ph/GlcH+s638TtetKCgz1jniP6o8owuM0w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lgEz+Sb20/Syw0As3tLsdRmvucviIYGeDJylwgde+NWKzNiVP+by1Maor4kKAxxHjnI5lkH0wLYs
PhqSC4UmzjejXWlU17tjRxtRz6BbrpAi6gmDH8SRbE1L1vIa3LM6opScw2kIKRT06DZ3npJLvb1L
GQYpSvbMBpeOoeXBKyg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cuBsFlva1Z5u1UA+GZT5hw/3RJ+t4o7i70J4gtLUlv3Ik7QI7QGdbqQ4mg46AQCjs/XyJI5tDPDQ
SIWqonbFU6W95Sa+82Fm2FOLny1XsFw2bfUdFeJCVtBal0R28pkG/kXPwJRvcecEIrS2a1k5PBE5
sZrJ66qcp7DI4wbfzpv3ic5F22QlsAxZqXZEB6lBkhSRHmx8sxDYGL3gz3qyqFuTzoFlxGj0D2l1
7IJKcs+gQikUKNCj4QKZQHmP0x55BD7tR2tDFNHuJwLQeErQDiAmIcwGhliqTf1RxwWpWFh5JUyZ
nisNHaWXl8SFhFbWbHjUNb33VdqRqkyTz+gZkw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49408)
`protect data_block
eYrelQeTTxdKJN3Jaa7YcfWciB5o3lM/3xGKEBNB6C8ttos6lt6QCQRy+xJD6wxylDt2hgxLoaZQ
ePKrWa3Fzu6nfJHuSvL8TA/0/t9wjEGus8BotkvG6gSp9KGCM/Qt0ujET8ZmyxxTFJpDb7mRb3l7
9YDJUf38Z/GQqsiZbRW9QIS3fTUjof8+CcqazPeWn8KvzdYIKiAsP+/dXPr1BfaTEC16JrxXq8Fe
O/CqpGbFVkg+oPcvwYhz80aH3AsJSvOPJ7/wilzAwymaF95AB1fsMlECGxzfFbbfUJ3jM2TiIew5
sMyGkE+LQuyuRijzoYqvQw8LrXb7QDR7BrfPPQ/nFTVmx4klG9NycqNXxIWMZLpAmU0y02hpvn6L
sl7nFiHx9PZ9xjXRCD0XYvzjSunyvtkTeGvRuABa29Kh/48HB2MwYizmVoUvIGkh5kqCSa7IhPmM
RCADhLOLISCjVt0qaPLsdDgsJ0JGHrZ558O2AlxmSgNsEVO5CNhifI9VEjLV6VjUilyiWgQi4soq
MyMUz2/B4xvIhrmB3XOLUXN8IJOvhYLw2AcHf6ZLMqsljDcPmLpRO9Y2ltjYcR7mwa/DKrfSyX+j
FAF8RvlMn7rhJqyGgrQJGyEoyLOUfFs9P3L7Pw5GVXggxSpxYqDeeqUIZv+EBoK7yb/mKbT8gjZZ
IGZT1/GnVrZIzni6b24I221QHy71Z6rl6eeDddHatxX4i0MtH4Ipn+gRR1V+xTod/cJa73FibTPb
4WlU3uh1d+RtCNobXDCsSd6gLF97l+mdWIW5cbdMbOVBjjoYpxIfZ0xj0WyTRCr+NS1N4Of+jXgM
rdsSZpNj+hwzEn5x+qsfyZTTCVOvAGxF8IoHnc8Ruj+3Oj7+ilglHeGJyltxhqHv9hCy5Gk5t9X3
QfrMyB40IitbSiTwXmrJsXQKlHXrog7/sn38gCporUylIsGTjj8g4olZy9/3x4rfPi1nDepmgTxc
rP+RVikQYJE0mABh8rYcbhWu+y/a5gdauMbUmEeOOBszYRSJv6ta3BPXvspee1E8LaUhrV93hHHI
3r9gkRm1f7VCEsBpz7XUy0oxYwxhSqywJCn3zVvHj16jH260Hb8cNrBBcdpH2sc2osAQyD/bG0V9
EscSQ/0Pd0RpHe5qDk4x610d44ivLBHGpfskg5NH5fFwaMrN7jRO6YZcoHJHVqzmd2XaBNiQ7IN8
iqmJcKqMDxf0/050Mk+cka6zRodJ53mOwS2M5RJMT0owqSv+wzBd4v2MHtfhRdBAws5YDle1P8IH
lfLpRWJ/wzzGdPjTb4I5F6mGrrqjZT0VtuNDHZV5lplGXWoK+ELfSHtWXP+mpvVHZ/FQqbozfVy4
uBZBpNvCKV7mwqnXso9hKkq+ORILNM35jAUjFYerSp+fV/B3INGZRg94Ymfbdeq8pIsx4BfHbIdn
k+ekEosI1O04rOEC3vsByDYBHcf1tTffQNYJcACPZ0ZDQMFkU7T+0OnGbFlfn054QIjLlFzeDNDu
Lh85yhPCFqEMoUhPerUQzWjBmZRXXrOWrz884kAS+fE15Ehb6JyJJD9ncJF2TYeN9RMuNw0Y9XuB
Q2qbK3vvqJUoY+6Mmvri5uCC7aCfDyEHyofe/HuN97ndjtWiaRSYdg+dJAoiQEZxqp99sWVcmbdX
PvFHLuEs7saf0E8xNc7YTOGzq9EVYfpym+Z37cRGqbpYUfKyryvN+YhzRAC8zPZ/1KCxE5V/4RVD
FW7tg+uTWRuW3QeL31e4NsWtxHomw5B50RAhI4tjtuEXgML1koxDzfQRH9bjYkKBvHDbJreukEp9
aK4C8o+h5RVKWniuVPwNIJ/UYps7nA70nlQzGfmqNM8TI5wLS/P+9fY3k5UauvPPbTpYNV/vdw7E
1W6BztoBl8K3jB0LAwVWGX3ppWLshPyGsVF+VyS8ueyY7Pa1U/I1j404UmlpyNvzcWcFTs3AhnMA
QKetu0U0f0KqADmdtnyL1a9yFrGg+P+oMjZX785er0YBPX6cBlozyiTxDg0M4tPBu2obSoQnV9ot
O/I7bTB4ppPvl8aehF5fqsI1isjmYp9dIFiNq5/HNraFpWyXyxK1IkGn6lrEeGNaE4F8KaZKcElt
skkUwbTY+6bDikHD5fTigjcqQ099GuTwJBBp2O+BKshM4/1DPvsAZUFbGIeFgaWKmXN+G5EnEu/Z
6AdWwE8Bw5CYGaYCauHWDGvLAUCFXsbWGmaNFhfqaxn3L29PplAtz/vrN9lboT4QV9dLu9KpD3Rz
M8ojXqGbqd18LeW8iEm+MKAMplDNcOH8F7hlDIJgwZYa2YMm2Opdm1yQJmNsq8CVB+YnWQAmIQns
6Awhz1TPTftDITtjxKT5qlc7CH/4iMqDRnZAxUardr7Syafq298t0cYU09qEettpmabDlQ1yBFuD
UcO6tboJDeeXR7ESHWZ18K0LzUDiWdlyueIuRu2ldzbqrWXBX2gPPNsTszEnzOA5QD45Gqj52SRP
WvKHR8WpgCIz/MQqPs236Z6xmDZmhSrfPH0oJnWJrip/6NPmNKaX1g2R0+et/RZ2sBxnf7meOrrg
9jILlHDQsc0Bwd/VS7SYN7Mpx6GUximSlLt2r30OC8VANLW8+6RQYSkEvpkHTO7xDO+bySzZp+5j
CVegfus/TZWThgVwHI7H3cLBU+SoWP8GPI4EDeGr0x2diCRhkI4p96hYqAbHRgmuhqXvqoozQblB
AEZrrQ5QhlhvIiEDx1kyOZgdQa31AWD6+7FAK6o9C6DCwESOykO6uQrmZu4ButejJVXQklJh8dgM
qFjrr8CLfzjOIHdYCYxHWZvqoztS8EfJ160ZcFYobQ7/b2Q+s/AdyQ8CGTYHIFBn96fmuB4tEW7o
GkitGvSXhmfxaKyf1jhdTvXEGl5AjxOYwwfBb54ETTRoy14oBoHg5daAqdcblNU0vMllAU+ZWJa8
ULdYa4rhyaFK54RIaEE1vTMoubG9M26Z4WXH90ewdFopZ5l5w5Q4TDOp/BpvnOLT7cdnyz5Flrh2
s3gw4fGTHU+GzQhBem3Sf3Eo8T0/kJ2BKuwd4K2412861SJtR188bkOXUwH5y1P50kiqWc1Pv99M
AoI4JoadGomAFjN9ZZVIjeTCGb/MjVWrvQUbFO01TDGNKtIOQjK3GZAN1A/7jSWCXjOUPBtyScvr
x7gZtReCSPfJA924IFlcc17E2VUNCBhtKR7tTSyeDQUh0uuQ5wGHNfzgQVzA6EpmEj9xsvytWAEF
xzKWYE5c5QyUTNphB+97MIFgXFjSJW/u+J4Yt74uil6A3LKPBBMhVCthWxih2o3ZDFkmtDdRIGod
dfW6s1MPhz+/Y1GjBEImL6OGL/TRD1LrGe05ymjirg+W9jEgV+8lDn4BwVc1G7aF9EwkmkZtfV0e
l/1YazAFAv30IXa16jZh5Xb3PlvBAO4AfzdjRHmGlsMKNz3zelXAvzE4h/MOTuAWrG5gJxbB8J19
tkP6HK89Fxrdpn0jA+BKfGzfa4WpyAwiyWybGE+HRwLLwFkCDlyr5m5ihPzyRXgPFRnw6Hi5GC+w
0IBx4xVnlJuHdatX6lVK2gfpQ+A8jDDsLoORWYYYDNZoQPf7Z0FbzdJdhKAZEgaya45z5gIGHHS+
WouVtWi6QFEv4ey/nX9eRaU+HRDNjR6z46OAkwmwH9AIothK9UdHw9X14LbjVtH1jW5ihbr3IQwJ
rGzk5808JSlCuL+PluZpBlBU6RyS8UV5unBwBShRhK4KLGNmknZGbP35r9sPY5pPpWXsYxpC8hf3
9uEL1pUE5sYZ1q6pe8MM7Jtsw2uKzPftS50IAzBNTE+pOMmqhnl3IiF66dDa/db4ZnnbK/qUN0th
H4Efh4z/SwjdmUuJ0+qrlqIazU1ZU7WUQx50RPuerBJBNzurNYEez2UuRRHTg1uQ35c5robgKPZU
f1meDxgCVmOkt5GDPW4kFFdj2VGWkPbxgpzuDV2qsiglMITNd5g+xed27zDcP+43HYMH9g7niIaX
4geSWpelnGSlzWNZnSmEG47EYRanDAQLheTMC9gCzBn+AAYFkcCEtjtc9ZedGPhIeFE3LHF5w5Cf
99Zr98kVs+PcxDBT9YftAhFyOCJBA+wJBetQDx69nDWMKzv8dQB7WyDBGhubDlDgVrvUqrBLByxK
l5KU1EVwVDptwTEr693ukUgcUvP9iZ/XMVqAt0bU3QP34yZaZl4x9kgQrzDQfa04R6vd2AYVAZt5
tIUglkEx2WzeE3gMPO85Qh60Hg/ry0buPKrEe6T4VZYRbg82b/n4vXykSk47oCng3WkeS5Afwcij
+x/ejlP8u0RtZjeJcfC6QqITuu76r2hcPO1R0Ycbd4eiwoKN1I+cPwaxaIhzYsmdwEd/HvfsQtS5
ghJmcFO7BHUohBl4UDSOpDsiIsc1He+PQU5TzVZbGtd6EAzVMX+AqDAYx11Q6sDwRUZ9JzzOvwRL
NQzGg4zDkh09K5wbjP5FqKyrwrIgqSlfA6gnmAwPkkCnzQoEROWEvuwCfp4a+qA0y7lsYX9K4UZe
JrkBFeMCsKWi91m5as5P4RoesOhYuM5Yj88meSev0t1H2LoaZOwpwVmiYgZGrzsv/5H2H9By1EiB
CuzR45g59WhUblh8Q+B8uTzadjUoD2wrsTYreEqOvLCDkEQ1ej+/5ZepbVyOgXo937uqt9kKZTUA
48FHAjaAXf0mUj4QEre3V10fjbCisVS/xqejA2ioEI/lfqqrW+1w74BVZ7pD74+X/BERXtMm+5ha
jPE4E2MOz9SbQAF6qt7onhF2rDp1eJ20FvGn/Y9thIVgdOXHLGOppgAYcZ01W3LBLooPZbmvferg
SBFGssu3P827UL6wl0EkI1Dwaemnf8kt+BZ/czRifug10f1GFoUXg6UEZMXqEuhsKoIQ1DAeqgID
vLJunUGVP9LJ2q+5QHflzedi6VXchKUjZgxLma5RGKQdolVjDVwzBTgkNQnvWGJRe8KxLbttbhTE
HnrvmViNXGQk63daHI+Yek20WWnjMALXE87vQ3xXsPhF32d3bQ5+qzdGUNrPVjZfT2zZgkt+3NMQ
tTbf0p8RTuclc5y8NgCWQ/ujM4J+rwVbAnL2DPq9mY/eizW2qu0ZiejcX9BLg55xRDWvtUfAYITV
t4TkzkmpWEUQW1XlsaITI5AGqgw1hRyLx4umKb58JEJATxAh5uLAgWTW067Qjhfz47nLPZapRdZc
n/F2Q4xWyhI5xjWi9pgyJzmtBraNxyGbkc1dP6RJ7c0/+NGh6/h6PcABO4LtGzYMMPG4DMtHsPjB
BCJ6BPifN6DJE+9gxDeEXFxLZHQ5hkujcb8u3DjqKQGZnMTTjG8AXfwVKZsdSNaiQhs3PIbwoIKG
NaJi7l2pqX7bhmIgDhEo+3MtKUUmNNCp6nJQAlarzP48sL2jpHRcF7vQBteu76OR2mM7Gq41Ynas
m55f44JYR1rb8q7efgzz2Rg1yU9QCUEpZjxCj3npTC97umXcKnhLeTKNw4anEukGt5ytv2uRTXcD
hCDpyyAB5n86DGYVKMRZZdg0K7o7ejULRciq6lzInmylEMK8MRlDZBD0ARjKt8UzGk5eIY74kqt0
C35+cVTtIFNYsuP/hQSZ8hf4bWcYg1fD2YvmoZ59v+kmaZcn738+9Uvk1Gpls/elo2NoMajf3pEJ
gqTCKf/x81Hxy/CCdzCVc48QYX+ECFIgYg5LFp1QWGA0NPc2Nh5qLYeRoAGtE0TmePVweMpNTAYu
sxSW3mVQlG3t9vw0+ni/Gtivg2stvSESjqc4uhVspn5sROxFTywZxNdEHZOoagkT3W8ARbLS1yaM
G2RxiKwhlcHzsP4S5vlXVJU4dBkv1zD36oc7lC1tld3d6YaoDzpqJcGr0Tptmu0mWFkMY4j1xyce
b0c8QLg/2cWkHTjL6spx64REwxE8sRiNjeUl0elQ/4V/xubAbaO+M0t3Bvjo2PXRXXi+qBzW9J3I
AXv8flnpOWS8inRXZKbb4ZjgeOjABtkq8AtERKKqTy2skg3OUm/iecMYnMx6xoLb6TL5PFE410lV
Iu0pbm9H3hNZnEH6qWjpzwrv/LIBWkgldOxpjw3aAPDRGS88MzCTwQLUrcMjDpXqkLELGK2rJ6/7
evGNgvlXohtKswjCXG5UF/RgayngCzaCnlFXA00ZPuauh7Bh5j7kIK237e2JLMnhJk0hHk/XsjrT
Wt8R7Q0iwnRTQIxJ8zYz1NcWpOmTxYh4uKgZBRg0XU69Hp2URKSUqNLr6TQph6aGhOhkUvTlh4+X
DMZ2xyV9E1aSs4RPMee5r/hpuseKpcpMeqatug9SQgZdSea+LXS0vTUaDu0wwzkFHsVn+zup8ovP
kWjTBkD8qwevMcKSrWxcnVK2yG5cCcaRooU22gTLI9VhtbXp0Jr/smnIPf/Fs432nEUyIUVM7yHL
oobFC5OJixRmAjBBXKYYq9aKjlrFQFOIGXQu2dGY+f9hyklgNgVGooZahibJOmRkZRKCjwvya1JI
VoF/FSJ+yiMgZVjalmQ4vHScC1eHRLmy3gEtGT71+4bkWDSpNNCNMfqIjTAlk4f9rlVD2arbmAaN
cK0REt51r9J8ekRvBPgOGGFKrv68lozhfbGm77HjqVmZX7cBffE9++rvjoUGhobFJ4lABP9YRydZ
YAvIJo3mStwyDOIHmW5VULJSoLEVpbX/QY03bx6dWKtHsGnmpkQlTnTG3C20+f7RAC/JoJx2qzmQ
UftgIN5iDRagNC+617uecOT7Y7eaYP9Uheu34rbW8QZBF2sgjXUEEpd+CC4yzQCaFZeJ3kJuvnaS
AttsPIbyNLTSNN+tz9AsznZCzILpYso3T7i9yk249nei0NDoWBeC8/nDn3dUK2JgIWFHGmrEvJcK
XSEam4NdJkebgCAUI127w8WcSmF5bCabfvAr11cSfk0d6PM1yPxGFkBdkI7QM39sO0hn3jmDi2pg
0e7QCTZo0cTsdDzFU6xU2ytVXmVglDKce4u2496T6m0m7HJwq396MNfc5AimmHtaCfci003uxY37
uuTdFcm3QHq35jDJrDkTkwtHeBakZxBi78/BRQbzQD6SeMcL3wmOhFrqDvFRitENTQ9IbfdycCA9
E9cKUKP16C4E2ATbroxEssPL5Stsx5rAUsyPSyyOAxJrq3I5Qa0uVlvT7n1AK1K59iCNZjxittWh
B5PtiWtTdHKDWXqQ7zdZZmC8gds+hi2zpwcJki7Kzf8/bfkmIMBFEiGxs+/Yr9wqNxke23vpg3nh
vJQmmzMitgbRx4zV9icuzI6n+pImMmgvqKR3TBvYUWj64HrBbIyBswayDnBDfZHI/cBfgl9Vaxgy
VrbOhxpW7aiE2rcSpRfJuOfyVvU5kLFSiLU97E1X6DXbMaKK9k8FjdiyMnymonDAEgFvO7FekVet
IxcnQp3r9BmHdTI/GR90H3DQ2kWO+2a2KORwjZ3W1kN0h010syIG4zIX9Ma9YsXBHHl7KaRjIGte
6WjxujKl3Ih56ysF6ptnSc8Jl7m1x+n7/XOkIU6MuOApDzgZWUVXu63XKbl0nA3hz2rU4T0dCqGR
RkiUDen5s9s/SDLKG4ad/GJq5LOTUCwj++lbCG2AdvvGGJkm+Uk6sfYAu+YY+iYKtjAEwy/BHNNI
QmZRsN1g3nm4Tr30lyvo3wXE5bIt+/v8oGXq9/6Wx3GmiS974sQxIMUK19unrGH2QQlaRng0DhSd
cij7IYb4HeaC2mpP3IbIQNnp/H6FSz/cTQPVcV2pA99ShseQ5wGRb/8hFPlyB0bQPTlc0krH1RPX
g3+CbMyG0HE15aBH6zyOMIUlXDoEfqhTCly/tCbCJUTMUhyaFTuxizSB160CFWiF2EA9XZGFAlq6
IPaRW03o3vdw+qPtNWhJdfRTf+YOm0VkV47NyUk+x3jgF0syMjTSPGgLbq1zZF2i0kbkzFbkWQbm
uSRrXqAlGj6bbXYKs2kX/rQu6vYLPxO5WcfyThi9IIQ1qJju1kRCn3+GdhmwoEwAkRqUVFuPOYm2
dhivYVx4qRlJbtIzgb3YN9F9OzW3zM0anEW78lZHmT4X2TeO+hD6ybdiGdwTNRek1zea/Yl1qyeH
73+TEsURbwQ1PYMwq7/7FYO5ciiBy6gq2EVfF9A7KAgLoRdvOKZQrPoGxGVLTd7V5Y2vLZgQdWxM
hi7Fu4ptCd2Diw9i3UZXQEv0Dw7vOI05qQq9GqJrIiPvXe4cf2rNpxGLx38pwNCsBl9mhgj1ex/l
U1OCHb+0pCA0JxxwYAUKoxVWdvvnP6IXNXi5KCP1XJhwQCqWv1QlMIVH1fDo9PWyntcYfJCep2ck
fNBZ6FR5dYgX7aj/aToNgambcF10ppWlZ4hYp+EDsfNHGuHuhlSRjqjPX0wO3LOkp8wfBkBaQevc
c2wucdagRFhbKTOGDrwPR/0DEkKPYQg+Z5OF4pYAhk7IDPcXjBsGfPYwT1ARDp7QiM0ZuCKcB+LK
bIOs0G+JOPwHqO8hxsSy0Z6wMaw0qbR4EQiXk0xCYggXuMULH0hXaDAZI7P14EMpgkI1wkeMxTlC
OBJMQiwcfax0s7PEOULTzdRQU4XvMz34maekwPeuTp1Y+8mvJKIgyQV0GSzO42S3TGZ5uCmgCgqJ
k1uzfBcWTAYOq2j8Zn+oa86GmyEdp6+wcGQdeZfJo1F1OwoZYdpgeMpB6HnUWMuZZ2KCP5o0/suD
tPqLJjC2BZ10rc8mbcVdQOmxbHMJO0UyclyJ54NP8z7zFHUsJV09xTuyEm5rdNrITw01shMCfLTt
MTu9byXC0sDqGaluowUhT1WEBAV3JgxE24sopAnYAlxa+I6dGv/CBLVaVixdW5pNrC+q7cbVw0i/
9x7ehazP5mCEmyENAO92e8Im90jUG6cHi73hKVzrjrNKmJfJyYgReWVAU5yhLOqma/sZZWus1gNr
bIEfRolM8qZncEQcxuNTaZL6NlUUe+C3hEM18+JriHhlPWzMNMlXxS8LjgGvMURc8I5+gFtb3RBS
+Dhw4vtHExydr/bH1NEfzvdBdU1ZFbYZf242+aDbYERumjZeWdVnkxJiAgilb+DbsCYhRehegu/J
247iggLBjcCwhREO6jUKPFo8BXSsvAu2mEnA3i/QN6iPldbmbzs/xkTIFIFZTS3h5m6hYOJkDeJW
xzBpWamMbb+WjjWTZcdrBfiqaHlf1q5CNFf0dyBmdz3ZyVenm1Qewe+8Zpr4MauWuzc3X6URUObK
DzVyoD74uGa+B+wVitwQx/9w8VVGUwDl7b9cAG51iqC3AfmCZ4uzmC+VMqbmzMln4XftbZaoHA0x
/I1dp/F7IXDV79jtYVocGlF3HzWVlijbusvjAfjdbnFijiNbsWM6HvunAC/2XbeLtT17jrKgG+N1
Hu2e5QEz2vVSsThFtfDvId6mcK7rmjKFcKZu/RDiRb/UOXx31Gkh3rhLg3aHeBD7o/vE5rYtk/yc
2Xw07CncENVc2sfTEscDZkC8WeWA5M46hLYjLEOc+R107ggRp05EAuo4YYdquw6OzKCJGUme2Jse
TO82HIdtAyT6wxPHlnHctzrLuycLOiplY41mlG4O2ToZNsYjH67wF5DwfPG8GDbMmv6u+0SXudXg
Ir94f98URu8bYaxwfbS1qI3ylr2TQ9VORC2Flku6bsPc8aWXSpBFJWVS3hDefewyGTahGKhkDE0M
kNaiCNdQmV3Z7Tjll+vLO74QZn1mefV766GM9b3/fwzVvjxHBRNzvQqoJJmR/qvk/O5P1b4X6Tge
GITD/D2jeX5nSGEA5STgtFsaOgRqA6eG8xwZ+5fGRorxa+uswKKuTPPnllwIzUTpzzjtiVN/AwEI
KqmEpcmzwSXf7wnEjwshLbZWYTVok7ESY7PJltTR6wGs1sboSl4CVgP/sBlGWAOu+Kaf+R/CL/eh
nWtX7QMABhA6sCDefuW1KByvoSHAVDVfqVTIa02B7n7scPNt81r/kmuecGxQjCjMulxfEyx/6PsE
nAsTa13JSQ0UhypyH+1JjF9Mbng4LwMRwcpV7AOGHo21lwvsnoOKMkBeLUP6SkR43MnWYRsBrRre
1EVrgv060DLBaFJG9uHT7JoIPFTfmoTaDl9GzpyZf8bu/zcLhVJ9KXAAtdltKMlTErQD8+R7P+wb
02A+CvQif0ZBUvrWmJbUw8GLhFZwuDIL7xdW8rrkqwg32HpMea2v6xNttNpZisvyA0P5Yqs5CJR0
tyUhU8NA/EUmZeBxSbLyX6EgZfWrKvY7BLPq8GO0arwsA3SNeW/oM5BZLmvepPm5N2LaW93a7agW
E85LspMQLeO6ccA0+zvDCp8p7XxKS7QQp6bCdA3tx5oi8qbX7BtQnHaK1JMfrqNt6Ymuv+tdYznU
KDIoy6ZNy79EZjYOOs/6PfbOGRSQubSQw/Fzoqg1zMWKmhMOhpFazz3LrB75RK4GMuuyPTlSJVll
/JbWGa774XKRoytvv06S1UApdazFr61eSLtdPWBDgqxTfjjRDc1bRvR+6FrZqkAr9S6vxiXGdvu3
SqsB/5nhzjya34+sgVfR0PJPHJqsAsokkmmO/vVpy3ll4aUGLbhbWcjgU3SRl2x1tkLmNML2e2lk
0WMrXyDLyyOj41LNuc5Sys7R8sjLXVzcxI36qBxTpl3rCo3bh0Jdiot4/Ls9bszq1azE7VupOrIW
lvKClyiJArDdna50gOQGNcqZrZytq3sT+NuRslfus3ZTGs/qB72cEIgABmNKft0ATBqrkj3KwBI5
yul/p0el9mMpfGKSxj/0od4bGZlr4MW7OdfYnv5od1lDwP/vovl6nZ/QwoMp0rC5iLWNSUwxaG8k
jzu2Zf8HOz/7cdkewIJnaO83hoqenZI4DLwO5VOWZlZ7hQN+DUqLbJYhfVJL6LIEruFeq6EkN6Dv
xTfH+UtDKth0uAYC99oeeqocNUPrnA8LxLqxsEf9E9Z2dOVduSL4i5+aQkIjLUr5FrNeSu48boY9
hUel+47WHCQeoz4YbkEGe9YhnMNRIvbjQ08PzrtdkkSIAnADj963RNUTFnjLu+0MAGZGjBWei+3J
hrTVXXPdOXtQJm1FHU9Jxmu5P7+ZuiWV0y2Siqo1bf8/tTkW7aONl5r/YoJ+YjNILnqHZD8IcwEM
RJgx4Dug40KG1+r91/hSbHtH0ftHPbyELf8YUWDrePs0bkJNuvEO7/jrbErSbQfS2EAvcYz0ywW7
KsIGynOd5C6GPl1ZDKypBQCHyDnn401tk6Q9EhBV1r9zAB+2JPSkishzYHH/89MhGXafbaKlgJWL
f4dJmm0N7deChy5/0u0MqJEJuo9m7YCb497nKLzr3SCZgr6jEMx/8u9u70bafg+zqT76TOjNf5uj
kmaB+MRyvsx2RfwclK4DoS7rz5rjzfq1Yw+Cp1J1cGnBvWWP0v3eyncx4qLts/YsI8Aw6/7fNNyq
2yQGJ4rWLbr94PkodV8sqBb8+Q2J59ibZ7mhc2ZULsL5ObT6bBMDrPmfCf5pnWLvhqsFosmid0oH
m71JnxR51TZTOvEzUty25HDsHnrWqqYCXvNv237ESEnNLbx68M/WY5nhQ+hPD3rjugyPXMsOcHpC
JAxBNaUoA0yCRIGMPJubMMnn0o7wXIogTTRyVZFF+8Xo8hsXkZOkUycIVH5E4v7G12Ixsrdn6j1+
8Z2Ko55X1kTJxcSV+vD8XsAuCXgv98hnKwtw5jOn6JTpXuxCLpWtZ4m76Rx3aiVtUIuIM+doF58t
f3fESt92jbD8w/2PW70M280ZzO13y1tIOgTxWRbr3PjF+tmjJD1ObtSs8jFU0YrY+1b/yKJZE+iv
F2ulDbJ1obBKEwtD53a7Um3JWr7jSzBINV4/K/lafIwn2Ft7V3NpybfjMJSHwjk6SurZxrj2PpLq
v0PgNGyZXP1i/yTNL90Te/LNjYbsCdeauPr9K7+OBt5SoAoFOiCYNvAPZHBwFcGVarWfki2vD9Mv
SJOJh4VuRgjLrPP9RXxxqZfeEEkpiyVH/5iFI0MaPAvNlU8ay/RSI0IqT5oQjqBtxxu6DAXfpNZt
UCdOfM4XvUsS6iWJWEPG/8FRjdBvcbRMe7g+6i0Ono+D0m12EFmifgOFK44Bq+e6CXzJHwLW+EoO
cfptNNEScGjMOcE4jv0fCRr4r491DrJnQ5DgaIo1EafrGZrm4yaG6iSGTUpGRj/C7DJhNzmj4E3d
yx5iZ17F1ADtuYqVDibxycU6QrG5f1sP+KgYnomPac2zY4/jt80QwbDV1kENpJoarp23IxugV3P0
CEqQwarFOmUr3XX3J79vk33XWE+4IxoBIyCPuhFTsjVnY29OhFqVc/lKRi4C68fcMlzCRTj7GRT/
dgAkg3WZRiXhHbylvD7Iz39fKsb7Y+TL68SE2Feml/DM6v0OEnONmeqxqy7F1Y5Nsi+wozGt/Aqn
tbsYLR1z/h3wVVC7P7s2Ds8+3T74oFZUzwIxEHKkJf6snL8T6emfuWhp/z92oSGLNnubgy2iFYQf
d49UiswoxlqfTS/Yn0ZZgBQge3mk2sAU/gEkFTOlXOcHRBHz1Xj9Z7Oz4ftMMllOHdz275SD1tcc
/aftWaxoWNRTduJ/7OPel21n65Tc7LIazNA1fSUtH34M+hCEg0uPM4lUQLvZsDU5hgFpchOs0VLX
O/cAOktaMe2hCFdNX9eJv9x6mRm7AHwRQ3VHJnLcZODuuhqnHCGpqm/n8a1FIpT21gIZmz+evkVM
nRK61C99ULXrJgnHow0gJC9iUVLHIg/T0ypt4gOEKv0Yud4avst03xzi2dvkBXZeRC4OjG+mPd+q
bk6KJC2nog2AynOAmWsdF3quI4WpoK8YVQbIy8lMVc9wD2/xzbLIY/p9ln3qf42dmg4XCKnzw6k8
t74FZZRTHEtL7NS1L8RlaIhUb5Ac5u/HpmtYAjXfNZBGoGSGzPOXggnwkJhKQO2JvI0hOwmvocvL
v2pZ08J4zEYbYJTDA9A68hMZWFVLQPDy+Ra/NIV3/aLN3GwEHXEpwDDsbpxQfoUTb//cVLbaHqRb
S1WXinx66OA/7fPgkCW9phD0lGKJ/b6KqRDuJc5Zor74ZozFE/r63RyehhCxs9Va+kP+fdi/3b/Y
j7790uNC50qrxn7Z4c2PjlflXKy8c9m6XsewuTVj+SuqX/kxLFwDZOdWExkgG4QDTSNknFXoePpc
K4RNtwFQHqAC0G4VFOUcacBxrYE31jls6Hwyi9/zqnFv7QPtJfmhRJYJ17yRS9UqL84R9HkYH0vF
C2t5FfD86ViQznFSh+IucFkoCZvQQ2BTtntFNoftUHcasXTKUAHYrSFSDcxWC7Lc0wBwMSMwbZZ8
JbB8fiCT7+glhV/4c75rHuNfycU5CBzugD/PWKF2EAMo7lEq9cyPcgLWLXuWxYKsabHwJqfwJ0o8
PIslAvtxfUuTScHA2d1MsTcLl1zzKepQqVIJmpnEC3/sg3b9QdrFFn5JFrHV5owKWhMF2/NgCcjS
eg5Pus8HeRPAe0CGNIFDOGtO4nUgBckliuheOcxWc/Tawt9dwdF8+/H2qwAlP689rypMlFuLjxxO
IHLDMnjs6k0drw3IEdnLgH1P7QU5naNRPa5uvA7EVNL18wd3QQuwO3I3iguHre91BU+ZZInDiZYi
ttgUB6iuD8H/cxXNk4ZU46VAP5It3uUCwMEgauxwiEcT/NnCvCWyOr1J4aMwYjQcnCWUBU7wEb35
RCM4ZEZqEgIlBMqyDEf4jOWYLVOXWdUbrQxE+VVYm1j3soKl06BBK/mbni6ex3Y9oMR/4f+oGgSK
rIl5g+GIABToYV79NFKxgq36Jy6TE4QEsaNvU280i4+FdhFafcykL3flGb4mX8MB1MPHKiqA+22m
HO0qD6INJg7R2Wxnz3CUr1gyTC6+rM8+5XlJoI3b0CH6nmW5xZOAJ8JCLHAkKQ5c1mJLmXbWp8DP
Mnf1+bXqGpxDiPiTn48FULe1rgf8eNGhYTH5KrENxO5Op7KKtc2lGSUtXmmm9Xe8gU83t2N59ZP4
i2pKyiGNyOg3MSXSTh8Pe9f97BI7NXnsIY4jK3st6ikFA15o9LMK+qiq3GYwk9TNzAdpV5U8ynSD
LzQHJVfR3q+rg0hyc0+P9QR2N+aBRsHgIX/6KblKI39E2uwK9X181nCe6jbpSax2lbN1jM0bQA9J
pVj82BZNj4G2LmZqYK98qAn8MrFFHi52ukO7ow/vlOs2U5CXv3zFY8eh5b/KctwODhKDLUZe644Z
+jRKjTWtvEHEgknX1Iw1RG670lMxQzAd641TZNv63FwF1nlUbq74yqJfCBP8Skn71Hmt/rF2dj2S
fRhTcyMbwZriwepsnjfl/FecfJZeO2H6C289mVcQE8q08rtoJoxIf25N6jEmzYdWsEtPStBB2fHY
NQ1Z9dtQD1PGZqnD2YwmqLxZ/cNyQXxho5Rqaw3obRoMO8pVN3bFi147gezhn68C7dheG58GE0CJ
ynsWeLB801TilZHssKAV08s9S257Ah+wR8+w2ZsTVMhBnq0qL4boRlt6P2gppMDzDbtxdGg/shke
NGMfn59gbOZ9pOTM3OWJ0M1LZUQ8ru+5hqIODyVx9mBEsXwmDp7SFfFlF2Nzc2+sDkEpQQzJ7NZx
jak/fVOZr9Nisf5lomKwVUk8llN/XE2BAbAQYNQqnr5FzJblnV+3a8LaBpOzHp7rpbF0yCivAbQ5
HkfjMOutBaOMQxGZfB5Ewq3sRUveOper5rSUI7ndq/t/l1rrJ8+yjnRQmxd+rvbBKYh1+N3Poinl
GiMEtaPMK4dV+47PtwWBn/1HmNmUxbWJRH3U3BQfPut4xITN0PsjOZeWmZSJKr46KkgsX8zhlbio
RBGafj11lhD4ScTYKMS+EVwMfSVDQFsKPbjEG1TlKXtzJuYPADW/NfNy3vrK8mxd2ZfaslDpan6l
T0DGv7HjrwPC8UOirR/QoxuPWmz4eGIPStB9/U+iisfUkEWtvA1Cwzb3MZC27xIADtl/2BtE0gQA
D/8y9VNcYIXtUcbqLTftD9uZMUIko+4G0lt8AVUUzIy7SCntLIJmZOX2nuAHTHyNoE/mHqJ2EviC
ktuXlg6hXFqBT7S/dM3WuCeuKFbG5EJ9ZMKjIcEVYBaPrBsap35E0UBhqKeF54UBk2+SHHsA1Ar8
sU8LbJio2euKhw6tDDkYUC538x71qbPODZmZGZt6GgE3vaaxmXMqILmGOifKDdD0mQdimtfunlJZ
OnYQzu8f+zOnD+v7RwN1gXHv3AmS30tU1T3HsLJnsfKsgmZHY26UxujH5+d+nO81NsMJRxRYnPqk
cqr8UVfz/bmf8LjCc+RH/OwofTsxDYfOcHuNzLblk68+c2xR0/HvYjtGfUxC5q+hOFRhhTzFRt1+
q4Or1VA+UqBrdp/dXtaotj84He6bVWYIudH72ItSnl0dsnRLKqhobm7tYeU0XCQDCIN2qLfHB0xy
CIprsAqNUg2cd2mUTWcKsrwGfbWw69lgfgNg5urJ/YMKgyxIq21qUddpaQxFd4cQ0qAa3Idfc0YO
YQRtFMyllw/sBxWnqD16vAFDbPB4q9im53Ljui2q/syay1PMgPEtwOL1vnAnd8HA01JSK+uOh2hU
iknpHALeyOIoEUzwx933IzE3BI/O0uTK/nFA1LjcZ+6UwFmWz7gCjoV7JKDKhL41i/YQnPJz4z6E
FlZWJxFyZ5UxtODScqAvJdC1g414ChBRY4o9M6nPWRzFFzLjSajYkHIwLank6eACGpIqWoErKmT2
Sk1xMW40AxizfD96JDeqEdOd8u4VtUqgmdUu8gfcs+1QHoNxu1T5CVjSMZL1RCGmaPgbluoir16n
G9m+GP+LZKtpl03SpGVx5zfDcjZeL4TtfUVXfIwlETAmX+hznkm3ygcmiMXB0XF/m/GGtX3hbPnC
SvwCWOsb4mHP+BPbslMrbpUKHsgZfiFhwlcZA/byrHvjTs2j0XvJIDFnEu9vXlgxkY4JO62XdIeR
RYYC0DfgpfG76bweQgxVnlNZgNskLAn8iIamBpJ+pMUxJiPVCiEobi1sG2kdwYYY/9tivNOE5kpc
+sJVJENv0VurWd3mHHzzLSxS4MMGjA8esmqedJ1FkxB9YG5296AGYFD5OokrCR8pHE384eVJale+
U91JRuUPJEOx1W1AOQZTDl+oITojf8ZjsCwzI9x6vCVHxz+otDtscAZDGxIkqT0EKfeLsLO5Pwsc
/PX0jF86Vi4n0raM30KHX7rbas8gCrqiCBumDaz/p21YGhzj+XjjAc7CcMm21oUPveOzabVA0rkx
iW54rjGxqMyZWoSdLwy6k2n1HQzpTtTxmohKFz9YhiQn2BPyB9/7KvcRG4SoD7zHj/xTUF1brHg2
R7ImqqrSvvfGAFwPtN7cnVf+Iiz3cNtcMMGpnk3sQP28zI+wxQWUR4OPweQwngPYZR7pLcNolEPN
9BuQdlsKwOziULMPq8Kw6NRKnERzkHMSEiF+Khh60vnTME1/nkp2l5yyNtSLzpmcVLSV3CbqMoDA
IO3xw00HE2nEU6TeMonDrWwKoV6Mc6BiqwE5BXhKCUkmqbXgfcV/Nk7Uf846a4pVMnhuMqvQG4t4
awr6XaUNYGXrRa1M94whB3pR6hA0sTGBVfFBpQWliajw3osTsLTYRA5dVSNiscYPR/VSxV4kORq4
iw4xocoAqR2ifipAp0OBgli2ke/xELzFGdhsHTGPNW6X03uIkKpj82rEKDEM1+Zv3m57CF699yC5
3Aank122vcsZdGOw/VOcIztYjhZn3aGTLtoRMVgMGEgTGG0FFCsBBCNza6w7Tcy1FFBPVahr4I+2
xH2Pam8M7hN28AyFcTnnJMrwMkN7HycAZnPJntxBxSa+M3jfNJEkO3+E/qK2wb58u77lvIgPmgmt
dv2kNpZnmIyS0R65du4/Ro8YVCM/Tg0VhavpdjZOGPwP/VqTLWQtX069f0dtG+7uwTtVsb9/nGcF
Kzdcwcq0c5nwYDRyR0Lf+pkAfVE6hsqKOUf4OzcZYFaUFve7mdWe0ZIY50TT7/sSOtgP5POjsR2t
o9PJBbUXNg84F+Ut7HyYqhdbllFJBvTdTb+1v6eTWn+1GqRDY4FqwGLTAA/WFzRmwgvlpKbfeU8f
D9XNIf+anyQlSEgKo/euhBJgRgaBFJXJWOnBrLXMAtiF/vZtKCqhdGhKK6XuzdJnusruVQkM4Rwm
CTdMGlaToFO/vLx+AYbbaxT4jbwglkXGzN8emuAGy0tRMqyJ76ZOpUzKMrRCSFD+M1OzLtecsjpv
dqtrvzavuaHeqdpXf5C4ZdXAWLzNGTLstbPG++P/bPXSBrKCxMYYr6rCQd2V3dAn35o/2DbTnqPc
WfjA4uPF45tS+k2a3tgIm+JUJFyCV8WiHqyCidYWY8EKlFQTG9UuvvPnN0jiM0p6lYpRPJcX9q+D
+6zvg0/jZbIHatHlIUTppzBdU/30/mdyMiJoFy1V8T6JrrtOlD6UkdWrd9Lb8j8ctPmNnf8iaOyI
9qWCq47OAR0oNyZWftSJm5Vrle+NruQLTMahyJQsF117psGN9Z/r0dmhdmgt9xPC1dyJgTJOOwde
RoUvKkAOO3K4PHGpep/+RMVlvI8oXf4mnzlE+v71WDlG2mCDMR+xhYCEZ+J28nfYVT1cMkEaAirE
QQ7qx1M3PygMDuM9x5Xe/0yX9hPf8LQQpTdeiFVn9hRnP/eBJkL7/9RqpCxUfK0Chqp7ll+yZcrs
Sj98KhFmzEUN4y3CQEdT0g/LdIR6UbSuX8NdfhdU7Qx0mpXMwQ8l7XNNB3U9UgAS/+rDEbNEJGDp
fEdvWPSXzHs+h50X8q7TYtGk4YCyvHS7/sTU/12avG8AgcA2cIjDtb9OxcwLk0cszeWkNtYwEBsT
lmr9CdKDuCJNluM2lxssruTI2wly3oxMFiMG6qabSn99hnCjs8y7BkY/AtuHLR958RAn2c8iI9fM
vfu1gVFa9rYWsTFMg8r9hR2Rzs/xWBpGvdce5g/xxI/A/mrDLEyaJwKNXd1zB8mmBPBhBgriwy3X
GdsJXSwTBxoTJUFj4uADiM8U4zcknoQ7VKYkIgyXFsTeUVLnbisEtffyImod8tPUGcq2idTj4rY7
6KCggcXN26swCSs63AGSYWu+f+6K98BhkksOGKmiuoySvxHsk7XLjNOuUYXcxeESyKgqbmEEYalW
dIkWZN924wDe+/u40NGX7mfizNtwvn+jlA/I6nfwCze+McWwPcNNdYl7zDb9/x25edhcULV0MgPA
SnAG7Xgk6L4S5Yh/5u0y688j2X4qZVwNKz+iruQBPopKLMgh8MbEJifjhl8pnVg7scqDNp/VGfpA
YypqFcBcVh8uGbR+nfw1Y4QzZHEWtNJF+NGQwdxAhxSqFIKWERn4Rlo8bS5k9vbdXoLgFWJsIvmu
plqBARKF4edf/F/ENg6wlhcRa22puzgzmTfV/vtaBVr5Zcl28/rFLhfRosm749J68jciHY42JzIr
2xNXBFDF5IQDvzM/CYnt1lKeN5fIJl5t7Ds1hMTq5lpEn+jy7QNpuJMwSBqhkeR4HUIXFr73LH4q
wTFkg5958q6gfVYFJ5v3EUdzzinvOMrEWbyhSDb2APkcm3pp0R6Iol3HYJWmMjsKCEoi/6wbGfNB
XifUnBWWuVsaWjdEswLxGc+FhtWiCZmzlSjIro+/DODhQx1xkErqD1/ZroY5kDbayn4blK7iMW0c
ghYu1kDIO17FeQa6pgbDDhkT2+dJIV8eQ4VJWbMN/AfWnPNivBOsZ5lesB5FPcSATkkGMn69kbM/
0dMjYmxdomnrA3zIyXXKrw08TdNkH87GGvc4/CRVDCEp7EhHLXIMW08TH0LJyspkjHYpAcFaAxlb
CcxYtMljR3nSwJamy6SBFzdXwekxVA2eb3jR+ciekvQsUC9ug1Xt7VPLRYI1GfKC0KzHpHUK0ZMF
qZEnZyZEXvyR+m1qce+Eupd+95HWKAFr2smEbocBdgA055QhR1LPaKMr9X1mUH+9uXhzJ7atWSc3
5csq8/JtoeoDc4ub8BUw8xVjoV6y5UbndUThrGsP9inE0Qb4B6oYa03Ku64rPUbKMJ+Xx50uC1Kj
m2eZth7n9EwXjCtNFmtZieX/IrmV2v4tY60o12EMobaf+IeqahybTOa6ZQFWqn6RCJ7v+PyN9DNB
CZGZtaRymq5ipQyembmo1vpAcJrgVOxdGFzMFMDNLPICPuDgr4hvJsV6HlMXt6d5VR697zawWAjB
BmpmAgXGTExOZqoZYza6MEu1poJNB0eSM9qN6kQaLqEHqRpPJEtnx2byQztIA1sabJWvSJtw1lD/
x9aGyVDT7lWLL4h50qKvktodukAkVuggwID3zC40YQ/BXnqK5o/JZNkkNOYBI2h3E1L7Qip09sJn
ZnFbie56CxY0Dyb0Gib5hoaWGMcdjhF2Wgzt+4WghvGDcOaNMT0OQWF3XxcHm040RxEgLFO/++t7
i6Za0ZRs69OCJ4hqcLdb5x/SsNDwYRWG+NzKYT8NwMHECHPCGPhko3R/0gOCUXV984zU7lpFAtkU
bYVFBwgNR4HTJzOY8CQoMsNEsmhCAwh8UFYWbZfzKczTGCuaGqrjNJMk7sHfZW5rWP/sYXCwTXBu
bFXRyu0XKnp9XEf0gASY/LKevydaqQ73p/llVK2hB1Q5DSPnLn3um2HHomuoN0Ys46hkH65zNaYA
2N64frChkWievmi302f3Nl+PGFoGMQYVavtsxrsHRfHs5rPV2ErpfxZQN/ZJvNFGmOeO5HNe32BZ
z8u+0LSckUcxm6oxiCoOV9lk2UyIH+7rtV5Ng9aaeobJd13Xsp6m5FLfGl0pW8P6PITg8nWK76Pc
Pf7XzV3CObREj+OCDylMmmGfBrXdo3Pd9gVNTNXHQ3kyufXHgBPb6NYttu0pEboHlqRxcfABRQz0
2SOPqLg+kBbbq41N3lEZPvfdCvupjSd7/rHZewMwHhenrpt+BJEFifwRussTazlBtsTyv1nYvfvS
ib2mFCpimz2FfrMuqhqlRE9g9FD1tnwqeNAFCTipNhq9oWayr575yD4cPFvB5oGp/oHkxapM9/2f
C+hiSwzskOjr92nvVKeC+iDftyiK0s4WYNC1B94o+90qluitlUdhV1Zrg8B283Sy/zY/GXZGGVrr
STlS82/tsxQux9yZPfd3TnctWsDg3rTiDLZcdmxBG6IiXJ9OA33WDTx11GngvfQBmlXYEJXEfNjC
LqZdGRHu8uvEhSzwZpCTkOOQIMRg00+dA8oz633YgKjWkmWAEv+SoHeRphZfvMHBaSZMGooh1Um0
YeJKrBo3oPmCXU/GVVVzmGdT1SHgZjOYpkyHKdcAT7cms7BNilOSBo3Uu1bQLGYp/j7ofzKDxNdv
oCh6q5YoFPaTBuFK/730CpJeuYuMPqoW/t7LevBFqOI4mMlFqw7wAnqMzLG0oG22bQPWLLVluaaB
gkPHnHCmIrx+8Qif5X9045sqxiofgUuGUi6GPSwTJyet92CmCjKbiXM3ofAQzt9tuzQW2foNhBSs
ctAEmzcWTjwxbZW+FdXL0F4yrMEmeimljZw0qsHgeu6p/q94c3S57p37C3vqHG1h4j5ABuONF0nJ
fLL1BrNiiPAhEdC93Y+BRtWHpjI098tGdsZwdctbQViYPTkDB18nHAQHPT0h+EU4y3f8pqPWGRZk
RACv9Mo5T/yJ8FiWTwhPswPbXaxGf+bWJFO8L5lCJqwCl4eHiLP+t0xlAv9HGxIL7mLWC9ukJqb9
WClnu63FzFWRslr7ouJWK+Ubuy57mW/1tv6CkJJoHYybibixWtO3HGHC19SNi1VVO5/aa798LrZ9
MZ7tXYAwj11bCnR30zGmU1VZBR1IPR1sLt/qki/Neu73vVd9j6WviFoJxLTl0nKZokKCYF8t5wZv
510KMrf8UKNygyiIooXv0pQDOsGrO2yI/tMhtr4rP4tqOR3dPBUEchXjTYIMikI8Dni+avk/Me2z
6PwxXCR/wYbQiVIMNXfDbj6MrxvtBZHlKfsFzx75aLQ/1wpdzZ3In3juFO1fU5vUtqQl+y1NZ4jr
VEQBVnV2NRZKw31f9pim2gHFDGecWE1lbqy9DxMjML5pqU0fHK3YaKnhVtNnE5FbpZpcLYAP5Rpx
n6BIH73j9w5+qQGfB5+nRWKdF4/yf8srtarphIe99g5c5hvLLPoJMEZA/onrAN2kQ+A8l6c71o6n
HoA4Zzji7AgN036KhnF3XA90186s5oDGoTuG2e9d5gvU8N9v8ioTtx+UsuzzgGqpoHqpek6Hx6xh
im/83n3NlxUcG21iM9Yp7XeIcp0uLbMLzS6TM/2tJuv4XFfUQp1LK3qpUi1A8hXaklyzj8ix2JOZ
En6RFsWs35qKaA9XwFxbql2v7kF4ZytU4ROXYLiB4nDeIDfOXPAQ+u//J9eg21ZYlnW3YMfBQgol
BOBem9E+Tjq0HQSgy/NCwhIfpRn6yv7wkwRQukFVe0pkuvtT5sIQt+875rwh2aVVp51DpZXWX6f2
TKInQYcEcaFOZaPtZVvYrJsl1rS5RsvajPM/1JPVyXG/RR9ZpP1IXFpwccDpjEq+w1aElrAwaM3S
b5bX4x4+4OvKHhN3ktIrOMyqBrPb2cVUUym73O9Ey+Rk2zMH3YqBN+wXvdAe/j5YPx4aoPan196k
ozvgLGKLVtJQwYYTEi5wI5Ru0agks9H4eUcH9XZ+0yl6VcbMgYdIUAtrhXMDeUER/OBWARi20dvW
0D5TXAwt4NK05D9r935UtHoRVSXmgtC3guBc3qz0HZEgfMaIb7nMv9Zbh8lRHL3OXqFzMCIKNJdY
5m/Y2s7CaH8UzU966C3s6YlO9PliUcMdPVJJAn08fojYfWICqoQkB+WRBAL1q/vJrFLC9j4MVOhA
W6WihpoFqHuo5AE/WV1S2/kmRugEq9ibwy+/c5e1qF2dlhX7Gfk+3iw+I8OsCUL/urD4mwKpMASO
mhUmOSH6bJVTyCOhdxd00z2Dn5B63SmfMM0CgY8yNcL2BaUU1ay0O4+sFVEDDDD10nEm6leggpXO
Kez2r0J1OILPEfDyGvwEsufiILW+PV17LDkx+ADTyoiu0vBfn6HbzCeKAT6pKmNCHX3ARJjM7b1s
QXJhDEWbfI/dnGqLK+xJt8SwVbj3Tb2/Ka2epj37nb43E/ITxEYonSqTQbEKrQYK9gU0ssrLvCNb
DmD+i3cCuI1wiDK9y2uM3HtxcNnjMmWuNo46CX2bm31j7ARdotTf2f0WIQljP2Z1fcO2KsNqee17
WxJP2r/vYS9Fxo2rPCf5ro4o5D6wi7mC0uPSwBK0xdsQPFM3xYJ7M9fZGffF6GuOFzTn7n482ztL
9FJlZrwu/9nl/xLa79LugXHyTsspc5z73sakPS5noFDE5IgCqA5dDIO36nceXqWh0AcuoNj5CBHg
JhzjHdLK0OW1sAjw71JmAMTq/KF/kwARRM92rpDnoabKRrq3VP0iyX5WmwlspI8b8i0W53dC3dHP
BiB+RHNQJeCuYK+EsvSbypUYg11mAqLnq81N5du+EU24UJQxXfikTa+UhiiUnBTGO92l8PduMVuP
WwAeEnolrqJe11BFYhYegTJyAg5/SCQa+9ApA1IHmZVgXArpWVdN4zAr1ciDJ2iYxGKFGcPW32N2
XwvQU54xgfVj+sbUzyxor1ZcPvt7MhO5rcY4z1sr5qsAg4rdlkkdxmhZGHvQ0V8pLsoP8fQLnUYj
gfLqIcGWNdZAvVcaZsfE1Cb3ejQsNk4wTgRjUREcOFMV/urdjmE5yPGaFfm4ubpMtBsNeSIl8FCO
7acBJGDXwgdbSyHyjbH2BL40HdpFJG1kh0RwAdWE66wQMuqa8+9jTOIqyJgmwnywpaQppZZI5Tpy
N9U0wA7dsP5w+XJPa9lWW11betjuPVIy2RxuF6oP78XWSOdfmT042VU8ggOL5aF/ETjdR2akocLr
ib5UCSOE6IqG48rpeRIQw43baGKgKPIael5n92/TB0sDsIH22534C+nKB8eBJdDql4jTootfsT1G
zqafYkR0RrppCKFdiGC15OUFNb0mCMjifFV368Yxp1wgt0Iq2ID7ZP4GylYBUZCoy3W7aNHWzD63
0NxDbCvNepIcszxO4zEyv/AF+uhoQGMdVerh4LbcjD6nEd4+ucn2uZC0UOVqyUKya8qXX9NR216i
3xI2MnbR88NdrGjTkav8EGwFpxV+RftcfQZIr2Vp6N4UvsfL80pM/YNLhUSwAdW7D5eueqifK9b0
QfnwDq+jRxbnc3f+YHKqWLkM4btlVG+qzj51S0IAApOzub7N1RKUHsqnQA5mi2mZdk2w6pGYTIBS
jkdX8ktwDnb36aUpCVZoGLV18aFAOfOBN37VALQ/XtPRDA8HgPTPdgE47tCgT0rK6GPhdjXc+g0E
QCd7pQWh5345RTFOTU5CSWcWdMEUF4cOPx1QMsA6j53h08zlL+0EOIJ2DC5qgBPnZoayMQVuFSu8
qTT6BY7ffod6SMZotL7Ac2IkHIlqyXZCdmQ3o0y9uFS6FvNdusCUdILj8tecHfkk/UNPJv1x41SB
pBihzCzH3SkI6bL9ur/haghkH3d9IF2kCWcqb8XF/VdKQnD4ecDSGXFEXbOcH19rqg5O5Y/GZ4nS
i8le8MsZ5pm4ZJeh7eNI/yt90bcFP1vsesYMfSaVzpsuHTfXH4664rMNgM4GG9rn7PrAxd+F/9MA
Y2VO1fu/aDMcqe5w3kTg3D9l0XXTMk/IO89AxXPvyPGlJ0mwRapu1ItQWkfo+sKyzGdr1050fQiB
QSw1wurna6PwgPSlC4bhSx/1qzknK8KcNz8iMxQ8dRnovXzZczezAOA3qBfJdsbnMf0U4xFXHdmS
9wxSS3LYNBKGLEGxPVRBj2+pf8T66gTIzAUWojNEPkWogdrN71HHcwztHd9s1DYxSfn7ij21jgOj
ynuiHv6PIbM2Lj5u1bWRF7nREUfc2SxzLKaMZ/IHrci2DszXmjfESjJYmLXbD/udoMhvsdg31ABh
t/QIWIdXGLNlMONeo9OQcqjhl+tGHGfJAUCqajoPHzI6k7UgWIWrDDSNqKKupPIvnyhMeWQsL0q2
cpLUAlKm/TmZnqTIyKQnq0jx3EKoT6cXrH/7b3NmiGGVnYjRjrHgTSbKaSReysG/uAXbgKfZFXZE
5aykcd52LInRW0/lOXEfkjS+eHqVOxrl8SVnH2SEyNK4ljv7Txr4ZV9vgsTbOoN0t5szQvKTjm6A
LLww+9aiUdzSLs3JlCgHFQYuitzAjRLqvtDX3mBu87ACmbOkaOy6oWPNMBHVIwcAaLlQu3AvhFDz
oc02z5ntpIzVNuoOA9+qXNZZJsdZninTHU8shK1sPutzT5zRE/an8z+6WdsyALM7dWCQqE4vUpkH
wZ4dyDpRdIkA3i8tdNdS0SlEj3N3hz7dfhFjFfjGJq/6tnx+f6f3jNaOKm947Y8euKPyxyquCKsL
9bFsW33nIL8aoIfajw2v67OOPy6hz7T4YsW/7Jw0fsgXI++wkNuChtaoVneIhv3ESg5c6zI2k9B4
MsemfuDsEmaU/LUQFXAbG4xG3WmJuwg8xIufWTjXnTgxApdcQxYr7d9zf2Ry6eanmNRsQhANtKV8
5VJaNsELjMgSO3KFTi2qB44bdYEVkbWrrZ+nlcMsW+ElEoMKoHfolE6WmjoVZpAQwfLIUbhqx4NR
+JwDLTnXSXaTKQfAf5+UIS7IkxrHUEQWyWEqp3b1Q9nXYhupOh+BKBG8eRZwok4KqMcFakYIiqSW
DKfowrc2HkVMZxhHeq1jZUNcOXGd15uxong20/NGnca12+Qf24Wav2dpPcrWyaVgyG9CwCAc4bdU
gcGESbgijM1y8vT0BWpynFF7lQe0bwPQjGN6u/TXYD+1bko9cRRZdW0za7DPeWlktMBbV7PWCcic
plMM/SnRBIXJHA3JcxpFlt9oPxiTIax6hZ+NrXXM8SMUf02M3cPos+a4+0GH8S7CecrMxrYuwfba
PW9hX/Y3KD/L+IGR4w/MIS0C0ZU1Qh29ifw195FKOLwgza4frgmKtjmDiIOyXkjfPwL+f+7lf2Yv
IW1EoMwSetLUab8LXz8r1hjxj/iO42Yyff0lrtQL2+gdnWxwH8zp9fpdQ9MsGyC5y2+tBOxTERMw
RWnP1w0kTzeT593VE4yTeRPaFZRnc+5ziBwBtK5rzamvPysBgDIGQmIRbob8nTlbZDZogqUJSP/W
z5iVlwPGIr1tGePu5vfIC6XATcjO7S/rvrauCXk6LylMvD7z2QVBHwrrkeAkrS7PL4CuvoFMaAij
dWM2Hh8dc77WR35HUp0pXW7wn657baB6FN9jlTyt5ozaC3JmkVdcdixW06j3Be0Pf66lzBtJynuW
mXsoM3JMfMmS3HIPofyXF7hlU7xoBhhId6QkFw2+KLG57/4n9WbdZ0LDXu9mlRhTrs4tKi7U4zQO
8nQyPT7PkJse9Qk4y7rq11xxcb23ZCqMue/fempVIkex/LTOLRXk2mcpnq0dj2azLL9g1HgcE8rJ
Ne1eZOPvB8RBbTbLUYfy4oPEAc84Qyvgt5UazjYS+i4GSkAmOL/rG84RJuEIBShkRQy4Ui6gjIQZ
tNNV47bpdPKvTK3FpxLwM1YwP+LpPui4Vpid8x3I+H7EmPiYT95w2QedcQePH4Ieoc2PrbiFNCyw
PtDNFQx2K6l9krImPcGJ2ZY32EuB+O+PSi8Dw2LmMeN6L+Wwj3yL7mCWgqmlRx7ORttvxO6nsTcg
Nx82xwzmr12QKUHn9w74e5xg83P3Q+w8vgaAX5rHhF2UbLTEp2ADQonWTVnyCNRx+kt0hvg0qroT
rU43f1iynf4tYQ4FriBjXdSY3u369+9X1DAjjLTgAi/IxGkjLmHUWfT7MJh1PE6KxKzawY7kOmvL
nca7xiAFj3syUitK3zLHtThlCqAl2IBmat77bVP5I3lZMmliOMqHDsdPHpPXoKV+BIRdM2W4Eqrz
xiJgt2Corv7SWvWgL6i9Ccl0mYyW34uqr+QdnUphLpH1uaLBT8Hg2ezsYGoIl22UI8ScnB9gwcC/
yLumiipTybdiUlOwYuAGIeZQGO8UyxdjhWQxJChBfJsEEKnRYubJTCu/oyBXobzmrme9S0qs34uo
borwnwAHJWLda1Im5dpq/peWdg0/9II8iVB1GXaRTwqCpB0+XvGtXJPwHVtk2WRQrLZsIjUOC/h1
5mm5ahW/tQU6PTQamZEKPwz4peRP7SYiI2C5EAoiKnz+uN1to7KmZEK0hVB2ZnO/1/VUvFBlM8b8
pWSg7zddcDSkrwEqN0quqK8+N+YnN8Vdi45SQfDYXKzctUIk0xdk04Gy1RPdMtgV7mWD7gQ3Fxto
eh8nFyCy+IRcmw3t4jSaIuWnntM0dOJFHiwAJuQOgLx+B0iagIeyIyAqwwd42zsetoKTOXf+ouhb
uCch2bMC8uTzqPGj2Epuxu5uwbHfaX0SKr0KekyHf+IH8+YO6hg6h9yf5i9OIefyHArXidJwR4kY
lWl1t2b0wbe8DKPhHkp8qKiCpngNMciS/Mx5ze18QD/Gvs5NTp4b9jHx5u0liPTZaPdpv/OW7AKF
JOb2GjSHvNNU2pGM1Rq6IOqqGiAbPN6ZUr0E4WcAOm4gurnl2igYLumDtpwQxDTuoKCOtFH2+qA2
q8Fs7LzfT7W7MPem1ce3lsP6ZaYKaJ20a98YkPcOtZEhlfxgOAbwR9MgmcQOgwlO/8tY/AyEBxpn
fo6ANaaLqQV9vTQhFyNNNkUt+4iTvRmJStPXS3YRPRSDxxyWin3m9ZDd9p8H0nkJ5gNLD37fcKe5
NuuVg4dITY/ugkLzIQk88AhX+Yx0a+x3Ek5kNrqHrifqHj+lixWUyU+71n162fz3BNtjR8Sizi9y
VqRVVs1WoICv+sK5ooFudXZyzQVpaWbP2Wz3Jdak29jfJboHIXgp/IsmtmBnVEDvDDWabkMV3E96
6SwEEDAosiQbLiv1c77xfzqt7cs2CWA1bN+wkSGADogdjXq4p2dFYZ5irQw590qELcf90+MLDxb/
hwVaxgWTkLDm4Ex6gZ8qRSaS5WOsnocBPQu/xRxKL70wwztEJkf7oP+o4H+h1RrEU4wpNu5jwSpt
Kw7ZBl07fatCFr8Mw5Warmr4hiwEBG/IIlyqZAz9QGrsUGyxbp2vcnF4vdiVDTg6IYxqb5yJPsgg
5yrSSqAlyLUjXwWkLdAUw+9gBshcEq+ZZja2nYUnyBeAhoM8D/Ii82RPfOwBmVhRz/qfepujxpqF
FdXFfXjbdtN0UJsx5GlxHx9n0g07Etw74AjPqKTp2xyOTEsTFAFhGrO53qZwnbSHcWDXPCIJHt9S
FdqfD2ZxP2RbD7j1esEeBCHpCpHYlx/BvDnORqpCHr83CHPvvbuBQa9G66wRt9tMIKBGG9vmj/a6
+DHz/gi4sccNtPCItg7tGzYY6Hvlew58BGU8R+QoZF50Qa0N1MsbXBFGG8OyRrbX+mcWrXIGIwdo
WMbQvxAr7XFPMi1nfhrG8UgGax2gSYkq8oPj3dqQhZZcWlQMM15Zl9+Cl+qiPMyNwtq8MaOwMtVJ
daxSd03BEJsp8qgDhLr5gUQIVNciN3oKRwhvhtG3TXAxY5F1WflblaoOVY12p0sZvkOF7HPAES6c
ZM4UMLGuPN1MUb9ObLT31dq8GBYttTPoGwmzVr86fXhMtZtzLtvP4RAI2m0iWvgBUTtJWvBM0T+W
KdGYhim83aLbANQTD/HyJ6BKns1GZDH5HWd5xQRxekyMLglcVUKNDxrDFlAYd03/Rteg7BnYrwkT
2ZsIvzAGzWmSKXf7xiIo96ulhKWceD3HO47DGDuszwmjKKB4cSEodEH+6S3q6Gst+3ThrAOv9R3O
DLEQe08OGdEvi31SbbRMzQDhiOkDWdUz0RV1UaLePPu0fopSYmJEmr+wcFmd6ZpXEtawT6hOSAx7
cs8pESJpZyhJGUvFdev6ZY1gBblw5ZuxM0XM2YvguBXboIqSuMsxoMxFbSOgQlvxvo0cemeP/eR+
UY09c508qacmmZ8w0Z4Ln7Dx18LTucaAi0EAZxcdW7tMM/3SK1HWOg88iiF7BPX21Eb6Btpvp2Jf
GKBMV3oTYZCabQwHjD0C1nNTF6aYBSaeSC/f90Cwq3g0CkI6oQ6pkHpWkhTexI2G0BzK8s/CcDDp
cMeqpJzLyvyvsnt4rpSlZjN0Nfqoo7uRvAuKQpgQFI1WysHIyWDBodVGgQMSP2c0lSgFmhGU0dAd
8lJPutpKFb1IPSVXNzn7IG1RgWK9kgVUnlCDVZi4d3jzEJmmlfAtvlTv5L8+pvkAhJorunr5ge6J
PqXn1M0N22kIZgD99VShr5WOHj3FibotE4IjP7HOY6FhUCSnGWD9falKcQ8cGrGDYnVXlwvltKsR
UrnEUEJwX7znvp0nEkhlIbxa0o+rR7YlkwTbLyEV302uvCvMKBdAUiFrXsRRCzinPW/eN6HLpHWo
1c3+P8M+LqIIn7lNaWCuLqM1KwNC8Ev2v6yZ9xMjG2v5ee8+yGqW6GKB4MZUy4DnUWPk4JC2HNDp
S3A2uTXwyO8uNI9fndMTsSJOl2gTr65VW+nRkKhUSB+XOu9TqAIydC1eEiayREqn+9hmrf9QD7zX
T9me4YhsV2oEQrpMQ9T+LANT9YpA/lKSvImz+ChhwwkjZqIwNXuNP5C4EFtFctrVHkiR9JsmKvoD
/ZmJoNRhUXZ5LKk9YrIagI+4SNmr9WQx9DVLfScIt//JFO9BgVShiic3yOWfBL/S+tdHw5zlU5qn
PoMp5bQ6eXS5bDCN8mcpEaBEQaSi8Qvvl2l7OSsV7CFmvLkKhCZEPlT3Bm6LchRoe+sJ4yOy8A9E
quUzwRBHIAFNqH3UDi45l0g1v2DPRjydj88zC864sPOSHcqOtIWBlfbUw7geSO9WzeBeXK95BRiH
3ZWcSkOzftVbwro/dGF6pB1+9btje1i9rnbtqi5pCSXJsSX5tAmYPn/9BYIWXAwaPWNlPczLwDg3
egpSD/3G23wTwT9jJIwCTRgcxtFW6BoK0QJxJodjQk2W0Fnu+7DCEH2OlPkcvFrgJuiwtPXezpWe
XP7Vn8PnY3GhcQORwomiaZNZ6GyN148nqqk2iVKOIBcVzx3dlnrivDI5bOR2cExZxhihQecofJX8
UTYfKdrWdz27Uzy/AkcfM4/KI7I4RAmCiz5IGLYwduMuDg+6gPJ+Dtik4+guxijiJUOjKGNg05SX
UrI0fjiFZTFdT164YQe/f+rCef5X2ZDPricC7guq1QuUZ7kANeVw/LJ0YxFfWx55CjsHKpr4JtxX
cHihXUBCnT4M9m5xCrinGPayokoXoZtrsXOZ5xnNvimK9bCxmaaBa7o63XaQsiHYGDobrIdCiqRS
CAiIludflnr1dJfUitjGlajCTGM4b48pABJ5cU9ZK1UMExyQZkCVzmN/WdwmSL2dI0U19LSwicJJ
lBffy+37GEgVgiSpfmCXK38XVDnuMK5TBLAsKJ9Q+Z97rudEE2WUqKqB4ngioJXKDwBia81aXaai
VLEoto3wQ4QRea68RSq/fPi2SSWqwEbz0ygLXHsVvWwvbuYOtPhG9R682Rz+opDrwNlTJH2NsJ8y
XTpJx0v+eIUqSnHwPaW+6oNZNDYYzFjYb/cVEGOKDX/SgvA3IulbPrDW+u6XQwh6mxR8DXokk3M5
MJiaBtalwcZVy7tD44gvOOlcY79WcxgPxWC3w2ZnLSW87v/HWBX29xgj3beBdYjwm1YX/Sib07DB
VFMS+w4clENAB8y7eIzINp6+LfxqhLsZ4vB2wThl0k6va5wN3dib9VRjDvegrr1rovxCmusLOoDc
uYDVs9HfjfC3EuZ0lZZxfw4ISoLXXrOnhuhBTqYVDCM1BtUBeDmgXQcvX/euD7ByQ1t1gHv5WnQr
/CCxSwhLqgxaaYXECCA3rA/CA+rNi/Q3Uot7zgK+xJFREn2HnFAnkjrQzDN669AO8z4eBrepuEBJ
mxZzdWTKFJX78s9XAGzqmQstB/mUFyWP/kZ9et7gUBGC/DTfiKXL7QLSdTLaZ3elAHtdyVeH+1tW
X2O62Q6/eoOKwcqKyrtYUVHNKJbdONQPvUNqXrbyWHPpQOoSPBL7I+TRCAmgnb3nBwz15f9sByiR
sJTG5Gos1pVfUuG9r/wjs6NctJ6Dsl38g3xXFutAgGNhFZNWTDRsGXZG1F5qR2xeXqJ6fJlPS3Ii
2l7nalcDUTLaou/5ft7EAF4fA7IYMEknWSOfIzVzhn2IE/nrfWUrGq3OHDnajl0hTDQdb/rWDZ4m
eJ33XPVlRCYIJmAYRttCBgD4k5w9afQeiSULTjGtHB5gKIktXuroxHyPIgYLHu3O4X3mJWHi3LO7
OcGg3I6WcX1YYZs25Yjui38nFIxDkvbbWNZhgLelmPEwnqWsWaQWgeiUNKmhdNQ90D70HSUVqEfe
gORSi5wlWF5uf5FwH8Kec1YE/K6/rJWzryiukqVPZ0G+dmESkXRB7wAxEqHD7m37EOMVh1IVxPh2
cbnSzOMpXjeD4uMQpnuXuQS5CtvZMGACrUUU4z84SLV/h/ncrtSDC4Jneynf9+2/XuS/pXcDle8U
mXL/S5QKM0qK5rExJ2SViL696HLhai+YXI/cFAbIemFIKQ9zlDZAbrMbWhvNK4vFd1gWZxasne/6
wSs2pIxLlBl/ZxOipx4cF4rgocMEj7/AQ69EUGeEf0tQ1ZAGfKT1sXH8jXXNx8s3C4nzsE4NcL+n
0Vb5BKWU9x/F94V0UaGIUGtFr3BKkB3JVEPCTGzSRiO2a1PKoURhhQXDPxZkLZE65x2LgLHEc1UN
GT9eCclOCXB66RpxTJAA/xJhGD+j+vPQP1gkleaDGEF0/gKL76D/r4imqObuQgnGAQ1VzCJCgbrG
NdnYPOTd0Y+LDWTLOsuJwOPjO9+7D/JJfyw8mTC1oy77IDmbvxscI14VNm+lN9OLbZmZHjvstxGR
1Y7jFHBq6woRxgVF04dZRDsrLPRzgW3fW0/WEbihMnP4fg1wJ6/lR8Ssp5BsE+qkZ4nY6purozWH
NauQFdFUp6lqGt0Bf7V78s3XOmsjGQ9nTaONgtJIJP2dHnWxLSVqO++ZmTwZuTTJ3Qc4iBHF7PV6
h//h+oL2sq2NBv+xRA73g8lUlBqAr5rpQzG+gfcezX0IhDrbfxin48wkAwF71ecuxt7lqw1bCMfK
n4zpmkvdzsni0Af3KmIJotzEBCg5ct4olA/RA3GePNBvRE34K7FxurF3KryW4bR/aChFXTJjl486
SEZS/7EJSpFEkf6TuZFAcza5tfxJebNl8Ey4RozgXpISMowH/l4zxv0t+xaHTNqwo4RBqKMl1Eyo
MAzNvWQiGGu6vev8Dde35vgbJsOlHzCipceLlRQohGAfSFtNBmywI310Fu0g4Siximu0S1x5Jyxz
29zWwmYTw6ilSHSx769eTzehG7ndoFYgPvHmUXS+vYhSawNy+4kvSYoM+9zjGFlUnhnSWXYjoo0W
duwFwDlEBJfbwCRHq9vxEK2kxl4GX4ub+yYDJq2GDVkfbV2laZvcWk/XCKAw1BT2UA2SlcMWubjH
Y0X6cHF509emTj3cws4pct3KptrGkuFiufNItJQ4AbHjxpvIlEgGBI/ta3rIkBXJ5GzQEn/FHnsh
a9L5BQqd2/gqd9GSIKhGnUI1JIeaN8XAKgSzAjPI11KQBWM0aNTPGILafKMvUgC/sh3wsZDGSlok
ieGNPnLw3Wv7IkVFSW69urXsZznaRm+NdZpPshHPYGPTaLxhEn4dtFTeMYwtgPrG94/Dq2Iybx1n
DlExvnAFqR9ly/9j8x7yW5QBuBnR1cO90UpRokxVqsoATAZHlykGFWn/PG+st9HsmBRcu862Ew8I
4kzGyI9MxZCVqi8deXdvzUOComd8XPlE6gXAaASnLM0GXo3b8GrHSavO1/arzAKS3pXqNld6sPLP
Nu0b6yJDNgwKJzGShxThu/jKRtgpIf+ZyvjuPutldLjaVjJeEQ5aYeH0gHw1/XqfZnKiye9uxMwC
D0U5lpBtMgen77QvX1P4zsoHYej7cX5Aw1wHOmPBsTGBPppPR3IDU6SBDd/Rnyc93txaRmRXbdmW
opr6a++oJSH5ts1YVJQlCCHR0GYmCOeQrBcrgFwVnK7DXtEJZLmm4u/uo9MbakPzZmf4ajm/wnW6
NN57wJGMMsOO4cw8k+EHY3XXjPnYsc9Ij5DzbwIb6rqscMRnv9x5CKPiViJWrUn3G3nDMLfZI0pF
XGIi7GxW49nbaj4vUhn5ioK7nr2gfeLJ3JZ6N8bIWdz9ODVXbkKoTW3uCbu2zBEyZhK/XM/AYshA
QLfyuLS8vYeOsVeo85NwwdfdSa7PxPXbN+Z+Fr/iEFKoiRZgdfttLA9drYu4fY9p8RdjXSV18hs+
yxAr14TSuRTMkB+bEW7Gm/uxELg325PX6ClamzjaizkBIidc4i4Qj+gZye1fbynjw6mY+76JuFzr
wr8xqJeoVgoaTQgpJ+vWUZQfStYeavxsOcssiNYKv1s1qyIVZCWeQJCA1SehxrKPfEHaCY7cJOsK
54pJXm6J6f8iU1hQRQwNNAZVnkrRFkZ6FFF1MgqaCylPL9UAwDVXw9mDGx9moRfO/6lezPL1n3LG
BTCRUGFKjGs8VIq7G1+pZe/xoGRwl2Htvr6lhPVkM9/Uv4qSzRHY9gl+UuDFH6OTKtx36mZ3Rzya
t3mpMXytxV5/ycUeFPirubYCl21XdhiDGIyHg6LuUzpAdoHeuOl+N9rRP6ZdV/iLI/Xueu9/idDY
5DCRmb9nCVre2x3ifDVgXcVi6PDd9TgMLIQaZ51t3ZKHHcEhU9rtYTRH57bDokAVr3xjgqr782qs
smVlJsWYnt918vLQJFsHcpNRgwywydm9GK/Zdlm2ptbzeDJMpQyK/dWx/Tzn+E6lPlrqQYQLBh7z
0GATFIKtcoS8TZJwqeq+RXzHMgIFvy4/EVrJ0LbQSrWYQwzAnYYqRq5mZIQ7QfroGyAwDlI86BSj
AWeDNQ6XqEQ+K1PR1rpxxG0G6SdbQuToLVDIm8Mryzc71w7Gxm1MzDFM6Rw0MSHFN7z8IYaIpSZZ
cs0ocfjlhQ2FGVLTC9QGjwcxZS+0oO48e73slAxKQlw4l+UvBbqx4avQPVInLa+BQHTmIp1uGXi8
T+Sennuhh0eKWeCg2L9YFbwx9vQvsYpUmWP7otRmSfUP/dGDEvt86dgfD2gloSqPNEMO1MuPdtg4
EtVoE6Uy8VPApbnUFhDvaBMuHKpirT8TBlZts6XC5wojMg0KFzSWJjzIpJrUx48P3l09IojrSlnZ
3pxJ5QGwkwidQCfrciU/rvxHMyiizmHgXYtoNgvAHDnM0vXDsGNYYFUjeB9iTR941pTSW6F1uAmU
cl3iDZ7ToCw1aDECMHypOFjEn6t9cB50TVzYgQCrdHdhQlQaax2xWQ/rS3PUwoIO3O4F/H2n7AkT
ejYlVBzn80YCAkBHGKRFdqWE2/3NrGeUyzPSOOrbGYU7ZcSQiUG5BX8t1ZGEfhDQbuaV7xcMwlom
vz7K9cG+3e2Xug5xDJdkJ1Kd9exPNmUlurNyhHeb7/JOcKzL/+d67qeS3XycO2wdSCsgzuZnz5+H
uHgD8L2c59DPB3iJQILteXUFSEPq4fwZfNwlG1pT/g1yGu6wnm6x2J+clHupQHbOHzCIao0gKSJv
aoSk4H8P7fJIltBvfckIQXQgbGt0Hsgg26lfJegso/yd716G+6k9r+quGIZ9SC03EVP0pL4qYoB6
Esu32BNSILGtmTHzvlWXGWxpDm/I3QBMYW86IoZgGgiPTPNZLWJlA8L1B9ujHyekkE1VIJRl9RHc
jvVxfjznTun919lOK7YCBgVwPrnOVqmzaIdbKUwwHW/KhZT1Y9Wd+niasFPtNR6BMa4Sf+ztAyVU
h+PlvYJoSkmHwb5sK4ImzdqlpFKW7IRCJ20JNjPtJY1+/sBJ6zMfWDl6rzXI1M1AQLKo9lewl+83
Y7BTKqL+IRnXo9dfImXflRq286+b+yQOdNzTKJUq25EPjtXUdr7IQHQ08Rfe6/sBi8YB4D4o2viu
nDBl8d5bJAEKal3VmZaAsV8yaI1RsrcpaciGMdwy1oy5b9xr9In+N+stbfrUY36Gct/AKqS3V7iA
MRHrq87mTyyA/ieXHmkxgUR18MODPE5U+flRzoKbS+I37637NrA8Y8oxbDSNlb/7sRDYxIwkKk0A
Rt283m2TY62dy82vlH28vMpRGMZc8KaDDC7fn1+QOHC6UKre6Bo7ms/P5NKqMRTCfHeCAsdrK484
ZnoKP5kW55N0cyH5e7MjXFvY7yBZ4+f6a4ackREhJnNpsKt96Mjps+PfK/1tf6zVf0uq+w9w7gUL
nr7tCh2AKG90pYnxOCLhANN/zdeTUGRxAR9jdElZMNAP+CprvyW8ZDsdF2lap0DJqbXpUn7gY7CZ
SLeKlrvKio9+EewhBQXtxTvVJMgfuATEsqn9ScvC4BO5yAnHL1wTNYJKBtobRd+Pk3fwUtJNHdLC
kG4vjSnhKvVInFdi6iZbMW6LiD+qr64CaN/iqYLbpLYxFVbLeFZt3d2N5IeVtxRu6sGUkMcj/spe
RdOOa2tFJK4LLTo7G4kJZDsOlQnxIHunFT2rMbmulpF/sQbQIXDoijjex1XrO05jkHzSnsSAmBrr
xv9ifySuiO58sqkgM2CysDFeZfOw7QmwROojZa80rkJ0EgF4liJlaoOW5qLHsLcIKmeKiOwTjoln
WPEQ1eIvL+hrzqOqJDth2R64jmIRABNn6ndZTxErDmupufMKZX7stMPY4VndVvUgFhCDFXqaBtZS
Jc1rR9UcatHoBB5g7BwDTjFqEQAcxrvOVQla+mUdYjaKHyticVVSXx5fBwcQtDQ0FAYl7+7Joy8F
SmnnMPg5/6pDfk8/q6MUxykXrjHM15Ch/UVu5+x0NuiltjarW6iHBqjLoldyMhgy+1XwAg2Xabyf
4Cp8T2A16FSeL+0g4574ZyF5htYurR+svPWHQoN3TeqpW0X6NtvwwqS/hjgQTW7ShAw57O2Kld94
z9DXzFDBxyVdnQE3X5dLajczXU4ssp+zQsAqTw4WEGMmRqCgbUwfZ2N4VE39f+tVzZcf/sY4LYJE
qsdwPoYpglkkneYjtWML/nuEGAW5EYK2zoKkq4KDXEdoRTI6eRhkMbOjvoCGCM8D7DT40YMcBZlx
f/48i1pt8AObmbcgm6h58kc2AwDOt1Bae+YmXF3qiswIPcqZ2bT5nLhly3JAS7CLUGoHxwwOUXO5
uGkkvjd4BuN0b6lC38thZ00QeO7qcWkIq+o6oEa5IkX89OH/+WbR0CJpGeE5jgcIkded5G4iadys
K8Nb/E+PivCsxgF8erj07nB20MHdnqV8ShImiNlc4ksQafkiau2LB2yI5V7YbtmGWrez1PJ49Tnp
B5SCvVDqcmtv4mGVQpCaqUnqQLb7SSB6swUm9uzeccH67gnrEa1/Nzyt3EKHj5VcQlk59KuoU/53
tRw8Y3ALKcBY7CUvDDEsgBTatoE/v2Bl4hq80Wj9Ejv4TAIGD5zab2pBRESoHq3OoYUxR3khuziL
M6Z50Kw7PTBHv2pGMwzRWxzxZJeR6W2bwXiggiU8Pqb1i9DqZU5sSEGwxhYqYaloqjimE7XU3MI8
TM5zVyhB2XOgOmoIYo0dwAI7g0lPxlQRL/1cFD0bP7u88cy2vAH2SBVQPd1Yuir+Kc1ylIPZGZZU
1qUXUGS6lvcbonC3udgB//9nxJSD1YM13OBiLV5Zlt0QiGQOAwwaf9vjDlR0FDaSaKGyGkWEJXCh
zhK3ONCfmNneUQN5P/GSdtyU09C5+5ukpLLINr2xuC9cNXnPDjfMGyXbAt1/M0Uv2RK0nDYJsNVt
ZhLLw1Ftx8ZBtSxa9Hf8VNy/044d3FtBtba4kki/f/AZL4iTFcc8I8kFvbDMytPeCTvJos+hBwDt
Ld+SSE1R2P4kWZg2kqsR9KbeLMu95NxW35vCe9RRbpLZJbU0Co2wat0ovxoZTjZn4YJaKS2NytVu
JwzOQCUvihSFa1NLYN6RDrHNAsSStv5m7FtUcVNVm9uKS937ppufq+aTbTi0U2LMZJBCZ71Di83Q
qyJDBVaiqbjlDavAnejKqiwjhQAwbxAqbdkeVcs+wzUjtNrDG54fIL7j2Pj5OWjXutJYA+PSnBeh
qozZMsdwk3MIVHJkCr7OtDaDSNaimMQP+wIgEppZ+nRth0G7L0GDfoPG/tDmuTik/iz21K2CNyQb
gNOBsZIaDCV89LkVwQDuW0gJGf9d2EBZuMpNK10AU/lEPCRYBH7W0QR6S2YTaGMV9UjutCLyBLj7
q6bkI306E2YZhjgyu29U6O0QevespGeUy58ENfqmkHB4DcoX+/wS52pn0TzTLJwYJ4vxzSZF+gWx
pPNvgJIiKFMiFlyY5dNNxq4tOZ6Z6+4zv/BE0wGU7ktXAytVuJZUwjvdl9blLM9eZvoHb6FKltJO
prKc49YlOmQVoaejPald0tx0WvDjwb6hToKxR/+iqZkiHS6vT1DXBKmnxOPrgmqYFagM2VISlCNV
lPn2LcrL3PBn17MCLAAi5wqTjTeBEwXMn3RhfRd0ePtpPBnDJIZ0EbQSJZiwZgD8EU9i66ITKBJT
HfJJkU1fCHzzrcI7D5NK6V99kwNoc88bOKJ/4bKY4embXUhJVEx1BKMm//7ORaLoqPSKyMSjiRog
+0/rzzh8FOM817xx1C2ounEaTBLIk/ilQ8vMgdkb5JZVQVABM5lkrtgxcqqjls7NlC1ewtAo07Go
bLE1qPSEdRAXEHSgqewprl3arhVUSlkKM6u9vvVZZ5xmeB2roSTJxg56kOcJ28I/s+EwvGF6Dk/O
qao7Khd/Fw3DiUZxT+R/n/T5oxoxMoV6Un9htkJV+UKoasj0/5LeqwixRxFFjHjjkEPSdRRAKt4i
lYfjMOBwlJPXqsMZHbZk8bLZW8fqyNPbtFvLJI57PBwM/uVvDVxORcEOy1gnpkINwQ65g6hwUgRG
3VsObMM0HkFUtxGse7ljUYGxjFogU6kL5b+tkgvGK3bzUopeqxJr6LHVZhAtNes0Gf4h/ulp/sOs
K+5wvd2ZdOsDvHuFaf+DjQlSCfrEGVVkS/F6KbHxpT25GzHM8iUzmc9B2VYz8emkhLOfgftKfo1I
3R6I40pfpwAC2b2vOWfwtf0/cRvaa5sfKGFmOKZRuOE+lxDAK2N7synI25aH0HXPmrHcfvvI56t4
3oKRaNWYcn8yNaGRM5OTr7IES53AJGDzyzyIHpg1WRUu9gtT3bINOGpyqY36W1pMqfSO//PEEpC9
5AxyqJ/5AgTPgHdyuU9zsgqlMlPeNSOsEjYlk+664WmPh5DEzCFgsCKb8qLWVFQDb7tXnRXx9Tgh
Ueex8CoOCZ/UBlfSdI1pNhRZfy5DEOmkFctQZPa75vOWf8JlQcqBniJQkW4ti/qvHScmAn+rtW82
aVVzsgHcjw2Bj91ayvCVGmNRiiqlMSSscMzp39vj6exgdLgbl6c3074TqMtxVjli9WtFbHL1BYD0
VNkPkply9sZG/buTHbctyzQPZBttad/jyT0IHdVBf9ud0oEFDPtdINIL2inu8CQ7bkj0b/T2xIdZ
ovd9nPdsBtQKv4IcItpEeNNsBQNmtQdfXJz77Wef5/kczVWgz/YB2oQUlpTdFwvSWrNZyJ8e0/OJ
hzm0g3Iw7SFCUDu5Oop5BzPLGeFjqxOsVi20WJ3U7AZM7mkFMtc8mWkm3OkGKLjLESIAs0baILBM
t6Z3FQh/ORWP7kQVDoYRPAshHh2PmnwChTDtPOfg+Xxqpx/kDXhoTt0et+TxDk+VxnVHaxLTcCVa
LodKU2ZPiuCOzJcvqk+PaLkbCL0bHnaPM89aA2YlrTUHa/ijoJpL+bnSbWo8CFV0Efnf+ZyZhYyS
TVr3m0/qE6x6wqlFfyEJCShx3pbJkdbFes5VVelFJCzDVVZb3B0ij62eo1YmokQdKBMhKKMhgrNt
7gileqcbEZMAEz/BvdbLSw8m1mRJCApfHPFPLdmyW/BxqaN+YnNNEdNbnQsDI30nTjs+OL+6GAa/
Rorud7thDIuaLwhQ9fli4WoILcW8XqR37dsqbRXdkpcAK7YYyP5dkmAdYEJgppGHCxQdv0CBgv3m
uDEv5S6LnRWDl3hmsNeTgmCD3eYWVZlzOKK6PUsTveFMqYfY69blI1KelMn3ZqmK2aKTyOrXBOvd
/k+fA5G5LhzmaYDYEMioPVN8SgSbnHAv3Qm9NQk3E/gl9oL+41IIe3JnUUWnywudvpYjG/nvZe86
LVgnTslqvtc/DNHthikn1K/kSv1QzIGzYZRv/N0WbqWhsfzzhTUHW78Kz2ifX889Oe+F2s6W45/8
aJfsxKaCrQlKoGwPI5K3dJocO9rr+nqP6jaCQ2Vu1qToskKybSGBF+HPMi5zFVz6v963K6VOb47H
4Z/2WLl+/YJqgfE0lLj5QQRdVIl3lVqQ0c0uTv9YST6442zDfk2fqH23px/SR1awXFaKPOq240ys
g6chGT+5jsVlDmE3dUR/1fvvkznOB3eMPZvLaUTefVSZL5w2UHgOod4qmETypi3ZFfhUOlH/5xoN
AY07VUHdpb7e1Mg3fs05KpWuyUQVHvKEJ21c8xyOum3/P9g70ytiA30oWdxke3eB7ma06z6ZrkvC
JJsGJq4xjYmpTFw6+xlTO2ePFYvSnHhJg201TckZPPXULzIqmsTF/n8o4AODBADoWaHBeSzin6r3
iLIjrnijOjvFJiGNjz/7Su8AtQhgo+iwjaIlX1zTSG2tjZ2y+QoOOqsGmtFKSWvF2q1Fid+fO0HQ
m+SbPkBAydvC9K3a5AGrmF1fGsW9aExqKyTxEspicvhPHNo7tZ15x2OPM9T2LMehHHR7zW/IikKN
wYPFAuDT1R9GV/imoDr6REL28YiAYoszI4csiSsFbDOzj5X6bLyIcO6cvvtewLJI6fI1xCjCYBL7
qhjjJ1/HjWZqIgPYyiX/BU61pNUXrszndoE+jUpNAOovsG5rHYVTXuoMVZSl+fEtMAYTYCmFgl+e
BzzrWyUxXOhFvckvvf30UunO8czs3YZlTLhafn5/Z+B1fLX1nqz2ExMDxQUWZwLUkMyn98kWSuxS
VDtWrI2LWhYBsRgchnyzNlImL92K39jF+X4BUG67VlKAl+Jj+UWMTiTbe+iiuWKKfmhN+eQZAyb1
Nm55nA8i3AGHy9/Yh2g7OMQEoVxZPlfklNgVL66e1NlkZSRgVTKqhexXad7xq6EkGJvkVLW+rPmC
FBVvbTReeQNnJXjMplqXTMOZCfjfCZVLtPmqibyMnlLdk5DxLseZpkZLZZESASqgasDgIH3MzPqV
s71UtVozHdsh9JwrYocP7+OST31dQhCBZ9JTC9YPu4G4GN2Ec8ixOabrTzyAUbPRZIG0NUl8hfBR
zItV71dFKHPuZdf4T9b5YLzVfF1NMj/SDxtY1GxvNDIWUXZa02XV7L21CTdHpA8dkBfiqXBpVKh9
VD++p3cU1vWzzc2iuv5GJzkpsPmv7h80rUD8XKmXrD6MGIbeDBoKYyapsTDw979Lx4sdwnw92pIM
SjBfYo443Utn79oGyJSJBICwI1RwgDFrFwtJL5wdoiQ2vn2guokC7BPV4N3qVQw5TSh0y5746lLz
qxaBePboaUcWAYFOko1GHThO0A7g1WNcAs6ItiJEMZufKo2S1heSnpY3sPdHfWja8tG/iv0C18hk
QRQ6rJt6dOh/VkibBOJR0GOJLiUnCtghzTLZA1ZKhKE6MXtKxOW2ivF6QGtcHXPvppLvcDgn8S6e
LBf2ZAR2GFTEheFMuFFCTOgHNYfOrFfn8bPkqGepWWFiLyEiIDARBuRR44NR92noBHMM00FiPDDk
WJJjdEvrz/YsdBNfEHSQiLkQQSleZlS/hn+PW+Pkx9f4TOGrXNppkaVklSva45yRLZ/INxRUacII
rHMEDFvkeif/tgzHKpSQrrsGL/QzQOeLEz1J3TWkIg7FtomI10a33Mm1L0E1Kpoq9wCkjIu/TJtT
uh2naEIRSeloUDYbbClD0dwDy3No5p9J0NnsPRHNke1TDsWc9mIyEQgAiFuRiWxt7jpeIdjWBM0Q
fwXs30wekhn9V2vRLDdeM8J8n1lNUFWTW5oUR4mjphKKbodcGXz2u1DHl7AEMVmn/VhdfRlnNItk
1U13h7j9BjvdoXfmQbXfwI1+LXFxgKgKK8YNPp9YOJzFXmph1FZH/pjFrY3gmKN7+rNJdkqv6wWg
HmzLWMBQivT1CrLVID2EyaK/Zq8Gn+nR2JFuFEfEijjt77pBw/zWmvXrSaOz3b6fjzBq8FCETyK8
ULdwNFuzzF8N1Fn79Az0n8Db3uEQK1zeuMs+5LkchEXiCjc/ovieiR0p9LSMVEAgh2vpdM2oKPiq
MINVrTAxOfS42EQ1kY92siYKwLRFQm+2wRuaGv1FhlRG/LhlK8Zr90ha2O21oPo7Ow8WtpzuNoce
Zs4zaBiy1jUq1R2LLD8/JIkWqxXFZqB9M70BPk5kjyuWz8k44yCkUZlXoQ/wGo7RXzPTc0Bs+27d
2oyVAAfw5s61xYFmcUCs1FpekU1DkqAC7VXBJL0Z+iO+ecL/fGwr2pw0MWskepRvIEGwvU48KIHY
Vn6NXuEE2LxhDx1PAspljzLoAo4REMfPG84S10lKGPyOc/JWZzsB2urEkLgaH4RP7HWx5DUDsFuD
UL2DPoDeTq71i2OPonadzo3DWZ2DTYJ4dwnhSbebNmj9TP2is3UxJ+nh/b85N2euuDNVJZXPR8z2
l3k3a/hvLtmStVjpweW7wh6Uke69litoXU+gAS/vmxTtIpkwjpK9LtHMOpu9t6CWAvl3UOV7eP/B
SS0S6AL/i4yCc13AlvrVO2Gi7XmxQpu/y7z8vuLfXyzD20SB9X4cGbPdTsAMGbTTPRMJz2vU8RkP
uuaOjiuPBIcjXcsNE/u/bnv0OpsvDvpbswvcNB30dj55GRXoKN1fp/upJZJeNtuDNdi+h3U1rQ9L
LvX22ZbKNuzFONIpBx/IlC6rhAPVuSsd2cWpPRarA4jB2JcisjUAFKp0BaFFyw4qNx8WqyhOEWyz
3xpc+2hcm0vTKfKyaP4L2+PuqgGev4OMyGR/N9rU7ypwt0KrTZi3ivIcnFT/tcIi0Fc32Dv3RtdI
1LAJXZPwJB8mRQ6qgsZJlKTxCmQ3FJhfw/viFhfMIx00qm4oN4lysbzBc3ibIUcCz1fr7jOn/a++
T4DSqLoYrwe5s4vTdUkF/Ui038silaNKh+AS1xBJlfyjg/d/fxi3i7cO4bzw55GfEY9BNmiYebnR
jze0k1x95Gov6Log4mSW7xwnIQH9wqS+x8V5xtYsRpqwH1obRZ/o/KsQZSbao4QmfDxo/8v04vU2
MK0QNpsB7pXsE5rzNt63HxGu0FedAj/vDXboeN1KTL/oNmPvUiw2mzZiaKn096eDw48CDno6PX5/
UVyf+CDXTwy8IjBUPAPWgFTeyvr6qihHKobUDy545ZkQSTObfS7ZWv+XIY2XlsvQwUjeaPksB3jg
JnGMJGDicFc4Ougsu9MKWUpUxfsxld7OxsYu7qbknbbZ01yiGX11DlmC9aeDtdtOuiBLguhh8yAI
9zbG8lG6ytWEaJq57YWXGYFUgdT9tsuFtQjogg1LRi073HWIeQ78j2qDVh4V2BNAQe0X7y+CslK6
rbw+MoWbBkD7ZG73mn0EVJ+7ajMbPeZyDhjAlTGSd2gxKqTwZE4lz5y2sk4y8N1n6YtoChZlL/qn
fmSwvt1aGZ79y+51wyZsd5JWCuHekYtkiW4jta3QtRrcr/FHHkrYIQh/ZL4ZOltBRth4FCuU55ZX
KrhTjsWE8u0AUQbliqrspbAxhg7Ey/vSQ0TPEdvCqSnFMzSRaaa9AbgAPrhkLPt0orNZUfadCf8J
rhInge6Y1f6TNEpcD6W0/WENeZsiaAZRe4GRW5+gTu96I2xVX1Bk9Ec7V1rrJxD+VBvuA4sawIv0
nE8WofA9EN4PRssEEYpDez+y/vegZ9I+U0YvWLh3cQxG2LAcdA9+9nJImoQuhRwGrycixpTQvU0W
D6//K3Pwirs5z6KKZODoSlsB4jizzT+dshZym267atxHs7KgFPQy6Zde2OaRq/43I3QMLVR9jv/9
ptYOrKodGZmHKswQtpi4xazUPVqpRlNF8qSbv/qeF0HUUiRCSROFj2AmZ1DY2ZMuYDdg459lboTN
XQaNkRzrha4ZxUy+7og0v8kOIx0f1Rz2ndkOq4gaBUh9wRN6ATeIsbivwljvUj40sRwEjlaTok13
albShPzCLHMBl4T01Bt8rysfE0M6eOXyy+4CuT/UQ4e6F8FIvnsTMk2IWWKllZllW0BtcDKIvr2c
Wq5DLpI5H5Dt7wmNsnzXmzku6eTTMr7mK+yPPaOBRQKl7gC0fgfiU3mRsMUF5Nb1NDls4MfnXddN
6zg1b+stGuXhcJj2GKsaKXpG/uMVYB18k1lxuPDORooack/Wca0IWxru42finSkzOvfMOJHWCtB7
z6JjjdsD7eDWcvYCS1mmXKyByQcT3raMqaVfWe5qg+t88u/78EtojfjK7eFdIjfPqQ5N89cQmSc0
CPCbW0knLl+X8saStjf/BMCwMocAkmyqFYSD+UoUCVE/VfBeNWr6Y1I6HgDnDAvSobSmuYG7tyaY
F6ICtRoMFFNdH7MjIppgEw1yVvLOA3sDaxnJM9dnQR825i672iNOgYQ3z1a+PALYtM4xdQoEVbxb
3osQdoyX3PzOA5fBYM2tFJeqVdF8F1HMSAHHXvuhWm9NvoiBEkvkHS1SmyrintwXqbNVHWjZzC/Z
YrdOIjyUn2MmgDcKQeo4G8o6I11G9uVjtmWtgSP4AqXEpBZ8qVme4uALyLzggLGDtdfjvIdJXGC9
CQHA116XAcH4mX1itLL8vZbKY9Nawy6TjfMi5wO4Gbv/K6HZlCJz2g1M2Pp13b7CYMMqubceq1L+
q5MY31gQWM3NGfz0x8DjGz9GD4Vfq9j/v9aANYL2UrxKbN9O4zM6Pel/RA7WGWYIxIZIBcECF/7P
c3SD0Ekj1GhXIGnkO/yZQhvteeBhSrLpa0XXOuJq1S6gLjcf4SeSRYbqNACan0TJ8iHhIaZwEqH9
tMEX45OE4RLbK8nK29aRtKq9sBivlq1ii/vqmCM7xNNfC+yc5y8bBDKAd50WoZmHiADYD9VFH8qc
OHxHsk9KNiqgigtsOPGR7PmMtD1LzLKbKse+Ehq2a2uii2dL72CS6bcikyfcgpVkYWCpkP4fgOUh
YqLZmN3ITnv3biUCnirSmRfAqs+oNvpacA2F3UH3h9ziOfHAEvpcGqrxRWZWYtJRg4CNsqEYcBRV
F7tp0KOPHBOxPhmoZ9Zj82CKXIYto0UOL7TNi5K1QVLOlD530U2/JKIQn1m4kRSh9JmrSWYqfwYz
A79dOoF2hJlBS+qscojWNfHAjPpUu2H047oJgBz8P2snEJjwqZ5TrNi7gcjmzhGyYLsrXUjQ4J9V
Qkm7hnoNKy2X0NqYo56ndG5CS47KNgmxWY24wlj6EqvYXxQsRJQNX8UctUANQhdrlVOEZBSiYy5G
LZzT3ypj2fNxqcqhfZZZLT+3MrdoH1IuMmtEe1f9UAkrV4L3Z3U6+luY6RJYlAfBdKMFpSWpNCIq
WbZek47Sl2RCASV8V97yjkmHI9E8mG/YqC3f6cAICthw5ODD42nC3S/wQqcEASq3evULcOJDuAA3
+bD2o63QNf7TvdfO0F69gN3/xKtAzk5k2He15Y6ezsRI1N4Awwgv5xlfPqUXj8X6/7uJXhPwyW9i
wBrA08Bo+9nxlEDjZ9XH/prLfDVNqGC/a/gIORXaURqHmWz4/zu3+G6Emgdis2rZS6/MFs7bWgc0
JQApeM2JbZy8HoW5D0Dx3yx6C2G+AK/WI6ndZANksno+oFuUp8mtocaeZ4DUyyeLPbIhGtIb0OlR
9/0jGGaSvT3aMU6TScUccq7iOUNS1LLHVYs/tc+zoeHH6k4+RyB+Dp60j6vNjmG37DcfnfoBxd3z
YZs9W4kqjqKx0u9pRmEK4ReJ12AWLzMm5881lxkV8JbKcE/poTC+Nid+yIlujZLVIVkY5u++Mi3e
2YfNAdp/YSLEAgdBQwxvpBUqjsPVhnMvoOd3a67uidR3ioZ+/cwLw0gk1tm1tLq+TSQoLoeXk1Py
EJl3qChEiS4xva/xr4QxZ01raZrGCiW8szw3wFbA8z37R3zbI3dfYkBFIBNvqc1sdJA5PdycPsV0
PFYh5RZkK+ivM9ApIaRJdXJSQMfZ/xdAZAca0PehFfCX7BvHMIbst8byVg2wAnotFCvHtuWhCA3P
vbcll9PZOSnLywXRcItNr6VEfXVEtUGjQcyWiMUlJD1hO74WmUeYyOrhhZRubrnImRhVeXWdZAru
vh3V1LHmZnyY/h22BHdvLsK7m2hTQDEKl9RRUit98oPSC4cDlKQeu5RWU9QFAVBleTzH6fkivKEP
+Fc6qm/pJBDyEe+/uBebCCi/k61qZKi/H6FWYrbIJjVt7BAGqB6Xca12v1hlAQ/uVFl5HPM4QThw
t+P0C3JQkAFoZn3jTbQA+GMpuKHWldXOYad6Ne6XIxek6NsrRoNGDrn6/836gAkXhCMguMJvGMem
AmICZSHlM5lEylHCZV7zJRBLgEsS90d9Q4c0uPqXuYlB7l8sVIISnM4RwcjBmWauhWVRI7++hBb3
Gudf6jOmd/ca02S6oKA05cy0hRR8DdmMDvtCVpGCfnIfZ+UekL24OYvNHVpofget4KpzVdRFxA3N
goyyg21AgeqX3cWeqG/Sem3FXkMlY9rihe9skmgoMoyBZd6SJ9EeuJJ71As5ljezU0/U8boJSJgq
o1u8lZqhgT8LlvaTaz1uGhWKrI5zbYSGyWiXyZLCLWtpn8QaqIsZK+B/znYmHFmIaBCIUCwwk+Wu
dWfwJJOEq0vdcVDJghJnMw59sI3nnX0m6F/8125iWQdwAk+t5sOAfiaDqe7+YOIXx2wihQAXU+23
iiLIFrjD3BdYivk46C2eXczAEEQfnH7RdFjVfxl00/PDCaZaLqqIB5M3l4azkw6t1bixRgn1KyDL
wy0ixrbOCIgrSyz8N9evF1e2qVuxDUCvsVq/liA/HlW9dLlAkV0+SYEipvsSOSPezVmUVKl0dMWy
ER7kUlJUvoiPCvHC17eQuQ+Q9OP7Ln9eOhf4Ni30K3cqhNqPF5/+l0j1kgJCxBLyeaL6t+F047rn
1VJbJA0UsOHm/XuQr878si40bFNRrivC/2xyhSGZUQ9fwh6LVQuVDollBoubvmkFlcFix68ozSiX
KJFWn48EX8b2bfbkRjPaEU+iAWrpsmxAejPXBL6X4kqELfkVUzMzkpah8C9zS7AFughVPYMhcECP
Q97rby9pgdpA2ujAH3H6Wnsi8tudf2YImmR2MrAYUDBBH8AFpWMuN+k172QMrhjHQsUtI6VvCvWy
4thavzf8DR0wzFhcjNBfaWwrRDazYXpHKf3hVSbg91CZHJ6yZrVaO6n34LpbaXzDJCdM3HS5oMGE
Tavjkihm+dAHTtbSdrtlc4CsrecS3YA1hnL/hlqN89kOhU4NRWHwswR5DiCTlMOcfm/bGbyWtAWo
C8A5YwOo3ciLk1aBkPhe89yDWpxvGciNNs3qfOB1IaWGwkaNTPe0PEtQoZ1v1cqq81ilm67yHaOa
mMBYRusdPTVpnvt2Z4yu3CQ2Xx4apSG8UT7m5mcMYsqQ2Wp9u/ciT9L03SW7sh5L/Id/oqL2IrCi
zwDb7+ji9zdS0VN2t/gDWoEak4q7Ux50RYntu0a1ZV6H8kLwY45jhB5UgmCVit2uNdWHMDO2tDG8
Y0OA36inNWNOCh3WsZTmqaMajCnJ55Wrn0IR+zApRZDl8qetk+iLp6F449x4ZGJO5yujgiousFD8
pr7vKsoEKYTBY7/NKPoPAhsjePsdeOlxUGmcijCBn1IZtcVEKqVXcd3aBhkNec6WNR2VaPXfMVBc
gIcIfvUQu1kOupEFKav06BV0o1mQjesPuRMfCsW7KvUYkJZ7gVdybC+HrbYEBgs8Ot55xFe2yd2P
aahzxI8dBrejNVHWWomU+Zu2BZJitB/1VK1lKdqrlcV7IjTn0RaOlVJI6BPd87JpRNS6FtRNQz6A
3kTCkLeDemxlsZIng9pXvf3aFpPtu5E7QU03Re4+n5LyIBs2FU4CnnQNRsoEUOZI8V7HjoGAhH3e
zNZTMiV65DlYTXMlrWtx+hIHb+DMAwAwjGpe0VnSnyoo77L60B4A2WDx1SHr8dr6O7au24J5EdhJ
nwxRIpwTgfcg5PnT1SlXZQOrl7brX9dPs0pGBKWmwX2o53OKB7bb84MqSs3z+aC8/I1Pa0M64SZM
yFwDTTuhX3lb74ofDPR9IpTSDrlFHxoUyAvUQNz52fAyaqSEqOunpzpOR2VHKX1yLODxygxiLDGy
K3mj2b0nKylSe71QG/zMe45ec+QyEISEQNwm3rrTjWLkLV3j7c/ymoz7ofWVE+9er8VxtGwfFlph
GhBu/M4fB4beJh8BRISygfcHf6mkBkGDNid/YvVpAJl12kvzbYtg3YYzSc0BbuJLlNKlZK7feg6h
/swrbqLu1e4K7UvkEPnJdNUSSXHqpSxAffIkU4TdkRPTK3mdGeK3EAZk4YrMYvlByuJ23K+8wbEm
kVyQXEwztD7pFbxQkdq2dUvO2d2U2ffhx6pvHRbI9YignLsTxt3AUXJ4NNWbdXBUs2apmdaU8cjs
k8fPX2cHhx4JOziVIWfr3Q9YzRzzdSBPMjlgiTPSWFhVXC5QSubrOqr/WmYKUVHnZ6vprg00BQjy
cipT4C41qsA6LLM03hD1oeOgrizg7NVmlNPjM6dvGIK+duc8MnktkvExy5/F3ygUfoNPl4PAZfiT
SxUIaRH5mMzrjsOaMjkzc2vV5Hmh36BwS4gp0CRn7H7/UFUGtRC6pmjCPR0U10K7lf4p+w/a8EL3
xtEZGByAM3TftF3jfCmOY98xCyEIE2Eu0Ue0y5N2/0EDfwiS0bmkFpIGt++7tKusrfn7EnXIUuUL
MdYbn7C1cGxHtO0cBmCw8lTsJquupVOTEEb0cQr3Zz0ilA43Of6GHWGMv4835I42wFB3vRDIwiPE
kr9j5DYUYgKkxZGLFAuS7F7IuDTGbhcvHV3s5AUtgmHe+FshgwVp+65ZXKPPQKc3LWiowBDeNO/b
90JO22ZoT3umLsdfO1sJFhSd/dcd2K94SuOC8Swh+/2hQkYfhsvBzTz3c8yVMnue2xo/NjQ7XK8/
liRQ9fjKq4Kmbx9U4QQsbqMCPP8reIzqWtDSKXVdRqo2sPvXjvYVgBRQgiYCwPQ7sMzoRcLNb5y6
lePwfdCEOT7mnb7/dp2tyX75bw12cBs5kHAW6gFlHaS1ATxAxGZTaRR+UsYdxnZ8QTKx+1ABQUDr
FOzNkvxpQs2ldUzzWtZ3CvElFx68Wa4A4G8Xng1g3SDl5L85UPXU2vfdSnW6oiGEuqXpt+d12yGu
I7CknjiDNySNnQnxUSN5JL+LIOP5x67d++xdvJNBfmjE1T8rAJkg1kbngQeaxn/Ti2FtovLCgwSj
k2q0A25R4IRlxaG8Qc74oJRNd+53ezdj8N8ehFnEL2hqYeoYKVx3EU14fLHoSePvG+vpRbrEJVis
P4JbeC+XL1HmkDVi/xL5oydxhrpQdbekgV1FzQJR9/18QqCVGCrQPy35UBP5qZI5RQpgirVzLtX+
LoEGWBSv3Q4LVeavS3peRmmgM/C+p+EKNKN9KzkqNY+bxpt/g65qLDOXCBnbzG6EeN4rxEeCc1Vt
jSbEGg/3rB9djmbdZrtmrlT8tiqU2oZdozwgWKFGFjlVcG2cvYIoYeeLNEuQBFN+wsEyZVYdpMDr
bWmQasxjVOU6yU1D2V8ARjpywmHw3IePqubpVWNRw10C2jMe7vZzpjmVEXZeD4vUahkivCVPEoqK
w9EEK3xGXYX97yA61zr9dGqVH2sMeKlgoWKZZDrj8Gjz3NuC7YaL6WJ+GQzH/awho+NsmEmDfToA
DOet8d01wiF6ZpMMo4r9mcZCIvybBfDrQyrMCbpO27R0vIOUnnRSd0TFtaRlpAf6wb9KGwSTbyJ9
P8nCr6lEDaHoaMoIgaspHhgTOh3QLwUXsJo4aRX+tYvSoHkAxMw0sWKiN4Ji0+PcxdY+pp7boaXz
mzeooPcF1gPFkjgEc1S7hUabYPhhVZNvAXkYI/iTw11rMlrOs19VdFiz8ClGZk2r4XH+acnsnjHM
MinzmFGRxach6divK/0APP5P4zYlWm8nBL/XJ+8N0OQq5bDefcZHsPPW7yDNodXHdH2M+MLVQLGz
mlCqzhiE7P+6wbp6XsEFLnJpWEWBadVjYjjjZPkB6Ktp4GbGtrx8dYGVxEKex+J2/5RNlLm//Kfa
8RZVpHAE4xK4iU4shKzrITvfoEdewJw04vgXn+SWzLYs6gAHgHkDGYjBIJSzaC+zNnTfaNury8J7
3lLjbGnKk12jfvfeutfNZ+Yy7lFohjtEZiQ2fOdR7eb2bcjVAj9+Weqj7j8MUeBha9JCR53HLJvb
QUp0br6JYwfnHY6wbelYuJEttwaePOjVbhbbo9N5G5is/xgpe17xtZcrYtTIdfpH4OfSt8fEd76E
zJA3teud9rm5YpX/yO9eIMNBwWGycn6ViBmegOQM0cuLfEvmmSam3c/w2f5wlf/9ugg7MRrCBK/o
DXhpN0xcrjw1WMi0LhyEIc++McGzXlowNlN1Y/dfZAa3srWLfYKJJuUUmMW2U8+bVloEYBsWhKs8
DvmoBV8b2abrP8cRrJG4l+D4n6xiMgMpBc1i3N0tg8eQR0UukLwDax+2i+NNedSamVk3jbNHUmWP
nP8c8u5V6S9b8sZlIn3Tbb4lP6Dvu/tRVjCl6qG3erX83GNmYm7qD1sUuPBG1n18N84M3ug24WUU
ge+0BeNPU/31mHa6E576WDnWBoB+dpsp17IksHzYqviwoxrQEjkv2bL++zgAgPbiZN7ZBc6zqqf0
SVFEUTAv2jmXWiItz0O8dbafOqNVgUmkF7zmV+3dNw/cr/W3UZvFq+L6ska+hC2a4+56TffK6rvQ
mvKWwLDjw32zWMY+5aIAtNO3vKqrO0bkPB2A2X9O9cWiLxBwSIyQshOgrXt1RgzZjzZxv5JlPprU
b/osuv6YhEzvDbffFID39SkcvO+t8PuGpJPo3iIt7CqA4rAoLCtVUNG8U7g0s6cX511AJCt9tIwO
r/AU42YgqS6Tk5ShCkfFWm663hy4o8PswXYBmzPS9GWacTFt3Kv1qdDWkPGrkuiDdPg2PHnjtII8
+5udsPGEex55DuH9J/Ys//GwOW91wP1uKdCX65yJyOfKjgy80bj/j+MXcHVTYF24sT/8Gq2GmgoD
my5FLHSSTQvMmn0rFcqY9yjkhxQfWqU1ZAM29oGL6wUX6s0oxLaJyWoipND4jZUUn7gxPNVRsIuL
CWZLB6hgozcoxVLHXtQqCpb1CkllL8c9QsRT7+28ufUKS9A+qnwCIRoMEdJdhKvtf6WQf7cxEZeL
azozr9xROY5KQAX4vL9+SufnvUfCQ6ZqNbcCCBnAmVzTH9HcQyRHligkg2LPKI725c5Rf+eqAo68
XYt/6K5a/sMzE04/r1y+cT1AWh9jZ/ai9TMC0KN6GQPkpLZ2Dp0t3pdHOHTyGb2/Kwv5019A8ya9
WXpakSPsf2EZFT3DLesXbWCSPhisTPMxfS2RwaHuJ7ERX6/dY2DBURMbow8lF8Aw5LH3KZmscz14
YFDSmp4+2drufx1109o5nd5RcN3PTv/5inILKbvIm4w2N/Z1SIkuUyTwDorfqbCcN5pBaU3ED/w1
VluZOIkgcJtN+er43VgaPl6S3rSyo5kWbW7VD+QxQlBOcORhIJt/zIsvmP6iqrQz6wdVKyzDH2Ok
ghMaZKN/XDrR07IUbJ9i+q/UcAAcbpwqClA70SJjzbg3L2Vm3Phc80S0XA6p6dugZRSbRW7B1f/i
h6oVsOCkqhDirasaJvsEoiSwENqFSDhoE4VtS6BXGptJSTFrAe7XfSGhh1N9FzNGi66yOCPJowEA
bksmjGH4PD3Q3HUscd19FXctx5Y5miAl49CfpRaM3yJQ9NitRJHZKm2q8zGR8m8//OoQRgOuCp/o
1oGrqwLl9n8r4O7+yEleQ1Q2Tk5esG4rVawJrkD5OQc95JMTEp/iSLcF370lDdJDlk7lNrT1GmqU
1keFE3ttmpdXd7NPKr5b3Dn53jvJF5g0TE11dO7l8T3vq5iWcVvY11FaiXsEnIeyFHzIEhdVEmXs
cZ7Pwn4NHxszL3kI9ylddvsRM58xzWDz4g3oZhANCmF+OJavFLapT2D5CYDi3lA2PYmMwTG4m6Um
Ji/ndd/Z8frEQiWn94+7aZBXS71E8Ty0ikAwGUeXGdaD+OdnhQv3hMv1kYm1056VZ+uiOT77Wf6K
f+mR0fA/x5ZCpWwlzMHB0Oesg8YK5rPH8D7Cas913KvFWhUDLBslvtXYrMKBzwaNpO+5Z4Urkjzu
yHRAlqHGfsBsUQKOOfNA88TqTSQbrxBKN6dR3uuoS7b7ZLZ6befoj0/qJYRXXNQ/GAwcrmWLX7ra
r+nGw7Vc+JNj+Gh2NTO0th4kWbvuLrw4AELscODKZy/KfapJKOPAS3nzHRkitKBWvyf7kyku3cmu
HkvpNbtKw7CUEsLif2xi0PYWpjXMpn9s/d6a+GGBdNVVWYqqXXfczULZUvV+EjnrO8nDy2SCDY1L
eHXt9Crlev65ruNOBgB7l5jao/UfCxCozq/4/GBvH8AsWxvQBc3wvNJYFh8N//JMfzAiT7AgMs7f
BywP1NPZsekfMcxIvxpEIMMcjrbwn2wr50v6O3WABOjHkxXOt/TWw1U70sBMyc0hYuDhmcVOfUw7
H3vNzApHtYjzmuonvLleZs630ApOi1gaahc+NVVPkj085ih8lUlhssQdRPv7JTNUcCaKuqbK/rVF
C/rceg+TO0t/flG4UyVPTx6x+xETJc97hFgErbCOi6eqV0yxgJ2rqYavOZP+0XGaUHzWGurH6IKz
vZEtHxiS7mRqIY2mH19dHg1d2Pc/8Abp+Rb/9P3Oo1JafzWs5TEKWR0fbzNoKU2+UdS30k49RIZ9
IR7DtldcW7CqZ2I7Aj1ExY0uDOFPwBfQjg4SohFHrJKGBxI0DpMVH7uLXL6XNDMSeN6qxsORjDO4
WntzEeTJ9Mg7SlSc91E62kw4tXnk/8rZP5/9JxGK9JPbwhvIKboISp2nIo4dVvY9dqLMYxgtcVNu
kkotmrvqS6isoVN2SaUe4KvVFezMpXUl1bu3e5Srn1+I1SB0zrVsRSBUBZde+/JUoTh2FtshMKHD
2MDBla4YgPhXLG3diUosYx9sob+kImx/1aNzYHzlmbVb/n6g+trwBWRZ/vQPa84d0BnX6z6Zpq8b
Y39C5/SZBi2o7gnjwI2jk8coteQ6cR9Qmnh9U3KstPCWLd0+SZ2gZLjQgzIRYUGwIMmH+6J/8tN+
hgUMUIHR/Og9PvxBhh+tjTgLEh/88Kzg05ksE8/nOZLUvrr7cJeeQZLruqIj+QESW0bEcA21DJiq
1tJdJdQazF8BpPrAZtZ1itl8+qeO31hOjTL3GW5T546I9zGjRdy4mFnGpldropHB3bRbvPgnU6wb
JiZPBDCsGUcmInpVwWEoICwT8Z6iJ2r9fdyo1r4KaxiW1/R2HJasgfb48htRD/SKyUY6o5vAgKc/
SvQp557l2XSKunRwvggHySRkaP9+nbs2EJ1KnL/FG1OozPoqMjCcVCCYDmxzE93/1tdu/S2tivYd
B4XbLHRMHFFdufN6AnnSc+tF1p2zFsahfiQa0x/fQR3L1GZZqRnB19De3lEZKfCNJwmc+wRhKDNb
rZigOIqW3qj+M0j3OEKsq20rNTg2FuaaiGsxxAPJCO/nCfqPU5oF8KB/c2RBg/GfX+P60r/QZkY4
Y4vpehQj5tKiIVwl65DCZTZDMvYMlGFfbA3VMiQgHTfC9KzHZD4k+RfCZca0WSGeY2dNqo1mXa7e
ywwuyR/oabhBRdLtE/JHGrulWmTzjQfi8lpyDs5++S4C880YKAcwLg07OpJDWxOrwjBWafpQzG6o
kp912cwXazgjfkmgn+iBtiMmi5HVbnUKK70OOxSkA6q/HEGOOrrpYCHAP5c2FuVDCHlBmKfa6fQ/
oMJFGdl4ZQxwmvpct0cnPEQSatsrCvEnQwx0x1pqbH9fEPf/KQ4i6TtcbhJWT1r+z4RXjPpfvERj
DHbrZ94ZrO5SVJkmzsdMmcZu4uGbYYd/hAGcd0fi5lAgv4k1Twbq9yrMnkk9hTVQSmOz7CMx/7BZ
Ukg90zxtmrKcY2cg7DJUDNSmDMUAG139bKXRij1nyj5F0Noa/NfVN8Qu0EspDTEUnT5aMwFvpnUs
u/kSkZZToOjCGS1F+wmO7k6TjhwHjbdZWxmr38xSZIaVSp890hAW2zg5F+DBDkmPAqLg0GeCdeRV
yrhpHElXdIshA7mTMJoiCq0qWvBLo4a+X8EzQEyoGb3J+dqMlRiaMMOqCzTlOQURx8TYNueyrjut
x04/YF+oNrMIpQWbErW50qZ4gzr1nyOPIHy8JZJ8/QnAuP4umPhREWdUhvIrB/hoBn1VLuTiC3z6
Wg3xSs5zVvUqOmWytm9hoHFwr4IZpRC/HUVg6LFrLRoHLz7oExGYB683kwyXnhgJ19o0SfxL9jOM
VIDWJFOoL/5dfp4x8WY7Amvpt8+GJ1SwQWZ6edcXFLrz8OrqIvNha6TTjq5sXdi8noupXjFt5dD2
petI7P8Zpdt9Y3yAckV/7BCcxdw7oUtgOHYOlVFcOK+RAJpGtRBcUjbzKqyjorECJbl7vUwKGBKE
v8JPnGeJURvAbOibb0/ZrtkuykViQZP81rUqQN178DYzPOnB77GFRCUa6WDsDI7iftanJcyjfc0t
rognyI53Lydv69l8q1uaqb8pA6NeDKuob40Ac05upQo0DVj/dHi26rt3oq/1C4NMgzw90FHe7/hn
7mj+Y+fEyxy9UbErZwGCYE1PmRRHz8Jl/FEy9ySavM9B6QVaQ2mgnvcItTf+chvs48LSBq9h6WOh
IcaciW6znejojitOqTyoUj3AcfD99QnfgR8nnnXHnT4W0KL+I2rLvIvTbSGTziZYG28FKNbyCsX8
Bl9e1JLIw+/82NOeqXKkqg0gOVKn2HJjUvR98FaoY1gNMaBqnhdHIHknRfPFi/pZqb7NFl7wNLR7
nk68z/79kSEmWUXc8gFn05xkcOlnpajr8O9vbg5TrI0Atw4VuetTtCcfsBgrbn1okAytTwTMpIXv
3+7bPWBU8G8PlZ0ivIhLSDs1YuneYXSq1gv+Jy5qNR8ufbr6AgXcKKsGYwZFdfnfEETSgStXXFbS
bozZgvHVaVwIJ4e1rnGtjY7bZKzavd5K5MRBdXQ4ExIyVxqrKwfPJTL+WY2cL7iphYqtvBFV+SGH
wl/4EKFxFOhX/L7o8IXtU10mA8NsECJr4ADunxPei9b/lCpcQgVAexjXwuyAg5pH5B+v9rQ06z/D
I21ExZWZpOW/E0MgWXq5A/dzb5Lccpzjc00UH4koCR5mJpbq5wi0BHF7DFuh/U/XnLDUFI8lcdm2
UQoUS+p9i7qHTXFdL/tW7R7QYf2SYhoJ9TegwKPIvNv9iAFGei7mqX/K1xHXlrafgIVAUgBHS/hl
LLpEhnIBvhg07r4CvpzM/h+QdVqX5tp8uWCyW5ENOUlLVlq+/mY0SOTvcLxbBDNPM9/gtil6sOJf
6PcLTJvWuIW9calJAMBD90GmItYlyoKE5beGY6XkL0k3ZDqtl5tbU1XakOUj7MHow4uw5I8AOaf+
2CjgIwAAkK1b0Qsa9MloBhBlIow2ETbwv2OLzatjYeWtHAZXH09rag8xdulUVEp+TvWA/ocAmfOL
Y22AgNQlacsUKBki1aJEWyA50t0sUMrcx2UKaFpH4kDh+Vsr3nW7I8rsFQ46bJwX67yu4cfdZGjG
JGkVMKT/ruXNCIxbmceRVx98vTgtjXHZoeaW54k2l59aQ0ooLqre8uYcUnYKZwDtGKdHjRGQBaNz
LwQWTQQeCsQOfhOv0h/CCLIahufvF5hzJxdGtfHwCn8QK2W6zpxRk3jPWFhaZ7Ze9882ROc+qCR4
WWqtM2S7jJMojhMSc+mexrKThVB/367HvpBLG61Oy1OvbSAiOdpMZ/igYunlzQBRSWK50bgTYvAE
pByCzeHbJynrNyYmW7L1Z9bXxf2C8CvsdnkMlH765eorsmPfgURNShYNQTq199TA+mleScs+Y+8m
N8V8+FLuAImRqe/LZuR+RJg7uifeBUSAmmY0TveiJlOW2lhKAEHRFAX/wXY2XC8J4X829WJxwzwC
WJM19lzi+SjhMSvSDWxfPRCDW/TOrE9CgUks8gVCONgZIvqih1/z95ql6IM81qROu+0Xp4hUft+W
HhxeQKVycrrkLPowWme3KS3L669otr/02pomq/SOqQbY84HVHvE8NytHlbuTEYZmaAyp461ythve
vzsU2G/x/+UfkslXOY9vyKaML744xTqOvnvI5tV6kSKYszoMsDg39A9LVJdsUOXxaiTFahmqt8/L
IBm9Yx2MvvuS31sd1zYpSmMpA2zPH44Kvb6YXe33n6FESjgbJ9aWICatssCPSdU2agLGjAxZDYAP
YVyr7hwizG1zV9eG56hZ89Liy2ghGLqN4b+hbkOWcETzrqfffBxVeITVjdLNva9UOKOAcoHpBR+Z
+iHY1sI7phx7xtMxZOUUL8yIVfs3p7dSdsYj/1JR/5ywagv4zL+pEaM8No8gPF9hEhIShB67ZOME
JGlqPI0/OgeNf1YuvEGVMGO7C+m96TF9vUF3RI96FK/NuN+W+bVh2b3I5n+vBh+Kk8e7/IUhy3ev
1l5qKsIDWqIQG1N5OsjYxP7FVCAIb6EUV8wSt5ricwCGB+rIRlBsmYmnpM+FzU4eLoyZ66gcDzDy
3wsKXRZWniromQYZh1TQV8dPgLrE9CMFTOS9PmJJJLmi+7D7aB2r0xJIAsicPTbUuFCHwr44Csug
gMR7+b9U/kiYYUs1ytv2QSilvoEozqOiTYt+E0M1oEOC9oUsCO3TuIftF2S2rQ1kxxrul3EPGv9L
B5VgJkcHaJKJX3Kbzpo9amCPSzZKIC30ZN5A3KmLd1mO2E6q4qAxMsa603BJZVeiT64zgogVd5on
gJ0CR8iCfXSGEOcpLff1Ec0p/0slo9T6X25kFRy+OoB1/q84SJbOKqQt7RNEKxbjtODmxJ0GMj1+
jue1HZUgFW3tKkd6ndOs3NnbcNi8m7C2juUg1shv4G03tN3k7Bl1CQ51cEu7SNyYNrTGRm8PJld9
Ro9zBpgwM90dH+ELM87eRYp9zKTiGowDce3FJfQ1hHbJed3MQTlChC7THtkaiK4MrdAMrnsDtSzv
DiHFGp6UZsuS9zM3NbBSVlSO92ZQ7Dpvdr9m0ndhv9qCgDaAbUcPZyJTTzijKk1m4l8yhJFO/s8z
Qp9cv2b4lsWXuDSc7KzOE9P07VGbK+VfZ3IyvQ3QeWTW9miInDJmPzBdVnVJkW1a2Zu5tMQBjo15
OsUuY4h0InWskeZqCUWLCUrCDx5AUAACBKG8JFkeSy1lScr84w7WHjWOkIIKBx8VRLKtl+kYvZiA
7jykfdj6F7KnanMJEhQH5StU3bzrFm6HAvjDrdWbSwa1L+++C006rnc3JhAgXWuISdbQzw2SN8vA
oeXP8/H0BNBG2g4RBsOnPFDdjEGGUC5krCgd9IcdOYJeow3RqvmODRIRFE4C4ZXNyl9i6Pe7Lgjp
Kiqpu4efs2nMGtlZZKZ+KKkHTryJ67Uqfjw3OlaAiEhSrTkimxXthukrebAskCh2EvktA/m2nZMt
AEkRSARs9qiXXZLPgTDUTTuls88YAQXzkxcmhe2LF4hQb5YW4ioNxvZxu/CoupaiDCs7k17RKBnL
VU+Beh3qsM7H6dT3THB8T8u9iR1GVlxhJaJJVbU/v9k70EnMx4HwgB+Bmfd4hJ+EiSaD3+55xJED
tfJw4P8tMnsbcxYv0XLNcuPADdSOzfhXwcAIuuT3qgWEp78HEn9OrnHqY+/KplJ3VWYDIrfqJZGB
SSdGVfom6f5AaPNGlhTa2ZHmIK22hNWppVDLzEUu1v23KlR18XhjQeUWqKUgg0RckM6Ut3VTPB12
4uY41Gi51Rphn650EYPQYhAHuQ7mMuTkYeuPvAOmCT9Mv6kLkLttCqFu2OMTWRdvZUXotKvgrU1B
AAl3CQrZ72IFPnfsPRtwtu1Ul2GSUWNmUVGWu/8qveeLsPGme3W9ZvS2zpxZZcgl56r/nCMg4wvz
RLA833rNM4Yc75jXhhdR5+TRBIF5WfMEL7MJQIyW59QXQvjZGFjseeXxUoDxMzrKGo9bCL1PqEYE
jFc9SanZmV8EjakAObbeb22yvogIEGIJX00EEqPKkpNW1NIRijvdFrgxVkIWX02l4NlN0SgddcjJ
KkYpk0yvsyDmBvE6xtbAPIo5+yfGuipKRd7ZszHEODFYLtRZunBMj8LLz7IWn+mA0WBm1/sMv4Gj
xG7zqEElsRDul03LokYP/FmgeXCHGYGLijlTfjgysjfLuK6/zxB7wePZYIioVxM81MpEBWJLUEAX
PSyipFoJehYBrxJifGA/mtAyfSDbSDDG72WKYyB4H/W9J/9mHVqeTsxJf5Ht9Pl3HJiUf9ndtFcW
10ZvVHPoeLT9cZdS8VwYoBp3Cfoxg0BSczapLDRWBqo9xGcBy+e8RHns1mtRozOV94OPXgryBY+G
Le6ETu/Z+oHKbbEyMA0+8sHzuh2huLxPE+32nnBvxDNxqMglNQXgfZIQCVacfsFHfqyAXWzKBaRl
nKjHlh9hKAPYJc6wCyBQJLuG9KDM4xbZI+qeg9L+ExRB2ggJ6Ox05LptI/1dWTC9ckxtlI2xxFh0
H65NdHGVe9wOw2Hqxkk8aqDeylTv7TmSGiw38ygOPqC/H4LCNxWItLJFvPB/4HBuKh0WTNY50rfc
KQuRnCKgdwgxzEwoPMKYERXXg6pmcpM0de8g085/pNCbEKxTilRqSWzScYY+QkU++pie3ensuhAQ
clXUuTFI38LUGIUcYagP6en5oBpFev6Zfw1Zo+L8dslC0bQnAaCrdmdqCkg4o2TFgxxwRUZ1hiMR
vzi5YG9UsOsykgMRBVSNrHmQAWV6MQxSMh8Eg/jbQgtz6GMwQRSmWrZJSolqzp0BCQWDxcs6UK8b
XntfUtRMoIoJjlAHMVu/AuuxM4ePkXQ9nE0X9U/4XOtnZFb8XVsKWVE2BxQJCiT1L4WUrcts2Hnv
UFrW5L0mnoS+N+joIrFNAmzHKNurBLpgTE8EFv2Gr51RcvyUTVG5EGTwuvtCSgi0gQkb8wCAn9MW
YZ59xGj1V4faYTnOyImpvJBNQOPssLA73eDZS3DAC6wL/XBzbInFHWJ28M6T23BhE7W5Z8N0Fhc6
nN0s7tWLzcBP4FyerHCagKP6+3FrPEtqf03TKTcJf8Pyq+nZXstQ7UhmI+sL+6BwhcwjlEwgkAMu
lwuTfG7fmyOH8YY7ePSiV+pedP8JwctQvm5V9w4EPZt8dAJby0vR9KXUw00Jh5wRi7DEVDp7th5N
uTejyqPTfuU+J8BE4A4znrgpjNUBD92OxA+yfJYGAhX+vPndJoq5T65bRFeDtlXW5oWKyNEia/Ug
wIQc7J0p0Q7UGXxsS4el8ziyHTnE997AID2BqQpMp2Cba62T/cl7PYfR+/3QqSKbocWuKUHEJWEJ
PG8htcjWIMWAgLHkA2/cdCVaDl+rc9i0t/sPa74BA+8ah67HDhxTeGJpopTyn7ESvRYHRxU8mDBP
f5MswGzIw8fNDMz0j9hlfCbd3D5QN0bMQOVHfmSRceV5Z/JqMf7Wy4OtXCuq+xnqRAkJfNYG2tCD
Sl9alvWpXJUyc6Q6hJiEndwaBBiWDAqzmY+hnmVaoQTxKF/a9gZU2nmdAEBTBnnrj36aHnfBKP9A
JkKw93MciplyZaaQtd7KCb9YeOiVKo6jXmZPpIicWKQu0eFMHq/XqMqhTdEJdQszGl0duvQML106
MW/aKaJCU238RBidDOajGQQOdc1W+YH3Wi9bdFMmSI6mF+aam0RR5U4Qqhqxv2gf1hUS87BhJ8gv
hq3FIzlRAxLfTmiqrSWSAVc7Vo5RLnwgbQ3OdGXCpXBkjxitmRJalr6wNgFRyQ/5RqY8xcZLIhQQ
qn3GTgqt9nKbZ6JBoMAMwOArn/GdkMnjk/x33nm2PkOO/J3ZTJyKpgZ758ezV/k3L1EponB4vKt4
HACyKsEM2NWjPxX907dIJKKhFDTcdqhe+1bbctVGW9KtpmSerx07mLNQV22pjsEcF7IAxlyF4etz
W3/Ol8H35NQwbnWZWOUtIyiXX2ykxOdBR+qwNGhFZFieDXJBK37PN3/5Wv5C10dz9MHixKb7j6rV
FL3ppN6HNxJTncWdutQpGj9Jw8qyEFe8hqpBomjtXwItxi76xRYHa7P5fX9qG1KJsN4LQU5eqm83
+LDlZ3YrFmFGgTI8Qi/ar1ZF+lS1Uzlhgrh7yVJ8ARufTtFgQJfY2/BLb5Z/AF83JKYKxtlhQve8
zRCkogiqvpDBemdFT+Z140UVlKKLQFLBDMXltrnT675lCWpoaiFp8mKkeneEhHGUcObFrhZY8mLX
BGaB/aeb2i4YDiuWK0KFBBi6DRaUKvAONMdfuARVY4Pcpa5kpuYEU5JWYxgwKi/sgftZLnSiUl4Z
7I9e6RNQ+YLQEpP4etUy4rOJz8ML2MEJpkXElJWuWoLgiK71xC/291w9OaXyMtptbcCYJwfqrQhx
ZQdfoMSx0Pjs/6MMIr0pCodRLrkE5y6dUQO5UdQR8StPbOgyNINIjGis79TV9+RtkRSJ0Ip/houY
NWoFef+6DZDrBC0vOLo9frwIGIJKN+2GLi63yirQiuSoOM1ndgcijJack2vDPIJ1BgrcqnE0Q7wz
EysGR/eEU2SdpgaytmlUQeyxQYJK68541ZVB6zHDXx5ouRr3iGVUHHihLvkkQdBrR6h0GuvyI9jB
nj/+qClezSVjr2vZcoeEZSsAihaBoSXcFE4YDUr2WbVYLeAJ9lZ0S7AD3tKMNvIA7D2EBlpB7+R9
k9TlBmVx0a0Y5AW7X+3ytOioiLUD9NTve/r9oX+bSEFdsVgR9rpmPmLT54xC/2Wf20yw46w9QS/h
nrkHY9Rnk33OzcCQpVcQEdjzcqcwEJz/PsNq5aYoZbtDAvk+oyNpuL/O9/XKSVQZmSM9gfICk4S1
VEIQHx8P3VYnLEw8PdNZsOLdvJWtTm8ndOIOuKnfNZXnIqCljwRf3T/EnlJHPA7StzMZyvAPMat8
7itSeSH7g8f5IMLUQpHnMqDuxOHHOCDzwakbzTH1RXAFAgUk6vZ+3eSZl26LzyL2/woTc/11cMtY
RvNCQAX+kOQwd8NqpqeLnhlB99iF1WH2hf6qT5e+544MNCR8AbgsVAJwUMobWbcFZa7ZF5tE3bXv
rv8XX7cAzVW4sbRNcqz9lvc+NqNs76IFM7TooA+6yastjzrKJm9PE92n70gnsaFYwsLa5gzN53c9
J29XTSK3u4rk3oa4SJWUvY5sC7vcT/FdpVe6X904qy4q298tyflQO6/oWoZIvMhJESn59YFOREiV
DaXAoxErymsJt13r8AhOf7zMgC1RYe+N/iF1ADiAy/W+zsWzbyMi18GuPqWypjnq0vo5MmaThwDm
C+JH+o7tsx51gqW0pfY+95uQsDU9NyMfMOWkd7Aiwii0i2zkQ8pmMSGIoF/waIqed7a1yWMvLStB
WZNP41O+R3k5t1DvXrJcKixsVYaxO9MLWg03+awpwWQ74IidccgAasmBUzQutOlrE9wKvF9KRv2d
0qHWqNl1K2Z/ab+F28nVIYIzoskGqu7+OyxsnPZE+Cfs0HhgChD4wVbNanD8eW1LcelTOxVhJ07t
dpY1ZcKmjKZaop3LN2bbbw0c22qD+WOgxkEOmaaA/dlBW9GtHrc96PmCcmbH6mrBkBbktvrBy+O5
g1spQzhAWuyH0vORpxCa59dOoJusAkRX+CLBq6LTPBQCIfBC3NmKtgrvP4HYQdPZCrRJpX420OcW
fcJ8t77FMIfS4l9uMl4YRu1MKceGhxBAbD8rwYj46ixcrStzz37LZgLiO5RZsyNmJW+ObOjG5WmE
QFiFrTq8+/6Ml/2C19Fr7I17xkzmbKiwgvhcJOQ6bHjAA1QFx8B9WlLkWIGr8jMcLbYaffdkHWXO
42LB1NRJsUiUT/U71co+WEVpcpPzJE0lpq+2AT+JNUEajQSqatMtwBSBfOzVf589wkYMchCF817n
lwOtRgC2+f5JGXBgQizyelTQPUedEhvPhXNXwy3dJhx8I3PrWvC69pZ4vG5byMfiAa/69W/6Gw2o
+Kd5EpEIT2dtv8XfcvFXxbq+0Ukr2Qq9+k8crP9aMNhqUKfUoBM1kgXwuzziX6so4eQfI7o8rfTF
PVURB6XF2BjUCrFUn1YOyJ0ChQI9w2KbnRbOX9Ghw6sSMS1kak5627ptpRqM9XyPv05oth6jiDa+
dM6sjk3N0ZJZBZAhZIu6NnsuEcGgcp2w3IWW0me1GZDXtXZm7HcMetAYhjvyhXQhNY2u52nm3GD+
Q1YOeO6jQ4Of+fdnvODFdwJHQgDnanpLrkfMTa6DvK2X4YL/u8RBKinXdIabjLJ7OIyS9uiZu4KX
DRv0n1mOGGHFsLAEWyUaIXuRWaN+q+eLixZaIUojSfSIZW2W0R5K0gk0/H+qWhi/WRq1ME3HWKpH
mXLvTimj69tGws2Lv1SPof1zGVvObqWHigsGVwawhMo609fsOc61/EEu7BcalmrHHqZAy3u8qooK
ADoO9CaTTzr4gN72i3SwOoGzyx/9vcXHa/XbabLEDH9wE5EL9eD2bhoWbWw5Pj99IF/sUhJe3RPg
W/rrQyQQ1VdJPNUYmv24GiIINg78SWrFqPP/RC8Yee1LBQgJcaYCZTQu3HtgAlKnDJtsXyvQ8e7Y
KXaFfIia9vEAXRauW08Y9D0Y37PQDyT0qxH/YWHtidQv7BYNvUuqWwhLSGGqLhCNPb1a5GMrqhvt
bfn2CL7S0f0PyzN3tuorSOQQiEldXmYxAaYF16nbuvXOSvHbCZDsNkKxIjvXAqeTAzYg6fFbIMeA
jiyD/oIlqB9pieTLQkVR2GJM9a5ENNw8mi0OA2FcBGRjHvBROgbKHjv6nh5tlH2SfGeBvIkdXX+u
JEdXmB4VV8FlIJzNceoD5Hz2nDdtvcCm3jgXLomiowhO/kSDCMsFHLzeUpYZqcIkxWjF4tRysRX5
mPqP/Rc6r/NpmkS14fzaEcV8TjxFEgfPOWBJeAYxB+47q1Db/OrJleO7LU0gwUqIFI/EpGqWgQBw
YjUBFvx5F2CVnHKbI5twoTTF4e+FGp/QXnXpenZoENhjNeEKd3xXSmhpDetMShVG5QCY6ULA3Itj
cgVSUzdUNp8W9/3TR3frzeVE/1wBTR6Kr+nnRY2CtH+0wwtY5WPgJY9rUUWh8ttITnY2FRDR38fD
9KZ6QpdGI4JK0kgdAvOuqwP/oJMXrtfxxDGCA62FU6LpZYKccLjBfX4Bv5rPoWI5EtNfM5v7s5oe
+O55INUoBB6otArwzSJndfjN+RxmYccr4xGWzq3vZPd/oe/amzxRP+RfvSSRZFdHiIu2KRnoiUsJ
ylcVthC3OmSlR1pVs9nteWQrHKqmrctnqveICCYZYdBw6gmBrWUa2zP7qIehzLV0yl/e7dzOa2TI
ZxYY1IDTSHLZizOiTGSdGQUOz59MVkmGcmtDCWU7uAZdlEuXW5gw/8EXexIljLmdfiSHNej3kuCm
9mdZY0yrDQNpJBK8uvYJd9mAAB00kABbSW5SMxAs/Vy0JVuNe1fnIdSJ39YDSqf1HX50eTtSPzcV
Hs+kmg22I0gVEfW6uTuEzKhxOGGi2xMHj/R3rr8ovYmGlQqDXJXfV6sjoD+cx7LdRB1u5x7B937m
J1PFm7yVxGuZSJmy80lOrAnyjBte7kiR/KxlMG1RFlBvdmLM1iw3Ey2YRRTHUKX4FG3YOsRqy7Qf
IUPeF3x2UG/c0idrfE8e8hFogAeyTK3ovLIqS0z1hrDRR16ZVOfOiWbIJwqUtjhSWS9C5zUPAcfY
MJhGMwonvgT8UTroCRjPQ26JEvIQ38uGm4ef8/iLp9q7rS6gKnaHIxJyiTdwMTYnnh2rdBbDFaYA
I8eq+3dHKdzjEa3BHXOTBAObMY4BekxUdPsdT/ZNIuX9B10PeAO7EkwzTeZkc7Us6oYTqE4CAqBe
zH1X7432v4XZo15RNKsHeXuwL3Btzv5AyoigL4uPSxGslnKljXadgJGbrk9EAO+O/wTY4+YoJqWl
THDT3hsSz79eOxGQBr7dAOq7TObOYWMu0QdtDnRzlFURRKmP/8MWv41v8y6weZEgLRqKSatDVpL3
rWsgQDP5pnbDGbI57YjIxB0cnYXURS91CHvNNRKApFNz+vDC11IixUp8PxoW0Ka+WpEkkM32seL4
L2WPMoiW1qbQl5nv5Py6Iq876anCunLvWsWHpV7aFooHmINnQE905w086cIKgPNY9NuzSW2FUKWe
E/mSQTNyEvIJRgzxHSwXlxcFCC2wzgFQt9/rYkL6P+dn02xwSiaWXeDOubDJW8DyEgY9pK/LqfZ9
8HNVr0JSgtUdmRyLTluEZvlpKBHF3pMtJdCiAJU3VStzx9BskSBMZz303B97N3++IRQUVShT1j5I
QOsM8csIyOp0YsFc5JHo3tcM0IdyoatLIruWWTg+TepzFHAVpR2M21nX59j7j4Dju8bb0XsqYPRT
u/LnVQnlbxSusPBbvo+ZNxBxSBRL46cJGdH7LcY3Wz1zWC1P34ykRUUtYchyJvZbyWzMgiPMKxZa
V4s8kHHLTJKiNlhz7FNZtrx50FDxpEfieRaSqDYV8SkWYfo87AlaqsUKru4p2bYyzeyONLZPiTra
d0tNqoI2pRSIb1vcN86tqSXo1jXdPt5NFYHT6xuD9fAT1MerZbmBkR9SJrt4twAse7MC38UoY6Ii
qxbIJSiyVd81y7qAkZI5bnN8ZMo9asTPhUdxBcMZUNh+vx116eSSyJ0rnxDDwZ4yUxfEm3GxXC18
pEdv8NtkmbXWzDXnNLnulRe2LIut79nvHuDMQYVmZEIXs+OFCY77mAdLBMybbWMkXV3sLyu1g9/Q
tz3zFQFaBLiBkn4wOWF3f+wGYdMC5b+F3rxBTeO1JUI5HprDyJg+d5IoLCRCp0o0PWwOuPDopHci
UK5CxyqMJMKFTq3vK2qAV1htkYDuGnyX4OgmIg9kwN2xh5ogF9l0d0pg72GaV/kStsuxM6ITZoJ3
OdISXUxr9LT20eBK++qp4G6VsW3atRFiWv5vDIVN/dZPtuSNBdDlpYFIgDEODnk19lYZBi1INTlN
Z6fXSZ9pRq5m02x/bd8BRQYZAnEN+gxq4EQKxUkellR6M1faQb1FB0zJ1a/nt08+LqPfKdl4Ou52
IaeZbg/rMmDmRHfHIfgSysoWI6AoD40IxQiZnnvdg88oDhtDfbjjaRmmilQ6pbk2lUKm7SNxbbED
8ikSGRENRvyCG79U+/aozeYVAzCV6V+jXf/IaBsc13xFhVklNhAy6cZahS+o+e306ZeM5HsimR3j
sJe6a9xCaSLIhmbkjftFYX6BZzX5kVP1G7k1eAr759sJgS26theh55CeViCF4QADUoxXWQnPxd6R
NwGcFjkQXK8MaC9DGSXFEvIj+aZfPoFIrtTzj8L9F9aW5LKXuklig4aLop/MAA9+Su0RwaA3HtkI
w5Iddhyqfb8wQRjJegWRbZIzTefYBzpc5+0RwN62jI+aKYcrnQBz+FU5slbptPegV3urmsOYcpxA
17EH7bkzguWYhLcNPDX1McoMzbFfF45tM+vXGAIf34ShuA5bFGk2kdg7vxejkjwdqoVAi0tycQn3
Vf7k9cw7q4R+nD9fYylybRzQA1K3YgXtT/2Zi7xcHuAQFAcSRk9p8T3tbeNRH4JeDQE8k6tniBoQ
ehFmgHiqy1/8aBTTtGVVIsHl+0WQfUDcx3Oy7thcxnRTlNXUzAlamwlOcelrdmxgazMUdzX15Oif
kGsi4Ox7KyBnCx91R3eRj8mrsvRBz+H/RQHcNlbI8a7I7VETPr1fPf8TD2hU+VxOt2g4K5yJ4iKT
ZXoIKQwsM6QbDZg96XxNfyALAwfZBw37q2tpAG2Vs/jT+AWYj7/qyDGaLEgaMdifx63Vw8SPLEGV
bfH4qz+TjH3q+/R3D9Bbc/p+cZ4pATE/iZDffA8OWNZMlfUm0gfc9CWb/q3ZKa3ForxLvQ25EZ0h
ZgMCEWLE46ef3KQcMhibCkRc3AAEBxcteOEnZI3AeyAAoRTEpbe2EB279QK7DfvQXwEV9smMNtks
U7N+u+A615Tf7kDAfcAcCpXI9NbZZFgzQ1QFmqdfSOGMbNd2DHBf2hso4bbzEwScIVAHtKfNhDQ8
5iNslXnijaYP+p08O9kFK3qXOFNglxS38HU/djN5q/55DiEzizfzl6Hzv0mrcJ62Iy6CUE0Wbp3s
00Pnp5FnbthuGoQLlp6hkQ0KprTzxcxgbBf4IZcMMBZ60nG4+piOk2s3UHTqbdk7GvPi7peMifPq
O//DbrrULY9IKebiDEWALFv2UbkqPugyxr7vBvafUO2QQofKs6vvIgjYosZRbNHcuFZb8MG8Z5KM
sH6dR2ixdzXS90oyaunR+ZrIn2mGCi5pwoQXDT1s7fBEOLNh5URBXXfcSk4ogVsDICN6s8x6MVAR
eMMIqFb8Kipe19tTbEluUQH1Qepxy2LQrE8mjYbEKJaicSFwasVdZPXGuIM+pBuGVh/C1WQZaSDx
vKRlCSGhIgIF/iu4UPnD7ZNpby+19eQAwFSL57zLpsxSZntFbyA4WMaqVmO5xFrPAXwFEY/GQYsO
X1RAdCTKUFWo7ADUoDXMKwrad6GDtDxCcy6U8diXxlYhz7mVqYvGOq1Rt9CyA2q5wR4ZnOhbEKyN
Kkdr+E8KXzvtn0DibfCz2q0zghgZiuGiaq4wvh7aO5HI4vxrqMDgS1i8JtOTxtm2dekZVeLldpJA
14J0MSVEBEnQmetezuc5i0jPiKCIgSAPHhXE7re/n2HkLmjTIIV2jSdnrMIppEi6CAJEPHWsZ5Lr
/iqo1plg1/btbvYcEd+y2YrZDDktxKCI4rq5A4qS4FQcb6VQ8QhOjjrT3yY4zpOHGt1pLNDYE580
aYWy51gs3zC/5DWt3g0jheWtq9vn7l9vaV/n9w1bYZQGOU8YNmAwHQF3Eivota0bvuOrDrS4niV9
hnS36on2e3W3Jy2PiQ/5F98ns/Tt0N3PoTud36ENrrH0V851hJSiC0eEiqeXRplDP2WyyM1ToUoH
S6IUsxaecViT8NuWhD+ZAmJIX2BOq9jGDwBQ3SPGjsocd4tK/2A03mLTk6uT4ccVI14QONUvAmuj
V46WUaKjnZq3loSZ9PCnhzBxR++M7NwtrBUI5TwSSuxjMF9EpKGzPCx8DC2QAw==
`protect end_protected

