

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FZWxslbw+U6Wgup1K8ZmbZ8ZvAwEdSXoQX5Zxu+YDpvGpSAvyJJdij56SPMVKmhf+X7kxMgvbsEm
5B5AiAyVHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ntA4Op0vLLt6gLQbdMxO+e0Bhjub4O0zQAgtU7SVthNE2o/5St+SvTkDoJ1ve5MFs/Rgt4JL1gtd
IBaLjbwdyEGV2JKFzmLfNOLgk4U4bgeRTGAx1e+I5wKQlcq6qarG8xv4yuzAX6jRFWecgDUKdkZr
uIZCcXBmuErGbIdhFKI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I/9QBkeb84dQg6xWUGWLN64S2R+IIBcNXAJuDMwqYLTsejjUFtntzi/OgGH9xu74CzmvMnJuiSkZ
p7NF+AufXfE0LUxVeYNmvB8UnCKeswDMIWMuVEpX3XPk8OVFRqBWCRJ5c38XRjldLuPPEii8dq/d
MjasuPQowI9n5pgL7s7SczhrYfNu0A0XEQTAwaUPGij8aO4+LpdeoyqZwdg7p9EXJlysFsw3bvdq
qHiouBqf7MqPbKppmCVMlrH1R0q5YlTlllFEZblTUq4IO2ZWi+5zgGnEERNaNBZQ/na3tnrwOTGu
mqAR/EaIPbn2R/AR26ZYNuBuu0Ym5XtWJuqzJg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jRGmdT13qAzfiT1K2NPIFkj82nI6QO0hHDoQ7U+cF5NSt11k+3KuVBnDKOWta7RjBJSeiJs3q5WV
MSQx2R9/yJGRUjq6DQS8PVF7sqUyuFjNc8w4wdPwxcG0hsCFj/tEGyFHTU90BhMVIeVjf2WlERXd
+UzGn82C1ATZxC/M3Bo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c66DzsXEGPMNOrzYyBeymw4AV+RpL9x7eTO9Hf3l3y/JxC1wwEbipw1XtleybcrcOfKY/ACDBUVi
s9qFxHBAPyb46Eh9l7EGLGzxXJTWMed4eJI910mZ+WMPkBgIF1jvUqr1JGStUHDdUjBjqP5Bbe3m
2g3HBNLeS+8Ciq924vg/jBwWCA+G1zUvjlqI48sc1XMFszL+AzQf3r5t6tBvdkd9goSPiuISrM7C
eaSWriX/kCtr9jogh2EYVx1Ud4JT59uRVRlS338jlkF39xoR0AXtgdhjpZa3Qu6PtAnEwyq9aWWk
FBo+MHknw9HNH3v+t/wWSpyyW9f8/AhQrF1o5g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12512)
`protect data_block
Rpo3wppsiM9HUzfYFWEz4xQgk/Y1V+qa4ogILkOLomXb/Go9TJCGjyWm6CbBp4MSeKelF0K6dcb1
LV/3oOQ8f0EKEYxPZg416FflsXJJFu2j7htTDh0Rw7FVzjP9y/h903lJNwQwDAau4SdnN2BTY98Q
MHV5lUu3IiXykZ7IdBQCBDWHWqMwvHC+l0LvQI3Bkx5oM8dBaRqVSj5ZsSK4TINdLTbgaPCmQ4IQ
6txKcs8YymbvLYTgPuSYTuIh14BsCmmQdzfhJUtS7pfG7usIAg2EUsDF69+XVleu9t2A7Vh408sa
VzAmUYYmbhIej2Fod5YY5aSJ6Lox1/GI7Lnm05lIw1HM/pSz0sKfkGrOQPgujHhULV53pBn79C53
u748VvVbn6XSQi8nllrkJ/IUwT7yOhf+u7X3P9JhlIpQXgZwcpxs2cALtV1zNWq3j/olH67ZqeXh
3hJv0gvszB9XAmJSHRIJDq+fkk5LkXbfJnFTh4koUHJ0Zh9hcrJmc1hlqLUCxZ9j/SXn7URIuNab
/SpQPgJsS7oABouunsT9sggWp6swKtse1HWUdhYClR8FJ6PzZuXCw7FYAaeWtqrfxzMhZ66pKWen
qRwfK9ve+GQhAh2nQ7Ky9EFaSVBbPsJ3D+92c26Sn0zee0w8rSowBezAPRI5x9lWsro+PkmN0Qdz
vqU15V4KqX0sa+4RK19+FgQK7hDd4BqzJTXjjNkOc3dx54PzXkTF5x5lbWioKV2lgoYFBQsKBzlm
9v3MlV+fxtJGp3L/RY5nPEwWe+X2P86Gq0qAKq9DD9ELgye+9lb32MdqQA0vSsWigPYIlDoiXIY+
ONGaZNXFuTBVR0oWQCtU0nc3rZtpvKFVH5NvHPvfZwzLt1rl6fidycQ85BxuOneO8lIrOUiJlImS
6H2BpwbPdj1jS9DaAlFqAqhJyJSwqgFAeNesxzTPLjO7LQ92LzbmZMeqwVvVgQaYqvSzPi4MZsNl
cro7lnP9wfXxf7lZ1CFLzhBM7FFfHaUBfAcuWzpWtXltUkPAkqlZjdBm5/mmV32+qklpAStxenxV
fD2M8janZgMSAAbfuPf33gQ9ODINUqyWfVRzD3MCN1xLjtEbMsXPcUhq4yxUBbVeeNX15cHE0xDU
fUVhJpzQQyqwRyo4FjZkqWthyxHON18GGlcbVGGhwZaLAvixDRIDvCRwVXZ7ihwY21Bj05QVpEMB
rGZHLiYm1iWdErjVmeHgDxZ8DcapZkV+J93r5lKltjyw4/icPmycDnoHGp8xFkwL6Tm18ppyYowZ
Bf4CLRLIomzokUA9HZlSczEmFjzheoeMU0Yr1QbT3eK17tG62PM0SbH2pjdA34s+L1QjRoXNK87H
PDjSLaKq3ktliyVsM1XqJi6hexkLFqeyDpDXghwwnOcgX1ATO0qF1mg9gcSKg+UHRAz8N2Q9YpTl
0+eAtzqom399T9ouh8EJz6MBwtEflErClTOyENYQ6TNM18O0l8oMnixTHmiQ3wSrPiOHWAiSkJuY
LWef9rY1EITGfRQrKeVVMdgjP6FjEkCyCb55O1n7tDLWxPPhZkaYJDNFDT70/dUG/RV/yux07Ki8
3tKpfUodGkGlDt4uo/QK+NtSTpwIFOM8ljeN0IljwexaeLKQoDDI1JQR+Pburdbg+8VCoCoM5QlU
megIS5wTzble8G0Nbbg1rIp8URExUsXDH6y6XzDHjBDiO6yc6QNet0kNPEaqYsAhuFGs9rC3Lj2z
YSOPi4Gb9yn41uld0TNV6IbKrtxDM5PgCfoIp7YhouF0vjWFnM05U+NUba08F0l7nnZfs3Q7Yagp
sjx07lVrzRr6d4KAVlpc1sCAr7zVT4eiXCDR2s//79O/fFw+L4leZq5VTKnsF9jygQ7A3YI2A8t2
h5ttO26BrUcjIRAdLyGpJVFvG6kbInb/Uvug65UzxPxZThSO1KFAfAHo9GhTfgoKBZljWPpq14p7
Ar6P6lXna2XuPmT3rBqCXl0PMEnmeho3/182khl46MkjO31KB4lmUwlfs1yf/j6lXwBqrLm5Yo3o
kbSpEGH1TMrgg71HujXLQwLXbv6oCaMDd5p+rr+EfXGsjfcPx+9kMfCe5inqcCuBao42EbaMPsHA
Up98exrqjrydN7DPO6NGXhrKhK9SwQE5Hm17VBiLOPi7+qNSnry9axbjnpBv13CoFvrZCH7+xWHx
3NqcbcZvpqXxq/2A7eakwVfqYNlzElJ87XT8VaAinc2YRZ+6ooHYbPYDnXTYgNKyToQgRHBkZgfb
DUNO53zyxoUZaAKkZ37SpvB6tRR29FDGSmpCU8zKB1Takp5RfzHIuSHrnFFy+ScDMsCyq2cL2j1G
GtchYn++EpPQr/d+e4pmF3/+PYUgl6npdW+k+DYPYSMLxdAAjPK7v0qzK3ZWz71VpCwwQvdIb+sL
umu0N1lqzzBV9dIA80lNokoYs3G1p3dZ6a6ODZHVjFvv3XF5mK+2mRiDtExpgosbpuLllmQtrQDm
qEsNEx6xzECY5C+ONo1pZ/PhbPuYMPrDUuvQaXa6TMt4rXKNidFatZELNQRDR6i2JsYVA2ITOIVu
NYkqEwKx7iGiV5tJBTcoqhjt6aMKUAgE986aNrSM6pPWJh1kIQIDrYjB9DVo5R3c/mpfNkM9IxuZ
16NnGBSOTA96n6A2Hwrud07l6bPx29hIt9skD3mEVXKmT1tv0z+a8mxwF+UqBLXjZXXv4XbRVs4I
e7au0U3x3DC9X5KyuLM4mFN6GU/6u/zfHwunDXNVA8PQAhiUCF4D3Jyi02+ZqeIHBGyGUIBJLxOy
ldzF94/05qxKxnQbJ81ET/s4Kse93Y0yMq7sHaEoQb5HG6VwjvWwU6wLP5ngCJOmVqghCngHs6gR
ZP98Za/smsJw4u9eh4baRk7CzTvKHoIa6dIoATm88TL30DTHLLa7RTYlgn2yOJA+qdAqPKUxRVyW
JCkrOTKVGFkmk4dqwEdGv6yT/bLxchRp0iq3p8GrqX9vz+g4O0AqoPstl2X71ZyneFW5dMy6xccj
MdBIFlUzkHD2nqU388u1nUnMQnkAFFpdJgggQ+5/n1nqNTfgJRlVXrWRqbtmbpoHNbXyNkGib3R1
bOZfX6Ex/KmjkmOpBO5DcGJN8WHXMqrLaoA1c2Hq7tB5SsMas0Mz1sLZdzcuYcytzqVHVxJYEoKA
R35dZzeWgtXAoJvarNRAJT2mWhfN3mXJH9SwRXk3lalPMjOZyoI6kN+GLHYJD9prrKwi7TRnzmLX
g3tTIR/zbFeU21d1sGb1RJ+JZCwTnBl7HnXKwR4iCt79tYpimsL08l1bY8EHdtWGvUC81oHWe8cP
OF+ByosDbRZEy3rfTsTn0z4QY4QG2ksFO5djFk4QszkLjGnDQ5WvwEc3dMnR9SiINVhNvUXZEcyu
Uj2NABo1z73lpoy56lfpJkpN6O1varddhFILSgCLsQ8mXl9kBCc3I3VFAJEltp73m8uwXH7m8wxv
UPdbue8IJFqum0UaFBzhytjMURfXComnn42yoOuNkFkyrqUdGmJMMDXlSqorQgrfpVsB0feRx5CC
fzPcn1YOU9E/hEGxCX9jOgz4HEEdfcZ0htscPIT1CsZqLvqG1YfrcvJjf8dntckFChAW1819qVuI
UFQv37Bn/NWmkQEJ968VeUJOMSD3m8MQZaZR/U6dOpcecVcDXdpEBrrsvwzaEQep62hNBc2oQ8On
j5KE4Q/zfHF67vP5ovR4il8dFjoNqY4katj0f2s9zuZ7LEIrTEipa0fDMA3JJpPLXZo49q0vz1ZB
VV/8mTpPMfx16F9R9Yf/k8HDoE+d32AYtT5SxuBxpqSewLW1QOU26j37JGzXjnBoj8wXNGKv123H
7IH47RWzRrkGAGwbIxGpQsVwKCx3rfdYDf/qHtFOaG00+S7kCJxCfN8ZwFdhnUH+FbEkF8h3XdNi
lGWk5q6Pp/8EfcyKxH8LgNIwpGa6bnsF+n17jkoC61KHreKrNMS9ybJbXI1ZMvsEO2fL/dOFwzSR
ePFhVLYlkHDC270Mf+IMqRJwgyyyFuzes9svxlkgiE2mQLnMNDidUU8pdIVYIxLM1FHT5V5Ba6Or
e6RIqUovR34k468r2DPP+nuVivSOr9S+wHQxH665SOttaFqkWQmKRnIJ9xrzFCGnDlJFVyHzBce0
LqV1ZQeW6ODEsg5jX87tVSatlcAWjdZ6Fg0IwVjyDO60llUiw5RDVXh9UOgo150sYG/H9tBg0Bvq
s2uJHLCQhJVP0eB2WwhBzMOpsv9YADAH7rV6sI5HBlV7Evt3aPLe61c9IZzNH8KmOIi4xOSFBKWS
DImeUOafsmBGKg4SLP1PwgE2C9UZxMMv4qeZ58AjieOEINeSM2+X3kpZ0W6pe9QNxlnXgAIMNYyX
YOxJngbEl1oB+k/nyvUUbCW6IssIH1h2IJhveOW44TKbQjL6gF4feJl/KHio4JOoy4HzCjuF3UAa
YqWX+zuUp+E+XOvAePvgKFjDaVKtbs9OzZf1AxhfDIQ4u044qooiOjK+iZ5+ddiz2ALIB9Etqvzv
8oa9ZOGX8JNVtNa+kn3KZ8cMuKTdKrWAcoJm2aD1Yn0Ygy0ITrXnKGAKuQS0PKjEwzYXET8+tbD7
Y9KECLCSaVVFn6p6645IHAGXqEECABMHDT9r/7drxxE/uwVX9hiaXpYDvbO9Cx63vFyhmIXCXPb1
ARmwFQwAjGu0YtCbpjhagVVUp9kMW82p/aK6ao1VbMUFxxpUjam+MDLv1uEXKW7TYOLqFwCPL7Ww
XlwjLgnFe+/vQjdIJXZZZ7tZw/BuCu/GwPJrL1k85bH4vRloRBcIF/Xh3q/8s1Y/aM9C8Ypaau0p
xMchcbjx2wltaCebHFL/wpeZs3lu6iaosLQOrT2YzwQD8dnTHCq1khvC4FpQkA+Sa8njXnIxG1xl
kYLwmjUQhrfBnhSQNDDYhZYVuevm0TItu5iTHowUoOQTtyuBIKX39iyyi1qmznsThO5hW6/el5UA
AUckATwcfCoog2F+N2eMsIir79/RCk602568hPI0UiMZBIhWHKxqPcCJRz9UK5QBpFZLUQ1yh+N4
b3Dd0qbmeMOR31Izfnd3WzwfetDfWiGVvTRnoS6nXU/4IPSd4At2s3YoCTeLjegh98nZIv0LRPoU
WZaAYIT4NzpDwz13zaUYJ/FLM1Z/bsDXwAj99nJ+8VuDV52EaAfIEWcf7M0+zVnu23VWo9U7YiK2
zJ819kFw1s+by17X95cr69wGzqtQh0cGJpdIiGfXbv2CrcpT1AvOa2+6cbxyhiLBD73WMJiDJyiu
GtXYYOD4d8aV77jvsPTgzC24j1rLy69OhGdfG7K34fUiIfcwJVIEjniirnCeGdb7Vus+rz0mSkUM
w5E2MrpmTDu+0XLskxuocWvdFZ2DOj4+vP6dnff63g7i3TaSKvLtL5OJhQ7EYpNlnE3xkKVJKJGk
K7ZPkla18kgQ5RugoOlq7zUDx28PjL5ED++tBcjgDHpzFuugggs0KSF302g9VrC08PfMck57jxf/
bqEZTzu7EtzgM/xXpBUY2tSFB2WNXAc+rpPP7OfRLkbShKlgpJEi7KRov/bjG9bEALsaYIO3jZsJ
GFlIReYljF1jLKcF9VM8eA7ctcIZQ22yKkodSaoWEpQBpycdQjB7W+5ejXQM5HnM/bfPCP5OiGx2
R01BqpM4lhbazWT9VJmbtOSzn8Cz3BSNjHpbPl+wbOmSwqMz6L9Kl6Ndq1w8OREqiLemVgtD7MyJ
UKps3M7+M3E2O8oQl4GjT+IsyW8xH//B4tnmLUBOYIeRS1+/GLvqkl2fdCEDRZ/GOo0Zn4U0dPdP
wBVXBIr7xU9kAp/QrBhYXVxXs2UAvj8YaL+9WOawFpCGRwOtRUERjznzalQmRWHuT7t0auDtwTFv
FHz4E6XY2oOjb3oIFELWT3rgFl6ABPZl808apoVeyoUhQ0oHtmOqYcge9NRp11VeKXQd9svcnLlm
0pf3nSzIUAZMT16T4/llyNL6nzHfM94EDY6GoIjr+lS94Iwx5IwqNfG1LWCybbNdmVbm16AL9Zje
+u8/d+Fmyf/qS3fm0biUdzjSG9I+U6vHz+FxGv3JSs3m4Oc8OH3wfu8oqL1JJqGginERtZZ/i15z
rXqy/Led1JRzkAHcvpnm/TT73ZwQkjg4SiuWTIJzigKmRMWb//sJSxlumpiyfendMcIx/0d81ZvW
EHONmsLvn/trEdfNKPBHyaslnhRjbegewIrK5mZCALRAPhIjhaLX53Hwi2gNXEUkcgWJFTNoAsVH
+QTQaryBvW+zIpeNBWqBeJ/MKNHyhWmlXH5biYkDRiChGs47GxdatzJNfOHtV1XZFdlknodI8Mt9
fsTKayHJ0euDkQyeDX92YwABc8VX1J3FOsPKYaH/UXa1Oshds1KpADdAlAbx1Ru1vlRYOr4LOcpo
+1Ql2Mo5uuMCgCyIiAlgps2UnoQfoKOZ09hS9sAV2evh6OTAjNSfzkOd6EHBOtCnd1AvW0Vrfkzd
njb+cMHqypCz02c26knplzoq7ez8aZtsMNIWPbTqvffjH0aR11fxKwES+lckVSsksldz2I+I6h9Z
dxDU5bijIVsHLB3R88FlIUTs8sXEIgwIFnI7kP5fdpLlTVBiJma0saOUnBCWor31dGCm4Yl6IUud
AbIstHPOTbG/c8ouHeA3d8bIrfwhD5iGJjjhDOFMPJsWCX/YIQC09egWgI9c1kwZUUee/2j0/MdV
gsWjBfwuC1UTOEbLpxcMuGJzm10sAxILinIhv2rpvodH5N5efA8f4JudzYUD/NU+cR7xn2+mtX9i
a4ca4OR3ANCpBh7Fx4l2pAM+2seQqSMJVC6dFNLeSr4OToDKSU6Z+TePCytTvvibF1mah7Wg0AHS
QNhGCuCbLPycxGIMRQbcIyYdNy1Wa3e5n/1Rq2uC6CgFRy+F1dthKkbFVOGx/8XUQ7n2SWORNI/S
udvdyisvMW7tcQ9KeFrBTW4PPJeV8tOvoChI0RafDkPTzCPGB3ieGQJCVekZJjB4nPHsvzQJkWm2
K/ky81EvU0/+lHZfjmzo9oT9lMh/MnSzXjBOrO/2PaIG+6D5L7dWN07aK3y2IAYLPLbGEjTpzeEN
Rq+x2stcSuMkUaIUjXoGDf4x5yTQ7gqakiWDnNyRKTuo4Odk2nD69ec9OZOJYfr0i0g5/48fMDYp
gW1jXEYoj+hYKKcZx105D1ixiRH5tMvhxRaP3TB1wyS21dG32vJ8MUf5NYK4f1TCY324WXCtoJ5e
ZYCUAcXOVGjVTuLvh9TTKC+pQ5C1SZ3jl5WT1ej9EuzVX9Sw6dqJYj0zkDYAyd7KvYcqRqGWVVp+
Ql93xrm01N6PaiIjPT+YpioSTGvrYfduRZf98dPNsama95YkfoD020/6u8eaDs4xkS/+p8Spbio4
gPlVHtg2JQrQiIyyUYLon2WUwFGAYXvPft2kCXzX4zLXW9ErT9Ja/AGtjrflxx5EKkq8UOWrtk7f
HocVxsP4J4FUJfsSglFFQC8veF6O1zMrewK3Ztia1uepWVFjifK2ExFK8Qxq1P3Ax4je8/nbEeHW
MXCWtSRc4769/57oAq0MufOKt0hYPujwCz9/DfeGJlQBhAZoLgIRIqkg8s3Bjsis/Inq5g6dgkKb
3eCbsTdyDwMNt6jJ6DNGHMbgpFAWrAyvKNIo7SZLu7yIqVq0WkYlsLCFTidQvPoGgJorK5mcxi41
BRdnNvVEtGlQh9V2rYE3KfN/2QdaZzFPO+BiH8faDk+LKg0u2GG0SxCZJBABIvHDrxeWWx3GcKPq
IWvZM8Kp4wPuFRc3x1E2z2fdQ/7C+Tq4aRhVSDdFn7aCWVki1hBL3DOv+KWDNcyFX5UnSmu5ABQi
0xpXNgYPjymML3tpD+kr6TW/qBIYViy96uqGB6D/X071dDo/j+IzxIkw0UJcG2P/AnIZVfsTqFlq
31PGLbQxFidSGoXneE8uO83y6Zt3FKHIv8gNXwJLoIO8i6nc8kry0B5gh36spOADs/M5yhyzSTG0
uw7uKFOQudXhI/EvRaK6XruqmyLCpFMMQ7+Z1DgjjM7x2Sr7wHxeV/aBkC16dTLuhJGe/FiQ4QiM
DeHiczT2sI6nPwE1Xh+zsPQ/mLvzeH6ja28rVMMXLf7pnypBV6PFyGb69qZArW/U73I62kEYAVYD
0cUwUhsMh0UZs/eNqI6wxOvgfP6rr6IevpQQy9PqfZYkYSukhPqWGcYpsCM/FeDqYduDVBH7Qk4z
cOqyzhyfVQ2K4rzqNhg5pCv2iD7y0daMMRC2U++P2q0kzs33XCMSeC503b86L3iTqt3e6Be2JrWU
9YFktSMh4RW2FbPgLzEzWuVSlmZhLIB39TqjZGVi0gx7HjFfmm4OVhNaZrxz9D1xJFmiVl/uN/ur
3JC1Pe9PHQqqTQk7g2ml1ukBNFN6HbjMf3OrB5veuCeRiHXVo47Vgr99sQKDACttJ9kf92FTc+WW
TNdUb4EQSTWS4BCYgj6qQuosX67xFdKEGHoY0dWk8l1FkiOQQeeFY9KYT1CsimyrWsVedWNKPwei
cBZtBM6t+44yOusiCI91nGzWH3PW+qKuGMQEUM5mMVXxbLNnnNGsVfZStnlhb1aFqDkTd2SqOTSP
Vqd7Crec4iSscGOecq2ft5rpLDijrmQUsaV6kqTukDM8mzNpSxVCUcY0GNV18cF3nKK+6S8rkOA5
HF+yO4cqelrOdN777xIaidwtCZ6NI+bkKpldw4zRVZwjxUEDZh7jpahMl9aHjB+oeApTNY6QE74z
MLM2j6opKaXNqtHXogpfUjdHe2kqIwP1hZRSPRrS8+KCIFQxnM9/WV4D4iXJbpFvRunY1JLDmzbF
7T+sX45droblzs/VbULArk8VTQE0Ebb/zskAJ/UfEl3XDubMV17c5S1ysmzjK33FAkfAl7S+91uY
dvUly404KcUmGxwRgB+ZrvC0uJv6POlKB6hZETYu9+kxaeRLXdF/h9pduZ8Uz/GD61mjkyCq1Iw1
mv4CF1/HyAOCAbapYqEtBWqYndsHoYBZ+XqsVLw57WrAGFUKw47oHUz2Ibr+He1AY3b1ct0lOvJO
Nv+F+gwItUsOEGWQu6aKoiYfQFZXvqrZZX5kkUOh1Za6+gvCgFhj6ZRxE+wAJy7kb4UlrzXIVn/Y
hD/PNptaiHkZ8Ckmi9SlKnch0hEbAcmLl2OLlGQC/EsR9c+Xjppms2mBdkbodxVlsRSi9fkOHOaw
/X+fCAI1AWk3Th7svsVAAVbvPln4bcvcyw++WnD/vWMx3+ZqzR4hPvc/XeZaga10bugHkjWJzFZC
Kj6h7irwlSa0bBJrwoDptovOt45VU0dMV1EFnq9dTb3dNY4w8YFH4/MbE4Ma9+jw31EXcSOuiFyB
hMONhXxIVy2TYkLRGCA3w3Z0uFQA7xO7rM/tdIMFhMSjRlIMpBhsku9/Szcx21dPkoJUVGu/8LNh
86zYlbQx3k9G/3gXvX0qrz6O25QrFPERRHYLofmLej0En0Zu0HaUP5b/y/B5m9D3FvWKFoMTVlk7
IFvOpAo/QshVHcTewnqeGBCIXIVqKAWX4iNQ2RmYPLr8VUHl6jTsF0U+IvWeT43jj4u1Yp0iAck6
NNDIyWzw8xFiJHte3LmSTYjOlZev09d3104yEZoRnnoxebAXw5rND1B8M1LWgPJrk2kYzOiub+QK
gw9EHqEg6g74brWzU3Q2qg3zmd/vmvZCEN8r6rTWvYZRVDz2AbdxYJ4MiUM/7q+UrdzpRaLr6ytb
SDnJJWwJsU1STEwLaFEayEw8HXT+VEkyhesAEF59dliuQI8BTMHWSIZZFNlizbpGuIPEFy7Vx+Ih
ODX9yM8c2oo7lzPK/4uWJ/9oNzjRMZwUAP0W0yyyGYlRdEHhClwbJgbykk1nyQHBjWlMQ8s87nYR
u96LI49YLSNWbGza2gVKPxHz/de4VcZFr7W4KGbdi80cVg8OwcgB8UPEgrsoFhY15pG79nxFiRJF
n97yxQpZYppJ7LQenFalswBq65IJJ17ckJQa5d+Tccb86UJdtaRwsG9yz8meqj1mqhJOsQKhJhRA
9vkIUTy+Tyu6lgRV++BYiUGJQmMmaAPqXCnmXRj67o8Bhe5f3kE+WRw6O/YFqiayxjwheXYj9pt8
Es4k8hT8xmkHBxwCwPSshGCc/bimyBWQLJeKEAs3Tbx+wAxrW/oqplC/rFJzHWSPGa1QtTVYEbpM
IFpc5Nn1t4k40XjnOV6Ir4fizLuE5FznvoHltP8NHBHjNBu06Y+8gZMDLqJ88IUAON8/teufYkJU
gqLP/72IRk6PlRBFCy0VXPrCv4hI11j9iApaWG/kVxJq1ibVM52kTfDDRyFXNPGlLxU5JBrGrPS+
3qI+tanrCPfEIa4r1EUoaxdgCoxQ+vlsRbZEic0mYqIIZw49LC0jB6xOkbtDwMrEUe2sOi0ah3Bp
uuppl78cpYmczDkx89tVaIhziUW/MgYGkUitTuohHF4pEoUzQBbp/+NkwZVlupVokr3ylYhxShv6
0cvHv68YaD8ksB60Qs27R/J6hRXCCPUYLcpaLqlSW+sHPOEpPhb/QGT0FVv51AiNtJWYhj4hGnbR
niQQW4Ar9Y3Mf3UKNhldZ/nry/dd6pCc6lfsYMLPBo0OyoHrZXlQ2qVHoQjFSuGCNbbYtNnOqO5f
3CqWlQ3viqAcAEI8yYHmWBzAw42yLwlg+CLETX+HoS3wz1XdcbBsJZPqRe0YlrnqzisyMiuHwA/p
sDopW4+d9EuqqyAA8LYuywsmiLTIeLznkajYl3IPTIazsv4A5NDO4EZtGqdS30X5R7QcKAL7LWIR
vZRXjFZQ5bnr9ywcJxhemQJHjaVa5PMCqQ4Kjd5y2lwcUcqZMAKNucFzzgYOHoKHbAZZVM8OYPHF
NruYyakancnal5Fb2/nXKwegm/PdaTfqHL/R6i8/raxeImvJwMY8Nv1Op8Fg6Qqtca5AR6GRaWe+
ziLvJhshGNmdbY8CgJysUXpes8z/IXOQrlX5VujpoPhFmCHwTlUYMz4CRYRlQWI2VfhizjMk/o+/
8DB8E7iaDe8FTfvbEOBP3xpyiUYfVKQ7P+6bHsQaHtZkF+WsspMB8srgy5Ml0e1R4xC/C9MiFW76
RYSorUiKIVpKQP+/vKah49FZ4ncFjqrPDcG4UUzoh3LUvXcoDPKfXqMp5FbYERbdev6nbjiYUtKx
tzn2wrD5kmhliTYBQ7Qo1qyqyM7TGNiSr4P+JFZc3m7i3MBRflvkOGOh7FBr9oxbmzdAQff4IiYC
X3m40fqw6WusjGH1kXk1oZyeQL/DnPq7H5wFdQhQYP97pc3HnEn+Ihh2kfdL2o0Js/VRAHGtpgfH
WuaKIMe36wByXARDiMNWx7gJYgcB0fdNUTlYfO1vXPkdfeL5UaE23dBXd/alyh3AeTfZskE29PLZ
UN4PJSe9T1QEY7JilBsAIKci9aW2q2aGXV4skLmHsVBJwofyuzEIF1rMaT02qKviATUgmY73QgSb
P5ud5h4yg8l/Q/ipEEjqxS7K77siCFSVtynb87++2wHrwA0O2NLUZXfl4D1xeYd1ph6LaC5H79c5
m5GjpnGDVdW0p6IWKm3Fj5SoEVpQRsVmc1VETWsIJJWnb0aIwUmqf91N1EycoTTUOPrDP3b5vTbR
qODVa0YaFlLpoecllNYe2exYYtRxHNAOT9kfauUEFM/wgAPCWn2ZoCMlrtNLTXaw6+TIWoyn6I+n
j2AkJWSikgvFxPFMeaDm2rUlCvNtE4ABcwRVvsJdv6+CA0ey3qy+M29muUZe5aDUqBhv4oMWFs9Y
i+qKCsqThToYVF58u1Zq/9BhwPJE3TaWAnxYoTvcf+UhiCc3HaoVSEXoy514reasM72fZ4pcNHzT
rHe86DFbQ28vIL1R/ZbPIbM522CHkJCUi8822vEcFpTY25Ob8BwMsdQCuBVUu7Y/zK8hb7DSjHUu
YP6e3jrXxtH3e03Na4pjJqtoCbN40H69nRxmkI6b04x2PjRFHSE4lnsMTpyuAWg2uDXSdPKI8X73
pRN2CA4ccVp3fBEWiCG2E/6pvYgEkIwyg35SirEIWvjiPe9knsJ2oSMC2HsBS8c5GUP/xzLq6nx7
JtSBBOwh1FXHqIrPT3ncW64ItpHGeL1qUNy22TMSttgkEsFsLObL0Vx+1uv8itqirq+ozTrmlQSL
jBH0fGghVqQTUBEOfJRAt00GHadw1uTPPRaSoz6IQO2bUt4gWCWgGDZr6FRetVIU8ZlwFboU/JbN
EEaDnzsml8ulU1ahWL5oF5r+xgycYEA/dpUjiFnLx1TcU8h6PZA1aLYwRcEO6ppjs7xs83UyK7Me
99JfxJ05L2X+Obtsy8NmD8MleaDKKvkqyyTeq4nm+mdl3vYq6JhFcuCcJmPiScDRECAlPcCVNAzy
TJv1UVtsjjW+FTpnF57yFd8gf4gHT7l1n7QMLlk4y45/Go9yT4U8L1F7ulakHSrVTXg1Agii8Chb
2R/p1BT4c6r91ZHufbsgnJ4pDpcdFiDti19ZhWeenMQbCzFF2FaAATVPMi0DGh7PKjgnHtFYEzyp
omq+qV2NO/ItIGcPU45ihXhevIp9djk3XgM13T4pADMMI9gLTM+V5wJjOVAN1NbD0MCRkZTkfAk8
Bo5P8/cvLcQCe9yXUPR6HEIehGCBTnCEXUkKOxhI3cS9RhZpaXb4kTOKHhdZ1ZMV6Xvnr0fW8E2H
jNFcDTAweBByQOwJT6pwblAY+SZiluHYdV8RiEXC9hrSlM917+weRK6nXvVEZ0hKdwdjHvlpmS1L
IIp3sopl7Pt1XgEoBqDEiz0Ad+wr8GTzKh2E3jsgsDVUSuIsWiW2iXGze0DZd8KVpLGbIdmj+qKD
02g6TmjmakbcdCPxw6ozWsw+5/uqJX4WSZ8Vex95xJdc/TsVl03QArvTNvCfqgHtu9wlTKNlj/UD
6V9uoJtMxV+8Df3kYjw/tBuIAf5hcIHQd/QGpeN0kbPT0zTClHut9bw0IENPrrpfVAtW9cFeL07+
EdDeWLWraqjNgCGAniXMZrP7WnhpMc5A5STu96IT1xbfLV27veV60gmFFFe+rUeQX8ACRwkezGiP
ciEh5BYW0ub7JczLsOA25MRlDENCjDVGG9YJD/eUZTx374XriWCIKa+/r0U3WZZH6lBm2lVyApOR
W6jPiXXTx4O+H/6c4HHo0B0br0eIPvZfoZ6OzEV7YsqxW9+c/1brSWqfB6CuCbZrkPOkFyv6APlv
d2y4R6nzKYDZyyFhxP0T3xnBQLoqpdJeo+kbolCUa6cmoRmiuvP/wElN9KL+ujF+exB1H8/iqThG
lsjOERBTUpswb4KQp4Pfcll6JhBhAKHRkI7/U2InbocOwIydI1Vav320iYEqJI9ppPqdNJJ5cGnR
TrQb/NlKaDjygHAWBRWRImn6D1FZ1uDDNkPuc/BJcIhLVwliJi5bicX+uyD/0whN7jvKZW53ZJxH
+D3ZRVlclkNheDTSxkkrT+LT503i6x3JwnwEGuUKqbDQoAA/Plb3MUjqhnLUjoJrnQxfdzZqfOUu
SVy7g+5lbuHTsk/iW3JBoLOz6O/Lp1Acm/2joNQXKtjsNsvWtdqjrY1UfgWX9eLGKBKDJ4H60R5e
BL+J/eBONxkm3I4mCbV2zAeOp8fxlo/SI14qMI7mrOnvO1I1ARyR4jRfBWDsTXYHIj5O9U7TUUVO
nwLo90l4S7UBq9eQZ7u+Kg3Bw1k0kvMmdWGnmO/ZT+fN2DuSrW3h3ehwDUAGp7ov49TtEWZtfouS
hETE9++OWL819fpPTLKEKl5Z0adsd7Dd1FnLR+PJTQLx4RXFkRWB/W9l21TvgUdoIIkk+jN9PYeV
JuEZDVsddN+J9FID1RWggVpV6wEUT2JFPcNqJn/35s4umb0ZMmN5MHnDvN6hnWn7W3rkGyUj5jzm
JW0tuwHewafkKd1GmI3nUpVA9MSI8v6JYVB3fUsS4uUCSRhkOiH05qdcUeBlboCRoszEpjlTAcqo
9Bo3SKRCJcQFTF8Dzdbjg1dx+CVG5BEkm5pHVgXZD/uVsiUhlhj0+/ZdJowDiajJGd9SSLTkZXxG
TL/BiS2G98l3n2OqyAS9O45rA7pyvOzhQLzNYOXkS2hH4lWZk0lBqEc5ggdIL1trdLOrqnCTbrdF
VT/60TjVSy4+lhKwVHmVHNfIC3bkO83Nrs6FjJZBo/SXtcwVEUKtVyl17W6eBLEb+qhBXakbqLwI
x5L3DK+EgVHvnVL6iqBIQnUsAvn2a80BabjOD04QD1nFlas8SCMGq6JquNxzOz/F18W3RvUH462X
S3GHVUe31PYgcSf3qoK9g5t4AUuZU98uFZ7Y1xcrQy71yq8TZBp2dJ95EohSyoq2XKHCJbDXdL2Z
pqWL7Bn626q59oXq0D0sr4vLhdCv7cL5xfNQICV8T5k0gIN5cT8rOCRyvzlnPGULmMzeeUdgeG6F
b1nFVes9bVibj3BpAjfKB2LK+hU3LjlJUgBv7NRbu++r9r/2g6QDN6i0PnJh9wGX1WT2I1mQIv1E
3IRz2mco3jfLWhJdNBmXgZgMcJCBojN9bsTuR30pKybBhViHCaEwp5LnI38hHAktoi22KsZxib2K
0Pkqb5NXm38B/vF2QzAaJv1u43Opwh6Ydo6g/9B2NyW4KzyIUcQaPvYqF7tisZdMXMee0JUDC4hK
Xlwh3rM7luzqq8Ft64xuy7DIbEq3L8OT6K1KXwcBGmxJEm13i0aj3+LJf/wF9AFqML4HRHtYRQn3
fBZtm3AOQuP9Zj8zHyBGbtPak5DpY3rDW+yE4FpqxJyfzypA1dNh5kEpWhR8/K/n++Xi9NNB04c6
0m6Lu6ieQKjmQ3flsRFFriehvlx9u7WnUoS5C0fnFL+h5S3AdtW8Te2lEjJe8QLqnTwN+YlZ3wwj
h+OXwFAxootTljzTmg0FFnR+//fuFMDNWBUpyAw9bIFhsbr3HCECfNodggk+VpT/DEsmsF/lKKkE
ottdjkxbwaG9yqmwc+B5DI25EP3d3Zprz8293amdrgZ7COYL+6ZH3KQmiPCWsaTWySzgFWdO7Fwk
7ZRPMtj1ag50x9lHdlSgKttxrg9KKtZ7u2jgo7P9zpT/igzEcGDTGDa8qga0SwH15XHjVhxk4ztX
+nGvdrGvtU5TQq9EDlQE3F+0P6EPXe5C2DE5ULLfpHJ7F/E+6C9f5LI7RrtXqmJuA4rftyPCHzRa
3BlnJfmUytehyNpQiemiAelcXKOxIxCgWu/IHSROTuaX8hA74e2yVfTjzPzzP0sH7YyL320mFICn
SFZz1iUFtBgCL48bRVv69+JZqK6Z9LMwwQCduTq3AAK1GCy0mnF7G24aXNoCRw5iDjReCtZfLYxr
gP9wcgEq62Yx6fBdcKegtpJQSEPuzThj1N8L5hh/bjkKuwfHkt63Fz8iVDN3Vet0voCjWT5NcftT
w1Cs7zDietEnJS9gOiedBZRLJNbosJ7wWPJo5kjPKkdo+iB3H4WMyZZqoCY8vB4KsfUHyZ9+vjq2
/W/qvus5v8dHM+Sp4pI/aB1kC/vvQ8JnyvTlNTQMyiewG9xGEQMNGhW5hx99ZNyGSqtN82hdHZhl
gZCwAvS58pc3noj7uGmTCj0tRKv5PK0wWnX8mjcZr9A2E6Sj4DrVVhi9RzKCuoJtBas+vTS+rXfc
3jid+cE402j37ATVDgBqcNGxGUSb5EMgjxMUeFAMbFVms5Us8qarydkAuQyVRv7pVORzrT5yY0OP
2RZBu0wYqYwkfm/kdegKNxMGv5hzBgUQkGfLXfxvwdzL9MMLXDAddb2Hw6hAmojhH+aYhIf25Ai3
a/42/5102WvyWJVfJr2iu4m8riP91DAg9FIoLanmES3zK8VdL9r4Uqxn8KlXWKrrkLQRvevHKkJq
iILqOMzN/fSR2/fQRfP5xLVIKK7hHV+iplgjGWqTUvIOUj2pkk/A+1ErY/CF0jtUlIIQ5Ra31Ltl
n3UE6YjstH7Uwb3eV24R/z8fsiyI3W8R8899d2qvM87ungX1iqEhZsYafHoXB4yncdS2oF2U+dyJ
wSCxpn4f+XaVQFKEyUoBIshkwKLfH8WsmEV1VC1ciQKvQwaMOGpG+S9CEy0DAjhhSADn4usHT/+o
hHTFU0ZmZFD5LDrBcRKeYwDL+mjjpFX22BjFrP8Tdmmz+mios6uZMtbOdOnUUUbqzif15FKtd/tV
60/0o+rNDFGcW4XTyTESP6ZQ6zPPKRWnXfeNMvO6X8X/sRxUQkFMxJ5z3Moo/ENGQQs5EWsQ0brp
jAFuhEAKMPNDt0GOBoRd6TZMZ0n+uYBWm+N/LKGqhWcvc4WnCXjBsOpDGSER0TxeirCuV/hoSCPb
Y6H5Nq/MAat1WXIMB62oCvKIapJkbWHGJda2x+QU5tU/43XkfCNVy0BwWuSsDVS+k0Qm2WMfMW3D
AbYOSNPkk1tKuLPy86VekTLTtdc49kMfDxfRqCOLWHrdtEn6Oa8p/f3UB97t+zcghA2uTtZiOqV6
cafX4/eUrXvT49uBYPOaLOH98LpRMd2HV5srH7YH+cHdFq4ZwSG7HN31amWX6vCbwKH1NA43Wjlm
b9Ph3SCDmtSm+R7t4XYoQA/BOu3QLkYbR7u1t7o=
`protect end_protected

