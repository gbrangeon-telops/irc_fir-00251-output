

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HpfjZK6WG7sYhkvMgAngy3z+9zzwD77820wau9oTTb6dakSkVNELcmI1vCDbEcS/48D2LFxL/qT8
BNFOIZ2d3w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VPnG2AZhAX4ivH+F+USmM4TuIe2lYrNUq3Xx5puxPaV5guza4OeVGJP6pYRxsBYzj3S4OGH7b6n8
K0l2LCX8eil1TGx7VbJh+Wd7uUD2r86y3rluWkRdWUlHXjFOxoCZGO3zP09eR4IRsG+JxbSDSiqj
FoMAGfR2zks5CEu7dtk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1IQ6dlJ53C6R12Hzl/XoBaoEA3n6gOO0fxU9jZJvCev68EW7XPnj0pNHAKpShucryAUuc2FQgbE
BwIwQ+0yjh3dOW/yrG6sHXOI8NvAIzuE1LMkRT00JCNCjyt9JL0PrhVhWC3cY50b1mAkSZBVfMWL
G4c5aMtB6wF50NpvOm20Ptquu8OAMlN0E+mHAN8qvWTR+CwIDUV/kvH/83yRaRonCOBULUP7XzwI
uAjFnciSf/F9eC2blbPxLHlWXLQDQaZnUw7NGNc2Ufyh7lsh0GoZzefU/JIhthv3ktn09r568XNe
kk/w7iRo/w4FLMicA3dbzrMyZkiVt8z4I74KAw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
x5ctSMYno/7jD9HwXtHguBvqXjqGDToxuRubQZySJLeTm3iuHlQTdlRRlvw3jNvFx8WWN4nEmWap
sLwuJFUESklgDZc8wPsu9plvibxKvIUprit+FQWsTY564IYlM9a003tG4rrtM7zZ9yfolbWe2MY7
qJFpoVf6XAxMMDrPtP0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JhbANRgOr9SOBKZDRGJGrZPWNKSEG3awknWUR+2QiYueCqJ0p8+Oq42E9W+XtOMQqS7h6dt4lJzf
s2rJvfuxWWYMk0rVRoGeqNzUfiVHbjHTaPdjhGKzIm4Kgu/QJ5ooRwBflBurdW1+74PtPtKpfjcs
79ijwPcRU18IbRTlWf2wzAlLDLkDUewye6if9pFfqGP8EVIxQIb2A7LmwWnM+VpfHc6KRQhcdZbj
LsxdBzKwdjN9Cdt40472gpQEnBtaoqRMW+4LW5rSmhm7vTXSum0cU3Afl+AWq9hUcVWPcrWeYdm+
aNrNDk+A5wRHt64iDTF82GsVuvkYpCi38y+ffQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12144)
`protect data_block
vHZSU9iezXa9XMKS9j3K7uX7qo7GkSCN+2di57rR0tn93ODqiYxh6rufe8Pl5WO6OUCfLrWtjk8C
h57LGi5vnO/yFwK3t0l9ZUCb7rDtDRN/uJmWqFhfa5KcCjvt3X1Azf/5K0dZtu7Ff1TkZOm+DJ4Y
mX74M3a1qcuURxYnzPWYhaVp20PPkiNVNyRyhKpGUjSbFQIOMYJNsoQgU2xQ+HaVWpgEq3Jb2hbX
W4NTJNQBnUkiBKIerdcKVvmPYwOs7gLIMO7r9r5aNhP/ZRY0QM4F/SRuRqx6G+ptgEih9DBfTR9S
hYTYQfVLHvOUSoAhJKBEzQSnbLfgrtihU+E2mhfcpTbMZtRJo+AVsw/LYCOH1iWt3J6AVlZKkbG6
bOw2OCFQtp9kf5/jXbBOURQ7UemaUVxTry5CUf7jcvewu7265KQXpz8On6h2E7K6MAGgjvJb6W77
+GGIXV6PRMe2EnPk+/c9wcBa2icT4kdzT8IYtmiHefqwJT6+/WU+r1bsBFXg883pNxohGcjE/vdV
ljmZK0/hN0/AL28fcNs2iOI9mnvGFWMxqlgpkEcFg8Qzhtahc8ZwVjkceG8WE0fBTYxjP293ER4c
PGmU1qNWTMsYo7yGvoWxHw0NuYs+tmBtK/hQa4DTyWWY/VfbK2NSQKEO9qDPT0Tf7nQ6GHeEqLG0
8xy5UNMSg4UzaCXbkSfiyiMKkPpHMtJXZax21AK2cCtDA/k4BmazLt/GWI8lk6FZFbVmK16cMBGY
R+L88Qx65KnCIT3wc+uZEly9QMTnaNvHQTCjQ2i6rgeTaYPCbgjO21+0d9Fp2KZ3P87N7wyIYGUI
TryANis+1gwf0mCvwfSMTtWrSSwUAwnUGvOLKJrXRLjRPJTtWLKleA7iwWThHrgquu1g/sJ4FUyo
H2uu5rK5OSLBt+OFyzBOfTDHsQPYITlPso8jHzQ3Gyb2crNJ3pAmcfj3rFc9GHLvnitSJsqoGPda
F/LSKbk68dX7Lp2ea0ywDHJTxdCTMJjW1R6W4KANABMvrfJwMU+r/5FQXzk6iafUIw/fPHAZpNJm
38FtYHFLGGYA63dsUVAKcoWvVZdFs7J8r/dM2rJNzTjiDaq7jHC5qi3CKnlUhb724dmaK9m4n0Pi
KywaGcTSYvsWgwS2STmc5BviL0z9tdehbhxxyGO6o9PEK6y9Bw0/U0g8m1g2E1ATHQP04hJybaLN
aYS80rwSomNy1i7WN6vr+K9S+K0tMl/A21CTnfmSLTEA1XIbdK+0qlwgo2E74lMT6BVH68NC5Ycq
GCp88sFAaWVAAlPTwu/SkH1U8xPOAxxtBaP91WCd5EqAvRtYBY/vnKoR60/2JrlWZ8E4GeXnOitE
RnVXD0+LqPIu+//6PZZSnqIwFGMY23w91W31BoUuGeOdx7FSOSVwoT9FVlTAbGfIygD3/pmhQIrh
lnp/KJB4BLu1uVqRV+UvrMim9Zzgp3O2np+hTLrYbYQyfqUgKIabgRiy3tHnP5fkjE8hHy9REZ9y
meCTyA5qoVTNTvag5gxQfaPD0okJZ3AxPvHooXctpU9Qw2geKwJwIFgyXO4KQY852V2CoSpj1X7S
wvBQ0DYCVSCLAFDDHHeuFa8NwfJCkZc78eATsA3tXQEJ/V+6lchOrDUavP8IJVEGXrolwiL0ck7t
5XY7irPT7tGxvxRqdq9ELCrk+HBiju6QrRn4etnbPTAdCcZ3nLgkMF6ViFNp3GAciHFfV0JwWfBJ
Ki7Py/mIZIEVSfsIdBTExJjT8OFbqC31zCi60wOP77RZn6rQGh01QsE61FC4cxQ4sCI0NkNlwnKS
5kE0EFW12erwQ/7xc7fPC5D4xJYypaD2/miewqEyNQ/x0rS/L+H7/sOCEWXBsEc/abFJXPfOGCw3
f6dB/00iyKPzqYl2hnHTnQQkG8eY5rAB30+SymhSpIQ7Wo1CtXBhL2IrRfnjQKqu827sOMeKj+AF
Jzyl5NPdgonMdk+9bz7Lof/gcY3U+AE8h0+wrYwoEWg0Cy0Ax122yqgdFHbQWogLIZOWoKFrEGDf
959/3NqbRtANHQYIrlVWHqdJ+n2CFW40KGN+QZ6wq9U8d7B7TWsAxL/y1HD8SKrZGG/DIc/Qh+sV
1086efcWoY9M2D8uSGpXkSquqYxBe4K9bfgx14O11wMluRzso0bf6nu4vGvpIfI6N1FZOshmpXlA
QIiaHy2JGe17VukxvjaCoSQHz2t2n4h0O8ssbD60RmszsvtLhWToOMcwQEa1kEvWatzeGlJbDIsR
4MWvpyqEeUJFH8iUWEl4kaGGXqFTYaBLY8+SANnfK8OfJWlwoiakojSgcbjc8Y8kha3Px7xN5xa6
uu6DYLVRgovhDXs8t6M41JIoOuOdvvDa9qdsGSPwJJzR9mXhiNDt433SaYFHM1IWj5YNI0vNiwyn
ZJ7vTWZDxCSoJUQmeUyqDIq77h/AjQ0b60o7/VAoIyD+LguEShMJCXdBLzhQ24T2eWVK6s3ueeDC
2BnF+6j/iVi20VcyZ9HuZJXyfQlCLoyWpBdTPykSto6O6OsUvBa7rn+hzlHUpE7pfmKJBTrgTtqa
Aa3lYCbExvmAxK8DcVica+92evHWc/32u0LmmktCcNxThqPPhWH8dCXu+ayYGcjzGwaFCW/TiTfd
VXLFkY9wORpsvgTHb8gA7VguIXusV3JBKllrGrtnehGiml30Sgp/uWzG7Kg8lww5mk9M21usqQEz
ZyTLVK9XTsNjx/p2Fz4yH2fP5fYcBncZR6FBq+hTV04pfCbstVsdHgqlN2aDJyzqWrSMszC633uR
uXoQyvgzS6j8beNZAOzflPmYx/H72N43aEDLwvdpR5bFpzaguxwJZGD+e5gh28AQg2YwDkxrHWLu
kNQJI54xcWdbp/2KUIHQunT32NhTj4xnALFWMCusc3OWV0VuzT9lC1FY0l2tiq+7ojK0icl1z4aS
mLAJeklzIpsMFgaylg6xdjVthlVMlTq/1o3DmJuVHewsECmevgDcGzQBpg0LIOJwOJrSjcgKSO3f
JDNDKQBfbL4Pwg7OfdduNW8rTmcLgeuv7nrdDyl3kmhhq6StuFgZNOdx55j+OMJumVIp40sNbXy4
5uzl4zj7IQgiBkj6A/P1rPpHjt6H6Blik3zXpsky7rdJ4zOFnknehwBjnV5sjGsrJuRJd3+ZWgVD
WQ5pYMUBgpGo3+pKwuer+wGM1WNh0qGtIhXsDLFgoP/8u2Tzw8SUJces+UFgSdrwzRxC/W3S4KBO
3RofQURmCrUh1rxq5lfE+PqH9bJtJRKsovCTLhoVLHnRdkNdcVUaQx8xm3K/s276N2JTxMolyi9e
VGggBgbyxh8pwjtpXFfMaY3ZyJWu00u8rkMqMkgnsoo4AYXNYh6T8NTw8tF9xSL8hDOZZZ5m6u8E
6oPq7hgXP7szPE5fjgK0BHogWsg/lfL0lmHqMybRCFOEJGjau4UEFmGQY8f0FE5vRCNHrWoWu+9h
1bFM3NXCXHoM+qR7Yb61csdjGKv3Kosz3G9K7m21s6/qSp62wO2cd2PesS/riTS2WHBOhKcr23Q3
YnYm6H6szpWv/EjcVAf8NkiO0jyk/RSaHIIFOUyJDCthxrvtAhTdRBjozd3/J1CQKoB7EkmKdN6e
jhU1YmBhW8iZqeMD+s6ko2ergj2eeu607UOJQRuIR6pU0YnLufP6g4YupU/yCXnxyfn2zQhhhoOU
1z3DnZ08o9VXGysT7WvfK6cFN01EquiJZ3uK+KE/S6C+lp2SjOT65e2e9jjCobqENmwscaIcZCTF
X9Lw+gz8XfZmzgXEVFiUxQm79zMpkNJEuvbG9xthEWFFp1XqKlWtbvqoPBfH2mKEUa02AuxGNGeM
BcLCJjmk/WkWNgIZg4IzSCkBkdscf+iPQ5GDk1fuK1/iwdNIf+wWvR1yJ3fKluZbz73+tfQnsWk2
y6tf3/Gam4ehLqRz27EyzKq8RiywKrOP6tPC/C3lX0BffKVgri6bdnVHlrVT/xN/Uu9n5nHQw0Qt
7ObYoYxCK3VPUbJtZJXbCe+6ubR8c16B5dCru0UW/yTxLT7fse/KlB/8VrrMJ+xKNMMC+LoY/zpI
vO1YQoJIbStKjSCaioWYVF4R/8vjC+buOwRhfOtDicllR9VuORAMwuNMyRpeIewloE8wpj5LxJ6k
fG1ygAgTSDIP10oibmcdWQ3kPk/nb+wr1NoEI9BkCWkyLHVXs+DoDCt/nFzUVES+j6iqzUHA2QnG
Tlkt/Ks+P2LuWsXwE+a/bBl8y13tuL9tLwplloc6NmxYntA6a0PHIHRROBhUU20BkhgsLlY7e/bc
f3txAzf70/S9qzihtBBYrTAlP7Wew65o6ZWflJHWZq2uJBHwiA606W1vKc/jSrBTT9xU/10LoI2P
/cY2Mq12nVXGfM55MDhOc/vD5kQAa+Sqfe4vmTFbcWIhZaM+lXIm9D1u7D+kUdJbm5HkjxhzxYGW
dLhN9E41ZYHSemZO//5XS7ikNGiTfDI6xHF6dvNdMIJCTeT2lD1ri7Pc5aIRLW1V2McYURaKM4xM
32wfRX3Scz8KpBoWwHXBy3suATidGUVkGEYsdZEVihR2mWY+qRbLnviRlvAxU5+ulDFv3wkiPE1+
2dyx/+5vUKFagqBGarNVvAKu8gs5hQjC6urpom1bdgoPxuv2R/CLhTqlvSpFl4ytF+jhkek9qPc5
F8Zq1Hxr/JuLLov/kSQlCwagLqbvwpUwDoHmLciY3RsaRiaP5m92zmt9Aws9i5xBFba33bDj4Kce
kiv6UN5STdWWnrCPHcpghVsHuj0EuZTvPwj1BEz/MYDRJOYop8YgO9wv2MwStf5mz0icXzEStyEz
SOE/4pBGL3gTGmLsL06a5FrzIr5MHHAQSjX0xHkK+8Y7pOfGL8269xNIYrwiPplfiNOrc/AOOY9Z
fmmVJEozeYhd/XQGfzaPxaQzN9mQwvUIhClEC4xCvNO9oTSCoVtQz1bw4FPFgsyB94BI3CMtJJyv
tR/2t2E+N5PzYGgI6b+H4lN26V3TsY4OiVKFYP32A/bqJsVoofYI9rnOQ900NV54L3I7eaHUI0Wm
pMo8UUo1Be3gaUntySQjyEJyIYTlHIjqtP3mGVCZqheocnicnphpqihpvIWuhts4MUaSoFL/C2oT
jErTyx8Wd1VQxUpGidOSGX3adky/tjr1CUzbrobWMjy6cB9jIap27ur5fJCdkBNBl71y8knC40+n
dqsNHWU+uzMRKkEKsWccEbSummyGsxORL7RLXje0zqsuugeHKGhP4cnkuoAlToxhH2nQkQyOjFqV
xUsFH0rTYPhlBTZz+BAfoYlYH6ftKq+oBZgSgQdrdFIWAzNXtAqABCjVYYEuo/Jinv3fENKuDgQy
J1aI/MXOceZsnGnpwE9BhpZDPUFQ8qGRRMZkU/r3UCK3CKY0G2SqnHkMAHxoGplbrvXy3Bsth4sn
RV+dHYeu2d9RxosQ7Y/SqODK2JHEP5+RF2XCprqIzrN9emCdixkkTNwUNjGDprHgPCiX7nfQbhBk
YhzPMDnMjPPMZ8N/H2hPu0QWeCF11Wgfscn7GhWtJTRYOFe6DDCSxmk3jlxKp3KCJl0YcYhgWcG6
fVsaIDxB7tNJadBDl7MZVIHtoURhBD/+cShUBpkLY/HELQdUyCUSdcuPSlhmyLm7ftn5lzt/oPVJ
eBiMizMJ7My8TSuWGgKoxANFj25bxM4w0GJDHVitFSzJkWaXann1utUGORXrbGTHzH+bNMRDKoZx
FqGKqOSgEk9BLNSpzvaY5JiXX+MjhQE26zU43b1wkbyRlajyucMyqMYdRK11PTQz25uhlXv9Twx+
RjgP9Jn5eMqJzwLCHtPE2IBFkZtDUDjpMJ3KpV3AgqJAASa1Gpt5SnSID0XDUCkZGvNOJ0H+r5gr
/mJQOEnu9mWeZOAxQwug1edolw66d/IyAKxHfw3XLV7S9IuVfCTuefO8gYQu+cP1IsVQqTHUFWeY
tVoLphN8g0ELCp9dZ8lBPj3U2CkKnS3s2j0++GzrBEy/xhY5R7Qo7UFchZQjlWGVjp3mDl5ufTfa
+Qv3ZJPTQC4/YxTuIb9uFFD0fAuN+WJW11F+0rzKIa/EgExnmyr4BToED+5zBfj48tF1QUPMlv0b
gOtVHOdx4FTRBTlv8+7VU3LgVfhoI0lKOPHE6I5wyJFBOcP85mzuW5ebYCOrp9PZhwDlJCOWl6Wq
7Gaw5Pim2XOixh1oFTjXSLoxotxV6cha54oVdmYlkCTpAg3fXTRWIFBhziNTrcAj65lXo7CgzB03
OvCXWfcunpfCm5CnXbiWeobOsffUGAhgHGUGRHD5iuFNFotYlVQPXuyyOTW0PPhkKLY8rqhwWM3I
jDCMAO809N3uAyUPxnon6zWqxAM4s12FjExXCzdRS4ouQBzXj1TEt/09NpWNbm8Eh3PuhVfiHCUb
6yVbwQQPtVbC/iJNo1fAGlcNh2pzdB9CZm1nfZ2aeqHwGbBvmhfGnuwmbycL5a0E+eZpdHiQblan
vGmqaQmQtzjL42RaDl9llVRrliqbwEJTKgtm2RLOUD+AYsp6WpxoZ2Pv0FCShISuLtuB41Ws3c3g
Q0TwE8hYCeO8fSOFh505ziM9gNtPQ8sxoV9VZWClvUxoyzC6dIKpzabxCSwVvFUKv2sguh2AYMoL
9LzSvaDvDwuofLQOX6bRPPA7CfHuNmXv3Do8aJ7RleHwY4LSYYeopNQVh3RYabDOCEcN0SFHUsKF
4DYlhDD/DTqI9dmYglYnpr5DTf3n5mufGTw2HgOj741m8i6OdQgH4Q5Ey/0Br46Uf4QZr+x8Tgxg
LAj97v4GoWhBR1XjGEFZfiCxIHV4CdYm7nKWTUHjY0nk1RbkGZRldWsVA17HV9VwnAgyGCjSAJFB
1IYtSKiAXJ9p0RFpUggekNJR+pRdE9jeJMnyiRDXUcXAdSjqD0VYEBCMZJpqoFhAoCFfttZF3JIe
muOIzVhYQMBHFutTGV/Ns/gb+aHK/yuyuedGRcPuQdcRU00ZbC9asduSq8nqOTArnIC078jfJAA7
m1yUztt8DA0t5rd1hwZDU/m3WD88VB84dIFSNJf1JTATP1doNo7uOSRswDWS1Kudr7j4dtd+2uZM
oEChHR3l+XbyFpliT5x3wyM9ISOHge8MC5pkuuXQQIiRXf9QOHQGG35MxABzaBzHDfWFQIjljDMd
wkpdL7s2vgVgRR+la7myzmu2s5QxXmZrdfXRqtIWThiN8Ud6Xfb0JDp+j7a5EN4QbOeSShG6pQQo
Wi02YuCcs0wHN6i56blThjSTkZBkGPDRknIWDJpg9v+uWKXuyk/9ICqKimnk3hqYgWA5K/VlvZP4
xmQKAUMfscQhmisZN3/JhpVv9rbQ6x13R6IcCEBfTvyRyWi7wgbqfWnLQ8C4eaQvrafuYtKdsisx
MxjwKSsJxNuWsVCrhEWQs1k6qNa8Rx7y4CEG8s6l+vUTSgd/WW724wlNZ2z+aj86W5MYQxdxvKdT
8v9Oc4OTDh2/Wi2R/unWN/Ii0TyNYnOzhUYECoLdT/eNUvQQED6KhyZ3kGZB+8822tW5QfORLK0k
G8aA+35ezKsNX0q36hxvEmpHiUDDNeTYc62rNWd7qEVpERcBU2q/qEcAjeSjxJZQ62XhyfIFwCIk
NBk94nWFoGsNEY3UGuweNSXoGfe6X77U/0wCqNhVvgjdi+yGbwUWsRaEj4kRXmMi1w8x0LwvcJAu
cTJylMIxGjoQ5P269CjvRNYQjEGVRAJ45DnrhkMpixk26Tfqnqj39IyjWrGc4bk7kG3zGtxVGFDK
CMUyZaX5x/fKVkxLeyO/qqnXZe1wPYqJi0+CBQv7313CnMcFFrRfVSeu0/OCJT5uZyKZImysNMu+
qKWfCHpeYYPkLA7BijQTywRe6WN7fEo5iu5snq4YmO+vbMdPAqBd38ATC1yhuobcgpoa+MV5aGj0
9+M7Drdme9VSTEP029V4cZZjV4LBdWfCScp+ZItX6ikaRkqPtZ3xyzG5FDPI9ZepPUj2PhQmu4Ep
fN9Ir9aNo15w3xDKy8d1SWFdT3TBc/YEYfqPrga9TKTWiaf8PLN/auuYbjyQ8gLfY5kYMLGY6qqt
/528VsJs58r3k98dnxSQS7oeNDZXr1XQVxi61Yhk9HXHWJ44ocGZZLLpBnXJr4QAzM2CqHMNEwd7
e209PZhHACqfSJsgiWQDehGiXxnWZzZs496PB63i08FPN/T9TzEHG86PIoBTssbpc65umr+jbmtF
+4tIeaz3+UVQTRaIiyVLsHzAKnU6KtnxmQ0Ur2OiAa+WSFldy5PTfX+r4Pt0tL5aqCDV/3JiaTZ6
78lY3HLI6nqcCH9C5HnYlJwhTDBaGjVzYb4t//fFWnbPn441kSdZW745hfbwtrDi4Xqch3JOpcnY
rLUJFhFuZuJAO5I6VQkc+QuBkrakcTGTT1LPocqk8R9o1OFxfzEL3T3IwLJBW9X/5O15QPcW59p/
3leXa0Q+gmJ3z9ubTUyTMYLDvpMHpGKKqRLx3G6HIv3y+1nVEHNoMIzxkWxohNgE+smJSbxwG7TD
gAl1bHzAOpBVIzWqdF4LtBtavCi55a6jhNU3CH/uNzfjuopdkPQgnpxiJ+N/2LB78pTOKok55yVO
r5Pv7k9eLoKnYaO/Bi1OGq6hLTaC4V5IdeZo3X7SbwhqX1RhEXYqu5Yg5cStuB5uqIaeLs0HcRde
Juux691n8gOP1xZd43JKgfmsD75hHzHCyIVykmslwbUs+mWzmdQ2VZWqnDHaS5vaYX9jAUrWv8dJ
f31alzY7+6TcT0qAKuE6IssW1RrXy0bH/FKDZS6tnf5PDhYLWrIFjr5vOD8KzWGA6txYaO/84whQ
R80B/i7D6ZEkSVTkWL70qBooAyjRxV4dlKLAILtdp/GWaZyc94Fkp89ANZNk6Lo1llPAJXzsEG1u
KSy2N8gwgHZiGr9HNppWLZQom9FFcFeVQQpsx+oWYPpqfKSUwnK6f2mk9T5TFkH8iYP6ULchr7A1
Z6zxKEdXr7w7kjX+r3/RV50sKG6ZDjWbYMNPbVJ8u16obJ8+OjschBRCKZWQMYDmJb+LxisQ/h9c
Y/vzpRoHTTAd1gABVHF2ZYXr4XefS4b0NzodYyIqZFy5In2yN6pMHKC/426XjLSUqnTPtmDnLHuM
TBGYpPb8Pvno5+2C0TEa646FOlFfXzHqJxcBiNf8b1V7wWhHY8tLTwwQ43MAM5eKnfS0jfa7HYeF
Jugo1rkUOmlopUr7Rf2ugk3BYAbtO+Ml3/MuCmahM3Dh+Ra3R11luhoKI3ydTLoC5YmyQ3w8s895
+DlgE1TS9JXY3I7W3nFHUtCPSMo6DkdXEFUJHnSa3fgrnKwiUKAtLFY5M09EbTjbDz/uRv0TL8U6
/lbTOi/yO0zof+EqH1hm5EONG7EvLJHanM8wg4JJKGjo1mnSD/a/DrRWP1qGVDCQrumiaqpodAJx
fmUj1TlCHTN5j4WTKgI0XIWqkgMS6uDtxmKvqMiZf67SqOgBNfvQFcF+sbOKuHKJvUwSyPXHbwFv
ELOUOIoy1rFFI/lw2KdAf0qQSE1ks7cl0CtbgqBuxmkeMiLQu/qJRtm9fycquFWhEZnryO0csI5v
kZgyy43eSVZlzd36HsRc8XyPg7+8+aSUzQZYtlPJoU8ackdRWnP0PzfRgt8W4SY1/4qONq/D0RTD
n6CSVrfziMsfpWmaJfXi4aaxAZC088kERw3uDdc6RuHGWafKN0WWQqebRPBVteEXa2u674L+yPFW
Cr0Rvg9xDATjRbqW87WMJY1vki6uJCjqCrD+tU8ugmgIHBfdhsGoI64EyAPXZG9kjnA+H+PqB8yz
vKQWVX7XuXXkSG++PDQ/R2U3veVeSZIww64LMmY8Z+07xjuuSoBDgVdb5inAiYyaKveaZiZdFId8
9gDI0NqO/Wab2RPrNrQ7HuKDFA/moVXMJ3//CfbYnS08/O6upZ4vXL6KhNvuXusGtMnf70F7g4Na
/UIs/PlMC4YrVR3I6TbPP0pdoT27jwRmmn62aDSzvhCDspyFJz9m+17hGbRLiXK5cIbfghimCSS2
4lne8Qy2y/g90JSEWUlW6oKbAzuDvWIw653n2VTBwRE62pMlah3VkctKqPmLBgqqeBlmCFHFkrYm
MeN9oKnu90AZTPBMk+rTqdtlTfsr5pp/5pBKS7Wj2kRxPBG1yTw0AwAN145dn+rsZI0l1xEEPWy6
c3FKMkzi6+LPO1MykbW431Anhs7qBRrASIW4+UFeNoLnk4e4PyZZrcskce/t61MWOyrqV3FN6kxi
RRSn5aNSRUt1lL+DUf1eNkMd/nC4ld37MzcHhFeKPC0Q8ap9x8fXezc4KWTN2vNhvXgHOmT2uN4j
7/F4gBFHQyNLBz7J+YAi9XR/pMFtW7qxy7HCrLi0+xJWmQLyIfSu6ezL5lYaF/TKpw7dJCSBw6Zh
4rOSsFf/OdjbdEbgl54LUbY9HAZFL2Zk9CDS/jmZuLNWmfYdU64isrwdVCJvyl6Y2PcUbLNKvB+F
Gtr6SKD6XnC3PPzNyMnlIvfz74bisE2tDbbiahckwcgs04rXYVu0VNqyJCHn7yGDS5GuKDhQYHw/
Bb7aRQdGTCVQ9gnPuHw+/yM4h2X6g8CW9MYPZBvYeJiwiQB9H2pAVNG75yI2LoPqv0t6H5W2bKQ0
1h6nvs9dNoZDCtPV6L+RV/E0uuHSChThMFnd31mQwmWj4Qb+enacHiwHWebhUApqpAQMdOBYD7Z/
cQb80H1oPtgL9hyE221G2uIEHl3+0PqBgc5Jb6KyqGChdKPe9XQBVHqoWZMXgFsF46BR6hwPR/6V
qt6Jdh3lJiuk+z7Z6p4XXevzyloRL6HOrYcEOUVJC/4W8ENBQYrUcfP2jxxtIPb8A7tTEM5trGxD
tJC1xMRwSJ/qQvdNxHD8GZ4GexvbSUoD6G0G96e0JIVD1j0XcuN8RzFrp4QPmYElmOOZV5YOGwqJ
wsjN9SLywQxRIlUcCNju+ccDPm119v8JA/n4HRvD0P8Ix/1UlkCsX740ozNHebO+Q6MkwLW4cKGy
eTw6d9f9vBZ2JiVzBcKUanirg+DMTYoQ2iDrHc5hCqHli4jlEDvNuXTtUKRaQwkq1A4ppVIaoPSe
8auz7iXkyxZtbokFeCUp6Qo2NHo6rWReDw2LfXS6COZnC9BfpsyT7rxpC7UcP5tAD3wiB83nKtlQ
ybieLEbiyLoI++4s95QQjUti2mm0XsCA+RiBaSN1mUKGjTdtUO+TYGncou1OwRRbnLzXsYwuiJMJ
ZqDCkl7Lc42fe95daVrpl8ja9U8R7v79tLI5PemhwddFYhyx/mhvFDF8t4toqxBkoPiksKafgm6D
Zoikum03lfVFMH9dI8nRkkZeLLf3+hYgYttMNTLOr++DTLWjE47lKIT7kRU4qE2AwiUeuDwKI3T1
yvvoPQLGDecTlpaHTL0OJwkZZmsf36UGf9HlZblsF8C4KkYgNFIo/g5JaDTabmuzquGEUggHigMI
qn+T2YViOv9TLqkNbS00TFZz2j4wo0K/JUWBz/s7HE6QmW2WmxlUPJe99O7IV05+IhrvY9pKmzbL
CecCAkePx8QvL22VQed4dTSbpRH5jDz+9TqRU9vSec0ekZM7iANI9JyJ4739rv4aUUSj/iq9WzOt
9mQ7t9GOydNYHc2LtT9//rt3l9cTDsm59A4lRLldQqEUByNUnrwtB61BjMd1l36VR5PAr2Fl4s/8
MkcTzSw2cVN2u7Jfq482gKWC6bLOj6VIuXhwVNFexYXsPjlIno5neEnJS0GmbGBaqPEBS8jAktPw
O1ruSevmZrOuEjpkgyrcjKQaup7OMG4sf8i1zl69HzcEm//XfhcQfHSQEPeFDv4jQAsdaikP3CAt
2PSQgG/9vlqa1984k3khph9B5MNi6M8lUElHsUrjtLtSg3WA3PFvWcbVn8rzYFYNCMc/NsnAFkxW
j4bR/Xxq5ZuF75VmnqLmQ3dV2o/Zdn9so1yREx7PIwlPcMN3LYnZeEwb0veW+3jRSoUY4J0GIoU1
b0HeWxeVg3IGwyWvwM3IHJfScTDi+oQr62MR334lNDUCLeeeltw/JyUbryIdvtDtvSpNkcBMwInY
py1ztmwBl1ys27fwWJOwrmeeJv10IOBmrNLr01k8itTDfalkU3aALwIvGW/koPQo5KDVDtS70fLw
7HkkTJ8euh0SFmIWSL6wymaz7qNnFOE83VqgAx9ahewtnb76Odsry+eEklMVXkkL+UAsvkdRmLJj
L4XM8CCs/WeMXvf4nUTR6jvb7fHtN0mvryXXmHHUDz1WtoLn31aIlCjUc/lsS6QRMUCarcH8X0WG
kPY50qjvxrJBwDOi1/zgiu5phf9IMexZaWgRls3d+91eIFVYn8CUgnNXD4ERC2+1K9O41mpldFkG
7Rmrn7G4c7AgIO8C5tY0PzFRuVn5ZjWib5nDKEAg3770wna2q09XBWiE+JkDHEExqpj7/lO88igv
xjkZR+u5RZVydTqf/ZOibMOAtvl/Zd9N6ekVGgiUCpzYd8MazVXul6TAKE3VjBax3fGKPycUTCtu
+9xP0wDujcZSXkbskccYwWtFdQE21rnJ+QhXOnw6Jy7qhoogNNK/De/8Dx95+z3Lb+Mq0eEFTT+Y
XlUGR0GhJCewRUnydB37roR0q48rDnsj/UA004HTK41KoGEaNKNUEVliaz6EMh6cMye6HMUurTmy
SJf2Y5ai1kk/XrGCUj1DunO0ZXef2DJWWvd8pcRZmVW4rjuW2RwKpYX7biH3zzl3yTxGbL8cxbxm
jymRQ0RtDWVEjxH0U1yyJJAAivAOIMSSReXFl0C+7vvnlf024gk3ao0+fggc3RoHsAwG8Bl8TvUe
LxZSFa+N8/Pp0bYlujZCeN7LYQMpfiDSHBv78jgzwXC8W76L6Cp/M2pbogGJU2U7Ep0whSZ/yLvM
jMluOK+kU3bm4fD0n7ellqzTFNvIqsTvPunMzdFR1zNt6dqIxlnjYvGZE6clbi9zUdvDGOJ6HmbW
wW/XOsliIepQCWUWT+5mnlScCdyhLGUgtpXpGiuwfuTT2SF3Tcel/WfJcyoY9ncoY10yUHxJ0HLe
iYSR009mkKwWAW7J75QMSJJopd0Y2gkHcxJKALr+sqbYgWl2OIVdnJLgJXymL59oHXAaaOUYZYY6
G3Va8GQE1SejJm4xpRAgabXBSmbAFxGYnEVtoqEW/2DLrsP3ahGFbLQI3+SwckeqPY1iQDdC7mwc
dhHLiW+dDRH5d1wDso+ZKVKZQTYjwiL2CZ5YitbRGj1pH1AP7UkS/l/nhMxSVAtADeGa2xKCfaU0
n/DHsfu9nS0r4AaQVw/HJsNFnjwgOko08NT/uc00yAkwmO5drdpieKhvYyWLuRal/pYSNvm9livk
4G5tB9kueBBI9MSP0qrLwaeTuxWHDAgrfbBP+gw04Z2+S82YM+bwKKbZ8LZozR17LIbhbd53Pv0K
/giP6Pfh7JfuE3OeMTcGXKOstqjIfT11Ts1ZGkXHbqD9yY9Tt1t7ohiNW9Lhw93jkbx73Zi5yQG9
6bKgzGj5WbDiAB9whEZ24ossWT/xf3kq8G2UjhazaXdjyP16XYIQQgLzF4MLYVaHhhh6LqYIq9xS
Gv2Ok0gtPek1TPKUp7IXoGffk6TR+7pIKgBi98LW74O5IRyRThyxO9lRMbnvZY7eNg4TrRZH31f+
65ZJAkMJ7qUDr6+AspwMcDUvAbmbS/IJGY3hS9F2U5flc+uepHfnhfL6qekK3LVWhkSfIgK1s5Kt
B2LwhTXlVumqtSA8ceK3nSFdHE1t6ryhW0WDgYGgD0FjuZRz9KnOdZpmBDKsnScnmpKDqqK42L9x
rEMZ43IBS2TEeKy0qeN61IGe7EtyGzLXEnFHV8kx2m4KkVueA6J2bq4zFpJAMf31hvFzCByMGvze
0Y1KTpdA87hKbU4ic+ELQnF/kXOdab7hQOgJ42tbSkxtrpAbVvHVe7Ue6AONn5wRlXQ7NrIRPQBL
iF+xdb533SS2EzaPtFqCDlLPQnBO6sVbJ4GXpzQaTn+w7qVYLilkJvqv/6Sy3oNmDk1m4NSIWcn0
ZI77dmo4KuYJGk/BfaryxTsU5k/wLmkrQkZ7rgT6M3PVgOkEO5TX0070wqvfSnEs2gfOCR7ZECYK
4Oy/WwRfkVpHH5+gCKrHxBH8ysErGA7ZF54xSg/b4X2ImU153B105t6mClPPjGhATn4fbsve9lh+
/TAbL0SD7ffVZg7MBI0Hx+slL46/7uMosAUv2+HRyrhuv53Uq4lDb8ZNXfdzJESzoPIAPWW8mx0w
1vkbm26WKT/Jerwnl+TYN6Gshlrfva60n/+KXCA6qK/V0GJbmn36uls/TUZdjX1f7temYSAsxUoI
O+W9Mx7jg4bYpPaSAFnZHjHELXPJ3cM3fmF5lJ7Cn0E37ZoRKNM+2yVETZCwyIRO7XGQML0fxYSR
9Ki+AEdzWxXvZEHfkgxt4ONSaZwy6ZaIH7wG/154m22Yl7XhizhbZq0iCgTvJ/ssb9MnxZiYHwrG
in1Lq95QbM+iptJUzVDy5VUalybPTHeM6595zEnRaMyXl4NUkT6lBCW9O7I1WVKIvADPp+j/lagj
tXqNB0ffvUW9kKvrnY2HAR10eQ7egLhYWBGBbQc6WrlDaMe0MZrKeO45oT9Nz+XxHn0je2c8mL0R
zwnVJv4ZKaYdB8kdjp1Zub/jVhKGYmg5Ph8AJvRjEpCYkIn3L4UDzMW6gXUJctRX+7XeRxI+93PI
nOtW1MttyPXKwmVyeRIfyTDlXDWWu81vnEhAz+bcu5FTYPdMYEKUKeqe3MuGlHlVtscYEKiu8NFk
TTBkim9tZJwXNNwpCnjXLUV2EsrTSJ/Pcqflh2uPut4M1xJzjf/8+68fDWunY50dpJHh576Z5I0r
PCGvbPXaTgj9NeB9jnwWFo92bKqJYFcFFNApn3TcAt0Z8bySyOdSxp3O4GeKAtn9/Sn/1AwxjMTf
RKKlWJaXIwoBloZhQ6w9cLNgNpJCKqW77e9zjbCVjfW88q6j8WCeCARLUcA0nJ2IR4qs6kyYSotA
sbUFPU/N4+mRQfLnDo0ZklFN/Z6yX6VFNDTfe30r5JROkN/jgMfCxE7Ea3mCtRDrizbGxeBMDAjE
HWM9ZViBpa9mt/5BGAKZ96LpCLEoFZN43J+9A35BrKlxfsldn7eSdOFxrRAbxJ7UIIyuHJ093Jza
e2mJ4ZsRtuD+tr3I6O8VdxkRzgAd81cMlxJA0ecgefShuKspLNSjwxINcFRkLinECckDoQ7BCxs+
qi7CfPuK6ZmcX+QUPjInI2c7MmV0HONopS85VvcgPkZxwPHcRoN+9x2qIfnWid+Yxi3M/wJ26W4I
bzztFT6VIg6FbGouBuCzF/1Rray6/NE3U/6ODeCKBrSLc6GAxSdDYTpuz9+whnmlJXKeHX3jMGZJ
XoRb2VPRb38o07vdcyxxZA2RsyAaC7ZLzF6wlqoe7dG/znEOTSeeVvzBIi4s3BKqJzG0IGaZg66r
sn/JY2mFRZ05mjHHbbvLeb7o1mnximxFNikm3+1XCrEYsCmqBWup/ZhuzPEaKofuyk/HOzMcm2RM
iU9poWKwAZNZmp75vjR0BRna89m+d+s+9z4WwYj+t4Nfm7ii/X5yEZsKBQhEedjSOOlOgivJa96l
wvhYtmYtCYEFwDzlbaNsbSnMifpo9aGDD+HDnU96dcfJB1oulMhyiTbViehRLOBhwSx4rWn73EMB
dfgFGqsAHCFusf5D9bpFpcLnzj642t0X5rFfitr3y/RQuD/BJOVqPs7tBYSD/pqPujqU9ML1dzHQ
vW4ZzxKUcdL3wPpOckemk8EyD9iFUHayHB3NlLFP35MqJpuTn98Qasn5wg2HT3sIcPqZ8H6fajtN
6osfcRJ3CeD7sjpIy8Q9hss+25jCvChmTETTSu11BOxqsRte9RNcLFkZNHnxQwJcuqNskopUi3gw
Dzv/KEokDSEo0fBjGqnTXRST+XBfGt8NihFsoTSpA5JmCEJ4bQsX78CF/wLxVZYEq/hDR1jVxI/K
knh6DAEX6IyB6kfgGw5ySbX8qPDTQgCtPNBetBY7oYNGX/OKeEKm8k7ehy8PfZKIZs+HZ0017cgQ
oykO
`protect end_protected

