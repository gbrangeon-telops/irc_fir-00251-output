

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mwxNacl66MFUVIMc1Encct2aHZOcb2pREujQa4vWHOpoY4Ryx1q0qOlrkehqJnJB6VdIGpRZ75ar
fafQO/Fcyg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WTY81lfpic8wiNg2xUTFY/9pIQI3CKsiY3j1Z19a6adif1iCy2STS25TLTe/dZhZiWj1W1FKdbVN
mTJAkstRD1IiixRw4XPUhHS0kg8DebELiBmCxBLwbMicqplV5b6X9QbZ+d65v5AnURtcySKvK9fO
g9n8up28DiiTZN5JTCs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wSJmxWNG9Vaz0hV3ma6xxbW6Q/tt4VebLF5ALUnEWrb0oMwD9MOvKTVg9bgiL2D83XqOs88TpeXX
Ifg7m/wa0qnVENMQDpzrbdsY0X541kchr6nHO22IjxAZU0y34IzPOD4wlt/LkBIeRhuE2oOUmiUB
mj42HGuDYM+OLJ75MJFObfMegkawW+dQ5MXJZAvaZb3Gdq+Nc//x1D0rUYdDzCYkIE6Z7scW8Wik
/MJTbyzmOPOK9ZoDJMjaYzyR5QyLAdSzLEdKbGH7TxDHRl54Q3XCa50pfJuN0PstSuaixGzvKQtH
Tl8qJKpy3o7KeFGSzvILj3NDt+zm7na/fYnOyg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TWs0qYIcIilONYk/cz99Kwd1RIRPFnNZwYyu+ici+iMJ2JCkq8jieFKJjspKJpdZ8Nc8B4CnG4qj
aN9KKPyGY83yGWxxRkXLLk1fDABMFcSV/QWTMe6VkTZV7rSzb+eWC79VK61VEPbjbvhhwl9UlHat
EKGcZET/5AsZpsdS5rY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J9Mi5TzDBer7RNgnQmNNaMr/oObsCpVjypskaWXDXbsUL9Tz8WTWA1k8rjWfCv9Dmq2LFoNWohyz
5PixLjvzdMk+0EAtGJRSdyjvZnuW2bmu6ekaURxk6HvWMfHmukxtVO9c/su/PcWlhTBaWmQfDEOk
MXt2eXdYnsY9DHX2xUQnYdQty3UwLIiL21L3I3SO1yyv2PefA4p4KfovFGDUvBPco1deVqNYRLx4
GphEA4vKS+OANoIaExoVeJSpvDGH50O+wbHahIOE11SE2zucQ8cWichU4yUJXYALRvrOZArC8ClG
ouWj0ts+fBWmUc+Q65XK9XqQ174/nPdN3w6Fsg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38784)
`protect data_block
0Zzz/1yHECrNqJ56Bj5O4qtsAfVKItR7dORDhx1AFPx9ECa26+PuXxlugkeJuScEYQXf0qrVPxri
9sMOK4NAW8q4q+GDVicNctFVFX+YkhxQR5ZOwG3IsB8KjXAWsuA8NsG5m8OVLryVnnFaBeWnGWnh
MycjB6kaB3m7xQZs5/zG875ztyjB/ZGOg7IxUxwE2c+pqKzaa0sqNU148zevm6CbDO9tl2hZjfi9
67GuZBX88Agv6MWUEcVT16lDqm7fNiJJfKWSJMY38AABvlmnn6pwJDw8bZNMPOr+o925b+r2HIl+
T6cxR1gtQ9kCg6Tt7ewr1Sbqb783Yv2ZFGzGMpLi59ikg9o4sIkkH7dEyKhyJ2N804m7xsd6vRu2
DuvFkmfvGySESKEMGri0+DV8vT0uG44KQSQ9C6lK0+qIrBHuZB5yqD1JR3W3ZIudksWwTW74nlJZ
2eXiniOYsjv/s9rjcCUDk/SwclKGplCgSQ0S7Eu5fylM8Y8xMrX6SCQ9DzvKDN9GtCjTKkas1Nr7
SH24VuWSMxj7WgDNE2KbKuDau1gwG9ukeV/pS98UvJSiuiIofU7j3+dv41313zopyP7bhnFoAaeC
FLEtld1HuoRh3YWxFxK0aMfSxfE4ec4gbQTUq13pQ161RPyzoSKzy6p1ysb2qyLXpGOqeSUrwsSn
h/Q1EqLGWoXpviVDIpE/T8BDgS54LbyWgYxxd5ScZTaKkssQkgnO05U3DL4ypYC1mqoYu95HqIVd
GMj9HMJMDbF+j0Wz8sP1SkDYiBo/KdTit0SvTnP8eiYzHTWaD+rC4jADzI/aqv1Jvy+mSbAdDn4B
hd8u29wIMOPPRZ7KHcy9hy9MCjaEQ/JaYll0UtCLMvadlfj0sJ+0AeekJexbaH/NDYxbzRuO1n5t
I728Ygo685NIzeujDvUU+NLpiSrqjrvKZ1Qy8wTaz8XoL7iLWWDSDHUnb3NyzBGju9RdooJA28en
oUyP6EXjazKXp8z0brR/dNefs9aBXDGNGq8+AwQsBpc2//UCp01Oaca8dohlcRh/gaxs1KQEYjEO
VS39Q2V5PT/YUrqwAg6RtYvAgFHTBP1RDaWGcoQing5X81Rqv0Zgx06BWZJnH6yqXZcuO/beux5r
j4DO4aJlBPdeLCB0I+2IcuXLnD0VOOj3M9B7+CAYchrDBD7HZeeYcHfYddYvMQmpXQD1kGRj28I/
gCnCjLKHzw1vi7ZrWCtomsKXPlwI6PVIUCL5Dyfoci4pDHOldh3srio0pT1QdC3zU2cBC/8qVejn
SjYpubISwXjAu+ZUVfcWOyaeqjzzzlmMSaR1w2panK01heWO1DvPAgMx7B0kF4qhNpZBdX1LJxuM
61MNVKCSUWi/bmBjzQU/84M2fp8kP+81nU5CI11mBimbQOPiFltGFuA+mw6zE0rtMCj1ULvMXPjL
V8LYkPrNQjVcaFFqazXHPNA/9zJ0EhO6yCbamLSnn05u6I6kePZfjxvWr3/AP0+37GpUJIbZ8r+z
8p1xITaoTf+cR4hEEd1ZE31nLTkdX6NszLzRIdlFMk3UpaxYPRi0oBFdLGO7UgyURkGBK1Bhg6Ne
RDlHV/Mqo6nvUfXYojxMIj2ABseSeWvweVdvzr77J1vDJydgzMUmpK9qyC86vIp5b4TAH/kLOZ4V
zmQwpPFG6JYeYSa9hKT3Nr8Rc2rVjv28qZ3GXy8TbLpI4fz6j2EhB8GKEV334X6xU1cedlLurD98
vlaGDHWOYPHmM9LWj3oJmGjXeo+wpw+xUNgfvbjR/BjwPOQToEcZHinz89E3MyKiLoyNchFkRt6u
5K5BQgB0ibQTkK/PDRGi+vFYulYtP0/T34P+TGwyJ9oVwWnApfDVCG1zZSuUN658HUUxqNsl5Jbc
24t9ndWjUpj/On3/o9LJ1BE39wFQCYjC3OLyNb0cYqL1uCqwufcdW3g+oSjcFyB27XEvALwpUlI9
PKbunwYup/THakMewiejJgYUqgF/oty3PJdZdVh/pXCdBf5o4WqJWqMZNA/lb8GZFSr4yds3lEqJ
hCV8u70vECsCVVKRqCxloZzyfQ7AzRcg8Uxu/o+jlqoDjnvj0L+tKbq6sxs4hYCkBeTt9CI9F6Lt
M4/q0dxPAkqQmIaLGHek3UIPTSZmM10hut+8uIHgouirzO08qq2zm8DERQO5Jkax272hLdPv7cab
8mXtlqGIiB2Vh7vMwzw7KXBsZYk55CuDAcvyqlnpGzLdmDLC0VUYWHVMBVOSIwGc3gvihXnQNi9H
PAjt4jXaki7RT6k0TEyVI8ZDYOxpykFBTt/Ga2uV761TJGEuUV8TO2+dIGJzYz8kkNEadGLANc3Z
TYESxuO/IOuMmnXJNrdS5gkhxGhp7Fr5j3XjhHshZHdBDIeiOeS2xzZTJHigoi+DJV+bqYnLgzrZ
ldmwbd16OHFCbPpomNvo2zBNuAirYE9+E8gfxZszz96AdHRfi1QLuXN2aPo+bkfsrK+PxDS7U5QF
FbpxCL1tPAHyRRtfSt4QiyaYT889VPDwwMBbBd9cmBxoGoYCkcYjpcTWBloLvNht3ZcgkE2BUizs
IPsiofEZsvX0PFLnPPLpXhTOi1iDqRCncU11Eec0z9Nacp/UdD6fZvMDemWRfrBEre3r0OSlX47t
6erxCTxJbcPNBbvVLMDsn9iZxfLHkZqT6inzu5IQ0tkc3chhj66ve6ewF9JELWq+FCLYJqD/OaI7
BdIYzKlgYBN/ekBaqAYNN5/PPZn3vVqnM/1Pkh27QWdvKcvfcdU6OSfkolsjvV/tn9AOUGzpOy2A
MFEoO7fuwybeetUBZWQ0CFqV0GlM9xa79CtCB1L8PXAmjw5Jl9qB9TIhrHRDaikzOLV9t/8XFRHK
JPlg3f/4jrE5I4uRRtgfnd9xND2zlrFb4c/wiy/g2U3HVv70oC8qGg/SRP+GMS5zsI8eU7+3dWxi
1eh/LaZKmNOQWZyoP8wM0ESqrNVQ/SlyHaX+J7xP+6seURb4diGESlRNN018Lm9lPaU95Xigbybz
V3W8p9EqDC7C4QV6Rg2TJmmB7cx0x7z7rGa3G5B55Bazm7KBxHk/oBvQ5vFEOFwleKj653x3ObrE
jrCQuzpf8huJrsgethnh5uVGjLGFyV8NXzjczD0XkZ7G/LvFyOOz9O3y3RbL/fkSNsetSSM1QDOO
47gLGgiA9Y2FrNWNULp9MZPKG7elsflh2m4IGt6KCGPWwD5R9Mi7iOaFx7Shy8Zp2sByYy3kCKvh
sLtC7k63EOJlWVMLVPa4t35CsZy/KAqYKlKbDCIh5p8S1NnnJElNV//qaYEC+6J9FvF4ThhZ159m
zB3p8iIcd7oHfhCnWcE+kzyYOefdJOSK3eYXCU6sC0tHimWQ3VFdogNa1aLwPeGWWuynMwYc5dqH
jB3cnkBgN+qLQU4WxXYl8Gx0cyb7g7CT/ZhnJLx7KShbWlysy5HbSUw4aMMkzC3ubd/pzpvVN8VB
EdD7kP7/RQwWPe7jT3GyKM+JmP2gRmrvL0qoNZc4XWuj+wqbdauzC12XlLXpq0rq2/MPzPc8NBLb
ArtLVj0PqDwvmYoBuSeqGPTCZ96DReJ5292xwXKfViByHAT+58tVMP2CInNA3gr9GuTDvgZtEKZ/
7oHJ2wlk13ZYgDDBOQy21nKW2eC50aCXnX9IX3m5yd37ANTsMDKc0qjpL5L6cP1wpjmxV5K3DsAo
fmqBe9mka5OprRShL4RhFjFSw/GgwI+7ET+hSiAWW3n96oRd8i1SECOWIcf0P5Bw45hzb4Ro9PeU
XC/li+54nqjVwCbeGOrGkts5S6IB1c8DM+aq1O58lc38AiWuxiKsm43KrB0M8/DKVXjJI7VTP6/d
bvO+wvOaA3lhupICx63Fs7jfdVGhdzYkkHUk9Kn4Q5mbD+xLud7Z7yVBaqrA3nuiRJqlnYhyuf7O
/+Pgn6FSJ3JQY7E2KuCE52Rx4Uq9aRPBQ2hhcDw00Ot4/AtqiTmQxJUVTTEBclXBKr8ou+JXHgnS
jY0FkLfco5k1bc3tqB8tvPMnxt6/NYFLktjkaGGAEGJA7mIYx6bVA+bX3vlmremE08Eca0oCZW5E
nzPLlmv4rMP0G7rP6h9351J/QcMEhuCaI7pJsJqSkBmvnMBZVncSPoIMzn3vzS5IQYEp5tgFj/mZ
H//EVRsRkzXWR7IA5mGwlp1dLn9wSphs1rpSTWTBepv7VDmHlkvbUETX/vZLtMeKjZJGa61O802i
ZMnXc3cb3iTacp0PBhb2Bky4CdTpXXYe6zACCWT65xZyLNo536YM8qKKr3meXU3oskQEFUI4ubld
8MnszO+4xtALbzn8isoAyvQOVVvKsumaqCzuTKQBUsj1pAE8Jwj+US0WCKt1bDV5Or7cr0h+CWzd
bNBoYEIoYIC9cgk5MNhnI7o+DCU4guc4hLVoPFV5AW9Wp4nvYnfo2P9+VO5snMzuE8ODU07R5pat
qLkx9LPdMOwaKMPNyJLaxm/GrVd9WT3tYHUX+m5pYoIhQk6wY3R5C5KAUbcAyS97zeoHe9z8y7ml
uT4BAQXKigRAj73R4FGEUPPgfLduIL4Kmud5MrCdyWBu3H3iyZg9LwUx6El/y1+UXzw5d+7LbyH6
0bmcj9UrjlshZ0tCsQhm0hSDZzMOWwBBNRL1+P7V24qWzEYC78hkFzjB/QxfxKOjeElJefkVcPkg
JWld4aWp2q6Uequ1bdXsP+ykRERc7HEuK4oqB+EMTs4GH6KugahyGhPc1KZlrmL3PuB/gEd7bKul
pPGJfFLYG9fYoVdMPFFiuz/4i23G8Ly1BGHHPOkupGG39OA/goquhX5gq4ifPLJ1+cLohJVCC5XF
X2Dd5uzWyQnEor4Y/A/58yAyP652oitf8rjIjnVme+D5t5GKoEcLW9A/dyZhw4iOuxXESm8Jbdo0
t5mS9ZsHthwtk2Iy8kpYdr4Ej66hAmUlj1hVn0StUpugbq9cxeFh8IGNwwq3M0Gw3U7cBAG4bYxd
EZhlqqNth3t88MxAczGCquqEUvClxuOCnRbTVhAHWimTqLOIWcauxXs3iPkPSDbt3lDqK8Y4FyMD
/rx5Olbcxe03PPps8ZqixLRKjvn0ZNstQyDp188WatmhU+LataUTKdM6QE3vnpgH2CW3l72jVta3
ZeKb30NzLB0IZn4B7PmKevSAjbdksR+hN1AGe4wrqFDRx02CMW9wR4mL7EG3d+Bza4ojxU1cvAPy
ALNbfx9oAg8FYlHG+RnTiGlq91/8TMMq7asUg8HZwC7fr48M5PtNG60M93Znf7fk9WUTmdoREFVa
CBwBtFhrZw1L1NbQRHZ1KibJuy1aNkLr/H7GvVM9V7+q2LUXhc16WqQBaQUV6P+N2daDMWJxyFMT
pWGrf4EV/uHxf3w4Sucfo5tAyudkF6IMoqlP6ZvlosZmcCPvjYs4HHL3EPaaMY0B/ZsFvVi9La7U
Sm0jDAnNH31FdEb656wRvm1F/jtQngRixcVBD99GFdhIhwKAB73QHHdqXt+0srMYDTSYbCnFlqqs
XIN8SHEeC2bp5OexWclSli0EHKtNTnVvQmI//JC8rq1Xx45OiMz5VghJKjqwKjlmMwDeaM0tG2Ou
eq4usCq7OKps4C0bTcAP4/xF5ZyjFnfb+waaom/B3KRe7QHA4AnhV6fhjyZlf0oE98eURVswiAMx
Lbu7qbTQyL9TazaEOlGb2AuOMxKUDbzBZpHLsgeAqAEc51d6m4fdbjh6l1BtMBK81o1Lax/rqi8i
V85dNzN11DnNVCqEWH33GT0g3YbE63dZqSTubniViHEcMTCwbuI8ktrdBuwX0TpUCwpqwSYAyHAP
6QIojqShd/pQybhxguziPl7cS+vNhc41nVmtwP8tJGSXl/vgEVC85YzEfdDiEsdWPZxbivAAEIvY
J+HPOWfQHkrVW8E4WjgyMyBhMPyBDg2l3pWvQWkM9c75zO70rmf4BAp2lZhxXRYpEowSltymDcfj
0nydh8lpjh+GIMT8anJiHFbtPXpxQ0XjM/nDj2ztoAOJAsEXTsmaW0U/2AC+tuJUe1+e1ffUpxPW
7U4TvTkvxPLR6Gu7L44pXc9FeQRcXmaG/POQzQ9IQBgVER3bUTP+Unn8Zo1UxLeasFyaqipKp2mv
qsdUrxmbVmpw/E4LM88X1flwZtRe3i5Ucv9c0QqrzpKX5iQCP+TLI7fSq/Ir/Et8GfFeGqoBAG4t
Jh6MtfFP3A7wDgSGZ/D7E3LMEIurqATfYgsJG0GAzCpClk9yps7UXH0uLA2qQAhxgray4ViMvxpy
GXMTaWhALKdYE5fSDoZV0FyfLVAWx+vLjxJ6zPRezVHmh2badHAY9te5W/MDJqKv9iMLgpHhEApt
HFaIlTmUIazrwGY8mFe0X9DFMwZNLcP2cOmSMOEbUahnMCNr1u4eDq2mGHotgWC9N06SufJ8+DFU
lf7RIuQvTRAZLTVJdjHDAup6DtDTXaMCcAFBB7nJoDuSrGvD4GhE3orith1yyIUGPq/CGRPkyYFN
QZyQk7FOU47T2hKMPtkAUDUsOIF2FI2qWt7Hqa9YOtqzYGh7nGfa6ntFCeDZIHJOnFfOYrSekwGA
cpMN03T31pNeMlwqmQ0/KQXbjHt0TzrbW0qJEn4UkXumsOfyM69QcOQsx8WIhupiuwmeuV61NcSe
zY2ZeeQIc6YHeVu5ziktmUZtryklhI1uEdzwS5wlTynit5ze/7qPy/8AOmbnenRfniYTDdDIauzG
nKn0pvTgY5tHqALrv/CTWcxHsjPviLb/sYohpSOa1GSEdpWJg2tkddfG7+Q3AZBRCcJKERe/4wRy
TKcFs6Yh1RcRMKc/mfrWMKLjlpfw/ZM+q/yEbSG4y18WCzwOKILG+SIlGjZeTLhWOE0xCvup6v6c
wESzUNLnH658B0vwXA/onnhZgRms+Tj1hLlOXrDIxRUzAYz9G9o/96hunLK53hHmAionzIx+BHWM
tCU+fml/2jRG6yeZB9tYKr43wMMMI6QlxOj340XxnMeSRfMgmkCD2NUxSaT2XWRYGGrQVC9QN3ve
a15/3E9AaU+Tfhby4Z2X1vd5HBOSPM65EynDhPZvb7MwZALnRXzuoGxvEM0Ti1llHAlj1WutaxRw
bA7rInuDDWA+6DDi5rCtF1wsUs3JCJgYMVheDOkQjn2B/8G5t8DPVJtz+nWKdcoRfwXC8j9yM0CJ
7OaOfTvAtA1lqcUOwJK8DhfgMIC40Z/GV5NXvndETDBFK99QQmLSKwx3lpLQITNx+m25R759kR4O
wno6BTsi9x0h5ViRE9EC3s61Y+ZapxA5SQvB9ekFRvaJ2lX9GoS6AcilP7xr5Lhh4uSwd2+PFWJc
N6rUxBMQi3PD4IZJWKvgPJz6n75SvRJI6pddmNgvb0H+Fic3DWuV3g/zObP5wuxOvLOqW0SFP4Oe
Gsxet3pkqtqbzTjNCgzrWDvkPDT/ErUmS10shagQiS37KhfafCBAZWWgJeK/cL9uBj5XkB5pM/ug
2Ij4lKWaIm726Jw4yNpLUzh8cX66LsBTlucmrbB1ZCCy7Tq/fPq31AMFfkNsJpBCcmu0Q29QMP1f
CpPYgzvYV5TSZc05t8ue3nChHk3fS1khVtrpSjmedgOrIB50aZG54pFAeA249mhR3hYZ9fw9Bl4U
k3+3uaQpNAcfU9I3Op99l+ZQdAF4CNVMHBFNyw0jVejTX9FYyjjqJT6duvqpyy/lVWMEO6b3KEIG
iCtV1pHyU6gB0tt5p9veCNNvsUN+B3YEKs5oz3aOwUWHuOMnCy1FtcywwW1JCwCMcidoB0KcGYQZ
DBQbLEsg+k+qmG8UL/kcMkka9QMNZjgXIZyUH2r82iLVCTN3YYku3mbkbzJ4SixLt3TAq56IdkBv
1r5zgftNyNvsKJy8I/UpQTDMDCAuTUK9pKSrlEPXaUj8UcKXf5cHzwuHVZhr+fHW7TJSQOoX+oHf
tB6FPIlVjMz/oeBcIRjkX5M9XAuHT8eZm7PuaAzCyy1oV//2bKnDPe7CECoOq3KKAZzef8sss3uX
XgvTIi235ryF6XZGrYPWmHy4lHwTa5BbjolDdkhUlEdMrCpREiXi+4oMd25JzJ6BvosS3+Mt1bxK
Rc5r/RsHw0JdgdhO3o/1sCEz6vVKOqk33ANE7YTbxKFpFBcyVrQn0F5aRfjVP9KIZledEDwlupJ4
ulp39c7hlXWxTGC07p2T2QdDSSa1rWKBSKMenr/ls3+TpHZVatFCcGFFlFfQFIbkX8Gctens6Gqr
emM+JvnPoqcbcFnr39DZLBQdE1Reh+iogLj5JQPeAcNLJoRyaXrVUsPfT5S8mYbVM5isKAWFyhOE
0H2uw7Bnwm8Hc9LgfPkNYI6ou5CwbgUXmjKsz/dElvvNyZsO3XNr66HzbywOcYmM/2vWnrvY+Suk
1AyeJS2ICnDh6bSiIzJtKtRo33g4tFnMA55dM6vbGHM/MidDl8SPyX/r5N+Ck1XFKBns8FW7xW/t
g/+GcVjwFLJAP7xvUPHvhtMZeG6Whb8+bR/K7JOJpsGXqEt8+PvLGuEvNMvQTCnd33b1O2cOEFFM
xKEUV++8A/itzpSbk4v9XjhT4/iV9UR/Jd8qEdUOHTiQiwoHvmrYlHVaxT3Yrc3614wqX6bfY0R7
uSH2RRkDt5i8rFh/YZSynBoANVgV+hLW50HycHIVRyHGPyO7Cr5yKGnM9usPiqkcdM4sYGR6o2FJ
SfjvghPxr0ffyAIl/SD6QfTqzQsdA0S4zIod8DjoAHj8qUvXgVTpBBAed41DIqNyTtGao/G+bkxa
ZLf6nAdIEn6Tb4tQguj+Mi2H9qVwai//XqXk4WgwZnYtCMXFEEk8vyvvKV14jcQHuf51jp2X6yK+
VKitPvO8Nu3nnJYY+XsvjeUEGPVlqRMeVeV64h8w1ILjYHTdzySc+9TnjlZ9RY6qalYCq3HgHvVD
L/1Off6cMZpgRZTXgbKm2lNe0R4HKM8lyprRv3Mue6YfpsUJbkUuYbismXJoJdIu11OsEU27oKTQ
sdKHB5AThgIH1XHE1+5CzaJmYeSXJipoKXCtWWZ59l8ZXmKz21PXtwlToro+41jfMTg8PCZhvXdQ
cPrWiJnJXqblA0SwaAfRRSZYX64kliTZMu+lSY0UZtaxK4Yp0jGLjJR9qtQ9onpokFtkMHCpWYvR
gNJ5MB73uakQkdC5CNwor5gi1KjerUHd/FFr699bBQ0QmCRzAopUhbVTLuVGV0SrfCvJRwXL8YUj
GAH5M7IQAK79b+mSY0PmslIgXZM6v/+22bM9hhP58/y6Wj5PNErGu76xp/jhL9T/6ef0GiXka5mA
Imsq6/rLyhBE28nc3yqgEUlW0iE1cRzoIk3QkUAZ5FfonTjcdBAlLqqg8i2kYaGkzQE77BvGncR9
BKKuqhKNwFlzR23p+DTEtjoch163ESlyQq45WvCkp19ZWsBilMf6OLpYxcRcznRErY4DY9K8T8BJ
ywGngAyt21gyY0akanjt8ni92VE35ioBvZ7/95+lDDvjgpIaTIHqPI9SFR/bCVFuJtss2gmRjpQl
rxoZZ6c1uYpQ4k2kfdUaQcPxGW7o6prVDne6ngzIvNWjHhYO3/Skm0cTOfZl+4gARab5mkXJsXaW
JNIOvtqfkdVXvPRyg7a0RD9f62CI5B3w6z8o/28UyN04I6mab5qzfJRu5jo07pOc9CLcun4HCA76
HHBIKc0t4/hQ21OfTgiLdMBzq7JMw8QuKswlnqTGqkIqG6xtw6PPtM45+SgsqlsihQQqere95pqG
4f8p5K7l4R1nCKWxbn+J8F7mkeUh7nEkMnqCwpYEWSRZxdqeypBAH7zFk3OrZBJJVscIkpn6UrDU
1NQtJpZRr9jFVUXgBq/EGtchHlrhNAss11p+MJEHSLxekOV9TwtpZ2NLwBVYlEu1ZSRCDwJLKHS9
ZXURb1Rnb6jjKfjhr/JamdaaNjbf5f0s/PTRnvuRMY+1Dm3ds028th2Q49p+GMo42IdizNtptJNc
SHn4G2Qsyb4RwmBSuXx16GeZ06zPF/aiOLDNVqDN2/6xsXr3O6fBTpEQPpM02Av6tyIQgI5ae1yZ
Fgs9mrkKozO8+iVyT0Fxrr4ceil1mYm9pbwVHyHCeZg0wL8tsEpWx++U1Mdv50eqzsr5lVsYkg0u
id1v9FzEadX+gF+JdKdDKMO6ZQ3ruAbRlTS7LZAvJ3/MPZcwOcbSRov4aGT7O+ikr3MNfVAmYu+d
3rRfbe75Bx4H/6JL7nGRYfv9b0ZmrtSx4jPf74UyBcXQRtLCvH2fevk67Xxk5zM3kcea/ePZYnLb
e2IOHKuQOSc5mGfRtWZxMG8l3Tach0pxMikvJrdbKkBZggupdQDGNVavBYJ73emfn+Jf//+BJDo8
9E8t7VPZFiFpExYUgy83WFs3uSXqgBOAK+KMYx7dVH2h69tDDkdaHQrHjB3V5e+Z7xrm8S8vPQbA
sokbBWzS8dwDaC2ZRaiePXl4kymZy5jOaOL7xSgYV4vX66zYGHgAj/BTANuLsWyrp9egrZKdHhiV
mybhxo7iVOMLlIxseQuWIHVjnJg8TuYDOoOC/Pgancdl7kDiURzgMGlga1qya53yk8q8QkpuygcO
9darc7Syv0W8NdwRC5bmFGpgM8zx/THlvREi7fqut5us99t2aY7oZVG3E6uyc0KIAYHc2BX529dj
C+aL7t6pmDf/R2MlgNBtO1U3AJHQdvM/3ov5DQRY9LmZIux/6O9doXxhWCsJHwv0o8JIK4IM99pZ
9YDNhTXZAmSJSfkvmTH3ehhH+Eql683w4Z2UBKJhvEluV4GQ82jByydORQhDnB2esr736IrYRPC9
FOZABTWXvtzDH/Lw3mzRD7xGJBx3RLXg8ePSdmVIoYXFpCbGdfFx7a7BsRrUI3TZW4sDViZpbvH9
+SZBM0Vo9T305gDECpiugx79d+yEm8DOavirq+4jYsXVHsxCRQXXcxDDwTSCDdNT5pH6Fpgu8uHY
u/sDxbqyLH4D8B9g1UEKuicyGHECQN2O0K5pNkd5kjS0KStmvsfvtm+lxBu4R/ZkdhFi5y21jyX3
QqMzjyP5H194POXDbtyn0CD6etHLs8DSXAci/J/+1Mg03DXcv9DquLfGULRlBCdVYgqd7Rj+f5zS
/kSHTHpgPOeMd64OzWdkgnCS1sDLh17M5s/u87tlGpVKMsffc+yKYzp8XzHNXfpyp2l/XQfaQ+Eu
uEfpMvR2pL0EphYRz0sX752qy5NrolRBm5/ng7sHn6L2V3bG4VyRVPYEQZFd87fvtyvirjbAvxRU
zrXW4v/3+jymLVfm09xZBVBcIcuL0/DPgdOg5WLd9lJp2H/i1XjStciXZM/xAHZElJUjoN0fTOS8
+EJ0wwfXQBkMlFPmNuRcED9K2leqY4Bom0XmGR1o7k86TdeIuTK45PuFdzA4QReoSyPnaCBT18G7
cx/rtuBbjzfRj9+fpkRUFTXGHwd0oJPVhs9okyRf5Te9R4c71/MVCN9mlDUYJgzdrUGKgZxsB1tY
OreBx9G7nwiMuhyc0QIKbrKRSsb/ZTWB7BJaiyYY1dEAgOZB3OtWhNMkfRLFowPAZUVO0nvbvznM
D7pLTjBbDoVllEZtwUPHY8yjf+qJhc5hC8/+TxULlXG+KuSzd4biGN7Tc78ud5w8lhcQ5KH3bRAi
NnHIgIWmrBgN6nVCpRcaNGRTuJ6uJY2YZIBM8SIBBBRMwCaYXLYqXoa70H9b70Ze9Ep91p9oGkS4
fKvgdxBKiWvdeRK+NLEtetjgNbXf6P0ihUrgtsy+eoCaSuzF9Ppw9SFiqmKnflLZ5AVnt+5CxZv4
cK4MxV8b++ml0ZyZ6+B8cJ0xL7XdEkfCSH4EzwcdKWC26zMQMJmzj7KtFnFI4ReFwEcreswc0Z5j
F53oSsbs5994Yvg9wcLtvF+uV+LI9rnrlwzFx3XJ+sf4uX50Ig4VI9dNKTkdvuDSPtXiDxtzR6Av
nXlpaGVCLwcZBjbv6XDQmkcAo7R7/VAW7gI+B9ogkjnZ+5YFibxfKyC25+OFgQ8R+L3L+bZrOwY2
Q+cR8dJcUp7RSubE+emhEFUZnTynZTP5DnK4aTc0cYfaNKTolEj9uhGKWW6IJTciGrUri7+wG3jW
P/x7iGGuM7/px0yIAiOizEhGoJGr2/DRe43uoySf+1SWWsj+JIT4/SgdrGdrXBgmu5ncWnCT8S8S
XHwoKu4ggsCAPmiypNKO+pqt3ETw2bx7xwjhBseY/89YC7At6Te7ksHrvvZ6TsX6kefoCoOwNmnB
Re8st0Ex4EI3Y9+JwajZcDqc1VmUNNuh010gCgYHRHvNPGX4nvBkfTiErmndVOzobGYrVBbn1xOM
eranMZOsy79IK8rcWgEtEJ/LuQvcCvgwR1y+/Dn70IDOavGI3jMwH8oq4puRMoJnm1XiycbxYw7I
ckPVuNXy71j0R7auMFr7YIv8MbYa8lLuobmldJpvxmbYAKwSRRwBYf15VHe5g9tjF7/KSEJPurGA
RxnCrD2Sbn5BzVNigntMNaBG6Paz75FR8EzzemTAQ6x+LpF1zwQGZvMpZL/XVAS4Eyr5VZsuc5Df
TGm8HzYK3LEEM4M00N2rppwxAPeXcT3RKKb5dzGa/3yUKmUwW316NqFKaMyD5MB6oeOLhLn4SueA
UOoMOalxcHkY1qamQKQCnYyEdA9NEi9vv4C9U57RO0LnDvC/F82mD+RBNuulRMVEcYP4ReQGnOx5
RaCtTjT4pn9b8E2EjMf9iaWSkq2EDOGQs5bTfRBYDbdpd2cKlpO+0+/e+YiCBX2+X5w7G2yJhPTq
slk5V8D3p1nuI6h3jl1nDgm8rZVoeCYhf9sqdnb0LFWTDpAdZsmUhSHLwsvHeIya1o85Uk3chYRg
80ip3pZu62oPmguKEV0MwOJpccbI1I2lRdgJFjwq2wt6MiuXKZGOPc1z2yUyYCO803hsJVKrmiYR
JUdo0xT72Z1i1Tw6FXNR00hCfMnR7O6O6xoBsEXcKrkA9WWkp2TaldbX16yzVyj7s/k60TCZKTzu
SUjTlUEyeniIZO8WO2KNklNcCEHfkaVpXNazUMl/2Kqumsmi5p83vZqLfspHEsrH7C4wLRDdOIaD
T0p7Re7eUk29eYNZeliFRcX8/6hfdy8H6V88X/Ku3coMNGrcJGmhCmchFdWANFeabA3jB9vCJqmr
uDg3FxQSGt3HUH47k500uDEW0K3zFH2x8mu98bS50/oh7RYP8ViLlSI1U2aBU95hNdSikVGZTevK
4+W1p8Uq+aF0om0J5uqozCMgvN6AfW3Swt/whISeMV1rE4GaEX3NIkk/aSsMzGWNaGMy1o4o2bhv
4Nx2NiGutJSzvEIMXjBbcPj5IyouljGA5VmWBPhX57+zuhQLr2ksd6MPmbdta9wHMKs3kzhfdOtC
6p+fFZUJsip3GOGOaeTi5xXCLahkYUiIpxB+cwjbXW6cLMMOFlys5tvvdMoiVwOpU+861wkWEY0h
6V6VSU8RbqmTI9IL3rEY+ccHCFurzpg/kuSpZ5UKOBYLnrJHN0D0ts2TYNoAxN7kjd9NagkD3eJz
saeJiZ8RdUixeqIiIqT9QGMWN1otJZZa0kEMlkqhA7bLge+fOAfFhZYyL/qNmmEXz8CszzlX/5bh
VP/rsIbERli0XfVI9tlporCX36c1Hm+5jC3kb/bAWxAbGyRge1utjGE4a408awKB4nNDAgQZOb1e
5mibFA//dPzvNveyxY7Y4JHFdDcdgyKyWII6i6ZmLtOhfXsuQjt1WQR1wukjH8tn11Ty2BicUi6M
pb82sM/dONguqBclfJrBhE5DAK0OhIIEhUvTZmEWnJptwPElk2GYnHfhAsWB8lf9tP+UqRLQZAsw
qExOWY7xpTEQLNoxRpPvnuzCU5g61B41Sc7UrdPQvlA/71rK/P//xkdAUtzwE3OBgiYG+QVB7+OI
dKwem3yhVxcALm8GpmeOGWauGqrl/B92Hb6mjw8hFZfzc9zm4/X8EsxgPJ2le2qiIMul2IT2XjSQ
u5qnxEIa39RZFB0hVcEQSQE4d6A+m5KdT8cwNkuENx/k20jWZxkGlgOWc+L/5w/LU4aRPyN6lyMy
2tDbpep9pCeaqQyFhrS2fF/zcSDBNI8jZdyrtpjvywlCAiDXhcFaLqW5EdXhBaA59pnkkI3/txRg
qHNGfaC/K3IsX/264LoKgZsCswTrW6SoES93J+LqAb1SZVEbdLJX0lie6+k9Blzchurkw/y38miw
Joov3KVxMQPtwpEIN4m/uJ9EQT72ET2mlD6IHx8yDJm0TQTn9mXVBNCsocgbXI2Cq3ojeiBrjHcR
Nu7rTmX86Z4Kl9DysmVP45Mxp7CTdIJHL78FgxR6EDmgClc2sLBqv30MOUHIkNz2n0Lv9dRjddgJ
QaR4QD+/Da0iwzyn6+oOqvj2r4YCQHYPO/L9saB8PqffMhchpWGlIRJXaRnauu+eq4uDquigqE68
qwoc5Ckn8VX8Si6bmbQRwgtf9eU/ygs4P2R3FROTybpMMFu/Zw7T9ztDIIJ3/ywTDwPci5tcFIE8
7ePFSptJKJT06m07XNsLvnCM/gDW68ycvZ9BFYf0nKUXX4MIO1vPoB4vhhuFRG+xnZg4LRCYFyIa
EIFYc3akHRk/g2IGtyZcdvlZhJcHepJ61MdXsVAq4+iyubjMUe6HnEwcvx+mAQpKeQq8dcZ1eBJW
yO2SdAUnAOcvIFmgomd1P5YzeYxjrM1fs7NHIdzJCQzwFgt78oCg/8i0cDLQQHVVwdJgufl12XQJ
93kj/jxDA13bRZmN35s3xGOaW0E9VAaO1sPRQPQKaxTIMKeO5q/pmDrDRYVxschchZbg4Zr6NC9s
ojkAr7jaFgghn1mLw9c3ew3kaZXqV1IzM7PDLHu9SJhEn45wHZWnHLg9BAqY3+AKOZWo2xvnMTCO
FHM+UhfEPvnGAvcejxp5BXnAxNd4kbjzlG0kAWw2dOkXGLkCHpxn7SnVsIEANpmSUU/MS9/CjfyO
x6Pcfo6N9MKjuas4X/+Wn7+CQYZTkmduQcrBQsAUW7n2e1mxQIQaVVMUQAvC70GAaNeeZUqjBWn1
zYCidEqaLaFMDZCles43S7+rhBaVHJJ4bapB2TzkfowxJbEilFZdzs7W+00o0vFsBSNKgqJJBkZM
1cgaF4CTqhdOzpxxaYwogSr5q6yCxpXMttcQdCfRG+kcv4X00Xvjsec08gwIZdkw0dtXchRVW/ht
OwUZ/a3nAybHH/1En22YBWj45wQMnJuMgctKbvYrg4vFr89FZpgb5izMccWJ14e516xYyPRpdExn
E+nCCyIdZLyq+LxnK+F1IWSqPyjCsp8mi9zOaEeW27Qkufzbpc5pyd1I45cLuR4zkKiL80EqA050
T30Zd+JLAnX2gyoe/GCpWMy13y2GPKQJ6qP9aGJjiT8l7UkPEsWddjaF71Mtnt9l0aNKRdyDvKtc
daB45R8/nMkoZWDT3drn8plFmPfWvYV73NJ0OdAsPpppkyPnwoMq61xJKPIQAxqRbH0f2l5gCMk/
KF3q0ligRW66+ArCrhttrKu5wbfOQQd7/BUnCmf6XN1RDoDtbguucKHcWPhR15o4N8YedvQgE602
B3qwGGA212YHvl+R22vb6s02K7Ykqf6AGf8C6kMYtaQN5rz0BbsM6tuS178IuA8yV8FinK+yV+Ik
dnhQjupAEyVTdY1wOzKt39oNCrs9s+5exR9mnKojROjciII+IaZ1KgW98T0cU7UQacqvP5RinLPi
4L51auox9fCz8KQAsqINGlWUr/J9r6cQZRYJ4qmCu4DZjt7OjHtwNt/CvZo51y3Ohx+4ZF5EJiG6
jEIBsXM19fAEltOjAuUjgHeJKSgxTjsv9thG/5kMzyCHaYW8O7RgIlihtLcTELtMB9Jv+yqC25x/
MjwpVpCQ7xggE9uDB0fqJ6Gj/TzoceDjpfiXP9pj4m4785BAyeESXrc16qmn1VASb/3jlE59606d
Xn17wS5sisoV1d/RXFDdNhOqPzK8we6LWnCbmBTK/TRFMUwG4MDguIw9G5fgvG2NdIE6LXtSPFDc
AdSe8otC5MwC+8baJPmxAS39QCseKo6ntQTPa9IdcdB8qtBXpsdYe0kNydNPkO6aE16GhNUUWINY
F2CVkuok3NpaXdUdVYo+DyXkQXzwsxJLr7x4TivPyZ2AePLZKTCKGPFZ+TvjAj9CGq2kW8DR4rZT
mi3WFz/uukpFgTyRRbLjMoanUg2mQJVqUm79/y8DtNDRa6Q0VQm0ITIKMe00/HhafJLPgp39hWMP
0Y7WHZETLXjTVqZVGHaudV29RNJKOlj7Gw4e8LzJqlXiFKJnL88GkO02SqdeRcDh3gWPbq+YiCjz
dzRffGjTZZ9fXdogWuSAmWzKrH0AspKjFJUMVAxoivkJ9hXgaGfTrpBWm2HuuWW36J1fpM6EEzhh
3sUsiIbln6FeTd1WZVEiTZ9mPMuOv5C3+6Ddlhe+jwYMGyx4+BfJIwIza1OkHpZw1ZBpMYDLPOgZ
Mew1PVhrSS60usDqxZvCi9Q18efReeSj6Sm5r0fq6CCwJTWe7n16Ow/cSwNNtRXiXctqusakSlCt
t2ArUaUj3j0Ruc/5WX8jiUrfeLiIRROpEXeoDJGqKmClq+s0McJnzowDJfBak1pFiVH6M8dYpsLn
BEU/75ElsIkmllEr8/G4IL6zLfEDelUZ7f0IWL06RGroPiwvqAskNvfuiy0zEdBCHFvVbhdt/RAF
SQnlPhU1wVC5okSUtZZAANRW6kBRwe1T45ubcvpy7BKMnNPFGrZSEafN0s2gnFS+JJRPUXZBiwIF
IPVXFzxi2uufKRuGChN3MX6Cu7ReGBfF2S/3LkdKm/Lwyfuq1k3CPqDQ6Oj9HCU+481mbNGfXbSn
f/+vFl8ThsCegDn+KL4SuzFNGnkpF0S4SxH6ataw82+5VeMO//27hFgWBtHva2hqdLwNadKBvkFG
Fm2DRfShzJ7zsn2Qed5Ujcq3hLvvjRFSCYzJS6yy2sszgkv8lWpbugvKzHt4jqKCoGkNNXfyXZa3
+mq+Pp3vWWoaos0tqGmkhBKq+leJcdMQd7iySzDj7LYytvGweXS7epONG4W9IWhAd66Y88SKBQ7s
QR306EX4XK83YT606AxUIM2o7h8rvqzzDPTBlEVDUso+hTFrP1SRuHC1DK2j6VC0m6xdn5mAl55G
8X8DBM/wYPacyVertu1uyEi9+1sHesu7q5jWsn7dqSEVVjmg7wY9ZBrkBaBkgjyOwwcXprdScXMD
fMAXHp93JhiMBc0P9lgb0G0azmri1W1ph9W4nv7Gvpg1prZCQvra59uYvDtRcvt7z+nBUQ8gpU4I
JsoBIVsTzXteVdMhSBpYzj2IU3NU7yhTyV4kf1G8J+ShWE6JWO83AcMkz59mwFn00q0kpZtroYnr
w9sy6sWNhynJuVzC1N8+X9rnAOHIP8Fb85HoMexvniDOkU/ItfyVzRw7Bea9eePeSIwGHaVwafZL
C05bE9J5Id1BzL343bXLyGfMIr1tOm5GZciZ0RdYaXO21okgcsnv59yl/AOKgnpO3yMK+vd0S0xI
6HkwWXdM2zM86Bs5/e0LjR/Ca5v+Y2J8YyR9llmukb/PdsRRq/IUPDDcw5WV0LLlCp8RVA1o8C1e
VXU5RXPcLKUbafVHXVd8GQ5r/1B9XfIrXYXd3awiIXDYeg6jVond9rQeERxB7NJewIIYoz4Oq/Sx
WxwWu6WJXuUInW/ccwPkPwxDSzB0YutBT4nR+RDbjkG5qL7FUmJqedElt93LHUbzhGOGPBmqOoJM
JUbkkhdZStg5sVe4HhonbJYjIz2F5PWT3fx7BR74Mxg5ckTRRyK5bW5pnVdKFIbokmmLN22/Ihbh
gZuvovWtyktBFG+kZqK68IvBtk6nfF4ayN7RXL3fym9+Lp3R4+Tfdht8u3FUcBtsLkk5S8AZm8lI
CnU523hIFSAgP1IUInd3P8DndZ3sBzjvDaUBgtHP1gH1oVXx5e0Rs1L8Rv1NhYyIkzjGK/PqnkZP
/Xx7qcPOR8PLTbFjDNp/ZbE01dOwzuWXSNIq6/Tbn3YoK9HHtJEVPqivkzfcK89AuYsSL8NLX9ER
J39AlfLbF451/6CxxS052+/KS2Z9oozJxFne5jRs2dk8nbUyB0jxkeh9zQgdQCi2h6sXjxLxnIwc
3ca6VInMvNKrpKjGlB29z9V5Qv08cuAXg6hhk0I76/h9a1NSGkFTp1zdjmbWcshamGMwmRkofjtT
3yrRLHTW0yH7ICsPUH/LGa70e9L3EO11uNN7gEtOif0jkmEo8zpLhjNSKGHS7NQgqo0sknYU6ufz
Zm4y18YTd7/PxfvRu9MQ7oVo4grNdvaQTgafrUHFvx49/IeBMcSCBWrpaop248Fd0Nl6zoKu+OtC
1WOLtTEtJYraESkmPBocO9CNH4stS0ZAoH6ky9Lu0AFfx+ojX08MDvAlTFhRUtPqCOtVvmewzcGO
/JT6m5f4ZjWTUDBIv5MPaudKinv6IBtopIL46rTrA+47bG2dTydwR+xk/NiIhIxBNH8ow0beFsnY
ShAT7sg5S0avYCslmoHOFPEpliQY1f7+XZDuIqAN5pXlC0cwL3PBLB05APPGF+/XXT8/wdgKKTM2
z8rmM+05iRw5PAFOY50ySNzTeymv9YqTBxZ/yrQam0c3uosx02D3xFyBrB7KoFw59rd7Rf6Hw2bm
BWZzw0SnCj35xweGJ2USMcV+x31z10S0gnpIhBPqLMS5KPQvVCA2OUxPHdKU/Y4UhfHWKsqd4zQe
lk5Yko5rGxsIFJIHWIJJcvhkBdprKEz+yrt76vQ/ssHObNojkrp8zDzvq5JdIIvycTYwefvKIeeJ
aC5V2RO2yHj6NxTlJeEzRt9QIlFYxEjUAxGAxYRWqGit+z4IYEeOxvXLfuH8+AHJTMpa/DnXNwy4
gbkr8RzxrmBA/oYzp55eLD2hho2vI+4GdttKJ12sHgzsS15M8eoA/bVY4sbPhflmMn++D+t5Flay
ZhwlEsMTCRJXS3UltOAW6mFDVY5iKR8yL4ze6cnq70FF2yn0r2+qEnHfsLMbYQih0whzgZOwzzfr
1eCiMed9UJteyPxZOfajtnMxIggWWviPZqm+liN8HkTMFbL5wc8snFL1diWD3/QakB1IL+iKaO6u
Az9Z0Rdo3BXPG8Sy6+CiSRjkAnJDH3tjIWNmIMLi/rG1iPWYtQHM6uMGP1M8rbSgAOrVttSrSFK0
PTezwdJ+JX2NRJ9Y+/3lurUeJwcKAmVBoeJeOtk9Xm21or+qIxu9zylYill8xMgPO9YmA/eq2rvj
fFX2IEWQ3pn0DcPL1/fXruewBvdMgxYoxgws12prfgda5O+62o9BOZTSznN+bdOw5UpuB2GDK8GK
isMoVk8loieTTPaby+GjXMuqRSkyUel4Ff/Qzq/Fx8LIQfdoBzVPBqBGUnC3sG7Q8uVZFYAAjSkZ
3kcWEDVw6b9vr5KwWwhFOcekD1qtZ+sV5+7qwe6SxQdkg8D+erTQ0rZeSdZT0a8oefh086/AU81L
5rd2Iq9OoNIh2ckd0QAJ6pKu9PltJECC9KKxaD5OrU/agZyCSWZfBejP8eQsLWOYoY1yL5fe8q02
V/3ue+wIkHG1XGc8bf+Kw449jl69N/Xyav081YHJ1Cg2mzOeOa0AUc9+7a1so5FwiYN/ti6cLVus
3H2Uyqa8lgp9dnlokq/v21KaqlLrsEN18AxT7SAbIxcc1QeJrlRn086cIcU+1OV6hIaEUepDFdil
AotY1fq1Z9rf6bMJv7MbyHzLdKiSA/RuJqIPFmTEy6G6M/ds2ZfZ8D7mmjio+s5sNioBvdoxV6TW
AqI4kPU2esLFiKXqx0Yw8BpOZ9NhnLlQHucoz6CYeVHJ2tnhks7ZsgDLpPON4cgiMKQUICXpxNGc
fh8xu+R97Ed6JSJYJxYMwUwxncdt18ZDtDokUJOWyzut844fCcgFfD1VwGWFvH7on1T3/2xsgNWf
LdGW2XioQOCXu0wmA+IHQq3drABUNl9Q3doM5WN2x7Mp2dbnwCQuiDYuAul0iedtiBu78KrDSS4o
BTbU5FqWm0ITP86onf4dKPwbUe56O6pcI/tLU2x7y50yyXYl5TkxnPaBQkeQ2VFWDsHoAAoLA0AQ
fPsjPDV+DXkQdZMSnnqfK+/1OpntYsDdKkM2NZR/Kfnln75NiEtCLJJSqmyvDkQ/2DaSxEebh2Td
LzO3JlPpiHC4Krs85SLqT83PfKirYf0JIVkQRFEDbHmhNjF5CqnETCeYVJoEqs0nrHaI9SVJJMHq
PFWsl/dPDfKUYS6hcqHoAYS0C7AlGulsiR6Edujlk2tpBaGLjK3A9KNdY2p+zgpaJiskv4qjAz1X
879bUrNVzq0hYRuiDHI5PMJQn9K37g6yh4nkf/FXvDqOwykdK9H/Dx9l8x5kQXaB0pCceziMAbCn
efuUCMG3IJxOItFVYNXrrbyMDccWAHa/voqoAQlQS+S1AALiE9hgWRJ32qXMNwn1fB8LIWwA2sZe
T518hzBDFsIhRsCQNYK/Cphj08gBxSzKtkCbRArjWnDdXEaqrq9mXXmVXg1g7d7TzEHLHaWa9Snb
bKfP4SzDfPAPzIn4mkb2Xi1qx4tZCdN3IL3zu7MGMHs8+soifTkiLPGGUzgMUuwKlIFR94MZH49y
Kocq5D0hZ5MVXRxuSE14F4v3QZO5CdOFCXsSTlNHKuUvm1V3u0yfmvojt5AM7VleNzd3q77aVS5C
gI25R2YHNokm9HbWr+aDTFy6LEus99lNffJPVWmdpnDHIUn5ycwy5OtPPvCdu7tWUDegIIfYh+vb
5xK37Y7tD2MZBaF2EwQt3ZBBTqERUfyNqzbIbwCsisDz7Y74WVDbEJ/UcHSg5pRx4LthP3XBmx0w
nU3Ia5knMeC5hHn8aNYa0L+aaThjsCLgguIya7z7MEtKBnx6TevDGYj6QcC4EqtgDv+RSyRhohA6
Uy1Np0HZZj+XPRKfm/t8tIRh3fMG0rSp0XBEm8YAcZqRfgn6wRMF8argtJi4K+LslmtudB1I6dVx
8sq8ixVedBEuuFBdTqJ668Jv6ApWc+wygxYAfkxGyTCmliq3bn9wGFOCWGGE0ZBkk/S51BK08qXl
Bpk+kwQrk2HsbJ90z7TmdGm/zv1s2TWQNjnVOnD3Oyyil2hFbBKpJOZxm3M8jh0pOs7u+Sdu/Cgn
I99Ky5PQlthM/pRNxHVVYZQYHj5xXoqDRN9TBL2ATheGGobv9nY9y9ldzSiwEv63Y5Bu5sGUPrrO
CUy0/tDrRKZIpmXQUkRp00QZ0B2BHA/IoBycpVBB05IUefIAGvtVkY3jwrNsz00kS8Ujweo0bMeF
9RzJRoULCuOeYBqs636nrma8JS4TAxH/xY9Et3l7vJnh12gJuo92MYMyiIOQvOmKm1QhUrcztfru
L7idUUXfx9EZfdy/mlk8vqootxFnlkLa5ah/s4YqtEBzZ4wPgUlh5HL92lSy1SBUi1d1Vr9hs0ck
SLwnhBVfTmtV9wOmdxRjLqhRJO6wqpAwP631sH2ZUl/5cKwPB3HWXpfprfeUKyHCxvlRkaANOigr
igf+MIumzUZm7qzDgiI2XX/OfQWjo7TuQhHGbWA4nd6EMnlAhVv7wkT4QQVlE9J8DgcJTOxCay58
BybUCNxc8sYTiSDBHd+xlA4HgjBPJevpY5WnnA9BzS+i8D5/TP5EYPU+e3PlV1tEGYMT2Acx6xbj
MSUd6GxeRSch5ijSthYYmzNzgDarppwecV0uvKXeoSpDv11mCnVhNGUWhHmGLaCj2cOHOiAXpV9k
l3byfSVHlpXz9Zl0qAmNvQtU/+8sjZId3oVIupmqe8A4f/FWyrKsMwIUIj6nZUpIrjDOBjWX1RGw
JvROLLNsb86Eta3QNJTNJgKTEiGghXhmAxrCoDlU7FG+gNA22mSRnFIPfmE8cy7eizmoSQ0WGjN4
LxotqsEdemUr/iLpgGUMZD7SnH9I47Z9RzuCatpFz3q+pMp38JwYEhTN7d12hhzIAks7lIfjfE3u
sljFF6kk5/jRAC0Epm8CeDzlZ5fX1xem+fwhQ6luUjNLQ3liYZ85qmhR13qYKJA6YPcEhzN0GT/b
O2NYplhEXLgtsTLQxGnTpJJXJLIzuU/pcYoXDkUwo1S52a9xwf1TME8WCMEShMP7Ofozd5kznBEG
Pr1NU0gqwgmSUqjUgJolBa6s7788VC5f4OCAcfBdcQuIUs0NlLEWBFQSUXxl7cN7qyYq8bnTXeUb
o7bpU8aIkGFyXmFGt4Y5AnT/19YuFxOZMBEMcwACc1OyPFzJUdG1r4FksSJI2he8tuFewWtvfwvz
Lh62BB0WHhh2+BXhhzQcngavha2g+3iuHevzipqvJOMpo7gGSYqgceNpuyz0pTLBj3EqM/dcSpEJ
fqeNyzlfTzRd7sFUmMIaCdyrYZjpqgt5i6jFpwlzm+xLw/KS/Ey3IdXpTjWwMYd2MaIDi2T9CuV1
Ibb7HcxMHWK3PA9NHS9JoB9y0T9NsyyPSQ3tXHCTKaorHMvwGcbWyT/h5v4sqnyyHRI96mYflrPX
c0aKLClpX0I2lAO0RZZHUtapyezCLIGr/OwXRcNt9P/A2ny6cXY+T0DJ4ubjFqYcEZNeNQfsyEpf
6kXR5cqL8eqVS8ndmp1pa1FcsewlLFgKp2RQaRnYJYdmB6GedKU4u1UtNaVfDdPMpgrMpuM7oHDi
n+7t1ye4T49nT1Ic3qoocvRZkeklIh8k2RtdFEE0ONd3nrPhn6JFV1knnipAln6xkxyE6ojhTI/5
xKiT0rjpKhaFAUYJja7+OGogzNAAet0cuuRjor3Qn4LRdXSkdM02KA9K14xmkEMDvn5g53lCrbn7
+tzjbJGqzHfFPIsKcfg/Yv5eLaWteU3WEZCWl/6DNvpr2zfho1MQAPc0E5PG7eQqwqcDcx8ZztCR
H1+QYJ+Ov5cC8rI9EP+XbDmu7foquSPck22fcXufRAXDCeaxJCNlowLaJdIH5n4ctKdLw10/knx7
/rlQRD35jWlNQ8mlQJdiEUO4L3m2tlpl9UZ43yu5YMxucsUBNFxeghIHqTutojTvd1w1jfq458lg
ieHPVd7Lg2vMVI7//0dp9Dt1ZTp+5545/GWN/yN4+b9EivCzSYgDTcvj4BqnDfnq0J9iQuUCTB/S
jMpe2UFyoCbkNAMU/u6//Z/RMxxGzfGjiuiTu3hhcbfJp+krpXYRf6GnUykxCP3gctY3Amakqrt9
uxfWjOIeDPupNbPaemFoR6sqLRudladE5h9+TebghfYqK58xKpyDOhnYJ4e5ZvW1XsR5YIznpr7J
nacjgFlpPUzD74TqiMXUJF9gUyHo8JHoIDYOrsbaUXKe2cFszvsraSVQHIRM4X7ZIYzeahs/jGQ2
NfMNKA0FENaC4cUXhQu8MOww+SfKpi55NJgoOREqn9K6xQEbHPLz1DDLavpJgzDFvIYp18jK5vfp
azaLTu7CLB5SDt5kY6FNHzSDDSn61w6x1tc2QUAQAIy20hCaWRFclUd5m1doof/YMY7rVwlDyIf6
b5pYjPPUKu6NfUICiCg1WaQX3iYzbclDot6GFae/29pOD+kWFCkjs3i9XZwkhpaPqcVRmIhHI2oA
7i62+kKgUFY34+BmB3BlzgYlTh4VQ56rQweay41rVlra0ShMc4AP1igCcZzrWyhVMWYnR6saIeiI
1lZEnma8KowfbyYlOWupImpbhbSSk9b6mlQJatVukLKqBtKkfqvcHVGT5I1W2yWAo9SUVCCyV8q1
x9Hqnytp0J1Hjp9g3Z3RoOjOEg7yr6hsn9OhZpD2mb5bWMj+ZoYvoo/+SOh0gdiEr0kO5vCzJxmX
k96WNH7rjCV4SYTXxCDU7PSyCIwiBS752i+rRvTHzF9ZZYjoEhXMkqbo5YPb+37hvvg/SpMhilk4
ksue1kzFzQk0JnEH5qvQaJ7UkzGiI9/UdB6lYcIbQ+aFWZW8FasxcVdXgS/zeXJezEJTaXMklIEq
ShFrnRiJcSUDn2rJ6CgmbOKo0i6utXjWO1SuBGhYyttCwdNiHsSTiP6jts8NHqd0ySAyJyd+5G+N
M86H+8H4gJ4SuL5+RcLvxT2z+/Z29CiLTEcvpQeDQ+Mwiefs4hbY0z9lHMHcR4cVPDbaR0q+gKtd
aNAyfuGC79aC6thBCjs1Hxtpyz3EcO9AbsWldyEpli/16gYUsjm8/3dd14L1kIj975gg3zJkLP7i
aJpIhj+bp7uSuq/MdvD3xknpXqyzhR/BIc/Ncdw9/MiZAT52i7+yi9nWmhL96L+lELoaPWAAjoxC
DTSDUA8PESY9mYqzKMMteL8DzWVSK6N/UvA2An6ux1GgaJXlT9Rq+KoVa5IzgXVNHvyOyg8Aw1KP
ym0ntlTXcDPWj1aC6XIWiU4q1K57twPwx2CP8oE+kkPj08uI8V4TVv6EYV9AYcUSdQyttnZbQZ0E
ygSsuhqdNvl+4vpngOX/MwiAhW5NcxgVuqeM2YCI1n+XjdGJXpzx2pay17WpHRyt2+yLXXEAuMQm
0yFiIMBqkPrw6Kjt2OxN/xr4rokRV8e069wSl3XbrnZahy8/SRppujprdpZfjSXb6cHGwrXlNQIP
MfpiAh6yBPd7TpSkVBH1ErE+0Om5ehu5SzXJO1aAExyyksy2gwA8h7IO4+x3fGrrhQ+Bbxul0iJt
ZuRLKz56P8ktne4RvB9DMIi3psyUx22+sLkpdyl9+7E1fsN7OZuKELzPRsl/A542hM9xiZ5vo6vJ
u9sYbF3CNi2YEQoHRRVe/lmuhc3vTiSgbTMkLaTdx+okzOcMDp4twpmVWWXItDVoESh7HtDGYeYW
rfITwgJCi8FJCm5fecJ2mRUzMgDj1Z26TMjwXsOcZcO9gHOftF299LivQwMp4FE/r5TvMSWovFj0
cKjoMUfpjVqTZRgabEvW/gza8ObiPQ1KlI9OBIKWUYz3CXYFCtItScCfR1YsQ4CtW5yzfY6ErX4h
mrOD8o43SdSBM6HKvY9omKXgliWvv4gcdotwcSKGiM9PrcZLxgepF9aZwGK+fe6ocY83N4lkJ/xj
rTx9Fh7ZFw8TPCfWFFEPf3Ogaj5Wkj+H/uLodsfkqXcvwnnLm7gzfXM02qpL1OFO/qTwRXal8aF7
KYBCOiqXbSzPlhE2OVjamxzysyb8Sui6QCexx8gHFujNzl2AcHS9ruRd84eQURFBywa++/1kGFZN
za/8HRdt9eb5VDBd0aFJX/KtgvanOBu5Hq21oiiPt3S+rK96gOIEBG6iKYQt4gRFSaKoZLcyvITI
1OBbEZ5Y1Ah1Hd552W/AibO7Ub0LZ6u197omkD6Ch9SKcLKc2puCgOG6k/x7WWgZPYPnv0pe3/QN
UIVQKppP8KpIqH+S2+4C7JEAAAdRlbqUOhmG4gaWtilPsCNKENw/rQ/L1uVh7MQF6a9ZwAdvCWIY
TETmyY6uH/muvw925XLz1Lywzh/A0kt4JMirV5rTVIRD9VagatDKmNQJIQkMs+yN3jXdX+/XW34C
XJYvl4HLiBaBSsI2ciYppeXdM+dHFF0lFMnbOxWS7Nvt02EtLGQkRNkfXfdpoXkmusdf3tfHIP4K
8y9Nex46dlM+/wrXfrAUEiz72f/FKqxmTnux06wBEv3FSSsW777Q5yte2uVr+mcBAig/9YVdjJHV
FsJBXnwUUWt2SWRS6tVxiZwXwPlK+9V4wLJmIXLIvNfPOGxOhYZO8mhnpSJarav6KKwZx1BVKmrl
GbHOP4iVAVlF3WEDEo8mKmvmBwbALbFrz8lPsBjJftFZ6U09bCQjrSVkHscswEn6tRjp5i8AyX0L
Gi/umQbWwG45j0I1llFlr6HPFbilwspVYh4AA6ZfCw9lHO1hxHzpmNFDooU0/1MN+0HMIn0wLyg6
HRNUZB+1R9dOOgotWnXsCl+XYNokW28AROLxmMa4XNQwfwGJCgdh9p0bbTVFezTl7QZ8zi+kiU18
DbF9OBCUtgxdziJauopNlI5PkoOsrMrZmypHpBNHrW/18HEGbBG9jhcJJES+4yJm4TUmxKTQqbSe
r2SG7X9CWQ3wI3Y98TtZTWN1UcFXD4pj2G7Suh/1+RPtinH/dpcqc3LMbPQldv8a+WMypSeo5293
o1a6/xZt8JhcGX2gWmirV5WM8J7+f8ig/9nF2FK98pJmC9aa7WzagC3B8HIeR/mZtFOlD5sXrXZa
F43EM5HMH7S2beEJOZzSG1JRw5fLkexuIc0fX2hwS9Wnc/Dxnm22/3PK3oi3IL+dEf+Epc3jcOIV
ko3eZwxy3Xh95fTTX+wx04kMqTt3djgOam/3OMnTOslX+gHmJww4T1IHVYYxg7akTXrjFHgfNkbo
O8syrUsIMh7ouQmSvpOr5Lxih92rNzfiI+z5zobksAoCuBsI7wPz9yd2VHnDmImIPCzVQCvsHZgo
53GjCqTj7/CEaNea6HmeKNtXTZm8vLQ/cNT0B9dqS9Bii3Hu8XMWaJ68gIMLrifeARFuowWXkhSy
WAdcWnHkjbP7YmuYvVCwV05iEnfpioCcXPylQ+m1GG4Eg78l4IBTPa9fjpTR6k0U6jIZ3gBKQa9b
NolHyNvt9SAmSX2AZ9MrYNyOtHeKxSj83OWcb0c3MsCx6eXKGYtQ7xASpRzujpNDrkVxdUtYnRLe
qcUpLIiuU4cN1KVnigxlwaEfZiVyEwX2ubJ46XgOR+ENqpu7Owazn3W52GVPqT0tQp8XJDSBRTFL
Uo8QrokiwXMOFHAq6phhjdZtO7nIJKtMeGOvBQUyUT6baxVwn1RnQb4rWU87ZPHi1L2pwv9fdHSK
E0LofJZm+AbCXL/3vDflasWm6WA5PFXKU/zlgpArkMhy5TPVqTr4JNaUu72GF41Yj3AvrrCP7Y4/
SmZ3Tya0UVJDYPnCIpMRAJtipVn7ykT7m8Tq11HYtGa7ZECTPw+3BAm2SGrlUqJmx2lPRuz7idEK
SwFoGCrLMtQ+nUl+tdU/3cFsqqwjVR+qZ1T0kVELVH+1XMnV/OlKhMci0ZZQtQ+uuV2EwDL7omf0
5yYygsc+/jxMduryF+oXV7T0J9fbk+yl5sqxK8hTCoWanZrJRNZmXegFt1gdoNLRpE/onE4en1Pk
rHkHw4zW0F2hr1Z+in/5UIFb2/qWkxG/A3i2yofn8rT+0u85qnfK44g8rjXZrVZhNP1Hj1YrE6jc
GOFmxv/AZsAl2FJSVZ56BteLYu7pf4IJ9hkvTuah8+GkZyuPYikxti4Nk1OA+AkWC1ldFFf0H6+W
SH58EDaF3jZJIWaMrh6YBHBs6Wdy87Hxnr0ERiGUu8GU/pZWChsofQ7QCYgbY7t1BsfehsjzUXOK
oGVxMaxBgIo4qPxCSXzaIMm80JyJaF7Ky01jnbuS2BdE2hUzgJPlH9V5/AQkR2ytcLfNsN96YeUz
Sf3QgH/G8PD3A18nZZwwM2wALP+i7chGIpskDOfJFByb0zQDbUJfsQ3Fi0jY1ahjDX6S2A6//Qq+
rOnkeApKxygNOfi7sd1ISwQIjTUncawAIGfbm45sT90zzEg5XFdRPxd/PFY1o3f2OYtkVvQfYhx5
qd5S+q7q0a62DgUzjYzd+qwx8JsK9QeJ/gn+x9OfgDVd1+Fzxy++mkUIXvDxzCUKTh6QZFYgshi4
G8rZGS/IpxhE+qMF5TbxkBBbG3QEZHupPDprSCX/zz09oi6llMaxab/oLOjHEIarZn5QqhWnhCBf
rirRWJbIvl+QtHWyFcpdscbzdXREvsqF7JLQ3rMEplKoJxYOT05alPiw4oVR6Z3u/GskTXOuwWMH
I+i5lfCyI88n80rrX1YipeVvNEGHKzBkopvdsHThbObU/lCM5OaRlACzDoE1FRe88aTW1mUXNDSE
6JNiLiAE4bNHMuBBPaP2+ihRdfzslghx0ABlElVPOFSbQIZ5it8HmFtEnPHCML69hui1S0ZfJC0I
GBq+QUWfywkZcWzRyn53Lm9c9pPlODZPL7usuen08RSGHXogxvEC3oVucZZ8Oq9YtkeClr+3x9aG
7GEyDTCLL6KYmejxkn5Ye89nrrV6KaXygoM6rUdtokG9GlkN7k5FJVNHmi+/ilDc15k3p3p3RBJ2
Qy/Uwzvidk9blNXMYN/y53+HqdiNvXAKyrOOooBgj0ySksmXQT+X92R/w9RLrn6qmFEmtzlS+XOZ
sPj0SRNDFLGFkInx9b2MNXh69v6dU00/U+kga1cskCug6+bq8pyTv1BMDGcy0rMeTJ6yfY7ikPze
7S0GuaMSI5PLYE7Gxco8Gj4l9Dld34HyM0YnE7qF4+nDCR2bDBdp5g147L4B/HKOfhtOosgInf7A
oI0CIFVjOyYN7ZvxQC6uZSr6IxqaXj+QVZ7QDAx0dKI4+6LLa/ciE7z7v0G6+woyTofS4oe+luUN
KtNM+me+EZ8Fp4E47+0QPDfrmKr5rq7Uwz7HThSR/pm2lcYKPc3jsmJRAtx8m5Sx18LXvKmCuaDb
djZ2qoerEpc6XCDGFSZazhR73NFoNtvvNG2JnWJS+kwbsX8ee/cf++uPluzyu6pBf/qzIJrDgozl
qhISiB9Dv1eGgc7E+75KKvk8IZn4gD7KF4/PP8HEcc4vE3jp0jSACHi1zL4czUcaqkLZR4hXaE9G
F1c7wFIGvcCYTE5DypGMsd5NMRdc+6IXjLxGBe78ph1MChbefsbtYDj0mP9mL4S1XATFoNLRDAlP
QbYHIV2+Fs5QJHXEMQrlgYzj1MQDaycCxFXbIwBf/z60TM5BFid49LpmIfPyCA7svHlGwCif3qGO
YWbCPs58QS86+pLHwt8NFYRwe43X6r+zSD4gOH8WfrFrTSzJnJE/9UEcEK/RMkVYSzKalvfXQWV7
Yj1p6ZAaEQwBVhT8Cw4F90EIVYZyIuuUsIDSwp8KEG007x+HQoupsDWGrxcHCy06HmpviYNageiv
Uch/+KPCR/pi0MRNAuv7biRXGAqPuQ5xxe0e0xXbNZ+0wf4MsSqFEUSmpiIeZvgwMhfokP089EWj
v+Ke3OwndX+7A0/2l86jj+Uj+eaBCpT4ncD5DTJqG55eDDWob26xBLBN3RXbk4Gr7WSlKfzItVEH
if0lEKbgtTUkoGGOUEh2hbfLAyqzWcK+1AAoMU03Zcgy7ZP1fq/kTI8eMxmVbcB0hMQv49vphxJM
ZjYM24Gw6fz/wSt61jorQvO6Gf6cBMG/oYTmnz2e0r2Wo3NhbgXwufiFuiS1EzLkcxyBHYHVB9ny
Ans8z/kCnfBv27mHw1F7JzG1bVzBVT8b7IpgGW2T6zOikRDwZAJcl3hG7IFGZLxU15P2ZMJVmmAw
5n9OLTiPq7qHWcKu0zO8M28ZFlU3GUlqnARY1Ubpz+z/pqcIWJEWdYux0+63yv6t8y5JonXsgFWU
uL2+sZBZ5W/kBEh74+HFufj+S4afYyB+avmjQvJKaHerUKBjuUuK2RBsEwu6cx8QruXh0qwTrKF3
H2QvVzom5xdnKvxe+4etDn9BXl3MlV/EXqPolV2DaMqCmNKbtSFL9phu7dOjg+MYCFGluvbEmfT/
Nr5MtY6Mhh0K109qzXZRsq3fdiTHQUQnEiCvu4k4wWNHClkqqKTt+ssKxoQfYdWWQXGqqczfgKYl
eOpxlF8Ozr4xv13ndyjwJdyfPPbJyvIKSBuXOpKoTwMT77nXCmUdYarUi6bMcjl1NdGIzJDzLN79
f/EU3gamy+iJ9nwoeMeTSfzcw0LStq9w+SNseJI5u8pgTlIS+HwfGIPo3IW0GaAxF4l71tSapNnF
WaJpDWeY3pXWP+cjF8z6q7BAdK0/V/NezRV61d8UdB0tmz0JQtutUS8/+xls49AeC5m9hJ8l+wvc
e0m8TXOhBuYmSJ3mWyxC6hr8HaweNFbXlkozZ3vFv720XIgKFRG7hFMWmngumjbnosy0VAcc1Gy9
vHLNUKQTvRNdHon1Y2dNYBHuKVhbm+MT80I04/QNHY+5BR//JdZqSYtQqwqgYVNN7pYCfg5x72xl
JxgigTmmW4quJVK0W96P7dyBIF+7Je6IJQXFd0JsJv/lrmc/g4VIvgeXujgLycZAVYaHfE6a3UG9
YYfNyVJaS5BGO/NMLLte78eACSdYz8NQK2GFTdNwwl1oZ95qwKhGiZjeUTkYXH65R+CvcpoXYMdE
b9cose+V5Jp9rkbyTgdejETqkwQRjjdR7uTIwMLX/rZ4INODdDbFHHVJt1qYe3pcNh4A5BkU4eUi
1SG6oW4LJG39xfFsa6GKSSGT4ElTk9M4M4lzq0mGQuLbgxHRftREUzZZC1texjIp+tJA/OL4IX0g
8arXStVp5M97jRS6ifGEOosLIQiNGgzOtrumiVDwJFJlHn0h0KfVmFzGRfFly1IYdrFEC5ASoPwZ
Oy69drQ5lzJXBu2wDs+0+WBamDpuK2X2pR3wKxmMjECY9E5vvIgqb17vfRhx/FUuKEAe7easDLdU
nYxpycSP7VJ3j7mxuUZqvAWZUzVlwOaNyRnHY887mk40AbetaBo2U6wlx+DTpjARnN2hIm3LkFYo
II9oNeb8JvKOeIbntUaEpFUvVxteK+leUEkWkEpa1g08zOPX+wTUewNUaPzMo4+5uX3VtP7lckPl
SRxew2MpkUI/pcpelXZkpXQQt+iF/qGA5iZB/tgx+5HlJroCyTRLJF2KrCkCSSJkmORaF51Eresl
KEMvi/hfl66ZiKTN3QLg+Jfz6IqII3Zj2HRBhlEy+OAqgkqxXWcdLS3UOR98G/QZ2cwQqqXNKePb
KXbKudnypqTqgxWlMxzKqYwLaJagD4ftk2HyYhbqJnjWjl2N9rzQlubXBx8gS64dRynXQb0rlUe8
VusE2esRvnF42YKjv0kQj+ojTh7PKKfPaSqTIbum12cvJRXWyCwCBCiLnuysQL4082hu3xHd9esT
5XLsMgsnjdFbdbHingpQbB3Qx3LqHRalQiqwLdz+SPfSyQuTeXbHNE70xTcAOjIkI2ne2IYhypQd
LnqqnDg5C3yiRKt1tKnZBvsBjHs4OgD0liN4FaGnA7qu/g/O2QsAUtC2NY+dN337uzY/IJJx92K8
j9y3pMVHXqMABle4ozTS3vGWLsHch0u7LcJOB66I0d1rw3tcrsOo/1dV2fxfgci0YM37L35Gipxg
4kNVo0i3o5uTXWToc0ZXhvBJ2/6HQw9A1HVko9230dYc+Cg/gLVSMmCUb070IQnpagvp6U96n798
hBAXam4mVll/E5gfItEV0ZkRFOSpvh6BqsSYlgjJlfVezUNiv1OxjnLjmgbLV+OtZSK74juVcgOu
UiLrLXAeWos9VghWwIYa0hCak8oWKHBAUXmVZN9zGuMEAV5TBJzV3amB1aWI9g+x3P6TROAlxrBU
rrHXLjJ+SMJYCIZRLo9M+jx5FsLFkVBwJf6RBsO1sJfA0m/Qm9CpPBFOs5y0OxKGM07/Gu+u8Yop
oO7KpdNnhMfU8C5k9ZwZyuvhL6LqoKfmF6c5sJIgJz5f4ak3O/14EFjo9TqB3MCgeWY+ivZS9XTn
pLvGoLsGxI1QjPLffNWTLHDYf44v3pWUt0+eSukg8axSXV1YYhRrIgGLx6RPeGJVvksMVo6F7Y7l
uLN2w2yGhMq2KBkwbS2nZB0dtSs5xQrIfqgu0CazwUFJTTzM40Fq03PyZijBx6QxpiiGc3b5ZBCq
VbEgeO0nx/SOoTKxvnMLXV9YXIocBLcZbs137eqQV5PrpUh11VbU/EcQkjihW/4lPOXhpJIeOaFi
bPrl9wJa/vhNUtWIFro3y8HVQLTMAvLV7qm5SwLFzIBZHf1U5tbCqVCFNAdqKO679ffob5v8ta68
vfRbIx2K4mdjWD6aXNqPXUdSSvvsIT3cWVTTIQR0glmyC39JVaHq2oXJkfWwf8/vCDxWZjuFlZmi
Lba68sULZsMGTr4wqOF6RhqqWbGwD5KfhBq4dNUwRQdHKgQuo+9lVRK9oxmtBaPyTanLWYWQjFBH
sFFzpz3JpiCMjRn0RP9VRrTnGCe3KFmokgqRlJ615tjKWLoVf1XXabU4EfdN4zIZTnq3Z3ntQo21
gZL6UXLoQR1r+JfUY72BKJajFjIXFCFBBIl4rAkHhu2nv3hZ0k0Up4DwfDRH3eNA/6771lzrxmUI
pNDB5AN4OjCABxSfn/XKudyM4aN6QEU56UrmK/N4Hp7KJViUGVLKv9QNRKYp0D+yKxPjGDgFNvbn
eL5bfacSHl/EnRVcd+tFlC2Jw/ks6SgXAgeIO4WhH4rVU6ws5nx7YE739ZKcdtIftK/QYZO8n5Yv
UWhJFl6clvBDD4Ol33nV6mqAP4AgO5Sy5q2bdPTxJBoxyWlw8eVDCKagOm0aDbulk+fnr9XrkytA
e5gmsvnb7ENViuEJTfgHDEbane06nSUt2bvelVfKqPYu+J8WiA801k+Es3eM0yIEQWFPjIagCUa7
/qyXP3mUWGrXQIBEyWP+se2CZu5azj+JpNLBR9Ar0Lhcg2ez4iRFdKW/Olp1iOOLsZbTebeq/Bvq
oRPMIVQ8O2H23nZi0OwoitV53RPoBHjhDgmAwV2BlbF2n0PNAgal9/Hs5bmxcg6N/wYhn01DnHe/
1A//3z5qwQ+RbU3pEhMZu6Gkg2BYvan4PiVDuuDmEw4+zCKvjCNdUk/JkXlPfIVGZHGNzp2ciwyn
qzd6YqAgC4Nt70+XTeUTY7O+NvO9mh0X2kDP2biSrWAOeHb1SMis8rHp4xhpjlmEZv/yaQzJqrVx
1hMNkhwUTC55j8wiFqbvKcTr4Dml8oUnqE9hgtLyfLQY0DzCVzlODvsRHEX7WEwQiXhvvkkRfM/u
y88kUpW6ooyzrpuyDPzICKpkWMjvoybhaDwR3Dfb48q0ucP/NnZIxkN23uW0cV5RCXIFmjvdqViX
00NvGZtCKSJGpTBEf7RyxmZqgcLPSgT94Nj3ee35aWAGntac3aXyGsFjqHSkITNLjQOmcjqjSVpf
vouvPRf2x03XqYT3Jg2MxciiKzoKWm6TbeIZjt0flSbsrHg9B4MhZojypzzX7MY3/Fo7uw5xhpqi
+v9OumbrnxD7A3Z+QhMPvrztjsvPgZtwnHU7R/IRK+yTfK6ERGRtvIXT459iCEV4yAG64k0ijLEg
KxPt7wxib4ouBTcUr0QfiFCX9EPNH49nY86YF96pgaYIHTq+AMzPrE9KF5fgb9Dn1DUj/B48EuLJ
9jehJcgfNncpL5ELIzuNMtkffxUgtp98AbVp5bEdUHvSKSuUuxgFghcGGfROI1EXG7re8VEQRP5k
49j0FtRY+L7dygrg/04ZTSyxeNAORCypzimfeedPfHdG6pR7A9MtQxLaX5JWPR5D6Hw93L5fq24Q
BW7Hmy9R9Tgk0FHgd7BkRR0awM55T+Kevw/+lde6Dftm6BwllQN9VaW9CXnk4qnsxkoFYLChJx9m
LrifYyR8i0+vmqNQF4KVZK3MUKwypStmTGQ8cq02zxY7I8iQyozhaFUR2Os8FWNHyO7BKhX9AE0W
+rVwf6iPpTzgnHSwuKjVGK5eLzSkeAk9H0IVPqOIZcKg+e9RdMndv3nUJJbM0NWR+RWqWIFJj4JY
ntaZVcGAQ+eWqO1GVxqLTbIixPAtw16DzDBtmgln6OEfziEU0pkGppKfnJjgMRZK43erLvqe1KJv
7jj9OFKb8JKtAJiYKvRSRjvOW9CYohXrGcBJSOGX/wZoYp633GR5QlOEtSQTGKpke9cIVicTCuNC
iU2wrlaYX3kLk+e7SNt+04u/AGej6vqIjuM41URZrs3C5VQnvnQbgAYCVveAgIykG7ddGdhsCoGQ
FoajYbkUbLFR1bzw44JN4XDmhUXe7C/q5Cb4OaKJC7hjD649peHSfA4sx0S+XYAmv7diwOgReJp+
uqz/wBsZkFw3vqyQGD5TWctKwl+uDC7kg1Xz6A9ZrOZl8HCqIPt9GWjY1xOBEMVhvUuSvJTTYy18
1pk3DCeU06ZDA6UeT2pguMR2+EoFK330Guppnu94V2RPv+wXJI1fAQSU3bZK4E0ziDNLDZO6PEkq
5oIQJ0o/pDjwHA6t7/JwRw8LRZakx3kzIqINZtzCv+srCVlocO+W2hh3qYzZ8e5/8uq2To7zSaQY
qVxHqW18mnXTBXcyhiyuodmJFAON3gBNab5/1Y8lfm82s/SjFYcvr8+GtvrIaMXKf/SFuuYBl+Q3
kxu1dCNhAGQb/3xWeZG2K6FR2CBAUy4Yzn77m/irWTsKoRuws+PF++jdAkv9hb81mPbgF1y0wmaR
eQE9GLJ7iZeF3BJphlY22YIUJu1OWIGpiVdj8ThJ+LeoAHVydi87qIoMjhpGb2qYSkIuA1JnqHWk
ZrGr7FrwWQQH3o9c6kQMb2riU+7AsrRE3vxoTz8sJmTRX69P/63Aw7t06xtH01nhPKnSBx3C+IAP
VkKgWDh/HyqLb95+f4nEa/CRoYAFxWjAt6qcUjt0xRCDcYIylMfr0z9wpgVqDYPInIqwaV4FouwG
ydYxeK6+4ZB9K4HFfeAKF9kVPUnj7dHobdaTrL0cBT770TDtjXjWJHsUz03zGIQt+60E7lkXbklj
ZBCbysM2GidvPc6GHFQkpMEKCz3s4W3NxdcEjd2SpM6HK3/AVYCSejILw/QZykJyLkDPdiVUrAXe
DQ/xyVh3SbstVUrn3p7Td3nY/Oq8CaIBxZw6csRYrAWzRjPXjXI3MZ7QP0nnJiyR1OkaAYUb8SSH
g/2Z1kvEo+oPVGwp2XRxz/pjByomPYeM8uocC0kPpdAs+FNRxEHljQ7RI0spk7ilEfbwwIJXlTrb
2cop093xzNq0rsuwVTnVzi6Suj4UFC00BKtbErepde8wEaBN3ItOrImPcnSMj4RsvTGOU45QqZZb
VZqjiacTaCEuII96N82Ecbd/H0DCtxdtcbiJRe3d8dlZR96A9eY07xF+m46j8s8GjOf5HBnZXkYy
uPV64AZpFMzQOoH5ACXyk5XAN/XeZjdAGw8l/kbr/tzNhjS3KWyKyr2mOJUlx+k8+cfq1jY9iZVE
vV0vdqRNJOBGrr6VXOuf9inUAkSm3r17Z51dt6XtufM2sa+SR4aZmmo/iI/5IwV84zb4CfON156I
MqIme5klGSh7N6FqMPEjjPvP6a+0KK6lgDlzXgXksV7vP7M8SQHqRVccuhkde9hTWMorxacZiWgO
8NaRoohzQVDdCiGMg0L8ObRDguEX7SD0aCBn9mmopqH7cPPOu2os/fvSu1YIZ7byJ9Ue26aPHhJw
4iOfGWynS7v/2FJnd3Bq448p4y8d9e8zole4qzfm0hv8jsEe1aJP2OMkRvWq9Uw9KIbthvmDw1nY
cQ4zPR7X6qBDD44Woclo4jgvBRRnSejI/5DIRzamMRnAwWWolcS5qJwbSgbTczf5x0uQOa/ay5g2
0gK6KCWVX+xi0yu1JOrli0MgyfbNo36jvBfGU1bhEA767myg8QiUUJyjgwS/LXBzX5V5jLS8c95m
iys+mC4MrtFaBhoNE6CwbryVHGIVI01cbGuycvGZZM/vElN/rKTa13ACJIcsYE9F428phsaux40x
bPDLc8Xgoq8sJNzzIBRxMJV50OjtKpz50ZGkGPimMQ4S7IY/vfzRIdPCKDKTpi8+iQ9WNmYHpblH
3ymlVola5fu+RU6mKrlcGbqSK/PgZds9u4MvMWiKBHUDVkwhRLF6bMRY3cYeI27YEhQuX3Tdwdts
M0qeZB+EP6fQe4pgIfhisH2NIvHwyVzWzGhL1/iSBYbqod7gVUbqhMiEgsovr0jQHmAYnsmEgfXm
P58BYUmHbsGl3GH8zXq6yqr/TeLg+4f1Tz5vcvaju6z2lB9fbSVAeukT0nGeo6Y2U1iHhB/gN4VZ
7Ejf9e0EqzbYeo8LBHzF3gkebMbgvsFmiDZlsiTuOxBo7wp+2WWesjC/OzRWPRpn3fixxEyPHItv
Lbu32ddMVTlnzA+ND77oATK9MxVtMLl0+XhLCvdJYQfUq8XSx6pC1Q1zLF0PLrzNRD9/b+mCsbuj
EOLuTbKhhgw67gaHcZtamaStqrZFcQj9YtGWlQ+EXbf/dMUZ35pQhSeyoBCV4A8gO2dKyer12xSE
DJekReB0KKTgsx9j9wnlzg+XGOPgB5B3QJcl03KMLZLlm+nDQQXFi4uBA3U9n8V6HK3cqvOCs8gE
fJ2KcQhkOd4tZozVf/spes/FW68ScGjJCWErGvqHjVoS98ES5YDwljXzxg0UKqFVEVqip+/C+FTg
OxHf78QZtXA1WVi8mVFD4T/voG31qq+oZ2lfR0i/pkaF8wcjxohsxV3Y2PoDS1rfM6g0PjbaLBZ6
o9U0URgNOCfI+3PWRN7agfJjW1j5pKQM4P1gss0Ib4e4Ayv7wA6XeKKh7GoDvUXcvUq/0PnJknXd
bSX74kval1C5EcAp6438vq2irrKJ0g7zBhjNSYJcYNMp2gVyRuos+OFTjRqUYbBi/tHX37klR8Yk
4AbIAEF0n6QDlaHol0aJNj6GT5WykwtohFk5TnYn/iIDzVN9TYsLu5z7NZZO3o/eI4gKJYlLjXLz
XP0fjcqs/abIFbuehoNF5N2QYWoojQbw1lkxliGz3CBW09pzio2ssfOJd/IYhRuOsHa49fISuoiB
np5I7AUjPvfd9vkWkUsmNBHachAada0EHPlM5UVbQdW+1pJWJtIBCr1ba5B2+RfSF2xP9Hl2cBDM
b90NbTERq+EmepKGERXyTUafA0yNN9GF2i+D7sL97lNexwufQd8s1tve+pVlmkQgtpTiwLmMp+dp
9zih1rUg6nyqaF/wrEqG1O8TX0HK/Y9NqWmQeB8SivAePkfMu835S8O2foIKvufPRN0MPPe9KGrR
Vl5extORwSLJgpEY6bz9Et/R7k0hiepJvQIDt4I2uHKuOLKftbWjAJJjcCXG8r0mQPJIaQCuQzUi
AATsqOweUvofCdChV19vTlpXoE5W1Ks6CwQQyC3Xpbyfat5dAZRkDwQcUHcOX432z7R7ErBp0qFx
SbBTo4BScu7ss5+EsKhLPXSQXHm5rH2eE2MMZ3SHlOTwaeNnKIRO1tlaD8U6YCPW7gVEx2g8Qm20
/E5dk1j6XdUfpg6lNW5CikdTHs6WZzK/0hyEq2+74aJlrczR/8xcAles06tVt3QQqBxDRUYeGUix
ySSFqrrD1n5ibH8QeJG3oH1dtRe8Jz7eHXtyxHBuhIjzkYe+kh9vnMLDQ0ubCqdjRFWHHpLlNOTp
YutX/+R46ejdi1G3p2pqpoIH+nLTMipBC16Y8V98MCihNiJlSa/kJ69hvdGfa9BfFjgj59IgphhI
rx8/lvDNUA/ZLpbQ6UxBzAMAxq/p/lafflPA9J5xH9hp2SmEgggNQl8/ezNN2ZpfEG2gD5pgPdZg
g6JwWOypYcFnTrBKnTcPBTo82jTuAD2G2uTkzl36UCdhSEzwdlRN2/KRD9h4qYr6BhsGSLMGGUEy
ovWsSSrkOG2HD6g0j7RwaeQT9aQH2BtA+vVfsFtUUp39+cbmGpPdriVu9wYETsC3EST8AAsPbTX3
/rLcwCHMLfqc7CIYTD+mUFM0fN1HCLzaJncKKNTlWhw8jCc4ZRh4t9slrohJ0shTnHjnd3KaPIJC
cqyXtt9nXanmWEmBt2F2qgwdzF2qx+Ujo4JKtNvuP9UXaGF0P/6PEOAWR2mUUmYdzLA6j4XzPQSz
STaz3ECXROHcKRHI0kv3a+j0Mu+1G3whyDN+N13ZD/Yr5Ja0MEjouePPNf2pM0/+EHzBSroML4Iu
0lV+QyVAAZqa8lyEAe28VZRENg4OYr6/yTaPbM4eprdIv+c9LFswwyHqrzg10YABO74AWXAbQZx1
/JCo+OGyCalIdNg6pBGJTqrSxjpNxTo1nlY3sD2edNDw7DvbUbNDqmo+Xu1emt+rt1uHgpK7QTX7
FW+GlUQIpLu0R7uUD72EL2/Ki+aYOEBE3bl5aGU3U+gmLAm3pxeLRJKtV5urxPQFLg8dNgiUVPNy
1dkgkCKmVVrhOTd+NDODPf0ufzh61vr31hZRM1VfkNxJn/9QpOsUD8+R5J8lfPQwttolbiCfajIq
q/F4e62VpWBeKlfxCLBa+WBTNPKX1ag/iPaJAJLEgNqnhSbtq5TsRD7d9eXgzR3hgdlP7rxuaMCN
2qEHjep/gr1MS3X4X6IfjV4a5L0jEohhFpgB0Wh0wGP0hMPaZlJRQACe91Pz6EITmksVWz9S1bf8
VXvBxQe775U+4ZOn+tcmtvQ+RqGBxeIHkSeAU0Ii4QVbt4pC/gxgJw53VH2DdeiqJp4QYAC8z3ye
J0ipbtARKihWJIdY4MFs30HkqhHNB1jnd5hmIVC9atO57yolchLCqwmcnU9ZKB2SLSE91m9+fymA
Z1q7QERtMuP4gL7mr5LXcScVY6fAMcBg1XLxHbGu7I7CelCSadVTkY1Bb5rz89YUr+3wlYcNKbwf
AVdfkXRTlYcWu+6L3IHQ8VqJwgO/8oT2n/Eto1/v9+E57/FcYzshAFFJqaOOrEzxtUnrH6+l75/S
8iD8jlTpxI9QdbVsh2gd4+iN/wGw0eMIXw75X8FmKDa09ANWYCOvQLvIsaTvwsvF9Spz0YY+78tW
rHbE37K3GlQFGTfAK8xmDcHb24j8j/hSdce/AzHtxdrEzBko1Y2UpbKzg7C9NVWZRTd5yEP0hS35
6TXvohmrcOioKxVHb/Ilqr7DYRym/T631StoVzWJrHF/gcIqGbs/cCtZkAt0/Mr5CVULE3IzPixv
fy3QlPDEhodUD0gx5/TUL9B0R1q9Vmdm513P8CclBKybR/W3Y+ZR2Bydxk8DLvFmrJHiZElUGpap
l6cmfqZXwhRwjdPMcMO/TYBVphAqwXnDHTA0fNeNWMfd1XPvnqPvL0XEeq4FmE8VDvsM0IgTZcPA
BwipszoHABcuJbTOsToKUZkktfcxdrBedtx3gkHt/eRH3Z/BnuF9ZeFppzCm+2A8tWP2FgWi+PG1
Hwrg1nmINkaMZ0wgfRZgKl8xWeXnxY8ErF2S95XgM5pl58kgJXQ5cykkieHWCjsDMHLjNHMQ3iMz
vqgo8y4FhuA3Krs9x8oPilyDrsMqF/JSAGjJc3lT5pm88Amnagm6KF5ziw1nx7aFpb+chL373UPM
5OnRcRgclzSGhxFq8IpJFTP/VldRl0RarlAiNdzBo2PgwqeLK+TonkbUmj0f71li0f+tPuYQDchQ
h5tKpdILp/ambgQcsmAJku3zOT4qU28M6zSPU/FvWvwNgP0GhVETaVz1Bo+LgbW1YNcEBJ4ZdXlT
zFqxGB/WzbhI4gfevtNcpPTdr/DRCrszdqIOHC1eU0jtLQUzlnxALHwPOXd2NJ5Lcymp1EJ6UHeK
VU09wW9pS3/xBzetxo789dJYY01LM0JlR/kyabZupBdYY9Zv+rB10fII06UWEoS/kN/GOoRN0M4T
/lBWZoM0zJLsPMfuDcO11kWCTQ+9UzDGii5FhbUnKwjGz6x2LdrEZoRudVbU8seDuq5l2eyir1mR
iFvf3tmCPUIJ+UO81WHJTrLpxbck9y2oer9U4Q6F9j37J5fkFZ1Sn3u2WRYrl8lJSBO5CyCk4cok
dxO0k18hf8eqxFSaWvH+MAyEFBYqHl50FNDylIJl4NdZ+Gfl4tAV9VXuyP2KVTylA1WvJ9Y2Kwf5
E3c45F4pZUmNLTC/D7WgPOOrNJrhnfrYkh+qtltHUTh0VmpwNngHYFubvG7mfb2vZPyyArB4uMhb
lUt0q9J+6hyMOrxW/5rQwHMBZj+9dBPWKAhpSLTdz1yT26dZPovxx1ZE7uHOUse6yqapWHw/vnVR
SPJ6hjLjECuuq0Q7PVvW/mgeRXZ09ZAuYCTdLcVF84dCqb42sqUZIC9A+kkrsf3CPTk7R2EsYynA
JrWaBMbs9SbXLuh7433JYbZ6r7sPb5X85L9bMEMUnaEAjbWl7MwKwVlh5jtfcHreCGgfDqlewQj9
L0OtJolXLwKc2aXWVApW0mL5XNNIZKQYj4CjpatT4N4BtXorq8MHNbw3UbZq9A04LdMsd1NkUdNd
GVDfVWi5fluprSr23610AIprKFfTldNbnRXKnqeRaZhdHxslZFg43cp9tRB9+TrEFYlRGwa6kmDE
QNJSo2Ac0HokdUfmMNcGCv8kJvKm6+cptRVeqxwOllcM8rNHa9iQhcLmtS4Gu/MDa5JP7QZBYnbW
rT4wQqTcVjHWzRnhiAi0gJyPUkUePoi+nUOEhRNho8klWZnVFHMcvLZasTfcpZv8pqpcwaUSOlnB
2sm/jUqoMRtJlyQm5fCLK19+VakbSLuwb8FKvqXFYZaczHwt+j/ePT+FGExepaNLR/LwDV2cVRP6
IgBkVHoLj6MFIHp1wZmdhTayWPlv20m9+HQDjJAE4kmwsTB14T24VbUbpmjSkXcVcjLj86++47gr
qO8OWlTyl3qt4myJUZUMOAA7qEFzJQ3X9dargcf1/OWouTmVb4WD9oXPWsciKUI5tQZ9pj+Qinqd
+hd0ZNaQ1XdhMOM4vaKLOmj97rr5paXMloxnsLogr/TcnLMAsaC4RUoVGM/926WHW8VjI8smymet
EfoYsgxFbaQmqub1JfSy13qlId63DVtRQbQjyUJ15gvbT7Xk4q/rumTh/606FCDgCPS6v25uEKY7
lRjta7Y86fpSpJzodlsDGxJwOCr7YcEsWPun50V1ttme8sJzc1zxhTnuqKeGAQvX9sPyuYLQMUt7
hSPjrAK3ru0y2NA3Lljh1nHMS/mBAiPwncQSkSJLFZrQPtC8s8KP4dqD3S42n2pkcCkolcTWtPc8
VqE3mmc8AdCOLli1IQyw1Z6WsA1uDbd0gJLp8tNi8Z4L46kHczY/7+0Ia6+CqWilUC3EhG5ZHZrR
I6uYRYRw8wvBFx4mzgzaVIXdS1xxu60dsTes2e/Kaz8sO3Cr48oiRbzNHiTH2rcWn+qgRKcCaf8a
CeNSed3tTgHiUCPN8w31dYefeefao9SOZ6rWnXmY/RJGXtetR3MdK7KLNUilYg9TuPH5dQm+I9zF
uuzDuMqXIZsyPBzjkF0xq9b/CFehtRjsa1CXmimdlLXoeTazJVEPzSgo0qooYJlKgxYz3Ympq8/o
2QkS4PgtMyGKyjA8d0qgCg+YZTwb3BKx40Fs2lLYvPMNueYRaaRhOCkJ9NPUyOH4yhprHTj8TMws
1caWVZx7qycEndsMaSm75nTVYPz3pnStgCELxUSFoE7FM3Y55tQAQUrwht4LuauEuMJla2BVOSVY
ybL5W3jsV7atbGCKxE/0Da0mVNuwTYdu4GkaLU36LGPkSJIu0US3OiTLO672xK4bJdjECw1aW6WI
dWmEVY9aBtqzjI8cLVaXQD9zLI2Ux+eXGJ8OvzBkhHLyq1boK/0XCHyWTlosCdXj7lbXKGLWaDET
L9LUwvjSt0RXTmWY8y0IjLwNaRo5WwmCuquAvR6bdN1IudD0FoWzODUsKWzVv9NQbSUnVBhiqMLU
iorr/Jgse3ld8FkKYO5F1AN/XeiTivu6e3CQmrwDBeyw1RXkeVMdbgak0GxBz/swq8MIjS4wAsDt
iQvhLwU06QH+r6ab3JP5CGLLcDI0FRlh3ZM1FLsngjKw+WMpNQdNpAdOcFgSCs+tB76bxH5eOQw+
no8qzdgtxsw9fWLatK5m25VsO7JdLEvicvm3wwOT4GMUNLFO7kk17JikTM3LHtT5FzZa7k7u5t2m
lqmtBN3d0cpzh9fh0o2xmFZ6TofQBl62gJ8as7zJvD730wBNWbAV7aTcY0kCFMkAYzLzmsYrusKf
NX/y1zI4bihNWcCNoGEURxWLcXabUR9oJnAB+dBISe9JpyBbhHjwpzXGzzNqqOB6IuWDPCvgcQqo
LwW8W2VgTjC/QrCDiRU4XJyWvrt6ltMVS6oomMlE7ZVuYd/xg8gICMA1WxZE0LO7RpabWr1VEm99
r2g/D9n5CEzUqvlT6lOJ9tQ+hLhCn/yusHPb4jOCzQnwANUeCXYeAR5laemjHkF7m4iwnL7jhwMO
RptDqv3H6LiIIPRtNVfTxNsb4tqvtBnGZzXEI9BSvRqY0Jgf8QeVpz2/hFcvKuYyNoT4uDpL8XuV
CRkfioC4aClkNRjWkMwqgM33JZcLWJIaJLBp0Ivi6Y/zuQdeZke181H3418b+osSDpI6ToGeOMXq
vAJ3iPgxk2VgxrHLM7MD57zYJtMHn8Oh9+63ssDglv0uaEuapvIuBc6zY70AFvupEYbut7dNQ9fh
IYuMQc6JbuGg1H5lCp/eSFh08M63S8fIkSxB5UK5OFcogIkrPQHkIIUoiT90k8uqDt0cALqzxgww
Jn2CfxEf8xdhlqU9rBZth4v+zwZLYKWYff2HsvOqYRld+R/ihkA1Xo41Tek1bGmLeRo+dQ4SfGpc
MIJ4JrizcADflzKaHo56ekwfNqcHzaz0mNWJgiWgBCjFIYiIH3Bg4rx46uGf/POVLp1Irn3Ql9+j
plYAcvYlDdktSkchAVxdXAn6lKuEww1x+yWECfxy2O59JmKhD53t3nzhc2wQAmk4g44G9N9jZ884
EJqLun3loIlfucZ12Ry8E37TCKW3ZqO3MIvZ8g/IcnzCpCVU8UK5ysEgkz3aE0p55TD1ZdpumWmj
ad1pxvLaJ9teAYdCr4B7POLmYJdpwwPzgi5j8itEARTME96kUquKbD0dGt95c5Zf1FXt/4G0qJDI
NszmQPFjNLdLgkKCIJCsw3xtxMGSpiR/lkAQJhNmVQkrI/VooGPj84rYkFVHr8HqA/Yo3ehIj4Os
7yxN8pZ46Cxox9hgbY8+WtEoax+omxalYw2NTMGV9t9QJWmH+8PTfnIJsuuvic+r+mZ0gPkrGofM
fA7xIsWj6amjlr6Y0BCDDzUQjpoKjnBttctQg8jC69S+r4Esa65H62PHxE3Mn502IqShqk+xpNip
AfJw4ODgjomHyzi5ATFIM918d6AZ0VjCZqM1yeb0fwZ2SkHqoJFrMOFvs4GkBc3DTgSGQ0QQmR7n
y7dG/9VSadbwhi14KUs/aWHYm2X3oX3JBjgnHx+JtSk8nEWceVNuA7Fis6VlxV2CaEqYPixQ22lu
AVoDjUgpMpkqzPP8Dg1jVdqak+R4teFqjO8iUiBSZOPXjQWHWJKDptm4NyhJ41N7P8ux2g28jXo5
Px3lbz0tq7dQR/rYgJM51+qUfVLfvt1GMSofKUFCp6Re0yE9yJ/loTyj9uOeXRehH3qL4oAneXF7
+9GwVmiR2CO/OQDhz/Jh8mt/VnI1JDaeNIWjzA2f/ERl0VScoj2aNBtYcRZHHXMk8/C4bu3hvOav
N4z5+VklDc/H04nSy/fTQcLz3ZtogcpwIJU8HsIp/8StKHq2AUMJiZcdkwILEdTBoCV9DgXtfwcj
g4ZE/KN8dm6wrwXpRXrS97knP3Iew+K0sPrP5Hgn2+4UgBoToRSzEk+o2r8YjalU757jJRhFSaJg
rIW0zNswu5o0Ke+G+a3EpVDJRX8GyHIuP/DiA2Mf4+2o01do8NLqysFGLAI/lRqOEu3N6+pB43lP
ow3GE+rHthpzfy5lv0WiY9Z+5ZQ2icQbFPsWRNCwWqrZia5Fy7+iw2/BmBsU/FYsoMPIxNksG+AF
G0ZD7zuIHkVn0vWBYNB3oaHnhQGAxvb4PQpdue+vg3Q87peYm9jMrNiQG1UqAmJnPQjuffl/Yppk
QNV2JrcA5GjWLQiyQ0j9ZmERSqWKMpvxyfIKNj+AO0T+J1+TCozui5ncC/YDwUBtNe3UgD7vWb/7
+YUdpF7VNg/rdv5+1OvYiKamORC486aCF0++5d3UuvWLyd5b1MLykqYFoEJSG8P5GpRqCG4EiLip
6MLdW70cExhgxpi8rlW1+xUagcT8dhREXvQf4TS5SeFcdknwA+v+cTm5nwxiFvET5FeUroFan/yI
/d+ZxQhav9GlTlSGaV7A0CrUWRxIzu6UE6Bgvls8SAj2CBYFe4RoTrCPoGFHpMm7vFDllUxiRH9l
Whs2xFa7wUzAL43uaJVziR3GCM4JV/x4ie1JPacia+Gm7M8jxK+os9/ypyyLIcy5h3Lnkup1NWPJ
sW1Sznu1IWSpux+Mx93r6wUMzv5b9Qth4QdyFDx1ZExZd3ftIEO+9qpHF83pIn8/UVnjgr23u05f
3o1PPEFqbHQlEuOb1IIvuIOEYQrgIDjN+o/9sxtS0i5u9SRD6se+8Iz3NIZJQb/ENnCzGS+P1Q7l
7BZU0ajFKQxxw6Jf8tyDwSm93VVWC9xVYbunojWsVd7ZTcyviW5+CncgzFi+nFJTFU0sX7d7Hdx2
9uWWBhb7lulcd3dV+69GWytHsoJ2AMTRwEh3SQ9bZF/4XYQa1Jgj05S+T5pm9CpACCapuDCTBMu1
SFlOfgoIXATfUhgewt96+wlLC9AZu0b6w65z8oJkjt70p4JztZ3CRKvv2jb31tQUXN1Mo8xh+RFR
xZSCVj6rIoMx3B8RiueGS2xSjIR0IDcdpDnisjMcbT4ushH+Z6cLeQ7K9F/MMFMkkg4JXSMjajpU
3jmaO9YJ+uDpV4aE72sl0ZMLOp9ua5idfvXmSSoFuJAbzJnU2yoXhLJbYui5jS88poIE2blctfF/
zVKZjI4kAptW5jkWqHCI77P6n6wXtwxQo8HkBs6G9DQajmv35UV8DMWSzvtr57uNbqJXyFISERGz
KTTW80mu1OI3FPMfcXz/eaLFhNd1cxOJ6XCiKPuUsRZOLUN9YLflrzzcBbps1CORNqzh4e8S8AwI
DWOE6AbA0raN/vrJhU+wJhkwS5E7J5qGGhBw0IOUdPAbSkyaA0II+kJ9E/85tp7f6emWwAhWXIH8
8MRl4hTYk3HXI/viTqBjIzoVWv0hwwVZ41ZHkogHVbDhQz/LLTpNfwbrvzyLU/GLC46hfnVKX4pZ
rSjPSn6qrT2LBHm5vD6Cd+T5/qXk3dQjgRUQ9efe8EQnpSBOOK9M/wKl2VmFX6rHlNVE4IPIUxtq
MnUOvMR3jXFUg9hD7snGp29B3vkpUfloB0u+sUAh9hZXTJHrjgCZVCRY1wCDniOGQ6yBAvudFqXB
ARbvdpF19miZm+QioxeY/YQsnZgjH3oRyY+ZEEnTDADygRYIXEvII49+moiYmNFL7fbAKSDMXVWd
UYd61V2uAOD7ML+sHfnoA3V13q++5mWoV5rrnL1QpyznPzv1vck9zN8a3M0pTAS8CIv2TohB7l5o
hqfHYmZA8RODzynihTyXG1sifv+Xc9Y+6zwblu6lMxiKPQNqJB+KXkwSno9bGPN4r926R6xqSaqD
qNJ/8Hx/rToZeY0IRE2ZsXNItfDP52IYPPrOUB6xSv//K03PfND6uYeSJT43S54QiHzD6EN/B7/1
ySMTwTDyoILN33FyqFncFSO02k/VDBSmr2VmCu8bj7xwv7DJ4obuoTFiXA23O9P0UqDvcmkTSLWd
PBN1L0a03TZE+aBGMOyRNdjVCShe+n26I38ieCiYos5FA6DRAJ64rTZ9iaX/kksBmbiAu1Iwc/Xu
5iXWKZBJR54liENepbb1xv4OtEqrEX3hMUCY/Sioe2Cmmf9fNVq5HzQFCEKVNWv19ajZtgQkkiZA
h/acxYNSKhyaIZ9GISoQZs3W8A7WeaUc1PlgwT85+npHlsWb26V5XuVw55OBXFFB67iAyyZ/mhBY
VQmj+17ghbYwZiHMCHY9XAe5Xk/UVDLysH92FVdVELsYpqcQTy8rZ8TKxN3nxPhndfiyRio5Kz3t
AolWB/o87vPFU/xWM64QnBA+FZhdJ8NkWmQc3GbslTV15BdDs2zJCiKf0ATgEMgXaFKCAtLMGN0Z
vBIbUKzM8N1rCH+OcTr6W32A8uZztRJ+ZlSKRKharIBQKxGcSXtrTtWDIfGUajVgiGRlvCxa+fK9
KKV5/y37d5nAIEnH55wH5JsLyn7vjhsKv5PW9+3weaDD+RPLDjRE62diZdY6zYwpBa0Y9af+m/pX
pC0oNIidhsm2EP2Gxu9xToK+wZWxNp5DzLPyJqr7UaXl6teU5sVy0k1tGLLi6z01C5fTk5FW19o3
wf8sr+Y37brn5+nySlcPc+9rORSty1sZkwNH/13+FyWG21VXrk1JM2YMmISU9ZDJ6MJn+udpTbr8
AHRIR0n7aAarFIBePzVKCVRpqYzz9YpsRlhMxA7puME2OoKCbJmWUHdzMAItjCew2ouuBjXJBYUS
HV2zcV6zNPovXy24tRKW6OVWD+f12VrzKbCiA+2NrgBtYLM68K7Z9xGqpLxUsEq9XQRIi6JiBPKZ
tD3CKZ6HBiLfU2Qut5e7n7tF8VF3MU62l4rHOmjGPJPo3VOz3M+MPZk0RlspqhEc/kgdH0MAy1er
nRXiBQTvo4H9uzjwOTqKxyHWz7odYndTV16WeAtXQ8eTgVUhpprgiCQVGGt6n5pnIF9VOGxXvLg6
8qUBh0Z4lNwxitKakAhAEaVwMx/TSNS6TJcEBXSb2J0K8maZT9rP7Wr8vnIMXMJ5uxpI2z9fgZeH
q8+SxvApzNlS9xMaIJBVuITVp3Ve5NBbA/iStnHX9lkMECSlJE4A1Go+79IWzEHT+h8I+OKWh5rg
SxEng1fpN9/tzN82v8wwxtRRl569gocRE/IBWMnoTuyoQGw4rUMlLL6lHHw+uaFEL2Imc/8BZkJ1
sOp2mIQTTXNHwxZEM+fBVUZtMkvJVw3LQLbeYy01CUIK5hPc384nImHGqWayA8gSlv0KO4Pr7Q4s
B3zZoKRqBAl4CBDM5bzzDmqCMZE4s+0fX5AHoQdpUyMKFwsW/xrX6JbW10Us+t8aSwAL1oNQ0dpd
bkE6aSYP4V7onNJTq3i7NGVmFKQW0m/knTOQp1ias1S+SNhhgTWn0ABWnnmBS5Rf+y3Ai3ohEwK7
9eUOyUnMtTNL9Y+OABxFrREjv1d/XbNR8qRZ9ejPuP14BcTooHBq/+McZlFyfP1RJyCabljYf0rw
iZUkPT6bNnZ/RrzW+irTb7/ZLePMGcDL1+E8bmJqRJlut+8Zh47icqLyEiQMRJUCku9P6FycLNGq
E8uHlcxAweaKBGNnEr4nm0ORfehS+0IvlP17r9nYH0ewQ1JJ+Vih2lrmvIEkIC1gsUtsArS8zWES
XLmoI9kkoU5GAJ4C3ZS0jytcO9ATkNEZyQpRIlQwOnfTtIi6iPGQNJ2eJabC27OYW4vCoI74J9ry
5KYG6a3ddMogU5BSrI3MgLEdewcxl/SdPXsQqzcmXNkl1oCOwTNGGQZs0Rt+x91dB9UzaGuF0b/M
odW8h/PfangXXsRE5yWbf4QRM4jej5hIOBi9OXB9G9yveHyP6AWev79jRPmRbmVoPBkoe/cUc4fp
AiVMIqogeRXYOxESsG2JuLR4YohjIe9LO+hHK79+94jvZwL39JxoVDlkig0PpedL0oS/hFS8cfgE
7ok7E/9GaT04co8B3HG06uMTGhtSOm4RrsF1yUxHc0U2l5MHHnOlIU7Avu/Xq+ja5WPn7cV7Tebv
j9QIabAdC1DOzAQnXg25pTCTiRsTt65sumxgUnRjcU+PqGCu5w9hGMP2Lev8ZnI8ieYja3YmExSt
xHeNlgf8KT1PhRBuJ0sAVA3hBbiI9nB3lhKDmSp3V2pTBD5SJCdYXFc41dyGyR+NHBbmrTLmADj9
jZ7pgYRgw9y3wN2ZjOhT96sZcWeSvE0PYck9mxBqUA3ZpngqSVmiTwZ5C0PZlYxjRnR+ZV5F5Y2k
fXnQDTrEelZqmfxyRv75SqLGz5plrKfmeHX2FNQauncW3PR0dnbj7ytQOg32snmjfPPJ9p+uoDx1
NhXKrS75wwXPUBzfTCNAyXUDT9oEOB2jMKvgtfx1lxCvV1EOhSO7/kCkUK+NBQwJhxjjMmfIPHem
Oiroq+Tkp23UfVpJ4cBJA0ttzBGSv3fWp+x9zpraSRHv/zxxH+gYF3nab0PFv4wpHhFxegfWyjWM
qH3iZRwne81xHo0YPtIrWUY+xzvgg4ter2W65UfLY/vH/7uOm8jXEM6nJZsRRzOT22aJqBX51RHb
iCJkeyNUFGmeGOYUhE31cruI2YY4OoT+MS2B5N6EAS4lWYfq8Kqbj04DOeS1K07RPZ1qsR8zoEi/
2cYUVMXrZjpyBnIVDiHQcwdrK264vYq0p/MwHHWLLO+r5vhU8QUGh35taeCxvcryE88sN0C96ahg
ra6ppUljVhTJxwz5T2DywqQk9VKONwAPo88WsNDoNiabxufmaaWn90xXtl8VhRj94sQqUw2gccLo
QQqiZ2tMZaC0PN8Z6/hAEwPQkoZWRU+KOcaDP8Nk0wFOAB4Y1yhy67/XKm21QN/mJ9Nm0Ov5eYSD
9MMkqRq9sOXrm1UCBA6h+hxEKu+PTYncVH87traRQkZv0WNd71S1zWg+n6rcMRI+bWW1QwjbWunK
Wzh1KV1CIdTczxubu/sxrs2l3F+YmQmkn4P7lvindxcBBlDSXAeWnBGokpRH1qtkkBKU9isNofZe
iizW2igSZtWrI6K6Segc2m+wT7w3+N/MH2HLAwAdfOz8s996h92eRFddZkOXxbub0AlaHW6A+/r9
XReYw+soxWD9flQx2YrvaMJhHAZS9ActcPKiFJ5pPW/482Gme4N+7j+YFq8v9lGW/G050ZgspWJe
mxxZRu3l2j6y+biAG+4JQs66iQDVo2wk+fAaUyMEKpJTnSsMDUKXkH5w4mpKYexMC6Gq1vDqTSU9
0Sa3fgSZxgfUvUv26Bp4D9ZSaOTR/oWP8W8aMYrSYdE3K7DS4yUbxt/1BSNHFHRt7Eo14WcY9MZJ
fa8F+tNYdpUWHPa7xAP8T5ypkqoSniflFgVpshQ2TEpU0QKhIe47VKIDWQa0Qo4bnUk5D4V1I0RH
CNlzI70TpEOev6wJadrQgXZIdrPTZm8lfFOeROU0gcCQKIJ4jv3QtjdlAMZPf2u1PYM+9/WbVhk6
X5yJcewkcjsVVoZnKe6VkRJBvOPQnigaStxw1EXxcWAINyscqL3Kal5KkZW/rT25+1uKehut20Nj
ih6rf+wmoAku0QQg52QUTVlfnnMuKSPSzXaWiGpqMxjyzuMEq0m2MlPF9NLkKXY3h70+YhJ5qfaz
uEfLgRfkjfo21F5hFNMd1UxR88AqgiG5CojXK3hEdy/qpqtgySBjdJV1YhpaG7G+AGCpDxLXH+RD
QBoDGeWyighveFFeCqauT+9/xKW9ZfHLIeOLSujMagCpDU/lxgu1XF2C7+7GQWdz6SJGY4pUBlku
qn+o3x6pQqpBflikdI2A32NtNT78ZfGVQLZVmhqs+JdKic9xKSfMaVxCzCLjRjWjWhRY3vdxpK9A
ROfKtckPbsZAvk/JklEQUr3MVlYIjnM5gojpXpuSOwesR47xfXmY5QvwiJDUxaesIFuTAZ5toMz+
fxk6d52WW+xbxCt5D2at/GjAvnEdlwdUe1J8VgoeNA02Tx5qGPFYjxn42nEx81TqkjI3PuJRbkLW
P1K2LhRLXk1AhzZR25YyYMoyUX0+Wo51G5bbwY6KuS0aa8Pg2FLSCeHsJ9xMoSlAi6Wc6jFwwZ1s
/YdDTm38h0hvBOKN/TLMVM4KfaWIaiCj6WoP3qHUGBGpH+tDrK7KGdDC5nzz+FDTwThrPLARjmIE
noTq6IuaSKrJPHbkK4M133tI03C56Uwsq4RdfDGR60FfufoVXBAsFDDDadPIMg3UQ83wQx0l0JCh
KiRmeXXU+dMUzMMh6pTIiuI11MCkpJ+0ZL18wgh2UCWKm4MUZ9uh0u5I3A9s/yHat6efRwK4hZSG
t3Q7t9sO9ON3D3S+JkV5/6iAcd0jTFI5udyBdGLHTnB/cge5wzD7FiCwntXP4BSp64Hp6hsj3AeK
sOd8t1N2iUB7VVFmP/Jy4giv0O27baexy4dMsZj0JXifQoEm9BZw+BpCWFAvDGlsTPbOdrfsLb8y
K4Mg5lbW7iXaGS5BmyfOCkAZsDoBtxG7pOKwZ+IaJBct6Gq85UwxAxRXf0Fk0kDsKut1dDSTai40
7WrY0zjfbfqJRLtKfK8u2D11iq6FiFMzkLNM5f6jki0F5ac+UB+bIi1WcnPHACbg/BLttgtiU2M6
Un6fDwEJkUwBn/S7Sl1Ezf+rCuSDN2i/JWYjhJZN1kARj9y+2WjXmC6BD8EKtlPG5lmgPJfWZuMi
2rZgL0rAHyyDrpMUKS625T62R6T8PW9YDZTjtksx8kDQkGjEpGuH/wtpyYUXXJBT59DBg8A7n5Cz
wKgkMOpl0dHtKIPL3cRNEcTGhFtLPst/Thxxf1rfmd6lbOSQwOIhGVYJ7u/8SCJROFuvNgv7QFto
CVCb6tPpc8eqgYy+gJ/EuKvjNmLP/bidZq5jjsK2azIlsBjar+easNxHMOBuLrXNqgMBplcuDH6a
0AtzE1Cy0Gac3ZbCDgMKGuxScMrQ1xrTGzIcVepDpLE8bXirrpw/ueR24vKfE60RzEYxbFA7R/1J
pvpHJMbr4W0vhOQgqBdJ5ypi+QU1ySM/rZoqc5pv4tGG8qIveRuRpZR8wuIKVYvQQaSeerbkreHW
q8P6UZG6xKvtfOlgO/9NCH3czo82n7sYS7+1jM7kqkwSNBC/NimNOILw/sLIOMH3OaJjtmo/gYz3
ODdQzkhTljnP2itpe9CIjxa6na7C+geVb+GdUazZu43Gq+wDA5tECtmw6q9wWu3W5HWmAAZ1fenv
0QjgqXcN0ZvQGDscw12y4OuPyvTRk7I1myqtVJrmj9dGGcJLqj00FRcLvtYjIqTetmW18PyyJxcW
KjRlQ9Acp3kNsGoUL5omtocn1Un7+5wrseTwWoBcfs/G/PrnlIbPPK6eWaYC3pdw2m/4nTMMeNrY
QPpcYr+iYrwRy5o9/eyFZ6ZWDjIzxQQJQVg0M0f9y4oNnVUs7b1VIGnHOgDwEL7Fk2Q2aXohMxjo
WNIUnYhQA5XDaTHKWEI5juKw7SOKipwI0FbR55KNKtbIGI0EBfpjm0lV2ZRhH+pPtLvxROPJ6Vy+
H1bcViwnO7+pXXrOiHbF8giLcPz4sTOOD3sipeIs05seOa0NyFmGRzt0AIv9sa1VYJiwdTKngi0Q
f6xiGwif2ro0TqeXN9rQv0jkZdNGoHkAAjOpzcdjntWCythoDisMP0aYmAewKo3UEXy3QBkbP+aw
kagnwS2mf+TpK/0M7Nu7egyAaG3iYS+3oiJVtRrK1PtUVJgkZBYqOJV8LBC4+YeeV7zI/WcWe9bB
kg+mRGoYkVMh4/rOEHXB1u6dyRoycVNTLtpm7QuAPVAF9iWIIqpZMp8CUamKVjb5qIOe3Py7mCsl
yRzdZHa91TLwa2vj+x5q4sRakWhTJhbEYsmsGRIX63n06ycMR4tAtbCVC9D9FvJ3/2ba4ewhVs6x
zXGnIeI48PHI8Jk1aDdGGC1Tp06U4zEcamk6rC0HJ0o2+uHBEO3n/8Wb7szhJZXFQVc8OGapKTET
7z0dcgioNz4qUDxnevhPIGS5ZWz5nqZaoNLnfeMqIpZ+/bn2LMCYoXyCU4cpzi/1qjawD7AqFPjY
8Y67LMQLrDXqNEJAG2b0dyp6M3SN7EcnzSozqgXUL07MqWUE/FthfXcmV/gqVYdqhUlA3GhOHrz9
uqSkBFIUgDvT/JoHDlt9k3oAryEfhCpj
`protect end_protected

