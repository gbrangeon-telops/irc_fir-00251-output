

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DoylSncttFMA3kx042gUfpgfS9f7wYF6CWxJheifm9U5oZE55E7a0/gn13EV1/Vn6tAoLpUpkm/0
hmdlNetDYA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nsjL1A4AfS+U1MlmYTovZuA+LXs5hJP3SunimigW7xSFqc+G1o1qnLbV4BnmOncmqUv9X6mR1dbm
lvuLbnkHJpdv3qype+E/DkwUU+uuHlSP7/5qiYqLK0/kXVQ9CK4RGY/33UuCkCUXhFP+4VquDr0Q
ctFJ3ADjSF9u4KfkLp8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e8PwETDI60MBXnrgCDSTetYRVktLV/+TTSXZzS5MByZtHEX2iao5JK/khM4FDpq/v0uNsNW0rhjn
1dIPd1mlQZEDfzGgZ7rgxmjzboNMUH8CMdtSuB8lFy7Tjd1hDXqhliwc0PhPBGYBs/YEff98J5pB
EaQ7x9e3Dm3lUX43BX76qZ9cgUsaVwP5tX42M7Z1CZ11+5f7kvoiSco/DGzJuhCbDcHoQ2NjrZeO
tRQwYWFDIi7vBls1ETe/q8cjQLCZThAhSFjjijV74aEYat0gpNy4Hxz/UN0rUMO/XCqC2k8lo74U
XZlHepR+ABhyrwVFzKEwcRDXuuh6ogUCrZ1mMA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YvHkp5oDmh1yxPKtyY+bCFF9nl00iIDnF4JnEfzCQKeCjt2Tok2cPb5/9L9T+H/cQ1x5qpJZSOJk
cf36KzabCPbu4/9VIe9vwmzzbE9Ndy2Ov8q4+HYXDGn/u3gDUJZcIYEnVlc3E6se6bxCrEZNyRYc
iuoolgurhXiPk/HMhX4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XZ/Rjfda7p8W+LhE3BcXwsLXrN7RfTJezMmvWQf9ZKb6JJ7gmlPk8WkUFEwjbu79kr2SMWbEP0wO
UouQmHkylGRubs4N/1VfavspwJxzO5pggGGBLKHkmxqVxAWJEQ3Kp5uoaJSKWxqKIRLzeGXsW4p5
F/e0YM5v9fK6K2B07V0FxCP6WuqrungKJmSTj1Ji3gWd+VJATYp+hkh4HPUA/aDTgCzwwIaJ6QWy
QvHMQKHrEHbRztbzfLMH3RPC4Jl5v7PMeYTnCv8UcX2dwujd4zD00VIt1jMD19vjN2WZ7U8Tl83Q
sPvYlUbNQVTnqIBf7mqYAoAlbAFXbg0t5zqPAg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
VvTIbzWWZBdeKFBM+HAhtndaXzB6L7JieMEv++WRkpdVct11BKwLgu0zyYIw0l9n40+RVTebs0M9
mnna5sCZKtBv6EB0V6b7cju0neCd9A3lJcX13oZ5pgJQcEok3nfcg1pGq70sg9v1J+1r1xHjYl2h
OEJT2r8b07iBtoL6Flyd6+h157260iUuljg2NKnVZMl++YTo3No3MbWv5ivJFclBu0S6Gqpuon7x
+HAQpRbocy9QiSCavjGRfhtKM+nfOLWP1l6y0oD6BNwy+sUHuyRolVfaqEvjVX2YAXLJ9AS9stsr
+svTHng0t1VzJT2jm4XcqYpctQjfHfBLoVF/jv7ObAFXa0RwESxNwcEa0zuiit0okbdLJSLlv3tm
viGc81jfNONG2c0dXZ9QlA8ihMcIrPNo+l5zu0DxFTeTjzlrekZHUG0tuYXTZwqJh+8MVQk6Cf+z
+6013K1dUE3Q5ftx+FbJAduU6B/z77Qfr+N0GMIOJfwenRb3/ycVWjiM34ZUe+LWyPl0O/eswull
XwW9SydjLxe1wqenx0fCTD41pZ4qX5r33lNS6GfSKEmJPlS6PagH2IyW2tj0dkRiZWvItDGpSxdT
MGjR5rEGz66Cqcho1ZAtLu4+tnhLrkDcoaHhCmU8tVwyrZ/LDyrnciP6oieMPm3G0+srGVvkbQkT
+5Ru8Sm4i3nw5DkRy+zzW+SrmAPq65m6mrkkYyOQ7DKgyeDHb5liLdbrPeZuR+g/V7hceeL/w2Ku
UTtuhGNjsgPdE6xRJLrHAL2Ic8rM3xdGRUxrG7JzkQJcx2tqpt6kWyskKzee99SeKX+CEClZ2sEO
ynksGQL8tA5MEfXAWTxSZuUW6FZ6QlVEoyFT9c1k4alaT8qr7K9nLQ5CzPHTcMhKZGAZdVQ0wA60
UVQhH+VV4Ok1x0N5tAal5fUZsfc/NML7FmdanfqyMAZUhbA0eieB4izwrX4QaF/xqq6DhNx0RZZn
YlbS2DXCK8SE2i5cKPRAcYyL4Job4HeXNkYtMi6/anvbXdjH0l08Rukz7aD0og9sNtQOgnH7pBhD
/34Vg/t74tTrXM12wbtTk+lb9ToDXEBQ6r/UQqMeaWb79Xnh0C+fw6gGdSrV+fUIa7MW0PdlIMvE
mU/LThKgnYAPo1CGALtLGNytCJTpREcTEWpAp1fwxeIXporUekGXh4v6b+XtmJi4G0QqT5O7SI7W
KWYaSJmoRSdgfgnI++04kJ6Ypt7GsdRK1X1a+cnfLRvtCT5z0J1oOc8xMBS7OfRkJsO5JeRuQNB+
PBVpuVmpQdkADpC28BUvuem5eU/B+1NXtMQgz2HJp4PBUjtvrdJ5NXqKkjR8IMascMWn0tybWXAc
SeJgGG5tMby2DAuFgYYuKD9C01jCKtIVzw1sY3lRMjSqy6229u2EIkfdusfVHfJNnFHBXE4PNJQh
m7j4Mlq+HpxxJ9Y5er7R9wwpVTS+TC3gAT9GpCQsjMGqijRgeXGr0l+zkhaazayoP77mTd/AYtw4
IBAqqa0+fDgE4HDiKDz4uQHwvri3c/ChDtKTPKoMjFaZ74xz50rFaJZey3U4kPhdoCUR7iJqxPhD
DxstN/cvD4TpCnunds+XOK7bt5bjk/3MRmyFRklFgHXXiZwyDjlLdgjpCvihMq7eHLinM98+Ft9j
fUsqOEG6Wy/hGgqWzyx6PrutU3l0dRGxuYI5DUPmdWFKa1d5y+BlAZoEwdvt8xfp4Co0k3qauPPo
xDYpnd4tNj54W7r/jRtNlqIUpLGzsItQY37l/r9fc9OqFcZdQZmcWymCrfSALfmkNO0+sL3Yei/s
ZwA66ZgLCt5NpDGrvWHmH+kgXboOottACWrLdej6nKGn5tVQMqwJH5367VBJQFFKFR5zBW7S6hW8
p1iFQshus2U9ZsD2dWVjiVFMbMbQ9QODI3jZOWLJTi/nEO86TSjxunzFcGEyAKgY8LFxeCaxHcq1
/hyuY8mtlZBSDntd1LUP9C0+57TKBJSJcC0vh+FeOZA7S0skjVZ56+39vMadNZK/9A4kOKcd95RK
T9C3qcAtHPCh0tsw0zdLPJ4zDx570WFiLnqI5rpF1o4vd4tNwIrvEzfDZCaD/KEXBCIcn4dUryWj
MZMySEr6SQL6nFgpuZtr/fLVlvu7wcBi3ou+FcEx75X2bnqUGkU+f9lidpeqAFL04fNkB9mgW1Pg
HsHh9AEZBOqkWoRG0tbA8ReZcaizMgt0uKSXLEzaQ3kLlHexUOP+s8nh+5S8fjvZfpZnGtNEJyf4
BiYyS3wOAy41/IJ8k+eqwOMrraLv3eIl/y2VcfZPcaMDPlLTFJuj/bKWG+hDm8vhQx6gvrtOB3Pp
Ou1saCi9p5e906eO7FP3LtOv7MAW+GVY0+mkrGJ3QiSPMgVTG7F0TuoMs8gCP/q3D7uSE3SvABjw
WXbRRLFADcAtiHburoau6BlOiwo3ewaSuhaopQStnVLq6hotuJA+LYYh+qeMaozorvE7wrgMY2Ua
3vaSoTeJKXyYGPUF54VV+u+aFkl6ZNeVL0JZWy66lU8+042O47e/IkZKl/KzrLq+Oo3FWq3octWd
tHcUlflHJWOXWHbOkIpUQiVpLJWqOaQeJKuGRrMlWK03idecPyN5WkSVY8VVg24smA3mfJnrh7HD
jAeMyTh2t6Q8V7se9JFWrDpT5bKl7rAJxoS1Tk5pkNAoM6/x4VSmpPNuiXoQkUY9BwEdEuy7qcVx
VaLjB5C+E281q7fMiOg5Qoz9O5QQ7zSJfkD2N9EllXiY5EvoFjdTWfuEqwiPxQlGefTWPhBsnqkm
MiuSLpoiMiEgpnAUJAXdTCgxNTR6gCPFiNPU3G9O5V0kgRbORHf4W+4Ib0V/K51veinOjxhzXZVO
MwaKj/qTO5sVzzPBAn9fzMh67x7th111GgwU4ndYVEMN1mCEOkPWKeM5k38Z9Rhp96I5qXdfWXdF
Cz+zVuGMPQhFHCedqOfFv6DhNMTv/m7jGnOjBH0gdfXjTdCTHm+s/Z2mULmQCiwwHn92kxw1jkba
GfdCsh7ZBrEQcCsW/QXoc5d8f2Hrrx03OLxX8OEpvWjjuL3CL8KqZ5Su+cqqAe6i7nl4HLfk89b9
CTaL1zDvAjM+AeoVKEDZLGJr6dazSEXuLLHb9yshZ1EaTaPqANqmkefH/vPws0EalyHDNgs8VAd+
d03Dr0nRjJKF7245+B2ha+V33ZADMMAvna+3RvBOiVuzdmBf/M1anVDMsB8rsGePQ4iRRZg5QCuv
ZD5XMVnJD5HlyLT3Tj5PogJMc9r4jGXmsFH2yBUMfvwtJRO9gRtABwlO7nzdOjtGjgq6x4iKoq0D
Tes77YjQ/jZx8ejs8UAA087gdPNnLc9vIyqeRcfp0gOrC6IJT2T2TWTgk1yBlg5P7bu0thJ39f/7
XflEbYmRYLRND/CqSPxazyU28v1NTMB+d4XZ/KKSDCzB1I6sGIbFcBOYiC/B97hvO5+33vw92gZU
V+aMzYxZflOh2FOn4ldmxr3YhRjndigeMP4hyus28VJGszd1g3Maf9gfMCzbnOJ3IN5+pQTKCEY+
WoDN3tkorZAVW92cJmaT13Jg89fZspUibAygUI7U3EAK5VMiU4DjRNMFvr2RYBKC4JgceCiBhW21
EtbObG44KYPL9wrTEwbqvw+1jXTJcCclQnl/Kx+a/VgoH9j10zxgPVTIfZKhdh/ExIi7FIqjqUph
1FJp6kdpWd/3c1y0e1JJxCn0tsUPKkOXqYQrj75JEF7rNs264iq4pRebOQxd+5T1a+0kJuTzL3vE
lK6m1st6nf3kMjhN3INzN9QlR76n8sSdcVLoEf0jwh1UOfiZzAd8UNX9h6wbHRM0BTA3z1LjD3M4
D4wX3CH7G+TIjl5oIiigX5aJib6INcbDrMwcQERm+9eBGqHMbX3vGhxeqO69RB8t3BUmsSz0TvY3
cWZx6GSlLTr8umJbk1sRMl2fcwXZ4Vo5BEpT3GFAYkLW9qmsSapUmZ0D6SEzW4+PIjA2N+4h8vlj
utIQIRNUJuaoiKKPphMnIHI5Axm2QN1iU2XKXK+gpOzIE7Gm9n3yFCN8n4g7dKRqxAQXeKkbsa0N
Yo7k5ULEj7t36/Sh7DMyqwShyKpWt0RqEs2+CD6sYoMUaUiuTfPe3ZXc8wkIY125wHNaPJ57xVMT
gOdWCeAuLxhz37rYm9VH+lloavGAGD3/KAUs5OvHBveCdA3Id3MVNWChTwHpuWN96lJI0dREImWo
sqZcDD43bIcBRHVCqrH2gNRDiq9MP9wbxij8omixg+SCN+1hM5Wmqp3xZEix41/EcpdZXwp1VrJz
Brjy0oToBHL7xqCw35Nyzz+KfLuZI5AHIHIpkriM4edRxI52dymyJpmHw2jJz64OqfjltIGyWyU2
8Z/TncnouCeP+AWr5MeqbXhaN/or8Sxxb8gRpcCTcK8Q7wTJRTYcSsiQru/3sZ5LXdys8BnZE6/r
L8orhnwk6FgJzVSOjwk/k2eycvfIdMMRN2DgMjvD7C3ZMlXKJzYUYAzcR3fnxHUTWeBCP0D7qIHD
Z417Hjgny/J7voW1R9wXlKNwaU/rQ2Dr7g/fKsJ2/C2iI3SlVpha7BHn0c/CInSiduHvMc1/Kaq1
vB7uB3MCBwmIFUYZN0fRcK3SqzlgHcLcSKdFkpzf4i9pKwhsTML/K4WauooqhVoKpF49OfT0vyYY
jUk+sxI7SB8BBVRWfoL4Rkb3giw3Hww165FO21cSVmhm7cYvFzrr1nLXl/Fmublx09Znnl6Uplw/
DI3Vai7Jft71A8r6XdZnHGFXvB9QyK7OfeZTALFWbVmxJ1p+SVn3OlAmAACn8Qzev+lu/3UkenM1
bDlo8mGgZfzSN1g+1PqgVRx3lianfm7k+bDxi6PIz/6WbqKXVs8uRXSSlN6owVnd9XdpqvT3AMM+
/zHsWLBmtSMH7Ujs8vPStC+3iwegB1yU/0EZloUlVYy61bjDLxmWisnigdG/QKXM6ovUJKUxrwzr
hBkxxMDFgojI8ftBgYRlHB7skIzEY7bhpcyJvZHjhXVmVSgJMsjSlNlEv9z8CLbayyHsK+QaJeoZ
NlmyeUQRhlxSh/XbgKDAcNTELOlrKe9VMHMl1DcE45u8f6UQcXTqelGqHrhGXfhYUbIMBQpQnYNi
UFHvPb6Tqszz/nwQKcd4U/teRvNrSupPGAA8fG6bRNRQgLRU/Cjzr+Tlfs1Ivw2sqNMN7Hry7T6+
ql2f+uk5mclWPjo90DYAH+aaE9mtXmJhrDnmlEA5qSm97rA3CnHo4QcWfUlq780VR9ZdEHIwZPKp
D/+Zk1DM4J4kyAGqXrTDz//o/k0F0BboxTfD5JY30hRxL8UbPuNeLjY+JPSuYkvX+A8yCwOQ2zwk
R+v3VoNwx2As0gZSe/6U3NyEkIE5kt+URskre5Y8a3gJffxp1YJ4L/WNQjJQwj0jufSavY2ZbdJQ
F626ud1ZmLVE2kp1R5+OTwPN9fsOd3PIqPhp8zNNIMqY6tpqJ7VpMnUNpwGIYW7gWKl7vp2ooDe7
wNBfQ6T8P7qyHX6Yr2n4WukNPH41TRSkc/Hz59SJSLfsj4oBaJz+7rABMe81Y8ZrmaW00zKc2af+
3OgCSacYgr8gaBPoIGeS+m1QiLmAzvBkN2icOUXcs64LX9lMyXVGTFUyBN5oSGE4rgSCZNP7b+yR
O4XHK46dwTz5q1gbo7ZSVSpGsUzFHr+a0XLMRM1B6fpdGBsBCoCxM4OHUnR+j8gZrJbkYTlCRv8x
h+6zJvuBuORtVqo2CWvj+inOtVlVOaoluevjXGPbHU6OGHtL4RRwzB299VLfGAckeUwslQe6eNjm
fGe7juqgFFnBfY/4S5de6AIAvhugLlWa5almqvQsKy+0Na/PZeHl9ZM1u5r0Quz+48vWT1hLgVe0
JEiw42VDyiNEP6SwTy2/gVSOYjpK+pz5DDS0IC/6ubabFhzNS6H1TCjW7KoLYcwCzdLnvcOF4VDD
6iSokfpilORewFKqSoBl68U/Q96Uk5zGd3juFoDedCmk/0khAVQFztG4588gNDdCY0L0Eqbo36PE
4m9hS6NqE5ntrv/BiZp9IYs6HDEMOYsavJdwHnRP+msxOIc+SeYI74gaETf3f5FWYKwUE+C467vv
ZrIB7juoyzpuGLRbp5cGrfSKmpZk7mxKdJVaWl5nSTg1XPwyQSbP/RFeTMS99BrRHMXqfByuFfTo
cxs7f9RQHc1bo2k3P/KGf/6Sbosu9HRTEZNIciuZ0lHtWJHtZ8csovDHvIu0bqAqkPR8zFFLrTYB
HDe+6pxdLwRuvMPRUO6hpAEMAfgGDcE893hKf1MG/DdpjYIo4RuwVb9uac47jrcCdJsf33yTaP9V
h6k89W6DEDVYrgm7fb18HxZ63T95PCiHZseaHxbngbwr5Ow98xpsGqrg9iL32Wr/wPd1WGzVbfM+
gIUnIPlr0N80pDYjVg/OxPwLqusGy9ZLz6qXGyVuM9bsi1S0FUU2PdChqCTwFSCo0SA6xFjvq0Gy
xFsqRD94yhUc5h6x4P3LXhkBbSWjh7aoevmpmPBtxmJnp/OER1AzYEeBsc83MnroBQzzBld6XxXM
S7vL40+BLaAtTqHBnUhN+QBIqbgGSkuXo6JH6qcjNVaCGITCRdGkpKXq+4MPvgXmvDpM1q6qnhmg
teUH9ubSjLfCMSpjMmoKyUyBT86BmBEG0Pz5ztH8qDZ4HgUA4e7+4HbzDXikA4nNI8M6fT6wXYgr
zC6AS+ZdOjYzgU7X+VraRJzoP3dwAmm48sScpcoUWKhkchKJk9p/pLeP0mq+RMA2qIM2cwkjlbRU
/xi8TZU0HWxVy3SYyJ4vo6Z7Ep45scj1rTEMvfsWhC6mCe9VmoD1GWx+2rKc67HxNZVRzKlG6WH5
FllNOHqeZzGv1g2iGr/NNEveBi6FIS1HhR8jwnjTP/Gbeu4e//Fu1jRaYMRQ97JciSyXvTLNgkru
eJlNagC4Xldei13h1dLNavEZzmNIJynDDRpSvYxSoR9/T+CcPrn4yQeg5ygn88XhdCXuB99V9vnj
8DivkgmHyZFt0Ghbrt4DCuNHR12SgTg0xxpHw78ANbog8YIvWqr57acDhcuJdmHhMxxKsJtfctxX
ZQTwwwtPp9wUNRf9hFn6AFgYM0P/6jLD+o/eLPHLEr/l+5wkYXLTfoq/Zzl/9qTgfbXfUj05ZbwO
e0uyHO7HMiSMO46Z5uL/AgwSRCg1ZC/lx7CzzO2GZuItuC4MHyLNM+PToo4AICvcTFKI5nmYW8nO
FvEhlQ64Z796q5mCkQbXpverYR4M2Db7vQSnEWJ0x45yHA/FnRFOnXEMUKIDw2eZUUey5hp/tVrx
gdlvIyP0DeIDRny1roz7p7NsfDL3GkEZC96Roqj3atdEN9uN3UuDlMYtIubdb+yuOkaWStd+WjRp
lTNx6wlbN3wBktnFgdnEF5ZXHOxL6XuT8HcdkXbODHkzsxHdaUygLDUt0+bOWiM9bQfkAhFGlPfm
G1s7aM8VWO+9Zk3fzcxrIjphz40hIlE1NpQjUxX7PRB02A5O3RkigaO8vMOT15vqw9TDhhZq3AFB
jFZKzKNSgB2VZq3XjzZ3VgGIJdQPDLSpvcGPx2KlozdllpzV8A+4co+CmjzTR8ZpodONqPz8TIhP
3k7PDh+pMHJGA1abvX9OZ3wPHVVodMKkm2GUD37FNZJy/tRVQnlK+Bj57kzHPFpgXesQ6UsIR6O1
jQUP6NSbdPJHklrymz3ih+lGLnwYKvEEfySJGAkJQxW3pG0wbYhHUWr7cmKMVt5u1du4BJqqvmeu
8gOXg7qCn33/C/56ju9mTmmex+qux1wdWouSV4oP1Vd2im6YiT1OQoXiGJoRweMkgAJICBSyK3yv
O6CNmCGmEZQWJPL4ax7fNiC3RwvNs12yK6NgeVTsBQZ11+YhAtCV/HSxb/iXeYALw89y20bRvt9T
IEFk0uf88FxxxNHC2Qer7/x8I7e5Ra547nXwc+kjNGJD4spm1jJaJv7cTAIXYbdzk7E6jL3ZnEOy
BFsrjZzLiE/XW54IUi2jO90HwyobVeb77dZ9CbBBcBbCoakrbcVBLbn/hM4EseECpSlwBQZ3P83O
KaeJF+omCztYEqjYkIojLskHBhf+CO5uOhzFRvX4Ra74djmnqTDsUqzeyNPSgxvCk7fNzigBIyaM
C2HdkbjCZRqPHh3kb+gNG5I9iVvNNUGbZU8nkKEJISqIJGoxLNoKGrj5DSJMXYKqwHcK75pMbklE
ZdJKCKZkN/WD/+oPdwcDJlj0HN5dC4+9IYUMkWuoMDlkk6Rg+BUigFJb0pbNHJa3yJv5nzPBmRf4
/i0vmhh7CzHelSGULHNuuvESb6YlmJrc/Pa9Ic0JCUrj0qRNp82NyBEC+g17LbIgYk1bRrMm0KfQ
duEU880IzQI7fQ3qiUIUzACUoWlqvO17ansd5L7qNXfBXtLA54Uvl55KlHZCAOZyvEfwwgv4EnqO
qQ3y4vAjSYmsMLnp4Xl/m1WQP3HgCyORuCsXspOvhQtMLFV7Bwz1Dvs1qVYf3r77N2H7fW5Ytg+B
5MXQ+0UNaO3p/gY49nezv/SF/0SuEZOHJAfpscNHEbkllHGze2TU7quubhSyyeN17yXhcku9PRfL
l3RcOZLaSpd9DKH1OTogO1hxi/mXq6uVvZYFhG6YputyOd/ZhlqMZBEQXwWWVPnb9NIbl/Y3So2v
H3NYlHn+XTdkL9+vj9Pu7+MSykua0u6ESjx3CrYCENrGN/OxfR/7j/pMJMFBkIjpY3gF5h1lzzYu
G5itpDgrrt/XI0tgxX10iFbL0KC069H5+g0U5aZ/CYIeMfO4OKM5ES//cHaYfSevM2q/bRgvDJkb
lQiQuDpV1LyEZaA25fs6WC7fzen+xUCdmGFIdc3XDfebEK6gt4oCt4VaYn9JCZzX3ctxQgYs6fO7
hew+kBJdgJXV3DcMXWNPa9Tl9kBPZAV9zxaVKyE0uDKVLjcvnDrNWt1mmd20Of3x300+/iGxrOAB
vFWAQkBv9EXn0m0gqZZb9frE3U6jmCiusGXjtNextVteGIE/ShXSRc0eXdMxL1/lLTXTNp9W+VP6
WoWDlFGImB3rCwxz3luwikHyoDDB7w/RqXy305jQcOKnFQCUfO6ZgqK29L4qf9WIXwBJUdP3LcD+
+tJUlYA5qpVnBPvGnKiH+gAHHa8JUjGJf6koBnAgHM7vhGlznUJC4Kbvh9IeIlhmIingRDgNDaec
G0qtzGgvcXEEk7/Dx7LkA5mUwIgRGYCzZIX36AX5YohgLgUN+UN5Jvy6YHH1VLWi3Xk9pBbqME8b
ZG4wz9FS9BWopnpg/j7Nv/BmQZI1h9ICpiVGNb9pP/VEg6/4VeZMtDry1ZGs6zMcedKODocELJm5
bYWdLKCle9JhSv2jokdzuLpfg1toSFBs5apgBBm30J+Q+3KHphcTX2M7Y3bTKZN4kGMowzERUW/J
M4f3rBfPZinW6XRE6PnzEj8DIQWBKVnHUlIGEHQprpdT38r5Nl274bMNX0ZC4IlkCd94n8nrF+1k
VO83YNPk9ICPdUMLfT1eMIeO9IluE1aqmp89c48LXJUPLhw+j2HVPdVJIYaMZrF35MCu1kWwe0nd
otUKOjy9BJU9vhsBOoVtlo1V2fUIuqBZBkRnabihFUDvohMgw1hMXy0HegalolvdI4b3Xl6YIBCL
Iz/VLL5ndRBBKS0W+XAdlUYIBZoFbOteL0uLjPhZcCVHm4GsnmCTlLucX2ZBiSc3rnslO9TEIswS
TYGOGgxB2BmzkGCDs2UZ/ign4eBXSA+FE6RFr9qDoAk6QH0dy71VKVBoKX4Fj7CWS0ELw4Q8Ql+i
8Xtcr1rZpNXTb1GOG/BYR+x3TBn7dLaQH7+WVhm/SZ0BAUCamk47H+II571k2pGgyHvDhSn9xW6b
s/Up17KalfKeZLTGfP5ZW6wAyHPwon/qNWhC7Pjo2mN0E1QFcUcvpey6trjAgev2PF4aSyWC6FfM
AFCgtgmK43pXzQFHTLz+rKok+81IHrgxADvviAO1/jKOceorCi3qrsR6CJxoSz55Zr6moZ1hrC/b
+VhNRpO5ZIOpVUPRCHukiH435Np3vpG4X/Sq7IdhETI99OZoJntjpoZ9HZX63muO6kqSSjBD7Q8b
3ENfbKdsLyciHGjaTsM88Gms+hca85U1GnXOfIHTBZJI+HbTl4SlaSNHKhy0Mxee6pSy+iounOVd
wEc+1sSVh6VBH02TJpvMfaEfjdQFd2ddP3zYZ/Crpb1Zfaz3sp6ZwXvaMaztycTed00geodalgdW
3nwrL40AFYrS7wkt9mzluP+Zu0DYZY8ik2b96oF7WBZwfwoBnqi+ocXZhdaJs+pKj9I6nX1Bk33R
dEGvlkQ2hDlOe/ytFFzdwTaN/C75hqwAqa+unvqxkzJYN/ATeIUpeIKYJnvV8t45i4m8rt+/HeKE
G0bEtNir94U6dvbye+7sGecyxACb+bdr327kfDNzare94GIbxG0IMbb5RM03J4kgCa5hfmiWbWLr
bhmwu4pTIBz9QcjB6tucC+l5WdbSiz7fh/ZU0lfEqhqnykB8DMmAvYSVZse6Icb76lFZd6Lu2lP/
27uScNuAe4UdV+e0oLmB6atBVjyFqbksdv6jNTFv3d6u7AVVybux63Zch8r+VL/uCsE9Je/jV/fz
yfUOi+Wwe9cd1Gi72lAW+kRLKlxY63rEAS5VwhfNtdyzyOzqwAEx+w9zI+n3r3G6qghFbRdaa2Ui
A8B1cKPBzvB1ShYKa5L3kiKvgpllzUduASJURasdzuyQDMIFBiugvp0PwrD5hjAj4/5RO4L760US
vMYdXmUGYdVOHRpRax7BPzGLqO674lTGCU6nsOQs9GJxjvxAJeq8WTAwZL16p7TNO0lo/JvrNMLe
JbnayyIwm2FzX9LiEJfWMidgdUAt1mHKf7S/DuoI3a7Qqj8AJm6fi9pWtxV+WDzXpRL2PK7QY8ak
ZBJCFoq0Lk7DwNbsSe9vnvshUewh2gy4ortDb2V/dv8dF/Luhf0evoS5wrmecbRu920KIuVL309B
2mSXsoCwFmbh7I3n/Kx3wOahJnnr2JRTb5D/A2zE+81wI67S3KkG17PtfSRQrYNxawitWdFlKDSN
eseJ9lSHnjil3zHLwgA5vao90SODLIYWbnd1eN8Lt451EKuBboVCxAkOCL8PGvxaDsLgZXOy3/02
GUSSN7AE3t4Vq656CWM/xX6YrxM1nDeNxEuslgmFK4YMtNW0ncusVjZBPn4Iykko9U7DKAV6cRuT
e3uTkfioZ5d71QA9dAN/wGghH55QbcTNM0snf3khwt/RtyQDZQeWOp5EZ7jbH/VPYVcV7qwmYsH8
NaBwbcBv1W8943A8Bv0aqQwZHqvJQpfdIdmZ3og3PPRLp/qcpaPqlZ+TTuKyVgx3NtRnHzWMDAni
WmOQiMF0M2v3tng6Pq+lxYRESBVZf4J6TuagDKST9eqcPKoefMGqT5ps6c1AleB3O5KOUDLl9GEj
Ny4OtRJIkkCuncjO9GkMM/kOkVfeIeo4bgYgEqOfkF/g8E4cysoAwQbpZzEQH+pHo6A2xyvEg1RU
8w68IA+stuKD6dbv6Xqx8hnm94ow7ValY2yWkl1K8AOjyoVljYGckgK3srh+pWFa27jsU7U4YTvr
5JiWMkjhmCvpRXVLn5MqBwI4aO9GVL5Qa6VssLf67+1Q+Md+9e3GKkMcFtJr/XKXy5kiB+dpDRat
W+sNBtDfEROOEF94cZnHHPcWW4VSJcszcMx3pSK6Hq/UgiH0CCgPitforUqk4jP3J2vH9R0Clhh9
a2iAQA1+KbATCwG2O8JQBcX4hibInU3eNp7mzX3KLMnGJt/427YboQdY7OFvkJYV+P5pC0Dc+GUC
vWuhcNIBfIAJOC8LpzJVaOt1bC/K70Tyf4k9o8kmxK4cD9wNIKNTpY4mk9xUqyQbQDLl5Yy+4mXy
Ef/GndeqVuTpdkielL3lBHc1quR9ZCyrcP4mi2hVvjdFCQlsMF7gQR1uPSKAHVPI2GGNu0IY1xk6
cnoI+XL8gT6+OifLNrNEkSNNxpqBl+x7Hdi+crT1dixdZZldMIjJr31GyzNSxHovAh3yfbSzr0T7
g6J8Mf2o/Zdnmo8FmcCX25970ElmbKgvUp/tF+54Z+DMB9EsgXLSPMuM5GeHtmEY8eiXazSJoiJ5
WdXFrwqWTDZdDPynbWiHZxlmBF/vBcy4zDzQd0gK5T+HN50mfoMzvHePsy5HvC+4n1Bg0MVieCDQ
zwfcmdko/QJcGueDBFDIzpv3l9uIwltNglglEVzgCz0JGmfwXDSXle6myh+EbNYTSYpKS2ogDwmf
M/gSU+5v127kXXxkD77hdbe77bd3hi8+P5Vij3NLB/uQ+OXQrCAmNJvtpBOvBP2jAnVkf9WUPzHt
Y8r0EWPYT5y1EkeIsFx4Zu5EPhVnOjZqUw/rrUTwlY4BOTiz7dPNdmSr1KerbfgpxqUf0sEcqZtt
va42Mo+zO3KbOm0ORrz2SmvvhmGI2jad4SjRXcjJwdA2Co9E6E0FYRuc6KIGhi49mdv59nACUUUc
FPFZSTwGDqSLmFjLTvDlQRxJUsEYD3SpSWdkSMbn1QviSiuL3+ylu1KZl4cDQO//lBYiPlPqOQA6
C6IeJyaF9N2cG+htU6MQtiI+VUqiT+QgsSX/98l/XSFP6fnZ2NhXKEnUVNJkBJYOzf3yJhx7gnnQ
g5G0lRwXrY7A/gq9+lfi6+g963b7Sy2xTe0PyxUTo6E03S4b1VdcNbHq+stGJ98XRyjAiYmMaY7a
d1r4taOzRdMKZra9qlpyvZNtPCH5CTCqRFXJJOHDMyAQ4wEvNTkE9aP0Tu2Jh8rgp1QIkuD6cEmT
kbg1NKKP/kcYQglWiljJ9q1KPc8O5a8xyEEbUjZ2xnJIdwpu4pLrDan344k5sHGI0NNoWPwHC/0o
jHy6MloGiXRKLW6+nouoaQft/8Sa49aNH22G+ZrRp2kDmskKlFdlpfolLkIyTLufMCGz2re003gc
ECLloeY08cb9jbpSlTtZUepLjr8t65DwuprskUWB7X9TH3zG/vy3+JkyagB8qgr3fPcPiebDkO7m
WikD1lZWtjUcah0GER0Bp+4UhTP4NuElxV2l0l0p+ACIP7p5w1TsBsBWvVbYaaHkyFTgJMO+dnui
0RrpH4sWJ0rvTJ9H2SjCoekcECXm+S6Mn5HFSUMO57RilX5QfSkMFAWz05Gjm3lNaJry0uXCQMpd
c+Kd094d1ilfESiAv8fcB/17+V6CV7lPgfGtUP4w93PLS8OJEtNKeYj5exv1gBlUHqCp0iStTfZJ
Qp0vxwRrbvhdV5RTcM+0noBkAhm8Gx7Ogj0fBkcJhaOwg3IbQX0uHhxJcwmYBc2+tMfqlpE12bru
/U/oAWW7yAOq7bzk+n79iNdlhawy1Mhy2V14k1E7hYPabdXlZ8dxd2pcguW5lQx8NbeiZcarET1R
KYnSwKEsO/EbhdEcY95psBfCeRQnDHEfJl0bPmU5G3TO2ptFh9kGzncWF36JwM5rAIu8+o3/fn/2
2xwqR4qu6RrPPimV14/0/3c3sI45JTVP614p6MLO6Ufay6qgR5osHiK62rIHUEP1vk+sABiW8guL
yGu2K9k88QtxrZKZep0EhPDoZWnXCosSPFTT5HKV2ulfF9WnTPYMI6t2kO6V9xdTNJPHqsLKy4cr
A09zkrZieiud7cYdxy5UJMsOi01vinJjdcgK/zj3pLcNBNVLHQRugRVZquJp30FTjZXxS7F4USiz
Y3aOpw8tRnDDfvNKvpWqlYh/BKcTdjWyMgfmZ0yoZddtNfkkM5RBw7xpiK7hbsuSGE0b1h94pX2Z
/3MQIarXTfKIRjdLWXrmRbeoruq00ZtPkaHyqqOkDoqrphdlSpmtZrnBLXPo/YPATI9CWCTE6AoL
NHQ9dIjYLibDDaG6wpkhAvjQMmWxPKrkRJHKGgBbwViKtJRIE623+QSjHRNB4FtSKJnOgRmbX0nV
saQAax40QjKcNCNoUtwDmruAznuaozFMzkXCU1zUVI6WqtgU/uiXPJxYQIUi/BfVQ4+zqYZaAljb
WWXgvJ9811HRFzBqtIw9pXZ9IBNcPetjPGk/IqN6ll8i2Yk/Xd430zNzomevHSfbe1oqmJ/mCAti
UZMA56YMI9ixEpoEp9iAGFiYzdLIbPfx5B8YljEP9iGWyIId8sh93uaBXo85ewirWHiDhlC9MCoF
2M/CdbAk8EI1PQBAKQb69PLa0x98/8DiXjHjrLbsHGs0QL48t39yDzfUJCPb3Z78SxdAwfbsDla7
UV6WvLF1pNVtdULmfJRoYkPmzglv2pAPPZ/dgwTdQIgwC2OzoNxwzkdG3//+wtirqVgN5UXUTtwh
2WkJYEdnG/zKuOzi3GQGmiDxGywioBzovOfa2Bux0rXBzPKoo5HrJOwlnsMVSZZ+KoPtzA7mPetF
5R2yI8j2lM1Ao+GDGGkHeG5ZL83lBYZsOnbis9kJnoaqK5YrKaqUGffGMoGAprBcgoHUujSMf6zY
PLn1vnV3EWSxiTJlFI1pa2hU5kWAFI0YkmpnWgvSs5TLFBAAwcKRC7rZ1ldoT3YpnzlG/T77S2/c
TPMe+S+5Fe/FGbnpFOiOQm1LH4bnCbxtAe7FkgqHfbze6N5Fyspa2NpHyKooRqGoyAob+h353j1b
8+pQcfitTsABDnQsF9fWLuOjp6TuKabCGRy9XccwlrGpMCpoZKUfP5oZWZx2vk76+9e3K/qeJ5e6
bd6+eH93ZrBDel4gWyFBn5+B6E5Tnyq2EyNyaCLyL98SRlinIHZCDk1JwUKCG6H2BBPhlEunBSvA
pGhLIFSOQun4U5+WiSa/EvnpT7Du3+vhyO2QA51AdYV7IRGTv54knQVlT0HGEs/rtVPpTKlQNee6
tQjJLPUisgF7K+ipbfwoJsGdYKGpbXUuShmTWjiVYukk114R/LRQHjIOrwGzhbXzzAKPigvgjXKR
3xyd1XB3P0TQs1sh1HqAXZcXTsE/a9JapV3c8IINhIQstxts4tlNcCxA4QsQBgmTwOl6zHa9OuEP
QkJ+g4Z18E4ZATino+DzYBBLTto8PC0QwwIeQZcY2EVnpKVb0qN+dAdk+4sNttS+frFN1h0B8BTo
EthBpR+TvD9cESLZIyTpizxzZ7krdhlcEdxo6+o+dyZwUopiDyrXiiN+6hCezFNP4cuLujpNA84K
GfcDqR8G6WvaH6uHEHutlphdE7IybnjIAJ85iqyMP2RK7t6DLXojGJLPjXzYmqwp91NxNCeLm7Ez
ICRHQJCqgZkMZVaJyAnMgoSaW9qwwgfQDgrOTWZrTvRWx4JYCA/1x8IOlvr2EZqLgUCwVGzJ2zHn
zsGEkZ+SlwBPmT9x/l3u76OY5jKhHnLD3QYhaw8F3VYX2NFnU59IYeAAeWgdPPOA4m8sel3vew/F
DZM0p8EndvWDT5ufI4vnZjaDWk78IN4Hf0+WJa243m5ZHiM9qL/ohS+nyPvVCij/y9c5V+RCLP46
hn9HwvMDxHZawKn5LnJX6C3i6TOgDCwc8R5tRCwdcIpZs3Wo22qfTrivDNf4HRt0g2SmBB11XTq+
NWKIeEIvG40ru2BAxG5UCD53W0lGCsyqYQRvp8uKZpOx23VZGlQ4IKSxyBFHzR5nU5AVemGmroQQ
dzPoBngQl/pdWsx4P17O842VWGiW6qIOJo+RjbLV7JBZqWf2SQ9njz+JsJJfUurN+xKeVgRnfxKi
cKzuXWW8AmCFRoHpX20E2YjsbF5yrKjY7or5qfkRiJGvvHtkXb06vn6TPHCETOMIB3QSJuE0fcJw
4/jQNllQRuRL2W/S4j/oiEop8wxW697wjc4v6Q/z/suXXpIQuF/uC/GESCrNkr72Jt5aNdSS6V6T
6C8JltWZB5IxL4FibhbwgH2zIC0n1kr39PkvhLjr1m0fWzZbImjOVRu23zJqHwPios2qpizg1n4e
8F/yxf2c6VR4Jb6Tb3MQ21U123njxHdvNeO1ahd1y6CO0Rd73zJTHCAmbu8BefM7BP5dj6mKMYvF
b8z9mEdRelxWEiqMQok8Kq6AKvJ8JO6ef/F1UX237TFSztYEL6qa+7rBmc3OGkCKzm2Fx3SbIa/s
2PQ+VTspxvwa2E4TJDAOrEu7Ehe0i3+boV2xndl28MmM3Cm9wbXYFPCeuwXeLY1Hkrh/9DmNNsqI
GdUEVXcbPZd9z0Vk+THQLEbZDLWQ0p2QGExY19+MoTno2lu7EVTtbF+Izl4OoHCuVyBLX0sD8P4O
VE2YiCjjeO6P5r5GUEOAt+Rx9dEsO4JvsxFyRVCZHhu3GBwApms4qB5AWzBMq8qVJt8DOWWPVQiw
PAdydX00LHCNtga/BhshpigY4D2ngeUUPX78FmlZ4Ay5CrxM1norg2IrOCI0jxMfMB64g+igJSjZ
NPOi+gYcc6NWP4ntwhW0vgvNsCHkfRFPXQuc/51VrvkmqqhU165CKH1eeU8lq7q21CfTl34vLBZb
YLE9bQLQ089CjvbNPcE+Z+VBQd7T4ZKxJkmy2Ns8s4v5/TSRejjnRpR7LHce2v4qCgoJkHPDWh89
1+EVUM9yH78HeVV2OuWRlGeh9pYPVfRFJh52qRTaWk5+Z7YO4fhqrWmNVBgMq7PLQQ79ZzFd7W5w
9GcfRbI/dVnxHPxgoLcbGHg4aQmNiOaa8k+6tuMFBBwskHZq4evGVMfaP0c7ANRgcCFo8tkiZ8iz
rckgJ7DVVaIaFfqJwPIPDi60wsnIzdjbxELOTTWc/5JvGuOipDAl4MKQ7kmqMPzKSSgNfOeTvhVt
rrpTIHXNahgbSJlHpiEzFapiTWOvRat4jjE7fH1Os0P1VHyqQaq0GpezLPr6x5mUkWuLRb9fSeG5
g9pu0hJjtDdzn6pna1nkR556lhWm+94B6ngxeZaMfh5JDVOS3lRyv4lYCkii/wNr9aO2kIDDM/wu
Y/CZLU5eyOZJiZeerVxf1FzVkUObB3JhDToEDK1n3vVOtvkcN0H1H2VHzWuxYPjmGowbX+fgZqYk
W9uexM3CBo1yygapCXuRd6EoyZHcbMYXal2+ilqRgYh42uNvSTz/xq4OCLYlVdIc/rvM4QiMdfNo
V+HKTgbCJdEylVWlA5m1E0llJYZ8RNW+jLS1FyAyHLzbPVystJxcZ72ZXxhY0lIasfTes+RFSPaA
c3J/2WxKzOMfSZUftGI/xu7CvfxaEik4qLn2AwtqnTyvX8fCnvTl342oKswiKOdpCSyD0cPGtawG
peTzrjEy0AcBFKozZMS36x9AZFmU0Vp6yifNqJIZCbeezMRq2mqqfs8TeJclpRVLh3H/Y6c8y8mu
FOc3JKCDL+LX79m/YZM0VYzZtnLtkKWFVaa8CdZUpLdxqsw72qmvqIAPpo9rRHjejhrW29UGyFnP
GUWxel6PwT6TU/ARpuL7eVgLvq4B2rGpqCPZpuJ7h3dQj5Mhzs7U+3RpBir1XO1OxAzNk1mJQ6JW
V9qntJBIhJmStVBmxwdk4RuaYD+WBdZ8iw/f6xClad3wtKZ+dgqdx1yhYuKL8u8dvxWGta4wbnAt
mFh89aIjfaZl9tOaR5uDmu4MUXQFJt0WeFGOoiVpzHKP1HaeFboktoafgAr/cS/MDVe185kdlpq0
D7Le6n2Vd/LqXXseIar00l4QSEgaveocc0ynSTgfkMp3QZ/4djwhRzwObbWnACKtFd2TsCKXed3Z
WdO5tkwEQel/HUuYu0Bd2viff4+29Y+hdmlM45u47639DHpDFyw72Y7D9dfS2JliySuzxspIgasZ
xm/wrFipxFfuz4x+LtRzssJpOwlUVEpa/TedFkM/+awkbCPIX8MjBjJMzPoyeMdPiDef9G14we2g
9wft53QV2OZcAkOJZ4Gm0N+CBwOtjaA+WMBP6KuJ6Y90AxC1V6ILKcSRRWDDNlbOmQ+poBIgqpBT
l728FHQB5ISOyPdLm1eQ4soewmOcbVZ0gFuXDJcUhNmtu8u3rAI67YvmZlWP0tI1tZ2jYG7cKp0h
HwNnXhgWJnTCbWx7WAvpbMZiL6hvsSWkDsa/kQ9XxhH2Rz+OJVIbrx2pR7m09ATjBcaQ+NpZy/tM
X7Gu8zpBHx0KXLoFaMJtMYGxeXwt/o1Vb1qxd2slNtea/DAKelAfpemRZWfwRzcqZ2hzfRckxiMT
d2c6wvfTCsYLjemeLQ7yMUMAnvt2DztCR0YXb8jvu0YuTMIjYp/p3SJXt1BQDUQkS3mS/CXX2xCk
FMYxKPL1RNc2/9HyTfSFg6gh9Y2JPlFHAAORveV/rZRuzbQdMb+UI7HrguxBhdO4JIq5W7hX4x1V
K5wZWmxAzltEt+7uPPAmC8EyeoJF2cS3wPGggno3pXfsETtczPLrV0rH1HIytmg+WnvZJed8ic/o
yhl9J39Hpdvyqup83LZW17y+NQ8+Tu09up4V7/3J6j/g15rEwBe9cL6f92qPu4Y64e3WdWil2NSD
oER75OXT8WvDnOEghVintAetg7O5zk5IGV8JAc+vyqzAkWbkfCOsz9Coeml/m8nEfXAfT1N/blxY
w/vJjWdlpdS6jD4lvhn1DeSozNHh+geZdli3SSuDN39VRuWSCRKYNzjKmA36wrDLG31LdviQd8vX
scIdqKWTokvrZ/4oOFKY7iHcAMbtDjQuldQoArklZFqVkNfScKy7Nr4L8s1goZ+0GJqCoASeTE5m
YlmFA7K16rT+78BO402hd1rEevxkTDkbcJCKuj5KOkwiXn9id69IydgDrlsGAqyNRJKs4WjtzCrX
OS4L9NA86HhsNe32KL9JpNOaOVnr4qi+66CPb6zn+lpelao9vCqrcQ8vtjJqCynq9SjDptNr3wky
IcZqLcJIDPGYYZaJmT+IzIC3/PPEdNpAMlPY2ZCc3vE/PipWFryIY3/kL8BwDlxkWR/g/n6K425b
iA+4l6an8IQ1i67RgI2ntfSDbsK9t6DolQr9jbx1obQh1w7zibR4LnFvMvFxXEGeZqUsF5G03z9w
QylffDwuLmnjJqJVAF/voVneQnVrPioGJvkDHEqDsiG1SykQvs+FwMu9+o5bNqDnQK6hCfKrbDjd
bqoHVPwUAU2g8dYcO2zZNxuR6sYaNDsLykrvYA6IZhAF/K4wtv9WiUMvo1EVqVF7c2SrRye4dY4K
Pl5rAove/CDV6vVz500XKRjhT3msljZMSHsmc0lgeqPNAKq5Ja165fyOUePVKnUL82SMQLVIt+Pc
3AvBm1fcHqAUh8Gxz1zzRaqxqYVfdQJpkcnJjPUzF2W71RR+5ZdcfB3w++oDHcoxFVYf3nbTVCxE
H2zYySbgbSRkBbKINa0c8mN0CcY4XOTWbaejZMUq6LnOxsO8v0Q6tv3LohFxUqf3+sr5GEsI2BXd
aCL9Qs3CbsFJ+QI6eJ6sWajelJUgJ/XvILnf43zuPvIojOdMeC6pcYHM8KOB+wIVLgaam4pl18h3
QMMJtEgwhbvzGZT++LmcBqx8A414xE2lfPam7GrMl+GUfc1sZzy3TLBfxsO2PddL37zK4lUAegcg
Jd+KmzrL5o+gUx+6QKP46wqq9yWiPEgrqpvWzoVdF2ZlKFP4a9JOlHT1d66XWNtR9PU0fx/68ElX
tP+4SOzpwJNR9aMXIL9jzbCBoJVkFaXqXB7DG1XxK7UsjLF8BExTPWcCjZtFzln0cA3eFcjenWt/
GxtsO4ZzkrJam4HrEmc8DTSjBVJKl5AVSgJputbFXowZMg5MnF/EiRtm4eZzxLqdSxlsh7kPF58/
FoRtgCqmQ+dGqIADqh+UHtMhwpREGtjxvJiV7DyXOW0AhjZJv5zE1L6Z87HO2A+FNJJGF/JLzzmU
WwH4BQrTiFhGIOC1BmZDMUQA+JSKypvUVhNzL5G/7ue1ZFwzDofkSlrRsRyvESom2PWlnC+VJKRp
mwK5mQzl7BFP1blJPbCBuvvWfNfklgoy2xsPrG0bDHEfLP4hH/TjwEpJ6pJIviWhdq8P3xjyIaf3
+xRk6bsOv9x0saclkG3njDYO0r78mSjhlxtcTMGanqaPccHm907BU1DzivWCJH1bYVYrW2JQ3a4Q
qMi2WW9co8wcbklkDlOdfMwgUXWymkegWu+w2wYB9qyodZgs7pXszNprXmE59CWM+5mGeG3bj+rt
ccf5FzpilLN3iCzkWC31rMj0KkvFQDiTYZ6sfZDRuuTuPzBZGkW98XE96N/ZtmOVHvAvMWkcip6X
CQMgzNpWOfLWdPnlyGZ9s+A4py0us+yiEKJTjBVQOjjM4o9Omz5e/sKcMT+kT/DGFzJbTzylBVWg
nomixDcio8TCAuF7zX88UfXSaDQ2CKlm4VGYgTQqDeM15b1cOzixDtucazu10aOv+OmYbLkimsoH
5bnoiJSEMesB8ucuIaJdNgd2DbbI9mvrdTgFOIIT/pq/7IcZhEaw6xyHITXF7qgis6p0BHz32slj
qiknCiROxDYMF3IqaQDGKU/JaRjsmfX5GYPUqmFgiOsWUmbvVPRMA7fbDka9EbBKj4T9OfS4978g
wm8WSi9qQkAbrI50qFUThYD2rb7KYqZYMKtnUbtriYSG7roGrymMyM1pGyZ09CJAL511l5c8MZ3Z
sIW83C0J0Lk3OPK8Y3LGjIDPnEjgxh23L3TE/ne6qBqDDreOzTitaqAXi4x3Utc7egfmyeG+i0T9
xc0KztT6Tiz21ftOKbW8tZ5W4n1gieg9gTCbNeMne6es6rlnHpW1i6QiB4LDUcKGFE3rKpv8Yxrb
WTFCpggZqM37D3Z4RX+RQv3O66Q/Dp/+n4dxQBQWmFU/T0tb58E8I2zkhyXS7EgaHQqfLgh85jYN
m9jWg+/G9Wd+U+iGqNtCjAD0ADChP4RBeott++86S2EdF8baXmO0O/iXYQLibhH2g20bJXibzrC6
kKRhdglfDOyW+3HR6GkJXTKC8v2qgGKwea/5B1wKsZhd+p60wvZuAkw0VgUr/aJa0x31SFryA6hT
o2We0E+rwnZfonggL1takjJJKiJzw6BsMRK8MMjADVKYQ5MJKMdQJ+5j/q75zkSEyR7noqC4nQzA
95p3TSCe9NC37W1RoIwfhXACVQdHB3GkOMq3tqBiokUepxhYQKurNlZGvHcME673ICyS40qzgaA1
57HRh5SVDUZKi1p1yjPi7uiaSPWh1Q6yjuKl2ElWPNHd1B4h3sig+pyPuoHmDZw0AaxMud3FQngR
8n5H5eKJSDtRS6ynCmfbDElJshsvsW7+143oiWkg5N4omOfJl9JBnw79jpsszuNb2cUo458nk/Mh
gjNBKoqGrwLVLhkeIdaIY+JNaG4eg0cxIQRAyygxWBaBw7p6w4RyMbLfEZLhU3OhHBVVCd8hCK/W
OgOcDhdKkPTP+M503Zbaie/MI3/zpG5Ms2QvfX3gTwZo/u7tMWpz7Gkkp+H4iJgjo360n8O/BiSS
YXFFMWErKq6uJz8xiJgeUESJ/BJoX+fS23cqmHJb2o9RhJmSZxQhwTG0T9EF72j+oEGjJPzJqoID
UdxNoQMOLqaf/YDCtc1iAWLzEtAfK3sy4v8PXrr6HCtxIzS7ZPAd7bVVA0AYwQHjqQ7k21jefAcO
JJwlAvdX4DXWUHs0E73q2sblpq75GZRbAE7qDOesamrw7BSGMtr8lyFAez2g7z40ZDRwDoMKQJFo
0bmlsAWNQu3mePxF42ORY8hk+H5RpId/dDNkHuHXCE8BpcOKBfF/tycDyCYPvOlaIDok170LVN/x
YD07tvG6u+EP90Tiyg8DQRt4GjDfmnThJ9+VLiJbyOM2ua7jd4VEK+B4rautKbVI15vjmeska2tD
uYi/QTofaiv3g56CXM+6syAmEk9yhN367BDVGE7aAYbInBDvGpHmiQEATA4t1aAyQrspfWtttkus
/9hqC4inGJgvpXHZghb3enlZ5nZw7ZgiUk+ETr8THVyPfsHz/8F0bqoNYfp8OnYZKCk9AapRao1a
eVlydack+oVr39Bl3AHshNgBqtvzWWJ5tgckXyfahyS1SJpraoKO887DYiIdW4TolRwRRrHM+L7v
NbRv/pdDXDn2yiQOAVBJCQd8uf12EPR+mEZp0EWmJE3dqBmpuX3ENRlJj1hgRbn4vykpRxBfcYhm
ho11FdMH6CcTh49SrTcni3LwsdssIyDrPik7xtBuRNq6HRwt1auLjQrb+Od63dTFGL4IG4H3EdpD
QPouqXUx4Bg/Uo3Ot/Yaa6HC4xqula3ZgrtH0LudOxzAMmD/KvlKC/uVP7o9+iqbyjaXhCEHMMRb
mVnFOtnjCfdbslsuucqE6HdD9jctef0f8ipug1lptIfmomkrL5C2uz0TS83V1WBu1gqw5qPCSo1g
HO533X/i3rR09Pza9h7bAm+PCAMDtESOwWN7ncABbE1QBw5BX7dsn5MtYcgZulCAdFilFXJiV7pC
gq8K7LYtk+5HRYm7iSx+kny10IMrc/c7pZoGg0X9vlgQIW5H8m2SfOOnMwGwZ73bjuIpqVFh+2G5
5QucXyfDpV3f4mRle2NcBbjY1y42D2sSTWO8+2zQbFDml/iJN57M8/nDum9m8CG5MK/APEw+vZ5V
iUC+nDgXI/A0klQjKdNjdJ5rVp02akr+O0QRmWxhL8dY18+9trccBgu/QVWF0LjtMGZsFkUVr50j
hsmYjXdNIzacq5rKflnCdCiKFkBCUNbTpjb2Oibm6TkyuvPQWuc6jSiSl+DDRUvTKqtuS/CiU0lG
Vc5vZMdgYh8zBCXJ6MmRWFYAItrnA1M4njYDIpeJldei/Ec/m+AzKiSTkPRATPLGtK4WB5p33qYs
k1f77+KHX1bIMwVuZhAT8X9xTVrhFOw0bxv+hhe8scxfGim15f+tF19yh2k9MbHenoNTF6pctCFC
PaMdymx62zIO8+cE5J4H5qCmpbAVNzRUxdwhJqnSZzZ9JdPThG10H/I+pfaT/LFHuLH4l++X/+ys
txatoWkutlKANbxMftAb/ml0V8bsYCbZlhDE0Tw2G90ooasbM+IaFgAyJ8FyhZNOII5nSorogjtt
B3KXlsUTwbqA3z7J52A4AVO8AxMfVFa6LGLMPBF4tgrsUhafCRjIIjdaa29tcpU3u5OEdtW4jbpi
Xdt3pHbJk47TXnR4bfeifU18LzPKCXEb3XQrrVYiLYIJ0jSQxLzt0h9WoMAEgh564eTzHKz9updl
CTOEflBUcdfi2KWOtKlyTsyy90QdumnUWYxzyHyLLSKlv0bwEKDiNrkMo+lVcg/jVREhJROkFk0U
fA7stU3z6V7C4Fe1NtusW2ysrmAA+ZTdHiJ7vNrkEycnS/KJH0tG2DWmWiuowgwBxxZ7F3aaSLww
uOPUrFUPwBtejXSFaWbEr/SzT9TuiOG9wacUW9s0QeEeQUlfl1lKIb0zV80tmQPKXsQ0GmXp+Mb7
JYUquQesYpuHVK92Rm1GDuobrYhLN6UvD442pR+xhMOKn0vODPeThQuVGLcO4yEBgy5Qwl2J3moa
qtXVVA4wbuRm4rmjZQ0xj1EKq0VWBL6lbCU/LtMJzrlFUENt50XVNjdL4ilyVfyGRDtaHuVsf4Op
/8ThDKoNTKnI3qR9vOi4iWvmxFno60GM9knPJ0JhBTBdUTUhfrNzPQRm7RRnqV0nBbCb4WhAzLrd
755oLimyMQa597hTgBJjV7IsJt89mMYnDYPT4uEzAsyFErBeE/RFwgKHUladxcSrnZZw7xT9czo8
IG/ovud8ZmpJ3F/Ooz9Qd0jvvmGNUruH13aqagQvy7WXYG2hMXyarqHeWGMai4Dz6XeFOOAOoZuF
MBeY36dopZDDRhAYSrp7ok79XfyW8TMXd6RTIqC0ELPbJbLIc8BpLUWZLqAHKXYa4iGZl+aIPApH
YJ5n8I+L786qt+IjC1L1FoXLGFYtaYAbRKUDZfpQ60aeKJGHSqb6fSy0FA5BUu66cwVrAgm2kLsc
lGvFD/fHezm9rEOh209gTxk3MD2gmnO4v1fvQX6cRjcd50/v4IHPkZNeDkIBwJ/TsQUAUSAL9t3W
1OdaA37EJ7kYLgjOHDjkT2ImutoJcT7QzODXNXogvu4DB0EfvbDXwAfL4UoqiHRJLCdrVR3idpv3
KAzquaX4Co1jOleB+lgROgF/R3R19+cGQxS1dxD3Ov0xlEZjLyHgpmJl9dSi74rLI6V1exA8UZ/J
Aeh+1Bt4s1EsJhni8awtyKIwbi6oPPc+o44hYccanMhph4CgfSGfgxLX/rEMa6CU7hUQgvNYByM0
s3gRforvBjqymza8tupwAT1+LMG+UdmxoGwP/OuG9fINKbc8W/YxwCbmboxHqbLjhpOyoyWpb51Y
BYP/5ADe1sJ3Y3FnwnrVIp+/mtbpYc4pJSHTqJOQ2JnFBWk6u3EOh2Lz79H5rW7FfkJsE3MILctd
K0UMfb7BBsaKNj2ZWPZAEfqwML1ljpNLcxRHc1R8yYQTqUNdUpuaowDve+43xR7fjZC/QqvH7Wkc
WHbWhOSRC6uWTLfPUZYAiseWMkPdjA4hWgHhMI0UQViXf9Ek/lzvwA9+OHVAd0ZBGTI9J+JpTvej
eJhLAOXLKXiWDVJDfmlNX9XIhf69m0d5RgfZokhy1N609YrCJI2SwFU/1DSNYbQAMVJOzW6hmq3R
s9dsFHBRXXjOsrhBCXMGofq0Up7zRogmupzg4HDD5hw1NvUztm9t2hgBxSft52vPrqDut0xPjAM8
Zo5I/9s9hMJqnKokb5yt0JsQmW0nrNjm6EZYL6mZQm42ojYvCVWLbC2mm9GZSX3ethMuBg2lFhrs
QQhTfJC1ScvcqQYPaSZNnltiNJRitR2L4oKQefw2rDSPr1lEHW8HvyBIp/+ybuW8DXhOjnyn9xmj
kKSo4HmRYhpYZT2L3tFRqohW0AdqCEWEhj0wC53t8wzSqmxntFjIXLunH7jnr4T1OJbEtM0RgOuz
qSndESagCR5DSJVHXNpo8kaCqMv5CVXX1oV8NtE0O6e+gDxEv7CFqvQOPLNqN3t2rgAEXSMIezhN
XwTLQxkHNzdKodh+jsXvEzcIiKr8FNksbV/voPdk3DUTbamva75qIOl/SwQVMwYtbDRzcvCnIUe4
wErW1ER2IJNQNb4HAz33FH3dc3hNutcTGwt/CCeMCdagvXM8YHsB0Mw6t/+/1e/tHpYoM7Rf7UOD
3dWS/igTEWXEsMBAtRpw28yAlNsYf/3fwwicg8aU+Xz/Il6ua3KuySQnYFAsUpL1XLDBm0v6G2nC
9aNdYQTHIsVw3MvISriBAdwZu3DFSn5KeSHb92ed5OT1vrSNZEfLjS4EzB4ITC9Ofz3rIoM9u55W
nUrkAmUqdGfMDwp1qYuF9DwrNOU8XVAsKhi/bP/cM0lpagE8NnIWsG8viN+7uCdRqcrH9HF2Dtta
xHTrwHWJ9Ay8dbuw3D7uyJBvpZQsHYkVOtZuiayT9gEs2EsR43J2nrVgDCqmaRe/nQFW32jeK3EQ
Pq6YRNg5P+tQKLLODhixvWGz7Z6HdLmBE3M0i9lHUViSfKCpJfaQepj+VfcIqj4skYkKT+sJrbly
eI2Bnf/MACQCupbxLyXm+P7eOqlrqDLfwRN7Nu5IPGstIl0bvmFxN+3aU5V4J/DR6D2XBBgzAmnc
9PtM7eYZS2jw6wmeS9XdbBWdj1aCAFtAsS6e6J6qHLMOxTRmALyQxQAWBau/prTXWukOAnFgop5n
3ox6vgR10UjBbToQUn6It1zzzwqOw/hgvLdO/MLH89K5XH+XqOTbrhvXp/ycePFdHdftsGlktxUM
AuZaV1hQO1+ppsGIpNmiPGxuS0st5SxwG3utDqLsGZvg9xAjpn6CHOf3lZauXA0d5BryeBlg3Rix
CTqPdgqPOCuggU/YkOkGUPR7JP50loRA04XmoOz5M7eCEa9WlA6T+xMPKj5a3sKhRQmhdqvM5g/J
gyUIR5Kaa2tfcebBQQqJsdmIa2dPJVVmJsg43iAy15s20ozDTNRmJo1TG5Msu5PD9akrSVsFlWkR
yDL3TIyoCUovASTyOSPpmrQQycmnRGemHjhs+nzbW33Z8Z2nl60gsRF2+ir4vBgTIcBXxu7OmPAc
MOYnEy3mYXwROFFMn8VOf5nQIfue8EBEffc0rOvOzchveubtMoGKkCJp3tPLwI5QYMKtOS6YTmPw
UPeBqMycoVpqW/89xUeoQ2psaOPm/c4LUMeIPKrBfNl6SvAqRSQg74ifsseA0+FcmmO9ne4Ealw9
WbM2RgL8G1eg5D9sHyOrPG9HQXZUWE0TsnhOGrqDPk8pwpkFwhV1ZqeDwVeiQwpvkUpUZA/PhFo1
o/rNHL7Y/8+c1kSRMg6tFT3DL0aAse98m0OqIj4eVDZUDuFJ8mTKVNXzIl4uReoQdRYQvKaBECB6
nMJzRL/DlVXGD9k/xJ8quJPa5Ll92Sps2+Pn72mSojWf6MndflgWi+UKoZPR7kLkZy+7MfgZ8tTd
BXR6iOgmM33ChLRijWFoLmSVz3uzS95ATS/zUd1BwB9FMPB3FN7lUN51uGMilzf5EOGwJvH/OnVF
ulaHZgdrCVPhRBmnAzF7K6xL+0apYur10FAYAz39JGpUM75k91LVPv3VipsOwWSX4gHHrBkvad+E
//Rnn9XFZWTgcgHELgAqdf1WdDtDhbyePCiDtuv96L7jaJlrImYohGfSOJhlQOQpnoIeH/81QYmi
2XZSVgSLEU2AV33+4P4ioKf+ywWNAABy+3WfDVLxM134T0nbb9tOHsh9V2hlh2H/q62fjolOmJ1e
c0Zs96nLv9jRdixS6dOjQnTfpB0QtbJXlVwAUZ6FFSa6qXRtzsrQO23rPxcm/NdUnKcMJxmEkNpP
aGD2e5V+rLfFODyZt597l2mVZKfSCVzdZT/oxGuGYcmOTmaYJvAPIzv1QFGiaZFwZp9kcuktG4yh
q9pEaLEBJEqbwwcHv5MDwjT7nawdhMSyKy6kUjp7EvA+WkzGQXD3NHo4Dz7IRuc/Ruyz4DdXrqg2
dwlmdJ1jZ69MuwV0H4WUHeNp61aGgWbvPxdQGbGFQDgVw/NLg7qWiqu5DUCBjXXYfCZ/wp/EAcjy
P85TbXG0YKiYdCRmDOoVEG8LI9yvshttiiN6gEfUn4o8UbMMrddQeJF9N1MXffuAq9zS2aaS88IV
wzuh8FMiokZvayx6EkWvTFMrNig61SpBajhXNZ/6DC3UgcY9jqlI4whMZ5cRJZ9PS09IxKpCxspU
SWU4F2o/YkB+yw2xtdvL8e65tfsmDZPub5eYGWdF4pTOZdoZ5R3tDFByNchma3hYF2xh6n6vGlCe
3fhLFMJnzRWhUfOehXkOwX73ina5MD58FTnmgvnwMYgMkkvofvIeo5HX04+DqlUYAzvZ7zigg6Ih
5ZGyRWKKPidyKmIkcbrvG96SeyJ3ve8UvGgA7T9+2lT1KUc9KLOx0XZtGOaSJDYcM1rpLIHb66QF
un9rC3mVlnJCryHrwupPVByadn67vAiop60QPAEUvVimN8BEmtbnODvEdbp1ywvLcdKYnZpao9qJ
IrZESJEGecxFuSbgNgD652tVpxMIppaHrCxuvtQ3XBjxdfAf+LBAKyx2uUilHpwZxOFdU2wapA2f
buNbTQuyKB4bnPRhh3PuH1ScMN0OnpugDHtXMgPVEysNM8TAZqvYDqSdCBXn9mJNbjRqanVxP29E
kjZkFWFrq8hVp0pDg3ZPHq4Qb+OknjfuWpfHwWtuOoIvIa5qgCTOTr4G9EjJiVjgTqPYyUtp6eLo
BrY4C6UWqoJqWqANdFIs9sc8O+yKS2oABVffukClX99ksYEUcc0sJMCoZpr2iVhjkxF+Z4+UIRhd
EAbVQALvPD7xGLWsIUXJQPtg21g9LQtwoT/zgvgVCsqD3pza5YqcbYFgr7DxOgygaX5VUbnQhX8r
JdZEbDfSp7nkLKCHiiGExGCkMRkq9p01mPfWGQm1EiCfAEud0jJtVwiyHboWI7BNJgeLcYDt557J
OX8suMlFloRylgPTAx3Bpw3DESuxAz18WJbZL3mu0bub1ckAG7TBgjwBJlR8Qv9Eqq5t9fybzHqE
rYDahjz/x2m82L5Q17v7UcoZKGsqioKLaULuM2ZoC/6ISXqAUAPfZbxu5uwGE/hggdze5H97SVSK
kpNHAhNvxtE8ZEw5rKaKL6cY27PLKd+1Q4cqR2HBw+UV8AxpDCuN17VklWDfPzPh6izffSFER8vv
a/bINHOwJApO0VR3b/jmXbyp0ltBEnza8fgQYymsybFsJsMHs3Jx1D6eaodJxitV8HTv8qXjkK6w
8+NGZ2dSWV1D3baqlHpqun7i/dSnaMYvnIQSD4NHAWeAPae6jZA9Tl0xzRM3xxhG6y2MwEKsUoAt
RrEQV+OoJIG9PUO7gywAIrAvSwpZCQE68KfytXIieC7v+Tm57+Tj565yfrrqM6a2A6APYo7SfZGw
LSHAe0mqGx+mXzA+IND2aTuW2IuU6GK8NgxO4grpzgyrqTKe6Q7056dBb3teR4i2SjnhHGVx+SGD
FOmb5a1j8Ze/hF3L97wd7cHucTVCujjDShCe0p8sOBpyLYHFPhaAmIK0JRNRp0k3NX2VtYs9OQT+
dkguIPEFub90zTJ+mryMuqDX6/KK6hEFeCiruVKdQ8sFI3pNvUXLEcEGOGMgvnluYJ+3kwaTOmhJ
NmTXszRs4wGdil/oWG9pR4QeGiHoCiLMOzrWyFbhgrJaIL0jBF18bPIdvItWCxERhhcikAYqWjZQ
GRNiLrvAnFPDcVyZfwL8dkHffLz8HXl6oMzeXcG7H4k0UmO/mng0OSo8F7qEcs7cen/HKSjRs7Ms
FcDt8X+JqHm5DCT5LldPQsak3r5kT8K2Pcja94koyuZgpNBUrNbo8EpOisNDKPiU6OFOoPtNrssR
pS+GYkSe5KzbzatSJm06wB3biQfecNh3ZrK5ysuM8Yp33px5S/NiyATQuwXtWRUaHN1/C6pgqf6Q
DnTApyM+dOl92NW2SlwFKyszf9tkATknyuy5HRqtGgGn5MJdkAVTpNSioJMmvC6ep+W8vXRYhGLm
mjdqzUG2ouq/3EBEqOUPjoYgtVkPwqWZJ5u3jSUHfaizsbajR1KzJ9qqMWoQg8jIXarnwRTP3jLu
arVBIXKccfW7Bht9auzDmh9ZQQbuXctXry6dOBeT/eSfPnSuCn9Mxlz7USX+4KtTTDVQ97Fbi9zb
l2zUNZdOVn6UypbxTLzwfnzG7fEsB4i+xQk+n/R9+bHPfizeX9/ocIurkl7mLqFwK1bc3sthUYtN
ofeq6S0QlCEzdb5VQwdyweAmKlJaTWBy9gykcXl8PQUvzGTsfihA1U/5FNRtqU8s6lkhGNPJQ+sg
iY+LTIl+dC3WRSsxFDWLuQlFsIfZ1gqyRPWj0YFY+wSvH02w3/Nk2jX2PwDPQkGsQ4yqFTjGpnJ/
I3tsnYxhFWOU5lA0KaQPF70LCeiYYjzl+CQb2cr+4c1eolc8H/dFeiVa776FC+6EkcW39H4lmXo9
dKHzuUeDD6D7SJU68LZuMRBtOznVJNgKGuY5TsTwbr32tNWVjSws/QsVcdbkKU9yLqXfbxvAxk9u
Z72JkAqx+3HV61vyKmPfYEmMNkIzubZ1Mln1eCPowKInihY1aGXhcVdTsNv4dx4HrjZHrGWgWC81
eFGNqfrBrr4NitfR2+iw0oFfHPS4hVlFJYRrJxQNC9BqBulgomMiwXorH+nE7GfySrS/bHV8iyTA
Exm5+7ujYTuolATVwaICRro4xoK4EPA6D/HrrcEwmCMWM4jn/T7mlUX0oBY7gOXLSQe3PL4fIurw
uTrAnXaWMPD99/UqvZwl7vUbwQ4RfjnDRXkMSdrU6t+AuD+2NYetT/zhBO0K9LcOmTPHyXev2tne
ZhMNZ8qjidYanz+X0YXB6blJwS94DWxr5LnXWgXsiaxQWrMWGjZmYD2DGRyOxzLmFvL8w8FnpzEy
TdxF/MqIq8LLScrMRTmmyOyOrEyKJYP5i+HV0gm3Qr7MQqlJAU19kvc3SXp3w9CKeulpP7KtOK80
p+p6vcHfn7/LH0RXSh37BeenuXY5glexsQw6Tj4x+Xi1qmbRbGVipnCnIiAdnzxjLNyEk18uvBBo
M+aS3BvTNtkWBr17vHUrGcB0TE0SeB4gMDeCuAkT3bCNDmA8RWztNZwnga6qmrhgpUjZ67Bbvye0
J1PU0ZHJDYPmSaLgMXv2h2n/t8Xis/F0Mu40rZyt/B/jojOSB7OstwiuV9TpYYXIzntyxAK32UO2
THoh9QEDNSYxXPh1xpCixobC6Z1A2dU5E34Ch9M52gB5ltxZK8kZZZ+ZmhO3sfX8FLE8gW8sNDMy
boZx2EqyqqoDPIMUdXLlGja/t4URzqzxz/BQji7qZrOp5F80BnSjsUV6osD1g11sNRRK37BHWxBF
l5OPLP2SdhP7wMZq3zkAcclhlhPNyaYtZTCeVIeJMWuhdbeDlMQvJ9+uQ4rvHLODIoKHQzUemZ/Z
8mpHWjoNuMlgNpqFo0z/I7Mbaoq3aIaTOYXlsOv/
`protect end_protected

