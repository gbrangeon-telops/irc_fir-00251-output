

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YdpNuWNv5ANxG6sesr+pii9y21Kx+NVDp0WoJ8gKKxKHNSppxy07GkwBsVP2aDgHIw9l2ULLZTNZ
WthaAb5amQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kEIsWLqGmgOl8w9T2kPb2uPP5XenCQ9kpxljFoCEGisg/vUEuVE5EQlDS3+mxviS53p6zH5m8hA5
bszDfKwHD76EbEoDDpJWL09MvEqH4hbAV7G0A9Qe7ZciYDi8os/DYZvhR8zjbLils1MINgQgL32T
+DXtGPXNuzJTAMDKzws=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NxGGOrhc83L0V7+Qmwb6+Gi21+qsbQ+hA/5/9jysqY4QYAqiXfCrWB3N0NrVsGWuuTvZXoFNcxot
Izvlkgh5KOucyz0ezFvnhsYziU+FkvqQYf1g82Syrsz8zvyVWXqii6aXcF/WSMwXtiDjm4MiGpFm
yTcu8CcJgBMXYGVZx6nj+IgO08YgHCC4sfTqmgIgkxkmBrOsiH76g2hPxvXPgVWaBlJF0bS/hLIS
Glmsy0cU+pqQlcfbTEV79W+sXQ5Q3KPQFXj7AhMrHHD9esRm2Isg/tuzcRVk1cq3LsMUN//vGrfM
OKoYOozZxl1/IflxrtIzbjclaBUaFr5bvZYMTQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dIJ+Oh/ID0KokdCrmxnp1QfFJ5QZBtIG4FQx5Pan4DTwhUxDWY/BQobSBBDXzWh1TT07UPg0V7Ui
zobKMfHgBNkMD8/PoD0AIDWLDLeXLvIJje8mGtE07uncec5mJ2eGa/WSy5sFj4M/Vdtk7C/Ab9LC
9qAaWZZ72ZUoEHuysZg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VglxNkzPd+guDL8DGRWVtgWGTdJbzbKKn0hBXJRIK4IuLrtOeezNwjLTIb0FIMSJGqYYwUrPN3z3
TVnjDJDaG+HA47egpMvivRkbnfO2/EAJtU7n0hK18OztWFzW+yXOUsOuQnFS20EGjEAN6HCMCAXS
ralqFAJsvMtY2y3dJNuE6ytT3WYkXmZUpTrJPPJOu2l9mCOnHkBU0dRG7RNYXf1tEMPaZrHSYyvp
XKWW5CTowIM6jJQxDVSVfwprGmWFUVJFtAmp+65D3ADXiHMcwre5cI/ty7nYS3euq41mrkrZyEF4
iH4/gU0xN9mM3aF9hBPzu3xQrdML35ONnUZTzw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13184)
`protect data_block
DH7dTensakM0Q37fpx3AicURbbBNLBIr3RHckopNVflBWVcnhPOYFPCl6k8J9nVCEeWqWWRshkzp
vHDSL4rrVPdRdaD4ZJ1M1up0tkIfS2DkR4F0l1UXnvzgB9fKLiBjJrw60rsPbBzYK+Z+poTkYyub
1EnJioHaDU8DVx5S6eALwcb6lMF78nqw1ElyrKudAznJML0ecfXxnl3CG2dQcj6OAJanfFdJABUb
WgINXtfQhvSBC2yDMuZPBGXY9XL9O7pneqW52D0SxARkgcNymR8mRiooHJ/xthVRKkgkg6JM7s9r
HVfQCEGDlmJQEIZGAxSRiUBIBN7Jx7BRAV5ggy3IgZ+CYYajAhwVM0m3a32G9EOGG/i6RGgq1s3W
8/cMZQ+EQuHvyDtsP6YEMD0raeU3u0rx+rP0Qe3NLMXoczqJ7PpEzMuzeqsvI4DEeYiWPJVbH8Q6
8IIuJrGC7iCVrLd9R/hG2zmHQnLE4hFQW5xLYoZiy3xROcEupGNuXlQB2aLtCAHgHHS8tcARbzwx
5vq76hAO9l/qtIDd1yix1TXwUiAX4Id4mV6N7i1xurZ1bu1f6I9+JktDUO0qW119YeeQ/c5X8pfk
1KWBvgDWll740WL3KeaHsI6ob/bDfTGMCCqS0zMQ5MYOpLekJGCeo+OibolpHKqm3rAL8r5cJDbK
IS4LXI3RycEunzM6X0YDseuTf45QNp/U6Pxm86O3rBCn7ul8PrmDrVqiipPRKMchxuYJZf2XiRE0
X+eU5RPO/lkCnCYWuuk/zuEhfLjymnbY5cbt8oUyDEp7JtHNKxJbqeJeRb9jPmDKTY6D5K4KzD6F
5rxwKY1Qbg755zniNpZ51oW9jAq8VCGZLy3bhxG62h2tF+roM6QkL+P2GxtRxNpeVcLJjUOhXM0S
Fu0MwG9hRVDGTsPiy3Kj2cr1/+HkjBYKlUzZkIZNM6XmjxjeqFY9UV2FyzDpYuq6VsD5HUTAPLmi
TBwf37vqvc8homsKmvnLwkUlAo+P/QakDMrmOwzsncePnWXnYA4g/BrVfRwT0lGzk/5XNhg8j2/F
zQlf0Ynp1M12QoskR9D+SfuAZoxWoFVT7sRMyTap6KK5n8ASmsskulNHdZvU1wPDqGI+VPdnNUOK
nVjBbUUpel4dUf6fdToiOjJGLy7V4zp83ARuFfTdr7D9CkdgpBbcngT5HhzlKXeq6jHBtdxm3U2R
cEk5FmcCQQhY/tcN8RKzjccd+3X2mQFeVBb2mauFxRs2uffk+TFFCEk0/QHAtP5STjG39Uyzn0Y5
K77+kKLQrxNvSKPCUvDWGgs0swKBAFA37wEGU90/B29c5X+1T0DuvfX7y1mIq7Llmd5FBn4mQ9oA
xI0j/kYenz+CYrzvHBf6RU3I8u01l3ToFmJ6efF93Gh2K8TNbYYxnbjdoXWbk0kOAUoAHGKAYjnU
cXC1JK1/3dhIh1b0amGnNOG7ecUWExfHjWSehJxeToSZEWOocRtB6bSmc6ba9TCV0cSA462ZhcUa
Mp98ipt3ZJBZIaja1R3IIy5BFvd9X1KLVZ4ww5boYOMTa+oUeRsgnlU6QgbH0DxZIM7YB4daJy5d
pyyQZwtO1WcX0ga2LgkdFbgxtZVVzPGGnQtTtVzpHsXoYH6uE9eCatRICymrjNpvXvS/4jKDRtvt
wZl4ewXZKjHiAbbRoSfjf3aSdhomtRdZ/oDeWheG0sRDT+/ow3ySfG+Ab6RSz4xIqDuWCYtxpLfk
aXgjj0RxplY/HPbpnpirBEAyHelsOkdnAGai+qIWH9nDrKS3KNTnFTT29n8ye7OK4O2Ztuk6SxQe
esgbOOLxFOWdIF4BUA2mfYHgg+tyQs3fz9q0ijcsE6qB6A6/3JHuqYj3dxbMeSEJHbVuIVd7LwVe
o6JgJjhZnTKJslHWrE6kVOKgDJR6n2YqYHeP2AjJhrery7vIQW/pQx5+r2VSQRsUGiEMT3nntrns
DRx5AXtGKn6gWOaZas/1pdBsXBKLBXm567p9RPq3dlH6wVxn2lq8IMO5OlnS8aTk45PmRX7WDXRx
qjc3nOBRFo+QqxILSWKOnqTX0q7X2q5IJtU+GSgT9DrbxjAEcLFsoqA+6dsDq7WKh3pDaAIuGIjR
5SCbt5vwhsgUQQzWiej0KZfDvm3OcyoR8RfmtRkU8P4V/+w/t43aNo6L/odzslLaRYGRjyjyBlIC
x3x39ULN4HQ69ZkT5RI42gEWDG0t2XtHr8AFtwOiGOI4Z93FyxTYu5nxCdjmvJ9hVnMnUDiHEaKk
SGG66SMIvvL1vaARN0xbMGn9lcPhza02NBiiMTMKXrrjHzEP+ouS2oPtjQdoNOT5eKQTycB79Usz
Z+uQENMLVf4F0Lt9NtruBy86f8joHxqEx7fP9r0YSt4aNe90xe7gbDuby0+3PG5Sh4FIAG26cGdX
Hx6f54cxrsKDXOuOHHGomIJ9IGu9APgIpcHeugRZ0Ad4OnGtqa0zR7VCMk68r3F9MBhzc7CtgBIb
bLsZocCXmEHpaChl0pdY89xEveWsa/J2hfkZXYF4higjkNDMdqBwspL2mh3Cu5hLI3tRMHTlMqlG
8tTO4tbRwQ9p0/pVQqROHhrElXS3d2NYXDKKx9cuUkDuCxqIDN4NV5bztZAO9Yp7kf3n0O2hFKet
FKYF8XiLQAz4nZDWdtBsT+eTuaGXMBZqG3Uj9V2mLrgK41Oa+g35VPwB/JSOZ3JI0ggXEgny0oa0
Z6cN8YtcgqqQuoAKkt8pvv4Z5NHSmfVjPJ5dq6JeWDXh/+oKU92nV3eM3K/a60bfYPnO8Ojz+t/U
B+QbVuqMcC66Nm1rTB/8kwkIMxzDkUfPkjfSNv3i2hfW2qPlDS7JTgzTMjiWv44hSkpb/gn+9Z0m
rlWVxaDUSYJXIv/xu/TXqS98QpjrhvkNGj6Cz2bJo2WEbNaAeXiNVPyir/2NWxEJtvGFeM2mX9NO
BFGGNQXLHatwGIKMc7XIejhIRJSM+gPIQd1vNYX86ZHz2Kny+x+Kym2qHz1Ej9xT9wL/1RflM22n
LR5BEAABY7G75k3OWE7yNJVIMbCwZ215iQTJ6n1FppB43Jwl0uoF4kVoic0s5gwoj3cSE3rtNEL9
fj5Vf7eskm3zezi9VBlEhaK3N3eNmrgsE7hQUJKwYjm1aAA5FmcNFvS/4ijDCx98K5CO5PLNU4tn
RPJGV3ksmcLmd+oe26XEa4nqwFTM+rN6lNpIV7QtiNStD2wsWfrcbhLjHyrQ5nlfoYXkghGzKOh3
9LaV6hlrG3Q7gyjWvbh/NmCHplmnHUpSkpuIV5aNhePU/Ik3CkiCPU0ndc+aAtm+Y+0gOoYmJvGp
jiShUQAP+oC0w6ugKSrNLL6ksMpdkigwpg1/gH5LfZs+8svef4SL3mPd2FAN7U1u02ZTAyO47RN8
UymEyS3h7g6x79uPQwFegzrjY0TBIYEPQ8ZS9N5JdENJZ4JJ1eEJFItgvV8yxZRpfqk/ESNbQZj9
DPVKhLENLUrFNz2LMpMHGtzUvXAAhpSTRiqs8dW4zUe39ws1ENIm044AXYw8WMDvzwp85o6ddxtx
iEsR3iRWB9kX5utfWArcUu5Rxq0E3deKRCft/MJAdGVdct/mMt1wrIFZ7EiV9NjIUKY/9Q7Rog30
2labAgTW2CE5aGnVMllYuuLY/USy9dP7HwnQeHYBeUBS3YxmLTcYN8OuEuvRAofAX+iZVLUoqF9f
eH8QK6S8FMutGPlCsw/+rsguAv/pJkt5UlcUZ1egmuNcnyMgMCGpFGGnJO+Cx3NiQrHjGTu6Kfuq
l1DWHSYJwnP7hoZY/sWtj70HlMP5jaH1eUKcItBTM/OOH4yucY/yZE/3o6Nslrl2p7ZbOqwQtmGQ
IK6sDDGnJW9+9nV7l1yPfS8eOdLgmIIf369zERN5RFhd79kAN3Vqg1JhzADJtA3H/88LVMtQRheo
jTqMTDO+Vpo5zrRLkKlzjFs8DJrfUF1Td/oJd5yDx2N3Z60eeuoqqKT0MkW0AQOBwYkifw0Rlfpi
YMJiz1yA8ItOxfcagnXJXT5Hq/PVE2pDYvdpklMDMHcPVi7CdTn07HBNEtZh/S0JiH06WNhLVlg5
O/Xkg8tWjdCI3whIl2aGfCEEJsuLBg7ON6tncVp10jyrKfOO5nQznD0E4Ake1jHibw4qUw9QDwcf
rwwHa2efqMMUBr6GxoAdM9wFLq1SWFsTVNNix0mggsfPurRm6BWZ8B0bJAPydLivSz9bCtkUuX8f
AmaHh7YBVgbWBxVpQ+KZjdMy7BPQkJtK8g8f0uZuM/m6wkogFM1l2BgYgJDFPkx/rRejaBanYvU4
Z+Vr5qsqCBCkbvp/MuckffUMlJMshqg5Z8YvZBR2vGFLwDNdzinEUzp079aMJvR0XmomhpADYom4
Jvkvuo2quAWhMp1OMOCwANSahg1M9FFbq/O1lMxL11Hv+vVvk551b+/ySVRB9brcO01A5HguK+gx
Mk99p0FhIXcv/cc4sCv+Ws0jv3/sh/xXvb9wrx5J/Jyg4rSihXO85VBIwkKr7m1I2r65+rORaSpL
6qVydO2kWYvHvOeWZicAMdFly1dNqXNFxw+z109ElkF+mFgCYst6PBp3AQgWL/lUr6yAshmXk1yZ
yxBaOVifSlFa1ph3/E33aE5XsueWfGvZem3mqonKARFGzV6WaXliWX5IpzVAhjplw8kz4iurlY1h
kAUAw8ej9meSCyw4VY9DBcAzadCY30J3fKHsSSpKL++sM6+QHIBnewRTz3BwheRNBJPGOTLQ8GCY
tt1ELBPX8L+GZuJy7D+8zcIiER18S1wslMzEm3bUtO8u11KOrbRXtODcgP3NXgR5XnuuVvT0QVS7
Feshwwb38sLo0vKPw5X6qqJ+vrfb7IKULtYW9yJfLJj6MyWqspUyaezhV+H2X1x+4pdlvdBkXSSU
qVqLYrSm5IkDDHo2kn9WFUUWrlNtJGUUWzg51zSDn3NiTOHa47YaHvEJuhe+5wbBs1yYNdgaXRwO
8kDSxk8b+lwptBEqYlLWWn/Dg1hHtwXiBDSNLbjSplCidHz6vw7hRoKaw4eFuZ92GwDi4eBfPxHR
7Wyecq0u8KmpbqMG6OUtznkx6V54QUyXkWvCA0uIGHZntGiwETg3znXiXlvA/UkilaRlRQ38lfV3
fD22oqU+jvGpjRGHiSEvpJIAOTb15NxtR5/wJlrHcCibbygDGcLm7XfI7s0Y1RHxln2YeLGlltOc
P5Zf9SRF2H9Wl3iTlCg6QIp8ALTVlSK4pMfdJy9x6y9O8DH/hukUCpqMbeQaJk1FpjPrnyr2VDa+
zip+55JPAP7lEikjsDh+FbbjQT6BfzJq0lh6z65y+MVXyoCm+jn+HsOSkbTRgcuMQ3PkIa97u+fZ
FtNVcdO/Afa/Wq9z+z8UpBOxBuUI7diDd5heP7aHA5opAhvidmFVPmejBJ4XidkNMuAH9cCirNjU
IE+gLQa0S1ZeOvajGiD6BaLyMYMV1pGrRw31/rrrHxv46u0mXiYW1LTMUe65rFX+CSIvVv+UQQ91
bpJ6i6kBzjGq10wYPajgpgXk8X9rcrmDpv4TIX6hVIk0AhSi9N26Hv+35rQy+nWq72+IjMY2Qkxw
7JHzSHCJp3WFLlpkUwcaFm1Gx/JCTSmjScl5rKZjFitpyF5zRiaoBpJb78xyI8K7ph9QPFt95F/y
PItTWHTY1kbMzZ4Ce/sUtHpnhkI0ZXsIufG9Rn6zSObGo8IKFl2iF/evP7jw7Bg/DW4WFXUUPusi
LyoV9IqgA6dswfBH0U4k2pX6PLSzqrwR48yM4+vL6phynEf7vh3EOc4s06VLakIpt2UWgrSbuRaF
jd2d6HAHQuJcIr5aaBzhofXx3om71lPpyJtwHoV6uJio2g7Bw4RShM9JVohj9sGB7SjXpVQVyWek
yJYbg8K4LiwgYm2Z+0zaU91epyjNg4uKsmvtwBJb17DiOHhI8wm57PVzz3m7gNrSitCwZnyC8DWc
/fITQr/aQxzUbhAUJsfFlfgavazjN/D5tmEEFeojyQR0wC6EnCdyuuzsRSXpSdUrf5AB+vHDrnyP
AaVz9lT8IjrvCfwj93boteDcNXfEclQ9a092+vcgfgL7q2ib+mfQSeBb3gAnziKob4yc2hlD2t9s
f1TS+xmGedqgNIQC58isfmBU/NOSMPQaQP1M7QiBmG1MU5OJO2dSkLfcbMPwiFP1l0dWprHSaJ5s
qYK3Vu4IofrRKL046JnVZbl9LmZUiv3rFNDTsvj8+VuhIdae25JDXQIsxpF0CoCEg7Ed/TPWgVZt
lGHFMz0464if22tiV1wVu5xwpfXvxbcVce7vEZkHe/Sc3LmIHLZIcmISsNdUfP3fBUm0wX2IVn9i
hZkO7O6bNOdGltYm7B9yFIgNgnVX3ErF6UYPUU3IWdCKf56C1JgdKQHmdf33E2ektdnN0LYEfunA
4tggb7RqxudMrJDR/QdFAObr4ZJ/51whcdBS460N5eWEsf46Q0T+BmFu2jQWlB2mgS0EL2EENJUQ
UF9E8T5ZSfBwqovkpCDowqtaZaAtaNQKCEZGaFQPNlRoW3hw69n1Frrdzxnk2H7BW4YRN4lKcZuE
FtakL8UP8UFwsa6pp56vQOGFhDNCOqqYZ1h+zrSS0ghalld5mWGjBQNDWm5yXEslQXCxqCDN87XQ
nWblh+ATZQPVxOBD4Ng6Kgj23rXuNS6MeWqXG/g+fnufbMNJhx2s9r/aJwhP5CRta27knzR8FMYN
HlurQwU5QtviIi1IyoAPQlhSdlK3QZnpwXXaG0xml28Rf6vo7ZAPqPUsHlfLBxHAVNA0HE5f6L5W
LmQGV4spGQ5Xhlckno+BfEDXYjvdtMHlgepFr6na8WbRlOH+O7jqrRuwuVbqVOkkzSXeBMU+pOjs
Ff1F9+O02o3WLYmgJXoxhRBktSXYBZVX0SRQmN4KiBerSv5aIsoHT6BFCIGByqu+Kd2+UxnL/g0C
2plRBGayuHJjbNRqOms289bGsfnkKWKERprajKyQ37vYRLByWdb62Va3Hl7TX+B8Rdd6AEDUfiQm
RLTYSuWuV6zbV3JTtZtNrZntDtK+usiqqT5Afn5CpUFeQQ885CZms15VjHeo1LMq4HaedZpWQpWz
oIn6uGUqwzIxUz80ztUj92p+dmYeHmwzr/9wZNR72D9A/qgMrN8oWV1BvaTo6FFzK+DHTBEk6vJw
SRkgVdP6rRPO+2xQJbwxBOrLxg3UtGoHF//QGDOE6aK4cn5tDqJJgd6iY95SMmYvDjSk4UUXrW4f
AQSOLL42isPQndQ8U8RCFr4ftL8hT30xGI6sLNGtu7PjqgFfwZhmw4iX4L9uxwXP48j2Wbd3ER0A
objQc8ub0bS3rxoFsvmLFKUA0TqNzaVQymdqjg9B81OlhE1CGGUDaBBErMnXYUx/8/mLAk5ki1sl
M0f20FGV+FNIotXT5DxRv+LTJPTKDVUtVtBl22HV594RGtppznulzXCyW6AjFtZMeLvdVFPD2tAA
AXjoGusaDJXQYSstbR5sRZgJXL6PDh4jAb274iSd1PD8U8RpvcV0d+4YynGpggeqpnpGz6+kvqOC
WcaAeNEnSbHO7qzIznna+fYAPX6qnRBhZCt696LNzjOUpJCx3Hv5iTWsVR9ki20jHPD1xsE8v7ja
eJiYseOvatneKDEQQQg+7cKaqSBx0/Jr+gtjK0LGh6H8eI6QhTKu5BcNkhd6bXYV8SidKW5co3eq
lDil1P5gI9c5fnEW902Sx8DyCmzWSn3c+kCDcdkcqzB0Pe/Mzb+7w2nhIgcssNdKIX9mGfXST4n9
uopG6QPgw4UJdBjgU0oMTJaowzehMYFl/Eyc9fCOvs2HoQXIDJt6lNf7gWuAtG9CQGZm9IZ0ifFS
ENrxpHw7qrm8z3bo6Om2cfsIsxODyGXtmqUvl19zZX6VZ2YJ1TsMXvpZ6CF+zbj++5tRu+Liyz3Z
0oa7XDR2rhfOe07/zTZfqaltSSp+pd2gZxKfT7j8bU8f/3V2rNaMieDww0Hm2UKGxtMyyWJIvqaL
fuuS7UcRbDiiHYC6cUyni4DSkTZqxmzvM5damIdPFoJ9tbIix4+O0e6MGCrtx3OlJJ8sajm2HzsH
2koOPWGgR5EySKtQrlFMIHujUKgePbPTZjGF3N28JVB393v+TSu7jML2vbO5FA7Fd4cZLkULeNSx
JxFSKgfoB3qss2aE5XhUhybqIKvp//NzdxWIIxdI7lUmvj3flLJo3UAk+C7+XdN3SrwnSn2zJi/b
byRwBtZJLxcy2df+QASE1yPiqWXJZ2ncRvVo7K2Q4Vqxkhm+SB8YEvUdgB/SdiNRfq2V1bbFbTwp
BtuYrMyHCfdqtaloyxBO002ErIrqwVA9APRxOEng7+dViwcN/QG8UGjCM1Y5zt5OfkCCEO67Y+U3
jr1irXFZ9g1oYXSOrmmtMQaUUV4U12kE2iEGP3C0+J5zDnoSW7XrVAmnA5pHdSqiaIVIbxnBd1Jn
7JwZ3eUp+Ck7Pb/0HL79vccwMtNTWUE+92W+BrpyTN59KLkEDQvwkXxS+4JYiO5tOmZ9eih8ols8
nu7+WO7nusy4bHCJlBsxszotS9ZI21eSV2YkYSX2PcIP9yvuTZ+lSerklU3uBe4rBLd9+MtJwRsc
k62fQL4qyGZ7eavZQ6t6SetzfS9HO2czFqBmhNRG8JNWkyhQ9+iO66kxIm+EZFQH/GA9+hxcCgFD
Z/mrfhp+VX9oggyLDEf5/OMes3BEEh7b2IpJ/LwkAjUvtsVmDLdvBAT+Kx/uJKKstif9I+sLjZ65
WbV9+mvfKmXugVSjNet48hreSwF4oJmNUeiXaaJH33GMPOakrUMIIihqNA5e9fb8DTJEfZa83bCX
X7Bzq11hlwh2PbLlKgs6Q4uwfWlbFNh1yv2XBrC99kwUoTgI6ICYfkuJ9C80XFdYHirZ/du8BtEo
DRcFsOey8+gdRa5b0GRt5hJjF8VD9Y/jEcHP6cQsfd/QD0PwctQzxET6/QrC0ejPrPuRoyHRWIZ2
UQWa7P90APXcfZfVMwxM3PHBZLK3xZNXNn5uZbnSTmFjswwtFG44ALaeqFyIEnyNG+jcVx1sGAXM
DLOw+wBSzDqGqYxMuSNThT/7pL5LyH/bGb0E2mBY3pqzC/cY1Icf0VygV4y+J11OkrgKWOOqU4DC
RNOYJUJQAWsTTffb9xocb/U1g+8E4M2Q0k1N9WFb7AY6hWb6+Ru+2sqDkLB7hnyQ4itaSmpOUuZ+
It4Kqk+KKJcPNcKIWJoXLnQo8ot/YKBwiZaFugz3cuPtO8uIZgzLhe2MDpa1uf+m9RPayidb89GP
G0/lFqoz6yIJkLcOTZv02EArQQyIi00PibESnbQ9GIOy4wJMdOMSzdITSeRN/zdg3ZcF3nnKG/1D
hfqcJ0L84C0Z+dFaH6c0xGpY+VSjGvHrHHmeL2ukeF5kI2S4BsuqGvrcKawBOlYqNvSfTr11yALm
OTeEl+X7MN9wHIkbaU6wLaZRdouoIyT3A5f0JDkNgp4GCJUZH5eDXrm+UPPtXwXPnDiToaEO2H1F
MptegKnix8qX4LP574XRsJ93B2+EpkuNHQsJwDHYspwdnYaKKgglfVdDlWMHpJBz3Ank1vf4PFvv
eMyZTZSkyNaBfO4C2qAGj11NrEZGyv/YtolxsnINbSa2+zDBkQjJInhpJGoIGcQGa6hSq9wZ4VkC
SBbBdMWzbYP0KYhNCExUJpXVKW8AwQetEX7YrChQKzeCWV/Dc8nOXFVcRjBbTaiOWu8C2wlsG7FJ
DO2tDnaiP6EMJJaYegK/zMb633MeVu3HWbwHepaQh1p9MnqBC+Bqj84I63ko9T5hKUYh8jdGyQzb
L06q1SoFI4YYbyHcM7xH49yceGIErBpPbRacPVR2pz6oz8fqNyTM7b/3ErAP3X9GPGKuOJZHewcq
+lzn2GuTgU+nd4HiMmmoN5dv63F+YoW6QUqZsy+zAQq4xftLeMWwILYfNYbHcpF+MGdY4B8SzbOF
bHF3BX8oxM8QyKok6ij/nYnvq8Ve84P09I1o9xJUUmUcT5FdOl8xivpZJpLlb7GT9JZDQsQa49MB
3sSsHJbRI/zcjakqbQzjV1SVVkeaKOQ9fE06BSFG2zqCZRr+4Qnupc/OetP7uRUZorugGkJazkc7
8cyVgVRu59bRoujLs6T2Okc/NF6kIO4LN4olJUGGtTBxWctLGqcZSAL1OyixXXzrHy76X7PRDwz4
ScyhBZKJlZTQdfWa6DN0frB+Pkn4gYX//e2kl8ba85JPWSTm59aerRfhVurqa4ASiwi9V81x/WDv
HHvZkvdKbYc+aGL+tZV6JnAeUuwt5XZzAtHXZzzOWJpRA1VKtrbw1v/BnJOy54gtUu/X7S1WMFrV
wqM0bXheagK3EZeBQpzf/oN1a6aw2rC9voyKfagsPlwgHz50kCAV6EGScqoMSdPZ/Kgctn0xHwVs
GEi+HxzdunAeEbJwMjf9rFGwoL0Y5PuyPYzCCj5BVpQRNM2mZMqn5rpmjJ223Zz0xoCx9McwvLRm
271VCjolz/hzQoDRCpm3QXH1LzBUWcI6Apky3nYFuPlZhiQNSXTZIXb4ThofqK3bnQpX4GAQDXUg
3MXNFrehpBRh48DKHUUQ6+lvjJgsu41E/jkoDsdU8gHE6Fmjxqv56zGR34eaHnlftFrpmIOvQo07
L7/PueRLlPYbiWaL/S8iYFCrNQ6L233T2rwY4AB+as0Nbq/KhKn9qE5yWkOsNWAYFYpSLNjYjHUu
t8ZtbLRXJ7KuniFAG8pkBmpYcvyEIq87X2Xv2uxgklYqeiDzSXUk0qrUXHwyvPSx1/kchYUS9i1Z
5C9GES1eGd2GS3iAgylWBz2Y60/TH2FxwVZOi7Yd/B83f0W1YbTphKJ5EBMhMUTinhAfHmWWmD0g
Z+Rbc3FxjovnIjNcCk16iUBXKoN7lVg2ZDtEKpMvbvkGaAhF5ybOynrjgsRXI8VFKCO8OArKF3O+
qSp4XKslxgSJI2hFNMrqQUxL1uKHAdW9PNxZosSjUrwBEMYKvQzWrAtxhT6+ib9L/AMfryIkKGRj
JE/WqpRuozavW/JV+uPJvPOWJFhLQ+tOHzeXl8kX4AU6DbIK0IZvRWyaMrAxjyBD3+JRFOZB1HRw
/v1g5oZ8/OdX5MMxsHHwORvVWvLpBi/JLbL/tkE967QccMaioiSkGanAthZSKCHvCoQEnKRJNGRk
wA+K+nyQm8zpYtg5aKqMnYkQ+ZZm6xTGa02XDBqsbKEjoLJ2QCu7ixR/cd/YxFqgBQpXND8gmf7A
nqObCVphLJrBC2Pfnx/ko/EoW0awXOgogtOcwx8i4qhCvL1+3llozcWCsXEbl+Dm+0LYaWuMouZW
JkZNiQs1WmygYh3plv0IdEzyWUWN4gTfnO/1MyHBI4MBiRbf6oYc8/9K/Xk8Jeeh7iXnZB+goTP5
0ZgmhMLBL807tCEPWmIBeS4FiRHR5JjMjifzpOHDHB+W4FwHYowWo58ygzfDuRkyAC+H6IZrgYgS
0FEWEL1wiDbXVwhJ/EvJm6HGgQjV4llwdaH+BO4m0ngd/ybghUpErStCz07zUhrrSID/7dvMUH2W
+m1/BgeRP+94w+XiSmwC9Ecu/wpDfcX0vaJLgBBwV5vq0qFRohkmTRPbVnR8xjwlI2bAVbkookfd
Tr1JG8dKYHfH532Vg7qNT9WQW6jYe9guKHwoj6oqdJIyKw/TjZJ4Crppp1cgU4095fVBlL7nXboA
3CagWLrrXz/UPxRe1tfdRfzXsR1618MvlX+vEB0+5Q9XVSxQEL4RQaoXLAhUasrXaFzOsrDjBf7e
6UWvlpBKarxmSkj5rdAUtbTC1Ey41+e+DMYyJh/pg0BpF4LNPXA+Ol0y75LfX7xj0KtI0513f0Hz
erSx8cOViRRcowZKO9p57CqgbhHE9BD57ocsF5+iHVeV8UJmerlUd2399rG4sfOc40A99rucCId2
LDCLDqTG51pZCieY/M1gwmFoWgRxJCv2mmb8ioWp8sOGqmI3OChDoP/eqyLCTEwi59XjnHqGMJKa
kFKO3xeBmJ/Ck8VApXTuI3u2dcPfxUanf7vGZLVGjAv0tXZi3alBsy2el3zKF8akzq65UAB/H0ac
jmlGdvmiS7OwZ60KIg1eU8GaGir4o+54RiZiStRddUOD1ftK4acndNTLmo4hiq3VaB3ZJnP6lcCx
LJS6nPMg2igspOTCFAfbTh8ennReyhxMRMjtpCov2vguecJmLiRNCWAbUrJ8W2ZOWp+HrePCK6Ek
kPLrsWde0i5sh+LGZHIyNk4RyR8yvC4J/mGCFssMxHmaHBr62qvSBSUJquU4rYiBhedrZnHzYOcj
FpEG9tG7321itEwTh8fVv+qe/Dupg9KJeZ/ukVa19x635wuQqlVc6CieAcBhZz8HHS3c62Gvq33/
jh7xZY1OkC9eeLPyPEvHyKkiY5fPEAR6fW7/3afl1cUNXIZAaVlJqV3MGHjrC3V3O9STNqCGiIaR
x5fp1PnYwX4F5M4hY/wlxmSZ/JaCBCLUkAnyub/OkaqNPpjRAQhBy040kr30GHYCLPgo+Nu5keh/
63oqSQiikLJJRAg1zvMrRzp1GnGROLc2G70zBROrf4xqcC4F2ikJbp7eatHFcc9caaXF8rgrYLDb
EZmPfQ1Zb3lSvPC+lSZ7Q3aDKKRiey6+bhiPqHPyExgoZfbHcmaOCs/8zJ6EC+Bcr4GeTOFjuRVY
hlIf4FDyJQRi5tzGaiQdeDmGXr1uf0EkzGFwGogz68R3P+ZyMfzvyqEKNX82iEk8Suh2AoURm0/a
oTYICz+O522Zu1A++7R/ZSGXpeoaymkrnY8Zm/+hFBXKa9qj8ttBRLdI0RU2yS6i80KzPLL2Y4iV
WQI8JnHOhg1jhmFPf6u6lP2pgOxkrlgqOrij8UlOCaMKoV9HgtkJBLdB4SLA5grF6TfPFimo6GEr
Z/lwBnuro8Ezn7kvQP8/mSie+Fx2Ceo/IfTr4S64REcupdHFweMTcBW0Dk4ULrsraNZW0LZuIBW5
PmHv9xOACmDMgvlW4x4YevXQGoxvhUWc8Ppm14ON+ZQmvGuShO7kjTT1eVARhPWkzaS6JzRhvAQh
LYwN3PZSc2t+BY08ONDM4ijwpWR5sceC6tvjQ20jVXFC6sO6DSH0ptB0k1I0i3CFgOyL5/KpZp2B
yPomCQ07iPu25cg50hqOZ8Hc6sA3p2Z0G+QJ5ORW/03+cgS/6RVHSCZgVFTw+TKMRsNfCbeRs3ur
rc3FtklTBOZX9j7h4uoVLPVv0hI1ZJ7lrDW1eQ+W1ed6JM3FOZ+sp0Yl/xUxuMp/CgHOUmUuNMDV
b5uxy2uwZu+oILUHgAsWB/H2A1sAyYiv9BLRU6krY4C8/JrpFWins+7QSoxl5ZBgp0MbxB1sbSH+
8PMyJ0xDvbUaZ2meUxsjAkpE7/7AnZstPAJ48l1UmwVVotGmT97PGy7Q8wqM6cvnAl8a/2KYrv6V
ESqA0xBwzNcHA4s8gChvVXUMguvmr1uOKW1KVVqoaCs2Rd5Iddwi6zUXcFUvaqcEUTvLkaiWKhi3
b0yf/3CU2h5TS9wMWz/9Nl8hfc0LtllRU7A4xOcCU6y7bkbXtHQqYGPzD12eA0BoL9pdDabe2HbZ
9gLbW8LN5Jg+MTHXfG6gqo9O+UihMbP06HUqVdhMMMsvZeZHyP21eDReTnaceZO2ECDyTGOL2D58
myeeJSmphHWJj6RKKxLBWjrwyAVXIm2U1ib1rqFO0FcYUOhFLB9rGy2Uf8rm5PuEv123x9Ko0MlD
MwJATa9CTavcCvgD9L8tjOsE8s3atTzbQw5GVkrzvValQkShaVmxAX7SElJkxXsTWfo+8rSAkM9i
RvekMISFDts9H6J8QZG68ycaz7t6hIVxljcIgK26Wal6k8vJgj+P5I/bGlsN1G/+HulKFSiT7ITc
Nm+J5QNpYFNNYBdv1QiMbKJMbFekjy2zsAGeckuBl2eUQhHXTsoaBkyJml3seVul/xgCryEyBkKt
c22KBmujMimsE/1yJzgqyL/lF76o7UVddl4amqAQUcW4fnGX6kwFSyz/DrAn7k7Tok2DuXuuAqKj
ivGONRIq3EL1Xs+sMXXsIOl9TSw2r3+JGUuBa07sgAeZZonMeCkbHftaduGE7xYKlTAPuwnhl0h1
dLztZI8T/Az2Rncrf/vJLMNmoF4cy1wUzRVtkjMoL/hCxkTYI4p6Ryu4X4C0pHYR1se8ijP+Ezcz
Yz+3h5XgRZtl+H/o/nFVoiaiI3uypxEny/Ymlqk+ibEeEPTMfJZbxJsfE0cOFO1m2mZlRuAqp+vM
SXhQIpDbup/k3N2lZ+MAoYoHqydog+xGoDisZwvuoV42FAVCzKRRKMDgp+MwsXL2KebIerfpKedu
EYZaA7P/KVoMUP/tfdQj2nxNthHvIF1muXSZYFGsYkpPzwICZF6rA2Y/Ba+ZuZ0lAZi42Wtt9lrz
Oe+ksOvYDUI/1u3s89ebiiDJj7gkRuFZlA062YAr8tPvN3T7wGE7BnFpcYBPFBXppl79LIEJDlyt
EAQeov4DhGTE9asJ6vWpLnHJdeknxtRI2mATyJvZiyCJjHO2Wc3c5JPpYWAzsVSiBJmEHaAMCeXS
uxfO6S37MxAE7s8oC2jbtPqz0P3s9z17qT1HnYA5oT5kOM2SPJmQaBNThmT/7pvR91sgVNf5Lbv7
yW1QDhHLWb0DG5MMdGf1MzwK9AThrZ3fnJ5LgO7kq11zD3JX2U25TCnS5Libtk8ifjI6CNaW10ho
FPBx0SfbRvHwI38aOIoZ3ZKuuOshOSwxff79+2w4TgQo53KFR1qQbn5k/KX9aWa8OKSR31AwpK69
riSHkmwIEfXTMQ4+ONn8Cx7l3+hqDSXD/eJio4/6FinwBqTqbMrv0WBLOk39U+cBwCS/Inl3hkSe
k6QELI1L8j9ybMs3cm96cs4bhUBxKcOUKu/lWNAvHUyZ0klqaAiTnN08bIr/MO9TpCW3yBcuPFsS
xcFOG4UPYsHm1lIpgV0SOFM6DfompaI4cWw8wxDI0WZPK4nPcLAkVagqv4sX8wKdRMKEW4IftCkp
az6wUB+MmGRThMrtYMagJkmNiZiH9rnisgU2jgG/oKmPrkknk4QBD7Utix9otBKdqaxyMuMYREVe
yLLXmNa2Ri+sYecYlCn1Zjm7kHhPjVCb+JqtZqpW2HtBQTL2aMSI9OW1D1HihE949+NVgdwIV6mw
fyWz18vem186HV8buHs/FKiFdMD3gjAGcwjlkTExt/GNNOOEreo1idpRJaOB/NUeWPNFmxkxNvQd
Ox+OhwITyxPsURXmr1VMZ+xF8jt6y4QZlDoZ0YnL+h3OAdbaLT3CQgpN35LdQNrpHg7Aes2zhiHM
Gx9xQY50Ac79N8pTQIEvfP/ELG9lEO5MFdWtBKKQSz4eSIvbWL5QT7iOQYYM6MGAjWgbt8vkHl8a
9KFD8I5rLt4F7FEZy9QsFmHWTb442yncRNbAH5VYoso/ePWu2NKRLHrRApfnzKVn8v3l5jLBmDsE
nQ+AxCm6xPZIphjeHvJZ846C0HdT5+AHwnW3Ea5rLyQv+MgaX5sTY14SUNQGxYKej+scMwjHebUj
xgIeU3TPSavd90bUbjEAljMXPBdnrWH/BrI+Knmtga6M6idzMbXf4u+j6/9mCmy8ez3J9ntiMGMs
uc+fSi4czd/XYhN6cOSgdG+AUoVII5ytObCaNoXUYfZYoc2oIRPg41GqEH/fDXacRoZkZlKVkVfE
i8HsqEG3DMpZB3iEL+pkN78ID7/W2+gLs05L85nNQnENTpBR0DG/1zjPNubiyW8poR6hz3CfzAP2
GoCCWWZrMNAXq3ZKx4nqjtqsBmIoAuG1z3vD03xM/3RRg8vmVmBX7WRDbkK84HeGAHm7UoRRhQfi
A2s1b2mYl2DYHX2blOTaqRuicAt81yFHQK4xhDdPvQl6JAErBPo4fQtWFXskt5zSCTZi+h6GTXDS
jdamf/b+HSXZdxmMkIGdvFQRQeAe5zTkDADn+jqLpgA6b5pNBkrLEL2q6A+CadMWqmrpl5zfbll5
w8KVM4PeqMRUx6763Bwa/xCo/N+GMT4lG7CSxm2+6AJj8wxwfl+BqFZ5ArBHTyqE/5SESPbFzy6v
KmBIXA5uFd3ueGWiH0julI8SSofvNev17vGcPofmeP+2xNO7rqVQnusoyYJ5bE3n6j9GFlQKzzVC
DZQh/SbOVLxsRpxuzNLl8YUNez/mVw/sd1haejKL9Sv2ZJGvxuopNwoz+JesievUdBsMJeTE8h91
bNzF9yciNuwlOwvYylwqKTnXQEzSV+4ztbEVNivcKNWEcARn3VCzvkMtirNNxWQIzK32zKAF6EZ6
Um9DX6CsMJAAfC4uEf2vWMzSIoe3JJBaATr//xrck8wcHhhCAmb4hwePujz7NSwmabCA+hRvj6Pp
O2yt1oxHcS/wEbkcIPQ23Nc2VjAHVYlU+MFlivzmQTGRBHwqhRGmotatOh0gPIY6SbHRLylcrPWs
8TLzsObrRsiGKk1+3/gbMJfvwu66ANhvD5FSG1zLSPN03h5fxvXb3DRW5de7OWAW+wulBsm/TbeS
1aEEHTO/sHnJ/tL9XMv61iEPMsoRSipx0EnOpKsLFURf2KHiWQbkdpxAe5/1hmOimxBqMRkyti/0
q/XKR9lAjDsrCp0tbt2GMpK1BXhsPx8qT2FwD8QkVD8g/eLIABDFH/DqdOYynu6qUVZXwoBwXiXq
aLEfR2EYnxeve5TN+eqXNFseC3WT+RpVmubNTkJZ/lykQ+dz2tHbDEuPCJ0C1QdbbeM405dfID77
FwePhKVYp4iRWZYekN1YXMFQCM+3RWMq0O7C5t9ewlvdAoTk8Bbnv7Ojst+wcXWwvmE4taFl0rmE
lHElfG+M3dtGbASdIWwzV4w3MTO4k7rkfKUCAAdQUyFehV6D98QBr2t/LsuKz+I1/h6NR9XR6sEQ
y1pjrh8o16t70qPpUHqYKY/E1lkcGUP2QYVQdIoYx8tfPZMUjS2AtQFAoh7B7MtiPemy3UuaKIdY
QPX80To2n4sW0dxTYKdqnOZy53kC/REMbC8TE/2qz5nbmkMPGsTciChWriPpKLHhRPpw6Rhq3YQ4
YRUkh4ugZGQlBrzfbLDOyxZRPIOBBJzgz6UWTLhaSfK5MTTnfnDoW4o0O6IGJYsotiicuA7fAXe7
rYYoNv6jQlgrquZEqgNHqAMmNxbvIU0iiK4XuNqoQYrdR0idivLmWU8Pj1nhr6jBMPoS7bH+ZBrR
JT2Pgv6wvhGLcPleBjDO7AKkk6n2oCqpvILj2GUIo1x45XGS27IwL3tPaVPPEznEEe0CdPPiYFuj
b9+/NklV0E7LHIDEVhjBymwNTdN33o9WXKQG6SZ+L7Sf+kYFojawu/72Gq9NFUzcoRhLAUvE+2nz
rwsl6QMixc5LxmjTfQYKRrTQ8T4Gbo4KZ7M8JDG1Xel6Phi3EMJuJc2ftrcYDh/VC3DfJTo8zzfN
5UfOcrCAthOJTQqJWS2Hous=
`protect end_protected

