

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Gub1VXq/9my70IMNYnI+loF5VZ7ee86ZBpAGzL5j+jwLQfPXAWQ9vuaGimuQWfCvI177d9QCmrcK
lRbHtdPXqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XCHJyRkscuJOpjxAlpPvd15b2tV4+cleGX5HVVJ/2Y6XWbVNSZsCQSUsTkLA7IyKge516I1wj3zW
vSbDpitOXWUELSO5CG6d5r8ZVemvSn2BJybpLquf/4fVeS1c+edRHNf6tkj5Q4P0LsQat4mBIGGY
5hCeyo5aPtqLWGIyMEw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RqwoFbaHoCNWZ4v1HvZQji+hXgCjT1Fmm8RnwPGBKk3/N74/TfbSFLeQsQ92UsPWvT9gifFKCg1j
7eGei0ot9ncWAfgeoFsw2zoynofNtXpuT/2o69ZZvCyc9OMmSHilEDslciAlUOrRZtsCwGDHNVP2
rJ/b+v8vvCejKLtIXh5C95/DXV+eEcsjEVRpSeKGeZ1MtzbV+fZPJnRzoH2U025UhnP55OgE68T/
nVfgRgkiVFm7ZUA/Q4uTOx27LPbQmDFQ6plepnrYm3dIFbr3WOiv7AWG29Y9MZiC/1j4MvPp1qqq
xE8dCNkJmOz9uD4DUQoSIb5VP26bf6BmGLvFDw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uV7zzv9Zx+u216Ml06an9UEqL4ajf0AMjc1K2s6n9qbyEnUVTSm6yFZ0M/IFYGglaG6jdDDlz4rd
W4zdLmcu66F6EUQtwXBmHtk4+/Am3fKB3kIu6GlcyUoJhx3DF0omCc81HS8JxypUZEAxz3C538KP
dZmq/6pOZleIRCziFs8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c2sM3Lkice55qsGCUzeim6Qm2yWa4rXMhx0Gil9+l1mRl06adQHebvNeaVnD5l4UfTgDiNRnixMg
t4I3MixM5k+/dqMphg9yh9uQH4HJHJ6CTIPJ7b0uq0QUv2e+GjaxWZa47ZVWMUHJwpscHTsz0hs5
a4sgfCiRr4cQxV9i8u9cWFqcZ4eu+RYLEbH+mYK06INaK4Fg1vBkwveCaGhKFtvHtOBXP2o42BPE
2i+HCKN5sLyGLlDI9h2MogiDBJsNAtjJ9geF4nPG0e4nijR/pyFXErJCeKppN9041em95AkpK0CN
GYWuH0jkznlTfi9EHnlKl7cj5ibz763zI0uZLA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10784)
`protect data_block
bxIlrVHqB8h7WVcBZuxcUEXud6LMDtwbGwMLCtnnMR31vCLzsFb6HrfnS/QkHnkMlolhVOvhq6/4
5Jz4HktfGSPeQI4ViMbR6gJ0vZDZTiF1NWx4EuUnKHsYYZq0m5rVRR4qS4qIlsVQ1GIm14Z6VZql
JCeAlgHsgtJZ1LYse6Iv1Km0O+KK/1JdZUcNw+JPHg5P0XK2jWqYk2LmtD7EtPzDMtJK7iYWImrs
PYGHejZ8lF/buCZBkPfpsKwsAMluX9srXIwYL6BzGiXzhlLNLQDAoIvqmgsBD1vgDa6MgtVR3ngW
sfWPKRi1zHqKHDKLBIScd/HBmudunhqvwRsXo8IM7pvJV5NvMeigcvGcQ38ow0MzZ8wBUCA2DNo+
GLyBJcfTbtXIxzO76wqI85hdByydnbsodWfZd5+qQlcCJsHdta4qJ97U3/gG5vlKxeQYE3QXu3qE
dQWZvwGErjoMbvpI6nIUnAFB89g52Tgq72LyyGa+KM19zsDc+9ECczyk1+eVS29/bVsBNavks8eN
vRNb4XNme/4mUIRJXMH3wJClKw40NqeIemsNlZ7Q7gpDVJdsLoO0vQZnBnSdgYcELvOQhMHO9CYJ
jbc+2QIaojvxPjkV8paJsDWX2QmiMIKC0X8FbOfGEA8KtlQ7iHbavIyPOuNmBpb/s2nuyKNTzbpo
OZACekIazGG6dKCtOMRxgdKKKP2cPFstD1Qm9eeqBPWmWWgWioBSTfo4fJVmv7GoqZ0PJt8f+oVW
w8yOv/tcOUuYaqS2+pLyEb5XJkJQe1CJ59mfmPrZmN0ZT9niFatMxwrNoTA/7mhCcSKYwfKtxo1A
6ON8Cf+MHHhS0lZHlJ/4GMBnafMj/GG3NecruC8qgTgb6/EEj4WJTd+YUfTIgiQGZsDqbtONpoO6
NRZjkSFOaYQa/b+DknGknY7f9Xl6gecbB2+cDwX2EZGqQ0MLpZrG1zu9AueytHq6xxYvYLJBWaUX
pCY7/nrt5YqunR1NZk5Hw0w2fxTBTJMmOYNTiOkNA1cUoiH8p8TAkDU81COdlwxE3J1U7Y5J/xpI
S8dXzNNvkR6mLRRTkVHgMayiySxAD8Mdgem6gwJjCI8916uevVL15u7p8TvmoGTPlcQm5KE1vl4y
kzxwiWaM4SUrJHj1WjRJVufqPD0atcmATT92PskzQjFEf04w4iLxr8U2E6YyiDa0aRiAMTvJftWf
7B8MM/jwGVJcprJFLZYVb+U6PXbdyUtnbbyLXkRH1la4IjcMRlGjhJqi4niQ9GWkw2riuVpnOJuw
WZWpW2BOjMiLghMEc7VY2HF7geBDezf7EUEuaJG28+qK1pyQIpYYUEibL59C1RpS9lC1XJpLw8xD
hZLN7uVLrczK/J2lsdmKIJvQXDY4tk7N3UqcpmlxODMY+S7OEkay3/+n/KzH7wLFVJtlGyhSzsLQ
IF1cLYsF2HHq8u/fNtommv86gut3oKPSdo5KSr9Sf6gCxtwtRIp2FaQ1JHyoq0l1Z1WfZewtHzAo
5e8QolzuLKpxGgggGjt3Av+vWZ9Qv9oRDFgKdRLptmDVg8W8a0l91laK02eZvnGrGSO2mEko5X8k
+jdms40e3lz1zOxbw3RVnywAT0Lx7TkAs4mNceKLtw4lmtnVvJmjl8+S46DLXjMzzcdVll5MFTXi
w8wKrWzxlYD21NIFXziB/LejLNdHOlZJNbmJ/UzgoouFoxSSjNA53fFlt2mSeWX7aYwSdIJWkhte
zwtkmPhivBFF90WOEfAu7T5w0h2sp18BWga/AeZW8MWZSNClgvzANtgBYPQ592NAC9jXGzC4y8dv
9/avVcKC2YWtStW3L/PwjEg85XHh9mjCkAGWRyERNoS4Agc1RYCcG6Hjv91Qw7q48pZuEx106wPk
5HXXRFMo4BOYcXNX+05O9gqJs04MjqLMEuiJSTZMeD6a6ddH7nl8gjc9ufzVoyI6D/MAJPRCKvWM
W2StpuRCE8Q1crlv4i34Qp5tLcs5//a9bEyYU8Og7/KNjNr7bQIoeoNW3rmJZN/RY4T2ZmfS86VU
NV96k/gWqN0MjtRUugWJQd1oApl+XBLddmmUDL2xACBU5FYIGXRsSPeXQuAKN6TAQAOkEf56AVye
aq00wpL5IPVm5/r/JqCMjUF9NgSVQwt1Yja93rFortsE5JxRt5r5NGQBUaZxXx9fLuILBEYxG2EC
DDm+Kl5m21MpVV+Z7lCYJk1DyaqUs/zvjK/wQOUK91JMTHaYggyNDkpJRG1ezTiGcPt2EmVILaRy
aKBSfvrR+WUmQyqZMbdOBjjuYOjMvp0UM7ixHR10kH+wXxnzmDUuJqYaKBbVMyxNGN8bggPQBMrd
nW+xUAdWrvuV9sZ0Yb55rCfJYDe7Wk97YMNKwxEPVKZ4sLD8eheKh3JzIuKhp0eqSuxBT1+0nw6N
7sEnWaf9HbWOiWeYsHSKh66LWfpJ6Dyu6ms5BjhxufCBJ60G67wbQRGdPyMPMopJk5jcbYKcv+nw
zPhq4i1IXVbyyV5RQHAOrI4rofXy2k9t/23PJ1eptzU04+03rriKggWDGPiaMkiw5t310BPSit7C
/s2DoN6fk7KTHDVJ7/eZHG0yhGRy6NjAla/tKzPp8XUy1R93kN29Dk98WwIbaQvUJ7MpJplXnD99
aLkfxeycRwHhBaZVAvdRvnxCcpYC4pmb3946MPdDuPZC9PvBJD2Df4xAFBaBmapxyXjxQEYhumGk
+Nw52iKgq71GlYMMs5Eqvpk6lA9uuiyEF2WFmgFOnk/KoBjN4yoBVh9ig7k150FexWQXOyBHWQ0E
c9cHmnzmBh5eS7xef1G6bzOE/YzuMOZuWkHOdxcTJTC29HFuDBzjlMdmuJ/XGjCgM6ZWJVzr6Muh
8KW8RTZjUBNyciIY2FqqLEY+qLTsFLjTRqncMEYFuNGuzcXSfpMUYMik6LiBr9uOryqFpRZkh5u0
VvNhu8QHyIxx6lVWC+/51vzSNMmYj0XiBNYM5UEFq7c5iSK3XIFxq01BUiNSfZmPKzqpafzl6Ol6
9cdm5FDBuSRDnbByCR8+UHUzVGzpfN09/9/9eqAd/41H0E035+sGoP36MZmDs6eBbZ+ehfiurd95
Bso3DL5Ovq/vG7VRbR7JkrGw4hR/Y75iOB0CACnOHrLquCJlyW9oow2bRf7ZrnS8wWD3wN2OaXqw
9qaTrpcrkyaAUt0xH+pFLsinEbhhSQBPzAoaujG5xzz+MTW9qYJtjT7Bd0tCdvZ7U8ktMBkxWT3j
wMDviMWT6HqUj4egG4CVIHPkaJAgbYjj1gGxfbfGTAaFqeFShuz9t9F0L9ugM5tcvZDHEkPRmt2E
U0pXyRiIQA1G0oaR8YzmaGtkaE/XeJu1ER6zIoblpJncu61bWF2EJlN+7RuDbHe/qmyyq7cvIzVo
C4Bktie0BRyhX7x9fgdWaBhpErh6FL4PnxWtiPcL4Uqq9Kpoyy0OY4OvDa5SiQmTnKts8UtsdGGD
UpQfdiQJl5OeLJaIts1jXvzqx/wfT0fGVeGa0zIxFdaHiF4qI+fJsyH/q8HfddeHzTeKzMTnnVyj
LTep1EHFL6/bO16zhnGmlNEgJYJ7NXHf35dx/AQp9VYiXZgZVMZU+v8cmjIFEPpKJUc/mDw+BPem
ylbryY5I+aYBtHRRp8TgU/fOiMCxfuO/vowiRp3eEPc5FnE/L4hXBGtrmkzdYidAYfouctCITVPl
we12+XY8T2TM2LIVk7BjndTCEnQ3YJ6Lmn/gADNItD4dqC2H+dO6yLgqADkTFGr8EEUg7T68/LE9
0s/m6CZeH1U+xYjxQE0YHGR7M+te8oBxatQND3AOBHyjzkrjg2cn6DEb4of7tpnubSDRQVFzcymI
h9wIzSppJ2CXfx9SGdjf1/aUffR/J6/WvqvSUuhHG10ui7PMUN0ZXgRi0HwincSXHF0tyJ83dwgN
SvrT0Vl3hNaytXrkqsCuFTug0K2z/mR/Y3Xj9NwBFFEGnd1a2CD75gem7YLyKdwvc58sfJwympjH
UodGdevUHqZTokWdfGExNddW1xSPnyil3aWp+7cyMDoZnjl14p5vQWy8HM4JVZUdi++3BAhvBeFh
PkG9SNFphde5vL9Y6jWMM/jkvjYRyfP+95PxCutr56iWWqS4ydXjWOKp6dNJccTZgVeUNBcUWGew
VE5XpcYwqYnIY2F6/k5T6bQYTVWaHR5UK/j1Kk8VYl+SecnDyouc3/4pAmbFHPd0hlhB781sEmUb
yLpNklDoVUwBU+m6aWYOB7kHFSm/HugizW0PDS1WFmg87ZLwudsaFVJ7xgTa5PMMttX0gokPpCOm
e9ZF9ptCPrlVuYiXcxG9l068I05gmYP0tOV3kxnESCG2/rtB2uPQ25miPk0q2keFDOoyrkRE86my
jWN5TeiGc9t+XrWjI3qCHDCB4JHZI2kRhvTMVK9A3p3/YrrUUb8lLUmlu86bxXTfTGFiKT5SAgyo
OwxWnfTMg2ft3U290cxINm/BTNKqYpg+kXuARwKBSdBVXmY9m+4lyi8WKlbj0BoWME9dcD5sTSrw
EkIel1ZFWITENVU5RzxmPlWXxPJ97G1H64RJ6M9GHJSmqLDo3Kg27XT66E5ip7XVwDUAwb/rWcIe
aZrTlGWxYD4HChdfCbCwT3V57y1aPDvFgfvSkBDxZQJne2/Haln86PIG7kOYS8qWgyuYnW6U3vIK
lrRjhhRixYS1olX3R0ON7FqnyaRt43QCm+opR7mokhFbsQIOvpOHWPwTjMMUlrPw448CbHLZ1dJq
6ipdLjYpp6LfrBm9FkEh3KMgrfKZQX3CBkSTp57wC7nCa6pPU4CcTC9G859wHm9AcrG4nOhNaio9
byOuCyTa8iQ4mneXTIgQPJK4plIftCmUDNftbOBpmiGDgTNf7qkZppjM1cfwmjAu1RjzV7e+Ulu1
uQYXhRoTTosfKk+tZMFiARmGgsY0j8zj20wLQ4bPh96T58/TDjBfT8Bw66Jc4o5Xj9ng+PZ23k3q
DIOoplGHl7RFvKsDUDS77rVgCCBH6h3XnKtujrSpTqXYzMxdDs+5CePllJZefp+EYO8jayf71TeO
E+uLax5iJVhyf83ONn1FVLxnzOW9C+VhmP5b47abAeYTzdbzK06aScjQtxnsF7Z51YbwmpiGAh01
+ZIkYmNHpfyOlGckmK/pD8HM+BxZblRW+SreoxPvpHmBmIpV2ZjU1HMWRWPKkJYCuyWzPCAw3UvW
VDGiuWrKHAXhKhbNW/I8qNREtk7gYllh1s3hi4Je/dovq/maRboHhMGjNLsG/vKmZpuZCib1xu3J
YjKe6seLIb5m72fluMHMIdRtWzoZmp8kXpMSsLJCaDmxfXfu7+splLmDSWa6qXSfAOtcbtwAltKl
6wvUmNDozSy+ed/t3soFWpCbe/jb2zLRgWfOXyEjbi5EwKLUviVELgxVWQV36WjCdleJwXZkViWJ
V8MbhPqV8sSMe5IG8h/nVJWFfFEeJYlKrt5RnvGHjYJhW97WLtblG6ZkKEOF7NvB20uYrluiE6CM
KAs/Z7Zp6AUVc2+9YAjbr+XnjlOXIUBB+LtPgoR82/x8V5Y4rgTC9YHIG27FM876E91zUytxNfnf
239RlJIj7ICpznPB0A/+eVYHkPRkKYnFrfiG8MTZlHvIhiIF6l84XJ4nbb4G7YftYCsUOg2tcrv3
M4EBEry217B2jZZvejwMsk1+f5vbyU3/1PVkRtqFZbuHGQGgpdbqmQCNX3OBYflDLh2+TnjbzFe5
mjIdy0ogRjrD9nKOz4wK5szf9CH+GfnH+oi9uIFijNITR9tdL1hjW9Nf0sR+bbH1voGZc4KczSU2
pMxD66k60lC3H+KdxDh3bGz9sqfIEPGLRZuRWozcEX675RqMC3qPd2isGECkUsFLXEb9GNtD8j+E
Ohvd5QhN+ypE0bmyc1qIJz6W+ze2/KdNGgU9CdpHiN77nO7jgKMTQFuVwfXVTnV/szjEJH7sS/PU
AiJjq1ZhneeTm+uSBGiexAuB7buV54oToQw9OSR4cgDXB7pohEF723RxnTk5zVId6DjV8JPGFv+i
PKTpzKNe9SseX7OkuD+bDkaEAg02nRrBQo6rsUpwjOxIPgeJwogRtOn3NDZZALkVtOOqVe/6HIHK
Wjxf+cPHngZUAIAuMdVqcsZf6Xaq2MvAUdggFw5pVDSXdwtAc/KuftC1P30PeufbEkWsJpVYJB7m
7kObvZ+uckVm09TAI2XJXGJFy+xfqZYFPfAy01JU4+LC0kOcKGE2AXAJMrYY3HqudWQeDefevHWf
J1hisy37hG9l4TijjSF3VaRdeCRMADhsCk/qDqbxm7f5M9Rhizgn4UPFuSNArlTOBtI52URSny7l
LWSf31aeTXHQTeQRvr+17e4LaH4y8Hi2Yp4nP7uC8Uh5tR0ElcE52DXINiMIG0G4t60PNfv2Qv61
LgyvhNkjh+LCPf1KLatBgCokHRBehnvJ/BVVc/x68QEBKUPmSpwcDqPbU3tl6OD5GXVtUzsM7gIt
w7wJ5EtCheg9dCFkiYZgdG81Wsbjo57Jvos+Odk+72v6lBcex8Kp1tXU4Bck9XaFfxNp+nNO9bxy
BVe8YU6vjmULTZhD6nNfk0NTQfDqsftaGLtLT9r58MasFsT3BYCvjFW0i/lgp0N2PXKZJNmxi5eN
TEaykywJ7LwdgzyPzMppPcLX1w0JYsMvq2Mlz1u6yTUt/qmG5Bmzpe+UMvmGsd97oYr3LpdQZ4iP
XUCgA++g1s0iJkU5KCBmoJ2J5+mAaXh7mfi9Cn7VF7Ne3QvjNLWvaiMcWH7ruiALVZnoXCcctoR0
ztrtl/s3xdmq4NqlMaNU+PZR4zw8+ue0n5n1yRDuJGmGiuy+Z5T/6F+iH1sFNqFG5ovrTV6hNNPm
Zvzi4tijr2nNcKvz/2HGjMF79A87EqiBG0mPpLb/1OlwE6E1y9cTHWu86UUA7aoah7kXKBjpRtR/
48Lxm6MJir3zutYbiCFpPTxemh3AH5/058s5Y7GH7LDg6B3RqQ4kzl4+ofBo23WlbvLP6M9pXRLg
q+mNBRNs/y+uFnHY1w2QqkZIhUK0oVuffMHfjuVqplvsr/8vNbLtQvnI4DU7Zz1AZuutMPy+japT
HGNI7TGpw26XIq/I6ju2vihNF4a8V9kHOxIs1Fn79JcyGWTlZsa5vlKNVlEhVvVnk/humxV25dTu
Ka7OGQ4CPmlw0o8UVGZxR/YrIBqMlnNAsJlEcB3WrSO2DUzGWW9/eIO6QwE/6ajcaxmPLmvSMKok
Ff5y8BeRTuvhkWcLHvTmOgL1qt1++FAtmQDn93Sz9pZ87+PCH2b+vUfWKZet1NNi1Xt/BxQz9O+a
MA8h9iJJbL6FZP/BtSYLqylvxruHWDYgDq9zYtq44k2o9l3iA9I/SZviOJxgOP1KTCGJYLYtmjuF
J7p272MK7o2I4OW9Z4u/3Zr6+iG4MclCNfAZtrJSTkxfYRsBgJNhKv5zYykKWw+droKulEZPn8Hd
wYPLubpO91q8J8T7AdUwRkOSy1x5eW+fp1z79CPj6aztzQH5GBhj0wChZ0Ny4LJKAxHPbeodt19A
uWFCazUPLLAvYs0y4onsZMVFR0QiK6qWogsG8hpdW2D7M23n9ARXo/RBHdDzOMkbejXao1hp8Jm+
dd3NJeFEoMlctDcluXniBxzj+vIWS57ZBifNhUTy6X7ed1x/RdDhvflLdDcWm9Knn0DJB1YbDAx0
sAxV9E6yeoiIq9gzbb6PVTJHObEVNY4BC+mUu2LZylWmLzNmu5lmn5pxDRB8TT2H7Y5WjvIWBvQL
Z8IDcrxPrtvMiXnB9I6oSvzmegukgQEOFYwKSfX8qS5vUk/G0rjX1RNwG5yTkCY3T2+IGUV+lwY2
y0ZSeT1szrmCgsI+boVfNJ9WWJi3wHIjh4KGQJhMUFUmrWSh7WfBTQ3Hx7doy1Utc6sFj554dHj4
k/AMq/QYvyQpMk0UNLsTgtaoLlPiBthF3ucxMxwJExNR8tewvNpfGcEUFZJ3T5WmmR4RVR0B7kIZ
yuIuvYNCYkZQKxAWiNzs9CHiOwlaFhomH3RkwOkVoQ7l1Ch84YykqXA+dnFwH7q2b7VA1JZdJFau
HlIVCPFO+m9Vr27JYJ+HYMj5tg1sseZ5qU8SEhMBFOJUSitnNKi0LkUUyXGVwSQ0sBUp9h8I6B9/
qBeQhUiJbMCTrMbM21/R2KVg8sgvz6CougWGTaReQXfe+8deQPrXR+5B39Ubsfjlc1FeJyKXoox+
dqPgUuW5HQi9OLpd7qoE3K+1cHMaobfBjdu/BcxGXwVeWrlC1ChhK6ximBXIACpvvN/TK4Gdi25X
DjzmHLqiEm9vFVTKemicCBbwB6iyfe7Hq4ZaFnuedbZtPh/fP5EN3V+6qgKRPgeIslZoBS9BnJUI
6MFQUuUsGwuufwey+EQNEuzhjTdmxa0fariyxNNuoOvNNvw51D24ZDXc3xeu18TksvTyULGdiDxC
wfRc8/de8pxdI5xNqCux+hHSc7fXUdK7ipka3qcGqhpiCoaeYRv9bvA5Oa/7O0x0iuBHqgybx7gR
g38bGuuZRN+f+qpUXMIsy6xighb0QhLyCgq7pw8CNHiwqh/TTnfzupX1S0cNGWN8E7ic5f9e6pg1
PSyHlZ9m43+M3zNkJDGLGpJ9RpfqnOvzrM3+x8974vp+JEgrbT6//Qnjysvpb+YPV/vTy7mIrn6L
OzgsTc7UjJueVXAYpiNPdSj+u04pUzk9SfoMVCR+fP//bsoZk/xWjlPRLH5CCj0hwM8l6HVRi+3O
v+RSv7gjaN/1VO10CPezjN3tA6zC4yii+fqKY+QQZMnFU6dAxa4gq9fAuiKcreW/6yisVnqkTvpF
VrxjXQliAhADNgbom7yCn2VODRCGaWSMz+tpPDdWg5v755mdIhK5ZN9rv2mLmPqFeNlomT8cSiGl
82SPAFVEpdRmmMUQgKRIi0gsVkQM5STPoAmP5R4EHRz9onPh1YjZ9m5uZwktcTFtxCmXmjzxWpwE
vyxuiJiU1f0M3odrc4TQmnAHxFJnJyI7iPdNmW/9ZDCFb8iVRzJLnESCVho5Bv2Gt00ygMFwvMHm
V9ulsEjomKA9s6cfVxycgFzOOASeqSYvrqmcYGt6Q5SWp6Y3I7t3KCCwm60H776/pFFLonz1Qzvr
16Ah3MWeHsy2lCMn9mWTem4VkkwV7Jo5ejHyOH1/AU2+vLPA2XMMm+1wzDMGPp94wRaPJup7uYmo
15ggwA8/Ry+Sg9rqTUvu4Y9aYNUlFZBLH+tWQZm4w+KXAMoaQMJgXndA/6UjyPrjNplgjBPMRwj1
by5XtW3M2Rs86r2XGzX9uW7v9V+97Pm3OBInoP6+ssaEhebplUl/YhTXoBTuzMk5nOwzuTDnfKyM
VI4PXXlKnFo/oOuH72FBK1F613AGFIVXSQzCIjhj5TGf6k6rplYh+tC748797wrbN7MjCrg9sp1I
BZk1tX3Wve4Yvvv9Pd1/ZSdaAB/zM34cH0sn+/62DOF81kj+GQ80ekoxxpzAKTkFQQ1e1ldWQkkn
nGmg0Yusl9M2MvW40jduJNJyGou477Y005B8yDZKIUIgPvSSca44MG+J2YDtRGiwspHvrDneieK7
WuXUoYtOJCJnaBs2cnaIrn14FjLKHWz32feMnN0q15xLB6TjfqV460/OGr1NlljIDJsoamthyL2O
ePw8wLD59RfDVgfgvKVFLsOy6NfdBNq7HQUkdILxIoinhYfX2wn7CiaIpaILYfFQ419tisJ6QB0c
yfqiJ+i/t24s8wUh1yb9RwWltDK2fOugPlRDWqw98/LKcvmEafolDZTHWlc7yC933ABTzezhEh3p
VGPq2oG/9hBzyhq1Dsd5U2Q8ZieXfQUq75gSPZZNXjKbZ0uC5qdzc3PoJh/36YjS0I+Xb6ok6mBF
y/6RdiIlhuqEXVEMJG9/9xLqaWXY1qHh9Sfoj6XZvfNuseE2UWZMWbzsDp6xvLow3Qm5efM+H2wv
55kHY4rqJPC3AhuZC47cxWwJJBLK4w6UshICHYVx5+vc2btttPs82RRKsb4QvG8/f8Qv9cCYInA8
Jmztf6BQCU2G/i5AQGyBW5ioTMQRnlUvalRW6NpPUz7tn88rAGpnkg7Xd4KXkjb4mjXpvLrBaZ0F
C8dhfaCHbsiv9UEZddCMeVbEQpyRdUJZiw+xQcLdz5lolnQeNBR4kmY+U8X70zZ3dBA7ADbBELtx
nBP8Oq9EQFtf0U0I7AVsZOPYysFQrGnqesGAUdI5ngImWG22jszvA7GHExAynYWIhZPkZEWAML1P
i5M5jMXQUKyEyT7IiRjzP0Swr16PZ+2cbGWSWtvr2B2ZGAceWL2Caan5GhzhKceMBgc/cvf+dQw5
DulCEGs/g+n0gtz297uaKkzi+wx2NQzWDmM9BgwxcS/3MfeY8dPTUS1b8GGaxmszjz/mp1xwdR/P
XFtm52+BRCqETD4bF9YXh3a2CHavV2GzYsI6tFgbvzq71xUkjlIDC3cSYPKPSpZWIENKnbkmYwcp
yJeTb2l/3vJwrVarhgjmkbznl9b9ZLFIMGqrxFQM8iAwpHXlkLOWOZSCyCCxqpshkn21NiYbMLnY
mv6bUsw/tzUaVKWDiQtB3AWXqgYQe1JpJxRpfNTRwsayWEVSh3RfrMn0c9+f8BuO3fs9LH5osPzR
1VqJaSuCUNHj+MG/HURdkO5L0Rf46NE9KXmKvysUOLI63q+RKxOaJFCTDsqFXe4BCgaQ2oUNxk3a
aYD3BWAEJn2dShtApFOGEDilLEWJcw4pYtP3u/7vau8kKW/+aIznpDI7rRZsqy7jCgfcVS74wwPh
zg2S7vX2obYCKwRlyWZOT0+5eMxPAHWvzXRcSqymhGRKuMJ2ZNphy7FR/0xyyBs6tOMwLbtC3sbg
MG1WESfXcI+oAs+OJw5mhYBzHU7OetSE/ojd0MYZP+3vMOMl4pzltKq5tetTYV+JXLHTNtXTANYF
9HIgXySNnL0TIvJHmfD4ezRirHe2aZg6eQ3C6+Dr4+/HFC8Iiy2ApNCrD/wC/7DmSz8g4PWk9Ctj
pL8JjYx5hKtEdo31e3eRrFnasuNYN26u3KUa1Kuu6+xjjItCSmJbVgVFBkq7kOC4QV8ROfXSoRsy
Cfz9GfsUhbr9+/VgIiVu+RyLTu2SC7mOG3eRt1BalLYxoZEcE6AxvhcifbgTVhP/1x+C+apW7rEW
4JzNOf4FAtlgUtvmkEUNkBsCldzJBvxy0UYezaEKLM7e1SR2Zui0wtPhzQEUQ/iT9ntzbJZDo6SB
iO6je/Opu7gz7rjU/HeUlu7TapIp48LRvVdgMi4aP5NEv9GCLqx1j7T1QKpdeY+Q3Kkg24Glt16b
Z5j3uyfEZAAL+BEtyB4aofnHOG1K8H98Uy5NOkKHB7tvmC88G5Oeo+OVNdZzfT8ce048PmDv8Csf
EGKKh3CG8YA12whYAbnsomtWoFaqoH3dDpU3ChppLoDaeMjMbYOCB+cJRD+gr/oWVYazj3FWr7LY
7bXdD7/HodOaRMeWUaW8H1pZEDOVPTTmfheBToZcF3dTmfkMcM/W9VycvLhbjKx2+U2sw5eeNOGm
YTeM/SUKBJWv2d5A5ITPc7/0iWJOVKC4P7RXzMjqcRxRV2s8A/bzu2VHGircPFWjG7BI9NwH106w
MQ/dXOf4KSQAOJNTMHp44mlHNtF7Nc/1NPyOohBXndp9iuOhjv8mLf/VVBOx7CRMhYtl2QVawFbM
w9ewjs3AnNnHNiI3QhxCmh0xLPnYAC2dEIV+ImAmE+ZGbPBHJcCangAEO3vRsJWridJe9w7XZtEZ
s/lPVZ74jCfHgL6XS4xgw5W2zfm776tDMoaHsy76rM6ChxMVGL2NhYwwiU8niJWLNgVQti65OJ5l
b3XEy5mh0pYX4IhydqvBSOCJbGWMfszxF4KgfqhJ3KCEiRHGnE5r5EUihR9jRYjZercNrOHMu7Xn
TFaThyngsEG09/3zWLyunYp95TGobtu+3efBJnOSCu9xw//rPVcNa+EN35+HuJVgOa8/BbqUXxRL
vnbimNHspOfjS/8UeDlYmAAW70n849SuMOVZFfo/DMt/9pmrW5XN+WCfPDDQY+gICxueP6dg6/+q
O958mQ9ZTeQX91Pk/LOFhfzssW2PoetdRaglkNX8LcMMDkhrvp8Anr4icwGW6i3SsADJtdYwxs9Z
eIfhoEi1lsoMoiRxx9Yn2zFJWGnD/xiyfDAMXsdWnAsxIh7pU1VeyjpJAdjk69RS/xgoqvI3fYN7
/Ln1K1W8t8EhtTsonEe3vLbr8KjAIoomZDfz+q1LO0JlKEG7vjKGS1PtqTAU0V2esCXCTcDqh8sl
A1UNSVJezJN3YhfDS8sibdPd02UWH0/L5lSdXd1p5s/4cu7fk53kFlH5KZ6w2fS1Edi7OtYEnJTK
gl9iquVwlg1OHWNiTc6loCVhj9Llmnyn67mpZwVlQKevgZjGvwJko+cBl2SASOKam0JULZejCzJn
v8wtCTE4euAJuvDbILKY9FVpCQ5SWzN/Gm00VpObItFIkLi+oOw8goDw76ODMOvr3ppE/ARxKbap
NtFWhV8WgmR6ETiueGEY3+FQ4n0RKwHfTglMdG2wqbvr9mRmvoPqY+vFaJFescgMKkBqiau7K3fH
dLyLKDnvkN1eF9vv8t7EBGAN2iX/HP32eFzeprfc91g+vSv9p5P8oAaZJOHCsg/q5/D6Z7FkOEyq
R2eHAccuLmnhMUyYk3I8UmBQgxXpcSjfLTXXwXqF1wDLJ99G1rkZ509TDbORoe+y32tjo7kUoQKX
uE8fOjuftjzGgsTkQiL8HiKG7jITJquJesjr8/HpFOWYU2tZGyu0h5aHolIhLGqcxyaYo8+xb3HG
yg93tvS+805xBsbHZKbEJicaU3QDiH0zevJ5LoqzbZN+c4iBdmhJYJ4SR3zVdzV3qrayKtJe7qdf
ocY4rsYQ8HRB/rDEpWqZsQe/YU5dL3yEq0wjW0FqvptDMDp/Z2fnPLjV2cOCRdBwr4PojRVwVg9F
2e9UoxKK1Yg9zc81+gkAKK35Bo0GKaVsdJufQvbVRJ+oNvIJeIl47r9gQg4mzd2AM9rf0aCIbK/Q
J/gHcNqpsryXjLskeRBc50DsMJWgEAz4vttsuHuw3y/P65FifD0O+nSpn2RXUAIebaYsr/UV3wOw
9T5EOxruB2bFNhpm0XJF8Ag/rjzViLpAXWtlXEXSrIMIIhGjXA+EnK7BGQSlGkYDTys32HgfDd6B
wmcVKaXqjk6Me1s+sk6hCaWHaKWwZkhkpSFKpt3kNM/hCDsFWdNq86rq+PPCBLMm3bjxHa1i4gXw
Zq6gJpW9Mgl7CbbHqtGOF/mvs6ScVYXglElHxB/EY71pYI3Lus09OVX+FN/Ncf+MwD0uv2hshL56
epiocTskw1v1XNV7vuJfZltzY6/8M3Xnp4obhhFHta5vzIqPTPiogvDczGlA+vXDlaWNe96Od3B2
j6sphmBIYUD4yzNc6rYL/ZJjpgumEq8A9l0b53so2TDYeHIzdAK5BTVKVe5gcol/HCEIumyUL14U
+/5WwIHoIy/0kJ7VRCtGELTXBFnN+8o/iS2lZkMqaTbyoRO7I0gqUmWwE9Bk9z36jGu1LDzIjHsc
xyPR33pNjAtazYWbUXusMf4qUAtHQIsdApNllNeuEFJAZq0ggyWkA8HyfcfOpiSYG7ni1vNE2B6k
l45vTNMx1XNDezdwFRP+sWc9vJwCjSjc73lG8jO9wnCxpL4iwORGXuEjQquoFeF1sDxUK/twpBNZ
A2GhFFimId41uQwjfeNSCLTECBzpr4G3pcMFYBFs5rHhhenFghTlQJYCZd5j9An3QFSf7ESoshDr
ERjTVPOQTInaKTFX4RP+o2bkYs8hUNMYNmST1k8TO6GtaJsKagS8bfNt4C9mKJE+7vxSKxsahj89
jeTctyjvsQML/5ATOfR+a7ThTWnRI8T53UNFHtbHtLiuILmNceBqVQF32sDo9BT2BxEPogaYfVNq
zWvJhzpOi3KxGTq8EtPXvkrVLfa7ZkQT0fjha2SKwp+u00+HfLQOlFw51xtbr4iNhyPMKZJJ5kVQ
6FpKTMVUab4b5u19EToV+NpGX7rYr33EQc8YhctZmqbT7H8YeAeuswBspj8krbOvJYecopo6x/OX
CvAhn730TN5I4f7zxOszBTzWTcy/aIQ8QccrdHfDdlHOQk/vMXV+aIOkM7piwkiWq2BSr64eDmz8
p9Awq4HgK0KKm+Qb6/0Xmu1IFmTHZNkT21Pi9MU/p/qvN2VtgNM0JJPo6vzc8I2iBX8dhzrGOb2H
+3eD0rTKNVg4zz4=
`protect end_protected

