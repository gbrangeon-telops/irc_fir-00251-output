

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OJrNPv25gxVf6MOkMLDXm9qPvzcLiFn6cGPtPoJyX0DRSMUs1CiCHluul8VfoMGYUnRu9NzC2pDa
fD3Q+Cro6g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OO53+YxV1fz+fdQXiBafTL0TfU0s578DnGOkBDgcp0ZiS8qBHyL1R2PISafYfK37QZ2xP9F0gTav
+sG2DKzZYRShUhSDZBSgMOYpY7yZxYTXlswORtjPSorUAG9VDaJFPSJUqemfgu4AY+n/BsniNBx4
zqFaZSDmDQebEViRgn0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qtwd1yFLlmEutFKAPe2eqNz2v7W0I1lWfaUYyRoJyXavTq0FDRoJFjh1vw8Id+dlXsCh4QCKBOe5
q6ztRPULauE2vnffEDrTLD6uStkKikAcWpHaB5kHv8W/IU3+JNz65HQM8j8hOwGUzUSaTQzI6Edd
Kua78SuOo2L/RNS2CApKLh4UlLjlkL69KZuDAj8Ds+wPTUwjY2h3tf4V0N6PH8lPAy9xJk9S3EgQ
ni8vjkjW6lK8he+zqjEtOf7IEGhelGexSOLg0dP3NDhMEcaxfcI7Zo8kOCl3C+GMy2w3TEyTZkQr
3WrfN9WllC++Z6rNtRNAqHVgNVA7hObPvyuA/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y5YBoFz+YhLFw0DE8aie27jXEk9zfvZg7zgS29dcVa80RbYJrtSDIAboa1ixJiDhfiME1gY5XfYR
MSxbx3I2ZAkTI/5DwNAjKseDEksXdqu1CBQcg+U5NxNg5wWuw+vr6DqkJMxvZoI9BhjAErRu+2EZ
DgyTp7XS17TjzQ/Lk3I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
amEW+kSm8JLnUlmLoRCPt0pU7eCAirRawwzTZA3XEOaldjEiNg3FqPsvTGL5ScrzO4MhYsVv9max
1PQJ/lU1FLIUBgG3vy1UPm9QWkUIWp2rve3mDkSCfvDRku+GIP+/ziqovgiDyF46b73fS7Mrb40P
ha2QhSaORrSFucLp3v+D7rdh8lKmMq3YY+qxM1KZEpdfbausR1NP2yVxQP/t1g0w2pAjiWQM7wT5
6xmmRvYxl+7EuZQkxaCLozCO1ELg5LiuQuDVfKRWPdTIjtVbbBvnn/eTARAw8sh6+JXXfmhauCWF
cGkCTU9noi1D4Z3I/hvgJ8IXztgyejVNBMRBwQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7392)
`protect data_block
L3UZk+638iqWN0MaONJvHd+rdk+vIp5BXbEnT5LnDfYWV/yeThINI2D0D9xRAOyWAuJgdFAhwIbC
aXKgmRpzC6XYSVS7KQ/7jN+3sKt0zuaskTWH1rFhcE1Vij0bWE7T3fDYX+vewDnDOVNuACkVhFg5
Z6kjQpX0/FaofalaitsfH7kNGUhkrqA/JP/S2SF/NEA9Qgn2qLc5cIrHedWGlLqwIZZ/S8sXrxwf
ab9vytzy16NhP3FqJPImhYTRuOqCIoua1UGI7wv3xX5Zad1XvMWF7Xl6Ohcss4MLORZUg8f2ju5/
c3qZVH9KDJodANSO9bxi9gnNVffjGmgIQfLTMa14muxBXRIyprJGjATc9y360WF05RCsBeOXoQMC
CdwXW6PrAye9B5QhF3Av7rv85R73d5Y1to4DJLfc3aarU1V42QT0sSArCZcjLHy6DePuaj0Q+yht
H6mNpATOYIX0I7h83CNHMPjPdfsENCf8/Q9T1/bWpRmaP8t5R/RQmWhWi3Sl2sTUxnbETkyXKJl9
EeE5cQHWFr8QGkDFgsqXKHlaMk+7W7Y31vEOVU6wTagNdbrSQgjxAEgDLzceSBzZl98TuWg4Qe+s
a0s4tt3ObbRpOexSYjpbeOxerDelKkuYj4f2ZmY1eKXvt6O2PHaYQbcmefELUTg8vVrXgTPeQ25w
fOJ2vA6gCyIiYk9g/gSlPb9iwigQJBSjv4rbedR6MjZJIZOFAJS0Y4IWbmVNglok1HsKwA7gBTYy
9THFpVN1tI+apdaS9SNbnvL04uON5RYKUIZiudtpQe0jGwe5SO/IzQvrnSdaK2sCIKw76mtAJJRO
X7cZIJr/xCtiWuOv1Bwx/fHOvGSxSojf9fa1iwV0TpXpTHDA6EjzGOWdF+WqxLXiV2ak0GH4BzYK
tN8ThFY5lyFuRHYdeq6GzbQhB1b0Qy9FCOhktB9KUpPfVhTYaXGj3s4Tfv0A/XDEkj3f6Hhjaigb
n4j1sbm4m/7kgaNv++vC5UbPss5O5r3MNQLj5lRL0URjlz6cvvtJ0R5IPpuo63Ck0A0eFpCUN9cD
GPuFjL1ubDSIIonmS6KIp0R5r6pV0zM6XNH1QxXeqFb0GJEal933WGtxSI4oySOlCgqgq2LX9FW/
aWc40YAiD+tH9+xinyNPs0Wq6DYFxI92iTOsFPIoQfQ9LIjrclCMfJlucCJA3SibtNp48D5SWBwC
KYm3TQHiU4g4yy3ztZ3+5e77zOhQ5BJZtiQ47/ssxC7kHi35Foc5klsM2C+JVULEnHKvrXAGXDz0
I5VUAJDXnzZfTbYy7NsgQp6kv+jN7ESs6EDZmLL0RhhQ8/NZv/X9lOCB1DU8MJmgmq58e3Gdc+Ft
6H0bYxfoEThM7NuXO2yYurwUbE0izM5REyaPe/L5unbZBL0cQSAm1F/UpbBv6I0WWLzDHKuRlzkY
2ytw8HfTNMbaFuPhA251KkeFirkoHaFKIe48EXcZ/T7CCtwenXYd7DkBCfDu5CNLU/1xVgZh7pAh
MZ9pHEv81K51Z29sDcUmAFXy80S9oo/okcqSIwhgiAnSQBZTF/FSYBhJfZDtRbhShyKwqnjm7NOP
EN2rWEe3T3AEpE+5QJJycrJKIBbvKWpU+5RBGZaxOiHwYS1CVVsVI5448qIXBXWbCaCx63SvSO6G
HDZGG7fm6fL2v7ZMBSaeVbQc3AjrkUUF7ieIaxm3S1SxIjLIlC2obrsMcesm9RI9Vo0XyHeubtQb
bs0VXPtPn/hVGGGGvlp+ld32mRQvUZynB31H9azra/nMzWeVLRnYIgfdD0q2g/M3V0Wz1Jjxiwkv
c3FZe8uECTiX5hIq/xLxZ8jU/dwFSv9wGtWg25Pj2nK49QomsAQDhrDEu2EMFftlncKUCnwLs+nQ
CVPRM0mNoiuDVBjG9B7WtauotFlRJEn7AKt/mBQVVg2mru7wAI2Vro4WTi+ANv3vm8/oF+YyMyvY
OjAH1V81hQ/tUKsMMEHEZC9e0zoD3uDCWt1cGqD3QeogWlAPI/6s5me0C2jUoPEd4+rmSPPNh1tS
IyRLDg8ZuajWnxwx/G0W+cA7sGdu9wDvLcmMBah6BlVUMuAD82HP6FS20c010oHhy9Glk6psJSqA
xE+6xl/I9EcCALI4GoF1/BP28TlIcyLiZ3OfXR1+X5ehcv7VdlmxDKSrDBCd6X5l7YbN8ns13u5F
Z/7EzcDwDtJJxXhLCRM853c/4w0AqPcpUDdpXpo3+Go6ywFSSo1jyiYM+EcMu7WDH250U9t/Ouc8
dzzkLG72PaptSS6WADn3oobUaGwDxfPBiKldYCsNXCeE2oJNjPWW9NYUFW0dyomT1Jxz83Tgvq7d
5SyRfCOdiN3Wudz5B86W6DZRfZuq7vYg8ILkaXpsNsv2Z/5FOuxwvSKjeJy8PVseIRuymOdaY+m5
sl2MmbwE38v2s6VRX/12+gW5bKLzQb2CGrrH9tlkDEJzCrO/6+M8TbCvkwkKDq1ctomM5kCZJSd5
ShACSREHP5hdGrevyt0KZl4GeDXVKllieSKyCJZcK1A26YbyGBQOjVp6ZTU25UcuyO8WB6Zzo9OG
DB4DkV6XZnvfOsp2Umi++u932HIJbaSMFSLHNVoVpMPEtjfv9Z7NxOeoOpolyeliV0R2Bl/5ZcAB
RusxFqHgzVaG1BzSVNl6OWZhDo19MIzEkN+wS0FXA87r7Xp920l/+ieQcXHDuQRrMPAhAk0dMl10
CC4HFw3IE2GxzjkZ+TOXycir7ZVHmLLLGVRckTsMnGqUOP8sbzEbc4giEkP3PxqBPCEWEYiy5/8B
9bMbhGP8wsOjJvojbZgG44XJtb1iI33kfRBv4WDcZuW0XmgWrMjpjWMi2GFrEj78AEtoe+r6Lhd9
oCRvI32PnR2O46leQJ7N3wNJWh38TdKDWVCUUdhER9D/YsV2zRJz2zvDJ2Dr5S8SILxQM6hp0aaW
FJmZKRCMsW8yv/oY0NOhaaLpJPmvBg80xDFJNjMlwL0vESEKaY4MvcT+Xum2iRKQFl5I4wPvwowG
D9vpQW+4+VrkogbmZnq82S+wOwaMr1Uz70T+zaCZ6rUMX+3QVQxNseSN/bS9Fy5U9js1sz4eu64A
S4Ghm7RojcXjtp8Thu4ywT15coqAiqMRfpDN7QEfTDZgpMnKF9+G0svPgAUv2Dojtt1nT0Mymp2l
/7WZb4uDv0fnUqtBdROWGVtSfZxl0XfdkDpc0+K4L60yYpaAcORQuJRdP/8LYxTzK3zBz5OZBwAm
XHp9P+djlpEAEo3q4heoRQOHD+9jtQ6W9ykvR2A+L8ojWJ/rVEnJsT7Li1zAEDLAa11O5DeTvp3i
/IWrH+7kcxXHVFcS6sgtpNWz8vlrxaLIaWunwv9XnY/fphflZZal+CksrcrJdnG85PELaP4C2V35
y48mxl7tyd+IwI2/N9tOr6P+TQl1ri6HTvE85yFF6vHRBBdj2kWKecPRP1VLUybnsnlmAJ78JGkQ
2mnyZmKI+hIHk09TiZi6d/mwREwEesTlK1S1MS9jG8PakhPU8wt0iIAlXLZJRw0PARli7Eg6TGrJ
NwlyYrWIjMGu90UF84gWrgNTEqyT8+9jnpz2BdmiIvVd5QhYHwhCqSzLzTjwGFx1yOv03KSRw6dN
xePWYmeV4s+rPZNIJGzIs+b4cFKzrsTZVt9TLXiCMF0xcHZW5al0zwBHZFX7zPR3RqtNW2rGJn5A
6bxIfs6g6mVEgZAnNmbo5e0hm3ujqGrTX0Vz6NoUnPZkd16D9m7xiplB3oSDlNwzq+0XSHtBM5f2
8lvGPcUCW5e4UXwv7etlNWpndtinBJmsmCbByjYq9iz3Cr7E0rWvToMHm2pKsm6qinvz/HQDVWWJ
v1MqPhOVSbNhrKQBzZXeW8X2sFnlkHdd6hRmdltK33fbkImCmVJKGJLBRMUFbiKeRIodeR5nTClm
Dsz+dsMdbvylF8rwjV7mmiV04u26mbVcEMtLzHST2RWfFaxp87yTP+0hgD/pM3Po06lWbLpmTc2c
DJeqSqgZF5eliYt2U5mNNOljdfQTT9W5SbEohcxeEUymLmmKc8cwrSygJUZ8CElm3mCUZ1XZG+cI
udMRcAnWWAkQgJ9G1evPXNl5T7ybkADC+K/Z1LPsl+6BpBpoOMYW3DW1Ic3T6tmYXhXQznkHtbov
zREiQw4jv4fleb/QttAmZUm6/Qa7+pk6kyyJz/hOOnGWYKcswIRJmV50QJjDUQ6IUzoKara2Iwe1
nhigyv+QmniS/TZkkKZkyNasnwXmESDJ0oA8PgAOgQC5QMluRWqLkJAcr/M9bGhxcYqdYtdvqbJr
iLbnn5AN1MTVZVgenkm6r86CCii2246MtDX2cjQo3Gvr6hVxz2UJLftkaO8ONDYMqoiMKbdTmjsk
CHOGTlCIzSGtK2iLXMoLmp2TBcuD/IuHRvZRzIwzyx448MWanS3b3POv+EX4P1mrVb5cmku87AW4
VqcD57lteDcGsjFKkMMcNZUVK//6hCrrZjVxmZjRfPb12xr8TfGiy00SmNwZZ/mzIwIsKvAl44ye
9dMhyOZ1IUcXKY0oBoAvHYQ10iE9VC6MIrhLvvyRC0Fqkgx2MJEzlmQAdHV4siqXHwDPD4Vf64wM
StvF+NrgDD0GNFfiGMSnT00BvNiHqpfwcTN03E9thdY8cvGC68Ut/1mi611LQj9qHpnVPnqT7/VF
q9uP2awD0g2+IaDNPhvycxEP0eq6oRjMqnuRCN98mxA6BZMFJKiKM6ph9LhSpo9KOZqOR+p6w0+q
8LwnQbjkB5ED33E8Kt0fBts8rnS8RhQAwa2t56XKnvQ3hOTlPDJLtFAV9kqfu1tL9EHUD0NprznO
LK1N/O70eH2o/Ik1rH0X2vAWwJ2DIgJgqRsGit1rzMWHXxuCws+RwWD1MB/fDNQNe4dqH0tLhIZ7
eV3uThFhOubHGf/S0ndMeijGME93tQRfdZ/2Wk2ilFXGR5Y8G6jZ6D6HdxG8FXURoLNY70g2TY8g
fu4NmOh7h/GFXMstelbf9ja7S2bQBcN79CE0BisxuLMqLUSlZuoXiLt87op4MXmdLY62n99w5p+J
1hAqmQF3VdHVGDiPyQz0xj93sbV0Pu0Rffh4dmQmmY2S8415sRpgYLYNHYsOgwgZABSW1coWRVMM
DaATxZvrPTy2lF0GXpDsX3ee94OTeJNUTnj7+2U9Gq2yr0RwZFMxDcLuK3rbHCZJ+WTvZea6sBje
WUfYKfdE1xG9iGrn3t+A+S05jLhyLWU/uI8doU0z3aXIXnD7BtrTcnnUP5DEKTbxVLgQGdTZviOo
xxpjqeiutOrrAJHh8nOlK5hrO2s295ETIbGrti2qq8dU/j0d9e8r0l3jeyO6dp0WLVhXxVQoNRif
R0sgxggPBHhRotoHz83wWof/5mWyG58f6x+mtDz5+miz5UlyrGlYmc/Ti7Sk16yiW2xzSdTNed9+
8tF74zRZj+NaQq73Qk+cPx3Yqwk6jCPH/rzQF29G5NCOGFwt2Ixju9S+LvcflRXr1Eis52VyGpTR
aPFGZAWAVljtjeWpwyFdyGt08WIExgv6BPRlBY65csn4+ffD+6UAAZAHGjRDH/W9S80VKpHd1lL9
v4dqcEddqvbBmuwVjWaBGr+KqSNeAdzP52EjoDFKpTkAfXoCLHI2baUldiyFJUGeIaKmKCQynV1B
Xzdi5ZKnEXarsgNp/9wI0ho9FpzmIiIatVPaTreCcU8NZLScPtAwNN01yvJP2gJ1t7xyiRESwikA
3hjzX6z5iJQDg6yPIZVxLpt7a3V800eKPnZX8gqtMbnsAX8UdzO6loqSPsCnnGFsAWOQvis/FKYx
smhrdySjc6NqRI1QTMHdRNsrpsHWCT7g+ANiSL/Ca/gpmT624RJjGaIzupg76MwFuMQNi0dg3axx
T01LJkLR7kqREcbf81YEvpFpLQsgoCTfcY1ltSUwNBZ3w8PY1mOvzxPNQ9Y5KUO/vvhuJuRk+/SW
oWIhoMiPC6Cbizih7DPYsz9rAZLQc/P2AGlotjfxBzYYOeoHtktdsuL+PipvgKF8G+2NvrHfg4dj
hHKdOImm39c11GRLUW9ztWV8QWJkkdPR/W8UxFnnKDUxbivOQKReEiX8UqXfTAbjKhTGrMSft8qE
HB+hfkusYBg/f6YRoFYIQcQSoPLdj6t+mWKGlc8lPW3QaK8vaXWAQoo5IHoeTv0LFq/jiDi19DKQ
ajhEqj6mjPw5BY00ZImIZyT3PbEKeSV3GlXJuMvDpfJzEseFWwigsEke5R1aaL7agS4laI/nyAv2
clG7On6dCk7eYIMC6dF6AK/FtjZMSQDv3v5Q4FVgB5Kx/fRgtSgTjLth5uwjdkN5DpvGBpsU0KVj
lMUjMkKJSMIZUOffNoR9Cdm2uvAr3WdayX7q+wF6lB30/n41ctykq6+nduGQC1ZTeStuWkbw+oX4
/8zpE22fCMLXWoJraA8yzQBJCoPts7feCqcA85EEiddTPaZBWuGjEwRkA0aYT/FUu3ieMMK106lp
atuw1i+rpv+6tpVoDAfxxWsXtVPDWIN3NO7Y5lptS8Ru2unR8szIQPiypQJj5guwDw8N8IxhB6h8
+J1cgkNya+rlkTxuej9sjeRDrwTUC3w9W/qeNLq9NFn1yMKWJ7l6CR752DRPGOQZDBXnGXTC5bpq
p30jJ81MEhacFDEL4Ad5b3AkfwToTwyG4YEgyRiNC6AD0Cx2ct9msWR3PAnrCOP8HQy6Y5NU73oD
We7N/YTb0vMxSVGjjKDa7j/c9OFngAjDe8cFQjbPky0e/LGsoMVjG3w6ZiomITN+CaHTr9gphL9G
j2ehsmagg158diH/vDONsMNq5cD7SY4p8zRjsojohDHIv1SXe0UVZGOJNNnMPgno19JHkQneY4lK
WSgAtyWOaejryX7v2xPecncuwEol4Zo7tnN/NWdw5+S5QK96QOMxpDlh7spT7xDXul6+G0t3eDJe
HjzibYe2qxKMbIMeJJdg1d/EMKD+KmADe07/uWB+UB08rcopnuwpnvbsiZ/v/kPT8U4+3a0VS9uS
JvwcT573a0sJR7WElYtDJtSdZ5jw6z69xPxGQKZHWHsrj3Fo7pZw5vPIVHzuSZfd+fvFhsDrlwnh
SVUnHSqXzxFlD93sF41uWbZSKNcQSEbAVCPJNiKz+RWAz6SdHGROG0bVwItpIjvUtH1U/Q/kg4pq
pp/dqbA1XnBQRuZsCMozbl5KAc08e2Ua9U91KcVxv9tbFxUW8njSo/sTI+jOk/OkLyBrUFMbT/05
ZwlohVtbFsqeCTFBiICbHRvNNHBjIhASlMp56Gy4nbgtI6lJNSIU8e1p0tnzednIlJQxhal+bUWF
7jDAn8lBrgjAWeHYcuytP1Xa5qD6tALJj/YJ3sd+wAZqG7N5TYnHQoyAA2W4nD+7DE/T7mmsVO2e
gum+9IzbmTS7SgL5QC/dW+GbL3AL3UBOJYgfr3YWWVD0/pL73CBf+XUsaHkN/RVGaxI+8BVA+dcX
C43H1zxBheIjEeScye98jfQ1VnzMLC70TcbKga/p0c0gzouzf2osMq0n3rR/PmnqRkRPS1iA/GR3
o9gqQRaLsAidlmGJayKyuI/edovRYBT45rHq4uVCYv4qDXR7+//1QENsMpbhTb82RK0j6X7LPlwP
/73bED0JJUyoFQDK76y1NRd49Cdlquakj6eOIOFCLdpbFAXTpLpcqogZvGbJqZ1vAL/Ajkg6O4dE
Uruc8b8RzIIiZ9sgyOWqJOdH8CCf2DMEtZqgh42U7E8BzLhuIuDCLlYq6AUVUJaL+jN/qt7ox+G3
B3EbxZfsFBQJ/VqsFa+dDZWJpZ9Jbszsl12aSrbuUcIvBMXTCJDvd3DhYyg7wCIBcjc6Op62vbbV
OZPqZJ5p+h3Bdv9VYtFG5Ev2n/63+eTTd0UAfmBgs6Kn6fi+mdky8wvKvdggW3/Gn8bv9QAono+T
ULMvkoCJmFy9oF0x7tZ92BJDcWzb5KaI7ngdOMXe7fCChM8WJdyF8H3RAc7/CgC7+xx1+C/C2VAV
/iBZUEDmrx16HMltWx+vqj0mujqTf1JRC0Sw5HE8Ogg+V3TQhP1bWwMQSaUx2s1B8JPD+u+lp5zW
i0iNmdMC0xhc7MzZkc2tfL/N6vNM9xo4GjlL0Irb2xXOi2s7gQTAu00QQrBLU3CoaKc/UTDiXcN/
CHpwa6jJanco6nF2emZgwGpJdd8P/m1RwEaY2MdJSr9/otPy16eqwqLHU4R5hjHkUBXAuvGNW2mf
L2IuuVF5Iow/j2TgjZ6c6aQhk84vbkadSBVvJ+WZ/n70pZi1LBOFSiKp3L2z3DjGt6R4G3/PyzVF
V+pa1qiRb4YaB8I14XTovSZPae6Pcz8IGGkepYDbijaRM1NKoqVSM0AUl3oAft3dpBQCfLJHHU+g
f5vpN0326jWFiN8vvacVqMa2RWOhfLHMYeXesQRAlFbQo9yBc2Z9RL3y/bXgWxLRfmzD9WgsGtXy
EoRg665mLJ33cM5hzeSTK8Z72f0ZOPXYyHDk0ly5UJaipCMsCIvMKJKu+WQO+4HrPkXteWFOYUkC
a0xTJdfpXRSjjyamAz4cC4h5elgxqD3WrY2dQ5kpJlDv4D6xqLlcMkKDxZX6RfWv4MmrQVrTwTlt
dBGGxPDrCZdC+DP4WGDbnSmOC/QdiUZPKBLZxUFbaouAXzeKhP5PKKGnwuQhmbDW3QAdvyJCTNhy
Z0RZs2Gj8scXfSJll3fB2OGvEdZ6SiIYcjMoTcB9+kXlp083Dh0ux73dKkK2Djo4FxQ2b6DUm/w5
xqEKXcgt3QaxLIRvW6OvVnqUuAeBg9SDm9vqa24LweqswDYvV17dGDPCUeT/cYSIDVGRS+rlCTBr
fhwNf1MzI1j7WrB5s0ypU+jYnsvoSCYadcCLj79ZipoocLSlvBcNUtUuCXZTUu+VEih2ZBDJPoIc
dvY22gKrYisTYzsUGwbQxFwU0VbK/qbuL+kj7qrWLSw6Zi50pyTv5ckPHheY5EXyJcP7RAOPZl//
kk0/o8RvI4kVo590ONgO99l0VbzDWN4Tbg/39Td+fUagFyGih426Z2ka8sJ3UrNbp576VJymrx16
tOuPI26NgVxQJOPi1xGWj0/SqgP+/P+Uatz4Szebt1OVdtir6YH4Nn/3kXVj4JLfKFzVQS76z67S
RwiMi9kzi5JmbxoWOuKFH4LNHut2u3EtgCsrDhVcNypvRrMHikEom8c54cWbBe0OiwBO4edxM+SB
ntaD78rTTpAW5XB76OdpBhfku0dJqs2BB5paJcd5NY+xA8mJXqLpTI+9GezoqsNkMu3X94GJrl9C
ZT1OuJP9fXWPdnM4b155MV7xNfs4PF5eNVZRvqww2FcxqW3JQo+dJw3q5r7iRPzdg1Ks5yJqNv+B
nvnoaTJ4WXG8dxyTIW/cQJPVPgUPKHd+9cS60pz3RYSmPuj4AVv71Hb3vwov72cC6whLZhubW+z3
Apz+xw7ushnf2xVSTcwLz4Is3J6CO8NBc5pZBZf5tZgz4h1vad9qLEBVU7zK+VuIoMn594hYf3qc
5fHEDcN/OqYlRnxecngJ5VVepGYFZuzuAdL3eThKl8C/pqu9DP66ycJVkySiB2Z5jGonuyfXZn6Q
ZDjQnYMDBQZ4LOjaFwfu3Cpm6sHWq8hk4pSVe+zIapCAtXfZFzZsWELFi5CbFCX2P8gKWOPBaSUt
SepttHxLOBfNCSQKyxIGWnOwXRXgGjxK8/9f2nhsv4XmbZnhY7rj2cWyLJma5t0jMt/tZKWTuVzp
clwHGln99vr2RYUW7pikuVzHOsZYl/c90RZgR/lwvkrFz1gw2Gue
`protect end_protected

