

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GuWEw077quLd3kfu8DABFf0P+6oHLq5R3U5znEygNXmkCks1DFRW7Mt6/jd95Z4sdDaR5vCLL2M6
FB/Ff+rNvA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jFvcfNCzhBWpeT533DDm5MsDXv4GiB5r4Bmmnk5Von/5jho0+BIo5IwIRMf+AlV4xqtSYYHC3I2k
BVrljYddp4kTGUJvHCrm4WaY6cktxQlEnZCt6LbtmRJq5bQ0+BhbjRb+yhnUtxVO+mqZJ8X5carS
6TiI+a3eiQyqjafsIxQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3uk2ioXVXgv772p2rHBKB55nN0zepBz6/NR5erkVu2PDHMiL0sh4KhStRZxPeDNzjzcvfXxTocKd
hKd8wwyqbvI0xJMti7Zm3ArPWxG9sxsPGJWi/HV3nwjRdbl8Q5i42ko8FFW76K8gPbQTkcXqEX+f
TMDFgnzTvHtLMrE1Xm+zXTsDfz2iY7i6oQ9oV094lrdSLAt80D9E8ysTFrLsOAY7rvOt1c8o26ui
lfC5xFONM+l+w+GytYmCYLC1g3/Ymlqj+CUT7JBGrc9OLEVB2jBY9OOPdBfOl49VdH6n2k4l06g4
tPQ+CDbASlaP1IKOpWeipcMMiP2EcvQEvzBqvw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ODN1qSeI0EeO28pILhOMZHx9bb2qYpmwvyQXvKPrPhpTBylybxluT1/v8KSBCRH/tKp0Ke1TAM0D
rxIBcEp/+xGCTqhzkt5p1fRCsGDy/1Kk5L4fYaTlJRk43uSfOTxn6cMlcuTzjFQ5x+FkobtNDSvc
hzmRwInNRUY241xhR0o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dC/Y1fV+mqTG5rOr6IWyGTQ8KnFRPeLZShUWaAXrkw+Ng+xoimVrmPwEeCnURpwc/T0yNbEjCDB4
bGeW47AlClSVksRroIGKMbG4EdH+85GyM7JEd8UxBfmIEn2qUdv8H40fYW6ndPlPBbIsiprcQqu1
BO1TrP+zbizezYEZNLdme7klmciNF64y46dVM3KfXIDNKQvoLTlpJYClTv0K9dc9pDZOVD/5ly4k
Nh9OSLv/jIhCDn0y3M3rX1DyQgZeJYBkDd4IBP3NH/wojvEFQZAcMKJEqADK3qsWu81U6IIzKfXC
PUyRFWat+MUxb64pAuTyWw3derZjtBnOfD89TQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54432)
`protect data_block
er6bfLA53k5mu0aC6q0HGT5o6hAJ+2tpOw2gR3ktInJoXQvDE5EquYMHXo4hCDQapLxss0ziMkTt
vpGfc6nkf3RCGXdjvo8/mWsVRFQE+UAr8TgexU8i23px1s7K63EcRwRlRpimFFofhRF9vqROTUYh
ZkCgCCY15AlzIQD+SVPaUcIG/Gcc8fSS3Yj5D+K6bvyHe6tzCtiWfnDXLdEV0nwcOirBpOtEFm6f
HX03EMI30z9rUYF3DR0xgDgRtltUO9F78koy0gc8BRqeFtsPzMZDb2DtWFhmgh5YQwKUThKYTVaQ
FwgrHIQQwrZb8TTTbLDJBLnJ3WK2sOyTPGPqrJXZSdKJLGfnSGCXEKnUZN/kfT0+fSlbf79o5IGT
3+tIYooQF8GtuyHbVHpvn/XgLBNpYY0Q9VYGC87uWPpw2gwVtWADCTlIFleJ5+aC/qlwLPNIgde4
2S1DehXpbXZ7yZVM/JKRnIwyc2vxpdm96287B05Qjsc9d41QFnWmkqORttZpzBOuE0WEmkYsZu+R
PhKNuPFw14nKNFDbcLQOHjm+qb39S+LU1T+HUalvmG/yHjPmar101uyCJbq//mXAtKsBKLlX2GWL
9K53sEa8LKXaJRnYiA7BAECPi0ZNwX6MvglddIkRjvb5iMJkirw+3GM3RRHfaPvPZ9DZxhtyJynT
RZwVKf/hyc0p5yAzH67BZUbUER6jf/TKd0kp84eOFPDXOyQInjQG1oE/eKnuto/94TJqb6q1nAc4
gh5h1GcWcAcyVWkZXxq4wRG9e+R2o1HjlYZz3hAPw19VXBUzB1tWhc0rY/J9Rj8DAl6GLjK/utqr
NlR5brDykl6MCKQ6N6qC+qtP0bKz49TG6u9ZKGHS5UHfoZKsdZQ2axUFhJWkDICrvn+Cr+FP0JXZ
/TfOnZ8a/ICn2hLxTfFX93CA0YnVlA64QWsOfFvsScFVG8wpqmt02hQeqBBvlwrnIWgBeLJ2jSy2
3kX8WQ69P2ZiZ6KJyreWfHhU5fVtn9DZRmbXNlY9D3Lpyl9Sy6HGuYsS7DQJXShgmjY381Zq0pa8
btosAA+zb2Fhjuxz1zzntm7g2Qp2oQX1J3LJoGLeGsijHJ41PumCnOsx2nYZ+kc4Vyi8fQH4OgNW
xlHGfo2ARhok39NvlXGNdf/7cmjLzV3qVgyk2LYafpdV+HcfLpGsdqxgiXGFinWlv3nik5SU+Gkw
oH/u1C9/iijVWSBgiU0Rzl9n1NvlCD5io553FRkedJ8MhK9Zj9n2vGK+bn0FOeJ1WSwrineWRt+M
r/704Mk9y9JkEGeYk2wDv6iqSBNxJ6WDDBWjNFxDo4YHKGJRSrdGNTXWa2GUXEd/ecCPgFNndvr7
+8GJrVlAvNKzgN9rJMEyNW+YQrOr03DyscoQ4F7kCgwFmQiFvt8XgpIQMIK7yJjXDCDGbaHBzh5x
Y4Xu1R+eQUoAK/cr2cnvfXyDfWkZ1zX4DceJk++a4fYdsN5PgwnsYxrJvk7bvsMVflPSyU8j0Yr1
6bYdFQB4n0Y2iE5je8IuKtwNbm2VBw9jSY5czJFyCJ8uWTx/dQlqc9tLXXVUZwoP9tnNTCFBWSOB
AJU2iigKdmUcf8/g3mO46+UYCOufhXcJ2yuUVUh/xUSDjEUKHmMtxoDNkPNNygxcUJduhTUivZ1v
DYEEI1xlTKTZ9nOBqvokAEI/BjLff6IUo3uRqwxATTEP1nIS/tKo29sJhf7hMOuAtMYRo4k4gmas
VEecmQOctS0hOoezPpLlu1smLsI2/pNq7s1aEcBmpYNAG2lNNd0GWPW/FUwofGPuJjEty2w9abz4
zD9iyFL5KzvAlF7UUyzBsuyrClF4B85q+bZkpCbCGOany5oXq/+T65l+BQofkTQ8XQKGm/XsqERp
HTleqAulSSXpHN3KbcXoQRVxZbDRQjQYgRD/QR6RQuCWqQU6rWr60fq6NjyyqL2xxb1xrXlz4Q5o
PnHhjxNSvVV6vKfnQbZ7VCIuarSblX7QcVIrvSIghZXyBJl8bjiOJIYIdI72E4hP6iNU+momL0Z9
SZ6+w9OTG1gQwpyPwZZrUoXyOgojifSnGfzaLnGSRT0YRyhUxP0BWAyRpz9CjcmV11T76DXmWx4A
0qKyYfw2aPQvc7OVOJIfVuxGglqmumwOhNsHb3QEablw+L0tanmTgusOUyCCcFzgwNFdPsvT/+MO
8JiJ/2UOU9xFHI9ljjrMS0AgoBPQuDFUyrvreCqD4kcorp8fdg+o0rf84wlx1JtofJS6Acq/vgJW
9d5Fe8t7SrWGZDxdZl4JpRZ0nl6ZzX6z13fe1OMdBKO1HtPpQIVXCtvQfWrwwj0yXHdvmHICORTK
S2brBUULwq8hvV4+3c0ogQP7b9lREkkN3+ruTG5pBhv42jTqnnFpLOO5get9I8J2gpx1e2o+7XbF
PNEmtZrGzALOsP8GrmkASCSryV4Dl8GUj4Y2dhcz+nz1zw+lE5d6smoCe/6Jo8TPDe8XeWo4IR+i
PaHp7alAdkAiH4lnTgchhlD22xRi86FGoAxLLvQuXHOsz1+2FljsTA4KnB5VkdU5yh/3FWHiTs0X
KZ48mJrAF+PRrYR8CcASUqokRnGvcAb5Fmqd8A5xOGMJ1moO7ViNAvyXCxRjEKo+mFwjAIzP0uUH
rRqj6vph2eD98XlN/eP45QcFcup/c0jX4E4WbVSrmKyf033P6mnqmmC5c0tF0Dc9Zb+AW+CAM0gj
5caeXGL50w/4A+cUgMZ4+Y0umiK2sXJaCjLwv6QbViRFGPMn3YFSC5esL6H2jnq2H8b0bD390nq9
wdxZLcUYhdlSMbyKFzv27xGhJoJm6vgvK9exGZaJ5wMj0qi146sOgf7OazbUTIf2mRBN8x47TMNO
DWb3gTa4RRvLTDhaVdJLRhZKL4RbY2S0MyHs/9FYodOwm2x8cZyIBdAC2nbNG6QMmPg/uvgC73YR
0mBgBKQ73yW1ja++8oUn0UPhcwlq2qRYbS12nxC1Foje+uU7JlEEF+RfewNXpxkXLt/yOPEIAEim
rq79qWQRu+7upJgskEegaN10jlT4pFWKyCkOyZaC+9S/lKyI/wvK2ugSkeUtML/3W8kLoaAtSFza
ZvTh1bXuU59RSsnWOI/jXJcckqkE4+ILyWiYFMYgC8dWuNnZu7dQOhT9DhNUMrUeruHA7Ru8JV8j
bYzwf+7G3692BNTSC4kLbBF3x9g3GEZizx58XmDbr9yPPGUsZV3xV2TziSm8vrvVsLubZUMLDElc
2tBDO5AgxgG8Jb6tpOzQME13MwlCINhIRZsacCsEwAuCkmLkdhQH6lmSVvFUifBDiVAIsm+mWXXn
Gig1phIA6kZF7jBJ4KwFnMrSRDmCjOx/0YQyZ3mgZ3Vw6SrZK6zaKBkuFD2VF3zjs57VsilMsaVt
MikH5M2hdZFB/ESGRLQcctQgLaRY0HCGlL5UmYVGoUy7SoNczA1QO+rk1GPLeAZ9sgTL25B2RFjD
ppX3jOBXRZ2wwn1My3fXrFiFzsoRX8Z+PaOEbDOjiGhe5wGWHHCKhie7Oz4X29ciDwU1Q8dzkAXy
KyS83dlndFjI2U11U4ed3Ae4BUQtePDJpTp7PcToM7Bqo2At2nnOepVBVKjaBjSS9o1c8di88nO2
MvFc+tZCYjkZ+syv4wKicU/QDdQRzua0g8VjbW7q5SeivN6gI9qcBPAwpHe26cUhH8IL4iiMVcjq
NbqrjhkZ4Ex8OIq4KiVvnLPfS26MPlTkeQoZa+gAskigiLBnCi6t+4NIoOQ4W1gbbjjGxM1w2V+2
lZ+UDX18i9HO61vEtASO5B0eV/DwNbMP2yCcJCIag8eLV8MzgbKobkJoBtvsFeaIQzUAUnKQ2DzC
LErKb+mWfMPAdoTJlOeTzyTEIAEqviy1E+lYztt0UKMUiIPbNgjAFuwFVD7aFL6QgBCLsdHOAHlB
7OBZ5uUolnzWbUIj3qtAW3sjMfuM5dId6bN/FdGmbzvcH4WljZSUy2xoMFEKEo/W0W7j0o9T89W5
7M7rqV66DWmkkSl5T98eRJLba6EkmaAK4k8E0K7SIikScrEI7h9qymySjw/LOR9Dp0SSnp0w+vQl
hSiY24+T0u9DYXjIg/UFMQsHulDmkQi6279s3sk9jEBLia3oEUInCV89vNR28jceDLgQUJYyTGJp
rIdOCD8w25YDHzMIcr889RLKlXALMwGF2L/pJX4cguFA5EDaBCCFAMUCydufYthQZj81ANLYyWmi
sMa6BzclutU+i+yt9LPyhoStzMVPvEHOhS4WNtzBqoNnhXcohXGs1B72f/XhS6LiiBSzk1aZYUKA
hMfL9q4+NTVloKCzWGWWcl1sUuO8l1kzdMANXw6+Ugf9bcRyp55khpACxXj3Fi417B8mdoIKKo5E
L/49llYfHdNQQUtWiKwtX24ltZR+uO1b0vhnYvkv88qYd6npl6O5/bB45zWHWH2rku0qbgkZTdga
drzLCQ3eN5JI/BFCg6aQrmkOYsHZGu34i/cq7eAp+dxgqArq8nXSfMIWPQL01PHfpyN74Avs/pG6
bBUjBZlFGXqga58nAsgX5euTQhqb82uhJ23IgwXrPkBuHXIoP0cRT1Pl89YP8DshsfmtpW8dmLZB
MZWXuEd4sxsy/ZPt7ZfjpJQ6VnTsCP+kCol8LlAsLFCHPMkI1yvxbf0MvigxroDXmFUNb2QCmZI1
8ziBsqtYYE+oJ9p1L3JrLijTRs7H77BuhbVBxf8qouWWaUaTfPvNeJ/GmpM62KoErFRWkVM0A4xp
Nrb1CjGVlIWZgZFdUwZ5FiOI84qyEqzsfpPtKIi7izPZZ+MMpR+0albm74TPRNS/TKqS+AsyCI0u
VlOhX6ZRrSF5LHhMfVYTMTveT/iOOr+vkokhKoKl4oalbik+R8ebhHk1tWj0NTBa7W/e3JSNzNfY
O71ap8eu1KqhHnxJk57luBgLLhrHfzh79zS+6BWXXag+Ho0SIFPcE/OevvOxGt4QBu/lmqV0yRrK
5aGJx656wPkmkW/OMzm0PtbNTNzxBJhQf4dafgInRsAbSkc619UbQTNwjgClN/h9+5CxqJiEWzF3
EGs6eqqOyyTPA8XdaMMd1bPlubySBzIxBFz4C/ogjkboSJnpLhXBoV/mCLdStRcK6kiBbU0dqiBp
bO1o70Upbgz20NuoD/7uAlDVBaxQDiK1dMaT6GtIAMtkisOxP58HXdufu76mZZP0ck1SPTxMv/oS
AIifMty6pcIvv4+HVyk3dVowvtsoiY9sCqwjEHibc8y7L9kNPfT7qnHEi2jnSmj8B1CcfB/VHlVQ
O/MM4xK7/cWMLfgHdfdODjIng0qE2R5N25XeWYsHbxwTI1H7ugfeOlk0HzZHvKQE1Xx6Hecfe1RY
6ub1ZZR8vO6E/gzFcEF4fXrrPociMEGzx5pcFOF/2xb2dM5HgoxwckZ3w0vKPzuq4JkJ8Al17M1d
Ds3cjYYBMpZN8xqf3xluwZPXz5hrAvtBdpbVbWXiaSTwB/U88ZQHuA/FYcv59rPFZIpBLXYs/f+P
i5f8FSKDfTVDK35JefBgfeflNFi958qJvMbw+6u1F2SKMhXE9BBrnSpcGCET/veUuwudMEBkKLwB
6lMDlf/nGDqgQiAozpWJzHS4ztl9iMPWauCv2H+vQi8ltgTDoc/M0VKi8ywAC/UFa1U7r0xj7RNy
zSUlTn27TK4E/ShTOCreTFGv2cK9M5S2pG+bd88dC76tnsR2v462NqaHU6ksCG54UoWfdDkCLRny
/ApLEd27j500NUbUgUAT08h/NAttprCcBmLmxL32ruouhDE0nUw1lClwgigEWUN2G0UoC3VB1gUt
zdXts1cNa6xuh6zJQXlwxrJVKlXF+SUllpEvQ1UO8wVjMhMT3jPokfNWyHxH8GxrHjyOZwHCNqQ8
4SvIDV15CqoCEQ+8JczquJy7Xuebuy7GtCTRo1cLY7RXMwmclMwy8RhxV2jSCI+6dELAsjpsJ5fN
eY9dFKpT7odCWBLJzwzRuSyelZVhzKOuKUar9aMW1bdyzDWuCmaznAQqBEIGD41H/yAAJCOY4wMu
/MESYpFRthPGh1r7W/lFJWG4CaJXdSZzfvt8TMQAKBO8Gppcc3ZEzQ9JsmZLKwrSwZB2e1Dlea/q
6YM2wdCUl0fFt+/YBpHJKFKNiZU7UFOChWxyC6W/JtrW00kT7yHHN2zgKCcLM+OmsDZyIYt0OAHB
vhhfjcD6c1o/2/syJCfqD6jQ2dm1MNuDw9gjP2SpyCxog5b7rma0S6lp0L/ZsoXlNlXwsi5RxazB
m/CDIsdrXoSvobBZy3G7VCcQqNdnWFdqemkmjS8GqCdL7XohgfIsY3BlIzaEPleUqy3OyNldHdSa
duZyog2dqA9HjfURy2UEYDFocF/2l8UO3zvmKjG4haeC847WdGsIA7QAsjVd9fw6lWgfNItmjNjg
PbSfZPDR7WWnlzRM1efkN9zf5iCwsN5gYyRhmx9m+It/kVLBkz9OMq+M8vehYcngioIF6HzygjXb
34yVUFW7I8JMpjd/gg3W8tP7VPv6b0w8BshYEpOWq4RGmq3QXg87y1Iuleo/ZUcU4+t+dJAq7ykT
E7Lkv2SubYm3cCBZzWL0nxkHS7SJrn3Wp7lvqHPnTa2W7GaauW6BoXy3Xo+JFgSW/NHBcV4rvgI5
/bPhH9aP1mW537POA0U1zgaqJQX5FWiVaL4e+euau8tX5jnliN0aJWoXKd1X31v3k/gkzgy4WiYV
W4fVg76QGWz/MSHQ7x1lALAmK86n7Jf3A6v2uGzvyNw/IRlndqal5ZiU3egWU9vmCWr+IU5I8QS8
CJp64owCaiRJZkkPgiDVMG6PAKQFTD/tm+owaU+CEpDMQ9RLggHpj9kQmeNnfYIULH0Y031po2LZ
3jE74g6rndQDR10SDjoW0b4jw1Jlop+M53FyRA6j4H3c9unPNZXHAPIOtTIYbNufm6Z2tC5lQ4is
I9m7rALLS+GOSBG7e1QXzYH+OtRw/FZ2oqLFyveyv2v2F42C9+D/6CxgAYVXen/Im7zq9i1a4Qsh
r1P56mEz43uf/HVC8RpvUvk9E79AaRJulnSHaQhJBeeYAjWQ6jX1anFVp0RjAUTKQl7QVw543YjM
JhNnln3XgVDqxgal09H9gS3xuOpQFMiUO2xs6k4kJrTj6aGz8+nQ3SZ7DnPjcVLrJ+c1/hmjEdE/
W/Bgb6eiahEchF17KcNaD+cj/UIJh6egmOIYmHCy7T4A5bCoLkbuBc8/eKOUi0vNfkFpbA20CUSh
KrCcw6JowduwWTCzglrVr9Gd1Tb2hp77SA/fuKLO0i1DQzRjIHQEzSiv3tdMXkOvqxCrBd0nzT27
5tgvVwsHm2haHM1esAV9i3N2K6XYwSLb1s7Jd4H5NrEeWvHOMnoFCyJsVetIP6ubqtPnHfDHVZcJ
gLjGbuxm5OF92dXsg+vEzbxWg9bF1reIaHY2Bcv7+lNtVC+0OsqWizy2jcPsrTengT5DHu8yOg2T
QOfLEPYrIYLUj1g5NpdNi6YhWa6leQEZJ4Melhe8hCIOIMeNGJ990r8Txl6rm7wVVUAQyFTxtO+d
2srTzDxcH9DA7fD7IN1LTNeidRsqJI1HISkS2/aTwBUbXkxVsMY/BUf3ZI7kjRK4mdeiyHALP5TQ
Bh+6aEbpfDRan9ZE/E1/72EwJ3Gsxtx+qUTE3JOY3n30ISohJfNLE5oG896LthPcplnIwBEQjGRp
Qn50BAYX0NdyNP/iNO6sQec2o9X9aP9d9ru1ctwOppd0xvXZpurByFeO9IYBddpnoTM7ncYynMJX
baAfCIL98JvRH7CHs0EJAk6W/fgUcAOtUSIMoxXtIXV6eEI0hP/i9FQ6LUHsoFc+1xLKcqYHe/YK
0Gk9/S721OyQ06o2iwFqfvGdpH8mM7UhmffNfM94Iv47Wmut95ELU2hmhgyoJQ5v1Kv2oVgX6ga1
VvP6mBDzsJDPzd/+StIbtoBiDWFMkZqLWASm+inRvazYfhLRs3vSwxy9i6uGHN6pR6/bQa5pJn3+
MH904fjV/Xxf4N3FcK9nxw9lUBrUV8AzKTdhWUYChS4Q/rbPUMRzBLtJDKZoOa6BMkh5herRKf/N
PUNtcrpTMDQte74PhU9wx6UpGrE9rOYx5Pb3mZW+RVXNfQzOALdOL8LrZNIsHUSn33YAPa0/6kF/
0kOLvQl9grpbVjmtZINNZGBMeIE9E0qRwLDXwHf3pNHusLHq+Im+KZ+8XvuQUIVPPmQUHlITuc1m
OCyhjdmAo9CXBJsrAgwCg8ORMPA4tjUo8l6TanFK6FpAc3he1gTOmNkfRR7iRG/BB18jR0BjLc6A
PEIkqELhsi04kTJNmStoboaMLFEwcLCLZf2gfUXLc+TTlAN/Ft3K7O02q6p2KvaD74c49md0NOWn
QclOG+Msa4S8nKSAuYnQq016fWQGkuHxH+3VrB1J2tx1Dt59GSPjYQTGyNag8fHOzfhGTUrFqgDh
5PQ6CJ2g1uoj2FD6xyR9rh208GgBmTyUDCgzh56hzkgMUishqVB9zqhJug1v56wcSl1vK94ce192
L5tyfLRT/RfktMCCPR0vya/PpW+YlXgFPz48H4TeE1ULpf0eKo5alCIlfLX+3xgu9d8iDnt6ITa+
rDYDRQad86Q+8uHgtwxxrcBH/MHOZrb/rA25kfFE+MZuZHef0cgg8rfbUBmaUzR45tp5VkOYQ6tC
dpqnHxEZfqXqWCSKlPNoqQqgPq22vKtlU4XhAqTJceOIV6cskFnXdOB0brS4gN3NVdr5Sqszk8ex
lqrjPy48KdxDHt2vBY2KXAEDhVmNeKgyqyh8euvdTSH5CwxhdD0euMjdKg7TQYaHiW6UTDQM5Gvw
RzFJQHYXcpf5hwKuyUFuhypXPzhffj6jmEvTKCsbV9nKnqgzkV3Jc5aO+MG51FmmeW7Xgggt+PXd
1a3QW9QJdFIdd33RIKCxc+NY80o3HZ4pVwZ8yOHIyMC42N+k94TKsZI5/nwhwblMjRWPQNXECrZ2
0/DX4dpgKP1rwAfoPBalJIrmdrfS932DajnEfWETn9BV0wuDzZBCfrIAI+ttH2Ut7V1Z7RgJIW7F
91BN7OTdn67U+Vkhh9autNUuFJdNKpZwb5WIhZY+eCMiDmKJz88Vfj2cO7s50ZZaZ//X17nM0ARp
KnJQyxz4CqlHDVu/dn3BQd8DrHWNsfSNmsJkX9+Ox+DBFckZn4jO0BakdWgAzzEuvq1puOBFDgOt
jlgKRfkiWhXyAQflN6KrsTepTGzWXxHIhdACTo7Xgs6KDi/aG+WN2BqG9FbGfxyqXYDZVGAyTw7F
igfVQbjb8CrJFolo1GuzXiXvlpJyl8D1IjFZda8MytOnaslxP4KFn43WWRqyrELI7ZXLc9Lmz6JT
K4si9ow4TD9miZUZJSsnrl4KdXuDwRbEc0PGDEWGbP2L3xeAqAyKHr6Xzy2BUEzky/7uaO8dbVKp
7IpC7gCq47DgreZkb9dwjB0YFmofd4MwtcLE1N4xWVaI/82aWTqU1K9T4hc1PC8opq+yhyAxXkyx
mU7NV/GnGapZ4VryH2EyelCM/hVODRg0TTdfk0AL+aopZugUDPxSm13XnDkU3EUf2o0yUc7VV7Nz
tfvGSPNiJ3yc7qJ3HFSFXtfQVQABbZ/JogxCAKyG0782M9B9jd3Tt29jWf+jXcNJOy2bADAugWLn
opjHSYLteIAxMu6k4lb64y9AKAfQbgq3y9sVu17O90UmdcpyuRq9H1NI7byCUeUXxTBRGVqGVm3V
LmVL3BcYEiRSAz4567DUnSPP8ChGrd+ynmdpc1ltptZ5LngYAuFvMueuMvGG9UzFdKw7Qfv9hP8S
lVJuaE2gw5OWLOHHuNZw172t2fkUH2Xzvx7bYIJA8D1s+RGqyy+lRYhNNXHpnj3JDpAx6FwV2oko
kQKEEqCg9lyC9jPUMfm/LmoYSSrZd+P2r+YcN4wHW9X1HtUs7IiEH3BkDTYKMIEMfhdiFI2W5bby
EjypIZaNDDLhfLx7l6tTKARooJZ/BgXKBOUpxbnGyfLcbUulqDfTavX80NDk16SM096qGi2teJ+0
ZhLeaDWJLUFpCImRcR1k6HxqcEAEvX1zqIRmxMIQZTFAN3VDpJP7bYxeujSjdrgtHHT2nX3uw4tI
JjDdsPx84CXg/iiah0eVwJ/N3OYHsV8SO9vhCN1gXzcufk2hYOtX7a1arw3/nMd+SRA4m4hM9KtS
DcbgPbt8pl29D7RHz3/HsflYLgsWASDUyaqvO1/nAlgU3NV3aaTN3Ox4nU2Ph40yoB9sN3BDbaP0
nAMDTk/FP0ARZvgNd9tNINqYPTHQTlNrtob0yZwnvw26G7hwiv3X832NLvvzrGITamW0arOIpmh8
T5LdU6fEiQYGGrUTW5Gsdwmttaz6CuOs5G8by6SaY58BlDSM5vaERbDi5uD9q9wJXo1sF4lWgJop
yhuEEVPDdPpGYW7E+HoEsh8iHu+OWFBiSNPRGp6vBJU8acqtYFxX7PYchGGQDCkfF3dJQuj69U0B
vgn5HCN4YAja7BCKWl+9P2Iwv+UZbkDjMMmTTc2ZavZkvzdUD1nLfoH7dkCHDA2fiPi6MYHd45o5
h7+VylcgIMHjIBUhGFhI/7VCJm5oeeSo+/kvW8DXABjYEdsya+vxXAvirxSZCOUj5FCImof3ZKz9
YmrtqL4sq5sxBgXH1j1Htvfm9A5ekewRV/k/AlTP5OiqWgw7WprcainI7q1FE92cZYw1rKvx8A0W
kFlW49mepvxHaYWL09pTT7gTREgxV4c6FiDfO/kAnLuO2U21GvXUg3+Z8UDlqEYi9XDJ0/QSve+D
3kV6jqLbK+LpfobTPR5kg2FceF0ThLsGTBiBO/c/tAxCrSYCYOoeVfUGiMDE5OZgOvNUNJjLOhlo
W4CI1InoMjqCztTzk+Mbc4XiCoEPDdT+Vc00j2JAjRGfJeS64X3/hedpL648czCk5mjJRyclQqTW
73o8z6OX6NBi+UuRtAuvUP8Sc/TS4/cbUkeibe0uKM9m/lfr9ro9DHv0yEMCt6+ctxlB0kIKPuec
NDlhyApiXGvKgYSXqTvHuJc2MNDS04uxTDp/eL+DkYV4KzHTQDdSP9xvZBDkJ5kx6FBfM/73E3zo
eVC/7NHJh0LZnJ5udibPJnMzblY4EnlWgNMqbwm1al8v1s+kS1ROX3uPGNa6ByjG0kje4SgUiR0v
VhjS2G+YvcMnbJUzjQv4LakxOcgoFSPxEInzRnstvirq3/uwTVxgOLG0Px2al46VgXDp30Fd5SiY
8MEOGnc5r+xVQDETrTsNYk7VQ3Ev1z2il4sw1yiXsQreqlUCCH8zLu4M4HfSP9QD47pGNlr4BRz2
bQWpIL3ZuuQaBk8q5vn+ajv3tW3I94UmCuaMT21sMsjqLf3gzowG8N0V8euLy8Ek9eLrylEzz6kH
XYlNnxua5bGDIwSHKp0+4hl7VSnVrnyWB+PNAYEEg9nv4Sep/kuHtRav9QSwifEeEz8QCJsw4EDe
Bly61s6dJTp2g0jwCndF5b6V0bduObq20/SsOEGfWGuBILzjBSZyAFyea5MlCE1vKAde2aoU9Mka
J1lx21bXNW8iB23UqFOyOnV51hdDb7SqTfObWhCwGf37Jt7DXGzaSrYqXraftuYCt4WThH63udEX
MK1UpJV1iM6gbocMyhYRhAgGUtNlMES38m0uCce558IwhntFrNmJvpN4pdSrDedLYRxAXFnc5P1u
rRF07FMZMQNtKUfxnygi8hPbKZgUGU/cu+Nq9MFLxD8ceAPwhzivMd764nLAR0Ni2uU5UA+KyBMu
GfTXCqB9sXUWfKvtcOVb9wMAwtbyPHJl1lKYWhGLDI+ds/dURI2qWX6ripMwlUwDrfxHZgaNuWun
x/kR9quTJh0o+khCXdGvJ+Cwp2J3FkxHZjxv14b9Ddds5gyYbpCnr/th7N75r1Kt12QvYeA/gbau
PXnbMWwVri/zCbim2RX7/9mIhkFodfM3GTOFJpwc5IB2PuHSSqTOuroJwt9u+Jh+v1oojT2zZJVS
Z/CiCCg9qc2LdjNLmjzKiikuaiTXYRh2V9uxUIDtH0vXMSw/sxvlg7blIclZI4TU2GALerDgLWPr
Wdw0652K4fzMjqvF7l4IRC7MUawjm1pgTbks5OHGEjSHXEoblT7tFjKKEIn5jFo77zWarePZ8CM2
1j4EUQRsO1yFWWSkHb2jSBTPJNUUuqO/jCfTPscvDCphLOtKJHZM/iYC+JcgTz3edSGfJnGtw0BW
F+vFzlb3Aunt9AoCbak98Z8zEbpVK/445S33+SXL8UTpL6DAnxhpV4eOi0SB0plR2ssA5KfEr9af
wRBqmrUrTkr3g+AKkJkeIA7XMABP1bYVXChVngmnlAqh8Yb6zbyzgm5/gQ8FTXdJNPeYEt4ruuXP
RsDfJ128bgLsk6lZcba8ubcz5WNIU6+FHBYWYlrmbi+NnbrQMAOl1ViXK0AZDCs7PEoazTYYhFpb
05dY6fcmCmd3F92v9dSGab/IjKk5wO8KrF9qAXPHHjOqOi/kXXKHtFGeX2jBCfZeY5R2ymwm7M6Q
wnhPPzf3i5shXIKOqIh4PrFElnpMT5mMySjRZbVIiueLOStCTwmTRNNCk3iDqMJM9zqoBo7EdmGv
LlZvRi/bZy0ftg4LKCTtgEuvq9Sy7vdpReOmhu4sqbWKvnFhYxTD3y3bGCClPR8UcBmjUYtGZSyP
TuozRDPnoHnCvDy3AqHgM2nzQE5CsHoP1kDEmYri3v9kwD1RsHzYhly+45kkjYY5OfhBD9ZrNaz9
VF/YpkUd2GhiuNwCrcnICWRGfI3yxxQLm3wXGNaESz7RQA1AvVRYEJII1Ovc/vWb1EYpnhkEhomG
7s7CYG7kYecOsXBU3pBCmxIQ5SGKo4wHauZKKzUhaw2wUKgG68Yuy0ORJAEyomhEurRZ4kEY8SyX
87uRjmQvEgKpzsuuu1A+xzH01udvrbDF5xE+1aad6498KxApVEIDnpIDsGcih37vw2BBnccfiG6w
6M2/Rgdl58XcKQsQM/6/VZsDZVCd/DeHh1k+ee8Zcj2OtPtlk/VAIDHEa8BaYFUmhC6wmkh08D6u
SnUd6nsHf8DztH/fTmx7p5ecKbmvzzvpqbj7O6Y3RLFdXHcJP03Sj45pH5zB8nPFLzoNtI2jbfyg
UdV2mkHxcIFH3PCHih7HSrKcGiXNBEhdohmodTKj7+QulVDVkBdtQiqXMhPB0Ws3LPap6oncjMM4
DGHRea61QnKgafzVZE1dtMWEB8LIk9VO5GijDleWrZjMa18OmWzGg3F1Kc4LcLcL7qtZEFsHu7NZ
CvCf5UKqdRbKQSwO32RGamH6zjGddCw05WlB1YOBjVRh80zWRDS5QZDRfvlMJWsJaF4XCj8gJDXM
d56JW1w8ABBCB83XPDCH+icfyGcOyIKnzXkkCQLx+TE4pS5gcckHGVVNZ7p2cOeq1OA/uyT1QB1+
RSi4cN2Bjbx/8jGJVYj8zvwpW12UvRj9ZPErEnLoeeKq9hSwXRcUyhx8eAWA8iTaQDRo5O4B+lJl
mTSKkWDsk+j0py2VkbI/KqQjW3hxl116GiktTWf2eqYWln4Q5DyfGFRIByNm1nMQf4fxxGh3Ln+Y
PMafo6TnmAdtp3GB3xhveNofPRhaYiusUePtks97TxmfyHYgYtTdvL9b/mPvlZPPEVBwFhIFd/TR
2hdoCLF03qLM2C/nMRNHI/On+elpGRM9YLM9rS40rBgBfpc2Tm/dxANzwedbeIzDhnidkqRwDVUi
tbu034vJkAp+AlhJA175Kx3tY+QH5/tsgmrgmDTXQ2yshMNJ1sMpma5VbR/Ao58YS+069RcYyxzm
G/Xxd+B2g0Ot7Tme6q7h3KVgyYIgK4O/l+YjTMtvupJDHa6wqjZFf2lvytUOfkjWZwy+foYxLqwC
7h/RBS5odW/fKpiVGWKkSCI2W642B9CO2lz8GlehqKBj6oYzBiwZArQz7RduUvELLqHHGWNewcTs
cN3PkIg4UAoGk2XgJnLZ6rr+8NoxUZEG77y8qj3UV2hiEYy5hbYytb2bM3bp1mUBLSOtE8Jn4D8G
FS4ctKWmcDfcdaIMVFdlBdpcUAVcD5bKAAioEnUOJePCdrDhcnjglmZ3VlfamBZn9u089AiTg1aT
mlQLiAsmeLNistP7siDW/BVs/142byUJZnJc/o6bKtExPG8BAlyk4l1XongHgDOp3YL7P797+/E0
xEdZZl+FX/9aQbaYzcan1vt5sc6k9yqRqciprKCtSFevspjkhrpaZOlcIOARSZjmuBOPtkwMg43a
Ok9azfwWr3NG6LPPS24/ZiI7jJTo4FKbG1kG9MswIVcpgo3kjhS6TTgLUXaKeNzzProKGqKV2ub0
bxlKqf9fAdG8Jdv9HEB+8baEm6GJFoYkm0IDbcH4i0/CUvq45vRnN80OQUYsDFoLC4fKJtPb92g0
9Sxip1u93Wlxj2BMMwncNzmcEYc5EOgnpsLu2DxovJtrsf5AMmH5BzJyIkTqkg7mbyyT7MZ1oJqZ
P9eXA3EdcPTUEX6bwmj8bMjcTM0W5n24MLOLwgopVVgrN0WGFaUHGkPGtSBfHdSuGAWniSHp4A/t
4Sx/FGr2uusKExftnc4LP7lmMXeyNcoZlHQxUkig4tfZJI+Df8WjlIDZFNUiFnB6uB2a508WnoB+
Yaj4gWqd6EAhgJ7ZZvnfu2kzBSiZkwE0lFRb8eww5n7ibuW1DaoQG9AKt+g8WVtMM93RB36opkpI
Q+/KsfBfdNkhHNatIV2BKNocHJsr0ekKp1EEmqbbVeFWZyLtFyUaOA9/wGa5qSEOEXZcM6/96s8v
TyEvkRezj/nJH2FbC44PNVVhXOyEnd8RaVHrL79/xvFiZ4g0hslMJgBaULtxwLBl5erUX3+mswoh
pJ5GkXxfK6vIVEbOsuQ9+qx5mMfIjCVArYJUN+o9aLysiLv9R2RLjwM/rcND2RdI6rffwr8/SbZM
90vQ9xzw/rBP+EYQmAW3QG+TMsun/QzeEQWWYo0cbhDg2ln6Q8/VoSzBj+YiaMT9K4JLBZEC2qrq
AC6p+dJXExKxrJ9cCG5FTzMwv/7MfSYnWrU1V+VljlZJKO3MWvYpti1zt8jqOAb0+uQlin9jMr2l
Noh+DXJsFdUfug4Xki5ceGr6roA9I/YN4WJBcTiQFeTLjXdW0V2bshTBlkMCB/+OgnuQHPmkehws
4a4hfmwCQUNWAMj1tqX0D3cDc8ZLMliPjZlUfO+WQK9BcGf+/jM0tHPD065TKqFufxQa19QNgVir
ENGwZm8JNA4mTwJdhU0Rgaws2+hPtdvt7QS83tu0AafW3rindTgkJNO0BqsyalPakFxb+ILwpTjF
YBonmnhNnIlSSlM0EzoBlq4FQuSd21DIyEPO1siqIBFFsnLAqNBK0H2D6bDeJUgCn3fvvCdp/hBz
NSfVyNcnGQym6QLQU1UOAMV6aevT7oBAWxAevUM17mpxwyiqA1+aKyr93dgFqu3vXUOz0Uwh1QAV
cdg4JJR0l1ztNItmG0EvlHDyK5Q2/dZl3lyc+ceacmrRCCB903nLPRSe0kKeFPP/0Pjbd7f0cYV1
JeGTtBC0M//c6gFUDvEKfgjsC/ICq19WeEJVm2AOcwS3ksJHkR2T279Efvdpcq0fGVKR+dV1hupJ
m0rxhASqNxVQhYaD4TTtBEaCVfM+qTwjy2djR+CFFGBb6WKjc/5zboBQrbF0biTkPOr1cLQuwoUl
npmDKDJ5DZG5syfM+nAZcgKj/gpK8dLSEvzqeYXnjiIh6Pn/py/zFzSPsd8plkVtZt/gN6buJm+p
sDfCfmNcrldYjwLO7HMizteoZCpkGMYB1B6xAEm3aXjbc/IjGHvk+4LQEi+1FK9odnNhSpXmouwe
sfRNHkezhZKguMocvVTe8I6PUGwlKRtwP7JXAgkoPULqceAHqLMaAQpwrRlty+q4/LixstX+wddE
ySCURCT4H8964vQkfvmkIDmQqTiaafd8pFX73i+FDz7trWsAnvyKAYUFrrAk2xDGj5KjSk22Ui0b
O3FdRZknPeaTEOztoeDF3y/Bt/6Rfgw6gFAHQnqfzgnyX0Yr2IlIXC3g1iAYoMNc9OScYRWk4OEd
D0jeykWMk++7kzedwyvHbcbfV9xV98c/T65s5alz75sbfzNeovs/UonYsdT9PSsr7IdjFRb7TNj3
yMJjJIKST869uxlrwVwAYS1oTaYlTOG6j+CrkFrkYwHasjbvSqhCMyS02azTyqxDvzB5qgeWNVLq
R/RPwHyGN3Kvc5YiPIPX49xcBL9lvdNp1eZzyrwIK7m439GZ2xO5FIt/KAhUPQXBbjBNXQqdGWPf
wjl3i8LK4EFAtoec5+OZJi4I+XUtsHlvWrGgZUq0P2NOp9Q0ZryG1RNRjex2F3f8jogNROwyRrid
NzQFOm1sHTsgOHpcyyUgUBJCpwAlDvM+4oUSPM09EP4DrSPdIeOwyXiYcEkDg7gM0FoMd4QSN0l0
9bAMiJg2WryHT+YF2khwqIFUl2XCbhmkBvty3rvKyJAUtwGYpMEdxhq6UHR6b5yqCwpmDE7KpkbB
JhF+4O5fclASHf1qMvZW+rFa2P4JFaJrzv+j7QFa+j6ck43dLOJQZhzxkXVymLMd/p2SjxrfQYJ0
ZrVkreuiFP1lMZKi9861Q1HQdqifg3oDpFrIuPMmC5Fhry24fVBwfNb4CMT6HWHc3YOIKgLQbX/N
YXjFM7pzxNh1jyMbAItWEhy6jf5RE380vsiSsrM7uJ9CoVMoxzE+tmfaP1hd4PlQZudSFRIrwPZZ
wzT8bG1fNTclTvNrbgGOwOTk0IUToEyBTtW9a0DDeaf1OybSrCPojMyVLoVU1xAMtUeiNyhntLR0
UlXWJ8zEAPDCt1q4tW2/tQlohabfcEYB+jsJPteebT4T9l+2zFSLZLmmSKV7UowMH9CIf+y/sYAf
DoOgHCqDC/G5QWmJU6knDz5kLcn7ddXTwjGaW1Jqpl4fjs4CSWeQgyGeL9vFTYSPltb2Y9h8ElGK
Jbd94uRPtz/9zzdJkC1ANwaUx+JZnn/APHzJMd5uovlYDWBoCHm5RffyqVeOVtw7cGQKpwmOTSeE
x4yp7aSZvAg1yzAKOw+zGyRHJZnorUCCW21uAyjGt7O2l0SEcXk2dJWTn0UdT4G4dPL1h4MH321h
65tvw2sr7jOAhM7/ZawwdSwez02IJqyyW45hH/3WOcXjIb3GsGyxeMOzJ9Yf2qqrt7E+kDBc6T4y
ofecyoLzSTqvWyQFHtUv8ABRG5d/wItRWPasCIt7BkEK1elBL/BvKqmfP4m7Z6EiRatMxf9fi3uK
zZSBWMlm+p8Uchbed5d247smDGG9JqvBWFCKuioMJ3AuuRLFZNk+5Ybbvi3WkG+sBWjTFQOeDfVJ
5Elz42zNQu7SObL0cbRLLRm5Ks+e7uQ7Bv+ALSb15x9CS1i0FgIOaYcC0weCZsHXr8tTv2OgYH4z
tarejB3wX1ZPA/6+USrSyDYTIpliAhswBwI9hShFa+/6CNn9zzHuFiiud90gd5gk7cvJD0xyXeXI
09tewuD0awQMNGzQkQhrA6VMprKrcMHZ16i2QF1Ous5DA6cbu3LWaxld4fd7rYiFQLO/nvjVVAQX
Q9w5LXzwKwfah4i8mSMehgZA8T2oHMS8jUbiqTbWuWywrw353Y0J/wJzFWfj3DSFMDcuS+hKZ9lC
0RZOW7PhV7Hivw9OofFyRunvWFGOyCg0IEOkAEaz6XsznFWmjcY/FrLE6yFjH8smB9a9Y7J9vPjL
fD9OUJl+9yq2/5W+jniqaf5q4pVnrm5+DOT/c6kqPRmEBelHtiZXnEPznLxRdsEBcMGoDNgfuLTo
rA+Fv9FiRK7xNcXSPfWZnilds6azYnrg4b7rCjOHJoBVr54nnwZbhT87YwOG3THfP+qR/jZOIfxZ
arxYeFz6MN46wNVQraISh4zq5G+QpYCkeUoTsQk0uRTKrXs9hrgolX9hF/EgpEw0BZHf7EEVB+/U
UTj1RbTnbYFWT+UiVcnYEbaE7sXrDJqGqbI9IdRYC9FOGlNOHn9yA3IH/4Nt/o20kuWUmMeIhVrt
WSzV4YX/Oyqp1cDM0TlRWIe3ZQ9Iakh9fLhAwYmQdP32Vy62z6p9ubBJDHPGNIw/FgrUraK/el43
orl5PWaTZYNcMJaO5H8qgvMytd4jx+eqHyYZj83ii9msurWJVtyMuBxt3SafjAWV7CPerYEpedim
b/smO7b5sfKsMz64Ob84N+U+7NWd6EY+frqiapYf1lZsppobzK8JPoQoXrOdXUwmpD7fLe5KfyPx
r5ZQsUM85SrL5GIBcIb8uOT7S+fVU7K1Z6PA/zhRmaXaELHHsHD+1AOSepV50/0zyVedpzs9BIUo
LwBCO0rsoR229jAomXkCWqySyAPG/eJjeY6RKSMd4K6qSLopCqzlr1SdCMHhHLrbXws32oBfP8Bd
Qjv97gTz3FN6RVqMh6oqLdXs6DyKvmMA7hYu9ktViwM0dceQPwvGYf8rFvbA8HgVkh5gzYPCUQoA
El8cmDAjw2glJ6i+tYzQRbJ+3N23YnyJxv5k/gOf+FmQUSgX48mU0adGc7Uq1kSQBKvTK/JuBwaM
00LJt6d7QjhBFoS/1Wf0gY0dITvSWPA3CFM7IFCl3GlqT+yZin0jXtSlXHyBLowtfBKsDXgh/cDa
RBkuI2ReoTSUAXX7SRMOrBx637AotcPp0IDvXkuXStnP9ZZThqQanxgG/6LHzID7vfZm5xBdvK8p
B1u79BV7iBGBQk7OYKy7UPiL4jnh6TnQy88SNdX+QDsDrwETYFo5avQ7RKXQ/Luu5dQEfy8s+GFC
y02Jwl6208lMW0sO5kRS5ttynNpTnSt7KHU/fv4pWUfP61dTYY/Lo6kEOvcITJPuiJcoTEHTmdS2
TtHenZrzoAThPJTaw2Pk1zzqbwWntJQDa2VsDsHhwYA8E6bCJxELplHANU2rNph3EG7StO/Jp7hc
tP8iMC5/qOEEfkoy45BXO/w4AIMZvoxdZcuGQlWxoQ4jc5xXZVVMp4RfpmM5veOp2D03SHKAqdGb
Bq6ETuXu61+wNzKwtYjl2yWIkYl3qcVcLKyn27BV9CFlGwoKS7EI9MZmVJmrgzg4/dp+Ya9HL7w+
9LJhAoJDPHnVCyThsWlrp7vK8BXTz3uimXgGfALd4t4AtKSDEXthdroGUyRPrj2gz0Q+or8Ore1f
wkvuOqzVmOxZDvi4NXGaAew38Lx4/1o9/m+FDt3war3+KHuwL7kJQ3DLD6lTqij4OynrPuXtawfo
lFENmZoAIH2MXla0+AtZS/F8NYGuT+OJ2PiizcPVDft4h2I5qFAuppSU8zT2wYdi73DpN1qclh15
wuQNUFFGUWbiFAGua1Wo6qlOizAMYF7m2Rw5oguFRP1muzcXOBj5IN+0nsYOoJ8wjpKeosMrEyyd
c4GnfmoAd9JhegbzSAkF5eKgJZPCgslxs+rYpYLMo3/qYn/NPNirv+EiOeggF32nhdzPGx+zuEEM
MBhhBtU2LCzNR39Td1QlfTtc2lxcAkImhRH9RccOJ75hOyYoM5MHekDeFF/snTb2nm4gJuHTgKI9
NObQMVPac6iE3gI6XveClTrPdlZmFcbgcPV6n95DfGINGvtOzlzESay4Ru1k8Uh/PX5JRsYToUy6
+FzNfHzbXpXat7R7M2nOfPjAX00ltcN0kaIHse4gSsHHH8Y2v0spzmNLPOY06I44qh1M7JkpYy/9
NTrFO8Ac2nF8ea4asmsw46lBxCUFSDSOWC33JJ3Bwq2FgdvRoS7kezYsI8a6LNE99Gkhajxk+auv
OG+I7Ewo0rDXkTFsZQIHJrGq1vlHzr0dE8hIAYp9AEuk3zRNmGsNkDfERye254zXM8ZHOg3eBIxN
3ExNQe72efv/8HIKKYJZGuahv15R+ntm2+q2gRm58kENqrNjwpS7YTIUWHsU94S2gnmFUNwIQ0lP
AAB3lJ58vbkNNfM0wz+geEPmRq0McCzwHjQSFmY8AkF5nYxMK1zr0okKj46KEQatTo+vpbyvJxT3
b/4jCvHy/57ykGreZK2BYcAmmZYyW3gY1WCZec/mbvG7OeuYexMTOeflgEmmqtZN7Iu0vqqpj8Kl
3C+xekUwC8RZ+SgEOW7YhVUe59L5S8iR0x8MdnzMw3heD62j2uIFKO6DAQLOtmqgQLykAoPThysy
s9ohw6epuPAVzesOQy3bMkd+MUPTO/oqXQb5QBrGJ7yrUYZphR4uA5Ug7E/hZwXx85k4nVX9w9kY
69JdtRuBCZZK2XgGZQQXxbzvfyCvFWtfFqV7pwnVk6ASHirDk9zCTfTm7Vx/ui7h6tVbzPSmzZu1
wqfm11f4GhB2rvVRjOaQv3T1D7kl9LFYzUS+ji9odzcCs7pSb5NgupsAUNKuBD+BMwNuhH1UzKk5
SXEVzbN64G/bRWyV5tAdYsBhNlf/uEtXJ2fQSgXc8AQwU9o8aBTGOaYq/jJrz7DGZNwFSGvRDBrR
h0D931OkMk841/WyNYIKntuYgd+0B9RbzU7ciWyetxiNudeL2koYhLC3j3ye4UndWfCS78vZP1C2
+/nNuTwt0aFxL89Jfz26RHb8kxc1NprDFbeVkVXJB/lMJde8hLgD4x4qYWko/lMk+hDPM3PzC36t
GFqo6EtT4d4q9IcAWMj6clAtXy16hHc+RlS6ZmCDAGRyNXkVKI/Zl7XbqqqJXL34gVeg7q7rrJkH
6l8+2MNG+BJP76jKmmXwuQAV7mhw1gAqcvglfLDUvagy2BoqRU+IMUjbOPHvhx+mmAs2HrmWEygg
3FrMjImtAoDKCeBVGZNI1nWTGNrrrbRLnHoqP6nWNrYhbowL0ilE9xb1/Ma8OuxAzffU+PpYnxu0
mTfOGMp7XPPY/foBTtXdmIqZjeIH1ZNA0XntSZ4tqZaZ+nFGX5O9TLQccvD9jPabSdVsSvTRFxJU
Mk8f9pLgwQxcVz45T5VrP94kvCkwWOh3H1CwleSKSbCOh7sgEO6YXeYGs6mxPthA04X7Rgrkrb7u
S+EVqSV5/LPZVy6r+2+hgSwpusBQh0KEH4s/NDXDwcytBzcsqT0+FzvlXeOjnYcwHAklkZwZeQ3O
WwzvasBvDEIIsHjaUd5dc0IE1NO+oVhHU3RBe42+aPFSSzdDzZp4VLqfIsZI7+b2kzlKO/yZEfcp
xxn8JL1paFT9zcudlSvgmOGIogzWqP+HHuaG5yUqYCkAHJgS2kl6pAqQ2iKSz1fO9MYELULeDbVg
agpeCMZG2a5+H8w6dDm2VXs0ObSeCEk2iztXO5Z5q0bQAtLzqH/zvSSh4VefSd5CPg6tOF1sQFaG
zmAWjerICNTj31TwN5MmxBjHhmGzjbLsnAhxAKbb9Mkg/5IHxg9WCUxaK3GMhvfKAefpHe7uQYWF
fVUqKEXdbTBbGtPNuMMW56gf5P+wj4xkSL+qpkpr8mXmXU4Y6rByLZqp6RzhRuz8LbuGnl/Wx7Q6
jhqbFQHcC5Mv45Z2GNBJRk1ACYNt+fzW70sx9YWMRh89Krj3iLMdT/4VwlPNWFwhMkqudIRITcae
I4zWB0zIcXmHIABZ24HA/OdjJklOtBYLd+B88lhe29U1TzZPEdM5Xo2uT4gnkOG4E2JCiNMZKeHz
LiJiVmO5Js4lphiGotSh2OVb1ByjJ2vvxJ2UFLQNLO9+4zCAaUEFhmN7E4HF9CtLmmvS4SDT5QWT
6ygEFeQl2KI595h/8u4rdj35ofc5p6WbjlNXfsC3ADSwoiICinYndNDPlzB4MhhFLnMR6R2G/1Cf
c9cXoCDCShCT55EKj+mMy/DPgSKn1uDZazijAYBItQs7yCQkHshhOejwUGSuVV15xxw9FYMd26vr
5RPAPixGxPU56HMKtiwIR13zSmzFgKD1OU/hUCu/h2tWB0kId9I9id/7i4evaUdxGk4/glXCOYaz
RzbNKZHGI8XORkiLsyqsSSiHNaPD3K1qr4VZ9kCyM2eJDUi1R4/mf+FkJp55aFet/lYJU7yrNOL2
HXhHIJ64uQbFxnv3kT/f4JjQ3LAGzsNs0G/m0rWP3veYz5HNpuXOUP70CIjCouKDdgIAq+NRUWf1
CrSzA2V5dEM1YgGjwSulB38WxO7IYfZ1IP7HoLNWQPl2PReXnK8IVS/8EmrFXqzBodM74ylNlXAT
zpq/f4x8O4FbFDovDjMgYG5qx8CZ2p2qW883DTgTPqsEcDkkD6j7gA5ZnOCByhTwaLN3UHf4f0VD
6dnYMGysMTOOpocbSX/XwrQa2LULmjtR8bWuIK2Za3nWQ31TkL0JpGH+LdeQ6AEZaFHKuz1dkeFW
IvMo/vvGDMokUvRxs5cWJT6W1V9vvbQ1zETonEZGlS6uty8qqWsElVW4fTHj9NVEWfJhwhyzj86D
BxdxK/rrUvkCJoWCQBL1CPmPFvk38VhpLNj9tIDC1f4XhvfVlYtQeuUDRFNTetg+tFey4anIpvMG
5pAGllew5MSREPQQhKdV9SF2GPes3pMhBKII7XN2AOz+GTGf758q0LF1wtod0i3YbKEPdQFNeXw9
SmCnh45TmMJxVXqmxO/Z1zKrjLbFtN3qO0OIlBZMmF2HGH/Ub3AD+GBX9d+NMElRWCGzfh27GalE
HMYSEfyOHwKdwILTqMLa7gt0I8EUDUVgyt56ihRbBn7i4UIz1HJQbntNNnd1pDfW7g7/9sf+EQ15
Ppm0pGL6tjZVWboAEhuUzyUD4qtu2SYQu+3XTpCKyuASS93JlMZ0Xb5wtjHMownGTOk3QsuBeq8S
4DmtDgBVKR9hKig5N2liEdOQUpdWZXVLTdP3bI3kntMaN1x9Mu6HHF07NF+quefpLUqRBfQerGB8
VcX/GkarZYCNS13jKfATqNKmobfyLur/foO8OAbHgLjLGlFW0jHsQmf71NByy6+ssZ8AdpL9nHU0
lVP3h3hTD3s1tWGaAG/60IlOkk7dFATswo4MOP7FtOipMxLfXfb6VFQ1ST2oHS4iiuUlyCzQ9r2P
dpliWSU3spiIlAmMZ8QxjPP4eZaSR3guYC7qtmrKeh/xte9g7z9wQ/nsMAvaNHs9ZiPrIvEnqY15
eJC2PRxHNqKBaQyTcmBC6D7AhYaBw9jTzvypcQnhL76AtwjOvvlrP3lzJkWzodRMO5jKQmTmiUEE
WhfwMPVRPSWUNI+Mvlh2OY3+yceV7sK/Ck9NOXzdph+cues110Fd+VtdjhX5diblIfq2TS5b8Xx9
fPV/KyySLoUS2E9foqJs17uNyer3W9W0WNFtFLSG62NkIcrfMoIxrcwBgqSrsIjDYhf8F1Vwvwri
W4Ocej/c/ZBR6vHs7/TQS+r40upHrTNiKskLSd9FIWQcMM6RJFNujF0ZgYIup+OO7ZpTs7h9jRck
J81GDLsnwC1tRBKrl9NblPUVA1SRAUx3M5coZlONgud/dQlHyO2OwxKnQg2741O9/nqeSfNQv2hk
GXmtvV5zv02eip7BkNGcrc928ZdG0/i3EsBivg479hj1z/Z8Yss9TnfUvJBR2vXYTWvQMWCMHq4a
fA+hB/s9JsYaJUuvgRcPMeQrl6ThJPH58+HGRbIwScrtksjKbzYD94M3U2oYjlE4xYQtvLCh295b
9cDsd/FtqwiI4hZ/ChEgzWIGX9E+PMws4gWrGklknP/gs560CMtOxRxmV5m4MnmJLaI2FnumQjNm
eR8v1wJolFV2c74gLean3bQ+gNwq5ErCFR5OeQnZQiF/iC//+vJPslk08xQlRmgOzGNMRow9fqaO
vNxmK4KWgxYj5o/9TXbdIOtvtzxrCFY9qqOctZiA71DTy2J8ucIgrQ2ijz6K0EeYy9Ak1V3VcxFP
4psTu1YXGqCupL0qVsUSmgN83RHEDFh+AodJOKGW1HhVm9f8xABtdzHG7ex0ZBkAEm/jrJ2l9ng+
dUx8SlQ3VOW7Z9wvK3yxkPNu995dItd2GPjjSAhQDvquSDo8qyEJgXfZmvxNr67gy9rdMTC/gZ8x
wVO+dhYXtqaa2Nt5Lo4m7iKpIj7iVnOwpprNJ1gTrgVbAhuh3SfkWoqRjaO0lg5esqLNrKqQBF4X
FV6QkpD5Nu2pQMbWak0/GaINYWPWjlbguW1ZLZ+EiR2GHgpGI5XCl1NnIh2RpL+eg3zSMT6pXB5r
7UaGXWt4N6KQazPTn5mjFgOa7tiidg2T+7VjB12QbKFP8PJ9ZhqfZsCwN/0wjd23jDS3DGj7rND4
dQTUSjNDO6LqbSj1Ebs8nwXtGrzIjAHvOyRRZpagzBHs5XBAdNKTKinxZNmqSbXliiz70V3C8lVv
f4zWPyMvDg8cAY00d1w2xoWBdDH2XfgZilov2eM2pU9bUwv2Nl8E2M2c+Src+9wxb85djqbzjvUY
+iKtLOWy7BKfxWa/i90SKhbw/kn/auCkOhEHxPoN6XJimHg/HhZCviNjWym70Dz3FUx4oaf86LzB
nBLKKoJeerZ+9DsXEc9FdLYeQVKGzro2ws7b8L08hXyCyUEgyu8jdoTdV59c3wFeMRD7OOsnMhhB
MQSaiF8U4HqYSYuxlIPo1F6RGBBKAfhZRXO9jmHZMgtQLvyeJQ9J0Yrqt6PY03tG9T6YELiFG8IM
vBrr6D4Xzvv8ojnk1LNCILBGCvinwyHWZf/GlHbuOL4d1nQbRAzn2jmf/ciy8WtKORfNY4HuO82w
1si2njJhK6LdZnWCBGLkNGieDZDX/AtL8Gam8aUdXDTzK5+ueQNUywq+Ivk7i6GMEvPZGzuevM4r
TUWsdhENcNuTn4WTQeaQ1KzgB69H0rLWlPIYAS+muTAJw1xmCK2vG8nWwVFWk6V7kmIp30Sr+h1q
GgBQty2OwDajKY+cReNbGh6Y1zlYJUm8FEs2rkUujz6FLnVVuHxbQMe69+vwR5Xs2Nb2H8yeXzjk
v1GHQYGYcqf893+khgp9WoPsOR9ykWHrsdkkvxA5DS7vMiiFwOssYBy3C3nQPttDsYI+Mkdy+mtZ
/eMtCM9G7pTzt9fXUiA8GIwJEFltXQWNWZFRpRjGWqc4LyACF004m5lRMhylv1TA1XPbQ33sIzDM
Z4f1yhzwtUVmJZLdnBVBI8oPIMpmS62Ylg4/1DdoFf7yivJ9S2+hmlBit3HNqbkpOyOnlZDuzJUW
tSVaQ1CxWh0Hvdw/ZnY3z1aKp8AL4R0BuknjoMCAu/dtjTcqzHMGwHJBATQbfTL+JZvioYwO7x+o
0vwKK3Yf/wl8uJ0kUWBDL/gqjCRM+UtXXCt/GvAjMNrHOK+S3TEvFPEdmPQoadJnmvCrVc4lDA3t
yoVMp0bx+/fl6nDVhk7qE5adSq0jbVbIn54crpMkyGiD8oGkB56ugUk6uhGFmvZRG3VMzddagTOw
xfJc8OkWy8Qv11ym6FU2ZVqAKZIr4jTxtakTp6mT7YFWp74zqfWqn8rXnxrc+VwAZVuNjIX4oP3p
SWgo0YqSkAx7yJB7z6AJww7NBICu4bhXGevJBVIWxYyKvDBxr6+b1GmD76TlPzpx9ZWTmSnactXG
VBMFLGMTwwvqe32B18NbRPpFz+X7i4CQ8PXQ9n0Js20wgufwuElEmiq7JSF6hHh3tc93QbAh5M+/
WwyiVp83Z7KX/ZAbxKwn/a1KSfXG/p3ZTPcJUCFl1TcHlz2x5nT3P2jRY91hoZB70vVYulWo86Xq
dKBAPvDf4zM04uMDYfa7d1PWX5qzckkR+MBFJxe+k/bX6HQRasmjl3xU52mSNRJFdRFvWpuSuh/F
KG6DNg/Azwp2YfN8HTs2dCuqO1zNJWs7GYAJ25b2kK7oIr5Lft10uYI9rU+gHb748jx8WoNjVX7x
hbwm6paFGBA5dNQDagZmBxeblxmhMfsgmJ2aCdrR6OU9ZrRUSBaSGDdCViZiB8zx04NYp1Q8RQiZ
2w4XW1okqS4pzFz9qF7FihgXsjeACU/qCfR2x/MZvXYiXNoOwYGLcBUsr6620JU3aqTfWbLd/gRN
rFZzQH10aZmX1fGPJRb7QjUVh4HGoNNAUAUIzkeLd7JkHj8epEMKd9NfOaGflCgvuBk+PXQxFtj7
+HIXJa//eyD/iY91/vzejwQ3E4FUOPlrx9tJLYaqaMoME2NSAZ5qU/M2btjmaE8bdm9mIeBLsSxo
oFuxlq3ztzuq78Lg9CWJsavV4QGlp2cjnCXaBj9gtjTMbKJaa+vSLCG2giIjaWuf+mfe9+3Ha1Dh
Lr4RPzmPpeqgEmQfqoa65WtU2Cm3rkKR56ew75hqJuYQvPpNV8uaZhb0BGX7kaRz8SuB3aMmlGIU
Ti/nRbc6XagrnmSL+wZWsYtAbLjsmCQ2MRv/7+ygGGAbLKiOIp8ZwLgtbu9afWJdHVHtdI4f4n6M
pa4FMsupMGdV5DBB3JDNNIxvEoQ0NqclRINeLd1LJyT9EV6MMXO+SDEl6q/NGt3dguKsNhIgSI3W
viNURce6kOa92ZYMoUo8iYRPSM6Nx7AsMax7V9HhXcjUJ4Auap8T2L3Wga4tBy4fD/uDgpzql2bZ
ijOO3907Qh3qTtUGCDC/JeMcZyqWYeC6hInourg8taHqS4WoDRTNrnXhC8b4UdDCOM+GoJ65zvYn
JL6v2uPFItfinXCMsX/LTQIO2GED8UuoZvSqQd/V2Z6Okv1UtYSz0btyK35K0wZhv3Npt8XWE98P
uxsTGsBYvzelRdu0c7R5uGJdQAH/L5/O2y1kmncN6CEAy/ac6UjqjFEleWchH/ZDVuZhEsJLw6Xm
1dHss9DYBe+Zv/kpDRcXpw/8N/TMsS8LnmyiofNe0Gg8EWS3sGvhkViaFJ9shOcn9yxKn6WNznWN
zw3IbQLCxEvO/aKXYwQ1lEuVy5wkgX5i7FbbYR9UIm3iaxBp/MVdJIwC2B/DPhbkg3qlcjnW4fVE
t6j8k/p3WNHK4ZAdSoUf9YKiY1Hl3ST8cbQdaYVjH5Rh+C9S1ONQTsq+LrYDb752Am2RBq6mYBkZ
Lld2Rb0EKHOi5FHOvEcqzioD8ZWaxtkgDrjBcXdoZMuRdG3JruifHCe1Nm8OqTdiBhHM3nV0aZha
PEJ/9Kr+1J34vCRbJsAgULx8Tw/oNYb3V9xktGDWmk5DIz8DqZpbdDM64X5+MfV2Bk/hVAJWXQ8u
/yBtDjuPOiKtaDqBlhKGbDtQf3fF9ZEQISHohmQAxepNl6a/qaISStvW90r+9kx4oVbJE3ysZqE6
IvhnbQS6etS1kQ/eF32LOfuskONpKGQORl8iQY+I73eSu0gahM4BSD25PsuesaWKshpRovihdkee
Q03Thtfinesue+5lAsmnbR3LWfxu2vVDxSMCOEpCyUTcWi+aTyvPaB1sMdwOG/uuj5XDo5y3uVHo
tIzbMQTua4H11xG46WGWSdjMSNw6iM9yrAckfDHTxJE73adhaSAgYcGCo91OQnGgBuvnD0nE6B4z
U3fZzWFoXpBxGDZCtxY5TM6P1+wbTX0Yc74Zd2cQdSGduFwF6FJah2oo2nxo0z+Jpz2V2I4jR9SY
pWBvh6fZvcjzMiSgw+T9NEp4o7Q2SWwj78AaAPGtTq5Rf5/RB1Cty7iSR72OkmS0keEUA2IATSmJ
Oo+pxUzylxnUbgxLfyHdJyf1g+y/QmZImiAU/9uxyXFJeUrlRoZ4HnI75NzIlnU4ZwBAnv+lsG8m
gK1QJ2b/mj5pMzi0cn0WFn0LvZTcAZP/bDS1HuJRi7b1fpqqynWkFjMG66quRvn4k7uYH3Ixh9TH
SoyVLp6vxd1osUu0Zv91p+jVTA19ia2YcRb7PoYzXRReCaZw3nEs9+yPgIp3FHIizHZNTZyZVzU+
fUCdSildlcWDIkDvp1X1/5HJZd5Iyabzaz8P1A6l3jUgWFBKg5DRYi1/Fa33R4UUbazNzQBrJ2mG
pLWNfosCLVRM5fBysfBKWk76MDfVyfM4oDpLbrWNSrQ5gGzeHx5Z6iP89o+RLOBisho6ukvBQ/HS
Jwuls6UkklkDdVdoz2WhYhT5Y0iGJfhVeMj/wi4Ekfdw3M04kLvUfN4akhGLx2rAu1Hhg8xFmMqH
C6dMVdc6Eny8/BAB98zh30IN5lr6YUcqHYc1IinC1AM0AkddfLLTeQ9J82eb8Dqg6jv+ArwmU3nR
lyZhbvTbFhDcYWOFCOEcvNk7zhbEuDuvsIKrmMrevexLJcm5GJHaALZzPHV0orsq3Ft7PksIlFpE
JpYJlVVKryzppczLElAaCC33UGukP0W+yRYewJA5UtvClq+Vh/jXcmMJD440YB/If63owhFxKWQE
3Wr9btzPH1oKMkFiZ0XxpScNphK+K5xQKt5mZdSCdurrP58bo27G8YxDTrWoF9NQJdNle87zmgAA
wtLhNoc7fbgM6nc4QuFUABxf9oEgm8QVO6QY5uz6XZ9H5qTg5oXTRcbWotcNhUnimoaN9dtwF/o8
lD3wtgObN9j1PxtzpxmsIbYp/Tt675XjkXy85Vfwml0YXpNihg9NmhRF7txayc5GEKUx46t+bW8w
LgfbgWrLuRr+yBbKY0Wv8qayTPzZGOuoIr/how2IHk3Vc+Nwtdo9dl33WV/jCc1ewB6bd+DoY1G6
nODCTK1n4U1RSSXbtsau+M04mtHMWtrMlWB7Ba8JgECYYMw7WeVlxPcWZUEo+wE+quDBGdb/qMDZ
lngMKUJYPE2q7FqI5F3SDO5Lx2PWxL5gJIR0asnr4Vyg4Qi1Ar7QLlkHkxUBVNdjuD940xyNlsUo
OCkbjnfyk4yHNFMmzoBYM1Ihr6/SLBuy0wh0sSqWu36yuKGouO5VMdpYMzf6HJ58dxhOw1RR/s/V
zwh/lElbtiKaK7Oi0k1Q/J5VakVZ8sbH526tJolAq3VKCcAO/tCy4InDhLBukSkMhWGpAq1JlD6o
3z09ywy4Smy12pOtx7dF5xbRgfUqfxgifMoSoWj4mbalx/SkvypaN+Fk+dyMnm1tSXkc7jFK2ymC
IugAyrJqwRg4h9m9KXCyztSD3FClWmJY3+2i6yMhbVyxca2IdbRd9QcO1EoXQtG++kATMMjzF/pb
Fnl75cSLqDI36PkEgosxpMQGd6NCExsSUDENDLE+VHrPmX9mjtvp06xCts7oTpJEa/bgEhGr4LH7
iG3d4fmQvllmMYzXjXAINzOvR/3VBf3diTzsoTAQ3aUs3wRyNg4N++mZxK0UJ76lyDUfWpKUfdp1
ckS1m1bMpZJ3UU+dXpP3qhdEgc0yqclafziL5GhpvhoANq45UOVjxJaDlj5DB2XQy3LHZjflL4QW
39/wGSgI1G0qvnUuwJKEXzlPCphFg//jIGyo4dk5cHWluNQZ6N4NflMr/rEEm7UFr84kfWpBrlsX
FWPh1jtWc/sZ5miOIgSLZkuL1a+ZItR63BOvoGp+UIQ8cg/w/S3afoG+US+yDNncettb4+xxcL0R
6vAcwrOmEkQJnH1KZmo2Yea194G71V/mXxNpAvh8FZCXfg9RxWUJXYAi0++XxN/pKNVQJDF0a/YB
ONXZxZR8IAs4ziS2MTYsrJNUTDRCj8bDJRPxU1PRhsQ6PLfbzWwkkJiRk7q59gj4cUNp6tFmhqXr
y3lcIsE7gFRMLz9llS4DWrGNJO5026FMeVTky4pZovy/CsBmu9iTL0GnWx1nEaLbf9KqAHQrrfmz
eR++tRRfqkwAy8/MDjnYPOZTF50dBWdPcKs22Ov7wSrXELRlbcSk2t7GsBQ8AZyQM4HDMEq1rQVj
1YBbOJ45YWzTCz9COkeQBGSDb6Z7RtTBfWfIc36Id3nu8M6hsNDNZEVgOJ8hvD2EB/f3FINlgJwu
WGK/lNvyJRzi08KrYCHpCJfji51w56lrwID+gi2s1vDgWpj28QmBhz4dhYyLK2i76lwFvAVwnKZU
0HRGoDec3b7jpi2pcrXG6Ma4L8tpH8AaOCH7UgdQmBTmXbEBWBNc+61y+wXZixrpekUbKR/iObyp
U0mfcoE/YMzGYVIYVlJC2HYbuvgLVjLie0pwF5kd8IJkKxeMQ4QAdmrxgOA7S4qZlhBVUJ/VPErD
1KlKkf/zg/SzyKWSdcfjbpFPtnq3drEyajSxabTBMqmk69JRL8mLOY55H4zB3a/HTuWKx0dNKw1W
uq9pPzwltXx3M97b3W97KYjd7bivKBxH3R4FU5ZkVxsKqC2DpETYu+FPHvW0abpWpolGlHkZcoSx
CY4lJ52aoXr9XkAb2dlNHXS0a/0rhKWfuaSn8ySIr7sm8GOqHA0Lm64a1984ghiETUCn4uHJ2ctM
3gzVsH+cibtXSC7IPFX3Z+0aYCA+tM+bQ7Y1fsqn150+ElKwToqHrELBZJ9es7PpB9sDBBmMxSs0
R69f7aq2bXZ9oR7Vz2JWh6DpzMvClg9xDkxoiy7tFoP9jH8uI4X2v1HkKExyDtK530I7A0MAkyVW
jsNi2C4ZG6Z7dhmMIOuuPfpzPF1XL2FcnRrcxGMszitf7YjOAC+pmes+5i+ume7GzQul/GRShMMQ
Cbiz3EYC1CO00kKunjZJKIlK1qEdYuT/Or7VEAzk9CBp7Hny7HoUYjMFiz+IODFhyeBtrAHY+nma
WocaYhgT1MCtqRVDStVzNwCdlq3oZFBPS3hbMvh7ldSD+EAUnJ5P+gf+tLwo8dTvJXoYtTg0BfD8
NdEz2FuPJVQIBqGdxLyw2FEKZw02kK9tyaiYr+V5T9iY6/MMGyNDYm0ivou3ACRovNurk8wNrtfi
xS3Hga8+Xcz83RteBdtzcimIFcbrRip0HzKK1wxYkl+XS4BvwB1ubpo4R4hbWYeOBsqazGD8B6PN
poeIdBbl74wJhvS9C9SiojnHW3EW6dhar/06gTpP5xKUVsArrca55QuCdbp7tCVZfQ/T5c8LGPex
V2tqhUvpiSkq0FBlmSdkwi5gJNA9Mypa2bzZXtpaZ7tYCC9+ysjsG++fmlw5YVU0jWfxl9hS2PJ/
zTcPEds77ceSdf89al5GBL78G9yHt2y8hRciJNVDL2GTYFcdHHPZuWDKd/IgQ1PAGcRc+ZSVR0G0
B2zbLQToNBSK43VbCLuThs+J5magfwzQx4VbdgRAixUV2xaQ/5kzg76VnQniUFvQQyr9iB6CsqoC
pHtEeVTgKJmXuY3RFyHr3+2OXd7+Piw8gq/3er6TPJCGiaAxAn71Hm1NVgDgKw8k9p0dXS92L3pD
ozQIXyUMejamO+iD0+ZKdL4jPNOEd8oWtX/WQTcMEhOn23amMHndmFK2KboswwFiymSHKIAMGe6v
N45VGqMBiYhsfJGnNhiWPFknkUPBnAxn0MNRqmVur7C0TXRWo7fdqUzB4hNRgUWTw0ifE7kc5ol5
BX5XYaBYQvh6NidyR+YvrYRtQjvDPNUCvoUSbFBneORCQOqxXKlKhXjud7IoLxwcuPnXWC/U8K9e
OKLSN4Tb43MdV08zG5BTaUhem5V2nazKgqmauhKOA9UkFproN59/RHMhFw8lnVbOiQ0K5ZxXhTC9
8/TVJ5N8AdEzVLgadlckmrW46G507a228MefTfAkcyAgFdTuIqOO8jTgv7C8sm+JCbYY48c/PGBd
HllsAlz+y9pSyq+wmM5qaggb4CWTj5BARByVpJUyDBUFNPvb+bYhh8Z+nyfP0O/pZ8g4qr/Rrd7f
fYr6Qw8MSqwzp3SnAbCoJsVO7jW8IcMII9TY0U1Okh84ZeTunStmRWPFAYS1rkRXwPgG0WlBzpKj
o3U5BEEmFqff2gl0F/bJvpgPLec1baW9zisUzVHrX9MhUvMGy29/UeslYIQtxPUskXHJOBfuIvUn
It+pRxL90kNwaelNyhUK/TnqU/Jp0moBvbylSwUO/2Tytao6xWD9wEF7AsNeCBvIApXsDfQcQ3a2
zb9I7pI2mSz4e3H2GCNxaTJVr1j/BQiVG0ZlHBRoDwVWBO47xJC/fIrrpRUZYvUwJ+80gLO2/ECq
B336y0E4R4Dm9HJ45I0cYcU3hXJj+ozW4YrIusNKV89SWzeQ/pBdS9/hSmUboru7Lt7oVcV6cf0v
BXr4KK9XRAC73ec2XLVfL0r8H5U83nU6CHkjkP4EPaXKuXzvElnm05uX+um4f+a2ZyIK/Kukz6Ut
BJFrXr8iIhmaXGdpqcZ4bDkrfmuFkOHTW76rwGT/N1qouT/TfdHkMn8gcCoCwAK+vDBQJD/Uf0cE
E6D2kK8gcyi4QGo813UB0ow4zjbOtdJCrCMTuN1WArDTF+Y8ZU+XmjW5M9VlJ4ZqDGat8MsMKsT9
aZh67XWCHQT0gIYxChm00fjPrPWTeUjrZD3gAmb7IxiqCUjz69sZlE08jwpgGGw5iDVVjBdYrIIP
ZUbZGd747kdNgfr+Cnm13XvrI2ffOrebQFczgZu6xD0wbxlcLkEHtEtdbvYB117O8NehgZWYQlWT
X+MmdATdRXhT0SkgWBuVfzx1PC3H47HHl41H3tbSiSLYHQr0YmMrxGmvCQbrVK5sHX1Ib1Euie7H
nLCloVHYvjiPPqEgm1+l0zoZ+CEe9YEd2+fE7Nspl9d53qyN40CvTwWTC1hEkzoUIqpO0aflTkce
1PdefOHfVqV0kxf0ukFzXjtRFCeBqNpaw/xcwZBa2DtaGnNVNyj2TjUwwozKMUxCSVWGY8fxkIq1
1LeNXL4NvlJJ025xkqi8T2nE5Z1OD9NIacUZyfzkWxDwSOjZVcB5z6jl1uhoTRoYs4xr7ljTIzXY
BNPfkWpG2u2zM7Yly7uxcQUIfIsNYJFFqVEOk9BoU9rSmI4XEGpSxwTJWKD34JMdkJ0tcvmLJfFX
mtAYHhnCPlbxT0xoCP5XygxlFlndaJ3KYEbNw/aIuHeBqLUfBjxLpdO4v+r6CJxZd+qyAQVUoS4J
x20BvxqXxIIf69M4XL0jpLNcXtngQneNBgphRFERRfxKphsa/wyfcxp2iG1X7c3ENujOvvyIAJOc
cODsmG5MqqSS/Q0veCzSH5bZDl7r7QKL3W7U+5VHTD3Nno4ctcmhpmLze/Q47HX8sV0xkhahkiQi
1hl/DiFF1BRbqbe3iSx/NGOzGyXIhvdOFel62uok3Fl/INw8B9mzpic8bHJ5kKeSCNXQAsiv3oDK
YlwZLshZ4CC1Jp03xMtxK7FW+S2VEv9MZ/A0dGp+8wI4fZneYcVTsaaGbSCb3tAg0T6WzFT6Y3Ux
fAagtRxj+ixCDjnpxsh6kiZTaVwQih2HYZ7RlM6//F9orub+IIEu/gWMwURQUSdNTYajwMdJeiPl
ndvIw9IgEgRV9TyhoDxmpVJV+rzA+Usd6m7PBaYC2KUOypeORwNJIxDPGR+u4tr7I9VmnmBtDnkC
EVBcaUCVLxPiVjZORvEN1wY9BrmyzEV6mGXVamLolG/V7jUVGwinrt2QXj6cGLYlLdVfWW4GELiA
+hK+SoEYb127BAwoQua2UdGtOhaLvxsmRkvNkGe701cJIKkewFGmZwoda0ebDLqPUm0xkewVuc4v
udlMFNESK0qtaGRFh/kkq1fkjSLjKAhxi1++AxDWj9QcuGLX88GqCLyEIKR5NyX12xLgo1iWtxHe
VYKleKiIRt0bFAmUgzCcWozSbEYwaUdefILDwejqXfFsJzCeK27NnSKXjJ3aOHm0I4WnUj41Y2fr
aKbzwspxlOwUBHd6KrdAe0LlrsDmbXrtxFGBcNxfxF3aSJXMUlnZDHwJKcUIqP1wMwI1uFEERlZG
pW4buvJeJiz28899lEFHQs7lraWBx9Oj4BjccCg3MjbKMB6kys3Dt3hwctopx4JEWlR4NOfl76Cd
6PEjB1RhVbBrS02pymy4HnBg1wFdhCaXdDFbrIpLgbAVhRZBAYaMuUQ5EN6aNe/Fgk/fxhjqDl43
kp2TdmgCtAL6bhfcBEFZfbMr47aFlC62flu/X1EPIVqXtUHGzBtkFrpXIUd4wwIE/BsKlTzk+9Zm
UHxs3a19VPo6uXIRX1HKD7c3Yij/X5VCAJno5e1ARdzmkUPC6+fv/4r77NRlKN9pUnVTcvvofRIu
1oDQdBbwwslnQo5deAuLbkTnLEV//F6B1IDTDfTWueMjaLbMbTn+PLJGBndDPmg8U88+KUhgOS9C
Rl1paRtzXENNmkPgMB01TlM/H66n1IbCZ5hKX3je5YbiduBweGJ0Imq6AeAmQGKxfBR0o3d8FrZX
X0oOvvJB+kH2R+uXCvEMb/F+ENvW+whAD0W5lmBWPAWpUq5Ebl7w8vUxuh9dDOxGoz6DFqfx89rl
/mq1jSgTuDNAQNz12i4fzkYtamj6usdqLH/I3OBwaikz/JYoAw/wk67J6KweLBcziiq33cwLVELq
XD5vEuXbs1tJi6rFGBfq0okh8DH2sXIEhN7LBrNMv2yIzA3ATMQqDhJcora1lEpcgoapyjY0diN9
We4bNlrm1wtLoao25emlQqf9VY6AmHXkLJC48XSBZ/PM4lWouWm5m2G8nj1QceKInn3o8G6ljjFI
pAkyTeDzFtrR8uykUpL48wq1LmX9cB38mkgk4B6NHMBVLDXd/dPh2eGjfD/FA4LggSVCmQ0A3iEA
U9o0qRM1CdjQNcjCgrjSeLQYwMbqzKB5XXEzEQt8Fz4j6f+39P09iy4aRt94grx6FUj2ZQB5qY5M
+1AL8l+PhRl5XtYA7v0mEZn0kRT2huqLoHT9mmcb5wJpnmxkPvH6dialNN3c6oFumy2O141byPRa
rdahG4gNTxHR9G54jx0n5UZJf6TmPsG3W4oXQF4iuHiP7vIbjq4n3B5m7VqQeX7Q9zCjzvRr/SOB
aibz0bzHDSDVVQ4N0ejWGbP10jQA27SJ5ODXAhmilcPkS1z/5/bmGH6Ic4gtXcDG5wjauhYT8rqM
c1QS0Nvup+F+HXZZzWaUw1dkD5oSpjq/6bVhQhtZq9taOMZ3cTXGHVNP/PFI1yHfeXRZ+T6ad1Dn
+qIICYwuA+QET9jbz7r5cUOUFyt8Qllzt0y1Ex1ufGmnBhJWLJ6Ftt/RKYJzp4rWOXE8gDUdL1EA
Hf38SyO9C6c1e/pJmgIbI1nor7wVSua6ZC/9wZp51PyZjXksMeh26DVfN2L5hmVqzbQNY40YD9s7
VvO+VycpLa1+I4okFs9yxkQxj7I49n1dnllAc6JDqmGIOpfDiP5XB7rNwhtCUxEyts+O4vYsbuC9
3jHEgurXE5uZOldSpcVg0spqsbwymObA9mUikbcdJjw8Kohu+EGlv2zBOtedliKCHH6YCO+R7Dpc
F110O/GoR1iGLKIcrXyKuilOKl0ActQ8xu82YQ8KMhyYkps+G6MN7D0r8VmQj6Wa5m4TdbzLFoUX
44/NHGQS9YNdlg76fdzxkGXIB+GeJVfFY8WeKuMcfKL2FC7WZlWYlbTyHhJ3d1m38JMaqwdj1rb3
TAmrOoD0+G4XZdX+Ll56aOcW5V6UIVdhuXqJMwsCT81/t8o2V2AwxIwN2ZtXOoW32zGZPIHPbZax
4SXuzjVUFps4MD4QeNuhsIxbPzgxfa1UFobIOKB/n7wKyz4+Vm2QEn+u5IE/d7ECG56Y0iFGQ+jN
/T0EZNQdUq8YWtGRT+OGY1DySI/x2Q4QQwQ0Hp0rEwOWTkUiP/+3YUc3/Ah2uhgNZ2tYFu620YWx
l80sPS0QAPcIs7/6Qd86W50n6rHfOzKflaxmvN8yTQNA5NTLn/vJrrMINNTTGti28KLFpV37Dsnp
prDIeRbUPnEQKtdPrruPVx+nzMySOSeD1y3jflEuxxnbuVAYsFR3mHUgaZrb3LovUEIaOEI1sCet
JOVRSQJC3rg2X0KCBlCwkW5DjFxTpKUfLSej1SHyseAvGs4B2kvn7mOzBfR4BYrdLjXvfwUZaOGi
eo9USmJMtuAizVVL8aHZOwdMPKb1mFeUBtC9id2mjTwllBNWx2HvlXH/LRmoBNBxZPab1Bqv5Y9U
f7K5v0DK2uPUR0BreAwWpyXF9qCKVo7eTazknUALN8pMO2lVGxjQwwbm9Ut6DAY80DXpqh4vd536
3ZdIbPDQIArWmqwzNKNBgVUDtYXOBxWLHCrw1VYYNSirSFO8z7vffjov6u3o/pzMCsm96PzaTJE3
Rmg/tMYnQYZ/FuVsdUBZ2Q00h4Pc1hzOYWw0bwZgjP/PkkOA0kO6jVZwzhzknKBwQ2cdo2JsUeAa
vDBHE1bhTAl0ErwJn2zQ2pF78H3g/e5VwF6D7W01h9C3JN1SVfs8Orledxxxe5O/rm5mRFxY+RWZ
rnA6LWXgPiVE6Jly8bCOOy8P1j//p4gYkq4u1zK/ADGjz3QmvXB6Nrg7FERR5SsG3LxPgJjfdC+T
AulMULO5JRoWYcEOfJ5Zk4PfNpQdUMiD6+M/eun9yCqA2fTfI3bNl7NSJ9zSiHRkq9ciGXX06dqQ
Y0Cw625Wu/ZSNBnW88DbwGdmt4YuRoI+op+AQtYj+PQOANeeLlDrCrdZF9UoSL2EL1VAhN/8kkZZ
CzcSPnNqAYmAOdw41hgllTk7lfVENhTTye4/py/5uUObI0fs3Yq9puoBjIcIxtaKdQ3adDIz8ViQ
1fopBiYmCWz1AZsACc3wtVzc/XD/b6fTzWELnDL4hXgFnbWA0GrW6cOWS2n6y79oABAjdO9MJTef
58eiW3zm8FYlxCaHDDKZCtvAhmPZSzi6pzIVMpHBPrg5eTkN1Ndaa4RHotGm8pXvQM6Zd0RYuwZA
ZSm/ruYIKjVY5H5ZJDhJ/+lI+E4oQlGTJ0nREXH9sQ1EykDFANFacL1tyOWBvoeyQzvx45p+vC/E
nfiJuBP2R3wr1JxdE0+tQdEEr7BU0MU877Wy3YzEk1JdrIWpsVH9MDsqDjEzeerJeVZPelbB56QL
K2HaURnNzVZ1F3RLp+Lcb6W2bhqVW/0TLG8QUD3jo6A+rWT1rmXAoQyv10jCGVmDu8SZISDYwFyY
OYNPhgBlLwFmTrxKq1VfrxbqOShEQ2w4BZRHPyRZMRV/VhCyMGqRX0tkpeMRx/hCasqQ+wBmVaJX
IS19Rlz8XgpqqZ2ZTMcJf2HJI7YRTJHvyqr0wQmrLhjEuaY+82cLhdGYeBhpxobrIpl2BLo8CN80
FcwphrRq/Ba3NPyx3gZd9wx49nmiRIDXG454V7eLifF67KA2INarxWyF9Jh2SmPB6B7JP9cfNBHE
cBpG3UfvGpPW07ZGmwJRZbnubwbKtNeqisj1ZZToXrhCknTCgUh8OK3Z+Sf1ObqeVEfUcvm80VID
UEsG7bpSDHxqy+Vg72ALM3gazvRchZZmkxreNJ3ocNX4LSJtmxe1o86RfZwP50m1Cc25DTYQHeYf
GIUElxS5BbpzhnWG3Np7tg2yCWz4s9vBhhmd0WX01WVikzhQt/ZSgvGptM38sssNMGNNpRtVpJjh
6WLIv4pqxvcmXM6wTUNZcZ+pwbyYb306w20froS9D3AwqjagYzc0q0q09wHFkk07gxTnzIJlQ/iQ
ZYbtBkHeZAGDXikMgWpeGl/SYBw/Ia+9bB7mN30RAosvQjx+jTfTus6WT0AWrNrQz7hZdpx6Wt5w
njFBC1bbdD8SYGzMej3a7e5LK7BBQ/jsBJJP9H7B0eqFI35EEUj8HFpxvRfI05CCxqCNOnjT0LEZ
k+hHTMHAWFZQHWV5uC2nDTzqKWxR/PpTD8/DlOtj7IykvzYND7r0NV1uj+O69QBx19AVIcSFhmi1
f/PkK9juzLX1U+L+WlB01xWmjA+CfOyhO1lImxxTFq1tKj4cMCO1AKrAjTAZ56AbrNHyj4/6gf+3
vs4xxb+A2145nvkJYPpRUdyMRDYOtWHgWy8tI/3tqzsfUFBp0/pgFPE5XwjpYCW7bznSI6NokVuI
6CyO+8ULcb2NVezLeb1HFTF2rBfwdWBatmgPaUtLF+engvOZMojXnzae2Pu729FW8Ci+wvwlj/bY
ZSa6yIanL5SW8L9x5A9b80vU/JFrZe4ALvIsHnv9FyE08NXEfi6Kr6GPmix2e6vn7TrHK39bEvV2
W3iN7UJEZZtyTsI9WTz0d8TBsOMLqd56voc2x4/2SekfXe0wDhhxqsXbnREkK6Nf7/GlDppmkumr
Gg3SrNGnx+sf05nPmEYJn98sDNYDny7w702rVXjBw+hsd47id104Ixg8iUaXZNNIms7XHB8pdepm
VbrbnVUa9+Dq7oJG9wbvYUAG7juNjDUWveHMjfcQAemmMAyfE2BQt2mS/aT6pbAZnhuDTntP2V3K
lROppr5679ufMAcZuJ2uVekRiDqh7cccmC0Sn2prau9Oa1lYHh7MKiTCdHdtkTqyIgGz8berGHwx
bZZiadVIzk9zTrkA3/5M//IN6R4i6P39tHfqgOV5v9Ez7l4EPm0alKlWjHRi3xKrGsnoIevEk7wE
0T5kujgckt83MAedtG+3nat+FGj1uRX8P4t0s/snFPFJ5GisFPWN89KQVUTsBUMFWwsDtVHS7j1R
azbBTwiuXhP7YYZs1KWG09Q0T5aMRKFRkfXsuu43UKUOmVwZV6dZYqicLMiC6ONJCWlm5ydBO47p
R3ZIwxnhq8Tp1rLeBAfJ5Ta0oKv5+ZTsxIp3L9SEWmU3RDDC8SyGnqlIIo7zNZGbfU8RulIB5CS2
hS5KofIH8XC8SOvgKRlyTQ9sgBudY1bPNMd3hv8muwLNPVaLdt4I/+Gx/1G0WNwSyuZWdLpWf2Cp
nShHw+iMZH08xwiFdBshxYtGhEd0gZHzP+KID1hcrx21lxM41aIZwO03UErkHQ1JLOPSOuYOpe0+
lARVCUThg82QEnxJRatUZrBddNiVY9i8eytMw+sT6JeL0KZaKJOnCAakJSLr0Ckc0lFfV0YBC+ee
4U4M3an7zazqxhibDFXCHiEqDlgAaI7PGMHbuO4HxLpTH0fMy6ZHSIWooLLEaGM/Gs3CpaExVlov
xysSdKKIyzMHduwvKUaSa3mougRgS/ammNngFdh7m9HwcryuZj/sKcCsN+ySX5kWroKKzOa6ccpw
wh6GpX6Q251N8EAxB1B0hKKWXHKqCvnw0HZhlhJKies/shZXh/8/rR7MyNvUc9efE+4oXHzs/IkP
IAsHfZc1m8XcXjmlHp6LK6bP4l6RamcLBc50qTCVU/dhlObx8nVQ/egPFVLv/KN3hf0rWyWEvi/e
WQ+F3gZb5b0Y03lHpmvIqQZ3mkt9yMc0KLZnuxVfwpr5SrGkvBJGI3tdxJzIVh+9qPaq5dQJ29Ls
iZuQwL43gJcQMyw9sW7k/nz+k2s5bAE8W2ZXinN0mjH4fI7AJ/ZuN24x6fs/XjqW65hjGkvhT8ZF
qW0PXWWqYK4c/j8CBYmKfKwrueaC6ouSREwZs4feSzmlHUUROSqVg8SrcGczpOg29nJvy768uZAK
dHJXfeQLXdnKEqZBYejixF7vzZhqx2uZvZpSuAJ16lTYtv/K+NLqxuJfJErzghvvah/fN0CvGPoZ
+hJ6Lrcf9aXX1k0FExB3SYWYjcAWGGFpzoUvaooZWISOfTankAXNeL9xq5dnmAZRxdXIXaHjaTnq
9531WH0nT1CaPA0R9dSu5ElK3EtUDyZ6CjNakKUlvnuCQMzHnqZ6et+5Y9x53dZ+OO/3KDO+qMad
SoRxYUA1FFoTl88hEdVh7s2sG0EiZRwq+O56xNUSd1laU4amM6fb4yY5+KH1UVimYrQeQTHfq5qd
u5hwioHn7IdN2NHHQYFo3TQVBSNjaEfIk2xHtb5aLhCemP173TnPow4PzUf/ZOaAImvus55ef02L
lNW++SlCWySuajOj68BwwRxKjcistPD+KlQ863EmIVSXzL4GzZolO5ywOchtL1T+4GEMeu9I2Z1w
71shjg2KZ4KYryA41wlg6M3sBRQrg7Nyro9ObnU9AE8NBnXV7cff3RZG6rY/MMfg9MfB/+NLmCF1
JhI1y9s3WWik2E9uMcNquNkYfCHZSpkuaQkZaOBnEYwfcM9x4IwhDEY8jUTFg7rC4XmeOv71TTvs
bCQEtRTV9cpUTaf7Z26dCaKRxhu8hbPuCPHzN9B67wY541AsTAgBoJXc/BktZo2joEjknuAMbJgj
7SUFvnhUVKTENMetF0pIUsFQQUnImi5HUVvIfS03RF5nyjzL1+Kc/u3oivIqzj0AhhuLWYW1tOqi
oheaP4PCAvXWdnmtEMAHn291Ml2OP3y9W/wY+WGy5vt7mQglt9W3AQXv4N8ipEmcT7jVZO9eUlD9
INZKOClB23Vj3UG/1qdUsSHuxcaqCDhMUjYwaoDJt5JLwt6egTEPivIHRH3Z2aHpI72jfbW28kAN
Kptwo8P1LNK/TD8/4JJnH7XDcf5GgOro0bzLYf3bLbivClIGzy7f2XVtwzJr1lADlbfg4qq18ayr
ka8LBzAqdby7oBW2u6z9ouNnycazepI9uYWGxVlNBKY5z3jy5MdkobIcpX0c0vImF5BwFY6yHNLB
mammWpoLni7NGfJhS0EB8uTaWXpIkiBFeQvesMymZEUVYufLI5WdT3m+zyJ+Qh6i30Qo5HKb6hDZ
HDCbh2ugokxpp74mHuUuw7/TjSbQUk9yzisv4QVYBvEkGrD331BZBPhITwGg5iWdIZzYMMSMlIji
RiPY4zR5Nm9+xsWI2RJiNTQ6F462lywHdgR5pftQarTc0Hk4waE4MuH05oU7MEGtloOh5i7rMsRQ
Yd4JTmUBg7oY3g2mJtJe9TPfh7/md3D+aBgtZkcBNkUKvaEBX7gwFj3emjCTz3dVL4osSKDtFThl
3FiihSWjMl9mx7lgFIdwBIXNFjhLli6t4AdB+UF+3az7OG3JGVUe1UFUZYx/VlXv8uPXZZrxncK3
sXK/BQeejgHcQ/Z2/z8wz2IEejMBPfudRRR3KM7z29f2o+QxIvZTovfzjU8lS9vS1kXC6BFrWwyB
MDAgnuvqNcYZnyWgv1F5xDvslCUMjShHifRv3hRA/1A814g42mbBnSs9TM4B0snm55DAEcgS09sS
MRAUQjtAEHqbfuV2eHLROl6H8CQSIxWtBWv6uApte5JSquF6Po7tETs47sfDvi8FhjZ58q9usHwf
r//wREA+DJ5Uzgj7PUDj+FG361J+GbFQrFLREAsmkvfQrkYcyKhI00MFzu1hFwm7XRH5blUhN6u+
EUGdZHJVc2HE7zT1GuBlIF9h7iars9pYf3GBGzdsqmw5Kn2j9B+VRasYylR6EBPrSyCbnHsneWVG
QYwTH+L4c3PZnTYqCi8OOfCR9Z+KKdeV5geN8kbZ5b1P72sdXgd2GF/q4GI6tVzcCzxBiSqFA0hF
1BS1iI6N94ET7MsnaQHp+/bBnWfi7APBqg/OzU4ZEC5qHEB4JkbW0IxxdfnkJ2jbhHAuaJpIvsCw
0J0h4MklAZnb3AD+hsWzL2OuMhzGqiszfxAU9sPrNeT4SRiY7J4gXEumFLoQQ0/vlZpQuHl1Phqj
HkadrKHo/EwQXFTmF3sI+bkl1eqkC0xe0YCjYzBIFEFc9xDKzCCFoq6IoEBe3xX9ejWUH6kSYVKR
EwWDCMqyNUD3A5uUqJ6wso1z2dpzfxQxZ+EHvBLZEVagQAiVni0P4GerdDrzrUdiMNvXCURqwfh3
EiGXZiiEGXR8go1yj2/I/1+37+Hj1DL4sLY1PegbFg1oGWO1DxoCSmzzEh72qnkAbXTApQ6vYnc1
e8P1HZyb6busb7wuskfDXKiAsDlG6BCi8WwriPxnDJViTWUh9Hg29UDcZswQpAF0cEiOMtOo2/EO
vZS9CMo3EHy9hGjs7J5TIhOMiFWxYJiYXIntqUnQ+lD0xml8iR0OKjec6N999dRmuFiS9msTrz80
M+0mTpPV6jD0f3/9Iu4a+Iw+4ACgiTokXwmQK/Qvupl0J9NxBTpD5rmbSz105ZC3xp4DA5MkT2vs
1fm34Sv2LCKaUQuj301K8en8RQE2JbNeey4v68SsI0NzrA1jdqbPxJ/eruwc3Nc02/IcFByfZsog
2h4kAsTmAMETKER93duA+0EGQ4scKsbAu2HqAjP4VwjHZmDPuNRR6Jwq0YDAfUUsmmp1IUfXty4/
52x8edAx0KcT1ZVZwc6/amGFmLu1xswIwHfxuQTEVZ1fbPj76T2EtoOjd/J3rFa6pHcuJ7PEntZ3
4VhsYZL3lH+4H94TcKojdKLiuq3jeWJP2IttWOqjS1pmpu62IhNNlrNF/OTjtGGllf1HiukYVHiy
xhJdEFbEmI0KdAf6zwwhxu+EsKSk7SuJLL5UMYddf6Rv5lvSwWy77oDaKo+qxx0c9C6CEOFOwaEX
w7VNMm2eJtk3D36INA9b8/R5rHClU5JEO3WwLdLfSWn4+5rAhpmZ4ghm4IWp6X5tHukGk9438M7i
yH9VG6tEiu3MIU+YkeF/PzxlnLkoDXarzwPlJkCSSWJQHukLIABhe6oQKs5eCLS9EjwdYHyVzfLi
eVebR9w1L0ekQrMhZ11BU2ntTgPRe5LIJJvXY3yQvRSb7+43RclCt+8FvhANIX62yZ8AiaJQmwGD
Au4v+3nMMAfEozXx0Geb6L8hzpcaKfxczWTBSFHXDOpPOQOdXDTGxcYN3iY+x5a8tXKHpF1l/9pH
nhlyr4PAYOzkDthznT06Rx4UJZxI5VecCx27WAhRvV1W7YDTOTp3Rwb1MMtb+DXbQNwPW52+TjEt
fq1s9FaMQalaRugJFpg79BRaAUKsLuZ7KrHQP2vXZMrlO9FheTUX+KWGWB8rUoZkXxw0LGddcMUA
90TgZqLlxhXsT3imA8FoQaph7goGOb7QJ+uUm8KPvtNu80RdtzJa4f7QXMYVTQA/X8+Lfemn41ee
boNfGkUGVwCWh8IBqZ/GRxTxYu+QtysBNy2+WWoIx1g6aypRaVhZ6AVIYNrD4tp1Pops+0+lhV98
IRGLx5L5l3cujkdiNf51Vg6aLpKTENsr2TDJ3mMUx2a01WNJbAvzUacnE/u9p72cN7jxm8PtHZzQ
nPeQ0rUKAkudu35GK+1S5HbBmgOUUSPF+cneFuc+N+/sqSx1rkewProf6j+QwO8GHCNCVJI5Xzg/
H+sFE17hNNwf+HJnpC+e/IOk8DEo4PEINWPF23dd8fsGPuo0NbmH8bO6/vcKiv7BmR5K2B8lmJTE
yOEeI5JaEyfyj5kZO/8RGSqRS9KR2CyOXd/m33voU82VIBaxFmUgbiy3K51/wjXeBO9lXK3Kn7hZ
60DOt13oK/A1wgYhZzLcSMyTm85Kof0IPczxx7T213d5vb+zMQzOiySYMv/O7KH0a3Vg1vub6OM3
94VgF17hb+mH7QXp+SOCh5FA6HltdUiX0Et9jcNkAFx/xwj5Uv4HdtO3l+BpfFlWV20Pu4xA2LBA
reSvHlI5iR4CZ3XKrCw6It1Mnem4p+/bYOrcILutaEjmeVRiyskLbNEo7wmdZyIdb/bN3rYJNSRQ
+97lIMZ6zgFzttl/q3X2ZhbpM2GbhjSAuKal0VxfqpERoO2dxYMhlpIUpdQX9rk8fsiJt0jK87db
bbjO4eijMBT8NF8+n1MxYqlKsgcVfa4l7dMjbVsy/px1otC2GKdlejVDdX7TNaZpQWU5pEtdRo7v
/6ehOTzLLN7COvNizqpepW+0vw0UVLKisOfaD3Oep+fVcEloHYEtPgUdn3kdjxLIXV092ve6Kn7i
BinoDjMnJML/UUU7a3bbVhWx9ZSYGTKaGJfjMcIXN8+E7abPtvNFAUZ/3Np9fTANAYdh7Oi30wyg
+F16C2RCFWGVoWeA9HF3q9qPAjRUB+k3LJSOP44GkTfpO4WGReN7tw/csXW18HqG2XPqpNdVTyPj
Nu6G0sujNrp/1Yyo2Qv2xI0HzbEMpQWXwh+qKDlHvHv7Cr7BKPSiUfbiWPOKsMs9mgZKrSfUdIU9
bZqRLkD1krNIJNhdlbGPKYEzNgmq/Ttjy+2gK4jL+EJ6aFhdXgAVu/TMIu3X5kB3ucD5/OiMNqx1
WZc2v1scQqXGGCrM8KRpCbZVMlPFvlUlwaJp8ulW3C0W3D9lT+Nr6aDX6GEDkz+YIfxELp9CxQ6/
HU6NXvB6ntR5f68kUwdEmzldWjoT5An9PuXXgHC5UfCD3JhoaiNLk70SGvxiSp9hzcVl6dP/hF/u
KmIHb+66CsPt+jWtP/dPz4F1QImoVKHmoLZAXrtJRIRZBHARwl/DhpYhwYefnTpLPtCi/81ZZJm/
tRgb1ydys3cRbsjvW2Cn/mOwe1pw1w62WEywZ5quSPv0F1ogNWBnaYMeKa0i7szTfGAPI3rKltX0
9zqZuGVFww3RW5LHNU2jQOpwZDEZQAQkYalEB3W6e7djTZVz0tXlWPlbIeQcLIRuz1DPnfjsUoAo
S26WLGvuW6ayKFcWmQIV/DKlBNVx8isZUHEnxYzPs7hdSyFEam1y/kBJEwz6/XoHpSAc/DHkutBr
uTpB+f5A29bhXtiyFzQ5CsiBIohgQCczqoaQp9W+ZOo4sA44vhXRR0w2MYFtIYn0iUI6vCvX8UVz
cN2dh5gQnAiMF4LT3/ifQJlnoS3jbS319MGFmVV427GNECosEwcR4Nc/4LQCEGccavRfxGu3cYDQ
gQQ5bm8bLWHTNokNmOdoGu2mmvWPxhNxKQkHRDIqgyd9ZnLsru7VEPfTPIPn/0pTYTy1HNbY0I8K
/243AZYbU23XZ/6y6hckd27G3FAG0gmiXUFxXQmIlvaAkiVlfaL5odTHxtajuz5b1J1HAijTTbsd
4xLLegxmNFA80aUlXVghMHvhi6/FR7njVs5uFPdEEQ2BzCBOykNlvHjnItOr6r37/78N9fK0yEHR
fna+r0cIwxbpQlFhtWxGIeEC1c0ZD190LI+MpD1K/NRwjA7m6yS/YSi2z+cFYK3vXSQxx3KMeUcu
5cS/2feEotR1UoLsZDEuz69f/czy6nL43Mf/mxTdFcGjkVz6f6kCZa/+TKHg5BArm6OqAGuq+a6A
2rVhsaHM5Gsq1WmX+nfNlcZNelLwXHwRcRmpl0z2go1FMPCLcokD7u3PwsM2mgny7C+cL/C56+ip
eN50IT0JhKXJ8NpPmCMh/8GLf1RwfvNB58n4bY4ygTD/aP+BD25BDMMqYXrccH/dhm0R0r/7e08I
QXJF6iqLzys3mfSVa0OPZYpCQq/ALjGd9i1QR8D2dl0ZwITmYp4m6SdINonmRwjcdBZ2/xyyqX66
LWWbapCKYE9okmZKI/CE+9Ck82IUzLFY4oGRLZIhvE4UchwhdSr3WmK3lgwMNWJfAVNczVlEHErj
7xRspZ93O1157Ze2CsnzZRRoswytbnmavr/LNy9WXMeU1Lh4PHYnfxYqRZDIb3I3YoCgZJcetiB1
KK0Jp0S3+C5TgK3XEvYHLco5esmcdlYBGqWpAP+embiAgbZjpNN0NgQ22EwN7zNBhQcCOl/gcILv
gpuTsiCTn8rsNSFpTH79s2YJMRbOkzV4V+MGHZ/wnCmoiHVsoYhqtpWSNkJrTfzdMo2m9b6vkIH2
vas2PX1S085t1oFWcWjvSjy0VBAi04yl/SjwtMJN6L1jj7i9971Z65BChx6NevTeCfSi0dqtf5kx
0fKDI2rnPZGIz7IKvgiV+8as4NJOU2/3nGMK/J8fPQ7NGi84HGKViZ2q8JZwFxnAYTxOBxah9B8C
TRojj8dKuOrSNsCxFNTSaXR58FDgXkg1FlFRHgjtnAs7I/FR/240ZoM7Se42ONZjGSId2R/Ugo62
SDP4mQdPI0Hf19sRM4M2TH3xnkE6ToIP+/LuaMnsoio4tea4U0WRwfoCV53py4mWIUAek0uojgSD
MPjNbm9UYj0YLc+1tuC8VsZU+EEhjqOb4UZ1LXS/8gMepsXeqfrB4pApNk0aXbz1ZoJwB1vgo/Dz
nwJBkA8SFVLEAmuN+NlkrLkjWjVL507S9HvqA7v9aQjo7U1hSAud/9q2qLaZRuNF9+Xy+ilhj1Bu
Z88QeI2LWf/uPEPoU4MeCFepRfc+3si6gsN3k3mz8Zqwr+GkQlAvqFFwgwlOd/96juFaWUyLZZyk
81pj2maOxjjCL2wx1fZT8/ut+aGl/N5ZynW0dWdHTX73ZiUiVZ7wOo4IEE28jf2LwELIiPRPAMAO
I1ykm1e4SGcnSO84YhjePWwHRSr1baK2olU1EY2/PUqcAeWBK4iamCV7+Z43dzSzcky6J8VioOLm
2ve080BDMOlv5ns6Y3qZe/wHVqWLM1Jba9BlaDN2+gyZVCq91UjRU3ym5fvKnCxgi3PcrI0/6SyS
+ymeb18+L27Clovk1x/SoQnaICJdXpipM/l7glmfOm6C8tl8/RwFJykhyQk2VmacH6L/nCxX7BrY
vQZSKT80wA/WDOAnPBdWHRp2WY2fY0wHJgclBYT3ZKGFgLf/RcfQVKjTLF1VCrlxublKQU7o0spb
PNPwfyd/DVwF2a6YP1sTbfWXojhWzJW3WIx4kwabnyayc94k7sW6M3ns/GfEDbzVSUs51FRltVb5
dxP+flib7tg3bj5xRCJBC3eaiBbMyv9or5Um0FYW2Mb27Tl87tZdq2nX7t21d4cZJX7zvtLQnW3p
C/YRX8fAiCIH+tbGiHSS3zaeJkEeiKP3Dv7g7WB+OUG42fonSd2gajmSIIzSZjqc0zJwJb8YteN/
lcw0xP+Tf8P86yB//kWWitPNPD3MnLeUKqVu2jC2izHzvHggDy17GFaCJz1JS3LWvraScfCYT3KD
P992UlkAUf4iDpp7WFqfWtPDreC9W2NhPH3JxwSMN0q0WBnhzApCNRwBoKuts346D4Q9ZO6iIZiQ
dwUE50RplpnSzRrHCYMCxLPwD+9feICAjiClifdklYPPGy3q7TZzQRgzidCX9/0klmvfzarHoE2t
I9Rewk2OGI//DMa2ayhQqLppy+wJRQcWRmkGtP0gb5P1XNL0d1navSW8sp/73pF7tpo73ksGhXxW
poMAtriBxpVmk5m4rylO7zO2+l4HJIBs+tsKzWrVMZ2E6j4WrpJfzr0oJkMpXk1orEkMkZGcWdWZ
yVp37l73heP5KPqfNYIOfTPkOpWLyL9m2ERtakhkiJrqg1FuEgy0bwDsPFiEhPdcWKRrUhl9EJyB
2lOPXAdytzL5LxEyzeLFCt2hw9xIzYGs2m+0gANLY+g7hWAMB6Hu88amr2cXdguGJEiUVuDAGWz5
nZ/9SkIzJVLAGkxHRmxDz8fMx+71iyhKttKif2Od0X0fY4hyfoe9uZSaavP6RmNtTWvKIORsllEy
oudnCECBpLyJKC9Be63PM60ySf8cebMTv6iwFrLivFFcJwvN15CvSly2Q8J9pYORtNpMy1Vcfa3U
NPPHpYcsoA71qyTNzt6vkeYHzdsyM+4LZFiWuWNYwkjl57o+h1fmZ0/qFGakLLaPo61LFuHw8J7/
9CGRV42Sxyfx241oPGtir7hjIlmSJe71SVyBrrlzmN08ijH8Sy3YHcukUJUYGb2AXBJrrtGOtuUj
C1BSX30dLUeIJMg4I4y3RV9/POxzs5/IEJRPNj1obqDIrlMv5GBxpFYvwBmndboAiNDHT8gK2JkO
Hiq0BEbNzG6hCIpl9sNPnhyrwUxJqBBUpS6SYonaLfj/8PBxoikNYkMD6IlcJpnb6Ouf9G4w9Ejd
ZmLeKwz2elwqMlSxLoBD8HjHCO++zrcPLai9oEXDeHeU7u+pmlDsSvjg6mtq1rTHb38w5aArb4U/
3x0ZFVuA9Omp6IZk0W7YJYeneLXKWz5bxgcFqQ3SmKcRf7CYokdvPFoXJgXwUxAciWMH0ILBdwPx
KtFn6VStDYd2RypWb1/IJ6NwEQfZWT1H9reZ//P1DLAojOFbLxQ+FHVqW+K9F1Br4SZXE86cXi9W
//9/gqwMB2ymInfiacG8Oe8RITkiX6krm+d8ZRfsCvW8zJIZt1XMvciMw6SI9ySuUQahARSPspRi
kekZzjnlhjErGzi88inGVCXBvZ0YiZssv+L4Qyye4grVH2nYrYIujdZS9FdRbh/WtOWw8LEqoPll
E6ODHVl49Cxe7vMVHxOQOVxljGLxHwVBG0ttjPMjpxk7IPg+k840T53XP9DuTpWMcOPz/6leStfw
m0+HtIDAmBDyEiRTlqDxMX8UhX8RtlK8AEnG9p/Mm/shJxbZaHRJkP5ozUOVpAML7ERb4AGpjydB
pxlIH4A3DtEQqZgM0ODClvIY2OX96wEK4szAyk+Fr62mHWiZ1xVaulswk85jNdvfxc6s6w7n6TZl
HlvJ0Awr7TD4oz8+lzTTl5z/xYBfeHOUTBX2gG6lDjRLwTaqJSpRpddmyTCLAHDuK4aH09GV3Hlt
hFPTDhLv5JkriAPnl6TSpK12MHHSXZcb+BGO2Nz69I/JrTz1tEVO1Jwstl0TItEFa56+8RCHN8M8
o/0KIUkj7Mt56jft4lOcmyv0SRHJ4Kv3JwhmxXcHPyafjzFpV+qAlDg8LgXz/gIQdBplmrNts8FX
kCK3i31+xEg+sOEBMVJvtLTIMs2SHTrAHEa4RrBuHR/ZT3fjTb9uGdkNG/eS8qHwgwkWO16BAKZa
IUQIvFujlVADJIEm9jBqmUaU0x37c8KT20yn3y4pEWZd1bNmCFcPxEDWHxkbj3midB3VgNflUdLr
9lUc93Yfxn8saorrqydrDS8PL1JcFRbwK+xbBg8EhmBIBdJ6opk+sjeKAKYbziFiGCKE4gLD+oXi
eJKp19te7n+wYbp659o8niqoLiDlVE/5QdPRQ8UiI1ExCMJy3qdxeKKg7WvBr1mVlzXBXCiAOmgA
Q93TSMOwoXxr7YoXXUM0Tncjzrap4SLxjE1e0jawC7HF9HIa2it7IHR/8g1vWvxyazyJPVVf4mn8
toyGZoUl0mFswRSd23sTOgpZYXsvqADvzNTs/xS8ofXVfh65Vq08+lkBtDqWvzEUaIyE7Z6T6QeX
Z0hKCttPAlKH9X0QoIW09VIK4NpmMiyHJtCVaVIfmEHxijso42TVJustli0qLDiJcyWJUvS+zrtm
otO3k5jk/4oWnhT3/1WQqaQVXJwfvM1wo2MATna1Y+AvrPYymrR/SeUxygDkcAFFuLppmEJ7b2iH
xuCK8lHmoT7tJymrxi1OalnEsvfCZbeiQvAfOPhhJcSrww0RwoQRFuBLeb6PduNm8kx8Od3Xe7/C
0etpvQbwkLbqzm6eYWHEMOcwLb6OSbu9W/l/PLbmL1NI0uh+MF3fejwtvUeKve4SBpvzXC7LZhOG
jAcMUEbrEn/vu4O3m9DyjD1uEsfiPZiDLojek0yXquFhkflA869g68ubaB5Kz3q6H/U1r0DRmL6O
xUJqb6kVHgkZviWvLtSkDDVYHJqyoAPgd8ysR6USgyqE3os0+WlACED2BgAXy+ZhPSxyOf1MqN0p
OJcxUT/dp+8lBoJPXmGtdIeqVMrsegJqQdVtWKzkXDQ/jI1faKEOUYPzQTjQ+z1vCoC965skgdmk
TAEkusFQ8WJ8d55xbyQVg0DwBgCM7ZT9XYmWwGCMQv44wCVIuwe/KhWndcZQf7WEN47jmT7YSNQ1
PaxzJswpHWlY8UFmURteuKIN2UnZ0MUOVfjgyVb9ynl03VbZXEInrRj87t5XG59jMDiY5kbW/2lO
LoKoPPjtSUvLPghdkz8o5A4bEACCWNdC2DuhcH/hNFvEKJr4878VkRorBoeqj6XXLMTUz6jxEAb5
laUX/cvO4DXZsyrr7ti1ZSop+y3WQRMQgnY0JGvL8tHZCVWC5YSwes0Ta5ndZ0wcKcyURftdaZoW
n+od4+1wauW/sGeE+43Rtmoi5/k7xVTVMei0H12fN6VCS8jF9BhBRUfrQHzQZaTzXCA7DGmr12kz
Y3OI0DWjkafFcJDm59XvMEe7dvr6YwlLT1iErLoPbE2USnn7TrmIJBBOl6Izmt8IiP8FFuHHA2Kb
QH+2UtqRSz653S0/mZ1mT0oRaZ27ZrYv3BWD3ZlUlkCBm6PCVonn4kD071nJIw3d3WLwrmmbazVi
SMQeRvSDLewcO68MOaVJGYk5b5fDxQs4geMx2+eE9tIHv1H8Hp1yq1KWNmHtNez6OgdmsWtScFzY
4GgjzZNpUCm8eASn1CJ0VUp4Kkb3FG+5USdKGcbZhA7LLwlnK+C/u5fPUNVAJ2K1BnmuTTW1H2YF
oEWC6REk5JQ52jYrRw0CChwbZNm3HqlCMuCCxYykg5BP9Kk9s+wXoqMgTxRmsmszjfoNOrTsZHyr
bI3p9y5b55ymGIp9yp1h08l6VDZ4gZy8zoMCzvkLwpGE495xea24BW6PERT3i1pJTQwfZJ57KFj2
pQsTqG84SNd449juk4ZcnzbXxTBrBrltzRWncgtiWw/A8a/FdLHLacGDlJCimSGOc/XILoz/CeUg
1fQBbZyNytqaXUuvFzBtOq9u/+G+MTEdYAr5YPHhwjINHJAVZFmL1stqJDx1yI+jEzMHzTxJDoX/
uYIFlyD1MNPQgbjnp04F3HI19lsDG8kcuGN6UxfKVOI31f3Ip0jKXh/HmH52jTQTIo80oI8qR69g
cBCM6m8Po+c7LQx1Qf77V5t/AxwJndo5IggHTNtI/FCHzYZAcSqSPZl8SOuxCMVlajmShNXZED9j
4PU8Xu11TiC9jjlg2L7rczXrSGk2Sku9CXnaYF619S0d49SDc8162Ao4I088lIVh7Y+Avp5dDDIG
/8K14E92ieX0zZcBHWas2xNdqbF6AyEx8JO/ZZzUcd2gqXPwiZwy+4V7znX8TMrbwq15QZ2I7yy+
73+Nu4REaFGpHusdZROvhRnktYm99as1zuHgE6M/wpT6R+nOcbGa3dP+iEuX/Ko5jx4X6otnUB9v
n4tpY1ND+InQ6Hhp1BN3DOCpt3hR31DpErqsmWZZxhuIe0B4xkFRDx28qLCk1/y9fAjPpPv0gWSK
ae+gXZKkwsR+963Wh61M0D2bf5Jgmm4sXOCQ1QTCzVEQ5yBoqQz6dhLuBzQY0mlTHFAFHzVgAGkW
dNeCg76e1H7Ylf8j/KjO3rkl1s94mQEZe2SAdetW2l/5dFeleBjdEKKR1HJm1s3cYTQsxo4t/IwS
Wt0ZYjsl9O5BXooTQtzm0OJ4Wodfou9MP/pG81UDDl/XdGssd8htFvuiMidv08P9q3jtztWVF/NQ
9SanZ98ga9hNR9+jxJt6i1KxhFNS/7bh7mBhi8CygVXRvg4lkoHIrbLVXOGrMvOSIMrWxzn0omcS
w84BeuBNzeLYyDrimNxE/gDsMHysgXlHqCn7TEJ1L+bfBUXoLVW2kYci7qqh0lvD/L0NLassNe7v
BVaeDShJZir3ERrIOqja/X+VTT9OBuEIBGZOObJWQ4/d705WECBVGocob9Qhu4JoFGk7Amzr/OzF
BwXjcKhrCHyZDnmbalyd0ioe22NJOmpZHZMcss6JRTscHLQqYrC+MCz42Mb6rcTB6da8GGNE/W4a
xoG8HqZCSxnyAlWsnL6IYwnChWjlbj3zB1zeet2JFTUxM+dwewznj2ofK9dLujmFRjHdo5QCgrdU
TBd7aLMC4QjfV857K2TAmyXxn3SE59UwFf2WPI/zjYXYZLWUrDw7v0BCKjIseP0SorvXfxYVGnvK
DpRDt2U5FdKgCOKlLsiIswxZvrQEUbdfozVt2s1dxTLDnev325IjBAs+HApYHj8schezp/kD3u5l
k9nzbGPp1Z8nL7cDMEnsGeGV+AMxLIRvTT1jBRwLBG++4bCUoF5ywhfTgCErNNfiFFOGs1T9+GBK
C8GES1iK2NxwViaABaRJ8NNf25ehpCmuXImP79GPN+uH/pxBDwNG/XowB6txi/4yDNpjsjilsxav
50luhJul+vRL6bWzHx+ftenMo0FkYELVVTALSsRp7CDEVamkp6EQndWyIT425RTu5xCfiCubzL3s
PFF0qRmcqoYxWZWybuxhhfj2PX2QLHooyJhSvH9pktf3fYADUBKlRbEucjV0yo00fV6onklA95aU
eAX/zkapGift6+/XckuQKU5TBQhsnIiQEEMklWvo4JW4scCcr882yFM8mxPVWnYIPxLGcii1J56C
0ZW1kiizASshBUkkNH01XGnY1r3+hW76vpKQLbKy2+J/NOw/ZOS/6ZzWLTcsOA3MfiAUQrNuWWoH
wzmTsfokMHX7uA4AYd+UYmsBwoYhfT7CnOP7YCHrSDdHFgnPoHfqtvRUN9Q96ovM0muGeVxsQEjd
6olS1p83cEry7XX2UcyhAKhZSrH9b54NYops9hy85KmWx1xFfYrH1sCB+bhGV2zFBc4AcyPGU8Q5
u58X+jkcI9HGB/tGgyskxbtP0eObfQ0fmbHnnLRmFoU93KelaU9VJgKltWCogEHBhnqi0U8T+I4/
Vhdf/kSwlfg790eeK4S8bcbratFDEhfV9ySDDtgdt4JC1a8YF33RcDPaLbpH8U4PWS0Z7MEU9HIJ
+PHj4ReFmhSO/791te2SPhdPXtMUn+l2wVvEZOn4RjVJHQs5eY4dvH/TpjTMqyOMtYx9+p7/rQky
wglNyxuIoaCglIPlGbxf5c8XT1Wh6vsYA7Kix+Nb8ypCYGjap5/gkKH3ZizcKm6lZvabJedTDO/j
PruHHtGhzOOT49/iq9EHxUVbeYMELAJ0S8EOhSfe8Nohg/iF3wT9MnloaLIdlf7fUhkiV6xXSzO1
z5G2OMyUTtIIJodiDmOYBbaD64OcOQGDxATD2GYYYkOTPvpfMcrQjiT5Rid6OHXq/KqtQAkfLD8d
6SGMIwgv2+k2FQysXzJ6MMNP7/B3LHSYHTlhb8EWSkVQqkcCRTa5vRvCjbBpl/A8i3Lvd2cGK3KG
TigCPzSFve5CYTaLRWECe6erOma7ftSH2nSjNolA4J6XsiHKrBqNI8HvIrN5yTaD+4jG3CfPQLg3
FpfHrHUgBZrmK+vKuEyMXiCHqb+hzpjd+6wSgWn4vUD8OBkSweEaTTdB+uk5WKsG2LzuaYLboeGe
AqzqnkR/OSx60qDqVDOFhu71SGF+Pbs5fkp+sgkizDutuMUvto3qWcDsBHRdwmjFti8Z4iXnnt6w
VUSkUJMUeNlxe5xCt13PfJRQqwq6kxqFvtWN/ambD0FTscEjyDUVxhUzjjt7wLrh/vKAQCjYOT88
s233Ly1XRvVSDjB4gkLWpqDfDglt9jWjfWbOMEX+OtcfOXwyQA8a5zT6d+urP3e263T2GGNpZzkV
QpvtElt2ChDhdf6bno7R29LjncwjfQ9zhm9X/TXnBtGA7jbYLML/SsQWecqwWORjlpIKxwXAh4aj
l4WsZonOOIuLAk6CSm3+TCrb4inVNJH+eFwAfFMxgMCv3mOSWP1QX9kj2ADMJQjpTGR+Fl2I2blI
qDSV2w4YYE24s8PnZTKEzXWTXBijk78F2yrW49PHIg0IlO78Nx9DF6cF9AvjlZt+GGgTKhdxfgH6
9ph7KymMcA+R/ZLswXdXQFNRiM9n+sERoP/rXi6W+FtJUArmfQ6j3OFgShRK5kojwp24zgY6NmGW
vWYi4YjEhd9eN3XBmIHGSseRCmfd1VECrJk68mo3CDJSN8ybnWE1QBm3ND502B2UfKrDfy7qDOfZ
i2bGZHlH3YJaMv5aMUmaEJnzawSKQ2LQ3UpdZLLJ1MXaRtkSu/A14h1EKH9ONbFfcpg2GY+W0g/U
Y1aEmZ8WiXESk3hBYXe8Qy6pbPy7zi7zd+7aGNCEC2NbdO0w8uXQZKN3qKoc9bOlsmd+DcLKSNbQ
TluLakEHBd3IEVjaG0rYbP4KeqIM8i2fUtkmhrWk0G4OWOFWjIt7ff3mKd9oHG0jSaa+0fiRxYZz
K2DjPfVmrEoaKJvXogiv2V+mhb9j0WZnS/2j5bF7wrS5Pjot/8Ygp9JMxc+OG5MY7KB55oDKAWJg
HjHVAzBxfVEEeJMYE0IGCepbcnepL+K8oIo/+BxuXEXX2Pc9pqN7yQTiWrBjJMXEWsH9iVkVn+UL
WxhapWiPk4zxdldaJKCmXkKp5IZFWk/lXCZRWCG2H7mPy+Yp0EHwW1Nwbtc6tmGcXA6lexi0h49v
efgfQ7uVkT5hMvQOpBGv2akuYD7dH2SWk5jjSNq6s+hw1rwHIesv2B8O2DowTZgI5yU2DZWKfBja
0TqRi5NAtBMbbisd6sDR1xexJWZEnyrsfJCsNdhbNo1I4foHAmqmucCalvB7IszBEi5fUBk3tOqY
UGypmOd19fxMakY4/CsfIiePt7SEgrCV0jGRmj9vMSGeNuJGdFJaP1Ii/0WSFzoVmwtmVLTM0j/3
p5DQfm0kE5D4HeC+zCLvSWOTlYXf2CyxZNb3xmLEttYFx4ZWmvRMznGqIp8vw589sSRdVDb3dz+G
JXe8YuMorLBNupO1MIOhRNdJ4zKYdVLPvOJONX6Xzz/A7Fe8RXke90UUisoqyq9zTdzfISi4mI9l
z4w8gQwc4eS0zBmT6orS2kFY3uagA0vZZE7uQh7IcDYpFhs7kRtdrXxnrv336lvO8qESIYnS3EWz
IcweQyYrP4RGcZQlDOuKF/CSU5GoufyMtJxwnXv+P7Gdfme83qsJyjzQvfFvq1AN7OdrzdW0xzzw
kpwIyDdmTX0A8mWwhdeXarHBWidA7GcD/dyk3uqozp+GmG/uH0mdDR8RKLuwhhtLaMn9KsppKn1M
/U8ie8vjEOuWf6ciAKqvnkUxwzb6YSPZQMR/WB48quaX/WCy61iLKTf1qJAtCDd6WwHbgBYA7Yuw
en9060U7JY22eA1WzspcQdSH9dvkS1DvqJpW8GwANtwHiHaRXr4jykQ4HKIbQJK2fIJKM3Ar1SDf
BYvR2nii5pQlyh0LrHZs2kA/pv6/jIIHvLAh3Zi7OIkgdffojQOyWvkwgRthB7qbN1S0Iuqh5QGK
imTGqnf/7J2K+gMfAykYYEwVrxM15XgTVHpUVSzo1fUV7V7ZA6R5L3MH0md0FXVIjuIqbxczjLfO
rcdyXPIP4wuavl4mpasYB02O1z+HouKpMpBWFI5fx5DFCUqKEqToxhglnE7VG0wlLpOjJttVkNo4
L14m5I1AL4x6OPZ+vL9KHLYkYyfamVHYKOT4gw2kk1ib/8R9FtidWT4zDP5lHepOM+Wnaw2VkWDJ
gfE0dO+EprXc39qRH7mvNCyDN+B/guPV/MrjuToL3e0oK84ekvnqkQCn/28xFXMXUB9cuou+2pTN
eA53fQXefcc3XW8MlNNVm2rSfZauA4lWTfBVXedBS3RKNz4fDu0kBWhN3fUocKcXKfpoKOb3vcP9
U1HrnO00WVJDxHe7leDTLjeu0EsH2YWsfeg7y4DnaBgDcfZtBjZTTrftDlSfi2dNxXceDQ1jdvit
C8WudIjAhNzClNnqJuv5QcbIwewPHH+j9gx1kDslltMHFpupNA+X2Uy/vQcXG2/VNnI+gMdjMcWa
CIPaNtoRUvC7L4DqcNSc0pARed7Ur2ftmKo2Y2QjvjXGo1Bs/BrwjAgA3jG0EFm3HulFMixh3bTo
jUpxviF+d0n00oqZT8dXocu02rAcUftN//RW2EJwk8iXSaSrR+7YoSevEPfimfdhhvv+RQH2ItQP
JXi6PiA9SM8RYCfIpEBIsdGqxNYZnUkaZM4Gv27LDX8Sq/X/4HxaI04KGz5t+rhQzrZC4UdDz1bQ
AIJBnCOk66GkdaVfiuG8mVwx1R0jR7i0bDbZE5HBlaRPZeOONO2jmsZ4kK0+dHF9oQV1jJ7B+/Fr
/0lt/F9xmPu95yJIq//16/xDytBUuRnAIIxn9k36ZuVPpxhH6Nkkpmm+92lLijjnmc5Me49AG9TY
wp8nCdS/BxKj/MdOmgzxOI3K2uo3yw60CPHcpd93tvrmHPFVHkLKJqru7l2e23UCmqrygcPT/Jgj
4FTFh3oVuI4Ght41Js7ursI/UmfgzplaqzSYv13AGLYP3N+OBHGsvsnhTiQbX53PAJSPPBJ+nP3D
2ZvOBc5QLsPR02iwEDUj22Q0uT0PrPdImpBQN37FDT3YMrWGsFzzN9ZqFBuSoCS6Zy8JUzQ+qUdO
fhpkbP9Z5mPwr/hmiEsX2maps3dr3dTwPWjQBrQWwRbWdge3w2pWr0wQ5dIoqwn44sp3t0b3jIwy
K2rHUi2Zmk6hWmOs9HEEMbyb3kr+4yXBY5swkYy2GDKY4kFaxdAq7oXxmaQSXfyRhHzCNQvaSiI0
wEPvlWp5zh7Ij8oJ8G2YN8s1NEGdcmBbKxvKWIeLUvlui1PrX8orhcnZC+8OQ0VUTS7Nya4Mu6l/
LB/xZ9IYw96QzLcAOGiZDtu/hr6WgxWmG8N5YAzjDK5K9v/UYKPWWcfkm4xJQDJiScJ00kGP0JZ9
sxNvVuz6y8Udqlg1GHfnKAJwi2YxZfwHA7X8bF9ff//vI0RnEp1M+a4/f+A8PRIUEC20JVxtBIU9
ggTBTxgeb24g0qjVDUu3pg8X9oHDFhZwc3CXXDfnQQ0btK/4yv0bzrUi71zrndbbP0VPgRXzPBtc
sPQhq0x5yFxYbECkSNFLr3sbD2TyzGf+eK4dgiExqqAMdyGRlqMjyuNzm0d2+DlYt6dmzsJZweWO
QqRTfZP86EEiYEwqDGlEldPrbFD5LVef4FC5RikQyFy6wVcZQuKdCQ36+S0JLYTxsTa8zOC/qHAw
FiA7H4djAvXAEhbV850vzXGkwx/Ye/t4gQkevQGateHnajdLV0vRqx2KSrCzqWH0KoPCMmbCHJhk
hZTU1kWuggpX5VUXBSCMs1fFT1vCEPOBp4RbUkdLWWH2cpLAE2FNLsYY/3e3kiB0rJGDfqmT5HBL
YQ2Rlke+uAXRxpJBKBNJq9+usoCLLU0ZY2skl2/Qpwdh99187IuW130tOwjaTGW45F9+BrJ0EQTo
wfKV3yVNdA86ruDC5IFV9WNaQAybb2H1Wipd01sF/iCGqCPAwsNYaxcvrpYv+zeB8CNSMaY8/1pd
ODBtP863SXX7+wCMkwcJJnh9CRMxinx0PGcs1oa/6I6+42bWVQ5Yx1fZ1kUGcHXxOU9p/MOVxxcP
1VWdIZE3j94s3NmsEGP5CIFXupwCYniD3SLA7prb/XVB+lzhJ04/4g/CVqWoCHvrH5SG/6BVB+z1
pDlRiRXx80quiAdSm7cuaYtEdfBzt7xMvJEKQd90IBxIDGjRNAH259il59nm4qhQ8yUOC/nYg35B
DJdOZurOzDk0kVXzdfjuufCHjfQx4u8DbaI1J6irUEk6PrZyRWm6KyzGzT+/YVpgHfRiIwdou2sD
28CDHfMA3uSCPVyia7Vs0of3ydblGgkRFXFwthn7CrlCdfvnq6LhOuOONNeK/lQWbiA/89YOP6DN
6YlzCQa/wdcwrV+AkfvRgYQpBoURwxs4AD0te1LBWsRd2+Tst+uF6VGuV19wjGb49KUvkTZdc/fi
wB2Rr4l0DV1MYZnSP1pCdNUJZB7w74Ury6nhjhUkV+izcMUSeER+DCh72ZPPF5v9ZfbJJdHt50UF
HPVewfGvBQ9siogkKe28ymu+zD5Os3KRxYww1XUkXHmqYpV7FLxBpSwK/bFYydAyJYjK08dUUU9F
eAexCq9I+UOs7DnBYzK7cx4DaMZDwDzQ7t30Vu/HQ3ifeC+9w5J/rxuUxtt4Zhhciyu7a8xYMejl
peBaFGYif+T3Je3oYVpJ6HRWta9PleZJXHVMHN6KqYO1T4QPoxsoKdZJHlIadfLTI3Fv0aR8i0+6
+NKzI1ZXLuiEaICk2ICX3C0t94MokIIK0Ye1Qy/PuKoRCgJoMTiRTcfTr/Ao2JTLSplM6+Kj/9Y7
N9uQHJoTXKvTh3/DNhFletg3YRz3RW47dOdjzeoPBALwPck71gUYuMHTNgqOfynqF/ixsNGQeKFS
6sL02pI6b0XVa1/75CQ2gpa3LgXgVWr/ud5YabL9zhaL7TgJ4VZxilAm+LSuXIoDwE03Ibxd+XGm
AJ2NoG3Ar2qrIwzyN0R2EPzF+wDNz8fQ6Mk4Mka5JCEna/F97re9ykKAi5FaEVhIB0C3Z615S+h5
2DMvYWts2vyyQ72O/eMVjhBIPoP0ixbrKcQMDxRp4QTdE/gicyMjnVrUvu+e1lc/Kj2B0R/yzeW9
ItHccn89Q9YETm1YDUEpZT7I8/vS+dEJCmdkbRBYQOZZI2AC034mlRC6lOUURJe7g4DW69xxyrR7
2NuoArNDRk9O0XLZDgLPzdaXFUENpaZ/h4w+h5/3e87bW76gGSC1v3qHj/bZ9TWJ869VBN+rGvPM
shLbrzm8386Vxzj3+1BZpI0ZjGlYwxkC2kT+Y+D5VLag5uec7txEHfRZ/qppOc3VKiGM2v7/dS1A
na4WEBgGU0VeqYTXdJyX0DK9NW0mD9g/c8qo23lViCc6aBlwMH0fIeQvTQVUVLrq+0PA3l9pPVOs
PjyUyD7ny042PSMFCAiKGhhjPf+KajhlaLS/gePZJPg8EKcjiJDgz6ZIfNId2jLpcPzNhn1jZs8U
I+Hhp4oekLLn3t0XKzBE1ztk2Lam6PGyCDkBD7lXE636muzGB3UUOAhV8FGJP6RnyqHbU34EsRr3
fL3by81uFdFXlZJGDD+SvIosYAf3Ur7cfjoVDZu6gdGFG7PbvcZOsuoYID0xql1emt7jN2avbZPh
E1Qjc6A7YPDjqRYKB5uvfqys1qsicTldhGsA/l1v7kCfT6p0jTFQQKiVJNjXd56y5JuQWOmSeHMi
KDDI9ASslOhcMbXhkCgb786pJlaC+84ju4nf8eEKIzSC8jgdujhPYnaAhsYAGTiSTcFXEoeaLiNc
DFUWpEnjuJM0HoV+xJnexUr3dmXiE9eHaCQEz9hwt5KMFpQfcqP2tZx1z5eLz+U8JO3pcyk8pMfr
o9zm9GsT0QoR1CzNEYsZGkSTbrRTJeoxw/lFmOcd4S2zyYTFVxFB8Onv/27zFAV5IpEU2Tv0dGI5
uiFXeO+NSTdSnfulD7pNhCH9myWn6TVXVrvz1bk95ZtcpHHsHbEotlSN58VHeF+s7sWivCEUEbUG
4AixIfKre+f5n+rMlR5KiVMZJzTK5pk9Zz7zmExijgiZ4vKTBw+zos4pR93acJG0CnFPfcrXoyqd
HEUA3+vp9f5VEgglIq8jZMUbOBbGzBEpb71WO/hclz7Nqs3av1CX3i1rOE4At8BECjB0L244StZ9
aYiMyEjr6bFWWfD31jvDHQfNfYvO9djxvdv4kDMufgB86aL2LuEX7fogIdtDQk84a+7XCA/PsL0U
3uyQGfEIgPGuM8ertpiwfeCyoSRSQsdZYwjvyr66vAyUokV9e9p1oIq3HmvAS/CUj+JXico7ni8u
/kAfWQBVoFUpXDBvwxS/urEDCln4lGEbXq8lm6OJwUXfFQ4y5rSb/ahhl/6xq6HtqEkQFDnP3or7
vkvmABIUq93ckYcqkszuNVTqJ9WbxN507BHNJQVh8l4aENOReYr3Rofxl5MhYUCMVXSmzPN52ZQI
zK8zFUfKB1nG1v9aKdPQpSlP3QV50TFjxBPCa37Dro3/LTPKhTUylc128s+LutSyL/QzwW7gT4W0
vJZR9bMPh7+ZB7jLS/Wpk9sT7PArnoKdY1IW+PqQGm38GDl/AfFVCxngGW1OUPuHNZhJGO5DjCwX
lhy0X+PxfJs+EVvuhnAsrx2cLEIz7VMNl+D/jh6NWJfWMthFjrYZfxsTyIvlnYdPRa2zzsDW4d8g
3pJU8+Ta1Ahy+dpRDGR5396oGMWkC4cYq5P2r12zXU1UthPB0u5bvEL+vxPh3DAuyBuH3ybkGYwU
2+6NthmNwqq3yZVOXMHq/gEXbiV7O1aKU1CYgH3K09MtYt3IQHCDlTncnl2LzGBMMvkBHeCDPwaL
/ApCSIxRl4vjcvBgpuWAaJJ/TakIO5+qlYO+3zRKZJ6qwHvV3yvW6th9eWqblMoVkCX3bpSEtADH
6d672PeMRbfx2h2xVTgj3opcjAr4HrjRmkhJZOHlV8nn4d35YiHoTYwWTE2EvdZEZuO7O8Zj3sfx
wZ7C1KrLSCzlt7JZhNOPn8e8LXbiPIFw6LTqhinYT2Ye+boRDTC2OUEgfJ9s5hmykwab+sgtHu/0
lZ50O2zuaUJKBnVGq+aBdF8OB/A9r/ZeYRxFM1Z3pxdeoAkzXtn0BtUBNcIxgaohZxNuMhjuijhJ
L7ioHDpKGGWNAxOHjfv+iAhbw5b5jSbo3G4EnJKmTShqEMvEIi3iouu0HVsY/gIpkJe4zOdqVBji
B+qLXZy022ZLH1PJpxDtCMWSwyv3KI0FYxUv9mNCdtdK0NvpWntPumBdEqLYoVCubX26BSZMXnkF
vjSLOF7cfdN0e1iWl++USp8GeMSX/gFs19hf7ovCJQ8y3IO2M6r5plMe5WvYjrm8WQMPz8D9jyfT
mYPCvBGfkLbZHsiyxjHsYQztmiwkaX3XPjGKoMNd27P3yZ6tn7oiK2ySgeu7Zpr+Rk/m5MEa5YFk
moHrX1a2Ucb78baz84qwkpQ90aV2AWS+v0YEveGAjXnNsbMtBf3z6dBvwbGI5fK2LXbBzFmRBSw5
hCyulHoFV8KjqOAcI/Beorf51k353yJPr5qeWiDld8JRzr9VPi1oytpL4loKv1BhN3lUW/iTfdBF
zKm2OVHl4PwY69WzbxaIBopxrLV5RxIu3TYTkuMse/LBUjTCL90axgLThq2QXHkepxbZzj2Bu8Z4
5dPZFbPCYKve9P5XGeye82fuoYz2glZwVAQ0tbFGPN6MpfViaVe/Wpn4YKIfOOtnY/phjpLLpdcZ
esEvonuXMhBW1s/HqVrh4KnPBLdSXPkpEg4WoIeNIWSwQskWagZbGaurRZfBM+yReRJxq0njujTl
rluHE9VDKS1Tlok38vSf8TWCMJvmn+gXhZYlmdpY+Vj3SMW32U8y9GcRlWdi5R0Ei8usncj/H2P5
9Oj0cA73U7PujklSLluyWy6QpMCRMQN2mV0jTMQZsrB9DN3AjBMkP6oDhsbymxaczHJIGXqsjkDd
x/lCJIZNguJg2Sh22yaFd4iaJslUkKo5viZclXBBxJSarcxSZMGyXM7/H/wpTTE842Q9pqG1F/r9
oBFLKGYpp01XiVGDSkgzmnpqu4vB1fgMWwpRghqdTpvqit2AU3/qE2Moxyrgc/cL8SPvebD4VbsZ
Cn505cqOfGNI2QiNONFwJw0iDoHOAzDKRwMgQVtIaJyUMC2k8SSICRATrws9NRlydHxsGd3QD7KD
XYXI2ZW52mAi7yT6tMHC4hRhjjepcIRGIKUMvGnFipFR+x5WgcqKz7Jj6oreuTuNWmY4Jfwm0ws4
Bpos8gIDcuExtuuqkFK/jskhsyks4vhtd4S2Ea0/yWo+6dBe2lqDT7Ry8g8Nc/BnC/P0oe+PCkBA
bJLSMjIlSdKY+s0H4hS8XCl0/LSSobgvTT9rlJ8OVHXBoNujp854XtrUSMsVXC/ZQk3r8dKNy7LK
cI4/sislAhm06TBXFympVqjjXwbMd9EfAvDOnta7gmOudHs92dCZsNHP3chwrTKNSKPIsQxf/utC
Z3M6f7fRa5047JxsZtxWIKUXltpHTO/hYVX6oJVhU+NB9KxasMuWxmVvkqszM8C/FDWBemPtJj31
Yz2J9EM2+IU6IvdOvn2smDg2o1Pk3GxACFap/oxNFJEGuaZQ9ssMg2bs5fk9Wt2oLZRG9jH0STBF
BFKgAUlGGJftzPlvYeuePQq8MtqpVr8D6QeQQDmp6iNkiXL5f5GXAq44qP1RdcUplieKiXPFiqAF
Lr56vxresolFLfddIEAjpwsPX/VJ9NsiVZY/lDo4k587JWXKxf4DBUe1paJBa/3NCA1yCWw/XsNH
shKVu6R6m9B37YlJSUpize7dPxZuerthSfa3CVEAtsfbACEbcgUU4ZOHk4R3kM8iMdDOUd65gtU2
Q7+JbQPgTObDME0VTqaaQtyMUgxucJSuygJcrgdr4+D2bmNgtj+vDERsUEVdu1AP3xwkh4JkAufN
6K5JglCyzWyaZPjHHhkTIVvxRO+7ujYUGj+zBFMvNoMpg92dSfUwfFoxaNk90MpcFouYewD6ER29
jYiMRIjvS2nWXKlqtD7PyF6jRGY95XNw4ArIqxAOFoqbJ0lN9laXKgkcFuG6a5+HJgUr4wbyF5fg
p8L4yyvMwXgKCIAVQ0MM1WJSY0ckUogVVfrb5a/Eb2cGenl6oVTXbYmiYuIdhciCbbLp4KeSmHAT
vdtUVY3+sRM+KKiLrwbRHExXJm+tSX8ezB8i5iYjLHmx1oldoEBd9rViXQwBjMhdTRJQesNXotz3
CztCf0j68SReNdWn4xqfazu6uHDWoQviWmMR9h5PMszWbyRE7Of08IC8BGi8lVuPV9scighkqYLc
9wKxLWxVBU32PCv+xWsou9Ti8IJMC+wq55sqesRhnu+cO9J1zPJMoBvsV3qCYnTEHohY23vFImKQ
NwCY7Qoe54tGajdwCfMMz/CWtNH/OjZerHSTJOg+g2rnairZrzgutcBhBvPqYQVaxJU2Zmu2XaG8
UmlohwW/dV+95cPtPrUESp0vpnD8uJZmrVFDv9mad8YPxW+ZruIo1NvAAXopw6rjbEC5ecb97oTI
UTSqQgVj/bhMq4xbiIqGxp8tw2SlUbJkL11ES7RSoVHjN+u7YJ7lsECMR9CzH7LsSjhOG2JKsCdQ
GK1VqIP+BWQ+V8VZ5SMoFJvPQS4wWcZDgo+igUR9GKp2/wEsKoD4qsrh21HeJTqCyGwPv+DA5bRI
+x+NlHXuodUBrNVxnKf4cHlQWTT9FaYc+GfC6c80ZtUOKDTu7Pf8mtyKCxMUkOSmRE8cjMWhCIw9
LaYRaqbKdkdOaWweisxj9D8fcns7Sze0lPDlPFEYPW9u/11glUzI1An97Yd93prPf+IZf9O4Sa2x
6h30M9cN33ClUDvDunDbuxaWLlVQVSYXUNKezH7YsSLvWXed8g4FnqTKBdVEy9KM/uhyjF3o0ZD3
BPVLMW0EsMuJXCy/M4Q2ip0BPrDeRf44fOSwMkvfRsDrh+Re2Sw7A4F7sXY60dBDWi5uF0ZdETHI
b1wJDoJUM1t8H4F650CO0WLuMd7B1HIw4mJh1tCin+0P9RX4yUFaOUV3bggvlzX5uJWAdTYUxIFy
Q4qwYtURatX5tImCEQzvAvkZbWwvs+BcnRowDuvphEYYTzqVO398W+TNfafNg3+nl1zV5RL7qUa7
+BwhhdxW/2rkGEnGhEtHMqJLcPSjTLWuHiJmnS/rMNUN0YGa6pPab+8Pf8H6/UkEdpcwwpQAaPF3
iZK/2Nv5pjqfQ7Hi1VrFxN0TfEWlKqUcGQjRDab89nXkcCZorIufskkHyzP6ziuBo6NyrlIaKHq7
ZgfnWZeXzxsSya9XG8s9zM7/d8WL1T9PCoWAn267k/b/NK+AR37AMfy37svl6mTQX0v4CTlbb7r3
ztr/elNp+ke0LXnCgnS7Rv60hf2LaaoptushkPAEDK8FXWbgSBCPfaDBPRtRyJET2fOThNwR+qa4
Dp2QBgRs8VpRB/h+Yn4yuOi/cZE8rvkGj5ejaxvjzN6uRO8Y9fPp1iFx67wVSSDkjQNfxnAxjaXq
TaYtcxKIEHA8eL23HvSlPlSv/CeWLvKcskklCRrIWS2clngk3ATZqzCwixsTkXgGJfogCRxoopvr
TKjW5YuL0ME2v/Z8ekRMyPDF65PMXwoZch2ufFVAr9escr/gx/IssZdKqrz326DVABX9u1VVqLmb
8HbB9fhcqpQXzYNLXmOc/ehal75PgZ7EA5bo2Jfss6X4PimH6/CpeSI6WcC8m7JxEAxt85oaxamO
BKyPQL2OLc3AzO1lHPncxXeFao2VHAAfrsk1FHqSuO1ak1aAGtXBcUQ3h5RfsO4sj60mlQ4pwT9r
C0S1OvseThU4bvFbF8yVQuKMwLPHugq+2uhVJtuHs+hvKysNIzm/S4pEiM+la6JKQcT9CY7SNQs+
olWMmczQuequBxrKgvQZijEckBNzXhEeH5aGNxnmSClVZXdIKl6wwQo+mS9S6YJ8ogp+H33p5yT9
7RNJKScgWLPJduIhRHKN+PrWt8fuc9xheaXFOAZaF8Npl71+7/4xvp3eOVmHEYu0cOciWnNrMCQf
IR4WaHWVPjMwRlI8/2z+i/x0UaCXxsPDVSxdbW/MviMiZqIGbhkGtpTxQ2/v94zy2baqiIZNNnE8
V1DtmC6hrEoXthPghLZkzq6YyaEPSHM4rNnDTGha1Sse3aOKRfzSqmWog2qUK3kYnz8cbPSMMhey
C7jPvwDsrN4TrmeozFiz4DtfFEl3Ohq8K8OUkcy/9IG8QbrDwoI0OEq+DFqZ2phuOA1A0euu4AE6
jpG7MUtnZS/DSXwiwxEMET+ostuCWvTFNpmHv0S802I3z1W8/3YZvXoStI7bb1LDHgT7xSMriSgz
7S42N6IRHvcr22LJedA+Vm+RKPt7wjlnliMYQFCnD6gBS5QvP/GE3Z6o96c9jp7CIAz8m+mVxoRt
YcA20xJGI0W/jNplf0tGqWKh858eAOk+U+Ngo9bZcFTmUQ6N3ABXSndx/f1wTT5w+YmX2f5P2MJh
cSprnasYK8/RY9g2jRbEtULDMJkcmvgaikqBK/X7jW4y3NaigvN9mT5caPnQ3U6hFUW1HxAtfUHL
mpYtdw1btvoB3ZCWZjVXZ+gpDMlj777GMYUly/i+VyVDr/huP6ZeZYVoEFb65pIL1aaG8xfrb39l
1nLslVLzloZm75GgUXWNwBWwWUY23MsM9kdjipLq/VtTBsA2FB40I1L5PILk7G7ZH88agR+2Mzqk
LQeNycZsrG/xvqfv+Vzy1kkOb3uaVuXTiBDXQjOBOP5KLf6reCBJ+zDgvmi2SKbOPUWRB2zwFDEy
3iwGaFoUyj3WC0tTCtui31TtlCWuDOOc5h9N7uUVkp8vj1bVqoLroYC4VaMl9mTOBJ+Bhqr8585b
ISxlwHddPwzcKAgL+hqOv6H7t48sZncrrFLrqFc9uySaQY9ZTV4ttZhSCfTb7Qr0nhoHdWD3/zzo
k0nKvglADWLSrADYbCwGSifEBkhzXG+crgjaKgqBpkuUgqfFnfI15zXbWk63vEFb/XxwWoS4qms/
P9FJ8JynETBPokB45Zr40eNC+XV6rusPvUebIRC3cqwneqb+W3q96D0EzB9CNa35qFwZ//KoZ7Wd
C9FJSIPy/rKoRGUP5BenmyZMuCndNjVoocUDgKcwWjgjxg/ep4sIXmg8+BCExXvr8k2qcSYQbV55
01+M09kikYqRinVbDB/snSKgeACmWPI8A1hM7uIi9eRUCVaHhpgQFW4udDnq8euO+t9Hf4jUNBUb
aGr+A7rXl+gzLc0jETFwBCw2B3C4ublIzCr3qg+jZG3WRPhJxucF2q9a00T/7+ypMMifXfq55Qg2
KdRGU80ZPs/pITzrWAzbT1CGF/AK10a95nkdSw/HkP4+KiXbh49xSwsyPLj9hpuIoQKcN7nRI2US
JX/IwypTTVNWY/g2XtCHyQLLqIWF0lhZO1DjHMXxjG5Ij0HtENDJ6htO4/S4mhCFvFYoCToWcb85
9blxgWip6Ht+sNE2J5J4ZF2ZXwKWIVF4rgs59BAjZFzwqRGgJj5fTygt8b8yVEn8tx90ZHrU+wp/
4TI6a3t2GfG7Gz9yDWO5PahmnEt76IOru33BjpXMC0pKQkLiD6oAocI68rIK6qOzrx4BeisYqtxm
npc7L0xZJCx3SVnM+un0F2WPN526DLoL/5EWHyE/fzxTWG7EOvl/QUPSZMDI8pxzJ2bNu2mRn5OA
xBEuRxXgISbpPW74IAi0TPyt4+ko/yuFmYK6EnCRSFsGG84zYCiUCIJ0w10HDDtsM0/afZ9qJCWy
OvMCVMhsJJA6ZETK48RdujxMUXrn8Sg8MYtFnNVUsKL2ijqe6wq/YxpSqyD2tYU30bz6/CUFGeOQ
zG3ReGQXtuXCG+hnhuexUx/sCY0E3VepuAHo4tAR5zkrgH+RqbJSgT+BEybbvnHo2I0efPWO/jFs
tT/+Ul8l61lBAplbAe5V1WcG8XAhMVEESlNn6Cl1IjpOMnEWL5yBp9V7MFS5KdUCG93E3dY5kxBL
EqGm5grb50CAKuqGxJIscLP44HTnHX22nSp7gIHcRBVxhFu2cjzNLqLD0CbD4uH7yQrLnO9O2l0u
kfGYoRfNP8fsnfHn/jA3J/FzEiExsdb3nE+w1TWmbApbuxjHVz8IJDofQl7ey04XcMTaVVEnpNG8
ub3S/jWhrZjIX2EKkP8zA6XDtiaAjxYZ6nxxY4mCCGsFGXk0o9gRiejO1SdFar7bpses/d3A4BiH
E35qf4aix6JHmF1wEa/4sPIVznjL9latcuDo4a9OfA96cmaGL7K1CqPobfHtKD/rcz7VlhFxWdHI
f/et6+HSrts4Kj4Kb2H7/AfqVylX8e2GjzKxp1KhbFKTKe+vf2ttSqKnsmVSLt8ALHoFzBzvUNCM
xoOQoGPaZ8FofCjBjm4qOXtLxuH567CquBS4vV4OUuwwgJqnlUNjoJcV4AEhBUuvldcQdb3wn/Rh
7le8Qlrk9dxKhdO6AXuEGXBh1xTAmoEUwhLlOUoK4fBOEExLi4lm0PbPb0Kg+XAmFBjOLwyOYt0B
lDjof8yk/qggiqEaQ+x7A+bEESLKLa2/LgSv4DTnG52mqMbzWf1ExCMq8w+pcEiYzNR2EfW97Rv4
96Hbh6K+wSk+f0fuZq8TgQneIfPgv8Q/EZcA/xl1FoB2xEPLkrRbNSlaMATXbhvFMJRAhB+/Qbr+
jHAEqqDrwoJNgMjvnHL4x9gSQsF0PwNwqD/y2RnZbdRW4TIjOichBoYO96ulkLnw+M3EJNCGIqfu
G82Y49irsccsukc65hizbYuAU9OGZkM/u8zxCT7ar2RJ86dGQeP0yAf5Hwig8XUzNP4jRS4jud3G
68wKhtq+1au0HUoZ6yXWcRQ7CvjEmINJoklxaPbDvhv9DAO7u1DaNiLogA03qy7jDqgvf6dylAT5
q1JOhdTIR3Z4kPrndlc3XnRGq8ffWIyLcNqT9z8QxSM7P2R8wJJEaDMoSGJIwGM2DARL59YSA76b
lF5bdgP0Y3vv/xO1pdAxFSxEyAlNi59ZVaJ1DsPoMgLVdeUwHr/qgNj7tt8juYc4DK5bGdgKSW4n
EGI3RG4sG1eY2x1W57BF+27ULdBuN7Fn1tKUO3GUAyo4gDf26P6qo+hsObYtOEuBOxJxjulmxW1v
i2xQQXfiUSlOBEoFBCZB3VTNKAqPy1HzPj7H6QmIlE1WaPKVUNJqlBWAsyWJk01MZXtr9DSWU8zv
4x3JA1M2dUdZg/ewoaD40MuX4lpGOjgq68CL6mMqAbAsnUD3SFvxtmqOJr2/QrJ0y6e/aMjUrRZD
PiTaZLEXBwy3VwqDr+Mg2OnDv1sMPwPwXzQhcdtIZ+cN7fBSbL+cHmFY7GtA/ELflaKuhadKRaWa
/deGkuQJFIxcz5jLrsZwLyZVtvoQwjVv+kGgK8cjJxTfjjEEv5a1+nBIVW9GNcjrvSsF2/dKA2IA
IZZhrvdZxhPJURiNdipXgSHSk4QgR3Ftddgg4ilD2i6ep+O6Kdq1WSwh/3ORmB/mDIXUGIJYSI0o
FrN3i2dsgUm/HQnaT4W75gDBlwNslKJ2G3DFaUg7hImJ2jYuM3FvAN26rMZ78GeucDM/JtvZzH5E
T9GKD1Mm2sZUYc0jroUc6sJKNjo/wRCa6g1unH6bi9RoQuNDrdXIA8y35O3g4nsNhLzuEUx013Mk
He/8RrhrbFP3cOrCr0iW+82q33gCef/vTqLCDMvY1q1wfvfY4Q2P5IGzrQzEyOP8gTbL0MbN9Cgi
ivPQFOnAzSnYhA02buWBQI/vfVQw+XpralV39T42Sz5PZbedXQsYTpiPuKhga6jseKXZyYV4RFo2
dLOXzjp6OABVgQrYhWBfMILvMa/+CrOEvkVg8elj7vpE0bZdjNbswGCgWSAyM2zowh83t4Rxz5vE
bi5dJ0qJqeXInu9f+/B7uuFrdc2yaf1yPMJQ8Qi0CZkp2dt96EFIZ7yqyEPFfbU5kXR+JZvfwQHQ
DNxKFnlpAwcg0/wFf/n3a5ZMnL03Gk4vS75/kTTWM7TrWeNwZ4PeUn+ebwZBNef+reniE5yeV9Nv
qagr8HdhQQeoyETU8JRCj5xpilolAdTRyJDWYg68bCeful2VieH5gmaSCUWLt6BiaqFERlYb5Bcy
n4inxC2rwyeFb4nviTR4YLw38QqmVKPT80PqfTRlrSYfGaLN6EsOSWPfxp9ouRMjwbrXRnbaH9yQ
7k8EHtlOCkIxVGta3Ta3sP4uqQENbf1qmCvvkWfm1k4uzQnSdUZOEUSLW2JyJfTM7qIBgEsx6E++
9a86zZto6vSrZukigmi/vHmUvWO9VvIw6eKUMgCapBDlY+KhUEn1PbY82I3DMRL7+4Ks14Kjc/nW
MbD2PjZyXBQi6jp16cpEUCoILpHJ5aVczB6hxauGFfd0EQL2ohq6G1tNZQzbnx9RRy1tkWhoj4cd
UsruV9M4GWLTNOwZnbSBTSzEBe1rf9u6KL5JwjL8dRHTEXkGQqgO/qUSAkc8m62bevSoYjX7NWo/
FytjuCWyBcM/yZBL/l6USU0Y55EoEClMVlNAzCA1vr0o5u/qrxGm919rO7PykDBTCCzcsWvZrpNZ
4CKc+4brvvG5Y0OGxsP5/NzGVGTHb4DKAvsofvgUEM/NLZqzzNURaGUsNieJ/KEo906RAjbfkljB
t1fPQeQL83BIh6XkFUBCnDjkHR4H4ck26wW1L2bR20xnr9ayLcRe2/UoFj606KQOgx9yMhsq8OHe
OFSPo0lXv4K+ntLfxVP7FDneGYFBuK0QzGu8h90lmilM6Tf3sgPrqkgGRPhzJu/lfMe/eTj1pDgE
sKhFesH7zbyuyl/FFT2RIf74SraywmIdGb7uu04TZrpvCELZEjm7/MT+2ZVTlijiUTXyCgBOalJ8
WuhBIwJqr+iZQFMXmGx7Va4YSDb69XNm+SzW+mMfW+DZHlMQMSFExNWfHwMs9FHI5hRcpYP4biD4
VLbA9VwlNDWDHeejjAPO+ha63GFIMl9NJ+x7NNzN64dsUlULmNF1rdr/KYTPRhgkXAREz/l6juJU
vQ/yMIT2vc4cTQ1tO1XkpH0tndeEdOc4fpyn7iAo3jl+qVPfUPxHGM+YwphZG/X71ykHkm6boNTz
Fp7wKx/QTaSOXYjZKZG7OTH3b81uO5EVLy31XuXKKMEcbUbj7CDT5Afhatzo30GjidHZ2TVFBqgi
qQSr7S01qbk37mpWyWaRQGs8ywCeD/gnC01/w9qdOq8X369+86oR1tPrQwMyLOu94eSn2/+IMF10
1fOhFIdSx1KAwqgGos8wM3eMvzEJmZBeSG08od+8X9LtSpOeA4/5S39aPKowbDdKZcCtGimW9Cgy
MHOQyHjNMsTukckqF5U1jzx7VSV4Tx9VLQrQ/5A5uXQK/5H+hi51b+bbLRnwuerfr4Wrcm0uHcA0
sFT9qQjU19SpRfaumRFiI5A7t44R5wa9Y2VICsxMrRsc3B6PPl1AwOw5TO+2HoaTqmCcMcLcj8LT
sYzL0d6a1W5DH6pgNYcsZawcnJ1DZ/W6i94bsXzYTWuSucvts7r+dSK684lSCG+fH9MvLoZpH5Us
Gey7TStKRnJ8M9BH0a66hMrlrA0NPH9dXKZN7Wy1yjrSc6F8Znw1lIo5Up5sRugCpfCLOS5TGrEY
oVLY+DRhmKZo8JSz/C/zDEZFTYpogHfl3FZxHGMC15XS513elIOB0MOTklIStVdF+Y9RGFl+OOw0
RWgsWKQvlcPFcklHe738AHTc+BOaMKD2HqAxvcRYRg/Uo9uSEOd8LAwyxQVQgYUdXFa4J69BuDW0
HPScsOA4jdIRnCjoC8D8g5YWr7FQm1vlIpR/gqqqMK998WtQPINKqavfLo4QogFOLsh1W1DX385l
21Bq1KbgnNohyImMr6DYjVKmPKVyo2zsYCor8u/dpl6tk7korh0SV4hYizptdyJlJ/5y66ZHbAT+
h/ZXgZ5tXqvT9ulb1dT/pvX7N7SRASs8XFh15bp/SPCrzH9vSJquPW7Oz9QzTr7/T7o910xoaRYX
aGPW/dGiKxGOlU7mm54IcHiZgvSRkZzTOOB9TitxpBuT9RDX2ZjkMZHyjF2g668AuF0UY1BPP19A
yYGPVCHhj3aGxmkToKFn9T689vq+sVTYNrx0qizpodhvY4DgxcDP/2yt24MYB9C+HHOGGiEnOznx
kBGTZvvJ0nDAIZj9y2Sn1VyCwaHOibFHCMp70c/BxNsuW2kvUiTb73i7KFX286zoCo8OENdk8mLO
J8UWRRoZheTuTgBUS3ZkwVs8bVdC7WD7qL9nQcyyUT6A6BTe3c01MadTNr/q6Yaa8SIEBNtTlv0D
upn3W0saUGujUxO2sx9pqYm5CltI5Bg62uqho6CsVFyfTQARSJo8UGeyzweM5JWkfliPYaNHVRuQ
Vw420slQxNnEHqHc2FKsaQxUxKj5abKl8CuRapzRsjsWunHFKSzPWhh6w1Soy22n6V7PPidlzXg7
T4zRlz9ZYWFLiGRuUxd0aKTtAIUdj9bPIFFyFZXdSz0Vcay6QXL0bME6S6xos2WBydX0lRpGOvan
XF2zROdxfrKVYvx9BzZyyGGGVv6NjLJu0Ca7sZanbeCOoFjzMXxbAmGLFDG+Z9Anwz/aMVfnnHau
0i0l/acrbnUFgseF5Y9PEUQmur24lmYnHXYdkouigLdaoDXp2mCbLJoYOWnb6bWZ5zVAVF8hLmYU
9D+nogkRve9QxMUyD33sV1uKLCF+k3x6l/Tq1czynQIO3XCfV+WDv/9WKlZXhRp5ij8oRKaOUG2Z
vrFcQscEkBRtX98lVmbbnY1pFrRVkzyTIr045wj0qSAXbMjBkmySMj/4Z/AXXa5/kzFdqLOLnIVV
AWHk8LztDinO8flSIhPVWO4cqRxeA5zH1/HBznLOacvbyHFuXCVrJiJqsOXd8b7A9cU4LV1KkmSP
cVmvhi1go77tOb8QCEeQU+o7ejjGTqvkkbSi9zx1+yt0pIJUeFl1q7Zs89PdKJB6zqoEFUq35snz
tBMIdsp78qcN2gYgXr5B0APuBiS00O2Qy4d/JgjYar+Idc/8F8M72j9idmwTi7CweUcOA4716aEW
3R6g1GI80NuXUCLfj6bdTwQHtj6adDcfQDFUDrOb39mbq7RnlcK6OuSZV/b3BxCb82DwAdl8NrzM
1MfgAmDM/PDc2g7RzGEtJGgIG5as++aqH8Ekwra5EF37gGQjGaigVCVfRHgKf4Gs/hPwzK8bo/7g
edyJztFoZMs4GfVIAfxgyc6O5yoyf3WMthD/jpRH58te8hNUNz/rtzZR+IrAEHT7e+ytXC090Zoc
BCSe5rFE3XBl/kdTvS78eb+IgzZ6swzbXgi4bj/CA4ySj6bS1IQj2qLcMpE9rdMuhXC0o3bLa7pF
fsHDz28I1IoAype37bOz/36ZH/iQRezS54KiaXEOcUKPMZciKCAUOpNjovccfpUs8SBNcjxbZq5u
cFw61MtZoSN7I47NGvAcJRs67ZmFnTnh1IuQ+oDa2GCctnXii0HwkOwqI3ptRZsKkurfBIOtumYm
q3E8xF69FTPNff01N0bDU9HqZNLmhVT8MObU6eDtDLT0mu3Wyd7VPemnmkB2Bhbnv6HeOE9yS7zP
djsuVcfAXjvd/yUpkJlMxxT8qhY31PJxrsQMOcH1Rlq1jHcqnQHldq3OKQq0PHIbR+S4qK5S9/4r
36TbY07SWe0JBsfXbWCv7LkTLkb2imzoBT1zMLspMGg3X2c4FCO9XEeeKndmLoQcg0XjxKndl3hv
OzSoC1nBWaG+zTQvlazw+w9QLqMn6vAbqhg29JSN+/wUE73lnS6D4i8S8nS3spvIbzF38i5VIKOv
EsnjYblvw1bMS2AG5LNQ76XY0zscvHG3TKoNxR8KD9AwRcd7UpRrAf7mEfK2lFJyDkZOBD5+KKxg
Epd81XAafG8QL7TzACNh+f8oJUxfsBCbi/XQtY3f5mWhJPVebA50GcO0b0yh+IVo1tYILK8J/CRa
ZRnMaB7wgc8uadbqBCDRITFfIsMs7Ha2DFkQUN42dgS8Eh1OrzsdQkSD5AJu88Ap8ClfpMMPVOIr
ANfH4FMKZjxnIQLVnD9ESLVWizDJ673YWlmJ5Nx34TnLlS6ArCmm9N0pBiKiUy+V/SKlajxD/yfW
9Bp5d1ISOOFVrbmzIn4dsYWgVtyDGqlaz2GGzps1rlIPc1gzLKUhAtCfqw/FwcTmStM59w33D/pn
vN8yAClhuk7RKwF+P8XUfTp5Pekks9WidDPRt0k/UrsyvyRA4trqL4pw1E08yAVMVVz1jS0wqWqR
wmleYZWVdpfYrNdE1weJpUYzChlcbnru2ib9qEQVEAihOm3wtYLBmkqIuuKWEo/0S1mmAhDyG2La
NcYcr6OM4TqnsOfKG3RRfN8mI16WyP33/2bMLIST7dxCEUnLyR/WHE5PIAB3hmNSZdzkhtbP/BxU
Uw35q7Nxnu1C9lr4KkNulych/leSIpvEXWDKwO6XPAkrF5oroY6x7h+4pNQ0VbG7GWlashoCiQxb
jDL4rib71HR7alGgIG2wUkCBI9lKvodJiSUWJQ/cM+G0kLZTHxzgrv7K7AL5AjOMh7MFbpT0
`protect end_protected

