

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DZrqnYwqMkKoBvgXgaWSB1Gvc9B94Zr8xHWYvXS3Yo2in98iiVsrSf1RUePWKa7hVSyhM66u+GP8
6zam55ovJA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
paoR3khjnzY7oR+WJ9YkW1A7ZzfFLvvVEXiP81AieLlGnfQuqZTzy9TqIBQ7d7KWJF2u8/GBJ9gB
S/XHVoSTyo6Jte9XVVsqnnFiHxvEAnWbM2e9+Vyqd/Q/lFB3TCGyLNKIFNdGxyml1xea2Gq/DUf6
P6PVaPylNEwivSbuc64=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IuseMdZSknnKUME+O/YmMG9MKbslcWjYg4y9t234jonRTsM/8uUOZLlJPdAz0Ojsb7gi8Afg71RU
Er0Jr7fpQJ8YMMDdLQ9qwRqf4zAR9ZhntG7zWMIroK9jxtC2bvBKKArJREVpkzOWU1g2+f7dJ4FH
ubSzqp/ur3VRiEL9rSTe80jSph04B3Z7vLg49YvLUGmYKlwP09xV4/46qike4zQtuofkQ8/u3jTv
rlLcM6RtgeLWfD/CY/EWIIuhTxeQiucCqPyYilV1cA55FNKfdMv57PsY4PVV/CwLFMYY9INUTcQ5
vlvEZIaCBXiBH5TWThAkm9erewSr/bL5DW9PTw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cyY5ZPlO3Eo0cmsRtMR6yuz2Eu2e6S2W/D+8CcC8VsHPfbx1fHUAOMrMRz8rOeXuKPOa7h1hSFcJ
XZ1TcAU5VIvCkM11jW1o53hK8qachmkkZZnfj8JtjstmyVTyWri5LmUnPYRufwJmQUQ0xqMJytkR
VTqDp0ZVnyDWp2/qKN0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WAcKeockg4TPNpKWNqCVvf1P8zBdM0HIqALOQnRkxsC2RA2Dy+P+XMiOG7cG04xrgm5iFejfnqcO
5lDRzw1y2vm9IxrTgVR8u92CBfbBU5si2daX0ciu3+tUaMvbyjjRBHmWEJd/+ZgwpEBd4jKx2KQp
YmRUDFYL5WDDgF6aGgbY7bniF7p7fSFQgxz06UbHJt/aNGcXnfge+DPA60LgmbiAZYAbqv+bSmqg
gA91XQkI7oyEKtZ35D6ZzgJ25i0EzUAy/u4ctGTC1xnExC071TQUx8Fakynqcki4h3cwrvs6RbsQ
1XULS0sNZpYYdAavNOXALBW23U6uD7bNRcfAog==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33936)
`protect data_block
awnwjKz/RlsQyOLwB5mE8iSC+LhjCMaHKoy45snzIjTQqCOS6C0PcTMwcydn0NsRX5kzVCyXS/cG
obgFQlVdcnIaOkUznA1xFdpzEX4+9b7tEWFutgxHPR0g7MOk1QzbkUwWCi8yor9vRnffvvh9XV6C
DZ7UhtTGLcTDytvoAOpnb+ZaUrqdv9yWQjLH28EiH/O1dk8OtMXVHMa34PFYyWvVi8CovX24QD5z
z6zJrW3o/QtOZaFRTo7wMRyyeSrxeAjtcWdkxfuzIhjRMeYzZRKCgGeLnX7XH6vZuojmdbGcwwV9
RkcxXe7HHYeXDVJiMGah94Q7Hvy0r7yxFRYTQH4rIRH1W50mYM9bAVWKjHxJ0qUn6BMSphYr8sge
9UbmEAXfnixospwc7P08NvvrVCiB60/uLQwf+LkQJayEor9IqiwI7XcSFxucwLhJ15z8dbI8lWVB
KnwMyrS4nfLG+6sMkXfGzzbW57OQwp9mqoqrEGP97SvtVbc5zfjcR46fs2OMm8ZIDbPwiXNfdY7x
/Zcp5zYDaQyhNP1rjcfjQYNMennrMtnzDgg63sp8rheX/8DgKrLXqO3NBg3/JIenpS+RLNDP1TK8
+HwC79hl0+v8Zlal2YWCpf52rIkNenn6pXy+lxcqwSKzY/1j/FpTdOOz5iSCHXcpX7/aoaHLPN6t
5STu+YnUYuVelBZpFKlNKfdqUY77fN4Cx26jm1yYFMCU375AHyr2ow3ckBj5xemdY9ORlJ5JHJ1w
OIAevvllucSCdQcrStfVO7Pfm1fGeepyAqMdBR1GfTZzsaeZScNqUkQIj7TJAX3SykdVCDYB2HVb
fRkFz8UKMCaeIjh6an8JwzB65snPLAyFaMupMwP+7JH+iffEuSzs9XSHeReSxFiVZSUjUDnmGsfD
PAeuvDtdwzvi0gxEBRTw8543V3ufNmHbs/VyMmGj2ITu6+D4vZcnOH3PqpmPYcbHr0UDoojfqfC9
N4dvC72koxwxLfN7txj9e7m0uaQW6xl0KxJBEwsEttp12G0MPoZtYjBC4xMubyxEBmNrxA5O0J9e
MP+qnnv3WRZJ8rDgiteJ15imwPQfyFRKnoaXA9VM04Rx+4GFN6bHGWtHPQMPFHm3xKu35fMka8b7
jGkc+GpOlTule149nr63qlqb5KbNLO2MtxdtouK/TyJ+sDcIsnxmCn2u3bqd9xSp4kkH6u0A9R9L
8S0w+OAiRX+jSfjXEvQo5ZTyN0hZueqgp7rBV0ggvMYhjnmAtDsm6LS6Q2x0PrXNsX+rfTA/nF/1
RUnwlo1/uwAchavcb4tOkfQucK+TGwMZgaK2jqEtTcABDaIcqUihcPJyQ5bYSIDx3yFAv337Bloj
LBDtqK2QKO9qMHmpjt2p2HNc3F8BM8xFsoMu7IFsg3sQcF6iOi/D4u9rhrC2cfyxvHscacoaDJ9z
WYKk4g7qf27IBogC8O1soumK+NOtO3YncMXbemkgGjyGCK+7csH/IfdIaiGrrqt0Z/Cps93VvYS3
BZFCxweBFwA2EiZIn/hqOJhFHuPeXYkF2Nn8DOkdnoCrd7zu7mt2tqVeW9aT0jQtazb1mhahxN75
gIio26iB+YerkrBYhoTtdtgjAOtvLMTAKoCzCUEJp3i4Y8EDoTiY43CQrT01DMccwnNgmZRdjSOj
l2EQQXZgjYoLiI/4K+MpOqtI4Z38Nug2CabAZDOPVp1YSx1K+AEkaGt9qMPgMTeJ/iCCwwHjYf4y
Ln7zxMu2zxfCzhI1d9xf7hbqKd3AZnl8ouMyF4KQCKP403mDZDolXf602rURFfOpvIXCU8+BdVYa
TE7XqlNOub4EIYFEMiBSXPm6bz6crc0y7CUElDyg/IKQ+eRYYfLfARgKfasJrH3DiUcq5pSgChFN
IeKC9fRonLtgZw70Ouio+S/KThBoMB7M+ffZAnVsxuhTWi+vgX5EeChZurhNuaawwO3alZher53R
dUPHBaacc6IlcOigN8pJYsbB9klKyC6b/HDW7yCiMKCLFQheKWMIl7z1jS96+mWeyZXnbcsDw9+j
huhuJWM5HKXJAm8dgClraKEJ+dS5GnZYQBWeZRw5la2FBFqN4uHOj7r1MZVFaTTjgRelZSxar0Ch
5Bl1SyQtGJQX+VpAe45yQUHd0XN8Qe/vezGCLJ8M2ot2LVaED4ClI8Um03xysCQOtly2Nx+CgOBz
vzR4ZMNSC2OhjVrU/WGjbFte9fg2fHuaNqU2+gMwz4I5PLtDI7d5mVacYvTyECNw65xKxKpAywEP
OWSWrwJRlbWOpEWDOxnkQMnyk46wexs/QUPMo9hYcv8yySUbpQcObG3Pe3bh7fMmEp9r18qHP0y/
PgHntKzEri4UwM8RWk71IOj7tBol6ghxarEzL0hmrjiquZ5FUeT3MZvT//0zMG52dMyxdO9vRa5n
hJXzVQKj13h9mCH/anroHJWwCgUqzf3hm6BZ9F3yYA5HEe1cZgwOzF+c7mrLCSFphcb5h02F1fMH
R0G4YvyZfJGzAPuCzozVYQFJh23WwFFIxxOPZvMpNRaBj5uhhMIzar9fSa7VMrNkfCFLw2wR7c1e
NJIYqoD0OZUb8xqrzsNLQOaO2Ya5td/BSGCBSTVW1TiYy0joPIopJS12GqmLw7OOAKwMDKWuofMh
KJVBW5oKVQkK3krVrsiUPNiRrChD4P2g1AsHuOeh2+EEnAT+8GGoxu5ujtT0Rs5DUclsAsumoXxa
rh7CDKJs3ALVdRQyhiMfI2u5ZeNCh3PJ2K/eFjU60nUGQuvvh3HL8GYsKZzbtxiYu9tcqYbch6qU
iZZN19fxu4T0xwE1fdtVRwGhfR+6BQDPBToOhQ/1obHfxXld9r0XLVvgh6EzKl7KSgVLlog3kVq4
zZmRXrMdI7Zem85t2560ZM3pkJ/95lXmsaJO1jBe5mH4P2swZ7WbIjFQwexe30+q21U7qOkgsLMh
OWUsKRwCGsEyOx6XHVTD/1iBjjuiJL1UPPifcOQ9o/UnjdLsH4CASwgkS5/bhGx4gxBAOkuhyHVd
+sH8KJq5Qee5EEmy/73i39ldJeFvjOjwK+z4bil2uyawoH8A5n9GT1D4oG3tOh3iKm7XrnEYd5lo
QfqYI8dNnXN+vFFWHQ9d9fpsyk8vWqismGgRTvsV7wMDxVDNBTyDTNSkHaLgCljTNwbSGFS4TFo0
HP0Eggd34nHTexdJWRPp0pOllOtw064RvLdk7v8H/Oyllk+KruyjmQn2arpQPn5eEb826ZY50d2z
iOQ2cmXSdksb7s3vrYI07zZ5vDIFym9u0o6B+j4WnD5c2d1L9UjA0+4+2LxyCuNA9simnPxxv2Pc
PCKUpsrxbW7F2roQi3oOh+JSs3BQ6ZrOP6lfAy2xxJwDAZvQokEtvwSn97+vgj78Prmd97cpKC8f
9KG4LfbI6TtHn5k0dU7w1HplNhvT7Jhq4Ww2DXLbbbVSuQRG+JWPzGdM3tqXPvYvaOBn05pCtvtL
ZYAbQ0187iAirguhQ9F+Ti0a1gbi8kCLvBdQJ90i6XD5RjHd+ukfCJD5UJY/ZFimu6ORtq55E6oF
4TdXgUEPklBYBGWFg3/ZcvjuTERbbazKfCRFFXyOdxewgCh4E8fG4r4CJUfBDEyqB8UTsGDWbNVz
mJ0aAEQKY5nY2HWi602VVFUJOfW7aYd4cm7DsZd13EvW+Phdu6jPb6Vqs+mBguoqvsj6eKwg+lC+
wznUzzmrnR9r87BrnRQytTIqcGFmU8VDekqhrA8UebWgOjP7+hcIe8LxY4Vt19F6eBa8cGwABzOh
Huh5nOMd4gIV3EDSKa4eRbCTvIizu37YDTGUqOVay3i/aSsaC2lF4dtBmy2dQHXnb5eXb1dKs89M
huvJ/NL4qt+3uLFjwEbRffmRAm6DHaVsoJGTZeRi/Vwakwp6+NvMSCN4Ihh6mDL+gt5DnFGCL8Hm
xmu5t0/T3IPF6mS3yQF5IMoZoc5rtWII9SWuEzNZPxMDJhJnbrus8mqjQLO2CkVmnD4D6Kp2dP2r
DtauWjfEn9Ljj0DNa14Mzd5C2Ec9kLDuXtCvdH5MxbRNBhmuaW2NpPHfHC9SRizf5fWOnhid2O+h
w1s4D5fiWJ50fNCCa6Ub31b63JudWw1Iw2gdLHma/q/h76tAzKzmuReKHuhtszS06F160UPVVzph
nUDGot7ZZBBlvnvE7+HByCGFABJdS+kaIGxTURhyXv0a/BU6ACdK2Ah5E6nctj8HZY1n46YrdP2z
uaRZrPnLev/DMYEAFhICmIlnpviPcmJJGZ4xSgwo6QjIi1Wx/JnpLx4MXIsMjptF/ClC1Ez5zECp
BynxD0r5enFmPmwD7NTVMjMGyBStCBcvEyrsjRHb9gtXnUqv3ZePUwo7YrIiGWmZj2nZbDCh2r4w
58j/LBXG6WjV6nMVUtYXpooT0P4iZyjkFvCCIVZs5rPiJZbyyueS8yXw4WLOosMPzm8BA/eLto54
Q0vkn95TQdu6cRnC7f2qy4aF62UTq9/Wg5JhnS2YnJEhecx6UZ8jviMyzki01ckg2VQLQf53fXiU
f+eJsqzver+Y5n5UBeMgfHswf1Fs+y0gGE8am7BFCko6/HriuQcZRPGxNtskO/pLmiGUgZ8mte9V
06L6HX/lDfh0OWgkCOqvabNkwoHXAs8HH/s1ic73VQ5bjeqZBcj1u6g7HNZo2OOT5ySnk4CP0gun
NsuxH16UEJbEA/of91MibiCenHPaSU0z6nTBGACdKsbt1gSnlYP+g0CtOTFGhRfPpVMtf0jZbrjY
EvAtrWcBaGHduygD9tuxHQGy4KT+iWxtvnqcAQJ7tonZAqCYOA2pCYXiH8QAE5RQeRgHgHR/VZ80
eepLYwsk01A4Qf4KS9EvacHYwlsBTakY5b2EXTms9zZWhrswpyXls4k5mSHOcLs6KOpl7lcQdqui
pbII+iTPOKrh+1dbVvWbqT6qhMfQ3QTX5I5ajwo3oqrhdJrwsrD2PRuXXi/JE+Xv0f4x0MnCZ6Q9
aEtkWWTOQbnMB8y3JJ9Hvy7fP8G+kT3IIreoWfazqSYbjIEnHrf+OchH3Y3XJ5+66tLoCwK2HB0+
5d2cf4COdIUKqmxhPikt6r5NXButwNyjO2XvLFbPqwBvnZOlbvOHI73TFcGKXRm7TwbMag80qz3B
76EjK6kv327snHxFlhD34/mCyjNOvFF2DULURpoQ2BJSe4xaFDSGg+2us64u+9Q5/hw3UHbCrLM5
4HePBfNvsbkkgVG8W0tpcdPhaipYl+2SuLIimJwLHUadM6z+hUjy3JDIt5kriC+fRPxM2nRdIgh7
zbheji2PyOojTJkIl6lrkLdttnqMQFkQ7VkhHZ6IGzF9asrwa7Rp0dCGLQQvHJdHEjakuX+RwZfo
PI7Otja5wu0H0kVmruOO2hE48XKHplxGUMvGmAfglevvkH0o14gb0R+dajMnuEo8H6K4SirMcN8K
M2PElEQlI5Y7EMJM9EFH4EkjYwWEZqpVcXTCkV9GwETptDXEgpvPTBNvdiHPV+RIv3OnJMwEeRo6
80ctAOIpKQAPqC0hmp3ic+jVXyCGnyZin7krRM9GZc8jt63fWSBw9WnrzpA2rDsT2gyIl4fElDbK
O1Z8/h0UZsHX3bQAWLV6k85phsXv6a4cV3CKTNwC9F/co1qxdtvXKvS5/j0U03h3aK6o+B/ihLah
R2ceKPVhKWRElRWzgRqH6fxP2MToTu/tyHdD17SuJD+bVryj6S6pcFxMVf0kPRUEmz4LdxQxIghT
Fu6J6N8BXEkggII0zlchbQNlGPgvtaOY5cMYUfcXw3gVeHedpm+cigU814X+9Xh/tbciL9SLKgHS
M1YdGAvQD49c0d5S2a3kV4UTcKRTevk7jthzJiUBZG+1utsT7ysOoHXBqDJC8U6Vr5/P5/Gud84J
Ei98SulNTGNs6c3OAZbEhdbIRdodLuNIr0IsmGXDe4OhFRa5RrIeJZcgvOHuG6bnG3PpvcgH1i6l
FqJOFGWp/kyYNzeJXTf8qkNvPtVuprDC8e78A5ud7jK+TahVfPXqqyNuQzLigJVaLvesNKcUI/wK
edz0eDXd5o9vMHMuf5Y/VL2ghRYwFvnt5FYM5txPOhp5Nln+QRsQGJLGM3ks1nnx22FNZ2jaQqvX
zLsXW4JoQuuRl9DpXv45zHHc5BgoadB1DH4aE1ynEBFkYmr0ivZE9wtYBFpLBhW47zvWqm7QVQM8
Jw4KedCID9wJwcpzrAIy+VWRgQjwul6NpwGVR8nRpYI5fCprgdRZUpArbuaWy1kg9rks3fdIP1ks
spc3EmQnEgktRZaQKDjA/kiLmXJeo50/k05i6+DoYll/ImXNkyyDrt/xY6E1cdNzo9clxaeoMr7v
OycPQY+KHyny8Uo919l1WlVY4U95WTlSSXXzRlOrrK8cX1aKAYKWXv72zZnlS3fgj2/zHCCIm3mt
WD4Q4IACYKNs2hCgW87P2xBWH+83yT0+GreipNxCoEH3vd7qj6Rvv5vFng+wwL5gXTdC0PiexrSU
tp5M7pqUhPJTYTZi4YjjCbjG9Mb9iKDOu+96A1sNtNQawX/eqpscWSYZOuvxgfLviQ7TD6c9EjPo
LxKBpvK9qfeVIi7qeass89ALLSb+oiitxyeFddXGTaZcsPsWpeFL+dRL6EX1OKGv0OQ4O4PmN+Qj
I4p9h2UJvAA5Rw8F5iP387TETXAyuxS2nw9cWg5GRxdiNXMFVg5l8oXJSIz0mTSgfFgYr+gHy4vH
HFYP6dA0CSWW5r7MKhPxnA+XPHGnK8Qg3kajXVo5+dUozbIqLJ8p0wqahPVlHBAfIWANuCy51Io3
Na/mcABtGXEChs1LmTME+4q2/dV3zQ2turqDYxNvkkk3bZ5G8VADobBy2BGPRe0dUqTyYZLDnpxv
bEtekR9Ks53c7+IPM98Ch2x7rUd+Ops2hbnuFXbh6jBhC4ja7tJ4Y+/lxer2MKS8xhExUFV9FrXI
Pj4ZyautQlR8utvvMChUwIE+JCfsY70grUFNtLWT8oUEyRp2Og9nY0bEPGa6jOs/YYm4doM6Zg/j
EEtcscc9soSRssX+dt7H5g6GHKEuh/tLHqvT+qPlqH7xfFvcsG2le5LQsn3JBAJipn4fjyTTrLAL
wcKgiVUMHbXRgZtfwXYkRIRPkwKFh04wIuAf4Fx1Ol8avL8GvuKaGCEcuPABLYUFqn7hxr/A2uzG
xswzgGJ+Nfvtp/++6JtncTaWi6gpPcL48joHuWuh6bv5hebNEB6fucvYtuJ5klF5AIthTDEekLqq
iXu95uHqV+Fe67emR7VESKyKwsWXoBzaC9YgnkE8PeCJVpFjrbtMufhTUXERBoNIQ35L8ukP1v1k
744xkP6hbXvChRkjyhkhqgEvJSKzL7spEWgONL/NWWvMaXW4Ln6l1glb5Yqv53p8tbGprbHHTkET
F5Nj/lxvex4145MIRsHjGA/tYKsaHthiku9RlumfEuE+LNsDftyQF2WViR4hUZJ7fd0CyJY6N9+8
/oDYvkokFLfNajGnFllGxRgifAXr0WKSoIzgYDKF32g1so2IeWtVkahb64WBBBNiec4fjufRL5x5
NrcBn5jZWsIUU+v9KY/wcZ09JfVIIPe+GIffqhw2ZNMjeHHjxDusLSaag96Aa4oVfj4sCTTyUM0D
B0GYqnE4TIUjfXOlZNvCrPAstChsmLTwiZT/MFbY31Z3oKQ1Z1nrPSNAOgdKj2s0p8MZjCeX4Pgd
S4H8nw5WCMVW+d3Rqf0iuLv+EX/8uWz5sSfd5nm95PY+QVb/yAWfgTLNOzwCNXF37nY+MMxWkNc3
acGKzYlHq0UYsck5LXHRL0QjnxANPhP63fMsV5KCVmUUw+1nJJmShToB8tA2RTK/Va94jzZsJjiq
1nLvEI93Na3dza2PDaRAIs6FOspN+r3uDIbegFRCOOaAZrYhLBapPQbD3cGMjegEJbTd1oiRg/mF
KCZPA9Qt1NpebM0/JL4AfeP404Ix6YAk6Ffi+JkyWNG9rpISsXix2GAG8u6nAs0UGfx4J+BEwTGT
fffAb+FQOWWrLlvvO1xUCApKiO/uKGRsVk0WBbojM7Ctj58ak9YbDZL78LRBV0xGO2ujv0sKUHjy
pCV7coRRt1XY5z3gsp3RdPfcYHjcKyl8vc7wv6qO2OQXQwKdmPQn8/fW2J1WEgmfqv9+OoT6+vU1
GQSDJ6psouF3GVyXNieQ+sDI3sA0oWymSlqLPxT8CeNv84ChBIDOrUL/BFLn+pjJO918JTUJA1WQ
5oILgsLAx5I66aqhjCcF1tlJCDqg0L5n0RMLa1y52andx7N0Qufi43c1hRfiAd+znyiv+iJDGDqX
nOLURdWvBOnDjQvH9uym2UqyXbo22Lcd9onQB2wC2bPEQcn1aq/fmuTCU6Eoc9iUaCm6pBJFmF6v
JfrQbmrK4kOaCo432zgj4aZTLjjzBQaPDkEdcg9Y6ggL42MQij3e+yrWjmnXmj1xz749SBRGFvSD
zsM1C8cK3198cYTMzTS/vVgGeZMUxB7HiFwUz4QVzwfow2zvQhXDPieLfif0oQFYudnXR1/Xg2Oc
P+8l/fn9N0gIfFkmISEH0bDU3+5y9GvP4wWgL2eROgFlBVGQr/SGGiNj6XNDIXzSzfpypPsvJTlR
Wb2NuxvQ7RJVqF835Uw3XPgr05ZMhvB6TtA73JjsY8SRbffEvDZw3h7tzVu3oMs6CcJnTmDlTclz
R6j0tLPh7jmUc9kH+msMqaU4f0e6WI8q/CWk9trX12fdax2XP5j/U62InP/sl4Ly7O8GHmyV6d+o
LvJPau8aPi9t1ZuIDCilKQ/fJN29+x1hwaUQ10721ZcziyUgrTpnGKDClycOx7mR5rvmxctjJHhC
T0vHD6aaYHzQXDGgK53ErRGoWddwWyFmFg8cRB7Rhy0y1cYMpkcnOQBP/OwAWSPQrvFakDMjkkM9
st9UwVas6HkZHnivY9PAooa1g6a07PgBXaDwdNjPO+XKwUYLUi+v0Klldri4O+ZKWAmoipDAZEvM
oaqA9kv9ydHfpjHX8axE++8Muto8aqcOHj6xXnmJ5S24mSgQg5ejQKU8gMlomt42xvTkil2tv4zX
XVrf0WdXGJ/2sysc3YSN+vLFz9gq8+TTd/xerz2B+4zmf2E13P10Y2y2F3gxqIEKS0IFQD7DtWLv
fF+sM7QmxdLNh3nKIePkmmIkD4DZSl7Tnnwr0yIiflZHC4kuBPuO9OmhXiZOEZgSUAPN6TDaqw32
0m+ibZPZTO+GM+3vp8Jnqi8HufWNSDeybHMI5NKyywiduqn25spJ1SOJBfPgTaRCTiWlYg9/YtUl
Wx4bTmnh1vh8+7nWdG06SINIRhj+pULBZ4zKi9f13bAMCe+MVJHyY2in66u8eY0+o1J6OD3G1mNi
pimyphEiiQ2o/6xaJnCh8mp6dfjS04RhAdW8q4kzvk6O7ZabE6PGuIArvRT6C8iYeL0QZVIWhehD
vXkFeEod890rcbZMjqYxopfR0T6fLkXyMi2FSnSk/O3966Wd9oILDMFIajd+veufvuyD2ocBVP0i
oR6IbxzFf4qFC6eqOqkHDf64Ihok1OobnYlziOdve4md8fnO9nIiUgLnQLHwytLXZoReVcxTWvFJ
LNPjUCaxYmBbVadEY2z3D0bVi0UqHycCUFP6UWkaI8Hb2GZha0SE6R63h8nK1ZcBioy3TvrUJv8b
OmS+Tqv7rsZ+Fmqce05q+BiEAD2QrzRYhFufXiEkxke1pe4EgYBF8pVnfzVRQd27ipO+XlSZscQv
/xqZNR9oRz4RWnPXFe0NpGx4O3iOfUEp8waKKbqoFFxAYZakMXeJ4zDrwW0wsr2igcB3EYZPPWIc
AqC/K0hpoYDRoYOrmYkWeMw+I4mYQrOGHNxg+8ecx2DCzCmclhgEfu1z+Qu2jeu3MBp/3NVso5sd
zQJW9Y/FrANM7o3oLEe8UGBmEaY9Cf6OYGotK6P8X/H9bSjz/SEksKTYNKjbjyTvE98+F25+xbOq
FIbvg7f71tHIfynZED1FetwZPNqVg2HuDKEOTthlOyohXxNjzK5DSi8vnB7+ZzqiE/IbSL/TNz4u
bd6M9OXGCeGK/rul6J4O29aBg2toWYxJjfCXF76VAWkzsju/xNTIJGiOLFaM4uRGU+lA/wWrT44p
n64KNGNl25NN2q3QeuJEuf7cPdIzGeerClfLTaGK3UD24R/gWtr1sr/hGBOlYt2c35uNGxV8zEBV
XTR48LAyoHgGCq15zwjDriy02ZGgsFBwCjeZnuZEfYKlryOVMcVYsMnTzDP6maZ6q7WqC8sBynRi
P5bsNM2Q/LF8iHk3jnwKz8HnVzuXN3qwsA7e4YCyOyMeny6G6LXog9JvJ0zq3cY6ctdiM0iO1n0L
9wp69J+oJcM+iVx4jXG4Bm7k9F4rQxuAsSZbikcG5rYJ1IpsXQxSKKIYEoZu5imq/1YOcDF/kG0u
2nFfrYS4RFv3wdU8JCK7RMkv/tXSN3dpT0ftQwx2J6yIL25GMGhMv4axnXVUgGlU0ArYh1CPs6y5
nltLmFq1kwujyKpEXqddfdMtTy+jMuoofZl4Y+84NdnK5LN4OiDIUYPghEFXqbH0XsBQyl2JR7PH
sPtMn7sxX8bZ/vbo/3d+IBkaEz/TwJCw+mp+pa9A27TWGrILIYL1EHWxmPkrAx9rWKLtawH6e1Rj
kIhlg1cCKQaq3SP/NB/J9e4P5h2d6K2y3XS9PoHBAXL0+/Gmw2S86uDyo8oJ+rlVnnfNz7v+nAkf
EEaRr4QYQsRXPVfqKiu5sV2y8mp8XQtjZ2RXfhHI267KdXz7AIuUKeWFiTkbfCLgclUOScaR1un6
v2nSitIWa+bpmny9OehXcxhQC7XClMoa+4+o/PpvOnZy62Faelf9JTRnO9qGXQ0UMmSULoNt4Mf6
unNA6/7wP1QGvZlo1wf4NnSXZJzVHb3YUfSsqPebf7PmfvUeYDPv4NPzy5Q2B3+pgaKPAIheyOP3
732p8QC8rTMj0i+YGe2+zOgqfo5vWDIy0OO84biqPC83KSH9oFH9n9kvMzMDItAU4v2A+kJgEp32
gKf5hMEmF3Yv1uc4uflRO8Q+YP1lbSWkKrywm3bgM9Sv1WGHHkUHybhNGyi6fny9MwBHcfO3My5c
undhEY6ntXrwJhkqAJhVMYg8YMFH+dL7lAur031uGOB2tbj1wr2Cm/cVDOepg3c1M5gNwfkxP6AO
crtVie1O+dWUDXEOkILWf+ZJKx9yCIHRBooThCkxi5LUzQyyKzGS3ByxIzxoUUCJj/gIsE4SnUNd
aN79PdgkpXFIjUW6IpImwgz18LwRg4ON1Rf6b7/lUyspMP+iKje1hmFyKGCup8f2Pi5/T6YyKzHp
o/SXBCcEUBRHvQQ4+M3SEEhokIEgc7k+FSUvlg2/zn2oIA6q7H5/kV8X0Mg/wbmlhi8e32J+pffS
hdFRdlMB0QW7YDaXAqPbWGlk3FcNqWJEUR0RDg/3cbtW6FLP7ZcnY5qrlCNHeh1fZOUIu49Bsc08
b0ycTy42kuZaSRJD8y1iXzmqtBZyYD3XroQw+wVZnTOZuRtB5C18BMfNyvtbPildr/rjf+N2BlOx
Lvz1Gq8Zqys6m/Ld8PtgVWm2flzrljcHtz5MbMICkDmjqiwZYxzee+iuYypdVK/Okdj0meXAxPuF
8vuR2DRXx2vBdY47vAVp//awpNpR8KPAXjDbe4mDyVYTb9PGSM03HyYOHy3JzlxK9NAA9W+qSVcr
YLNDB/wDTE2puP91TSWRW8xwYFmamMqjaKgdPN1aTPvCylQ1krKc3c6hbD9ikvuTuIg4sEC4l5Y/
9MiBkkmO+ZI4YJD3yNOMTQs43gTz4Jiz+zbphhvoZfAuCZbo3h5yywdNI618uWbl6qYqPSmwGKUZ
h5BiWYifjcpZ78Q95F2/EoezQQ2j3v5dJ2FQ3vDDVGZtEDo99lvhrLv/0llOMUK1h5Ftw57+/EYa
3YljAJOTlctACGIo2ZJGft9mLPr24y7gMkgU6KosclnpYLoyWnyla5i2b3U2RtErxfd35kC/V5ZN
kcYwf3baDC5ay1P1wCnLF+RiibgEBhBSmHt6inWtAedJd0eE+hTx6m0MmHgLC9yGy8cNmBqp3FCG
oWNXiZW9wtAeItj0uncEC/Yv2FDZ4I3skbODkTZPsZR2VxUmtcr1TbDWUVXAvFObePVe8orAO7JG
yeJuLBi3pZ2Gz++EMRZrFPks6l9QdrKzWCzxUXUgEjef0b8OhQjYbjOIIWx/AueAu5TDGXX5Ygfq
2sCX6TtdMGrwednOr7Uy6D6YrC4beRZSD8EyD15RRJ+lAIdbK1aH8e3qXw256VbHAmH0wpLU5d1i
N/Xeec+ZDi+Ne5x7LOLbi2LZd8SxuWSaoqFvHKBA8G6ec8TyU4KJPR9iphLq3qDWyzf1X8ma/0mZ
2DBgRI74Wiv/8iZbcdz1eik42RVZUd70yk3S4HMezoscbtFAB5CZGRom18g+LDoIscGS4Qz51cle
J9Vhq94Mdt3pACBlNzJX+xo5J9lHVXOUV3PsJTs+Y3zjMKFMaiSTXqsSnjPGlJgVUGzajow19ySB
nsnlW7gQcugIZepunZH/6HHaqYj7HIfVzeA2rPOoNdcV+IkzxqK1QV7eZiD1aPTOzulmIrTJ5Uzz
KLF/TW2dMB6tYvZD60QXMu7dTcGO7Xqc5EH3e1AGtL6tKNNvGqN/FqRW+yGB8A+xIc/qszWDWGvi
K+Q0KCNnCJzHM/HN6Nn8T2d0vu0j5vxkcGtMy10UQwbr+iE80EBtlB66fkZoD2QKySqc1w6wZhCK
TniSEoMV3+S5x9raz/GdmzorG8iqm+WNYLz7ypB7tmZwZxtt9sEDaBp3PMvg4bs/ReC3pVEq3qMO
VjZhwuNWttYyJclh6M+ncq+KkDbS+8o5iAWJnVmyQOufaJzprgfGRRt8Ff5OELh8mwqP9ljo8Kg/
Hn0UncMvoVmwmMdvzxpQpWNfUYwhfn3IgYPzmwNQhW3jHPOADUfRJqfzombAP+LzgWMpveQ3rWbU
NhGetHPw+Ckg5eftB4ZWpr8c+MhjF3ohjm6huxl86vAoYmw4R5Go6MA0O8sXc2UUHeSRDGQa1UPh
jyrx6oPBWG8aAtxG4q4IscmUV/cz4W6jD1/ai5an2EPleoL4rT8pp0sOP0pnyiqghedE1qq7eWY/
lYRTG6HTKZMHm/gPPN9cBS2vxdZxCY40zDEMXEwQxvAOobcWGvD1GWgFua/kUpt+j4TSfmQUzJot
nTM6MNUeLMOs1m4+9VuMVW9p2VHaqyZ7ZT61mjRC2q3xVDHbFEoxw0JwIy+4RUU/ld/aDZer3zYM
M5lZGbBEYZiEvcDO1mwAwRbPBrgkmtyU0R9Kb1KeRfnezt3zH7ykRsFF361RTmGZ86Ocekda6wjc
Z3vniNeJjurFRKiqybh3lJKx/6ME2K5QDhESCpG/WiGC1fiQrZNfJnmiXy0JKkur7sExNEpZA7f1
xbl1xqGiMJvXwM6u4JNXUQQrRlsylflVD3LnSuYK9A4EtoomB/Asr+6/9OFzIgXBo1iHurUBlwpG
u5M3b/cM5sNHxqxARMXt/TfdgT58a2rjzJfNDWoBeRRfcMwd7+RS5OA7KoBscOkOAvV+lgYf9N3f
GmEoz6+Zwp+iCX0HrNoQoUgR8AzQ/ZZBcVPv+9XLGN5Y+Ghp1TuVbDc+O0o6edz6fFhrrOdLGWMk
hrNUQkvizj/AheYevOyijcpks3tS98pwWzC1cJudgdvWWKn5tBBtd9mlRk9aYzu1tAZSIQMpBNRU
tn7AoGwh2njtmVUtepdv6gzW0hm0P8k+nlu4LZQWn6YER7EdJVPQsjPLxQrr+aaIA3duBEKsGTu7
x8ts/m0O7H9TYjc42EPZuJpObqju3U4BYWVTEc/uq8rDR1QeskdwcEwvEJQQC7dtZBry3x6kchLU
XGH+43B+rvxU9aDjv7lEe2dV4kQ85nvIxZws843+GGOXx2G0+54kaD4+kNkHELihXQrm0tycgv7p
FZe4hlq2tZ6VN4D9WuPAr2tjW0ICLlOGWyqFJBT+2EOXUgY3SqkzoIAbueuvB2JpYBU8UZIsnWr5
v/uMwnUks49jn7SOSXupq9Ddt4rtRgN+/5YEbHipLbPn8JZq9BG936Z6s4FzORrnYJ1bBplUAwvy
vqSPgvx4lc1Hf9NPeLl4yYkizUuf6wPUdqk0xxQNJisL6D7IWUem4xO3Gf/GGNr2e5uX58LZDqyb
xQx26QEiNsd4NgK0ZrMEEuhlmBCFHSQjahGFTz+LaerWHapaFIV1Am6Hpy7RQJvC1F3VD3XHhpWL
yqV8Dl9GEfeZ7FDvrcHrSIaYlLeN+UTebIC42lbyESIlp0UGaVxLRkD/2EIAQLKY8GFRx5vDDSi1
80qaFVBXiMgKPrZdoh4QuT9dHPf9Wlxq55ImTctXNoFnIPyYcVuKmBfSCqHCRWuc6+iz+YNwUiFE
f7o9gDPkwaj/PO0SoRzGjj3UJ6DSx1SmXukuPWfL5jrtd8fzWEytbuRG/F0mZk2mmxOjZTR9H0u8
VZbeZphAR6EaVSOsUOJTwGbilFGhICcwoWAs8t1hI36l8AxubViA/uV8ezrpycrIbrNrLcsm9g3N
ovb0cvK4Ya8H6lWOMZ+qdVeesi/76Wyu/UTc1YgO3UtIovA6CANu8aEerM+UPuip4f3bP63ZFNGs
VNN+FnyPexrR8zEHKSQeb+mfh36dnrBJr+cF3fsUCTRIeGNbeot9lUy43eSeZpAGsH8Wbw/jLDPd
TfY62siz63vCCAYMRJE6Dc6Xmj6UmhfbpIA47LkPbVxe0HGeKfEIgqfshK+n3tnlVt8LyrsGespD
D4qSUc1lFzbusmZEG1NqtjrY5fOrCmdMOahRXu2xuhjUKPg60UdgTBAfKwzB2g1NKE3kgkntCdcL
17Jjw22LAkFz9ExodO5VPSVV/uLo+21yN7cHxc3xoZ2UEhq+PXHd18wsM7GLby5nQeNkR6akU/R/
16YmNuu20Jqnf97KBdNsbnn48JKl5sVNvaH+cwgS0Sgex+71tevxSaEJb9C9FMIHQS6NTAweZcEC
uxck7oYZ7q3Lt6TY1hiJOsKSvl5G4N219GKkQZsKFGzhIe+M+fUwwyC+fwv2YHo5sv8p9ERXNf9d
JDq6IYUfES2FSEhwjQzRmkBfG9pXv6/hp33VGzrFSS47a7YlRtWTuhE9elRoGADOZAel18NpEHC4
K27AcQwj3MgwoGQCYCIhXZgmBHgKhCaDbcP4InJP7lPts5c4ggDDmQohQ3h776BGY6AOMD8vpKcU
PNMPN4eSz99KExjUxTq7UzezBroHfknOqUhJY03HA8g44SELZ9QAVTOQ27CAm/IdRmcB4V95csJS
T/e0b9yi1+V7cqSxrr6xl63FKt7zlNBojyS6LqVJK8jj47PgflF8pLVVdS1nthTm0Xu4EQkdTn5z
As/2ExadWMeuKsK3KT2OZavSpHeRD5hiGyDcfdaCihU9T2BCX3R1OZbvotUrPxzVRWx2bM2PdMem
xZ4UBJi3o8/4boGOKsacD2hen1MdZ7cMOB8LFwQWHj9j4VRwaHQjGESRsq+wu3/LoZMkJY/aG+/3
yhbNtepRBYBvQlaX6MeSms4pGJS8Yks5MJ0kT+Lf+QxHAB36IRrYkjjpkOSJQk031ixYxwuo+pdS
U9W0sg2Brn9lIQBoU2djN6E3jHXyznOpb2LzxVQ5dNkOLannDD2wUNy8LnPXSKJwkAqNtKuGoLG6
3KGSVEOTd5Cz2B2UU8tCgX6HRAsKVHkasD4/4Ssss9u4aV1IwsvU3MT0aLWrXWaFFFuoc2PrElUv
vexV6sZdixS7CWbCqNLRAwWr6+gfcNR0y2AvqKBFGeFVo2ruMQcNGpmPCFWJX4hMmL/UeJDaCDW3
x3df19yQgxnPhkQx0RNIEC9mr7KlcDQGQaHzsxzu4v5ZrtW5LXG2MEwt3+0YkPxpzoPQA8Qf8NZs
EaNzerpqcuC93Prnk5WN3fRsY+VqLKxQHNyd2YpCvmBjd/Rzzhg07RMcF51OKgwgV5sPbY0iBuW5
vIMNXPy2HtYkb4SASUA1+CP97pnkaINFKx77W7+ZxwyRzVlb2OlSWg1yFuRG33J/KdvjeQRXURQ/
o1kMC0Ogw1XSV/+lBlL6Wpif7ZYR88iuW8jpCORPHgCHfgQRkYGF94XhsBnexAQERu1C+QHiXZv7
UsgFLfMMItkdPgcOMuXuruTWB0ztFqdMTz8Z6zO6IwlXmDqv67SjZkmk/LgjZMwcw809gG9ooH03
ovspypz+EfQc5oQBELRCrYCOn+xooOgT3aiNdPJgAgXubpg6Z3bxkNHt+2bMH0JDYTho4k9Nsk+L
GfxmyORuxLFYH+FOaAD3lWg5fCtriR1iwImlSDKjE6ZUiYd/VI2H46e0fhp2JSo7Nlo7/rWvo08i
qZIhhZsEBTcMFiVYymYg5IzK8DSJfGU9EIdtkgP0uHBMBEaHsjWIzT7rFdbvzfHcI7jHlKNtcOZv
2D/wqVM7fqEhTNRDndakq2iQ4Psv9dm+C2hcBDoEKr6GhyIYavLQCBrAoTuNxeCmgl1/Lji2VbHB
cuZAvy+NBs/ZTz0OBSN4QLq4SazsV8vX1e0SQ8kHc5zSAKSIDU1S/oFvuxPr2rc1ugzTzjKoCzRq
WuZ05sopJC2lciBARKL9okcTqOEIfyHKTHDtEwpRgdRMbf5a1n/Ncp9BzOv1nbOd+A5tPZutvkYB
tdal7q2mwYvu9bLKeR9yK+G+pdxCuOpnRdGg32OVMKBbvXmYBocpWPxHkomtx7L/XklLWyVpLbyd
boA9qO3zQpH1qbXO420Hhezm32LGVXdRaqaIxqXyDU3O51st3DCDcTaqpYKPjKr5O/2wNbvbl4T3
1NGR/0v06KElzZ8NmBRoxROycXPJajjQYFMRrcfmbiWxiAssBfMh486Ba/+cRY1RZLevzFTIr8ZI
tUX7hRqJKX/tggMZBVUpTWPDrYmVpLahrF3OhYZn7hdkoRuY+jbcPZSJLjPB8YSOGT2lKJ8ts9/h
VquDHgjWpcDnIPctFIp7BHvSm/lRfDjh44cInW0gSTcY5Y7JwvBPBdF0IlaYwRIV1f5+AgPkS14V
bPSFEbuhdlcAI6/cqhLKUOoDMWr+41ZfMjm821ce7HgXcEFBjR/kp4IvONDyLc0rxl/HM+38DaDw
vsC4GWQZV7lzE0j8kWgZKRRKBvuNPeRVkQxpQ4O4kF7KxX0SiVvRnu2sKNAcdc9crfZ2Z/VmiPiT
Nb/JGyRiIoSmSWv+sXqfs0VVsoIhxKH8aW4xBX+qRnnN/WwmsF7Hdtni5PdURJzqpuYqF4l/18f2
eOwcXL9OS5pEGdyDbURexZhhk26r+ZE2Aw474J5UOkAGRnbTPZv3EIqg+DlG4hRCTfiOOz9P0U25
5kSlwDv3lo2KeHLOkO0x2Xum+nsM/FHM0OHJVfAJvPiVCASedGgZiD6gP9D+8kiZ3ja6AgJ3ujcz
33kLcY1A/RQQGcopbyLkym0cS1nZPAxxasGjtAzbTI6Z1FXhgltGSCevgWbito84eCm8hATxAoRU
kezVRMpSVeVWh1BY8q0stD7EgnLM5en7CiYWA+RNzHCJw6ZHeIubF5VjmwukgtkTZX6P6SOn7k7g
kyZlzzH41tn/4WmoNwn+wytRF0WQJ7di3dxqRkS/iqT0PPnHZYpH1NVp0/CyqhjwrRg7x1h9zph6
fYGLLyNNKKY+FyjJsNfP/3K2xD3JweSW1sualhwRx8hcslDoPZVnvVnyPRzLxZeXz9GlF7Dtlel6
NO71GUyxNYDpxxHwCGViqOgOG7jrmM2m6xol7vaIABMF7zZZsqQbN71y1LA6fI3tAiIRg1YEgYyx
d9z1PYT13Lk12ShDqZO+hZfsJWRemX1dHcTWKcJFSKluk7vzjhTgi86EnINBbiY/Kpz1da0ew9HS
VVk10hQH9Gu7d0Xx4YakDBVNdt5kIT5cxFnVKVPc/ozOnzjDtCGam7wIlOubekm0IRwhlSNOFZE3
1DBNtmKt1Ei/iXOLfwg/YdpOBW/O7ljy3EZhDaMdau7iNL96Zl6YRl+esIVWZiwQHW1gxKBcTNn9
aSeKvgK8MjY6m450bd6+/hZRbUCVciuMr9nLHhYjA31RJPJNT8UOoqqOAVFcv28gI2+45Q9TC51L
ETmZGXdR9a3SsdEsI2NUU2mO5JufSs7QxHGOHRz25WTM3zFVH3792WYNud31VGb5dEaAoM2CcIcl
cDHhowX9ibfkuwclrIq8yPiUscqnLCuLMzDall/bzCFiqjlev77pvKLzWCaAU7Y8dCkEVIF1swml
SnEcE4onU9WPD1Ai3DUBgNR0/byhOCzNRCBVxaQc1Abc3GACe9/XsaWtgN/XZxi74/S3qpTDqAsr
xkwYduBy5Tl3lbPTjnxWlpK+A+187hxD/hdYsEhD6UCHLBmA+hOhhz3YUV0fJipRV41f7MNxWs3L
KLKPLxABVyigUajhElyoEQ6By4tp5PBqyPSputicNuu/NKbdqmlMsBlBLijL4kN/Scki8obTyYOL
M01ApdrurHy50ri5Q056a03+JitVzpa0i9MJli6wyysK8tNpXxlh4jQz4cNKmXSF34BK3NBQWd9I
IRC/GHkvwPZo5xzYexKw61F8dbMisAweYvfM+bumEtKFb53F+WpXBffB256wJfShP204KqqGJ4QG
3c6vjWr877f9ynpF9ZhDqftctoHEH8e1Osb4Ie61+XRY+OnlpiCDjG5C1GfZYFasGXS+82HI+WSc
hDkp0+JZFZ3ZMRj+oHsng0WSZSq2ZVcNVdCKeFtkfyydY0E30vNplohaDzQh0+7L0uwW6OHCxxRo
PK62FPFimXoOjyPHIvRS+xsbjMhPlHhWtaaZLeVz5/CxYrC0VZ4fz/4iPdvqAkqFABvd9nQ+//AE
3int47L/IMxdo3YY5Neb2LBkHsZV6HBusMpgcccuET/vE6GoIcd18gQ5KAOlK+cbG4s63i6CPdTE
7htgisfibTvAlK3RF+Ugo203wAnexMWFhJVKHxIDKMExgqKyQf2jyYvTpNeceoo/fOvS9VGoV19S
2eJ1L5VDmNLB6U+samB5xijSJwHvfpTjndZDPIYvGu//rO+vqlYYeAEhRJ4sOuNNh6T0Haicybo4
DLBPX3Imhx+sOgx7IVwxzhUFX1Fovx4YX5E7fTEjw/HTxu4KLfIY++jNN9sjqyi5/sT/W2KYgDrh
t5eaMospCoE4ji3NHzx2z1lZLy744RpjmaIqAvWH1B3yCVMbUHIRXeh/UKnj7rqaTENAagnBvWsp
CFezC2rHfkpYODs58bi7RaENvCZ3ds3cfb4av80CQI0JYzjCSeeXWaigkrI9iqgVNrKBKuCaDMr6
NfqnOr7nXNdwioD1UKmvflBiAqB+B009dGTykRbERzNbPKRMAkLdEwQe/HUeHwO4owR/cXgzs0SD
FUPMnA4wmq0zKYB3WNgkYmbN+Yksg0ILDmq1VfkCs0JwqrgYma7K10kuH1IaLv/BlZaAg+Y/IqzL
nsLPzrEM1idRL3Olw7R8KWDVdswwmWo/FXKxcQfU2Yxm/CMT3JCF7W27fASwsXQjncPuWszXydT7
vPSN77YJGdz+ADK+8L5YyCQ7RovnKnDh1EbmVqiSyhYoggGsa6RradfacG/p6t/+/0GOYR2twk2G
PbhIJGIkUh7r8tZtuP8HWKnHn8ZewUttEIVwBxJXrTA64ubjnQ3evqc0FerMtprfnNwgielR3LQr
oiEflhxHbQZR2p1JLvokWnoTTcgilKmIX+zn+rWBGjLPMkEIQ93qq55n1/iKOGHzS9ABSl/CKlL2
rQSZM4fASNaJ38Wck2PfznVbFq8EgPWyMddwgpRSqbEjHSoWgm4fX0ba2ElanB77kMlx4SSh9M9B
+3NlieRexf1EL7+hO4luB+gElhk3DdCk2H+u/MvKL4sARq9ZHsSjgTgHiqX6IgOAiXz1TSnSEikP
PZJ6lNtVKxAMKtgHw05HSxsO7fcPMf9dK2GB5gXiijERb9s4Nbs3jaYbkKZmhOFZcPNVJVPWIVeu
GqHCn7+IWkWfDvetxi5d3aKBrJ40QZXQD/t3jjCqkn90PQye80r2rQIPl9mrsu8Wb5BCZChlgVXJ
lCezVjykON7CvFWV9+FChoP3lTZLLQ99aAA+O/+raT79UJhDTE736gPj9aJas4Fn1CzyJu5PP/3T
ntvcQJIqfWpBx2GEOcCoFkAaDoq9uCrxZqsNSBHwjKPysM+ijP/ewNYZ6wLArcCXjHF1hP+ThKAI
j0vMg0W3/R8lzkcJZgWMxeK4QiFaWM9U0Q7y+7pA/iBVbxdXvtGg4YAmOdd6z245eeh6WY7Aw/Ce
CuM/KlUwvslefi0Y+ksn/0c/FnDCiPmzdP0NXPcmIXYFhSqPRUcsTghrX9vqQIdhlfbfsPxcAkqE
Qq6IeP8ZNffsNfXxIUCP25yPPXUwWxHE8BqPckRL06oevukcK5XrDZoK3SOdlmymLGI1yx3CGsMN
lhMm/TlZe6K4VSssPkuuOMDL6ANhCfe+3DPZENwv1J0sZjAQcNlHrlkYpzn58krkQu9ZKj3Rxrc8
losCKrCWGpfLq6jrntNibpU+GOIzBRGQLBLcItcQcuNaSbZFghg259Ql1b/n30Jfa3iLW9TB5bsz
8a6UAymjf1VQX7o1I3dofYJvRwa4EEyaUkQ39uc3ohjsA0FcBnTg/PpBH6DjA8RPWecOSdr8af8v
5O6IG6GRStjZcFhEvauvao6n9FbFW7SXOgpmWcvVoUJ/r7nhBZcOQdpMq81p4ApfIvgUGEH6qSds
nuZRk9vg2jhnTzXV0BhKXSA9ElV9fp7pi7JUDgmoYeqr6d+qGxKA5arH8MWrRFuAMw0sTtLDiMdS
26yhqJ3Ab1wAQq+tVzceqbqHq6Tb5UVNE7+GRMYv5yGJumwfBrAvLbDTz/DZw2oV83PZV+p8Tq13
OAXzV56f27nzrzK2yrdzx2G1c1AOQ+9O1QeOTXz+6clzCIzyCwu/7fuKH8dAkMAMQ4aXdOgSyDte
XK9F5514a43icVn2z29BNc4yM7ZtR/x+Z+nKH+kfgY1ElQxK0HB9Odd6Lxq9z/9k1SX1YZWG2IUr
buTV5iVS2nN4ydgi6wziPYViIzZlsTa4eGbCia72eev2wLbEO6N+JyHHPvN/wFT5gaK3RW6Nmlas
nhZj4YSWZ+BRXhL0fIHjkL72ELxvP+kiFO93pKRgFeGFqVd0vnNsXIiSZuA72rpbp4hgmmYEG4Z9
S63kNIiyUAq1MdZy70Vri2dJU3EWP49ZommXYu0V6lya3KWU0BqBA0gdYF7hkFCATfF8XVMBcqIT
7r02gMDxYnyDjGywNMoP1D49VlL6B95H5AqQHAwzsYQNJ6Xk1DQZ7olnebn1TSFkqXtBx5wHr6yt
diRTeEHumZtgqYFynxcosHxy296kdyuWCLo5IazHz8kSrXSShHROJnUOJq0nDLYMlXTzOUdw3gBg
HXGyYzdAPySWFbxRS0J/FSbBDjiBScKNMRrrLR2jBqCK2q9rskUIeLGMza4NYEswx82/UHKNHCqw
FE8ZtA5xqhhQFIsiii8XraoSDJFk46kcXBaozP+0Ev8PbUYrhDmMkVbICMPmYS6tfr3TTnAGlaxL
En1giw8Giq4d9/Q5uMAFpjGt4kFc+fuSrvgA/5dH3J7hcGSn3h6A7X25Q6sSkT4LbOdMBOcMyGji
7veyjA6Z2tm19L0vTH5DI1D6b1NJLo+g2LCggteLZMdjLxsi7fYhSmyBhp/3zv+Bq63hKoKoSpYt
HoWH66cBiJlvpvCOccA8m7hUgF2DaMDn0LsLdJaQI+tx8YNLy6aT+gR4EXZKP1YPuKTITx53vSk3
yVPjL86OVaM4xBZdTb7MeH5idPuj4/cWCDMlTX86iQLl9CnSRbE255CBUo1dIt786xNxRvA19f2U
GTwMwAxyWk/Fir2Z1bg4wIaIYa0/RT3EmNrGNVOyuarurjE5lWYolMujGH4UIkpZ8NQbgns34HmQ
/1vewwSQQv4+CNwnBcdRvFMdG3XZ+lU0hKE1QwpPACEGALnRQs/96HpxmlkYmgeyYEcPC9e8J5DW
M0usy3av55SaQCedh9CS9aFSwEcb97HxQWVchafu6uZ9ksMnr7OfAu8Y9W3cS77FhrktliqIEdji
LRN5sLdlHyyicmPmURf+lqfOd+FLWuKQDbcNSMvQLNupVVn2E0psb6jfPVp8c4rN5QNt8WdJ4+CG
yp/nAXyi6hFL0eVUlG0ARECr9YVQpWeTwj6QcyBQzM0uREM78pXOwjZJz71xLiGeaJZOkIcefXOA
cqemUhpk4vtao0d7do2yMMUWKnOFuhsKdPdxGUCOcixFcKjH6ho4heSeDZ6x2zxL4rwcYz+zgSAE
ooBfyHMsIQnsYSBdcqA/LnRCzGLpVyBvJjBHxS/zDuQKMt9RgDQSZUueCQSd4K8GACKRc9h/j6lP
QhKKeR9hWKyJ+ev6SaATqMKjaLleBN7yJ+vxRArYceRvSgWu0ekzIMYYFawJaYQVqBwmkPZbvxvt
jJi/qCoChkWS0hzKJctdKIb6UX1fpF+bFsIel7pdlViintsHBO+SLBYLVnsSlElnhQ8fY0OkDRxF
2FSf2Tc2UXZ9gcEexp1Q8YwXUu55EcRYGeyXDU3XhYrYWj/XHqksrxnEoAcjKs/W+Nql/1G7v4VV
qzpMcSRJ4u4T6KoTpxDq1WkloKI+eeXt5ycTWhqoNs7kFZFXkggjEWfgWAs6FiCxW2x6QChe8zPc
F4ZNnr4yTQlrG6+n3IJvtgJYzdcYCzSehhUh0M7M+0h/H0ajm0fdIM/F4JmjqBJq+FPLhlWT3qOL
hKeG7yovbsttJo6O9RLD6ip1W91x9trjoN//xFDXscpJgen5X1yWsgA4ARis1G3toq7gWsoQjDq5
dsekYYzu2y5n+gFtqw4jnhMBduHWg1SMbA4hBuy18koShFpSQnIdVRVp1S9Tw+NAzs01TuOiRaTo
Y3/FnuiH+KSlZS5c37EgKHFr5OzhipibDiI2Sz5meLj7p8wofZ7M8/9RLS99WVkG/bgR5DHuEVur
Upa79q/7dWE7AniuoOWaMQmtNeGnFbUCX3CkYk2ulMRUjF2+cH1HqU6rs+ganqiSg4RrDsvujaAC
Vypha8RfBMrOdFUjwStQJCJOFUnlCnFroD1UKwlxmhLpSaaeQrigfTQnI9Lln/sTW3v7t1xmXEYU
ZrmLfwargkP24xGDRx/DGnN8pKN8lC4FBiPH6gFSMAtEi5iabsHpiMlfrErG7Bcm4XtiVsKVmEOH
6y+VnEgmKq4WpemgloRDVA0Pr6K+Kc1CqQ/atGytf1IuUFQMznZK1fn0lCMU2jWolscxkbJIUeG0
5RQkTZ/qqxDtaQjJe29FOHCcV+gix56P6trsZ9oBlC06bXM4mg+vKWQdDkMuu5pLfmdv8kYE1Os1
ujUUAdDVANlUXYoMRRJuUo/bsBpn+25ta1NkdflWj5F66NilJurVkP5KLKYQ2YENPF7K8mk/XTbF
lhtvpRxJtwKEzIztaUWg4RqUDrw0Z9aLyHS+KgR7941qf078QXGygcEY2cLpHY8z3vhMasmDA61/
QpHWVtlee/0ad/eIMC536vSRxmkipMy59EAJXJ6On7mfNbcFEDdqfhy6zpog13t7NtY0vYVXbwRV
CA0/+bthwu4igSie1FSB7VCahlldbSq1r+kLm40f2lR6yB6SEfAkU5ozSQ6T2UriAUWWoG//yMqu
eYnYs2kH19YJ0QOk7z3L6gI3HASW+LR0J0fYSUJO+NJT6Os0ed/59Nw/3Mottg+ixdz6J8NjT6Se
1XyEsRxT+JyWSRl/0hbkLgrnNIdnHmqfuYQQ3Qw8cQf20QCi1rGU0LE2NcXM6p9yyCbvXqYI8lYW
J+AbY/WfF6X2ODQ8mA5Vxn0BrTJrNOhyZzX12gE6UBip//Z5tDznSCcWiGDOsjB0lrFFohd1+EGn
+L1Ikv6w0Mc9hqCOukWQieZYMsTqeh7kTPw7EnFekrdm6L8n7XyiJSBL93QWPCSLiYrhbjQsPRD7
un3prfkWBmhlRNkL3lR2ZLc5LW4PlccXJHLVtB3et5yYXtEuDlz4b4nDMn0Pxvcr3AlHQfvvmRXd
YDob0KHJQ59jce8buEVAgH+r43Y02rZYfPNs/GIgRcop4QFdeDXitqXymuMGSfVKpc1s8cOvlNm7
ouHS51+UBgYgXSDIUJ85yXKr0nq2caYLfttUzOvu1A+8G2kETnGJ+1Czh2pmAFgc7C3kCZG2xKxv
chycJSnDMtHybJIZ47mkGRUB+bQrvf5btdp3Vkx+AyL+PIKnjafW6uAUv5q06C7s9CsMGlPYgx4o
YrdnQqUjE6K/pY+zQGzGwia4hhhfZMfOuMIaYQIYnAKlHYcmWGeEWVqvzw8p9FpFgpmWLpqE7t66
Tkm5Gvp9LDHZMFrrn5DcqxbD5HAiEYt5KS/ET2qgNLX9iAyy+KvoC0IhvbjykvngbKDxp93LB7rv
ooqc6mHPyv6bsHsvnHFhMZDD4bxdbKEglfHZhDFMIFnmGOCwCKYXbRv/VbNHuxoLZCZWOXzKpYvY
0Dwv0g7/y/uiJf1trbkDVTCnIC2U0wdYv/tQtvxuRehQWDiYjfakkTgMKjDSIDYRK/JXxhTu4Ykp
Rmmzvdvcch70p6bjKJ+LaiciM4Gt0+/ZYxxJhhZD/kvQA1Ab6IqVzClu+jO8SZiOVZb98QHEy4qy
7rDJNCmyuJTPa0MLFCLq215lY0pHL+QWTZJdQ8oDUWIdur4dUjDaditiLCRR0vTqmsAsRoOtK8PW
Ie2cTaHnCXZ07b7w8RPj+PM1qrTV09rAqWDySqIB2TAh+Glaee3LnvUI4CdaegwzCprE4C9gdO6I
34lP2iYFS4SCJDLHwF33qP6puMAh03t6T7gLhSDXYC4e+8mXLLnQf1HP6EPUYshcWS3SmBQcryvM
q3u3ifaHIEaAewSmvoLJmifO6x+1YOIbww4GuOT9DHekF41YMfKrPLesFvZMg7KBkOOUYa352oLT
TLqxprbhwoO4o4s44bPiqFW3m38XUK5idfQshyj/gbDqUgfai64YbV7JzjN1iGEfATU78RmC2gfs
2DfR7zLq0ZVzW+Dzzcfg/y6VGPSq32A0qE4ZP6Rr39DiRakrlMS1F6tDWko1S/TFUu3jUzIIANVZ
t/zp/yLTfIRVrLeK8IIzDtCSZ1Wj209M2k6VOu/kmVx0k3TAZhvDjMlzfKEpgGpiYLaOoBW7l9fs
50wgoqEF2SNg610yuU8DjR0AHLyO3siFQWsHMUw7Wn+EXef7J/NEN9aKPnksBLTDe9LnyLXbp4gd
d67L8KeUw1X4kqF+NUxecH6VO3OGQentz7+C1MlWaaM3B0fWEaFoBnk+pZ/Ae/nFNW3ClR+odN5r
FL+sSZXU2Uf/QTGI9ySxQiFBTZMf+Ue1bTK9Nh5RmYqwBFnj4ae+PNodptCsxhuo3rWOy4BPWEP5
9cJQQr2kyAVH95rSqzIcWt7/WsSH2EZCpdLpJeA8YBVe7RnqR3E0x9urMqxAtXdNtUVOL0RFKooo
/ecDt7lAKTb/EVkEaMB+7cvLw072d97y+vCifsZdT7qZupqn6FYMaRPqQkPuFtrEKGHabwc1xFlm
IHFreC9r7nTVxO/9JUuvNGwt1dTOxbVIhM5Q6iTi+iQ0kJsuNf+ccGzcq75C/uHPZQ2DyB3s77KF
/Oxzdce1tuTyY8XHl1e3Wi9OvUkZw+0BPbQkqM9eGDUctGc9VAfdWH93lCDEE/UVhF8qB9yExjAI
lllxW2iGxGO2kedOD0ijnXn2X0kc3TBFQpTqObcbLwCXjjT7RYrrc32H0vPafjHvhW2x0JUxUFiE
MbpGh+eL0TcGi1uHNboh/2rRZTDMd2NhHfWQZ/I7hLDTzqw7W/ZIppWeJLvs3bEeMKKEwrdDCwtN
/It4dTm1IUPjKoq4uHEVlnmMVYX/nD2Y8qBvnzr1Ix2kiB97coye5lXBPitFJf50eZu4LI/8UCmg
f8dvDk09vCIruXaOzB7uH3pXv/64MuNTcRwQDFJFFeXNPJjBkF9c6bBMAbzwKUFKgbao+3rGpcFV
kYebTOTU8EbRNwmukVNqb4ehTWQMq+eznJCvACmUjcLF6MN4dn6aYfnXbdvUo5dYmqbouxFEf/ir
FjrKnqziRAryyXrttDRShmxgEXYdkZtv3eZ/I8YJ7GB/9/DHec+1OcHmWWzo6/HaO9nf4V5yKyAg
uncDRX93AqeFsGTlsPH9dn8VTCyt1Gtr5hKo9KZmuIRbTdR4+jWlvY+dfEmRsqgpBDjUw409tzFH
su8COyU1n3Tn7mWzqFf2zN/+57MaG2nJey5jLP1nrXLOuTFOU8DVuxWvKG+VqelFIl96F8xiGKlP
VBiUfoEWpLlzio6GzyEU6zf3+ZWLdc8Yx7ViJs/LYrsf0xud830g06VSI3O3G+xdU4MiZCT69D+I
i1bBMakingfZYdtIhv/iyfYWWPFki+usRFEXAf+4jFrWPeYT4pJE6lQzeQIbUm5vWrZO5r3hwsgi
FjaF7dJ55d07JgYmuB91gMPTAIpAuPl3Rz/Lr2iIoCqRUrt4h5863oAAyn86XTyy7EAcamExqpgi
4UXXDiBalKx9fo1lfw2hcn8QQU8uSgtmvP+Jo0+MQdATzKDz6Z5uwcs6BYgdEWSkgVWqLZofc2za
4LJZZswlaZFvyiZfdza7vART5iLpGc5YmcD8MI866Vk0TIopJnDSqb5QeBTNAODOyNbOjsJl+Gbl
mpiJ1UGoivx81AM14/9m01SMEzfPXCbZtrkE0zD0xMwsZDT4or0uzzHqv34BY29ftNwXfFeHtR44
VjIxGxFTFr7I1VSucwCCOezgVAr++rLjtw/J2G7+whDli+iHqefPFYARaJYCubjaV6KxP9RVTrlX
cJZM9zxsZBzhgXt/wsCVszFtt+9YuD0ScTcyP8Cu+z1KkHNnZyM44EBr6xlAk2tQgJD79TatT0BH
leXgm+Jx+QYNzgSKpBD9OPA/AMAmrMzHK37CLYZZ3z+TpUw23yYnQ+OoSES+qF99n2QjLOjpqlJS
IXZjgN9g4BYdCcBFtsZSA9Ljo/80kwLvNmIzg9Rp+n2B5USD8tkLFfnPIzNWcCIdC+8UyMxsIfae
5L6prPZixPrkOpE+8DDAbh0XGuZ4nbm7XRn1GDAlwoOIglGUEwG+CF83u4Lu0A+iXa9cHFo9nDSP
TLfBfj6zYBF3l5HeLUniTo485ijOEIdOH7Y9Kwhzo5mP0DMot8CuPEHD/F7XX3pYeowxocLIeLUR
nL6JsEs6TA3v+G2igg3KUw8SLRU+RmHr9ImUhrBItQeNreCosQagmxC5P+dmgW//DNQPOuFxFgTI
GXY5CqRNR38sUbEpJy83T1+AeVCdB+qpBFtL/GsDxSQhl98zHkW1Gd6m9j8O/jLianReRSCevvwg
paDRDSL7R/NTPt+Ac4cSbZ47O4KmvB98rnMB0yz+iHs0u+Ri2aQyFRSj+IHnO4PHQ6ZUAM+bac8K
tMuKsvjyajWrM7pRSSThjGoYXz791eZOrFTJgI6S91tD/lukwaVBwhdVgUejrPnuyZLyYUzhPPJ/
Uc25LBKEaPz38kFctxB0XAU0fSWd3D3iX4x35QVNZ6gWHWkW2iCD4PAATEPnKAl8RCLqDjXVL5Bn
TFnKh896hmZQznvCnBVVfq1KrCSKTMoOL1r2shTCUf7Rg4Oa7GVNmAjiweN8B5r542mMWSeJsXZX
OLYSm6cGa79WROkuBgJf5yqykbJKEjCDZjeibajctY00X1XKA/WaeTLDyOy1RuGu1VKCKwQQW5sf
va18dxaP7UO7ACOW7LLT83pP+T3OBkePPuKceGsbxrz9edrRJ98Yi6mU9oEDiPDkehYI5uFDSHiL
AbEM6DEv12lkzBqGeSjlPtxN4zXymMU365kTim8ATx6/93U8dde5edbsSnPW7sv6XcUTSQLv0Znz
2ZuoD2u2Da1RbeBp6lySOrP8bDc+4QqhDWxgMBDh7Z/VzvsnVJYCZdrbobC0dUNwFLL5NIvbCpym
EVezS+ObJIlnIVyvaY9sVmRg2TfVceuWw0GDQfcnB3aBWGIPMDguez9X8pnu23oj51YtECwWBBbb
maUinvrD+VqD3no2oY7XtFXP2sGM1xY+Zs2+1ATKHlKo7wYvfaPuyIuPXlJGmKRCw9CFrFHvUvoO
nOpjtHTDHlT447Oh9VJN4rGLUPAnWj/UwdjpU6in9ffrY82pZxznQHfNS3WM5f/wwvDvuddVb9da
bCRi7UE+R11G8WjQDZwUVBdoCS5wHiadXss1MywzEZWZlZWfxijptj5jrxLQ6HpuCzWRTYtXY0jA
V/NGPcQmrHj4ptc5QtVsheC9QwZ03Tj+pvX+WeTeyHVPOVA+TW0hYPceINhfEZrtuLvPcLbg7RMZ
EPHari78Npe43L2JNJmo3YlcUxB2WX18aADtJJW0wq31iAwAKR1ZWKo/9kU52IcM8yC6gbH7+PZR
T+mXiR6GC+O/l4bLLSrKpJATLR7qjRPq48MPq7TANPhy0AEIrW9YcPBx3aZGfujcIiQrwLDk8kjZ
EWAnBHK4h/5puzMZlukK1BjYxFpzbl5RL6lb3fJExr/zWRoOLF1XcyDdYwewRIT2OXN/s4QHm1Xj
9kWM7ugsGmxPfLPCH8OHJaU1kp/xCNPm2XDZ3ZAoCAy/TBdYSzYz2moN339W0lQmZ+j182m75HyG
KLPxv4kCg2y+4ENVMY16u5fk6KkTpaTYxz6ZqY/LA0VuJfI63+3OXbrCCYFryAZcMCf6mhQvtpGE
dEcpyB7CGcayG1BwIIC1V0pVCuaGRyL/mFyF2ZLNTO8Rk6XGLbwMLPlkkP6JKEncOouM6dKEaC1g
acoJu14vBdZ0DGMqd75ZJfqTEqsGUVJXfp4h9MtAYpYG7fxfiC2OB3KsaNpk4PyJt073hnyp6w30
X8om6ljcECVpf8yqLJJs4v1+6kAZhtd+v5OneeMkg02ZwAGAiDtIsrx6oLVd2j6MMuoXbRtpgu5y
31A1WXy3cMKmeeBggYybskT6KFSeiathXXXEU0F5M4nOYTjjus20aDJoGZ1GhzMCAVgN4pQKhLt/
d6E8w7Z5LjpPsshQRK2EE/EXKZLXZVwqJOIaKu7KK7auGW/rLPdIm/rUVyWSNmMGWvYz13z7KwJa
dhkHex6u06s4iTzCRJT+S4hC+OnnTT1baGKvuy0Rzs3X7U7foJV8LExfS1YxHT89ksax2CnVcrIb
tneg1nAMGLyYxLYUplae4V0wfjkad0Z7uXq9gkLWu80OXcJVmly7VvkNYerbY7HQheBXxkpzNmpx
YQck+DOQUnKHFfertKpeIvxdpOfPkwTN3b7EyD1wCjzwKrTkinATjx3VcQmgbjoGOV8Xt3weeHxE
A72njUMoWjU9DPZUQmP4AaoJ2QrlT+pIVjJTFTZKS7VAdVt8MDYFywFqZEIYSoNsY5HL8TpxRwuV
biRVl7DIISyAoYuLEtq8dPx+WWdc9jcZ+YCOK3DLguiWhkXX6ZCaO8QUyTdRMNSkaFvvxdcQUXar
YqiqPA/jUQ7XuHWNpoLv7+99lhq39vDNIkl7YECTpGr15ZTsSgrP7OCxQGT0C3cMYXL9QmcEEO+Q
aQIy68Vr1sHJfdP86cfH49RhyM6qHtkdLZa9VL2V/mFt0lvVIF0lA8h4AMeWElGplpfN4+MIejpL
eJheOgFrTom0d00nG7LhAcZj4oqNlLj+FrCYSBDC+HrlG60BNaua0V67pFmbmZeRr7TUuVyHuRsz
2rt2xMPa6sLA1QHfmZu7LhQNi0o5xV87RSslRdqICPvTs8pvf7gTrRIkeVSYqGxBZuFigaqKppHf
7KimiyGBqPlJNrFxPTNTQ1BmTEUZz96Nnzp2riJI2V/yvtVjxha4wNbCiAzbfy4G56Y6rHmrFYd1
mjUFbLVsAEs4I0kicLYdueuwgOgZ4ipTlKikMox69Zb97ALLGplT9NnVibM41juQdT9dHp0NY91M
q9AWwwIwD+nC/wDdm5kSISySFowjSPCOexhxn+FZqCB2vAwfsNuqe+jgyUkJolDo0315RAruDCMG
sMlhUVARAFBFOO4QvvsYCr/tTD3O/OCtg0dvwj0aus5++SKnxWYrRHegDG6dP6w/pqx0dtoS7TVv
iF+FYQG2tFVH39sXzDLQvAOc3+CwNxFGNLT76q2GeKEYnGOw/GGuhzuz+EzUm2gCq7TvY8bk+Vvj
KBOiCRPECFBkZdJuni16wLLm77RSlM3X8Bp5JRk2Q/rDL1Zc2IhsyTE0SdGw3Zv2ETbz5auZlSje
VQ20Dod0ZELgysALdSWd+dd9rDtEXYzldhezRr7UmrNy/8aOvGVQN19LffBbvpRniPnGraPelVnc
dL9l6U+S+PfUTfyeyoTGcZz8utDqxjA+vIx+wA3y0EpMXDp4cOoJBJ/vfdKiURMn3RxXPxTd0TLa
R/VDLc0CpwpReYrZualo1eWj4qmzVQAi5m4YwkggH/Xb+YU6jvxFx3G9bAtBcRk2Ewa18E8frzfB
HNr/BEdFR0GnzHYXRCrz+Q0qxa1w/lFKOlXHNdYTXyfu2subeQvuj2HnQnsUYCi9rCWsWtO20ipK
tTNpX196beui0HDF9CgkfLqQOfmadfrBawqXv+FFL2uVzEMmhng6aHhNsHFCmqxMuwXrolgCLt71
QUW6LMrrk6K8lFSzvcj/bMjhANZLHC4sMUgzgdvzNDaVLxroDAG64mCSsI4iBr8xtQeZUFmfZ8d9
S0vlsbauxwBnZxVboseXVRakUkb9meTHt1zhXIhqwssld2mcy8MLIyUVFFYfYEdPzo1+37GxDWp5
g7PbVdZcz7DiTVH7VWFjt7TvB5nlYuCsgEm9lqhQgzNA92AwYZ0inqOKCXpf2DSgrG+sumdr28k5
u0iLn7cG5LaOZ+hWrzi6/vxRqI5yncSmPo3e57+htp+mZv+/Gq0w1a4KV+I5MGJ4WotlKhisPtF9
ZZW2/5M0I4rFlfQAxzS0hvqnUxmrtPaqHlli8YJIw6ngJVnXgVofrJ0IH54vwtWrCiyceDGBsF9j
y9aFW8dqm1RunXo5mYQWutLH3J2yHuVDRVDPuonuqGKLaGm+vKbrFtW4Um/Em7Zb4dGJdA5Bg5mT
pUeL3jKxKaIyD1G+HHRUFRrx5vq9opK6qyPEBRaaPZEyjIjSakZE+cl6rp+CoyO8Xf+Gy03TmFhu
Mzdsd9NDghYd6XJSIseZbbVUwVyG4Z45oCFm/M8tAQU8O06Ghm62RLEvQZqZH+4TtcwzD3Tvnp18
2zbI9W6sUmWMrA5SUdRgCzbSvMFSSFM5BQ/i2OscmwSn7ifuVKUDrVgmMREBDr9Zx8kSyzEP1+l2
14MvzUJVZPhhRJgAcQ68UXd02McglGNDQ4YQbFyBVlnIlCUwZDxNyIdc/aAG5DaLWbwz/T6yQ5d2
Ep5HcNC4V+BgLKDnGp/95Aesk4B7z16OU0g/ZDUFdeTaQFymIPVQqIloezLT6o1ZEO3aiEQ5dlXN
8rLzVbp6sjNrlMUYNJmH9PWTcPtSTnPoaXrGWFVPm6PonsNAffAyJIQdIk5da0XA3awXRGmPo/Fl
uaaQBGI/02e/jT3kfJhPOxTU09doZX8nZTk6lR27O94gSKQTJCi7Y4UN7XkflV7NuUN3PfOysdXX
PZ19KALhLMgYy5u5X+WmaVz2Z6iDCULWx0kmrpg54jIkE4I10oHoRitUO+woLG2VVEyV7g6xZpxU
F//UYPl2v4Q/wMWT9igGO6JGyvt8+iZiWr/8CyNxKy4+QQlaDQxgpmtMFlqWCReRoBLSsPCug7i8
Uh795Mk00ijSFKrF7d2a6xZwGKrOmSn0nsdVDp/XfmYkAyCwai7oePRjPLjpjqnrjvJytQMonilj
eoPJAzPRYUbW2fcqBh9dEO7dt+VlXiRxRaHqSj2IvIVUNYEjgdC2LKbc0Zc8gW/R453EmCZaDG+k
xLDMFf9DFA0QFy/HYRNxjUTH0W4dLXit+4Y1C57xOGO6macnqYbUKPRUpyLZ7c2v+LQQCkTq02pf
qb7MeYjcPZwfDoxow4TPy1fTJQyjmyTBVw6UfPxH086A4hFgNJFlzqVpNV7CjsJKj2O/mXyeiBOa
g6sQjTZTKwRSK2Idb+R+sdoZuOeJRgn2ijO84CC+pVacpsxnqFiYwyz5C4oeMx8ANfzKrNugXjsc
ZODJBeoJzdVMkuGvdRFZ9pxQnQpDXGdAc+N4BDOzuYMQlHnFDNz20SQ3iz1xqLD6CdiuIi2lRrR3
K6E5er2Tap57BTJ/VDEdri1Ko7M1TFHriJXi+R5Oel6P81dmhly+WJbHlMoetnaIIEdhnZhb17g6
NQYHMr7dxcQTEryZnGi5lC/PHDS2/8J7CoPgtTgUdl9uOyk46btgH8BIlRiCIX3qvqandEPexF0+
ZUYsHJksGxk62brjGQYqA+yyvIjf+1woLgxa2jx6OqXs3lOJGGbOauoxc+Ld2oX+wH52raIZFftl
VjjAB6mtbH550QJUo5yQlRLzw8pCdCHjHS3jBuiyhGnxxjUgpCkTOCKXy0jwl5vLq0ev+PvT4qBm
2ToYZPZO7ayP2tAtiwy9NRfpL1VvPSLjQIPJZxHGyVPxq6Sp+baZHxgwfz3vPlJTU3bJgMQm3/rz
ugNAxWpc8DJ8X7uKTGjRezw53lVJSyRIErVwQkqEsb6EDvMo2G4WHwJnqEUhVgtoryPoJhiYOQTd
DP+GV86QOUWoNXD0p+qi/1mOtaFu04KMNeXIy35Eyh1RwdOCCIXr5K+Vn+bUneb5azd4p257E5ZQ
MbdsTH2Cw5wSst3Nf1zbqMk3HpOnzzAynlGGrILbNgoE4NymKdxLbxLI2EflN01rKslnjwpMMwHo
4kNCQE7QM21LqsR0YnMIgs/tsDeOmdDyJ2zqEfc/TfRUq/q/qprRapir3vFbUW9J3K/GXQUuQnoG
Sw4EePjFC3YwmLWram9Pex2IFm/hgLZ+XNuGbihuHZh44Y68Gz7eBWGRNCu3CTPFg/TdXOPC8Ayg
NH6C9ozX2KljSKShO7cl8eqZJd3CKXOn49J45h3zzDy33VypUpZkLL2OQwODoVGLVRobeiOLo3Yc
KHUj4Opt+EqhhR7HfjXpQIQ06TF/pGUvAMxRiTN05lyEBPt7OT9KUkeXEBkS20v0YQt8orsDtKub
DUkSEMgW7r1lKtRfn6l0lp87twaN3m9VXR/XfLgCerO1tqgJvxWksfiMgs9+YEY+4hfb/u7KyV7T
RE9BBhKYPgUIq9gBJLKdU9PWzL4VRib0XhSNfs0aCCQkjXNEYjtf9RVkjpYcvjLJo/e/QramZgqK
7lRp7lxX9yRqWKxELkPv5VaLbFwJiA6RPnZWjDpa5QkVcuDn6Y+sulOeL7YShtAB9GOoNKI0SxUh
zQdrPl9TePg8BNpATfTAjTUkw6iLVmS0w0L9qN9aX9GIiFmRH7taikV0oBP5Syf8PVbDqKafuwAO
fa2seIEglJ29lpQ7JHokNYTuDlcLuHIYwrbL+dRY40VIeWWr4asDWFK3v1upN1CYY5IDk+QAR4vL
2QsVeRlkC8doKYZc9ZeNOD5mQqlUI+ia+lX54oMg2faZVd4dPoT+RxkAqtpRhkZ3yW4d8i/vxOLx
8KBA7X30cuIwo47FfI94T3P3zTLgTrPjlxCE8LxPHZlXZ4Te5dBmn2oRuqXM+bKJ4BXsipu/qvSa
UuC8/FkajYgDVC5nr0am1NtOr9FBnhqj2dRziZNPzfA/IywfVkDo9qqCqxM0mbWd2Hs5mna2UKUA
TMiSWkze6cjbRrVsZuSSDcL0hYAfYiXKxTEE6r3vI5v5kZ6p2e7FIDlyySTO2UIpni6YMDtDLnSW
WRQG6ljWte2xBxYa30FBrYt1IPeoEs3NjVVLFODBUknhVk0GRjA0h/Sa/+tQlxNJH0kI9a8yPMEy
VsTEVoliigXSQBF2l5oRgpEFnfySE9x1Vu6U5viegs9slnf4/VyUUeCujZQeJzPlbH9fgqqy+4pk
cbp+QVFKcKakeD2FUkww/fUlI0hsPbPi9vZi9XZmb0b9ZPcY4a7ZBhvNyhf3D8OI6Gpiuq4DDBri
9aA6YKstS2lKI9vkOMefaDqIU7IWMdh12eHxmbE5hJlOxKMav/yCF/wjqvAwXKm/2+YyWs7Jvv+H
d/0q2VIk4E0V1x9uOGlYxlTGwLUQpJFxp7sO/BfWUwnHX5igCkeEN/pgOSFzaQ+o4VIZZZ7dbiWo
6jNIcU4Iy1//XHAP+iXejCzwYvivrdMnWxnbDvjItkFWLwdV4Y/UpzbAcuOvzDPMl6Vk8ZXvi0vC
XM3Ypyw2XaXQtO3mvwjhVSb6cnK6e7fWIPHEauEBrYw60BMezhd4KR44dpk0iF3ZGDwaI18k91L1
nKIWN1s0U2J5QwM3ctGoE9GIuq+EsH5+Uf0sMbG4tMvqCG5bqR58mxvOAFfc9k5gvCRAbvS1MfYw
60Si/SeJYJUSdie/yGBvYe4iTWP5zimcoSmB9QggQkOmXoCiHELmFhFA4mDPkL8pAKx99P4JoV1T
b4lNE1I26a2WVpsZGpTCwC7eNyewrqJNaIQaYcueUQJcRS4AGXuiU4cjFyko3VP5+HLayhJwSvz9
RA0yVt/99nGCtlu8HSTh1KKpzH/WkAwkRmFvgkP3lLstJe9Y+QBezpRGlev9imFldC9PuGGwvD7w
3VYaZAbtHFqkModQjIuYWiSxoOnr5FX6peM0prp8uJbXo/bUU9GfsVvxDgy2Eow/xLIcLbpZ7/+2
mvIo+wz80z8DiYxwJl1u+EIZ5631BKRQK44kuAKZqEw2tmOjuq2RWwBgTlgq75lXtQL/H3LsP3eX
IhiJ6aPegELOZOkwucM2TYwq2SlzZgcH84sNOR1vXrOIYv1GgCkfXhK1f41PO7bRdbHUQ6iXX2rq
zSG1a/A0NBS0TXnrm2BQe+VNEkEn2wWn4jU8tdg3sYb/dRPKmuBiUgkbLaLWPnyb9lJYBiRAO+7P
nX4qGJ9gTMj8ERkmvafXEPtRy3SvnQh1rOrSDzVuYD80OsEkvEI0ehJqETq+NBenCggonfj+lPqo
lUHphXNhql7r4A4Ws32bz+9fP1HeYPHZKnDOJn9xBDq9WcKUH6CCe0f1cPt+1GEETHke31TzeXw5
rvd6FnHxDKJ4g3sFdv/mnAFVffwQLX3pP00H51PcNlFYVxam3ftuUe+KM4awcsaL1CeDxlki3WJ9
34Zv+GHyiYZryKAOUy8TJyxlYzU5RdyFHd2u2BRzAlV3HkmkGmBZt9ViKsFvzIu2sJ3J1gl7G9/f
CM/IJZJcAX0SR8Jg2V/Xtk8jRmd8K7Yz4s8Oq24UdzcJ1vYiqN6qqDs+afFZRGklESAjYoOAYwlO
/rvt7pfOxDoA1p8hcts1veYC+b99haxRcs/k0UXQB5ss6s7ywbW7mmprE9JJHwlbFAsHnBRLWA1p
8TU1UcrXquidNsoKeqpokZwvpwz2WLz1CAMuZB3koLeWz2McIyi6nxUAIAZo1XPZ0zyfJi3C0pzY
N1BOTru+ZAWW00wddNY7Y87ZKDMF0Imk3TWKpMyk2h0+a8rFRWa7Iy5ULIg/CGySyFXr5nhcqiqn
QL8kE8rx9+CJUXzNuj/nI2Hdk5o55MQVx9vPVVZooV9hdMhdvE2AEmU36o53O+e1eGU0kLRjDFTU
8R72d2jIYGC4bL9VQqnOgbLKkzTF9EkI03n+ehyaymlbthcUFDzCXdRDUx7jKdlB5dBmplWdnhYw
N7jjWhRVHRbUHdy9qHW1fSssAT/SzCIQqKvRia3nONQ9WxIJZxsSoFz/Jjhaq4y0oS6DC/ustavv
sZKLo1FJxi6R8VzjfqPcSbAKr5TZN8op2HTv9HD7HUcVsaSAVokcq0LEhF1hsni26FPAO5B738g0
kx9kWLHns4rVzN35Qux0xa/R5/leQFuJciiYRMg0+Ep1aVyng7MbawPhTC0S07UQprx9aqxO+GCn
6sWe5mHl6NjJz0lAakI5qTJ8iDeN0IVlepRLHE66V4hRJQAMQLBttIIcdirkMfnAUiHXAhau4jJX
9RaFhEzV+qoiPG7/UTJ3zU6fTGSkpGs6Sk0Up3Crpv1HttYq3W2EjT7BtchRjGLYr44I7h8q317B
TdH/Fl9fDTDMukTXvld8Hh6xs8afHR3r9cJqaolvRjp3gXFtUTVB9uMNZK1KZ93VMFuCCPnxgmQZ
NPzvbVcCVrEzYTQjys6xoDk5RfxetOBUFcX1Q2Ih7xx0mB6VoJgDj8JLM7drgSsCQcvc++ViVccL
IV5TVBBsag5EBLFdbD+eaEssvItkQAvDpavKPpxEk8FH+zEqKcCSraQhnfOybQKFefcArPMj2qUC
Ktn3tRpum+yWuDPr/YLNUQlxx2I7l7jzGMAtCX2lTMx6B5O+XXq6uwzITySHlVOzQ2O781kFNGUi
iaw6lMnH69+QU2ZqO1HbB4Bwq8/ahpYg4rL1RjT2Vt0dBcXyh4dJqtw6MVeHHhVHA/tTGNciUynL
1YSMDuvPkgK9at2tCgYKNDOJD9nHlYG+e50wE+K+gXJcbF7C8AxACtoof7JnNXBhL6hkFi179ReM
/joYUEC8H0Qebtdmfvi0SAcbcoqgsvqNIyCeWyoHdYNyEG3Axkf8/ace7ZylJeCrZ5HNSQPpWRmt
MfLzMhZpJNOyrlDI5+X3CbZj7hL7jBbS3QbcFvH9oKI9D2G1UFEiphiYr0/m0QzU8rccelU9kxHX
zyezhQ/QEr+2k/R6ft98q8zbFm8I+Nqgm9PfQpgl4n4+JNVtzJufs80JN4zT6436ozhvHgi2xibT
3LLY3GDmrhml+PpEvvHMJqP0HieF7wVmFi2OEbufFOoXFx6yu1R4GklgWnI8utLZwFMid+oM5NtV
JpFuCtvtxQzT2dla/WeKm7OHD/I4rD4uAX5J7PLOJ2CtMiKSPS2hhDSKn8lam+uac6nWrcAaDZN6
xg7xu0JEa26vk2dljYPtXV3KIGD9AbXFBvjInHbsfU7oRxLwInEC+gUi4nEDX5wKTGqOLzywYIHh
tDKExhW0v3Nb+cDyR66uJbu5KYYzxuRJDaa15tuVM0H/mfsGdldzGsP6MdQ4tcu/YobCAPOsKzQc
AILqo8zOggLfeMVJYbWc8cs9QOFvYFJWd5CRk8pQcFI98G6v2nqstTVKPBiyRLGqVt7466UOMGT5
zyBQQUFoDEeAMHgMPsEr6BosFYbpHLu0x31MguPiUkdaovB/7B3b8DKl+BGaMMdn2APzmjbVPDbe
IUDouGsMQbJLEcLdidv/sHqQRCa/Sc4BeSAC++BkMYNK/nGyGz7FvxPjVG6GJIDBHRx1769dq3lp
jrTpbsAsmwB1GW//1zvI7U62+4bX1HbhQf9yJSFJTH+bOE7heVKzJ/gkOFvzALN093OrDzHshCoi
UApJFTzoyZEr4qIxHIG0Zaq4cUkhxz6Z/pHrahuJO7D8QSmnYqv27zBT4tMPTaceJmQ53tSKbJ9t
4LwBzCqovYK6Wvg12mk3rICbiIrncHLjxV72j48H7Ysq6BJQlWavInlybDzFEmyBQS0r31IlpZju
551TP5k/AnrB/gpaPYJoDxdhaI8FYmuM+BH/XtIa3HxMfzoZtjI9yt+dVcBb/zRgJLzPLNwvtY/A
caknfWVqW4mVdTdmQ6oQFfCOpmFcDA8JW1OxlMXZlr0h2yCp2VnLoviQXrkMbsE/LVoy7sGnIOPD
2jPBsL1lFGH0on2Inm2xyw7hoKwtlMndveWAyIuqPRQ8AxxXkmjyl8GhWzB81S2PGY+VAcJoYwI4
lw4RMG4quUxJOUKOvdFvYeglVjICFzbEYabh3WxwmERKhj+AqW7bEcwFb7U3ooMeigRBnOMHDOHg
BSe+EZF8cG2h3CV3zy9PUImxwHc+bBmxCQBREVE4w046nPxNpDJFQWK99aP7qyDL46aTgIlb7YUM
yCkkvvV88ioVtB9lGoqWCXbsYtsV8O9ypyeEGo7PwO6gGZRrH8hHQ4hk7SOERDUr1vTIxtSr4pwv
3nb1JM5qH7UV2YL+Qyr3VtsEaBBN46aKNFEc2M0RhV/HtB/xWf3rk5/sHMYe0+7w3ytXPbi/r3Pb
7UcFUvYx/v2S1G0F5dWgb6knRI1enxyuwYKoOcla1xShHHh5kJ0SbWLLt4pocR98Pftl0wrBc4RD
z0Bdxm8pC/wBIZfV/fSFCCHy2PKJAvQYgFHTYcfbWpk9FDpJXvbiGo1WdP4YspopTJuK5WWjluQs
2JM45FG53WKAoWx+8ciCcoivnE/SA1hnxi8bVB1bENRnFBvUWPD0DCU9j2c33eYbGHVFtFz6NiFD
YkZlykiEHiFgWWQ887ZY/TSHT/NJubLEPcjRbidS/Je6LBi0oO5OwvKFIISryNTQv1yppIO9ZQyG
ZPoldF0DGr9BmoIUFxNhzd52ImyuSIp3zm/uUQUeKvtJne4/4yGiJR/Sf0K4Jc852iX51mqEOjCD
CI1g7bInI/Q7RZppKDTWWWQr9VcHbYbuQ4mTQWFFzWwp2DabaxsrguCjGultNw/El6JklwXYaSG6
hmTl5UBvZivtadqm6e5Q1krgIiv0oprtqori54u9GH8NeNnDvx/73iusPK3jf8+p5rYqjXUp27qB
8SYqEOOrK9Tw53lkhBIF+NUl40CuJxE74NJkiKWSewWJ20NwMbQvLOOr7uIboSGxCxz+uv+RjLr8
aQU3WfzSf9R+ZeCg/UNtWOEjUJFYY17rOY34pcaqQmKJ+ATXmN9ea2sQjYV/ahBMKOiPfIooAByq
x7iDCN8NIJgFWBAZ7ohvKhsm8sRZjWbnCqciNrqYXr/DDTp6bG04xB/xL4vY78f7t9coNFBNMrb+
4sPv5eb990qzEZwiu66EaCQyIzTHYw014lppIZWa60yzJ/d7loP36Y8KBUz0bbxMIk0Az5vJAyFk
2Wvff6kvvcquC3/2DOBiyrcQpH1rewgX9xbXF9B0gfNP4KhmEWrCFVjIaXHYENJIWG04GO/iHW2k
tUpp6zMEjNaw962PMMKYqxinaPcjgQWrtuQeoM1o8gI/+ZSJoIzP9iy0PMD4iD5WxBNH8paURrwT
e/oFc50RihBmrOhTfiHHg5yfCA4H42F0y3QfcUa249Y8eKw4SPBzkBnLBEy8g95FOfYNZrrXibrQ
e8d9/p/LIfgok9meYoNqdN7dAlWnnk7FNI/getry0tfrZ7U2Tz0sDIl/ioiZI9rFNJKcZUv+Kpjm
PbfxFAj2PhB4qGa2aaPugBhPlGvpceTXhyuE7VsrVDBH9iC2QXQCfwMy9j2+w9OwQ8EHB/Ko4h8N
6CgRX0YrFrWAIgxKU0fBsOtRPGNRxXkdQiyb8A3cmzkPjyCnXRBMi2/r+fE7AuLdcbJUxIGiyfZr
nVm4I93ogGd9eYFsHnsZoZE9/Dh1088AOVV5dJljebfQO6USBCpFcKAgv9NAL6JpDRIcTYHg9CFi
SgCS/tiRA5wYD/lNc/l0eNN+6cDa+vGfCin1OkfraZ9YNYFzO/K1ZIyPy2GdmDS5vnr1PVfoQz0Y
kjju75w0/sb5W5u4eNZ8LzyiW9TE1zmaRv+L2XohHKWjKMT14hZvyHHWiyQqkhr1TzLAAP84R8Wv
eTsaXwzZPnWl7Zm8oTr45YZS1Vbca9dgogt4vnbYKfeN3G1YqTWcP8URYwvCEcgkummad/HsHD6Q
hjNDbR9c7yPQfVFXONE4fOGfdSQSWBsCaUncUF4eqt0JbBVzbM7bVeXjH9zL2e128NkAfTVhtbKV
FR6nmhc2xaxRYZ/U10o0e/q3hkiGzQtEqf5QJvploa2pG6CFC4gO7qMfPkUxDK6MPNLk0RamBi2l
mJgE5WR1KGPfwH57YkLZFPltUFPaEsEstE+dujxGL6FehTY7qXB/ktPcdQba18vQSG7BlaZF7KIo
XFO3ucO3liLSjWNL46WfnCv+V3tG4VIY9zrITHn8CckXVcIXLOUyBDT62aShxzFluhOnc36qie8e
HyzexK7xbFOocN+C8bGhufrvS3qikLX8bTrpoGX76MlFCyUn2pzffmH2xu0jjo2ukfyoc5Lx5yo5
ga+zeH7M8ErOsdOEpmEtpOdfOxI9xZYRkbO9/I4KdwgA6g4d+Xi9WYHzamRHK1SfEup31KnMoM/O
N0Zm2H3TOx1GoTo9pL28iYMNRfrKCAKXxKqzcyJf6C2W8H/q6PmqSVothjRet6IUrvjdT01wmuw3
qBl9IsYiYUgD3Jyx+OcvrKCYyXUBx0wjCD8ZMTP8pGbcG3Zp8EA2aWPn3klO/dI+ThQNklIHFLQp
c0rrE5yvERn9uWgLDxO9Tn3ViJryJeQDbdqNp2Ab8uOSMNLHLMP8XQO6CsDfUEfEZ7Q4zz4NYIIf
JeFS3iQjHTBU5N1RdhQl4t2GsAYYqDiH3+19M7CZzO3zH8Ar2WJdF7cKr1v4C2pdmpOibojq2t90
ztL03onlXVHnyWQDtLOURR5PJfPU95+pxeO0uIlvVhJDu8wOoZMVonq6oG0nu0BFVKRgW4WptnRg
l4elCStxRUm7bQgizr6fNcvYN20qYe7t4H6KZE6Vx5BEF1onUlLDf5PftpyeHVPR6THcYNIwgeMb
gO3qtuAF1eDbdCtSaReleVmm/1bxpbJeR6KhIZU0+55Dr6TS+VANiRdWeNgLvWQslAVIKwXN+AHc
KH00PLbFWq9jPMhWsNXt9WQV6AhDxWhryfNQ5evWktmP4y0fk+pW2DrmbVvxU8galM3cCvYjnCWn
3pUTUtqM8bKTUCaDfRRll+1npGodjYdOAzMWmTwkIEv25axtqCZdjaQmt5WE7XUpwHdKxYaqPnWc
LOquO0mN4W7ZiTuPiZYoTcN+Pb9t+g4ftUSFrPeGoDzKA7FSg4cx+q+/Nsmm5+9/tGRNYfEYnUqS
Bqenu4Al0viPDw3q2unXf7kHz8ni5b2hII3At+OMDPsgQTEpl8aPc+Rk97L/rJnKEeB03bpUmk3j
rnoJJMjfq4ojZKLAeo78ptbZG5Agbp2Ytw/M7WTDWHtPWP0PGdp0tjqm6d/HUGIk6FSQt3LmQTss
4jJoTwkK7EnQoj5Ic8A+bNbu1e04OUFJ9Q/mqxgTKQyqXVKviDe41/uRRuhb0jzl30Jdm9mHrGDT
L4b2Setw6uDJKlfNsYLdEoFY4JT8f99C9ObmXrISgHSbUil7OmVNbqSshuIJ26i3GbAoJzPasVZV
Db9E73cyG0s31yWk14K5Clj4e2rDeQ/yHjjyG8tlppERS/plVsCvxTKQ/5vfGWXpTWD+bA4YXhQr
XHXuo9Fa64NcOjEQWjL2pQ3QtfYRoFZjm8BFERcMH6eS0FQ+STx4uCEHRIgbUajJlvDrRFZl/23K
6yzt6f4ooAcUZClTXXhuWiRpnUi/lzplEb8ehyV0OlldKb0XeEJfANtF+csuGu3lGlHEZ1bDXRVH
MtBywS50AFsj5icfB97BBy6DO/YvXkfzrVrkWi0Le8T7s2LRHFCC3xWY/L2QoEQ6S2z6jtrNRXQl
/vBPYkAWVyeAI0XmdnSjX+0JH0BdgaDq7sQoaniE2Yz1dpj6mx7NgVbYMThycXjLh/O3B5ccISoW
oyyUfXwLLCrElWEUZOIVpx9vEuZy49Yj+LTo9o9mRK0qvxyW+pjx0UwWTaiiGXk63iD6CvExi4Mb
mig2T525nJa+2eihM+ORa9A1QESi6hj5mKF/wjIs2V1i6xsRecs5/NX0OKbgB3PrjWhOSzqM9rri
dP4/lncvtxHHrqJsSK8ZBzWpJw4t8FkJwy3OkipnO9GOozm/2r1FvP8M5MEE2cqtfFfjbZp+u1D+
n7VXIiIqpzvL+hPuFRD9Pw9TeIMAclyaeNUtrtJXCaV7NLG+NtPZWCP6NDtDBV+U1sc0NMLhau4T
09CIVaGb3J4Zl3JcML6H2jG35qr5bK881uv3sjSiUGVbvZMZmtbayhj7aqmpgNhvg5/x5zUImP5o
cjV/d+g4MSy8Mbi0tKdMe3cH88UZ9l3v3/uX9noYgoYmJ/R1MTqJI7UK6rwE5avQ6a227eOKBsc3
eeiwMpm4twnQHjwdWZwIfHsRBhdVn+rWw/pDT+iBqvDH0CgXYApiy5Ak9gLgJHAHmieb/7EcBYMG
lKvDb2xu5wA/4bASgxkXpe8cEEyrZUwSJBuETM43GaQY77qJ/XCwB6j0WDajkxiCAw/pa4MUFm42
q0+yYBScCgtzdbbdVfacy80WII6L8d3V6YXRKAT8z3XqeJspwuDIx9u9Yu2vmwk9c00DaGiK6Abz
GmdJUkGfxynKLmc4FQuHnlzO2zmbllpmQ5PvOFRJLzEyXoNsoIOs6vanyySK4uzzS9soQ6+mvwqj
RQR8aGn7eR2sZv2im9e4XY0b+FJbfKVFZMRNSaScTZHBwISNaWbWICWD25Aw+tYyZ2UmZg5Nk+2s
fTVB95G2v0ITM5C1TgixbOxA/4v1q8f8x9oRfr4es/NHwPh1ciyoTY9IjQEF6S7i6lGLSMEuYMJT
0YxXGhwFux9DlKgEKTrvijTn1ZCl8hzjA+0r17GCxKq21/IXB/LUl2ToDnZA59nWg1wi87CviKmK
3JqPYM5TYMVMoTjNMuoMG1WiQWNeIFPprvz5MUNIrm5WoyC2nKHKXZN027f2vsYrlxV4YUmsOJAk
8yN4e0Xd+TIeoJEcSazuT1AELQ2w6EPIAC3JmWcenVorw1PL/Y3nqOpHgABIsN8uORhAEOFzPePO
vgnpr4mwOSnwWHrUZn/ZpZpL+OETQhQX0W3n8vpc8u01hoYmtpp5PkSxs85ttz/TRSEwuDwGFIDB
mywK/NyEP8ozlvS8B/suRuGHB/XyUkuTSPIHJPTwbbCeyX+7llADOcf0MvOYtHbWhjBfqBVsgzwa
S+IKBnLOJMN9An8OdgM2EH9xPeUE5bADxOdpFXa4ipJXeFRD2XjASFUTAnyZ252d3tgViRbsY6YZ
jQox7WzK9nncVctoLnUj7EO4M9NwpFXv1T0f2CfaeMLGLqukEWwfJRtYVnQkGAtBKvohTlHhfwfX
RknhUF0MATQLo8wA/uVTLtRw+/PAXSFzuj3j54fUg3VkqED0ZgJrLgoz6eWOwb2z9FwTLtDgCPwB
VpS0iTUoCVY4816GvL38hK7PnqS+8a48VL4X02xPkREGTfTlP/H5V7JDQke/dMW6f9HlASvs9R3q
BNFi02TH/x9ygVHEtdnQLquGuMIRrvvhWepnEbH9oWY2dgViGjD0DE5jP2r0l3XYhTiv8BG2k5r8
lr1rEhLF5BEwQEiJnaoXf547n2vgxVVB/BmNRYY9BAvlSfaezcos1x2mFPsKGyRpQbuS+bkWHfVL
TZiKNIe4PjSaPN23FhqcI5fJDdpzVHcj10vNbiF4QDWqh0h4ZBxBI3DzvzCVsS8li9OTBsBuu50e
0zqdF+nw4UrvdPHLMUBXoaPvhXkE2r5Q7xs5qQdZESd0HPJAh0yC+QMoQTRGsJuJ/NHu6ykSyE3J
fFEyByk7AZ3KHLUd7/ymwWlklJJjjeAqDYrqRvT/+sFw123LBUy1NIKUyRgvfJCUztptTyYjiFjR
WhBZI5rySpjM6EDsGBiDPjzAKWTz9t2KR0vojNhZxLdJQLaO4tovvp0tpixJYrJ6itJ+ZQcljNqc
omvpEwZMG4ziZ4nQdTGMAxfI4lIjLem8wNu+eBNs+VDGRqsAx9odeyQL4od/QoJmD36J2ZUyYXcL
Qj80qoRnIR/wCCGJapbmogHhajD5KqsIhFw0UVF8sYbaW+5sqdOzl0PEKUpqbX0AFEmQYfj3D4R+
oFzkYSJocwoBNKurutC/PR/PP4X7s6tEdSKHmYpXkrIkgjESrR0tyPcOkk4OJE8by24bdjLSWhdr
EO8cQWhPp/qI86Vq7HODqeQGL3PJyHyYKwwFRy2R5o7rPe1LjH9GjIoOemFap051qLPePNYxW1qV
IEGZnXumPnjl0oTpT29LzHgB6kWtUkJPSf6Xjfln0ZlEmfMNxGJFVXv7Qn11LYzb+EMreI1GC5c0
ljeejB5hxevwIan7/4RXh7d/o1zIiNpmE6bZUwgAZgmAIxCRmCqmkD1UOJqWmWvnvw4UDZF/4OVo
EYylHRqIJ9yU7plt7BIp2uAN1RjksqBrU2+ZZ1lMTY5VSMaWT346tcc5F1gFnDoSUTIlsxES3lCM
xfHi2Bbc9K/lDg/NrXQ3Dx6iWw122NHRJh+BpZbGotbm8MFAbehbvHgzm1q/e1IcX9Gf7IZ3qXQ8
Z4GUFLbAiuTR2IRZQ7J3lyTeRPPqmEtYIJ/DPJISMEPQK7tUnozYMwmcWDxmElDzEPuns3Z/EFrf
IfE+LSV0w2VZw+bYgib+Fw08KEgezErqX+nvSpCszWY3tEiYNTyhxvHdKSLFJsSuA3hWuNJfK602
vm9Ux9O/s7z5TUaOKN5KJnuPpEiLYc7Ml0SDw7BC36JY8m8R/ZF4hlJpTRJs0oD0utyRJgIXAwPn
MzVSJ7S3YN4YKS0XBbmV4qr0PTrm0e2wkLMBLzIc8yRc4vaHaGajtmD4pJyi1ugclM7hOpxnODQm
s9KJe41AGCmq/NYoAfq+8xr8cnCr4wzSCy9NZAM5zzBoEPrFTNIyXNpWb4jkPzW4ZHdMttI2Fri1
0d91gjVAnfmJdO3MbAYfhbFdFKdF6SEzXSa5u3sFcWN1+rSW+PTWjmb6rJGrqE7cbzyTe/5XPe0N
VV/MvzcxRXJRZHV8vor2pR2gpLJkuIcAletuyXjnxZawHDanWjizsDGCnPgiShGSUvhtk/1UFVmM
n+3v5lhjWkRRTXzL11nAxSyNSYJaA9y6nljgJgVS1Jk87rkX+pLfhlLU9TS7OT4qgRzvDjuors+u
SmKDRrT6RE0aTM5JWIq4dcpF2N6Oa04yaV43sRja9rFGemzXrYe192x5mmjopYdg0LssD4Jf/qNW
Z83zDgEjG3Oi/QkRLPW0zhgGZx20tNfPH5/2lgnLh9JXgw+EMiwcJi8igN0Ar9DhOu6PhiHHzI8g
L+Yc9gp1et57r+Hs7XQZfCZJyRdR
`protect end_protected

