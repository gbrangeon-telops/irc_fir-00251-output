

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AAcalZ8o/jQY7YVFFozBN2W4CJ7dtDMmc4qCXcw+X1HsQOWsjlnqJ0ExLq/9HwwPaBdBtHuX8sNt
9MbzT1NoZw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eb9fumGdx5oOSTot8dVQVSjhrvPnjy5/uUjD/aIEqv1QEwLJo5EU+m6JllUu7ONkl4q2pMcv3yUD
DaaWMJ5SKNM9IQtYV21pAAxck+unqu58lsMHcSYeRXYcYP0huhB41kbacBO7fQsq8URHfGRa6NSF
6GxQzFgW9OWA+QBW/NU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EWQNTRM+yXYG4PYEP5SycD9fkQkTTfcM6sgjpG7m3z8pRk88pPYs5UwluFbB09hVSCMPYEKLENX1
JIPX6A6AjJm02cmQD/SZk/c9uIP6nVMvhv4HT2PqiJbMwRsRLnp0RV8WJNl5IwtzQhAltPQm5tcZ
c9/ABn7qb82RSMRxfzibhF2Uc1QWD8PnV1j6nVmyG5zwtPXyKG+iY84QCANIn7Soa/s6m+bpOho3
0pAI7CU0STIdsIAbeZ3h93cun/ow5TnTga8aw0A3DbHVrLc+5xM9M4rs1eiVbJSSdL5Fc7sYK0UO
cAQhBC40rZd53OFEkTfLRVfwRFeSU8VoPsBCag==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EUZqFPEsLcyFBckZdNISKg5E9SpkAkJYhYdYkwRh/xgSz3PN8kMAAO+ttVMn672EPHPSTTeJWt1p
AvumrJCguaLVBM7NIXSVbD3Ckha5a0glBfzxCIJFFOPOOxZ1B+rxQ2W+YUfoLzcw9DE42G8bHsgh
CvpFN0Szn2edsSc6Ou8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OK0W/E9mRq/arn5PVxkw4+3w3BGYpl3KNYb/ZgKXRQbbZBHdfBtfu0H1VHCuj27qhD0QdkPpdnd6
gHcvGTEag6clv0PLJ5PHHHzcIl4hIp/MStOr0nGLUPNhqZtLAZRqiy0IB5ktSoIvGu4wUrWu3P7t
D9RQYPlFcbj3tpqdazX+5GhWSHnpe6FaCtaWmer4ZDmYZIG1oGk2h3p7ggKQ3amLtCrg9RLkGQQj
yEO/bz1jhZ65yzQA9tlLPbVh4inksrXMkvmJzspRm61mhZF1ey8gENJN2v1TzCuN2XD/gXtMbo1u
8igS7KocN9wbd7hsHdkLAK4mTBcgTG5pa81agg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 998320)
`protect data_block
md0Qsq1p19ihJGK5FDiONLil4FktxpMDGLa+YF5Q4BjmIAxsKLhMSsiqewSj51SNEW7L3kqJD2Pg
QYqF3J6wm3GcsLvc8fMjSq01+ULXsR9YZ65VNWzZiKUg6b2SGEmnfiTUlE95xnDtnkfpFxTNwPK1
AlyRsk6Wwpspwl8m/4Pp7KkKsypoCB9dmwL7mGCvp0JM3CYlFoJSQ1Ib8+LgX3izXvQMEaTKL51i
sv8ftjpru4Ae0nhMKG3t2SETJX3QL7w8/WLNyLUyeX5gJNTrDEI+zp3W2TMpqsn50zHg20noMKYf
kzghUZ6UicngktE6InzA14tnfWJSOwHeEwgAAHX/KS4qESvungor6S88sDtD9YPDCSYs40cqB5rJ
qHr7W8zEa6fSuKDYHbOTgoSJbDuEXzl3wu6WW//wOfgtgsknvAFMrnf5qwXwF9+kfA0I7O/a3z7g
4RQ45T476228G3eKR1FZ2YrTqyd0yzy5G2L1SyCaipWV/lq67Pvonr5LLQdHzcU/6A6PBAPfHo13
PctN2nocCEGylDCmFcNOSK404v8AeKIm7eOxvTyhQkEBCfQp9FuBbzaIMhX/CRrJogKxV5chhE6g
9Yw/v29PSXqKZoiJyFLQVC/1PNZq11t240u5EDgJgCDPWZdWRiK1dhy1QkxNW/JCK+7ala95Ghns
mikwFEbnj8SoUbqTYae+OVUNSFbYMRRA+S9xkbETpLKQSkj25rsLL/Bqn900NZrRE817Y4PY2uOg
gpsUQLT5NCyqB5VtsRifYYc51ziJvuvgxHuK14qyJc8oMsP36zJvqHDxKJPk5W60afFj+u+bzJ6T
vBPlxUbCCldohhhqU34uiFkW8PWXIGiEhcM4XfjP1lGEOdfcpr5LTzeaMhipOslQVB6oDBZI9i6+
Wr1DYRCkv3X34ktxHIpRg0MUYp2lQ/cJu2utX1dk0ZrF4PomgPMmvieZoJ39SnxwnQU/S+Cn/uYs
GA48rGxvVSyGoQt9MB0nmgdsFQuWnm9FI7IzBz458Ma1EajmNGofAQw31pjfCly1AFZl7kWruiW8
PN3gPXgYJYdbFNhzjc+hqIDdcqxxf6RhShVIZUQ4CEmGo9PcL0PSOSV7xaXGCNXZu/AWmG2Dt+IG
B/+HJCUczHrto8jQ3lE7IZ5w4w6Rh9OROEfQvIrVtXmVKCWVXvJk9sFkWUEUNrxZZsuLwHb773Nw
pZw8CdvNEiOORrpFss187oElVxI97138Po2BW71Hgv3EkLnsSM26v4dLK9QQ1bJ1fwRNtnfSPD5W
wYL1lzSGEv71UCF1XNSG2NIB25wfSE1TbZ3GgI6fq6YPDDeu+hw3ULGVBRAQOZUcwS8ImRVtkdIw
/iX0NuszW+EdIzuVisSZsiRqvcWDZ5kVG9f/r2Uj8x9xn+F47wSVakxwMk6z0TJ9+wZCFXCThc8R
7icoC6qiAuFVzvjn1xwiNtwhL1uHaIQ9qUBP4oQho7/g4eGOhTmgZJZAf3uIfBXFy6IzGXOTKiji
QF3D++UpGIALStk9BOIJ5RcczH3pCggibKjsJ+AOtmBvKxMG+yDPXgyDxjTADZ+svVxdkNpwctv5
p+00rARXAC3jGD7sVhG8BkZb4nXGLPAJltVQ2M3kw3HKx6lAP4p4NJcu6bKCzHYIC2cM2lRBFu0A
ails4H3ElqDW6JNmsGSjS/JtrU5Uau6ph/gRGnZXvFIJjVCVQ1Qk4q6I+2IHnwR/f5/Ej0GZrIRz
5CUuw0M7TTBFjJE4Gg3hehsi1T/YaEi0JfvkCGu+cmPPQMJEw6n7jE89ACYL7KLCW59vAn9MD5ki
LuThZ5Ft85B94j9HHF1h6EVJiAcJqXJHP0Hcn17GcSxbeJEqh6Wx86SJ7/vgt0nxkhmVOSLHPo/o
YZz0UAih1pfitZ8LxZJXKUvE+vLaShMUXjEOfE+N7sA5mu43Rk9HWUppOP61ZOfLJ+ejy5bV5imq
hZKplhIy3++6gdb6s+uts9e2nkOWBLPt7TrAVRG2l/4h3uWdx1GSlh6FgPTURxESQpcgHs8eCVlD
vhgTPk5PMXytwKua1JTO7CBD91fM6L4tNpzsSmR7WmHnOXe4yxv3jyIn98yrdUSWnKhDp56ffRdO
8m794wkRhmGWEipg+dZwPTu/+x2MnxZp0ke9rwX6j2Sl5x8tVWlNTBOgRMbT9WiWz5vo6iC8Q4kr
FeA6Dw3Lz/40hT8POF1gtrQhO5EIUpPUbxal+K4+Ct9zivYKmigtI+Z9RSHRp6DSNiY3xd3LLRki
jkqA0UYde9l0x8JP0omoRDFGPd7pxS6jI8Db2mUEOWgOW0o+iGHiwmIHJzLvPBYOsK3JsbGUQFMR
u/XbnV4DhkdDqU+8nacfi5S7kEE07zWrrI/3wRYQnmNILW8UuzyGE9Uw5IPDVwcjIConbZkAd5Ww
OttoRGLhQHnQyu2xww5UQo6Z3JwjpjWTSWmm5KMTgfwmX0/Tl7Rg9p3WVRLRyHSTNXQxCSrC+1aZ
4a1mJTgbWtQO8V9Nt7wcxYyLz/Y1mLewJ3uQixpSocQgm6FC1SeXobmk42KLaOCVggdOD6Uad30y
boMfTJ74QjX5lMHPI5Zr3WA5JbshIHwRr/r0KkkczqKcbPS0w7hLRfv6fkd/9+AeLWdZ8TCpEnTW
rX+hvZcQbdJtjnhtw4DJUIxb1qBRZBiH/PqPH1ELn6TIv+WZnIsKABvlR+g3hxWBbWB4LgTvyUgF
6U73ageZxgyUzLXNbS1tv9mVBCsAU0s1nJj5QndFmq1BjCwcK/jm5WiC888QShPsgzxdgxi8nKDy
+kmCQv3BvTTi3QG7fhVplyw3kNHCiJCWw4uOla08acCuCLPNQjefYDhVJQAffv9tKUjdTtsFWztX
dlaM/BRSGSir/WrXpoDl+razQ/FDfqlSmTyq+7POwuukQ+zMHJbUCpgb0gPP1k+AzYh2xcm9z+kP
3hm/Yi5AGq0/O+PaT9NobJlq84Eo6B0xaIRf88LWMUXSlxlFwVsv6qOIVZEn2Gyw3NU/JH0NG3HT
jPltoJGOlDEqBkNUNLr+xyxTMIcIeGpHiTJIa2z1QpdoyZwqD7gZ0YR6L5HcVkES1Kn2pEjS8xFD
f3Kg4/lEty5gU7WVz3LPbrjDUloyV0KdNDWo2xkciaDxdlBlk87kM2jyCRAkAbi9SC1Rn856fDxq
ERFKIqN557TGT8QHICPLwRCgGds4A0HP9E0jHi8c3tr0ESBm4varZiFP5FqEGIHoa4DcGozbYjf8
CvLUvO19V9yWAOa+vbJoJcJPNyAglAaF2uaKNXxr7olxzKi1dgzh6PuQDrLBJcA1PsHmpfiDvo6P
ygHIw84EfI1vnEIAOzLPHY+cIauGYGSTwbQBuIxBXjPo4CNSLJ7ugoCR4B/3BKg8zU3ruuHdGGp1
AlXEq5yDQIsXuAEDb7q+Gpf8Stk47H2lp7hCBgkkGwdRp0ng8k4Yr+uh37XUpOWA9fOyDezxVZ4T
JUVFc8ty+zDsOz6jvnxScLEvEmqasXJszqlxPWbRWN3K8Ra+34ivRQi9SCCeQpU2W80Sp9zAq4FY
2KwXCBy5R7WO5EggRsZsH8s4+l1/O87o5oaEEo0NBTuQz6CmcSgagkVdYZu1PGPp3WMtf5lvK6dL
VQHDxoGj1WSfRw/VbT/SzWjak/lhTQ6H8VCAGrjzvhfUpM3R7kFxtEtEpGoqPfqpYX5kyEdYopzk
w5HcEchjiOjaRWyG27ylm6gz4N03FuqxBOdKkjuquEGZecT4RI/wYP0KQ+9uFF0NxYPnmi7M4j2D
kxOPmbaitvxMclkqxlIc8wySzMfyeAzu0lMIRxH0kZjOm1DPpws9DNZaEtihn7Hn86gsBxMNR/HH
ueVWReXHG2DCJAxNFKMJ0oh5eZt1JZ8Gff6gdMsmyHPe5BMXxnMLIzlKnwhL0gYCcmDxq0mAmCxp
Fxq2/uOvgQkVtyHcoe0/GKNMHjpwSyWsmjK1n5iTNsl6EV9xYmRSqHwln06uYFfMLK3iTUmmn4w0
ym0dEMPQPMNQJhGtFqJ7N5JT+iZGIijb7v40p9lQZmvYQADj6IgTeS2dhoF68ZzyPx3w7hTX0tSZ
jlHNigJbQLcMVTUVfUEX0j9Zgs+NUwMXg7LNaRvMDuxL39USf5Zv5BzvhRj0g0g19Ia1ic9Y7DmN
BFcEcwMT55OeaWXSC2wQmlIpbm9sfFp24zrVXqrSSq67C2Eifg6V/YM4IEdajc3XOqF6sR4nCc7G
XxhBTuRMtISmcCKR/6BYuPWxvunLFKJmEtdqa+5wz6W1mSh46hUjrvMpUW/i5D2j7k4Lt38jE8EG
EvSlZX+Hdcn0m5Jy7OJJsOnIdCCe8l+ZPRB+QH1Kmn7LDDVDNSgmByyuoYTgazuijmZspaSkh6bQ
zN+o7piGi4erDmt4E3jcUvqwcqy6RAQj2dwwLnypCim7Jxawnij0Kyd7sV8Ppk1Ip40q+AWrse+s
gBnGIJHc4AghyGi6eU65Hjgy0KLo+4wIkfX+B8s4ljSRaMgbz/sIUpKk9XqGkSG3SMUvgMvJvEzy
E+bhCbWq/KPkacu4okYSsDje9nvuao93m4+ddgAjjqBfr/xnJ6sXGGBktvVtqvwtpJgI2VDTokgt
plvKJx2SYuVd/GMkTGrU2jD6f2t1PP+7RzUsHFhNB12YamB2YGjiywNibVtuUOcJR0P6cRFItfhX
xK1+nqomadqOrhVai9Zi9dJKNLv43tXpQjAvjDLcqMGLYtcfQA+9wljraJ6AV40paUh4A+M4FNQS
dIEv9UUK6aC0a5k5MqwrbK+PXUTrU3s5z9OcKoeoHr4GR8EUH/p2YRvnoZU9+ktcZV7aBQKEzxGW
wp16opkMU6WSCN3PdnxPnafVLhh3uMw1j8qfRgPYMNQhSazLHBk7xV1dfoyyNdMobum5OoJNQ0IU
78NOZSJqe2kGlEbBdRHQlcFmKlS7KoL8VixyKpI83P0eTxceT9uvlqwSyl3h5T2r1A7ptVAjrEpy
7y0Ld9OZiDyFWu8p7SX2yW9OvPcgkc4cGObAJ8oFnnU2PhZt1F/anVT9GmMIeqo/7XrQDDr3GO2l
6akZSuuWAbpJpWf6wyNDg0nLyzUMGGvBCg3jxHR/O9ZgAwLBnU6y3wuCLqGT/YZhUA+FzOOQqXfl
oLbA2lX35knizDbAUQEojex0D+T7NPLGsOPnMaNNs2KbexEa0eS1+Diow1524rFl23tQnX7Xt1Cp
/AWe0CK681TdBKoAnSUqzhzJhpm/YndUm2k62l100z9vgQS4qxFUDmqcsJR4YToXmvqPE7BLskzK
8ji+QW8SVq6eDkHyW6LzyfmF4osDJPygLem2Ew98YrS+7xyMG/3c4BTqgH7ufdI9HiMPwpsS5TcY
+MhrW9NH4PxnAi9NiNLWKP3uCc/EQlk9H7HD6nCsXI4U8FTJkoIsxk3O+px51ZaWhOWoKngjGRo8
L8WofNWXOwak9NSUqFDQleo+CkMCmmvroJMa6ltDxRXJ7sEv1keOpQpcZXl51dKqfBr8sKDY+l7+
KPssPEvbdDVztqEvf+ZE4Sk9N5vdgYLOrUDRIj4RKOqOFacJlVuj0TPD8dgVUJozbEWP97gViBQg
7Wa86J5U7K05juff2KF/FjzPkGuiUwXbzxBZpQ8JMRlYrfBDyYedyUwZ7Ol19CvDC4FE4IWA5Idn
HvRk20QAE0ehlrJWe7AwWABzsWfrWVS9741gdBY1j9u9AxAc2Xo+LtfXX7J8CEZdQ7Pae0j5CV8C
18DZb09ABeiNt7z1TtwlmlYibWy+Y9OgDSJaqZ1IJOfcOdBereLiVPZfTWaRSU2r9CKDx/5p9+4g
JyAI+8PsBBqURsh2+6VaWz81C2/QwjDyPls6f9COfFBkUEKQrTOHABDkh/9kbnLUv9uAfo/WUTSX
IS+JzJkp8X5wsVcKq2kTX0P0agNKGNkW6c2D24Zx4GUg/PhMGQJF62duJvM9HjDPpUfMTVMS7dDd
mz7VYh+aV+6hZEH5jvSw3TVJbh9/SaUTPgSkBGauZ+yErprack/034D3dGxfbanTTELmFNDOHVz2
qGXNogbNKRGp9hxDWjRF/E9UTjHTYaL+s5p2zx6mdY3olHAdjDr/6mwlRDi28qJO+kZfEy9BC28W
sfOJHidKYc1YkkFHTE80gf/3qTHpdKt9VxRTo4vKEk+D9umYd4UsK33dnShacbSyK7v8X7Mnrxwt
VTiQ51MaDFFzoFi281SxmLDBqkeYj9lCOsKuYxHpldln2HKHf+Yf6cUQOP53M7LHMqJ2JpbSJqNl
zyF+dPT30C2VyBt9zEkxIwr/m1HnZ70dt8W5unqa0h8kG2XP5dnE8TeRqPNtAC1FQ46IpxArLTGf
d6nDbKjiTkUVvZu+UgJn0XDr4SiCQbw8uReld+KhQbiySm7MDDPki8WdYW277cTU6V6dQ0qVVFnp
qChsFKHCFwaxinkr2AmRptgmrP/kcCHbXWthwYFDfj0eE7Vj1z2SZEZPotE0wbzvvZPyrlgEFyAW
aZviI+5jpCYBWLCVsM51DXScAylzasxpCgVwnnIP6MNthdK7hg4KV2bl8iPjYqW5hQaMYlqOD90a
Yoq4PcJLFFOwKEfC2gL5cdM5MnSgfjm729uq83//h5UZ/a8FQG3DIEbhAR4MwTnV9SRbS1CySt0R
cRAOlSY18IEAaI5nAiPOUL/+1iGsk7ZZKbrVymvDEBVm5SyVw0AVxsZadxXfsCPvHj2xeqD4/KCP
AdmmpQ2fyArtukUfTeSOFfc3x55D5xZ2skpBF+WQUSrDrhAfmdSJBbT/af5YkJxICzFJJdzWM2to
GztBXxTyqbDhubHO/66Pr/FsTqcWrb+aKGrzQgDQncldJugxK57m8Dx3CGZfJWtHMNLwS8YnURyO
qWcDqLZ7Z3hAADSHRJOAdTDaURSmMjStXs1i3gl7wsBsppmAQFEEAvKzo51ZxN02k+GmVjy/eSEu
b8ToJqdvt4yXjJHLxz/YGcGxmBvA7k6Bn85xIejd6SSznW4tdClnEKZ1UHC+qa0Ks5C3O4sv1M/U
zZxs19Rjd/d2kefD2saEom8OjOSr17rRIE5A8ht/l4Zqg+kEUjIW07nEoQ6mOLdP7K4QLA33EuLa
+p6IE9Ank6qtIB8CRW2H34i5ocas+97X5WIRLv2+FhJ+VSX6PrrV6V2sJC9tso0XZ6EWjD91tX/l
EBMOMkDcAWe+aPpJNzBd1gOLLV4wHsp1rYdcmESD52zuwQ6TNfnhEy82ZyipoHD/QI3/63pTxnON
79sr1AS7NuRLYS1syR3iAz8FuIf9N9DWFWWy682HXGhk1JYfUQ4SdBOKSbTFvvaGUgHW1JbE7LR2
apg9ogaWFSOu0beqsJHLHupbUr13asQF+cpn0s5XwxijAXZZXTrgJxPFnxSmPExEni446K8jF7bC
/9SlDnshTlS0DIQUL+eWKUOI61x1N8VwmwdRw8v/nIvX4xyw7UgJ0/O9E/ieKjg10Dli7aU33CE7
DSeUSuQbo/NpQ7bfSucNmbRFDaa/MmVo4VH2x2QitzqvrKbWazflW1pkseUUw5Yev+N11sdibihy
BMin69mHJeh6bLXOsszhLoLnzuDt/vzqZpLIDDWRyQVRSWBOr7P5/XNqpiii0vvRrKSM0xOEGHRP
o2Nn1tSsKOiP02E1dnVbKSYgjWV/4Npj3viQt0NgzoWdH0bkT6TCMd7NKD6RopF663KsmpjlcnCE
ORayPIBmgK+9+Q1aCRtb9ScgQJPeocvcVHpKr7aY1dVUdDMdXbEfv1FTySbqomNLarORqhGivns3
uPwccdJZsrYd++4rHbAoFduyLJ6DpcWo56d512C71tY1kQkNvi98gC6m8hJgJOdP5NIXQI1aH3nn
FlPJMe2vF+r5zvp2762uGOdtZnduulDdXXCGsu2YMHRFqN5di2fLWjr73OxomNSRdIZsXICiWJs+
M5G0VXwF72eRUSHkQEH9Bt2C/BGBOLxunM2qFhDbF8MjxidvIPkjRemEfgK1Zzjr8jroZ/1SbMMh
xSF/vEkz9OxXF/9/S1pdmJHnMGRw0L6Bo49SWfLqanZSeQuid6lFXI9f5AcZ0IbThCOussJjS6qw
VDNb+fjEcwJpNwdaGOxZMyMO+48No7kaCuP3G+mTRwO69Nozk2SC+OrPec+sOvu+aH6sIF7+djK5
jXzELDpLOUSUUtqB7qADqsaazaHRx97IBzMeM1Ds3hiIWlpwT/OtlghQ7+WFvaRiYKvHBD9URmv3
4Mb2/W2qwDuJmFXvL5sTTMuR7NZhcen0vKl3otH54uY1cqHxzco21sNNVKPz0LBOKNwVkyCGuILt
clHkOkm7+m5ZxgEpLr9Z52k7b9waSft/gU6wvv8p7LwuGTbb9ZMB1oLXB02A4FksAqk8D0kj139O
Qo9OZv04RF461deK1gMeM44nAheDg5K0HBdBmvv92WvegzlovJNy4bFFJI+XMWXVUwbCUnbrGsEk
WKq6DkGy1ZICxXc+x0A+xOxTmzsDHrr+5jcviffm60gqjjHoGTW6KYMQuphlqKrNu3cjy/928TCF
ZD2dWNgfYDOGB5UMdeCF4NkewEcw2r9IReKEcpZIgEjABAEDLpAOrUeSKM6kUJT68dgiRaFe8qkL
PWDfZUmE1JZ6gkXC9Ky8qCdVFuwAg0OEc9gWFRcGnWL2iEU8wl1yajPvsAEjLGQ/2C4m8vGS+9Im
dkwTpXmC0r8wGAxv7DPIawusNL/zTu2ksoDrmL70+Ibpj91rQJqRdUEwpg4UkJ5B8F9SyKWQZ82g
JHV9SztgPbdtXQTqt/UME3eN7E+tZDxy9bT5Iv+DyIKyfthTCX8VsSPdCxeb7cnFeWFdhhvZr6Pu
eECp1LU/Hb3L/l3x7nN8hU9jeYZgO58+jmMojoDQAx8QDCa6YMXnkLlIjjLMxh4LbRagLGbNCtvp
rb7imb50tB0uwEnL0eBXgDgGngM+z/mwOkkL14G5hEerOn/Nhu3WW1zMeHvp7H3ojU+PdlfjOKgi
55iRSQLWsaEJ4ItrRroE1QzWsWa95OA5EJBYZ9uHoGvqPte0JvEU3DUzHj0a8738uhdUz+pKqNK1
ItEvPRoOP8pYWnmGEnM9dMHFa5021NNToGC+qLndSCBPSbldW7ZwM9sgTpzbUBM0pPKXf0fQFRIF
9hvau/1i84rE7+ABE4VCZT6Gv4yTIcs8Ns3MNNeOdEzhulobOK7idkvwVqmD2kcWgdMgiEUBNBjZ
q47LNAxYtoQ166nIrOrTnRB7qPHc9nEtK7Y9Zon5vRBzH2D3vWZhUBHUWMTYCnm3V31rEqfvQMft
3ekx8ou2r4uMufmYhjLfT/A5Lq0O4Mr82HpOfqkzpBPIeH/hLNFu6Fo4iAEKTQCHju+oHo+3bb7x
MKEScToSeFEum1OgELfZQcxlLvgVGHG/0ivXPdRxLTLLdtB73JTAl4jLXNGzhNybxMP4SBt8+vHp
piZM8mNi9XWX7is46qqbbvGj4krg9HKCg1ggMDwPcxFQbCQrRf1bdUdCJtAojO08CSi+IjwWZdFO
vtrT9cGQLmeRTeWi5bx8yC/DT3PBTo2DPvNVIjlGAOle4HeSsWr/tBqehmfGNO4xw05Tzl6pX24W
66kbDccFsCQCO2mVd+J7bns2FESI+loalwjgioToHRyX3njmMF7lp8DRTFIuXYEKJNrY904Gj6mv
vr8IHI+2DcdqtIQXXVcydSM1cPKuYdhwAo0B2fWANIWwrXRFXJ6xFQQ53cjLZV6eRi9frcXuMmol
CF7ZVqXvRlHnFbQbOu973ZuhSZwC16qvvI1lEpeG6ZK88isxzo9KbeumNNf9aRlrmeHtqQeX/8DL
lx0XoC9g5Y4N0S3p8J27FaGFxZei20LweVkS/xBCzXQc0bd9gyKG/JCfkI+oo1eCv0k6ZTX0SNYb
IZQ1Er2FHX/nVLENIwqMpD4+s9S0uxdnv1cGz0pvCEVq7f6eByHlyz6gxqxINtNdPQ+6BOzBo0xa
nc+gLOrSb4V1Zr5Jju79cc4SJ+qv56EcZe45sCz+Cwldtuj7iql8ALAV3viSvd1rBvFJTPXqmgy1
OagAJyBFtlLuFPSAUYVsAOeyxeBo3HnlJX42sll9m1IQ/KW4dvyqIyaBhn/vvc2eQbYQraAmIx/i
JCUDSN1RKkSAgwtUHT2MqmD9MqBXuN+TApQV/8D36YVhPSW9ppzXUVjHl3hw1XxIa4oYyQVUX8ka
tes/1o3OOUOz2We5o0QuAT+o9q9nynmarN+JtbrCcXlBoXzbfGEEUq6I41dsIYvNhHa8tPAj1EC3
c+6uegZM9eguSFnIULl6w8N2LAOkl6echcPsKzeAGbNUQKFGMUxp24jFLWhwKt5hTiXXg7QAfGgs
HQwBgQ0sGOVudI6La8/JLj8TcgK70qm8jLA20m8y7Epe6OFj9sEGVnA7M9SJ0+ifXG79+9KvAWZp
zAmFGjQGvQqaMaAsIOQsNEl1XHITgDMaubpf8MSethlb2BPkZOdGLJghRxI/PqQ5tjIuUOfburDF
cGYXWiMf6V6pvJbW+Eqt3zs3lB7nZOkaNsr2ZcrLJs13ewoT1r2MVy4zXChjIhtWu25gaWbZb0tR
5B9hwMnpAvzY5VkVdPHEhDqVOrhQgVJmoNSpDC7pGApgK4UyT01xecqrqYB8IsIsrD/nTLWqokqc
h2HtRAha8mVVhFJZ2dyncrI/gMwQidpmWSHH413bRWVyRaIwGLDUN7wuAv8VRmCQNxSq6wVSTmYb
H5DkVAgz0sRGYG0xMEBwFth3MUxWRPHCFZMlQk2Tvg0xwlyvCXLVylTe2UTR+FrNQV4mg+gR7aGO
x4Jh8hkcjZ5pwxXk1jqrCstigX8Qm0SguguCBk4AT0kYP+98i6+FGgKJ5IehAdYjZZtfZB+cVkHT
Vmdf4E2i7pBCBxOiI1z2zg8ZDL3ooHtq1KGeWwN4M10tIbkYKEXAF5Bo8wxxPhlwe5xm0InZacU/
ZRuryLRDydUKbmr9M+rqfscEb4RG5wYxPu2cpSmLQ0SV021yD/dKzRO/e1xpN/1mSSWsZwfulixS
Z6/g+7hWysCdnqkDIEz5x9Dle0W1g0sTHs8QrrhEmwdVp3TQI0+BLK/4GZpCLpv1KGxXEFaSFmFg
PY9A9Uo3SdaYKWOe+mwtiNrpavXWUeeqhe77urdaaYEyoccvqM0YSJTAvUgFceFgxO9OstvRwdt7
pnonSAp+IZxZCt9tbPc+rZA3fyRzSVkHS13xW8ahROVKthLo7PhjqGdIgeLybFrOI4Cya7/SBHj9
FfLNbkjdBBhdCa8wYRglKHqJprrqe7XxCAxTh6q6bdj8GTyYn+O3hpujJCdxW+AKG6qVmhfywUcO
p88qDv4lByMDZDSeFfSpR+ssB1pPEctQdnyw8VEL1bSdcXtb78Ix660vUD+POv+dMoCR3HiWfWcs
SX+ZBuploKprLogOGCk7P7Dm4g2cwKxgyZLjuBnZszazZdPBw6dXEJQsCIfAtCiHU1VjrKLmIwtl
oOlEMwB4gNsHuYDKe0ESNBchOmFkDJMB3K6cF652GZ9YCXdbJGbUcjQY8Tj1esOpojOetNrmHQ9c
mo+sKXN18AjDNLtK2fB0cAU/Kz1z+E2aZO8QTAGu/hdBKvMjLF+KISCh68Rtu7qEt0EOV3nwu/yF
GKMDLN45iojGv7ALmkSLwBaXFeZkaWH6911idZ+NBfcRsZckHWIuIr8s4xoJsTz8/hOT5YhuWcVh
we59C5M3pLHiSCxikY5LBdQNvkhniXtDgtIbkTSaC9fdAsSxFTK/T63kVn9ZyA0IDYQeOYm/hyZ2
X/cA8nbbIGkjl98F96lMz6LB3jOAZ+wRDDsj5UzopfN8XTeKpZ+KQE+EKaRCUHGW6nzMrHcWS+tE
l3uJsZbI7gS9C2gnXYBYhTXt3zPcC2BW59Z6vapf54aAKdX85lXkksTxeVpAkVXG0zZzs0SLbcjN
IKRFvc1/QcUYejReQxs7g/oUvdj90201pFcT+bNkVDb6ZEqWxRZ7/o4DDW5FyA/uQ9O0v3HUDpLx
B2m5PKKgSamaINmhriYOQMYgnUwSgjGUPa7k110d6zrQjUrh4ar8n8g1Pc6n9IFS8W0VaVtf7XxA
5/cBhJG3+uOjKRw9f7k3EB5CEWVT5uJzPWcuVyZGQqwG8So7emPj8bkqS5PY1+kqzjHHnJapVgJG
P5hsPNlaCxCEXloOcLlKQl/P42Rp4sn9z0vQNN357/pcss9V9/ubYRzblS6ndlpBxVueZ3ZkGrwt
71Q0gR7t1Ki7Bi/20vdOB5Syna34wnK2fn1TZEX4f68Hp5AzjbZM/VsEV3s7Adn5XXHMCj5TvV+H
44CTI/HyXPn2+TYleEw1HVQAh6Gep51WHkRWHjXLsYKZD9Jgs9d9Bk+yDRUggnI5l+V7cxgFHDPH
R2/ZClAcOT83a5qFNoOzbH5JmV1ao5YdUmejYMYcXcitkwTNqkJ7IEIwmT6OeLeOJSCminlv5vWv
jEc0l8/mnSGw57hr6IoYsC+5InBN8Jg0fbjjeoow1Iq+y7mT04GDKTyXY/qrU4BbHu7VCH47qEZE
2sa+Yhsdba52q0BP3/jBIs15Ba7JBPKS1nlxK03+v/+qXecUVa9AOeiEynQyWB8sYi/PAkeOjhyD
G6r/HuzW0MKN8fPkYaintS/B01PZ833poxdGOthbrmdjdrRgIprHrJXxWQTjm4uW2THdRX6RYVTZ
muvJrT9KFdYlRX8418dJpoctufD5TDtRoNdB6QaMmu4iCrEU3TDy03K7jXm7M84MLWYr1gSGUs5m
81wJ4PU9YEgkTR34/0M3xD6QBLwWaz8mv5+WTslC0Xg3RwaRiSX5U8Y75dEV5wE24iIq7JDePtJ+
sLnA+jfBymAGhKDse3sD925OxEv18sTmtDowdT9WDLkq1eAHE+VQ4SmvIbge4A7N4N7Q1Uq+AMCj
8dFtTb5T2NTVXJzr2ICT6arXpznP9atRz0VJnv/qx2VqGsh/kd0ucdRVZFai/030ElkwKpFudszZ
k7lPLAfx8e2DiOYIYzA9VasUKNHUXUCg83lSJ7CuaoqesqFgfpBXu70ZyZyjSDtfGv8jp3AdVPJU
ml3Smqw/T9JZrLVkYHUtGLAqh4o24EMNyhM5ppD3fyoacXIjQbsfmrEZ8671c5W9tphtLmen78o1
jMMID2+e8O0uCoOgNDkMmHp66d2if/vPnCSGQ9D+FM4UhAN9DxojeYYyW0Q96L4vh2NuyUPSyZTB
j3bLcn6iXXPhm8hNii0P9nZ4RjFaWNJ5HyVtX0HiFezeK7cYiUf6kKrBa99a7FvxVswpc9zxL/Ph
fbQdDPqFZGRSUfMnoQtTY/OxqJrrhlbhVqJQOZSgBMvRUBTNlbGM+6vFUTG5WvaRFkfU1JwsC7JT
aeMwR3U8CoNbLxthrqLsEoFcTzhEApfaQ5NeM0ZsuQibjoNFpJMNOF3AJVMhOMwNAwO0bM70Usme
NAPPcAeOb+nTlu0V3bW5EOssBn4/FD3pwwgXz9HI+/r/4O7covuDgtlUn/w36FtVMnMn7Bb9qHkt
A9e8XMNbAEDFU5L3qSyiAQ9JZXleI4MNe1QJI8kKteC2rcDiTeUESll38HwmgPMCSaiPS6We6cNr
lToqmCc7CmNKVDRcaJlslkq/2ViZTP0zqYT8Qucb35nvQuRaTaBaQepvZHSM4zN5gJA5L/oQNWaN
BGbLHV0EYWxrAPZcMW0N4OogXxdtcjltlHD8WXYIloGgUuLDrfKlOK9cm4b7XVRVZYcq8LbtNy95
xubMZsLrsR/O555/YB5u8Lqb9UhzH3JiH71gzYbM2xzAqNeNwWWOpISWWZzPspjp9/1uZyVonedc
b9uAxinpHUoqWEyWCb5Q2bVb3/qK/8S4xXZUnBfQLyJ67wdR2aXnx3xXD4bLmt1O32QoKCHXWTZL
ilMtLtfxydGMvodeE0qTlHHY1ko5pJau4u6hUxKJMYwFMvIQ02B3J+5CCMlyMBH+5ssZ7EjnTli0
SxijlOxMG1qL0kihi0eDEuhQWfTMydpl+ILGqqgTjeugqYWYWRoskoKyxI+/oPPlo9iCR5w8kdPo
WeHbFzJpC7xv8K2iaeJz54ae7P7bf4p1y40aSbQsN+xdeABvC87bfHbBZTyN6IBA1RW9o295xLpI
VQvJb0U97xQGIjWmxtx3fqUUQLsmuBeDnL9TRwaCssXLndDPYKSnw83V6jGi/ZimKsNKpg3Q6VJ6
jGsV+oA0/Y2uJcaGFjTfX9koobgTaSShEss0/qzU0cW44Rmz+jPMSNPmtIM3fqHMQZP2LIPEfD20
rqYNNAxXPobx7pUF2xj+1W0+uPNCkZGA1ppd2vYBpZ4J8xYG8owPKO7MTGF0VoMsUG6Ww5n7UWs7
wSuoAprFC9sOuhqe5OKhPT0Vw3nYZeXjAuNdqF6DfI3nJ7cI1m6+b2y8IMuTmzyBUvaPXqtHiik/
Cju0CJ3sOwJGjT43onl89d/d7o5bwHzaJySX/x9woAN/kH5LVXMm3ofMKQG1wL7RVxFcxKGURJSY
/FiAJDeOCgkiKSiz0Mbzer1T4jMA8ZVqEi19/duJIRj9Sj/wB9CyJNU8CU76ox0pDzelUL9xfXPG
WsEKCeWE1kT3T3Hr71HO8NRrtsRBQUXNXD+NI+aoi8kiw9qIJV6GjXmdJYLCLrUdxFBknbhapHGG
YNu5n1w7rYluNiSk56FcPlzyShMQkyeS7A0AZhl1f/eZ7GJItr2vYkzaJr+mZLlFOKlG6fnPGNUk
fZNqTxHQU2AKawiBYiU8ql/L9YhgVa/jAPBnWx+ccpfwEGZ7yCire057ep3F6Zw4hODm3uS6vzmL
3arx/+KDQmFKzpKO2LB95nfyp2BrnfStl9G87G6LtW5kAn60Klau4ptFFLVengHJyqZJXkOfIlLZ
oqt0UjV2dinHXWYRiNmIdGz9IP1bv1llXr3C3XdRHRz0uV6rBiPzYdo9OfExeXEJJcidwaLm5Wom
TQXTZbUpQVn8VekWq1Wx+4BnVkqMNkS14tPfxuCI1mRBX3HKFEskc3wdl30DLsrz8kovyYdCL8IQ
ZCEwDUNN9tADWjv+/+eikxcxzOiKaOWj1WSQG51KK9Yw5O//ewf4F3+P0GbgIDMNExfwHlN/AcSj
6gnlC1FiIcwsVVzkm5ULMiw1yeJKhfD87pMRuHWsDdzdfIl9HjlrW9VEIWjAu1lq3DyRo/qzpsIq
9d5BI5Q+fTHdJ5Gfh8hjgNVxcyMk8F+kSeS2VWdTIRKprYWDoej8X3U7cue2fARpxFdCmetSpSRs
LeJMgoicc+/NJP40iwO+50gVD8gKvkEmgG/jhjyhPNRa3HgD8Sx5YrXaYxbnG39i42A0MqHhs0Fp
WgwiGpW7hPxocl6faF303+yA8oJ7IpdCqWDZyB3Io4NNA7Kl/5iJk/f0ybhlB+ijpoZHN9n20vn1
2KA5l1xyZsxrdEs7T/gHFVsp2Py3P+t78B680YHdiA8TksI4dpApYF16JFNWFHNzppfjV7m6pmhU
O5R5Yf84ZKevj3lAnGwQm/7zqvjNWS4RXB2o56pTQttDFzS+pL+bYmkhnmpxzxAilfNCKYjsaRff
uOCTk99jcl2/w8mFyBFbaP7ZQHZvRFXShYr0y3n8ruP6sKqiiL8NyX0LVemJ1++fk5Oi/HNzBGII
fN7LOJnTZcEFaBi/AwdZzBq5Bz1YftcGy/2Tr5znwyx9JTZuoeD2MMxIUx/SnuCtWFkOPGy14Qwj
YqF0xTowR5gSi5+c7jvcZKqLKOEEhJK/53PSgkxSGxW40noAEYQCy2XyaFqpMq0cDNpLKzC6whdr
p0IlNXaBOWsVsT0keS9Xe2IqQSURHBz0yvRsdQV7yIJgYfPUDohGZ7gUW4B9R8rKNqMmF/O3BCii
DokxJH7oKNqLc/KJ+MkJyG/lPsuaIterbwBTRTU/1dVGa7j8S5O2SNHfBhjdBlckVDMpuG8dcVtJ
/piTUtnXLgc0cx+aA/J8VCykSdtsSuQTLO6hEZxmqpa6Yf1zN65cJw25G3BXEJUFs07dnSMJxX1G
HHD0KNwMPzhoRGMhZ0tKdvyHNth9QOl+Y8lnSq0tf5P4+Fc3U4fjOT5NLLyCkN5Qts+9Xe91mDbO
47DLFdsKANIa+2yG5EX4X7JhnVee+k3JGYG6XnUWiGtkZCBmBAyiRcW+o3P8IorIwf1B6MENpWUC
f53z/HWPAEsJU3/zu5b5GQq9u7HZeO33IsmWaPyh0GSR826hN3f5CK3XotkGszt7kysNCx4TXCP/
8ArbLWiVKyK7WJavwdNvlAgY9Ihn+IUzyXtM8KAEq/XO6JPlMMaoD3Epkox7EwsH9WRjpOiJYh78
2Ozv3y6Nf/Wv0jNP7BHqnALkXbXDf2+tLxBVSR6mhc+JcqhM1m1+oOir2RVU5ppTK0NEdHh5hoFG
UH4cKuQB1C8Eg70yUR/RagTjmGkpFRXGlysRw9ADKG/BqOsB2BIYSwoo+5ZgSF2J7ATM8Vuxc16+
PheYgPwU7KFnP/ps0AMdF64xV+Web+19W6tMeHEY/bep+1FXTenG5tLUyLzVsct+kVMKJ0ZaXRZ5
GOXIljE2ki4Jc8Us18RDWTF7gp7DzR8TjiT995zlrVUH6FEwUHlf47vs3asHUwXoR/sV5oBezYJY
YRRFWYf+EgGRysSVn8zqJFhapZ5VBRnYCu2IqRrKhX/3BLXyzXnCvy1PJv2LG2He8GABt0prLq2g
nnvJdtSbqgSeX8FTwtp421lhzey+pvsAn0fzY/eYGy5Wfwru8R0eTdCFbsOR042KF2nh1C5vE/G8
PUDRyBfpDNoy0SIdoGQmRABoyBCbWx73sQCoEFgJj4G349uOflB10ZEQIID92NK5qy9HsGCtZ5OK
OU+FRl7xJFtUvzNxWvJnE7DBnGhF3pCQUH1IGKTVjnYiLcNYdEGA7h1k4IUCPoHUmnbqI7GgmAeT
DTww37dYgRS7SSsOrmEFpThKU5guqxUBieiwqGGkXYdZK1tB6Q5Xeft1/Kp1jvIW/mjZbTjGvN0x
V3yvCPOOfNhJjWAyyzJo9vhP+1bbkhkmVVq3mPF68AH9EtNaf0V8Bo32vvYiODd1jZ/xBiIZfCP9
leyLD6Yyx8OFkUAPhHx5ezcQ7cRrQaHJROo7JwVeT4YQnEN635HVrWKtrXK3ubtuVA17H95peGnf
pEnpZ08GHHte2toW+aRCRJuinD5Yn7l/dNmrRzSjilD5LK5CwOuzptwAzmpWwhz425zzDeEC8Xri
VhNqZMHpFpeALh5xCWnK8aHTh9q3IzYJJbS9mB3W7QwzQT9FhTQ3w+JdWcaD9q0l4t0bAKhm5x62
h7rz0ArFoVFHBdyJ/kyu8+/CFSd6npd2SafOoWSp5MYddsiPW1XMYdsyti51id9M86sPfO3bAxvi
79VEsSVOAyLOGDWwtG8BvmLM+Hyjjxz411m+3w34C59xmqqhl05gSzhCkxGM0tGW06jSd1x8Fa8e
hmlK4MkA5jY8QW6utbXt4fV13YPaJzMY6z6CNxwNh29xK/ctwuqyFg9K9gazEMc+dnua/iAd9Ddh
vG5Dq4xYtBjt2d2tHLS+Y/sn8p8/i8DvtD9iOrxYYmai2Df9T4mjne2T7rcds/UZskigfag+hEn9
Z7RwGikXfDt8KVazytsLYYojGPrKK4XxENphmQTy5aDMLp9vvXCxnDX2eb9jQOT+V8RJkfZZnFHw
LRNOkW9y1aAJaR72GaFeqRrS0JwaiEHc5BXYNVHBzf0BGaZ7oNapAKXK0FII3uf5WA1GxclsmRml
Qje8UZrA/6oKXSO1zPWcSGxMGHifjmp/Xf/8UNY+QCIOSCWLurVC0pQXpTq0lqTSSfaMRuZ0GP5X
03Xd/BfABNsroz/TWUf4qUOc9G+ALJkldBT2K7p3zhzCaLmCikHvJ7aVzAE8X25NjYmpR2yZTPjo
/P5psDq8YkOm4W+qCZuKVmDgfkTJnMQLqQ9COBasJ7EmsPQ+9YpsjrKORNNNmOAc5067vydiZpaQ
XgMQeivQ+fwlW6jwAV3cfM/axYZmSjAGMYOlQqaNzUQkRUY6SsiHJfw7KvInJPMx59SCgZeUTV/k
utSD+MuwERhxy2Me1xkWE/6+MrrzzEG/Liw+n5KkpL5rvcH7mCTWYv78ByfaEGe8HptwY6RJCOE4
xHYGTCZC7U5lqXaFH8ZsnRajtOOK8F6MARP/gle0V7/61xo/slbocI8pLP1fHAm6bq3RIe88XoI8
8xRC56oJeuYwMmL/fT2wtJpeK+7LL0PsXDGV/Rgv6xsVpEX2Tj7UwDANRBtZ0QK2jwT6emN6HNXI
OvMNWMFPflprgdadVQNWTqPFqP2pxccLq/DXZegIDikHPpIjhIIAIB3o633gSg3b2MMwMz/uZBJi
pNTVv2pgmKcAOICE+I7d0TuAhp7w2LVBJsxxM2YaeqUemXTs2LbyM3G1vpJdpmo1RzgJ09h7fotv
dBNFmaXBsNHN1ZeNzJYUELIt2/bo5UwcO1MBXnL0BTsSDIFopAYFl1sB35XgkdUovt0x7RXtnx/a
VcytMTpEOH7pjVGoE7weEpOOywd9O/jjsc07zStKLztTI5mtuFuA0IZQBOzcMSrERl/lpLqNulXW
49dbGmUzif9IRVWoqCsjC3kZwUZdTd7/jtjFNf5ma/ba82Yf9ls+c+C9u7dgNZ+ZgX61nAualNma
gAvXV6upnmpGOqpiAkNiY71WmLPb3LTccceTtdJnP9oAmiQ+QtmF3xFsZVJoe361IFmUDCB9ELal
ueKRE9UsmLrCRDMsPtmZoZVuxhOa3veZO3UxG9EPri8UyKjwGeuKHJ+GUB4E+2wGqj+YSc5Ky8fE
cvGMvs38UwI9HmmVkZC9q4TkTQkd1U/GKGidrF+vNlFmnL/nWtYuaJX7x7rxL9hhdoZUOgCOrpwE
EORQHK8m0nBnloOxNQj3BmGNJmpvMGbLUuhMLt38twUBnjy72wc33VSMNE3GbZLHEHIKUYC3gGqZ
XgzNe4lD1aPiIIU/ohbhFpmIP6Zo/5xVW0SOJX/CkagJWL9JUSQGcaHjDddeamjohWR1OKPOQM1p
dtzCBt/9L5dIMxXtWc+u+KDHJ0WxCk2IXnXmujebayZCLWZxCztJpI8s7EEhvptttTgyX+dhhlYU
kMi6xPOEbuZDNoNkKuJsUxNri88deK3V7WkuQG3MG3pWkc7vjIWTjMic8RzmD9SfgFsWQt7O8lNN
1cWNl9qyth/Y8suP9VoqAZxUV60v8Swno+nZir7AHY5TWBUjyImpg5O0uC0ZBFYk6biC5I8Ri7Ib
nm8A2FCc9nJNWPZpJotNEuPH0TBgOKqdD6/z2hu8tGeslgUcam9TQAyS1iS+2MFEWXC5UQzmI0YM
lrVjIk71lu5qSIGX2AcIlfU0doc/fNCRP3Iz9Ty/8SCS3asRq40WSuOiARWX1E+qZWZvE2M4eHvo
4y6xnHOSURheLI1HokfJViMglXUZ9mbNzD9VP9bgN1IARDTn/xxZLMHGrceM9zZs62ZcP7A9jFDO
IROYg4cYEvANr4/QIijhiGYAVgMH/I6BWJwm9OwXa0IokkEr9sCtTy+OGdJ4LzowpRghh/4MsuFE
M7JsP/jHFBQKVtCVKe6CAG4dYa2D5SErdKo1u6YwDEySN2CGdRNvC9ouGkibCEkoYsrordGj78GH
fhhXiaOGvRM8nSM6+YmEhvx/e5Iecwi//nhwmcOSEjBRRHz1yZe11RRkm7oKm8QQT2txEOdnHmNM
OxiozOa5OTdXVyTBwIY9zkWT5ibvsH0gaCLb7b2N1+9yxNeX5Wpfls8AKIc/VxcRd0q1WB6xCSaW
2i2Sja8FkRJqquD3jGWJnrsOtC+xBQbX2SNoxoUo5bCIVk7Ju1WnFh2tt2oVTf7rANMHkbEkSMVt
m33zRbOe/Oeg2MCc+WWRRn0f7T2tdk8o2zzVm3PvWqmo7XOMURhEIdICZ7h1Z62NmlNFrlkSdBuE
rwvpgQnooxySiLim9pBD9AR/hIDzFOJ3uE0UK2oyDV2PB6kv4vJpuod+smiB+fAGCbrdl0rHJKpN
2Tfkas7sTCGcMBN35XW6UmKv5JxyiwCpTSPfX6Yc1r7SkKQK9qlvH9IWrzWAneJVsRfwSBmjKKiX
Q4vJFeqtcm98twycQBQ0E5fDtvyYCVCe/0RAVs50b7uBgmZnk7DILv0D+pMNYN0VOExXfLwztBPW
K99Gqa+ZzqtL3/BvDwqvffTMzwMwfLGg1CQ09+AYghz+nZHnmQ4yZV7saMPmSnG0ljYWzGjdO7VI
m0eN982l8eUAIiSUopA/OX+XrchdTsVtTePlz+eQUc9X0YgcaJ+SDB5ndg8SNKZN311QiI0mLpDc
RXL/fWZFO/9Pm6Jl2/JOn4qUgbWUhOu0RMmvfseXLMAE86GtyBOGURKusvXoeVfQAHtdSFqWSKO6
E5VKQD2Lnx2XeMtOU2Vy38d13TQD83gDOdmyJ1C2i63cde9XOmxgACGs97mxrLgLZCViQSn+Lu/+
jbEAOAwJKrDUC5NqIAFSCCwpTHrdcqORdUeEYP7KTZ8w9Basut3Al7JKJEU24rLvmJ8fRB/pxVMk
ScaPyDiYOhnZe4Tom39w45fdPtOj1dpYflqsVmiNBHWhcKd7wwI06hHL+oUdKCaWnoYwYuKk+kdI
AFCOA5Byx99/8mf2bsATkXVtkwUOJ8wNjfX03PTCD6/csnp949InRH8UW994guLYjxhcfuoGeJVW
Z/d2ahGKbagi8JXpJdU1k/7hzbHzt1tlN4mu/jDGxi80ggSNWgqNJ9/jLkvBLGLQ5tlus6nkVzaI
9uusYTtdixopnBNUAnUsO3ZOyUwHus7Acv/q+qLRJh+6ZrfVeRo/26GsS30Qh4D6oX5WM/JeTAo9
cJS8STzbmrY3X7bWETUFhEOVn86LXHp2AuS+ZUa0qyneifrzJyIJfb1VrV9HIGwmFSqvyoH+H7i0
xDoES78xVAw1M7m4pZ7XsebEvNlrpfcHtighfbFjTiIhOM7Gq/tavxl9ITwv1LV9kRuw6ZZcaOLs
O63vKEF1SHeMaRXoofW+udBJasoEdo0SB7ifxRz7uJuT8RN2sBi4pVNkDEpB1h30MVuIdNYVtLeK
ORvn+oQRLkdgJX7kTRAkcoSxDdPGVmjeo4Ub1Fx9Jg+8L11OTCUBAEbYKM6GqR4TUnqg9f9Z+vL/
WfgU+S4zQo+ckS/prED5IJWLdg2/R1V9iGB4JJ/DI1W82A5SqFbnk4dHXHZpCAWMc7qoRvNij/rf
1oNXk2taumOiEOMemw+AeWPEPgPdabhypvPGm7FHqkZq7xuiMWObLvTDA3yyFKVfDLqT1c1FbjsK
nVfztcho5K7V0KFTa6b76e34YtVCt393twF8MnUYbO2B6pMOG220/UbDgKZAssUp2QvedUCL3Cnn
0clBnnf2t1kwymH3Rtpd++2Yq2zn/E6c4o5e4CJg1iGm60XBlv5nYev4ZyqsQWVRQbJmNdP1TYsS
mb/psdwbNmgEqoGFiVIsx25yQWvmGBeaz4U6z5ncqPoR1ce0mrlwNnwi3Zs2k9ijJDBxe+IOyXw6
wl0zzQkGgF9tnBpFGo41cQrF3IakMAqBN6nX6W/vmyRyOx8cBlQUBTdk6sF5euvcpk9E+EOx1JuI
BBSy4EcIj6BLY6gvwAu1fBsjT64Df4DTO/pU07vzCp/HpgjnMW5DT/dqW142ckFBEB57MJelfffJ
wuNDh1nLaLY4gptCPn1/wnaHB/ZG7WEJSEVQnX//MTSo09+vvANkKwALmyTcMzUnEZZIweb9cVOq
rsuhQhAWDuRkapiHuicMvoxsQl2arGLIbFuo6uCERitkvGmDoBF8MuMZbVUiiU7aBDJevZgys9aZ
PHKRs/5d1V/pvd1kv/8vjQ1FbcGj6qeSa6N9LXxYqRaZCeW0w9XIiz9NU7zHFJRuH7my2P800SJV
7hprb6ZFICse4GyVxEgUdy6+YjChPMFrDxngJRuj7xrGQpFYoDXdv3DeEvG+OpupqpTibVA6kB2e
Zm4kH/6WzAC0Kh9BFS82ulEXv4LZaV/b+ZJa5nSY88yopbNRx5+IJoucdWvmPwUiE39BZoq4bbaW
e1GmztpzGCyK6wiwmf7t/HL3lWBgbmDau1EAi/xwohgcaaFe2ChlvAl0W96oN+SktSHLrIxDRWpA
ntq8zJdlFAPfzVyFuXjBfg68NJr6mcklMDOrP9Pcg2ul0zo6N62azQQNR81xFt5U4WBn2H5HZ6Al
g4kNhJvRiAlyltn9l21MEc2v2IGJaYqF33PvBRDna7WN+D1QjWb4FnUI/VoQLxGIYsYjZ1HFGHDX
jxAX7LW2rUbTMJksgZ1iSmx9pryJELUSOFJS5hvoqtbQzRFmubF5+0hvknH4t3SDCym0j1pEf+vl
8oGx7eVkRhqOFgoY8CPYIQyKIie6KVJgVRhBG0p8GQgjabMkqXEP8I+W1LilfRMsg/xrY05vOyYP
wITnclBF0hly17OlPAIEM9k2G6KrbxEAsvkRqoxaM3VGRIYAnxkDAdXU1h2gqqLciThk5sA7dsNz
5+0scbBYLKIzQogxycLiAMdIMSRBXrVRXc6HCHlwwGncINRWGccb4GtB4zeFtE02DaYQjgAD7I32
mcMy0O/ufFotm5SdG/sVoZIOgqqijWV6Y/1qCUyBzjnglYnvRdTje9BxIiYBoZxAIFTXUmHMX+ws
7Unsdt2P5EpEd12/1IJ+wBOl0GB2UB4xcL0RbSc9F1X4CjGUoxs8+A4SxWUFRPAEgqbmlYKG9Dlm
YVjvvi3QXGtrYaoLERRPqs6EYSjVweu/5jXpVP08D2/p9MQRMbTz0wt6z9Wwwpcz1kEkqbA9vu4w
FA5LKCXUt6V2I63C8JCvrJiwt3xjoIIOA+dLZvqrPS8d8LYGD5EFEiTXt0LBHDKGPDGWZF39rCqx
zKEaFpw2Mgp63GSHt+IwmEgDW8ikUn7eLSILHnIPm5lz7SNLlxzwBrg0vhqFnAN4KX4haeE6TmMH
effEFLjKftt5C9vAx13pFgO4w+5UH4HtYYHGgawLSgpNBQCni/QxpfmgwYN65aRthP47/hmew/C3
8BkJQ+J++EcEuaxhr+COopQ3z2MVar1zlLd3UTvi8CB5Xyo9M0akMudYqC281ddu412PiBii6SZB
h30DrDQcvAYpprRFi1mD5QT0qq14C7ec4JTuUkgUPTPKqLg7e/e+tbYRt3Q/o5oaDNWldULgKEr2
hEncqH1ER+X27KooGni91qDOUw1+dqepFeRp2gPt0Aa1lvoF+qdww3q8M0kVdhrAay2YrmXVwaI0
vmEuavuXAd+UfzsxAvYKTltEGngsOF0HwPjcpGMNvOJIyvlnjDv/zRrsiJRbHfsZWNayH98Jkdkl
k9ix7hMIXBmU9BhyEjS5GRiETivxZDV+KgcBUg+ekyN1QuOQ2ZREmfU1CP8I37iVkXIopE1YFqTQ
Ur8KVw2S0VE0mGT3pLTbOgcGJt01ufy0acejOvfLejVawqv6hXktzTG2//IS0fFBPF9kMTt+5gQH
Z06jH74ISKGelKfUIxPZxAYb6DlzNhV/8fuZkRJUWhU/5exhpxmCqKMZuVGzPMOYLKHZdiGXDqsM
aeNTAp55+yyZJsx6QhmEQXWqgDDfzfcYQ03YwxwNSUXWhhH6owtv7X/Ea6jRC3Kyro8uZnRsJuUl
v1xrEORro4taEwHerRJPlVfi9ZZRbuiXM2FXV3rQlOxYSbFv5sfrf2L44da73Fp/m2j9Gh4MYb4r
yoAZpXdHDjxvHoJehQo0Moo4a9aikw8oUGhezY1UidGCrpMtfgS42iDZTE+0j8saT3o0Xt0GL3mT
FRP9gyEema/ibEbSWK7FJPSSVc8Ulf7KzXla8iWZgGZg0hLArIAMqlWUb0cEWqARh8bFINBdzvkh
+H6JRiopTbwjfcaswTtAKxQcSoD1XRMv0J89EG0o2aFa1ofv5+fadX4E862Wp2ydjmH3Wr4lqU2J
eD4hh/I57kgEvUijOILR/KrLuMoaZ0Nwo8ic9D7QCXfCFrbXlDS0Wti6euMNNUFlGBiHof0P95lS
eAX6CqpO3QCcgWpbHgwMc0wdwU1ShoBqUNRh4UBuMx1ZCeL+s68uMDmL29T2gVqx3j0/u5GBAoiX
iRVL30jX0KyYI4lAVsJ96pmg10r7EAw65YtJln3KywcKK16koaRsyJs/PDJcbX47g9jCfGknTtdN
PWFzwfzsADByD07Ii16VhctnCEKf9LUiXVSy0hzbrWnzznwSr1fVssUcGLCXjn64jNIoF2rbSOlJ
pDUIJaHPcySyXInd8RPBqFdALoiifpBdUGrvFQQIyX/6t6MMZnwXl8xmnWaaNMDEH2N8KFL+T4Sq
MP4tmMtj/EMJZfNn7YyiYcjNH/+yuFsQqtEOjSudRK0rI/WMCiGh3zAv6DueYlTbJMxlwq/msHNZ
qTZyYdq7hcqI26AH7rLddXXSXC1+r+VdgFQsGsbQFGiusoA+TRFuYsuGTzPcEBaRVZAdiKoB7PDL
KLTObvYGtPfEcFIF22K057ktFm5+5gJ00w5soJdN14q2eK2uJOi2YV3Zs9ZxMd3o8I2CVAnREs6t
61jPUTTXzMkYS9Uq9ORpm0AKAj4nSHwZ0BgL0Z7ywDnOkl8JBhVT4ChxL93KcnSgftSqMTDBBIuz
vv9o5gYIkePGh9xFQcQgySHhUaeg+Q/rrcr/3zOMJBbAiD4Y26e2Zu49EyiI/Qe6QEvTsoI5VDwF
unL3OjijKtFQC7RBkWFtJFoO3X4k+5rEJmBqTIOHD/G9i4yjnG2/MVA6y40LTqXiWN5NE/uHwPxK
Lu+WxyulvGwO38oW3ovp1RyhZhneH8v7KJosT8/gqDlQq+cy4EmXx1rGr/UrqhCpuepdKY9CDPlo
o07UzrAziFdB0BmQFz2vxsOFMtqo6yVkwpPK6TCznrl32RsQUuoGRFv6MEZojDnpxHP6zy2qiijN
jrpUpp8oLYRJCjh26jlujuo5iRtxulRqRRj4wcuIGArcrB5bSXQqRhQ2It7l1KJEIDl/ICAjMx/N
/NA9QdQwbsGj1U7Hypmvc0MKBMnS3frM2EW9XZUqcioc+gDmEKROUc/18eEX2zKvbO6V0305cwhp
aCUxVi+afLcVCSM8kJvXjW16RkqpI46b08oArYK4b6iErIOpbT4KY8RyRvOVAU3KNN3P+qF0Or4A
4LRtiYr3jbnPKGx/vzAK1sSeXnRSvjOYNf7SvPwK/OD/K7RbDJ/cJKqKCgWwUoWsd02KffNS5tWH
6U0riFLMXhTuyLS0R6N1TSxKwNOky9noymM2SxDwRIEqwtvKmddNk8UJCO19Y+mzB6raNNYTDDOd
GLobSXXVz7hnwwxTMTLhFaJDGnJ0B8FQXfZtH6SGmamr+mJMlUwhd6sNJlVyksuu+AzyYuRO0uKy
XanPDhykNKictl8WfoIWLWGBjbVczrKpkJcbFJVkvW3ot81l9vVJOAbbr+Pjvky4G8Y3nXajYRk7
niHcLomzv/bjxRQfkhg5N868yHqIoZ6jNUIWVZ3V2VU0mkAQkqTDsk8fP/hINm6RGYlezPp7Lha+
f7/5UQPkl9S+TuninzcW2xgbSqEQTak1WVYm9PXueOMZsUT+35uMkR9hqktkNmI5Bo5T/D+XZA62
opBdfOwSixV3f6mdcKOZvJLmXGmWn/8LPwFp5256rgEQcssltw1QEKSNRXZw2GulrTreUppOUvEp
oY/J0bICfavJbA3NaENnpNBWSvybx1ooK/tvbGDeOt+SrM1Jov9O0cPlFOIr4pBZ7gaxL5NF0Met
OltjUG+4TGerte7+GV6g01WcL3GUz6F/t95lJigcPGtLxEWq6DbTLb0mNy8eoaOwuL1Gt4NH7j5O
vahLVwT7DRD53lrvhQJF0gN26Mx61/h6xS40ZAQ52rWKHR76iqKAV8OJ51R27lXoo+2gE9wRQYvl
UREJ2YkS2ENRyW81zx84JVg6onPVBGwol5v1X80jkOuBr6ytfLA3B+R10ZJMdZN5Lq3Sr1+pDBCx
kL9ZEvoc98rHe1MmWjlP7dLbzsTC/e/2b3TLKes2yAZSOHMSrX+i0GNF9e9IvhLenD7a8vcKHt0X
sfh9WzFgC0mzp71NF6tuBfSKcpCo97WnIqlwu6J+kiwIZmu/DVG5cbkJMfaXdkx5Xv+/ewHSh7HH
9b7tac802xt54XdT6fncQEnhEHIUogd5kKAFGoDRXigJ1ijdZ0yegc6T8Qxl6aOsUa04s7YfVZpD
fFPT9OF4XAAC7qDlEmob+X/trVtKCmSN6MMqY5p0Ywr3ZXWnFpBH4keB8HUonug/LMgU0DRVyoFm
KjiMBpDGlJ6wo5upSeJL6bkYg8bz3Y6ciO9byO4kr9HdwWhjbn6J1CefRKDziN9HxEOb+AU2C2Ox
EJvb/bmIYFetH78WumwJlXnet2Mlz/r7EoRoiePx5D94PBt4sJuxP6CsSqpqNqco8LLhRJ6GJIvm
C7CjIXQZQsZ0VBH6AbiWuQ0uWDirpeOC8U8sCESmhImiv4E1glLDGmyA00vJrosBr7jg62mLB6/m
4S3K6m46GXRWxtsSoWkM0+AOnssRrzaUzMo2s5DSwkws7o5UNFD+AFdUFfXvxpS+E6WSFM3b9GDY
97rT/j9IPrXn8LTyoxQY9DvKRETg33Kn/Dry60VW19nLYvrBdv0uIeTrt2EjKeD3C1QAq4rJ0cde
qsMW15U0wRtIkpqblm93He7qyTZN/fkkMadAZqcgGwDVecKS78LrWdta//JzqEDYq7QEqSSs676r
01Ur2TiXCjDwBkQ88HJbhBYfOIAp0USTXoVTTMMJVUi6dCmRGSbaRiLMU3ehcZrUBwWiQH4f2s4x
+Tn0Q+sh1X64Iu+ppNu8uM+PyITETFOezXEGxVtKvOGIcas9AZcOHEXDpG/gtim9LHTELyTNtNET
lq4DZyGEqQ4HJX2ITqk+lqb0soXY6vonIsjUUxKu2wEGXqmwmhk6mp7UtRN+zOXi9voU3ViyY9t1
ajaUYcIx9SdZwhWFyIkIKTCxoB6j/0LWrbRlpXKHh/NF3lsAfDszzyJEzpM5iekGXz3fhCpBZd+u
IZMpMEXCJ+mytMMyiCXHQfVeBk/LmFbpQ7Cn4zt3O9jbby9G7kaJ93+Q5DuiufgoNKDXGnPE6UMj
GaMlQj+f1Fgz4w8Rj5Z3kDXHCH3IKbOeR+ndL0BszBpWM14lFRwTFr2hWbCLt28/2vDWw9WbIovv
z0iQORPifpE1MgU+zi/U+qEofp9c6sSF2j3G0s1frwkjlNbZ1b1Ou27IPj3bBcS4IaF5GHs6ajan
cg+0cmFH33NrzLNRCW0zES+0f3lrFPxwrunQORVp5SafP5FTREx4Q5YpQeV9qyDcF/fT4LpGiMAr
XQ9xPG5mmhx7y7AwDsu8aVqPsfR+nTHkizLDQe+R5fIJBbbfSVkd+3roUjsJPZM2nRwWlGkJ5OHr
TO8el6uwAnU1ZhAHIYu1RB/T5xLjk17Al3E+LyU84uODQHi3SEsSZoSAcuUWp6N6/evkCRvOfL7K
mhQna/B7kqPpuRw8AwCAlk94M4CVVBP8nCflEgMsmWLmNsH9lT5EN4Z1Ybxr0Au0zcvf5eHPGJwL
L+YbO6dbybDJ4r+Z7wD1aS0Ur9/fmxn2R/1g5IyDcN59o3ODT57vQt8zIEDeM74VCHZN3Hhd+vX1
PID6zSqCetoLF7RY4dRLnnSj5q+MjWF4ZTGqDJiYDnLgf1reD0WroinQRPf+Era+a70vCiqlSxA4
IO03w2FctCyN+PgdcgvBJh9srVmO32f0oaxLmOSMdv5sThj5YCdnjV2mYNd17eVltG3M4HgIatm1
eBfQ0bQ/ski2FUCprU5sBrhHqrTs6wqhe9Aa7Czjb+r3xtGI7MhOYqF89y+RxT1veuoVoB3H0mf1
m6L+G3K6I9T3xJXd9hxbTzPN5ivhNx/OdN+paoXH/RSQJmkHEE0wR3SbaskD+CxmsuS07jNC/yyh
c56yh3TcrHPDkHjjyB479SYcBB4xgrMTazDp+BmmOY3V0GXLvsvURbTmR3BDdG14jnghB/xO1rEc
cs9CY3mVbHUNMahSPsUai+HsELdw7JHiGHBbnh559jaizOq5xFxgBAqfrwrrTLvRyLAuRSeGTt/4
Qg1mgorIC15awjjUu49PBVuKMP3tLIi7HQKZjPWCmb/qvOuakdi2LR2s2E3K/Su7BJyxowudJGeV
nYslTLw3JqJzRQ3rxRitcBcSiXrllREpRycfad/5s1yf1/fFK127J/C0hA+sO1uu0e75Qv2V6i3T
5bz+SNoJWCk6j+feTZYdc+97Gig9baGfkmnh+L1Y7wMBbWv7qWNxuQ9t+DsDvtMMB7LqyTTXHCFX
nRPRrIYVpXlVtmd7pGyiuON3zeEAogT5skGZLU0rE1gB7hdkU2pBwC60Daatyi9m/7DCUPZogNEj
qv5+YvJf/wnSmC8xbl2+OOmzj3qM9UT/MLnczqB40XNw+0dZQqzUQhNyTSoMmmD8w6izjmbEDnXc
aWLzz8f/cPkt8BhMReHlxdYLkPOA22zzdSwXY7pAPpS/2OOgTzL3ADQsHEQIEueyCc8yHbcyfI2v
uTAqA5m82GKj6xHUi8457fOiSYLbof0VDM+Ouh019lI+kbl7K6+OEg0aofNEmeYcoE5IbnOYUSEl
GybUFej9gbWefP/pLTWyPhZPJVJ4WQvAnZ6O+StY3qShI7/HmvwKN7Bifz34BTXbUndpCsmKD67t
E79bR6Csi6Z0i7nalQLDjeYFGi9o9tKEd1Q2CpqMOjhPn7/NwMUcy3NJfoB1Wi4ovOtufcPZEGHN
zdk0/mp+0y08AYHwbuqb3/urTqG1Azisq+bNgLEK/UrMURG5R/s43fWEkyZ0Vo+Yx3IMSSYZ90hx
uIfeAQEaayYpfWSnfz8R7soCReRgV6YFUcRipXcfNccqAgAnCoLUnPQBiuh6c9esYUUBOJMmJ2xC
efqK1uDtkpR8pg1t6EDxyctLqmGvDOSaCyq5kiafIc9WAQJzbUs8CC6rj7VjOoSWP5JuF4VfE5XE
/A54KQ1eHCHsZAlTROt2yIdUYSz7UgCRm5Gy63TV/A82b141lDbZpgingKHDOBlqOFkTJQcKCrXm
6N2Ll2XlTL3dns5ONHRe309HuXBFIdkVcB7Junllw/VObytN6X/BWVdtv/BRaBkeKWq0Qj01hifH
eNot5pnzklb52x3DK9JXHEtXXhIU+9V/DvfTVUoJ/1R/DlySp2du3sVP9s0hmSOBuZFgDy2tWuyl
/ApCUuhMs0JMdTVEuoAKe+92Izuk+rUnVf1QDQ0m1nBnDC/+Nx3Or6naTcu6jhquBsinYacgisdo
CVu0W063o4iCyfnTsCr3Gyaoaa0SdcTIgxLpDgNOqZZcyTVLywt/28RYo7rDeRF3QtzTOUEViNsH
AG4WDcsKCgVqYzdh24rjnI+K5YhZ1I2jbSUbmNGGIJ0LT+BD3f25jaP0jGbuH/jd0daJLM/yqiHM
2ImYHEDID59YABCc8lavfUsytzep4V1dqZQf3dtS9V2o7pfTEz4Seu0XyJMcFeMha++yUyhg6k0Q
RSsf6FEIROFt5TqJs+UQBnMrLUxRsP4+ltRrpFJ1OCbGrDiri0F8oeSa88RNvmZm02CvoHaaeA2L
dbMX6RgOefsHJ9dIxU8MaHny7r+lBewQmdD+y6BG3L/sRY4TwF8HjSxuKaDk4YUfItaJUeE3EF92
AvGiqKFxPvcQ/uLZyzhCYPiPqQOG3Bl0bwKJsxfB41u6UHETLz3+vOdvvV8iyRFdOyM6g1oujJAR
f+Jm3AbTQ3KV39jrDkvR7Kfu+xh9I63xLQooCMyZwReiesESIKLBb4jfyM8Dtat/oMfUKAepOdCN
bKdOhEIf6iQaqhOPXSQ9kzmXYrQVoQIFpkRQxSrRo7Rdu5pOtYq1gqPGhFEH/3YAjfzcdb/rV12y
swwaSwK3POAnDN1wS6G1Cibmov/LPWelaNDXwPJdsWqyHCzEsX7F+g1wW+nhEgekbLHfbj1pWlNv
vbX0PE0zxWsSNlrLJlk6tL9Jdqa0rsnpFKVrILrtShrbiXMxWj/f76H+lYfjq6AUPYgID3gZUAsY
pCHq+FFSfq+w4lvU+rK0OGwGun5Pv7Ip1A+iwPis69DJXvdIqKRMnHwOTumiZJtQGUyKVoGrhfNS
yNTIb89YOrlnsaVkQf83iNoLC3d6ffZSd82t9/oh0SsmtK5/QIgHCrCc8P73KuICPsqU2E4CGaH+
qV/atki6dYQ/wNBBniQ5n32yxBaliTeVzrFSV1GPZp45aFJncFzvBJzzL1ei64ZCqeILHyo/kQUI
cGE7e84jWxaqhb5nxJTbpL9EEwo80fh0FqpbwBWYWyiqGQWGscxi2lIW+jAVbkxnjG50emJB7WS7
L8OjQPVuTCrjpKJNLOXI2WeFyrD80/NDZrireE1r1YnNLZ6A4jd0+sL2B4jk2LwI6QmDcv9E/P2g
/mTHc2Y6LN87NlVu8w/fGzGwVmmYNb5JnejQ1dKhOWEi54a3TWvz2XpMOxgfbi6pfWrL4d9Stui4
HF6C/hdBnzG/uwcmbU2QyM1o4Ix2kIUIsgW4QfC/I6U9spFkFmbrpUhlJOHPef1Pnb5pORk8rPGe
6iyZngWEeTIj0YU7e2POFNcYbvE8X0lYexa7EHDZhOdH9oxpWG07rq5qwcUOtcOWgGthH9R9gDk5
BjrwvJoh17NwUOWR52iVsoiVL8HX4eIkGUCdZw6h6n4inoOgzEivSiQCxomKUbKexSqyX9rNmPpH
49vUq1qCd8HYQVyiOkPoWSdNsgj9WMNkN7dSIg6CZnr6EtD6ZH4oEsZiO8u8ogqpPa0bEC7uNoxj
4vC25IzuVMyLTPgwC+2QmtnNUYJhS8sOteGFmIJ0qMhY7WijRCIKTEOT5q5Y7dq+S3H7bzJWlIGY
5lq2IZHRVRh29OdX0o/m8rxzCAE6kOnetRumwakFs5bXMok58cyfAzOrtJRuD93Y5O14+KJRUXil
ZImoQN38RCs5/iPEYC3i5tMC8YfYJmQ6KlJqcIYa/Gbvh+5a4CfFzusAGfReCz//TuEXa3/otohj
2ZmStCqVK8/Un0Wlq2bKjtiSEZN/oxkma0xir91hxHGkV/iBbGSNW8h/PyuI3AGtXOuPF1S71cRT
dvSnL8+xQIO6Z3csJS4L4/yZPMORfP4LxUzxwJzfLiOk4EfOWi4EUzol4pE8cuKs8CZ4U0IUL8U1
WeCot9DbGUtq2Tde5GP5jfUWfLzjvl0q6IP1oHKkvHa9N9YpaNdkogfYnNduvAUVQSSAoqCNnRMr
c0btTv88Ogs3sxCTMKqmR8JjW+FleTo9fr1LqjP6SHavhi8fU/oDwia2ABlMKJST5Gg/i3PLBX8Q
GGIGlgdmq2IaTFOAHPk74ChW8BTeYMQKyonb5M9wcAI2+/CqfvDAZoymvGbokUjXSeFAiW/Jg4Bf
XyBFNECiGP3XyJdt4yX+H57Zq6VYkxTAMs4Sy1jgZuNdQ34pmttX9Aessagg9oHsI3fYvvdu9Fxg
x4eW1AG80Jm92n0IMwCGX/tnOu4pngL/AVeOH9kzaT11fJ+PU3PN4LPtIaZ1UZeNtOKpBgjFryO0
6RjCF3i5/qIHwGtaPCTwuIAKH6BtT+P+DVvXuHpJfNi19cX4/gk+Zyx7eGOP0GlGbmKyImhaul6y
RKjTuw1wmwtqcDyR8rqDi1NXjBXv8AzkfYZhUtturoZAuHBo/8n/vTiGuS8B2H9r4cqzCZeAMt0j
mZFyiQ1ndi2WmSVYvW3Vu9kCHhdQZpW7QmKHaVZt5Rhi/SP2Jwl1VzkSao3alKPWDmXtmMuCVdGb
45+mpHOvQIYMLyRFw8ItzhXd6i3Oaq6/9FFYusEMVjUh1SZlpq3/A530oyA995ccl41tJtgIvQEl
2KtcRwNAiwFRCu5Q/JAen15rT5AIndfxq9SeRL0Om2ELPerVT1r2A3l5o4HfaZfhjVmcZM8kjn/X
1cf4X6WVpbot6P+lu0//p6q3tfas3tqiHNp/IyDBctO4Qs4Q8B25KE568VuJBaMbWM9QLa4zG1lU
fYuwtQi6+2L5P38R4kVpNKJaxJ+8uB8A2Pq5VPxzT160nS6vgEKpqWcKwAmJPrw4eb95gk2Nc9KB
SJET6nt6dPAcZGlZ02X3MCDN8Fr9zSgm1FfrRYBC07VYegYbOFqDOuO9zkWF/Na6E7SyBDd4/q0Y
e3cTAMI+pU87Qco6hPyQobrbC0ou9h9zOIS/vaNJz/Ut/5KUsTwq8wxMd7Sp9tmdqUj3wQ2bAMYt
8fzI+C0snwijotrWhY732gKW5rr2uafLcWrHUOGIK0gsZy6DCGEzPl6x+R0B89PQzBLjcbqejMd7
LLvIlrTvqGOLv/kQot4PAkqDcX6ou9hDQpRvyDJDxD28jFSgJZjPk9e9bS2QxE9u9FdOxO6ReXxZ
quY0TMd3Ti0EGZi8Bx8I1g3vpFkkWRDN52Bd22e+PHYzvhdYjK3akz5oA+frkCTPlvcwrLay0eTn
LMahg6ZLyZd/yxD1MwMHtW3JH2MfjcHeZPIZJR9+K60CaZu6emlL96V/+TWEf7JMsDrTuQCmxTcw
f8oOKP/KSw2PbPcJq4Neg0OkoiQM6f/2YPMR7l2/yx3oDMyyT13rPWpDoDZQ7UeW9mTkQ0Z98qkG
cbg41r56Wz81+mYrnQW9TkEoSNJf2RL6b3zjcAX4oy8K4irFn0rPfYkxWcMp3UBIqkPm6bnT53e4
kpcKq9orIW5lsevlWD73Itlv+ENGQULKsHDEo+59TVusFmTCtzbITxi7bWL6W8n/B2UuxzuxpXSX
BofAD5rcOp+pb0STfCnpPEAbnoz0+LSYsrDPE+8im5pZtGgHnMyld5TT9ihRXG+bnKxmWyaFmcsb
gVaa1uIAMQ6yg9zZYTn6VgRBi1EtkdWqJZ7q+xJJPcQKX20GMeUV6pGN/UATBQ/RV+vialWw0gTV
0x1PjYzEZl1mUP3cbFAAH1qiNv49ffW5EWtgZ/FpWkxlf77O+n4n/t3TERSbUe9JzNoXm6lq9hwR
1SGV5JFU618NuFX5hnOfjtBzdgZAr20xNSAS0wf2dS6SYJYu06hQ+udSktQWNOrmAGFs63BE338z
uvJzHDnMRSa/9QWWIJFCKNEiKNMYlUEJOZkVmu1SHedPU2dCv3FHyNeT6tx7D3S+GCMw3CJ6aht0
8UtjOXvWM3EIVcGMj5u65EzOc/L851ivgBB+KBTexX1mJHE1S38C3oN94Vodi21IvAh5UbLhX2hF
peCcDU/43EVHqnH5/VpOKVMaPRwrGLfoAxYAgb+0trofiUQGsWz40fxKflOWlu2GM+LqMvuNGGVM
hGeZ5ui5/kS1/I6DcSTJnfyp1VfWWX9Nt+KeFBDK9aLwkFrNBmtzPdlzIZZcFiYVY9ZXj7VAmrcb
Ie4JKwsgwyjyVOWieBzWG2lvfuU2cIN90UQ21kcyR+bhVTYdFTMbKKWiNpFQFMSdrRWEuN1Yt4A9
8zVTAFCuqNud+WRIuYpvX8A+gaKgYfGh0GNy0+nvaD7b1U9NQrX1+Qr6ufRNextfXwPpcTnp4x42
EP2SwQtLDmwoXTlOfb/koERDJlz60tiB+Y4GwSL73zIpADJZY6XGJJE+VKh8bl9mbpbAmxMaJd9q
Yd7iHRkefaR2cHZr1L6uMdbFGT7YBHdt5z0kNPEwzjvq4td7KqFrKu2vTpPJNn7GiACiTcb8/Fn2
A4AVyYG2cByEcpPqWAKP6+O6EYoibddAhfpI9Ql3X+c816K+1On6u7Bo9dbLIgUiOHNkX5YLB3JA
I3W+WxXkcqF2PhsQJmREMMzMzzxAMGviAaN0ltP2SLTIF9LYNr3y/3OTK5qY5fhkXwPJNxqpeXhr
zukz9rrqBwqhuE9ftbIAIZJ9kbfKHw61TvwMd1hxMWupw8bwHU0SLa2n2A1kuYaWYbhZcPm4kVq3
R3zKr0aHmoH6901yPf9jFAMnKjREuOy7C3Ai6AcLDMLHXqV2JxRBhOe0AbcSNcbZkafnFpeUkMBO
oICgGQPJLuV8277r9jQXpTqpgX0BFuiYX6JJEQn3frCUG9ZBkvv8Urlg8cy6grLZGynYgTJV6xTJ
0N8an61awJrmi7YO5ceKz2sUpnEr/pFuz71yhizHRj77Bgkn2uYb7f+53ytvrALFpnvHkUwu3JFM
3sk/PEGSz34jr0kpJsaLKs6kM06BlfA3FVuHJyMhOSbitm7WBQSom1Y/WRSCcsIEvItEivvTyDcc
a5JeQphRFGq5o4JFJwraLOc+bo4z5th0n1KdtsyjMTcKxltBhOsVBp6mxDPX8jz0WgVhfhYEni7e
94QW/eksh8K8Swz7r7FPgimgoLvBwQTIUO6I5ldtg84ABuMrnOQ1fbV+n0MT6WHQ/v48siej/43n
2zGt81uUUkj9Ei9qzfCAy4UVH5WdEq8jt4zNkGbPP4jHKL2OetWzDxHUyqaLTqa0Vjofm6VANakK
pH3wObtgjgUCWDWNzvmJQ4cbVGeu9PcO2VWYyNY1uATGbPPa0WFPj65qnZFwsjZz+mmuanZTWdTU
ad4X14Dcscb2LIP7c/QIhaUR7bVuIqgZ8xkt0HsRlOZlJMhon2uH4QWZ+e82a12pt8GapZEWijXb
JIEuYUI4sX004PZu6vclYJiogNdMxzaXm12/i6LrKzJPr9aOKoeA8MvjSOVBSDNZ7dzNCuY9NvHr
GNJMxFZEMqka6iFWriMCAyMg5UrnyOI7XlVj+FwTImtbsp+bUZ/Si1w4eZpnrRQGqOl3aTRbg3gX
HQdne1L7X3t9OBu0QGMT5iTWAElzA+zuMAebuZU3+sRVJeS/hpwYOBDmJJaoYw3v9znI6cLwYNco
waPQswo14HfxsfL7J3zcIk6Rjns+dVtALPc3YQzLkuRfTfyco0pEHfgFpUJ9Nc6wjdpaeG08SW8/
sRoPj4LqhOa0WUgD6ErA8AioALdsGSCtRU10MCiFcj+5evD0/Yq5fXnSK+bU8RENlsApqqcnVyXR
6Sseajd3jgUAQURI5y/U9bqIgLrykbYa7WLg0U/C4BgBmWcxmXfzlOEYtCk3k4PDpbLHglReUE/j
cBLb25Wb2o2SvHqaaf/6Ep3zdZQszf1uH31cj7W00Xct4uVcuuq0IA4hNmPr51zm9bICCr5wcVoI
Mbh0ILj5eqSmVcXSLxo4P8u5Hvg6yiYC9I41IuYPnIGYflKyj7Nzr+hsmzfbE+O8NbkPD9Pk0GPH
IhQf/ousRDNyiiFkg5HVRuh5tOSvsKVdKjbo3W/LSbEapcGyVleuKdCICi6GtS2xlP6em0QcG946
nM53eYeon0suxoMfjkkhQiG/Av71jZpln88APwchLAW+qOyUzNjTnQwDXtWZUaj3M9ngx2j43JSc
o5UBh+udvE3i5Y9uVz3scc2UHlivAIU8hrL5/H4GkIjXLpVN68hvYbrcgW565dSevijC4gJUE7WO
dIpstaA8mHhTWquoTX3vD5309ht4JuRmCdwuSF/h9GXTJJfzeRJFcGs6P7YtZWanyRxMa6V0FTd5
BzB+Llsb82Ijouazge1QQrwK6be843+xKzTKnuEynKC6W4lLW1Zw8sCEJGv7sgXcHI0hecSF64lT
DNNzTZoUIcc2QANnn+ahYs0p0/1buabDXxWomUyTgXlbiBNCCzUNAjT73mrxAKM1VoKqtaCoJQId
x27RnWRyGxmnilxBaKZzBAu0VHOfyzwW/yA/v2enDktscu3XUc5E3stfQL5viNxrn3acIIs6an3P
tCswFbo1H2gAGCOYFU3oY341dO9q+eTwXkUZSZlL7MgP7UqLEFFiLjsqnxp+KxRsWR+9lyIy2d3X
Li4o+6pJUMwGPWTPdgZghILOMIWG1pwxoyka89JCJPcw/f2VMdK2OmAH8H3QSbx46rrAC3mYiAc4
vRgfE3TZYq2ngFP7PMH5tyevLCJyz2as33WselT97CJXZp+ED4DWRE1pZkn5dFEAo+H/f2QYuk3w
dUYgdwKGKw969FpBniNx+sLEk+pOhWIXacSykwM7b1LnbnWzw5nsDL/Bcr8WO00A8Bij7e5z6xsO
01h768Cxs8DUvPuYbUGX6S25cz1VptFUxYyXpWBbF4hI/YpNosKni5F2JqqoudnEi5Gkq2mmVGiH
QnZpnXdjKnbzY1AEK2szU22GRWsUgLV06GDYNZu8bgkqy5pyKS7PN1L+eWE1B2iELUVN7Je5kqBp
KWUfsaCtJc+u97bsshbiy8txofucGy6/Q9+OsbhQUH30awyLvNbuO74XhUmzHu4Slu/FOgrOn387
/yYg3PAIiU7uOICvJcFioaFs5UBlVu43Dmb9AsqQ7uhsVv8+A/eGW7382JM2LhQLIQVfouCRXfZp
fpJ1UY759GdGNhnDyAxMSrbtfdRHLO3ojo/DuuQ997nDXLhq3v4k9Mijv9aXJStroXVC3xC1UKUh
c27z5p4WSGNQXPlEVayGBTV+FzYUZu32jNujESuln0b7ISq7G6O7kZN8v0IqKbuivzOme2C5LxKT
iuoYPBJNc15bir1prTDyR8MjQgXWsPsvPtt2ca+RyHBYml4t8uukeKEfiRfUYuStbJku/dC1o7MP
syL6wq9xP+h4BNGWvnnmcZiw5vGUbkaBukRzQiLZyXl3+kLSAk2jf8KIj1cRfTioLa2NfaPwklYt
+cFIJ70eQALd/JfypQE8mfgg/qOpBVNLxUgiojMW+Lmm91ioSn3VJg+xxmjGoH6MNaslnmfr/+1L
Fi8lsIj4LrNswhOIKEgJU3+wP1t45/RXWbsHFdDjvPjDbkyZ42Ophpd6D0xmg7r2KDfMA39K20qO
FE4ySGyGWbVCJWrKOZJgQABZ/czS9udxU5uPgpvuEIb0XjJo0nKbb/LqhoLXUIhQzZl92djqXm48
0WyRFgCu0/OVS7tyTpWBvFCxRfW1KltcBltzITf9tyxz/cet9aKZ86UmHLcEYU9mptPm89Ck3wti
+ctGs7VFHaKZCCmsEnCl132yhaPRMpP6iqCTaFjwmk1OSmHJi8c4UGOQ2SZRe17kTP5pgn4Vgkcj
rFCZvn1fQM9k8ATG8ZcbX97Ogrfo670ZmA14rnFBfZUPxkjXj+A1y6Bn0GiU26jEPLLizh/f+anG
b/cIR/aWQru5yknIdZBmRUhHtVSRCmwo7aYaTcFn8bVThoobqT4kWWZrai69OWhCCGlqSb0cMEis
yqnoRaILCI6a8EWadw8+0f52Xy/6yZ1g/MEbM7HbbWnC0otqRxUAlm1vFQyFKuoIwgI0y47nrsSD
U+mjDHDRfbT+PpYYe/qNtd+PFs3uLBK47NYKyTho6hZxzSjKneMfcSTUjN9f+peuO5EQkH3jlJVe
7rM6coMebHaxmIs3ybKvAvNG5yuhNxAvMVHqQmAmyXPJ1Kv4iR/6wzikIsc6uEyAOuKw+/j/E5ps
dsfOjC3uZik4iv6oGFxFFDgD5teNRVuDhfjvO+lKUFQDIce1xJvs+L4XPcHQ8kC+F1rK3Dq8IWrz
4uiH7FjSPjEY5L6sNSGJfRQRMXzsulzoPTYAXHsSXI5TAM9uy2JteNzFUGXjwQf7audL6BJJdAKQ
2BN4pJQs2YoUatkbryjv/dUdaGh+NUz4NSduUHTQhywiEd/A24Xn75ZXFVhZ1VMNvafvNh/35LjL
a6bEXr96LlpdCBk0J8HnRQcM11d2YcM7u/aYERTiQD+ZdDn1crIcOLpTp8z0tKeQ4I9Ly9rqzXdi
N729syGuguJtdegd6zG/ZolOD8n8CG91AJ/rEyP4ECvB4LTFyjtUoC7D+KalcrufyXcp+2A2ygUS
dNiCeBPkFfIlxDL90CVc2V+vSuRDjI5doDsRFQwbYmleI84EqypafZdLPNhMB2xTxl26lMOefaQS
cJcWwFiekN/p39uAeVLs32dups0C/jUO3nvNo5mOVyf971SgWkPytPBpuU9qwXOddOP5UtqsoyGu
2BwXt/18qD8hi+ntAiyRSLEDlGPSMBY0mBCJXkh3KFcyn5Drqv+YPT9u6tc4F+KYtGxo7RnOPHrQ
+wuWGd8R6gkJIhsX9Ynfyaa6h6uNrSs8ggfyUVShRWRj+ZgGocoieIZRnZ8YBpA0NrAlHMU594uz
auV3lc5LDA7pfjDSckJCWmJ5kNYZuW1hRYWi8Aa6Yp0fgFeYE3EpSr695zHG1wShBub0jtCcolnJ
dr1UHImEdlkP3nwbLu+FWCqI+lLUoZ0hi5utLvVfvO7TGjp+/AXAuUbufPA2YJ+KpK4diAg7WdvO
PPheta/DErClCDphjQh/CBb5XwtJJm9HpxmiuePErWsELN/7Wo3tAPBCkt6ulEcmiL1c0H8MxAiF
TRMC0as+aOx8iz8ci0sV60jRI9NT+St8GY2zd0ji3OT5L5X+UvauAF/Y42Dit4oeYFx4zBnrxknc
k3gOHgltZCVakizfiKwNojWOuhZhS7ZF9vBtsWwHB8sLbCx6zxpxBeijI+IVSwCEAIsPErHrBScD
27QmNPgHeFSn7a2plO9SfKPOj8HTwgdQg+0xrkg1/tkmI0C36gCjIsDnktHJDuYi6xlijHWX+ez6
belKd+t2u7KKSPn0C6cZbi71bu1v/JFSsRGVMYKBfT8eHm1Pdj5QW10yVY/WzUZcp9MK43QA7GrF
9XQSlxl5sefwr3qhHpdpFImI6lvMj3XZS2URzPLMLqZqmDXL0kbi0QnrHf6DeI6OIXcTVgllSwT/
c2RrwBc+BAJIDS2t1z6OxfdBLFxLVWpUE4vlIgWpgsMHpusmISz4YhSFAG/Y6NVYz9v9CDn1MR4I
zyBrU/Qv/G2o0KJTV44EFXqzAHDXGOqnFEMHywYE5UlPvjKt63c5UTwv91F9kdELCgZB2+V3vsiM
iLZSNpqJh4gcOaG0xd6D6q047su2swKevk71T79VI/wyucoFGElGNv+xy4PiMrHu0mmQYD0EBfID
DGTkwvOjAJjSGjE4Kk2th8vPTwyMNaYU/QoljCS1TakTE9Mq5FGjJgV6l2idglUWPqUZBZQVFpyf
1CSLBFHWbk45y3tX87+RdnhoU148Ea+K4KECMt2uUUmlpVSv+N2/f1N2RvnlCJ1DSVCIfDsyu/Cd
iM+ppWVuTLfbR6mv+Xla+r0sIfOEcCAzv3N3ZLwBTVN+7UEGGk3FP3jiDOWYnQOfXZGjk7JFv9T1
VTdB00NCrYCPkYqvdNA6vOYvU6yOdlKJ9RalvX2Xcz2NjUGfegMGiRIwVlSidWU5YzvCGWi3nyhf
opoJQ/CnyoSc3I1xY8dxuDMHrdSwagoiZHxfB32TPWzAEZ7D3BlfszUAzS2vIT1FQ5KSqM9NwNIQ
Vy6Hiz+P22srzMiMa4p1593GEXWreJWYX7kVYm0GisHoOjMJiRqAoGycESrpKUsVMwLAgMOrHywX
rcCQEYVE4yibIvkr5swSMIEOG62J1nZJJ9k8NsLxfpL4A8O7fV2l858xy4wbnlDoqKPJ+WMjXip4
VXNylPRJAvfHNJtIHhHtHcAClx5jNd+JfxIx12RqIoXL7WU1ffiVgMY4ki6BJELW4Vor+O5WJ5XE
WqoMdSTDiFh3fZN3Dc0R/WznnPSUHd+JMZSqYyDQ9C/U+0HcQPeKkf6uar3M/bjPDQc3z5gzooQx
6Fu1WbSxBHoUZVYjjxluP/PQ7Ft4orBMPvU7xtifyAbdfY5XlUUIaDJNc6uR3gUDsUBi5fcTA1HB
RKLxEFxwHbhvT2kJbs1Q1PCnxkU0G9qXAGtGgPIJLqAZpiZrojkeYxNf8qw/9JVKOrlCHxYVfP9e
RAoE/q9L7lOA5cDt3Y+BDwokAFhA3LIduxipTHoN0L2YT152LLYcin8q0qZvh4IVbyqOpCPJXAaS
0UP6uAOi13xs8HDXG1OmY5ibTjGTSwTLrs5uiI1AyNo6S4fyrvyJ6hV0pRQ5HdhJseULbZbXoxft
jH8w3Li5cAuKw5EzL/3kjhWIHxBbhmoqr7enDWk2HyFUjce2F4eT+Ic3eynS7c4ruaidvO32GO8N
Z1Vcmk4vE+Th9wI077wmRSuqmG5p7Y5KYo8Kco/vRTM99+IemE9okyKCGaQCYMzRucA5a8xk7dhC
Fq7PAGGsnorlvntjuYN0M4AzJLApkzXY8DRAiusFncSKiitPbP/3vX2Ycit+/xhvvS3ADaVsPRpg
FMbEHipnaEiqVGwVPZGCreQYcFqIX0ReCBgKYL/LqMoG9VXM9v1QxAZDYvbEBpoPsZ2l7hatoeqa
YBdXgba5O3aAqAfB4RaNbYF0r+jT7cdhzLXbc2yKrFCl2lfSYWs7JFHTH3BZ/ekMrr0FI2dLvlOZ
gmQEaH0aD+hegM4/bhU6+9uIPyTxBsIaf8W5fLVG+AeRiiDQO7FukbNC7H7hQyHaJS9DLD1XVn2g
yg1dtO5puNzKW4/kReTj7+Q8eCXTkU378elMiwNz8krvDw9F7IW7kASCV2HhhhWyI6FexB6aTShB
EJh5oCjSI3+6dml9cAW3d1kl05UnF/7R/SusAeec1STV1x2evyo90BRrG7909VRjlOaRjFEt46jI
DWkbJF0dXGRcN7xCst1ueBndBGFTpIzxE4om+JCrP09/SrMvM3600Ho+FRZdVZeoYc5FqmY+rsKp
TEcTxltJ8zyMyHSeKhMky5ZWncY3452sHgqULp57H4Eauq+GRveA10Ga0naPVwD6TXKD8hjMmf9K
ZytdQQZkK50VWAngiLL3uGvy8IlJeCJahbEB42pr/0TmsUY5oSwF+3RKmZqt9vUAZdgJNvR6V6pG
v3FUwl8qknHeSNKKi1B6Gnwa8LiWmiqmwlfX2t8SOYoV0Nca/c8LFA89lVS4RZwlOe6pC/i/t7pL
Nxrc04Gx9/33aZvQ3VwSzAEmzTul/DVtAC6i0dmh9FQlQKpGcV1xShKQ7P9xxNVdyPELs3dhsNKR
Sefc15y+pX/3Qt9O4JCR/xAAoEkI7FdxK/RC0crCqrtj3vUG1LSBOltoLTK/DGHfYDLP9ocVJL+I
aUIV80hGrT8ad4BzjHdqdWjhw2pkC/+ZPhqzCr9UUWPs3em2IxH181KJKnzUKX8XeyH6urTibaI5
WyZ18x1T+E0x1M2Xst08sVJFUxKy9syraGa6XMTlxiF8DFPfwUAPW4oScBxfHXMdCnSK4Z61FCa5
chXEWxIFUTTrL57xxBBR9THG2x2e8BAApdEg3DeU6wgMpNYvbLdNt+dKpUgiBlKXY5mxpygIlHyI
C1MLTiEKJQpxu/ant9ahpYhusdUdy0i+NvWjIatwDuWhtQd7m4LZd05aaHbNf8F768nIaS3UEI6E
LvT3VD5T/NNljhgGGKppaX+PmEzbgHj8co6935YTYTR+sJPvjWcjMonC4x1uitc0JsqSZwonz8QF
S12VdXiDpFaVBIa/qrBsKhT6wOJn/8TkYH6OdlrDTF90e1GSuusqXpMUJjs/Tk2fzJ0NwFpl0jl0
G8Pg4IzOSiqRY0EKP+kO0d3cDHOihlq9/GVgsAimaqnVjI55W50afh0Tzh91ya7Y4GPWF6iGlbxM
hW0Rwf3xcFCgx6qPrbXSNd74qRsagjAHcCsHBCwI7CG/9eaY5txtuJYRaW5Iqua5H6Ah2tcb0mq4
3/pONtrJFmzpyLRZ6elCNfMeXDf9+3YY2CAclUYkxIGWko0/tE/jK/ya6W0erVv77uZTcnNHZ4ng
6Xy2XMgl/1DtfWm/5/vQi0rcndyAMZZFKHjGfAlwV/A7SRLRewGmJtA+XnfAfkLBlu6lf07aGuAn
LfQ6lFIJMBsE978iJIcwPUNmxle76QACxM2EDLF7PGlwlN7zv3O6fKyFjVxP5GclTobzon4zu+YZ
GkZWriHVOJ/zA6yPp6K3xKTxdtLB6UOD84yfT06ZBV5Clgnu0VV9IyK+GosKNzB7yjqgXwywV26+
431CnZZfTHKWUJxYZAFd8RDWv1PF/6WzGS5m+k8Q1h7xfjpu6Qy5viW1IEa0oFPOs6aw+j6rnLN7
SA1RT5ETUTqfRhI/9HVsYJ+csADacAxr1kwlPfcEmnq1mH1E9ZSt4y8HJyBwXdwEAXonW24aHj+L
9nXt95ne50F3isneJ2pEF6T00z2j+hPuBpRQIkzVRyKdWBCWy+KqOaZpLdhwy+N7qnDtTHNu9u3k
ATsfA3Gn8mU/0pmArHsab0PHavKRQQ4Oz1o6B7728UiYCFIYz32h0tmTgDKhTK4nooXJ4wzkOfOE
72NUxEB9OGjxL2pDuVcrYnW41jikWe0HeIeI5AiOUr64+vMAIs7ywUrj3c9T4scsdaqKtcGA9/A1
lY+ZoGgSgqaVOkPQDx43+5iJaW/MIiF9IsyaQwiQ7SiV7m/VVwR3doQY5ogWtMONQlPVAHh76AUA
SP+sqh2wLZFnOyzXBinXu2uBXzYUFYpDOxOqsMzdF0qX/yRqetSGNmdmT2tAyh9AB9FB865xu+II
xLeJ+hlhkwXG/uFdB3YF/5dL1oupZC53pYg3a/UJlL+q79fsiKzA35WqkngJK7afaHnnv10xxaJF
GPIxiUYZIvyV6v/kQmL2BzIGiUtrP9Flm8BLlr/XpYCo315N1IBnr24CgOcuOuY5Lub/DvAS6gwe
7stlgX1MzKNuZX73lHEJfmrTRHSh36TceAw6QnasFzno7FMTTCrnC2gbHBV9KEMsIN9zz9vKBs3Y
wVkS3sq6lGd8le+nIh2W3j/ALleoQG6WokNNXia42oENK5RYf2vPFkhSU9KWgiQLTqggmWQrTL3H
7tXzXzcMmeSldzq+T+Xfanty9+bBfVbazQGT2ZCtgCRzaXZBoT/SEl7vzZ3fxIUc1dwXL13zNkld
XF63SBzjfvHWPzBuuv1Fdo8j3bUnKE7fW66heuPr3LNbxhWlYz+ChNjvqIxUYuryBEwxdbq8VAW9
sYpQ+juP1HqhxcR3i1JKjrhQXKHLrPnNH0ZatYsziD+ODIaRwy0IRleuhaoj+2njdkCVavAjCYBp
3Rq5tW+21QDupgR1efW7A1XGnXJwjQ/YZmVt9UkYBdmNWBBNUEmyipxCDJpFWsB26zqvXl19Qaz/
K6kcK7eFWwMIOrJURPzsHOqEC6HPTjJtyx/Nwa1xTzXhuEDXnW5h04VcTApIQqQk/ZF4q/2UOo3n
AA2be9zLWB+eD4kxo9WkRVoZxUwDB7HdglgLYHfFs+YoKp85wzLIfTXU8y5hhYXSsS8036Sqvdiz
uRHX54jZ6nJQNX5PpMd7RCoMJv4slo24TTNNtTawEFIWnYrIaBBfokjQkHt2nYthj0IDUP/12o0a
WfZCkyRelBsvVMbyBAejTze64uOFsUzW4D23sMHzg4+DwsONPT9iK1dx2o+EI8BoTTHLoPQHMT13
YpHXchH21Kqcw2rpjJFQ21EupN+RJkH7Gy4lqDb1ctPVz2gLNrRprVceWQt4DkUeG8vlutEPCmS9
S3S0VctfsOOcJyBs2FNadmd2Kgm2HupEZy5MeSH4ZK2nPPHkPcKvOu2Yp3vDVPIOj0y5zzQiB1Yb
bxjs5+b76K2Ib03NbUVg7aIutL1eDGb6teZWm7onkOJAcpy4vbnvTk5Esz3A7KX1VzVQy+GolG5+
d4TY58qHZSz7DdA8BC98t63QY09pWItXYaNCLuxychJ4lWGteM96oVx1unWgnDu6B3B3W9teKXRx
S9eo6YYgdxy44KtN7+SymWb2yVHiYTWoo5D3yAhMaoDY7DPYVIi8j2hIreOhTNiFQoRkVPqOLbkB
9Y6FELHjbtl8xJeecbCxtXxRrpPnIDT0VHk5V6q06AuWYPNxA/QcaxJIp5D07tWuE0eenbW5EOwu
ZNOlwuuDp8Jk+fbsKnvnikEj7kHH5JvXAVay5yY2+CRfqKzBToiYdOB0KCjQhWqLBIpSOWisRnx5
unLZN5P5JkBOtvi9QJrY6BKpbfZkFmga8inJ90v68iMl/UHReRTDsmyg4TtI6Vem5Zjj5ImZWz8C
ajBX+AKOU780LEXUsxmKOnN/fhRQZWoaiezzOMdjELu5Dfn3W9f3HxBZj896eiUFa6JxBGs0U5h/
hUa+wrJUG/5Ldnhr4P3H6FlGSQtG1nUySVNGcsCMMLNjb9ZHEviRIEXaSXfrAXIlICcbN/cHm382
YLr3NgjkbmtY/X1gvhnYPvPCKCKYwBELEIvkRc9ajnSuStu+PR89H3aVrnEWUa5IwMXn0vg/wWEZ
6glZLIcbXhst3DaWuQMO8bX7Kv4b9MRM+7drnfbUbewvZlP1lptZyiw5lcdCGNofkqXAZ51xlp0A
D9r58d1J/CprIcZInKdGQfDD02pSSsdhZV5tlmvVCOK5cjtkCqDpKCSaTgSXfO6KabKeNgjcs2+b
4BmqnC727YqjzGLx9Mr1e1jv018+wAJI+xo0yb+V/oxehSInWI2RxYhJt+ZX8ejSNZHA5pMOh0Io
UiWgTMmbg2zJ83LwFQNM/E/RZ+HoBJW6PgKYThY1AbQCjjMaSbzbrPMXiy7HDUDIc1/zKHu3Q9KA
b6VG/hNrDkrF3oRwfPx1pEZTBvsxvQiQ5CXNfKUpJR4vNU+MTNV4J4kbfiRGkfxUgEkH8P/iNmTC
0L8mAYdrZF5g8GXjWwHg3tuO7M/o2OiiLLmVcVS8PKgG9Blt0jQf1GKjbO53levJtzOSAn+gop0O
OvQ8659iZixfKzPaarUCRWl2AijJ4X/7LTgu/PdaALn5+Ux04AdzluqRm+NQsXS6h+aXJNhlIMsG
Xkk5BGF6ryYrR+cF9ZggAiNx4leEBAzj2Sv1PfHK6ifYrhGMgooFc4gaqSz/ATRTDfH63JNPFRsl
KsHhxHXUaXBM9PMdDjkQQ5ELwownklSRlZ8GmilShljRrSkllgnfTtk6pau7woQd/yzZhzheGTfi
Xir8ty4aApTFtamwc6CrW8F37owWfr+oLK0Epz4IeOVArx6AMqnOuJ2QmH1yD2OfsEZ9XYQSpxjx
giA67fN9Cmb2HdjaagGRCW/HZjcXrNxBMOUc+6rMZc9sWYLwb7tkpDc4s9scRDyPskVdcz1NAIR2
8HCAZTFlZFWHcwXVKCf9B8bb/7jdsKqTMGph1Z3u3EJaNvfyPkMoSR84QP+xBZvdNAa6shoRi8rt
TJrw1o1CEVHkD9zq6G5nja2HSftEOnEd8K4YCTC6IFvFkcFja3ASGd+AlHJX3JNZg20eM2qYopAr
hAMDyUCVMKABvRrBS063S52zRAWPLC3UJmw4blIhDHvglCpuGszMnI5OSXFylKbOR80K+VndihgA
9obbwpCrU3cZLI2ECQMZ639rXAVTvL2XfKiNgMPXxTyutZDlmA5/r61p7zG6MNB/30Oym/D1oiPJ
iZkWjENxp/cjl+Rb5LUB/XreGcQdDhYdbIfBQs6i1Y2RprD9mADVK+q7+j+Sbs8GPB+TQPfzcaoM
5MC3uKh5f6Mad5rsujCJ3SHVSXYnGdI5yirQ/w3hR4yHm/QJVgccR0sYlZ3jFGh2IcvHI+zcYWJJ
BRfb5CofGiXcM5c2ONkuvjqo1nuaVKMRMXNJ+R9JNkoWvZA3qchiBj8a59OiXvmlWeGf6S11RhPR
3d/begRqo85SFGX/h7jVb0MUYGy84X0t72JRP1ZYn7uMrtY4gWe+crwWAGA5A+X3ouxjEYw+tmxB
AAvrzsQr6PXSwwz8USMQpv0sZ+SSGW1uJLJX7X4Ij+Wtoe2Ol2vOLMEqSylLYQr41EiT3CGgvgXS
d1Ncv3LyKSLA2GRdvdpJIZ9xqsZSncxOg/3njen84IMxL7vEqTsGyCd1GHBlxyatMhIREKLmNYuH
SE7jRnKKGD6djrBynpTy3oWAo/5/fJpg9SsMM7327DpVwYgSfA3EqcSmgZDfwlE9Cqqsklx1NyM2
pDw3CrJlSv4ffVvc6VZHEpBwotZu13Oicd/ZHgh8BEQpnBH/L8yIO12gkYoIEN230GV6ADEZ2XWK
5Y0z6JvutOKEXsyGUOTvAArIemgcrp0o/sC82UJzmkUXwD/HvDX5fHCRhTajsk8lQS6Oj5ORGupK
KSviwT4ESY1eZgOOmAMXJg6LzqwI1hyYoFaOvL/8NHQj9O4wmRgcFh3VDuS5wHOv7CENyH8nCsbF
JI5JeYQEaGjOBBwIWBz8jFkCvtLeuMiTHgRhE5E3VCthqrPhF558uZ8vcln9DmQVIc0cEtD0K7P4
zcEMGu2j+hx/oYRIzlAL+93BHgk1+dMwM6j89S/+e2hroQ5vVDAAS2nLRk9p6mAKvk2YlDHQnCxH
2iu9BDojvdcZnwobkrSnGNXzXEf4tsW/2B//etAbqecaHv/YjMXYnefHZtK+T3Pdje07l7/ufhj0
PivUqVUhJZkk+TPpAabfLnA5WtxDeZRwSS+MzjhcmOzHPwfn5akX3IUP1pTDFzscjOmYDvR0omkl
Wtt+v7crEavNqgGZhHUrnVPS47UZ0IxLNQL2HYHAqwRkl+5Qq51Roiz5rlrimm1HWgtNjSLR1R+M
ip+g09aCQy/NWn1iSBb19z53ZsSyXrYSxoolmQxmTXbRLiIK6tBTaDImsOoddXZkHsRMMmXf85SB
srhQl4EIsOQnDGQQ9ftnM4a0IshJM6U4Bkz45fT68cPejEVMEIsV2jV1n3yPIptMmW8dJad/iVk+
sepy69NAP6TR62IKieh99Nk9+e2KfkoD1kZ0J25026HOtMxZKbBbL/Y1KpIYZGrL2e0qYl61EbOU
Vu9Us05K6i3FMbwLU5k6eAsfBzbtd4zRaMbd8oj4MV1pxxddOc1ODdUrrTA0sOhW+ZfCTqgJfzHL
ooxa8mCkwjGt71syOfWzRhrxZVSBSsq4sRow4w2bVVaCssFvIh4XGDQKwI7RB+/7uoOfq/L/a/Wp
6Rh+CviEJ7mR+niLfViBnu/uQaENfVnW5UbSosAxwhUFCer9Inst8Hit9iDuCN0EoPYLrVmlPIL7
M0OxOqrl49Mkpn1txEipykFOBIjSJbVZZF5Qh7ChCxv7enqUoObSZxbBSsdFQDxpmeCEmPEXtj5E
0Cn5iLGahm+6HD5X9y0pXgq16ApkCqRzH4914LVy0mzCHyrXRKCxikylZLCN69i+Qq2LWzCTyMb+
iCIvdYmqVQZxJ/z5fWKMzolXrZUTlPkHH8twweK8Ayk2JU0SjnS6M9W/VuyKd4SsMihy6yTMKNJe
k9J8skgQwVO9LW7S5kgj2ssv/95A+Ijoqa6p5yk25RNqnqni1TOjlHxGku1MqZQk7w5RGaCOlheY
nQ5qYFDZRkJiu9Al0VSaiGkpEXk2Xijkp/zEfZDOwkz0mWFbCmAHAeF9qlzUoqrRGeDEhrktXi7u
VTczTqwZPT1KHuKdPFnmKey49v1eClst9v7Fcv6Gz09TuWl5eahqKy0aqGmwfr6r7jmYbWweEjg9
m0vFuxExWaYyOrGBX2ChQV7vRf06GoKmQnX7ZFNaZnssV6ONbiNdzgazxKO8a8AizAns2Gl3Ch4u
bqfev0oYRd4Pw5rzxthRgK1T8mYBFSlpT5jiTfMR/LBZVRuvNA9EX2yeADNaN6wR7G1AenS+Ym5C
gfw2lWTGCFsbImSpsLE7cBElUWmCMLEGCq3HMOBINtGO/mHMB63mlVLj6IS8RrTVIGA5yHkdAr3C
esTYdwbD1TYoDa5dxZA1B/bEnpZIsZ4u9inP1Qqxs7RjkoeAoTS7MCZDiQbyXSSzFK0+hvjc0EhX
I/PDWgXukyNiadV+db1j7FsGNv1gj7Q8C+AK/KZ2NfLuhdb8D8vKs/KhHZL9IXUTsDq9qXCSASOf
ClUwRKaAmk3JofMVwhq6z/uY35JohW/4tdH/8qW9MOO3I5O3+7taI1t2rhGxS03WqQDB7TcIxoGY
APtKpB7wMEqi1wbPU0nB2tPitfPBoDsx6POd8CFsPMNTxyTg9QIOJtcw0u0RlaONoUDJa5SIwFBz
GU9Yhy4YdpTB/yFFaGZ4pJFbHwm3E8frkqCwkaSe4UwKfQCIm5eTyIYrKNay8PeIbFKbu3sHGznF
ziNEdxf8jZkvwv9GYSwu7RrtB9yO8hO/SHUdC5ySdec1ODKIA8xrViUoKWoSwH8LFT4I5r/f7Lji
dT0j35Yya2X8RmJTtNlWwq1jReb9D1LO0mM/PBwG79rSqU84fbt9DEKUhkhHxv685sRs0MXdN1aG
2a8BXf0JoLYBhDvogEJ5MP14lL/OqgXCUGml1nz46tqGiDTXKgLRIvkXPXP1MkkKJAf2CDN0C5rc
tmu7ddk8U0jJWH65a/u56V3XL29amopv7xifNXtzr5UsVE0bwIRMfLnN7FX1FneCdFlC0Mv4XgFC
/qOp4d7rnhG0oG8ZXyanaaQTLjunsbTsictr/gYsj6aOJeknXodXQHwnrR0UlGNRplIXwKglRqSa
qW0lDShAZ/np7GTZQ7bIEUiQjpyhd74EkBlxcDbh+ZELjCWYndJbx60THTnHjS9X9mL1OJH82u/n
0QDK5QBTzmJyeQT4EPfXMxeiQlg+WjeiNAC2rPXCzw7zL3chQkICxN6WwgNWNMojfZFv9GNacoCY
C48cH46dcBBbe/0nvzbg3x8blsH5BpWeFwx/P+fZf95aPcSLqtpiD7/wn70Y+Ip1YGG+YwzaHFkC
PR7CQR/1IjAY9yUgjZ/UHzz55giGAlor3IuOJCGFj7bbj2Ws+54vHwJsjmI5bs4XG1kPb8P/CKOr
sgTiTfEnJQ6jneFumd01/FH/3k8Jt1A5wOOPIviweUVLuO1UCSMURYRFcQjsE+zC6ak4bjPXWJBH
BWILeepVavwO2gvHRx8vHmj/Sks+u2E2/BxmyXbWpQJSQbC4MP4Reuh+ZqqpM5g6/ONc6kzLSou7
rAnHQ0rUgyrMGLzDRp5OamY7WV7uNt76CRB5789rC6XSNsQmkNjeUbv6cHU5rL/za85WDZ32K2Tq
Re3sXuVDfHRuPn3ZSOPLUE5qurRksl7JS9Udg9EsKqc5VFDonTshYnvyK+ymc2kMCmpurfrMnz77
KsbCuytR/9Yba75Zi7Gcvo2jmlpFBw/hYrC5bZnerc0NVLeBZ2S81iB3GPhM5LJHrHecbqa0HCtw
mdzTIgew20ej7IndbMtRBq7dolgEEMbvjHMW+642ZL+471A8RkNDVS9f4PypWADyOgBXPO63gh8N
a8/3h4/eod+r5Lzb1gaS/5SjMwSbQ8H4+klvOlIA4hFeSsdNr45A1IfYqKZXE8ZDacK74oJFFPHR
p9U6W2b4tV/foRBmCQfxcoG89cVLbsE7hFAk3NNb14jxinSVwLNQALNKy6c2uNLJ79aA9fQgbYL0
ZiMM5RaqpiW/5oIxqLY/dLl7GxC8z4eC6e5KlefgRGCJLk1A8vhKeIlYjlsccycilenpodIu+YUE
ICsnJgHlus8hrbMsmDXTmL05JdkiZ8ljRwvXNASWxWVK2VHNGR18ZdsZx/ThNUpjp3pfynDCedd/
gQbwootZzbR0bWQG0QAfXXY5RDhVr89wP5vAVRUR9s2lBjQSa0iPXZxiDW93wLfpk7Badpzqpllo
gLIxn7m8lvkFgxF1n3jeie/4woQ3Ktxoo4lGjPJ7EbCDBGmupU/yc9JqyazPbKHiCRgLeVd/e24v
PNfQyRvawEc0+OlZsn/8MhZRKVhlfxnkbpnbDTeoqXioFmUB1I4GVEAbDIoxweoy98udemMOyaCk
kF3YlOG4Z1HprT2JydJzK65upGhLpgsJ3A0jTe6xPjwKRKJfOpvNw2VNS5fR6KmNjIAQ6pJ1KQ/3
m5ikUlbtbYRv5EZWMHDkFOAlmIldav3/JtUdSXkiIZ32IjFAV6ivrPJi5Gh4zpSehGVL7fcMvuGW
7GWPadLtk316ZUqJm2pzORgJn/GFK/A5Lcjw7uBQvwOrNJvUWh/jOFZ1wuDKXMDlW5Sw65/YSQST
NSaJb99z/0EXbyfvVXrUBCdtaBvID9P6sBjWUp0CUh1XYbb/4bk8HIXDvYMVkDPGgKqfmkoI9kHc
04LVzmKnhFjW2t1Es1OFrEKBQUqFnAMzo76G77AMgXDrSW8/km8yvQhTP4c5OjV4dSrW5W5tcp7P
BLODzB6yGjDIz2y9x2TdAoQ2v5ecdJ9XVvOI3iE6KQcBvuwMtxnnrW9Kav1Y5LWnjtUBV590ha4h
k9m6aswe6Jea1B2nUJTwQv/fmjMbtZSMWk+QVd0K6isE1KofziahUaO/NpPgNnnMMJDGYUS2q0Nz
Bg4bYFFaOSiRbYXWDPkX/Qqu49m436ssDv/Xt3aViDRtuTUVkDrAOp6ikCPDEk49SYtv4NVsEtxo
6fHgD1owiX/oaTcuqdvyo4L/6mnhQRfcXrqM0l72KbttWaaTMetmCRwiYaARSQJrt3U8HdgcaFtg
VVv5hZVM1TPSLC+G3VlkpNrx8LjoYGIgCoTH2dPpzlL9d6jW/XHsNlSf1JQfMDA2M5V5z0qwjLIK
2hewP6DmRslTL9wtQDbImg1sYD8LvjlHdDVPbWtQ9LoEW9Bsh9TuZZ3xxp/Jn08wfV5CILbmUOm4
7187vpc5MPQ4tKUeaMXykIHiZ9Fe5zmxSFsvgSmR+4y1iRH3rw0G4O430um09nzFn8T9d/uxTHeO
IZwQvIjHlMm4uq1lww4R3zwFVBt72246ZClRVaMrT13T6Y+B8YB77ThVyaxPCl3IJHMmHSt0TvBr
84RqGmAKojczyCBcvE9717J+ikpNFgCez3MEJERmZMRb0nypASmEPBJCq4Jl7egFaDWd5FgBzOdD
gJIzGCqluA+MTvGDL3ylqnMLd2VNSRFOZdSdS32PvY2ua5hhF3qIUKM0rfjvY1Z3x0DIUYuEnIS7
T1gKkHmZdilpPsMOSXdlDjCfj/J/4gJMTc3HNPIeIzK0cr9iRKx4U/AwAAcalLnP7R5hd1dxEgE+
lJsdE90UL6ANaUOIoBCSKwYZIb0XfCGyhCBHtN9F6lk6HWyubesdJKH9oPYaGr3LW4/T5nOrja3I
DjjVB2mUW5A+PKcml78fRP1C42qaNrRjmEP09omz+vebGZleRRDZcSISscbZeq5GeSR/RLONsLV0
p+bujPRhXf86sjp///GTVJClhBL/jEWO9Y9IVRRrRfEiIdtrv4eqiijxLCriH/J5RxjpjibHEEI7
/GffCY77izgKnLXSwOE5wyUX68vCbGvFm18sp5kK61sYbjwDwtMmKyEeepw+mc8Yi7ObvLNG1tNJ
mReKj9MPvpFXsKsAmZHxY9KsmyKaAN/RmrYsGq6ZX1N8LAvSfV8aZAOv4hl9QWehYmjtBv+djz+C
HJGIQCwTpqDx2qybk0baERt7HA6SBHQ+BxMfJFw+uYZBHup6Ae1f4VeglwUUQSFdJPsim0mDHluu
c6kHItuOKHOq3AsWRI1OZAgNm42eK6uejm3bNbUgDr1IxgKjI4noL4N9nGq3etp15oUwx9spylHz
bsu14Cxh/B+BK37fkdgeACtXPGpOfaka7dTabCdAJPJCDofD206pvl0+Bsxe5KEjrrLKbhfzCSTs
xg0KuaPAfnO+CkOUKcwY8EOLwDQ8OM1DH+xEBzEOcCXGCPHeGXAWGdzKQNIDVJcwN5/MV9kFNaDT
4pxzZUrBwp/qh7ECYzzQBlnzo5L3l1dZ0wRhViuQqdrrjVDjYsuj6+KjDY5UhpoD4+gqdYqbx8g3
94b3/5+eSf6q33NXsyvFLzee0EizYNeFgWNAwBIdmPuxrsIHpYSEfqC3laPG0qofAevhnzvofoqA
szMPVXc1kLzckhTzdC36uwgjTHHe3L3GQzo8VJG+peQ1em1B3lZD+3HkAJEZQNlpdxO+de33/2fo
IyQ1FKgS9OIIgOcN6NzjXfIrojpHo1t3tvAV6I17l+chbtBz5UFrEnA7LZWVjZ2hC1mzjS0HQ4vq
s4HfPtP+egunlazrNP/DngMFPtOS9QIwhBnfuyS7c6IEQA+pRAQR/yswoBsXlHnN6aLGP1wIy186
jgrdYaYdtu8WHl1xwST3MTeStzTO8nyq6QyirM74aiyY67nX2xSOORgckFyTV8V7SKNt08iLJRUF
2lUoOIMXzB3SDrHVexCsrbXACdQnrU2nsI38xEFFBXuFKmaRZrPaHwUjcbbL3Pi6hegaw5TQk9cu
J4MxgLju0bsCR0dIUDbcVgxvirE1LybxmGYRm20hrIdpU0qiUofPEpHkQVf0FPfx/CA38kRXgq7b
n/rYmUoopGSczeTNM0Le/PSKRbcVlxlKgYM/3DZKrSLdFS5+XFhY3v5Yg3Y64S7vO4iasIsWy94f
VO+0WBwbM+61VRtOLmgaxBBU50wI5xW9Exg7npV9ezShM9Z5ivSJUL3mSOgNdki/FcNBdMe50UVl
XJKko7POPejiotpy/tFPhRnmBH5ia5Qzsux0CkQocr4145uPwLwoECfUsCp2JnQaDyEZBGs7L9pm
QPGM7/DftzXIdhBO7cMsF5m/Nl/YtYwW96ROHPFaCzkf7m5wJQp0Y3jJ1RXfh3YF+4hl5czcGlgn
okSKdUuqT4MZTO+ppmz4AY29dCUe/IE80d1GMpp5Xz7BDCVjRX/BCvFEAfJB1o8ppe8o1b9sguoi
R959svP6ks62CNGQAnSpmKZm3/lEYLShVxicvBt9miH7RQ8ZkVCZBmNL1haNZgjQJmqf2ik3+Gh8
uNTV0fqQmi/QSREzf52jXRMJpac6V3wkbutUoGV9z9aRbQ39KTOLpg82L0WZuFR7cf4zaZ70EwMr
M4fdtsl8KTZ0aYwyLVx9+ZCbyxCSS57xlnFw4GREMI3TzGotugSygAGgH5CNp5KO/qGd+x1/CdEZ
vmmI9wqYdJb3SHEkLUQF0prNgtSFIvjESMj24Wv2Nuh97lGwBQ+7aniCC/wNQ9pPHqHeJDcmMg3n
koO1acKU7Re4dfOdHE4IJsWcFfiV5NSfTyE7Mjvyb9SLWVFoj4qYP0O5Pft11wJGkx0ePsaQmW+6
kGSx3ciUXm26kHC6JPcUevsLRAqa/OePsdi9M4uIQquLwONi9qxCRup2r/aco/L/T1CagLErhD0m
MtnZPyIzY7Q0eyMEijwdPjhzkbHzlosST8fVodLboBJ95DA7DbLccxecfwhSgk9c7RfdlhXVXcbc
rgxAsNZno5oCjDDoz+80Ddk2vz46R3w6P063T5MQs1Fr2zowzk+feOYzsMCzD22mgXYnpQSE8TgH
nC5JD+Sy1F41p2TUjmO532ubBrpdSOdX9xvtcvH2+1KT2RIvOilR4dznWuQqA2AR+zhIfNT+6U7O
J70rtfrURBh7mpDz+U8E93X5fBFXeO0VAAbhtYYB9dJ3AtwjnGL12OOJ9snT6bCj2dxdNiYuSdby
DxFGveZCJf8NS5HjFw6E0Ln9J0T2M10Nq+xH31OCqiH+QH2pAmWCYVUQM+hiEqtlXoHkJx+3drKf
zew8M7yn8BCwHJBFmSTc03yISmzoNljY1G+INRBqyKUwVBAbT0GN6GiDQ/HX3h6TILA07yiC+R8U
yD8wXj2YT7Gdp/Is1/+VE3nMcyvQ/rk8Q/asDNUHf4ThnYtnbg2RWyk9fp1Aql5qs8KQ9Lze4K93
7Rdm0+xmC6Erq2dfdGJPG2klfB5dnEUoe4bbmQZvELaKMmRP/igha56SrY0COGquaNwnduPJKNgn
ukAATXnaMh5ZobCRt/cijZt1xCqFIxo00tpuw43D84CL0AollUccLEBqcfH6uLGUEt3dvKeGun3R
0WZyUCPCilc9DE3AkOUDYwP4kyVmGgceHX15uCzyF3LR4mv6H13ZO3On7AzhZ+CAJ5g83nLDYrZP
Jwn6Mjt3JsyY/tF7saILuMcTVgoev5TCHTEk/RcPj2/l+MJYZDt45wIv90IFoofmqbS+REWyzerC
Xb2f34+VNjaK/B2eeablAWnyqmoxVVa2QNHugKAzTfta5DVR6ULLJhj/wBtVVj/USzsjWejD4Dge
Mq5EB+sFkQkQOpwiAoH8b3hIKJFl9hQVNzO3BJzrGvTbnfwHwbGtrHGO3cyEPXzX7M4lzv4ycAmW
2n8gaHL4+k8M6Jr/w1c7T6P19Tlk+XKqKI9MOlqu8leReyvZSXOCq3+WtxV3PWsInRN71iAkSpcu
t2l77n6ie10viKHOe8zmgdcVcelyV3xa89hkAQE3Rl1YTi5lVJSMSwRNnX7waUWBpLPqXzlqgk3h
uwWBNf48HWETDk647pk75S3c7kc87MbD3kOy0KdVT6OlYcFSnFMCB8nHFsWa0ZlU6lE3vtZh7GZJ
KyLdoghRznIWrYSI9Xl2a7CRtUqWpoSXsorhtjbG67a5h27pq7zaVooFRjHJXMGvEdeSYmDiINRd
2Tz23eSOW8FW/RWay1s4hm8LkWnWgk/+rHiRWuDwEs6FkK1rBzWG7DVKQodorFVHEzBFUPPYNKuD
YvgvnGUQRCshBRa6K7jYDYpmP5Rvb9OEHw+kRWUHDOUtngGlMKTBNAiQ3tQjZ0VU5bIinz0SUgrQ
5z1AiP5ClW8DjsNzYm2a9rfwDeFIXKRNyrTSNKJRO2659yl821FazpUukoRu7U6yAo1WOJd0YnVb
7gaxrSuM99GKlUjrqDfM0OraK9bxVaeKCnEp1e9yOaRHJMXq2Ws4+UFRD59sEUTS3GQ4LurQ/h12
0otnaZ6gHOJzJuMKvCIt7azhzM5/pCyHIJP6MYwjQHpE6IBA8YbSjhbLFJxNdtUjj8+06EZi7WWV
073jSlIbnBLSWX4F3n6+lSyka7M7vOX3RRTQ1Br+lWmjPaHhxWCrtr/zBTRKTBR/6nVJodQgjHUR
LvzVgTGni3Fm+vCoiXYVII7iReGg2Y2agSi1o6FppbtobT926cgdzv564av2arChgtsOMwmmERZi
QSaxNe3Y5BucX1THAin1ikSlv7s0rByzzUYyxyDh8urv4oFFK8JeMzC4wGeXH40dTJUxdy8iKWcw
xQinxdIudc/gMIBhOibLTXZZUMei0J7wiXuIkZau3i+G+MSVzYXk2JzGMaB4XqspK/lH8ThfI7Lr
7xLBYG62WQNkadN4uDZcPCijZCh55hyhcwTW+tOEp+5hijS7iKCP+w/Bob2Op8ogzQWium9K9n8L
kSajJ+rOoJP8BIClVuyM/QwBwDL0PEdMGMRkB2HtpcuRpciKKE2P5+d7RzbpdjouZUNjb9B3Lt50
0yG+PyEvEuYwjVTKZMZ2PsbK6siZhX+WrDtl5v/whpiIStx6uK+kETX7UTQMU/tPGQwkEkufWxgI
Fn1/PpRddsp95kvysHKv/DNQari/1Rc6Knb+RJ4ELGR2kCITTuFoXUriZNwQCAXNFdocAO9aSK65
GCR0yqVpqFXgMjHsTQ+prWLRPH18+lpYPoBPTEV/Wfz3q5CbLoUg4lU6sXMOBx06AjZefwYOMkIR
8XW3TAYwU0TSlRW/7qrKy2BLmaEY5oWEeg4G5gDgOsmvSFoSI/JG3oskpmVWHx5xYT2sNq2ADkiL
zsCevAap6SrjCdgJoprP7kiPbyTZCiefFoS27rqvVZQDZGLSKzgYptkpYmPKGCrPhuAYs8Bv9dxs
qRGYa5T01qW73DRK9QPeMtGkkshf1SLa6eIjMPRTCFct8DtgeDh3c49ZHA7cb8fzxm4qQ/ygaA3k
c9ekoXdysL6tq98N74epDY8nmK3nUmeiq6oEEwkfYI4fCh5dydKzznhsFqAERVnPyC+rzMaOFdPF
qwqWer9bZPRScOfPO32lhSS8a+YQhodQJealQA8ddJcCcNjMqPL89zSurgoQCcz3Tn2ghu6IcoUc
e6vHtifbVLVZGR2PqDalEP4BkKY7jXKKC1lH7UsCqNzUQCba8rl7NKSC4BCkbYsnb3VhSy1NB47J
9ojH6IGyA8goJH9kgoNjYiRH//AwBdwhsLVaUkmFDNqq1z4NNyul/QhyDl0CSodhJh8pqFBGxdm6
fqEuDQschVM2C9tnSkDkQReEgw4QIMjvAPscl9oZLdWMzzuOMk1X1GL1KGma8UJpfdOlEpwEsYvJ
ruuY0lcwyz+XvpYJw4+yy+YYWI32ml9FIWkXtmV7K3PEnYyDegg49AtpfGhYtiYJ+TrGEJrgyOBE
7BIH91p7Lv/1YnQ81U5QN50TMuIuD1PLGob9D6vuaTAS9yTXbj4YmHmQzoL3Q5yqbOPuIBzL80Tg
QDzQnFXG4m39GBic5onuC8tvCEW9tQbaGvZSsgDjgweQ1N3oDNP4U3u5ADk9o2pb55luyW/rt/Hx
mYraYh+uzYvpYpUMCCx9k+mIoeOhevPt3le2OYI1M7/un4KdL65mygAJWnTRq0URzrb5sRH1po9M
Oa3eVzjrkFgGNFzZNtAOziNJ2CZgVOn5XbqqsHSGHUNUF/gYscvv0IUDpW0ycJwfsX09GxWXWl1Y
87vC+2ZG0Odn6Bz+fQMm+q+bR45vv+0KbNRKSTuK41GXqDh4HytJn1j5T7sVQV6S1h6W8DQbMEO+
IzPL6AzCk77fazwaYIoLSvWCfkDB3koEpc/MvQuwptnqlB3QjDUvKEvR47x5HLQRFc6aA0UT91+3
gQbVEJ+lWNwwLy7XcqCHjA9ZMjS9S6q+C1llT8bbgFwprwDN6BO7V9rhTjWQtbvdtxv3gZRYB9B7
vnuCUE986ksbf4Z8a/Ls9UCDCssr5Psc0OsGtiRdfz3nQK3AHA/KZPPhbxsfm9aaWQOEq+U5DQ+e
ueilJ1/qLwxVL4lnVRElAngSK0+MF5rawAWiAnh2PKBY1JwGcLa5IiDZiCvPz/snlLFEbNZ+zQKi
qSWJF5HjaDJsKsSx9Js9XY1zSUHEk7gto1gjWJX0Lqej5ZeCZP69BHW5VhNnLPEtk7vwobSSO3Jr
y+77Qyryh7+BEMpZF6zeEt1X35OxjL/OjRyH7NJ4aYH1eBz2ySqIU68cg1urCsxb5mZNYORn0/9k
DDTQCNRNmwXnHXeg5Da/fk0Q4Ukq9CQMQTh2ZlZaVo9YDrcGfAEHDAeCbGpu4sWmrahHOACpEba9
4jOwwHu1zrxEWq/uV5Q+ZL7x8DIQ1sMVyjzNq1+8+KksUFAgWcleeCfh1z76Z+x+Efb7i9DvltaU
yxFm6uMHL4w1540vOPOfztRpeMaFAIjupBPl8QeHKjMWpKjJJ88LYofx0m4wL6M/uTwmr6xiLqdq
w10LOg6e5ZTOyJjFgE3JkkGfaQoBZwS3ROKgUY99tYFFcdkQhjI2p97iG59RO2LPRZtBPr1DTV4A
iB0wN9RBJ2xWsWzpvPa1/1OfMUm67Ro8ACiNAaxNzA9BlXSPDevCVNJCRRXpkP+Cm8bh0hxoEKDW
s8eGq5TtQoIlpQgbvMtOqYEHN2zYw+vgENUTVEzqnO92Bu/hdvedMUGqr0heaw5k9I7HaNLBJhLY
hNfJIuBTfUPcFWV2j6T4osUh2VcBviPqEyK7Ar2bSyJKJlL2uVJRmBpkC02NaBt9MvvygKO/rvo4
C4YPQckA821tIioZ2BQN6EQTeKFSF8/ZPojgWjAE8s6BWKQME5H6wf4sLDC8QxTaq+0VJJXgsTVI
hxaIRGFnqqpac03Do/A1qq3Ow9S0wzuFDaePtcB1GMbSdNaazboYrEIH2OI72d21z/VopPuRzxhF
/2Z7tJN1r3x5HbaHQ2VYbzxTOLRuqix2G0LDMI9L6CSBnwrxIY8sq7QdEmCgf+wt+D6O4KOumOP8
qXXwOPS7NTmYqjVvFiyPnq56qjAXijrmOmHh+YJq13O2yceJ1b3RjADRnxltAQuFgAx+OAGh47ic
hTs+4rkFPtH+Peap5Psh9sO4XlmQx37n/ulAbxv8zDIVcWP0ZDqQLhIVORLwmMUL08h2R2IvuVg+
E/5bcRP5S6gXCRA+OTeNAW2FejZze81CshZjkwUgz+0eHboz/ACvWZbCL7H9bUXaa6BLAb//ghNy
3Ek3B1JK40NIqIButIXhamWu/4faoasQhYlJWqhm3NQCORttJjjUzppeHmMKsZuWE8F9gvJcrOfR
FS9V1yy/GXTBQ1t8zuv+aHSNJHsRoLjxYmYTCWX9gDLgNwjKb8wviivZHYjAKUhFYMjlkFLQhul3
PDvgbI0+1/SG+cFYRfSUmbKznTT0/eCuO1v2TX6d8thDZV5ZlekCfOvxqrkUc5avaJb+S8c0Zl2z
cANuLgUQPRuhresG9wkR8DxYIOkX6EoL6Qx6QFdKHFeWbl6kjcWARlBt7Ye/DUGYweqGQv0CMjnw
uc96TS5T2ipNknCvgDrEmFBjmz7+uLEhQfCMZB5xjcjf8dA9DEt9cJKw/HJleAdacvvr/+ws31f6
kq6Lch9GgZbtf4Vm3UVqaKTJA2JS73fCWwxKTiKfXj+DmxAz5LmwWFqVsW9ecXJ4JxIjYqOytbOK
AeBEC6UhBhd05oFPm4sV3izJipllQhnioe8pPvaxKzIn+1wxjrlpLPlt6iZblgrGv96u5wTt2b1Q
JsUp88cx8X7XejxFm/OR6sDS/D5m8dP+wMiD4eE6DnG0BPpC1gbQYVioLg7Flp2cPd30avaAw1g8
fmzVwRyj5AcHa9uXBXZ7UHZar4rZGOizMopCDrCucvNjHUINuTeTeU5O6m4A4zPkv6dhFErfaOin
X9ytEQjNDjZSOiOnJZBzPdxSRP2RP7bM+ctfkhuSNyya/zI2OXKvI/3EYFpSepX+O/xc+cgpYzkR
PX8SALEsQpvb1IkSnAEYaKKL0vvpyjqoWtWSWMLtlEo1JeYw5Nj8LtO/MiAOhMDJAKC2GER7jTM9
9iz/z3iNvRhsrk9HjCSq0zhPKwpSddrl0RO6YmDWIL8XB8awQh8Fw+omfo5YRIOlpIoPJX1Sm6EN
DliutLxacr8WSNfl5mTA5Um0XGDe5Qo9KB7H2hXZDWxZMG5M5Xor5mfUY30PXocwW4WXNT3po/d8
hHfVLas9i7AsXn1HfJ8yqLuO61DuuYhuHPUpCfOjcTAmp4X0TjK/iu4TMRdWk4qUV0+ODbuybl8B
1OpNadX0nQB+gir1i54AsC4Eb+fUrjXOkoIItFHNkLKQKemr9RhQzILEt0smo8epRtpw/t0wgchH
w2TQJFlbJn7TBmmE5eZktkmeKxN7v3cMqaXGgXykNreK4EXLMHOb1G0+NhiWlRV9bc9+iP/XElSX
mpwOCByhgFc+nqR76edmH5mp1T9quozbIjI5deJ1mCgwR904J7pOCfM8kVzsPscXMTJPiX9gyEuC
zKlKjzAnCwgfaXtlB8h3yQ75g2wCdfUkYXdGFTav6uABvjNvxSGzHRlyQ/I51Y2vqOee0+2ni1sT
Tp/tyWkWr42iC7CN20yfSrDq0edmjpzsRUQZfAjLaXwDHjGqThMci8JTU2DwoccHl6aa5oYQ33/d
fIIC+DGiymFE5IG8usKabKOUggceA9wbI1wk8D1IzyQ2LejVmtE9mtEdZotwdCu07OsHEo53PT47
34Fne6Zg7SbEguc+CBZeF4SZwpf3VLdWs7bXtJ1MVq/NT+uMk5gq1jk8iFG9ewwRunrSfbhHMo8T
Y82YpAE+dphU5wr6KLkVmYuBE7D1Il3aQ1rC1dTMRHcb1ABwW5kfSorRhJqP5Lyl+LdWHJzWMSPN
T0Knqom7KtQCHeZCktjOzvDWo/uTuqnBnQJzscnVSTU0EMvJ/y2bA1ZH3dB1VdMJo+Mgswgm2rfR
AWqk5Q6JzNy7VXSKuQRaidfqZcjW5cObt1pVs0fZ2fIOcHkU2pmMR84A01Oa7JiJLINNZsTvePP8
+6cIGQXhMo8kculn2Lg00rBI0Yv8ENWss0V8CNKmj3P6uYCdBHk4aN4w7j/q+wZhjCAwSTUoC7Vv
vwj56mxCyGVn9/gas1NHvHoajMY5TgkG/qyOA0S+yVo0BuolvdT1w7DVL7gyw8UCRjxc0rQdsjBv
4bMo/9IdDLHWutnYj6h0hBPI5fHR32zEOHGF/PdxJFwi7rqUPnNjWkkUjKM1tRqjhG+UchIp4ViG
Wc6YUsDsdgHRSXTcO8yvzUrFpG+V4cf7mUe6UW29fAY6I/Z21HY37jG6HXnVxVzvZCm41PrktbCG
0m9mxL5KrFCoxMMBMfJeoKvUU35DWIDzROCK5kmaW072swyQ3OMXUdzFty/DCnLugtFiAhBlDxbs
sundzCK5hEZXr6lRHgwgqZYafQ5uidDIOyAdAI+Anj00RnGspYuTU4iLJIi7ySY7546kyP892++S
zPoO+LIUdr7QlW+HDitBBRdIItCZwz4gHvC1KiG1+4rllgzbSjGfIRt3b/JHFAV2krlSg+UaBXfL
JWXreFwIilpr1i52vWF+uziLqIdiwdBhcVpBoitn7sijoNRuqXz/2eADMvovhbGtUxLDtyiipQKl
wjgx7BqHfwAwKAqP3yUjt8j8z3DmSfkRkTQjVpHpNFXiq2p3s1B9EK5PwkefIeGmU02TrlNnw6Vt
WfmqEpWwukL3vIMwQ0zlIX0CM7Rk2YC7xZxSHD8fQKgBK+UllzESzu1VNo+rUFBi/6rWUB+RJ1AP
dgxO5zolp5suBGOAtBSgqVtbog5cKRVcx6Auok9f5pJ9m2VbUclcS10Uf29bDyH7TSw7bsWq2GkV
jRk4/Q5bXj1T15R47/Jb+B5YMShh/deZaFTWQyHlSl7Aw3pGfzJMuIYUQ1/92GB8okZQsHR7Z7AX
RrxkB3PBkaiJuhs1bv87IJifi9Y5+lezPJpPuZH8WkILJwaBK2AlM1EwLvUerKW+Mb2QORwH2nei
Zs2vZHJDl+vjlu/GTmiOutmoRnj4UdEbnr1SGNhEArYXUMKlR+B81dAh1CefT9HnGYEK7yGtv7JO
/08Qxj1IB7JQNctcBWg3HdRp4sswl+eoJMKwQ1AI4+12X3Lv+LR7/mtIlT69c/6R9+6EbTzC6HKs
NEvHUBRsTdEaeJIi+3Bj6HTIwkNEjKpo3lBNtUl8W9B4rSGkGPC3+Kx2losZPXFLpH5marROd8Vi
9TfZd9aY4TwyGDKW06xp+1l1WxIHTFGv0wiK7nVuste4EwBq5KJ1h8TYYrAdImNf6IIW4mK+U6kw
VRqlV2cXxdqDfy0l7coSZrZwT32SN/Ojl4mEd1f9O2luHmh+Sy3+gA5XVJteQmCtohhlFVEHb38Y
f0iDL9PGvYSQri4H0oADrc9CbnFL13gopbl9kLajiR6HOrxncpDsNkCA/SNzT4FzqvzY4NzJ4JkK
gC3+Cj0BEjYQDgnIcHXok8MvKrEJzrdasFq/AuxtH471KUk5QSD1t9wFz/FJgsK4yQWyp6LomYmE
AWuTrl6C8QXLDbCsRJgAAi6LbWIIeshJqon3FbzmNklWnjHjONbEQRMDn4I51hkh9mILPiZQZSpw
Dob+61jiGwd40tX2W2apfwmkZ2TUDjzJT1hgS5fEzSBWpzmDRbFosKF9E930KKRme+RfG+Zne/pF
kQdrHROJeSMH+S2ejBSmy+giOGtKUS0PueGpnR8OhMwTNHvfw7LVs0OMQnnvncEmbs8+PU/wFSy0
VwcTto8cUqN4Hs+7+zI3dyqsEs19cAgWFMBf61GTQrua5hBIznBXpMdtp8P0ZbSmTbrhITzr2qfR
J3+2yWE3M6oVmyIgn8f63YVwgMPYM+jy3+EpqhaOXa5B/u8Fyr5XXCL1N6yEuP7J0mKQvGONF1aT
SiJgIK1CrP0bqVJ5cM9GIELJHeJN1PAcvlVYtejxevN5rzoEyljSFeZD5NnhSk9h0LeNfX0LXG6/
UNdbcbiEa9TtO4n5NSqMZ3wofbJ25tL/UmmK3MoMzQFFxrUKMktj2DIppPNcWV//GlzuXU/Y8jC5
zijgxnZTKQxDlaECKAD1Y8l9cD36nRlcPrQZOX/T7dewkxQ0VJykGFYnZY11sGXFsUEKQdaeqKdA
2RjsqpRBPoDjrKsH92i649xp0fbAdPRmZ0KvPlfLwsj0zmsUO2jrwi8fduy4s0uUz1urpW4PQvpr
I/nR4y1F9FzTojWRVWparw5oT6AMdE2Z069JwzLNn5G/wwoJ2A6jxuTq20UKG2wMBk0EVdV6p3wE
g6e1oJYIxRo9ugqDnnV6hXfyzTUeXQNj4KS3KzrH+nqqXOOhQFf1K7kq3KHAVt3yZIpMtQJoWjMC
fr3T6JCBl4+lTJZtfPJ2e/hzH7z2ebfDhzHiILy5TO4v/QtuYmwbu34nzx2nIO9XMa2pkseZGQnZ
xJIeGpEdf1lBNHorO+yUAnehxGU9wiWz66Z/GzbKkmiMU29UmPbubFvDSV8ZmJ9HaXmYlGsRWdxa
624UFyK+1+hxkXx+U8cH391b5SCZdELJuWiwc6lRtfW9wuTb/aLD7VkveEWGZwv3pVA99JbPmvli
Wb54zGyeKUIHKDH/lySsCwW7w8dBl4SCXUe6DkpIqyd5D7zlkssrRaFkwcGEBDw+accW2dyVFdVg
ARcj7U4WtWhbxNwKfVjNGi6d/3VSh/q9E5dhdx4Iu1KCDZpFSJPdHkOP5aO8hC4LBXgi/rk5yIuU
NUfNT1aVOwawTcOVJ4Xsw1cnt6jn/s2ilG+sqtXZbYimgaGKVP4PStPkYdSYjyn4CLC/oaNOU9gZ
Am+iT9HUyaO2n0hv6+tfb3Ou+ZMq+yGiJZYNGjOOmk5/bJwUaiuNpFOi+Liy+5b0XLr0bulX1ejx
2D94zqkXWfCU/Jx8hENnqCfwXhAOa4gZ6d59yb5HURrJNjLEHlY/kw7bxAuEzto5c4X3FfEiXJPz
EjBrpcV5LqYO1crAZSzj9I1QzkHCwlgjNHd6SWdA+jmi/+ksPi9vwcW2hjJIeXj7SEsqGqxj2Nw/
0ZtFYSfDGVFwWeN9o3E0Aw6OO+psdslieYOTCvV85PnwC5WLgGlqtpeN3zwSj3Uz4Yiwu3PCiLwP
SGLFWMsgbT9209VU3ucJ+9YuONNknC/C1MT/iNqq/jQu3VIjnlQ3StaxLhRIp0jT7rKBlhzC4TiI
+JXkLQ7PjJW3J5NAKGQ8HsRb79wB6bluLylmFJi/FB5auZE8GvsG5wdAlp22j5PgTIZSpCTTsOYt
IZqlnnBA0ZuVQ9RVyxqe3CsCWCGJYaB1D903ISG7xMNDYLNPEHf8LCBiX2E+ylsFviX5//CsGFR8
C1Tey0vXeZ2lCVGuszWYB5kUuC0QLPei+V+6Lyb1z/Z7pasnxWA2v7f+4yc19+XIqmig+PUbMc/s
RUz7ySqK318gwh37Q6sYMJRu2EROIcpK7IgvFyLCJvWw5Iz2T0WnvWUd9IqAq+5RdMMqm+lQRRHQ
XuStDI/gFdqlI+E1XNL+Yog/g3lKPCwavguhe/5B5subm1oVQXeoxLavk48Eeiuq7LrvjB+vabeH
HL6tukgkaQjeQHxJTIWvf0ZOlPGUDVGczoRoTbVMPvI5X2kJu2obDEgWkQ+O91uEbXL+tjMcsE2w
q2oCwrD5rS/3N6mj7LJwKpHXEZs5eYcb6ljXVzM+rcmxC39TjP78BrYpFgxVQtNgmqfToVMPpIQa
9Ku3i/m4LgIm1f69IJWNyFFMoxHcaESzSokB2mnkKcHNdpTvO+9Duqu0Nc2WLfGOXvJJRbqeVs1W
usgjjTrcNo6M7XohFJJsmVFEVV3MYelM6Y4B1TQJd5i1AURNMq6dpai+Zbq2x9hUKZUHHazTt4JH
RnUenOITYwOEsSDhgRhCrWcby7u2GxNWtBqftze2lS3qv+xKtQagZq0xGYnzDTc2vDzUaYxxvlvr
UsQ0IvXG0o+uVdFx+CMe3PVos93jNmVu85f6YoPKlqoDad2kFDn2qp6xPCzlNspOVWQycE8tZvCD
FAd+NUigx1f+TkM0jF5aDuxerCXDYwsmjMxpEp/HHdkNaa5U4UbIwJU/IiPKnO7n9CcUX6Sk4yVk
3VyE+r65zBkMBw9f+lsTkRwD2NPNCHYPX/jE0ehsCHetrmEP0FMoRB9CaFPJ1NLEWy5ElSFdyqcM
uNoIuPqH+DN6LVbyIW7apkKaczc9a6fGiu+XCyyaKraeC0FyeL2/isbiZffckPZWAQBEhsahSgnh
9S1eaD6DfkiK+6ZYD/kMDbh4x8XjeKRf2BjfOd4fsiYooNqZMZLs9QscDaGfaO7Uo+ruTZGdKIpy
WQpt5Utt8/RiTUb6JbubzehnWvNy2rf2HnBJJh1UEdbz6+X+QPc/YNJNfrii7E1JfDF1g3kXIEP4
siu6YMgE8igb/w+zCmaGk+jgJcFiSCm+gT0wSKNqdTx1xBZCwYXSyNZ+KUwdq8+0nOzJCv+vBRjs
J/UeBmf3UVhEoCQZvMe1HdG+GJYYyJbAfSGKIVYNIHJX0nvKPFqVq+i9VvBRZmxxAAuQuFP0hEVN
9HOBnPYXcZcsv2he1dqY650IJldvZkomO0e/PBRQxgALdKP/SH2QU8uetl8EyFy7KNl5ZiASNMXw
lGssiC5a0ObSjpA3VEywjvUPFiko0n7vdOhuJTSseaYbQhoI2KvMZYIHQt2pSqP2w+nL9Xe4Ddvg
vxa7xZ8NwwcX7xBet7qP/0Va7Ti10PyCMB/TkFHof5kD3clUCQX0ULjw5FdD8ZUVpJ0qEa1X34XH
2LrZP6saFWacTstlXyhEzGcy6pNo/vfkNNm83QtfpC3e8Mrc74mTw5GZCZdlgR08JDWIj4ax/86P
+k0iy6+Q054YERfvBgPcSXvNBAPxSxe5AApvvG+nOXYn3Ey8PKuU28utOO3WQDuWHtlieSxAgjG2
sbJCth5iJ1cD3WSEnk/KNVa4PHHsmZsUtyKCOBgZRxtQ7sfA0r3+8fwK/qGxQ845dyojdJ4CY5fl
2lDRuNXpPdE23TalXAPA7gcvXQ49zFkILMtvGGxbmwvzIxAJ4p2juHNYq80Sm1a/SOI1kdfHX8x1
rn5fp+5mUaXKD6yeh78qNub6WZCksYc0pj9rnbyaLSCkYJ0XDXdmEeZ8AMhMMEcu5DHrl4s4WoVk
zQh29966ydHSuJ6qg77Sb14lXpelHPWzZbhcKfIiEV0UAFfM4yaY61VWshT4QE4Kt0o4765c4Ind
CKWyZ1dgp1cEMSgj1gxRTm+dmpnNvKKvbXMuB5j992lFz43zYDZx7djJqbmUqzPYBV7HMzjw8s4p
5UBd8ZTIwVw+Muy8tY6vn2lm07jJLSCagDvDsoBWQj11qv4Vo7HBbmskVkfL5uLN+UgcWJXBq7wr
2vCt1HcYZSHq520UDQ0vi/lEcG98wqxj120c3CB9lbV9za0ZcNQrvgek/BFIDcED54aXtwSXoSpC
9mw06FmTSK79K8ORui6y/OE7pcZQ18DJvOCmP4s7pwsJ4Q/w3JQCg48n6NAdsyoU6DfoMEbXtzZi
CauNH/YCPF4dE9x7CQ2AK1FMRtarI6wzrVXqglPOE9Umq+4zzTAXVqzvBs7VVf67H6mJVkocyrWU
9zkDtbAJfxD+QVq50HjumNwinZdca5SAy663atSlOgTSZhuiw5XJTjkS2ukz9m4qnWDTZ2YVeET+
AEX2UbsUFP/cGIGkOKEZzLcFc5hJn0gDuFfWgnMH+UGU8Taca7FUzFUycQ5dY+d/yJbkxNNYrcXb
er7QiKF57RP+O3DtP/PHPLvBQr8zLNQuApypP3YnrnC//rGG/wl0sfK2FUvcQIbjZS9+/3+US6ez
c5kbknMnzmq2RzB6oe1/298jWzxD25m7M0wXUNkygQUNFk7pNHLjqK4fWr2ezZMSYvOdmMrDiY64
UY5aZj0wo6uK9RQWVG6QuCEejd1QNrF2F8PFWuZ6UE5t/87WOFAZVFBL27ewSnrOyxAyNGj+EatE
kiRxcZ1P836sLcGDZWBaDZW9dfq/FM3Hj6SAvtu1fgNGsvKat56mZbxewEPZgH3+cgi/FCmxtlyt
0tX50nvNeo/A3i20u8fjqiRfkCRGcbbgVfGdHtoyEsZXSf/EBrrlSFP+ukiP2iaPrZEURX+EbCo4
/dBLx9GBPhrMfb3N6v6FsWOyXbqJGChZ0TQiGG/r3cvYOZ6V9l694t4zJRZKEZz8NFSUjKsU20Ce
75K+KZOyy4BqIbMjaRqK+5872oMBTncr7T08z0Qgd36awmmXI5KDqB2q9opEM/53DnKkLBsnMxiA
dTF2nqBM54/qB/8/IHokf95dPA7Xan5ozPdsMNsl+ICLYOy8Ck4wee9eIe//8W/zfo29vtdkPfWU
Dn+ZVfxVyYufkNbDKqoeDRPBcoCMZnInPQHVxcpvphZgItFc4Uj2tAH1nSK7j1YCSt8VDls18CWn
dw9IMQfdP6/5BJi4LFqc5B6HCnbS7IYEfyumSsz2iG+sFPYdDW0eA8L9DQVWdHP14HeobBGGWx03
YF6JQJGxnYBGhIzrdexTc+ZJt3TK9e8Afa6btEEixf0r0oyZWQMhYV6WVH0EbhiLoKwZZ2sQ5Vqg
NgOm2DkoQAY8uVcJr8SoIL/FMSonQjwJsRLefrAoSaJ5vG9Kxt+YUoRhdUaMcAIHI5GHRDu8kJQE
H+WwQhv/l9vWFb2BEh572jxCjf6/ZOvN2Wmq79EZfuNOaEO+iSvnhk70RbC+oDE1G0yeaTEm0rZM
Q+a3gJUsUekXQSLjNipWJOdfyL21yvmwboUf4WVvHJedZoVdN1TwK5PyGcBegfkQC7/85i2MHS1q
d6KirMN6Bbe/B8GauZYIag6JH9VVtSHxXKpItG12YlpRJTHUkNAKhMYF/IM/oj+gYaRKdvHRlC/v
KUbLwOHf/xQtIwLCcP5sWAMPUHk56iqz5vByKOFRUUbgHTJAdeZE0KfssQBcGgwCk8VNvLGcVis6
mwQNeCcLlUUDM8wrVc9uMYJNFm1iCSI2JzjjV1FWF5aUDAVHbE67qVcB73yJLvotkEH4+SThMOsz
PjZTxAGvIIXxX9DQ9i2C5Q/hULcwMm0EooiQmJq5OVP2ZMwBQ8wi8wSWrJw6vvbcpGGFwI2dZ6Mt
6ZgNlYkfMdsDksFuBZFtnxH5VJVUCVGik7fqipFdEfP0UKTKJWyTF+kwP3WdLUhtM002EUjdI28v
fRiutipN5EnOOHWB07JgbOF9ztoMpvU8xph1mVUHEZGsGiEumFM3U7OS7Q3RtzDzQp9DqlF/Cxzu
qrxADv9kFhMyfoGiMb5qQlBMu22YcMo3rBmhOcekDsyPcaTbce3BfueNG7AUhZz7WU1/0hfXo7RZ
bu6C6zec2wzhISi8Bco1ms8dmqm4Dn3Gj1NAYZVHq+4Ird5UYrg/No4hJN5pPW+zP9TH9sS/MpBS
V9WsVZl7fq5mzzU/TqYtz6yrkt6QcwxewOIEhzYRTiqFaWVhlO01wjmI2aiJ1c/OLOTnNoU2Fq3b
Go3ldxGD76l9bWCJmj50pi4D7GWetiAiYnnCrNLAQhVU2cghq9sacc8RsAyZNaqU3I18NBfM9gJ9
hPwc1Aae2GzyEV9qO6xrENkDfevQfGpu9z1jvOUMbmUHi4SBNWR24L4Fp5Bku/IHlPaivxxrJEwD
YtCIPWZDBLStj6pXf/f27oasy0NjN4miDhSFeMf36zTHXTagXEl5U5dYAl9VyimploMjexTLHDjB
ZDmrC0/BCsTBrOn1npnK2ZcE838MNUYg5yC5aL07vigwxcrBSK0m79pg+bAfra5yieugQJf2l93r
vEz4AyFwBPqtTi0pnHDhbDDqji+itTujfNE8jotKbl1eDaxdADrqb+lf2JKNuqCN//cikfAECt5J
SCA06yIlx7zdzJBz5EvVUGTLGnOI1F/q+jjyvIqyjImM259eG/V4Z9CiFK4ZJvjKOejjFSt/P/9Z
8o9U82CnNCK4TzS8lCqWL4fauCRHrYkU1qu+ZQ23KU5841VnOB+sOWhdPH2i0VxmxhR2uGJfmXYJ
bbfRVg3pDqfkDJ0RkRcn4oeMai0EwPCHbnadwKZfkzghVDiPtFbIkzD7LN/GWfYfbsBbTE4PHy1F
XFT7AdziVo0g4xBzkb8nupVIO/k9IiTEmSmfkFxV9uuircUBGqeLNQh+5hVQ1AKpDuKz9gjz00gu
2FRNFyqnMvsVLN40k4M8pQKbuwffzD3pgstXHK9Rk8gBLrJoDg6Cwo8D1kROpxXPnOhNKFyor2LD
QUC/U0emRIOEEK0b56vSUkc18zJTVkwVU2qC3Sa4dmfUco6JHRJPkQBKuM/iqCZZsP/MR5yIGN4I
q+SOEmvlLUiTVq+6xZ31dmQKKtZXuZfzUJx8MkF4K4Lm78uRdSL38Eulo+GsDycIp8IKPtrisPCX
llF2Pg7drbuF1L0sq1B0m/Om6q3ApIT3QZFS8d83LXSo9IHEecUhw+7S0RLWKqohfvgw4eLYANij
EMD0Xixg7PJigE5hmod5tWTekYGS0gPFDox2XupG8pqISNw3hhSB0iypew8ByAvDBWKQwlwQyRxL
z/+abh44797IJOkCla00S7qMParz4H6N+YNOYzq0I1Mm+h18UxpDo/pu1kENi0rgtfRVPJk+fVZy
0PBlEsRVmS7jyioYDLz1km6nNBeAx1Lg2EXpQnSuIyncOv3GFugQpZtkwvNd9AHA4R8xN+l3QPdb
ReDxlywHCFrqVo6EtmrUObZ6x8v/YOCXt8ZZKPofT5/xSOzaBQ1+nqXuhayqghFxG5dm5tVJktLG
7CTZB9rYQPEhAPbBItNEhk+QOpbH84CqPtc6byJVtjx3NrMDRANrUEhOEAqz3oMPAruTZeSj8a+u
DFYiMOlOdg34WS0WKFeBavlLy5YPs28H/chDtHtQQ5kQhk/NSuunuLvUF2CajJy5F0WsObNljLQB
zAGj1U65VGBFBOae7we3aOgaT0gnRP44ekhceobigQ1qQTOxa7fA6IW80EQO6ELujb34aWdZl0N/
bPo42S1CRTNWUOVD9U/QDA07NdHha0Ua4USjtz3ZpD83wwKBmw8payS+YqDKajMp6tdc8y+HjIFM
S6nJ0sviSnHEe9xZaUHpoVzsxZtQae683IJCWlKDOBFpsz9POTabK7KLHQ+/rnCTpJo3wqhoGVBu
wMMgPfHI7fdiY+bbAkt0G6fwAWcRGOsBn3Fu/6WjBRO+tbaOS3qVKvAZ8CtpPqxqnzR/HVaV8nhi
+BeuG6cuAZUsy0HFu1SQb87UZ1uAKXPv1qbkAQlhp1FML6AhTWv1idJcuPDP6ACGDiNc8wxQ+ZTF
u++jIXvUC3wWIhEJSxkVonMmyBeBULj6rOSaBB1IjYjDMnGafdDjYIaMJD8Awq0dliWuXLneAUgY
ecGLfmcEfSLAItJGsXqiXQigwiPofghmykLutuYF1uOkjTP97d5g8PTsJCkYfXvtenvkHSkayeIo
jqHHijXBhrc5kKsE3l1Vuk6Q/i33ZiOAFgesENBiWCwR5swHgxuwnu6jduqJUq94GU20fI6Do6uW
pU56rGgLrMgdPdnIqxzjZZXdWikLiZwA4div1OnQaMFQxG59OLEU/6Y3ZsRlZbeLGYdNBo7kqVxY
TU33vSVCE/aPAGtR1cj+GzEvKpgwENcb98kam39swackOiWm1wndd7oywg4UkK/Xwvs6LD6Oe8kJ
/W+tWa1qcl/EMkKk1L4MOD8/wZb16nNygGtQhsjJMIeyabRo/bO3G6CfysZ+gjDNagecI9b5sZy5
FbF+1X3vPpCXRgA+AMtWtbv9Bg09OjlX8Im1UkONUXA9ih9plPtcuuk919pkeppVZy+1Kphi7yb9
TrV6Ub7qlG3IGSalQe+mBtt+DBB+m5Qzx9ujXD2QfFV0Oy+Mem8rNkO9awZQKCdnzvK0BcpihScq
2agwKE4C2dlUyUEdoNSEPTYRtk67jnZyFw+pPJ7IbzkzFI/Uh92sBKKX0ExMTISzvR4dxz5oMJsh
REMyv6inp9MV5AA+pNE50dLd99AjKt63dSF5uGYqR8trD+UFiQnRJxvJB01ggzpxtzITYj3p3E6+
wgWWpuFT6Lhz/UNJQx1Cjjqbs52IbbgyxowKDZ3+Qk3vzSHH8dKgvD/DDeboLhKjwhN9GNknbj0J
65imHDVqxzpStuVKps2ir1qtE7jMPLrh+JlZn+ZFlGE/4dNoX/2AhKe561e2g4XkEbeaX+vIKR82
j185+sO2NNgJ6j0EOaoD91SXdGhHg4VCP7SV3x6r/80SDZYOb+Q/X1h9CPqyOMrzFZDWH37eIX2b
MQJADw6t6kF+ZhynxqGdBgw0J+EAyB1/LJ1kqyTA9RmQYkcI/2KywUih8wttqX+yEcr8XR7giPCi
vys5mqiD4jRrsLNuW5vJ8nRg89YbYD2WmUu0p4u0v6rVVgCF7JeJSuCotis4XvqBkvVk+5EjLrO7
Oa8jEmbuZuIpDyGMWOoMQUNnQdvC529u8I/vL5FcF41KHet7T4uVD0jjrkFDHG77XTRnuM6/D/tg
xLYNrwcWqzpwMvE/T12+JD3/BCrEbse8nM83sPP8FPV8EAbaEJ4X4qD4xtUc57y65fE50HpakSDj
Ep676M2Cr606qNEJI9CBg21B/1w8KPzKqUGeIrROVIP2jlnt1uxDDeCbAPbg/X2A5BRSHIoijc9L
LXvMBAWe6J0Hq05Xyv9GBSBMk2+ww4TN8oWY7RHuI8SjvrrSOGocLXND1qrP6FCF+kioWsiTOYVI
WHu7+e1Sky69MI0/cSXeehUQKSFrJ9vMfu36KX1biDuGI/KTQASc7LJExa6ZiFmq58aji+y8f9wR
lI6hM0BuZRerIxxRidYi6rLLvOXheo7bDsNI0eT6I2EtpsyTju8v2pTSoVyjlsp13utjh4OGRigM
VlvZFe70kmWYoxCexVZEAhQxDoB6EVenGiBOcOkEkbDgxep6mGFFyJxiVOoG2adOEfuK8QSu6a+g
LB+XGcE2FclSau1r/aIw1/3SqVEDDN41UXtB1bwWYhdBRHdD2Mi6TMRy8IJhuxosowLqsn9oUlcr
Vf0ejh+uJik/CF44RLra2fs3H8AcM8jEJ4GvNqIuYu/HrH7+3/ZYi+mQlkS6WhXmiTnPHFgAKPlv
0Ul0OFKE4j3K6tT9y5C5ofubo7F/WxoCCskuUVWOQg4J+J8UkKYKh7869ETY95uMA5YLy3dWjnsw
kQHa/EYciJjG5NeZWaoytKMiiwVyEi39movqgHTmvcMfbpkd5+dYy/igMGIUFqVQXlRpgAu4No5l
t47L9tGHPTBNiJa6nwi5b+tKrJ93e4MVzAWYuKvFxFnBcdXZXtemNzD1bTIVLVIAnDjdAwzTAVDV
8293/kjXn5QknHG1IyCkbxdpJ8ziIhbI1evRCkPk1lzwzmz/RuFTgfhmq/+CIGjlg6sYscUINT0z
fzdtq4cLaRDTNZTjIcBcajcfB0N1GNtpKCO/+CjMZfiTv2bmGwds6dw57X7Vcio52QaJgbcvr5r+
zyZajsARAd73a5LKt1N4uKKuCSArYgGaokkR0stDmwk5wumvYOO7goVd2GregySngrXPXJxmzt0c
Od52ci7yaaMrPZxYvRWEmnFyk0OfxaazOKz03a79GEJwSel+UlAp42y60RZwhtG4r8A02Tlg+Vgm
TUOgUxIreILNdMajA/R2t/Goh4/mLyaqGP19cISWapIWLlxvn7d4mzN2jqNV1vwTYkGUzU70oUI6
6MnknVrVu5JFQqkEyy0t+J+z4li6NtL9ZtNCMwqxfhmKUhBQE9S8gzeX4XqHIVJH/rFydojUB8XQ
TAdPIwD8E4VxHX8Rv9Jaw92VAk7oWuzhP1TczoEusLXtsuhwRtMsKoezvsqDaxSYxNgS+XuEA16a
np8NM9kQ2T2mYxCe/nfkvRXyAQj2LzYsjjRXS8CVxClNLKxw++YEfElwJ2/cLnV9ip3Dku1+bdXA
edn7u+3uiKqtFtwFdYR2C6LvSLxwCCMtHx0Uh86qiKg2gdDaKDv3vLZuys5pz8siNEwbaE4rQTOk
eNpintu8PJ670kbjZNCeFEeRmTsIHoJNhXTvhb1iqqbwc9r4qOPkxS8d6q7qICmxhpo5E21QSNst
xqKs/nRYXhzeGtsTbT9TKdp5iZskS9bMEFHXM2SY5XdmOafJVJxmTNLMpcVxkneHRbL3cz4D7Nlq
IYDeg99+kyHnU0uHSHalywYQ8fcW/Jv5AAxQLZxKX/cMpZVbVy9s2KYn3Jn+OTLvsKYSQZrtixfr
RTl8WhZeqh/VLSqyCwtwIHzIfpQJYmFKnGUrT+kbtOynxoVEzZhpp7g4KRlBN/pqh45hNN8QLCuF
/9lcObWPQeN3GifQxEe9KaCLwGEnFLOZ+PUJlpVJeXNjLH9k/mYVF2RTsw8etti26KvdKQ7P4d4a
hzpFvlUwsDqwC1Nh0qTSyJJWDu2ynT8Jp+N3adt9URxED568yrc3s8eNR/Ck/cn3604QTjPxhANv
I04qYSUZu8BTS3HukEJ1O+esW0BPKVSs4hE6vlVFnDhoszlmIL5PtaYrPX/UhKKaKBleoB/hB7tH
dUMOo7h/nfnklRRI299xV2CzJXd+NSZQug0PtefKo7lkT5bbsxzgUTsKpz/UgOR6ctRRqcb11G4z
S+WS/cDB9e3uVPAKoC5hBqhHjDhPFKGM9g4Lj239ozdWowul6gc/zoDbeysItGTF4Nas/M/Npk4t
NXaXyPQ4eLGpG7RuAo1sJ7gW4bFrSvrYegNgmebHD+5j2o7lrldAcYO39T+8YDCOwIwFlj5Iu8sT
3E6Yldmz+mgsSBXmIKvO3/X+slWtbtDkPIs51d/JP/vmExxewa5LcLegb1ZpcJluHYHY3qX40Kop
akyGeY2tHoPd7NuXAuovr3M6Z86VeV8BK7PnbLBFG5M8CWd0OQHa81nc2Cen3C4FBIO0M6L1twt2
7KQGwP5/rL3pPOEqX/2p3k8hADKuPVooZijTV2ip6AA4Blwx07qJMfeafp/V9iaoSX/ACyFE4QcJ
PjWCDYcxDb7+81PHf1HTIJETdoTPXHUF1SXZBGT4qkMpV1oW4nVoPcDJEH1BBEKs2QSfOl2ykhA3
UCzJyyuqi8Wokx5HhjIUYnmiZBjvrvCs4cXYJKrX6fFe1tjB/1M3bRDe4tK9BVI6Ksk/XdQBZddg
S0gxg19UoBH94q6L+5PoogPRJf0hE3LboFEJCb24iT6SskVzIJ8fcnnz15bb0bIx3gxojPm3Jlte
CMYPdkbWwsbT5wUJeSRFfMTb86KI2DMxVmaLdlS3ZY2lALgutdjJiXpHVZByyhMhy6lP4MHuO/nZ
pgXw53cLuGyP0+dX+Cz1WUjq0I4D9hL8IggmgjvHIC3tFDZhpynB78Uir8aBiR6JmasudDwcNk8y
dJnmh7jIoCfLEHPnynxxm0Gxl3ArUD3vmwhXyBQIl3FUahxz6Ap6LZnBTx04Y7TuroWc84b/gsQT
gpJQqk4lBnzL5LeHszLweyJjRg1+hV8odEpiGFDDEZXmkswdkqnSNjtI9+rLzh5R+RyrCdGv9q2v
Y2fvcQOMhRy/aud55JmDvoB4+NGdPDJRbr2VzuNr6OFXN6XCpO+KE/5Z//oapHn9DjV6jbEn4zHR
uli3cpSTcYXI0BcB/BIFolyycrxKZPwR58Xz76eBdbfYt5GK1gmvWuP6d1eo71+AC+EX5KEYB6Rr
EOP9m8i+wX3DGmu0W3nPH63LpXUlR4Mfgh3pk0mCJyyx41qsZk88RrLEOdYGGxMFf2RYc7y8Dxbv
Y8YZOjFbflf0DwJ4idBCSS1aUzmMiDnBE+a0HtqtemsiunUTUa2BsUBwaElk+qQZRMjwPgvzxmfJ
Y1A170LtUIdweePor4Woq9jj8epiloyZ9huUHaIoeV7n5Sa84tLbB7Pb+6kIky7YTe7BbmvB4m/G
LZwvUBDQ47tS/laxTqOIdRLNePo5pyEJglpwhypypLE2jqbqRPdQMcWiOnefulmTWXL34prOoag/
ZpOq5U14CBGnrnl7vfyleI/AXsxZAjNKvx7ctdJpOnWLJNp0dHjWgAUxfhc+xfVH36JFDua2WWzi
ymbD58XrNX1Pz6Y8xcJ7/+fm2QcHUtq7kYHYbd5aFzUdOLtWz+S6A1M5m3pDANcglsOwYIwQn4Ja
ZojgkSY3fU4XujST45YzFN78DQJXlJ1eGhJYyqcnJfJ8hfUmm8BZT18Qh0jtQOHROCHlcwSWxcwL
Q0vXPSLtzjy/qNbiW2wl6eJOQZnnW34mLizMRuJYnY93xLiZr7RcAzJ2KkjeY0sHtIZF/gOVnFlK
EqMx6BJ5CsCQ1JCLb7u9OWr1lzNec/fqtzCz2xvyJFch0521eUy52sQjdqoApfKEF3pxvnkUl6kg
WCdX3Py9yb2x1CqJOhUClDEgBagYzi8YYwOCBk2C0oGiDTbC/yfUWy2TeKblM98kXtQLuu+muIxQ
DI0rDb6A8p82mKFULeeHLDXwCN2cf7bEkDTKPZtw0fgX5O+v3BixXzDj/YyM34NsrxLQcJ9ZVHi5
DzssuGtf736SCb9VmgIIBYjpC/hkQZao1mq+w+WbRBKrG8vyd0iPDX9Lze3JGB7N8tzyYU5ChU54
nNxzKejezkQ9MWz2NxoaOp5IO5lcdCMuUwiSC/JtmMP52CbIK4XTPlylVc7DolcZeWd+v6xCoCHs
mUOejVHUfbsEJA3b0N6WD4ovnSUuUnVYo45aZH7NkZnyXjYYxIwKCTUc92ZB3ocXOQnzq/UbdwX3
HYvvgD75tQzukZ8d5/utfR4n2fi+Ab9KHHIGYa0h3ii1ZIrp1qJGPfjIV3gpEHb2YKTC+7OdHEwB
1hAESXGyb0vnJbaFih4z6R+bTNcIKeh9c3GzipDA9KGE9LHyg2sx/Y512IimXBSGlFb7+Fsu0Xzi
PVkvr/DjPudfqmWcSswUdwS7OM13LfwlyPfE8TlUywR3Z83s7+wCQ3zuAy356uDr5wg6Bl8do3P8
PwlVeEOrR12C2xk4UFKto2bltiOOSXjAQqXgM6OWykClbaE6B5qruz0u6CLNaDOxpCQHqAUXRVKO
GRSR71JHEKWZ8SlFpeqYh9CiHupFP+E7evvBWzmS7735JIbbDigjtJUSiboTXewsFUiLjZErYtLO
4S49khqvYYZgYhd2SXtNGsRyAPxryAPWDygHNRMshL36CyHLNiyYCzl/pin/KAZqeGz8fdkKUVrw
i6PDvYsvdxmiKWkkm91kbmyXn9KDVXJi/OHV9nIl4KD1W3yOQBjb78T0a/ebMigsYOfYCSCJg/Iw
GdCN4+2+p8JM4lJeKqKEDVNhEHo/Iy1CceReRmJwBG+02eywBU6lSzUAc2HcvozInI6R7ir83tNO
KRPF1JXAvCgsdOR0Xro2TRkG2xI3CCnr1snMCuFqKO+/IEUVX7LtrVwEgfb74Q50Jd5Q5WEnRUYu
7/R1MG21dbbY4uXaOG+jaUKVs88e2yDo6YiHvNMPq4C+iiOU/oJTOtbQNNT6YJZF+WvIariDvbs6
5/2SCAXBF+2pQb37YUrTU4rgBDoQyTrU8qlENTQvlxcxoVzysjElmVhsQ9QHNoAxO8zSIkrN3n7V
LetM+PGQXEmlTVszzWqrjRvfZ/IpsqhBHZ+gMGWegEF+I0A0nVtZo+s8hmgxqNZMUdUnTCMPyAkb
SKI5zqOUeyHjfMGZph6dl3U54D8rBvYGaXTw3rWOs4tP5KPzxoz2wBFk2CSupG6v2P0Z5x3lAnqw
9bGv1IxdUoSIHDMCRmxAiMc/b0PkxUmVVFWil5+f0Hz8TIu/G9XU12foIgC2+QtDyTM1d2xXdYuy
Z50Ik0v1O4xcPDZL5yq7TCr4G7OQb5SqipbqPxpAIrUXxT3qtWOZxk7AGzCIxVnBjwGr5/q3SIRW
gJf7sdwZt+xdIy+D+E3RmL0DTlAR752oahwgqZn1quw1JCrcH8+XCUAV+isJr95WHqiicv60xrly
/o1IKFQvbHtruydJs0qBki4dYxKF4g/WoAkEfCJyaYa7BEkSHp9+KDT5iwRsBO1/iOCJbvJexJiO
B27GpHZmhlPNjfpVhw3gL4CnKNvzFqAK45mcKO2kJj4/VhkoY5eUuzNu1BzDHBR3exIC2eSg4Rxc
FHyj7EQ75W0iQ/b9oPAN7FHF/hF6hXeAgF3jbBISt2c2e8iun/0Oacr7JJJ2SexmlD7uhxNlluW5
sNd/A5u0o/GEorPOlDxDvA7Vl5W58aMw5Pmnjq2c7ko0Wwtwqa97gIa9IbBP5Ed/i9v3uMdDMfra
uqsXEiqRjxs0QzC8eNxhLw3YHzNI49U7m1pDHFKvN/pM6Cx/uXnaT2zMEn6TauVnCrNrDsEKRWEA
vpPdp43cHoJOSswHKXBYiQlr0vV2PE+jd1oKe5r3rJtVZ5Lh4OdU9z997ABVV6/KVLQ4VgmI3ZcI
m6Saa7Y89BSVLK8VpGjzx1cZaMY4bDywkKj48Z2Q9ZdsxCyltuBtHTNkRdHbO0Ys+9WpKHnjKTGG
Fnj7cPj1VGuDs3uOHqLbutWd87ZN4RoB6UABYbMoy20J6tmuxpp+iEU6gPux3Wj5MGbOuq1amfA1
6a0b4l0+X9D2fyNygOsbCWNPFfNkax7ZFRREuKzVmNtOOmzFm3/rSGb5URi6H6mg8m6eUovoum/z
4pSFY07RPV8ZGhjq1HdGnP9uRREhbqNmD/zDJUrdDWnlvjzuONxpa5f8ByXrr3oOX2VXUK+hEahY
7AqJWn617vsi0nww8lqAdzlFp39tp2tF2cPzoCAcVhPe571ZibCHlAMbDd59n/sWKbGvtDyCNzI1
A0VXRoOdigdorzNgCAtqzVs9Wv4yTELNSaoRm+P0HlyCNqnLHqkCluR3DHhNmgUImp75jNdFJX8H
wYp6M5JFfeeZkylNoUU0TPHMmc4XntrjzA+i5owCrFcO/GHDHkLUSuET0pK6vZBajd/fcAD3Ar5t
vb4vf64FyiCG+Qe4SL+vog8qq8T9WY4vT2btFB7Zi0E3db9H6LtkxEgQLEeblru/anarDr88Fblr
sfw3CFJG3XXCGFJ6SzFZ0LVJnvVd4vOxjbGRiV/gD5Nq8KnUaO02hcW9SScu6O4GW8jx/HcIcc6M
TRRAnBvaN7Y4IW2vFEctXfa3OvkuxLTSxB4m55aGaa2JcnoMCGSW/Y4iXTQYwuFrQo4REybVGiJU
qiYs3n0sL+r6bzS+zLOr5xYgWCVtY381rtsXEKttgdiRXEYAeJOhj37QdXoPK2NQwd2rkM4Gb6Ay
flbO+nAZe92bkfXn1rFQNjK4EXfmrYY3nqxSQrAby0rvy/bZ2UziENQwTMo057tsVme+GljwCnhJ
dxHhAiwYGgWSqf4aZov+sdSaxp+l5dRs3ZX4O+Kc8Ec31eC2hh1FfEQYayM2u6bCByKp6fOEpCVI
edzAdGTGB1AayaoSFLhc2D7FfoCMdoPjVgqaaB08ODvtypPAgKEhDXTSsF3GpiCiDWJ/Ny6R6tMN
v/KOD/+AWG7utj46QGm8LR7DKrd8MfspVmtvVUtF9clOTArNt7aq7u8hgg6aXjyRJU9cMqlvEeo1
GkRhDJoXOSLBjiZnZYTEM+ewpW6qymwTQwASmod6VV3bQbgDGqoxbZbsNCrPEoS6GGCizlfzLgv1
ipc4Np6UCNknIXrlaiqg7/x3gLhWMaGvu/Ed0l/EU2NZxnWbHHo6TRwVnvyahsxYSJnw99zJDlTe
ohynpzU29vy4XoB0cyrYX6lAzuigWEWDKg0mbdn/DDgEnDFhlGWY8O7ZV5Qeomg3sW2dTE45ugnS
FFf8VxTqFD6ziybDUYqTKg9j94Wg3khh8aRu3cz0sOV5hq77GTtbCTU/nch3QL18mso4WPIcNvZl
2cCKkZ3GReJZ9UCiZV8DAKHGtdv2p4tVXtg07c5tJ8crujac5y9ZcfekxIhbhEA1GUeYZayqdfLH
wFKEmRIi20h/XQRFNEr8tbMDwgsAKj0HX679uT4MELjvqsu9hIuF7WPcnVsTQ31RDvDQ8HCDTI7m
qbjpSi6m8VI2ZDfL9uk4tIzt/lWT38t8OIwQ1BgU/4P61B+7qXSB/BEGfqdLpcvMHqZULqzzfHHw
GePVuBJFtZL0jwrtN+KUQza3nYWmcPwOTRADfq3yKm/iVtA0A8bKRLmcE65RDfYu4+VConWbZrCH
afCQMEkuMsMYBcbMPjIWFerj0wpTxbeJUUMR1xu3jHNgar37gNXOzzoS5WX1hEr9dEl7jfr565cK
0nTjVi7qHqIvMF23Z768pQRDfEgHRuMatFQJ39ub+ct9DpbNQgPacQJemNxmyxZrwi8puXL9jeml
M1DcbWFlberL/n35Vgnm7OB0w0lwYnsMLPW2jwJE1temlp9t98Q1mlcLzLQghkXcX1v9TK0nQdKn
o1HSdOXWtgNXXJA5XLJuAROxzZKdwb+PnbiLw7MNAIu+NiTeNG+Z2U8eryKlsBqvfrZ7/BXIf7ct
q152U0CM/Ma8QicmvR/qyz8H5qtsy6N+0xricLYkOjOZqEnQLuffI6luNFf4k8gfaoB0bLcClWhe
uYDQrOpT22QypN1JnvZFr5S/wtfwPCisMrTMDZMKKFmDluesJhv+1XxJkijk7Yc9oonCCgRJOxNX
9J9gNigsFFOSOVdWw0ZdTSpCA5emwAcxouttzc4vBI9UD4Uj5t1QvwW8JcdUqPB0ymGaQNqDSzG7
lLTktEj2mBw3S7f52ENWGqBTraoIgXFg/P8XF19joX1MHDsNS6Ihq2t6YHVdPUhS5NvP2Z9q6ovy
tpH/64iEU4rsCMVMipRQ1xOij7e9l8cB9taaBVGOOCCljo1JzIcDhjU2tfsQIJkePwuYiBY8tRFH
mFd0L5PaKqyUfgxdeI69cJc0m1TFz2hog2ufoUU6iYvXHtey813b6lXDpfq685JOgE38gw020Gjh
GrMZoNqHQE66aNxFyYTrbMifr82SidpgVGwUbRWUFORBo0rLp2nM5Si6jbQmdNJnUxF94Kh/XFKq
mVffcJMA7AI5CeH2fQaamLOgtrvnNYRq9b2FF7PvUDa4zny7ZB32Xmq8OgTqxxGuJ9oVgeoS72Uy
W3mXoVpfPYvlLvAYO41L6y5WpI43QsIBbgEgLhDovaU+doVSWZ9EQ8Pml/ch9Ef1lCFs5DpoZOBw
rR5z7BinZDIRyxAoOaSyif8MWRdgi5KtQv8o71Ymjvfw2g62aD+RLJQSyt2Xd/ChnbUiAuHL9BtD
ynbPWSF2NU7rKIsH8pmDSMf0Zehv/EYtqUCATBgaT7OxT2cdH3XQ3whrNhSCX2vGneBJgdunwFui
yYFbFCd5JAxrzi4fUnqUMV+ZRE7ZMCDiUPTzHqtJpDo5xVLBuVt0kThfaWmQV4QGZxmlwPCd810e
EBGaQ/C58Hcn/c6XfLwQbZj2bIw95FaWERmAN90Dt3M9Cz4dZbCLmPRuqOy8Y2ej8IBKnAq/KFK/
Y9u+3wxeoBFzciHFK12TWMGWVIjVtonNrOz/ri49hINmMqrfe+JdLPHXRPxgJbTbyaKQ3rBqF9Sg
IJiPGwxJ8DmlrgBf6TGCaClXZ1l6omU+6IM1HEs986KpHK8qBYko3zDKVBF/NU6RwNFE+hciIMDI
Wynfe+UpvhOiBmS/RQhQiLIlqEGU4ePR82pK7ayuA6NLVvgkW5aZnlzdKXTMIV/NlwyGeiNZxvsC
WXPsSFNAq745QHUPUlzuXV6Leu6lAYcibyqlCqwR5sZWdU6BnQOuZB7HnFtlk6potSwUBMDnwBVP
tJyR3aJaPDBd720/5hXPkjJUGPM3qVbN20eHzubpO7YPOSvWeZtriz5uhERY0DlaPjdEUFzcm/Pf
GnV2TNuEOafg2rXcTtB2Ey+a+UJTgA1stEB1hSZTN8UmVel6ZOzp1lOC42BM2WosI9KbxhCV5zzz
p8AylZ4u9DvMOR1gU5Jhzzlqkny6HuI3Wk5oC97ulBvfddyGh5zKzEmWklnUXr724gyFuG60cfga
3V2gjKUa2ENcTJNkPmXE9/9f6J4apkjTUm0m477F7yQQ/RhZjI8l0DUOixpFJ2jHpBZ/LrH3mtn/
yQP3Q0DADmHCx6j/BIVO/LNiIvnCVBYzHau13dkqhy6jpjl0skVsVFg7KHQxu7X3OvVTdjnnuiYV
bfSc/X/yZKF3DPGQVm8fnpjauaanw+sL2iYXOYtFmOxAy3aS3nD7h4O0JdIdFG2Bu7DNLFTCzFAY
MZtfqT6NcYdul00Ixqkqc+w3dVWDtrdjgAwhRuUVtM9S/7go7oxjH/WPpwNaU4BniO9VGT9qO8wk
KzsRy0YhBSK9+AP2rLek5L63PuoTw9FtvsJl6UnIbJAu91XIQvXd0Lc9pfuQMOaSjDqwmMrs73xU
ToBx/ANyREPMSY3wvOAEWtUO3J7HIwRwT5NZTMs59nUFcClgh1KANFNYN8ZeIzPXGYWnzRBMf+mj
FGpBqJx86ilwxjuMo6r7nPgt11L0dB30U4V52IcPqZKySbtWyr/f3ejsgubYFQ6DbSOzADQc1czB
nX6bbUh+/4IOO1qzV7RKspRgozHft8hLgNjXdI4H/pBnJYFOtJlMMOpiNPLgyIjP+RrUWCyxssOZ
JSS+vawpP2FUDnBeE8cj+Jcy470nJW9N5r6ALlmzzD80GWTTMNd1QVnct81D2gAJIoKgwit5SljQ
ZgEmGvXuomGaAJufYepHEJN8itI3rF+lLxz5HLe6FcJ5kkcTM35jUreKgrvuTG/OZdnj6T8QNdPo
YAcQCUOsrh+UHYHxSDHsxiNIxjm2tqRPjSs+3pLDaDV9AjIoQCskA60tif9VBcLG3vJ/66r2gwmR
LBcntiuiTL9Bn8d9l6YQ9MZu9+ZP16Cmf2k2Q516IAIBql9G1wl61F3YX20Ubay33fh04A7+Jfgv
tQVXgI0wbhV1HUhqzOiaoiCrg9sLIyAv/iRuFNKg+LRijf1yJ2H4f6he3TyK1HU54PNv1cgQVYo7
553630oUCy96DwHv38VkeHbX/Wnu4yHSV1sBvpd4mfSyk7VD25N0Wly84OLsgDBWA7wEDgLz6ttY
BgQGkWxAkLypjakqIGXRW8LSqXWWfkUxJDIde/ICQYmzOQMiSy0U0O8YX3Hy8WyMPkwo8HYy2J4k
05vwL331a7F1fVrYzRAzY55qzp/05oJu1wCEiJ5Q3jKvPNpVMmKfbPLZt3uu4BlOAIwOHWEycsjr
JvhSQh7fNVmladscoqkoFhdpXbezljblATVnVv1CIeGgwdnDuzZQtLVqtvyAAZFtTZXpvjAO5TnR
qO/S43sqRZrZvxy/0tdVEUHzjALqo37vCdbjxqhAiulwA9vsB9PhraChgyJBYhJehBihN/Q3NLML
FT/A2xI/3WrZMpZrAc5HhniBQ2Q+V7BKnbMuXrF1OHl9GVMRpeRW+xCgJCl1ulCtHrUKL3QpZmkE
WA/d39vKN5CBDzY4urqRdmd8IlXRRD07lbPiYNLsS21rPKxpzEH/j7fn6xJQIHGWmfceqY81HFSM
aJxOxN7bX2KETd7x3uwG5qgKf5QGi79oh5xnrZ0rapaq46qtjuFVOuXO30BXY0F3wIQOtJbMHiwn
wo/+9IZH1PsRH4D9UOfTnR77fuh2RVZccmdajtKqOAFrie4yqYfy4UrzxwbVRKUFCl8HaiaTodhc
0vxZUSkk+4QjwLG1WodwFfhaGz0N3GU/IAwp9UtJIyr16jC81FJC8X9TQwUattsmNcv/k3V80+rw
iHxdIc4eDSv9ZDznM/TWKGLI2NHfleJuSnYh7jGpFHNgW5TgJs+2e2mPJjkfqGemKW5CDeYxwhVD
NkxQ9IjGkYZ9BEgajVBfR9Wi+YQaAP12mTTQffUxVnmISuvxKkDa3VwWaIKujgxFy11qKV8R5Zm4
MzFCkIh99t8eW76sWsYmDVaNPdbJ5L/ii5fgDdV5vVi44Q5hAcO8nQp+L2VbywfqvXxGuxzXKoog
6Hm/a+VEB/7VKK8IUhztQQx6V0XuV5Y9hcSzCcUoPSweIM0ufh8ImdWTWychrVXjB4qyMFMbHC+b
rBpykuG0qJrTbakxuu5Ch7XOq32JZgr53/wRxBg0WKM+NiojDK2RMYRHKZ9Nn7II7gZiNWbAfgI+
Mrcpe/E3UtDFRJ//EMsmjPPVDrqinv/FBIYQP6AQR4b3b57zrxgtows/rKb5qOFSG+mO29sDwgw+
REnHBLMVMC1PHK2rv9Tyqhis3MhLjUf52waFylSXvWUlVsvW5xF7QtHp8BEyWuBVcRHe/7lnpGfY
OS+Ohk5N/WIs5nYMnZXD99odg01H3+zF587APuyktvWm6zMV3LopAYCOYjJh32312JRZeqBw+IyP
06kXTqKn8P00+1g1fPbcQhTP52H9OwbIu/DMUSv2PmVRd2lsrKXRehkTTX9W9dHZJrKapGq4HIM2
KkQG1p7ML6110bmolsxKCRwbRECKYUGzK0oePuqpgdSiUkErhfS80cnG0sJOB/XxH+v+qrpqJb+m
2qeFzoTR4EfvurIZuhguq3IlVm87HXZRzzdDnBbasdb3N5KZwiUA4zbeU9qTZrUtIUCerAl3iKKN
ehYrVTaQKV18xTtt7tcchLUb24kLVu80ac4oDFqnmAvvBkhqVXINvZYwZitVvlEpIw6hdGB4eVYa
1pHYognPr7F/bszY2RerRXDA/6a45qh72z7yutctrHObOrFueR3bFfaiQZQLjQhSSoPkhIwoeHwF
C3tG2cCrVfe7xPHiS4c1pNOykBtSAkxSBiNnig4vEMQp8LnkcsMGgTp9ErOXQDU2qgXpVHbpmomY
LShVn8XsFpRRjRVr0SajdBCJNAmqNd8eSDMy6ALz5L98p256zhdpJ2cYL6Xj/DhOyVUiMP0zsVFw
BiDkUm4ve89ROPBIi3YYPljGqFcScdZxpCuIW6NPsKGl0yrVx6OdRrIAMrR3AwpzwQ9NS+HQlQm+
eRU9vkg6x3VbCE2C/hfSL3gPhTKTvYlPwxdiJwduG3uCU4m+1dB9bxNQb8wArG8uBWtqNJkBTF0S
NZDA43W/fUKFeGe7OAhF7vVSquciDmOHZMyIFJMz+rwMjXCFPm1meG7zyk3Ix1uh7ZhO2Jy7jqgE
N1DbVJTFCLL/no93so0SbRhuIOTnDrEyFyciUkDjaWb+SsC7RCWcjzHknPHdIdWVRuezaQ8d0lTS
7ga35L+ClsjFhcqHkXZ1x9IZsPBTpm6a6IBhFXETVN3s0Uhvrhtn/C+oSBN+N2yzr7mm1xdSBAz1
lStsnwD9Ktm+hYd3AhT/gtyZa61pvNFjwAbP/sw4fiX61bPjIyvqzDe88wg6qHiVrOYrHr9+42LE
mCynBa0MDvEwMOI2Wz35JmE5LGwLALsGFUQD1Tv3Wf3roqvjKEQ1L51CglLaeE5GoTUBpibAxUhl
oX3456v1ySd99TT0m3bBlfw4kYE0AeSwOP77ggBAyQv5KEFiocXkdP+R0tOJx+V7KnM5SVzGK7Ku
FVJh8iKp/8tPkoST3pkb4jSYRREBLWnxcf7ultU9sPibPQSsete8djfsb6TvPTsUJCQPHVATxyf4
OUFngi9syTmW2t1RMYX1vKakBLAj9BffDbBISw5r71BrZDY/vljMVr0/nYfG9VWKUr0+yixaqndZ
Jn1I8UJPx+YZLQIvx3OJ0Ph2oqVqD1WDEFi0BqtfVPoI2T4axwqoey/1Slo7mvmoLTWijQAYNI2g
nyNARMWrz/vI+X8Iy3s9MrKLfIVJqb5RI+R6enC0lzfpIxkP+OH/2EsPJ/Evu+jdnGcD2pP0qlwi
juBxAU0O0Xns3yWWv7S0kYPFcyVzVdqef/pDd0zkIPDJsvzRcTmKgYcJvmzkRrDGip5E7P2pml+U
bIo5uLIqLbV3kxGfngRDF/+BsFh8JzuuHUK+XmCb6eRPFkYalANjd9oDO1d5xLRzA3uQu8eCsC6g
eg93Wrx3nc0ky/Zzu5LGa9Pab4eB01IE80ao6AbS5qGay4YUty2RDB6mjLWsR1GC11kkE3XRjrwC
UsmtUtvSMG9+Yl/kdwjvFK5HQU7Chv9WkNydNfcCpSBwi0omH1ByqZBoyWTr0wyQ3SuwL61A/heh
GsgdYRUCRkewTefQGUJSvCWue7G6+7fv0f2Cq/cU+n+18KzPOGPaBJg7xQG9A1MZw12OdJWaBAVw
AX2FSOPp+ZChXlBdjAC9GvgUWwsM63fyGMUb+MYc0DdsxcbjP4anLPeI2AOmpGnvHlpXXcEHngkg
KQ4F9C5r8C6sBE4WBelMvE7PqmME5PsqNIr+J2DoZIR1YbkCK9O5YDVoY7HSkg1cyIMi96M2jZHR
1gR6Vud/GbUZpXi0l3NRiAD/LiGG49otNNUc0NMlyTHy0lID4gEUsasjnrUwrwQr3VXECiseOxWe
aI4VgmaZmJB3zKFqk/8fG/P8c6vH2hwj4xHPglmQkg2IuffiGbYtAVB0oEqI9VsV1cjD16m30/R8
b2fPLvBFKOCTso3bSjbSpLdc+0l/+VjohpKp2dR1eDeY6M6xZB9JOOAOyrs+jygcmyCdLUHdpfMR
MVrZRYsYXc0ahqvmRZi0u4c/CCCVu/98SjiStdvF1mJZo1izxtnKAN9oe3nQ3SmA/Vl3nWgQfmCv
xWQw8BEx9btLpnDsoCA9oP9huYci40qEtL6VIGaTmONd52lz3Hqr1HsQCz62W5NQ7/z20pqFAPGs
cGtYqE96w2BKVVQL8zlI5suNmAbPn+1ueQKNlpyfeb0w4bFCSNxWbGJV5pU3bmcr6Jmvxb0NtKLf
mQ0FpsQcack9QBDPitXxuIgmxwKhTxyy8xz9MuaDcO7u5U1Q/7hKnMC7PsJEHpIG/7luyGeyHJHG
mG0vUqGt60tO9pNV2p6wW4pCMhAf14R3o4SmBVcNARaFw2ZGqyJY5wF2zmrn+sOu8vsbHwm3PUd6
07Ih2YoHuydKPzxt/wXR9+fLDtD+TWdSXbIrc4gUnBT8kZrJBkfLAKPZFlrizH7AAjfGcKQpsfnJ
nbr5xiu/A4+JLjSUY3MuoBHjtxmiimtlA/cjrDv0as75lg4KD0SzNGCNRZtR9PzjsFZY0TDlwXfN
gOJwQMJYBWIMPYiKUb9qjde4C2GdcDyBqGB1G5HOcK/AZfDSxHKqBdhKya4pULZ3+7/XTEu7Ae01
u/VJB+8kLy8x26WIPWS+vG7xJ0sBS1lPtO6uau3QpZThSfqgKxkJlqe1zom3Mo5wPDjMoBTqzj8G
W0Pf7SLn64Qe5WCJmJdVWeczU3HVa+KJM+wYVEYHT6ARsi0h4b9yeKVBJG8ZuhAod5Xc1CrymouL
V1RNFDP7egRXbV9/TPZIaZ1evEBdMUuhN1SLD0ZlbomQNfBVgnwM35UaY1uvMUbm/osSXW6x+Xbm
SAbNKoD14WbqGoacJ0Ae9uXqptzVNJlbaDjD729UaW0DQ/KfWQXUf3o829JB8YrCsEpOzs1RglAE
3YAwf0TXNd6LZqWnjZyEuZxmCt05JdypnfiXkZnvHFDaDSY+MiljPqE2XigpsTPv8mKCpFYqKaEp
i4vvdguTB3IhmMjh7oHK+BLkxnNMqXb/gN9nHzvH22wCNGjf+dIKhH+Sb7E//tgKPblk7siiLmN5
ba+t/ZEovPbkcIHvGPC/esYkKTHf2r8nscqHcs29mUgGiUxvTnsAPP5TS+vZ6ltRge0tJTKeeVLF
Z8FQLq4I6p6e4OCf4Te7wQ3PI/HrRPT1s//XIQerCPjlcqDNHOJ/uqd3+TZmPMoBZmIEhsZyQuAt
Ls3ZiWplSg16si2kGrmnrDfxJbfxyTFgYU2dFBmbOVn1xwxI2at8LIvSsQr1XMMiSpgE0+PrXxhr
nx9Z7vC+9TgMC3FTCa41MV3K0jMvmQFudjsVqWiaradBtFrHOEUZnYMqV0OLcnB/vn787WOGGSzA
Sv15BLtE+N+OetO7qmlK75VDYf53tWnLyLX7vF45UIskJln9c9kRW8OvD3k4lX+h5fVNlFLJTNlU
WoG5Es3qhqAvUVhTzPNgV5AXIXQc8p6meNwq5LC4r67zxdooeDZEK1QMx+pugOGautN6JQlDYvDN
5sXtf/O4gwhU9/9r96fkstneRCsqn/1auWczWwfOp4yJm1BOltRlJhworOIvN8dS8fWgHng9RbAW
Eqhruyrq5mxFQ4+CmQ8BVJfyLy7kWFPNxs9Tq+SxMYWaZqv7bnA2sKA+mM5/rTV8zA3SkezAycwM
8x0z+QLiEKjPU8m9N1alL2Wj46vkn1vgP1oFHoBRk0BA7rN/OqwRllpmy5gavFitcj1Ay69owrDq
eQCQoA0ySGHSC4Pt/TZBd2IlBVz7jh18yWoNqyAeD+X+XIhzWfYdGxvhSIDZdqKaPZ48UafsZ4ep
s+oPzTyYzD6Ag3ef5u7uQXQpIOtNRSds05IvkWGNfDuQ+N4czSRhHLCnMz/c6mISxEs1WERJLdh+
HLDb+Z1y9CXMDKn+Q6KkBSoT6XIsP/rcJRO0Anhk8zuUBpkXUL9GbYiaQtoxKk6ySnIe7KZMyYT0
5xngEVFHD60NEa39f5eGCRn/obVLVWcg+7tv4bf3kK22knrm0bt/OkMdD62Rd9IGRdp34grM4sCA
qVQwPMi8/Fva3vrofJnWJilRLPEe66AP5TwQ6PbRpZSJ+unDj8YKktkPyYW4nyrEECUcuE+IcD8x
yHfXJTj3IjV1BidJ6V96Hyy5JvORRQEOMg+jStRMqMcGKltYeI8V8vGfLCMTk1X7v6lzkoHvUhYi
OvaYDIK5jIr9Fx/QZWVZWVsWyu+c4ddPDwksebPd59jJvjiFKpZk1XuTabJD6dHEzJfVhxNG/H45
wA+wHlsYrd6M+x2twOZkiaay78/u0qb02xoITurxz5/jXTVKB0UD3wVI7uumN6UY73XzVfoICl/B
qqz1sF90sovd2Hcee88TxqZ98k+5KkWa58CABCxjvlRW9nQP7z3J41JxXqRUZGxOH4t/OKUHNdwS
+VanWKNacmT+9EsqzfeUijf2iwkpuBMe+XL8S7o6MS3dZJ3OinLHiN3BAOuVIBHJE6e94+l8/ql/
mGVIEvSuHYjgR0CQOqg/N1GbcIh0pf9l9eYKaaVdVZNqw8+FOM4g1+vqvx4Tq4SOPHmDxehtA93r
8YzoL2jDE+Eq54H0Z6p8Gpa2XdatT6s9Ys2BXTtycFAIfPgFTziWYNWLcnn2tQVL1+Om5ZJKGduT
VG6WsmGFNPYuBOPGTRs3CtgPuEBZHIzsq12fUbVWdGNe/sRKjB9gJH5SqQNBbqm6I+GQul13EP2u
kd57fuZmgbKt8kiEJOM+NCfke+F2GABDWnEeU3nNDCbdfKIgq1SxxlXCYOfZLrfkLjT4cNIHN4w1
xax8S+y+6qiOjHLCyAi0u5WnTlg4FvMQVct3Vwh7ym/1bgb2KuW3gXt4gIzDuJRSB/LHlMkO1k1F
3OvWUfN+09pnuIFTl/ojP0s0DY2mLRRJ0XANGS/+hLtuPPoIFcKblWlw11H9d47yvnenzaK7V7Uy
eMMhILZ1ZwD1WnNZERTiszf0NdHj93kowSW5Fjn7qVa5m7zf0AULgH/Kh7GOT+yipt2BuG/P4rJu
VoenNN/g5PgPugLbK/hsfEeYa9S9GMgCBi3qJ94HF8Sv7PTGo9gujkkneHLZGmxUqBzqoHqQzR5o
XfCdEn7pZOiZuiwCnDenDSluIOkKtZUSVx2pEgkbIrBfFQvGA34mN31NwAgLSr0bgzcsmr7QEBlR
I1vWXN4tSvxXbHWxjzOEESsbZFQt9cyRtePLczfRZ+q9XjkR9+e6O25C6sgShhQoDf912g/VvvIc
F0bLIoAW7HjhzKXBGVtCq3yfB8i0FVRvN5bM03AE12S/MkUPfp36Qx6XHM6oUqck2VVMnWsRgLJ6
0qIClzA4+dAO9P1YQcx3/RTaiNmRCC/FcZEyi0VRnMDSjWqxqCEonMc9X+UFFphaEjK7u6mmfSvz
f85431Uyv3kc8R1flad1T7yg7qysKxIXNWO2/9OhNO/aFkF8iph84D97WuaR1lToOh8L+NDQ0JTg
9YoURDxHrXRbOHpvVW324BB3sCIVCE5gCtT7LIXf5RIJxuf8Ozuol1aH5lmhBTulpO7LQMPlksSo
7QhR465UmFK8F9FPEkELRNJ28YNI6AVVJCzvtJSmtM9TXRWgbJEzqsLIvEOh36RbrDyfQh+bRNfu
nYSJN0J6Uj2mf4suydD6dVJvobYf69MVjIRMZTIdPn47sI3sgYhPwojagtyEmTTmba0AA6fsRz2/
iHfO+lMT5NCOgkZNvR9YlX98Lftvo6x7EZLEmaElPBSvNHD0M/HJfkkznqsARRb539yei/l7FyGM
TKGchQVBqK3w/PBq8nynRH9qQUGnOGwUADu84u6/VQBCPHthRCcAZTAIhHdsN+KQ5+KJQs2zWtNp
vuPzADQe2sLKzLsB5KnnP1Xv5FmE7R7PzhDWq/5XrQXVwVWL+HGLMsm/cQFhM+K/5cFG0Xhbas+C
2Q44wIQm8nXdoqUnG7CxrMy7IL6FMWR2c0pjNyc5U5+0HBNV5ez8kBCB38ZVQAaoVr00rT+FnZKB
I1s6D1BOMk4S72x32g42j+w4yVO4/A4/Vc0lC/d0QyL/9LmxD3d+PQRyd2OxC7DNToJ6Wvia7zpA
kQ2uuv0TeH62oo8RtnCJOU6dS/jdia7btNvMHLNZn88YnwM12hiFhfRLwOrk0z1teHPfWUTiIkpP
tnRkAQAFuVU/I17ZivVUHRzkbHsCql5m8yNNY+fvj8/JraMQddBF1h0rvrO5HZPugOATx2QtNc97
YxY8XNojsvKsqYItwx5U2l4uTj/QTrUG+VQvLtmP1JPwYgFRkQIcTvmlb+AyE2VuLIiAE2dDMfmN
eHBnXRQXiv+a4XbBCXf9tIjOtQKNxN5/Por+UxwT7U0HBRk/Vzb3NXC5gYrKQ0fYkMXM4kU6rpa2
1XeU7tz8w8fdrgSonqoe3gm6ABzr0SjfUBMOshWTJ0Ddw0O1nu/KTIy9hY9bSRSGpM/ts9tLgTvW
8upBd+8KHz7Sb0MlfMTtRmTXr3thOBivpkFQmembnSijrVskl1fEzNYaHoNPUIoFriM3fHJurAvT
CPBbFSUs7WFBhtz30Mv8kJ2e1JYcqwEZhYIcTBHuYjRoKMTZWZi0Aj4CwrEVsZqB6Da3PlPMNfV4
ljgYsmNP0GaxqmSIvwn6PGTowZxRKYWMCMtizJm+z+MCrEx3/1BvUWM7bNADDNGAF3AQ7Vm/vQ0H
yl8PJj+BPs1OorLhlVF/I89Gmup1kSqVerJRROrIZYmIGYitiiBqa2hN9nhUhTEa3USAybSkjnJ/
qnJlHRApKFLF0+Dc3bG8mEgRon+RTpW/dd7tzVtD9IdGlJbWwUac6ovDdagqW/P/nhoZTZAUIFEQ
UFYN4w0NosWb2ExBiVPUlMIcmsh8Q1irEg01xDvAZD7KtvIuOUwXPJzXiqlwC7ALHg4UTNVkcuBO
vk8gfzr204cyToMavhDQa0qiBffP+BfyBYs3UxpZdLebxbdtQCkHQUuQlld64EPpQR8MUxs/m+Ce
oXAYA2Eqx2tAIPLqm1co28NgoUBxPCfYBb7A8blDdHJJXry+sYnGWs2m1bj7T1AQvoxD0T2UNNdT
Hj57/kQXXGLzlHNiaq0xj76xawr1RINM0sElJJ0+sIdq+e6DQHOUUW6ojWFUg5zaEk1wfgScskst
ChZvk8FiaHYnOeEvCTeNEFEHzbo/0p+U9W1IbwBDFh8sA/pIT4R2YDxlmlmyaEYP8dqgwzPeyCXn
G6f7v8VBGmhhnK1cg0QQqTzMKq3U4DzWbyjRv79AKAiSEBweNRoZfjosCxR9eYbO0+q4M+DOUNhO
deuQFEEwayqsm/wJ77NYTr9k+oJJUqemNYtWiaWvqr7diN5upBwH6IEieVtocJkwOoE9Gvy1qtJf
8xZRBlTd3sHfXnHof5m5A79KMPGpyo+XaowGZyiuT97Ndmr/syZxpX6+AOzwWrW2cm6L6sULdiOY
RAV48gf0T3r7CQgZdSXs58/2+Bpa0afQvUXb7udD6ncdT2jevhWIqOFZ1X6EUYyJXAO5xivtIi22
J9/XMth/vhjzu5jHmH6M7dBEWG+g6DzPer6nvWcgXMMkhYqN0zmfLTl7qkccNBY11l50d/WewNzm
2ZIsv5MyqeinNiauiv6TtJD4q7uBQ6K/5XtFAwBAdH8Dkg1sbleDx3AtxGIV1+6soYVasfePSS0Y
ATCeeyWeoRnG9CKnzNPdFJ2Y2JtxYz3wQDS4+vj4ovfCNksfpWc+hMFLdl6bBcn39BELTWUYU4Q+
RzIZ4AUGeJ+Ijs/2164yqNnuZAFKa/FZz0IUPLLTktOZbJRHYiIDNWcaLvlFQ5/A/LBdqI7b1vYt
cPTc22pwD00VL9jzGT5L3F8XTmIAwY29reOyRgDpT772PMCWLRCGsKvtlqHKFZFre2Nkis3QnBjZ
s36mD/S64qOuxRHlcOBZjR8XeBPNG/e8mq7fxoHXqLTkFHsfkOuMDkvA6yM5vX49PuAk5SF+6tqh
psg0YnpidtsZM9M3dKrgEusUWuWb3SwEVDskcio6ROsMunPPTSvXqO60ttjAyeG8wG0+09su3Y0e
lxjgMI03R+za2nPKv+7eXPsfYOExUKdQNagvhq3A4AC2CkGxzw21sPxyDeBbtwrQuyV61dgf7t1O
OtqYEoNZA4eZYFsGPbBDeyhBCuzkKP5UFt9Gt6CW7GndNhw4LJaNH0UXZ8gO540dQ9uVAufSuJEr
hr+zxOTRk5ns/CRbouubwXakWXn0g7HeaAohgoLMUcfOHuefkPcu3pNCQqEY3KBixctVFa0Hbzkh
kQcrKIQS2iEnNJNJPr8OoRTAFTYclS5hfCGRqE6fZmd7Vv2/jSXdkBwd4Eq4KYP9uZKM8dHxN64J
mF1SjjjRousCTs+2O8TpGp0qgCeHB8NjjShAuvoDxnFHGFgJ9eNHhiUHWAvySL/1mFJx3Jea0KX7
gheskVHqy71DvgMtk12fEAlVfRya3nJkvEQmF8qotR/qULVooLitoUcLbnTPwXL0Z2DhmWoCAtNI
5UstSkkutM1Lw3Qx/nhHGJwED6UezreqnDMzUFzM0FbePIyi8Jw89FdM5W9zlPaykkmPZb5lTTO5
z83c8gYN2m+C41Sl0hRcrzWHU4nvwOOgauQNGgQqL0cKfLLbOa+By2Uo7cZp6y19fwx4ZuFoekV+
QIG2NofheuRtWWudUhWZB2vwB6trlAfYV2ypTeEG8WiGJFHgsldCbd7sQb3L0Gw3q9fZ1dAMkxHW
FCVi9+YfbTUdfEltAVxFIAV4Kv6Mjpmg32wvdsMI9tW01j6YCbfdhxii+zTnzuT7arDp7RoUC0NE
O3zwNr4Zw4jFlpwD75Y8pz++/GnJAwHYmQdxTfYZ5J5aMlcRphCW1TmqDcDL6olCzAAMCTpl23Oa
KlbWRB2ma5nqKTJ/g4X53fCFh1IlC8W/By1K8OqO6njpJD7gs9X4KmVlqFHJejBrSmQJOzK3uP8x
59KL8yy4cTvYODY5WFX3z1aWDqXi7T2WCnynZfGEVLC/WmIv5XP2S2wEDlcbPpHeD6ebFjZaauyN
jfkba1LCizD8YJfHfDjeD4MFAqCEAZxBKXX27OZa5ZAzdx24rU7yghQ9LTh/uIrGHj/Q8y4kG70y
pALas0E8qe+I6g3cMBd7lw2eIPhzAVHqPKNX9iSU/pjv1EdaAIVKt5OYklA7zaEc7tsgiP1EvHZH
R4An4V2TOrI4x9ka3X1MelaIwp93enUm9HXIZmhenSU/3mlGdr/rpqCknJSbpoO5Pv7bPcyhhxRF
9FxZmcc1/9SkpEJvV7ZhVCdhUcV5uTt6fTv3Q3E4SDGF+CXYzvcg1AjxeRaNXmCHCWyzjbDe7uq4
V1sr8i5RNhGOSWjVAdPxLtwCIHMpO2qukhDVtGZzfy99HnqVFfTy6rvP1WTi2c1MpjAi8aIWwh9p
u/9Vk4fpBjikdnYCd1JhPsGV8xq5a3ezTmcs3lsCyRs/Ln86Yp7zlhYqY68RqoanZcr/2/KYrEOA
DgtR/4dyvyzigRoktgob4re5C3baaAiMEyAKBWcYj59aZG34ySikQG9HvykFdgsSUYYxg8O4hPa1
LQbJj3bHnzRAdDSA3ze4nbyZE6IuTYYh7qH4jVT/JPWbP+JWSn9Q19K2u/cVzp99oROYTPnyketh
R0kT+te1oIuN1PkBoDig6UtZuHBqJzaj/bdluja3Y6qOOT77TsJdIsPaE7EtyBRACNisB0bsYycO
M6Lz5Mo3ECrM16SAunVMNt43SyzSDwOyeFBVq6xPhFxLQMOCHi6iOQSxuejx0y3I+nMveA7XaFD9
dkmhhA0o/hDzaA2AgtUCbFbOATpmHhWWO4g4OFOkdt/R23AbYDAzwOUzucQTQ85M5ScK7nwGe6G1
6HBtfsAQ3cLvyFl+2JnvcqteYXNpeGKpj8V9YnKrUfboKh961+LOywJEu6UbQoTbIVFyJQB6LNIV
UfXI7Sci7oBA9cu6y1mW61o794oO4dH2t8tMq5zCI6riIzOX1Tk5raPY+MxUwTPaw/xi4qi729yB
Hea2xYBrh8Y0qfh2gBbQ2n3HC1rZ+vdkkfywYYGVii4uTDARxY+iFWv4pmNCJR6v53f31MnqDf6Q
tR8H/jk67HqSFzRKhjxFjsQBDQDeLvv7WO438m33x0Pm2ZPEGfcn2CgyeZkcsSXxacOm8Repeeyc
ZlV/ZaM8L+nuFCupk6+AxNBTxdwCWqsW/bB0LPtvCFys7lEhhiX89YZPSJ4LoLMvNQZw/HdP6Txd
YO30/x8kDcr9eZDgkQWU0BwWhGW9NJFSXtKj+VDVfI7oPoXMJQClphYu1tcOxFrKywO3I3TKTPNO
vkhhmgB4A7wzWcxcUFGwXTcDtRzd+14Lc6qf5Fe7a70dosoeS/hw6HHp3d2LmvBXRT4ywpZajzKy
VpKcOxWmCxqbqLwwyMRLzv/JsjV7YP9fsvjZo6fUat7m3khFUlUVLAGVajYCStLuglbCKS0F7MOe
uTML0IKRCVrdDr8wcxEEjKPoVE4x565OZ7jUx5skG0KM26cSaEERZrRtDrw63CfF9PgsrDriscbI
RFtw20FzSCXvEzYaPeMxFRiuCshsvwamXzr7rDUp5ftgcwo+jJdd7m0+yq+rWbfrmG5G2kyBIZYp
OOTb+CTxxZVP4iFmS7d1NfPYQkZnqv5ssah2Bgi4oLdL1U4beFVrOwjVV3MdSHiqVaxC/u8wpWzs
McZLJX9z+NZ2GfKoth0n9QrVTIPuTrXrePXLtVDP+SLl3Uj1vR0ApTda59E012n/K4YRoM+Iph4+
U2jEocUKi7MiG40S1homv2BKP813TzhdeI8du7F1nTr2CdFPiPkp4aT4rdoXetr3VdT2G8jThy1e
+9R+eeO8kdJyJjFVaKR22hXlxslskjpNoqusEojrZDw7ikyPWQiEj5VzXMwSagHMwRv1brPPVSb2
zHVvSpW+yMSMnPGbFInaJMPX1CS8xBlqda0qyzWTtJvdVyoxbs8SXzUsFsFoTp255B9mqFQcbvdy
4ueqATkawLehvZA1xK5T+mtEpvV68MBqGR3ng0hkHXLHQa3MvDeCym42KtJN5woiehl19Wd6Q3Ix
j50JkXZv4Zf5ZAtYJbrZ5ZS5CYHBspZibN0pa+r4fR/vYxTaMqG+yZzRbRq0/MFrhh/wXpCgqITk
GcGGIb84Ebo/Redk4zhr7n9crZfG8TgIXOmJY5DjUtcognEYuPhCwcNA5vBDiumsamJqPIzqH2Bk
N3htmvXqCqxrF6+G6GDWbh3dkPse9z0Bl6yZmDguJfu4xRu/Q6KbK7pMGnAyRJwMt9tAZyzn+2JO
7Q0eKgO4zSN+6clfC3XwMIY8NNtAp/cjOqX0juWJMkb/gFiq3UNvtC3sV2RS0+Kc3a4sCkul/Ffm
odridEgklWt9+JRN+Hn6+dOZTfP/sZAX7oeETiBCnvoTDQDYsRi4Zyr4ecrlWDHKZR5VckCTgwHx
aH14zIN2yIJIKAjUjCE+RKb9Lz25ikeuFJpU7wfsWoe5Fzy/rvCBp8pmdZS8IKR81uEN6Q++CsHi
LDznVLRMY2IitsdyJNoftOgCkRwMU3vz9NK0ZzYGHxxbQO5lFyTc9f024M7fFwiBKOWqdBfyRu6o
3arO2pUUTPGg8WMzOISJstWDypbWYwopH0dAbOcoi6x/u+HuxhYpiInWwNzOqDmMBNT14Th2kNHl
0qjtmlqouwkFT0Tr+Bth8hmmk/0GIidTOpcX2vjyspS5F/dXoXPZHVFxgQDazmVWkw2CrlpU37eA
kAnK1MVXd5dwJeddtFdi1+/a9C8ZEy1tniTDS8APNUbAOZDFufb4iur0j7UgPvs1tPY8azEGoVT+
7LxYLZBQNsCn3iCY0l5EkPbNe8YMPyKp+oWFYHJbAVLsMu83Bg0Hhlt+K/rc8TmOhOfSdmx8mftU
Qhx4wQfMAB/YYT66joPk4mIYcD0xtxy6py0rMdWzDWBCpbewXf/9EmBXbnfZLDci2Yl5fJhtWBUl
6JVAP082ysHpQ++LHP9C4g8HZe4+d1/baZ+ItQBjXlg+WZPJqUzt5jjuhUwQJq+MbNoU+bTRmkBY
HL/MSjAMeVLs5bRwM7wZVpmO56Iyq2kZex7W25mKNVZXnlv2zLWReq8LgOq6+jj4DHFnRKHbHxxX
O2fBld+RzUWoTNLbdgQI1p4m9V+PmJhsQsOIWgECY8nZBcDY+j+o+RU7KIAXMIYT1DVMYrxjr7Ev
xyjlKnmvV/wrg6doPlg7uUhhvkuBP1AmxMeA9wwKtt9raNnRztBVM7tj1HYY3kkCavz1h8Tc+I2P
JGDEiV+jFAKogzADKmXg1fxRO8fZnU85VDmzQnuQxmHMxFxpBD9R44T7g98GtJBjTmLTg6IDjb5w
8ZM0Du3vqqi5mi1A6xUG37I5eXtfaSCxyvL6nx3RIvhbfWtmOUe+XqcGnGeksomGfjm5GKWEF4TG
WS3zgbjpS/0dF1ApSRmjq9KH6WRUWW3WId5Kp2WaZaXIy4t5DKW+uPHXrmXrjV/JZUXs5efjAYKo
L+dBZxxZWJpPC9r/oiZhxyqDVFE5iZaBTKtw05U65FlzPb8TizAQUIU8wcFr1G1K+cURBRasatYK
PcXb85pexPR42g8+SdVj4fBjWIFBoomSFyr0TEYgsYbhX0ZcVwE//h9t9mt0UmgG5d2j2IfJv2/h
yi1xZRlA4zdxt4znb7XaPnFkkWlzHlP+zkRyeMo3FufU4WVinLGE3n0M9QJBcs51ICPxxAuTvycc
yzbvySjRxcLVURkEChua2t998lodtdglPU/7371Uw7VqfNpHeqqZJ0MN6tsbisBA2X0zPdCB+e81
zxyWe/rTvg7jM0uOizUOWMO4QKQr2aF9gYbSuKlBiiYuWT/K5g+mAs3Ps/2fU0cP3t1cP0GRzqPd
Kr8u5jwhNNHxb2ainL6NTLTmM+o9wr8SziBCvVYgVlJAz/bXuc7icwS6nXH+yLwHVtIzhwsq1Mz6
fxU6y9npE0SzE4uT98UskyQ5cyVDFU7GQat/b/JnHE8PPiQBpRlQsPaOvCdho8reCY3sWTnS2hSJ
dhzVk+I4TuN1H0b26BrhXNqO8Nz3WuzzMVutMAWowHe/nqzu5PR68JLpVFJc0T67wUFrBcMRwOKa
4nH5cIwPuj4piqQwwsJ1GjvMpS5GWqysvd0eri+ySMO9rVdV12o6f7UmrVRjpP1AOI4ATpb3ya8E
5LXTu8pRNU2n315zDE8t9Fc6JlEovSzLo9mchAVzkCnUF3JC86XovgHyfBzEqbBixprq6dFl5uZL
BFrcRJ/W96Lw3u9UCfCQM54m9ZSM7Bl/Ib7QAizZLjp+iCIwxVENLtcMs/nvB4xMrp4z8N6bhn7x
z715vLLfsuSlmgyAYsZBW+aLXPVHLc854TudKiZ8LdoL8CVRF7AuDSevAnEWSaLmGGyj26KK0T79
GP1OtAS3u1/25Oo6nUtpokcHuywvTtvwuORPNs5J4dYNfX6L9p9S7giuDqm52Lf+paIH20sT6cj2
lV7Ya2X8sbzfuEHMjr1+lsg3VJ2k/+QyfuRDMJP+UBAFMqiLaml+xypk72IcBvEfiTmzT9nilyES
yvhIbay7RMkOZ+/LJu0sOjSS/beVzf2DssN5/owqWK845XJzi5/G84iiYAaM2f4p0naSdpGUjvdg
/mTTgv7XCLrjrDs+vfibiZoCPD9BGRRyCz7VWycOnSpbuhLUCiJEEgKzx/lNarTbZErkY3AMfNCk
XxT62di8G0MmP7rmS4uYxqKRAITm8RZbF/QFm08V8fg3ODjNnGF+8VZowecNSgegYZIMywpfLzHO
MD6mgDCC9TvRpELRzE+tDoqLRbkGB6SyqXZvxOhCHhsnUQgQe1F9HvfkkO27hVc8Cxfq2HzwxgHa
JlMMKUKJI9HkYmmVcmyLdZEtIGYmCEtqLPnwSNitMgL4sM7qgpF4VawXp753dYW5kIHKYnoEoTRW
R1hYnGH9jXV3RhrSXuou45klYAiT70WF6bHC/Br/lD6Fnxi/TrqxhkWiqz5xNDXwXqWlhQ1O9qKa
RDSsARMlxHvPk9L3bEFMvDX0IKyhpUsrP8iCbAhbLjpP+x7bWrpSlglRS0WPbkcAurQSmFgW55jq
4O6YX15TQI7r+tk6LZ6LjuT20eaVt8N4AMkd01hruT4pscO/kMX8G1BNujIs6lMyhuSVPROQLhoz
ia2TMiqZFYdC4ayx/KRMWzjvOkeA1fY/5kGUFPgooNFPAg8RqTOWNY4D6cpvBHLpyaGz+0BYz1bV
2N12u1RWAy4kMuVKUcv9P/IsifRbp52hazhBBb3+ikKnrRw2qFP9gOVMp6FoKwJeggbsvK21RiDf
MabOHxbeZBL72acv2Yzo9g58/XWssuKBIb2uFHImEGWPNU++Ll/3HmRHUkkSQLUaR+DnX/D4FsV1
HnzAJjsjy50nUaRCv3Z+R01zBj8/8btQlru/Oh/jhAJrDUbh3JEn5kZzJMYYR3d+j3mUO5t4uI9j
3FLIPFJmO95cdLfgNlU8mCxmjukVNNGM4fXOTFXFbx4T0Bmhm0/84LizWSFpTEpay901p87GwPqP
DjCzLO2eox9rZjJy1+7tj5CUU2pa7RT54Pa4BF6TAh/ttJksxl7cctNunUd1GnPTEOTJo22dTLe5
LH90lLeUDrhyWvaLMoqY54sJ1sbkhW9rjDMG7Z8yO8fcKcoWhHAT/UIWqXj1bKDJB8lDhODUWSFS
oUPie1vzOL+RUXEoq4Te69HnOR5t6z77uvXwRYwv+J5tAxfJ/S7poyglv3H+bYozXF0N4uMzJm87
I1n4l2tKGuiYIySrzpOK1BWK8nEOdDUoq/J3yzTQ1L+UgdoebG1qofBrIjWTpqr2M2zRdjtmK1+/
yz0gELdsG330kCIYdRNfrY6vjwevD1MAcIFTvFuyb6HgwB2OtEM8zor3guSSXio4GYx2GFr91W3F
S429vJ4M7M0rR6sxoU21USpZSVGzqk+iIvhvo2w7uFqKruXeLTq7gMtV2z3YFx83BDtFzQDgmPAN
/Yu7MkZBg78lqbqn0RCzM9p9SimiaY9coBrjmisyY2lCOf/bW1cZp7Am2DwhXFG5WaZL1w8u+5vV
RRy2r2aqUuGL7HY6vSgNZAiYxbCFYV9BUBgaOB2sgWeHtoy5s6dGZS81tRiBcbyb1LN2BW8oSRSQ
wFgPgXnWK4tAKO7ajNVW7FEQLmN7Dhk1l1fGhGkIo9MVFpv8GVdbd45JmsYCszIFd0ysiZD6UkBb
uKAfXzQjoIw6MpN7fbjEePm0RPxrHoxQZy+kPclddijYQiFqkNeeI+xRyPXr6osdx0a+LvKDeHAK
uKzHnRleDJNhMwdic6wl0q4FJd+aflFYvrUVDGetE7zMz04B3f3zqzwFGoMCCXNHghVGmFydfjjn
+lGd2w5GnIEOhjvdCvNh7Is5M9X+UVaMH1wWR2Qk3uuZWZ90UlgmsTZmH9p7wJs7tq7K4OXIo0MF
nDr5Va3D5yzCVr1j2DIGVMosHRismhvVmTPnoAhhhZkjwnkuLFQ+H/+EcT5NkA331UHWkJnI9AeW
wEYy9cNgLrKVHLPFfxeSJuMlqa3CNpBTMlocy8az6Vkn+hv1jO3JUvqgWnGW/XW2fd/GjMZ2VMK0
l+qWIrWM4FY9Cxbq/GpvnnPI/wQi3FaioHbKUTHtAhiZ1HvltMgl3lshAg8EaHNEyJU/KkUb+k7y
C1giuHacnHu8y1H6NF2fFDceBdASmlAssTXEZKBcg03zC0Qtizc+bV4xW7YhHe2Dt18paQ/uFhOK
Jp5QKlxbxeWcIJeNmdVJqw9bAdTPph/zSjuDtXYWYcN1Ww75VtHqfrftoHLHbjYsJ4wuhN2oZQQW
TKembWpk6rPCBdbrl7AMwTUR2071IJhxYa8kusyyilHYQw7BLrbKVqyYWnJXr8oVTZSOH775XLDq
VnVR3C+QGdFopKQr/YvQyClBOSSW9bV7V+mc98HJfNB0Pcq608ukrSir8yshtoYTJHqXWJTf/xON
BTacIcF8O6sjNDPrDmQhv5zUfCM75EOA7zykGJNQxT0J1VU7LoSHpXJnekf5+Exli+pZ0J06z1ze
gq4LWDfZyyO6FXS1c83UBnBN0sUMrzndxFirKaN8fYrstOxYz1B4pHFQmYoVejWqaeTLARX79isD
shb//z/TkRW8YdQaemagNrNEN+nyI15OtKZ2zieN4I3RjIqJ2+Km8Is+eNcWeeOJhpENt08l3242
2fts7QjYnRTkE2hPNsvdS9BcobCO31x6ZdyXzPB4qrheSDLThVVbdc6puEHq1ZMQ0YvBSpOoBgxc
3QeAgxQZ5clKZ3dn2riwbW8D8mD9pAXRpZ9C16AaCtqnZqQk241UB0Rfzz0sooD+fa0RWo1ibxeO
Wg54eOmAObvR78jInaNEgYodLnutzDggFFMiPkNgedB3P8CqQCfAUE+w4dpK9A7npZamkjj3KSGR
I37spYhMGVB2LQACsFYaRqxQaXGth/bWPdccrh6OcTKYXpiLGqajw6M5Khwq7U+S/fKwhgnsHwIH
5FDGvmU84h8zcnWP1e+DG0KU/iaj3pU7P44AeFQyNaatmBNpwK0ZujFIhjHr+cpl3SuvsB7KUSsS
qCkH+93S01wOHBzBAi6akk4v9sQS238DwJ+bAY0//7JQ//eSx3mARCdrCwTidPQzBfImhLW6Z5kx
Q90ClofoJyoiiqN0zz6bwxy5TPKT+RF4tyY0VW0IdOYY8Kd1VPX7Jci4F2Y814liNNjWrY3k/u1+
2kZyGKGHNK0Zojs/4UXXAzTU5AIo/Kfo4p6b9vXjjfdABlk3L2nlSk7B+Q2M6/Xz+eVgF6V9Yu/P
HLtwtSRQ8uFlwdQCbw+kIcW/iNc2qIQSXUZKOGsjp08503PspBa3nDO3X2cvYYgvXUW1AjCmEyvu
X6aDGYGlrVk6w/iSjVJR1XLRYpIsQnMoM3xlpq5XLLIxAsBLzBXRf2GEiMlGny14u39EHz82vvYK
1C6L36iF0+AdSLFNv5+x6cHkRvk/BOuUNV+CBqQtW5qKezluNUcmadat9N0wNsZxI/IYL1iQ91vf
W8ExWVK5js8JOslGyTFshY8ID1uFBrks5a4ArY92n7YHX2Alt5nSiNdVoktyAwWPcVZPTNhuh/N2
NW9pVe21R7dDaS/qwZSyq0GqxySfj3CP2aMHH3eHzcCDDiO+OrYLXas/AMQjL5hJFbd9JPBmr3X1
o1vgGyynqQCCL512jhfkXYdRSzF2sigqll4WDZzbzSyUckyONEB70qikBF/6CubCRv6Df8ZtzxV4
6ieVXOPfSx1DoR9gpyjDgzlx3VAoGCcEvL5l3l1Px7BIn/HTzxdQIEM7ZcfVSOsYLIydt7x2E3SJ
uJyjAKTyTrwbCFLfugnLNBoGsBjQq9HiJiL0QjMFAfhFBk8YDF07xIar78CVcLZ5GUkPqpn3ZYP4
JT7XblExd3x2P6hrfiViY9MCDq6qD5begEYLg/dbSRiq8NNumuGLMUfEgl6hkNlJkv+G1duXmHMz
Pw7MVDwk/TYsmV1JnCbtOQdwMVoNIGT7+exEsgohfqNQCnko201ZPTREvyB2/ywawmV0XV50o0wa
AQWFf1/AqgqkCEmCgq13UCCURjdaM+hu79B6imiaP8nKeAyTZNZ4gANY8lN5VTILqpq/ZnTccb27
LT39RQxbfCuVumbo+oYaigj3IHyGw9BWJSYuFzTj7dxrAqUJVW7QzJ+X4bFVCUT0Oq9O7eGt59n0
BIN0J89Cw324lwFDZ5MEQDrJ1vRli9C1mtWn1IY7E1VHibdPara24wkjDaVa5Fh09A8au5f4mgBj
9ZrrX73PrUrmbJINjJxNvSlrZhgPUN4fsd5uvcwUo2nsTjI91LZ37stKw9OTmFu5VlRPv1R24t7D
Rq0Oh8g0mLiBoZNy0/Bh/Co1kmQ/GCVXcavwUpqdv/zmWYov3bXYWEmZQ1cFU2lmXsmYPRRLEI76
V7G4PJx36/ohD4i+DVYieQ0g/pHrmcGTc834d80CfAQRibkou8yZnmhtls61x3mQoMZsMNN5dQCu
kItNQP2jgT2X7UzZ2p7hunPXXTRvxn82Idx9baItXSOXFYZWjDx6spJm5nNNd0Yt6HqFNuFCghiz
swGqUtF7J7vrzZmoR6lRJhENi7OKJGbMFW/q7QcGBD/LQKpEf3mrqjgrauZShVcqONlLcqk2EgoS
23pTPDSJiUDAe6lVhtcuoL/vn8peOW67js/QSoX2H/6vY4GlfCuK0E/cFEb/XkLLwhPzsJBBVGoT
zvnl0WW9wytvStX0D0V/JLHsVdVVUWJrx5GoVY3FyRGziTeivpKN2gP2P09V2keiGzZy4YSoCLEC
j492n52CvcJztiy62OuctN5bGvQVRFeNvBwLowU3tB9+5s4/vhtx1G+MWqXtu/T8ew0DYJ8WqJft
QQz/m4V8sQ2y/m9DpdQ2Y7I8qZQTnIOLHA0U7rwD2cIeHO1pRYrsXvrQl32dENPJ0jEXDo/8Dqln
xW995knA9IjPeBEfrM1AxmEAStKrAP28XeESaMH1oQx7Efo59yxIhdztFcrmbgRDv41bh6eG3/37
qAt6gt46B14vhbDihdlAsv+nbgJFUrE6Y8Q5UaYBwQeTHiXjeFZ9/tE5YZAe8ReNCWcPAJztzUXr
BZBbrmSANbv1YY+RDmdIC+tbkP3YL0m61L/HvzHF8rrT+ogG6hvwNWQS6rVyB4w564hVWSwwNxS2
ykdmNWoTDAuabjDnox7vTvM+UVz5xtfpMy1jf5h5iHzmijHERhm5PyNob1XsZYnwmiAzbPPJVIr6
GWUtYTTYaSKu4KLcuQYfEpiOmybrfq/JD8RYNNnI58CzjcM0ySM3REN/IaeP7i7qmeDhV3hLpeBS
ldSmClPt3bWOH7ZjkW2dEvtP7/3Ha0J+Wji7FTuEOuO4e32mS2RU5Zq1/if4ZHio/xAIu0iiF4oo
hPEo0fprgE7kyISX0KxdErQlTbK/YBVJnR2MuyDI6xh8qc8wDnjmVzPrZA79s1hwsKbC+wF4BvUq
xUx9WUz5PmdbqmbuHZNX1uL8El00jydatoRJh1FjTAUqOLKOluh3iyrzquwL1wm29IoJaGIBOD1N
DiANe0Q9pmwhVdmGOKdkAAcoihAZKlY6j8ya97VKI6aSBLwCu/R+r9i19IMAUi7N2SGiNbxaiyUn
gw9mclIoLId56Qa8zj8a+Ju6oA+xtMPc4qumTz3xHNltlxjlSxOq6hQ++KkDNeeYis6CxAF61r8F
N0AeT8VX1/7Dpw/zyX51OdqSwFVj+zlyOMeLPggL0ykTVSh6xjBE96K1S4hR5Fjl7lqHmNzTxDzW
oUhD/fH/XzvLz1B4Igc+KDQhK7VKEdMRiUZ1+w9iMQ2rny5zD/47Y2awxmXgGo73rPLpVUVvMagZ
UMXodQkmuw8DGcbQMpHImKw0DWp2388+BaOgOSIyZ3tsW7XBfIIXEp29pQb8IurvZObEa7CSf/Zz
xEuNEoNkENvQips/xrrMz9H0guiGf+xQXQkA+C9gAXuuX6QeyDC8YcLz3aLia86rv8xlLpptzGI0
EuV3qQi7jjbfE8QYpiy/4+Iy0TERW/3GLuXiapMWHML/cqIRQ3mgKFlHt+TvF7ImGEK2WGcprS1a
Qyx/cJOKI/IPWrnpRb1WqBxyr5f11aw2hRyIsLYJkkYUgooEnPdLx3Luad0sDCF8YC7/6xSsha6u
wapuX1tdQgRpm7Ds3Gk0/ZLI0gCujQ+22GFz8WXtSsnrq2olQ4cA73jugwDQOxFaJvojh4JJiqqx
EbtW4YHuHlyeP52rro9HXfmmYR5Lew6yr1/4aDfapNGA8lwhz9SXvECKS+K9SfghLJTfYqUGIVou
babBsfZHO5DGX71Q+3EjhZnMY1qqswZ7Vvhz0UQ3cKOwhw2XXcatqWpvZWB17UfnEZA08gPCcyAt
XaJHLbKfClCVxyCA3aCR/HVkks7ZIe5cZ3Lc2b11ndVGC/R2clFBEzVqnqiMdrPkz6sTsvpB2L4l
9TjA6Y+3H+y3qe86eSv9WeCqbH7MZjySVVKhUAM9o+WV+7PAzPDunK+FTVdDxeoADtSgPrgxVcbs
KxzZAO0troeX+c6Mh0A/pojbNYN3ezxv+ON7HYHJr8GqXuSKEiaepbIouG6a2lQfV60eKD34ZnVq
rgr5maajM04zvTAGWnwXmSSJRw92oHr0WaW/6KlYTGSvXqUX38+zVsiT4FuB8ayNweq60Oa5Muw9
ti5sd8GtVVrlztGvyB86B8+5TOVJ/6sj+cMb4QNsWzVJl6R9Cl/CVtsyZ4H5ifuZkDRZ0lAO3NNM
QVdmTGU8ikmH6zXaYvUl065QBrUEqFmyPWhPiet+JYizYxLeMiq4LDexT4RhfJaWXUb8LYZodAxd
UV1G0FTgQlcILbi3BSg4EzIrR6thmV9vt8gdeaGGxOd7QkX4iqFkdd9+oPgL4m/STGxBQFnCkAwR
D+xs0fCxhhbhmdjDVs8BPqGsOmfrqgykWhOQDuRPA1gItG9wkoeFGJ2ArRtRGHd75Zkxd9PBMt7H
ZJG36TifEyDt45pGaPLw8GF09seCTMM6+sTYFIh4yGhH+AdP4WIrdMsaZ06RD+2IK7tKnV5wb+05
IkWKfqkSTY/lHePuxTKWp738iEydkqgtYaEAam1d1CmYKrnrAjqBbGI9GVuxjQvA9p8RXIXXLfXN
8xwkVWuy5f73mPxjEineWc5Rog0y7gA0YtEFvo/dCoYdkkcy008wPx0cbiuzD6E7UhQxKYiNprPI
Cm/47I9wrQPbY2G1cSfRvIXPyFFF1sY0kCYxu2raljkjSAn0p8ynrWd1RyeGjYhMjOBtxITkuigB
bQGjWFjAkqSJXjFr4ciRIq5NqxwpGRs0IBavO3aCv2gRZnUwj65dIKjEzdkvB29eamlnIhEOCtmt
O+8s6b/LlenL+J6KEhs//ZSlblsTu7f7/kFUXHaMWXG08vzvPuS0mGfh0ZGw6TsVquAJNinCTij5
v1eK8BlyeDccYds75XDm0KQMWHI9z47lIMQRF1f++GhM2IWMdKuA5gf95E5l538t1f1eNbvR80Ai
Jyou5ScbTW8+Nrre32Vq0i9qt7Onduz9bmrvSKKsvcYTJbrWuB1f1uu1ExqDQ6XpxObn4BaYP7qV
VVErAlfq5BFQBl9nNB2+o/HEwoOIa5VQUG9pALSGuTJLQRhUWrq36ZSH0fIyfKD93R7szhK7DK9c
yDFK0jxhi2/8eFamvv6etwatTOotaZ5hlkUAxL2YhQdzSSggul0Js07WwYBAo/DIzRJEk5uOuT8Q
ksdCyjVHGgkJTlTD0RVVSKsxopAocz7WYvLoyhGwTbmQsFJa4IiKHCt2mtW+YQuQxWBV0syqIiGb
j91Sjj5PL2eLDbMyQs71ZF/KZrW3dmITobw8KEcKmZBIYPig76/9z5qqLkgkEICnvLcERbNaLxzX
tbDKIU5w1sS2FM1Ik79KumI5w6kxpOw48q8dXHSypknuTKqpUGCuw2BeLbZiO0d/Yh6yj2DSNfpV
yjAkelXjPQT7wbgFXI/yNOjma7GL4+n0oiBsVxmFMda5hPYZqx6UvhQUFUnoH1g4KAas25/g6E8R
tzOAn//bwMoaADJc9U60KQPypueDs6HWMEumh/Jnh1JSCc2kC+0D4rzGYLYmE0sq6G6Dfn4Kg3Xz
mrn88TRn4Q96CsRwXZd/x424+AJzoNOyZ/46AQ8oF7mpFhYhRnXEcEcbQldJvsGQiJKNz7HSRpRL
WsLrExmAHxBj8FFBcB4SMYSr+9FyrUikybPt0mjfSVIcp4Xy6A61sdspIuDAvRmGiDYUCbYiuAgD
lVRGGLm7wuUhrB4CZ+VzvuIHai7Pikst49aJhQ9ocCZ0L3Fw6UBXF6PsMs40sV4iefQTFbkOMi9m
fPpyILJGaYsTY0Iwyb92vnid/3BgOWopqypvAiGnIcElyl+dABNs/wS/OIjXNWr6SP1r1TEayR1Z
OuMd3Hn+5a0iMP+KMgn3VosEyMN3pp/lWznsL8KRg7egaQzUcIY2r5PngA/4pGBDG9TdvxFPhUVo
aX5aUTqoW5I/JHX/uB4p/g/VlBP7F4MuU1u0cHHRUL0lSAtPvWGvLGGZw5IH06cKFBz9IoABSKaA
oqTxE1qukNiePu1qDdS4WOQHPyYhvw2bw52jnliOS0EUZ3PsY+6wIYFs12PnLP8LM2SWPOt5kINC
7DWK5PWgOLVqyu+MIAjdTN0tB799iL7IRmNt+teQ9Qm5q4NxqlK83IW1yvIIwZjJ0ikWgz7NS69W
mfGZXSRsmX5drm/prl9WoRskf1LPfukraIRivTcYqU2SpbZiv41XCxkBb5AcbfvFP+SWompb5QzA
ZzCcyZEMQrxWxi9aa0mqIBvddVjyULXwkjHja0dhB8k7ulnAy/gLe42f94iFATo5SjBPvWBEiyPl
knYSUKZUV7THofgM215BKnt+xuu/nXLjxxd2rk7Gxp+euMgEcrqDPR19IuqZkLqIEDlHAIWXg/wv
cRzV6asuQsk29zy2Az0Cs1fNDmhSucnJ265Fkk1pkaUuc/ObIreBSpJr1CGL35AoxIZwHAeBU3pM
1JOUAGRHYlWCRC0vVSuSqHDRcAaBbgaiK/7xLZGkT0rrqVVXTivlhWCFR7InE3m0WWfBvAeJtyFe
dW0irAkkIOqunyRCRidZewoLegK5vQyTr+V89O/K/MEcJ17ficETLvUVJ/0QbiJU7IpeB0vtUtTm
MOoI+okvhYMde6s9dhw/9W5loNqvP/5P3l4ZPO6njUlf2igEgigskTm68TeERuezuedjdsr9bUXc
AcUmihFsccJZdeBTyENRQ989FolQ/6jCJR6bqigWles1RX6GL2SUlNqqJWkCaHuQwEM7/nUAHDg/
EuhvHkZjDWpzt6LeOQpkr07eVhVhh7BycwVkF24MCKW7Q9ooYuSnq0IosvxVFoWbUQslPfmCjsNt
AvKNgNdqOWKbvEzRXqw77nw2wWsz+/RoYIN4xxm0vWqoRlH5Nw946cB6QF552/xh17/3G0tYjTVZ
D5GRXwEzLwZoBih20A2xz5cYM/CHeoM+KRLzcA6TW6Kod1RXSK22PRzBV4Mxjs9oGSQPtuwj4i28
q00x5OlQrU7y8UHNHG2XVUVvpsg+7YdayYkQ/60KkEwdOGElKe52XMgfqEvhDfZG0AEsuFOEWW5S
LkU74Xw4UZqckFE49Ujhbv24KUTFugCGdsnH76Z6+q162VwehtLuZIjwBYRy26ZjTZp9pbFP2R3n
dt3Gq7970elfprJqW3Wq5EOFTMyKUBiKwGV5NGF5IJCHCc3p/huHjH8yHTjWkDIY2RcPXRJ+XY66
OcKo7pJi9dwK+N4H3j4AGIQHEDubbaPBstYT9Dpia6iOlhR3ShujE8rMp0WiY9nLqey7/X6fesDL
UGJMHvuyOzgBxxzblZmX4HJ+cmtqRNsruzbBUlkV6Dp6UouFg6KZ4cU3pFNExOgjLfX33y4NYuJ0
6Z3ZEeI3HvmvhSu+GoE5FsOnTLohcK2y1mdT3nOPbV7BSGU8Yx/mvM8V/tAEvEIAQ0RzhJqS+aCl
UuuMN1rPtIaPKjZSoJGn5WoqRiU0u7BtBFCQUT24r/mfGXSIws+1DEbugo7zpeDBDnRHEfCd1mmR
bpxoJ4owwzjtufNwJjAl/vz+pEW3/oIVMQPewGq6G+9csQLUWAqXwGJnSFX3T5/E+sIw7BaUFFiB
zyG3VETq7W4ZhrCdItX6WY0oJ+FybX5ppMznPsaXGVUkFbdTI/YM7PMTXLm2asHdqZdOcAZdkL5K
CXJ0tEt9AT0mARRlGLJkhiAlRFT4pHCG3IJ7mRqok56vJZzOriaTYTDFpTOoZXfOtwj7JtxX4D1O
jR9IR9QLO+dCcBI5tsNFNiE+xxk5UzL5447pNlu/AdyFVwqTqxNa9vZU/LcaNm7FX1LnnbyMC9Xo
rGgseYPOjVqF2BwUIZr13Xo+Dm7ugugbAAWCWK4PieCXHOiI7pTfAwRNGGtniibwiJ9HIRJVJSGJ
bdL8a0hkmEqj4qXiwFMjYko+qk4gbX7fzPsKwBy998jQKB5tf9utwNdLleAkGf20sFJcsrtM19xq
EfSVKi9JE9J7zzQXE70HeEq/H7YbRlQJ44JVNkSvu4ta5PolJ8WJoKe4fsKVAGzCZhGAm+zw0XMm
PC+F19uwn0Sep8UudHQv/6osRxIw2YlQ0AzYXcMRlEfmmdDeYtb/ME140eq2QQmA9slJuqR2P9Ei
n4wdyqOHqwWZQZJMhnWr9r8W5UwpnateGrt/YKxk90KwPqqfR6eI7z3txz4UZQZDiFzQpPGIU0qB
5cnSvufF52bpko5RIFXVIPKOXDf7dvVVe6OlO//XMVMyMGB6FZnwTroQRGFR59ws0dWWFsA0m7if
ObMLZDDJa74PwWqVlVxXHQljHuPnYAxmbiCxGm4O7p2d6uDXT6zQXVjW4FTW65xbH9/e2VGTYhO8
uwp0EG3DkqcLgWyWQ6+vzvPAEGzH5/GJrt3OgrRUCOHDgJ4+M4kbIcx/c1fCNxU+WUu9982ctEm7
zSrqQ/gemui9wBf+I985YLTinb78CmBw15pA9FIeUyM2YSIYkbO27LM6cLqH1WwmTND0mlTp4LIM
p0YgYjC6BKfSHrRstS36KLQzxyBKvVp29qsImHghNPT1oM6UkQ0+uibdipd7BF0eGjHzzfqE6naT
kel9vCyAFM57ZfGTR3S6+vGJZ+EPOoA5uq4OjjbTq3/LpKFh620seC1AenRKmAEugJqPxMSNxGmR
KnuzBPvmBNzMdZl/l9G8HX/V8MYsEexrvxHIQii7uXoOM7oiXnyG4I1wMR/xgXdgYuonaJvYUdKr
m+IC12gU2J5QMWoliFLJZq//bpyGSnb5UDx6rBKp22j99hT2azpwBuY1ASxi2Faz/GWGYkiePGX4
HJKcETBkc7xIx/u0A88LVZ8N1ojhdkFfVZ6DK62fQ3u31QfeAuQxsJmykE8NrOLGTcGOXGE6SWEZ
V6Z8nK1ZklbDMBUn1vRFKKyw47aInczBNnoFLCc7sQWFiMkZRKUil1Yd3fMTkYFxm57reCnpwZUm
ztppL8ZyfgitwrHC99OqjGbsKkYLnoeTbFrvsruTLnSet3li87Rnshg/1NRtiO/tF0nAlSJt/5+i
xlJndn8MZPVMJBt8G58HC2t9H3v5yBZ4jMO7rSpM8uWFOXVlPumpkn1a0lZ6/LURDfkXDesLi4vb
eRhvL42zqLnb5pHZ9YvALhv0HXMt1axPVm7/O+Pi9Bxd5sUfvnhTTa19HOXwK4KNBSH+nI38EcJM
rLj80hHm22eDKK2V+bJOrfgTISPrcYjxq08GrKP6P5dsz2fNzfO5P0+Ug9HBXny6qNLO8plD2GAy
EsxawTYoioGigIQQUecSIf53KXu1zyNuSmaVR/jtytHZBo+7A5DRz3+Oef9/u1EapxeE3614OUty
qnnUCe0izt7XMSVmWsXk/D/uwC5W1lxqoH/XCDzVxgjadUj0a5EP6OD/3ViSzmQAiviQhrMAjOmx
VcNTZCasUoFF1OKWHKZVOHqIwHZQ2CGtSUZA4yyaXDkFxOia+z5wxcolOwXWLdvHCZs70kIwqNdZ
AMB2RbWS74XUC44UfcrM3MXcniMwlWYzEFXMQKCaoggzaR4sSk7bHISNtfuFtJr18jVtsQron+U2
DeCJwwTkgeFZV517GN7wxLxKTO5GnJIK2c3y4wGhCwgAO/QW0+lhHukd0KvZ+igQhFVGTqEkEkpS
EhyL+KG1HBtHquknmiIoZJ4M6ykbWxzYypxpXJuYmAlR7tnUdGvvnRn7uvQk+U/Knx7uq2pnatvq
uCCh6vUYmC9C5gjdwX8MJWALcWKEXyaKJB4jwG5OFdfiMc7jsbaVUS+Asw+Wca0WupkJ4RuZC+mo
r8nZEqB7l7vXIBoogO1vDcKlgtaiDHaIkMbE6CnHM0YRGv/0p3g0+JXiydyfO+gPBcN7Wgbh2BP+
B8uWtFguxVozpVs/MjUC21qqgrW9NDfiH62FR3VT/uhI1X+kggLP9amHus5po4AQnKJevB+RWg7k
V0oRTpIGSZG2aAZbFfv8kppo5Pl+NnZBrfZ397vsavEuJ15wblK+EuBfQ1ioW7l4S9CdM+Nqn7rj
yi9eEcArpAkLbmNWFTH4bVp+M3raBddrCmYqHbaHO8OqWVp7a0oAZgvspuoQMZ5lV61rYECWp/eG
QXOEwOCo82DZGgiKPgN5MZtC5zOwpYNRwpb+og7lzS6oTiY4H+xmBrvbk1T8YexrPK/T11jLZYdt
VWCaZJGMyd+wHndZOGuvQw+UGBmZdefz/OjeIO4R54J5yAp0c/sblyeF1OQbEcczX5zstSYvfsPY
q/1EMGdrOR4CZQwEaApMO/XGSQ6sx5Ur8wIsjJWtdA/PPyUSkRRh4W/2YJphXYu9Qk5/yRn73jiS
dLB9tOEJZxS0PO8qn/qEDyJ5LrQVxEOOvNM2F7s86K9oLR33UfHipsqj0Vs8MEozWTNn1LSA7Fyw
GXNFFk9L49aUPoueAq9AbDs7Eo0oFPZzJPS/P4gzjb7vHonF3R/nsqNfVj1G7JNQXSTVxaDM1buw
jBKAJc75+nB/Dg+CkccfLOFCA3Lb0WnpnbZzK2R34WUrvKd6LiVgnymzsuqdKpSNkyyhCHf+QONM
uJXxp28FHbYy2rg4PoyMKDCXk7Tl0c1sA1yYwOTTvK6E2XeSgbA/sk8HCrWMGOSmviT/sfjJQ6VQ
qTVc8OyTWzLe9xJgrqCjun1H1VOi2ERdo2ytxAlnKG905F+a/ZUPW/7pLRI90zOd5bkRz19G8jCW
2eJHQwdbReUDFm5xS2D4mAWTU9Je77qswjW4J8RiF8vWNJtJuvuLqODkoJX9rYMr+j1UM2I320YO
7bfvRWhmPgeoRAVMeXawOj4mof+nT5QtJPKIbZclckoKHX+FJURtddgOkS48PrwR/b8+bIuLfoBb
68lCuPSBcMRWaykFl66WkhDNiHgaZvNIo3Lr7XaOERppinOcrt6XyDHjOKrPtRIsCF6q89jdGqAd
eLqdl3rpEMq8sOeyKStHxJCyRP1k4EidEzxaeRoy7VInSCdZ9L0eip5j96gUdpuP8YGvDFko3/Mw
tZFvnD/QC8LR5VgAT0hzgJyMSM/iduUCqPHk9QexWv1NvUNBt361Gx20z71U228xZ7DSiOueFpfL
ZNWR0gSU6inc6i5sGvFrblaFdQcDnGNyHnBjhyjnhr3RBJ7P3e2bFfujUJgor3TOoyUJ8lvwdfBV
j7G4c5lczmI8wOw+qmVv+HXLbZbgz4AdInLyQ/47uwfZfZQfOjA1voTPCpPDMLPdE1apdEKvtFvG
oj11EpfD2rWTSoipdMw5xFi1teyNm+xWbQwneKb3GhsjDlT5u52yTAoOB07MRIkbkRGxqgO+Xgtw
tCvr78fjOyyF/V7dbpOysXDxENXrXKXG3W1nS6SfQwe0TVbt1UpPbrKssvf41AgdrmXmgWoM94pm
cY+UXzmNsneVVT4GeXfYYLZuGHewG8YVOlBTVVNbnYTYHvvYujUl7S+XiG5DJ9QcChISflqhHFUm
XDeAFgtoHGmKQGktqPbxMpTLVKisWd7b4gtLDORHlFshO9Y4qzk47gMs2Or4ffqZSL1V91ewLL5g
SwpOPh3PVAYzTu+O9Nwk0B/gW6W8I3WKGeatuK6z/37nBXyLwzJHqBUrKc0dVJQxmX6z+ZLm50JP
01WLWsujqmzy7e/FhacNBxXQT/CMuhSmaM4ui+AuMZSq3e/nMX8mImu6broReYfRB66cceZ90Gkl
wEJ048F7Hua2fiPBHYAGHhvhDk1HtaP/Q4Fg0dRQ5Dv1w8YM2vOflwg0knQTZVXZHkPZp/GmfT+7
/6FMJX2fDlAeKGeJqFkszttJG9XHM5sBwb3efObnL+QTrKhMV0pXXlDuOb2I1Ktdl8vfl9KI8g03
GMLY+o9saFuRPUNEBTJSS1Q2uLbwCT1W5rJkCYl5tXr+DlVdxNLu38eCYTBum4ZrrwXs3BX/qbLl
o0agHiDm3a+nb+kqCqvB/dBQ9gndNl3ALRURGOzE1RbjykMGY12jwKvXzaQ31v5hCP7LiNfenKUY
eUWHFBPD5iYAWpLIhulGqezCGqH1DcbISDPQH2qfClq6XOh3xtcLZMaT9XqLOg1CkCuZjqtSDBSF
Iyk+OqHbPNrUEDAJl6EHiQ4lcHnLgjnL/GBkhVhruUyuovGcM7GRGCyZOugvdw0qMmC4Z/M39PSL
L7Pfyl75ozg1NRfU7WWIJ7zaDDBxWSq8dzB8IY9YCaTFso2xIjLrAeZJjLAw+iPQRfTd/Vn+1XW8
UdrlFIXDUlRL2+B3be6TMNVKoxVQaUO8e5HF+ebOi1WQC+GbnHgqjuJE+GvLLQxmAz8SQE7620Nq
Glg2aYyQneB302OzwwOw4fw2TwP4P2JV9enJLh1+w1rmK2n9XmKiujCTDibEHvI/M8QEJrf8+U3L
Kj0ynj5daui8n3EJQ8o81wXg7B2tdbqfLfT70B0/2MNEv10UnxapNdpxP2mCZAPddHelqgM+z7Ic
0qRN9xyEGuFEDp4cl5PA//1u399RtE3f5npkJk/TOSkXActqyGoRvzsBjyZonVCJyEC6JpnZrfM9
bprMavaziErw5JLSsRLAk/31yHCwYBjbHBC6hySJTbGFiuMyEwMY1AwTeBUG0I5oE5pZFrCRj5fm
l2ddoHaHV9KIevzzQG63dXtHE3slQ6ot3EKlKiXEiSCycC+xexaqI7pJT9heYHx6aNQR0qH1iYCK
1/y4OUmusTsd1vc+qPSADjx63Nm9RAswgyKBWrsspuyXvlWnSZ0rsXNIAAodlMkdfAKV4qnKgE7Z
4Teho4RHoui+yfmV2OT1+GiBc93bEuvQJ4PTSeXvMNCNJdeYxLGBUajrMmJQlE8FZeYTi1rqMqs5
xFxpD4sPVUF4J3n03KZx3CSoZFs17bHP/K3eD3MdD6uGEr5RWgwR+X2TMpVItoQr4ipzPVR1C2ea
CJqc8V2Rp68wrrCuYxfGZR6I5NR4FBGMufjPBHnFeT5ebsJSaWJmksAARJRHmx6mQRUJnhPnOFlI
3GDJaIoRXkEyw3gR5hK36JejhkJTBvjPf5KLi8RGamERY5RLvul+yfyu/tDo5OHLXRYquLHw9nCs
/QZjY/f6mdggVcqNipLgdo0qjB0tXWqTOl+WvNlYRZ0kqTXe3wSFb+LM27ZoNrV/ja0cRqp7MNZn
RGflU+Ks6G5Jh6375AOiAEWueL7ZWeR7zyIJeK6sedVTBGwpZTTEdZ1OBWFd/dKuRl9fpnkHSm5X
DCKBQo3W4MuvTcDm+ikVcXLHKG/T07upKZj8tMT+VZQ20QueuDQZaPVKWZYdImbVcYP7NmrutgGS
PFw7u0GSxrD0dF0Us0yO5o8Qiu0jGsrZ/q/D3eWXTpK225FjpdUVwTRoc9Y5BWKomqRHFmnw9nPX
UW6z8cb+at0aFdQ02KJJUbFXCN1xASX9f0YQ/y2ehCOH7+g+JIobUXzqGv9kz99Zfv32oKkHJwgY
o4KhYj4SxfRDdKGyAnnzf/4ANz0b6MvU1xhy5iDG5sk2YtahVj9n50eNqWSeHxMIdpZopgVs4g9h
r3oCcOcCg+9qWvy0/3K/nhr949hy3aWZ/u8EkQXhIN6rmUZtNVA0BjVBUI2teY0biK2N/zl7IZFA
Z8CNq3wKVWOSKpEkyyjDGoLncUg5CkhmXxpQstcJSjdapKtJ13rSwX9kfE31itnHHTCvDqPsSve1
vwe0Muc/TbBmwzxhzjsj8CjZ73blRwn8LpI0ObtSoqfof3h6LyUzck1UytFOCkS//Dn10W2/Suhe
jQTqDyUUqt67djLbQbPEjsa+hYy6XBhEuIKOFh3NP2egvtv8quE2XTaQku1jQTa3+lronew82MSO
MqPowc76Xh/Rne2TEY70iOHB1O762CpJEslbztxURGDNk7fuJ8deMkxPS9VlugrAu7LxK2kKtR66
o+po2xS9Lf0g3oJd9Sh1tZ2Hj1CT4T3igxCF8L8CFiiPSjUG+bVr7R8tdGUj8vHuKbd4bC3z1KNy
O3ZF1AUh5oQTRWCEnzEsBNR1zz0g0DXiRVR3pd4x9O5XvC6mfj08i8rWbb/7TWxh6teslaqW3lZR
zmgLtk8CBo4GoDxG7w//ffH5JM52kUj1MZJqcl4cK/PqCQLSP0pJm/EV88wkjjkNRlEl6M/2SWms
aDg51iIB1RwM24rALWhiq+9J3drKawG7qtpKMZKievRYAuMPkGZ5Cc+FTgMewafkErlHHIA3rlzp
41FRjILGyWtt1NbstQ8TNfpEeDi09ARx5VbQBWUjvTpjjj9N27puy8Co5doK7pnwov/XsG/RZKWa
MDo5qSeLhCAiCH0jtXHi8ui8i38EzLNaHERhowitSBt+u/viAJPynM5Kilu7Hyj33fXvB/x8LENc
9tfkzt2fjOWYD/7Lzd57xiKPDpdgmueHvMRBVyvnFY+tspu/VQngHGgZIV3ZlJoIxRfEgifvT6RM
VN2hxaxtk2O2MG3UuMeuMQclOtE5bngR5busNqEOL055nWxNRBFlA1OeEmTUCsE/7+tbUmD9spaV
gmpkiJZoy7mKl8UuUOkZ/+UFfUoW5m9gHSQREwkg+F/tM0Cq4huN/mAH8EU6CGit5ctVXM0Rz8FI
LSCdhAHSBYb1wVQQ/l7a7mlapJ6f+O82+k8vt9cYPZkPGifD/LjryzmKorOpGHOvTEp9hLBiON+D
yTjwEbSoQfDSqhYTeDjv6aH/5V5xq2VZsvyNY9+8d6e8GOiLMMIIbwx3cf1vXc87wM/engXlSfPS
BRVh0Ehysk8HMDjr8i+pBqX/8Icul8zcW56ACr1Pquvk0zR4ocPhK5gCKS28CR4S3XL0nvUP+4g6
3CRueeNArrkbyWdRMkVLiD9JKVnrCYNz0xXqaCqOapPc6jDIM74qThZ3HtH68fIECsR8Se5u1Y6m
4p0SqcohbIeA3ihoFe92yajMJ5cUu5733tbqTNjjPN6j5+5827Bu9KdewUrCEGPMswTElMWmC3JH
jj3vLtcOyOkktrDu3dewXHvtHsrPLBQYj070/fXJi2zdmlU6pMjMtipksu90/CyLfeSl8Sws8WMJ
MtsSSnpAmUAhztQ4vnCvJFx2iwkoSl+aJ8ABrJYxLO/3BK6Pz1XqhV/2EfbSfh8N+xBi2XpPjbsT
2ilWWzGQpnQWwddBwl6cPmF/L07Hz5Wayt8N3fkG7AueMcuwMwxIpKxuYrHhXNhOXog/jX/OZe5X
1GKLpnBZCim9K9zn1zrJMuFjrfPeZpXPrJVJxxQVk8MjFdKi/7lDN6jT9vEvHIr5Q4ewkmDnFXXR
+j7cPsa3nlVVQ0ryQ7kEWp7qm54048gF57X45ZoinWGxORza0LaGfh4nWjxKDM5V/uJZuHZIqIv3
GnIdGfkudZmdJy4TmBEh7Bef+DKqrVWWTUZgLl1zUCd/C/oCF48h397NMi9gc81JdRtCGfteF8Md
RHnyA5Kx+WKdeCcdsrN4U3e7+QomsknMPtH/7kBnT33NiAoM6q7EWz01mNaPo49G+yKxtyKMz1hd
efkE8kBObhNWYCdNCKZ8jcrGHaRUSgRL4xgKaKVTdgmOt4IYkO0dTTESsMTKapedDpQSTr4rJFpf
pg82yib1B8KWFpOs6xYRujkV0VJ36WZk6JSwR7I+n9K/OdkqONSRTh4bevkuRrMU47Rwoxw5ltOA
Kkvmh4jjD2ti1PmrBOeXTqbjh+q1cxwAsrhL9acjise9wa4THC39owuEgGloAAsKofHzGAXsn3d0
KYpMA8thNmDwxrKqw96Uz8AT36yHhJyjH7lfuIOJmN30OFDAivDoxkjupRYiXgzWPuQWyhE1dttU
bbycDEIOvRGsIesJxhNeAYVCAPrlxIVGQydwBEl0L9dpPUilMEXeeAc1wHC+u1dJ/pmV/qGzp458
t+ek2fWobMAnQmS6BH6UdN3KBPiki3ScYzST7MfWD7Urpp6XsfaiP4C8hEaAU6qBLJlVvMVSgOdI
0bveU0FyNDqi6es1HENziwBCQfCgs1uTlJKPtp/83/rmjYLMlyKriVvM+Cff3zBTp2e4TyUnX173
IUUPetjFEtvVArFCu1uxpqD+E+pXb1lp9c3QUAO0GCX0iWtbSYRWuUFxGUzB+3nNz5j9/tKcoWpW
mZWnriXrnQRp/0IhcQanaAfKRmbMnnKtmpa9n0exqg3hRWd6lQYzFnmpwuYydOFBEXJLI1zh8L/6
NLsqS6rVRQURlicFdQsRkGs+LqFsUtio047SVFyqqJS58mMf7y3CwyKz6EUbmFke7mkdj3ucGbNF
n5VN4GE71niU+K8GmnwDuZVbxWn4ZXunI+MsZbydpoqPzg+yHOovpq8/3ZsOR+EJgEHAcoldc3NU
sPNJyduhx4VWpi70BlCedC81ompPakns3271zzb+zGROQiD2RTkeSjyLxCCvseq+jMo3sBmMmxFR
B5+ORRcG9hp95lsSyrENDK84uZcqf6BMGyITymqM9JhWKQVVIlO2G2abvpFdN5rHGmzhC6ObHgDp
yppGsDRWctYCJG16j8jq2Yf7m2lldVW4PNaK0al7zg7o2RUJ6bTAng/3rFXfDLuXfjwj8l5YDtTX
0HWW7AhXyIZwAnKc/LUB4W9g+Z7mvwnpC6swcwwhc4cX4q3KJr+/9IjwpJrbGavjOdbdo83ffpzt
4TlDBpgtuhgs+sQti2MOCE5uzIUXeARK88qBVSjKIhTTxHl2GAiR4rpeX7o426yt9wZOtvXlzZEC
m9KMOv4Fzq5hewWDqNsx0yCNyI0FtJhXNDvDBcDDgOQ4287BfR2I+FG12XPaJTxPkY4GL17esBYV
P5OD2fSEcc06sTWlOSGAS3Ys9MT7hg2NkQxHoyP6zjQUTKzxjN1bY6MBYn2AS7HtNVxlMoV03iuQ
+S/ryGzuPDGsJfI79CWfXnaLcXWP/8nH5OtP19fxdyLqK6n6JxRgVI/xz5391nRul3W7S4ABtXwz
Jd86qp5ucvQ4IApYP/qBmuSD7zKgXSIphz6J4m8eLSOGiXuzS853d/Y6V2kQIhrYkDc0V+x+w0Pz
XbitmRi6+e8Q42wRizOwideY96WcP/nZpZnEaZiIxaZMaBBx39XvK+voTWko6cu1xqouWXwpKjBr
EBvVNuSdFf7/YmgqOq7Qh8nVzasG0S2Nfr2EMt06SuyhuyoCj46D9RHSGLlaCgkN0y/+w55Y22B1
1Yg/OFHSl9DNzeth/i9L6OABsl06+KFiunt6KtiIXufnPmzLVMPPkM5Hci6QEVK8lHAcbimQxfmU
iiaVe49WNjCvqjdClBNuEgSjvhzdu/AzKdmomARFKlr3kqkYogZzw/PFP2NKp31lUb2hjmxQ1M5q
xKZge5yqO/GAzpFkt7zx/OChYaeV1N9ZRD356FjZyyA1y/kgs6wHyY65GY+h+s4NANCxGsjvjf+7
4vPdYc8qXBfQMeF0dpH7HH2tztWmmIsqM8vMCchd10Lc04TavIC0nfNFaEEq3jyG47ct/QpjhgAQ
adxFLNwnuazkD30nekY7dP/pjtaaR85mFzXiDnp6BJ5hgPq5mnLPm91k7ka6tq33WMZpd98ZBRZu
Al2u2RzoTom+vjp802Su/OcksvavuDadB9gsXw91H874Ai1TcXw/nKY/rtdL48JhhRvtVHUAgJy5
npasCr4Oo/nX1J3JFaTFltkgDAPAda+KahdvJ3smxjic2PMjA6VJ0OB9CM8ikp7PN7T5iajMUdp4
KXlsyu7uXwRDiJv54+AjzL/QqsiKtuKRPiEh9EBaVmxw4n2I1y3c8n+DYhDQjQl978R82dEMe1tY
MBbRuVXLyzevdajxJvCNVJqTDEQXWPFldl5CuYFtir21B1nDHYWa1s5ypI92JjQ9Cl5OSI7woLcm
/U7kjg1bWa68akJ12MxNWPJCKBODS9p67ylW7k6XLL5bX8EPDK3FBvQSJPQ48TXOnjCS1Ba6dS72
1PH0U7ZE9JVHjBaTP7/UGFBAHTcPb9/r8Z6XOCjcJw33yKvSAqK6bd/zYIYu5G/gwFE/aJykK/Rt
LS5dpSvomeJocYsOwYjOfqd6mXqN0hq6ZY6XM0qDKOVzHkpzgbeplSoQ9GgCU2P2+FIbaurfpNoH
o0cIaWAi5Q/hylfd7mXd2z+V/pitt3cf+gL2BYUpr8bWfCZrkCsWT/EACkY+Tfv/O96zr+lKI4da
vcMDooMrQitz//6sZhljt1lUuQ7wfx1ioIOVO4i3rfymlYc9Xe63BW5foUQSewKuNsvAQSW4Gzgr
zDF/0xGrmhiU0bSejGPAhnxj9MMon6yzAm3J4UE8oISidRaWVJiD5hOZN1JhxJ4OQKXwuj/LVsqU
V79sRXOTX9FDqFN8WPzFL17MLWbBm6blfbHEMSEko1wMD0BAsL7I3gVGA6nnQKTsSjoFMuGLeAvf
gElNwNz5AD3mx6fNBLW8lRMtM3vYeb3l7HAsHarA6iv70SCTz5NmWLJGHEpZHW5+0l47DG2GES/n
Bldi8feunA5G/8eeS0dzdxHrIkzZqImpdLH5GnV7iMhrFzw+qmuZMzVxAbXvgk6N+tx4IReRIuM5
LfKXeIhteQzmr1jzrRzP0p7MoEJg1awvuC+rKLyY4Qp5M7hNkBH7L7Fsi/YniPru0FOvnTrIpcyS
8kFgIDNrK9qP+2AlliQaASK7VeWDMK0VmAKRDnCkLHLdsCaIjTkkeK9v2oNoJ2y8D9/BGgMgTiOX
ZJJlytTZFnnGaXLPVDsonRQoe6JZgiFlG7NTVLvma4ocPuduCBeVm/DspE8n+Kc4yXxF6vj+1iLz
GRytsRBVCikDo+p5GCBClUdVI1v/HCg7lg2BHYvsOwm8U4kfODHi9h3vkY1wNWRCQf+rkClq/HCl
yVf+eF+4/lFNMIl5i++nVcHKcRL5cvkuLWoksIifWDIBH7kYmh2nRjoiha67ENF7kak+lBgdHMfw
46N4KIjqoFGQOtO4yB0WcNpT4pfaxCW2IrS5WU32VPAtSB/CY+1qxfUaGqVph9l6bmPl/o+PPgsD
sjXZyPU1LeHvYkphzpJV6EYStAbDU6eWy9h/8Et52qBHClKH9/ZUvfe1ZT9M1cZCB0NUud6TpeoQ
edHabUCyipJp7DZr4EULrNmiQp873Wnb9bhauCDZNIEuF45EShHwrXdFUr48BbMEWIngYIEyhJEX
AHM0AOp6YknF/6HTucgOrdvUiB4MW+CkHonlI6zB3azWw30/6zAXbBxmY34Ofq5GWtvLPw57xEzF
pG+4QeXTzhgq12hx5GlFpQjJ8uPjDXHuY65Xuyzfmu0R+SlraC2PyKrd2xcW+B2FoVeKXt2EgC+X
PVfMXfg3jrAPo8Hz5E4i1ptzRMupXRr4i+1GmYRaC02Bje0y3QzzaUp/4WBubzM9zKoqFtSHxIS9
W60VFW7Gkyf7FtTmqZfMsiSZoxtWfpxzSwlNgmMILFfArpkASrhT37v5WLBV0yJ5TGH0Lc/+r5f3
+BFCdVMfAtqOWipUwa/tr2LNpPWA/TDd4nFq7VkaBERiQONlCMv5vz28KEDfdvRLmmZX2IxKPtvY
6VkcOhD83gYsODWBx4WW54A3VVNH3709Q31pMfVR79AjuF6jk+XRrkapuJ5tPVHMUtzoR8U6B8yP
SE8zasXWKZEezag9LY0t7ETR0FZfyNU+npmrBftM8GYpWWFlibWJ9u7WZ2S+8NUGTmaMrph/KU+K
jea1OFAMWdgf6B5FFsTyKGBE3L1QF3b0av9fTBTKiAofJb6w4pFw7DNk5ABHatfC4gif/OSJpIaA
Qh9O9+Gg9h42KKdP2SHUofzdpQwZLcIsuLYuRWOYpN0tHAxEZ7IrO5rkeaLPxVv8ZPO0c39PpMEp
VynA6LOGSEVJxybWWmMJRN+fHddRXXt/tbggb/AHiDReUAv3dwUO2w+u3OBJmZYFFAirSzTs59U0
cfz1vuhO7NySCSLqDTimjxp+NJ801mxz/wcAJ2mDJo/o4SJNeOsuTOcjYp/bUOq0qhOSFFGWUAue
znihbco5tuoCYGNoYKrnE1VFZOReoTY1KDXC33+jjvf7KEZ/9OX+7xo0aC+gSx0jWuCrF5ImU5Mc
JgNcY1Yz36h+F5r2Pjs3Du5ZI3HU5RVFnjuafoT+fCSMY8GQS2bmrh+iLPLUVVerdkiyPGoTUcFp
UGk1g1SpKvfyM6/AVBTZ+mguloWCC+LnvYlTav9T7+NpTPAcuzoWPMXaZKfNeCw2tfl/5Q1km0gK
luP/svDK+x98CHW5dRG1exw+l7jQYgi5ciZgMBF3iCZ141Z1jrFwTYnBYXzU4cYrqt28enyt4opG
/7glfOl81Tfx7owd6ppdE2sxDPPHVrh1XVruXanvYPYEykOA5gXteJknX9+HTl06+INalPNNK5/i
hB0yYbPiFALu/4TEND4hovpJbglufs8v4Ld4JS9mbnSWZ3Zd30WTMPv8eSPgBy5+6nC+nyrIp+9z
vdfivJa26ONQlSQQ/BWWeA6i+mp3TXchsT4fqs1WkhkTJzVdMxyDuEj2YiXt4kld7qDRaJdvDXMd
T5W3Jd45nDdeuQrqb0VqSeLiuJJC41RQQ3Lp6b7gsdEpX3TdmbKHYQqJoKrFa5/VndOEslRmW94/
w/A1uLXW6L9WpbIjn5kilrna+B5n10iKNpHEYfhg89gArAhNEyJkWeTgmlOk+Mb2WCKEV76lJn9Q
3RNEXbrUK41GHwTYobAwd1+YV1A7ZX3tEhOY+mv2Merr7LegGuN6Ttdto7Asw5ZWwkYGmZfUdZoN
AUKwdRVu2Q4FM2yvRP94d2QT49W1wDifKa+Dd6mARbaeLc3Yf3i0qpkOqkdVLfndJ59+Eh22c2iM
oyOTECRdmeEbSYzUFagwhw9DegW6hYTpRJkOahS2s9EoZwPAUN6HmeL/y0/eyFR37FFXv4d4pSv0
H8NnLvJ6LMk78uPfX36y9toIjLl1NP77a1OlPSK20/Eu+YVWWKHox26iuBPP4Ggh1E2Qd7v1WyZH
g4QHGXekJAZI0u12zI1Z9OdFZunH8w2xeNbsu+v/zqHYWB8cIc0nc/9cIDUHSTGBxjg6tHRXongY
fcE8/rRa0qHJM/UGWLbHXBSnqU448VhigCmDLgcAsYe12ObtGeJm86tx8+c+pAjAx2NIY0KaOsMm
4LN4RoRplorbiNZVpXA9iFmYA3sfff36+tLlwQJh5wIOUiIuTmyb1Yew5L73VMlt8VQkTrmg+qdb
4l2qHU9hf6fFiMFEh4oWlE+/utfJK4ONNiHmXJi8CArT5VVOxRXX1j+iEKcMls9BvcI6Q5gkKv0s
cDvBJV1TD8GTZzdVAM9dOa9e0iNId3O2ZhoLdGvAEZKrCg8lsdeEW9dTAW2Yh5wIuoU1EGfwHvJZ
P0II8Q6iwvIP4JI+mfgEBfcKcPA8DcbQ/yBEB5w2vx4S0VEP3o4bjdNwDMu/FZnBgskM3dSkD8Hg
Pse18F4R3nYlkJesaS1KJ6LHBbWNi3jzO/OMUo0Ssvd62Vk4SSjEb6ybzAVkodz0WKKnYY3jqFT7
KALNEsFGa9WJnLQ7Ai3/syWrwQaU4U8Rmm4WinsELtHg31zbBDRxwTkwH+4tcbRkn24rXADOcPZy
08towjSTXgyzFA2KCRwE1yj7dAVV2fE+nvLK+c8kRv5tSTYazn5+mRJHR7GxjgXPDGtrnsNAkPof
ysMtAVqamHWwij5AieH+JA7aFnsWX7PKLpzJ1hqIUFFAfO0sCZeo7F/x4WXL+YFj10Ndgr1gZTlK
X+wB0m5wGCfFEp/sXxrqDuNQ84Zr5oMgTt8HDevkCnKQ2OYHiSn7EsSFIT6hfpjhX/zmgtlUl4gT
2hrQ1TqhWcuDdHliotLDEoUutboxI7/P82WWRMQRSvkJEfu+B/iYFF8l901Nu6PdNx1SyP+g1/OP
dzz+tmeYo33cluz3FfjkgHy6kNQpzInfFMpOHEv5KRRX3JXS2zkzZCjtQSF5NHeO1BAfLvuhMU6v
BvX1NR5qnq0E+czWi1P9UIzTXNuILrZsUs4N1FZIzoCB6/o3pudwd9wLctmiUi0SyVnWrriE/7HW
kGu+67TE3yqLFDjJlTduHH9haJ0XJWYQPWwGnsfHagJPX+ybWZSWmxVigXgyL8cULf8NPHpTmM5t
9O+l+FDA6pdCkZfT5UWHTPAtSBatEu6bZ1Vf63XrCI2Cf4ofMAJ4CIdGgC4bwozZKAqaDY8psLJT
0leRmbUYthiZNC6srhWgCWLNY8dsX/ShDYJ7OpjxdjW+oRBf1PPlPFcDPZCBT84AyPjerlt2PXc2
5cLD4uOwo6IVhgoUaKzB8fWCKdVAyq6BkJIrqewKD9Jpz2EqIZocp2dXXfZHpm4CYD4sOkqCDZ8J
OMCsnbYP+Tew9gKQaQhRGgnzuMD5z3INASTXSKcuPQggT5hI4GSBiQhnvkZZO9fArP4cDt4jMMnz
JtBdiOf6icNSfTlaWasJuQy4YY83jTCstGRnomVCfUkaQrYrib0pgfzp0dHVf5de9sS0zP6cQydD
0dda8ugXvaJJtw7WkedWy56M+bmVUIfm03bRu/Jo2xVSoNQsMwAGUrq/+tABturxRzWBOrlLpV2k
RaqASTF0/f0u0EoZx9onKzjw9AThf1wWTRdsss3+UVlfpA1+X7VA01OOlxblqMbd6dEOEwcuTM3m
vLArdufKPJrzL3nWZc9mMdHY8ka4KZJe1QAyK4VYMHBJIGw7WhXQ9vdeQroPFBHvZAZfbf6IRrb3
NXrMNdeB46ALa5q/NTB+YrYzozcD1tZaTkF7J6uRqsU4/MISiZBr1wP8VDUljdt7BQ/AUDmQLhP2
cbJJgoshspYVuvmPpjlbVmPRTmffTNV3AnYWyqZhp9+DlsR2UiDqqGZxwWbCTHssxOY3CXD6/6mX
jw8Un9fc5K28Hn+LbalR2TpurPNLfeC1qauCM/nzx3rI4znOtuP+v+mRSHL0CjKViuLsuCMN3SUN
3lbppfsfmzwTzPIjuw5E1DTfbL06sDM04KVTL1qMM+jDBoUxH/shEhQvZygjdD8B0RYwFtdsgZZB
Qb4aql8kYnI+jtkQpZqyqQMq0cFeq3sWZ/lULYKMaYl7fmB+9EMK2Az9bmTGBJwmurExB8iCV1ra
zS9aG0Fn57P8JcFvxxAmb4jsr54MqrVB2QVIjCe3mU2n6Pp1kdnl9Iag7UNxByeGCSFRjF7ZyT88
geJJMUn4CVrFnMYfNqMysQEY1AeiqYtJcwzrx80+zJQquDZ0Chpm7aT9Gd9GluEMZcA6x2C8fdSL
eeJ9JXLmgn35Ki8zRevGmfkj+K+fFLbt0GVo7M0rmGvJwZhBBIyiPwinHgVbY+P5MNUrhkaG/U2b
CzECCt4npFnL+7NrHk8ac0bsE8xHTgbnifL1U2aW1jSEHre0ma+ZqCKLiWTzVgYYdKrGnyFVmOFY
Aj9pMQtfep6jHBQvpMdb5bdOcWMuBHGbb0mFHaO/2NcdDhGOIkQGE/mFuBgDH+m94KNwAPrfVbBf
cFrDxoKlHhmBXN+qr5/PdSID1itj8GFDtWH46SzDWW25bky3IDfRMDiS1H5nIyuhlJFl7GajwxBB
kdpqOgqUYe7tyVKoackQbN9/NAjL7u9ZENCm/WhEBt+uczYg7aFH6NSF6yIwJ70YKTk1tnz3+ZX1
acOZOKiMHHPPRUDr34TD+O1TN5e94lUPqHp/Rj9UPB1r0P01POYu6bKaAMu0dmBBLp0Tdsttu7Xx
JOcVhqfJOvW4O51qCqaErqEqnwGX4QCu99rHjVmMPtUyFKWQz39l0uIXajj6FenBpyxDmHHLbjR7
m9+D2BxAJfeLFHDCG41o4KXubXU+Ozod5zVz6FArGRtUYmknoHjgmSeskBv+LtgsjbkTSMho8dUw
camq5EHBLQR1aP/zbB5899+MiU3KJd8GEOzZ1Cm9yxwABDIq8mwj8nWhUfibGC7NCq4hJozzZMp3
PW/4g+KC3wxUkqZyvBaz/kzbfVaoL/503Rj+pVbtyvxNzGdtPMQBTUxOB2E6j+x7YxDs0VQ4MZgE
dpbIgyD6oinRfgZEUAQWabgQ7u2ZPQUPDiHTBn3LOG2E2DgqTjzwk7a8yilK1tl7P/BEKTR3PQEp
ACNuVL7neK4AYm6Y3BBCRDVHhJAKwSclBC616eXW82rEqI8/3DlB+RR8o8Zh9Kq/rq6HY97KRQDn
TevqPCpSRBspE2lFyu5WkHwbRxBR+nlHxQWPrNA2RZKumZ9UwagHFPqwMg7GDnBPNHewmTTDeMaL
RiIE+rbW4zbqJd/ko4WycF2eKeC7Qd5WRrcmrBTqJhWjfUlQmp7qHiybZhscXUithu9ByJbwpvwT
6rZNisEx3yRSHwHY0Ojk9K4v+A07aSUEro0AZKBSwSdamQt1qUTyf7wq6dcYbynU4uErYxwLn0le
JZ3pboCyBh48yEq3zITvQfP1KLG+2bAajnWsvs31UCXmK6mbDCkwPKAm3TCRwAhbF0Em11LVgme8
la9PcwzdnNnjzrK38uezyQPxK2FlMnukcH+UXrBTEt33n9KDV1/aEl/ng4FNsClyHCv0ZU+7gxu9
HO4Vuy2M3PwBJ6T4i99D30w1mrOOOIEolLSEdpaL0r6m9Bz7YonryIscz0MHlYwQNIWCaFU3fqlK
+1INaRtaYV4B1awfHrvd3yjHMUKqQKalOcO0Tur4FwC4W8GxSmsC9X6FnEsFUiORLj6ofIUEy5gK
Qohj9yZF9qmqxvb23qBDyuqDGARmzcugEtADXDOVWV/YLmVHRG5Pym3r7AXcqJZren+ibR54oiRB
4eYuuI4UulyXeUwFJsryjOby96HYSCCxlaXuhyIfVMTepMFmdAD8UwBAPtNm3obmu5+5hoqPHo26
+F1LSjV9NY8oiDLnPO4X/gnHpXshP9xlbnWcupSqcWEkg5h2hPM812BySQP+6urcT1T9srcRoQR4
MgB6w1xyjcPw+9HENWn2Q7ef0kVlLymyekogH7VNTV24K2zZylPFgCA3qKtU/iTKS5cPSoUK1MKK
1MRWfhPuznPsGMqO9sjc5k11U33MtVoQG3pDaPzv6YVKPwp57emDsLxm5BjNhBSrnjkWFmHwjX/a
x5zYPhlWfXqbRK3nx/m46Y8pD/o5jU9xsf5BBYVtkTRMsW7JTjL5CB7yKt7S12XkSG3/K/ziVYah
cl1snIRk8DtjkA7dwtHRmbvKg97AJvwk6jttqrP9wabRS1iK4tWWuOWkVC3FUnSuBQkShgj5vHBe
bWNGH5UkudZFvNop6fogBlOIADVG4f7UUZOu/Z6WX+TSNDCcPhDk26F2lfljnxmSWJD0ydCu1Ca9
zi5GDSkbbZ/HycC7EFILvJeoAvMnEwT3cTpLXgshtAframLrlv7Y5+S17aRGsWYDhHH+hNoZyrA/
vE60MG1d28QWzcS8grZgTHmyiLc3Ygu/Np6PPXCMCAgNYLjPtbHF/saLSLwBf7ET1CQ0EUAyZFC3
3ao0ktmwmNoF6zpmJZfK9AJqLh29Ukpd6cXhtIhDObVs2iHZ8QsJi1wCyYGk+AID/0PbhYWuawJn
d7y7AU2c5a475XQdtM6REN9993tpubpb3QOgw9gdUVH6Mw1GRzXK6YeQWYy5lgSsiJWeLP5Ye9eb
PS6p3bUmLVWZ80p02bdo0DgC7uFpk6DBW4hXHst7kjMX/QINVi7OlmYhMYwmX1HygUIqRvifmDMN
zIJ3Gg/C+48pciALqDrnteAkjkwkMRiOTxMOrXkYWilVDhEjRSXV+c1E3PullkUE0JtOnP26gGFn
9UzFwC5t3oO6SfQ6KOMWUpRluukykSf03N2vst11jICiNP1FsGCAaRzHHQ0dqL+xCSr7wvN0j25h
QNB/Ka/95omNrKJOMtzebEAb/OaAnnLltu7yFdejNvb/Wlj6siT2JoSGSFI4aB4LOCpO/qnQ5Wj0
2RVb8/iUcWaAcw5vJf0A5g/zyizneONL7yEagwuxCFK8DstDje8WTZUVe9s8ijIpMFepAg4BAK2X
eZABmVNcAm70A/CEONlb1O+uE88Hq5HQYignix8+K4N12vO6Fa1R3aD3WFbQFGNe7sv+wkHivewA
VbNbQzML0aGu1SeQBYl+Rtue+KhdiBOirk7XcFzjbElhgEYFCk+NOSEusaK0diIUWeRruPRxrv2o
P+5Aqu1qUBQ5/u0riGS11gaWKIC9WxOkCa1IlC7xTrQXoGq+zsTFiC4GrD7VJPVgzsUDRmRtHVLv
k+IAVWIuhbixRbDakRaxTrmo5v6JP5LJETh4rzTc5lBk5oC2lE9IXMLcKe5wkSXtdWxhIy3eO8l1
mv9hHFh1fSFQ4JOtphM/aEsGIacMFh0MUe8ch6MxWZ0dnXY5+ZzQoZNAgdmWQ7CgVTWxeC7CwhNP
thEXfeWajzwjzv3JPtZqFJ9iHUMjPflaFTzDVpBN/Bty8DB3h0+xsuCskZfGpp2UCU+0bRHceXSb
vhWGH2QyZlNfnYF+n2ZpJXJ8/73nlw1UT+i7PVORe9QDzbYRABlGKzK6Y3MFLAxvpeF2VvsjyVg3
hxfsXW2g4TBS4idgeDyakgsovAWhne/mw4AlXv7ieYjL541w4fEY0F88lcU+CbW8wbsnGmCAKDlP
f1eCdL29PqJorNbDQaY2YgHVx4zB4NlNXwE5A3qBgOtT1RU+gj1Ytpc+SkS3qJPW75wGlGkrVdTU
rJcvwWwJvBaODhK6QZ8O1ZPDCSI7NALaiAJ+lxj+qeDEg3uIf5GeK8Ol//5x3MQqinP0mt1Hoxp7
6ElTO6uUpjozdxxrnwRICANBQDPNFPL5WAOxZ4wMMzkWK5mglu9NhyzOO1NoL0bTr6uZdQA1/FjB
DGp3snYJe3jDT2iw+/7xG4aMqA+BNRD8hlQ/dqxKAE3FZYy29eCtx3qHJMFgG8zJie9frqAKXDHT
JpZUujFYeFMPv/KwG+usg94Jt4tMtDNSfrcWr9az6Vk4UoBd85H5HjCfPL/+q045niQ7NRLE7aAz
LGefjnov3MZok429RMHT7Fay7Ng880KvWrJtfQmA2k7+v0sASGiMfGi1OqpRg0nOfJDYHgm8iI7u
XOfCe1Xn9snsf2i6gEbYvTZkO7kBAkdYXx6NjP8OclPcrFYMadvnjpuJklGG2cLQsOQAKK+wFrnM
+4MuMt5DPehVt9hGbVuq0wF9ekww8yh7W1r0Fe6pa6tjk1Y+P/DhUn4zrNzkRYo9CXLKMwz4B5cS
xXZOUbHcq3HJ/TRSZ/tbzI64bF9pIbVVbgHBJC/+5vIyH42Uf5tN/t7gbsXIRggOvm7SouxS5coO
csX9IbvEDNM/EXpy/kL7l6nmlRpf2kJ0aBoeEtqorEo4eacejMZhK+T1WmKe27TCmQto3J5V5Osw
kBu/27s2dfVTrPxv7sPO4HoAfwOb4mKZXcnd95lIcOTOu3cZB5gZMi5ff+gpKKEKCnfq8OCE7Lkw
SWK6Vj4bMK3R7uFrWxhZOCyIlgUVs1LoS4XpW7tM6eawmeOAfiCRnXSzAXkF3tPybU3SQ0rNwAyu
GV6o0TCynBTu8RvLSqpvp2BFvM/1HQ6w/q2KYdVKZGZpbsdmofmJ7iKj6gz4P9k7IbWuAduSBOTG
SRL4HO5RuRfqCnyNSKe9Nuk/esESU87d0OzgC4efjayyN70598w9jqZNG9mnEtBOpHNOJ6ycubDJ
48NmvIN4a22jgHam4LcyrcqVxDhR0K7d0/cxgterGVPHRuha65jP8jpKBw23KFmcFj/1MjnNl2Wi
LjaRiGsdUhlevT9hq9tVXRz/gSJsp03h97s0ftBxPd7ahH2v9eFrWawpnKNbv2pCNZy5b9jtUoht
qofzseVujqWjGSgDhkjbWQQYRbeSsolD+UvIBYq8SjLzqRIln4Tc/TUAvLL9YwlqLh9eaT+LTzHR
NbW8vRnkrT6qan9GNK2YtjxQgWCLdZdrGGtbpbbDuLtq/TF7Wr0NUK+HfOo//u5PT0dGkZVB/2RP
A87/XRLnQqHzvc6jsxS4CocsfcsYwtEjXZK3rLoBcgWEWZ+1tS4KYJbsEIT+lPu4SFst52t7l1LT
Gy0mfHniPtEUtuF1WPlIB6nmmpCqvUvb0Ak9KBxXEluLXuODZ9N7zr1vlgFsden19i+SHe7PgJeQ
N87PL93vb4p9ftlr85WrjSk/S9eWUifGmeJnbTjsrokG7OC+EeO1Xy1WQmFAhMUZ/komODQ0pZ5a
M+FVR+sGWl5HE4lggwv3heEoH5OpQ5EIosak46KQ8kSQYk0YjnsP7Vodp1kx2N0wRDUXJ2lwSpLP
r5yubiV+jxBNypAYNr/2/hHe2/MQKbYfRw6bCqYd58kbKWmEGp2GkHmZeUINF2h2dSCsHHzy+jxR
33GivZG8/JdW+EhVR88HoJSx2hqOlIYC50NB7mkv3giKpx9Qk8G1yRd0WdVgbnQwZi6fF1UZV5F0
QDfz8iS0MOLOuNf8RG6wBZCaSdbcyUifHdQCIGYc0+s+KVAQQ1IeNeMJZ3Li0cqky5icsjh1Q4IW
7HDWpFFWUPTlc5c1qZQCRXEQEkIUk8q+ClWsCUq+1SGEXAPspJn+ONwKUkqmqXB1+F9LnqPCRHzw
ujwEBkDXTI8zXVuhUVBmi9ZAUMQj2koRhlvTgyZ0NXgpUB7H1YY5S1H7drrGgeozTw1mtJPm130J
W/GG/EmEeKdCylL3siLnTi/7JTM1SYiIhlO12sTyjI5GJbEYX48LSU2CrKXuTLVpiQ9YgYjvE3JO
HHEVQPA+qg6R3lpZ5Xr/2/JCnq9Vh1ok0jzU5F7JlLJPz5JwWUMmJ8ZH744BcW77gn0JcL8I53Xe
vl1GqJSpiKAq55aVAGaJzPw/NAYIXwkYWoO+eyYgRmiYiDWOTYP7am+qsF8X0Zd/+nIWmPssB6KH
jaCNAgraGkuIOcGOMMk56qhTGmp+ywy1oiTF/4pIXuLAXvYvFXC5VA7LUE4FGVaUoUts607wiLIF
PELs7WzxOo1qr6YuiKMBO/QZV6KEI/7vuT13oBMbUDOl/uoWOot30vy7BPO1MQXXOLomefK/ZTGi
fFaU3Hr1p8gXTrUHlKQC2ZaUbQKMIhkSloMBT25ijZn8gp+Fr38hiGH9MEKu4DMgt/VghUc+KO+Z
FqOcj6ztbMYqjx1nWeEdElXUNh1jjgp3nXaTWmfWDZczHPJCcIsUbu7RGJmSuEMJwV89oPlhBGSd
zlEiXOhxiqz+ZuPAz7KpCdYLmeX8DQ9XYtueN/8hzYmzMF/z2HnyFpsAaxTvRv/oL+5HBg0V0bkp
v/ovdDfrvJo3Fv2UrIKF8HdouwC/PUbV/xQM6mvOEXa0t3La8bi/2X/fIbn9naEffz+88GSYQe7e
3acAtqEZaCOUDkmSWjrQfvVhw7AUng0tERlphxcSNGoz5yqavNDJ80UIHnaMQL0ahn1N/iKdbIp7
O8Hh30ae2BhK1WLuzHdWVclCUu+rH5kuPRHu8Ix3LZ1d/bAMQ4D2cabjomPziQD1uOmrNJmOXUdu
0Rkkv+L5gtRMkMs0ozFiJWe4JV90PUausgwor/FCcliXhwn5GHJK8lFYIFi0U2841vBDPJhJJD/u
zrAAoGUnkgbeRS9WKjHhtpnqm1MIA787nrAxH8IzzL9ipSWgP+z/sAg2FwOrvMNVZ3RhzleaRYfC
WA1c+NTmFMaxs8Fu9INFCrEvhxEdEoY04AYZB/4nahs60pW99k/a7B2WYSkPwHmNXNn2JlF+Cj0r
KUJdm02RxpGMJ4nsWzAThWRtFRz2Su/Xyc6/i2zSECoEe3XGFTJ8XGR5oyd0bx1uJYy5laZHSudk
LFhVLGHS6dTEZkSM6+fYvjq5lEmk96zNxhewug+yphmGE3+VxO1/cBCuxOiT3ai5gIV8BC1HrMOo
Nx2Po53Psg8ckNy31+us0k/r5mejkfUGJbT96n3D2JUE115J5oID/SAexN3h+S2iab0fDMZlXoDb
4HSK/QI+h4grn/kPwLFMCfI66I6Qo8167CgaCZ6RR68P3KtMOy5j/8aJIarpSFp4RU+Gp5iDt79o
a3/dSHRRP0D0RUsAwyv7T2XI7RKMtyQ1JWQdwvzWcWuJDNqPbjQVHnWjQu1JrZtY62fMoE+hxneG
BG5NiEwOkmmPBze56eh5DFY69iG9qav7ZAXGu7uy0rt1ij2hzo8IY2nOcVu5w13xQnoi+2FVEJ1r
QbqDBGM9k0YvDeJITV1rmtslZELRTZA2hjoJ9HR+MYUlVv0/PigQZziyOE9YLFA+4qX09TUjcHqi
z+wMXFHbZKwvBqXzfpWH//XrMQoNPEFRe2g5se+h7tzzV1k8YOi9Hakzx3ECtWfuc1YS8YqIK9Gd
COlse2xH/mwH4kzCK7tnl2d/GSuurynExmo2c9hmvGf5FYMi11/G5uE3rMaEiv25fVVK3sw6NOWp
EjCuyYhhL1xwJN7+Pg8vA18+Kx1vAd9px1TCRxvWMAVFD77XjWE1bH0BAFxXFufXCXISzS5QL/Sd
fURF9uLL9JNt3Yj44GAm0GZx8XiQpEPiul8YcZocg59mHJxPJQnXxGW5TAiFw1HDTjKRnZV52+2Y
2QSspWBUJ0e/SDOO9cSKDLO0IFV1GYjegYAq7n7YjZ0/g+4Zl7na5Xj4SGpMEWyeMp9/vyU1xqH1
G6xeZqR+2F0OYPsr+RxsH/YOHvzZba7S0jxTKOzbPfApTSyv1IWcfmEliHE+qkY2qs75LgHkC3oj
YH3smWSu3bChjI/PmjJL4b5+GIkaqsm+5/Cc9NmdsUsR1fM7CoQ6YbLb9Kk1Y88IT3IB3edZDgXN
M1icu+rJf2Bt/wU5MvBc1wAnEUeXEVW/lrVBytwYV1unLgJHAaWsRkBY/DDBZ6AFZZKhu4fWvR3S
IfKD8TyG4QqPzYqYjwzYBqZ7OGmKHxWMAZRc5+Ewpk7Vevs76EGi/10N+MEKVT5dP+pNX73GxgD3
U4SXhhGzu5Nb/tCMPolvcaK62KgVq3FC27rpKgNsjbB8CO9j5OWBBws2nEBPEkRNBk59iDsBLL8L
Zzp4CjZbSgv3nIOJsVLmyCeLdC7pLOBW6uLBhxJg5RNZnu9RsKN6Ap+M8zLKS4zL4IvAsd/W5zyQ
ztDKnvHpz7hsJTdUvWu5uuxDbG7KZtLptEzHV/FPpgAYuLWbI46pXnOKqYUWSDkp9nZCfTOAo+gK
IkmeloIbYs1ZJ18Re0pMW2GUdpxrVNmpC26psrhaGEke+91N2gm4OEiOjYOg6mh3CgiyXpac6NN1
OSgpewj6CuCwls2N9K45hpCzn54/y7kn8Tni6d9JWaa1OYdHahF7hENIAyMrA+fCIULI9DLZCwFc
I27s3svtxvldwDXWjcIAlUS8sBu48TCzbVaoKA+tkWoFxrnUTJawZZCWb92qkK/vank5vZcQRewl
Miy6+nRKpmULDS5PRbL4me3Hj7t0JiiWqRsWQhvTGIsRgJG5IGu6v7fYI9Aldw3tbxKhnhtjeW25
QSZ4Dtn017V5HUxEhBCLXbTpuz1B+y+H63cXCsg19wMCOD4EusoDAByL5EuZI1ynEnSdjctbPsJ0
4EAi5G9GYs/5ymO/kngRqt4fLISUKr7yV67Va5c+e57X3lF2G8M4Nlt49QW1k9ziyz714kTw9JQJ
eT28vZZFn5hlBmzA3v3qOx/HCc9tOuGAb/CV9ocezz7Fya5egj/ru12KCrmHIlLSN01LZBsHL4ZY
/9X8Xj/+oiZGnPbgq8t3CTky4YSlBBG9f7HrfNcEII2TXud7OvnqcoVZTRwEVJ0eReavCuJJK7Bq
n99g/H2qMu5QWVU8dMyeo0oCkMljr48GCDsONYWEMryb4T3ZCgyQNEn+1j/eNO1XVhYZNR7VaW95
tmpFdD3JFa/UECMcSLtVGggQ8BE91aFnBICTyreuAA/Vum2GcNyNKaduOVtTw9uRnyUpp5sgh0jA
Ky7bUlavDVypWnoR47suwaUPOyGS+hlwRKtE6IVu+XrYNnC9rm0N8ElPCClFPSI79kzN/1JThnyS
Oq1ZuiiIz+q+QkwFqkiW+OtnCAuXKYdv/G6g9A+ngM6eTPX4kwjumCi6e6RLyrKRaDYuqEjZrNnA
pDg0ZB5LwlDx7JX4Nr2yLym2rikzMN+vyS9pswyE3FUEXK0kQjANi5LhuVSPXgvo68v+LYEnJHXJ
iQz2sQvusCuXN6qbUdNr6Oj3JHgS3Bfq/cYkUSPNCieY7pPX5lpx9IRMmgmEEVK5N6PZdQJsz/Zf
KGrn5GdAhH+ScxpCOip2+CrR10RMCVQkSLgbQPVtpvbN/B9ajL43MMSHBKiqyOmu2VjceJPNSznw
dJOAQ3ZCAaRkT2yfqnsrax1Yq6vlegTmpD6eV3f+cUfRYm3H3AW/SpMN1sjc3fCosDU1xgZFRYV2
BCmanclgzkvF/pE2LGWAqqnjzX24gZxz1pwsoQJB1xyUuBdOzVaQ+Zlw4dzrvQyyob1j5K6JCIYp
CzRGJo6ldHCOUGgF53WU8kt1aS6ddGaswbzMQrhGNla2tYXGgWUfM50oNB2jMyGab68ukrIcax+l
QUnBOxQtC0VT3TF3IucWs+QJ6qzZAbvammE7AkYssRJvqtiiukNFc4dz0zsFqQwhTZMuP+SgMxty
/bnzfpApV9c/ac6NS+8uTG5KeDkebzBUzKDLK/znTa2OOghY0YCVXtJalIFnl+ntVx5w+X7se4va
yq3jhGkRvNBQ6YSyU9tP0V0LAEkoqXofyOqISNr5EA1JV1QQK6S1ew5HDi7xpFGsSaGA/l4jTlG+
VAzuHPCFbdhc1VtE58vqWal5FqdfKEYHnNuAO+rANQ/OjftEZTUKtXvnJjzEE/sl9z8NshuVILcU
LNBNeIc5ro+GeznTYV1gVwsV2Q3AL4rNSezov3RHLN8AiftEIPBC0RsIbBF/YI+KP1x7sAwj7HXc
Ffffg4uL8TEzXvb+U6LAWfbeL704kWwCFz5FUpsoAPVlJYgpT0Fqv9smnsFo5LAVB7g/SUqQbUHG
PVySlxqunZbfentOQhhtgGBGWyzstX7r7ngfJHp8aNj7B3rzLkioOdAL84x1Amz5kn59q+X2CkA5
2d6ze1gOVfmIMt5DXD+JmxXw4uGjAjBq4xHP4Yppga/cqGag8A1l6Flrarb9v5vSqDBf8bIkBPqS
IT+TYNODVv93SN23Rctm8QdtmWZkEk/27O5lumCItc/kTpB8ViqM+zXbi00sRSnsjmDY1vK4kI+K
jWvyi0NZdniWVXKJCewiNZ7DUawn38qHmlfR72MfrtztSrr6S81QS7MH8ub0l6VLc7IYVFy9iWSg
C5Z2YaxbhLWpgw5+1yBIs1IQlPZi8LQTK96ZRhROPPiOlPWTZJ9zUl3RsxDg66NHVaa55N+erO7H
e6MtsohSpPjwjCdEtJmPoWfyhXw+yCBY+W5WbcAq7V3hqD5ZdmBapIEaTY/bmS8Y/5J+UGBwKVz6
3qYq312bSN6dEw5ObCqOFfL9jGslioWCxziR3Gc3mA4AIsM1mNLJX5TKXpw1UkNxjyelG0A/FF8I
F4bk8OHsxmGqfZzkRgckYZ0WkYst6o7wDcFQGPGW9Jb+hxbr71EcGSokXW5Ci1U/GBo4BjmvfE7L
mf8P1pMioLGe9zuEEO4iUoJOtf1LpBdXXrY35WCctw3TQAKEDLmYL0tpTMTzMxEjxLjfx7nctwx4
aoifOzRlYHH3/O1C6kR8KB2ERsmm751A4U4RiwGI1AOPUUSOHVvvhLeYVF9KjAXlb4D6Na4GsZ1a
vB4Wo23n8aV+qyqlKTVX9X/dGW/uUl6fxUzxCll5Pvn3VfzZ2I2dsHdsLMcmD7kPeAbCZoJeDl8+
N9Xt+Fisrl5/55KKn05FN7RWg13h0a8xomXaCiVqPFYpDdPUMRTcAauoyLnzcifcFkjMcWQGyirI
ZgnnjtS5UHDanZWEBoD5KairKNS1UuRec9Mw93YGdVcM3/3RyuBH6nQKiKW239HW07HRlpia65v2
DVBK55zJarG3xCwFZEMuddoAillxmnDjXziHt7RHQvTr2WdSnkqGTh+sM9fDbknzxodLB/pb0F6I
RJiZaTNDl+VeBOmVGVU/JmkXmvnDApLSpRmDSKpJEc6tL/BfAJ1apEYb4ZRgHndXEvFj3qZFjPBm
iii3EJTIrwpVJ4F0WMDOtG5tq+3btCGPL2CIHH8Uk+oCchWM3OH5ZNOPqqv5vf6Mts1Ed5FBt0rw
v3RMlyCiNyHPP6FJYb+HdWHRt0xKu5yfj6MViSMLNpZ48zxqw3vzHp6lhn7SgOkQR/ej3vfobfeC
oRthcu9eH2W1QilZDzkJQV8sbBahP0JpXQ6kzkISWmN8sCnmUSmx/W+JDrBGGmQdxg1n+Y9lqagA
a7pvBSdEXtydPbVbcCW1Gl0GOa9NwYuMLxRnhR/v9ouec0uHi13ZdCJFo8SDG0K7W7rUMik1SEo7
G9hboXzBnuKU2DJi3/yiwvdoqCWv8yFK51zq2Mf/wivnPFuhnOu+JC14e5bgfHyNlL9s4BhKJy8K
Edc5f5+iwKeS/CM8o0le2bW8g88g620UkecbnQJsD0ZDIOyHcFHU3T9lfrBXemAdNpVia9Iqc4zc
4/qM/I42gABuWzOXtSnm7ygIjtm6Wz11woAT+4zV+j6jM4r/cPNQuCqOf4+ohkHZnFEijLOw3Cfa
8waKeuT1xZq0Mok4cTFOdFZWjBxDXyvvrx1FumVES6AYCGxbtFA3+WnPQ0s703pJia+XM8PhwYoU
AlsusY26snJ/CrbQ3LsvFWhNrvNyXSSEUD9L8uDBSEsobw1A9CDV7MBjQAGWWp1M3HBTtLnFNXf0
n3CBQZ8IEwORwLgrkXfeAEQymg9hr4KdXvZYW+YOv3TQa3V8A/L2lhV9qe6sHaejv/BFHWAdPmrv
TXMLVfj91ilRWM44Y3ZiAZeGeHikOTCmJC/m4OikAvaE0Ak2gANqXb1WSSdO2yuzSDUEcAZyGsfU
7opy12C8ON+oYjMserM+V/LKpP48nLDXCEQIia1ZoeOMiqZu3naTPlHoi2Nh1Nx7vjpYsVJuvgKW
S2pWbXaqditUrpQj/OVVz58cU6YXMqZ1dUHbYcObbFRIffGk/XencIeGEVJ0DIr14nLji3Rjh0aj
/HN2Hi2+b3MCZHT6N96tuvf0s1JxYknNzEXhyQEfHsBy+YaQzeMcDbt3hmeZx3KlD+JHLAfPrGiq
RqF/L+pdnA8z1ql6JtE/GM42NHiN85xpR5fNqQhUdFBxolRRm4Xb2TkChESlAozDaJE7rvDYbdmZ
XM+DT0Tj1gIRd5DJkbmB6ydcn4WHii3lQy/xonyCpUKtOeIVGbzDfghqlbe1LZmDEVAPjcG06Axm
MeRDE+0gnt3yhKIQdOwIxb/Hq+XoQc3vv8snJ5S0PqKkApe8GmmsOOQDTXY0Bmn7Nodl2xvoCuIz
Tg8h24+bvvM1OcDgYVexn84UuHjl3W4/93hR5Lqgw9QqJu49IlbToz9l7FMLKYN9UhzcvMxtwh6E
wlC8w/Q4poj93gGfTMyo8X4AwGv9VG3DEvf8yClm4xpYgplqeN4jGlJubu6e9puPqL8RV2tZ0Qsl
fyUb6f6+py3ntSsGokEFPpLAvCL2LJiECSaSqxQcrWFB7NAr3HzPpVwEY60KrbOv3z7E5pMZTRQv
3LP0SqreJjNB0POyhUOANnrYrBZQ83pcJqFzbf+i0HdtFr96ZcdrfuzzUBmVSZrlPpHNG+R3NVej
+pH75bP7qvQLbgcVWO8vDKufs4Qg/M9ofkB4e7ehLAXRek05pZCDvb1MIO3RWdvf5oYRAzFubSRo
AOgpGIMjZ2la+GPHtRSHQrRqyJtRykOKndjv6RLUY06fTZ6jWM8wsp6TGgVvXoqixUbgl2o7zp4f
Q60GMs2JKdH2ashVDb1H701GQg7XFbz3h11+PirZsDv4dM4dvjy8DnnPP72Wc/+WCmsyA1MV8/Nd
6YRteD+j9Xv3HGgkoI5nfz6rJjT3d53yf/1cJkQG5L+zs4dvg6sRqb2ahJX0HxAQrWG5ht7X71UE
oQ3t3404yFvf2l3Uzl8JRNxfWbDveMqMJ+0YS5Ks/e/NKe+z9Z7AQxBO/suVuWfQhmVaedwXKeBD
MfoOLsCAKs8Uz++jYcw2D7vipHqg2yDvGOUU7OikczYgpCqrH4sKJNc6R3pcx5dTPvfvTTcIp4Fc
njR0PiNMmHvxh7uGXGoJVxZfnomYxC40mKpbhWvAwNd2/USwsQwmt0eyxiICX+Y6mc8fI/aMqyYW
ng495LHs0e7sfrLMPueWVu0JEjfztD7hS5YbZ0/z8lC6E5EfyadVlLIW2UmHLjHYns9ZHPVEIiVW
DBcBN0Rs2KQXae8FIQVW78s3YB5YWEQ3z9ec3uX/ie1AvwM1SYxC8VWbFWFzYZl9DhzZ/PcT7J62
aAgJUXORdtoDUmO03NiD4tO1P/WrA8bEYF74ESF8i0N5liEREm52wR15CP5/G08WlwaeKOAeIoqd
O6DXtUqNkm07B9si+IjPvZkQbFJyn4ZVKZvcQirYWQ/TNP56YUtOpdt2nCASDjM90OOExOBW+DaR
8k9rdaS8YROLXY/eHw6TgLroYdMI4fdvEoCSiMR3eOtJjqn3hGW/haHgyELYNvmwnd+uCzZ3Pgw6
0V7i4hkhbyGjC4AQcm8fO5HSGS+3WN6yUF/6UvElbCDOpIamnDvREvqE3FSAim+C3fb3eRkSab/l
pBEtw6yzUoMUGF+PagLlBFIrnwUOKTM0L8L6OwAhEBf0GTz1m1TWM+snN+ijRy2GU3XOBHjdq77v
P8FwtLYS6HUuz4Po9jno5ZzHqR4+ZRjB3ES+DYIj/SVB9NEKE6J4R3/tZFpfnML65Hg5RQ3tQXOA
kQ+tBAfvBqCajw2YKzLQ75MTtwXpkTPJDf6Tf6IDzDoR2Xw2fec789sIH7koVdTWR+P/L/ddItwQ
ENmRmwMlVKhrqzFFKaQqrwCfWyN6x6iGfFn3EnlcQ2OD9Z16FokN7r861KwVWzvxiIthKaPlTIRz
29ISTFrlX3+SyqLtOrOAGHHuWW4AZpoSwBVCuMVe4ugP1C/x6yHzCtFkB8wbqYCRwhOlBaCDQ/Uy
pBqrflB/e2ofjRKTwi3OQUouW3Axl8xibnPDho8V0/JibnS9G89L1PxrfWJUdHQadQG2CzBXWbL8
GLmmwRyNv2uFx60ZjV77PmYSpt6Hqn+dsXXKbRF2k8bgk7BZvGxC2iX92ScE3ueYnIfYTPlxoPAr
IZi12moWBBcxTrZjcbtNWCxR7wFFd8pEjS+eY2WJ1gtwgItjXF/DRM/7lv6GUG+tD5zwuZU3ihkZ
qcybe0lgXszlXXDPIMg8/RbjA1eaxDt126HSZlaQOc3Fxbv4HeRSUhwbqRKnmy3hurWA4KMMb/RK
AzW1c+w1tpqqlfuM/rVqFG7IFBh27TGlSlX32JMxg91uLtdT45c96asvdG+KOPJoMqbV3dxpnxIE
f0gY3PD15kXsC+qkRyyh9zaYSOZ8tOSE4rpetxBl81zoFN/tZzkLsBXM5V1XtTrdNxMZV5PoCt7i
ma+UxjCOFUWAYRJMFuFfGAgqATYi7p0J6Xw3CZe+BoTayYt07joH66/llvQwbEOcf0sYIq7jQUXV
LFGxn98ARAucAeL5lUMZLQsz1Q/jc9b/a97TGfymzLc8mJHYF6i1ykCnNah+f6fEEMYf0NDfPl4x
3xDSVUPTOCPgu5spCzvXUh3K29xpxZJDIPiojsBW1SeQ2qcJCApx62dgmkcGCqn5Fmru5MZyOKM/
20S02aqB45wscC1KUQ+o3IwA7kz1jnmW6/vup3WDVvWujWZfwjZYEafE/tbK6N/4+Ts4Y8YC/2Kh
VYzei8iPG/WbsOt/ZvgU8Qxd60dQddBnP03q9cfDdZBAn1993JaBMqXLMiZQjLb0Zixpx2Rb7PcJ
kBp+jUDpgnScr3omOoSC7VTPb8RUco0Ofj2JJvxxKs7gIzRMyANFiAa4XVNYEwb+X9LX4DcqdrVe
hxwYtvvFFkeCdb4h/v6PBrrLyp/AuBSn6GhjIsQX0D+DDEJ4GSmBo0PUhpuDzv+lisCNk+ieiAbZ
jaxL5JnwOG3FEs1BMvsMuLVLFdzk0Q1EpcxvHZ+3qPKamhmG3T+GB+QSXZXgg3gPhksTA4WOIdp5
JDrRontq6AviFbTCz5q1NVk+eOfN3aL3uY707U9qjHZpOI8LxE8kDZc99sFbxeuk+WjMHoNe3scl
TLg2BWrtUl1XJdUh2/EpfP7HS3ntcoWFTmc01m51vMFQuBj+I9wCORlk4iyBDA/l8vQIguoPMryP
h7udPUQp2DyyPYuxO4a7cBpvA3Vij4pSuoM2CtFxEzhl4y5R/+wfrQjakBBR4G6hYh7ZuLj0uXEV
Z9UQpypOnVsJZNAuWxfhkDhID/FtLiAmVMzGv3xoheYW7XEci9VJuR72KTBJk7smY5HRsMBxfunZ
rOceOJDfcGA8QzHMhXd5PL8qBkWMzMQGYuwOdn/rpViM3OiP2AXNbocTScmx/JtvM/29IDF//aWd
A++lQ3gTSAIkXsUJcML9AF2tzZQnvDRP0pqjMbwydH9PWUDBcV37BJRh5WUQaXFSSsWcikG4hpgS
Lo2xmt2J0zaauO8fB331M9Lsam25wyH92OFLageEfL4ObTqJL/fxsQi9Ypm6Hu2g2LI0IbmD6Ccl
4Cj9Jp36BvhkvLCx/teE+WdeOd2LUDhMw6oZVI+JN0zG89464v8kpfqpwyCJ61xsjv4+9xzF6IlK
hwjnLd/GXaD+R4PFzJf48Emi8enMXc99ciBCDK0t+wfkgluyR7cWzLPtMIdqq+wGTm2L2wOYNlYV
Oz4QdCyLWeEJ4p5LRiazE7D5N3039UX7KwRDuBn56k4dx1egBi3Zgbu0C+UBLUMQ6Y3GzgTuzUS3
p+rVGKcRJwB+Jc/+TQka2RqI8ar5pTaV8937DefQMnuuNi5+ebvSzsPjQWi0Wzlps/7FhINj6iKW
uczJdzMMPb7mqu9A6bFUjzkyA/d+Wrd/KL/M5ot6bv/nb9GrcHg7aqne+mazRbLlWoquS5CpRhyK
pfMec/laqcileF+uER2AsblvGn5ZK2FCTk+Hh56LRCa7FBGs9nfZPwlFIzAqQN+uXxmvGLK83fPn
Bke/bKqt/TbK6D2O3huBkyssaIKEtpYClw1LwR2LJeiPPCjVm/6Gv9rAUurebx3riTf4+W3IyP/i
BPjmpgFkctdmR6RZKbpgIsqgIh0gDw1uNH1zYZwI3F1gKCdSCzswHeiwVqr/n9b6qhZZnBWyFIH2
Kweh8pId+/kaZI8Ky5DWHMe9r5MNpfr9NzeSiS3W1QSSZ7NpdbEOTreWynNldQaZFwmKoGzoxqaZ
kb4QUL6oULgkg6qPC3FMtsRiLnTL0TarK7faimBsNwgTcZSMp+i27vFbp9bOyVm2S8ulRq+1u7uq
T89v+OnKvL2NMerpJLnXaPNFzOTgPfY7O8bvw/bHqWfxfdFbFV6l3ETDiwce3MCqMBLMzxgK+VVV
+ciWCQTrCgVOKp2m9uRlP7J8+VEAI2HpHnRzJnrT/Fm10UZU58rk8uy49uKw35svanPXY7PIB2Gk
m3PJIv82gaI3j8w+X080lGuUKFztucPrVtS/rjHXqI4dzpsNn3McL3ue75bQRGMSFJvZ52oQlskv
S/DjlHbmikT5NiNom7sk+jcQNOo3q+p/d0GcSbBgjv4mXNQZVdPkQ6ZgCh2RhWBTI8Etd8n/MIcr
YPaarXQxyiPRGFYO2Xrd6bqnbd7ZIW6pvQlFbseBTheGuqGF5tmxBVq7Qm8y55nFXkoTC2J3dQ+B
ild3MfvThY+Te45RBsNSHh1IoiPWs0V11W68L1u+kRDH3Ap1XZNi9j//1StHuzvZsU5k+rZP6gj+
59ffuEuHnBKjrznkZL36M+h7VDhVzWT+hSY0us13WjUZO+KiWVAED6iIlPm6GDiDatEPr1G6lbu+
EExjpZk29EvQjCj/m9Fs4/1lQfI6XOD+ZNuwLe6fw9XSBpcPeBNMZHG0L55qaS7kUVvHHQxPKsTv
RhiBJuEvt6SmvlPH3T428jn/6aOaHX7stAn4G82QUOgaNnkmbBWuznx7JF02sTAAAAlVrkRYubeo
V5DWRzg0j9U+dr9mLjX09cZVPF56FGMsDokt+553Ly9U+ikA8WeLSdqnA+bO9ex18VDJJCOc+NWt
McQyZhwvPhG95mr/jam+jDmd4ecy3dAgPzfPs6BgluGSdKiHiEpTTPNlWmp+SqUThYbX/SqbUOFR
HOWoU1jDfvSX0Llyg1IymzsACK+Vk0noAi+oas469cDO17NwBZ54xvpLTnbDSzw27NO2mB98duGA
bs/x7ZjjE9tV328ALCn5+cOGapPdSTRULlirvEZMx6GtNeDESoOUJP84amfd5W7oqDpU1RCxOjjc
ZWasEwWU6YC5vq5MBx9hyguHVir15XzHWuZxNBMMRrsk2OLI3erdoih0Mr2/IOgN16GYV9pBUQBV
hPpxRZHJXWex+dcAJo6iEWXTB5Byu4huTaKplUYsuVZBY3fHo27JGmjeZCEn/Ci6mVrReQS+XJVp
aW3DHsIcsebUAoVLRqWsXGCCwrVcYp9c/ga8vMAQH4Z1KxT6tiaZuFlg8HBpPoRvtIosaxRT3Qw8
3+A3yRQEGD5LpMj/4+AxOKSaJ3K+RnZ3IUDV44wFzBs0IqVoLCHqMSDW07DBjqFiRTp37gz+YmLO
1UGeLwWQOSbtmDF/ghiPN7yXf7wEJb5FDb+fI5aNTniomF8+j5+w3boNr1nprU4jctjwfrlZKDxr
wtehvDtQRFI9X7OR8GV5Q9Itwl/tFereuSV2aKA7AGjcibvgvddi5JNpRzNnvopD3vjGI+x3Zyd1
zQjYfnnWS+82PSFqfqmlLNM2vq4yKomAhMerMb4gfKBBfAXp9BtA8wjc+OcRCrSQzyvnRofhtLRr
XE/KE7s2vPmoDqqbiTs7hbf95kJi5y2aA38StX6demFzCrufM8XMj/jqguWP8xepsvZ2BB4V1e12
sbU/YixRH0qF1ZcydoE3iX4XMJExqmQwWxQ9WCDlTJTPycum6v1QnedJ8NwN+jnqUbwSDXprTpD5
j7YiC4uAcXFi4u2wM8QXMJE2ItwnU/502dLiwgdfbUx6u/kbb2/1CPmwcsdnVRnbcSqg2H6ty/eE
apxHjKckzcikwkpwWHg+bQ8IAGXrm9axaym6nEpchJHi1oZJPb38njTduTMsH/VwautPVabkX+V/
UTRKioShnbWOTLuNVTDV6DCHpY+y4S964XvSrmUaXfhQFGqiIIdEfHSSbjs83uP58udtXssvxAA6
W245hLgQHbzUadlOY2se6Prxc81/i6ZpqZSS5l6AqIVWnS8Peqt4gmlVhk+UE516f2+bbGQuIvkN
oDmPCRXKv6dpdq59swwYbnDG68lpXpGtUzxxQA2cEqejKuC3IxpK0NpmaJAfB12v+CQ1XyIms7vy
q0mmXHiJtEHW30hUOuP50BgmiX3+ZdiN7fLIJz2NatLJDorRtNe5pgWEY0XKYTcgTk9Duc1BzFCC
qReB9cqNjesGIwjx50rYi2MGIGDfjFOAogq3VVxdMEX2AVs43yIk8oc/dz/4D2j7vAXJx1aO/D6c
7mqY0JQckeGR59Xlr9d+HM+a4SfXsKHuY62SvLgpTZaImP0SAAYZZZNTQtUxH/wb+V1BLqz2JCSO
VrAvF2yAsv7QMDRs11R9E7/CDou0mgyR57EgVgZ3pNkGBxeggbB28Fnfaa7+N0KYmB2DIoMbtSvu
kqNGsRHCRNcAXbqPJLNcSkrUjrL1ngHusmDDHEl+dLOdHL92+cQ18fEdQaJFsayjCSGnp1G5anZ+
uqczkEJGOzXnTzsxL5geFfw/DLviDXMuJCiO39SOt31S1Na7xfXYhMer+p4DuxQmjmB5RUEKiKe9
lovZRj1Y2iRb80iRYRiKtcTfnszgHmFGcNkiyrfEFw7EZDQHUu+APeKfFRdeuAVT7VowWuX59fuX
0fR6fp20hHhCSsj6/OViNoIMiszpn7Jek7tyUWAWhi8QZZptbl8JeOG0mzbkg17ZrVKr6HWjdv3t
MPSao3bNQKitzRb9b6gvIo7t6e3TsGROaRDU+APMJpGVjLVrUYDid8TDeTAl47odmTINxp3Ewwfg
BQ5mCVGzQ446INpJLTBTFpf2InJS7KgMxJII3p14GFDvAh2SBA5uEuvwTKVR0H3dgBraoBM4FwAb
NKSSJGiuEUyPt2sSPJ2ETN/npvvcZmF0dN0gVA8N+KIolwVbFYozRELiaVzoN/P1I408q+7lz/5q
9fAORk1FoGeDMtaYjKcN30jyXCyekKMWe7cD/g1svvqco1G6vKWkGCBpr6tLwE7+3BXBlVMaCfIe
Ddz6ZhslEDQOC474o4hPQdOgjB0c7feUkoki3UiOoRgwWDMiUsgicZcRvrUqnOtiqfkO97j9/qsS
noXTP2h1iLMxsm5h5BC/DSwZj1J3bPdl1LSu//WyhSDGrTYutsa657NT1zRkrOJpuUqxlLuVMAsR
Q+BeK1CliVyxcLpUjz7jOlWSJKsiIL/v1PKEOFXoNuIMkYtlDHahAYfj8cy4LA9EtoLzRCW3dkum
jn7a473RvRpbtNCVUe9tfoIh4kQLSuXnLasU3RpId9lpo/Yt+RhMKqujTdEjnHvrZQfq0srbVg1z
M3LT908LcTG8wzxzRS+gDI/NDkQBPWpe3J9JKHQ3Xa0NSwASfpR6CPsC88eywzISASD//50Y57R7
vzpkwS//E9ZW4Z4f02pBCmvjDT6X9brloEO/ssGpP1PtahI2GhGYPXQkc29vPccKNXg4tfPauqj6
mqftUwSGOPOxIyZLMbiosW9ca1hdwYVSnSSnrCLWTO5S4NcMhsthxzHM60xx6dxXuMICrxsFICmC
8JiQDnH7+HbHG4XydrLUthvR387AmHBzn40i35ZHVYKDXTUzHdY65TUVpALciCiknSB6aq6fhAld
qVX2y/n1sjlfAhWoxqiAClli0f5T4wp1f02ChvKTJtUDcZSk/tp551PBztOQzZzzmNPsLSTABR1n
vWX5e6CWASeOb1pkDG+MFcbtvsxiNFjDPAR2OEH+puQsnHCkDKwNXvg3wUV7bbykbyG1wYEzKM7Q
p14MYlEaxBpKvxhjcd3jjvRSXf7O7+adFYjcAh/MBNOtzqun3VdFhlIUtR1hDW2skQ6J+8sMrVY2
nxCH+8bnP4KDaIbLqI/1qZ/GiCrZHE2fb7doHfXgUC0euCGnwzlhR5G5aOosR1ULmHLgGvL/+e1K
/1fD4//KwGg+cXTOTd7CUg1pUQwj8fqniwZaQRCBZ60afr9hMEKG9EMi8KWl3lGXuFh8/c4BpneX
ZPf1ZoGjb1wYuujfLCN+KVXWOToEv7WCIRk7DQOx/HhDSbyw0Pt9OgnKoPJldA83whjrgaOmjg35
KUG8mVDF4+K+gq2BPu65oIn53Cs9sfAcFK76SNb8Lmb171HHLdSmpgSvXLn8Q3ezY/TulggTpwu0
vpyRvHk5eXsG53pEbjiV1crUJpmSyZ81OfYeNh/o7hZ6EzTvGkZEIcv3VK5gxHtoMrKKjr2pNguB
VXkHG5IpNAEyPsRcSHdOEF6hTFChTpyEsBeVWfoQD9x+T9beCOV/Aje5O3ozGH6bcJbiMRhPMY0q
+ZlbDJyelbIffqIn9oUHpj6O2nWzVXnfOpMFbqifs/2SdoSpITM3aI0K+VYh+gyPE2mc6JBXkbog
iuRBnng/Gz8alOUsoiY482z+zOq3XahiMZqHCU0lehcG5igjMb1iRvoOv1oX8arbUwIC3O0N1SdM
6e9oj3Eimn8puJh0rU+RKJzDndLhRBIodxmtavAxHNRJRrGQlZNWihPjJViE+IgNeNj1t+U5nT9z
X0nWrLgLwGGziSFeoW29NLi+bU2rCLLQ2cNgzZjFS40xnuAYyerFr962hAfVCrfy1osfUUwGiJgr
3Wan72qxSJZeAsITBjhXzUCdmomGgb1uKAkpdcTRpOF4b1Oa/2ozAppi7Fknbt76XUNYKhJyXnyJ
f3SRc8NM3eIC7fJZfdwspKesCR4VNd0xwn2Eb8uvPyafBTDb/GV89iYzpXps2Iox1NNs6VMeOXKD
VUYTR73tsC8Dn7jjcaiSf11TOU2wbCTn00hGQInAMsS6vPfgwKP8zoMnIYMxsuNv/ZE6TbFRGHgg
PfhgL8qUaSmNuzIjj7OnKdFcyCBxF0aC/5J1+A3/tNkxMPSHF9Grn+YG2zdmbtfxbbhohabnRfX1
l+2LL7Q/9aoffYSaZfnuRdLu+ExcpWhjMwtN2/jba2Rk3How5Z9P++IpN9wctp3Lm59loLLt6XPa
W1EpCr0ZFfsmUKuhytJaYLn2ywqFt899Rly6X4G2sb3DOxJAwkF8OaUVxzyltnHT9msXIblsd1JM
T0fApz0n4ASNw5oNyK+6dmTbzcJnSQIMNITLRmV6g/PlVx74ZH/BX/GeoB8WpKMnlG9osx4R1IeR
PL/HiDA6ESg6U93LK8d+TeXjIv1g4PabNuRLCmScQjNMDTFT6Y4121pIfIbY1fGa0QJVUn88X5yK
MXIZAAS7tln9ywzl3LVdAmSFw4drkkFy91C2FJK4l9tvLs/L8Ltct/wBwHJ9+D+4drxKeHbygBSU
RnjRibSX+f/T+XUA5SYERMlpl4sDg1Lh5xboYvPjZ0Sci2oaFTImUrwAMRiyMdUWPaukRFABCECc
5UXLMu5BoUcmOCGfBnmjlvrr2V4nS8k2ONizcIhQEBfn/jhp3cSRp/H4LyRW3Vwy5rtqIETjTsU7
6GzDDeDMdHvtj5KGd5Az5rluX28iKDcyl7GiJVKxn0k9HzClgUIm4r9aPUudpQhujPn/zh1aGfC/
tzDlOQeV8n1pJbfVk96C05XVmuNXmDAdJfOcwBHwg64oanVvoqzAZKEU8sYQ7NCpNhSp6LEne0NF
lpVioh7atGG7Oq0BLAhaLmwujABFBKztj9GVUncFNvPENIC+z/DeDvBMFWVfVNRZsRHDZ5ZKySaq
bGfaKx+5Q/X34eMgoJ3i/aX1CNtEdGPxFthgtCVJmEMCCEeXf5a45HpyfzKJi3tq+RgAi304CLIf
Cx15TLhQthaaMSRY3+XvXxjPRoZsO3KQ8ig4UIanEDdRB9IhDtruMKM7sUkyQdHjlBPV6bwPzPZ6
WHUxnUdIEhDgJ/eTReRmj1M+pb1GcO+z3jU9LZM4EIwrydP1hOdK8XKNUEKWgPZffQ40dOwzNdH+
XyRbJ3MAEIxC0wA4J/O9acX8VRp/Vffd8E4v0igChwGxI1J9wgpVKC51f67EOGO+pBYFaARzw6JX
vEQ+VhiqQMpKJtSTCp36Ar0AOgpn9tf5Tjab82Y6ZZRMohmHgFTlg9hWhNChAXBWG6qEc2lleCxc
JxHQMK2kxz2AIrJ+Wl1nyYYVvZdES051fb8uVoOK7lLdG51S2mCgaaUQzccal49aS58S6+UakKOM
albAEhcE5t8Dqy0B6UgS/Aa6+njqJyYZGoDoP+Wm456KmEzVAQx6fcppYzmmXce1xDoj7Ep7cP23
7a2iFB/kC10ldIYklStKJQZ+0jHsSOeAPqUDiMPUzC1EbHvoyYTi1bKGpPQXkhz2dD6XrFylDeeK
bYd3WHzNZHtm0RkfjcY7ZgAO3OLYIJcG3ktESnuSszjYBGbXaJaHiNBj1juxk8W9x6kZhUNsJSKH
+6hvbBEBUkGinX+IkblfsRU60mSz9TjEDlGQeh3pPmlcSDAARJVu/wlMU6BVUOj/Jmgk40+aIJLd
h9AlEiBdzE973NslZuOiRsXJWEBmMnmMzYH5Y4Qz75bj644xrL1EDP/HnhUWDwXSssj9LybY1E7c
ns7ojCqvtwZZLBf+GjrAyLbQ9zOoXYIP2Obro8K5yzeZCJtkgw8wxzv/Ll9XFlxUxJCe3/KqICE6
aO9aDD04RzRvc7VOz+BAlmMNrOeOic3Xm6A8St1gbhRt110+c0ylAvjySbqJzk7y1CbJfsvDGTDW
ftxtuPzI1TnDDclKuiEnYgUKxPFFv5vr6OBzY3gkJxY/cAZpTTRvfnXJc3Vrs2JdXbeRat5ypQUl
DpbMGcPx5uPdSTp2I7+sl6+ONNhidwqgRJ1QZPBq7G6eqYnLptmTuNZ8dZA6mFpnZqwj2pKQRpbo
GMqfur3jJ950BNam3GG71knOSogDQCnyPY4n5xxStzhIa69b8+JhN2wJy/hs2zOrp9jzCSkHYQdr
543UrLRXHbeTDGGPGG0KImG9OblmEysPgpPyebmllF9ZPY70mnXDDNytFyhKe51Rlej0BsneiZFb
AMd0Bsm42C0mttvHOec8rfW8Y3A/tdxPPmf0AcJb3gKgq/1mZtLCLnHM1oshw9jSk4oXcfFV5ADQ
Is4lW8acxxxE1yfSagm01uYjDuLsNjRcwrkfZo9WvwwxUttUSfnpKcGZPzJq6RDJcAfmlovbNNkz
HsPpbnojUO8OHx5lZX8pwvJ0SJa5wGhIL3iXBIZTYUC6wup3VM9XiAezvKe2XJpiiePQM3Yw8Ve9
AMTxvlwt/v92diLaqa9C7xbCx7KYsR9TGdzHmX/BE5EF+HbEr3mn4Nh/UsgpVRoNDZqrc58d68Ls
+5hBM/mNo6ro3urVlDRx3+uAdoYGagLiWCibcysS+3wFdFQtWV+JXJOD+reZoH7x8SFVZ1ujF9Kx
3hdfUqsWMN5pyXdPYh91Zn6b/Nve+MJzrQUfO/FMIAGB7Y4LRgpYSrJXnk9nRDiroofA9RqgsQnb
e3SD9jYsm38PIggc5/rZQ7krxpa8/B8J403lG2CznexdSrHVrlQ4FSakVwzaAD29pw8TVuomAEH1
XJOnIw3y/Yq2sj1aJMdLEb+bpEC+/hVtIwjcJESDqp3W4JAeHEbYvbq7RfgMrRMzQDQqOF8bXpDx
UBjqdq5qtE3NDJBI3jmfmf6w54NWLncxA6kK2o0x/yeFseJqjOerYav0Q3/CBoWPgQGiAG6W2ik7
s7C2fX3+V1wJe4EM5TuA/kDO+8Y6JsYVUuibEh13Z3uaYLhGzI/b9I0EL2x5gKwBC+GVbF4cxlVE
QsZp8jMmdavobds5PSfjB7tlsnhfyx/aLsEG9qa5ioj8YStH3c067kB3Hp/je47H1kKFwLxFJ4+6
zG3IaqBg72rMKxvwkvqdey87HekYIbkM49vnLXzMFeQHQGFRNF6pQi43RJYhrIeYkK4j/Skd8Ngi
03xDENNLr72sibrl0aNHv5mjzsEM/vakobKcAyw2qzmSGNeUw4kwur68yFBPqyOEUUWCkA6P2Mch
liKNhoJIKZLYXMRE6sksl6XODpakMuYQOVwLi7PNJYBHQAYo2JCUCZi8wIiAq+fVbY/3nEMsApaU
pPRfS/H3J+OqIkSc3j8wH/jbsZ6cacj3srI7V2MSMfYJ8WEEfgG8GVeH7UQgcQ/zfZ9x+IO6Z8mL
J4OYZJm3iSv0+qvi6nLol96ME4FHNSPV4AC96CKbjTZTX3MYepeZIL37WBADYgCqwZDrQ/DEAtLU
zpqfAuLOiAPsfz15sBKML58aEn0BfQR2OZwZMLq/ocp29PNuqF2bhYsSkZ8Fey8a5COjLHYJqMZx
A4bS52dcZzfOodSrgDeJpP9469+l7U9Ofp0yAMcpSoVd+HZDTUvj8ICteypbU19VA82BIHG7/xsI
doUnqcsLa5b5i1etsthRG4ky8nHgTPnr2sNu+Vz8YICSxcsOHzwhcLSQsrn/IhCvVGS7UYSXtEfG
fcqwMxdIWrt4FmN3Cxn0kM8talhbrjaeH9RI0DobDf4DNVh7QISyRTtEyMf+skrXviA/Oqk5bJRw
uHexEXd2rjtO/urPQrDS3S1JFtIcO50kOqB86AO7OnkejkSNYdY+xrTmX+xy8ZF7LH/vl7J9Caim
k+wLOhtT3uMnFqxOXh1CcXb6UNzat7u/UST4kpIfg8cH7tBI3vDnatfOpemyVxWnHip1mGamV79e
cSE5L8FyNImEA4TxpoCivZATIxT4SR+JIen2LzDTM/C/xvNMub9hfgKh6qD1ySWUgvy9gcOcrYBQ
mHAQVVP0fCXCoj8XPVcWlSSCR7gB27Ngc+3cRBdGRhx38oYcD6cDLZLT16rFmye/mnswktQ8z92L
St3jz7mjMHLjhGfxOy4LJ8pZ5HIAqBnXIUaFf+iL6XUz94owMrYYbOH6elqwwecI4dqaMU9+7PwL
AEpAs874b3BV4eXPTyXRyavB2l5fOswlw0dSFAmjcGKV/hWjc8LG/RrU4dtIhHpthg9VyCTnWGoy
6CnRtBlJeAJOAyudERk8j82wR4G7pNNAaWTF0WpfAaMJIDfP6KBoD9my2SaU9Nzai01u+F5Gb5X3
ofqCe77jRSsOYKpw6drqERuME/ILH0+ZDXFfoW3mU2UUuDJgECH2tpYufXdiZXDIp6inXdxLVUdW
wg7ufMbP+LPVwk5L1B9pncO6Nqtqs1ptjF+tuTwwT0AWquptiAEJ5GkFEiHkdFGdbxJWSxIWLGTO
UQWsMhJupRB0qWce3RqEHSdx6uWL/6GEBzuOf3eEsQj4wuvnLD690WhjrgLa031UgBvMAFBPU+I+
v+Z8c1R/erxKU60+PW4j7bP2RTDDxZRYFAZjW2B30tu7movHyHtyewj4fQeB09DLNIcm5kLWXd6W
MhYcMvtKnZkpYfFzNAMaP51NFmqJiLvCe01uoWFo1DALXVygwYAqE6Hzba54MWY4KkULAI07kyr4
BGKins0I1p/Vys5b9vv9mhCP0Gc5HuX07t/QesqmBPGUNm2CLh5JDQXIzktUMCkZQHlgMWgwsPpr
aTRplfGJTODJ5IQOhjwqx7Ks6VvpZv6yFDIU8qJElRJXLlzUX3GcT52wDboE4ezdcyXO2skxpy97
jd5dhiJtisTkCdlDRpRU7/rv3OOJ5kgQtSrhotVmYIRgRW109sLXNRntgUvMPebXdpi/7eaxT+W4
/TK1fSqyL/KFZ+zOub+9GMb35/fOEvt7Acmdl79IQBCwIh0eWfiqYT5NWwFk4xBri1DHA1l0pVVH
JR7SgXOeLK8Y5465FVEKALZaHfybubYvp1TRaB71Vrd5F43ICz17pQGGlytBPokcJ9yXf8RrLs80
BW1E4W2mCsVrEDWv8dWGo8UMXJ0dXg5oo/R0HMUJPZ47wNMaiUrIMGK8YxrXeUcQeJBFTkK924Uf
m3U5GMkhnugGYRdWLFkGeGhr20z5ZY5s/7JosUdlyRKZAD2xxmc1QBJikrLYHrg+gqQJKXFFJ3eP
juOwKr42BaZ+XJn+1f89mim0R9h9VnWZVu9FqhINWyHqEpwJTbgR6JxOn3Y11/kSIX+VBbko7Fe4
tfEVx05H0R+ecQiZfgAux5xxbtdoWvBeJIXzgYkgCuUmbCZySkgbIRzgLtkyYfq97rY8aPW/TfVi
XusV5Ofzyzb5l51FxEEBZyUsEX98PX72nMmIqXZn2IBRqq0RehaBklxHv98dB7jVvdfGSarT5j2L
kW7lAZgTSu6IUAyauBGGphy+ESGldxKoWOa6GJWcHVxISkQYhgSsA977c4UPeQuMR/saKW7SGJ+Z
mg8pgnKhz3njXb+i41FspZ4KyIaoBzeIR60qPNYSh9I/F2qpoMsNqGo6tulC/LiWKDT8aOaAus0x
kcKofbkGyxpZdxwxwWmeMFda5X91DdfcDK5Si2+6MDOFtWkf3Kp0l95jgK9WmuYicKFAD9yBJzI9
OCcwrMX7Kpi/sSWHHQlYBXg95k+RazzgGog9O+Da3sH8Od6+ngOj0ot5jAVUxUicwYSn009uQDQx
nABp8Fcj5h8jZSr4rQXmSx0kX93E8rB6CBIcirouqQnXu8DQm0KMiPb5U0drYZoxIOD12J7Nbeza
DmNu48jUgvJ19g2wtq5ZjofATL8KbqHpwcDz0GBpUo2nVr+UWnR/gC7HnaHBneW0k7aRViLtXaBl
m2vpLQ/Aq1iG0k5ov7BN9U9EpSxU1COOhhN/odtapZxnzIMTAFC33Q4hxhnDlE2N49wmO7jIpNH0
sRDyAvbdMQR333IwcC9gYl4Cen4kRar69R7xwkS65aTQAT5bTndtW0DpozESueaksnFiz7qErsgm
F1KcMAYnD1JcyeBu5bu2/I+B5prHOEGd8165tZq2/fP6AfY2GaC07h251keizOH+pHvUSMI0glWw
FCstH3LKzasCL37Ak5+xC5wZSQpivFjdnEgGYJS7iHd4dSIg4EHPl+umQFZLmpG9MSDinzv7OqgU
Ss+XwW5izkXtCWKF7q8RooV4inockq3E7WFSySk/PXYFsel7WARrsimYk7MNZou8FxaRowLrGg5A
nmXB/p+WFFqpGGF7reLhQgsi/F/55Ilt7ZTpScXPRrtZT5P0phb59R3HVeFTQLLjaSUV9rIOXL1G
MU/KQGdtRQQaV8BHcTvNV0esTnckb7k1yPVesksvIunreWUbF2+LokuORrOKEKSzNC3QDTUW+HFb
Tz6rT8yJadpn1gs72GnFAnP6eiqSmSZEAorhRbKs1EOmJSgezN5x8FWooOYMPxOWMgLD1xIu8ZIH
3UqtbEHqN7588N+mxByA+Pvw2TFMP2VSIK5+/FMIPNxJ/Vh6rx6Ukl7W+Cmu/YOSeDhBzT7ZXuoN
mRQ8T/HMTEBDUA5+7W2Im789c75JDXk0Yq/fMasDOe/sNcbBHf9t6mHER3eCEYxss43Nx1RMqFPu
aNwd6pr8LSh3D4u/WrTpztG1Z9ss1FkZAAT23Dyhs6JXyBfHKOxYxgQ4m6cCrSUNg9Y6+f45naQz
GI60Oni5eaHxgTtcZgFMmWh8OSG3oUbipRLveW9Dg1Gks5+BqhKGeAA/bb/8WBC6DU60/ziEHUxY
VqAMPlTgPD83zJAFeDbhFfJPJ9MfAVpSX+Bem9CeERuo1aVAw5YU8J4tqFqVJhChTcfBMJdMKkYS
Xat8CwAtw2P9Mpppwy+/4y5q4UXy3fA76mMacAdurdJszdkZvDMRnyAHZIApY0J+m2Rr8G/pVInE
IOyMREU8GdsZ5M/gT1UinsdAHvm3k5aLE0QmhaCSgZg/QYCc0UOcy1Ck4kkxfDa7CbBbaHggukq4
u1GlzSWlvrVq1xXuqkhBa4+JVbTw4swtj5sRfci92iqZ+7ZknEtPyTCZt37lQQyUd2j0NUVKG1LP
Nv5hnmppat/8Vz6CBWChvY8yLw3gOkBFdhVy7QPZTPropcJeHaeZnBr1+dtKcOrgJ3q3lnQ2qIJ5
cw+OXBq3s163kHNfrfwRJUatNBTkDMzkmnFDAU2OVFfrdf8X0+r9bS3UryqW5ZQ+pX1w75NUP+Qa
B49JP6dZA8Bz/t3FoDY3Gxxg2hkgNUWXaf4a5o1Phcj19L8t5fXVexplMpNdSMU2EUoMmbA0JApD
0Ab7kx6sOu3erGPWYZza0KZ4GY/th2LdgLmdUfpOLSZANV/j5uVE2/t1DHfvggQYcOc3ayO6zTjh
e0720LD4cfv49mMChEmUvddHJVLpuxszBKb68bxGBIDFSQaRDt6d4ZX+ZMV09SO//Ncyczdg5C52
RNDCS3Fs47K79c44BW4megRwQdVbfdlEcoKaWsNTq7I18DFW+jQT0lDTIZG5aF0cutY8UtI5gkIQ
/v5V5ZH71ewvcjzzN0xJaR6QyLLQz3ihksa4omnN08VGKa3ad+loOqS7N6s7HzcXMd/JzSnyvS79
LAw0/TGbSHC2x+axQz/wihvv55NHrmguPXaAG4lScATwmIxD0T0Smv2iV3D96Q2fmMz4G06XeCdo
8yWpPdDtySw1v9VEHraUboeQ4d+69bLBjDho3FSO0xKKiR24Wa4SzPaNQDTs0hikGoT33Xe39ZZC
Ni/JTOq18vaqtu4+xZoc/JlB8hZl1URo3C+3V/4hxz0oVGoXKK0pAjAtAcoGmHwrk/7g9IfQwEUb
8eIlBVFDohDgdhjRFn1AlHOPdzQSHgCbGTaYefgg1jCe4qWTcdREn2eBifOcSbXddhVLNbOxJ7Xc
4NNHKnFZf+eEXqYxp1io+oBhOBb7MNcJHOQe1TPws7aV+FDlmyklkm2LSVCcnYzrO+vXarPbVHnS
S5ZZ8nSAaExlIOpW1IXRk6gUTG/eHrqSWM5dFpR6JvabJrNN2huKah2c5zyloP+Nlz+Z+sw/aWqW
w3MWSBp/tQ3BkWwpy2W2Muf5fNUIK9s5YD6R2uE7LVCUPN5InpG9mE4KZXbuKVWAFnOk+zXo2ev9
uKD8JUZu/ZcmFKZlAOcWnJkKrrqDbNa+T2OMSgohsAfyJtHIcYBopGqkZCtxo8JIb6DHQC5pruyN
04ed/C7L6cI2nYIJ77gRihUx4kX6tWdOozBS+635hRdJ7VIaaU3ynNy0q+gWilSyrPjzwJRrVGp7
S5ac06cbS3FBpegaY7AS5SVVFhGgg9592OHb/9UZT1v7w6HPTT8s3OVybL+X/DOpWTHhunWnFK6S
beu9ESb4BBlRaWjIhiOlVd/n+d4w27RRN5aoPTeyoRJzVnhKj0XKsu/ZNzU9mhKjxibW7XbrVAwO
h8y/m9UIv5gxURAbL9v/90GoBzKP7o/GD5yI6U27FiH3ntosygwT16hAi87RkzLclUwsfhJIbhc9
kKUfT49FSqCCOFckUEFMAz8tvmep1QoBr4K1eMj1IiUHAxOchX3418kcBTzkqSCEaL694V80t7xG
XyGHGD7wdaOJ3GsFA7AUant4APeXHZsB1quqZNxo6+37H2frZlgWN+yv5fnH/IzvUJ68/7jP0V9c
Oxy/oGPlVG0RnVCwbewRmGX8h2yBRJuVu8j+HK8HdcwFGUOCOk7P29sSiJZ+gmL7X6Mhq5KMdn/N
nmXlbxaNJSN9oVz664KsnpjLdSUeEe6ADNgdv+K6zQp3JQHXJOv33GeGCkVp2ZN/sMN2zJjQQVEJ
RZe/uaZ2+ziEfOmek+Stwxj7Hac+aczIMjDB48UZ+0cY9XmwYt3btnz28I4uGqUW2snXwgCGypKF
uDPW1tTz/l22tZwqeXMUtbAI+GUMTNxw8AS1T0JyYx3EdtkhpbUNIAZNkgAUAf5QUnBSZTRAgMDH
cB3tNeENNnJVtaVDP7TvMK1vCTf8RH0cKhE1QjIz5+2Ns9iMDmR2pJLkoMVUYNTD/dmss7jRsRK3
4zLP93uydSyo3AsLfHBtjWW4oHsZiFRagzxa471MEySEesLA8UWF/QirSIYW7r9CEOF71wGEVC8C
vT3wUcXR+q4yWz3YDFJ8n02umAOfsZS1ES8buLSPnEy7zOGq0p7RwU+vwS+2LzLmRtRS55l0BAaC
15MFcAAWEPA6Ab+v/e+jSF1NcK/oT/4OBifTp8GI3jZXxwPZ7RtL11E4YKiPpk8P9IIy/wjUE2r7
4Xev1FieT6ndztSmxti1hzaJCNnm96e0BfVtHH437LYxS/7ZFBxwAKnsSlAzfPl2uWw0UK3cLn3o
6W8pm6reLv1/pUo6Ga7OhA7RfqF0miyL+vQk/eMHXThxUgVnKtXh4TcQHohMWOY83E0W60Lb/oOV
B0QVA3lS2hv6SlS63dVEI6+P7ed2xYjP8/z518mlxwzIASKtiLyGISQpLfpzDt7dabzxLm5HndEg
VdjbJsD4yirX2S8aqld5GzDh6wyWago4d6PtY7MUXf49NFzGZPWPxPo504K2WI7ko/UaWr+J+EPY
hyhP/b2xJtMRQHc1UQjFLJgfW6j3OUd51702/nW8toofBqJ6mW7KPNGKM321Heln3Wfzsw9V1ZAp
pN3Il8xUwy44TUIszpuoDbsTU7Fj18cXsMqidfjjbS8GpcnESPFd7HORPQ0lQlkGAB3yTX1epNcJ
ZlesmL6MIx9EyEk7w8A3epYGor5+QEdv3RaoBvRN4+etnL2fK1vM8Ex1xTyjn26Ct4o6pDhTZr9b
ieMGNn+JDIYVuykXVKo8hQrfz6wrOHXMBm97mz7YzLJZmAi6411Pot1jXIacq7LzXK6zqTcO8ryy
LsZJjLyP/paMLVz8//zaQ5kB/EdIO/NP9auUKHpG7+6aeDPNLPAlWwM4VIyK9Tih9kbmHohBcsFE
G95HrGC5u32SkW9UQ6Z9t1oEpANKw9Gag+HI6W9WF8fsH47oLSazirlpXo2d0+v4Pr0WnDHzMvgf
foMMtBrWaCyrOV66nT98sC4/Daa/sik/ynd9lDDG+rqpCSKl4DQey4zxVBfWEPK72X7+7pLhgHrk
MA7dHMhztgUTYEQ8KW572WZrqvD//55lHlUTVx5SEAgJ3c1+mnUQ2ZmLLQIfwdP6t9FtuTKuDhbp
7SQUXsQkRjQm73bRvWgL7CLNosd6oBdyo/bJAuDXLpBr1KaibvZlt2Ytj8HbWnVPkSzYO4Lv6Lyz
C8sNQoMuiv2vIf3Ond2e6ECicxHPc+Y8xgKDolEMyCHT20/ni5thXH3TnXsHcfCn0MWWRAbYBHom
6MLcjb2Hnzjs+HlePQV0IbKAICx1ensNWHl2Iaf0bEI8ZwXkoodp2xC1e/Upb8faznQw774//7mm
/zRsIRBlc659By/Sse0bDjc677b/ZYPl1uT5hR6cmt2qhTS8nICHcp7DLNlWzuH6bgVhIupXai+P
W/dkChEGwz+mRne2v8Z0FlOdYMMtJecXCnBcatPzYmuJsZOSp2dJ2bwOf3nP8DBalYZ0IUiRKTlw
xRqgZOf+uK5DKNB9McMVDfaHHibXk2ZBm6IGr4TtKpWkNsym596VoIVC5UO4uWTdermnJ8Y0d4eG
p0tIXAKqeZcNZLwp7DrtQWn3/fxFjfHmIvcmmtzfazuH5TMqtiFuKgZr6iS0pmxeYq+3HKrCFohH
jbXR9KrCjH+3EsT00FiAup0VACZsHl8nVtRCmlkyHqNxzZAJfhhKcIpWxpoxbZcdusx8/1fKoiMI
YA7+SL5cpQ9UT8O0QFBT7Is+59HXkTJidB4UIK9I03qcGqM868qI6QhV2VVPHAEthOAsvyX4F3bR
IqGmgSUjeLLaiSyh+qEjyMKqv3u7pE2cU8RMqAAdfJM7Mh0kGZfJdP+vD/pQUZwYIowV8tDQs1A7
XZ5Xfj1KmBzGgI4EQF1bjkb3oyZs1ENo4p2o5c3urEeuAZR9RNKLU1VCss1DJkNEbZD8NmK9D8GB
nQFTDhbLBTydQ01N0vwQ+8tDN5FBhRFgdTJlQwy3rvyJPvw6B3PEMEqkyIUxrKShjNrb2iZrUExx
6T8N4a3JDSx3ukYf6ruLvc7N6ThmT83L88tkimT88eLofdeFQoRugUiQ7IuMj0ye6RIsOPX3gr1i
WoTM7PdemkDRH5YH8tQmUzDpjX1MSnwpbDvKcd+20qC+kNaxOAQTBjNbNaJ7evw7Ibf+OUa81d65
sR789W7WDMx0t9Q+LWRbRrum5IKctN27dFM2hxUbX/GMwO7kyD7WUSfSLbwUhDcPoT8kNVYX8iAc
blGY8eJor4ynEj6EzqZpBjTrPJzyQD7LOlJZr8k5ejyDlHHO6uL6hHSt4koTLwY80oGn0HSZ11nf
Jn5phrCJBUYv+gEsEICnxtE5Foe4Al1OzPvS060X3kQnl6FU+fcmc9JMqB4Nx2kafQgujvcdMO7e
vo98+hDm4v9ZbepjJ91GbbllcZS2lnFd+u8MqsrePjy/0zaThs46hnBa2VWR2F4KHvZVhgUg09AT
cG8QqNqVqS85v31JCjzcHsDTRFRvx43gSIlXkoyqxIobHy7IdO6U4iO4JKj0E+3juwvTIDj6cobq
g8T4fWC2Y/Jdm7kosGwS2Yi6iokSKOR7RCpBkQ5YpbftkjQq/nsBPy9TnnpmBK+2Vasbp8PfDH5G
9eKeoUPpEkOoS0qP81Z037lrS9DDdFw4R3pjlTEYf20DP3ogTaXj45+Y0ZdgvjRj04W7+ByDOXjR
na4S/UrtFr9jKv5J7a+hQwgrEyXDEXQSniuuIAAeDvmlLYD1BoeGvx5eQvsKP4+HxMwxW8oNdPNc
T9/AY13lNyMg4P9E8rXRoZ5H9zOBF4WRrL5Y8nKgSyiwj+1LTYz17rqGfFHc6hIyRSISWUQaQWLG
y4uBpR9r9cHTI6CIRp0Yg97unF8X2VR5Inkz70jU/P7AJIMtjdVmhcVHHEvDoEVlEra+pfgAdoVu
s1HH38Q9yKoCMwUU3YDhnPVgvtRpK1tjKXrd90f6N9pnmU0FQLoeqsUInfobXLS9LGWS3O1az2YT
GKcWeIvJPbzokasDGgcDss+pLGTKxUvztIpaWqq96/uM3H8O5OTiPhO66sEaT8faBpXxXg22Kj+Q
LBMLoW5evq00sswcfM2efsQ8lW9Mi2U4bV9kwaIZSmZOXxA0sXBvnuo51ijjJmyy49H2SNqVOS45
mpURVcckX4eYtcFp1vZEtIeMBRC85Cu14mnub0L3ACPfbZPpYItVR0nyCoZGPc9QqIGdnq9x/1WB
pWJoZii173jOnBDRJq4ZZYEwNhNkUZwDnMtS5WZEceczbxGV91cxpEK6M21cMZMDrd88Z0ZGf06U
ar4MnOwRspwm/CdYKbjuP9+1xf/4EIjwM3tKs3olH5k/o0lbjzh4D34fT5+v6jTMO1MAmUAbU4sS
DQFjAE+On87n0CsWT3gTU8LNCDqjTjN6WB/gBggR0Y56m6ddIrWXaG1hvRxCoB0xYeYm3n3zg4HV
kDkMXj3awXtcC78DW0zmKijU2r3ML5oqkYPyJIgoBY7JsqI3Al84YxWnwg4vTq5GJLCkYplPptDm
RRACTBXNoLvsyRcMaKDbCIqF21gaZ14e+04J0+H++m6Xfj3zYEzPQjzeMjyEKtCBCaptTqNbkRUv
YI6cdA4z0hY8q2kArPxx2skqExDBUBOKKG9K+XIRc+0iTUuvsmgRidc2+m6YLp/9dFuPNK6099oH
eAm8/zHuCI3rKoC1U2ZHz4qIfFpgbKAtlpoEYT/cDKP+NXjnGOEO6B7oU1VUH28cHoAMVV5OqivF
R+vi+8IG3vXbYc5fdpylLNW7rjZkhT9aGpbjXsJNcvwN0JV5N9W81721N3eTQhdwiRLPbHGveZQ3
j5yRtOCrEjp9XW4XRG8M5eDHzIrZpzcI+uiVvZt9Agu0oaoHgIDJNJ7vuagjX+j37UN0h7QxOR7d
f6LWabagF94CnKg0THQKTpoZVYYb7/+mM8YyhhZILoMYnAAaTlfQsaoeu2sfQCb04w15u9M81ci0
wTYdLWhGYyOTt6rk77wuEPF7J6umY184VIcpeIwEA/ALpRkOQiVURdQmCf4zqpmSU3vp9/3GlcNy
ZErIvlr2YiPLmLY5Hlrg3UAuLdM8HEzI2Vaxr9l8AY7iLaQvlRvUU0Lfbxo6+N5LTfNTR6rzxh2N
sthwgzwExJ06Lo5p/zK0KVgxge3ESCjtdqS5aMk6coSVwY4eyedO1bcrbCAmHIcLzrytQGn5F4oJ
R6Zv/p+pLxllMMHY/Y3uxfgRmUP0SKJSKm/Nh5m+4QXWzsab94lMj7NZl5T6UGVWpufSyyPacUke
g09tztCR8g4njSfa5XpQxVLoj6D8sbWnCzIgcVXAaOVvWVM7eDzGWObe1/8m1nX603BfNME5e9Dz
vPheudjvJeHQ2AFb2+b93l9RcXcWP5+W5qxq4g+LDQX/VAmZ+oIAWCjNeA9dWVYr+2WudYaA7XYF
xzvESx2CdxBXg0yMyKiYhHLoijO6EaFFHybiuzjW0yDE1KkXHnynqiUdP0BLhFRIDlJaOO6z6iY2
6BC4LHI507pcQ2dtfS6H9xE6lgZzJxaMDjjspOuD6Nszhvh3rfSmAB6685I3vQj4HIDWparx2sUr
rcmQ0dZLMGgWTwKUZK4UkhlnFFKqMw4b6QVcVoZh7gbYQv0R5W3QsOiwzF+UKj6jrPN1VChM5wav
Ohm1nsmF+KwBgWFlTV5BMNW2KfuV29ZY5FJvC6eZNqfHAuk58JolDr26jN5vR8cmc3r7Y9nbJG1T
YPKXOcTOD3ftAjhjChYiIhDQENMuJBgJXdMRPHZpNoqXpH3PAQkw/rmnunlwKZuMpcBbyoUyEJOs
T0d15M2MA0zaRXl21iC1wqp8zgq7Um4/jskydRkRtHLDSU1vDEUhOfupkhk6NNGDAQ4aGre+K63b
LXQ0SENqeTaSDtqJndS4IAS/0F0EX0HEM1r/FrVR6m5j5xS5XQfJttOzwbNYfXeBeBafxKlD7eTl
ABkJk/H7jgGq3hTt0ZnHQbxr5hi7KELz+grahwfYgmn3dIYM+doeLgqsWFkwFiz0kpZCbus9f5SS
9Uvp5HzJQGV19arECjarexfYJaPCqoc1cyEz45p3TTdf6IG0dcZExI4bjJtjOStxJ6CWh5f4Uysw
fV1YoW2mHWpuBD3TXcBgdNN9RuzyTiCGEeBO5QaKuhADGao3qwBMGGCWJzGyuhcIf/oVnLIqtgsj
FImpiqEsS8JZk5Fs4yOwjRiVs+dQb40yDj52n1FQa4BuDhzG49R/u5ZAwn08qe19JZ8+RsMiZmH3
3SAsjX6RxNLpgQCKNXPktn7S3U+p8H9E/pbuHR0ix0uTd2/M9GWlFVEf1Psjz7zi6htBrcHuIZwv
vBsittgDgLW6bXMRqahRZeHjOrHx0XoneNnr4M9ko5zlGsDme3a019shG8jjxfKO9yrv0bHzdazN
19kHt7XjGK/2U5T3IxOpbLZjq7Exy0T+OKOZW2rCC9KabLFRdq3UsBhfbmOfeoTNPLQuKcNRqbwB
E87dU2S68GcOLtAStokuGlwAKjQEabnHnZCXPRTImYEnknXpPxSnBJ1Xntb6w3R1xjjJ9y/KM25n
alrcTvHgjvkS6jUr3OGK+sIxf2XGAvqp7qfvzQ1+Tur0geLgpCygWC8QT/yAJ00svP4CzNmX5brP
REp2I1lRWu+uoe86q0mFHjSJwNsXCvitorn3VqlDs+4eEc/6HhwVMx+ulhvJYRUzUhmvnHUG3wD5
P6zQMmwPr7NLU71rrN79mDzsqDXVM6tKO1MG2R0PpUIGsYO5SbjbJPgVg8TMK6wuCAEZlSCkmC4D
WlLd3+6ctaSiQkbD7SAhnLAWvZrn+xXNSXzMskdn7dJyL4Qx1aRCzjL2JkU2cLnVW1RtE/VtXdea
OlTnrYwe4HFsaDhK1EQZnGkgMArtNQAXrCaDE6p4lb17ufzqM0TyatyZ4wjTM6S6aagVZ/XkRdJL
C0MjhnTTC2v4dhwTIC4FpbVKaeb1nzu9nH4w3bgHgcnYYEEnJorMh0huFuqDwi4dvMANx2zmMeuI
2dtaXwTbyHHKwCF02jPHvuMXsdfMlF+jvB0ohcorOEqFXJbPjYiTObigZZ8fI2KbF8B6E6DPRYVs
930s62/sxGlLv05ga69ELHFSqWDxQb4rF8iP0y1Y56W4JdkcynYog4AdSu2+JNO+F6vfnG0VoHUD
2niBcfCzoLI/Gb/eS50NuNQwOtYRADVAfz1eGr9n7RFYIQXJ3P0I0m98G7HZ2CUIGH7J2xDoMIaJ
eomX4qSzpGuHis7nN7CziI3E8V/QBe7mixQ8fxRzrQoDXYtj2W2NvCnSF24RoRyyV171SuKG/I1R
GK8iKlHay/ztvJuPR681+94JVJu47g4jMRqv2/v+95rdIC1l2flU2+D6PaV8KSmyENjPfB6oz1by
vlBYtZCY3jlVGtcqeTmmu8ZJ8u4u1/wOFvDD0/G2CeFwOc0SBM2ZWaWha1nMHvYS6Akz1rBOUqN1
JG0k4djNdh9kjIQj5d+KCcCK9ljqvepw48nH2N6C9pjBFbEDCX3s/9FhzTFv/CS8Fkyzbo3FAOLt
9+hAh7etp7Fvszk6f36sBCzsGv7xvywipZ+7SyPnvxtpS7rYDBjkgNOeYY1OgegzMHv2IPjEzgLm
Ts81f1TkW/8c2fWo5YxzYZ7ODR9Lo8kq6KvC6Z/4xFYC/z/P3jd2ZQPgF+mdizsru7Z44Ooo3XsV
HafdSbdOtFFEuPvZEqttn9bVqItylsypygmmjWY1ky9xwstmYQEwjJd54kj5sL/bYX1OABfQc7+7
a07S1DXNxDlXyimKfL777FkYHVcaJem6rRjHmjK8NsF44GtNyrD1q2o1/qbZB68Qb8lF4fDvdrKu
zYXoMRZr8sbpWoAxY9HcHVZN/XQr/FhcofUBgfbCzk3q7wHz+eTiYVRdJxjyURj3Y4En57si4ucP
Yji2xL8KSJaf4l12XFkNIuZS40BtFz0oefLLntHcUsptlAcUBSlYRlWA7z0JkzVwZC0JgtksFNWr
b9NFH7T9Q68ChUuCgxDWFQJNP9Ms+Qn7XL2TKdK6L14Xnyc+qsknmlJAusToZpZX/UkWbYbBKCuM
ezisBmJH11SiR8FxW2uxPj+mkN4WMUu06/gneCYqYDKbZFWfNyS8CjWzsJs5ByZJCXJN6fcV2RC0
yd9aAdGibq4h553esRUlWSsq5G4TecVSI9/0LSSVRiontT8xqvOfF8AFXedOwjYG2rJBApmMLJ7j
CE41NgpON7rYkIsQW0SzPeubGhQXviAXFH+k/PUzBUU4wzuT4b24XDzyzZ+QjdLcEI51zg8b7Tc7
LVS8N4Ita/GxftlUVtG9sGTsxwL2Ne31wL0g9t5gcrfgBi0ASmQU62MSRJhcKgxpLIva1hvmXc/c
9lZZ9Z2pcTWEFp8uH/iHJXXGfzAnnv6bn8Yf6TjMU+n9irOgZdMAo3rtp9ChQho5IWKr+3z5d5th
bq6cLzVCI9QO17DZyPLiYGrvOLs0sQQmREH9Q2/Nr9y1/ZxJiIVZvZWQtfGXSoOqarfzzODiAljR
+S+2ZQCJ64kIYnVxVjCY1FGEAjTHmgD7veJhW7aO+dVkewD6lasxpKXRsoLDDt+sne07g3l5FoOE
kFFDhGjhnGe/08ijqSHBCV4cREpjuzr5J+/2tBUhLYJLYpaUg81drb/rYSuNYzqFrdQJbt7c9PHX
1Lv6BqR/VMV9jDgjVmII/mvO0qeVaws9DUNUtY5jEmSR2uXAWnNCYZi4D8Fey4IYG/+dY3Sm94tl
rZ0qqToLkSNNNRk6t9V+ZPocJ10iPZMTAqOCdFhhatghA2PN171vVEks66+Q91f5PnHtdLnrYjcZ
+CiLEDPPSkqVevOtod2ZDI/qo1BAl06ZlWHLVGHHaqd4S76CHGJGGje8cvh9eRNiLsO27ww3gAjy
T/xpFNaqtck7/pS14AbNDkBzWJE8phgRrfu3ugXyNx81GOoDbGeULDicdUamPRtAOlwoz04QP9i2
58uf5lneMP7R56hf9dCxGSNSFejwq2nxxTVWzDPhE3teLmmC7xjQ3tud7rFyXt8mHLC5eymwjceR
Kiaikvb43G+bP1seqiFK1EdzN0VvP4ndfzVsyrZE82B1VCeWfykay9u1J4+vbJF/beqcFw9U/Ub9
vBlDsRP5KSG1LGx4cdPy7R9VvtDE7gJUz+9f38qdixl9VJPvqtnTVpuWicqjIsUcqtk6FvygcW8x
Vz81SG5dbwpCSgEArqclsNWk3os/vZJxrv3ZDJGwbeJVaRu/s4oDVtIVEG5HV4zbRjvU/NWDspDO
9D6sT8Abc3/VOUeCZyn4IleUKnNFo3NHUOMUj4A7W+gc3JcZshiMpuFm3Y/p9xemjDrqTLNGBnIJ
DSYNzMPPFykQXv39Iu5JIWX4201lLNG5C2jg6DkHsRtayAEjysg6f8KrLBk1XImcbAq6xIUyJD8S
kyolu9YUZu1L2+WJvLhzMD6NWy58TX2tGCm7nYcbmAGq+4FvrlMkCFeP+XTtxz8hrXn/CGcKGlgT
2FbE5301bdpAV0xWb1fkD0i7BA4BAHVqHBqRjxYhYTScqnUranjmEJ5z6+yPXMcwzSPhlov5CfIQ
prH0Np44d813B4bCo+++2KMzLediFoEBp8yxNYErLRo34+RuSI3TWDLEt03jsPxN/J8z+4hAyLI1
6xHpgsHMaWfqE6egXKvfbPqlMTEHxu8HJV8TrDCCDTYMMm9JXSfTd/MyfSmTuqIMWyZck2TiT872
pjyhApdsBmW6/F0kv0VCJ8aY+/PejG6mUAiROqFFH4vemfJwy8n1rRX8SJFKXyCqtr1OBc/nguUr
2z9T0ikDs3krM39ormq1bA37vcHqULMQZZc23kAj578ueXk1T8FY79Odt+5Wr3sruXvA2d2gK9tC
/oPLQ+soi7ZPkD2UaNjhEmdlHjFF2JdlHCKvRZytJh+/YOKeBRvfkkFWV1i9g4u6S83KHnbE/MUz
dc7DFhgJ2VGVThnK+oT38q8Pt6toHD/laXZVMqBkK1IY4BjyMNIp4OMA/zQTst55/YdOqUbwQs0r
B+rDtVcmL0/IKvAQxpNn84Uqj8hzhL0PasUpxaTyQ8qpcYwXR9iUH04h0mMu2M98wYKkaSgzOJ83
ZYe9ZlBqpt3h6yn5W6CXJILxRh48zroBM8PSvWjij7hKorrU5kcz79C+0w0+v38R2myDrJ5LKAu9
LmMYm/1fWMsHO1Hds3DXYXkjXXM6wsipRzWjVA/cFLAEHAv78/1z3Dl505CeWAKnM0IzHW8RTIs6
7N+PytA+LkDN16wUQcKNQ9znsU9oh91nVmhH2/kUisbpAcUBp4eplYAvy2zz/1npk55LDqvsgSIR
SVNlbu8uzTeJz0P++te4yGKFegYzdC7HFDqZDp1L9hY/RIJTDrL99f2iATA500E+SAbwHXftQkFT
P42euZtyKzYIUoszpmykhunLWp6STxT0IU3AaMnc8DLRBkDtyj/6HwPn8pJjg1xIb9eZ8MSQI0RL
+JcbG7nFn41afudHLyDpFhYeVsunI96dIRbXIDM0wT8O+0IsHYhYdrRnikM5U5bEXAXOu4UfHmRa
yAv4ZDkozlzxfR5UZwCRpMkGPakqz6bWkcLz9F+Ud7wjg1JX+kZZfuYrRe1ZTioYtUy9I0hmEA17
gv1shWkTgk8vSbO4KYvAoTyixRErA6bdGwR9AM5rle7VTRocfrHOqhy+KBhpsWcvvvXDdhDXXJp1
P+kdcno98JfRoRzkEgoky1eCPOYHnnBRVzC7lHSCuW0h8Et5w3ifvSnnnxd5sgSXT6u670EpQCsk
7HT0/RD1yi200RZafAmUxf/xTYfe526EUJ4SCGNkhYMV6L4OZ31ecWoIUiro7XTfk2RLUMjqodX/
MhIO44JV30Nyo9fVglD10X1WxwLure3uc/WuEdiR9SsrPXQivmcy6ZZLSqpD1D6gFDVWCqIw99Xw
xCxfS0WECQ3J4HxMHIKGS7Qsl1wutsPhhQkx9c8V2vMvnGaT0BpYzXFsD03oSlnU1GOsLc1jIyDh
aSs47ezRTBFONaiqJQWJAssYRF8vLLUtF58c8nSfuJuCwRB3G3JeTE9TXWwB9TUwKu/W4ifEL9La
QozMazLJ4zIORfnvhyzu1+u2M1/Wk0k00J55DdyDpLfKNqFsCZqPn3bB+nQZUH4a8KT8ha8JG+20
OXgWYdrJi1o8+E9iIKI4igmJArkLvJGOGRT8vdFrxQL5RW+NyVBOLRA+g8OoO/lDTDpBYHQXdFhq
r+fl0KbsUxwS8f2r50tk611E7jMhIKQo85MDyJRqZS4TRLpmByw5s06hUbrb4ORe7p/ZtGESBcFy
BJxTrpBaYh9WgJ9mg/r4dWeTqB/cyf+FksThC+1JoIaser4B12W4PaMj1ayeJ0lHkkSe6xr8t3xD
omj/5/3Cd/ZhLRXZtMXQSagERwkKwMVZXBpS73yGvSfiLEa8AllI8/Oht9hFQzUdBImJ6xVmY40K
VYSytGitxpyW8wvKeH2f7dLmF+JIPtGCCDQKUeLsq3bcLf3oK0ug+04159TL/7WgT1PXN/dAPu4w
UPiFxIuv1C/UZM27t6383FM9m6JSfrWvRoyCorwqCfo4bVl9JVrR/QiiTMM0Linpxze3ATYdG02k
0nlZkqX/CqHCIueMgSFcjXiZXvFk7Drr0hak2Qd8/v2JnC39Rw4ZCZYfJ2OLFT8bicLNLQaTAC8+
yI+aqS72Ek2p/IBwZDCS15RVli5Hi2s4C9RIsEhhUvSe/WaiFgGH6Y/r0tsQjzV42Cdzhq/Xb2IR
xQaSpRrobTo3FEAw3nEQxhCgvoqjXNxW8a1QgoqW3vjjEynZIhDeLHeyFPr2jXeXYqN8dgLWPbFw
rC6E+Ul58cpJ4JkBNeRIwCfseYx9mg2QyYWkfd0W3JZWSpOuI6269+2cR/E+zDyZoxJTq+jsxNVg
DIhD5vTbJeaNtmZdLss9GX/MroC7U3w0wSUpldbXuiqIv9ZWmBOJd+iSZYYhZsPVm3BjjhRYdRGR
/jkdP//2bvaC+G7Qug3DoHcyBBqA9vzqHpX2xjjbvD6YTbh4WwtmlVezeFaHECCIxoT7Pp1XjRPB
Ns7uQq3j9QDqsAvzk/qPgKi3p6367FZcjCjJmn2JONyyPOedMKc6LNybZkl6xmUqRS0LwmDeg1ua
3HomSrFeaKb8O8gliMZS0F1zaCA5tZZPBL/5cTllLCPKJnvm0K2EQayBPV4uyrzcLzPHE6oNAJv4
zTZuMRrcx1J18ECP1ICaTVAM2vzt8CH5+mtRwBh6K/eRTeT3DHSIQFw0IvKkllDDmrGDnl+8+J46
i38PzbQCKHgPL1UaPxpbuRl+138Z6yuDdoUBKsJWCtChPK3s+NH8f6AubehqMcb59b3GRIHos2UK
YjiOM7n43wv8/NWEXTG+s4dQOi0yxzAkE+86UVuDJTtS8pe4qxZz/zWLBqSPVyvEoKeTKddKkk/c
vZYRHqKdNfijQgZQqhQp+Yhj5gUIinROgYpzYNpd8bJTeh/mkIQbmGn13VInyctB7WDbU5yVNOh5
EQdk4qA5Knfge53YFE9vV4GCKM5svsD7v7+EUgJFtflSH9v8l5e6YWUoZGkng95lF4xWXBaVWWbe
/pKhlNDO7NEf8clRvWPrOHL4yuW7EV50vBfVevkVZStlJ6ZytcUgMlPplyb69qZsHp4buTmsN9IS
Bc/4RVlBmexmJ7nCO4V990tOz9K4439PhB4wwCtzmsUMyTZYwuWx5Rxi73EyxokhcGAD/8mpDXGv
M65X++v7GW7kMC1T79zPgRMA1lMuuO++raSiIEbYq4xi2pT+c8L8Ku7+t21or0TBm2KTi7NrFzWV
nM1Feel836yQwLoOFZoMu7wseEdBFJefQ1iMyHvoPLGpMe/S/Xg5vo+/V7nXbap7BPkvo18Qc5jz
xC2ws1g31ICZC9LFFMRi8ynk9sbnUdjROGujoGUnyRvLqYlKDryCKPC31naBLNS3L6o1AtTHBWOh
B/O12iffIzAahlzbmylDUP4cTo8OGKYmd4InVRlBwf55sBMD/hPohiP9sLZB/9ez4ENFmgmu9fCR
L3gxpIucW2zfouwehc0Oqrr7ECdSjklrbx5oaFLVckUlckLRSmPBb5kyJ2+6pldB10zoPnJDWx5W
CDOWZOXPgAr0+P+9IGNa3Mqkqox0sF88V3M+b/8WPl27RqtVlcVUHwdLmIF19/XP67tO0av1OQzb
ttVtRnvLK+XiwVKO0aW8d0ZwkwJ8uTeHDkVPTzX2PKQ1uQOE3TLgESE2WH9rLd78IBcGyUOC7+u/
xwqKvjBa2go6jtWmx6MMRy+OyRsuBAGoA8CXzFbkpVLyCEu21abW9wypt5PumOg2gOSQ3Re/G8x5
wR9QKQngoqAEGLRHdL36lwmmK7GLjj/3mFET82UvgbQfz7gnzcVDWwPpRaI/73dyzeIOZD87B1eY
qtnTqcXUMFnfWBAHZ9f/o5lOHEuhq78cBLpsTNGdI9xsJzgkvHX6DEwOEfMmTnQMwwwHUP0JZlBD
P4beNPG6yeGziinwNKQahUmOQtWuqaoPWJlIlHoHz6e1NtWDH/USAjb7eBjch8E/d6uORY2tTgq2
u5T3o/d2Wvhb8GJIN3lD2jJ9xSZJPGl7DtpFPPiT5o/JX2qrq1/an3hn4F6foE9IYW4Pfc8fJPS5
bqlwvqWcg1nM5hqT5gTrwTv5JQzvLoJjTaQHdXuqlct67hZKOGwUVoIWeXyApZTTQhGKSsQCgB1o
AF+aDqclz+6MemJQMXRMEdavC9ZIS/dGM0ruSJWOmbCMp9/aB6e7SVKL6pxy/jQ7r0Hp9+jo4Ko7
KnD9TuiVywt8rpBazAEBq0eZl9/6lFFYbfYtyXNAi4Tq41EtJJ9fCd2usT8JP0wSPCF4zDgTRzub
gRmDoJpRsnEKpyEtc2ugr8gyu+uquofe9q+TeCZittf6KdE8CuspKADEGs9jW76tHwOPcMF2M9dF
fnCmjRP6vtei+oBy96ZCOvlUZqvm/N2iDG6elSBo3T4AxsPqtrl39Kslk8DzEggDgf/VlFUqnkqw
GeMeez4u8qs7Ju6eT7qGXb4yOH4Bzr76X5uM0TB6v6AnHzG1UGUaTgPKkI+4lntttJf9r8evfgqL
k8+HjKdZ6krsN3FT4uPgStiMoaFmYFWQui5fmhfHpEnYeDLKoYVkHHdWe1dusFPGuXvDclyld45G
wYNfBOd0Mhp9KsK0xUYuQ7Go9L7qBIwiWg3GQJibEp/7z6nBi1oAHynSNya6drGSadgZDQHlqNTP
1WyosJX2w7KnyFVPmLjRQlS9mAf0nG4eThslnDdCFFeV3Y+WJLPbUdJEtN4RWmgPleEVGQ3RY3N4
9Vg8eF706xvwND38Ri6YHpUAtLi30gCp7s34nctTyHb5xhpCsPGn8E8OjX4d71dssNnXJkgfujBD
5pACMAAPKVumrzsQKApntJ8daPOBLMmp0+BC4F4NVi8uvfHfhc3BOQd4t3B2AXE647DHIHQsqXX5
PpO+qSgL509IGID8cf5YvBZJ2O8xrDe9y1dTN7QTj4iAqiRUSLBPd0om+KlniK9hI7+0WNbHbyJU
TU+hzQFL55gxOhRhd/vdjtHKfJI9TIiiUUVi06q1roCIxx4s0KJMFYO3ErwueoKbE5llU35sPunY
MMgqkXmMdPd9pZCSHVrXb6cHlpxw0tbI+UDKJ5GSdjPgiqUNI3y/qRSE+BUm0pRqybQQpN9sUhsJ
UndRa+Cy2UsN+4WtcrdF1DMJ3NCbENX+cBmNtjmu7k3fEDd3gf5m0lazYHQRqdIaIV8psX4VNESq
lYZKSRetK1tJrNEM0gPVlhHlXWdLl2Ho1NjUAJB4/DlySUXNuAIrP+w+xyEC2Fc0KILdIoIJQK+f
OLF6WgzwC16py3TeeEpf/0EIzUWZknakwLJtcktEEbouBAr2ZCdAzllZe8eDz5UedL8TcQqxkDEf
qL8XiUeHK/WwiNwWkb6Z2B7xPQYt1aezNFP/7oKjX9T/GRhNGMM3pa/6JPJjGQqAxCOaHDCpCwXN
LrJCJaTm2L+vFH2oesDBn86ZVtigKwDJOrXQcRLIoaECPjy0KnRvZojFa1wN5OmuOWogmIEph8aM
pjZGXVE5REpvTEVRShpsp+dfgJEBN3KQZOh3snSxwMrkexfWWcpnwaX7x/0l9R1mJY/SNHGNx4oA
GboK0UPX6FetZwyJCAHA5OunJy4pAQpNaAzlzkuxQn7K1+fpw/89vv8SU56Qy1MyaBMewGkfe4T5
k3qbu4LQv6577cvGFUXwcNU1MkcKgbxil3kMdPpjGdsUccFQZ5ZIGplFyZBlAHL156IowENU2cik
YiGo1PvBMuGfEJTAjxZjLsE0mna02WrASDn3zvPmrg0Tw/ey5hCjoJctv7IP+nUf2cVOmil1U+Z3
/Pgsj1GRGWhO4phOXnXTN/K9mD0R7gEJEGHjxbzfLXtSFQ6dI/nSK0jDXW2xTJr03xAQewZVHaj2
6x6zrtZ+OHp8/bB659VKpnNS6tU4FYP2S80tJAhix8S15ojhPpLtQnb/L12Ji3mcK9m1wkG6oG66
uY0ZYQPNXFqaovExr3G7R1F0XGhEpbMaxkN14uv5KgMrEXe0jXv7FpZsBp7TWrCIr+rWfFVPkbWn
5DG3H9b+imX1b9XZ2UNcogGwB3l/bpeMXA2+WUEzT0RwVEGvAMQPymc3KKUXAT9KrzwDhJz2IUih
78oGB/lyp7Jieh3JtqdjqAouKAFVqFqweyOwIFfR1vNl00CJt/C/E3gps5C0VPlwZVhhQwB/Oh1j
frIxvkEzmTGoN9xqgl+eDOZAg1XwgsXCWqj7pvs+f6Ip+ykJdRpslg/4k4GtagMb8SocBQUpuwPh
0tV+tnSVv3nE4s8LeMY97lDkOLR09unLDJeD/AsS3Ij2JZ3YKs+9Xwg9k2QzwCoDrvGJoDvOVvvR
+5YmSdM156vwAljkmpJBYWigRIMgYk6lnDLTlzGqokxeMzqQ+lnQ1yqQciTml0QzkQ5HYRSfW4wg
5TQPBCh5Q131q2Mpg6B4yW4azwzQVdnMbHJ+bVd2UCB6sVP9R6KD50prdc27z0iz7cxGHQRGVE/f
PbJ3iFyt0fqdBE16Thq590w9Mfi6qorVnJ4eH16phrK2aDEjtHqydQBqUiPLmQVrqLytr+Fn03co
2n110O/xEOB6YbX0YlKtkTUh9U/Vv2aj3v2KMRNZdcBMYVLCXo6jSmejEKEKKwrKI1/w6PpXzaj/
m8WawAAVulVm+dHuAjdxQ7/SV5gsrjGAQm+NS3CRS4tthe98wsOuUSLJTM99rqg1EykJyM/J77C/
73egY6hK+dMjl9Z8bVhES0cD9+5+fYRa8xacnazEX1CDbuy3BKSRFbLODWsG/jPoHnUf4VYlvOHE
vCdb+vXgtxq94Gn6vyxE9N+IB0WZQApo3+Xq5uFLOGES6FIZepo06bnGZJt4ajd7l1K6MiJLKlhg
IXQz1XDH5tPFBMZkq+LK38KX60C0JMZnqLPTH6Y3er02K5wUYrRfTvh7raxGmiQMnvll7W/zo45o
ROgZQpvb2LsWPflQay+fE6h+0ORE7tTApVfC2IUR8dXEv/oe77U5bR9JCZwHWwNqDxOWBJ+Xi7gp
9DSyNjORC2jV3fDBVkQ6Sz0zGrvU2e/3yzZ30AnzXMbVyo4jFAuhwm6he3S6xrdaUCN7LI3W9YJd
otXS1KkBIDhMfWJn3f2BoRz1IP6DZZ6nqMk0l6ND91/WeimiR3V4V6dhQ7sKY0kU+w6Y1JK0tTB9
ssOhQ3Nx4/Is1xYJIj2pZHbO/7+fZtBiclOojh5VsM3ESr34YemCIl5cdXESFSt8uVvXCSUv8wyy
riPEWWVxcaeAXsdmKQYKBz86UF+0BVCKmjazNIGG7+P60KYb74w8pQfnsjJ8c0YMrVX2K4cL1Eda
NHvRcv1D/XiRoayZHXon48KX/BNsTFwOAbh1OK3Y6ZC5Q0AEpJahhgiDt/57Ia1zh9ZJS5MdS2jw
j/WJC93wvthm7buLnLyd91E5PgTLbZlczey0jR5KOF0U7ZbgCAqPSQ+L+WIdTsPrXD3ngjlzjXvz
cNSBxRm6AUafBxELYbmhFdFXE9DUb5fdQgHfq1YtBGCCY97NJWIib7mY57K7ETRnfIMJEQgFi5L9
r7XxByYnMVbhee11vJ0gZzBlAjI85291MjVa4zJLCbr+0l36xOSMJtAxOZbWBHN9V+my4U57PvAY
tJodWORwcGUnH8/tl4tdEeUQWWL+hgKsKgSTHpQLPQaoSfGT5hnMlxw0o9w6AgfVr13xr1tceVUg
LBoU0yZNpksk8C5yG/aYVYDuhl2pdwZsw2suSolv8J/qEFu/PLwy92wXKgFi6kOpWjpArYCz7bf/
zecSIov6dyll+eMjnmMw4o/1BwsVsfxqZXypMj/s3bvDiGWp1UXGsgj4F7tNO9e+4wpXMDLN5liM
WYr3saNfnFjYK+BogcCqHJhtkuYGb/MW6GH8zXtv8iCtyG6fOe6ZgB/SlrREwUy2KFe3RWO0kwEx
83wNCXXZ8j4W3kYc8SsGwRx/etqbK8VTooS3NQQu+BjFTJOz4g5G9felW5MIhOzgJ0RM6bHCDQNT
gzrX0bjAxzCFKYp27GYkhvJ+Aab6Ns241IdAyZzQm5NqAXn/JnGtqI6i31163Y5TDnCOWrcUTxp6
wig/Cw027w7nJvGgDvAd6U2/JnubvnuWXk9mxN6CS/Wlv82DDX5BZbiEf21jT2mCLoWfWXdBaX5E
L9lnW49xgOATB3KblnkyP6NGKPNqxqQAJ0uli3DqFIQ4naZfAUWxLesEbMmuayL2Gg2LUMM5pyP9
FuKLgTF32ojqXVDEEvQBTXWWUAWJa0cgUnEVI/W8iouMg16A5FU5WaLXiEkhgVA8pIhN76+c5iZB
Gqoc6N6jP4q/sVugLDlYKbLW47/4ur41rLG38oy2LdU6a0o80EJ3okX8sy/vdx3clu6jSxjEJ3Pb
IHJODZkhsQCbw8qMolzSulX6pYOsGinCH8n+1BCL1PaKJMW9DqpONZxZQGFg+EzcoY3OpJCu0EBK
9FggJffIDvpG+wOSN5cBwfkHKVvKAaAGFjaTxPN1oG8AEEnsfb2sIWIjvmQ7ydTnGjXtRks8OFUV
qvr4uW4FgcNvb9jU056h0RbO47cmXTH3ydXWXXIGNZbKFNuBzfZK7hfqe7iLH1+3wNsXhS1u1Z1S
aPd2cpKYn31yHFpGO6oH95mMMlywUun8X4dKxOPWUK2+qhy6yAEQ10fODcAZEv3cyiS48eMTZJKk
/smWcgvchVujNWTNCmo3AsXc/RopxlvQ2m+ZBqrxbL1HZCh4btaXL5cESYRNtvKrO4x0DKDI40X3
rR4wD3ZnRNjk9ue2fwq/btvRAxTOVvqQjkRcE7rmbxcUcYkpqDRGja55fh92gsUNNR0pvxb+5ct7
1oJY2Sh8udUXzqt8bnG///c7RMSO21WO2fkaEF84Ksp2OohQbwZSBcRjhBOHUblRTCVbzXIRhiSd
GirNJu7LFOaTsrsds1ltbRwrR5f0OpWvXBFE/u+YVTMGeMK91zi9pe3WaNk/0eAVO55Esb9vh0Dx
CQLfHOyR7CMD506h9a0T/kjVGOui/HIF6qgk4VCbLH5/TOtMiayQhKd0ES0QQWek60PDj1gdir26
EJoFvRhASo9i8GI4151XPGT9jmi2zmb51gJRRR699fjsbt8SkEhVCfdhDBqZz9W82r2Is9PEssm1
UBVxvaiaByWmk9aw1yHmdopKEyBPD0XZfgM7YlfHhMmRyqiGjbtTDNLql98t3hnPnqhHOLgi8F/e
pqJJMXqXdXQvaOj0uOkfp67n8JS0KNF/THiyc1ihH/9bJK6bTmL3qvF1AleaIF3UTIN2/wGWTcNk
IooidTazTYsWJlTi+1IzElEnLlQkf2nKHz61hliRbjKwiilV20Oi87U06wQlG6zjID1bfBxzqqBM
h7nxc9T88/VYwC5eoOkUGE8CuhmauTHjAypr0Z1xqQ3GbZhPqEo+wSLRQUZYhOj0ccNfyqlG2F3N
ufrvW8g1n4GQrvF5jF02ZqAhW1U/ZCcZqFHyZ1nfCbx2BpDz5vnhuGIFViSk/Y6NIVz9un67DoK6
SGQ1Q3YuPdCcW2G+e7vMSpukvbDyCERoMuAcpI9BnVRUllktCKBAnnsOdr7wtfTx6feqa3s0PLyn
8xiImEErA/DXTiaI58/AqWF2YT9LjtStcwJa5+NQR6rjhBy8AiXUai4HY+6wXVDu1Lrks3zEhoXq
9bQzLcBv5zoPYMqzbc3uTtPkL/mJyzCpy9VBo7Whbin3Tf4ClZ6NkcBsJ4dBDh3TLtGoN1ncuUnY
IUfFLATAuzUhMjODQ94QgXWbVnqiaJQSTgKF+rsO6ke0h2EVd1aB0U5UmOS3l1GEsYazwNvmVvg+
uXyubPSaPPvoXIJRlB/uNosxbDP65JR4Yxn5/5jZHlIFrbWkUk1F0ooz5l3vNO0Hsv2CXyK916Zf
d48qf53oFZVXOcJ/rjeEKeUN2csGt/2GVD5honh8hBAaoLAJ2yfxwp531HqiNVf4XJquF7bLL3WL
gA1KQ3pId17C3gvYE6gOqze4kuMEW5bjDwCWH6PwZv5dqW3/4C0O6j3ycGuEJsl/ZZkRitKqyK61
Wngl4DINjiIMWLOGjdMTgHRRRb+n3ad00H3/Mv+zfKMZnVdWY8fMTwzvrZGJ085tXKF5ngVZxJN+
vtzbCGDMdyTqvJGA0F9voBYTxwFOF72+5w1ZRutwEj8LKaOHiNlyJujNeYQYX/POcrlCvhZpWMGd
ViP3inMQ4n0ioejAke1B9H97dcc1VfWYQ+cXCkrrPblavGsoyUB83ay1WaPILMaSScdC3knLEhHY
GI47FmM8B1GFsOLCa4QtOZAAfoikJ9YdLaLV3AMZ01gI4wBghfHPyzhq8gBzN5SlPmzFEA9aH1tn
UAmPdGFlUaK8AkAF2DLTxNXWkxR/8iT+IeVy/o5m/yl6qjcem9fv3eLSKV3eKg7Q/AN/0IXeEGDb
sVyNfiUWnpTsCDA5xrpau+df5eLIzcgIm84ULAXU2mraseVm4DijaiV7DMzHesnpo0q5AE54mV5b
Xbyk5CVRkwNSCxyyH0H9o6T8iV93Kt0alCPrYLOSF/Z1LBexyOKgyOBDORh76f1/lqw7eekj56Aj
dwkNn7d4kFIcTxukPvWoVxVzW6AzSxl2jdN8YHlKhFB1HE4zezUnIVeyqPEwpLU9/58YcW5FgpGD
P4WNnd2mhYCiKJz4Dcd3FK65ul/2swox4+pQVbfj2FHJ2i9ruLJdDEQ013PjCK/i6ye9qCBzkTKT
wTE5FmGXy2ey4hRwUztCnWx+5bEh90YwY9TCGLS5//vWLWLsaTsspofusjX3F4e2TS2Hh97vQNFh
xJ7P9WIkfhujSpzG0u/AKNnyBcvr2fhQRqfXmhGKZgYxMCIIADQqQJ06/GbSDrXXymEjbV6G5X5J
4vECq2qV9Ecj5iNYIAmtFcxr0G8cz9bYqpzYmJDcf2qrmcorOw2cWC+LyVMfhhI6fABJRuRjBvRZ
ch071HDOYt2B7ponnDgHyocfUM9rI1jQhbhTY+GuafnJO4yWmTPMMlKh22wRLnjKC0+aZHLS3CJE
3g5CGsI57rmmpte1rRL0osycRHbULrW+hAy6SSt3wRRHpRfuh+J757iZk7IXbpLHEoNeW+zMMMLg
NSpl3pEjqwDVMpEHcaJMtT83FNTASWP/3DujhWJfxOt5sIunZO+IMK06E+1zVUAiBalRFhQG/DQG
g1z3F70ASnJh48d1Z71PTBvJoI09rq99g7MuPsRwBtuR9WwTI9lk/EAYZp3P4waYYO1Eu8KScRjB
i6QNZzIJ4Z8YUuUfpDQW6dXhW7aX19V15YMQnOAn4ntd5d5LmbOcWBNPFr9zFCsMJVcmyqUQ+dVZ
oGE4YHDPkONfgkjNTBs9JWi2tq4iYUNgeRipccm5dPQ7Vkx+4li30FoaiIDOIyrJU3GdlssuauKk
f/xRUzdaLwkzUhDNF3UvZZCRRSQrL11UfB81u0H74VhzWhTNObni9gSomOyylyC6m6whQHOLA+XD
XVBQqjBPsBmhqwq82YCWi9MAwgJVO+irvVTP9YbHBoVVhZOd84tzEUPfiSwOP6PdnEPQsccJrnNu
7s3ZOKilS1m3n1lyNS4gFOmKbGQ9BZsqPYRTk5gw98tDX70WE5PHY4R0F5jXpjX4Ec2HwvlhdMf0
t0CzLqFeRwCgix1PwMI6LRDFtkgOeKvNt2mh7MXNlrTV/qFmcW/+5x7aZUI9XYgq8KvgfmhF/Dd6
44OuLSyv+r6QcJR6mRqM1pQCHvmtRwqkaPBzOOsFims1QfkPMf1qLIp08nbrUn+1GTww31lfwL+2
wLbXEZaZ8qyBkV4172NsK3pPibEcfCLwaBKbWYsmMnccPWlLxKXMcOaSLGc6z/JJ7MYxIGeEzY4B
ze5pqWbCaXWdbvKXjgDCKkH0cWF6jwPWOVG1PL76hneVEfEgGG+BAIEhVGhFj5U68rtcyjQkBouN
slhono3R0fttJlRgpQ6+avIWzybM+u0AFnK+UdLzAna3694biOZUNhK9FEmQENVJt/KsVAWn0JDv
uz3tBQdkDEuzF6yd0T1gCPdRH/97/8YI0Z8yNEETsvYmRvOw4tDr62LihzReRoPf6EPs68WKBAik
Ahf3iUp1kuzPgDMPpcU3zV09+SpKXgMCoKdZbLzWfET81/CGZZzBQ/YiuRqDDJIlNvsGMewzuOJn
zooZp6wFpkGkOrJhRTpY0YIm5YHq0aSKeJUR7QnhTNTjI490YAiWHrD7Pco6FsD0o0ITKuv3JDpj
unfbcyDWrmqYzqd+rG6wHj+XtDjjvMyT3EvVR4u8NUJJTBcGP6zJmZE61lKer2kAar155tB9ogif
n2/ImryyUsowcQBnqI6A30EaLW94sZiUyHsCRK41UDhJ5JQwuIUuroKGxx7D6DhY9TsGIXDzuIk5
omRWn4T5hzSOP0ZB2TpStkw8zWT6+nPhtQ/IUYMNI6x/WtfVIv3QAAiy+BEFzAwIbNlYMkLyhc0c
GhMr4x48R45LKq5qpPYPFOCOy58EG1m/Kt+8BGUJfT0eoz2PGXef9Hy3qdHIotJKMAlIjCLQQnBI
kHNtEJWiKSGpIdKSjQG4jppG5n3um/+yWryTtJmQ9Uqql47vPZUAF4NNd/7X8Eh562bPLIUUThCe
cWJ7NJGX27VXB1UKwSdN2FkGosc39ccJ62InL0zMPTQzJY+9wFaNnJb0g400l5zyfttn9HL5+zym
XrQR0XrGZkpodYlo0gL6ljEt9XadlfYDTQ96pCNrQ+uGgm+qEBbMVsTUJLKO+Azd6Dv+0SvPGwKV
IGtUX8x9n5G4SAUQFl5kb8hHRJZ4sFzurwyTwTtgtpoPPQ3UvmKeUisE6K0aII8vupMpVaf1Rs8p
yaLYjz+gaZTBdda41Kfa48bgZmpUVZ7p4CwTNtOm/eeFm6Eza/pE6MKGjzKU7VkPMtZs/0Bkr/Yn
0uPUBa0aJ+Mkp3qBqmnKlWDb9NKesgNhFudaxdoptVYAJgZvJ98hdPrXaUIoY4nnK4OfgaHui2VN
UXMF+Pj6AMBcenKxdZhyQJKMdDGWo3FaXJKUGl3xkomjMrLOy0jhmxZH9hBBeSsoUW9ORrxOdltx
0Oif/OMbxFnhHRIy/zOx72AyjTDfLSA2+3CpKmBzFDEHq+g8FcejAj+nctwUaglCm7KxJgNw+9gz
IuNVL81P/oRMJ0fykO1eCtc4sE0liR2tTO7gdn7TXgik9JhkGjKAl9OyebwfVf2hnGSRgsNNrJxI
+mpXwHaS57Z9HR8ij1BZGlP4ESlwNdjvLdRWqeGfhagojis3LfeZWZ3CG67Vee0PDWV5EgqACAsU
DetPddtlNHgt6i+YHa4X0aAOXeE3ywPxRAlqZxbgUOHL9ax+4zoRBdreTYIrhGCoHghLqr1ALPTU
G483eOUt/Jm0s1H53gKNQZkKNWUeeNP4YUWAmF4jCDPPI1/h5efSvhwd7Jng0XeSDvlpuZzmw5Gg
Q98IxNOztHZWS8A7lC9cfHpwZ/MMzt4ibggi56449zSMCBZvCJ/8FTdy7XnIbkUc00mZiXJtnn6J
ewnNjFQmnS76X0dU7mxgSE4ukF8ZGk4voeNa4Gtb1pIFHT0etu/vMnSL4BcIQNXOEqTQWRd4C18q
dJ75gBWka5epZVUzFjWxP2Xyd6fK76OtuNt5xD/WSrR7Fvxw4d68Z37jw5+Az1GqzcPHQNA9FZHY
wCMZxjUKep9AJzEVu7/Ui+SrcQMiGxXF5PDc74al9a3IoD5Zbyb7XhpSqs7FfbI3L5bAvoNniUWv
zT+mCYu4kBQBoJcFSjuJMAEbwca459vPCXrAiErEycErx1swezeGkIMUfsTq5O8Tp5Mf8uTUN5yZ
Ngdm7pkpfDu2dMdr6crBjQoWMWi9ClTYGlf87JB/MPF6Myu8fpxK5tPPobRAKNxyAL5yRPVHGyQk
qn7s9hhq5T4GikmxDd5aieFafHu6I9dWNoBX2/ykehRQNo+/znEPbBtt6RevqFRG8K/im0NS9HqQ
fA8DfmRli/67JiOkARZ41yn3ZnPllpPi6VIBqsevJdF23d3Fxf9ZMowNTlNKyZmPtQeucbcwLpac
mXDs6HrYM7e5jMtJ+pewKzeJsV3mvsHOovAILTd1MnVfs1hSmMfg4j6XTX74RUDA9Vo7lHMouqnR
xTmnZXYAKDXlDtRx144OyNHwZEeY6YoJqJNMitt+k0u+l2SjDo3axRNqFyqU/hJTzxNFtKf7KyJH
ECM2AanySNtfucgnQKemgnSdiJ9P/s9I5QiYqSJCoFE1fgZUzAkQF+lCilque67UO/5KaaLzUjrJ
OMPD0d75+czLqalB5s1TQ1KZFa3rtFSEJMAA3zMPunuBKJyZAT6Ca2+pJwKc6oxPTcSaDaZiNv8q
MeOta8O4t/losFiNfbgo/aboddddydtCCeTQsif5oBguWEQkOnqzKzFG0lTkV6PO9TWS5Cdb+94B
SysxMLdGEeu2ItV6QSzoGobXUYKHcasePvcmUBPdpIAe8yklSq7iTQb4IZwVqmCiY4v+v7J4+/Pk
XUW0HvGA6mvhHVNC8uwsIULfBxV/plEiTkMWAFgLqsenyYEHBv8pI1ovB3ccOdAVkgS662OTQ5z8
Y9YyZfWWvSGfR3UbHMytgkPr8uNqN4RviK5M8roB0lEHl0T2gL7fpx0BxSpggfHQX1Rm2VH1l24n
AVqy65OLhY22LW18e0Ehkcm6msEY3rZ3FBiN4PVPz3X8LpcaeZG0o8+jaZjPXqxJGt9sdQNntu6c
vm+NRjss3USHIoM9vbdEQsrENOfol8LEbYWAA/+f72nieZu9rD2kNZg6890GvvxJnwt90O8mtmN8
Z1OUmC0AZjJ5km7ODuVkHfID6OjX1hv7ZPBjnbeyDbTbHfKBmJa+PI5VR1X+qrOC+u+IeX9P0nze
Ly7+SseTYaUnvdagIFRX8fK5SfILEExmeXZh8KB0JvyEFw7QtOA3HiZBDbyh0DP+dPQi3SW5r71z
xNLWQ5NbVEVxY301FAzfyjlybzTWhvOj9wTausv2l7iz1ErxBbGtr94u6rrG00CSExRmWetGAQyF
vZM0XVRdufWMEERcnyIcxDJhcSkw15ddOhngfmvwQlzo3ezdlC7r0gH8DGEPMNojasjZyXbv9lve
DkO9p2DFHq2ooly91im9i516bJyyN5S98DZsxXNsElT/S0Fj9R/opOXd8AkePuSATuYzjpMEk2AB
OlL7xTyD9IDhdyQGqiYX82yJ+WR/eYAVU9AMKEnJLwcDla9Keb9245pgQJqkq9MOkdG+7JCHcxdS
mzWjmwJaSnZMMS6IpC/Wq+KVrItaDqmg+dZD646zFiaU2AirIUgsyX3JdFOqTN2P5rVvRkiS+9pH
v4Ncb/0jLj64Wbmg2Ni4bO24SauxRJRaPZmhM6zJqP7q5ENCWOEZK1W/irv3h5UBydKUdc/rFrNy
TXZx20qW/zs2lgabdgEGveAhi4xrLkgFIwRwJA/vxOzx2agNFmZZHGTrJqq2dTat8jLh+oBJ55Qf
Ldm/cEZH34Rmk9mjW/mmYegULFoMUp8IR5B15LPrKCPJh3ivHAhTEqEwencgiwyazC+xxpl5yYB4
kvp6x3pMYbEOfFM1i7u5wdEjDBpYCAEbRP1e+akyxShlwJa20cyM1HOYDQSqUYCb40yzR+SiTgaN
r56fmtnfWN0WddCT6+702iLodk/wHwxUOV3EriAwR8cwruNNUxA+2eVmiVtd0sNz3zKgpB1PE1O6
L3SjjRtbPhPjNxCDF10dS6kNc8Ql9wmCTjv/gkz8rxLUVA4tJ5qLesMPFxbDL+jlLQaBroMY5snx
hra1RzQoo3s6a+21JvLhb1eTKwszyYXR4HEoJTvQQ7NJ5SshIr7f2cbwpPE+hS4dafcKe2ZfXgmq
eTHEfh/RyNtdBzM7HHVCaLmF+cPkvOaMFbb3SxaZSDPfY0AH5/zlQw7V8GGQCNzUkto80rtcfJtM
Uh1BfQwQ3HavPm5ONoRbfK5/h6o+xTZMdNf2bToeFoZ2hte3lJ5Lg7Hm/ygiDLTo2ubaIU9PEGiY
S6nRvDIbrbDM4oyhkV2tSY2UituEfNNeGKHmKej4aerr0OMgcyJNsQKROg9LgpoTq7Ht62TozkDX
FyFa8G3WV1hG8UPjfbIhneTWuubaqC+c+/o1LF2qcJ14kvPWFKEZDPI9zIgxxafwc6Sa+FWKDDMY
hJ2TDPpDdDcuXF51uTFwZuRLxra24guNJFMw5Ygp+ilIjwizuUAV6341Hl08btMYePxs2AKB20LA
WSyPStHafFSg32rVyDHwLiLN7DfdIIGP+15SuqVJmT7MKePSVpGAsc98Y7QvY6w9g0ExIu4ZiODq
2hPHQNlZUKYWwGLdz/r7mC0zjuAchSGJvOQncmwE6n0xUxhTQCtO7pGTTzRDrFHzbKR1ok52hyuk
+7BZhTYMeaHFa4XGjLOov89DFkXa5fIdqjwfqigvDXOaCQwDNEpJ7xM/pQVbFe8aUC4qj2evMEgb
+T8m4kIxFS171FZO7jBW+EOdHpYDXweth6A8MiJ2h5SzmLZgfHxXqBkoVURdlgHJjA2FhW8XxGKh
4k6G5IA6SS+IMjB8pwzh+SxBgKwvZv6dJTOabVuJnXJUEwxT939/qS7rwd0O1kf+v8LqOCRX1RuU
tkR6HtOg4Js/ydGazMaXcBjA39TqBEpkd9oxoBPzInwVZ8DgxGVmHwRZCHcE9RvY/zlUCFvo8OZq
wgwrzOjz8qHxdxzIfzCw2xPowLsEkBXx45Lv+i6kvLrZEpOfYsVg+yOOtKCsnXXY1P4cRvoo/U8t
lEY5FjQYNoICWIXaKsjCoQYzAxWltYFD2izWlm7L2yvy28ygU/MYuJ/OgnBntC2Z1R6SwA4UTi7r
6KVOZ77+FYMb4/9l8f0BbzmltNDlNOMvo5ughZMqt471ILjOw4zsK7/TbZ+fSi0dOOIZzYlbQv7r
xJdrjJp6Ztspsk/YWJ/OtmpdJuRKK+/ijLSOdBcIIFOjvH33mjeiBlDiZmdTv/gQTLuRME23kQZA
952zpN8RrVGkF11EUViVvEEiG+VouyjHcMS1QWKSN8vTyQx9cSNN/rkO2KcNPnQ+U8XkQb9Gc0Ib
J380c6LQYaRxYxqs3j4S08k9rnFwHJhKkm1VIvKVh+WkcrZWtK9NuEkGc2RFfxMEssb9QzMIKT1m
vudn3Zbo8V6/Qi55CrBWV70hqo5Bi8XHjY4fCieV8TrXmm6Tz7EcqF0i/ad9WXPRE9q27hg81u1g
BeUhNY3RXbZEa3iXEY3Tp8yYahoJfjclae3KIWj00zHHWtqpyLfyqr7Umb2qGAzSQ8mHux15+Vd/
C0jStSNkjb0ocHNpt7pzOw06GXKaMVS5+BMlRMrsz6IbwrgEyZ5ox3uDUQvM8qq4UkVXHyqLFGtE
VRC+dZPL/ecXW5TB+RcITb52mfrTNNLpN/RHOpEvr9pcQtG4rmPN1MTG6KVZBQqP7apFpZth0kil
TNe1hyXOycYB+oIS226BgvLkky39sf7gm21+pr32nzAZaziJqmPQxqAGYT+prVBx2lxtm3LTZqkr
NDAZyllbvQmYBACaSCSufk7dhoKgYj2bQfRjiI/6alb1RcJp0h6XRT7UHOteRCi589HSYgO8g3ul
cg+M01wl9SGRZCfvjRCRQE9lT/rYPkpbWP2ExaWhtmRPCkfZTMTjHRkarcagd1v2/h7Kk0YbmXuH
eXbpxO0fqdD1RivkxckR53pCQidc2itgjMl2GBy4HRgTRKfzc13ZeP8uhsEEPpF+PTY7Bgr7bRHm
dVU/w3QKFaC8ufZY7GHljtRid/4RBUM/lns9cByT14Dd7g826daBSCq8cmephG5kdCd90y531D8J
DVTH8nVsDqUOUE9d9i1hHooMFkt3GJMWB9MpnijHWZSoXjnbjdJj+j4jIcwECQCPVLekxFWzSLEW
C10SYk+6/ZV9vNVX4kxPCWUuKJz++FsacNqMLva91lm8k0uoX87bOX4BcmQJOfPlIoZJylfhTUes
jqADnxyvUjKQafOkfNt7QCyPceSORkwRYAXIcCvF8FoaeKBFbUQRC1wlJAgVS4YSKe5uE4qMdPmL
0m3bkoiRkOyaOboI6UU8upogKowsuEC42DeGgQwAxQ19VjJdgRXSiLWluqpD1lPTNMTUixuY0EA/
5fKfH4pRtMRIVmISchM0aKtmkDHcsxFI1I/GPwpsjKvdOA8xKZ3IrbB+LdMNkpAXfzZH745695oS
gXKLpCGOHW2z3MIzxhEnS+nyI0EHdTXBd98Rv0ZDdSKPrAyz/gApY+BzgvtJzDKGX3nzebItWL06
CTaPPA31qBZpiLuDDQ9GxZZGm9rkc3GuSHkRA25bb08z6h7opig22T5XSZJAfQ6HJN03xUth3YkD
qQ942N7kjAxpSRQLPGn2DN3oyVOhG49OJnA9Y/Ka8hO4R1eVvIvJrvaCKf1rjjEtsEHYo62wt/gR
B/DMOy4uK7hu07auGcfuco7JMdUZMnjKWdJyXpqKLE4Hcymug8HSoBkhUQWpR87zNUgDJLB8nZqo
/xp0dJHGndCBemkL+TO4pLabQUEl1fwO8QVYpbNZ2MG+Fit+0MpYeWdTcYlNR6aFP9AEqRTwtyGq
PM9OmQ555ukK3Bjp1cT0uGWzwd5mlUavrsnc4ABPH1LyQkZ2DNSqbwpXliNk7muM/aVNH/a/WgTU
QUTZwAc5LxIp1TFaxF6YzMd+8jw2VCDwkK8juJMeN2C6KX5lmDIqBwbhQ8GBuYcJtookt9IUEIXR
zk+EeeGN/5TYqcwdcIRONsyLrJ8uLassIlH68GHDA9cMDp1Rv2p6Fxn0YTuUp6hkn4/7/O1E6NOd
rXuuzYrkPPRrzTw2jjEIo5KbPApMHe1AK3eECLw32y0YM2Bd9nONwrZ8XR+JVhb/ucQDu2DcdBPt
tfCHFmvtFB5+8q6UjCm/aP+FDJc8VwhjXzy62a32p9lmtaSQTTQtojmVN8B/OtkynqKNQRM1eKtU
RGRK6NGdPl86A2ufE/6LvBS9FZE67rpuKC1SVpGjjZFOhesEwdzCfQ+b0hN+X6rjKaoNMZY0EcVs
LjpXt+xm9mMoqdQBdspGNrGzcmfZPsARIqEi3kJaXQoKN0HKnvpmVjxCXrb+eq1mDxuOGMLWVbbw
GWv+F6iU7w5ra/67HPHQXnPGxDJ9XEsU7kjoPCuRK6Z0tpyKygTeyAbv1DzI67G+eWR0JHQ0kOjM
FZAnj9Ho/mvXMQNTSLy0QN/ZJr4H9gKJjmL+Kv9+G60nSkhz/dMKznpOs2/KMO2z601vmqq0NPyI
9AvIz1aHFgKFJLsBN9frtSASHQmSeb/OxHbpxMu26Qz5aqMEWE70zFmtgW75q4G9qQubkc+jHu9O
byr2hgfSmnT+wLDKex4QA5cxjfLNdGj762EH7Ax0XO7W+/N4xLItVurDCixAR+X7ZxsN79r5cfAp
V9UzOThuxnG2qMNBIKUPP5xceTFGozE8NxrnxitlwhQiDOop+1DCDS1W02dXZZVQqaAtwait2XDK
94M9c8YZuWI7gMgLElC4ezqQ6XKe9HjHd9fHH+uL6poVTx9NP7BYhW30Dt0rogqfs+fBqFOkVRjZ
XYbs4SFIoaeWbpiOsFgcdUXxIjlW34gc+NtFeAaFm7D0vL9rmyYuSDP3zWmPTfx8d2vtEv2O1jq0
iQT2bErsUzXtUQX6YbJSXmKqmQCoz1JqGOXhhgMuWrReJG2NiRu0Ha/BbygMmgd6n+0ePfhR+28C
mMI9hSSkNY7F5mRsBX/u+hgFsz9wAJQXCZ5aTxNtM5wc0mnow5f/KUXPtKx/DoZjLkkc08fD6JCS
oU6slr0jk48fa2Jdy8HFVEkggB0HBxGfla0mWM3CMDR2L0xN/tw2HJr0LVIKKKx2bmJCZgB5OWFn
iEXnElBYiksRuqsg0vL3q0TSHUodWzF6tCuK89HZVEEnEvTruQyU6kH8ZFCc280mg/kjRn0FAZA5
tZ6l/7e+biIEjABp0THVI5cXXxPlqkSTsZ4ccm4ZJTbFjXNtExmXz+KWWf8yh4l57A83JD2slHtI
CqmSBZ2fjpF+kVWLna3mN9/5bkBRzBZuooafmEaVv4fnysn82zLFJz0O1fDze7tSnaCb5ubQhbXF
4JPth7/tDf0W3t44JsFsAR2fmO433T7YxOSN3KZ23gw457jkxLuW1bL0pS9MROXKQLKnb4GZ5+6R
UW3WyjHk5TA8YTQtsOvO4CVGCsxmyiBU9vKQdWJqlcIsCUAfRlhtssk/iFX+Ba/7RhECr0FsAqAn
xf49+fObOynxURkEwSLxa5ag1woBRk4ATdOyPz6Ht3cnpP+T7T2yitMPrvitL4X+4nuEAWh+AZ0b
OSVBL5Sdo0TGtChRtNR0JvMhu6kNdpctOkYoMFQfFATdQ/jm0g4uIj1PME0u6j27lPhz814XkpYQ
RebTX345KR2FM20w14JJqKZbruMRmfm8MHQ06PZBR5wIPp6cF5jMSPxL0IdK0DiCWyqerhRROrXv
Q3OiCbDt2V3fVspY375oxN+01ckI3JTxXCX0itjr+cBk8klEdOBRf3tjYnsmNBJEbSSkCor72S1y
1x8G/iZF4rT5dOJy5gIzfobsCTbnoiGhg0VYiIs2JjIksnyjgZ0rR7O6dKg+0tLY9KyEgaTkX58I
yb6irJ05p2ao04N02cXEPerifj+koS+av4EqPTzksdSatEcUnPFoxRyE6XVY38Z1x7QWlMtBksEk
Jcgj4O5bxKUluhYiN50cjIgoM/3SkvEJourhpQsLQ8N71kpmL6jN85bFCun3s4cj4kWhhwAlT+iV
nf9YnACeAr5uLGbRD9ROnJTikTvoBpw++UwNXzQqibWnFd78rWEMiQj9BTaGu2twP7GoQkw0k+0l
N/2F+6ZH+W9JvPSSs+8wTB5MQUifjdcFYCNP8bYtALimXIfWGd3QmTgDAeR0t0dtBscNvzwAuIrI
3o4H4EgksALTq8Yh0FA/XkNK2AabW+GDbhRWgXtVC1bQQ1W0RbgJ5Mv8LhbAQen8UPrZiYNlMOQM
qe1KzZzGezt0zEnazdrKa+Ux0HkyOXm0YWMflfPRqasRt/Qp1Rc7HPKczG3hTIBDq5+idL3HuqqM
Q31yIgm779vYRuK2PfRu/8KK1DGc7Qhn8H84J7o1CpcveuPuFmVuWOUszFAvmSk7HLv8Hx3bv35d
xx9TrarB2EY8HFYbxrqDBIyJXouS5fAZ2isQqKhnXFmEKnwuzBdrRMpvnQwVCkzqNWU6GNFp6Zqr
wyQFT91jRAkmNZOtpMXdjQUjC27Ehv4rCPHA+7D73XSGjjMyq3tFYFfikk2K3duvQD8IIIOnQzTd
/mV89LcQ3KxVisPT8de4KrS4P6nwM1AgbS19qzIBRA93f7MQ1CoKvqq4K51fXjmedwGPDyhSZv8D
253V9zqll8f1qpCfYdUkN56JOFxT93hKz73lZdI9ox3rpTTsDKj5+QoSVVXf/jMV8BegmroWbr6+
f7UbOyl2lwbfukHjkSRmfrCku5Bzq5Uf+zotMDtCbgJVuitmTwNA+NdDzhaNBM0KXAeDrm6DNW0q
ZJxZWAMqG+nq0snc2QWcBjLGuYJU9VCz+YO4s8FFBVx9G07VjC3DLEZcPWwSnSlZnKJ7s/PorMYc
YaeyfXRgudooOdaiodZAmuzSmYqWiEzKb/4UAHkTseWQ7NeGY9Zh4ApLK1k9czeIiNAN3rmjhS07
YL5VIv/P+czx90lSwBCzWQuwMF2j+zwzC+S0PFVo0ml2hW9wx3k2smLkW6WJ8Nw1yIH/hIqfxyGp
FQ1dv1WJeFZOZmWbWP25LoWaGD8UmO/a13B7b88sE2XYVKjt2vUtGiO1IFhS8GZQC70N/D+UZyAM
XiNqeABd8wrKSQmk4TNhjEjR84xZaCxnb/T6L1aKMtaxvcNL56jEGAI8Ge/5xg0qagIE5Rxbkcez
KdENN5cM23FQ+dR2Xs4Vh4IhwF25mA2eCi8FvR2rO5TWMNrmDH9PETntoeeVVrxyhyv7TtwfsS+A
Pjb20qwFu272Nhmk7w7+yjtFSHpgn3FitYI+e95DidwLEnOGi7Gn5z2cQ3Y4VStndM5ioMeHfhyR
H+tbPNHkEA5YmOp8nJkT1ojAu5Xz1aGmLfo6/hUq+krdjafDqqBdYgb48nMUwglV+ify7IXHx6A0
mYmnm3QU80Cd90fmzXlQHb91A9bCNssFGaOl7SwBzNUnKyRehYdk03XuFlIBd3SGkMtHt5Z7rrYS
oPPHZg81MDWl0vokwEp0SXrqHqmDzPFn0jZmao4BXCZqUp1V7Qlb5j4wp/Tcudtdgrlc4ZB3fAAF
uc4kuQFLXoUoJjCHS4Y5/VF6XfprpgUI9/M3ZfbRjX6sA1CVGa2ox/VdTQPtaU/XyJ/yxeMVTAJq
kDwe0LtIn44uwgnWEWBiz203ZWlSfKFxRZ3iD5ULiSkY8aYmjQfXQsHQS+xk8ZS7ACPqIZ2Nmlfa
rYyiLayKWv4ZPAGmxnlfLgasQGJqDjHBpCfo3c46jH85uQg9aaqiQyCu3LguvBghlqPMsYoCb/IF
ENLHdENu6CiP14Wk5XJtiM9dBfC2ZItYWNteZBCoCWswHXR7CYOHxuB0KsJrngZhsS1gaGRh7p6m
EPXyVN1sEAwX8YDwKSOBLUoMzLMZNxivLUN62Lv5p42O+5XjoJ/5yviFgTP+hKo5+f/su8i05RTb
bHSTaKdZC9vTUIumcFKD2rL1GU8NoDqkZINV0RNnncZWh4BFXo3C/4J6yFfn0EL7MEtMEIdzv56E
sILDGz13b29jlIcYNbLLw+X0I/g2moKU1GBi6KFgAzAxewnWUfKTF29VN77TfQRCBXyuvweReKHT
ftxHhUkksx3f7krxVTzq7NSaPf1qk6iikJ9ya3BYR65NlsZoJI9PV+GRjdGdss50aVUiLMnZRXe8
6II0jHh9V9yrWFnat5bYq8ZGqAwcDOHoorJBnxp/+7irt8BrXohbcEyuT/m6wc9yv5sRt+s6uUlH
GmreG9xBF5bQDJSroMDhhvOgZ1CPYfuiqhTQQi1JSyAs0x0Tgau9D37XI2L4p06b+aactUXN9nLH
LNqifa2C13tVMhZ7RBU5nivz99wk0iayyIbR3tVLrV04mY7bpPGRAVuW5ix4wESXrZ84qFUvRCne
hASB1kPgwess2NCyPDicfxdDJntCp53ev5VybKj61vhTOoP/lUxatmn4UI8OTDFBtjaRFPz2YJuj
NQT8gSjKCP8h7Me0GOsGHq3ftlrRTYSdhxp+h4ZJyVtcrfzcJM5WWNdLIUoXN6jK1bs0rSaI6OSG
2axGqGbsVSWAifhuNLNvbRSuA6RTBxtCQtvzGVPUr01bkn4S2EgZ5cYskj6MGo582WnkBYVjbhfM
7GpfUv4Nwh3JJUzMp31d3R8Eln39xt8eL497yQwdEgvH0J9Zkk/qjJEcOkQdt3dE0MrtScwjRoQp
WCSM4i5oKD+f5CVueVaql9ZJXpJ5cT9tDTtrzwoM1cdiT77B0yI8PApzm56V7cCX9/r42mmgB8jn
uA3wW3D4MGSN2J5yIuImDgX9vlpHOqPXW5wvhUBonn5w+y5EtvgTrVDhklXNZnQp4lYKNjk1DHyX
nfWDvADKRzAtQ20fqAJshRyJTQvhQlakwcdulZEACSpwYbrL1lbSO3CmQBX5rqJ4yIXPLEvCovDV
DMWcumtNfZB2hrgGggIttx6yRYMU4hDia7wixDYe/qIo3tOWTE/cBV01+0Avl09IrHPiuXO+2lvC
6V/JgK5uGypVdNVPAPVNqpx1RDMHa7CPaYO04x4vLU0ReQKU2fgwys/HMmjPY6+uKobImd2xL3Hx
MJQ5BmeVOi/iYY6KYgtqMO4GQs3eFIFmTCGdrxPUSnUZPJGzgCWviQCerj70wEnS2p3M/8J1ccV2
+qiFa5GBNjc3yECozjGxNTRk4IceQELRT19yYR9MVRm9FGEzBX1TaAQ7MGTCPXf/z1Ze3tuc3emU
2JyPginHhQVrSJP9Lf5epthnMsRKjMYKJzGqvQrZOPtpXD60ChfuahsofJ36SNBf6OCviDHNQDr4
JnYkenwG3KN4Bjkbo2sJd2HAOUVewq7SE0qixVzjpNASHUya90AQR5YqNg0Im0f4xFDNBLkCI5U3
dZlpPeTK9wd2PfMAhcphbc5Frf43sEV8Y1GUPkuF+e6G6Xr0yzQKClC5xZytNLhF/sSu6cHw8e8a
6RjZygHUZKLvIpDOSboodVI0dZX3mH0hUBWFtzQl8dtMmC+AzOdUF2W9kX7oRDiHw3oi7styWex4
HYr+3d2pOpHYJT1XVYVMFNYZKvx/JTewUx/jvzxhmxvde8OB3QRwr8Rzd91sbW8FeZ0pzK86BfDn
+ZzuFI6D0iHuEjqTg3eMhcafDz7wCMIU3aAjsgQa1b+IGNIf5IduYaT+r/qzzAsOUirx+8NaFbVE
rmNUjaTMc1ebNcC64BodIXmBQTyii7loIO/KxB3fHbquDUf6ogIF4q8UYIjmmIRMwycubu1b7yWc
5AseO8wSqM96ILi6f0GbSsU4eomVd5LjaVKXzgJMjd2TQX8mzfPQELmhV2ZuC0Hm5Umcp6wvWjnQ
WGfxcwVu9n4ul2t8ODMfCBhcxs687LnOTpY8BPrszJlUNQLYPfkdMDMEM/jeNfz3XV32zkMb4tn1
KJdOvkHyGdFixlGfPGEmphKq6oZ+tSUk7tt+GpeXf4NeOU1zjMmBXwWUCOAc9tgd2LZZcPlTzUco
mr9pmxtx0bmQDAc1pcwvutG01X1zonv8EpknVY9NMTjaV7Q0aHc9gvD1U2OAH1AmoKhoMhkqk9Wc
uY2PxMzyb786Tt1V9O9L3DdU/27SXB/kisZFQ3V4zxFbw4t687+DWAg0PgPT5prl1vcLCXoKfRvc
Lkc7BJTNc3kNId4EfbW2pAQKPAOWQ4TTCxTaPGu4rsqJxe5NLcTfpGAc9oGpkyId5vp1NKpCXbZv
dXE4mlOsLtqqXeMnRUux4nvHaNutFW/vl0TwwrZ0hAuabEdYHhCYqYrp09o/Az5LvKg8XimYHmk9
ohTblqphyvU7jh1SQKN3M6z4hYTiQ4swzmj5Ob3HYYuFN7sflvzFBX0K7Dd15MpfzGlFf2lmGcUm
d2STFF/LFlvkpLYk9unofWl67MBtafBgeN9xnEOSMG1YknnhO8IEMWn2mK2z6JFcpFhIHOe8Txw6
4+CpjwuQTegHt4208T9UlD9viAgL6iXCoyDPJzsKsv5wYEqrd+o2IIyM610rahDEBanLnd4MXQS1
towzhZt4rMjunf2cZl5rm2xJbJSE1jV462xcaSYuJaC/5KTL2IsMlEgqYOoK/wGXlQr2/3b9c6es
YekBuceFw73ebCbpzA2M9/+hDByO3ul2KBPYAb73xO2msdSV1By6o4dyMtqiUmIJYPRNMBfs8FdC
K7Gw1Z7yNyMgJwUmX1A45sqLiIxqj8lxswkgOHx6OGu5Gr4+XNSkAW8z1fcYbCle6SrE5MtAPOx4
xZY+UVUUQf8YcidZCt1VfXr+lvV+RnB2Z2hLr3Nc8c9atqJbJnQ+K+OoNg/u2voDwpCihRE8tiSI
wodbArFtLfhq17Md60x5K/kr9l4oaO0+2gb+4G9AG6JTwOWwx4RdrYs3VgRwocDhvuEOEa/9Hocw
pTQdQ4c31PlXUzMjgNy/kg62k7WujFf7T9AuAgbmYlPBWyzn1ZnD67xVSBvK81Mjb0mNsqV6UwuJ
2m9xlTQVeKU7D+EP9DG1C5BHeUfQjDLc7pM0q2vQGLjHvSRjrRavvytvgdG1BEZiTJO7gLUSHq/6
gbO4khbxkxIlu9wWq1S4r1c7uzdRF/DzrKNQ9TrOxUSrRuKAk7gAz64kIy70tFnkZsCbVu6vFQ3p
CQHVIouu+iCVyr+JEgDdb/AGvdhCvI9MYQt0obiz2lzoVlixKGE1JoXmsRngRKH09vtygMg5Wsub
lPxDUlOlAEcQbTggxMjdREsEzIYmn10NZ1abM0gDxkVWzwZs0ev436Z7FhqIIetvsn1Ql7qAfw3r
zeFg88XfUx4FFwClhcP9fwwb554QDVdRJjmCW4froZKm3rOjiJqQ3urxZ2q+cFRekvUJrDyRTj78
aFNebUfdWfJ1UYxj3BUrXxR8xHsyQDfEK3cr6G/dSTh4Ietl5ut78tYaOpVuAPECWDHv1+eGaZ6j
mBzgeqdbYOQMdK2eQvIS0amUylxuCbRCELDBORaphktSQAFbgKE4JnnPXA+P00yTHlvLx2s1xT7D
4iGmtB7uORm9McwM/qCnBaLnxmx9d7Xx7a0hKWuK8yhZDO+twYG5KPUcitCjWL96PAwwxOTtKuQG
SRnO/E7s/2XyYnxVMQBqwhf8UoT9w7h12yI0Ld6bogyzHr3PGlflRK+YQMpUmDT850e3RFWZ/9Id
fqrAMZiETIA9hgiPFssuUD7nUXQlF5t6nAAk4ee/6fpsulXkoJ+5h4u6PzlovqliVDnEyxA1fe29
l+IGksK0sQVOqyYR241KdV2sjen+dDNnmY5ZaYqZg21MFd9gP4Dh6qIcVOCqxIc+tv3rr/dGH9HY
KNE/IQiJUqhWP1WgJgzHOdHcE14BNk6FCI7KUKCWmJrmY8RramMPYUu/VPVMLff1ToSc36yJQx/D
Ilz4sGZLFbIdxvXluBIikB8f2OYGpyvGcOLHRD9jZnOOzXPak8ipe3w2MrSSVwqUn9+YOR3FWzkL
t5Jg8l66wLNJYd7vfnwDH6VwVVFtmhht4uLeKxjX0U4PJ3h8PHoDJFCKFz9HsgkJ1CO1TGBzmhm2
Z1tJlljK7AggNqiIMAxWPBv7HVRVg9dEg2FllIAhbTcBynhgxvpwILJhnyYxHGOm9ybcFexCb6Jj
K7X+lLYzJIs4RHtyhBMsaRgEh9NG+5HWIJDL6hXHkwNLgY18NMNTBTOvP4d2lD5Yb5dq/6dDezsJ
UHsDityazGkTdGlpqYlHiODd+ZYNkxIPdCUhCR0s2Bm9jQoCYT46iofY8lCIeD55vDTVaeb00sQg
PcAcvCJPtFFbAMu8Ju0tWKdRG17oDCHEJCZoUT9TtqPzck8d6Ut+O+sKRd4Zfu0itCAlViL5PTwJ
urj8LBDmVd55jExkPu33tBkqLll+NtGtHoh3lKDZFmgmgHpWD6dmEGwXwyt7QKe+N8uBiVGwgzD0
ey2g/ALmGs0Os+sT4WCPOE87Kmyds55i+Vf5OgXKX0ezl922Ox9wnh/RN9BTzdTSNfi5VlDfk8jk
202D3rLNdqaAvbSUH88T0AJuElsf0mr+uHc6pJ9XBbhUBjVjCBRquAf6TZ3e701a4eo4ysUvimkJ
ta7DkQgZTpnWgdBokQVnCSsiJOah2DH59j4zlcPYECTJSXNDpnSpAm2yLESRLYeFwWV6f2bIBI0j
M4//7TaWu92Jy4yJ+WHvuPFMdL4TegtFt/gmGcCpPSDl3mMCTtfqOXK+0Er/2O5lCG6dIMFOK6Y2
xt9qUbKuL9OJISkCHpOql1UKbbsp0vzuF28863Ih66xoqJzswSTLC8cVobEr4btyrzH7RXpyui7d
kdvubBVHZCEyOJ4PJTaZeaoORVu8YWbNejJJruTerGXgDw3Czo1KWao9OTQI6yeVW8UBQsKp6CdB
YO6YoKKPsp3J3w+vFqjFD7tgrqeTSxzmbhxyTQTvi14zba6H0LMxfuZaTP2fKROOw8t3whGliNu1
syJBTaudOmPry2qHM+mUMw58mj+7pVF4ADoZd1MqS/RITmSd+1Wi4vqlYok5pdMzDtX8+fzgC2Lc
nXUsH+fiJ7k9KWjozB7Y4stFSkK3KaSraEASZliJwNB+boTIEEFD+DnBFzRpRN5H376pgbmusHqy
hy/HEuJJLTWmpQAxBBJdZev4b5IWtDuSlr/B1cbzBdsAweexGmeFB1xhcs3Wtg2xpM0xo9kA135y
jQOQphdjN5o6nOzQuKChzSeS6ePC98bsxRpoeN5TObRNN2kQqwl7b1mncGyx30jd+NIC8ChOTp6R
q2eqCaHTvo22bgVB7f/RhwDuk+R6PxU4jPmk59m40GHFnhGbSImPz/Wu62a18H7LC52jqu2C/oIJ
MBp5WR4l7MYpFd+CRA9kVkx37moCsXrCSTLtljL/VCnZmag4bRlq/ofP3kwXP5yEJ3NuSBKyXZk8
6vEr4p9M2DA/Ak2S81XRNQQ6ycpi7lOhcRHT0gSgmCqg4aOWCEifWgquneCp4sHDdh1jvvRQlVa8
Sg1bZx8os7kC7s/bJ9JJVeIKUuoCXbo+16ykjOjjY8K427c5jzijFzjfGmufhC2eUOmo67SEDX5f
nDLHJO9pDLG904e6CXrpteSH7t0NT4uy9HatLhatN7aoE7PedsKpxXLOCa/PNTTGQc+aY5pRVfit
oBWoGK12o+ifAY/+g+gjqresBW61LVaCs54YE/SMvmekX7BdgIP3KkhXAqi9LVD38NgAms+0ruGA
oy2bRWuhgttUJG116RnTyGYyCjwMcNTR1rFZHEFP0Lq0Itkr3OGcNGxz52BBMFVH4lPa+rbap9E+
E4N6fTiAIvo19QofR7aNtuuoXceFpDf4Fy0C2/xRk/JMLO2fYjgNCfBAhz2wlBq31xz2z2M89p8n
1GtO0bQOaZtd0l34cKoXg7+2vvBIYD41fJpYSplolEK3pkTyMf+kcQ6ZB5M7YwFwIoVeTYu8s/M0
MsbScRL1t5p9Q2RWiYQUqcqtrOQodIaE1v+F7cMnYW0Gk0hbHMZ2WjwiXN5p8vPbti9xYAl4iRxi
F2EL0wQx8uwEFeOgIp3I2PH0YKTjeRBZpJuNXIiVeEhXbyEpCZ25kRlm5+XbI9Vq/7+p4EkJXys6
F8804KOlt/1nNBj3LhH13Omqabpx7qz0SMwr+FLqGVfQkmcsQJTIVGA0O9dOE46paJrQyL1mZmnA
XBW4kBLj5zOZ1STukB1Vw5iDvN+BaILmB7binU/wm5+t8CFOoHN95Ed36Ps964DMVyvLIVPiu7jj
PUk+57HIy6cPhGA8GjuwfOr7dCpbpt9j/EeICPIjA1pXU/V6Wo1d9/8ivqwHjnxJVUt/b/6XaoaG
Ge2eWG9HLBaT5CHNlB6e4e1g6FGrnBA+ryws2xxFBdLTYcGsTTKihwNOfJcRYsebQKjAnceJRrA/
QB5yHZkxS0Ytee0okGPZh612/V9A/7rjt1OfXo64Cz4xizZhqFb+weFLS5IK1qXDL9AOcl6a1trQ
i6N63qIVJsZ2Ief74qdv45JlEmkbMkosXUsO3Kk0VE5VIhWrY7s/ywvMZ7v9X0OtvJpzH99aM83U
wfH2KPRZCe6mZl0ktCxse4g2fhDasorKMUWFU4sXgnzTbXOjcl0uMHv8tpNxzhNkIgkuXdHbzJlX
7GnOln/UCTye+zAQNqRbykL2pjlLhbcaai8fYv8RgOm4fV+MnPJfA4avCuuGW+GnwQJzqhMrUe9r
I1ORerUsK9Bif3uExmHJ41UpTBYoRCkVln2bAFt48omtYzykOjyM1JaHg9kpKJY2bvKRs8WCSQE/
1XE8fjtdP4iEDnAd2AE2w0mOJzwUXcgx2rq+8tRXfDKzUf1IL1DLMvDqUzvKjja/fVi8TlR6ILWn
aNzoFQO+7DV7W1vPv6M9nrBpUs377qziPTtWGH8s5s4hptbPYkJfEv9rZT1iXp40LKwVPcl/Syco
e+olS8qy0Meza6LgBcv1t/uxgTYQbpEh3QoWQbTZ/ntsikdGyns/ZCH5w8Zso00hnoB28qZpcQg6
D57ufqajVa6heEimDPcwe0ThpumJJD4af9zuigvL+xigKWjqZdbjJO1fyn5fhHx3jqin8u5HCGG2
IMN+n2N1jT+y74x9JcgVjzPtuZYTzclLZgtRP2oH+OR5em/FDrHDjMvtO3gkgjVVPf0bKM1mdSTX
ReTwro9KMLGwCFNrSZVu9D9hML8Lsq0NH3wnqqYAFeeVaVoFe7ZiPrRKpdDCte2jmiFNmc78WnPj
hZPXxle765uGrfLKo16U4HXy/eYaywXedZuviYDmrzIBkqiGm6sTsrPJU2MoAWZzVJ2c9uTrCJve
gJ6cZBeg3WkGIGHWjQ2V2B1IP31HuVJxrw27dccJ0jZtMvhZw33Wd+0WXb28vrjZwIXvIFaHZJIj
rP9d/k3xZM6ZtZq7t564F32prXx2mGfqgjU0Y9Af5PmNrzIvDBT4PAhZbcWRtU5YFo1Xs3HDef8s
52vITkMIDc6NZcKVZy1tMKsxqpfO7ZwJ+bnNLocOnkacwCzuy7CAONeKv2Z4PpEnQdOLM8xkydJh
17ODA5XoH4P0JybOR+4nchicD65oQaJmQxFogP5+a62E/CTER9PDOVtVHSTLzRxD+e25h1joei4Q
+DmKB+9cu/arzQFpwUiIoEBbKY8iV8SHo/xx7syXp2Z+AphcviQNo2nAFhWn7pkwsDe+t6JcMUO+
1T5qzFeS5hIilrdZRc+RfibbQC7RSE1gXx5WqfR2zxnGoqbXOlszeT37Lrq+GtEe5fpwGWMMiPim
iy/Qk0XzrjSYGJRaR8icoY9UDqgGteUzOxLw2QmYPimmIIEItJpXzA7j1Qi1uvpmZ7pHCJIIxrI3
y8gCeMQos73Uefr4hPkqh11LxB1da04v+vg9zACeU4C3ggM626fyyEBJHuhf3w87qimfacHuGoG7
S4sUpT1RlCjvfWpMK3zMYSVzUchwzRDSUigQtLIbBsWgqzGRnHO40/IR4CPc+06RwH0kBoauJysJ
fUngPZNpXJwyi7xwOiorrribpMda2AdL29uq6D6pSMz+3lM1QuS6veibWnK99RxZTgOQ7d1QATAm
3WKjMwgN2QWO5oiG8je2O8FRvuL75IVLXTrGgIW2cTtNF/WP/JAVgVZwlBNozOZbOaxI7MynScIA
/Eyh6ZScVpIHYe0eu58IOwMu4DC5BGVoUma2QOSJod9+VLpeE+PQQXWFXFX7wobBK9LuxD/9rfuY
dFyf6WZrRklZydNmwTHhHReOP89UuCoBJBGEprh5QXLmzxSLdP4BIIq7Yrn0a/yefgzNIPVQmBae
mavpakWDdzrKH1LPHFcWeLRO/YeeCH1CfU+EfUv+cg0D5gon7VE/eeD5llCs/Twi520C/dkbMf0W
bgL4e95+5t+6/2lV5ssH08nlnDTNMVokyVWrzZgTzOpPgPi1r9HPti2oAzlVWhVCiEy5PQksS2O/
2/bSitdCK2GvRGAWpRqy04atUacpxfKUl8tw2qgf27Hv8wQdCmwWI19cR7knibGWcTl3zFpRIelV
FcdRg1H+ciLlh4f6fdvT2Z+92t41twxv5Fdg1w9n/WmRG/JOaeTGktrNQhh6ccF7CQC3QtE9o1YW
bwVx1LlxGor/nPZOAJozkGctkI1Iagx3E6dO8URI2qErO83zl7unRLFwVCvHgxZZQyCnh6zbl9X5
+Cw3QwVM9p61o+Bt0mgPnunkDybXgEbz8QUVjhALF7i4+p5oFwSwmFlnicE0K3/fRq22O52Mexr4
M882aTS2OBKWkGohw5u1hJGPitXqLMCr5INOr98CAahppMOJDP2zVuL/wdlINLus9UJMIA6dVL03
Fc/EbxEfE4PPDO5phNGEDg4FnohBMmAg3/8TiV8iOzbsWbKDd25L1mCPT4O2uWGp/70DhXx/TDlT
Vk5YzLRmDwUQWp17SsspXe3G6H+GyC+B8L/68qRhSCnkHZpxperx7+CjOrFYtZ0hlbcGjlfVLljJ
Cqe1ZCns5Aa7861po2gNsgVyIQw5dJDnkuuHEHNAAZnIC1EoFzh4FUn8JkWMbIMftbcn18KRC9NY
EeDqUftd5Wzhg4ssKrTCyaN8iQY2qJZVebJRpP3vo8nTYOIuLx7APtkb2pvBvThJ7BKlKetsrksd
46+QycqMSAGd/hUcxvFkhbmvCHHm2JRBq3ojiHCZBX3B6VRjoiCgsmsgB9CDqTjuGM7Pl3fhuUSV
EogVOUVDZQ1Kw+sq7OfUC2aRRLEj0tW1SmjIGm59iU29mCnNDl2MZpvPptrT5X7s+yF+sz6t+Z9Q
pNEbst2W0j+F2vSRvMqzD8iP6SsSdetOFDw6coFrUPsd2NytMpdGnLdVfK/qoYjaGcDcT8bQs+i1
I8NxOeYfJhxv/WyVseNJ1zGz5ACi5SLca/jX1JE97031+aThS+saGczNEOmMh1YsFk1Ggt4Ic+9Q
6iPi0EY6qDSiTB3ERnR+cdB1JxAwUB/9zwh+uQRcvEn5IasqufK+UNx8HhQogeB16tVECa5S0foh
CRvbI/X+QD+SEn0fTWJPEsA8HbDElnJN/IBSGw2UC/QgxlkHstiaoYJeIXK3MSSNXfanjytHq1aA
BSy/nNPSPyd1IfoniMX+Z4fYB+IBm8EtkTkCAwdthfvBT6Ouw3iR24BsVNOQRREwFmiTVagWSNFe
MGAojRsJCfv0bBnXQpk2y01nRPzLslvWXWXp++ZpRSYRTMOBjMpJlM1MZh/LXaIR8W4IdkX0pDoZ
F5A/+P2aEX+cWEXoE3jOa9moVYgCMcDWI7H7Jg83BaCdOKxUEb73wSaHmUoiR79UotvEVHcXzeJj
IiohQPcP76LkgyLR1k0wCnIzhtgAj5bCaZPQzwSws0ucZ5p0QNMzjkhuMHoE9w7GjYi2tyRRURlb
WAwtHTNF72xS2iTQpZqoeWQBngterzceBTYhaRd6Kz90ipZZPF/Ia4Wun5SppDLoWhm62RwtIpHf
WeQM9iUitb4uyocjYfygk4JmX2wL4h+L16UoknXWKxfkOEeZP1yzxBFgmwPdb4oXHgFve42G4+g5
mlsfP4umxOYa/PX153XQ2Yk2Jw9vTUP27nb4x0zcXlQUKNnI/5qsOvStABvATN720vx7uEi5inkB
NtqRetWptu2u6uicrfYLQWg7UVwVzdc0PuLB4w7uN0syYvIXj9r1Lf16bipTOl50awv8UMVC0w+t
73wqZh71P/xXbQ6/QB3ceYIHyCZKs5j0DGMjobulA7+XDwItbz00KFxpeGlyu9zEmypw2xZz9DlP
i6kmnbTch5OIcXqU7ev83dNB5vj8nC8DKwo0qvidwEcJ5xHYcNLT2K2Mj/KeOPr3hTRrfTnc0Eva
Gcv+B9I3Re/Mig7is2Upa3LNqIZZFyY6xupVSwduYoS13uQ2uNxAmFb3oKofe7nEPqfA5NNhC8TC
HHL7BziA4bRiYmuqD2QRGPMAlz8GmLFR0OgQRc+4ESO67pinUNvUzSetcAGgiZzBFjDuwsKhqhGm
tsYyNXV4YezWcF6G0+Font5vo9y774UVVZoCbjfS3FhVxBR68jov43xt8+q1N/BNxNF5cNptn9XV
FkSKihmmk+FcL1UuSqkcKiTt7cQCNgFApkErjpg0Kh9MxLByYVkZBvSq2f1lvUDcLn0UL+0SBHY3
50rg2ATXu8w3X2oD333XPnOkF7yv+ovMsVuMJUXLwtsAUs3SBdN6BJJzmHGTrITRLW/8xTLxSOU1
tmbOyanJakC33x55VCyFbRmwqMGAp6x+oZLX5e1UGl5DDfCzNcU/YnvbFmgsDc87Z1jIUbFBIomU
7t9a9LmPIfx293D1ydiooaGxTd4R+Ntx8YwsxTFdC4maIbY8giHxgSv4BrTadbhSdKwv3DXwBLXK
Y57PI0SAFM/vcAmAMiQ38S1kDoUveqtbqpTgVBp39eaMXyyE9Eqd7SyVOxJQO4RIfTBP1A2l3DOn
HqwOS1Xo67FSxIyap9xSWxT790QAoZgpZrSzHMmSSzWkvESB7WE6D+s/V2Y50TsUS8KKzK1OMw/K
lZgLnJNsJAUF3oMiVEacj7wNWuDFTH3780QBxIF7bCtv8uoGrhBiostjSMQeEkJJKXoPoiERRTHa
YZcqId2oNPg2NpOY893OrcYeKF0zZmHMEqVsIZQcr++5sh3pqEARJ2CUwC/s23Yy4GJrHHj7DdMq
SsewRhu2LpY+0wnZrUrzoD1HwRnfbWbNRr2rpcAnqN0/7lxYdXCnVQUzckub6X04wRzefk8y0RYz
QcXBFlR8AdynticyTyl+vHu8mumJbSczzGJFj2oJIx09yOTrKL8NaFzW7viOqPk3lKSTUyikCDU1
HXXOMQsfqdi1CZut9S6Fs9abwR+jTBdIFbudRnEiu4XNVrCE60LQoNbGUEA/N2qOm/cWGAcVqrHA
s+qih8Qf9g3+jUudPJ1TFsF4H1exKhEueSqotvzmDaFi6GLLRrTf5YlLFutVaxrOrjudRVnFGC00
bZYv7UkBZbuJM/DH3+bXT+EM5GRN+dksrkH5FtMbHtDEXigCI0I78ASSrf+WVMTWF0pNBJSNpgCZ
bWUQreOHz8WGN+nQD1clGccRE1jVUYPrdrET+tUHydBxUILZcvcYpKhEV4XUd7g9BAu1G3NGY9Cg
0Hy2a8fN09q5F+PNQ0vEsBcq5PTxxPRPesWXrb97hZj0tL+2JvK7JSxQLdBVZYVmTPQ9s73Umr5T
booa33EACMZVUgjdtLqtgSWL+RThmK/wmM+CmqOpFwORIUZnk51TmeN3SAS4ixQYAyt5S+XpY5sU
qnkSncS7bjMrRsjkN7um4ivJK/qCN0Z2iHbGa/1QKIiDVD5Zn96Lx2X3qaCGX03JhpaZDAvUlDK5
XA7hYEu/DifOElVI/fsbhXGfTvxQrgKUtRx2HMwU1/Cbo4mGwsKgxF2FHpfHoeC8j3WZSNFe4VJM
FfYOBZmkijORbQbeowLEKaaiKsHf0cM4EAmsVvogmmwZDZ7BD5sb1WZvxQRNi5HYMQpoaABhF9GE
AFholOHIc70vu56b+gmnlUqhsgFKru0oDY+w755U3T/XmvPTxcryCxDuwpWv/Fly0CHKJYKWK3P/
DwVM2GJBx3Y+VE4XAiHy1wUwUCDmtzOrBweoF9aRnvpHPV7Z6kY3GsZ5zgelBGlNq/Mkwbdc9I8E
71qSSc53f3tfWB2n6uZKV457dD1tWzH7UqpMeJV1QM6QRqOA6+XZeDbVrO6SBhwo2JNC6230ISew
9K5HNYwVLL+qoF0ahfn8B5JvSRvVqFJ90qtBLhy/n6vEacChq3VlmPLIsT7DH3jZmQuo80EyKaty
3GItaTgE/gs/w3E0bacrO2MH1xr6iGM+45kzTIsWxc2Abiu0pEpm2x7PSb+cDynkqlLGAShB+QaK
fkg3IDYvdD431UivJh7QDH8QQPB8lkwhjQZV/lnAz+SWxj2RN2GfiAPIBH6XGrkZgbPdxMioEUNe
pwNJvaOQvn1wLhKe/vqYu4TwtqzSIqvtzkW1qdWAzvBzPd7vTi5JHrDBEb3/KEtBk/83JjaV83v1
r6aebyMMnsWPFMwhC/wpKNQsFdVCMujdal4HbLlSGi3IwWczSQs7XTIQpgHSopwlQUV/AaCYLckP
EpAghYOGa1bNc8Q19zyybe6SwGgHQ4Lvb1tJrcCkMQPuSOFkLQCE3eMe64/Zwa4JJOmxmKMHWlhR
GmPQ8NxEKp2yJeexnSnrhYfP19g4HbiUYXrXa9ai1UcKJPwTW0WhobrPcLvLQeYXhsk7GhHxGGug
yLZmsyctzaZXZLgLcxWE9oX6VYWksAPYKCDAv3S3AbcxkremzY7NotwBzUo/NL5igmde2O0N8pxL
VmTqwMDUDzaGO5TT1y6ZdVjbIIRdz9fWhZuInFSUJN5Yib13ZeMBlboRJhCr0gSMYmpV11k2naq9
A4RFQt3zCJkvAESGq01LmweE8jYV9xhm9nfqxkx3l9VwKnTYdCNgWkqSgjkgxfZsYXwwDIxAjZIC
ZzFBqz9N7oLo1rNx3wHAotuvZGyFUbWM//BSpwVLsOxcHrAkreM48fJWveM/7rSqVFL6p3FIO/12
ccMaJ2QQuvSUgyeX4WFpt0ON+UOeB19iRgz1z08SOMmTKTqnfByDpD+ehpDWpJVaSR/9ODcC1EPM
OTaoToHv5gRLCltlVkfSKMcG1M1Vu0JRuZK2qWXkSrOkMRQa3Gk3aMGVuBPFgE6z84oyOLTX//j1
FG6E2TDIErult0CnnRMUwhM7LnNCeIRj5Vvk4gsMzIqcUZX3Yfk+DdaWLjuRY9Ou3IroYAnLPCxU
1nn/cgIeeYPpFYvu1QqbKQel+GBcZWR84ZAHqJ3sk12JTogGPFn1EHApjSZ4ZhaEwqvmSbEpGo4i
qEOchfWp+KNKGsOEyZnrmbF66+8hDdnxr6XX1dVJoIqu5iKk86ImfAqDsObfdXpIZgzNdmJhx/18
I7az8R6c5UkrEg61CmghJMstsK6+pCetHIJKOA586TXZ6DyzA/agW+7xvh+KsduDhUsDmX4AWbqY
kuX1LaP3coAgf4Hj0jhNH4nLxsi3mHCJpvdqt6FvGR7VRDgJ0GHUv9z5qBJfvp2ypX0CFLG6NRMZ
lwzd+g+nz+33S6/bfouQokdYaF4HJkZUfUFfV/K1IpxP/fksJDdCVP6yoCJGqyllutAvfM4BNH2k
cp5Ut7ACyGUL2WH4OHQMZHdpwk5/mC27JhqllH7G+lCfgppVke+HADB8vZbPtcPwWXWdE3KPzAio
FhCbFxVASXLEHJHrQ/u7cQvXK5JtGJb8Oxg6MS5Avkk+JeY8x7d+rxgsy1A3FDrGPo2+gOazLLhR
0aJQboH/2wZRYHQllI1LHEsJz5ai3PMoEdkSyYQxB2J6Q9JZW7TYfP0GbT49itX8OHs6mv2I+umc
X8XsbjTnPsP1Ok2Vt10nQ1UyFAZ+vWTZOwTDhTmRNEgSQLECFtJvzRTUUXNZRbd5Dn5Ph7b56M9c
POunfI+4t4GA5KT6ds4QmBqKPphKeTVdnno0p4UvPW2qIlrwL0NX8H++ciwMWuhctYq+NM7adH/D
usVaMznd+jWiWKCAaKzFDhS+L3RXUMS8bz2GonoXz2tjokZq+fyBAFFPmmgl91K2NPA34Xc9VD+S
2Ycwiv6mzjHlQ109vXDp6dENc6N8qD6ZC368Vngc0rq1MaIaEAlH5ZY4mtSJVoH5L8sVQzRJqi2D
Quwx9uIA9hMrzP2RaOjMmPLHMNc60vPHgzAFmwfSPlgrwAufowVkspJzRAk/eHlwZU8V32QevVnz
TZAo4PLubGsgwbHBMky+qN+WWcf5dEGsqhrmpRMop2PdlQk1el8nVskgs1S+35zQzXtK573wENEb
x1rxlrxBtH+FKl4duuxncU6XLUNPRyFAfj115fMciL+uBfRMd32gZGg7Udm0AJYWKNuxip66nT6C
wWYa1kC7R7n4Zpro4ayzeGvI4yqFRA0KkwyfzBiv3aTAh+UoWwd5gmm32AEppbjkFVmm0JQ0NeGL
5WT2uuZrYE4FNiWeTAAaCdTr62+Iq4KlZVS9zOejj/irYQJTeJIA+vGlwLKIkfYr5IFFBq/B6W1S
W9UCoEl41yhMzqVP+HzLIi+vsvYdkQCkCW/it7cVhR642H9XsXUk/WF4c3TUIbKk1AYnmo5IhaqP
zW0NhC7ugf7Q+f5svawdmXYyexbRWrMaN0fDjR0MRuFz82MxZwf58Ot+Z4QcUt/n0C8qtb7h6q1q
AdI9EJGm8YbCwGHUc/WmGhSIlLQRppYli5z51sJgNeXRx9DXJv7AgR9bVEuslFrp0qL6ROo3/nH0
ZuZ9D5MNf0VBMaXNLUdla6RIaLs9O7GwsUn4kRCbVnLtKtoNtBK4F83fX8LAG7JsaqXdNCYQUaPd
GEmuRZEmOqqi/WTSiA8TRx6DUGxtH0pMhdTQGTZ3dLjdR+iJnoNB4Ks9HM9n9310wsfwViKWa1EO
s0PVb66jdPYz7aPSmsZpiiypJUj1yGT0KHFYKxdtC1FHAtJ/3seH/bpQ4p9HL17tRzn/jWTA1wxe
5VER0Dbed78BZSQQYdpY99jZ1jeXZmnv+2QMe1Tqsf635PPMVBBFFtJnPpJcJn2UlYfb0J2zt57x
d491fFvGwV4TMmvqfqKcgomep3+aUpivPiFub/RwbCWa0G8/HBnuXEc6C9Zjhe6BZ+VvL/cu5twx
CZeQPAoNFD4XUSONYl+PR/1ex3zJMj09/qyyjmupAPKV08pNRDfafOX9MDHkTibYKdSg3zgqOV36
Imdno+oeLVG8P8NorFWMBqwxjmZpZzz70tn8i4llDyQsyv8qNUUKOpISbbw8BWTclwt4pMYkBRKd
ES4iiMbfHuiVwmEDQ2FY4S3tbgzwJf9rA62p1+uyihfWn8sS5Z+2XOdwyF3dU1OJREDiVTzjJlxR
keQLufknaMlYdHqC19xjpMwK/5drMsazVHOK5wbS5i4TdITcEYWwQ44XXkyhN8saJyhvgmU/cujW
uw+ItfUXClTMn6U0xXM/FBoXsF2IakHjVGEZVjEK8GxeC/zXaM156kVhmzaLG90ncvJuZkAwww4E
H7PU7gxDXw/9nSGTOU4QrR0kkV1xXSpgrgdOdhqR2RkEp/71sgLH3Eck2YOiwfW063eJgHLARJbK
vQz3lVS68jrEJWIJA2VYvT7BKYChmcsdkrhYV+hI0E1lLkMjcBohI2vhzmJW8Ty3E1taCRHQR2Sy
TRT0cfI0Si2H0YtQPgbGZyPqKnqWu+kSgT4fhpkWKlAfMIMjs/vx7LBmpLZg25a26+JeGykcI7pt
gjhG10R02YxpflSLgKgibqwVqgRFgD1wlMsO2BEtBbnVIG+NlCXB+GiOb/Wmi9kdqjlVWLY8g6Zk
lnGjckvQWgsihzKJWA+zMdPg93wt20jQVwOZIoE1jE5k+LXXuJmTzgxrh3zA8jsYadRRSml12bH3
Xk/NkoGeuVSKikaYgBgDiQJkM1VO4L4TiRD/cHh+sOu3MzVt26UErjHywMKk8XMbHZEQfalbdBaU
dHctOkWvUA8tqJmzzWa5DM86EO5u033sS3NqhdJsPXdaD5QPbO4DAA777iE2RwDPPSMVsEXzWpMR
hZq4O897t35c0M0S/4H+en2vCLm6DG5XDYj5/ZG717QY9WHIrMnHVD1OuoIDLwR/Tf5ei5kQjbeK
Rtlfw8SLsdWs6YoYnPrzshyKgvlWs0SZyjtu1vZd9mPU8olUyADTObuUCYqx5qZMcmUNLE96dX2t
1nPQFH0Qb5YTYEKAr0ZOMjL9NJfAdd2SRbP39XSeCmoetjEqOJQY1C6IfRFizBBfcWKw9aYo7dGF
OupBEZgvR4Bebt0okjl9r8arnxcR8QKhO2vAYSGayWaa6OTrhr4CNBf/WwBq43M+rKZmt3md7YcO
m9IM2HheAx7Ug2i+yOTDqhjDT2v3XhYFV9NjEv10C93WbvV/nnb1TKsT1f8MN85REBqI7WomScyg
yjLsW/H69NgzpcqLDb0VUNqKtuqDtOK/2hnyxSZrFjB/MLbsjwSZxsvk/fYEjqFmMmDMXJxOukQK
nfVHUE1HPJB53ukansgep/tpKXIiYYAZ8LhQXUAEh0xehTn+fA9xySgvdK+coU0lEur9WL3Q2DrB
/ufaExVeINckVosMLI3MXMKSgTBWavc8bFg0oFDZh+gNUySQeB6/HQsKgwIGSmru5yHbgfedKP6t
vNLA8+NLIOUBXYkHgyWiLkqLARVPQdvWQ8LMBikkW0gSm9xxGQOfnIi28JYMIrS4xbZlAQoPr5WX
plsNMs0X3xlQgRn1EDmKcpzoTU/pldvpoeEMzw0pua9DvsGArG49vFtjZ8E6roP8AtOJ5QmwIAeO
n5XPGK6kkO59ye35OPTlGWKLkNK3HhUwmEYLUahJGRLx9hFiJSmLkZnzaLetsQMV1Kt97kHliG5U
oyiIr/Cnnj6yJfhr/KLnAvb6hg2VYvzruc/06ZXXnBNAzPTJk/VYWtYtVgdY0PrbK9x3Md3H9rxo
x0rAzZY9+Nux2yjMO12WEYFlP99cYeOVE0pnbKUCNwO5CxVzkeSUUHZ9PShOEAKuxALwXrTI6sdA
Q7h05e82mD3QyK0pJv07yoCMP8M2kI1ej/idq2XVnei2o043KkHZ5JnjZto0eXaL7M9BNCcZlk/N
xaqewXMpIMBsuUfodfTUejNK0KKy1Cmh+A77Qba+YZEYAEOqTwWc9TTviyBCkowlvkoVFclq1Epc
CZcvnzPMi5A73HOmOgE46XtdrjfvA1nImolym00BRVJgp2BUZrGx1A9M4LVwsSWKeso+rrNW/Nd9
lIJ2+dFHhTye8YMZQAb46xq6Qanq5jhXHWD9D/lMsl3Pf6dGVBFqZf/pf5Q8Ko+VWjFrls9MsTxg
PWhZJ5AvRCvLhYO79x4Fx50IXTX7dNsSFv5qCvY7fwngVrRS27qQJYzh299JmYVRoXGOZD3AUrZg
uEoOnNNDWGXcLSCAPSJG/gFXEH66C7IXEby9P+IGnu+wP2a3heJHs8w75uZMMFm0GlYBQYlRpmOn
QjceAG135lgxFcchKJahAF9I2BXi4wgRqdYFoT81JPnScOPG80BtBCJI1NO8B97ygnv69GRR5JDl
CcMR6ZiZtqmPs8n0FXFllNSQ3N9HHrezslANYw3/LA1/1KcMlaFL+PLRVefCnFL6kUo27nN3eA3g
S4dfYKE0XSC53Zk/xZtlxI3CUnrqzBhc6VzikIx9ngtZfainRqP7FXDHv/9+bZ8FsJ58RO2z//fi
BUKrPnQcctFIfCrgQSbOGgK87MteCKD0MUXFB+QusIKJCV2EIx5uUnVAiXpad32WrzykBdHSKH0I
0NU8eR6XJbJdyA/X2T5S21kBc1muaLtN5s0RosKTD8iAM7OcwtQmcBbclJOGsy6XeOPbknZj/O5D
PZlveW4JMDlIiozX7D1WOdPvW7ic8p6OLiLFdrp5ARt5OGF6r97BruNLtmKzGdOrvPnHVwVI/Rg+
8T7zssh3jClNhc6yAB96n+7Xw8iTUXBacLB+NpXZoiQ7P2KiBhygdydRmfwC1v8qOXOVeM0DU8DP
tfPFh9hAC/tk2GZWDTEq9q3wGgefdjQcw6p9bSJ5IYNiuqu6NSjwJDM4l3q2j1NN/yMenChtk1Q0
pAeTtXD2fYQxg48IezQ5ZqjcI4lea1Oj6Q3LIk2YfeOFknpzMnOeo6EeJl3FgmI1naGVHunz9QiO
8w64wIC7s0aKEmYTxyaErsoCv91mf4HIHJh4lzyqVCaF6KCc6sjHfQgriDFtxzNi5DHK/RrxWDcY
W6t3cfpWWYcDNGyCm0vMqlrmcayT5Ouq2piKEwx7sMGOWn9i/oNWapzUI34FfRloURbUQQuZEanR
NdahZ0V433MwG+agHNQhrK4mRl6Jdw03xoLHRixprWeeoRKUytGys8gCg7rjWVoqjj0OQstAIssd
ZtjW5UDecNjTDNNBQNBBh3at1bk8m0Vwq4E1h2QCZ9bRZ373Ac1oKYW9kr9cG/6v/Oe1YvcfeVk3
uA5xkeVK4dlpYHHyWMW4eShmsil5XDcZ+yUwa2ywbR/eeiNgJCl3OG2Ue46AmAG/TGtzGk6L30N0
IpEgwuXY1eB6fI4kgXI6k19zWdNuVAsLVHza/Rw+olZbMhVSZ17hBT/C5IPB/SI6lttspxb/EdWF
lS57/tKHSrzj08bvMKOSV+EKrxtasDaZk13dmUP5ZkjCNyxcR3CK5QByGMK/0l2o6XRO6gnvCyXP
x1dK3mFKCSvpM/HJbsdB/mQWeDCC49LE3b+2hHxqEN8RY3ATK3Bh16nyHG+ynumwo2X4REYsJNle
2ySG3RyVoq6Mdm9e5kARYTVt1E4dHgNGCS/KjQjajw/eqFIg6yjiNNr2GyWInAfoyvhbyxNpyu5D
Z66BKSlbH1gKJmRmhPzvmj2ocyhcYwy/wBMACPEjrIrxGBnWIyOgpiTjK8gmkBfUR8RqO8YjPrfZ
WcydT59z2hkt0hWZ1h5FVXtxP2n6VbWknSHaUC+VtJB1kGsx4IUdBXpOPORK3yc5/kG8NsOI3O/j
lGj9ytYh9zjWWRrMGUZrBEkXntcG0DVAcXyTCe2fSSA4M5GTAYeslkZllmdM1dARAFbahjDI0awo
PK39hO3hKhrH0Wx9ejpDx7b+YppuIvGABpRdEkBQf5f0IBUYbpqWdT5t0MPGTYdQhaS99ma5wI5X
g/7C3LBS9Zw+zz114qmLCIZII41aVVUWkr4ELJBzE11lnxime1cHVXK/I5os8WXfBqBYR/fKBeG9
uKvxYLbfTS+1+QTtvlbf0neTxIP3DdgeptYYeB4bHJZc9X7Fjl+RwPvs6H55mORNxEcjt2pIfmDG
uwC3CUsL1cL9q+A7DIeolME3cHUrFMI8yXCf44UovNcu7sRz7ttEF3/Pua+qo0I2r1BEsjZBCLzb
qDEZBN2DheTUtD2PQnMIgMpNLRjZC84zJwvPycHUOPgFgrVs/GZH3kVizRBIQfMzRyReDbJY838Y
GhzbaUkp3pjsTSiyU6FnBadtyYUhllUQ3Io1IsBIC+UGNlkDBif6gmL4o3AjqC1qXvw4KLMzrc9m
qjU65FhY8YA3eqF2JPWM+IpX6GRn2iUo+8IlR4cCb+GgtgvOaRUMmDvcOd9wWYE12J2uk9oPtScx
GbII57bjXA3S/5qNmg8goofZxdxz9kDOG2uA4TJmZ4EjAk8rab1gZBumXSkBrIj4SpPPO/8zEgXo
rvjF1OqPaVcxKfktll3hZxVkqo+8qdWk9SJfgY4BmFvWBIYkU4xL1Wn9blWcDmq884Npq4t6CWvx
aNZ4XFWvPH5hRIB6kWHwmvVaxsndS+ixhy+OgQKhsh/BahoBakIr7O8GgDw3vUkK17wCaCZLqs62
Ym3rRInpwy1LKjLHW2lGJ7jWlepQBEItcf4ZJ3yTwjUjmP5B0+3oJIsPHJtLnS61oiiqiX3DtK5R
o+c06xzaFXQT8Sd0sdvX8X4MlO1WWDjuXoLgAr/MMTbDaycMxRRk5FsXQdrR5GAtE9ypYSnX0up3
J8IKdmFmElgldemCw6CgdsFpGd17XjIUAAATcPgVvKNz8I961Y1c1gs7ST3izD63I9lPHrUadIup
Yi8c2arG19FE46Eswy5ZKbmHrb9YA1MuuMgaCx1o3bYCnPN90PS8mvQtGaUlgN7JGGA3RTFr10by
4MGCipHzVv10hsdjvdEye12hvEGR0E/uxo51ModdaKpVD+HTsYzSTc3CbXtqwLOZ/CWfeRlmTe11
+POIUvvQnlSMpQxz+KGdvLRSF1IZq0hdbEkXD2rDrLjWsG4wt6lSdqmVel1+1h1r+39gXy6jGUNp
bg6l1ocGIp6/SeehR5xAv8ZKustkrJSWiIcquQ/8mdUsLCUwjKVWQ6yYcu6XhTRyTU46THEVZRTI
mm5TiG+mjBWq7eSlQT/opTaFwdIh4USNZaDS15Axwmc9I3xkBdScZckw5rWmmxnnl3rQaNBrwX7z
M/4hs8HB3SZFrp+HRltKAtS2JVupugwWBtXTzjqgDVBhI9iAOFWsOW+EgAN0dr7kXHMSfQ+xGoYo
+pAaU9vDBlC09SZ/k7JeWQnCl2Vl0+NCr7WsbLSeCGqPP5E7gcYTBWc9xK4mpJtSdx6BVOT/2afY
edrByufFIj+sklQPhP+0X056hVObpe82SPq6envmfiRLxJRgRlZK8KG7QV/gb3VEzq4ShLntOv23
CFZyd5nzBpFaAxHZMdTtm31YZ9ZP5dGXSyHvGOrE1GvnsytWrcetf7r9lhowysdKVBUoy/FE+jtI
SqjyYHuLUbQBKn/7K4UnDExChQU7M2EAvytYsPgeJikP5oDnsudLxDDTyUBef1yiaUUSOInUQ8gg
IDIo7y0KkSDwexHtRANljZpKDIcCBR9XTejUIS9zsgPx0FMnFB5rZ7K+NKs4gRBrxdGW6l8PFH8S
22VN/CTojnyYRUuMdDMpw6Q15ocYg0Qr/yRBwZ2A4Dw1vs23yGRAErNg6UEnvEP1oB5kpcfQ0+1b
GC43Nq/hp8Fcb1dmf4NHy9Jfk2cak5ZPZ6XiPuHNLkHyMyJcGhJ/GaaP75eswtQ/xUnXhyVpcnnm
UpNxuSYkAckRkUW+TLqINNPb1+MK5XoDy1ILiouifV8+65IlPZ/1Tt99P5fe7ep4d2wH8Mf40qCW
uX0U0GkLg3TzcDm7xK2bp0b35hBF+uzdKASfDobfKGZA3ODXcQSw2UFu1n6l42zSyK6nKPSb8TvJ
WXYYRUeinU/VTlaUZeB3+POG++94YuHaA0PAohXSoOcqNXh6+xwAxRIbbmSReO7bCD6eismg4Bkl
BMGYDP/eTsHUkdRGlzvbfDeiNy0G/epnN97rBDC+Tz0OxpZNMzyiv8Ue2F+WGYTVXwPtrMTNs1kF
oPKqaJ/geBO27KZWTBeOG7kocTIw7M5FyUvASjkJFfi5+0p3e9wLxqMyswqdBh1++6t9rJ+j3RHw
CW775gWfnutoul+76RCvkOhraJSDasi8FgLWKhOdn6IScf6JMGSfxfv2389RuqeEYeKUrtz67f1E
I4HQyxJXC63cOLJFRNPZgWVLy70AZC5PlYl/haekPXCsx5Kl2HT5fvjK4F+5QhDpauY5X8Tk3Eh7
8KNdK1e8EYarkN964CYwimCzeyR9BZohbrWJowIWeBCfMA7lThB4IecCBUlUvuy3XGYfxvbED06B
7aYbbvIKdXHlgJ904eCABUGCz18kcaEzSLuukmJOS5e0qR+xCHg5ZRqNBzJJQVs37bc6VqYBqsSp
xLz6TlTL3ELRK5FZRoDVd6/wyVHBl8WNtDaZhXLRMl/Qv49uFXPKBCiTjp6n4mnrnWOxAaXiG3OY
zdM+fc5TWgpl3WdcE4wG/85h8FCMjhQP6ue995AfApOxwpLRNIqFeyWB8T/H0+u+A9S5rVCTxPnK
hIZQbrVrYnsdaQnXdSvSRr2HM/O0JmIdLc1p8lp5HYXG0VEWpH4Du4vgRZI9Y4IEKhXZo0BqJwPL
97mlxTVYtv1vLXcWDeb3usccmUaPXnP4SjiN2VjatHm2cDlq8l8jRMq972cxr8DI+eYXCms/CXs0
gjtwWDOgE6cHkHPKVF7SqQD5bB3epTXIzG4r8zC5S/DXJLQrS8Qij/LxcpiUUll9IoE49IeG08ll
jL8r8RBPfPvhQfX2NBQ9N+CdLpKxgQd/Ad4QxXHAaBk2gnzbG+tHR4CLmbdeF7c2Z3UtgFzFWjl2
m48Z8zPjyVRmxg+FxdZw43dRMTcl529X+KNAmvj0IYBfQmzxykWzbUk6smeD8eg/BgqVScmq9B7h
sQ4EaiECtw9uMFJqNg6NrdJesx9IKakRwP7ij91qcSuvOJnV6n485Nnr0osfJMTRzprZTgXeFFJp
pVBhX6JaqRSEpGdnDpF4RZvkCqs2ZHW+zMUGGF4jJDqK8F3pUNkmlGFzJcwe6aDj/6pm+0oMg3ER
N79J4hf98UvtJACwQmGKEnLuT4rLtABG8o2ErVFSP7l9/NvxT0S/LeRqe/ErCmkhNSwSFBF1P6kc
M83PbD8HNin2mN+KPmNyltSBWTw/UKyECt0QTZUNebvXDfjVkN9u+XhFUu6RojH56xYuwZ1MTAsO
5aHzQ715tdfvCba2AemWgj94zF6ElvJARB42IUcjxcQ+tb3nV8YneeHM1DYqe58xw4+IaTh8yMXS
eBclZv8SL3nz7Uc5mewdADUCvUiIv1b++AcBnbOd5Elnnsl/WH6ZQvZY7cjLjxZUTLmPM8EJ6UDg
D8u3++DX58EjDkt7HCojmv0vuGO57+HXheHVo1BIkuumHX50i1NNlu1jhmZ55c+hSNK3SSeJl7Ao
Lql2fRJVaQuEjVaqX2S360hezS/bl2WrVGu0ymIulUlMvGa6byI5QCEIuo6HsWf17+oeiXDv0igt
1qqwJfyFrDFQ3DmXqhZ7hhZaD7R/0S3j87jkIvu/nK0rvoxYrZXZVDwJFM/0HHs4pviWuHGIk4Gf
OasNnwDgVI9krDdpgXcJQd3JGdKzU/U1vM9lXo+Mg9Xu+Cu5ycUcow8saBnsEyItpsp1HI9moj0E
+VE3tXrBjPlv1mFMW7TTM/G/JJE607dgVfID8nZ3MALqFDtSf48rwEmkTXVtoZC+AQAZxqugbfOU
nfnMhAd4eZWCjZA5Y+PGNf/dxESFX1uXAdRQGELZiboI/9rxrN+XrEsf7sd155ERtWJg0Jp29Qul
ptgjHQOlS+xE7QWL0Dx7OkzkQiINqyUFr9s7kK+5hCNFIPFPYn1MmkKhV1+d1z6P/ZlLcE4I3xo0
Yo6gg0INXTl9Y+lRuyfD3dASB2B6ylhtYRggotStdnF7sWe7FJx+flP0FFP/2VLQUT3IwP/nHirt
KoAO+Da7Hx6jt/h47XB3pH7U8EZKG/wEEsHZeTmLcolfRoe4LWeMP689+MvpJ/yJcK2XMn/OR1/L
mtnjFLg+G8sLp6ox/3jJirIdL6ACLt9q8OiYjSTYf7GrtQ9LGMwB6vCVEoWVEGYgkGyuJ0/w4ORc
LG1BRmH9DFqNRCrozOQSq+I4qoazXxUtu/TCgik856bjRsCJIpXqG93h8gFBNLkEilZG57L7bu1z
EW38/7EIynB6QQwj32JgP+zSb8XVk93fwrCZksFteFberoR0EY4GtJWzRv4zJHD5ThfW6wx0n8Ly
4sB+W8Q06n55svgNQYeYcVoAB0A4cHGOqo0Va/ffU3lOO+f/RmZ6TnB/6YO6S+zd+FFOMSh0TiIs
peqfP/lG1wXAxHzQlNffhrK69+iYOR3L4Ajw8JS3vB2pHB9lwd8JNYVCd8uMS6rlwURjuWKNoaMV
Hbcb6o9fcJxpCVE/bj6JG8OJjz5O+qtB8fEWvcSWD3h2mlMqojDQwHY6rlQgH2gQrddc9LBL5mBC
I11BQpvCP1Y+uTwgTg+9zwRwEJObFV76dUBwfiNf+qnGfZQRMmTR1OmD7GhN0oSGj+yaGN6QkzK6
rN6qlEitWTnH5DE8oXnzxXxVhamcNenl0ek2LL6FoDWp+1ESYf810prYCkfqfTg0HBleDIx8vtdo
PHNegIH5VX5mVYSyQfpfdRqTIFFW7d6heWX37jFJfPwFl1FJGCPnKk3w31PXQcXjdQJjj/sKlSCi
CAfCZJge9UIW9vyglmZfVnx38UDtHaJlko3CKjBa15NnXlaI72eEl/wITHtiwnfwjtWvf6OQf6iC
QlUMYMyEeg7ntQvnZ7Cu1+g4ar/Be96btQlbrsFWzW2F5psbSvu2KKyBFmypRkPT7EgocTbibrVe
vg+XMaCpLlKgdb/DuOvZ6hevedX9LKRybUsDwGaJlRpkzL0nVWvby8zqX1lQu8dIjiJrxUU/xGxb
6/Xv+tnasqvIpw0LqQM16t1bSy2SwZ+Zsr1RvMUdBBvWjpevRmfHAxKC/X/TYeHIGDOOtkQijgrz
ifsQpYq4RJ8yrGDxvJQv55wkvCiInG3xEXevtvdTe0xKY4l1oFICM7vtvPYyhbaKhlsJ9Vxuk0Xj
jTMo5M0BeqX9CbiRRoKN2Mi8WJXaVxBaMpLpTq3obyymhxvayECZpUbc2BefjR4BlYb/larqOZCi
1aFKkDDJqURl1Rk86IveZhxO33wx29cMvQqAYvBHTV/C9RA/zfDtnSKTkd52liV+hGGoDd5EgvyI
L0lVGUNmbawahuY0T7Ij5l5S8gcgwIh0EqfxKar7xubO6oWwCm1ORGx7GMDBxMQZgmiFdimN7jbR
9dM8b6lD91Vpo8b/AtsHsd92YrV5ZvyR2pnivmvK3/HT5Cw8o/0QI9jd9vWTTHTac3lVUmBi173e
C3fq21ssixjfD59zZG/1f6yCJxfPU1ghHJf/oHO8jInMUcoCKUn/KesOKSs9ew1CvmNAB6C2JfGp
lvifryaBqAATgPAm58ChXl0RAWXyb1EbqP6bNGmcM/bBRBRsgKgiIKngaCP8pMqJ//FoPQ13edF8
ICvY4s7atY9LEqQBVKDXb9lGLFyYp1MNoCSyoJYAwVY136DIxJmCbf+P9/bR6NpnsSjoHOdYyr+H
XO10fRF3dWynWzheuw7WyJdcINu/8PG00UGLtYAb9FyAURBFuJv4DxZ7daFjFAZpfE1IS5tkEcHB
fX/7w8K9vx/uswb0LKMuuf2SRTSd0xVP6EUonySeTWmezDUFW62lX1aTnxyp4WR/cUycfXb8o2XS
OD8lcxe1JC/eW32MMzMGU6V2hl8/sX1zCNqWKZU1bd8r6DfEHVwsKsuN9wkBIa44k2BWDqzrK61e
phRPvtJlQbIvVQtaLy1Y5KNuvCaR+JjmDVdSo5shL1r99f1WBH6iAF38yrq+U3MyC/XmC5TaUoDa
73j19ZCKaYh9zDpUS6YGRGyHjjESU2XkBpYEB8E8xC2yVL1LGvrF1uVc5vuzbd8TS3wZIKChdYRb
UhBqWB4D0+Gxhq4GczSPEFk5SBhK5rL+UH3O0mTYTF0UlKpgsfV8PNlODh8Y4qPd1UymVb8osNmc
Gfb4Dl1h9+f2hDY3NZQ8hqyHtF29GZWqTjZ9kUsilFfNRPy5c62HOlp6RBQbuRSoJ8ObPyJBwYDn
ZoF5/luBPz2TnKeyYWBLuQMlqMAAzdwEPLCVC0do64/bCJlsbqCPNMsH8oj/xufkvqxPcVV9ulsp
7Sg7x2XHP3cNMjtHjqjRfU9EsjLQKrTW6usJRNA0hLJYImxxV0ZXrIOwpex0+1oQP4nfOhVv25AX
jT9HyM15rlRQPOSkAuAv1U2OhAf2cuVQUPd+SLHeX5cSwXnoGira0L4vXmkUGFWMVZ6ZdT73iCnz
I2ap0kTYwH3ZGBHP3b9rDfTU+c5ToyMpwvxU8j8vuyp76FHJNkT2+EmseXFWmJNYnytTk0vW8R/e
J2yh3exbzkko+8+s5tnpYcvyl7Jsz4iUvnpkTqcmJ8LsaxQYWyGMvA61b8bMZNN7Go0QJmXk3wF4
7I6rDSR1td4j+FTNkkelVHAMmqf87mid58+uNSGK2j+G5SuZ4PKqQWWbQWERfaR8RciwrjK6A2TR
vJZKLbtXvWJQ0hSuiUIltC3Gey96tfiS1XHJ6N6cDeVueBcKP7OUtFXH5MdEC9DafLp7Uvt6Kydy
/Lv5Xe7pzQ4ilauoxhNnaIfr5smWBTxsA5VbXEK3204HEYC3N1yZED28OrmmSkK18w129Pr4EnW1
YfQzkzF7pr+tYiaT5uffxVdBGYcu5VFy9KpZS3okVLQ8+xJ9kd8sVSewUjRc9bIKvy3yVLjIP9LH
OuxlCgkRtaGRDG58amDkgft6M6HP1OexKGrgPVTB0aQgvupYXaaVwa+KnueQTZTw7s8Ix6LlSNSU
VQojGZodbwH7ybFuahcvMxI7LJ0KavrMGbLiDA3PbcyeNaFZRkFe9R190on76bsbTLZBlbUWE6N3
fVPxh7Nm09G5lyk71ZG6Y0pEVjApEUAeSDyGXhP36tTCH1AMAKAiMZh5pokojlLOAF6Zf7RBOyS6
pDmzN3RENYg+URZvjFdEdWi96tmqLGjKtPC1d9oj/U0cblm97MpOJt1NVhed5U6f6Ho5RCSEqCI6
LD6s5LsZz50jOTM54tUlRN6UEzVIesqoNgHdcMA/vVzu/T4unlQELfS93tTZFsCrVxycUExRGBp3
cIN3xAA9ZlRHeLeHSmLWc3yt06B7fOwwSUe2H4papCWHwZYvFCqdS7yOfyn9qXN2gWdECKZS3jIA
kEa0mFHxOIxtc/tRVDnBuwuUaNfIDB1vO1PrH26igIWydxmpM1g+rIia3rx7PrJ5WmkasOdMNQ2/
uJi1BF0nXMor1g3BIeCVOQ9xsXagrHtrr6NKuFRTx3r/O7foLbw40YE+HTTXKdKQF5QM6F/cOySC
T+UTCSljbzJrzNapB2LazIkKSYTXBht8ns1jgAGtUJAOUYG5jdqeab4gNSo2lhRyDQThsbmwo372
ggyZP0V8O4rqQ4C7KQuNRH19PSFpNI4S+LEdeg5/+NjCvbrxqyofR4qByMRjD/ljJP0GJrBWtIf6
L0L6U6/uuvOw9R7NDwtZFb4pWGcqteovqm4LtNu8i7cgwLFsQRL/sMsoErsEhxyvEvGXZVb+8xEI
X5ITo1H0n7Dlh8+s24aZsPdzdJ+2a8o5g5Ga4szCP7Kv4H3pgEjhrEtZeTcGqLKaQeE4y0TnT9in
gBlAZlrzPxzK7t6oftsLDinKPRlA3r2vrslqM3ZsEmJWZEdCtuKWvu800FNB5yc7oyeIMGquMJdD
+p1HQp2SnIyjBUlxHS6xGrd5YlrOQIZgbgiNJERGoKCusZfcE5w/RAloUJK9gIzKaqUv+RAeeSBX
+zdKk4WE7T6PqYo6fQt49QYwGv9AIRNwXMwja4iGId7kv4mIt1i/SsWiyajPBMNmK7e0PuZ6zdSE
OyDwYgisOwVCku7jzWEVItAfKiQYZ6mhW5NUjvUAN9lXtgPfgFPfoxHx483rtPM1m/lt0eENw7WN
l51x5+NbzD4ZejulFLhMei/nZ4gT08XTeXtf8RarBiJLgHIV+Vg1GMcHLA59RZabWgPlwsZsbaVq
nhQvupOwrw9uvnfmw7QALHIyqnDzd44r762ZpNM1v/dz4UfP4ChAFZ0atcClTegZFj5w0G4T6Sn/
djgI6CpoF1t2GfJYfdL+i1tqg4jkquX0S5PR4LmSL2MWDmig63eAzr11e4hY290D29+HszQAJUkN
5+0EVCqQ8XxFIYOyEvclqoAvTYLDxu5VZY/WjFohERtUyJMTElxHpI9PWnqfGiaH35gW2G0sGYge
fQbZT5Z0F/Z1EFf4deNpFuK/ic9IdfAY0WOtojQk/0dHjTAk4/s7g4+ETHnI1jdTWc/nv/j34Pup
NpNlbFGVLyWrRF8t3Dl7X5zVZqqPRITMZNUoApzgsQFH4A9lY5CpA726Beh3eKZwPbVdeYcffnlo
XgajydFVaF5RsvTF9g36dwXCucqfiazGoRXBP6zXyDqTn0Y1yWW59dqY7AKyhsyjz1WhyyqF/2+L
m6qEUcihPolYYs2CnyAA1LPYK0pmBwSPftm1t/B0lc0WV231OVZNmeueTYBBOfj8k6yEhPxmM2rb
08a2zKosPYOf8HrVwbRfFCp6NVSR3zChjqu+mai6qu5n18qr0HJhCDLVo5yp8MRzEI/LI5JJ8TfG
KrB5vnfoaYGfvIjUgRQkJrxGKFJdq7QR0BNjN6GK+km294l8l7EdUR9QZwTeMfRMkkkWtYzNdg/j
8bn7xGb8em0OMMX75aOBPQ2X8DSffw8bk/dGzkh5siQbPWwtQlHiWTcbor+VsP1dRNjFnyOesgSl
vgO961vwxpadw9L06UkphqjZ429FPzxFy1x0oIppqknFkbODAkdZeJpalKkITJ22IhHpq/HnFgmo
ZyEwfH64CfrGoe7m3mszn/9jJejpXOPOMcjw4acImQmOZ5h7wWOD53wXpx/3T/Wp14xtLf2cK9HL
3TMdjkOFK/7LPksBBpNgqq07RLVIXG+7AlCK+eDzjVkgfdju5f0MPsu9ekh2Ssoxount1tw029He
+2QVl7/TAO9mRO5zpvRmkjt60buIpOexdplypYNrWYskbzqDPe4AZzWc4+wANP07+s2E+IzaVaWY
pY9hWfDGtv5K+1wMBGGbAN8QvfjparOIc6Ro2bPSkSClcETnUV44P5e4s02t5J6gwOeWuwybGLIN
jY+mUJkSFxOVzfNBV3WM7D77UqkhR0QfRr4CNCL/qGJU/pSFHiNrqq+jJRN5k9CYZ6pDP1efcf4K
a5Hw+lnyJV+STLhcsh9Zp/FF2iXW8584uhHzDo/5kHHO5Czu3OP1bLxKrdNV5nIHRlF1pSMstBZO
3BRmIMDx7UUevU94vRg6pkI1ipJVAZfZGwQwPExQFt1t9RQ+LsYyvG6dLYu5A2N6fsYas9Y0L33z
ZrrnXhs7XZteu9yy0yMM77Q6BvAUB4AJcMJHRR7pytjQxiicRjzr1mYaz8LpiHJjT/clwIDsMnyt
D2S9pxXQz4ZVWpDhgEqBn/r+ZBQ5d7+CcHBh3sR6dsaXVEBEo3WaGFueii5475dl5gYttQ+MdZyp
97oGvO8Q+SA64BDq2OVprUIEco7FakqXQUdiwaBQ2XCReSDKt4D+O6JbbZX5XhknN0dr0Rq+5lwh
9onwH0hxFHZ5Mq3OO5OPGsRqw7SXgNd2eFdvscUay0nqgQJCkGDfg5hgKbQYSa9CW6jMnsyNID5W
5lxO1YHhUuvb5bz57Wp6N+nsCn1uyNIvVmZtCS8BlfjAKUm6mUy3rMCiVA+nrOmSQYLv/Huv2ou0
lLq+f2pt04jJPZ2BZNR435tZUF10k5vHT1DF/nVHxb2405wvhDsE19NX+YoPWYNwWxZEAUXpJ1jH
2V3AuqZfjXnAbhm1i4Sh+e+Av1cVICNRfczkmSGHKaoMbU29Z4SfVX1F4CmE9Xoz9mzHzf52ReK0
RroOaZBG7s+dT9KAHVW+aEiqL/xes946YthbCtYJf0zuqnVpdO6TlfWhrMwdW71ejGupk1TRRg9o
BP+1WXe7bVU3GFsqtIUrDs5VoHSAdeyudo/2NWggm8fH5Iu32Fk0e3vVN9yEOt+huvwCKRLuz40H
lXzjm1YhL3Lh/8GnO1DIoRlPLLCieJQE1J3HD7gpCEeCtRstCsWsmCPouHM6e5TKVHNFxJJMeQPE
XsMakNbHCQCdOakA5OtuI9hxTUqR+0jhbaccu05NDQz+T4Ea+xnMRIaSYZqwB0dypTiTdfg9ZyN8
21TKpKBN5wFm3QJ70GGYoj2xYf9i8jsm3zh63Sv4TrmYQWKLa9IOv1SRP2atR3EMeX6KW3eHaBV8
NLCH61uV7nhPnRSpaa+/RLCBsOEuksmUfw72bXKpu2668ymDOjy+mcDVLiPFxpK0iuzOXO+h/uie
EbBe2io3lEhpziUxuHvDY6+Y1gE1FZeYe9XTND8rQ7Q6rlqsuqSDJfCvBYWP04Z5F2CoPWziLsHO
HhNiBwHiCa/kAM93jH204Bqm8pUEJtgSKZPWgnuN6MGX6Ipo2OxVxTPQyz5g8UZyeu+XaTUKuoyv
P7mzrZF6aOaPP+ZkN+clr7GRkni2HB6+hIcJHNQljs3Z8NWG6kX2LLRtnW8ZCgE/Ji4kWGk7lGU5
+W19SvCdRyUmc5dvzCiIyWn3/Q0/QJha/Xa7fFfejou0d+4yfxGSe1AMQY+numxr01TxtYHD4t7Y
fdZJQAE4h0R+fQsDAOB258xaS4gf8Jyv80uoC0kyu+KafqBxeGnCvbs6iEShxplaKTtU1pY+EAgJ
rbn7c0kjDpQbhZUYpoNLlfmAkl4FDK2CuGcrYP7d4ihCUpZjhV/jU64gUes5mdeFSEU3HzhwGdCe
Ic8CshKm0nWQ2Yyy+s8N9uTSikY9i99hgXKKp3BTdkrbUrXKiZ6dHQLcmvUmilq/iLZ0ioUm6jA6
asnDXMXum75Z3VL5Zo6qlmdV4TdNdL3DuM3d8k4vUDzHO5J3U/s6Jm+T74cwJ5RafyEgndWQoJBQ
L27k9ZxzdO/tJo1WZ1wwtNGq9iHhtPzGh63rc76bfUG+GuvyslJUwjQarI/vO8WqIrAkmXKKqIIt
shlae3GG94T6Lzon0XCGdvhlPQjJV9hEQJWdSEbviOqjZysWF2GwnOS/RoFJ1VNKj7y9GfUapJyK
LNQpe5m6NK0Jdj0spR48mnIf/I5e7hOMTyTob05RQHSMjmqaiwPBd0KJ2A5EdGBRZjG+1CeKV7a1
ODrHDoHE0jZ9WbXbsaSq/cizncv+RWv5f9o3yRAuggnjloFxLk1UXgtLUb3kOEubJS3FZyNqXGLX
GJGYV57dQK6KiDvt1EPCueHrJlbxH1fOiOnIynlUTqNEA2F8SdIk2kbSYpZbR33UmaITwV8pxtt5
BBVJZ+p5hsGSwWeP3eQU9hYtD68oz70HzIdImo0CGeXAo2hrKQmSPTPeErcCpW7doPA9TkDLLNkO
3uSE2VBmOhWqC8ZQvfqY++QqzntYpnaC+LqBVC40pKySAJHp4Mdc9ZJFAMEiU4gjYs7t8BiNYumX
I+YsD3f1CJYI6I3CF1n6QYxihBHk4VV7WIhL9tALy2aXqZAslVdkTFQF1GnZgwyFgkGHRwJUfL/V
D1VVMZwyCv50F05mfT3a8SmLrM78LJb2Bcdgy/j4px1jOrleGBEu4owuaDcnLChZ677pZ7gIac7g
RnCJDabUNmyUA0ux/XufnW+Iu66Sn1CAGi009S/r6S8OuoLHoQByu+8fMi3q6BiJMlTZyXh7/Djp
94H1ZvNqNr9GMvnn8s+66SeGLrAq5lSeiioIy4KMfSjI/res5g2BoiqV4jUQD6Fc+T5f81y5HYAp
TCCgpA/DXcFRkW5fxrrtzjUYwuKJYf0W3HhaV5Sni1m7BuAvsjXmhPvjzec2OoQBrhJ041XKuKWz
AxHD0lDRJ5K8W8Vb+Ewe/vHihZ09F5H7Pfe+TyozJecpo5bPQtxDlD/16p+xIf6ANpFLBxxkl/zl
CqFw45vA62AFMvM0LxGwJytjIdOTPL8UQdgiERS+JEq8WSFnbmzckNrb0/BboImGMw0gSdrdtXyD
BWtLGiPbQVZIoSGcgsKlEp9qyq8rMa4sojnMMNN5DNzOYjck+F/XLPZHyCN2RuRSSLa0XHnHt8Lo
ZaPrQzWM3mA6rTEBGlQ6VhBoIzONWnvxWqqpZLfKICBz0aKFxZtY+UrtUFeeb0jskQNSjjKQF7VO
G46vCwe98D+JMk5MUvYPFYvdyLVCXcANfH+awypDVYStmAy92DpRaAVp0VHOywbOheQviyjqZ5MK
KvyRqGbp4N0ewIiJJH5Px310tpflYGp4QPPLqyMPmEiABpOFlUYpKQ0t8S53pL/uzHOg0D5/e/tF
cQARQALGPIsuIVB7rTjt1a+Doo2Wdzk6jJFDfN9bCqbTuHEj1kXK3Tr3W3iYgRufhu7Xpdet+1UE
2a6pBa7dpx0TRD6JR+XyYPNPjvAc6HQn1+cZOqBvOB5BQ+VbXagdfzw+/L+ABhuifhoLPGQr5s3j
T3YS0SZPmRBqb5b/JcqE/oP2NOqCxmCWZq/EN5kgcOIzZLI47JL02j05c4Y1fSMGIouqzfYkEEqp
eygL/mWjHWKs9hLpiPSgCRxeJnTZwUXGnVcMEUgounsvgO4ctd8q6BDeQewI1e9ICObGgPVbyZjz
EZgEhuOrJOEjTni+RhZ/P9IS5ujVdNGdAtL/IRDyEhI+8GTWnr7kj6ycMyWSB+TiCuOpOYvf6e3R
Q0Froon4TkHG4UAj+Km+M9ULJVy0WBapmcy9NhVmD2zvgvAY7D/ipJHx4bv1nwlkMoCKFHqe0dgJ
ReZztJbtG8sBzf3zduTRtbLJIoB6+edImYUP5X12IA/P61Bi6hK+2zsJj58KF7a3tpk0uMLAnNZO
+UwbVbnktcMuOm3PkPxjceCT/VzmP47YTtJG1MTelJ7qQDJ6zXwCLOO3UB7pvqZdU1UFdyzlQ59T
Lo1G1UL5w8TvBxuf3Q0n2JuLUEZz8X5TJh3n9xtJQnl2wUwFkCJvNJjLiSZA6yN/Q0pGVUVjDGX6
3IgKfcqqws0Xt0mVnbHzSCg3+LM2yC3PRsLcKfdVElgGHk5MS1fk32ybdNtlBFurJDlDPGDsvKRI
DD3T/qbbrHO0uvLXyci879kDqJn4nW+qQQrAGWHfZNbLMtBWSWMZDWWVaDde/hTo9QPlWN+LDQR3
Q9PNGBWRSGjYQacgC6M6DTXLnC22ShGET6SXp6rsesh+7rIf52HeqSD5lz8qAc7q1LBv+bVTXrPa
cDgEKnYtUkWKL47F674WZkgFHkSqTJZFx2OfMr58orMp9oK7vN75fKMPIqwxmkpNXlEftQNnZYh7
Vq8Rzzy6bFMqyH84QjWc2f9mbTaJTa25f9KdbuUN224zaAeMWASLsYuCmMGSfBS1mqJ6fGiGBEvI
BM0R2KaWv2rnYGpm5yIkyeMbPH6i2SPAiKmD0axzfsisnpSrtyjFMdfPbtIBMtFbWY1XAXEK4HYr
82mB8otS3MiGedSQfyFmCFebG4H0Ga6kEQ1FQSICd33CmFJ19hzAIudgf1cz1rLFDsdwWa5Z/GXh
/zSPVypQhyDqG4QydyTWJQCoWHB3qYkyK5T46MbtDWJANECRTCs36T0JU8sKVBQORVCwTmkCKRlE
mMmIgxR0e8VKTnaKN1Q/slnXOQtFZCXjY2NFbdQxQ+ER8Hcp22lezYmkhbblJmZ1INnalR86m7jL
G8yA0sb7a8CRaaWuyGYzx8FhybFrYgX1vrsyCbDbFIGxEPL+HlbiWsfDPF+6Od7FRyimN9/9a8Sg
FoQKt1GV79EwcrXA10nW9tebS7c5u3dbL0TjytwJdtX95rXKXvgdcfM7OFTRFr6OCSkXZuFlOVOx
lO8IX1020VaFa2GUTZi1rFIL5i8VtfZfDblGdKHZ1VShQR7r1lBgWkaiIxNmpfO7tDLt4odQDBrn
rN4y+sHjPfoCyRrbavFdvASswF48ABiv2qOR4qhwQAutM+lkuZQ0vzDww9eFVWj1WB8QwF4gSs+3
EHjn/4d+d06CjPNdtfAHRfrDmDpx0K3svWCuzUcwx7aVZLUmoBq6hW5Ry/AEOTA76CqjPKJdz7x0
tWwEVdElgJko7gTKUmJkcrP9CqZ802zn2mNOY43K+j0guCKbBmQ/pmI0HEGCeLAqM5Nk2VH46jMf
5ibPqgh9a1gRziyaN1Ai2ZK1QYL4n+ycd5yyEvpabGVT+lZ9QwKnvd9L9qX3iLRF1sBHdmABlS9R
1x0TjJgX6ywszWosldYClapeKK9gMOruExD4PYl8zyDKXxu46IcVDX5znIJt/1P/CUzQpIQIFKsQ
z+4MpoezvsKC5tMpFB1KX1usdBqZhth5K6lUlujc6h7GYWuaEPaKNdmUbPGW44oR4NHv7gDVKDus
xI1D7cQuOv0552v2RvZuFpgmjEL3rC6HCSiPjQf/M0wyNKn/YPjIm3aa0k5QryW98XFDH4w99EvV
17/SKS7ULT1QorYNNY9bJoWE1Nw66TSNrOeCu5OHhE+0/LCBj6m15Oag1AaCnlz75zJSAMcnbV/H
HWiAa7AmpKJnefnC6ntdKgThhXGZZ3DjzZctvmgXtiArrhjeLgCpRn3pBsnmQZ/aZWqGhd4fiz+3
s3ZyQd3utF9ZS7+u+3068PS9a0vmBClGcOjK3aeCqFl0o9EuRLrAaaadSOHKeGgwvlNF9/AIFycl
u+8AjR9XuuvK1r7bdnElm0FC89+2WxJMhNDlbNjnZJhnlCud0Dsy2Gndqk4J+oXcN4v7suZqBMTR
UuUlaPWiRIU9foLiFuFiSv/bXMmuwY94w6fmtxvvljS4HcsCuXQoXQ3laCL97O6UpERjNaadYrnB
0q3GAYd2LFP6LT/P9IpWkk8Rs0a60RaMtCTHTSwIIIQr+PW2z/hGPpybfcQTHNp45dZfXxDQUDIg
oWiCEnSB5B5Q7u1kZqjyRiNHgTUxEkbQFzXBP0AsG3Vvdmq13l/A+62acFbz76FoVsiCxkCytmju
6MSzGytfAlEvBEsPXZxAQ3TxhdcNe/P/20cyf4tIlmno2O5gM6lz9GW9v8EQpOxdPU+U/+fvum7J
QfByhUoYwAh2TfB40fD9B/s8yaXd8JnhPQ0+EsWPm4nrRbG4MYyAgRohR58PUsTiqaj2lY2RDoaA
I3agYziFAAOtWkLsFpV0s5+yTs+72WMW1uPAnTE3P4hjrZcW3yGPr7z2aNLhrrp3wSif+/8mFyR1
PO7MvO5nE1N/Su9OeBShZdtk4Ncrko8XHAsw00kcRpVSkvtrHz/9Gqn2wMjNRzNVx1WFCjIG/orN
YJnRo6WKaWVgIqsInhZ6KSwloSS9n2QaFuzHq9vLq4Xk77JFOiFGsKLWPI46UT1qqgQncYm1YWOp
6oEFFrNlDNUR/B5IWvAMI0oJyT+T5LWYOnfE4mdbwmm4FvCEDxlcUJou8ATs8GBCqegOars9AY6Q
VLoI1McuDyZuw5PLfix979Shf39MhiVRXeKpM7waSL/AVWTMBxP6LSEeD/zsEjBZhaMpdXG43Zxn
6NX/VkORXx91nupy4AffGFIwv+jZb34ucE6nlqEzQwz/WQlaozuCvxpa24eq1rudrlmdBxhxo6Mh
cUDfY3u1aTwx+1M+sHpSIbQzCQBfIm6P3n8QtEa7Hs2jAdl4nK/Wett9QBx8paT6X87YsgnALcO6
dCXOTdVCHDhuSxuJH7vTiUIyc1+FHPjdglgg8U54Fst8CWq9roTZILBjowbYQOUaPZL673PhxQs0
6f6l9uaFqJVr/m5uVeQp6loYwFBch0vIl2bwKJMSe/05xnWpQPe7wSWbnyt6Ac0NfKmHPUSzVxms
GAPupJvJy+EbZiMAFeMTlzWmdxJYGoKcIbeYgo+DOeBHI+8HOTZ3pa9/+IdkPHerdeNCw2aowB7q
gSlcO9OliXNanKMKq9m4W6h2W6nNzpLyJz+p0T60g8go3XI/1o/y51M0t5G/uQaE4jcHxC5HLgjm
pdo9dmiQs+54HgPLd/Mf8kHQfZRgiQuwsQ3m/v0KJw8gSapCcoW7c6VeBbmcxPXebh85Iqd+vqCJ
knYVFjMaBz6g050y0sHEqaLJ/tMba5pD4XPTloB6SmSg9tqGPApqNd5cE1xiliLdX9PX9jntqYsm
CqJLDsE/quE/3W7euUZ3d8xJXIJ4+FpaKt1K8NCNBqKP2xhmEcau20E5rxpKXUf+WHCNgRG7wh9v
qOwrVhx26qrUoNt2vWltDqbihBdcRsLiUI+S/MFzCN4TA5xsFuKRvhMZE2pQDXBdAD61ush4NYpY
bVXlLV2sT9Snq7YS2quRYh+B+wIWd3mBIokjuSc0wcd1/RpZuAvZ5/cdSVZ12O14YNCoZA8SjgIb
J/CtyF+avySwpUAdqM9wDj2Zv6+UKgg5YF/QLEmap5VUuNznlLh7L0xex5AN4bXcx9HNIwPzyiEf
yBX0Mq0KdwRjxt8U+yt/AwfIYK9Y4bHhHYXDg1IvELUISZ74TJZpkQ8Ei1kCdEnc5sNKXL7LCIYV
umP6zedZYQbXTRZe+AXy4/8gCdyrs0fRA54ZCk3jaLaw5/n7CLvRbyeTWUnT+xvlvZzIGjlFhuP5
aByFihT6bJ2zNIO06RjURvcEQsmvo9nIsL+hS9zVFDeE7b23dyWQ3UBcwZmWrJHL7fSuPt6cJGPZ
7HjKkj8xO/s5N68eItVvtFSDvLsj4mPUV2xCHIV70VBmYuljvrzC5IQlx9tJ5o+GX/EIy8t+V6ps
GiSVKjfDWn72eCOae14xPRNcAXnUtOghOLFc9dQ7WB8htKk13bW3/L/hEJXycJY5pCcBosCtC0iO
lRJe8AtUYm5lhVf+NmUvNpVtU34XqPbhknwirWoqe5n+fl3VVt4Kd11UuGxlFskD+ua5I45TMcr4
Tx6dZ8CHFyuuV/zP6vcAg91hSPY4RSINu9/8BLXAwgaTKAFidVY1yj7PrJ6tYiNTY3QbENfBJKuv
XSdvaPU5/VFakDUUxAPQKlGehCx15yhQEIBXlCNLm7Vx0yuv2awJS/bgloKZBiUZcnN6E6lPV74m
ZetEcsbwvxvWjI5dIgGq8Gj9FowPi9rRO9S/fTyLw9ZTjpw8oeHbrYcOvUU4JCnZQ6U74CBBWcPU
wy1tMo4ulgopELSA40LE+xVouy/cLdtYerjMfHzUCyBxfmPjsNVR4oHBlHSKz6OiOo7hzf2G6Mw9
y4zXHijMhanKw8t43cc+xkrL0MS31+DFSGsW0I/9GjCZLssOyl/fY5rLvuvEGbmbJijN+/saWsN4
k/0Kg6+LjR8Mf6W0XXep4TBS2ZLrrini1Dyt3BVZLN+o92h+zTQsVODw1Dnj6ITaMnpSs/KGTGOj
IhhNdl5R/2+lppc6h+lIB6eFlalMlm1BtXQ4vX5SzXxIWsjl58dhMUWa68Ig8N/AI8JmH/gK5s5d
tOr8Tz1fXcI8b6eUMe1wyFQCtvRnJAFu79gvNweWXT/cVtYN5arCasil5a7a/aW3zcdGeBzdvs0/
aX0tjC7fjJquWmUuPm7vrPSX3zT+Tt8FAhMRIvg3vKCZ7DZjOkJl+obKIy3PdFsmUKx7HaoIH2vP
FGyXa+aEXoXv87D4iSRMqiXIifpdl8zrL/dGFziuSv6OWFyHKzAiVddGIqASJ+SKVads0lmyIej1
K+jJNeYbtHj0FF2wsG8yzbcpGIJz6rXVzoHXzm061f9rpQRnFhGEXgpTWwmPgigcvLbSNPSs+L//
0ijfAyYPJan0O2gCt1Yd4WMHk1KjgaD6YKqb6wWyNoM7xsjOKUNqXNDgNpLlDoLoiNM9gq9rnkl9
URB/0v0h1GOF066bZfr8PDwism28CH9kplqwTAYdrhr4NbVjpTSyidb+C43a4bibPheSliqzvlVR
CbHDwLnA4P9e/hiefAH9hOx0XgtRDTw8sZryKMl1CMq7qP5CZIZEDub+Rx7e3xPfeph/fQxwwDt4
yBdFvDkVUz9LYL2gMALdU0F6xxwYLS4z/2GYC0h2oNoAqY9C+fFG3uRjYk1qOB8siUBlkSFCDvTV
LRluv4EYp47suW4FFpavClLj6y7kpB1Xv+J+X7junLIqcBL2p+gkePEZ/axP1E7+zXCQLOikKoiI
NRYtb5q1vpXvHcZl1VEqt9ehFnWNzWdnpvfoeGNuMTvRXryT//Yn/c+GPRaQHym/rxSKlwKC8F67
FphUW1Z0gfHwhdomLtxc/hUBbx57fTIBKmtneJYE6FhhmZ24VNUKzE1AkQo/p9S5yJsSGkQLBXn/
Mt0u7FJ4Nu/J6hVNYuCizfWVzyCcnWOziHDy4m1BnJzXuCJdYESVoVjEBRwzAfqqHOBz7v9stGda
Ufrheq032n36lMA9wca+1UjwZQVSYk9GPIiyA+5wh1V05c0M4Lm0wS4xhG/gJXQmL65AkbviYRTq
pqQXUCqEdIz/JlfuApdz7wG3c9MJ+Fk/8QcDzHZL3IFsf7yDofNTlWoXfam4Gjx1mVOEi0fb2tiZ
RjUsP/f03wIMu6zX+Vtbouw8luY7eqZg0DUb928xobeXX/YmrP6YLdNcpILN2jfk8hzwJtanAaLD
5kZhrYYlkuFPscfjxe1NVVHMBuwMorjVkU91Lu21Qj19RIV3IGLjpnAKHXpYrHIkMTSJXVZLP8HV
RqWhdROXwjDz3E28jLbffdKyXMb+fqzhplxkfTnZ9EQXtL0GC8myj8UpBACAoFHM5YO3knKtgkd3
rgI139irqJUWN/s36AnqHmYllVaTr6deQIEJAOhxSXfpHm9VNVZmdpg1Vkoj5XIWqeYKoHzl0bwj
c8Oinj5QC8tXapINNiDs+5bYrZu7D6sfihj6bXJFJEhj6YbNhA7vIvYDoRqzIdyIzAC0pyzMhjWG
2PzKHDWxhdL+slVap/zWl/MWbdDX5PYnHO1eAb73tQJn2V0vN1r/FyFt2JL6hKtv9GDBsf5W+c8Z
gaG2+dHDfi5ar3Va/FaF2cRJHvFOFyAhvEl1ErWK3K3D3zFdtf/xIFLwqHU6iTHRUKTS48rejfxD
yUcpmUiD+mGN6T107WXDpuCAaN/xneN5KNa/1oVwW94fip3osa4ELq6IdrqeZ3HB4oSxXiAFZ1Vj
aOMygMLnTIlQxSs0Zo/LyPrzKLhgMCvoscaGlCRMjkIJcIQhZ7j0MeLbGG7QZgp/lXiWFiPi/Xgh
04VCwHUwoOobrL5jJOMvmZeRby9KSkcqjnFwfS0ytcGrtLJs4183LuJLhzhQZivJguTtI2S2Rv2O
6mA87t4277bA0gH7oZ6NnLcN3UfjhbJWpsadPA71giqjWtnERDlyvno91KvLfJ4pAI9w1k7ICptL
8Rm1X1o1oeKVZFMryaNnIWCS7STOaPbM9ZM3x9hktrLAm8i7nrledm4fIRvnbiPVi7tiP0gHU6Qb
ehca7f/TSLfHCGKY/AmxuztS6BEKLTZLkdae/1O/dejwiYAkm31oedGu9/EvDjKpT5eyF/B28Hyf
c84Z2AX6A7vnCScsJMSXPioZI5f1/QUIVaQlNruadOWeK8wdAWAikS6jrT9cokyx5ajDVffYgCE2
aLzreXTRFg6RMM15ugu9Xmjw+wx8NCCYmof7ST3v1eY1ngqU4mWEiFhmBkrWEP6x67cD3tOYUqt1
MtIoSaftIA3GsXc6odUASUdP944R4MlP2o0WKC7LTeL15yvZKb5UkYlwlIjqH9fuCs6ujbIB7voU
dx97xt8IJ/mviGamgxQjP+puSlZUv6B4N7WGWV+ogT9rlyfP4hiQNa6X8FD0R5lG+uAFdTpD+1Hx
3qLLRIaEKLFEf5Q9DR5mIcPqbtPvNoJnKNNGNJ4WiphZzBq3VxBFTgxm1MhFQt5qd1JZp+/QwaZK
6/0394+wIhK+yJdDR6cMOBjAtRK9VLHYMlvfbJrjGE3I12hQKhQNO0/aPmWcISOVu3xvT9BmJWP9
i9jITOxshKbB5x2As3sxAi+ulHRPGJmOzMugfNEDiA0UXS7AhI/Vlm+ftNFoU/B9bkMDXNJ0S0Mg
UlMXm8FqzfsGpmoXPHrWuG9CfwSsROgHPLyF9XmZeT/7qUqmN2WDZcU6DSdyECp3AtHoGOcVKMHs
pSeFg1cELQY4xaSn5DSgH71BOEzoy5kwK9blOskbmlfoSjS7/ALOBqyVpSBNuM4YNwsCvu0W819B
B93wFz8K5e4nHWNkUPRdgXNsJmhdu2BQ6PYYNS9i49NhEQ3cDjUZgmQOABTnNpnSgVdRC+wH5lfX
Z8DxNskLABLovxF8mWZ4THgYy22DxzaCFFjfslbpdxnqnWYevDPZCMFbtIT7whi3usOig0+F2J0p
LWuFHrI1tU1juaFpsiQ/VpxHDjAgn8ST46wJPzKMk/0vQ92VFOUElf8VmAP3kstfEz6UsLH5cgnq
eI0YpHankqqAdexRk2d5S/Kj8x8DO4xHlDt62o7chNl4hPHRx44CuWudX/2xygenT4lPZSbdQmOU
T9NzmhRNf8CtmW9XyFxCJ8gEy+ADG3aDqmQFIqjnYxbz+LRw2+igIGqMgljjFInt0GibVGBdCE/P
a62hsV/I89tLFf3UtxfW1+IMj9DClp5gKav+z5C4AZIjrs5dEr13c3zc9miuTV2Is34HwOqH5v2j
Yb+zMHLZZtmJxspBPsxpdlLR+gurZzgbpAfBISJXJf0hMRMtpozF/spImNBPV6KXWRzGaVNCfnrb
DTA2RA2T02Z3SvMBY0rQEEam9MCm31Mh9PQCZojXIevvLIAJYivIBZSSqDIL3mBwwABiGCGYmZK4
B7SOk/YVTjfsTl9j5OLKKc3k2JRqDlVEroz+PBRbYKmhwIo9ESzJ2+WJcHPt9NCd2x7UJLNvESg2
cS9YVuX6r7qJunnZ7Szt38RvR2BHOlUQ8pOyY6u/Ds8SMurhQnIZTKTG4VUMQbeHkx1HwaGnS3G0
GjLhxGj+0L6txqmEm7fk/5j48N1CDiWv+lzS117vCzB2LYy1GNCUxgYByX2nqUMzI2REkPDFFlP3
2UhEJ+iP6946nHVnktYB+3uIZmB+kcPSGiJXSnXrpSdFnDqyBmrMcIpHp2KJGvorRnMPLZ5F4J/2
Z3LQ4kwtvdqZq5fDLhBqTr7UES0tRX10ud3eEI+pWtP/Ax4bfaMj0/lXUz9ktbbjXQJry7P154XK
JiaBa722B4nXsKJfUys6ryums0Z1qCis/n/5vlUCQoF5aQ1aCdJrZgEWmr9biP1DsfVMvdyccGYv
dth1xyTKe1rU/6rsH3V45TszlXALkStSNV46H9IcHxxKew8Bod4N1+ikMYLcqvJnoAr4qnhNKlzZ
YYcikBvQx3HgjTmZUPPNUC0fYSERv/khoQNLfqfNMQOmBbnVU63PAmw/vE4rGtQCs1h3cFTBaAcY
RLh9LuCRy/Vsolh9y3kSIq0Gasip/kNYyeii54vbgGZ5FlCtuqIlp0lJtvyZ1byQyE8xJgWs2nLA
fjri2Cb410Iem5VoLgIYloe6GNDGW5JgMvQOgyodSjJsNuBpsmOyAJvMgRvWuoDXW+yF2pT5U28s
qLLMCDrM+Gy3sioaWhZKfKEytME0T82U6CFSabRsLJr584GKgYkr0JRfipDEtbSlZor+ZBEfkttS
omLutWrYcWxW7EsesFvNBvk8b6OnYxKDvUn2XE4dCeTG+PJvRzaCOQk7FjLzhdw65uf1mt0AycP8
LfF8NvfH9fNGJDJYvX+nr9dTqksPtc7+PbfAZORv3Qx6fnxGGesxwWfc7W0GdfKkev7W6wRzSnVa
dJ4168TjJHWNR2OyMPKJ/qtJATBXguB9+Z5s/y6RVz6Oa0oq2ykcDYJnnbsAjHkhkzYwSpD7GqtS
ozQe70rMDFyrP1nRb5bYqrMW3QolZxdqNTqwwPLMkSHKYy2ZNuW17WyTWxLGJjTmTRgNxlVvn5Dm
s9yYhONaAb1lLO3U0f5KFbqUk99tCKsp4UsDQvOwcw+Q81KsOynPjeJFDtG2Be4p8to2nBL/leul
o8msIWfGQ0facD9bU6QwHdrnEZNC9UkUkzQkNip3uykbdk/R/N465X4M/F/Ff6IrnYAXpsCoEYc5
qHCrasQ6fiQ3OxRT7QpDaMK93DulPMZSrr+rXg9mjN1n9oNeAE2qoxaKyVzBRKK9QuCR8vns3TRW
uTajpH44b2wyXug2AQEDdeAawlaw7RGA6Ew9Wpwe1jcf7qYUPoiOR+auR5L3aGpuB8C2G/XUI8UJ
QRHaihLuexXlxsEaQZKXXV6SslRhbA7hYWlofVVLUtmB4j6plPoU71tjttj8fnnisxFDAJLBlLLX
fGKyPVQXS73uRXb1wAi/JQ32smbfR3ohz8C3jBoNyMFyQzOl2b+FLxtVrpZrHurrDcAGCAUPYFBF
gCuh6TTm3ZH7g/IFuttuUzDpie5Ed3G1dvWfd1t0D66XaLEk0KxUqjGguWbW/znglItqBz3IZygs
PcT0ytWUeVfQ5oWJy5S8E3ef7DvP/PavbkXETbNmLI3aYwa1+M3/FnENtzxeuclNroQLiGQpuA+R
GCUfadVN2XvJ6pS9CD+3eWN/F3fK2Y+FpDbC0cHkLNwOrvzuIeC3ihdwpvVsFmoOCkKjNbumJW6s
SwEqIXOCWM2ciPacB4Nb0hZXab8CECqfUuOcT9aABExcYvvRtb7M3/Jr/h2AoE2so0i7betBwjeu
aAPcCbuHPR+w4RGN/S6V1iLtGyQ2Uk68GFFv2sUAV3Fo0x0Xe6clj4VqqnHr5sHGMn6WslRrTI0D
t+o5xh9IlwUTAt8yYj1deFOEYbyg9jLYq2twX1LbMDSQkNXQ2h/c6X+AGwRriPLinOh4Yi5Zz9MR
hfa59d1p1iFF6gRo9ZPDPWDHCVKvs0OWmpvy8N+e3PNI0hQnwJ+4i8vCqQkriN7gjR0BhWWw8S3K
0IRoK4sMbeFoMNHE4qX4XrrHD2K1h2AsSlUT0awex38AlFQl7/fTp5wA3fGdopGWL6u1VcQUgy9S
24TQiTdiXwZkPqH9zJRiwvTtG/uJ+K2gsZTeg6abJ2y+OuXhsS18k6XbKKu00hNKGwgrsyZhkjf4
lxKAoBgJPrZFQqntmeBG8t5x22JuQruUm9hTcPzOBMbgvQLAaHIDLeHOU1uC36KcCOGVpb6JCPXY
p+wEm8xR5qcJ9vEXdkESYaCgy3zpvBIWe7usWevqeLN90BzEy4E2p2HZUGRFspuy5TZMrpku5M4F
UYoH9CMPk5gvtcM7G4BN6xF5OcqPz9qNuVhDa3mL8tTlR4mFUu3aiaND/gOz79as1Pab/cXBlzC8
PfL7PIbRDeg4Init2enwcUTPbp5i0KPS5Bo1C3ri32HeecUmYq07hLufowU8wqx2omK6S1HnFigv
iaDCbmZwbpohp05gZ6+5cmPSMypj7RQc1b+uMDM9MY3dnIE0uuct6ICGgDSCS5P6svyzGsSVkoZn
4VuXgf13rY10zHLODSOhGr5yhQCejkBnhExoTk04Axx+2aGE9Rm3zgtjVVbFV1kJMfWIHJOCAWvg
eBvkZ25g4u8VPvpIxOfB9Tc1WMuVv+XUau/01i1hsK5G22vNVuMHm+aGlUvsyy/Ypc+zLFXS7Fdr
jFG6g0sKiAIUfBLtWCWimXHMQy2KTciYBkQXjYssfYeYCX3SkGO6o3PiC+aDD7/XLHL8MMpWZ6Ej
b3kUehJFXK0coo+eS1OUFZUmttH5aQ8KWJgg85B7Tb4yKZYl/HH2oFA6lPiAkyf/9N6B6ockmpGI
nSh3kwcAxMmjycFTwRTyPXZ3DzbtW8kj8SVbcdNYsnZMY7ORCZrsJuKdaMAPbWSKxESFpx8pkMCr
3XquitkOLqnPzDCxFSAwn9+KjeAROjErj0UhJYtAY3qViH42Cr+GdEz6m1CtyWLIKQTzB26B2Fk9
OIj8kxLxMSHmm0Che3w7latWXVZ0SBEZXW2Mqnvz5FQWlMb3XHEdpBqHM8LswcQNt1SV7OXDrUW9
iPURXYhqZogotcJMYF29AlpUlr/C325wmc1W+rK9LORK4B+Il73PiF/TFxBYEAZZSMOQA29SDb/y
oJ3zJKOY9ZZv1Pq4kcTPWNSYhM5IE2+HPsBAM+6cggPUV6mQp/vWrCnoWInLVYUFgZAlEQMeXXEY
Y8M+N8l5Bv3nm4BeQxDbNBnwn0yhTgovnbEEdYdsHa/RIPV2pJZOaUbcYba3DO98VgXfAOQEeBNq
shzOgtd4foyDC5nBYOlGPLvHjyJT48xCLrBNOy3E95GZho4TtdhhNHcwbKQ6Q4L776DOrO40TbHW
NNzeT4tf6cBjb+fJGPGx5dNXRg1dBNlv1ULwZzFBdGNQt1O5+ihpX/g6bwoWbEINV0Q92YVx98Ar
sbfYdDFwnk/EJEJfMRwl/oylkjnO5BgwSB85b7eUL8XK1aQggSRLIiQELtyRfuCMmMD5Q0uzXNPi
HcsXf9kjAkz1YPxkVirDFZ3+5P3gtTU7l7HCJbE/XmhydDuubdFReMvh5R5PIbvVAhsvGP2sFpDP
IgVCGVNenBeCmmqRBuRiX2+wiU09CGArqoqMnXIyIfmtL1z3V7LRPgluXUlvLl/hvDNkrWMnhOjk
hAvheeCqwA0V8tfodrT6TX7BJ+k7ejOgIM2j+6H8Namgi47OCsRzQ2CxGFSOUSAedNjCWr9f0Q3Y
LtoXQsqEI/BR+otFzHipiIGazzTNc8rKJoHSHFONOBadiJdkqZoh9R+WQLLtCd9ZunhDqDz6sggm
zccwntxHQt0h225cIHORVby8BWYDXPweMa8nNqJErHHeFCi4zGcVUBB9sRcnaGri7ZIhp5FromTk
sbtOU+jNyDWpYOIHD5KqyCAapohLe6ZgOQ6OulyvZkAh5cQ+r7oT7fntwOZPoZCJf606mkjk65H3
QVr0VkWSHPUYoN9XVviGla0NgItMEIG+tZV5oSeVAW5ZgktW3+tKHxd+pfg4Nteb9qsIC0P3XvEm
skcd1WDDVNesHaoRPf+r/erUiCpRA/r58zftta/Q51s3nu9+elzRpTGMkorwCwAkEk0IXYVOVCeo
RCqBsDfFgmQ2ZMpAanIgz723RQDEL94MmE1uSifzETJf0vfnnNIBwtrHKBnkjTJjpMLWfCbGaL1O
vNu/Y8EDnidennEO09krOZ/cH1qSBp/d2kx0iY+xIy5twajm3ALJwVQXNeBBPr5nZnkFRauAnqUy
gFYxCOkk22s+nnOd+s+qKfdFoaf5f0k4tLfZbuPvyb1hriGZTgV1aVRGWD/IYs4gEJxDRimUamIQ
8tgXPlQo8nYpZDFfIVGhU5HN4uDQM4rBMDvY44ENW7YcLX8WQyJ7twuocUaGmIgnAWDjVCb6oUxc
+rDDy/rlN+WNBk/GwT408jGVnaxTza4gct4zByuZoCCFYsME4ge8bxYkobY2T1EIoXFmwu7YdMS8
xhw+X7qDlpW8rZhkMVQs0ZiTSdC+uIx5OfbgG0lB6SmqVQEm9L27t+VAUrsZMzw8bH8wpuIuqjsX
3IeK8kIfBmU0kM+7PNwIGKJc3kGEsbJph6XkX7rel+Wo8tTd5TfQPJ+pJkJdN8RypCbzelvylzin
nZbCSef9ZpFS435ZBJSIjphwd07f5cPTDZGz29zYhtLC198vbc18vc1Mx9KWJ1GYNlcRqiqoFU04
m6XyBRvX/Y5Tgk0l3t7YLCL06k69QqsrUwok4uqSYO4mAgeqYeU7/1FP/hI0fhLa2qGsI+OphtLh
P2CmS69zZDRbgaOxzBRu0R6CiZ25UWFFNp5g/G4zKGQRMbDrCpKI/1V4/jUYtaKKuwYtpwsV/AHR
7/eyFjhPOrqZ6GGVMewkq0TezTdgivGfwGUHD44uRf1zqlBPWop2/yRpxe2YSoex9YwHDWBE0r19
qRiUZLSfWPbi5+GirzoSwsl9cgy8LFgIJsJb8GtjAGqtTQR53zDnCixvB4eaiHhZSzmn+A+gV61S
w013m6843ZdUigL4vytcOznLYJo3irizElciTwGHu2DXqbK0BBbao1W2kVYDZPrDwyt8800QRevD
Z4lLPrWlphOhYynwET5orQj4rmGQ4jJqkrsGFn6z+9M7LHB540hk/SDKYQ4j6ZJLLEzYZGxWfdvx
d/WQSHuBnLy36EfWska3/oE5mcoVl+Tx6/PFESl0AZFKdtKAJ93tAds+fjh73qm9nXJ3SWDlQJ7R
FqiaBMRTPI9jv3RlRi+2KRRkRRqMeKjCPzl5k5NIdZVNlCWMML5UIvl6I6a05yx2E2X7BDrXb7Sb
+v6chkIu9A4vrnUs8fmUIodactswspw0tBjm88WRBcbJbUGvfz5TubcN6v0Gp6Nx2K9s54ci1UKU
C+F/2eC4ezfTAtLBoY7QhjkU0SK3HsTBs8Mi6+Ac3qw4gQXZcxdjVnpC5lPB1bSSGcac6YP9KKEm
W0ii3ukD60HsEp/9lv202+eJl/nYLOWASHDIBDy8VWdgedOkZBpx8eoKlH132+Kz8MaICXqLZ95x
ovR944E18sGOwHBXPkosX5+nO9bqAJdQh+kNQLzmcAjhXtQpbpXrkdXRayibNd577Gqkteh7doDz
Kojb4l/crjYi0gKZ5ZsKYqmkisPJYkQiHi2dLdZ1MYsCWYggG2SWuprOVH+gV4A+ZM9l4IbWJtp6
3omOd9pEgTvA0ewCgQnMjnJCcN6hkYEAKdUL5vJlodIi2TUztPLY2MNshJut8C7CC6nn9kibD9UA
r9R7X6HNVP5RSys92Kf/SUGLNOlU8aIjHKlsrdWM+LagL0J9fSu9tjyGcCsq5MxMZDyfHTDdfmFf
aBbykXPrBziDhBU9vRocYtOV0ZvHyvANN/QHllF4pcO/81u6YjNjgm35yDEmrCDKQ1LJ0BcXw60/
kPZTGl2w9N390hQsHqaFAFL6z4w/c83PjNjS0+udQ28GmM9rgNwSeZORc/AHAVcWULoKsBzQ0DDx
HsmBfU6y5KsGR413OlNyHn6OCdluuzu9+9gG2EQ8y1JJLtcO7xMr/SiLUHlWmpFxwGXs2puCwvd3
5M/5qH4njeV7/VQqHSXOkUzBmA9Urr2uxfDz+2T3X2ztWkyNh1cUfsl36T9H8BKl9i4B2K8GAEZw
NcpW5CyNGQmTjAJp9gWG7lNv2Zmoxv/2lOwhzWbK7UbwgqhHvrCDeSInV2qNBrAC19AVgINySMqp
DyQajagcKSM6lI+A+tP/TM4cofRnPQCcwHZODybKsvJqQHrzN1GGc3+XTRJrB2NOGtAsNjlSob6Z
UtjtRpdk4W5iRb2yFzLLEkD3dOwWXn3snQ09gy4fbLxCsO3jJDgg5vN94O7feE3pjJFLRkBksnUL
OWqVByVlKACrJa7j2VzQhdKGxwcfOqtnZhQlxOBlFnR9obtyioGqEV9foHnAFiUDuslO+dPqkjpI
F7S1QoBHrv6/nYMrkI3IaU3+mR3ElYK02Hen8C3LaWQoKGCK6fyTfzY2k/cw45YBwNGoY5in2mk0
5jyqPVqY2HxvmWyvo1YD6BcUk08gdyim16017ZLQQmIorB/iyy7XlGaEnmIyxrwLJDXpP45dTSXE
MzbE2Fx+kdwcigiTTPXxs6CpWQ7SKwMaFZtFvrzr0Q0tUtKXIsvezyuICpRiBShHpgLvKkHqB42W
e+/hohMZk3Kaj40w6iVkk7NFjA4qpOFYykIjtStlkJVB8xGPsErm5g2+cd0r2xUrUCA1lwDWOugL
z9dJnjkB2KyawaFTMJTwWY+M0rpEbpa1QKq7uhHK/aO4206S/g8GcTNwCjnfqlS5zjTKUcJa733p
EcBQU/NJCWhExQniud6UoAVDdNWQrxtPnczIDwyH5m4ddQ96egx8DuKiob8YytqkwKnHIx+vmGqH
8fVDINonM0u7oMk5vhxVjiQOI3al6WzmGbVT4+aeU8JSlziG8QqJEFnYC3ovFLYYFop/9FncOYyZ
WTNNl6mrPd2sktkSWAKtbhel1DDf8+efDfmvMMovXP6IsWT01itbqzet+Qkw8vLEGxvpwze4V33w
dWMPGjQ2ALu8SdQIMGANbveNk2JvhVAV3Kyzu+vkVXE9hfNlhlm+WFNRKcFbZpwC8w7Ih8Qc7k+o
zGPrdDXkuOt9pKBdGfdDDNpqOvSDFUt1wdkombNpYnOrkSANo/v1GRF123osIInBuTXZgtB+Qeef
gDsFXpid9p6YFNq+usEY7tz8gvTKcQ5FsHHA/BNtmdN8jk1LAtBzc51Ofsch8fANG/n93vg2PA/u
J1NCtbb9mqlx5FjfQ7hz4EOMONwAViGN9tWpTMVrKGgbwBMUbDRQTyQ0WhiQMDatGFksPfO7weIU
4eEtD0L+lpWqRdmO+4YNTBUpeKmQzTR4eBA0LeXW4Ih9k8CBmOmxKWTpTw5IqhWUz4nOr/6oven5
ULkuVnQ5AXZKM7bkP3rj+q97MBzw57xAnkyvatHMJziNWjzunbRGTmD8nSUnRTboBUh4kr6tVifj
crTW2LZ4xPUhPPpZlGiK9jWt18ObjXOQ9f0557RQE43N3+RAQ3SJmqS2dGfxr1qy4HtlrVyE9Vjp
XVj4Giky0eCUEl45eCDDrUbIgZLvwegj81IwBiUo4s2FQJVVBlmuxwnCbpxfohQFR7bC/qFCEX9P
3pZsXBPebWOGvYiXWyjwQdSOCykssaH3DIMJ7+Hr8EXGylrQGArgXgCZY2RS+KBi5Qhzdaz67uyk
qGdQhY+cS3nH4OKnVyjoxJxXSNzhsrk0RyIfUL01+jukd/ZABeO04Rij2fbQJJ00KqIPfAiLV/GW
zbMbhuDv6osyp0ddB4uXaR/z28XIOmFISfHUf+Zdv1XWjvuIj8ijLKN8KyQyhJcdwQFn7cxCAqDz
XVam9Cpgles0+962qgMbUnf89W6eFS6e3FDRHluvHHeLdfKYj34iScs0PmrS6aP8E7SihRQRmxfq
a4gMhBif6P/oxkmu3xnY3n9tBboyCBrnkL9zkZbDXUraROniQyDrXZ0lKS+escg3LxImpg6e2Zgp
tPx1KoErBEbSjofAHkZVLqQYzNvq1pdB/uYML4ywE9zTMoMpYXsRx/p3zc6quMDH0PkTbrhVUElT
H7EeSpKBkjfpclOsRrN+OcKw44pR4OtbmhlvIT5saNkBnvWNG2Rs4Yduan3LYPRWcfkGqHSttN9d
r7vpLfPZpUE69gNH05UQD828lULtrT96P1UhESKHSOQnq95wlmqlKkoSQOD4C2jZl5msX99kuylY
nIBz34cYbr7G6VcgW0tdc3603ll4wHt+aVBjzlZ0Dz34UjG17mJqvWfVqIP2hvn2lvJxKxBA1Mk3
Q4dVKd6FZJWBLmCtWKEAjphb7Qqos+UIunBw6Ag7AMxUvqUtxwQexCaEBXFUIMVWWazglTDz+cx6
kTVv5CZ9BdGOu3YIlLDdOKD4SG5DjGZ4IkH0CU7ArV5Pl7hpxmZx8V34imiAuLRnGhymqA5xl7XD
8GfW5mSKyfo/7Yn9Mt1e4xGMKZ1DrzXVSLVgnzBt3Mua7VymTlikZog8vTcHjH/k6zx+Wv8uCmit
WUGNbeFPKeFup8bZQVwLtEJyf+cLswIJmf0+FnYHQzxwUHxhQm1fwr1Vte65SRts5uakcKNCmv2Z
feVuNRfwYuWplOo5SES0CMzmmfAaFLlMSreA6jtIwytUNu4dccCqAXp6H+eQxf2ntR53txMBOo8P
AxEXosnX8xArw0HS//NnCJRuYr9SkgJgERQOI6zMdyT08gBU2gjRMOKwX+BZIEf9pBR9ZLEk9j0c
vHpGkdHvG5b0YG0PKJGfz1C3xzPJCrsik3OKsGiEeYTmlgYTFITHT++UUnXOPl5ipbFauXhaLmTI
kirvIZ9roRnb81+WZ+UqL1TRTgPWnfPzSCVUF50V3AOifyOotdcJ40u6k6ABxCJPHb1M7eYm5XlV
g75rCuns2Y05IDQfiQgTPsNP/IMLPzjaYSatZhFPQ5N+HFEo7xQDf/ELUnF1a6X77Cji+XTJmBGV
+s0j4/O7EAzr6zBSSCBE+i+sqiJa6ujV0ouo7XPYy1gMnM033FAaPIaH1Wkfe7cAdurJWSVjAsdN
922bPYe8vVj/SjGP1S/HGhjkdd9Fxn4hmdiYSd1gBFryepzD0gY04jcxuCaG1+xDvouB4B0IIMXl
3QtbqboDrXFV5bX0GRsw6LF8Mcy2pB8K2iMsao4wvbSUmaMhxYXU0nf0rfnW84sJNwhhcyWZr49B
tVkDNnIowrI7Sw+vuVQqavykuExawi2j/YQj5MJ9K8W24JsERrsCpKl8DX9tuiCu6ZwPPZD22j6w
6keoXmMySIjY5M/6RMsPsCAcwn2aSas5//0KvV+fFJQaHARrjXQpP1B2BOwTyM0xEGbCPd8TYasv
uwJ8NBY1pGcj8L9KMJcKKmIoDL5U9+799tlxD3/9hP0De0g/h2VGwmenFEi2CGWQd4JqMjZy3TiW
tlVLgQQ6RvxqYJYuIVcUhF2O8jTAx0AbQNvOGNyJgbdvlHh1ew02Dm+DcclsFoiUCP9B5Cmc7qo+
C3o9Zsh0qQskcHri6DxugdH6NpWFncyPNCBGu4nYW+C9g2n05ld1NUlBaTeiV88/3qVqOL5m2xAL
lb+FiJSpZlUt3pEJINtOF+Vn5HSnspiNoVv7jusMzDZFZu62+6js3WgYklUkEtRtQv7QkKDbxz2s
xkQ7o1/iTuAOuBiTmUsruS+6xNO6JfSK8CPWk5Ziz+VeFEQjmHvRwg4/45jyu05zAY1H7B1ZHNQF
n99I6ZO+FxcZL+1gDxeTxEoww56CPSPJ86Z1mVgGLcn2CL0kZHbo+pk94FnKhMFna7MJetzsF8wN
jVrg2pJQYiEHEs+7QW/Yc3Cc69tzCOWi/ugJ3wv7Yda5WQ7ZMCnZ7oljSXZ3U4g/n1YiX9h+Xsa5
4FQ8ivomcvFIFHDlFcXuiIKNYb/xBmLd8s6wFys4niPa5Dldn8rzUAeJbLSpPSSFnSLWURpQ4a0H
JNsWVkjdC6FeITM0trpeJqjx2P+EOVwAhQ56pIuNKB/8eaxOVfLZ7d2imCZEtLAIRHsgCB/Rudw2
XhI4YhG0nEQH/hwteJGXWgHnqR2ZqCRPAeJT3OiCI4rzEcTDTGViHfbgf8XQDV/a2XVqG255Y/z9
iOeM4G2YuapvbuS1Js9OQF0MFfq6R30ouPgIfMfrNDgo6mur3V6FnKxhHi7WX2QP6OFLeFmn/l8p
EPaleE6Mvuf60rvfCBiBKOnMK84kyRkI0qb6vRW5zHGNjb4JxVHOm1SZW0ZACcym52PavHwP4xiG
6oHAOyAPsBmI3uGGON+gmbT8zDL2uE8TFHsNbjSgyi6jVphgIDprs377U0mA4r03GK9r3ZaQoNPl
Xn0/0TMS+NwKi7Eq4fRl0OMm3FwrhCIMq/dljdm+RuUYZusz6H8KRd8q1y02SsVi6kascqC32MSb
QkyebYJW3oGrAnBCyjYIwUrmQImDlkYdWc5DjoFdK3bA4hWPbUcVL2+gwXRXTj5w5V4h/vTDqx57
HnQf0b9F6CCr9ab6MEntaXVJdhSv+mS17Zpzy22bAx2dA9MDWhHBJNuN6y8XvXpBTpBSwnlWYWxv
YuM7q1fZVggYaAhI5Y9KcmXIAMPCYzAkfFXwHpHCT1PbR29+AHQ90D6s0FfHf7rLCe9Py62nUFSP
NxcwzasqGX1JWPHDI6VmJX93qSQuYP3r4zmGek2gl2NAsAXc//id7YsybkUOqSHWsqXpEiTKLvTX
yxR0KHaxgi7uOA4TNrmTdMURoKCkW6CirWTkxuv5htbI6JG5E9zts0XFyi/n85ZV8twnKwDr79l1
Ks7doJLP3d4QJesuQkxxVvehQ/F6b+Gt5el1m3hkE4jLyV+nPFMbcpBTw7+XXcN6XbfHohCy48n3
g+kNhfU8UYZXYFEwIOBoVwi7jeSz+KpTDXrUEuhn/9QgVEv/BAIqvAmRJ5tZjsqHnqzwtLN3RB7C
ktdzpDFxttjbGRKh36fsLVd9OP+8qB8SmmkoulJWeuMcJGesAyw4ed23o8UGu1nmVdLId/OnRfN5
rL0gY4eg+QXLn4Ir3n/z5tTgMvzp/nBnunfTcjAOtAm6Htu13IGgaz6uESnhPk8tJMa04xTlKaXV
9OW+n1eYlnbtl/halcTihd2CZtF/sa5rFlVAVUldgAWrMpYQY9Jwar7/VPnlfJO9DQptfaWT63nK
leVmGi4kNl7FuUq2QMm9SiwrRL015cOAWXKDwMTiqMfFp42U4NDUa4LJzHmK/WttIn08Ho1SQBFW
yX6eDTwruSxsU2AP5vc9ao36pNLX4VA4iwrkrh/BcqVaALNWAO6GmkwkQTk9Lfypxej7TTJa9HMu
NwkkDjDhHVsc4Mxjj9WWV7WjUddpASUP+XcNm/Omp/k4V52MXbmth6GElNOxsOMXcaPfPCuTT6Wa
RuZw0eHrZGO41ieN73+o2ejVjK0KC/wbRrXkxG6p37wOOrdqmCdziSLZHA1W4avdRX9o4pUM/NYe
/LgT1uHcRcQ08TIWabqtQTIRykQAY5fC98A9KajHoqEXrhXgohzbu+NeeYyekJoTYZFvCRa2dkNW
fB6ntCqxW5ROpkNWyKkDkYRGoFVIYVyjr0m5ZDGLM0k2v30OzTDHHS9T9D4qbvyZQNZqzBbE6loi
OeLuo/kG+ukoDUrO7JrSUlrFXnKGbhvyDdXLhE6L9R7dQmh7XjeLCxZsD/pq8ElSB9c06pwrX9Zy
0WWEXQW+YxZ+ND75ITxsh6kNEyuHUUSjr0L96PJhWg2J1zpuPqB7gQQjLddaSg1yQ1wJjmZjRJTV
+BuWw3tZ9aw8ExxO/2tRXCYNfyLrdSVywuLnLK3nJRlMyluriMprzCbM3SI1j6H8mzTinvA7XBGU
iwp8XEou4BeczQc3HNdrd8uTh//3c4cmORhMmwn8rIGqbyO8Ac79zI/Dkgc2BxUhsOtzOUfATEJl
cvXj+IyZzhOUFsR0s9yt0ThmHxPELXnWp5D7frB0mgU6XQcjKk4b8qZz5YVuvNxYV+KySwmh04Sh
zf46FG5rd1KZfir+bHWsBa2VfIJRHcBwS89p/8z7xkStLdGuJcVWQHlKlx2fupZFf7Tv6AVGXiKS
5QsL4FyhotJy8OYuxDWcBdtq2MXj6b+vltgFpOgHQmUu2bhTDKWFPKMoZXhW6RzWOVvzRGHBB3Ue
uRf3ttkzJ5qIEQAE75XTtZzwo8sw+cdxlomBXGtU81uP+yoegX28gtKNkogPq1aN7E90xtKzwPSE
hgctuZSp4X8Vc8vKePvnr/d2Cq9jsJbWJWOvwih9yc6qDKaQ0UTSd5GfNgsZP4+6Ag/gye2ZnSOt
dNOV0u9NXwY9O75zGuPoImgss2I8XvUH9DmXx6edLcBFNEtOxRxMKHKIlGep6yDHmIcQ1hp+ixr4
ksDrBjFRec1LCYdG4mtbkHzSRNdXRf8H1/LoMss64VKdTVgTO1lCXGnPvjX6LMKCUJmR2mbXgGBs
YDwc/bx+8LS/rc3Dw7WFOu8AJAzsRq7UjbvSAYYM+eamprhH3znm4z0mDatusWqOFDM1jlI9ndsb
mXFfhhVY4enqoyILUWHYk/OKSU3kiRVd0Voq4F1j82U0P15Z3FmXiwJCFsFN+jmfMu/BlENHf57k
Vnib1eXXnVZjg5PzsiLXkf0oc0Rtvthj8XtntgFe9PL7Tbzvn/FkuupOXDRV9D4+j+a82S9l8vMk
6gGdor67X6NRH9VjTTYA4vIT5j2Gd1JeQ1BwzM1SWTLBE6lcHKLumrxTzxGKOXpWYd0pmcT0ivPp
bkZf+PUCnUNrnBPtXk1oCFmwsxLD+ARtRzhCTooHetomaf51nZvK77Gj3PraBnlK7ux5+Y1h5MD6
4c7EtYUjw6jIYjcDZ9k5/Lgg6t70Idfq9XoJy8ihbT5HdlWDI100D8S+TtUdKIyFpkvLHorTBK3y
FqwjB8ETiITjblhbDFxT0oK8kz2OcLsncfeSlqKA1MmzItJl2oTA8gL5HzYvc/JpGi5YyHFTeEMM
4hIXjK5vJKlHpdkKT+ThTtGXoAl2ahUP2jEuKN4ahxZvCa2ddzXna30hufA70MzIASB6HwNDFtg4
EjnxWbvj7QnFNvnQvS6EJ0MCLEFvKlHmJXgMnnsJHmZnCPnIF1j+jMJ8K9x3+9FXaoiRdXsDFXUm
70Vo2YA1PSBkaWJNVFLBnndluEs15S2SM1p+oS0QX4hOotJvVfJEU9LstWYKXv/sPGS/rL2qttIG
mm8mP00WVeA/d7RxyUXf5ejdoyPXqtpKQdBBnE9zBpA2zTn2gImaXA2Je0gPsoYtWv+MRuxPk/E9
WkkRd2onOlrle/mzvGEhkQcIwR/goWFQI2ikL2yHnAOZHH1+z7v0xLkRPEUCPfuMJPB36oXUnWUW
5Uagoqm656DGFHrUJxhwJJmUakKw9PMGmUuiwNvyWsh/PlHXQOUKv9GdX9XDe7htMXaxTn7sDuYd
ePxNUukiibv4tOd1sRS5xP/XqKBbtFIGRKuerVkUDJPEtOllZAa00tkA0TAI5y5yG3WQRonmszXD
u+BhPrVbfCPI6WHKdYoucnHywXejjp9VID1onNB2ZyEyqnIIO8pZovvwtfXPNODwEbWoQQkLTzgX
Bb/wRE8+8hPi050JPJZEP3vkFhU7CRVpw+9ecXSKxPEbwWRsvbTn5yfaYglE+1LW7MO5XuZiN/OH
7t1PGMiOmAvA3VPFpaUA2m9HkDurLhmHPLvYYVBJg8lxOuUv7W1FVsD6m2W9l4wntnAnNJYpOrIw
pjoJKowjJq27hyLgrqCwtYNGwwQtZsuoM+SqiOf5FUDCSgE+ZGRaWUyNiu+7rR7+UBImYiy3MdT1
dNMTFSVGSWbseV1bzrmPx5e6fwWS85989pSHjKXD9f0OZ956+BdMxYxAw88FIvwhdr9oTpa2xeDJ
1/1Rlb/C2n3utOXE7I+eCc23CnwSwjt3SuAzY7LZ6UEaUey/gRjliaYsnjOU7NQFuTYsg+A8a1wM
VwtYHwNUvTYO/fx8Sl0mUtQl/i+pITZSnvRVtNsaHZQHTQK2uxu11ANw7thyC6L9FUXvVAE/Z0ZC
rJ47yRj9rxvs+ii1QcC7jffXc3NXy6aeze2vWYGsihHElPuzINwxxxgKJehDDU5TDT5WrRU4EsI7
ubF9dVf6a0g4K6sUm2htRNQEGhaF0RCEZr+mY+0CKAK3MBUEzd7/2k2E9KLn1YJf5xuRtyMAGJTC
HwIHQDvZPc455+62Ht4Ub6SrZQm1yaC5svU/t7Y7b5QwmP2NI2nyLewUek+tSYsYvO+BKvseIaiM
keWKIgjF7SeF5QJ955oc2d3pS+4k4BLqMnDoXzpPvKF4Ttp6FkycCpjmEJhkuwgAlzksdQPKbgPz
f6SeFdnhFnMkf25sKtSpRbZc8rltajcPtle1ZxQl+gFfZEdX+XvWfF6p+tyzBTvyTdPfn5/vGX4W
4nPcCxJ0Hli+DwzBTGpc8J8rrcobAGMSHFZG6QgXIoangaqKj7ceOfwhlsM0p02k6s9jYTPl50lE
Eu2ol2B3BvSL3dsrPaMJD/MZk3MeCKRG6i6aOW9sm1cEZ1X0vEHKbWDsv7TMt1gmqhmvr1xcGcEJ
IP6KVuZKG2hrsy6ztiehIGJvrsDm1eEFQ2cuh/FKui1g7MB0PTS4J/qUV2oaroaw2h61WfnJa6N0
rC3bodpEosMgOAmSKLqORK1KubgPgjA2EQqKbVsnaX4o8piqEkXa0bQNACHngbky0Iuc8IZF8jyD
4IXN6RrIMFRIuSh3m/0Efxn7UYpTIt8moTCkrUp6Csnv9S4wI3uMUBKo1h2z7O6LgI6hSa6BgNnV
dDEVUUDs4jYw9/Ga/t+UsxVZTT3ngYZ+7SlHGgPRJ3cV3UIKxMYSsetYKkvzhOtiVS9lCwGnuXhv
XnfMGF+fGvDhFkwEhf3VcKe+yCOY14VYk+lZGQMd+v9RTM3s/ptkEowXUd0xSshg1bpIGMjYgOJV
8yhGSZwwJu9oikjCsiGhZnoYFTCoE6n1P5FD2inPDwgdblOLJaHWShgQTOG/ArbAkSFpkcFAI4Gk
FYYk4K8kQyIYCmLjN5SWxAszzBFgF3zyoo3znNXcbTaaGNNi1E1hKqq4aeAhSBgPOZbJVd6dwIj2
c7+LysCP9kk88ogAyGXlaLlNp9SZhvECUaJO04eg71uAy4UMS7eGqnmGZTJ06lPsay0FheRCfdX6
sjLeKlHv8fINaJDEPIW1UQEJjRING0aUK1Em8PIEaKBvqVdDal8gwW2MsqmWTa2l6RMWpI+xKKpV
EP7P73P3rdiw2Bst2uYYL5l4aoTCpsogDqefcuTEe4XW+od701sea0GgQR/yWzADXHp+ReNknMVF
0Zmblfq6phNih5sua5vLwMsqZh0YxneJxf+GZz1/irUSu2+I3HJ061dl4EjCJyjean1ylE3uFyR7
vFiOUC6dX7zVgZzQwgocPoCVWClr7qui+2FxahuTi2X0cSgphPhxokKsqt0+Uae3Q/h47XpwRL03
oBAX1NH7fL+EJ1CIDMeCVVEq5IqVdGh7LiJRaEOeJPrfZbgkCfDKhH/633V/z7Qc7g4dG1/hMUTD
gMbjUVWxcd1pHgEPlLlE7sw6Rlv8/vZ3LfCKefLqTf240U5djGUnhY1/IkruwLIzwxn+vjOVlMOJ
LJDeAbOBTtXoKsKwXP5sbd8SqQwYk4gy6JQFNZfKybqkDW9QWIfA/1N3ZMwlOBzIUnmsvsM/SnTS
oL+SqnPmzUhWV9sEIuRw76xXAVbrt/mFE+p+RSE6m15vhIm85VaIwxqk2SukaznGXsMRU1/Rd5X8
QiD1j3GVmWzOJLdRgWXIuZIIvWp6MQ1Dh5xR2jGg+bX874BpTGgMchOeYh6xk5leWoeVVF4Dvkpm
ued34TZOlpYQBaY1CdI20U4AvrJX3ICWoaDgFHklEkvXwTyTXKhVNmVrQTNo6/A5fTgLCJWt/9nK
iTCFnWJVBtd5hFfjoFyERUcmo/e3RSCIogiowUdFWFrajtrN45rIlfQWS4qiDfnE9LBGHh/e0kp9
5JEon3KRgdVqd1kFtEcwtApJenpV829bmykBstcMElVxB8ebvFtlN5/uPudfCVqN9xLIXanQ/IWq
GoAwHDOFes68DwsWNCR+LVEc6lDfclc3dV6KozDGI9huB/2d7/GGvW8JuN19Ic8UiYrDU9gq4irb
N2MbfgAQeURGdFxLFchCgUaZi8CgXfihPSlFaqg0rWc8TK+LACpnqfKPkLp0WGIr3VamyWuixX5J
1TYVn3m92GHkuE7rJ1dK7WlQHtEKVbDf3zvXPYLPli7pAyC01nKBDU3DFcN2SlMyvoY4+toECuB6
WfKqKJOpqq/cY54Bh3BgBU0hQSxj9c4jDtuqV0r8xS/8/Z1Z0Y3oE5l5JtSRFLDBJLiqeZS8VUHF
f1/2BNNm2af13p2KpteILq4r32bn73CA3N0GSPC1/Jolw2PTGX/alSQbtT9dhxiO9tkdLTvMsQy5
oc9mw2qkGkS4SxM+A05kT//N+IGYhCr3LU72YCKFauZYxThaycf6RzZb73vKVI0eG3akpqq7LMrK
KTIlVa6OU9eTmZWHBRia1utjjXMUmNA7izHzFjPwsVfx1ZqIYug1+Whr2XvMeCRrQ3PqPdQXAru5
zF6DD9bFQwvv3iTM09OtS2nLKa6uvbOly/DKeOxjEwzqg+9JvqiyZE5yCHCyjdWfS9iw4+zk+Ver
3n9lTu/XmFd+kqnzw6d9mVSkOPUzKfdkxUdRErY20omNuH3wF3WzXG+c47g5IIUmwu2yXqoc7CAG
shHzjYUkEFt+qSANla6vyBBpMVW8oRWOHgK/V3C0VoJkJ2+FgWGD31eUQItdamcychpezke3H6Wk
kWSUyroGfLHBXaON54eUzzXe/jGnF3gLUVCDux7/YMLQA92QpoX3xdhsIURwa+KzZZ67Y+dYyf3+
3THHtt99h3db6MTNvemTakSAEqWQ0APx4dSpSh5ReBUVQC3OlXnSTXo9MHg56ezEhsOU66VnRk2Y
wANbocj7BF9pGjE44o5KmrqAW5HGqD3vD6b92YVRfhZAaXIgtId5V77vDM0Q1xKIIDc0E/Th3A8c
zuw2eqT4dn7u2cI6YLOP5D5MC9q9dIJTBbCtE8woL41VLbvZndg0C1vdxoc+T6rSuOHz/q4py7Sr
KVKLMKof1xO4sCiqHYCIHD/xlrY7CNaKQdkt1AlfYM7sLbfxi3zOaGpKStfhyjYHOg/PfeUhoQIZ
iqag+m/+Bsx+EBBdPVpiZTImvBa9Qd9jye/i6zEg6VtkYgLn6mZtBt2JrK0bXVD9LVBNF+5hXtAh
AKqC0VNMtZziB7H/2u/qaOGooW5ykMJW9Qq6EDDO8WoSNCRVCvh+/g1eW/DJ7yOHLWhvCevjsapy
p5ScAyFbFu+xAXcN3rUsuAT8Ap6sNIh5Z4NkTdky+PfUnVPLrMKcANPwchoC+2cxMvrDOh6LJhSg
bOjF9kztJTJdE4hSXGaf+nNr9DzNAuhOkQR4ZGMc7rPhvbwjSrgtN8qGAGeExlAmaTNCTjuYWU7+
I3akXWw7zb83Lg/I96fKCJy7BP/ITMpr2H0hj4/M5ZvHS/4U+DLmjybiDcowEi7korcMiaaZlIif
/wP+RlQ6RswqJC63ggo8F2PGuh0l4TGyxK8IKPgfknDHCSye8SLundRNW2FClFIP1Xnw9ivxOgvx
ic/YT/PtafXv89y2oNturFwj3m4lneNxcQKfmMLYkWSMzppCkBS0olcntljiDV0eGzIBuMC/zGpR
TmHZXBPZIixX7q7hx/qby4+GoI0O0JBkJIPYbuYiCKB/E21COqgJNUCQvFGJVRgRoWxqzhiBF72i
fDbaTl/Rs7S29C4w1S8Bo1kgj4PUJkkHcU6v7IoKxvUyQVI/Z/51H8YYxYNBeDQ6MYxPS+2v15pi
urwtzclgOSMosNI3Mm2aO9cvRS7fvYf2GIXC+g42v5upkHZnW9OBRr3RZNCRkmsK0wqZ5c2J+DHI
HcLWL6N2GNjcCF0vQuW78QUTd4BS6fPTSjROT0wwQ9guZBUXh/BR2z3V2g1EqEW+pu/PLa+s6cbP
oF+ejps6Q8LUhj3NQuslM/78RaMl/u+1Zhr2NQrb5D7qMYCFTPpHKp1ps3UqjZEfESnijffsqcbb
AC5k5xot7G7h1gfmIPGtjs1zrPOlJPmC/5YH/T6gITlGGW6E93WWhkRq6T4jmt52rcFrXi6ScFI1
XYPoos2wqeoURr2PCY9jxcj2Vtb4oDYxCyq1ErvubiC3whva44R0lG8BQ9lv6CTX5UHo6ghJUsej
X8wZYpNSYvFXL3Bs7Xmcyf5BxhdTCnYtflYa1Z+oVW+/BA77w9kHKUmIxV7ULKO7Q+umQlcesYMe
09IMkAwGZ7INAPhdkrkBzLeltZ6wWkRYJFt5L95eEhseNmJFSnvscaoULUFL8W/uaLSF0i/H/gfq
uyphaLMDKlcmse0hxy+rw4QfbRlH95XJebVUvg26C6W98lfrbUuoYxGAbTpKVk0vKDiHu55SeC84
sPfFLd7+aRlOCqxDAjd2A38wEEtSDFi5b34RiAwFO7UXvuQ28pnQ8V2VEwlmTBFtBcQAM6JZ8RT+
jbaklhrN9Aji/yeAl48og8knLEvdIWHt3M6WOxFCcv3D/jcyKpLzcAPAl8LmffqJga7cmDoacZNm
EA8fsoK0ybBLQwvoUV0czx3BoegvAq7b/uvzjf+0agv/cLvvIzniQROLgX1xbuf4yl3UwtJe7ziY
1U5aBW3lMqZArxYxrtYaVl9jUiM9ZJqIes6y85YcRE5qHjc54li287HviVGmtG7rRyk+7jJpDZbE
Ylxe+pmNasDCVrIGGCc8XwyJFoCUraoYcPM21NyNkYgUX+BfpBiokT41dx+zgrybf8PgnD65Y172
4/KiLiGI4dWpMJ62cxhyqULcijOGsGpEyDfuduAj4EBJQTQ7uWmFn0zaFrlg4Qp3Vl9E2Cz50msU
KcAKIH4T3NkRJQXA05nelcV9CTI5v30oYIEMQOFMwt2vr5qELr4VPEmB3fzAob+IRubHFFnVYesf
2QwaaYR2zBAn0q1d8c/FYNzbfz+WqSwsT71c/zI83wn/UnXVm1aXWfZBVUKuHDGsX6EmziHrfzvL
tUnHQ+8njkBzB57DvPtDT72tvswWGhd1g9MxRTIDdJwS/UsLAGVY976dkhGUClPhCj6VlAL/3JBf
bJB9NsXZVINF1td0FIXbCqlUae/COSPoF0sxQtuzl6aWac1/WniVSBulZ8RMcz4gFiFlPA223tqs
MeOSBYpIe00/U8BvoJD8MuJgzg6FHNt2kl3/8tdVl/I0l2DlQUR8uIi4nMihqDiuCkdzaXCzOs+2
yjwaGSSAsaLnmHAlLdno/ELW+aOOVYmR/wDq9d3F1f8G2wSFpYQkFiYNqjOvsJeFpDHrfJqst+YU
+ED+OYRwcuMAgxfL/6kxIus+H1h8UGI1QbYyc45MDuGV0KajvmbS7LJ5EUkM2peIezqwYRhGn9pg
QIK2KKJEEGcBuUNHAUn3Id9+ilO9zF36mNESkIpcoRJYd7KaAY0KVDDkLr6j9BHaQWUHQOMPhTnO
c8zKINCgM5/bM6ySYyqTxDIbeHDxi2jAsGU1X6EmWigPyO085Kcd2LA1ESsyHdWj7EHkjmIVMrLK
yNZr9t9NhpP8dUtkfjqj4mPG1uyEN0m2plG9zStlbZgvtzFVvi/Po5wRY3h3+7hujYDtJHbqeC7/
XWc9qoYIK0vrolaOPJjTVJ8/lXYn0TsYPAlzDhEKGwqAIAGY6z8rIQCTfl7yabyl8W/CXO6QEC4o
pY3PkZdsEPZdJvy7PLq9z97mFH+YrLFiCnb2mReR6ouPb9Ppr/S3sq4oieTpjyNmAzBBIONdEX/l
+eY4UD78zY0tgLJsnYaB6K3ErZPVU8sV5s53kXBdpF8QZw1vvutunWV6GvPahPvnwD5BZDoeosqL
clQXztyX8BP9nLZ9m3Mq4hhIC1o6C3PJzuGVAXQJ8VgbEU0v3Vxlaiwt+2E5kogIVPxc8BVpl4b0
H+KEabjo/svNv+wZCZDpOFUjyBXhGJ5nVHg1cnBuX2MVSdNI3C6cN0AWCzf3Y+Mjp3WDtsfhkON5
k+EmaR4kES2geWSrEOQQU8rfPucu4gESPB+QcChVuh0gescoz4B+sd7EBUO/4eIDhMENbZ0y/7Zm
1ILYLjJZLgtcjCfcLbyQX4q0rfbLnOPHnDuovSis5qzuSNi9wNDKHkq0MGsOahiMvKd2qsd0cKYR
Lt9UrGCsTBYXpyA+BCEVepbHOQqcrnq46pmndh52RzP/Vv9R/iBjivsaUHiKjHq8C8NQWcRyyEFU
E+EyPN9+IYbxa4EOtxu3USI842sfkyUb+W76dnbHwSCFBmlY1TZIQlf2UISoPrbpb1QceFK4UXTr
zwsKHr92L0ouHKlhaWq6t//UJ4TvSTzxQb2emOt+Ymfwjbg/rQf2CTFn+szodFwdz6hfxsxaSiOV
NIu9fHux6ZrdG6qwliGStzbrvtJH8dr4kRTU5Nu4oSeKyqrzq6uCzL3LQEkv0sBLf31e9AxzTj+8
jKrsCWHJY7sAo1Gd/5IOKySCAviSXC4uL/U8AGILqgeppAw8EFAOyzfrW5KgTYaaKYkOekC6eBxO
pWUJxbRlldUCEkht7Zv46b46r6IdvnTm3dr/FuCwqZg8NVbAxqTPVSGehFzpoMVxbUCKSTF6HudI
CBhd6HR/mhV0xLhrPP1S0AgUhvjzOGSfezozw9kjsCwYhK8AD8OXuD3R8hqAUDV3/0YSWsvJMa+8
Jw+w3la3YiyYohLpUXKt/ZUbQWCJtG0HgRZgJGWsyZi/fryg/PW8AaLWx3D1OtARwvAiGDIVrtEe
bJR99JDmPibFxLjzDrps2IWJxJk58UJWtLkr0MPDo+E/I9tz3CGIkNHnF3xxfMZ466579UnCWAXy
/7tJXaozlzV/PUPqy+tVGg6kWq1hjUyH1uRm2cLF2mwLCKfg7SBLTQk6FAlJPqwzgeMRMUZtJi8b
tGrfAQjR7lJC0HebN+ANXN7T7+8Q5+/giRk8Zw3umdU4NFnA6772u+vE7iOSDFFVUeuRZrCsQgfx
jMprmXYWA6KZSsQ3iCWgWH/uQrmxiXGj7LBJW+9dryG3WLOp1a54IIhs+wtj+OIwW1BigZHixitl
/cUDRxsf8+3AYgpJsTOVk7sSF1FuhL2279SU49BGUB3xfVzjv2TQICWe6DxxVdU+efQuyt+x7QEo
EqjiXmxcPXsgOVy2XhbKVOEdNHMJzpBdlvoMhM27a4txV42ZTOxdzy4Neq6NPpwzvaPH6ogv316A
EnyI9DEXcoDIY1QzEH4w7pk3pOZXaCa48WgtPKivhF2l0hX4byXt6v+ETpFgzkpRH5t24TR5Src/
29/4jAuO8LrtlRSVpgvmBSfY+wJpo8CK7P/eTEH2rWchsfNCRgFvWkKBleSuSk8l6H9fBzfo/jtT
JbCa0hDj1JtYvb1jxgduN2mBR26MNFpFlpAOWVLXJytFCO2DGqwWBQCPAm1SZbChGLcOuR6uJzhQ
U88ueFlA5Lwwukxah8CV3jOcKJ7+HEpFCzS3Lj+5vu1E/7JoNZOkgMdY6W8JSO730CBBjGUnVUBD
ATqzGQAxWVczx5YOOBoY4WQWtqj4V2p+hbimml33Zz0jDy40Idbe+6v3Ue2jgnXEscbvwN+opfiM
xyRfkhQRghoHWk6/acQDmCT/pWE0GEo7DjodMKhscrI5hyZg1fc49TjZ1s0i4EuIlWGZJ7QgXoxr
nbhbSnyecTd8c3HxzefN28ulazWbQvVgqH+e2YcULkLLSjo9bymJLAFzq+JqYQ+PJrkwJhEg1gp+
1tD7FZKFyrpHsmGHLBjPjeEmFZQ7zCZ0V3FiJZC8wqeGZkP8apiJp3/N6V78KGjgibOrX5Zb7GcE
eE/hecVWdruEr26i5GvRvxHCy+trzZum9HoNZFZZMIhN/+DoB9lRJP7tgBahmYk1nJPEWU+sNQNh
rE+I6GxIbTaDMsAkOm9xqCeX5dh/YzIhOdgft+JsweLmonGT2U0Hy2hxjbMpPh4AvEOUYmMovif8
eSZRxe7P38ekOn70AU6R7tvKvybOxQenOpJkx07vFVBcBEtbTuTxz6iGnFG6nWaNpQwZBRNorzI2
DZ4M0NWnwIcsH/xsLo85QxX+oW+4SxaTsxn5pOjCQQLl0qcBE/KsunaX7nMcSUMrZCRG2EwI4GOa
Dk35ck7MIt0ZXikKAe3bacf7MV1lsof83OieVA1QwZ0iHn8di3LIgllVfPymwfU4H1ffS3/ISqf3
Cou24Wie1QrKwSiSY+KgmjNPBB4E4QwMtX4OGTapn8coksYDpiYbzur/GE9L6Q3H4DZ8gY0K+ne7
pINka1XGNueSAtV1/dCUEXrySmdQmbfckIWYrv3VAEFOgbwklivyqBiQ/Fz75f472vlW8RoNpOh5
YTU5xGnwDrXUA9ecf1uSo77Dguj0wxv5InOxjJfzqOACyUW7IYjfR+UARsTv171b5xaiGJ6EF9Pe
UWPT1BRP3QAXxqNm1XRC4TUOls8uoaGmf6/rB2wHfXmJSjFVA35h4+3b+JyoHKZ9b2rsohCZPIXo
P6XIPJuDPQAfPSpsAwSFL/A3NzASE/K7V4EJPG3UWV6rRaTg7kDHzqbInXniRsQBFWsfa+J1QR8o
pjoFdbLPHxx0bJxFcvLti1wtyq332MGgeLAwfs4pVjeGf7ol707+0fMwsN76lUaj0oOH4j92noLR
7Ftiau1a8Ux5zluQtvzkgVi2FoMZ0BWrwfX0FixmnlM/QZsfV83dODWtsK6gW+3OVEa6gK/+vzPj
cVFOvFh4CyN3tFCZnmNcRJexpWEyB7kXLBJdRBtdQoCf7Vf9iMNFKP0RQBag7fMBabZoxbFPZNO5
PgvHDa2KHB+b6kbEsubLBk+rC234R9JdvjF2gAQCzyjyP2nubKVAhlggDr/7JrGfrWVZN+yDqTur
URa2Myp76BCnpUszVx3sO0GyzjnmYaL1GzIOOl+PR+4GdXRNA/c3AcKkFQwD1bQxA83XaCrSNOTu
wWuHEQwDjPs+7JRQW6sp6r8OzqyjTvVjH7Exsk8JaMYR27rAR7pmPn6zCYq1zyibZI6nQAN6gq9M
iVimIJLwJKERkVGFyEbRIQz+MB5QYnmCm1bOzYsaKaK9nk5BzIDAsltpRHJj9LnZ9f6aUh69b6z9
zC26z3Oc7eq6NgSZirDwixbOfJLJVUI6qH2A6olol6kDo+DV5mJav65v0thcNLlkhyZZp2IqAPLl
w94+o/wEnVJW7Yt9s0qc9M3I59QnuwD5Id9ousbcEkRZ5GE9X8Puaxq0RK9vq/4m3IyE4j/JNoz3
fpkkoPCEv000wAAwkLZSGcGBIKUmGSW6/JQTCLXGPKkvmhtDWt7PCZQCA1zsJa1WTUwBJQgQMjZm
dookxlo3O6y9ObE2HCj7fE+f8jmfbYLTN0UJDLtVHpHxpsezKY/QTJkTfqbrV89SQ0W1sYzK6AO7
vJhiJPlIlFw6EoUmGSSl8zzolqKcGeVksi1J9sxS5hwNaRhYIO4K8fEZyU0Vfak6FkQF/JcK4gMI
D0i4UN6llfpv6iFulPH0zeVbEhtJPKaBdFpCv8tl7citFv4rl4VnsW1zuA+l9nEw/1eid88GxWoE
c0Q/I2CMMyGeQ+0G+p89wN0O+QYfTO7U2HoXt6C3BTLZxyv4cUTtJPUGu5rZkj/f0+UWim0rlhDQ
DzDYW8PR51C3L9PT3LqSZupoL6ZMeW+tZsmAfaaa6+xOg6x733bj4yZs4/1URNmHlmYZWJ3T2N/n
Fwx+ZtKikI5V+6a1KwV5AwBAe5MNuZWkeMoN8jAGkRtTFiJ0uzI0BZhIg4UxK5YSXGt3N3opYLFw
DM/GebDbGR3jtrO9Uk9OkOERc+9ypB/XBlGECIE/tAIIm4Y37/WRxTB3EyCmnMdgcrKhqapPUJ7z
3FDH+H+Hm5vAWElkTFCWNpALpNOATToGv8E9zIw8ntZIJz62KMh6yVVB27OY79Fvwg0JdVvH5Dz6
W/DEu3VVFPw1XGmMEp5dneT4HSMgxZkkTg5M4UqMAShsPNhEL0r2fNcdm9eHqF2OUZ8ol1rbVmw0
vSNZOcEwHhHdefP2wZWFmyBLKZ9M5PM7Yu8kr/RrQvVVsJ2CE4VdWD+EUDi4e9kJnW0fru0FzRYy
luBp3q1G+Q05dgrYGMBfpxqmR9oboM/szCrsDPDx9+kyUL/3krvQ4iaEl04KvKzIqoEas4cpV4rP
Bdtw2JNeJK6za4qsnjNd1e/F6mF52MpRMjPA8ULxeh+xb3nbklvc4Lp6Xp7dOdGaIT4chRu1SJkt
+7/Cpx5cJTjXZ1nzMU8tJVcWzAmdvcv04UxiXaqZFx1wQKHwK+L2AOVtTglvaVI3dkM3StSvPHRz
CaNMKxm2v+dhW7/oSiqaCobL3/zGYE7BheP4MnDJdgKoJDndYfWL+G9lv3vxB4Q5AltT7rEvryi5
kZICwnukX1XsvkBP8ls7lCTvxQPx0Z6eYhm4wdD+ClDV7xpOSHtTe0XYRbJ0kOvTCkRENCEAAfTH
zDLL+lnis5y7Ez0cWEyTU/I17X2E3R4HcPBT6hiCVUCtZgQC/ECzpFqasPShW87d+tFFxrmzEMBC
AKcz3ZfvqA79CWgThXzkOjVFTZCdzdiOg5OcCsfZLWuYQKGHpD/94ZSPPWidrF1CFdJJiSao0lty
mnHn0rUjjHoNCwiaXqBufqsBAzZ/YyAQGOpqbaUBWkYQL6/G706F12iV4K9d3gtKkUswGvjLnOH4
5eVABXlM2Ho5R1a2mYKtdJ5FT5R3L8nKbrSV9gS5QJD6nQVGW4nJMj4J9KYiaQyrUjZ355w0lCLg
lnUzCCd3gB4nwb5Fpq1R/8pXiampRoBItUJxfrxWfl9BZGE0Dou1pOeEYePAoxJGE1OQbF01H0iJ
7qcVUL8a3sGsm6R7hR4ijjy3zIDbaihqjjQujFYIlnpRk6ErCrZWUc7lYS41YrtePDGd4SmfuiIi
Zuy4i+jqiZGZeu8IpTRkUTVXP8pzLqizruysTTZGQuvdFevTH4+TUQNBsjbYjTnkS2u+rJUglIpw
Fxa9oby1xApHYDPRLsqXVPiFB3FUI2dx314so/zAKx9k5TjUT5Mm9EAosKXHXBXZpjFdChA24Ab+
54AFPRzcDCoK2Ok6skCckIly0B/vvOrE1jKAotXOvhqNalx+/uSZfBpXNBo9fGl3uS7cQLDiBtbw
e7qRT+0up1BhWnuswiXC0IT0rKQbWh7Klg7EJVaroBVqTfBaNA/wkVYAv5OW5JjaiDlcWXri6pTi
qXnH5hU7azuSB/Ml0XqtMDahopowbhDu7QeKFqYA3iZO992p0+7Se6KjFMjM9dPxSZZZh4tBuPnH
C9Mv9d87sNHRvZqJDGSmlVefuoqPqu3QOA58Bbi+gmq5Egm8NVus+qfKai2Fx3qiB2wpB6hWvvGj
VbHopFGszP/lzQsIfCcuPTVyhnBHl2wraxIGPpn5hwrBNTQLu6jFo5DyjyFQqc0HT1CTwMk6+pqz
NznRVLiZScPF+9a4BpDzgOiUNdNYqkcO3kps7ajQnFMJPsLxbVTJxCuR+oxUR5TcHSC1uf92T9Hr
zo0aGtz6UCELT99fZM9BkAeuEEV8vgNSBMUlFWZXrm0lCzzD04baYyVJ2JVaimcNGfSVg2G3JtSv
qhp7hWWfLf0GO4iTY+KglWkwJ+hC+9AupOTegundN9CEfT/ZfS1/5LjVq8AIZWGPnopEVQJ8scio
y04bqSY1ZsvXRu7s773lri8PCPg+CamhLeoUQf0Dbf4lGQMQvHBn4ktMPBqm7CBlYdpNsSIkY8RX
kVvo8TItHJ3XFrFYPePNih+SqfwkL99YajKed3AIadhju0UZKwRWs738nfK2GLdypWIh/0I92rjr
BVfdkLVoRy+Etpu96xmSMNBWPuNIKBILmWDDN8meUtpmlNgKJPz9geFStNpUY0G8GXsh6xsMc7Xv
HZ6FQenUYIdDEOoeaStEKBieQWPzhtwobGaPpeRs3Wfgcq48PEDBiROyuLubn0x6xAdeLcaGq5/+
Ia76BsSdOPGrG9J0N/xv7U++ih/6zM84TgNtKmWTcK8RUSmi3O35d5kV/9av5ovFmqx/ON+1Icpg
549jPUEDSMvYd+Bxm9qv52ojL3U+deIvTpWRle57d1MpDzEJ8Ti58DLDRHxNB9SWzHl7UeQxan6Y
bB8hZYOn9ygf6b7L1YYKw1xR29VpstQKuLLa9XXmpLrFrN+gqlZM9rx9tGhWr5NoN8z6Uopdjr1D
ErdQly2f2+KpiyNc8eAPOW3K/jUOPdGQwm971XPbIfRoKaaw+96GAM0jnTjU4LXNRAD2yGE0+MvK
A8gYZvZHVDurlJ1ypOX18WgX6dYj1mrt6/l+XXD5+L+1244+KUvjI/p8hqyGYx8V0CYBDk49w/NG
gfdGAhTHQtQMCOl/jZM+rpl9mgVRgqa0HFVtWd8nBHI7COS0Trc2rvcRIGIsjJ3T2wbeKzVWXnsH
5DPM6xMAj1iiewzMZmDfTdx3ktt0wmU+L+a6dMjkbFGFmYXdXufKmvFBAX1/viTrSb3mvPOPP8Ho
gCcpb+CWJo2jka7ITRLJmDeE6vP8e2gGRwL+R8+KtIbDUeZEfgA8N0tUmgNF6DHHG5UURl24YP80
YiOsDOzBMDIFpayK9HETCJe+YBLqdtJEYN8wBE8IDbt/zEEvjpwzsQJ/kd2hwiubKlKoFWEXdm8+
TZPLSYNBCVfdDr5LjonT9zk3aD/pvx/ARyTs5fpiYJTE2O9FSb3vPodyYNQcrJdDAyq0673h+wsH
U/jaFW3V2EIAGPJyortS0NGyjA1wNeOoovn1aD8oJRHHX9YE7u8WLEQeok/y3iPA8PRrlPVkSUgt
fdQ55N32FT4I9o/bWNeFiTKuXQMypWczauMly8pnmN8dIdXttL+lvPQi3IREJudBNv4CCARMf9Fr
OwKFPENYWiKiTVnTDwcUgqV35fQ1vYe7RDiRr8EAe7AEQoRkW7Ci+A9q/tKJnIZYDZaoN9DiLdTY
tWh6RCnIFjxEb+wx3cqUarxh5T+fPqBHd4ANxJXp622DQn+BiGPfJLu8OgigdAEEI1dB5F89qkoj
OsMd9R1VszeOqAGvftDle/cFLnKZk4sMBD3l1GQ37jhl7Bor3V6YwNDmPQJECY6Q53CoVs4oHlpR
qcH/flzC5cowGLwkFTGUhVocR4mFAWrgVREAIPlAccl8Z9mTrspmEq/++qOSWD4r8CzAMIWm4MJ8
Do0Ki/NwNqXcobUDZBDbj/W3d0J+sTAE7346GBlKAo6CucZCt151r/OggT9tmDaEjUdjunJRipeu
FamW2cHsq+XBut5vYtPic4xsSBfxmW6cwNHPjEEcCNHBIsph7bQzCwov82zl6wqBnb/0uvlyXJLy
0CEzgyuJoifruwEn71B/bGIeo/3Tk6lEypN6VVTwEeSKSM8UPp4GH2mlZX9fWWmTWHRbuw/3PHD8
z9/lmOWl/2jgYliw7winCHvu6ZBCkUsmUwsJ1N8cWe3XG4V3IFEUPEvqJ/S45ScuKDL2NBebX107
68+feNwEjsKYpiv9sRkTBftnlTrmeiok6vTdYVng57b+8TSrXFteoJ/eitTu5tw+5J91fnWiRB3R
eI94ASkcqkNwCIApuB7120WDERBvuWr36tFSwmZgMuQ+VUBAFOBqp8xNwRofU/oqR7a667AgmmUA
toLG4F6r55B8COIbbmlKsn4H3WQKYxeJzJnTtt2Y9XyCm5wUotNhz0QAdOtqoLrqmx4i4n4QB5tY
T8YcTfGJhfWgKpWRGgCRlpa6RgNdxsHZSwNXyAUisCfLJCkaOF73eB0tXs29VzoEsSaPJ4lrokcm
XuSv9E5vz6UInu8p3772juLlEh6aOUla/odlpdR51zUfCtRouFog/Is/5q8kHo+0Bk6p2JCIbqIJ
ZH2Zg03b5h99oEfGpFddEqAWhDUVvE8jEJY8myTiqNH5FqvATX2xzTe8qydB/O05AxHOI8Oh5Go6
4dPAlc3N1CzwC7AyPiPccDrOAzQdKkzyOLOXevR+80c40FyMGRg5QkHT4hOF+/fjknH4Q6sr9y2f
VoMxMjBCI7Wx4WGeOkDSk+65ENi917WUw1RzLjuBEXnA16ea4AJi36IlylttNRecmVopYzp2kF/F
lworkOR0xtpeSpdP0BDQC7OyQsRDbWhLPrKaov1rv+nNySoGx34t6OnwHTnwrTTGafo1v4FQrp5D
1hEAl9ps5WaTIF/3fkFuE5LwOlZYG19thVpIWfhf6Vd3iKVHSpTn5nRZlxdOLSENcH20T+zrw9vh
8fnJnAYGopeVQ4+sIzcNFJ6BtqqgZpZ5Au1YK1D4DQbqi1y0vuBbB+AF8QhfzBHScdgTwpsL2xvg
nawazt+/nMrevIztvyPnSFscT8k3tjOUTqaA+koqlqLdJx4H6SPayABCSmeU3mJxpRj1p2U6w8Rz
jKBueOfC/6MnxL+h+tIdRsJyp0myxwNL+I4etDDs+hrAQlJ2nQW27Ckt3lMCsLuKnixFsfMjsO7I
2y+wOk5pvGtoHsITe15pUDCZWigIlX0Gd0WrnDq/gStEwiAhCoeuxlQFnpYbW3tFnbR75cuJHQXr
PSXGCfGD9rVof2KZfsKn98XLIQ8AdsTcLG1mVcX3FSuk0ncCNMxBJ4J6jtNw76ccwcBQkfvHpHIO
gJbSwAdiZkILMP9aTDFBHN0Ylb2bY7U0DpNmFdpEgpOxuGcJO2huunrQfpu4SlmHjr2m5sUomFN/
peFy23aQ7JtxfF4VsVnt5JQBBCrdRGNOnUZrVeTh9CYapC55HRwYnT6XxNai/j7i/2pPo7sI3Jn7
UpGhdgqn5nkgHif0V+fCcpINKlKVl4vjghH4JdhDrpqWJWHO/RZyI4WwLOMfHEaMXpnVIoZ3o+G/
A44HERK/jHZPb7l5LjYtykb362l8VRi18nTjkxyGDXR8/19fo2/xpfY7G6Qam3RxqYEIq4SvD3yR
C5wWmtIUcRVOb6t15OKVPDrdTkoR7QDxQRRBv19y56Fai0BTVH6BoMKVXi8MAjU5VE0c/S+/8AJH
FoJYuM1wb4dCjsIT68s95G7Kv/OkPwDJ/+BDXZLUBTDQ6mGVzV05+MFLhVFJvRsPl93aYtpMvBvZ
NetBeFISWOWwrDTgKp/O8o0Bhzk8SmS/BwxL+V2UgV+z8lwdwYNWkmHEsphxhhQL06IXJcC8MfJV
MaMPcjCvYGfKnKFIUgZVjnkr5tzAaRTMBmLusKa28E71/BUIN7/5Z6SvM3vS98UC1v9jqq4bV1pw
8CwGsgH6e+vMlT8qldhz5p3/zeJQBbJlhyESXLMQ3oI2XViypCHarEOEv3pyra84oomMnAcI044P
uo1WW91YVEknxdL2vIfFCxCGnaLFNsZBj4XMdPJ09EHNEvelyRsQrWHqa4othYFrwMx+gsNAg6gq
X8yS7LEZpkxRPx/owX+OuNUUvkvQk/Ex9XIYUHkTptXprRTh69zE5ESMKl2JBwr84tRUId0PC6ke
Jg97CWZd6PAXJGqJ5D06kglJGHi7zkBpGN+in6gnQnTOc/VEdJNkzuqYRVbCy2iEt+Nhu9P+EgUr
lajQcRShM4gzZpITT+GIqok7cq8Oh4YjNFME9ZXyQ+dwlYbX8TLDLfEy/fRbZEFLDdKKhIq5EHQv
U8VbFTLt3PfxCtgcCBlVC7rqcxc5xzOP+Al0nS1c+49AaqQ3K4JSxi3hwLB2/MX7OumX7GNMyCqP
piEncU53d5qPS/+ufwj6BvItZgkO/Z98MiOc937FuivK4xV7I6TZkjwr+qt39mKUl3v915+Yd4Jo
NL0uRaj4myLb3n97EjyuKSZX2AzJ1Tp8DtmIwtc0yUYMyBPyVy1NFwZUdefx70DU4fw+LScOAPzN
G7ER8OR3hj4rThSFApY3UGtgXOHVesB4nBHKoFiyRv/HxbeFwVLHuf2KKIwUfV80PrRQ9tXzMBfm
yh2jv/RTI4vJ7KkDZr3DuuTqtiyrqL8xhDvcusjR6q5CEo6b89M6jbcpIzfw+jMjRj28GfmoY7iW
A1NwurBR4boswiQCDe9UpSQbpq+0CWSL/ygSSoLA6jlE0VPDMv7DDdVF9nBh/hT42Yqy4DMtR9dg
czK/YRXTecmp6i5ObLfM6dW3p2n8Jn7W7oQN5S8azDYtZFhi0OGPxAAOq7Mm6/tSbw0LxQXCxvUj
mBOFp+vFGLl+5D39KzKNjRVawuM6/+IHzpGokt9140Bs9MmFIRtrRlz18Z9tbzBR+vzUO8jInYZ6
RL6XC6kru+WgnyfzhloyZF5oE2anHeZOPeJjeGrTPA5Df5aVNm6uGfQk0a9E3MWoJRUGEg/tS/eV
MZB2TS1bilpJp32sBW5jiNnGORnzzDOZfrdgouzeceTKsji2MkI6W+PTDMhrt6m1A6+CsNW24pge
1QM0f/RArxmRL7T3wywNFvNlWuWeV3GOTG8ci+WClRElykooO520P5jXSn4MfGoOr4mzU1kOk2Dw
fp+ZKR6089IPiwlsjKz1LBNo8D6jz1EHrsj6efSbaTO0UXqdJjOUgD85JFQqDYYC6M0a74KZ4mXX
k9ivvCIasHb+7WhP5bAPxOgGAVuecqCKPfeuoi4kDqv4OPACTCLIqXx2mtJn1XzFxcXTN9L3MeCX
FiduxZB1kRHI4ex0G5/SEIRw98rcvb3uPlHh/vIgosnNWH87fD8u6/LPFkoNNAZnom96fYBpMXyS
jZDOgXun6tCzM6e6vb0e3Y9nRmNFGJHDtleSjqPqtgyMvrZpqG9uoKMEF9hSEhIRjnyalsgcTtwh
ifWPMeKLTPlSkT06FKkQTxjT9KBmn2yIVbrFiN3UjYYyyLjfVKuhWGtjl8esoT0nP8Ug6cvi2pHR
XWEZrE/VfxCGACGnPldSD5SWfoyuxyTEt5EFPYReZQTnHrB24VZ86I9rKGPmKqAWw0No8XMBGLd9
dQJQhdmOC4Qj8uwD2Jh3ag1aKTr0ick3z2BgC13ZaXpVMxkZBtaCBG+8iF5C8xAtNzOZbklSOH8c
vIBn4ZB3J8xQAg3Gv6QRFAxlnVsDSfVL5rfbXMgQYcoC8aqTEw+lYsg0fJAFA752aQUoUU+AefSZ
+QdH7Drms0zIevbxTTzoEV+ybDuYyf58Is1Dq3gJIT1bgr+BxNbMzPglgq9/XwTw3fXzaWDkyM64
j43g/BUeOquWOJ+c+v63HEPn1AzukNGO2OzOXKC3Yj94pYqAaVB9fW4FgXzV1qY4jhLB8jcKRI2h
0hl4+pg6AIb9laj6D1JgFKmITuDV4+dOYBu5sXQ7hHNz0m4++OgruW/Lh8REcvYvt+nJL4l38cLm
SKWZeYtDDgbx69xVW3mLuKWaxf+mFuGQ5ON5PcofRPCAPdoRe+J/Uc+DVONcgKFU4oxV1jqHK4qT
WNuhU0LhU+iFiNzWZKk5vB/OFygUTKXrKs3j3ypKYhCAorxL69HlTnu3OcHugPNZlQcxKJOb5pXJ
oEvC8UeuOvfQGvyx0OvkAVI4A/QtKncCnjtlV/gsDvLVShca+3LvbdxXomIodNTOHWfb4ThLJy8B
5iVr9mUhyxMSuHU3Tc+qO3VYrFOmWpsI6aWS/NrVy0gD/8A56dUcd/D39P63rOezoScI+gXLRAxD
osTfjyyqqtCCjVMKHmjv+sCm4Jgcv6jnxmIIjvBa1MRjg95KPPWzuMpiSv4+Az9JJKxl2KkPFBiQ
jGg9UaFGCQXNYhSDaacH8yttux2WELsGKbQDVjYF0Nj53prrTSGNjNyC3gO3+Usqe58XsDR5Mpp3
Nl66EkhuiCWgak36o3iXovyeUltmixn5v70EupYB05ud6zqnsWUWFyT15YWP7PDB/OLIu5bmzhCQ
KjTZtOrR9KyAiiyypb1N4LoxooRy08x4d65b48V6e24iMbwYN7v46rQ9INpH6f/k0oMH+un0YBEE
rmCsNgQauOmZqYxRJKa6Zk9n0SWym7Gt14r7fGCJ/DRG6Lh9AnMxYq5UoiFnEH60cKMYhpYm2TY2
ShzHDxxq0ExUwlPH6LovJVduP/POx2ykehka85/Uw6NGWzbJjibKN13jCKSVUQO+M4UT9Phfagtt
0gxgXMjIGFk2C3l/+TZ5zU+wwZ9OuYyrsTOdp+/R7D6sp6xursf8Xpx+DJqsDR5gKY1qchSOTueO
t2dDq9YNVZjaxQRVUgqM/EYUA7pQrRVjqMAl/YNJoFryQlYRLQoPZ64p1eYHbBcVJW246etjAEF3
u1yW2NlNmNp1dfuD3bVl52OJtMCSM1lBqzALpBpI736bNXq1Vz6mgN8OjrZXSTwnJdM94URaQr+U
ky4uHXyXyc4ikmn+Iki3Kt62/pOqPzjCvfKIJUsowhIod2RpttxJpQ7/fwcJGP16axo/nhswbQw/
z4QC5GJF1JPThfRhXME1gVqORmLQuRknRqL+DVpVojT2LXMd+Fa0WJPGodZffRbAO+Yx49LoPm17
awESEwelJrF4erbaa7pRc5eF+4Ns+esxfmaIEXxd6Zhemjzeswv4sPUUzOdD406DTMeGEbSzBn4C
raEe0nc3gRFFddD0kkIIj3GrvKzjbAyT1G9pT04X0bv0Dd0Si9gEMDSS5ssjmLw2fvVuOcBnDxar
DTvnCAHCb2a5wu/VlKMNVJRZwYJsYt3fQcIsuAzHy3iF3WiFeHVRY5hp6sbc/ijSVGmxx5WWi9NT
w1ewo1aZ5LHzQTBB0WweEhFZjvtTeBdHImtbYo5j5X93Uc4hY4kjnK2E3gcYyd4xPrTDYwCsz/7a
vCDF3ErQHgJRPhGs2WwkJMJuXPdiLiDEmQGNjmRxcY5UrjpC6+ALDpw6QXAYLlK6ymAOl69TaQ8I
uAammrad3sQaizYm0tn3Yq1eMiqmqY2ZU7NV3MVQFfDMNDPPM9rkH5GBIW7h1jXzdtRM7wMVwECv
X0UmVv8YcOvjfE/ayQw0Fcuo6vga1ikPRqFZWC1sei3kT2z0yixhYvNuBK9OZt9yK80TFC9PRJSW
pYcwA0dTEB3O9XDVBHMo+yUtx/ow5PKIQmYj5mUg4UvzY0+y03twg61buoc0MeX+xHDZSuHefdyT
dmvLF4iPy4thvNOhnnoLFkKhBo9O0p17/N3tZoQ946krTGKwmS4dEbtZ0DpJ/t+nuwm53+X7QhkF
mPGMR9Doupr75dD9lH7orK60x/2JRgKaTx07v9IyeCszeM0vFH6vHp3GmwV1+zyYfQKMmvy04+o+
va0rXQvsLGemrZKw98jkrU+q9kEqenlwMc6xLU2ZZGEo4nBoDuofW33Y88OGul3Inehq5l9Mpcww
TncujNYgH7du8DhdNkF1FrIDKiBh1dxTt4rahjkkyrAVnbgDUWTTn2wD3F5svFlfkaJkq4JhF95Z
FvBzoshdHaQYrhykeY+R1rPm60lSlIfharl4qav65Y6euB6P3fUbRG7EU5aqleixlbvCcmwxsXB5
o1BJcoSqx/t6VYvH8R2HVYRSGvJDI+aLz9ZNkLUpAW3YlBr4J2x7vD0azDTjz+ierylWADibTkqb
l9UTwfvfBgecuYubRmrm4qZJTzY34kyk5w0SGJFeJMAS4+ZIkV6FwRXeH6jtS+XUYZgNBIOWnTTr
700PKnCZi3xK+QDudsSydrXNdHO/atMoNT3mi6xctIV3ux93APIVEgHXxAhA+VpgXfGSYaloCIDF
N/q30AQlXOVOdcLLhv5zmgYERO3J6+dABvJqW4Cvf9x7B9RR4ysFcqrgmL3/BtHKmW5CIWUIZzSs
fqoogzxSTvVZLwrAfnC8Itj22JWV67iHfMfnFH7FNWXDRaXHSqhB7vgxebGHsG5pPeZ/UkjP0A2M
FgdOh0LmY43NHv4ilrfeNWNAYNbFwopEG3tWTrYauc2YZc7zQRQdqSEso7ufalyJkU8XEh4zCfO7
cjkTauT+gKfNxE52Pdv9NESzyXsA+9MKkhLd9udniPoqldzGWs5jupW0BNzIg3CEkbmc+bsM1yyP
5SmAETuoc8XMtzlo3yWTxdikzJSqK6br2kzkZ2sEilzNkxYF8DJqmVuW+y/io7Tpj38FkAQaPZOc
5V5Ikyqr2KmP0C0BhNrSnOfLQ/lW4AU6OShkM2EbveGIB/+/R/iKxcqDFvYmnJU64N8v/aamb/SI
MmFoqdmL30W3uqGHziAE15/SYOeasMQIsYQNul6ZPLjj2y7Lz17Akattiyvyqy76cJw3FOB1joPa
D4EQKiG43wt/BtoaS8uD0x+sy5yR8FJYewg6HOGRDrR/uy/Ok5cg4t7dwXRbW/n6K5drkWHKtNl7
sUA7G5b+f68mJAVw1CJDqqtYp9vEgtFifjRaDrZE6gV/rQPR/p3BxqsqScYxNWMXbvIwFfDCmZTZ
lpOBecyZrGD/tsk7mznvqvLmus9vMtdZR1sIM+mW6uF94S3ic9r+xou8BizF0gfgoIsSEy1ihqpg
v52oBAlqnmj390ofyJXWhu1zpxb+8midfRBcDLZnVnLtNJa49xdzD9NnscFdaOb6vv1+ibAkLDUG
e8ulm6qAQcZVDvuOhQJSGu+ZgZ1J8HAXd/OsfVz2vW9eeXO5sh1ukbZcP4C/VbuofKErOhfi7XJP
3dZ9QuQFwm4lROO/Rb1WFzw1GCzoCFJNL8nrf4LBbZ0xgOs6a1NbHRHhHMPtAPOnwUKaW0EE2e2q
YKu620Fg1ileYRvT+QOtqbsFopQ2GRCdzBigsTvT30zDJQn7z4CmTo6d6dI/nMLrCl6LGT3A3qra
x9UmgbSy0tMMNX0rRmVijeMzQJVqNcY7fL3XJbdTLoMA04JtfL/rJ/EJSNHITbj5XFRECT/bzmam
pLYCR3dJheSjdgjUmJJry5ATU6lTZPkw4F/AhLizK5RurGmkoTvhhMPaQv0f7mf8Y6SfppG79yWb
O04IOq9c525qax5rzCjvZGFJg+HFqdezcTXvCr2cacE2ZaiZIjA+qk/+v6nFuxhfJfBBweSMaQ7J
JMRl714VvH2GxWxGkSYUgT0uQYxc3lapB7qOnUfoImENtXATRmYCb8NOOCFWhepB8Chrd3N1kjUK
cuycunjWmsTy5wSZEhHTf7EAYqeCJVkIgi6bcP0cGnBkeuXyJ6MmHlSVdlW1Q9cSEwtvCfVIwJ0b
u/ePAkobafrorNcIKCiRvbGt/i0hVTW6H5bEcTVRx/78HIBzJBpvSkyeT70o1JCKAzBhXS1IC06C
0Fyxw6UnYBl5mvJqeb7r1DLlgB6YBUDJhn4r4Y4rUprIuvgavq3HsE2SwljGOi5NZGK8BBuHH7bL
7ugFzUqp1XgOH8qZJNMiVA+HZTaKe/BDhPpKb3A2nE8SfZcQIJKS65dwmRBrTo4GdAcns6Ww9X5o
kUXXA23g1Wt5qUefAvU6SS7yF/qb8y4B4GGlYPZEmusW8tIUw5UJJ+jAqOAJMw6Jptvc8895lW5M
Gs9TbPQhWqmxuT0CtzM2YAkOyZgv8/allrl8IpMfd9p4otaRu2iJTitF+A3PEPEg+mSOfUAWtAks
cUThW0aElIffMc8qf1u8dPGgPUFDem3Q9FiUaokpKLxTovej4AnOYwQaHdbB6Zpf8gi07lGL0dIQ
n6aer7l/lek4lytL635SrNIKm+hKTLLRGs6uoxn/txS7X1jyb1XZRXAaleAYQSdEUQJfqOE8Tn4u
vXZOKF3y91XR1eWSBsB8rIzsDmmu0nhz9aL6/EWF+ZpjUf5zsTodDUOkx7TbLFn7XFDYtpM4FruE
u3vsgh7fhvbFZstOxeMREVlu5pVlKDduWmkn9nrShHGzQE1C9P/XWT+WpkJKXbFmrkzQWN3gprWE
Cw3nLMn0ZuVxxtzUKUfevGTST8G3mpvu3H/yezYoTNtq9De13NCBPuNHR9p92fqPdMjfrAZhwHV4
NMUQtNlFAXVoaT8Ga07D77qfw7IZHXYUtvKpvHYry5/SFwDkCVWdtVAHycl5VLiLN7l+0e/vxzSn
I3/Af9CDRDNw3cw3wvfDfS8VPiGlzoZIt9xNDmrrH+Ye8uoMQS6ogbUpR4+gV5rJabyeOxQgmxOg
Uo46BlPxWKA7xbF7wNHxy2f73nbT2eZ2IAvuHY2bpdFK4cZvKaatr7+bNtguTQwiQ5g9gXUYsJ0F
4N7QLC7XmiZf4C7sXrtiqH3bG36FCUP0lTUWHhEeFulrXfz7KErfz/4lAH+PrFdru/ZO/qQLm2oV
S4OqjLNivlBh18h/MWHuyF3T0m2spYBS0wkNgdKyHTzz5pwVcTPq1+j70y3QUSa6UD4NZ8CqEoeW
lonQTaw+KhcoOPmc/Z0Eu/SWct/wydGE/RHu3ehBelGFYmr65Sshpwxw1YoA3+GO3nBtrLAvszn1
gBsJ4qR7cZ5K1zLNyQt8rQMBIN8zC81BoTqsG7TMF/1G0dLDRCK2eZMnjgTg5fDGZhHRMBclZyNX
o381+/jz34WUNq09rMMvp1cBOOoDWXsLJYiME8wsst6Tsvn2Wj2qHlMSKf0HO310PdNwRW874j84
lWh2NPYcvZFCKnKr26FI2IH9mn6qeKAM6knnxIm/XRrBEkF8zecesc4sCgzigvQ97m6jBsMDblGr
HSvTeXAHufKiR+8zbtESsT8D22VeEW4cTtO+7AHelFQhy1a1KXja41pfDWGhlppW9gJyrKe0Iqa0
au1vPQL3/vWyP76no9BRYzywFS/pndiUrOQ5GMD2JqTyUlTl9Hd3zkcnxxST41gJA4l6b9NNdjpU
mII7t5L50HekOpYtiVnE/YvibxwQizzuYkeBUREo+36UQnlQFwoyB7e5I/X2TJYpj0HosS2L8U+P
626mFxXOSP4/N5ig1BAHMt02WVdawS3RQw+dJa3O3QyA2GOROfhPeBGt6yTreXnoyvFE3sP6zz3Q
FdGfIxVXk/mGHfV7Kn5/ygmw8nYHz4XH+ZNpkZMXv/qaCzvJE2oJmheRnT8m9jDL0yDHyqx+1W5z
eJ6bRufgNOXQa70jeaWV8dcMeB1CB2Zo8Qby3IxOF+Kuu/IW+o2uJOu+x+WtpT4Yo7fs8vEF4206
E8lgB9Ep0//tcccZEbyNfSVnsev1YLsaQRCf3nHn1Snfd+y2+zjE5Pyk6xd6C8w3AWds4On6BtFc
Tlv3cncRuinVWhihk2/jvNLQrV5l/B4XKRluQUdplVVcx72Iehw7DSF0g8PSm0PVvuVEoKmPXYHE
bt+ARLVgqNHP5J9Chek9EEe8uc4aid1aF8VT4LhM+3KZP07JLeNvC1LbuxhvowKL2ubE7nQEFVTO
fgKxFOcn5Lwn1q9q7nba+5sPl7tHhsGtKnj/JETqWlRoH9TrGmgbh6BWUpxSPguCOhL0EIZvy0rE
DMvAwp875d9DIRSx+/ylDncMmRt0CfoLVXABsei47Rowx2dWcUS29rWxUXMGBjCxEo/MgcHZ5aBi
34Doc/CRNuVObyJ84mSGTw+c+8KL6MCuZgqv8dmyIhK8plRMglXQrAYf/WnlKN5O2957RIDkMOlz
ux9RBcrBsQuHwQsytnAodRgx+ElsYOsJETJWBMalxOvMZxGSnoaOT1NWVgoSYEfkR8dT8yElRC3+
W1hxAidjBZk5PEGBdNEmoNuKKt2FfCZS2Q7YssCGA8SMqHWolcsS9WHw9kqSiTjqJ7wjfG7HMLc3
KMzsBWU0lKTYMizJHvzx3hI+77FY2V1tQTW5yo+cHMUii1anJ/us4B1zajnWuEGQUR16sd0NWQQe
UbqCyyAcDqC7bUiJdBNUP7iL9PJ4NjtldketUGjCVA08IRRsxIgGRZuVtdaDwn1RB1FylUI1/2q4
mpCfzCeUI+pC96wWJE4JLhCzXSos8OTcvwPtZFqCZ2piHCrJxkssWDu48dxVcWyrz9t129cFhJ6M
1polN2xZAUFjZRX2lix4AGbVxMMAyZYpxUjuZU2Sfg1k/VLXIf6B93C2LHucAxh4wO6bntMrjwAb
88KQeKUBLLKfsIPgh3HbiW9xSLsoi3otjwXdDMtNrpZlHa8e71QeDNxoHOmV9GL1Eh2ysMeOiCHN
bRHfHOa32rNNfH1IEjCVmIjAIXf+M7I6UOlrn7I9MpwLZABp8vv08sLM6R5EW0KoREka9C/ZQqx/
h1Is+rOJ5o9YEDADVm1RsxNbTb0Ks+Y4t2bwhhTC6H7wsCz5V3/3M+Qs2OeZntk3mu4nLkS2QiYJ
c0o2vCXha+aicijfjfPXADrJ51v+hWdljPBppz1e/8aWazsv/ItwRfgh/jF9H6W3gK/q4necryRY
EXr5ideWcuybZpunWpNyAsK1c+bi8OeM4PmJjAaBTY+Y1WmQtG/IcRY4PEHg9F6hyPOSQqBfC5ot
fW/L0/5/PyPtD+BENEKpa8bBJ7zyBSo/8ETPfd6dx1j1G1z3wxiUEqBgiMwJOSHBCZzYdAhZIhk+
wH2i/30eLpWLByVX/2yBj9W4vdZlYbzKjitetmZt4ivlE9lWfFjytqaaJxjWKIbj5CbU2ikQPLIf
1hpRNPwAVjkukroGGOBwVpbfgUXaIMgMDTqp3oB73IoIOVKFA3dPIcaJp9c3t88d+wvKQOddUaam
qTaM/UqwZA9iryURQTWwUm6IlFaAGOQSRbemRH8FFbBTGoM9EOtYo6GrkqdKvcmpbFBO5hayMYMc
cjPDg2KEzM3Hd5i+TU2+1YE39lSzXAapvAAA0GcHjOjRz2JJWdEit7/Hi+tDVuocLT/AhGl6gcj7
UJZNPCCftbjH/kXqpqZ5J7YKkGQ5qJtMtY6cvGa88+T8tzrlKR7l4fO28ETFtMgZSZDkwHFObd7E
M3f7+sxul87mGKgJMXlF1uGwG4bNAtckpMb7y5FT36gJj+QX+lTfiaK2+pxB2q/eaawDrTV0ysVQ
rNNUbs2X9TYywTgVYaSzQ3LeKH1CJJUQKuhINQhaEWL9kFS9vAiM0dobODgbJOe5J1VvzkbgsoQd
2og8cI1hxo/Rg/mhzQFx0ECCETxgt+Z5wRQlD/3DfDCAD2b4m6l1MYGk2ainvuu4sYv96qPtznrI
aRi9fx1lY+zNlMcyjyEsKjudNxi9+ZN5zv5ZkaV6mUtC91z0MxrBa3sBg4bHiPJJf7OCGlLexpmG
mhplEsXbzYxYvWipAvZNFg6tMs90HGvqeShzdp4Zb0AnUt1XklPa7Yc8037xOxRIavvBvVzllnZZ
SJ/YFTT44fBIL1BDDpata98ByM7WIUMg4QAhTMh2PrI+M35awLNaO+6APPt4GTqyFxoC4NNqyIGP
fTnfrPGLjVBmK9Yah8ZEBoPgq6dCuyv4G13kgM4C8buT6BtVtZqqC27ceZ70nZSnkb8BYioS+y/4
fqwSlYH3n6hvZVvcpOtU41IM8qb9nn5WtAwsscyzm2wc7+ehs+TksmXS2q7FSlDVyCwzGnMDG/Rw
EH0YldMGq7HIdLDlDjoSiNO8TLdwJzs238/v4MTJEVDAyRkpzlEmVGbZtPI8LcuJDBMssY0A89ah
eOgg1vfXf3bIYKKRW9qvdP9tZd91YJsnixpFsBpslsmF37X0b7oNtP88bcgN/o0RFbbK2IPuDBYu
gMqF78gch4eiffhxNYV6cmSMbqPXvZt8UZWG5WnQ+V86MCKwHuh7Zf0hzsmNdujVlY7sd1th4w43
3s9IN6WmTl9DTHUrhuu6PBfu2qw+22ch6X+VsgHSl+vamY9UFOQBTZiGnmv57EFJta0cA4kTqR+0
KohMgRwpkO3GlFBMkMJGXZPmxd7ZdrrEs42qEqpbHkA8l33u3J7WwHe+mwkt6juOqpzs/domZfTf
16dBFYnTy8wvlVLPMPPNv5ZQeLWSZsIxLWPox56vTgDI7SCOFaIjq5fEovQfoSfFljuqVeL7HOoP
P+UXUcVYhXn/tx4DiqoRIfRdPX/0+qnxgjKHfVEeZlrkFxB13S1eAfe+yMPOmsRdWDJlSkLojI6r
YE5yVXAF5I5UjAUTDxE2YIutprgL4C5SNX5MBhI9vBQJD9PhF1L+ld1ktixNKaIOy9I7WtEulnoP
bVPuHP6mXaEhkt2SqLDNbW+IfryN0shNDLsTFWMvGe8lEMk4BFDa7r3crI8u8MEC1PM7ww2ImIJ2
N1MLNlME38ow7ZVBKjzWprI3hklljGDIS9NVcqyqWmCIpZEuYq+3BNJhub+JQINVvmMU3DqvOrvS
TbL90i5u3PW8Mw2J26tDA0GdsYSgh24HJpjOaKQognNoMa/IXS5Iv79QpGx9hDvRKgJBJe6DSrK0
xM1SQerWef1bWkMK1sEPn5RZqJNF2kQFE4no2unA8o/38Gmc6EKwu9f8JfbW1pn2FIXsv/Ciqhq/
JrmXX7oGqk/+Q462QsZ6cxI55Nwe0UGq+LWz71Z+tBhFK6b8bA/69AP1cPZYqbzuVh0N34PAiVYL
eGz5ys/H1Pf72ypPT7yg0b5QjEvS3GIqgSvpxXbdibHIltHKECar8jzupy9p7mPn/xItNSN3j2gC
u0AQpDTm0e6cebiZMkDMos/b8divjaZdBjcKF2fcfidu/x8dm/kXeNeaOHalEYpQWPjIvaam+Hv5
R2w6yPsakHUaY3v2rIIyQ4miJHOtGXo1Tm2DkLsl/TqrNiDFN4jRJGQNyUrxAQG2eC94yJwJyfkS
PsTefTV6ykI+rw2VNGWSUznvu5YJ26904T+1eiL+pAZoMJ3389KDcHYaYHjHfsmho6C/Et6v/XaB
HslqJeiYLzumS3vxTp9Yhs9aD7PMmEm9IfdRaNUjGUcJW4liwIK/4m+lQhPcvaLKtDJ39z+Yf9M5
OEtS+Uhq8kYB9ocOJYr8rl+faFEDSB/7UT9zKNAapWr3ey7oghJ0rjzu/nEmxGCaJpOTvVvU2eui
UftcGM+ts98teG/3Hy4DO34IXpBZwWFrqJ5rJFn62NRJ/g/sfhxzovs/HOZhyU0trgbvm5SYru9w
XpImsK7bl5sQPaFjeLBMvWGL0Yg7E3lGep0goICuI4q04Nysc4EyKJu1kndg7zbX0vgouai7winu
DmKdFvpLONkLmGU5JP6zuLKjLX3oTT8owMeT4tCZ2mjcnkgKMAjyy1fcr5KDEEkePWcSFjVVu8wy
moSCsOwV7Zt0OTkHDALdZqz8Xrq0a/lHOUe5N8lulx64zjjvyrtLLbJXrfQ7tovRqbsjPWK0nOYa
dXFMIeF72qz+RyoZcsMNqF5FFFfhUS+bQ0d2tNUj5yTyVfrXb731PXzVdzuE+gBS+sV16OXdhVAy
I1YkJ53Kd3QmomJw7AA5FWywZ+HiC613Kc11QMQc8QiFrhzMrCSBo+Ns3u7/smWNkTbZrloV2g5O
xETrqEMeWwiIq+L77MNgbnwR2qXpmDjq2UzVT7S3PUiLdFZZfPRXxPZF2dttJHpxOEQyr1wVVI0W
e9Vc/2wDk4f34Jpm/On7NHfynZIUlfSoloNoAdBE8aLV8pZZGoQMG4mGCDcEL5BzqR092QyO5hi0
qlEi77T2yMcLrl45j9TIjSnE5j4j5H2EGt4p2YhQklPTuiI/BJxFlgCfot8ZL1DpP0nWM90bznDH
oi/ocqA6MSsTT5S/TILCrdu/AWZ7iDOsh5Dl3eQoK+gXA7Mq2a8JNik3O7z5+6AdGaaPCgY2qNdA
41GjH9y+KjiOGaAjml9fMEQjaj4qz7FUr90aqs2ct0rB6iokON7Ytv+76AoXGZiZYoRFuZT2TRkN
lcgcIF3aUakvqDez/4rBrO7U4jzX6CoLnff4ut/mqRg6YYw3l6IeIehSaoQErcB3nSufUEZdT40S
5msYdzbCKLyAPsydp8DN6t+vZz66M8rK/UjLGDuyh+UV6VIHsuXvB5datr+gxx8C0m4zNsX9PUQo
zXRSFdCTwZtOY3W1KkovJeqm8uyDDQNF779fOr/QGIcYEf47C9On8z3r3Zk/EshAMSVYvmU1Oks7
0wFDwby9FdjCN/gO/jgR9H4jJiWSJTR9IlQk7PShtMhrEPJ10+khGAWZcr7An+6UTIu3QKu4zkfV
0ycd9lwn13IXNw/3oVkAUfQ8yVbna12+cQ5UCfabbyrg6cVeAEVHktn5H2eE3/fhdDjdr7+Ot+mH
3iElwS5GkOnV01e2RhA6a0wZF5goINFJ52XSNeciZ4j+UGZdJ4znLG7goTUE4QKCpMnMdqe6l7gt
dYfrNy7NDTRbDAdK0NCXSINPH2RbMwblc5gL9+FN0YpA/lRNWkJwjT2KFD81G0W/TojRF2BpjIGN
dYc0YxSIU4tH3B5VBakmZYOWw9f8d/zW5p0EMYgRfOyWXJf73y8z4Yyazc3z/0+WPkKmo1A1E2sj
+keagTfUkO/zMOlU3eQeXxlrOfRdiOPG4GL4gbBz8grTC8XXmpcG08ewRdgqUnqOz/CCNlF/amEI
2/vd48+eIjuJFddsMC/8pp0he0PS0DGAtUCDFI08ruEGtI2JBBoFwz4ib6EVyVnVLFqXvIfkf2h6
hlVBvaMsXLihxLPqJ+eVWjdon9X/F4IvqAXHl6Br26n0BUtiz+RRXll7gJfWuqLIJJIApMOePbJ3
xdkVe22sORnOm32rCu3QMvAZtE6oZBY6Rxo/t6bYU3zCbXFcp4Q+ulmXpakitx42R/a6x74Ac1Vj
fuZXKED5VcHrYRsEA0IWLl0EtCFOGD0m0pTSayFjoeA3exiRGBuy+3pXkVYRKzRpWIurbVww5O1A
NFgkp/hPZ7KW4m2vDlynYGlXjCrsx6S7cy7ZQ9cZi1QK3MLu0EtkzZQcMjNea7bI9f+y5VwROwru
MKgC7h82IjwDHWpnPMOMxnDyKq1eZzqBhFqcv8hF03xvFjEXr8w5diPsxPaNnPhwYeUxG8i/K8EB
tMX7m/bBJQekD5KwBiNsBgaOqQgHC72XJ1AfHDgD9AS+HLQf/uxuGMMqv2cY8VZvN0BQOWFg0cMG
5qHC5+tjG+EoHncEiB/aUFqCRSj88vy/DcazMAmXqsJfA8vpuBj0zejIILgZtRAyOcf8hjV9ihtP
EV03G9cbf+c41vYLYRIIHN2Uf4LMr74A4z9UreOcRQxGoc86QZ5hHtXlR9GZj/Uy4ByU5rMvptQW
7A5Dya+3c126jWhzCW0Pvkrfq01Z4iyHq6N/qzEPs/2zcJfS2CqlVvoFXdWlz9t7d8obdJ2xZOJ1
gRa0i8mWwBUidvMtdDb+jNhiz39lkiEaGFa5+eHPy0KSWVKHZ6/Q3Ifl2fZxqlkQdAgunvMLPOFC
n7QbS5iLBiESUzqAp8sZEzWzJxEsMVdJ+EaRzsh3Nr9DmYErFQ1cY2fdE580mh4WUpGdapcraFjA
/7DWOnyzZyqNLb5AGikBq1rZSPqgUE/l9yW11LJ25CpK+6bSOc+1RWwt9D1mN76hIO5/oOkpGjGF
7PwW8iUV52nm2ydSneCjc2BB/1ibC6/OBlCVyGZJZiHBJuofLwwortjlDXh7kPWtzNNKYtTQ11eO
H/wSMblCH3f/DV69ABCJ3hwev4s/seURS/zU3ijTiOMVs8Y7QmGHHXKNgRjQ1L/IXHu0kwwLf34m
3UgJujAmu/Mb8/YvpX3uUgr+EAr8Un4AJ/vuzfvX10MidbnbLT4BcecrIx5gNsCOxk2ytoUjpLqj
FN6iOzmo1yvMQZlLZu2ynO3zve+MbhXt1iu6R81agt7y8UefM96rw6kgSmKCm6+12fxCx3O1sKmS
/txFllwnkiw+DeBnWYKBlJgEUdLg3Rlj959axcmQ4S5f23Cfytc5Npd5SlFvm27gTm9wsSY4LsXR
K83LzOWcu8f/GYYZNpkyQNvcWa+RBgKQ/9b0YnJg82gjOf44pEkECO6uNHbJcsyAhnyjyInKjXFi
vkzBh+hNFeMNe3wlKVm4WgsQphRyxyQiTraPHeMR8HOxyXpHyxqTraJW6p1kuMnnquBxW6FU7bLQ
2WBABot0Ho7W7/I4Zok8U5p5fzjP4FvEC8eSuFPNfwejyLbdc5EWGRmDU8cxdyqefypGRm/anasq
X6zwbQB7E3UoZzLJk4C1jkm4IVc/gPDRRolXk96u5OWr8Q44HYhj9k88Xo8MDeCVf3E8ZljsieIn
cYEk5EUKUJV9nCgkCaRC9sZVxdyyRIyXR/U4G3jZ7C5KwpBsvKobSHYVPE8JZiAurf3Xl4GCBy69
qc9OQLoYX6mviFdBQsukrEmlFd4t3rP86+gLxQgF7IXHDibWTvAfVUW/RQmGINRtg6HK5UnvHZL0
4jJw3cPVTY955O4V6iFnZNaEyOkMVLAaiARi95e2oVR/6XUndGX6p59e+CLLxsMgXMlgg3gDJhaG
Z38wEoKEO8xXsRTPq17GA1X4HNjvW54o4+FMYcpFFKKZOKtvZgn9h/1IG0fhxT5GPs5Pqhh9GH3h
2NJSaxJKWnlqlaZjRcz09tosWGdCIPYKJCmnkRAWtPkWismWK746j2jdx4H8fJ0qvrGXbUWtQl0m
piTukfRJvFq4BelWDEVB/N1apKu5fX4ny4I58TstG2S8B7rJ1UPMx9EVV/ywjVTIMoiqfI04ykLv
YsSVXa8H6kxrzrtonZoVIknittN+UaSbmX3H3xEU7btxxpbSd5yOJghBWDzf3EnwTIRBOPNvJjEF
FYDL37Y9djkZ+LXAEsIRLPYtloderLJpi2oRqMggV3FsOkOCCniJ+TK+VkEtZybaXJIwX5glMa6q
UtsO/pn9YBgtIbWU2QSQVIF77AHTyJrGSFSsZlfzWoBPoK49lLecQPTmUJtiVSyFFX0j/Xphn3nb
MuaA0Btqhg+/rFR+Uy/IMSvsS2Gnq1A5Sv+eHmgyvYQgX3Mm6v18bv7UWU56koAiKMdV6UWffA9/
Odi/m0tBKwB3givn8mNLh+Lr+++MAT7ltWxjdmSSe0bR6EcU5cYFbAaTXwQXW7BNJ80oQNkDEYe2
WmqFXUylAmgvDzku0tX/M05FVMv/neXIkSiY+PqqlP1JRCL4NdZEBM+b+7i3T9i2PW+sGq4NXTPr
jeS1y5NAfA8GwEtd6qOUrnWAQ6sFmqGkGmqZTF+V7wbSjJ7Bg2TG4urMcdw5ryZslq7EufhuAzr3
8GO4rlPQvvvTkABr7yDaucGGwOmLhuimTUm62xmV39xOQDdB8Da7WkClz/A9Cjr6gKpKULS9VsBy
DM4E8woeY5014bNoLdvKGxgb2CFLxJxwo/BdcBzm7QYypuJKzPBp7u6jUKXGhCaOtaxGSJFvZQ4q
7pL2Z5K6pmSQV3s4kRRTS0wAHNepcGJLn8i88u4ovNxJs/eCEYs/8mFqZ1odNJ6wkn91xkdVzCbr
BBj1pKw9JzBzdIE9lR4B2oBln1nmNjbSDBtuCFS/+Qh3qaa9ovm1He+Eyk57hXxXLMs0iLU8xXvq
pgwiOszZz8wVl2CglzYSMTDCUe9nPcDGwPODoLkPgkFuXTQKvT/qHfK6l+8rbKeIVZS8QC7//hiG
Z3OfQ6BuV3YxSkKYG8nWPhtWyOK1T7VZkkBuIp0EE/IGTjv8qS3DsdPQRdeFzWJWqVdiKV0HvDz8
3boTpwBbAa21qX1t1pBeEYD+ENKtj+r36KMZPsxXi3+V3kz9qlt4CM0c7lCkmLuR2yq9t5fZ1aOS
k4mWKZSlID0bMYDSvVBUEC1QD3oo8cZqMDWI859NOma7EFR7fjZgcWerrlu/089FoyBCZI/jmpdy
i9k4xBMB+5XVcyQBTUqZS5uuf/U+pV/5Ml4uCwaPpcSivv/pgp/6b9wg0+omOuaRJ8TvtoSguYYp
U9FqZwOa8w+DqXb6FvCkH8i0EpiUYMnPvmJzkYbir/GjgTbqBZnzK3gcLu3otOx9ezz41jdkyAcG
3P7icqoSccsPBBBS01UTyFlVFm+Mc6v823iomhYL8svmGHpYDsYY0pAHsXeeoGp7d1BQBonUQQez
arQG/CuxQqLTO1ud/cBzQCWa4KhRMWprWTFFPQT2bZn5IJ/kzGQpCWVyXvovimWo++t2CGq5iDh5
UO35lCnbV2olwWK5f/Tm72IMfxpl398ZiafGDF8R/3e4Y4Jkv6jVxaaflhlZgiiDEWfjaWL0I/TE
5h7sdIm2bWnOstq1JpF+F6sBzaZfqNKcUj22vjql56KTp0hFVDfryXpnyNDKF33SB7vsWyTQWyrp
MWIukq+p23JLGwLov8jN6cDeVkxFTgTVKfp6m7oR+ZRRdfxHkWmHnR6BEyXsWddzQjf4Mp+dRWlG
AD5yMPJjRm+qG+m0F4Bh4yT7Qt/Tk+M+zgS+wOQPpinOWteuA/CsWcX/urwge6Sif5Q3ThBYFxKL
p0LAI/pCgYFTIqVGDIs4P5iTcsGlnpvL9T2Ru32J9E7NEFto4pM+79gNIGInIfZoHG21pz/S5WPp
85osDnzU+TK+z5aKlb3Y11RKg3tN2J//36B0kpXhEu8VHMvXwc2+GbPtD/lHE1cxeE/wFEgm96TU
cMjMMPE15QKSVHWqrUw9Lyv5zLgRwr43V3MAQ+KbgG1ZlEx6mDcvHQSAYgeAPuCEYPUqK/lB8e00
PacIMxFxoEW3vyBNdQUQPq0CgbtBoK/3qgSmXt/StbAVDI7fdhdejecR1+IQc5pJsvBq0oCSEtgM
muulF2eVxAcgiI7qvHaHFfOfLNdK9IzCFj42fghBkHzOySGvkOhMEYjZ06iAsNERVSzhkB6pPfvw
7q5+OIKgndaBxlFMh5jDIhuUt2fEJlsiJ1E1v+ISbt46Fh2ipy4kptc8Fi8BCeFvx/26jaiyByze
lQO+JFndzSuv0YrgZXQbU6LLJbD5c76RYveXOda61hOH9Z96aUNXl7Qvurd6r6UUJd42Q2dsjQ68
AVMA9uDATLGUGizAuC7kWrIvSvddu8ZtHvxhVBICxXi1SPK/qsxb0+VZ5beamvpFuHVQun0OsDQh
0CXqj7rWf6rZlIflj60cN1NbLoghUt5Kh8Gkb2LVKM5vDiFPp64rKtl6er0ao/rb7Lz4uo+Rt9C/
8bJsJGcrKU+AChRrg4rLVyCqzuExtTIYKtKW2FJLGC2l6LWqNUKPwv2Lu/+4uxZEZxq+AuiOU6ZA
ToNEXwint9Gy5ZiFR7t1UAFN7CH7V3csPlBauyYXFLwsGLcIAw23vNoB+HqWSLXkdpAc+J3uG6V1
opkOK8mCo74kkIWFwVqi8ZyfU/nY/JqklooatJ/X+cJpKZhhBhpcD9Q50L8pNdzcCoMb33FI3sak
gKefZd/jWP5OP2x1NiLpzgMIQaTqOBNSyXIjMg1NzyB3ub/OR3/iHZHaZNx2TY9iT0Feu3ozPIyl
Cyde1DqO83tXWhujWWmIc4BI8WKuJyozaeDjb0LV9f9zC71cJAwX4QQh+kdYFUMzQ2VGROCNeKOW
NKVv3JrEY1BrBD6EERspcEt+fuZQyyDFfmaViHbKxykpWkwrVxWM1jcBzW1JHdsFh9w6Mp4LxT8z
gyJwY/YC3LK0/4wB/l6qCriXLpCLpW7VUX2eal87gULt0FK+3Z5OEZylLDvlivvqAVUBjdJ5H7vd
oStRO9lXbHrOXSXZklvP8YT3/A7dO1Pr07gYnKYk6xAX3oSzilwPXj4YRNPYgoEq8ZcMlYQQytcv
XJTx5bo3kp7OU+EGMOjrCJui/9PXqPLRYobC+iFNliH0nOIguHpoy4H8dwxGPoGTjephhJpYXvL1
oKpikprjOAcvT5ZyiJiY/MGqwu1fl0p24P283SmshCj3TraPpbV6848TonLNL8JAJaMs0ReCUJgv
1c2UY0gCsAXRpLux3+Wl8H9cpLXPFrWlfkpRh0H7+lWRK4TNV30QKedZ1nxlytaQUGZJWo9j83rA
qvAHfz1JnqpSlHX9WtLHmTIwcvJREJb2+eJQSvEY7z+Z9sjLTD6iw2S+1fongZca9WBN6AMsKdY/
mZ5B9Ov6NDJU11keoWDHvOD8Nu4Zb6Y5KZ14vyXGluEQII234vF2LrSdzl4myIZX82Xy2uyA9D6x
0Df54vOxGS5VEhwmMzF2JlecergcUA8tta50kKIulY+aqTZJeDjl3NKl5w5GwrCOnKWUVG/MZT8f
6FxmkN4UzlEUCaSNd21TnDAwslfR471quaqrGr7ThjtQa0oHWe6ryo7pq/6MROzUd7dRc/1NwnEA
FgObnrQmGRXPwgUdg1Xsw0nEW+ptY95vjzuufEKl9+21E7DqgnKXKnDvaOO2n7ZhDriB60W97MGC
lezDi3/y3IKK+fs3TIeLfEfZ+3J41ZlGJ00nN0nHiGerrQDynkXTO8LMnWdu7Whp2cl4Hd/sVeTK
wA3txqNdco4OGueKltYauMKvUw0NAMsxTTUbnt49JBRmPS6my7uiK3IkEmQyGpmsaRODmHi0wXQP
NGcfX+DWbV0XoTGRYCpBbwzV6liTH4TiG2N3DLl17P76O0+/xYKztcSbAlHSf/KYxH+X5EM9XHZA
lXM8nkTTFNJHg8v2YCsISDbAoUtCLpFupt5GrO93AIgylKa6uOasNXLM5tiJYy3miJlH1tZnxqtC
iP82puH1c1kKFogvJzVt2qC3e0VzMecbqx00Gctt5a12/fg4yzowWhpwJxOIBPE42SM221pq8Cv6
8Jrg+Vy69+E30dTo+dkDk9kHLx6fMDzEBjkqIVieA9O/uv7oidp/XJGiav8yFL3UZ/eGl8ROS88F
+AIWFCH4JrJ0qoZsgqRqgWYs101u2CymZKsN2xtHWbon2Pen20igaCuQO35Z/dkhX+34c7Hjic0p
znOqbDyRz/aKPJvjTHjEwuCDhdT1sfZEwBAtFVRdJivHsa+Ev09FHTGJ6O2alOARc5vPsZlDwigL
7mXWqC7+oUIpeonHpS1s+fc3fs1yCsHgaQTG4Xj+00Khb3BnBulPy30w9xftL6SRPhsLFGA8Cu5w
AkQmg1uhzFcIsKzLcncn/ZXJZiBQpm4WduArwb6PVt7YhC3785eyiaV4UFf5HU0KffjIY+r6/PvJ
MxzYmimSkY02ybOZIiqIEYMeN/1aabHCFxv8f1PAyU5NN8vTt5jWD4BXwftDV4DIR3QyhKzNjMTy
z6zsLaAtwOc6/gWk2O+BsS3Lz4wfvM7iUPtWl51TG19HIoJciDkf/9lb0dniiDxAW3dX0aPUPvhm
jfn/MRt8QkEEflMGLRqADPTmq/hL8aFfwxeUt0cFq1cRBVJSMd5+r9fJY6Je/XSGKF4B6snA4Ngd
7JbaHjslF9BjVNRdsuYYaHtcJ1OmIdkXYBxYisjbVDOaG7yg+9T2wAPGgKJj69I4S4WIGuWxDHIM
JQtwvssfAimTp14Km115qmTi3UJkC+olH92kys9FseXhtGP20BwneiWDQzm0T0I35HhFfaBwpZJS
FSyhoRs9yga2cMCJrEwrDVhNw62/nWhT+5HoLpdOrrJgQ7zCUn/A0L6OYCJ2oIqtVghu2ZTLaPZX
tMFZahVvSjDMzklv5ZWQFtWHsYWFVyzGBGHvXW15uqgRafJ+lSysXGYUV4qMjW8tsXgj94y5xtRH
krL0Db0oGba9m4ZeuExs337KtVoUTSrgf4IP1CmK4RLNROO4HbI4TKCmbD70a2d1wkRl3nUeH2L8
4vc7OQqBTVJNJkaUmqY9UCWdqSDoFZEn2mmM5c6maR6Px+lqrsVYWKGjnvteVYaG9NgKXAQwWqQ2
mNDtw3ACz6RLXsbaez/vNxgAZSiHA2EGBsVZZDLzyxfabbyj+sD7H71Xh7yqCZgykOtK9NOPlEtF
nx39ixqGu320ebL/etZunPPML4j6eDys61R5x4QAov/uwy4OmBEks14L/+zX8AJ49d9JoRn0nxx1
cCnA8G202pbXY+Ro8v+xulTrvBwBS5RSY1n25xBbe7W9P6KKBUA1m1J7XJEAjDy6QfKr9TXDs2bK
xtbpBciH/IYFx2cTya/uJomOZf5mUokDsnaDlQz7/tEVLC4sJchgqbEMg4IM8Ug7v04VS1OCbkLF
6WQHy2G9MC1SwDkRS2LRfLyvFq1rkYQM8PhJ3xAGzGKYXABWyG6Vgpyj0A+UqqyEHOQ+5+4A4doT
dX9Ut8HIdngQNQrLFlptLunNlfhpa+gxtZCwe2XQBhfZMwyR0/MGhBZLJzqaGAT7dD3AhxbAHTZd
CsfKwf8dXi0Wum8n5o7LBIGNU3Qx7vJAdTGHMTwFQRGEQ961PiCE02UEaAlq2yJ3E2Q3pSbhGsZr
W0nTZO9nqRT9A4UVFd3CZATJnOZqxbsUzoxL4I64JsnW9bvR3ytNXJeQQVzA3gSghKdIjN26FODB
PdgvikI3EvCTjgQuttct9f4CNpYZcfH98EqSFLSXtrBXYj9CKhiQoz1Dd4qsf7lOM6nxDdzrj+ro
2W3TSGt9FALLoUBATTeYGChKRSyJEOBjlg7NE+XjChH0o+UYZF+nG+SPCkazefc6oBdz2Un9e/5n
RpP9S8/EEgR8rJQFYrovG1fphHZWa4t3Vh2vuvMqYlHhZjswqUjGBFAPEwbh/75DDznD7K3IR7Zk
U3bHewlKIu8sTEyG7Ox4NGOxE2qbDpJLofo4f6eidn1sihLtRnB1HNFnMMkHMOvGPgX98LvVtJmd
iXNcYt2JOUw5M7JnmM/GR5xTgK11Bl7ixsEH6TlNhveOEwXtdImIpGb2KVd+k4KGrVlvOzmNUTnY
g5DIQWmj3eJb0LCkce1qR7wUnUF3pv56jylZsBqAZnJSDvrOq9hZD9SXaT7WZzx8YbERolfISKI9
muajs/IpWCxj/iuOQthnNp5TkVfEQYd+AHn+/O3m3k6AlsNFFIp12JSFcHLzfRuo8IEerdXEsOY8
H29qdMBWU/A+uv6GXNHaRQxjniLVM3pMPk2aG4zdFpRyMsJ4D/iv1Rw9JI7EcdxyQPOJlVIzy8S+
QwEvF/Svr1YLJWJETHIAcbMt5mR9etAecWb6wlhnzuaCUG7ua8RNSgqTjghr/xkWaB8C5WNLi49q
g5Tf6txxcy7hB5AD5NeuKIDDOwJ13s4Gi3/db+xXBPSR6nCL/Bl/gyJEe9ZpTo4wVC9q6eNGIWaD
PAi42nlCQxsVuONpO7uenKLBsbUrDm0I1Fdnbiz0M15FjYQ18CcZNWVwWaq8Sq/wQoa208dRFkhs
TWraMnMC2lSMOvKIf/AXNOKtuBmGLUp+4TmZOBn90QWbhd30L1ac4Ul2Adi6IKrouUuAQUtjOqRq
uE+kArZRnUwqyZy2XmOnlmafmnNYpy2herYLiU5IfiqJGHr5VTQQ350SlcjUBia1cTiUC/M/+x4j
hlbdEB4wbRjOABVtGkc4VwhYu2jyp/+swUrx2/fECYaX5HM9cfYDcsBWPMzodmdziEtxr80vMDyh
KRanruhO8gIdU2rYWUH+YaG4eJXtEmo83fkP4lCXNlk+dDGRlSpCWjCQUYvuuXi60DBUpqDKPQm7
PDo5Czp0XTF8A015/lBJcd1fTsl424sBD0L3frRqQJxA7m3GjNgSjrpM3KoXDaNXIVT7Yr4YhyIf
bkid8MWN6iSJvzQ4v82G5rJfHHeW7b61t8bjxF/T6tNOB2dEE7/5rjTvuT6N2up3yhBKB5QzaR34
tUK2oGV5xIB7hbPzKZnRTnBqL+Y7hbM5ZRx1oOqCK3g9lzz2FFB4TSnnm7YGgmtOFjQYBdC0OiKO
LumXoG1vcQ2JnD5+A5UjX0ikNtqes4MUi0PqF66S+xYAfOfxEUafoLLmcG5jX+7vwjXp8K3iEFTk
W2x99Vq2Re2liuaMAG0g5M/zFCO9nzvGtYXhWh6J0ga5fy2AER0yegsb64G7Dk2A2vVtEZTZKhPo
kHRTBvmH00lWBFQJFtRGjHfXI6ZtAcY24NnKTcGgArHKM1DqGljd+XNDNwwIxEgHwhiA96CiSW2k
FUHrajxk3g7Ovj0I0SdAHcdl5s1dLwXrxvwtx0MMBORXHNgAkC/X/7z4HJoBzUEV0mf7qiXHP8rr
ROHEPFYNDQlXhCnu1o7O8ZAwiw3V0ZySTdNh20mBcsbOsb0anY1kIFHMFOT0KCh/LYKfXykBs3SK
saG1cuDd33PvCP9575tevR1hjvuFT//RMiYNzmWMSQ4R/W0xOFlBFVJlNZ8v6pUVr/PA0ZzCxCwR
rHQYeoRcxwtX7fWeONzRF7oSdnIZHP/0YazaxLy39vHKjUpD8Ht0Y3i9bTXuWrUoNFnjl9F7Hu1S
N9vPFAy3inmTGObW0UWlScshl9mnJZdmxGChUylUiy2UoQynVSww+5o0JYrKgru3e0e4AJaLxHPm
RGBnKK7NH9qPXkZvXEOPmxT8o9yetTiwFknlDMfZXGMxROftwDxPqvpISpddKyRSmD/gUbTdthJk
xzKPHXXHFJ8NkkJZFNU7IA8eQYXYM88S3xFu/hAKEOWRGfOn21WDZDlmjSZaeeZMFnu0048tO6xV
Cex+ZdoGxmZFOF/ZH5VRPSz8L1HzMP3zDpQws/B4X5Rg69OFAEYEIBQCWHv2LE+2emSQQG1bX/3p
/3CIExcY7SsJIsNRgty+89j4vwvsvxQCHRpsp2r0op2k5YlzBrfwWFCaG+wl8vFDMU2fRe+xTnQl
2fA+xMNnkJf9y7FFv5eaHrCLsYrplVijulhQq+ytX1T3pgqwP2/Xzvq2qnchjBAmGZPGCPVyG1in
gTEn/ew1GYD56qVbsS02grT34m+Y0ycp0NnryEGaS5PktDL/N/fgqvsft/FmsOnnsGXenF/jBOkg
fja5SCeCoZTc+owdZlXkWtELVSvTG4q4s7RzsqnaJ6higLmzuasfHhV0cVbC4fz+MxDBzzjEX3yA
O5eVzksPvW1bSO2IBIwYmBxSJZiCVGybbmsctnyGYCjwaMzP/NyLApFCGCo08pFwvfq6Vk567cnO
NVJj1QxXruo3aKcEEWsKlW/L3HaP2gC2542Or424hbpbmDFjGsHs8G/ZLkuaOvgJJYVe3o7SK+pr
kRa15Nf9Cx1kf6vfLPlWKB0wAJNCW1A7wA85x9pAu0LiG4dO1x5CmXVung0lmLXDRoXAMq1VgKJl
OK/c0IiEVzwQj9J8756+CvBEin4RgKcOpSdPoFS97wcTcKOLhuIXZSGOxrFx9T3X2/0AOUePyLVo
omiYNK8lMrOXEZQJH1YJsjbDEv0t2f76Fb4faAvayMQ7ozBAytZEk3/f1fPoBJzmaX6aAjghFlHK
MRvXfpVPSZrFRsmjXJx2QqbNw6HS3x7iVSKAAG26xCC8xf+9J20u2MEfK5SqwXH4Vqci/A3Axub2
WUazCCW2br+BOQ2hsZwnqr26J1cmOW/a4axmycb0lHbAzOtULsHXZC29vmWyxmhKdAu3H9PjH3mn
piqrIDK0PVruR/HD8E9dTutEftqutqsAU/Cdw4Z2E7/xgMTPZNBxYaAkqsPQltoIC61bqwIsIneW
+hHl99r0gn5z4JyiH3c3v24f/w2py3QcnG1Bg07fo19dSFogLfKWcrdoX6lIBfnI2kVRPae7JqdR
oFV6BMgszPPes0TkKPBOoyjnAhvNtPRmoBxTp0UAO4ctpNtvLAzG+Zo1+wzoXJ1pijk2pTjLvf/e
hS/mRjfHdpkMWRDnRPVEDzepJvEltHsz/18baDviwxn6GYKWCNIUPaQBL7C6Whr6v7p222xMJqqc
1ry3WlfkhlyGc2ab0mCluBhAbbyQgCvUMp6l6CfqCqXcyeReDM7uXwsCTIenUqtybZzckN9blYOV
h7bMF9/zKyQdD4XLrdsnwv9K2JbWp9lyaiSoTgOa3fjVshJDPb2x6lERKQ+FL0xfjG3Ngj1qu0av
YVjJc4mkZWsKgmUxp9uyzwbnwNT8k4sTvX/54iuZGbMkO2Ln3tV9arSGt919b1ouHnAzce1Y8CUf
o+HVnN3BYbzv4tuyEp7lb16U+C41LSpq6G9F7rIDP5RuLHBTBXMU07tE/ZTmSJIykNiS08RS0Qvr
fcZGOP0knnjlwgO/8CFsokAfAkpBnzpw04BNNOEhZg6fhLaZANrzdv+n4rMZeffjc1nx3+vL38DZ
JsqcObQU9cOTscNOPu5hkqfs7QtQzszqreFxKxXFCL8iYfmZrihoUqfODad46QjTgR7dZHyoBnSc
gcj/K2n2U+0KnqHAeUzHpFn5pXzxJj/jENzLu7G5zZBM3mucsxiJPhnCoR7nJaes0XAQZzfFh36k
N/zPxx4YNIdrdZc4qS22JH7Vf9wNWngrK6EOpUnUFNQfb9BaAUQPM7dKUj8JyQ7LBBc/JcIqpmNo
dYhLqUnjTN30sb13fC9pFTWmALuXVh/bt8tLtuF4WB01arRjKrNEbjEKKjPB9ugf7QWUwbmirTm4
wJOI4yJEMjlYzl6ABEJTBLOxjBerpDiY+Yzco3jagmQHn3SSt+Tru6a/XjoeInhQ/48Y5yb3Gymz
4qV6yxI+/ldrMggAHZmjnHpc0tDrQjLO54DLpNdpThwB9MlPI7e5paHNZt8VcTUq/lsltXuG+/l4
Q0bABiciTQ5fUEXQE13k4bQcGp0Fg2LgY5WalzDjLcnNX+jOkzgJUTVIyKkYb8YGXbRfi4qLjB0z
t7tkkMWq51plh63xQNU2jT258QihABV2etqwXfYXivaedkr7lJIc0nabVWE+5mCjcxuvwmmM7u9b
PqxC3akztk5ylQqcr/JQ8djnmBdIQaEceCFTmqXgkLXTtXVOINkbCt8OCjzO6OWiTUzRBULq+si6
3v/8eJYo+LI8mBFpLbB22KT28b7LOXHe4S282e+dPj5+z/uVaT1AOQiHXIrG3H40gBTwp0bQe2GN
NzT1pnbNC4m6C6uedF3HzoE4TucS90V78H94I8T/AltMMDZdPQ9l5+oFlBmtVwcRMQXHFcp7ZSkR
mT0Zct/cOKQEJWoWtWPvo4WmPgL75J7QUf9fTVP1GCUeC64g5va9MrU0JuGzIwgYqSj2JN6TfFT5
UjeMSrVB2kWBhX465m88b8Fn9Vckaw5bUdhlNZygD62Y/FiJwldKp1PjAojXfPL1cyRm9c5d+F+w
cNgIi9p270glYMEq10zhpiw8JsBzwhjoZvYYwUfyHt78G3NP3KZNpSJwzWYoYMgUHdDJzoC8T2cH
SlQ8CUZxP/Qzs/yiTGUbEQZPu//A6T5lyZ9PPw6o71iReSLT30jNycucsM7SBmKuis8P54dA5xBP
bheynEtr1Gg/8T6bijro/pkpLqU6f1SSXGjZFxagpeKMNspA6By2e5ECEYaJhiRFIR2Ar8OpLYCX
1EFt0hSeM8a19XOVkmq5mNwfy5vEXabu2AQe/m3CVwiQt4ZRQwWf3+/20KbIHj11JEC9RnLR0+ii
6nOxaDcnDWgxSkgV5J9vxmZB5GFTat8lSlIGqIuOTfhVslMQVuyM8kXkxT1UhjNqgRBKGV81ejGA
5Zwzrc7rdU5JyB35APENfHSXpIaTbNVIpsyhhaB9Tku8HnTOBNp93jn6FyefG1ctRs6pLjf1ZVoN
9aeL/ZPHlhOWX3GskPefCFbjiTWKZQXAVQUFZ/ChtasrGjQ7W+p2Mev7D2GEBiQqPpHE8DZXo0L6
FZJvHvmAgUVN8/pSEIAm05FNlJceZiUUV2TAl8q+PWLMEct9jGubSiDgSjzeFHU5zyADru1yWFAl
n7SHBNey8TzqD3HxFhhZChAS9Czj3TLgG6YcluR/e5jN+gMBlLdY3i0zpxnvtMUMYoFo7tmHn2f3
SVAC45QwmWiKw9LmtF318AFZ5/7LHMlUKx4OBIa+f2WeDoxtSZ9DLQs+xlGrBJFXY1x9kRtHCL3H
uPXX5lo86n3A1eFCNjZwn7dYoBDIshp4YDNBoi8kTAIaIHYw6s9X9sWOpBY3psCiNVH4nqNz0NKV
dJkjwHxAHiL7F6AVJi3XDWnpJc9OB2233u9MARmIRlt8NKSuI6IOgXiHbMjC4Msak87m3LyHJDnO
gmtA8jV1SDiEQbusFAYa4IafkZJ5EB0HNKazRHX0aBtKUM8Aohh4JCZbR/Zf6hlKf9t4pAdktB9Z
SbPZUG2S8+Izq7Nr24vOMM0RVauMo0q/oyCCJCW/0PTanfYA6E6XmSIpsk4+yZHcnGgytmFLopFI
fEvwQkrty0OFcvmWpMypsgabbOSA7dmDjKY+O34QAfOMVTkzgjyPqf2xpDr7Pw/vFk3WVlu9nFhf
4OnF2VVdj0YKZXFy1XgIO7s2ElL5/6BVfWcV4R+FiDJwThThJZpZUm4gaLT00v9tm7vb4y36CqdQ
YEOX603r1EXE+eZrOmkKm1gf+UBP0WHM6mXfSQwhB3Ov9ufHey6mQGDrGmirF8YKZ0UPaHuLhTsl
l1tb77ibC0+Vd7uqSCcIpOg20ZvnQ516nkJA4Bu6hxfia/VS9S9cBXXJrWrmixfCMZKEpLgIYQRb
S/KAmy+k8fORnOHjpKmq+8+8ytaF8qTHo5n1GaohWvp2M/DSj6PKB1zilLAOP8WZcnxEcLi+DhUs
ryrpZY2RanPTkb5BTVk975pZoxKvckWc4IiV1DNlpgtWfeis5csVwnNCB2vF9vgsYQsOMf42/R6t
VVBJHj8B/n57fIkhH53FBt936DWFwmpERYr6j5G3lv6PH3YMsgpQq6EAYAcYrXLPh4oPoLkLVqDP
sEfy53E5cd7IBVZLuptbuq3L9gaUGVuQ0H8+NGcpVOvtVqhIHFYPu3uK/vnTiiqlTT4QiSnbwYMh
GEOHG3tosmQQFf9GNFIle4w9fLOzDCDso86FNjtPQDGVN+lIdueyFkD337jBoboLvKoSz1VjTw80
jWKgZ0zInpbeYGSBgQu5t9ZrKA8pA+yYJG+sUE316uMdi06TAd2w7UtxfnCV5Rx6UaZmZQ6P9xgl
MjXSUj6IJPPy89kJf2/BV5aErbeTmaxaxWQcfv5H9AAIbk150qoeg4peZsbF0npbp5PXMGEYW/fJ
tki14jIqxqmgv0zABH70U2CpK/6xbstnVU2gatqFmmJUDPA89qexRq/fh8B2RXXFFx3mQunFF2fm
BWUlrOMpqxE9zU1Bw0RzVFP5P7H27NAtkWszq3rrMYVEo2vG2EzTyEPYVPT4LsWLckmsWLX9GnMJ
jGWzepOTwcCwoIG6b4JJo3XpvUZ1dLj53U43s0iXhmnbYe/HdPZkj2U6ltLnJ3DYSEHnuHIvMoPF
4sJEw8JouwpwegNJwUzBDpkqOmxXO1iz1TTjnlxz56wS9kL+JLZZQ3N1nhEITRtyQ1ul7qM8Tkas
wxXM+fxJQeD3KGy+TzVb8t0k5Frs5Bi40JrQzQa8VlCf4n4DPMGcs3bdYm7uRA7I7PDJHyOQ6pr4
5ULRYe0hNSDw8INDTyuQNg3NyugrBkvay6lZRczTKCLoXBqEcEU+VNA8UEA2jAxYQCwApDNGIFVe
uTzMmOqa0WJIY9EyPkYbgFpbVjG9QD1VTIroajh5S8+QaBehi9tB654W8e3XgCoyiG2azMW+f4X3
W1fukrQflqiEoFIIKsAiOvQQv9OdX2btwxnCgzmQZNlxDYhcqHSfi0Ev7WcTCjnNTB6ugmW0memU
FEtwedWT2iaXBNgeQ1WsfMKwH8ig8KkYNyFbAg+r5IGPCQn2CnJ42ffRRbS8J1ydYNNCv14jePkw
8yIvMNizuFpcC8o3Av1bpmbg94AyMUADjqFdF7/hg0Kn8VcNcx0VQzrZkmbaWTq4PgX99D0IYWE0
Bg1satgPr6IXtuMxeaMjA8NjnszDs2AcwYt26/eqfJir3PFPhlvEArwR7m4GewORhw0lTixDGMM1
YXhmcfg079ol3UmqrmEu/FVYZXvJ4JKh1+cpE1bmh5qOlN/IuPaIe4Lej2PeOqGAcPEFzzn5YqOm
5+2UaK0Jz+xGiSFKnRHhBOg3vCkryu6ViLQDPzoqrMy9tUljX1rZQeY+KB54HmuC6jwC+SRWdQky
fPVkiCZl7d7jvKC2kL1sRIy598mBQXkcAwe2+mwQ0zQ0SYDaOEDdhie8F7Nk/y8R/FH7ueDEuxMd
l9KVFlM0G8V20PXTGeu1PsxrLB/pMWpPGPQ1AC8RIYVh0dBOAdYKRgN23S1IdtKf8tYwynfa7vdv
mcH7wxX3hReWbVKlyF1zAAN4LL09bBqVWgawS2UGemMXYD2ge8EjXn9aPs3HuBXsN36QnYpjKW7s
uKSqmfCd8G8/eaMPQ0qt+hoFEOU+GmNq5erCTlVipTENUWsiMCl16dN/7hlF96ihvZhJc897SZsd
BoHkw9xvl6v7fzfV2s7kgKKyDESzQ1F0vpULahunXRo4X1XYDJROOZtTt8IzTVKnhiHhmzUesd3w
0WsEuYWGvn985dhsXb4S07tSCSRRnSnXejc4V54Y+oaDYhqG9xxs/YrV/J/9TCIry15TrzCu1QWg
7lpWi+ULWzXN8sVPTeSpw27jB9p+L8/Z+qjcPATlZZKVEJ5nb6vy8lj7qBLRo0SPTPlxSJZt5I8w
YF5nYOlbQ3ccMPGl/SXGPM4nHX1Y88afXpQkUs7wLp1ZR8ugNivNryF4OeLdE0qWNVp45JqmxcLp
BJHYvrf2brsmavdOBUwJsAC44gSdlOZj0OeTT2pEpygVYj7BkLAqdJRliWQ+3hSrOVW6EKxf4xbD
7abSakOdFYBu7B4Z4KzkW/KYQ8Wv5NNJzUK21freY1DllDAqnqKe/5dZ9G/TLWjfek9qQlbYeA5s
8PmW44YD2Et8ylhKCvPTKFGWd6ytl+BpsocTa7OhMgHTkv6FCmBvgqoElMQpEsgjuHWIHC4jqm6P
V2/IpC4bGIOp1SiNze8Wr44BVClkeW1p+W3REEg+rvx66s6PN+8/tezcQ1WeraciMG2vxOuu+j9U
htv+ZOMjmqfgOqLEVoIXDy50eYQ289jxKxXPEZs7zb/wzDQgAkc/KCJqnCbCbRXN8pZeXh4B7tiv
fEQHH/qe/bvDhFnzof9IS5FhEdueeYfumIUDsKshTBWPMyEOdzhZ6aRNMmHLEjlkkowLfIg8pmgS
LGhlH3F3vHm7MTUwtRM7Yv1BeI7MrmqMor+0e4ZdKgUb5UyDPBwQSpbpns6khorlab64imo3mnei
yVL8Bp00P/nu7MBMDzXClZpDgbk46F+UDRHLYyv6/9zbOS4flB8xjluRRGKS8dwdExZFZ6/D6Orf
xYKV59SLZAl8Hhy/7Nu+BeoKvbcATctDN9q6MgB4BlDDep/N74VTD9X+5TibuZgGcBmmSMvJYFso
aQg+AqvSY2hpk1mG2r7ffGof2nYOdXvhaeayKtcqROvaKUwwaVyq6VdEIRIcJUyFQt7z8CcLg35Y
k4cNtY02u9vpmfVBkOH4xwfbaqkH+SMr/iOBb6pJxWuTHzfQq5Nn0CuHYwskNZa866ZZXg9VF5sW
720+ru9ph7zfG79qCn+mgAanEFGnYVDjxO7bnMwpJawDOqljIV+fB6n8RzImWz/DrnLxhye87V0F
LYslBNHQGynVF2lCn8WSTH10N3V26HjdI48HfvhCy+lCkcwJCBHjIZcTvRSfjbvHdAr7Rq3fDZxb
xAa0NmtCvUbpztR3QunMR3ey3KWwTxJYxkEQYCKyfxHm8thdYAU7cEYp6iuHaKp44lcO5O+fICX9
/f067Fn6klusmfnPU521Z/ONp/xJBVFX1gvcK0ao7Qym2eXjIl61tSGEDt6+ltePNgiWhBO57BnM
Btw9yb7UtT972/mXDMgdhmTVw6i/azehSoWm5i8oKn2/tJmcNnl7EoDN8ePzw4PZGnfz4LL6MSVu
imKvsYK2LKgd/0o7YczxpytTtQYQ5gsEZVXY/PGDG6K9/D9448PRCkav+/oEmkSE8b0a767FrZUy
vumR3IyGozvlupUGn2v8EzrxQ9sH6MlWe/A8OYE+9ZaB1y7DM6aDtYpuNw8HKVgnfKgfJomnKF2E
nQpqRFamIfl+Dp9adqYA6YVKxaVWZTDtT/uJvaGCLVWY8dTdAWVcu+Ythk7vMdhX2EAVqWyOOh6I
z67NscXyIJpY1+OmBLMZjNp+ofQU38eyFZVXO02DK/f9OQjtfcfm8AYlJMALNWIqGqnnGhOC5Rt0
/ZIYZQi/8C5Z/z9D5CJQvNwzIMipJPiXYrXlzLS6RoU2uzRw49SQFbE+BRHM2yLncVt+szqg3KfN
jVBP2ZCaU3qmVHGM2oHurgV85psrcps7tD9l76ER8NVOuTjLR4mM58QA3T4Rz81MrQad2f6ZL1YQ
11mzWBjW1ytVpaHAIB3W4QaSBq+2SNSbcx8gWW8DNJOTfYD0bdIR1WNA2SeThDMnnqYClZopRQZX
SV/W4vXgMp7JAVlJ/tmK8xQWxYmzFb5A2A3Fw2yy1M4zOdtAjiMd8H8TYChIL6ZzWS09mFBUrcIM
AAcN+zX2Q+eFkv54/ojEvp6amATObuV1O+/VhgArV7zbb08KYvdrMvx8aiuRHtIjbBUKNeISWl/f
Kg31B5DHD90afI8AiGUKNMM0Xpmo+MyeO1Na62LNXCIOilf9QJ7nufg3WKY56o6HIYJpU+5cp5zL
enzz4ZLYC6Pl5FbzgofS6v8NVF4oZ9fOAFjFAvcJQaIKAoPA/7IhxCZIrS4GaBrj4UE0m0Weca+c
vHVX+zMMMLP8rPBUxRMbmmmMAXGe2oD45UqEkf9ypjEMpeGntDO9Jyd3Ws6DWeaMpk+FTsyBxslE
gwgjIt9COBc9UzGLZjPJ6dPauXZZv4L+rh2K2sBizA+mJEl/bmpRbV6nCHJrCU4rpTeo1JiOK5vv
lCpC/kWjaZaJS0cJizXLsLk8zmParihj/a88Rv/T1mneFJJxUQ8dcACE/E4WaVFJDoBKxGj5ZYQQ
13t7zsJUIY3B9zOu6dVCVO8uLLxcBXGvvIbhuOWsZRPy1c265ysYUU7X3R8My5E28Wz0PQ5D4GuH
UukEbPLqQ0pRNocMFVqwF/CruTESGf1DNKbk0USqKw1JVCOYPoH1kx6k5drf0ggEgNbkBbZZ6fnE
JDy4VhAIgyPmluCLj+rBMTATUTTmYYYjX2/w01d2pFr+91AnNZT1GqFZCN7DyeQ1HRn9ofG/Fq67
4cSkbrrbVCwpehTSpXWG0zsy7UxIp40OkKwi0u4s5sPffaHIjKfniCzPcXcoOirYPcu0mV3hflXX
OlKXTOrPzOW0g6BkAuDWaWKUfTSY6cEFz+nqtykJTehoAco3dVL0TQzCdwnBaVVL7Rg7qaGSIQLH
Qt9Fz5CUyOXpNohOFsrMBaw1mfnzxUNdBJcwv4DaWHwLsR+JkJVcT0MpD7reeujkYlfUWcKHpcQO
csUlx6zhqHDAS2K8xvj/XZ9/BWynoGpCaLOU8yKbrtbhtIyeeltH4+bSREZP/72FOCCbHnYoUiwy
SR7Q7O/1TirbLDUb4RzGjKFiUHCXcJ9eeK28ayvz+Dls7vUEMt1MbKMTMbT14AIsCA+s1bGCbRLy
DiPFnQUOHqprfh0h9ut5cRz9r+cR5xZmzdQ9FCsEiZgpZCHa8DZGtaJ5lQMu45/OjBRdzWN+4iBa
s4p1R67ntzb5aIPJv4nyIhfqNsEhAArarmg5BdMNjgF5BCzgFwxhy20I62i0UU86aZidGPgX+gxd
gj/BB7+RK+u9SqaLnm3mVeFnCfVaG/3MUt0sx0WS3nA8gxIRckwdeKf+V7zJoTYQ7JwuGM+MBk58
lKd41GLxlykXQ7gqPzCWROrGLB6O9/JEpPy4xsM4zQEikce4JZ9/VvkURV1+qcB3+McGQHzlzD+r
nDiygfQ/hZ64ll8sOIG58BsL4QWOAk2DYn0fjybIp7ZdQSwvGB6jTHEKaG6nBrmSOUlB9fPdQn/i
UJxrMox3etf7Mja1H9CVpgUr5u62PbfstAgr+vrGf4hieG4s9YV3nck8dzarvEurWsprGbuyjFWy
7YmEV3dvJOw0k9wuyW/Fl23Sg6o2QkP6oQfwLfGKOVtuL1oFX9e2yFFDzpPX7jd/phxxthW0TgiU
CGAqNxCDNlLtFZ5WoQdskfxqVa40P5DEE6fZXSgfO7nkhXqpVlnEtq5slPZOAwRYSMsNXd48XMfJ
nPUX7ck1vyHRN5PT/NlADf55uRYHuNnLI588OkuJb4r8ZkjpfL6WhlljbQ1wEcdIdAj1kLudfjtO
xNrgGsTYLU5je+sMtny/7l0tgpKtSCDdAkBAwGN5XeDukyGwoSbEVkgLo/ShC2Hp16sitE3hFKd6
WBn/Z4rrWF++PO+oSj0ihMlHdZsKzK/phDZ69j9vvFu/NaeaXJrqpD78ycrxo6JuLkASMqD3RmyA
jibu2ZMv0e4PWq6Z2UnQYzYO/YXJbYGvEy5b7CKKO/J++AeFQDPU2ZNZkWz62fqtUJz26uJtmrlP
uin3enP7SjEO582asITU6G8aoZzvqg8U8YZGeZLAYuwugfWvUF8B9HarYnYTHNHJW9iXIOqIoV+p
75EWccgpG5m0utiSWXID7gF9sgvh/jFT2Z/qGHMlOgipzin6dednk99fgIp7RSSduuGUghize60o
mMxB14HGV0YcQz4YwjuqplyeaQ61As41kMEUIUAOf/5+6csCjK/lzq9AsoRZVFSHaX2CAvt98b0b
VULSyHyywQKQuW7zXzsF3JlQpK1hPF2AIX8qUxxcbv+x3z+G2iOGp3z6fL18WM80Yi7I8vML6Ssf
cUpOwKb+92eN6u9izsYHPnStpOvD7tB4fvkQ2fVOvyZwUFodlymapzY3CojXqJeKBDUvP5qCLimM
RbiHTGjgogKK0yP2FR80s+18+wNlL4L/ULaCS3aGc47Dck3aOjoIa+Qgai+/SV+T/HfGEkIKk+tV
yUmNxcAQXtlD1wHsslFaMxpsvtpSPXZu7CxO5FB1c/LPR5Lxk1+soy19n6WdkOG6fb5yK3s+iuV/
DAl/HV1A0h4Gw7ZSh54yhXFoo8V3IfUWMNIgU6Jt6Js71p3KAROAm9/ys6IiUZKA0ivPdhU9YXiQ
PdfxfUGk59LmOV9D6lfVZzfwE9EyYfJduzFUyN+LVmPOImVEIjpp+mtCw5ud1IKhVzXtpHxiIsvQ
jUFKG/lF5rnayHSFZ8+Bx0/dCG6w3EpwS0vzbP1iFuXBzyAT35h2q21yfa5np7KV9oCiw7syfMmT
7qNkfkuzJYXt+c1saTOnoj+HtKzDm05mkViL4a6fXv590Eq3m3p0TdBJfzII0pn6vVOyAlqI4H0A
HfJ7uMcyCm77BfBcBzpMj+NoTGtqEzxpJjP2RDoLedUGS61fnYfvuqDS0F/ZGfd81FaqVLPASQGy
br8mcA88Tvk7riFXgbsuVmjdEGYkGWRzuI9kzCklYF6vID0T5K3WDFjpezTrhIin3vMsPHTRO0LW
jzyPfTyf4zGhSEFky2v8O9vgToLDSOY6mQnoQtWniNfTEo/bLIkbMwC3TRpTt2ZoF9rKjTsiWbOU
qpcBueKwdTXpA79bk9XR9F44HZdx07CtoVwr0+8sgxWv4gOm8XPf6Wb6V/eQmwqmQAEQTWyD14/P
QsLrt9MFp9vqs9S+d2SyONnBt9YjUk7LUzo+rcyH92qChK1ED407gcP1fxSlIK7icFdMN0e6Z/aL
l1+t9C9kGkbsxlMGFfQ9NyZGIiSse8MNYvE5wmjyrMEMPVMQrL8ga8SLkOIrpoEoa4GdErlE3mju
I8nm2FUgdlTbp/nmFwImV3X6CK4YlF6Y5a/fN4jrZ+0SMKF5cICevaVk7M+Llx8V1Wa63NpgY995
0q8xQ/OiDbr2iijR+nwpvF5zhwWaRvybGbyvNtzSLr0XPlB7RO7GJbyF6zoPv2KrZAan3MZQt+4Q
dMWihnMTIOCYPoztyvpOqHvBv1etVaqJp4DiGrUevHy8/H6SzkjPg+/CRql91V1fjMKklUS2FV3U
ZlAWEhL/95rLQ/rpZsqA76KTmOYEtPFLW0qOExCHZynvX36GE/0fA2EsVr8AF0kgDIO6ZzQsW/N5
/fDPygpwos6g39dSeU30w0GWs0JwlgL8C5eT/tu6a9PzvIUPyw8YSyh2n4byBpW+NX+y/R7uH+se
oH5lCrbQ2EDF7ZyBoFCsql4NzbI/1vDXR0HIcXavacCp5NHeKqGe+0uA7nFn9Gw3PaXEiE5/bR0P
nkvux6/U+Ss/Sfs6vuRbXKv4oJdNklYoMSQjS+FT5UVC9wokSU1vBYCdh77Ia6j8mUAi4ekSNpWY
SdP5A6p3bZkXc45NptNrex59yBLYzEf+i1SNiSIZNvF6XN4dL9HVf8saFrgRRB+dB/tgLtGYmkEL
fM9gcIV8RZpatNVjYHHSoKDOz8R+pir2YmQuY9M59d8z7xynOHmP1vxBXL5l+YTEd9PheiZGHHBO
qII2S9nG7J6Yar9A6AshDs6VRviEm4kuGlH8GLQN/YCx204c4cgVZExbIh4+Ij4jOC5zQTvYAES0
OUxHE+4WoI4Kr33I9icum7nd/uG+EispUHyHRZsU+4BxAFckZjJ9lHfPZbt4yv1+HBXeW3rQCKrc
Ng+bt5DVXNOV0WCVGSQmQG88nx1D/13L5e6f12ehMlHTm6Uzbovm107Bm93u37TsK5VdyNZbPEId
03w1jN4nkcj+tcB5GIxSoh8XED4IC+IymDqGSsWFOmPKmPLaS5UPpHsvV6ZpgI8BficYw9kxx+2c
NF6xVE4yZiX6xp9ZuETGTuF3V9v5TGAL2bIol78ATTGJmuWfjozEnrBPHV1dTk0Jj5QRrpMls32i
XBoYK8ucI8Gvsv+6Fww0qPQ+UbPXiQyj6mri5yRKVZ6ceyj45U2sfEU2h/kpCbaAEmweqZIy1/jT
NjM3eS936Di/WV/xDORN63TISbLaCoKLRROO97f5vEk4IHLG07da8xRUr6Ma06CpHt4VG+8gX4sc
i3UyRNSkXh0yBFe5BVAEmPbpvaarfU9T9apbhx6IhMKqgzWEJUwjPArafRKpMZyKsJuvvlvCjaZl
1lDSQgkfGkqm1pwrTEdwJTr0H9/omnOwn4ymexM/nBOpZZv+XS/jgpq1MIEvHYOgwZwsnBPjglA+
UwY88ZL8nXaazatwPN42AEQmnk2VOg9TKYo+qJ9V5mcoWZBJL4tsq+UOFo5JUHkZTLv0cCbZraKA
E/knvFccNKmUxsWRhx49XdDeZ6iZo6a+VgL0tMz+u8FGIJzNoXm5500/f98O1kv7DkGi4XgP4U3s
6CqhwwwFDQaYFJUWINn8/JaqWhiDoHE7E2ezefQ7QokWG/ZZEwfgxa4K9FMo2gTo3jXHAHEgZvIC
u8c1CojeVl+eHwRVHg6otVLu6BXGds0jm+zN+5fudxkxRpNI8lhSUkrrbTtvllHvNGi+KFg7yBoT
YNTlqlLdFrxYmkCddpLFkVYn284x0y3Di9AZweNncjT95lKlPUv6DKjR6L+XBMstCttEh0HFngqR
WCiqdI9N01Ioyz+0XIpHaZqx7k5L7hd/cR8oi1BYLimYrIWr8QaT93MJwKmGaqlElVT/sKcVlFhQ
zEvESsp5Ub4yqWXn+AQiW7WtZC2J5lXjbPShWk/FekME+VyH0xRWPLgpdW/A65MUwfc9fnCkwj29
5JjUagLPs8eNI2RZ/+6n6V1fwVQe1nR9c7czQfNUvkkXUWjqmjY1g9Y3Wh+rnAW+hKosBMPTAfrd
S8iD6dKEpekhEavHJESCKVoCDPCjYhSDw2eT1bcUwNRO5xlG40z3cIcb39PpXSun9xA6wxFnNmwa
iwq03wS04SWFf2vuPUfRPI8Z2UwovRMWjPfjaWflwwnl+GAM6MlfHbwyljDC5xvLJAQsXy9Dfc18
7Yr+wKtMlhQLodpN3JJ4or1Qsg3B6IhXCNGHFrCp56ApDaxb0r0lyqRULyne+I4kLXVF5kEExDB3
LaxqigRI/zmyFZd7zafGN+AjviubYU0udQKruiMqIGXOC91XRwUXYa9oynV8p8aaDHnsxrkJd1gi
jYdHI9a7Q3kFj3WGz8uYDJJbVrKb+MHjJ+sH440XBQHpul0z4WFJPaE6zz47gRlyOzCNS0uw+81H
OetpsTxZZN8ThEnd4v7wBY4Sv1KPbFoprUqQrLtZCczgHAfEfAfcMXWQs47tW0YNrbIPbir/a0O1
wNi7gQdn9mWkztjM5QkQvmvbUZ73VpyG8aI2Ya7mZa2N81Pfbv8qPg+VRSaJvYWk1hX7HPiDhUtH
YL0qvNEySdAZkuNVhGct9UKXTBo1RP5IPoC5XY/maYG4zta/X9NVicKhUDvgw6/B2zvVlDA1CG3Q
3HxEx8GXbTVduSlhReYiYCITrnRjyopL865vy3R37a3OBx7TW69cW1GDR2iE6QavT0ms6FaMReRv
eVJnxBNP+geLYaFyQ9An1QXNJ60xHVR+bFUxO0AayuayRQ4Kgm7n53pgqSVYFVFE9EB1DSrMfnFU
ZjCex1UcAid0HtD5m0kbdn6s54/RElJtwB+uuJr7GwZCLiRaXECn8DAkJr1uE+cJXgLSLiI7xQQ9
p+GIYm4GxacoSk7unO/z6WoOb0Loo5IoK8MuZme25Ev/cQ3zL94ffdrcdwkSI+ZFx0jNHtgJhxBQ
mGqL3QnbAtO99EzFtrtPsOlJua0JZ3esA1/etgL7uWXoqTY0Pwrmr2IJSjvR+eFSBCwUTpDAXplY
m25JcUzb5RdoLFQ4m53q2pUdnEdBoZAxoorOex478GVL/UHgWWzoxCz96XLZk5MUGb5BEWVwnEjz
7ChRvigCgKJbEqWErYmdxyZm/Y760ST0kFaKsjHf9Nm1BiQROaE47kuAmm3v9iqHhtv+Y8AXb3jP
E8TefLQ26yPTTqgjLqU3nuiePs1WKnhqQ8BRp3DYSGRXTMDM/GPvgE1Y/QDP/AzABq/J97t3G/qN
4Aa5/TwH/uH7TJgGx4o+cRNdyi/Vcyx0Sf9nDGyyK926Vv/aBcGag334kVNizYiHewKxxWS5qw+0
lQ/UUEUiBUhbAM8+ZZRyzuEXAJWvvj6IeUIBsFbdBCtbIMEkgTHUp51sq4+Vy6VaSWSAbKLT2EmS
xUrcLCdSy5DQCoMQRLDWdMaa0F2c8ZHbJVZPntTIMbseAbJX79APGR8YIqI9280d9wJKppn2tTQZ
+9js7BLiOc/nPnpQbJQfGzCJZDFQdmXGgofhaGriFmaXhNyjihF7Vd9/z3KLqHLga0yNpE7UaPtE
vHw/E8+1iZLa+7PjekVFrDVUjFgGTaRBL8oI25Z4u0a/rULOhdCOmj6Fg5gLmJJZt0Zed7aStX1O
+jDhgxfw0l01iQ9jJcTTL4gl3yjnh+Xq3IVaUiswDg63zcu+r1bbpo1AtgE+cHfg3mhaTAR4aQdd
OUZXE1QH2IJmAiwdyur/cPI6fqE2EfPODR2UurF7ts8n2HvQ5P4WnWgSResG5OHknc7V6YgCFdIO
E2dKz/rS6JJJhv0hi64MXiyKhYi4aRuiJ8Kn0PTzjRmBzpYDwcLMDqwFRtYd/hrP5eG1CRPreB0Y
UuDfjsYhsiEV2R0NIDmT8wgRb+2jD9QZYZe58PGi0E5tlr47xuXjAtObavesmscOM29G7Ds4l/+S
mNxBP3nCcBMXLA6jaAdh+UTWyW7ctY3zc2Icxu4aqT98GiL0zMYdGyUv2N6GWjoKhR+5QhrIJt40
NmbkIprzJG9Gx3/lM21DDc4IHvh/riyX/xMOr884MoWOsa9yCiBaOCeQOo33wGSR91QsEDnhSfL1
OCR3FqtWezo4zYtzlDO6vM8MzQlZybAIiLPb2v1dPiym4wAGXZaarfhxSu+LsDMZOFd4QKUsGWgD
9p6vSKkgU3AQyCT0dB4+u3nwyJauFpREAyYF06IO28PhLWjFsPvGzVke8CHe2yyP84UwtfRxT/Y8
8dDs4tDDuRguwhwsF53Edu5QpbPmVpEohOo+TXGvVDav6VKqNJnOTZKlyLpXYsv/JXkV7wsP3P7y
/FW6iFeleNHFQgIXabPThoYeoc9I3E+m16JDiQCVws2N0cDIaBjZXn95Xlg8HUD3wee6ABsX22v+
QEK14f3dqscRISTEODrYLzfyxGWI3lCxw/P7uQrzU89xbXVH5FtsQDqezxXXdvyQ6qHzr2uV2rEe
rvfpcnBspBqSICj0IFtay3/g3Df1I6JnQOY0woAUWJjoS+Qi0XDshKcJB6LERI6BgfmFAMMIHfJY
l8EMCBwt1xvxfF69KxzajXibY3viFbVlkugiEj6mn79/Y6WPDl1zF44hUlK57hOSoVPgfwNzR5ky
fsuECeEvpNlz7k1gR6OZfscGUawVEHKZuZA3Gua4Kod+bJvMAxilAL1yR2WCAAjZAOR6WRZ4XVLs
G+z+rghpJqd4KQLnni9KYKmyTTE9/TUDCXZUYoAj1IpfaS34l6qDUcd4q1cF57xt6WyFBK2OZG3A
Fgcj9bm58rxKxgfA/OmS+xLBZ6F/x4QEb8QWe3ZHQk0669m9/DvYfMRJXikZjlO8Ta0R6JNuHunn
Yj/xxi7o61kSn1Fz89MjSDyLxhemUlS0OGZ53hJ0ZgtlwOKjjZviDjsF5iBicg7Plx28Ue1ecLnY
RsEIEQ2XvfP3Ki58MmVQSjkoIeG1p6BavtAGigncPNkmEhpdy3QfV1uEJ0PObvt572Hvxp9/0y5B
gbNQAEczU/4nboLbneaKf0Gywy0MYqJXTSWjhVapl8Mw6uznaJB/oWtT0qSV7AtBGOHQ1J7pEacR
9xVZ8CPFAkPLbCRn8ibwgAaFrvtMvEyQkTgIOmYsZVT48O4c2MXe6KORO75vDkSirLYWPZ2r9fP3
EYzcW0Uo+Yvd+/UXGYFtY02hcWJ5+ScaZiBpAlSL8t29CLxXTYdcOPSgCflwasVVPWHUg5zx1ADq
HUy/st+jFhjlN+W0rtTXKTEgMCNsSTx3tpFKPJbPIPGluOoCEvb4+nL5K6mlT8dzlatmCK0Gvdtc
qej5MWmTMgGzGmOh2UzdbhSPMBiTFqKEBiW7MpLNUsyXX3e4ScsF0x4TEHyrg2O/wfr4zfbwjKou
jBPLfBuwG0Ao2CariyRe51Oiq2MEk/qAy5Z1Gw+T8BqpPF+dDUh8CDjJwVjRlvCGZ/Tp5+YDVpwv
elNe+epeoqZxriF6//ioEGTNi8CflGLG/KNUu9eW0s/K/4Ks2p06qKIbt3JCfa5bynkDCJNJ1Rs1
CNNZ1v6xo7DYxz4aBUXIf2znTo5PU9YbYNN8BsNIDiaxysDA+jfj5ZxP0ivaAaZHVpjt1hM2AjqH
2GWEOgmV50ZYZ40wjuhlSy6UJkuUPAPiDeB3Q5Wp+Xkd9tJa7flOz0xuu7MEcCEFjKyeMcPeEbNp
pLZ318/89e119qqEu66hXMPgj9P3oj/MeDg/B0RJ3zZBxlc+XtS+24gv7Esq5vVWpSRGQUyl7QA+
N3LGVqbjipitaCajqreWnUbUKrT1a7LpO5PY+2UJL3ElbNl3e7Be72AKehaqT8sGQ6wsSgqRmnvx
pXB6FrAkF+m9s4bIfjxc4AuV7xchuMii/kKS+AQm9mjdLVT5ytBevbL4v/duPWDZiB61qdLZN+Ai
l6j2So2akxA4SedNvjGY02QVdSKV2Uz/sTCBTZMPf4EI/QYQTnL8AJHPEjnhAd4kAG4EZFsUJ8Kn
3gLgS0iWs2Ps2RV8RwgXi06qRPkPVvuWuAmxvQBZReR20vlmNDwC3pRla1+pCW9sQAP99VEZREwv
uYPUy5YAicbO4osHLklGZhMMtaRkAnYEUmSUMgOPPcAFfI/l91RaB0WAi70bsOypFWwJye5oNFjG
dnW1+WHBNT3QnYD+USMtAdH7FbjbTol3Z+7/9AE4IH6qMzhJW7g9LVG27pOkV1Q/jRJoMui5W9Jd
vH2e80Roi1zd4JOZAA3fteJv5SVn5WcqVBGf0gOYzwikajH6J7raCHl7FbFxGVFOvOrRzhNCe+ma
8Pkpv/w6u0ov/d+TyU1qBxVP+63DpqvXkePe2WL+w+6SvGldvVhWrq1DuuYhNDMWUmE5gtjyHy0e
tshkrq+SbWQzFH7jO1IRXonQZSBXnxU/EsNs92d3klnH9xVdqovcu4bVminBn7wkgtzFAb3gFB9K
7ZaKT8bKgobppz9lVStlaJHmMwATNKMC/86ZWAicgpk0FOUSNohagj8JwLFdwq4r90snsjUs9htL
aNmK6w8lIUM9u840nE30bwfO5XaxL1Ubc1UyixMStCaW5taBIiD5UTwCfTLkm9OA5oCYmiQ/ziPx
6vJNhX43z6Cut0KIG163zOlx8GfCU12k9Q+WGdF88o4zKhjbR+9D/eesXZMOdVy5UCprssQb2EcQ
ySHrOojQTwmh6Fut4oHUtrgWo/I2uLRCpQbxBoE4NGA5tahq4D779SeVtFjnmc9uwx7muhCRh5df
DNB5Hbvl4BKtUJX1NSerX27C/mqEWzUHrrs2/vv2oNGJKxxvB6K5NQ0v9XqUY/6anjuBnLppIZ5z
/kPXyQSv6TkprZxOoLinDtwM8vXvfZaNVvQaB0sKGRkkmZy5kapwgMBvvt2idTS0vsnYfW88w6Fc
EWoQDRCBDMwJb3VXlNk97+o31BdNLiT8hx7uxlsZ59+BW7BsS0qugd9Vo8QC9yTz+FmsVsmkCIhH
DoCaowMv6bqebuvsca3kQwO90qRSq+GfplebZdRbLtIaGbq+xYOBrbkuBFKgAlWytzZKiBYN5O0j
let9XiOcKzzvAasdd8x//Zxkk6ZQYyVWT5GuV+IrCrv/DsiTPgByaThuril00PRP+RNDrLFuyBcA
9nLrzKLWUT55cuOiWYyavj2TczKYYcX0fbU67UqltDukB3870LMsyfiYS3PASqhNzA/TGaDAOGE0
waG5j9itkaYgFvyews7NWXQqGTlF6g6XUso8qhfF4ghzGypq6HeATnRyRahKX9YiQK2lgFlVhnZI
vc3+rW/0ptEuyomQTLse+eyJs44F58vKhmacCgXRIWNm+4kGhKgSgoT+AYm47ojf96q2Hcbt2Eiq
cdqZlJiCTjoka966GQ36YESkX8yiPYDfibeVeKg67sHgv/uj3Rb9Sx6CO1n0L64mAUkQJm1wnvHB
9E0zojcP4YvegB/Y5n/KpADk1fmCA+JtlOiXAEYqDBQITTdFLMVtFfiQHHauf8T1YxBu4+QG4gpL
P0B3mCQ9eJ4yfOb6afu9Y7/AMzdHQXabjrxWqmrARQSfUZOeC0d94hdIDDgB9g3QNTCI/3r5P8hR
wXP3Nzk9kEFouzTrWy8i6PoMtvMSPhUsmKe0hQkwrGaD0yE/hwnctkJNjNPFsycM1omsx2KuD2ot
g7zr9zpq0oLu4zK2NMe6nAlorGxyNeYubzQ6MJt7YOs0OOLSdy72B35eZYLo2MHi6DBtZPnvUDMV
QEnhjBy+QL7IssTCksF9uN5KkeDaAOQDmtddMNWHxHq8YaIX/iHBxjM8/0RAcKY7GDG5lOFvqlZs
nK0txos54AqvM3KyllbqKiO5iQB9sAderPjTNLS3MALOtErJy3CJTH2S22XyPnECAKMi9dxzMTBp
GjtC8sv7NtgDoyN15QX4Ti64ey9IkkMA2Hw1LErN3xAcUaMbnyu4J98t8jk3L3kjf/yi4pkNFC95
s51lEiOsX4K2shkxhTwEA/u8Z59x9x5N2v1eYfSyR1p7ztXCwudC6aZLjeaSkXZDAqoXPuBLZu6+
JBqQ+OcNc+vC2WFMGjJVmwTnUxE9Y29tzqXuApTNjXDcZe9PKwHCAYSphycKS1ju57bcZtEt5Hcg
5BtlDn+VxUQRiIATuSE11cPc2Vdk6FUGeIXIz5NSeUiiJAiBZeAiZSQN2HBhBlv3BrrZwmyAAI5+
721CroaeQFqMixAhd7hFh4EipQorXCwyWvj4yTltqzc53LnUjMhq8xxI5uAwifNi1f61Tq5rI1Nx
iJsi1uG0lQBPoWC/PnMN78FgDaotSfkrWl81lWz6QNwMDfTUkc1/mSJqTCLE7WKJydpIRymCGxY9
u11ho7uKMnvab56853MvFnZKctqUzMIvSy24hCc6UAMe1iZCi9wfSVDmCT/aMDXp5S3MhMc68a3T
Z94ZyP/KCwQiSVQN+X2xHnQwAcM43ro84LMOGB8ZHuGpjp0mJOaDq8O/agB9q4bNFvimbilcIwmT
ImNoabXmPxlZoTeCp8oyJk4OuxbF3X4C09BrXqWDX33UYiTiCp/rptnygn3dnf8sXPo448JPw41Y
uDp2xzbJ8Q6sP3STtkueZhpeIlOJy9o0sWTtEyTDvVmldaQQZl8GY2bF6iQrVspsB+KzQbO1Mk5s
JkMbZF7R5QAlgXLmGIw6+nIg+ClyMSE1IKF97tI+YKOQTTtV7lhuBa/4M0zJ56noEtwk2pvVVJsU
F49ysiNPjvcv2GU3npq9TloGudLILcta0ZmZCVfUcoq+bueXMt4L8XJObCk/qjJcTXDH39lDPiSz
QRWsLvcK08lWxj1HWWOtTpeQN04NKvlxwyT0xQkgDu6W3aPW2VWCqZAqMVPjf7m6567oZAdar0Hb
7Q79jeoMXM17+h8kOiLlpSY0I6MEdqjiNfcs4Q7/C0epxmrby5u5XOrUEsyu+ilUfAleZXMCHiKi
5Y0qI6gsz7i477c6ax4oKHCd8v6mPwfIlUneH5naolwBn4u3dCWdgG/f0unR2pOWnhF/tULHo49z
8yPZnSRg/htMW1LT/oY3w58Fi277+bayK9dtVRd1N3kCRTjd9zTSusUzRHyMcvzElpNoKRqsW1cG
0qnagRIgDBZio8jgyf/dKBH3cCF72yueZ08Am4UfqCcmdHbnD3//Qz/tAcoAElHbnBbmG74HLgtK
pOhyPx2hBL9JvfLDokf2fE6jPB9bsI0I0ei6wITYsTHrazkfrfYuU+qcrsmiKmdVOE4LyHkH5ubd
/CQ1GQ3RHRshtvx+x4SMw4pMWRnV5gtrrlTgPOYnXLukm4HwB9DRjmx7AVCb5xFyJjfDSXAAEc7Z
FBup7AX2rAMm6sEzvCwKmJ2fU2GRPH8CHAWTOzAaCdABQ36A2f/sJaW+N6u9qOLATZaRCmombGUG
4GNk3wMAfzU6BoqPxMg6noj3rIJxHsM41KcecEE4FtOufKhKqE1WQ0gJDRUkY9PVyNpnPxWO613N
SA/B7/hPmwSqn4FkBgcsVd+5L7irPOLsFI2RseR6kycWaDSJx0JHqdJztf9VOv4N1mrhtz7YkV6h
c9QfkZQvRZiJhO6A07p5FGtFjD0Ilg7x2dhQbJJHz9LDGjLREfmVfuqLzutCgDIivv8KD9+QSPgv
n31UUb8ICbwyxkVncPcDGGbon2yv0QuzJE1rbzCEExr1ypOur9AmoFlNFby9IvuWcCXSSPHawnNs
VlsD/V47yKwXBU6vMsuatTu3Owy7KjVUgnCGbTH0Ma55PQ2qM4Zl1+oX+4c55JNO4SvDun9Bubed
S9PCB1GRZwi/MWNTYq+WaUCj9pC976qyyrG6CnEuW5o5m7xXjHMf33Z5p82SBqPxRkVD23doi/JM
g70cnKYDhrsDu/PV/UDm/UB+sK+Vh75+QVT05IGsIoMQTmkFu5xij0tStZ7TcSDUhxPYvnO60rQB
EpWrdMm8aCN2aErxoMO88DEGnivFF2votiCJ6HH/Pg/iu0IlgMmDomRruoxhGuMtZjGE4CSpkGij
xSNUDfefeV+PmFXadJ69vEtf94va97eClZcUzUwDjQaWNnKeSCWIcRNeyQUkzBUA0oPFMdAN1GE7
mLH9DAfdprtd8Xo6KiaHhKZg8TAIBvGvulqztLVQ8/7+4rx1Ohg/6S6PMKKnf55qd58pLMYXfuJM
zE0jqKd7aMS+EdIY+fh5ZEHQUgtrhcSKuciu9YpA1R2WB9Dgzz9fyOjsp1rVCOxYERt0nixJbyha
0fvS1SFxuW4oWagTf/Ywow/yJYc73Y1Rt07l5h3aUkdiZJReFArLm2lznmmr2Pk0h8McQTf73Q7g
95A2PddmPfu2OArX7+onUH1OyW9OxiidN6LSgu7Y8s2ybRjUjZ4ahX/OhPz3tdYqdvoombDjGznL
5rPQpHm9/ZoXc1ZvN8vX5C+GCAhJKzWZJutyZZRYZ7TftjC/dpeXhbotcPpFDHLVEBT4MyaI85kq
9gAeaE4Y3llPJxTblKk676aPUnMaRhV//9gyz/Hz+aXBAmNyRNfDmyvDEbeMViaQq/+BEnSxFuuV
D4ohhbGUQY/slOtYwJaAigAWkXyaXRbcZlIpNKGmNLFOMFfcbueuRmvb5jUgvjFaCqfBLs5rhad2
1XBJ1OmLP7AauIQXyoQm13lE0Gt6UA3w3EsV49m7LuNTkmUqnj1y1L64VVkkfndpcM1LPGpHQhIA
3DC9HKSkk5mWABEOtXcZt0MLevwh8dihvtxKM1K0FboJPy3N7pOfc4+B5MOIjdWWAP3QV/DHaAoL
xa9mY4P6FYpIWjJ0uSrk0YWVLJ4SScyC4qQuvPj5+ykZGACpTfu6ShFMUGrbdv1ffldnD2fVd1ep
pVrYIjHaMx3F0mymc4tckJMhn+Wpaex2IabFrRWv9kRXvkrpDPNBp+jcvKN2njbc/qJxnOw7EE8Z
j17bqZvdn/ckJd0fR2wV5f2FYfFYZKF2bs95dXGVmYgYXNTWQswOi600k5qxKw2y3ZLGLC9LBL3v
j8CxOtzUl6EpkYiPg8TGQmQdRt1VZ8EBv25CIS7q91WiCTw9WZjaaIC4uS6dXbVjJ6LEiU+IHTJk
j03c//0MWiEHmovBkYs2DFRZXlnwUw45VpxD/ZXSHq4qRKV1Lxr0x4MRSIiBS0LPniAWQ/Z/l0fp
JTwhUfpBTKX1R3u6riHbHyUxcVmns+tTEingtlQLnkXYqZIcujI2GlC6E6r2+DFu3IJV8g5okUWF
nXVeD5NHMpxHj/e7In2KCZOuHz+12+UTz0p6M1Xt7sNIsMgITFvX/TF50lbO4qGsXRbIA9t2rl3H
lNW4Gva6AMwnA8UyVai3KYhH5KIBbgaiv8YsRilERpR46b5pjJ9iOlryPDIayt8OhgbTaqcMwaDj
pvqeQEGQNW8xB/GUQPRyUr4MzwdiPzlCbZ9cX6tx5Ro1gGXH/Oz7/8+aAbDJhTFoRs2MhConcHWE
uAFIGEGHF3X6+OmsrBWaCYUNAIWLYW8PlENT5SY3ALztqzP+9zv5x9M/Jl/WAMJp2vZ5V1FQF+pr
ZYJARWuNYknvmi2GR0bN2Y+/RkscfJeK5uRi7cqOO0CcrQiL+GSE5W/6IwzhNiKuVVdXB+QpBB6R
9f/9FaX6Ghptj6yPBvcxg2rJO4BVAIByIXEuC9NYzVlxhv2QkSxDY/oYF7KkozE7qtx7rASTBSwg
nFJzSbu5a2MqyZ4tRljlHoyQ2Mc8r6QPBEr6ovozWy9WqyfYKG6lln7z5LH3rLX5Odmem8tFMG78
f9hXSDi1H9H6UzNzfeMxt3M4y9uExURyK2wJnJ/CP0etB/UXP3DEPKvYu44D1Fu/d9te5v8et/C2
gfwTrocinQo0TxtZF93mkPAfVir+hLzhZ0JXKqmFPzjWD9mtFPte5AyubMM6JZ6uI+FKEQQndvWk
lXgJBpKufR/oHudbSeRPTC/2a8zOxk+HriQqo8qmn/9fRqcn/nckiHd+fBvQiEAArasuYvt1t3BD
7kYiUaSoKDuwQptT9f0pAPYgdLHF4ULURNFAQ92eZBQ5B2oaARCFySFdYEWmDVPA+ZA8Rn7a2RV7
IdZZRJTLl2tB0ZfoapU2dD3/5QbHnz6hf9K8VB/UyoIRYKaSlP6hqSXIIuD1Sy/A/Zq/iLSmZGP3
+h5FDIeAlPQSGM115AkFdLt5ECY/04/eKg7pwhahOIbv5YH+Yf1cp9Ek+AU4AZgFUqnDu8LjwO2n
4yXGgaz1c/l96N2RqLqDqNNp6de4JBhAMAFPgq0q9h1tiY4lYOmuPUOCAcnx6AC46kQN8w+g5Npl
RoVSbvvk7cxubaT31Fx3j/A84XKt/VrHN1js1U9ecxmeR/XPalpeposW//Lq/iKrSkrz9yeHazxZ
aVfkWe//P2CuKYGA7DLbdQ3ZSACTpJ5JV3aIHB9s1WwV8UirE7xb+y/F4pEm1Q7DBUTzCtuRpErW
hSAg/lBZ4WunJafSYJq4hPvfAHhy3HO+TPj+jm48ouUAMrEZg9kHqsvnJjaHPfMpYRRIL+l74wVj
yCV2jQMWT6ge0DWT0hps99uKnz8mSU45T2UcpiDbAo2OKJFSZgc3x+ouqZvglSI4S1BsXuWrKLUO
Ewh3FBufFHeOdz6EAov0cfFovgYDLcLzWureD2ghtAGBpffo07j9wc/T2/u6+Ix4zQuc9EuPIyqo
9Dcz8IPGf44wWKfUmd8igajBTwRmiPOMq+aIUcpl9voSRPXH9avizuAg9u4q8M4fzUbMdKasd4We
QiFcOw6zFBNKRPlcb4qVt3EnWgDME3Epymw8jiKyx/2BHURG4S8/3yhCzneGs848hmA8A3y9xe3g
qI7JiTFQHrV1OBnXtT1HyMHU3sVTRV6PTOWM1rpUQ+KArkwpSxgQvHXTBY1WVPppl3FzqLM5tH3f
/DTqfoR3z+/fF+bIoyHNCr6Ds96CSnfwo7GRsSFqI5koVO2grc2o+5I40xbDhL1bZ1Ce7bpp0U0d
K0DFwKfNf2ca1GcygpD0aTbhUV6NxUOKiEQtYjBqw/GlHNC0/Rz42AjR0/7K8aFCO0yKa5KFLtrD
JG2EkSJ6Vnqf1JcMiiEOaObIPSAoVhnALc2hQm/8CTUxu5Z+RttI6VLXJugimml5R38ZimbW1taP
2u549QE1LgZ19cvLSNxqolEd9XyT8LfyqCRWBOlQdqvHBmi4eLOS9X2wN9Nqe82jCt6NAHT3+Ei8
akqjb0aLJSM7wmI0NWEgogIl61ttWU4xR/pJEUmVxzjQ/xCUrd8jkwfLaSvulnsvVOfYkA15VKAN
jvDK5t+cUFvTmqfZYrqSt0lb3GfT7daCXgu1BQAmVQeYb8oJRWwVhIwj3ICJ4RQg1FqEJrd9hDNL
GRME+u0xQ3aa4ndMqgcPvFEfQVFD+5SuXvtDJ4EhhbB8dPZTu4V9m4f0PTx/uFqDzUWcXdlVow7u
1tTP6ExJ7CEKS1/63li0++qm2tjB7D1348YV7qDQOv6nL0Mrpehf0Mge53H4fNW1icZekGc/PGZM
Q3P+dpx6O/cH6Ehq7h84ZsK+Vvmh0N/2GgLCqpaTy4sSFcK4pMLKgNDJJBppZdI/VGMKwTxiJUjL
/fb02DlERAXqWLMn6PXnsiPRZJasdmquzg0EmRS/w9QGc9i74WGjmHplctAVv/AizJ3yJWXtYLRK
Lyvxhw91b9h6N7IUajFj+39x63Ml3XtiZoYuX7WUljvkX0rO4McgAqLC4t89fbzfJ3ZVQ4pNX9we
4GubHTvQ3JryvpIJKMvHV2pB8fdjMTCwvVG4I3A9XFutJeOJ2kjbaKDL1WFxdi9xRdP4QUQmQegR
oVOQ2qm1iBMpXNRrd8l4WNSQEU0ZPcekg4uFOUFoapXB5kZn2kSxEHH1O+m6+YKdiZICP1Lx9On5
DypHtL++FlAM+erHDTmN/2oa98+0ALWrjgtbvGEyRAcSIpRYqmjGIXjzfGq6Z3DKAb79D9gyyoz7
DIMUcOGIFUfKOvPgx4h8SuSOhsPQQiJAztDl3GOGlrAJkERvbELdbcV0iXuRo7YrWRnep/j+zy89
I/hILAN0rxR0JnmD/Y0gU7xLZThWSlyHMAb6eOQTojUpp88sthdUqbw3A+AK2yt/exK9S/0roDd4
iO7WEUdayd/StNo1oT1k3CCEBgwJihvPK6ZpL5Qd7WxEc0Xjs6LwaLlUSF9Dp4wSWGWZb0m9BgR8
pZWtuQdvlg6iGche5txJ78hSANvBSDDPNk/jivq6okYkNi9oFYSPb3S29sA/tu4xmkiAy6VIgRz/
9+Qi3NBRg3780LEoRrjZQlrn1syb9Jtg3qHZex8IL2S8HTmhhv1U2tZJVGeDdsuIwKpMOiAIC7yy
BdbyBbmdx8T/aZ+Co7Zzr6RSUUwwhh0DqHfr3S4UUh+WdZu7SkiAEP1Ht/BgRVxde0u6h3jLGMKS
jYI0ETwWcAsW/aQb/IO2fGzXFASHCBw4D1+Yosut68hT9vLpiQr6ezzCnCFvVeh3/+Hjbwlif+fC
qy8mz6Q5mV3q/Acet0LQbCnb29CX5d/Tx+Xhljrvcf2v8CC+363jIv08GytHXV8eqZ/08aPDcQAe
SvMYjUb5G7GsSSpFrpXEqkdVhejPF9p2WlknM9ciiOJe/668digAF2nM//8/2LhGJfuNaipjL6BI
o54lUBG+1cmKFxrrfOZX+j1U3UQhaTXuVkWG6BLN2jH2f6HtJnj3c5W/tPX0/nzFXf++Q7B/oro5
sOKEzHIz2BqJCVLipMa8SRG1u6zpR787mb/ZV1M6JCJZz2vOIAGgUFho59lyQXwQboY1gFXwpzVn
/GSmQgBzQDm6ad4hII3KbND2WLMAXH6rVzLE9ZxyYoRRArEiF1BHAmCAjmggLa4IMcoT/K1evvnM
obbprlmpjJyIPHjlGUfEP/dkqPzAHPWEKl6g3pcgxdmMtvUIEDtfB/sR9B1xZFNrti7EeaE4c9na
O3AlVltcFt5eVzvcgavBoyZHZyhgxU2PoB5SU935/HFRzYV+KXTCeRODhMPAKPjtkUXJeIM8YlgG
U+EyCFVM/DxcX3deAY3WNy/uSLhJeFL5GmmBEvqLcOJg3m16AnSVowJC8d/JAjwwkpM+m1Plba79
MAfgcCOHQx8FMC5Jg3k/L9+Aqm6eqDjQD365a8L/jTswIzcpQDvIw02/NKnX9CGA+TzbbU6Lm+CN
4BbyvuK0Z7cGovUKm6fw1V+/MfPif8koJHJnQaB/+1dnXz3HIPs/UWAqCVa+gmpcn6q98nvDhknK
4fsHgK4LrCBjt/c+7s89TomYDeABnxRogVTqKXeIRGG4OlRhdm6lQFa2mkayRoHPVYn8mlMjZpxF
QfNIgA2Flmt2iChP4tZO5YCiKm+zJe3C1elkncSPVHCPwYm8QywhnITmKOZEfnfoBAKX0tiM/wHB
P6al464Z+ymTAPbWbsjtmKu/8hsy0h9h2/VP8AOL6tm9YKj/JYf35AhQrqY0qv59kThbMMZoPb2u
5NPImCEjZNBQiIcHvDDpwt/NCo6D+RPmicDTm89ZlrFhGC9Utnjo2/dFq5gE/7HoxO6iIy2X9KEq
VUrOT7se6AvSkxhRlsEG8N8T0Hp21/1fpXDzdj/XlDOHJjjTMgqkQ5LykcHEVKtE7SqV6CphOsnG
z/XfShDi40uw7zOizaOmDv3s6jca6FhsratWEHuxKFRvKzQvpCLd5KRfYUSXOc9uMPno5WqJbgfc
Ca7R/EwlNo6GPEElCrlT+rNTJCQEtmhdh5IRanlFGhgo3fuYayJOdo//tnesdlvfe880wnM1H6y1
xJ9wm4MT4m9MZTONgGYwgxKx4SPiHtzxFgA3uq45o1g2GHmKr/10gKImY+cw+397K4h1aZeTSbZL
0qdT22TzjVPhgsugvQy3Hdv5UXZnKDFQiHIPXyYf7ZRC9Pblsmkup1OZCJYwIY2eSqeyjIwVzlZM
DI9JpE7r3DY0JbRCgdRjDPwBjjgnbUkCL8XyYMYCseGV8aCy/Ry2BanXNyB5yq5XmsvX/Wp4yWMY
HXrKl1lugtuLRoB3+DBng7wPqUyMCdJkOO+hW+M8rczUolNON6LVARVYomXz3hg1g50XnJwAj22m
PlL6ctWpeL1ZjiZj5Nzjq9ts9e1WUU4RJUO5BZTg/Beu3y0FQtHmGhdVlH3QI9G4DQ3MEWrPKvW8
Ifxjyoy5CwRLbutsBJO+Hsk4ARqbfz34cwBv7m4B64ZboQourbmmRH9Kc/X4nzGUY9qpFBmwcH7m
gLAX/D4eQZkQJCwCVIUTr3RVmHwzOs2ujxO1Tc/bX6MFsal/yNgVe/AD1aWinNx727PJkfGmw2Jz
iM1Nv/+6r3KJdMTbCBZqRtLekSohUMP9uvOHmwQrkHPHBJVRDZ6qzT7vhxVlPY6Hn7W+ZnPlyE5G
WIMI4di1/mSBad8HUvI5eb4D49PKCtcvTNGNZO9ubAg4eOepE9gzJ+MJ/w67arh+HbE1Jukwgd/L
rUQ1DA8m0A5vyptb7I5jvfLKeagKs8ZJdnJwbdKL6IK3jY/2dNJYSx1EcWrjHaPkuFjhuuSbo8Al
BZmVxxgXSRJwHuIA80AiH8zRcVhSohyqazy+fsy+8SNOe/5WAqXXL+oAhD3/4WrXg0M4g6yiq2vW
ixgKiZg/trG66XbhHT1ks5SkMte1wpkBkMQiG273+v/2TOdp8tnqqaOCA/OXeqiTEfvFCCvJAlZW
cEDwieaqDupBU0XP5xELo1OQPBATSQxmY12hyLiPN20TizrBqxgdHFuehubB83tqtmKljtZeoo1K
HPygLUwExynTVbwUVWdWw0G4NFxvOlz+84FH+A9Owuja34QJPqkWG3ycvv51H45eul1JYwHhXsaP
vgcODsbEXWAkNFs5DmIzvXkGHXoH8quhjUMCkgAxy2E2HIMTr9tPhpED3ALOOcNkIsWYdymZ10gZ
z6mWawRiUTbt4KkIxJ/8/Q5HZDQcZGhvFcpZO2GsIzGMHGaEmQpWpCtvngPleJT6I+iWtbKctkok
C1EWGSo1r0cnrc7JMwzA3gWQVN2ekXuRajKJfsw/7cjT1H1w4EHlZjD0V69/F+qkXejjy1TfhlPn
YITpQ1FUQ8mu1nGiSujqlcYxXu/+xRiI3FObWAdsGBj46RrZ+EakcrQz/irIOQDanOCJ68RvICJ+
paLByckfM3KQgxHhai5j5DvMlz5QXZogkCNUT0vddnGWWx+B3qnvLpjMp1LV0h/Y0NHRv7tW4fsi
7TElRBwZeFyhKThc2TE1NCrSDXevJeE7BLUT4faBqOYaFpcCaHjuBJ2kAOgS4xlD3RNCAFLcT9Vf
Bftl8pfQUaLszyDE0qQtY8O96ljOmy9+9Oc2S62Pps/ilmPAsTVINrISlXAD+1Df1T5c/e54y0B0
Jc1wHXyvXhQNF+UgMtzH+YeBFqrypcDudbRRTK59S/FT5RmtZAEkPVU6EPJAXdRr8Ty1YA/H7MXB
W4pJM5xlmovZNBJzElINNYEsIONnp062XysFrz8EwtV/l77Ycx3yem0WdEdJnDVefTCQ5OFDU1MA
hx/GQUKlCv2ruepcVKN1k0XW4ms+yT/RT7aHagf/MBgXdlh1TWddtNzBbSbzTeK1K76VJ0pKGXfx
FAzmkHDdi9+c2aQCqBxVivTc1JlWQozYdnOnJ+nhd6THxsfJ1Uj+1i8UI+Mco4MmowhDTBhiYoI5
BQN4kOwNjkOLiWa9jF6HTynGvpB9mFwFcGHGwrzKIkwuWmd86n/v3hsRckpDtKTHn7uEV88fqDX6
B2IY9nnOszSXwX4QSXUvDh4PrlDDgFS05S20wdtJxsJLTm3B6b5YF4ZEbdzdeEcCi4RDh2EHfFQD
1E9gLc3NvC++PRAgZmdz7oO3dRxmMZIxxT6eOaABf/Nk2P2wukymCV5Yn0vYT1TUYDlroYd42y12
Z8JD6nAFcZdavDtXgQWv/EPMtzrDkKLbRUcnDwdasLPMpaLBAEb28VvEv4l+QPur71mClSmztYD0
A+HphrTZnBQ87JRxb+LqpsUUUsL8uj9HfVqfXxvuenigLNuPd8HUlbgwGQwlfijGbWYz+LxwslHi
03dyQgsxyIvW5TEGRkaU6YW/MLn85rZQFFtOs94ew86+w6CGRo4GLa3vIqLyURlYj1JCAQw9qie9
F+e9DrQXKL7fdoI8+x1k+O+QwJqDzm46340EsQVmtiz1HhQ6Bl07DCIzaD6/kVezaUSC2Zxz5U4D
aElpBff3zBYjqYDsl1858LqrsU+FH7k+PZkixuLqNCeWsfyHvZaPl83020oOHZL6h/8sMJgvI73K
jB6oOlwsRgKsqva7no6C6NDz5Fr2yMge2Ky9cSBgF7c4HN8qnbbYJ1gTxC8NAQdQ2ntbamQuuwlh
hnPmdIBcBudXmr15vhpptnTl3zShW/N/S2VIJVn/X5e0Rno0Nw8BntWxHQnnKZ/4MUYdCsdG2oz9
ZzUS8ZCic8D8FCZdupb8hsW1VCaKzhH6q50UgtH/L+ksAn5MDLKYyiT64PGRtX0QvAb+oxffTH5g
eoW27m64XHOjf1/liFRd29fco6XRwSSje1rWjtONPtHpnO95f9t9hyXJAquro7wEEUB0xU/9+uCE
vHmhwP9hKPTyvwDbzMFse5zV5823lyxg2eiaY+EJCI7auZooajH4APxPa9Po5V7C/WR54Jc9auSi
gqkdvLpb674BFoDUb8RAHJLTFPMyFbYKe601/B6HOmWM+wZpxyfyTdQnjowxIFRKLKPfY185cFIc
cFsc71q365PF3z7r7z5ARx3Pn0XjVXFY6mCNjcECokov2swWbWX8esEPLU3duVCZqfPTA3qXiKGJ
wKSuNxYj7KOOXRLHPTVCUGNdryoob6AXrDZqP0QPZnEgAk6gaj/90am2QsfPONX6PTI9iLodDwM7
pLixS3G1V5T0qCHpPaP9h15+8SVKfeSrQ2rv6fWfzQv5NfoerzYd19O/a67srJrlIOWYuYMs6GgN
4TzFmqjb3yJWU/yMutlnWDl55Xxryt+Ot5N4447Yx8FxcWuyVPeI91nM3k/CPcDFUtWMLVgoUGUb
gpb7KlKsxeCLnWFfjLpnadPz+ChZGnt/gczHXwkV+poGykZ7Ms5lUUK/eIMs9X3ZQD1Yba0H1QW1
MHG+SpgmTcVPBj967uKn/MJUpsYQBi27OtzRJ5VYL6JwlIhJ7hhp2MMR9h7ZfulUNZP49Y9Jo6qD
L23ldWFVWisfKlgVV5wXByg5vReFVEP+RgGFKzC0LE9Qcgyl1KhjkrBsAD1QGex/I90Bq4PgNF7J
0u2uly1qwwBsaVBur/XzSzsN2562icQ1Pe+FNu/etZg16xYvpjWr7TqiW6D3NiZUcEzHHDvLNzAl
0odjovsd2NB35zUWvj70JiTLqTN4MvViNGPItceGxjyuZ0tOx9aCGGoEj/3yHRejUkGtVglpHTCV
qbrJUqCM2vhh8IC81Jmw+yKo8kzPAkl0xA7zDuzu356KhF6y+h5V3E1ZXLXxbiV7f0JJ7GXIzMq4
qGOtl/SPa0X88akKAZ8dCROImMRc8VYJlSvDmGHeQSt4VBedObIL2Kry4EJN9IDZ4x9BDoOJgO5q
XTrCps2MvGd193GoKRP09aX+wKXt9XXs7rnmGXi+A3VEe3tMBX2jG5okLXzNa7JCxvEaH3SlW/hI
prFLKzqA757w3isY38TRjzZeb6dg9Ge6In9RjnpYBW4/GS+5aezGwyV+6V9po4BmQfQ9wikCpjVP
chIYs/gnCtfV0bFznJsXz47uLtU25U/cbZiLyvrjTyfqLZLQtYuyxBHK3wLsSzndzkE1nQlaOSSf
b9bDQnJ3u8gGT7wqSE6kedTlYJJN+uxXtU53X+KOD+ZaU7lS94nvMaHkmIgF34ka6PFpGufg1gDp
1MWmdUGiuK0VkXYCopbejVyT9LdARwX1pUY2hmmgTkJ2sUEWGzKBuW7vkb8M3oGir+l6p9HFviPK
0X2Csc6LRO+cxoy4fjPNiuKsf/hpgRMScPWkWJIZaY8hE5P7h5J0NAeOUI+qXa0lJU1fUY3QJSD0
D5kVRyx44WaJ4unoBm3Uv4icNvjF6MCasNNslL2g//p+kGN1isuQ9JYe+8slouekpOt+1eRNTIWc
t1y1D/dgt6tFow4VJ8Qn7VprDtpRotAbgV8WVR+v1JVNMeyh8aHalGSpM06t9Wdeu3HO58sqVTrV
o7XQtKG0Cy2jUTKKLpvXBohuJnm94nX9gcVeaazm/eYgqNMMdA06DJbjD2miVF8Yuh2GYZMVQSlc
vnBi5e6nrhwoeVG8B1o3r2m1TJudEKLKATKlg3APB234667SaVVcEE2m0myMaAuFpPqVH/dPKiEg
95JAT14hepnTpDier0konCRgpw+zZnkvssupthON8JjyVE0Zb0RaLX+m50wceXEGk+cgvqvs5zhL
HnJyqeEBq1ZzPsJOYc+hrDbuTBPjM5fN5fNr8IavSoyYXgGr5l0Tkz170o7BRn/NRQCGEkHFAa0n
D7bXf5g5Cl+vEzY2CK5RopPftWxGUpSfw9nGaDjxsNZAC1S3dRnsnXha5+xdVOPd7/C0KHcxw1v+
u816HLcOvXZ6uRCTBhIVO43ZddW1KY8vxKS7LRf5zQ7zX55iy2WdVfFbqsfSZKBnhmi0lxSxPxiW
qRSvXYCDjaYxMX510v2ZHJ2rEqos0jtuTUJ4s9J5I7xBsS/1FCCAVMeS9wgNWgSiGQCYmFtlm20M
i9Ob7VwoCan7Vql6KWrLMufqsUUABtBPtXSbQXPS7kUZbi1XWk0sIfPHe0JMAq3Fb+YpugQKEvnQ
Tifstz+PTYgaV1PdwLhQGATasSrNJdKl0irj3ITB2I4yGs+JeiTxGntIlpPrraRh9SN97zXY916r
IHqRUWB9YCi7OtbjFJfWf2bxtVP3WpPZ5WvThZt13ZxcTjTR+5181HE4/Pu64kN/LT5HHxkGQikJ
lDy6PLrD0R0OUg2CxfzaXM6jxomSl6ap3fqXUpF6hrmCC54WEQDE4zDgcw4956AFFdlzeXgIv2B7
5GpWtInv+YMXAGu5ufIXuhdnqliESAJFqEwUEMV4WifBDJ9WVN3/M8VZCdeS3sjC6uuWzl02Yu1T
/qY4NzioBMOZtA1josck97loV/fQ7KDTJYD0s4lF/kSDwm9y/Y9PNs194ak9WrK9KyDrRWJcYz4D
y+ez1OoLtw8DCvjcxX11V2JWm3joDGZmdz+4+7guSvGsvPe6P0XEWHlnkgAz/jYa582MoD6WN/9u
CbIa5Q+dRyyARLSqiF4xusuni4Cldz0TsegOwEbjSngjwPzQQ9cSGG9VXPsyhGnq9yrpgAS+7EfU
Nwu5r8fBAMu44isV5SSEOEPdzGYa4anFaRCL+XCXOAnXuTuVQMXEi7Tn9xhA/65JWfdcmqw/FOPf
CxR9VF+u/JtsR/Z4sm4fC6Wqd1dW7TT7GS72itqo9rTMwh4zwzowlEpacTMstEpsa5C0PVwPN1gm
7e/NUcYe7vGBO/yuvVOMrvAiKCJSY7yiFl4sV9CjU6awEal5bPamRUXvxzwvU3XRFXtormstmYoA
0HZxFXxdcQ5V1Kv0NiGNvSgYJBDAGSOzRun4mnXZMr4jGbljEN1J50LiYvR9MP5mFx3R4+Skvo0I
Lh4tiQJDUuRCqsXmxhsc2K95kNCyiGRPE0RaH2zKzf8zJulSGA+YMHvJ9ENhtVTMFK3zfUZHkimm
k9ibBf5t/db/7AuGjN1o96P64ToxPfJHp4BWBvNJwYANdp6cYAsVd/pvfDTtv02UpGI/pVuTGeh0
YhVexlFFutXK0qL6E+vPEOMO56lvOhvjXOgtp8ImLkDe0xqVAVDW/KrOP3uYOUV7xazyayq8fA/I
+xcr01pwQ4SVL8UW+6ozfqEZGrCds936XvXKFZAGbIiA9WI1SMIT7aCVTg8L9DeWLpK2ShOoTjeP
NfrGfbZsybAOwwuKs/0phj4QXx/3tXKY37e4rZZPOr5QIdXxqcjPfn0h31am8ct2JesCqmyrlSh1
LslvryWgPPKqGuPBp5S0L2oT7+OW6Ve605GGQkXJZohpFEDhza0Dct173mGwCwoMUQVg5+EtVBnQ
XVVeIo4SRTFfOxa52+DiRZqIxXs4JxfBwzADYyUYNFLM6uhDM/azqWNVZyQ2R4cOnWZt3/RUof2t
njeyoQ3AZBnpEAyjmXyeRv7K1BRMKJG1YZxbjzSZGGYjQimVyQnrFnQ5kGvBhBSyrBz18zmoaKqP
Jp66gcq53kJlHrG0KpKvySVs71xlGglR+cK6b7r2/WDNaa889l5KBzfzfbxecOyZxdMJoOUSPEzE
n4emNowckJyaEKFjhrydgHOzh1Th/pErZbYeM0DyWk/vN7o2e8dbaVpTlz/09G34O96rkwzSykbb
FcqjiuVo+Wi92w182heCNHNB9TrXTmuvg8KSWd5qKEQ/b8aXSWbNK+7guOksPOjY9SOMtUO5EDbQ
Spzh5icOpmFDT6jkDLRP4xlErYxik/n17cE7K6Q6qIBH/KSgQtEYX3D/gk7BywsKl6abj72XDL5Z
kzZq4lGPx+2CT0TEotpOOkW8iCnec/7MLmOE4H4q8JaAJA6SNR2idClBjvQKonugsOoqrmOqLdKD
9g3JOZuhX54tP3IUV5T+I8JbHn2LSKwpERTH+IPuEBKfvFDE/aqSZnHJuuo6Vl54IjQ0KfgN1NdO
smXHkfRMXhr+vy827vKNZWT7zp/vMUy7SMo2NhkAazieSLTIxl8eB2+aiXdELkgDOI12WfU0w0+8
kBAJ614d88Iyr+9CbogSfwLwy2nyCkna042aLfoFAhbpElTpAzsdnq+Eow3Y9X1MJoWuzevbAxh+
9uMFcpVono6d8W/knbELiCW3X673wSeLNJPlAUucIs2fRUITiJ9zt+dK1bp1dbaM5s5PPNU1gCcC
fwQSVlH2/umvQorZyFtKYl/iA+237XHQvU237CM6tuS1FYfqYcRAhIAMIjbG1oBpok3YFjpGBlsw
76CqwVvQBJrhpEZrKQqdlx0wt+qNXMUZqMngZc9mMpWIOlO9K1wS4dXEK5QeSJeOKPwanF1ydQuu
jeVoa+urriAKF3v9w5ChjsTRS0GCOgpNO3l24m9HB4+1Gk5cecuejkrFqcVF6oYJFwdD2YPZUzLK
PoMh2C3H4sBNMknoYrrWa/EVaG5vUhR0r6D14D995kkhTwjFXF3dm8hSk0m9Kb73Jo8CbMuTAz+f
L6u+GPK3K8xriv6MUcBfDzsUeGN1AC9ZeahWli85OIImGgRFoIEWmt3smWRECFv8rSOIHlbpuSOu
UYDOC6xNfogYMRpk4SjV58NwTjoK8uajPMLOy/ksW0hiGrCm87YsX5rGzYOBpNCH3KweBgjDfmjY
PiWkTiu6//mACMvqtMZIce9BrmZqrsI33xTBYJ7DoWogpWkaFwbmNjN0aJpTlQRopGHRMES3j0W+
GnsrzgKRr2twVgHYPFyf+tLPAzWdk+geTtRGzjJH+w2/YejJWg2yfV9SwSX4ZpFDe4OGXOQWqnh2
mh91D18heS6uEP/RgilEqALVJ7mCvhKvzb0QhSP6zfSmW72hk4vhgIIHSYrUX0OyOkfK5o1fcvWp
IKFj4cge8mpiaqimb8UV/LXK9EzZkg8mKKDb+0MCnsSEYgufQWtgAckuGYtytiAOuTZg6xv7QXBv
oBCl6M5dg4Nn0gVqUoCh94oC38Vcy6F9bUK4rusYnPT0lFW/+geKdzSCU0r9eqnGd/Kgw6TkPITU
/NS5J+dEF6mquws1ESryu1SdLQL5HShF+aJGqHcuXddV223vTfxpckQ+6NaaXBGX6+DV5dH0dU72
/bigghe4Gpiig5BaRq+8pnt7mzj9NtsXNLerFoAM18A0w8tU701WzFOqlpI/R/Y2kveTDEWvVtwB
BBqBmF3A/g9kH4FvlPcBsm07jzzl7+1PsjOqCvvHeJ0WXKj08YJZ1+iEptudsAygJtqzKqiCzaGR
3ZZHC6LK6/l2/HHXhPZdVt0DbGOKsdjBeIqinygz+tKu8SVCLSrEiU7ewktcwK8P+Nff4VWl6GeR
0d8SxoWp1tEpUbwuOQMQWdBCpgQtCsU6b2P2BEp6h9KcFxWWIwhqlaIRZxCRxXdoEL2nLm3149rh
wtzU0IP3c4E4YyNXIQcjc/EyxS7HwwJfEOAuU7UgmSuzS481tUy2/DgtPIX/cVTEWhyi3eHAdeNq
Rn7BbfHNalO7RPPdK9Y8+L8Eeui0WkE7zEoFVBCu/MtBeRqDuV7XJhCDfduiEjNf1jjgwlQVHj9p
SMohFlDIdb3cneN0kRA7IDneM8zVlIGb/STkblJnS3KpP+XvCvhFXKNMlx8AJzlyjwWm1lMMZuCz
zp2PIM8gpRm2d1a8zOlNRtos0+rnYTTiZXKup9GVpIc9EIgYjPartUK8NPPj1S8wQFT68ypRYD2f
fQitnymI9/QzWjJdres2PQsbxBZsAuD3HIplNO7J7sshxORWTD9iWGIbObDL87FowhJ5dc6achIa
GSjaUbg7J9mmc/x6gR1+IPQ7HyZMhebINqVVSaSXDm56iT25D8izSi01s8jQd+CzzOBZnv9JHoMW
wVaqk+x9JMD9/ifoV1aiWJw90rXM20fbg1Pa/ARwDPmi9GJkZjta5SQhDIdCj0qlDCt/5/NgqaWq
Mic/yrhV9AkeBRTRGNU8p8iteeJU3Y6t8Ph0VzcImYglPBr5fkpSLUh9Vy7/HxIYlpr41DmxrXoN
LVwy8k1/jOhjaosubjjoIFJ/L8TsL8A6VGSUW1JcBqggJs8b84rdti0a8O9SEehxZG755LGnXfgc
kWRkSXPqQY26QCTrBoMxiqzGNyO7JKX7gBIU0CnqzeiDLYeH56Y6dylXMdCSJH51nQjxV+QsOprV
sVhLmGvJEqHao4OfO50vhf4ARTTi/iHQ3jfzGYyOfMgpWVWBC2594P/0N4pADyeInSAt/sdx3NOs
2eghNMqy18Pb1uUXuRsK6PoFpnTl0uRcLa2sntV1HAQjJUxGrQP84hb7xVO8myR3QGuqSBKIZobi
N6rs2W5ZMIq+jezE8g5H5D0P8qamEsF6IUTL+QbiFtvWac4KSf6xl+w5uAGnPP2F6Nd4sjIb/M19
fZlGNeRXHCSJAqSq/xG2aNP+q59vaH7Xby0kq2To3AC4wS9M+nlkM0/wuMxOVekCNjKeHxyoOvog
m8PwCYa9J2OxyMo/GFBX0LphoXJEFT/ypiWdWLrtHn+yhNzKsgqwKUNChsB5nJrNZsM60xPmLrZX
kACcRG2ca73MMpjO1ZZt2MigGLunGPkCbsytLtQnnULGO5HYooyONI3pf+nZqX531FQhZcy04qsE
tNP+putcIYtMrQdYvKjMBMfLiUJxeWW8ziroo74Yc37ePX9E4wM9OTBnCZ/BYXp++631Ufrm9jPz
9vExjkyNPLgJ6gel+fhnl8za2O3wY++AI31j7dcWrKacbRPAKEua2yqhbwWmCgKYzTLZoaSQ97ql
nBXCStKfDEp3dlyrZjPUj2LD24t3mHaHJG8fnmvahb7pTKMfK0BjOejtoKzNylodyx2UhttXrNVP
HonATDkBs82KXGVNsXW8HHDxnToZS3GGWMIfYeDjHrbMgFAmbbmco3B8qRBfmV9te8rqTLf5rLJe
fv1oBjlvFXD7CVznMosAIwBNzkYpcik/GkTXQl9CpURn3IQ+tNetKDsMnq69F3ckUkOgBBhK6SFv
qL4LP0xPlYa1amqOJ735Z2Ve5wQPZoGIwfFnNvU+3v4MNS4xs8S40/LL1/vU204oLj+GE02jA8Uu
zHukDWr92Jm3UimeGX9tITvVOZtocXC9Rs4lrfH1GKlUsXNdvGI10HIVqpJx/sxSQEk9xuyAqiGw
nywnx+loGeeRm/kk3DmKj9+WKRwmFRvlph258RHHCutrOwpuKfltb2NuqDgQykB+EMU+rJUST8sA
WCKAit2NAlP317So9mvTWG6bS/1Qg0XbePRgCuU1wKk3PAmbcVtovr48GTwHlJOetmsbV92lL/o7
3UP6yVvy4diIrrpZD3lVjrFBq3bqvlXagvs6dv0Vvmz8n+1U9BkX78Pr9xVBVrVoEgYvmenarpFy
1kz2WGNddRba9HeBBBxApktc4sUnf0cIMM3IxA1u1dyY7/1is/AaA1Nr4039RCYMpssTlaYsjX4V
QTTIWyqcIN+NVRpUJkVRXGfvKwnCcRxjtjWWkYr2VD/IuCGNCUvr32C1LOCWpwMXdc9lK5soyTas
EJoZpLRDJVKTKwVSfw+7OCHj+wgVIbCdwK2HNCubuLKOIscHeosDaGD8rSN8j/BhLIS4X8/czEVr
rMjEoK6n2Zy/fZBy94MRm4ChWPV57QOBGNVvXQ0g8mknJYXnsuftv8zILU+lAAYhINva7yuBAraZ
icryy1IV8z74vxmII5SnBbCTKzzqy5rMb1JMYX7NJgXOweTOpzziqqIk6cJUEr7S7oqzbBKeTtg+
/BOCZEA29bHUhVjmJ4sKtKek0C5WYubTQ+Ycr+Ri9la99ZmJJHPIF7oNlEVsmFxSMdVCJJD9Ax2G
eZAcHDrXRWzekrQQUx8eakknEgRpz2xkcyKFaT+itktyW2QOd0KtV0ITe1ID9zBK9LrroqNeLiAJ
5hVZxlUUYfEJ7OHJc3j6tkHfK7BnIdGA4hfIcB1hzBYXwbV2kOBYNGNOfV2WLZn1hYTYZ1oYwruw
OD4fKgfjq2O4GNRqglmaJWAkHdffwGmsQx5Nbilg5CjC1EOjBzxr5SpJsyt0/2wNr5V2/0Jh9EyE
+lcs+ITVZZh3CpobDyxlqD09VK54rzt3sftgUQz5Bd7OI90w1XwrPDrL2zGk6yVZJZ/7TRyS8+TX
UjNxYPTQk9cmOKO/GhJZqEoM02Up0lUGqE5OXZcPjYh0BQM5Q2MobTvW6T2TDjjSokjp2cM0MB+h
RPeY2iAqpxT7Ec7SBRfpqqsl85py3vtqqNILdc0jDYKIEvFGEKs3zA8DXeBA30PzYJo5z/Nt2f9k
3KqYRrUlGmnpV/7K8JKAwWN8GjP5zG1N1IrqwDwAO8S7Z/9JzQCGa5ZIaHg0W/SFAheaRrYa2UEz
+2bGjOEjNUdS76w2+8xwNdFI/Ly3ctvHBlYW2JarBMkkje4Wx+n5hx+pC038KRXIqGrkwV9GktvS
H3CDcCxKzGrOwHdRzXfZ2gNc7UKE7NJyFndUAWHDouGkqqtRaebPcHaAIbjpwEDkOLuTRSMpSb1o
iqjTuWP9SCfQBPF60JqV+Ory+dQHlzvONuWKYpt0pojy3rtKm1WzFgjJmVOlw89Nr/MskktmQqhz
YLfNlIUm19a+qU8n55pn4u67S/VHqX+sprRKJpX0dPFOW+03w2w3Ao/ATr9l2KQoLdh3JwBBeaxH
Ga0MkonU/sBJrgnD5U0nT0ay5J9bSYRX7Zhh+svCzZuSOgVeJNF3sI+qQYQwPBFWEIEWcyJ7qZ+i
jou0QAgI0KcOML+HuVtIkaUcz0cyJ1on04kRDB1KKrh/hHcHqri0g0SabMUPUBHNpi1Jdxp3lEVH
xh4dQ4fuph/Bc6Ch9zSIdAYUKCMyOaRdBFsDldBjh9UOZF8nCHPFn6XlwXsinaSZ/EwGHih6f9SH
a4lGKBAJa2LD9hX5nZguqng0rt/smbX6M7rL4DwleuE5V+HvZh9aTUtsY+t3bdxCdCkpMC/DGCxO
ZluIvBo5A96hyxWSgDOZJcEaoIiGqlL8WXnh8K1hOtoc4ApXTDN01FHL+VHRUfVR+KUCfb9T3gqP
ncFTUKU08Ft+bWVhmMxyqlbDtYGfymRiKFpdpviTR+HVnj9aBccCNOo1sHejPUS5LQ9G1VutXSPy
BgHrzP8k4gtaLBFY8sDzj6YlTZhLodV1DtN9DRAKZPMtFGMxVBOhhiByOvDrRLgWEVoCZqh2rLYS
yPNf/ZDv2bOXBgqm3808LofTtmdxUWYFoW1orccHpk7G+3mli56oTDNOygxRui5HnBzbzuRTq+fQ
DVYdltzCxu8PMKBXfyDkjQEnOu27I30DL0oWuEWXLoL2Ipf6BKDrcdIXjraUHsDw35A+gz5Di8ag
qEZJAiW1DfSbivJ7dShfueVhpyT6EWqKW8w+5Xd90lzZBmIlIzp5MIgnJ4VO1hr3iAZkkVsPdAjS
UjAgJfYn3h1MMZyYJQtjIPUITLWBh0xiQNpBos7QdH1beLj5h/uAZfVyAUdXZnj815uK8+hFAEgU
K1YTEMJa/3eeJjjkJFgwBguqweP9jBgVrgFpXKC7+i9ebdfV4w/YZ4BNxMXhTPwho5Y4yLwJj5ZN
CcA4Z2cgivLS4AKRSBPVuntPRSzu0mvlafQVQ2S1ZYwU4sNlQMwJPKSrvISz8jnS6aUDJIjMY8Oh
pC4uy7ZkypZJ4EsHhxaviPMuqD/kZOtaLQHz8UUQ48qHt5wtWgpZipD78dopTPjrSPdCUtNeqpKD
hQo+qCu7cpRnfXFhLBsBwOg/zqHsNQ96uiS6NB2A/jxRINKuUJIPhv/Lgze2Etq9fY9dWrwihcdu
O4W2vkAW9nNTe2g2+afSNX4uamExLaBxYxW3PO8ro/CkMZs+YEkpo1ysM7Vaz7JNk6/1XU8E81l5
s7wmimJxEkChFgCGkV8QjBegKJN+h6YY/yUy3U5WpUmg8d8ij8JAMY3mK/Myt1L2qfGTiTEu+FS/
XR13AgrxgZ8cVJI5/3XflhZI3d1Sf9CTSKQX/UaMpOQ3Bp3QyC0ChwGoQuKREU/E41IwoKdfmRdx
dpTQWQhOom3DxNyCAYt7CRQgXgVkxTLk9G6ex+bzpxyujrm9YlMinEGhwur89KW5OjKqxUTAIVvn
PK37R1L6qQZjB/g3bsDq88ngml4uWhKKd9uOHUoNl338wWtCX7cf7Ky7jKUhfY2FMWiOrd0T/WLE
CMOru9/09IeGoof07GOejFxoL1ryKJUjlaeBld4ud+UbJ89TtS1xYrkIwFJ3bMZt7iwcE3iPm5HS
cBdPeMq6mtvV1EXU6hkWsV7Cpm+dWcC4pDBx7KrxnhvZIchMb7swUqWn3jaCUxIXRJpO4GrRocFb
7liXz0EkAavDW5H1u5fnrd0ul0953V0UgeimlUx0biezJQOqdg6GGmLhPMShe9izfjfap6AaYDgH
C57B7bFOo0VnjDSD6+eUZVY88eMYJyZyTsb4zuhvxYw4mKelxXGhUusumq6CTnimXXYfgcuJYVNG
GnHLvKkktnKz9jZTaN09Xlm9ICP7BxxeV7gNbSiZMFQ/vokxR79OzIlwUQL98whp0zEPNGKmVqNi
0c87f3JBvhd1Rp2DP7iFtlBivQI6CK1UvT9iM6iQMQ+LKKb5fygioG5tM51UeL8wxyPN1+ZlOsmQ
/xyocRGewAU2gQb0kubRc51YSQCB9DtmU/sKGMVnrz50JFjTl3lrH3dMHtFpOO4K3wZK35QJpYg8
w3ko115OT3TdEZcFdLHi3wTNxAy+d6xKw85P8IY5MiSRibogXuXs+RVu/K1qpPxA516xrcBImiIp
yBCoEpVRd8LBU0rWYDXcIV4ZMUMxEzZv8dSBNhA3L3Py8TIoaSEy8y5E6eZAsaNzGCslJNAKXz6T
sRXXURvIE8sOHKbW6M16Qny9P1TVvf/X9/30bT4r9b2R1mi+kvLaYvB198xvADOn1kStWsugHYSc
zfJYTTmbrqePkrREyNpua+/+h7Bu4pZi7aWt76HT4OunQCUxU0aQE0FQGxN41/GpCKpFcnziNwaz
PYEIsbsyf/DHDbO5shZ1C5Hx+BlzAsnmBuqAy35pvh3IdbBg0N/2wdMGNrvHVvafIu/J6Np6FyRL
JfDCUpL0iVv4wpNiNmInp6z6eqktff+7Li5JW6XHNdf+Z4hHSSl3RGiq7dqXYxKNO3sA8E21sESL
2plaYj6pq/GUacmZZD6i4TPzhUgpjBa+V7T+e3OuXHGHKh2Fi4XO7rFIKuuggw/Ty6zxWAfcsDjV
lgYLlDMAIFCuemByRNPCdRfHnmtzqXX3zj8BOScFxyN1Y8Cob56M3Ccki8Ko66uuFBa+/2geuWZm
khv/+bJzvjLJCzNMW8EzCS/TuzmSmk9fWSPKyzwzTlt2NoOoeb3KfTROrDV84uFkWQ8vRO5vbNe+
ck675bWa+VZ/dVMjgAqijYp9sKXb4PpFIiabA7bqH4GWf6/p4rhRXtrqdrt0mCQXSn3h7hGWuHij
ANmcshZZdKrJmEGwnbjD4pE+0lVX8B61ZzFvuUo13nQdCndM77CL180gCrjwJsWlFCMPum86hXB9
Lrz5uD9ghxFsX92whH6bdMbTxRjZV602sG2vhPV73fhipZEPKQHGDOWyZgDkn/urhpJYzuvGqiiE
9xwjiKqxUNnGsO7zZ7u1oh2LV88W9B/kpI7kWs06D4sRszx3ENV7vruirhkSd0phgvlFr2Ivzqfg
/B8twvJj0ty8oM4oP4QclDDri5UDlik9LouF89a04K1tFvXhO2ID2Jhq8jbX2/YWNsI8jR1jVAfG
u3emmKgwa6psj6dPagII5QVslYyQQ5lJb+gmZFZW60hRLrXJQOBmM5wlfFGARQmcdyoetXhxvUls
gyRkPw/TR5iNauHPVo1uE5VGs8pIwAkhlD8CjY7/ANNppBVafP0qIzhHviaLU4cQyAx/u+AAC6Lm
acD3AaqtS3VrqLFQ8LYYmp8alw/Y/MkYZpwXenT5wb9Wsp0TTGoE9NXUC1LdNe6asKF2sm/eseg2
kG/VpbP3b3yvQddvC1Ans7/NzCiywSUkabkJAQAea7c3b5hE5t7d3KJaxhmAzRCh0/YBEq5fbmUD
AY+Gu/ICLPg3IjpAgTBg0YKoYqXKpKWukKIt4Og1XxD/6HZ0KI5iphsemSJ6wd8rgbuvZLqAQsRy
ssY0q3WUDcPuAFNBwDCzNKOYGqWGB4JQFdSpT3p5XNWC9ZeXP12XiYHXHaEghC79lPCHB7EAa7k8
LcG2AZVvsBF8Z8bDfPFmuuKKQQ5rzuG63uD8bmt7fI2c5nUuWsit7+blrhNh6h7jAnIy8VMRyMmu
ZPLz+aIEmWlQSz0Lfbih7zNjd4elKX+yrgD+TrHxGR24q6nlIdaLJQCoN74EtwysZCASQ9UTJyJ0
EzjTEC6bEK4v4hIf4I+Pc8JQAkDV8R6aTZ/gVbfUjAscAY+uxUUZTf3ldNLvb5/WeL5X3+J7ODhh
iftVeIWynCaGFZm9HRIlBAqzDKvEy2uy5G+yMB+BpOIktnSTEeaIJSgVZOAHizRTWOAYU1qDmP28
JKdyb+JSpgtrno1ImDUhndpfZVkRJl2wIpVz4peod9UjYyzlSWUTbBRgBusr+0XiV+AtAP1GdQbn
W+4DbtpWS9L5xDdBfIcloIekMewISnN1spZFx492rh/iCSzQqbcj2ZI8tTGQN9fkU8lab/bJAiEH
kwYVRVdJrCYzIiMRTERCsczTIuaplkobe0lTxSjy2QSJYCJVJKG9ycoDFhKU4MD0kFLJ2EEi8Q4T
A7Kye3RNJqCU+uODMEXn36ilU+t+t8nTnkT+u0DV6l14LMAW6nAYyTF1wFcHBSy6AdYVkkk4JXIe
5gg8rujX8XXt5GN2ASmK9NvqO0QIOeksEOJ41XBCRRBDAEJHg0aCDoIjdqNV7gvwIbAN+XhApnTS
Zd2BlKynDaOBslG122XSk9pQCxltCrJt75zJhrxQSaugZKc4bhsOqY8/+p47LLMDwoEuIlUOiSB+
d7chJVcji4iVU3pFd5zY24vUL+KE1l8YCwlC3B4BOzvGM63lo07Jpvqj/jjk+k6MKYfAZiFTdKJB
lMnAZB2PvFPmPnP46fbSp7ChpMyVN6gabk4BTtgXduCrNER6hDYzo5l1Vz6tuuyEG2vAaUe8KDQ6
Nvd1JPVFPgIgltaeS5GMfnyoF1T2rieoErg/D+JYVLgQVF94WGf7eEy10qtZNhLxbHwgRe2bx1un
TeNpvyrbE/oLBwp89wmz/ZN+jHX30puTL8zjAkGsMzn6IXJtQw7yhP2MzQvp5ctE7y9hhORfWGaU
OuW6ADxgnC+IvBwzqjrgouMVDDoU2lIgCnnfusCdJeK/HX7CRp4VcrLOPTrYbHK2NlH8xmYfv0Qs
zT8jndBd8300o4DFjmX9j+bhEvRiUkeidrgyISwYyjspqGeFtf0puV8kTkSEX212VpyTrDYF3uMo
ZiFCGYMMQrUP/AuB8TE87eFyWDkuY4qY3nYlmPRSPzQG/7anMthm4fEz2MVr6WmG9c/6AEWno/KC
bjuM1xWZkjeqg3U2jDeYRYkAaJhUKBkppCRRGObXXOJ33SG+ypMxdgzX7q2GuBY0y26Gr95tvEid
yXHJnHIMerXRyI7eITnc2QE1Rx4zcPxrAwqkyfiyT547rNL8ib1YC+LuGnkFz/8H6TXnydtAvXg4
bnxuxj3f5sjjgcWWcwAK7F55Gw6kZ2jjmuUl5Hq4mtyCj5a88Etji0TP1SgfZ8nSrjbQHUjUb99q
eIJ+AE7tbzV+23chfRBGcpTlLiyU4p4LZw4w5jJ++1Hr0F5mp0q1rodmxgxr17jcTNb8EaWBzSjT
fLIveY80RP5LmM4/MNZFtAWuUje7CP2nFNOtQdD7vH9oPhTePgClKXKFvVUHFTaEEKu6oCdqj8H7
/NfLbEhSwvVUY/Xr3lFlXirCMTNPVvaiC/HXAFj+d48+X7DwkeSlzZgyolCH53rSf/8QwW7b6ka5
YsN3JzNRnU/3pKCSC8xgb/tJ1uDp9zinVrpSiz3JZJm5dYYGsrcdNu63DH5T86CVxJfH2v/EHCLO
8xSWZl6KwX6G72s8r5O3SlEdXfKMB1Jsj4MuD1vCUOZ9E5X4MfDiJ/rzesM55R3tQkpAh/FZTTv4
V9pbFIwdVjWpjImsRTPxbQHHft+OCLV6PDN0PNbPhb/VKWqOVmBp9/iIZ92PvCcQDk+xGAYe6deS
aM40D59rQnYWLb7W9ltBe8WotKk0ZFw4scjkuztQSappjLLXdVXaTQp2A8XA9hHfNEkmlN2WzxZl
7sS7MnirRRuEyrixz7yOi61NJrI0Olmn+5mBVuG5zwSg04zEl5P7+9f08PhhzTHvRxrE3J0CDjn7
VirKrtP2QpAGqzNkuSmLHKXK+g1bUhlnrN4T8LOPhZKnYUdV4oCVrTtwlRwXhMmafOneO4g9nzLn
F/zP0u5V79n9hlQKIN0cEXlys5OXnjymqPbzfPO6rGi9I/29rujRlhQZw5deOKOKv9EqyDgZPvlY
0hiox+TtuAE19A/bdZcc3ek35vo34rzD4WpYiNw2jt7aBjSPGGwNHOKwxAyDuxyR5yfo6UvUqfip
CoT3u/0xzhoqcz6YmVjVJoxCXe3J7VYRqffZZruLy2036QAc4bDw/lgblR93ShiMZX7L47FxoavI
MTWJhLwaM1RyjiKYO3ciwy42gHA87dNSereEY23jlm/sBYpOdYlcaGFKCpnJ4jTIRpCBY1Zi4/4v
lJufbfpwflLQcPFoyZKnmIZ+gbPTVomQg0PJTG8CVaMY/RHODpyBAGsdUL7wkOKpDrPvKzN98oCn
4+PE7liLkxuVa0uMmlpUqyFKhvHtcaaglSYnxG49DeGgAVG1CBd0zbJ/w1nvJIe4b6Rvu3V+G89f
WWlg4DEsva6RpdksJ5yzdtfNDZm5304gDtse1ILZrnLno2jgBeKZgOuSWKjOCSHeEdE4W/2bxfWI
xi40es2hPWFyeI+c5JYKQjYFI6rvPo1a5kuxrpkisUViKv7Cxc1nEg75pW1sIZ5hAOiE6sxn1Zzp
gr0DKSc5ReF/b6f7dF1bj1kdW7RBUYSUjrBBpuJrQE8vz6ASDOejHFjr86Zg8+oIV/QB2VY74JFd
hsgu8lZI7MELn0fm8z2/klDq9WCdnCRM6W/9pwE2YNu7BnspaD6q1zXSJqrhL3XKPzMmtkUNlTjs
QWDy6xLIlDzBlYwUR+pKT4uQPz2zapNN5nsemg6LLX8Qr7Clo+3iCwodsfw0g8jviJKEunslDj2q
SO3LK/hp075wQJ+FY3GRj9Ec55WncWRrHYxUtIBBJq5EB7suSvv34KNWHRV/c8GW2mtErsNhpOn8
ITsZxD5f/8eEcQXHvHMvVs/Uc0uVDoB/CnmLcatB3zF1plCbUfphfsD3TAnWLLt67m0U+q8ztu8e
+J40B+AtMjEBXaBwvKYi0/oVTWvmFlo7q0MCVpEIoMXfsnpM4nadLu9imHzHsvwoiuqmmezrCPvM
/L0vSSOCPIMd3jRrmzqiwHiZhq3NIUcWq4UXnV8lDy8QiLwa3/nO9QAouVbPKJuJW5xfGyOXoSCd
ZorMQYxdkwn2p6xIMwmsNUQNkyueaNeNsIMgt0FUC8h0ClvxlXUt2p5wwZ8p2O0g9gXFUYH2eAbZ
GUE7Wt1FzzzT6l0QX8Vdp9iux5Wwq2zN1AoVKajgZTFvgnb0+XJAZNRZJsHlx75GKhW41Wm91O2i
esG3WqHnr2pN3xzIRCI0MnuTwuFXnVLlanNx1qELfElHr0TAzWyYHYkzOLHzxmcACLwS146pHLj8
Q5eoid3sYPF15lUaxwWcs0EHfvmMN16sJf14czCNceprzPb3M8dDnNhMu09Y+Yi4Ymuw3kz75zo/
RPCV93GVgf5+ieweXEX9N2PcO4eVT9+ucfKM/cY2an8jUGmPDssdn08pkLYC8V0/Y6LDo8OUvZm2
YNKmQgiZliaaK25ZTR4HHz6McoWR+smoy0xz5pM2os+MchH0eQBlvaE8epSqVKK4hDxE31/4eDxF
XljcWsiMcf86+zcGD9zO4EmVo9Il6pRXngbixxFZ3J17SajkTrmWzGfYNdThpfSNHpvHlklq/usI
pvKU3HCFE9Ml6mrE768f8L9ZFSaK16mcNigQ4BOrmY+LmnUcCpeuNtsjFgeGVbvnhVHltM7/eiyB
BIg734BsAahKGddS+cDKWsdut9ihbLfYVr0C/4Q/IlwilqzbTA7eKF7lE0UL9+6Cf2tPDgnik4hF
K9sJg0oIZpTlMAgpbU/PrRQZcVUgyTVCj71Sts4lLqi3D//gRr7NE6FYnaNJGByW2pAL/7IIXVOK
CjxebyCjV7qf4wiQtedjO/amTZaAlCSBgHRiBtYugZJIonrN1Ypdh1QUHAXMSQOjSV5k9uHm4Rdm
JIil7BPiYPsIjimkfiAhXYE+WTQOiH0he6HdttTpvnYmsgYdIv7nzc7JxcFXHbzzH/Q5gpo7+XC2
bIWEeZfEucnvCp8wAJlLVcOnvLZ7WP4L9gZdV6YUpfY9Mxu525y1OWB0+yjeu/jcfGY+8Q9TV4mX
wH4fEMuHjzmUhStq/YVQxtwYrCdU07mfJ+kJZyfQmfa2sOdtv+nV7mvmOPjYKggcnePbicSxwkJk
UbAKRiwvBYwtt0acmZHYl7vy5PNZERuNRaf+sAKOX8Z6vAYmU/lP92a6sxIUGu67tRxeqeJmwUOn
zUv+qiQygGiinft5RH3czdZMV4RomaAd1WVYY1MvQnUohsX9lZHJocYTSjnFqkszyNiapFsFeSom
+uB0LXnzK8Bo/9i+iszaO5tJKvTxAre8rgvEsi0GI+zSO5DjpeFf6TxcyVe0MQxiVS4JlHDHn8eV
81RveIpMyC7k4SfHwonYwk7OPccTm9dTBskOJ90AHU3OpgerXogzK1dcF/JHdqMJdZ8qHjpraDsc
PcD6zi184nD/DzX1zkrPjoZ+vODDhZp0j45Nl+BGaextPyMjNK6BfzK0uCwycSkaLoSWBdG6BeQF
HKc0PQUBdsEiPkXGj6/gZf6aOsoJ7E5IVG1XyQfXhgyL/2CzoZizQVDOTwFSERFAw37G5lb+mVct
jXOnHDKVz5P1xXs2Td6UEORocug8sv7FBmOCYUqWjfiIppHLPnWX3+gVuBVTX1k2efKzuoNXMlzC
Vtc+18cnnJbHurCORwuGPLDam0B2kFPDNkPmmIauNjPJoM5pJqqGQDPKomTqdQP5TV6fGn+sIqy3
/UNM3Xgp9gLiDmDF/8dijpAKgBQhMOv20ZznvWndeFfEeGpyO0BjC0jkxCHG5s9aa4vqmScB/jeg
G+Wrir3wcFZ7/ZJlBPYlXjnDu/ZQZFCY8zCQZRO3BXotOgMG+WYf/6m81pvNUN7VP1DMHYnF8AII
XCE06oygiElUhBx6xbEOlHaqiZ+AgdaMnficGg4B8CmVXRvE1GuWiKkoD4CaTuHbIeYL76/h10EZ
+jTyYYvNrX7OUMjmZFSpL8Q5aP1e0l5slPcO5xNi83anFR6wHlI6KDtTCqje7L2isdCxZWLZ5hiN
Bna+CIMmWyTtpcBJugpAjD39SeE0q9fWerctAh8voIhvJPq0WRffch6qd0RDUuNgOEpwGTxB+27g
9ZwYyqhPlQygagOUSqvc3j0r3NuEZdv2tVTrKFF9cSZCxVBev3khVQSBv+63CLdiyGvWJsidJz+2
6fSnS8IokhvVZmvUkrLHSR3rtnLLQP6WOTeQW5Um8rzBRyXoHWY/elyzlU/9sO3nR3A6lxdi56oM
RbkUXQ6mJy3vaazCcZEjh9OoetQ2xR6UkdFkv7IwjHG/m47GxSxLhtwq3iX/ysgpmrUc2dyZ5Wdl
k9E+TwpCwY3dG+nuq65dLpvPB7zybvG/P7zMXkhKm3wpMJNNJCXHC6QvFOE96Mm9S+pr58e2dQYT
8kn0xo3Tu+agoK8qzuVDHEyUrfrPIhsGsIv9v4O+1z8tQnO7C1RHFXfBIzYyKgE2aakH21hV2w9M
rU4cAafGMxiEqmjsB7OtRcSGVfhAkLvQX8s60NnQpAF+3YNkuvpZv4WBb8G6diz6oi3qwQJ89z89
Q2yFq+7LVxCSZ5V4wltrAYjEdzYyX4gniY7mRoF4TQKhO9qc16p9YvafprU0XGVRohq8Td5RP/sZ
ulQ5mqlj8KsKNdKepuUfVoOpOSDqoe1a2WNlzBaPkVEhZEtqGzLJEtWwDQvG6JMuRxTOfxHWacaC
zOpkuiAAxo3UT7JWqkcyOkIXsVDBhhSKZxEuQ1mnAVQcLWENk4ZrlaWibTSrs+5panZm/ZnNe9Wh
XPd6KUrzWOaIzv1O3xTK4ovIeFdmEdpzCdC3tYTdGcGwTKzTdhBAlsKghm8aK40pg80MNfL/9DJ7
d33e1punKJUDl8l+PA7sLoCguFrVQ/i7VcSk+EMecpEcrnZaACRZzQNQo4iZYHdYC2YzXo/uoXW2
PC8M1qPzbsQsiCOw8m5Kg9p7O7Qslvh9hme95Rd4JBys8n2AHdIPVgzcqq3PoRA/L7c5BcdgzjiF
noXNDx4Kwa91lI1j9oXLQ00oXOH2Pyq1h2FxSn98GYB8Hfl8VnNA/UDQx1Df0dDQwXLhEvZFIfNA
erbrz7Vu0Zzjo7t9gcajrlTAHjBQNA3uBu5gW5VBs5zDw8v6jaLAdX+DnLxPSvhP2sy8O+x6mt2Z
+j+BdKut9ImcofX/cbPTdHmBPN+Z4PQDkMiRX5XJV2kFeFQiyDOr4wPAybm7BMMAMoRMLpQB/GWf
QvZk/6hzkV9y8Rl5+2+Rw79vl4hHZu2UWB5kWrDsTvrgqytH3Y+QiFroh1NlQEvcZG9pjALq3smX
N8cIEDsZ4+Mec0EQ4PWjfDVOafdmx0smQJcTosg2LuP1genS62fmyRIzqZCBYLM9HBhJ+F3fo6BP
tYISb0sYLpx8hd0Ml7TCdBBym34nCLgWR/DYsRmvWCfpaZcyf1BYBOalBzx+iBLdMZgoUjINSJmE
O9Kr30WTGxjVrVAJLE/mB4ZA02Mm3p0gB5pcC3JQRD1JLSifdbhaALVlIEApaEwPaPFTgGmyupjh
mMO0VP9klXrF2PT3RDjjQWZYdONXo/8fkIfmeGuH49TqlVD5TWvOiWpqph/JiXef9yDHA121XmAC
z/D5XaOvN92/Od821OR2szMD0EUhQXebljgvGQ3jBBZa3CeD6xxcFbEwxVilAH9d4404SbM+fyOV
Q67lNTVztF6HtdYWeiYFZWtEUsqjRkS+LA276kPSRxYMRL8mgYy0RU64eaSaAws8rAOp25d4T8AW
tdAbqGhFi/s/Mjb+opQ+P40Aew84E3MATd1jQAwrmNXls24orWHIga6ieE0OLZYyGKCqmG6uA3Mq
3leWSgK1bM0OO4uno+vfUnr0DW3VM9fE0Iua4pxbFed7MRMsTqKt9TmyzSDOkFxrEF6eP50xgbE6
vyP++CDQ1jXuQvytLTLk/Iqygq+3v36efGdnxjMhOce5xmF18T9SOJPTWkhV03qId49e1p8xbPMh
qSDN7aVHYMqbVhHOyPJx1exKypPCJne9H6t18O3uImLav+09Nb4OzPCBVo6F5accKS9h+rAjg9Ja
btBFkDgAwLXHXkgtd0JrZA1E0YzNN9aPvfLCBGTSBQKGdgaA1IAkTjBmVXu5u7f+zA85RgHv3V4M
58OwxW37b+GFLPV4U9sPskgQnul+cG/0N2OG4U2XGLVexRJe6/+1xGK4pWtrPzdy1J6Do0AftUab
GOiCCliLVR4F+g+Svx0sGSTAxOvkFNkwySAjt0Jg+hntqrxVT5wkzZhSlYLR+Prm0dqUI5Qw8/Jy
tIKkPhuKgrIRYqhbfPlzTcGOlOqhOK6KwKjPXzTShP2ztPubWF+8QYfhgN0zGsyF0kfW5JSl+Oj9
NvtOrryqOx5+EzoJpn9abJW+1oPgS+yumrew48ZAoJhMadR0tZa4GE/QrF9a797T5zE3SVmWrBzx
TYs51QzwxKFNHDT2wlDMuNDIWY45ZMXI4wwH9/XmlWiSpmLugU1Hideta/GEqui1sCuPPpUN9km3
ENcK3I9XhVfnuZMpsO9HHip+TdDxqOrbJWsi1xfW+UNJGhzSRAf70T/Lsz0EvDXbbLema5Ls9jT8
/LLu2toIEz9Aq96uRTG0q6+BRmhyd3sF1GY/W3pLJR58Q2lCma5CNBCp3RVERIf2pA0Pco7msjSB
DSv7c0Q5huxcnbHj/BLs65MUiyCfUaAku347fZxXybivAIlkB9+kpz1HPZ0yLXKftDN/MoSJ1M+Y
7EG51QpehGAGHnzDnImcF9wv6ASVxCr7oyXh9ThUD2t5qJaG/x054gBkI5kkCL4NEEdDNRn50LIg
lns0zS3JV8vDopHi6BcIGJITCVtmVzkGcQc09z9GH54ESHfDsNGAhjaa2iMX5mxP7GOWJsRV+SrQ
FsZ0od+k3JPL+4MkmOdoc+RAh2fee0XJJ7u0wRJQfiiFwLy7yooEZhaNbDAGz/t0MZ8C07xCEpfW
GQwevEQEWHX1xDZ/uVHJUyL9sV+pD5tRok/ww7cgnvDLi+5GA/R5A3BJyoSiHkGYUsjvMdnsEltv
FRk7ZPe0f10p64qWVLIaqrL7EaQfwHSISDIXjWmgrZ8aquMqQLshqkvh4sUjeFzuJ3kl+f7zTvk3
13OW6ZPhsnjUL5do0zxHsMFh1z78hvnkdpEdbL3LSq5C6v2agOB9r5NPfhn17kODCs+m6Xy3Hg3r
5IA/OupfpRSp60RqwMI1vObSpVutL8LTex/O0WNEGRFtQ+sFqAEpdUExFfINVbye/EyO4t2OS0bY
zueGM6XMQMKq3lZYF+RiVj+h3Q0mBaB5tc0diE0UFEKw1XHtO3PO5WW3ED9EdUh7kVqL7sk7OF4a
yCnHOoZsMQM5nnSGaHkpyZPIziL2KYttxFhNI7yi/W4oZZTPKCOaMRCrC8f4WopiQIBXd5DesMMZ
i0AWKCjpuhg4wCKyC1y2P0Pan7L8s4HkViwlrt/MGAAr+mT1ySTL+mCpjMn3kxpiWyECmvfKXSvv
MOSdauTlK86exe86vi+TqxD/lGShAolrjAVnwVdPUwkbjkzig6z61cqGhMpipIKGRN1UmF4UduSc
YE44Rf4ysoG72pxMilng4j8neYtkR2isPR6O0untQxUbeYXP+mQp3TFtazbdIKCvG6Kv5N/sKDaT
wRxcVb9GJFb6IKdpGe6JKFliDKkGKs/k8NnT8VxFI6PfoeWs3/8/Y+lVVPpmeZGFdo0DF0vk0hVB
kV+/4B1CRh7UdEd+bbiQbEWWHLD/+7qRW2+N/4LuUmxkJTP1U74mpKCB/5KErKzHCMAAcmZiRERn
xQ1gDvwKl5xIPQKX98HqM5oY7FhSLEHoWmvxM1F5JxAeG3fnR1gAFY9AKsNTe1cS9Va+G1jmi8HT
G7wh33iNj0syluSkJSzqshCJz6mYqKUHIzJpHlMhBZz4dyTCQC8yhH14+o0c5bRKTbcidL13Eblm
5PZRhouCyZ0H5LyZZuzQf8bMNc17rIXtTe1LJGg0NA9h5l19cCYe6NyGlJreWLXLiEEQpCHBG05V
n+3BfmWtcR0rr/EBFvkwtubg1sIHzTbCYQctHpaZNCqOfPQfYDqEiIx0EvYeoyRaS3dVK2HDHj2O
QTjoD6yb8WoeuLi7oWBgwfUaipPdkm1hB8McjCMa6NVZ91Q+R+2Fvjn6bJ/KwJnnWzLfvnX19QmQ
kzxnh+2AuOw72kNbfZ8gLnGZqFToXghScqH3DQTDhab/A6TqNwxWh5vZAdecNgwCxeojRuvA2LfC
iU2GVlJk8xvjsDfThjNtZQ86CeUn09vlUV8CTELd6ICHw+oRqX2GlMf5sZnLSFde3cDHVfF+Fui3
AzjNhQ5dXgxHvT9PbxeuOWpGyUZaeiajLoUb8PUBBLW5aqkcKAxwZsJEZXvVENGoQ3+/9UlozF/8
6NnC++WZrPTxOmIyGYbicfR8BFhWGENHqRD8SvA5/Gdet511rgbKK0aLQIFXhLv1J9rzgEiY1Ito
ac3CEUTuwFzdDl7NIQuBfPh2eqdhig7uVWP61XZRaYEG2XPbF88R/ZXgmyPE82xtRHQ5OTdMi1OV
AN60UKf/bssqGkY3jaAsOmoQSuw/U+rtxEnDrMU1APgc9Zf6G0jndaRK66o3sm2QA/YKfCSJVcvQ
SLrrr8+m+ByXLRKjVHAnd/FKSezBdnmA2qBQ0RNo8MzqNNCMStpxV3uhRXhL6T3LTfLimAuxRH+y
E1SD/QCnhK3EwiRzDKkfuWE59i1dJas/ByeliUyAIlc8c2+lne4e6J5RJeMPUst2FUIK6Ja4rO2d
E5CmRH39Kp/RBSAQIgkeKHcP2FHhKvnlMZ2ihLBV4Jo7NnvGZnPBgj3OkqhovVMZvsCFDU7FIaY8
v6bE5EimAnp1/iabVmp2KNYdOGTDqci32LuybmUrh7EHDxcWjvoHmBBcLIjDcvCOeMDAqh/MeZj7
8WkvEGgIaitaQ/61S+2hdgK+Hbk7p2qSVj/rbkaPVlYuvUmZkDgq5ZpetYYERH2YMjf+z6GQuT9h
Tp2B3ARbIx0bszVnE1D9OBMY7YfJqwV1j29SRZX/X25bpinSrpvh2Md+IKAULiBisnfHitF0GfQz
csc3iNcfdRDGVYqccOcpfcp5+NZliaf5n6j7EbsdpEnokxh/e1NEl20S6woZNnS+cqoQU3M9ehqg
h2BsVHM54erVivmZwgZy6e+unL/1Si/fVmHV/g9gxaQH5LtPemfNDTbT1Q5AMm44xgyvb1mOG7hS
UAdr2pvhc7sQjRlBc3BUjXIByEXE2CEHzqy2DLvNIN2YiDjyqHML5lcM8MXmYuvlBdXF3Gy1da7/
OO+F+JQZNXxAcU13TuR+AFZv/XahVNXh6hwIwBfu5P22Nzg53towZw8wFPaYro+Og9ev6lKCLHhn
9k6ISc03Db6XDfmxvPFIMpe6fzc4/9Qfvm1xBNXsAEMNaam38gv8AJwr3s8I6EBQiHW1HzhwTFvq
uKZfHY/6up+Gi1HfTzn5qmRhJnfg9hWJqMfF2defERcTYoO1iEsLQdleul+8P5JaFk7YMjqnrYpd
zocaBrpy4cF+DsgaQaZkmydnKkyEbDwooQyednZdfYXqm0DAQ/9mXBWobOPmP+m7wOCgfdY8iUPy
rrd9HErZ19i9QAKJaGbWL+9Lasi7sY86nE5pNonVFObu1IVGRvhvkwbeYKFhzZbiseYLbFVxdViB
PyrwspfzKWwzjM/fI8Prueq3SgJrrm9DcSzr6dSSit5g4fIN+bJluvtWMcFGbQ5F4BU6LFJSzFBn
5KnM5S2j7dygHyRrL3EyQKiCVq4c8OOmVG2Kq6rphecc0ijLyCE/ulrvX7YVQtXrVag/fXWZ7BK1
8oC5Nq/uV0GAmlfOh8ea5HB6dnBNY4zxev5gdE18yHJt0j5bPzryXeNRxG7jTLDIcCbQnmwhgijn
LYew2EprD1dPm3hesyputZZq3y+NDVTnF46WIUJH3TB65laHpVV/GtB+KudPhU2O7OyRN8C0Pwu1
zrk9jwkkifK+J06m7mRs04I7s2Xu+/Alu6fDu9veQ6QTk5aj4upEFofWZzPGA8ELKQ0GpzU/x4xZ
w3d1LQvAdOAqGq5NxAZyKRe8DEoHAmyqNHUe1fI7T0fqvriJGMM2vgwd2Ra/4yfIh+OIhpE6eMtx
/2eK0LB8ElTTme5Ub7ax50gPLNqoRB06kJ/rzt6cVmx+re/Qzso298yFL8yZmgV/Oed0/OWQOK8I
/P+LgEmzKKTi5Oj/mUgMePpDNZFPZtBxDU8hQJcUfw7v1UXyChlfObkcVzcw5HoEzZjPXg/bVdm2
pF5rXHnLEyBgkqkRHLUh58hLzDThJDKWvt4p84VBGYIDaHt00xfQlouXTv8hV5k9wJik8JQqeZpa
kpWeA8IEYepgfalPeawJIvKjm7uDumWbQ/gPkra7vc5FtI3fEkOK5JvvQ2Ew4p02sL2zPkz4660v
KVSWqazqRXE1Q8vPTfQrW5Gsb4UIM+lYS6B2smhWoTIk5xBdjltAWSoFIZh0JViZRT7MXnHqEDmQ
4f48rmGk0t7hRkfUAXvlnETjIAId1M71DGAYHkNfkPObid9GgSpeIs+kVk3TLzAzGO4CXn6DSlzR
dlIT6TtA3/ICKzxOlPKyt0/KhObrklqz0ZLZJ+UnPFPzGMgyAJK+NNylqPMs0oqASxPthyuxnLm/
nONje5ze0BrwhXoon3eD3Xu5yykctt7oP8dm7vAS06AAEVsopHoLiOvV6im+t4+A6eg7iCMH3xlH
yMoSVtMZgngOESeJrSdeFBHRm9ebeYSogYC1xoKxvvP6JB5rlS+TBqz6WRKkMuXAWejRDT6fsFJA
+VpVVauKMK8mHuxGR1xqpGGdxwqeo3kdPCTahw3vBY14ZTj+v4JF5TDhRVo8p0N5X7ngY6/SY8P+
cPNvnmbjuQkUuiN/szroKFMKX6Iybp93K28e0u/N2K2k5eRXSqa62dcHuXJCUSmen2gUHfe57kT1
7THSRtW28OtEaxSvTffW1EqH16NWRagTuA+8DHXddffKWTMPwOIwwNBMrFTC4sSSvc6kRm6y5rbu
nbBggJwmd52JHL1IHZCbSPFpaP/T4WdYyxF3Fi2GU0Cfavqv6yvSMddYtGD8o80KiB2cStsXCaWl
egjyp4lqFgcGCMbwquzPDr0BwLQJ/vZ5YCK3cBRhv7OMgVx6wWH5mtf/Jd6xDJb2j8pB0Ctl4u2X
VnZT4Ixp1U5pWv3cblwj53bK+Wv0hd0Qf5oT0c9BPrpYiW2d+WTN9zBxhMI1WZ0su+zmFuhIiqwO
DzGpbUq2yymLSHm0g/0uCuEs7c21nK+aKkBgG4Tb/mkGQECiZ3hNpBHUCLi4L75R8jjorb4G8S6k
UFsBluWm5fuFQ1jwB9hJkaSbE13Q554drcp+8lr5zUIN1KhlI3NMX/04mxQjD7bzaaOPhHRqQgDq
Qppgz+ovL2uj3QvRdWUanMXrIrzMtnNjxXsdNo2WFgOamlLG4AvQkxx+CSkwPeLAQNp17t7tWgz2
b/VrotrWmcLCrv5UAaaO+z1gc49nS0ULceelPmBZL2S54n2Ef0E43CytXJi85USLOVuQXg7ZPSDn
fqIiCROkMWOW6GXIE+BHfKWYlJhiKP0ITNUnFcmigTX9+lsWU8twtd0tLIUHiQUG9c69KHH9ec5q
2Qi/Ae0deFDMdl2fGeskdj13BbSwlOQv6dKhAuY65c+rAFO64I1awQnifQDpQgqaECjRrLL/LQTH
LhShUtK2dYa0Pzq8cSbIHkaf7GuF7aVgzT6qDlvLZJKvi9r/aelyrs05fC0GD+ayw5CK8ONjLGe6
kKDGo0gZvM+3UjfW+zq5NUT63FvRV19CJDsY+JBjUwk6HMRVq/kRTFpZcmYlo++rOCADd9in7m3w
xaZisens4ZRQRQVBNg9LrsfyWXvNpcTXhnNgRkVyBfODSMEvGbtZDpQ3SC4eIfSpsrZ+XhYlDYxw
k8soqpAttGb+47HUm1Jh4JB0A4F5G7/cYz9mu1A7I0SNAr/988QT9Rc0guhWNYa5NTUdmPcuErWV
8X+SWog7tQCty4bF4EJnzPurwJoWoLF6ukj/+hVX+3osgzN2cZyt370yC8LjrIyn8DYSnCmV5wLg
nKLiJSHfgBDvrYb6kE6POppgbFN4ZqXxc8HKBcADZN1We/TRBQ+gyW3VXIm3MYLpFMz2dK+/pB5u
BMFQBPmIsD1klgeVtcHMreeHt0H/J3mxMq0SWw3Qz3zEfqFaIDh85m17vs27HPkRyVUQu82tzSbO
G91WhXb1a+0MoZJ61eyRnqVlHEJa8gnTaKycdJuRotEmjoSkaDXfhqMXpJUwoI6eyXuheB0s1Y0M
ixdSKcp9Af5uOx8k8sJcdObXMShbAup/xQV6MWG5KITbj3YxMiuvGDccyLCadsbgdv73l/9Sw5LD
gKBRCtnieEDWTzikpW1CcDLglqhgRVAeR4RBCYFTYpd9/ZVKBFv8vhhqEqot9lw96sMxMRoLHyAI
hbMSByCQot4DZVlEWeJwjR57DDVkNZPSMb4GFekK+u1JUuat/6D8pg00nYF4T00n9zlYu0iU0WCL
RnEdovWBNrcKKNfG+z3ZO1GtNYPgqWz5GeQ9Sb6ow3be4mad9xU2ZaT3nALtZuNRoEwFW4VZ5jbT
VBkivFy8r/VdiYrI/XamKAaKmXaigbGrWsaF2Xk7Q0gpeT3M91/CC4F7XhCp+r3B4/yc7gyG0new
r7D2BwS8XLc+NHZDfibqDZQcEgVCeXbw6vHwcqJ+0SBZFXSAZDHLhNpZ0CfQh2UWQGmi0PW6bXlr
mlePVW8nvNA80EMhl6yMDi/Mzsao6InoMKmwPkP9tvJOhr6cFjWIpvVqZGGQTkqxCgBMnl6Xr36W
nQl1IO78A4WuSnXu+e34Zmimqquh4TOkMPZd6YFWjkm+aA6CCmQ0dDrA9spr55Lpd0daC9hzI20i
NOT6IMO/dIWdiS6MINP4PVDxf3GMWLJOeLYoJS58Mi+od6sQjVILtKtArBy28pbIHNCTwI5cpEfE
DnIl6pzPKjtUx0zanq6UGvNUodTQYJE8pRMFZ3ytVkPiiETkTmfUZlIKXVYR6LU9/nTAuSMxOeBn
6H/1D1G1ShOfdAXnZNOM6Gh8I28owO/ItilgUWytWFnGxyR2Ldc/5TUb/mcVo5QxOh0kb/yqSDKN
0SILY7C39E01YoiaYH9nIOwULwINhgTEHOWF9FzYDsepySrX1XZnZXDtBHvQ+GYD5RpRRxFiSlQx
w4tSzaO38VQl6WESDzfbywwoCqeEuea6XPzqAsMHgjhiZfZX81LL5IGKlYolprLb5P1qbKjQWQT8
lC8YJFJqw1Yv8ckxkeu+wa+MWW+gNp+TOiHjlVFzw5z64T2iXCVtPJvAySJqnsONb0dkdC7GDr4L
rRCBdYA3NYiFkIMh9FvLVEhwEmhS/40h4tzeA1CNUBz9lNWcHGTWeTh+OmEhYcRXcNwLRvNMbVdj
a7TGZ4+XQlwfzWrMnx2+aFkGPq9VdFp8gcQn8ZuvikYr7Sv8yBfRIp8IZEJtjaT14FcBVBZCdIN6
bKdEb5BIsppbNd0cQ84agEwIbuFSbnt2h71l9Op9MCBocnFDwblPjQcu1hPm5VOL4ty4wvtt3RML
LyxTii188JbS99pO+codtGt7y08DuIzO2SJRb0vgGGliv05K8cTx2YD26JNnWyL2QyImkT0sMZpF
Zqi8hOX22mT2RRUCGZZIxW/GwBBpOPWGAvlwL9T52Z+gIrrSZy0r6uobTMf6vjT7t2g/0a7YUNd8
WrnZ8fLH8vHVXNIww9m6NKLeDhvMe8ESRYTw7iQDbCo8NyHCB7Wgkk9uAkJV/4/ZQbZdwmq/zf4V
xM17YhkENWx+i+tTVTFztOqwUOTmICbN92AW1iOF1IxEovMNiVfrWmWtTUomjpyrYBm4cv4TCAy8
MHgD5BrqVODbosGLbWaBas+DE/+U0tx8jq/szFDbnDv1JDuqWi4DbFFDBsX0id+D8CnJdaJBNCss
lCjc7zeryOPwmqlilTVHzyud+rJ73qMaS9oI+qTmaOXHgL7KaPaMUKsezNYfHIQ7g8FzsVruXusS
RL2iaOsJwJsY/kjEOQgMjUa8O2RUPmSgKeESRQdyxrS8nxdMq4cCVsJyn4lj0JlBpi4PmRk0vkX3
xogFi+q2GEH1EKGWRQYBUZHW4zGMwzFdwElUlhXTbdhPS/vqy1Uawc5o5BxECn88lMevwSQ5hTAY
lXr+zVJKOT+Vc5rXwW2ahxOhvn5ERrNJNfL292yXog/ivpFuH4jMugzMUgpvwWyl0IowGLxRvBjx
CqkhcgWVukz70PheLFSidz5D93agBDh073alK49rfPVLGN1oCcS9yYhU899Em/N/NuQMrbjVKVMl
WLyI9SmTrKKlODD64HLWxrbItXi9IVTYQCLVDylcGgMB178SrCOF/xx7ulpJ0TTas3+qI5ZGgLxn
2blkEO1CeAM9gdAzaW07XLR6xB45pfAt3ubWxz1iq6v41ZytyDSgtf/aCMJiqNlPPnOyoIfKR2BF
ZMq9+iENjkxpo/OcELNFnZd3oL9JZGzDp3uEd0PmuELD5xOolBB+AnOHtCU+xm4wQyxLvuIPpfHI
ISieIPva/OkrK5HNS6arPj/pWUJ40ONJ+j4C+uzPNbj15sqab9inBiceQu9zZqhSCvb2ZJuRPSdB
/3X+vOFtEtjcxT4srHxg7c16ZveJh3UGIXOW9Tz6Gux89/668NLyUre6jbv292MVAUgwr/tJgnZv
u5efkobbvcX/Tsh4IPbTuNqhBeBMrSF0EiVow5rctP+dazxutF0bqY7NaIuURiA3EkWo4mQVa1Tn
ChO/eL2bPBqFJErYCJPjd+hiWLlNgkHYZ0PFVc++TwTx9fsbYADAX1pNv+RTo5gb5I7S30OAYR35
pO8VJQRZYe1M0sR/cXJr/58ww3XDyRpoU7DWXJQ1ty1wHWlaAvtizLpAgAiStcOOnOukQ24YXpiF
0R5ZZ+zeJ1EzTC8nujfaPqs6nXqb4SWc3ZMzSB+1xaWRzbcjpEw9FEDGFbpuCyiYidJRyth8Ih0W
xsvvzXSGvlydy4d8anNDawTrJ/09MqACAQ6tYDcnhbt0axz3cswcL4NzKhkq/Juuju09iPexzAsC
nTBVwxwXX7tIRwMoQOmFmwlD3Y7/EUaEx4tPHNl6nzHdLORNS91WTPkZ1y3W0H/c+46jsWO+yRb+
YwRWiU7Or1EDEoARQaaeKVxfr7XEbpvISInDzOj3CU9IPhyFm8bblmohlUaT4uRCE9nt052WyUT+
KRltdg0W/TzgHhLEDxqmUTbl7MZwQAyxuVrp+BlPWfcwSMDg3UQOp7BskcnNI/3I85AQOVaonmzz
kamgAex7KI9YInVf26WjsCErVGxU7yVNUBg0nmxbZoknY0sdcrfUtwFAHrMLxZGLMNuFH5ux3z/1
CklHGU6Cvl7xAWmdvbzSVswpXLgBKevkyVCv36CakSrltVmTjwfaQXs0Jeg6yXI+ShxOfZhOh4Nd
vb99qxwrx6IQ+H/eJIMwUJk+QetGqbWNKdiOs5ucjGfyuoNXBPZZEQBY9P3JTCqBViO9Gxxnb5pV
oe6dZDKtQyW5cNHpSCojtezEYrekg80fXLpLKyQ0CADVRReEVnrKr3rOyhHBGN/vJxe806DwpyZu
9tEe6YqcARTLjypt2i102QWWDLcbZvjUzeDvQQxw9Dp0J+A+8qfFqIkl5obsYHF3kKDeQHC8/Oj3
4Dob5BOXanyu0FaGioXz4/pG/TwqrUs/xRT8+3nlgcFJ65TF5b0nkC3U8a27GXEt6jE2JqL3svc1
jxMyJ00a9rnHjThrjCVb4uBU66Ekwxx5TaZMJrCGUgVqlK8zKqj3QDfiDummlIyRlOy+VdSqwelY
poXr7qX6jVf7aoQelXRTQ8LcvavDxTlMMbxU1O9ZfchinYvjV0KWTefs1gLYJfOHRTnj2rZHxblw
bcHDGqr4a0NAMc6d6fMBgBaWnXaBP7wAOyYDM1OZXAvTFSTYzKIYlPpDskvl5fu5Dpo+AohpBHe7
RITibusiB/+a7oJhVFYdffkWogEhU61jbCgSWzNC1I2DHxhwc6/e8n1RuRXDd7LFEX3T4HIWiGft
jmMUZFqDkwAPvtlam/QEzma/JSteYnusPrvcXn1UCcbp/Va6RQ+9wlO6q6bfQ7ho+NyJB7WEQmBA
HxJVl8QSRBqGBGk+5k6VSY3xNh8qmxuInufaM9rKB9CEqmy7PvRvn34P0mmrRCm9ZE6RyqS7WwLR
+9I19PxMZESYpbQm09oxePpmpGiBKnfTyWr34NuUEqiJebmcldKIIRt/8K9WvgMcBIsYYw3q4Ylb
KpeLXBR5fmzI4wpn0g99GjYak6EY8jgE9redT3ioLjKS/3vG36M4hAX/lhUvOLT1h7O88dVNetYk
KXVFFFk3csok1R8lQXFOOmtxuaWPTbU0RP1fM/CIRfvrdy/Qxb/YULocIsBx68pFbTaP/tevpgiO
4lBLywDpGmKea4WgtEUvUWVk26cnTLiFn4Fktdq1cvcSPCaHrd+BbZeVSpjgbc0ZhzVJ/3G4CF6c
Rlx6GT57JQbh9+d1MbKEbMqfCkB/AXp/uGWbfIKZMdQ9GFuy48gDPXtMlkfhushRLmPZOaTdUaX4
QAV+QyXDLxrtXIvqG8c6/ZbmZGPTUHLP8XSnZ2eOSogp00rP6rOB7Lgdv8YmrcZz30xjoBlt/Koq
/umMW9O+V4CuCDalYWUV60cJ6iix2UDkvLUs+fzOXmhq9HnkehY2tAwTrQO3rAiaQqYc8s5ASUwf
E5pFkbgs//XSho7EdfNekc1U9ykUx13KMGSC0fhj9Iq0aWul9iNpXijjsqjCqbseCP7y5YtGO/ro
A0WXBJmfGf0H5vKIynwUXy6eOIIhiefcG0KUA2VZVOve4vBJgs2uSaj7rpW+li1yGGVQHjycOdEh
RmAqA9G9MDhry74zG3TqbbXEuwejdsxwTAxtzeq4Nd+UuR117eAr71qzfN4bePStWlWQTqc3b1Ki
/YlBGsl7iT+q2YEFvFoW9K6JDzHqN1J9Y+IQgreRadNHRn3bJOyJt9rD4FuSt6UqK8z50gg0V3T1
eA7QipKm9Uwn/zlBirnC+QUZj2uW+us0KXTzeZcQbFyKbMgHmtkZGVl4PJI+L0bgHEzePq16LK9q
2S7V7N5GzGWb7qpXfnOcjWef19z5jx9nL/KOdLxG/z+vc3DRcSRE1XmfT6Sjc1hus52JSagpkFIM
AvE+BvkGAmUy16R0gHj6zMKysiRdC70mh5eW8Vbjxp55VxWBr3iS9TBz/w0/G8/cr93xMav+9GGm
C74G3eGggVGGH0y8aS7Z073TZpIL7qSex921YQ7x1RhFUPuvCgxr62Dr72q08bZXKMDlUlXS4qi0
Taj5tGOYFQx2Bxpdk10WuSO17Z1CAiy0lceB7O+zPgyXgGoxD5P5aw3LFW2RJ3+6Mw+Uho4nQpUe
R/3WDMGDVlbTHuHVuniGQqIOFNDzI1JfdJyg2xn/bPIpPZoR9FQhiKE3RWm2TZCvsdOmozZ2fX4R
LKxj6s6JpUKjY86czOqPh5ikTB72J1QaDRc8nhaRyjdarHQ39Pj1zmQUkCY0yW3qS7l81WEFf/x8
aexOWqze1aV/K0Cd+s2Ft423GXsqflrdfkqFFYMQJsxNCilrtPzkpmKrbR26q2HcC0t0xIspYIQ/
Xxlm4edElJ0hzOhOo7me7Kk2vJ/eLTAcJJ3OsFzlk8Zf4FpeSupm0B8P/FXV3uKhvWVseTP6Fb0K
fJFPNKnRRl04EPrURldV2yABLRUmf5UtLiHeR5uIRxXB/5ERwTZijRVFBugUgpgU5QzuH/HLisCx
eUgM65SdissyW5ciBu7PDwmXUnp2xtki8rCn29s9ESMXI3CwD/JrISHqIRGna6Iim33soRhJ64mC
hn+YTa8WUow/HY6Mz7jikJCrXatjKq9kbuU0J8OVorjuEyn8Zm+esz4oUuLPt80GLBFC27nn+/X1
XE8D6DL9hFQ7LmJ4x3zWVrRxcuy/2xhPava1BOQJFEKM0/Xz/oYPlEZ+nK46JMOJBWBxlsBIqmF9
6WKozVvAoDFY5/cvyz4a3h1a2/ZCOoMrAipADz1OgYgcRZvwZ9+P8Pw2p8YUespAAhw9REe1efNJ
aJECyWZ4d+5/eDBXwhlojpMpB01WNO1pc51IPrE6NHtNJTOdFTgW70GLYINTbrF3k3e/w/PoYiWZ
caBtS4cIp+6AhYz6snmVWZ78Kk6okAQCQH0PGommlJVUdQBGytxwM4q/7OlKTmesd4ce8+Ytf1U+
99E5v2asHxmY7o15+0LT9K88nQi6w3QK35vEGxAZDtJol0a+rZ1EEWn31gmNW6ABBH4wegP5WCfW
tX1o468KnC/vN7p9afjLHXHBsPPNKD3kak401vnzbznRg8fBb9H68Co2482m5vbuxPNGbovbpvzK
a7DRoOqlKPNRHeWAXKTtB6p6MskdIkmXX8JeDRWXXUBURFs214hpAFX/g44ER/JUzMTlW1nMOXWt
MXW4/eEd6SiGJFkZhKXYcaz9/ogMFvWhGWds0iXS9PsvN0h/M32pIm6m/lmBQ+EmItbbxaClx2F4
lXCiYIyPbxbQJWdUGRnGLcUR8ufDIJeG1kQUVOeZBT3QqrIPnwHb1ntzV8NSdemtTxjpjIbJasER
FLEsuw7Z60gGQxzWcjlQk10nkdNRmIfXg17f33T8mSqSORr8ooOv1ZGreMrLgPZzpDGxvKpa4yL+
ebKqliqJ3ZmTZjnPvZWsalsKdXz3eqZO3Z/GQiHdriM0BwiLQ+LtKpS8sOLk3pi08MSbJNO+aNMN
8m4fSBTHIsSLFs6MPCh09KkDJyHlygI5CrSrcBAZtN4NPWjVplGkvP++K7Pp6MdCjQV4iD8cv2is
H7NuAMssePwsPKXLNz8fnHU6Ceaq7coollbngHYjefljHliTi08monXhMK9G5a7S8ofUjQ83zSSl
thijZhMCPQk/8VrOv3t4fl4UtG2txLTkzGxDzW/SbL7M4R339o4EDBOrv2WGSdavKrhKejpfvahp
KmDrRktHFKARhRa01wYGO1GlOJg4tptT9UNZOAvCCzl6LmfmnfEDF45KoblEMdsqMxy54b0VcNSH
ktDwx7MC+op5qvkBupCqldyPnyzpdSBoIwI9Lpzx64xHrcB986LDc+CKTeFcNeLJ9Ku0OUw/+P66
xddZktBO5jzERSskZ5er5VhtRjvkrpX2JldAC4WUZZ0wVoeTdn8ec6c68DtBdFXA4y2YqusMVwL8
dgUvGT/3F+zAuPhDPW4Hl3chPYBVx4WIKzGvjLsH5fY8FKsi6a9f3g2YZ10R9/92D+rYaGmDxOD+
6fGbYEDx5K5ZDs8ml+OrtYLWJDmNBbKHYpWnPUw5o29wX4QPJWMJBxXefsOJJEg8F+lGIthjxwdM
apd4w01fhBb7Wd5vRp9Cd3Gmc3KWWDSuyYs7fzN7qjpZ2iaJSoqv6EXv9vfAnI7iagLaZoHmD9nv
7Jx0Ur2Fts3x5t+Pazaj5IQT+WtI6kj3f719lzTtxnYRNSXG42ubAMldgppBPyD9hPZ8W7fxtvBB
FIPOSB194I/Q68z7K9/xg9DtPHvWvToxHYCkst9IglEgssOqbdfuoTNXtuUz9xhgA2hEUfFJOriF
nKC/GqLMxlLoEtJ757BSExRUC5t3tqJpMJvyuoPu3z9udkWoSS6DkQoxgPeHGA1FS0oBB1e+hBVr
UEWimSxwr+3SG53mjgUqcUY4/v0AUZ69uL3ieVurmwP/mJ5BnZQhxqZSYg/0h585pGKRj4FRIxEr
M/Gn50Uma97Df2MghafS+5M41qMstz4tK3zjvaP7S4CrKYgYsEaVwr/pl81xpXN27oKKq0iDLgeC
x/xWNTyBaZZFkBxVuaHy5NagQD3OZvTjjjySy7D/q4arScP2tFYzkaBMnnyhSFW5/uel8kYVKaYX
qtXrE5iB9UvQMmDAcHAFBZK0oWGb9rZfo+U2Ht5rPa+P9z5osFMs7QzWlEqqdYk01J24fgw4FDmE
PYwg8JyEhgqpeDQNBPd58aion3k7CqCX9Rwwle8e5ZhUxzU2/B/4s5/SuYdDTFXf01mJrX6z9Qci
YuFPgqir84TvTyl7nQJRXIijGIjZLR9+S1TV9lVWx2uyQbC3ntnBO4btVje4M0mkM2PVjZfid+kE
Sa6kcdUc9irvKVYWQh8xROgFHTcm1tTBS66tf+Q+80dwqUw/d7Hjo0+WTQvTPIKmQDjzsiOXmz9Y
9Ygi0tCQ3N/TqNAsJVRWz03FMMRuxK2hP5pR5b5HH0LkyxlP+ncDCndBf2CQr+lgkiC2sdDCQlVA
CuxGcQ+RkUWxXIsNF2y+3rC/toyAzDCmR7Y0xUOmQOodLRUlmYUU5cM5Hs0jH7eVpSm4QdjHY9GK
Y1jA7R550PkUCnnPq5wZHtPv8Nc6c5kk+oJdHWeBKZCeL4NdbXA7UMYD13E+z/5q75ItXsKoGV2Z
U06zG0LKHg2Av2GiAYw7/XHO2l7URsHe83sAUJ46wI5Mz65l1imRExx0QJBzEMZGbzjlUSpcNLIx
B9E2sJVQz1NXEr5sG2gBWg/oAEQtUrAnl6x1ZkTKm4Uovc0FTmaWMFGpvcBQ0H/uL975WQ/4yOoq
BRgkO+gIis6Q/QoYlA/HZ36HOCT5a52gY2SVADiEOBhodatp0FbsBUvYvYpfwQSJoQZBzNiiWq6a
Sw+vAHyks4S0aYBSlURNaquA6swCZq8k2rPWrRFh1JqhNr93e3wM/Y8A68thI1nPG0x+K9XXzB9W
lQ6l3Kmwb/GfYHlq64hMbXYAYERnF8PVn4y9QHN6JHPZiPPL/e+rHeI/EoV9+KGZcr/udQEpHmd3
zfQC+aVAYEvGEkh7MooQaRQCishXW0mstEujaytHTdszUr58Ko3jTFSvfa5RzFoLnwA8zp7RRAp6
L0lLgI7pNu0BjSRCTLYgj6w0201Raa/waIe50vSq1P6N9y+s7Dlz86X3LtTeBOcQ958XkDNCFBnS
AN8KwxXCHgQNSRd6YGQFVieDX3lt9jusyPw6/W+fXu1n6F6M0tHYBsY31KXNBt4rEhaMNoCDdsYf
XgjmNsL8dbYfucDIbTq5FCxs2aexCooQ6LWnBQj+amF8ulBpqUl9BUCyJVwXoH7pFA5WxGAQ87Z6
SoztRdduTk/yuGobU2xHRdQeh/K2a1tlj3IGOPQ/KZpLvrXHWLZ5z6O16FMy7013oPxjQWw6csQO
plpy3YoihzJyv5kOUBhEHMERefdJ00chht3N0l2s3ox4spfbJGdlPsVTlQ1ed36mApBUyIf67FlU
5rTVl2FL+Z0KVJEXh+Ud7icc+8SBYAiwryjf3Eoey6w3dmeq4FwLlBrn2MdvexaBlMqx72hip1dJ
PwDd41UrbqoAt15W/SThfDpoF8qxFb3hW+GyUOJXH+Q+TCmjYAExEQPu7Nl6bKwnr+NO1/7ABsog
H4rytxVmMUSwISV+n605vO43L2a5TQs2xLT+lkgIolcSsGZZ3CU8cvNNknSoEBLIEE+9fQwMVjOy
/u7zcqenbZhWe0j3Ru+yId9ZKYJcXBUgfRrV0DpLoZS98/DAclGOFzlfJzmDdSq0iz8ltISYbQ8u
Zmhr6tTwARqATwqHVPZxos5vwimloDZbdIf3xYU/XnZgkHo7kvKPwKUi8n282vh65ydBTrqumHe8
rxcM+qwQE6ztDUXL4F7hP/aXQ4fqMQPHIigEY3hQ01ERSyPPi5ZBcGHCO260gKavRGvuJNr8G5yf
Cho+AsE6tclPwZY5hM9oUWYAFK2k3c9eydoLH5j5/RU3A0x0RbbgE07c9eA0W1tq1k22kzQ8Yelh
t9aoGYr+7yBRvzUcr3G+nFnM8TikNRtWQscqpSU77c0Zd9GMChVNiX7zPLILfVwtU9zqXUQiIeej
aEMDZTC7P+ECCizkkpdacgyoL3hqu7sVt8Q6O5WDVhWyNt8QLOvoixM8TiWsEnHMbGUUsJ7Kb0GA
OaR2uL4nERLOhXwtoUBmIJcaSVBEflGbTEnVyhRHgA0ZMcVICbeqWBZb2eT8o3Y2q2SjfdX1MlCp
2oOO8dEXFmZeUqHf/MQCbBo1+AcLKhg6IS+92DdKYFuuiBd3tAIt8ClHJpmxdgB8YT6pilnckC8n
cOgjQ5L/oujvFKN3yKzy2l/4BJ1VCoy/KtQi4phSJfEkIjKERqCFvbLMb7KDUo5Ys2XV3CcPMR+C
0nCc5IWMgAPt0NqvByVZx8+GwTOtvSWIIE63M9H0M2TGmk4evD9oUVraTD2kMqFE9KKwUNBsANdh
ccCC4g80hw2qepJSbmGxedHpKv46wbZZVUK2ni5d0SsAhvjeJag4ouaXclVAzI+aYbMw7xNIOM0H
HiKNJ0FHAkEYh/QSdAT1S1ylNDtSNg6PI5lVkGwMRv7+kdahoehTSVMlwNJRE6ourFJrTLUiCbkt
S3F7jKSkSb3z50upkidMXvCbeiQxFgdNANHCHhQqBuoWe++1ZtQ8Vkb2C6hD4TqRq9G8tMRHeKIE
UM7GOFGoZIRMaq0w5GbhxwEwcVT+o1k0mC/tGE+nhAWu3FaZtXcxdN5jl1YdG/2CbYPvAsk7Nb8w
ffcJkMYFb+OC6Xv3+5CaA9lYc0tA1kApcUG9aUm44L/lTuQWFlglKe7wxyZmzwl3WxbTL+k0hlGV
SQXuXvylbUGg9uCdi/sO+xX2lS9WZjqDl3Fg7csQ5x7JKG7gOm9hduAdGSQ+wvoMF+8+BEduTQBF
vJl3ackbYurefaqTpyKVgVCvCc51BJnSLSVQkYWfx3XxN6lwKdSnxbVK6Ne6V3zAGyW+P0m8RN89
+ru53BbXOmEITw4jrIwEshuCSZg/yQmwchbJmUlSmveb303/QqCUOUEhqcvd0RVl6RcIIuxNB2J/
z+dsjJMXuP4qGJXUQ3Wz9idW5y4i5mrxCox6uuJFxGrlna6BpF31EmMlTedQMtk3zfWFK3VoHaG+
lKRDx3zrSzlZ+Sqb5B2/e0ZbWcwKzVggMCb7X8febDWX2LrgE7zCiSVIMQhnHgDSCxOLnkyWr1gx
PSGPFmkmg2bL2kVe6GS7VGE8RHlL4xRer9/VZYCBJPwUKbHjLtt9qc2eVFS4Ww/8kv+6Mt8PtgyO
bJOYWxqPYLGHZcFlLR3jVW7yVn9m3ZKhgDR60gnmG/0thg76eJ7NTc9t0hjyKP+s68QinGbJwkFc
Grz6rnMsdE8K+nyXqxUQpnuHx08k66ypCWH2/fxw6I3SR5nUXqXLCdwOYUyNS1QfcL8nTT9d/7EY
pj3Z79ujDQjQEPvESZ3xOR8n9IJf8B86x6yKR4Wp6GHpD7iCTkbuuuwLnR6CnmG5DdQPiAkrgDQQ
BFf2dWtX2+LkHC90p6UB9KxzQQEgj4bpTZU+fgHMt5JN4r3IcbgqR4Ru88uPcTbOVqdAivkbanCX
VC6QPZTc2VXyGHpwIbcFGfyxVxZM4j+Qrn6C7l+R74amyI8VqCRbVaqCNVspE8rycXw8A4mHCFm0
UcS36Scrn4fED8+KAXgeohKN2xdKrRlVw6z4vO9rxqRTsSqKi6wHp19VfINnpkB18v90GfbdvUtZ
T4N58FXVimi2t5JwHKGcgb6QQFahre6615lXw/yJ1hsym6MUBf91u5mIfid6vGYXnNZzu4V5Fl0p
+s/jTNYz9/ecBMEJIekVuvKjwdFGwIZBdcNFzhi8/6vE03QSysTUN+8MmoVyH/OTCTBbEovXAshg
DIhCSD+jAgxAHMSa/YDMe+8g2SpP2+SmbdrHL1HA+w6UCRgk5vtPHKDi5WwFJuBO18Wyj6N17PH8
Zt6fx5/yCJvqV47PhAbyXX0MsM8PLVr6RDSkfnQRPj+B7QYfogkMY7XdrquFc2nhFIRPORTmMLCY
Cuk+VRsuCGA4ss+eZLcNwmuG8tTB9illdL6fxESjim20jfRsbRpp2pNxAo45mv+pGGekyke5PmX8
nMRBRsN6Jk83VIjF+w9aqrf7DEGiwH0euU1omFIf2qL147hmYmEklTZN31HDxXkmt9oXQZABg/ip
K3Al4uO1WzHC5n06IzouHsfMKm+7O9ETlD9gLQmwf619bfQ9TXhQLQnBLjI4DWoGTU5qrY5YHv0V
7Oju3/0geyqzdYq1BIdAfmvAatRS/yk7eTxDYGeKMzGBWxzQvurMWk28XAMn6HjPL5RClHtRkh2E
cX7sSBOBFz6VacEQ98EfV8Pus0k1jUw3Vj3sTrfrola5GX2iHiw0K3OcE3wgQ7JnXnF5J57yburI
feeiCzcS0lUqdRLvJ2WoULAz7rNk6UjnzrIUOFjfaeHAEmOq+eckPhqrmOj54Du+Cq9IxWzraSp5
jfPugPyas5QZYH96koTR+2s2rsANLI1hhvbXOLDAI7ItykYN0eeqJuXRSI7KTR7i8WLnMq+3QE70
7iS6Krs8aSuh9W4yLreNZsmuJPL/VAae7Lp1ZPvn79q+kjRIgErEsoUUYEhV/8fC8UOXEuQaHP6P
THFFe8oeET2tSm9BRbO+ethLz2AK6TPG005O8Z1UUlFO3tAeB+QBoqvsYG2wDzXhznKfP+T2zujw
2UzgYkTPnRwip/U5pcnTBh1tJSnc3CUKFBUHtM1rf4KefXMatRki35ef3yJUZZR3gKHSrNWHuRDd
vgvuirQrYftQPggrJKuyS1o8xbF1OD/nUCxbd4XPTn5yRpUA/lTYTQSQZT0xzyTxOW80D/4PNHG6
ack+Dp139/2R4aCPJB2oJaNMuZHFPgUL3ySZi01OQlIvG2JECgPP3voXcFGIwJ2QSSlhVN2QFU/0
BjxCjbhyBXNnwfJxQLsiCuqHaQ3+MmC6KFgsxR3xneg3JUe+FDQTmoQhltrUHHkRARKEZeZml2gX
PtPq3/v7ScCk/DWyLsisZh/K2itlr4e/bXW+WZEFEm28e07ETqARrFxpur2Hn7EJ+AakSDQw30gs
CUmQHjujOnndZ/4B33d1HDZw8/ygxrGcN9HlkF7/qatfJW3cPyB+DkQEwOkQz1WJo5BUKmbb39hS
HdO7iIOMyCzu0TPGQmB+jFVwBuvs1XphZJChFldn9UU8X8HinYFDk05GtvRtc+0knXqhNSanmZzk
AGr/8O+Y/eQ7mWRP7AE9bes/iZaZXSzuwysvS8i0NY0eSC952VnBQg73q4Z6hHWlYIKBlRo1geoe
M81FEqdrNrQEHPk35tjbfAVUo2mT2IQ3S5Xlu2J3WPxI7HtwLsX3yhv17IN7SIwaskBjbg7QBWlF
5Fm0rjSC0qjPWlR9wC7QYWkA6S+OyGp8n1kuJTOs65jTBVwXSFOHSgc4nJFG+BHP3zsvHKrcgPuA
Tnohb7ZOAfYCq2DTUdxTT3b/Ns4kgJSjd8deXzwiV0NYALlL76Qo6kAd/K6guP8hRlAQy9zaqJdV
lH6ZaKXqhQnQFEgH5mzJMR5h1zah67l3vJgnl26U5+v4Idr9Mss4ChXvvIIXrB7cRLszMxEajR09
QkNZfs1SsJJjJuHu/5p8F73f91Lj4WhSR8059epcO5KokUInQ4BGyxk+SHArANxtthv8pDSs39uQ
aFzy6Fj8iJHOAXrn7f2dbV2tySso4Ypq0SRm0Xse9bodOQ/EcGmcAk/Yr+6LQH83umRIwONPCsQs
ODt2ZWRh1NB4+nzJ3NSveDBzGwd7ynWHWlEqj96D+NUxJ3NjPnaKO/UwwrTgna5KzePCiRznY+ri
6aPJCdbFjj+ijILmh25xaUi/6XgH41F+wD9pNwB6rHOMisLV4Hg75dOR55uDfZ4uFBBCEurH0e+m
02pgO79tTuouXVFiodiuwt9Q1LRYlQueGpxWvcXhYvXP38A/86CveP5M/FH8paLxbJt/ZgaN3A1a
tcHgrQwfsKdlBqXlQcLGmjXro+CONgcuVqFci0SUS4CQWUKc3Ky5yTIiZH9TG+JSAzrFP+h2IoL8
Q0TBAS3L1h9XW5jdRhQvMLWPdrOT6RZdCiSl6JWjWOycawZSDrmFicEXYAjeZoJ4u1TYEMm+tbS+
QCo40kN0LC7asxaojZaLr5Vi2oCNiYHj+d16ReYIdgz2/3vGuUcFW+Qt4cIPdKKcKMMqVNIU6adt
eOqbs9ATvjrWDvqoO1I8hpMQpC6qpr8hcxehoYpYEyQLMTsjAiSNKcXUX48jGnowleNJfYPgLnHK
8wYR/KHPV6zPHvFjnRjg4DMk0y2VSWbHiACTASVQcMkrNZrLAVvzM3DT7QmcBJIoEjXGCpj87jPH
zCbIhgl+zeeMZqzgk1LGcJhXDinDpL/OdIfjodREJ4EBHT+72OpBype6Otil3RL+MxO2jL/Ruq/u
TazSNpLamE4LIy49UdPx6qNqsufNfITPm8udX9gYTBXLBpq4ph3uPpx2eZe2H7b6x/xAXApwZfd7
txjDO23/tx1QTpXeUjG0C4pOZ2BPj2Oxrb266cqJ3Jz/PimvjUAAWPijQ/sS00byyWc1ZJ6J3FEv
fDWPxWyrakT6zZCL3QFtMOGDm4a/knT9bIXcShxrWTNKL9dDFKFAiG/UgBphIcmnts3WY/8+bF+F
dJ6ozvcvliJHV2GZqROwRzEbTDkH7lT1Wu7PnDq32XrP/hL9VdY/ipoYvE5hE24I7KEBzcDimQ5G
NYs907cdyFEl+KMHT0/BiW2Wrf+eZ1HocHx2o1eUsZQe+yPCrAYxXiSgDWYVxSzE4eCIFmpn2wTR
nixLqCZyPqsuXY1s0FCsorGcBi6i4TJ2TBwTI958quGIWP4xlfivs95ReC7OvQ0+0ocwoLS1w6nP
XSgegny/CQqd44msP6Oz1i5WpF4PhGBtlZ+mb5bjX8ck4//LHqKPhiMvr2d0Fv0dUUOp4OAZfgkP
SLTIKOxO/3UL0GrsT8Thgy8wf+4oldtY3Y6ZoOdqO+spNR2rj4n2fIEq3YJA6uum6l9A36vvnY8+
6L7y7jdG6JgCvuShrS+qRdPSjzg+Rifc3tMz4mSY0lc/R/RP2Xz/FGzVny3qq07Wzuk1NtJaQDPp
1LOwrAfy+oZFwhZwQmp68QD75FBqD/ma14EwdROhRzQm0k4Orwp5OTDPCqlsOI0q0PEZ/VKDnFb8
mmY5/4d4XmPjCfqUfeFCADxjrAugRHApyunwVmbk7mPNFr/DifkRn6OUxJJljc05CkptZ+4biUQ9
02vT+//w0Rmd4VnWcsAynFVwLFJmgybGnDhXWMWRrNhnMrxa7qCB0UpJcEOFbm6jCD6eUMKTCarD
C/89jxsr0WNOF4DOjleyW+zFJ6BXCoghmFYlE9PHMJV4OIOZ/kmEtEcDDQE7kfcR6sG7BkJg8sbN
s1P1a993hzLzP88F8BrxkQOuRaGvjjrFMlWwVoLj7941jsIkHG46bj3SYxtxCtiSuOqcO9+H7xRH
3D21f+Onsso87NzFPn4Fb7L0PABlMGtzENBCbqxy1f9dg0lSGdVzi/8N9CJZ+lT3ZqZDRJlGF0Ss
H92kGXVoT9xgxioQvKkDva36L9Ob0O/7+zj77V6aO29biwyHVzjb3O3/8FDW2CuAhg3q79bLTzc8
2yKDjFeKYsGwrsjRlrFVPRa3UsJkJ72lWm22Lv47WGQJmriQ3ujgVA45sN8XQIaZKBA0bF0UKcG/
3lM07qGyDtoL2XikBD26wUetjy/qAozG+x8udQ/evRgz9lDkU4DO+kXbD0tWCPKfUmPY8unJeYNA
DYhW/+4rveuUImNHuVcQRY8v5wY9nXekCVDkIvCSgpB2ivYb5JC8pj8CVdBmpuVp5ovc4ZIkI21c
IY8FIcLz5yVM4BztQ9ku9CMFX0/N06HHUNfhLNhusAvkR76oNBVTx3CFjIagNjYhchDRIwd+aSF9
7c3hmzy3XynaT7/mxMgjvvkBfEEPAOpewQCJrS6EXNSNDo6LUAoQUMrJZCH8v8jbidbupmffRR4L
FkYUIFIPOf8eAX+z5g9XOn/g5pI/1AqKaeSPalb35gPFI4NHztbIDl5o+XvSBwmuBs+3EAFjq4SP
2FuTroqHRi2AcadFqLRqsfkLKUGOhVz4N05brwu1bDQhSqsqw0ERtgqCmA1+wY62Jp5pVUH2LnYS
IG3XgC66cKcK9AaMYPugcEhi7IDo1cV8w6IXzgyaemX9N9vwUVGIgaI44+FWWaKHBebr3EXygEv5
isjtUZ5T6NxzaySofS07g1IIcgrbNnAVWuwJ5o5K8YR3fqf8B62UFGokue/gDh2CoY/Id/HZQ/xP
nhhGq07dAbCSXWPkGSE437NWRtBg8uH2Ga1JJfia1xY8bO3PKhwEkF9xlPkj8Us68Hk7yOfUBvt0
/TnsUEmjGu8g/2GVuqD7G9xn1kWulvjfcHRIq/SQq+Ggy1sW1tcX/wB3gS3VE98mWkaxphYi2if4
/WmtLz0Tkg/KVtptC3lBcir401wt5sZpmac+z0fHqmSvZksRfST1oLjX+/sbu0Et6RSEHf8LQCiX
ASgbfg142yz9W3W3O9W8OJUawtOib9xa8/TrplzmlY9i4uHUQAIMMKWqSLazMnzSWUYRmtOOuAW7
L+y9sHouzfJDWELAG4kyOm4h/U296dIhaTNKQrKyotTHDe525jp69idUuEtzFVFlMsFGHOvqdnDR
BNA6QaqtNnScFOGNcxLAzH2n3dV0qgRL6gP8fvSRvXJVh8hRnjDAgq5+K9aklrM9oDKaRyr/N9C9
A+4Yp7sC+ASzQcMKBbMHyrDis0EHsGd4nSa8gl7XRlOW+iK7XV18DZnKQ4Si5yZt+vTUdER51RcW
lSOeU5VE2BUcr5gSr9TwWDwVRE/89t12F8CpjXsCxFrX8ZPcOUdcg2MGCTrvkOSkvT1iEkDRkPjr
ihs6fIHv5hRLmho6nOppGPQ3lsjoQTl7aNQdK/rEmns98TJOM4M9nYrh0/WIDWMPmyVJmxlwIfQh
uFauG8V2SF5ZsfMoZdBqUlTVNcPSIR7Eu5ojo+T38990ccAM1Khq9c0jPPi5V16lDkIX5EW44O/G
XrzBa+LiqrNSqKC3Hx8WR2NCik4+bTYQrKWMIHcvyCUlfxman5ZGkbfZFsOgsoonpGMb6YG4ypRh
JE2ZtTAfNGqLadWYyfBpWuPWckUaA/cVcv7yaVQ1hYOqSg7wo64SYlCtJUu37FZm75bnXHOaPTCk
80pmNLfXmGhZ4FAjhjMbf+TtcB2x68jGoxYwIIrLdgifJ9M5yDQixIHE8SAQmsIFTnEa2sTDh/to
+C8fZigchA52KZMY8iYpf0NFceX2ZZHnFIK1vQb3Sr9UmUHtImFfztchnAW+xrLFXM7uJOeKtwM2
KMFeX3xZyXQfIDClllW7VISmrHTZTuDnnZDBgqMwjdEUOEepplbPkKgsLOceo9AtgUvTMDfF/KPl
c+vj0p/AmaaJK0oH1EZChKOM5/RFUxKrcxR6eY7Q0IqKLImkAcn7pPl4scnnZbDUtgXav9cNCsEo
2U4hnsgKQckKtH97B0S9+THk+tK3IJaY2u+WpZW8TDwzImlCaRl0gzVXtdoIBXr03TyXC6MaR1eW
gV3egBVL2dFgrWEzTiexb/QEEeftx7oKJXn2TuIWI2i/gVB8Ct3GLZchDCvUkjFd6j0jOM403t2X
kv/WQIhM1YweBKtwHLpne108D8hk1pYJm06k9jMwbiV188p8hM06FJBW3WcNoadpvlXj8erCk4Fq
J3dXQ5vixvxIxRKFmDYzdNsyupp9Kkgji+xKrAG8lS7SpfbuKqE1K+AdZtkC46YbJkoBtr5x7OLX
CzLdSbhEgDcXgKI0mDCj5HEtLjCVRG4Ds7nsheDqdymLJmKkorDtaXSaTPxTCU2zxwup/E5mZ7NM
TfTXQUm1FkLEXt891jGUhs/gUIROpIEx9dTX1w5fistCOurzFZiJRc3g/+ELTjo75VCUoTnEV7wm
j+w70tklpNDpWA+H9skztnetL0zRHzqO4v5U4g9uujXuFmratkVFu4RCnlVUO77xifM6EYmgFnhv
4OOTmeK4657raiOab5Up8Qzm7qB1dMF7uEWckR0iowAEvMN2lII+pzGotk0eHVTrLqo/uuULV9Ou
Jl+UFL4NlgUvcTSRlD4APMTwGWMBL69tneIa7sMMzg+h0FwxonomQxftevfY+6SueW6hcaK1UzS8
6U0S9COXQUcjo22mU3lIjeVZjhv1Z5zxPQ78mZlT5ohBSq0fw04HiujbspXhd3siSLcitGfD53fN
9TNev9zhI/BLZmrbqlC3VTnWv8SWf6nswpVrvZQeBSVvt3tLDlh1f2GtR+hC5SQJyFPiw8mySXCr
NjeUs0riUx2Rtz100+4zx+pVmV7oS1VvMfCh6QUDklSPC+aowXdPtk1Y8DGYoSvxwPULeQl9zDxM
fvTJ0wQ8E3VichbfkT4VqVFEyROGHd1tY21Y0K48w6Sy6sTrELPF3pAO4VdHS7O3UeuUFYYaQ2uP
JageNYQ24I6tb1Gcrbu7tyJDywuIzZVcV7Welli9zLoxJZSliuiUEFVv3HQnwqanMqG14oPuNpMc
x6ZKpLuKvvsEJ48L74hH0p/zYgi69CsfY7N4gltoFqmzrXooNeRLPfF08r+NK02nyqnPFGM2MWpx
kk6GaBwc0VD+G/id/M6d4oKnTxykHdljPx90PCbTzQmdEktsJgIq/VkYS8dAzlOh85CKmHHCY/yD
L3URZyJ9El2e3jBmOlM4jyrcqB5/vUc5eMkqdYgo3SVZDXpr2O498AsGoRoc+ExKy6aQNB7ZvwJI
Yh5qxkjmkXFLh1ey7aZ0c4zWcAydnoJxl0wHcGMDh+TfCel0zynfJfEMYq1Wu4JoOKD+2ArpjUxn
mWbo2iaqQiKogWfqcuktzQJpYTwrWMRAlr2tmF7a3yTGYkOMuB18fqTp4sYT5ONhu+rqPUXHwJBQ
TFRD6oPztdAtnbH4TDfLWHJ8VkLWn7B0yuH/WnX/+Bq7r0AtYoHCiOZyHqACJMwRN835QrfTt3sT
84tITuj+b9nj70t5vZIN6+1p6YXqbJO95CAafJcNe05dfpLlwzxlWvkP2sY+cG5qbV95duRjm7Th
Mc8P3N7rX4JV/Fw5qg/TChO5ZOluyxq6XlpLuWGPzBO7B4q1HuSNNTZjVA9oBjjSzRlY+1POq0We
hlX5w+vdEBPA+vmbNKgdIRCIYtT3UWRX+fvo/j1COV11FJ4Mty8xf6LmtFK2LxA4oKYHOi1cLHIH
PvK5r4poj1KYlKurMaZ0nwJ/ydrkAAmuCjq8ScEk/Jr6dC/atepyk1iWQ5UbTDSrE/nIjMbzBxhX
kPMkJumlSZCCnoaEdgBPwcnDI57lhky/bd6jS3di2yR8Vz/dnf2VJlvysb8zU4wbJTbe7A5Igfzx
2TaI3QmanQHEjova+peuKbLrbpBoatSzI2wa9Z7qIEDNd0SpGmthU2SGbTf6jUc+dPyCqotsYeF+
i5VzEIoUmRL9c7n1DgC9GUWX53+lmeTm6aX3FjoNKzhc1e3905+curk0qlJWfkq+tSt1AdEYZOpr
HmTB2tAZTQDq/IAA3zB7YwdPoF0df8Ls+wVnB8Og6guHRNNfCoLWcejzN/0FgLchbS7bDMvVcDDH
F88MQsMy8W5tXRV/MLPF3yhL0PKqcUCORmCZ+CnKdkhk5QtM1PmT58c5G3oSc4n6kTU8T1h1HlQi
1JJQbaj1NbEkzOiwRqkB4YWy26Sm0QA/mO2Dd4C9ECYMwv9oNWINk7etW3K14Ftw690OVeHDhvNO
Z4GDfirsIiLcCfa/iM9vlxmDP+A0EHuY3+gr3Ji5BXZ9glELxQBwb3ip5L3VzD5Ney1YZ5MExumY
EvHqgz04ePHcgMTYO3i9zxPvvzvKO3tNCZf0htVmrXvcC6mpxgpz9tCeBQPCN7UNqPeFigUwzTL9
1uZrx9yG8QxiKx2mwssT6G3gYe8VRaQht74o/OaqdnF5fHt9MqcLmVbyeXBott9A/ecMuQRnw5AE
WEjrvuZ9xDorT0GlfUgsFWUr2AiedpOiahAq8U2ggLQd0jdaROV6W9ZFNK4SVvA/uHLEmB6jXwfX
BpCQDWttrD44ZZAvqzdGFYH3JlZ2G4jJYEUul2yIUnyX1yFhBS8SSIiwttIGbO+JgxTxI7L/VVu3
BHI1BecWmUM23RbvS5atK8RfALJXuUlnmAJPss1HK4gAkkr3cHWyarWXuNiMcK6AI+QtbH0jj1U8
ls4xOMVMg2ZhW+Yqs5WNcAn1eFmMgXgNxvRlpawFhVDE/IaYFQU+SY2Gtb0ExsAcAS7MNRD63TV0
sWDfSxvLrskRzJpTH8qKKZOcwA8R18Q8MLWHFtznlLdbYjTwDp3fVm1+GjGTHpZ51eWF6u6a2yPN
swwVCvs/gmWhjKcwfEy1PFIa0kjdeEc/PQxDV3EicJmc11KnFJAF7AeQRszH76A9iXBfbssNXuhM
l4X//548PcExMuozH+y4d0rjJ4fT9sZifyQaLdk/dzS+U21viGIbtVtxlyqs5zFxwSpFwiQsIdUo
9kgmot9L88CzucOq/IHHj3SfugHtYAzBwH+7Gyyi2G0+oW5n09/b18+n4Mc22fnt3gylqcGukvXb
3U8+0hVs1kH2Mt0ZwtAfyAnmiBIT6Pz31ulfYRkWUmhjq3kleYx5GgQ6ROzF1JZAZx5o5x/42TM7
hUY//N/8eRJZtU7b0MapdOXJ6YbYEAcO/doCiT9QY1MJEsbtA0hs7r/OdzQepEX1oi1VOpmJMOha
KRQ4Q7s9+aNya/Zd5Z3UjRVe06X7hUDmB4CokgpeIYewDUHWNN0f4Ao7JrkigNFFWDJWH0zfGn/B
BiQ1XGXEiD8EDHueFRgqnYoBGtRUNYt3WwiWgJqSmaXzp8NW2syxyrqmzf4E7YM45Phd8TcjMib1
hx2Droax365hncY5rXKUSckGP+JUWw6U0wOOOVePGU0hKprdHX/4wv4FECUrhWs4+nlZzkQPa31q
6PJqTuFa9NGXSIRh/MbHLMGrjJifEed0v0sWYaxYOspfHxm43S412z/lfoeou3YOWRc3xWql8vK9
fsX+D559R2oQE5WhvZTwhMvXAh15oPzkBctfWnIOJ8RjZGs0tYDFDDzsp2XbI2597FEwaVhisqU6
TJ0JwIDMEDkiY0R9OkTpSgRc99+/JutwtpmhJB5CI/++amQUJD3R4bx2uBRU+R/0gfi/sV+4dscv
CrxFepJssbsm0ILEqHl/FOCY/X4zpv7aDRzrMcyX6ri01reUcgP1rj162LLkxUM1Pke9EPvuuhSg
Kd41nAF164reKJ5VAUYHsc5Kzf394d8tGxASI9cpqK2yodh/QCRQZ7aMgpalo9AT0iyVzPXHboz8
2k8rmRYFhdD0eAaVdN5vVqxhAXt1AKKEk/PeSKcX6A8uGW37i9CMS7p4qrdpnEGj/j6sjYwtNdUB
Twt4+Wmo3ABbma5hIzEeqi2KjrHItyOpwofOsm48ZA1wGMgiE/3PNZi8uZt8IYv4ywYLLjly4RZc
1kTZ6oAKnBnxXEgv9Pnl9hLuVOv6xrJQc2cO+0vutGOCpBZgTDEoZzeKer5ImiRNtUC3CxLuaDyl
5M190ArX6lfVCRdQn6gCBAwLhqQvKTjJKpngEIHusANOEwVBD9vACGm/dqMnFOwLdusTWA1uH54q
F+wFrI5xgDefaubcF2exTB08wnhPp1SJkBHaaV7Vy1+32SIMLVIKR/b6/XpoCF8GY0xK/KFdtIoh
epFyClRn58h2bGeHLMkyGfqRkLUWgN1FHbsBlexrGv69wN/M8XWR91EfU3uC7k0a+4pLsxNsiVtz
6Jo7aO9gxD5Vc5Rywm94rAeCJJlNZMrc0a4aR7NIFrpF89LfTKWbJur2zA+Y3wV7+6vGuu5xQCrk
kwQXHcoMcrRlNu6w4IIqMF/H8VcQRulLFvaVbZzzgTAV6WQ99HJ+vCvk0LHwsSNbSEcZ6ui5mgSV
MNQNUGKRsBitCZZCu9bAL2sTcZnA58v76ABuZvOPkAhC6d52GSCvUSISEu4LWg77X/CUOXHoIYpe
Rkr8BnG6LtBLiOXqf10dIK/mBTdyw/NXgxQRV4aAA3dVwB//nx2qHJuOpuNyN0o8QQ1PWOHuUkEs
7PLgw4vpzIMJsgF8Jrz8yMiTmhNlu1wX2GXZNW8G7WmV4B0tKnLgRcAHQBNLDyUbGBVTDVsm06nH
2TDhW4JuXXyDIugognoEAkHLtWRJKZTDHmPUrNjx7TV1LjOCpErAzk2+YmgBp47SDuhCX/CMkGUu
kQOAZ9aMjhu5OE3E36fn13oqE6JQUFfRvzcsYdV3A/FP7dRTQDhjXVQCk1aybyeqilDMJwMXK79H
vzfkRKKblXauwtm+zUNdbU9z9m3V+yMwFsbGVLZ2lKdq6TmgTWKTfakxVWW1aD3nFYpraIMSclah
JLIB2X26jpqDz6g9Y25pwM/smZ/5ODef8WFmH37UAS3jQXIGCdpf39X3mI01CN2UyCiEMuaK1pvA
EleVbLRfoL6M/sQzBQ6jbXADv2fq4ODb1zH7GA4MtgcOfeDpEgGEKqTZhrEV7WOOkr8qnkW5ve5Z
KRPd/46z/gvTSMBZ3t9P+DDt17toZHrjthGFsWcKvleCgvzy8/pGaiymSinONMLHwXHmDVyHQt7j
HuXISVdWYObLKhu5U71qCftvKecQ2tIRg4SaeJ39jQWK1Or5cXpq8+kw5SMe+RxlPkth9Q36dVPI
9JCZnuFF5WtQqvtHj3j1rvSQ/WymAmDilfg5F5DgB2213hjkyirzbihF51AcGYkAtFmx8p0iZyhY
jwHItll2D1lMRA4e0/KlXkccqBy1N5IpjxFhMdCSc5INpM6TAy1ocEYyQPjvPrgyUKPi4vfH+Xu2
RjPw6Irw8bxQaoAnPXfV2L39Rm+CAYYbi54ojn7xoSSKpRtFyK+n1VqA9n2zUFHw02nqZxqmQan6
PCctUVUzbvIWFpjs3H/LGpEURzpUrREcmZUWjkcNcj6nOQw9JtBudVRwy3koqLJm6MTjI1VY3r/U
vJ8NFM/zB9bBCLdbRatN8jaAPqvRFhcvB6ABvP0Rd1Bksd1jZyRs/QOx296Q9TyyJmxAdU04aJMy
TIMeIWtw8qP6fl38XUPqHKk7LnpsDOhwTG3qjioV5ExQaXCTkxYtcjvvjpJMHcKvpPVPCqLJlYiy
tAdxGZtiPYbpL0GZiaCovOSw8bo8HWhEyYgJP+ZCKTcy4Kk82GvVVhtINjWIYEOqkKW3W6WAWj4X
jWwBTxBBkhYXBVurKw+py11UoUja/PlwbrW1MesjwB1f2otgVD7ayAbhga70JgGbw7rihsFoM3x1
8SkMeDwtkCuDgkmt27RrCKIFalA0VB8rwBlqFesMegx497gbtnCjgA7WWlujX9IBuIVoR8kqSkcR
r+oTGehKX7hvPyuXT7JVZfot/fyvSRgqjZmxBTvZ2XiIEN1hQkCxbAH/GtW+y184B6ftyxtHzLha
LYV/hvhbtjBMRFsW54JHKoSk+OIxG90s7zxG4wsVhgSPISIgVnn5K5PnyW/iWcrYoruHaaVwcYYq
YFdI85PSOeMTf9FtgQpCzVepkJO2l6KYN3SGQFsUHj0dJlCYPj6Tx8K1sK4N6IPJwLzZNa5Xnkqk
y3lNyLY5B0AmVehIDhf5mH7iQzYtxMeiQx+XQ3Vtoe4n47hLff/goS4EecPS/J/wHJhdYm+DOv5q
V4ZcGzy5TcWo0FkHqr4TOLzZ6PK4xbfRFfjIz1gi5QWUlh4BrMZx3BUAJK23P49k2SVIQ5XqkDbE
8ed+IxZq27TJJ5mcD8C/iLSEuad3L9YSWuSNRKykHD6OIA3h0xHNCwpX82CmWhcxVAgBvNNgqV81
vrvDJ7nxgPE9SaCFtucRcgSRtGwQYvPyo+D0ubqsQyBWtEBQF3fo8LVO1IWXrv6OG2DGdgNaWXO+
fZG7M4H6w/kS7HlxMFB9uppoJG3SmbzSzXsvAryCLL+RIbJAMdWFfU/eIxvC5hpR9445w40SMNdl
4kEBkLWqSIVWNBYovM3esaAcd8LBwe5jCI731Xj1nLFkTUw8Zx0OpWT4kAFwVTw1cfjL12ubJvCH
SMjvuHSIp4IQcTqf1102Oby3D54EqemFamLfBnV5GzM0O7dSmtG5jzQutfl30EnIIm+25inNGgLb
oFWhq8Oo+psxbryx9ZdLDygBrSlWir0Dj0glaxwHafLDuiLGivZS5NdKlZnRrAIQ3yGutaEBC6hc
TRis1+6Brl4F3TI7VRBJNz3LCIGQ2NBIfuO2RnfFGKz5YYhpC8AbqDqn/MgTjaF96lfKKfPmDBRh
GBTRBC1DWlyM8OutpcJYX3RGZ2zZYiCNTjNkp0j3vwK7YXySXp4wYlqakjOv1KOXNHnUFh3U+QT4
W0nLyOCE9hGbmGycYPK2ojoqPPN7cCJCrqecA4zrnWMiptaS88VJu5yZvxRlNUz5Z59BFMGLHP4G
VbtX+ZgOzmgB+oWH+GABZ9lw8nFJ5HPr1mcOPmoBzgdWlrmMaorTQ8WfWQlNJSCNaDzHyqj9r+e5
mwPAtg1cxra+C/B/Z3sLlUlvTA7yey8sIJfhmWc04afaciK/WzGmoq+5sRxjXU9hzjYsNd0Dvh4/
Brrz/wO7Di2d1mtG8StNf8mVYskmxKcFTBWCi2njMbwKENgTr5P44O81ciKm7ZGnvMYhCbClf4gH
JgCMocCUHMIC8p8IcFy9rbOC5EdzSHL7oGljZkEhH9AYnX2sxXoFLMUjPo5oiykobBVbAcbwYsiJ
LNgRYkVxPz++O5a7HfivA/VUwd1Uq8FmOpsdF3UxG7xYLdZj6+8OIlpJct6/AvQVHjO7qYcR3VQn
m8TIM0gl7oLBfiMnb7l0CASagDTQvkLmU+nGo/PSUpD8iAUl4sgfP42WUKiO0qRmwuWAUf1ydb7Q
m4Qx7DDsT+ZEhH6I4yriLY1f1cTKZdHD2BeR+RzkoAiv0eVvFPk7sZZ1sPiGnhirteXO5VqXi3cx
8AMZ/MWGPoAhjg/LqXILHfW1UYI6SQTYpAE3qIwz2JvyLtkHd5VohDVeQjQD2OuUctlUtA6Jqxru
q/Zz8rt/9jhWFPOTkM3FZz91c2kDOKhNmkqTd/sOXMHtNkpHTOm7QArDZyX5CC1advhnbcfheAYa
xkAxL7giTgQcNrKRxzeaPUqLY//dZ7X5/46WN2lq+kY/kN6TszVn/VfcS7dzmkwbfxDmYyn8lVi2
w/RtkJTYIdhfhkifJsLwNjJy/9Ce9yBdIcALQnqKvcV7rO7S+cr/3lqr5pDpKI9M+PlVvqEKxtdw
wyflYR1eH0WV7FH5+Dc4thO456bMI8aLK7Pd6U6E13xuvNQTDz6iHqWIU1tXX2hB+Qlnr9nKVyci
ryNJCB5i4QkJLpH+xTJa7Q6Y2oe4VBajDCzB6Zj+F5y5aKPW5q8cOJkdJAcg2A8ksVM5xD8gewLu
kUE7GPFos62S1saG0J1/+A130QjJw7Q0Yvp/Fe8PWiMI0eHCAdLyt2iDyug454UftxfGfAPCZI46
6AcdlhS7uOxhC0sdRdtVVt1JpAgpEweFv14i0vSzo3653UWobBAXklzU0tU7C9G3LL9rLp/PD5qG
kkmS1+y6zTKOJLD1cjRWyS7W9J8b36Dmbx8/lk/gtRJQ88kJivy/NnID9ByOyWJBMbO1BXhH2A8d
BmmHO3t3xH6RR6Aqaw5sTWcmMXOaMzt73XixsOBqpJAgbumYoL67ePW1+IvnALZTxf2xrV5cUKeK
R2bDNRDSCv16QtKb04yku+K4sTlIJv/VBztYn58OoCWKVSFBzOWqg7Jzx1HmtCTvWB5AriLhtell
MY5Z46EpJvdZ87zZRWIsfsPSIbgOCHLBJ6N3Qg4HzF0+BuJWDrqvEeX+SdeEyF7Qhfdp0QF39x9J
jJrCF+2vMB57SkqvWGKLBIkema/p1yxWWcST5tlMcXgLjnFUbQOrqrcBFXMRZ7p0pu0q97BsX6Hd
rmlzjOd72Sh7qDjOYfL58Hhk+W38XSxTYntV9eRyXdtz2rjI6OtkTuCsBeUvFNtbvGSe+92u9jLm
QefcBDuTom9mknSkzBmohi9KbXf2nTO3Lw2mWJfYwyYNrIWmuIK2mSwlkpShNCP0Z32UISCVNWn3
cZNraj+69ihnRP5gerMas4+jWPBJs/2wPowEEbhtOjeuiWlCogRl0dkl7EemcIOAy5oIwiJndzWm
cUeZa213k+37ZOQqno9NKbWZnOS0CfnD+lWEZJ85jIRDj/46bfztcOxdJixPJ9eQHQAlXYf/ZOws
YsWTvhiDPz9ftiMmoKg0nUrSTeRxSubqjzZcaJpAdkT3aIQele+nsSGGGU+FVEctPX64038TVOt7
EhgH8ySczir9IL2gblVtpv1rO9ImEbNldRi5CKHRJn70ZqP5SZ7bi04dhyQuTfIArsXRzmfVm0+D
9d0RZXPLoym/eX6wyMszcDeeEopn/Sg5+JETqjSBv53NdLhXTRv7c/2tm9dwxtl0QMTeermEi45i
7F68KKgoknjWgY9PLd3qs+H+DlIQ8Dzghal8OuQ0WsLW2kT1kkCZGgS/H7Y5opIy0h5yLbWMzQn3
pfrL0njTSpEFNRGJ2QKk5G0AEmM+i4QUdzI2rcXB1hSddfcECg1dIJfZVXCa0Ohqz13l4SkvEiKg
wAGW+zXQPoaICaRW5Z+CwaghTBDD5VJeYcSSeSLG9CuxZ0HIxvt0QbfxK5rvMnePbbqXJHY69i+S
R49xY45FkZP7MrKr1bw5h6GvGIbgT2x8rYpJXTvAli5YGRtqoxFFR6Jj4QFSU8WUgiPjiuJ2gLDB
lx7cv9TGwUGIieyKZV1ofA72VF5FpUjM2Uvk3Jm6SsvSlnCnq3J1jwftNsP83Vvt2QFyMOhxovv3
S0zBUuJK8ANzCfVL+aQFz8Gk9wtQ1XZBuBWgNoYUlRJjVK87VUmNnMN/Nhdj2RPWnCKUPNarx76d
awFfqVIUD9U1kmSvX+x2zUfF59zv7RT/duGaht76j46XzMR+RdnaybU7vsm1b13Cu9GdeyWkm+J0
W27pmrB0BqNdcjbDdjlxvxs63b/uh80mdDLIqy60dLsVAlTkCgyd60eyog8IiVP8A/+bO0wsHtCu
iyjzPxMpgNo/CPURp+9h0nhPYHwODQbBVzHIc9r+lFSBf5YIp42oIet6f+Bkf1APRgs29whMLru7
pDgDCOOuDfUqY9xkfqvGPUHU7WTbBAcnby4uzRoAeGgK/AwHRL4WMJNoXmPiA4uKB86i4LZIhAGQ
YE+nVuqxJVy4oigmFrpMmqM16qDPK/bTTSR5eI5R/BY43WZbcbVPkQC3BGV4CBfnda1aM9zuGnvN
wDN0OVBnDObWQTmmzudGgdFmB+sb6Fuq+aFG/vtKp9NqqjPewWovPgMEH7s+/b213q6aztYaBX/i
FgzyulPqzJfND/Yp6SZveFsziIuIK8anOKerdKWFshWdY0LjUdC1MZUp7bMbvTWpFztTc7o2NjXB
5kVZAP+G93xlv3l3xfOR3+jqWf2b3m00FATug6f7kragkgXHp/uPhF4k7x36UnkKHF+0HpEHetBJ
DGzHOjPascPWizsIfjEFVmuOvjmUsX8MtZFgi00IO216WFl2RKJRRyfKWMfwd8g+Y5MC10pQ7QR3
fKkzrV2dy4biwkJESCYeLl5EPYSQHoFXZlr2srS+XPm7LRT2S2jjEJNNtqL8qxZd2kTwXtaeCIWC
McDNJYT+V+XvccBrcbMx0gcFtQ80htCzTv4WS3G+ZXIRHYTFEutXd8tTqdWGg2uTe1Ffpv+J6+yn
WKdz6XbKuZzs7JGjCvdWUkVz+VJUNDnJaAX1+qD+0giCiZMjqQzHh4Wtw1PXtuhTXz32hog2seLP
rNIhmCPjbjbk9NXASr0L4B1LlicGerhEv95nb0OdWnOZsL8Btm9qUaNzlfh9fyB9VZ6rDuuvPHNU
ykEbr/pBxRspjEpGEYb11u0R1/C5RnRenBT5OH25e1F03/17NZENm7bYV3/GHm0r4LM+iozOBTqK
oE4CvIUVt+uiqc3AlGYGy4bSL1HoeFWr+6+wQ3bWr2WDPFyAN/CT/jv4K7qk/YNoIyJd8ry/UU8d
ecogQmRLC2PMxzSy5k2UA5jpvX6gfg5ZLgomRcmvZLr3fp3l23iecAbB9lJ5VBmMxsOi5XQCTXOb
2YXs5c24iIpLO1NqlGuSH5XZAYuPoO3wzkGz0ZAurzz/cjZxU0Iu41Yo2m8vWQXnkqfgkSNC2tvT
Kli/PSrbFDNDtQ8kBGdjzZDROoxMizY9mWBxpn0BDEH2aKqsdC+d2ChVn71blEQNvt1+d1y7fiDF
4NCC74iqCs4k1CZ10MPzGhTiMc9/Simuafivvnu0d4bPwZGlOSV7fjuGelzoTFYOkdLdMGPkKNWy
rk2bD6+ViYzy0y9vLIs0H6s4HA70OjMI3+AP4aMQSYyC6He6lCLus0vdxndwM7ku98AGh4kVtI+Q
jHU+b3BRyfUjDG1IhksAKK1wJGu2svXCmq6LPeouCMo/08/e+aImEzRzk9D4n9kcI0crafMqKnBi
FKEw2yOuhGcXGL1ERx1bBTuRa9eJZ+cH23W7xIK3G5h3KSUuhSxr0nuH/+yy+/kQFfYqmGe2rhoz
bi5na+wmT3GNugU+YWdx9gOW5bbqH/OcgXOpVNxc2Q4B1Bgk+91xHfMn7hr7f0Lu+mMnssczymvw
lynSuix59aWzm92C6/j0Kj95Fv6hRXnbm4sUE0LCFJlgh7PBN/NqAJ+KWXyZGHM9Fyft+93oqxoI
SOk989bUOj7zyTT0vTXcIrg+YvhZB2WZgqsRnIG5Rg2gaumrt4P49EtoBwtruyF1XYIZxJScJ8Xn
fqgNJ902WpzwqOu9M0BsNGTw9H6M0GL6gNjtfnLa/3Q5/8DQQGXE0vE2Y5MgFkOEgp6a2y8L6iXQ
WFhXlWMMzMypksoXIXRGIJqipL4Ymwk1raEHcV2o5Lp58HHbWUtNX411lY9ga8SV1PiYrULYGTFV
KeLcTEw3C9gxSZ+bbGvpyq6Ai71zOcBFTTSf0Su+jNOWGPpv4fJgVq+swlTVAsy2EOJ7felbVH0R
7k5bH2Oohb/UTUfKq9GIx/xzXgpRGjNdlnsKopUhBVooNMcL/7TP/95/7BQo3z9ukBW5UiQvu6J1
HGvI/axQFYWrSjQGhBU6wFRNbwF1WfEghe1cJyyVUD0VcNehwJH6HHGV4ywTSU10M2fW9pt3/K1O
nkIpo9R02CwysVrYvpFejKCFhtMxkXeHsyWveJgs0xVYsP9SQ7U76qZinIxUK/Uybhu0kwNyCGDf
8gqbx+9rC7a2lJ0Jf4sPuVQv272S3OheyaKgYTceB889egaDNIhpMp/kBKIaCFtC8QvK+V0SCgVB
6PnzvISyysY6K8b6iCDlhQwyEPIWZCgZzgzlFavdQqhJeTJIQlcLNnbyCfUD5+pdDebmcDJx3zbE
X3/FoHiItuGr8HeWNjOygUMBIN1ucQbI1f2ECIAB5dUkNSCEFuI5O32tPsLqj6ofiNC1iI+QI4tu
aF+wF7dXsBYvQhmyVguADytQnWxaWuZMlF4LFP3gP2wPXanARmjR2yxGeckrYnZ5LV1o4r5t5OzP
/ok+0nwwn9g029mltXkd9DOVNopWBiuPX9b4jJgAA5rv7wNAyjFd1wdR2zJ0f5HQblkdbFEf6ltf
PvUPCYbHbPipYfZfreQrGTzd1/gVDlGCpyOgZ84qk/skcR5cO3KTwKCbzzzbhzQYBtAP5zYBocZ7
qT3WLpwnGvdOrhwYD6RoLZ3dkJjge5tIxzyQQSPn+Crw0r2WG+IV2LLR7J02BXKOtXTH3WafmlaB
F9QSQXaAV48VmJSxrz0ElEThGTqCxMoDgX4UT/oLiKBR6Ayo8jKL/Qlz4zA8qJiG6wkko7BlwTH4
nhthCe7X5+QB8ryOU/zTQkKum7sfUEwo+oaQRETwkmtEDVsPpvYkR5+ONUMFJs/bLL32G3UHFwGm
niPyPiBJoDWmbnvp2mdLJc9ow/iKaqnKafuJJph9hqM1lIW1r2zE15XeBUXuS+4yQxe+VbPkk+5L
gJJHwCWylKguspzwd96hYKlpcup/9/9SO9cijiokQ/MuLSj3RJS12ZdA68gf/SYXWgcIngc3GFsJ
XvG24IXVNzxz03ejzatMRt0n82qzwUKBlfdE6IuaRieYdnBYjjEEQ4NcNLSi55MDyKLtOQXK1hFX
JtIiEwzEU1lb8BuMgi6rZX39GhnOPwkQN1aeKoaT2InWmehoxyhM4iyyV8bjMpfc3DWSAOb7IiBg
Ns3m+/fbwKLu3WBtsboFtX4SzkEUKiDcbvh7vnP54u0kRHEHHz+xAzyq7ApDPezGUdafxEDpiirq
iq21K2kpXmZD9FDMyHSXjd8fhGTXOlzhVHK/0Ujc9Gm/31ID8XQv00tOjCS+ezlZ+N7ZZQwJ4JHz
iwQrZjBlZk6N8Be5zhHnpAfmIj0t6ox/z7y7iy1jtEFO2zZ60sUOBRtzKUuuW16vmiIsc+5xkY9u
nTtA72InMDX5SgBNy1MdBb8GFOJOmghLJVM1sok1axoSLJcU7+dgf5AWUkp9qkTY1IJLHOYWf/A0
VHBcncLoSucxMfNn69+AA7OF4PQ/LfbsXHnobI+J0+ysHquhBrdFLrtceJAgCo4uNPObW7OlhnzG
haAk3QWw6kuo+cDKze5GTAsNtkgkYHbjAW9/sGphe7V8hdaXq0V7YFG6KTYuJVSAtYVDYi8z+Xgv
+ZeroexTBaOm+2px17RgDuMgJ8dLXWA2BqrZ64DOvXluXZAaOiZXMd+hTm64ldp3qPWhJ2GkOeKW
fHGKNCCJ4AUYFAChHRYOqUksi27muTPGCxDCVMxGheW06BLVaBZvT4U7NsJ9tRE6sXeNfWgWOCJ9
gO2+itUjxzTjrn5MLEv7NQVCX1aoz3oI0RfzTJOsLZwt47FXmpS7ey6v3A73RfbOcp+Xvmf6rB12
WPXfiQcChKThSxF0dzPRzSzCEXsh13j6LDQHnCAoQWK5JosjpLdpi6ck3ahaCOCzSzBETjn6nq4Y
sk93y5LOyjEuolkX79Y07YMZycBlciT1MvdIVg2WWMUaJIZ4pai7D7WbEt5jEAxOo2CGO4Ow2mqt
/SRDMHHAeHm5M8SWf2XQpMmlvYZ+LyCDFyLx/AXEqDKdD/hYroYLiwSuMRt+pSN+ivI//1T+Vr6p
5Ox6EqWKLYJYMZnH15ctJ7FFa8OxyrnHUtR/2eMFaXV7z9wa8Rvuv4mhfTMfDTCITsTODZhOxpFh
7fUAAmWfdbZ7FppgLIBChpOyOO5R5G5yKSzlUBE7mtB1ibNsGnqwgGpobG0rNedaFTIekU3dIlV+
kvbfQvVT3xJbwk6/PohBkZUoQjCUulk7a1Yr76aEvYKMGLKWjyM1nLc+fOBT3IbI/AV27KpmzyOz
WXfLJmya4GN3a0WZ+6TFTirhE/zS7h9RWneBM3LuV6ATqY62mcdw5zRDPBUBSceg2GrGfrXKrzRW
YCaLSXpxRu+Bwin4EDpFPA+I3REek4uMFS7h4kBngmq0LT1pS+PGXSJUsgDRXFbA/QXGAKcsa+0x
l54KsSHoBDubsiPxEGuPUkQ01Tltj7z2cs6c53k/OvvUcV4PoPVY3je0pF5Pl0N9pyt7+XZ6YdGE
RFZpjn9afgULrlaNSf1+C1ZUm+9APGGz7MQouoiKMapi0l5GVCGIYM9LHS61d8Sl/BXzLpIMTvR9
/UG5zRu8vlkyrGO5tnMSTZzxzAF8ePtw/Rt1Q090mhbwqZwV1UWZNWjm8R22QPg1Dryq2f+1693H
kuOdoOSQWbTEKDXDersGa8oSXZn4v/xQ/IP9w75MCSF3eUeuildnAqD4OdQ032VEfiZgs2kAA6f/
81dUXsZNuKdKwNNHgzCuczmSmbiFVNtz4vZjq+sQuKx+w1jhnulxxCEj7jBoE/ESkzM0FAFA1hSV
BBQVj5WYx1E/nyzZT7qr19mIS71+w75HuXHpc5pMsSYfBMT8WqfFXKkwQUGHry/ttqIxUs6j3Mzs
rcez+xVkhJotryukoD1+Oaoz+jHAFo1lp070ksRZWL2up3nEoilhAiku5ulMDaD1MeRQ9scU6K11
nQXRteMOhho2fC1ApFZ7wOFDniAP5MT64X9Nh5krsXkVDT4QtgSmxhLO26CrBxwQTKIXj3gsipfT
kx0Jl8cE6g1n1JVoKk5Q4dpGlKDvFULdMYbGCPmxdt3eOA6SkbuNw9/N4HNJIwaRJq0+7uYNXko9
8aFSg+kxmXBkRS1IlqRVtJtMLx0jKlKOYBY4qKoSm3vYJl93e/sZbU5haotPptCSllzGgAf69OwH
S3NeNDQdaOxfpDb4JmtBNOFwGuqVpKsLxmsLaAW19Le6UBO+4TbQ6S4mDZ7SqrfVEYzdfr912LpN
jvQ8nlJSazzPig6i3scg/0pnnW6htrXUTkWaei62zYxcGglQaELdDtBmBpTNc8Mg9HrOngLTNNgy
fopsr0tEAGCnYhtOhQLJ3o387pYu0OB7+qHDsvh1e8HgjX/ADERhuAmx16tglD4JkK7l6jxEVvcU
es4BF2l4+B5BQe/XJ2Led/y8S/Q7S7cmWP16UZaVe2dr9VYEHosQmJooxghVSDPw8SnZrpPzv56d
he5gqJXdPYboCwib9syOOUXwIBjVU8Hde+QKMPR0NIiWGwVO1q1/PZAGQJITUvD1EIVyEsOQLPKV
x0HQmc77zh/zw4eLQ9DVr6DUJbwc5tJTjkW7X6cSMeNVdgv41ZULZhy/mHEAjZZVi9Q3+j9/Meyy
nAHJucXKx2OPhsu59p+JXYG1PqJBh+S7VmtPQMYIb2zKvfmsQf8W04HuTPCQzDqJrKe4mqZLlKO+
HNZV/EPPx3iKgXti4dSnMuSYg3cMf+d4exEmKf8iT1QXjtqgsxiLcSWa4U2SQxQzZSYicq5MeV5R
RjfPGt8hHky6qcpVB6dBsK3SeMsDtTtqmyN02dcEpHFBNhbGyhJedMDg6v/KcorHz+t2HIv5rMsj
EB2SBix3ybXObDvvBunrOX5PvCKiL3rR69067PVOEr9tPLoH8SjJwSBHLVbrlyPb6TATmgQDDFK1
XH9igfq1dnJvdyE2G1HYquxZFuum1DmnTigkmEaor7RzGYQhoBNsOPS2hpc3h6y3mkZ6Ndje6oXU
z5hSQt2Z8VBqqBxCfg4LdseVFpsznDMmBCzeAwu1DulKl1BHj7wgdP6z4vlSZq29A9M1s70nwJi+
GIcVHRn/nFKLtKoxeKVPjFW64zkG6iBCKbsLNQ6yiu9MfGfdLHCDtjSKdhfyxQ111//maSkgLQDp
rDK8SQrQjS2Qhj6yj0C8ZLAtclJ+amnLNURbco66s8vb/db2Lm/024k0ZgU/ezds4XClOy6GjLN9
6dhHb4W5OoCWC88atT1CHF/8D5r13N474UPD7STcCzmluCkXivYjpjmK7QEtdgUfyjK5BJWPrI7l
xyqHMlEJBX7zv5r15Oarcoysu8tIYB3i6GJlM2eg9pZVEyCpsptJ7xKEVnimI9ZenZySohlo7+EU
GiOAOjJRFTI7vezjxva2zb7pTWARQsYa4h/0bIZL3l+SlP0s4nMadVftjJusFy/z48FhgxfrjCd3
q6s9vn6YmEHQvdEakpLF9kbPI0Fh2LbLgUFrskX2yqYXABYqfoDbT8TBUdqXtm64a79AFWNmjnYA
i0dOU9xveGqhLMiXnFt76oUzrV/qreMuuuY3eBLw5Mu7PhW+PTvSgs1NexZ2EWzvkSloeLqkS7as
MROj7hJbCxmu6gtEalbubmLQdFCPmiWnVf3p1gspqHj9DLlQ9QhLHp+sKqzc2Tsra0goKl1NecU0
IPZBlcVinK1AiL5qlX5ptueAdUIi7fDraViOZsa0SqYz1MDs1XMg/aTSTGxRtyfPt7O5ZB34yms/
MKWzcbQbTUxqAuDmdjkBlL2gCaMvTHT1lQu2rj3lL32c31RL81HQ+IvNmkkWvjvXwN/guZ69sR4l
X3NimMboXX+jAlV7xQUFyKCUeMwmM9s0vkP1tmtysZRWVCrOFI3IcNRUXY1SaluS0wxMN1oclZ2s
TotyO/Ig9hi4kEgle6GpU4Zg03FrVOTRhtSNXIwlwEmD5VLdDoNZ6r40ek8y+IKM0JJo0JpZErFe
dJraqqISrh1Rlo6DdbmBmcnGWXSe15Bks5moLBV8Xf6vzz+8pNzaaz4loUIe2+H0r5wdTiVDjL2+
pNbanCG8PPcm7qCdOwzW7FIFr0j/SHcqyR9xOpKQYB3cjUuCULlPj+J52JWJaM0vDmSRtULbfvUP
wRBoUnJ18ohlvyZk1+iRR1Sl3u3HEwXg3gT6QUOsF2t5hAPlZ1HjErRCu19pMQZwUmbya5oeAfvT
sxKha5OyZ3OH5A9GmFrna5OSpUYql11dX3dnbI4ibHP25oh5p1XeEin75lsDNgec/qe08xgo5Nef
c7conPzXLMM43vHK4Cl/ocjd1N0AuCU/O986Wp+AzeLh4WoofnmMYDJjzz5xju1iI/ZxAzd6hdrE
QBIj/nTe6/5jzoTG07pBIcLSunOmmFr2wvxXGLuU8sM4Ldk3T63DmhHdqz3lAoc8T3bQH9LtlzKG
bC1Yd1jXF4SPaf5qZPk+mzxIK7wdJQsgZiMNw7eNgOM4c/Oi5RWQu3KXTletHRzTUTFTune0/2hn
uTKjNJkOHXczq2QYsLO5WHNiOPSFsQzXeqk5S5CCWC+zT5eIIAfgNzvoWXpsYzqEaef6QIDkZNDE
twSgFOR9ItIeM9KcXV2u7GwbN8hAFhSIdaW0ZyyiD9FeWt8ATpF3djTPiTE7rLMc5Ew/D8lBwYlG
cyu+bYXSCT01PiR4QZR63HxHvLpTJ8ygp5dbPYIbQC19NPR6nY6JrulKNC92pbQAh8Ka+AC4wzpv
86uzZdJv2p6kK8ZT2N6xmoDNmJrAeR+rKGoQngR+S33S/0IO8Eam+AkypXOxALGx1TkqlKwIguVy
+vck/GEifwppZOaM8gsQdF9AC4ExBV3MiYH2UaJV4rmiu4Qu5ndKY6cql+R6L9g/8/VwWioOyFiI
TjIR2O9RDk0FLDofPfc/No8nWeBRecinJ6Nb7et/VSpOzodSD2C2cxtgYHxcRlh5yZmfpa84sjZX
B32aXwYvUWvt6UyZsPEepLAidCD8DlnTESwi4nZxdBBCe3vkx5uuPqtv0C6m7PEBq9l0DNgb/JBn
02reXuJdkVX8ls8x2Dn8iu+ittZ9pg7d72Rt7i2/e/nOrESIQuxds9ASXvb2Tu6+dTIE07saoE/b
YHT3I5m551d5ILAd3IlIJ2bYpwzNqmtEBvDa6Gehf6Lzh++T6N608118fWVVBqgwwdacshk4IIeW
2OAeJpr59s6GWvi3+BPmNaBCYWnCDRVIrdSLXchKYidZk/mrYubE50Ob+w3e7vj8ktfhdHfejUIa
983EIHUXLqfNS+JpZwl5/8aEavJqb5w5JyYaUXrsNqnu4cG4pAwt7wJR4sZlFR04XOAbgM9lDPSN
Mxlv7NpoLjpXzmnwPxkrCndt0vswaRGYSx8eb5RMnErOXEFB36QcNn9f9JZiHk4UJdWXVDkKGZ5B
mTSPb0Gafcr4AkGGcKH7hbQSKS38+CrLpA9B+u/8GB36qPrGGoG+F7HdgdFeELLGyZGxparF9dAi
LwgZva1VwC1rYbX5kJox12GIctwcsZGegubCV+WpFo+G2M2PpkhXdf5IO9gQr13PbC3TXRN/ocOZ
IqUGaiGRqSKO5lZGgvF51/H4Yii0ZlrntBde7XclIfNC4onZUlnYWw2rlG25eQY0937C2LvvK10V
hZOgE7roBVqLNez1fMKD/0kNZz9HXRvSpycwtWo9T2BkxXK5Mg+x0tdBT1CCkyaUTS9dWKPKvh5I
jTZrnLGmAY/bvgW4B2LzOY7gfbFvjztvM+Dtmqk8CzOmbkSA8U2LOPZpaGeOmQTp0fUexbwjyObf
Ub4+A8MrEgeXyjL6FTCdrmYPgCKoUIR150ITEnxCVQJ+ZVCbmt0qFQ9frt8HF8UBa+aeo6yrb2qt
AsQlH9zWikTTDscsWbWBeG5g1hGVO7VoaNIhxPR/UiotwZQ1A8AzE7TNfJ3JA40BWCV9SG5Gbn+Y
6RKv1DLktSGj1OToG4yqT5Ou0teQ8aaa+I7noL71IFvI0T6TDQLGNsF+Qo84DfZFaHjFZhdOPskX
j7c/11Zi7GIJ49JOHpjPrFt/T9hsMODANhh45iRGRWHxhnzWN4ainEoDlebY2DLqvidbGv9fvOiZ
RIFGYMVGDdwaOYyc8MrZW7p/HyAwgbpXCsEYb7Hty+NQ7dki4SUTJo6TYPyM+b1Moulfkqd8Dd9N
jhGzi4kvdwiYD6CBGaUopM8+Grvvyz2cPGpAA00om+gZpIAfI11kmk1k54rbZjFzs/Ok7O/y3RcD
C8ThVEujMS+iI7fobkZYBeC2UcP99foY0+xgL2rVU0IWjzXwrcE/HzMW6YJSXXgpjhlQZ18M/K3n
gTUL+jk+Mgoob8G5+zy7ljhhrgWF5ZquBHY6+5CLGspfeXqJmiJvS/WtmSP+mbvrdLMGZR+9qR6D
yQBabXlFBou/8RpKBHUiiHPtlLhHOrRFX/c2IPkiG1hH5oXiGwJausAk8Qa7uoNtEttenNoTtmGA
KTQsMQzy+wY6H8ZCB9MwFoENSl0muVEeiMzPf+wKmVpW+o4lXtfXzEgmW4/7nYDTgmYHvDp5kHAl
Y3RFS9A+XvBBklFsB7MbGAmP6Ee2KVjkK0aShPbMaJY8PqQxACbJoPxV0fv7iM90m1qodxTeE6AM
ZExMNk2z2nIAGkCqF7I1puH+uWMUsskYyZcRE7pZcoXWTJk5dfRu6lEK51ECRdUAyB0OHaqkwgUC
qt/Zz9sZQ5l0wmpnpnFk9QEgZGTP84yT3ZI7oucikusa7ywMV5857II8QtIlveLTqxPKn8481Wcc
vPgrtM8nRqbc9qMVVGz7hKSTYbhKreF6S6N1yAFRzo3e4fL4M0dfTDJxfAUQM9fIqwh4UaTaThmT
Beu2AGjI9tAHjKORXYQAJ3BpZflONoRqFW3Hiio24i+6oXP5roj3r1jb7J7GzS1sVMVxFLw832FM
CRIb+tbBNb/ab01pulzXbqXWcHvRHyPqWQIp0x7ZIpyXdFhzbt7NrdfL9rzsU4yUc4RgvimNMlbB
7VaUplSM3OumhQala6XudQCsQ9U913/niTyK7id8CJFjhP92Hri3ptCnpyalFJwFbWVDDG3eMBvs
SODUYjOmYpSaRhu/N9IG2T6qZCxZwQkgPtEndalegQ5lg0pruzSAlwG256Gx/yMTgZGpdt2pq4HZ
OIUrhsA+usScCURII6vCOeak2MGbaBgYos4ou7Ct+oi+8xmgOEy6EPCFmxJm22kPGCdPSrd9hYD3
cQ8EA896DMLAnBZXLENyMatrdkcVrxDWankPEzM5V+w1Fx/JymWITKRV797niywmkgXVv1xFtjmF
GL24Q4gFAY4gQoVGYRmQqw/z7mOrnEXJyECd04tCgkjDqoxeNrnIaYFSssG7E/8o2f2gHtvkgaCT
YrXdMsD7ANp6M1bicK++7kRVLVfCRG15QgbidfAuhROp4ZgVzy2mwTtf1pIfMQKnGI8HCFq1O2zf
g9SsPHt4YUt3W3PN4YoiE/0pd0URarblumnk0BLPF/CUclzWReMEVZKFl3sPjEmWAf/Bak4RWPDp
BBC50RtsPP6iMkX4YjUPWARxkpihwPPUAxYOu3D+drdkMKerfV5iNWOUNbKnhsdEtIR17ApiCIP8
cGRN0A4k2VA01nKt2/NX5joP8TJ506DlBaenkpMfJQ6tHn0fVLMBQN7t4H7rk7fZyGG54A+aGSMX
95rq7A1r4Hq7oQnJx2tBshC2nc/CCX6Ea8/rf8l7LDUuVt2olGpDn797uIV3A6RsWcedVSkYllc1
xuPz+3aB/PkbnhAcJgbaK/yIqBOLNOEmUSJDO2AffMdSYU/h/AZFD/BfiPx80Jwn2TvaAJLBPFhu
CJyK1ZqB+Y9roUCye1vZDv3YDksVSDxKZ5afdLygrCwS6+mk2iCaDfuFK/QMagtQEUtF/zQrBTds
FWDdqsrszIstnFh9PQpvBH737svDHjt+tVuT5VaUoo+UjA2d+itpK5hy5N5bPuxHi2waqvYgqGp6
bN81ITHiDNrfxdMC+BRL0y97pltFRJep3GCHVRKbH76YU2NK9YH7r2hApklGCq/9rmnc4dzmkAR+
LrnQWi8wx6/mYuivOJYZLISaxfvYX9EnwVASg7Q9anpPkILKRDmN1ydvco07BnFs/oU34gbCl2c5
avWlyRdSwUeU+F9xAKPNJdbMT0EgYZ+Hp77lT/KBXaeP7cGMgxk8EB4PQUUgz8Vp1b18u78pr1yl
oHcUBdIXhLUKvv4XSzR8BeFlkUMzbRGaHtCIuDjpV5LeGOSIlzse0L492q2r8GdNLzSDMEpnBCBR
btOsE94Zr2eMSmoUbWnm9Br6f9NIep2P6a2CtFXEOClI9TbGsYW24Z+34h9NWWqZtBRV4HSt41U6
r9kdhbTFa/tipUjvujxcmcNG2i/31MKzis/+8I4PbOuBoVJPFFiLy17toOCTweXkejfNbXq8QN2H
7XytaY6ZHe89YzGIsc0pLNhNB2g/qTUyNiYmrIxLr2PptaH1cRQn3Xli6p19mEgiqxsxeAT1Fhye
o5V7O9XNxJjCJ2A6C34O2nt4fm8I3zCBS/U2gqcaHrn8XZhFbps2qP3RbEn37h9XXej03iMrNuEp
eZg/qDRdCnjEqVymDlQGSbK1x9M5eCb5r1+Ubp4Jxa1HDRt5Asg8Njt5Us0f31hqwD1my0GjfPSb
a5zMw45GZ4tQrPI/CRT6VdyYDQW7Ylf58IVTOiLhBd6MNoVx1QI4bPcT6WEreOU17TcmGExwSXC2
m0LbV1YxAgX0tNyQbbgeEcPuSOR9T2DQGBNaUXpaCLs/9BoF7OOP9X0XRXEM8FZDx0/WLndQMWcA
dextwOxn9NtcAI7KslQ8SUqwqJ2cxyCyxiNUyIt9tS+TMTyGSXxyuu1TZuSrk4BZYbqDCgXB3XGD
BeE7iZifFu8XssR6kmMK4KTaqMouQwJwHXxHvRSYaJV8EBsnSVpqV9mPXK3aAzezhyeO3BzWPaGN
b8ISZYrVEL9UbsxwKPsp1ldajCUret+gtLkfHQUwSApuaca33EjzAl1JXPe3bT6gyOdhOgllcjfW
BRNlnP48+VwHBS3Yw6U0D2xm2eLEGIdQzwmJKMadRW8dAkaJgiMrpIMPAq/2oZezMGW1eD1kUZ+q
W38KvW/v3A1IJyFUzHoHc3TcrWSa5b7gB5KUXEnUX4koVc/LQ35FRukyjNWhUUXlEVfyy1ZHzOrz
ZSx6D+OOCJuUtOHTiHo5WdgkrvfeyKu9HaGtGqph4Xn0ct29qJUi6NzWcoeHWLcqMmHST7adU6R6
PV4BqNAI6xcg0woXH2X9x6n9RtYHOFOFd+IYYpkPHqhtkfYUkd9eblaBRWsprnQBegikzgExioPN
RnURvqTwU0ePro/2z7mWfmz5+TpJHe7zM6nIAEQnL2z+AJye5CAJ76Ehm+XwGbVuB6/tzkjs++i0
+KTau8NPOzpFDM90NjtTWmv15Ekap0t1bW2kwZv17hk9LK6jrSjc8G+Kh00HKNVBx0Y0rPMWOCkp
BiB0HR3JEU/9bNI93tTCyi44lhMYoVCxl0yS4/eQJ56O0zLnS0NBxvDezjhFvZjefD/eOjEadYJa
1SbbKG3pxTlj8iHpR3bJO29VPVILS3F+RDY1T2W+xUxvxP8oFZFUZDW3s0/SHKV/pU4YriEkAMff
4VLWmQ5cCZJhnDuBfW/CXgkX62tnmNJTsFhB3zf4Dp1vBZtAstIc8kngBgvDx0e2LRioWWASc754
7H+aNSIjUuS/s26ICgpkThBsyMTDTzFLerfBEyPpXfRdAelqvbGR1uAUtKwGM2sjDvdrI3ULZ9rH
PEtApxtuQnUuJKvNr6bdPaUJhc0nJARbst8hG+fGhiifs7e9uCYkuNuo+9SCvyv4T0P0uqSFBgV9
5O2v83xnpEP5Gdiy3wSXzwZiQyDVa/Sxh5Nsq7xrt4oGd2Pvv/bRSWyPLglI1kfpLfaxtne9D1Jr
uV1upnyfRJD1SB9UhYzeG8cXPxxdfWKVTgdklGy6K0fTLJTou04VofTBawCGKcRmkerMGqT9q4EU
mDG6bWRcTBGmSRL4+F32jgOsJABy7Ls8glqeekt1ObSjag60IKopnT+IVXi8UkiKXuWezONY+nOF
xp/+GznqeZtWoinQ8ELbWOOA5lUbgTe1RhT9oc2unFTHD2f4bhXuQhHCDty3AEDZDmgbGe3J5R/h
T090GgeHQ0DoJmv1n5/bk4kcMHLKw6Uu32nND3j07cARFCivsLU47NpBwgXT+4PLxj2LthlI5bod
XuSXH5KWvGwwVl8wLxPARRZsbgnOMd28jum50UywjQc8qABkB3T5oRta9nzD1OMlh0eIWktTQr8/
QfywGpCygntuWzcUBe/4pegb03ThvVPjea45Lo0tPKkp4D7VjmvAo6QoWIgw+fxheL9DaLRIsnmf
dP8np1slpooPFH751riVGY+Mas4zB/hr6ufdN8q8j/qzn+7ZiAuR0iKfrL2weGtMqmZp4X12LwST
aPC63RmmpkDI92kVfDsz5ePWKIAxQym7L/rUgnFhxW0VdtKkqVWH0hoCaCkLMgGIj3WBvUitJ0/u
ZxeVM5ED2vQVkYho861iZvrrhl+vUyxlimFJJDicIwIUJ79c7TQWR4vSMNyNwM/nR3xkTAHpqapb
mRd/3HN+rLU18kbXihoIPos/yiTXj8x0bHdocfheaAC+rZ/Zz0aaCkCIgSeBX8l6O5IMblnDSVTx
rBH/SQpOkave7qfPAiM3UWhzlmDUxcTvlMiPKuPWCcet7L5c3mAQQYbKS88Qcb281OJpe/iPeB12
lc19xVs9UDEXO/xzFPxOje9MbQjUqb6jd26MzSF1vPxVMgSAHUeTF7jeYXHOOByt3vcN/JY0ISnc
cK1sIujT2tsv8oo3xwC9WR3/WY3CZ0f7Hu5XySAPbjuQD2Z/9Ks/wn2CG2cqfeR9zsAHr5eS6WCl
a65EUphGDp4sighf08csDOSqRDIQegDmGb2Eb2K4HxkEHrDxcjmQzsUSH3/dtlErgid6OHDsOUk4
TIrj8fpm2depMo32l6AEYyoGAn/951ENZDIKXk013R22ZuBlZ9l4k9ULZ6mQM0oR+PorczNKCGhK
YS8HdLOykyisPvmN5634FKDWYDVdCd+f9EryM3HOyWpFusm/diJ8xR3ObES58aJOvVUYO5d0V+IQ
Vl/EoqS6V7rcPdB9+qfRWS+ckZ26Yg4xZC6lyeqZSpdkfpoUaGCGi3dMhGscXLHxWkYeHdvjnoDy
+G+L61qyM143t9kuh39bHtl4hd9c5KVhkaqqBMXph56TF52Wm5tBP8xtPYwkGBI2R/1+dkXF6BOX
fCBuCsBLvRndKKPJATYxsSe//e2VzXXsI3eoh5/ZZLJqTy7KiBvamd6swqmmFUoH3z/QaPXw7LWN
AoOuZOmvIMVNj/EW/jzqDl86586tYfx6XlRlr27ZRKhq8gAOgpa/Eq5LovwQrBOcmerKRgRNycAj
u5PojkAeO+WYIKBXQCQBZYsBm9EN91sifovdIzG90mbtfltvtQ9SzQMhPrKFf7ylXcXiFvQFz9bB
08MjvYZa3XBui23MTuCmbmVkOnwts9r4JpzfLd4c68dlLFY8RQ+35+xp795mjbu59H2QSxubextX
HgEywGjOgUbRajnzbsojJREvcbt6aUDYJredpHKrKmemFlGEHO4WwIZegBsnp/Lstmf8nBs07pV1
0oUFClPRudB0wYwEfkg77uxhVm7OKYkgiSGR0dr+kCHRnnbfB3gWboPFYCHBsw6duqbPJ/2H+Xah
+NbMYEIlO8ske2RENC8ZpTPn4E6NQ3Hg0/onpqX1iBiAXF0fetHrRVnkwxB6eWMTkY5NOLPBelbG
vHQeVDsV7z2RMVT0VSdIYeYeT9HN2EM4sRWDx3lpfM0j4qvR+toLEWZNwU00VWGA/d3b5OLVG/1f
nzx+BENuo48L0SRcpVHR3tNpA1H4lIsxdDYu/xB7k96+FafwUYLxEX+lIjhsTsoN8nIVHw9d5Fvy
wqsOyk4QZRI0ZHUQurJdlff9rGIevkWZwk4i/HaCVkp3HNv3ESQNXy2/qUFTbFHPZg/ZpqKBF3Au
dPK56J8Acmanyh/HElNAlaknGiuH7cHSRHheH10x7/KSfXfC/nlW1ec32yEqOKDaCSkk8iKEAwXy
VGpxvBk1yZA0iaIGvA+/MC5TnwxsJLwt5PqjooQH+HaxUV47aW0eAbhCGa7oZqdvXQnvLHwcZXm7
aSa2cD0gvhzlPcqeV86iZvI9SOu7tIfl+mukPmnd+hnUlePRQhEKL0e7vZGYHK3nM67loHTMr35r
ztr74I/ESBRQP/40hBSoBn5KEyRccxt7Dbljy86KV5yr/2MyxVmFh8jZwAmyDdz6rgOeqKXFkjiq
UPB4OPnfYEMOqboQ28RCFIC/X+0Yl/O5fyJgzC8rmPtNBa8c1510UsDELE/XMXbOLG+fFgDpKlWf
2JukeI0G+VmLVDgFQH9YXl8zB51bMMJoOrGfWdGw8MyRV8/U5YDbdAuScCRh/CRLYP9HH+t8fOnN
nQpCl4yXMm34JpT4XyJYvIFszKAQ2EMO3V5YS8cX2R2dftX95AfG0+2OhtwuqFxAHeaSZEfUVrR1
ExxImtQ9s3677d8fL2Ak8D4O0o4IXK/m6McPvMUIdq0p3SUqW/ghyfj4B08Ig0BrnNhv4O6ZxDC3
32YswbZwF4kz/lqf4u4Gzx7qyDLP7DFFkhlot8vSBGc950DmD+RcIQ2pQPHv8tok0GIPZ4VBMl1b
jKsWZzgpb6BOp1qdWpwkjx5/XXk4ImdWwnvMyWmQP4C6GuulybegPOvnd1iB9DlpxkAgBWCnV288
Aw4Qu68SzPuD7p+L2IIaulJ/w4pu24OAnM0nyOKF24q5JHikkcie7hALo4Nxmew9gEqIa7TTI1Eb
em3RM60icMMFUwKG0SrTp7L0JkK/pSF1A6pD2ilmIFKQFh6CwneYiZMOF0+VZJ88di+WUY7jCVdd
SBYgA4+7LFwMnkFvvw4ySljheLCLpiNwcEwoZvSQjoAlkFSNcH4Dwdi57PtZ0nolvCCksIfK1YIk
x264Qczirc8DQOpDW5MVFtC4Isj7u00QHBzNnbwGlG6fSoPb1LiAh5ssXJ2LHl8YYKkk0hJ193Yg
QtUML77fzNqk2mTYvH7Lz5GF0nE71woxbAS3V7JN95090lFvQpDEscefqPPC/pR2wnurP3m7sSXk
qxScVgzWxWrnicgFCHZYJkncL9bFhA1HkXlFbfZ5LZSjWR3+0CVxWKzERk6pgxd9m1jb8pNPYWTa
WpAnIYaB9tLoG4swxrbWs+YEZPIibmwwoID/jNcFIk1gLXuQcRLNxZY8Cz3N1MrSFivRURL0K+CM
lrB6a3y4ghIWoG1b30ECCV+8hu5IHLq/SZNJ6xOtWjNgSrFPhTEtg+lcC/vcMX7032s9rpsCAA3H
cGer6p5kSdlX2Ece9DxUL05YnIggLfX8cpqXKuubw8ypdmtjh3b3fznuJMlVOlaAlnBXy3l8fP3U
kaGyZrihnR76NknJ9RABnCH90NGNDpzDmbJds3uJ4iqMOEmGfIIa156eljBuf5FN9yeFWPmPwDT+
u154ZJQVul+YMTHlALNR+hkjF4uOk0WvD8yZAEfGyRmXqYKEwO2AWYCT8dSVY8atJzpiR7bfTzFh
7TQZ5gYHEoAdNKsxQL2jFTWpK9+sGhtXtEZjyLvM65dea0ewj0e1M+AQSK2G2ffN13PrZHYWR79O
zpE8FMqwdiaTvj+7VsNvqWn7uoU2C44h/dzqpWz+SbDZlBlBkCEOQDS8sn+sYDc3zvAY0zGW6qEh
qzQx+T9kjKNOVl5G8i5gSkWH12xu9nOX9x46vMIWqC/JZnCjjCHxWL/LmDt7Lof++UU/DkOlaIOi
r/GL3WxfZzq9I0G/w7F2OwXFX69wA+FIL1vnb7sRdz7stp3oH/RWRq1ePPmCHQrQ2wYuY8oOQVtP
b19Ai+K4E5iEeNql75NJcyoZonbUdfZp8r9/2NurBg6dUwzGgXHrfVUXJ9IffDzgN+XOHIk8+jas
NcckrOWLKO11d64+oWAH/pwsAcYS3cZHkv5noXSWXG8tS9YRu4oMPaBfjfZ2iz+E3A6gKJ3jZesp
VgXPXCSqL3Nj4832fYc3Eht7FwariicDWLxjlfVXd4pVcm7qNGvq1u0Q5Cq15zgEAgCgsnb/Te/F
IRTP1NCU8VtGUsLt3UzO6WJCC4ouESs1arVqEoL/yOoGCTpjNvT8Tqcvz/gPg0Z7v4Wg05OTPOmP
qXubF+H4hPW31R1xpM4qZrhdGFaooXutPSm6eHUkyWByd8zH8zpAax0V8sfMp87W8mAbtjHmW5n+
NxQS/wT8TY0PbsInEB+sPfHMLcQ6VyPPufzpYP/OccIeFPWz9B1BrbeVfj5P2WK8w4IjPCcS0gRP
jIpmk0dz8ybdEu9xYsbD7RjUYrFMLLB1IEDmFj4r+R+yF60elgGosTQaYwc7Z1HMg1M2zn39WCY/
bGx5IZQucu6FDm2NiOQ2ppa5o35hPAlYc1gaFIe2MZViotxa6xFFC6bogUmBiIFk5iUoWQYgCDuV
YCwpf0+HwTb5PVuQW+YXr2Om2TJVmsfytBM6PNndKvMu2EUPweGZr7S6cI83IL6GImsMMI08KLLQ
ojP6SGacjHEHsqZWrnKV9SBAPHs7gbhlSJbEOHA3k4UcikmKNpliMkdL1cygDbLwhUa3RgTv0hsk
zBHi7cLriiiII8Qyc5agT4kwXkXKSTgy664cxp3q9RseIAhFL3+C/CF0BdVB8DMdYX4H+jrD4X2x
UR7O3kvRlop3n7T6IDoWOLRojS1GK8Lx3qvBRFpmQDSiJzaxkweViWrOx+2mSPT2qpXx/PNqOMHp
a+CiPQ5d4Wdq2nPCVoOZAAMvzhaVKa+a9IrtRwNZLgQgAwL3XyGsprqcXLLLHnLz5E3ZgMSeaheG
kW++GCEvpx4jYF6YEChe5zGwVPwCS16D4Zywq9E1l+OmqIloenXU7j8+05kPJmzbAyuQV/1RjHsT
wXypOk09vxe57OGtifWOs2L0W/OCSZQTTj5zQwXlnYQjJfTFjLRA54rpx0MAnu0++TrsE3+pp/vw
+KBmSwT3i39LVCASUs/nOemFP/wc9oedY3whKb91W2MlwYkfV1F8mYwg46xsVOgZ5i3c5dNCv8J2
NNq9kxlOGDbcPxku3AdJAuGcPHUyhX/1mfD2JZ6+YD5f6D1ra0iVuAZVXw6CkGxrGV2VIeQ52V1u
er/0JHjNY0AhaaHDQJOiK/qkvfUSWfUbnCGpkPZT402qSGUBN+8KxN3MzFHwbl6QAPmAySDUJc6n
/8t5HhkXTSgcLqJN9Yw0js76mxYsNj176y1Qi98gJhK9dV8u8HIFDcsfa+0MQHFWMSNZm7SNMuvC
Kx2Fg217b8+H0tBUaIpBvmv4DIa9KNhvBMT2aEbu/LtGRbJEG2gSqtVgBaWdN2/8HC+tmrGrfVTg
zjeXMV6csS6O8BVqhJaSvNCfKzIteLE4Bb5SrGKLgpE/JVFr5ZwZJF7C7zTPqmBDCCdEEysPE3xm
NjTHcqPbhlTJLtAXj2YXBIopNDzPe9yxepZKGJNmHUnWxgaYFjW63s9jSNG3KIjcynfLb81UwNgm
HPsdFjEgwsJodhGuGfTbAFugco55k4BkdRmX9vzYSbDUQF4yeX7WlYPY4JB2F4zRJmEqlsJi1+Ty
oni2t6p8tkAncr3fPpuhql/mCZhFa4iQ7YR3YwDQAYQvt9pJu0notGy5AXyKPbffxTXl9U6ABCaV
O2yPqgb7YR7zpyXjZaMCp6YD6ryy/h9/J1tIXEiFf0Fn3bcpFAu3FF1Vuezz1HdIGSLeJ2c/ZOf5
eMiTnrmqCMozGZGUfPCUHl5TRj/u65oDxj1MgvfNPtzt4xGPRIjOfBJdbdThbLrKVPIFbeheU15k
A55C1/FdHeBYujo7JbK61+820nOXuewKQ+iXsrZqI5wZ757jlvL+ETHrsqrEjaXyk2KKRAe2ZfkL
eQ1ZeULeaLrqIDNUMizPNd9hnL7R1RTTc6psGTENgmYdNbeClnTpRtQOJrXg4otrbVcqhNIi8HXF
7VxNMCaeRRjGYQU9Lv+WoOjD4vJwVuClcF+XTLAGOGfwA/Zzxl4hAKkW68OL84iwCMWQnDmeqQTG
IiEbp3Y9MiyuHUY4Hse9iTdBqb8aKAnYf8+1qZ/qmosY2Tq3VxBBRLtCHkATT9MRNRT1fAuoHPMj
/ODw1bruL8LZ3a+lkKW+CBa1Ud7g2JajzqedaaM1uWxu7hP9qHqoG0PIMHdOBRP+9X4423nziHBU
4QwDhAydlupf7JMXvGCVdmdOiX9JtwhTEC5TL++PUpkN4hqCCrAlpP1C3FsPmZ0iY/+5tZRr5YGi
kjmijiy7060eXjR2WLXMwW33H1mbB3MY7H4h4lR1F9IuvnKlX8m2nhjbkx6vYzRhHNXQ6hDwMEnw
vH2Fk0b96twsRC4g7/a3c4rdNvlvdjJ3W9wj2ghc7R1uEDkyt3QeTnkYaxxcr3W5K/wVCVnXAoTE
4CBHan2ifuiST9n1l+prH/7aHdY0AnrJBcHLVYqRxc1nnEkygKFPPeKwn1s8BMWsCTN/Q214GOt9
Op+g6rtBohzKaLENcGNkHUC0Fg3r7bggy5zOlZCNf6dxh13RxZmtPdMAYGCganrBck0vCAUwymWr
piqDECymdK3k1tA2PWh2eP7+KA/Pqz5aBMhKka7mmILyMUHxgGDvfJeMxmza6gUbh+bgxNEwFuWX
3NzNQ44mmfboKH97zXFosMV6BMN5fZhTeGEnqcdL3FbpLFHpUWO1hb0JtFQbmMnahGjrmeeu1krR
Bp5HkQy2dwpddF/H8pEu2fMQrvZjLKRoyfZYjzzO9amTWRUP+trISKEN7tl6f9hilAftPHHrYmDX
4pQqb07Yic6JKKyko3cB9KANJCwiEOkf8wQxLbfZHjn+HAr2kUj2rfwHbfJsW/y4cFSsDeHhHhSJ
cWjusJDt5b1wjRtwZaRufzIWJm7sujdJMgkOzWytE7Gx4+zSjjp7spfZkEkmqOF3sap7uqnzFYud
bYJvAGsS5tqrToaVtD7Klf/oES+xX8O9tHxmQ3B9GPhwZ3K+iHwp5Qsj8zIxBszq5bR5PQvKyAp3
pMKjnZUPIpC4MJqW7uzhRzgWsRLVrPwfCb1MBf6atP+tvM8JsH2jtYt6cEN8mTVwM2OQ916NgIHI
Z7doJSQRxsf8bKaW/khAtxo8EKKX08EIuSXcHuVneWYj8jWjo5ywfIJikSybwCU07nfOgSC00RN0
S4Bw07ScoFJ0tfjzi/7uQQKoOV4ucSG/3rPmWt2bxfVNNlqo1G8uXIUWO+7YUYaf/VXkiGnBj5FG
o6rdxpbveOzciofQTZitkMglH3tWtj91dxuQ6X+3cocuXsp1rdWTIixPWBI8rjXVZQuzY1u6q0IJ
yZRgMe4oZ8w8KEtx7f/EwU/mCr09jz5c/HK8XIeSmUt7ZYFRdT/Pi4b79S6IvvOeeucpxYVKvIKK
E8kDpGpYuHsl/MmtVi5LuV8FsUvaCjaMfilfmFjkK8UGI+cwb993DNsFxoGcX18LHeb9N/Wm8EeQ
f7fkUbb65SCLq53RmzMEDfXx2RzHcD3k+Fo1XsKVUT3nrZJTliEVzJrCfkDXyj0O6v0KZ+TrQxpF
WcBE2wpfUR8JuwjmxUJ137OUrN3Y0Jhv0she9CMnBsJoZ5CN5SPRsMvsohVarQsVOtoDfHOIT51m
RnmE8nYWHuG0AYFXz2onIjrS6umjW1JiLP6mxUEqfSZ5h9A75oQ0z2HwjPGg2RYSb5VK42pyKV72
NW4MO9WGlN1AB1eYzKZd7y0bFpBxKbkEPB7GLzUBB0GvfcZWhrFOz9gIqww1rQSbrwkGuJV4Ldlb
oQBGIsNgI02nSrl/CUqtmV4X75l3wa8CggW+1lnOvaaOeFAaNNDcwM2enDvUblufGEhJGz0vndv4
rnSIPZe9c2+ieeDW80mkofGZKEA6OrXHP5b8A4cpIXq4u1ppbMhtFS8cX1GzwZURbf0NUKOOlfKk
VdRkSw1SVvpzl5b2OnCOOxFFElydpqH8/VKeZFIcVjGyfIbZpM3D/DkXGt4g3dwfBGtQrPHX65O5
ChvN0whdR3lOMCFnOqy+aafGCZmbsHiryjQkon/difGReG3T9riUekTLF0aEe209XBKA+bz++sIl
ChQmBpOegrBGDT+lVZOnRWB+Ofi/8Wxp241dDBhURM7Evz1SV2isVuyhvupT78P2j8B192j1Cjvp
BynR2Zq6/aTjDAjpJbknAtvsXIe8S4fvc0Bz+RF4PxFBEOKEZdY+GeY4x44R8BBwt//G5JAfH4Uo
cMNLeeKoL5y4imaOMANo6bSOztvdlyqixtyDoqxkwoqt/bjf2LfVj/H8jgKsBjGFJkar7CVarLY7
LLSIutSOjCyrD19RoAAJ9cyeIjBmrI8Vb2BPAFPM2+SCoI1ZNl+fDqxVdZcQTpHtRcBJiVximvVo
f/j9vIUwvUy/tlqcEcaAh3lG9+SZPQuGE+/bLSPgvl9D0l2rsQdY0xy4ycgcXwRxjf/1Qu6qCHMj
kjj8x72S9PaMqcL2NyWG03UYdRcMeAZ8hVVYoFY6+Q0XxeUI7aM/FQirXXE6g0JoKvqXHo2SnqUI
K8yEoWCLYQS+jpeTj+NYb+ZkOQrfzbAbB/iBqmgK6HmIWuHguXzE2egL0O6qot4H/8qse+sRGIMe
zdzYwV1LgTqqryuStFedRCDW+TIgNgfwQ9bOH1pPBW3M66MB7JrvVupNtZZ8M+uSGptLeyZMeni0
c/jMlrrc8iD2HUOk41ISuQhU3NfY9eaZNuHTfdb4UCJ+kqtLKtJ8dLcBTDLQgBnQ1ZjnKmx0Gdea
3ZrNQ0BrtH4kPQRMaIJaO59wFPTpMsKmOkkqyII39TSaNAlbY1haf4qNnrWaKFpVp0qYoPPQJtDy
Enjf38lSWCaZzuMvz+2dYl7vy+q6DKJc1ak2J4fNnrJBszAzsDZQ7PhAYUc4iDw2YRQ5ztqfDodN
dRSFG6XNa3MIxJNRpEVVUk1g1dLABbhRpEzZV/fbmI2scX3JFo5uq73i5HVaV2GVfGKZ5dLo48hG
Xf5Ln/HtBCBf3osArmtVVfb2gdKDorWfEh3lB8vUCiIo126Q+FPIA96FlkLxgOSrbupOGGy5aYcD
XGXiz9JSFlIzozfx0l+52sZt/pZYO0dAhBm94Y2fe/1uwmLT6alOiywJHB59tNCtDPsqL5fYrH8Q
wNJhgZT6EWQGJFVvp77TBnyjPAQMjm4c5DtFsKKeKIREyuqb0N4tUsmKzZYMDR2J9GyUSIjQowLY
n++Gj08wp8x0LyGBMef67SKMFoGH72FYuUCPoec4flpWUnxMdd83ZM4GN7IZr1k+riSQ3ANx1skf
Cz2WrEp1HbpbAvUzgQF5c5h2lgfnXP1M4vWxtLlx5WykHHnhttCVec1ObIOztquiQW2OiNpY4wde
MVQMdX79tIn2QpK43QrxYOuplZ1yMEnGhiAAPbHbecAyOqSmRJDPZAXKOJf61NTug/Nde0IVk8GG
GB/GJDvT/mu7ZneXYuCyUSYYXBi0+8ZCmyjG/LVXgMLugtdiWTrF3Sc7cboy5ka4D1B0vxTSrXKN
7SzQycmrElFNNs/1JDxdyXYU86BFSN51un/SQDPR3L2JzyaJIQRycoULT73VbvSAnOBbsS7eVsdB
vADK9eu48VDljYcD+V0T30YWXL8ZG0lbO8zzoVCjinp4hbrdLNnH2Y4NcdJW32TiK8ReZlJfasL1
jbFbRstUjEdZUrjQiJ8+veDof+TebBjP1J8vJF9MXXpsajPJFRKy4C5+SxDOM2FeAC5ds9AkWVdC
QiKX1d2FPd/tQ9LaLZbioK39nTT8U62RsTO5NRyx5Y2wXNqnFWm3U9eYG8UT79eyyd5OY4q31JLH
JTHR0S7s8irCowc5ID/aw+GoOOSx5jdZ1je8cshgKJaxOiFb/kV9G0HOPKaKhDE89p15arH2hiLf
IvhSfPLsE1I+Oc3pJbqXQse5PEl/KPBbnGrNLlfe/BoxTfohB7z3nTaOZgBOY+3bJzGvrpHdiRvo
jWOpotq0bWoF4Dck214iem3CHKPW2kfDSMjwLuFILuXQUU0tbQjXShW3yACsPqGnzQ3/+8vUPxmN
7Rpo/JFghRPxtMzZME4sT17kLeIksFex9hH/mwasJDDxMi3q+WEVQWEPrFAW804mzhJllJ5+rOhb
0GrBlztCsiaM0guU92ji4g5Hk04gSFbINZLKrV0HlApdWOH/QcJhjNa+Jl7pW5+Rfje4RfXBl2Bo
JoOP0S651Z883XbpSUa3S4dNTp6Em0OHOSxAXirFMqEb0t9w0Wi1r0l8FWwgRAfc711zpGO3Wa9p
OxukthhTZQGPzkFog+x7it8zF09r2H6G5JDNkclHsghr7fyQncM509BuTdhmaTWOWwU6ojDOVU92
q+hYJeFRONZvEDJUCXDvbd0hpfak15GviL4P82i+sgs6e4JVIJ8dgFuH6xFjuU62eushHJ083CZL
+EIsFwQ/494AZXO8dpX6lo+V0xcITignQMuUuCYdsDWN964mZj3RTl7ogVRHAesx4jkyT02j91QH
t/zS03MlrRM4IPnurVeWd+iTZJyEzLT+nkqcw0aQJ2qGzFsuWs9IBR09HYa+bGHBwgJCHx2uZQo4
r/01+NoH8kvDSZClQJfWM8SItygconEv2AZ9oXFBUZSq5FN4ok9BJgaR47rxSfd3W0uFiJElpFtG
TBTv49pQti3TvTvZu18uzMJWMO0cA7Ao+beqlyDH+6cAcxmbSVmVhVGKCo7kxaXx8xysWxINBvFO
JI2chvxwfiytPxv/X4Zz2gKF56zRxk5Mxzp5fGbTSxyGZfSxY+SDPlqUu8Sta4Yibg7LOOQCf/oq
bysDKeBf00AgTySNbSoKYYhxtYnb1P5UGE680kF+2JTz1nKg3zJV94pEMoy/QCT1sO1Qr/52iRKK
CeYTduDCQr0+ir8sTXKx8Lg0jhWDwHejcYi0x6aMRMw5ARLGzFPySZXVfpz+znKceALJFbyBKbSx
1dPPYYs36jOEPANAoQEoegMTVu8dA7y/7Hn4ekHKbTnRGHwNnMdO9lHUZnDYMAlhdcYtTD2niXH0
Wxz/dt0mbO7ry/RxLHXtYSJEUu7Ovrn3lisHauSBYb52iLSejr5LkfSeJ6XH93qRHsQ8bhtRXqXt
hYSAqEO8G3Q8oDAluW77pzoNQ3vGh6z9cwul3GKFcRVFz/u83fptGhhgIc6ofb5glK2aSbN/+8sS
ictYC+VgXo6Ji6lKhTXVOeVvP3ZpBYpCml/ROfdsospCI1Iwz2WNTTApWt8OBeqmDFfWCTg85A8q
n1rt4rH3PYRUjlqHo4IZVr15lAzeTLUGnBqd2Az2K5GVhbPQ3pjbCYDWVlF+5GiQXqFs2s37UB72
p47y0AdYICfQmQhM9HlPufXqKH8V996pBdHN2IiTd22K476wHg7tZPvEdBhogFcChOjKE4PMHykY
HJES0+rmMvS6+qDxc1x7ikfNhVlxuqfTDbvnibrFLxrBnUUj5uFNVI7pxLzpAtxq7IUDUE8v7CBe
4aIvyELZbTYr+8adZgEwy+UMo7So1ljCI6y1EWIEamdF1ybZhbND3+hN70pfb9Bu1JenD6Il6/Kt
cjYGOF0LeCa7BB8fmUz8fI0hCpPJgNWb4sJEjxPa2uTxEgppitzxjvnyJbnWFi0ffBRrJAO4KnF1
mrlJHtcb8B05Bbsv3vaBc5JLI4VkRwXCtnVqD782cW26zbmWAZF2cYCnbxjW6jsMp+uM/diun+uH
0yQTA5+zz6qriJsKO4cjQYNOoMqJAQqSWC6hUV/T1Bw63BNq5DCl00zjiAXn4HtP4/or3tTXWQVg
EtKUpK+ifPCQ5TpTQKFCzCSeUvZyp4UwVwBTew/cmLj34VRZ15MQHHmtp3lU0sm2HZpQt8iQ7UVb
zx9O1MYx4o4v2/Xt64IbuVPAzPgqc4XmU3/owGGh7SggYV4BPaknHSTn2RpS4R57AIvq161tMRj3
ofz2eBYIIJjJrGfBgJTZZgdqieCYu3lY9ZtYXipDeOaqCrwrEsUJ41GPo7qrQDkwCxX55qXS5PWm
vCl3/S108hZcRcurwW6UPqQ8i7W5SrHagmXUFmlwi5oitNxbX5qPbpmm0om2WFyoXWmlxQfYaW5m
G/UlxbQMtuByq2KqrwlgrDUJZyr9RznOpjL0+Hgeja8M5xvZvPrOJVpuFDrnGOBL36cSapB+x2nQ
151nEEksJDGOlYPTu5jyLXhX0Y5Ksyak6igDnzOc1NXYJ3tZ97QexvDHall+IY/i3RXt925XLBsW
YS3uNxCG6rLiG+6mUi32zQJVqoqS9mUqZa6Z1U54FjhHHln1oHWAftAEc5R2AQWaCCV4g9/GCx0Z
EH4cni980f798C4QvDFS5Stz0Oful/Qhre9KbW4p827WP2umuDp26uH8ujmb1vxITkPvkDlH9bTv
kyLQUc6ZPJ9x5rKy5l+Ryt/YxYoNPBfohY5OtCw+sc6X+kUKhLP7L3qkXhyv1PD/qJBlQcuWL/3m
vEfjE6gucrc/DLkGJ3deSYzw2StL90gk0tubPPh6IAl5C8yXsdes+MBXDPK3IqsWp6aNOxJpSZb9
/wy1KXjqyA4ei0bTUXbHzXuvtKaWgIWnAlFWs2IKALZ4ue9nSJ+7Cd0/tgueYomoZ6QPw8okaTra
lZkuOLogqfE1hUYzLiPz8Ntff1oF2NxUfLDxmM7jg4/mr/NlnFZXAHKjXj7zUrICCR2+5aT/wWoh
1CFYZa6s1Ylx8CmqvZierO/xyWVwp2pv7lW/7b3Li6zyOe6QKvzqlAeHoZb1rM37LrrVXkmNusfP
zbxlU3dUcyCyPapXbT7sEe4LcH8pONmDA/QMCTBm28U9yv1AFPJ16BH9PXaQSjqhF/fXBUk6QITc
w0mIANbpwXgX4KShL2GLqyHjUgTEZfenN2HyUB6vKfYLQ5/k0Tnjq0M+xD/Ahe0QsMYCRxAJ+ZmK
VE34s7drV2XDsYYdGDwwjw09d07WYZdsNTVauXeMZs1tts6nNKdrhY6ueoq5c1RHSptFg9Um5Fku
xXRjvaNBrwGRsEMSiv/+bkJBZfFkJHIoPYiqd1/ukR+YnIJwzvr2Re5WOYha3Uj+IDolD3jN1JN2
nnvDtXAdCHMr1pMLmgVVriuxpHezFIIfWtqkZUlrP9+XRey96WMcQBa3t0kCZieArZn4xv47gf7A
L5eTFLvQi8/PeqB5DE9sajC0AE676lR8SJtWO6lXkm34s695IeLeYs0pFN1/MxWp8wb7GDOw4wu9
G7dIETVADZ0c+hExIAdQdq8jOOf7GC8cGVqY6JIFxyvrHkxkdaxW28lPCf09a3453u92kVDvyHsZ
qUx78Xx4EfrmnYMiQfCDohZn2CxX4BEMVY2n/41PsD211hWSgAhbQPD3DYiyPYIYji9H8qvPgwjS
wZyRfizcyYDwx7YzB9YcGLdvvahVH2tOykc8794qAbLvKwTWTKS++kiYxmHeMl9V7taSCa086lBw
Vs6PW7P0e8HtEcSsrNrd9SCMFwb6vpNiEbQSiOqHiYliL1El+EEFmPbT4SNuFZA+wODB63UkjFna
1uyjezOq64+SZMHpUZUDSc1vPLQxpnHyAl5XmBVwFY8aMi420cvV5VTIbz9ZEvVBX8pz/Y0cPn3H
UGnAYwkr9CvfhMFavCGLDiFURG2wEYaZGRE0VO+t8nGwoyR85FSGEpLnoNBY0kkkb1UiV8Y43UhN
4hTK34bBXX8cOFk8/DRjihWt5AzTxy4BKpWEx0tkIdXZa+dBPx7fQXCCHMSkc2V6D3I4fdFr2DxB
4/HhAHmkLph7opI5lL828fADiEkgAX8b/VnQO0IR3NwdSMbdIrFB5wwrxuXQjKrXpNpq1lS605wK
3/UbAuhodjlffVdTTZUZqyoB0TCTbbP9TBrgEgwLfLgLwJ6Ff1i+SudhjksOANcsx3+KUNdGanSs
6SViLtypSK7sShD/tNNST0Y+uLkUIVjZIxhkrTVnz7Dtygq5V7gjS5PpWOaVbkBxbuES9UXHeUAZ
oRqac73ExyWeez9CXD7z6HjaCDHKx5NHsCLbQt3D0pFjMhHdIvUTbhadOn1kXxoWd+iQKTo8EZM9
vBdrfjetplvpuMjFA2wEkvlzLe1vGK/OgIMHear4Ta41t2FCAkGvpfhmtjt0RAWGRM1hHC29E8gQ
FyUm71UmLqiKyKAa5Na7X6XwrTEo5E6UM4L09vt0JG72Nss2zttj63Fj7pgzfury4npGKlNYBWj0
YwCjaxow2g9Xa5fxaWayEig4Me0qnkmQedeMq0KcOQI029bCTdunAl57bMEGNxqF+EblJS0cBfYw
L29Qo3K4vhfgoPl7GbI9V0MoEEE0KzV5p5HMq+MbvsRckr+Ftign/QpZUOJREIqgx6q5w7KFPRyM
XiPeEkUlfp2n91hfUKtnL9Dpv48LY0gYM8/dl9fejmNmNc/1nqZd4Zl1AhOuhLOXI22J9EjLZSuE
2tmeMYCDlomvOwZ7N7gpQ6VZJcGWDk//BTqs71IFbf9/m7LBU0Q8tF0igAcx+hVa5jqyizE2DUmi
D5xf+4O5+6DHOOCX4gDH+tRXugrvqOCo0HFWEuItXS9yxL8x1xVgUaFfgYS9H9hJ1h7NdgbRLen6
DjFGOwNgorKFJALcxy6o9hTGyPMOQHSDZ1g0P7clcHEeENT0cATHDCWg7zj5U8sY1YCZ8wH1in91
ShXGrQd+5XlSqOJAJv9JTBDgoAPbeQMjB4nW4zbTt8v9CLarmJ5qPzLTegSm1PGs9ceuBJ/GCNX9
2aEEYeW5vavUuOgrM2Se2vsk7RpOM4cWFjA4ubY+UUT+0EbmFfDR7ZCJ3DvqyOvlc14t4R7AdaPm
g4rXtZx9sumGZUnERlL7Bu5CHYg7U7NtIQj362DGDMjXLm8j3DcL+m/qWvu/j0tlCkSf/pWIYHTl
KT1bvDuwgfxN7G+90QH7uQBOLrWDIgJDwwUIN6eqjiTroGyczL/F3h83ZasVlGKSHheNxgHP+JaK
uDGEILu2ZcvpPNzWXePdgLASNwi5tRo6UbKWnmsLbMYFFs0qm9gpCe12Z1ubzjblFSqR4UxTdB9X
YLlzhjPCtHTRL4eAY8/gBi/7fb3WpqF3xFlgMJQkUSsta+2pJzeKQfjyqnXWC3X4QX1jwBTzIfCy
Z1obPT5CevgiMqR3gjr5WuBvedLDxRDxGn47MWR+zTmdbT46GCpqYgAfOodK0CxZ32K+XuZpIQuB
K81zDEGWdjDsMFjRgq3O0koULUfZjFw5Tf7cMyMA04kJ9vYNCviVrY9WOlLAT3tZr9LgVUQomQGZ
R5ZNKZKHZpNKamPX2uxH9sCzvDrUB58WTfqlXeYr2VpC6emURz10N+IXkNBQtMTFkaRJt9OHyZ5E
K59bBzmUTKQICs3MnfqYrb2gDcX9AHx+iD1mgepjJn2pjyPbqie3xLvSQ7il2NbObEK9getkFgnp
Cpgyevp8CdsvWPLjhQjMgTVVMjTNAqdoMJFpMAmu3ibfATQY8kjaBb+WX3LHdk/BKrVdReoPWfms
f4UL57qMJFJs93xP7c8X/uUYnAo4JKr4YE6/SMIaJqsnyoO7r3DQRsCXuvvk3BOnnPCjSz2tFQHj
YCDk4iDEKjWNJLbvWTPRXvXMQeAT3bdkQX9NRfB/H92bA7mmbSp7xNHH3OU/4S+DlGfdtWzRRxhC
geazGdM+Dm5SbBNVNTyUwXH7PswVgMyFeB31ubD7gKPL8k3pk2lFtie0sOzLd+1BEtCXEmBaUnqO
DjCozy/JogHzV7H3OKEzi6J6bnYcsdF1ejN4LgJTrgtXNb1Z82IFzKxmwlDW7eFuxXdZofcdD2ll
oqH206JXN/Fjm63mb+/y8wUTgKz3NlyaHOplTgc5rfgSESmjp2hOhNG/zcmcDIPnC/lmuDMtv4LR
ls+PMw1SkHqA04PaIuzhVHaSw0sDtgm2bMdRlz96wplBIF09KrGTEJtF3Mfb+Y5uWUTp9ZU6uBqX
yc6gd6HyBPyB3Ip1/ER09nPjVYYl7MIefB1Ywni0CFzd0mtRW88NR+pJuW2i0gvQzsmwGSViM1gO
h9KrDML22JttdWfQVwf5WKUiF0iPSdY3T9fVuhDD58NPrXdQgyt7itjpVsXa81sL2UeDStqmZWU5
SP/norxCz0AWuX0wHYvqxhKiV0Ixc6+Yl4ydoOXhxcGUILMRx+vtBb5WpmCwigy6UM9c/vkMKbwv
LjrQxcPzX6FJTavjx43diCtCs2qZev5nG7d/uYRXk/oZE69Sr3DIxQgCER0dCb61Jzkqsx74gM8c
RmBZaADWmjugS0IpwmDyP5NXjos/D8f5nnWdpgxBGDTaNRtuE9SFHsC5HSELP8W241MMKHLXfklg
iMmU+aEkW2jCDmQMArTRwIS8rgMDuaM1K/OpSOKqTA6MQ5PIXQFEySe0oryg0daqYX/+mCDT/Cr8
PWW0AnkZAPEAm/UPIT5DM1sr1Y51SGH36JWw7mCHFkvOQ7Z+4Ek+Unga7mQaU2+zfQ3z1oIJX9rc
/rc/qAo2w0nul1BtWJ5/T5pXBxVET9bgNkl52+XcLHrtI+pht6wM0loJTYHCAfhn2FUpggqbbqyO
fDHWAB2//xGqyoZBkj7l2Dr/5H8mM8aVIqCm3/jCXPb6xMK9PUn4GpvKelbvu8rx5Nj3FBe3wz2x
lvcLVbPKNtUMB02QRprETaFK3fAfgtoW7JS4zS0WeY1twhLHaWPxWkaYLPP1mHK3cA76jFxBergU
S2tJCUECN6bd9cK6WW4cfPPWmuNGp8VxYpYAj1REjb41l8PK9YH/fteIGPS8TrTTvelN9rYU07UH
5WEtEr+Gcgrow5KUm9SroiKYcJHbvD3SstX9lEA1Ypos4LGizGBe00Y6Tovm10VhdB7hswHfrg4U
wWEvFgtXJ8JzHIyupl1UOeOuxkXHOq8EREGvYrFfOawCf6qQDnVu0BPw1iIpV8INeeH6KURJviu1
bdlztf/mR8X5a+Labt4h1kvlNs/BJr/k3DDW4AwVFx2zftSnCx/QKvrYEOtpsmDovnaoXluX81jq
UE+lOa4t8EQp+WxzI1sRR9hUPBoWUK/Awb8Y2yUOQWNjptfya/vnvynp+Q2Njj5K8CnmQc429SvF
neOm73ToKXcC6sLj3tq4GPuuj1d6SQKMMCq54s5CvbH8NxUgCsp4wjYZN5TgKRfrpQEMlUoJoZXc
KT1FcswP1cBu1ezX0cyuw59I2NV0HWDCvia5IM15nkhFhLF3KF9ANTCUmtKBPza7ifCk87ZTzW60
yPxLGxhsh18zdo4X72chneQLsSJtkSLIFk297nCT1WoiyAMhat93331jqnCrd6Wh9j43KXQdviOE
K+6byUrqPQyA0Y2Uyu7lSM3hwPmxSR24+uiQDyisXZ3SENX2HKoaXDdeNFnpa4Ry7D+ZWMnCkmLi
sWqyCIpLjwuVhoM+xMy7gvuUkcsQI0fSdqZp0IE3fxUNUG2cGkxhP4nZB+EKwQOjhZHlDONfrPDD
8emt87TU7hsSgxAhBCVaXe5DZ4Ma1cccH9gN8Tm7BzhihKgajUvUQ1V49XJmvvFkmuUNiSSx5QgH
NhgYoHQ7CGvVibd2NP+4YBhHiW/HBrrmS4zCvhQjEqzC9BuDQru1S7uqoKhV4ALm+ZkvzbC/7iyS
73QEldbo8gUodv/knNwGexXzw1a09knsYcXbn87esmUEhM2M7oQ+X1MkkkDF/3fF33CR2ihBR73j
hMVAqT0daL4svdTHoEkb6TE/XlNnJAGn0kaXfMbfo85qjHvcmLUxbS0YxYtTNePp6gFVpDDmtr/J
9Gt4bWtoGrDdmc9p0wLzgvVz4B/05hf2qMvtR2F16kzAIzKnx0hWkZ3nibG/gNYxFsB7llfgp2Eo
8xL4BjFUeePF55lZGa1xwxorrnoXUyk1MTa2re1rnNJwYgkxiW147n6UilEMZ9Lvmz/i5VvkmQh4
dB+n3uhkja4fRMAXlz6hvCWJbDAbnyqxiWXjkBvTTGrb9hQ/5QQX+uA3ACqFuh5fsRQUK7oeFcYl
9ejW3ZAXZRYGkVkEloG/Da0GD4gCFubb0iUFfe33cpKCzoAtaP8Pfwp/LH4aeuVZqInY1E6bdJ/m
MiCg5OadioC2m6BIXVpmsYMIEgtbIhw8k68knYbomz82/aUoC4InZzLrEOKC5SgecA7aXzto0kxP
6BoiS2Qg3WFjPegkO56tJwL/0t6PqptwTU94Ix0UiwULYKNf0L6dbRkoFpKVFmvbSzYebJGVNVA9
Bxl4g2qc11GjZD3y9CQgKvaLO6yh2hSdJSzNWkAEPfIKh3ZzuejsGHLck5aOMSPjtSVieSEujU3w
ZliX5OZ6CNNS3C4zK0GaDUxJpKBas6rkL6EZ1rqLxS7e18xu6J5j7KOLvLTsEvzj5jMFmJw0e27g
3lkoe22xES9eS3EcM7AB5lLE82V5FqRrOqmTpqRQ/oaralcXv9v1MS/7ofp0ky+n0Ir2RsFhNZ8Q
gLF6PVWmsCNlIhHFeOU+n++RUqtboKzV/IuJyADj8Jw1h2du+1FVRk3IE3wS9hCsR7cCp6sjrs7O
0F7tAws5A3VZaXDCWWbrEvsllXXHe7a45wY+53mMqRF5OvbCa525oiNWgf/GaPs9u253htuBar09
wSLTtBakcJJJMOkzj+9vt4AT13sIao1rX5d+d8TA8I/MItKhGW3+TIJEWhKomQ0U9nTMooKaW0XY
CDxScmYLVv+/pa/V9cce8t0ugNpV+dVvHbSDIJpieB/WhSiG5NSJNZfdQZDwxctegvpdgktdOz78
En2Xx946N0lUoxh1pBvvkRgilso4lKveKxgLPZbSCMqDiS97SgxoTqQ/fdhIPkn2eYPG3qjFTBC+
TKCG0qlWVzv9VnOWNjUTM3NQ0zv0/qiV14CVqdIz/hNy2bwPwqnK7v83EhjjCzh826mEFuJYPIHM
w375/qjYsK6jC+IiGHXrIx9qfrMaGB6vtgUYHrDpU8+Si4Q0nl0h7G/pgzDGBwnkLucLvo/iZfnQ
B7PBLLpjSR8kVAn5gFI4b1pW9m3/MpDfyQJ6MIDa8CNgPErkrQecjFCLztk37Vi2pDOd830rZYDD
3sV264wKfrE2O7Z2g026ZeWVHp8JKHz3/4tkk8EQGzfSDPnskI6T/Z24Le78oNYEMihobs1TzHUQ
xR4WVShzdQzcyfxxaJJhI7NQHuannPguyLX8kM3wh8MxvdkDoAT8lPIgGONR5yfoPV1qwpHO4B5e
z2UmgA68FkvClLA2mwocWGzTD62hNxKRH9l2Y+UlP+LnaXg6Ab/uUXcxqsaeqUNqEaNeWWMwnPG7
NKKEUGWruTuJsgrjNH1M2RoBRooOJgfMqS3QOhoXuvgbs5n00QvaAsBeg0yyvuQt62lkQPajcdqZ
2WMeDLecuAaR6peLzqw8ePHCG6TK+1KeVX1fF78W0GhdApqA9qgxTuZFUHnt0rrMWAYZdzhkroMd
ek5K0esoOkH8ajkFJ+SEqpzlflfvp7d0Ca2tId0PYB1WLkZfbG8I/jPeH5aFwJz4MsO8eS/JYV5p
8C2yUthXcSjf5o1Jsu+FtYmLpU9Tc/oexGdrPLdyc6+Fv9x6YVL7S1I0RWxS28AQ3cgwQWXfnbZn
HqlrNIX5jOlHjZ4JrejQUg51taBh1xuJOXjQsOZ5a3vCEWT8hgh1t+hqe51IZbpoPr1OkhhVILgy
3Ai+aiUHMpiSeQjuYOBk9xpXiYEdxDwa/xr7/STccsPYmjWYZ45i/papSCpzzu5R4hEpXc2BAdNE
mxBR39d9U8jH1HCh63buAvZJW5s5JFA3biMeaY+axgeERMZeSDMDAIVz7z+Eahaac1bJvrr7Pc5O
iSjQOWFcxRxWcBd8KYAK/00OpoNdTBJPvZ2OYUZg60fYEmE5IClXEXTbKVPDterIsZAbBqwHrhfz
cZkOkYLK8XGwm6KSgzWxcu/0mLoGisLWCf08iOePWfIuk7Br/C/CiZdF6CHVadpb8+6c09T4ZsNA
V/RWBcWbHi+RpMLxtP16Q5INESk2m5Ax+c792ebvYi49SZNSVXiS98MrcMCMnyl5GVPWNaemQbZA
YAhdl5p+pVKq3Pqu6UcLc3ygg4mt9feM2+9ouvJfsrYRHusSjtzyuJcuEt8I9p6oI0xuuj0IM809
6bsLIVRUEk4Jt1DdcMCUyv7jyuMzNzCa4WTfcMvt2UQ6ujlL48/VoAf0SBogO47M8dZdBRtoTGlY
7LXsjbYAulUtibWroZ49caDqgkqXbyGr0OE3EKUXCDtxwfSfLpOf87xB6rUOqeSuMLUQmAGZFL3K
x6hvUKfdzq0Zv8gA43M76k7OjXz0tEBG3Zl8QSro95Mq743lHDZoF/bvTrTquGl73Vztt0ODxSyd
m7Jl54ClXrQy5J1VDHnxNFWdA6tZx8vkDC0K3pClfSIuWjEOgPn/Hv37707Nm8OEYyhaj0+EanK9
/65v765+8ao/eOmfD2iBwZJKBZv57sYMSuoWqfggvXs/GOO9rpqqTy4H0vMn94SiDcO6T4+OtIax
d7DRturX4z/VI08/gwvg6i3OGhlTUCegjOqA8jumNUuogevp/WWPmCuqDZHwDB+DZ70XTrnY9nw4
d/wOA7ET22v4RxfRF6C7be9mOyqvg+sTZI+2AcCOkWByJZWLQZQDEs2V53iAzAm3U1M7m9jp0lHm
ENNdlaRF0G8Lx66Zi5LUtVZv3hPTuHW3EkVlQMe6zU3x4Q+lBV9MqwLRXEhGcUkgRW4G0WkBq0ug
4PsnsuFvUaAxTa7rhN6CJ1do+NA4e2FNzk5CaoOzAtzTOx5nRJO119lXiebNiVVtWprGpJZWUPXS
21+NJpk5U9bMegpbOnYw47hr5u9NyxvGUwIix+fyl/tTtK6YxUe2N+RVvef2I7bl2cFk4lhtEk81
NHc6qTIa7wkruQbGYV4SJXxGchJrm+UoUXEw0yU4bd3+2ykSRX2DQim7hURZTVlRnXY6FUF7WxP9
9qF+LcSfyyu2WC+kOu0RO+tJcRapayowJOllA4lc80BUl7BGafb/WJXjV8OD60iqnVdjQmuOpXdH
5xsZkUnKBPg56aa/1b5YYjMgw7YtnMySRIZtvpmoQtmaNbc+1FpdBy6FUss2UWyTS45rKyZAwcyZ
KcnYqUvGAE8sDHsATf2B91gWvR7bpCU4YEei4qtEnFEiPwGruIjJArImjGG5NuylMsACmQPVjF7B
yOQO+KmLDp+447SBZ63bV7OJmLMSCy4Z85xEW99eozEr8IZd+ncAzp/NCC9DWL2C6lMx/jwgSWE4
S0RV01VMLRHfSEty8jEnnt+4+gk5mT634jQbzxaUvnQSa8rqebj5wPYCdiTK+q9DbFK5sEXCAON9
DNuHSFruQq60RU1BQsjSlfKdrN/LjgMs6KaedqS/RL05E9o+F13sBnd5glnyLM76HTw6MbMyPuRZ
TQmNOJquFXxbgO7Fmh1CDw/Q5eicyzYYn5zKfW3vVoBhZy+IbHQGH7iJKWl/mGvwR35cAyulrKKk
PvlHFrvaC0H/Lt6pYf0u7nUSowTg5dJ7QYHSxSfN06JzEbW2c9ZYN/+C8t993tFG91PYaRhFdYmv
uuq9Z95WUqYAjBKMwHvK2QoKQZjhS+I2+fa9bMiEp9n0MTVFCWKl3oRFZL0KWxHPrMnKC3BLoEM4
DD9xXRtDAbtn18Zk44wdCnJYXNtZHoG4Hk5r/OGuaLS0WKTCQyCdq79o+NY59SNSuUhdkDGrez9A
YhmECLIx22PbFKj2Jolg8VyEKUlDb8is6Bpr/lee0MjbgwSnMBcfciCcO7nxDVEm92xgxYD1QHUR
kPBCa6DgA9A813+wrUnU68JgGcmQ0q4xWmci9pefnIMbb6aBMJEE31LB6qYgxmgg3iCr8XHqG5TA
lL69OLJd7N3kx4V6gBY7zoepr+5A9Pm8ecSG6RdTMJ2Dv87Qa7hMxBSFkfrxqjK6IKjqKLXAZFc6
uG5KrV+CcSBa7BOTWm3R4mYm7EpcrMrJ2MlHufXk+g3pu55Uq/QF9sXurJA5l6sBM7Q5/zY7V5tt
BzrmyBsW3DNURKP7RWEwQpjqurCGzY3t/djcr6bNIn+PLgrhs4SgKywcDWfSt7g2xESIeBR7utmu
H/ASaUcB54i6LIBYjB/1B7N8M+xC2DxSDFP72xwlO46REMTLX7GNsXQ4r1eeRdmVgPfUk8hhNIXE
BSpRqVBvWDGgivO7xTrfybU7vBkG6A+zRLvVK4Wc4yBt0Cqo06bJOE7Qh/jibKJCT2L8f10YSaoi
QNfPYniCNrcENB6/ufwycdawh6GzB7cf9WyCxextI1d4w04uJccQEMXIUvgKoxouTjnc2B7qYQiR
lKpfP5cGbK6ygZ8tLwkwwKwRUy7pKxd5GplpNnvRxLlWnvt4K12TYZz/Vr+0JokOoPqEinc2AloI
UzAJTJHV+H8iAyQHUdRgCCHYWowA68QHG4loThTqe22idX20slQFAXJNXv/3600sjOcrP8AuR4WI
FB0Sojo5QHbG9umVE9TV8rg/UU7TXR7oBdTH7qwqCdKrx0ITN3Ntqd+IL88xLWQwFswTWo/xTUaa
Eai6b9Z9u6qulrRRbJomF8R2qXUY5ClvqilVkWtWTDThU8yKGClOi0KZVV02Eo1RgLi8+hZeJ9/g
L/3OPj3yytjc2Fr12X+rgoGXit2OViihNOYQoh8hXSbrbjEykuN3o33oxMCXXPtGanZMJp1YfgVb
Ad9sTDaalzfjQ3UxnQDuy6HH1iA+FwOkcW+xonaVBUB1kA834r2G8FbLkKbamVk/IekTDfaAYVRp
xHHhGin+BVb7x8ZT11GUEyS+KTFobfGQtU2P+HHmsojWrugZUgtV1oqTxBbEVG1X3tTO0gDFdAoc
jJo7CLrHySPVrKmNO7yRKHLmR5IIRrkhxqgKzVXaKZguq70BYbC+zg44olrpB4cCVuuh9VcmwyE1
42nHKV9A2SaIqfueBZ3gYd6FK92ecq6RYM+V7CfXWTwO62SOL5bOW4/yRMn0g1OWhaehj2Gh7HTk
PZQsqmp6aN80/0vDKNOoCeNz25Dj6kPaibH/CXWRsxdg/cCzcf8DeRXW3+x4Lw2T21cOEkcKuWo0
RGVUzYMZNnjU9pZ4i/IoHNJYA1uBCMiZyKvTs86wSPdBLOyu2P0fL2e1utFadCf+BDdKUoyeK935
aXbe1+xUuVlFE3d29uEbgpYdfGaSXGo+owtKjqc2lZF++SIENTbE8h9NIhYLX/H8GjTVo7cjDB4g
wrcb17jHw5JEu9nCfaLBeP5MVtvknTxPv9GMYfocgkNDREUaWcRv9CDTBuip5T1rbzRCt4/TYCFl
r34RjetTbksxRNggbmdPidxHPn7EHX09EHmuvWVeZJYrPv+81rtIfP+XKT13QjqcEPgCVfF2zO6f
Kx1/IwH3X7n85eW5PoM/Z/0ZI2lautaWy/ouO1Lq5nB1WNrNVroHJfwz4lqoXZbFIg2JtZz/33DM
cGO/e9pj4Kg07cMgMqJDvZp3wh8zJvgcIjHuNRpa7mobJO3WraSeGFZPhjInojRmF987XPkcCrEM
8XbtIs3CZhfx+XvOsjh7eyL+csp7fb8E8LPzJArDdAwguzxvhQqTvE7RehVmJvwQCBmvigOc+yVR
WnXF3tJq3uFDZJfUcy+nN1Txf2eDPcbPZTt9R3/0T+iVaQCbG31fYyLEQg6GqFI7ZJRmehqTrKti
dQTVLJcMWrcTas4T+xrQ14rS/gwnLTz77q53IuSmIUZfnYVycHinx7lQvZPaFUaUu1bQg2p2QoS7
Nk3I2Q8LfD9rJ/1q1CPiA2dCvpzV23EwB6Vw4CkK6qf0fMvJogbE3fjXbITYry4PTL/Frtj9SrQs
fQ3OyZyURGkN+JLk6mowS9h2SKPxRjxpStZLOsayYwaQvzQ0HPS6jpX53wfsrfUYquNoQlN3CYEN
dS+GILUeGdPaVtaVxaF1lHWwauKecZP1dMvt2clPHTb8Nr3wtxET5lKx1lpmv9mN0X0ZHj8eKbfI
tOKmkPvGj0zwhIe98qh+s2eITN+Yef/sHxRxhrjXoZkT6U7XsnrmzNlCK9xcxTAcc8hgvkqZVdL1
TsKo5VviBpS316mWoN8pl4B0zEbgupBB0B2PnnJHzH8Wm+p+rUg+aD3RaWzDOw4hVjQn8AB0mWG5
ktiJjQcd/1kf1fFsLnxlMFd9+jeq8h+ZWEPTYlpm1DfuuwQnoLr75o07vyPFQpWBxkXB8Doa+op8
iLBdpI8bPzC2i0rS1bmzk71cxoFaNsBMnChNSTmexndb1zQSVxaNwv22P8h5W9G/vnO9O5BBOUhn
86wMYFE6TwpBhhpKhsIxr0Mb9oNNFiqGSv7yd1ioHPB6MAkLqdcRMF9WXULkQfJyOZgMAzOpH2nH
7LuVM4xeQcVHdAr9NHJiP0lGzPLaKE5/KWi6jN0w3NdPZUTD+0U8kPrJYe9h+dHCyFvuyHhZ+Msl
Uf5aeibZSC3erpmzaHqkGI1fRdVRjlhRc2nFAwdDLJUX6OVXFbi/56BB6wAPDAEdidMe81tVrZiy
lbB3ufqjKJXXeDRbO5k0Ph1lJr067DnS24p4sEbY7pnT9yw+QN+1AykXJXTtOLew77BT7lzzCT4B
FLrSClasyho1Kjb4yUmznFeTrdSGtmphwCN68vpViXo488dkfqdvgw9Zd2+gAEx6IBrD7MpeqJHS
ifQOCHY1QCvYG1RxhsaCuwJz0z1vlqIup21Egt+m5MUbFSGzeq2bLIMsbpxGv+Qqp5HAZ3QQlgrl
MPjO88yfvJLHr3fRjWnXiYnRk/khnHLBtz7MNVEslkbw7PrXjUPaMM1yIEWdmNH7BnboyQVGsvWS
1UvjiNGb5SOgilN2oAj2iAqWt70jeGJ9S5ENs8usv7m9YPBO7MzKXEUcQsWOJ3SSC09ND1vm5IO6
hEO5yzFuQMq3FevPwa8i3F9CwhxZWx6BXB3GO2/5M7LsoAHtDlA4JI4jeAoDPL2ldsc7vLa3PYjp
xO80Xp8aZJG7D4DAuXWvHT645xVKR/UKV0qKDToTeIscoBvmvIoyyZjJLW3oBGKwvmn0OBupISwY
yhGobjN3Zq7i4gX2ktsRyVGMp3DSjxmsMESS7mXzxGg2D//NR0bRJ8+VeGUvVjKQi30azknCyRKu
ZATSSJQpRQvxLK+WL9J0bVDk4h6RbvjJVtZ1QGqHAzbqfASYmtrYWplvSTDzGnFFl+Wahg50uv8O
5VLMAAjy0Y0HSDAhfP9RdR1RIZQcDtEVeZMtTyXpF62UQzF24FIdLp7l6+egi/T9Ynz9GDIj+bWk
zVWcsHuZhP3TW10cCMbwlbNjOfYbei572boMJx/2KAxD4iiV4m4Rfy/ZHe67g/3lhbA86LBpj7h+
gKx85YbyDebVrWsxzTmzHmmp9H6LPH5MbdPj09iKtGW2EWeVBRK8e/pmDzVG8pJJtkzaPfBYxny7
+IyrS8O3hKXpqv35I9IYW5ZTC904ThZYPKMUhLagbPLmaDIRU1nYzdQvPzsG5xuw55kDGhyWHSaT
G8G4mQYF4Hq/0P+eUpuWSss8q01yLNmCRmtuCCOUaEW4Cw2hO4iDOMEMPtZOCCTzvQoKYffJJlvz
mj+A3qh09yXZsCmhyYO5XniXuxZAsW69ZCl9vig1GdFaPWO5qiTpIsnESMOPobpYsi6gpw3+UarZ
ALAO91QarT5wQe8PPKqnry7HfaeLrdcwkfYxtOh/VT+1GQgDlY2Qnd3bXLdcgiZpkjSp9vxlnmPg
yMDqeMEByyUdDqMXgwBPhwqiLHUvwHx3bW4ayN8f1eocgfMhoXsPq9baJrfHL++2dPNm0JB0Mifi
M3CvigmR6jgdp9wMkgWAWszF3vt4D6GvejBfbLN4uccMoBmhR7dJtSMxa3RWH/rwEy0fJVbaIgms
9YjTbMrBXYcdMzm3zQB4SFjdW0mDSMiLuN0dKGkFsP2zIaMvbR3MiwsTdnRI7/lCMxrsrdXjH2/1
n2Y6l/hCMIYPNhWrkYHOsg2q0Hjr8TFTgxZvD1dOEDz74bA87mBfsE2/od9YbKFv7dD+G0CPqL/K
C27F3INPXhusFjdPQJks/kZCPY3QqUsC2RQb6xiuQg3E2jjAUu4voCNBjNjr1OqchIi6f/DpfTOX
Al6SWaO3a4oJ91EhiJIbP5Pk78g7f42aDZljGxVhclx3vPSFMfZ2rHlMa7Qjo4yXN88GlpErjhaJ
Ml7VpHSsXY1sECvJlFMcvps6ENPmzb9Lj7n6wXk/myaDTSx8EuIfjAy2Bp1QSq/g2bw8sO9M2Hun
8WGBHHiAakQmTMsc1nR312W1HnztzirmJLoyoUX9nq+/XH/Ld+8UVCGSYXLj7tpjPr4E4WP2pD/H
mwYzzRUd6z5jopUs35/WCitGEqLSsbx3ef3exsXoRVx8NAVQdKmiP0+dkoTogciya15pkYm/H/HF
PurbkTaqtLyQdVwGvfsQyCSK1K6wFnC0Eo/1cuSzUD+nn6dlGDY4yIqqGbdRdBIWP0boEVvifnHP
Xzzrx+iMiM7vvdUvPtasCA81wGQEuOuuxfFpLb0MfUnFK074cix2ZDlvbvqd6qA3LWtcrKbPMRQa
hVGybTuSDNJkD9kBFzh54FKzPBM+fqxly0rui+eOnfyIWc3aWzaW/Mdfwx/+7fov1x33whZFBxgk
JLU34qh828R4yQVZwFVqZtZswSzOAQkog9uu/O60KKnQJVd2PI6GhyTjQMFGVVaR70lxVordpi+c
iNndPjdp8TVYhrbJ8ewGruV+dqTLHrvVHnPp6tUmD9EVJzwnUitvZg/EM4/2WgJjCeus1UrpdFl9
an4iw9AkKZl84m/hfC0CMFtWicfJht4yi+1Pyo/YTXG0pJRyStDtv7iC8fQCIUiGvwVqphmKAoPX
ACTBGSZsVtMwmlshAKe6yzoIhwdxi8bziDfLZqlTL7uuxj8+b3SgTLAEqpo5Ci8YpArOEVcNZ6Pf
ZnUWW+byvH4Ej8we+lsNLPq4aHOmIBRBbR6rB/9AxVFWWMvFp5/1yDe2inA7KJ/+tdyYNDf0a0sF
Zc0jBcMrsT/Y+SOALRR2lOXvZHIWWGyVByl2yXFRcm9CW0HsBpIQyXFBNFt7E5rxB7HrvYJIDi/X
WKMAZRU6yujl9dAQ4FCuU3m8dGpmwJh2YwglD33WiBx1Lr+w/et4sQZun8D2NS/IxZZJi+Dm1nwD
GB0x3O7JYiEdS3hfdZSGFHiuSMXjBT/6IAFqpee4CHGaWFA6oWH5xrw+phb+lOxJlv+S72Lfj/qU
rSio3fKBDKZTCMZV+D4WyHXlvHVYDenbH7skGIp3QkFYorKMqiz4Af9RwIjwDNGd1JV4OIzL6BBH
3lVg9Q1/pS8PE8ZRW5LTm8zcF0csTtSqFVquVSIzdxtRa0PcRXZ2IF+1+3dRdI5kFhXnvrWbSVrc
0DTQqUIazT0bkA+A47tj2q36ZeZa7JrmwYUN6FMg9Ui7pAxHA+Yp5LgwxenUhizgYSKt0iM+Xepe
uIW9xUuc7k2X/7ySBY8kc5EpjNal0+1qJzZDkTHM8e7BMpt+0pZMraol4UtbR0fdn6q/oVwDrbUK
jndwXf06GEPgNTyuI+pfZ6s8dcinuTotEsMeWDNHazXNjhW75t2/n8w43IYovhQoSlBN0wJ/fmtD
j4XtONzIQfY7PDBLjYl1oowqoTQBwTC8Gij7W9zf/xU4fwHy180n+EAVrExGVuhyWUbT7knfVoHs
i4QPOH/L0SPAd5G8PPDLwgsh3CxXN6/uG/nIBhn6REY1LRwgOuNoir+TGuc4pBfw63qx0O8H9BzZ
ej5rKasDiFTB88YDeK98IB3hMHw+MGzzWAGVJbOLzMTOdqe/YBgaBMHtPd8AtWKtT4fA2mf1VU4D
541aUTGaDZPneZmRQsalVvqV8+ZEQtQ39lkStCYQZ0hMlIjVnrr7iGGSxbGy2ASbqYWXMRMgmARs
S7wIm2DNtuMdGN+/bM3rBDAkrLW89p4riumz1gTNB4vshrzN4UvqklnNc9wNbQuiJlNRETet2VCA
iYE4e5QrasnCthb1Nx/bDH7ysSBNAugLo35+DjUoMVwXtRpIOsrgVzq5LDwgnp2zGqoEQFnGeFS9
n4hKQZemO+87MCDb/svgmeoVJsABruNz7sgd9hHhf6x1d28vlnfJ2hmxjLhDVLz46aiY9eQ2o4Eg
jeXRamDWqO4v662Z/JK14SLxXYtCUg2tJCgxtCu8Z3Fx2M52XQZJr5WZIaw9S2QDCdQj9tp4ri/Q
MtM4+B+FBj+FSfUsZmSBRryCQW5FCj4VWqZSmDVXPhBL02MfgL3JX6yJxbXmXb21iftR/h/ZC23e
jqLGE8xczEcR9zBFrgF4Va4Ue8lF/pjQkvTBrFp3tkDACeAq/dpP1k66hUSVk9LSvSTZlITrTNt6
AwEvIBaKr8WJkgjISk2GPlvWWOveGp1lNqjO9aP05+d4RSY8wR+idi6aL/Q1wqK1VWBn6+LrUueT
6BS9ZAyYnjLJrPGGFeMNabDCRORTmjSoZ/h/qtZl7eR+FjBWg9fI+GfWx6eP5tUiVA2KgAYKVM4j
EECNXb8I8+nBDQ9bfyjGTjKcY9CwItebI9fO1C0zfh+Vq6Vzxx3Zqa8Cu81cTIJ4NNycG3NH878Q
1omNv7RxMhz0yg4iVvL5sVgGYH+K3t7Y+8QPgga+NFT5AwBFcMScZjMl6DCoKJJG9oSRNLFT8U/8
hE2foLdyV/NvafORSb9NJ/+B0fJ45xGErNW7zv2OAttvAAJP/35MTLxiGtv7dGS/BGTe3B/LUySb
blBeEe+izx97jLX4u+xhmSju/14YaDkKU1c/0W5qDc9ssjqcEKuYtIGOQ0ANorlHeQgrUDPvK+7e
lAkOc/qSzqdEEt453412mzYf9GvrkRGaXYIjGnwdlFw1PKeDKlhKfc1ds5e8ILRGvjKtxdEnkf0U
ZqzZ468xA8GSdmw6ElaFodQjE/GxGEp4ikb1YQ77Fx2Yes8igZ+kX8mCT3hmQor4UBMFm8nfgRpz
GnTJpdS3+e1BqF967BHTBn7mYqTNNKNAXbNbjb/Up8DH5SNDD5yO6n7hJRpCbDI8fwmtFNKYJf3W
k7vQQRKFKZp67wCqdeLFWbPV1ZEpy6vFK1H9Eo/2ZzCrp5rtlVwoInSANVQecAtnhGFmWUN7dki0
RCH57oKzxqtholP22LZHumhIc2tvkZ+Y7yiLIKzhaJsK+bRsb7vnCQL3H0LdD/CcuscneQwDcrF0
cY9BbFQpm4KQuvkOgfh02Ko0Pp6MYWHYwxfPosXW/j0/88dpLUVpCwF3Uvptquwkqq7kXOJ7DAc+
odY1YoWGfQ524+6DTwfXD09kQna5PrPr8EamAWpXejoKvH8RZjXJPzJqFbqQboVSG93xnDf7rgYn
7QnB2lnRnFF0Ii4oHOSThDx+uXTF+VA2/xqeUB+dVIItzcCxS6czJuj214oPG3wr6EkfLvMK6pnL
yWqCiFyB9U+Ac4IVzxmOEPr08r5oHjPeNmzcGfHggnkzTr5bi2nShmsSdwqU+zEpRRUgebnTHTvI
55hW0rZ5c0JzKD7DL/kIJmnDl63IrBme/b27+sTrV25SCQpRRtjpf5m1NI68SJmJH72uPybDR7Rf
zNdS9kJ8mn2VG2YUie2ofD+JvjU2FBQEt4lRbrVudTX7tsU+4zsrMg6C/wFT4d9JzPxzLqqT3ZV5
9IHzx8hAqI14ro02uUYw2mEFBekLg0oSlrXJlMAPQ4K9hvyNamxCilDE4NViw2iJqs8wwNw/2uso
+bbx1Tpq8n020LFRJdLh3vLeQW+dXuOabgcwAQd+vanRAEdJVmeJ5uKu9A496MEsgjOf7/s79B1w
sp5MTJ5mOR8bNPWK7Q366XX2lk3QqJ8qlQRCitfO5KzJBDzONxC+fOFmio4qAR6yaCaSRmN6Z3pX
ZzWI2U7cvVRdiYX8kr31XUfhvwcIbTMPmluHap8GRc7HHRWdhr9iPnAEZemH5mNwEOl1ztpGmHFS
RpzgQ63XL02gCXlBJClgQz3G939yca44U5J99nfN2818RzOpJSvQnG8KlNnRVHox1b8pCjoEBbHV
PinchcttDR+86/mXWu0dwOLowFKe9A9FZH5yW6KYM3ct4+SIptV7xUvmGDIRJhs/Q/JfqH2fDkV9
JWrhUNUNJ+WNlu+hqSlWMsb44xTyAGYkiTiVQuy+r1SyzHB11zV+mWfgpg9q8BMga4kpxnqL0AVc
tL4UVJgzIaQ4CYMM8KSPAdqg7f1b96MbcvVo58aOzIwyANAnKKs1VSeJnG1WsnRCUsOQke0fs5l7
bIJsQnGw6nJy33OpYIdnP9eEurYLyN6uH8fB+S5rAX1R+ntkztfZEerduH9Py4djGDS+x/e48aYx
U82rAYkLZKnoFz9xTQ4sMG4SfzfS7XKKsWo1Nj/TSs3pUJmtdBhHl5FKejNQWUKOYTVSVa8dQ94D
yBNT3mozCcIdX1e8qbq1EcJpb/LnDzEpEbhfrIdJoNSbJf67TLIQK8w8HlUkuI8EXYx+9MR+QTj0
j+QPyGSLrIPxGw2kohvQR0Xc9ZIl2kT96skfqaguumX7s5t08WgPGpbZ1//5TaW3wTfGCYpIFTzJ
wIMNIkX7cqpM6bigHOVClaN7wwRGpdp7IqD06mxkSh1UbWX9k5bwkbxlqkeiPt0AqTXUUmt3j23+
F5c0pE+Y5lMhcLcrNaSe0bsTuFwZPYr1I3mvngKcLOUO3oDARtLLsO2OV6aV9e6PJvfMsaCIWqvK
rwJxbzn9Wj4m4MZNQ/Pik3OTa8+sZXccdGcbFqkI2CIN7IwSvkWPfQv41NN37duCc0+vxgfJl2RC
+aapSvNehuuEKnRs8LM46DPOv3NBGXant60LZUEcdij2tHmL41ggaAaeeCFs3eLClSP8/NLDdBpR
GE9UIDZQmJbsyImttRo/K9n+h/+UrYYqH6dV0cPbbNjpgW8JCKA880mOy8Fela6yb0CUEWd0AbUJ
FqRIvHF0bLFpqCNhmSZVPCoENFY090LO/L7zTL3F3d3LOSvi2uY8Fw5+6PaJK4pssrsDo/1IjwnE
UPiQ44ON0ySfDqNHaIf/ltYC8+HgkO3JmNdlch3bDrvlxT7Xzn9NuNWXcWVmexQbhMeAeAJkkyHb
zZGUdojpSP1OUhbLKKVNvNJI5NgrkOz1RBRlilI2ejwIT5sdspLZJZWb5Yit8Mgd/+x+2J2rULzJ
Ew50rddHVBzE0Snfg4vqXo9LSHyybJ5tf62fB7e+h7Mf6yp5UpGU8nDZODc3ytPdLnow/HBUfrA8
J6eEO9N9lU0NPSK1OUNZcj8OjWufJoqAxYfSdxFi/34yphmGx1w8Gg57jrTpsCMBKPA8L1OOiPDT
ZxgjPTRsmKJzZoyHEKeDKgSuxEIOhA1hz/jTKFpV3uIFP05rFnR8sxrA2mUMfYpZaZLFBkp1RSP8
GBomzzPEb85NwGOq2KOewGCkMrVYnq1sLAfPNj+BdVJqRN0evpnxXTffdDBdYIajpmd8Be7jyElc
WX9PzJHxWmwt4iUrbpoLZEsvW7qvj5YdZysZKfCulDMUYgcIKrbl/DpCzFWbuGbVQ+xiuNMhTyJ1
1ECh8etsf6sy1NWIqHvRZNY1NtZqbaijnkvtVxnJZhp5jSCz12h/aiKVIuq36juxndNh9+XSw8YH
FQer3Qul0VVysPOcoRVlV/mAGKukNJ5NLJe3jY3xH2wOHC6AbW5ZEusjyLcx0ZHbSOJXUBiRGIeF
V72i0tM02ubp2zP/0FX0GgwScHiix3uyfHUKUlMuEA20LKG6jfYzPn1bYcCVX8W5Rd0kO9/yZsix
YtjKmLhZv23Gn9wi1DRAswshZh5c5MJBzRQvuk/CZz+gTHClnTiZw2+1UegtZENzYz9LdZUbGYk8
0qirto1v6z/e0zBGE1FJYUG+okquZ7SnmrvnizgAgJ7/hUy75Tom+VDP8LmzVPbx0zlrphysBbN8
EBEaCY3qeBaA1I2Kw4JH2+mDievI7mv3dWU7MT32fkQE7zFhSlpGcU2rXgVh9YonhV6n+gxRoRTw
QnAVvFkLaUPAkSLKkbWBziyqkHWluH/X7tkoQtGPA6C6YL+MTLHghF6X944bIH5N3VyU2cIPQ53s
pKNpBngDXpdaOe3ETf2axIGQC2fNP4NVx+nUgXXU+6xGABUxHhchTtAHircHPTiKGjnX37BB3vnM
muRBOTCgwTT5gvkEhMfAepSvg7woulHUfvrjc0gM/K78uyXvjYu56ctSYJfPQEbCM3vQIzaaZcrP
Pbf2mSQ6bUd8to7ma1ZpHBT3yHwjl6IeBJxzA/vtUVWz5R5Sl6nnkQzmVHm1VsrYdWvNGopeatCG
CUKZso0h013afkXxLDnVu6baqt8Uv/A/JwplZpV12/s/TWqOFbd3wQ5MMZornQ2RjcRfBrG5efal
QARtDAi8wow3E3knVpRIAWbGBGKybBiMyLr7b9+mdEXF1Gr72seo7gzFN2M7iIjXeF89k8QLe/2Q
9NSG8X7ChuiwZwrdaRTc4qC+Iu6Rq0F8hL9hZ96T+G6Suk5TYRlRVSz4LsQVgLbfykYSZ7BEJCVl
gBN8fYM1NHgqfzePU2NlC+5fZULMzMw4xIuf9KPedJMIMs0gv+ua0WUHRp65Z3pnH8RjZ+fSz3O7
K911mcOgvipGqZnyMnkz0xxLFJ85AUWaJ/RAA17fbPPmdfrZgy5/idUx/CEESO8X9UJ64DCpdDtD
S94rbVDchaAjdylCvoDiCedj95FIqgG69DoKaOBExwNjLAHQsCVeUpBiAga5ETDE27ILuo4ZB+oh
Tw0zM5923KzFpE1E1ZnovuqH7QAl3ghMs0WhSfUIZNcB4YPTKAwZQb4pjZWv64Dpq9s2gouTKNNO
PddfQ8bIhqp4VQ0BdP/egFNAeRiWqPbTo8qQuXobFyUBeW7persx/UT4ZcP+ukS2+cLiUtKLz3fe
IA+eVPrbnGTiosWd5SX41nfwDxE3LGiJMhS95i5zK8HbDSFG5weanI6xSZIWONqzc7VE2UWM2AwM
lxycSkzic4/v+A4ZgEtQTBG4IAhnnURZklpzVj8LkeB57ajls/AvnT6oWe992hyEuek0SF0uOVUa
0T4iAnwJwQEgv+akmVCuUVy+YgsTIlL0R9/Aq/nZU4pZ6BAwCsCa8XFQNhd6364U9NTshjEL85bQ
TKxv77CCqUcKyrrozIRj3sL3ljile34AjFQgRNc9JX2kQZCt0LHJ92I8FIYnd4NUtBf8W5813MHC
02p/oVtlRCbrBxDGY++KDyhp1pC5cdwWErNFvStgn6YY3bRSGsQcHH5skMknZZxMWofIullc8XYH
Mviln2UE6pxSa6Qx+R6M8dzJFU8BQzk7+A9pBLQ7BjnGhrlVmPYeWh2Xv6uQySc09C0JrKdXQ/eI
WjWGBZCR7YUFxxNTBDRt+AZqTtEQeyAfOwV1ULvWKFn8FpNPWkaNaaHYz+XRVsWtVIkXtOemZR4x
Zus5KKpydgOnSekDoyclGYZeh1OA1QzdS2uGj1F1srykQlgBWx/jl6YanjKZOnx0798CrnjSs1cr
VivdluHPuXFj5ziavsGvn2JHD3TSe4Ke11GAu2GvghbKASCUl19JXQZOkx7jVjMjjwheB7rYFtYv
R5XVwSwbjDucK5biqu37fY8AIhPAXNQIBogChwi0Udzf92+fcFpRdFscrR8AwPATWIWUzHwtL8tX
SGT6vnOSfMrQfbtZ79D4chCDQUG69YTYB7YbZegxTOl0+21e843bxLNB4K3y+nCoyl+F+0L7qO89
RMy/b11JAYs+i1A7JAvVWiThxOrRCyyqL6fvEBZojXrm9yrdrq7lLtob13jugiJfeFDGSfo2b9em
0BBic8UWlzEtSYkZnyikFSzeT1Fv/Nc+tGmGxvLdgc30UlW4fd1BcXqXguhaWsMjZ1wKLUMeWM0b
3sUSN9IE4H1tz1ccjwTroxrbRx3pIbUvmrASb/i8DgZdjwyuHJsc5sZLqD1xUyRYTsBDogAF9LRK
A1efAwo2uo+TbPzC9bdGJ1NBy+7MR/2Xmhpx04LAFrXqKVdGvTvv/pEZdY2VzNNaTiAzZWP2mDAE
ZbcXy/g7TnUj9llFAFMXY9NjT2UPYE9WzLuNROpEdYSbkuDCPFr8/4/r16BUWlbWqLv338yNzQY/
K9UyLuadykIL4s9/BYCVpS78BG/QjnL8HTMVtJGk0QXFgCrFbYHsIEcbLFOqElHiX08+dlJEtWH1
qQTIxPYPwzFdX6rNQ0w3bgOuhBio6O2cuMg1ctPGjftWyTv1cVzHdwLJVt5fiTkLvfmN0h3CTcYh
gm8KJSZvBRqdG6Cm7kF5m7Y7h73SqyHyXhtL4C3ZC57n7lJvYc8fAtjUUqwDEvGtZw2DLgEXcS1e
8aqg0g0rL5PS7oq26M87tjieHLA6EuxrghY6z8UAiKtIfTQJyd9HitSdxcvSds3ku3bPXouP4Gpr
RwcMdhvWzzXcJzn/DVAdO3jvAnG0kYBFlvsfrzvk2N0ZIjOicCzAO6ixlHAxImoHJ3v9qE3Qi+Am
gD/ahC+Kb7ZeQzjmqa3EwAm+4DroY5yYhqMHaEWoEvhzOIuNANWsD1yl24pN7Y9x+B9aNjCDd3Yl
FITrHSSF2eA97XCwKat46DRQ81lOMiNE3ROLclGHySO8CEfus0M3+KtLgAz2f2B9OpGO+5hWbylM
sWEtUNjwoE/asJfumTOSjcooDo48m23fLRKqQYbUa5z45bSnF2EWinUnexqcGudRScGvTbU9A53R
I5JCZDA+sTQVRFoleP1xm/iGyJ6UDeWGOjnim32tUAZXyIf7Lqxe9I4D2gYxABggASqOboeRqqfk
72gyDZ9hJA8vaGD00tK7qWMpPtSgqevT0JuKIpCKDtHRaGaKPoP+TsHKqU5pMqH5wMBT8MGfpQZi
IpStNLd4QGpxzX5EL4OnmYgTfmmoNoE0csP0Deq6pS12FpKU8hdLUEe6g7DKBMsVYMA1W/ddLg6z
ptsExVzBXkDdF9/1PdQ4byaw4R7DYq67wxOKTJQVX0vOQRC9eV/MXyhwuYvUeISlggCt0T2TKH7z
0iRkNE9WaREGObTX409HOhZA3LvzxmJoI3PExl7oQXy5JmanZx1wMm8zu/DCPsDyEtPpr0pbszRm
8KBxK1v/OioVzaX7pGh3+bH3bdWc7QXxT5Z3nQB60U/F7coVU/bUJIEltTIfo4GJHYAq/t+/cyF9
YCdDFbeOUGt59ncMMh8otaKxg3gROM/I7OYJtOrZTtXW7MAExht3WDaGoyoASiIyYeQQe8mSSzAS
TcR8KJLtHEIlpDFPqwJKsqX1ycOgF6CEj3fDrdkefJzqU3s8U3wKgw4Kngfu+fXGdEKIuVBBZzKW
Pyynq9fph5yr3zrlwMuHPNd33W5n9NhPYSsrPFWjSJi2WunCBlFm1+cl2ZQ9gB2q5VnRKMTE0gZu
/tolZ6FIvglQrURT5z39h2pZ/79VQ7KPpEZFRlWB1L9AHMNpcRx164T+UA+VY/AVBDMNPIq9n474
AjbUqMt9uzuyqs6UZNqwblUFmBnrMS1dNfU3jNesoCmN1pK5OYUrqIrjblheIGYuROt7xH0syEE6
PipWDPUJJa+CL4HfDQOVzgpdPL4KoSYfC1jMgJrEJeHpfuzgt4qxP6Ftb32e0JZwcIggSQJr3e/y
/Xxec/JJqm6SJz5exe/eZNrmObrk+4bU9Z5nBbhKj0qiS7e7BMy7gvuQmRxba3fEf8S8nKGSp/Gr
bNh35oPdt22j1zwbq5nafJ4XFUMd1FWETeZ3w9Wp0078PectO740Um3ldqbKcWSqrRvRZ4aMKqNe
zeCpDkswsnWrC913Z/wqsrCaylW+7L1/nTULX0VVAWBZ16N7dTvLT6wRRXN6RxqR7qOBt6qwCaKI
xbaRmZywhk5B5D4IXB8svMzgng62YGeWhaObAjRjfg59ruMOHqYz/ju8UGNbzeffoL8lKtmpSpC7
CWWvvN3JNH3LZGUSSG3df0ugm2/EtQqIxd3j8DlX8KS6RvIVFHOGbVeXobl3Ftlpn4scvkNrBqf/
nFZ/mxyfC/gFj+iBBtlF/9mytG2J+enR6eglNznKWkYGYZ4AGU9toDP/q1rs/TRhxzQb7FXwmYXl
R/6NkCUwNk4HcmL34IoeKXVuE0PZTL47AB5xIdwi8zI50yj3cZciRyiWvaDT36IyIlxOTdFMWW2l
e8bJJIL6l+ZQNwHh7wmbkv+Vuum9gGOoiDPRUwE9PvJcvNW36e/7ZRENu3toeK133z6wNVBthxNl
Lga6s2RCQBTRbfzGPTCUxcq3d2v9wpOQLIAnG4f/1u7b9ISp2W0foFL8tUIOmR2lPmA1OAiKOgsQ
4RJ2XuKi/q0xggtHw/ThZQ6UeAdt9U30cG4J2ZZRPd6DdC+tqvHviHd9QJAotw5r+0FiarP6UJtY
i2sGZUqToIE77JmUGZdD5/oxY2/Oczn5+MpG/YI3ExwuKEGzsR+29MiYXGAC38u4muiVtJ3za+VY
xWm9GDp/TF3S3t09L3T49qJ0qZjYq8/M8r4dKE63Qf08px71hcsqqQ2kqUoWI6aPtgQj6i/MnK+G
9NdLdCu0PeT4xWBYWUTtZhhhtgnCMiey0moeuItKz9Q77zAAjTQepvCKwTMBfJzAl3mtaCoYMsTz
EzTCqD6h00qMFbKT7ScwohLBw73YX6hrpclwbmW80pIU6vtQG6s3RN/w4oooz8em0pi/CKyXRxX0
X3w3ANWCar0HMoJOYhwuDHfYHxrajXCcaDKkZiVKJMwQf5d2ZHXREtZLOPr/bNoqWBVOk24utxDo
OdqpQMF1xRuRQ62BKGJ/5XLApwoDQVw0T5wEzlYRqWgE0Z0PAw5iE2LwUInEXWbYesis4H+ZvLXY
ezj0DpbC3bCxfzCYPt4Tuma4gVhwl9LcPX/ok8bfOzHIME0/lNWYfzPa7X5niId7ZuXY255BEWIH
+YF7oBxx/AxqGgEZG3x1mu8/BIrVK3dm21Z1MrI4odvpLd89qX7pIDy7BTpCBqUxzvjCi9HtTIbS
eX5bFspGzIOgfkOWPuX8XUsDjq7oLHJk6o94JlejdCmytr4aJuChtsQ4tbB8Zrok65qrDwP0qB0P
H+3/zOLG04mjFbAISfKsxjxvEhTE+Vr7ncxAti65VUN53izoqIqeLECS24+GlahNaMGfTvk29fhX
mN3OtlVAwGLonRH/5RvWgPx5GH/p4BCcxemBMq1EkzNer4nNCIFYk7cDmP3U5gIM+D+FXDU3d2pP
5OV/o+Es0iWasr82wLBGWvbSmK3dAWP/E/q+Uc5wqILuDJD6PN4ob20v9H5YyoaHELYUurjq4nNS
JpdEJzQOM2cHcNe9Pu2wHslBdw8kIazDbwVeE8YjXtfr32huffj9S9VQ5O7C74Q6bd9jbm10Ebfp
BvVpRk3+gjKlNEO1sHRFvBMXcreihHq5WbZNHSGaNDKY3WUyr1ftIeOjXokK7zvF3ClRGC0u+YR0
Rsa7Mz6LAFhZblPC5oE7Xy4Z3RrEbiavonULl/ZnA6k198W4A2+/7Ts9oYwmMGZdJshSsiXgqhxH
5eo04B1gdokNwR0SuS1oNGLpQaBw29bOJuP7C3Jn1qjv8zaIubIV649zSBODa46ZJorHbtL3qMct
wVycj8ccKs8ATmg5YUmYPfzHm+x60kgTEY0I8awK+FK0T08CxvDa6QJUA+bkZY4LdOn+YPQdRzdO
FUaCnB2V/Pmso/dwiQb58AJbdicY8dy8+p7GFoQnfaw+m1PPUHttgqFxWY8L9niRIxUyOhuzCweE
1r90dx9mC0E8EU51Ocn7nv9SQBKQZw09a4KcA+7pid8FReXuWMP8WW7Y+GEbAA/S82m8lqNgY3hB
6O+kSr4iPSik0mi4iJbkvx4eGiUbAYBdtpgTzYZqP0vPAc0Ku2XnyqsPHI9MKr3U2sp6/juUcFrk
g7vgv9wahgfd8srzSrqoUD1vZO8D1jFMkABc520sKhUE99V/s83V6GAfvZvBzgK3nmx6Hk2/yPH2
X6FANJ8apaGO0z3k9fezmypDAGLcOvVZvMt47v2v7xnINDQK9u4kgkmVonsCwkrhm3hvT5RO7zX6
KGFXKsw/O7tXxDymqNnratYDoXtk3ZHnYH5wCXcD7yNxxTTxuChc37eONovrwBGEUtTMKIohIIyN
jVe/opcgtqXvK9pKIwByercf2Mjb5aUJtZ60bpF0o02pHEA0MgarsYGNysnHpK9fjFJ5mRJSzJf/
OXiqq1d/1JMeXB1o8xUSGWQYY8qD/sZWTxqr1WQ4SBXdrDRnGz6XKkUEmqgbNDKqiXwKulJjh092
PyTqIoGj14YFdwv9aMKJwB+3ElPj8qU8MIJg+Iuu2jmZsxrhVdzfoP0muM5+hDrXFxGWYmUhBTG+
gJelWFtGR/GYpClEJoto/izJMNjruc8fzAOyyxDnRTm227ubwZnjirPqxLg/iO4IKYA7PsShx23t
C0YolMMLC/alkOp8smcez9b3/IXcQAS+dHWUbHdvttuf2TMp+bl02LOvvury60QP9nsB/m7gAict
TpOG2ceW3Avuw3lwZ58EOJcZDTK4Qp2WaJR5ISqYtjhZ+T+Rs6ASraWktVssCPX+1GWZCm2pv5fu
hBY3kllYmuZxnzCgjENAwuDXRMBb5whWu+zUHdI+avsszz/W2Zaawtuw2cXnlIqpVFcMkesOFLha
Hs1wHbKzozCrN0w+pOK7nSUQ3CyFnfuBqeZ7zh8wUzAh8j1/bp3T1CnLOz8ZrIwkvjTmM2fUlXKX
AmR0HeZwOAIxA6zXw4vRL05iCu6EfhY0aSWoU+pDrzQq60v9q2uovGv/jITU9k+MFV/BuzV8VREX
Yop1D1lN7We0AfTWNrD3vIQkO6UhSewf7OspOMDXStlKPvKq4siTKvqAcgVCxFTVbE2QQUfH3szD
B84DRi0XnjqgZor1mkpI7aOOl4c+kBnA2nzZ24NSFyHrodzemzaHVwUtJqlWW/W891tdIENIdjYS
h0MjDE3DzQXEZ3BpSF15Fl9/109P9IHITMoa3/2DKlfeG1kdHdb+91fc33h9YbKxIu8oNeqIaPHw
HtRXokTsQ51SKG8Bc6R20MyDGfMWaIbfstlQh4ZQ2gpSHj2Q4tPiEJJ8X+hnmWpQx60uZU7VaKKj
vUqWqQobqBBRY37JTn+miN00P5z0jlAxXzhILPQBd6LbSohbv96s2Y2fTeEa0h8E/wpV25kHhars
PXVy8Kg3DIqya7Ntx0HxBGZcz3hnft9HRm6his9WlWydlV2qnXQGMKqy+bNDTAfM4gbfqqkWlydj
ouuz/ftjdTUaXkBZgAVA2lUYdf4CxJ2cXmo2J2Xqei/pcNsfeOdSbxUoy3RDvVWBfGZ58wmm3ZbS
AhtSR+jnjWgukEjMncX/OA3vtLo0ojyvQ9zdtyYhU2l7Y7iZqaDSgxMgNVCbBcH0W03F4isRvibt
4GjAwqKVqd1CUWpoC4WMzEZuiQcaiJ0CTLjwqVLhB/Zv1tQYb7KuYoyjvkY88USy5HEDfZ1ul8VH
IYHde20CfdhN6Dw2CsEDLJogkimKFJJb5jDp53x1/E2iAJreBcS6M4LoUFCtXXGM1MF/FmrsLoS5
Uyuo6cedBMi7TVWJK/yg0XaDoK5qMyzNmnMbbHyAyRenXz/4+GTN94EsmpoYTeClvdfD9BgQjYQm
UJcgOKS3Y25i7LYLAsmnyN5PEocJXzGmAftdOSHc++8TkObX9d6Nl1eSvgEVuM4krsBEo6HhWBLS
iyYCMXZLFrrimAH7+ORImo2GGOOt2VddQT0wZYZwm7JzxCOxXlZ3UauhvmameOpmCR8dDM44aOGa
7EH3u/gId5YSwe5+xBlBs/v2t8/V0XgX53R/TyNSsiuIiIH9BlxrXrSQm61vbp67QnwlFZjhFjQM
Wwgji8n4QY/HRXtXTWzf53sNT2kBX+e6q8CWT4rTwvJBpJv/gQvI+PzaJz1BIyIPTeqrV84Rpn6r
cJ77yOai2tq1XtxkEG6yY/flYrI7sJIaKC2jdb8ZNkGlOyUqyw2BrbZRx9MWbDaQD3awYr81mIMf
8+U8oilQwv0EFw1z2+lhpT+W7Zjo5QObGKci4Gf3kCmPaukpoV6sbH5Fs2ZHKLz/axvIW4+sT1gL
IvnhlhE4AAmY4X5av1bNeXihcs3hGZ/w5bOI0ksjAXWB94eGKSqJnEZATU/Cm+9n0czrHVBaUV5o
xkfZ3uorDH64q1ucc2aQ4UL9FUQbNt6vNPWEXPuy5JBiVMHnB0BAgjGoG+FkgVok2zqOhVi6GesQ
u/5VRyt5iD4Sdru2/mwWxtHS/glgKMy9eie8/X2LNYjXnw7nvGZApG68Sy7tmKgHERXIP0HIEstm
NS3rj8BGgcvC82kBYlNXfXYDZ/5hMAmGGiag/xGkaOoutX+l+7pYacS9tFP7nTURV/QFG8B3tjag
xxuPJfil/Kk3X9mtrOo9tSoE13/bKn61BkcrAduZWu/x+WGV8LpRithoDhgMsSb7VzzFxtgh2sT0
QxHKNp2V+7+Gaj3K9m5j/pumssrzElHTDkwB6VGNgwNpn8saC7bGtFkO2q4kYyyJG/XypKBxJfxn
I14hhg7xYGtMqoT3/cpPW7TgNgYHWdHXDoV+jW/45qTI63Lh1/4zdVVKAqpyAqnLQqhaXtPnKOFj
W9yYQuf5wjKecqhLXtvoP9GEisSCM7QGx25iNc6sxxY/WrtS2VA6MiP55E6/XeQBO9jXMRC52Kn5
I5NOTvzfii4fyineOq6sLfftWnXD3DepREZekyTh72arze/cNsx8hfBIas7txR0qfwI1THRfvp7s
tPJxbbZ5WRcSEFoPIkcOXL3g5MDXCTy/86wnvEmA8Zs3lll+QCaSNigYJwQhmgjL9T0L4vMdSe2S
Wf13CxgRtSZO6H2F4okTo/muNjQpRCP7+V4ITvRhXsPe9Q/pmb5vuTl10XQ+D6aXdmywOfxInI77
BXPiDbUFgBd44+izfROUT1+GruRm7M2S0YxpndxyMXCzvbt5/aBQBdzvU9S/cV+NDnBuuZDxU4si
v+XuV5ZuxAPQEdQv9xf93ddZd7Bm2pzlNr+kA07MCLToZokUkR73pCqxEIq3AccL9hRAsaO0lkgp
bNrNPeLgSqFF5w/CDEG3R8G16aYeDPEqOrWNzWMiDBFH4COPhC86+n7o69WmjjBjSq1tYflTxD53
cehPBL82JH1XK24rKvomXIgiUHF7WS51GYlhp27LaTmglffvsEESJzggf76bKlL0C24jXemufowm
5MZlso6WX/FQXG5GuI/3mgX0wvy706H5BK2JGvxve1KzbhfWAC+ZkmI9GOXJSbrE6WFiT4zKEhsJ
jxHzWu2K+KgVymM0QU8XYfFR/jA/IC7ghgMF8KZHuFMMLav8zq11JFEkI2MdTRWe+JwmMujNqaBa
Msr/63+lJl4upoM3KXjzbLLeSE+l4zZs4HP/ww/a/U1ELqwA9elx46AoW+TBV896NHnTgA8cI14T
Q1CmSsSzlPv8ykmJtUIGfF/lChLq2C1yGz/Lzd3HdwGxA+c43NGjL08fscVLi+n04TN7nO+SWGPV
qfv6QkH+bdzPAZjJL2E0YKP7P6GZ0+Z0Zb8HHkqMqFKx1UxBahUCPQXsf7TV6KD2HTDpTGCGV+r7
iPul7q0lk6KZ8ScQGXltQc9htqssVFYlF97LSJakwWPltFnz5KGgfaGPJ5Wyu39ypKe3vejk7nDg
HsDyNU1JkvIbOeP8FELRhXiktlB4IADqAgPdi9Cc79setByhSmr+MzbsvVewR7Ew9kWlnwTVGvDU
49uAgbpQfucKB72bpzLKQkwIf52rxjN5TYrRsDvkzqG9tEk047jxEpng+2zpd9wFRRq2GjjwQCXD
342aSm8ntAxYlOOSurD+mEHWWA5neyQSOtyyZKj4hoYlWfMOYcIgYhO7YLhXZ3J9ktr4kC5noAG+
f5IFLGyhL8wLtQAlY8foiwA5qRCC6ONqUYK5mlFPo8vqpvEeArTn3K51O/Q+XPjOi1rWez4Vnvsb
8kg4xeeqTw61y0XaGXWVynQowFhiQBPR8Br2ps8gYy8zKNEwAqezlyfHdTHxOq2eLP8ZaHHd/v43
KAGXeqUI6X+5Cx03P5tY4iIoK7wpw7M3pf05PrpSBMdKS4yISrdtoOICK1rKzNx+k901WBZiRByO
VyL7c0elCmspbukHKTt4/GuYSZ0HDaGhkDdOjYDn7fXu7yZMstzU7e6NGKyEMOx79sXDCt9BfAex
X4leb945Qbf1+3GzgHPPSy0Y+CeHCOKmbugV796ei/ZFn9c1pinFlTAl2cQAlobSVHLxiovWDXDc
HBHk8FwhWoUOz6lhO4K7WbMLvqwgenSXFg3Z3p/4Ql4V+INhgcM8/MRZo/MSFAdFBGAuciohJ1RF
qdUQIf5EemMwK4VIJtu6yRod5Ub8Gfe/9fCiiGVFy//131Q0bxo2ZtT720Tr8xibPD/Z+JTabC8T
nO+0ND0UtSwptUjvZdDgrRN97PL2DHHBFbwvOnI2CaehLLzdAYZ2RDSvtvAbaVQY1rwwH03NbG1N
mgJuk8U5TI7nrHTrs3+rFY/IVHqzMzNOYz7D4BNzSCYA343rEUdb9z+sQ9u/TrqC1mWuB4UMl0G3
OoKhprvRi7scF43StOjzjbHVcVgqWw85sFBdnFIXY95wOcpSV9scagx4FBSPfe5PKsT/kS4JSjbJ
ZshmquvPr156sryOfPX90sV+uvJ+tCZgvhk4C0yMHM2HCDbGgEuHVYLXL2gqhhYck+zKkjNS4vfl
dcsXD21Rb7tyIl6cIDGv/D65CzvQH52ny/UcdZRaGl9sPmYEt8I0z7OUhFI7NuW/1VVnM3DYhcE4
ADneaFkXd6rPkatrs74wTws2JvQy8iitcaRkZCPrnlwT38F/aNBlcrruZZEEfnJJZTWIYtKfFgFf
qYExubvYzwzOiGe0r610M+tqso6kQ94JywaqK9Og5bU4KefgPcPm/ceTB8F7F/CCRoVSBosHwfHs
tMjrPR4JrovkcryhmpJyoP0IRjV4bqT8XbsDrL0sAOnYejV4tFg9lmx190th1aeMEiwg2D3zbL8G
n7O68HJ9CFgoRATGzKyAeP7Vn/5icbKlIe5MLnYF2RbhTHhWkafLDb4/2vDkD+Qu00it126oA+Fx
IgdT3ZGX1qpKg6pZb/gv/NvwW5aVVnQGhzVmvXFkwOXdTWWEctUBj3svm48Y1b1M+zEXkxjkPzNn
anCJrxvC0UbijVNmnYNDwAa4nv0sRasYJHDTe4UlewqbirDDArb5wrJETv/D8FX33fR6/+4kEpgn
pXGRbWM8Cc9EJWoJ1KIMR0bZEjGrmSnVEVgL3y5WPtJ8Si4P7+PvocGn+D/1K86A3trTvazckCwg
XbKSa7W9s5m8sXdcxRpyaT95+vqY2ksXQQOZUtzmdjtOcvk4ivgHfWsU0kn31CENX3zqGKXk3GNC
4wvFqTF4X8qk5jBDuAfWfu0PxKC3uSOG+mSzQBSzfxVmrZo9Z0lMtRBNjdkBvUtnGMhAjNQEeFvf
pWj8solYeZpoB0RXGkE8mao/350tzK34PljBdeAn1mLJXj+Hy5qI8kRudccHxU/9YWUvipSwWCva
cfrK718OQ2SZByglW448Uy2Aci/5RKa8SBsTQEn3bHqjNpchTzqo2HlrbfUc2yVl5K67o1e/0JZ7
WrAzqyE+bOv1tSi96vAx++sbGrRIcA42a+9V6e3RqCJixrPjJxGPWQmtuRSV7ZV1jRY3U8WtGXAJ
xVZ3bqrVihcFvb735n5TnunqLWokZxNJWDnkB85b8BkQwcFuSLKnAoVHt7hhugSIrZKs3df2pC/6
hpUMDz2E8NrDDPQFHt9TWLMWP3/sizgHW1Sj98BDGlPJoISsBle5+rv65SslAQIokq9gkvRD2q/0
ouKmN6NKXYLMCI7vhYXIFxxOc0LD9D4UbU4FW4CEqpDUGTrD7+TwdasCLmn2srVTPuTxVWl2mHMX
XkQtyhWgGH2T+DQWfGJCPXlPGDHyHgu332h3Y79VnCtqlklSCvevvkD+qBe4S/w7mruoZnL9kcr8
OaZBFRKYsvuhzDE0cvpT4pcDO4PJVhv0KxUA/NqC6aDa1m/ECvYscvJcD28/16h6R4RNSCx+nfZs
I1NqY2v+FvU+7dctXwLL9PvqNNjHWpsfOT9a7SJ7qxf7nDC0RdI/btXqx73XcEFi0hy52biZeQPB
0lsIQgnyD8rGfQ4GXKp/loqoohKOcXT3fsZi5K3Cv2ImDMuDqZQD/9pE9I3S2s4D4DL7rl5NUkUX
jFDFnqKFA0I8ISGGUPm2xnayUzmWwCidMdhetgmnnbHea163LlB27iF+v8JXmn2H3QVhu+5IYz0k
lVTP99ssNpHrvdQ1wdR4S6sHNQIia5/qejnXtRVMFHLC7T+soZNDTsI5g/lD/Ctf5iPy7KmcEAfV
TclECEqJkIRNrQMM1+IsW7wZi7PNH75A949GxDN09yHhlNZ95bklZIvPBK4tsjMgIV3cfL1cIl9l
VhYr6rMbkC+Q5e7RbgcGofgwfdAn5XvmKNrz8xMS3HEcuXMWIUxpEjSEe4hHuG+wSEvNVplnAWLH
BfyLve1I0Xshpnts20TgOa8eyBcILCwoyhyJocqnVPgqfFTwvFSUh6YIwuDkSss7XFEQDoxTFAZT
LrBpruFj+dKRnnlkQ7OiWVaBDfrb2m/rt68Pv/y3ZjXTaJ8IRjWhKNlpI9GkevuHLpshNj0BXXE2
41iQjVDsN4t3X/8o6Jvl1huDfnq8yCv21G2D5ZzTkhjdj4Et387MznZUUaMUuCwRfmTlxMhsWv2D
HSEgJgQJxpnp5fzBg3/idt1ypC6II0X7YFJBmx/qQ8BZvUZ3g97DOOiuHUFOra68zMZpdIs+ig9o
WVjWMkJl2QFOLP0+0dHvRvLNqoYexYblzKd/qprYE/DBJmIRJhs2zfaoD5loKP7A6w9I8XCJOrtc
w6mvZrtkC1FL4XlaowsW/ughryhm6/gt7/TRS8gD06A/wh6SOetILgVE85tvHljkTTrPVFwVWLEh
+gWNDm4FbDuYldvdj/VzhuSh9GivE5BkesvPth57204QMMiRCC5cWxinNC6SrS09S8NPht4iLMLv
R/ocHOJfbKDqCnsKNJv+vGfaDfWDvYErlOCbRi3mYYvnURqtDchNXqY420GzSbkLX3rIUNRYbJbP
dKhESbTL3nzgYpQiSaQgtQiVS0IznptALOEHDjkl5M38jV0AMcGwdz7wSCPJlBQmz+QOqObNroWQ
lri/gW2Hzju/BM3Dg/pXeQgRfinYxSPQvvmXmlHP+3ctp574UzFMugvoP8qsGoH/v0SsyvWoLMAf
t3xXn5mDQ+z7KqkixWVhFqaiSCYzXg3IBjJohuz7zqOrDr02JYFd56lwkbWdDOQtu6yNiQK7Fs59
I0gXVl4pP9YmvHwVSpRzKcLhsWs6eRj7T18V+AOD37y3I8YxKtV67vvdr3r8IjbJncRVvjww6oUD
8pChDB/vkLApRdbw/BF6NIvj0lMEtyJcEO/bi+LGyDYAC+01jGk/Tr39SJ3M2NnikKu+EOwI7d4a
VSKrMltxbENNpEg8RWObFtJqbCabAu7h8IuiuRGT7+B4YIZvsUn4WlhQVyU8prWNoZb6OfOscKPn
ADrqO1YlD1thb05cOjT70966ROnb1eXgot/9V6qg+jvKtL6wesbnOcXiVjB4sKviTcaICOcjzSKg
03vpZtuowIaiCj2TsKOCf6I+zVHLzu9rpsGy4d3vdRIQmIn681HjBwBN9Qygx64TftQgxMmWKrXN
QI5jHtvN7IavvGUI6N/XIuLzXxHZimXk/S5wFjCCkR5LrFKkX50WyXCExoOdoGf1kU/Z1mgrBPjm
0G7f2O7uKrdHfK2Rx/BJp7dh7mYAC+o0KXiNsSBE6EjqXoHNx/knMIGDtX0nvaRdkFACaP/eMT5A
v6qY5mXHJeLg6EXatqnBn79UqFblsbUwl0E5jXxKBGHYb4RcSuuKzAtQuEQvSIc0KqQJxRAT+4pK
IeNbHnbHmdkLC9kbiRNQuR6cK4rIGjvatyPRso352axi5u/ykUlvytcLMc880IJcf+pSRRRKt+8T
jzOgZHG7FI98x3MG/bgHexaDS4jZ6flNPPRqBEw90WzvdsTz4PRJcmVGmo2Cf7yBAQ0CG0wIBejp
Z43p0o6uN05DoEJMVb+72p5sgVQIRcwE2TsGXbEqxvsVJOfaCxXpRarhcv9dIG+r4TvZMv/yYJwp
4l5W6GYYMj8ySX9FMYynuWXpOcIfaccGBsuz3vIRpew0ffkpdNilTFRcq9ANpjQm8BS7xwBPPBXK
9Y/RY1NdllAEP9LrEyBOp5n+RwS6SHa2OXlNA1loFb1erHCOnnwxYsfYa+TruFA1+wfSwmx7qX28
WWaUuWoGi97hi6egnAh6u08UlvCRhxszG5rawM4/czk8l5ZrVCWYx9Z8kyWdt6sbrqDcBm56nm7T
SAOqOlQ7GUl3r7db2ZRkM4mt2KYr8KGs5GkVKtUA0psQkV9X/DB6crmGAkCU2+RaxINukBLqJT8Z
+IafVQW5CCtfPEspqkhzvSx1E8/6ssyiPgCYLvW4u7VFuvnnzPCU2FTwCcb2V+VLUC2n2iqh1OaH
wLz0sSkMJJCApobfA2Y6SaEE5PgQ0ddMCMrr9FdrERKdU2jpckRrWpTbU+P0GjilthygfSWLbk6+
eSg+sOWsX3qTIvHQMrnOAD21e10wgEMEkvM2DEE8znQqHFfYIPut8EafW0v1G/Y6MpfiKZLVFf1l
jOn/U9+GWCNoxy+ro8U6aStvlM/z9qUNxdPqnVfWzyO16eOoaAIdfHcnOFyt4W0ZfAoWsMU6Wy1Z
UQ1WrLOrJ0Bo3XDZx76fObSAF9TfurFPOM0khiY3kKSkEROoDbIM5UkNLuT1HWowYwX2agQc/eEB
nxTH/3a8Y0zYVvx3LmsVu1E65Ls8zK/PTe3sjBPE9ZH1aHeoYaPeQdcfO7N8QCLINMGx2GCT//GC
y+EOqArfr+zXiSWwXVyU9UdeX+xpknv05/yxoHPYyszjrUFPuJpjMfm0HNoTE0BAfH790VtN4C+t
enuHtISVfDempgXnudCvtAde84kaDxea7Ki4puG0oENsOhAaUOeMhpSQTURyrbn05ykzRlys/ueE
ujfe9ngmIGJSnWjEjyF0NVoLCFgFtzR15hSw07lR4/B9KVep5Hs8Mt/aGyVrKlMarrUv80tu1Kvv
C679svGpVU4HL8YnNxDRD7HW2KSnTxThYAxwwORHudzsoTuXZ6OLBtdXT5PisQnK6nfq9kmmX2mR
I7oHbRL/xrV27g5n7enA1X8ZxW7Tbzvfnhxc9QOYjk+zsAuY78AUhIBjV3sgVVWDCmj1w9miXeD9
e9nRatzceqM3ZGGLXv1W7xa5xdy+0ANbChvP56Gsnhj4OeCU+mo7LRbCicV3r+ySfhkhhjtDOAdG
d76jJmaGOYbt8954rOugAWTzUEjzWJ+2CGOKq/A7Sgzek7DiicuGUXOHrM2qqHM5EaZzKRpIkHBU
nhbNoRuT1JHL2uj6zT/pApAz0BQh1GzOAF3BV0Bq8a3nyS9DyLwtZ3KJO3QEsWyAAb8YvDefaRjm
mgzI4LenBuqe5mz0GM8iaufqVZyAx8jxYAkzWHNCPwIuJl3s9/gjnj0s+kSIlepilVN96fVh+FEq
YUWuq2NK3Vbacfc/UydTuFHTDyq/CknRRjg7OSqeox6l78ftAAej8JrQ7axE3cP8tYv+7RhajJwI
eTsv9ns3qK6jn+n64qIOdnUYXhbb5YL5yHgYC/P+2LM7XZkGS/vdI+PRJEA6WkG8ssk+deI3TvtV
vNAJuO6SV3I0Krj81vpGdRLFt6GLBcW0mgr8Kod0ddduJ0DRipGaDPgRSqqMt/RDAFTyQKhkoZwG
d2pIzXRrej7mXI5ITMgT8jCZY52smmGtEEZu9V7soOSeJxJAw2dCMckRl2jOU7GSFhs3T3rwgO7U
PHCZDg6tOB0xl/3mdYMqRqlV563PEgASGBLHq4R5fPx69EI/fKL2ou1f5q5wzEL1ELOqr8TgwFwV
rnITIgijZTSXVlKN91G9fnnpJfZAgN84YCpQ1QHzMex9IQTGlEzQPqPHrQu77Ibr8BFUJFxHouM0
Ld4zhrDG9nzU3pu7djFJRhv/hOuQwECiTYwCrCul1dyYKMvjshiKT3I+eWkncUz0ye4ocafJLIaw
sl+Jtb9bcOGi7c5HVmHs2OsZGXeCNTYGoPqus8MmPXQdNmJmxbU2RNfXENkaohkef8p2ZVZAZWyo
yq/y1/WOhwyS2Wn9hWmELXQpyfhGmMdZxVJFqjnTw7gBTLn/074d8i/ImnAV085xD1FLN7Q5Lyf9
nR8UPPEgSIQ4Z///LpnQ7/UCWdugpUgPh6euZZ6Sp+/Im4d91tPBXgzOSrawlUrf/5lvVUzSc6VY
SwnvZwaoTI2917KV3obq4a7nJlRRkCB1P+HkM2tI9r+SJq2xHTsPeRgkJzPwxe1qguJTUwI27kx/
R67pikMYI5r0kBNpoLzNrWc39v3Xs2UfP3VQ62g0cY6AvUFGRR+rC1/PxTWsuLrC/hrJWFTWZS7J
nvzanzE0ja0MnO5gFaKT2/03PBWGmff29QGdftG0B9VsaW/AcHFXgtp8YViWAgMAQOwvg1W03IXy
u29SX+2gV/NlrqTONhs7WTQAefFykgWB9rE+m9tKwkJDkgPjAsjZ7ruTAUneqih6vCHuHYB1tEhZ
DCO2iOx8i7uw3TyVp8vcGFYT8sg1ZNWRwDAx9qia1BLc98Tjtn0CxkfuF2dqwHRKaiNdCGL7qVAg
//LzhBkUuyQfKqK4Fj2c3X9oCNnaxcYoH0N303apTnl0jQ9KhozAI1+6mIX33AZ5rJchSP958jbw
dPYnNNVO7+lIT3lJB0T0gkR9Kuzr3voz6vIapwVXrAJRQ4FAiM1+vdEt0a6poFeOgRY3N386yhlr
Bj8BcBCbV8CCZh6j+w4/J77mNK907z7e+wR8mlI2UNbidt6FtAeT10gOg+c+L1r3qnrexg3yRg6s
lgQAzou8cpt3oYvc5YQLNwdwNeTh4C6EFiDiY/GDLhnS9JX4NkmwjkOpZpPDH2s7Z5rxidQ/Xh17
KHJQ1EwW8KnB9wokpGDcIAuHuUgt8WCDqAOM2p4KtRZli4O2/440xxt4z2DnUPp/GGM+nDWy0ZLi
ZMkFnOpINCo59STm37vd57VJx1PjRS4VZuNQ8kDSkz9lVhmMmTH8Tg9NG6ALFndXaEp1JFHNRUnn
DBXaAiCGFr33jQgW8MpDJKvqX2kRW5qn5Uov5Gmzcytoj9ezSgf2gRSBoz3KhiKwCyohFXryhZEF
HP7Xd9hj16mws3tbZEEWXhh+Q9Ago/U2gSFLt40eZF189nV2z7wECq5C97pDDSQoegA14kzriZsY
hg7o1HE8wEo+611emSbE9rpLlIzuACypPb8mNcfhb17yJ44NvFzc032EoR81dT66C/j5b7w0mfU4
Ps8ORqfrVLhQQEqrV+1nAiktFfm7syNIj2KNysaFu/gKUUtMrc4/q9o37e8Oge2OPoeYz3+VDJMp
xw7AR4sEdwWOmNTEWE0ZK1IPQuWa/ybrJZFHH0KfAK5boOLtcoCV5LM8FjvpQC29RatbD782p60a
DNgfgs9ioAkmb3GRS3zAzZsFolCl/xpP7PQEHpSDzpR3EcEAgpHLekQRwlISMyMv74TBU8vYWU38
fSWVgQ775tIEnCLab8/VJWtk5K3b0Z0fHU0HYjEkoPGvAXdoYBUq1WVeshqUyns22vuyRoXjrUIa
MG2UIMHVFCftZzD0+IVXs5aueipNWxXXb0xzR7EZINYL/2l8SII6RsuKYez8ZZxPM/xcpd/9JdM+
UQg98bN8SxF5ogNRTcRoSNb9oofijwDSfmkbXYhy0g7YFyuENylDNGJtlMeCWo00Yrbg+FuDulEk
kVhuGny2bS9rVsH3uJX2CHpqqVWUNqnUo6O2rhz9VrQbbReNR9PSnvmJyE0KuK12xeMTqN5amY9s
bNbzdrZ1DpyYhw7qdilat7JHhZ3ung9r/ViMy05/vdEHb0qE++5pTgu1KsIBFEDqNKOYc3berBDZ
Bzj1nUrNcqjpG1KRr9x8CF7emY9jihPb4F+jqYEll1VfOeAIOnlOUzNCm1HuWVBUbbB72G1L4G2E
2CzKp0CElzkBCb16mucF+IbfFRtTPYspKSOOR1DfCBcaxYHNCwJsp3OvGowC3TsBmYIF3RAgkwEo
DkR0+ekKa9F8GG2n/GXIoZh2HrqazimJFl3ArtPHTZ3a4hcM4X5EOzmZCEExQG8kxUUrzHeN9Fap
9Pi2nxIcjvlHa5bPWCECSQsAPSxa93VNNIxFFE4r7WW8dCAJpbhGuwdMBswjw3z9vizYqCfIXmI+
Wh1Q7zWY7y354hS0M6aSBv/u2FXRfnYqBXC0nTXl7uDB7NH6uSCoAb9djQxUuIG7b+lBQAmauZoa
bof3Y53djDkhgeNyqR2EN6DiSf7NrKuLb84M0UZCRwOFuidFnp4H3dZf57tQK1kA8tAIQn2hlA+m
M3w5AgJiJpjBNIdV/3k/5DToinaE0RFpw8sMdAk9pwl/9gN8+daESD3EX7mhjGl1uW+MsW4Y60RP
o0lJfap7awkgLyJ9cE6oiopj+5bVWl1+/vyHq4W0eniUVRXFDv+E2xsp9jjEBORqCGE/sBJcfpSD
/fa9Zxrl1zIA1tweG1AHXXrWjjgJf/dSRKxmDI3Ps5+t+/6aQDwtlM25br4/fyejTWv3UkNQ7jRt
snWpNqL3+aaXx+00bDL0cuVKeCS74ParhbsbkBLW+ZQ+hgKxjyG8eQPw2hxdTcO4jD1JB7ee1Z8O
1LjKlMX4FVOiOOshIrOOXKvDn3YzAZvoGj+kZ3IYnDCLGcvZxzfir5Ugxa5BiJMFFlhuebwGpnbq
4RBsWLQnak6u+jzT2hVAN/eq6N2tm5eECmA9TmAjEKONK1/WHJ9EhwksPaYNbCMRrwd8I/egXdVE
MjHBFuL8OxSr9oEJqpPFurI5qyVk3KXhQDVkKBlAzSg2t4j6gLCfn9IW9tm/j8ximFYj/9t65Elx
UrBXVudQ0KYUT3B6RwPnXyUtbLPcczZYFrwBsMmFcAJ88q0IeOehutni7/d3YZvMeYWUFuE0LcG4
GOWp5V3oyYCq135rzZI6Unx4IxKlwRzeY15RM5IwEDB/ACvsGG4J3oogHmPw2UBYG9cN/LX+1r/c
yhV9A+aOMOMmQZ0R8uqFweHcWsGWrE6cpxmkQlqBM+rP95BanczsnkRnV9Etc5N3aBBR82Y678vF
MyD0AhASW7/ERFDFgGfzsrYiBKTz5Q5Scbz9fo4eXwAFY+X06HOXYVCpImikhrYKe5xWKW2Dehd2
YiGzKeQX+HUk0NSpTgIbzB2cOtpnF9GdLX/rLGlZscpr/SKG3j9qbr8IE7jDiSn8+mQQUygMnnEx
iG/mfCjj+EkxV/E9XEkmG5qZ1+quFoAn32otsvpjRTOIMZbpvWOBSsCjmyTIu02iv/OTbzzHhIoW
WvoYmktEvtF4yLrGOC85oo+cXjh7YZWSJhR9f8A+6Vj5zKC8N78OZruCC3qmyjY02oB0oO2DyZtn
L0sdpeH7S484+L+iBKPLcFDqqgpzeZiIow/48VBuo440p539PQPNDcXWJSiVwY5aiVZzSeiCBaDL
09nKrVKqP495SpPLEMaE8PZbUHeqU0VM9uXNzaZn2Q/zR70Wec3Fc+/X1hHCier+ZQhVGzyk/DFa
5NXZJcwhhIc5/DqP6r0MF/w5L3s/kRR9eu7zFRJh005e3L3b/1wq2U38QgTJBP5k+9JKQTBQXJv2
7sQ+rxriS1znLjFmRk5EpqVvLnsVe0t7hJOTNnsPp6AP8CdNAb1C1ReER0lcFxR/PCic/I6+myOy
CnrnbAOny6VXpjnljfhQmTgNgIjlI6UOEo53drzMDLCKWhvVrDN+OEonpPv4R//WJjzVFcs2WaRd
YEQP2XXdVOcb0VHHgDxGuWbdGZ2Dg3MR8acF0KYnAAUSrfU9NS1d1270kHhtb6r4rVm64pLmDjRB
tN/9skG0BC0yB4U+XJakfOnF6pkA3d05Nhn9A6dw9DRuhjxV/Aupf+IyO65pmaeW1h51I5RAhA9B
3mv3g5JAGDHiS0eNWidCGgiBmb6qVz9dk9+LtGNfD/baMqmjTpg/+mkYbYRv1Zdm1zbyDk/+SaDD
pxhxG+J5t0MJOyP3Ag3QPL7aVAdHpYIpct5yBWn0mUN6b2gaJyx3BRbVeKeGwEE/SGn/orQCpghk
fWQ1iRzxCPmoNsjKqTbTabfdOnpXoCW4Kqhtm40+bZH09WvyipRxSNqDkG+eWnU91J3MD0tT2Ix/
KcMxz+3TZrM/TAehA6Hjz1QlVreJkmYa6adwZEe3CuHYNoZjcZraeMKmlQNEbNwHGp3nosy68GW7
8MOFKvfIwJdu3AoMx2B+nbs74sGHXMfICkE9V08iBKneq9hfI2Uve0IlYJXZKBwXQzE4MRNpRvJd
+DdQcUOwdcftlBjoYq8ZfRl0/JRTv1YzAbTFRjMSprfWqrpOdQrA1VOloDNJYqPmTu3tXGIqO/5Z
SnwS6SjTUU/TwvVB5ByQKNqNz40rriMss7dhTSTsDSYnVy4tGXsbwvQQcpJMrtsEhvvlYIEM1b/k
NI+x439ubrPFukM/OQgehmuFDVvnIXjkAFibKIXk1dl4nwYvn8Inw8y6tJss+72oI2C+bCwncjOm
CEaGFvU0noS+elRjdizwYS9VcI1H9YL0NWvimF+IorqqZWEMSOgp22MxS3A00ILpaqvRmf3TmcDG
oE8bVO1qxgK8dL2ESf7lL0bEYe/Fk50fNZaleZ750EVsxVAnmSLLUBii8Pf4UZS5kxOH3+3UkHiE
6S0Z83ZdXabvhQBDlBiTl7y9gbB7rbcd7OvvTIwJJ8by4ZiSRxa2b/L7xxm7lb52p4pPe4mhqNFQ
TM41Vii4XLsh9WeyoOqYniUMZRiCS6KbLUbH26JVqnpuwtqVQ0ldbfufbtB+nROqFchh3S4xZ3OQ
PENlik982KoHMG7HSx1X/IQYKEqOIHI6K8LEBQiD3mI8FVA9o8Mg95YkQcu0XDT4HpAEIus9Ru66
XndCCOfWxfbSeWeTzM4FLJfKBtkCaOXYXP+JSsC39XY7tskJ06PDHKTudCNN402aDJ7dG+v9Ecvp
UZFN3IilTu5jUzw6YBX9NLw29x/bp8IVn1aH4goT3CfS+OUzkniCsMkyOB+TSeXIpmRyl1rDccgz
3nA9l5LaBN6GeLNC7CIuBB+Hu0P6mgXHCftIWKGxPN0pkLwWgCTBTUCU5SzQzI2wLhL6/1NRh5+6
5mScwCf8wNPC08uFiBmoqe2ZgyzoYXl2CBcY4Decd1pAW/jBGdgb8xi9MlsikcastXJ9/9/7/GUk
1Kq6zHkZmW0g0T7PhPTubkQa05i6QtdNuwbHORu4Bk/TBpvuO9rrvvPdy0Lh3I6K5dJkdVe68t0d
dGIHNiStvSPZKXkOnS9uIPN7lQsHloiRDm6/jtzETw5HTc+hj7DRAvvPhT+Tepr09Iej1mvgiE+d
f8/RtMQX7ms0QSlTuDiaVzWYKfSaV8UHGtwa2/06By6s8kMhQ32Au7ritQf4tghEp9QZZgfwbzf6
evgTqJkd7uXTO/NZ7YpJ8bWcw+LXoqqhwjapMBqPEcZxomYjGiADXeas/ZUivBomuhe7yFmuQtSn
NqmKE4kkZlt9ibdwTTuMCXyYUAS5LHcm8h1CYxudxnT61867LfOFWWfyMzpKCGbtOCmoArzQ6F+1
3v4nMCLF4gXBsgqPlUPM938MOU0m3IPj1LgIRMqExIvGNklL8mP8xtCav87baweTkrCJgKl1YO5S
R75m+JOR03rQIF26DFMa7nx3hu4oPDQZ4cnj3VLGDuPx7x+eTkfH6HDfUtgVpBicD1NOCdECOWIG
yi3VOTt9o9xpm1pJwMZuIaPA2XW+vnZ+O76yzdYMY/jvew0zgcwa4b3lvbnwIosRpjPvrz2VO0cU
bgYKjnAQ1uUOn31AlJDeEVOdyNnrgiSG07Z6sfLMnXlskL2HBbomJDx4cBbPuNbWqwqA88l0HCMF
6AjqECW62B3pzSGwVxhsDmiWW4SyEHIlQNm5/K167Z/GT8tobrB/MOzAa0ox3b/GzSqFz47Q9JFk
tmiduZqNlDs76WbjaNZ1bDbcxJcvICqtCjEljNN+25udT945VBf7Izy8iW2tpFtLQrHIAiGyYUOC
rARHIZz0Wy68z3CKiUpOF1ApnRAmjTs1DqC8snrrcTZF/aqzdrHzas3ptJ2lRvryO0PT/Rs1CsEM
e2AmxReworys40yUFXEf5FjyFecwfeMdx0rfBJdn8Jy0jdXV/g4/QsNPcRxtE6gyGfc7/gz5QPPs
VugGDYgbbUsL025hCnAxVYLmPavnMC/xbXPS/zjFgM9l2W22Zzi+KVxmEsWUss2xCMvoOWGKYQjX
4ox1qTfoWO6/Zwcge43NqLsw5RjwHNnHibXIcnjPGipQ5NZFDXgCtE0jxXLkKU8rprq+7ezBKH+m
qIe1CfSofXQzube9CwsRO2fYfThrOqpJwSsZh/jlb6tv4IwFnWhEkfeDmAKU9goVTQuz138+lJHs
jCHaVO4Gg4LQXBrxyt6o8XvR8E5S1b/8/RKnNUSHmPIeI103lVP0ouuQm5fspE9sn5R6Dp3/seWu
ynz47XAhDqxA/PUF+7LrzI3V/nzTKAjRxCTqZLkBH4w2oYROIjC2S20CgZg5c6ylomdTFfigaEqC
oVLvAuoHNjwA6yx9p7/9ZDSUokFvqecGlPF7SsvjFttjCOSIoFpAIHtqOQInzsd0dmI5yJ83Yj7t
gDcMv2Qn5s68O97k+utZHncmupWZfCAcEWskdV8Ocu6+/AMJmqdDugKT2qW1qRTe8UusWY8zja40
jxLogU6XpwFu/ACED//hyMKPJvf/3+pUDfGxU4SRBDUJHkJAr8f01QVgof7AthbmNQ2lTAyhXTIm
8UMb059xcfmpEUcFxIhsSAySEvL4hG8Uc6kCNkfs831M0pZl3DlzqRrUc5lLVPzej0G4W8GVgmyV
7/O46MU3/dJ7/lLHU89RJ1vIGnISNF82ceeIgbH3xuuvdZY5Dti8FoMl6XU5gsjy8k0Rlt4f4FLh
RJX49QaZrkPdPL0qSJ7tG6CKWjEbPSl3tBkwvpxQ0mXaIa9YgZOI7Gu+yHsk3W0F3MrJj+Z+w899
w5Zvh/JSB2djsIRr/9/9ouM274Ykw1jYd8gtXQA89RJKXtNlOX8i1cJzNf7oZC8F4oQhZJdmvpnW
bhYmDnsAISEfcliJxjMU9xWClHvtby3UwWVfP0Ssm4wenW5TVgRMnJpt7L55aBW3BIAPdLafXT8m
YvwmX/nSGmKvFi7rwn25SCyAN3dq4tII4sF94G6+f9yqo30iADK13+2X25zn4BbZVwPJwxzIVKHt
YasKSgC0NdDBM4WYAmiqdVP3yhSzvxteeK7xvbkBAyEEdgnm+3jDxoTiExkqsCjbtwZlSOAHMUwr
ORrphVX8XEF4XaS/KNqmWg++lZyifoLermFlwaYIFd0he9YpURiRnkIxp4Xb2lFjI3E/+aA1pFg4
5HMw1E/cfWJ3pl3jCWhW5qtlPSgPcA0BJAoNcnaptNsDXZ2qRymULKYvArMK2mTu4u7BenLesYRK
wp5VYqa3IxIL3g6k3MGfG1o9rJOFWFvPy8FknG12rjOlKaWAPUgOfQ2S7ED59T+9hIg9IXyURatd
R6L7X5kt4UwO8NtzTxU7tZNVh4CN397oP3aGcozRfEwIY2XIYd6b0wCzAfTbKCkXSqU2qOv+hWDN
NpIVAIBHSiJi63Ty+/U7S52UahkYyHeoVSSPBIJmMxbWQf2eRZ53OJgqNnmRWktnPYBpC8lD4Bn1
jeBpnqxAPTJ3k32fSxpoGOEieo9Oer4XCcNxW/qIDalABUTnFhzfOaahDWu+QmWw5qX3CvHHFAgb
dSMS4LJcC+A+A0HAtkgDdyazcM0FSBmL3Mf8rpWMF3F9pgtk9duNz37Mv4LXjqk7OJf3eUIyxQuv
GM7UqGQxTcmKk2kycxDqMPhaQBCh37K6/Pzo+8aRFIwAdJ5MogMYJKFQO24qaiSf6peBAtVCiJMV
FGolSyXS1QGjzvVkessWPHbjyWyw8HLYK2T9syMDBG/pEz9leGovNWsGexbdzFgEt3HX3NjacsqP
sg/l45yEj7YRFWb3LDhLf4O/LTnL5tX2GRB66ibgg3WgF87qNx3deusRFnwKLFQ91TJKUncwHvGV
dLveD+QJO4M7hoqCxTTxaBvuThEQg0+iuoXKjA5qMaL4UQWaIDKlfD1oMKrDbUce908CFTXmVfcK
e4wjceI6AU6OIPwxRr+L94LaCofo0RNGW+y4lBJzt9QFGxzyxFNwyXMMRlL8kmaLXXj9sqnfm5rT
OzwPPqKJ3HX0vuowd3E0jFANxA5ulZsXNM8gfDv5a71bHxwIueegagMEBYX2sb71diKYiM1Pc9xN
Hp9XvlXv8l2U6gZWN1UbT8FrBZ8a4WCvpi7g+R2dKnRz4TMpF0izNiwOzNCLm3+yuGhlkEsTtsCX
Hnu5KK7CryYQKDAx/um8XWiMPwzFRum5gIf0sm+808ZUg8gZ4V/15Cp5TIBQjm+omannxsP7cOPb
MVImBBZIDJxUpjsJ7WShiucUsX4p7O+j4m50kDWBOKiV/2RLCEhpIGbYidyHhHHKLSgbUzHim2jJ
LlNhG3DhIGNs5MLkcrp/TWpbc9Z0ur67gzyVJD+kslBrC0kAgeYe9KRR22OvFjxAsRmq/1Cju5jb
xbwWkXCCr83zvr8BP1I2he70OIOuiZQV+yqCZhj+i1uUoKrCd4pSEfI7vjCttgljF8t7VmkuN3gi
vZeMGv1OFamwSaSFaEYlRA4j+uzxm0kZYhBlWli38/VgorSe+nc3X1ajl3hGDHhzjfpidGc0r7K9
yXS4HQNQPnAqwvVG/ICFVOqGM6VSJ/buSPtEvPBUEUovvkeFy3IAWo6Kqkw9Y4C7PaOiYJ91uFEB
m2Cs7IxLc4Vd79QuPRPSSipVZrltWXAYm6zZVPSJiWjg7GA/9nBoUdWDWhWLEDXDRSxAtN/hVVLK
8CoMpcbCJ/ah7ruo7gFs7GmS59fS+0vCFJKzRFUzjENbMCzw27QAl0Hp24wEARBLxmJ8GNy/eBrT
i5sTnp/da/GbMgdc7Dj93r2u0PB6OYpMF/F+h+M9dcUArsRnVAo8EGCkJ6RXB2ectuOWksR9x1VF
toL/NXwb9/wLtWJ6lbLQfhiMJYOC3YHCHTRReF0AFNRb1gUt8dGIW5kCccrIyYi1rKAtExNcL5/c
nqv+G72YTav4skomnpXtgP+MLseD8rbftXLX3STvLA8tZM/Va1i0XWBwHN79ftt7xST9PxTNUqHt
jxD0yelY3zi1df8E/iPbGtL6XZMtnjaYH7o1bgnNQa+KAkC0XNvf+fJR0BwNlulCYk3PN2duDqCq
ik3cFxhr6nGU7gRjT486yAcu5hQOWrWCyIXFAQge+7W8uH5Qdj4S0Lukjt8QqX4yu7/3opp5N282
K+lZ/7PMTexPw0oVQZ7Viqm4H6uIrP0+uDDTsfvUF/FIo/H7rhJd3pUUYAabHeAAgrKawiVePCHe
qyf0jGkdAu8wYCRrEHIPCTy7a8SL4zmPjbSP7pUwAgH0Y8rFEbCOdMDnEXIXCtXWZB532obIVTfL
SJC+1GHDUfbkJSF4UwbDnpnIBCPM4fxQStLeEkYJpkptm7o3YxZPR/wUKj4Y56OsHIN4ZJ2xBXoG
+RhdaoQ4drYclBOz168Nob9j/8hAoiDgFjBz57xc9lAfPA/IurOna6/uyUl1VhqGKkLpLjBHdb3r
xQ+zufYAKRO2Wiv66wwvKQOLbAjSOSpZFApqtFeVjoOOe5W4hIWDFxkyeryaIWsG0zunC6iWszR6
r2bciSl+XmX3SC5OjoKbbU84Enw+KuZXkBkSxybjVALYVtQqClBDjatFkjf7o5gIEQgf8YGA5xBh
jPA7XNGNPFGi+xy1qXKyf7MKtKCrx+BOuDO7U6OxNglTPabjEJA+RCX3PEGWZzmfH7wQV/jz7mXv
1h77RgX5SdolaNsyM0YIhiKYItVpXbFKTVhKnm/rvCqLV2m8lPXsUtOVit4mcM/XYxy9b8r5p0sC
tbNUERYhzWrSVeZwnFaIyAAIqH2I6ec/qUyFjXUu8B9mZ+us+m5fhj+iuENq6/ILx1wiDm7DCifZ
APAXNnaJbB0CHEonoU5MXr8pIt0Ry3EMdGWkABpWG+EmoTvzEXHzL2H81zbkE1CU2e3WFgS/3WYL
XjbKVS+ySowpmmvzE6lF7Ol29BtiVrBJPbvVxv9q9DMSQbBZqWTEBQVAJNdLU8S94zSAzQPszEg1
NswlhNMq8eH1NTozDPYfj+s/9J7v/0o+15HGtRb5rlsGuFwXvIJk+tdEgQp3SIvq6IoKMW8XnHZO
wYZ/YviZWczrwgiC9yxjCtfntkclYVtJ2qFIoBbjwT+B+mu81vjyA1tSY5i84xNHZ87fW51octQn
sHpO7JrIlhV+LzMvHG7etNgAMa1+7If7KbJEjt8tQGEilu6ULCodQd21Kz1nZwXjvflxhYK6Ecy/
HIL28P8a3+N+a/kBEn/LylVIkkUk84+E5YYerqaxwZYUeo2dvfAkl4U0HGO2i6V6kkXaENX8b1CE
BVbIpj9uoyP5e/s/OBh9fH+fYyJFC134QwDtPAakDAfVJFgWeyXwA1uV1XNzZfHDpUuHYA1OiXqL
xRwkZHheqfbHR9KuJ8mMcnmChtByLaUJeMDkPzeQ8CbOFjgZAAlZxR1GMaLnmAQgba/rHrm8NctV
9tagj5AlcXHVjPVImUfWdvRCvvVF41mu+1Riev4TYGpRSMRe3alf/Tfe1syHa1Vc4Syk46yzTxY0
TljP8F3BCu3e9D/X1foEmfk/Lsax+LRSovpuN/D3tNZ0nnIIf/O3tD/TnleuIB96UH7/JlZB2isz
va1HiHE8m9AiXk/vY46Z7PKxWjDFE/2AbP4NoRfbgsB+j4Z0G5Jrhpob7V7P8U9NSwnfEnBgd4Gf
4tg7qSlpnvgwWzUhp/BxIE+yQTiKHKByb/jTdmFTnmn4x+G62mkMgVTO5HSzj9C2WxMdkeAI6XhZ
83zE5wufjnJsD6yGd5giNPGh0/+pbgRgsxUG3Fn93C+wp+BwjlyxLsAdGNOchdAzJAnBkklYZZ23
k7tw8159KTebCykp4suXuPl/paweMgGJsFEWjA+2BNrRAQ7NkoNrjN3lDs0HanMF/Gg6EtFu0dEa
/VTdJqeZgqfFU6pLiJOdm1GWFDlUv1xP3bCbYtRxwZFjqxaN2K/xLdisK+an8Vuzl9SWeERKfjkB
PLo3HxaRgl+wTkaUQoYkLEAVLdJ7+WnjfkFAdZ9u+K4y9229kifQKHyFP03ycd7gTT4Ph1fjgl8v
/KcHV/knjEALrWl2iYx14HSXEbfbeoFNhJ1GSzLZCbMQiHjLhUC7+geWrE/DRby1gmkBU6PWFBY6
5pyG5w560sLyNU1NPH9uFzYEAgoFJL4Whs15KJ0e8WtNkzd+jMkC9GmjrQmkn0/9e3jkxahYg04e
YxDBCa+BoDGT5UVlCCViry+t9+VKW+lR2lHrPv/VhpkdbCMrUsKoqE4KrefJYh0xEegq/+rYCu2p
PVj3N4s9DFUEzSyIBHpz5jDN/UMDPYc4rCPpBq82NsBq/QhgEX35/1LVhf6iiO6RAC4BY3WL2GTi
H/h6H4qTZ5pwSXuw+PBtG2IHSgE+i++dc5hGBYJEKgi9NMYQjo2tLqcpH67396LurPJSVY/agVjO
ZhqrLX+eXHTSxaxgwf7TzsrmG6rPV7QEPxWJy+qUmZ9qr9uyU/s+rLhkOOPdmgeYsW3Bqm7EsgWz
tF33EbFBtZ3YRXMfMyq8vU10nJfJGC+HSGo1pVRBLKPuSr1JdwPUFV7laJLRszTOsZjHGAKSJoET
RsmXMG3eb9Qe1h107ZXgMHLIOD5xNHRvHxUYshtJnMBQzmOjcwTkPmhpkEk9IlW1tRlJv/niaMbQ
1C3lK4bD9NTFBCORAVJz9zLq6c/yNlvyzc3O3zAttT6bUOmKytHnW2wp0qIClMTTDXdzTDi4zVae
/NB53UtmC5uNEbOBzAbMKMI7ygN8C0Y8090tq4CFsDSFl+nzuD/z/Z98rnqOkAw5LQCcP7Qj9IZa
4w0ub3GVAAFr9D4jmBdWq0w1ofKrfeAsZ1OxUoe+f4Mtx8wNuqPLTSJl8TdXfAy7QHLFbNnez3Lw
vg59czuJ2slelJDGMVfZFwzGqfbZss+fi5NqlopHfzYlVEczaoSfmLXZwj4jlHI6TQpVvbjorFFN
EVqu8LA303sxxXfY6tzm8W23+GLuw/FPh+6o+TQQj/SzFlADYbqa8brMcrHqm8eTk6xvUN969Z7T
whoHz2N2C3WsnKLcoJHzOnFlEuG5pu3qKEKG8yAKqCN5gmeq//DCDCOpYCxWPmWWtEm5fostcHAA
GsOmkvgPchO2zVM2gwgO4NvZfu5DrseMDD1XH0LL2IUUz1UhHgYnSstfOCJhB2IM8JJYpwO+ztwe
jzv76LbSfoGa+2A8c+SMlMCBZhglvMV6bLfCM04TPAL5GE9ILj7jqtBztY2DEnL5q4zl5pWoF452
90jw0i3ErnbOrCR+H7jTQaXvO6XGb7mInnpK3Medc8eCeFk9CGooWqFNOrq+KUptZHY8XA3hI/jE
gHOiXRoqcJROpDssd6jFwQ+/MzQ6Xndm4WnJKw4JEl7zt6x24qpnrTiJ0fOodtajog4q46hDWg7q
Un3FXhn5aiHek279fYVZpTLxBaThZrKUoJ4pdJMPbn1sOWSV3CdCswj0MK6qo5Vfg11dKuozkMWN
Z77+BmKi0aSPd7hCkz07dlXN9973WJ+gjiTqg7WNhmx/2ZvJcEvgGyA9a5w5fsSo6k5snHVLPyyZ
CXug0QCJm25V9JwED/45/R/P6hlMxcgzOLXYZQ6zIXPZ/YHjzTuGFRmOlP+fwumTeyk4Jx6ay4d1
lJ+kzo63tE5WV3p9u8SIU2Iw7FckE0KkJ2fK7oFLOEMtxUNCMuwaRUl6tBQBx7/5L7PRYpYd/iCt
/Q4yiF9YwvFg2+ZRoRHcCN8UMXRvtLsjJPQuZe0YYa9N9/YqX9YG1vi2EbO6p9BnHcWE9Omw7PLl
eJVmve7Uh75xA5juyb6U7pN9TqvDhG7US5TkIdzcYlQIgSfBpHxbw/9jD0vswFhzqUyzykeSeKnA
XTMSgmN49TGSiwlaZCm47bcpyAJSIJ899c7O8v8WsOpI80soYViemetJ9vhvTFA4zSh9TNd8zGCf
+f6KCFdcPyWkilRFcvNs59zUa/AHn5PUkv+gNcAeO7/r+GTMoby9Z6pZVGW2O8jFm0HTj2HW0UL7
9y0HDBUkGUbZMJrmnnHxZEWd8ttSH1Va72IePOWxaW3kT/Z8KMnhXxUnDpGrWRqKw/Feke6iNs+W
3GJqpAR6oX54Tj+MN1C50Xb7ETbqbNfmchAb/bCT8pRQoGpg8Epl4TCoGmhzqmUUtlHc/PpnfGgO
tyKsv/mDApQSO8GxWfdcCRYw+twaqjBXX4l2k+2snIlxkDrkHMUfqBQWvVJTQ8x79pacW7XIZbu2
sot/+CEs3I1w27v2mP7Z+lc72pZrmd6ZL+rDYTd/RotrcyC3rMrYUBiCzKNJ/ktLXocjO/JSWuqT
f4cjvbrf3nqVL9i70maOADyrcn/TfOzlz5Q7lBLdbwz7URyV93/74/WZuwrnx10FyU/hmC6iJSm1
XtRbGOAwc/AYv4DYB3EdVYtbo1tvXJ61CZVD4F5H8tkFnC6cPCKt6WgtsaoZwmyrN38l7ky3NOqA
WQN7I2MO/rpuvC0C/Oabe9ZDUMNVZdSlsmpoaTKfn7TFQDK3/5YHVAnHUaF2Q5LW0XxWjzl4l7UX
u+U3/O5ls6avUnDHyXedjklVvyqvJF+8P/FA1nTKALgWf4k99gUxP9gIUTV1C85ism+Uc8CWCGUD
g91zwLiX9OfxAtnODhmdaHVnxhPGUW3Yp4NjSKBFaTSVini8CxQGJw5vYderiNq29cU75npvE+4I
VxNkkPvMA43xTbUAyCy5GAUA04UhsEatlRIeNNzho4aGjt8JsrvtJ39cw9IdJCyt9IWNCJ/df14u
hGq0b2P/BSi3QfatHzYvt9ME67A2Ak7FCM0stTj0OsCFGiNAwenKFQf8W2+YbbnQgxX6eAgoLfAw
JEnaSmQcpF2YQfekbNJExNnYe+z1v2OycNevlM96lCsPrv07DyZkhJZRalJ0tDqonbUCGM7DfDbq
JmGtoUKtPJtiEqHyR7vSO0+xofwt1u+KdRkOTH78RTnFTImrC77H1/Xrz5G0wkbLXMFODXUpruYV
GUyUYd2XV64zVVzwbXbAO9SHZizjezwgz4WDBYK/1LCg7S0Vo/vRnUVMS0dvWJlWW5zeMs3J/UBA
QbZ0xT8j5BSx18F7m4SQd/23qnAWW2MTcxjFvrr2T2KaQ6SEzyM/I7LrxpDuaq0Iq+0MUd+cSapY
q1mj08flGE9ugXlLpLmcPIoDHomGPesce8AJZLlXHy+BrAgLsRKBaaH7obdUbfAnXegYBn/9Yr7r
YK103o6RckTw3fDGg9pqKY6zDoaq4bwIrbRrRmSYT+536dHqI10GyqQUz5i4P0xEQ1MWTNdZa1Nm
YCl9p0ZY5KtE1uvcfPuGfd9Zlb0yphlQVyCCsIsMkkM+143dFxFYdgoVaGN0FTJJhhvswJfVz7Bb
snwY3TEGpxyCtrPHl+bkOytZuW+McQiyADuC0/IhGdqT2eRjJ4fIGW5Mlmte3is8yhvPwk0NM+d8
i2TaPdpZJMrzpkS9k7/L1XlXOfYcaHZnQpzq7nNzatkkDYQo/OZ14PBFEYKz+PpMYXVxfosIRafv
wHjzsLVUcnWedHHEJT5KNGW3eht0ObuCD9k82WYWbPRX2Ovyhp1brhYvth5CBVDc/gk30Dn08l4g
nveJWJEZC3VowXbuiwK1ap0V1ChA6YwHBuvdzbik6ieml/p48zngy+TD9vMQrtQ+OjXxvBzTKmGe
xfSuUCvvoBPWqQaxc6kBj36XxPU9Q8aNWAreNnfUYdZiHgiMS7RPAGt3ULnm/+K8YyM9c4M3iSu0
GIkNCx5zvnJTSTgPOnmkUNE65yK9NLHco1NJNd4wOTPRbM2LtV+Yt+BW1OwLYKkFEJepTbVZf2Eo
3FaFZhoOiFPPb63KipizhMBvrYtf6WDy4CI8medDRQARFBCI78Nzc1O5raK3xoDWQIE/KQOAvjGS
c0RXgu529Bwa0IF5uzq97kaW1ah9jETL4UgJzvq8jf7AS1ZVvqDi5KvhDqqso5Nv3zN0xo9v+hOm
rZYjvSb3LTQGu0I7xvEPhgl6HNSi3ARCtwJ7rholSUPBk8cufNb/24U+jfRJJ/RMzuediPd45b40
Al3UfyfVDVg6RoQVGiJcW0MIbwLVOLSf/6BWLZlmWt58+JPSPuvBXl+XGTxgmVEHfm79IelaoUNt
OXQRAywO0oZMDjTozNz12SnTCwMxvYo+uWQ4LrX6JA54fQWk5C6i0xmfOvhB2BRrZncIkv7shHM6
D+vyJfqafngvDYnoQ0V84e2cLNCEK7aLCLekFxNRDLkL2NVq9cS8Uzki/LhIx1D5jxpEIzYnaaFx
JBzrDuyHzXSmCY/yJ7YDv8ZtqHbEva3gCsnk08lF7zjSiC0IIHsVM1XC7Rtm89s36qFtipawrgcf
2hHEUH+KuHUK3xdcgpZc0/U5zvy4c7xOTOifCjGTMMPeh+ZPg/19W67nEZzG2sGikMtZV2sisZFh
QlVxM4Felfq6WgDQUpPkzRaRfzH74RPhlvsAqGs05YjFQYuHe2/hSbodGJHO7CRnQlqNyeEZKJfv
4rOOFy4bAA7J9R0ghNV3rACJ0gdgh/F7tdc2MqVgEvV0JbRVIyVx3pWy6sGqygsSR6/haw46dotR
FjtgOvUkKQlZ3nq7/7WQlwkP+v7qUqUyiG7eDtrjEqy2BuH3PCqAOUsGkPBngQQSSqI3bTMM9Gao
zPsTvkMoHrMPICN5wJMvHAQGy8Entn9UEz9YuD+CcE7zupdRAkeIXXXsl8TP4AMeIYeeFa69b6cU
T2LJibf5UYbGzAAwdOGK+QTCPm8HhbFoTcaZbQHu8CcJN+kH//zZnENU9JMgjTD5/KINF9eTiq25
yZw51ApmJmB4kC5DUnIW/2H1genFF6RXTXaQG8dicghZhwKYiUhyEJo+wDvPq5RaorWAQ7a7TWVw
/kosmx8vaYGROfIy2YgXMWNspH2Up9HD53sVtU+sTXO34i+7l69P/f7bzb0wr8Rzfs+4ob+5e+3O
Fm6VTmzEyvHjbz16IVd1WhQH0xvx4c1ksE7Lq8ceFDaMVlESVFZf1aGDEQIhILpf8kxeubWVFsyx
idMgiydqdEjZ8avqsxVt8oenmpu1BowsvEZFe9zHxThxTzPF/Xj27hiCj+XT6vEzUF5XcwUAkSq1
DDJIRxH84sj88iD/3LqQ/imFJhOJJNfMqNQUlKCMGhxqTpqoJDp8x5/E4JPlXzHoe2vGlspdQe4k
S+C8WQUrUheaajYIExvafU3CQMfn62hW7WfD6md7x0OfxcgXND+LrwET7zuqpJOT3t8MNPFDXYCZ
DdpXO56kJYyPzc4IBzRPZD6e2ImMSCNy1svENfhFVWjzs9KQZYYe22JB60wOUO3cONoj+WpbKvyP
GdSTXSn75ZsLrBgEIbZXEeJN+4rQeLJNRhViq4fo6sw+Ug2K/E+9pbspYzQSXDskHhtJEYDNnADb
dBAnj3I8xmqpEr2zBD/uObGJCC/COXzVRXwjcKlOS1LPuwnFUVc3CuXYpJeWc8TfLqBd8qXPJduC
6DvJsLjUg1eu9El7p2pYtmtERW7kT1sudccym7cvYh+Jc09qqC3YyvFosCnhhsWYsTvGdOo7JMyQ
890RbLiMUYL5E94x7/YNpKlAx2zZjhKjeyh6x2U+mVlz7Gl5Ev6/Dg+VPPFT6XHzyxsekN459o9k
Qr1pkLAdLjH2JqnEmFwMwdeYv1e7q9cjzOoS6Xs8b8L6nSXhZ3spk5mxU2MDcUoJp37FqDbapOAe
OPEOZY86inPYE6dgRh9/ezfNV946KkXClVY2FmbYn73zq82L5oqvHKri9PB0nq5w/WdZnt+A7GBd
im0azffSuRiXKicfLCBkqsGMUovKCsnZG+8V3D/gShhSXC2gUC26yxmiCZZ+Cl50a0XtfYX5hgmQ
WD0XjJ3QJtzSwDN8WbcHgKmGfWcBM8rHQMi05XilVGRorSZ88DnQDrwwYJywUky96LHOrYqQJ1kp
fkaMRZeeMPyJeOK6g9K2sEIdt1eGUNhoL5yzItuiGEugIRzUP2lIE/ViHZf9E8yX3KbEzrahh9sH
ibAznLDy2n660kLfKTmPfNtEvRXudkOf6eMZ8Sf7Lp4uioguvcMT7w2tBGLofQWacfACxTEDmQhr
xago0GITNzMUrDokN7kcWDOgyE5zk/5VWcEPOvoolM6fHomK5kfX+7Us/Zp8OFhqbzUPuUiWwBKG
aNZG76a16tdkB6OJtOGb/L3GJRvmsZaxdhSWEVXG4bT/yUHEdHcJcb+rpMmALl3ASfWb1v2zXS0P
axijiPYcUg/ZZ31UPb8OQEMcNzoMKk+Dg31ftoVtPmdR3t9DX4s8JUolnt38AlpW6X8DN2qIStD2
XDYoQ4rf6D9DB2e8JtyF5XrYOzhPy4a64E1BjOIUlT7ibl8wj5jHYHAXhi6dY5qCWX5gyffzLgPG
gordF3t0nJRSg4KLrec+lu5jRavgHIPhnjU9FSSRk97+3N6hp7DFanb46awQelP35qUJTFh6Rciv
iFFzHDRJoePOng/52dkSLFPSn87bM+L0oAB0oW0uNHA0y8Al1deaM7zmkhHADXNftKEINJKFEPea
EpKOymR9KUTTR8dFa9tIJbydJwdxYW7w94rOOtgfRxr0kxP6B03kEIyqw/huKPa90ZoYUJo0XQ7Q
9LwBNnluQNcx93kJPbMjCY9z2LrRHy5/VLELK6ReCrmOSm+f2lPbiUr1pGRc05qsgw42NxN5zkTo
Vu2g3sjCfKabyzfKtRrHqBrPs8VtrwpsJ1QNsDlLnmWm3Pj4TZHDMxLivjkb16vE1pt+/1cB5nON
WOJiSSkB5NdSz1IfqfE7WSpV4d/E3t84QqqFu8tNoZyr6BtOpDWyT8YPKZkIkkvQapUHKZnfiYk4
viRhT/dYWWwPYuPJQRMDFb3/nguFno1X8o6rm/UyFYi7LDuAY80PmLuWqJjN2gMuMyXIriHE3LwE
hCBhC5btn0AINNxVJC8wiynWvHST5Em6XvJYM/vYMKfK6y5c6/8+0t39LpCDJbRswK5M/applRmZ
25dswoGJhx9zok1Quw74TwYgjA1wApWANz6r8LyF76CNd+1FCTKFROCB9i+X51Yy1xAvHwmDKQQW
Hhn7+4g63i8pHhY+GyA9OGrNbIF0L8liJC9Zyew+CG0CRYCVCZEdeFYsFy6PlDjjGne5jweTW50i
9I7gmvM08G7F423egh5kMcNeaUjymdRb8WW/dCBb5/0/2+F/N2AsKd76VAFDQFmz9MrLE1zjRwQK
Bs3Bq/CnRKL4JHxD/Lpmh/a6qi/O2L0nSqloaHxpjcdX6L9t1vsMA+IAmOY/EGJ76Izg8FBCsMyN
s0GslXWaFIZD5u9fF8Z/EsAy9G1v80Sq6qvaASWPyDO9jMwpPzS2AU+fo7UbiBp1/imPoB3YW5mP
r+A16SCTDjVrFB8qweDAtainkhmxTCkDqbG44qzg2tge2MPzsmbCOSLDTqoIWZ4eIJGD1+IU3rsx
1qsfETl1ORq42CXHnLJZiMBVT7R0j8rIY9uGfTlBk/O3o4Yqf9O2c/0DmqgXGJJlKVwDz9p/TRU9
sowtgPmqUaD+VeucXQ/GDEKYpsMPV5RXhdg2LpXVJZ63N2Li6S36Rwocu1eXa3iTRLiqIJsBsY2S
c13ohrelSxrCgleemTfOof5SbLEnYAdKK1oa/kJH0EK86pqlmaGLj/XAUO0suwFrm87NSzdjVUl4
mq5lDVgAPYSc7/G902rtEl9v4gBbUgkIPIgyszGtNhigsg0duo4zjDFA1UN+Cbb8lRxuR5uX+sux
EtC8+x55p+W8a/PgyzkNJQ4YvBOx1Ry7nRkDVrgHVMiCl2FZgE2emQAIpuT+Y85p8/iY09bvwnnH
QWhhabJXvFEOUdwl4UCp03xi2inM2LY4/PCa8057xE8Ww2V6UX2kd67UkooLYZodQfk1SNun4JDP
Lj0HiRKXt7nCaU43N3Ek8tSVyQJnukU2Knl46vbmIoCE7mcSNAiR1s9UoHdsBn0b6c3hhji+6OZG
Re617kGU7m1PEcRHUNsGyn33HxoMhzPPw1mJQYrQEdC/yl3/tT5kxJqZ8t3qSyghk6cvlyEe1YG8
InPfOm+BNfJ8eHQRgVi8Yk2S6fLl8VR0tA0n0NiMaFTzI+QFedu7u74DyjwdJRURlNEQ8jj8xVpT
HLjsC+uQS3uTK6H9gsbxkuaCLtXGwdWROZztuH2X2JruY8qU1jUhHkUjFH3knWI6wVAyz9r6u/DS
6+h+R37GivjVCrJbWHAWI6wnWWv2JwZEV7LP45NW801942IQ4QGqRbjD7DFxcYbUWdn7Q3hGCT2Z
QBh82fabTPPceuFibquL966zG9gaww6V/bVXvDgbW7emrc7+Did0y5Jh0J3cPLDCbv7LY3jOHdMk
hO8tTnKFLxkydM7bY/HMq9gUP0WNnpkqYfTh+N3ajn4IR4EEUvtLjcwPRU+yzLFsODkCjYkaNiXB
9p8cc3X6jXDHg97brZIPi1mEb1VeG58aUW20zhtjElRVtwc3Tn19v96G2ffynkdq49n3U/M8zJt7
LA9XGICzPGwEYzzdKFrWhDL/8v62j3lD+0LWg6lhDra1UiYr+EnLIEfO4CJ8yrJ4NJySuS4XGDvT
I5p6yT4CVDFSShV8fXxlNen+gVkNCFeRAlB53zoms0OMyKXJwmAaWZ9pgQDZSJ0+5NtjlkZy1iu6
cD7dKmVYQ7hivi+ZUfavEZMwrFzELrdXow540ErEspfTLSY3nDfYDAGKGHVJ2JCf9kgmA2xiCza3
h0OxbV5eTTAYBVluykBruJm7k4XJ0xqWkkU2gj9aqCwNqopWjWayhr9Z4WA/k1uLWlt+jprg3MAD
DN8LDVP4Fxa/palrNhmttIBJWoKzI1E4m69uXUcW4iaNbtFvmUXW+FxI9wrAS/OiIcR8AcU374mt
m4buaD3HJfHHUJbsuANol+QdOYKIoQmI3gVwe8z57LEYniY8ZeGsAViT/q+lG6RTCmU9NlYWaPr6
u4AfkK9bVBUk51bDn1amIOt+2rrelT5MphplH+yU+UY/oj9A3dj2L9DqVukFTTm1RR7ThT/TN8Bu
9JpFW3+9fMGDL1KL4kDMPclD5i76uQGong1DWQNnLy9OW9NvUJ3/TZPfKMNGJsHvbs62/ar1M4VC
SBvJmBMh13Hb3p6Bir2OZHnhB2nUHnL8hY/u7jPuTTwz1r2GlwN59Cabv/FsKImQEIkRbpBvQVGH
rkLH4pv7oLTTBUYPQeltAC2AH5Dy8e2WdIiWVV8ke3wvcY3whKfQDmnPgEPVaxY5Wf8+Frbl+KSS
EEzyEZbL0HCGKpwzhDDLK+TfHueIpsXW7qdUiHuhfAShfpCMzr7oswG2b9IuWJTpYJBHjVuwsiN/
AI5uC2KWT/bAsYDKsU3aWEaJiRO2Ha2rjPlCEXlWoiJHXcB6ZKYsy3hVGOlyGBe8uElsf9SnCCN+
cCFcNVv1Y94iEzZWCpeUe4OMHwUJSIUjxv2S6OFOmULykOs5vdgBhtiDVhSiS9e/OYZwONy81Zvc
WRUm64CQUsvJgks11eiLsJS/tZu6+z93zHKqn/36foum74CuxYnw21/9UmE3uh+QFomVnWEHwzYb
S7/9Qg36sP4QM5umh8MOVrFPQhrfbg/6IF7PR5qTW1TxQ6q8cuAfSUnAc8HliJjMenlwKOC+MDcs
NPZYasNw2C6Ien+LoL8rrpJjrYHB24p3dtYC3shtk/aRRkRSfFLGU48GpOqD8cdRedfcggYfZCgP
/C2KZZwRBFHOtWiZThMVGMv/0jqM17LW4JSXXC2q66kTpNwtSeF1IBBtOzMqGNzTrlIPgvbB+2TB
xS1kXwl9xxy/Il6yBauri0QeTaYmYVEzH+JjcD2YjfgHIRZZYPAixbiHyx2I4lnHbaLqI027jysW
1M6hrouCFUa1i4JuwSUME/aWYv6jOF6w6nNebME8UWTxqu6QvTIIbwcVBoD2k8p/CqePPHn1f3w2
bCV+qrhvYn/dzEBm/Tkg2HhMfMZGqGP9EGWEGjp6Jk650lkA3y/IMtsVYTgeN9YQDRPkpCSDVxOw
xMDZo0aZ4rXjJy5c8vKKQM48Pya0E13ZdMWwD+2vFA4kB1x1weARLgFw1O1coIVHCFw/MMTtTAKb
UNUDB2d2jJ1Ay/PzrFOsnPelY1kjOqz6QbQHIAKuOGKvrciqhvp0E0vrO+WRddPth0sT0PrimZH6
cSKpyoRVps368MpSELSa6DsyVDBF2gCEtiW8WQb8s4+OC+zWnerbWzsfx/nMQ4IUtJzhLzEQknzn
kUBrk1aofGHOUN538CNT4xMnt3oXbnxm3+bBywbyi1O9ZjNZpPbrusPVTWNqhkgGShhIxaksIB98
gMzbDgmyZurZdBlZa8o39++D1qA8INiMamVfijAGVi6bpgelSJ6B4oXCrnFMNpqhqxyTU6I5F2XQ
S7laXKdsJBA0uaDek6NsD5YTOPrlVQ3sE3bR6UQ+0YQ98B+cjfToVQi/i9stMiBWDMlI2j0Z2DNR
eKp7JKbJ+dC6VBCYJPxu8Fo+2Edq5ZpD2cMywZhGYHu4vErgCzFhCe0v+TEiZiJ80PlLDB3QHuVo
PeFeBVpUl1gcAZ1EwJwVQXPfjaaJTn0LhFHv8uUis15+bFey6LpGIKX3dtlrqnhWeBV6vDH9BB7e
CTfTnGqsBHvGsY8T5WUqYFB6fflCP1XfI/Zn2stRMQhsZecUhFO7OWyCQ6q+PbzLzs8SqeIcFcXe
8clFztRslp5ZRbDMZXiZ+6V9j7dDJnxDMdQU+zZlKGMAR7odZWOMD/g6A1b71rSAlXDkerG1vHcw
7wDgoYpIDW7pfKX4Si49TOfZsAOLcsqN5jaPq+n6C8BTZFXr3AbvX5KK4KXc70JP2ozeS+9nPU+8
aMDGDnXeV4K2ADKZKpSazZHiifR2RRbESXpX2YbKEDoEr4C5Wi6mSmisNcE+N6L/C+v04oDOm/Uy
G4LK2kxTLS4/ejHIKSfvgbF1iDrbtjMsHrlTJKNq+fcHM3oztIyzOpONU2SdhtCborC7enoLWyug
I2bXpG/JKey9XT5m1UzkQwgxgDDPhPG8tKYI8dm4LsWWoeS7350/4i6EAn7m2uGQDsC9IOVM6gDB
ELdCNkXBcXOPXcv26/qWSXKJIuaBvLSqZV4ypJdgR5kQdmix8csAX70FPxQPsLGwW9XExu+b6j2d
iYaOsjf1KaVeSMdU5eepMBJWHgH6VnCF4tUOdLgElf57NzL7NC5a5TsSukE09FzIgqSf2yjK+IuU
9qU54kZs89n6h8nvtFgnPH3f9n+B5/H0I41m4Toz1X1+pJX273pORLcxtelAAXREPK/UHggwSuIF
pXFlETuanwS53IXKXOciuc6Yd5r4o7rZiXeQjxacCdNlRLQtf+MrFjNMPLk4CktuPAgF6mmyD827
4+g0XvqL0eERi0pNA6AMjJ4j+AtaHAxiu+9uOssmkymgVBPNqPllgeukkbouhk5E7FWzr4J/gowL
Z+HeCqCVPcZw7Xkfd5XMsA30X2EkPApGPgaJAnbxPLDWx9MTAoYhY5eYZC56jNNeULtOxEy5auhV
wyVZ1TG0JdOHsQadeuriq969yBMrFQM2r1n50x96l+LYX/vXnLzsA+3Q5oG2GX+NGk1AMDDYp9eO
HJv/xMILLmdKJZkfZIJH7I9U8yhraVG3J9NcLs7bRlJZiK4Z9CHjzE1S32xuTNpVbN/vp+IEXCxz
PuEQSh8viNCVGJ7dfs3Sa6JU8HtIi7JwvgrCVywMlJxHqd6K7cS7G0rrbjP5JbAoMxXTJs9htOGv
QPkkJSUQcMXSRbMdXuuWBdiADn2M9WMFH641Sip+yAXy+DjEbiaXvzeILUiKeV+gkQKIQp3zfO7+
NMIcY0FnSM1PM1+xa9BO2sWkt8BRt8sOwxggujwbTDqmLHkB1JSF75dfeAxT4uRBQ5B7OgVImESs
Rhc5uljAB5JTT4TWOgZhfYnjJmgJuWyE6v1rP16gV3NwXPSozmA0oNs/e+FYZMGV+YDRW/w8Sbll
WQzvA1+XhY3HAGr6LH9fQqb3SQcZcf8BO/ABH1eL3fSP3ja+owJBPGL8yZ6f9ucoD8Wa0zlHbT3o
W51tkF19Qkn1x8/GbM7J5bz6qj6MDl2qsL3rYjOMWrZyUEOL/XCTgJMezoAAXT+K+RtIaXbMmn39
Uy8wRF5XbmRYCAcGqZtby28ac7eABlrElaNGtlDWNIdvn+c77UiPF3FiZe7Z8NV1gMj9nm4AHDvv
SGWC9Of2HT4QAnMFwn7BZlc58fKvOdF4jPtgkLPXPQ5RyIk54KmFSPrN6heqcwrzndGmt/TzF7cb
MRAVi4cJ1oenejIqWWYZ7HTdLq09oWE2fjBODVfRmYIrbowgViGbj/JnPVvZJFjC5Kvn4ggZKn1R
Pskqk1aGkCyzL9ddXBXBkGZHTyRG233qvGny7ShOL6+PsMyPQ3s+MGL17mQwxS15cjOWXDxlBIUP
q1HmlWhkRyRDDPXHyVNNcHzkHrIKTyyXEPC4JNJhdkN6rXO58VqZlaQAlkKk0hRhA8wJ0jU686Vb
2dQrJ5EtmPuYwZgXxSj44eo7jjxElt7sIgedM0oMGDsvCwOVH1GK8dwTvDmGJA+4/42O4YBySe4U
Pyl/CeTXZfVRr/SLUk5rzuf0FQC94A3zlGcl5NdKDNg8l/GLV47Zct216hsNcAsXZdKe297QnNYm
7kqIWQ+BLA04nx5BBF4i+HxM9phl29Q5Qz93OUdzODrTaAuRcmlQp6cu1HzOr+RtS3UnLyRZ6a3o
It6GH0jtPY+clWcesfCWEB6lRFaOOJryDVMWh34SqS+kRXHkJB1izElrMaI25ZoCI7rjAx4Gcb7q
rlVVg1D8TXrBQhk6qnI16wKbacr14I5jG5nS8Adl0SnxwlSqgnUPp5dB6gcs46DN2IEnZOevUDAb
CkiqQdu1MVNCO4pFr0gWBEt4eh62vK3/e/3xCeGGAyM2WR9Rxcu9SXI6296mlB+WoORcdwYWUSwU
l6lHDsYLxKZVrc0nzXCIqN2L8OTUWd89tcQO02k5Lss2p43Rz4sjz6/Hb1XidU/gKc3d4y0RYWPo
uLAxO4xzwFtqqX7zx2X8vKsHVHLH4m+VWkMPTfZhS172ZGUsBbi6qZ6htdqZboEWdHnnQbxTp7iz
DM5xkRc9b759IKY3q7RsKAGrJJq3dP0j1L0nRPBB1tmIGk0Hc+tHpzmi/NLzKwP0Q6yVjiKABcJI
9SV+eT5Y712oczL3vkCZg7t1N76bt6F0dXn+6NCjw7kiSOEOcpGKFV1jZuwcUVw8Ma005iR6UTIm
Q7GB+sOPAWe408G2zk/wwoCNCcwOjTiFoTfvNgcjk7WS3bj7GxPHzR4Zi/Wa8zLYB+3XkW2oXIxu
0/lTyBQawfBWmOTYnYotmFjOFNaUnETJ3ghOfhmBrU302/5JLUfWR/1Zp5FFV4zxB4sExrid7dpi
lx3CwrjcF+PLqPhRejZiluw+WbgeW3seBqagHliX/mkDUn/5EyyFv1ejddQjnFktP3hvKG73RDCe
5G2x/ZxOaePeh7Jc1pyK9KyGTFxS1OckLtpb06LA3wbEHn3dqyJjV5PzYmlwRDbh+Q2yjlzwltMF
c7bf063/6taw+hrZG3n7gvuUrcc1ZOH3bSuk3pKGUJeoT1YdwQ8xaduC/wbj8uEJZRGHBYf0Bio+
idIDIEsYC9tW2ayyObm1zKBfwgeFS2u1pH4HPPixcsy3KFbiAkt+HDecxj1tpVR4vhxKkfGkKUS4
rRPXqZXr1K5Q7fVgxAFphFNz53vh1gKV/PcHWIf9ah7XwH9RUyuYG2tuxCjmIWjLACZKUFqWV0I6
suCRj7ru9hkDIMHHMJ0DAaqUnjHNu9V9ar57Z8tc28O0KImogZKVyfg6wcEjcVONQNQF/qLlFHAC
bXCSCmHQQ/n76zSXGHIq7KBQ32pwzdcVwXcBBYejTAu/3V3W2XObZAeUcevP+nOF31nY85Y1UJg7
YT9r7UoL7/tCa6IM5t60x8e0yzxQ1OadmikNH3TS7DXIo1h+QO+GFTVFMip/z0cS5k5b8w7e6o07
RKsJQLeDSqYw/xmRRHcQ1qb2hfG8VYstnWgrMP/U4u+pfmcQMivfh8Bvpkl4IIxA7nSLiqBkSUCA
qDLhluRYNn2sbN4xTG3hEM3TeFi+WizV2MKLpdmCQn/zuuhpZVtZv0DM+nKNY5upssi+AK6ewglU
DJmosYRbJ1hpawomQKhefjAR0LA8mPiSs+vuvBdonqydqZjGvZIR4s+n9qZLQL108wYf1gJMjKG+
E+Kcj+0fBdTytTLk7zAuAjNOXzFBC4iLhhR8V0Bnt1cGITsjDfL3XmpbBwoO2RG0bJfoif+pnCpq
Z5/i3uUD7k5GKgNKpJpmpZLJeSHikbSfn9C4QeCRNv/lHCoPPuwFJy19gcFx9Gvcqj99E9fav2KU
Zis2Wy8AM+UCJK4fc0W9O+4GbXiV3yIno201kAZGLSJyLrwTaW1P4ifm1ljIv+6xPefXdVfKLoKn
gVuUz0dhMZbxvVaDk6+FYcrJ5ryd675qZGbPij3uPkS7m3jW0urSzmpQmmruo9j18fKjZbfh3BOa
sDjSMQMCEvM4dz0lyPvyCwH/8ooUxhQBAsxEO6dRHLgFVHoQ1N+6U46qKyWLuwUDpMCuNDkY0r2q
G+7lRyJCHlTSiFG9gZ6ftNGuXvxIBGnAne+96gdvLwgYOyE0+VrMuydSSyrE0rekzT9mLsg2pNAb
PxZrdkKdtoBL11an/RTHnx/RnYzF8feV4yz+gGZEa4Q9/b93jcVf9gzS2rBssVIRK+wtJWP+Mys2
dhMK7urRWoggCn68WQDtZdUffZHWJkv3bC6JBWXqm0z5KCN9hNTcq99BXTyV8ioOEIWW7yh++0A4
V1+STSQugQshJniuX7Dj6IhYOV8QcREGrH/YqSCqB7/4FW7NHWwBNULJjxoerGr39tAQxBxVN+Ws
ZMr6JhN9blJzUz4rcwN+Fo2O8Nq6VaLIlETohJFIv6siqW8ad1hHVfVg0oRRtrmgkwsBVMSlFm8T
QMMpj2r5Eet7w7uOg38ljOaYBAhTuKE5eyS/Yw7HpoH2upmWOOmUmmgHdEZsAIkNVbJPrRXu5M6p
4CbsUP/LLaQICOa9Tnsw8VUk+xrwRyfVasNRniHWPkiMWrrrlEAln2b6D3Y92+uw9CuhxGkxCM6c
9rJkrDLAZn3KecRurKO6KhAQFyh4SYbl/3zVCMf50a2Qhxi0e3Wn5GEXo3ysVfT/VhUfC556K8rb
Crrauo1fsnEEadMOhsJIp7YVxLOvzB9ioqIX2GqRG9aiaZQzOosgEQRlHevLf947Gqb2OfDlbQxC
xRSRaBA1BeBcZ3vOpq0EEiYlBO2jEYNkaFHa6GkDzhyduvitNU7cByruATyp2IylQ7bzKh5yuZRo
4LtJ0bTS8kS9QQL+FiCxUMIeUCBcIarFOE6bqV/PPm/I9FNPWpjoU/bNd7VVsC/bGSxqx+CpqL7x
fx6yT1rNW4hsr7cxKg7D3Cegc/oX1abPd40/IIhtIwIP4pB0WHO5ZhnEIPFyZ2BEAp55vocVPPt/
xN2xTmvo2FXJZTw08f0GD1IysjG6BcPccFZ8AhMbqx7tucX0y08mWP4Xfdq1654HO7wvKFasRH4x
YhRzUnbzYYFGBbrVLVSR1adKtNob+Q2uD7XClunaAJhb5N75vI58aoHmWbIF9GVXQ5dYm8ppETte
aHft5vy7woe0vPTWMN/V7CI6diT1mlvd4WeoAF3OgiTeZ70CQcMTr0hMgGTmPY7JmY0tPSkmipw0
I/EHkbmNRqtVVuFm5SDuEoWMcgM95+hX/UlmdZZIicbcTsqghWVRhlepnR7IRFdHPXNlTKUTxftK
UuOvjGcTldwR7KwgYksWnnqj/RCPzSyjzaJuN8QbhGmMwhm/oW67mZKaorUEoM6181SxFBkOFVz0
3hHJ+77fhxUMQtOXOqsKxaQbgXZH5j6Fjv0V2KeTRp6PcFybk5M7UG//tl4RjiC+FJSltz7Ytvfd
dvLAM+uls+peS+wVdC8RR0E4OwnQzTW02vSEEXkqfKWPzlT0wqNP19QE5zFuzsL4Y6exan25TNbL
PS1vN13DHJvNKHl108T6JpgHRyjQEKe4G8k50qWxng0Qqs87rX39T6eCgy5NYFnqDwoPj0hKmfcc
h7zwH/2dm0vyjbYW2YYs3IOE/fhXOoy+GEqdyE9aF5c3sskE4/APoQkiIQ72u99LbnJRIylWY35x
rbn2xTFTXVvRRxsDgxHt+g3tDvpna6D2wTfDkSga6Q9wTtbIOMOeK3eNlAhOqDEy8MAiBZ/kHU35
E7bBMKLGrWAnY+5x/tyfX8czVSz/NYCQzcpEt4kMSdtWvgcT77eZTd8IXJmjGAjVlSBg45l0F9UP
9DrlJbfRPF2qjYu6SbTFFjO1OxZcwrOCPsvCsTxu9vGya0RrujFUjTx8hxY3BCVPJYw/kZLFhexq
hfqlAmpFxLSWHGbt+Clkg8mJHZ+/cE1WyrLUb/jrVM6O4xC+bt5/yfsPr4yTR/HDHHigtF0bSaoy
tJJWMjTlo52ZbofpenZIwDxbpH03pdwZw0yeTOxOpqp9D0RGUkj82IIvUG88WIUj7zkrFky1o0U4
ThWgEYqF/17zu59j3WlhkfDaIhSwSe/JeahzMw8uILc8kqN4smZr2WfVtYdMdwAES6vCSj+aH2x/
qtl0NnnbMUgyXQ4WKy6zfzHT9lvncOvgx1OHgN3yCikOFeV6eMo1f2Tnmd4Op4RGKS6ZU0BKPQ/K
hng8ZTRBhtnwNz/X+6UqoLxWBngxO2rm39IJXLiHMS/9zh8GtZexgwr5dJn5YHL7bto1NFP3VOvf
6IdZE1nf8PL1EAi1f2numcdiLmsQgbmZCdEwUrGbmB1ju/wQT9FfIAqQA2Cgvgb6b4x3SJze3nhe
pE344V9/+j9n8cz2tcPHDbFIXo08pyrTBgX2aC/PIbqAsv0VENSykv48JA8Khq5+AKg1xwQzaIHg
fX9jXh9ZqP6SnlaLsAsUJtVHd/63YQGyG3ZJ4d4sln0DDlvFzaFQzWDuih8SaIoDAhsecFzkt3M9
mKHlpZatAc7BHpF8++TlMqLiHvt6uvc8ic5AdLzNNfVJUXqDt6CdaaCrDlkw41hK80SyNeTgnnAD
SsHzdI0x2+pzwBFpkwUKkqP0Mpw7qAjbntUjyHJO3YAM/rA6itD+K3gMTk6Z3D46cs9LPH8TvsTR
k7PpTmoRSbLTw2SdCTdH/Bn+TrZggJz366XWdim4f0DKlBsv4A9omefqTTz1JRatcdW9wPKup7I0
EjtJG6S3qdOQzhGz4v/h/MgZTqm30fBC4z++41TqxPTeD1OFPaGaXISsdT2WwLySkk1HOr0OHs5N
HDT0bKfAPTFDja1+mK8LCuaop5W3x8hkCrlL7wnMUEQp5xwKyoTILZsmm4MDciNx82b7kqRpjXZd
DqE6oy+HltzIQvEqN/Gkz4mO0dXauAvwelBgI+WT5PPXtxfKD8rC0hpxAdL5zMSg/S5qXqnwkVpK
OLf+G42gILwbRkVsTcH+SvB+rORy3zSJcu+3ud5r1t6P92zDEJEOYWLlPNZu4fJy2EV9VX0rqsoD
qwbTW5AEF4SWA1ZvYJ5gUQHDhntwGunkX7fNVcW6hU31bjJRybWQr9isFwMT70PmzxeB0ORBlXLo
z6QBdtGp4Vu4dnuct/d0eia1CkIgd5hIUaF4XeAk+XeELviT9OKu1UoUOEi5iNr6s/7IsrxNChFc
NO1da35apZ1m78X7vgoc7Tg5dsC3In1n34qfp5MJUdKL2T/dUOv8alewwJIhJ/9FlJvXOwYmxBJi
jyWmQ4tQfYsEYZhi1J0Ba/pJG1FbY1rXHvagW3DZe2S8tTnWtYahE6Lk1gi0HiO1Nkp1b5PZOGjc
RzIr2Bo5nOH2/PzLGMFpHGkeRQd5y9lmkQeupccPFFPxl9UxslkS1Nj7jSyZ/0ePLn98xCy+Ldqg
wolWBqfH9ACSZu4MWOuXTnbyw3rjk88WD4HTd/2+UB0zvuFzppH4ZtC7nTfwxpIWbyveCrum2Ugz
5kZJ29bhUFXS0U7n7KImrCkrdYgHfCRwaldWdavvWYUTfzxtd7+GsvQSwJ63Go6t4ZSxyyQ/fcKA
sUsWpBkeRRl6LNge4STmYSfYnUS4fYY06arwG+EvEGm1kI7ceWxfTM7mXkM7UE7gdMw4pGQ9rkUV
xEs1gx9jhQsvJn4aAwZpp+sedlT/42wNLOv64WVbQFLdKK4DZCtQQmo7fczDsTAcIeXdA63iryFU
bNH0pXcbtyin0qXD3Z8Z3mD1cT6izcJNCTQ94IwjqO2c43TXYLfpDzhDu1cl1zLjkG5XBaxpfYlZ
/GvpLw3ocV7aXiHjY7yDj3n4d4fG5sOaDYyVAyYX4f7xNIauu0EMkAuQHATaeAk6tvRZrxNOA+rC
h0MIk6dn8poqXSx9b38XCcQ+ovhYdhbCrHg0pj6As7e/Bi8FratkNBFVWWqQ5P/0fAYBUTlUt4dI
HCVjdQNP2+AfXmM1jfW/tnGm8gTsRO8U3oEG9Esgc/6yZxSYWzbhGhOwIWncOtwD6HvDDMJuNqfo
x1U/ACi91ZOhhdyXO+o+WVqH8GBO3o+2aSLiIoaGSYYCZaEb1SARyobWDQxSMqXrOcfAz/2Co8BB
s07ukElPyDazzdy0+wwusxPSmJyvKxP2/E/eHB6Xsz756qRJqse8WcRFxlA3Mdm7ennCKAdJATUe
C0TaDd/CCphQXQd4vyP4YTZcK11+r7n5pAWZZvxPY4tkAYmDWoDo+avFPUJbEJuiVgVyR3sunw6Z
B4fFaMYtu8WKfvPmAF9yQ3s1f0TJ1/v4tk/y6oTlVTpan+0UKqvlEWTOLPfJRTvv7q11tZrVaT4/
xcCPDQjIzGHlSevMY4iBZG58OFFQbXm5sgVdyrlTvNbmoNLQ4ILesDyhLa4jSL+YsZJmQDHt/jM0
XsRzvmB1ZX3n/qLrCe8ko0MxSpl8GgNQfZi/9+PYGoOht93aGjgqsxtTxry9meXYtQYe6lSicUkB
Bzwu8lH0sxoMrRHgUwadE56v0AW2AzB/90NfYDJp+cYpi05axz3UuNQIn/nzSsNtxJ6AfnR/UcFC
CLGRzj32TdsuM33eOvEFu9ZE4STWlgD/k39o61zl7O8741+5dmMOLZXSN73eFLU9YkHVxx3hT4qR
xzZ2GQrAMijUWEn+VLJiYmRvZLTtPvXj/w61GUtOJX6L1wQSj5JZYltyVjBRLv75UzbawmEprB+i
OqxrkY/5+2BSScA8ve9+3kleeMU5Ax1GJLWqzjbT5sbA/wZAGwWrurfK0kCaeOoRgRthX7TFlhwK
v2kCRrfyI4J966KKB8hSJSmhjNYEG6Ahk3Ofziy9KXp5aeIGTGleQvgPr4wchzU9Nrl8SmhFsr5a
O1riTe93yri9qlm8T0FoXj6gf13AccIiJ2muUPj9gBOHSvSfCtL2/KuqZwrpoCPmyikwgP/6Y6IP
F+W2Dvob8RsCrg/pJNsZGWrVEoQEuT5kji67lIOX8cxSnkq90Yh5nFhdLhnUgEdDUfOhI35kSHhJ
QG3EzpGEnuEH16KjprFQN1qEROekl5cMHngzxQ3/ZggTCdaRyHfPFZEpUU8xVmcbKhWOuoMg3lqN
4FOM+GWF3rz0BB9rREPdMHMd8ny2IKwWkA6fAJRF1r1pdiNqT5TM8ZuHeaQ+xVWeVHg6i7VXpQdC
0b1K6SwiGeNLDBfrWEaghCA8BK7yDVN//Q0hAZYNmvzKiif2H0w7hgijkhlxcf0UEQiUBs2MsEQm
wiSZzZfifLgTf1Zns0EA/JsJXpFbBP0jNf1rgvfruIrQAWpvivSZSzBSiZJAg059EzacjviHGjJq
InUGDszP6zne1vv9r0kURDqxKmKS3kPa+u5JwByNsOl/Nl6x4isGt4vGsfjtJruXp8kCkUgNii24
uAHQJMlVjiNJfnQR3Kj7Uqpw5JGAl/shPqOZ4Ggw1FUkAjY/Y/MTY7hOJj6HcdSoLsMskfCrpGq+
4mjMkZiuYmldCqzH+AoCnXnDIOAYjFLWkjCZy2+EoZr/TsTeM639mqGXnm3ghg//6TwLiyrDJKI8
Fh6rrhve2HVvA9k8lT2lrg5tW6V1Fp1oKML3BESUd7vpbWxXN0OdmQ3ySFb9OdBw1vG5u9Y8wXna
FKobZm1zJSBSzNcKvq/JEMPglKxvixZgU9nRpW1nQnHZwj1LNffvI4esegFSKh09Lzbz/ELcBJBG
hesVePF7WHj1OGJ+KAw6fjoNXAuCJqywLj6p7z4fOxhBSZn52AOtdpGxta5yyGRFf7FB2QBLxhoH
oPMKbD4eOXSx9W6eRTj1oJIUP92BhEkYN19/cxJANY5t5c+y9Wxue5VFP5FCKNma9B85/pyydcZA
DlHykT+198EeZtCm5Jx2LJKM9jDaE4MyFD11IgzSFXrzOy/uv5cup9p1XN8AvYwEiItNi18fwRqd
ihIhBzEp8DOmsMTZ27TX4Hh28E58AlsduhArZyR0yb8LIJceC2unqN9r8nI940WBNOCbH0+eOucJ
ZJzokMHv0nf3u+NTnnRpvbOdq175RKc3ZPmbjeFCUMWCDPo35Oakb8IyQcFfWvMNvBFhscmp3hk4
A5fveXVdnIQ3r5qH4/XnVIUW42MDUSPp6qY2582iuftCQo0HVy+tmGa/k9IvjO0y1/MgQnXR9lRZ
6mJ8MOvWQSwPOSrhKEdktuczLT/TSMFZ+k6Gf/H2OiwR7y3+J2RVG60O1vZhtpSonImhW4b9QDWL
tfW0Yzm/G/CkV/6Q8ZRa4/Yd2aNxvv59NHq4TlxW/d+o8zGiHA0A1BlKJ46GJP+CVVUWA1WX19gb
hmTWXX27Na4hjBQRXCkDFmYCrGBnZmV86QIQRhBtLG+Sl1DBue6UoALSyde/L4GE7ON5HKSfj4lq
Ocx9ROviCwwkvUKvNNIGFMXWNmaD/yggFmTqjip+ykwjuRnwhD3FqqUGcAWo5nuoSzJrwiMLBJyh
yao6Oy14XRAjjRNr15orFm8XHIAc8nes3F1RweAHJZRbw8sF95/qjvwmFqwpDfSr7f/g/38uaY9x
vMH7IQoDWVL5NWINQnhbs4LYUKDpM3kLGajvLzX2VdqyoCeNN6LUumxTVyhtwo1cHS088tpo29U/
ITtaZsw/C5pyra7Cp6V3MBMpGTYWHQiQ0wv6tFp87kAJrpJ2O79KbgG5HNPhe/f2vKIzq7lfaBCx
iCccYJg+KmlRFhd0jCIsbtlD3LIBivtc9a6zNUsvBmP/YO/cdaL6RI5a2mhFlGEroW9/BKAfiKt1
2m2Wi2mSt1sBuLbDVX2xljdQeZdIbStNZcBC0iXi01v8WNENtgOZhWHlxxbOne2NR2166345I/DG
kDDM2wfK5UZ2fU6DYtKy2klUde4i+655cZGVMhmshIGaHMfDmRCczFJvCJdmRxNvwOJKvtI0/sy2
tWva2AeX6kzqwqtuX/8aW6I6wmxtvvIWxTH3jGIU6/boQ3asoNqHiVecwPnaaX1OxvoXXIbvW1CL
K0brd9Gc+6ZOlChGdTUpE9xsfRuJ8RDodxzpnf4w2q9FP13KyF9Y8Ibry940VHV7C4ryGf8Xu69z
CQWpSabEDxigLuj5pm629X/HUtX/qJhz+fXpUkp+gUfmZPiRBsJWxOwpBXDmFVDgf5YOislpfrv6
Z/4f0aenDukQ2XWoNFBO1RVTIh+8JX9aUQjApbq0kQpCC2TAWvbNtmw8LhTmdHz1SBi1KvjnSje9
t5v//Un1mhPeJY5FVk7PAG4HmS8n6lqpyUAslyjf7vLABRCIYl4gCGcHi89enves6LUkUxwKkvvz
9wi9gI+tlJhXISpZoYXaW0nsFOsEfS15zGLfgnq9TyXK9opqaXVS17u4SGIO9JXcJTYTG3wIyg9K
3Y8IEUMLmxFZZZq1htdWDNRkYS5HpiMpNVdGaThqJIn0/XjAk3XCP5VTSLNxGwFLtowZshBZ6b5l
deBH9skZcfi2l0gIdfYKI3EPRH18kSZ9PZibezSR4hQfKmnSoXyj/P59Kzg5XQEggZ3gKdwflCjm
1mfLC03enanNYr1BFEJPn1kJsdIJn5OtB3ZhBfegJRPZr/3qur0IfPzJyZmeWHoo3bc/zeRYjyw/
zuboCKZMkSmE+A/8WjyBrDTiAyyQhllXKmg9I/QU3n89ex0BFlXYmnd6FHm67PQeghlW60Z0SeDc
mHIbuGGAlij+ihIheu+eJ1nl7XWXhKuEEDyG2PE9JWJzguwXbN9I5+34ShRNCI35RCwizZCFPV1c
+9EBxhBo/jRY/ayz6PUpp9SXJJReYQRWUGdLQwqq8D9/dxxNcA5WUzQPgBkPjJBowsjaQLp9QQ4g
qCuAgb5MQ87Srq5iuaPBd7ynh+QjtP8glzLQ0Q5B8hJATDOwmStvaGaan8qECrbV2zhurVaBUgjp
t95KlTGSnKrsGWuIdnZEHSUPp8AiNOEHpgDq1jjQcw/Ykvv1G0+TQpmuGU1CP166SmVUA6jUFYsW
yVSfXwucBjiYBflS1J8TE2+jcQoHcKBnUFxaR9EhvUGOtgnYjHw2sfpgUn02OUyvjXPwkM1+JetM
flWLvB/bzfhyWPEx3JQ8tnNkzAwPUjsspfeDtc+bjbC9326yCOifqg0UqqWxhnWJmWkXWxtJdDvo
TtZDHPHJwNfUKshXwrHbxFfR7Nejx8TlqsHPVAAajrFVEQR8S00bMmQ1abUSjdlbPHO/8koXfh/0
ckI5TwsDd9Xbcq0/n+SniRCddiGDBdcdKqnEsbie5ybF8HoerkToKjyB8gyT+SBKErVmDAysRJUn
CavGJrKqJy6HMCGdZ5tKi2If8ihE7/k7sFR4rTS3VAoHHPw/44VudgqdjXf97/5ZVtZpctvsr6yP
LTA3Cf6lH+JcRWaPlJb28VKVC3sEgOl/1HLQVvpAPnyFx5mLYD9vV2J1qTb2qw8ZvJyqltl9OmAe
vrD2VgDddaKciKQc0VvX+ecgJqc0/VTMQqdTom83RF9p4uJK5C2OkOTQflsT7WzG9WXDM5QQNKW/
J1jMOD6ZdYF4bdbiPhyFPKOhIWfMz54tyTJDM+ycCNCMckwdmLNu2XTuHGhCUInuYGOnS1Uukx/i
uoinNBfrRzJOu00Rqsy3bMtTs/i3D5CY9trm3dBUkykeeWE8NKmIUAoDrsm8tp7Wajyv9WF5UNIc
nqSfTIVaTXtaPd3M9OPPNckhpxeSX7JRNThlOxiKIssP32irg+9MYCVaDAJ1XQsALcLTioPMGR1I
EHPXS843r2E5I4prwmqXRBpfBfWW6/llvPfFKbskzoGvwjn1720zk+jXaz32vDJv2V8xIMOUG1yu
iPcqinUHSlsNsplKAfBbAzyUaxJBOaLU3zGfZt/M9uQ2bYK+0X2g9BdV4I1isN260lZphnXf/iOs
he2jqxpIyyAaSa9ACq1s8AP49+MtiVpunlplmaqPKfwX6fF1MYf2rXnGSaiYHA2i5m0SzhAOI4qV
K57/PrzVT/zwACjvFOQ7xcXBDQ0g5WijxMVHKhp1KcUuTr82FbNSQoAnCPI7Uc17BRxWJWfQvDA3
+/gi0fHjCcf7ZqeEAR+9f3qHJaqjimMDfce5K1YgVOukSuXy2mvqPTCTLnPVEG+PEwtCb4JrHCkf
5Hn1q8YN25Aq9ThgIY7/fMhbNhIxmViWmHnRywoZXnJ+uTy5Qk5P3Qb4qIYLAzrEF5Ev/Q5BNNQD
ckxSPDBWjJsNrY3sQyDZB/qqSqS1p5pKaKlnByDn7uLC3XbDv/vzVfZBshHTiPi2JVnB9Hf5DZW8
ury3gILzwfEnBbg7nmDOflqH77U6riWxTjFoU0HrpD807ly54bUNTzZvMZaXRNPlCp8fZpDyYQIT
sQn34eLjVL1Yw5RL7hykmGRAKMmRbnVjm/Rnrgpe6WMazqH4JINz45C/d8Wao99yflNI/ggCK4TK
pjMLgkIl3Zvc8lCEGCDS5qWlFxjIwatMRHPgs6hwvGFHMYzZzdD1RthTsCEYHG16cyB5dnZ1yc75
4Hp9jOCMxkh+d4+eNmt8Ztkt/v68GjuO9IzySQ7/qAGu5WAfBTE7ks0fVBDPPlE+e21VQkRPt6ZW
aEFwcq0pagSKK/eju/QN/jn30Uh8zezDpFV2zzERYPmKsNLZC6DzIa4lX+7gkm7H5CnqSnsQHCY6
n8cWgvOffMw4mgLP58u5LJq0D+EyTf5zn8IgFhbH4PyifCjse4R7tI902+W8IAzw+Px0pDSnpqTf
ZRhsJZoQElDvhcCSsXRQmoX043KR1K/TodHHMA68CzhuWDtFJiRiVYpdlXuHEgEwGuXtexJfirSh
LrHf/iKgiMdpXjidoUKjqy3TFztLrtTifR1c1IVYbdY5fUQoj6HcYGE07xma+3czOF6SAZd9U7QL
uPmEhqhTt7vdQcc+jDiAPGXjyoGrhEgT7wwgVqBBF2UWusNRt88ICdGP18cTJQuAALRedBMGuRJX
OMDVw2F9SKSw67EkmT6qe2ZxXDxGPk8l/d2FIgWfn+eHAn4fy2WeXNvXbISUf4UDzSVttyHSBt5Q
SQdQ0eQpgjr/dgTGJ2q05cDYlJiaxNtozOdU+9nR8OV3P6e67GDTkGPWy4phlY6qk74tlYWj+4qx
oyG0KKXO3HD+/onxwTwziwu5QqOvLP+GalkEavQ0A37aKwyCtGf9Bvq+2456/0MOfXmhd7zK2pPs
5klUzZXQ0sxQnpzCTEg+XqOkgInb17MKFO1Ae1Lb5W3YbAVlUaHMp2ZEZTjY3wkcnl+rI6ToEOok
MmrWF5MiTvntlckaY4eenRxKoX9yQcFMUx0+/dsDO1wxj9cKK3AUnhUdjeyej1HMR87KqiWs9QVx
g0RzmNGYGlYAH7caf3CVBPSB3lDvX9MDXLRGU7ksf+hScbXY9zmwNWkVqOW1YavwXxndshrit1oz
momsXKSBG5ixQs14R10IwzPFke/jrCwblHEE228u+YdfWXkcxmQX+rYMdeDb6C9oqzlrZFeDf++B
KBxc/T+CKTPUwlNUSUNQx171E7ueBUZwdGK7R/QX46hbW/zYh29Fe7lM7AFTFwvUpH/c6Cmo/rpk
qPfL3abMKKCCkuBd5b3+upXHBGgCjcTK4a+PHvQn5fmnz9o8Gf/09TYX3MjU4VFRDM+Jo0ds7vgt
q19N2T0fDyM5CHDG7qrdAQ4vHW3343mvxb+QtmxX9ie8m6JtocSA3HLaINSnyHKBaEsq0LP2zRz7
u25TmAKiwv6K5X40my6naFMN4grIHrSO84y635E5I869YCG+PKvKtuImT4RP+7eiF7oyxJxyEmAK
ilj64pSGDHbmqv4ZlV3VoK5hspbAkRUIvfLAmlHViRAo/UtJM9b7YRsT+NMvMeS+eYgBO55E3yUi
A8VqFDlHvKdyD9YEEH1BHLJ9XuEGU3bLh0O6FKiKXgI0vlffVzs4VSLDuEHksY9brka+BnrFrsY+
5Yx1yEUo3PCuCpyxp0B1USJGjYJ+5IAB287losyzCpAKvhFVl5NlK2lYdH8zdB2tjEKZYRb5RTqK
dRXOdx5PewscuNbE4uVmzHwloI/yIRUEihQ0W8APrSVOfQal3znFw33tj4NinnKb9jwFubhDMDd4
Pj4Gc3Jgz+CK3DSl25fbn+5ti/zGmTTxRMYeZADb8OlKPW2qB2PvWDlt5MYKHAgzDo1FC12JWIDq
aKIF/d5eIwuKxzvYFU+CTR2FrYIxMEQCerNkBVTEc9MOPNb85mxEPMwLOq41AbEvrKfY4FDSu/NJ
hfl6u1nddIALb6XDgjJdwu3W3gqnZucc6hpRhbHVAoIodxb2LE7BOPZLITCfAPOof+AeWJFTaYbB
15pd805BJtTVvQktBaf9oqjZ7CNxGUEkvS4o8GC5O2kykFWuZw/WVy6mgs7kRWuasN13lzmDjd3R
/kN+P+axb+mvKZdivuMUcUGE84vIk63jVkxUAHMjTLABOUA45fWyYbR3NSSxhIdQ5uwQWr6sKb7i
T4Za8hgAWeAa7QpySkvwDFQgtiRaX65E+72PZBG0y+j49a+YX5BO0mnv6hwT4KFfJck+lzyBr25U
WPn/YFy1Lb9Vr/EffNwXovtVH4p9A3klOZGQmstEh8rlOw9RXQtkMB3TzXzhCJXEB/nZXKpceQpo
HsFwKjF6pn5I4mcLcRCAxldKDXw1rruhPVGcKxIcpvW7DhKrJTOSxKJOhlXuXPXHddJazi47b+Nl
euSs+WhiMf7x95RLcKgK7usnwvB5Q8D0tp57pATtuIySC9rz1ipamr8BpjeILY9lmJz58c+elnho
zw+8ls85k/TNDK+EKT38csDRvFG9wqg7QwbITIf3C7MjKTJh2cim6cHNbjcDTZj2xyLNgzFwvW/J
CBcMp5i/RKEqqeeC4E8d60dL7WsvBMiL1asdp1A/37hU2gqdOXEvvbS45tIXZbopcCWaQEyB3Dkw
XcHNDFdTD5G9q9bwCq67SEduEBsE2tyUln2dg7Ld/MQ7Y77koWeb7csCO8ucbaSSGDNPUA7xJ0NN
nOfgQ74pmVZwsPagr6k8oThqjanZJPpXyBSgXkvSmAur/EQQopJtOwjPll9MNj3OBF8QxDu+7S0C
CvW69p28iVetMApkDROm376K/Pma2RSLrAdapfnoELP4SalmMV1WXthq1NY9fg4ieyeaZCqWWhek
gq5J3UAUcDtEhYPyUV0gIIuzPxxhNGTP3XGGc3tmgZ6dwb1qn79mftzRv1ZiPxVKC+KWyaOiyMtw
QtMX5GEiX14evx2j3voQ8QVEim5ep4RluesRBVqS6y4NzgoNa9NqU6aV9nbuXBIb9ZbQ8J7wD7bC
+cLcL733wWsJr6F26PKY7Kf+hEoISftVA6VFgK8B13SLPGaRAkZobZsKVuiLzsJz0zbFlN6wx1z9
R+m1yosIjR9dTsPPo1zx8yyKnmgiB8J3Tf6g5BXUOoTBLeXK2VXOVuyiUrdjsCUF+FhKbVHVL0Aq
fPlSc1FzGdZjPrsc94c7zbmbvgcN5UoRFxZNneNQ6GnilCX9scnwrwAysB/UChwzID1jF8f45y47
KDeifOExn/3DD2rAinK5Us48z9b0eUNPerg3A2AQZfmu7uYZPTEQMIFa5Lfkzwco9L0fSjQq2bdR
xN8ylQQeTnnI4qH5MujcGeMuRwdHrqqZ88NNjMWt/1jtBkJaGhE4GypW1cTvuwN+oy05EBKRk3TH
NDtazEJk+u3SInEZ1UmkEco6AFgN3YYHuSghjSeAT7MY5zkSGkp/0jxJr3KOyvsjteAvqs+ECsFz
OpFjQJvAAiM8HqU2TiLY3Og3z9uWpEFDe4+hATb9RYxmLR1TayWvsRLI2khiY5HApwJuFo8cX0l1
JWHXJkeEow+alH7HK/36ZxG656P/P9zqT6X0YXRApvfn4K/uacgAflzrLaOowgX20ioLpN9+02ku
98WvTrDBUnoHDs96Ox8xpa01oradgNPu9xUT9CtLeDN2xz4Z6jwBy5n1nH1HzlNtfFDq+7beUbNC
+e8eeW2zFWKHiUfD59WYAAawjb81+PhIEyWP+vy7DSKccpdwnrriv7/+zo1k4lLlaxiaSpjv642J
dVVDf4PUiYGrZDtfM8CRmvuCh1FHB/SbRztrYEsA5WuefewhPJna8fCWEKyuYezY2pK2rDGr9LR9
uvEnI0dKbCO/simxHE0EUf/GCcljdBe5OO1jcqGk82o7ZOz9eLcgs+NjAdEyITdbH2PyUKjSg2X2
BJDH5usVtjySLXMu033idjzZpL6po0f80J9U+1wspDm1u/bd5OD90K0XI4ACAQ+MNaed8As+S54F
nRO2mvHJWR0dyz5riIjtKnkJtHXQC+N6PS9XU7KahDy1YnAN2OK1M/BKyte+rw8L6XvJLGIoeIzb
AFXS+pSKwE8833RRLUJINOezvnwSSQ7PjYy7JVdNtcPexOrKE414xy+YTEvqBQDR5gK+sjkkR1Cc
6Em+FewwN0AWKi54H59hj2a9o4SQbGiNhlEK1vak7u8VdzAXn7qreR5etFAtE8LREP2dJ/yw3Kbp
ZG9FY+9R7CZgZhka4jMBQXt4bTiSqcwmja9AoWLpqZdbcLTTtJBAecng97PI2a5+2yvJdnKsTmSR
OUExXBWDWW2LRe1cLNZebmABiNqVl5niS6lJC5WI7JmtIixTHBAM3d1CagUZyRUF9zuaNfb+F6uZ
aUVaCEqL+Kxz0NF1E2fiEXVwyIs5gLTXThTweaLSF/3qZC62T6ZaQpactFnAeOOU8AVxuOj034G+
TaFVKUBObzxiIfV6mFeQxWKLz9JmVSePFxkkNlKqO1FoWi0o3j1/IgR1JMI5ygBAANMy03FUkgnz
QauerZpKCxXKOhQCfuBwWNzg1YyYsIBYsp1OcdLAVDuEyD/Lnbbg/RYGbfYpULp5Mw66cOBrUOpz
bRSDIV+ZRPzJ97iQvdfFH6NnCAi+pWTaIcOFB2XVMfIpTRJ5mk34sepkt0BNnhTIeRKL3Juwdoh+
6TTqRoKqZeJq4+e8Wouv99Y2eBWL/uuBLRVphwoO0fEOkqgH7knKbQBaw7/GajCLsyo7QML6y/vO
MtIzRROMtktRyYHvJd3OZUnWtysPUDK85Rh1XPacSPi4YtvqTheXbU81vl7uiXMziG/zypWc3lrT
8Lf5HZINZipdZitrOqrqEycKnhXGPDABWUY5JeL907XJZDKgpm/LBbLw3/2IN31j6nZyN2S3zSxO
EhW0XpdWyKtZzplccMLoXREokp8hHgqD8RT3YLTwV8qjqlRS3n2WLiqnUxzPEXef0Bp2aN6dX9ap
Rvs79UEev1MZFd3lreVt7QqJ6rOTJ5w+ghV+S0d5QtGPnpMejM14COqbR9kKhHoKe+aMM0WR5Gpw
OZ6nOP2j7mLkm+DfPqAmRJGg6L+G/9xaFd66KbgVjCGK4kMphTpNMb30DEOKX2YEhFjWV48Gfc95
mw+BMYmUqy+ZlFwnR8SgD28G/w7IpdzdhBvHWYJz917xsQ2Tvjz1gAfWnP/TTXfmXQyVXavMHteA
R4J40riFlAV3qxfsfQ1b4iiJnXGUcoxmokeBKDXpZyVsjXY9YzPdsLnTJP0hc4lQPOFgp6KVtHd6
gVAXXaZDaGgQPnQpMRTzg+5KMVQVYgxJzqYbwwbES7eOku20sSr2Dy4wC+dSkYFfDDcDwHtXmXpl
mTsm14EqF3nJBrwLMMp4b4ioWkskevRPHKsQiLFDjZoWpXY4N2tpoCt4S9xXk0yi3EBqwq5DmgBb
2lO2Q37gG9WnPNSibXI+QMd9m9tlL8h8NEBCTcoSg+Q16RkCAOyFrFadxOSN0MpYe90vmkPGXsTz
j6+/ALoky+ne4IgJOuDfGznBG1dT/9ifUtzn59at+JwWP9E+W+4hXFeMIcLrBisbnLn5lo4JxnQ0
PaPkLCJHBDdTUKAcN8EkPUyQGoCk+s+F9aUAqY3kffB7WdtG/HRqvE7z1QZRI+Qd5Tm4aFfBpGCz
cte3tbviedvSa+SHK7IluL+JwRWJ1SyRNL9eYCv9l0kh7EV5kxPOD1olJQpa4On8pPKrcExogIxh
c84OIAbfnq4U4NPEm5Ir4dpKz6W5ejOnLznZDb8GOIE307qISBk0JC3KjFIy8jflMuCxr96JWiFP
8iMgNGYaAR+0LvTPAS2rh/AWJfrDiruEvfGTocyq+8NbuuwXxanTY36IGBQzOuu3xxjwKzOrfh2/
oXH/FOx0vwZbIV6D+olxXrzl/YX+j12F1UVDeVTLut9KQq5SAv0y5F+FqwHHdXbdPJe3sNF46z4B
hIogeBNGFbZ+OTgH0jh2M7cy50j82r8R7JeBrCiWlzr9eiR1N5xnW5vqtakrKIBhwokGHvaA31nT
5faOk+iLFESXq/nT+4Nd9q63mcCQVzU1w9uSlT3wzTjgxwwP1EiqRjgMSRS/CnXj798UBH2vg8AP
zpwBCc1GHSJdRJd8Y34IPtCCLOBSkGsBBfb1TvDDnNNcC/E9IJXLFhnsH0nNYCEua3EysxIN3Xvy
rYUTL2MUAMP3d3Z+T1StDSghTDd8lw/0Mjy0cLEQy5Y1hzayJpeOtq8klCVTLUS84ntjFQJ04GqF
g7qubBZGIo29k7lWQBGTJBJQvQGBwJE7MDG2OrFqXHvLrDK6C9d38FRT/JxBffon9Q8Z6cz5d2XM
FGPeE6j7ekcQwf6QC3wlGlzWM6orPBptjQJTpSssAjwLWtKEGsh4dbj7kQTp0ism7BAoXZ3e+8DA
J6HMpBc+qDDbN/jIgt7LlZBcbrEkO9V2lmFs8WbcnOZ9XrQPydcRQ8hREatKXj5rCxwJ83WAD537
wwL9xuklZiS9XRpd3Y9BsAc3BJnxtRJLecvRdXrsYyMYlsWFm3zP8FWcBtUojbqYcBx7w1srQ8fG
w+Xobn6M1MNvYVjO94cNf1crook4RnAe/YG4l5oV2EF9pusIG4MOCO5WFUtb+yrQPt1utJ+hcO4r
LP9pOWbIDyT4g33UMdckhiDmG4aVQk/WPaGYq4qbK3x1c8IdzZb9TqUpcFlslMbKwJTBGYDrYUNi
+0gke7UifzUozwAJdAiJhwxfip0/6c5Yy5QUHu+72bXTudE/alpbdjMtl0iuhIXIUto4nayC6tM/
2jZ/xTTQOLH8fIsTrLkXkxCfFDWFyX673etr4HSZMk9aP4n8D0zRE4OpnvcIqLN8I8q5tL6nVCdb
/+KkALnLNsOkMtb8uZqesplStiKZk7OTVPZ7q7h1ivSwrPyVclE1Xop9NkBgRFIx8qOSxj3wcB85
MUjLaifpPwQNojqmjdWmYgHyfS7xzwZWjifsk87vPZOp4AY65Q2fjEkvp/7+kJjxXGJ5M42zCdEv
AlOGjuysr8zVjTwOlI2QNnqcZZvptAOsvinVGmGhnTu8PWBOtTdJrsZSJErQ0w1E3Z9Ath56y1IM
zRRpiWiY9LKTYXGrwPgvBCa2kAGWPHr3/zyYseTIS0LLF0ZoRWN4aAxsboXCBTVAKuj3JC2G0iW/
S30gifawG2+636xuF1weaF95Ql5bdJnyGW3LzUa0VDQwcVchP4YmteD1RHkYFnh77f6zDXDHfbTE
T4V2RfC6JYGt7C/U6iA4A7qKYvOtL1qafUuqKtpClIPHFxUnO+HZurzS5v2FAsDJZOn1KiY4Eiui
1JW1nH56OFBJdoDvAFQ9EBD+Cm49gODrJ0KwAfQuvoDEGTKYK52+BmJQzGDfNviZnZg1x9n02eD3
U9sB4iajlbkkzehM60QfvTT7Vkb63EesqX4QR3m5dFhmtZgvqy2tqGZXjN16tJVkpo96lQtqw4Nc
aIKcwwSRn19ZRnOM9XnYCSOjA3d722qeAIYC6LKaoRxvTb3h13l/Nm1kHbh4spS7R7JOfV/Wt1yY
jz6C5WknZEvns/RwBmQg5rx/gvMI/bu5NOzrj+ThDjn8zC0Sh5GBiglup+pCApVewomLbwW7ugCy
jtX3k9lFmwria2WY5EnUeHN/lpHSCVytj7PTMeapMvnhnLQPIIRZerEqBAIErZgsAV7X2tc41WE1
NMlzAx+Mo0NLLnZyL4u8gDepn/ASbQ9MbVPRt5BZr6FKAcABZkGEoRnEyeOhqwiOlMh1D2hQ38bb
bSLYkO/6rUSMyDUqGAvzrWK2m+V0K/xXRRNDhLL1qTI5dpXY6Irrl0L2+t0No/0ztJnX/BzHaSfO
MJRYq4P4OFBsk+w6FUVkkb96xOvYV50OFRRzNIxyJSOebO0JkGEkDJ+WD/PHXcHikKxNwx7Ced9c
VOGele6eyMYWb2MiN8Cd7rVdlRWfJ/oqZLLjcXa6eon8jMb5KHCYpTwvaJt7kA239BITJpJUs2ry
4uXyV8Af5kz3WT8n87zipU29Hj1dj//QM15CQfIyMKygZhvDd55sCxWrj8IwUOvpj5Y41r7NcWXD
WlCMgY3BokZJAwNdBtvqGcHxFb4fYyY/nXUvNwTULVC/fTbcycq88fjVchBreS5r0pb6HXPiNAcG
suinOZXI0Jkjszzw7rgOthXSwaXjbhd+7uFiX2fb2AU+EOo5tWva7ukwEU1QHfke7x7j1j7EDbWG
OYV8kJdC8bhUpfkRkFSRXPIt/kybtu7uoi+/4ghT2+3ln5eSlmBPr7NqI8DM4lql5362ibjKvCOi
jI2j8G4OWwVQPykOItlD0nrxG/EZTzBLqJ7vYikLuBHSqnI59fUWwPvaGsvFyPe5JtJJZHBh4+0b
hE3RdZt4qRkeA2kuDuas1dpqdAkWVQXQNrtGcq4Oi8qZ3Jz5VJ9L9029WPR0sDo5hxWeQCzsmEPE
bmvaVBOhew0qhsklsyE8Qsf0QWPRnqfUTXUs+VxTErMU4I9cKjkEqZdJrusY6W5pDj7DriwEH6aN
W88w5I8EhMWFSl5hKMuC7JQkMGzEJvr5LNHgU7hMP19iRtxtpWKKfeTs1XLdfEigsHEBBqdS5Hjl
xWfC+VteP7JbQrEOgllYIh47OSkL3l9Ew9nYmpr5aY1hTZsT3bYJRPVFDZbXcFWAHypYlRxQ3m4R
jZBmHZa8BrvVl/O1C4f4FL5OllpjXWMC+HmqPWSfCB46B2lmb0006iCN/4oMT2FYy47AA2o9s9fg
iZYvMw9XU18ou4qqhutRP+iAwxiJscEb1bCDhAuDEGRjrp3CXNqTfjEWZV26tMzkqYCkUNUJpIAU
HdaeGZRMyF1T8DtFPJSkVqgA5AmxdftYt6MwovFw1tuSqUpLpslVdDxfWDTzRryeNcgnFiFzMSCm
Hgmi0DFMuwTzxj8GN9uYh0VuGph+HEhO83GLB4HhKT/bWC6OJeOMmDLhYhnPiBt2jfciKtTM0O54
gdwx/MDuMmPmrUmuaDiICjnIkdMnf5iYaLPlg4UrK3Qa1le0tzdE62HC5SulAM8oXbW7HOsAD3I9
dxbgkIILOeFVSkSa19iSaUWc1IemAPl0QDMwIqZZMR/tv1lex3vDub97Cxi+xnmZnzTNKOIS4BPN
iIk3LG5mndKpCEWQOcTNehvD6LfPdu+Ihnj2VKfRpXm0NwWThCRIMtKG///6UnEGXfe/HUp7PRVR
3FDyb5NrgTBO3BaxAHJ5ZcW+f9iP7vNty3Rwxcl4bwAUAwqtejXebZ50sB98OSO+FuTB1afptdmQ
QnSYbz9qLxREzvsr//THqUn2CNNOP2D9D+yv6v6wMDg2fsZDoKs+g9sJnnZ0KJtvjphj3qTiaQi2
InUbI8ys+ZeBgjIiggiKr/GuWhMUsV99yBwEOWb0HJDnM//jXgAv0Z34cjeGXlkK/0HtTehWsxTS
vbnpdNdZ/gXygJ/JLSx7MjNQJw2y54odXFziTCK5jmmhck1TH2e7cAREn6nxGVzMDBRcOWF/4Lcg
bDsdUVtrEI7i/z8k8wEHR9BfUNnDvEmsuZNKCNwlThJOC5ZRvWBp+NShOSMPiJJlUV4qkK2nYlUH
nXAuEISgK33XwVADtN7MG18XryaG4fY8CbtasceAQlH8ARee9ljkiZYRpRKIsKKJSyQYYtLUWTO6
0WxFuZHpluNMZbDf9AAulD20UYNGMh+p0pUNr85MZWcQYQQixSviCfTBv0bx1v0BIXPeXcbBH3Vo
oHf3asFAdXPsP+SSVUoVatGemy8Kc1M6M4w02TjXSx9wizvOi6XbdB0Y2vK+8L0/KuxigTTQpiM9
Eua22PGDQmoRqy8nz1Fbq6lNyMkXaTnbu5fKvgr34+THV0vF2qs85ojF03wEZYSl0vX2WSYfk1sk
40Al+hR36adh+Hd5HP3cD1OhPuQmYdBpKXE5H6fq6gptfBKPhLOM8acphyAk30ogjR+8HzskQeW3
SuMQmuN5s8hZqxiiVEVL5/GiQx03oe0T9boto4xc4hO5pWAyWSLB5NSd2bMvSrKtQT8TwOH89i+0
XTdRt7WL5yB77NNkM//PTAcH8Thj/NIIwVZRukPabJ9B6MsHlBvhOdgi6T6hyaEg7jNRxt5p2ci0
3eWcXJNNnEdIOLWV/ogpcadg5sDc6KzwgA1pIJNo9FZO3bI1kmfhJUonuKKJzhV99ccMfFMFdQtV
i/I0In+7sPyB+ga+C4xxqWKZrTDEKXqklEAzTQHDv5Zj6IWrsYKgSvqsf2Buu9vxzh7SXK98Phw4
HRqkRKr24ZDV1MxVb+oAu/qXWRbB8e6r46gKgujKAYo6sOtzd/zJQBwQ1VnqxOsSgdlV58ai+2rj
LTJLkqY3WiMgq/X/nIjUCX0ELb36N2nLTInwmhn/e+HuWvICbsIrMpTfQMs2kB2s3JS2XXB76/zj
dPjDXf1isWYvl/CT/rsukf6IjonAwSUDPqsxxQ2oBbnwWF8T9Rh4ma0mP14pTqbB2mWNFnelkuD9
q8KHOyM1B0sNXxT/eHH5Fu9VmV8rjV+wmt1iC7tj6hCQFOUH6FlKL8EBWVyUcHCQtiDfmV1YJKJ8
Vb4K+ny8ITdPBflhd/bTjBDbYwdhRZiJ6FsvajbggQLAwRb4Pp2OB8jySFGNMsfPqKB1s81pF+kl
B57g6NcpnD2ZAr9SbWcVhbm/3e8zmqFWF1di8YSonWHc1PgkxUObQ6YZdR0MolYbkzTw4IxH+yC3
ygMbO6x3og0yyMKh5LtwbiEZVhjCjMqQdBZ9svpZEDCfluShHYAzZMfI3ESDwWHKjI/LXIKV4KqW
530YfTYkeCGJ9AakbU9Fmykq2Rrbv2pH7lHr2AmUwNeJUU3uxk2chxFSyF61Umuv42zZYle5pODa
iwp4AImdk/Mnb71sSLhs3jNV1CjAxBDnnOpzzlc0sespdYu5HkN3G4agF2fNv671J565z5H/3W9X
MzYiT3Xsm9pZMWfyBIFo7aLwHQUBhIyWvO+Is4NyxdjF/bfl+aDxJxbiWTAmw3s8sVyr2m4z8OIP
AF9m/2IcFfY2x1rcLHx8m/J6jqum4A+utWjkWc44tVAvKV021TQRM3w8q3Xig0G5omsLRKeNGd1G
cW35XG3X3c6CIiQLjuPJjbzWihuPmJEWwK4wgmRd344yuh3UicvZKCLR+B9nkJKMYLK7KQulka5O
6ce24TAakLH23spudUaP6ZqktLOrOQvQ4uU1yomREaCJ6imgqOoGPNvEMCjLCw8uJnS1mv2Yab0B
IcVaXwB0S1BHYYyRR9eh+Cunj1HwtYc1rb5ggwvxN1dED+GFhgvllWbbNUPNeSZrWFEcQ8ABKV/U
k+xe5DRnnxfUBU344OQ1RB6PRK3eXiL2SVwNEBFqOTb+wAS+JJhykEERv96dBzi3ZfsVcxl9K38f
qzQm3iPf20k42UvYt9EL8ClFH9fmueOYiPMJgepIg02KTx0uoeBoaKk4Uo2UjqHMBm8+aJpWkPHN
cHBXripVxfjSZhgD7d8HRP4UyI6UIrOagwFjYaglh6AgUPP8L+Qm7iCv0Eazk7KJKC6GcNuh/Sp5
oB/xFpbl5BAbX64pKWmghn+7oecIK6XN7WzALZmR4vzPvsUpLeHFUEtzh81hPOos1f08eZYbO1aR
cWdStezPbGu1qmQ1qlv5aMbCkl22RcyhwfzygkDWj05MyxnSkNP0MDGYke8lBqf6RVOpx/cvwHHu
wZJvtMI/+2hXGmY9i/MzO+Psf4gH4RLUUh+pLux1976R+kbo5F2r6vTMBWQuNHuzkOwDQSaOff5o
Rvfcki5PgU5KQFqXz1nnLJawst4KDz3VpsAwjoEBUrgTinyjTdcopzAeXNoD3Cv76HQVCW6TB2Kr
V+yjcZ75a7RxtuvRfJsfeaq+3sRexXdvEiKrAdo8NV/rbkDd+bx/y3iw3nQi6+pvS+mfo0SbSIvY
2mGTpCvyUSXZF24aUKNeLgMtFacJKG2iX4bu8YtC5TUZznN+drjQzWFxgaR+7N4Up6l5Rrrh05of
yp8SJO3MbqeGsJYcyltmpsSv/LxspUfVo7KiYNYITvlVarbpzJaKUfzMHMcMbG8ldGR4qBVZ6NAd
OFnFL/rFe2Hl3mIapRhS9su60rSH2ewSHC6NXC0N48XXEbH55aYL5nfpYd1GS3FvrU02BTjLoXnv
hZ8KIbx4c9VDum4/vGOcJ09TSnrGHNCQN59LpBI0WhnivFYkTjy7TF0iucJqHsrW+5noNiU5RHnE
N1TUp+YOhce7nZgussWcEQBi7kUi9aj4EXRgI1LJvu2Uoq8JnuzQ4TUmoyUIPcEnKUtae8r/EUVe
454pT4PBHWMwR6H4XF1TldhDnnfxGVOq9FJncGo2ABkXZJCdLuqlshbGAujbdM6gffj3e+NA/MwJ
oqx2YqbmkwuWswoin46aK+f4Mi+sMNVgjTGHWhaEXKIHLoSnTzFzKnh0N0S8XmYLFEH+5v3hCJSH
GTbyAc2fkF4dqfDn0tqd7r4XqStVpl/tUkakqLZ5LJ0MH9YmqD6W4c62cFKCqkLyAOtNQNgyk4HN
lQZVBag7GMRPfjEuvsafZKt9DpiUk6idgAhTNOwsIw/nasKuP2ryU2sCBfmaYGe3pL7aBG3what0
aaX8qjJt04TksRVF3MkGYv9R5TkYq1lDZCAKP4dgK4cogRNYXaWp7nRUKKR2kkwA5TntDdPvRewB
5cXSfkc9P28CHuhtyXtsyAIWQSi/s4a1HbBG4cmHTcpAY6LatCG7OOUVZNWgbwsj6VKfYv8SHGXL
uw+4EMK7bpfBCXRcAafcEao7LFOyflMMo2V+GDO1eB2pi9eII1K9bXrDS8zM7mwM/1W4Ari0qdWm
XxZdUX8yZ4lk6XKtLSnGQHAZx2ngOuiOXrKB+e//4u4fcyB0ivF/haqUagGMMzBaRvkJvBg4uVCW
IuufFTvdBIO0Kmie4OuFlIFZDK1rrgnizZ6HWS+ZmLu+hJOX8RqSk64PtTKqlhNtk1ogyx52yYBs
DqQtaa8Yyj13w3Ry0LY+kH8r2fAFiBk3gsYwll6va6MyPo54BVekqzNwrLYvL8db0UC3dlVaoLNa
/+ac3I2QrfB+C8swoHHVUZAxEmYXEnk/x+7CJZeuRkqt+g+Vg+CHgPIYvTb0IbfRhOJ2/subG0AH
H2mV35ppcc39s9KA8u6Xu4LHSDWI/AKAD5ea8iIsZ/9hcstQFblhfS/2XtcJWtmMWTWrmqDvA+Ea
csnUmSQJlDf1Zh7UoXfjTOHCbC2O8vOt9tPqZAebNVYdm4fk0fIev4Agv04A4bZ7SzjdIgc4+jxk
SK7jHeltjIAsqlKmnfM/zL5bSQuIfWsMFUHV5QiEmSKRl+dgL+6POfBZZlUp4tlRZlRVgsJFBjzp
SazcPpSZMlgr4HRg0vsIbbADbyYoTDdNNt0jVAeqbj55Eeok58Hg/bjre+om5j6yga1Zx+zyyIZg
pbEZilqhjlQP3NFMywz/6F0LX3RM9fBIkg+QgsyD2A0Wp9ClhY2Eog9wgI0Vj56m9iGPGGJoe4NR
mij4dUvCEb5tipZLPnFu2YDqWXmF/Hwf+uiVHqUl2zl5lE6CQ+perKIjlPWYmz/9ocvXIuNqykXc
x2Sl2L5j2eK/ZDtdHMl/29u5xCNHtLDKAmD/ujsxJB5r2UAlghgqpHGF+2NVZLkzGdtNYTn3tx9N
rvPnW02ARY2j4ND976o8YC1wPS9HQy3hDSr1ohaaWFw+HjBapCCmLrDYAkLprydJAYWMAnMGQELB
GcttyhxWu7sWSWeCaKdz1IBz8EViX+LPliUknLvcC+nU2+WlW08vNStShVBorBeJFWjJZ6qC0sIr
1y7si2qBGXpGtdEjYSTo7Oh4GlKnvhzf9qagnZ3yo1JQ8d02ZhLDBXscePjRTBimye8dEjmj5jQy
dBpP+pH2grUSDso1lEvunZaEBWdD6ksNlM3U6TU/uiNPVuoy+LAnJbnp4/SkiiPe4YJpehI70NVt
ufnMaUfYubLKFrnWcJ/7x8KeEkAzVMYgUVasd4Lb3TOMhmvlxniVDy1wSFU9bdl7sPhxJI7464b2
fZvONxLDfO0srR35XuAVA1LzRQpcKPEH0qY+bbj2qw8uCToj0yMGuT4Hx4DUjdIFJBR/DQQZABb7
lgK/c3UWqJpCnW6vmHTuums45VmY/bZ9k9zGj9gRflkyaul9Qaz/xUseGTTqaOTcZLztb6mLO4Um
wdbnV5NIqRe2gHzOycW9vu80NCJfl+iHk63GIZnzoXGkisjl/PWm6H69dGsPoGpA5SWL2PWw1Wap
qlQ3e2Heg40d1FLfYAvtD4y0Fr8wIYTWsXQAyXlTZelG+9HVABK1uS9THI/qW9Ei7WnXHepcRHkO
VM68eFi1ibeZKYctgo87VtEqWjeomOQ1NEsUMretBhjXb1rci8xBO/bwj6Wvd4SbsQsqsVHgD6rA
RTOtuoteFvQlvuIim8LHVrJx3gvbC94iwK+tgt0PKc61Zbq8uilQBXQS9PYV459uVGPGQt0hdV2b
/7na70v38YCzpMBuvYRtdbu4B101GLJTuKCVeZAv9KGIaOX7wM5AR1hwCGAwTzDFMzOxDlm/+VcC
cduG7wQeLfoogFS+fprmmCXHMkFUZkWsscfns/i2ljR1/Q/N8f/YpyN71JLOiGyhtEyjC1ACMyN5
Pknf8+67rXSNBBsYRo5XRu+2/kb5qR2BEDGyvU7cMzOqK3fQFP/HleQUGwIhz4GI99AHGStYF8bC
rqixco9B/3F+PrWXkCpJciVn4j6Dy2KDab+kELbBHiopyJhhuu7/B6yrJzj/05ZaR9uanDk9Y2Pe
zuw7O4gtrMBEq9YlS9rk1wvYuF94hIsKEkiDOyitWTCSNzj6RPMC0oVxhMGj3ozD6E1ChOPAuiBt
ZUSytAWkNc6St5oh2GkuG7nLNsKWdDPVlb3xstppbeX2hplcw2Bq+aNBPvTTNKfk57ndt2yR3bQB
Fd5yHTIJco9FSVdzFoRdSvTLNldTq7p0zw5v2JbyiwJDVHOBoaIgB0HpjhRkTjORinucvbOjG8c0
8WvRRDATJEqJv9/l6eb1lZ6npIO4IzJUx9yqtMmuOStek69qEp2OCkduxhXhklPlnpd/NSbNl2P9
AScGD7DKw4UNaxnf2kCSByqRbW9f+9kNhjtMS/796M/xQrcc4faxggMHfAo+IsBkv/1nC5W8tlW7
1X1WZNZQUcbKzzwBUB8+s1OuCzlqwOb1iV/StBBfEMJ4E9pRzGluVyVATNFMQWcpqqxdCJcB85th
z5tBB3TAyAAUPAH6OYEk94a7eWLtCrJAz9JNwlNc2ynXzA8J3l8/E0feuQRQXK+0Xq2AEpwQsx+6
WAQIIqmaOQq09ZN4OM4yatuSDAnCyMCgeu22BJgyZa3x0rL5M3yRGO/LsLgrPibXS/EHB4/axLAx
R9pBSRYiukNUS7SperOyMvX0TBbAP9+w1yK42d+Eq6pONX7bDu/AB2wrGzFRaEJQ9GDDBPKKZ54O
m7gbsXJ5ROP5qACZw3DaH3pAe7ce6MyjZa3jVGmWzPmAYIga8ail6/sw1xhFuwn/r2I94/C3S1k+
ts74duokwVnOjVIb+hgNyA/H1sfRIt6GV1QF1+bTfdWZsEOddfl9VRHctHrKsvhldBi7Fli4ZAwg
WgdeGRckheS2l2AwxnDkmqpIiNkCbut6qWufkjfYpetAciIhCpWxW9H+kE8/1m4gf65RAau4o1Gc
dcJasl/tMsmJgJgLvLMltLNu89OwJSRJCEEclIjmRsc4xJjVn3NNOiba0lroplg9odYCQhwoh+Ar
505SZJDFIOGOqHJacRQU7HciEqhZ8gKhW2vbE4E0a7sMX5VHGg6vKoySPCaK0WHv1ya5xmZebuC8
6rDeAJs6qTUD/v4Xzq4uL6MZHWOtJGvX/FEp+w9S4fHjSuzfx3fHbdoDzHfDcpdd65s5V2oitaIN
j0Ddkgtx6odpcmlvbtNlA9V1UNaH1owavKUy/JQDEvrb45lsAsJvU8eL5i90dwk/DgInGBM6E8U7
mbrwMW8nM8fE424IBYIKDaL8G5SBvIf/39pSvkmOpEiFGZTzFzUd40RpTkllGNICUEsf1AmhSiKq
nUyJWzAoGbXQQHdtxCLM9IBS7llP3BblXI9IGggfhIm6/aT2kkSJ9g3fZ/DWrLSgyaB3JAmdKuVG
JqkMSswxSRA/bZILGaWcgJwfifXRb3U/ajIlzJnSMWN7+Nzh6BPMUPXpX3SmA5E6LY/zDSNI7HK/
jqKgi/OJZNUcwlaFJ2ey1H1tpivcV/iqc5NNvgh81856cpsh70TZWn1diU4QTbQ+YAHHJ5u3sY1P
2tSZpc2deCTY0GEf70XBsv4wAisSTj3koRvqncay5DDpCJD1WZsoztDQTzngMpRrQgEPVknUTZQZ
QqUTK12gK2E31bHABpBjB6OK2HBs37qDp+ALrQMtz+EJtaYztvQaHDBswjGxxD0DvojB+IMi1ECU
2gJ15zlseFITJ75SD56GYf713Oe6Nno5M3LIGyVjIyb1/DGpgjr/uv2TPo9JapFTHLOPEE7PwYHd
pLB+MuDwQxb9IVbizPP9U1duw9D8cziYrN8guLQLTpTIN3PxKghR0C/P/ECbxxxFwGAeQPtwlUsa
6BhoguFTzcpXpyqDp/DtYUoClH3prEepZwC5zCGp/4NaOvDNk/1KkV4TygQMjwmQpVtfyqxBiKXQ
oVHsk/AV2q0r6/VPZmtUYglraYwwlSHBBrhs8ICojYxTQDT5ykuMfuH+2gZlhI/xDuyxZYZtzb3f
gKiromJ4WTXbwhR4iiC/Gp/yTCM8wF6uD/v42xIqMyP5PXunRh0DjvS8h7k0ot4HWBUPdv8KIAA2
h0tuUsS93d0f+AWEGrd4u62bVU7ppzV+5bMfgvzcI55DoHNe+3aIm5Ez65+5wU5cpozc8l3/8O//
Cb1mEIZJ1svCKU/P4pqtQXcPihT45Hn5wcIHZvNokDn++exlebjmmtLLOwVOXeBDZcSQ54QpOd0W
KG4dPGFllO5amAoXGtMeGP0LqB5KT59mVHAsYBKnVPJxdHhzeW3UXAVpj9B0qs85YH/6cqv7sZdx
WKvHKR7WktWc7mQa4GYvSd+qDWnBxEVpPK6q+EvWh/kB28B9s8D285Wj7WV5VcbP4hlor23IlXtu
yTGDgqRHz++DsiFSVyZ6jknf9ENkuWNJtxlURVPoXrVUusJvpKJalQtbSPsfGs45l/FA5DI2WaHI
IXgQ9F2YpMonsAkY0JPN32UblA2Sh2Sv2bsVtrizB/KNpIvnvWV1kZlZ38OW0cGVcufUeLDOa9SX
i53QHPI2JL/X/+iclInpzpLiDTNqrVbLyWmU2V3InYkdMmVo/FkCzSIlfqaMMVhihzYjkta56WZD
G/Oym7pTkgjmGoGv1p/C3yVbWpkzmuI+Jq9Sx0OLV09tGaP9BXVONYPJ5AaH6muIE/qKOyEz0dsx
dKvn76GY37RMlpU4809ss458eWafY6OVtIBP4SYBgNiPWeal75Q9dqhtLzmexP7ZjVovnhqGFGYB
JAx5SMTGP5KS2rtul9SUMlacvceaj4GQp5WqOLqESHaaIB3+s4apub6h4PyvaMPoyyRbpV1fqYL8
7k0VFlcU7y+HbIYao84rODu3Su03DkgJ8DUwBuFAtrmCoD/ubUMALDMLb+IL9aVFq+YdKr/GASW4
1mOhXOa7RGQyYtSl4F22P7tZdhVYR1lRjfrCvmYfscFxbNiqDBoGIAZ/K6i43FPtZKvNQF24clt+
Q/Zwc8OxYQIMOhueSYJJXcWvWXTnLDe4H3tQ/y50DaQPXXXK+XwzI/fer9CniMkpBKvPRMVMHRyh
rqrIpZW5fU+xEyFArd02uoCN60YAHoUdhJ1sC0kccBuZf2VrQginZRMCOLjv2pu8IcfLtUYSQlIe
JloBj+UjPFWGaAvflNypOtmV53aicl82aEXG7zYCkWPplA2+EjrU0UYTYp4vQI3VSG/dBDAC9+lj
h4CwYRUlgBW97J8z33A+Vaxn5kBAP+XLuV+QAFqHCjMN84kbJe4/bEzbIBROodZzDO7+yQFDBVa+
kPNdHS94EGxhq3jYbmU1GfQgvU9LYv5za7nuWWTALG+A4slrt0lq0rPStNd+6NhMS/AwPzUn88FG
WhaTvdXIem/BLJrZb2PB0JXG3ACHLl+X4nLaVhH29EW1OVnqJwu2pGq5/5RJkAMVAmRvaBElrBVN
Z8caEdRrjAZ3xnmgyKepS8LItGSDtREiHuMJkaphAU8hwy72R4xZ5fBg8V5dfp698uOQMcIxKfBF
d0VxIeWwyz10GZQ13Yp3IqWb+ZHlxcjcKk6dPK5BB6ZyEymF3uDPZbn60IhsVK7tApppNyrmqx+b
XuzGdvkT6nPg/jvDKgelNm8D3FU4ekMq4u+Mi1WxpxvKsax7aKI66zuRKDZabOOz2frSTepbmV+I
mwq/g+ehZhcOO/g4y0Qa1C9FlUNwmI4/RAji1hh1gg3wHYcxPDRCcjHzwUBC/0Zfyueijgr9+Xan
FIgMeOnJiGtaeRe+MAAU5q1FIkqYgpUmlS9ev7ttmFtQ03X78RRlgCTw/P/+2gMV6RJOtrokZXqN
zfXIObwmeqSIpD3oVPhXA+SBLeoX3sFvF7OOt9jmeW7viOItGYJ53QqQqnabq4L3UsWwOSH24xtl
ORk0r1hMC5CxTNUQ9qXcQ+XF/x8bYLxEeba9patfexlbra0IW3T96G5zijN8Yy0y81nfWEfF8T8V
S/mBLRN5nIjr/T7E/lPVeomCwFydbN+383nambsn+GYHGzVohtT/mVjSyqjOwQAt/gGjBoIUR+Z6
AnODVYUwXYtTuE7xa/eZ4RC6uK2j7+WrfMgkGSCxW0BGUihegPe3kddtxErryoOiXOt7cury/Gsk
Wbj0x6JYjymvmWb2annnVD1gSRBTfoQdrtv4Qbn97qoIjxGxmz1GfLYUzeHQDiT43OfImTeruc4S
j0r7eQTYjrsr74HUqc+fZ8Gbzv25b7c3wVFSyint/212/gtec1w7CpJ/LJ3WwV8lQQLnafD9z5pe
MAFsM0aMzYjvKDquAZIvcDOIzrhmq/vIqcM2nFZW0zQONkPKkYJj/qPu9LbtMJDo7JdGuqaDlod0
rKjEprXNZ7aclkkGXhhsMgUuB5sBnCSTNhr+fRJ/rIS0dL53/rZCziOVtT5gNS3zVWd2pve/T7MW
47Cq1+32h1PdG7a51Fmd6IZRa5vTlxzKdKhVw2MBRgSDkWbysUv4txcb/u7MzoyjsQ4PnBls5vQf
7pNagn4L+zhDJixG2GP3OMnSeFmi8J+UebzYDX6Lc3zSsVhTCRCZSGGrqcf6JUZFAVslXnna47YQ
Wt2sUcSUWJVfiISKdICqKlGZLoeKO9ql9GojZ3aSWvDZ+mJ1kd/FpsZC6/SzJh3by64wK87wefrr
wAu/nXVUeKM/wWeoz89H79ocDkOekBx9YBQIbLdsvtQfpig+HTuhZ+6v7tu/0e1JXs9xYy9TAtKy
v9kz4pUnuIx9bqrLnF6ZVRRGhULOcO4eEDse/r59p1nZm84MuXZu2jYG94kWqPFyPI32VB85t5Ts
ar8hXrhCSYnXn7j/VOXi8dAIhlYpLNeXASrtXNZLOoKCQFV5SqFQKEUd3PUNcygpW6qwGnQDZA2m
cNsy5XGhbtV8e1hoZKpzWb1Len9vRXFI2sLO+DFkYQkSVZQcvfLxxxilUBYF3ubQK40MBwDCraoU
zNwNJRafVnaDVWvNf5p/uBcx6y3trWlh2jo/IyCg4bg24fj8zjDnOsSe/BOTva/c+LOKbxGEHOcu
9FNF/AAnQB1ucSB0gvm4GqQuYeGzQ+EhrMVgItV96lF2Lhzw8lumSqK7IsUZfGK61Y4hnACL0oq6
PV7yXt2ruPWvIfZXn4+J6q2QKAet3/VhQ6RWx8tiqMgei48FwIWr0zCm28IBQTWqG6OTgFSTQhlg
SPn+o8axwKpeIzphERZ7Cxb2HY65LxLDaNC3nWofQLOQX+Fe9rUnDt3/PbqDhzYMSYHpNWzG/xEx
fUd8/iGtAh8DpQnVQXbBYVm2dcVSe0VfD7ee1R7LggK3Ne3cCRC+AMHYa3AOR0dr2WNGvpijt2CX
ekWZ81bNTudE0LZyhXQTzk3Qi626YKczUeyctiaNGb7Ybkzc8eJJb+tu3DiEQ9q3PkuAFWhlI6xP
DqzM0e0FGY9y4odLifvDAGIIJxBJn7AdmiQkZwH5Le+ev63L6DF1+CYDh0fC1spX/b5qcfka/roL
6wCcfjT+P0fe/tr9IJs8R1AD0soTAeWgzsiBQZTONGyLGtShEuT9L3piwxVDx6Q5SkZNj4TeHxbO
ZEVPELznSvo/KNatdPqpD/+nqpsAlmQust69zwp0Jk8sQfw0/i3Blu9BhND099y8nhRtbdPjMGft
HOpjeQiXSUmwbdmg2xtavrW2P2tOLM+j/D+thWEwt3p9gPExg5G+bdga3ehDIALAcpTd7WNpBB2g
0PmKF+P1Nr+0xqBpzu4duAcViylCRl6Ja2fKlXBfcaE8CuwsA5bRohhZB3nlnuvtRPr3ntnP94c1
xcxzCse7OrSAJKxGtEOwoLmqn+1rb0vNY1cpRUDncw7AbR18DVtFd7WLekSXBUMy2d6B9+16Sjnv
p6Bb9l9kcMehHR1F2uQknmyQasF7ED52kf+sIQm1wDmGgeHbsfnmgrPno3kRskruBz+83fAb97Oq
O0mAR7qyPzDgwroW5zqRrjfNfxb/R35cejmUkSLB3rTfslPeDKrssMYEgkcfmrZWJCVhPKE7FO+X
Y2pagGQFpqiPWzXRuzZAqSM22C7kYf92lfGhePNVed291Mf0z0V4IUaPs4IpsMhsZ1kVyk9ziVv1
j/l0WpJFG+/6QQwATmYZQNqvVF+LD2GgzAe6KeoF8H1mcD5SFoDsq9JIV9mEjDhsxsEzDz/gcGEI
y+AwqdoifCpE39FmsJVOX0dT13522MiS2bp/BuAHTBzk+6545XKyL9st2cA+Y5m8iDWq5x+TUudP
voGSBM5AK0WDI270D31mtH1pOIQNTuOQ3ZCCfhrRIxyDWwkFnn3Xx/rVnEIQj6VcBpMZ0OmpWvR8
UyA/nINhhBd5QcDDaSKHAGY0maB8JoUm6H6cSXGAQMLvb93QZ/tTCntW7mpetqeSF4Fg+AIUwzFt
70o5BdsbjIfrwgT1I/K25S7lmLURLDxJADtigpW+MjZsd8LuspI8l1SL7r0/PR2uUFot+3d11p1J
v3yV9OnuADO/gBsrAgGaXs7D1aa++6ajETXp8setLVjftLxcwzFsQkXckW5WCnDc0n5d479rK8Bi
tKaQvBU8kjeK86P7pN7njQqmWQO/kWIep/23FkEIiUTePe7qdGqtfV1Id2noGtcD8h5IqD1uExFQ
QgyZvABZJ02mtApwcvyYS72l8qfjVcv9e6jqecKsmVkVR+jiXnVhLxS8CFfn7oCrz1Wcey3AE1Y/
RtFNOgwsjqPcoOp9JEu+RPNAuj+7Y6r5Min/fzf4yJ6I8P8bz4q3fUdsVyJ9AdFqIgavsp5nZ9Bl
ChSOZgGbdGCKMg34HZefI5TbDo/AjUyatauBr+2biDmS7ueW7Hodokg9EE6OKtx0KauRfRkdwKNj
PfdE+AiOssoIWfsakRdpmxnOHZErWrqJjZj0GungTM7kPpH/WzBF/AqTqX2FsTnPspcC5k6RQXI3
K4QY8/ytsHfdhYcLscvkHkzyLmjKNFxRyeMlU+r5OgZOwEms0wYtQUPWV1nYn7/UpI7q/qUE7j9o
8VxtQbF8kdYgQ5UIpTAHUOae7O1hNKzzH6kX8FRWHPyhO7vZrYeX2PYpW6cnVP8iOveU0DMXlWOB
/o1Bwi3epMfH3mR6zC2XiVuG5Tgd57cRLZ0nS/ssF/xq7xJSXt1ZWrAhwXUTtaaJiX8RftTrhfv+
VwWZKIfnz3TNw49zZVnvWTXgkGonjLOn8yKySUk4t/mB7q/FDssvVWwbKRLZgbTKeTj/rTb1ftr9
rm98tGeib76AXltCEYsYSut+I0G+ARS6bqdjAArwFbCqqYXxRf0YfMv7nG3Q9IbNPqMBzK50Mqzr
FvyLdbBrJrB/eeCq0W3milb3TxgeJQVShD3NVAVXpHJlNV/OtgQwDWX4beP+7O4hgJfioy8fODZV
KKG5rcEnDM7ZDggguzqiDTuAfSaiZlMW1R+Z5wy5gjXMuspFjbqZDAXr9918P+qM3OgnTdKWXdrd
w6s7ikSNWIOUjpp52g2jhb0HAS4Cn/IZgARN11edhM6tuaQ5HtI/1uGwoECw9rJwaoEb3k8KPta9
vtU5jT5RoSq+qeXaQGkzRuW2FwIwrlyd/VMPOAoh3Rru2P20vz7w6N4kpqlmWu5jrHTQ3Wa4RR7o
ZSFpyaZspA8OFut/YY7CEiTDwm/tRbuea5KJwyzRs0shjs0OCMpy7HpZvQe1B6Bb0mcvWTc/1G6A
xhBuEFg7aTpXJcUknMlYBEaadx4fmfzP3nQjsf8logE4cS3zK2Tw7ggMigH3KaWSNGZZvC4cin73
naOkng4pD+GRhaDHH7RwMwW74MGm6DqJmC4fCjc/cry2AFs6zWh43OiwlG0E+YjC0cN4k7FzKK7l
BIchlf5AutmTJN3yefUe34d6QMDxxZvGa0IYy3NH6XMRP/taIb1k63HNR2vOAOH14iQmbqCvDl6W
CXr35kTgQChdg2opCOkNdFv85HZz5C9eIAkIvJKLS61kbJV1tOdcqN3b92oslKbYK+Nt6uYFKo30
D8z9DMBCmtm4Dp0PxSDe3SMrfl2CA4N7xbxjFMKmWwuA4l5MOE4eOhbPBQp/q49DtoObCBYUIOWj
duI5JRC3juP665i868qaixvneV+INQSb0kYggjE0/wfcgbjghsgh+16aUNZxPYl3w3L4ZzSDtaKn
eTTzFS7s0QVHiXiVUOKg12G4bZAutqBlGbQsR+Q7mFDJT8QhDKUh8Xp4w3fJGsSehUmDpsHb+1FU
/h87O0cQzvY3FY8niS2mzwvu+e7g3zpPdVm1721QLSVKyBeKLe2GuxP5LuY+yyObHCeLqdNtlHSN
F3r69Plb6t7unNqH3av6Z/Au0BUJ83QbZ3XhbKWnZFYYxzf645j55sSo1hnzwV1eMJ6XQ88Q+cBc
UTW14kjyU6qOrMkGBOzSKglIlvf4xenzARHbirAzV0hTvd1KdnILvYNJOMJpMEaEZmmepfxsVDTu
dqN7niV60oVVPjYN3J1DHLC3xEx28NZXYZGmos26Ju0u0aywsKmhAyNF7O6HjI3TlfBDQ6fO+746
s/jFQleo6d8MKahRCkEbBqIcjSvjJBiKHOxQ+sotys5qHmvYR17wen+Uc/rvoaCr20ibY0QwSVfq
5s3V5Mg4oIRw/IzhEbFc5bXqESkxIX9tG2kEbiQJiRt4X/rON3gsDk1hgoUiqE1jXTlP41D5fxWs
1QoORlx6EyoJnL3/l/O7a4qPZCM8saGFVK5O24kHauSjk5uFd5iYkb3TKi3znOrZWDsNxELhe66e
D4xAWAq8eUe5+omutCc2CqhLUuzFxu2424ybp5OvNWy92gLoOrD6CexYVY0F5Q+rQV6QmMOHlloa
ErP3U1dh9MrnAf/M0ZSU9Ll9jL+spDBCe40hbUrjNAn4Jjg/Q8d04WGuVmNI7f9nmZ36P76fDqWk
Gomz/cVxoVO2MqequLMXRYF0+gx8WB1qnTgjmRHJAEgqdfbgky/NmAnp4jznHXljrZG98FazzGX+
C7ZcrFOiTB8FrC7b9XRjpr2MPB+u9QvAHvxHasCFdyyWaEKy4SUMPvkXhfy+pXCiNPRkoLez46VV
RE69TQuaC43FYyTpwzzN9CSnaYaLbwabJxZyPNK9yQamVDT0spxt9YvMMSkEMUhQV+Z6ispV8z0d
pFsHDmo/GH9CAg0tDYeGJDtREexwiMT/vlwXMnFqgszC8gLibSEtNKlqXypdP/WFBfsybepqzbMY
LQ3Kt63N9tx7gbkGIQxY9UfnqDET1mheYuGpVEgWsNzPRAVi+tj72Xfv4qNUy4H4XHc0H0O1Y5s7
uE8EjsJkdlnmxcQ7CzskyUg36Cj1EnLE6AZwJI+59+/oF5hu7i/MkC+RgK3dX3MhWqBdYBgzrpEw
M6KeT4uf4Y/XXywVBXNsG/WbspnQA9cWmxbZj8hHFzkv+jjrvmswe+W4vXlLfn3/e5jyQBPdkdfy
h7WSLXx0FejkeqCHEj17jtf1EFaRV84zKFNx/f0Jzuwo6n9E3KwXGvhFvePzD9JE4iOnrVoawyfV
j8tRGoIE4UvWq4F49gVutA/5DPVJo9gp5qh4TMvf8nBNFgtDPUAzR1XHuMyuQAisscj7UxkIByFH
OqHnt3O6qJHs/yClsD1nY1E8O21xzOoB/8ffpWZ9lw7858UuUl2mC6kPjT7UtoHnXBAnfYmK+7b8
kjM4k3fYhABvvWdJVB4wuhKK2jc0Qe7+BkUTx8bpn3DC2QDmymam1Nt2aPBtq4wOpbsFQPkYjAHH
epXMn7/Lap2e1LdK8XhhWPki2bWzeCDdTors95a6K2MkCKbykcAtnyvGYM9QmgIw5NN1RzMVr1jm
TvYcwMmU+ZmlqWosR+Bhb6/2hUW1ci3Wn7Sw1z6D84JrL+FEWnRURaXxCPZWFcHF/8FcIgfTN5jK
F8WvUfHEfB03xFBtJCNWniQTKzE+CP0ISPpLPfDdAyuQn14J9RPkGfY+VQEeDW8q+agwO2S0jOcT
cdREzE5bexbsAggVdZ3g3SmxOP9tY6Vd1crM0RBBJOMJQFggJsPa1PgKVT31NcEppQENCONLC0en
RH734g+pgfnRa7StBIDILodQqPtfqNR3PhnFyN6UR61gOCZJur8HywcdsZOC/jmXhid6cv09pZR2
+w1GQvsx09aAUyJZNaydR1CCR+jpeiJYxAqKfIP4fH0DdmUVSqRvPzZTTckDJwj30JSp/p9Kkfm3
7SkemoGLGCQ0418Pnx2mziNG8JSKKTBjwsL38nxFL/HTx4Ju/h3YxSrKyFcPaaJPEyWTS/dhZiYW
hv9Qo+ZJcpSx+0qRIwnZZmX6JEMGdkVK+A/xXx0Pbs8ypLJ7Pb1O2LMlL8U6gOzqM3ImsgOwI3sW
6T2NwxxdgJfGE5iWEMUzEP10lgJz0aBbdKrWUCvivlIwjLbrVn/GGg5+W3Hzz3S6eLUpzAAQphoi
9lOWvxqGO4Z7UNHjp90Zi3TVQX5fnt08+VgH1Csh5zOTiiiiEan2hMB61ujnagwC+OY88xE7NGib
V4gRLrVB0rk9Nu+8OjcB1zin1sVehvlVesET5Az0gfo04QUpXQXyzMgHQluhxWd6kgYzsY+blSiH
xqyA9LPyoWaphBcCMV+j0ktTx1w4c2mj92s+agx5ylNuS/XCOFCnNQDJ8R9Py0/CPdOd2XlInSbI
qhOZ0liht6B96OB4V2wFJBUUJ623ZdEFE8IbgXKy9mWsc2SWXpPjvUor7VjXY//w37M9KfC10sXy
F+Q/baoCcW6MVTUOTYPrXdVjNa24nLcw8qvUC8gXlIi1hGPLPR4Pl5CewDWuBOUDp2Nmgou1bOad
8c+TaHaK0QC0u1rKTnldkmggddqP48Q745n8AO8ihjeXMyF9PoUt12D7I76RyVr3sJmhOmAN4+tT
JA7R5t1/XoBdKlNZKMnU7UWwHHbXtwcqaGqZnNb+IV177vX6eoQGIszShtLG4/ogsfi3DH1fceKe
y6UkEt8UyCk/+gmbOqOkuB6XLkYRXd0VwmTxNeFDIq6uxpgRMxFS7wFVD0SHd017IGUxUMjnTxo0
/IpEoHx69v3zSxWY87tg7X38pvRODPBwwq+BYV1Frf74KDT3Y3okZWhlx5hbIpOYEMDgV0E5nvif
JPGBIOHfc6ZWbEJHR+XkMBENMcQs2/bbUJD8ykl/P0VUxnIwtNDqOsE0WsE4WIqsIJknREsTxbf9
xsC4cLgh0085NgBnLMtHSTXqih/9gNsZ1N+t7KgMIHBq9h3TJ7+aq5hFbGsC82EDTSQUpdnSQmxh
A7/jqvp+Ng5zDLONmK8j/g53Fwso9atKG3YMLj/mhCMfOHBUGdkMeW9+RHCzTXk7wsxU6glwjEOY
JuOKPyNvnenkAMxrsiFjKRjRo+HMJhF2iUfg6lCVwvYh1mXQIhnpdTw8qmcD/pA1VBF3Eo+z0f0c
+ZcOi9ytYbiIHx8RJ3lmgLGmmTF5zYQJC6koDPhm4GorQ2UmYlX5Nff3Y+ZdVCuo90WBt6MxzxrN
A+04FDXk+P7NRLN3a4eeGh1bfbrgj+5jgJInr4GbpaEiKhBBZ2XHu3PXI0yypA0yD3ZjaaMi9LBB
24UpQQVPc+APOFOpf6AcdO8hKRZXfQIh78xCT53aKpMsawIg9iP79l+T+6nugquohsEev28GxSS8
/KqynUC+3dWzlT9a7ygNiZt0VMgY3/X1SMW5t4oGIW+yUDgziap49oTLgZYdJzyoT560ZcRdhoii
H+Q2pmlb1DW6/GGa4GdLv+kICNlK/ILDNE13hQcZpKnp1/7Po8t3SQS3q1HeWfrikG2JkMn1Vpec
WnC9vk8HzHtZ8Xt/MbSnVUQXvu34YTzba3x7qnwrUnq8AiPkE+obC6W/5cJPBEwcmqnHJGYyrYqz
LAownp2c/F+UB8jn1ryILCYxKFzL18wZaCbQn55TtdaZkgJBEjZiVA11qbJOPw9FU/L3ThfufV8X
qPa9nbSGUuDBT2t0CwJy4nG9YqG63DTrb7W8urWGSJiw8cQBUISyWrhzVA5he2cmIkCl2Q6HkaVe
LFkZc1H8oGMlhCQKGjUFgmiu0Kq/JFQHZrLSRcCfS64Gy25p+oybDCJvh3p8AmePi8q48jiccznL
pmEIAerxkbrNK4S5C7N5/lYZtLbYruDAG1jdDilPPR+vEP3fO7iTXGyf5kFR8yfhXyZRX51923D+
VZwkRhW+wxx6eACk0RR7fNcxNwUS57uAeqHMfjbbtEQ3r5Fz/c/CYvvMhwWS0a2Z/EwIEpnlzOh7
dpP+vKAjEyzbeKDPPNDnTZxUF91vWhOvdBBaXuKIa6JIdsFt1DLP17DOsoC1al8X/BzUS3kKJ1zN
397yDQncIRoWU5+XMT95IiElbwpKmlREnHHdjLWB/qaGi7iLnjmD2aHkQ9Q0hSQVWxzFqrM+Fq8k
KGwTsw2+ZAfdC2xetX/1Q8BsBrJ07Ziz8uNYxWlxHy+RsM5kmz34BomNJr+A8dvvGGJ+fawL3QiC
E8pIYXTXQufsmb0JV4rlGo2LxhZE5I43g/gRu5UqAISMbSl1zI+sPLVdaVZAwQ/b4UDExzdjTguw
dgEzbvfbzOXZK/9572vSPH8theeQ+6lq0uIpSkGImdxXZzVRVianNbwM4qMPQ51NJs+oXnuOOLMe
6dYiAuCkuVdPdA/6EwXEnbU58nhSH4ucp6SiZ2VSVETb+uLZSK1iAZxATxN0erPxe6k8gutHQ5zu
eGlbhr6l9bbbctIL/SevMBrAKSchqibmY6SRF8LNzq1k7Bd1CUCdEnDzR1NKXYJoRG/qUm+pCK1C
Fy9FOZxFLWxNhSMhUKmUR+wjmAbQmmZmKcnsd8EIKm8vqhl2t+XOOx0QVY4TJeMKi+zLiIN8h1nI
aMRUzQbpuWi4k+cw4eCUKVSgmLF6GHmHaXzDEJv2Te0/sxfCe1tpXYqQJ+aI1egWcAxUL+i5I+cd
vEpw72X1steH/JenLnhaNWhdcDb+6Pc+p0BU9WK48Gl7//lhvPz3qQLMAWaHpTbJgCFcaiw5ChQa
AH40AClFxMa19Nsp2xpS6nwHP9M5eQ44EQwypKh8CiTjEO9v13mxVMjAV0eD5L7BW15qcqKKAc0w
MqLaG/6YpBKhKZYELuZ2/nfYWyY1L/KxQzwCaapXqUYg3xnRd4bbTH4Nh8MZE9rtMAlpkhiTIxNV
Uv5znYXpZ5DcePA3Pntpnhdkj4gtzFxtP9KqXz3XKe53yxbvBM7EAvFqFCvCGsDbGYdgnRHZI7dp
QJH5bioLmHsiTzUpVZbAWj98jrPzwJG5w/5XG7Pxd3NaDdv/JzN/ifbHgsqhhhlHDiqCyl8piq3/
aCB/4YJLDFFfKxP+T1wO+tybzjc7eSgQKlsYc8Gbsx5A0l+72GdU6pZRYadZ+6NEbkP4cwiMzMDe
JRm5mp1w1gsXdSQ/qnzG6r8hbI8nbM+tzgPmtvpou/iaOkwc2uZyNqQZYhyjdNt0n7L1hiYYcs5Q
vZ/iLv+DUe7qn8HwJhEdWqG3PL55VcO1eZ0apkqL/6rEc0T4QBG9h4+Wuh4u1VOK/3jjbTsiNHmt
BAaifpprQ51GAiP1HGRE12ZMe7OdXTGUC1Y/QJLadfCpMyVteNzr3cacOtoCnA5Brg2xDdn1x8Bh
FBh9R83TagFxKtEJpbqycW4RlVnmO3Dkt5DD+IWW3ZkBIaYEgT9DV2gsKxqONs0wZ0cPvKOryGHF
N34visIWLd2XBIKJZ/bxfZFCqwc3AC4J9sTKJKs88pG2YaVG3m9960hXkRsCjX7J3tFFJewb2uRy
3VsfbP7BAEwSZhSfmhmYUb2EtZehi65ZqIqQlqTJ2gbT6+f8n7rN6Ud1FM2kRjth4FkPwDaLqKbB
HTxuh5aJylerIUthl8WoJK6jdu9UsRE/y2BOl6Ivqhc1r/vf+3/1UAs3LNNz6n/geiiOIiAkdzKs
8OEOCAd0xveXIwfd5aPTxzEVmcaU0w2FPxbjIqDqrqwS4aRSC5aiYAM3Ca8RsA/SImrwEM73bkYr
9s3xZFlFT+2V0VCO0TMXRcUXEc3gad7XxhLA3cD7zHIjLpiqPfvi1RP+n815MJsNhibnA7iG67F7
oOCZn9p4J0VtU6YVC32wQKt//V6B5/P9ofNqG6tJpUQa1k/wUxsPXLVMu0UC4+fkweK7X+xQtljF
ZDHZZhWP4dmPk9P3bHKqbgfVkUGtfc7jPsx+uO1ZHB+mb/0pSXoSX7KBuExCyIYNv/v69SQVNpsu
d7pp9GBgMK6G71PXTP+jRlkH3wno7wDB5ZES9OXW4PUl1U+s+Og6UPW8vzHvsUodnl6umr+xF8B7
SkroJM36zpFNxezR6vxtm2jnAU5Vd1iQS3DX7Zj8nurK+ZXbpMFL/9eZTR8GDGS75ol6VFEXW9zh
lTsNOz5+u/fjAUl4HQRB9T7vTpdAjeLmWxwgOo5BSlOzuSaw9T6VR5EULLdGc6op0TWFIoi/izxw
SHWinppzzzd6yBuZu7eqRySh/7T0doq9S9Apq6/L9JoviwyQg9DZ+ydEj7HRt4lX39uAkSxyGnFn
O4uGS2dBcFyXWPeB2doHQB7LMgGKx2h59gRQcSAQmqko3r/X4rFLYi5BbZM29Qn+vVtruflMSrwT
fStIxGID/dQ/SCnBJ6HaAmhc2fB1VzhSOF7GnbuarxS2/IlqT6rVx4Le64t3GPAsbTBREShjk43Y
1qKNikttaS3r0ZS8F926Sgd1tWuFdMq0e716nNwDEH3XZ1v0ueqx7lp9S4/DI0ou/SHMSnTynFL0
FBxPHrAcxZhp24bA7Kr7E1MmzSQ4HUEfVQAZ8/s2C8Lf8I/9iBUTbW6gzZdCGX4w19R3jh8oJnGD
mV/0ak+kkwvvX4m5/HfLpbPayY37JnGEsRr3zl0jj4XSYfmGpzvcMk3B6D408slgZvQZyShITy7K
HtcR2BtssiSUhrg3E1T/+ZjTENV09Tfnfwxy3BzS6EEc4Kv822fjhHeCkPsdS3KIZKqb1fm1SC1U
xkfd9Xw9gbKdGuk8sCjnq6zRLJKCwACaan+rRvJys2tikRuUzrlvZsM0j+8Dplrev29UCs986D1X
iRYSuIBQEZwzjC5jsB0pxN4mUKV11xeOZuHiuGLkyDFTlKPPlwiRqKeTfAaoawAxfCa7/2XL8ZpH
xHcl5Dg0ArGlICEC95ENB0VSXSVOvPrrBkjemb/60dfHln2iNif0MpoiP4ykOUt2o1pKC31ub4AA
kUu5kuyD6l56xSgx9StMeK5dWsKKYYqbLVW95LijV3zvre2XfsfymH6K5fXIapPo9uVUjnK9XAR7
kaZ8aRnrCOIChI2fuo1aJQWRGeB+6GRxynd1YkUhXeVhzcYhPJO+poskKI132ke1TaBkfOhwm/UK
NVE6zHgHFSbdzJerUX7RKDrHdPMIQGRy/iu9wFLcKm35tDUwiB+fF06ntPp5qXPGEIpMv+gmqJHV
2T7N2/ZNsQdbIvGNs/3+dDVwARM74JLES43EXmjKsQUXapB/s+5V9nEnoWzwDU6zYnDZy6GQ2U3v
nne9xs4E2e5OVwpST+UxjVj4DQ0wTjLRuilSvNab4pn4w1x0TbrCW0tZIkAkq50zh02wkijhBznl
e48DfJTI8DrMi/n52x6CtU+sUie9cLzFrdIZT2vrOxylLrbErAl/A9M34QlCWQ3twct+rFKBstoD
nlZEO4y8kIrV1lqiJ+gbsh0kuO4LqOpzY8sAgmNDstwH8eFYn4W/bVl3EczcvFgY1VRwDAcMmJnq
tR3W+CBwXsWf5WQFsw1mvBpDkx2wOlkB5+XLbpHG7XWH05+zrH4Kw+AHxCF0gcZr10ZDbehkoUjK
5L0e3jZnfZsUS8gK1FN2vgAJqV62XEL1LLtg1ls+8xPkpHckIzpmlgxfHJo1eK4sN2/fcK9OOtk0
lW1bki+rpY5cqjBci5XO63DWT7IPq5MeJ7xN2PF3qfLrTVeJFyHJvGi4z44210tHpVrCFN76KEUy
LqsyIe3d6o86IJTJ9sgNZ1+h0073e02hvdm+ulz5pBY1/vjLfKFR/oo3CtiiBX2Q420gCeHQSC65
flQj4Yb2FwRVApzDiC8WIMO7dIIKBIxVWIpzT72aJJIE7j0CrG9m5uOgexn8pfWOMVpcJrAh6J9y
shWZ5BgX2SAeyvCEYIAxjHxvs5k7zrhzEm5NC5SvM41XfnYe3LlKgtezPgR+EbN/mjq7hIUK0lmK
nJV2NkjqVhan9v5JnhQECX839s4JQc6mpXpsv4i03GqRpJ7B8GzcRmNqwEUl4q+9bcQ/jDhWKcg6
YU6gnpf7WfsMEovUu053oqOpkAyeG6ZsjIcr8zlsV6DZZJmAosG+EcKsi0EZLJ8ntQjPbCTxNoiO
IBXDxEhD5KKlGAunt9aKL9wWjK4L7D8C7RbbyDU9O0ZOe9fc9wNw9rlGujGIkxaMgmWv/WzOtIfV
Fx/EZ4DzSAYPsTtCE5tGYP08dwOcCFYeHQmm5Upq8U836hnz8o86EyVtCNrdUCVc/RJonl30yrcN
wARPBs5pYHiyj6pLGfXr7MKqhf42AU7EdXJTxiGEgk4cFjSbL51tgxcg4VHxjHZUuAo3gaaaDmSD
juWjG16ks5hoazeSn77EqwlyK9eWZiHFZV1YcyyI7uuPYHXSAiQ2svHHjpsyVSz2P+CAUX589auA
SmoIdJEwcp7dnc40Y1MsPok3iLLAtP5uC7QkMXg4N7O2IyGEDYlZ0B2zVXnVL3gblP1wGMEqRogS
JwIUvP+0pGWOTvKRA09T4TgEZTGAL6oL1/LaGw5M+j6qqzxFbrQeJKA+JmV9CFvYiLjK9vQWbFbd
ngu7D8z9RKxKxoEkQ9CYxVPqLTIR/EsXnlvvQgcFB2p6p9sQOEJPA2ob/+HcBCa0SHiL8CQy3af0
pDR7jxF4PWFrdMRxwyWDnIVWsg1vV4kTztGlk6y8GydwwhfWjoBz/aepyhzgGcIo0q6Uv3wcnUx9
KCAKYAbfG8sDYYkYGpCEHnKk95RolWQzynKapDjHTuHzZ7KBagFdW4gBy27d4+SjZrFZ7gk/a9rP
++6HnJJfuGpYCOPndalkZv95FoSSXFfeUnpx+9at+Ebq/osRJ4NGDg79nUl4gdG1ugOLC/SIElWG
o4J6l1cr99nt4q3bq46U428LTDAqKK+Mcs8txZL2bC2VHRDyeohCrLretrz2LIzx5qQdoYhF+V7N
am6wJIfv71YagchQE45hpxpQYLWxWNiKPrdXY1KjOuMv3vTQRNcFUuRIZqmuSp+tYM4ZK+xLvfiJ
CFUDmsq+fgYl1vNcZlgifanjN0iprLNUH1hZqZFcqlEzsEanNeMa2QuVkY4QRC4J5Qi5xuaysd5Q
TnlwcFHzBUT3nqDZeQKNxCDa936/WPGj1gXmcXF9dmHsb4BF9PMlhakFftttNoRKylf2YQm4aM72
wkT/vEy5kJTssuPqze6rwOG4mceSXFYJeNCesl3UFNHfjXBAfUEMa9SSeqHEgvFpSZjx7/BRr26g
9USaxe9z7AEkssfrMryaMpeqA0Ez86QB11JQgz8dExZNx+1qhB4giHPkVc1W/58r3bLx+9wArneH
TgwPJJaR5lxLTVmglxSDjw9m6tvIpmOcDbxh7CGlUzc+mZaS5/pgFqLdq1WLGOjJnXBQNlvarnXq
uuyL/5zyLNUhCSyn5W0yrgIP9Gsh88abEk4mElMT2Vkhf+3IEV4/Ar7wude2/QYB0IM+YlpfN6P9
A+bA48UF/VVNfA/hFxRViyVH3H6rpbrKMW76TW2L1AtboRCyPkFEsrAqa9RvBdfoGCOpnGgYWwU4
TUDvnrGD97TwzE1BMRWmCiI8CPDibhI6dmzE1zGLn0Ee2Th3oZvRwHnjrD4Esp9KcXtSuwJ6Sgss
HaC9Ys1erfH7awqHmiv+76CeYuvA3ubHz9hWsMDL0qhELA0vxeCMYNY8uQbGGiTogCA7AdPRLiXv
7/dOSoizt1pbdU70gZ8zt8k9VxueJm/PNqVBscNpEhdL/g6oHRtRIPB6M2jpTrNw50C4jyDEab0L
n9LXljBUfrtswcmWXeGz6nVO9IlGp7eDgj6aUjRZerumNH94+LTvTMvgfHyOkcqFCX2/TmcR0RNs
wP+9i/5oqt/e0w+VgepCN14I8cHpxMgs3br+Rl9Bq8jzOkhHlFSL6aKrNzHLVMODqc9NXhnMgV/r
wzJ4MTAGO3RN56yE3RHeeeGv9afXQ6k9LTEStPbw+gpFzIXh9DlONYdR+RcPtfFkMQKJefduJOG/
C4KWyS3fNpeHWhuZErg8nfz+y+UAGzp/m/YUfdSeNG6q/oeaPffsoJ1tCt7zqJdd++P+yX6Bnqv9
iyacQWjhNHJfj7VgF8UwMfbUMe5vOK06/rlN5tDHP688FjC0NJD5+DKQzMLwdbmSQTB4wUAIz+IL
85rLcc7eMctrF11BOkMNv+OCk0QUsjFst5bX8UbXdZ+0gOCCnWDDYtl4Wv71WhWm5rt5Rkia2Kud
YB8qOtxrSfsDzkzfzKLQH9OT9bXuAQjgBVy3jOBkmBNdFLySg9WVEkzWbsbNaQ1zn8FMvnSU0tCM
2/FKERpNtmmiCZ633TZTUC2oxTA5mRHB5Oj9h6SwAUgAwSYKgKxqoqONRLG5U4UK85OQhMI3DwsC
gwNLrbIsD0VG4Y3mvj4UIeFZ/1c5utC32a9yyc/oBosTULUgfAqelt0sZlzLLh11o08N8Q76YbbP
0x7r4hzg9U06Pis3ZkWSWYag/9TBKhyJ3Lt0rLDS29JGl76bps/N87PihgFdVwkWz51AHhlYXLg5
dIPhILR2YrCJVKH/5rOAMD4xKDfCqz0n2GH3M9NtarcLgSAowCh4iQX2LKpMoDC6/OAhtZSwkw2X
FPbNQLMbLZ53U7+3cyJ4qbqTc+wOdaM4R6Ku2iYw27Pkmo9cz2RjUOOFv+ZUBUOScL11pUMRi8t8
wZgiS1B5l1/r9hrzZXmI/fiDeo5eGv6YFjWSSNjmF3ZuYOJRBAGQMCBtgBTRmSVMKbhhCtiA2+Kr
oOTnDxDK9sQBYwvUL9V5N+UnDkQGU7YavUrT9gJx1xNww5g6bKKihOIMx3ZS7AHG8YgNzdiFPKaY
eKliF2DL60gJ6feQxx9KDnIj4qhCX/SBce09X6yJMmna73xaeNnVc8bZaOMqbGnTbKAKWrQffGgy
9cfrwlkoiqqHRehXDg5NkIpTU5au9utYaO3M/NYSVt4CAy+cELZb3VBvNC0XmG0g0uHeIbETbSh6
rivv+tgwIGcid3rOyBsMBQwOnw1K9+Px1Pqkq2dLzb2dEV5yu9m7XwfZqY0V6iPpNcK4AQe9UZu0
Z7UKI+58nn+YEwDj5TT6iJH2I4lxWGO/FLAstBxvWKbLfYrF7Zfg+24TB52dHurp4Pz8kOnkVql4
4ZSSDtgrNvwtmQkwawxBTeiU0f9bMKhm3t5g0pZDz/EftLgnMxffdyb+PUeP1E+dovB/PIr+M+Bh
DyNGAKi79h3BoCvL6bZ6bG3AFQGGoSGXUzpeEJntA82OVmzmudZNE2pZOKvg6PwtoJ6tR+4+jtfz
EwnTFmsWeQrYlskOMfn2R48JuO5mekvhP/Rz0YTovqAApjtVCecT1gQAoM1I969oKOr3U1gTcMV7
y84+XLKATBs3BdFLwGuVIM7O34xj57m4mc8QarLzkI0ABNWcl/0mCIjP7WjkNnoAyeKwyGIN0HHW
2XwqWwelGQpNgPpF1fKorJR3icVHNY3fJygCoW8t2mk8rB8i1h7uyuLf/zfdX1fNiVkFcNi2YBdf
EhO4GYRDxROr+48szo5L+0AG9pPgTOhd4Z/6JSPOmoxuVNT5hHU1jFKrpmWIYh3w48ho1ddqNV+n
2Z7gPQ3PES0/yc+s2eFMCs917LpFFPHsRRPe07olS8O70MID+RJeIJIp6x4dYIfwVuT0UtpCBO/s
2ztL/5i1sTVNqxgG1KLFnYKWT/hvVnGgWLmySr++gl32FoktyKeTy6lqyM7Je2+wYgFDYTjiwr+s
f94fDN2jYxEsevXBzxqFFbZRcfHgkl+QQjCeCMVEuHKTSU6IvyztSOpFybIkU7AjW6RyhEvOTGDs
kugKlwdsLHYjUvo9si3EOwp6mJCZMFr68NtZ5tqdds09eDq4nJdLxS1sNTjp8R/C092GoWHxHHe2
m4X+l9FAnZrETVFyGA1H0JDIyz4b0kFl9JLHh6hRX5AH46NWpY007nLc0M3Mn4miWN4ysWQb5ht2
om54rrnl3yMhMC5weghzp/X7Djj5X1CVNOdbTI0ewxi2WFCGBYHBbocm0paeONPmXa/g319AK6cz
XQzjXKT1/lFdPQslEee9pHGxhOWxHehxDdxQA/2d8HEJGBV5mIZFmqLCfXUXKUbYXdp5nzf8JWAD
zGierjEWwTj291X6LjybcFDJo6wWFvEhn2qCw5/0YUaq3BM3ZPwq6/NO9ewNjnTvmpzFaBsA6NnM
fnqWflRW/9wMdsRY+o9uqHM8cKY4yfExviWf+VKojuWTQ3IGxJ84KyCoyJGcF6cs1JRVGvhBu+h2
vo8+COoiPDM8pdaxaiOCVUkxsaf8r+TAWpI5OXwsJmyF2DaCHGcPrBGUZNSt4UmcIsulYVHT2wao
94T8iORNQozrXJWr0NbCqWHTqxpfM+sYxCHeLyWFdrrAfX7f7G2KnfSs4pBni0YaTHJKpMOuNHHb
DdhS43kS2DIHOqRYFE1tidSwnOjAaTWG8vylCWgAyYWUHqfj+C0U9xD49HmQeHpY9h4QW4gjd5/o
bqUJxu/SGOxs756h4INdLI6fsuAH1EYPDpd+6mz0ymz0tIzYUlX3HO4+3r4OVR81jB267XhJ29q8
hlw7nmAjhszez3IWLRpXdWcU+1SrBtHbdkDrrgLiiGuhBkXYiId5mr0lrFHq3Rk7NoZ5joGG9dvV
5+GRaMbFYPfoJSM/+knZDsEZBlnbuZ/at6ijMNdZ1Jbcr2afaiRI1ck9cqj+V1NzyN8xqPek8ZJQ
VFc9+q+atedS1ZLouaduZxNtwp5RLhTe78QM5IPVQeWn2bQ+26nwEbFsDvjIseYObYf1XG9pMdMv
Ig96x1bOM0TqmTT/9AkKz77sMiGttRKP49y3ZvES9zAZA6ynnYfxpGNZnJzukGFw3LtYjXkyABsi
BjKLwPM25909E7Cp+/25Omo5HV/VQ9l/5iBsc+RsdjIMqj2v6JYxwPS40GbYiQQnzmndqzFngQw8
q1PSm83tipdncrt+7jkJwPL9zp5X/YWAPit4YLjrsr9Ow3ULc4U6OCNWCLRjh/KFGrOI53X6UmCh
VytVgzCPx7hw0XDyazBHqlZ7F78pQiS21kWioXT9EM3/ui4cNFFb85SuypD2QQeUo2oW6GpuB8Xh
zZULTiTv+TobiKmvGpTlLGg1fBBn9Nrq12OGomP64hIZhFw50HPH+/TasRfPJ1ujyYnzu+9BWdzV
U6PrRbxzbzGXR4XJB/C4xvkj5Pn3/1N3FJjUgTnYKnUvfi/Wvn+cv1FWEWg+2RxHOlKcENoFyZX9
PHrtveiD8z67CpIw2kO5uP2HGtIfZYBMD7/Xyq8yFmENr0+tkip4Fp3+OifPWlxBs2Islg9US0TB
SjLXsE9Wy8oX9MJPkF0OMO4fYydpXlLKk5iGYx/ex96bqW51DffNdVoCz4mwLxc06C5JCLWMW+3x
xCkXerXFdqWJp4ZaJ3J3eyymPm9v8CKr0EKT+HAb4KDX89etrfpZaTxWqnq2YspHgNn08b15RdQ0
9u5tu0IxEFZkzS7NPbwSGtAmES3pHBCivSn4gygmP0titVIJJ7A4220LbxArXg1ckXF5STxF90xS
Tj6Ko7ZyHwzpLJPwUDkkIS/fta426VHGp8Pmr77vkuOs2DvT7YjtSVNQxhPkE+rvOMDVgm70uRpx
2UoORG32w2fvqrbVqf+WA7dYWjLqYhackl08Eqh7MVwxgQp/aCtdefk1gIeE84cVLxsiFy3cO+Av
Sqbdgn1kOd6c/d+t3P9RkTFkimKfhaQSlc32K8Q6Py6lRDtpaLxZH+lBJQsyAZwUuxjOLjttdlZH
CK/5wMD/EgMCEonxoeqMZl9BFPFipgvimwgH9IVv54t04Ckx8SXbpVW3rr6iXaMeKmk7C2weCFrr
DmBmBf0mYMKpzCyEzr1PUV3aWDNy772bgL5kG2LN+qt29/gYL+JXlVTAaeFzczU9UEXs/4nnOCjS
t4+EGxCuuE2Qd7QyBtnZ9y6128wvO+5bLcqC8eflGxKWurOVlI6AcQoCnNlC7n+lORLQGReUiuAi
ZEhVcSbbpoZeD42bdhb9YsSfMyLEHyUIMf1BqaanRMttvU6kGzDWfpUoO8lyLcxywrSn/bMA2raB
MjLAE6F7ppGKnGQf9bwt0PnsHsCmZvQHoGw8EV8j3X8bg/9rWJrlLHfFuIErbYQGxgljDWeG+H6O
kRX+m1XjNZHGCZyfYMqEAfPKzNmeDfpM8IdCdJwPs8Y2qlGmFvcXa7tM7hsIgG5cKlAWlbttxOyN
VzqKV8JC4gx8Z2FzTKtJ7W9egZTj8Sb5KHvVmq2SjnwGU318uTr/vn5B+Uu0P4ttPPFEgKCV06wL
oI7d9WSOBvlHIuM575nt91Z991ByqEYGsF9jxdwAluDgTvnv9GEjlnZCzalS3oS/p8OJ+/YNwRIQ
kL1OCJBq63vpIawd4VMTg+3CzDsTI9/L9QyIkeCdvwHnzp2cRnk4BmPySyQqIBeo6F15+yXRC+ct
1kBQYfnS5vRKeGxLZFD8x6jy/ZXB7eWok5zw0RakI1u/N+igR3fKBC2RR6s2S7YS7U3P5ENVEN0A
CN7OjV57yl/M4G4bEm9UW8e0xB1KJHBgRodZURAmijubF2J4L2M4YepE6H5MRpxOSuvjQBk93VOv
754vsVWMjogyDd7omvs3H+CaUUR8Vw9481kb0JNGXOvsBM0XerJMK9TDupik6e77YuXL1LWpCNDp
NsFHGdpJdOnH0B/3o4WA/M3Zm4QRpZyiOd0kqdvp3ojNnvWNso317Z+eyT4b6YXJ9kcKJAzB7XOe
WUgQCVWARcFdSL4T7+9jMq/TiAcV4FF1GlekoDlx31ayNafUuOG72u0A7nFpbDXiO1l/XSDco7W6
ckUskwoY11bObcP6UYDYb1vx02UW/Hl8PeRBDLEqetWu8PBnZwaDG/I81P9ZvPrFMkYA+Ch4m9me
5BXfdCH/MJJHoA54SxViFxWn8gfX5ydWVUvnNpb6voovwBpgRbel7srJUW0sb/YUUL5YRdaPIGpa
BM2Li6vQy+zDmS7smbUe1p6dtDwh5NYBy6kzYzwivTjQQOl1suP/WZC/2jIgZYbZlHljP8FoEzIK
rUXpMQRO23SuH8OV2Y0ZpZfeizJea2kgLtgkXrACsp9COZW0K5fI9CFPhISm/7MapLGDeavZG7Nb
EjE0wWbYAnsHSB0Kvp4KoReEn8AJg5mUHv3s78q8r7GJd5KA5ngOYIFh4drECdaVxqhfyCsgfvGj
7zqrEnCW21K/6Jf1JPwHG8XwiL4TsvpuG7lj6LvHc/c0twmjpip2Q5K5YTlDF7G3i7lZWz5v0A7Z
K3btJllA4+/hVzUNpc8ireKx9r28d3GNO2IwLo6STdEqPitqJfUA1UT9SabcKIk1+dmU6oBowDCT
l370a79aI/BfM2QLJLIaHH/letZuRWY4lEZ9/eAsbOg3oW/7zJRKrNRfzEfVUqEs7rPHR7WTgNyh
K9HnZBsRbJcVAj+4gEedVoQ1Zhj0mEVr+1h3rgscu30KcxRtytrm2BypBFJ/I/4xhQEugWxhWLFO
pJfVpITGaHMSfsMtORU3R8t9zB0StJvRKYv1Ya162GDN4ZGeRISi5xC0OIcuUVqMGNhRaontSJaK
zWncSMVVKEOWvVNH/8V5rp+rSJoJU/3bkbaInB3B4T0nycU2lsskeNubXbmtEr5kPmVQPEBk0nQO
4RAdA2Qw5F/fP89uxA4g4X56Cs9RgQ9gwQdjdpDwLFWx2odEfX+z02x7OvdrYnt0Am7ttpYOPT/l
zzkFwhprIFd1vCbAZJzwL5Xh334rizoR2AJtoHUG8nzx+FZ313UCOHSvMcAa4dLCupA8h4eGvVXZ
d9IXROHQRp7UQaGZcWR+0kfV6ePgPjc+GuwdwKSyMzqK14idfFwE1AWyfM4Veh+mrfu7XI65vZof
2vI9M8Axt0d8nPxvloIPgRt5Ebc32D+I79VFniDr/zhS7vDj7YxZx2TxIxciDaot3wuXNgz/Mfzx
nvdlPIddKy2/QhkKNr+3k/VbWp04IxZGOr+45Tqg9Es5PQWsIxgzohrtT5QxmVpIdSzYK2Hr9Ajm
91oz/Uvn64HJUfbWAM33yAEjVtBannhtOzZnDViUKmWCMIqrcMW1/4FUQvgPzo1GZfjOQJBgriF0
E2PqtuYgvjSmwx/UcF/CI5/6F9wsDxwJ51XDGRKtAAiTGaNM/TsBkgCUXq2I7YIYYfFHagVn/r7V
vUDvVtv03wRQ9NzSThFjj1w/2zAuT2YGlrDH72nlphw2USu5EKw+Mws/5fd7O0pvOid63rPiiW6l
uaUjZshO+985P40IiewWQR/+mO1yn6B7UFIcqhYeX5Zdu5cUT3QmjenCreA3UKJXkaItMNYILAeW
18C+gaEA6ODW1tOOMZXrEj4Y+bc/RznkF7ywZrmOemyvRb7OkctjLAFHcLhdOVJGJ4NYPt7Sc/vc
IA0BLtlFu7ulECwmOq8Bw3eywsaOJKUwCfrcXr24ulp2+CAzT3DRk1KE2G41fdET+ONu1etAaLCL
UowMXF9Zsqhr9OE/i4zhioh/ewwVHvp6MZCR+NQMtEadQBn5BhlvlDOE79ij3mIlsvUE5NjmEyle
eNRzs57bAbyNhCY8OMm0okz1ewI6Uq9o3iWGvqssfISeg/k47xP8rESI6iHfoUntBiQHVAeRYd4R
qwiHVPvL8LZqwBwYK+MxjEH1tRdfDaQvWiOl84NXUvX0OIejc/Y6iQ8e0eMzjXIl7yCxxWhi52OG
QY9jdLc1aJLRN2SM0fjYJj2jmrBI6Gl7gY0KZdJwQBtOMeHfnZrt8bywwfQExHC5p0UUVA6rbiDb
qEeiIyDaR1B4R92M1HaBqjdp1zokxRv/FJ0RJs9SfM5POOc8SOnJ+Vq7g0+2IFVqz+wuMQVGwRbI
53xmrp68U4YQDZJb5uGP5jpUkdFBIxmlxGQZYg21whlqJ5roNhVWzUDZxzNqxSRmOnjfneU6FCm1
hFHZrrh6Q8Ljln5SxHFiXgFMyOALvonu1X52Qv/Gwntr1y8uzrvQzo3AoM15TSIyspUyjvFgaeKu
Msa5GN3GaBZ5qNv/zL6Aa1RSqlOgYNXd+9Epmj481oQIBGV7lEluGl0tni42Q58tpFS7cL1DUDg1
nf5l7ZITmVfapGbO9o3UL1isNsG0Kfr5HZc3ha9xqkRHUFRtsSrjioW47FmDyGDzsbFqOpKlWBNU
1uyZZby+hbb45niGBRvsjnL8a09oX5YqUCPIlh3Q33C0LxGshWSJMKjdP0WDSW+Hyf/P8GxtV8aM
BgrDkXLIicyRg16+g2KPh7eNAztWdmIz9lrRm1+likQKQlAtbgl4MlUiCaQ49wuM4OYo+0Mtn+Hk
cwpXOv7M7nMOD5vSWCi9LdERHKu0Qxg6AQfTiqF6luRYwDic7yvx+tIyiuNK87tt/Wx2X8Ma5/x0
W1vvhu36V0MqLVcM7Rkxm2ig1Bqyvy2hi79uJf6PnTU7rYXnLVEpuwP77VB/rUcIjngZr+jz+cMz
s/g9WWyk4DxTTLAsLL15SFbrTMVqv6vArZV5kmXu8g9WHiAoOLuslEfPu8/9SYIYP7Ly2t7WiVMg
Ri1kuyJL+Xw8rqfSUqtyKLx3m0HvAP1QanxuRYETM6lvJFAxg/5h1B9dxqq4IgZaT4Y2mMMI1uEW
2b1c18T6P8P+eC62YGp3mrsWzTmlUz5YLHAytmSL95VepiEkJIipSxFw2fji4p+TuQC5Tud0p9u0
2GpG14Qm+iJThC13pM+j1Hw68acT4unIVFH+0oVOMtZQSVrmAP9W2l+SBjli+XMJcelRxIthL3P7
AfI3BnuARi2QwWizcnkhX5NHE51ec4+QeK9cgFAp3KVxUcocUHOg4BQwNWLEQCkzEI51j8iSs5SS
jUH3GlVcOjViUH3PXTvVb/dEhyGSYe45DPDt6OI0NDZ3a/Xf/Ck5DEfxTSVd2rBxkyIHv3PN5eSk
klRVa+mRDICawXCyXxPVp0oAapsQdm8tGk+Vcq3/kTE7C6jUL/ZkQ5A6E8PC3fcvLitD4QLDd0Ci
RpfWKP3uq7ke2zREvyb4k4An4L3bCfAEfi5LfsLPxHJRA0QSLUhnoqqv5bc5DpJnL0XXs+O2Bll0
984GTPyPVMruPL3S5O5Ii4i6zOgQFbdoXY2U/sxyuSj+2qKG42JkjVhR5TrHoqXvzWpYO2tKMmlT
kV/GIViVO4RN1PHXZxMJvwgfY0GdO5lOJTsaPTuYTV8q4xJfeDlc316iNZhizxOUH/d/ts942h/m
mgZMRXFhpuJahhq0tjyTD0b7dRm0BhdoMUESgTCS/huVWWBzW2106AfiZkUaxeQsge/vFWYqCxS8
PmVr+wzdEzweJ/e9Pcl2fmGTWub0WWpmlR2PlM48MeUSmP8HBwicDp01S/cWav2B9yuf9HZYm7LT
SFfDkf672tBJSNcAZVa9Il8qh2BHtSLymsnQI5jfvMF1ZOpkJKBSQs22/4ubTTb1yS1XNBpL3ugL
pzfSkW3m9R9whXi6R3LF/Ce9z2B6T6X4yq6NQope3gyp0xAwvhX4gOGjBMDQEie4iojCKnUpLBU4
9yOvCVIVNRk46IJIwTHLk4z6CRfnX7K7TqNivvYv4neD6Ah5XJM6s3iVm/aFoTxWC+HM8xHcOE5e
r0FftATGxR/eR1PMz2qxyHl4UOFm8Ukb+S4fwrDMooPG7q40Xo/xXLUVrfDw8Sx2jOb/Cqt/Q7Hz
vqK74qRo3RLNjKHAwaJ1liqt9shOG35YfcC7Qkt1YhjdNX9TlzGSgd5QMpqZbpo8rixameDEQoUC
tQp2L4NIyhXM26NI9QUYJndaBOaZRca1dnYYLco7vGP74SqIVRxt640I7PQHFLog49FZUpo8RaHs
p+rUfQcR2EDd+78Lo0zELpPdw8sjQs2gvNTXkseXqy1Q+25QLe9c/BgCxHj6kmVZDsmHXZhrRfX9
rQv8ozYIVAb37kHD7TLa3qAC04cwtC1wiwZTZTmwKUakAVnl+YWwm2vwDy/Kc3dfhTsZ2ekkq8uI
61y6M5qbcm0HvJoOA6MYcb1Jdfy3qsL4RDytAZvCxQxMBn+9DFZOyvgTAoYu9RIs2Pomw2PMhhbY
DqAqsD14aZJ6z5C1V8a20tMoebs46akNaGeY0Yp5p8uCoAn3DH+kaJxOjO6sW5s4WeHn3yAvZEjm
oTDn040Fsv8VBVByGByCHU6NDW8H65EYswXFk8fmoaR36BL3tSlLtYuqki/wr/O/Rwl+4S48Mr5G
wssF1HUmkH/2E5kXEt3KnNzB5MWQ6csaH36qLC6btfCPV7VrzUtbRBV3CQZsoqHA2fGK0D12/a65
wPkPUxvWTcXoGC3FSa+ayJ0fr7FWpeKCNNfvsZW260oWcWZdtByLObCSRjXelDfifKA59Z3vfrny
t65cfjaufttS7BeoidPEPrwMbR+qi8o6yR0/IQoWcy78PnAdU1mLO5ZwYW/cxatMVfn0Bmkcmnbi
Rt8kH3kRm7IB/IHkKf5xqXQEGrC9KFqCAaA5t+/IU6YFyuU/MfrCTh8eAtL9dyb3xNXf6iXdMcT3
NKaz+xHL1DRnCCTM1pFzY6Pvns+Ze2HJgR3WqRURZZMP2mPpLkdPWNhuEAWZAmnNrKsw/1c4I6oY
eSAJqDDkmX4PYMFrID7XWhpp+lXtqwS91sGmMuRtZpIESJgD8ow40wv1P/RuXR4PLFmKRIW7W1S/
gao7NW3LA0NigYJ0gJ2O/A1N2YLdY2yEsfLyc5+wBY22Q65Sj6r+O3qMzT5jbCn1ZiM/Fk5f9o+s
xM28pj35CXjCE1zoKVY6fVpZnyTN8YqQFmSjz2kXsHq7qxDkwwLs3KpLJnMP2hyIOA7ztqFnI2OM
iMDZrpes8LyX3cxuUeGz8+E38xxSuxtfTVb6OqwtqwSRyg+06JUX+dXP7ks+5PxH5SeNnlEJz7Ys
j9j/w5YAa2/CaKVyigIpPued8zWQ9zCxy17h8VFA+Y5aGyQSZgvRSO8JUvtolHEZVgljdmfo3mJz
H1rmodGuW6kptWDURx+E0PyjxaHqJxl4dDlCC8n8G721L42T/PTIkVkcCBVL5Ux3v8IMqXCNfEqm
hr77QSvGZmOSarOSNJ7HDu/E20PxMv2uNk8WCftidhlj+iC6UIKGg9Cw/oQWj+VZUxPz1wNYUrJV
EAVraBqb9+v1/UmbR1OUZe010T13nru68lFESod2Q5bhTILn/KDdu9g3xHHm2pbRLKUy1aFgqH9I
nHlvHkEMCiNmRWPApB3lTqbWat7RaLZSFeZ4Ul2aKf0gpaiNFDSZo2xtCPEwiaRKvG1go+aoCqPy
qd352Gf5yqUY7jBqKpnSk856yufVb0gPbPV4NDSBu1pAPF6i+SQwSffWnsx9qbVVTSFKwkFbDRSq
Qb/9/XzSwFeXFqGWxwQOX/XxnknuOdaLHg5CbRRXRoz8D+mFkwQ8ZqZkEXZSw7RbAdqzIRACyrqV
liB+VnkuhiPIHLH/kktlH25PvSPRTC3aEVWuZgq6XjjHJbogpzNEWhZpQNxqVo84JA5vrYDi3hnH
DRRfqIL5K0LoAUjzoG2HzjK78OIZK7X+xKzEQMU8gRGCPMx0kpj7MKHRbOLbBilidRbflNqv83/E
Yw9YdVcpfVT3pKP/voXhBTn54ac9zyrehz0PnyOH13nKHGY2hxQEaxRj5YH7J3VfEBRrMn+MUgf7
ArYGFBIQ5D2UmF4sOWpb3IIcSdlhMwcAvNnFgI4FQkZWggYFF71ICpwgebgKz9CHrIGakVPcg0b+
uO71cp9N/jfh2W++kCRnsjeRcf0zCijefe21VDLvuBYEVT7JtUS+xmv5vmaTV1NHQNfY5LE7SVnT
ghJPAzoYPF7XLF5CF89XiD7r3ewOBxDWuY4J4t2wf4To9JbW9JgxMylRP9ZyOEGsg/Z3B7XBOwn+
Ew+yxGWKkvWefhu5nNt58lV8dyErbne+LrHWmB3q4kNt2vxwyDTn6/JRlPMX8DapVEbhp3OIgjvy
1KJ896rq+OEazTmn/8xKBCB73S4CHpcp5HedSsXbjCBIftI+iGLlU2msROVB7VTi3tue82AFbQZs
3idtM4yvakZnk62+IHB5Kqyt3zY6479sws9nDV0xoPbjJw072YVocHe8u6uUIN1DEvRYkEbnurKw
c6I/O2UDlvU8USpt2SWYYXoceFcENGb1ydn/EPnVF4lpyDkzEDmEfKP/pAuVzR3YGfWef0N/VrBc
h+hstpa4HZVj3tDdEiUy0wCL3iSm9N8vKL+N7RaJzHzREOcUXQWLUiUAMD7Z/D0nFvQE5gYVFdn7
YvICMVi3UqEzzF+Hd5dHIwZMaangOuIeOT7hPPIHIa1TFgA+XePIT+Vx+2j+6KESdZ5hXsVYv1P2
tZ/HXGFynfhezU4gYgu8dEJA33UnC2q2W6XPj7mjJ8I1q1orRaJNJ8PUle+PaRXfKJG5py0YKNcK
JxVWsIsTm1Ww0bdLVMa0KsEuKqspLyUbLBe7WT2LfW4ju5GluV9Wqx9jfLVfYFoDjnME3oy4/iKI
jvKtEfmVvb7qv2wewq8nMGCRnRJ1ANgW9Xtg/38qD8dA9qoZlQ/eZ6m8qxPTlopg0pR7f3uNlAql
eEpYMwUJqnOEiXqYwPlTB20u6VLip/yogw38QmVv+VaIcnvh9gCcpMxdJQT4xSbyxaN2GqdKMPYt
7lDuF1FWuchgmVeCFoYPhlSCdLRt99SzOs3UC54tf7MwnHHNpTRSTArL4LG5q6kItQMiWlm1f7cx
0mrYEjljQftncU9wvNSdZ5doMyuURyj8N28txX4lT/i/z2LovFuFCJSSMPJWv0b64/gKvKgIyONw
r4TBQwp+RBVw1JyHbfGD+npdqVCySqoS/LEp8FTf/wHfXiL6jVf1+mUuuPkDliev4hdV3xni9Fi9
4sbRo0YRRFRSux3F6iqBNQ+5jc8m4jk4qUBer7gPuHfwAldnyIn8lReZyM44O4qDQAQ/juenojQC
xBHcxuXUHwlflTZhi7A7MFwD0JMQjwialKlm0FJ4dR44FJyzkHFKEaCbyMDAsi5n+oDY69CSPjVC
z7SeZzJy2i5fhgTkaaRsmtU3pFkzhS1ssgizb8HOam9yIoW4fNilHbkXS2ihRvKfAcOKrv0ab419
rCRaygxeKBG4Snd6JAHH45pPBKGqfmLka/yAZRobMLi0QqL1tfVkJobbRCu1tOAEU7mpck/jdSNq
SbGAW8SSKWbxfwadntovQlv7wQipMlguZN9vBxYMdQL9HJdvF9sBi4075NaxwCc2CffqJnmDX4BS
jOk9FDx11MCFxmery9i9VOulvNysXaT2SUHZOkqOv5C0uJLz6RJJgJ9hXZquHxCvzL/EygvxwxeA
2CW/p0hkpwcLmVe8v2QKj+2UuoY7FfHvB6Wg/QHXMYD+vBPmsVROwaCrp21t2+loiQSk/J7b3Uhn
0h6g3+jzf11RLInXG3fbEmrnfv3DywLWhwKDaALFENu4/7TbKa7Dg9l8snFCUD1Qq8DGz6zorN4M
WWm9gj5ZfSBGM9g0xCk8zalP96KBw6lZWP1VQw++R385OAC+kmANQhhHNHiulRq33hCws/5vihtl
L8oGG53oSL2jAcE4UVUKzYRbtOOGspSvpfAo0PHHDIim3dG16ZoFxlouf6ecRbKJJrTiIz8UsF9e
fsbKw2UmMP4ZBtmfYpOFj5P+nFU/t5320RKbcmhZHYdb99Srgs5Jklr4FL1HHBcRtHlvdr9veVOg
v4xWUHLsshEhxr+HS273dXPodnIYP3k/tBHQb/1XWueVjTIjNmbqVxdGrJUBG/FuueF4872rOUsE
UrU5DDsCskpYYgM0Ixt9YsG45SXKB9G3JOY23NC9FnA1Za4sTlinP3jgVUSCScS5dGrd6NvWHV0J
1sOle8bE4QaQYHEPEszqINj9V3bZYqfNJPYuIaoOpLPCOQ/0x7YQcMb2If5VQkjHPKdb6UDPBsov
f7tpOvzVeUumwDC1Zpg170nCCifqTxjMDv6rX1wpYoNVfXvXmrcfs/7qCwccdbC2jDHMaVWG6sw9
cK3oMckwKqaTHE+VpV3qz6NOpBpIymmiyRIkqNOWmyWsPevxGttQLDQ3kO1PI8RWrRPLMW8Lb7DI
FQfSNOCOFgwBxzbi5+vL7uKJumQknQ841uFOLZ040hBvNOjNcdDXZpsJIoICAbtcKZ96e8LnGdm0
VtmuG0GgNhiQRhzHNno0hWGyTvQ/Ouc7Muh/558+14n+A4H+yYXlURrYOSx7xxR15DgIbGKLU8Nu
5YNwOnd6TL4iuQx2gEcJrGARMgPtR2wnvH1sXquuuAwMxRcg6yyqUzep1dGrKKGWZXP6ABKuFQ1P
/HYKlYjtqO8UYLL5WtrkhX2BcWBb7zl4gw1jTaXqv7L0jbHJkFtMmMV2VBYkeU8MV62OHHOZKJZ7
StRUHqEppgUSCPHFGIXqt7tz6eJSBmooHDdkYe2Y/pd1GDdisOu+Juz3BpL3YI7zOYHy9R0YP0kR
E43WisvP/kbWa0zJcO6ZVWiztpVUQVs6rPgfF1o0d1VKy2GmNQbGyQADAETkgIKlOT4LEjwqBcdU
musAlTab1RoSYain7dOncsRNd9tzU03x/QjUQlB3HDrWeui0pe72vmfJsA+XXZJgiRwuSrtSv7a7
s0wArcBo6xGBC0fp1aCg1X6DkSE/CSnm5fIKU1I7DP9nlyHIwgFj4Rjsd1vjOxLC8nqPWAMC62cu
OYKpkRZ+3rRsL6hSsQxvXOozWvx1Za+Y7E7OvrPNDX7YkFF//cAeTmanPw6bzJdVWf1bJpdbv9A8
S//441IIoYeoqPMfdDZ1MxqslTwZL407DayjtM84mGcJdo7SHTPTkqBE3BSxoFXnjB5WlrT8wq2+
dwyLeXyIKqztlzJ0v1OEScooctx2vv9Ysjs7rYhtYA7BnsqWZpVxAxTs+nyZVAktce69XNFpFVSi
lqFbEyZ2RzFraG8uUlJL2jU4HbQMpoOuPDT3yHJjEvqA1k/vDhmwDseDzOu/nHZaLz4+qYRJhayV
nqhf3nJiZu3R4I1TIil/vOlVPEmldMk6R3+PYRBFt5b/NyY0IbMqLmjanR4TwJnMfLzx9cdoFE24
oOAOHYKIehDTo1f+L0ChZ2dfeMWiLlNKM76+b/Z0D3f9xCi4l9Go4ZDwH2CfD5Z/ZSoZEt7nfsNe
LPMK9KfyzVHFI0XCoYtk0WLEOMIrZGwQbgeh13GQwQ2k5Hewd8tD1szMina8qICBG2YfKJkqdHLd
1X6VOFDfI4T3gPrz6bRiG+vbS/2oFSvA7EwtNYYWiYez4nPnTOJyMe4KCMoi/DfrKWx9KWYA1Tuk
3LBetNCDGX7j/nCaEMHCyhnNkAONIoPMTPNPXh2n85e85TND7EDfiVj2KBHfIKTIaC5FjR598dD0
OH67uHWWSQRmTgdZ976DK0mkpl6qHR1TGA4odMGqy+duS8mX2Djx1Tryc2Pasqkv6Myg2iaDuRh9
DpY+x6qiPYzzIhC5AYF6khsqklP6GA9masuplJu++gWn7nNqCOqeD2ggmSQNjCpXkxDmAMY/LI2z
gNhHVxUXgwR+S4PwdyG2HSL6z5lXgaf8vHllE4gRtAdLVL9K84fOx0jT+dEnWCGTKobqGgL//8Pp
Y+Zh/Vh+aDfhvbCbCw5NFc1efrNQUZ+IT3jsPBdIffaaR7iMV+WNVzUKJV1b7hYtCc59+YCYcDAN
q8zMnJ0F6TQgIZuuxeZ9JJDCAOpldDPO2PjJIVYxLjNyVPBk8NIok3PHGSaEp8tBGTnptFL7dyC1
yH1wZMRQL7EjTCPQFP6i7aXPObJmtoYLfWdHLvN7NZKnkAV9k67H1sb0n0QEze2DykI0hQDQ5rvk
zYV7bIQ8fiwYtV8ABZWsq3dGYnfcJMjXPj1X0Cmhz8y6mYFP71DupbprQA2jobiciyND+VvCqq9b
ELb77t4wq0l0LXjBeIRR0oqT1NLcfGpRdxK7WmUNZLhc0gpw9OPFDPZ4PPswJNw/d7ROAr/rMLZk
bBYmYK3gGYIXdcb5gV1l3Ub08vUahfWfKfwHCpPz2sTMsxnTnQIFor7PY2aL0E8Ot5NqJomBbobo
+DN+GWUzhqCC6nebY7h1064dNT0Y7TDDZXIGpAc1uLWkY8NfvoU1oWPAHqDetpwNMwY6/zRyb/A4
juifhgs2Hhzwm5iQF3+4QEk5nilhSgKvIcODHax7FSS5+IImdWpNSXwE0snMA1fB6ktgjAtjG5b8
dwt532AfZnG4fx3qfufazzqhkzeYPzW7AXxExslhpwr+p1wvKFN0OloBugjjLcQnlUztE9qauyED
z3GOjbBqecpZQZBSeYaxVL4ymEnz2UYPCWYIVdqcDgnbea6BbUEeCysjVcsInw8RIx8CtxkFnVDk
1alwjdpX4+FDOr55H3gajSkEi8w0+eZ7eIdcZRFWiXZ94V3C6cf8epzzOAEq12MIk2/20QbDUV3Q
7gqtBxm/PxJ8gECsfqWSFZ3gfze4yWbfO4DzpN1TKcCXGRo+aJY4qXoPtqybGYtzecgS9OprZ6ev
oLUFP3gvWBpSzcmArQDVd7zStzw8ox7Su2FIB91Z5p4kaycV3Bn96dLIv9kitSghzMPgJRRHd8xm
flaKsfnY8PviS3paiFok9sRE712YBX5DC0kJ08YKShPpkuiuzOM7s8IxYSDEmyS+8g6kM7+lPIhq
ZBh2udYWB/id5EnI4h2mDpoKlcJQV7IkNet+I3mVLTLnjTnp7Z9N2iMkBl/iZoBRqTqOna0tGf96
rtS2lLLn7lWH56EYLIMJKVBesp0reNlseleMAIxjtkag8CWYGqv9rJBTf2t4wLFU8CuvHK6y8vNA
9tJikYjYV37d0tz9ibHqxUzFUcQj6MCvY8pbe8+C5yVf/KUOrSipJvTkXBWXOaIR2VLet6/iY6lq
n23CIxGRU3rVAtiwCC7WD4lpUfqL00BSTfCkAp+9/Bq6P6uBRlmsgBBmKXRQlC7gs+M3KTMZcVU0
dkABRNdXyOCq1/jgPkZsKUCALob+SD4zlqp+J5XueOLHQksgHnicEd4rpuCITtZBX+lbjPK+XSpU
VW4oO8p5Hr1LGWZdHTnU4Ppm/5MA8aAx6Ulgvdk1wN4l+9pJYEckbpQ4knJkYmVrrzm8hn8DO8AB
PowZBw1A21Xqte4aGormLWPPsQsV+UJE7WJ2LjCBmg0yW1V+t0n5840SR4Ec8eFRM4VaaFW8rRTb
mQi/Nh951Ys8RlIFqTAgZgxsAK9ZN9Ce55k64Y8eekQPs8eJY+FNo1D1aFM6yw2HhmgyrFKSDHaa
FTD1gOXg8i1Dj/cLXLndjK2c80brbBWgUKEDnA7D5MsqC2PiimIGvXQe41NLe/cwyluofO2P2sqb
uyKL40bTy07/jsr9QwXb2DCMmkAB/ifKd3hfgItMRiLqy/ez1l08PQ2WL3mZ70Vl5nzAscvDdn3s
vXiGrtAZMg3eTE07CoSG2lQLT45donRLlW0JejZCiAiBbFB1Z1ZqC+qilUDT9R73qP+DL++lcnuU
qoIvRvqQO/8Qt9u9hK+MZAa3i4ZR5lSa/T8wR+NHUu6P01VDQdwKLZ8QF4oKb5YhPhawmw/ARFNA
Sg4EOfCtCKOw8hC9fJQlbjGvYCjo+J5EqgTsofB7Bly+YLMn6/3UYUA3AAg0d1+yZst+xFym0N6h
8qwCnkAoZpc4Y+Q8+owS3CXJnD0Ofb5qpeop+/d23ulELcz4ebqSF7Z/JK3/vKCVFO6/0W/m3WSR
417HZoDW0DHavkqdqeg58QyBTqt5L8cxmygYSs0k4ScxYJfgpv1rGJmBEOZ37NX00JCwyIZv23Tq
+SU1qDVBMGsm02xtrv1+JOwbI4RIpB76AA0gjKdjYI5tug43bpJcnFrriVY6G0bXIesYc/nyoZxG
TXjLSVQQJkHGKkToyC3n/LmLnD9wc9IcrZQTTG3SzDMGXuF6Lu3vw9V6HsCCLqmqiCDVqJXXWX90
MPEA5Xboop5oZvLbEhU03NPXRNrEBpPe9rtl2wjZpv4YAHQiZ3VgONHNroa21dP5yCaNtPHyzqgQ
cOxvleni5zMoxH5DgW2iU2KiRvWiUgxA7tbu11nEkjmkheSd5coiyuCHPrYzXCzLVburDysfZe9f
WtlNuhyyyZWBd0Ou8LZG+QrFaZBco1WlbO72pkUxUi2eiXJVNchPFZNNhSPFPfGJfuRL7L1ma09V
9LlTPOXNBVkO4kazZDVHS5i1PFhhKhfh6GF370XiP2zt8TVAStR3P+JfOn9APfjp18sPXcG0o76Q
gZB8NJt1fAsGuPEokeIcNzcloaSfpJ/whgg/Cxpwk+PWvRhlgy6SCF98r8Nx8qbj/LXe0Pj6m2Ir
kAp8VWvnC4AsbaWAmjghVAZPPBViE8LPvD3hb1lwRimI35n5zPkZu5tB3swaRQV6e+PFsbhNe6w0
fZxWdu9LGtWsK44q4ZTq6mQDMnVouCQ7KmYW3c1qKvkrktJ5nkmBBZMOYVgzmqWOZxYWB7XlEFZ4
GFTjy4ew+iL2yG7yv7HkUiZ8KQRK/PiEz0r6dpqebCqBpsghSyPeODCzQClSIbighqJtn2DJZz4c
AiSj4EYTyQ3XcR/Ran7SR1YiXVh1Pf8f3cU7KjxDrSMJx6RRGF1Ip1T6TQeAt/Yy0lLZ5S2A4LeH
a2W8v6KMAFjotBCIYd4KO9EWcQTU7nm6taMaCaZatBZR4O77O2R5qd1pdfkrN/WfpV6Mjn9GTWF3
g9juIKuQnxC24vcpQ3twOuoo0brmPz6QoVMbVafvqxu/zcPsf0KqM5KBIO5+XMIDW4wVOOQwNLyA
FKZYXjlQiS9DF5DvdEoNdL+R4srNiJqXZf3UwODHL9D69kLrY0bjJwKv3JUlb/qxewV8AgtBiIcK
9Lep3yq+28Qk3+B+UKNiq1kaCgtjIMVoPt5tE/1bNq8XnblmPX9u4NAklGkErtyI4TDHJHZLoMGv
Lfqx5zNzSp3K8535XSyvGOJJh3bPU9Hssf0jsZjTpebABpH6r3DE+V2nIzt8Ix73Pj3VUU6YCzqg
Rq7cFzey9DLgHhN1gsaM8XaxMpNQ2YldUHwgl7D1aTEjkj//K4eC4IZAIRqWMVwP7QaTuBiZRt4M
W8XvHGZn+scMRikR2k6Ia9SVKxKdpnzN+3sv10R1RPjNpPMxnJXgbZ80yVYJDYxJZyJ5fh+WSGV3
jaIRLKyh0cgIeLOJQo6qD0UDudQOLUI/m40cN0oDhWUFWDa/uHSjfdX3lwaHrZjEP+bwmKwZOgNu
nkK11S88yYi0denzNQ4lji1pKin8YOr5E5jUOI0iqh/RV5e4d2w+LmVQQHHWMjpmFteW4s0DpxAq
8rgEpAHb6LLdhfh27D62uoWUR9OW7v5UnN4DSTnVz9K3vR66EbS/OwE95nbYksdtzGuwAkom/HxT
N2XWRGUVJ8aZNoNz0EEUM34xWt7cLkOnUZEQpXZKz0PGaX51zbRb7zo/k1S8/eESsKkmasdwABhA
QpaXMzXjSj7RWaELBL7i3wil2CBWyFfoPOnfP0857q65pJDoSCsilK2VBcb2vf/pXLkUwMcRZm18
eNAaJsjtvjczSMWknKMJP3MghWPvezjVPSAekAiZpujCVK3otHqXC6JePtW9WydQzpna8uoPXzkE
X47+wZ7GANcj12RWClTtHu3UQ958BtkY4hU1DjwH9+Uu29+cRG1cdWP4FBdtjQSg3uaJk23IVIt3
s5g2OefbfxSWpyJ9eah+chfplhRYTWGk3KxmMEArjIU+/B1s6qhtHfg/jm4uaCmKhqWyqWK46j6Q
cjAUh9uQuWCdzuQn/PI5+gIXFy+4qFEiNe8Y1Wg5kAMEpkJQNzQONTvllBjM/rIkNO8VJamPUvts
YyduLDJ15S1i0PEaLY44I0jJioaquZOC7wPfcZvmwfL0BkYBwhcMh9ZlD68URxOxcqQi8aQYWRTK
DQAu4MJ1RI0e8czDmMcAvGD36WwNVJJoPX0el2TkF/nl+dOTIirRrbZzwDc6IXGqE1PnurRsrvW/
S6fY9uiT6TYyEdR+PYIFMdh519qYcHbz9HDH8m+KommYTSg9ObAR1CXaKwy5bIy7pa8VQ9kkMKMe
b7gxSnlqgMUmQ3X1Y4md88i1gm66iPCMu/4xf4HZlGYVIlTSKPAf2sEburD8fcnUZ2S2XdZv5TNh
bVCPyfOHdek9j/eQunDdCKIegZJrnAaoSibka0QZ+n7ua5kX8yTLE+QbqpRGwhbuuLwyMS4fw++p
YpEb36RFaugVgsZR+3R+6OPmsLhfGXqGagegSHs/h8fQIwPR8phAqTTaioUbA26adQzpAzP144fH
4A9p6hymt0ZfNM1wJrIViFwiiSN92e40I3TNcKqIBrjQNUs7LwAGmOhTbakWZJ9BUbdETuyesI16
XBMyDCwX9TkJEBAUQogxjBPSvqXOmOLwg4bcbxRCj2q3oCvwGJAgA4GNmM6IgMsgJ7XsBawhCiw/
/YYAoHzAR5TDpXE6eOiWFXmiQMvBjtVh7kM9k4C3sx9Jqv5Ah98MCciR1GgAK3Io/ztnsA+WIYRM
CGCwntgVJ0WD88aFpmyGXhMrJB5IWNKKPjPgaR0jlNpvLcMqtywFXS6WiUOy19q1jeU2qxvG8ZW3
sAlpF/jiW60rNk2ICbMfj8IIcfu9mpsC6gkn8D8ucoUkxd2Xjj5ffBq8v38csyXpdkSSNkge4xmr
pPaEtxDINeitq6wor0NNp7yynfjVhcdzsjovMDLj2GLN/LA8Mi2dFg2RMJCnRwuQPYpKj6aHxO9U
EnwTGrqA6P2KopFXKxHhfsnpMpPNfdonRgJm5JJNo/veT2SdmLz82W4AXx7MqD42BzEGWZcwRhyp
o/Hl8ghSqtdRfvikKbIzF4LfmOyiP1vjB0g7rOz129YRVmxpgXj5TscHVj6Vw9sQk6hjQ4EXpgYv
0IP9/EOpI++1FE0NXpSZvkS/v0IjlMz+F+Vb6UTjsjXsDb3qwXS4IZF1WA6+nSFjFRqLDZp28wzQ
POt1mA+bwhEEZXawYR8cZjLaZuW9Ur2cxQn3TTs7+wmkGQVPrQQ3WxB8SVe1lcreOOjNJqSdBB5A
sCVM26FHtpWTtS0G9dLrIMtEgSHqwK318SdigCsnaedShQnbq8PuCabBLn5zTBza6SCm9NbhImjT
I+AyYc7m1AkCSLOmiRMJGb77JA9A7CtuZbC59AbJM3b8JlbzUIBfjo+n6TcWWO62xrIr5Ke6mLa4
nnLo81PUYc9OPzG+Xw/8wIoRHolAbYKdpYzIFp9VoWBTEVr5owko+zRuL3wP5f1hKdE9KwigqUur
0EQR+LQiL54qGbBigtl0sTuybzACwSMohsHY6PInb5GwuazGTaDUiKLy66xksvsd8XgJBXiiUO/g
l1GHHiB3DE8+mdf+92kJ7GGcuGcATVnwSkoSMhtOGML7dBrsp1iwLZjKJvzjbS4/Q8kTvGq27h4Z
bMSQWlINjtu5koDM3YITw4xaJLztz3JWkkpq7nYsfXCvQFdOOY6v6VKWWN4mGhlqhzY+tY7YNsZU
pVCQpAgwAPbmg49CPTws0i38R8uZogosXYcRW5qOsc7vFphuZeed/daXN2z3iQNUeJ0TLWJNvCrq
lZITq4ZY3r0aV4DIurp3iq8srGaGhDNh9qTZr7x00sgFJAFmExhJrHj8YEez+Lu4psIwKDfFrmiz
I5ZJVDxvRAkYeVeiDclXIjSjRv40ahkHr2Cow64NZqpACBDp7rjxjyxiDuHv+VxdfpPTwMhc26W1
S6D921AhgbEGevT4aacsUgpyLQiuzSZS8FVOdwyxbkHEa7LYyBuE2pEtgyEp/w5pIh4OWFbxxPnG
OQYif3kxvIZYaISj7QTLLy/FRkxSZyJiiQ1IR8K24WGW7p3YrBqqQ46cx95AlDSjD+GX0iqw1QnW
d5KJjqUIzdRpTOemd/KsK63yL2YOuG05x8a7y9/uzFzJd5g0yd8IJbLDlOTGgcJ+rCG7XA7Cakln
1BKiAkJHQaLdsqK/SpBNQqwh5wkxKEoO3dJ/uawLqMBLSp1nytVgHea023YJ6Jm1IHSZ7MMec5UI
7a0BP95P8mw4Aa/TKRllpNsQhoIxXgeJYESCC4qtozPR4wc1XzEOcMGPLHAjdzqpxRXMfwvx0Ft3
paooAKQqpkrRSZKf0giIExgntzTUKgjWs3vS64XkbY0BArATS3GdCZyQ2MvAX1GQOEsUblQItMEK
F4tMrKtfIXfgKxpCMnn3AHDFGrrzggYsGZVvMYqk0sYapZsa9/ihUZVIRjwfkyR4ZyIW3ZGxT8Vv
NM/v/zaI7FCUqdD2htQtfyaatzJnl6cP3m7TA+02diUDui8uN3hrmarMxCQ4UO9pYUQtgVB19YqB
50TQ2w5hVHV6cz9E+VfPHb6yEmw4cLy27US7IW16hws/9YWboOgZ7/Q/aN2kqxT8I4Dhe5sNTZem
3g6X8oCC0Gn8O0aQoCbF4bkrE+yp+znzIWpb6BKVH0z1VgAL+9sI8Rl0Jjw61VDoWC48awiXwbzO
ANAdGYDCSzWu+p/9MStYMkz3FkH1IbzXDFAcRLgFmrLF1//mzOYBJtrXIIHF8po7zIBvjNFYgYQ4
cTga4a/MxxH7942xijCqaYC3x/rzxL6e22ihO8ei4Re1vH2PEGMDzYpAfAfNwwLP0vrjGvZ5RKXi
RoHRDlNTsWG0u2dqhEJO30ZjE5PRxR9cVYgAUfYNMmk15Qv191yOZDTMMoZ/2JQCA/diaWw6e25g
8QVGuujxbmVd9JvV1E3WL8nGblmSStNotvKIMYmxMvo/MI4J1a+hQCP/p0H9blH/1MTe1kcO33Pm
z6N6qXASKQDfXLqA5sTBmCx+FKkZJDZCPbc3JC6RN9hghoixOSZGcW86LuEglTB+AEFdECC3tPZU
GWsi5WSHeXvl7MgfPrtjYFqediIzQQYHWXoS0ZreKA7m+X3kFvOKHhox1bV0c7+ExcC3oydEO6fw
TM1ui6AtXxsTTgh1u9lu1F0cb4NZkZGAHFTQmN/XtNZ1yQnPEAJ3VghdnXALQQ6UweClFgKR14E0
IsFqtpcdA74RWvF04L33I8gcW8sGKlRBPFJrddHIbIK28CdzDlUEKroV1q5TyJkWAVLJimQiD1qF
P1TfUKX8ckI3TSKDgbD0V+mLG1z5xCKhA6hE5VmcFY8F7gCUkyq7UYcaXh6rQaokmiq5YnHwwORt
dFwa9yd5abrv84iVVUjc/kx6MW9ZqdwzW4LrthesqlLgY6HsIwcqWr9w21GBimMEtevBvpgbVKTh
mKJZTMn8Cj4C+0Tq2s5+H7oRz5CpMgLZ6x0p5f2eSwA/4ejlOnxpyBIoEMkGnvpe6FZ5al8rnis0
ar2Xta4S+UaPxYyuOLPRE46DEpTfkK6HChOOf0wDEunvQhjJSDIKBRQlhbsHwnLuiPMZf6meEDt0
kgOws03NNTiUhU3AYntltb1jSxL/F9OxF4PQSkEKcfhwNZKC83lbfThs2V3AvoBnfvKnhV7o5lvG
yp7mnoPqJSGw4MM3zGaejq2ZoNLIAaCjW2wTTNgPNJtdyUeVF9bIAThtwfSS2hAA8FQSi1OfDdaa
YMG7MyPX+hS6i4WcVU+17fYeExkg9MMWDF4/80oqIpw97y2JPUSAflLEFQUyzH4tszXmeQMly7m6
H/CiCoVQ/Ybd+GiLRH6Kqjjn38vEsVCxKohug6Ub/WnJ/mpo1EAPV6j6seleNTpaSAKP9jFx2fSM
2OqxGxnbrruWn88KzJRoe89SFowIswyMOrQ+Tg6TwkbXwxKiiJGEZalWH2+yayXUhxEdg1U3GYPX
XU28uIUEzIGHcQak2tiJP6RzdS/IG1lesKYm6UWTiGAgDDl+wz0/OePJH81cPtq/2thhqgI+THdG
IF2u1BKrseK/jOAl0AcuP0uPXlehdhZPSySct/D5FmwtuNA64VrHvTalTw3+lUNJu30FbOOTUNLf
dAYmSrSttN3gogAqv6zrLZe9hZD8JzAko5ofnODlV+DGpDIDVd74ID3nMfwwRyOk3EJT7/koPtjJ
n1o1Jq/rlV/FW9CmOB1MSkF0p+hxIKZrQYMIQqmZjIy3wMsh1CIv77DG8ilXGfKe3udtEUGM+pvr
T2nAojlnjrZhAJMn+FIiAKhScYZDiwNdnbXDKO9evo5KNdgagCw8rNdd1bp51eoj7nAjU/EmYwy5
OiG4XeSpmDIhxM2l2N1nWpAfFiR1WHipZxOeZ6AdP+gh0XXLPGY6Jho7odfrR46i6QajVS+XApkT
lkpGTtANhkqnDxb3FjBWFXn2HgskQJjceSOuKFj5IXAmmFN5yA9CBUDjZJ0CEkTDwS3HNisJSQFX
apSXRCFApus4NzR4viUcg7TLlSD2Xiq75n+VLXb4uXNA/gNcIsT7A2+nSBOI7/atsDKQSepsa5N9
ENcmD/7Rw78TEWVDTVjlTMh7HO4+D0Qy3PIVUWW1zwCb2duAZ043pnuDOOCAK2vg7TLLOTW4/HZd
F+hDPzTIH818K+twF5FSbrFsbHm75aAyevGzuI6/2lyMz7EZYa5uUr25vdmkmCkJF7oGRgfvTMTe
F55OxzDLXKDLiQ1j5wrhA1x376n7xQwVbnsz5RdEDoeyLYzYAkz7WmzuuSp5cUbkviLZJ4k8OLhN
1xGDQ95sxN6AF2+pwpUNDyTThM/mfQ2amcHROmtp4p6nqJ9pnGQemR1hsfEzCLS1gkd7lQtOQ9qQ
WY1OiWk/qjXaCwwftZeSk+R6REyGOwJyxzYR3opGaphYVc/tGFTlykCn3I1juFu1xdni73vVD34D
5yq1OFbcLMU8bgRmZRt+J5I+uwhJpVnzq0e8eGsEdmht7a6HXOAcVtHGNWPCL9tKIvYSC3zRc0JE
00fg1t1q3kvS/LlK6d2pa5GTHK4PytpPqf8COVN+bBg75ylLVhtz5mT8xUyjM3WwIyGsDRHIzypa
pQlLNxaeSV2Pc3Xjrfz9UfwWT4KMrj5J1Catd7ZekB2VqiP9PZtjm7V3iSlZTpsWTHusx/P2xsul
hT+iZfbYt9qj3oc+XEte7eZgnnmSqrm7YOcgB0ScoxpaPawU05GBZ0UfUkI3TOenc0PGu/bGXsQh
l9IiLY9TZlgGSRcMadN+URuQnl2KdpnC6dFpwvxRCReaPz7DdHBIm2i30HoCsEhdREXiTiMD5++Z
quqPyeJa8vdCtig60p0OzVdfNwLAwYpULuFSIIlmaFgT9BYnS+uAla4lFb0nvQFTqFK7bMnikc6X
W+f2IMpx42FtA6Njz2KjvyHcOOgLYuJRiRvpx91KRVXi6BmsDlcamDcxIL+6OAuxWeYP6KGz5kho
58dRbPYATwTDybpgmtStUbgypA/fLCAfHuys7amTBisaisaXTkLmR6I+1mFFRmScl/Jdx7495e/s
Gy/twpzDyLhDu2qKER2AF+6PWA6Z+CswIliMtXwxkGs+pxxl2GPvnS3s/+VwraoqHvnM8exj5/mn
AZDQEzoWYJOK5/Ay1yxQyuUwS8ZGHhWkB1RAifeJJwmkRCzhR8KR90/dh6R4WuMOApjaF2PjSxR+
AQWQ6X53eN+MaEOD7+ExvrTsL/GbPexVtde0CQ/jFz5cyS7l8D8Dbn41vBRwNAymniYtaaRrdG24
9mZBSk24a9gyjGUQXU2DsXJpKboaMbHTFItTdThunjOXGWC3mwH6/DYYTYxMlzZHyetJIhHxQ5GF
WSghT5G7JSe4EnoaYCfQgtGSwBhSzm5ZeIuaN4QLBMv2vsPSK/Hplt0HZPVW0B0oIfy/nJo1Xkjj
UHM/PzlBkeRo2uGDjL0/u4lze/Dhnzs4RdoLoOcrJ9ocqLfHt2uJTTQNKd8moeACB0OU5KFoJSot
sxSjyvv6j/8nv6bqy3P/Hdnb8HFnaxjochR4PUwTQdXK+YNxuTwFByby6NlnWcL+dzZH39g+Pu6W
2Ih1y/ikgettx8WWJgE0UL8G84rUJ1Yf12EZrLz3tLOU2xQpyiKK4VSjhXayEl2CT25EjhLizMN6
lCfvgJmylMrQkPkfjX6P7pqbBVf+IWW9v2vTzPHj/cQx6SFhKpxtlNjWMpkTRi8CX0aCpscONd6I
c2yoyfCk465xWv9K90eT3fsHhHQqwLwfY7bI/I+wzLzdIzp3oeUkYo074Yg3Zqy9OnimJitghd9u
5D5QIrxbr7NdlqllzV3XPIUm4Dd96hgRie0EGJ3tmDeaaW5Mf+AzdgpKtWiQfS6XKoRBUcW/6vPh
CCs7iZIQTE6SS0CtXFpBvDC9cLPzKhFwRUJ8gA1D0ZN5Z+ja0V19dq2ZUVgD2yPT4Q+JIIQesjNo
R7nQaGaa9yc9a14F5Pj+CwczJEofTfTkO0q0V5dewnJQ6Qwq1pNihOXeTvjKbCLyznfu3i/6AD95
fyw4pgkIRtuyDETnX8odqsKI2GVvZpRY4520eUoCGwJUVZ/LU5fErSjgtAUfXgouUAC/+MOTnsMH
JLAKnQfD6+hzGpU7laiDbuOBhqQ+hcupqiGHcDfbPHeCtVOWJhw1oIwJyADFUPWuZynrBWTuhQCS
MDmpBTsxq6bLDbQqKp0yzwXDIOZoAZCFPhZdzHrbq2abdJoALEXXsRQV3baM2ZPgm6mlB3gRommT
GffFpzMcU5epTP7wRDfcEc/yj1T1lACxaZvOeiae9LHaT749jHMdYSiKcJ9ksoF3h8TrmfUnlBQF
Q4CgevAG/ekwSuLQd0ND0okzkvEvUEVqX6k71YI0iP202ILkr6xS29GIndvCaD8SyiBUwF/uaHbd
MH1m62h21+59tZgMC0lNVJEIjuVvhvWJmK2pkBNSIxoyU4M4DaFraRxeF8o/GHmF5hlBneOUifVf
0cwC1ybWFp98cu4TKiHc2T/o79Kz9Z+fOjVquAPwN88oPnVa1OeEvEMqrWoK5izZmDyK+55WWzgG
u3fH32hLXBT/14B2s7va+QcP+8kY+BYTV7cVz4+t2GNV0lXGY4t1qo1k9ZLG438YbTMrVI4bt6UE
1i4iY+HCcwxPgrZvie7HKCIEqZWgGqQASSV5tePLrFDzT9AKvcgDd0BRKJ61eGaRoUd8jcM4Y8Z5
JpxhHpfSPs3SwjlUnFsg2+djGOv534W9FU70DWuLHd/6hqUYB+o2QVfL6wEUpcLT/AWqjvSzTyzE
iYGZVz3NI4SOA5sR6ii1nXtmkFafLO3NGC/UmaLNKNhSAwZ5PhOTyTsvw3u9693xPpRzB6tbcGtB
cqF6ZVg4nGFnsex2BuqUsNGEQPaEm8Dy4/86ormHeoqeKIHLKs6K45GQzMcBUASVVRNr1qKreGec
qVxO4n6LS1sCoLM4UPky66iHTKXSPV3XflE+DJHtqUmC0oKXu41v2wF8Q1rSqOf6lkeKNuPUPld3
ZsD4Pg5owD7uZMyQhBKYJ6emaPFuG1IyOX0zLqL/vH0pcjoCWs0zzW7LoJn/hzjiurVjiwin7DXT
7ZZCzyGt9ERqy64VIR1dSmAz57bPrBFTdqruW8vZqiNl2GAVGz8lsoSFIBJEjTpGBUCn9m56u/xN
40MDyLd3BAZcl/Dtdh9V27z1TqOBqUYuHaw8BkLCBDKe420jawa1mwpusn4yJrDoCcsBeBnOuoJF
vTB0bmy7cvZlnilFg125kUFmeYDNzAZeTVihH4S8kBd2xjIklLpzU0sgGaWQF+yiWruWthiw8a/3
I6cjFAS/vA3GIhcsEFyQ4N4ZJalHFqcYv+7HuOtEfEtiwYOlw5khpe+fT+2rmp/Qd32Y/oY2hSDO
nBYtTbazAN6GlpzTPjh9skXpxuERO9yJb/Onz7IH+Cc2YogrIfKo7gm9cAUKvPmjgVn8CMXe4VTw
jfVbFqYIB9vw62WPEkgQQCIuuY+yYSgQSG7LzwfEvhw4WeMk1sLXX+zo7kESH3YTzxrI7UF5Fxun
PcoC+1Pt36KU14TI6P6Fmb6VQCaoWoE1xqJiGh5HgXILG9de8rQutgLrfuo3a4lhsCLjh6n+VBLK
6K/td/GdnsJ5XtCwvWKDpmMjN70CG3LsVqKCUmr6aBXZp8R/89yTeZ+0xgdHauj8MRhPXJ6YfV/a
AA+HOAm8UFhTxU6ww1lfLpslV5MV2DPpB9CVXhmmMgfzYHvTsYPzB0rqpQMe+oad5XGPDtLbddUq
A5eTChOPAoZxToJooOM84PVQMjr0bjzaoIrYno3hniMx/c7RY+CbLQ2jqxIbI4WpTibIyDtBJAkC
zKa5gyCQcL9Rw2Mup6G1vmta0+oBZbsS6HvKWQPBYuLG32SAQf444gO4a76fpO2jHwj4P+AOeQ0a
vlG7AYW/tG0TmUQM2BzX3EgiXyNFYA2yApXFoSwqt5bMx/xQBGTr6qS1jVhbUKvO3NUcLzeGhdv1
L1Fmm8STpWjPuZasbiEkPO49sg3xYGMcspnsma7mBgC8koBGyaZppb5TTEWHJAFKHMqz3nTi6GVs
jL6ulM7dsF7ASKAiqNuQ221sMAqMQ2mS10vd5EDRJN/NyG9DVJIaX7Is+81VihOTPyi9+qtxfvOA
Q+DXdUp8CiyhnqpOxnkpDAs2EzV2RBjDDpeeMlMS4lrBvO2EuD6gmFY+sbn4zFoVYC4OKu/8T31I
I5uBPQ30SKf/RnZWvoeEn5aFmEdGg3dvhWxna7RoIuGyWpjZOsJJEgNujxomuMAP5RxRKQM3NmR6
Yo/IXgdnpjVa5GO7z6KO7paTvAhZs9/fJhlrE7f23KSb0V3DRzcrbb9m+T7zh5t3iMJeRKpeWx4b
tE0DhhVcdjeSi0jk1tJwRYy20AJTVn66E3RDuLgZBXlboA+BkyKPaxJUX1s8AoiUxltPXwzv1VMf
/XlOu4semmqdCKqMVmU4JbSNS6GAmlcZvjrLQUeaCpQ/s3Jn/u0qzxb2npZRJJH4pLU8O0bHU6f+
gxZIDNn6MAtq+DMflG68KUp4u8C9V2/KF7gAXVX+tM3QRhudeWRni2bibuqy+Yy/su4bd0DawXUE
vPo+2oslsbhtinc5Ic4vEt0d9wTMOMfYLVELGwfqKc9+pTc/sfArsTkGnLbsnf4V6gvkCunlLiWE
OqJUiK/fnSD+DmRnD8hKH5I8HaZN00Cx3AoNyjAtZIQHUS+7Lov2wSoRP/PdQqizG8Uc9f1gJDw/
tF4dRvRzqMqk5opA1JOFAnBA3LJ7KbKGzw4/MKMYoYCUy9cKBOX3ZLDj2OfLnjngXgNpyOiQ6Wm8
/SSrRyeni8DqE7m4fMnK2gpWNAlVF4JgquuEeI7jpaEg2I7UlErXPrKkrxjmOCf6+BAqElcXv9Qc
KumZDj9crEZ13TdGHNEVEYlFIaay1Qm6D2Uqn10VLxXDsrRKT/NRCtAQfhE4VnIqIdSA/bhrp/c0
J58lmpY+XEk5Trqwu1aQKoZQ6PfG2sR8QUyRpzdh/Vn50dzvKpfR01qtuT2ou29MBhrsFkjaWzd8
/rr6s7LrsoRZS1MP8FQhwtMsAx65ybNTfhrSrEqY5vbfP+nzeaMlSjMtpZnpSBDw24ZIx/tehWRh
RHo/WExkZSAAftBPXQDyr47RMxR76lwYzJp3RQ5MN/Cz0D9ugQAAk1Wzz8mTzvPuMLk8p36tbJAX
F20+KQuGZI0/0oe+2WVfWEXGPCU1gQjizjOKpF2qA5VY6NIsbwVCV6nm0k4W4aP01QYqvrPSvL2D
rrhIxO5604NIJbZaaI54eUe0CV1YmDhy8wKyJg3vAfX5f2huu5KoQouj3Bod0sgnnjmYIGCXRBwm
0YnTDUobBmE+34HJrSB+1sWV4kKuPWrFaw70TYOFnNZr2l2YX0OgU2HX/zVYzIm1VLBFoNdALoHa
p/7hoSgixzm7zGKMVS//RPMC0LFGC3tBm5Q7Ps7XeCRKCbEU1p88j+klq4/ydSVmltUcAL7jK7aA
Vqe33PWO+QY/niKnSzVKswA+sCfdKXdLl4iTHde/SQ0V6EW/+91FqzBXNnqJYlIOJuXBU3QZidE1
lU/oFKQu7pyhykuJz7vwUxJh+uB7ZqXFP6KSS6tHxJTzKN/HkSYxhpJ7PeVLq2jiMoqveH5izJEm
xFzVcXZd5ztPG0L8YYkMzTqMbMbicwvb+bG/dm9RBfumVHKZM8xBb/XixbgfyAg74b4HfiMBnDSn
pcmcL6bQrMeFRtmahri2AcFh2IsObgeJktIY+KjpOq2H7FONRpjRjwoz5ahrWLsfaD+WR5qU1X/z
HkN7p7Gd4szAJuUrHhppaV5AZc5qUaQS27DYYey7Pp2ObRtSntHB1qhC8nfFokdaqJM4C8P1ck9u
wiIFdKGw9rEWR2En+X9g+zQgK4+DTB4ig7+5ktkzoUpwuoNNKd3IJLQ/DtW8M0b8yyNvQeijAE8w
3BtDYXGmQo5u8k+j3HzigPcjarDfmJZqj8Ago16KgO3kjrrqnZut1JsYZMG0v1oIVvy4wwf+K+EN
anbE2Bkm5AACgXwoxv9/2rDsv0x0S1/S1FcMbVY6jpdFUKuped2KwC/ShwZunBmpU8bYw/qLVd9T
6uQOHTmGY8gzOCNvkshBkCRJi9b/NPp55e+EQdbJeOlnlC/GjYx0fj5IOKNFGzE2JNiwdyOPKogg
DDFOOw/70GBSllYzP5e3wQ1mXYY9UwHg1f1uBZ6mKgR+6uRSuQ4ru6n/5kF8nFaSXD5Ellr0YS9Q
9zlJt8KwJtoChIfCI4Pcqs1vmnq0+mglResSk1k7Fcp8vCv5J38nhfyrh0blJpgS8VeJBviqzFAh
pLVKBCLkozy/WKIqOK1T3SYLsClIfJV34/o9hdXlbKFasd3lZU+FgNatyvPLWzFdUYsqgMkHcpJp
9L6rQ1VQev0AC+v5uW/MejCikjgbYAz9BSvtMJiTvrEuHolcXZs1h0O8bvHfStK0AGQI035z+4nd
aEmGLHeX4g6hI0F2m+GOcaZlyINPohTxILaTQ2XZzQW0mH5p4pLqC/HLT8CDi4kT6wsbeCJubQva
WdNvdkLZMOgiXO5J22MlI6ct7dvII42E8zrYZFpd2U1HsUsNP3CSsEcPh/43jsVXPJOhx9OULkS5
mkUG1Sd2St/YBDVnc7e7mNwUznelM0+xQz72RQMqak+Cl5GSYZs65TCbzLfVYWAagQEqacSp2uoB
ixl1EClu651flUoYDZfGlHvHdkm1Tsbt0rHY1aj3+ytapwY+UFXcUaZy+tiTrBic5AT4fMeyVVox
5rdEKlS4Aiqijtfeh1lPnM6bnlbmZXcSrntyt+SHA5ETz+yjxdo7loRfZApeq5g3buobGbTCxHg3
Sd5zSY6u3FVN7NoM31JQKOWFuNt74PUS31CYvqc5kLzQuAN85e9FHz0dfTQAOZWAYpzd5NyRtJof
bBzFJTWAxBR8biNkO9T1yi7vEb4A2LsG32dQd7KcgVt9P6J9C9/qaxP3f6cjYi2OZJoFgdTi78e4
1znn1DIVbUYzzwEDEc4QkCPcT/ihehB4pfP3vJoEHkXcxOko5cFAtLzB2OTnMw8LX8Nu1wvKFw99
n6qsgRhGfs3gmZYsDaLhgqMQL7iLSGoa5+N17FWbAiNr2UOZdZ92JM7/3iui706vZ4D1xIkgoUiy
C3MFPuOhScSMVU1ZF3LT6sKcrSG2OFOKK34Kc7dY3BqprwsoApim3X4ijPD93t0zAdyqHmTjncvm
CZpS+LFsQuM+q3hWNGr4xoO00N8rS1iU3rqgFsy2Brk72UDzawg9qSf4vquRjmbvN0gMjEa0Et5C
Wi2alJtjN4sRdM3JDM/0+b/7RzvOM0nWxu/DglVpOcvbz0qy/JlL/WdlhUAu+g2hF5OjzgUhUPzm
mUEQjUPGri6v/9qHITwRrc00f36DAd3d861TZFSCw9UvPxFPLxY5RygWgdGFLYpkqLBywKIYZaR6
em3wLP3GMj9gtbSZFRoijIGZI5dCj54Gxt2VK8C2XMU8h610/YiemQk+IAi35QlgTzA9YYUgXH/X
s57v7GQEap5S03i984v+WwsX03uzqer3Rf2CgmL61uCWi8ms+16cmDGVHuM6MbBsTQ/OHX8L33wd
5G8R8p+JsFe8etXzN5ug5ndfFGt7ThM4CMy2i5S2BNr/0JwRXQTArgSMoI0jwrA9TO+KAYJ5tpCr
qGYE8rff9zXk0pzK+TKsBGTbEX4RdkfJVxP1kS5AfK+11iQ619fD1+71h59zUjI0uvOoUycih4pf
2VrDEjKOMusmJN8ymavS7cYf1lUDMTwXysPo25hrqvVOwYmowX2nK32YySe6vOe2AIilotjgnf0l
oiWElFVOz5rYSb5QFP8534j25PQZTkPDIAlnmTvuBr0raTa84UgzMxbiL3U/xYbRFPs6+LfCeA3S
elNkiRSvpdBIXZQ4145w0sPWR7YjrmBc2HAGFl1VHDo4c25nmJMzUiklaO9AS0tl2KUgm9wUpgUn
aYAE6F9HvQjltsknlNycvszEv2uyoWq9gPvf0fhInXxiKGR09ZvcpmKMTbl7GHeg+InnT0XROtLw
nachz1bqKG8jUGnJ0blI6i4YpqKPWKcJGN362FeBDCdB3TmRNCFpQexi4/r0/PN+QwwIwAxAjkZ+
B8D6UIHOiDtOno+jmyCNHm6jAG/Rc4gcMNsGOU7vYX4uZekWB6RSJ4JXodUG1VdaTX6ZDNAhZtM1
5hgPGfBYsjf87bigMB1bcqDHbkxqsiFkJWYO6owBmgOkP91eZ2lCK9Q3THXc6tOdUhjaqIp2fSBF
v2bp4I2f+HhK/XZu2U51ow1uuqbCqOpybEBp2W2ECK85HV+8sE2hBFRnMKvxwfI05UlkVvZ4OlLm
bvxtOW+sxa3ugFUSNJYqFjb7a7Hn8iEFh50b9RS/08NnNKe6VQ/Ka2cUoRzVM/KtePEwbvPGOAmX
nzAk4iGCuWr0SjZbsL7S5HAuptobcNXKXQvEe+9aJMFWZlXoXZUITMX1RYvMAfAdchd4eIA2Gct3
GfMlJsu1yQRgSKgFeV1/Wp7DqL46oHKIbCtyWD/r4aVpqwCqGXQ0GPjI9UIzj2MFLTOkbpZzP1i9
YeoFAhqVBBuV+TfEhpoMyCIljFCbN1igafKThs+mbWsEPmw55feKc5YuW1scq/AOTvzM4SB0bXy7
djDtKzQeSq/yk1vOcAcl79up37ukOQpFYFMPXH0SQ/a/sdU7nhMh7aEhcde4wFPGKg+PdiOuZWhH
ZM1kF75hpmrHtAzjTWpyQJQeiIHE5cvjKikBY8CFmUK2uG3VK67drcqaluL+UtEZnZnTP8TsymJN
BVKJRHnO1bO44PWQ5rfhN3MbiB2p/C5LiKbp89R5ViONktrvh0kvbL3LX2jx1ZpPcw6tr9Ss2GKX
YcUK5g58Emb6YE06uGuqo19CzQKYiiaAW9aw+5GQJvfgzsshKWGjexR/49X5/Q1Lh3scfhY9k1cZ
dJZHA/Jg6XU0fggJTS113a3R+3bQ6vMqZPpa5Rc957NYBu0fkB07MeBbe3/Ar+MpDcalMLxhvOPw
8pBVbz99H/ov3YDKS0KaePsxs0JrvCW9dboNpLV+UQDdbECDwOp6o/PDYjQ3dOdk6JpNiq4W7P4l
gyKVNGsASnf/hazikXjrdelqEcUThvVFNO2WslULcyFHnwJz8Fef7L/97txwyc4h0VuSZDAlzy5g
y8/MrE6OdDFJmlsEFwzJzAEc3vAen/2K/nXIm0lcSDq+KnPPxKMw4WYj39BHDS8pv9OED+wL/N/j
DBjekgStXGAV2ErHf2plmCd5mrlOrfAPEl47MAD9CurljEaSRagArVU1ImWln5nfgvPNsTZg8FvP
UB1wfg/2oFv44t3VQZIWOio1YANen8+9Sc5O3AtMz1WVNPkdep7zs7heRucpslJIoEQhvGvt6ieK
g56dcb6htIfZEAJo7p/VDdxi9lJ0V5hEeOq/UzzkBx+ZZlgqbNtdkblTJtPHVQR1JF8lpjQaD/Xx
LPxdrSlrczsAVOr/QkwOHEBq5qvNjcN0hGGq2EKaluJDCYEUamYVBoFXX4qXrzafL9pldGRdgO4U
AYJ0hqBfwVq59M89vP3mdxX302mCZ8WAKQQa7cVDYAjXkwuaVQ1AY4TKMKxEZJpMVCxYUWQaJtiR
wsewfA6wFblEXhPln6viaJRKldx1ejSYrzlg7lmC30QJaSfFTOpe2DFs/ddedYFfGs5/osuyjnSG
g/ADA7qhZiv11OOdam4OE7gAx6SPepTno0c9We+tcy3nfu9cfppxUHj/XqH1L1Ttuf8h16sAhhxe
7tVKkHVg09E2x0TXuhTwcvo0UF0YWMkfSvtLhfD3zv7WMMu1S8ZFyB99HJmZpbQLhAvWorswpAf9
ma8OAWJ6LqtHuvMMJfkRLIP/UHHpiS68DHlOiiwGY48kNHUtzo6scWHMPF2rkffkbCMwfRlwxAjY
nU0KIrpXiIu4wWAedYZxTNMumU+r3Xm3JSwvPzO5LBTS/44F7ILFP5vzeWI+e4jKd9tjftuu07qK
tWcg11KqfGX9i8Zz3T8WsOkNOl7PssvelkVzemvZcsHVa2lE3y+YtjvZmF1tyItxGqx/cdFG7h6Y
TghqI2GfOTcToouF46kO4c2RF/HwLuFo/w6fV6cg0ah02U5tnrUpqPBJwTu4vyArNcVFKHJ97Hs7
5PSGkeFzJxV2YK3Dfh+xuaww/dmKQYDozdlLtb4FcxewVTvGjo6obMWg6lXpgvJrGBetHB0L/L8U
m5Pbz1CfSYlwIUIPfNvzRtEqqgqwG2nxqGn0pQElMcxWXWfIdk3u5KVJLBSTGZ3l0PIGQS22IsrO
Exv13Fz1tmkUnbmAifrNmhy1fRbkdylOSYhWzsHkrMqSBcM1gOkwt614zBmGQhO0c8rcRCWSE+r1
TNl0mQpeEtetZe4JUjL/XzG6N+8P4JrxapohK7K06TEnYu0xVppemCDpAZMdrAXVo5u7X8+1c8iB
t0iF2QCW3g0Wn4SaV40eLVmkUcS1ex0mW1L1OF9NuVRpDODgTuGBILi3VYOXTAhgRkP0Gxcf1AP3
S5m5RaMg2f/DrpOwdukqouWxz1A8MZOhcpKoiX/DwlH19PiRPJ92ebbbey0kEB+ca4o8FrhRcIZf
jnbeAeEoNyVo26ejBHSeIuj0sak/kWmUBHqVEzBBzBQg2aZSuVU3Cs5YrAbX7dxr3V+3Kg31DhGU
cWfUWAwti5i//JPk+erMf53zZPizfRa7PdUZ7/+Mi2RgqNljvY/k3zDxt/IhnGrBuIbfFjMhZ8Eq
BXWH4C86KlDLvgXbCwmy+RDoHoRWegBWV60VgaMezkKKa8jIzQ/y7V9k7OcE0/ocVQCFDaMyNeUG
IzcJ4R6FCQutI66FCle2Sf+OfkAHK56Y3mBCD08Je7mPrhHHf0qn4vU5IkIUZjKlO/HxrSCfYbdy
nke9kSxUh2ks4uej+NMmjEA0i03oY9bbdMbE5F2akVgZDNv1ESSWFnI1A8YYyJ+L07us71xd96Hg
lsdICNDEJ70W1hF4AVWD7VnTeNGtG/TesYiblL15Aac24AGv9WuU6dR61WdOr5ICghpYR+n7vtJ6
GIlRpIYToRh8V+VTx2jWm/CWfedyhlS8MrXXfecaDJndHIvgqT8F9q26ooSsygbJEOqdIOxEK1I8
qzaGxPFdUvbzwSbi0bKXTGMy1MSu8Uw0ycWumPc7JGDdkK8JmlmajP3r4W9DY4K/+a4jfMJ87n82
6Q9rcq5gUfAauczrQvAyU3EcadGbQWI+Aq7qoy/qDO7L79tVDDcEQYjKZ0kDozfzXKGqmStuWT9M
dsOhLGana9nEPlUUSaj89CJri6anrrzVPf01GNop2L1ruRupK3jpJJvTKmMqgXuC87ZVsarXoegn
bAZa0lifwsLa3zgEnbBMkgbFyY6fMtfiXDWqnRbOW7JbDIT3fOIoHXBNEC13hU0/Wc2tthaBHLxA
SiSqLbZQv2xLx960MzxPRBf8fxLXfDVJrFNGP2CmiKt8lngF4Jw8/+bn5TL7sFXBvLo/NIxBUkT8
TKpmDfwXFRCVb3ZJKwQOHqCSTCh/9G26aYk/gTj6fSViFLdAqbpEBJgpsGA8dqOWXMg5C5MLTIeq
IZaQFlG2+fSgGtV4PZwYkGdvHdsTQiaCiZqRF9FdF+SQsBywK2ggQZRHlYXILH9mxj8b6TFHJemk
nBdOnSf7ywpOZNSXQJcJEdMrSqXiduSQkLe1Sj0TT0BAgpXYZyrQRP7FxGCAV3HWEGDO6Vl8nvCB
kVcGYbQSRN/qEvStRd5BfZw7XhgKtyUuWyEuqsShIcf3zWBl0ewvdUi9cfOK1Aoj4m2mAxMOtw8u
S/gHrlF9p4grXgk4TqX4qUAdaI4AE5W1CcQJAEQme81nX3ECfX1mTH6ODM6X9kftsMpzTAsgVIga
BaomDGB2sjnrhv/cckMFsYnw51bpg/gFBc8reRUMTOXAKF2RLcb6J0e7XCvNEx3C5qJGU1h37O6+
4M6tJs0GRntYzxgYQWMxJ320KZ3eXjbxZC2OqSbLUaYX5WvB8uVAUaFFlY2NV+PQjPIlapJfSP5/
FTXVDsUKaNO5Aygh+PPJ2LUOnTD0Tij9FnnEZavFWkcx1iHleLJJQHd2uEDxrRWTcR4DHPbRDBSj
dyyh1sBvtD2wiIUZa5nbiBUCpUajkSOKi/UsP4FVR3YH210/RLkQlRt9WZ8HQ57u1ZvBjuJANY6Q
OIcBBhHa1X+m2qE21jfboRHij4z1NUHqyxdvCK8njPZNpqQwP715emvLJ/uavO9hDaMiKDfwIglN
Wx4ePH62GmHB4K6Li8PFDwlltIkQCkFieoEUSmqdHWYKCvo2fOPpga3nlM8GnBzj+D7sOwKifxTX
2th55ru6jy7eV50U0a/w8/2Sd8WA+B+NRf/WXAMReQYf5knt2NLk5PsVrDJH18S+oYKkO/QVNK1k
mKJeoAXFmgZoyFLBMBjQQzYjtUkpBmdFIYduHLE1UmVEwW4Qz7gVM3P50X7HGlmDJAA/9qabe9ZZ
IYdCw+gdN04w3hIoSmWQrTFTF71rrI2UNw0r8WQwEaZWn1TYR/zZa3zGDMf+oi0w/8RDzuN2MiiF
gX3aE3hnvvOsuq9vIzkAGwxIDuUk2MAY87tek5W88+yphdbma+RmWy3TYNw9vPNqfooMwRmxlg/C
E7A9K00e5iQiPbbkpSFT0Mmej4OSv9KU59MptvXd/ZBwjgPa9lEBd5bBmMzL15nfMBJUWxNAfagw
ae1cIP2N08pjTJo2o6KDtLEhXb0ywzEZCn6Imhr2bPaLN6sWITTVckKTpKeRPEJiiv3u4OGi22GB
6hxlgSjYlEgDDk+G78lnE3qJMIGY2jheoHPADwglssTBVWj5bLjew1Vd8eNqZUT5ntdKHMmCWgDo
1qjqBn1eGFcGxkmgEiy4OkN7fO799ffvj9sa+zz6IkBWk+yt8y4nkWy6rzNN2XHAG0QmDvkt5DOD
1G7DAV/J57JcNBnbML9GlyWKHEKD1QrqKb1Pcxh4nmETJ7YpgIcBY+upudxXzYnMeimsa6rC1UWP
z26ViO3SEJb51QaBdOo6bXk1HkMpZxusSAX07Y1bLB2epaBcpHpYhKAjKn2J+9xz+/gZa0ywL8tF
GZ1Dv5f2XnR766YpPBcVshkN8zsFhCx9uaHQ+Q+ZcQATsk83+3IRDiIqTnXbOVBiW34IVNWB4Zt+
8V/ZWkpsLnx08lQux7TAuwwCqei4tmLlm8Bb4V7ZVd7AWK/s7y8/ZHFjU3XR+evdrDG9nGv5vy07
fje7RCwDjOqfbcuwq9h1tSG/oF2MNaY0uwfBln0zaquYixu18Id8TmJ5RlEzPXJzQf/+kC5EE/yA
I5Cli7JZGhMQMQUJ0iehxGAg690u1WYDAOTCdCR10/66hEcZso2RCEexhZElZ0TWRaEUrmDY1FxC
GNIgKtBx3L8TeGQ/nfXcg6mmpoLMgu3XlgW7inma8DIgMMRRrDQQq36H+3u9lNEpPe4/gseUq2Ba
REHQLTmTBz0izP1rMIdsGgnY3lkqGzEiGOYr8V7yC3YSp9am9DNILNFA+ljvSp/8veaLRTeX98A/
pdJMQTQr8pymamV9/TQCT4qDNv71QCRe8Mp4PwiEl+tjzHFlVSmLngHADNKIdlKSiirxPKOLnwcm
frmtqaD7+8f9x82ypWzkjrIB8ygOskV639tJZvact5jfaL1LMqXsoW25ACRdpxYGHoea8oZIjmEz
w9rdwey2FYneU7K5G9wFbWrsvQ3DDe+1zPxpNLCxPVcuJfQJLtL3OopnKvaN5LX2bFkgbU5UgxPf
u0VcGwDlFexF8sumJ4Qdq3T2IHfOaf7vmcHK4qxFD9lLijWEGkLKMcYOmOd4ygOUwpjf8+5rEqvM
OxVv0hrfK2rCMnukiBdPR70ErCYhABNd2tNdIeviygmXI68r6gN7+PHaGuK2uMWgslRJz4vcjxzF
qAqJwwFzy2faMQ61Vc3fzA3G/gefP4JgI9vwW3irOcen+mGOAsheQops+U2lZoZMbz/i0VRkheCr
22oaj2SGv/F8w4xej8kBhlRMeuZ4mXygLx6CjnJyE+/eaNvttCJkNMAE8Iz+iyD8AMToZ3GfuiXg
Rk0jlJMoY3K3PuC+uYe5eiIVTxvp89ap1H48BTybGw+ieomAJIqfPJeOB9CGzPen6tP7RlGyrMT5
h4VkrGgULKgKHf50lN/UP7/1pkKNpTZw+sMRvkeB7WyWJGcbifkHml29ueX8XRs5DsdgXYq0cwWq
5pgva7ewoL5Ru3CdHcz0BlZnAITDcK+4ce/cKIMhL1JxA9knfx1Wy8+jtPaD4bT+ePotxlTJytGF
qiin6k6GNqbJzpkwIO9PbpeCA3gMulGyQ2sVHY6cxJxgdl84KocEIjeIUfesUGK6/pDNMhL6UQd1
IV2CmUNOdMdtXeYIhpbGrT/PL72YjwfKNSXdPcKrLEAJV6ltx6zasufjHhblmRLMaycM8Ze8RSkL
sxhenYKcyDjpfVp254G88Ax/VRmCXoCE8dSQGIMeBpBU9Bl1Q00uD51seLzAqD+lrPFFBdShF3eW
c+9eYNBFW1Ot70Rlbxq4fu7wSGvxEO7zIgOJmq8yv/rdM2qmFcfHTQRGPsKdu1utnzbua9/8Gj/E
t5Z5K/koQm+arJtSPoyTyhxuaNhmNIfNVnn6LmEpSieFGdvv8ZYHUqPG0m7ZV/hkMLBgZrJ/P2QY
cs0k0rIORylZR5H4V81uzTOTwmAqEv7BJvlBjvV8lwWSxxw5YEEC+qBUOOmA1A0gFIDqkmUDa7kE
aP+88swX6BS0oGEkuOOlQty6GTK+atBdq7vq4QQ8hKy4nQcUQ503kS5BskPH41nCh6aRCXAfXDBE
8+Yd7CE4eTF8gOs5NqA+0Qqld9eoT8WAYxVLiXuM+HDbbhBO/P88/hAnbaQsJ4yAxTNbRArb4Z0E
z4zTS9dE1bp5ML1km8S7PUe+lfogJYMfZavX4srpyyz17OefsgM7QhoQhChd/4lC6L6c41SEDmG1
ol+3NhT/q7BWc/9m6rSHWdK4f7PaQMKkhACn7LPP+beexwsMvN83Uwaur5QHuQpsq/VeF5cIX+SW
qhZ/x30/ADqnXQR3OJvImHl9kvWTTmnv4RsQ4B5DkUXP7V6wWYcyWxX3+8Z18WjuSp2EMqsgxhzb
CT356AKBzNK73quB6AFoKKmVieajRMYFHVdcvH/EOCG+rGhWY6CVTKX/4/Vvx42bCjzACsqXsRcQ
7DoxsMcK+yq5Bj027bux8u9SXeoQpFO2327dO92kSu5EubSqC0c8hUUPGYpNQ5GMrkS4R1gwIaQP
3ilNHH99GcrXhyRhHuGmaoLrQEh8iqekEaW93+WModlwwT5ZPkesx4iTebIBCC3lpmw2YjH0uWUH
jL/8GWkRlZIeZSvss2B7z/CbvVTjb0ejLYS5HpJoR1N7ZZxryekwcqUwc2bDnwMcnENpMcMTXAro
oeunDi16av1oXe46ExfPn994G59LC0U6kMQRhZUMaEgxFbLW8z4Yo0LA8hNcy4QDhxEpp+OKi6L6
I3KX5N9Xuwy+k8w3FCfDEKqEaZ/H2MB/Gb0Y6O0CzwrH7Un5c0idFaMZWwi8C09mfIx9eoO6M4J4
6tOqR37ioc+XHUFq+cVTIFa9xXIpZOP4L6SM+XfixtrtH80FCRPCqJORppIoep+ZmDy3AlW0hxJ9
moGQEJI92zPHmeXivoexeScJmykuO4yCDn7lq+t0tJy6Cd9QN+iWmOoFSAjhGSX3++4UpEO2JY3L
yMU4JMNCpCyB/6rB5WUnbuTwC1THzJYqM+GGqlelLQLNbWr7mUcr8cxQYaCwqLx3fp2r/IfF58zV
Joge1IhvgtZh4Y26CZQ3VjpXPlzVzbkC9rcGqYejHn5KguH2sWC075/tAMH8c7oehyWTnOE3zZKu
aywQlHCWfW+hEh80wSFVa8SChI+a3gDiKpotIUYSj7EY8ZB3S6M+jkklSOxRRRCELWiNTEYLNcns
KDvMVp5t6VgeIAo4YaYd+0PhYueWYwBakfhyRhJhXquZSjpRHXwBwFq6i1EizJ2WgIMkXlapumAh
lC3bJj//rYusiSMrdMzfaPenhrGTh3W4uuky73fxI3qa0xTVDBWUhjsfNlPjmghM5zOGhpOi3tlU
AeFQkHEnA1OGCosNTBj/9Vu9IYDRYcUZpVB8MmjMkqOnVb3llRhTHBTKlTdAD80TdY/iWFlMZkYb
hYAbPl524G2aySY1CjCBb+gsw6dEe3/i3ZP1s8eI/qtH+/TlwVXAnmxwDgMVTbmhyShd8l9XlBhO
8hJL4BXqrvFVLtI9BWIX89+C5HASYNroreThz2vtriGlkbn2g/ABJwSrZ6VBnS/hB0+byJssI1og
iAlX11dZN2RiMRyjR3SW6H1MrwA6nsAw+zUiIbtKNDp/Vjtc3gFYVlsj59UU0H/RcbDEeVLBfczO
SyTnWpXACWZBD4saIhsPJQszx3F1vaN9InSlKbMOqS4r6OD9A4Z+xEBEuQpxNtVn6pJPAFfdRARk
4+aV4rhaUfZAEYcD+fv5MQlj7fgXTYBwlDr0jAcNWSeIfWmOAC3xS54/XfX+D5xcATuNZbnUx0Q7
CciG/48YmFpeduTS53dRQ97t0zHvDwoqHCZbz/bfOYw0/gUYChFX0JmUFzWtME6sepCPnalSaG18
4z9Ozotot2nnsE1GKEU0r1NlN3iV/reyjmItHs5E9cFvPMHoYTD1mGH+Bw8Fj1f34ynPBJUpplvD
RvO5/HXak1T/agWHcew7n+d9YMMpuJD9WZbbFKHni25cBQK0v8FrzxGpyllESTZg9HvCQn8j4b7/
RNifgJOYbAB2bSBQaxW9QcWcTlzJGMIvNs2pRADu4bYOer/cg7y3h3hp0YTB6+eBLyNbWX3mBMZR
4RlxZpsLI5wxGAaaemh3DhPXoafpRdf6sM51crbcMcoXutjyLOzc/IWUnyJNi0cA3r4yiT3/pkNp
LemtP9VQd5n5j+d2Q4P/KwIdWWlKMnzWuzvFqSH9jeCC/t4BggCpUPGAYJGSj+u961398iPVrxdu
DkaEwFGYDOB6nPBAUCkBnTrjXvpV9XcYLUh5VqZyu6/hiG069lGWqbEVXkdvqQ4NPC3XdpHAONNl
tT7xw7UnyosAesXNFYAldvXq1SQw9G35tBWBr4M1OJ1PGaIaiNArvnc3QxE1xbsmIAmCJx9QtRdb
75ysprRefl9gpETXIvNtwGAUJQ2kj1uAaJxbEzqPIZ2N8UCbW1ba80yt+PKuj8paooM4VnS8eG+a
tITisitYCp7rEk2vapNUhQdRDT5xGfI/ytOP1N5bASH7Jla241p0H/z/yOE+R54oNEkI5azwhXIX
VGrMoUQgl12Adf4MMOSOHJdOwPTUvLZBCuDSi16C7xzZ/m5s41xb9zUTTp29zuwKL3B5Qylsns14
wTCFCxH8hLhkNvZ/OmIiaWmNG8cZ9lwT/sczRHp5HpKGQXYwOOu/Qv0apLSo1Bwk/cxyuVAKKbls
w7GlTZHeTNLNJaidQZIbD5WGvs1lJS91b+fnalDke2dAHlEZIWT8mAoKoLAGMkP02TwfLSYWW4PA
KFooHnE6aK08d2r6TS1BJKkI3mEaWJWOPoZa8wt1naePC7ZrHdN0kT8+0/bzg/8YHi0OEfLqt13n
1rSD5pVLXvMGy6QxbM2RIyIca5XWxbaYaN7QwyxHBLl4CFShoTbSvn0KVyf9zHZFURK88urXownf
EynlwiRrRVhBkeS1iUwA1leCe/OEf3X9dtIdqoHxdOkHfvT7XAM3/TYye2KW+BORwAPpXVEdChS/
eoccaHFw0i93sszS5fvFzUc1aAwi5N9pfCACE0ydRDEHSroytbEdR+UPpRRK9Xj0tbFaptQtBApI
e7ISEhvIRAw/Y2y7G29Fzujn1XIOKk54CvaJa6piWeVdfyCh/8h50aLBgdLhIAk5c1DK4ChVWnIb
AnAVfx+5HfHNlnALXqJJ/HlsYD8N2Kr8Rc8XWmPVaUTpngXLAlE4XUA+ExdSC3XgmK1N33mCuDSm
2BzUwRJQH8kTYCEDnAggI85b1FslZsWQL5eTfy/3g+UlDZFlSBvzI1Cd6BADuqOg984+IGZj1S3X
VWnyalmN6ZbQvCCRIdmkfqPDnvjuJRjFZGl9ALyuyeUB1gsX/DsK+7I2BC+4ZBPnRkT41NkRj2Hz
bATRtuN15m3L6sgtUGCOzZDyaLUS5jkPtRAEVunFEW/X82w6H/JEcAq9kc2eaqO7K/G+WWKObIVr
EY7Vh0/dpXAQN42GQ51Mw1blLWy6JPX/xkgwtyNc2yTPTOHI6KHZyMK4HRKVC7fXABjHgBdciypK
rVvi8OGCd0mirv3gmtCT4l5MBR/z51aJZOVaUcCIP3HFF+queqyROAmHBtS+bKDjGfOFWsq9lkB8
xv3VeBUzPZv4vp1xrvm47Xofveq7IP3L07p3BdqP3PerRCDDlqkJIvIFcrcVsJ9FxzUN/ibsrdBj
stNkUvZrbTSS5sytdQqXeehGHs2hfstGF3OWWsKBteFlYnz+ONkzOnoxciyj3YPM8AB2mNuWO4mp
5WSe/7n+lL0aUf50/N6NFU7sna85QHuqOHrj7dwfPZY6czHGhxVXDqL+s+fGiXBC3Jfkh/dlgijV
FeDbpxOTemYEuDvk792HIhLTLIdfBulu5DjbRZiN1fIerVdF4+YnJHGebdnQSMMKwTYN98RluEyB
b2fQDW+A9pOd0tXdoJQrHEPYgON7/dbtOApipBA/rJc8BsqemYGt2kvFz1NhOqw7Wszo4eZw/i35
7WHHEFn8EuscasPQ4bD6FHL+KhB2pJKh1XHUXGUG3ufvCIit+de1X16qc/YWitrnQ17MxfdxfeDe
6jUbHTj1NTgwKIRJ6IFr+bAqAgA1kkKSV4VwWN2PhM5+TVtX32dHHn0pLJUl9k+53Dohj1VBH7g+
wSVZthfQL936jowqiQRIqd3tsiqW7T70JGs7V29ea7l4TOhC3rw9MfUsJlNQC94NPX0P7mAnmdeK
NsN5xWOBynViE14A+K/PDSPHsxZqsdL75G1yZz+bW2lBkCYIoH0heUrhjpJEI/5s7rDlbviBYBDf
KW2YlXSOciJ23EQKSmBZ2QfPBbH6zRetYe09T6CfyVZVejbPkKawxqAWGn8kdRkR5NDm4L5wmEiW
rXz6eYxRQXjJ5Y8MNmGc0eo96KEJuN5yQ2C+wzG57vqyen97WHBZR1z2iI9QoJxwFOheArMT/oa9
1PbJYTwoXBeMfn37qXLlLgnNLOrxIDn/CsfAuiosTnchmTAzr0Jwrm9ITl1OpRhz1yGE0J42tUtU
v31yYX1X+F8i2ey0HSD9OsKMGhsJ0D8D98j1bccB7H+fb/L1922E1aJ74RJftaAbPcfviiM0Dz6o
5fsBEQBw6PQ4MgPWTI342zamHo/u1UbFhnYxL0q2Esbvu2a+a6+9kCoKkG1GYp/kOL2rOzqU/0Sq
smz48jhYRZM8vbpooB243/wPV1BPAP6UQOXgfuPFU4geXafDYV7pFQ30t3575HLAH6at5b589TEr
flYvTlaACzRKYJG9HbxRlbjvtcfCYSxhOA3wt8svszC0cCnqrpHTU0qPGrzMsgsPVKF/Df8DbUE+
t1UWXStYw0uaIJv4oJOtR4aSACHLeCE93RhkMfDGaSyl0ElGBsB3cQiIAkvVRnrFotcBzdaeOrtg
Em6LX7WIYcmI026HJMbYk6Kmby8HDQf9EAU4bee5MHcpiasGPXJ28DBxW0jGVp1kooyV4e3fMkv6
rab+K8mHRQ1jRpt6ogbWqZJQ1yOixGgUGi+JxLoRxK0dARt8rLwM030kXl1OnKWyGz1CwKQ6nByp
Iza4uLpcFwUM0VLOzWyKy5FpA1V5ri5y7HraJezxU9OYR6Svdf7MnR779yoZ7Kp3Q05HzdxRUDhq
rMBWX3y7bSuJbxMjlNK+b88HtwdX9L+Gb+VlAXHCOdDhVGlZQZ413QFl5tvpyaLAVuOJzHS6miRa
8JjXz+2HVcab2CHRpAodm5yOmeDiaoenMEs6R914AFlckYEOgcU0LrlBoQkSuzhw5PKAP4gxEFXP
/eYTIRN0KXcC2aWaOw8RHxrFy/NFeJNJHKQ3mfE7sJqhUACeqxpn6ZrS7Xw7GCSSKK6AoJLP5GE3
ljbp3NBruh/fZKDhjCAugKzmf5KIeMMfTEkoB4TxmhYhC+/xiyrP6V/wu0panTtOz0g+am1sC7vr
ow8zJ4go39vLIdWc+MGSxYOz34tgCy54YB9Qz5yUUO+VGNnHDxlU5vVP3dwKKEnxthhNDsmOPSAf
tAU0lhhtHMG42qg7/EO2R8aQGOlAZInejugPGsCJgkpbu2dcSfEjjL0/WyEhGih8O0GNET4O0Ov0
rMD8jDqEkxX5mO+Bw38asTg48rUWLlpBWzyCd3dBlxVjGRO9/RFuCM8gqVMCFTreO8V6Uax0UTHt
2cwKAS2/DZGBpxiscLax4btOyrLLvFMOKbXvoUm/hq2s7kGoUSiQajn3dpRZQUD4TIsTRRbD4PRQ
2BTbPPOvcQ7YhNgLxcfjGYRCpmAbZEAEIK4nPCtygt7/36mcSfTIq94yLCRQLChLqPc0eMe96uHn
NuZE14XNmcIWv3e41+bmPkFDpy8fkV9yb9lbysglZVf4n2lES9jBa/erauGqcs5g6ImravDZObJZ
3KCXxH3kucgkXCKrPVGYgUpgXzXUrWRQB+OND0wNS/v4jkgI/k6qisa2WRcDPsUv6HilW7I9znAE
FgOBz1WTN1cMiY6OnO8N/GmUZx1kfqog9yE4zn0RJtG5z/Rth2vLPiSRWmh9xPOVvxcON2LkmPSX
Km47BnNOs6Ll7NhDBDGBSP+EtkSgVfxOilOKyrYvxF7aJqcZ1fY9zmFe9WMnhcS700+T5bNedxyC
CJM+1Lj8PWKWJlZSkE0MYLXLzyic5G05un40zS+X+g1GgiyQVbcinzmDomUIBEFspj8T0K31aq1J
KQE9baSIH+9qcuu/Hn3I8GhV10DY4Hg8kLmbh2VKHXgrmItSyR5Mnt+cKAunFQZJRLrSqx7Fa3hy
K7988xa0Zf6F9GdHblB5H+t3kYXKMbDqP+H3EdTSjRbtGqYKdnzvbx7FQoL7iqheh93gBmZAexmf
2JAfCcE+8nPdABdyiAxL+qcKjWDzeG2ww+YF3yUzDPfiwTW5pio6DSY3tJjAGhojoeN5fbmWVq0q
FH/wzyTbZvxGjDtqalUwpKZ1fF8ZybpBu/ZXq3KKQs4hmutXNZ17rH7FDCs8CW4KXC9rkfqI3wJ4
HedEBs/ETmQFweHQlCKmuvSDKi025JcfpMiFqV44fQdqdrMpvErylbZbvQ1kNyOTtpzzgrVEA4Bl
O0LoQJJ+NeeDMULEM9H2ZbU5+E6S7Pwry8HTWqRd5lUsRzPLUE9uJdVMGFXAopf9cHjodGLQmJT7
pcaAP0fndUT1w8yvOTjE4e0O6+pA/ipDYIdchW3YKvveSyD2NROOpfwDYyjpAK7nUw0BRrAXUhCg
1l/dHdOnQ1BvtAcPsVokPzhtKzc8N6a7iCBdkyQL1LRLKrWNXxH5pCN4ZwsBsl5fmX8CXhHxKP2f
UVOgbOCFhOqEPitP0WyWR4zQ85JkJoZdYgVMqjtBsE2U8NJfWfLEVF7Ob7lfnq8i3eEfZvAzIMIM
1z92xzL4dQyz8uY1Jr05MJ7oUsyeC/H2h5DA63KdW+lYN+aOQ6Srnfi+gggSsW/YW+V4y08WLfI2
Lo+sOJFBpjUHxIXDu3+m5CLAqu9G6ME5fH2wvplhNbqndxMFy+dnNCZmiekgtktEROQZgYi295ZP
lh7h/hiGyWnHH33EeIsPHy7uH59Ng8NafbG+K8KiHgaHhiImZh0hiilNPJrrJa4fn5/Kh/4YrryH
GMHuAoKzKjL0MNdoPYjsHn4t1ndB3D1EUZ3L2rWQOWi2kudbzxKIxeUz5wINMZiM1F/rROw3iy7l
S5thzHIux4zGt8qwCuiA0iLmhLtkN64L3m5fjmTukB2GZciNF/oR3knRKbQnc5n7QGaykrCh/ZLw
V+qnfICAsjCISU58PZBRonyDxVSH1Y5tQZeAW0XW7mOI9+qty7VYj0cbgcPOaDm0R3EIqpCSMkcR
6y2nudpttCPIEKWiGO1H9N2r/FEN2zYhLeTVHolcviVOHEhczRB85k4o2Q6vV5DcFhBOs3LCIFBZ
kxQlIrQx2OFShoOLp/df4wt6OjBZHG4A0TS4NqNHw/s6pG3Yo+PS0CAm1rBJ9Tz/8FDCSqozYvcN
vR5l6+X5mwXD3Jp4hk20U7u1tK88fEv2+zPudvzvKebPBnF9Oca/Pchqi6jWukwhlg/w3Zpsriqh
Zq8cznddwcYhQ7CNpgy0j5kSEIGA4I2ot+Nb/LLp4a4S2kUMae9+fjnyueMfNADgsTKBLQKyNe3s
mYyOVyNAGd4WttagJfamzytZ43QAh++C3C5H3mQTHTTlCKtjVPlPyQROSRxPPb9AaIaVxN43UmLU
hHSaBZz4nUp5HC7M3x35NmE9lKWwnksvv1OdbLvZ+6DRG57G+T7Riw227gkHeJQ25AssvUtcNgt7
D/cw7s3ue9sG56J7mtWry+y11NOfuZzO6PwgdUhVyzyN0TyBr6+pMfide9IweTRgsnrnF78Ts4LJ
kQGiPUowVZ1Tgo9G1HgTu/BQk9PqqV9XHPnCAyN6rETMHqsDAEZ3Fv9jzRFj0wbmdr1ls3VDBf0i
RR/aNwYW3UACyAT0oTB8GoLhpnkHG15P2027hxEED+5tsTzxmwfR5vSNv9uWqNt865jOJ+SiVXhT
wtbbEmemFgImDkQyD+hOZ9K71Br7GQkpMBoOJKq+nJrnQDCbyWGe+qEg/sANU5usebaBioCKd8ju
5d4cuBjbT0o2Ux36QIsGCBFTOG2Qp5X1d91MfKamassE0efvlyqNBnQ9obaIoZqyh7aosU66klbu
6Y+tbz/selnjRq5oW6t4aTEk1NFcPL7fmQO7wLS22wEn32aW1Kcx+bFClDJSWmXpBIwjWn97LQME
GlGFZd9B7rxgU6Hp65vdRQ2ZRSrasmVC0w7D013utZJZiaLzFdqW/K5NpmDX9HRZe5oW0gnTIzkw
cdD0czeYi8Lj5b/pcCjqbD1/DF5v1JycpXHz8W3nfvSEtRJw+ZhZT1gYYNIg+E/588QzGr5Clv9t
XZ+HNhTYjgmojmP5Ps17TKT9n36uDysXJ2VAefkX/pyZGpXKGVVHqU1+qbbqrPN/0JJOl//kqucz
xcr3Vz2Fm5M9sywnFfbIFAbHGJVi3x1GCBJ7rjwp++swpbyx12E60jodnDgE1xndKyTwThwsn1zy
LGBzBgB1CYYMeBWCVkJt6YgGj/XmILHzbEByC5pEnrwlsXThDD6JfiMOnX7958Xkim+gRvrlm4Ga
vytVGd9ApOPnuc/k/WvAuhMzn4uqVeI1393qQwFliaewt9aGwznHUaHMXdDZ/kPSzr1OGxvzq/gX
KqYDlbMDksvnv8Wm1zlcpBElqgAsIxvtVLBgtaljOD7wMLGXEyQ4Zb1TgghWcWA53MFCNYKq49lt
jwM0b9pE1I1yXEUhe8TGgZlbhmrlRehawfE9vqPy630ro/LMP8sfnMIXGHXMVEpOu9quAFT0j1kd
hyMtVz65Z1+wGDQ1kaIFvF2pXrs0pWG4hvQeema8l7hpc88tDMsenYn9HnDZzHl0Jfdxs2/2xCai
GKY8s/fXFmK8YKteVq6vpEBCR7+TbjNpmJyMvD1WTJsagbtggLoWeI/BCPqBLtleVZKzfvzF4Gdi
z/NmbNBBY46JoGIUt+7xriKn8tayse9Bs7hmN0rHbgY0tUzEEjZmmG2vBV8c+pweJaQFnZFNMvVh
MWPMmPHTUGyW9ypvZ1WOKJp9Pq2dByHWUhDRsEDvtOv9VC1iuif1r/Obj2xyiSRndRl/IbQONQyQ
aCV5+wdbOujT2tYJvDtYwk6GtyZr1rwAVX1XYvZ898gsF+Ez9EVdhkjwN15B32iFHQiVj7uktBHR
3DODQ7OQ4Yp8E268fskGrHEPuTu8I2h+Qmzjnw5pLxNonN3hh2KVKXri6Gm/7Pe0jK+HQ8ZZ0yJA
ACfu4iin7XEOpqe+yaPI9l7e+QeC/QfL+KYBmBVcsDsHEbpfxnJOAaD1C98QqB61+KUFU6EMKqAj
KPq6BxpRdIKt5OdU99nd+eWbBECZ6h/HFHqE5OmHsslzoSG2tXPw7u2AKwcwamA6GHFzAT8EVC5T
0aINZ3jMnmFYUlpu9cZeBpes0uLWI7dG76xuUX7Bq2wz/NKGGGNDqALy4w7y9zowjJI6uzjombl7
+DxPI9ZQaWSZCFYJ6PO4dleErtdGrI+2myhRO3iGfeBBFrTMHsEipyedIxNpMNCK5kkmAzzvkjUZ
xtgZfq+VSKhTXyvYnYpPTzATMnvrZQma35wa17Of7wp6hiyIJepT6FygR8wgbUbxbrlDejp7Q/ji
HjNcMj62o5wOty8QyYR03qeMDNCV99HfCQQ5DrGkBmGtz2my45LxYPUrHhk9RlAekB+czO5Rr8bL
HP5CLV+bNbwI26xCn3TIHVxZ8g0+m5OarTePWKg6HfVo1ZQmg5U1GotdrOeMLTs26ehYATjAu72i
c1uOI0Om/pdgGA2mzXGDva/AGsjjB55kuxf9JAeqvjpFlp9FTXR+h32ERzpg3U637TycJiV1k5Zp
hFBNhh8DFs1/apQKqmUzPHRGkAvD3j2xyOkXUqNhsLBzEsgAzmMDWIJ3Dl5xml5ymZUw3CPDPDLL
5eIoRmuqJK5Cy5aTKWPDoX3moAf1HzL098snD2uic55S+acdVa6FwxhqCgp5hZGn2Fj/Skr+T9r4
rbOUQdY8H8a15vIAx3mpX60LiECcTvlsG6QMfTMxt6nwh9k0NnmAdpBsqjJZYNZMXC1hDLyMRIV/
PtZi7Uyn1QX1PcFwyJkWN+gIig1Yz4F8BfV/o1X5Zx81M/YZyOO5fct3Uc8IHGMXp/7D3dY1RIft
jQ8S6d/erc73eKomT1pcNX6sca7X4gN+dUBV1t4TKYW88/IQPm2vXaLq23H+v9K6klVcVmAtvzzQ
Vq6hK8fluwiLK6Clo9DNnw2LUss3kuTZIXRHpBzLPdw93qa1JeSwdRptkYGuegTedBMWzS4eK/BB
eyqnwZZhWRLD2X3x6oEC8DhRBKPM7MvPGMc6etitwTcuApqDk13GKIMD+jUsG72rqUr1T+/hWJ+z
aDcZkFp67+OEFOiDNLmw0gzov4YDLboudnaquU2wwkw/xHf3ePfh8ezUTAd1OvSMhP5sZnoknX9O
6IjZ18q/5D/n0/EUiPY/2/bHtJFsqHvz8s495VuHqHuTfiQHsQiTFW+cqwbH/Bd/XEqUJMBqwfHg
kf163yuU/tenYh+01BDAaOb+LY4xNFNIFPGCgujytWU96uSxSUG9RH9h0NI4mI6qVJU+XavimGE7
COyaPq5ZzD58AfnbobbOHfRHhmSGYtKOPwz+5nd03tEzFBHK2GT1hr+sletnR/nev3iO0SXvpVIw
Sjkhv+I5t3l3+VS5pOLvDt0sLaHIEDNv/D0bth3BsRS7FHJKUu+2wCfA3rpGWlIdGhKstJySAcQo
cxHAP97XoWq/N7ZjdK4T6SIZjBoq6ygG0LMS2BlL+mL6YubMkxDa2E71ndoW4Wrrb3K9ZmtzK5C0
3wokdAOBtfEdu5520ztxFAd+xHQVRulrX15NacoSM6d62Wbk30zdbnHCx3Ne6YJRmSpIkIe1PPvk
qZtbyanzovgJJI5THN5h/opFDS/PfMClJHSWtluI0hlReo+F13Unz96DDSpVQMkMz4jxGQzwEeSf
ymANOmRP6oR82Dnxp/KnghLC5newYVKtojpQt7LBOXZd38y+UiX/O2RxtYd266MRWWy83sDMSYLR
CC0xI2F5nbSqKr4M9THDxgL2xwq+f5oOqkTlZfUOVlzGplu98sj9pfXIFFlMDDEOcxnXIpzqamFz
QO9tt1WK4YKaYDynQsv3ID/HWC+T/gVEsYppkDCifwTSvBO0ClywJ5UmO+RgUE8Oa+qzqgQyap0b
15wWw8kYjwh+sMPMq58liSOVYtU8pgM7pwIxl7z3meXts850CKxGCIEgqj3M6VCyF7U4jNAdpeX5
1zgFMP0t8/i8dmcF/YveU6JLvwImoIma5xE69tOsrb5MkuTxtIS0Gb6t11MiX/5w6jw16x8MZ3SV
DgpQdqFxzqpsBKdwDFv18y1XJvlrfI10ANXs0TWoFx9ZLOwluGowcsKYggxL/sdHu+De7KvVWUyp
yuY4Mbp4qK7Gn9ZEoUaFl0JW+ys1CL3hUM2tBRRriHh9WqFe3w+7upoJPD6WSoewXngix07CNCie
D7/BL7moIMn8maLD61zkjRf7kJr6QTK9KhqRx1M4SUU3rqO8q7zSunJVRv2o6OAExLzWhXllNNoC
vYh0YBKCPGUCEpR7bzkkKZnp/JcZT1VgGodf/4+RbPSvlLMr4/I4bnsWroGJoDY9vXMmBF2YPNZN
RSvbCyyixvAb6PSaE5JglTn+yS/+LpNcZGHOLthBPi67C5TBC3hVd296tR/7vQf7AcwjW+d5BOb3
Q6aIR9UA/VRiOEJj6cQHicjmoFM4dGef3IMA96tF9d2DHED5I2iYUYpCJKLtcNWdPBsR1g+ob9gH
LhuAbrVENZn7g9dbbU3Zruj2TRwpaISFdiCr++2blGqiZoPob9ykxL7THvmIOsbAF9jgE675O9tB
UWNaMkTMyhwbisIdtxlbPxbYD6XEpsnprAfbBISMtT0qnrGb6RDz7D3atbJ/Fn/tp1Aeplhh/olJ
yT34/tWY64wb5cK1fa09wdtlX3EqJkzRR2TV6PTlxQhyQImWYE7onRcYtBJr5XM1haUmpypA0wz3
rGmurVofwwQrYftTkOeHu7AKAUEALM2DrBUDyDBzZ+S9BpdOyeqyA0wRrEuSd4x2DZj90GYy0sSM
ANNPWXJA6Y37F318y2Z5M3UHyvNQBoo6EfR6YlNzcVCG2Jbif/nwDOs7558yNN+LL2lKiK2PcH8N
BfouApa/odRZX9Wx6Dc8k/4RkSzq+sQzj68RFmkNCsbZIDOMS6pdbFuxLEuB1Kjq/zcYB52Eu7l5
CNZpeQaCtb/SE6iEJWnST5SXzS2PoWmnqjvlswPDKAqiNNq02hADUI7RinlACJCow/JNkhDy+93Y
s++WuGk7X/Z/O7m9sESaXqLW6FQvB4UQEuoiVQIeWDPj03lzUd3nlTmN2qh3ksrdJcf6tPqxR9Fx
QoCeyczmT6oWlnzB5RgNPkehh//7YjiXA/1VukXTCIm+XPtr9SihRqVETw+wleer3Vq6zr2IpY1l
0AFUnZ5aR6JEJrtQnc7AsbEa73Q5vGteECjXL612rLwuXpvqXPoBpViY05wJ8GKZNmXEt+iAxiCX
eukVtHI8+dGZJ/a7F5XtDn28EjTFqSxVJ3hV2lQNoMIo3B8LP1wXBwqHw3GMhRUi80e3nfdbaH+e
E6uZ/NisKdvYlj7o/YOUo5GWq5oBg5KzalmBOBnzQT6j4nTSyfpFgb91XqMaR54OfG3kNL3W4Rvj
z/DNLLlBzt1TUMtWGk/rzlRJhOhaHfspCTkJyRDqGH+kGA6hD7EhH8tuzHJ1Y+4nuBy68rcxL/jA
NMUwOtdx4FG7WTYLMCe7A+4gAfELUetthJO2QvpYZz/wkYNx/xMiM1CVV5u/Iwx4VgTJ3BPzGCng
g3KmArbKL5HRqr4pET1MgSwleAIWwoiUjZqq3ayM7Kh8jUVm1hQS0nqjX/kkHDCT76EgNQpDQZKJ
/3VEKf0JzjdsAn3vBfk8nH7dfS0EDFKsow0j1yhNW623z74c6/HugcHMCCdWH/asWKnpll7iknB6
GWw0omWqWMRSzWdGKyCkZgGfDksf1n1oUJr11WdRCH/SrakusMbbcREOup/zf0NVUX374/XunS2M
+LEHeGG6dQS2C+tOprivCyrcB7W+2C7n8+ztCBTZJSp/acBKujmF+frlRwMtIlstEIkWwQYScCpF
jI75jw8G2xXZ2OzDjpn8/vJeCOL5grykvA1zoGRfr71NWkX43rD5PZdxg9rrCBNwk/Or2QdwbAv/
ABLaS4z3HhMvkRHdQvxMsEtMg/mBiY7VaEkxnoekikKJkvmcB6cf0wDvrIQJJ0iCybnfUuHwbn0J
dvaZQKPWSomdRA+W6IMjUReWXr/xa7U8BoANbppOUMccNC1LgmI4GhnCc+cNUCrM2jm60gsWLHJl
l+SpMUGoFHcjhZcVkC3CwlNN+FOHwB655U0sj/Q1Nz6baab6deT3oO1nh6jYSeKYdRm3AzA5TnAZ
9Fctlbn96GMdAbuKbSs+5tJH/vQ69QxDctcZqOgMRQnG38V5vO6h+rywVEeGmVoJnQmdSOmCyJCC
dV5urGPMhIGkmnSRq8M6O+BvuA6nLuFEl/Uu8bY4POdSKe53+4KMOnOJ/1WDgMIyuUWp3rUK/XMh
b0YEZxnsngHKDKBCyH1bln+vo4vlelaj0+CAtjiJRRiJis5oED1rVvovnuvCQIYW//FZLpiKKoNa
x2UAHtj3JnxGqqLRz9Rsdse8tFuJcjS18eEmp/kuI8WqkKLq6+GhzpNu6yn7CYQE2clJV7/rRTgg
3jnqzNthynqeq/uK0gQ9cthR7i7Y2FY+zJef4QgBJzvfhms//TnUVo6wf6JKs7o1817HovobkgMo
A7ZaaNmm+uDa1PHfOqaqU+mpuTa9gudruv3NQkaK8BOv1EdqNVisVTBTu5AzS6m0FJfgsNi/SSu3
XhTTy38tk/Ex3mClpD0M9Bj4zUbOHvEenCsXoS7bUKpwdYEM7XctltgOgPaHpIlHkkU1kcAX402e
8+5wtvKPJyZICtIcjUM1DEvMJ54JiBdLn5ChUU0yjw6T/sjPud7PmQb4nwll6ndYzrHtsznBnoDL
f/GiLZ/Qbg9+8GhBxQ51Zxr8SrUYhgOAV7ZUjNLCk2JisXA6kc7H4qcfSm60XPD++C3fcTaSsqfr
nJwKegwgsYwzb4xFyZjdEoBgAnKo0n+il+KpOemK/yIexDlcDis93IsFxbBh5eujnhEy8NK4133i
j0gqmwRl8YMpkyh9XbuOc/r9r56k7Sfsx3GOs2AG+m+2NCrEd7SPHQCkzAozBbAfYN2U8zzTDwg0
QkChV/ZxHCaXnBlx9Lusw/5OZXEDYTnMejjR5lAbZ85RgrXidQpxOSjD951uXmnlL9C/8ZNY+K/1
+vyBUAi/9VoI1HqAmOfzdy9sJVnCiNBsBYqwRyc9TM9r7OjjKiYsaMaODKyBS5mdqVgsEZofnJTW
C6omAaLUi7rS01PtWScvQ1FLBGa7oX2iIeXGm+aPxWfHUiMxzG53upPJ0HIaBjIOFcW7m3BZXt0O
zjBg354hqffZXkKMVfteJJGPUbcmnVXnAyVoozI5cJrwYtFYpUKodl0op+FBKWNGL+loAmpVEZSo
ds2CmQM/O6PC4Tcp7UiUHme/DnMl8loHcIsXxCfsxiL9YcjNOy9oH98NV8mC3ZB1tqz63lcwS16f
rU1yKTwBbBXPjjIYe5+9iLFLDMndZOHG5U2dPGE5zySCAI1TgPEBvr4QvP/PLImV+l1ruGGnK3iV
PXHjuwgUSNHhxyQWF7MSYbiCvOvBFjWkdT0unQP4+ksWXFi/GshSindYTCcmvKtYLbRMXEmoQy4t
WEfPHXXe55IzU560BuHus7AE+Ntb9qKrYAXXA337MnWie3i7ZVkflarQqc+ozCC5VR6TN65iAetY
1QCZlLnaEnZRr5mKvYzkYWUQvtBSU4woopTtRZUp79d+II3pnfj9yWsGaxQTiRVLHJhwkAngCnoH
zyYnVbD0hLz9XyJq98ByME4QiYAYSyDPhZM1HeWaj0o/tjAFo2VHns+mMktpcuCtnr44vl/FnW1t
TC4Cfnx/oOv2WylQrN0L4sNIqvt8IS1pYQgiIKyIqKeWtF+TspQMreiGm/nL++a2SrnumNvQC3ez
VRdFOMMhhN9Gbfm+69Gf27b9Rt/wM8gFoUDDOtSGAQjQLo7vnS6tdafE4/+kO2LiUcBaiSUYr407
F7yFaWH4vztFpnDBt1YlwGkd0L5DIwY4ToxsYvQvgtL5B2G+6fHnOakziDLvCtc01VTymt/SL3US
TZJ+OwQstAPunIzSCNepcC7H822rQlIDeojePkmBUqzwshoyraxKsCAiK+yvDOw0xIzWeIZZanIE
H0PTEdOuYwPcB/6jJvgqOtJY05lhzNxnYFijX786ahQBBjJf9HaFUdhvgKV9YIOQeg3Hj1nvub2f
yrSKhifdeLNV9ioVsEG8A4UcE31OQVQ6BMKpcRXjzBbui+0jmP+ZSyz9buT7aGfwYsLazPsZ7SSu
xZ8mDRFPBaapE42A+Ts6sNXT9w2waSgWE9PoOlSowVpCCQ09jtM/MKTqOiLx2DDUGjQ6Rs+JSO2m
Ua/W+1mAWUJMWLddfGBwddi/fjEKqjMazBkzvtrakd8v7BD7EfCdNBhe5uwQlojdIo6GgYrnJfln
3Lu74vx0Pi9uxmTHz9r8Fa/oNOEcMDh/N/w9pmhKbNdW5da8fqnR5kg5iaSu6JVua4JsU1qMUYJr
yAVkDLxUZf8/YKr5kdsRuKNQuGg+EumxN13oaIahFOaCeUlOVdase7xGAVQjWh+3BzC1q2ENaFoY
1G7DanPxLglwjlktqzfZL+W2zpBQQY9/lx7xZwVfquimze6oMIBsCXPPNsFR1MJBC7txfTqE3Xcp
Blux1OPB3NfdoK3ByW7VcIydBmAT2W6e8qAKGz8OAtavFf6tP4FvNvscezQuFksl/LrNqHtIIos+
mZDTrq7SD5Lh/U9jUYzwbXL/lrkFxxZAu+0vuNTtsiiW6+SiRBkSmwBvczpCs72B2S9yLqmkjO8a
mBRVkdiqFaOjVHdEZfom/6YFISQKz0YxiOKAS5kGhsD/fCbIuBhIcaLZQkaIF3d1LbyuiTl10Cmr
0aiAcMHDhRvWub1KynFCFxG0tRpm2QH6xsnOQnfAbE7/XHchsWXSNo4EKq0/TK/G/o6Pr2kMwVlc
bgpJoevyj/4uZNrybTWnhmkbHE/XvYMbrWgC4uBjo6BXX5Rp8SsjOQzAeLucbW/RMRRRhub9jWu3
B58iUIpTyNBgVbmROnEUUAVwB9iUVxWUfGS6eKRe3+Uz1RHzA4q1BsnqfqafPBwkekr7fZ4zdZf1
ZpAq6ItspTei5F+Ck6AH3oNW2DVi/u1NkK6XfJnlwhzyYC24329enAr0qkLt9PXLKCRMytcUI2+O
oCrrh4Iq0HcGHV2r5zvEK3BQDDEpZHMAlq3auKChLgZohjCAz6SyIgbLol+6bApGtjAX5hLpR4el
0ETOW0SSo6bAnGAehUrA2wI9zKa38hD/3vTKiK/5QQxQbueFU1a57t3RreU7+69Ny3kzZ9JGHrAb
4/P9Ygqt7Soj9Z/SR9yyGsM2l1vozg3KaZIaEBmolrCri1RaEX82p7N+8bAokzfUF4cPV7GuPXf+
pCXGR9BRxlLesm61S8gnMt6GiWWfUXU6OEvb7o6jZeGfmK0hfD5AR+3koEQ+wvASs9FnW7RALRDd
liWpaH1M5HonSl5muZEwqRBjxfoRcUjFNPSQhfnm/wf95MmgLVRp57Ggq52kvU24OkPwV4wicJ1S
9vt874vmD1vmBh+tGJqd128F1zZ+pagtvyvWoZRChk3QAV1A3QSowMTXrKv/EJ+9ITWgCbZFVCf0
aLGtk6dvyoBle/1rUHVeKWtTsKT2HuObw7wdXHTrC6+b9frLshzT9k5ZWRjAFCpQJ7mqzqXvas5d
vqIpZj5lDjsAojHvV/fUkm0O5JRQW93tGsjBl5TNRAkSWB6NmMDHQOurJz43rDCY7QVG1ZqF7AFQ
VPAJF9ova3RjJ5dvJ/do86mpo/UAnV6poOqBJKaEkYmOAAls66fPHIGMFm3c7xT6filogcpv3JBp
MAYPZD34ggcPqLN2NG4O6uYDacOGq5u727jymP0/SsiE33SLcGNMfGh9JhUlCM1hrU9cGfJPQ7fL
440gF/AL3TAPGnKWEMMrbD9ko4pslsWVQWOf6oSo8RxBRsy6KrASva8iLgRkVfMpYnKBio3qZF/V
d5+7hMvAwTEZOt8VXRl46JLC/9jR2Z9piHbfra96ShMfDmB+BT2MxFabnZ4jG3IBUsDl0JWVfT1j
TRppokX9W2rji2Cm4Lnz3bYQAzVXnZGmwYHl/jTLSwsi5YjxmoqFEFo4abPcOgeToc4y/bc070Sh
6CsN2IHC1CwobzWLXr0CCLeM6rwfvn23oT7XCZrlYzhO0/jELDaK4RW2xO+fXm2RclzQJy6qASLH
KQrPBaM/AOxu2LgdcCW1/cxTj/biLZlqVi/3IM2Nmz16iTyQ+GG2k9aR0vRcNykPtYLilo8v65Da
AQSpY4Toc6UTST6tVmsYnvqNL2DiMs/HGjZwWytIZAx89Qg6HDmeQK6Wwwjtp4joTWC8H/riv8nZ
1pbMkXn97IFuUD7+eQorLIabnhRcLdTL51eh/A6mU0VIHfHIK0cNuyaxczymvRsPRD4ykomP+Voa
Ccsoeo7XksV6+yOluD+AGJHcfW6cZhEo4sbG6f9J704EQNEkfebTkZIQ/0hr8roLAhbpbB9HUN/W
irufm8iiGnaUD3JEhYAVDBmcHC+DOXX7bzOqtDmkMJuZ32ihw8kiZj7MGLPCHsRknXVnZyf/TFsP
ienPYmuIALN/le/1ZQLotG8Szp2EmFj5kmzMUUitHk1yjxMgnhiBG5tQCIfSuOgYVGCRoOWgLdkM
DreRDgN5qp9keLML/P2SkVFd/Wr/MbVAzVAMr+pqgLmsGRaDKZ99+WVONvrIg/q6rhaqUxT1gmDV
0kmWxZ1Vsk93FzYLt3Vitr09dyGGXFD2uANA2d2U5NFMeP2c90cI0vm9SmCD2BBY1TIbsXvTAGi1
egSrK8FMzuuA0BnJzayxfVDE3kY07K47wu60wklTwA1SAjrsxL2GKmbxz/drMR9ZJgKkK2Gjpi0d
aw7yBmql6eFAShFm++wWBCnVYDJ7RK2n8p0q1166PhVj7cUKebxcEACqm/hT2ScDB0VE7xK6oEx1
HCH0Gu0gWg8JnLUecaqPloGXfbmfGhKBDZHafySENXMJmb7xsO+LwxPuN6/bMhbEr+N+E7WWlO5e
O6doKn+W53Jpj7jGlvklX+hS0ostBQXIsafON/+mUh/b9PQ/XQDF2L8vLDckbpk2r1CU9EVX1ecn
EwHhKJOsr0byDNNKLVIKOrNrm8gYC9kWUXgrtkIYZnK17ogahgkC7IOiigCaBw2OFhXV2aZK2GwH
MXmc5EoFdS40KBftNnWo4sX4In3lD6Jbmr0Ql45j4BicIRC7u7xIPgK2rBJq/JHKcI4+XasFbs0c
7aI4Yze7fW6wHvtnE3xnjB4kTfNtxAyEEBHUdawuyFdcjT9hFd0mdBPKnfL5vCLxhfdRZLvZGJS5
Vbo4SMdS0pXGSlLiNK6rI6qBmWajCKOKIteR6QxudhqYSkY4HH3BpmdCQmuWbJ4gdqen8jS5GrFj
Q6H3sGBYmzZOVEwWkawcCttGhsxLXbMQ0u0aGPG4x+IQPxHmImLxX5Aufc8Aiz39pbo5OhJM8c/6
bxoRX4QrVd82YsR6MIvyWRtfpOnD+vGsuEzMDolQv7Gsgk0ndPaUMAA7YhY1UH381h+VUEdBU5My
OzXzewyUdePUbreYHLYq7DfTPd/8L5aZvjDJIGI4+hTxZwvOa7IC0kuCuf+A6wydOVQCSh/lE8ye
FGlzHATkWTqYUg5UcxahAH4hf2P2cwchOQPSTSLgoTBAR5SwKIKFU/V23azJ9rtSwxr9nVX5tk+S
hvNZn5Vviuwa6Bn0jre9K/JT0gjZQBayY6+swq9bQCrCsgauTmn/Nh70RHus0EJ7ZYLRxltyybDr
eKW6gouqEen685t2EEY1dda/o0kpiZr6loafUMCpOBWsOB/f5LlTPZX+zFzPaWi7g+8ptJV4d9Hy
3vBiulbI5khCya8PE97nkO2QjHDfQhajBvLm7VkIQ6sx4hjV4tiwicJA7hFvcZbTcbPVHFy5yLKA
gZw8BpakyNAm37eQhY6H9BUFIguDrQP+fKdLZQHTZ8pAkAT0o57hHAm+7Ey0z0DVw3qbEHOzB8P5
N7wRFAUkTdc7TUCvW0dKnk1UmSapalGIn5IMs+cWRC/6vltL8CAXmXPl8IZOCoESSFAaY7eLcOK6
86p5NrltJiv3R4mKAGP6TNQ5i/OVng0mj2sKbFJsPErzzI8GvnLOKf50BIDYMWUuZvtmHkQc8Mxt
m8rdy0ZVYc5TQhauQrGvtxREK55RV64iTWWLcjNQSXDybK6xvz3DoNgSWND7TFf6A/Jopf3JiTUT
qucMDQMPEj/DITFDbYZzvkVwTM6sV3JesEdfs39Zop8+uT+4fzwfGWZQJJM3VL6SgnCfPd95iN8v
/G51NPVoRdr6inoB3uWt4in4gCJ65BGZ5SKGT0zSMxUUKefXt+EN6kU7tGKeJfxxhZE+L7nD+fpW
H9Dz7v3f7nibXwyPWP2ZNOAuGqZgWyGd1EMJO5OrTNU9xbVyGAeAm9yvB5kHQDIhyp9/h5UBBcwj
/6wiGs2fvvMuJJm7GJatCT+Az/tCJAtENqVpu3ufkW3BvdLiHQrKqoe3ubja6ixI70Q1ny/oRVK8
3yp3uS08M1T4FneTZNh1HYsTf/D+yfss32hQyDxPIIhABduLkCksa5PmWMqjdO69qf9vMW8mOrzE
30l5husxskpsAapRcFvyEs7IZdw3FOe2dPr8Yf7xhM2te0tZX99x3+42p7FCCIxeaLNcBOMj3pWt
5ll2hFoRBzJhgIeDPe0relJ51QYn1HmPOW9b46j42IXtiueK8z+LsiHgLv7kZKwrTwAgQ7XDSwa4
BNr6CIpEm+f6n7Yd8gjGCpA2K7fajWDcHSJz8fSoaBK5S4BNvwP+skIM6GcLSd6B+xo0sgFEod+z
N94k34lha8o92lLttVHT+XpLk5C+CptTwSKOlfSEZmrcEcItTJCMTwBsoUvAhibKr+Yuwzi24Kmk
KYqEEAGn//eVfGz9rPQzMiUjDIEztGSYTvrEIUV+7xQV6Ak/IlehsE0/Pni3JSdABaU72zZfzwNO
rq21BRCBLycDfcatYbMXOQH7HuRbkrosYlaNxraO89bijDEMJBX/GZyO5fhIWjs8I3Ef44UYMVyf
natuKNE5HZ+ZGNrzd39iOSZPUAiv6KIEgSm+EyMKTZk3WpEswdnAc7HDz3u6KI6Um50d6Iv5EnUY
WEHVeFwUbzukvu/nxVcg3Ps4si5536DhqgFlp7Duxt5WkTuLkXzepcN/R6HpGwoS5czgGMJ3G3cU
I33yzPfE+R2t4xs14Sk2Cbp1+XPm3T30dmGBi2Q1P17y/zseu7HNzhLC52oEopVc6+V6m/955TUN
8V9VD6Am8sMBsf+QOS+q0zi++pjY4EJ0UKzrRBkshNKXEMcTO2o5V4WbFQ+Kjhwl9ttMQdKnypZh
rnAWKclwtxACLpVZrLRhom9IuJ1JmIKJ2DD9iea9rootNIyMlVYD+1GnhZB2YSPuYSrN6OIdnd5E
F+qwiJ0Tf7wqJyCqGrQ/Gv5dlsSe0unlJHaN8g2fKGqx0Yjrp8VZ7kelrB1uqB/Xxm8K4u3mUMg2
UavoD4clZEzhhdkXJONUxx0eRokh/BJo/AurVgWa9jBBYYr1mQZ/uFom+in1oCryK8Z/d9sHLqFo
7cffoHRsDHJq1R179gc2xicpItG3/utrtRUSPq3Hv1rxAAerKTbDagBWFmVn67E5r3OLfidX/5qQ
QGQrLVws8eJfxYhj7mIbpgzph44TrsvjxW6ta2NjLMInCL4tR/lyYFeqib5pb9SOa7u2e6nPL20d
F5DfdjEtfRB78BVNibgk5WqShseyrDBYZCctNkZCJo7uWFeQSupPQcHBaLQIDefSXfFch/qmBux1
axMbVAFbjg5IOs7ebWKXzZOKg3uCWoHoKXP0Nkt4wpSJWNEO+xSc4pfqahAgaqkOD9oVdF5M3msv
TZ5J1EgQ+xAsIQf4kMUZfTCvfWXn2RNZW4moZ41W/CZ380qAAvU47E48fzjf1armaOFPOVWrT8r/
Aq0WNUCY1nJzOm5YjsXo6nknFdQGAZSB+Qa3lYN3jYttS/+y3OHOlaDBcPaFre0fsNgvj7d24hQv
fT8IJOPMeAU9JICnvndrUTuYkTpcrdQnIKay9YsbuOnMZp642vtfDZ/21nWX6h2xqh09lMOvnbj8
8SdnpDYVXdAaOX0xOq+QmY5PoyGSmD+Idfx2Gej7Fd/y81wDPSmN+u8H4iXq8pFNkh+i1bFjLAIA
+3N+oi8dTJ8yKDmvW1zBOJisTorsLokqQXimTtqTcIbdVxUmVAN9Vg87mQ6NjBzP9LggR/3qEVkX
gX9gqUfstzx4VURQiDNsKEOZ9mFF1R3oRWKIDmRpPZEhIIxN0M6W8WvdEt8WgKT/sNa+ARTKcSUW
N5TdB+7fVrHsrYZZ3z0niY4b3aN9RkDGpuYhCwJS9lDR2HdKf7NwqJKui1VQ61h0l2C7XuMsjqnA
nEVwQMJg4d1DBTTEHvCsuXR0b0A+lcfxNAIXt5qFDdul4uhvVT7xxKWw+2mgVzkGdHZoLxl3tglu
CSEHZbOJnM1dcSf2Mjz+d1C6kyGuQEs+biHB7eQf2gaC1yecpujmUNmAT07NKdZ0icBbTjgcMIkw
1jZAph29rphv3K+hdGQVsvxlx78Q8JCFRmxJbLcLNgtsi9LMRRpF0DyAtwKGGeunwxTfsAKmCKYM
7K67JsTkXDkVox+U4BTGCJrGoGzNyGONPKq2cYi6qWItB7yLyGezqCbQ0N5gdhOXSeGsGcGY0TfY
SXDVp3lG3XKwPr5l4RhvxAYpwhz+r6wvQbx1tBS0nT35uXJOXHdsXxBVxGlvI0uBttvvWnaN+PRP
EquKxYqxygrp31IOZfqOsqxyQS/XOR400EHX5+oTSy/y1aZbU27YS3s8ZMLcdsROx+ug/JK8dXFm
xWzXywTZt5wvNgsN0bgmhoNw5Y1o0+QiVSVl9RKdHIx+lE3W128Gwq6zG2WBrsRUOpuJ/oTL5gND
NU2xMWSIvtOc8hRoaNXGu7WxAzQeTMxERKGnNt9o5hxBLX+UYPBeCpwVv/y4/CQ0QcS/e64S2VUt
CqMGVgKBGJhfF3yA1leHYTWmO5PF5KsKkqw262YZPf02Ih3ON8y+BDTFxgAavYO9FpfX/GqTTPEF
Gbd0lX5KUjiPlkqEVBl6lL33+hEsnU0+YPEAJ5bkXwCEQeP/1g1LWjBl/bFE2zDBzIEiV0cljiId
iy08BAEjawsqiibI8GwDjrgnb/H8oOHs9wcid76qzii9tYv1ZjTBSXUxEQImPZstxdWdW+Jdjy4A
eTABZnb+qyTxCV25Uk9RnLqHKQXjiZn8bsj3RubcXO0kwpKxhLdxYetkAup4uMwCCAo4nN0OKaN3
xyALfyCQ4OBxyaQts2BLqBmYNFBQYpIizJhDp2FSW/40csI0YIleGnLjYjYjHhk5eMmSUi4T5Wv0
TlxhQMcLd5R5QVsBpfrlCJbaFeF+Pn1zGTh1SwHSh5GhdN1xjyG0wNtXXjI2oeakKPG0T17rafiI
eynF81A0WOagkL+bztQU9nidW4tAypG6HBXq6rA3FR2o6LeJRplb5PTo7cNHT9pbuJTqHiKBTdPH
4TlvJ/pwTtjjsrApDq12zQKGAp+5eZj3+Jb0KW9lfRS2LDiQ+/QEUGr7XoTWCeGllQTgcnjHGaES
zofPY1eFTVK12wQDqIqp/Uu6h8iD4DYduAwoRZIVcRAYhJwyU9/c+C6iv8Bw0b5DrkfknlAKeLi5
81P7FMCxK1KJDn6L3Gfqc6Pk2pHnMvSM4AJG++UNGl4lwBoBN4/JCy71+Za1ChzU/aujpZbjO47h
oo3XEzd4aSi2fMXNXfj8TuTkzdWKFn3t21BwTJZhGvHvb6cqQoVVha9yVFE4OUIHoTulTvB7AuEZ
EK4paQSd0wutq3A1om7C7kR4UlCJx7PX6DzMUcOaP4bo8RsrXSAQtaSlZ2uUfylJ7Dl7sZS5AbIX
xLrHZ6Qugb1WHzuZSwfu/q4nCLIosKdzB179MK56bv68MO4cBpFPdJN4LHgbvy5AWoV83+2SOjcu
dari4PIVQl32Mec5yUc6mjLBWJOEXB6EBf8YVPizkPp/kQYB8KH9p5Nd2mKY5qAApseLmX+l9FR+
sWaV+mbOnPwupSRvz/se6NAaUPvkxffLkqwTKRkLDOVDYOshJ9h3IJ4+fokLb7OZJXuyGICRVT4q
FX4tIa2ey6hAtKh8qlqmk72Qtuwk4FgfNgMLHY+1pJJ87FF100l5UhmrunapLjaCOlyghhWVVeJ2
naJQpCJopgXJvTwwWiswFp3zxvHOMcm+AcigThOxrzmYRvKrzTde2ejqt0heKcv4sd2sNLgMKbBD
aJqTPmQXi1IIQ4MbO4TjH0xgajsW7er+9ZKYHb0+3my/ic9tLPoWL5ppTsj/+gHZpUw6W/CJnwdL
aGR5Y5LHOk7LLBugcxcqq4AltklpyFpzgFII/M6e6x7Zt+auB1BCWW7bpnjU5eJxwg9MXlN5ozAB
qMMGeX0t3NNplIGiTpTUC04sMEsDqWPDZky7sMbVQ0W6tqUDooMoDQ4tCMkrPVF45UJCjm7SEuUy
5d6xpUOHP+F6YHzFZ7VnyaphdTXwzTftBS13ILsqWY8ohsYrEOayxdtsAcb31Ok7jeW/mHFcQTpK
ieA9sHML4qLfFeFpTcKT4eWiozfLaSaf8sZE76NI6JIz7Xy7205QksadS0upy1jt3mE8sOyPC7MX
zmR7vHgE7PkcoNv9rjiMB2Lkhj5vLsF/P179rd4k5bS9kZKI7C9DppliSI5yFH7JxDQy1ZrLh8Qe
FJ+3EjWIGHDl2o8A4zVgTe/a5LYR6o3tZ/5YbHs8voKaSvE4vbhneqYr57aBmMyiekX/H/S8Pd8J
5ieFmT/IxjFBs2xZyBcmeTd14KFUjDQm8BzE5nYZdPOH3wWrIG8XiCYwZrX9K8D3Yp6lkYznPI4Z
PUVaDzdNdn2IShaox6DBvqv8Eq1+4/lnnAqIItYmYIn4O9c1kZnCntuU2sLBaITU3aGxiQ2FXfGx
Q125uLUpvm3yK8nEhziOX8lVx3tsecJ80GmlXKVcnl9nC88ILnu1d2LIXLo52JiqGP3vKu+ejJWu
FHMTXsuZuq3s1enDaFHbtNnrDP0BJviTue+fLQp3jbmy6z1Yto/6h/wh7vjGBEKCx2Yp1b6YjXv8
0nKYeBW5SwHvtewZxQhMtpHKT5B9mhs5T7fybqyLnXY70Tl3feNEeL2+V/LZWSwXYnkik0jcovHI
cPZkMtQD9gtP8I2THUfsEsaQWE1x3cz0SQH3M69fNKajr91ypbdS/CtK8J7tlTyySPEoXH/5kFnZ
A1QCBysMgsrGCZLRlubyW1HS9prc8bxSG8JkokKwzWBJx8yueuayD9117POPczdaDQ9uqHJWK9IH
EvujbVc6VL205csm/ocHT49ItrQteOB+XHq7DU310PJmvlqrEf18eAkj5OAvIKbmJcO4fgb7VrCO
ibDCC8G+1liGIEcHW6ZsGjI8kRxtb2RLNhND9LQ1Dr1wSMKLpvs9YlW5kRfohByTTivysBGbvu47
bd0hpxAuJuBsNkWl2SB2ksEQFmWTtFt0sq/aiXiIR9mr3YywLwRaEHXi7nwFxon+adAVmKfgYPG7
jq6902F5+0T7x5lIll7HdDDDXnPOu7RYfq69DUwI8AjpPIP98zdZqGO02hPwPwtNyb2k0vin3Ofh
xLmdSSw189euwxZ+mdF3TZKhUhCRyKxfJ+Fe7UFWXu2EL5Iw3scwG2gR6E1vDioT/rEbwlhy8LrW
mTKjlQmd09azTHBd1NCWnKXvLS9n/5CfApGbnH7CGbtbUsTt9Lhw7/F0loHsU+2x8vjFJwa5Q4SO
0JH0wyThfao1XsqdhwXhVT3lT3/qkPZNDb3+FQNVu4y7LIQrCn5EcJoKaSWK4VbRLAhrNh4/gOi+
j8/bSE2IUjiYz2uzO4DYFVeuZFTsjPkFA8IDywtpHm7GeqVtkUeLB/v/K/TRZNEekDDf0YtTnZH3
tGItZsu9rau7KUka7PXEzkcnxxQl8itGS5hZooTTnQ2zJX3HlKILtXs05BZVdo+nCcE/+V0+a55D
hG6ntyh7JEw+u8nr1EZ23OqI12k0kCriGyvTHqzMosy2Pe8uCZG3LYEu384x3rHurJmSszC+HPL1
w8NGyC7rTfqROgp624VeGeNsgQhXPfW7kxWdy80RGPoC+MO8VnIi/QpHhfbssZvYjl25eHE9PfKE
+oPopT6FqINwPL2hzuXuACr2E6IZm5vlZD1iRdt27hTM83a+UH05k0Bf2ont4PblMaU0j2AL2kSe
oQVt37Zt2MtCFisuubjzC4KXpCoZKz0nu+8B2J8iFHSLU5jXb9j1CLoyNibo9aS2fAbN8A/w7h6L
2lnxQI8R0UfWqmETtis/9tf1SLIZ6dG4enYjrYQUmTyK9yryjTcQznM8YLj8xmwOh3Im77cvttGX
zgAuLBQtXdO1S2wXdh7snzKGzsQ+7tebtFzNhBoQC5WNWGtHce58RYKTRgz6pN/XAH2UlbHxiH1h
EtgyXUuxsTfDFeFHmWe8Wt733CbMGuqR9qWvMLMYTYPfZRE/80QDEQ8SR5UZCxvplqWIAuOhzh+c
61rQ46FlDHKAdoKw+TcCvA1lDvEtsMp6/r5mOBCqfN5liK0Q+nvNXB0UbHQN0YhgsU3b0pLmfLo3
qJJRytImbsBwdVSVzCv413pRVcc1s/i7qcv/npoMcwUXIev+uFTLX5qzUrYbE7LoOmz+7nOWGLmT
hR4UukE+Wam9VHIyQwu3OQtU86ZxCwT9C+ZIVTSb/dWismbvxzSKi0YbHqK50JIKLHm3Q45i6W8x
Q7x4o4BfMp5XrcpwJQK82G9ZbYKpK4uZML5xsFTQnHJRbgHzyaEtyE+ZBYvVGS8Ky40RKFU+sN8S
QIavnWE6PqXX+xkXOdJTDQd2efCNA9xcvKvlfyLn94PG6t0DiFpCdWqQyWmMYl9UY82GXxqpfkZO
ZJZm6Riq0E7/ZnsW37EJdsLQczybCXElfx7K9jmm8wDxPv15efH0YNLEmlMEaT+AOhF2/jdECH39
CEpZU8v0APmsQ2+cC7bc27KWOrwnOi4Htm6d9FAA58xGxXqWodVxQ9CxQem0x4f7wWxhT5eZ2K6P
NX2aFuzkLOTYOTyNlYNX2dPo7SqFVSd9ppTy70qB1cNjMJDqm4AtE+7BSU9LeO6zZp2EfckihAoR
HwWE11G9oBhe6cgDtpY3BhVunEq55MLCtCckcSY4dodx3SAYIUtC4bM4/wPkOIpdzeWvt1NHQlZm
fEHKH3k469Joz1tSL2y65TPE7tQ+cV2G00YmmRhSQr76T/0cECp8Wo3X0fT73APGvkAZtWv3/GI0
zzLjBVYMBy0BmQZbEO9bRYmrfu5dOjRrPa3KEtuVn1PFVI1EFBSRYtthMXArnVhOeAuxB/p499oR
dFp7aF5nSZyyPEAKtatBQjAxen6V48M9lVDEvxQL91FaUhAlmSaHyRRpGo3w/fOMZUgjGs84aP/r
pWDG743JRqpUUOoodesEZ5btH8Ad1hVAv3Ev3QCZx0hqVz7VrlcSpzNg2lu9115EfTtxRRtda2Ox
xKLTPORcYOCmMZAyU7lf2q7nCvSOP0SpvA50G3vEbsWOoG9oUvDW8ENxiDu35LhGUm4RjVK1VdP1
gYL3d2B+VsoQj1M6GLGgfZQjf24N4HwDf9/OtLuLUCMn06uGnbjnJhPwQu28Iz8DMSzFmKzeaoWz
1cFlKc+l9DpeACqTno1ZxUiyD1ynwlHLITBE3fK2388upwMuczvzWsv1ozcdGo/4ZPh/UOCvbJJG
h4rSWmoBxxxyJUYf/mJyA911eKrBlrJYjKk/zGg5/4YLILjGpUR6qZvPsyGNU1vDE9tjgjVTmVYt
0UYIGwKrDGiwCAgC0k2HxlhgV+qVTTMMfKMSAovFMp2OJGNmP5+rWLYLA9YlIJEKlOE54z+iDem0
kFNVehHu0euccKgHiLn44uk4/7I92mAw1EF+oN3DDFs8SSFP2ye2aw8mlmSzWmbEEi1PvwYddjR0
HDR0XQe8oUI4FDTvlqHit3EkhnUwzCVfAYmq2quQw0+pg1Nb5FiQUnPt+usNRq32UZCqFNnwbmH8
AU3iRLEcTVUymNzz5nUCANUoLMTW9RSI990dqhhys3D6FDWUgqJT1yE3fq4cRImvRHiuXunVOE6z
6F/9g1C3IQ6oqptmOeDhcTKjqbGhuWKvaGuRkcPzGNyjSpq77hx8lj319qKCiMq+5s44qzg/wbTZ
vBmyLzKTAaQTCizKTtG5fSTvXaBUAtL2xsLjyojvNcsPMwzYaShiQnGjnab6iaTdatZrHUrDpbHa
jIA/2b6w86iQg8X+f4CvELxTlTgWo0BmnbuP7B2meEz5yeya9HpPbs524yXKkMbJOi3QO5wfFOiO
J7hKR8GWATn365GlajtoWM2+nil/089kgkxZOkK8lTqbdLq7fADyO0L/8zs7bo/lB0/TyLUUZPGj
GoXw2eEPG4rzRq8YS//j+7zQOb4UQG+MQTqiJiirO+CRLJ/HlR0yVPGfhM4paljN16f1Ym7+nGTa
Wk7QPcqevbmF3xp3/Q9emdR1NCapnFRnjEcfTyjDkrJQET2ie1Jk60l8+nVnN4hsNZ4yr+MiLypO
XiN8/aPwsRuGJq6sGRKumtrH7zPVmJHHpNbnz1+mqm3Ixa38dR2k+xNU7qCoGhxtMIc7aw+Zcjwc
lxtZZ8slbdhNNPEuU1KcsjjuUL7ZpgY/PLSAXJt89VszpnrlayP2iuQbwDJkxw5pahooyZ+5/1i2
jX0Qkstdx6yBMDBI4Qu1WG8RBnDeIxkQQTqLR4KBooBREQU6ddKog43hmxDx6L3mNjGQP5jDPg85
W8tlBqCLMqI5MJKZrK5NI1UpBFYnJGXXuuVn5bhcgdjQwXJ1n2ztPP9muWlfUif/ZMBxBVALfkIM
ETmu5Er5Blwaspd5Eim8VSflq0flNd2aJIcAG7AN/ycK64XNGf7bx5hB3cNiMxRs8Opk+EJ8EVlt
N/b8tlOg5diTgNwyfFlIb87rJDv8/prdxPvXnjkM4Vbd+7AAwfWtOVGfQNXIYBpNEJpNOFoMdwop
eUIiONevgoYH/sFAjwUAiNzijJiRD9qQq8KS+7rhfPL8q4G3ZsQPBPBZJKEPFR528nsUlSW4zNJi
AIr2mlGUIVeQUOGdePJpkbv0xDtX3+xEc3/OJ0JED/JGFXhrrWe2dPLUNb465Owq17E5KM1a936Q
Tv3rY/Od7f1xq1XmaoPwAnDECY547ES2542Ez1H9DTL22iK9LtalJXGQFD8VHJEfS7TVsTHRple2
L9P+GEVWfd6oQWidDPdsOG3svmHaV7ep5Q0yaqxA0z61t4pOOQEgYKxfzTQAT3f7IDF5FZt+HhBH
xPaO0d8IAbXx1r9QT2+prnF8SyX2Dg4rM96huF60igvztQtteMX31i7V0YKYe/kd9dUoLYvwqmUw
mR71n9Wqp/21lp9WSd5kMSZXJ1TSd1fTK8B2rFYXPZCMl3YBlfnzj7stF/QvwCHk/+tuxltpFS8u
fMN75dWymj58UGEP5+n8/pw8Ugi31RoFraEC9GLc5Cwu2gPkJVUE5beuYHvIgYKFCTuyjyVY1dlq
eF1VbBSRsS86x4ZyGWOOh7MqjlK9N0rn6O5RCFUA+/MXTVxCjzwGhSD6XRpZ6fI9jxr+qAReRt9j
sCrey7RvU7lm5/zOkRsKdh2vEXLJR7NEsqPdziPLPa2JO+oyG5tf5HynBxNrveHV6rJzDIcp5inb
6E7mXCdXq/8Uoi++EVZglj6x0oXrYJtrZ6K8+5bc9aO0pifkpChxsaB+mOEyGaRR6v2IBRVtYK4c
Y7ZaWqAEyAODy5WOsIhLUWcekfhDVy31vAzLkGnCbADVdZiAOh+Fe0nwI7QYpfsV9kmtsIhBYu9T
1cN1z5TObC1jadElgOtPdtkMLDYPD+2IQtmsipOhMAONQoVrw+kn3EGHZB8vpnoYCmkcQ2vq3e+w
LBwSqe2XvTDMDj6hx2VrZrvEPu6B254UUBRURUjF5J93d76rvmrIKf+7uynPUl1dVoSwfm/YFs//
BhWDAAWrKSSOvpTSss+X3O9FOcd0tBhxSuboA8pBTtyee8WtqC27EOStxdxOqOCoQP04e0jWknxa
BdTE8/g8Izsv+7GAs1hdWMQDG8sYjRW2ud1HAK1W0WtBotlEJr/YrLC95L37b9hs9f6eyD1i4YCz
w4mXGghsZCWGaIsaqFKefBcpDS9ZDBQEvQAaefoQloymInl9hws8dyInE1yxfXLRws4kIH6nQWR8
vB791ZSIlxcxqVf/zgfXQ9KJ7Tw0U43D9Zv/pSc+5KEeu6NCDtbF7XPMpBhEHLZWAv1W8omHaGe7
7n/JHqsQCLLOozPMtaBaxrSbiAm598PziNMHDl2N/+8irqPPDX2vMv1EVYVoDWlRsuoMzTfNn+0n
Q/O83/EiLA7yN2P/d2r9xf2hPnmViNMCsj6dSnWT/PVgrQKjTtjCY2bNnFVzb2M0N2XHiZOCDOqf
3i9AWJf8wJr6Z9Dva6yyy2DtSGGb1RN9+c/Up+iaz5Q1SVFzRVe4MkweV+qufy9Cu2DdPh++TUel
fH2F1A2NOmUUGtv3jO7UtBK43yzs0MOTD+p9EsAaUooUiXyXCITpSOQtzfHhxuOx7iBmSQnw5wZA
byE0YjiFmSgDJlKOJNO4abb9g0SxJwFq4r3fiSk1+3CJANp+wJB91w/1gk7gBYHIAebwbjvqvgDi
EhQBvUmVn5rJoOZ07zrlAufKrVfkA4DkfErhi6K2SWLiqrkAnh48QTYcpRPyyZg/KORAQBIyqrOF
t3K1fEi1cJeTbJHpEDAqgeYsoW1HHDlZvfs5ZiYD//rKNOdbXIoQ4Uflvxs5b7WqbQhwvbkAV1os
KNJY5or7OV+h5ynqKkZm0Yjss5afzkmVs6bdCPKqrKf8co2o6+uaDZMbqcK9limJ81yLwVlAi1Vr
auq5OIuHrJ82d/5E2CycEYPdOnWXp0FcmKfZQhgxKKa416HNNJAJ8nU7JKkoeFOSpLl1VteTyLZf
h43QEgE9jALgkj8t4ADy0Kj7An1+NBVGuFX54GX9fNC9QGTvkqhDaOTQ15fHqVvBYjgAvhAgUOPF
3M15LIlk2kUV8oxw1Zp0P7qQcYlpUEuXyC5Cro48nKiZUR7UAqqaeq72NMKEd711fb3GmdpYJZUu
JRli7iJm3uTBMpnRK3kLT9KR9wLDDWBMi/L6Ix/W/mgkZokoKLCLxndL0ltXweOxJcK8M67RXMuk
21MePCVgnzo7uaM4VJHQ+X22dpekeuC31eO4099OgSEEEPH4YQTWk+dWd/uqaeOHph6XcwabTIk9
J2JA2sqinCJSr+dhecoVYgHashrcxV0MlxiZwG0xf6wtUxCeHgaN6GsddPNTaAFXPs2wHVKaaLMe
CaEQV2YpNS39oU4UXFan76NJWqrRK1EfB5hXPjkb4Z8XYwhldVD6nmdWpZE5ZjkvY452pPwi1JSZ
Tfwbd5hnJ7vmzpQwsUxOs3dt3IeptS68rOkAZvId15lNjFcu7k76uqW+dPs3XKqFqmugwceZVxQj
aEEzghwnCUb+Wvi9tR3ZXcpZcbQz5xRxAeHFGsUFqbdrUfLzjaWeb0C2dzG40OcXYpr2R5/Rn5TZ
1Lqfacaurzs8rrIyyVCT09AuLgcJCtFiU4ZL4vOmCGH3O+OB/tbgOGfdjypUS+aaL/qPWdSk4Y2l
uGZzl78TEB/E2+yMEOmKenMBFP1zQ04BSokhxCIQtsIb0SoE3yrWfePkBwu538EfsE6Kio4xhraw
ta0sNcsVZw2h2XdJ5UsQd5ETtxiUaylHi8XtxrJpFW8sqxgM4XUWuFasEZBt0FbbQUNBCSlta9p0
QMkZzwM1fPu2rrxKkaIoUdtz6J7DdBeoWOhCdC+DL47JcnGfzHzvfCKohoHU5UeaH3EAADx3xRh2
qS6HZLqsl0ACPobNXA+fJDH6lgBIEkAQ6J3s/plwBWrXmDHdgFVv5JdfEXP1Eq7gxtifhZ4HZ4Ta
9+raeOeIExDac6Ea2EfLR44XyZJNSyYn0rXKcGOq/ZQ9pqZuk/3K5sVBBLLI891+czurBP2uJM7X
GUBNqHdJa5TUZ50wHnFhixm2Gb3fB0c/0bzWVm6lTpZz+ZwdyY/WekVtr4XaPS+aQHM0p3F4QM2k
NjsYypPA8yu9qP0Ig04zlFwr0GBH2K7JlwmP4zNlIMYFKIm+YKzKD9WL8Ej+VHgtwEHCU1A6yN0T
z7LfEHMV+UeAiTCLgTvybhIE4o0jlKPunJZhbGf69aubxi3esDL4ZSf4FoHcMcX2md3PloH6g6AQ
ja07fJnHqB2UHKWjZxIU5SoUGiT2F6D8g/re37wuDe2O0IytVVT11V/KCL+3qgXmUg+TESYaWhWw
FtNm6LwaDbjMM/DIYrQ+/wI/kj5L8/Kt8NU1klpNMeRD3N871jVcWYkTgTyc6jUa786OFFCpgqzA
kO5JUMnW49pfIqq8Lqf79lEGrc9+kA1pt4293h663LUFw02N+4i/1SjU2r7R3FQlg+QfdwH9n06B
VwaJ8+ArFa8Lf5BYTlsS1BozcugKRQRRw+Fm5ibDDpsphpysXvnzoRZuE6J9I2HHO5Q4B2a2lJsd
vxovbtW+UyHFoRU7UmFBBXBkKSDwufHoTR//av+fUH5UtxLp15gEGYU7Nf/aQgAL3EYNmQrbAntc
FJhl22DjqwKWv914KYnWoCoufyXbu+R+7/6ouPvF6YifZ0g1eV/V8X+qD442Yl1RfXcuTYKt6PHv
8ENjqs82zCsY3WwNQrNyMV/7SPqn6Yd/bSe4Dy6gEulhnvRtM5lZzyrhM68Z8cj76GS4w/az2R4/
A+QhtmV2BxmePwlYWzzJ2O1ss99n/XZtpTC1lxL6eu13KcWzmm5K4CiUx/89VCh6J9IdlPPD5+Gr
qHpIq/sC3bPSwF7NRUz/TVCxsCCDGp1vmX0ww95rHS1pm9q/rAuGs4Pf0fBbPHJ7EfXJDvIDZXrW
cxxVXQ+68hQv04GNrWdnLRQtMWcM+XLDy7E8udC+DF54OkSxw6SnnJ4g+L4PQkU/dNw0U5Crad+/
Oufq2biPvIjnLgvg5W4TN7ufY3La6yzBDhpoFy29lqxuxtGz1YYUZxUrpI3aDUIpPY5o5N1IwYpH
4BiLa11f7/gSkRmM+zSvXfdyXdfXRoRVjvR3A/2+R+N5yu5SngGRykXMUTGKeJzsV0O3oxU98QTm
FlK56c4Hbbkh2Ld03UIys3idQCxSCdbJzm/dQgDsMcnuqyGZ0Pp7acY2vctt/bhgb6o8zPujrPXf
Pdkx008Wv3rY/DM3aTnzx8DytIpVEpEjCzFSU22RoL5PA72IwmlJ7SLwNJn+nfobOhdFFGMjBq8E
7Y3Y5AdCPO+kBHfo1e9Yc3CisoH7GbPbytulzfJb+NwXn6hiOCgdLaP6T4H1EOsL3Vs0Ykkp2IG8
7XHtVZPCkyqB+h9aNcbMOeQrtXvLWa67Ss1Zkx5uUoYidLULPcO8awXsXf0g2fx1AiMm2ohMXRtO
wP9H87WlyeJJglfvBaxkY/+kFIX3GVWyxOBlinSocbMZnOIrLqeIGdEYcXfZBxyDFXrFnWa0qI0s
jala0t61bG4mIQD7m24rcMiAJeuk+6BFq9sH91LCSHtoUU0xr2Id2pjimGq25ArOpRCg0k8elg2F
q48Ym5cVVplJoHP4jBVmU5H9d9P/gsVfX0BBeByZKDq0cBB3ipetK8HGOwKBtBrfKgotzRAJwWi8
zSgRpls4OXFfMe0faPpxC+MFKelRSC8OerwKOLcu3tK1/0LF0Ge+kn6tTnWooq2jhWFJO5ZqkIkL
e15c6bSNc9ymzTPT4Jino96D7L+IuIwXC1UPFAEvjufA1EHc752CYp25ISaPCac6YOWQZ2lTvbG5
SB08bo3e3dSU/ZnLdGrTDTMqsYFV53HWph2nlC0w9aSzB6L+5TUxCLMW+wNMSOE/0ZVdApYxYAYu
iC5OhahyPf4HjRDY9cPWGH1+IH1Z8SbChDjO9Ev45PzeyYPpGr4f3DJpCmakl+x5tb8diPFLbECD
HncFtXQmP9welTOzZpFVStuSG0WBoMuaacCvrNI9srRR6qjTHVg50qTCd9w9NMJId6vU3dS0OAyh
zdGHyEYV9LXpzoI1oMUPblZWn/4x2/ipJ5qk4v6W/51cP9jbXONX8GEuQ39P7GMmtrOXMm1Q6YjP
i+0qKI99Za0DR/who9aEud2WFDOzeXrc+KkIpdn3bFdveyOyVTtSp76umc0cGeIjwpJASwDSHj9V
rmd4uMBgj+ZuHZ43ShxNOBuFgFJqFt9RIwz7NBi0QwglDf5t87hco8n1mXER/U3OMlpxEPrXoUfa
l1tszNyx6g77xHpJVQxlf1vE2w+JFoAsdGzjrO8Rf5/ju+ds1grZP0NQyNtxyrBo+/7oVQuadhqX
jsOWgUWvuBFcCraQerhndsGY6Qs90lfjrSe6OgZIbpfJxz0jWX8xXuHc4GGo2hyvcT1VRNOcPXk1
kxUyAyqhbaSjsuJgeqJW+RDwAbWBXcozPFGZ9/A5S7yHpm2oymRPZgW2At+v8Aw6ap5s+S2AFpuY
vBc9Wr8ltsfcF2CvLlW2gfoEjKJ7v4kIFbHSVNud650Oa6LC2LdFe6gfiNbXnZBoTzQT2xjyLwGT
+eiiCspSmSQ1fwkfR95f9hR2Be9bv5LqssxlUWDP9bt1Yiut5f4FsW/Ree97clmwMzjIaCEBi2pJ
VVmCobxb/vfPwfn3xMaZSipww0lx2AAZ1kgmW9QSdsVgq+gJ4rLla8DOScISMd7vpI+2CupC+7tV
pi//eVQDEjaFJvry9+SdDdrEklEbCQZr1JC7tWUd+gIq0BwrfijGEDaXKNWspZnvbtdyXS3bOjq2
PDCB3eifs6Xi2PiM5a4Hz/F/Ve8YgUBNvU3SN5npVnC+MdeKbFi8g+HtenXKyLQE3IO9VKI/7TPI
kkAvJeXrRRYMNqav8ELXN8Um+Dh0xN0Dk+TFnZF15UbALqV3pdFD0O2qHEP45gD18Z/FDoogiwPG
tuFbt9diM4IgjhtzAY9zS4C3WRp+9iOSLY7Bo22iU9dvktEZ9hmI71GVSepf6iTLgOP7WgGGDC35
My3NZw3P7n4pV0MP5FNTztp8Lz7LQ1/AHQU5uWX7eKLOdNfDY/JIYrEuaGrMSr76cgaV1q9WQBDw
uBRbwTcm1o1izg+u803Ae4Iqqk5tZE6DhFNr14Leyuf5qtNx4gGssO/ZflqxhU+G0twaPDCtsGr0
3SKJSTqkrfbv4o4T75UGGmKXJ98KVFgNTfov1DVyFnjzBdOgLLtJCAidddndsG2zNUS6I+9iVx7u
BKM6QGkRsVj63aV1Louz4u/M5H68EZWvZBPeMi+dg9FbTj/GDM/Cz90eep/i/WJzTcXqjM84lbqI
RmDXv1EOpLu5O1ehcLZK4E3cS2iEdw83/uTWgEEGvwVwuKYTOztnAJj/acwNCivAtULZ9rT0m6sy
n1vnbZFUDythbEEYnO1Fcj6g6H2MN4JYdghSQG5ASiSo8bZd5hS9QDlTEw8++WDPIgVpt/LQsiLq
dMwpmPUesq6qQY/hi5gONzEZaqI/cvt8OvStRvNiru1WteV5KkZ6iZrpfKyyFzoJw6GPHOvIQufS
z1l2h86i+gvBCTDwXPgiUduERPOVizEw7KqmMKa3UQyLyIVlGnArCWKyt8kgvNhpUgMo9bxWhtsb
rj3ewWGMx1HNikz0/vWYPCcF560qCUfb3RRPu6PxkGr6FCPtIqLEXTtSq5HJYPuuuXUNLvnc5FDs
HU06tdTiJL2ToxJu4TjG8bSkUi7mBtOLny/ENUEpp7vE0tHadFG7VQgQnXku5R4G8s4QemiMEc53
OTWiKTatyeI6vfqRFAx2We3yKYzWd/VjPCQE5BvEJ2veZGf+KfQtTDd0hnDF3p7e55jo/l5V3MK+
8vKt58gIPWxsSpsDOr7wt/rrL0IoDO61r05gIXxjhcY9r/e78QM/NoS7fUj5OyCpyG72o2uBVhYa
WR/ZuDAaM4DyfYzCB9lg8xD920UCDgDA1IBdw7MtTmkgu9k22QRSMFwA/Yf2PHavL4sp1BLfqFI7
i+xHvANPYWwidwmtkn/zMeDTM4Q74yb9VUjRAGVRXttRezMOqUrjY6k8LAaXm4mte5E+Qy7nBNKt
YTJoQ5jf6mszewcXFYI/Cg1NfhMAJw/9ucg07Fto3De9CrEcYwmxiCrTIV0lKVuyH4jQ8dLz/Egw
pZWZ5sqqIUBC/aLJFYA+agu3D4gt8AToajJQ7+y9g0QnOb+rC45/z+s1M/s3HHI+bAFjBWEpa17d
lTa2Pw4urOWt1CVvRcwQ3OJhsUP6tEUZN4kJIrM1csjI87SQZQoFMxHAr6HHjPlKyoVfy0t8AJct
9xaySM6kbuCGZCyWHcpVA5tXFK77KMw90t0kHcvGThYNfSM89R+mFXrrq9Lew8c3phEkLjMb9Nq6
MO/Ud4iQm8FAonjo5e1L6kGdLmCmrJeuOjjVaFUtYfSmunBL1VZ4N5oksoHrv9gOYvFNar9GFMh+
pwIDPQFqxWssDHfl+YMnvPQ/KP/JeuouAYvC+aQVAETUUfK2Wmq8+Jh4kqXUDx8dbHt7rttc9U27
i9gk1vyCLg/DD4hHkqlQKEMYeli7HuY1LtjqIeVpkVaovu1N96kWQTH9bhws9gfi9V3bDvCQIxkr
Hh5+TfDFIsRHj3ragMyIimpxddx//UaqNmWvJ9MLMfxegoM6/aJiXazRAaiIk+fNgiBSXYSKrZJE
Or08+V8kUEA5RMs58Huj7nhM+d637AEC4bOcsxR+9DRAra0HYOtPMGMC3/4VpNMxGUmYrGmbPnku
X0QAHru3rVqy+946KZD+TYIOkBUidF2mUhAWfZiPTLqozsigo7/ieOs3ccbQBaQXhc1nrApTZW6q
81WwXNpCC6avozYW4svu9b6kto+V1g73XTLLMkhbnEG5JOebcFymzZPGHYlEZHneW2BRzGv62K8+
TaI974roveWkEKlb54Q1PJYwA2ux7FjXHeAkTtU8ca0nmYrrWiLIuD2VufsFkDtLwjk+OaQNtO7i
Q+dTHuuREVcVDod3Oxhq4lDvXC4IJ1pX6iod18VertXXnjUUDMyCGeutLtSO+X6XPurCSCzSJIjT
nA9R0cnxJaB7bxEmOkdXFimh9AzL1Avr7EGkIODS1MmEdkqtrCkIAlGifJZk8cBSS1dN+NXR/IgL
cW7o1EojfOjd7a5THIrhRlPVNxh0S/BZZvpcD8RblsJAKMNOFikuxpc1tpKOZk0JshLfB4Y/8BvR
kdsGmigdkcodRkKX923RHRftyQB+llPvYuW1vnR6xt/IT6Hz90/6qAln71vA9FbylHtHsnGAqbw6
pYJzlywUll6y4sv+aTCfwmb261MVGb1RGmmQi6TM5ddpV7NwQ8P8It/a9L7xV6Nny5d9zjk53J0p
o7aOf4oaStw81STFl72VpsA+aKJygFz/SG7SSWu0+bCNfKabCrjfrktaDe+DA0GvW5DGG3xK1FrP
Fh6J3jSmtxKG6CoOR3ZqIwyj+I00x1xVMl4JVvZ3I55dF21tRZGXE33o6CncBiyCwlnekal/YF4h
E8YsCIauR9lRdPlVFDlklDvWzJsBr/zQOhcqNUWijlYclw0j9KVr9xvoByyc9KTyOmB19mNG9zCy
RRSZzlbF0dIaJeoQSD4u9RvDRzPR+SQeJH+bk9U/t6mJ/EjM6gIfbfpJnW4VoRdGR5nf6hvv307C
CJooKLFuL1/nveT98J55eWxrA159uD/hn15U5uv4+pOdWbhd6H1MSrJKClJsoKqo8wxM6SkuM7I3
KFD3b6MC4fPXfrMK+cRigDULiTltgRxBNOfpiu0R4tmQSgtI6kcWg4+TGBDZ4MIEsf9lqG+ULDQj
jiXDCTUoQOAGYpaKSJgtrWY9cAW6J2r8ENiqR2w/XQ3ofAa6vouXhGyUBuP2HHvu25zbi72iuD8I
40e3eJgXBEpfLqTCWAzLeZEqv1w5lVztXy5j7dox4e4AfmVzfMlwWT9DspdyulwQZvLHPtmbfJjF
z6+Seoe0xasaN6WqyHVLwe1yoQRPFWghHoZ5WOeR1lpFCShy9Y9fLLcUH6Z7F26L4YCX3AuOS4nR
oFFa8kRF+709APBBQbNQNb43oPmPSCnodibRMOo1wwpOgaCNtGAG8GmwzD+Qam6IBNzYX7qrhkkj
jLQGcop/lg9EJVQ8lrfwboEy+7p+3WDvyTqu8uqs1HaaV5OuKR97CdlYLY2X4ZeDy4pcw8ohzL/j
IG51u5ojyGXthWFm7JKw6hoeVFzRk1rVa8u/AoQJmOiTrSb9dkynBhcevdRNMlNZ4mgjFs/luW4y
vkQEzqumbOfveMEvtN0qEEdzMA+2pzxxSt2mSRjAq8iNmx35+1oNydS2VepHvSWbOj/xy06bYxbR
8mpm0eJe8ZD+p9zMTx+gbN8fmXI5hl+aIAILIdAES+Eo4PSp+yCwYCiR1T9lUq2tyDVwPsrNJomH
hADrBEtbKvS4ZS/NWmScYy/TMtEUXqUARxEnFWdvIk0Ub1VKi11ZBYs5pAVJCwIL5EeaLsSMUvZf
M2HomXp6MqYzrhc3+TxOjBlVRRXxA2wE52o/Czj5rGMUJxYOwlTqX16GTSX44b71lv4nMWq+fItl
27o/aBCga8zYPr+YIEXqTlM6KuHnZRCVy9amaPjabyEQhx8bZ5WgVW+Kgg1xggM/LGqeNw/JG0AM
k7yBXREKNLI5+g1LTkfawN5hgL4dEzacj8dHXVJ/KJXDr44MP9jkgsLqCIxzUa2o4Q+4C9hyEykk
I1hGTtdXfEa1wZNWZEh8KM/hPDSj/19iOSHoOtjDwlscJtd5/y5zxHzEpAJbW6HIU9k7z/z1EOxt
sg2BvyTujC2laLAunWi+ieU5NVFv9FWzqLhgRrps5weEnP7Hb5IsH4pWLfBpc4s75uZsAXAiPflQ
D7bItYep7olFqqR+rFHNTNIx4R1Tnojv6vX7t5ESPltIBvKvhmDi/B4CZ6pS3gvNsRVVtIVF8jFB
nb/7VNlh/hZngAjCBhc5Std/mFgbGHhOtiqsHaseHJKhPcDVw1IwWRE4bhXMo/dBNRVi4zfcoV0i
0dekDX0G7xvV11FmOtZeVsPMlO3YcermC60/iihMpdw2ERV0Rvloabff8F0aBxll4tIkeItZsHSj
EZFzub82y1Na2mdjwxhQWFRWnMQ8drncl5BPmsNZoBbNEXDjiNvZRfEbEaokd3lQIX3HsunjTWcg
s052tDOQMkZMTX/eHZQU+JRXt/Ofb4o/+CO0euefp/4XwwSxLa8gRVzmVUxmlkH2FMalT3qHMT/2
t/BvGKSslaYxk3ggjxIiNUxo20QnAZQRARzIdxw4OBMtcvLUwZgrf89auQOQ4/diYtqz5qjtIeCz
Q74pW/tXuDpNgP6pBSyk1bxFSkhlBF3z1tU1wJNUjMPQOfY52/46w9nj0ocSSDLnpR8Fu5GfkztI
b4ZBRVKffkwgQQNKyQYA0u0fWB1pmUfpyHuIrYUnuQwYcfbM+urt2bbgHoiK3tB3kiAura/1NPhs
9A0qu9XuJYE/f46wZqwoMiOmWAs7QuxTkI7cfZYOPDBwXB+E+MvRTfUtiFz1mRjviZ4U2jH7v13L
owzWr/8pXg4ekWRgZT0EgkOa9L0jsL8r9fl6Aa00Z00EDPGhbNUUQ4CRi2O9J+WEKxzxm6L/FhO3
Gnwcj5PiNG0pjocItkPrVp6tjQv59npbRpztXMnwlj+rPGBB3mzgeCfip/Q9cmEs9M0NtKey3KmK
Pi0x6YJu5ua1E3fhxe+GIi2NxxPfa14r8/4ep/5sAtdg7/w3UBg00YCzrwJVryCPX24ikZzJnZSk
9WEUyIpQ4NCOJg4vHDV3W112SmGxhZlUr7Ul5RpkRzldFki8YAHx6ahT1kIchH6pPSu4AyRqKt25
NsNpOMfO7xsGIpGjp5VO4xx4M0kTQFUb7oE5+53KSzq8TASvYgHhDm91z9vcFKl347io0heTdFz+
+v0om8N9iTCrg0hOwliYYKCzMz4pRSzBWqFnzYxx3Mm4bAA0wgXxd9Zi3Pr+wfjUqCZ6mJOrP+zB
WtMKBTjU26t7XU+8bIVdetukyM9YtX6XzWrkJzEvDyaK+MVFOChWDyPFuZNTY1T7VpMKYPrJAWIa
tL+6iz0Iz5bnNW17QrKXPMKXKifuQu4Ogb5FEKSxBU9CoeZQO3WGH1/785dUubDvf/oC/Vl5GKVh
puCc1bCMEodxtpj/utayQCzVP60OWmqdf2DoipGdGeIomJp7ovvG9NReJWMsJ69uHcr6YXVgazr+
2wd6AMRZQIGenItMgFVHlyinC2YMSjmXT3aV9qJRJczfgcnnCHgk5wXflLUPtS+NE2xj/7qdiRy2
zVkkbFNzXBMy8ak0oz8lKkThcYCSDV+iWOLCd2UltRTQC8eezKirTVpegL4S96jBfhJGxcpy6OHl
+ED/xmS3DgxiG2ucmKhmekixXQTLkH0/loOBjlK6hCSk/4ABqMEgV7RBRQU/aJUxx8FVTZ3gf/Gc
8Nb38BzN4k+GL+lsGuGFjs5aEvo9hFruxrtGXql6ybmOLLXW8dkgPTa9mUeh9chBHRDjxwC0jsKe
WRhln4eUjg9nNzrEwFlkvrknzwK0ycLZbCwfgkMzCJ6Sd0rIaKdGf+kHgjSv/B+BUGRVD3eetose
hk00quHWtndQD/a/IaEKjwz4Ay+LzUWI9hJ5QJpDoSpm5utp+wl22P/70iWkbiobD257m/k94Bn0
zUu6+yPFHT0hCv8091Wj3Mvxh22M1NV3bPA9voRrt21+VDTrsNt5MnjqgAlbjZikjsA4Meds1mfs
KRE1TBLqWxmMzJG3VwsqlgK6J+zOTqLWTVJvjfY/H6DuAeQFsQXoewq41k9VKS8OnPfDorgDUBfY
JNhw1QXJZ+/UREyyvZaJ9bePAw/yHCTyU9aYsIAWC3SAdFp5LAo1icAswsW0T0ygpfNnwUqtH94q
pQaGTD3O79blGN3y6jffGFs5sAZrPxhmMqzqTGJN420IotvUHhyzdfubpMExb61+mLQe/5JUV0iN
6YxbF3MGxYZrvJj0NBWfXWdYBn5PV5cYRG0b8qDa+8b2xq/b4KdM7nEhzDKeG1IqkJi0b+xNdIJX
8p4FFJucTNV9WzvVgkv5CXf4o3nmlM5zVgP/5EcNv/Iu+JdBZIjC3SpaSLzbYN2EvGOIWttFV3bX
jR7W8MRgVYfPOaPidJXlzisJGyjEA6l1u3NjUb6gPTk0sOBQ02hS94fNRgFiJDQFirc+yit2+Jd2
ZWVge6WyiTAVrcAjLh5F5fyxC8UhksamBApGgQSMGPubimLBtnLTFfZeXSM/bThWTIK2OQBT0Uju
Z4GKQQxKGJmQjcJZvfi5HtCMSamCKvM1y9+iERNOdml0JnaS8bZ1uS5aBtx0t63HFQI0ZmDfa2V9
iz1p5tPOYVVX2KqbcxzoNjZMacpZndeRkHZ7J/5SZN8keLAgNLkmDFcaO4wCp2FLzta25TeRMA8M
MlYdwP4EunojQs785oO5nh6cDwsGxR5Wng243N/jSBmbrPfOGj0y4YqC28NK0bkLTAseJOfNsLlf
3wzUUHceLDANTzEwSQ6C3zdYfYbzBdPVXPWWScpfSO+asb5TQdWD6C++iOCG+nNzyk25xEtBoKZp
gVAJo1i27m+sVe3xrxtAwKP++BoXNiIXqea2DTtwo3IyWYnqH6FCOqjvVtNpHYBEMLMd7dBNWzIf
cvi54e4CsNKMZi8XbPF3qfngxmtjQfilO8z1V//4tGX3oobiHmVIaRP/wJKk2QZ5j6pYi900x+q7
YZE/fGyGxb/JD9KN8Y+BILyNf77PnU97/lwWDSGjxJh35C87m9HBF33xb9Omnhn8MVbAIyPTR5lt
sfS7sQonCO3yiC1VTOkDSZJ74NfI3GiqxDzf41CCVyeC7JKz2AYtCHjzenYZMbPG9kFyDZ+bvClo
XJwoq1Yw0ICQdGGXtid3oEXsU3a0WXgvT0/LDVYopiVZ4oxyZkR4FLsEb4gdUpVSCUZeTwwuNNJr
LGUZ5dA7YTt9+kDaHSXIjL4K7p9OHDx8wUEH31D1rqKy0RvFZjfCMoQCYCVlZj1ksWuqi/VzGfXc
youxRHm3N0jhO0IOXO2NUmW52NVJ+72fHo1ONpUFLfQ1NoV9M8T/trh7v1bKiuvMRHJrSr10LcAg
sia0FHtj1OqN8kQ8ElrV8G7Is/NNfCoegTCn9cKcsrfsKZlt5xCjoU3UAb72PF6vIWwv9M8PXmUI
UNo5RMof7nOS9wg1TM/LEiJwk6QlaX/awnpYdWE2OVeqwwE64ovisbfHEHv/zBrVSuiBbUduK/uP
WQ9HegN03/f4g/1zu96ixqYrjGX3b3zISh7p+6tWGgPz24FF/BaGDnOjWj7etEnzj9anouQ+lakb
2jHKaPi13c2+fktsQO3ZvVjETXtDHGgsqTRFU1HVgp0/a5tdtr2Y/YE+Lt97Do0DOhllAXGXk3Fa
banqwMmaXVe31B36DukxdwZAKFDPVGlbbN8QakV/2ki1SiCupQM8FoLCED9kd/VHLN6kOm+onD/a
FfwIhpUGf/7Ac0fq2+N8+V5Ioti5NrRfvELOcJX2UEnPVrPnM29Y17PB/IYJqx0CpcVcnBwpNg+f
VH1o/4vIJ6yM5/Z7SoO+2N/VUicM9irAjYK5/RkP1JzKs2hkcex8iMkjgXCFpG24ij4R89dyuyRB
elbVEUNYT62b4KUS1twECeQr7eVfnH5s/WNNtlf5K6a8oop/Rfy3Xcbz2NO8TjCgpeWLWw1LwV8m
xioHWcHI8CWu7/FGol21KMWGTY+ZW/+q0ujRJfpfZPvkJIUROLW3wuxZjCoRF3/yqwqP+KEogDEC
uAlRFnOFH801LCaaMzJM/4KtWQmyAgbV06mfhhF0Qc3HjEr6squullicEZ00uz1ajVDYdootYHwU
t8DGNnQ4w1/fLUNwyZW2KL2VRArVJQrZZyM3iubowO7AF8c3bevuahmFGTQXQvjjXN1k+CKjsvAP
lPjI4IuGmhTbKfWqobHhOhm6fx7E2sMCSos1g5ym62Gwhsmx3GL9/n0JWgP+3XMKt361d1vtOT7G
9OOS8LPqTak5xisY+qoE5qQ+1iZjvfCp9kY29LqAyzpYb/39CZZ6EobzFqVsBr/jbtY01fRlGRMJ
bFlJlPhfsRhHdH+bVzQzOpeaX4yzq+sU6wVSPJaDYbkzDtWO6qiqjNRuLfh9cSDLhv+Wtl7suRbm
5ME42UEFw82w+7S/HBKDNw6RCVKH8xioqchQnieTSnRZ7NMQVe/NZv7anBDXZHNSV7pJ2Mm7IeFq
RnhzCFqOOlGB3CrnptQHK2XFIPJdaWuH0fQmSzDEeEzYyN9+H3t/YXXaH03TbI6z4iU7fmZO9vBw
68OVQuXAZdQ/imEIvmd5f5LBn1UXl2Btdnr6ixtrnODSYc5GxuZnj6W4ZL2XlzrTL3lebXLZT8ZJ
uJWM5CiI73+eEN9yV0gk4m5rVoosvaKYtnJ/zudnAWDHyuqB8xw8c2zZAeORAcVv05Tfyf1xw/y+
FuxHg0gKdsi0ra8sphcEAwHry3oFdaK2+n7cI8i1q3phF4k+2iN0UmhQH5WAHNR+xpoxkrzSF8US
NXxG+5f8LIbVljU95Xe+zXeUH29z8aT9fRyBZnBgLoUaa+s56vQqAA19NLG4NYVec61cm8Xsp2aC
rQGiQa3rI0950ZVnDdBBQHEdDGaBRwugcS2tsBOQiPyU8Xje4EK5R0dGU62HcIu7QudcIqZ8U5Cl
M0kl8lj5n9fDoL+0bQInaidRcxbOFGwD66b+ERpykSEsL1XCuneTSbjRSHmdKiJfmgd281kQYvwZ
oRE7RzEZpd+nSgUvu0eBGm6avzJ5bgPG8s7OG+EPlDBTpEbV09JlB61kxyapOT3Z32KUUs4BQV2J
4lpsQJO6d+YWJDayOBibOuTowme9sUdcjV1rRd6bEAkP00a/KWRm6zepN8tBsBvgZW06KAKxD1xf
GwVNI4Faok8EBfgcndBv6KvMHcGo6sXOfo+Qo09W35UuI31DkdoVkciDF72Stv2FXMQIJQm3F2gJ
9CfUyxaYUBgf4zhAYbprAMYRytGS5FUz61qI++VhXROzbhucOLDBwFVYt4rtj8E4+MPiWPGPFEVp
QrY5hgoDRKzgnccNJjMv1s+LhAxL57cWwqRZLlNOIbjzfAvqjEIuec3fmB6MZp4yTfJNiMBEeInl
FxMCrPdwoypM/MNAf76d6QpYs0zDTaM4k+E4I8H3itY6eD3rQgV6gZLBdzEn4H4yfUZI8OVDpiIj
vlYunnfM5Wu1y0HSJfeMbylg0bCkaJgGEqnbYkve1S77Vvb/HcUFP/iIcHCVXVED1STflhblwgVc
x+an7OPd6+WEgIQnlfHPBmmVaeXdZqtBSurSu3dIMtIRCOMVjLktbObLrD8WLlhJ4biv3Av8aUSe
oWWfiL/xvEDlvbzLSr7nsMQPW6+bI6vKUVvNJ/E9AJcWb7LZrkMD3f2NV3t0iw7CszulMvRSWR12
nRbfNyZhva38gGMvPtSsSu/wU9RdNevveWf37AONh4gRm0zSwx9Eiro5cuBhy+NtudmfrkNUfN88
c+AIFgXf7yLiW8fSQLKa0yC5JFGOjwWJrFgRzDctXEq2yrd8PBvcjIogMRhf0wwnx7W78iNjf9u4
M+ZF3BbqTgl/DidEIBOkYGTJ0XRTZ9UgqyKHkgCsM/HK14U2WeHzJdqouEfPeC/b0YX5Ondzc6UI
a4hShu8nbOG+R31h86coV8iYIkM35yrwURtU2UEBLGDgnFwJmRcoeoBkv+z7PTy4eEMsMNKZiv1+
LRjsEC4RzIH6Yni4PjIpnCkY3/1K5TsMF8QRluvKkfjYeD+ZZO/zOQtvnLmoMdoUFwI/0ou0WJI8
nsKfye0xPdF55x01rzskDqHaNDk+Ao9gYcIWqAYnEjy54h2BPBbYHSdaXHtmsVDH1b4UZTomzh04
LKTYing0Vv54pnXkg5uU7tTIHv1o3fHzAU9tZ4rXb4IJb3vWWBGktSaGNdjdmHvjVTIhfR2xISSQ
FsdUg3VHjYz06kgSlUOECA6qaupacfOQXO4H7D5WqBue6XGc99wAvlers5Bt8Gx8iI1gmvgdt/nh
iQg7ZIFLpkM09op4VKhylHVkbPTWonoug5w1LW8rYSDnjNDrcQk8CIG6LIlaKGl83ZZdM2XpgIwW
bpXFDpwcgi/aiZt7+TuWaMGVdRlZsG4jez37DDQLeQhDW2AVcVxBYeTy5qU6GM51Z/Womk93gnwh
Dhz7dHp9LFmQHSdXmJUFJStVVUwIOL4oHndYHvj6sg9RBs0nNBxVx3u/sFHcl/tz3h5WBWbQin9U
XldmUaXkUfcOOmeJF64lffluCe6NzKFCZQWsVVe5SZBTQo+Erbddid9r1ffjzeXBsuCz0JIYMLPZ
eaCjvVwueu4t8xBP8G2Fg41PExgL6gx+knFc318xF/Bofh9RzCpE6iqaxculfSN1QewB+BTA8jGm
TbDzIwox3fkfo8OF5pSkPKb+SDOL5OGLzdGnw3WbH9L4QMz7Ds4wqzQmqvLTG7+yqd3XbGfjqUm9
8Z1pHHSiGcdiJHnJKd7ZEmD+jGSMrHtRPFt4qTDc2ArFCZiwwgdaeXK7qSLvbe7kgXhtcA3Tft3K
DwCXj0bL5/CNnIcUys8iAui8joxSNSgiUl2dDsmFOwKPcPUxjLq/h6CRDTnsgASwDPMNXlREPzgN
kqllghSrFtlhcjzXeMz0WKN0gDXfqV4rysGnU+E78zJTr6oFEVqbR5EDusFV19VO3v6Ct4NosZPo
rjhm3z25OaXWBYWx3R04q9C7nT99iW7ppt30WgkH0JwEABUXRri7/gzsOYUIEm4Vvgf02DmLwPbk
lw1EViqox8DGp7a/SByvTH69xw7CS1zXK4K7E37u7/vQ0TkO/vGVcjAwoZHjpVpDGQDKEQyz8gDU
r/5LwTkSnnIRvxm+dZ8JKgWQH+f80/XFNonGe9rbfkZCBEu7dbG/DFwL1KvTzydfUiC4ZevXNC5m
0LFo58q2afn9GCoUIlQVi40q3pYXBM54EcDdt4oQJwzbDvQDK4M43AO4Jz4nCqytMMivxRIiohyR
0DDqZ3IcL/B1W+zu6yIveIF3I+rr5YwZth6xg6C/q4FO9/zD82ZBRt53AiYQH4F1DTX8RSPTCYBH
Osr/eKUpRt7/22/a9B59CKN9jBX4HYUeZB42moXp/SWXmytaAaR1DkQPLWLRUK0QdeJMWuLZx1Mx
U8cjPT8c8YgwUVLMEOzKNQE1qWOULt2qeQX7trosuNvNbkcqL5EFT4Ueq7xKOSWffetNtzsfE7WY
hzG78X2rdfNXj9VkfS1alXHZfc1W54YIGjrv6qAn2VrtG58EEZohf8bK6SClP7QCNPtSmXC2fvQI
4MaCT40rm96PX6s+0c+g/O4MFKfzHfuLbI3LpUuDupe80O0Xg7W1SaxwZXCNaprWP7gVWP+xSiWT
gq+Pm2u+8MjheVTJzsbDnjRVVQ35bg191kC2IJJpZmlDLtUH41HuKbSlcJk6ubxAHJTCOXwZTZXc
BLyryGS8XR0zbwoy8WxFWJWl6FJJD+ZNRAqdcJ4xfsfN5DC8xT97O6Pe+3HOf0x4kVkJJ8mNQcbX
9MeMJXwZlyVTYUSg/BbMUwiQ5KaT3GWJtihi1qHeyUIHlQ27ktSbS2WZMCZiXs847TmHIvt+Wz+z
wBMsRL6Fdeq4M7s0M4QVYB4AXeZl0pdf8s1wfWKVV4UuMICLV4yq030Khv3UapcKm5KuOYdvMIcC
MDjCr+oqkNZ56jb8eQQbCDq7jTReqS6qhUm3QrDVl5x5dHsNjxG/OxbsY8y35ncKraJo6q2twxUM
R7YyFtDQaoNOa+wgQazpowmJyoE4Z7Dh5XmXck+JGlRXPYRUePW50WERDOkQrWGFkJ3qqC7olLN5
E609sJ7W+W2Irt+MuXCjSs1SsELNw2fGXcjomr2GJ6kOwniR6NJjvKPJORvAJeGV2igJseZHZ0V2
tq6MrPIi3DCNMKyehyV0vhzPKCUv2r2a4h2RizzfAJWG46sOTClEsXwdOdUZpluAic85kvPfr0c6
6P0qum/Jwb5w3OR1ghEJkp5c8BfuRfWZGRYmBwbzOLR5F7wqHyC740L6iOfSr4FuDpPzpbhp4YnU
/HkC+MO/E5T9aizv/WR7N399+5CLEEnOHO7m6pNk4aq77XvhgexkUJa19qi+8Brxk7ZmZbSPoPb+
+iVsp0tAjhjGWKI//XBh0Lhv2S9C0hBS3gvLqGwwDa9U0SJrN20qJHHDfW+tW9fUNJhxYEJo/QgV
x4sb36Wkw6i2amlujZB3n9Uu7hyoHWJnx/5WdlT3Y1D0J8BYMp7OoZCS/HJ+VYU5HdHMr94UlOTT
Z6kbMFyYnDSnN5YiiLZSgQr7X0behVpBbCcrGTD0MponCiwtvAyziqSrRKqh5MIwJuN02fghjDsG
4VoOxa6VPAPNU9OW8aH8OHZnNzjAoHp8X/3B4lwM6WZ8Nkghru5xp8M987EfNuc4QWpb5znrHuBP
r96gJJshDTfWKrDn62U/PkT5xEs/d5UpdKvUUPywHJiPgyIa9tLiht/3ASTJpIh7rOaoN794Uj6M
OsMd/+VIQTenHrPVAZAnx4aSEHZlRE0BHCdBLGKCSJPXLbPO8J1j9kWt3rPosuKhUPxAir4BH9jd
9xnOu3vRBR8lcTVV974fi/FfLOqJQWNSQz0/de+zUCIoR9b0omGz5ihYB9nhNO8BLu4toJS2moLT
hu31rKubboopg3xaZh4iHVpEtIECU19HvVfO0YUS8xxu1+3OHkYyrvl6uLJygFx7gT+kip4w2vPg
b+lBglpOVW7VwYpkqzK8Jc/SaAnIiDTTV6Z9FcqdLUbek6BV4DerwYGO/5mF4aIfGijYPwWt3bNu
hrvOfxOpZJXTeFRLgoPfoBZYErclWeuLytFWDt4ed9CFn0agUjbZV5FXnKp3fP06ao8A//dDOIq5
duI3S3LpBHLPUlLozsaymzZ1MP1l7B/9M6XgJ+qpyMIiLpqTv8xUy19Ya4dRp630eREeCna5bjSZ
8ZHZSx3XnYxDG+gD6zXUoDKs2mZw1fhcSMzQ9QgedjVtA77vo0PoqY3vwmRHb19dXMfyEiLcxC/7
lhT9tC+wHSiNEHAUnzOclPsrqEe67A4b1b/gjZokL3sjLj2Q4PmawW9Pv0AE+MdbS0yDy/Kqrg7y
gAIzgGhV5eM4TULee8KY/LZvgOmrSqik9jsjn3+gIP0HY9Kx8l4pP4kuIxJKL+Zlgr91ZYNhvdVy
LgcytvWTJCUQQ+1kwj+4msmZs6n6ca70qdT1R15fo7fSFlk5aLOgfOn4ggLdcj+oQrwWHBWPc6PJ
KlPMzIGLOnjOc0w2ykvUewp5qx/54WR0ng5PKCBKS3HMFqGoEbqc6rDQuNVpc3MmqPnMZc+9865c
1fJ34aKSRDeanpOZqiq1wd45fC+CJcoT1QiO2elmgUmYGbZJbf12/G12Eb9GLogZX3gjv/5Km2xx
q7qRZ2xRa9ApARW1l6+o42/Yv/xbufds2LJp8yoqKIIxOiLc8EutG2gtzvjdJ//0LaClb+49dzF9
MTtSa6sqNHeP58ueeLVPCDObhtKVqz2HBzpnPQ9o8nyLk/ZEuHXrHJ1oLVDbL20WAbeYBn4FXBPD
ElR+feWWd0rMowBuc5V4lTSs8W6k+Z6e7mUnADwYgMyMYZUikEv48jW7vcINcfPx3SOcAQphbKpS
s0BD/HHorXFwOCurulP8WLwJYksuyRR9SP2mojC8yoKFxHvWO/4rMwzbcwMakhZuIZiq3thpn2i0
W9ViWsH3bnh/T1HQR5TmSpUx5AupggOYqmfZXDS33HKpEOq/96meb+jXcoXp4C/AZfPA7q8COYu9
IJB7JxC/RhRobiHSlb5NIRr7iu/x6duTTceuhE6w+FjPN6m4rKZ65lakqoRaTqFnCK9fQA5lR4FJ
zPP83WOVatLUkIGduU8bOGzhbC2L8F06x3CQEgBVv64xWbdqroQnaY5aor+MjVzWMWx2z7pIPPOs
oke9Ax0lvKMiJGaeyOW+SQseq7BSBa9DgCR/KSvrKz/s1GKIggEVSUJAcIjn1b26bwNNxtNtOMOp
FgCaVX45l7bCsLfuDihc/MjeQvWVM9GLNYH9hASbxbItiqMFQpLvb0s6n8TzjEI12iZ8gck0BZEv
WchSoWblomG7Biiz0tOjpJtJ9AtJwaeJZLGfRtF+IwhHGeq7hwfkQ6A8azTo8wy4kAGYnuMNK23f
i3bL75qOlFjEh1n29Wkw3tbOqgZyr5DSIZPSRE1x58Kew03KmzCXLCpbbN9f96FOeNnBn5DFWBKS
xnkBKtr+CtPVtp+rEWjGE3uO6RASCXmUdCjB5xxdgMrZya/Wc59Do0k2do4I2t5iJeccHHfXZKvD
f1E3E9QqepEX12XV8CMYcU1wUBkVm92QP+zBConQib397pXyXjGkVAq1kl1gBp9c4fCEDDPhjumy
45SPit9JNI5kpthJQMj161qqMs4EI14c9UwvedmvYJgd/MGBX6pq6htJZl0UA5NvND01mrW3HRoY
PID2HvUMo8ihVvBVaEIqsHFcUEKH5p7bdK/q6JljguRFP33lnv6FS9HJJRU58VoKCNUjlrQX/803
kxTsET5hSK1vW1Qaws5qplcJzP+x3VJCSCONIkHLwbK8pBYdpRYkYUbt4X0lrE21j26gcpHaro/k
XDBeTMUDACmIDTilJvz5wvWMWUA4vgNZQnZJSc/u4PzQro8lAW0Evx7utJGXc/63h+zdSaRPYNZq
NgiDUVTM70oqL4cVmiiCHYa7ve7ZcOo1otrbjpRr095PY+4VM4ucB7izRDQWR65p7+5RmyXFPEMQ
ux7kyA4h3HrATcuFeuxj8HKuqYtcyGP/PCt9cRPTrbc8Qs+ZAm9jXkGSYgO+3oJzPzs7c5FCQZv2
25wF50s35sKXueEfpP4JQIKUgk4z0H0mbh6G2Y/RiXkUAEb8GRj0E8f2OytqHWZAQaRgw34IQB5T
i8UmTvia5ZwbPb2MVjlHFQYZKcWr9LrKYg+M/z3o01U2v4c9bi1YGIB67SnedhDUTa1sqSegXcOi
H3xHwPzKxZpocbocdNM32PvvKMFEc4NhJLeigdHi46XhNU+wU1sO7QBBZeGj+72ij+xhCcQTn+P+
hz1HYPVC5nMsaGR7gimZzBn/P6ejMzUUAjVcVcCxUF0yYTolCwcifM6jlToh5DZyf/vSCUBjlY6S
DEWbZyqSkQClv2bmbn/G4yeUjSniuO+qpcIbKN+Dr/rrHMWn9qHCMVVwtf8rNHIV1iULQAYjeiJW
59DiVMSZAywnTebC090gG94wE4zfIRZmQ9+iX4DJK4hT84BYLPduaSgG5DSezp8z+OLv7Ziqge5w
sjjof70RAY0X/CVLCe9fFgSd8TC0eFDVvmYF0EEKAGxkvymii4LtB5LQbXuBjsdRqxO0sTQ9mH1+
iiFn3lHBY+YDKFcp04x/NSB6gakqteV8cnWsP2e0I5Yy5DW85FGkRDhlaLAmldk9DyO6OC9XOR9Y
dbtj4rSmmN4mgUzmhmNFRXv9gczphZpuhwhVtapo7UZeZ5dtO7GalJt0ERkxliN0zbPIlM0kDoqH
bM3Y6TwXYGYkdTyLaWGa7qdxK7DM8TxrAQvToTozZofzuIH7OBDkRBycDhilvJPedlCVEoTlijQI
0N9ler2FYivDuB+PqHUigJvACYgAJmrkaSagFyihmdFJjcjP1IKUVUytJ9qrMAGmnUW9qEi75eY0
qcUJeeFc6PvRYwOcAELy/Xqx8HsXWaY6GEoa2uSx1K0k8NU6eq0z2Cbak58+FXw7nm91ZMhIiKR3
zLZE3QzuzryvzOEDnInZVUR/vy+uEaieHOxwg4tUcL6NcXPkYmWy6yNpSNSMOsak/Ui4pTJ6nbzZ
wKZouKWN2PJgEJnZsyrk/xayBSpTBBrtKX+OzelawA7gNnAjCvj48tcGouLzmahTSmuac3Dbvxdg
Ud7VH+wIgp30QN18Yal7ggEVv7YNWsF0mddS9Qgvs4lOhO0hWOnwXokzgVBk3KcaXUNcddn1xIhB
K4e7F6ofdgDFNyH4IVmWULjXNeB4EubtBVHwjQmIxZBtEyk8LvjrGwbtvGHre9NQeCzY8U4Ee6Xd
9UjqcK5BG2FrGlZ6xxohXrKQyQj1SnNKvV0YgBEKBo3mRK4aYxaLDV0Y+raASglebkXZF2VEpxEK
pJqphPuhq7bCU0p4AULY6VIuj2eg566JXf/I26yCOpohjUVCvCyCi1v5T1IDaQvOvoFubfi0Rcod
ebFQY7qw1xMGKBrs1Fz3enA8o6jrXL8sLlxkzjTbEaL/xXijOLZpQZjYOouWuwlnaxRavEC7+MrF
O3h7rcrw95iUHZZ+STrgLw61jE5egBNgcUtrfTpe/t3D1epxBCo3l2HKVYQNTyVJiAR3k7RcwbhR
k9UH6N6eaM0SlSBhRWZIRDhKNCOD0BpwonrRqwniLaEbfOhrTbaONEWH8iFZ/w3FavgFI9cRylKM
df8YbUt5FIrhQry/XHRneXhYq/uEHjkCZ5vz98QaZbUIiSS3LROPvDQkKztZfsXHxCmLu8Cmp8DM
CnlNfUaqiHishLZ5pKoCF+fboOnVY6nGXVvABU4y3dHNOt3TuegqUcqAGBJ6e32NDAndvbaww4Qk
VYn+HPGmt7AGT++SP7sCY7ij+9gGW43mtIcMZQoDG3XmvgLWDNkVN1c2+Mqbq+h1uNchXgJi7ang
chZerBi0CdV3HNiQ3vvLfL5uSxOMCVwQKQu02bqPBmQderhcTgmMXChaY3BGLGL6ms4tfY+NFhdk
2MoRaBXI8Pczs6VbVAOoPoX6+lF1OFD2Zu+FOwyMOyO7XU6sRPcvZFumHQ3KrkmewZAAOgVu1i8X
sgr12GHLm2wn0fZSjwq2+PaTM1RHqHtiezYJ2joJ9w6KR/Yr94N0QZ6PMahthKTEFfEIokHEPKmY
Q4NQVPi9sJjTFA1xbzyW7ofuZM8JJLxB2EnphIaP+qzrYGf6aCh4TjyH+NcqoEvgm7P3Jhlliabu
Y3kyhLmwud4ObH4EPXiRjBrZ6CRL6J5epGSpjCYJrmfv3bBbZs3uDwmCunYZXKTR343JMLi6a/Ag
t35vbFXwxWExofDYtt++8/8pRCPhCsynPYfTMELGenLXtsGtALS1K+fo80NogLYV+bftJWxjNQkE
3aXZ1AyLQjPZ1b0nrtYlhl3q3O1b5JTozFSyykpbsCTlAUmGW+moeJor69HMQV8PmyV9FgTes7ua
D5wKdf8J7aXyrvpSC75NdKK3w94w6aZ1INH61GWDcIxMI4tbLCoWJRASE4zcGvPVqVRqkBBiavKQ
322ELDnw3Otj7bPnBkMezhx2+a5YanZkzC7XzqKDm8xk872L8dLAIoBka7zBGdJCxtcX2qAujh0c
JMRHVzcARnfLYgH8n+q1BeVQ0c30ihbEUz7Eye1UTgAlayRG+gRokiQjECNGqT4DlGWQ5oEukLo3
Ere1R15UEFYJOvc9mXuE6YTRX4To8MlEQzp/gGnUwBmKTFerkQ6j81w0jOUNvS0S1PmN7Si+Agwl
xg27QSBkK1d8oBF43xsO0/ABdxI7Hk7Fks2w05tddXVqG9s2NcNAH+eKbYW7X4UkSrKG8VZ4hibY
fxz0U6byO8P/V/ksq3Nx9bTDrNeub0POlauV1uhdVzvrbarg1WEMQ6Oc9Tbig0lkUNflXZlsL5hZ
SrwKIOEUzpZEiptxqLC+7WWhyIsVONOTuHkxDip2tA3zHyrK7xP/wkD14kzDYkITH0hxoSLH7xyC
hOa9182KnpzcQyWlbI95A8ncgiXSHhpNMgkvEW7eU3AkIyhGZKYo/2q/g7d4gPDwQGrZZA/f81zL
aMTGIEFu4SJatmsrkWJ6NH5xpTXyu6/hSw9Dpi7aeOaBrrtyc+m7jEhy64ZwFBdson9JR5o9/kx1
UbhRVYVJVQjMw70R6BpwzUKedTilnxjJH5sa+V/xz5G3QdAP/ycXGbaU94i4mwqXbD550521hA/M
6UCv1lH7miueXJgt9ee1+fABYp8xfCB+zVmvmZPTQKY1mSH+4LQBp8oOTYMdWeNB1hyVZfdPCW1K
J42fjeH9OLqnH5RcuxjJUNMo9v5yGARlO386Uae28K0DIb5R1MJ7xQE0d2ZAgLcNh0YOanVk2IPW
/jyZ2KqdGhZhmV9dgdGCObna1XxQEmNVqLAAnFLXmkbU0OCToOM4TCf7NxMf7ikVOh1lQ/PibwRn
T/COc2SvllLe625MKUIAomgt4+k/QWivmgySfq/xz7Oq4X4j8X8T08UuaZHtBD6/VQGHaA+ptfq1
0fD4YxO2szjmRWnJyIZozyyPlkFUyf9mChFCTuDpBsnner5isvtYI2uNIwLMEgvCwHmy/7tRMAAD
ataQW/GL768CUB8UI9Cau+RMLalLWbGfnsClgRtylVBFPo6r92dGYgt3aQmkGqlg9S2OroDZVjBN
2JQ7dkitLPipadPTkfOoGgNaQemysLUAgfWM6rl1HlhDL8QVN7Kf9e/Ow99gyyd9C/K67iWy/2g/
D54ejEdS8TtqCUYNXJpp6vymBpuBRENN/IKjm5zmaRSnU6rnPOuec83542ymEBUml4tCojjuMK9l
nZxfmRBLtKo+SHTIExPYZHFlBeiaf65UcinVP1ZVuXMTetwDzDKoYD6KaT9FxlbziYSmAmPKvwyO
lTShCP5hu+3ZZiJkARhNRuiEj2c8pq2dhd6wigPTCBxDphylRTLt+vMoNp/cRbpdh9vXdW4KSiG9
UpiUSWL6lQt30PZ9gEKYhfs7+ajlj8ilK5bhMKniDsa2EPbp+/tCyJftDYIt+PkLs7Ph4VguSKNS
QVjT5ROJ9VFae0fLbDsP/oNdjdOv03f1X3BRBqt+Ce0jeQwZ6cLjZcs9XnmFcoWRDZP36yVqTVok
Nr2zFrudDqB8PvIbx3NGIZbTTVNCXXfV5+4SLgGTDmP4fb5O9WAGLQYS8N2g782qEJH30U++Gdif
mAP89Ew4uB5HL83RXTXW11Zyb1UNPpC3eOcO1hxkqfNqNECoRJ+JPu0BsRxHdicVZwuGOcttD+Wz
nt0Z6/pxp9nRd1E7gZ9ICX7Gri81+VWHqF42KSRG1q2yP2oNB0IaxvA5iKhzLQWpRmboBF2zUEJA
D873zuT7SWJfpG+S7mIYm72Z4uUmmiLChGBLpeAjY+zngvwMhDgiLIP6XiliGRHZH6X4Fu0+5pMO
jv22rEpesAxZpChQAKBRP+I0AS82ucAW2r23Qur947OimT2JjAOgt9BqCXscjZ1kG1+n4QmbNAqW
NVEUwFh8aJuw7XEqWZy/lJFtbEwZhv7DgFXLNFTmKXxv6q4qJ4dmu37QyaKJzb+DhUMZsTgJa6as
FXxDrAgUAsIxRR043gYcr/fnfUjIVtAZerXFEW6Hx7WJlpPO+dmtvir5oifIyoxAU4cKBmWuE1MF
l/a4HW2nOLNwU2iMn624BWuHwdhXyhg3zUAbyUKxGijTO8/wUdhWyKYQHNQHf6CHi+WmGJZxNgQM
pop/LsAe24CrIGBsdfeBcscMFQVakrentjlHQu1akOgzHLAMFxXxWF2XI7s66JdfB+h/D4O96GkT
FBof1jWCpNAazalxDV3xDWWqTXbPIPNhbYWvbRllWadsylFstBbb+qAUETAKTge4SrfIXup6VG90
bLn45nRINlomZtNiNGnBVDuXViJpvwDwi75lrJi6JWtX0ERec8OJG8zkbo3An0snmOxW+SVe8Ttl
oUNmfKKwjTRytXepWFiuaL7nEHgtisSVGLvUot4TwNIwLOA46X2BiAen12+B9sBJPS0sip4SkupN
sLN5+QUY/jjfkTqRj9dhxLnxZgbEEH52UBG6QlBjf3WjJCxycmsmGOJNREudJ2T+3w0E3ofNgFsU
qhcCEhBJIU+YfojkoQRVOXTM4zGvcyWTTfqy8ZaGFbCBruNAt8fsCr5Un5NSKeLdTmhAfHwRTTp9
imi/Pvh4bcEYA6sNSpwwD7FOrhb+idmYledqqVRIjQGDmEBFNpzEuHPU5gEJOIfMzUOerngdY1Xa
K6axZJ4Xt/XftjhsvtXG/j3PJgh3969QL+R7B+xEu2WSeG9poMViSdUMCCBy1z4kcTpxIsGU93z6
SE4OZJJT7NqGJS1RqRBMZTiUTv2xROqtLkMGZULVJWJMhbU8Z3trGB67e+GORAhdeqk1zj4mhLBd
By0+/8Z2uFw0p/8aDSvcXZt1F1IMTNv63NU11Wi/gaqc0GqQNmKhED23Iqn8AV9jCwQqGlEFQE4o
IxBnyNS5s1IG0B81LUoH605e3cr/5ahVjaF1aMXEsmy23feuJrfl3XFBnzDMLvBJkaCFDBlHexCI
MvOtKSxjfpCB4YSP0HfJTwzQJTD/amgizmBic0aN0s9hNidhC6NntLiR1MxNj+uFMwMliK+5OEfh
xuoBV616CGcezhEL2kn5+Lc/xa6C53eNkooMGkieROZZCUX1vfAAPP17JB9FpOrHXtH1p5bxbUTR
3lYs9v2iaNkId6gcJTGGFOnxlWXBuBiRCjMV1x9dXlGF7xLhA7jWj3WFqLgNEPnmY5jyg1l5H5oI
5PSapKA+hxB0SAAl7FZWGg6lcnIjVYKcY244buKlcXIfq+4t9Sej2SvyZ50YjilPLjb2b41FidG3
7FmCYxnrR+kPvU6BL7dqDvhFSfGyyUmJCv1Ib89eTHOZhSZ4Ks7Y7Na6spJo/ahRHpmiXuF+fFEC
BFKQbr6DVfavsLk8YjlnL1cZp372oMgv/WYVQKRC3dNLZnakvVmmuN18eR1XxKpRV4klXVCYaTeE
VXJowM9dk6BTU91BybrvqJ2hJ39j9qK/FJwJkA8bdoKtlS1JzsUNZV3xpv6mG5L7taMfRt0HXqBH
jxipgkIGbJxn2TwMlIn3XF9elFYTmM+B54nMc+/5PSYZctieimBrzc2I4H7Ummw39sMpLPgVd2xc
Pv/YZFpqy0vNlErVYjgocEV+0nY6y27phMDUdlbwqN4YR0firgHnQRiwBVwXl27Rp0+nsZbMWRtR
g7iDwLTtv69GK8357+hHP2B0eGSQkFEF9ZGIwRXYQMjEBxUqbEW2keyZWZqvpks79UGHqMuGmIxA
iMwleJr611Vk2VN62y3z4U3PmGrsNLS9JdzKacNM6mYEZKksiPhhduGU+84Z/XcbROQ1SjJ3JQLC
UTm2i8wnG8fpbiTG34qCcbgXyqj+g2dP9a9lfZRfXc7mV5OWhkz8wdMSv5ZXAZnDyRQLDpr0M7Kx
89XQ/f3JVsaj8/NQZLF8GNJeLpciwMOn9fmnrr+N9+626A8ulB5KPSVYtw3IuKCTtpoesAjDYl9s
KC62L1hGojdbNWxYAvuXmyLa9YdEfXdIPUGeshdR0h4cLtX81I7O1c9f3hplaYdGPh8E+BgB4Jej
NcUzp5BOeftGQ+8rQqEsBbHNf/RbHG40x0HFzptwXe0aRsiDTdj/yuazQJngADKi1Poq6fEmL/nm
hsj+XBPqeoD8TfyOPWmFpPYJyVKnFzPzUVtuc+Z0QJDKsqKfIb/To+HMBPDm3h/Msv+WlI9TpFsG
HQIfBMr4AQNfPIyo+yqmM7ZWxBE9b/DnqWYik3bIRLcHm8AF23AZSwXQk2R9v9yPQvDznJ3fTJJi
zLymVw5KNBeMz/d80zcXJnhZi7Ze8Dj0zMYnafRZHYh2vfVzFVki4RHbIoBe1O6bwiYdL+O+ntGX
7x98B9jGYPsZC601C1ye6k8iBYMnMx5Mf/Ig5qan2MY8uC1cJ49qttYSV1Tpc1YgSxeCWpT/ibSq
tJRr0+0QXYNlEAe+Ru/EfUDYE4QJsApEuiS96ylCeVaqFLyAFiof9peLfCosXI3URkTKKkNGY16r
9Aw1oRrYpA7i4ptwQFW2OX1HGyxaRX6Cf+YOx/sA1cO+JbskYMrHcMSJzFSE50sbkRvhYEBJGYAx
S2rVVzIWzboVIfJMyfMJBsZfsJguvdsTcB24cYPD9F8Ntqm8lHIqby01uYgSygOdb7E6HuQ7d3VA
ChxLyawJiYE4+Gaym828JBAabCIpCFG3Q96RXOaWdiDPdRiogeI8a6Ar8WHaAFJDUYU3wOoNQaXh
RklgLO1kJEbvPn7fp5dO7cds0rdB6s4EBIzkhXIcZQ2rB0SjQhtKL+DLD0YEvEHkid9K8bxtCPwa
htTc7874IIWZTYcp1F1eg5SbrJZ3IDZMoTU1Ox5a4tA0OZmH7f2l+G3U8ztIzWnFZTMHb1kuhRZS
uXKpiRnIs+1NtVmX6grq3GGmJQaXWfxCNhNuaePaQNjtTpUKFLrHuv5BJzoD4dIlWiSQ6KUsJ/kU
x68pjcvnMtcP7Odpm3nyn9HTbfT0Hl09O9bpwSWAbYaKJpGnsLkN948O3x4MASjbJO0zvqvO3EMi
iQJ4gTC8HJ/QDiZK5l4f1l3lVB+x8yeUxiIm0BCHp1uqhCNdAimo15Jz8u2LoqGEYX6pTJvs7gmY
C1Zocb+AHYqTHlAKANKXYN2gbFBf8M11CFLFVTxkqmelT5ai+nOftbQCBKMJeV8AZG4rYxpeEN9Z
UQ48uZ9R7Wv/rQu2o0isqfXd1/+ZWL5SqgRLctwt3ykQaM9ECTsaIdFyPFmh/87rCIaKVwcTxqBe
icKDgp7fl2b4E1fmDXaRLx/B/DW60AgYWwJlbncIGU3HtOvP40ShkZy9NVwHyeq4EzUGxf2ziDai
TU+ajLFu1DHfGOEkAxOhZUP7sL4nmtHVa4AUZAUSFMiD1FosCfSEI5gUEkNfG0DZx0v6Ai+jhcCB
J6w5BLaAKbAkM6SfLld72cyNeT9kZS7/oXboL4qQ2UrUPlu618SgbA5sJfBno/axE5SYy3GMuCdu
FZOGdBPtQerFeZ6OA6E1xS3IyHCA2CJ4EsmXHiUMyLCqOy40Q3Z71jeRalQqB643fXUjEYo1Yq5z
nqCDNGqoV3fkRBs2u38ZQYZ6QNAOAZ4Ci3Ejbqlyxoekoc9lWutyyBpk9uCGvIpqkjKgBwaDMuMm
NnwhqCM7V4Jyv8X71pAU6zyo3uvf4gQvvBDTvXpSv78XZpVVyD+omtNS1i0hv26W9ViSFn5gFxHP
ekamR3+ry2gQ5oQtFpq295LA4XJBwaP5DC54pXYNajoHw8pHv262eY4rfeCMq+gw3HGcGh3Vv6GV
jHL82+m0N4DVsrXj9oKVosijfqZHYMa682Dj7u4SVHVfQmi09Zj0VO/inEDVfXHVBdwtmfm/5Z5C
9X1i+TDoIFYHLMy14XdRx0IWHbzlUlt91wY9tmyH22XMd2OUu/R74T+EO7PKw6vlOXXp6gzf7Ae3
/93zYe2dBBLkg/sLprr/TbF/CrD8gTFrbJRh8w1tbXJjTdeEtCt066ozzYwjgXuI2U+JfqRg+t+R
c1viuf+9mU9fZmJJUWZvOWnFE6IePC0J0XTgnoer98Bx2k582F7OftE3R9S154dmSyUF5Id8UuG1
wmjNj/YQDdrAynu+gBNgH1qqImbNg6x3xxmjN5rrcoy69bAByLY2R7WEjNseGwJ4M+BvTMXOAoev
66KH0+epq82QGPA8yDUny6qOraXVZkSi+OF6/BSb+nufPkjunYsktD6rizvYlhmavgdFHEoqZfbT
Kt2byXl6Jw1pGRivvhCmfJbJPz2am4komDsCuyDjHE7LGMow68ZhWuktqlSth4CfQ8mtkG6yURIW
UrBWoglp+K+9XXRqUXo/6beQudbarwjl8bP2Q7FR8Z0hxodcpz+8gKWyVSAUJqHjxY/IEGW+04OO
wsmLXPOvje4LjHcXHLPBRUws/oXodhGBUuPD+4HwVuawXqebAcmxP/sGOP/k8IIWaRsvm2fyDEOL
7bDwKFYJr/nJkuHyBXSBTaLAT6hhoirtkvyG5ZP3QvmDCy6plIIifxWl98t/B0lAup6C/3TCYZdA
v8Qhpgd5n+/vNZ0UIg1Q8RMwK0kSUETDsVX+lF7rPUVIdNIJjl/bu8YfgDwg5fruQhVLIOygdboZ
dm7qFwBq08W69T4sTECIIKFk0IWn7m4fyHXtgfPRGngf4O7/WS7wlNEPdWW7oGiBMUeqDkhEc/HU
41lUBHmYU6qtCXd/NawgYJPNZqCjEEI/js/PWteNjCjDXuHhly40i1gqnhPDoO7fAvIIrAmuIRiV
v3BjRK13DGxo8lAm5+oPFG68qLagtdG3XLV0FKUQdwrKBuVB9NAjcQKJgXuug4+Wl1lb7hqpX+tK
QxdrL4ZmweWFTR/50MD3JKKptqaK4KZGDiuXb7HKM7jDbLcchts5ZQ09pVNDjBUoqKpDz8X+qaOC
z54SrLD3B+E7vzA9i+G8/ZGVzCIIOKu/utZ8lGIzmoDdPCRqTaJyn4fFqu0EFWJBjvTEvdeKtj3C
3x773SljCdfkJiB3Z4GxHdLT9Ahfwiw+uOYV3tW82gjaKJG2i9TgM4RfBWEEQfcXo8LE3cR0hmNe
i5WuAMdSClwOAxRtZMDXWYpB9GRFW8no8GW4qeyUdGhDk+0L4tHFGewr23lGA4KVLMMFpmY4WnC6
7G1yNya4Bmv9xNMPHSpVzk/z5+9IMPFzfZu/2pUbWUvqeLN3mIW0SPD7wPIMo5qw7KzQJIlrUU3j
yJopX6W7TO5WJfIPfe9lxvG1HfanePN0QwcDKM/sK8odyF8EbWIvoTOdXFENxjHrTObVx0FaZbsE
BOcyO24dED6y8ElS/UoZla8IRd6XLJ7EUgFaNKNEzaS+5VVjMEXRLq2PwKanfFh2SLXwapqth+Ye
5nHthZd5PFQYOL8FY7/7+B0T4OIogdI4qjP0cTiIFg4tW3m3kndYPKgACIo5Z5JsK1kh1LJglMkC
7xGUCqizOWJsj70IPw/4oDxaC1ZOBWF1SQkS23Hxuybt0MSkwizulk0lvUxZsZjOm4tuNfLJHx+N
8B2TcZgdeb1yH1Gw1Qdvi3wwBTh7FCUWONtx+rASB81+zRkC8sbcyfce6a6HNsGWk57hmvd7UOR7
rEuyCChu0+Rc6m025jwbgY29PvUuGQKJUy1wnzOxQHSiVpZaW65kVppXERHJONQcTvswPCBbqkW7
/yKoRkEd9oU8wd2yZhNDAixqoyQfnbCjomfUXtiK99uazFsSuztQMLkfcoZjh+6bHBjwEb4gIx/2
B49eHpN1vMRgif3UrbFCH8JYpgPabE5rMU7v1zzryqi+6IeGL0Gois1gu+bP/+SMBfecwpp9SZbL
AQqbWjfRjP84Rj3kGSy8dTWaCjBf6U+40YpeOPtjhjfUve6aoQ6E2cVjCuMAKygPxi3Ilo6aJyIK
sdJfT7wkXzLTtHrtHBn2XAHLp9N5bov8UQtbCN2PiuYcrg5dAprZQ6bskbhetLXBS2kR51kmlGoo
j8DWggunIqqTe0rW0gdztwuC/nWBLkvWZvL5Daw+RIar4xnMvF4tv0XO+B6U7eDMAGdcAhj38pbL
M/3xP/yv4aEkP9LBEkmlgm+8vC2DFzvdRgjtJfOs2H25xjuqMYO40HlHPYW48knbvdDOSCODNARJ
KItyZGzYCFR14cdmMZ/avdOQm5nCgb6kYnR2Ph9yoYNOQrsJCbGW5ICv18Ka32IE8chW2bW9axsv
b0riakdT7kSAgrUCkGJh6M/oxoapYPJQNP0mkIPYS/NFST4/AsSYtODu6j0HlSHdkL2vhKRAqTqY
ZsTPp295Vk7ROgbz+h3p/L8fwZiT5myYkWiFrEs20+t4ZDqXEhkURnmlSd5aAFUshdwg1WO+WkzO
xNlABTmg8vMTzMgub7ePmWmsJRj1uT8X9K4B1b2x7ezhie21pjjy9WEJNalG/Xo65+KFaSKSia6a
jUSLxICObt8maWM6LVyJkp2+/J8fK36bRPk1RnbCR50Y6zF/3nZbAKGma14hfPmS26e2dXOuN4AJ
gyu7pkzk4Ws/ZNVRplFrwz/9SWpTr4OZ2C3s0Zw7CJnQw3KqShVxgPmOsIPwY+43U9KsiCZHakmk
DqRCno1aSwMkJcr5XLwL2ZiFA5GujsUAqyex3V/Uu1Ey+7dTSre+YVD/h17eQ/i3shMQdB87ddYp
tP64KOZ+2mYFOmG6hSfYu6d1zulyuATnZyNFqXBS1ke+L6eF+k/LCX2psL5w5xCFPE9vdg96N/On
Pr/Px/mppPeEIG1p44HrIFRhkhfHp/xOTEX2alXQPo0awrakpCG7ZIdv1K1B3IBfzPHnaAiSaRWy
x2QLJIlRcSuoRkc08F87FLGY3dLCuetXhw7aL6aeIaXf0PCsOSYuFrOXU+ZzXp+7fM+O8hU0/efh
WpGUPs80CRLz69m1c/+bfBK3eRZYWOCZ+KkBfK2rgHJCUOttuwUNZDN5myT2J12zVGAXafYO9PAZ
QXho1mP7DarK7NpZWlFQTNbYQETuWOvhaLE1UZF6/W5uoU+xhpiqIoJIEsWXLEdG1sGGtIbz0a3C
LWXK0fR3lxm0o95Vg6gehBLyYcMP2X0CBsUqDNAc7BXhp14udD94cOF/KNAK6sp36GB4c/nFd4OK
ipI3U4dWpAFAp6DZs4hRgal9LCqCIo5og8w4cWoX+gxy6+Z24ULP8pBsBvYVWFCWLuaDmX3CwBNh
KXtSYYh3ereqFdKM4ArN2K2BV2kK8e3twO/s9HEUo83BG+217JVtiTkyIAevqFAnDLCcC36xJunJ
Ocy/AIRU6z+4K0kCKTk0GRgCwqAjzLP3OrnB9XiRV8uXfM/5YGxZBspHz/K79X0rjgb0m7pYe0sq
aZru4gmUtGRRNGCa2UBRVHDRIB+Z0P8KfBCGs0cIXVnH+xYRCwPFFrStQ9/eh5Jj0kmQ3FMSO4bI
n8OrQ41WQl0l7CTXi9Q3xDkFjQDQfpdkdliyPib+1qdkPNBiAVFoOv3tsFXYCbtI0551QJgSDsxu
iMynXt1Doul5pGdjJVgvtQn/mVzceZZGmXaOq3tBv51E6hqLabwx/s9E10yluCG4InkTVc9yFKLX
eFRK8gnYZiAgJc1wFE17vaIp2jDmAwX0upO1feTC+y0tjC3u4aeWypb7YR6HwWGRNfRbH1rfGEP5
qF0JyrKwAE1woLbBRhytg+jLCj8lY3crnegAzMP/2NQAeVPkpZvFHDMkcQQeHXC4d+N4eZriqBCZ
S5rtFZ+en9jdgK50FKcyGlWP+tldVnBneeMWUSNnM0auIsNqUsOXXYmLCY2cZWLgtNf6soN1x53u
3ouuV5j5+byPE5XHncl2eWJ4WP8/PqBt4KUdpKMmEZwLcL6rkvByOJ8/F8YX2+RtLL+Z+xo4dLza
UjN12LPokkLTZPber2eIgwfAeyGcr+Uk/EzcWvSmMWlXx3erjysNNCW2Vpn+7wwx5lfMSYrtDpyc
5z8cIVkV6ZYVq9ayWseshsptkldZHViW8SWuIwBNurMEVETq6XVXUQ1Db6IHUkWvarHrOhSacPmS
5vqCwG7f1wX6BTaAFINTrBSR0ARZ5FDld4aBJt2FKY2ApDClX78AuXLhtZd7LJjfALMm1kyXPK5A
+GuojHGLU1vDe/h360HiUFZzq18fDbo/Uka4aojyMj3jKzXShORYMpczYjGz5L1z8ygNVraOoWxF
gpmiz8BQHhXaXblPvaLb3yFwczaKDS9AosFGrvdkpeGfSEP0qY6TuIfqDqo8S5wO0V7HSjtdwPdo
WADHpkD8U+sJXG8jo4owjjSPyk7MkBpm8yMbP3KScb6ZjakWN7XSwkfCvUlQc8qE5JVRkcHWys5W
Ny6Ha3hb69aoe+LzFgBsPdu5+KMn8geWBhHVUMTHv0h/58bAUL+5ifnIk+usxhFcABHuNXNWGyL1
zh6HLnu7lbn0yhHCj9e2TK8m4lj9jJWX7R9a405NyFDeQhWmG3B/BkceDkgW+2Uwj77aTblqT58A
/+sYbzsChvq5Rmbf4dIXTVwmX4oQnIo5fyrChubql7Wj/aBSktiagpiVzLJbcUWuj4MbyTn5oF2P
wEuAm8cNAnHXfIH6MywyBsOzXUuwjqeZ9yriJfYxYpKCtv5cZDlrwlX9agGflMwqf9/IYiOs6t4I
VLPizAg/xB4Dzib+wiWFAKsuSRPvUh27aPwa0mtM9gFVSuHT0zO8PmakvahpHAogphbSkINx9JD6
a2dOO+kQw/riCxZ33gp/iFCaazk+5/uWPQ8M2SCVsXK3RnrL7IW0QLi4IS0vXW1KktZzk5PfTmnR
gckLx2U4KwHx0Q4WqJYWC2Z1IqYmK4QK3mq+Ouh3Ym0B2yteMPvJkbzmRhGyKQT5eBeH9qbWFMrY
LpiQwzhchv15PUBHiSCNPA6aJbLHnfi8NLEVvuEfN/WLzHExBjCWEhazORUQZCNiFknmNNGH27Sl
+3cSv4emVY7mdJT54DyieeLri0Bj1zicR80PkOn3nvrXD9h7NCD2qcdW+DFbMvz6X9pXqJYJB5OH
1wxHpQlRxn59wDFEEBojcdrFaplVuq66997Se/AuzVNKHbhCy9Kfxvuc98oZO5lPQd2xsUNdsC/1
NUr/kW1qMDXuRrffnPoiZGR1rSx8j6J7n3nlLJT/DM7rjSUoO+ipSbqTjLeZHajTwZhbtGQ4dY30
pbpaNceaBlKvVLwgsxrDnaYvxRnXmpE4GMJcmJWjx5E27MqLI/Mu1gEGZS6eXSpPigUJx20ZMJ1/
OeWrtPdb+2YVmZ5FvuBZR7u0epvx8BvOqGngy/SjVMQf/1jy56V6sSk/vElhsVOHEewMs8F2hvEP
mSRJ12coq4rbHxUmRoMtPlVqsyT6munF10xwgjxoagsz2wIFbxLP1UHBytOnltnCpt4INFw7Tn77
usBxVYyoGQylrWcIMoabo3Rj+Kh6a+YDnPySN7qi9f0OgY6XrZXQiA9HECF0nGL7IetOhk9+Hmjj
kbRe8Tu4WYex94rK1+YRNMRSKtSJqojHuW2gj3jecRJ7oxo8uHr1m8+wzMHQu0C2wco/E8fCKlRU
WD2uenA5T0tZHRC5dPrZrtFPQ6USJFqeG56Qe9p7VjZrE17IkmtWfBgA3LVn0IVhpbHDiXzjS8OR
IUfoRTnB7jHkCHLeE9t0naQgSUNg5aLvRci7vMToNrdSIbtbDbjwpARJ1xVCYJqLx8XQ2CaRBVuW
ku3DyGRLMq9ZFaBgxcjt1QuNX3yIpf6EIuRkPwiVxkoSTEYPYGVjlrQPKWYNS6mfkBuoVIjRU1AF
xJ00xoZcIAne2SkPwfBdkzjrkTLMG0Ge8tsBql3bJJds83+k6sMa0c4L/nQckUB3XW94xyrP5aG2
weAF1MiNN6JbNULPiJNI8K07+Bqxr5ub5vf3e+QFo4jD8XeCbpVfmYvpcK1qtvb4Gl6Z1p/Wo7kj
TuWyrBBQF2d/IqANE8xLi0ceXz+5L93kYSsuS6jDS8IVtoC7O4jEk8iNL7RhHIc7lveggbLKAFrI
07OxsN4QsVLuvrVsRdJ28Nsfq1bUlEZ6xLpTA1P/2vf/T3f3oaih/BpBio41DMS0AZ1/TJafzE99
OYAfF01EK+z6y7ZRLvHKyHAhqFXXk0muwYGPuKHRcq9LI1/hVfwrcai/FRysONHvBqcGLVC2tXT7
tq4vLwoFfb52sYtQF8mS7tCbyJei7zgLTjptiY83SFCzYjyyJIFbnO01L9IArRL0kkrpPoY8TgoW
S7cXlhGqL+/sZymQc5Dw9gKI6b1R8EJKWt47EiDBJYUELtC5p0n6qxhwawhW0OwR/meMCqoIYfjO
g5ZZzaXXCNP6Quwq7FeKsCBVeixK3LtspcKmmzYFjku8H1lUnnjczj1WtIiLX1bd7K7jueVEpj6v
MOGn4kjNxVT9Dd0FQy8RoB53mkhrQTDI9J7TyxEgxSYFlhUgv2IcqHIbQ2wxRcdIYE5FPZedrL6A
kGzIb5CmjUDdoNhs4lBD4y7w37U0p+beXOSQb3bJ3iWoHUgJZ6UUYTCD6zZsOvLn/XKNZLUDlYMF
cCpjz6zq6RoIErVZfO5fEa2w03kvtrSJSPwlPdhfFWj4OfsPvTNS8hZyHwkQ0WYQgCvMOoBX+OF1
mOlQVsrcdTm7asSPGWgnUvEca9yrsgbZV1DltHpv2Kl0Jy4GMM6NrLKeB6NZdc84AAhWxjkUn6d2
DZMY7Of+4ryZ8miM45O7iobxCAXPJBFJ6kIaHwFSo+iEHiCThDAYLQOhnPRc/JRaxZSU/sfi8iv7
ZH1JgQFGH5q0lkguylC6ST4Beh33YOO3+onGLeYPlsLmXfV7Y5iPqukO+zCjISTTJ9qzag2new/2
T7PQRWUEdL/a/3tjrCEFUHHlCmOa8SixD6P32pOattAkHdm2gdozUkxml/QlY+2JZqn95+0+8Wv9
WBt/dyU6T7oFmPMkU15NMNg5FDAm0IQNpAlwkNKXjucTZk/7QX+MQ0VUbEuYG6oa2pqPl6zsNScS
xE3D8rJDu86k9GJU0kWv6+t3lwYBqPDgrvypER+KnDZAiubMSmn+lehEEIxEuI6c4x9Cgo3hxY70
8MDBstd1gHbniIDND2eLJR6I3RUVZJM9O13Upm28uZfQQM32Z2ftMR4bM1QlU41TLMK1wp4JOl2l
mwW0o5wXu+vF9lfapVh++A8KjY6edjHjptps+zEgiIUcjACgPnY32VUDpGB5WqtPKRhchsEJkz2I
G1uunEabmjJ8gFQq7OnjECS+wJ9lZYCjqq5EoZ4B1vTht4sqB+Mh09EQzmMk7Y8bPnM6N3PCWJu5
M6idISqkKsYIaixTQu41jRJ/39xOCXstJrzczinn7j5Oo5DrqbcDv8Ii5nTFcyxgR18zclKrrWDM
WUIWPETk7TXSHIJfLcHmAB8YdPza3pylYgo/CXrZkh49lq3DBiZuQyvhO0kZ37UzwjyB2ybEJ2wG
d+vxxyJj0GBbVUlixGqayCBbGboOjRu6FsmCf/TmSThUxrecj9jqGeXzD3sD+MATvRnJ/An4JtIX
C8eV2Zfa/VW62UZXA2hoFioS09TARPKoJcvIFbrVZXphcFO1xDxVLhl5gwZ3QNmWJ8htyNp6+4EZ
AgNgZAPUAaQh+GQ1r3ck6bLSRofV9DxVLWr2aMELg8ag98K+MhsROocL8wHCESMke1Y82vx6omdz
56n8SYIYJwp88tBzZBgASgLXadMiR6nLCz2sJGZrA03q7HL93YgCkFg8FxaD2QQujkye9HzQ8YZf
0NXB+ggZ8rfiGl99ewEMO6lGE9jrQd2a9AjTB98T7EJxWsQ1rVaESsO6/kdnFWu6Y/FopiAOp+bN
fxGVUNyvUaAkzaozFKocs112J7KVh+nwjuXnjQQiVL5f+t0e+czTSgEPlO5UrH5QR/Vfi8CKiAMf
TvlVfY55ZatoQYgVd9kOIOLwPHQbmIRAyZ+TRxUpOp7N5xC/7nA1d9XtIzZLTEbwErRnpO+zBk5/
iuW2KtcTJ3UOEy1kWvi3EC4O6Ntzvo+Yyqwpt5gB2bl5KptUrQNb69c79r3tsa4O5SZ2Vmgneq2j
f7QQNmxkjxVeod6CJ7tYSUYp1Af8tyfV0d7P2cIpZfH+RR0qRyxEv/GApVS/PzX88KcZEd6JLRII
6ffj4t//eoLhfvk65KZZ0gMLJRoSGnNu2bZIfPMm+pyP68jPGvJtHCqijDAxeBZQlUvyyoJKDpSR
X6P2+/WHEkq9CNrMKk8JQqx9BBr26EixJa3PJ3ok4JAdBbmxaW6uHpelXUeo72H4lxVlKjTJ3O3b
xE/huv8W1xfkRBI9WEVJf1jYpttaPcNS9+ctCCV8pYVO8XakKgX3HFz7P1OWHoKItTqa3W9eum4h
25sO64bm82cduO1jkCXVOInBBe+wCv4zOHOZy4f8vHFAdbHm6YQ0XmLUPR8Z1kRk0IIglOQM/smv
YDwVsBvaUorsQnIHspjsVFz8hev166o23vdbrwrfmEwtI9iNdMYMW48oR7uKuajQKfRGEKI8NAOE
qU3f84F3aSCJXP/XC7u1oLtg3Q4xO5Ec/NMbwkT52pQGpKtQr8Zyby619q5A3vQFP8zlsN6qDWZM
aIUESAkm5obXasxbFZWFJciIFOVdphPnyhcUfG19JBg4RADu1yOxddIcd/UwQQwWEYJPr+IiFdrt
GYA9ZCPMo990Rl+nigXdE8/Hc9LHXcem0xbY0cI8XbPjWDP2eVHiMmi2XEHGXD3gGdZuHM4YetPr
MmA4DvIAEVpRqAZ0gZl78+MGanUZo+rtqBGaLW2FIllVQlfYCPcrPy6IbYJFCrg7yJeZQquvCqRK
r2hi45r6dVXWA/2DrWH9Y39PRgBa467Ej+xWsvqa4TnXX5zZvK9KEO25yv0Cvh1LD1p5NRMSsiEP
oJE0JEmMGi33J9SBAie/2IIBf5RJApZVkApLu2hKBSSYvhNyAcB8OiEDVlu/le9CUODvSaCqzQO5
QnbZMUU1ImHWhZPNI15xaepTA2sJDcdT2IllUUFhV0OZtM7bD5s+Lcvgr7Br5tcyTa3a4PjTSV3h
KqFfwu9qTSOOQ7Fh7xzf/y5WaNxceMWG+WVdtz7bEyEOyH2tiVIglbMj2Vdw1bhYFINF4hdFsQjW
xRR0WLkmplLFso1GZPB01xrVMzI2Tm6L7cHKdxYeAqBB3hCE2zn5psom9Qv0Nk0wruo7MrELHAtf
oDVR97djgT7y0kYo6Ohrr4+ldER/8v9J1Y4Os9OYNd5PJuGfVxdhrq3ng6MN4may3QJkaS2ze8GB
lOZdIh4S1vC2HbjJicxRH5hJbnayNOxmOQf9ewVh1t0r7BxX8yoPIzMdQ1QJlkzXuhobnxA1G9Py
+QbxtUIs8N83mYllcXksWQb8CMvh34PFiny0o+JZx5JL4IdPQSdHHUdehiPsU4Jn7waR6DZRqgh/
L+s+6MPa7IwhLyrUgxtK2hAwcdLKuT+4CNLqurpaH+KiOmJfT/XuLAlqyLzPAL+RrWFgB/MnB8R9
dTrHNAgRvJoh9ZYIsGEpypsNpok17mGCXtAIxiF7sjKqTbgcgE601j2FzMRsiP1nVODD8R//OUb2
hiHvjEC/aE+q6f6jfFywuhhYsj4u9meGQlpIvrUPQDneMrXcuacTOCMMmOkraQXmCb3hOcIm/qXB
1eLNel8ZuVno6qB3tCYCZwvnjPjIqql92jtPWkNTjPeHMgzT/47N0FSS54NTGItUyA000DPrVh8N
spqrg3YfGy+OUJ5hq013HQQhbmLWylaAUlwPc5A1lHno5lX7//IOCtFM9TXML+PhPWpu0RVh/DaK
zuExnX6j8HsDBWy49U5PbILnN2geNHNDHnPqAVvUQmpk1Y5LRSDksPlyAXzpR3XN8nbaUgiT2K2Y
gBQqJsuxBgzwj2nJihPP/6sWGhK3m7nFFm4E13AgyUJO+nGrVDp15tB0tCtRcxF0B4FoMUlAuT0Z
mGZLU7VOe5jE02wV0WidYP26pGINm3n0axJDH6gLTqCcozj96co4dOAIjrcyGNjKNBGk57kTzLd4
EKdZGCGFxWwoQCLDmT0RyrppXsWZp1xmgqa3t2Dbfk/vvmv8YzwPINYqQZ+uM4Cc884FGCVzIt/z
k31E+4kiAmV/eEJmdRFfoulZVsCoqvu2nhgs6KE3kt3h71TsBHrDZR37be5cZzwZg1aY6FqeFKS7
uaDqEHwM64LVi2vKkC2yiRJvWbNMXGpMVKiewz6iCFYo2bUzqlZq+1WxAPLdFkiohQ8aGp3XhGt8
ePue0GY8JmBvv61dHCol8T3Xyp2nTYZpyhhBqwNI16og3ZnOCqkdAXcqVyB7DFaHg3KXRB/ZHiJF
QW8gHCUBkZUXM0iV/ZhUw2izO/4YkRFH5r7ezkvRHt1EgE3dH7HnL9PzIct71iKouoOI2cHwfuwV
YfTxmrdtB8zh1guG6dfLH6pKrCSpOgrRC/oZ3jjKDmC96zUHMfB5xN64rFjcLCVjUnPZSUZiQaxJ
6ClMJ6QtD33vKZCd2cwQKf32cesXk9KU70lnyudpod1SzgtjyWIEOp0IfdlctPLpf7+urc0mtV/I
82PxOGWPoAlzbxteXKiP7qkgvwQQB+QpeOi3hd8rsWZbS7ytBC0BBJARYvtWGd1s5UyC7VyVZ+P2
lGrf+x5kgaB3a+dlEreHz3T2a+jtlqGpX0ckZdNXq9WA5jnpcw/pKg1QzbQqlZJaJ5gThuRgyirw
mB4DGUBD96rBoZkKE4hAG/yfthJNT1bgpoopCxtsKE5lw8XEj3fqZGXT024Z+4k/TObFrUj7pQjw
QyFsHt/EtFZp+J6KbOppnmIfv8SDGkdA/PonYR8CBJdQCjKodNWs/GGC8MtHh3SCxu8hSVjwTCpJ
bSUnxJ/krQt98OykehHwvg8qsINSzr9oTvhrMLQ0GrvheK/z1JT2gxjNAasJNhV8MSMCznBRzCwa
B9Clp+VW3PrfvnzlmK3wXcu4vLn7Ht0HkowrZaT1lz7MD802Y0B3vwwqXlTMbziyAH07xTcvGrgJ
aQVrHuUrikCkFdjDxYvYoxYTkrcN4F7YO/cQtoZpWRtBG3thAI3L0u6mq9FSbzhe2Z95mSaaRNcG
nkepRB928JwXwnJYuD8rN4AL1Ry6/4wCYdvvvpme2iJUH+SSKWID6Sf9Cgty4h+nKXAilTElWS2f
62RSPATctTCVh/9BoJxkmEd7TAqDhjw5kFb4hkj7tO0WyNTOcTsI/qbO9KjIH39l9WQsQvSNVXmM
uxWmLpLVie7aFHojksMeA0mRghF4mkWZkunHmi0aLImPHJl1qLgFZ40vuRzGdEGqAeEQkdSlwy/I
7hWUfGwUyWguTp9XpeP1Pmd8ubaKyNzpbTz8ooDoC0OJPA5L966S22M4gRUSKLRPuTNikrrN/5W7
y9AoMB4HvH2cSkAorbnGHtxAUvp3KV6Uo78T//gx2Dy+Lm4DGvEdZdyO8w1O5myYuVOPTul/oZUP
JtSYuYgJHjTKUqjXYYsE4sxBEudzcFwi9/w2zw7jYd+KYKWd7xp+qnW5DKG0l9yFdzqg/boOVSFu
umIfG87iL0gre9FjX1Of8pFMmyHbKp3nM23uRypPCbmdCvI5om6b+h7WXv2beb0Y/04Ur4eHfN7y
5PhUNC6XV8azh9x36CtnpyO1S/wkS68eHxV+OaQkAsBCPK4VyH3qYubW9ljU/lz4IFST9lcSHW/A
Ff1Yl0mGH5as4M8H7W2uVtAyG3N1MFJw5PsKxNrSiRVeG9YZn72x5iRKK9KwaS83p1IYJVb/qnYO
X6eqyNxmTHLPoilLnuVoSyTepkm48THQhDDRRHveNGc+mPwxhqS1i4fyBtD18eX3aIsqcwd+86AJ
aoCzg8/nvEm7VaDSE6n66kqTCgQLZajC4Y3WSGb/++OlXpboKJhcfbSoeaWKzM+95zYQKHKN5Uca
nsVZEGRfGJChLgPfwhdNDQ8K/biyL1l5KFeLhibXJxTe084hqgB1/9KqwzBPXNttlKlKshJ+2a4x
TmVMowtfuVEH6zrXlsNgVu6g9DzYOWvHWpyKwqwo1y5Ou+qKdBJBGXahh663x51P434hSIFGAz84
O+8AIQVqAElyUKgyurTmjWgp3H9N2q8wQAV5PxV3CpDGBVlPU4MDsz0wtgaP3L5VM93ZKpa2s7wZ
8O/uA+BTFg8LwONUKihQGud2lrqZiZoARd4/0hcDlBnzRiFu4xh46Aj40g/tJ0EKAZ22EO3Ff/OI
VBJkwRIDKemqnrFZq39DGlZeHnB8GSFJtbiLAyggE82+j7Utr75l7Z+MsG6TXDI11pvf1UdtnXeg
v+tvRvXgiemuJQArnsmCDcgsMpIsMsIiot3v0VzeuWEvVx7vHSXOvJvNNBqOHjWpKtU/l6fcbvhb
nKjgMPRfZHLgOYdjS1pCA/u6B1YJYMLFgoa8rc5WgU+4wZk9Wdf/5dmIY0oeXISIVZZJgZmNCInM
9ETwgRy04jO6a+MWRvrqMId59Vf8p5Yhh92FS6QIOR+D54QVLkIhnDA3+cFikrt6/D44EMb2rAFO
ScXasxM9UHSINmNzW/kotD5uJEzYR8mHCKUnu+lg2e0yIAFpXe+VK2eryipJxY6RUWQHsV+Uszgn
pTW9W5MICbcnXg4uONFnNa6AaecTgMUMtFDjK96cGANiTfP6/jvZxJn2fD27lLvmOy0nHd/xKjIL
Y2r7MjtrM9xh3LEsGGk0bd1ZHjQumghas58UXDABvn5jjm1mKdvx0psKr+HQxM0ezIY6lnjuoNQF
278YroN8Z28fI44YheT9KcFNqCzO5RZt6q4UfwlsvgQ03OkqHGO8b+dHxRziMcXzyhZggZaL81er
aTQzLVom6S5rFb+tlDVMdBN4dGnzmD63YcTAnksm3fj6npUiQ0jIBL6OstzAD+6NsiuvbrpGmtwg
kK1gZinwk+4bdqOYn2fazxBR2hU+NFYxV3U7qAfNYOjO/RfrdS6c9dlyzk/JCsZnSZWJvXMIWB7v
bOMZq8tpn8nXjUN6JHybDPNuOypuqYFDADE7qkPYsHqeMPmmG+FW1jzIxyQpPT/uN8DBdARBHZZi
uJU3LpGPZn7eCpmHUslkpbPRO6kWy1cOdplV/Fh8Hv+Kz/05+4hbIQx+KHHfIsfO8+Lj7/60lgnp
83GFxyOJSqVOc6LFqf59/AHrrApPPZfmlbTTz/LGE7qrcTtsYybktBQwpPD/DK3IjqhWMvYokcfv
hBI64k1nMR1gFQtX47HFsPtMzjh7lCGNr1z6a/yOM6gwmK/1udwv8o/8kg8j0qkmo+vCndpE/YqN
0upuGhYnj1AdeuaE52p1Udk9eEL+v4qgO4hNHCQmniJH41ruALEMYlTReZJ7/54s/g1mrCzqpl0W
OHTBjsKMYsIK7hs/vOK8G2IXIr7xDlq+fh89ANbuoUYR3BriMFeL71IH+iJB6MuGaJkUvp25IVNo
0oV/tbpOE0C8TguQZxBRW0XSO7LVyWMvoGljbOvZ1n5LFKNCo6gdR84hgmjwcKGipTgYSZ6mICwa
7wATsfi5xgTODb12xPujNeqgeSEZ013x2rDefCVexu+o/1Kphh8PuIhh7rJjf32H9PReCiqBstMJ
z8rVVn2ijkB1jL1OiMfaA9Y9wh3hrBMDxML8e7JdHBhLEdDf/azpsrBqLxaYslGvqkFX99wut7zw
jgK8H4FeXiwESSKQFxLYDDHTR9SHOZ/jGfusx8fgm4NJ0/yUKH/b8UMYhy41HSvdQ8L3M4MF998y
vfsypSlNtpnjXTXQ72uogxkAj01BGkavUxIz3keOMyH3OL/tG1cKqhHb4cvQPh+nhYys5NaZHPfu
niMe74qV59xtLA90iWgr9Z9t/OMDD34SK374y2yDXQZE8uMUplhKVdmDRi9RWSNyBwO8OOUqzDqM
jdKD8kL7QH6v/ZMETYrd4wDxL3bnvWuS8Wzxx/HjpgoDN77IBTk+ygVlw7x1fkoCh0O6Nmermcqo
tXnsz0zAR1IzmbXAgJ//QW6R0GeRhr7zvlVaeVgd6D2Eqst+G9U5SW9Q1wc1vjwcTVHGCmDhzd7e
8ibrxGyMtFsqGC77mi5GY2m6WSq4jyVMlFV77kchTAy1A17A9LydAunNXNKr84Dn3w6M7+Ouk4yO
eq3D9gZIMQmVerIj539rr/dmsBJne5CYrHL+N7/YnvcoRWliKf1uJjoZr+MzsKeuR/+/543fKP9w
+2gsoj5kQEkdCkzBnKwg4AcL/pqmHInVFKUE9pPsnVYbe9BiOnSYHebyB/2MebWwS39dCBVATwti
s62i4wso3Kv99w7o9g3K19b2nZ9Eai84JvwLPr4+bmHJsRoPUS7+nWQYEHfrVNcCi9m26RMM9nnC
fUTAmk1ZutIxMum5pCTRKcA/UoB0pZzWA1ZhUQ9LB06dzBKu6RJ5AQTSOZ1tmqp8A9Bbita8W5vf
AnqNuHlva7rvx8HI5oIR2CD8SDOlUQPOLUNCbryal6gFTMnG42L1OsI1ZJEh3dpFsPF8z/NM1TQ5
g1twLBe9fIcXr1Nj0aX/wP1KLN68OC0uIQI5jYHCxrpGWYQp2mJJrt4z6o/gs4Lac+4KT2p+YDQB
UGgAbXEKPzqfEUXfWvoZiC8u0ZdO9ZAawTbTB1tLn6JuiB4NMwvuK9mIR0XyGRhXWrxyn5t1M4D2
phUP5Tyz8HXh0q+TzkAG1u90Ng2o3ZvoEGvkWzwXCQZRWOnCHZk6LF5VhmHO56uL/bkkOwAhX8RD
7tWGV/7TDPsKBJoDW1YbUJB9ivssB07eP/qRNa3KwBsWRAml2AxsXeeUNu7SxfWQ+TOWeGygfD7P
rx4e68H1KpjWcqciF6saweNtlBb3K4kxNn729wMF2wsWctUJZplS8xbqnGyTK5hjrUjLZmKg5n8m
7GDvD2tXUEIHgV9gidtFezQ3ARKdBNcUlFV305m3IfytqOhx+gOi8LnZhpOAARagyIqvhHo1Hn50
y0UXakdfpUh9Q4fDbtYzaJxeJSuXeHR66/puQXBkKMfz0B0ELUpSRYdvOqxxhqN2i6u5fcynWrha
jve6ohirAb5F4eatcOVIkqBG1/qisX0nehq4777til/0YsFisAlq/ouBmdloPXodmcT0hAQM3Ztj
hd5TfJ3dDWib6ljjsBqJXmqcTx1pLF5V1OtM0E+fTVhvDdKdbMuEKXVA3IAQBZpB15z9dOImgLjZ
0ynWV4OlWjE+UL/M5DIYPQ5aGtuuZZkvOcM1BiJE0lpY5hneQ7Xi344oLpDPOdME/6R8uet4VulY
6/iJ3Q5TyedATlj4WSdAriOOfPlttNz1yMmGK+3zo0+zQ5ZfMJWnqIaQoZhc7Ou8d9i3rk2hF+Ao
i1hl7CC3BcEnE0UxjTgDbGWT0j/mFJ4C2VUcm3in4hfLI9cyuEwDeHLOOOBZV6NeaEXookb4mLEL
D9c9e80t/6ZmVfMnFb3gAthDIe4hUTp7JkmdZn+rofDuyaf+SQw0ZC+76wKem/tK64qLJJ+eUvsY
s8y8/JgLcRVjBwK5DgrcRlc4WMMDnuFPz+E/kLe8mejduQK0ywDZfdaTGyLHsY3GhLPjlt2eBRQQ
KlcVFcjCPKN4eBOiYXTNIGCgKhHgW+r3pmqcIzk2/7ZncLMcVE6bWRk20/jzmUmQA6qOnDF6e/zt
PjFId7t1D4NbETnsjLoXeD2lDhVs7r5NdIT5H81k/s9gGzedgUxBUM9hnrUiMgPiQr0whShGhneU
6Fo0BEzebsNX1eZE+BAFDf7fioSlsSXlg3LDJyJlxWYhQvhz5grv+azbubSrBKvToUCn/Myhu3aV
POR2SgE0Fmzzihc3qGOCx7bigaupiaXewO/hq1rdbAEH80VZ5ME4Ut80x2RxxOalmXjZzh9ePHEz
TC0C1EK4Ulq2TLxQkiqcLbkKLB4PXV/+JFEFJfc3LJ0diIVnJB/N4wGBAohAaAcvH5wvBI4QUvC7
yypPJOeqibYUYkV+BH0OiI2jTVd/pw7b2JaclIianjjTLgt3Hut/a1BNvBaYwuIVDMRo58UVKG6M
mIPiQHZ58+KJqo4DCK6pzjWFtNSwM8Pg+i4LQtCjPcEqsZsN8szMEWnApSLYsDcO5SmXZBVnrPpt
4wGd2654vefZ1Aq4bwBHPbZDWvQkAwGFwofPoSKLTI/szirr/aEOor7d5SgwR4uc2GzFtHCtBujO
wgnQtfibgDeWLb3yAPJ8nTYfo+VwQq0znGYxoFQG0N+KslABA1zUkznf0KDtrcftFC+VpilriKU0
QKslKeySsTvS2CdjjZsMjjsma7oHSYhrqHoLsjOcVuXK5bmoq8+elcB8Uam9ANhq0ESSNq6ugfEA
xmRs7QWQKK1jFSrlWBYKk/oK7bM8H+vUBC8Iv6aVnmjjpX4kTsy5GIK8P+i7OTsp7zI9JiqNZ2Rf
WZz9oHCiPdtnI+Tt01hbcSdZnzrYduuwMkgGmzehhTX7EfWIIjczvBMhN3HAt+iAYORGEesmUE56
iyQNOuFmzR81sMgKLembwqy/2Ba1JnSgueUAqj3ts1ZDZvbaxU00fPEl/ZxROz79wpc37+ebk4oR
vAKSMXgG83YrnYZANsypDXFLwXowtsERat86dos9+zG9C9OfLrw/Ubgdpg38hQeyVa/MmaKq3hC8
fYXz9GjvA4t9vMeJ/mgxWxKW0V9qrgHF4ptBYNENuMsFAYMqqimizsw9FV4ImBoqSjO5R+qF/bF7
tFcMoOcgsAVy9llSPturhluxfAJWnt2ImsBcXCOvp7Okm+MaP7cu9wk1WTlXlsYKaGULCgbe18ir
FXyBdRvBFTHVMrbm6lPhGdd41VoNLlIiIcKFeJRqjZ70yliXQOelIuerAP7OCbDYmd8J/G5VGZGU
+YXe6Vj4p9AtNCsjhYYdDUmxRB4ndDwyhWNz+rJJtZTbFPxUomlzcmMAHAJplFs8HN+rX2JAz/Av
5rk6E9CNoMJ5y5OdqJY0guk+OgFlIRhBOAIVU01hxq62TVsWj002Lh1F9UUxH80dPvdQhzdq86ZC
nEmTYgDinsko38w/HzOmb3tS2fFIwfnnKvqzl/Tqzp4l1gfmwdOeOm/gdpYQQkbkbfgxeY5ClFZ4
BoecP7nvlNY4ceFbsGtk8gj5Xeku4dr/tj3DDFCujpHwHK8Ld5mhdBZESCrrD27DfL4M+q9ENQ02
JT5kr+uIMsmtVz4NP4FLr4RVC5l7VZZZTEPxEEsr8ArcK3ZI2xOscyOBDZNltXb/2qkK+ES9kauP
gMvCkXiZTydi/vq3+dpOu/1MBq6Ppej1agkXZ7Ew00+rTdA429Jiff+fBq3iYJwWez+V4ymq7lZK
NN12JND3rUSbewOybkp31UyB2lGXuPwsKAXcskZ5+Yjc6AWAjRVRHS5IQYfxzT4F9/gCxA0x7OFX
J0o6zuSBhaKCLY0a4cQS1WeifUg2HQan0cdav5rV1dhBOf73ENJzTfK7pQFAS5amb7MbQVyTVTo1
6ppz7cBk239Q5FAO4as0OC4tQzNVhoAoTOlTDvL8Qo6i5TTJQIMTl7l0PCNSszJq4cV9IGBtlWTU
Wr81VozQwFtyR2qczg53D68TRiZDr0ZaGh1DOxsIIc7tHojrfsvrrJIG4OUepEwBtdAHFLZv+WKD
tl1hGYSup98x//mh7vZ7pwCckm/cfKtI0HMdBy8ibDlxKrLnHwvCWeCz8mme9atrxEG98Izcx9Qv
M9/Mbbp2xP/XBooTehwUN0w3T+WYOZKnD+9B7hnLZ3Yc1XqmRu3qb1SoRkYie6NWckYhJNOT3ag5
Pyvd/6RYMpUxl6RxXNzUl9fY4ZABgTtF7lzs/SW3cZonarWrUDf7zfoPeXfhHynHng+w3NUHJ0C9
aTX+r2WXKc9l+1dEuvZQRmLuhoKuztJXi8KHT9metU5jxnzkCTDyiCByur3zKypHP0aNGt+aFl62
3NQHzioUy05PiZbjwtfrTZYeBMGxBnuFTXlpiWD4uvE6Qi0jjAbxcCmEGc56Q1lKXFme4/CCrZyD
ymjmvzt/zB1jpr7bbUVDPGFjQvOQLnl4E8plVhVOCj/5yhrhfG2qTCHWQR8u2lCyYSjCn2WCJHSm
ANPfYH54pMe9P6oRvkl7RrXhTJN/6Kzp1ryvPp1iVLGkJIELSlEPZuaY5mi7UUWCs72mVYJ1dswt
2gTdTN5emEvon5qNWEPibYPEf/VLqMw/rlT/LS3/ZPZBaG6zukuBQCuQjSjTzJXOjUqY5n62WykU
GiD/Ep9fe7HOtpBIBbeELB/juVzEEC9jhE0+B5WgLfbqDSbeIxIfCjoOGp/iW3hqvTO/H/D8TGIT
Sc7rJVOQGFRr1Th/XK2kWSlMUP36YydmRLyK4RxvUB7fj7RH/vC1xaz/laTguhrxHhdtvJC0dI12
45caIw6R5a4MuTxZvL/LO9T+UhvgMdSX85w2Dm4qmvIi4MYzfQFmH5kp8z3Gt82ugJoRkO27+CpU
udtN0IjbDO9CElj/Ws9YczlwL+y/OGcB7hOUTQka2xaprhvhZbDFExj8/8JMt8mVzclXby7M46GE
J0FxIYWkO7Wd1atiQye4XZIt4M+cKgXeqKk1DQ5R5Z9cZIlHLrqN1B+iKuPruOjY2gTVcdPs2CfQ
HUxIDPO1JV2lUeegfVedgg7jG056NXgrlMF/mapNsIVTe/rgPSfT3bQnBM3OoHNjREvtDGW3HKfR
JcQ8+TFelSUu15eNmLTBNOfl/RTKIaXx4LVOh3xIMadU4XnpXzakjYIWq4hD8oJ4cEMreN8fYTXk
IPFNw/eQr6U2/Kdr06A0lPyIERPWZ2CNwW7X1MljcvX0200w6hQuK23vMr5EhnDGvKgzgwZkR+3F
gzvwsjcHppkrURURua07rvqr2nfFdsQqyF9EO3SS7KANe3478Scy4WPMQpHO1XcPYNRjwY7Z1nnR
cwVKO7xeZVOGbsODFCJv6BhhVYBcSJY3b3mDz77ddMKbwVtA/nij+oXlaaUXF85Zf/TFvP9+xXlr
j8PYxfzJDhK64k/PKZABuUV10gotXOAN6pBV6Io/CckqktlqIMdOGA063qUfFrZktDLInlWt0T7b
jRGwS1AEiFUz5h7awozzRG9onW2zk8rU7xy2ozZu69fiGkPHgZwkmwNQg+xVOu+3ARg1Bzcv/yhZ
GduJAgCl/Ikw1vaFHNlzymy7K4Pj+IXGQseYBJQB+Y4VyF7HLlMfwUtjhIoFhrNuiRN6li8Ms2g2
38MpKwG0X6feGMTRSEKPyx8I7F4ssrCVnhXTYgIzd8C+Q7OaP7R7ZUaATnUrd0LNrjbcLtLN7MML
MvKqbwA5j3iCl/dKEtswksSiuaBc6eE6QNCSir84PYSQNzvyLWbjZaD7E8ZwidGEr+c51UJ/E9kl
XemwRejrV3VTv66LDw5rcolhHp6u/s+TS3RPq/D2iFwr+fVAktfdB5dNRUW1TkFxk5tewiBOOn+n
FEOHVQOJ6HQcyd2v+1TtWWtZdupzqk2eMh0fJ9pW/viDhON21MztDbYmMPXIZXWOdLcIMu+sIk94
iOqLhviS+1rgg7ePCzi+gE7dFcLMq9I6QgCYVe1sRjL/Sk5SvOUbo4Vw8oV7SAgN6IV9GHIfjSn+
AuhjTxDGq+ubTBPqyMuZH6PGToSuxS+uigQssLYvWGeJWVodTdXiHgpn4yDJd8t6YnF+h2LMeXlV
bGCBqgTSI3F0mM6fiRrBJ8dUCKV+mqb0kHH+JzNy5hAi+r0lb5VJAHlC0A7Zvmt3kET+B9l1teN9
PHJ6SJoURqhad6748vJePv/cHwsJFoTEiKK/G5CouoKsSX8hH7lWEktJSzJLWBHOjCBCW49LGvoq
RB+vTLG416jFbFmr8AZhqxdbMQbHseYXHK4Jes/Nb3BdkbbTI60/nTIOznsuKCk51ceNx/Zr28PJ
I7kjTIAXWgPYHXbFFZCk+uDr9lPTK/v6Azv288YkwjlMyINQ2cxX5iBcxeEK61r2RUkhUiTq2dRM
vvyFeF7+7QWPQBpIuq+hjQQ560AeYY3yqwXJBS+jZupamnXI5uN7fAPz1hyMm5iYeXL1ToXEMqTt
vVB50MqiAUriLsp4UvmzbPkJpATAYpevFRVtbLwaBezUnMy/O4OBxN3YCeSbxNtRwiLXHHe34Cx8
Xv/E2RVatjlXWRAMGxZGkYZssuPjSNvWB1a2jxngVfHwxrH2s0aaWGGQyVt+fAbC/x80ANzkxIZV
GwUgoSZTQS+Q1yP7/QRkh59xvQTbGpzmO0/v1O7KCDOTlqsAc5zqZFB/S9x9FLdX63QTLE0QW9OE
So0Qe3dfFFpD4bRsvi4Y4MxjyCQPY+HCyuTKxJ7VRKtQH8FyGJb0gE+SK3KAzRmpMT/TC3+j16r/
ggJUSnQpFsHQ/UhG/VbDbIOjM4LyLiSD47iQB06h++rbztVorxHsp3pifP1etC0JWHlRKTfKUJSt
t0TegiQufUgKzeHoKGYS3L73HOK4G3MP5ULdUKtWTbIb88H9o8kAhQP9fVzL7WofxziaeiunBrOH
EErIJlcsohHXLqArhjOrj8wf9b9QCclPXLaGZd13Ts1KnMTNdTsCu6/qv0wLvr6Sw6feZEEeVmpX
f44GeqPSzrIJZ01pMaqdqoAvQiQ+qfC88Ppot0UPjm5RiKPl1noqei9WIsvZ2FGSvhJjl5n/ajjy
twLff36Gf0/hurzuaCrUr/ivAoGICq+CT+SP+LrxwvnD9SeTcuWISv0qlCu1AkFEQRNLEChY67h4
Q2fhWmYe+XmPP9i6nd08oy64Vvt+2yFn/JDtNPYn30fsGtExyvjmDHQkWwoVcP4ThIEtdZMp9g4b
PlqSjakLWOQNfICFd7PGDZ+tk/mar3XKTmX3eKGa54bGZ7Op+CahJ0DLocSpWoaSLeNy5eH9nWQT
ofgKmTDYlje9ymbh1qcpk/ZQMdY2nwkpLgA00ZHRl764tqX80NyEXxMWB+wesIyIEy1RFfTZByKs
nH+Fre8JuECEzrqpVb8GoG90mzSNyfWcy0rb2B1lir1xdPhxXeuCq4desYz+ZoakROvzPqRLBpZD
F1tFgkd9rth9hNe5UH9fPqnxrYrAhvmZQKn2VCIuwAazKbRgpu/AiRxEV1iqhlM9wOBPj9GL9jpU
xMTgPrBPJM1P3E8wV0pcgofUm32s223iWCWYiDafu8IXKujlUvTJCXcVt8L64GMtGImQpbh2rew9
NunE/NQ9bBKBTPNVXNKMRhC989bhvWAEp+i7joNYocjBK55jPRZ/vHq4pA4Qo7MofbZBS50krQf+
WYoS3kBcNrz4l0z5xP5wDthxXsjv/wgCpfLx6pQNCKZGmgxN39Kehdd/DQMF8HJntSaMQoDUmJGV
Gl1OCftdnFSSHlG81ajDAROMpjTx7xBC4gcn4XUpb975GwpAexuTFCcH+rNcd9w1eS92/yscNDZe
LUTwMGlzZJuPxbIBHq+siCBqCLozegz3DdPBPOsg4QI1/zgCfTUmSdDTO/C455JLP1ZjZYzpI5It
4aaMTOewOJtGBaOfK23hlj6niduCwgGV2bqSsWRh1+PS2YM26sfNKxH8mSKpvRJUuZOXTcqGVE0Q
kheXNSrgXTw0fabKyCE33Mx1o9908xM8loleaGouJKdXG7SyiGX3bfqJA6BfnGWPoTCDm16exn8n
OFT1B6MAFLeaHgLE+cwQksSikVcHwlc7hqgHJghDy2KL8pQVDgZFIvAMai3HdbSPQwki3QbNJpL0
GyQBCa50b4MIBHrB7bjijEE02JojJhqKA6eJttgfNwMEtZOzga2H7TTpmm6U08ui1R0VbXsR0LpR
HM6GWrGGCucH0hoA+VhIjkvXAHxg7D9HWVQCqQL1XUzllvw+kRmeNiYtJkJJ5ej1ft0KrhmkFmOG
geXnStL4TnERE+/cwgV5iXn+lLTOMQV4zh/a889R7dYzaP7qnxX6KblJEL/rrh7u6+qc+EFP2hGb
GPRO6UL3Grs4mXH6dPwH1nkLulHbC5L9X9rflQQPa/a7789TGzzh6yZPQ3M8GWZTD7I+LY9x7ZBf
B3gRZB/rl2o7RLFrAIzHoDXr0Fa7m4EPmcHoXIuvR30lVRRFcgH83rp9PBNjNCpgYeUb3e9d+71U
bBSOFXUMFUaiOwCQSHR3rFgQpHi5eXFAFaR1EdDbUoZ4pRCldjvOBxG422t45EyUxRck0PNGYjwz
e4x+Uggz/Cwml8UJ6Uio1WrVLbZeh5GyHvetl3bcs+UVV1ABpx6ZGRvACUcs+lmZkVFZA5cJ59l1
HuyZm4fxIsZTM92MpAjYRD67WOIVFF5t1CtVXriImEeaGBkhXlBVD3yaHpvczZTZXVABlPH7byN6
qOEVVVWAlyFZUyQneOFjjuYz0OSrZjdK/t6bCjGDwCn2DOQkM1m5pbwOqEVgSWSFL6sw5FlOPbaW
bpn5MqkFPuebD2pLLlSMP/hRs5TtFIvVws1Z3NU1+J1kASeOQGUQoQzk0AOhWTIkxE0CL7K3pRHp
4Msumm9USPpgG6UcOe/38K016wV0gRF46d+I5LqtoAqAfRN7p7vmX4FVjf1VzpdwjxU9NMpCM9po
PqnM4dsxQf8r0hlo3BdjsmQFGMEgvTDf62mxeRU7QK3hvijYy6FZ+U51s/GyOUDye5y7XdBKUwE7
c8sEWUy1zXXOOc7C1kPqaQG+PD846xJdDvmYe+Di42t3xskQP7Pz3bC0GoehYwuCFiERlDYG7gXt
eemr0cRj0a6IFsAgDs4NfNy6ClH/BQvdg6A1UjR8g2X94P9TQzSJF5GBtl6l1Cs5jpRGVz94vQ5v
ZVBeH9gLTAdLnCoFtpPH/naajdit2ZAjY2F7bZkrHyk3zYUrhEwbUrtJqn5rAGHP1Ir3RayOn99i
ZAdMxqCn0rDOEUuQe4dX57Pn6JIzKL8iX9GsnklH/cLIB3UlzbXyXqETd9uU8yCjEsTMEft2u+MN
VOgPc5Cdd0klHrDEmEzN18I9eM65VlkFnl1ms1pvVa7HCpcmjKr9h6xXiZOWycLlB8x0oaWNYCuo
pvAMk2NQ1NMDCFKJfZcDXSSAdW9rI+HmdaPgFj3c4g2Ut94L7SRZ6tVD6Ife7FC0KuI0YMf9jdLM
YbP1gLEGEwqEW2izYgB5/HKjUPuIuUi5pS+2hI/VUVCHC4Jq4bctTUhpyi3YYkfz74ea1xgQOyxB
wnoaFwd50njKMeCPFmH/zNUgivNVjx4qnV4ePycy90xlgo36aCVTm/jAcBSNm4do9Xb/IpXNZgyt
n0i5RVKTK3FX7ywv5HCYU588zZ/kBuOHf1492i4N4Sgl3xPT6aWKG0ifiXdxOa+8whyOeHnYOIhQ
Qv2WKsnDAa2FnpKWjAp1wwcyGgyVOrIC4xLgECS7UdbUPqfJY6h7cWrXMbSyWK8ZAGPKT5bfxAh1
gkqzxx1M7WN08wcblkidxiUGpGXZUWp58h8Xh9SaJKFP8o0p9LsrnVJpb7/qS2OUXJn7fU6b/D9e
hdpVxijPXUgipNUuj1jv6Gr72uXShfdeX9Or2RRQUhS5kktDSMJN4S/Hrv0HiOov4kI65lkgxkv+
lHLpxhSM+y2JyK1ilLdmrWZPW1KJvWtJ5ffuYuCqriEtdACBrV6XSf1NJfVHLBA/mCg0nEuMM+oZ
H2XLI1qkldH3jKQGxTdpC3gaFfiYXCLcfCwYBa8UXt4q3sh2L8MJtfmjlTp1SWoy697KUwTDCtBa
ttZcc4yLzbjEQjQb9QAO7CvodUoBMZHWtXC0y5YZoJaXlQGxtrbo/5Pk01CdDP8iHUiTbFgjD7Pj
ceDo0poXVA9OSQL3uj2ZGZiqOWOMMIHJnwN56S5MQqQXZ0ANlHGuDzwmJgHg93Rn4g7I1g2E09ZS
cOo3T9m7IOmilOueEFZMGHa1yDVh20utSWXwDZELEEsz34bOXuxodzpU07lXEwVRa2YJUL9Lo7WS
hH90RN72pxiBL1S+YpWQwD6upi1j7CD0KyPTzblwPRzi+E28nzcMFBnvu5KcW5Ggnm4aFjmSU9rh
oFuZghFsZIGo9qxgWSV0jBULeOMlUjjZHmZ93JxOWLTFqe+0pPLuJ2/UhNsuTf7Zrc10qOXgvpXm
JoEaVPzcNygp1cZkdUWK1MIIfkOhojXOvB7nsLFsjcA8qHk7T2oKsVzQSvqsrSay5xHul55Q+I4+
q3vMmMB1YfPhu9AbtSWg9tjsIX1ZMcMX2a0mHE5Rv1HYgzZe+NYKI5mr4GIVU9izYx2vmbCexlEH
M/3vxsKj6SzAcNdPK+yTJ0VQJ3UqvTWVcfL3jH8Y8dxAK2R0gvKKMS7bOyOltaug9x5NQeHmZd9T
hZ+KeDTs9O9DcgbQjOSbARPai+jWd2ktLE9AL/FGtmGRbj9rcDm3VLt0vba0pfjKmOEEzEo+MABu
g9svvPSXzoI7lo8o/DTDKLUiLGXTJ61Ijv8BCC3bIfAzBWWLNRKv5YQifnsCfToWbkNlcHHNQqTj
k2plTRl2JvO/Blge2/ua395u7iAjF4ozsnBHxm1tyr8mk8OT5ys5YFbQ1yrFH3aRdihOEliNhjTu
8BVhNBONLNyvhC+8EYedEpZrPwGLifbD7YCaUk1TjmtQkUEjKbYOonHIgcmtiSBZser72gIzu/5O
X0Z+f4JG3fQz318kg0Jstu6Gh3UbE2keHnlx2TtxvQjt7pw9K2x4L/zQeL6zuJQ3RhGl8DKRoSz3
B8+QV08zgpYjpwgfPoEVQJgKX8rQuiBZmcwDo0gRlyQuEKDZvax4M5tnz3WDkcxPgLppQQncdA3k
wTy94Otg+GGNxdMCAdy5YPwMmrrUiB5bj8Bog1xlMPXYcr/+OsTs7M2li2IzCjNTfQ70u3xwmDe5
0Hq7TSEYOpg9Qlgzn9W5Rz4ZmUaWoTPEm8TMeYMuzR36c0sgMUBOM4JpQPXA3qb8blEDu8O+E6rf
CHWh0mddW8TXb4Xf+GKwwWbGj+p/Nc8DTJvCsQgHk7UGeUR173XXQ2a8eGKB+QVjxK6CNtgs9ikF
jGYD3nPjfvIQ/LZr7nodneiaAOT3bc6YqAl+dMFU954IeTyEyFNIuFPYfj0ZzuEyjjUiBq+CHCA6
psbB95sDC9hDwb+RNCG/pYrAogTvoKioZDLbHBzCvkfihH6OP+SnnSfN0vJcKqXSl1yUeTy5Okxe
L+SGEvrbDOTP3zOSaCVe6lDOXYrCQCDhb43q9HlEPvU0+GmEfA3l6OpimwXAnk5Hqln/vunpob3A
aDblduE9Thwx2L4wkCaKU+4XnWfNL3ts/Grnp6kNkXGmyupUMN8Z9nd0ALc2TkXrH6aNltUdmuSz
RsX5iyp4rBTpqoEQJ5jFbqO78coYvf1XA0DVcVnsOEjecjqlXf/A/j+dIdqukRKmBzcP/2QpRiHf
kq2+BTaZIGRnxWJG1BTS25Pt0XlfHOntEntMAjwhpGimNUK2aC8mQjiBCzYJBVPSZ6ZCXZh/byu4
hzuqzJVFLOQcf4SQ3ijJqmWEFJAQf+ddaaViD1ekLKsGf4aH6HZkxlBNUCuK/REFOY4WDq761Tj8
rgvu2ovUa2WiPg/l20xTW6UXNqdScdUsx9blYM/+qPVgM7M2Jl2tVZHVXwTHFw7CLUEQCBAZdJ0Q
SWi1GpPsT0pXwMCJ1j4ae4c/crCKE4RN1SrZdlnmb5GW9sAw9YvAykfNhtJEFYRY5KSGkFy1S9Di
ilKOZ2bgBxQPh86vxzS5HgIk/FPh6G6dPZRiEwmLd9iW62RoDipGYzGStJ1MFAGSwy1VQ2pyiyn4
WG/0swfPgrv47sEWTgqlcerUn5xLELIZu4eQ7kNlCpz7KHXTJNB/9w5lnQ5+LWeyK+h/tZ8bqrCt
YF1cqXSAUl7xwnb17jlFWQuQ+OHtLue53i9wm+lpkw232lkHM5ud0iUkurAwyeUUDM3mgfV0HWyf
ue/ED9WI2kppgwXJbB6eSnQRMqHxruDJDYgZrPfP9CSU5tTaT/z2YBJdEWgajXuHSclak6k8tNgL
73x3hVG/803Z/3f5ZG+PYUYCrfv3iS2bBI6DUN+CQa64oO1M0IP33X3IARcpDTMZ3OledCG1PpF9
+v+PfggAwQG+fYl4c6gJFUP1Q/HMAiIR1crJKuY2CyM8EJ/ADOYPsJLhRnvj1s2+ryLWdi8SFaeh
cUkkyxJs+U/LWTOK9UqUwFn66lcglg8vL2Ch4fdP1NKxKP59zA8Wtoqs7hAhX0oX9RUE+Zr1IJK6
XGW6E0O+saXFemPB+lYzToBomv4yi3OQVTpRkKx8dZcFE1VH74bgTavUPD0ILFL5WF7BreCxmzdy
YBtLm2yiKAqRF0m0yhJNG+1T2E+agtdfnhsnEepIW0SZCYdrakQGExMCs71S+DrjmYf8y3QePaqT
hb/DkOq+5l8JbzxdPLTM43q+2RLcLptdqU9QmT3z2+KRPSsqkjWRtihW1AhdR1S/UThbKS6ZWUaK
rhw6pd7FE1lqwRoYzxSQesDaRUVPqWdX3yQzltu1bm2YvX8OlJhWhLvdj0WGKxedqTO/qNDSPwXk
llwE28KNhpWE+OtEiETNPp8cxBS+qyf0o+DhueWlMoZ/fmHqp0nVaL7Lq4+AmaYDr/NH2Njiyonn
ygVFUfxAwI5fTikRdhbajKDLnkUAa7rweSNbuhtupm75uDxL3BDZOKh0D9wG4jMFl6fGn7FYu816
NDPuzS4xu325Y1Pqy+C9kYyzwDRRxKgU7SFXCgDDWwMRu8GDWdkpqhbjyj+FjWN6zhGKEklu4ssh
NnVCXsVJjex9+rY/Ux0Sc+oQIQF3qXcrZqrCTfv3T/bR8hr298/URE17HFLZswVoz0gdQBcELtaM
WnSA5Ptm2Ei6F6glLeesd/hHUzrROM2NCrvOUxw1jCRKgznwZBrhpE95ERosmhiDe7sUMkrtKAgG
YcIgmwSTk5j7GQU204qYGln+1I8kmVxPekyIg3vXLA1kJ7c9nvDJeMlVcF58jh8g7nQo9ZeICHe9
r4wxRq8yaaCmUn4QIaJaXi1UYezqEENEBEYt5tfKnRgJjComCpLOTr0qoJUCY7l9gzK0ZX3rbe0L
KaKj7T8Ipalx2xMsBHWUORysN2sK0472n3UOS9kU+9sTCQ0ehQelEGWZ+iDzTMIB1m98wP8urj00
xM4fx/+2dcva8+qc7nwB5FOuY+ikzKjdDA2vRfRJ1QHGbPoH8nJPth4mb5lYsoupsCDYfjJ7b6OK
yXMVRAI7tJKUfeKVLi1j4LMLwUleYBj4ifBwlzuUEvTM3gmH+zmUXWZ9KkS2QrD6Rxkw6AAbsGDO
2plX3SWl7la810wGtQB5Lm1s4y5Mdk2Varw+woV6NQaaUsrnt94MlNJJXfsv08/iLgu1id5rbS3l
ztBajc8lsKzbisiFxLCZALQVjMKjeW6acq8edCTCNsp84wQ/IER3KaC2VFdpEkm7BpdJY6srQKqb
yJTX6kx0J5BEyPuRXf6OPpgLntn6pQmvQaz626EnIOsG3eb4erSLv8kj4fETAVz/CQ4wxH2VgVF+
pT1Q9QPH0HUYdsWhjru71y6HXpZAmDkk3Mee4lj2DSyGbsGpCWBqYf0MTcN87fqny/uQr2mkgvQ5
T1XnJ1uBK6iuFEtdLOI8pWw9YmkSrXC2NRFMpXiIg9I+HAZzrKv92Yfi3tJWTxL1PjldnYrEAOMO
JWbDoRVbC/ClIW5+7eRc9G7nJCkuYMmXYD2+CzUoG7JxglZpISGySiaTKzrktDp+9rcKIPd0Z5DF
PZ1gJhzYMz6VD1cg+6Hl97WvflqTQ4pwy9fcBKNGDWao63sLR3uqwlPHUdOo6+yF/qlg9J/jGpSr
YEEJFP/nUTSPDqvHe2fbdS0bgpfbFPVQABnGMTPV/8rHPTHbey5n3wib29+nOjPC2nn9KP64TsJk
bmUv2odoHpneA+MQoRD+8TAQSVj4+O8gYzv7zbRkUvoD4Lk0Wg7pYaq/QtWbhAYKwEjIOBuUJqcJ
p+OgYpzxaIRUjQwWFzSZpJKWoYmClTKa1sFATdOeGZP/8ie1u0Q1S6QuexZI72Ymx0oh46t0a5ot
apaxMisIHfGGh3yMawclNZyddkarV+g2HyoE5fWAgrofNyzpD6+jFfLXlbUzBvvOlUlZbNg7DFb9
yg8XA8Vi1d6ew6ZhTh7v/R7ad38bLWrpuTMSM0iHF1eDRLtBiOV46Gyf/Dv2GsnNQHcLUGuR7ZDs
Ndobve/NZYIkytSK0WglEwMDXZFpFd8RpoK4SIWX/jNtrneyTpABFshEKP0m27/ghTrJBKaQbcG0
GO2jBGqho+YPmk3BC6pgIdO0loDjeYdkFXpvFxZZwVQVzAHvgKKQ9OI4WAIkbuzakXHypEbFhtSA
qVer7myDwXh1QLC/lTUoKkUOg6SyrLmTTRoHGezmJlRumlyeJapVp1DfDGECbLlrJd2WoTZoQLP+
Qb3IuHwYF9up/FQ8WsGGMeR2vQErQCy8m1C8m3Ugfz6/Ddr43q3zCKrzzfY8fYvXjqvyDYZCyD10
H9sGNCTiMnwPbtE0RPxGyNlwVmFXPnClkjDz+2YZjU0lxMUgXOiddD2BFotn6FoGUbvlr9xgrWUc
JzK094/57H9oxYtOG3/MQpZZpcSqeyHsujDUU/FagkXCbabbgOsoG6z4dP2XLLLbfjrqaGjxyAEv
oEmTrnvrnR9lLHiw3jtX2gepNj4yib9cTKWC+ywjgsRyE2TtKNrp9ik30tbIWUOmBhVCH4qj+q0k
l+RdovWN5Whe9I/Gilgv75YW1UuJT+MbiQdWhwpBjpEiFnLiPaed7qYvUnPfhwYyQifiRFvFDgPX
8ME1Q8a+koS4qapL3jZGuebpU7r36pGc2DGMsVl7J79LpnwpzyJdcfyMdEoK7lPuWZI7j5mAnydi
C3TAJcgaoZAX9/DFQBcrkBjuVmgCKvZNk5lfBvSvXd/x3naSbj99PX8yuu3y0vM/kYZbxT/dYPsM
BwDO4pULQP/u5tfGUpt5Kc14o+VcRrbCTMAFJf9U3du66bX1BFt/jygpcNKDutlP8G8ynDbJH9Yq
3cfGRNoIU96P8LfxsG1VobunlVPjLYgfiP+MxAiw0joUq+57b1VKPZsuUOvGvNmpKYlzMTT5N7Og
iix1QuIHoQRGUKs2lZIOEh8siDwKjpE6Tn0GfkBE0h/g22RGHiIVINwn1K9ZlCJMjnQtqgRytGaX
wbbipqVodso/gG2JtVYlWkhY0rsro9lEzzK2u+N4JS8/iokhwRGw7qpMUgvpRkKP06pNQbtqUEpW
+rivKJxtG3pgZEkhY2iG4TZlSN1FpoTEz5soEjZj6taSTovoBK4Qa8xji9i9qj1sg5VJpAOz2QeC
PoQ0fqoiXXb8tBhbKyNHLzqJaRZmpiHbIIM9wCOufpE0RfodzX84fgUAvzcsQU2XqR/Qot2zkcPX
wmxefadB594nvTA4vIOPDSU2ploWzNtNR5zpZWVb3Eg4bZi3jXkTql5NXNanoCIouHbcsfj2BXkg
TA7KmW2AG3q5h9M/fiBJv9OqSbKuPOJvdOVHEwN95LkoU0biSogTI7Yx4o1s28S5R7F19BZbK5KI
attNvaYdiAPoRsnJVTbXPzyeUOX4zCFpCQlKSnLgUY+qKp1wmB6LVS8nWE9UTLJoL/dN3yBKPJTg
O1I/rcLRwZzQyj3EOwUfwfdySVSEwetcGlq+fKiMVIOwVJIYsRJLSGgeBzkHEqQ7+rL0z+0lV6RP
MMOb5c/Pi0ycwfLSXO9NNIUbhh2CzJ7W93JsjA2pHQVIC8iL3pdGa3GjWZs9EsXiV1aY4DrPz+HZ
q82Kf+GUmKyfS467vO+5ivjfu7zus/5l0jdU8HsLZF21qh2PereC2qCf6rXKZu3HuXhY0Q7UIgfq
YVuKH42Le3sqqmkKYllSgq2Wi2NgDAx6YZBsCak5RFNhNVcTNuwkhOWImwjSNZNOhka8QMdkkWog
0jgsHtC4M9BT1BUYbBNUkc3YEUdthf4/EGcte0w0oLE0KP+QRGHoYDpezATBjkKpaC9dGFIyagPj
iWzOPNGj0Us6+A/NiiaUcAqn6Ja81zLPUNQFa4rg5tNnb51lussvDsIiZvlGFkBYrSTovBnEstY2
lzbdSDFVM/2EEkrzYd5wlLifGceeGLWjz0YdOyTxrSF1bOEIltuwS+C6L5CypmbS/dIK2o89zNbw
9zhVZTma8KuBlQplcDh4WlFwjkjxIL8Je9pQaxsgnbBP84rmEYvyTT3kAM5xM+xY18w6E6cYfB/r
mLzqgBejNqPwIrK8/crPpRNt83eVgxHdx8Az8G6ooT+pD3rYCxCVxhmN8pWrziv8AGxL6Cey6Kco
fDxuofFkyLZOUs0oHL8bg5VdmbU4BioM/MFO5hNAgnkLhkjUwxvE1iW8j0GbG/b/TLRDZIZpqV/P
Z/LDfQioIAppszVSlBC+wZ4sOu56TZ3/lKB8Xqnv4G/+JlwpZqDmmmJSe1R0e9Vik0tp6cRm03ZI
kF3v9/unIPHrgl8e5e+VFaY2KMsGcYjeMRFGN1aZ2Ll2XYpRSWTuy/wRkn6zkKrLBgn0CFynIPyv
mctVgovRKCmiEFxeI4ur9qHZ8ImGaD2Kagchfu1AkDz04mxIpbwb1Uyp+gskHL8jVstfZY13w6Sk
Aa8P+fdreXFHKmPt0BHygXZ6/+tIXd2K0oRfUZfIJKQpBvUugl/OyR6t1onbsz87IFzkmQreSKUt
dY5+bjQ06MW3SpEZNwkPoOwrgArAgFciZsrRZRXNYBmH0DtP2m2wSH7nuOhW/0Nb6c8FdCJ21Yrv
Twql0cHbTiKV/YA5CmHBCsnw8KdUJDO8cB5re0wf0YfyqEmXPWAt4qBc9sDI6/CA3LEvaKZdbikj
RgnL+RP4XzbwLwm4fWSzMnDLFf8oOfF9Q5zrsHB1MHoQX1uJ31jEpaTVh6Gn9qDaUv7LCOVKVliU
aTaFm6V2oKUQK7jjHSRy9VktL1k4hWAMfCkPZ38GKeG4S4JBWE7c+Jp/79vDC/geilcPTAv1XI9Q
Yp5O+jTVCFe6NuWBBXmd/CuHuxqs2s79vSj2yHL+DBWpvXSspo0CIU1O03dR7tcdEFCabNV+NB6G
lRADYLo9XAbvKk5YZGR+/9d4WAYSwQo2H4T6mNBWHAbGfkanEDEskFfARFQdEBbTQki2CRYrjUL5
A8lT6sXzHV10vPz1O1oR9Xo0ylIo7OBcv9S/iFFsMGfJd7qtX/DKYqfv9sl8FDoYLJAPL719Nt7S
KVpct+AZXenA9hhc6avr8GZafovDCfB66u1C+wZqLF2gJYs++VOMSyW7peDwO4TyTQ9KdLzCNjHY
LhRTS8y1LxRhwd5XdtgICP8kk772PjMn3dGGuXnAtKz8vp/yhdS4P1PxEmvQRhSfSuLGHZbWjjSY
9HngXqr2gmT+N6+7reHSej/GuXNof25coMmjeBktcKpxJKi5bUNWj5QSZyJviiXZdK+iQeS8v1Vc
x3/52qY+Z4ZYO6pXtMVwRCotAcCE25OPEmVGr0gQMYqGMp/pWTs+udnufyI1ArSSBSyq7D+IJse9
bk2FGwBGWld8Vmhl25EeuOymrYoftg38+B8MiokUgjekl43i5BFcNM87nQjOSKcDLAlnxKU3w3ej
qme9QYb5fLdoDeGYLUeujQFDCDUzRLQkZ/YXmdhx0xJ+Vo/yaVBlf2kz7FEnkEoE8wwXcBa41l2s
KzIQWf9aXlUWjgqKRk1KyfhcLk5Poq8mohWsB9spALK2LgXVThQqjHLLJPEz3FMxHhromJGc3tKh
5ZrQpAU1XJJ9rIB3364dBoRctgmNqfN0uS07qkZ28QSpXJ/ygYRcBDEdeEwb/ZLyxYllz+DwFI1I
kNbC9KrX/x21y/whva010sHwqYO0UbXxv1D+cEf1SaO6mPx6qeBoMxQA2hwAl+mFmFkhBuZ/gvga
vZBqrBJrZ1Z4BZA8bmJN3bKXgXEeV20A+KU3KbKe0OFSGEvNhaZlc78hiY2ab5eXIfRUPUs4JlWx
sGqnGX+TGEgFqcNNfimJOUZSjGVvMW4pQLF4RBjTkTpiEwhaIsp1h70zBBVoTSLt6+cp0NJU0RBd
BfmleSyQy35EP0jHRj/V8TL/9xSkQKeHKM5hOMJeYxsEGRX1TM0259cjqy5BPIQHDO+qOWlfPm13
aWVygUZZ92UAJW+ICpvyNoEfcBwpm3Iu3ytUoIJphLeSXAZWOI7ilMWjJ+ZYL9GzmP49oLutEtB9
vUwflQr/1RGDIY1oI91S/1Y4LuI8zVpqyIH60Ui7Q+6RcGm6gVeB23h5R2SOYyLFmavdZitCnu6Z
WZYc0kTWwzm2YJPuwYJv5dluOcc4a7dvm720HGx8rGnpvzMav/TjD93SoCF5PMKUN8/bvcxoO/oM
qKmFh7goerAkKxv6RkYP2OE4q/7/grSiiK6t+cMHL4beRSaWQ7VQ/agX+mYt7xUwPVa0fVgzEJia
eNhVcBOQuIR5XwlXue424oci/b9K2+IqMHej+swEXy/eV6EZYjCF2vmJVdXtwiVjx/1XYu4LDJXq
tCywyjNWCXjHvxboTG3tpIDaPc/4EguOA0uuXdLDkHkmfmk2su67BCGyrEre3ggB0Eu5ZONCzbvj
058ExSqSNRwEwuxJAjN5/zjUtfkKDiMr9LcKpIEz3AtVqtS3vGmtthK3L9n8HMfSuGoCu+07VfNN
z9Fx5IIYcGSCANIJWlErKHLk7cxChnzdW5xqpQXkc+mdCUF0F2hpogJogePD1ob7gxmPD9C5JI2o
ddEbNrD3BYXWhLgoaWVGx/BEQjF7eWR7G8/wBfh29bx13w7NWWoncmLCJ2TpZJ/3nB9BwhgGH/+/
V9+LZbQ0txFiyHZL5RGZzNoqn43jJbXvD43kfAkuBLx83OjFV9f6obAWCFqTjf8NOagMYVva2xpd
mZTMMD/kN7Rdq9aULRKBU2PklSArN/B647GC/zO/KnUy1Mu5dIGuxxBPOWMeoA21+N0s8lbivrS4
Jv08O3/logFusF2fCkkuC5jKFK5V9lfi5XPhxnQYvpcGQCIJ5+L9ryEpUG+adxpDKRbekVeQcAke
lKP1O8oMr1oCel8zYJisytSIZAGY/ObTpcnFXn4ohWBD9qNRtDJHMcYm6IASwrXfeoTbWoGfU7i4
xocqth+XCTs+SCrVo3fBh239HBdsSB3Jevcg8p1p0PREtcQq48WgiQ/IY3cVcOvyl+Dcq3wHGgCm
XXosSIilLCubIVBYkbgmAI2jf9PEtPa5BK6Xu1LYLo3fEcmU9eSYb1TywcMU21/jH1sxgl1WNWV4
mS6aTd7MHuE72ThhzPU1E908Pn7b3SwZ0MSif65GyLSSulYysgipglP5lq3J4lH6Nxy1RwEma7ke
vlKpSARzuyHgASfNK7usOy8zxhGtkcm98d4K+KoBsqu7H8SvykguGeXC0bXOA276ryV7Op1rhGj9
/VaGO11q2p4SGEnscm4c6PPYaWQWIbqe1YDvuKNOjkoZkMc1AbjxoHnji2N2YfzJNItbm4te8rgV
OiPxz7gmRsxahRu+5S/GvoGMttrjy4fqzg2P8FNlnkP/evLIEdeW4iwtdF7a+3YkqMcZufgaWueI
HAxpz+fNw+pYprPT/jPPOYnZ1t58hHyjPdvZ25KqXcTOBB7zr7jjHc8wXIwiYS+ZJq/2ppEL24iQ
OWstO7raZmNi2MLAgF5TkOxmhKhoRYo5s5eocJcXH7XD+dUykKjeYv6Jt3Th9cZ/Q/aaFOVMplGT
IFLHJ4nZjN5VuN+doePlQPgOZfaGa2XCq3Uug/OW0pm0nbPBcvymZkx7Ato1JV3X19sjAtncPvt6
vgp6i1yZMgcTKlhi6PQck+wQL2tUmMzeP4EZ+P3DwmAXuAZ5ZQApRy2DOZ2T6ELN3glG0s/7Y56y
eSpOyJvEflQ5Faitn5GSCinbWZFSDt6+nVMkNxftJSETDlMZs+e+3UzWN6vdUove9N0ccxdbWvLj
ULE36OZnpOH4h+G50FuepppTReQf/dzHX/VUpdCddR4o5uRPd3XqKxafTyS/HrDmwkg22BddO5l0
igvrb+RUMCnwtTcOOBOPNxBrNCTvZBNG+y1CUPinhHsvylU2iQVVC2UmTDjp9PjEmy8/V0sHcK96
Fcem0/KcwBCRWyBrqtb1v4QbEQPGrOcFXQT3PSwdi1+oMV1mwBjct947MKEdHxqPA8z3qg01p+ok
ZM+hRCbaBIUxlaz6gZadYdaIWKcVkdZTiWpUyC2/Q5jMu8sWN2qzk0xc0jhk9RZKJtcnxrSOYzkt
RIGp7kCUNuuHxgwHurGMiGNNzmDZjLKZHdWun/yaEI8U/LflGWZavSWq7I1EvLDtZL+ZJqnfQ237
0JQq4709V576J4JOHAsW9DLz4ffa1f6eKCFF+3bTDA7X6byc9n8KsUzEDnpUYK+whki1mYqn8V7s
QBXHBup5W05dC3y5JDBo/Ljb4aM1urau31S9ccJbmmu+J/ScDXACvqQ81eVXr3WF9cU/5Hi35+wT
XME5+4Fu+rXfeADdEzp2vcLFDDZn8qr2Bbd2EFOy+KsG12e5Tt34CaLF6QK3DovwiMyUN4h6A708
tKywKkAWIAM8DP8bhgtLZWeV1vi9LUA87aRtKeDiAEtVwvg6muWHqXYKr3fSh4lP9CCpBHMJRinb
h7szlix+1WWgzp2+2W249qwNOaua+GAfJQzYhW2DXCU3jJVI+EUFU/HLtJKqn2bmfEA6khhHGKuG
pz6w2x4dDlZNQaliIiiIYv1pyLLmmYifGnH7PXOn6hx0aPgT+tQPPIA+qikIErkMDBFnQnvgsit8
V2uWJpatNpJS77flD/+1Yhvpz/Xnt0uLRlCXi1S1wr+gn3XTHbaLwO4wwatU9zK0mpY/hDHPRV5Y
goRlX2pkyxh3EAOcc8H1eP1e4wByQSky7FiLckckjr9YM7Ga+hPtQzkWJm2s+6VdMgFod8RrSdmG
I/zWN/r1D3slY1w3AM/8boFF/43iL9yCxG4OFqhdbUEMsU5SOe1us/qXOZKq0JBMQ5/EZf0Cqz6R
IAXb7Vd93lbC/3caTanWWboY5B52RRBlfbuk2aR7ReXzBHa+K4eEgsWhBX7OJk/NvaXxuEQRvBTH
GynD0MRwMOsxBFKc9TDCie4UmTFovqRiOj5SCot+AycGJYzzuw/H+J0rXn7BQYw+zybNwd21V9yy
Q+S2LyyET+F62Kt3C/x69MparIo4OLNqkcqDuvwVGncoiCaLhc+12Ylc0r1wGT6xeXch7lMdOXuX
lIoP22vX8KN3U3gXPBZVkOgL0xZZk0hsbIbmf6XFVKj4ymp9HOp8hh4vOxyrmFnlJ951VG7Aysms
vtLoDm6yEx3cTnTEdCMrzvsfultn9B2nNq9rcj7eSMS/DOBMm5KrpIqrPXK/4Qn2gCuNnsf5YepP
wHleIj+S+IF5JGer6l6K99xlUbSlK43R/qIM0n3GRQETZ4SOLv4Cw0zs5ZPZF8ENBSLBtTqhg/Gg
Wn4Q+AK6a2V+KBZ0BT2VOyzNG5Bb1zSaycS+2B19Mb1ZZWPyIixkUkQ5fopJPJsFkBQ0FtMENVyz
t6nbSQszcF1uQ4qKdvkWhat71ZPKrbOOl6KrALRkB/xv45Maim7CqUdcaEPFHg7gqJcw97ObSH/x
LNOJaJOwkqA3WfPUamf9DqxYq135UQAWsvSZB25BqqPsgTK42OZDatRaDtIJ5AatRVOubI3DycPg
ICdzK48GH0RiXJICpHOwJ9vWJTZ5MGqRaDnnJgrxsCRYkYP7TG6B9fVyrSwLIi46RpKG/lhvkXvh
W9ISz8u99nawMllZkb6ekRe0Yzw0Wbl1lhlBcJ9YoubSesne1GOh0/9cnqtkFWuF/fyVW5QzBEZ7
iorI0mR8R3qp5I85ibXbtDO5IfzxUhqmk11iD0qJ4Sxgvrrcc2xS/PkwXjU7YXa34ORBuM5Zifg0
kZx9qLj70ujHilpIIjD5efxO2OwLVs7q9iRiLjQs0eVfa3xdlUL7DoWUdU/VOw/vg0fDKLbJncdk
BAUOFQa9Ae5gSVo6S9A+Du2TywovprTWjnQIjvsZq4q2sGy6jGxp9Pwg+XwmiwywiDyif4wj/l3I
qqGTiFtoYncuDDS1m874lLs4tg1mR1QNyqVon+1U2dCJkAETLjC8kK3/jZROFbNTUM8hljPaQZnC
TA0bM/4Q5Tusp8lOWEpPXi1d9pHLnCNDEZY1CYYEOY4Y+O5i1NnvDZVEWPlu+aUbXVIeO/0Pv/VN
EZRq+XeLbG+Euuu1xMF+SZVN4gMv3fJN17InSMQJ2gcjQOJwhnumhSUcfg1MJH2nn1MfSvHgQWy/
vFV5I0LRVy9AiqLu8h+V4sqR/MVEQwnmWjHzdc9igdXIUgOWwbuOmCXppcPYsUOteA8Kg6QaUYX/
x/8/NsFWSp1m1DIrZ2PNgeX4AVG5OeHtFOFxh3rjcwj+OS+ZzVOrLWtYWTRBjmK+O7fwumeZAh41
68iVWtnCwP9Xb/ThmFlFZD/AUDLrLu/72XK4mOlGMWp/f+s1YlH0VGfo0kP43gAPaSiJA8Ec0j2U
JLRvrONL10JeXVHCtYC4I+LFYADjXzrFm8pLDw/HkHRu28TK/YQ9iFYiYqH9/WhTHZ263SphG0Gj
GVqyVkN94LWlecbZAStdolcDlQ2twGQ/G8G8LyS+S0fqrFAYTlADTjPP3fhyI18C5Cz4GqoPBECd
mdeaB6Z7SmpDgcSSp5G8yS9cXx1H1OvvxwXAdwz6mN2FehZeuhuGpi2CREe0rmyySgkqNKRsi3Mo
4y97g/gL645DtcJwAQx9GKx89FIXno7+OH5r9TqeSPJblL0sE5BugXQhpo0iW3U69AavYp+SlJH/
9tfuRQcTfaPq/dqdZPLMTkqORXYD73xtlNNOwNr98RlU1Ns7B4kizJbCbfbnPralQ2RlF/TEA5o0
eVbB2Juxdc/itODOrqbEDsaGipXDEYbN7tYxjhqpJQCuZ9NOIL94QjL5j9EBPYwaEKrOSvLr1HV2
JOHFGRWpNfcoqLSmMHd6r1m4Ap74liyJSMgakMY92u0K580xmcjYbP/Bndh5kSAtE1duTfi+nn+D
G4itVyx/1ip1+gkLFAiKV9J0o9Ovk3FfTz/HZzuvbdU16AOQpCAsRKMUde3IQRO29CiFsDVbw9uz
JMUT17IrPtjoIB/gRV2w8nMBKYrrYqsmLQA8nyfhM6eptkjG0AERz1wbTfox0FlBLtevyKBtvk9D
jmxGb3Y0VwnjxzwXl/pWpLEcKnYV5Z+bfJ6KtNoh0BADgiWI5b8XWb+2SCC9TX6eFTKsx/IZLVcs
lXcZAqGJX+JZh1t1dvN7CHJbcydqSEaOoYkAeVBdVTOkQQTuw1IQtUglmxQAEofxs6gS7gVLUIEz
yxezXvN14EA0DnBC2Eg/wCuIbYfiGDzUcECl5VGZwO+RnbQhnrnLtKUxmnIqaq9Xw8za+SyFctx6
hJbcLVIawvAWhE62tVHyUI9Tflm+ARnd++ANpuB0JBM/2Ti2eb21RENykZSoHSH0ZETuINMjXYjy
H+/oWYX+EikRZ4AEqtq2Ld2rO7SB3xobEZyYIizj65hQ3i15lSqEN1QVkrhzH30/+eTfwjzTwx83
ykblVITeyDW4zcSEv92IRQDfG8K25qwemNMOXlL1Ewu/X2WCKBxMxG34KLVln/zwmuVosdld7JQW
x2hz0WmJF8MGqCbK3OYdlq/ttfSgx2wKxv2AN4nuR4GeH8cOG3A0nTDW4LLQBF+QFOFZZP7pqAHQ
VqY6GvfJCnm/tbIRwUsOpzlVAEuBoHbav2ixAdT0JTzvoq6tOEFV9+kI/PFeDO2IJr+w+aF4jask
zLD06/rJDRXiFtplD51A2W8UbZQWDyd2zKzU2vJ/k8W+XdEmtWRBZFgJcEYjwKCzcEzFMyjC6C4R
Im/VAvJh61Z1/cbRP+qPi+EUnxRsrMxpPgaCzu+MLp4k39j2eKYSvzxZSJlKHawtWwXMpULP5Iz1
Mf5UGbhHuzXn2Ems4bSISI/P7jZfd4FRlOZDDepmz0n9QWHhhPiPR/rJq+wWXm24ZfP8CsmB55ZS
nxUa2sPQd2ksiCUXrrCNZ+Rpx5aSY2Jzg0mLRKRAU0IqDndxAjePNN6T21SAhf/iTi7/kAvH9AAl
ksVKhicn4hB55Aslts8LZ9I4euJnht0UeknNnm9iTprzkIMlPKO21vCh7qN1p9NyJCxcSKdJJCrS
z2OmCZ2vInbRQnu/mjOrLw8nwACSy+zVLUQXn/I06UX5uZPSCVGZIYwVdRlgmaUg7LatE/HzYepb
/N7IFJPfLoSOlJbEx7jicImzfHauSOr+a1WBQ90mLnIvLZNOlqDghdXmiqZze3eqQ73ZJCJc7rF+
TZ33glD3bPeVIK2HSI6xk+cSBy8sNrPee/1LIX3wREgKKsXvnArhyl3seiK7nQOTwrcnZv0lfHGk
+/21uAHSNID2N5H4DcNMDFTwzni4sCGwcWhr90HzT2YDgX1CzUDB8YyDmGcD9DZIyttksU7D3b7Q
AeU/Yrji43r477VKQY/9Hc3wkZ3iy+q/W8yTkOnlKnUTNMhMsB2RZ4zWV6VCPHjVeA95I/9N8F0v
ppybCijG9I20gjedx5IE//CI4tvNTINS1aF/2xtLNsvsw3EnaHL4eFO/aV14nYuUBl+qQrHqjE0S
tYEtbE28Ui0ZhNv+f8fZCwstq0OpyENAtxA9X9UcoO5/dAW1sr1aFojda1OXGnJjfsTs4/C+LHXT
t3icjLhl+LNjbviL/YBDCIadqUdpgf7MieEmJqRXD7L4ov+ljkhMgJA9CbytgzcgefhbIjEpOhig
hU3RjRWmOOiTxLu3SPuJJMBekeXubl2/nTcFYQjuKLLy5vZEJ/ADtYstEBvSHfWm0bzfhBwfMtzi
G5RAzPzYEE7icHFNxvAaU7YAj+1XtHCZg+d5EEcxSBf4KZ7SKscKKjfHggFfNs6jIyJQ3cF4nvHM
q68nzSykTzH5wnKZxrxnCeceGnSrWKjDfnI7CaOmqoOfBQogTjzvuY0b48rnYbTezt8iR3zClI/t
8V2tNXd7EROz+fiIJQt+2lnEH7IOOmAmOneUpz5XOMtxQ9EHrHdkT4ZMzyA5LcnhNjhIJ85l3D2+
xnjL8OxuwJeHh6oKqmuurNOqZS9trvXHSmwh0HjTgXmOTwrSl6eDHGCtGwu+Jlt+diwkwMzkAEHD
Hqwx9XB7i0GPSd7gy2xmhk3G7ltuGxrMwPUFw7qTUnZX+vsRWIkVOW6S78BQOXX5MQX9NCccSdIl
Tlhu5A0jYFf97ZcxkWUIxyBEIN8PUZb/Mw3gzrXL2fRlxANEV07iKs+tYReTc2YUjPtleVh3RXaf
SkIefHlKg//ZLur4SLQBacYD/4Vy+9jvzr4WbAtC/aDjYLUs4QDwhGDsaKX9w6MMdUONp4CojXv4
lgfowlX2dBsaw6fZ71JGtgAWeWlNO/2P3PuExDFPQbEyMAxSN9lHbcFzo9ub7+2CBioDm0OQOXdC
8VWfIkGfCoPWPmcdX6hCapDPGgIvjl50vX20belKTvQleD+y+t9xcJPNCWCCETbZ46rH30gs+Ybw
EXwViOlSXPgpk2NNOrXQn2CAnHpGAlexW+HYE9HoOYswUUnkbcBokESOO+u0Vfj/M3HaCre3R1Tw
CN4EL7utSzX5hdzE+uNtGbqUGmhrZSvPp+3yB5JQByXUcjRZS2JwaqHGcLJckdtExwHKpa9+s75Q
8nR6OpKbXkyxywIYUW3Cpf9/joCVnhmMcY5Gm3JfeNl3hKqiDempDbEbvUnGJqHcAPwDsJPenaOw
5WOdZqIqiQUtUPFiersosbiib2Ae433UiqlPIMSfbZxyqHv1ch/73h580m3Ga+Lp62GMgaiWi6RC
p3M6ILx7BnxhjXYOqTLYzjGQVmwgNw2ZVj19abp2iHkdDOQYAYRVN8xWMr6FIcKwVAutVI+qdwLU
KCWk0ZoHhQCm84AZ3UsZ8o7d008J4+8MeN05jJqLfPrip8D60pJPSeBV9onUPmRDSsBj9TvJ93wO
j0Ot/KKxrKbRsekhbe9pr9kvNiYjjAqGrlSzXWtlOyaXBgNv+WdUDK2KVWALB0jC1FT8A42jMcuy
9WN2dZDlaKr6rv9o3/Y/A3hxnnPd1XIRAEhljokoLfCuqHdARDrbxWKcYOksXr8wGJQSpe9+VIN5
RR0AaWe9kaKh3yyjZb46BsaQEiQAicslPDPB1obd9IPK8boI+yBj3F0/ojE/Xtx9l/qqBaLFG1sY
ufyjw+jNgJE90qSwhT4H2sgMPyk3SPi4KeelEouY1IU7aqiuyicTq8Nl1y3dX9G/NFpI5WZwB+os
CLn7I2836xAXbn6vpquXxA0xo5tfkfWL5HywDxc+3DRqYoGU9NPZI+djb1FG6I+DsGfQg/B07IbY
XGomuiZ4UHtwmyM0fQnEIo6zfXeWVF0BXfsJR4BepCjvYyA+qtW78kiInv6/2kMt7DnZdOXiDS7M
l9WZmJTV0zKM3RkaY8TY3SsvkRp2YzZCX9ugMEyURO89Qu8uJd0FxZZKh5ngh4W7FFMVqKL2GzkD
SVNs2S+kYHM+UKoCQu/77J6QSYA0EoOi6YxezqB39l/eUtpNJN1LvzMTXmhjmrV/cP+Q3NcUWZwt
X/FI06mcU4p18t0fAPscEOS+byi9olGTEdwXhQQFP7h0m248Sbhg1bAIcGRFVwTBw95UxSVuXfhJ
fQIyrWnpyT0lEKZp6bjVmXhvYjCcwBWI9+7TVBGEgwEiQlaqmbVldktj11A5BPkiRigDCfkfYTTq
+UJgCRxnSCOPuAwWli+Zwpm9YAx3wPqI9pjXk3UyZ9wXpaYhZ1FMJwos+l98FTCO8Yi7eECqJF3a
p1mcRCtZMi9Tf0flZdfg6QLbKoIsdF8qLvBXTaiLssAUISYxcy9elxbPQfuBQOLuqYVzlp+eX1bT
tdeeOPUQ3qA8KCVWDlNj9soh+GPI3AC2YvM3IjGRDcIh+f1TYBFX5H/IXAZ68HezH+Qj+FCzHMCR
aIq29KdXazQ8HMBIveke5kkNvcEJXi8BqWZWbA1BpudyoolnhlWMLAGWU1ZFO4OzxZOL4qFQoeCi
84C2RYasF/8qUwYMT++Nn4201u93okOXcdDU4F9La3oJUoRxEalt0u2ktmTNdPwqGWroUzviHAs8
PxDKRcks5p70U76CUi6cTPj9cxCkb8JchwPHxJ/sqqH3aw7iUV9Hb6bmjcTnXu7xBEVH6aBbSPvg
dZ6t1wVGDo//Xlm1obMI5+Qu62wOAVRoYp1ujF94AzXWc5nxCkK8N4/D16zqCtEcklob4k7WakWD
XoJRX7C50chFDDB/dfh78BCM33Gvw6gTbQH/aTp85fE+ub/Nl/QTlCrUdtChIj4dRaVnzZemXl2a
ARcEcn4kvjVhTqRT6xy+6la8l+qJQ7L3KtZr3vxlypwTPuKqBqsxhEYWUVpnSUwzgWZ0EfDhrosi
DckyAx0pef7AKn72kgs/h3Kp+XnsegmR02gCk9aWm641P3K9rRCnXPTnF7wrGhmZ1BF0G+QRM+oY
jkf0R3qZyeESKXOxD2onMuLi2XdUA7sKcw3NK8anNU07q+FL6Qxb+200glpSCESevG+J0WDlUYb0
LfHLIx8G5uz1o45X0TDNPEOEqu24q06rdF4+xMBki6b8UhKL5ZXIX7JeDBghhy9Iatvru0QH9cXL
uyO32sT+R7exiMWe8AsMmb304s7Ej3VmikcBVH63iie4QoO8JEBGAkF14Gne3N285rqgqUhnUlH/
FFJMHBNIin/m+Ra35mlc0ZydQ2rhdy1WfvwJ36cR1K8K/dEuDv27bhBqSl7UU5R/c8NbTzrHrYpH
HFsRuNKOA0/sjgLSa2lVXGEcdIHaCc/DEYXr0yLy7dQAtt32xnF6UkyaiRLrjb/kV4m6ifNG4p6B
HrRWSiU12ZymGKXng8/LoH/cTmUwXAToTG/uQchMPpYEPVoOCCOJSEVdSMszZgIp3S46krVWCJ9P
ANIjgUCOiApfFez2/s+SfzwSfICagP0ESywZ/9O9gh2Cz8eML7otCPd5ZsN4jmNSXZ78TpZSFEFY
CJf5s2osTpYKqQQV12zCnmKR0JQFlkjeG853oTRj4fwTfo52SDHFlFBpq7t++Gg2y6qtxEXChOeF
yjiPlzXaDFIMtA4BA+akpr3f7bEwqCcPM7Y/ijTH5xYoKnagZRjqNmWtBi35EiS90y5Ukbgne314
YGfar8ZT5T8YaAfFlJbn+EUPnoWFX6z0vUpZDKx6Nszk8GF5ODoD+lohTpUetZRvNU25W7aiPcxR
RvdPGedUdGMEjdurEKcn8NhSRJYjFTq3P4QbmenKMi+FLYw0nfTIMkv7wHXu8ozEKTUe7HPL4uPQ
4J4jolpuzo4YqPkwclKKjlah9S4EVfZP/5j/DkVvwvs5rCwjwQwdEEosduw77YCNRcgTjSxqPy3f
YNfq1DGvcZpVdAFJ8Z1EpUFr2gRE9Tph3ib6cWrS5ME9PI/qo235zWEpRL74e8hxzZXRV6Hmsctp
6obsfQYUNV8CDyIWptWQgAh5YYV6RB+toysoj5dGxVHsRRbGmSrxsFvOkJIAwrwHKUbb9SwvyD48
FPG2jTBX7INp63zli7Ehrla801Ml21xum4A0yAopt2XoyCBC7zQY6bWwsb88R2g1TptwgkwYiRw0
o2lJLUoZ5wAhAstDilYaQ84py32kJhkJS2i4vTZlal048jBp1qZRLbyi+LRvlMVmR/Ysk6wRSKR8
vp0apYLfK26c06lPI6wGcNzy9H2U1x9GtYBtHywNFtXliU8xu/05kwGAI2XKJ1cFgACBWhPa/WmI
VZuGM98nH5cK/lduV2tyT6cPPGsVJKFKA0xEeBi1kqFp+dqBmbQ34qX/ndRZYMDSFhgItBL0bbf/
1s4/TJgyFCgfMkY++PFvgnlkLH3UVtoJaC/Zj351szzoNoAJXhJ+pU+FdD/x3Wu+UQE1qbj99T5A
sIuy+p3Y5KTP7Xlmb3V0+8igRf1YUZhRJpC/I3ndCjUggFJbQ+3fZ89HrqmKGgMSwZSzyWOhPcPP
856pLiNFDHyW6HLEgywshN5ON1It7UwDwm5H67MVOSdZGxPB616L2QtlYZyleSRJqCJMgGU/E92c
yPk54JEkx+Z/WqWUget35mJUPhLUMZdzIxCdF2c5SVvuQ8ltdojaVs/qG+XGZ21KRYFX3npeZoSx
zXIRfp1zrq3DmFvP07HxDwP7ouqVeB+JWpIEnbRsdjXwVVmL1vQfKwBgCLqzqTXfvbOWmLHABh4X
Vg7cmM2hiIhyktKZ0IMB7EyGbrVYcFu+jSrW/dLimJNJ6BAmB2VCUm3FLrR8JS4GqlMR0x49QUCS
4IDtS/orKT2vfVVGhZbeByLfh6BvR9E3OTvBwPEgJy1yZcFgd5AKaDCMfnisosbYDg1kH508G4TE
qind679AuowQE8UpHyPKjvSpxQxba39gE3GG/khoxDJHlS5U/pTuqwXB8mBUl6K6wwwxUhlZ6Y6L
yN/x4m1SF0P7E7e205CARhoQm/vxK3gBLeJetRAxqhHcsjuYjChw3uihmZtWZ8icU1aUIZP/N6zg
oxuqqUyM6CIIwuBfHD8Zgz+bLL696Agz+5rR4lY4wkhVE+Gtv3dmMOlwOtwIzlCGYJl2M6rQv+yD
WL/3Cb+sUOyUOtTVTRQPXFYGoqY2mdxPy7r3yUc3hRIsHzoKzIRlHfWsK2lVpefW6uKfTD4iq4C9
pwtNoE7CxrhtIx9mQYp8zKdkXvSjekDrStop4itgNzgEZr9s3GKRd18ffPC6j7RuV0kOYsDf0oFT
MoNH8IAdX8OeRE96aWRk9RGUlSNlbHAQlA+W5JxKvlk6Oi/7lJxhxseMXhvU6T+9shENLHMPZw6q
8KQr5va7Rr7x8lu2i4rExZmkUh6JSnKeDkyIEd4a6GEW8BC6iixuy8PimuhD6JyPqNRSu/UkZt6r
EHshqhxILAa5uYQwgFO6MDOMCnMbLLTl9EXONdi/mNiR2TzElo/uCbXcCekoZkzjgixV9P43746P
QOmyYMY7LPYFMWY3UYGlx0mmXndEwMISoQawDroHWZFHSiHrizptbhj/Mk+IyRO6T840VESfRCYn
PMKrRnCNolZySFbHe+qzYsy8JNvsCXcBC9rSDwk6r9rvuvpcvYnHITv7sTJk+YPMAP3m6ogozr6f
Kn9zEF9Asvt4PU1anI53rgst7ugdLFw9c9/u/xjx6hAo1fX1bdzA2viEkUuvnciR1lP8lD15Aux7
ZUA/BB6gRkMhYO9rBWPmaLlRATcHnIH5evgnq+lvxUYIx5imKe3FasghVU2by6pkUoIf7GAAMMnF
yPVG1as0/TRWOalZSftBGlSJlJCq3he0jTR2S5yA+klFcqSNH6nZymhe7xjvJUAsgVYO/ebMuqlb
zQlkcGmHt4N/lr6BKzxwzS3basvbU4TvsXRViW3sC0Jiu6KWo8dkW48LMmoaM6dpiNompB8XTKO4
L4rdvk2r1EY+gzNtL0AYAo1+BDLkIwqfuwoltEF0eGBI8gHKnlEsem8naZwUWTy+bQXkUlJ4dRt6
/lAY0ZzV6At/R+J/sbRGbrUkJF9BbQrkzDPOy/QpUWa5R6ZFa/JHDYs+7P2gpG33OIQ8i7B+Qtfc
FdmHULp4RLTZ/+Y8J81yshTt2ENYbJzMRKsUUpTPup540PJxSPwR2yBJj98lN3Op/CxqeTNFvfSi
rMAW6p3ADPedI8XSGyctz0h64itNIg9ZpvRkGYbjG9ukIn4QsTNs/KPTwAW+hLA+Osbtcoqsn14+
O5gn+xgOOXqotWI9smq0S1vIDb6+v39n8Ays7FOmNAw2X9Ql80/2JwtB4Qe2mzEobgUGkzP5d/8R
emaKydTGh3BOZOjDQKLDT5Qmb6wWv6dEe74I5GRPGY6koVhbQR4MhP/f5222cenhnNPPt4N+0VVR
1cpu+RzMGfIPQOUQcynZzNUEw0eaKaGSglY2o+iYSq4ABo61oxtMd/NWNi+htaVGtYjyWNQTLwHG
DoF/FQYGPc9vuYFBktXk63jyBG9vbd9kbSPBCHZAnfunRr0+vb+U/unHQ8qygR0TDbTYPaCCxUi/
6rI8KlblpHNi1WazR9sxCtcf+kp1WqjBiy/k60qwfqNpBsSQSeWg3bvicqnqXKuTMod0/GAwZBQH
mCbn2IWGD+qqS+xh0lVC/CKwjtOTjnifq34MMD9v2bz5b+ldW3VMdtCwyedRDTaWsj8uMr6jlooH
31u3ptrd7S5a17P4cGFywuyTJ/Okzv/zZDqgTC48nDdlVuEDp45ET2yKCjLeMduKHWex/onbo1XC
Ng9yPsgxEacuhg82WWhlvwKsPgG+gCoIi6RoiW42I5D+GXFRy2mN1IxwYiarTL98DPub5YpiLcf/
scmxpvtVMKKxzU6dKUIlml8/dHD/leeEX1Ee0nNyIIZxB88T0VYmYSucchsJK06C4GCB1KSlk/nK
M3cHHP/SIanGwzUA6dDG/lMBma5nar6gbJDRqkdnaFE7BPOlu6fkFZZSq3R7VZg/Bck/vf+T4RpW
sDM1jIPMieGmSMeVKBDFHBJHJwU0A1FWdrNIWFGlRYDu74PdysFGr2GJlj9J3L/4Jao4h34TlC4A
sgKUjCoAes71QEde8ujFUx9NlHZRZDcZD3TEFIYHnAa19voruJ6KFYiZfxCXNCEmakuZ/93ZGx4Q
jST3sYdxWaN9Vgzpt0G/VQtjfelOK2DeTo6x/O5xUpX9MmFe+HqvLKZTytK7Ra5Tiq3w8j//58LW
eS14N4jgGJm5i8L9dJtUtA8NVWUDGI4Pov9VmcGxiiX3IlQEDfkhIWIw77QDymGwzDcBCF+tnnLe
LmqLZD+bdT393w1kUavR6EnQSLF7+CjZCyxhELn8ryl3USGSAuKTYXUgKIrtr3RzYUS5li5+Pxh5
mUlXA2eIchl/gm9H+PJK1bq8oPWsk3w05usI+BUC+EFJ2eU9UASUx1iTTP6eaqTlAyugGInlvBJL
5tuD7YIIKhQjZiAwv7xWLxFjzZdOtMUoWUD/Kn0UAIx6XmWxZAmRm6hieykiyAwOHO3OQ+qC1BkO
p61bTcIdTWnfJR2W4J2kl1fV4g/qMxTg9mxv9kci2jaK18Tn54icPtWtbShJ+Ug0EEB+3G5ZoKzl
xKK8Cnglm/cuBhwZ+CH/VICkafPdImb8ZYUjI5/4O+Ny8S07tfeRz1Mei696ji3rHbwFNoFFHxOp
caAB972kFO0L5p1sqywko9Tjf65tFgTmjbQ7G7hSBzrb1sk8hTRFbxaiF3+RCqYcIDlrBj4UsxNh
Jzps1JRyyU6uaq/tJnEYPmrW2TN67OwIWVKlhI9ZRkWTtynDM4Ivvw405aelUtZxZdUTzcWd6qos
AJZB8LT68FNWU4qvGmEAKsWerAOg7CSFIu/qqKr8ZGKl++tuNZToymL2xV30Ko5ujUlBM2+XmrtU
IThij7RoFxfgeeXwAEzb9ayftBzv2gorIfCMdJun+MjUwZkNVQSab2P58o/AHkfsoTDvG6+ODT/A
4FcY+oWEzGIcRvQl26AUmV16tGWv8FLOL4Kxi3b81Pk0EZy9ObhZBN7ohGTbEVF2iXjMCGxafCO/
C+wp5ULkV/Nkk0IIIYdaTR/XltOXPnBaWH3UKMAvAfw2fXJ/dpuFEhgm3K7zHf1PrZvwhUVf54Se
FFMxyI64o/cqhZ9H1nE2186sATLg2lmFAlVjJKnrU2s5hwwgY5ODc4Q2KStX5cyyW8EsN7pB0Ojv
oFv6y6UywqXDHXfcIPgUtSO1W/warVjiNoWQtPcb58+J6U9qDs4eUGYOzD3I4XmFrnYe7CElQwya
QtuEseZ5VUn10IYZ1/q/+qmWfixECPao8zWBVqbd+IK1wRKPtCoX8AVvqQ3o5jMjavZkm28JVldE
ak5tiLemTImwBNRLdgHKIgIfh3sAzKKlFmW0w497ntiEe6NvBY+KDfyRv+jEnvR/GzaFar1UNb6f
Hb0nAyY/wjO4HIbSSgPxFGVYWQIN+Pi8F56T3uc7/lPrjwJqFjk2tHL2reE+sVL3fb0KtzbgUZEc
x1vHxfgAH19w7zJkdUpN+F9+uE0WBnMvBp4VggCGAoO0RGdYMSyfqRzHj4R+RHqpRHhy5B4iNLFk
vm9QhKP08xlhxwbFzkJ4XAWjwHEwvPjAfWT+rTkmpRcUCXMlGQbDHotGxZ0QdEeB/yE5/lzYUNGK
HGrX1BX8sj8XrF53XYWPcEIH8F0fQeyK3h5VOTcQ9Mu9X36nBq0S/dABmnV92F/ZLS+h8XmX0JMF
JgW89HletRp2HydBMOZBZG3j92NcMWRfLWmg82vuL0eLz9DVjlg7cdJNhDY3GQhdpk1afHxGCC0T
AYSBqqY6TpB7Q9b/89YirDF0+v/8FWD9LTj2e9xmnq4QMWVbCAvRxQN4m2e9hwZBN/Ck6dUS6HgR
E8e9eeU8mfXDYSrqjGOL9uc3UZdJaP06LUIONrKWscCsLkYAIYYX2sw+DzIyYLXqVdjQhm+Aj/eJ
di0m6vZ9ThNo4Pqc+X09WTwE974NHlMtl5nrAshd/D94gAu9KMcCDwhzHRg6V4Mt1Hc0P9nmIi2y
au0dUph7sFdvHD+J2YyIrNlgioULvn6pcxb0RtLx9wSrWwK3wV3G0dDwkFrte7XAkm2P+KCVt4G4
ywIOgMO/Yt26U0pyNWnxhatXT6O+I/DPiG1sAp/nUOBxiNApLm2LKs8D55Xnd7WtSFjkJpv0gprG
LFVlDJvY4sj3luE/sRqtr438lhxR0H/BSwZmoFC3Sss3VIJ7jRla/rWKeD2oJH7wYf46VjE3/VuL
sEMqi2D3YHVkk67WU5wIiK5ebteul2zixCNMw9bR2mm1xNR9oY8SsvQ7c3E+YPeJUppex/Q8Gspz
T0Z3VC9P4Nz5XvGLRHhzGOG9Wr46CV7OGvNsx9m3QZF8yXOK0sZjjyuZkGDfLlWqpwqVa91MLezt
QDgyOh06nJsUZJ+G9Xdpv8TXv5/fopzR07iPfLGmhIQjsnOvqbry9y8Z499P12CMETGZ9fidle10
NgSF7T1+Icpp4EedI+dqH0s3BQ6974QuewXx7xMjbOM9fTV2gP5078SQEgFmD19Ehgp4i/SiuWFT
+OvbD2B3q5BRK7RLyFWM8jMUxocL38TnAbaqTrJLW16gUkNnxj+HfhhRJV7FB8pbgof6fbpW5WpR
fE+FRQrq84n2aciuTrL+ZRhbQlNpnt9d3jyYgkdx5G4Yv0wgZMM6J3leSpHCB+qY2NJBM4mR+tWx
BmkRBPZX45hn90nBBNa+8+RtxW87n1YvmetQ1gMwfxUikE7ihRnZzCF9uIfU7ERtZ6hexAVOeJIN
rgJKArpREFPbSepychh8C3Y5yknrw7fXQjtwXd+FXtieMiWWK6efllBXRD0lvfQ3gR+fJP55j98I
rO4we87SES9mtIIia82p8tF0N+au71qhHEzbTV7ZXggmoWnhT62eHtFIcXWg67qgT5l/TivZOMfT
xPsHcSQ65seyCiCTyvpO3yVy2SXaMmi8ArGrDiU7bbkmax3UPQKsd26PMCBMxonr0d8kd28AlEDo
mbqAh829UrTRkJwuA/hzkOiZG/outG5IFP05taKnAYrVPXzAQrCalGZI1aOFqFUZN/9mZsKkZ+2S
aqEyTMCM5ucE7wrWQmCUewsEMFxyo5pJFsBc9kXK6fYlC9bMfSzTzTvQNJMAjzrWS6yCjk3AdxLn
zqlXeSlADmP12EYOAmBDflQLCahO+lEKH0edCdLJiFMNx8k6lea3pmUCs5e6Ly6lQ3Eim+LBUmeB
f7U8L4DyScpj0JnNITNbFdY5okL3c2kHWsuV1m0aKCLLXwIsbuoeaDDEVZOS96iCfWqmY2FyHxx1
ixxC3GsZqDb0erTxJts97F9Fbx19+G7ZJxpY42J2I2TiJBYlyJNxIhEjvFujm6rvyYFbObBNGbNd
8gCIXE2VcSkSShUDx7aSNls5ybW60CXesFcdr3U6MrchA1I5+7hgQj9gp8Y3bhP81AJ9SwtwSTS1
lIyUkRRoqUS411xj2xiBmSZbjSBl7OUzwm0DTXqmufW2LlzSJfJ+/u6BU6cYKf23yZDljQv5Da2+
jARB9Rkp3i5j74ghA0x3awt/1vTzVZG8c11zQ6O294Y431ri6VFhQr3xXs9GLQKjamDtY45kNBHG
TO1dgpx/aeYj82aFuMCibrust1Kg4IG9Ov3TyI7ON9Mi/9gY5fHZBeZbxwvwDNrV8HfuOb4s6hvi
DisQrp/fT/JUySBELtDPD1iDWtZKNLMI1cEXU3Y+Gv8w6fCVo1AGqJol7wDrNHEi4/V8sBjjn+Ex
dg10CrdY4XL7watZ9f0IbPeOP9maUIa6GZkIKthvN3ie27CoYASoFXrI09PfrzIWAe5N4Swu5GtK
iQAHaHRvFCn2dY7TCX0tZ5X9eb4ONGKHcbrQUi7jpDqReGTMM9+5YgDqeFlNF+mJJkOzTb95qXQB
PbF4aztVQw+s6PD6GqFcrHDK0kZK02UVnwlIPpmw2ecjoKm/jVECxLUGTuBu0kXbhuNWaqftmSEX
l1VuvMXBAq+yjH7sdF0gmmGOPligc4HWX/IxvFFfsfHl1D7HCT1uTB4sGxQ6fpYW7dxcMRO7HnAf
wfwJIGeR/MmxMtsWXaGVvV+6qij7/HYl7L2HjL7sgUsEVgrcxD7QkTJCvA2DWrA5r4Zuu2zpIqvf
XAjdqgdFz2MLqpM+r0faeE3+WnW7R29siceaadL6j/PqbPEap0Te5BNBQFaJ0W52M/4UaX0j1vzk
MKHqZySEYBW6iS2ybugp1ZEalJCRc+64v/B/ZxD8KQJ4LLPGA0sh1KKaGEpVKgRGpUU0c6OhjXoy
ofo9QdU625d3Yz7u5U0/MjAIREHitCedO5l0OpvJjimf3Q6sxXGxPn2dhQMCErf0x0u/XX3PoVrr
gfoARmMoxK10ufQqnvujekoJEQ3VM2WxVZijStukzcuWRBnbxwScDtvP1BJxDeMgK1s6+FHUphXO
m1CjJ9RmQiNs7iXpoLFMc5uzvN9M9yf+cBEX68e0A1NyeaFVWMd793+i9ywq5f6Xf1YEyYqzjHqz
3kDrJw2ZkekSOEXfcjgml+LdGt4WNTS71tD0/OtasU9bhgdKVvLjck4hQUoKAl5UfDVq0EoID8We
beRf5068SfKx+eqLHsQ99mEwUd1KLNAXQgWyOabEPTOrMBMXXv9VWcbzY5043UuFUWAeErzabNfO
UPoIQXp8mWLQJOI/U9YJZdaEMA18Ys91QUURKG3Nrf8N+wZV5uAP/XgWf0ZIXps7bwU/UI8kXf9E
3qACXuPJz6m2nkY124kaOmHN0K8pv71SMw/ISUm5tc/am023SZrgBz5t4OsEtf5KGreYsJ7X6574
MNH5OGMRSV/+bxLZdRb/YKnjfNK+MlrFRRIXU8Ufl2yscVgRfdbI6cz2zT7/aAff53thqVc3Txrx
IQqm99Uju6PzvlA9QlfENOelhjtFINBp3KiAkFCpffKf8dyumAieXZiXjxF6S7aO6UQEStvhqOel
pInqOf/Qd16nhz8pc9ExLuy5rh3yDPVEUm40fcGZoQ/IPSb/GeNsigZ4izlP7Ij2W77U4P4enOkg
ffSzfCgYT6/o2r0hk3AiPWafRNdteg0mZOhhVkgCcYSGbcSH2XBLt5yY3LyOMY93RJSxDG0PSEKM
SDklMVShE4Cyp/ERcF2tnAQs7IJY8ZaDZ79sOWlrtYSse0i4O3x/ik0xHatTRrWSAKclKtTLkBNS
hDrKu5pBcDZTcayGnSXKRA21pYC48YTbDubp/hM6reWFjV1A0ILQHUEd3xLTPCNi9XeXJHV1G9Hy
MRG2lRlWyqcLiJmXdXJepFx1PlDQ/aHEdfFjKLtZ+fQWrqXtuov0H50IHwZHcSPEI4KRZ9xqRjk0
0E5HyZS3psmO0q0byJpiBhwyWW9hFPwMwZeP7hLLRCChbm1WOxSUDdHSvfAtP25RuxqcrETqXLU3
chhZQ7Vac3F0t338gi2gALBRDioe9YYKIdbEf7XU2cA02Xh8fgR66u6XJyBU4hfMQKjepmKr+6Ka
cJTtNHnXJYUQJ6gMM+rPIoDYvGM7oQj7zWii2e05VekFN1MMf3FMjbYY60RPPBvIVtTvIeWg8agw
oJopBUcQqcshI1Ckww3khkBHsW61CbdKWfxTlQ5pUGmkljawpjRPRs+BQPzDXd/yoKrR2RADy+4l
ehZeyM8IX7LSSyHgnjL8Vi1Sjo61S1hd/W9dzz/Q1fUG0saXM5rD3bapsiN3pgOAainnOtruSK0Z
2qBpFPL88mIq5mPa4W2sop8FqntgLhrmT1w5j74nSSkD00bI4bBfuboYr8Cqyxbq7vQyAkRscybo
Dn1YHb/0UE7O5k/+B4VIoNyqRcjz97iGi/0cJO3X/3OCk5+llUhVkKcy72Nr9WDI/h92xeK5qw3M
cd538f3yJagwEHRFHMdDG8AkFHM6GEwjHR0Tfwh6HsNdkzAqerYMA6X8ltR5mnMjMmtpX2/knsKw
fqKyoF6mpc/9MirEHwZKubpc3rWjwCAkSVTr/YhArc0bgOFwmfC4k12L4y6EggMvGi9M0U6QPXAm
GGMyfU63UDKytStgog6gG9cUJUyZMDX//JaR4OFvtKGWWIqZYwNabExeawmMoS+6CqCi3ldyHR6Q
SW3SlF+MsG7TZNAJy1eI839Iy00b4iIK3cqSCwwAuB/dm58YC0/VRbWKnnqCu6XWr1E5yNcf0cv8
N2C8R343H0csW16sRZ75bMunEuWe1YK/aDKiRMqsIMe0CXIANtVNilDDAsUMcCX9RTlG5WB2HMHm
K7HxCdnyO34dHxYBC/hs2clrHnEcAqvZ0sq+OywErqwseJBqaqlwB6rwCiTSLUztRBhePmcCMxJv
9sIURnDzc16ctvVfdqa6pKtcqEln2VpLIvC7keY17/4gN0F4g6BMEPAwgZg4JVCUpb2GSmpDddeq
AGAHODlqDmLQVW3RM20m7d/IgshSubPmYl+c7e4txZIYkOg+gIh8LAkpvaCCO3+IZBc7DzijXFXs
tqzNUBlJWJ0CoIqXmnroO4aWY+dauQ2gSVJoEwGgLYRCSzrAowxD9IjasFF6Q/gmLMmwLMKNNTiy
Ns+rlcmf0E74d6V0y5ciTFSYiwXGYTroJUeVPM9vTy+c9BbFYJoNuWZ47W8u7xl/uplFzMYpfB08
tDx7rRoPhcpeVlTIsl7Z3AQ4hUvsGxa4OJLTckOHpXvHbxJo1SoH7Xs180oyWc460WoruaVbl/gG
ATDQkuQiaMoaLCcJWD7uoSAuahmbWKKmttA7qj8DnOXDeRFNK6H+PzmGrIM1fb0bQ2PoGabAIdCR
QhrfMd03CFolAciMnKZAgs8xhH7XNmyi8OuWaAMppSW/RsrXOsfBreVkaVE4MkOPw470z/tHKQqC
F7yXzQ2Fra5UMkALxuZsE+eHK1em2ovcLibSqHkUU6t8TlW/Nsx5Kj9vp3GwRPfWYBuK+eJ774VT
7YYxGJr0JZuTe6hYER8TZrXuKdWeQ4HVWZlPEEzz1qBEOVL9LPNstjcCR4+V4H360hOJ6wxwumgO
IA52oO1h5R53VYdQMDAJons7xfpAqLFVejkA/T5EVzmZvRqufN8qUWRVtAxZoIil/aWY4ak5xS4p
DKhSOlggJCs4ONt+GkCCaA4YHHOQyLEIy7w0DGBFz1PjzGA9QaZv1Mjg6Eb03rVuXvEFTpLDaa3O
G5S8nzatdmEadk6JUhXO1PBFW45eB6oN44D/UTw0yyr/97LHvTGpNjNwWKPDDApt2mgnvuEK8KP3
t7KV3p00QrCRwQy7lf/ZP8rVcw7PO+vM9TXMU3C/2FHBaU9RaHq3yALVnT+dctfJqnx/fPMFC956
E8KGOdXi/2wVvhVvF4GfH1jeOr1W7/iHPen/gs0n6MPToQk0JhU0JZpiiCV2PeT1RcI1m9+XT958
AdNAwU3H4N+CD9/zPv1tIN7Y9QozXEVQ7Opjp9d8D5M4LyxiBvKsfTccjIdLmfiuFhDYIJ9FVx/H
WtVxG6tBxDZmr3ON0Fv8+OrMgxj2sHmNmkDfFaCC+EJyb9KRxg4gBD6RDU3H+RlA0pmGetE9hrR/
fuoySzl3SuxhBRhDH5JI8kLd1yb8W3uepFbO+TIM8Is1WuTMIDGUpbNBLxkwM2+G5o0fWI3q6Yg4
Hdk7CRZKuOee9kQCswiyn7kAB4p7trLzMSRtlbwYIe8hlEoAmUF5LhgEa66xCrMxrTLTwuIK7FGs
AZUrQwVPnVxT0en7cLuTllCLvLN+Z/BAJjjmhykXy4+g8qMMWzIwLloBv87KtdwPON4aIz9ofy6k
XCQ9Wei22hDDAggaBz5ezvqbskGc+ySz1VUCsnOPaJR3s9kOYNdyLc2AxE8bDB4TSUdgbdTLKff5
42VInBfAZZqNd3JRECOBk76cHZyGFNfVOmkUII7iHN4DZmeiVIX42ej/M9+DEU+T7XCOg261UpXo
IrRigkt1+aYo6x/yJm3OCcl9HJQ9DkEtE3pMbjDqLZNPshhEmWDjvhDGuaST9/o4MEv6eRVuiTAo
z4gLCavimMF1h5PTmKpSyV/4AXWGi38R3b+wycHp8srEvdvik3zSxEOGpBwGzJ0XNLGKcDOaVdZr
NHZPy9jf0eno/VB0MkAQ0UjyFxH4c0hkmQybQf20JQVCCG0o29SE31+QkavPp+LNuFWSzOFxPc5S
A/MQYyINFarvqhwK3a2YaA4dOn+9cmFK+fcXSxOg9Ntg0lfaEnZda3t/dTDNs7rdAaLqzbWaUKET
JuHfUfkCL3o1m9quTnTQJ4Fe4RQBgznB60jBvNHBNRppx7Z7/tdBvCbSoTOJeGeQMK7pa7A3HgA+
rXeL0Vim4+Uj1UcVV2WNLsVBBPptbWGa2vZ5RbkQ9ld1e0gxM45fQ6/yJjjDhDsWb6IYbsk9T4M7
m4seO4JzEQxNFchZshYzf9V87Dxf5pIenp00Oiy8HG5o3Pt+iKvU0+W5kU/Axc8cCUUn2awxMm4q
aE72T0F4Lj8gO8MSZHdQlRZHUdL6iLdJc/v4uYYj6uofcnwljzUnB5/r+g00bUxki1ZCB55J5aby
rjSSJM873ew353TUoT8LMbEK0GyIoCCy2JIrqeMNJhdXR4QL+q/wojMVJ52kg3woMoFMJIdqph/J
92NDnevEN3XqvwMycianGCSBMUurZS2EAhGT+50tUMKBJ9GuxBYIVZ6/ly5aeUH0/1VyMV2u+7Au
a/xIxNaeC/94EoN9Er+zK2PA7jNnkUS4vJnnt5rUxxEVTO2XaFHRo4n9ONkcnf6ej6uRxJtXRP3K
9mAGH9ZDhk1RSkFUVciKYUzAz8XjjiGenMu3miTp7cYixUQIMD/ag57vMWrqyrJ7CKHl2LtUkzcQ
UGSCKDsjO/DCx8QhZnPeITjLxZ2d6jSL9Xxib9rpfsEapnnn0o6X10qN8OeH2YGLsYqlkj4g0eNJ
n+T/aBaIfycN1XeM9OKXx3FiMMMgoRKhM6klifWELWJsDJHdWo1xBDFxr4EAnrbmcdKZ2oJOteYk
bw6gBIZpOT4KOAlYEGMXrnAWUoz1Jkce/xq8dNixUcIpuKxrG37oh4kOXGM6NhhSRFso3+yxXIow
U52Qb3ud0ukV/mX3Jc8ccOw0EwQCWd3dpl52UrfIYXfgqJ5U9y1FvgFpAdusLqh84Cf5GNj2X9A1
X1YGfvQpa1QNvb8rk4vWhLtm8WmdDF/R1nX4/wUvWST6hdZT7IWVnxrhI21noqKuntrawpf/Wk/0
HzlkGVIypw2TLRDWbSQjBP2TUAKmZkRORufnNsc6SIdXAJdZDxEEk8J/dYmOaElavqMjlN2lwj+u
3AEiur6a+o3zZPhjaxKcyPl3ClR1YoiJf+KEtP0iysSWhq6wrzMJN8uGaR+hJSSxDeX0urbQuulO
XwWWYcuX5G8cQV9kdB+I5VG3ulnptW2dqHyXAmruLWlOmvTm/3opCq/pKrL3XzWgFy0Jfqruaclq
msii7ae8GDeYHEOnYpy8cSxmph8sDN7fNV6HS7FL021P01HgjhOGaXlTv+TtCf6Lrh2rjMXsIsfv
y9TvSVmyqqrbILa4UuDeq7QPa+6Sj3qx3za7RI4a1Cfx056ThCZLCbg87zKXwo0fahtkCgzZb/T8
8qzLFKSHidyfbADa/+Mr6ycwGtGZi/BKLXPJ49wH4c7vR/dfwsRfse1C1/RV2QyWp6ZZNVGon/8B
72vzp/zZKJBp/wWnyR5dJenabewFPEbXPOQfSubejsEDKNXKZtMVjkDiEXB8ykmlD583zln2l8WC
HGSTH61NSBnpRw53Q99gorwb6jzF/EhEAc+L935Ppzn12iw5I46ahg5wLd8rACJ8Vk/LRic/ZoPq
9T4VFGbGA7/fsdesrqMTP52pmXyudZIN9nbHDxqs6cZrkLheDE5djJ4AV0Y0bL589nyjhjBOvMti
aXnhrJycBw1JoExIXvMJJV5RUb9V/hc8RtOpQp/ks25iYgxfR1ArtuIQx44wulpMfEexrSpvk9L/
8xTWw5T5vy4LjMbPv50x8NAJ9SLSsOjTyw7bJ6iLaaRQtJ23ys4voL8wt22PDKRzrb50l5WUHYmw
2Qw7W6hx15/0O5fKDdPH3cGWRX705shaWkqUhHQtieAwYuJP9mj+4PxZectN6zXvBi6ZpbzGxbAF
sFpOF4N8JnSX+/93CGdNLUKYgKZOntOJFDVGYHT6uMSCJnaLR0WZnd79Qb26BRcqcZKuXe/PRpOd
ZgvSjW0jjXkAKPVlBXaXj6rkSLbV7PV+OZukepZANSfqsWAm5S+ou0/VRFpxz+hP3JsOhA6gfMkV
IUQOH6EPzGkiLuzrKm0N8EgNrxeoqIGiVsoM9Kf64pX1aaipMaXlmHIVh380PwFNtkCQJoy+UreU
0x9MHp3DEmKXk9ZPWse1U0S5DlsSP6ktZ6ZH8/CLSIyceAUeRbKSscsbimTIGYfA3CyMKxV0UxOw
Rj7mX+5c97Y48sOrsYyTtwT3B1j54dsnOlRWNv1elgwpsI9M1k95geJW4MOh59EkzPjKB2JxNg+3
983aMwkMcwwzHClEyq+Em7v45B5a0IZ5jFU65BNAuQHx6DSxPCzgKN2TePv3vkkUgUr84mp87+Pf
0m2T9gooyXon2NfCNFmdH7aX3BEc5FI0m9h6v780XW0FOaXNHArgLVYHEcgQu5d9ym+bZRE8STz3
XGxHQidDdDo+3r2VzbVvV++dRI9dg4GNqJJqOgqcnj4RmmjhGi0gcX6XUj9CqyjoNhiFCxCO0IwP
IOqu99gJFLca2i6sXZk4C6yAW1kG2s3jP3ZbzMVeCxGwpmXsr2lsKCOJW/gWeNYXbKqGTNHHiIRO
e2gRdflEFV4FPHfUONyPA6OYVtguiTshYZx+plzK1X6WhYgBPwNyVLQEZTY8PaCk98Q9LiVhPqTh
6/aVZ61i5eovZRSv4sxmyeuQ++Bs4ecQcrRVv9hUwGI988xY9baYqbIfP/Dx7o7qq2ngtoSb4iaD
Z1d1aJs42qlX/jqB0DrfMBuePMvCLG+VC5U8kE+yb4OJjkJgDusweCtIz7AsPfFXshS/v+NeLT7N
YLhqrEBrUfdQ9YxfxmzELs45ZtCHgoSQMT6K2Xlh+7LLsJhc0vrfcQD5VAiey0zrtghXAKnBZwN6
oagm0iFHPD3f50MOAtK9T3hMWQ/pZ8XBMioE5RYrOyVDZr2iLytTuiTm0KGdHsUnHBZWN9PlJh3/
2uxZlbxWyQ05Lv3JRy8w9/o/ptDqoMw8XHn8goi1l1n2UI3b15zkD5kQgtD8EvwBzTJ1roSjr+O/
FMEFx2eEo2RNnnQ056W3HYUn6Oo8SezabY4vI5vrhn8WEqhgggjO/O9eZ7tU1ISCUUuDq3en7bQm
Fps//frNr+jvZJz9XicS26hYH6kNhO2+Y/Md34g6Zf9at+3PFjDMWgVe1fChZXV7lG+YUtwqYSTw
uiBtZVrUMk74+5f3CqdFqHGEUMwPAjnTpXYtwQMowpBRqkQ8xAPsWG3h4iHtQVYnPd21qea0Et4d
eSlRXJYsjXfdvdkXVz7rIPwJmy+oJ1DVQAQzO66YPdPxyjHae3+mTnVrehj7eldz5DLJACs3OABw
Niuvg+xtVKZkmYaeA029D20ApefPsaUGelskklRb9oZwK2nEa+zEaCrncKctDnguso3mCU4+9dBm
2qpY0sDCL7YBCq1IHvyU/sDnCZzk3EdiqgfS7VeUbA8mX6MFkoV79fApNOOghHNBjY5MoWQapTEf
fHoxnW0cCF6jY57K4nzUeOTbkhOuCqhXkbqT5xzmwcleYJaHWibxHEc8dD/ERLSG/7aVMkQyvb+E
QRsNS6x5P4icjBqpCSeSQ6kTV7cTV9koLwe0LRiryc1zwRxjzVNKwEf4P9GDLTD5/Vpy+Mv0bRbZ
Aks8I6PFFNQv8ymErx3ryLlzAoZtBUfs+rV8Uem5BOgjupMFK3so4dhmXxiasw3FsFL3CSTDVi7M
rA/qgf72/ZjNP1Gx3ScQrSATtp/p06nKIBKfF7TyshBVpBxiUv9BRRg5ayj88vXG6KfD0F5Ksm3+
PnVaY2k2FhP6R2X04quv+hssPJpe+NFzSU2aUOqLym2foodJY+9WS0XD4DbDEaJckqRUlYKqWw4k
GOcraqai5nfR9dHdR240Tgs0otZqaB904AUNV33PdAQSiPVIBzXmZoWRYX74pUNIqwnPqxBOlk+2
Tntm1oY5l68ELX0+xizbEO9vL2IIyjGbA6RZpsEz+zBglaK5T89zbP+06CWgoCTG+O8EoUaluB+u
My+KCaQL0DTlpRMSeTM3cFHUf/leemR51/13PRKaezaXUYVI423038Kr9Re0mt9UWW63TbkMZ3ii
ce3BCQJZKWdMwNIzeAzj5Kd7aKstBqYK35kBPeR5afPMmio2WMJU2RyyKNKXFU81Cf20Ns17zVNF
y5zOEgY9hSlH2qkCGTfXmywEFGOGOaR6kGJgbqVStSGkF2nNG6n9fKithfgGlTTZv/K7j+IYNhrq
SWq8R47MNjGhxx/xa70TTE7EzrdIF6ziIf5YljTByz6/x8BMq432SfTWal18dBgKZ7fz6witENzn
NdB/1/IlHTTEZ6Ubs//3hPUXzmmKbdEXKtRMNal83Uph1vYcazkh5z2XfP6fwaZj1Sd+aJNXaVe5
ZRFx3YMqtyvzDbIwfQtFRHa2HhAR+ulfR58HMY+E2dGX6uqmoJLYtmi8fG01iU0ez3ysgLW44AaE
utfJGN5N5ygYnpcyXBpwTM0XHXuJtTWbv9p7YridBKUnQ1foULI8uwCIHT79MIIkPhpKic5dMkGH
NxDgUUQTYF9YlJ2jz2oiTcKDTgv2Zs6+4PQ/V9Cpwz2h3t0dAXiNGBcV5NOv7yp/wcvl2hHqbDfx
O13eZzb+U29nyEfsUkPyS2qVhwLYjgEl4CmiqQ1MSoyOh6kjC5ZMibo8XzddAvPWRwaiBt4lkN5w
2wScb7McCDLFug4o2hORMa51x789dO0IMEHXFroewG2dkTuiCZ1o7CUho30CcYt/an2AvPpGIBmn
M+/upNf8zyGh9l5iXoW3XRZPfWGf2TvXa4rBLimReo5WCBwEJf9eqTQ4MEVXVJGylK5NCGcfr51b
iltErWpkmTppJgh17AeLHzHoU6UPJWFxGBhdtHsK69vsnW9oL+wvtHHXwE0eZkV21gqMHklmd1sF
lAyjViwFpzNoSyAszcYAKismrpm0f5LLrOwo1MonktA+4q+LkIV3MLZqFbophgKLvll/cY53JOIP
k5NPq2Ztp/a1hPL2Tvqs7vh5jlIUjItFWFMUSlgKWSc5Sril1cAe7L9qh0QqiCXA4Cjx41+IoZck
jRVUjAI2lqZEwfCpCj5QibhmhXYt9YOFTBgzzroGnFDS7kYlnwEUZgREnNlOx/ktiy8FslkULqz/
Mqs6rX3TRrY93n2f7hfn6p4BOVEYQyPM0CgxDPB4Lmyq4iAt0BcN7B7afVD5BhgSWBX1zLZ9wDFn
C19uB17hCj7oILYJ5tI/YyPPD6KMAdaMMAMA/wZJU5uCk9XWue8p9VAj9X6ToawiL/+Tjsf+975L
eht9Q8kebIOJpG66bTz/+Vs5r9fayU4z7RzNL5bkwYUOM1veIRPnxdszr9+nk3mJLtJS13qDVR7w
HO6clcA3+tc6WTabJ29yOKGeayGnxCnTD5VnFKcU8/xzjtlDSv3L3Q06bgXHB3pFYQbvFaJYIh7H
POeUE7NL5KUVmxBqgDqyJbs9Par1rTUk5WAma+7yMMvYgxcKKaoP95tXIOe7QII4MksBg6S7qQh9
bXswQEcIcXdX8wPx0eske+MF3IVfP8UUSJAy3k3jNxHgYDXx6iTrRjxYY1XS4c+LsB9P3JGHKzxB
GzutwjJ5XeW5qc/pLNG+XCcymGf2MFpsOKaNTnFzz4SPrw1DLgHFmNbKp00E0mHawyvf00dSv1Sw
ZndGp3oykeXSGCm5aAQVHB9ooW/6qn09z9O18AYmtnHH1ALNvQvUMWKeaBnp4+Bi6OQVUZVhHfcM
INKF8szkIC6NkXah7SfBMnfpMVeoKr/R962/b441X2oJZIf9hIlXaxf3PHAA0YAz9iwXKiya0Rqb
idWDNVvO7g94kjcD2GOc3ayX6XKQiECgAjERpvIHXkZx871JlTSUKWsVb8jYHJiYHTu2wE313Gh2
/NX/XjWcxK1/qszgBQL2xG+Hv2jxpMt5iK/4qY4W8P2Nyx6n5IjsjJ/Y+7FGAMCmFutYGeGXIqze
0V+x+iFHtlASxyHKNOp6uZi8zlApLoAGbZdpwODhUMl7k/uZ2OCQaND+Ks6zw7pZVgQGd6nuyaRg
bYScNbYq9HQvtFO6c42DI3cZq1IYndvMXfx2MCxTaA31d08mca2qY4vmkxwmQzdSIBXMUnIzx+9V
o5tYfUowQcB2oJZG54QDsc0dPPkwJtikNBiBYo9FtoZBbbKof2JNSKrBOG1ORblU1y8dEHNJCndZ
42Zr60EAv31kGV0nowygEqCS9HQFTuZZUI3Pl4kYUQNJh8V94cWxgwh8lHdfK63TM9STBBfOoYhd
NWkNbxNRNKp1GDiQ83KbRwKrGCjMrLV5vh3FGmVTtjSdqmcpi1b+ZrrkTk4QZoxyt56cEzU5KveO
2J5QoyGPyuxugfxiiFpTjMnStQDn7fTMeAIFiafpDdJLs+pcmYcYb+CnhhbASUllPUU9y5c1LIVC
8d/OOLhRdYfnm4TqWJdDxMkklBsO9Z6yAlUIMzz5BfI6J/kFjGlXNOARMREX1RTT7cNUu/mWvGQi
sy2+HCJ5MM4j5ecH6S3DrDQ1NRxvK2emdp/5mAzjaHsUo5wrOR9FgPC1OrXvTTMJsmGivrGROsg8
qLBQ5aLGFzCfnqzhDcpkCgBsx0Dw0bjd/sofap4dofFdiLYOwRG1ggWyIQFyClTe+vq2oNLtsby+
2+pKkAOXiDUVpzTUwqfomf5qETHbAfcGMAtQokUbKFZRr30y4Eai4hiW2dE6hQJYRKlxzq3atf5R
11YSb3TP9HYfvBgfFCTAgdvxb6Ytii1IALSPzQBZJ5u6fkKAt9uhGFvsy/Vyzy0z3Uu7SO/88gBv
AEUMW/aDsoBVRmRb2a4tpknkLjAgHkMe5HvP0NqwPrniSoPjAslXGt0j0y7jV046Pn73mOLidP2f
igalSrzqUuY8TjCnk4KmIFdi9BBfk5ZzPfHZthCE6GBlRRrBZD/o+A6XOjpuWV/+E5pLIMFsH/wM
0Gbzx+X6k5DJJHtVV1TtpccIK+VRvMsK5fBWuISH+sbYNjTcylIxqefp4EPb/rF5jfXUDPkT91Md
jwWc3VUb6+5pwMlMtC05D0u9DNnSdKOM1diWojcpOPCIT0hwslUslnY/I0JRKSe3XCN9I4Sk1Y1L
VNJ8UFO61mFCXd4upqCEuSkp7qwe9peyU8eqPFjz/SRscUuyWvJBd3EIWvHMbz6zuyexZIIMKR1+
T8Cd4+d5ZszBGuTecMpWpWDjeadK0eH8rJn4f82jXWzzxwckOp0Uq8/8aByoPmBAfMQ6Qnlwwltp
oSqy/iIcJBOOLzVX7eiE5HvaYqILV3Tgx4KpIzkaI0Snlzi7Mw8KASvoQ/e1quV1axkwYbFHh6e8
+pzJH93D4pbMJRJml0JKewY/faJlfTrc3e82DHpXJIW83/bmLaqkV+rhnMIkNn2m+he7pckJnG+C
zqJJO+QiWKPqvibIqvJXvQTVgU0VoosTQtrkw3PVjm1kLV2FMBbJrYdi7s9V1wboe1JiHOe9o5ag
D7V3Zz1Wd+s+2vCyygW6jyTAriA9cawOvWaHpTToi2dj9LA4oSPhhP8+DFG5GzZlSKEatls7ibev
vdhnNQop1MsytfjjOtEW6td7YNWu3r30mzttzOeHX7AccAHuZsHDCPzTm9zlR3LzGHGJaxa0P6Wa
ETHhpohHXzGwBMNY0I0BU51kOrNlmzpD36BG6oz80VP1gUu9N1JAjUvuEzwqkQzCVKHmAMuLujqP
X9ntgUXI64L78d0p1y0t031XuR6XKXFJwVPUIXMFPt5E8KPaKfZ65a9PRbnYqZQGGlW2vRCXDnWc
EQIAPOHLB1zkbW6flkoQZ/mwb7rHIzgkPnYLvNlgbEgMB8aPprFLPbzyrlUqfp5lNWOJopB+vUvi
4TCrD4DcCkQ9+mGz5VgJYxtusCBtWe5msHqzpwTMPJ+yNahRaYVAPJT5xI1zSzCugzegGeNlhl/t
omSRYIQak3sifwCbAk9KY16Sz/LwMmfqkoQN1EW2ckA+2l0IoMDNiaMGgxIHrmD7SttQ9NspGX2C
OWgvJbjJLQN99yoNps3FwvSP0YpAG3QmmTV/n+TeUGixTyuShO7dd5dcJkGeSDCb52tylhcCHGiy
BDoXPvcHhWZDX6njCXsH5U1L5/2ug1AqHSZCXlRpf/3ewrtTQ6Mc6UJ5ex8o2eSXCLDxMxv/Huby
l/P5URW47NzMW5cbxBZ9Tkb+L4EUkv6+zZLuxIrnA6EZaS9KmWKOZypZvFxXUr91qwr+HCxxp90C
P2WJFeAAb6hN6coRlICVwkOQpok5WvyzI8NdFp1obNr3je5g673yLwy3NkGoA9mPslT6R6povnce
sJXHNJKIkeneK+iW5j9++71HTmFtWp3LdeueAzW+WEQ3Sb8LoRxxj0PK2M5oHTytYP3oCu1aCi+T
f9EwLIGjysDr65uN5WO6q4m17bfIy0Ca8Ugbs1MvunjTVXw+hq3YojXyySmHMlejaJbYT1pxh99n
VOifLfdbHz0VZ7kJ2uyZ2Cj5MQqfdw/tIbZ7eyaz9FiAfpMINR7UwG/ZSh1op+K+6dW8PK+/+L18
rJwEuIFCM0q/rn9iGov8zL3KEij33V2oxJGtgWkGwfjc2NmyDFrK4fz5z3vX8tbRa/KoGIqi79Dd
kmyBgkHN4BZttA7EOg+H6/xCiTuShn1AYVgsJSxo29Qc4GANzbCJkps/Zt4Ebwdh82HAxR9NqGrU
ktClZp2v1Db6hpJXQFh5YSP9q3tVynhG/sWRiQZJE+S6//HjDy9Tk0TnyubKBStsm8+AwJM63ErX
1kkjb0X2PxBWbm/YaJnKb3i0POb+sh1YqN2pZyAdsg1sh3anQ6hBOxCRsb1bBT48rUpOGRHvcV5w
chE5Z8V6FU+02WzWqeseIkzFWiQDYHgAWQmmIcO2IFudO9pYRxLsvabplu1rR3yIA0TpyLW6dfO1
i1GLml1ViO/dQWpaFPwQrLkXsr3O3YIrtMzTCD0pRiBIfJKJU30RxvGSuSNscxzq1yZP3rIh5h/B
NiRiPhVwvYgU2nFDgc7fY62KvzD5gPVO+V7g49lZYUZgGwZvm9d9TX+sU4nudI+DzWoggfzUe8Kp
IU1RjblGZee12s5B0dtKal9m82FD6gppYncKP8qsDhf8Jn5HI8xYAoHHJncL2mcCl2CUQzWnxE6X
rl7km+C4yXi+yQ1wtlm86igGPrwnsHFMCxpaYgJPr4MaVNtomKEiJRnY3vyg2My09YPh/GWmK9uf
CI0x3jJDG6KK7KyJw44QozLfKC4RncwnVrbuQUufJl6q9XuyEsFCpeI/SO0Ayo/Dj58ErTj6QVG9
PLtFkByfNSL8BhTHBNlEuLUtJmby9pbapCt1fbviENrdNKARyaY4qdRFUoiL5BCRaOokIkkKyYHn
SqyAzdNE03JTODtgugEC684A/bgUXcoSTW4LXLiET7zTaCyLwJGBnzV13roKXtJ6xCNxHEISWkVg
0pc6vIr0pN1s+Nij8C3kR44iPoeKDD9LnbxMqzdMrYy9UyVmOLPXASRrKHzfPtafSZ6Jskbfg4Yr
DB0T3KuKpB8LCTRkoa7uinc8L6ktmWyyF2/vzAk9Yqzq9+xwUhbyvwoqzQ4ixUeIeA1oZdWdPfsb
TMCfppkj0DGqKUHlKzSvnU3ktS5jW7CWhrSDZ0s2HEhk7H+VeOEa+RurEDZDzffNCvGXd8nmszHc
HjGgR/7t1CexnjqS0YtjHSFP6qzYC6b4aVG1Xm8wjhEW/imDdPLOZ3IEANfxrZiiAnH6fJhnNIzl
FknwyqiqHCVzh7ULDfuBIpAJZduepbtQUQU4kINI6BFP0UhxweuhizQWvg94H6dg8VgEisIGC79D
XtUBtOkJjQFwVvABjVhGLBYvE0K0FTNYkRlFRnEXwfw+QgrNyGbu8pw4t4skq8G1KuIfBIhEVLmM
UGZrWt8F7XPJGOvO1fd//ZZYtM4Q9HZRfk/R2FcA+98tjl0tfE8BudBCyRXq+X/E5Mhvmge9Yfyb
H3be5wzRsa/UTBcTS7FVhkjnfygPPVbRuSDpvVZccGmvcj6bUg8zmiMXgflJUM5rvk330sD0y681
Y1Zd+FhZ63S86N1DEnOwlX2eT0CMzKKyMGBJ/dsIUZNckOHt+rGmjDh+hpwquFam7pTNi16yHhdw
cczrwDQbjkJZZFBEejeBtqPee1GIpZsHYD/OVC0dXVo6Er/PpsQ4vJcLAJ01H0C6ecc6ix80pa4L
rrNpHAmvW3FIPE9Mxbo35YMd/vSgbMeEKGRSb+7/o7P8YXZrzN1Csn6Q+r59ijjceoeiduzF8Gx3
9I1viaqhZSgGSw3fkufl2y6t9MQ+H+wwcYNwPvkXQ/iL06bcjzPaVMuEDWMJxbsSS0obhyCyTGTC
aqLUTbsih2H3dXoXuOJPHmUeAMzLWU2veiKzCm4XJrmtbcHiB/NaY9YBS6n+v2q+zHsma+S//Jgc
/ZUlB3qi43SExffV4TXh5HDaj3o9agEosrC+YUJZdFVwKWty4rrXPg22WnU+/K/NwKcNStOp8JTp
IMkJQaRD8GrlGJIGNLjmql3PcIyp/OsZ1wJOmVi+iOCuitGH5tLnRdLbvClS6gE08QRIwSw8SVx0
Zj05bVJUIeO+bRj9QSvrXw9G968qv9nQaVcVqM1czeWviaQvnCZbXszc6NNPu1DsZeuEXnrAp4OX
x5yG1AuI6LcOUlKtkBz4chiPcnVts/m2B9prGj+2mNGC3MkQOCLQMdaFvfgzU8r+nF5cytLDh574
oGHZrJEnOIteQHqMpBCI6DnbrlUt61shxXu4iizum0/Prt3/NBFRpbidv/ggMUZRKi8qGMcuQj64
3DQVuFyK+Jr8RhDHwU19WRnYV471BE8QyOPT55SpPgeZSlwRpsOZOkLopn4X5NZsI7BsC1K5K1j2
q9um8wE0iNs7btprEeCpQ8iuXhmFYiuEtyXeYUiNU/3l1Ht0njeWfvoi4budibT7oeaWC70RdAN2
bpRrXY2abT1bhr6V9th+UF/S3qj4ahO6NhtI6LE90/5UZSlT++lW65a1AwhLR+TssGUaJOZK22rs
sFIc40PJl7T5CSjoylY0eQKyRoyd4sD0EHNBsQL5mhVe8akJSEF8iWSXPVxqGG7Ncvf9CTHyeiJA
f6H+hzUgI4rptlS3fRk/ADEb7AIaN/ebkKHbQ2B69oF32eKdz9LMATODaZJg9TO15KDUDFNR7oXM
tPzrY1+3dvFHRbNw47nWDVBh+soaKVKy4x1s8PCZAmsnvbysHqPAIxpDb2mPUd9AJvtfhfH4iGVK
Yfi85miqVaywEg9UCQMaGCioE0/FEOArWVBPv9kLrhlipJY5CdaYTIjRsmtekhYyiRlHu95anWIP
nBxcDsLYQDsCwTWDckGYlYy4hFBaH4BbXa3nTj0jz68JHGq/eMDSgu3dIu9ncGZVnOHbVLvwajpw
HsZ2Ixm5LABp9KewJ6cgRFwSzAShGuYLYACOcSV54DytEErW93hUGIxpeWRIYjK2AOBqWVcgdMtC
LzHCQviPLddFr7bxEn1eY7hl63gOialVp5WTyVoBVi5xRoA+jfYL4m3hD8BDSQ1v8Rqa5Y3PA7Cf
kiIp3pb7/b93A4DoR7vLUlz1a5JDzWtvon1OTiHvBUM3Yr/q37TuQep31sI6mvrmjhBWaMXGfeW9
OEl8ZsZtnhsxERg+T1lCoyx2WlGxPnxFTH1ai3ADGFknP593UKAsu62Eii0HKeiWOkZVkMsQkQTM
Q63iqGl2vVwhqOR7FdYe6h03BEzk+jMVSMPMvRQd1j9wka9lpZczU6vyDa+fChs2S0WwM+vSiuhU
5s1IeMqLJawwVsLMVEbJ7Y139F9LwvoCaGrSallBRYsjr8MadSf+5o8nf4sWue49S0igrIEhyRaY
lpmyFw4UeYforcVmDkjzXnAgzZ9vs9fWLLQ1eUq+1WHrDUzG/WnNvH3dqanMy4Ix733FATS3KYLV
ih+/W0/BM8dESbG9F3uTugRpa6PCm+fuhjJrt0Lf0NehkIS17N2G3ehuJbRsiqE+9kAZ3iT9bisW
TjzD3ORrO3mFdX9qInJGoixKNyb8hd4OeKSh0NgknyJYyf8PglYW+GxtM7tq7mzrbNTTeq8ltG3H
LW4YdkBPY0lbsDY5O6tLhBRUG3RJ3zdal4KXxkZeFanKCIrAeeD3LmSWGQ7c1LMlnZCPcZo604Kr
soBFZFfGXUx03Nrfir9baaiI3bQ4xUuAFrZceRdTU+FlZkngCDAVwCbSExl/1lqCJ07ZjHU/ScEK
ne/nqxtvb2aiU01trxJX0Q84AiFkXjHoSO6KieKAx2/jXiVD7IPom6X2uBx01B69uVCR0BeT9efB
RgtGz6cUG8E4OPDN8FHfWPokqMIelWcM7IA9O+3fFj9ShEE/GqLBVLet4QBS17ctMqE8ZPNT0ur4
2A/mzJNa6SJ4MBfu/+zytZFaI2EWnSFN8EnT1DyRDyhmZR6g9F1EZdNewqFkIqFHul1bcjlsx6k8
fUlLCqLVd2B0WC0uYZsx2gSdX2sL6nsTf4YuYeRNIJavxcaVaxJcc23hjBg0xqia/W6yqwB/viso
ZIg1SqMhMETK0EVgm2RrI8LPLw4vjc0+OAXfUHP410rD0DcsruAPCfJbqVVhB8U2bKKLJcw2MWmi
qlJf+nMrsCHzCFNEtZdTkzQeGWIe/8muMt2ZUNT0vzgfPP3AcL+FrFnTfTmW/0JImEK+L2qBDc0M
KQ4TL0lNUYkp989jWflpXxCYMjqDnD33mq/dtCspShgFkEbDn+wmOoVDIKk41gN/o/OhzL/2kFPX
j+Hft7+dZYzmQIqrU4SI3R/nnO4mcjTjQhrSb9sppCFDYB2Xu+PSE+oIBeIRsyXW4rwJwZeQWgI4
mBNDPTqqos4eDXC5MiCmpxEyTBoZm1XTAqX2VnpFx3DJlc4WOPeTm+XeOJueYFzsk6FdenwLSjbf
6i9kxdVjCvf0c9wG0LMQEUgwr7XiOUaggsFNv3YUkF26bn9+iMP099uTPUsTF7fzC8no+UCqRq6y
DibgEvjzrzHwrpENtkVKHrROBBOI8a0Ywde0T91h3mVIoXqXDvH7PCLf4xopy+0zOFmVuqRa3E3M
j4LnWRFgOiej4yOcRPwl1s02v+9vvbxBo616uhDcZWkl65d/o2m28bZL4far8mkEYC0vbO56+jnX
fnLTZE4uOFWJDyo5fUMARY6X34rTiQ5q4f0JW3OhveWwF0MFKgAo8QbZtZ/2jCaf/Fbv7+Qhs0Yn
Ml61qrZBQ7hpS54FEpW4Fy6Apwj3KHLSP36SDozuSTVvR43BjvkEGNDYtDNEAqIFpy5eAyknCuJR
vtl2iH/w15DDDdr9OB/uVSMj7J0h1CLuHQF5yHn9tqhhibKJO9hkOs9qD0l0F4aFIBWJLBtQtx3p
5PrvPDz62rtuReANRoSFQ7Ks4Uz9mJVsIDeCcqcRH/CY8Dphp8AmwbfOAPa0sDtxIBl7LM+xJlOQ
PvRyf7S2lJVuiuuc2YRHmgt/kwvXGZzwYDO4siMjopVmgNitG7H11CQBnEcJzYdU44R73EpvBSdM
+oCTS8CoPQaXRUagVV2rTcZCSgZBTB6b5uCrWfim+OVJmQZ0ZcSANKn8H+5eyT3BKQaYmrnQa8Du
S1xxlDrcpsf/EBQxAikMFnr3ZwVv0R8IWEeKJzdamLMTxUDYrSFok5biECxkQsr6XPT3zKiZHDOv
HuEimpGdfPlwEWfAuMrT8Y5/L7EeVIDSCHrUcg791Jwr39NgzERLijDF2cGN2FBA6pcBoYRiiMF3
J93s2TLYomwmttN6FQULT6V9G4IWgnS6jEsrxp/Jdo6gfhuD6sRVJV3GWxNRYXdHLtj+mL3jOwLI
Y0J9YTzzXp7++PHZAVQ5wUNlk9vpB9YzEb8mHkFXYYE73x6j4aIGgyK2PjzjPy3wemxZyZ7z3rK6
Z9aF/9++sBslVOY5FWlWRl/Qpb4/HVLsd71O4bH2MFPr/+NHVWZnvR8iprimdbKqHADDTm7OFh7r
FKHgiOZCK3mp4wphQnzEDE2FlvPXR85a24OG7DxuwJg9KHbxmk7+O4RT3rhCT2/BKKhfxDBX9oka
lop9366SC0vApE9kCDXMalqUBZfAPoK/v00nmyt7t7f96qMpDHIDQpT3/a9eo19LsfNEft3GHPP7
IOI4XEN1XwQhOxrgskEDT075h3qdAoZs5cJlDWdnVKXG4YrGodNv4BeT1oPZV8ZiNo4P8ZBBaHkx
WQSxe0pXG/HAVkA4Ala01D65saczdyBDvsiY+FlDlPifeE4y3X5vGhR07DMkGdW6j6Jy64u60PmJ
fF3pJvMAROsKLIGIsVv8xR2BGL4VvrCw3Qm3t1TIKdP/yB6bbdbfDIgCxTueEcIttxTjIpoHI8eZ
X/sM7pFusd0VABH8ucvvq0cJM4EL1LUsT9J5fBZsq3olhfmYTuo1iXisAVdjXeeL+hJnUEWlgRFG
/aOGDl+MbkzGE1mtFL6OGNQc8CJJsqZF66AGQKH4wn1XW1WV8vy6vqsgJ7wzoZ0OvQmtjU0HIn0Y
/XCpGynHihVtiM15C77ZQ9palptMRyFg2g6R1ADq03YhsJi+MbxEVx34UnwjJCmwFZxArLFDE2e3
owTpyuSptzgE790mR0c/GnuVFiGRiVyFiaWZMCLtxmmZnZlHHtY6rslUAKwRysKpNNzi956aLv8c
BKx+dOkC0z/yRuleWrp8J3Sr32orDyFqRw2fEa28lCaIsdT/JRINEql3p0b1UoiWqspa3TNnaoyg
xVQLUElqUp7htjkAUmMmANNOJWtmX26brJJto/F1y4XxLWz2xN3+OKcviZ2ce0sr2SZDfoyLwBiM
0MMj9gYOJ69DhiXA1bYuqLTtyAMIgdWbp5PnzFRc8nHnaNfTNnxeohBp/D5O/L0cRGWwHLHj2Xnw
CAqFS16jvHJUuBHI4IKhjHy3VcLWDZpZZ59V+g8VA/E66cL942bp1VcLOybtunhC0+Gr3loiDGU4
rluX2QC8TU3DqO8lbDK7/yMtNQv4myvEQrjfRs2wgpWy41v/lgdR4ZjVtXdNDs5ZHoO2JHdqfn07
t4qWHoGBTF0BD7mPbie42kWUYnImikUp7HBIDaScZjVic/tD9KfRD/8vej51kddPgr2z4y/zS0cO
mn0VkxxEXvCue1gRj/eHPQ1zDzjDyAvBJzs7WjjWX+PaHUpoFcZht1UxV3umvncg1R3rKmijtBNn
LVm62W8UoUvkHaCh5FCb8OfCbOWWXI7HPmkLP+PgQ8u7s4oqr5UCxLMdz/vUbiqDy38tUe3otVsY
YIeuvAVtIjXgONO6mbzAmAXqr5YARBw2G2MnyQFJSgKTAkVDocWL/jmbIWEK7lJIptjQNFIT/4/T
Cnj0OC0AFk+mFnpNQMt50qaSD2VSy/LZIkUQJc2XmQbqIdmC3iGqN2nKIgqgpyUMUMijYdt0AVnl
kxXhu8By/6OHJ9nl8gfu6rlwAu0LomZ/XUapr+BZuB9g9NOiplsSuGLUiuft52ETUDlnJ0TgQ8jv
0IQYboG44vlZcdyVFdfNUMgL2i05j9myQ3PHv0a+MUFtbW/PfLGdCTloyoEOyEayEquz7ghjXrG6
fs5xWHg3vB+zth7EaUdZnWTDdNmVzjtzF20/BJ5+FW150RQrdMljcXv+K6a19aAnfvISkqI/jDJf
eRkbjsC4P+H+9fJzqOTnwEfLhkIfXj8VH5Z6jPrwdA2k2yyByhfSzlYqaDjBcTzkpcAhO1Ipyohx
6+oF/u/Y6+1/H8FuOfYkiGcrEQbCjhPqENU7wynqphl/XOey8Kd5Is3a6IfgFcITVWOg7PsRW7fW
6SqmUNk9dj/Cz9sw1B+u2X+QlgkPuUtCrCT9l7rkkktn9cr4rm77/J5PfpOVfjQ9mjhXqy0F0zNe
ex3wrspntuy98FtP58K7y1b0QSDhEgJUhj3S5X+pACd9uE9WOQam59f9E3MPt8OcHvxgvVNHuVhu
5xN2mSjuXIUk2Xr33PPtqc2lDBVbjAFSny2r2Ie8ceQ9wrCa1Y+xAHlHrfB8pxGfqU5dGGhRhBOi
+qpcF5lboktGvuj39BBztqZQE4oXIQlwa/jnmGR1egY/N92qzBAxbBRglMrAOcMmDdcLalLAhc9A
n5nalGh8x8e3PCNveqlCav9phPBPTAqExZkALgbaBAsTKQk0H5B4Vt67RqTnk17CYpYfGwYEA13C
a/0k2ofMUFggieL1hWTyZasM6NSr3rq5F8ln41X0djoQfVmhf7HFR9mzUYXAbSoFBN5eDtH8tJf0
nbrGX4R8G8XDI+9wTC+hsvdD7xQJyw7xtcJhl/f7eS6cioAO15Bgiq02Hm4zvL1zuW6M4C8JmX4m
YH+WTbVQ9AxhA1fm6bC3sPuQFzpCPAsPKR2HGb0UHnaxtMQEhMfOFVJA2mB/SbpnGwuiBDxri25G
PIzeCVYsDzwHTYWekGiFYdxaXGXJfz7UCneUfLcrSDk22KaqLa1CIdDME4/C/785uixEf1Q/fLTq
JQSPBXn6AHmqbi6sYQ6E0031P5wTWBze6WjmjvTd4d/UHqismd6ah1p/S8fmFXBeF2MdZTPRvvgA
P8s7+RUeWLZUIcbgpZh3nLHXqiK1hWWuPPZACiXWZUy2X8XJ9hUf3Gdhrt0H4S+42HAD6Cs4+Wgm
fiMQDI9GUO2J73MVDAbgzxhQzQ0HCb78oRP1GgH8IBnNy/fSqMkZbpMX0q+kZ09/0K4fo+07wQnk
NOFNoz1vmm1PFIsRI2cTPdVvsC5y79s5879jmpbZCclJNQNVXMLDl6BiYYOkqx24M//XGCnTfjlh
f/LLAVRzbb6Nf8AUQJW2hG2vroxqzz6K4Xz7b7L9rW+Jh/9OB6UsjX8tqIjuHp0Ha8l0idNk/WzV
kbyzf7HsLf3tkj3f+2UvlWYgvx7e9DF7X5zI/pYWTzTBdhu/+S21/GkaON/BjmEoaiccOBOFKbYF
0C/mOTFMRii3tnf2RTzb6kpvH8mvlI2Pr7kMzlnFIq4B356YZVIgSW8t0A9ha5C04mlZIxmEALPA
Yixq98quRbzK5Da8OskzHdx7LhfSw8/9B8ccRkc+DyAndbTWPfM3hTdcTTCZJVVt3e121FgU4b64
OEDRPbc8IuTb/EwjLWzk+ImBJoT4Y7SsrE++3eyBPcgTIF1BapJVNTsxrEaXe6g2fSAlzhH/xHHR
XzkIy2xJoDRamp18glyByb+zNsz4oW4ciY016Oi86NVJUH6tyKo+9ak7i0SEmsOwmV1hSBEoOIe+
lm7CVpL0FFdih2AmUvzhSg0l2ujIgBQd+oEtUrCZKQWfcmrsiWdn8dZP/B0NiRCnirg6J/MGOb8P
8nSs6FRuQvX9R2IQxN/B79Wke+zqdGxRSi4K5uzitW7fein8du8V/JiSDi51qaZsen3Q0Wka5VS8
jJxYStDVxOTT5K0/k1ANKfVk7+NDEoRpyyoVSCwfIeJp5Q+uyJwZvFbdeT5ZEWvUbNkQfyefaBbG
GN188EElSzeVSMcbIts8OzqoRaQnMcJrRPqDGVKhd9bomNCYmBHSveROeNEILyJ4yO/DCVw6mTO3
YxjlDak2Mpt7UPLcJ94MhPegx1Za5uBaa0ADUG8K/C8317m9iwOo0UD+e6f+BxoGWcKTOddquj2G
7NXKKj1V4HmlbC8752T8EnWXQf/kj7V4v6mOxi1JSJD/vR5iVsgpwhy3k6fOSVBBLHKnjWCZ33CZ
qzd5Xx9gS2dN6IjP5M5Mj1E5myWAPtdQDAeKFagAeGX8/jzIXum5UUaLngN3+haM7i3RDomfLdsw
XdlWxOV0alW7XBN4DSg+R2fMWbAWNyamQnjXxWZP0hWe/GFxCSTxEp8y8xI4/mlh5QZnIPXHfkny
1NnELjZnMUIApjZqHQc6R1Ryj71FizYBa9N0fymyPSCR+VCUhTu7qnIW2SXIPTlV+W3CB1WuBO78
YHKBRODBtAvNk8tjXv+9AM4iVAgH1BmcWI8ibZmcboNguHIfMaFJo5/fMvad+m+txnLHqK7kqgg7
Qc17vH0K6VXzS8qI1bfFefMBYJ+KttbKD/r/5VIBid4Zo38xlaA0Yz5P2zY1DPWAvLK1MugnAnzn
CewpTxT7zC2u1q46ouJdiTYBYNRd663a1KVUeCUNfnpgFMI6u0A5PLoLGSCbh6VdPjZ1IEmky4RP
cuvlN4UY3sk4t6y0yJ2I4pGham/2Vc5h/s1Vq/aUhiHxiMGBTZgFEqySnzK3k51QqPCfF7Uoy5yZ
SlxIbEgPsOBK5vQNRP7ZAhH3+gLYGDetu9FApu6AI1XPh3J31q79hVlj34HKCgDWbkLxCKp3TG4E
KpQJX0qU/Jkn1qmhCn20vfxrHIPVaoBTEqYGQXxuZMUbgkeDEohpjV+PfR3u7StKEN+akm3zTsgc
rN+p7AgEaihP5Rn9cthdXQ21+Am0PMX5ZkohedliT30lPzZ+f6v9BDMirIBPvBaKQgnJilLQEd20
q+fBt0yhhGCkEHFqHgLSVu4IiTRMNGndyUsfjAt6HCnq4mLF5vc2YwGlfqcQ3uPohVCC3Ogc6dNa
wU6hMlzFB++iEsW70o+rLVwP80NqFbi89tFoQRY4fX67pexTB7SGfWbeyYTfFEPVJGjBnmVsR6EC
vgHek5d9SvU/vQA58FK0O6BcGsryaAttA2lBqNpKf7dGfPuNfIaoZfLHk68EztZ0Rfp207aVSRq/
/dF95qUkuIUT8muKkEY63bNJssYFHF85+6/WLw8q2WpjaXMOeyaje63bW/Auz6zJgHXcKhK16CVc
tiyU1KbeZ+ky/FrqjJRUpOtyDHFppVaEd/AL6Hz/4Lm4rTnuZhOWwv6NDpYh3oNHGeaGDBgvj0f6
goKrlUX/XpuBngr31TOiBmkZd1cF2Si6unUPko3sh1bNIftkX6rQBYUKSqTtOm9sSrHsNXuYgXsJ
pTYg92KQ37oEXy+xlh3F9AyvBPVwerhagiheuYof1lv3xCKjUhxTNL3nGJke9FmKhbssW5LoUICx
p63O7U4IbOisrVj1x6Lg9tLZa4EAB42TUlKGnQcZzXbGVZ1QX9yCyR+3XFROk+3HrNQWJqkrx625
SZqyBFecFEx0X7gx6BOkWyUERPtjTMO9keYC2IXNUAOVFyD8r8csrmnIFf041HSjpAXCdMzbcqI1
2915mptiapaYG9194fpGtf9dPuQrhAdcXjE4pME7M92grAycQlr4CB1pcgOaPDrvnxariP7RcEd9
eqo/wKjIFraxFX4fP6hG9huLVIzEH3f/Al06ELBNQDf0sg/Qq8nyTp7vTG36IhwPMK2qtKLlVyCj
AA6E5bGXe7d3fjWTkDdP4pWlGHyO4FU4V5HgQTG7aTThHXQzSXZs0V7YE56G+AWgdZwQ80heDUQD
hT7Ckb9nc1aMd5IKUwusQ82u4Vv0jMpyH7wftwlKAb69b8954EYPtoVXyTdkKlv0KxWdvTmO88Jn
OduVJsC4DKkvQe84SSfnCPprB/xoMHZunpEnizHoTyj2YeE4Rs3/GawSuz7/XWLch5HZHAQncSAO
mWlB6HY0xgELGzV5XuuWhJhGqhJZjxJoXdeMBp5g3mB5CvAdtRrgdTD/XuIZS969rcNSgQGEPpmu
sK2JEeRJeRaA8ksG7x1C2MsTmeB3j408nieiXTbMDHwUBXGsOn5ORjYziL3N7L5+xggf6qztYRXr
3l19ySDx3d3AEu/t0Fd+cMdluuHCib6bJwREgS9AdHIkS7johDqtkmYpGmL+HUV6X62rdEDa1DYP
UVux9cLjeXf9AS75Vjj1n704uFQ736Ne1Pp2zCtg21axTf4t9fMMnZO73gCI/Mc9B56F3e3UvKrv
CgfhDleF00rNfBzbZwGBLnQEzAowDpVAD3tW4KFd0iQaEh4Ran61hyMad1Y+Kyj57ZsJVJeorEnN
fzbpBBoVwU+PM+SQc8+rrCYELRtKYH6bMNYZ6JM4Vtv61hSwTsBMl28D/LoVxXyAZ8Ha22AN06jB
GYi4FfqAhWlQXYaiYkxFJ+o2MA9AG2h9/KqhGiuf14riD3sCqCNGm9qajEptjnebW1MKVGnHP0r9
6WRh3WS3UWXkkDDnxxuCugZdi9iV0/PaMBP81WRS9f77tonlignM9zBh0IeXQP9U1u9dY65SkvfN
pmvRazj4nx6jM521nNX1ake3rmqEDJu15XOSZlzaDsP25Se+PykNlCy7R2YvXLlUXIgQKJsG40EP
54GXS2LYe2A5HErThUKA7PTw2QVpF9LTbkBW1QV4ronrls2nEIuUyXY5425aJXz1vif0guGrHUk2
eQTWBcepVxQUAtrpBkvqlMggKnGlP6A3O3msJO2qP6rAkX9SYOQx1irjoiiX5SrGDgutZhvatYmT
sxohY/ZumByXMJ8JwshQU/4W6WU1GaBoKPKKGyJgFbCnRkwoGZS3mPsPe5yq5ArJVyRyXs1b9sD2
TBm6WQezpYnoXocUE5JKyD2ANQMjxBxl/ked5jyArZ9dE/MXEmRL8ziZ8xFJyje7XyQOqWRd5qbI
IOcHJNZkBcLRqN0aq0pk3pRElG5WvYgnTE1WqGHM2plwpQzQlY/5Hgi/aJBW934sRP/71CaJeX3P
8I+MSukPX/SVVlfxK+78cj6cSrHjLQWO72qETxdj4nVJ/smr6qwe/hGUuYEaeva02FXFwxo3i0V7
fsbqgPu6OSR8a1APC0UxthA0YoW0Uwc0gHW7lmgxpEmeG6/equZqHWlaGDNyGKm0wxxkYDW2Phtc
1MvotqAC9rUs8iuxNM2HkEoZ413zSY6dLSlviq6M56C8Lu8UaKPMBAISWjLAAi5NuuXfTga6dZ2B
qJY5geg5Cy4HZXih3eu7g8CzSKsEtVeey2SdY1B2tMXP2hXNwcpq5PKesUtiPOVB+EKq1NFtij6r
7wlalB64NdOy7W81139sI5zCyFOJE2LSkJROVr36Q48GKWQzwt8WcrQQYP3mt5LTiRRbn8YCshee
tyvgN9/kNIJJo6UqIiIeJpJFIooYw5rJzKIiC3uHEscNLuBJTPf1SMcjrAp4bYh/wCvyNP+j3trw
/cN15sS9ow8G//baIgUgPpO3p/PHUOlklz0zLRz2oE4lUBQVtZQSlSro09dt/LoGuYQJTLMNY6jp
691nE9oHZhE/GCX9MCBKFi7X3nFpKLgsVrLJa/prwwVeKofPz9wkwf/ta9uearCG63uXyvuD9jbu
JUqd7DHaLYVC9lPqsbjoXvYsLJi3mi+jxhvtsb+GXw9i/R3XTfArMS1NtkcvZGBjPEW6u5rUQLid
Jr/qrl5YZaIj2+ma9iiarvG969/Y0giOYm8iVp5TD9SR5Cs7DlkeovibvEhTY+F0KYKZfud8+y6f
XZsjVVLHceK0yCysi+Bk3fd91IzKmZXxfERKkF6fNIniDIlihx9S/p5NZV7bW5F5ZIjThrPy1yzZ
zTe1hRHTO3gqEQdEJ5RhQTvpMEyz4UI/jsVumUEj0BHpv51iR0HyeHTQerxDhP5cSAPXFiVfD8fN
jtb0xi2vreSPf9G0Zr+X5DJ6gtF6wirnkm3W/erZjRgFfS08z1yyN698yeVILsYfdHXUrYWILscB
yqlY+N3cQmmX9RxL6OgLYHNknHu7hlmIhA6OVZsan3CPXnpTLKzv0CJc2D/Ci0FXJpag9Xfw5SfF
vWL5X66znl6S7v3BVhFMbaMkuSm9zpaAwdvzKGxx5ebDOjrr4EYq1HtQqPFtfDtTYwueKQJ3pntS
9oQlNiuCnxjD4urjgjIUKqNQ7lk6S/jM3mLTfGd4Or54HsDpzD77lxXix/9w73GL2lBXdOrfkfnk
S5wUUybq9Ie/yKWHG0gNTKyWsAgZF/l/jjl6/alrNbMdrJY9NeSUXCVzTrK8SlwTktdLaqvnvkyx
3DFV6BWGivg3AcjCyBaQI0lGbuD/SRwucz9GdjgicwFEllZP6PqpNV7mxmExT/JcF9+Ebp4h3hbO
iGHiiTJCxFB2NKTVf3w3Y8PrUr7+2gMOrBh/Yo9Cu6Tah3Ze2j9+POCgS/IRoidnjJeVqMoH73Y7
qXU5AgCVkSB4r7/YiwJQ9l21W0w3dn9FaFcGcQihg2gSqqs+D1xx8/ogPEmXLmd45unVkzS09Q1W
ErYlumksaJXfZpomRVZP1glg6acG4SlT5tLl02dIYkVOx7Ok7nKNDlLYxQK4buQ7qMu/5TeyCYNp
1LX8RuJlxJt6ep3zUx7Wy2PCjIhi82/yjzqAPJ0yHyPm1NNEYjf+3Q7YfWBQIKuZrnTurwftmi/i
kjpUpdgPWpMvL/bNiQhDBw/5bfVjDCDAqERqjawSB1p9sfHuX5yGpwyDCg9BWVJtt+mAztVIyMRf
1KPr/QFiRqhBv5Ngcnu0eCP//Q8uq+CQezqACKW4nLGwmglzpEfyRgD0ktpnhzJMRyZZmByw5GEf
zyJMbmnpPPfE2tMRYtqfn7wIUlXr75JgwbioihLxCVllIBCizZ281tdMxp9U76i0DKzb+4snpP0y
Xeg/Stcao+QxvDEcDAj4yxc1Xkv5atzGowJZ2Zp6FHe+MYZJJvYE7SqxN7aB0+YwvTYzPwTx5ylC
54Gl1xrvi17jmUeD+S8Dslm9/12a3yIJoIOHsXoiUn/u1MqLhmdDZnt7fbDxY7F003jbZvIIgdbr
/5UW07bOLxe/3Rv9J5wKjL+zjEAQviTZQAdZE0zxPr9SvbfiPA4aPB2w4+762uNW96qvi5cPs6uu
TkuBj6YAiJBguTwYmPrpXIS3j9jdwT3HvCussALmrJBpcvkmxFEcokimChhVM1AjyRzNOsyiQJfK
OY1NiiLMq5tQrlJRGUuRYlPUWIiQiJv1URyU7Lvl9V+V5kEon6jAl+6byvtUvBRx+hIZx/yUOB9i
64T/4dxeV+rLJHeDWdfCEJiYif+4OPTx1i97gzmqOXOraIkH9m4gIZKz19NzMPypBldX3Qfcx8aK
p8V+RSHItorXtoXQUsFmyLcD+Xn6AdA6lJvd2eo6rQ0nSi8c8/PmboBeRhC4BcsN0QKAzUCNBwHn
HGPUl/jn1znarzJgU6u9gD316od5IArjXqJhIhxI8jzmMYWEyWxp4GHVFAqIZWEZUhrmHwNRXi6H
2ax3WN0a7Dmg2qxnxUREX8WQBGMQun6YJJ24ZUIWACfSpvK/dYt1IUA1nt/7RqxaIYHDzgY9suTw
f7r5hllf5E/x1H5XfI87rQky88PjAjN67cJDC9+5QvzIzpIIS9W3KASKIzzW3z8r+g8sU5tqTK9+
w5WINgVRGfbyRiJYdQsbSHlGBZG0hQa7W1Vh/zHg3x4OZtM0/kbIcHh8AYSD4OcFr3db+IHqFyWk
FtVVVteRSQb8sKKLK9dnT0JxmiAOAqy8/ngliHMxJoXk+758bh5AjRhJnza9484TL5Mou1HpL9uk
rzrJq3iABZK6VOy804zvBGLtp6qH1qHW7f4NSZkst/Owm70M/zXa2aSWGDOGe1n1ieBdZPxjEBjP
hApzMZusoD/Gq/d9XHhgvtoTQRC25BK2DV3BqV0AY+ojZXS3ZyB6y8Hsv62uGFWUb6s6u4uthvbd
AVUeGaaU9yHbG0w1wI96fgSlwCY7S3r6syFIqvjBvmwfMPWPQBrzkVY8uZ6NRaSiOv5RiYdZZVKQ
67pRg2V7amGVPSDWHuKVAdyiCXGZ2Q0+JYo1qRoi0oZ5aCvyJoS1TDZP+hpkhKpnk67oEYq5V0WJ
z0YPW00UssQ1bGYZEvgp8Jy+Fbk8L7vQRia+jPatNqMApRygNcvfi9R1LCZmFP/oInBlG299RxLb
T613n+pcRhZEXnw7LqHdLDHdN9q7bzQVp9qHvqvvIrBMCvVvOnPZLNpN0pP6SNQ/K6sqdra0kTJm
c12VowsVESKaskXXDvjgGVktdtKQcEQ/tdM+ESYUvDQf39dveTHUAzYFyRMd5/f6Iz9KL3CoG+Xz
JehqKovL89KFw1X2GlxVuTEE6qzIcRvo7PbPv7s1OmZiddeXeL/ZY3c3RKnAO2njhJCtgzqX7pi4
MnkWqGHvxI0nVAJ3wL2g++fAT9ywFz3q2WHKog2zL7gR3njo6iWlzVm3wiCPDYcPVBDkY3OgixKD
fbcPEq/sKE9EeinVC+ukttpkzYOEcGhBObSqH9rGcpmhedGtNzVsREbNRietp5i/0PW8XbtB5L56
0oZd89EBcI4hCU98knFirh5Jdq7/yjBHWZFtAsnv/zkS2pXstBXwX/inwEq1vVWR8l9qYLBpUFDW
xeQLmVU1GovPxyVzdaSES1Lui68FDvct2QVkBsfu6NlMaxlyKjk4DhXzn3VFdoZ/2SqSACg9f6rn
c65OVKkdPHWumyc3TOL4k3ezd+FpgwhbSU7jjcZXV9gVVnMaN8rBotKY99wcnfcZv7r/F0eGtKe3
/KK+CA2b+mtXROpZ82E+HeCnjKwMmvCRTtm2UEzOYerAiOKuXy5H4py2UX7D/kVJRFGMzNFMXGS9
casqIc89WUQjo2wgeLXNjawe7+AfCkhYypeMjiY3Y8U7NPFb2f/iqyxSLFd+kaPRssT4vJTB5DjI
hEvzhzKM5CJHEJfaOOTSijIlioMOcaxFkuXr5qxaUWvf9kpT9+uu+zdm6uqTCVDYtYND7dja3PkT
OFKsctmRMW4mbzFCxwuwyKDVtPDKVQkB3HuCQXJQTIhyV4IvW2uaBDp3NMwiYXZKMnpGrqQXnUgn
OyHZJv5ms05lAn3hbb7Nri5NIDni5I/uvkAm1LXAc469nZG7xnjNUIQ4WgNx8Qe3rJEOgVhiTRxw
XA/rRvDjG+WvP+1oOSHUAxxlD0EnkrQt24DoNyBaENtpkTHecrXRewVOA/JIU5RQ7AplUDVabt+s
ccMGfdc9juS2EIJBz6gdf/z9MdEgBXcdbZt6/BvmRJgOL7aTVAmOlogsYx2sit9yCdvWPoeTu6qt
kuDUKG5cVjhzAUetbzvWWyiFTeCujruoUYJuNE5IVp/zePw9lZr9J+Nlw8WCQuRCiweENv4/PbuD
1mPkvUMHIxqnoJcIsQsrO7g1EKPRVt8w1A+vorVeYVB1EwbcIEG+5Wsufo+COj+yIXy5nQqtgaG4
+OCJ2ioEyUBSP/cPLAlQkKYr34tz5fgl7T6/D2hsO0T/oVBpQxijDUDks3hcwWC3sWhklHp/gw6x
Byb6XkUQX2IkdIX2sPUHDWc2geFgFj1LHMe14TAWivXXVMFNl2fKhxOcWgeZfL18I/0ob453VwcR
4WzHphMw6J9U232drFvvCDzPdE0Ixyfdxp90/Mb5HkVsIQinGYGeH6LnA8vS1pu5xuSnU/tm4dgX
+JVgpjocig1v9tgzenDtjQyE+2GslvoMJyyuSxEOdygln2WJV+xoKa/sh7Qx5HSMGHPIpDbNxNtt
9hWPMnVtYCwK/cYGCvX+CMFXx03UD5PU7oUDlLo3s1cvtgOaJFnHgNI3ilWt6/SIRjw3zN2tBoZj
QcJkwuNxU66z/RKvGiJ/QCaJhBn3UrZOqUSotDCGDNd9M9IbW6mZTlPRo2UDZd5++sg0dcIlYnZ9
sBDcMTteDNgAtbx3y0iWPNbsleEL91KbPBFLgVJqygOchduz8bInv0AsOKZjTzr5FU/517caU1xH
aYJ1p/Pwpw6eBkBDds9pyZgKrZhBjuoQzDOVEt0USDHRzRxLvFbUGO8eAGyaeu/yO81X1VvQqXoP
26d/8pdZuk8O7JsTht4NwuxK0Y9ldVmEGXd6fJhSJ8GL2X8P2tmmh++wD/N/LOG8ZhLdhwyfWZFC
E2t0MAHiPsP7BSpwPwHDItwuiza6hAETqnl+9y/y/kGcaQV9xg4Pm5d5u1nLDkQRve0V89Ifl3/z
xQbRyK5qOftZ4VZJc5CoJV/vHbrn8tnpsBsK2aO7z/EPDrSX17FmvN3DI0LctvJ9KjpJB03VNlqs
cgkTHPcGbxBOpr0qPQtC2KAVZEzHdguW70aGmaZn5HBCjWbcD02fx9Wjw/CT9M5PzIM0FGyxkZE/
Fkgt/8vybdV0utOApZ/EfmNysvH/inst27oLbqP06On+MXF5cgdXjY2uP3mCnOoDyQ11VeGiKFCz
SuYhtcpYaJMAo84tU9+kfw87ObjXhfSeaDGObftJTGO42Lg/Irts9DeMNVLSaNN7UCsFLrAM5SEy
nBeCoURSq/vJXHtFxslx+17BTzhvAbi26zYekyaI/TiDb3X1zZe4z5T9hlTXBBedMhfTYjllMoKg
m0YYLSVxrB70qBEwoeBpfwN9CaglH5W3OWashcGc+COyeXyfnmvJNDNvqv1z8FauK7HNAdYH1BE2
wHB0WQj3iS89LjpYaq3JHjyK+kgRHe7MpgI7g7fOZM8nHH/9dctdJ6uUeBW971tPWn/c3OgCbvtA
Rd4wtISA9FNoJm1+ar/iyfK6/rh4JFNKRD/9I4EwONGCMVFn0eQItlm3SSvtpm2oTlS4tFXdUVfO
v3QU2b2YUvshj7YVc8JuoN+02cDFwMrozZHGAhB7oCBbauJfpRHe6Cb4ehXgTn1FrB2Yi+mfLkZk
EiplvgVo9pTk947ssMCH2FkQYgbREeqhQAvCYlX9hiMD2+gDLvPonIDOnuyMYhC9824O4NRrzTNz
Q8YpD79FgWm/3Ujgny8oFWnDKpd+p183lDf9It0F0SlNoZtbdi6+rUPEBIlAhD5XyxQj79yOGOvQ
+/7JI7zAtLgDIRvZnstgXivKV/KkGNI+QAMESg8WsHR6dQfKs2XcSM3xw6YY1JiVYri8enfu6+AQ
l/cqCR5XvaCtN+4Jp5Lcq0lTdcvK5mG6FcJMtTS8AsrUe1JWAR7rpGKWfs50M1Fr0+3jYCXGfHaT
yEZNeU7Wnha0fpbFwVQulrRXK814JmbaMQSTlpHxERF2Z4LF3kn/Sp8MGRl31BSrsyz8NXTImhGJ
lDUD+jdivQP8c16i5anqg8Y+WKCGbbSkSlJLiINEPt9aj6H3s67cbx3lFr1+Us1iPix5dX7Aasi3
J0wHQ+P7GKwV36nMVtq6li5zx0LaHL9DN9aLiPo3QObQH6GUs3zU82d7k9STejM1QluspXaFPHHt
EyBb/jex2TrbaHff8tM1c0+Npz6dUrBMywBG5tXZE4qN5CoBXA+5RwGVhlx2B3fIclISXd4PKY5t
UD/A/8CIpen6na66C1Wxkn3iRWM4FnmHSbVwMHnuWf2lrsUE8ywQ5VyS3JO7pI/UsTK+lg1H1qLP
coXHQI66W5Qcd4rOWV2zggno+mE0uPqv/p01/m/NLYmqA7eTYS3wwuVqjai6+Hrngz0ONQ5RSatT
Lna+3Bm1qTfzIjovwi/JUmRUx6vPl4kxGhS3CncfDO6lPCvZA0Tu2yObE8wSLGfVqii6tDr8PtyK
aOez3T/vOX7R6lo+qZRatn/mQXyW3n/pV6jiThuxG8j0dPM3W0nXw1r+k/inxWozqwYu5mc2DkJ8
LrBB1j/HfFyNbyKEd0lfBdI8BFXC24b9owyQzlaEUU5PZnMRh642akoi6MgzzbBUgNAxL3RQ7PWb
7+qKGAe9Qf2M3FbQona1GO9v1fBfi2a1VHIM2hqAWVpc5zj0lBb6eqsmrrWwjP+rEITbcxhOY/p4
yIhFfPkFKyZ6+kj5Gh6rIPkOxnbycskYsYtPOkEBnjYe9G871l8MyytyIE766xG2QvqRFbR5ruoR
qVfhAM3fClFYmE7Fo9bD+NH7IF4yNanqYaHRHt/xLkEZSnF8eaTsvSguTJ/EpqFJchkCuu2NQVZH
WN/GpQekXcNf1EZXV34zVCysecTEyg+3MuuFmf+W/HvI6VTEBAl1up1rF8hPxQValgcXb7vHdg9j
24/PzL78Chq0IQ0CmwN+Uoo8xOEbYDaMGgiwttYZhn+3pMRgU4/ffIp5GrNCrQ/oUPBcUzMdJtzH
SLivqw/BJL46oHPp8348wLG/OeaZPjL6xBaNAgSLjGLhTzs84yx87uEjCWJ0w2gnGyDem9SxaZyw
WpV/KoTrzWJxdG0HZYic7HYHRTnEu8MNCLnP956bnaYbprsdbkvYsL2t+oYoIQqdbT1sxJ8AFZt4
0rECcPsvziLLd/H1ZbRRlI68WNakbS4MYVD/OZCS3/OsLqPau5JhDVrPeELDH6i1kJKTgTGYFzXf
jBcJzEKYo/Oes/fPqTaAu6QtJ56IIx1BqSPc6Bm4H0KMJZhAAY50RofPvDr0tnQdGv73XuxVFSEK
LMF2RNEJ2l4jnHNpN93AEYbL1RmLjWr9874DixTgBsj/NQMEgEuJfeRf5YkaUeNiDGpR9iAv5nkT
B16Ca7Z9CYpAGFwLJaUsnYEdD8Wmyd+qwshEhF/0VOy56SEITYU0YRYF28U4+2NLQWn6I/mnuWw9
jGzINPG+xw6DcSAtI5Y1Ion3tGbsqv10CMpcw98bBkhQ5vakFd5o00zEMwZOR2B1viADgwWHZRkR
xzEu4GoXGartiYfi4AGuneu/2aF2Vs6ohoeNJQS9Gd+UWnC1zQ7nyfwjV8ZbinfGnGR3qUvB3T7z
vJjrvQmmNq40AUwPI2d0b4WxpPmtUwSP1CUqpFiTk5rSbtUuGOZjVAs40ALeDAzuMODYDnLpr6Ve
lbAAztVLJOo3p7FJiMDcb6BiNBu0Y5j0BgmMCsII7a99u6vqgJPRdRFmsbOBWsLH3o656U96Zsek
RddeqWw92/DA2B4jjFrx7Jeu/JVtMda2Une8XSa4rkguQVTy466bJLaeXiO2L5P2pmLzjBxnWK32
JNPAbp74GfwWVt4OLZsmi1Dxxc0FxYsIeL36f8Gppvq20uYZ8UDI7IkcUUj/Spih8LXMj5e/2U4P
yzpF09wsuJuLJ9NQ0aTKMc72bOnSrXe93QViTkmWSjK+KUGGjxo/LfGeVhCXU/sUwip6qim9MwWg
yvElEXo+oJH9uieJ4kTxg1Fb2nX9M489xh3v0/I1jvNsNqIxwMrz87h91JpMhNxdl6dytcPfgWSA
t1zYI+2LI0CfNSm74qBULVIyaogP4ig82ZA+ZYpoB6L+JSR7k5OyUXWvxrXtMf+ECN247/+tjeCj
4gR4Kgaey5iGljRTWGYtWlE790WG6+R6LzkJVV2lvJbYRToE93yVMo9Z7DLMc9Yo2LPaYFt8ea2P
jn46tY91CrU1VmO3CU2Zhn1C/t3CN9X718XNkFG61VGOsdp9268jkxeuFyOJNlvlyNkwgoOVRqET
Qb212BIJ9Wz8ZpcbRXwYyL8GC33MeZ3g0OMtdZlRTg8rGD2q6kN0ITXUK9/9vlVoDM2iQb/F/Bta
cQcMJtw9RRmOxRnnDa0ZbvmOGM5FYKVwjP1/kc2B0WcCbMMAAt5fOgC6d+MQ/Au4y7YzVtGLhLwB
zrwpZCCJIDlJETGVXUOJGniyxqi8pJZcwknzfNGo+kyssFxgRSLXWgWa+3B01HYL5e/leoMtDHED
KcP9jczpXoHihfw9/TIrmytE7W/4FWpRmzmsfumDCgYJcGqOViqJSSKCmBdIp+CVX9FIaF8f+eQP
FRopJ+1YjwiiUOA/WDrQqYYhwfVKt0teMfmBEjl1+mG5UmUMDDteFvB3J0nWDKEerTX1dCtRMQA8
SDwryjwjbWj5q0H+0S1wfOVskVfjEGtkcKKinh6TEjWCW68CE983rHn2df8aIL7nHaIfWvc/K2nL
qGzv/PQuhDB4vK9PwK4MlHvzWqXbMJppKpOtw2cXHmFT8/f/nPIwbgJilHph/Nkg2ZnvhsdmkSUy
HOgGui3ObkcOunYE+Zb43vMyUc+6SmVUGYBpnm9kE50YXpC4mhDkmmncLK5Jv8gGCsW202/GHHb5
puIbfsTyT4yZFu3Y8Zu2u5WJLC8/vteG2bOPKIyzuopFJktHfUMntzgUOpru5Gpg3eVO/sIqKwht
6UfwXAeIKGBO3aep4WCBmzRdOYYH3EZUEcbxuNbmiohfGYeLUunfgpFi+sQCxEZsEx3zAKqJyRjP
N7o5ZWQE+P5/IjsP4hMJDkI+hZpfBS1yVq4Qx6yk5hswt1XtSmnilHW31+SbWXzGuz76LEY4FZgL
xZce01nHKLDZVpCAWVrKOj8PcI5bqrbA815mzuHNpBmcrqBmBDg1T52X2YQTixe28Y8VYIEVZt85
o9zm+ifElWpcM2avF0kshA4bTkt1vh5MPhgwsiviLW+6VUfeTVsiFMmqT4OEbOgxrKi1v1jWmyHM
qn/DSqYvnYyF5ygKy76u4H2g9OQZCZ3wkQP61AjT2IpqGAfrJt8fsmaQMk6jcw1IrEbFzC/i1v0V
RJDJQf7yCyRYao4sN1c+ssB/81JDCPgnRH6dhCas9uMdYXYMOpQ962374WaaW2v55o85sh8wao9L
OsXDzC1YsAc13zn7hjf/l8pLa4RZP0r+cyBDDvlYGMfx0cKPBUVFwRqOvW75tZntIhR2EtvS6sme
OBgqkU05K7ygJ/jKzJY/+cJ387qhuXENKbbkupMJf4L47CNm3jj6HV1uc5NVIPvaFj/ghI5hf7HP
Sz2EIvuL61HMmtqFaSEpa1+AOAo1sCjHQlo82M6DDL2h604MDrYRopqJOC8eEnuNWGrbGfigQFe8
6DsyHLUmtdAk4Dd+pDml9sBAibIczIjDIZVhHC+YoaGFEoCwXNMsFGnhKswkIJkIBB+GbcTtiHZv
Ajn3teV0Ed9oITU695WlyWd0JKEddYilJ3AtCCt0R3iFiiWf9TNJKVbF541tL4THmCcwIdC2YBum
eNrXm+spQWUS44LmkLJARbiYWAwbHfpXqUBfYJmzTqlwhGRppuXXRc5+c9khwBEqK/sT+RI7cO2P
Mvj5Aco53DPw2eVSVTeQkm05xMB6gkiLzUTcWa0G7c6iqX/pUU7t3F8sl0wtrCNDu+M1LPDhbf/B
tJPazuogJDGMhV9UOmsHOkX7auRNtJ6rq6M3M4+9aW6nd15haBFsbvhkLbDnkiWTWcrQzweNx59e
1FrNpqYWPR+bv+XXabz9kOZemeOFdLqAULsDMOJ4nHzAsNVXQ6o+OXCQGymHwLXQ7aJ18KNA7+E8
I8NaWmsXy7fiTvzE70rUMkNHZUqFd5YLEvD89zETABPvfox//n6Z96emJZ8JIfYslAyWhxoOQB1d
f4EBdUPqEpKYsALa2n5mivywCNx/5jInPjPzl+iC8lvmWrFURhIucMcKAd6FZkVb4XBG8K3kQChQ
FaMrBfbDjyXZYCJpzH0HP5Ll2V5Gq07lJhuqiSfWilETMkt7QBIgOjRCwi9jggPo73RXb4RoOhD0
THDO1XzOyTWGc+WKtwjg8RKpEuvLSB1ZG3w9C2ah9pGM6592qQa4aT+C8ys1dh7nQ8t8/jDwWhZs
G5NiTb9FCY1gDRxdM6Zb04Y7bQrGxhs7IXYu46hVHrvwKFb0T0apAVLvxAgddh/VVUZKu59t0U9r
GdZEKEChR8VjVNxwva/vIotYXNWAhcm92rAJBohuvz1ruP0rKlwOv1DUNl46MfxcWZSZMlYAz4DD
wIJuP2CKuO5L070gPM/uQ60CoYj01k614yDpTNBJPlBI8mNiSjGMTNy9tA6WTXJxRvS1hmmFIzV6
EbFl2l82KtCyr5tDGMAhHmVsq37QJRTF1NM2k0jCD23XbUXLk4Dvow296GeRJOWFxjsOIrl9aSU3
uxzKq6W5trHSSbFs/fMFuexITLnUMrJDfb17yAfXymCXf/PJCwr9mxLF4rfM231Ijztg9Uky/6G6
s9G/+N3hlvL1Az16ldsoWtWao/SVyQVTu5GYIFmEdstn7djbgKvLlXXMVTSIjdqZ7VoEhyKUMGzz
C7MPvn6u7bK1SK4MQOtRfWP46ei37KQ8PYgeBuEQNAqD0uUbA9K2JtQSLMVsLPUb0ZqSSGoA0j7r
vi/hgMMnxEl9RoqdbtylSKLmkaTFVdssJX2KuLkF5qduH5nhB3y/kPvwl/fEy7FAIKlGvpSDVX24
aLGERW7Gz3mgwsz0GeNC/HhK59aGSAADeXTwJ0OZ4luOK1bEZEgiWjQTmCcA/j/XXk/VqTcUP+yN
N586bVYQiP37yKeUas9iyt5MDS0G6lpXOH+Z4r3Dm0sie9eWMhDjRWtBMX1U3D2r22LouB9pyKKV
tZMMTZr9iJdtG4lN3khowt2Z4eGmdKzKmui155xJIehBZN5MXBz+kdi/3gNJZ9SSxikM8isIvr2j
OV3MjE7IoVZRc27CfVWLZ7ZxU0TM9nSEICFmxVC7YIQMa0/t47JqhWtBuYBgqKdJRo8oiykiUI3C
OJF6y8k4IePkFz+cHM09l+mVZ3eg6EBi7Zv9mWMPc9dZrc+QeuA0nlkXJ6OG7qwEVTzeDUD48/r1
5hqf10QnN0YIrirJV+++ETcTkKkIbBcpFSf0EuuNXRByNp6XWw5dVSiVxSExnMzKcXU/NmJ+LShJ
14Z/V7DnhX/+IoxDG1kwvWXyzqxiNUymTocQBHItuj2NPTI4/Vke0/ik3rMCJI0IbxP3+gwyAE0d
DA9aosl8rJOkzzal87E1pAbIeeR82K7fDKrmaH6qqmDdJi97kJpXMq+COzoz9Duy+e1g6/FhArDv
uojBKapVN/gfDytr0LcYwlwDC77IEzk4lsqUScMXyTNYxjtmet7W9fzxUuHIK30VZRpodTKMCWak
VCzEQIDSXUu3xELh0ok/B44OXzIeMAHRZLM38FexLIE/nw/dvPF3M1rPBwmXk1eFl7YlfTcoRPv2
8Dp+dO4/MMQcjJOfR2ftEGBeYQl8vYktMt9UtDksNwBT1V10HNU0rkrHMg+TKGCFZmlKJdUK46Iz
k8Myxab+KUgamtHvkm0uqU4Y/YTXZNtOfYj5lB0ch4blokGIgBnP8yPz1r+Icz9x6xoLKGvrnDUH
89n43J6qPACwsWJyX6bdVdbZG/jDM8n5VPCZ2zbvfOHPirwNWHeQW9MuAuL3yYL+X1cSuFE0OwWO
R5S2DuL5uMCfeyeRvNj2w2PYnBpEmrl426BHvHCj0pTR7d9EnBq6ZVPjXFPHLP6QwXwgBDqxKAKW
qOPlk8VzS3TjMBztZqRZi2md7R7O7lsiJelG4eTAhqe90PkrO4SmG5HWi/dcv6XJN/fihjkeaTM3
skiV6hsPd4w5VQTzlIVvEdB3iOv3fc1fj6z2a+tz3+F+OOTHlEw3FEEjHYkCijkgiqUygh9WC3Rp
E3f2AuXTMUQIKFC/28Wd+XYXMDbbgg4a9Wx3L38SFrKN6LBtarLQ/qnYYUIMY7mTQFRRnLRwafQo
0saiTJ8JQfq4C3nhBif9/o2mPY1qtJLXez3dToNHvdl7p2TP8utXi5j1jJmEME1WjM/U8sZbL38m
r3DzBPIRo0aw9MgbSFr5Dheq4iU2P2w/lGcpHpdVfXQjPm5iYA9xvdb6c8obq39ELM/yQxvT+tGq
Htd6OAEBLpXfGc6tXIq4PKLN5CieDRUIqgu9xvCqz91o3n9iV0IbAswABDUcfC4Xa+USzI0Z1H+A
gD6LFl/yJo0BCx67myjw8quz9zcItNHpkOZCCnMCG3oPqd9reNRfaY4CYW8yHrNTB/dUEdxHIZbV
x3/RULtF7WNzSmGt9MuKsSSlFA6TzqjyY/tm0tPoj1zqBR38chpW5JTVo13q9sMQ4vzkPuZmU2DZ
AMw1zbtczbsep6RkDNP38x4KohN/o3P5YAd8fn2uYEdwz3P2Jn6hScrhdndm1YodNIGJFfWiTyoD
imASyfgY7x5WBnRul4eBd7Ar4bkLekW5tq5zeIon69WBIDbr7vr/Ukm3KGdXIcoacjGVbf0Q2qU3
E3G8/hCWaj+6Q6e62TEk5KPxFhqkkm34EXP7IWtD0GdWS9WCXpducpXvoV53ta71W7Jzqe0kmrxT
DSJGn1AKM2rmmke7HxoUjw0Hu4qzI9mFWVHro3QllysLNlM3krxTqtCCXanWcmtOSNvtwIAroQTJ
lLbIQ/hKMZX3h7dZL0R7RhFs8FSWtpm5csDiMJszzaQIeDyETP03nk/dgzruSxTAY+i36aKYDlRO
2b1cvkXCQHH+gvRIzP8XwyXVji50I0bAeasq6E0o/VPSJFEf7jRh5QMnVzrOWSzqUQ0m7/laOtL5
Or9yFWiMuONlPLuzNRsggtS5xErzrGFk7m+OuUpyMJ8UeyMB0qW+EK+jGAUJq9hO+v4usGCCqgCj
LhmBjgIEH63BFH3rhQXMuu7dbv2NRH6SkFGk0IGpeHSytMM0WdiLIQohxhtaEvAjUE+Pww7GWfHt
BGAIIRwMp4yH4IjGJHFEW4yBGyHaBRpsL4TVF6cM5ahQ3Zw8oOgsIoML8d71IL8sVMQFqyupGPQg
fuBYkgBaxtWJsL3oSGTKZAtxG+sElfPcanhumSaBeyfwavuuIJJb91tGKcJdOXp7/kGIJSFs0KiS
XpZxzATRJmRNQsSc6iPRvMkifCpjMjTOs82nrF5Xe0TbPV4BC70v2DpT9Q+6A1kQqg0wKc9McMap
XWmR3hso0C1wZONIQW2LafWMxcSlfgERaYxlO47EE32p/9lm8uqtcyHCom+7UXQSs8gt2BBAJhRj
qEPM1slzyZZFbRHXUo6c6cPOkuRC30zMiW+bzN/+9L+VF0cnlv+ccRcBktpNSmLvHbxmLaEXTUN1
ux1JMqdiZynklM40WZmnBTnea4rUzAhfv7XaDMPTTUsBtFKniIa6H8hiCSKTD0DElIK8hQshE2UY
CXA1/QXCTdiVIDwmPLREPt+XQ/wVphulFCbVxRrBTUo+YpnWx5jccDBnwKBciDGIvnjAna8d6x2p
9fle5cccjTOl2Vu+EzPa6JkpXwVwTTGiEDwB7XQmWNSFRcte0uU7um7Q1wDe22wDwj4IJc1NMw9l
M9WUGFEgVXHK6POvu56O0Oj9VSb8FJ5gQBVACCPg6U+k7QXwn5XtH/DGf51iEw3kcR79L/lusXhC
qw6kZh1ktqiVVJvp1fL8vojacQsxjvZpW5fx3RXAnK2lFSYWrto1AXsNjC4/FTPc8KLzYNHyFmPp
q4ZNdwccCd7M6cX8jRL0zNFzki1qfjIAeBE+bTXaNtN1gr7SHeJaUfRps19NUtGyzVO3VsA1b/Hk
L0cPGJmWoAlruc8J9m80FDhui58fjH1DyN64m4KDleLn087ne26SajatuWZbGGfnyIPm3iU8jvqp
YBHH1LSPjZyM9eD/FbKfA57qKsbOLaYvOqwAJIUHqq9Iers5NEwhbbunqvNxj4IeQSYR/xsrPLn1
wws+YID9mMt4K+3v64AjkgLPdVTMh10A0qGYRUIfnVCE2wdkETWw5tLch7DbBZRD6wnglCbWdy/1
gpR820/eePKbgsQshAXDU57CuxwLFDqdH2/2lkIVHcvEk9YFeqH/XFDGeIYzylGNC+B3GEjelCCt
a7j/Oy8irDk6PXJH7fqKxcSC/M2yNSodl+Ikvi/ODaGPpBMW0ajfBRxBiXlpchMKjiUWySZEiFzY
MJhhsBsOVez/j+joWRMvIxZ3siwGUgCqQts4jM4AtLTuN0I5q8sVLrChLuWTD7LZvS7mC2eCA6l5
3Egse1mjWwQCwrnnhKTpUl+Fk6TzaphBpNVOOHEiBSUJAa7Skg0eWP7Rdh0IxvBYprSed+LrEaPe
BIEaeWKGxs9xqt4jOQlFFbgk/d3UPv4U+zrvctZ2TVgJeBN2NU0bcCS3Q3PLYwJkEqXuqwKpgeW5
6BYskAzXYTb/JVmTLNPXvWpP8msm9Teaw0dyxdmWAFbGYiMRUPFXjt17jG1isaZKDfa4eRc96L26
vnFDlHV8ovxHwF5FURrCzUk/k3I78WSPj7/v+E0yK6qXEx7nO3xhvfhIPkB3EqsKP+wRxWK83vSH
nIaW94/SZ2jrujHgfAO3zk+paLkBiHhIJLFK9sVw2ytTjC+KpV917JUO85knC/chQeVKAbm0VI4u
sZbjaQPZJkXtpEhjO3ZGPjQL8RgeI6MUjmA5sK13phNPoyWNFCFq/hTgiIkQnVoPz2ESFcrlknhR
PfFHVspbz7W3Nyr8oPtlDykVFNNxS+Cs9wtKFOGRsxuoJ3TqtXP5qkLJ//nSHK/kMz1/DuNC530I
Vwp0XoO74GzaN1xV30lszOmrSA23+avGRxkaaWnZqlF1mUoEx+kkkpb6WAMi6iHRqrA8W7CIuUBu
MmrHp5Oe/fn89DW4Qqn3Dj/jfiwvxNtEP/5UUdh4W4FvSHRnIgsi8Sowdtc4wy5izumrF+MMHx+A
fFt4nL59cpp/Zb7yQSxh6RiXjKmHjJs32HLls7DsusfKkAlT7pTiJRJ0a5GRLXH6SDpQ3qSQz8LR
A+FcKp7sk/7PIbSqETLgvdErXzEH8YZ3pKMOkHCBdpD1Y+QYXWK10fMY7oIke4c0V6SbXoexAIya
KEdrA//mFneMIdQqxI6xYHjyop/KogJdF27qzfHq4mqIdD80gQWP9zLrTSUyZfLkxhxoMPh/y1vv
qlb7TuEIYZqlkfZZ5+Qd1JbeTubXylfR6UkWYhlvfLjuYh/mQAmbyh2mtAz6VY40L5MqJ7m9mSfj
Bq4tNlwLOLHi2Zyb3XKPHqXIjv0VZYbkIL1rHUZbCHhIzyau1PiBuMU/klXM2hJptOpCATF7yzzN
d8Kug67lUktmN8SxI+Et8cNgNzSC6UbEmY9SOJy1ZG3IJrDB0VJhd+5gMaTvzLo/KIu41qcq/qBg
jMqvd1mpZbYFpkxwEyqP63PMmyCR+ev4iU32Pk1uVWyKReM+Wr6824pkV5IbueqV1lLR86tKUOHv
eFHClkoJuwgyXxA+zDLEeMJTbAeT0rMC5y5ztXtZfFUPwcF5l9udiycrseJG6OTmgHuQIjNrBeNi
o80PAW+i0oAnQzqemEkz8egRHNAqFHEPiTQhc5ZTBPgqE3zWZGZmJ/x4WUG9jSo0wxIkkXOXjx7y
iP+XjPT6/M+WD8fN6IwK3ONWvZxl3XfTO84Gq9hZEfXmxMc2UvCgQ1vrikS+rgapdb3M0cBtbsp9
4u2G5eLZZ2vlgFwMavroKq7+4fAb7WJBSQOHP4VXjP13RVyQUEfUK7+ikT7LXY/nMq/MGEoRhjnY
cB+FjlDt+W2ibUSsg8vzWWcUeosVConA858y+3yml6cIJ0Zqiz0t/mVKv8F46ZvYx9EmvL0mVhrG
sTqL4awEhvlfLkCCS4f2zh6LqkgBa+MdPUWTXm9Mdbe+tku7d5kAEXo4I1idt5/WIFF1z3OI33EH
zV2aVBaVSDhA6Bet/d+uF2UaZ62z2Bi6W6Q5Qz0fTfZcn1ZHqMhTWuE7W/uZTngrlmuFB6wosDPX
xXlSYS4vSx1533pRdko8/nz1zqAaGp3sHN8QM7rNSfXXc+ySNmgBKmsj30OizLqYZKUpUEbPxaiV
4PB3Zr4OH+4bdtqp0gNPUBvOy/kMKi6FWQ1i/dVYo0NYqwbRP/pPittRHBrTlTIzdQZSGfEV263y
DKpw807QOWLXXBxDnqw348mvHmSSOinK6w2q5v0tBpeaa5D+yPscQmKs3XfRN6AQLlODFGLPuK9m
isoE0tpfu25EjL7fRKFEkdA3sb/vuJjF2ZWrVmpuIahyCzSrv3YCYKjOhrEoo2/q0x9lpNtcec8w
UE9lXBAs8MP4vsw+qJQxuKsTEWoQT8F0pjJ66FOHqzKLSGlDWKCggnfieCk38xNvStIiTxdEelui
xevuSMH0g3vQHmpQF0tP/0y/7UFiKkNInDQrkslmkDftfUocb6jO0J6al2rtvngXNIl1LHbltheZ
CgKvlH1AHYshVpd+PSuHHOKlUznZiEbGNjHWgVy+RjP/S2/u8QbUN3foCy83pEtQgiwDD4a1Z93l
RKOTAzUf18j7llanD/8cp/IkWKzVgb011RblSpgPoJm3rVGbD2tEmTmyCKuhX2hlyjcsPBfmzDQf
+0/OFdcy/eJXD69Zq3b7BJ7+sRiUBcX5FgquxvAiMu0oWTxix6XgHu0mqJhpvQZ2GFKM6+Ywcl5N
mw2z6uv3bBQpk88Adw/4R6gdvHdz4ubWNfmWkRMUaORkOa3ykoavC/Y4xR4TwKd3gyfdaBcT0BN8
yTmG3e0NL6erhBMvtcVhMy4vuZmCjgx/iyAnfc1HMYGOSStTtrvp7x/1U7S6wPSm1CibhnqW/y+K
dtOSLCbEwmbVPiSnNp/f/MSAsOHOhR6cRCIy6pmw6bUnzs8K+dCetUfRwufQM4Vwnhpnt6vaX8SW
mMj7idHqUHOyFWV4/KP2unk/L222wt6Iue1xqluP3FmL4U2zYx4VHMPcR5OLeXQ0YWE2K13SCIoq
NKiUn/SoR017MP16Ybe6rP9aABGzvy5XTotF69iFuXgKgsknqmS+lDDzNSiloMHWzpg99yvZ9dBD
zw85aMokrm95FH96AofiwanjoPFvMyj9jxgoPPa9J3nV+fg/6exKIO8+j8iDCTd4O65qZk+igTRI
QaF23NuldCs3vJ49LsneqtSf+1SmKj5G+Sk+wf4bVfHuJTt/jH9pm8+2vUml4AwAU/mlz+Z80k8F
eLHrxJsy4NtdcQ+ninKb14N0TLlMBy0grAvJxP6mqG2goymx+H8QAZBqSibSEUOQ4UWek9ugWSt8
rpz37W9pFkW6HDSjGd2qpgVX41rPD9Tabpy8Stsip/7vrA1PPO3XAhgObIl8EtuOT1T3NdnAX07V
e/RguWj29A4S5nDpQruIqZRkZcCFCph/EDkaQTRd130tVPGi/fj37flEc5E5V9V4iawQFUjjv6wj
g/pZk1x5tu7fqs1KXitGDzRYYFcjfq3k9h9KWel60+TOeZDAyIDz2HO8cOJq/GE1/cs21eLEZKpW
fV9VP2MCGV61yE15f41lbqwi+ozSo9p7fupFhPM3lsS4XvASW2nnPnuBk77UiVGPX9Ttd+Vm760Z
w+ogyAtpBZrDkYzG2VHky4KdW6KW886aoO+IOaGO9hHp1xdE91UfLHwp0FzJ69en2YbW2CAznzXF
Seak2B1mcaJPUQsJhlslUt6Y9ChJXUZ9gBiQJ3AaewLWPTqiqJ6koh5uvIsymx1p8XCOJs2zI/Pw
YkM3E+++ekzmGe9jFaiRvKX09lJPtolSSd9JOsKlWCAJpMsUAxiFzLIMfnYWYbZom+eedoXjFMpx
dePckqbE/HyUN3F0Fr/IdP8E4VqoIaNamJdBHxXUvVuD4fiEJ0Uep0+mxtt1msCTx/2zvw7Ne5eV
VwirBDVDEsE4f46gIejM/MF+Go5DWr1Ls5jZyH8LTDJhEZdeFbiK584teNbRmW1iEEDKMjGVUysc
ytmY5+Uu9427QeT9HxKsTblLxknDstqzAZO54oToNcbiirTTDTytXWXNPaOC6soXT/xiwC3X3RsG
JVfIcYZAJ7Dpq8uI7ce1hyAQYPMCM3iUqFOcrA3Jf5bHTdhOzk9KUkHEVhc9LsppsYiwujjWyVi3
3RWuRvoK1ssIp4+DyxcCZMqJZgVjiiO7zyYweQjFOizSg4cYCKCzZ9Q7PyK85tRpxr3xNuDPffsI
155LMe9+seCwnuwmVDceadz+dL52jApnjJ2xHQqodJ34JdIlfgx74pfOIbcUPuiWjBnBaYIZ2vxe
bl0ogwRuNIDG5qW+zMJLt73itoSacshUZ/lYuhtg0epJ98LSMQee6RZFVGBGMvGq7oM231cI2TyX
mKOMIjE58QgHmGtJnw8injOkJUa8zKZso2Qtg92EL9w5YFApm8B8pl8Ml087GthNECV9+3aw1bdt
1C6pNvFyablTOxrVhbpK4mgy0LaIt8V5OO4fdvMU72cELsOTN+KZdRqFBgqKAqATtTBKRrVbwpGe
tIAKU7rP/sil9SvvZqtqW/GZ2YfihGepCug8ZN/+4m7X6CaBGbXYkWUfsjvBFslEG8xT3raZNc01
9XtXdnXZxb3MR0v0EWnPo6vj2HEYam9Yt68V+vwUTJjPLofo+PKHkGWIMjhlomCmNg1zQTzerlAQ
8NfDETMYRlP443MjQYrn2YF23Yg1JIaVXQlVs22Qk0wby0/cEnjOcixWJTbaN7KgO3wJwL9deCiA
ZdU0hMxIgi7Y+Bk+Oytw4Z1aflDebxdGDkPf9ClalWQ8RF89eoRBhE2r3oV4JxViUouKV1Lj3xya
GeWq3ZoCtG6aVU9Fw86Ndq19/UAOLoE3WUPEiG6014yZxzG37qd2fO5imZx3OUmqhVYSxbMkab29
vNoxBQ06Emxd9qenOp964N/NG3ziombDib9Zc8yBUdeiJfDyP55emhSMq+OWuZ2lga2l0aYXtw1q
QUUiel7F7FlsEX3cQjS4OxLXY7pmyuiVHpuXJ0H+0lZVfiJc7idd+JZTjtoxJAF46Z/KorzlKebZ
0DhdC1GoXtTJfrs332VVlmymtaobWflxDiwC/17KOpu5ic4vVNuCfvNF4u4ZH8DruZb2iIndvRcJ
QR86YXxT2Z542tByO3ztXYJ0hir1aYY57B3c3W0QM5K11lFNVG2ddvgEYl+UW5Z9i6phnJW5P5ZU
qa9DGolASpQ6VQ5qRe1JE+8WzyoFXIrJojEA2mMtCdYk5gHUMM0R/3Y2OS+HhjgCQQH8q66N1dv0
a4DB/VFTnaVNp7vc5Gu7eS2idEl1v7SBnhzbrGG3wcAna3+RCxqX4sN5EoPrghnO76470x1OEfTp
09/0fbFwphs7LtXuXxAW2YHhEoaCntdOGnC7KLJxXNL5RCQMYCl3qDkb5+hwI8jdcgrNLcGkHAfD
btyTPrE1+YZ/QtVJxLNa6RwEShbj2iCIP5ZXiap3OJSFRMfbFagKmB+hbW9/Ls41APb0tmvs8n2d
kcFoPBWMwyBOfGhtGOaW/NYYc3Ibxk1ZJDIqjVNqDT6FjsqgyPaAK39QsTwYGv1Gcsn9ypFRq3Jp
/rAhU1UMOynM37cLpPpPBxbuF3JEIyt5vFdOJXbUvzkJYK7hcTTinhtOULL2fiDCiXVDzAyMuIUd
P7kOzgEhT8yLwa5t2A45sm8kTk+YL9oZc/FGuGFaxESPSiGxuOMlB2tDE86ZyF+cJJptU28LtVBj
x+TP7r6P5RysE8mZs4XGaJhXvI8gDWlnJy34nxfo+OjQ/DFhcvA6WVHxrZN09GyR6kXdc+EYaL9w
L7mtXdK8GLyV0nPhbLrzb0sssuV4HKuOqIm6nunnKsjjn7EmMVxW/QwdbiRvGV+iFUOyyo4Oimwx
D6PcPt4NRBDDuzBSF1ejzl+hIs3Yt/aItZEsfB0z8QdoTyOC5LVHaxAYcG82MlMOtsfD/Vyka1YL
mGygL+FkEhNiN2WHAtvy9ntnZIhUEEf7o3hb5fVEXdIVb4kw+YWyOxAzQad6bTKFnWi3fII+nyYR
VIIrwJHtmCCVqPJvyt0kSJiun4DMs1tGcE122Od+5NQWA9TLFUxh2QXhhz3CJFAjP+uoHCLXIRWL
gXbINpssWu+enTjXtY9ePCvbG+Q/UImzhNOhqa6n+uqXUvExZoh+iGez/LwQSP321kaR44a50NIi
KX8k8LTYUMIME5OFSkmpegzDRGnmv1EtNtMSEmikh7sWVR+9UhMecZd7FVwHN2sNQWclbYBwdGQU
b6GdWpVDjh23SvChFgKZD3TdLFTGCBDt/lXDTaCBbrKpuc0a5m+xnMn+2KM3oYDNoJEasFi0XV22
fG2YpeZujs+d7wEIZI4JVgIuxPdbIV3kHfp/an7YUls56y9Q8k9SCO1cq/Fvt0YONKAqM4fPLWjI
4yeHNBxOeWl5pIREF/0kjDqzraZOlSZZEDq80dfOlrsotu5iGiXn64/P9lsIhlCifOAhRhtl4Ku/
6jpTlUNrWBYKhBoHw2HbbrC02XB+h83yY2x8NAqwWo/NEhRRkE5AEdwloBpcqeYd1ndhRPkWOUN5
B7XqrKYyap3b4xD4kFoTtL6WyGEGSQw1TrtwbDiJWIV/M1S6JTsd7l1GApYjos07Pw3Cy5InumDL
Th2lAYtA6ex7fqIRkfrbpGCMWlRoMsux5rD0xsPkkD6L8WgZZ16dWXS7PjeB3yICDa+iMUNDOUmv
zakNxC+CY47W080s++hHoz9oNizElVW8Kw97iByWuxP0L39Aw3pE3LsBbDU3/tENfHEIDR24rd/N
ivFIRK5spwhx56W1ptk+6MIlSnHvm9t2IrnyQ8uC2CVNpPQGwrnEdJQV+ckSJDUI+zlSnufUtEOi
BOAXsG7l+SV9GVr4rq5pADGpfqCZb2FyGf7aY2PJNIgvJ1fOndbJP0PmvGdjPiaMW5AfyF5HuyzX
XhPjRHu4fC/M3qa6wtCYp4/2p37NZhEG14Z3EihUyIxMiS8xpw1WwxhPsghB9Tbhpom8BR95VyPJ
xkLjHGxkwUZsPJxIcDrUZPEs3QzMb0yyQfVN1cY23JxIL3twv7WX9H4tlymKRHTSya2X7w29S0Df
I+UuXFpsA+yHZY9j5cFGS6eTga9HPjb3nlpdw2g2M3uC57gVfZrelQp7VeyBjmLwecnTDw3JWbF2
MLgyfu5z3lp6+AG1bbjIoFhdrSouRep25lrB90V5DZJxvewA71zp0EV2syBw7B3nwn6ZyF/NctBT
i7JWtIFIYQPWKqmw+c+4Jgj1g/PIZbduTc39YleUOUXL750LH0wZSEZH33sk1BBgpFp6/fdsbSTy
AQBcYR04gMRWhT5iVpjQo1xmpW0WU5u18LtTSPC0QzDyRWkKoE0V1wIeAVUYKsxXD/InGYufnI47
TRjTHrrBPAiWqRmQlKSHz8UtNmeHVmYkv10wwTI3KCxdaX4PHlJxVesF5Cwq2d9eF1oPbkruBgsI
dUxsnRmgKL+VVCJNtmN8xLOHoykrOQb4N5ZYnygoXUt7Y19XonKIEDXbmn1uSjiUJ89Oecj+RwH0
s7LWBMylA1EArsaTM+vy5kcpQ1diy481QNFEo+BYV8qI5u+s9ebZLnBz76g+4JN78CEaz978frln
xmYT1JhuOPzYEN/qY/hQx3srcz4XIeYKrFrpjsJOWRZU8VkXbolZXfTPCM2bh3YsTnpf50WUEky0
RP4ih4UNz/KSIy038dCeNdi0W756ljX2hiAr4qs8V1rGz010F+QPDcTosLWoe2X26XbzwBKi/cnq
zHVw7fbt77tZ58FqHCfxgIweqBGejIYDIDHPO2DFKodp1Ls+MiuMJQnXxfzd7QoX4AmIsZ33jaxd
xhOALCtt6khC9wPWuHOWdfSDPbtWQ4ur5Kh+xXDDhEPB9xgp9mjHVRTImWPRmPqAQFhzGNeW7t2+
YxUds5aaLD2zqkJKrz2KM6INAfgi8PkapqppDWDS5OsnOHCv4Wv7zLhVSn9KlHTf5BuvdITuGe0t
eTGPG7FLOparp4hgRMx3v4goemNhfv8wMZdNCZz1/GxUxIKGoCU9tYjizJqke1900sRthGQmq0kZ
Cnhy+sHyN01Q0y5ybTQGxYMxvUzWYNV8JBOMZ9wwF920EV8RgkkIc7eullSoc+f5CTGnjR/VJxFD
uohfPBd0g7ZrzTHfLKjiupCftBypqOsHOgYLXFl6qbAA81x6q3AEenSyN9S36Jfa/6AmgrZU6N2m
gYKxpNlFjYhYNF0pdEC5YE9GwvH7pIoDi6Fe5vbJClNTSEniqO8lxQGe6LcqYLQgGae8+S02RZXc
xl3g/kZBw6RFRO3nWUX9F4HjQxA8n4D9N/2iX8FpPCvugm1s2cSPfPYIB4kFnOyHSRW40G3Ptk61
OnOC7/k7XHI/CIzy0NVo4cOMi9Mz2SbWL7r83U0RoKGihPoVLiRXPu1EGwIHL7Hrnrx8bZY2l/mL
icGntJtGZFRk7Pu32Q5pfIqyWC2aoVu5z2VVIEXbYzcVr25t8Y4619pzXODequNQ5KNPq0QMEUFR
x2DmsH6BDw9ngw1OtFOuna2JODH5c8D8mZC2RuPb+o6BS+WvVpn3TXhekbXS2EbsN2bV5aPf521j
b/7Hw96mrzp8FLTkaWKgq5KPTL/Hp8jmAzdaePwsZGmvT4OCB+dtanuFEX+HuzV2iRfhRmemR8Jp
RCwEZ0kl3CL3pnq5omB9dpeoVaecFgnHahvuS5CW4EoL8HR4P/xF0iBFxtGdel+rSil1JpQ7sCjS
XEjnaUCJL3SPK4yAXt28syRLufT/SDp9YKDLAWVAFNtj1QrZ9njjn8gbee5bCzWCp9x5l3tb7wV1
z1W7WHNwgbCVVulC35PBG+feAy+EwnMTVedtIME7DGhZ2L+2acWwaT2RAbMeJXp5OHGKK0IfptHv
Ylugxfea0TJoUygpQSc8UJAFHkQlx907oFmTC7jzcrGWtq0dpk0CQ8ngwOY7rX3x2YDHNK6VWixZ
RYlD6M0e5MAbdu6N+aKRLyuty597LrKArqgNSn0o8QG4pfU4r6DqRtSmGxEyGxy/LhtxhzH08dn6
c1omYTcW0G7Sat6KcnwnwE0TBNBtslXmE5NLWsOSu41VhQNYc3NUY/aB8mVE58wY4XKuDmVxoPzW
/0x/AVOTJitcIK6GPNW5sxz9Vlv+52sXdWxX7maTeXdYvp45NaOd/Rt6ODjvdAeh+AjcbHA2vThK
nlo1E47uFnrGoCDRX/MCTgW3uRUR8QfAw1GnyM1VkqpxmInuRCdVgl8w47C+EFY2sPU4akSUOr0z
WpBpC/4Bj98J9+pphMrCwnli8jhuLgFSclV+Se2SPRFLM81qdGlbPZtV+BqwZYyTp4ahknUGw9Ae
voZfiR6Mr/ywWGDXsA+sJf2LXxFSnNR4ZKI3ZD/Q8E63mIpNDz9T9lTajp9SzBQdLQjWgFs/6m+f
3xDTiMxZg156Bg0TC0BP2LlpHFjoHyRWrPGsB7JNW3N5gZV3to9YxppzNpaCQMDREi+Fi660Yx68
J5dJTap8uLLUlIfb5jwTQmCXRnde45/eypunQwrBp4jCXEk5AUqNPIhVC+M06fGkeRRw8lKHc7+W
5pOQxu5oXY3ZVRzXQvm88LXzd9NdPJTpWFzzwo4rp3RaUsWOu5dCygGxmQob9yEFLMbGXQ0lCV6G
Uorvqbk7ScgYPpbihUHZR+ybW7o2i11V/t+jyKxoK+wXZtEWnWBBYrs2YCYGJq16JXpZYwBQ3p0F
tIsf0fDgPrnpT37slj0T2rMe8fck0sJ11VglEmMratUWCDs9c1JfkF1qNNu4JHq5biruHz9aCB5d
1jBtUADe+IxygbtFHaAkJ4hGU2zPujyLnVlgfIGDKPjuv0oV8oiLzOOewv7rFNol7urb/aZ9ffJk
GN/xNqwacwo4k1hDJYAL7di2FTcUBgf2XjPfE8QCRweRhoZzL1GF1ss7l29vs61evCvROKzGUB22
a9NUFQ8d5jNKduQFORPZD/OcbZKHCbAv01cqxVCTnz/cpv/5z6B8uzAH9dC0HkcMhD+NUstLIQJ0
RZwa2w1szlTNj00hnnFfTDNzJRNykS3JdO4rs5vdu9LSUryPebfP8iyjH5MMWh2eb8D3EBopQSJg
2gPEfyUxglKFniqirdVSVzf6/y7F9qh1H6dkgkvXKBQ9Rqq3kwHjapGHlzPRRv//9Ba8qT7WDVgS
FzErqx0t5ExQwxLJppYhQF6dY1Yaz4TwMNH+NdUfbI5M3Y9QChVkfuZKsTKjk3llCJKQ20O4MC4W
QjoKdmydAqUGaslcji8LrWyqf/hdx3nvg3SbNiBRZNtpPGBU4PaqJqF6pJOgX1VB8TXaxEuR5dTx
67LtkizaAoD/6yqDZkIuzEFCuES6MTU1sxDLzKow+Qb/Ex9yqXwuUFRH0svT3z7PutRaoJUEPHAx
phBl25XErHEbiPZZ6loYmO1OzR/kSWGlNwnpDQcIPhPiFVSQQs/H/RWp2paOMSD4ImfHBWzfMLm6
kC8DTquEi5/LZXe9Hd1WI/K0gI4tmE1RKYKyqhwDErAdquR1u5Qv6eXdycLNPppRf/KIjnuaxohu
iuGXG8GMoDicti/1FTBbKKtgmcLUdyYESk01c48rTorIjsNg0y6wA8AHmcYuGCMD6c9xfKV5Pp9a
RCFw5oQh1heNQjRXyN61Xnk1kp024zbNgdIJt7Yqfap7jNISkNuhy41yINIwD+6AXtYW0boTsg6s
VP879p4HJgLeO2DWk89M1t03dBHcU3OL0mO40Fywg+hLSRvLfuaqo8TcE4MHaSLOic9iF1XVFsiz
BrAkok+2Tjb30AxSh8oQhXsBn9353/QegTD2WJr2FSs5CdTbM7qas+mrdvBUdruThP4dFk5pm0Yd
ivzYXxMZdknSgt1Qo5FJmqxcGbkEJzhpPbasgi7HI1rMJt0nndv4y0WlVAF7r2iI4Zz1b0ZY1BVP
oF+7nts6kEnwaM3NHZoy/MaZrz9bAyFpfkwh2I0yxLLmm62cteskfHUhdgmiITbm/pW7rY7Fh7bN
l6bhdnN7DVmtaMs/Xl+w5sxSWaKVvlP/+2ZXKS+fvY0ShNPSuUD5AvDM/2WBvPebAmc5If4NoO2S
MvXSgOyzLEHAYRrymznmKF3BDIJ/Sc/u+AcGO5ts2GX85a6aCb3u0VblbrJhFiXiyeWcsu+GCdkX
iVre3hOTfkEAR/+aP+cO3NPIGV73IitICuG7O6Fh6vAsqbfNmxH4lj8TceNP9/oBsQ17stm4pNfJ
/kMZv3JTcQmOuplaYWF7PEMbN9ZkiWXn99yEd67EkSzUkk+i6Zy36rXSNJZukNDAbW4ZPwcDY7L4
0B5l5veBjHasB9VMtNdU6EVOmHFZotXqwdZ8cIvyHUSqsroxB/zhJHRQYuuB+JDCHC5e0tuUh1iD
hCO8eq73cD5vDUdH+VOnEs+Gh6viaAtl+IffuDYcO9ADpIQSOzJFbMpdhEQJbt7tL/6RSsZScfUY
LjPb+9BTtA4h+BCyTX//Er/mP1qyCR0NE26e2dc9yZzVu9FlDWc654pAdPVRN6VBA/6fboOOJ4jv
Dco15Zh7FJ27R5RIXLfYJd0GKcvNogxGhdgoWEQoexdyYSccvoKVrEOEM/LEkdIofqY8Q5ZOPT8K
oOWCbUwy1H2XYX5zX/XW21lDYROgot3BIB2zpuNx77Sz2YXOp+V52G39M5ZRsbj8IQ1JnDk/bbr8
t0I4FBb5n3cd9ES701csMWyFJihBA1dhyEDfAsXH137TswbY7mRVVy0OkuB8I9klP1r8kyEGUfm6
PGP2XgftZgCF8nfEcciEG3Aab5rcs/RnRN0+s01XQtm32Jp7Y4gbTMm/bODScJBUNCJaAAFvoR+L
QyfxtFWMgnmL1zYvGxU80JTiOioxbCLENh2tWBKZOkzPL/B3VqNO8HW8j7TlWZ/RhTlqeTO+70W0
u/LUWX+orWDOUCZxF986gnAsOzCMS+LwSnCTMhG6mADm/3Cu0l58z/O0+TjXg75Oe6+lzN6Ds0NM
G4Smo/xFwrV5aouAqz4yVPibd3D9kCcsxWBhaj1FGe5LkT2nrOGCrZDPOWCWSrcx3H3UHyJBwIek
uas3SeyH4agXEl+qRNKmsoWpwHiKe+IsYnt9sNANJ/wtm6r1De0zzukF3W5+RCRB6LPZd7LbrPmJ
4r1nhDJctMDd7T6u3jIuG6dSM5Gu+zn8CEkrIA6XC67ziz8hh0hTSaopo71bAv1K0oBkpzVQS9Li
wBsn1g0BvoGP/Ey1vY7HI+C3MNlMxAwXtGi1mFkEkF4Yg9wUwrdS62xYh2HT1YFoLkQ1W5UpuE/4
pGbFHnM27rSQI0mCjKyBhxqVMpnu1iMZRAOCt4o26Pl4wDkoSbv6yRTpRwv8obKMtEs5l+m702JY
ihfaaq95luv3BfdByUpZqpHm7wFizgCUfJG39eBZCYGmD4ZjWJ/oqqxmIzp+GydW0YgQbdyyfID4
OB5rmfbYjKB6WAIXdH0B5I84r32Jb3ykRuK5JrAtVl78+uGuXVxvu3E6sP19uC+lc3O3uwuNW4zB
cuo7ArzSNCbGmHVGvusHMRLtqX6obqdnwDY8LXZ8D0y5EFXK0V1AuBnNKHQ3Dk74tr/TLAb5gXWB
4IW308JHOqENHvAn9A/sVJUchnbMtBGcAJ1/4SOU6IFc8Zb0re+jv9pmSJQQmACKlXOUacMCUsVI
MjZUO8CKfcR3mLfRuxprRdOwKrJ65TjdAvxoVQOJAHjfu6BPz3UTqQO/4sMIanvsTdY+16qOblMZ
ncyTWTImsv96tEuGEIxIxvSC6ZIB79f6iecc53O4KnbU8OUCMvfFh2F8SK30BFA0J0xiQqsSe7wy
g+xXk4J5OZ+VL8UdMpI7ZsPI2X+XBkeJCDn8WEC/o/vGAE8jPknwgHEvMp3HK1kHRygN5G7WIzqf
fVwrgsjMq93xwZZcnF60oEj9/kKJwbppX8yRkx3jj3s7XJPkWkN8IlTmWczAfkSjcJ4AYq+Z5aQU
csObaRS7zGSVza3i+YhtEq38MiXI3adLjcItKOxdeFS+VFKNwKpHpOLQIuKws21jDGHCzjplJsbO
az5LufHkznVw1FQnZauLEstmdSNl+wmEZf0Tf/3yv9K9q3Prd1tyf4/su1l45+ZwMIzb4s1QcSaO
t9VkT6HordKYAXDzfl/tWAovvNVgcAMy0vBJmrxgAANSrhuLuaTXykDIX37Vq1+5bhGtfA0zfdLc
UTSc/8HKTGdaZcIE4fEhzm8RfZnzdUopjuBYyOKIqLx/cfYz8PGKk/dbJBXlTqurqh7cQjc/celP
6peRSguCEzdBfFbxKvCUtLvzBR0BXBFQCDdhu47nrRD/zc4um06Do4JUGQjaX6xYbstT0xqqS43C
7TRbxkeU7OK0MP4K52p/s846FqPR5NH0lUoN6oixggqw/BbQRYrPYP3vrJFmVnFJHmaFv59nL358
tPtGDwRUxea3BcUTYL0OEBVlXocBkTyCcGy9qOFekIFnOaXhS5Gmu53q+WZcUR5EkQR9vPEBc2Er
NK+DnVYiduxkV80f8NARGmS75tcNEn71AeDrfFIz1xB1tHppHqEe9Fc2eBUBd69/0tbqIH04pSk0
xDhEAeGXyx3bmVBdIHtSHbc89gYDql0mtrSBJS4ts5a2hv/d3dZaweIxLPf474Pb4mEivtWfkxYE
PsGdythvAdrSOR1CiM/77hcU1a+1fdFHSvD2a64LZyLxsdQXOgHIV9kgZNgdX8bNPMY12Dul1RGB
+mac01+dO3dKMZhLJbDIRfFOs92Al8bgWWPy4sRflXPHotQgIkf7RrDIrDQ2gdQKZl+UQCdtIVFP
SV9cDeZe6KrTX74FWuHKdwR/WRgs1c86jL12nRoj5YxxvHbfbSc/lgrpWXyEorfymx/RJwweLZfd
mUfYrL71+7xg8YZEPInCPxT8E6QFMSA2z6dr24/VGTZr9x7qenIxCLHyBmweEUZ0cLPMFD3Hy/RY
a+8PjNU0U+ntLdR36MbqYjRtOEfLtkcPQevHWq1viJlbKQs412YkrllODkYYXiWaOnVd4tFPkovc
B7lkjXHrB+H4hdPqHjpNx8DN5WTVtRnG1fSHUONEqAwnLTr1A+s2u2A9OH8Q34i0brcDNSnqPwVz
Rx9VxHgsQSe0e9s3JhwaR5d9NMSSSpQwju8HS4Q8PEqp3mhefg9RLvkjT4HyXFHxb+LhzPFE+BTV
uD1cSs7qYYHdpJmxU5Yk8wpQ/02e+kxexbBy76/YIjGhORRUBzyZwyR/ThDNRAdpVUpH5yKT+O/S
1g4/JsOUNn7FnUc6tpjcTpYLu1c7Sse1IhZ0IO0C0el1RfmcFOC/eoOn3wbMIfJZ6qKFOvAAPGVv
nRr6DmtWsbspcWHwPYE2rW07D8yYUhPzCX8QHC+kPQYfQXdHeFPPngYJKLdrF8h0q7UO6CiUG6Iq
vlCCU0bdlJBL9uMI/O/vAM1CEcTLMbONkY1DDoxlBHGKJwUQRhCwrV+viVNBw+kUwp4ReZR57igQ
oaQyG9Azr9VNpo+vR74fQPQqSg3byVBsvrnZeqyMKJQ14hlz/rcba5oKkQJabm3jTnnnak4w4Bfg
lwRXDZzoTZGp20r7tixQ2pV4muSJ+UXbROChc4xGutXGI0y02j8v0UKhkEx9mqiMipeY4SnYJzr1
GzRxpUGn+NUrKQKGRsjecEvO+27Y1rXBfzxwuBlpezF+f6ICrxChG4n7ElfIpa0dgF73gKZJQqnx
uKc4hN9n7ACR39w3JoWuhgpWh0ZwK2muQlxWvTvSrTZ2Vq68Pb++7NlO2Lm8YKQjmQLmo8M1JJo9
zWNnsVgo61dv9Bzdk8Pmmuc+YVGl3uk2yxq5GeqUsVdswrYaaqcMoT8FH5K0PWgIAsrsurfAzZOe
L7IbTIhg8xYOQYjBZtDBxkOrRizdwTNMpzNWiKYh7iudXe39+DgX1CoXGdIgp8iKYkrMvX3cTQ0V
6h8V6t6rbwit/WII8QlX1VnFNHhA8TIZP/q0H/bqNd4/3uhN6mt/VeVjig+A0dzUgDoujBhJtkHh
uqIHQDIxSQG8f1dxf26Tga74k5RKav7dBhbdiBWqrwPii3z8a8H0b2eVOERMBWZDscG5YIo5zV30
kWw1flD4W8A9kYDcG6wEjmjbfLVrEspFuJWmSvh17DsnecTSbjyKH7ouMr6rBQWxG4tfN7FUn2pR
/Jfl/87TO2Y/aLMON+dA7vRj6e6dcEDuHwZHznwevCN8hC+Lwi06ydJrTC1zRoTTacHyIh0yJnyS
TOBc62OQ/l2D209FXPZ3Yt4kTGT5SkSwDDx9bCe4BupsHW4yw5eWqFGla/M3li5c8NBy0PxtnAPS
OWUGHIFtAWGFPE7fJ2AHnm84VRgOQZkojvacpkG/x7USl0tQ8CiNMZ0FxRw7LH8P5qFB2w3/ZJJ7
r7+RZvP/8RKk9HKbUSi7VcraPqrdbfGjJT7Vrr3N6tqy6xze3Itrg0z8XiK/8QwDGnXEjpA7EUu5
ZEz3Ttdti8z5SVJ2FvutptDIzVHuCixvYauNFxGkhw1F9WtsokLEag9SVy884KAtJUoiMC5Zdvkv
FxBCbUIYC4A692qmnGTL4d4nI5+0bR8sk80wB0As5We7kX5dOW6dmh+Ek80U/MXi88qExd/7gY/M
6YDf4oSBLXFuZMmbPjDWWKs6FBJkZBSisalvdoJIy+cKvHOWtQQvc6Qk+m1GnHwse0pWp05jjGTz
9UrvXMXZ8rDTJo/n09zMzAxPkETuxyw8PdseKXEhW8OKD+zorGDvCrTMjX/KawzdPe8YNbytkQkX
8G54dHQKNHbcoqdL8KJGWThibjWZP5pFD8ciAWm8GEqiJptSSpjSgZYVvhHnxX4zTL4BoWK/34ko
YWH4VdOOOa8ETxxti/RJ6zBY/v0FPP66YS7f/p/ytJxZNCpSDYs+Y57ngqu1F4d6fdBrAiFseYHC
3OKKLRMB1yzXsz7aSR3IHWz1MNbey13qJSzUcxUg78YkguRsBdZvGbp+HK29F3ASFN5/xHyJk1Vc
uAwIimuf/kLVpEpSc0O1Wli5W6HN0jAlcSOJlco3ysSuV+FqR3a+vR2c/mHZq2MYZgEf4CcGev97
U/+WcJEb96IAVqKI5TGfyMR1RySht8Tatreqy8kZ1n/dUd7CHl7/AFngTnMsASblOHDdd8IRoBG/
PA4IdHCl1Y114bbpDcOR7PLsz/wQgUUcK0P7lOukktpwdMqrybaTb3H3/vGO6tI78JVEi3Uaeq04
FTRwMV5lYISE1wln9R9Gli4Q+h3nSPb2rZRPYh6b3MR9QcTiUnwYducKqRVHEFTVjh52q8ovp1hQ
1KLYo0H+RK6/MSA/mCUpsYcKGLZHSC/6rfywwDXAAV5O2GEYfYdbw/0ccVM3AsdiAaUPdPv2NvQ9
KH53yLWTgZbRcF+ZSQWI9dZ8xJ/SKdkEC6Esw6Gi5J13pnjfTxSr97lngPZRlwXxou0UKdkCNJqn
NgBCA8f/noG/8nkU03/vGJ6UmWTJak6BQihnSNnz6phpH4JP6WkBnN41BRKMGacEiQ46MvL64P4i
KrKdK5J/sZxxOzXAh+qftZvuO5dvFGb5t1YJYncboiijETFHU7iVGNt+rs1wbmCZjuiS7YbN2vjJ
1Sl7nepJCk8/cfEugdQBi1OC7+97PuPPeo/X+m8cD83yAq+mRmnfD2ABvkUSEKpOydm3gKuvUGmv
9B3LWkKV3YclHbmTKUsp9N2b9AuzmdzSDvRLMIjy65MrrWCEWMsX6lSnEN1FX5bIuo+rFTjExbIk
tFqA3E+KHiGqes4Zg64NCnwZtSgjdePZkzsKrpYd2e33n0ZaVezyJo/OowrQo7I8MdrGVtgOquYA
R1xhDAJ0jyNXjRTGvODdIQgvolNfmxCSOFOwUuYayPwdfDy2W+OE0r1U4O1fintSPn8J5Y8dPCRl
AVZflED1Sg5a+apvrh7EVEK7WKDAwV2098B4LEEAAiMFqdz4jjME/fbwSi6LZvC0gGXoZN/UeT0z
gtBQer1CF9pMfI3APj1zPbCuaRhLJIecX45f9fIoIGmXAm95vmQIOog3EMYzGqgU+C4LqGFEsQJ+
AQXHfhYHsiyyMToD47jd0B41l6FbgA2e+OasHDUyPT1uxQJ0yDoDFRauj0x2tjxIj5IXEEqvMBfB
BNUfI35Pj0u4zoBAr0ymrfLrst/PmUoRFk9UKbe9j7RzuHjlAxDlUZDpSiIVeejN0d596gOKaADs
39HPGgikE7QscMjDK5l3DJT0CcdmfawTmmqKPYCzkGMP9oftwbqf5f7HXapXLu3fdxqbqpfnDskH
1Ksv3H/PiaDCOECM1lX+nzG2/6cYf4PjdFog1WxK2VGKRJkdZSOj5ojrZKoP/diRwheKMluYGMXG
+upLoqMkjY1MD3K/Bd762Tc4gtRwPPKCIOuMcio9ldFHEwnpUzMrfH+ecE3XfhSiO5Jp6GPe5/vv
APZ8dT349uM5lcg27Pdk5nLATRyaZ9ptltOJfH/Sz+PpLGgeUWVwGfxsVpNwoRnazaetpjq3XAYA
QLCO2lWrno3jMat1r02ZgXgTEpTOO2Wg07N2g5gftg59hmsG8B41M0CYuncROQC8DWq3j2OHFhKN
djCowMoqdLxjmty+6PvSRirL7tn1uBuDBw+rmsZF6ChvNdRxUytr+kWaKuQZ7ZBCN774MfV7Geuy
ZOP5HG/b4UpMDaXEoYot4T63GDTv6OmFQqxa53/URrmMckbI7vSK5C+LvfmAWwrw9JrN5XV9tsRg
UV4ONiEoUz8LYcOoPOTfwlxHo0LzHNOuAkAfbLWBnB9MTZ3sqt8pXWlMnZhNsb84xoyK2Szb0Kuq
rJRIQofUh4LPVTVcT7NU+Fd8tT8f8afeUcK6MFjfEEXiBDYjNmp1kJLvo4d7VLk46eFU7s6bBWiZ
VcVGrHvmW9RtMmZJry4/SZUerfzaqU9u9qHcJNeX4Apflf7gOSkVh2zWWPAO8F9BvuUxemhVY0HU
04HP1+SFiOYNhd/ZvR5GnOunkFIzarcpS8cUbscKdvGbke1qBiB/+ocLaMR61rLG7LVOYo31ZIvo
3EXISVcZMiIJCYZNi6Y+RVZdz5rQEv4WPuhMpOat676BJuENVmpbky6ZoyOS6PruHNrwqu2YaLVP
/tz5aKw13fDoJt+/t26sqXxFcGayeJfgHuVl2pG9TIZABknoHys1klX9uUIowuA+Too7JM+9/28B
Ef6G2gIOVxWuRy4beT24dnea30pCjFj2IaJOicw7gsN60te8D4bvcwLn3LXBKB9fpls31BGYlfXF
98boJhxpTqjfswSv+19iYYNbiArCo5v+ce5YYiU/oK2AwjYTbJkaO2FRSJwrKFt8wsLLVFDFqsBy
m8Q3OVbUC+jpIqxuVDeHuZdLGcwrotmeFhh/80Vw4z54rWH8O6ArBBhTfetYIbTXVVJmTutoMKwR
FSt4OvZywaBJ3an5Wv9h8zF6Scdd6KqRhNKedRAYCh5wSsLwSiYljTqne+c2dx83tIUOaD5ghvMr
qQJgclt904sa6T/GWywJwkwAdZH1fW8MRX8UX/CZf6d/eB+0qtNeogtXijRHJ3evNPMHndimb+Rv
R5/JzCnSV2RRXK2o/NKEmjZQlLND2WEZ/lzgF+dWph8M9MHuzCRT+VznoVO3rd0wgVoGOz+65eTk
AsDUrYeo+KIq6K+OguKPbMTPdjF8/b2w+XWdl/8CoEKBdM1+EKLb8LTjtK11+PWtz7W1DZlkaI1z
HSz160FkpYACc/BtjOXUvGI0RM9YgMtxIbvCaQYXQaeC4G43a+VYzR7p/iJeGQVJ1KAEgs6OslF0
zvvgf7cCxm86wGHir8aGXQele8EDXe7aFqWr/AURVoswDJlwM7V6FGwiGUe55VLYxXa3oK6487xt
pm/NIb7Ie0ECgB6iImAtbTcJ95+EdYEP4c5F9q4akRf9FwSXGuKhQ/QD6AJYx6baMkfJQjOKyO6G
mtciyE9SRS1tPF1qzcN4un3SwZQBen9Onmed3e6fN/AtRuDmCr/FR8jQA9x/PTS+voiuBQGoFTor
rInt6VW2SykMYfuu6spVdtTFYOBLkEmES585TqUqtp23DK7k2JzGpzya7x1x+nGMPiUM3yc/Zug8
47Q3JsJwqQHWGOSkyuZDvXPSsH2/RM7h/QnQqmsisiMJDQA/yk1suNkJ618ve9DxWK1/DsrnCe2a
kpU6xaIERVa+NE4lyzPqm6c/f5dKG3HQoV9K0KFrEPe3a6rFAFM7UgBpthzhyroGm48o2Q+HKF9P
hP70Ul61/PsrUsdbENzoaQ5i9BZTjrVx1MNm57PqxOmXP0aiWhTfApjQB2jjRzfJcfXCiXuVUGPJ
Y13ZMjoZftwFdL+fNQedZIsSed0X8ZaSIr7Ku+uJCNZergXBGTC+1Rx21e8OMcV0Bc/whrsMgWbl
BMvvnMKnUXwoITQrLm93iVaeUi1XEh1XAw8/TRIr3lThxdfU7l8bpSzTcyf4M5tPzBB6Mv/38eiR
Hom8gAIBFFj1UlItNfdNUdCsOM/fB1nBdsyfQcSNJ6hb+Fjy/vgcSA3lcdhhYLgrLTSn+nEic4vF
bLTxbkLyviTpAUCZGi6s/ypkTzEBVGzO44T1yeYpKEcKxvlPjYjyOGpqE52vwW/Xn+aQtCaDtMar
kqB2tQUeHE4fwvaJA8iGQwI7iFivjb7iHDGhMca3WMboRvZO7bZ5qNBFmbzXR4X9BSsaNbL1jWRa
uAgMf6UTBmExiqNHRgsaL8w/tYyehq6Pgs20j6Cubt3uR0bfpDGvHB6OnDWa54mU4DL12fpJNexk
+zhnohJYvEqghuoWK3WZLzGOTCS99AyRomxs+j3DRANWiXQdK8l+4YzCrIsUpR07HCcypjYinoaa
ZSRR1FoJ3AQphxwc6tAp4QRGd151IohzwQuVwQ3KrR8Z8oqmKEYfhcEABRhVa6GIBqCeiw5x9OWB
553rLCTdDkLN6KRuVW6gZCWHpsHDmbtq49GQdH2xzpLRoalufHv5q2FKvA/E65iAU33Ck0y3dpTR
+Nu74LzXexE/6ksZoZjiPIzlpos7cRd8H+lBiooLMTndLMVO1FHa92Xrl1fAB3Ukrr9gCkZrjRr5
Nzp/ElZLb4dmLLznBZMMkVEE/SINuzcsqwYoJPuldCCSTiRhoDXVUrQTToydGgwT4+Ffy9vJ6W7R
1w23vZE0nWkYf/ikn0rtjc/u+jVzZIW2c7whZ2Ra4zbqw7/giFGFW+3olLzfoZ04wKYHdbQwtLcQ
LuPjZA7+/gTmzEHz3OpIaacSI0AcIC6ISXY3HggDtiKEi77HkQoanPimx1nz66hlEt4wKD14E1rg
hOwJ4fUt2fKb/YmpckSmHH0KHcDs291t3zBRFklIjcrxqK0ZCMgA2sHwZNxCV4o4n0aci6Hq6hAE
tpTbbo0v+PwFDo5EWISDUbeygw9GG0fwchcI2pnhV89gxCFO4wzOnSb4TpOuiupAAGcwdU8Tb1vP
Vl7qOoZaDHa/+AjUfSCyIitbfrqrYoXSQON+w9iWhXktQFOqqL88GkLP6HZ0DWNFd2egTZhqV7Jt
tTv46opmCSMLL2yDueGcNMMAEPublZB7awJOZOq4/WSmpMvamEQPwiyWXogoy4plQpBZt7OTKIQr
VKwfKkkeXiwLSoBxx7MbUUhG0ECGztZ/kf5dCreN7ZaMWBQk0T8G2lZv27AFZ3drW3ALWPdUVTml
naRKKXMnmnduU/45sr7jSVz6E34F+U3c8UPPAuW+IVuYiIu/Iue1XL5+NiP5kLKoi/79ZN1llnTW
R4ADxMdEUVI1XUsuxQJrf5QuEz29kwcaZWT+q381d5Jiyjvr8mXgCax5XOGFVprwdFZzs5iQbN9g
8Arsy7ukQIOnUWJaCSoMs5m2HJbJlK/L3m6n1dBjB0xGGW1LWYu1fADyDRi4ZahOhhgRFfCO8i2y
Y0k0nRnzQlt83uS0f8TNekFlQ/5X5wkbUEHnOsS3rwfr8+gLl63+B2DDmOZL4c5+fdmgNclP/18U
y2GSIxkdG3dQYCOviDItufSn7BkBJ/qDMTEveWpRZA9b8CWUPocYy8MCM5wa9r563VI1mO+LkMCw
UU/Q/jXS2fu1c5qfndacT7ktFmsPLD+rxb4Hz04FvC9VS7Pk2PEozymrQDI0GMnXoyTKpfIpomRF
wOtVX9/yOu0HpygdPA9ouPCupa9gPUyhGsfEclYTS5LprBKvvW46yS1U8w13t1HHU1uAfjF8cBLH
2byggOcUDwSp7fUJ3JwxdGN8XychSQMpxYLcPqx5aL0iKJnrFC39U6J17B76FjyloFyoOQmwimvg
I0Yg4ke6dUr3FAo6zaDz7VbH1E0BtgusLH99OR1INWmB3CMjPHPwF82Tty7hz9sBjGe0Jih4Pm1Z
8jk+QNVa8OSt+1/NsGr4JCxlG7Bo4lRq5iy0QhHkO6wxo8UiWvOdTjjgCWCJ06dFJkWo2fugfxMP
/HWyVk+/dwcnclXA6AfHp8EqvlGdiwfAZf1EWZoVezls7XVpUSixX4XUJtOvgzbvkk1m65xYx6r1
MNmqU/VhkOKT6pZKlIIDJLTZ/24UxpKTHRAvMzD9ykJTC5LPenGYx/lviOZbJ14cvnwOsa/vmsiK
IL+21G3bsRDDnh/nipGUm58jmqhKGzqemnzs3xCQbFjG8r+9wuvgn2IyoZLr+Fe1+HSVmLLCmN8d
aV4QBDsm0bkaTYMg/JFnboJ0yx7ZIe7de1yMiUP6Qg0YgAt1EGR5toQX14cgbEBQsQTmrnf1kHwb
M6EslrmtI5PD5pyAfhGZIosea0QJ5EvOEWFJx/KyriYVCn0/u/KyxeZpNc2RUsQVaOaa4eXbxMB/
oUEJgfxsrb/FZcIAUAJWKNMrmB1nLIhDPjvrRTyQtG0fMWm9XOJ6AXbdmlOBPO22IX0dsAaWD3UH
jimDM5b1BzR32eIhADM/yCRubgaeIGlLTye8UcNj6XbKlrArYirmXdgZoY3Q3gDRJor0MAins1Zx
3+aD0wYTQe3addrAwqlZcRyWFijDTQM5XFeYSRIz/bt/BhjFME98cZ6pw1qRLg6WRwWryQKMKb4i
dgkcscXZG9oMp0fDdf7WY53kJRuuIMcdBumMiUxhxiYu8vEN58ejXvEaLmOCu7JmyManm3C9g/6+
6O0fDLpO5qqUjoy0aazXZ4fGotdTQ9P/h7RkEyY44KEI2iydjWnD3kAMksBGMMyAHB94+L9bE7FS
nFjWGsR7u86URDguRIWoVTanLu4KqAH21ud3g3DOtIKH/CWJi5ZUCf9FwmmSbK0hLrqZ/9vNjSBn
vU4ph1fpx1YQqMy8H7UxkFFZU32X5Orlj9+/nZ57exboFkxyKhKCfWdVWouoO5btyospcDjGhzqv
BHOwZpq7IcKA3Wge1CJEreXaun8mbOM2prEn9rTn0VNT4umWJcsXIY/A634UTtbsrduaWV4Xb0Gg
kjPbg8ecgtZabFXFtB5Qmw/aTl/RGIOPKzv8bTaWX7wmjZ08E38/7PosiUxUSQQy47j/l2PG88Xu
lBBb0Cq/7mt2Aczd3CDB1uE1BnHjjm5C6SpcF7haDQIKwlaVO5U0M+MPrpmZgi9lXrjvKboIrv1I
SChv7Sa2+23+mSZoKhnbpKfJ3RnhrrUnBCg8KprnAb9PX1Wdc6AlSyUOckGnuxb0BowKecNbbkU7
66zmCPy9Mu4zm2WCL9T+Ud38Bez6y5cVMgitC2M3yuzxM5+jUymVOc1T1heNqlyj14u7+fMlM5cI
+GdmWPXIK+wuUV/8S8jx/X9nGK4eM7n1RWTSd9DGZKGTobESfN11WWGXDhtsHGVTpygdRuYNyB1a
f2WywAZ2FbeSjbFuLtsCQMbQAkMId2L+iEreI/U2vluDsWIYCxWWq5EmRvLRSd/a8MdLBuGgSyYn
EtnmQB4gosD+dqKwA/k7xbmK4+Ur05nv8xhLT/LrmQooQDVy5OZ1EmjcQNRbXQgPrKKArPz5AYjn
E0x1qmnklovy/I8D0sVT9+yY7BmVrJvLZVvRiiSVkZwvpmPRdwPnGHjTuLGJ2BpwARqInrISgpZv
WqOobu1SLdU36TlFFtxHp19o2sdLlTfrr2I6kOqu5b7P6RwT08mrbEzVFHYKbudIDl2fnd9OfitW
mcsk7kA802vhAoRuV7on5xQOhLy4eBDnqwIsPQBO7IYs23nxvetuBuADqV3xrN4CEzW6d7S7l3+e
jPlGyx964TKptptNDgw16wpCCDUfavT0Zdfd/sXsqZ9wG8J4rod0rHyh/HqVzLMg0eJLZE0GyHIY
q+Yc34YpC1oYPKm8uxngu+a8x5Li7FbxNJhjg4bkaoq/hf+BfdvtBK6A7UD2WJ4RHx32YsyPPVGi
ilxD0OdTY/3h+v4cnOQaPgQHnOKvVdmtArZKt6HpGVW9pFAVdMFJp32eSonzz/puAHR6eIjpEpoI
ZPLGp9j16WbfpbKehyJBb8u4KJVVfBGMuB9SlT2EylabKgGxvetpq8aCcZ8eNiG/VM2GR9jzVuVg
Gk9WDGuRh1BK/lEYHBsp2CNyQT/5YdFtgsAGjXKQUMDC+HzUJzhwcMPrNTthmOt0pp2+bDpe61H5
wEqfsfFgEpxGPsgBfULAUxkdGW3xFJZ7R9yWSnEnfxO1jUnVrFovT64Ce7BTzKTZqo6SoILt8GHb
P9Nm4RZ8qu22JKNovjiEJyeUbMqyfLlIXMa22l8Uv4ohse+LLT1bYF2G65/MaEYbpbm24MKT6i2x
o6/zOottKBGAJUUEl/CSnUzJ7RWjy3YaZysRG5n5jUQge6PcAT/wgFpVje8F2S4vjT/+xeM7cOSu
3h51ToAGWJXDCpOLd55Lgeyh1GKiuC3obZbgIQVwzNCpF1wjlG9LtQd5hSDUt1qhqy2QtOPMpGOU
Y7L8OskRKKsL86XMD8cN2XCjMEv8DG0aQQB0d0oNd+f64ZZL/o44wxGX2HJ5GXoyP+UX9/K4woXV
BHRMCBdhI9p6HKPRnSPbm7R2F4YBbyRNSDj8paVLN47YtR12bPV2TkI+uE6pL2ajXsoEVwFizXgc
rl3sz6tTEIKXBVXZ0HhcOGxxnpUDqjWb//gDCrGOq8h+i0O1yOfKAq5RsIV6kLW4eFv1gcTvzOPa
2Y7dUZhF+/OT1+um3Hg8Cw3wkKgPkZgyNHitw4+lKlFs1xejJ/c6EbbDW+lVmBVjU8G0riAgGkIX
1rZlzLCg6GY75F5TE8AfC5O6pDPGzcoS4OsQdNHWK4Rdfz4PmuzCIlsM1ecf3E0h5p3ldLYAJrOF
KNGChbN+9oasg7RNVcPJrwD1UyaRuFcu14hPtICxVabntQkO/bQ4kQECsViYNihS/G7pw6LxT6X1
uVNDgVKuWG/3UrqxA5kgmuyHHS4NYcx4Eo2qs+ZcX1HhiGyw/zv96+8C8hzC8p6Igd3Q5d+s6Rba
vP503c7sDj+dMe8ysY1zvKHmq2BmICd8x2YDXIihcgPAfkYswKD3SdhiJahT+fBiZvWHJUl9oxy6
j5AZMxW+gdFdM1ZBvrf0CGgCSCye8Q0V/HQPu0fdSPhX6O4eSf0chgWbSbubDBX5vvnT6XYLmUdP
wrabBQqBG/v3Jf/u8ofIX7sJ4iOQdLJZnBZc7VH4+rVxw1UEThXTyURCQcSvHZhPWv2ltU17tMlT
aWg6ZlbLF1L39j882rI2kNpjt2yLPaFGj1qCKr77xK92/dUrRUNR588komrkm8ssTqleU1rpwlm5
PE/574jU5RC5ELxeqw6c6kmYEcLJ68ibh+o8QuPaZ/uHH3pwRgEUy3clAEyXZUPMW+ljVmSO9Ywd
2aF5ZKXuoyguu7D6MW4Cx37KweGqbSlmOOkxtM30hHuH5nA2feKFZdznZpKb8145mMfp3HE2wa1C
4HrxMOCfhyI8h11U2iSFOuoJEGyDdxSPQDU0ieLTbBtEw8A/7d1xrNUDkxxQNTpMTE1m43oxOE0w
0DOZITQI1HLx5HsV5mWTyNpEecHVoStNBkmC3/XGjAjD2trxBG6Q2GWfQCErbO/fvn6sTXXGZkL8
WPeg7Ngh4TwY6KyW4OzfELG78rsd0TlobUOSjuAh9xD3xEl0pv0oUx5Kw7sDrRR6AzCOKFXjxFFo
QHFWOx2s6pBBlOVeIBKsX6NJ/BZbAMNmvbxLq/WuhAst1MzFIaUb41uI/MfFrB6dwnt5FxWe/YEu
F4vFLg5Dww5th0TNvOdXCv/2indYSGoZsrKwRUoVmXwLIN7lSafQcslv2oHj6UeJyPHMyITr9pF2
d/nINcx5gPKpQ/iQc2S6+v+FTaEm0lX3JWplmxcLTsSdKmlHXB9rsONKZp0BP31muvzjm+pl72cP
WOp78kbq4BbxOmeJYSWIRZ5LNE6/MZSlM2VY5m9v4aPyxhmZJZ46mu87We3d2qugRGz+EpWkCGk9
t0dkVun9+821vsAfRgUce0xVV21zuV6gQ/vRRRuYUBIEeAXVK7sd8FDYrgCgYdcPiaI3WR8JR4bf
h0/fWhV8hrJ47RFB/r4NbErcyvqbJx3ymPY8m85TPt/fQuvLFhJ4Nms8gX21FK3ThyUP8glOmmHt
Zb18pjWMiJbJ5mAgp3CUsZUvzGWUs3y+Z6NoY895/0TxPHQYKUg1AyY0oSbDk1wbDIDIo79eX7TP
we5s8fkWMvFSMk3KfpEvHBnGZGhxcOVHFJeY93YiAHdytNy9ns49Iq+jN5Q8BN4FmLdeehM153eZ
tNZnG1wuUPSQxXtg5lY7CZSvsAbZhnwh5l2JIScl1r3Z9fknFVT1VNIE3u86hCgJntVGQmwxgyBl
H0y4QNPR10DJUGbURk4iSVNXMum8fM+v1lwYaKXvYpPJWA74snEpeVpdwa5Igr+xmcS5UmD92lRo
U7XjRunHwOxbEFOTEtvgKjfPdzHkfqs7X+kx7mtNXzgZAzMecpuPFCflkVjh920hc7dvD6epAV8I
JUFmTtcW1S51AgBKdata2dDbT3MW41sUt3OvhJ5CZdWyuh/A/VNCrbxwVn9u0hYunWo6BmFinjBG
md+bMMSPnvj+BaAbjrtMjHL7T22W4C4vlmTtadz1aTpV19djXS0fB+IzOBmKCP5wa5w/9HNX+rUg
pIqtszEoK8R/CE7kjyj5j3Nzz8PaS3hZYr7n2qDnKeX3xrGvItfRcnQsXJWhM+BSC94SIgFjU8hj
4RCVGpy6rNJGJtSCR7JL39C3qyEpbEH0fxbADMIZxD9YnKyRFmfTMiuNDtSnaJu37VvYBGbG/8/C
wBuv1dKy+GuNzo05345H7QNvZHYuh8LCQh2DTgJBR0cAHZ8PYZ3NRf7NG/UBfM3HRRGa4Ov5bkav
Bh0ddZPjV4mC9y5ekS+k6VvJ3ZgVfgFKV78tXIZW3DiMqUbWmnJaCuLVysyDVNTKSWt6aZmyaCE8
1134MTHckt9ZhNzdxTRK6rOhlVVvqe7GUGVE65CRJzA1OUqflU4IDo3y5GUV7ThIXQE14jlCDBEQ
b/Xgk+W3ATdgSrBCyvHv0Ht+wVr6Y9h8juXnUyxOjN2fJgUIQ/82nnCDnvgAwTcvmtUnmROpzquk
ULzNZYA0nNvpZ7RikdZzQH2a0XFaArozvPrzsL8zEJRZGq9ia1SA4dPbUbdYSHxsRVLLku7jF3Ez
fyrn1hO5mE+CWbzsOiUq63OKs68V/5AGOX3LwdaBQUbj9NepShjn2mNjx1shSTgdtDxgV/s8cJAq
8vnAmSdpzcJGRoV5+TlNozxnnhhMWsTcCGNmejw2nS8k0Rg4qd7BgxXezvb4tDKE2kqgpdbwEcks
RG+FqMchLioFOWQYbfPxa4WEAq8RhJdGsriTY/2F4yrDkzB83WwioWCGI6WwFZTgwqVZ+Xc6hkp3
Zpkcv0P0ryD9dsbgT3IT97vNjBrMebPACOSyt2geA0prZs9pZ+wN55XWxfm90LdAGa/LGByc3Pb7
C/ms8uQELO4fMBmtA13aQ6r/O6KhWcp7acsziOtrOFoJipBbucYSOeH74Pz535Q530r6Xe2m9pC5
R0ahe4ISVDjLOTeEs1BTnyQ73Y9MHrjjK8GJIRSZZIenU3p5lNoPY+AWSKELCjqlX26urnG9I+OH
ozRVpPIaINOImE7m4imR1a6j+rjbgEJHQmMovFmK9nUbsW/EG+DLu04OpIZsdm4zb1ci5l8en475
iGfDNP1D8DCyxLKNLL6Uq49DVJqe7vJSvjNe5SjECxK4j/OmBM9RmRsvOxR7/xYRifHfPN2tUT3k
lCthGr8ag1Kz7mEf1eX/du7Fgsh+aFzoagSjFjFeen1t5FF7cbNPByqj/jrPcIvrrS5L68lY7O6z
BNFlgdsPNy3C1Z3kF1K2G+ikqMqSr/C1SoDHk+FGYX7GQKgAU6s5jA3SSM7XMROYU4EPOtcodsbr
iohIOGCqpXfUR8skmFzD1i53wNexwwH4yo9p+PlFrt0pzEtVmVYO3HuG3plJR4zLyXTUjsPWY4js
o8uZbYi92OycF7HEYQedjyQeFmUbPA3zi8tzzHPaXtFruWR0aI7icEwPtwiCGFeifxq0jfaQ3s3e
SVl4qrom0GcmuPm6nBzh8pougNuLGjVTGTYQjnGPBDS+98Yv9hJ7mzrTUp6mCWTj3jKmR1r37Mss
eeOAeIMSa2p8/v/i5ZVISAGt64awTm5JZjzkuCQi4fDP1vgMeyIY/IFChrf3UxQp7iptw0dG9B8o
We5QJhgUQ94lIPPMrdTl03rk0olbfTyOJg7TFsdGWQm/MVNmuJ/8b+9FQpKFXw7HikXwdYXs2qmr
iuKzJJoT2Y8an7KhVwKrgo8+caqIMXlf8dO0zBgO8Ps/WNVVunwAEq7fqPTsng5tUnw7u4Q0vgYp
hjOIZaXcNegxcPIcDquJ8suW4h2pYypHqT5GDC+wjtYpWzxbE45xyUIPRu7zTAbfE+kGbnVDaN6f
7xgzLdakqZShzHi2wwweVJv2B75KEEC+XX7Rg2x0s3yHVSFYqRB/3NuiC4Q2ph9sLXs4AA7OF0Hu
OKz6YS/NtPgo9PPwhble8wqexeQs6sdlgP2Y3IOqQc6JOx1TzlspmsMejXvDWV/ZvPeOM/CnD0aN
CVwohFjV6+ZfcSzLuTEGMX6Oh+ZqOKYb5vngw0FvS3CRHARJk9lIXgdVoiDqfO6BB6tiYJeAytx9
HqEot3lLl7E+bDB7DvEs4OEAmZbUviGKHNwGXCqgmIKKXhEveU0vrk7BDIduwGKno7w0H00Vt6pN
LXdVO2Ijod9689UDJvdGTKtqa4LTsb6OezGyJ2wDqGV2S4PddMStxE6BkUXTErak6r9r27d55JM+
qI38tXOiqejwYvbWDGuxvq0raETNjMjXjUtrmXJPbaJ+IazxiS2N7bmxE1Xqc2Hck0kHDD7oEWQp
bNF0FvEtgG1WTn5a0BCnfrZjPTORa8bE+tqf3S2Vv33NfhsWmChZu8EyN3W6EbxMpstmhn1sWlw9
OA7vQyOqs7f6uGU2dKVvLg6UGyRPfwAgOW3YvDZsMYcx5tsjqhE1g27pnX5JrMujTIcmbUsMBbT+
b6F8gTtHIHJXazwFZNgBdnQXiJ+7eK3+jXn78pJGtKXfXKHcltz+lR1xQ/7o2hFGf71FQ6IGpO+K
Ry0kPXRg+cmziAkiBOW2kraGD4FwzIXnA7D7AMwzhts/dCzbOpzx/xKidUqc9V5jTsEk/J+hipQY
hGDeX5dppFd4bTCt01KlEd+6Vs8MzjJKi3RESOXvNN6P2Dw6fhXhb2edD29f8Dq7Cdx8En2RRIn9
y/lbMaxhXOIMnIL5QL9TcU4iEZYhthhRxvr2AU8VoBUnLyUg2J3HnSolhJlyL921jz6Lt2Q4DMnm
Y9wvNRwnHGn2auUPWA++6o4AVeggHFL6xci576wjeHvpcJXP8fuqN30xIbnvQHyPeDDOdHgH4yFW
o7LcXeoPlPBBuiV/fxODyvEw6W1PLeqks9wToS3rqvM/S7mtnFkuzLGaf8h3tXK6yt4mMEtOCjV4
c/FBH+X2zwxufmqqiR6mI7qMrGkKe5AfsA9mujSl8vjg0YJVnE9z1CvTLOr4iM57FE4yBSCa2pBM
W2z/rk6Z4a/5Gdd4vXP3qoQPqEYUXTv9S2nGL8m2qjxFJrBJy53Vl6X5PO3CIpN2aJzB/Za2Un1F
9CMAI9pJSXU7SKMaFJ0U+OOHkCzRpBEZ80qucaxW/dtDuxutNHZUhrOOgbX3e6tEQt3Jb3m6FL+5
VZWFF8M2RyUz+P6CiIDYstonI9l0Qd1MqmaO9EOrahb2sJH0P+CD4MwpqSDI1nyy6m9ImZri12Bi
XtzvSCH+Xt0cCQ3x4pDRjillJbsq4W5ZzCzlgT2uuJURnU/sl/6oKDW9vVc1BbmVVAKO1deF0X7S
labnwgU1naJaeoiMGL7mkpYDuIplBHOTeNOCd/m6VLEbL6CjXX/w3xk1p0NHm9SvOa/LU11tvo+O
T0OOaiNu3exbCEPXMR/kkrVf6WU2yDfE9/NchRg1vceJV/FP2Ts0jNImbch2acLFbyh4lk99EPeF
vQ4S/oPodJHW82PKCmg1u+QiUq6W4TNLfuHKgi9F4KGjU6a2PupAhVCnZKKeWMWy67ifUVGzwAxk
qHuDVEKs1tKzmFLkvo44D9+tS4Px86RpigvuGcVa9pVhYzEat8I32M1dYdLJJ6n85tozd++0AWFm
LaRaf5xk8tNahrAzOw0NhtbmN55lfTsu97dCzH6WyRdiPxg6a4HN46zBK0GxRk0Vpe0eeYxDRPdE
GZ+fkSr6F6T8i20mZ2BT+V4WKuV5eTAlpaweaa5134z3Nw/3snTbHs0YkCvbWMzSdXFRr5uP4jni
13UAuICoe9BPBh/KdI4VJeAf3loUSSm+OPIcAGjkZjdZnx/LKuW8ghOKiajdC8a4ExYrm29aN5n4
Hn9QOGwkAORR5gJ1HxQqIdEHEmlHtL/fYGNzqSPA2/wBcDDNVLDamh642r+63WFoLSBYiVMZ9Cn/
1sriQYfTVYGHNuUqxHZkiIs4tfT2Q9DMflDgoq515jXQ1/IOzIaiRWWirjpCYClfsXI1Vt8MzZUp
z2DSkZVOqTs08j8XLKOo4MK8tZTPLXmnRLvP49GcPntAg4yrhO9OBjMxQYbHD+6du8oHZnsWP1qP
CarDaYQ0S6mrOamSitGrUnYASgOTRnGaWggUcUSwo9lkWnw7g+W+CkaeIYc5jBaULGO69reQAN9T
8fQ/UwlnJkN/Y+FTrzPisIswlF+8RKKnn60auz6hm+2yFge+nC4I6bFaXjbpJE0K7yg18+MOfU8a
s4FDt+/qNE/iH1x3f304pNdQJC1een81RBOopcyWeFPjSh+zy6NXweZA21MgFf2Mf2sXWRnzG8Ux
YBaTIbuA8gmFiELCMs/GjrcARfnDSwMdx+xfYUMul6f1fefQk7ihaXVeenlZiyik9RScRSR4C3QV
uT8r0sIWPlBszNHd4/2lwEDPx8AW4jF8LdcbH1+0ZQxmX4kGP6JA6I27Anrom2Ws4Lf4rSpQ0yWm
nVZ/+SxbpP5GeESHyZDgq06BLtDKQCUtVm8qR80ITM1K9P3Ptm0obV3eCpvOUqnP4H+0Zc1dye71
mb+D2unTPBInlP/6VD6EMfSQaZIaw2/cqR0A1N6yX36yOY/jiDf7woh5ASbd0nCC1WSaL0AJy5rY
rSrl6Zljwh0ca4KBmEo9XS8JhVGBfRGIufC15JhAGTK/d+DDyd95QM5hOMIIGk9sotYWoBZz2PW6
4AwBJZ4DBHVK6Wi0sFSj8MgMNMmh3fB9tZDGKm4M/N2RntTRY8yKMDYKRzV2RSm77zIPyfxWi90S
GDyows8NyC42ydizZbRJ7LxX+e4ugRpqnFb08xgi/8qn2/XGwfU+gOWWdpgYpxVBDMYKvHl5hBce
1fgdhYFC+/CED2svQVOafQVyXFc7SFP6Z0XqnMWlaP/E8obUS58KrZXRUb+3a0AQZW8qqRvchMip
5IDMCfb9eXGPSP3uzbC3tMk/7V0XhVV76ZV3cnLcn/VkNf2jEV0xpEYuUuB37b9NXf8NcpDM0XH7
Znl/VUObqPXP7aQ7RyG3Gz9SvSmI6ry7XdG/3m2+TIgeqOLwmR8naUtda6EfamwX/Z4Nc3RKbW7K
TLWKBTYslcr0uE3SZb6A4NiaNXFZsgN8FLC0O8n9C2Q2WMMHaOLDwlQ1KfGec2uvauhkw48jggYO
I2f9GCRPob50U7SX+6lT7Z4JKhh+tlz4KaLCvio09wq7DAE2PSVK0XJywlcvdJkR+gOWdQN/6IGD
NlbHTY7m9jvSHw9LXgks93jWnjyev44VsjwTfa45lsSp6ph3B5TmeaQ5FSI6U3CgWgo5SovcuFSo
Fui1lgAW7TlcUuuG8yZt/s92hIdw0E4N/X53qQ6tuFxfIsLPMNhKmoe6oPH7HUs8apkObJTdWBz1
dw+kxgm07NfffnLoM+woH68tFUSgJyB4cIm4w84FWmZAamsXNALGBmlj8vCG0adZzeE1R4O4rkFa
hD4B87dixAKlUGPRN7avNxpx7MiIFvPNaUriOu1ZbWzjyEPPSL/PAOCsoEQK5M2TdDoih/jMofB3
Q5j1D8tk6Qjerfm+UpEgxUN8RhPqi81aRaU6Dfmm0nH0QhJ92B0NUT5aJExXdVFp2a4rgdmUzKkc
XxBVAhrLkgQYnUrdhLCdCT80EHdnJtnOGbGADESQjUCf7ktdaal6K3KjnP8PK/TYMJQoAt/kId4/
wuOur6i5XCzbLvelVypZOMRT0FbwLE5xtuC84LS5X+3T289Oa54D6TQBWVzRC1HZfBq3A3CPkpte
iIhEgHb1IoA646dorKwAT520Lk977Qhlr1AuucxD/r64eMz+KvszMUmbOeD3V/lrA9arLufjOdDP
TZKP3tgVJtJ9I6t6zz27t/bG4GhfPqELrewwZg7vjClHOcftMACpB8JfC0DQoS1gyooUztXW79YI
wuxPSpHhLBJkjrB3dC7hYg8zTHbt0ads6/b7VjcFnDxgnhJxCleHInChgf/nzZGAIb3Mp/0MZEGL
O6SZ6M6VJylLbqS/WSnfq5t9VXmqilE8o5yMZdSM9YPdCsuTLRkW4EBxocCIDsEYq+kik0Mxta5j
sFOr19mG5XlfFp8p/p3dwOG1/O0O5t6MraOfAMLW1WKLAOV+VOxRJ55+dBm3nUrV/D7dbM1p4vLY
wYAkcVa4OqKodcgOPADuH+U6Mcoa4BxC/ftaOEEZ5JBtWMWLo4BTzWK+cRK2b1qUGfwiXtHedD5a
o7xqrIr4J617bKxILaNCCw8VS9XsWBj2mJYzNzrkTkbIqjrtujcUvKxYggR4diNNyS+gbSmXX5Yy
gnRAB2GTpdwde2bOrZKrrg2UIT+wkMzXa8IcAK28pUYLTHSPjTRHvIYUS0f/LIG0gsxKrOkfsazP
FXVtUaEYiTEOKaF31PPdWKN3KArB/4cqCleMV3Od+0LY/D83CcDpl4qGnTp4moC2jJelMRGdnPq0
MNM4k5LI+4pKZFEB6E0TYyfS2/ogLK+Eqx+B5JXb1rBTe7Ry5ZyDXmk9PwsL648Lnby3WeH9LLF5
KHNndRZnLmbumk2HX1FfBnz4Yawx0jO7/eNYy2+hhf9I9+ViEGfQQpSBX61hWQgflOl63fmt1CL7
RYTjgpADkj0UY8ZVxHoGViidH1m6Lq3ZexCYZYemJOH3v00OVCWLuZ/pCcx9ydyYAlv3NMfks03y
+/weueKH9/OGZzPj7BXXxW7EHAuBE/hv6CXOtoz49869dgNvZbvgAmMw0zf9pLI7XIunNt82eb+T
R8zu2gmNT1qL7PqFWRlcZiYMc13V/jITwpNntYwiMsx7Ppf/Kly1i76zSt6ZbANpSd5ZYu6wymc3
v1jwhkXP9hRa/fI1DEdBbgd5cLFMEoxLbkBtlP1DgIX2LJIlObNJfDMS//JBGpOHDGXSb0t9oMYS
izICRTjpkdRjmBIhpWw6X/oOFE/dd/zJPZL8ua7xmUJRtiS+miRH42cvspMNyHsszNQGIL2TQn7w
1WXAtSjuyCK0vbOP/MpW586JA+4QjRx+rwVIz5K0rRILjK+G8pZ4S5ZtzExweZP9MWbyBusGnITB
bMqDGYiPC8vLNHPTME3nBneoQCP/31XSnttgLrdtpc6mb5vUXyP8mcfRGxZ1AkMWatiVL5IvqaNh
OJgTeapwdvHe4bpt+HNOLMdCZcnfS/45JPsxV6z8NsiFe9J2OJx4X8Zt8PQ2F9C6bLiB42F8uy8F
qQSUB4JGhv9Q2IbpyTDIuOCqApOlghFi6M1oL79XJ7P/YyskAQY8tz4PhzzcVg+RP2tQterIDoPD
TFj/cvCtH+jCdhM1YoZkj1T/X8oxKsbwQ5FiJRSQ1Wmpj7idStYDyi0cwDBnavfDToMpVgqAq8gC
RQ8grI2elrP5fmYtM0DKbZITMCpvtM/d2xQRy6SC6GySEr9XO1OIDAG/hXQXGkHAaBicdsgTOA6L
UthhHRsmeXdeWXRJMjfSjM6OIlrZEWVScWo90igLlKRWHMZq+CswWw8Y2v0YRwRMrahKd0okKqWV
P0G3QN0PnOyFkLCZjXQO+gJzc3ZSL8aydFkhHYCKFacbCeXaHJn5Ex4dr38p9WUzIcMXnJqFtNVO
rSKXPOUrVfddlsBDqloyah39XvlHpsBreMSVMuSIx8L7qLvjwhVadztnvyddY6/AOF462UxHd9+4
VIYEWwAp/SKFRYKPZsaBJ5uBTjN9jnFtm/tRX7Fz6Y/TJfmkaXpFt9qqTzBDj7KcJ4TsVU0CQUY+
T6UaSQLJFQ20D4LOdXw8+1X74V3EOW6JdqMyl1xh6CZx3EC7WVZeK04E+YQnOqnRnTrSlt7+HjYQ
iz1dcJXSEwHAsNh0s8jEyOajSk/aUnKgj5yUtzGSYk7VK+rnnGyhV/Neb4yp0jDktZE9ht0rcFWW
24p03IOyZ++3HZh5TO9dlwMDw2aAUcZ3lknMXPn4YWOEBkufgdyg0Rt4T2A+jMMFKIPl3jcbs6T5
f46rE2/10iLCYuu8+qN4vOMM93Ewf5et2cqUAx8U7YX85SgwA2o0luzpN5lDeKXmg0cJksoQDiFv
CxswhbFvlL2oRq0x2hukMCH2OGzBXXs8AqTLUKZIHG1LbnfkZXET9lvkcg4sulnonUE07kX7GEQv
7ozXGPY+e4Eew0IJ3aJa4zpC3+28PWND+GpAA8gl8/Tk7EwpmHCIJyebaHOVbl21l50FgBDiYorZ
tgwf5s+YMdaBV+U9VPhd6CnXpxbCFovUmhUGxh8NXFtusDX/1Xgo6w6SWL0dpSyW0dEDKmmhFbNg
HPB1Kom24HfCfyE98wQeX07ENZvxIdorXRrtUgeXpLAy2TJ5mqYPEtARMCWbAyVpDQoYpHPKklc5
aX5NQQxdldXGCXQ/6tBXW1mmPu0bIqMhMPWOtw7YnzEo5TybNLNJ0I0BcI95+1MHgubYlB6fGvPp
hU6CKO+aNyRVZnN7nJ+3V88IHT3uYur0TDnTZBSZ6vJD1aPZ5B+CGF22rnsB6M+2WPBigsyRuL1F
vQnP078+dM8UihlnZwHe7UGnMuYUV+xH1QlSf09DUTwe093DrnEb+pCmhpftJbGHAF6+Ouh49HqG
c6nDFQKQl2fwf2hEW+Qepl8RP1m6mgm1Pkzw+tPhDnqh9VN2cDG+sxkvhAgQTK6Zcb5J/udnSQGX
W4tzFtVufRj0M4QLK2xxijsmwcgcruStHnIDZpZL0ksiGZymb8TtD0l3QrlDG9HJtDa7tK0lz6Sw
iql+jjQ457mISgZ8IfHK7AjjhaqCuN0gYXYK2ZrW+5kMn/fYOIdHMPoXGGApBkgny7uH5nkw14ix
UHRo2FsWmBeHBmq9ZHpMg5/6nCVfg2art1SDR4Dz0zrNXnQ3gTbVybtQLdSMqIwxECit3lmrYPQe
LSTjBviI/e+FrpTKBfvsA8UaR9zMtr8niEcvdepJV8iZQFZbtizlgtM1BcgCJEXB3snIcGpzunjA
N4LuM91A2Iv4VpL7MrZEo07hqRmVXa4oCF4ehfNOp2hSU4lYeAPa4wVlNXuZQlrFkus3UjA31PFu
TLTyH5t/9DDBlsQvbAb1UwD0QvPPW+4LC/tKqLjdImgut7imifHSV4Wc6G1s6AhWRm4drNfuJb2p
r42dKQtzV8gJ6LMjJUCxrB+bvKbEgmOhHrEVOK5B7j73G66UL6Te9A5E/RKyTguUNd/IALjJOV2P
3QpiTjGQhnOYgGyGtcHWZDlsBrH+MJ7fgg/WMspFEaRnksJHuAnRei9gaMw8n0pVWaIf6vM/dxuc
/Hs+0MPc5ofWIHx/MGqmkfsPE0BIBvVPRHziCxeeGE0TCbH8klFT1onSlxygRE6GYYKvS5ONsWbe
BLORIQ+2v7K32DoSZIc8ilF6cTcLHrYWQ29Mimes6jV9RZkiUFE0KTjpaZgMUZM1GIT+da9nqyIT
pQgQqkHoo4tFWaD7TLOGQdiZ6PcWd8+Jh667uVWfZLw09gdzQviW6cZkc7uvS/VPL4pJtpwuxe2W
c8MIALGV5KuNyAu41j8QUF1w+vs2Q1CozUL5OXP7ffd9OEXwg3//rUpK9kBplig4o6djgzYUAWS7
psgsfMVsOWcG5x2hKDcFe6jxM0jQ4B7wOYiMpDi51xQ+Ok7P1aHHSytlgoyCwyHEZbi+uAYxad1k
vYBRfVWKIepe+EwL3/pE3bEERmqcdwn70GAGFHVwqJP/0VeUtGhw21Mk+K7sA4hMVlcmWkYNXEYQ
NpodOD1aZ8ZFGdAV35v+Trui3N5Yzp5NlKxGCinROHqJ237za2nynIElhe5491NnDCuPU4JpZEs6
ODZKFbDh233baMJburwrj8mxqZFyaeOVkhafTwT+f7YDhFoha3pyjpc/WmDOtnS9BE08UrAJtIfN
bVFXpjtf0y2PfrF97Z3nRSncqg0pTr4Bm+0Ab8L+MRCBOCpLu5Vn4MH0jrOFRcHSYGynWwDeHEno
9p8tDyttzKVvTOf4WU3K4/b/1sx/UuY34wNWNjSX1fngbkqvcPFbjvIBAsvtMUXFu7aIdxW1uGfA
b6zGxK4ie7qn7t6lGblSkZd+KtLhMLdGi3gqloQYqkojv2rFoiN6Pp326XUsoiYeia61+RpOclPY
r7BsOlvHWuJfgYD+vKaHJV6/lbZptABUysRxvMKg7uq6UVjfVfy2yhZ0YcjdVnj8ajT31NZSNuTk
mgbRpi+Toz0mNiCZVGLTWBqES3jL1DklhSLmobW+wEh3Ub0AoG1Zh94v4JRaDnrl5BpNq4+ThSME
TijN3i6PQuHP90vOsECqc6NUG7qzsA1jwfvHkx5O66ymSfKBoJdvLg4/HD0olVS/1F2r+Vc59zF5
b8y0Pvrmqm1fLlMC36+Nvz9z1OaUiki9pzWEBkgyELqLEpU3JwSy4EKnUJ4wt42UFqzaANonDDUc
Lh9fbfTagGZdtfkPRwTPNujQ59BGUszvsgA4wzIs3X7JDPn0yVCEx21XnurcS5u7DaKCilnLrc0l
N0T7WqgsJwnawm/j4T5TlpT4G7EUMUv2Ke/WhN1ZrZ5qSf0LSDlOwhQjwvGJVfYfyGQcmCweYuUN
CBgkfyjaqsxaOJR6WeGp3zw6K/zTfslKUTb64CfAgMfq/tsfBI/1Od9FmtmFzG5+FX7TnICG4erG
hqEM4GXeGGz4k1nmpWqjXpn+le3+w32+gUZ4kW5dun2ONFWkCU03U5zV+K5O26l49lKKFWpZxaTq
rdbXi5Y4v5t0SsXWeEZ/2K88rZQZphE8+Nwns7tUwptUZ6tUPJ67BbKIcoW6fNAm9/b7Utx29Vzq
wevVhHKOh9+tCVerfX1kEH0Rna53sBxCV22rEh28DUzt7fBzRysbher2ynlWhWeWizKz5HyDXmM4
sumVrpbqwbuzmIBah0wjk4LphJ80KOYcgSpNDJQGTu057SdFYtefg8baPzwnMWdMqAHXMK2Rf1/J
3i72R3QAA0z8GpgdPf2qSgv4JP3Dz2puYqoEN/jfn1Fthr5zFbfQAOB+ymy7mVvCJrWpOoqSPRCg
yUocFLqACs/zmDkV8/ZjN4iFClPN+6T7C9n8wSWybkMDp01S+6WhSMk+egHODGppsHk652JWSuDE
V9OdAdp4WcXda/E9v2aYt9rRlNyRkxWwQ+nfeWORDiGBUUzipWYULcEGfVAxkAjMzH3c5eufcB6s
Hpa7Nui0tgTGHBKLexXQiz5XTBd/J738TKAqax+WAUTb+c3SLTyH6osav0/Sbp24DC1gyXUNkg5A
aR9X5+jxrRZe63OyABGn8C8hnO7eax5RiMiEuk1TivcPvRjqY+KmIWDzamQ4u9DV+tvz1ETNSfMu
DFeLNIkQ8+uVRWnmaV+q27LXBfsJ+lkbFgHL4pN1ygJOefgaxsFMOBXyfu/6XdZfQnZqDF1rej3d
7nK34ZWkc0QX1CqhWXWUizddnaZQYwzcCesjyZbArH5IkcQmUZNjxo/RKgB9U4jd0qRMKueJBREy
OiwEsB8n7APe3mvcV8V+8p+Rt8dIQ9WuoYcHw4eGC+CCi6BUPKOw0lnVWc6iyBYztUSp1M+dCdV6
LlwqLsH+Cui7bPaYzbsJZm2XzfmDFZO/UguUTrcB6JP6k79k2kVvhXaIcOZAlS4vad5jBNAnSMgl
TeznQiunRYtlato5KmagRumFh/Xstdx8A4HZL6m9zfhFuR/zPCl1xphrixWadXaMVkcReekdmpJU
AeVD+8QlbzGA8PmRRovKj9dL9TZRSGQJrVfJFEO85jO9jqetxKEO8yVUqz37f5a4XRYIAFC2zb11
bCJT0AIz2Lzp3bQUj1+01ujxMdEMlBkAjh57ur8UPIFES3mNOGpILq0o5vI7aX0ixY38fT9DN1bM
6mJpFTPKaKFVQ+auYsenArSm88q79dO+RMF1VCuASI2WoWlAdlAHy2RHXSYxEmuTcuEX6/mGgECe
I2BTM+1ha+Y9PzjzJP4iT2nFfwQaU6VkxyjPsAXLWkE6MbbNZ2V43+Vpo46eOK+pOiIQlfsUWzep
JNxOpA9QHytn6nNl9izoOnFTswtHZwD4izFUdqlj3WBJ79+ope+bT5Z9MTwzAczfZd9gP77alQVJ
7vEaCp45w2X3vUnsbC8MJxh7qdeIoF3mk6D2KXUABOlqpMhPidWkiD1Fv+NvKdpepZHygbaknXAJ
uK6/Z1rSdHb10gXkQ5R27xnzGzjS+l1E/HwOZDf9xwFMoZ3+dKovlF339eNM6GhoVd0EKhJl5xe5
/MwcASK+z+cMVQE4PL4hCnAJOk6IVnMdTnYmoz9rXNR94IT6/SX6EdzTgdUoOUf59ez641GKYNzh
sYX1F5ad39s2hVURfXeRlg/l2sEYJWEqfGrPxqyR71A3vppPQ0DMcVB9HGPzlJgVm54XBhNGKabe
jAByK5ngH6H/rIYG5FQkGTTpIP4+W+UMO+fVwVfJ874vRM5wXXiVYezH+c6PI6XKplGuXp8sLOQn
m+hZ+N/6tg95K75ewt/i7YdPzDbNgWoUqj3drNpP8QYCewHED8Q7MKW6H879TH5MWC06o7rmOXWA
OptNnebZvlZnnZJM0lZVeYQFIlwSXSMOPoOw0efhViszL7vtV30LA3VhGOuj01sTKKm7rrTghdGh
GJMF3LeOe3Syr1qiY3P7MGio4zw2LhW3Gq72MpJdg1Tefw9CmwgCc/DBYh9PukqIh46OIyTuiJHk
2bVh1CNbFoQlhjVr9v3k495XCXcPplgphRVkvXp+G1vzgFXrz1arDFtnMWqWNrjZlpWpg4rUfkGJ
NGGsGlmKRDrxpScYKlQcNemrBVxs19KQ3gLpBNRokoMTeFmDpO5UAkKWpuPVHAi4wafvTEOwLhW6
wzngxlQcRXKQFYR9WvKFhib0mz5HadAV2T+JID7NV0UF8Ydm2Y7APoYg72oBQPHbYdPtOFzq/SyK
ZVaEPFOAfKKLuPvplTfLe7Ze1GewOIPD6rw33JBo7xIqcNPmE+X0dAh8CAvYxaCZcllZ6IRs5s5F
OtxOK1wo9UvG+jvW8aMCNYbNAhX05G1Wc+RTaGodLSnA7qhIg+vtB+nOTJbJiiUktiZvZ+IFsgPm
TISaldD+f1ooNIMnbXsSaYfh+UbY7ilF/qEIrvNsN97NPCRw0J2CNFahvj/JTxPAhSiZv88y6XOW
RfUL/ZvHXfry53IND8N4buS98sgEdmnchg6P4jimWGj/lzNhNZFCxfOxMlLyZUZlFBuCmXl6Sun8
OOQ+sSua9zHMbySXHukCoTt+Xpea3DiT9LChdmwZNOkZvgmrHmfAVr06BveKsCGm6GFyn3jhpKD8
bdf/l2DgtVYUSi2RYr1yz24orXQM5munLAyaPo2gUqlL6rsFjUU6zi91i0XRk3qBaypsj2UycgU+
b53yrhcrKdHTUo5CVlrXWOqWLcImObwufxoZr/zdBb/1G+CajXvBjcSzKS1WE9f0szuOoF84fp1m
JwcDLBgJQJJI4Exz6s4fubRQxAhLs2Mg868Jp20qw0e+iSGfcKNYCW6Rs2KWCxpBoJVocYdMeU8+
RSYUnWtih1Cr4QdL6GbyBpoi5lK0IwpeXua5/SvpPcd6mNF2Et2GGbTGVlojB0k8LAEu5nHmmJ5B
rPrhSr2JqE19jC26Z5StqwIzRsVf1T+/cdJeeFLPWy7wpno6ToBUGmWqcxbqZA0r1r1ifGXeHF9V
KUv/+XJYTk1+kMG4jgriJscCuReK5Qi3+xFr0h2iOkRorNc2rZJhHT2+I8/gdMbTWaIWcbMYAYcV
H9U/yMgsUr9NRmCdmbphI4ui7J92QXQtBLqDUWs+4R+0xPukpcMFl6AW5k6ermlywULLzFsBuEHa
r891nFBfrYuHLvW8PG9uJbEIar9zzroQqQ0Ybmtac1YbSjpz+ijxypnZfCCZP0WdmVeL4QBc0fBS
tdtd6j5uKF+F9C0vt3E+/IezIk/XG1ns66+f6NGJx3wUAOc4wqhkqhOK3reNmC1r0ndSlt1t49xe
LBKRzHiWoSHp0SKXY76twaTn+zMnaiwkx7urNY/OPdGan/fy1gnt2kTMNegfbWsMZ/kecNgkjHH5
f+/2f6HiLSxEIqB8z5GJ17CG3izsYyTH9QqFuT3L9zfF+0j1z4X8dZOnCGekezwtJ3RrqN2NgN9+
ULFWSolhnRZzFbamLFeeEL3xrb9YJDVadAWYslYD/z7DZdHaD3P76EcGSoQ1P1qBYCFahmOhycqi
7YeswLdDa+Kz1XIORYdzxpQdnvDD49MgoTAO4TXra/aOlnuokcBEsoVsSHhp6ds1KgYi5+uIBY11
kFM2SdYwwabiCPhI2yj6nh59z9Q5s/I+cSXPpU5CSf4VvF/0N7cF8B7rBggVJdxyV3nQuJp6cbsI
JxTb0h3LKoaiNiX9TVmZTWWEZlXs9bUsPCkq7UnVDGfWyYp0+vQN4bf/Y/2s1eiXjZfpvwRacjXW
+7YxL0Vvx5L3lTrytAJIXo3aWTYbzC+ZI5U93QAjF5VQOyeQe4J93hrXij+2UbnFcnY2kU3LbIC8
h3wUQa3l4tgH8In0r2VTVZB/uEuuLpBlXM2wcPvSuR953M/+ApHdAXtE8f5NiEjXKXt3/h6T53bm
1A1JRkpt4LGz7jGUbYNYh+wH26af9bRXhliWxjCbj+r0ZymoQrgZQ+Bc19H0grqutmgCkk/miK1G
ThJo/gfVuqgHJDtO3Hho5RYr4EGPBEdi1iO2Vvz854lJUQd9ndWJfFARzgH4bPfzHpgUuDhBwInm
N6+QaZ5OUajtnmk18NL8ODhMMHMfEp1WQTAC1xIDTSx+kE6pLaZs3S7YgwdVJu/dgsvUyQHQ7erM
ZnHbymRWIQcoOePQlvT8ydalf6uy8tzIZIUY0z2JHDlSpQWWvjJH4oDTPMiEQkxmbES76CiVJm0h
/YOIcOc/JH8GY6V7GE5AEDoM/MWqbND5p6h/Mcqs/FVlXdh/XabVhazR0PzYbzVIgDCutQFoLjOD
FgOU/J5aX6NSYNFL+dwzCvsl4+GVjBMLtE6pYUZ/+vObnzJ47vxQNcNP0O2W4wLE9pFp1VP3lBFb
F4lHOLeqfHp8ribypkEIujRF/YbxDx+W3XvqNVZU0x2MHQ8YWH21QL8YukJ6H0ZHXA82QhzexR15
eHjSjw20yvpt5fsnW1uF4Bsv5n0upxi9yiVODX4vziA1tt8IGkfhmsQtwC894OZlhkRkMOsebrgf
2N2csP0T4I8C3tiymprXp9r/75Evy2nnBPQrY2q0WAkMqrS0LKtCl1W/AsG4AcpxMljs6g5M5zag
qrH5AbX10SRHFHiNsEwHAb/sK0x0e707TYqoAjncb79M7aN0QTIbYnNgUHr1ZF+U/xM1lzgT9m/V
DGb3Hii4BohSP5WqzQOIpWu2k0tBX4jKE9ecWdAQkiGdQPAsvkZjpVISRTLDZQbQ5rd005tRCcPX
H4bDNSDBhQp/mwybv3wYKSGeG1O62Pu7KtM6RRj/RYZSiw1s0dYVF+eHKjbGBKrcjpIsgXfHk/CE
ezzYuvztCudM69uOpTaIiF0kidS5na9S7n5/qarBZkSzEN3/mWgV7hyMPBSkm74r8xY/Vy8BoBvQ
7jpjwBqBZ931i8bkIv5G28yERhCNwtm8WeTBDlQ3gKhcjY66oAlwoQGeCjtE+ng5fshyArNzbKl+
QKzcgGy1VOWUJUmGdPLceORx1aBrGv5QrfEJFL5SSw4iZSqLLRiKW64KuC6q6Uv0qOSFvvi5qbcf
NUwrI6QcykLR4m+iza+6IfSr62LXGyZXw26EZ4CP+mDtz6exvZX6BMXQJj0LE0xTAzYreZZwYdXL
EDibbT6kioZnMoOmheayNOg1w5fTrUNFR9W8r2mfI6zeAgjfL2LSmfKs6cV0sANr/2NBOqwPjdIE
48xPuuTGeqs1NCggbNq5cUD262datJBhuZ4jMYsws+hPUanmYiJi0bMfr1C98IEQ0iIUAmSx4690
VFn9s1SEGujhDjV4kdRyoYUt/0adlxtH1m++D6YV477dIzJtStydyi+4vXY0+W49VglpOQNefk3D
QwXJwzrCPmXRrnlToEw6RtIvJ3102bfhtcvsX1SXaFdlA+Ec0WpB21Xccc9MwaU4WfG6+noRt1iF
eBG3axslFyjlVchhNO82MyI38+n9WVpwZpDC+7zj1Usj8e/ztazdARFwRzhgWERTFrixe5kDmagX
jMfeDmpGzaEmbLP6mpJZwjA88sQvmK5YGUyNe/vZVioZDBfBhJZs9BS3KLQ19Z1IxKHOFfELQCOs
WhY9pqt0AEVObCb3PuwKy/zWttIMDKVTw6pV97E5ijBp/Hx7dClxqZKljHu1QG8LYtok4PA5k3qT
lrn6xrby3MM48dopYauXhvEvhWBFkltBAs9O/VASnYJM/i+ZdU9rqAQ7ATvkxc5d6soUvLPQTjWD
c8gwUHwIvcfjz11wumr6vdsi2Pt2qzobBTlP/k4H05su0fY2NRWnGozm/7AM9/R7Uw3Y474IEqW0
JKerQ3WEJMatoRUkp9dJ4ioC5DCR/wjl818W715aOr0wBNCRHT8kMXzNm6IzvjsADAZJJOOIZamt
bjD9okiGpzJrZTMb03kVymN5jaj0ghUK/Ej9WlwvWjLJuW+K3TMxMUY0NTa8Xglor4mUE4mE0U4n
Wyb6hVKOEV6iCtEEUKsaEHyHOh/VqZ0V/7ALeTOqqt6/dzxnvdk2NICXKnmIRzV84MUPsoKqJXhD
gUagdi1OwcGuPChco155LtfMX51msjKn8kOPa5bzaw3Ff1WjiMaQOs2e7NWgxXzy1ZdV37zQEGq7
XZitoy4rOoiI7I0rjZu0AFiU/0Xfiom/Wbq5vD1+KaSLAkkSFQsb6JjsB1FC/iM0wHnAjQU42bih
PJrUsTfbTIArrRiJmAWI7Q7jRC8MiKVlUHXo5c/kWO/TqBp6P4zA/bLkJ+YMMfv9p0acRqL7BdCh
6rINgpVg0IZb/ZnAJOqmObdFgKy4ZbiAL2wnfihv+FTviaeRhpmEQWJM47fThmu1OLNoFrEW/lfK
EAR5QrFOMI04bY6yrNvy0niqU/Xn4u5vX//D2JOJkzzCTtlfqoHvyEm6/pf+7ebyZh6RuusSXXDD
wOnljMtJpDkD3UZUiebkkrAXAugAV/bBlt3a8sIdy6+TzyfrpUxzYLw5Z9BbYgSgf2Map3fJ7A5T
IhUuX/M15xjFQR3RqI5ZTxdFzXUXff5K9HMXKI2qbzPUpL2fkMnyYE0u66/NwFQvGWGd2N0c0/Yl
Rg6rB6+d6cWCES+cYUi42e4UEqiuldWFj8J6rGLHv2ZsaRSHMUD6Qf4YFAVH8S5x9EoL301jS9xV
a5SdQjIu2+8LJXpYopTiqmE1BBTU2MlyN4LHxpf9nplicvbZmmMQF/ERTsh8CEa7/m8dcCISpGE2
XWevzjcV9FQIOGNHXc2wpwBwEQNVbZB9DqsVK9OLeMWO3GMDxA2aoCvo9RChIYrT9ul9Q+jVB/Ld
IlZJ0DbxzYPA4P5BwxilsTcgrxHkEbQl17i8iftVd2CxtowiyJoB2RZ4dCbNz+YYO9NOyMz7K33I
7Exoca/KeKwh+FUqK89ANQpsoQQ7Zb1i9YW7m+uI0kh8CHVovufjGtR6cW4v+LgeXDZKHGSHQZ6O
LsJub5SefVMboGDImjbA9JxD3x4cfv6kqQyJLXc5DNtcs1RogAjn7/h8K0Yyx8/1AoycYvCEQxpR
puvXA4IZdaKs47UuIYqM1xafJyY4odBr/LGvDEIPm+7Ot6ZYCpGW2hYojfwUIIXZhqx1lfWhnQ9s
sxCQ0WX3KjOqIwq9pxfkZJ9uZuVRlVYvFAAPpTTUNkohsH5HPyUs6F2KP/mbbf2Nl+i68OiNpnrF
wy3hvoWoE+6AlC+Ao0KzobkzrFG5JHkbzJXUI+x2boh4Q0jqZVwjny2FypXpteG+2w27nh8sg/Av
zOBCp5KRchuWm8BQICYnZEBS4Lch0c2mC1ZfY9p4C1yeTtg8IdGRDcvjd3Laue7xUhUkr8Gs6VL1
LcdAiDuvBCSlDL2ObnL1G2lJSs3HCQ7BEtYoJovYcVzfHRzwAyWqkHODPeh+HHEfGMN4TmK/BmNb
l+fFcX6bBwRj68vmd9cUHKyuoUbw8p1px7r8JXBOLVBIyJqKDdvutRMxFjGb2lSI0z0bbvUcEPvL
FvEPR23DTt6BKZaGT1D3lYk2Rc5Hll8v5pbYzKnFY31vgcsVCVYaUd229XoHKp/XPVcg4vrg16cW
kPTF3n2w0tPNIq3FrlcL+R0wM8s4S2pBmBemYRxBTixGzbUlG0XZYPIQuVs37g3PP7zwVLu/Tqbb
ir8Unv4lOJk920xLBRF3mFMIiNOoFNAzjWP/kE0D8MmY+JPaI4MDfYKeU8xF59NaCfKexteB8Gr5
/0ku4QltDap88VKfMNpwCCfacB6GEwWBxw9OMWlB3FwIjtHYnTtFZnxFeErrRvigBi9pKKCophUt
aLhNNOiPLRlHp8xXOAmIEnb7VzVytFGP2bD2Qf8Jk1aq9V6wF/xXH2pp9MSmvhUlQQGmcLPvAZQw
EHR/2NuyEFw1n5GLE3o2/oehNHtv9/KrsKDvkoxnTxBuWEcadwtzls2foywX24eWdFKA6a37QZ4r
FbZcrnsJzBWbiqv6u7KmybkCUcWzT0Xh9xQqBig1t99jS89lWwoY+lCKwDCsbGBkC7nZeUbqUD9i
DSaEYAhRKY8UQl5u8pguoUITKdZ/77mnhMtHv/8MfQEXPD+LXovcFZRrtZcFLjC6octuKN8J3zfS
yHP4kc15m7SG3He2aoGWt2zMSOIzGnvqG5VbgKY7Pqzw4eYqweQPvaZoE+Ncp5AMQ6e8hO2ztDFz
87eTOyPqPqFN2lLUbeRk81OCA0Nl2AurP50B/r1/Gn6lt0ifbmydHAElzRwxkrRJRUtNAXQEGm9+
vZPDVPSXvnE3Oss96s4p1Fcd+NOaMYZwImhzHx4vG3UpkGJlqYEufhf9aT5VNeBU7h3yLaSmv5vX
eY5ipQWzaCndqjJb9rb3Sn46r8v6LY4wSS4bIQlgWxNAC1tFNUFo8xwtrHOkxhGeDtzXlaNTdtwr
cymy/yMbCffaqkeRmKBMyvB8j2999dZxBSQSw7fOK9cBacymEs4gavSbmgsG+c9ZC5FALGQ0ue/d
d3DzZWuBQFb1LiJZo9LrV2oHliu365I3gRGpXMNV18lIRjcuzpxD6wZF/oiUFvdI+3/vFEXa1PW0
Y9GaUp0cE7R9oDarIITiUnOFBLiLmz7bv8QpiYGzj5sZmYGadsw+b8HsXVlRLJ+ecJAdJGhMLRl1
gQmb8RwZEyjOCF/Gv54VELUF27f2TILesKnpiUTLnEdZa+E6K5PICKnomQVlKYh4xmNKjjfESIFF
P+2FubyLhxDWQhwBTpVp203fZyhvsn5zRxiLB8il36ohAyJrO/xdwAmjGtSHcFa6eF3vuc8TJ0/Y
fnVvMHq9lCCeaPQwauegmj/h/0f2/VmyOgx+euU+CQ/lbJv8QOrcCS9fNs9p8uZCy/um7CWX//hs
0Wq1/9CCWwl2rgOEpryVnmbVP4+IHgh/9wMUdEqcnG9Us73S2I26afWs32/oXkMSc8TXMhmrm8yi
PiWU24kLwcbc+Km1am7wbPGRL8TwLeiq6pUqd3KEkolbyAUPV5GbmyLZ2vSkYGEsgq0WSdMSkLxg
KttA7hWQ1gR3wpXr1DztzHu9Nxd+usYNsabX1ZnAji6BixNMyQCzkJW2Nfk4uv1ptEEsTx04fos6
zObt/4QiHblBjwCwblv/WIK/84AwLD3ghOfMifvSFs9vxTJD3sd2RAfAwt1/QIW9Vwk2sz/nkdkr
ekx55zlfA+KzFKaIyUt6St4WFXPCMw7e3RoSGwFQHGebbVWwJw3B5YAtDDMGz4rHUQ7dS2ZDN8MF
zjFRIq+cjtaauOmLKRKIf0pswQznAdykKBSSuag4ZcEkJVahKlAbtHjs2RmYycSvXWE9vsWybKaM
2B5fVx0ngKrImhuRSHKOD7PGdv6OAKvewv2yADyLKeytXGszDbLKGTqkx+gp4jQRIzoNAjrKN/bl
uNuedppnm0S5cxu7u/VpaNd1qoP7qz2aqAYWYogMgXZnT5bn+V9/8cNvXSciHwOL4eA4gVMdu/W6
O23Jh4jxVWPXFv3x+R8XKQ8948n3igfPVpF2tLc4NOXj54UVS4IsqOT2lbAw9D4TDdhlrPoW9sJ0
dJrYnKSqnLMEXflJ4oaR60wQ4ud+lnq9LpGMUMgvkzK84+Qz7eyNau9aMtj616exrzTJrfFbyK9o
/jE9HZ8c3RTQIWvTc4XpHLgPT5/faB7wRKU4lqpok8DBLv8CU1aYXjWP7ZQOza6VPV4GoX5GVUF3
roeP1kl6FTfP+aE+Dclxc/5m+XBPqetUPVgG7fs6Bw4GZydc/Enu2dKGMcEC+D+DajghwFSOG0jF
ghzwqvUfJZH0b9KdXRGq1ZouR33KL1LCl1+fhqmAVwSLtAXw+JDpnSpEtJI7SZDLGIAcUx96bklm
SiBWbGHWIqnMVQ6N+iu5SSmKETfitDNYKNsPuDXFH+Xk11SS0SvQo5ejJ/f9y3e6ZNfdle4ENJoi
Um4xCC3JGtJ8FNCim+2NC+ZwvQQkUxlhMyuxirGhYQdO3RhRXxJ34KOOVghWIy0b/BWusVz9foUk
HIBXQ8jfteevpRLFf1l5acd+0cuUFiQKNXQBEmAj81Qj2hPdhIHE1keJbMWZAn4UC4KpAFogxaK7
pNT5/fv/9dlBwXbynTsLaJtyFsgTMWCb91zKZAqDDqKNLp7ogUHtSViuob35vsOO0oTktgWbGJds
usI/LukacUHS0LdqTbsIv/X3kYcDVo3Z5lIna9ntmr2i+j7FHN4R1Y9cU/KKIUUYolrxeSwVz7+m
0BjtOkCz5aZR7HsILq1nLIDiwrpHbnz8HBJrxIqF+ihynm5f6KeOIsuNAOF/ugkfh50hhH/ULG6C
UEWdENjtOViTyF1jBzKwMqBizNlwzblMakVxc+iKBnFNWoHZjWcL5vAMzS10vOWDYxepK9tKQQ6L
y6g1rxo0go13AsYSFUe7CJRJC/T2befzeOIwyVIXG5Lrgte0ysFkR7r9khIfBLmOcclwpRZvE2Oj
SLnUjYcJDjZgsiWbBytiFRbpwK+L8cJH9tqfIObpAXqgc1YUQ6Tpjy/SJrEs5QKdIEmLcYcq7F8h
pC413wS1F+NSlR/YgAwkmAgIX3nOFgQxR0jnVAF0eS9K+v/PJL+UhOd39in4SHM7PJ8SJCnDrgjO
mDEB1QDkOTZJtEpwj4mozuP9En3asyTmYKiYWVbdpacqRmTHDPbQAHeT9D9l0x/xO+PKBf93hOC7
PnmdI5bjinoUu9dAGKMzZ5xKJOMqTqGWc51WdYK6rT7XsoTUB2uMvw/1Q+2x0+Up1jpKrbCVIzB+
oE4Z5MxxDVELP62VLrcgthOsG0VLBjaZ5JowfMF8xLYnxkQ7sSo4rzPpia2C4DdH14Zh0Uojnwse
uYtTlQEnw25yjvJfIgiLuei6JswJKTPxAQNVis15ex0e6j87m390RKCVDo8L+6gOwrB0nHZfq202
0ztAd57c4Jao086MktAQ2XNHYY+VqEXYAyJDGK7MrMxC6A1CJQt42etUX/lOkDzYJxa2jQGPj/+F
x53jo07UDOXQM2HC9ENHJ9+zdgo4KMy/9CNW68aaPeQfeG5LC00+v5dUgYZh4GHgsvLiCOthaEy0
2Bk87vB1BjTroUO+IiMqUyE+h4UYxbMWv8Leew4JXyDLgjQsYubL8TGBRtTkRbxBHJpGk1E2F09R
3Euyz12ZhJiJ6SARZucSc7brtfDjz/jT95aSF+UUfy+E2YF5cqTt0c+bHbjVAwwbwtKRBLrNB/Zg
pFAubHsL8UpKs53hwqR6EiKhfExpAp7ixcQ4B1uBpn7TpLHTH/Pl+8jhUraYWU+REJkBLnMvR6HX
bJm6NTAD5BHBglVwNDY9Tj53OPCATL06VwcVttsw5Fxi+0IBnrAD6oyRRkL7AqD4QVXFp+J9rALl
67WsaW55EhEd3++JD+hG3HOTnj0kUQhy2jxQyV9GJ3mVknTjH2ZaRo8idoHSP0luu1WrZAEz31l3
l3EISEGf+6hUTAaO0Fpp3fpWlqjMP1Gyy8UVU29tu7Ihp9ms5eJJ4jlUmQO8ThPXvRePCsZPe/wR
l91rLw6vPWDzWzEqLRJCGDma2B5jbBadcuANx60a3xnlB75CM9hYZW9kE1yPZT/lx7zyNJBdmJ8M
GOweZpLVeoD/h18N/ENrWFEG/Dc0vJoWVlTbUtcn3ifVZwFLiqtVskMeLdi+WedoOHna81H+xZTB
DtVX+nCu2fNmKsxdfI3gh7dmGeE1L2hCLYWB1Kv3c19ohozs+X7oT4x8ol79BwKSUwrGNPZNfbk0
WNkqIpFrGo9uGrmUh/iSHLAnI3W1vn62eAcKPsJ1d13NMm/uvrS8e5uba+2duDS3xU/5Xx7R9fcC
PAUgUKqdDb3Pzx4wFas4pmbzE/Dqx+/W715tYZoNRQeJ8ANZDiC4yxjwqvFhW3cX13Dh7j1xH0CS
N8hTSmGGuJybwjORNRbnpTryZIQv5myrLYPFx716k4lBv6NNa23t888wYJEeVhJMo5l23YvYGEJP
gaL764PaS/R1u5jEXI1J0rhhnIVrH5J/RefAIGPDOX+rMkazDEz5XQyKPZcm+7+nNRZNFrrqpcyp
0gAibIaTRgveqPuR3PcuAh1cHouIc5hJFEHmqnFwu0mJGZ+ndNk21/vEj3E7pwPUHryRVHJSt9Qm
b8y8I8W1wsFgytSzzc6h0LfZFZbqUGJidtFKq8zYn3N36b/VBqyGiFuZfAawsIYycQ9L2zKeXuZW
V9w/vylzaMfAb/RZDGmZPVUELnanviZVk/hKXtTkWIiAh39Iou68Z3R0FR3K4B/vKMLyC86pVUIW
sxCw2iiNUnFoY+T1sPXxCCc26IU5VUwwloO605t3YLkqOzDgw87wsCIHCkHUtuaEds5FcQy2Arwl
HtE1F96wCCBC7gpKewAJcfVh/8yHa+aLC7nuXImLo2dR3hVFtjLVCugHKI23mcfrYxiZS3B5l4VD
5kuQSooRUZofoJfeb6ziNPBaMvz8krvYnmWTLtamr5T/hGsEfNYTu1wWrHfzTsWmwqChEkjh0bxV
qVRtltaRmEskt8+QZSMHkm+yRYF/+Viku8pCLsMVtbyrSY27xzN2X2H3qNfAXhrCaEhC4rI/VS8K
GRQUp967CAIjlluokGc5QFHqdr7sg5357R1MTxsx2OLsQEAFcG4zecSiW/zuaxOhW/I7ddl3nXSE
PJolYVDNKGMvJtg86T+Xvyrx4H7UUZTievQ3NDaJlAPnCPttQDGBTrWh5RE53TAYjolQIdTl2WCq
mN4UYIbaTmlB2O7+ul97sqkxJ6AFdtBAtOci8n7CkSQSQZTvZ7B6OWwLmxCzlATHgKIWKL6sC+U1
a31sWN7wj/Zz4MSbRMo0PT5UhfnqK07JmhHontkBylyW4wY0hxWKnWwMjoEqHTNqvq9QPQD+KH5G
MRgQhNJfCAdpdGCn57yTpz1kmx+RCMhlCHMdWfgonevN4yVV50e2Q4/xgjkxzvvCtulmfXf7xGHy
vRTyTkd8wqKdUNvcAx3tZZ249E+pHSCDZ9vjD5X0V38/dz38mf9nF+SjJZB/RQxYpcDxm39OkDyK
6qVq8STLboi2ZGDD93XsJg4BKP++luwYriaYEN9hRsQxm/YE6wVi4Cfyc+NBH1lBO1Bf+t/JweVF
Np7kGJN06ES55+B7lpFPxnJKUNmDEJhbSCZi0Q0Out0do8djjWNhl8JX46prmibK00lGCl5dr4Ds
33xV/gt8+dLxrbYNwKjJeTZn+Oy2n4VgzhCOus/fdg/1mynZoGYOd1PjyYwbo/4AgJ9LlXY51Oml
qu0GhlS8Z/XFBFWruwkgK4TbIkJ4zvXBgZc3IFIzILuXOnmMBaEcqZjrcpqaewekTV4ec9vYKjkQ
8CYYgSGmLbLoLciWLSd4yxCxiGFbtiizakWFAAbxJ3zs2fv8e8pV1eLQtmIztwCm8RO8q3MDkSLp
QNWbCBEyAcrhxuGTUUdVACdxtt9zEGMYE1MyNOyWtP2ObQY9UN3mDVpWVUltfW0OkxvTLxkupMS5
WGQptwcyqx1vRdr1IaDxKY9stVhi/rOl8079Lxc7ap56UOUbCZcnCse+7LNMI+KO7Y2Dlz0iQtm6
kqMJoHdRh5kL7QD59CJHAe4btzjpc4UAwEjAJc540CJZ9pY9F0TQlLw2CeSkba2+eS0Uw2dpGzV3
XwJA9xkp8gOfPKGObhLtJVMNGN4PO/xm+Mw0Nt3KLyPJClSZjtVo7QRJf6xkDvEh8dAk1aHZ3HfX
0YAR+QzpvsqUe6v1AcfFQG8BVQZgWRGOrzKWnd2efccMNL8OMpSmiPQWtIeyti1xRCBhir1zRppS
vnnPZG5IE9E8jzoVr0aimVwqV1Qkimg7olwiJT/X3q/0tF6IxM7o3WKdrqofTAiyXngEsE2aqff3
wbD+G+uGsM7bBuD/WkzF5x6sCvM2UtvYV5wmawDYQRQZ+UIWA8qxSqkA9IRB/u1iEtZch/LHq8cE
IbfMCQN3TCPe+MQLa/eEk9IRgO3bFPdmNdPWtV0CQPQx+TE4KjMl/+0i/MQk0VbhVAwFaTBBkOYX
DltxJLPOqE+nlj5/n0gQJUMKWBOfZ/NoS6XqAVy/8KrtM4LcGlP3Ip+KamlChY9rE0uLQ5EmxYGf
9d0IXi1uQkSfNbFw6iOVq2MtbMu0HoC6rqBgDthSJHUy7OrLAjG7ojgkBrq9UJVflady1RO6ZdPY
9WCSnr2kQWEQdUTpBtqcXcJEhL/zNNP1PzRSYNpGOppOvee7qS88VSEn9jYRJwzutWTpwgS7iT55
QkAnqD0tgtce2XobH0u4rYzBA2dTaGUkXjWw4IWOvZyWKnz3flDXZajdCYDr2LbzRfEQBPc6DxQl
tXrAkz4VhJYxMS+qSGkj/qW0RTJcUQjznDesPQTH3V20ZdKeYiiGR0Ou/lgoYn881udoYLwmDg7w
sTLci8e5lUB2cgYQruB8aZ8ZNVLgjaDDCsOdvhZvLtd5vYlJTFvnAW0MRSsevIR/ftO4fwwTezJE
pHm5K4yamdMhFIFwpaiRinTZxM/jjWZVF3DoD/2l8hgeB1v747ZHMGnbYP+tu1dNLDtDxADAhCdc
4dKHSKGGmnJnj6thS3whQFDxjeaOvu67LmfTKUwquWVeSsjLtW35HHIhxG5FQef1LqQFXnswDTU+
o4Imw5NGpfrIJurTNhswJkk1Il+tAJJbYAr9RpKAJD0eOjt/xsn+wNRaXT/3H5X24DvDj1EY/eou
dXhW+Rf/IqRsQfDiPFnGGNcZ2YZakhLFTxQzl7FrPT4+2iGi0qGxMSDpwjVXTs+g7r/zITbV9GGf
XOOENsVcqrSG2LhgZFGg6QZgS+wbFIWD4lqeFGze7GR+KkzteWl8G9stozQZBtyAkoWY0kxzahHj
S0nAzb5SEVYZ22NhdpW3/H3ezu0fZvQ2qN6uq1858cDCQewRQzr0v21EVqKFQNReUrXVzAx0kA3F
PiTw6fMf63buXo/HBakzDK8ZMzCbiPick87DqD9MepSsMm+p27aBr7H3Qm5GaNlW1BMCwGppv3+f
cYgcYWYltvmdDuE0Ji0jSfHF/luWIOFba8vnecv67fsVmGVCqeSZOu81hblnATmRu96eFFdqIxoA
vRbYbHcQvktppfY3FIR80Z9LPpYnSzJQERA0L3ELYy434D7D8nGunmJl8vxNFzOaAepG+/rlMpkV
EqkPXMxLNq52Au4tD8KRWMeKEURP6Oh7mhTcw6H2DkC7IZAS+7dChJD1ZuzwlBRQOjJIjRHwSWIz
NkAnYd3uJFy2g4ZPDdnHjIYEgr7yKeKNDsVoeAA92jtfsFYG4ki7+d2YS5sHawiNaJn09x0Vv3sw
YnIWohZwQxjULFYsZzTAZyUwAScvr5ZyCVTbirkUrN8Qh2QXczybSnP0TcKUDfYeN1/xsGEUxhC8
0GTyfKodXCsV08FYj4lpWq0S1doMQX3P334AcfZubYqJjFPDOsDXZcB8TQ3ZRw8XUipRTT3UDINJ
vywBif6Ux6jmIxJNU1fMYf5ooawA4k+A496g+ulYFB4Z0w3Vs4wk8//55TUoGXkpdTxJdYBRa42U
vPk8HEKCoxYgDfx7UmmzPdyQ8UXmfMypiVP/p3+MlticA705ctZyNDIC4HJI5C8nvKyaq1V/JlUX
iVNPdoDUUUiEkyEcZoz3tUFwW5V4dgS3uAgrVo4tQVytnWrVdpH682bkfK+CHWri+5kNSA+1LJaD
mbVa9pXRF2udXH+kr87qH/nb53TNfUluYhN+tpKUMz+tdZTz/fUM4UetUcqiq9E6EuT9niBlfwLR
NIMB7uF5qlz/CEf766pgmZCHcyKX9TZyKyjvRzwd6eLUBTnBCSAE1WuD/0UCWeYd3YC2RkZjRS1h
Vnizc8Sr2bhZjkBEADLuOuf0XbiplrcucYvl3YWKGNPNWuHOWpCLlXrHgITaOJs4SgQBY8y2V+bI
njBTUTfck0DmXbtwy9wOjjs0e6HnwtHFxbMfZMTylRtcgo0/S2iw3gX3DkD1fhsraJFXQc6nwSuP
iD5t/oUCNrgPrbGAFyVAmavlj64oJA98sZI1eaD8P/E0GeUR1krqCV2gB8qjiI3HBOl5S2GDhfkO
xB8N1lhQdBeLRNCazOG7TzUY3NoQijB+XXhGGWCP9uy/gUXLMOe5OSWJnF/mwN2DpNJEAJwoY+Xp
qOLZGLjTh8InyTImqJBzOv9zgggKDXc6ZmOIYqHrZnjMsUNP4iNVNerXvlvswG2jrnYlHxyafCPn
6KZrXxWjJgrU3wbQ1yUJ0fhnThXzQQ8rs8BwJVJYjyz0xrGGr8pmk9ZCWgsuAj/cIe2ibn0bvD6A
H3hlrrRUs8kajx37XHdgbUpNF2t0fcmU/BygvcQOqGwKXvj4g2vuKXTFTIo11m+V3GtkcpsG2624
gLRzcAZeG+AsvAzi0BDmpf8hmxIs/pwR0aIw2gc6CpYF2/AwDsU+K252oz97O4k/1gJ5Lx5cakrr
p1OZSRfJfOZ2netY8mwfTTX7MiM6jkp/jeM2JHvzXcNO8MJ/sQUmrhCyKjKXdq9jQlGROL4/l1SI
ahrVVk7EaEvOrHp27WwU+DVYWb73MZ+xzeq4a38ngYypEe9mon5dejJpYqALxaHiiJrdwPkK4qY4
Q893yxpgdEGM4PZHdaaq12B3an6Ev3Durdho4JHSsp8VMfbXmdVMhsVAWf8ajokQInxXNHtdf0Db
pjcjrhMCK/OrHLLPG1UcIAU1L+OO69WTDk2+68CC/SBtdVOxDu61yaBfUenNKwFYei+9K5x2AR7X
aXaseub+JmXnx3rmjV0dR7txYTmwnCfbchXODfp2hgC1Zkv8d2GAQS9VK1O/M1V0NTwNvGCL7p6Y
V7wENjC8KbG6HoqGuO+l2kDvXX7yEPkMibXttEgcwg9nm9UNhjiu59cf/51Kq/MET2uACv9NIesI
USaHaDSdwp1x48qhyRlfyztNnvhVabizLQ/n5Q202M7/VAUkWXc3ipFXm1c2Yfy67QRApH+ruFBd
tQqBafRt1LH+PFCBP7VGyqmhgm/rJosPXvDMC0j9Fh/g8GsSQ2n3gxy0lzSHGXbjHn6Jn2dUF52a
LWRSZ7H55LBPK7tpzR+XkYYGVPmSKjn7Gb+wMYja1MPPY9nezZIi+juAp8Gb3dr15uzNo+xBV1ob
L9esdwhqdNfkM2ZYLs8olpVTGpIVIT3AAinptQ9cWkK2Hcf+Sr6YHAiG/hTYKX2VesyltdE67/La
0gDAJllQEEi/r4rxu5KsfwySzUgQaMYXGXq/y7NxYrHbw2lLENqNMlDU4Tq+WsI9yYmc1fQABg0/
cCrsORIZPyhvKm3XVB/wB5llEByIHFCNVEXy2bYgCpGUbIrdqhHqliyiQbo0Exx7k4E19tZW8225
BxuSj0QfTQYtSEJ5NbG513O4YeIQUMdA0vm5rm3+EmlvLmkinFX2yY0mYTvAk1ZXTxHDU1XoJ4gN
cNJL4ozcXWTMgBgZRUHM6wtx0oQ2km7mimnf0dmNk3Cr1O9QvU13YOND8EGUG14fKF0eHwG+YqjJ
mdlInsyGaxFeSmcjfUrdND2bpZ0SuSVHteZ6JgistQ0sYmkPYvt8j/FJD3aQgOuVqH2zE6C8DyxX
KyTeJRzuWkEdsPfzF2oD7KbJ0754dKbJJT+SEzamwRI+uKcf1+VMTUE+QdQFVOnt3MhxWHIl71Fc
CqB1Q08jTzVw+fGlpUIjkMskHUwa2TipKPkKTrQtaJUTtVvSlgiIQR3yarBCXszgElj6EB9XHg/m
YawQpgf5/cvSelx9lydFNmkPvIYC0JJTCVtfsrZ294Z8twpC7sjjDvYYYbEtErTKtJZJeDZGAQQI
xZW5axSTvvBhPp4VVhAdm/L+rFB0JHyvazI2V9WVxQGbtUiV/PTBr1lZuIMLs9dmzIWWdJWevMau
yH9yanIHpM2Kldh+Y8pxXSrMhPfGeU/A2XqTgu3V7Be9QfsC2IR/vB407KAptiO+uBjbERnWvWi/
EyksRdm8S+ZAOijS/lk0dkAllsi0bVPji4WdEWonsxMf+lgCazFqj6Vu/7K+4OWUuMk4NVYBkloM
OAvuNmkjGO5vfBfABqBEZ/or0s9ZF9CyxukHkGwHfKIva2ycO2cwllLjvucHLOiOLmvQqbRuOS0m
WmWdMx9B5wCCFHIaH3ZboKsR36WnLgSdjEmUxIlljUYuFFF06oStGdzNrgYNt3Id5Bbo2MIrmSgC
tpHilQyt+B0PeKUGg1bp1+GwC4EiDwXRrr2+rWlVkB05CrFiSkZxhvdd2jDpzgfRqc28juUSSO/p
NX0hgUXnqyyIcs/QCV0ZLGFmcqLxfwrmWx00xuMvRqmRoBl9k8T44sdchwBUttvf21h7NUtbSEId
qsNjOMUXXBv3R8SsSZc+06UadliWntGsiq0ByS3J27CXZdnX39GA1urwCIjWjDxe62ol0O0UQ7y/
BTEJHSCwwpyUHqi7+etSR+jNpFNzp/N9teOqtjQY0fJVZ4MRcpVuKPo7cYY7MNzrZgaWA1fCoXxc
lMVs+TRw/QQp4DRAbEw/H+EjrTMxCuyAlG/KzlYog4Oxnkq4UZPUa3TvM8wgguvMXSvc6PCucsnZ
C4del77/e8w2hiPE/aFHn8IWPoSq81bcvC/yo/QN/o3e3dSMTEdgQDYF2h6TZGENPFATSN3S5G2W
YfolJpcNPFRMF24Zg8yZ4xBwAnBQq+vTl65Gsy95MdscifgotONWKG/GD8yLmf2rR8hNHG/4pjci
vG79Rtj4fbh7SZo2NxkhgxJin857smkbiuqBFsjXMzxhqXsn0iQP/qmOUFOFAD7K3ADVUORmYog1
meQdfC6p9P02MwOCRdmlCjPh/lFljDPaJwBbG5CMNN2YDfzeGGl6RMC+Cy27z8pCxD4rN/KKOQKO
2Hwj6DxADsrwsj4bd4cqT5Ax/mfvRTlvdiUMMUsRF8r6yNwdAZUpYHkCr8yADwUtcTqVDKiuCeOg
TTwefm+LmyTe/z3C4shBUYVKFVNqxit7KgPxIWHeamSjRDltwrose6OitrZXLgbCCrbygN8reUm2
wqa1e8TbBHjJEL3qCtcM0ZrLMihoKrfyCMVE2Z1jfKrKwTp7wF7V3aTLK2nJrC8qkKVoJ3/Zhhrj
RdbKwvFp5n0WLmUQLo7S5bGLOMQqa55sw78OmYykzhLfgqB6d/sq0QILG/FDb7JPQ1BmSwweavV+
iXHPYjpGT3v9JoeKlXVoNtsDzlUsK/H9gVFml6MMLkUdoa8emdtboj/VYeQ/YhEduXclFPRkVZLn
+NXjlFy3SxIBkhkExcFWX5bODtYF+8XwEueCrTpIF+UGVdIcJVM7EaW5hxo4q7Qq8WMXye/dayxm
1Mn3WdVGRaABS369L5o2uoHdQmPl40fZyxB75DdZo5kvUWqUe9nxCAKgxzBxO6kRj26548aa95T9
FywDAi+Cv95jBNDGTVIEbSvTopyzXIaLrTxqX3zR+Av9Z6A+CWSa9g/fpt9kvONhjfLUSNflhpaP
lVl7XbLUvs5SFug7gTb6MY1bW6lHzDi0tXmfFdEofZNJV+a6gKPozedSLonL5q+ZCXDuF9Iw/K4O
8h0Hw0MCi4H276xOgRIkFZOTaLFcWSWGdk/UMkraeHeRXXqnvRPeFnMiABhYiX12Q9J8n1RFhqaq
bGAs39aA4kRU9H5XDvfdRQgUrufIP+uE6fuzMo0Ce59HT5VZoDNT/BfYJ5tT34HRiAKnSxKZv3oZ
ffyRX6hRtujg/bVj/IzTMMhzAoDN06fNwxD++wtjUKRmiGiWH9Xf5cCWV7cJ3HwVwnMs6JrzaN8d
j8HScUFzaGdWELkveCA/pfsYuYwUBHQ7oqZvgXNOJWtubUAE9aYbipLVtMrcSGDUST4gUQz6zMlG
0Wt4I5EjKanaW75Bn9AyfYwLRXs3wguPdKRv6aKFhQSQDx1MBLjB+gypOBOVtu9UwnfIJyCLuk3D
m7780x/D/b7zyIcO2bB71zNcxWT3mkTDWoNDZM22b2L5oPaCmueKCDqckp2wz97nMZh7Kr6h1ny2
+7sOYjwr4Jcl261tU5jPwwXn9QT43QHJ2ECQWeG+BmCD01G6y+OVyDnPB+plukDZTh9gMTXkzQuR
2lP01UEw73LPSRdBYuChtrqvpOVp3VBos3SYE3opvaBEy4zOtrucA/NGnPcOE7i/ME4wSME5JpVZ
11gH5U16mBSYfaYIsirSsSeo6lSscimGg6ez2VmKS/9LD6D+NjE+PeSEqz+2lOdbqb/kJuYl1BEz
8VjUPlVB+g3PgdLspRwm133ZOpvEN2Y55+g8BVVsGZO6QAsXDJ/URJZTNHlR0DQV5HM+qQkutbnO
bNq7NZbqhXnK0lCY6yTJPZmdZMovACV1nb+gQ081m5hnY0CETP/f1rgNvk7IkTNL0M0c3sU9SXKB
AGVnWFKUkZSlbW8QDp+HjoRBUMg7jD91eN5wQRZ2Qm9yh7PJ9u53Uj4xZub746Ta5u/m4K67v3sI
yJNEZ2tloovOr0OQzmMBdeWnrTQX1LzgNjeaYj0irBQa4YShPCNxIEtL94RxDtTickfI5avhFYFa
KXsgndKvZzCm0YbJCcPG4ELyod21epgL+5V7CeVRFYaG+SV466zDalZtDn6rBlQi9/xd+UIAGrPW
r03+VeAjfiO1jm/MjMQEhLaU5vgo8CZGDaGShY4H8DIe2/k2uhMj7PxfWwR8qPNHJA48N+aRcbpt
4pYEcRfAvCqrs+QmPxrjz3HkWuJTE6o0kCTrbyjpCx7nW/n9SvJeVRaWCIYW3AlalaYbQNGR0Rbz
AvkEi1NI2AxI2AkjPIppavTeGqNWW//gZBxWs6NIw8K0reao79GOsh/mFVFMXuvYF/u7Ox4LuPLX
njG4TSU/hxYt5rpxE4X/WMmMbmZKg5aQv5Wz7dmoYqLk2Bwa2PUOpP/lqsigmZLD3QL83lzXAX1q
7CebQi+aR00WJGduoZ9u7BrYGvcNIW37YWYdFx3F3uSAHtOp5uWgLeGrMwGXA/DPfQQWG4hA6vcK
ZPSP0FFRKcbGzluUa1v/icwTP583cF7taSkFls9Di85cxm9iBajG5S2R6GrXewAJ9FXlufWL94TZ
aOh/Xq3jp8F6OfY217gS2Yt0I6OWYPpsbjeQlhUgvBRQYYGZrlQXs3qllAsqxsoSPVmJ8cbg6/M8
8vhg1N4uktzj5LsMjBJq8hs5u4xE09exJ5dIuyuDafoqyUOynZNySPH4CB9ylzWFgsfHoDYe2B6b
onpyWyK7SUo5mJJWRfWZPsJ4UOhlEwSdaY+ku7oVl1KiRrBhB1o43ywmxkp7KtnrIo5bi5vrLVda
X/5lT3P/FcCBZP/OfsqJf5FbFFe9Hkumym5UYLKDZab+CD3VYmOCeNBcDS/slfDVjuR2996d4VbF
Gy8uNh4GzV3XaNs3dPLZKdQe1JAnxbNmu0WqG6j9r4+BeP+5Tu0iJKmbbxiVYd0ikDySUzfYC4+I
YzYSIg0AGZSUBHEz/w3v2OF3PCPuQjAQfTRf/w3w1yuKxA6DS9n8SBb0ue0nCaOqGtdlEkObwuvH
EwB9BR2UkOQo+hX5reyKgzGDVGz7+vhCrw5JzXkVfdD37NEybsDd++AKbN2BBTAB8LA/XdTxDXjx
IIci+DrrmHEjSPnRcNc/5f5TGyWOpACUnEI2mYb+bHS/2JmiJ4FbvUHq9umSYtKogeEp2BOFLGWT
jsz2l6YO+X2RnB1TePAdJt/ulXnvoG+/t94FLaHr3yKGlTB8P7elx6WfidSTkWeLdZeKUxoodgry
GacdYwap3BP69JV39wGPUY5J5EAF3MqyKBc0nHFJ/JrLXynRTQZuD0HGfr7APKhfCOQ84XRgKaGd
npOx2osvRlpK47CclQcC2jrADPAm1dsPDHB+zOS9IFS0WMKjpMBz6/kRGr/68MsbgMD+Wq8DJQXC
xJx9WajgKHU59XsPa7bpNzTYePw9N97vN1ZNZWU7aibAp0SCRfz9NTB7efWoNVL5p5qjL4Z6eAMD
kUegVFL1qBIY8ffiAMlK6AmbGPi+UrSiuFnEhzUkgDBud+Bvg6BQtLIwaEwNIB4KYV8zpH8+S4BU
SBBebU80H/KUUYpr5BcrfVc/hvsLTfYl0CNr1N6g4uIsKoTFt+MIoLTPsfyoH/OImp3fGb/tWDBN
xZgwTT40AN721UT1T97TJi5qzGeoOqKfoNpd2TLWjDwXgOV+RBavoEpEaxuOZFk4KOHCfvuZPie5
uKfpbh43jk9Ul4frCadOZSojgH8RwzvelRe1M/KAyuwMnlr+BC5Htra2QvwwJsylfAEmFrbms3kB
zPtqiCcXm5y2Ta9aPP9dunvEga59PMGSFQgI3+uO+uYHoVpNxcTGLhQOqZSP7TF2ZlKHTJ2fRQgD
vO3E2QoI+/IIZkvEQmmnTB+TB0a2SdKyU26gathPxDtudG4LS/urqzUMsIYOF6ZG9hWdhc2imEW7
S3l+GVzHDqsqC88GarjxWPFGOmqfCUckv3McKZI7e5CXQ93Zn/EpqcTacWBdXSYWJHRRlvTf5Qfh
TBF1ZQ+gpRJeRWY3kvgRK7Vphk/0hoA9MtZQ8+dGOILcSd4OgS1LNJzx6QLNq4FFbBPzDEwkgu0S
HQPwjmPCPqViDiHbIU3Y8w0H5rDX71f/UfUtLgu/gOwzCbdPUPrkNTXGA+N9ywqjmHZD9otv/6oI
NpSDg8W45oZolIJSUD7L7ChH7IoFvzlOQVQNBnizjWfc5EBRwX2b3G+LDAeXZDAmfz+GQLiXdJlH
9ISj0xL3vzxsxIM6jcLS6HMXJblzb9xHQy3fmNLKb1Rj2Mz7HJKDnvm4cx0ruJF5LigREQPuQ/NC
Zes0QeljWgsniryHph4Kg9nKX4RuExXLFxUnb3yqDqsCd5wRwtThJcj+tmRE85GcUtLNtf/QxK6+
wVoXTdBLId7euID32WlWDgrpcM3NkMKEyNRpoufSpCegcmAmCUj6lhc5D54LxlrCVeCSzhKqOR0e
52sLtGkhAP5ff0y6thuuIuohpYM4nLxeLKAbu9qnDtJtFqjNcG/8pQfK6UNtc/O2TCzMA+DaZAh8
E0Bp0xm10oryCX0sDsQF0HiCloxtoIkpvI2cvYXXQ0o2vgrnmQAadruFTsmTEexY8bammztC2Sdq
KFj+9OI/e2BP3BJ4GCHR2CTDnIYPgC9q2SKVbcJNoMHmKw/APL0iUugABa749iTjKDG/90xy7Dr1
U5tKjBgVe1B+rNcukvCHuYtNhrmnp0JnShuEQAufq1i2GkudGWw/aLSHmLv+itNikF0GxUsfytEg
rC5TbGd1vOQkAgNFa4fImzeBt0U7sKqHypfdNHW1DCI5fUOwu75XCZ1mgKTntwDTH/AacNP6sSW1
TUgHSIa1Es5fLRL7vqQRf0IorSHe3NpaTulMM/GTqs5gKvtSQia5ms1KIvY89HfDKKYDbEmQ1xsx
QlVZhuf9lAg10UVYibSSVl4IxlFgE7CK+/imCYnB2Zde50kj/AjcS5YruNwBWRMi/q4gTI+MPK+r
/d00iuN+Otdauza0ZtCaJyPz5yTc+j7UG5/pEVTvWMlNK7/l9V7zYYLhk5qiX59l4Gp5JLLUwGia
wfCrJqTNdv5K3oHSP91UXZkxaH5vpgWgxQiHTCip5QruPZHxOk3+0oDGl2B+h7BkGjXDG2ztM9F0
zVhg1J1IHazOhcj+rVHc821YF4zU4QL/15W51GK6AknUP1EqAIEcgnbgK8jTXVKP6fGDVsKbGLUU
GLTkMRE5mt+Gq3hiIj08fFHyL4YXNf2oUrw84ZPC6uE9VA/lps76a9nGhhm1KXVQzOP8NPEFTed3
TogZhdSd99KZ1qnSklrjdhWwE4wUPfWLK1PHlZ7IJv1Xm2klNw9QU3b7KNSC2zlEFd75zxH5oCRk
sJ1B68LxzUba756n1xMyGkjhDWihwKK8XVjXNCkWZ8FtIewdWWj47UFsTxgVMF9JqH+dXw9zOUxa
qU0FUPgMHkOTkFRxYjzQwltx4qF1wJ04MKDkz2XZOdU/5Z6zt2YpOm0tiDrSwj1A3wJnmVvEB5Ah
Bq0GRq/qctZlxPadrwphEi0ED4teVuaAm6jUBcwnxACTnfJhfVUKuSo35sRyvA8/30ed66AM/3O/
Jvru+iIcWrblLTmYv7g3UWi3KNEnCC2HTD5T6IjCDFBj5iDmTdXJhNdNRZlLckemn7pfATm3oVqi
L1yvPl89VnfG2BjsbczIvjpnzxfg2MKsQ6WsvsvB2KB46awfUYKopeTdi//a38wGT2HzQdJjq3gf
7HGZYeyM//hfEyCzKdDFUsSjVfUjgKNrBFhOm9Hh3p2hHCyfGc7TzyTOOvKOu1GmGO+ofL/ynqhL
/Mpb+D/Wj2pDHV3jFEqblZR52JkkSC7QqucVJPRmc0FrMdk58Xk4Xo7KlKXzpjsWFmhk3Vfje3lZ
gu8Ne4QqznjyRfvw6sRF26ZRQzfMlD9EaiEmP9hXIhKXXLWMen7PcBLta6sMMLo70zj1EsrkPAHK
lJ8/4b47grhT6O78bMyzuaYas9mAAQkeZnGjkGRRnnFl9rLv72ISiHAIueqeVsIsiZ7dQi8l/MsE
iERwm9hIbntalqG0WfuJI0yo27VFIWXfPAa6tiLveMa4lJnaaQP8Hw5dkc36sWJZbjYZ6fFMH8GZ
7cuKy5hvo+3VpnUccjFWhB2LP14BhbVCzLafQ5ogAI4trgHrnD+E0gdI0j11vmmYpdpOA9AmYGlu
49R57U/D7cZIGbuYi/KPUaXSfbcLghpkqZfVXlql1eCFlj3Bvq3mObX6xTWZDuhZ3+doBRrTOnsO
tDAZ7BAWbo3RdHbAwnSyG3lddndyI8eUzpZ++kDmiIUGCChEM7kLBHRpejEDikc0ektiSCw1qdpL
tqWDADpV7KXxu6hoBA6f2w2P1FgpIR/b8cqh8oIhzmLqO/SW8MkP4wI3pJlhTVA0JMejv4Gzq567
dDyyfrhnWYXgaHeDtECOo3aTKTVI/YQFHLM32rJzTANj/NHkSry5Kff7SQcHz5f4zMqQ3TfoSmFZ
OuIHsOuAo+K5NumVTIExPlGVkQhN9JplYoCgSebNPOxwZpT+gfhtjnQSBZYA+NHLq2JuQ66xxDpq
Qxios86tdKgxeuqUvzypjvaxS/7WqAjMBpc5Nf/UHXCk6l87yobMTSmR31kZ+0HRRPmxOXJ3R/yE
kfw8me242KvwzKjsDCBKFtZMrkzBYkknBsx5OxbcaXuiElSlQzUiULLxUpwbNll7hIyaQvJYBdDy
be+PFME87HeepnVmUfQioCyDKR1WSvIdwqs5KhdvKoD0RaBk6Y+4nYfhU0iL9uE70zMEbTQlGiN4
XGVRPODJOn2iPEgS8NCrYNAbuuNnZIWp+Age3MiR5KwK3B5uaRVFXc5HNlJY7NSIWX7CfGC21cC6
JJy+l8Hf0cnWlTXWdF5VfeEU6OQ6izfxwiR0S3FMFUgRR1HADMST/W8+ORsZc5Hhs8F4hm0jL+uC
QbWQqGVKahIuzV5PFfzvSYkg9VRjUaXNXttxQyYkX2kbgrv0QyCensEQTvVoBWGFj5GA1V4/t81p
DGlaCCEpuw+7JJoBe4xROKWUpeK3OgS0ph5gAc9LUmtDoRS3cRM+veSU+9Pfh3EpCueogdyx7afu
fhy9rDeIK+awsp6ytjUB3/DtVLynOBaOaIrrO+LdYzi0bZ1VaJEtO0l/4M6CRZZdHlU6UjETDyUL
3uoszkmuHQVnHeTDznlMCT1/lETOex7NxXZuiEb+WjambGTPNdtjhvEr3u+IDmN62rVBp+zM535d
1SZT09G9JUwclqDqf50BuX/HvWLjhtjfjzV6w5G8eIBMUVbt8mESVU8y8/iAhPrkDZojIqqtyHYA
nh1siu2qmFi8pcfR9norSCzi76S8N/FGbDzWYlhQJ2+vKuoEmPILNp1Tci6oqTO9aii9F7e3QxYj
GYiN7hPcGHI2LLcCOzcUxr7jC087KodZOGsfrqjYueWD1jqap9sBTjLOwdXEXsHfZxFlpehd7YDz
xYhNfmRUxE73EzXUawO5Vsz77UYLLeOq3tbx4q8kvdiIV4RFW08f/Nt3ZeG2Rb/OqcjKjFI29Gz1
dWO09yi8TIFzScsQgM+w/EyVRzpUXPGjxgt3OjWB7sgA7cvZlBwN5g64+4RmA4q1yVAxb12DFVjl
BKbI4HhlK/qjb5Wmt5/MMpkhioou8XRf4BcMXnA3TgajzH6/tjLr7L9z6AA7grMCZaWGPniwmHQ9
cWnjdwj59mrnblg7xHnzO8+vTDedRkyRmKqumV3JWglmfjAQk9/F0UlDXrXxQNcv4QMHjqqbbcS/
r25/z43Pelo1DhXYPlALXATTIOOAZJzXEUo6TZRK3h8Vha/FbwL1n45Yg6NPxKzf2ZcEx7YbCcgY
FwTKzDeFgvQchRfRqm2zKAAJRH0WOaGaV/Ziq3nm1QvLaEAs+tl+VekIzMrNKlXUTGPB43ZaARiP
j+Ovwp2J2MW2w9prFJLvlOesoSjr0q2VLD04GZQBEP/1fw94/s3hSziEEWJxliPY1t1mApzrkUtW
Pi++v5UG5j4BXdTaN8q7hOgmBUyZ30k0Z1+lRmpCyzoTMMvWQRTbRLp+GvQuTdG5rbbuOCNMgoqh
gPcnHrucrhXKZM+oQjcU/ZQn6Q0e1tvEg1KmOsDHGCnNMbIdSz64P0UBv2/0azuJLw37Y9jdbcqQ
6eh+/0KXaBXYgB5g/ZAQ04a1jG8/dtxrQNYjnoLRVu0kjoPGGvBmnE4ixld/Lr4NW+z2G0JwZldS
9lhqPSQYF1lIT/V0b7q1vMkGTkz07X0y45uCIsmkujB8Hk1pypRUfIaMyAoV1v4T2vo8sHzevV9D
keqqQ9vk1isRNkhUGPdOL2EQ8WAau7jQ6yaPymBf/hU9pRRNO4SToErhqkMAOrG2Ua/G+EPwXkC2
gc7fm1KBPryHPiNG4bLsUR29w5yMa8ERwVLwwFpeEphHeq1WoZmt8SDHi1quZvpsDaB/dAdghI4X
v67i6y+wt3L0uCqT8uK8DJ3OxLd8fbOA8IBVMipKNbRrnYYxniud2G9BtBSuqyHPblaz+YKz86xw
jJGPrE+e5JPPqivFQy4UwFTC7z9+dUD477SwriwUDqvkQCOJuSEL9YL+ymO2te6dCNdtshUQtr4L
wZNyK2IG9Mhi13BEKMAqrw4X+Bl/ZXlMiZxTTwfr3S6I3YF9KvuORafl+JSOdxMlnhP5HdTyVcKI
nSTk3n2btNRzrJ708gCzI/3H8fqbRhHp79QiaTp1cUECJ8lxscEBKZFKWnXzf4oBdvH+W4iR93Uk
yCppkkmM+WqBMkZQ/G/428txBipoGM0MPIqVi4A3EvptlrSbXLs9JbNVPGHnAhimykdv6IoexGxs
GKojUkZo1g+o4/dwvsBs0xzvC5tqR6tfzDVIEafb1C7hXF3Ag8WnndHcUh0XCcyfdLzAEf8DgbPO
Rb184gDl7WSC6R4rXRbmxb/CJiaWWdu9JIZI6M8itoVONPXsma+m1TFnABm0n2l1Qb8e2Id9IilU
w3UG6GjgJ5ZhA04Dq57vzKJ5qPLetlXwF0kvEmo3vP4j4xeU3PWuFdpwCUd18qD/fid+9QGuxCoo
a8IXzkK1HbbDeGb5E9XzRtfQ0EPCcakjsIkRzte04cd3xXXMTaSYybmNr8CIBDutJKjEoBip1Xvm
RXql8cAkQstxzaq2wmrkYexqJqaezs7DvkSKwZfMJbPhQXeiIy0lPshLt+781yY/lsQIzZKb1Pc2
JgKL/coh+BHm3KnE3FuF80vaTLIWPDc+Ti+gNqwlcr6nHwGhG6SkD+iacs21YCYA7nmbUFmem/6V
SGVj4+kMnlT9B+m7/tIR5IMUcHt5aUVU6co1Dk3H9Ua8VKFJTEruHUiI005ATHu47W0KVPeGh3Ep
dCJ8YCAaKl1tby0XuS8ASv6Km446ek6TBG8fNTh8G2gv8joHxNo+N4sH4EUp78+OW8tWOSHQZmaM
JyqFj3vkYA15gANMuLYmF2BEq/H1bFcpW7bvNWoAoCfbWBKS8JFNwxSNyuhPMvVN0Wann1rLLbmY
mfdTLN2Qunj3ZGV3tR9ZHBTEgj0BNsWU/c02N8Oo4l+A96VZelNlswUSZWZGmA7/onz0RLLHZaw8
KksP0ZxQfPTpgAEQP9qjcWFk5kWYM0Gc0PWzZ2V2Mlvk7Yu7yFmcVS+laeIaTCkQBKZ7fSekyoIA
5kD3pXdS9rmYWWUafVDfmbKBqpSc3vKfDQIfFLwWNkZ03angIefytumv+EyPbC2OHoRWwPa+5O8q
Ng/ozHq7FR7O5phW/7QrI/itIYxN0paVKJJUohlHSQir1Xuzt9H3FX1CtmEGL81oFgazopK14QbC
ij9MuszYIvin2h+pg/uYqbwq3p+E0cgefmYEqMqBwGqXZJZnFYf/spd5fMaoqIHnvX8+m643EF0W
GxE+uXHpS6BPmb4sN1HxCmRJQDmVOOLqJpGLLLwauSvWDNWAH8rJ6iRzJkfTbtvvpdNza8mTvMyf
5V7szHNI8ybjzXOsx9hs78KflJUP8SmFls5QuzaGY/IpMB4BuHdJjznRGGOFRiuImHp6Zd5khKQL
my52R1v0Y3STNuCeA+i3XStKe+iVQ0XGSce/RB+Kfc5T715cCGAVNN21AmXEGSx8FER/x73CEdc1
MQiqj5s6pIlO80bB4L+S6eFY5nkzCW0CR+QFgYtq67wWQULWENE5lvCf7GxNRjHfUtQOLf/azLGS
+lMLUI6oRKeY0fLUWZTyohtP6g0LyYzTHHBOppHVLxszuw2B17LJE4Q5oyDNqDSzX9ikVMK8MHz2
8LJ64djqxPKJjmtKRDy9hLf645vWB3xnNRbaxI6KoZ427bOWX+WqErMChKVVbTYEb9litFD1WOzN
fDTd/tL/IErhE431U3SjnciSSipzosTJzrvypq+JqWxCbQYJf+kDqBZT4TVh/QFRuQLvOeaZkd3Y
c535aCIBrpxZ5eG5E58c0yNIM02spCtoSuN3QhYXCZLnYSOEV03yHInG3hn/SOJ3UVil4KvnEdCw
HXHes9KzpW7QeqQ0PhNcdxBSdyNxeFWBC5ZoJ9QshW8Whflxnx+WB+855q8dt/kg0pjzgzvU+uzn
WiHepRb7OawDU7Cc64jln4OO1sxxB0XPZ3xIgkZxn6apPCWic4aWnf8CUw5mScVAmt8IN/JXzrRP
uK8VGDwOnQs1iGVmw+Xu6csaO8CbChMy1PqA2rWUaAk+HZ9OKz97FGJwLMj7+9aD5lxb2IssZKnK
TtTqdQN7SUd4fjfvzA+YPwk1sRI24XODo0q7618jNKLw6W369I7ssMXz9ja0zk8qmmHjR/l0FhnQ
KT12gffZ0tv8ao6YydJOJGsRVryfWN+H1RfWa+cEblJ6SR4nDU+3CtevLGhE87F7OlkkcsqhpOxF
7zr2oHfXsuw0qKVV8gfdMxPklzHlyh1lZvZN4VU4esSsuqaR5oa22AkKh2ipe3uZjHCfk8trnjYx
8B9HuvOR45Aco01ne4nXKg9BN1LZtfq+9DCJf/SZzAzoWc/tN4utOOhurd9zXVM35BXXTW7azoMH
n+fhMq2bbxqDFltFHW95rb1ABFxjsaW92SF1FOCgsUhA60LZZBVX0RzOtBov/sRlo1sFDuU3MVS5
2UwKeLnxgu+I6cmZINvG28zMC9QC4UsuQcYbor+OWvfRZvzupP8kVfCQU2OdU81qzSQPmORZNpFL
Pva6yQ7iOgch1q/FtSVTfE0QXk5iIKpY0L66KdmJqbdh6nuEYNJSPblmX7p7ZgEjlFr6dPUynRNH
tAFHgTjh+b8tgXDzSbXRNoVcVPM+7weND6KsrgSx+0dKfaj2eCEEKiyNwxqCcIUi89MBCwYdEaoO
vl5Dt8CLlww3e3f2h5zirV3vi5NjiB020y28LoBiTqbdUI5OS+N1UvRuEsWnXOdA2m5bYt8FUJCz
fra0dH2QxBIzgCkmOBxwi029Vka+O6GjP+OaS1QwzUUgSispTXkivo9SgoLqIZPL/s3db1X+ZMI6
6idM8sdhHTW5EKoj9hV6Ip+4Koty/RjgHZaqBSrUPkD8Z8GuaMA23fU4T3gjanCNlNCPVW53VUk2
esj2EM5/dukKNt7kzjSM5EUrE+yzNUohF0rnxy1Qtb4S5L1nnoeYIrz/17H6bKf2d7oKrnnLhXdD
Nw3vkAhgEl0XMIHthKr2Ggk54kL1xryhh21N5gtr/lHkeaS0VjLB9EnFPMsCfy8lE+c36LJrlz/F
5BFzejQf01Bz4fQIysqr3kTOThLpB/+pf60lSvNcDr8ttQJdLjBFD9mfcQ25004nJZNL6qOf6xma
Te/ILpmktgxgJvQuzha+h4SXSCOrI5xrF5S8IBGvZegOrGfSn7T8U7FxNwr5qqbXqyi6MzT/M9yL
XLf41wpJM2a3zRJ1XAYMwym7GfkiYCfVOYsUK6OEULiYRuNOOTrsRuJFXO4RKmEqhMU38vRE/9R0
CfZ5vwMQZdjkcAotBRtHJ7u3EQ12sM/ku1QU5sALzrDEejyA8b1jhrwCgKZZqYLSy3b5aNJaEAgp
jrGvD9uD/do3h2tWYsfXG6I4rGvIsbKkYCaM2GIR3CjJHQZ7Xefzje4DgL8crocM7ynI3Wd+KqKX
SQl4hrFOfuw9huUnxdOC9UmID8A0LYc7G6q6PEVoMW0olrWuObhcfBl2rIIS9Sl8pz9PURNUe3sQ
yVPJ2JpQWCkO9Zbkx1tzvy/NCttTCSxDCO/GuVnjqcKDpxWbXnvkakFWTkrzXM+qLNybkVHtDL1S
rcTgldZAIavXdkuzMn2dnIpJH2XDIHGnBNpcJLnZlLUztZdsR0tCyoGTOC3O46fwbOOAagttuaE9
gmTJPqjrNFd/6pjkym/zFgKRRNGI90V4H73/c7A1uFJTvvdX/wAbB26/lFCsxBR+run0RlASnKnc
djN4+99ImPYLiAmhMxpvy5qqV5CXSC/DIRlz4wL1nHM/OnyIiRmxjhT7yM+knhwlIYrMXAFAleJg
SY0y1Z6PDLUrdySy38FI4q6qDQxm8QjIQuMqIlZuEMumO7Tz2agMl6c2YmApPpEEofd80CLUCziI
s+jtnD6KCGek21LO1WpXJ0Yg4s/TZRGHINNmhJBlK5IjQ0DYAcLow487pSL7weVMYQd55RiAggiX
xlIZiir4LvHQCDK/i8P6FIf5PXhc5qURI0WVFJmqTrRPd1VuCvZWU5j3ocnDm6MVdrE6Ibed8Swg
URsHQxbJGc1KJn86xRsK/m1qny3BiN0DhvqC467vZ+hqAaS/eogmoitChOJM2zqp8X9bCr6CLEkb
blG2Bq4PmKYzBzOgGZ8sBlp94Z8+9fsj5kQFPHnLCYHW8JSOp+EZ/uyuPkudTjjsKuLQZz3B0pDO
zDN6tUGOEGZd932hyoMOne6r8E41CbyCxF1N6k/HBorOlRvDbppmkCEJ2H/2ozPBVW67CN+yXKWB
64BHrAAL6NpEMACVbTbXaQK4hJ7T59xtMbU7QMhOHhAtPpIMS1kIXZMYo/ISuJqQqIKZ1NEw79YU
LQ573qBiPyCyCqo3JLS6gAKCfGC2shrfwaoW6UEImnu7DxSssVXeZHEIflfsReVdPVlJXLSZCWlE
X2tYAqq6Yq2uSdgya82xsN6C84T/EYLUn6egpusxwBPibBHuxzxXvxEL7Qvwy+rv16oWyj4zsu4w
q2annuCDf9Z6lqN0/e4KfoZwFR3AUXKieXbrQbemJ2/l7c32Hv28TIGCV4oIqtENJ97+z6LdHFQ3
J5lJCgDOeaaUW7Csvs/FHnn6Lj4jkgmjqwoOzJyIZiyrsx09jbDJRgCvIB/Oyup27MSsrzgnlB8J
dTo20zc2ESBLRnpptbKHtOEQCzQnEIsl4frsHXhCGcKGYEAQwOOlaBSX5ofp1oKD2kQbE2kBamkb
MmKitfBkHThL0IJwebFtomeMBR2EoQkj3H8F0XXhQxAEX3RTNTUlVWgAT/jta7uSD+8QfhLTH7yd
RHHncR+uYzZxREI5JlSHtDfgS1R5N+XqnVO9SzMkW6P4vPlPn6UlrLEgZ9c8o5ZFU2l/+mLHTuZp
kO0TZRv9UYYn3PeS2iobb8bdxVtnaaZNswhY7/9SdNaGVIdwuLVT5Hai7XKw6t0ifZuTeMdBtbi7
49/wayaeOuNeP3v2tlbhPsPdgsXec3SoL3GOfTuIlIr8lLvPQE6ehfdHhpeGdhHphxiWs2IMC2hS
7gGi9wlPPqeRqU7BUzOm3+fVKxlnI0Uqqeg/VmlOHUewR3rTm/iJKj1fi/TfgJHCLvgf2w+2X0DU
JZdagS2uUIpeK+j3ZjJwRQvW5opNLAlmHuPKHivN5+M4x1YzFowL2h8entL4EKMMEww3Mf8rxH/s
fHXZT8BBAoU9iOqBB4hyefbS3XFBH+ML50UsA0bir04pZWx/Bpx17aXFtxFeCNS2CepqGx8q7guA
TkyihsnrcK1P6sZaSKcfDXbwHzr2y2OHzxryOTe6LDk9kbRRs5yreOLEKEmPBtQZtmLh9v+dulHW
dPtcWx25xZLb8qrOPgJsKyH8GW0kOrn41IWpqYqqd9aA9HzwF7sqRV9yQMi1mXsQieMMrvjdXZYO
MTQHabi7mjZDPxAx2f1mPS7Mi12Y+P9F6HGwpgDkLYfkXTjPehMWn1wyx9RcqvkaY1YAr1YhJUna
yyMIBOK4oXtd07/v06slaTr7BV/GUmZc/aXf+XKdUiM79i2xFGUVwLLDXtRkjuoXEWGlcqhYsp5b
3VQsrhDKaaCd0mPOygkMn63DUHrmYWRSCRc9w72WBOppsyYmiuiddITdSyq29kS2IHN1iLYk38zD
5L4+NSQ+X8C5YSBCQok+05Z6deKUlcabagPDMZnGp4LL63vrzrnaJNavzv6d9vqTg6e26ZMhjbeM
KtoKRMhETX5bMDsX8h6y3OD5jNXc51gS18TvEObfVOSbASWez7ut5etszF4MEau5mW/8CFGCiKm6
6xXxREYcwMU5j24c7Yyr0iB6y+qVfgCEH4UlkBpl11ED034Vya+6Eupl6tY3F3D+tjo9aBMUxWvk
Aedzo5XoMdc0Yv88vSsnQlhz9UExtQDtYRzpYfC0vvnNZZanN77AkZIpDMz5hNJUGOcTukhXvzGb
7iV+KQgbjrdzzKtwhfoswFq+vLT5KWgpUjUU/rpIqKyO9G9S6X/4c67V2cofxaCEkA70L06SKaDh
aR87ugfycWTmX7IYnnqr82nUpbbEJaq7HyP5hcGGh57tnleivpO6aYTSd0oL/Ov1B9rwLlJwtd1w
3k34BeDflbAg6ECw+PdH8ElUYrvamJxr+VNm9RHynJK2vYLRCvmiBh3MchG1ODA3wJY7cD9k7m+t
HDuSWr1rawP4wFh0LJzFaftkZW1SyuSiLeJjnLzz/HI/Ewh4/A7f5G1w5+ZEriBvGEWu6oy+ZduT
pMjL3wzZXRcJHVyO+58/TosziXMA4xS20YTYcaMPi3l3/s9MFmWOlZwedJidGtD6FGVkaHc7S0j6
9qO3ihSs+OmFmYSCC0Ui2QJ4VjlGndxW7jK29e9XEeK7DyuGYWSHPKWxq+qddlIHMGuBZu0lWMMX
Rc42srBFkhyMWzDHvQ26Yf6MnLfp6/e72Y3g/cFdQ+Mkr2aYsnCtMKxnH5php2xf22Q41r5900qP
K1oXsGE08Qhb7cs8VB0D69x+6aAJDAe0r664JXiikuoDYIeEcVNGvhH5edVfWemNFJlyk+iu9WGj
rpPKhZLoinNebJ4Nj4L8AKjZJ4JlHcz8lM3s+V8+84EwAZ5zTuMfR+0ZLG4j8We77wGyDIGt4igq
LOLkAmLO5G63hy/DGgmQtF8txzQfM1ZzS7sZ9HngNCNflm9N8Jdaxq3pBHzFEtkv2UTWiI4UPvxH
MBI8TddjYRfk/P4IqslMqtPbpRVVQA5Hh8JwcX3jx+NJzpJdiV/1vZ4cjZT8XvkQg8ydCiGDFLDQ
F8grr0+GCMYYEq0eiae5zBGqf2M4RBBB/+hVLRP1ZIc+PW6KdirC7GoumhEZoNKakN8UlOWiQdKW
PRAfqkyOU+BfYCoRIt13j+VjMuPwto+vHQ8GoQ6qNIZlS+kpmN221hmzkTaAerYsRLyFzO9B4ycl
nN0KOx3aFEOWeWzxL/hRmysrO1bqmOGqSnP8jYEYA0C+XLVJrmxuoiqGnE22J2/yCAoiSfCNZAK3
X/ifCv1l2bGfIjkkzNy41oyOH2sz6rOzJlzZT3l09EcfQuTORyeoqTEc+27njtcxthIwc00cFu0x
lHiuQVT0aMyZXgCazGes+ocmR7L0oFPJPWaNrcNxjXYIQ2zIVbdgscYnNkRxuUXLFlnRP22w/QLR
+osjLECSLnb9a1k6ax0JN7nI/LwETFkj1uiWnwxAr9R7G/OwuAgFJM/44yF4ien3WJgeAGNx37RV
0Ydk9N+K0DVkiI+GfPaxO/3CwLBCrGtu63kimjyRS2tjv/5Qg0h4gs1S2q+XXD7JrNHzX5ojg56Q
h8tJA2kVlidBQQt20NLPdYUufHoEGE88tUqfEIeqZ7Ubsvdxo6mWrq6MEVYK8sKpclp0Y/UPS8/b
duSQhnx1lsAfX5Ml0lsLXh3psMf9vHTEPVlVqJgIE9INJ5QUhMjjt7atDwiGdcBzw6acQxdU16zy
ra5902q/VPm+7pNe1iglg2gsfFqzUxJ/4uPokrp0HpYsiGcmA88shqQp3Rqw2BEkfoW6yXcD6lQl
fYzfG4nwTY51I9Cc4klHs3sH/eMXy5InxbhLoBg4AcPtMjZ+EuSytz6dCJhQ/Wbd3uVSbpciOoEN
XihFM/bUIJqkOC3QWM2KEJHWVeUeHmscafXKdWkEZxc4jFw/2sUfHB6zs5iKjbi16W3HMZ/7oJl3
xT+44S+Vb6Lwm7BBsl6Uw/hqYETm5xqL1kFmJPazrRsv0MMGQy9lBE/U1mKEAk2Ezw5pLuYhWRY7
nURAFciVONFjxD6XAvh9qAvRy2DnX9o7KEfK15+oDdaBKdpYC273eSQoun6sINEDdK5M/b/6gAwJ
F2ruwEd7b+S8q1/P2VreIEvGyLI5BiqR7lyMlV3DnhngwVHSas0/rog4h73bx20XqSrWUOllX6gc
7aMjb2DleujZs11XwwTwk1rrBOdUlfVrPnrL0ZBJaZl0KiUxLAIkYRcbsjt5Y3rFUxOgKadiHhDI
R/jYhQgZJU0l6spog49s5nIFPHXMQb/F7Q32S7Aa0A5ufKS1DAb6xLE7ODcsckANh6U7Ei9fzOna
CDr1WZ+pxQ+AK4Fm66iQrDlWpm5d7zmTcxBFCYxpa+dSpttRdKCCztU7Dj6RHX/aBFKvR7qpUO8V
Acr/1vlXs1nRT5yopj//SwxQzNr7KATjdP/G1jnDw/CoukTGZSIBH7Ey3tIsn3UZZ5cTteAVYmtR
RCR/KepePwr9wotvxSNGeTNrQajFHv+MiB79kvMxtiS7XhdlIAM9F1ysdJISoAm8Tmoe401gSXj6
/FyxghVVBiDd5swUqWsznbwI81qUQklKR95IAEf76L/EXsWR0uNgHi+DacG1A3rBlJm7OFWxdBM9
h9wEqUbt1gKkH/4Gqm00WCBMFEtq8nflCYlhT0iCumfMegLDDHEKlb/m3b2FOpRB1ZmRY8vn1xSx
+OjBaQFwKkPU768VhXZt0gL7mOeASGA5vrQTftVGnWe/gJTJraY//Z2ROmh/RnZOcJp2AQ+aTFCx
1ZxkwHtkXB3p/OeeZymPiwjpgez+pIm/NZdg5VGaZi108BGBKJ0SPKrcut3JFq0lfyU+aOHUdUre
iiDPLGQtWAgsXKpMNOvcuXeD1W63VmbTZJa3Uq4gl4J7KzbaErgc9/Jg9gfgnAR9MVnj12MO3xTa
mzv+bCsDD3z8wNGLVFhCaAxC6p8Kuh1P6dpV0vUMjEDHCyMbA98Yj8mPHIjb0JVF77yt108ZpvLK
6uF2AUC8aILdTCD83we1OU/RNwrWIuxg41V6SW+giwjZaNzJkl8hszv06JDvnV2Y2f+iohkDvFgR
OppC6QjbymafM6kA4JFWYpK7CbXgkBGS5N02Xk2UwP4V8PKKh+idyVOnOuYD9usQ1AU0ajtwxmiL
1OTU3Sqx/yasO/86ousihd43YKtT2qpqrqBzrZZ7SLji56mVfEElvXZHx0//bvMHa7IMS5jP3OmZ
KPpXb7k84N9XBrH5HX0h4jrgHAXaSKMnsSB4QSInCuXcZVVypMgrO0AXbV1m/hNFfVe8yuZps7lE
iPgc9XbaM+UrU3Xy5DDa+AHM+gqJIpo9IF7H10wiKKegHNOjd1xiiHtvyD1QZR8PCc7lShICYRCr
S/1fDm3rDML+QYbJ/QCFvJ1Cj6JK8Wn07U/jisF9X0Dnac4pJ+c7bv9ZEbg6DnUOZLxIU9hY9zKk
RwJy7dVfsafl3k2t8hMEaszUzlACdPAXQ3jhFnA6ssct5czEUuok9jGi0IOGcgm3vqfBlnWy7M/0
VBZw3wy4rILiF8w2OlPY7aWaLIayXJbV0NsrZP3+fDuZWTL5S3sm5tQb8JmrzDYnJk9Lsq7HgGSF
sTMXvPH94R/Cr3IvNUQDsyn2of0G3NVfQ71a34Tdhq/NR+VxFr9bdhHxaCB4OL1lfirnUhuG8HoJ
hsEwjcWZ4NWI+znCj4ny/hqLls5dN63CPtd4OkYKacrlDzJeq+ndAgSvirk2GOQ8ABbkEzRim1X8
wE/PvdCUlf6Wnx/enNiYDcD0337pyxHOloSjOw0P7bkNwo3wiIAInefn2WkmNU+SkIULhnUckTxv
izty5ngpJ3Y9WGmRfWE7NVERL9GbrOO6CcRM5KDZzHHIVZm7KQHCwlFk/syGhq+fdVe1QP8s1ohA
TbuXYSMxWhYZ0IwlNEqAOcDm1VPoRIcyZ/tS+ghJxIiSwtoqTa/7u5FVG+9L8qu7ZkLblHf4N7UU
uEHjR/iQAsY565m9aJrscPQ+AMal3LBIJ28eOY5wo2PcdtewK3qjjtL3jaLEfh4/+2EW+h2sq5IB
aQRkdzidwIQNsayUq1Uai7081bX3GBMO7HIXIv0Ax7T2WjNNl8ugUre0FXKNQad0jihR8OHT3xFg
L0ElkAacEC4LgYtj0XBg4g/ztzf+7jZpjaLGaqfWj816E+czc+U8IPimxoUYq9jTevUGvt3hWr19
IPfZz8TnvK7KjlZk+KEUO5ct1lkfQ12j32+cwPQG5Qpm7aSDReOnoYp9IhCUKY7TmNFqwX4DPL03
eKOEvMdLNULy848dOW8fywjogQLG1kagUzQOgm2HYZVP1UCv/5GoFk+xmawHnRpqOiVdIeDDwYJ6
j2MVhQDptAAnVZwXyBolufdFpaNz1O3sB7j0H8qI1j9dKfZJCraIYZv/u9jlwAJTjqbSLHD1pNQs
7dw0PBfe7fef059w/1jjg3UlXiHihkYl6jK1u8Kg4PtoBbmSY7AATQuwT2ZeCVVnlfSzm3aIV1ti
lCZOrnrQX/zVEKx7QN59Ta9GEJFz2BaZRYXyLSrPZ+55gQiIUW9MTZBB94JVxgmSSuJ8egNt3Jmp
9MgpZACGFg2XP9cNDGdKtvd3VieF3iarTVb/u/pQmRQKUJ+ar7m5uz/lmDSkgz5NhtAIAvFT0CDS
vzsAmX0jURS5Ckpi+oS6+diIvfL7IvWnGmLUyuxfI67gpQ50MhQwr/daKcAh/5udJXuE6y+ZwwW4
WOnir095hMfpfCQJTerDRNeRKy1XCZd0O38GhS23QKVgD4HYTK72o1O1lWR72wBCwBC71pwAFrtw
O6R/SSYXRw5RufYdRXv8P33qpr7f5ujx+MCLrxvqaDnxEsvvd60iauba5tND282nJa4htv3OqabE
nbTOwUJeL7Mf+LmXSYfGDvHSCa99trWvZUuIcXXKy38P45BmYwtAaArLhkwNGNURG1C5b6z/Tvis
j2UHTfTf2Ze12N14JPlb2lg3k3GSXcf2IjraeR2b0cPJkx9ctaHZOy7mAPAIwYr5EIk6r0KaALsM
kxvjW5MiRcnQ3ZDlEWBSmyWpKY7g+4XCVYK4NXdk+sZeivaBweXsXUpqGd91ltDlC+TzuVDf9kg5
bbYMJf4kSJioyFJ6MST9VcNPt182oI9TC7xhIjaXlVmPFDEtlgE8Pd/BpGBumjsofeH1au+eygHL
2+VrEP0hkqIk0xwMxV0eOrypd39EIsGNycMqOwkRoaiEUVWN2Cg0X72w4MLXJ6JYjDo+00XTslkL
YFNn5CXjkcSRM761+B5fr0WY3Bjk+EISk6g2Pt3mJBDNMwz7Stq1SUOQ8bCka2oztZmsC9vraLsJ
9moHZs1zGtF3P4EY2q6I+0JfVpS/Lf3Tq80v2DTPNpD3I8pC6K/ivUHC27O2VJknXFLplZFaj7ju
rYf4oCnfUWfPTUg11gDuG8n/8iLwFaNJeHfKdn1a0vjfrl/+SKYgRcf2umW+7lbasJzj+zzDlmBY
Ora5uTx12t9FoWIwydiE2fVrQdaxJB0qHWs298Xq0vQQpO6H/qgbIimvkBMgK+KjbDK1EBoqw+zu
cI0Qr7az6FUc0S7tkgZ/rCfxLhEPPqvIsOqf5ZxFAYq0Wt2wk0WkQNqGJQhsY7x99oEzCQDRW3Ic
5ncsq8sfeyJBlJGAhYbeXYN7V8W3zGDhvp5EP+d0fybj/LPZezbFVksQfrk3DzpSo+52xoNc9mgW
MvLWR0XnZsw/oUZGou/y9oNJ1kLbFXtzhtmTquEMd+I8pKBJp95pSw+HCQ4PALaWD3Uta24KBPli
T0RztXtbyWYQlEEV/sSJkSw+7RdOf+htr1wwuHkIgLtN9Yho2f82PHt5N+AGRGepzovR5lK/ftoR
I2/m51XGJRATCY4tdlN1a1qcjjyQqbesHRh2vRjlELubmyQRLUslnW5Z56Sgw85OLI3L+T6EsteR
4KQpbSi2P3yhTO6NUXoLneUZL4Paz9QuT5mcXG/3qKLkJwb0uZLGltMcreL50u1yhXTj1642U4f5
u5mZvLTBHQcystW7SHXQfM8dSL5QyWyLswfe0FTtBHq0bRshICVcp64xr0BLfFJoZjKyepyV4tM2
NLfJPjSBz/paW2FL80W12XPkFWaHJeHYyO5LG6FANXtPDI7KPaH7KMkcUg+0wyRuNnVPzE6F29/n
JXG3oCL7WXbjdsxXnDMnZhxhWf0mEt66ogdXiisfuHNci+PgfAbAeY0VYeYRYbbNU1cGRGAeTnOV
jypBmxnAcmPWc4hV43otDTha+xrtSUdUmG/RcRkP/v56leokDlwG1Y7XEgf+IfCVez/CosilY7z8
bbGg5w8aqWymRpq7XCHgKSibqKDhTGTui56qdS8lGFQ+7loEPp0sGWWz7KK55sqIzES5tpvkR4jy
QPqgwqJg0difdSat3Ih2OcI8dkEXDMd5yTPq++NIZCXMGKffNVcCQGjxgUndHdOHepQT1jAjkmHx
dk6oU/1XH4j4uhgNbb6nxyTkIO8cc8AfCtk93dlfCBw0rgzvKRsYWb209TvRuCfbaD1ALA2ZP1VY
8hTDnvZrQd64SC2KLVxlqGnAk+7sudfQMDp5+xMt9a0ztfscLEC9U8VUaTcS20djDAAQANRcXpV3
rat/uQu+XHDKf9hPp2FN11DM5vnGvaHUm+RB4Dldp6/SHYWBjRSSIsannEGraJllfibVwp+jWQNS
UxST7eCukEkoRLJXOQYVoixDKLInkHlm3jFWatOMvc0TXB5xUukHg8fh6iegVMrgXZP2wnhv/r9U
EusWR/GlM3UdAL3yvi48RHPV8QQEU5IWZW+xcRNMDIRIOQsT9ttEFThJfeBG1UqigrPAUzU2Sy29
nthQuJSkh/k4Z0oMrR/dYFi8LcjYny4ZUNzMEpb1n6n3Tyw5enCMAFsYGJH5ZA5ZQXXijsK5id5n
hcm7hDK5ELPprXk4QcuAJfIFjogEU6kK+Ln+QTMgMLpZbAz8Uk7JVLmMePRrqo44/y7WskB1E/RS
KrtMb8L2+wRqXfCZNVbIOO5BXJJdY+oQHcFajrA2TNv8AbL4yhKyfX8Bb0gTHyrYyvFuDjkhthtN
cfQLSU0LkVWRpMVSAWVCSuzxB+6mxTIGpC/udSIOHcvf990j2oUAgBPx4HmNPsDaWnAaw+W46KLW
mnMVSnJYUceKeCZjUnQdzoUrE63pAscVqc5VcVJba2jGRx4INSR7ZrkMErf1U2hj81VMOudAR3GE
BM512IwtT6x9Tk+CnFhJpux8iUPedVRml3L23BDWOWWcldrdBj++imD7HUnF6iZSLA3KPxbBiQsA
pZZL4FJ3OfjG8sqKQdt1CIXRZojEk4ru+YPvssVXR3GCrLNk3SK3CelcHNRowYtU3szfqKyiMyoA
KCO2bdAFSSHSb5Ie9FNvF3oEusSI2BL7D/QzgGWiUZA4/yW95jiXGhODMQ6pPA0EhalyzXvDWVYo
ybCZ6BQ99X98sGNvvCRTnz9LrlREbBKJcKy/OfoLsA6OX7XJgfr99vJhb8nihCqO5pTBMO9smeIv
jfsjqnq6WjDWWF6pfjtmUc1nIa29jWF8Bio7olMU6yQdj4UoJNGdF2RXrmPT7M4B8xb9XKIjDk8r
z7t1ZK1mt2/yjtkhOq1HKH4GfgoRwr4/cV/AvREN16R6qqDb4iKAf9+6wMQtZ6q9rEKu+ZbPJp1B
+qm4lP9H7R/2jv59T8Es+ldltssHyZ/JGUYYe9IcnMAlqQJkR+bDUIrFe+DM24THey1Lv9KBKbMn
GRVJWWKyIf/PhOFUIOlB96TnmfnsGkgvBj1WW8RWfyPy6Gr25epOL3AsaLNFMzbl7l0hZA1r/RzG
VaUKG5JR7KoxlV7TLTpG0HW3+8C3rlbVWQKl7W4C0lZRoAAMQP9keSwgFBj5GqwBGksVxsxsttUD
1STWd48+zaYy0XsE0av7S35JVaVHpSam2BDA15oQtM7HHjCgk2IiZeaQB6XxF5PK2kfFwFNqmBZa
GpORT0xxKFH98IIbAZZrD55dprpQfwy4S90PjnxfHa2W1ANom5uTNgZtH3gkW0UQ8WiHXTbAxnVt
Ok4+VrH1hWyucesOsWkLNxcLLW+jPHtF/qLGeP7irRggzINDf3f8e4sgObV2vWhJQ3OLVDyALeZu
WYf4PzZXzyMGpcLX4ELSAhS23ouzBinsK164CFYcsqthiDFldbvBBUU2y4S6HWsLg0CDNU474EZE
pN9N0LjZ+oLDIJEJzcDqL7R4K1QvPzkf9RGzK168UIF7MSwZuqId9Og501rBL6pOc2xqRVZevY9U
dFc2ty0wMbag9mqfM2sgvS6kO6w5pn+myajQR+Vq43RL5qHFZtHvbkDEDHRtEiVrN5xK8Ia54rmg
yNQb/Wr7URtgMpoV0k9JnB6Oq6APfbMnOILOHdtnEV6agRCDcygj3FS5QU6JdlOQGew+pbiv6IWN
uRJ+aRUqlieqcbaZuxat7xu+sp8xjsI+WgIRxS515d5Z4zzUyAIhZ/VavcxEywc7kRKlrLWElwo0
8d3hSwJJkNhIkPIlSti3X8GAsMd608N2vlmlH1WXeUgBzJjhJ6Z9ZaE+po3uke1rmh0Fi2blL/Q+
fGCFpyIPBAiTsvwQhe4ycHoH22tYmhoyRkIV2DmnWpzS1pomZJs/aguV6F5UoN14Y+Nimuzdr8vg
l99aRV3yNdkY5ejs2kcir0ZdD3k7b0mFDY0zwCq4NjPPtDXU0fEI8/q6S0AotKzmYjGwUF1Y+vl+
+w/3oEcR5hpHosT08b34SbGFu88OE5PhKWAa+Jf67rUdxwORqbMfZZE8wvqAJzvWjhTIh3ys0LdG
vmSG0FUYBENUBVcb2jzjmBIXJ6oDft4pN5vDrZU4ySRoriz2PUG8GCECXfix3tBjfsSxZOiv11ze
YssrHJNgSPOYAZn670nC4ONBCEYe7ZBBhihaepw3IeDNh4lNO+rUP/DExpA61nBluiw/CUGhoblL
vuBEQOZwxIBSpSNRBinffoyHgetWphB11ZiAnPnakaN2nokV/tfYw5OSv65vBjUwiqgZeyNokmC7
yoFB/iQrp4sls8wVbewIYW+oF1h7yqArbVIbo1RzV7BbF+mTGPsZQS+QY167FB7cEBUHMmgsNlbt
KPIDqtLRt4KXmjJcOMDBFpDLI/JUTWnC3s1T2PXEAkn8DNjroI3nf2pvbg6wA7T9QafB5dHjOz+g
Fn0ILkrJAlrweJBmJAPR0AMM3aYLeztoNutOqzIYp3v70XjqFU+1qbyHEYiaIg54XUMUvmtIf4jc
1XXf+NBJLn7Z75jI+bJ9J0RbX2B2fh9iQwePgN7NHig/iMzvpwzrqlMnIJfgw3Y1TTGWNNo9Y0/m
NxX24c07ERAo5Sx5hU7nNZ1uU9lEYb1/3gyF8PWMYKbfRM8eLySoPXcGK38xHnaP0ZndLfiS/qLc
xvf3vCBxPC91Ce8pM0N2aQW+/VhgzJcp+g3EZn1G5GXXRR0pK8sZ3wNPxJw7tW0GIXUrM4Xg3qn2
7gI31VRoiV4eswgPv5c4QrIS+QpXTMWgHKkrupSMPKtkBvszpCo4i5N/Bdf9TVIQIAvajGy9PPDJ
K/OqkpYl+H49DJHpVNaLMOeDMPoWam18Ad10if/aFcAyhWQ1PwnhrWX1B9EzzCPwjVm89jtR1hD3
LyMpWXwtVB6wHA50EL6/VSRqZDHfLlPtNcYHLLxxSEoRhoxQn8KkiO2HB0FHmAszFCbCsyct0AOp
oUYy+rxcAbpuBrV3OrkZhfnH1AqOYg4BWgVoUO2JjcMnPNPltGZ/xlgoCPszkYGxn+RLM5HOatnR
jLPt58Us45/HMeT1C92u9nDF6PEg99a261T57YuD6KgevftKqDgc9+Ep5/AWyu0YqhjMiPqttFVj
9rGX6Cstn92SiKLwFKxrI1BvLJJRjr0GMf4eX8r5KF89fwfpyzhBn6cnubkTiNj7Vy1/fpMDMB9w
MgUhpnHOCrw9ZDhVtkb4sJHRdw1dzp4FOD/+696oGlhX8b7xBNuT2bbq4cf8yhYvphyM0MTqC5va
BjtyvW0oooEKTDdNIqUIqvbjoZMI9FSyTRY/doGANRV6kVvxnUhBBhsm1isXA6SZ9c5yFi4cjamC
ZwzI4b+FmlSD8EkdaVgR8mborRG4z9Pa5PKAEzaYwIAn5d1n9oADvq5I76GOHNse1HWbzjn+e8AM
atjdxd/FIVMpoccPss+X0hnMrvIj6SrIQ9lio2wGGraWsyRBUcMhEI/w53/xTqmMc6nyX58NeP7y
eSO1kPsE3yGMouj3dlLufDvU7h/jAuLBBxKXo/JDBSNVOo3NFHjNzD+gRqkkCrhxgQNE8sTX5S5F
2xL7FMEWhBlgAsfxALX36lMRgqyHOyq43QmAooi/bdUkHT+53JuoAEjDyOwHGBPLIMMqPewNxS1c
5nZa6Fw/VGFRczdRLMYUZK6L20LmebM33lh3+mVhYUTKQoa+wO3D9inl8r3rFJ2U9B2S/sqLSjRw
LBzrJt4l5j8TJlV1WEQ9WL8Ciz/FYJx47C1E8gFMUEq+KS+TKnmERntVoHb1SQuIMaD6vAhalSXn
GbyRhBTtvoIOMsNAK+uXzkSPjQ3F5qjggY300pIJjQOng3o+vZU/eguj3D+0zuVOHdHvlkXNRhf9
wxOdL+Qcp3p1MXl9/1C2FHNxHhEstE+O+0KnlE1B1GlW/T4/VG9ZQvwLILMbYxNsKfcx7aa5ObN4
vauMvBfRr+dmXntyeyiB5UJ01ssmY2tfDlbNrk+7mGW/7lYsO34/ekpjkZbBcbidVSgl944+9ryE
1YPUl2TMpT+qu8uZRoA+g0EsDmv8haYBNcpeSx4F3z3W5h9R7xsFztZfliNUPjeRzgLZq3Q0R3kS
SdIeuTVXjvPZ+ZiROa+eVYVoJU0Q/RUnR5HahsXbTiZKhuzcLyOXwcC+dRHFypSBFgL2BIxiiclJ
1qZuxNEdVp2DUGuU/EW26L45yZJUIpg8gPMorbLQvSPiQuaNZxwpaFRh4jUc+K/GeRBiu7E0XFj5
kb7pz3cWzsbJIacsGFvZEk7iWI5OJEobyupEaqaXAKcSMrAj2p+7cH2DlqWlNK2DSO6rwwxnXvyF
GYm3grkuDYFWU9Fr4yfdvKb1SgU40nQxypXSxRDEILz0dBcVA43Ok0qBGDXcYkoQkjqIAcvOekL+
ZD1EbaLogail2ZwdgjetswmNKUUxWTpjGu0s3VdpfqHj1UKW7qvaOZfHricMqCfSsW4BJLa5CYkH
CepwJsm5/8MGH1lshMzxQUEmUc/aApVKtY6sQDJfIVVxvdz4ZbaUyTsucrEnh4XBm1qb89bx4y0w
Sj9TiC27faeZIKOwjwF5aVvSAWw/9YvADA5/02wCHkYpHQCFboot6Ug+PaxV/keHqSvkmXB3W6no
OPKQWM48WfibNmE8rPpuQvoCE8Yxo73ye/W78wOG1Gv4yHHTEYkd7Ff53DGi/jjvb01Uarwg2r9O
vli1/ooRoDc4urwASQIOtSDNgRlQFjH0VAsgfTe1PSEwPSWCH8lI/VAXpkfG9EoJAJvAPB1WaII+
ESesQNxZOnjRLlG1P4HfiZEDu2pJ5v8H0JWy2LWyega95IZjU8dDTCnL0TFvh3Tmxwk6ooJbl4C0
TMpvb8BHYWXbJG/y22wzGs4/7Cd+N48t8z9h/gLJEdRi33G2eD7p4psH16Gk6kBi8Dfrg/331F7i
4x1h0ZNNUnset69omjXwqsHE0b5OCdizaRu87BEKWA+uEx3JoX2I9T+bgimHfExrscSeSWLC5PmN
Qve3eAwot8lroy6on8qs3vXXsYYcMGak9cPwYzctd36w+jOBU2JhKpxbUt9nizEq3R1bxe+xou6J
ByHcqjaQDrCBxdgzYt9BArXXW3PIKlCzCPQDqbq1u2h42jhkNOBT5YY0MtzBCJN5Eau7kRlUOWRr
ANQIfJhuHQaRs3yr/QahlgubY3wD1GqFF7Tph61HeTL4tdtVzhuD6PQZ0WRHpiiomTtMIm1IgdGZ
yE3+M675wxhUaNpJoKskJt8pJtzSvMulWp6FAc6VALv+mUmeyDusuknwgKy1l+XBxRzvvnb6bPPA
M/3JaZXT4w4KdUvbZsohwHSs4ZxTrQ7JIt7LVU72qhtk8CkVHF0hX3AKGrXJ+nUPqmVr3MvpUFAa
JEOCihrR6JFSBX5hJAIgPPltNnHrM8anVzB9kr9OsSUiZN0QDf8uyHhyaai/hI6yar0POUxtfObK
Xa7KmFG7GN5zD5FcPCQ6JpnfI05q5WsvU3hzTTfbu3AIiclEyVtVL6ImAIkHmx1+9GFCpwG6kIXU
o30hr0pPXwkzZmsEbPub+/Zrj7A4a5+RMWUEhPE13H601KGWTwthNAtW+61FPKzsq5L3wHpcH26t
1i+wiCzmP1Nedc7kiXJ61vPwMd6filKfDREHS9zv3cEfty/5mFuVVbGkjRzyyDBpEKBfXwXPGrvQ
t0uktkaz7UPkMdXlk+b9MfuHtcpBRLVagbq8Y0XOs3BsxFlrWCePe6RtMDr4U6CdEBc1GHDA/b7Z
tSHxMz44CPyHQsLduhdeCkQktV/d73yNTT6NUZPLVeO9Ityw9Tcu4pY5xh+Vxz6PB/kF2u3gXuvR
Kpl6OP9drT8wTVnA2fEMBSO1N+ojWL13LCi9HyaDPyW7Wd+iF/DdsjHn3OK9oIEJY/pmjnUJYvFW
37bF1SBVSx8qUkAXg2XU8xkIQjE7VhZMla+wP+32LtDEGEyWkO2ic8E1IGdL5UCcoj15IsXAm7R5
rxn+ulUirfCmX/ukcgA96FFtYA1cVv0UNj38Yfk7BeFY7m25IhOKE5sS4pDWQFas7yTYN7jRMlmP
jouchOJxN0OCq5NMlzwmlUkohf/5ntaxUKS1k7ODvD7vZZzzr56ohVjw/6D1sQUvHpjyxaFw1IPO
BRGBHoO3AOJ3ukh+2biovxKyr5rnuIRsd/sCmyXapQwH4Vg28Q/33Hb65hOg66M6jM3cHE+xa+Xu
EK6/8M8Z4GvAbAG1sQ8+genrE+138u1mN90NaipMlXfXeMT2Ss9YLvyetBZfsj+fHq95z3jsFA4w
kFkGKaKB6TTY1VnHD0HSc3y7CGLTClnQEGJye1SmxfuAAkVG67/VZA1zXiPvs7GrxsEaHqBPdez3
aE+S+UWrlNtDSWt7bI4vgilYmtwRkyo1zGaNVuA+mfaANOhJWDKDHexS9bZz+O7cx7I8qJEStSoZ
2KINzEAvpqMt69/VgdDoYOCumsnHHjkbIBINI4mJ2jHxfp98YdG0toaultlX2th4PGxmouKL8UU/
TER3djG6xfEn/6C270pSDenUXsyO6NhrU0LxnKj/ew6yTjVnVggtfc9xoMkogaqmJ3HkyklapXAU
7XUJlj+awgCp7rkf1o6U9OyFAjrXE5CQ/IjYUaSw+pEfoJYbZWa3LkD5laJoaiPEpIzdcix7Lavw
GVtouKOjJ/5H9zH4EACq0vSiBEReb8WPrFEfaYi7ZAtIKaGPV2zf2hBVJ/v2An/6o0m/GbU7hRaN
ffm/Oc6l8KoZxCkJ6qgU61I65O1c0OD2uBBGYAvizR2frHRnVJ0aMCUBZqC5nljIaLUhvZo9e75b
yLpoAniVkWSA23fEOuhGpMBzgLgzXttcF/viiG9Febxqs6mLcya9z2yfQIusBtCpTmZnsTfVc0ge
HPzQ/WOaYsgb6P/hu/hqFBDhKNj+l58KBfApcuOCZwInNAR0pxQkSzxGTaj0LmElyUQa+94D3jMd
aP1ZNG++GxmUXWHaCRQ1pyPB1ZNRTh3KbEAWmT/fFq2bF1CE7hv4+g7Vak2yxyLa9b4cONbggzQA
SF2hPtZCmVdS/G2+8VkAtv+FB0jh/P0ALGkvsrwkihAB+RSUlZwMkmEoTKwem1bC4AfnYPAFcKld
7N4/GG3bJpgEGLjXNIsdTYOMfA6ve7NmVhHRP5tJO1XVoOr8qvsP84kl5/97el7j7zKSANQZWuXh
j3l0LXHwybNdVuY8a0fGlLz6/FBKFAgN3VXTkqXwSxqFSgF4sWj83LFT3IZCYpZ+B2tHMm3Y/OEC
E7MReRhgIQY90IMJCC+WA/pSIt6RVuJhNvBwVg0BV2IbBO7o4OWSdMo9R8ZncwBPZHOaEJVQ6fvO
GZaOFQtqhdsYdeeMTeu1Jw1lTaEn6q4mMK3exgaLsMsQPWyL7h+790M1tkyOQwUOD6jTRVekJQdR
BxcBiKeUw7nmJgIli0il4XMsYJwGEKHY2pylL2qU+C7x9l5jaFHpRBV4DhQVWYB9vTOj1f6qBHtM
umDbegWEYVzMKZXgzIs7T9+yYHq9oscBvMjk8RkbTBJfDkfIjgi6WYYRiTfGEo3KazftS7hSjl5o
QGsU9YzcD+J5DXCL32NAIZnUQXraca5eJfgJzOCD6mgBMUkAE4bHa7GyaJBExiYbyGTXoy+pWbPQ
1pR6RPzYgTGX95SA1BTzYuHSwLWuiReg6ZirtsSqJU8v2NqLLfTA/FVeb+MGyRMP6O8LGwFJFrlJ
5oI/pBUCTWFKZYPJnwCrz01ro4B41Tj0F3dLGpToFdHj1/13xj84HCgEjjCUy8xEpiv2MJC0BVJy
8YYPUnXqUwPRWvTV83CSq7eTG+Zi5D4LgzPV4GoVHc4f/b5rkK0eJtQ8OmgboQD3zyIPrjVME4s6
e4XSCj6ZIJReJ6sB38fuXuYfD3Cd3RMmYyQ3H2hiQhOedvvqLW3R8MnCoGS8n3kw+P4Cy7faHkiI
aH2H3V0r4YQxOlZxfogaM3kEUblHbBv3oyr8GbRs0wH4x32+FUu9Lq+7CCMEzsyE1xZcmrXvA7Qm
5YTGw4xUh3K9gQ+iS3RpSC+d/K2aWiyfWwshNAYGAxxF5pcbcY8017iweOjl0R81VC4bIxbz6BKa
MG09hdYpW8tGMcIxaii2Go6JbDEetgExYp3aINIdEs+CnHqax+KIiYiP4TLH46YOcyer9h43b2lG
RbQyk+/kC9jwES4ADTweg5LmraNjZE1ktPw9w79puOmQ1At/uCnXvYp83s7xW1IuHFkqLVzyXLoO
aFKKKMdGTV3QlIOmfvgK1kjwsB8Zqagto1py6AmcDg6pbw6F/rhzqu/DbizTJz6ydTRG/zdEmO39
sioDdvYV5fC1H0izeFFQNsMzq+XKf+hA9i7Z+madqA+7olg6t80UXDrkHmaexrGwBUL16G0sNox3
t5jtxbjHo+f2uKOrfpBI2zW/ET59KFv23fkbxVO+5AgW7isZczE78uTY/yZJCxCwp2ZiQS2/jmgI
ZTQwpdi9TWl0t8icTGOQfSaj1EbX2jHyw78Xw+4bIZs80EvLc1+QpTJtAAOp4kTQ/OTa8E7rPFrU
xB5zJrJHI2y5UtrXKurnOFwei4BDw++RRfJti2nZo21logONOD/8BDmhUuXj7LFrP488L5OqCDiJ
AvHtmDHwRBtp0g8LptdEK8gQcSgw8pUpH4FB9kKAf5mXMOhfbmCcPrN3ep+1R5tQI39ftJASTZh5
ZrZaiJgUQ6u681DB9fOfEt8TVBAUjbp7I4zD+NXxvbusFG7LewURn+aMaIr4Nr+jbM8GTFBZ+bo/
IXmOWgkDb2Tryb1U5Fm5bkaHjaq2JUfGQaC+L05RG8Q6BTNCLxThspbPS7kty/l69YFZj3wLos+C
SdaxvViX3p3C4wlx0JIA1KFH4XA4+xmURHPSbxSOEXBKQz+VtKmsGsqaoNwQ+hbtt1arQ/nGHy/+
mwhnM88VUtz/dt9/+/9Gkq+C2Ip5fbvWu0bvK+/V1hvRIS7PDMy588lQCed/GJawKcsU+enXTmOJ
MeH79KScAFJx6rZju/FWCyoTNHuOgQVoVw+zlMf0OafXFwm47GMTN1vqJslL1nQ/ilbL8LUUfyZS
ZV2IQTChILmWPKxuGslUq+P9qtcmmoAlpkcAq94uRlN9A1qEM/ZAzk3l5r4Q5pZqbyt6hxEdA39T
Usf63SbW10ne3Ubif5+XHkpT2oHpNyZJQdWMKTi7xn3qKWmlqQXy6HVRmWujvQmXFN6GRmJw0eq0
0BAsMXUVi6Qr3XQmEEcdgSIomLC3GXkykRaOCy17ODuiNUMlOJfFvCfqaFC7uvFIUEozw12VwIUi
UHP8DHtIiP4gyjgWXAlosKZNHnHMfu7p+yKo1+d2Q+dJARzTL5XzhwnPrPU7JtXQt5OYESkrIpqU
62PHuDuJcuAaBNrDPndQhnBcVyfpr50gdMdAT93cDaJthmNmox/Yqr1bUcwApTdmBiDIsx1kRwVq
kyeZ2UThbtt2zb4Lh0USH+3FITVTE3SHP0Lrx2Q4bKoAvx/WrbyTKDjrHT+QZM+xwUj5g2sYo3ka
KTLlGhdh3MdjAZAF17lSHd/iQIBluBRo/RdO4mESEbeNzPiRVx8TNko3iMQq0FWPmoWVfarFtoWK
/uf8Wp/JIx9DLLcBjCd0P6sX+YED6lpeUVcFMJqvwDb3gqqXfIsgpCT+vK/Uf8bDBTy3FSxfmuLo
tqB2kbiZlbx1/MtNo2zjWcimv49P/RmTZpCl5nZEGf3bQsrz/NA3EcIbZmsWnMTD6P8kE9qjQC8E
iCCh6FBvg6NW+06t6LQPPgbTX/ILnnMrMjCjWE3vThdPsNJeJ8rwQGVsJaGRHFNBsakb1PZRguNl
MGy8/fX+M9sl/XDXoazCmK0trGSsnCPFKey0hfe9eVwYfTiQL6J6wwD5kNFZVP+7gFgSxLvKc8hl
FZ3H757rGmT+LxjBxNMuhAtJm3/jMFBAANNa1rwnQupwNs6t7ZXT9ji+sfHQN/c91FlS1G5zqh2t
l76W+Pvp+DthjzXx3nz8fMoWU480SBsxLSUrSOk95MiLCLd3NOqSn5iexNX0ynCsuhEq/+7wxXi/
Q/Isrx5ArmQeSzZKmRt06cmCFtWLgFF3dNaETQyUC23fODuMu/GR8c7YlT9bEmVkFKX3Wx56yvnw
ns9fJsc3FLWYNrXYnXVSLu02NMYkWEvBNYl5LVcjEh9eMlnfV3/ltck2/a2mTNP8jc6GeTeEk/q4
b4l9FSgYHDm6+MIFGneQqREqtvXPiEap2XMFVWDhMj5RfGTDrTTsnZe+DIsun64rz2jtLmGW1pht
w20S53TdfscCuAQf3s/6RyjVBy1exbgh/6T1AckjpTXDcecvJj+PtVJK8URN6OZezS/OEhQin3lj
Drcq7JjjeSfCVlaY4BLu/wCId+sagJgze/rJrGKaY/CCmZFQH6zGFo+ETgkf4Lu8FKL9ugfrbdsP
8HGY6xbbHwJUx+953rmN9zta2BJyd/agLwLWRniw01XdZZ1RWEZrNu4hp/DX/DsT8Gsv8IlWBYbL
f3A8h+fghu/5ONdJb/yYhsRFs9LdSB25RjeZZHEnrO5hQ+pr36yMrCywKPu3dlEQWmtGK1JJTaJN
vhLGFz61GJny2QfHSiuPYkBWSrD5I8XcneebZ6LJuT3fLYS6uIfdo72nMg7g3TK19oZTu304Izks
L0RI4TD7lekyfyJR/gOKPOVkR6ZQSijd+GhBmDmP//djClOJe2Kz8ACgxkBGHiByidJSFW+36JDA
txfe7xbiVU66NU1BHIXfRbzgx4AWYD9stTFktVoFlP3htO5V86d2h8TvI+NgRp4iRieE6pny2wfX
D76Be4jNyWU9ggma621zSK4B/zXtSeU9nt9p5mvxCqO1hgfjSKjzd/nTzbkfPFsdCEq13VSAzWEb
9BA29GxSTnXjWj5n6AXf5t7BVkxjN7q0B6jY5IPuSZvgRAORnzDINeQVR8y64XA/OR/+XMKrUJcM
eyq+W+8ji6d+omgNpwXbwY6SlbuNP+nAhCA6Y92MErl7xBnpUUoKF6P05WhaVRiKrzVUimLZGBik
Jao5zLMl2pnMGulcHlCOHhAK+hlxe5jt2Xnpl3pC4UCJSstWfJVdg+CTmJUiRyxM72e3I2wvLF4K
qFUI7wFjPkLbANI3VsV1Vr0qLT2j2NoDyzdKNM/Wk/zdGYqsjPt0j0AZPfY44sZEU0TGHSR2eF7N
bPT6H8Y1pQ93T1pPuYozZ+F6a9ZuVZ3qN9q2nMr05bUNM9dJnEe+9LUcb61gyZTbH3DViqX64d6R
QRO51qnn0Hd4D3Bliauzukzinar0LhNCe87ymaOHoYWTAs5ne5zY0pkzTmyL6GI9tioYOphPBK4t
2+zepjreM2VKAtMiTa3pFPbejClEL6ADbRBxjE5EteYpNRGgNNiG7wPg+kEGWTmMv/mrqIxAEZQQ
EwcDatGcaKEE4j5UPq2sIkl3lsnOteTVuTuSED4pKAVAAjPhQPKnZukDsrYMMtMDyOgJgOslPVRB
/McNETzFGCPM0a/TSitF4nQ4EHjpLngFDg5rosOBk+d54tYhrLGbI/EswdGszCGUL+UNRfwHa9tQ
wU9A3bqa9KUKsR4OSk3YMSpw+3CytoIXqwnVL2g8s/d1V7jlxeisucK4AYeOy8Wjtkp9me2NSX4C
9Z4eVMJXYEu3jYkpZX5AvckFsAzk0inQmf8Q1zQSst4/GQaRldYx2SFTSCrCQkhgwFZ4nLqalaAG
X25AeCERtdpdNuR6IQrD9VxKeImfuVfptcW6Oy0eaOBlk34SJ1dPMNx+lgCtKDma22J6pHlcm7VZ
KfpqRCYvr7MmrqY6FRao6oZ8Z2OTL+XTxcY6T4tl+5c7NKBEUB0EWfk3MMrQ6d1itQLNg9Qsw2Zh
ULj2WpTUW1hi9OyWJFQgaDCM6mJS1MURaEHl31zIXvjuO3qUwnPm8JZixJQnKdxWDXcJqIeqQPln
HPpZp70W+gWDjNtBQ2WjeMgFGU5auIE5uJ+Qa94RlYQZjOkIPtzaGD+UxIwVs7A7wZTjiT14HNwq
kW1W74oYKZUn2JCcEVZeBM6UcSo0Tzg07KdJxoS4NaCtfDM7tIANdbezSRsu2PLy2FNCcbc2EeFX
TMAEKO/Rn5JwsA33cdsp/OAAhKa0ukltBprLkSwpUsVnvjerQxAkeS86XJDs1VS7Wt6nxzrwvjbW
blKOTTw+IvD7+io+KSxcTALkRy5g3JzKO76mZS9mFcA99GN2BxWw18eGIPCLtL2G3VKq1cEbdPmW
WFoC9r31ITvzbMLoA5VD58ECNAUrc6cBoZyTyYOiUwlJHbMRcPNssoH9SPNESAn4C7d1EP+lOiF4
PrRK+kpn/77lvn4hvdv1ogu12IV/CQ+8s/eUm4lLZSqxH+bMXpV1n5XFBD7lOf33WOfQDj++V8Ww
4t2JPJAQ3Q6F/oWmtFvtw3gt25C9TqcgOgimOxMW0CdOLOihne6LVqqD6XrkZ3XhxVjJ90yIySiV
BaPvYxZ8eGGyKHiHRb9kXIh8mTf1rs/9ZiMD347v1IoMz2J+fWZUI6Md5prUICK4LkI26G5IUZzB
nJ90tLiraOOcn/ltIXAuZsLvo7zaS88LcPOP86t+1FEMlpGLF7DV4YdAeEr5yqigNVWDWjxmDO7h
X+6LPk/K+ptaDxx9ffBXuh9HMeuEwizxDpmYxvDst9286x62D6DstenFeJ/mg7+gtMyMKX1QiMH+
liI+VWq824KInCK0DYPNzK/KHjTVT39lZ6zqRmLQqLX+FAfCget0eBoH1LW2q5IV2dE/B5heTJsh
hsKHb6xUbcds74hOtNXkIYZnATSNUJBQzOLI/nZe5PRd3yAxzDecGqkVlyH2bjm6GudnzkOrIK7N
W4uJlmrzZjyambZT994Ntnp0jlxc1K6EqTHBWTvJdch3bOmre8NTaZ8Bs1+f9LKfk6kfYM/kgj3q
9J+epeUzGeLQ4A6eCpVeJ8398l5HQZWpJZ+msL59ZPd1VvA0j7KbbZrE81OS95q9gaT/kp7294T8
7qWMHtrUDypnH8NmpfbqqoUVQNnxNMRmsel6aMHgqWdjPG0OBiFfAVlrr9nt2W7BaQ83rvSrrkiy
ZRWUvURM2D1ydbFHgUjyoamXRKlGVxbBfMMiTysEiys6kXP0VCJvWbDFRJh1hra8WtOzaCfsa7EA
e/URzqHpJ+URajuG89WoNHi2wLAGcWT15NQc5VZH3NxZPE8xil1KqzJHv5NP/3Qbe2e0Fo5BdjkX
/X8+2ptE7I6gsd8XlxP6fXjRmZd+jbYleYan8ViMIP0kiJxhiIyO2R8dtoLuVLWSLdoIGXkyw1Z2
bJHMUESQneLN+rMThmQJUaZqR51xSqh1r9jkEwvNZlTgrlL1Q0hNK+CWGMxR7C/n/w+LUVE7JI24
wEySPsw8n5LxbByCpOb6joAzvULjLWrqrlsDvERsqnxN0s7OJHLxFGrG9gQVX4lgLODhqg+VYpS8
sdjilUTRxu8sCGYjow08STJOaMHGDTvlr0FhPgPwLhgxfbAsrnfv69VRb+BaEgFSjR9rfbyMlzrI
hE8MlPrHxVquPUcQie2GpblZWqZtQEqNC78rVh6Yo/bLtl55ofp1iZbxR19AafOanubQH8gx7MDt
uQh94UKFHeXdlTU315S+xC1MRovcINVkax6hveYpKreHSY2lKK+1hqSyr5Z/Ic9o4tmmAKZhy4nZ
hnyMIhfSB1gLeN8grMj3Hpoe7eigGo/UmqYnq/GVwtpq+eQTovjDfjPSTus//fm8G20yI9ZtA6jV
+6Oi0qLE5Cr+RDamKnhaDzp4kYVrplp+UCFq8oWP3B7hAJGO8xMbM7Abtl2DRt53BMLJk4wIH6fn
Mn2othjTMhQCSxHAydoAPnxpDve5e3kmMuD8lnyNH4SVBPzIYs4rYG2oCaMes3TWbNo5qI8VqGmC
p1JTlKdLwXzPaukIkwZKBalloJQi6EZLhhk3/0G9DderF+r0YsW94sdj6O2VsX56/QCFzvDJtwMv
oxbLxgADihVV25+PLDMFzxrFsRgVao1yxCD3aR15g+uriGUlrCyceYWIcO2t95Vucq48fU/VF9jf
ulb/MYzUNfIlNNthfLw6hj0eZLSJLV3IMzt31nxd39mJ3F8R/G3PLLobYHyfZbfcBPNi5aTWFm1S
PV4h0hvBXEguikaC1BamyMNSMK+rzw7rKMBxEvF6MhN5wijGRO/iN1GmefjkQIDD52T44ol7n6d1
A1mOPyYSjORSlDMD8nOIJCDAMm3pAUqA7NO6H5y3uYAfGxY7OiZtDE9AlR1f4v0r0Ogwcja27PEH
HLfP+bq94HJVYFsmlKl4eANzammyBb6XMfK4F0dC0zHnfaQOOrgGddPIjrJeRA/VYdDkst0bKI1p
DoRK6oi/BhHoeNttBRGuzBATlrlQryY/6WcMWUhnzq+Gf3hMNyTmSv+QWi7Cd/TQTshcWWhYULPj
GXfORdvvELEm90eHXItSJZNhZuaxbXxqNqAvsgtxCqSnXX4XPxCAlqZFyMIhm1oUFnxFPSlarZYD
zg3GMnr6Ulp6JSwiBAXqWja8HQjq0Fx/lRDwg4dE6Bdu+LTEOhB2qedzeJWikzZRIH3fXk9iNK8f
wSiloqGfWO3j9fI/y596E4+TdUVO5BLOkNKiSfB3qhKzyOaYtRCO17EeqnnoSNAVLRYRP3hGVOzS
7ivgt5HAyy3x2SMNDqeiFQMs13KywJPtuXolZMlYfJ+87MpyYVL/exlRZCjHu3NmV/AHCMo8lhoy
n+n2nKI36PuLR1kY84DTEdidpwlpQcXWjrEXPpAE19XplL7CVfOgLLRx852dRmvXXVv1aVR6EW7k
F5rafwp1oJ+MdQ7i0959nJXS/rrQ7tQ8iCzXCpmO0M3EMrDL2jXCmP/GI7A2lXmKTLY9mXJphKrq
dRGCmyrtia438unj7StsQlL2RZkO3UWLN93hPe2j0kfVpRZRPnc6l3o44EFmjiI6JOIlGT239FJe
DksOdIHpuLXw5M3d+A8eNImYIr6+2ia6D+DZHMVVmvarQGjTYW16oJWFSB6K53jVvVVWii+hK3cl
xQFtYh4Fi56jmWn5OSnzYiOaFwvYY+73Zm6H/7g9PmqPS/0EqwDZQxXkstrH9rDgpjxepQzHqgMn
5oYAq1YcTc/thqhgmFoH26vT2KFH6SrExCzmcD/UrX5b9QTWuY5EHd0WgrMmjaprefx3c3s6RLbQ
/k6zCsBpOITJGFzqFRJKDPqyVOozJE5QEtXlHDNzI0gzDr7gwsOr7L6vl4mQoYDBgoycAmFDL152
776e0Cgk6Cra+pHLV1ZIlZoknxg/mht/pfVGoO8RWyO6PbxvcQdtPRHCr7qhllcHt2jZAvDsSiL2
byDBwj18JI0mH9RF1Ocm/asbjTzblb7qkfbJxBqytuufgv0Ml8gYWVQPDYdOGNhyj9KCaGle6tkB
x+cskEsAX2GmSCX4ZSaG8tYHXzPevu8JcNJj+uFyeKu+bDDH6s50P7OPRa/HFYVfQ7Ni/dq2EgNF
4pGSczjJOwTnrFW1PKMieE4FDnlv2E1GPWsSQ7UpFulOxDlKGe0J0Bhw6jqG47JUhe0HRleyXk/L
WErrSPj9HdwZd3HWfvsjejJgKhkDRljIk40eab1fWMu9EcZN2c7FETNE8pGCQnr0Mmqz2qpueL3i
sgzcH82ob5AGdhyNsg90JqE0VMq6v3ntbSGKXbNkNxwG6c0Gaah0GADEbfVQnSV2oUQVaDJwKq5J
i5Mjq9TwSjVXKIFy8qY28foPdN53d6yb8OaNNlCj96L001/nb71Rx81sxMF0RkalGl7gwqp9pHRQ
6bS+jfqNrhzY8UofawikqStD2sDVUGIqJ8zkUtXj5gQz2Sjt+PXMvUCKBm4rgujvAW6U//KUs/y1
16Vw7stqhs4CGK1vR1WtnRPd1m6IuCJ+VgyRjtsOAvok/6EnGI8Gi9m4VlM2oe5ChOU/4zwNoybJ
1n4TprkmCquH4/QeYtRFJ5GR75ycnCOHAgBgHrVwIqKJVaCzYTf/8Dv8cPnhgMg+SfD2P8uGn/lh
WIy4oKjEi9oStqg0g1TtfXya9I0+36B3RHtGklsIJGGN/Ijmqma7AgVU0MTQ+McSdlcWoIJ+aakk
jCl4piCZTAJRUfmGa4p9VrpIxueOfq0wPyLOGxsTm1vPVi+XTkG7f2c+SLqF5/VgB6t5/EyOBQBI
bn9u6KfOnaGE4vE1bKY311bhtVR2Zn5NFdLmeW1eCGgH+dVcC/pTl5dxH4zHpPeG6zvLUtckqLpb
F1p7gJFtFpA0ufqpzf25ctfyfaXf24V73EONiMKnaxBeB2AFynyDUmhpaRcblOPS2dCn6l9DvpDk
V/UhPnrIcRPFPHK2xGRZCitHK1793n1dW3wiqhmrbwzyKyMBEjFPlZaxkCWYWCRUoULjNb7LRwp6
kdbCDoLvuzvM/8ouS/zDSy/eRCyxDWufLeLzsOvnVmWhWxiPOEKkz9LAxDRv9rFrWgaOaH8vfZpM
JKMDpU7/7cBxCUuCLfVFJu5qmIDNpy+io/NSvoWOVQSpvu3oc5OgbK7H4uO7ub8rvOxHy0TJqd1+
FdkbBVixLFV1keEM0LUbNVr9zvl++RB++vWHxGYgAflBc3wN32SoAVj4w3tHYU2nCv7AKZJ07KgI
Vlt0wR+8pqT93r9CghYj8TEPd1LtPmUVfkSSm2LdWlyZsRDKyfmVD9TdP5XVubHAn0g9oKuc+XGF
fpU+vpDJMQ9t84RscCYc1M6/78X+1gsjXNCRj8kMEAE/XS2SIocxsjRf451YwC6mqJdUhFi/TdPD
LZ9kRfK2qQW3p0li640dhm+xXiowFkGf6OUY1ExffP+rLnByhnz8DtQiGguDOEOgkJj+0TuEgFEr
nvCCtta5mee+PVG1CWCDSpKyrSB+yJfRFdu7qO3uqbxDfE0NaH3IHGSJVH2+TwnwsyLiUKc4xjcx
+Zb0HRgtBWVh7tE/gxuhab2OLgOzJDKXuaiSGKFPiikwFDxVXQ8i5BrTXAV4AKyzkDgk4Zfh9VWi
gA0BhBWamVjlaVRE5BfSvTg/YDwQAmMHK/eI0ufrbFcUZ67RbxmAY9gizJ+WIQJHRSuwWiVxtqyW
vGejjnnbGkjiNdd3cEkktIwxLZ9rgKyfnABxsG1JR1hm7cbgKB5P3n9PRjeK25V3Rx9msSBvXE6t
mjrRzdTPLXPXvVJbWzim4lcPt4rcJSziWCWKdXNgII3Lz3xcbZXkCApZypw/tb+5cUaDgGqf20ju
huYUUXuqnS8n+pxqaoPheGG7LADF3AU4d209tVH1lIwOp7CWI0AH+iQC5q128SIswOMV8dPSWkjM
YgbHgYtPxnLMzndORS23CNEl7RFXg6Ud33LxKZ7uXOs2hWYDHE5IFnoRSi97pKRpm66r1FGRsPPv
9TxbGBZ/6wBwVXqSGV/aXOvyszHVsb6giUSyrF/HpOE1VgNyoJLPewryh5tDjczfLIusZvpE+U/u
tWkQ8JZhSLajQTwpvcucOHl4+qqaOV5y0K3i0GEU0nHsDVMrzJjOS3q+TyoDZ2Dsy32nIH3nEju5
018h4DIp87QOTt2hbE+6mXZBAfDaMV7o8Qje6z1Js9BBoASeLsin1R/Pjo2N/dUw89DHFPazI8Tj
OPdZk31rnGNm9wtvshOG7tCsVtwSKbMHGYb2AON0vUxBO9z0XEwZw4tMjig4ym59JqHCGnS7E1W+
3KrzbJViqsbxYik+0di+Ti/HR5LorMS2ILFC/18c5o1UQnJMwj7cJhqgkKyAPt4QkpeEERILZKtW
UIDxjpNTTWleROBX6PPK/Uxthz7Am/2LT02J+zzwbvyJYAMChBKW88rGCZ6CSocuscfITGnZysUO
JWnadZXtXL+0EiCG11DbNs3/J9HopIj+67A+6OGJ1SXnXpvBcK+G+9w0uiHoNMSHZlRsZy/aubES
2LSIiXxGGvRVAiN4Qw1/jYA0PyoBputG0Sc+rm3l44oK8V3HVoCs+2a7sycQcSmYC4mzmBABX19R
CScw9V4DVEJ3NOLGA+fYVQ52Vv+uTFrE2t6PkkHbDPav8bka16yDtgrU7n0ax9yNB8vBiBCNc+WT
tCE9UttRgfcAVbp1ndArn7nqwFCxOFo3OzKviUuIk4qwu4AIxfy+nFVo/nzH3TcrT9EQ2V8mVD4m
eLE/KYDLXM0DvwFSWWE21bNYs4r2jYseE7HREBJ2D37pymjeoD+UB1M/Oj5vLB4f7O7VRQ4SB3kI
jSDhgx565R0rzaKsFb4Cni5XzXp704BSFbi6X9A31AU4VoKSpa92rBK+TtfHnuXobd1tbRRsBiuD
mOUQL+eLuWbFzDHYVgiqloaViPgW3xSJAZ3DWMkTYTaR5b35iWpNnGiroR7UlMuOgQ6E5wZm45Bt
K01rjhJ/fz5M5mZXMPfGzMUkhwqirK0cO9VEt60WSqYUl8ZEptlQTG5fwykp//mzNQ8y5WT8zLJH
ukDF3twFUaoqF4SzCdns+YoDrGI0vODM8tm7pBQLVbrIf8gJnypxj5MrKEFm8aKP5piHardKqlFj
C5m6APrj/lUqNBddllauiwLupiXDalVhQiIzw3HiY0rqtHEzsCT6mllf+hubNCeMdwR2d3j/nrjS
wzWzivTMWJJOlSAgyi8LQaVnUn36ADQz1yboYAw+fV+1SJfXQ3XF/hp8eQdmtg4axoP0hknzNrYU
VCtZv9VttTIwPKvDAgb8rsBj6/bM14GGz+qUGtVRCAfCDMKPHLUlRc8LNQkzD+zCut/Sm1yJ1vuD
p+0ekd9NfIFbFwbnR0sxvScqSPoqfHkjoKrK/v+P87ET+CH2jdRXAWR8yodfUixiFeH5M5txQGZw
INV+58ULlV1+KsboSqGYrkKAd9Agvjck2TOSsPENZbUm/IU1YQrb+Mjg6z2rsDNgvTR+hB6k+ezS
W1VuyQUyMs6Py62M5b8nEVfxsvKGFmOI1z/+bjBjGPEpBMa9vCZEumjoPJIf847TMqN/YsWXLHmp
XpD4v0DpvemwHxiQnrbgP2RJtxwTK6gqOumwmzaLmvJzuvU6TNCfEtUF2kGim/5Pxun2r4JcSBb0
uIKUYl/8r//TyIBjvhpJD2yxD6OowNanSS4HA5EvObZF6n3ifAKXx0aVWkJ01iW8TPmxOAm4mLcv
hoFGrCE3HFL93xbZ3gMIz4PzTsc0KyatZhBcw/3dBLPIwVGSqzQH8q/DgOfZdfVpFcUTpqcSJ+e6
syTdxIIq3Z6+9cCk4X4aLf3YNuVb+DhkBYipIvl9lkT5BF9wd0JCsLqhhRnUq5kOOtgn+kld5Vfx
AUf02wdtoiOA3yezTV8WUxQ2QnO0WgsK9VuUu4uL5VfWs7zS7Jg/VYNlBNPpQgdJep475oH/2qfH
/2eiVWImGepr238uFoo8ZUTmRkwmEZ68r99Z45j/39a78yIKEJxyuEGOQ3xxGM2YrtmkhTN0sznP
7oo3vshzZyxsFr+HNqBNfYoVL1KNDJtf4o98BvIZU0CZYtxJjA8rm4QhgmBFEk98ALkhkWSqNhY0
z8Plp4EamYKz5i1sGMv8OSBSrk0wLoD0wocx4/n5Qv5Whzih7IabTnzFJrelFH4IkjsC7zbi/MqB
Az9uVEZsFTt6aT+dMeHhZqNKbaWzN2NRaJNmK5GO/lgdBxqvXeGFNBUk8bs376jsB32FHmO8LacU
8hIgzBz4S3QAqzzZ+9pbrrnHZi89dfrxSUAJXla3j5kiSoTDgBzyBj8jWnDOJVgrgcgYuwjMSnM+
Kq9ivn0gf47X4duEh5srXnjdsLMq7uy0TL8TUiG8ByMEwT5J6adUykWdZbpbnW6nyMlQpJg2jwNq
BCUbG4nekOT6CEMSO36t3A0Fw1znPtdI57zBDjpfklvwT79vi1Xl52jimfukVB/EmZqQWfDXfgOL
SOb6U1XTcovWUwaSPvgXcugYabYyDNrswEuKHpwraojDc9Vqkx7hrOawILoSwPTCiuIV0Fj22LWo
KcdVDfKscHwkOt091F1BAhyPeNsN1S+RC8qTr+tT/FI3hDp8EfAqDHUfhuvI2qJ1ikSizsv/vF61
XtKxubGtsGsau8VGehavTvHspBbFnfOAY5A21p5oqKF5d0vlHcy3pBemXaVthcsDDVT5uxmM2iJ1
0B4gTFV3D6UKxHLbzICJO6TI7b9lVK50fTivwlX/fUj1vBzMtghpKMuJZ1ozyWT5apvEvXKu6pli
QhUPtYqwIyUZOkeRjHBDIbhRqEExiTZykjMR8VIKubJK+i+3t+4drS3VL28vQG8d1Cdfmw1/zQ6x
Yxi+pH9OgtRJk+t4lxQh9X+gagvpE1f4GDvEhfEehwgf7JuoLvRGRZoNLekV3rjQtmjgf4ADFK4k
JoQHG8OfJ7N/xH4YUgXtb4tVhU45aUobGXbJ5uuya/vqptz4gyrGcth164rwEZwAJBIYgC/mwWhn
IyvZSYsSIGnCW9dzf3rRWrQ+k/Fbw+24AaQK41ZO4FA1NT+obsll1fKBZEjao5BKJdnX6L8a49PY
k+Pz2UF81/jBkfzzO6AaR4wjP846zLuBUoIWhtQisvOGwHFG+S8GTe5D4+kz575q5B3+nBJK5hBa
oCK+i5XsTI2htyjK1RhzNjCwNz187kzGxYtKst56XKNmERMLOu8fF5FkW80e6m3qVTqy0Y9AQ+f4
Wowx3bRXotX1+gXY+b9Tbvs+t7XWbZpNpVaGUXziuxjoyuUB4UtW1sCP5q7tdSrgUwa/PNgoEkVa
whYXzNRCr3vPwGvuk5qTSCw1wrDtQ8x9kosL2qsL3AQ5OCzHokMJ/vGAEr9HGto7F8a7SLqTrEpw
LWxTEG9XvEvDAyOTtmdz3PeP3//sYebdzMsJbazS1wywpC4cytWcuTVYeVgnCHMFSOV2TYBNzlbn
JTGTH6SZZDF+DVWjHT1wIWdaRMmBiTtOftyhTJNUIUFondwntqigvS19QKj8UX6iW1XUbxbUzmyn
3nCj6kwfElwXaYAgnklSVYopVqhFruzgfsnwPaezMFliMpwAtLZad9XvRLUkflACRzWnOKED+ukO
V7kNWxTchD8oOGNQltdnrLDl1XSk7qEw+u5LAb31bOhFfQwoEP8ku+TFr5xteqQSYkDNWaONtrYo
7JrcrC2tvXrB/Fs3GNrWUTEc5bRjCvINhI6cSWMPj7+a0uk9+XjPk/+NcrSj4+gfheW0NyCjPecP
xZ6E2Vta243rv/jUcZqLOXRIdsePn+dsTygeBdpwI0+ZBdWPIIikbyVc0vKk2No+RJqoosEZdttn
GQTnNLjZtaErlrGdsUTDIy+DzCzvwCed454Ft3QMLg1IzzRflsCvUererzJWqmWHmoYxW/v6GNba
X31hUXYyoEWgzfL14zqXJs/GolCpOdWNsGIxOtNeNk1xm6dhDjHPHSjZuaOjHuSCOyo3my8vu0ev
9eib4rArzDrIDG6l3pgbAoc19zxCFr9UbPNFmwNIKGpvF23K4tDckLQY5G6jx76+/0Zfp6foIqD6
M36xlVQA93H98Hdv03pbNOJXsUO4HcGRRf9ZV1aZxRpettfnC7ankUF0Um+wGQhIbGfqFcS7Br2l
MYCLcVTG9XGjjOIdr2gWtZ2gn57EqUbal8Py3vzctOpypjLnLSIyKd0V+rnfys56fnbTvQtAVU6r
82/da18ZcnLEOyPJNqpV8S8rrd53v9RYRfmkTr5gZDoACd5Ve6IHKui/0d+++44Im0rpyxsgNXLe
QcbTfXBql/tf24A6jYOaJIid7mk8LWnhibWgblK8WvZvQ/h8mB4pGp7df72l+RkgxXFjwFpBbIAw
S+7MvGV6Fm/S+XeWJVrgrZKp9ZWFmtCGKHpsGK5y+FKBH8HhQAcBf2Z4D825pifBd2QtNMVD2oXc
k1aN3dqljc0YugP+aBVk3VyH7ZK3aboIzlprN7Ii3tE3ViOi4vfse+6W7SKFQ4o5bDiofPKbtEad
iJtFd+LHMOY31CdBz40BntZksj8CGlqocax/KtfamE+z25QdiRb3W9hsAKroiK/GxvPGjfvYdUwu
WTUTgUWbMi93D+8PXvwsNlJENwtfpv4RiltqqozXUVS/PiFXKDKqhEJXQYGwiJFzkzFArh2EhEsh
hy5jBPo5pyo1G1CaOrPBZSqu0JFUoKNTq+pHqG9biEhlAn2tqwXDdKkeo1k52lRHRI5F1gQdpTzW
+Fqh3Pr8RZR3loe4OwU2MK0Nhh/pA1WKoele+vO2Nv5x0OwJXE4VyajR5sLcUVHpI3yxfoHHE4FT
OHblu+JZp9ZFoZCupiuXTin9BWr5+yVOiaMXnCNsxb6nbQhI/inMr60+1ez7F3JYZMzGSzRooMnr
IXvolLMymmsMAk4OxLA8wuCPo5hgGkH10s4jhdCfeOjtRm9teMnqeliNBC/Os/IZCEvIIiR9Ju/t
9PVXYEvTFimwranYcGp3fwDWuOrnhHqbGHW7mVn6VkfCCMJjGLvFFWFuhmDohMtosncBTw+V+fHy
AdHqMoJFrvfE4831Z1rwgpxV1+uwlc4pCEmZfGjsvZzw3SgliGRCOeEYdg6w2GRQet6BJCBqtsfD
/MrqYUDhZBu7xXzPfpy0J7LEkejRPXtYXqO7QwWEqgxE3Y4edHUOzWEGx7yKz2X0Dlo/mLYz6qfS
e7e3+o6cJ9H7VyLTMJYGDNDdXAbhf8Tadbr33AR00qpDCIYqxi0XGTeZiWvoIof6pwvf+Y7qRqpQ
yJ31v34iAnQl1iMrG1LqoghZYml2vqVFjST9Sjo5IsZLAx7ZEGkUocGoWbbWZ7414RNoSXP4jRA0
NKo/LowoYTJdOi4mFN/ehjVLScLYQylSlBbEFrqNQ+hsbEjq9RTgxXOxlVD9OmiJc0YIQ2iSFSnx
7m5PByZDXxHb64f0d/rDqfNVSdK/cT/9b9BfBHGAEwvGG2IoLNnSOLim/leMVD7YfE3xQlkcNYkp
B8EQK45a3PZkzXx/ivsJaXONgmInvGAkwIuEeURRZbnnENV6s2OcAIAEv2qZSpxUdtjXdjDpZOny
D7JNjChx4feDsSA6Cna70KNqV7LPKimkvMyvJ3gypruKzsEyTBRaKDNd0M/TuQjfO3vO1YKvy2X7
WB4mFzfFzd8GSJQKDv8iHjKewFyGESbMdYONLPPYtjw6zXN2+3WtECndp0URGLI0MMNWHi9xq9Sw
FoJmEXNnUFSSy41uNxU9/uPcJ9vrNuRMwT6zlYH/Pv9aIldhM14p0kNm2QyiCd1nhhm6M4Q8jR2i
Wf+561u72dqkCYSjsSHY4hvkcKrWAG0SLs9kaKjE0Bjc5XAz2duRWFYZafu56Z0pcjYVKVEL0Tkm
sMd1efuFR51ke8cGWcHQn2/LUyNswSQ271hxN5JWj52XlEK2qi41B1579WlEkTTxMn0nBb430uWC
TwQ6e/xmTyEuCNmoL0ZjIyINckBafTj5KeiFsLPpGhRcO0V+QgIhvT+mL8rKNv7hX8a5m2oITGZW
uPHMSL6dT5doydw/RypOh/xZMTaeB4V9qUC1aP+zS0919/KQTEuq60pxT9Vy2tA4wNyoCUWk6B7U
Q+fYIJRxbTfsO/ovmLFhdO5h613KUgX8oUDVOUdl3K6VYiT14BKjtShdcUorIkv1YjYEEhsNaxjq
+PS3wSD1AqfRAniTCefZ/ufo5GJgW2fuJFs9zTy7wLoZLqRhES17NYolIwqjCzbnR3gf1a18VywU
qjiH/H5OwW9onbbYx1LhCTq45/LjoANb9iF3FLSIlqsmNgyK3ioguHeEkJHARe/I3i1JUAOIABhz
iVa/qvyrMX7UFJANNfD0TgYibdEnHXhhb1dRSRt022SZKWwyYKSMHbIqwwgGywSk7f4v8LKjGRff
t9R+fQHAcbgCbo7rPBrMQ1ozfpUET6MaWgwQJjqwGOfK/QuRKw2uHwEuZzZsiR+Dv11MHyUcP0CV
0UPoCo0FkIFZ7rTLE0QMoYq5VYOy4ods8BDb75BKSr65uY404pSE+VoAxjP98v7e5H3ApnaDur29
rPX2xqpMwVizng/dG6VZNl5el4umh41LA2UiTADKl6v6YIJ7/ut/5SHTI7IRQHEd3xNayc582Qjj
4hGjVtbkQYU5c02+hPLEp2FA6iVyvrmu9M8bENlQ1jEjsg2v/jl5vdChcVVjYGZNcCPNVi/753nr
ZtG4Ufjbr0lnSjCFsGzJXm4MjXjV1eK0Frv5IL+Q1HsLh8kI92FKtdwT37oYX7NuaJ4Lq0N3VnfC
dkZj6fCMTTkI57w4+BjJPi9rjdokBaUjkcnf7+TgWmaUIHEKbnwSvuAM+67xagDRjk9e98LWMmjl
7GcxZ6MyORt9Nd+voy4EWeSGauCFErqXSdBzh88knnr/ilALvoVAuNcj6+N3lumYpMYT0b3SkMXG
+/7CMYB/jyFt/E8c0YGzaqjST1Ygz02VM9FkEwQS8NgHVqKwzxBvMjzC7hs3RZrcBDAdx/dUmZuw
H8nEXVWqjANtJrIQ64dJ+qFk3h4KY4O+X6IULokVk8ZXXxY72ZKYamlww/QNF4Dg27bboHGJLVSM
gREDyzVDp49joQpbztnY/+/p2CdHlDwNcGHNHqHU0bQHzFoby1AYVksMVOsjNOALoFB7e18jNPEK
20XF+sAedE4VH508XzCATcAR+7WodBsoz3EAuwVy8HMR0o6cjXtBaRKR32JTmRqhbiDOROxwnfFZ
XpC0K5AVbnGLthsurb7isJ9DetED+t0S+o4QgNWl0wM5fznXOVwXIGbsetIDcH1v+0ScA4EpUhJ2
gEvfajUmhoZf8N3Bs+Fex6V9xgMUG/QJ6xKJVj79qaprxDbGaPt0CxxwrlhgxtFL3PsgTHSMRqKF
1It+YbM0vBzR7kQMZl6Egj5aBxnliORA53UNfDqkJpd+9qOY3ZtK8Be/ul8l3NDCvVG+MZ65ESCP
tNrrWb9j+qBzip3DnGyNlW7b6alVaI22iJWtRnJTqL80e05dpozI4+t4kYDf/EfDNOiTyATyqC4t
8OqJu3vKFbELQhiEgWkRpOVv04DMz08QpVYoKPzOCIlJZFR1ivB/wPwmAVZ9kGIoC3C9By4igIAz
HUEbKAoIes65TZnMdM0KvMCVxYURJphf7FqqcT9qi0aJ23/DHhDQgwP5Oolxp4o2MWEvkqCqYUaI
SUpDQyQNsgVeDaCPQfG1UCFIstVYZ3TUbGuJbxGfQkA3oCKOb4GIjlwDXVgGEOncxssdvrhnzsSw
25hz84zOORP1s7p/flvVQbDq7gNWhwYUDu3PvSusvaEaKYlPAEIsUJqnXcaukuYpuatP+W5TjTQy
30BQFPg15S3Tf9PMvZnFz7lWVqRbS2oe3G7kiMRHKV4mzF8nxd3PhTPqGpvqnY61ytQ7rAKkP6np
yztQkjVvhg8ibrqbW7qybUd6eDdDdSGQgjK70Eb/9eY9zIEURkJxkqLHfhPdEXXTpE7RDcSdZoYj
ECnjKdzm0vQ+Rmjcxr4NokqOohaDLRvyGTKjsLE8mo70kDMaEgBrbOTUD1ucHCBPq5KFmH6WrVa/
qm+SNpHJw5E3DR7CwvEZXjLb32QVQ9RFG4tbU3a5otiUv5ttWGj9sziFu1m45aFP1wNTUlPhI8ht
lydmMqzVEJ291HxpK6fB5qne1cHiKSti54TxKOCyoEEiKYUn8nZh5B8nV1W4i63iPq3js6hKGXUB
eKSwBi8ZKPvk3flgil0p1sIcWJRAGzQAOqfkK83Z0mrem3rCMDWowHJLsexz/23HhrXREpODwQpS
UTiaabVmux59eebhA3ySUrUS19MQkSingxGa4pqFWmwPU+IgD+lEqrFnb983ldoq48Qlm64TaMZr
EonpOEg+8Jx3phi7Z5lAtJlfmKDDC20GdGJ8XoY/zfsrOZv5qOaOJCndCi0uEvT+efMul9dMrTNf
PYVs/SwfZO9CZznoIFGzGFgQ2QWCcAloJ3Yy+SbKeIrpNw68oG/p//njniAaI8iwiBls7btCdxKj
RBBZHfQqI29kStwZkPQy3n1OM+NMnnFTs7TD91w2zv9Are0NHKSCl0Ry623ZxZT+dCePEqAJpJ6C
OW+uf6E1yNBnxYveaN3iOydyWmp3scSnT2Lyz+NvVyWq2YGRtrC4IjxXE3su3tmWdFLU6KhMzX8x
iMKdWVYEKh/0jjo9nPuuOMBTvYcNM34SFHEqK/ryDPRJSfVPNvzCTbwEF/G90R0xEd197Zj0J9md
BenmnqaMWX1ulT+cAFNLha0uMcD35JrIaRo/VM2GkuSgAwoAzuAmV2mPPfLXBbumRPwIEwVhPP2R
YsbSPrasA7JuomAQshL9hV75RjQ67bZk+DbPCDKs7i/xe4Vw7pDIS7HvtSku6bp5TUNyBpkQqguO
AO9o+Slf3EZYe8ok9Ym95O0WZqvo3h8o/f4hO8fCOq4EjTkIAcdlHMhIZGfI6KyyEATN38jQcFiE
gMPDlVRTrPxgkFLroboTP7yq5F5r4mxYKCctryRf83MNAFiE6ZMsNzy+QI2SzMa+ggLp4Q5w4AwL
yOCZhMY87coxoDTcHBZqqvo6hpjLDvzJFpqWGS2SzYFSMLjPU9/BiA+laU8dzZK30setAeHFi0FE
eJwsweFTgU7O9I0I7XvGmBpopqcODYwlEo5o3nrVGutLD4yAfM3QZ3l3P3P6ls9kMw2Ih2b1Nxom
hN8RHfW8HSrpiHc53vpHS/V4GTlSVNtk/htbUdjVJ0TpL/9woKDa0kzSe7tHmJLN+0L7fqajA17q
+Gy7RzF6lg48BegrVWdXEwBWS6gjF4DtjOA+XmjbPkvoxTFZQV8z9Ch0YBHYJ5i2h1UwUFsOMJVz
YngXFh60nD6Z9m8A6waT7ZkdQXWREctAZzzn8au1Xr33ghuEVIb1i7lcugIM4Spu6Xvf/OwHqY/G
qT7UFvhdaPtgOpB34YcXBYFVZ/YdQ1P/7hNYr2RdbvzHdEGPMzUcXEwyqgjvL7JhCMneQPSRuHq7
PgeFRYLv7DhhzebmabjEspBJ1DFf1z6TAfG/BzvAAMpbatrTUIE650Gjfwswja7s9BwoTzoB1znL
YDUxqaL5AbT7Sd81hSkPveLhJwPwIwtjRmBUJXO4kZXMVX839YEOeZY6GgkfuEd5a04trfa/n6Q3
YNyCrKM543BO3K9RnDvyko5GpLEwo9Kv4nUeyLe/UsY2wRoij9a6gYxvvNdhxT3amQDy8dLGZfGF
9Czq5vsNSYqC08Sg38AGIZgZo/trScd7uKa9W5f4cnYCFgax0NMypggnKDpVwbkRguSBvu6QlSW0
vriEUArEdZg54mzL8xdKAQGnDotVZR8kKsaur73Z18uZWvLWXwC5NM5ZG5IOXFcBatWb7X4weUXY
I95+YF3nXcyGcJf1prEqblsHu4OdGsKsMWdgjrn0ZrEbG2j8GV1BAG5n2bPBiGnJNub4FTMe+Efd
LwglOEiYPQleETH40jR8hAlGYZMIo9DWmUQfAaFv0ISgbbQzJdYGu1ddLKDM/YCW29om0Hfb3/kd
qoFGxv/916dUh+vEYBCkYdixLOzL6FaBpTyR3x9DFTinLwIYftbihCGN+44GP5wgs7Zap/jGy4Im
dvCZi+rsrOhouf/MlbjfN+KU1nvHKWf1vqyXJ8fsRR2tGV31yecAGHPbgMfYL7Ll5+8LDKITxvB6
ehz0r9r0x8L87bEyqdrsfCOPY86z7jR8Y5zltW/vma9LN2WQndkObUUtNOWtu0Gj/XMIwzkvmnYO
+aksd03AfZKwiSzopF0g74SZBza76CKqd9qDumH0e7hB8jnx1jUekSIw7VPDeAU2D/7chzWWY38w
U1sQIeC9gV05StxXP2DPKsTpAQJfHMZ/orvAPENFH8EOuJT7iGPyFUCT7afIQHlwkN95PKc1jmPZ
XJj9flDAxZ0XwIoE+3cpxDen5etO/4I/X7xUomgqBfwEnH6xviRjypME9gk6ISLo4Ij4p4M+k+jo
wOyz3AzCFBRbb16/VxZ+pI1gTR1oHLYW1Qes+Qf4AROazEvhO5w5JPyLRmPaKbX1ifxDONyWhVo0
MjVpSOyBCAXejowF5fQqnKaQVEwSmDiW0FagWU4i7RTRyKpP5lrsdwYZaQWxYqmTvQ8tVpN9dReS
81Iu+8tflP731bq4yVG1EhvMW6S/5t3ZhJWOj39riH3kO4j3kZpRICFCNAwW1dH9ySOzbSoMCy6D
rKo/W4pJDcMrv+bwnZ+7aA8ikyAWT2bmFH9gWLgnKkPoIIKawgj0ApUklXslv8faO3s1D+LoIrM5
2w2/F9AE3jG1tZg06IP9azirnxxetJdzcwmlFPQH2Awv2ajrwtzseokzF5GuWvOSYvy/r2blwXha
zwAEdcRY9ZsRGDiMwsAhCNb3G4PeO02R4uVK2oDLRLsTwb6gIUUPDt596xCCCrbdzjJjanBA5ZJd
40vliNUeVHuvwGIXR3wMXA/dGzSqzdyewCLTg1BiJii6YIHw5C3u7oEodfAzSHHPH9PdBvPSR0b/
ZxkeJQz6D5rvO136/ZH4vFc2BpthMLAaWs2A7+5vxJ1xIkisPZurTwq3PU9aqcWj2XplcPg/oKMZ
7VhE82KWHe14P5xugmrhkopU0dRhusru+Ek/dRA0Q3k9f1+uDc6uEH3m6/DQoNk0p6MU70CxcXdv
ERIAC52+l5EywvB34DGBNU0uA+jjFjW/+Qx64yCJtiTYr+RCx850F6GW8WB6css+kD6ZoNVNrf8o
VO+Pcc0tULSfZX8hihDhM3iDNv/+QAwbytGr9DCu6oWpKI/zvWRYIBvhCQneiLkogd0y2o9KImNG
edIjBcldK8zgVzdc5ivlqm4fKNxs1Swe+sRBWTAoyegAZP/kMhBPGzqfsNs3FrFuyBTy23+PXAgI
7gb6f1wlZ5apxx2pfTIL79G5MW+mztXw+/gZGag5b3J/yEKKxE2PR7yQs9hhTkdZKns5Obd3lV8o
DoaDdpfCW4TncbOhprQxtnOoGCegfBSDbOEswLA0RWa8EXl0SBLHTxHNlUYchu+pkYCeTex5VWIW
WlPf9cGlUKOu7q74Gd2uYJJqbngWawDfZAVKGSzT9YGeJN9T6aUPVGWJxIVQ/VVOH31y0270Fvk/
cqfLEOh0pV4WB654JbDQe9ZNTSrUtdjGGeGcZAfiv9TD5FAAnGuxiei9+tTXv7TRM9lLdWVA+PpX
MnzsLnD9b2PXp2LLkld+QaE9mJpkL4/Jm3aeyFEHZHYCxC3PKbS+bYQ8DM9Dm7BEWeKcup8mND2D
8b1ddj2whfQ2IH9ZM8VptkSFPGesWEOnQoARVvwJEBjQ6OWxo3mwp5mWPuK7W9I6frvNuX6TqOLV
T95YVYp/dHq04V9G9USPuyiy5j0R03pTWthYR/T2pYRMfuFmx5wJaoZpp0W/JQbG7ii7qNcaacOF
2MF19I12+mgSiuKIsW+KFGv+JzFZja9D/DwNg9VNB6w2P52UbPvGw6rFAg+NaoS9AjWAvjglP7+A
8qH5Fre8KoE3AHLnt9Ge4tz0ua6q+jp1csiIz9aC2BqoWoXpR4MN3nL0yDWVTC6V9R2HsG6B/JIJ
/f75/bd6IgTgXjqpdRlfvAk4XmLog3/Ebncqfv/y4h0c18g+jyxYpeFG3rZrX+M335X/JZcLAUdU
Q82hVl+gJzTF3jO/qZEUl+6mUpG+mDalOM+LqYWnWXdwgNKgMgEf9PPjH3FbwT8/FXvzz7S/A4kx
BwfzbnI+soYEcpqtsTSlQvWekHQRwklPhvtuGkPbzEUjA8JFs5JN2pb8UMxphWhUA/ylhGQAnAVO
xvc3vQdIy3ctvM9ek4tVt2yI26OKKSy/X+ouzeevp79zvgIpD9mOo8xGEbC6aj9MIyq98PASNVfR
oIkq/gB6Gf5y8npx51LFgehrE1j8kO5lF40ddT2RqtViLZ0ZHt6Bi9fYlcUFY1Ar38oQrBPMSGka
FrTbSu7yW0Fkn2zaJAEMuUzDuHMfHQDGeRpPU4RfM7K/NaggBiGAzlNw4k9oMuaCf7ixSB5pdTlI
WHf6RvJKywbTAe5hRIdFSMCg2VhPso/7Hj2aniTaCN54s5/aAeq66Zb2vVI/OlhQFh/ipLHkxvQ8
31Cgxzf123FYZRqBRdDEg6OuNHDSxT6SaaJ9kyShNwh+3AnSZYN8lQP1j4ebKFvDy7Uu+fBRCh+N
gGV6PBv/5qbFgB5oLPRXRXCtnjBsPYBvWoptLis6pvx7s8J+rVVsJIwFu7ipjrWa4DWiq2GB9xAt
X//FUE841WhH9wKAYHQPiwPS3pbZPN89aQgUYPFT4sdz8I9mu/JiB8aCjGy2ShaX6/2NNJNmNsGp
AM0oX1hYbUKUbSE8ATO0xC5wV1z9+5QSUlM5qEmL/bFUxrKjdhh2S/owU0pIJ145QUZ+DsH0ILWa
M2WP0fdsmKmDC1Dxr8gyyjK/UZoePOGSAPl8k1ylA3ye5EhgYcERhe0DyfHv5Php6mfDGFBkWKVj
lRnJ2YFuiWmZ9a9G4UIu+W/r+apKKD5iarc67nMs7HKElJkH1HGIRMQOQS8u13jaUSU/yJ2BJhJs
eyuydIAEL6geLTmeq1qAdiEmoO2JCYlLzoSaXsUfbSLloxLVg6qgBXlg7EahzSP/INHpqCOK7Fiu
kOfvpckzCQ/CGaLAPFz5Br7MsrxCHLoRJHlZyX7+m3T0veHIAu8zE8bvIPMUOzGSP79JwWRBJcNu
bzVYvrhWWzlBV4KQuPdxkFhmte2jlxACjlxO48ZMS06Abm+7Zipba44+y9NRGkZGyPYSGK4muVFl
tTIy4+GMhAh7wq6AF33msrTKN9f85i++OjgXM2DqwJAYcNQp8WxBOUll/BrexglRKuoETTTEPHtc
q3jUvuMCzCODEdm9ny7t4+FkuJI8AoqPM3fIUh7inJ2DRBNSao/x16rn/8zHttjTrnY1NIJ0qzoA
SFfMtQEFS/mlnIbXeEgyOf1C1D0xcPYIsW4dY8zSmO9LQdiVKxKlR8vlbtl/Aw9CQ6ILy0kRbP7o
GHL1loTSotSCDuydErehdpREywlWt1iDk/lLnqxuGFgp0sWjH0JKa/Z64M7ZqJnWvN39lGvtmLu9
SzAXGyQxgszCSWx+iTMG82OnahKwA02DekAZfeQ6oRM2OxHoWlWnKGYyxEDZpQP3H1JercbM/Ai1
zKHiYiqwzM3PYbI75odE6Cvsjv3ns71yCOH/HVTSYxjGS4WmUddWxmVEynPejZhrPUVuGFeEF4D7
rHSdGDO6IDOzxnw5AUMm/44oZx5r663CAVYBwPvrdhoabL/CBZRL/9RPNgOFeyvZ0uSiCxenwPYJ
oe+n9B6TMpd7/VPBeQhgjDvl79RuYUre1vEah2UBbxQngOASQUHzC9EiUmsA5LMd4UyOjzf/TZug
y2UEpFKjhLuTFm+M75WsElHC2phU1bY/ihwifYGVp0jY+Fqn1D7TKqSGG789qEOJjDWNMeZWr8QT
1lNDXa0jeRdg2DYC6NhX3PhRtDdH0PZywkHjTrlRCKyJLf9L/dTPrfwW1kPkBpANi2CeoxoKDaZ5
w4aExrw3fPxpPWdZm9wHfZ6Ug/9p3I01qpslC4xnqJSq07SM6tFPNG3OtApkiP0uCW+tmpsOmFOp
7+hu+7cq3g53AeEYu7QeP1lEBsvq/+nbz5NFehCEw7aQOCmgg4Pu7J6sfb90VaRv3XJhBYfI3Qwt
sg9GkZva7U0LU1+3zIbG9Sf893K517mioHmpDVbcDZCuOwlI75Z6+J1urWddrMADiIIFtw8XcjE2
aU8o6rpUterUvdQ/3gqM34b/VlUkMRfcV5144s5w3agBG0DPsDiT7+RqG1W/dy0S4mc693W504Ms
KcywxMS85qhLTfamPrEXLclZYZduBhlZozxgm5PluhCX3z2MEKddKUtkqTwPY+kdcrfKUt6sLEAo
Q93mGNufo+YDs0ESlNKzdJPn1lgQyVLsKwJD6iRQ6b9MzaSkCFFYrQnsRXbuuWEKGr2tgLYrDGyF
c1V2W6Hu4dN7yh6KtBhWZt21SFDbIwhiWyXY7PgcuCy1Fa068AoY29NECOolxNWXOj1GhliEp8Pt
krvSppv5XK4ZtrhIbtAoeMieZCPLPPXUteiw/JeHtdzZgUsMiuF8eL4eBsbZFJMZ7KlQtHppQOV/
RbPBaRrgpblPpH65uKlXY0M7O+MuIsdLSrCogjqyEFdlntoSquyUn55jDg/Zddtm/uGWqQ6tTOZ/
cqkRaDpNdZyoKUqiVE+atNMhwCcFsQckVDOVFUSy+W+rrbMBAdyxda2Mr2SepPrThje1dZGVrwuR
KMO0zdpEM2sMSCn8zYp9TXo4k9HjQgn5lti0DrcpUPEfhytPxIH/0aD8KnPwZupyhYJ3jy9o9QsD
PFgfJRolhaMnhyNwrrV2VjOqWDQ9+ZzVO8YUgBcPar2zX6tQf3wJvkdvZodF2GwjuMoRD07KNNAx
T2HrRgMdIMOa6ukbLzMVfcWkv+TMCh9PMqF52g4eWErrquDDmkvNq5Smb3mIHWyKvnn69j2bfP7/
MWNwdQv2b+XEf4+k6CCzkxJGrxz9ecQ1p46JRGfBrk4imfJVtVw4weBCXfINjLhFWzxh1JnX7npU
UQElCozzT5750grQS/+YGwWrJdoGg2w4toqYH3yHCJKUa6DxkKJsHijsQcJGpX6WYVTaIJtGSfHj
/vr3L7ZRI6Co7m6+pJRk4fkbn6Rhn+qnBLY3NVagqXfmO0Et4RkmJpFaYoqbUsXuE/0AJR2zuTlB
r/U0eXI4Vaecp/Ccv2nnlpneQHYux4WRjCm6rukofKYfHoHpCCLhnk0bQKeJ39f+W9VtqJsMs+6e
8WAMBAgoAipC1aaW7BmHeJlkpaJp3OhfLBt5gW09DQI3p7BnRvHj3Qem9R442TO8O86GTz5a9sKc
MXxO+nLXMEwhtepSfJllGbdpMD+kBAri26j1xxjfbGdvKyjbGZK6r2FMDJ5ON4MRxR+POkgBuZt/
ci3fzlpG1NRBioO4cfu7ZmsLcWQC9Z6XNWe08EotF6p0Y7EKCUWzSiP+GGF2wPZog4t6bLrDb2ej
Ai89MY0yo6T58aI0D+LvJ2dWw03YYOq2sjxFeGed5A2kk/OCFK0M3o9zN650ZW+0UQHFoPj/VRJI
J5hXARYEJkwb3UggFVcLvDLOqRQNQ7dRcrUcES3WLVslHc6CXULTKCQ6qnAzADC+wxKLaW5t8l6B
zWCsSp19ZUbsRssu4/PptkBu4Knk74FGej81UZULLI/nNx3Ie38Hy/3XlrM1CDqTdB+JxiKLlS5y
/J8FjeZBoYMeRT0+qkfK18b9CVRZuLTm5bKU+98w5nlhTYB9WzhhbZngiv5NqQ8Xw23lWV2xkIjg
ztHxun0w975k4ytSHAOKxRK6VkrzsVz/2qrEJQATkQkNildtRhaEMSFWeOnwtcIlXaQBlSLbX7r6
uqPGidkIt3dkW+ynJD2HYMFwz3I2oRiUaq1TmpgWDDF7bjm6Ie2EsgF7gKh0aq2o5Obv2mMabxWK
/3wy9nw+slGVv4wx4yWK2Di9VIQ2VU5OdjwJ47+CI165RA5J5/y+RawA4yJOi3WoKmCo1TmXfm9s
26i6BjEsLjp+c3N208WWSRbYktYdC+Pab9/u6B4Y2+Xrcat0BFU9fNN3/r+kalU0WziJ0bSAzUgb
Y6wG+JX30M5gA835V1FohT4o1iGdC2yEX9CpJRstGek7Htg1INcrEW8twT4ykYtnJnZWC5rx8tuc
9Ipk0BU9cRz39XDADsABNibQSH1egC8AibBr0t26WuzbTdX5ycRWKaCaSoePQtgVcGsY+7FPu60Q
Aq7QNwDv2u/PlXo83c1fxmpCm02Fphyzt1K/vBtOFEftz60aXmvVUZktlOD1qSmUUxzYs75p4tdC
5bt4xMDogMAcqUq2eudFSERb+dr23iQ5WDELZncT99xPDJEOQHeL3nLdmWBzzz7RLb/8VIVWGjfv
TE9hmBxwo18CBlesVKK0hMrIKPE+VdytkMLb9vpIlcOC9NFpluhsmvzzmSf97HquSvNzKnYlgbRy
p41F7+kc8llLTRxZyMuVHCcMsXmLzs9vgFP/BqN7Iy65MZU+kXm3BhAxcbFsz5Uv26RY7PIh8L8e
8uJo/E66PRelzCiB4D++QVn0iLO6R0Q+QQTjXT2hzaCAUG3nAqg5vD7v2znedVxNOblEyH1ASswI
bBDGOo8HJqCCE+LhDgsAU36u1+h52jFac7v008dMejyT3NQBPYobCBbG1v8vkDl7hVVa4GFcYDHL
noOzeyi/2mOrcsRezic2bnxqKOrE63CK8nNDsK+lLOw1S1vpUWBZhNuE9I7+5Wq9RuCBpefo9NyQ
g9b/Zfuqsc2qQhVghCVAiZXTGUrFjgznbQ4/+36UiXTV712MQhRvvJ1JsZxBWCnWABVWc1YKOWfB
PiROJnw1aoekesaFi85IiIUGOLc7svrVfxTuXh1s9XlQjXumxhAfQ9opE8UuL806tKMvukDifRUq
eL2VpVhDPxme8Q2tDDwwTNAESdopltBpP2aoCTFa5t/GS2mxKYG8RuNcS8yVp4AvKdSG5YiVgQFK
TtXFR0IwjaZnyThBBDcTFOETsfm+ad7z7IUdPR1jrpkoZWs8IAqF8K3lRZEEuQOE1+C7Z7lJOe6c
iEb7tkqgi1ZtlyT+eVzpVXOBMyljqmZqa34ovPN7wXvfuXmyrs3wE2MfWoAJv6bKsIxGEhHEduGi
W5pXLi4FEFsZqb9j8xYyBiPwMENHNE62URaL5D1fctBK+gvoAQ9a4KLnNVS2ZQrds2rqUZiBCS7+
misYTj+eOxnNdRT0sOWETHmleN+aMziJzkHDOAbHHs2k81+1VyLhlFX8NOmmYDZv3g/NppCXTZKB
Q8Dtu7lLzL2BZVUSTibj3Rw8jlTB5vtGTVSrjE01eJ86PuB7nB5eK7tcSnJYtUhaHtRxyrwBxPuD
IuajcF2ApXyG+ZPL+tlRWQDbYZk7Jne9E/45YvoQkTgrDZ1cGSCec+cp+3yswVTpFuxzrnG2GBzX
NeHSYdetl7ILs6UL/JVgr0vETFLp0X/kw2jkWyR9YjSncYWeqTMycezXMxHbl95IFW59TaC6ACRy
IeYSngKhwyVLoKtJb3nTd9XcG1LHZgioBAonw72vxXwms1Ea9zzR2vDogWknrZ67VHhlG9gBNGZr
EYYI8MXEiisxps4ZGxveXlBX9PLw6P3CmHTGN76ouxCDmloARGER0AAFnsItokxGPymzdu3S+SDl
veY6Byu58gaHc0NoqdNKLyDwR1m7IM3U4LZhcljMQuKRNFkz8eESg6KoVFJxJsXgRHzVHGlqFCPd
6PBFS+Br+XobBisfAxaUKSpdYKwrL+abD5bbfYDRPyfawUrZArOyuD0XtEM8P/fzayqkStmzk2N8
/EXLpJGj5RyrV6yD7zUn0AWWjT2Q0tPC/6BgWIWil0NdcEy8BLcTLsAxQqU1Db4/Gksd7BRp/I44
bkyGK+dx6hBGGLQUlx/ovPV/aaef8efiyKhDDCWCddM+xYRMRsj06CEFV9yZlPcwwlk0dKUtE6lT
Js5sTDlErqNtLHV1IEeNlej8Cj2cyEf65fUAY+W9kEEBA6QLFA4S8Q84tGAX14TeeRH2Z8r6/Zsz
VL9nxrhC+bDkTA6JQKk+mmQeifD4AVw3ryuhEpMeEgxdS8okuwZxz3PrDBtiPYvcTGlh/ytceM2A
RnpeYS6Rh1R9npp1f3F39gEZEyGsdJAYoztMe8jPn5s1qUYmnkzBjvFbwhqrIXKggCNLrOI2vA34
mYIaB9qr+7EOJ8nLzdSmXKkm4k6NSsbdA8yPzIpYA+qBV9KzOEK6CN/S2vH+rhfNRWQY8VlQBSi/
C6EXtKNncgXZfwjIl9XEX2x8nB7GQEYjyI3g3h40kV/Hn1GZxbBhMW3xdtbv8XkO6bCTJwOwg777
sLJfphn8MH1G5iu0DGUUCjFSJI/uZYfHGJh8qPJvTi5frJ+y+VfLS44lrwkrUjRTOADI6xSTevxF
FGspFfzPcPhWAuKITIMhakz0ybTJrwRPMAcmpVhvLV/ZbfQ6xO9FPhEdixNfgsMJntoYcHVz7DIa
eLMLus5GxCA7Rca1dPmYbClyfIyct5CAZ6OldhsfKH1AnHS+Mh1e+6l3ieYy2wN9GV+R8t9snpmj
QW/tQ08qLjUtJOxgjBbqZj6mtE6+gA1tHQuripl09V/R4IroaU1FMb9a966EPaNwk52WRnP1xOFQ
YvbIsy+1Ity1SKqUPAqSrGJ6oMeL+EH42DnSGa6zh6fwCs1eMvS2rbyHYw9D1KkJbd2uiN8tADR0
Irm6sww7rcQE3hxhsum0Xzz/hJyCrWA2gqqpJ1JzXDqmzqx2f3TQZv+wh0QZMeNGM2KU6nGqfyFN
DEiqiQejFFNmODHT2tpkqCmKFqJeW9Umb/qZIKB/0Bfh5WWJmh+wughICwR5W9zbTFNo3zrnd6o5
jLKmo5ATjzhEBkpMMzWDJflo8hr1AYVhRp9VorAaQPP03kpSc7KC4k6n0zXz33cvAeA7yhOvbdmt
5OEHJcuKxfxF8FH9CMbgAMQRo3T+TL228/D52S7JpdvHVUr59WUZmZw3/A8VUVCqyj3rYy0/lHGO
MNW4yu+D3SC9MGBlXnfCPywHDmaUOq+9LUTE5Fnop3OQRGcq18DIxlxQJ9t/HYEGpgFOaRtrS5fL
N8omK6+7aBAv9tD9ZzNWOT29MLXDrMANDUqQCroJUpZF6NE9yo7nfZEqpBIpnkhP0d0ez4HgdcPe
AH0KzyrDV/w5acgvFJ2ANKT8nJBu+fhJCOPbLtiRgZnJCeMnTED+ufC98bDDObzDqHt02xCNBm6T
zZSeNRaRAdDqmxsnX0cEy8m1NJREXOdVCbJZlzBHMAmw/ruTwPpS3b63FOXUaAM1m+fo7VKOdr1G
VRxvWNU4n856ZB1p196v1v6T5SkGfkMWMbGO9EQ2WV1oniPGdf7by/J1/4v0bEbOumhz8O61VZww
zZ45M7RmxMSECUC2fbAdvF7HgdGuhddpb8TM+UzwDXXwQxx93jZioK79dwWSUieeSf8IX5kRkr05
TY22tcwG1uNRW4cvAEP1dohYaVlvMeoUrs8XEV8bwRh+LBls2AZ4sXbM0hewR+sfwQP5q4Bs3WUF
O5KiCxuZB0BStQOIi7Y0SJNhNfOFsoNXVQkatoWlMxrm2a6xYmycq1nZMgXsIwxkigEsK3O7kYdH
WrToUExjHFxkYGPGXR2KkUzL05yw2PpYzG5zn2KaXMwtanhM2b7tIFcRQgYgsg1a8/vjRScJaaiH
qZZgAOLZOpz9vCK5nxb1Rh8KsaRY/GBBY2JZ+WHJeXglgq/xMlq3ObFjFhtTcAuVk9GZYVosIq7K
MDZ2U4Tfz8stEyAGbOsWCwU3sjAWNNp35nGHvVTBpYA/bABcmGGizmnANJfNNnULGb3+V93WU92X
gnk0vonmoZlMAtUSsYr/AC8hMSFKr8qJc6XJzeFxhU+zKO6GflX7wDaxWg4Nt5sRv6rVYjS8fg56
lp/PdKwNwTROd6JggxGyiwDiBNJgq0FeGI9viwUvYLcM3dlZUO/agv1AjqechaDkYhX4uPq2Gl24
N6GR+OYhZWFuwWEzGdRwcO7LWlsvGSQTYutTML8SHCkAZiLqdRCK9L3mpEy55+LABiV+fkBN9mEZ
Fjs1Sn1cFkCMnA/2omTgmKEOSdKT8HhiraTSsKFx8N1VbbYrl7KpVFkLaSdWgZFhkvDW3sDmSCXT
BopNgOtE9RRrZc8UxD4JkOF/ao3abiY984Kx9Wl/vHHeGFMi3c9AmiLHNc75ErvWB9zijwxamPMi
MhCHvCjW1PYBZKi4YfIoPb3qJ/2C6hMFmKK9k3vd0MiGXfvOrTK7hGFN2E9A9z9OraweyfDVc5Bm
HQzyGC3jguGgnf9w/fuJWGuW6LM/1iPN2IQs4E4CRa40yeM6inUuao+uspMgv8u4fwR5FNLu3sok
/Hq//ZWqtXsa6oN4KWaEbKndIPdGVEB3AfkJ8bmOytS7rp7utAdVArFyY5kglhIM8ugxmXHOjRzn
SfGeAUGPBiBKsmvpzvAE/WTGlWRfOF6WIzuk62g9yNrmkMTqbRxJLLBHFs5k0W2kvk/S9VyxxuN6
GG1ofWNmFIPqOhDwL6wstRV9OOGbMJP1AckQ56r5HHZbwPXrF+vLRZk0CKd7hv70h+CBg7LQxSBW
ix68Hp813jaNt9kcYQfOg5DcHaZnVApKUOhi9nlHWcAnb083QVJhrLGBG1oHO5zt+TzgSqFE2mMi
FV819enjabIawyLbrim9m+ZhioC/S7hxYqv8llrZwSKiWisNDI+oNhh6aifTVKb/tkJEj620lfQE
EpAeuK/GUKkr9Y1C03go7lCM+PsQ1nllpsANT/L8zB1i58cM0lYyZ/Tto0XKRl9axLZp7BJM1J8U
HuXJZ0vuvHs9nBSctrv1pzafvLDwV7Z026qPKq1LcOkoeTUZal/PlDOEDfSP3AdNlZM5d2lBZyhw
FEBgcnftgKoIyVSXCo/0abXHJWgM10BXOA6UeLIgpzgfnoB2sBLWWVSzkKaYfNATUJmsS/EkaZmP
9oi1uz54W/PjVLtqeK5dH83dae5ZdrQTHhL4sB23vFT27WIoKAMNLRKtU7oexCZcXC5UxPOiSfZO
pyDgWIXSxp5DqUQ4mteIHll2KrP2KHDJ+JpeldiMh8GkY7HDCmtAl8V6JpRCnUX1exJNzUi1PopI
rtxlql8u4boH0OkeglI052ZgwM0lvmYxVSeEDLq1jRziOnLCqas3mnubrOwRvWNV9GofS4/t70k8
k6k3nRplIz740svELeaSUgZ5XgDr7bkzlauce1p9s+lDPZoyl5NXCwAWzNO25czrcPSrKWwLsFPh
Q43hLqjJJBpPzD+NE6L3wz0xyrUwOWgshNjA5CE+d8kvgqFScmjN10dkNmNE+m5yuB5kr/BeQIlW
kaCDTEfYbZhAl9NDtSDpRK36j5bZzIlxXlEtICox71Y4whbNxkwaE8v0QpwR9nxqSpYSYiccACzc
Q1/bK8Y3VJ8/aPGxn6jLzyK6pn7T0mb7G/HBlTxJmyCaV9jUfJLHm9zw3RQAk4D+F+pxLA0hU/ZT
pgdxveKMaer8HFZxXVczRPkaCS/qgFw3Z38Aj67qkm8gSlUxmiT6NtiW3w/RU8Hwt6aXHlMA70oj
WDXxUIPTw++OtjFCyaEL5LHDuEyY3W2f/BhqDy3zzKGZRYjjEQql3JkPzIIGhoS7glWuVWhnDnLL
98G2KDGzwCXiCT+6Zsx9axpKX0dNcCa37t9kggC9BB+Ct0qOHT6H+aLn4oOsNKoHbUTmB6n/rUAE
oBdQBA19Y7DkJWdwHafNQ06LoGtHxUc/hpppViwOcqB/9LCo4LUtRfba7rQnW//Bk36BrrzjMApS
5pGkk/PVevvwAnK7OIVGc6knXDoM3T2ibLYU9sx3R730yvvIzpti0ydZ4vtuNObc6VQNqWCAdxvh
Ek83xT3cVFI8sh077kjwkaWh46OFmcsME7IBhcPc362o1YrNK8Fbne5FdqhnurFbP6GmzF0/SAAG
C0YsggEpP8xDR1vCmQh3Bst1X4UKIABSuNWqueIFYuTbefoYIjh0/psbIrtKShoEe9f0B5+PZ6of
pNzK0SDN43tiVNo8IdRamwq7FaSYxo5kRFKVEtwFp/r9kSWUQUkW9khx1+iXeG+jce+c2U6lJufj
K7sOuX8lmrOROnrkn609h3YEkM8g29k4gYB+bmipQ0IfZsbDnKNY741iaSetMtiqX1Ldxusk3iat
lpL2km1q9lsn3Vf4ae9gONIj+loIlABWusUJAutmBhpisJNPk3ZJaJ+c7jR+nQSNiLtbtJQo10am
z9fK2iS+dA9TsRFXkzuCDRNfic+Hp3n8hX28NJ7JYCyMsjWJWmvRt6TZ6qEtPTVihlwloc89/W9p
vnowc/gVluDu/WAzpUXwaY8gl2Q3NtDoYLKGifuCouvQzOZU/uKjqv+7IMNWU9an1A28JWwsPGQ/
h2qOxJTsN2bITz6zhDC+YHt7TzbY7qPXTkzoYf3KUjpq5t074e0kgQ8VfmTF4Psz5h9uTqNzfCbz
uRKSB2yaQ8brhNLB8V5UKHLm+jCVuQTqa2RasmNBsIWcRIx/28XxQUd5rgyeYMgTA4bDNJ1HLAEr
41SyV0V7K1AhSKwqh4czUB2mx4cOKvommf1+uH/gNiTpO9gpbtLRZBMDBtFIIMZV0IT3UTY7/BJu
pcikSQkJfzPqm+5mBViB8Gx88a0BPVkHwoM5Q8mWgdD1AMykkq6F83bnlvPTve84pfeP8/9hp2Nr
bCybg3MTRzitiw+KJrU6Ysl9x7CMRjcZOsIXKhWXTbvGzcvtjIEzShtckc3R5YaEUAA4Su13BW6q
MPDylYHye2Ek0h3cMoYkihShYVhGs/QYY2HnT/zXCm2HHpQugW9vdt0QFfwz7bllcAhhI0MJXsRJ
WaFFgiHKLYT63pbFMioCLZIdxAOxm2tM7xWMqkcGqlxOvuF8JzQA+AMMjZSVRNuEf3ZKUDZ8jmk8
nUgItU05vBEtD/8ylaCmFiW+sfPdbTVZ4yorISU2EVeTc9CjhNaCDzl0rcQ5V3ulBAzZoDEmz8V7
vPWVGMY0Uj81bDfVWhTSNjJ7zyXx7NCbIxghbecA6ns8LPDaVxOPb4J8mOpSL8n03f18kflYPJgm
yKJ+a0VCXqtf6lIZW7W3ZbDiOgUw/T3yC5KSDEzZaKy+wHfyZZ9zyY42jWQsUNeg8JYq2BDCIAtw
Fsdbg3urgp19qVz29enL0YdQwIL+H2bEYszWjlMJAaRC4JoOhNyYlJTXCYFn7ZpKU0flFgYOLLl+
9qyjc+EU9oshZ6Wczlf0g850aaXP8I5uO5jX5i/HGopTL5U137gNeI0WRAgh4CXQnqUWNfBZfKcQ
T8QXURQZDOza1icQfIuw0WvTaUm7MTgOcNGkBcRj4tfXqUFOaVlgxX4GKnjSUQWUw8e0es+jx/US
6fXTiH+jvLth+Lb5xRM/aL4NfrQxhVtSH5uX80kDSB3aYYeD21HrNTemRQLw9weonbFyS58G2NTI
ebGqXhfg4R0BoAIToINg3tv+qmjkXg363cvIJ8tquwguQvyFvbni8yKiJB+QHi6wIkZiJw8muT8c
8tcOR1cNqJHuhhqgOff2EFcrwelTvgyt08rf3xTyWqykB+gvu4niQkolviWbD/C+YvaKFOD2GcO1
Nn4dS9Xby2fiGR/+dJEgwcoA3TyNwfCKrqFK27GZ0a+Wc118+ot7/ef9wQsLoOcO63KtpycJiOsd
3nGydeBerthv7633qxiZUhs/F6nN6EBh319NYNBbGAxF946OVDcwNS1H7yt7OCED0BxD6jCiBnGG
c7DiFkdAqrki3Htcim2x8AKjHfyZsN5B3cFtBfqqj0JEzLk4746F0yI7drdEvyaBSh+j5dmlr3le
KSVskE12NDRgEBPUSfGRZnQPxV9LqVvg+E1XIFXMqgoFg7evbJtnGV28wC3q2jwvCt7NDeU6LY6U
GPCP3VnnTOFOY2Sqfv9lCn76t6fBaawKfryVs1ylzzqX+8SARRRpBUCGpfwJa08awhHILWpXUglH
7ftWm2kfeq16YCWwJqrwKTF7BsG62THqh1NBc4EYZDsZyMO6K9nfwW8ffUR4akMLuYMWU5xY5QfS
5LdvTzSSpfRZuSCqh0MhCpL3bOmXhAtPGdZu/Xy0nFXvjTT4d+Fl0wEXWqoorQgbMSZbw2/FkuZZ
95qM+X6VFhrqkWdMuDH5EbfQlsKlnEIGROY+OvwrtAM7/MMCsUqV2PX7IhOR/aiO3OA6PCaAvIDZ
zFp7AKbQSlLATJ/1oIv6EmE1jnGd4A9uUOxlquBxQ5nVzYRwjSu7FSjt4gVGf7LV6FiZJdJnatrB
TI3itPAHX48CUEGe7ln6Aso7e1PaAI+q3K0b6CAzvaFIHC5g2vbKX4dYvXW1ztOEy9/wyQ6zGNKS
/RZOm0mLiuX/fctakDLp/1M2/LiOSFvgYWpHzNsJlfkUD2kGBUmdlgxd+t3f/OJ0ycxF41jp1DpI
eWHC6WrJmIMWF1xZI1dwJL6fhlBt/DNQg05wXhG1ni1iwVU7a4CNnqGw+N9YmW2N8NjutSl2WyVq
IiEBHQV5CzvQ83Zqn9Cq3eu4X+g+qMgTDswzS8vyLQoMYc13D6O+iptuTAdEnxNaRCD/tsy6PqmD
LKGf4+5OdX181mLH77+O5L9Iiu72pjMM+/Tynx1SX5XndVZbMoGT2gN7TjOjYnfadxbEIBKSyAKQ
4LtQom3BMFw9dcXUlBgfwh2Yzx126O7ekA8g49LzvTdxbz81ykTznC+lGFgw2qQ4mSI29WZaNXZy
CQ1bxknRgWmJ5RDQWzE6Uh+u8Q/euKsEqPLJz2Zg4jbdcvYznFsdwT3nB3Q40xbisC05ebLda4Ys
FVJ8+m6rQka56Fuhs81kMJnkyKoGEHbG7EuxgcsOsgHZMy+shH9oK7TA81Xw6IOOavv49vq+75XV
5UPbI0W8Nb2GY+1kN83nh9R/8wK7tJs7Vzu2Jul2tl3yKAR2exIH3eHA5P+aOFKfqv7N0fIH6Dg/
P7cpLy6cRYPQdPWYNvB6mHFJQEI5Xo6TAfZwbLd9k4D/DVNCg7Y1kgirHr3n6pzbMRnB/kjl8GS2
eRm/JJ8xug2IuumQ+kceMEC9iTsculh923Ly9XsWr4NjFlJgR3hx0YOeNNGOmMTM+u/ryi17hrs1
79bQ+eP3AqOraf498lagwMmNq+nAN9MayzG9d2nWC8/nKTn9kxvlqmwHUyspNzT7qXWpq5+CDCvo
X3LPDJaIlcv4x5G+wEy2fPIuh5MNp0s1SqvnBI6Ml+R9G5RFpB0aV8rAq4JP8GOltj3A2DrsUTXs
jjS6SxGbZDOlZmE4rfGHgpV4MqmeP2EF8iqi4XeQ03pWwPdTGj0xBEzsOuKKLyTOvuZ4HtZ8a5AZ
9Iv7eyBy0DuW40r7nHgAD9glraNqRbmirqBr60UZC1m11USjb9Jvikt8GmBGDgYAztBxc4AVu/Dv
JdNcv42r22ONv9/JB5o+3RTkyqZrxWSJMfEmDhSBEl7gM4ydK6RD6Llj51n+Ri9InCjFPSEkGAsc
hwRbN7WIpb1uL2R2Rv0PBSgXnOoUpI7RW2sH0x/Jsx3B+Jr9ZaCI2bATjqweuUE8n4b8nooTSaNz
e/l5K/rr59M/6/Wwz5kcKbx8J7Ao2m0zfXn0ZqzcoKEYIF7ojyiA9gFKprQ5wCys4nc4cw7RCByR
oAmO1net8F1QgN0s++vmWaRvkDsJypfyLFa4c258qo/PewDCrnrehNmy9hn8YnMiyMWmS8Ic11Sz
DjSL2ArRenycjzdUBLv5vHbJwfZjIALXEEH9xsNDZaHpzqb7C+tOO8NVWWqdBMnJQnM9vfEFT5XM
lYWhEdyZ5IRnKErvi2t2FEDuILa1rjlR3S/HJwAgwlUOH4rJGT5VoV+UDwm2WQh/C6Dw8c5TDFuo
AFqavd2lT8oz9C3EzShW1zjWvzNl48J8edYxn9CULPJRxHL3aq5We5htXn2Mjtg7WnHflhDKtu7S
TCmmuX/gkvmqANptXSiEaGxlry5pApJvc8IMJLHiU2yrZof7Zs4Gz8oHvPoKIz6NqMJ4oH2dc0uu
hgTzI3jQ8civySyW2NdDct/ZE/HjPF41YqDMIdSce1vEQYIJ9tyda+vCH9nMlql+hGAx3rj0Qohm
RpDr9Q6pkMbGTyXdLuY0eLcucUSqVtrAPQx0aqc8madMwcv8Op1nrVOAbF7RqGgIdzWYDibJQON6
9oeKsX4a+8LyEQBLSUVxBMEDi9fqQ7NspYrrdcNixfBcelZkHII6g8thp8urzH0gmLfbaf8v3CGS
aCYNDtS+DZ1OSEha1orkAd85P5+HdU2jbhi6r4zgaAM1o2A92YY8FQB7BpuTGkUb7uHj2faBFc06
uRTlrdOVc303bya+YtLBkl0EOUNy8tOJ1Hz9Ne8l+7s3F08bMMgl4R3thEmQ1bO2o3NvyZO2P4U+
BgZr7o3yQKlm7CN0RTCzBDLM2Hgt3TfJQ0OiVIOeRh/1hUVXToRrQSaOYQtdEL6c5Dum0c3QbJlO
YkTucE2J7sQMQRbQqLnJCOFKOYfv1u0ijTaQGt+2vS1XquSE91olZfke3dV8zkMXuVXj4T0JQMNw
62OH/Pyg40Nauy/vvuYddmh61J1GGMpqyFo9LH0pTjSEKAHHYMQk9GKcgtHC5yJ+friYvJZdKmWl
uf4g9Jl7p3117WQZ26VyVHJLQa+orxD71Is8DOZizYkXFnoVfRNCWPNLN+ndxcLxrdArFg5wwj4T
Ghi4jOitIqvGvbzcrpX+hj5rQK1eJSM/j9bBY1XygmMNBK5crr+aS/bv1ovFzzWwYmgtIguYUrZj
fBYdhljm41HguH+VQqb/8AN76PnvlJyCoFGUnmd+Di5Zb4cuKBP3V6m8p8s3qzWYaG68PXX2P7Ie
bVWDvh81fke4WRiY0NqIePNRkBY32zuXn5UhmobtZJjuxvIOyZuFPaO8iqK9AQrRVm7BbaTqemFh
J92NXH9Qj54OuMf9fN7KejBYksylrzfykI92/blJKu6YzfOvQ+1g1GdbDUI6axYJ0/M1Dqm6LZOa
RwZD7MO2JBsEVXQyvpf16x0rsjk1qK8lUuRYUKimxp4MOvcfIn1YmYTsmLSuqCsrZt3E1YN1Ktbf
m8OUuBnxkrrc77SyDW/LtejcJi4TzorZ2CNKtjyjT1WF+jzHmL29s8orp/f6crnyg1HZ4TJEnLG7
nLqnsnW+ysuG8iK3Y/lHgekEcxRIMPTbBC77NWnSpd8bchARsQyjSKzZOkzKz0EwnZGIc9QnT7Ml
IdEnfhY5YEezi+JNS4ZuU720+Nhytv4x/N+1xP5mnGxtteBe+2xSoFMaWj+gVOs0Mg0Y3+CGZbH8
cbVivo0r3GDmhVgKjPhvJ+avMzKwRnTHWQVGhAkhJKaxX3Rz9dtwdlsyk2oQjOwFxc4M1PR7J/Nr
Qw9jrja/06AbBKljvgvHUqyWqAh668Fca2CedDuSQL8hlSth8Z9RAZ1/HV5eyhUYzPce1KyFBxJT
imgbkgTurRJ8QVFUEm/ZyS1cRSzZfwB3U1rJJ6xZ6Q/yUA4ksZZf5XnYdvAhqmRZWphTkfPZFFUZ
vim8OAFA1SUp2fiqSdQ6JwNIQvp2nPjbSyaiJoYh8cBrT6ffbOgaCgLqk81UfxQDkH89Soh+IWh+
qN2fIMGB9uCwBH/UNscL+jQSLxNbi1xKgZF3uy6joGZ5I63GsfSiGkS66ZMs7LhfoE/N0KIoXI7U
AC18owK1tZS3ZYhgB+5b5dc1n6tb9UDKBkb28JO+bbdfG70YIhskeSAcDGrESLMH8B+LZNKA4pEQ
5KcmuBpCVBKnabZ7dODrCum40DNUgXZ3BvJlWQc0/ZDetWrWfrHOl83Q4O9gKrvBd53WJobkyIev
/JWr4t4K8Nh061DVbtCGdBkAJGmLbtZMZQCsf4ClvWUluMHx1ESucd783axIfWdiEKJe/Eq9GRVI
7dsYTglCIw9Uick+eQGu7zclm+2UjeObdmtpdzTzD39nJyawwXDvxm7LoF/2UnpHFZcxmhZNnjm+
/m7KZi0iwsmsN3Hn/FV4lc2rxBuR7X/GfufSBer71adVRwuamjPtk0FpqXz12ZsdjD3VewkEcU/l
d2N32JuOjVcbX3DdWZRe4+FvZM5RnQQy5gcapQ0jZUwGDbkdtjuN1Axz5/lvoPX5NbFUi+xIY8V2
dtupQJU46/CWJ4P5+URAG3eGEo2/HCWGqZB1DDD1dx9YsCSzPg0FT3Y63/aJSmo/tjUrsUDh18PC
f0y2wPXPgqkjqobekuDyUBQR4LYLPMeWmEtsnknprXc/8Q/4LtFzxBScDtUYVD3lnR8PBjrBZ7Zk
bq0M+b4nyJA3z1+u8z6ITn/gUTcyF0iIt49x90zhBjFV2KScsGPGmvG9+sIVCNJuF6bmQR5JIUh6
HJOR6TVbBBa7/WcstMyctwaYdMJtpzxBILit5bnphO96QulJGdADSRYXLXgC5ahBzh/WNHTXQX4e
RSvFQvBDjbU02GFfim1SZ5wdORx7eJptLAvgMlKknol0wzlWFczUv1wu5ewUKvL6FgNCPCzsolLj
EbIA1wmsqCR/ecOHs0Gb3GXhhjCVzqe3JNH1xryIbjoPBxuEV1+xO1uSuHoimjIHlvrh73Wz4E1M
clRWjt4MykYFC6QoFppjEt6uwrh/ZnsnCdmQ/vghkzUQPSjpnlWE99QZG6oUsZMUpPe2fTWcV5Ft
Rxyry3lcUAXI3MrLcmzqUUtOYTwvkaWVHV/Lgii/v9A1md8SHgZd6fM2sjaBPoxOrjtzqZb3cPq2
JFcWsacHj5qG9c4zJRYF01YqtzfgKvLMBeIQKh7wEwlvv0c3Nt1a6MZC1b8l+rhon95yjSCXOKtM
jFSTiaPawR7MUY8wSgdE909/P2aVnKAUx3KklUMo5HXs+zoXgZydXTYMAVl7OA04pTCPV6BHvsgW
NFLSLnUe7/+6JSO+A4WFZZz044H3eRB1DGczozmE3VXratojRXsdT8lSlM/Hb6hPPwh2mg7urQ8p
UcXXJupR5IiamEoEvD1zEbGJmd7GfdXFVe4z0NUAMLwu7OmMl+u7Af0sk1B3qu1FxE6l/r8sPw1p
AA1NNHeX6QKzpk8hAl5k02tPtw9YT8DxJeG8Bhj28hHE+Qw9tBZtpLepxpY4mZK5FF0bPGTdBClH
j6AgEOww+q4eEcqGXF7t9zOS1DR+yWdxknRQ5DCDwI+yp+pjBBIvYWZ+GU5pzZyzwG4t1a8c08mS
A/dCUKubML2QzMJzWNSmzkr7FPot2JFAAGoX2pBrUqB5XxJNJjHGKHqcCdVCw4U6EofPmtXo1zxn
IOG2TWehcDsthishgKEN9ezSankZdLzWL3G1vUFafV8stX2Q4LbIgpNn2yCW0SywFapjzLykJx1c
yaUQ9yVyap+KxElPWIv9ZXEHqpzsY48JNgZuBpDq2CjIdNU1TqeyDRmM2uhPFdtQrsrmO1JEFfnh
fyCFxBRO5gP91EieZLW6KVI3zQqhLBHO2VWJijT/0cXjjpfNTyJQe0wu+uyfRst5ANsZ6ve16dJE
eloYXmdosoz5613j+YySV+A29N1lAQU+1sFEBgUX65zI81bE1ltfje2n6DzVz1OtUZTaT+oeTJpN
28gZSEi451UPwLMClIFrcNiN/BZRmZC5HEvDBiR9foWWMzUJ8rt+4w8LOeMigqrlbSpEFrjD3d68
q0uITm91oOYcASQZcFsQFMJ/cWHe7NyYJm/++5r9V9KPLMtoQSDxrUDHUlXojGSjytFhpiiZ7Ke2
98DHfca8njIwc0ytmXOIurpO1JH4SpNQZeU8W2/41lfjHV+E7DTa+oToeyhGE6SoeEXdohNOGDZu
OxQzTSCn6onBEiZrffNjPAWQLhfz/zkYQBMJAIk5tJTmpv+5T8vJY1edNVivt9PaPUuj7PHl0egc
ivLnp5Sa4rOZ/UcaMXwNyyO/zPQgaUSpehP6FsTWOFXBviatgTEuWKkZS4XYxODqyITpxF+Q83eq
Y5a1okKG4JuchGlHktByy9EIEb1+6hIZ3yt+RupZi7emaE8LpOM0O22hU8CvXaNPnAlniC+Q78/Q
/9RBIXaxi52Jflh1tW0y4O9i1Ey2c8IjiYPLJvQv0h9raXM5vpJeLElhXwm9AtmJ0ei5Jgs1Rj7c
k90cxx2bCCj/nHGtVABM3Mji7WlVhRkly6vrRgO9ElhEBJNi9RLenvVmmNPA+WUvGSAuhLFK6Bz7
qW6h1JbHoXVdL4AqGb0pWxHMbKY8pkrTnKLm8dUNQGc3/Vgp9y71OThxB+hj6JwlyEERkJoXR39e
9BCRIN8KiCAR+n7Nr5UkyIb82nCh0QKNEAES9orECdlvqwXTLRiDcCTjt6SxJ/Yy5PvAnIVr0cIc
Z3jaPuRkM8NdgONXWvKjeW/QEL9vpBni4FYuSSvaW2pJV/cRTMeZnddnDZGh5DkpDf8iFeDUXT7T
bYz9YVW/CqrbaNiJy7SbgS+6lLtfxqe1K/hXQTHLWxRWpLOD4CINRzmB/paEY7WXXdt3aFgPCh9O
Z2Kqg/tGcK+njparnTtjQhyA6WLpWrUJdi195HkiV/iFxD262ue0RH64dwEwJv1ubsjfIsZU6NpJ
0sZMoTYeP6NHcoxdWDVGVqnszmZHNi1uDeS7UlSDR6LBT473XBaEdhfSqMStXbR+ZAFvZEKxQ8/g
L5hRgRON7dCvnKMxUu4shk5R+XLlx2w0MkG0mN8oovXt646Vm9QX5bDT9Wq1hlIOboovxsVAdTTT
QFQ6hWgY7JQVxrxsaucicZLMHEPEKs45Gxwdu8mXiP2CVO37Wl9cL1i/iMnMn+Xn5UcYxsfbwSwE
a5Y8PAZN3beeGhnf/4ARBId0NqduMkFJNxFxKTAygwpswTCOCQc2ILRvwR/uSpYWQocTgjJJB1vS
nSlZi8WdAEh5+Tb10AhBwhbkuJ9/aTYgGvSETIUR8Ap2CkckyP8PUUZOehrMm5kLlmWC41E4Ojf1
FUSB2FmuKRZFs1Az3x7ngyJnEUL2mbYSo58zJXhH/06gtQL9xJCcHpFKBm6ZZxIkB18SFZ3PDJwP
dQ8NoKq9pZ98APA2Gns3FrpD45q7x7XaRj3gmRCwf7nwDHVPOHxVfC3Dykbmzw15RDKPxI3rfAbk
0ulaFGevVcSxfBJhAEGgD5xrInPjDp78VT+2XYDy+iFqlJ/PsJJx5ZPD+kDsBEHW2EmL9iW2y2Lt
uHHqc0ahG2+KfxLhFwN5xBxxjOJCLsSTapy9ZWeP4b4f06llzqq3OQeK8lUNkUVbrBp876JCuvXT
djcgl4OyW54hU6jKMRr44jfbcCBXmSFLnNBWA4oz8ULyDyNBZ29qLQjNGe6VSEfv67rDpOInaBDT
L4jXDhuRlf4PsQh0aDztcuarKwVUL4cef7UkdMD/nhDVQfnigUhZNR82SGYWesdcJD98yYSBe+PF
WTyGjekVDj6T4J0lZymc2JUl4IBjSomRNgCwbiADte74v5QHBxfmvnDJH99J2as5Sf0jWMp7ekE8
rJztRkS1oPuHUpSVpZiTbUsGdsFiTft8S/dwBmHpIbzYyH4n1zVbtiK9rcqmP8iOR/s56QGZByth
xdp+szh6JLGMBSuO2t+JLCdsnJ05R9OloZGpMfD2rEkeSUM/2cxvzxDctYvZ11zALLONOr8HZQH9
kMXqGCtxkzFsJ3tsxyC0AGq9jcMOENs4DEOZGX5nQA5UZkyOPX5OXNkoAQOQYVxA+ZIAmBZWLk9L
//qohpLntdDj3rpwjcRo2Osh6+Ezmz2scVJpASu8evadoLOlE8fRGlZpwDkEMvrOW2GnTCGPaAjf
1NBxd9oVlDKPKPvq088LxhDQEwmxVd9wOJHZMsNx1tVy6U8Heu3bUezr/wzw7tsAX7WPIzyS8OE+
cx2p5eMvRNPemp50ynYGhxGsVXXoFzM4mcnRWhlQz0PxX6MVTK/0/S8+PXThxLYWnGNTdThXMuXw
gyrkGykCfEFZ3TMH8rYpkVQBKV5nYmVxAqMrigYCM9Hs521kZIzoMlCENtzHusaBoSJu/X5lG9id
AK1IzpyDZJiu3BunfDg9BdiFJ0UWMHl5zRIrNHs3LffYgGf1WHxikY2y5oDGFxf3o1LEmCF1SFMm
xy6yDUi+FqTuA0inlCi7jfl+vZBW1zkrfjV2dNpd2fmRG0C/GahboG4fPg8CycA+HsipHOlivOsr
ILNFnC3mk33SjjSDIwAY3BISW43q9tYs11XNcwah9mvTx1Z3/hVaunbeJNUH1Olj3SEilfhQcukm
jEcHB3YvlcqA7Om186boWnRv5AnqNSF1zFuQli8JgQiG5t/X6d+oKtMdA4RnV7F6EFCzo2bGqPIO
dnJLqAWLC2zH2bHTHoPm9FzCupZ4HXsiFIaWevBfEhUZzRawrzsuhMfQMMq+Sp2JZvY9lL/l1md9
QQfuGlKRGePhpG19HS7o9cgiyJEQU6f6o0dkdVNA+0D2D5JWgXDyKNcmK4+g3CRgStxLT4Je3zzY
KnHmB43/BDzfFH8eKx+eeWxpEOd7bgBQzC8sTLM+4lvL+5bhTeBYu37MEK6I2/MR44/a4xe09vlH
D8okuVz+dA7hB5ghLms1GzEfajkHn1rmHB4d1Wtq85Tp2tgG5HFvF4sGCTFMpelx7x6rl+WtIUhX
NoCtQGPMDXoXgmX5kMmAMWt8uZRiMlp3yqVlDC8Q+O4rzmdtY7lvuP2ibTXo7ZD8Nf7DmNwaNboF
r/vcCh56FhiBRqlKeceotT3FteUmLDQbs3LZQYph3LWwjdLOm15k2kG4sPb+g0wRwBoprYHRdzsV
oNta4d8kXZ05XYzUZmYslPm6GSVlAZped+LBNPWuAmawksfu/UsGXNV1SBwI7Vpzl4VJFPWyZZW8
BIZ3cr7HGx1OFGTR9gpnXRnJqUvPEHVT5ZCeq1BQcQ/SFBfjdOF7FjhqynHlwDVcLewsKhiAyClr
LRd2xGyQzE/KjBb3x/o0xpuo8YW1iNklNCK2jEilHsJIlF+zyidr/lwgt/L33bA23AWZe84fS6wu
5LLBnVN2J6z7FW2N2dnghhaHjXznzjOhAfv8epRA+W94dj/pT4i/Cw50p9U0ROyCHxccmPyRmMNS
reKzjb7d4QY5QtRtWkx9yPPWFii8SWDNoROyul/uUIuSVQnMRuBOOnZPsDyzzZim7h6Jl4axMqKf
6BN8IPMKrwN7bK2qOs0n/4woWMDhUUIFkcOWc7BGfF6QAcBHON/HR7vm4M1FfinEdFoD+3vlJdig
FaprIozsdhGe1sFU5Z0Cq6hbjrR67REF1EZJPM1bD5VRM3HShbrpNfoPhZxYK5KPN9F7EnHw+DYG
3OzKXehw1f16WdSGfmalnGvJEPKoOCT5Y6LTM9W4h7XDbSwk0QWkRJkEhDu/EL0uP6ZrsHskh4zU
cJbiT/cnIS2WbuNhbvrhO8wEVcAPXfapHK11RFRyX1twRYcMni37KGya59Yopq7BXTiENxF450k5
Fp6ElslJmplMmRPXA9K0iwZ48aJFo8I3NP+dMoFTaFvBLpDlUx3NKZ3LyUrGmjHu0HMCwSlFdSNc
o7tPPKSby4UxIwO4pC5nvIeDp7VzqmhoqoUj8x2OmQIkxha489hR1TgWhXwrtVL9KxonTslaYzAq
r3OvO89UI/PC/wMqcdmdqJqaFsHa3CEVMuQ89qekUPR4vCzAXPlislP3OwOYzhGUYWGu+xm5JusT
2ziicfR17BYEEL1Hdm+Lskfk/UM0tCv88ib1ci0lyTEfkdh4fOYjHH3nHJTKFhoqlAxTklvVGuZK
HspLhP0H/rb7BUd+8oGUPy5M0u8JmTTMxhvpVIhQmrH4tgGkKBNUV1Eu/TW7rBIxZXQ3Gz5rIbkU
CnfTzrtLag0M3oNOv/osm90xWiAKVKMfmQM0Dj9cLBM8yF2WTVVEqqiIYWXihnEBRJ16vDMsoJhU
8x2q/YnOQtdbGoNHHq+RdDcjV/C4iY7dgjIPA6XlONqwRSRxK7GVaH9cQFPCcYsN5W3GiItycgOA
b9Mu6Zy+IfyROP5Yh+ls06s1cr+KovJK/uQILk/CcbEeY8H8WQx0yWrkX1InV53oXcUo/HuOn0UQ
pqjN3ALyYKDY2E8RgDkhmYghkGKVREvQfDF0kvB6eLh6pgBQ5rjb0tabUgIzutXtHT1i0PS7oIp/
pjokAerSLc1WRTZw98CP/wYa+uMrFdejOMqLaN2Bwg22GOmeJrv4k3a5aim5E4XK3y4eR3bCnYlj
3EkP28QVgCbT3Piqry+pK3wlU2n4ySNvc5hI8qkCA9B22f2rb/b2cA2wKDKCv4po9EtQpQGISND7
M5NCPht82Zf+t6m3vpMhhnvOxzlU757m4zY4eaWDFXPPxGrOVYD58MSyyO7wUUMVakLPcKBxns8o
JMXLZTqaJRsNrOafrdo9WbShAzLzVulCRAkCXzM3lcqD6XSsFWtcLPuisPyL9R8SvVyXh1n5VUMe
sPq8uCRXgiWSwXvGabOIY57IlLiZtNxmunK7F+RKzVh8Wb76yPVUkp/QNzW3D33fPwWX8NTm+uQu
QH+5XkgFZHOP51kCyc/GDQRi3cTPSwyowClHAvNsiJ7o+AkjrXpito8HMXuTL+ese9ya3+0Vh9kO
ZgbbQtgmxcLlj73DkkBEyuTJQq3mlBEYyMbK7nw45CFaJfDqv8JnRLCi0GVHNfePMWqvWI1OSxCo
/DdhYdoHSrc+bu8joTyBYe9sMvF7HhWyReaoboB6wbZVzR7/oQKd2oJzPtNPVUc9Yj7T18DnXX2j
VrsC5XHvEfO70PrHr0CfwIoUXUrN8bINSkdELwAGyWiyiw8DWYcKpSXQAS/JV0qlbYflcxHUsEZP
9B8sbGP5mIn1GGcrmgB2OCZJwkMXLDpwmcSbWOt5aDMVF7HJvyVZNXFyWV8U9CrEwF2LPe+LJuDx
h00VB9YqcCmYHi/Gm2guvoAJeNFh76VVIGwn3olFYajBfeKwr6D78YI6fpO+A5IOlOiEESUxZcxU
AvyJfdqEfLdURfCW2Q/q+1AYDPQYEEBS83zPIJemC+/zm93L9BQFxFT7mQZgzueAhkvFiBfxY6DA
H+HA166wLQBMzFLwf6wO1O5YZyFoIu03AyhUCmIrY/xBAfTpjD4ATs1hZD8v+uFccubWhUrkiBIg
nArn3Dpw9nCRRAvwURMkRq8l8T6hkcBhWordq7Hv9WVBPBuNBTc48ramT4RcE3ooqi3EHEYBEJ4m
mIB3taI2tQM992wYiuebdTHd9Th//MJuNeAxw4XjbLy9io+ReopDKlcaedRmClG2woMY2OPzvr5S
fkpDieelmjd4E4NkKTEECMkA7ZIvRonwgH4RFvDGJKIMHDSFQUbiZgBWO/UuWV1DZNAj+bKOTAQs
15LWFKkHfNkNLA+9S0IXrG2/sIr4VxT2pRjSpxbHNwo4zGfYwGMR7DJ1fSGKrsWkbWoOpt9xmCYt
DJsD3mJ8+3q0BxlfzDQcqtyM+XxP/i3dkUxZytfG9M6iug81vHZO8YrWsX4mXAtL/0V4uw7NwH8K
LKu1mfJZTMppebHcmQKRmhdV/sU/edYwh5vwofy9842v4Z0qsHtVgG8I7kTGVxLwUINmYVU7RvwW
MRLEUQIKW6itw4eW4Aau+CRC5fxS8zCrdnpyh51mYrQAY1NwyR1SDStJYzv1C0j2DgGeAydiS3fT
GMjUDM/kl9PHqADgeVZtqlADJlwcaUvtq6pyV8UMUjeFcnIDgxoee8l1+v7PaJoDWnTxYbCxgGgw
H4G/0OonEAW6EeJyxUSwUj4XVvGu7uE+RJtjYa5+VtWx0eA1Z21Psn8d6kDq8LQs/f+KZSuM2C9f
I1yByK3Xogr6/1koHwCjETZSuHcQEqZGcNVNEp/w+iNyaabiItzDUZc5IW3kBbfjIPKnohxzKDqe
oycbl7stEdc/+ABqn4+kMRdeAiQHGCJDWsgPfY1GG0zg8IUgqrqNclwLX6njnsxVrms5OjTZf/04
NPe8TCdWqXPIJDe3WIHwIIArqB7fUPndRoO+eNNqSvpN1tZdyGnV/nY/mktjQF/PFeS1yK8yfqlE
rccEOTqe0w9RqPk3eWPiysPm30YA4UcqbO7Ah4WS6hkugwQxZYqxc/qUNROaxVrE01ubYm8ptMQO
fVjCTLEQzVXH+n9kr2VNry7wcxJmh7LyGeXHR5I8BbzGrVYFBvmDkqQo6Bk0ALDKeXrh73C1qOyD
f/YCbU4g6Z5s3DVcJU7DD4Uf2Zh0YG5cHsxPnEGRa1gxWrB6PK+RRLbLV/yhgCRQU/lyxcEdLx6r
zJbvGczYph15m9qKBVYAKWTz4XVo7jYuPd3GfuEMylnZ+BywgIRRShIarloQduiL8z6psuffLYKS
06swBtiA/D9gdyWP/soySipB1pd0s2L4z9vJoxUVcUR4schJODzFVFLWxGVY9yZ837WfYbUtdFnC
bYvVHtHtfz5SwVyiNpaW68NXYCXKwV+zdfkA2c8Ea4TVB4RIxtvTw2sV777ZnQX3WKgz2G/Iy7yb
nX0HZqFd3BxWdEbTEf3wBH5oeYNgdPEZUvkrAz/32GO60AaBI8stDSJUh5sCvIGEmA2QN3mdPGvG
WwyEMmDuuzGTHvwqJOSMvP8mUf6rSeXXFCy/6+XpJ3FPv1EZWI8kEN/8xv1Ihyjqd7vJ6yxdyUXv
ofWNZD4jq8KFCV249i+VHkS4H7kjxu0/yrSPB19PxkE/iq8e4B1p49oBBJohvlGHrVADezziGxtQ
cVamVMQTfNulAFCrYnpMqYtznJVcU9opLZ/zCVaP0hiXE+dNyXmvEAB4PokwBgnvxswBaknkKleY
q80RCwTDXCd9M1SjQ/vQjL7z2TH7ELco+gUTP3LdHN5y5qG8PMwsm/4HtJzCblrqYYdMqnf7nMIy
zg7v4iCR+M3XGmon1IFtdItdEVdy7R08epPkU2eaBCWwhv6Rx7ri1/KqvPN/EuD2QBap8PAYG7Fb
/41dyBDmcIFbpCdTBvhfULJ/zBn79DjU7eWE5AjSXVAMZJmti03hOH96HddVLXWBJHGC/VpZFEAr
QfRunQgODyax7sSEcSRao3/9AX4y2mHdw4s20dbdnV9rMk26TDUqOT9jGnuL5rz82W4xc92Af9bP
zy0aRa+lu84E9fibwq81jJZTUPccpqFL1ME6Kkw4VzoTeMjaMYVCm8d5EQdOLsXO0zQBh9cvJnKT
Oz9Gv0cq1Tbn9ErGyFq7Uve/9hWaJ5v7J5/O9t5VU76dvIPbAl+H1p1Chn8JIdp33xTx0Umf7GGe
SwROqSjo2EreOuwRY8MAjnQpK4OQw/qijexsE2L1aAQwfZtM5b2MDKl2JxIDlcxBdfV6YhxYHez2
c9rwmXNz19VPc/ArCE1uN+2SILef6zLSLWcZgJFw5HB4iCZwxeFqnd/UIdaRiLxmYmx8hXIC9UsX
3BE0PVZ7OGUuNG05SloEgER1ICcZmB3Ja3ICOgdO2RvYdAZhG1pyKFKvVYrc0kDXzUDSH7PxKTZO
eTwSATpSf8yWdrtyOaFAKR/nVpTK2FAH6sKn4xA08EGIYiO4DcrBi88VpUYFw+sOA9erXjsWdNN2
ss8PPL+gPsSZiwgyjqKSy8Fw174/vXnEN52SuqUeBoGP/hy9cHqoRUjJLDkWW92DV3vUhjbMy0ze
hXRi0+066sdZn6fnIidHtnxYPIxt559whzOvnFVMSSyHu3yIYKUSi73j/hyaDtApp+qeR097fRma
RtDWpao1K4CArC3HMkL2eQPNf4V4KFDFzFgcDOzYaxpAWi7MfclP9fMN950lLic8L1MUDgDDXEhg
nDx2mTqHdQxnqlvWv+7LabYOvsTweqyLwxgybGpf4O21bosFc7ZJhBmB7G24paH12EwtkGfd+alS
zCuqNyZKwijN0OKSWKFVUtk7Whf5eOm4rMcXOPgQUslpj2kVuspwavsCzsDxjnibOh+9QR+ucrda
VzxBEpxfvPzC0YZD5z1G7EhpfGg0saJGrEqvXm2JOYpyyzosAPOg5UF9pjQ61BlRV5IYzhT8CJbw
c+3yWQ2jc2Dr9pMOS3xO5dWRvbQlZmv3jeAhCC+gdfY6ZZ8qkAvmOXixxibEkvj7ajFHKOpSp8DA
KfpgoyabMIzv/10omxyOj5MoGXwKsazsomIUG8nCuvGCJDwryoE7QkLw223y7WSTXXFQFqedjqeQ
ZUgIYS+0seRSUFGJKndxzGfzTYFQ9xSeoBoLpZeyGGCiN0qOjk5wOc+1r+Be05T5EQR0lUVN3EEQ
m4SIcghuQ+8JvAIjtix2VmGYwG+TMIglpEnaLSMCNjiWAsiqoj5+D2UOJqYVqZaU1uPKNRCJXiCx
EoUu5dE8as9nwmMrTdmuLiNPeLNt19hyeWgbsQ6r4U8ZMSQUOQfVrpxwzmWUpdwi7GIvg+/8a4fR
9VDHC9xf1OjqiyE2MUI4yh3CIJdQZdfCoH727O7sLF3TCKPvRqasY3tglEDmZ8lzYvn9E1s8cJ1S
1wcWjttuilRWrWj3Yf54dnl7wJAKZNHbyJMbYLC8Ge8A3Pb54uXdY1ofsb9dsmX8vPth+tcuTSyx
ypV37fLJkD7o6Bt5xvA556PnqYXy333qpkJlUih6RW5tGcscaOlCkW6RH+wh9bbJKl0dvmYlhI/D
xnZPKdenhcq9ijT8Fb6SPVgMLj0hAGQ3DFVtip/Oy10FD103/jPDENcn8FtXzRPUdwCYX4ULDYCB
F2aYjJSoyWR92PUVjhdU294onFhxglpL+53/1y1FUfJFeb8EuF/UVtybO3SN8LU9swuUMI94ENHE
9aR+qRwOQPXd+VcL7gdqpsw+ulM3IBbRnp2+DEw2ecqSVwu0zq2S71+NH9/qH86FhxA+9bOLwIJB
szHWL5auL3G2l0NTTZ3KeLK5OSKzvncoX2N0YcXogSsTTefWdu/LPxg6Hs2FBP/Tv2B3qCWgwMuW
4KSmFnV5rZ65LgPIFodu0WZJQIs8/5aSO3X2WTSmnoWFYdLSQ0GGrKRS2ih0I2eU+2sdCvn3v7Dz
GCxeO33efcHDrjLdJT1ZQoOLcFH4lnW9lwDB00TExwZ9/8BimdPF4pu6LRKS6fm5fwboauz7Ibo3
/5YHtaMBXYVGALejR5vvJEQPiEsTPgCAP2WKIsYrFeclqJ/7vwPxms0Xt4oSlAg/Bo1QbWwjDWLi
agFEG1Z8Kw1tuaB0YZkia4gd2xrJfZtZwAqT7sNo8VO95BS57kBrw1MJMpCnOxrnZA3NPQ59s4kK
FymXSMTscHze5+y/69oongrdESCD7kXnXWoFNS5dbCZBPqLIg/scB5XrVp7zR8bZcm9PXahl4uUp
pSv/7D7dDZP2Dz75qmqINWWZifxzkAi4Hsqelkx13sRQ7OBuQna1rtsYpLm4UhW3NHoZWr2LCgys
UrnIp4WpJnilpad2bk/FPQmPLeEak0+LG4/kirQMnvR1NGg749jMt3/SQ+TNc2gbZzJjyU2mUHx4
q26T2Ndg3bMqUyD6Kcx3wato71r92GLHw/dJD5s4cqiAJGL8rrcU6Ue/W/szb6Q9AMZTbZ1OALnt
Uv2g1837IUrzj6EsFrS8GuLpBWYFniBh0Sj7FmMdM+Kd9Y9rlt06r8DK4O5UmHjL12x4yy00OS/Y
eeHH/PXCF8HCY8EFF43Xh/cA858MpUNFdJLO+SnoiVKs7cVFOA3OEUKygFC5e2D0LWu9EI8zE7M+
WTwiy9Tva11jPRxUamv0PIMh/IxdUbYwDaxRzJSeXwdJUWp69IDc87Bvmp8rVq5Yd5rwi5kt7qLO
a7doYpdN5PROuGpojCgkNIs+azHSEDui15Aox10tJPXmcQR+fEHi3HvBdYKo5i6D+GNTyxdT6zpP
VzKPIHRO8CHM3h5CbeDULGG5MlIiGThO/Y/Exd1l1MVJe2ihsrzBIhhza3qUdqdHMR0hwTMWwtL6
i1VnjFu8/P7jWMMUNCAHkxpAU9Hvcp+p5IJULu2PrVxD7V84J8r71PG/bsvfDUdsIwO25GL06wnq
6ULWUNb+y+VQr7A+zD9RIVaIep8kxhB91mmb5FNS1sj3WkrO/9udAhQD+LbTrXSBy6+s5nq6O/2+
GNnz8iVR0WFkq/vDqgJkoRcksXHSSsSrhD0Dju2327Eoc2KC79/UUhY0DxJKmYFOz7Gy/58ZzToT
Szy+JKIoiy7t1JdtcPO39YRccLDFBO5VsXnAntD6FYZ0TqBdMNAEB4YU1asugdZzm1AJ1LI1gcwc
TqfDCU7nsVS0hkA304rGiT8o0JdkjV4PG9pTF/u9rNGx/TBiBPunBBX/aar79LeO5vaPuAQB1tI5
Ot49HYrVQLpjHMlbyM07/++I6DPnjeFYUbZ6NtwtEkQyvfdO3wVId+VzE12fG+VUnfVFpQePovtM
3Qpf/z4o/wnXfpS/nVVyoXEQD+22oiBrK4q1wZDuRr8BP29ij/q4FnkQeMG+X/1C8ni93PcZb3Pf
PE0JPale+8Tb51CC2dRl1nway3JoLbxQey/jwgSllCBKLIIlIJj0D0wybf9bcTdBF8WadqM0zNsW
u8KeiFmtdhPr+cJ75wh/czQPQsOk3LB/+h683NHcTy5+DKwSi1FxeRA162jWEMvhSEZzfWNaG7yu
bGP8lDf1377nkrNw6Tpns52zyRAutknSTLkH0k+vsYOBnfdPj6Oq03cMdKJRhazjEiOED4TFzxNp
lCs1W6ePFMf6a9/dVH9w+bfwP3hc8aYErbIzA/niDqpqlyuYegJ7H3HKdVDTwH8yhMwlVqAoHufg
P13KOp3mmp5zoNAj7RzvMcFEgbt9F1uv4xNJZcdJdVrK6BuqQFcPcTTBRodORP+avPwyq76WwVyW
5BbUYJH5WEpIOuR0gvv6syv3HZN/l2tn/9RHw1yZ+SRq6zRFo5gSoz+KRiPvakSm8JnFH+L9Eojf
m32YYfWcy2ZrlLNgLpGXAgBTMJ0m2mRkR0H2sZWdDvZsn7EqyL3Vy1JU8/fWRgji8YK/xGMkC3mX
UHH2fIlGEebbLGaZi5L5DeT/XNQmCgKxtK0mGmAkhgBXODnQUNDO7JWI01XfcjsUpqk/c77eG3IF
B75S+UDq3iQgsztc2Fnq8Q7c6WqN9MaHVysV77Jx0sYZxW8z2+BSKOJJ2UDAzqVymjEXOJqWJHXL
smPFzEk5TMqXA4P6IdBad+RUzbCq5wkAHBmRGSuzZKR1pFJvaKEXPcPJRsNUT+b6vvO59pK/2kCu
Ph83i1IheQu2D2jOmOn3ljPLoP85nC5Tp9kJ/FTn7mopY5qMJAu78pfZrGE0qaZpXVLwxmY+rPod
MKNWRFZ/0YlxMwGnuAnzMNOIW6yYb2b2DiiXNEwOQqDE6igHNTb3n4V0MMC7jL2cdQb9IZTsyzIb
Y1aLmpI5/RwF5Uz3ftKg7G7gZfPku9V4hOGtvzimTAPaMBZCM1J9PntRPqqcvSYK0KtbXlKlEK8t
4LBZA4EysrHHuQay5E+0v7QbboxKBCV/d5xmgeMBk6eOMW/hvoOqmkMQLBt1iZdrsC7jgvOmd+yi
XKSg34ZwNBT6hsZW9UwRzMKT0B4G2e8g9doeiIvhWhUMlOzNZudwAMxziG49d4mPY5xWLd4VKOSC
fNFO1APCGnVD3JZyT2RbkhkJYIp0fZ8H+l/algtIbIICf78JJKNSnWIsayhSKrZupoJNApvCuY8h
SvjSaPWoUBLE1dAOQGVKJHgbhznlMylanxTitJed/e1Ak+sF9KGBsxNhWC4b6n/cbMI3E3vDbTT1
o1I6UZ4tniz8lIgIwvtFiyeOUVht3R9QXwK6+3Yjw1r2SL6ZlK9Pp0zvYC7Zdejwh6BFO5puxnzu
I9NyVd6ZXLZVBC2LQ/YV6deGJRgqTTEshcp1Av01Cdx7koYPb149mL9b6pO045MNfNnmYdBeyXXZ
i4wZJOkNsKoL+NBT54ZqIv7fTmfZ3geUqWlnsax7eRuuK75Z6Nc7/UPVCugHvh8iDbTqdCX5sBnS
eZGs5V2xdddiuptm+vA50zxCw23tGIgXKzhxRZwZ8HElGYLW+8znxrkElfy1fZtA2PJRWqzxUKnO
IOVJqAT90tIqxyyb3zdvvt/nXjk/dv0zBdZQUUpDYBI7MD2uICZNAlDHgEcFi3VjY1xikm6GVg4D
qec1bH1PubEYsWiJgUWgVnK0YJjgdqElxONpr5tuj3YQATgZcWo8nypTt2DTrXfnh1uehXAiha/n
858TEbiVRFSToPjDra/wyOqfGqa6oM5XuCQe37YIv5yWYnxy6mZ/bbVF1wSoHGSPmv8WAT/ic76z
zZ/nZ3ABW3Qm6UZbeN2uejTmXYg0ikjSm/H6JcdEJojCjWeq2/kJbEbcl49OnhwViBYdJgLiokyC
6dJDAlajcazTLR4BYIiDl45kOj81I6Bmtdu6XFkWh/KXd81mHw2DAax13SvcP9NcamqjgjMAE1Tn
M1v8xxQbyg2ffKAPDFMO8L7I1OOS7dV4SZ3yLGQoMlyLz73e3/cJFR7RS01KWogFiqGcee6lqnx2
1LlrNeL8LONUUxd+Us6zqdsOde1t2GsS+n6OeTsSzigbO2enhpXG2xgwLSVmlEAObji7PdmuE+9L
Oe04ngUV5A/CAR4ded2QQRJeb899nHJJFZkbZY95Y1iqAlzX8wtmYx3aP6J+jWx8NL2P00/PPnAK
LKNblwK+UFV1mfOMyWocdq0MCnCPikJXMxPbEHhQCm7OM/wjoI+ft1ApDd1Ack5l9VUYOQuRS56W
qGQ6uKvINd48LHoaS71hKF7qdbRvlXMsY2bxBeNRvRACByAULmbLUqzdbdT2ajjRI0HyXEHSJNnV
0NC1ns7eWCZK5YPEg6h7JbHJSco585e38Qle/7kUEq3Q1hFDxJ6QV9A95ZAFgD0DFR+MM6zdLdxs
QxitXjLz3t+5COTxKmqXJAxo6ZG50HlONk2UFJujOyM8qZzQBu08PQW+TaX/+PfvibAwfc1VNh9U
AjXsY680rhSID9JxzvM3f3ZexxjtL/ZX+YHtSLZAFg0szRyFjDhOQR4OB9OcQg3msJ4Ylnz/8BL2
HOrhLLeVYJKOmf5zfIxOliPbXwqBtj9m3yXjxM9hnIkamir4KLQkgUFqYQzckGMLoZ/2nVrvNaIg
+gYC/B76X5UrRl6Eqxd9b1ufMUNUKqHh8ORRgtzI4ARD7Z1aNQU2KPKZ7XKhQ9r1Qht22nZ/M1Jn
bPRTUx7UXtm3RaTX9HfmZpfCqERQNUThaJh6GWX+lgITnQqYyTaXpOuEqNHlPJUbe+BRTuoyzcLX
mvm3hVB1t7z/+qw53ECDtULFEwyALHij1yngGCRxDeTAB839Y8n7ZkH/clQA/mqWjAkL/8hGjVR2
o8TzVSo6sIzKO8JsUz6ehmee3s7L+I7jEi+KszLlgJ2w8+FXZF1JIMkRq7OScRh76WHyS+S6amnO
KC93MbmHmjjN5qXEzhF6HFBX0dqIuBOKAnYCj3kfXhUfw4n4LoyNXOoJ9iap+XGJLjYSCz3eL+VF
tnZEPsT1Q6FoLzy4vgFr3JmhVFwd7jEqgAKu9x/N9qiPdPS3fH65CSFiJLR6B9Q2k2lM0M4SAfVX
dXmLPCqLCrDsrp6OXlBsz6hjMONJsks7vlZlGeg/80OXH1WUk3nekJkIK5tmROPrsuNDHxhsPvjp
xcRRfwix4S4EPBFyKwPN4e6Vawsfo37sN6Ncy8B82SSbCkiE3Yxsxp3E3AqXcocaopKMxb11zkQa
hfklJnI/dkW7zfM6dN163yUrJlfqXI968W3PVesaqC1PjoG7ChoZscy+/dD5zbiL8En/8kqbgpAe
T3WhHOe+t5miek2HHP82S2fb23oTXhswnb2/9vymoq9eoQ1FtIARWJdl5xBnsOLMHwi1tn1OfB4t
fJ+meFjZPcx9u5JRjZUC5c/miZB7XEEb0FBUvhgM+buQQREKGxzvAt7U3jxteGYlhIXFHj+Ovwrj
r2gNyK07uCTpdjSsJmZEfu97NHqfmfp7HqSuQVflnYQppF0D8kRqZNMiriWICjjdXHr+DMmtdE1r
bR00xhV7xnayxjcT5q3tIwq55sAe4KCBjoXKW8lAz8ROjKQTl6vRdgs5T93SFWd6zcl+XQjyPYER
gz6egPcy3GFA7ReIgOi/EALD6ef0Q83J7MfsMMnY2ipQtagcNsLAX6EtAGoyiveS38in3l15G4Vm
OpHmkpHskvBrfivqxaurBhcdzuHxmt346lmp7bHXoYE4catlyTiiGvO1cS1FxXrfLYRNkUR/zKIe
kkKIMbS5cZXzfW2Q4Ggx0EztXGDtNSIs+Yja/GaHvGW15+Os45Lql2D1DTeRN9YNsg/tHmvWjseL
cw7fHQvwUSAn0WMXzdS0f+wn/U4Av7CMt9ID5xIzfiivX5SZOc7gO8h6BhsLM8XFTCV14SiQHl2t
W7IFSUO+ogbC0Ght5o1eFWMWU4IB9KSOVaQxCWIaguKjayBm8d/yW+dbkpvqUzRX7OpfqIfMhH1H
sLyd9RBD3LnifKAh2mnmT2eo0m3TE3hIup8QGQocAk+Sy/zVagU+ZmLM7TyKsQOAsv3PZy3Kl9vl
eLqDAigezoOo6jm8Dd4ziwd7lGUwJlqd6DKrv1bADY21irGkWWLSLX6BbT0fjUSSf33Ggd8dxKA4
o4YZkKgvKflcng7Yqai0A7mK1LEmhyIFLac77Zl782zgPEaxDZSUiq5tGAWJtDk6TvTQe24gyYzK
zSe7+KmiqVPG9H1FY4meRE/ojGpon66j3cu0jdtuAx8fO8BcjX7Z6gfNDYVvIR5Jj4bi6alqAW1i
DRsjZm3V86Ia3bCdXto35JDklnOmBvy3K2V5JXSuMJKKVODbS/nu+mtmTHai2hH+fpTdFd0Wgm5b
ugnbVI/tQKIBabkrLVeKvu7VCZvoXhxGt8HS+Co9hu/PU4olmk71F0YUyEkO7y2EVfekfvPtK350
F1O3QMokwOqXds3N7tcNoojBgE2sac7SVs8yFbiq9WTBLbfAHY+2ykjsHm2d2WtvCw9GUBnEVea5
uI41cY6HSYzb32rfefA+ia0Mnf1lN5HVFS/SP/MAJYYrLolNOo1YwAZJZ6eBceJxeTGD1+5c8HtG
eclYNmwChbsxGPlazodo6ly//unlmx6kp+zlbZx1g0Aq2EDQNJ2HYXH5u8l1eScr8P5tJk1yWH8o
nhO17liGBfuvlwEVPt2vy4YyCW72mPJ3yvRhSQ+cq5i4UKsKfMfSPsXm4vFSKqUUt2PG/+sdOiSC
z4LeUUI4iqC0vWCLzcleQ8g34JmB0gdmEVuE2Go117MneBKcJicAJBeDR5Yk+xpyL+It97nrNBIZ
n1wM3dwGWyZQR7fu0Fc/KLsmstT+bb3BLzc4JPolU6Kjkr9rg9wy2w4d4ME4Yx0jGvcKC9RI6lWL
EibF7wbhlqP8/yh0LXko73cXIgrDv0L0KHTALbJwrsWHlatm4sBA64uEbS5u03asRjFxSCW2L78m
kSVBd4ctJv4ADUkjX658fPrlkqmkW0JkazimLwWItgJGSPgqtCIq74Znv19+lMYt7geQ/Fy29QhK
m+W2Q76vX8Hlgll1vvga7MhOLQWK8vegBEuHIrCMs+dyKf5I95pR9xdHsvIwG9MMjswTro9z+6Lb
8mkZvnWy4FoUT9eAYUnl2K6KIsntQCZqC4hyshZW8o1YZknHv3Med3/DNdmUhi1o+BPNZccW1wTu
G9h3KpKSW+SU2KR27lwe6Ca4Sptxlv7pPIm1TF7LZBspwv8oBGISvOOnhmr5mzPDEEcmPkhH+h6n
iloEyBGNCoTXtQQutMuxLYu/rfVX2oitC8i2LU3QYUlMIZuMq3AruqSenwUSYG2JqJRfbLcfKRw/
ZSxJSUiudEdP8QgoHgqgQjT37NiTvkPbXhgtH9juBRbXeVEEqlGf4fZ2U/df5VZ/TUXKQYjBojhr
O3wX7v6z1NR9uLns7Eu/ifY2NBiPiwgW6EeXLBciDsFbokBoSTfTMN1KPAKTFMVfhyYefZJAtVzE
N8IVc+LLYTNz5BOwE2Z3nKmJDc3rzhDJSFypYlg+uQXSoT86mQcd1dY7kHbSRqrldedamXFlZv6C
reDIgnEarx1zbaGl5HEuOUgFbOBYv/5gLrh8Tpx9Maghvw5sSKRWcnCqGhdtlhoc9l9nKgq3Bd7J
Q15eibksLA+viLmJa6spEHiR9n84+IvmonDsK1Gd7l0TSgeByMtPhnTVJ8OQbmW2VZR4Psp5iSBr
xcVKjCp2sJcv0osstZg7tiuNqzCT8sEFEpyqneLnAwgqF9fEPKBgRpwvwoTr8P9kOK8zuve/4HVA
k3Ym7pZkrd3GDYj+cqoRCZgHTFD57b/apgXKudbY2xWwOzW/XDXULL6PQx1tmPzCB95MXxcFCo3j
MLZz7h9qE/YqYVRQM/z9CihkRytma8OF5W0O9/dd9n0H+1JGBmFjwrDouWuZSf6+44EmjzOeSuX8
vNuZwnt54ScaIoVNSdigvNLh+g4NDHBt/R0vtVBCquPzUl9zj+6CEIvUM7JGchYRUbQKug8QRlFK
QKk9Drn9NbcLRjqnXXpV0kf3E5jElRWlkG4htMUPy01xwjjxOtu7kKBSEi4jHWrz8Kx7iedUBmkQ
d2Z/31VrXfqQd7Uv19/LeSN+3D1WKbFYZzyciGDG2D59af1IUg5yQV++fsFpX0FHbGh27fExT2sg
0yTz1Q6eyHA/T36vxncRn4HnOfVcV5Nt6dgVljWOIkvaCdDBn8UrliPhzHJb2vv9+fspcXCostqR
zCaaplzGjuB1ivcuufvRJEj8mb4m9erA2bvF33KxZgWhLS0S3JYb3uAecati8C6t4N5BRY9cnG4s
Y9WPqdaPoqCG6FGlcvTS34yiTBs0zl7Z+Z6JTCRSMWEZM6cnPvXS71QgYfypDDN0F/QGUkTbAcYB
WZ/UJEIWVZecMRd9uJd5gm3hLYCKEiTzWU4F1hXhCDTWROVnnE5K5t3qyiAMu5KeQ636AV9QDAoT
WQlSJ79JuMWK+oAJRAyC0GdABypG+GNBanRiPCjJQ0c9pVF3XEFzZQAo3MLeHZa1jYIch73N7VGO
vJmKepGVMArk4sAiH3gv8V3/3wkAL3lrjKzAOudiIDXOVvzAOf2DQ8NbFSmmMv17lOEAOccqGPsL
YvVrL8iNOh52iSE/fyIrcBJn3NdHXl85ovqbc9oVOxY1P9eVeWG2tsPDGhe61EaAJ2iC7mZlLWBF
wGe5MjXZgrWaAtW61bYqJHr111dliFE4PFSJKqz3/sbpVIRKSzUUH9VlXvPxeNguMKHfc/enehml
ffNzrivaI6ZeMLpCSLVLe8xncMytMnrJ+5Z4+o5sxWNHaWYfVgPY2if5XhYMDUcOPSStXUxOrnJ+
2Sfkg6pWIGq2dFpvxuot1D6PKd/0RyPDPRyKunCrhoexhPpgF+Wb1jJXdJYr/+h3jz1jPqp9lJ69
Eah0u4bvOmy5iogL1CL/CjEDhw7OOlkBlOv5jIwGO+gMtuqGiM3/tlULm2/MDNHYuGLNpZ1jaRMS
8Kq+SBxycZwE9qBKC3EZZZuNT2TVM6tjdg/Me7U4kh2SNVVoWqaBxQ+ph3e6EHydMmDnbnlKYAh1
5kvn7Bh7vBmUsOtDHlmjKGm70buzO8o/JCcVRGc084Z0F1uu1dwkjaNW4bQVj7AqP/dfLD1pe3ew
igkjKIKmCOVm3qFWzjX9T+ziR9QgbGCaOp+kktYFU1YUAGqbb7drMLZ7Ckk2IrB9uLKexnB533QV
B6BTLjI3oib+YEA1IDo1NhukZ1rIUyn5VSdnig7+lvU7o3Q0ChTaRDv7Ovx5oulqEnkOoylhs6v4
LzXgR4PXmX15Unmxv775mPnH1eAdx+ZGt+v6SFV/yBY8pz2wYHh+DIEBPQ95Mrko1WodJcmqLL+k
zoVoNe68+BtXn0mcXIKOLZttFrw024WLNXwZXau/RsD+aBfY/vywSQkir4nM6sSP+LfUDkQxE5iQ
lvOYzmQRgD21VykkH100qEPWNrm7iPVItXvixYYGJ7uBVwTB4TvqPSEXcFgSxplA78CcCOobPK77
1QuTKRWfQRfGI3UiV5jwPS28np+mau9BaPrKViCB1/TLPwGhs/evV7zE7x8IgwecwBpqLSNDiZfV
438Xkv0SpM3dCxav+mlsCTXMZI7NrWWXZ8JEx3zkhFg8zdxzIOOhQzr6+TiwVHpN+4fSTGzAd5DS
c+vQUSal6YJM6sISe7Wuw+uAGYkG75CXiONdep66of4D/9n+OJhf9aAp4HYsWJjIpQhTvBIqXxDG
jpTG0ULB8dR2MuEbzAjLuGDC3E8+KwiixmXeJTn+dMYF7i5rWYK7BmimJAppNmUjPFNHNUd5H4Gm
tr5GfSF1l3FdVqzNzXr+ruyDzowm7x+DClzioP/fF8CyLRGbelSSUCI5EZOyipky4pahvgYYrQow
KXn0PQVSPdDFtnHAT/M4R7PVDjltbpnoYY/vXkVvMTs6BDALx/B+HqeMhVNTfqFjHhyUoOR1Q0zO
q0b37BFj6DY4GdU2Fa4hbRxTbfKPa5owd7lAzMDdS8KVS/mnP3y0wZYcjjxoVv//pIjeMsEPQlta
Jdf2GMlBfFrbHl6K+4qt6k8b4nrRPogx38AbpuuQmgXQmAHfkQq8drccQ9dorLnjzzr63esWTGtl
O9IzSR2VF8aZ++hnja4XeUycuLL0Pk6fQIQqeVLhvvBSVbHmDZlgxJiPmkHGuJtil13JZq9quLNh
BrOA7C/IvXlRvmgSwAKnQhK35/DQ+Xxxi0K0TFjKh+ht3gJFSvqIYghzmqFDMICSBKxGWDoODKFv
ziAiFVIq+9ho3qZUIl3xdYEBzTX68DjJ7lA3PKZKa2ZAOIA7nHPtT1Af9lIMO3GkMgaW9mE70Ngj
P2095VfRbO7TTNzCBr4oH0Ns5dEFwtcZ9j9qOHpH/EXXGmwF/PKS0NtZU2qSqivYb646f8ZDiv7h
IdeMYNin5OYoRBXcA+pnHI2c2bX9lWUm0fOYx6uPTgKWmZ61llT7zqwl/iilYeHCj2So+VqeS8dW
J5blYeZBB4NRb2hZN+zh+dD69YRRqIWr5Hk/ExxVWKI+RcaywvlCWfa74MHFUTLEOSwgzE2orGnk
qwDh9kj1mxvOWAFMW8CHXBOFcUb46UBiwuBnkP4gGmdrFiymDwUeHIWAghnk4iGoOugiOwK4bzTB
ZI/0v6z1MqKXFZk55/zZ///TYaBzSWeOhD9WDWBhrMo3GMdzojbTAi3kZ6iKzcDlG3TgncrkGOv/
LiG9hiVddBPyocmI52KCllZ1zyclnINRiFutXk2Lc6jFbuYtfERh51B5obeYA6rA/QZJl2/A/5Xy
MjrlAt4AUOVUeLIKeAgYLemji6y59UmyQbBfaZnN83Lw7Ld6gWsMG0Jn8aX0mgOIaEMb4+VjH8NI
7RrCw2JGL6D+085GsOnUlkJUQW4GSamImPbPC8kNoKs+ozcr9Vkun6ZkRMy58Mgs7UnS4K8p4qQw
AFtiORSt/sMrzMA3VvyNo0PPsw4g3ygTLtll2BcyfHzkkyGz8e+LkJ7OjGKhgG4HDvEo3dq3FdXu
XOGtaDO7abKeO3kkjsaBnIDbszpNom/rKyUVdvu+jNYKW1xzD42HwLymaMit1kXuTognVw371/jX
9SAsFokkvEq++hGrFCkGuBbjDtP7ZF3Z4d09Bwk71jFjWu/TEjcBcx69WNwcswt/jhKR4jcSh972
afxdEPcMcKrCX7kDUuBASGPaSQmLfA6UizrsJtl48FKoOxs9miH9e99L7QZQL/qEuYMrG4qnQD4L
cV7gZe2PJiVJ4k3w6GkHgiZMHcrVXlETle3SB7Y7tuC8EAAsgVbJxNXg9Q2Um2H99KNlpJJXGBTZ
pjhbMPEBZTIf6MlMDbX9zjynXnVFdL/pbn9fDmZh7ESKmq+7ohWKGme2n9TNcn2d3ErwP1dZbAMY
JTWYBn/W9na10XIR3N/Kgv3/WXRNCCWGi0hoO55b1jqK2ZO6ye97KTSqIk0gz6t9hLPsaLfdteTk
Emkk/9Zjlgi+azUo33Sdd1ICyTm0XRxfPyRiqck1/DWHEUrT3ZRM9uO2ZaPDxlF/LcHotbD3oCFT
RiyClMPelwnQtEmU4hsdufbLezwvKkeRBlZjq/mRwGhz4RrnPziW/QUH+PvlPNSfKsukuiWQUUam
09i+rwriyV6PLtg6jykJQp5DHAWNAuLPhuO+//+8ShRdqtfg14Gk9T5M90ID4C4QuJ2QLdQWKsHW
ytGcdvyduIzjxWM1lr+mA7Am6Vr2DdXWeV69cqHkCIjRdum76cxFZXxGRvMdKWiZi3SU3H/ewTLB
0uvoPFR381T48N6sEEz2M39DJkhYUJNidf2oJodUJPlQq+DvgAleMS+rc42TqV9oxqXT0L6BGXUK
uHUHzgFiFF58w/D1FI+dD0ehczbh3efW6DcKS3Fr9/NxKANF/83a0RqM70GWhVoOLcOjgOiMqU3l
9cHCD70yYclZ6LPjzKYyUi0Dvwpd9l9fR4b7Y93PigjGuasxgbf3emB0bICj9wD+KeiySuZS283B
3T5ZtLjuQrdWtwraEn+q1eqeNUHufLRGBinQUbK7V3+BrFImyGHQ5czQjVikTw5wxHCRVr2TIqYQ
cjJVypz1rGJYgiGAWiyPVX4IDK4AzMas2J5ZYg45S8l5eXuyh5R3eCUTgJmei+HfWA+KRyR1wr1u
vlSEkX3Dsw+fesfN32kY5SEq6j2Q0UNDFAooFOOkUjtkDvyvUtFo2YyCQdpo1vm+JWsRvUu4yaOv
pleG3cG903TZDQqwWOOa5Qknvu9kmGkqgMnQA1r0+TTwz2Oci7779ACxTmlZgG1S6Yl/34u1k5uJ
Tx2GLIHS40JGSNr/mjz5GKPrJCL1zgVSdKKdLc7KrIl5QIReacJ3h8z44bUa+XEVD+wJM/kGOPQO
W9CgO0gYhFrbwkhOnmDN7bV/MD4t1QxEKu9jDXf1QRx4PxCmMTKgW0MWUE38xqTaJ5Rzqx4gmQEL
g2JDwUaO824HPR7LEeCpnVBa8q0c7DLd/BKClKlCtdlDzX7ngMBgO63NM9GlwoaIQOtnpPv5WDaH
8xVMZS4GxOMRChUZxhJlkp2rchEjA5W/ZXQLJH6wThZd6VuQvJSdn6K76o5/8RriT5GdLubM3Svi
pb6C6bkfmgss4mUeZlHe5ggMqMhT4N78m2jphBqEGAMw2PRdCi5ECo7Vp2N0/wvEqW6hfIttAG85
XcncLOv8a+Nt11YXb730SpypFn+2FiXCXCa6CTe5OfB96ZcBXHyFPxY5+njMu01ucWrQxN476GEG
z6DO+NCkdZVrpIQwb+FQnR6h041DElKMXb0Fts8hWMNG2x3IayHYaAflcBR/DWXPnxEOO5VKFA7F
LHinJ1zgMjjhnxlDf9yVh7fk1HZ75iMim1xBVUhX/2gry1WJHL5RsCqCjKHtNK4l9bplBgUkpFGl
BgfCjgDrOnMu+pnY4C/paddVUgOes+P+kekI2wgn63XD8L2COzbystaVNzPenPagGvxzjXlz3mBT
1qxGCJm+k40BukCZVILT5V+ohFRNfiHYuxxn5ZHkhQCNJpF50dNiTqkaUrUPt9/4oYqSa6MirqqO
gIGzxdDXliLXXHT2NJB1UsikwZGkF+fdFWBb6u7A95LOQNYdadmVXVTlrcmFEuunuK/KsvmHvtM8
R5cPuVb45uU2x/s2rMoe7qod35aOTKXDrtyV1zuOOrLLFOrJG05ckIKN2v/Wjx3d7qhRhRiPOBEo
PYslYklBUvLbJgJGTUknK15bUypdkx9sNEevK85a5l/CeAYdnYjnUXwxqcKbHrAPps2y6+O4YaH8
5qw0W1M7oU+DGg5zcgViosg2bRbag1LVq2AINZbJoUDanOYPQcE9+SpZjHhTvvKY7zUdTPz6n++S
0Y5SeltzfzEkXTxgyJ8l6PMcIvjPgE6WDliHeGm/3VUCjewv1jeDQefZtZwdgPmpJxJWah6Zt5OG
bQWywRoFJNMg6aXBHvFXHkF8G4YpNKPXpsHM/zuggCSvUzGrHTBrqV2DJTTpPPOjBhNnNSpxrgDl
S3ojewQ3ete9kG6R7EHvImqMo6ygKkIKMGEtwPse1xijG+WiVr3Z+k4r0DEJVM588+lxxnCeeQot
X8hopbND2F1fRUSTrZUT6MX9CR5NOppSTayCOSCOAodPlPGRBSgeC4rMRpQO5rOPZPlYZGW//HmE
eTHyyFFCRUj/C/t89z8jarAIUPEfaMlsDFFDpCFy5eRuUYifPqz6vf5VNgH6oOkoCM96g12sZWeW
dNzymwQ+YEYDiCVQTGnZoXuCX4TuCGg29b0EjRYEiNNSzAlEbCqBk5747SvYfZ63T/7JqO8vKB/X
H0K3M2QfkCF0o8sL1N86Zr83AeijnGmfeSAYOjJj8qkUNmRW+I/SG5dLToBqI3eDElpp7jTgb3cz
lE395leUbAq1dkftzrck51TizVksFdqEy74kPCvRLRyrFp4k8XLkEgLGW1syz8d2u3mxp/BNcAsO
g7w5Z+aQw4YzCfu2YVXA+geUxyDfVo2y6l0/sytROmdwBdcdIhQ7FMh6t4VaxlnfovTrw4hzEfV9
OZFdVhTutsFSnD5DgsxXU5wfAP2xWhVcPQhNB3tFYlmBkuWJtsge/wuMsnsCUaGfyA55tVfUb5LE
d60QuKPxOmMT2+v1hYh26o2yE2aXKsfzcTt9orA3KxvK1wNFdUzEWsKSDeGLnWDW6tyFCX0GdjWO
YsffF2quu7QP0+uZx/5Vw+HGxCAj7JJXd7fDaSF7Ae9GNpgAmpuP44ZU8Kmi6SuOldOpRsJtiPeV
idp2UVAoN9uWMvUgt6QyKNdaa/YEbZEiu0OrQMWjWeOqHqJxXeUUBPO3+Pxgj0/Wx2YlM65UXMAV
599UKvPJidJYUXUySSpfbBRIkWn/A8EqVI3euo2i2jp3bdWebIg5J7bv/vTxNgK4Aeo8kua/LQEJ
Mfbw+KpC0kVimoq5dIAUawQX4ZywUSXoaaYzpJqoaY3j9Xy8MivDYQ8945mX7XnM3wcR2k6kAO4h
hkI9lwMQDA6E42+7XsmEE5+lzqa6pbGTqbAAKMruMqywR0M+EE4bJV3kXA0oOMPYTGRN4nTM+B2E
DSCkgUfMpqkvOAX443D6eoiWLBkLcrFx/706qbjZFMwsyfL++FA+gTZux2QbZdvDiJrszZ9zN4St
Wsx1VPY6VN2raZtqZIYHr03jNMa00B/gerM1uHVuAiKwxyV6AxwCU2c/fiSlGuycDXl9r+r8oJig
xqEA6fKIQYuqHaCWFkLi82bnm3n9HKTlXjEXIhYtyvtIIVJGw1IXbf6bojtW4oIg3kCuMusL0w0T
kg3IftWMtxUaWgwLTjKimlbAue2B+j9DVsbL3NmgtK7V76sAS4+s1SwK+IXuaIIsuyYBDmcIIpQQ
0328cz9ZBsMof73bzCSaNeLtgoV9+NY/fTG17kPOZrrb18Jj4xAAETTWMuleJT9gw6T9nUpsmTGl
RJxbcnXHaMNwOL7u+bCoiUfVYI+3LuIp56X1ulA/WCULqNPCPQLZiB9+4wuwa95XDEq6wEIXTCPa
2p5cFvMLEHUT9WVbEd+sW+Rqrlwar1H2BnQlA9MYpPRPFwuWcnQEb6yagR8Ls19/pKPDYVGXbJ/9
XOsvTNubpwee1qcRNAUwB2FHYkPswQ5n9SUXqTCjZhLOlhe3rthCAKEM38mL5nZ0WrJmFUZd3L+p
5vgDHef8mzAh6Yr9ofVTYamfVjc4z8N3LQ48+h/5tUZm8llUouz08tpDAjP5noEwFu4c+Ph73zqa
8PQbD4eaP9iSUDozDcaQgiWVYOmzk1hKPSLGXWS3osq09x3U1yls0ncPshiF/kaOZyxlFSI09qvz
9uYc/eZBawCLlOEjxfqFTq4sqOPjEN9cw0BnHAweNhDq0Ltp/C5oT6hUE7apQv6I5hFuXcoax9Fm
BhpLKYtRt0QmftZyCwD5bHn0FYRLIJZD60SuOC1/iNFGO92ZZ5onKMAYrurRs9H6hI/dK+P2P65P
H0KONwk+vjlJVKxs5hqMKz4BsKT2qGF/a8TpvrNDVK9TWMwy2xGWY7AwVN0nbHJZsBbgyrY9vCTt
dOkL+lhMDxfY4QzeZYrLewqJbaTyLtjMEVJo4Max6uWo8w9C5/WQiyvK8fgG3971g7wqHUOHD7Lr
Gen02KGPd7MCBQIl3AFBdOVtlwMGvIISnMGbxE7ngwatwTY/9FxojGfGDHIkWTIUewoDcGfThuEA
hKP9+83iZg7I37if3jIata0JaaEsPTHOiMt8oseIrr4Lvx98hcUG8A6REcpLq6e9gsbyvic1bvFQ
R3SFkxgbFTVqbJ85l+vybIDqDA7zHUGa3yWpe0a2I1gjNhoCwSVaMRcHQPLYFiCEONexAbCQFw0D
LBPcLzTq7FAgTwD3mKa2uGr9fwJxWLKut7C7WIFbcAMZqm5DaI+rqTyNN8q0iHS9JCBuxnvocyeV
83uPDEZCdsAfLQ8poO2Lz2lpbzp5azNLhsBiFGxDQjvqAK7qnYSh/Am6qccJbbpDxVkMUQRreGmE
YKDAwW6gGKJswXPAgjhiX+IDQsWEJjDu+TLuVPxq0PJMYhIIrFIbN7oeI3enMkOolglwlQo2JO6u
MMMQJYzW9YXxJV+XLASYC3BZ2hUe5HceBlrqH/TvqYnNMPQHt1k5YLwhWGPGg1LOPBqsxKwqqjEP
j6I1TET9TyncbLpMWg7XkIFzCWwVXfsjKrf9CAn23xpS4F2NRDmF+x+cUFQfhwrfnjxhVq4qGRCd
qsPefuAoFOBGsnPbr8tsr3h4RLE3oAI+UHXxVPsgTWvyE+z2UwN8jDWL3qRl8fz3NEHc0cD8LjLy
Yzpn1GyjbUxHDPxbDl7eXkQIYtiDkjN9VQP5KB7N5gvXZRQMhHcp9C7LF8piwwbMr7BckIJsdD7L
c3M9kif6gOpmFZyOCnATvjrnthYBT3s+uc5eQtvxN0NCno0veuYf4U7CW7PejeeExbC9ZzMHH4vY
ZqTDkPQ5byHEGB1nv2W7QChRzDRE4bFA2IUM0uHgDlV2oHVjMNkr12vc8VgIdA2YgEwUBakbNysY
pIAR0FW3872JqrARkKEdSgpnK/FCI6utmG9zrpS1i87ufsmBfrSY/iepJzoyC/JXpeYhQlUFqe0s
zQNfVHNWlmy+p4qDDYIYpkXJV1OPZX75uTGkNdyvZEK02wh8tE5yg2lZLp6HbMTbzRmiCWA+M7Ok
78wqBmND3urcB1dBAFMTyNvzLIwBFItHnHAzriyqTwglabb+6rLFp/8slLblTfo/fZpFz9UdkiZj
bb/kWVnQ5xZ+9eUUykwFq3ydmbYnlnVVNyCozWsxU9UgzUbCOw3fpKjHczFgnWA0Jl7T39MfZOJO
zEnSoZUBK4arPFGeI5gsRzsSp77N5t8z4s/Go5L/tWM/RDp/I4YCS8gYobauCPnAg9Nm3bOBVCyH
lwbv5Dilo4V5k8wFuNXr9TTvjleJ7esF85a/PK31BE0ls+MSmIWdTpvt1kuaQ1MyxUSCeh1yfRn5
586UU0GyzqPWIFJ8Vvgs84HPhUwZs6zqhYSeghUblLB0nBiOmvbYNwIUcjGPqf0kdSZs3ovgw8N/
+6yWzCILj7mau9w1Tv5CoDBXeeVVLiYm49JRQDb09hVQRy9vAMrskRoPvniF6kplXSoCSNK8+U77
gzeLDJt57MqIOXo+6rca8OsM6IpHI+nXEo/SRG8+jkMSQMq6ez5W3LFl04oo6p64WbRPa0DxOMSe
4XvrqffWhbgvIpbA7quzVU/6Gya9JXY2uIyx0hkDNpmy3koX4T/Wogiz3elcpiPhxeA8Gmx/7hVf
wfwwGF6qNMtpbFAmumBdojIe4ZehS6vspwmQfhmUNXZVszJ+7S/VSMNwnBBxsjeqo5b+6gRPMJbC
x8G/kC2RlSjuDk+Jznpgp72jX2ZqXprgBL+WB/3b01RYd95P/V3AgWbvVHDUKsSneHbIxuehYOtG
bEBggKj0ywEhyfXzcW8JuaWTRMHw1pPsnPNBoA0uBJdZPU5f+r70kp/MIIT8Jyu2w+Tan0amQ7l4
f6luhY+uQeBp2z/jZinry9Km7zGNzqsswdiPuDrOoSMej5sDBS+cnvvyRmECtJCAYz1qSvyEVE/9
V358tWn4Xv0KkffWabDP9mAtzKscwdY59/mqbJiZZeUbWe59CWRXkGe9kyuKqg8zXG1jVj1hb/uR
wXXf8tWXuonbjKKgsSgLM1wpeA1s6XnRkmGXyLPYAvBRDUnQxwoPEQ5ZOuS1XKcytWDHS2gvZLkF
1Bq87YO3pjVJyZtUNLHHLGY87hsoDLUvZ/BdR1/lAR8HL3oY/Pft8zHAfWT5NCBJqyXStdukjksm
PVkWZo/Ux8acbkCNJMnEHgITzeayE3IuurxfgD2oxfChkNitZ9MgSScCQG59dTjCk/9B9r6G0Wtl
A2evc04ZCqOWFfBz6Xq04vy1v4e5KMHWvPUs5tbC1j+ugXcfx14d0YkeQExjOsxiPmUlN14XPjwI
pMyRb68SYRIGPLWNJRYne15N+3is5soVDsDXoBvsUKo4EPVQeUytW3oirMv1+kiT98kWKAbSoZmX
2p1+MwgO3t52Qd1ROFiNNAGl/e09FNR40RZRncVH0LQ/HhE5vo3oBeH+SETYj9YuhiMBGpRgAFxZ
d0EgGcY3eXFDmreFWtYZmeHfnOggt9ZMdwddslqbuKnH8+GMY64BPLZez0rxsZRFBVYcI11LGJsW
xK6Tif4oJugzffyVQrun3Ac3qWSocpIChVYovL0LgR9AuzywTH0/414ovEd5K7tPK2evdW9nvRJg
KY7cHm8T8WSqgcsCEVZirbVSqH8zaNQWuw1WId1TDi/jMkuGI8KDK/bEwWzcT7wlu8e2nROv1B0v
U3qz8YBOSRUp8odOD/jnwd/VHX+yNZj0iVKdvWbXIBEheAS/oYrEMDaUE5NV93AH/xSupGPdEJbd
vjNAYfKBFf/j+TWwEoJktA0bGw1/16IoF/OlvlXQgoYeEbA5974njDQdKoUdSvsKZiwiOzjmUTOu
aNipv+Ip6VQi2su9Fv3oEAuGjHJUnGXKCAXOS9KfximUAZRtcqgPAoo1wTqWigVfOActu22aUmb8
h1HrwBb/OkzlNQhlhm589iLun5lwek4sIN8uzgi4Sb4uzJyyvWvId5F504r8gvePyNOQP1gfI6MX
XJM1PJJOOCfyX+XVXd8hVFwjhBU4fYAlN8k5si+Zs+PTsFb+O/j78hdZ7reWMWR34JcEPGJoBgMg
mUNS0/oRuGWgXry0zivkN9zcoj5laTCSG6Sh22FsW2GnRYFXY2ApHNH2Zw7R/BYPe9V9ofc61qWZ
FkWnosey4O+oKkHLOXWhsbxjFeM5aNYGY89Qta0dBGpAsfQqddlABYeh3NnFk8XuPVfgD9lPDvF/
TkOrzsU1iF3QygEowQEOPDEiwzsBFXnVP9Z9QB/yi3Wh1iW580BwI+0QppDv6Wd8eJuhLQ9tggl9
mPDODSSBZK8n2RkqEh/9KfcLR1iwLTwHTZjStt97Ww/7UM+CicTyQoPIY+k7KdE6PKwMbH6P3xGM
3+f7f0n3+KOV0FfzWuKFYxsWn0FwfLCYZZoKcPr7y9qGDnimaiJoKTb8YFBZsyvxSfVaSlCndOA9
UdB6QlQ4tfMb/T2TyQ1NUu/t9zqIuAAPiZ+AO1DODTKhZHsu2u56ujkdlbli5YfKxNPnlwnve7QI
i+7aJsqlF+i1EyPs86sZhLsVlRxLJT91OrFZmgP9J7AdTVvrPjyy14s9yX5qwZPatylsqobVGvQn
V1lMJMFEBMskZ3DhuDpIAPpU+7jmCBJYZ85GF+IWcLUc4oe+7wCIUhfp7lPmQp4ugW0ac6R6+eAd
5I3fruA8d0yvOgZXcaK5zcfnrnf4BgOm95IQogjQ3FbYNo6xHqJUi3iCq0r9753eP+ncRKKh0scP
AynCqHMz+1GmR9Kv/JKrqNlHLfrIB+6LLC5u/5Wc5BPGvFSNXPTUdkLmahDtMqK5M7ux80goTSn4
AiTTXl+cMQTTJF8LvBmQpowuwjNCbljfmgbFV39g+EZrAOgmCZA4i3YqWG0/tnR/0ks5ANxVLD5a
p+keYAfR6eLrnrO0mm5OPxnIIHg71BPwyI5K7QXrjcOK5daGqK+xSjchhUEP0OHK3RxIZo9M8Q2D
07eq/+zB0qNZuUjStiwzBTb8XoK1AYOWWn7GPOuNohbT6Yvj/oX7LptmYY65ExRPzTFD8IYp7hZn
tc+/x3zP6w9LVQV+2ppJJfJ2Ak9IsK2ocTjZISeymtz+8CJrA9hyTcpccCqikltTilCcVoUbZmoJ
jbZtcMLmDTLnqvKXsx2kp14NeJv6YrOWIqk1Lf0XAtq4F9+e64ZCcENkQGN2fZqbdc/4H0g9bmBN
s6+5ln0T/nXwGvs4KkzSAn4YnN2IAn6YWBgejSCwjyH1P7QgUU10as1YfblifSNoshbzagSS6ArP
pvX/7bg5kTQVq7BtXtDhk/GWYKbYURWobSv1bsYKbUXn1vly2BvSNXc1T7xG6eijPNBnpCPY9P0c
jG52KPiIrVqB6VW+YyC4TwxnAuc5BkVPIx3jniHmbRkQGbghqK0U0hTe+GCunNDph+p5wZUorkK7
JiKBEst35vfH2YvhvhUDJq0ABuXCEaBHg5jiLBwvQNGsogyOJFn+7IcOQpHI7RoGjeYoxuyA4atR
rKBTHA4THZymfvVUsZO95b3eNftAJhxoj5/SVCsn/aVPzeiaXtDhLE2gV8AHYScGxdTIn5w+OLrs
OgMgCBp5I3ApReIuA+LpULNFfcrRBRzQ2MivXRT/FZKI1kBQpjCxiHnIeybXUs3A0MK796SsHaLE
sznNn8hzJdmENrgaY2K0v4EJti0wUFq9Re74PtRcDeHnKE9nMiMqLgsA1me94V8fyCbzpOvBjjp0
aLnkVCWdZJgwISVnAh5x/ecKgoWmjSke9+S/H/YBh2B8SXNZda7orT72CqFzEV2X2oJeDESgocmD
O5Hw1vOEt2rt/loEQamDyH9ypSJaxY2MtMu+LondVrTBkQ5dbrSBqL5IM7QCbuk276jNCo35YuTh
bFNr+swgcne6i+zreuWfwqRsJtOEXECD3wgkSZ0pifHUhSKZ75SO0CiFUY/Xp68bATaSakYFrLcN
+Ss0K60jJ9fkZkvzmBaXg+Q+XcajQrVO37KGKhx4G3G5nOoiXG1rENT4xiPl3yh7cwNeWMnEcGee
FgiAHpi+s21W6b74443wH3/cV/OlC1EGNXhYqce6RikDvWAx2ghhN2I83zF16diADOYLPC2MStJg
ZvAO9lD/E4Pt/lea52Iw4IfU+ENKJWcklBUVfA6hwrQItd1w/nX9M/9p+2VVq0wksmmlKkAQ3dHn
j1mea2X9a4vY/UkMg4JSJ38P353uI2YvYNdvI+s0JxAYUGiQxaCq2bxxXn0VQEDqZpNN17JRTBNH
s00Y2nkNW/chECO5ildMuP1FFq5FRbEQMIry4Uw/AIYw0nBlobhigUtG+BBYp6DsWlw4wNRkA5Pv
e4vEuf6asVeiQKCqeX7WtJzUUbv1cMObj/358Qms4u98mBJV7irs15Iqdxf+xLFcgo9bFKUZ6F+J
IXjZLeWPDDgLa9l3QaV2OihdRSxxn9diFmAP2qQcXPdRHLO3duFNSdSznZm+sSGFnmhvU3+4RLB9
clq4sTjHzx4GJV6YY1oPmqS2Mgw8mpnAV91OCIsZqAxdko0xO/sDMr3JhuDgJ/XZeNvWfswv7UgS
iCFyupJOa1Hn5QK2+IIeEkdrutdG08OxCINmmMqlSK7Aud7xTmAwJNrRq/Hl1u/L6hoGIb+dveqn
3PzBhYZaKQ5E7ix15zmLSl6BhzWQ+APYZ+XhNcNwQfTUIJrHtN1DsCtdWPZ7dZ4eREPYTREDJ3e0
5Qhqb7RMSdWfkHIPV9u8BsHDSwxPerbG4R7ZNKodjjRmfagyN3bbVU64WKpLcO2Pb1KLOnN9siUh
J8fuovRzOWtizhN1gDyk0Rd/QayL8ZcenLaCAGO2ESjNOkPAfCxllIdew1PQh0pSTHiXf7ARsuCg
E1OUtn1XUFWZfwocI3rRK8Q3nZfCQGIEBhyD8zd6LBT50LPSTTj8cAjSXLNSvx7iES7SsxzpeJK7
9VBCet2MSDemTO5IRNcEccVxmdGR4sMvrToBmcIBBYWGNCiaI12/G0ouK0OV5i7QLqsltQnJF7Eu
/Hu7PNCNRRh7kKt++HqeoiiZYqzq/S2X4lVXuS2wxew0X9EQJOXhmAo3LZTwxytG67yG5ybkklzL
ydrd4XQskjMCvZy9B4JxVAAnrVWLznQ//ro+39cg3Glk8Unqr4fU/3mwsdZ7RnBKxgDp9mz6zllJ
btR0RBKLasl2M9kn8D3qWu/aIW3JG/uVADuwVyMwZnleDXF1ea/aKo6bJwrtd8NLtVFCatrUEU74
wAazY0L8N5+EGGQQ/GL8pCBGwG61uQBDo023kaHfdP2KVria44ard9PQARHdfltWjAKzXOmo1Cw9
Hq2UZ0YGiyHCkycJ2e+3KfHVFNO+44HiR+EzOOAc6LSysPVxiCcYn4apRhkMvgTqsGMqjFv+2fyR
9QrlX+BMcy7WVBar8Vj4rkj1GxCChhM9NbNhRK+2CWN1/eohsehXxCByWiZjRFnydwvtOfCIGYe5
slfi3+dl19gNstbcTatWTLhPNHZdtVrIOM+Gk+1AvmR0SBF55oL9U8iY6I57+uevz+xLr/SMmiQR
hPpCvK3UC+N6U1j5PGDYCG5VNiOUZzWfV5NFo+QIuKJiTctMe10mRQ77zEhNxjEFHv2ezqE0X+m1
megzwXyGdT+eQJ+hQA1/0ZqyhZZHXbznTYcn8PSgL7zD0bamC2wFr7YMF3GKJnOANxYPdv53RpUd
nBewtDeluEkZzk/olbSP8yvnE/dHLgI4vl3D4KJ9lBy3tbLkojRkf319kRcotDLXb4yb/cbngyi5
3FBqGHTKgWekt7t1ayJcOiInizHyGWPXOVW+Lt0f3QVtiJjgvDWhD8ldse3Jh7hcV5OGpA/teTgG
50Mv+4VXGH54u+3YaBBmwCGn4KBCU15UWBtZlGTaEoXZF5cZtv81wloLfS143Kpujn9D31Z/zDtO
2Z/I9hwDxpYdBRLvsQZhwl4ZAEm9IWxMyoB6DDx2Ici38C4vMIBuLzDrFGKx1e0wnOCLVNC57PTu
m1dogmJkfIRbsmRnB6S4U7gqv56GC8zlNLKuavgjpg0jULCuVHhtjlQPYH6kLf6mNZMd4AuZoG3J
U+IJh5SFFlQOspFzYI8idb2YM1ScmelY/eiMvGfArsifG7ZHw5XER7yFXBriOreVa2w/XduxpQPb
OVhoKlXBY9lqNSWmBab7TI0re8gRV5VuiOFkRqMdeEIMVXKHkCD1wxZaC2eggmkkkN5Y2U9ff4gC
tCAmEpOzvAyHIXPnDcAjcyI5q/55juh4fn1SDaa80LNDIkKWz7pXPdzJ+TtwYx27slP3qBm4Z9+x
fklGj8ZKm4ophXN0fWBwRr6jxwMndv5agmmvn79gu0hrDgrUGLvZypU+Yw3Uma15RVVKJW82Zrh6
SdT8RKfImGsp6O4ubOr3tum58e2SBni9JiO7UeuS2MOLUcs9XDB4x4WE/BWyjPFLkvBsgcyVO1Si
YsVhrSoUKCIpZn3Wn+xNwClAZqrC0d3DBCNrhKcIBv2OrBobJjUH4YBx1Sp2e6fMAtyFWQoyhsFW
ekzK5hYAhqATjiws/y7OVsHrI/EBWzU5HWJWabDSOcSfZGqwgAgz92LMVqrtP7bLV+y2E1V+Z/hW
0NTKj7+90rn+h3Ui8eNBg9N59jNXxAyoAgCVvgSDteOiHlWbu0eljDhba3Y3SwAaVqRX1culPYGn
xGICYMJH+3vuvkWrp/JhzOJQQxv4efGexCO5OhiwuhFKTOOGefLDWG+2tVedtKKHHa22/oKaAGl7
IAa9MOs/oLupNPL1UtSUbP2EE7Pd+OFCa4kmcsnqWOkdr1pQUBgBp9a4HbyYHQcTf6ECYkQLgWnQ
M77HUDjfILRomnfwZELW71azXvI0HdEVsYw6fulWOM9m6rQtd7mzG9W9WvQi8S2aXzGupbJyJyvM
nBBKZGDVcDN1W5x1FKWlBzorkgzdU/dzxOnbZGqxYVI44sXH9JNcqsKScAMbqPvDUNauZO9YMnTg
e+HsxprX58hSBeeC2qXT3aq1NlDL5BZenICPfhkQ2Ix6K+sCou7pml+Zlboc0+4nCY0NfSYu4E4C
+DE0AjHyPUcep9cJgpd3tZ9i/lJjuVrTPT7IlXOmh05OA1FqYo+hG7hV0b716gPgVo+LQOrTQeJ0
y4jSXQE8/cxr/TyBa3ZaWjw6eLk9lGERFlt6i3TSPzXM1Ucgbd2O7vThdCwKcm+LthZCV+45iNRv
b/1jojpyfu2ryyS3lgv4jwGYNQHYx5q+6lxCll9YeyrijrFuVeTItxtn0fO3hH2ywDYSAEpWqAhN
bccKNvxHrvxXRiM06Qwb6xDrVyj+IkLLjuHngOkdDqP6VOu5LnsEEsKxoEx+nfFk3mG0OoAJ6598
BBfbyLsA3eBnmET71BfinWX4LqeIfvMcwoH7ng8i14d/cVfavW6UAoL/N8AQ64BfalOGaOqF/fne
IDJJHKthgjLb/WOp3qiryHTMD0ukPU7W+h7FDwu8V1n9+2bvyd8K3Ey0c0L5ucfIRg11c2WMsGPd
jIvCOveuMho9UUc96T7O9N/cipQFEVsxPY5+rON4qODpZudA0waGtgRX6bQs4XQLAIL1DzaibdMN
/dZTDw0DC57OpT2SL4n2x3i78lBqAIlNIHApodNENtbCAAn92HjNOVHxQ9sfyfktiFHHCiMXBZZj
pgCofLoGJo1hzmlbpVbZypXSSMJn3fjVVCOofDblpwbPv6Ej5TY2eZb4Hyf609o7FqtQ8sJzQdVs
o0nmdNgv8VMmlY/Loh3G8apgLN4zDjdHZwSThiyBxCaJgmFJgQbL36jHbVhz75ugXGzJUn1On76k
19V7Cd5H5PIHjEfWJz89+93NjFC9GjKTJ6RbVZVPdxwSBBQu8MXbdjbHrcgcf7y1pEBFYGi/Vw7i
AsCvsOOrrXwM3Yc8GwWKTfvCLxDoghvQ2fSh0iQSGDIgBCFNqEHM7xRRMFqtQrrC2imfSfwBfvtG
G04N8K5X3HNBQ/5REKt1oljf98cjUPdRBVreZG8lENUWXAZc1VbdXsbN9FDF5E+cl1w+2Rqp6evt
/0arvYUGBQg9EZ7QNqhIl2OT7+OFXL1e1jsfOSduR79NbQN+gw20AYhFF8fUgb7pqYHjE9aYB7z2
uLh9/ledMGJznCNfbf7fzX9G7wQL1rfZnYMrmg3Wj2lAJWZjAJe9I337jz7exk2i+js9gPZNnKt4
a8dZFDuVH2TUQXaqPjnKaAUydP6YEEzPJyVXQ0WO4cBe7wTdFndm/ShlqaxtIqeQ4hDBDsnQgvLs
pAf8AnQmnf85IoYLN9QIVxgpDeRNDz6Db4OaHVCZx7RofQfgoMOAI4GmgiQuxNVhJIpRGmUV+/EE
zY65IzgeABBMpkJAajcugZIgMBZuResFeGluDsiYecOoM4RYOV9xaQlk7+G2CrDxzvoCh77f8oWR
OJMs33YWVp5psCHADxOHOk7La1T8v3/tQd4wCNXIV9FPhpPvK6gfK7p7BJpYAHD5arcu0S3Qw4XG
KDZ67lJCXg9E5puhU4DAcI7NOk1VaSNprYo5jEL8+y+9apDc6H8EnarhBX3uQBmqnffiu6Z+O1JG
mGrFcLUArku2I/ipST8iNGcXGl5oPyItK7ESov2gGqkSz82YjYQy+FWYHvkWFcJxYkUt7+aa9Uy8
RjDliMSSV9JpJ70GR2ug0BgZpth41QuwBH4sxYFB1Xa1zkn4X23jKq5B5g8E3VL8c5m+hyF73Stc
jBSVDENFf8QimteK5QLyZ0fWZxaupnPRlm6hH7gQ9O6BZv6Eu4sXBoVi4UPCBOTrS3rHq9RZCvSN
GK1t3kfpxyeiREI8R/53I2eMELvSd8m+uGXJCV4xqE94GMTTKhvv0D5+F+Z67jalgz7W6DREgFa0
WaKgg+q+9yLnxL/JOboJ67fmfRN15TJbkIuGIxY0JSmUG6QnHvywD7aG8W3dEh8BY5skcjHrAKxs
dvX8ZFhHGbQ91QH3AwKBSViZGSXB+/cwJc9vivw3vTiARKBmmoBmWAones5bhgvaFz6XZ6zRqpkV
dpa7HtYzpVyxJtM85KYxZ6w8i60qQ4BhutAHeO7O4+XaLCZjA9riqDTfvVUpS77dAHAKbSLvWcvN
8xDDYg+TYFsGL83Sz1BOAKV4H3vdWyxX/wkxOjVCJxN9WPXhTwpOSiZjI2FHwLJhZls+ZQ0s3e0Z
3gC/lyc1q0XsDfVE5Jh9V9Mw4IfKf5dW/l8yb8GyD/YeVSYxgHw8cZ0jK+7MHKBL+cbp8h7FCXDL
qXcYLBlQxwqe/ZDrBkeRtsSFHGkd40Bib/DMGfYZlQuyFfRsbJQGMNl0mwSI8NimSE5+U2TzB4HN
OQLWpXUtriHLhu8QM43cc5ymj4ZyWtCri26nT4v/uda0ZOXqpovoUNBouAAsZ7eIv9U4SIQDPylm
s4VNMQhXeyEKuJ8hk22RyFFy3Z41NrTDvth5CnkJ5WeF1mL4bTOhzPLjwUz9z2yzumW5ZFas7+3y
S0/670TPbO9xSVySAVbBh7Bi5IcKzYjaia6QX8L8pnYOQrUMKvaIbLsCMk9v9ITUp4Sz4njPqOFP
Emd8kTNyf7/wI4Axf5uKf7SqIZwAb7GWthqZaJyCB+lRE+6AUa4dYY0faTvP35GMEloZqSrAL6eg
HhO0TI5QDPb8BCs1W/wqDgN/STG7PWegL7LNaK7XiCmNPsSaH0e1KXJm/xv70iVdUGgzuF/Pu1DX
End8xhXen/UNzG/3ZDdcdMRJBaSKVPuImfEsQukWGDTpsqcHw5Xko/WvvxWt4VD8w5XJ8yHZKC+L
Adj15Dh43X5albM/X4IOPVaaANgqEL0aWT8V6m10EltmM603KVdASup8iQEKp7MsR45TstRrwmZr
XvaeMddAUJKsSyaCW8OBFHuLX5WbEM/PW/DUvw7pkIJOlzaASwrh5no3y7SKbHmSxKzMtn5HiNqM
++AvJqC4suMs41ziQdc+D16PFtAEi+atAaW4xuNXBZNeFMMEqTuhBI+jMe2ESvKrQ8BRK7Y5IfRL
rOW9tsHe5uxemhDfA5MELbZRm/NhtYRHAliLMc2U6lwhF/SwNEYNxpVtbTaF1i9rxctK3VomJxrr
sUhBByhYJwY8NW8YaYUCcPvaDw3A9/s9Pzb5IQQjOeqxcA86KaSCtaVjL6KuLoueEohb39+kk/M0
+dIiB6Aer9pIjsqdbFzJhY1kAZ/VpsaeDkz8oQ0zCCwy05Yif82pDMKEgdS4XRYnI1HP5oVS5mBM
okCQZe04psHfSVenUhxEZqTr1eoi4reFcecounOckEEloTRMeHPZPm8G+Wuns30zM4VcXAvM1vux
dbUMXH0lUdanOxCsVyETLTgPFExdNg8bg+M298qzvWyPdJ1cX4FXE6OmKQB48e8kM0bUIvRb2Apx
JvqHYjiMww0CDsULLZGh90T5FMd0mnPWz4/r99yTiKv21ojlw4dvEC+Byi992bKCTt1Ut1a8Tqk6
0SXpiyq8/mhxIXYxUDeNvm6E/iiTo6ofCOAbie4NNrb3U99k6ctOoIPiLedJ/rmk9KCWM9eNVw0a
a1g8XYNMghptxztVzrMNlwPBKWLWDuMAHCrVgCXZvvNDWqvuBbx/886XqVu9ys5ImUfj6oTHqj3+
d1OqG+m04HC2ExHeef7pHeFaUA0dMhJlhYeduzTfU6h3EmCaFjij0FSg+E5lb8sBJ+HphA0j3MTm
3z8COjcwM0LC7y0RuHo1mhfMO8R9NEAn6cy5JllFZ9fLRfGtKLGljf6v2muPkdMZg67CrCnI/gBV
O2n5qUSwTBOmvQoE25X/vSfqcIbRYc8PIjZBre/WqmKDuaSyrvn6fehbORlTVMVOWrnqNJDLEpch
8M/L6ZD+KXTtQYtEfxEs3hPu1dwUNnDHmyqCKDFpxS916XK2kBLGDl89x/BSRyFuDlfOmc92gcQy
S303XwsTIzJKJ2ICIr8PZitOI92w/RmErzmF5L2hvHQO9I9QhhIZ9p4ASC6i1FmQ72cH2QTvse/D
A4VOig+54BLRdMJw/ZFeSanyr18jal3PvZNNXx1wH1Dl+PZmYws7SgxtrHCAEuMiwYDob6WP/Mj1
IXK4IwUNwYuoLNCHNgQsAVMh+33ugI5V9+h1tnwHDOymxZ8c41h/UWHZozNVnm9pi+RMJSS5W8C5
6gs6Hmg0mb/qOxnUiYYnsMR3PlckGeZ8pRiwaEV5cNqzig/IElPf/6B1CKvKECz5mmUNN8SfH300
Xh/dpK+BtAI/o294qsGUdjggDcZH+pPawElDSqOlqlFEZZWzRn6tFrgaDe+Dc358SpE7u4op1XrK
C+91pZqWUxITGagultDCI8yrbg0nnfAOyqPEVRExnsJqbfTiUbbi2FmJgC7s0fHcI6a0CTFG+X1i
BWH5UoIqXrFV5T0NVYPVaj4LzvjgauI+KblK6MYfOUm5gzT3ao+Z1CQUmdAJn+7SVnVdCY7dTSRz
MrQf7GtysHZfg/joAXChZiWYCxGNcwk2RC9Wv+MR+m2aQUWuALBGK110XJYTv/Ay7eZBtuTQILG8
WuoalRqU/W6rF+w4HvjGSnzTfn0i4CrygMHRuBlYMmGCJDlSvazYslwat9XKfnk3w8ihnuqeXE8U
2Pz/MBOQtUbw4TRw/KwfnuyolKl7oZOnEafwnvWjM39DM0SfVwFsapL6aifZbFEO0baz6EiIKh5l
Pmc51ClAv9JwiZp52w6sYmYwCqUXTF8rTHPCE41/USv6PQyh8o4V/p7+1JRFXvoFm07M883lMILQ
S5zv38Ke1URESFUEOn1fb75huwhNqcKwcSSERtTeghCz/+LRH6YtoCO+lS996k+fg9kd4PkXKJP3
p4g9ZdCBSI/OYo08LWT/5Kw50s3WKHeEwyG5NSyiagmpiVSNV8IH5xeJaGkvhk4OC4bffZg54IcG
YrgLcNYkEgSOrjBF4C/G2SkdvOXTFZmQZ0LhA7Z6oKhxwFtV26SiV0BbqLWn1ydgZy9CjWsGDSL2
ge494FS2Djj2tyNUBfO2ThzlHyUagEsR6msd5/U97nR/azv2KTQnXyDjm19LdY7+bZ2HOjZ3TeYJ
pCUcZ+3btqu7irJawxMFX93WRupYidFk3vttmgRI92tdbYSiNYaJrD0MV6JioOiJIsJcH2rGmdzE
r54YFO5e3JdrgMX1Ch8NzjRL/qnJSphgz6mY9i7HNDlxkQrmL57zJS0EwRBM7VtkotKe2xztOYOb
JEyLwPk9po8OsGxnDOVLETLj0rJeDUz2J8jMCt8fYnIOYH1qKKo94r9wCANbAy/d5mYBsanHiHdU
xibmQcBf/E1vcdEAlOUKOjkuF293wBzTeG5xhOVN+DZP0s6XBR/cw8pqK9b8cgPvxjqxhNorrkt3
ciJlX7kJ+ZkF5cP5yX2PjPqh3ryUn5MkVPx8tN7dtkgs8EqR1N6jYcl6gv1WyBGNoHgexLoZ0ViW
wJ2rzM49lRH5HBfJBfS6sWvr3bxF53MGvS7YcG+DgGXJX3vjqEM94AzKA9/nFX/hojFBhcVgTNEn
IUWnP9s2nmA/Tvf1cDuWU4JCWzPXuDEQ0Op7M3m5AFQtXeD6IBoAJWKYctMgN+2xPx5XNpCHQGaO
5w7RxvxOByywxihYxBiEDyqk4pkPZ3XvmjU/C9h0bJAzKdwVGvrCZ5N8qZdSkZk6gcV84OAnU9ox
Lvl8EhO/zcl3EG78E735RSmHj6lp4HGLUhn0itWGsFXhudc2ph8ZyIFjy3rb4OK0h0jwv8boW0jw
WUiHlfoG8doJse/uWRGWScTQR+DmeoiZNW11NS0mUGMgxUk6dxiC8hMSpuXUYCVXcKXaIL89X3Mq
F7qohQMn/FGZsRTLq5SWLIDHL+XfN3/wsk3elkhMLfKuNeRXRZy5rlpRS5y0daRGi3AV3v/VsNtX
GhonNRbenjoCiClfxP5zvTzFE8WDaRLiFBhxMrbsvKpg/eGRWC5p8pf3K5znW3+m0NmAj7QhmGfm
cZ5YUc19q0Mj7k201nYKr6bhIycReUqwl6QlyO5dD1U4yu/EWd4m152Tw5skUPYmtDmW2Mz9oQXi
2IwdOk55VsjZoVquN12POhr/zwmMv3WoDthf/gJeMRzhRcqH44NRN1pzOqBKm0OGE33IE7uXCEuD
akJ8W81giBJWnAJapCJJXSTMFWXatuqECaHikeXtU55sGhxG+gJfLk0MXlD+o82ZGzlnL5wU7xHe
LWZQqDKlxVbfrsp2NhLOtUxLODJmtGRavIX+JeXrQMt5g12lXn7jMaCEDuXxXwXXHwUkP2raUoKV
SAYEmYSms3i1VxkvJvk8EUOHwS7EFjj9s5dDU7R09D5v3tV+tC7bwK9+j515gDXhvGru3PiekO5j
RQ40GYRgybDZyS2zVd5lIj+bviUqS5muBHf1IyZe0IQnx2uTen1sLPqHbD/9G4alCGwQTr3Q5Std
cP7T9J4Y9DM4rXUcqN5RA0jxA518wWfbqMi7Sr74r3wzdU7Sb8yXXUfVO/8lXlno6bO4SS97UjHi
rmJo4VrLeRsPLIWBRORVRTNKdR0u/P+J/qZHTU6lXlGWpL+HnzcQOa9CqV7oqJRYY6zFmiyTdRZi
Ngme3wVt29wI0AbEKFxKL+h0ps0yKLHC6CQ0L9TiZCIlIAmqolIMYY9+J1BMgXNSWf/ryFcN9BAO
W4Hs+GacubBlcRHyCs3UWbcC9Ps5KfCRbs8Htk+g19RIwYJNuYmzM9cMsmATue0gB28XRLBE4hKm
WEC72PzMYnJUeiYrVt+A6Xxsz2RYVme9+yHc7eyJZ6L/fRwvBGJIyKm1KjKXw2FQXOwtGiK8Apt2
FY4L9h+A+0F/VrSOiCowWlC3j5WinOMK31KYPezZL508Y5578ncjKW1mxS5fWMz8a/uqPtbELnF0
BSkMsHxoZiwdZseVByWLYv8voOnQAewvsIhpIokM6D0kf7zCbrRQLvRv8yBvkVR9mlIqft4MShD2
T1weqAZc1lGH/cf6YoG5jbxbo1QzS1/ECAtd6YzLoHHdW5hWqECeQ00CtjTJni9jjvylME/iNErY
aSdWZ0nxgC0qgvdSSCVQp7sniOmKJD3KI/InU7vzH8eNP3vvwm4rk0FkAsCRQ01VeXrkvrDHsIiz
9jSr4m0UXmw67MQAc3yuCgEbHNNppsiyAjl05/51zj7PCrga95HKDm2gQo9nuI0iU+SABrP/1K6z
8bkpLAYm6jZCH/qhPA0VcBYFYXS2QBDxZLGjyXg7vrb/dyxi9Yu8Pl0tznqIjE3KiA3mqXd4Ag5v
5XeuZVSScWBxArFpg6ixQfzYHuXIkkxbkVUqGUJnOE0XBHfoggmyP2+W/ZSfWzTSAM6jIE2bahEY
3Qofh3u8XxWySBV5b0sRi3FhtW280pWyL45J2ClE3M2M1eHTy7XUF8KbuOPB7bv8OZP4TsvLPD4C
UFLTbxsCv6FB7HWJXzr6/lSIYcE++PrSesXADJbmm7FyhNNHr2YgGORXAdV3ptjOOxstSWQAGHwI
il4WX1gHTfG7OmmErTqVkXNX7sbIvLF0eRxwDKoK5qs9uGZCv7fWhu33TF132uPm3qJp0ZEa8gbQ
5/S2SiTfG7TahCpyTy9yQ36cduz4XstFqkZZ0jG41/ES1RnmBgjbhRW4HrkS8/X5ofBG+pfOC085
ZXtEBiet6P6gVKnip7ztx1k/hB2H80TPZQIqLnvfHV46jozMH1X3+oV5RtuukQxKnd/sZcB2CfGo
1Qf2rLdvguo3ww4k1CycVFEkPimhDvPtjHKH+fbaFkxD9g1nG+ta3+ppEqLpphZuJUUxRbE5Hs8d
9zcyhULwAhni3qypr66+r6VSeQ8wgcx6pRi+kCD4JWxMXv/71RDBf2ZZ+z9dQq3Sxo3cv96i23gk
1Zea19C0LbcNjNOGQE22BIm18RUD4yCmaLF6dmaHyhGzhbQbz/PLBxuOpXnSvKlgCslK05w5VssC
+2t71j0Lb8XS6aR1mP1swpDXN7mmdx+G5FgwBXAekxyxdQJA35vPuJHmmWGyWd8yiXRLsY0AS8/K
Gfn2y+R7oTYQQKD6hxUhNBC1HM6Tjvyp893avMJkxg5Hepw7erXoNo7oFA5pZBmnN7ug4Kocz3Eo
RMpfBE+EwcLKRNaprA86E1wFkURq+oyDV3eUzu2iPnWz/Kct9fkJMhsSNflamWkkIt90ZhuuEGt/
5donIuiQvEmyrQW57hxPT7j+St4GRBNrStiJqRdA/NAaezVSemnPpCHhT/2Uoma7nVfxZ6uO3I7X
otW+jmHuJUcFLlyMEx4sstctNwmxWycMg5daXvXcjL+Xsj+vBnL7kIklks0JK+1Q+expGIgJHK+x
YN0shGMDrNFp1ZlWQjomZARh1/r2JmkmcvmKjT/UD7BDwDLJCGE6dlP+YYlUwo7pSwCNTRh+8l84
TQWYyLvHZNHPCEEhLSEPnPfh/qXmbV9EH8IeqI5qujBp0W9MGqBxQ0anooROSCHwxFE7iDCrHNu4
lisKXvlhFeI1bpSbtIP24VwXVCb7nHPb6Fq5xYFwynXGohgPn4KBKRaWKOhHmuJpQElC/CXbAgJg
oGgDOdXemVwBSPcx3zS3cR89GjP6m+exRjnnBshypOKi8eB3et5cIpLhAnw2V7pWzTsOAjYoGPxk
4iKPWF2AiVNBdTg+7n+E7E/W6RltJwYw+Tb39CG5qxc3dShB7uIIVV0W1733UZ3i9bQH+eqY5grD
9g9J4kG7GmyOv5Mav9teP3tB+zMgjC1bUzQ+pAGMnry6mTkZA1bsxolIHZyJcOdVO787tIvi1qU8
wFwIuqGyn6L5qeKTVS6YIMcF/UOHJDIUe9YP0yYw20srLT8SoNlPfGhJA4Qn9JE0VDDxL0I+NmT1
cF/J2M3Q8I7vgM5S2ar2HBeLxBYSg/CQDDUvBu0sekrfz23IDr0WFRhMQm2kww8XaJEr4o6Gcz1H
XQN8sklWSmQcSGeFhD2KG09dVVggS6ZkheJBrp+5TxI/pY3e5Xc9fXYoPVbiqu8toN0ZTd6C3NGq
Ck0XfZQKMBOJpOxNVASkZM6ZeKzkWpZtol1CJQ2npv96cr12IcU1kQTXF7lCnVZ1w6OD/1EjhcC8
pKU2f4aDUsvXg5UP1Gy+Tkf7oFeKA9NViinXcAALfvJrVoqnRdEV//EsJAOTsWWiNafZCdynzVBS
Qd88ghqvCqf+5tNfpimdms6V7Of8smmmHHV8XC+X+4yS3hTNR6+MiZSYN6bVUkhZyLm7Ld8TXt74
b0VAoHlsqX48tcHfeqBNSIaQAjWjJRye/w6/od4GfdYK6/62ZCTRKrbkKxoObnFRvBitnKql7ypq
FlSphqxJzoEEZabCZL7FbDjitQUfOiyKsPrIqdiwPPfR5ndacbmgbCSPA33TrtlM/J6aVbc2Y0gC
vdUnNBC9eNruXT4WHtMYl61HZtOwFpAM5hAbd8mKsT6j/QBxmiT7vna9S9vxeH6vRvvHyFgW7Efm
v5QosSG9bqF9mOizVcl9uy4LdSkFN8+BBHHUPkd+rF61vTGRnZ9+2WnTZHgpzKB9Put4IW2ITxMP
787keonazaQ4szSisTTAPx2pmTJBkrMap3s9/Tj4gZUhn99xRQuTQnRA0FUQSTJlexy50KKFBESw
D/7eEENXe+0XmdMvZTNnjk6XZid0w3wk+/QGHolXGiZQ7cC8UvY7v41RnNLi/S1Gwt2f7j2PZjB1
a+JWXeA0LWc98D3EFrCASUQ0tLP7yVNjuk+oeFluf5P8s3/4o0Zb8VWm5zjQPMNxmKcNrvRz++BV
NXkM1LNj4Sz8K3ShZt7nVJdTkAlKhdXnefMIRYjl6ImqsbRBdgy2hQ7T7QMkZTKYbvlC05Va2b8L
3C6xrdD4H9lwNgPNsa7L60JCZxXd9BLqnsFWmoYRkSKCWyJmWEPnD3edgCiiCi83Mxc8URIwUkXb
L4biuZxhJb4xegyg1AUwcs9TtICXSzS0Lhro4s7Ba6eHz+SdiM1NFYq8T2khy8N1Y1sMorSi7yxw
wqNO2H8zGvnjver/Vx0Knw+VM0kQS1rwKmHMk09Rdu81rxwLOQhLRUJqMyhdTvvqtICHAC6dTqRJ
E52RqBh7rlSMo4Ldcuhz8cyKbHajaNx4eCx4ePuy6VUpm35Jb+z7BO27wXeIybidtcAObcE28DHP
ItB9bQphHNAIlXEbyzA+JUGCF7BDRZeB1R4TiTgb4oZsY0taLQmjOB/q3je99a+Abfgxj9ZYSsL0
AifOfq38OpiHxZNVSlbk/7QthnI39v1uw65JlzDQM1ei5WxY/crwjpUsJRdxwzegEfabLB1DpJsb
0AMzd0iizupDcgTC7Y/hzCM5OKRm29uWwEYs48nJ9F4jBwC42MXfhdrZ4nCPXNgfLkr4pDIilEtr
byeDS9aOFCl9BDdj984TzUFOvdXfx1l9Bmoh5SmiPUXXWDoyBGS99xlDhJo6kq84jBhrwlZ2JyFY
mkNKStQYIMHcQ9NFoX6hq3cVemZKYQNCOU4ZVIN8EuaEFsVsdtNb691t2mfuWoCv81g2g1bHlDcm
ueUWQQ4hJU0QuVFsVbZjSdENqTlh1pX7XXX/hyvTRY2chOSTRBzn9zGmE+Fu4YVHRbnD7h6PElhW
eiuqawMbGH13zTRfcdC/gdnIApsYh9cv+e7nQUdVn1ft8TSPTKaC2LH9c9z0TD1nNRWozsMGRsss
nzQ2+3DeZyVCwuoTCtiT5bGjrF313xwB3cRBW+ih8Zy/l9DYDB84Nu38d2t7XctOMIiZi9a6xLEv
SqHK/c9+iix1UNkXu1j8FCA4G884SnjdNXFGvmXHgjZP3SubYIzk0VD23EcULXkJR3eEZYjOIeoi
m854QN6nqTcqp+xorPIUmbMgT+6dK5zwb2fJXUulPNLx9XTRwfUIh1jLJM4gQLwHBUfjMZ2mS+8C
YWzDRIOO8I+C9C8j1UxSIa6sueJEWK5W0KUD/SGkHSyF8sQRnJCJN34kBN4GzX3ZIxFtw4tZR2Nj
GSh1j8P5RUbv2d4e+vrbkGwS7CKr4knus5hAAaLn8ppFcuMd7jazwK9ZRFd2sKThk+JU6WxIN7CN
qGJXqnzB/X7KiroZI1646/8OKXjJ34NbvdxdVTTmB352FAqQGTQOIPQCwbSSc9+KEvdtEe4EJ7ac
XNHiDCbSANP3HpCHIHuiZrIbVxgWv0QCQ7qhU2PRZqZ67pZB8aPLSNm8D7ajNN9AxV+3MvDeu2uT
HAjIuffkQv53QeRs9Dk83dq3xZUtBctfgN6aF5/wjSMqHvXBIEsRSkA5iMPHAo2L4YN9HHcuWWTS
i7ogv69VI/LcXgpfafsaaNudKllh6JaPQbuDCpFCprQMQGQeBiD9CmB6y84w7IIzXnAdnpVdETqx
YNW9C9gvZXnso6dRZAUjcIz1xrwQg2XC4XEinr+wGai/JYYv9X6r6dJi4y7Xh34TAVgdIcECaiMQ
SWXpRTeS6Y3v5k2/TJBT8VjC2UzHdC1xSVpusumLYr+MKOQEAPQcWrpA9j+PTF0xNxZZda6g0dH1
4Tq6DNmuoFHaXywqgGLeoFtKmQCJTNXz477bGQYzvfuU7qgJAhavIXcgFbvUltnXMk1pRPEKpRor
4D5w8/+NOEYLpR3KU2kbsPG8rFNFp6Kc9s6Yj8TZTq8haEYsN92H/yhEK7+gDRkTVvDk6Nf2XfxN
31G/81xHphlHZfBxShhOaaFWl9fRgBHIm5vN8t6ahgxeAg1H14xPT2I0AB83tX1tja2DW0Fv+sVt
csxxbclNGy9Pc1kHSeR+L1KH4VLOl/SmGwiXJTKwypRB953TOLZIQq3umzhqnv84WTdfL9gb2Ahx
MOnsiRO6EJ67Fyrppe6oheiluPRPu9o1ZUMnJNjIg8icJLwcvoEzb2fxgRWCvLqjJP6wg/YoSVac
B4FMGYIrSaVEoY0RZKaUX0Rfbf8GSgrRcBbWnDTbK1NXGPV3yMllkxzmGgXEsH/x85BwBLQlViec
JMrSuB6NCQP6T7RnwScOQGGWFXZnMINfm0CyS4boFAkIvT5B75okizfmyesicnVMVAr2q6yCP/Or
LkNqoCoNfdtBSJxGNgTR1y7e4Py1E1wurz9wqsHhVd8DI79G3wHPUqCCPzlA5kqk4Ais8TAUNj85
OyDIhixXKg+nprGhw19Xs0Ui+Eu2UdUq+FK48yUzIDZISF+4m+Tq5/D+DmNaYU+IVbhO7vnOTxmc
gpzQ9S02/3YAOk+U4PaZ94fXIQpmTNwQdA8WZ3SatHb+Yquzvr+F0oh/0clMujBYSLUeY80FAfl/
l37UiFHa4t1Di/i9dNaLnhCIjrj1pP1jGNSq0Tv2CFYI/N7FZAC8mzY/ZaDAPUlZDGy1X7lR2w+O
Dm6uqngAbiFGCFkng6TMoKW6vorUnuPnQh9Jkg/lvqI7fqjkTygfL01fe64m7a8uV1R8cBM1D0tB
5Cye6ZxCTjZLymbYK0JXQkqhqeWeByc6fb+/uNDOFyekwgjSsRKUqbMQwFyQiOjrSRb1Os3negou
xPJ1VyhWDKhyjdj9T/vpAQ77PE7pNXMOZpkTNtQc1bvoMXAiLRI98ixokzojPACxut27NHIhYRbU
7rJEAJCp0VqqrlGU5cyuRewoyM3FxIDiaS42SZZiAKjdm5T2Y4WEpNAaT6Bcs6yyoKu+yr8Vef6m
e6sIU47B5IaorGUzgxsveC2OtxaS2QD+RwD3eva6f9ZcD7eJl2Eyor0bKGOYLLzzMXjYVQbXZ3rS
hV+DXSpKfFEq8xSNfEgQfaiSaH3i42Mune3TsfphQcpiapOALhax0n17+aEfyaLIfJkxg5qHiFVP
Uvauo/6HBsGavw6Q/otNmbPy2mnvzMiDEvQwQyKf2Expti+UHVUajwbEgmqfYzC11uWt8j7K+rYZ
DvvevZNMxYyJybO63qK5ID3ZPSFcLqbrKouj0PA4WVwUeQTLtz0+IO+4Cih7P8JmFMu6+ilt6hQw
r3CeykNvrT6i0MM11agD6sFqDUlxFBQa0rV6BvXTJx1ic5T9yo4ZTTzapGMUAbjdcexY5dooJgF1
bWasWXRi+71Jt8WP+qNX7B5P6E5kUAH/Kebw/P/H8X+qqd7oqBvTChXk1oxFoIWKRRRR+UR4BvWg
yQv95c4ECf0qiaESlDeJ/9t2KzajjgBH1MVhtiC0NHkY0diAUYVMwp8ei4liiVL2GNnfniWM73MW
uOJBwBbgbHK6R++7kwogKKze0jIjpH3E7r/ZGjDAnOTv5qAi0ZQHsHxN/nqZfhptUm6Fuf2VJ8gs
R4HmjkSzNHYIRV+iCsrjEgXxiXzj+UHWrNaeFlgo/4+RsUdbVwPLwSOqL74dE7DhFA8/Fgpn0YE3
lJf8iFAoq/DWzGdgv5lwBfQjTuyM4KjX3AVF7ybuifBYsmsofVaLV28fAnFSgZ9/ll5VNvMgWSU4
0xV4fNVViqUr65wJFmSmJ7R9e5UlbEyVwRg3sGx1gW4LkrGVzzyyTdEQ7db1tgDtRNEAGWJD9C8q
oCxuoBs1e/DArZTAIW6h1lZFpR5NEyKKCMhIJyuc+D75F9EttKGfIQC27sXHfbKpaWHrv9MlaXDy
FTxH2DO+62AMj8yRJWQaBwwGb9fBY7tvWKAq/dNCuivLZDoDNEZpwqjsQolhYKLGrng9NPkB7sJj
SzjmCrp9K2mXgYYDCrHKsypPK8+wWZkqeT0n/cvtjMAggeqQjAZLe7NRb+LZR6/CIBlHAE3rE0bD
HwMZXmws7CWVitI/3gd1uxV7pY+OUpGZ6hVGgUOqVfbNU5dabJiN50P2YSE76LkCz5qMhVYUD1D+
+NQG3+s/m/O+KfVVeLxBXjX/801n7MD/1YsClTD7V8QSCsgQNYOulJ3upTARNtWlLFVyx3wbLbe5
13QJyNlXGpFTJ0bKW3mbfjVNHpLPOsQs4AkaPnmvpzbe55ehDf79v2e6t4qxt4OQ8MPoG7a2ui52
MxP2wxnHZxd0aZhjZEmXW/fZGQL+GnVLj7nRBrar4A0/sNF7Q1kftUiDhojkNsgy4AAwMfVB5zvE
8EQ1WpwSY5U02eXHlDdPc/8Pma4ctDhLOVeEq4JQN6XU3N1mHCoSbkBE+6dm3b1BSf4eF4P1GJB5
jX13g/89tDJ03fRZa+BYnWklE7epHOYk5lXyDtl7tmwIUqbF2AFL/opBlbdxEi6jm5tucFEWb4js
04yBAbNKgF4y2A1wdDXi9YB40FlalaG58/i6lLCXkctJ3CxSf0EFtcFMhwdYPYS4ffiN6Ub1A6Od
lLrCX6ZdKyzfhcvt4Q4ADzSo1zvq0Po7NCYfA4OxO3WAenUL+A3ZbanmYNURW+pymLLsWiGy3NW/
bMolUCHlNNyq9AyWCNcpHVTdZYRyx7ElJqzc6+V1X/Djj1DMlpYpHTblmN4zIydxMLTxMrwMRp0e
Tf3TsrK5Z3OXZlCy5ILD7R0D6BmQLG+p3nhIrHiHRe9SMgqHEjFz3k8kvztqMIoWSZ15m7hAE64U
aUXQ/J4mSFtPzsBaBS4Eyvds4+HLSRUkUkaFfOM/BiEa73Uoq7guXVZBtwVJmzZtx+R6MDofT+XS
Vp0WwxiNwnt6XrwQCuOsGBcCZQ1NoDeOMGS9kZk9frhcPhPH0NlGiLTJnwmpkaHGJreomRZds4QB
a0UQlYXpSodQsKUa4cq2kudf3G45bxncY98bwam/9lxrJJ5ZGgEcAW4UNC7ralz8gnQgMtBEfqBi
8vopFqOea5oOXorrIvoGpwLyHP34XqSbNBKyfuhLN+DpjsucOkerp/E7IIsUsssqj/jqrgdYvM7a
bNa2fuKz7xdFf5BFW0VgXMcnP/oPn//51mPpOXBFF0KhiS/DzYfGkOKnTmdWK7SDzPpRLpZ8WERp
H7EFnNhdFxw9+hEZg9gu2mC50phiITaKBlOxUsDJziwV/HqsBtkbjGgCn8A+YeOWtoeN0NNHYwts
ZFK0fE10g75O/9/kjTmIr2hq4lo4De24a4cehg7P9M1P4eFcS0NCMZSw0zB9xnh4/PiYY/oLltah
V9h0jwPSUfYolWpPNn6Z8xKkTooyrsRgRqofjUcfxlBNcrbksoHf83ZmOAAvIpbWuLAUBbPNPtZC
KslDiQDoxiXebrJbkMwZrzOGRdPq73u/+0EhXdXVlATQEAh9lkSFnuRdl8MlqEOsUPK1CPzrpF4o
A8IPpTEuT8Wzri465bG83JeTddAwp8opwUSrDUoYyQbqm4ZBygiB6vUMHj+fodKQiV/AeYRW2/Hf
qDogUSHaCWjdGPETLs+wg74bRpksvoXaKjGE5z7XlJJEorvA7/6ujeCfBcSp5cyp9YE1uZ3ezHlV
v+LJVehF6tDQnohIQpYQr3q/7uoQeGtwIa6fN7n0cuRIJdGznNEpYx6bSRu0CFgxnjlHLe2pP1p5
CXCD+nXo9d9rAGDQB4NBn/7G0h6AgMPAFPTKj5E3tXjWKfGziRsJLgm2c1Ix0+czU2avmLO+Wg+D
4MZsi1nwhMPuSLu/LQh5TvJvQ6JlvUqTjzPL8cPnTaxYT8YeIDvLhysJo3tiuvwOQLeM75CcUt92
HD+w1xMrwN09JnBtXL8aGCpanovXRaHExiWEFvY44ao/2+A8c6dBxTlQIeORJxebbTduwvBARvSr
jORnU7MyuCnVzub7bxTY3rI5Oy67i3dkBqV6e+G8qReN48MjY3LDS0l4/45e8TCCVIoqxJglWQ+u
c5UL9WqM2ECOlH8j7ZCt+YPzFWEVV7D3jNzqmuRGzrvEa3UkOmC+qs8z4Ix0g9vFFVSpNeRNc/e2
Y3/RExxp71s4y6YEPndiis8sMSfkwWIzjVFrHmBXFIYLygwi1ef9KBejUWQNhcKcoa7nWZx9LuBq
pKxXIbuytlzg8Bm7r6Q34PSafv3qJmSNlKDakuLBlcbPB9L6uVqfb5lcKlEIyVVuZvjMLypGPkAf
HjWjdnBaOM63pNPE3H2Wx6akVNMTgIfymZRiZxCqp2Acha8/ecCJs5yJAjEGbRbJLGuZKlrTxdHu
e/D4vxmkjwYHT4dzzLd7j4UYRPy4aVw1LIB3Vuuba7FZvDz/pG9Net7XXQ4m0kgN1FUIKiU7W+g9
s0ouYHIObmgNoo0pLOhZG+O1sn9rMJO60WzGTYT8I0dQA+iCn9woj2pFPzgJgr4/KI7KNd6TC2LR
py/IneKhdULJYbWmZl3Y+YczAwQn3TnWO9cUOYlXtHifg3aHUUhuWcge+yhuvuRcZvrrRkZbk1OM
ADeNibl6Xi922t+zhrc+9LGnXCOO841HvK7lUdY6rug4i8PWOCOmDwlJmxmkuMA63OxKZLcoioQb
J86AuktNa4uavyQ3Us1FUEfocraA+ZZCoqK9toIAtTWpucCWVUtfsBiVDsdC/oaBm43F4WYz6bvp
yg/i12KCvXh5ASD23EOSPKwwsIm0oOmUXdwwhHeJP4U4Xv94gbs97vgyGx1ycR324d+ow3T/L4Jx
8s60n8lcIPvhYKbjZ5LA5BmVQkt+6p0tgMX+q4t7Pb6jqvk9b3g4E3bolnde5pCU3L8T+oQfepAF
sDfqGdm//BNEnpdIHee6C333xAJGAkA1mADRDpzHV1/cjuqK0u910sOljuWhBuxWslbm7pU81ksb
nCRgb+qtVUc28ohYzQERAhFIhK4qUfJvQtWJ1BSCUngG1YiYzourwj6VtPmHaXFIypaaViT77CX2
x7+HpP6+H334UzFTqKrzOuZ74IBsp/N6UrVCfJnnKBsDCS/uAo7bRRqmfW6hrE7AKRPBf9uOruqZ
vRuzmEaVnfZLACSTXBUD6u/+HEsXkjl07vBISyQAwoVbhf3xvjyLu0pAG+F3KHtUy6gs3IJgkGtB
CRA3uZhKh4SeW81gpig/4M8Q9fJYDg3ESzIAsDApagvnf9C8ASWQuJ4IpZ1yVxeGIzYWWbVYsA/l
jdOjRLCYEc9fZpMyJLbCilCm/gQhG/LBAfKrMsxVKHpG8IKd+vtX8eK+HAofdlsCFQ0xvlDfwxNq
TYA7EAdg7bNaEtQpVcW4/93IIOtSeHkuTz/mt55HfqKuFCdaA0gHeQnlwnJ8M4oVAhpJZa85gzru
/lH8z4BjuM4PRoaJ1MsiM1OELZ9aVru4SswSxEcNc0/MbaXQRtHRGLV5W7tYFeqvjPpJ35LUxoKf
mH/mIeJfPG5nkx3jeTD3JzESLZdVwQuVNE+ML+apVpW/I7Ec1fvRbiTsJANnMSH/W2kdS2khz3Fc
3N5eorALfV9KCCkMOXQKdeujmP6hnvUlKpk5KgycORefjjS65hMHlVzEL1py4ps6OlKFgYHDucNr
t2QM6cClA3APXxFterN3XV8m6JT2RRhKEM6BaIcK/9YChpCYvLouW2o9v9l2rylwUw2X8nVCXTK6
mQf+wuEUkV9FMdCBM9vu9oPW+z8JXKEsMD4yyC7T+yBJHkb8wv50NvGCMG3iqonNLlRQozscAfQ/
4sbI7OPRZOJ1bQnga4ksGVQ375ksiRbGlZE2nrsjf0vOL2tI9b4pFFg43g+V0FsusRsaAUlXjLpR
FHtwX8f3ar0Au3E8e9ZFdhaKduw2tUkkLYTensHovsSYuxDpFNbDDQNGuyLO3tqIeiy+n7ya0zy+
0ZjDepPAAoA2pVuqGtDc2n+DKoYDM3ZPlttDiHGAq9nkdjl+mMVPLcNBbTFgLXOK5KjG9jNhgnaY
7kYAvqDhZ6g6U5nvwty6soSZKWierNqL5Fo0Rhe0I6+JXhMmcjNw8aOi/a+rG146LaVk90gmIAOM
F+r9rLqJhihlATzPZUC5vjnGXggiaNTs8qcyJ2D3YRy7m5eY1Zpxuoi+ja0fTxaKlEoSZAeSU6Zl
qq4VbQq8cX6mbiALfxC6VjkjKegojo4RlWJSk0VATJPCdA8st/O3W5l139rDTkLh+1fl5QTqGArw
0KaMXr0SsDiq0lO8pBH6kZarv8O7KcyBm0Q7Cwd059ujQ0x6XMMvdwccmGZUYl5orpXrWlW816x6
HhLIDHSjwXc964Z9tRoS8xp736OJ9rxFCvde21SmlgniAejT2h0zo6qifrx3o3aDCQZ/d9yyuOP0
A3VYQV5J5onz50U+M2wXv6tGC5z3VCOK7T7fUGakUvErlpME7q6XE9r2CIJrUSq5x8EZURt+DrOA
TfQwRTj5vU0zNPUtM/YS0t5Xd4FQq0wXkMg+PQbEYXmSgBm4J/I0q6u2VGqxepgwMJPk2l66KnM6
/7ZsYAWqqzl79XNs6LvgROATQWz2lco3wRLAQKq8zf2IUef5Ejdd45gbI7zMCYsvGl9eqxkPrs4f
5ozCv6q9T0PZlfBK9AGAeR26I2AGc8Sh66EYagrl1bz8uVmg2XW35bQ8Ti9cGLPoUBMrSiefjbSG
6zZSXfnn27dhweuudQMlRx91s4BTx9cHA4DCIE6JslMdkJuokb8Kq0WHjaJZmDPPr7GfCVt0gFTr
E4n9Xkf1DPZXctUojCVwMtXssLitYKGi+gV80nGiUU46lgCBXSK/WFULV2knA3rIwDlqGZIguXG3
pZjbZOIvYtmJXvKuhh3Vc+oYN0t8JVXT4xBRnRrotHhYdR+L6bzAWvaSB4nJ/YM/vP6GQziXm7ds
ZhbmrD2kXxHgYWuL6cRoJN37A848VB3gath2EUDa8Pj4ohbmaWcoe0bbQsVQ20hMPyYDB2UUBvgd
gX/rS1w2NPZ6RGMWl6MlN3fX+RNOvhwErH2ytpbE77L7951YAu9YsBSGxYEomfCDgDWW0t6ONT1p
cj0xsQE+y/4e5/HmCwqr9XhZjTU9O2UHajqehlNOHt4M8TnbuuWjMdwlQKgYOi92/xG+EbiuUf9/
KDuA+NB/eRd4FtYtFdRw2YnTMBqwXiLkys3Rm9K1RUgIb4H2uSSNwe9NRBn+wnetBKzmHr30bTQJ
6/aeFsLw2JnXC517VP2mrPXBlsmp+3yXiVOVkzcuSi+nNWh3ser5bPFEVCYDwcDZK0lXajFOUXBM
U4wR7crn4ilQymU2iNsHCaKGgPudC2QiXv84/Bpety8JZqCebXnZBXnoOroa15m27v+VT3Ih1Y8p
/gKOnvaBvYRmKMA2BLvYGDBzP/7/36Kl0P23ldxBOWgYPtCOOxoWLKH/BoL67kFmTxqORbcoSbk4
3mY6196JGP8xrZ1SN4LtCYH6iOhqZyQqXOZvikPni8LyNBUmFS0rLGzqccyyws3r++RLwm+lxaDe
6PD7vnzmhusDPoWdM45gjNnxuIb/e1Yxg3dIILzUm7FEl8Tx9ktgrRmChtmOkRdtpUZCeRQeHRu5
J7iTCEHEtIrSpcTmteRV+bRPoUrNEzYDXy4psdV1Xf7RmArmFTc0bvJNp5w3oGZpb/m/qHo7CNbL
uo/6Icq4LyXLoUHcThYzHu/qaaiK3tOV7NhOVhdeMtm4VMbc9JI2u6c6T1tVBh7VUwymJxsJMgLR
lXOEI7RmW8v+v3JVAqLE/4cxUIOlEKl/4LfTKibQWKO9ylNIH7+H9/M/lJkaDLMJBeuWjsMPZC6j
zblIbv1vdYz4XdpfoEuKPy8hBOzK4wxMWoVbpo41H9JpFZ978E+h4MvRgiz5kmi5ROWOzY0ABx1v
y7ul0gO4ds8eS87+5aJ1W4IxjMqaGC2MLL3e0cZBPmRjlQOrua5+fbWvI/tXQkZ+HmK4Y5H3ARBw
5EJEce3NTc6kNRhuBdvsPhhqn/xMQXLKSKqhTt/wYKSeUJbDB13C3Hvfu8HOwgFf3wW4zs64msf6
NN2qBgSS2FJgsRAmQryU/TXTsllPQArYEw5QKKRXGT31G6N+Oi21GOuOZbO9Vd8dLG/+QN2iVjBc
u2ulijuvw5N52oOxhCi42RoBjzRHmLS4S7FZ8B8nlwRv2nJXKlUEK2ID5S0x/feQqoIKe+x3b2PS
JtCJiTPLVVQHRp0Qrwlh4SjWZj7yK7nqQCogW7ObwndK5hlh6JqOorsJjsJbWBO75xEBP6FhtWDB
vK9QhXMWwNcs0jwF1YMPjKyoWzD/o/QOnits/Sp5xsPmbi05Ijf7yk9QET9bcjcmfecCBwO17WYB
FMQfwZtWjGA4Be9X4o7HFn6E1Jax281MNHMPC0hBD4M3KiGVVKPu8KfMfpEg5HcF3X7+naEjxtTV
ZMzhp2GJGuyahp1gphS4MBLNhstaUZkdGU08h8vceKUMNZHyJIXY1RI69a3MLWCIhkClDKjqnXvC
YeZiPdfNDL9iZ6CFz153UtlFD7/oxzo/l1Ev46Qwt2XBFj9E3SaD7wUiKBD1FP6SWVhjg6aGrPwy
exXvTd3OBGkDeplP+GYzy/czYzfHszaRDQaQFS9J3TnR/NKAIcYA4a5l9wxjcWSjbLuSPyczSA7A
4kofUedxT8kW8Plca6/hM6HUCkLhvlamlpsXxqIG2yiesko6UIdE2eymtlD8nmb8fpFBsV4Wgus6
s3PXfI7xiOWJM1dDczkGi81NNquTzG0dto6CWgEgrrB8GS6v5nXYq4zr/OgdAwdvxpZOCiQ4uxDf
Tfo3+wAzMhRpIHPNsb24JPTpXuCTqc8KscJEzmA04/EK/Orr3QWxp7mOaIqZ+C+qT3zJhY/NkUNI
WXVQ5nnkaZ3h4xLcRtbXz1NtlillbJvPsErLohEL1PgNnllUG+euuNGjsbuVGWXyL4egFE3YTuWn
rkYtgK/YFpfYLcAOH+BdB2cNjxQrdZum0Pz+QaPfulBQ02NbECB+YmBx7MaDkPtjNu/6A5z7yrFb
omd/a/RJvxN9ao68rqDSe5OMPY9LNU+h45BULKMVw8RveStnzjSWxgzNtXOENWUyrcJzntoEACPd
QfUSErsg08iO2zNYH8kw7OR6ZNAjhkLCmi4ojecqZ3eK7jIkgIWNB7JnBlGHiSpCZJ5JR6NWeeeG
nO6jCKg9UQCA9EHqEsoUER6SReeQuc+A1QSu6PANEJRsufS5UfndRdKu47ZLccXHVj7VrF38ukW+
UjgTV1BYPhrm9WP1djI00puN5JL4WyhjGPuxoLc7MB9e1n78sQHU0VMPF9yKI9Q2akLnoOgoqP4z
YKhfizyEkwFRy4cD77We+cvvn+LgywSZLIHJE/vRFF+kpzOnjtASm88p7KeZC+gSX6OKFHMbt2c+
KOJFhoP06w9/uXlcAdq02VX25/7qYbxIzqK82fb7pygO+LM0njd8Eay9CT4hrvHzGMkhKKRzqSK4
C8cPoGyb5XLB8l9caHhyIh3FGfJHyeqgjI5gV5J4rqxhSfh1+xR4gTMzbgNAQBmfAFpi0QyepdX/
aT+xza/t6YsVsa3efcAcTtR8Ee+fkOnYQapG1H/c/s7UNWLh3ZbispFSK3LBn0/UHH/Gy4jafP5i
dYFc8RkV8K7c6WWebhFYuQ8w2Y/aO1bakPiXu5HkUkZnOf1k6ripQuAtwhho2nLR3zqbOXx9eUWG
vsWnoM8Qxg7ZK88RpM+g53Bi/7o5h91UEP9sAkgEi1X0kccXAHnZolckGRl707OeNMDFTIEqpxLy
hWrU0W2U7a6iD2o5wKjsK/zYuqSk+dxjjO1k9kCrNT0nPkw+NdTtHIAynXp7jOlAn9wPsXcYeIbx
F8CBSajnv3YNMqEOOdgBakVSuGlvD50tamIOoUfXrM2k285/aKILfhk7ZJg7E7Qxs2tEDWC/q8aP
eT90IDZGQbL+wdj9FAdYIoXHrHHyD8ikEO8yv7rOdRZqNeHekDmyJXtFcfuxqgtf7LB2AFqQAFsO
NpPhUUxC691GdDmhJbVrLwPRxFoPQ89/n1rXuULvBbzj5QzThvy/o98ccHJHbHJyaZTi0dvY0CPs
wqfmmp2BsRWirWVtMnnwLeriPu0utPLl3KntNwFZpwFG3zbuIXVhIbjma/G9spXi365PQkdO0tel
lWI22viP3mj8b+oN94toxSgzSPCtGSkpoKmIP4Nsdv6D9AbkTHLsH754yQ1ih3nGJY/29yJ4G8Ue
2ADZ8afcC5Ejtbwa9AoVTV/c5eMs5q3jp/zm687ysuGq9VF7VhpbUbewNubkYa9K8trsn/QuJHDH
vcXlNEpcTYrmLy4McAPN6W0N0DdH3KY7Gf/51LKvGmO+GLbZqvqFKQmish3p/j/TbxhgIPZtIZSh
3i+ZmY2yoWb9lak8JVRv4bRHFxurem8Ek88vBJaB4jgjsI/z2egL8eZLv4WlSzd/NBiF91o+LMGv
287gRn4iANmrnKgGDg86AArdA6NNGyEXw6AT/aOPNYiySkZ6HEC3eUZOnzQ9r7mwkDvN5MokWIXy
8X9KRErAyUc8UnDXF9NgXe0Zb4KZmrhshZzETt+sZvGZnNWYBVbX3LJt52mfybYaF9DzTBHK4Rbs
nVng/LpmYnTWQmqUOfOom+mRiAnOW5H2OIjCJLvIKlE/PvvIkiGaOShUqhRuUS+LQiho4LOgkVsz
RkUbvPY0BgF4HCz4yV4nITTU1sfxE23YuCEaCXDWcvTYf7aFz09KcUMfYdXpPZVFA3xO6KYwFDJm
KpwoCn6BkY35SQEgL2Ur46yjWKGVWgGMS9nkW4sS9tpVPNCfBgMlK5L2YIWbb5RgBA1s0XxUNRPu
Ra/2Z89BCJpCoHZluw6MjJpTM4hZLqPqoAFOCdMR52pQiJrANJraCcJ5Izfaf2WIcztnFlWXwlCr
4RPe2juJjfLs3sG+eyoD4Q6C1/GM/aYyMUaUxy4wGPIEM994BxY6ZUyfchM2cgiuC+vCZ32Hb9Fq
nopi/x84kskI5XL2+cKeZSSeH+MS9qJZX/OS2pi1ztcFtQqvn3T9irbvsfXhkt7wKCuFGMdSkG+a
gKZ8d1NCCuDxxOnaRmHy4sgXDzij8hkNVc83ix6l5RVJTPNR0NMtk3rYksUW/4x9W9wVAV4MEdnH
qO396ibkj6E/8SPBabq75xpCbl6K65KtK8UiQUS/dJZ0mr5UcxtcYbL/0Cve8PMKncLJiCahFRnm
9DNiZ7zWnEQRatbtGNQf8co9BJqx7U/CGSb3ov8C/nIpjQ6QrTMRuow8/twOgDAbbdi/rMpxY/NR
4Duy9y546nfsPjjDvz/60hMskrdvlekYhrpUlvzCbDU1ow9nBWg1RNhhSIzzrCmHFfnEqv87xX17
Vdadv3UzSfASiNsO/v5kWRo7Zy7kQD2S8i8rVF0tqYQIbxH6AlH0UUSkFfkOLGEtRHSPDJdkI78i
PLo8j+ltGFpCXyZeUJ69yMDP/iI99yA8xNP1YaroEbLS8awqek/eoaPgDRKcdMP3fgZ+SKfalRQA
mxiARYr87tpubxuwRh3vEc3jRM45IKGuhV1fBE+5Lnrz0fbmSRqFVLQJNhw5ziy7WqWq5126I/iT
sHxCtrADtIwB4cH9FlA05bw3+UxzhbTS+lgDb0NPummVDkICOwFP+DGH6vhUevcUk4AUbIA2I7Ag
v9gIxblaZz6KGkmCn4nUtsCIFSsBGUfjHzhqSCz6vlDroo9A5neDzQKVjtkCe68SnfVUc5wu4Kx3
6LGg3vGyBdzJY0rSd1ftLGvl6amHM6s14opu0/tRvySrCowDMScCoRIYdcqFYWbmRl+bRBi/Ev5w
UAJ7lECodzQ0my0uVkjpJE1Y+Tp93kpShp06c+YMlG9Ypzf16o9zbz00Nc5Hys+a+Y50TXgugDft
+DnBg6x6P3ibbF47GAbZcpZIAnX+iBt2wY3VMSAgz93ew7NfiXK7zpLCBJA0zClJNSiUjUuwTv4Y
IFu0ZJp/7vGehmb8E0xJXafsP08RMnT+jwuwyLUFzvnRLjLXfjckfumfV58baQlrsYZQsbi4hc6d
tp/GMz1bV3RTkz+wDHyNBtkNXQ0oLPqGY+XO/ZiLZ4/wpIJ8+uHRlyEoHH5levDmSDE+Hdl3m9Dd
lgjoRAXoz9ej39XyMDuYF/+ovyCxMaePw958OrJbpESOLCYKojtHTKeOy4xchqNj9A8DCW/DJCpZ
vkYth80A+uJxruST8mINBMyJrY+PqbtKuCkzdasa60v7mRgYSd46M7L7mViUPtJcPCF/HpjbeUeq
kSSNGNl7AJOPwFudNvyiGzAxb1jwC4fOLBTzk9QabTVR43uaBiRqFIJOE2ogmZmw9DHnWp5Juq5X
nTyklc0zL8V+LSh1cXZYU3yOO7vVoX2QQCZ/QnBxF/2Ex7YUOPjq3T7A8Lnb1unV+P0E/SknfCLL
iTSsMQBMs9REfdreRUuUOs6SxKnR9ANMyGLOoyxXNFL1NTJiQAuJ1eiOUKl4NNU7dk9Lg6VdfDpr
q9Qeqr3ML2+tDOD1xYjziWzk7R+ODlxYpAm1QT3tg9Zc3Neh9HCvAzJx6p/trdZV08g+IsVF5VEG
QSJWFFpa3ztJoXKA0zrbxC6lJAiw3hAU1wLxT8/VtRSd15f6Xh1fW1tOg84RYCbjYIiZj+akYZXK
BNPG7zEdbB1kJLBdCN5uZu/cOrPijPRr7sW21UfrKCu4v9zWIZPtpykcSw9SSQMylDzN6M54Fba2
hfzMUuk6TzvaPotqEqsG/y5cwQg3xaP4WLBF9CLehzUEziQhp/DzdQm6dEG4FItkKIqNFdg6Hk1i
/kE0F3siJ38TcjnuBzHAe7g7VGMac4bl1vJF+0WaY824ErdTzj6lD7WXccE9n5uXRn/0irNGFO6k
KXVDbjYir1yxvOb54VAFjRRZsb7UipqN8LpKHiYe7kymtYJT0YFnMyJ6FCOwo+1I8wIFuIT4t6qn
bXp1G5OI3WnxRVehNf92VqFYgioixMvuJyVW9ZltyDyW6dy5A1oPNr/2Qz6S9V1J8MI7gMxbyQP6
QSfdGX08o9sWnY/DxM/a4ohf/3yS8pkf5vT3oH82AczvmZ5QloFjRCXVq/YI9XgiDFY/3vnbbJXK
5+ngTty7qhdIf5a6WoW2ZkcKJ4qa5b5IACPp4tLrPyiueq8JMY44t7FhqtDBxVEb9W1yu4SO9G+V
uiRSieMVK3I9JWsTF1NUjvHHXWAi1KfZK5Jg2qPu/aGUqi4spmD12xSwbw0HmSqx1rwDWTziaYzx
vrUe9AQ30h5fduDhiGj+/MA5ygDlL75LTk6O/rpPbWxoeRVztQMoeuV2NkHk3s24AK5tmZWUnYM3
CF3k2Z9VBfa0midU+jKZ31Dehp1jNUMQm4qMWbSUnr93zUm5dqCta2KlQG9zAxqWfk3kGDb4SnAR
zROtJiqHCSvE5xcjhqAVlPgbVtD+YZ10r+0z1YkLfHadOgTq/9Ve+j4Spc52FNPj9Ir0YApcSdmE
58ESD2gWu3ok9bC0TPciFGIhG3k2M/lDxAaMK2K5zvhbJvf0UxAJ//NhgJ6L2o8Qfx42VWWQS8bZ
lyIG2ukx8PQZ7CzgdtqOTirJZsjDXM10YSM/oc1uKnGQM4R7ukG2LYFGgQTypn7ST0kBvLGdsd2O
2A5GP1Ek/w617HdeCaKFMqd6kassVdavMF2vWzDcR5oIm+B6kmU3cV7iEiX7qqzdUY1kFEwbfYgz
eYH0xiIH0q7LkIEpJKobCGB94t2jLJHLKJMDfvAZUoX64dvAmXPiPjCEvea5LsXbdy9Ku4m/d/EW
dCClPk2j23NadAN2gvkwWLtX8NkyBzb2h7oa/QJAWPj+1pgCQdhZGMpKPNF3xBMOWushiglKcxmo
wPMMxM86kriUYRxsrO/XQ4oe/pE065kI/aYkElW2e4R1VxxoCnhLCx6F1+oi/BuyimE/MsKj5UmK
TJCs4L16T7AXnmxs5ESyhUz6nJUNtUMyJEgdW6RMqcQn6VlV8lvtmdxW/wJ8/p4pi0z0ELXgvXZZ
eUTMld3VdcrnA4QJ2y0pQMW/GxJfp3eAdNcieYGXhHk9LX6g5eVRZOosn/W4Sb052djerRoCBNJd
fqDtzJq48AX/ExLI3aQeFuSIKX+bPDMvFSytPqJxsmOxvXAssgcuuhkiCvWP7jIe8kghF8bM4yrx
Ej4WLwb095EmtS3cpyAd5QpRYDgs+jxmoC3VJ4pIZCiFa7zFCZpAFzMbl7KZLLxivDXzexVe8JXz
9F0ss7J+XbAsRmahQUtDZHhx2n+V5xDEw+PGZHCuLSRYUtJb7wcYi36T5139lwSHYsA9Tq6/59f9
Avk5KKtxvwkhdwYL6VR2baFJKm0CFt5h0yftjyOKu1vGlw1WMw537+X/Y7EBL8yU/k8F/+Wb3UKT
lohOatg4xDLDSVjrae+tjASBw6rvabzj5FkpQ8PRonDqN3p2fmHttL/SPNg4qEUHJTnC4gVhI0QY
w5//UHlQglclYUES2kcrSHBn+OneNZjxr+RBkyp62162/fur/s4fUUGH6NhTwkF7L69/SBXHeIso
fMRsSvuXuaj9UFvPTb9YCdDKLMFG+FLzwf429h29OSNf1w3f7pquF0Ugvmjho78jvKu9svjtVrI7
eNJU0tBxp7srzYwwnR76g4MqoQU+NUeDvJkh8tgQfx2pA18gaSSQzo3qQ3Hu0a83SQiE1bUJsMYY
tlKwzWTR4XR91ntrY8ujViVcRduE8g2XpMcMQ8fKjThmcRt7ZW6eyYUxnN40mcBAqZYKtvgVq2f9
6ZmdQZAzAapMP+TNJmOOTnzwtBvJ0mUTfQIMIZXgYxtO6SuCHPz1J0H1x9GHNArK5VlBagMXIALT
tZ7t/jU/bXRTBCFRJL57M6kCpI04bIzkEO3tNsweJkqLNjnGY7sgS/PPWDcs3PC8BK82PohJgdP/
6GsM728q0+/E5LrVnRsEAR8otYA5afnIhZZkgsiAdl9ZfF1Nu3on/5w+R9Horumml0tgyOSIsyrY
aabzYQu1SAeUDkPxIAbdS4CJjitoq3VLUAxfCLGK8YNL9ZmiD8Ny7qITBLizNenqAos3g+a+P2fb
u9Ej7HzBCKd8Pf+yG636UEHVkVKSl4hrpqlyiRNP7ZhqHKsiks9HlSt9BQ9ihU6ydiKwpCFaWo3B
5mBa0Qem/VUenSfaWTz7LUnv352MAm0gzOJuotgoSDsnap+Y+E01IpVaT6Up1lMvQdbvdqfUqn7r
vw/6b5AcDRTrPrM2HHamtDnGHV/yOAMPUy6awmgq8q0EwnD9nNFEyYXoSB0nns1gK/LfnnRykW05
YtcEq2xB+o33Yacyi3k+BQVQ1f6cKburQkRPS/JcXx29jJpkA6Le/6XRyaykrodvCyjry+i0FLfX
2kMBsrCPUFOKX7j6D61D3nduLVnSyJTjnUZ5GIea/RtDAHRSdgz340lPosLNRf0aG5UAX9XPzhk3
jPQwhL07zssaNf2a2zTfglag0m+ZyHBR+ZRnfE3R8Zf12FT4X8K+QjBt3ciZrufzoVv+d+jk9r2c
QxToLt9pfwmY4EelofIcmSwOcoIXoEbFA7iWZCQmEh0TpgI95/qbv0jks/8KDsl9anI/HH+gXYUT
tNRIHmHm3p++JkKOm38eH2tRgLzXbdgIxbObHUq0kBX4sIeO53d5ZwCN4ZUoyOFapb1bDOU7OFR+
r35bom8n9Si4Hm+4MqJm4XtIz/YJfGgiuA0WoVje+F3kGqcqW+7EKiAvbVYJR3AdfstqxD/c7DBz
eHLQl3vrF75s/KXaCyMt1pVrtemG9Vj+ombXoo0uhuvvII57Sf8s1k4sN6+CLo2lM9/2/jR+KZ8x
kR1K4anIVbaa4b/bEtPc4rHA8r++ryJsuuwG09w6vxXxe6cV+LO4JfvFcJE2aQI7VNPiBwkDJ0kL
nINshdbzxM5alRyrmI3u25IOXyJnRLdsIJfAcUA0+hZDC7O+t4wQWNvF5n2gISEWY52gXRwoP4Md
RhWFsXlABoMRw8pdLe4ljBvP31Nu66FADL+cc7oElvNBVYU6uExxA3cZC2ujHCPFy0wkKjyHur+g
HN2f8HobZUH3/f3rwz9f0dd4Emvc7vF+Q6WlI9M7lKA7s2FY8i+FHJqdbVtxUVRHxvB3jXYlqE0B
eM5aM0AmffWJavIYmIFFUnW9YprUxrFxmd/lCT5TXplVZUbjhTWruvUGOcitApwg7skfZZM1DNcm
kHshc1sxhZCRmtyDki8P7JUcjuoPc6RjH9wkTgtZBVbD22khakeB7tM/ThPdZThxtVxLNNIc+IP/
KOGsw6Vk9WXv4gQjjLR5SycvEDCQFr8R1IwAa1W72qB3oOaXT0xQiNY9GFJFeBHtulWpjiq0Wu7h
iL4DXn4SxDTTOYr8Rn/wKeaclvwtJEp5RikOLyBpwkI0exuQDtNhPeuxE2Oz9JEQv6TemHAEdhT/
mEtTyus+GBtwBkZTE9/Z5Z4N99SU/zAlyRXpDaEErC6ewGqnVlXhbi8syjtbpYkBdJ8dQA5Rh9g1
sGOPGigtj1hj6OSrcIuxnzAOXUGWX5UOQBLnOzqLQWGAwfqCNm7Ms14X95zjoHWCkcLVh6+6XpoO
YWmX6bUXwNfEnt2QUxnp2Zw/DvdXgK7ogx2D62v71hymbzcGalsiEfwN8ppS/zaMeZxZsqwPgjNe
r55YRJxm0PAmr0Opm6QwNTkkCVhWHc/mumYqMRTmo6DpxUVTcvvH2V09hjwQMHQ3AWT9JNv2qUlh
d+CGEhk1rap43ePQFPZy1UrnbcgOUFnoojFut3nbB8nFn3V471jUevJSTO2dwys9MQpmNCxr6UvQ
sdrtxw/bc0EJe+nOJNQ2Nh69Tmq5wgNn5/LV4Q/uyb+RRF+TLQ4tJWrhWcPMKfx1iYB7+8cRbjDR
DUQ7MTI6Qepj392smq8cR4JkbLMGhClqDB+VizYJliIxEvDu89DmjmGJ12w5xz04RG47X/iDkCJf
H2XZwC4oeg8wiHqFjFIiUnzyMcmDnIRhHlyxGaCOT0hAtNmjVKxNPjf+WHJ/a4jMkgc6sztNWIqn
HNWYjuXsxEK+8FKksGNd+K9Y047rEGk+8AbdLHGmvgAInr6e2Cg8bHNdbBjXSg71rXKCUn+ikEjl
9Ll9XGwLRIhudnFq8rtbPoG6hTSNHdyNCC2REE4fywpgvLsObKCyGHVLvm0jAYWmwu9NtuAocvBf
xAKoMxLWEXB6EodojcxuuyQFJPAcfhNFfMCsXURKvgXAqJQlCjS1/AaNptUxz0nAFgcp+Zcjc2dG
goKnGNsIXp5izYucVONnlR4piQ8Dc3tEwG1aB+Vl7ySM/MgUyqCEzOMfMtrZpS35NmvUt7NOUA8x
5S2NmE/p9E5gSHF4vZdCXhcNa2FL8F+2/TO+Ltz2MGjpeGhA6iC9X0Bm6pn3yW452/ZP/UmyFvxq
AsHeC3KhG48DQ+L1C6nuEeCq1Kps7ndcfIOXK+QkhsWaEJsy634G+b8B/xeD5f/DczAlYcovjVeI
280GTucPDTDRsfliL1xoF75RUWkCNsok9bOfytrdYtxh7B9uRutVHfcx5qqPCZ40xLBs/RpCoNzy
P02DOn6ReGR/I6skG5KB6EKnoGCu5kv2ISRar+urdgj+8hcWfqMt/BaUvb/Kbk9FWcKmEx5eChD1
UhCGiDuo1J6TpRu0GkHlLWhnOG63BEBq8rBEsa2dmg+6T8TcdvOzhZSLcFzU0B6Jp8qsEzZQbvXP
MhvqvGIW4raXPj6xWLImNx5ssqi66MEDcStQ+JLx7JtKBF19Z40Mjkf650Gu+a+4WdGMA5NURKFd
5EmwEwpvnHsYAg0B/fvUCbMb1cJv99ENtUPikXIVebzu6SlQ8CFYZYPjH8PQjvNTu9wQG7/tzjtJ
4DoBXsafWfkzJLbHPDmMbj9Zwv/QfR/S3x4r+ds/1vK9yvBnNYzjojmqQ9tMxpxlnT9+QQk8mAY+
GiroTemPAC5Ia6np2E+KLfMsR2SpiqSRt9zjXCdPyESj0OKebbtFWP8hE73kygU08dMIKEcsySuF
6YyUtW8O++vamrvhY8jOgaIbkJCbVQvwSPTU+UPGpnrnY6zb6/z3Ll70yVyQGqV3lCgo7bkGjxZU
5UJ0SnLhzdNvQ/iJKmvSjL4JWpfxUaVz1sb8CUTakYe1CsCTDLV4ep6y3cED5NWlKsA+ZWKL+LiG
oTBGsAqo8J8y4cXWlM7gZ9Bri26RZlZg1j48kLl5uQIRH9sMICBHMAXF0S/gq71HMvLFTdbcD2jw
/1yhnW9K8bi8FgJRkJTxfj8jOPKnWF7J35L8yRCbhx4SvsZpOtMpHQyuqQjYLkc48cxyspp3TZQv
endA6/XAzbAIriaSI7yIdptLgQ65qoNCyT7GJFEfeYRvBY/DaIbILxVs4QJj2rjrjLR2aGT7p+Y3
/Q6tY8cXH4QjhfVyCs/96Nf7N8qe9q70VyT7mKJAen9sza2MNVjbuG3lbYqdzh3TczTRgchawDWJ
2CprCaTchmg+yQD0iJiICF1ex5E5cRZzPHDneJeEyFVpzKv4tIQmDkxw/ZhXV26aJ+jynkz/ZCxK
GmiJa5fLcl3KYM1VhV+lMM13XDGJoexGGb4lH41VHxlNfwWnWrFUCtWqys1gXimRjrVxWc25KtNk
IxO21gSmTjp1LGRnrpRaW+PU2dzGTGSbk4kyUHj6+eG8x9rkSTT/SXPdjX0FU7xf0vASpcV8pnF8
9y023D/6T/xsMpxtsUEmxBh+ZJu0smZK1SJ5/eIkj01KsiMaXmT82wkfhY6yTULNvcn5ln5QPnnC
tw1Ws1fEHQNXJAjdvUujCJUnyL6p+sPYqj5XegpW3JkXtX0/5YUmErtWI9M6QygG7aD7xoGb4CMt
Zu0NpoIyh3h7RauZGDnis0FqFTkocCJ/cQI8rtdcJsR/mLzCrOa9DSiJcu6XMxJBf6E64oard2jD
9OlKSFPXKx/msQ/6aIBiUJyrc38+Q8bah3fChmq/ijeeHLNPDyIWT1oUKIc6CMmx/qiWpTDmgJhV
osuionUSDI49391jn+nxN2H5o7iQmeWBAnK0qJ2uIEEf3cdirkIBGDuJNgMaEkzCV2owK5V4V7aD
jE/ZSTOT5TzA+z5ZMGiiWFM8ttMRFSA15BG9FJiHAJYGsufwAmk1HZUEtPoftIMo//IBKyVL+wDg
+C7sVRZw64/pEtCK3jCa9v/MtWTgaEHA+5Hrey62V0WJPLhmDwREtAReHUkuw7dKx/zaM1lUk04n
IXAljSQ45NYM7j3KYMCorYHMki/4cY3PlbRcstZEwbkJYkjtPqauh9B8LkzVDNo48c09c7etQid6
JhuOc8Iseft4q55OMlsXgo+DR/fHXJsFX03crzVLV+o+V6dBnXUl1ekYle0q7XWCSuLumB0ogn3q
kznxx/v49fEslXNX71Oh6owEOrqWxLDfLve+3eLv2/CWeD1U3+4FpYaHZtJ7s6tyvZ1/DoZtFmBT
GORFZw00/3ZBtmA9+GHqiSEn7b7en1FZELeZhrxakcMMEswouGdrpqW3zROR2Vlvd+a6yj/4owv3
rgcQUaPbnlM2C+12+LkOT2pllFopnF18oWQwq0rscPZWuZo3IZgP58XOMpofCLPwwY8WBiYdMb6Y
JLcTPszEjA0UEHRlBdg1O9zPdRhvLXIb6qQksG8mQxBgxbR9cO6I/a9XjOH2ZPucd4owe3ARv4Ju
SH7WWlvmzm+q/yBAGz+OCTYgQ9cPiFawp1IERVQ4RS+c8je32avL7hiiFvIPIl8fuAy12MPHp05y
X5kRfonm+tzf5Avy6lpfXMQ0MZ+2Ju7brEJOxMoWg3tl9UVHfyjbeNaN+ozhU7IZt3Tv+lo82dXd
nWAU2pKwPvnwAnQ07OM8EpMwWGSI/0LaX1CDmTWcytsvkCLorKOR3P5yqxYHUL1bliGQi/E0upNx
mwby0zdG+k9ATbDQTCICxwRLbgLbyNNzDFFMBavOUF+S70XA0qTxlz3Wj8V3q5NWEzo7WO4buG/q
Mt8hyLZc/exusun48JlPzPdATNAMmHc9sYCQOdZkO/a4fxmDj7xmzTjFAAbnMKSlYzJozrtesox5
bU/3cVUU1HzRCTFbC+cwWEVPiONc640KC8MReX1mgzVK5FQI2BzVYQWjBjUZmFAeYBAKaGu5MZYM
MkVrB0W+0q/NRU5xxqFWO3PgUmzFiFx07/5aXUJsgu1vbGtwtx8rqZ1AadttAkRxLmAzmewooR5T
0qXqMQM3koV50gYBUReyPv7dHgy24gW67BUTaXtHBEMXNjTxETt80G3vyFUGBHPRuFB3pXprKUKK
DQJanXA+kbpnY2faDsYhiPSi9uGazZTh0onohbfkpYlfEV627ZY3PCKUgj/nLYoUvFdUPab7vzeV
qlYOFRxNgVk1vio6GQQWtS57KLVwHrnukgoJdgA6ppNaStiFSmUUus0Q+R7ihIG666Owm6+67Dui
k8g3ME9dn5ElhVJfUlUwNaUXu7XTqFFiIFoAMaSRRWutLE6MdFexygDmmxg2OyQib61ckllFY4gS
nGB1EsDpZDhV3YT0Hud/M/4Gr4AjB6Tl1reHCG+QD3ppye2sIdAPkyfH7h8yVf6RW900owC0gvut
XOaYSB2PhdsxGtulzTXAWTSfMJ+62WIWL/LkGqlSia4NLnhBjKSIel7jWG/LZbNFEeiESdJBm60U
kOHc9S66Dm4N8j1xszG3w52pE+FJmLapUSzWYGii10Nwr6BbLwJSoIA6OzDqimX80Ph7qEBZ5gLY
hrxZwLA12qAqSFZQNwtlMBZJULrS1bgCks5DH+ntlwcq4JECI/QHj6QiGWAl3B1ctBOhEgsW1wVY
RA/4laGWGiWJ93RrlqWN8EOCHVVh3oc4cktdEZ2FO7W2YzUa+C5s5hIbhKGsD+08BLXm472Wy4Y1
hO8tjR3NGngkNtbsADc2cJIbxo7uYDUYrn/yBuzXfUkG3g0rAcpKEz9HvZiTe6Li+56NXLB2pJKB
b8C4RDjo3iccQtP5ei7vLdqhuRBgnAiPsUN8GvSef2SGTnNNbrMrnwsRBiWEuh72PM24VaxDo/AJ
MKgHO+wo1KxNw/qNy2XO7Kf+yruEcEQoOC+EyZ65BAnG4932N9eMdtCLRYiAl3Kd6qkIFEhcceK3
FxwXDlabSFveytqMbD/wE0jZwsykMLM/UEpx6Yx7+pB1QtdKr1e2uodGM/G8utRTIrcN4C1Uk6Vm
ezqKwn99A9wdur3gvul8HZYwfO9e8sNK7FJMV642fEZJYPgiY7gTJcoE7DCuaQWERlPJ/XCLOgeC
Dy60UsH/Ki1jjoAclwTeOKeQpsuidhbdQY77DobdVZ2X15NQQ4gBR8Jir+OwwFyaMM5sM1adF9an
gSinD/ebzciVc5akPU6fZ7ph4Bu/CjSAZ7dPpO4+f9dw2n3DZ/Gb1WYDAlZD6qJ3XXNV64yexz5M
KzaCCWVc+4OrJ772weNXEhJR0ZrH3oebnAhUHTMgqtsgv8KHcstNaopXf7TGy9nTt+9Ortpzf65e
IEEETfyumyK5j8n+At7l7QAEV2hWphsZuKdl0Gnv005lTW2gKEBhTdjkQKFpAoZQd0TA99UeYMzc
2XX0ahDi64TtDJ25iAsrEW0Tlhwf4LZdm2i2MXz640Yj4jS+Tp8QcmDcc99J7YuGH+8OcOIdc9IO
0giNp21PWNp6i+eo87zXYD/k7hcLwJdS+OSZJZbKrzjTkntxMwAhm6GbVE63b3MCY28fcUMy2gyS
Fn3JcmogsGJHeomWpJedOsLQoHWuzBNwxu33YUbVkitp3U3C3/EYVgdEk4XLLDT5Dk7FtqBUIWoL
/kuxdF7Gjxrk6pjxh9oJ4wXCuGar042tEdOO1ZQcss05BbzOHzEVdcyQBEY4FfanDU8kYxrJ6Fdq
ZqQEkGBGVcYhCUFrt5lBJ2qdEXoYMqy2m5QP20LLbYxHYEox9RG9XS2iOgGWL+TPtk0OEFhNumx0
LCyq0zH/eh17O5BKFO8Zf8rtxrd3PsNZGAPlH7WAXD0jOfQXRAgYc1Aymi6DhnZgh+lwsUS2eXJW
2cnAhRB0PPacVFwx65NOOQ0fNYEVJGK0b8olJ3b9S8+8Vk5drIyWzVvEl0F5r9h/bDR7J4NZv8vo
2pp2vB6Ex2UdkfVLbIcvw9bcmpCZXlffg5sckwYw4OtueH3CWrpy4HAyebWdliI9eh1YGjQcES6V
6o2xXwT/qHs+Q7sJ6Q2TnBL5d/zm36qwXYqiXtbawyGiY/86K2S5nE/SbnNBpwuDbXde6pR57Zzh
hqMwkq3rOKKuY9p+WwLF0jb8hspdtEwIrUpJLxojOC0wtkyw4Jva02ITVHtc7I56DXpaAaAIWtYM
LIEW+LMOsz2qxGfjXeLzI+J+SQJKyGNZ4EsmSsJ1Dk4mLSJeAq/n51L+Eu8u53XVOTiC6s9BXqB7
et0wTqTF0afST9j/kNC/muCp79baSlvuNJeeXCOLR6UWFT1jlSF6p2XcDurmSkicks+Myw6Q/ysc
dLRfB5zMusqWcSdIQIjq1SOAaK8DaMXcYIMXcFPWqOqUb56E1MJgUAbTz3KrAHuQaY0EaHcgbPA8
jTe5evZ54MF/jb2W0fwnJmxxpbq5T/F+U7xrth6uBivfnDTAE8xwaZyIs5JO30Ig4DiyLrEhWmak
PoMNE43nuf1QRgc4LlDJ+hSCqNDJjtH69IDHOvx3mYyhnTmC1QAzKVijoQOQcbQ0hUxSrjXDxht/
y7yROZzOyD3s2+Mi3fg6ptgGTrOsBhhrO4YlhesNi/eHLDyEDYM8qIuejOMCWpDFfzGc1fKBYS8s
3RvMPNsvb2BVED789lpZ5Er/sn7q51GeTAYoFc6NjAhh0VUA0lR+e826B7V1Oh4Azm1BFaDbtpIL
QieV8IRxMJ6yYPK9yIk6mjVY2Ta+rpjrRedGJR9JJ3aEJNKBt6D7kE/BI12gtA/U/lcP0XDVDNMQ
hwrs+JVKMZ0abi4b3AMw83tt0lflPHeOVeztaUS10tcKBjL1ezvDkNo4FSzk/dpfjPE9gao0uiDK
4b+YTO4HAUoejKrbS9MNXgtvH5u+YCBFKTC7DLG0i/1ZVnwRFLDCkTufIGFE4IbrxT+yFC1ZqVNl
56Mv8epfGGbQyULg9q3OaLJChKiEMIc5AXVObCzLRUIGQZdx2DumTnOlP3v3cdLbnFTp9IACVAz+
fFarbZie7TqrytdXK8YA1IU0UdyFVw1WiPoYeyk43NtXu8DD8JTPSLTOoVfKDg8EwQgXBxPoMHTI
fEb+b7VdA7CYt42wRNeeyFbqqkTRi4qN5UEXO+T837RLiaaqA9JwbTB+CzMrWktq81eMuWqIUxF6
nof2Ip4otk0Aafmg5emoJ+vGpsGYleyM/tNRUvaLzYFzJk9rnIY9lzzV6x+UzOtX4XAdKBUhfptj
Vo6M/ldIpyUa30lKi3CVzkPx+N5ZpEBmmnvqfPJutYWnxt2+gxVmtbVQIwbddt8oO+CUS/dqRrCi
mNfBvklNe8ai1VWYPL75+h1uFBNJT/PHGEDxoPZGiWduhHZcn/r63Mr+nLuDgtXOgay7ayF81D2u
YtxFzOD1ctF5+kz/ooZhSWzLhe5L/kkPdg+ALzzbTyCgj9eH/BM2wvI0gPChw1o5zOt6SUXAm3QO
C7kRDcFhdRJpem86qKjKVjbx/3jh53zmATzonDElgKgsFT1UlNWKYo8E0ZxFyjQRnkuXJtn6bI5N
GOpPer3BwYx6DQhcGuYbcvsfXsidI7WUe7bza3LhOcL9mHoy4YpN0SdZz4ELfpYllVhAtmbC2CZe
gcLdBkb7WobqcVqfNL7Xhrnc6i0LBwgukso0dhI1FzyoB1+xqmwXi6Zly6fNJXR7ZsBF3HA3kk/Q
+rGB9vQq/y1V87lorYqHV7y0DYbdxH14xrz18FgkOBV0EjP0qlnN91boJ5EKqzRbkyMqX+/BQ1hZ
iW/QM/37qJYoxZxS961AlKd/H2hOg8LaVZaBgMakI4zE0Yqe0F5+vmXTJtQRtiYm77kTbecpq9Xe
FJ5SxLU+YCUY5q/f5prVFmbHyLzV7VmNWIoekm0WLBUd5gXPvtacLWcOYWEMLeiKZBMBQ8n3jT90
DYuBU+yrki7Xi866f59zjV+LwisruTJmaVWnRjw7DUm9TVBK9qoluI6fhnPn7sAbypXvtkF2HvgN
N+dKvK27LGOm0xh7daoa/gmb5RaL3RvAh7T0BBt0OmxR1R59wzWB5c3QBg5U/HXVHrEoT8xVTCMa
zGcoQP9MqZZNSWDSKn4LH8AMt7rVaFz4aN1x12x04r47fSFXOSjaUm3iG/K4MCDu2IZfQ13jwhQD
KMtPN6//ResHZyn5213ZnoRDCJP3CJG6y0P4vuToCfANs1TylZHExIA3ctW0VNoN/KpEJz6mtugc
uphk/wf5nXvl/tMKH2Yy7CmTiYTyiXiCdcWt3hBbsnr4cWBZlDJ55YnShgQwfoI3B8TzEiQeoQXe
/yoeZNUdB2smzYe2QiG6jZ/12s+2Vd1Bc9t+p8qGYLVGJ3cIAgDligsO+Y9lnwCxOU0DYpDn+55e
4fh3iazCVG/ez2n2EXtVIC83/lf/nVgkXZ7oBoFIUR2i43tOCtl4F+8T67TVyuTXgArbmF0oB/kS
xGH6lz+V0IpEI+nFah7l2y4r2RuBJ0zW3W66VvnylYxhboj5F2rqrvIf6+MFD3DkOphKtUZIL63o
8ambJiRNUM8R5bWY6jwsaBUJ1K6sh4bLkhCJ/jBbkQ0JpENUA8ocve/YuuEJKILv8KZQ4WveITsk
uY9Yf+6liCB4ked8bb7MH1w5fKaULEHUbqyH9EcGTYi7Lj+IDpZ4ZZ8iGntR0Feu7AXrsp1pEhkn
nobcXba0GgeXDhnY7SoxthKePi2uPUSrKJiOYXzDAHeGeZD0wSR83p7+I9XUw6gqmpEjn7CP1vIV
3q4+NYaIKC6UbW1TNSArRwC/huHElDzSemparUc9PbRvAFfaEcYKMf63oWgfeX+DmZDifQlGxzBy
480o7KxHvZkJRw0xVeCZsUcF3SR+72aJRqh/cMCIqjxO34dKsRJJ9nk/2sopSfJ0hJjTsu3GGplv
Xi4SgQqxhPCk8SrtVF5so+ZcT3ryjK/VsfxkWRujGBwocwIBa2wSsDUE8SdMeIImf8s86CkLwLln
G5eh2m+xxdwQcXdJEwDNxXBZpIjpWKaBdB8eYSV7lq3Zqph+oHQ5+bsoCEVVtD5q6HSuorvNWdrP
zvlAlIV4rLIHJDHnvvORf8dqeQMhda5qo4XW+6Vir2h42rVMuBYLH46+sy5Jzw6FHQa+5bFwMBNI
EYCq1k/LN/hvP0VdP0vStkmgy09vhJOTZ05kzaE2VvFNtCpDVbcacJC1lHH0D80i38SdfyNxys2T
u9Jra2IZoTL8Qm0HxLa1NeBbryb9vlDouW8bevA0GnJ2IJ1h55LSsETlratnaxRHPaurMtZA180Z
0IPi5EDeT6ImDfaM0kmpbyC6W9mZiH7cSbjXEBbZW941wbq+umCXd3Lqq7ZMtVTbDXOpNy0yE26b
KbUnp8YDg/UKL9E9o3oexouhL8wbzD3KQeSKnCFNCdz7r8Q9Sdzyf9oBT6eoF/HHeK1p6aP8Cf9G
lXtJjgdW/ZG4gDZurvkAjUO0jxH6tT7rcIXTcbFPyMs2Ktv8GSI3i3CEgckKySY+WDWjy+C5bqfC
ZM6xX0M2Qx+Syr+YlBGsSiqljrkMtTuBlrC8UGBu89NHnpJPfZZDhqVScXBu5aZA1zdGEgwHjAUH
UQ8mgRIcDVMNmppL1PMMD9Qgfjwn94fqN7KuQj9dlm7EEcBYovPgly+0W0YsjeMDvj8FbRz66CMq
Nw9/i0kziBH6Qg3kzPCXZ4quSBTqTPiQmvJXQTccrCEjYGx7VFDgZ5bK9bQLd38L/5R6IT11fkx0
qA+f5ywdKIsduEU1IyCBUhMx4sT9wCZ6iDLvDnXa0wGWEf5CkBggli9peYXmE8BZ8hmWFjGE9SCu
RVCtw3lHluQ7RLDIplGp5fFEYMj1QDLDqfRwUu5BcLY1vIl3HvpgNRcvK5dpUQ7JYhZh5Y4U1c/M
2+uzLxO0mAGMAkIXUzlibaqyfOGl+Ij+g7k7wlbZOgAQWVSKRvHhwTp0kPN/GP8UMRnc/Vex8PTI
tMqAHpsNN6JzYde/MZ0uD3iXHsBZZMITKIsxklKzixZuijor+WOdtOOL+jM5lcOBsuClbw3ucI8h
NPFK1WN4b7vH9bhRv0AW7qzDuTxuoFdrQbnRna67Uk9Y4ggIvnydJiAmyJwnEQTCq5mBFzE6SZKw
TUK4rQXzb1+aE4k7l9/odALa6d60k6Q84jMVN+btbhSP0qrq42PbxvG7qaYUqaiSbYc53ukeWlES
lPyiQ7wfn5yfI4LgpL7/1QEgNoBqtr8PJgo1HAnmI4IwhSxKgSpM6wRaqCUt+5nMiGOa/qWzQMFD
BE2hVu7vD2q1ftlzzOqxas5OlFgExUfGv5q3EzshvvH1qWKWcb0MD70c0OpJecvb5+0TWVkxZ6vR
Vpf9KjOcqfoQpw6sg/pH181RwvBkO3C1usGMWhbusFQtxggPm5+Jqu5hdbOJzhjhFarGjEtky9D0
vvPi6vLJFc5UIGoljq29o8VFR7Fqmoo29PZRlLblxIDK95EJqaGfqeGDKsyhzH1GD5oO5P6lltU9
5LtMqEHC/TsXAtoEFGkhQQ0e+ZBZGi8GSAhvd/6GeCCTcLyCjSagGW/vKMuZC5Ldb5NEUE/fNFUu
hAzgjQ6hRY8Pg33GuNhaFIRGpNco3vcbfyy0jnZb8LBxwLhPQR4WD+o8FWee0me7ML254y2cSjrr
KSrcD/0mZwkYcLWrkuzHF9s3riM1cUj4gPYDWfT4uRbmYeN7jS0NOPdGVuZD4gRfndSivA+7LZwq
x7rt3u2wGLyurMPceyhRCSaNzWf/SeF2fPNk/XEpZozsyrLQmfMDMmMkq53zMJN3khQcJHvHkENl
rbdBKVxi7paOX5b6Dom7bTv3a/8oZKYp/d+6ygdiHjFvC8qTBHo3h0LhwFVZBW5KhDaU/P+XLSwe
FowE384nzhRwMcsSohTd7VU9Lfr8kNMLl9Utr1qTGpF8BbPGVk/f8vBwgWSVWI6Iyb5LP/G0IV1L
RyyKzYbLpn/3xZHcd47peVpHLmYazaCPYxl+EDmSVdCzwDQQe+DBqwxGvbX4FLPr9VeMy6HFzbXE
/vk48eaIPbIr+1P8hkD6TXH6q6uYmr9a280aTF4hYUI38qFm4pBnACDpjLTaj4YbRDDAM2WM0uQy
XSipuUB2UKOJaPl6q3NDuHtdfL6itkhPAbeOQtay+MMtvq1rL5LkwKFHrqh2cyhDAKP+kmIkXN8U
gaEglg/jyemthVezmq1NvhZAxvBgsN9N+dXnDFmOgeXgawC9OcR96ie5HHjTsqPstRpdo5umvqVY
Ez+Y7sWgrXlqhslifDTM1Om5IGlzKbM06aTA463BfFjDaWjDpXZdi8qvhhTCv//YSP7U8xS5zIfd
HKLl2whUf2m5O1V/ZJGHkhW4J8HS5bA1sWhy7jcpN2OE9r/hXK0fOD4RbUgLlZrTa0gk7BzIvkCe
S+yTcEiAwdpYjpgEFLq3n/Ram/k4bYySgp1kfGnnQm69JkpP/pI98uxkJPbewPiian8siK2rlcMA
vx8442C34/MrkaANK6x54qPnwiOBZrAt25Yce5ITzBo6RICL+2rzVG9Yt5CBTDbfP56AM/zqtjYk
XSWH4Rba3rfvj0Op31Qcya7YERdJ2YcWf+GCoySRL5uvDZp+zQIJ3g09Q49c67IJa44B/B+QkFN+
bctTn8uLFIFVgY6AmEnNVBNq0B7jNf1Z8dsGz5CX8u9uG1LG2Tuaun0yH29zigAyehFZV7K3MNpF
ghUW7OKRsmaii2jc17uxc3hUWv7wzbS1YnXPeFr9BSMVnoWXb/LLuau94DGBHHlZOYwDLxlpiiX5
yXWnleVxqcjlJnUE6TOLTI/AOOzj+6+YvWfHYUZDASxbn8RaUyVsu0L82aifcJ5VSW8O6rO5U1Gq
okhUPQ84OSmNn5/PoU5R2YES4LesEhI2H/LsyXiCk8UPgVQC+Ti0niEy0ktA25z8HqIoDzeyEGXW
mrg5vMRdHbcwVskXKEVhx7KBbQqz4eh45CiQUL8vovduPPaLe2FV/WOGvwp50UCf9iFlFQuxKPVN
KFD7ujTuNq/JXITUx7EdWXbO18+1md4i/Q+VVnRQhZnBW5CAmiA3Y0/PZKe+FxC2hfOyF3jFSMEX
sHDAMMtIcDIP/Ssm4UEYkfHh/2uVtuSXXFrTN+Txj+G17gWXjdyDLrp58LyrpvyQY40yEqbFFNIB
N/vLUUVV0DtYsdMRwBtONMR1LXU4zLTdLwCzoVs6iInX/jUnWs1KHtW51g4OKSvfufR4RTsSUomd
6S+vjGzCh7BEgNDij97Dmxh7UOPmwzwVN0u7Hrvk4pobd85sEuAreVWG4wY3ofTsyJLu+dJIe23N
mo6PfADwYFVDjruw9fJ8DXxxbv8/Yyd6AvxbeupQnKzp/3tHOT78HUWRd3k7SiT2U/cx5qyYTKXU
sxj140TuJ26jmG5gep76tasy0/lngnK5toovDuFKK0S4gfe0VL32cmsU29fRtBMsTgnWT7fEH7WN
0LWjG+kcCOh4GXQBORGkWCGAKGJt0kLNDg9Kj1ZCXQVP9qpM0k9BHplTL1L52NVJIYscJKQoNMCF
Wry9QrjSMKq076VKsCK23TbL6Xoc6xKh765vqDPrI88hpkvhrteg83YDyXr0UUBBv1xPybSA4tEw
Du270f6YVRzPtokuloSFJZ3IAl6FC6apJnJOooEojqSElXgu+KdEqGGCse04596/jT/KlUrFqUU0
KLZ8XmyiPnUTX+OtJECEU0eabCxEWd9CYakM0mDhM9p473vnY+6p3eP/oj+QXdpkhV5srA09BA/I
l65PAVQTC19XNN9ndLGjwOWZtapV8SmY5qYDbhSdJ4hzMImDDRnf7eYkhZI9N/DMDa0AnmSWFp9o
EgB08j/1fWf/sl9A6YmFc4Ur0NyTTjgz+vdR9QtEGabM8EyoWmyJXlGnU8f6AKeQVzwtcKxLE4or
mUMVwwcJxkrwz7DZ2VidgWQxza6ZwvGsa7PjxQHZ+wqdnibhmbRwkq3qIEiISHmumPx/N8v7cPZY
rR6AS5P1zRhK0dZ6OsneiLou+z2OA4QauBXLL6xLFJNKhgRXiSkuEu7rCiC0ALq4awgbUZ1aC89D
3gseaA+V6sdNtB6bbjuDl2uNw3YnKcrhINu39XBS4HDEJRw3eZsiMwKfeivijgbJl1+0PnMvRY/U
rNjJ/mUtfNfRio1Ss6oGzyWfMcGnDpmnjGMiOuYg6e7D7YIbUJPgT2GEzUXG5OaVy+TO4cQYzOqN
N+zLAyTt9FnJQX+VwuuB6Y5isL7JIGCsN1j3yMX1iH5CYGONR2M6TWcT+G+iA71bE+uUQgWyMKc2
TwQHASd0SEc0d4YX/2YfC/HXAfUgkXCbPV+R6IXqDjCQUdnnOy0y5p0QAu42tjFXkWBRAAuxw4vz
GQSFRAIetDksKDxoBBAZN0kOqkJ6Wij7tgOJQFIRNSpuRYqsj7vfB4Cm2UE+mGhBKiezUAm1t3oj
5S4a0zuwBUminfwU9K3Y8eLgpebU1BNOO5jdxXeqaDPn5V+sqht+LXTxInNF0KAHoOu/eSNcrGxk
z+Mwp7JAl5598TIqp4WR/SipNghhk/3m7B2AOU2oEcjFHz8EOmXcqwC+2RgJoeG+sH8rV2EE4UD8
1O9k5LweQ0wOdzu63vrEOP9mm/eXG3RTkmUfb5pgGj6sb+3VeU3INb7fclZmPcrKf5spT17pJ4Ts
SecOw+Yx1w+CgFxohfGzPYPC7NZBaLzdFqAr0B67kgGVofNbr3lgRu+CfVHxelCZjh5oXdCTInLD
iGMVuQ0q1/hmHU/VMKkSwipYDsAeRgKtnXpwV1J86t/1XHK57y4H6CS9qqXTWABCGD5uxcmakWHC
Fho6Jjj6Ac5ckQrBvnsnqxjjoWjeUCrvM5qU1T2SLsYUn+znj0bw5rDBGjPA+03ICpTL+/6PCie7
KmJeqAvaM3ML8Mqn/NCprHB3XbJi8SlaIzabHEqt1ym81ENwMIU4hWqpLCawuaa18NyxEGO9KbIz
+Z+fGqajQPRWlqJCmL5h9d4IbAQwyFWerutNMWbVsS3CjQoidGtNPIzDgSpi67WkFHva4tcdzWRI
eAiXIGrSlUXB+JfR13FIw+stCwX5WtcF/z6JWP0TKphBSQqaMJRSLdlCemAoBiBw1D7aH9YdwHJh
GjIO7ttTqJV8jNdPOOrKriSkqOWkJkUmfle+PtrmJyJNQY6ZXEhgmvdXMU4L5UgcbLMmROG1GBBb
XYvIEpGqq9yZ9o3qIKdZUWjyqGQFWUOqYjc1jk7tXscAGapX1mVlhgfC2I9AyQytAsKgegLoNa5n
Zt+mGS415UmTYl17Tks2dMvP9wuP1Y7+le1pWDyqLX7dLDHGSkvQrHQFVxOiVZrq+A02XQYtPey/
yBSZvRiH4PUsytLK0KRZYRQOtAt9oV/TfV2+C6MWoQjcqN+1kOI2ulhrLg1RSyb2qtUgKF5tQaoT
LNC9/0NLyhFvkbPjboBX4S9uYz8e0rI8CUD/k28OXoAmE8S8wDLZPjZ2Dj/hxQ7Xtqezc3LsggeB
Ozchpu8zgjZFFNM93r7LUW9O4BMqDCZCBST9fo15ugOJnrszoG9Xu+UIdxvujgMol9Hyk5ucfhnr
7XhjRQ1L/+wmkQddgZEdgunQ9zxCAFhoRQxw82jc+uuwrP8ft4bQM+mN7i5SKAMfzmdo0wm8UPm+
HNkPqlF2Nn7n38Q2N9u07pro+LW4D/G6gNBIQbY8+5SK8uNFKY1/KjUCvSpHxvZUPmnskPebiVb2
19NqBibxr7Dbiu0tc+Z4rCdL2foMyjb9mut/8N1nyFgS0lEZNm7fPgaotr4bcqciiZQXR1PIsAAu
4oWSyiOVVgf/VDIyWhPn/KLHhWerc1++y3GCADFEFmikA0nWnrqn/8Al7R2DFdjVIF4IjdVDbXI6
7pBKcs66IsHIv56klL9Mp/d4HdhOw+VRsx3jSjmoq3RsGb5764Hd5nIf3vftmSdOZzK9ODPYZsUO
xDyrbg1y2VpC1DbfX+VZzQIp0y/nin1+PPAzuCG5k8V84a8lhhBmkeyFIR1vCWThC4XzEuZGTO6L
x3xpXwTNv84gK8oJevdQpi1WEMbmoWHgJXIIXhQYBrWKnhLyu3x4omDqB7ZHf6eLPkSMAohQaxGE
8KhvQAfLWOKrT9/zu3nLJXIDd+RAknLyekTvFU+Tn43fgUwRXnsIt47LyzGR9p2aI5Lg9kApGHtO
RX27SmMK0oUJeCzYeFfaWdC/TGDaNGxPyHfTbskB00Zxaajxi7HsbPjC1R8dzdtApjfZ2l4nYFVi
SqRej6p+Xss69nE8ayynZ5TjQDdL0+8HoVOM6awk4OiEkPUR6Jr5rSolnordRQUo/FTwHaq5/a7U
iZUGFlB4ej7WBWjEklWswQ32Imo0Bjt5DIh6+nRnHHFtv+XkTbmaKgtCwSU0F9SIt+KPnrbCS3Yc
TZGhZNUa5ulSsEJHU/Z5+suhRv1pposj14CwoAbwBEjlMP76SBUlZJjXVPf7+QUKaETUvD4Tz51l
p87aNI/3Oa7TU21pf98o38nFHkvFeiWcVGod1Y8Moa6yIRqEhufx0r4/Ppjl3ncEfn9ixO79NdKV
FKIq5Oq1lx/nYSLaJo0Hbg4myUgtZ8/q2RLlikvwskvR2P8PpnFmLPHGhAjCOKS/YEpHSYRz2TCZ
9Q7KZLzmuSZGc3sXjm0w/kgwgPYSs9sDjN/rfs0OUoVgw/LtBLHftgXLHb3+AzylNQOQJIBsmF/q
DpI1SVne9SUczdDNyuyXPNfM89LIaIcAB+/41NMYlU+Do+3rsXIxLHq3liMJVlW+rsrhvoDmj30k
UU/AX2u78NZlMNlCYw8IuPqICWs+q9dLydcp0Gc7LIP2bA2F5QRnP3GVCgzmUbF6mtyDsjmwcRhM
7BiFGfT18EVEBwM0G9quv3q5PS1ofp8qRpmDyOydYqOOB9ZXKGCpzzmtCYLX3oM0/xXBHV8qxID1
eSXumP/kK6Djl1ScY41ITPiez2kERsTtT4Y0JkNjPdSPuJSIbHyzFlV08ZQ7p5+apz+fxjzGYCaT
NYn7YXK0OxI2yMNI3BVXYlUE6ESRvIudF4s2D/73dT1b+8MjikEvsI9HdfJpYKfVMLP6doHOwXXI
2ZnixwlRHNjDeVsIZSjEvkuDfHRN1DvItGm+mGRkxHr0bvID+m2Sc8P0XpECCZXngbojvPDjmjxk
AqVi4eetVUifzZA2LWirA/GG4QE9My0RBswWyzhdT7UXWDLn/z7Ly68mROfPUdBBEiGThwfrBU4K
n3qiVshzZaXwFY/nEc65KHujuWOcuOMDjRh2uXz9TD57Te3bHUV/JOnLZVDeq3GwQNhALybSPSCm
91zXe1C29NZNF1Abh1eVK481xkV7wWjoriAn3zmk35vLDcacZhIwXrIBgkSv4yuWsxqbstNVQTmH
bFbjmqw9Lri1tGaotbXkxluq54a35AaK4QzZ+srkjqLZ6mP9TKT19I1OwzadOWQ9BvT6TurXqMSM
Bhi4j9WP405ocPPgTZnG++KXiXop59E+eBO6qCgVuqifRWEgkXUedR8IslrIPUXssoF1fwOp5m21
iPC9vWRCPgkXFCDx+GrS99Pe5Smj48mwUzL4g/hKbRHcaXiavkh6XCLtQ8HO57osRyiUR4a3/e6g
EqX7cxc6yC3Bc6DkTNoebqJWp8tXIiY8moHS/HM8pUNg4kLurkSrOw4DGg/mxXokW7ct+wxozoZt
hwwkjMcwpE0hLNGmUidkn+U1ukewtYi1XxHhhKXVF+dRR3sKt51WY4SL+RX3/fEmAyyO7J0hS/hT
pLiyFwDxGreYWevFdCJRkI54A8PGnKxHghr5jnhKjloOi13saT8cgq9eRFBffXSYgYQWvpPSvyd+
z07ul/Xj3HeyQOSlqVZhkvzXRHo064dJpuBnOxmSRUVaAm5vGG9VAQAvIUhIyliBhIpN8tYQMPQx
v0mudoYHjeDjkYE88naVYfx+SYWixjyc2103sdn1i4OKQw7tRvV8KImYVQdOrhdXkXlHAKi3ZRX5
1yOvI8msnXzf2BnchjSs38gyvu/2q2JsmOuuB/mSvIhdIG3nXD1JGs80zaAWwP0lTSatPUfb2FSp
HMaVwMQO57HAF9QBQDf75gYTaDjHbU6eJps1M9zdEHTWYi1RgdjyGsb7Jb8vixWl+Vtv+6ZkC4gR
K+1sW2rx0OFlWybhuIROc+khUVrfx96MiC3Co2sPXEMx53AMKqM9p/ilZcwlpSMS5oO906RAu808
RCK7rg3Raytv7+2hDK+dKs9KR2Nzqe85Hh9XNtArNTJjSQGhLI2uVb0clE/R9Hc2tmpXv5qt0XW3
NjVSwatxQLUCGNrj+k3sn5To6ooaNwVCtVK4vgK98M8PY50RondqXzGwTtWNYWYj4oXvFMXmP7KY
qaLLekfA/XjNtpQdLpVeJwEX5VXwfwmjcsxMvMnKWJkdZiwFBHdHUOgUrA10lviT8PatZZbnuHNU
Wm2PphaW1Eht206UbHPxSZDKCBVcB9cvsPYEDtCXLv/nFmq1bkNoEhsjJxahqMA22vrPEET9gu6u
kxsICaUjegUmij+Qb+a3Q0h3/6+yxtOFxK4rY5FOXjZVLgcicaoXXJ1t6CIdG5++6jGs1lGBds3L
jWPAuu92EffMP+RKE+KqGh8lgux5ZqA664yeOWzolXMGxPZLs1qi+H9U9ovEDv5dp5aE7d4Bliwq
kb+XzXYczyTcs3koO4+okn5/gEhmwY+lcbbBnanFDMmTpwgU60nb5USjnC4rKd2UjZHBsmMm1uH0
HO0gm1aeV6BKJk/GEtUMczmXp1qQdJ36i2L39gSeyzPcYbDHXZOf9yIwtPvxxP7EwYcosqMD5uZk
mU6p7Z2XAEw7B6LlXJgwtYXkD19T22p1wETkZTlhVjapPJFRNe4VHY0kQLnlVi1Tf0dYfxiGS6j/
F3oT5W8EMh06/DubuRfttOdl/r38Jb2p21f77CZLdr1mIhSIkJ+5Yc+/k1hlRNvvo7owKvkkkwBJ
hUDzhiWOyBx+ODajdCHGsajo2f9NyAOc/5TZuhNNZ8MK/VE+hnW0qriKqfsA9RwFgcwbk9L2c/yR
k7mIPGu2kAapgxHdVrc+WHm1y/B5lW5a1xv5c0AwGuecVVnc0PWQPZodmV2WghIIU1t9a+8iCcAx
f7PvxFkz+0g2VBIUCUsdRgZh4uYujsIWerJC9dz7xheIK74HI8FWqjctgTcpkKwI/U50SqbjsKLR
Rhz7wBB7p0G1/pJ4dVP/VmGr8nAlE2AGaGN9UZDpsh1zeYDGIFGMOpeL29f8uIkhRUQW8oASShU/
QlFf+856stZ7eWfum+kuRIp29f4usanxVIeSI8OA0lw7yoPa61Hai0Jcju04M9eS+Abak+snuWba
MVOi1WZfVLMEaWFumYlGGvfB1LF6SeZGRoMn5Sfl/5rRqqLVp0GRDjDJ0r77idUvhhKfa3Jmv/mJ
ScyDYP8fvwYK48+KAUxSNceYTbOlDoA+PBHOFm4Yuf4/pQowp8yL/Y5Gb6YOQbkK969Ajj97+20/
yQzrS4dgJxBFm4A1LCFssFCnkgaq3WVPtvhncQ3oXyTZyMQzHB9XEjP97cTlrUHxIZG/2Nm/wqdG
r/kAHhoiIZOYh9xEMmjw0fyOYXA7lSnG824GWyWCmOyA7rzIblgCNz4wI1R5T7o2KDpGhraqPfq7
U9Ua0VrdyXYvZTG8tLHXQNti56YLFiZveu6pTjcCmtjR3gvmVxPdu3+CABDXccssKVl5Z01ZC2++
fugmtBUI+QAxHznZRYt8aTYINDBDyDeZFvp6E9xASLJTfU3WMj90t15dEgbbD3CbfE3VUKiVCpw4
nZDmx1lWqReH4eEoKnOJXldxPxOJ6aHawpIOHbejXhnjKePo0wIurkIpwWNK8Lx5YNYl1u+cBAOI
sLMpEPF06NrAh2aN72UYIuPAhvinDor7l4Aq3fw7AVhatR0smKyzkK6Z4rtnd6hxdHjXSRmehPMN
oEvxB0Wnimyak//axPJkQSRZwqwPtxUsgMPNKkkT5/IptlrCF5lvZW6ONXjSXK9+NIvL7hOVgfnS
rdIXHxj6hxuyQSTGscdU4qQ/UG2taxKDvbypTb594rFS+IOzjqyi+e9ilKkq9Y7rBVC+CuYDhKYc
as64L2lqjDzTQEQRjh90Aoa5pI9IyToNVNtHBmiJz6Be3Qd4TKYUO+nNYmacbv1bT2cwaMElriZG
2YAHF45i8LWS8i6ru4gB+7RV4SQjaifBHQ52P1rFtwtF1UjATxvMtWjZVHk5wLEsWMc6W71b9oUQ
NabiQT/Q3TnPZ02HB/qjTHO91IMAczJ0jzgH7zgdd17ndhoJCNyfWyYecVI6YjYE+h3jcC/3XV4b
lcQYkWJWiIhkOj71TGkgk/Kh4nCgz5e0RyquUq6GpOTfTa57sTWNXQtR/WFXVRXTKdHVNoqbKnOA
KUo3JnH+Tufyojd8BtsY9aUoX2TYTxqnqTVlDyJcStLuuOnYj9DGvWyziraze5TU4Rx/4MBXMkTD
8iARrl/aQLAUn6Je4jwZCsy+o+NQXSnYGtTx+6+JjsyE90TpOHL4GGBsmcd/G4s2acy0vonVT2Am
xTo9uOa8KoU221gP0lkdPXgvQZLqphCqGarjBts31JYs/SALLoveA5mUA4b0VPiLAVXnppHMQm9x
YB3f7knd7H/LEnurat1G9flgDTT8z0QOtOYjh3g1h89tJAQajmLrYqFietmK5OzcfRuWen66EyNy
sJAzQwqMCG/kcfP/qK0wjvbmOpKodyPX4xY9eBlopYM8X1yOSeCdI0Cq+eFIEYhNHT/FIO2Q6GEa
wzfOxnNpVhAKadzQWWS5ykk+y3hi7Mli4UQjci8T0Y75oy2XgGQGNBUbHKeYrHQtmfmz8ojc656j
ldc4/igikZTQjyWa1FcCNeQxdPf2wm6qmwzP9KgDm4ihPxl31kOjUvb/vg9kLhmtNjkXzxjrXFvJ
8SgTRNSPVm4bjkxrjFNp6U17yfe8NQuLXZSQVAn6Qtw/5FRDQpuJJ72G7fcVvD/4HnUzWkNXaYVZ
KyZYaCHKwqsiP4nCbJs8ZQjZ3HWBW54FXatvWbWmxvk1BSs4jOpyD8Kkz7s93WhqkBsSJN33uMtQ
arcHPaK4ILfrmrk/4lGdVmJigEp+m1RnPqmTTsK9WH181GgtY0jiqhPcvozbQtZUKTxx1Y5SrMWj
tVyxyaN0BsluI7fDsuQ2Cw7xT3TzObCNi3iz8u1B1gGhfTJnlRK7HkXF1LNG88ZS+9t429exjII6
zJqdhtCZTV8UPWDy/k4kz0Ey2HTxbg99NJeVTS7hwV7LBpOEnrfbfttFG7F8bQB9YXdbiusPbNSZ
KtlmdeV+7QUaKEN/NO+Fp5SsJdZpufdgJIP20GX5lZTgJfn7WGaBKNJUImFNma8uEz3QioDvra+R
Eugn2xmu+rNhKURbzxZNTyhDhnB2bESp9F5lKnuNutt8pbiSPCF2WonD/WA6A3yfVKGaYFX4tk5l
CPGxIy2M6JTNn+Ov1dZZdHS4i+z1L+4xzFyz9nsN4MXYv/Z8AlfMRyybahoonMPbHzG87Em4b75K
uwQOQzhz5+cP0gwlZri1JkqqyfmDMqgMVL1dGY133ZDHPULSU23chXR/nsz61IPzqn7jIO7bo2cM
O8bYDZkJ/93sP+4u+ww79eIzQgEvZM5Y3ZSpwEjAbgHoesZabM+aUtBi0fKWurB8lHUWWMjt8rAs
TB7qDjnUhc3mtp3wtMxIaNoixDvBmso+dZX6El7ia4RMNd+98ulXC0huRdvzaFT7gbOnLrXyXJBw
z54If99NbGup05exq/wLVziLnIiOZeHN/1fj3qCfyTRy3rl8yzsGNdW0IQPyo0kRBJa0NFcSc1aV
nvrJNg5Px2Z8L3wV3LbESL5bSn1TMvUO5BtWgLxb3DBpEki7PFRFMqbF9KhhownwwVLm/w9WaSbT
rgrSCEeru3HIyijwCEDBkfzTAAI4gmHRRZGxBgiZXtd/8CUETsnreukaO9WdYEeJmtHQSe3CgFou
0UyA5eZBk54dKCIWoWDwqQ2Ds0x7CPYTpfIQSQrONNhSjPOLvAwZxpDEzdYr7y8u/T06//dbD1I4
5bUi7+7P44ZZVWxVbOpWgvWAudpl407MyLgBpZ6+3OdjweJE51gCtT+u6eub0F/waVLFTG5EmQVu
eKztBDo1snPKtZOHywr4hTMTgvHUP75jcb3xAcFdv46noxIfPBQUpQwNbJ3hXOhJgVyiCpAPvyKD
nA9K1S9W7qjv3I9Rlho0RkWOixyGrrVLYUlqpmpsm1F9mSbHp6sUzZsxdDz1E/vr/GoOq0XpfKD+
J/R3LoK8TSSecHYmR2FyiGTzacH6LGibiUdjtsMUOX+5UTXAP/DPIahV2pdbCamG3oq0V/7Syan0
U9qc6xaAD4xW9vlxYonXZ323eiE5NjH1V5LTr9rf/mn4IUTfwfkkeVMwNs0v7+j2Iu4RJQx+k/y5
AvZ8UqbSwYkr1ZKnJhElJanNwV6v1Oaewu5L4YLZp/+EDR3sxy9wPvNiMVmYzfn3PpnTuQmFB+q2
oao2C78ahCVTbk243vAAX/VUXGjg+sa2DrAN9xpmClf9bWpQbWg6rX24+ikDAdIGqV6zBku54Lhr
N1h3CM6NJ/77ARh/3n+/Ig6DufQCM7z8ZzhsF7hPKRaBQcCg5V3bs0wlA1kPOgZG44U6nfxnBvr9
gGO6BzSuCpeh1o/HdrhneHLOB8AWi0CiNDG7Y32ns0h7krkMDnx5DYm2o5JkxC7Onxbht5SECa6+
+bXxTk4FD5uM7cXX4QLhk8wbZowmB6PIHRtuzoFoIKeAZblDLvrafxGBsiTvvZeQZL/p64kJCiDF
mTGE1jYEQq9Dwoa3gtbLzjNgD91M5QLSgUUA6DX0ziX2MiV3/F2XmibQ/3KfDMucR1Ny9/4djPrt
pRXz/yN1UATgMLdHAuzFIBcB/SOTd3Ee1VVcVSrpb1i124ovbWqQHwDON71rXhHd9Xza1jUnXsSx
Sn/odsGs91ClqcxPoIb1N57yEjfBiqgmZMKgvDl6peYl7XEonD12Uek6PIkN07oD4eD33ZambeUD
zFFlU3fmATQYnfal7INW0EU+cGbdcmONf6OE6NIlljKXNKr1gahQLSGrC/5l4pIrfwA3X686bp6A
fhrkCkOiG2FL5HDhUhHjACbVxUhdE4IZrruZIRlLrSTuYfNbWthVcQbEKBWsHYsNMpyCDqadqTtn
SlXwXewUvKPLi3YyCIjfcQ93iEe8CaOzPRNo2DOBwb/Wg9fbCGKu5ZdjhfP597WBILCpbsAXHOGI
JHnAkp1ig94k+n7PSMTdMOzU0N6/AlH4el/BpLsxSQfoE8EmiSBWuRAWWUHlbbzbRWEE5vYrVG6F
zuRiGY0TdnzUNxlXk0+UkJqi+Nsl1yS37csZvzqellU24FUj9tl1lk1BTgB9lOzgXi1VI17Qd9Q2
HFlM+qkc99vNFGYxUEIXM77yvQwOASf/nlFp4voJKnu2VVnP2M57W86QgWanYboUy6wUr60j1lrk
3jfJFVQV8n6RHYMqUMJ9daPwGDRrwsZruks6Rrz3c6Vbs8alyX1wtlKeyer15G3cOsp9p3mff4Zh
0oW0lvX6stG4MAFuMw1a3mk0KXL+v5dOL6vWlFldc//NONrer4XmVVR+022nxgZ7+3K0KBGRNQ0G
nBA3TIlNDg9K4l/W3A0kK+HBrw1Av7VxpdWHoUVnvPC4aBsGKdcDCrAw4+VjE74ATCtGFOB1Gb/r
epyH5anO8gRcF/mHvRnhlqPGOTlgVBIGtj5nu8fXeDogp3Cf4VI931GiFhzJngzKVksedd7ItGDh
uYFr8s+mlLAFLHBIkvBmgAMz2zUgnLCkRRbVLkN43jdv3W0Ek2Sv9xcx2OugBfa1EFgiCZ/R/fzi
CM7K2c0uLZfmfuX4ehxlJB0ddYLCqSEwtSyjFTbD9iIsvJpm4nXokgaf2ccJwlDu5FAUDmy3z40X
TeICNOnBvkEai81JueKi2oAmIbkbprA8PTmP0v9ihSJ4qGTdZqr1obiP4yypMyzhVMO/yum5+R32
jVM53wyT4s9GjDqG3eoM/UG/UzTSmpqno9HwjoPwae2v+rEsRuk48qOpHCa3twrnCEjsaDuYL/mf
Vy/kW3U8M83whZXaZGbiSEpWXpNe5q1aasfamIfhmCPWU4hUKuTCjVXTzgZjCGzW3RZORZJtAme2
6vaq6R5V2CH2i0OPnhXk9vkZOpl+xj1cr4uoNXZN2KPBU4TEI3Hw3zOqWlySVshc9vqbJuk8iYzq
n84my5KWBZDfO3AZeydoX6J3yrFITSpq7YznrX7EBQa/+AH/mGA8aAoxdP/AhAz7zWHqIbwmQVaV
CngbYPI1w1b6vcwz1kvyBK2qK7P5S79yHxxwfBlSDfRPCNKnp9Rwbmd3nOcPF4ue+tMYyqwUCOUL
/64RAt2S3kADiUXrcPojpIc4+TAS2nwOiv7xbN8l14LerkQbFR3NrKBgBCEjD4MJ/Pp8l2eWvGnb
XbkxDVK196BO1F7tlaZ7LcLSh+smbfSEpj+bfEPLsqk8EUUzX4ShNP2N5ekHdyxNToaYBSYubeBG
GR/nrO5XlT7jzxCwyAtBO59DxD9ePNqeuuTlsTSNq98rXr9a37nloohOanF45LcmppIu6CSDpWTE
27DF1bCI/TrV0B0WP6BlfzSFpvUMT53gfXkztX7cc+phdEVvSILI4Vd4K01yBpblWG5ooZ8fpAHk
mO0r6PKRpis0nBydOyKP9zr/b+milaWaFckVjQvjnrB8q4weA/asCf2qSr43fs7AqB8wz2uWeUiS
T3f+f2uTBZnrdBIXuphX6DqRl/XYNsH3Gq8IuqaNV+t+OwsZLKIe8F4HEC36glt4thcxGX/nMzDw
jN6pc60HqPG0XoUkfDQ+ouKvxJV5uuxyXBXaWVtcoc3yn12ZNlBqX8zuHXlv66Qo2GMFz7C2Ixf8
5CG83Dr8c7BKLX7CbJ+D0i05sECpFbIeQA3HbldpMhLtHR2FhGK47CUvkrFC1Z3s+3Pn8aLheG4/
DKwzhsICR9Qh04/Cc9+Lm8Upf+wud0geX4fMjF2piOTXpq2f5aIvJJ6dMvLASbzBmgIBfU40bs0j
a+38p8OpWluqo94htbGwFtz++rvibUzeuzxIjoUdfye6WAFuhtAYzE8yp44G9q/lJkWjyFNMA8y8
6kT1ErpJDI3GAu4+Dwg1UisK+REdxVIlENrM5h/3uTQvDe2Tw0Ubs9hpZwg7KLGoTSfbiz+jlXim
dOJ7H58Z04vDCv0gYaagML81qWCYxrG+JAuabFmj4tSaxVfpp0VJAyz2trRE2k2jnZPzcVJeCaDJ
JxDYS30Ic3MPlNL6jZYzkrM8dPIsvQWzjcil0B/GVEaosi08W8NaK9aUJ5TK4oF5okgXHjwuc48P
7w09OIbq6tkjaGMtc/l1kucSUlOW2IM9aR8LIhsNavIwU2nDhkz6UO7jo/aEYQ5b5YsysUtE1dNf
DkWqhXyd4PLStAaykhH1g1Cmfq7sGyPtze1OdhgDIzVuiPiyt97QmxeLYr4mmmGu/hDhBRlpkmI2
bs5YZZ1QZ/I4fN8rpAqaCsEOLiRlmeT9PJiNh7NLlNS0WZ6w88RRvIh/tR3Zv90dvp2gloe9wevH
JO6l1ZvjkvwJRdykpg16mYfXNhPuPtQlJfOxK726mNbbRV5NWMQcdDYJHeNJI8kiBip+dZpbtRub
nuVVJuUOrvUz+1BwH6/Mryiu374NxKTrhMbvTARXopUaZYOh6oMopn0oN41fnyS/OJqi6TcO1dG0
mZBHOBX/NkZ1T4uqyZvmRCA4usojbhHv7ACKpf3TeGGHTfa/10V2MDuM8lA9Dt+RRIlVyDvsN0aj
ytmBOxYnjKa3zY5OWaxC58Q7WD3ZRQsmOrd0lI+FBLfaJrHV12vPXDO/X79ARu+FgcJxzW4R6IAa
UoF49AzkWPmfIPsymkmf8v245N46DkSY0FgBMVi1MeUCuDA8NfXu2E8zGCNKzE1XN/DDFrKDmhOi
vXfpeYrktgIZipUvRSIizV96/gXfqQYi9J19tcKab7q8VlgTOwe6YzYl1p3r0n51cCGvArTjCEFX
FTsm+UQcjOg2+Ebqgzz7Zi9Gm5200M9lWDZhIAQqDOa3ke7xgvN145pJ4WHYycj9wOsDV4QDZdiz
o9yum6md0lujzU40biW8kJzygaTa/+HRMqcooxGWUvM3JkzUxKt/Zp04GA5A6Gt0evXvk+X+R5IF
oZfZCyZdrUKF8beTLHK0CSTKlXsLI5AwD1gTUkM+i5Jguvehx07VNxRkoHVzVuxriJAuxz2/EA0n
VNcgPlHvb9mbnvs6x6dioVyci2PFjsk05YCFL+g8M+ACKg1S+E3wO/RsCJ5dBmQqCT8bnha7QSBL
wea8Mkf3q9S1dXbQ6kcV7NRomtnI4MIhFWJN+c9H1YCPGNDoYAo0uTDcN0mVgG9yqaMYMQu7WQ+6
+8xxgXQO/aBmVjKuaC1MjARXDnqHsf8V70So+xH5vNaYIUB4XY8KniuJ76X3DBOmbg04eRigCmxD
PvtVH04tGzBOR3zozJnLMds84ll27iUwi93qJ5CmHZoieVwD3NEkqjmbfyWoIe5MT4loWBi4v5On
2fvonAhGtk7x+UaKaF8/8mHq0mpVVE2yvAkyAEXgHggcJY0DBA9flZTHmTHYzyTLQLLuVjpUxAWu
/EzrmsFg8+ci6tbmcAx3AR/dUsRzYhCvfI1DNbqFOBwXrfg5d1y8ByFi+8P3mXij+TYPd0vZ1vjB
SVc5Gu9UP/8JQ/wO0z2S4L/t8wzCsPGUsxwAI5jmKfo8sF3u69dtPlGyYmeCddSMhI0wjGN8NxRt
h6zczNKVhH9Kvkzo7yReI8CAyaMiVQrSmx8w3CNCqmpzQyw5N8yzXk1us+0Q9S4pKobDtZ1i8EgS
eiLMwmRuXIm8wXWHaCIjcOOHOKzIEdDZ5l/gAngTgPrBQ3PwWt0gjF+KZwl3IspauIrSMw+hdqvu
U5VpAJYpU1ALA4e8HGZd/f23WjO+yy9LaiNcNlJ5+35kxtlK88/n65VuTbFa0DdCk2J60lkZleh5
ZRMQkc1K45ZznMWdnzUyZPayi8s/haX8EuMe4gFfViyu3jd+bEwcZGHWCFoBFZ+y+J8kAtYxFaQi
hq1iGzbDk4NeGQVowc2AM8vnsW8ltl9/wTTlMZBCqJzbsn7RanIY/g5CHp9jdLMQICj4XwkHHvuM
bGu0x4dQuPaLxhllRHNAyvwm+MGY1i19lFp1j0y2ED8AZNAgbHLFnZvqE7BHoj4B2cKR08XV6ljj
LOB0hU1YLf7KB6UJQEk8J8OU9kXj8NHAmKVf1bdrOfK17kto3EMzz6bzKlYOrRHXu+SFFhNyZOGL
756JB+od2y8uC/6YjMWlYy2fBvvSD8//MZj0QAOfH5Hl7WZf5NPOHJZQBPul3I90hxteKNmxCKZ7
/GsRHhF8/IMX6BPwZjgcCFSWpHeRMApQcHkiod/if3ZQn8oXSipI0IWoTxO3NQPgJyM32xA0l7Wh
HV4A36EJ8nsnT0hGOh8iy3nKR6cgt2kzqeSe44VdSybp57jGgNJLft9HUf97+2WFKiPksvBEaTYy
avfruBWV1qLt/dr/TNV93EVBm1YiMX70gmsXcVSb/4EoXN5jrr0uVEaeNsR0gVc3MtlqdmaaC7YK
LrI/5Pj/R5iE+bGsRWS8wdEL/3D8Qh+gw8Lg8LapCV3Uukp6vxdWCNcLN4qZSAqPtFvYSz6rp5CK
IkfNxm0GoH59y2lV3bDmKM2PaYAEzj6Q3/YEYVdwWyUN3WWCwfxq2WkCv409dEvXbvyQlVBUFHPk
DMMpV3TC5tVBVt1tc7TTSO/NeAH3LWIispmAZUCd6xIunLtnFs9MR70Hc1ApW3yCXh550sJtSyE5
o3566MYUJeWENKVTZY6TMCJ24NOCAThzb3laGuK9zgsKx80j9McEH7m3rHVCYLSTTU2/ZXPjLvof
tBGdaFIfT5UrhDRKMa02Uib7LrSDcwITbzmuRTNfo153pMAB+1XjF3Mn/qe/ePO1RV9UdQ+lJbOy
/yzF12mCqgrAXW5Eb5ZgB4tTss3APWDFe2FSztolyjnYU6rlawEHCY3gfnypyew9kIK/rEeo7q0H
G85zXriMKmvMqqhE6OxIPjW05Y/n7ROqnUaoyckH/0esuiB7cveFDtXALSOzRHf6pgE8CH39X3qq
iccpLE+vhpP/GP9g7fkmOirk1hmpwSVYb5dD7aUHdR1yXDgQ7JR6euDi5jvEYdlE3f+qyEzafzxe
6kl4A1xWgHcpb/kpbHJedfLvSAlGhvMAHLb9NsJob0ACDIHov9hZoQhagF85gmNv+WGuFpCnexNX
aaKWw/vBZfUdD3MwPca0anD39BmJMczVhuLYnJFgXZi8b21N+tmyJzb8M6SeLsYbn52ppEu3e0o0
u+nqPfTmq3hukhcF0zhHR01Q0LZaE2q6NQsFgWbd0LfB52sQdVWg/qu9xkg+T9Uk/I9Oy747imT2
HzQw7uvks/o+1oSkleYDaHO4FDjm1fg8SebmCWryHnold8cefalfGVEYw+ICFiGimFh2fykAjqsC
skCuuwJNJibmufLSS0B/Y9WxXvG4cyzLnt+ovynKKpuAawd87xXIm6LHK9rcNu3Z1sUD4jnCckec
JxZyw4yEdcDvSUBLytgcdt543lQvIm0UMWYwR0fx3DzulK3Hi/yjYWi4l4leG5Waa+pltdZqc2i0
awWADW1GYArZOXPnbnzVFcSyJSAbzFozrQQFN546j05TNtc1RKv/TSkHo/dCUD/UnwP952bYJTLr
gahOOXRYxvNvKyuFaSL+KvEX/9wiUPHbmGQr3H6dSE+ZTUhv3aB9AbQZLv5OZX/e9cD+R2oTjrBh
DtB5Evet6PMJrlaEtupgaz4jwSOan334ReWZJwzRmOw7LMryhBl8RW/MZ8w1LLMBC3wX6JY6HQpD
TMYzKeS4UY+5yd8XtiorN334oY/SpAhjEHW8Rtk81NOmn00M0Q8+4WnlwYUCd6dUmh8U/6ykjLlX
plDxqgNnGP5GFY0muQmPhnloOTjQ4aK2xXqdnuVfWTtrbRC7YBRN3SqVEyWi9zbRmOqhTCsuODZV
gvKDyVCvBRceTu5IC6je7kNKVpvk4WUDUdGpTs3l197xT5ABcBfZgwnRCuNclazH3wyBoivdNvGo
4y+8mTE6fdZMbDcF2TsXO/qp1pGXP+2Y9y8tvujPPb7Vt/SfAuGTRl9rWRPLEdr5w4hcFtChyGAD
VnnGAXDuRLJ1tZiuVfPp1r6FLECgfPRWhlYuuKoDJwpb0MmlOnuNwtorWv1SdQhw+6np/Fu94iBy
Vt4TvTNlgGSVpuLt5PAhFAaTvkgIabr9M3lAEUVnLnbmj587+Sk+a8VaBi6U9k86Rk7HL5GMf9Bc
+hItLeEZ5CtOcZNZ3FPz72JP4hinpkHHDVrxKSSpAs66bxUMUNQfTXTt/3FCyk67gkxDDiTLxYUE
lCB5qYiOGJyJ7+F+0Dhal/VshaC9x7YtyhnTSWgUAt0mFgeGVFadjzxDmsoEHOrulpXiUAGxfMNj
y5Nv9uhiKmmkWquEfI+CnTBlFT0IBnFmNHmd2UaSTXjzaSwIBO0m9gVsbrkKB/PtbDwJk1bI07F9
EY3QsKkkn4XbM7By7iovl5fKqVrkZHw3yCCAQBALFgAPRHdxMJ38/lY+1WERgA8QXv9ZhlVfMORV
p3SGD/yZlOxic8WzA51lHSJIkG0by6CnlpkGTTRXK+57zhciNQ0BLUjUgIYsAVbjDt4ydCrz7JR3
NN4sDxfx+VyVj7hxdXeW4wItBhXkYM3v/JOQ9Slmi+wDX2jP70nOyEHly7/NQsXSrQRhQ+RhThQX
mVEOIimBUofIzl6XUe2vy26Y3QgZIjorjA4gJsCqEKCcaF9VByezfo88RNW+70KJlCImG6JhJNjk
OzfVhU4jrnCzu0PyhMyOAWJxe3lbj9BV4E0YK6pppkXeqMY0345kEVEKcZPV6cO9qqznxvagnWru
YYi5ZLTktEFyBR7YXwaSaOB+5te3Iwf2RvtUR0785s2cqhv6EDtzKfeiQ78FLBQyOAxHJHLf9c1X
sEhdRyZkZcVaaVeGZJNq+toNxn/CaAGgvO++mlGS84rCaUIWmsmwhAowkj6xi6DELKaO1n4aA7/F
jdraI1r0I3oBzuergk/X91NxigtSL3Gmwqu50VRUBqbDFHHGkweocsmsyKJtDbR3WG6sYMf8bfzk
tM+Ju9tTs8OEVXOxctymyp7jcZeBCIzRs23qQh6Uz5StJVW6ebr3Aid/Jh3ghVjikqS9GaivSpF4
uv7Isv7VPbR43FZnBlGY2rUQEuyXZLY2FjZHNHz83bEi73zlv7kmd05GdQ3yKNfXT3z38xj9RUNP
5A1bbiJO8eDj3dX+XzKGeKluMw+zTmXPW8VRVp1CkFnJFpXHfcKVbFN6mm3BrcU1JEZjeyl+6rFX
SOXmw3K8CkIITzGdHhk1uhK7kaJhy35+JhCRHyZnE886iMyyLbZMwFhFQSAivwRmdgmZqbaoXfMi
Whew1zyyI8V47HDlgQcvwNVHpnzKI8195/ekcgvCGTz/kmKq/8Mrr9ZULXYZne8vqa1Um+ew/2PT
Eb92Qp+B9nMrkMaNzI10LLlRcdLUEdt/LsGQ92iu2e4RBviAD7g+CqDOBeZni/DjgF5UL/A3eMFr
M0N/qDyZNtgH/ZTznW6++TGYNUwteGUfhYFZKujyfMLu7qmXxYu2QHDdpGXgCIbj8jjBEfpXc2Gk
RO+f4HdSVplUMpx2HOeAe9jL3BQxgc1LyUqNQnAk4xHZXqHwdi9vcskOwamR+98mkQdOoOqFwzSo
lk8byw+qywOBqe8uGLpqv3QgsaZ/uwL3C651H4/tpcTvUM48i24DWW0ln8QTjcicM6cjdODe7EEK
Iv1LkokQP5Hyy86pjBU4h+rWMRr6tZIajnu/6kJkV6QDdMAVzsCWaJQUGq5UYuOhDn5vm1snK7UM
RAe3o02BvS4Mh0AzGOT+uU6ZcUyIqa24OXrY/YfJ2yznskBFXz5qGsHg/EKP5x0/L6FNceU+GJD4
gO+XMce/NshYBw3qbkBL4BR7rxFRW1s/oSdxYldCshbAif0INU3tcTjxL53J67csPdFgSfo7dcDb
ytIxBQR0DD0UjrnJo7C1uCfkb7IiO7FxEAJG8uPE/7gt9j2R0hLl2ddf/Y6g2AkqZOT2vZ02vUkG
we712yMlxBMz6Vph1uG8Y5oKM18ueQK/eCBnqH7/+DDtUC/OEjituatks4Za9VVBBIGZM5+ulK43
lkQH4w2AOwyewo+0B1QvqguDKAmHvqG0y7iuncYS73C67wNUDne00WZHN8QeFglSw06mbQU1b0al
ItLvFv/dBX05+CckuI4yZiyCDhjzBGzf9NraVlP988nLDtRbucTCGK6sLwasOsf3JE+26QzgssvB
hbCePPO+xamQ2useCtM77gJM4I8W8MxsHLeneIA8Cqr/RPOv2/8+/5JL0ZuRuEhmgXUNOPb6wygh
Ya/UCfmk9AZBWGcsti2XuaFGbQdp1ul9qQVKNPtWlokn6K1/8Y9NDMUl6IPm9ZMt1763F8qLMowD
OxpgmW2BCPX1w/VfGUfU+yQwZjd+RXflWQL9JoNGYiP20PbMkntWSTtVaLRnc1wJsfDs0zc8f1R3
NQyrm+bobPtR0XmkMBRzTCNrYEEmWwv7CF4rZiqIyqlzFBKtqeb/CnXM1EUgdTgtuwbqcWfp3h7D
OHkLjD9Bp2bmJj33n0RH0012HkXJODv8lltAVvF8dEsZjvRHJ0K+akrhJ5wg+Zls2cgYLdtmDGGo
Vajs3fGV+QD75RSt1wyRwOXcCyShfYAXszPYPjsskTTDRFp7QlYd96FXbNU9KG42YiJyu3GMvCOT
/OyCmWTqT6PmoQYOVfvfmcZpYcuufLvM+CJkdAgdiR14FimFPo9c4anXWWXm9yl2UeUG1WLh/Hq0
F35oEmjdWSZg5taQ7gaEoVuvyuZq5E3qEPAUqE/dMH/1SyhDNHeifPrNYiDgqqaQsd+qLcdeQqFS
v/6pRxSXmUAzCyTQc6ocQuk1JsKKC3f8Kxo+M+MYTyc39F/PYJY+m7Q8tq6FqNr8CtvLxK2Egmc+
muLDwbt+hByoCMePi+nnpF6arDwCuboeAmS13BgOqL2VFdne6GgjIukHiOXQMlbz5q9JYEn3HrPF
baqggv8RFstx3HhOuKr0hDkJFZDQ3Vz61aYYgzhsBsa/c1UBh9zJIJhqIb302DLthTQua9PJUgfn
zy+8ku+hQlawOd6MZPrai/l7Ta752RsXgO3VX7MZudDqVEIKoPclx5eaaXfiRQLenmVYu/ZNg/xB
d068B0ajAHqD0fFe4NYcI4G+wwFR1Aiq4GknTzeMDWp39dZwTOSXB7/sC2t+ma49WS6pbVWHMB2C
j3+tYxWymw7WxoQSDffgUUYocidJo6GSChUPSxZCZiwU9NUHYBya7Np5mmxKK/P/8Xkr01eb2b4v
41mN2G8a7EKNp0PUTtmVqHP5ufcaC02BFtaEieFXwOoU1IqV2gKqhNKGb8iP9dCKEjqKldcNnSbO
8uXRZGvdfLwf9wP4OZ7YRNzLqjncvrIhe/atx+yIzfhUFlpctzW9+CauAqm8wz4WmD16PGLr5axg
b2kavwtAk8bmmKm/8Hy7fMyMgJfbnOgMKgs9itTZTCPvnT/a3Qk2bRqV60zQWhc9X6iXoDjXOlgA
+RaHYGBCTq1OtSSGAcqkDktvx3TkihdhjNDXK7enpEGPT9FF82GWHRYiQlCbNNS/1ej7E1ackvxX
OD6ucEeCKCDAilqwQ6drvl9quhoiVIrqQbHPrljVWWYkvuO9jLDoXUFeTZNNqvBBUUJ4H3aoZfQO
78jH/a5mhJUXiQLttJe3SA+2C252OSqVcJtBHArt8WWtXFVDEC8PiiWHvMvIpcRIo2WG7/8UgKeV
lnGhhThPSdoG0MpUJytrQYWfDyGe+mwcGri+fu9SDOL79I1l8wZLMzI+GTO6gl0kn4r/WNQVS6LY
yPugTVMD3wcO5U8lp3rOa7/g0HPRG4e2wsMmZe1k/6Qwl6j2mqw5bdOG6+u1GFVTE0Bzv/PQRuSU
6rVkJsCxLMP2x37piaWaQBn4oVQSraT/MWEJqQBn13nBXBBjtAkVSLC5OSmhpYycMbtg/U5eJHbw
kuDyzKjGqQ/VAz2giMGf4f0laYYbLZraGvUllUhTnoAO12EISSVW+BzSitXeBKUtXmEQWTQOP9Hs
0Gm/DYUI2HpQzFW5qYWSG9gGrFU//QZo6SNFZAMDaysvq6OhAuRY0Gnd3rQlq75AQDXE7aRhioEE
ZmknHU1+P6LDAAoEHmXiWnHIKdlyccKQEjFkPrzS84Y9SJMfpj9S6WoQjgT1VkkrkesqtJojCdgt
nCKCIQ3TdMk8fl82grC9ACXjkbjaVdJ5aj48pM8NhcxY1NVr81Bx8EEejec4qekLUEs1RgMEUMuZ
XuMF54EyCqa97+PFaqAujjJtX0QJih6y1rSmiGhOaN+2ecRpl1UGV38O7336kZ3rOpOarhDU7u8q
DI7K++i1Nc2oS1d1JRKeUxnI97oZnNhH0h5GLH9Ugyp+T7Wq92lMCakLe+kQfST7N8yoJjskUOvb
j8tzz82Muwhq4g4Mwn6m09YVALwbOnTgltht0dJgyrwAwfepbquT2xCRSchhVlaTBrOI+s8BG8Mk
rYdNlK0fsArjsvKgWiA/EI5t9TfO+EByw+xD7FXGcyooliUmwGn1sDwvPJ8Sx+G7fMdnS0xF3r67
ZDNos9UZvZe+6fMtn8ymqjlX7s2B2BMlYKb4L3eOxuuyg/iFsoVGR+1rYZJtOWUS8vURZV0JD8KZ
MsNsp0g6wIw9I291bcyRIFtiI7SK5AhD0CHeVKr98ypJ6IcCukeoQZxYHIPx0CRZ0g0enghEXbOO
srMZCFkdXfWSk4eBh1EY5G3G/k1LqjEpUs9iSq/quOuCZoOrgnpGY1BoqhIKMtSzzg3FHVC/8i5e
3CZP0TUqO1XBRaUvU2w+DD7oDw0UJ6/Bg5zhN2WomX3ly1N8GbDP8ANtlHeNtgBtHews6+duT9ih
E71mS+6k+95cyjIA914obrhlldCVRYFNI2f6jiOVCmqt3uz+hIhlHJyEFNGxqEnvzJHbS8bqN37I
13HC/lpm4OIu3d/CmWLT6nTR2ugXipuf0aJq8w6JRAX9/4PhgyEkQWw1kxuZeNpGNBGcRcHLPAPc
JZq6oZBCYBNZEvNNuAL9ObcbfljXAHXfvS3mgSU9rhYJOTGnOXcl0ADnnGfPWEqdWcFkJf9b9zCf
CEffEwV3Q4wRa6sIwqqIvFHB3kBBQCcaSscYgMwa19omwEHPD1iALothR7iMWJ8LtiIJmMcEVz2l
7ubkbZDfokxNo/wA6tap1o9YQmiDPu05caRV+2Ug/ufbg6pW5Ed7WMaJ7ycI2BIglMI7dpVEDSjl
BXzF3q1OrQGHe79Sboj8zJgvuZzaaeOqqMPJoDIHsWz8mdYjZoewv5GTVoulDqeENEt6Bd7eNWG5
qP93mzL1W+u6wl/pNvDpkZtlZ36goHUsqpZhOwtiEPlQ/vHYBxLNmJl8HXfEikpeVMs5wlZUNc8Z
pc7W9yAVZYEOHZIbECufZ0ir/kPviWiq33TfTXCXzgAKf5CmS+7sJtU13R/i7sqNM6qxKo+ipzbn
tTpWTsggYOpkuB33ya6O1h1uQQBQLwqzpBttCeHSKSoWnnnL9wGaj90zkeRbOV17WOySV6hdOZFw
icg4AVcbPyb48RF4yNes77IqS5GXQF/fbu3Pf8ql8jaJ9vXmaLjt1tVK/Sq7MYJ+L91JfLvQX67E
V7bOx6Zei08fEq/KmrhbIRO3AYq4mx99+/YyegU+VEYHtp2QfnU5cs9xD4qD76n30P8TwabiEgwO
tV3KmqJ0yt1oMLFFqqQSJJKFF7cjkrhFBLkGBT4Ch08k6xy/gkSE4d6QG/rBB1sZ8oAU2SUffuGn
qlsrK6aYbEMIAJu1cKdZVL/AwVni0ZKBd3Ostm7ax3z0YIxpEfOzcfwz0GOcGU4OtjkOium7P9X+
+Ldk0qatt3tB9FmQV9Bd3svbEex5WzKuZyMvXK4w7UrbM31yB0/DEdYj0yzZPI70yt/YT7Memy1c
iCvqD+LUsMkW9530oaU5HCsXeJTEAYO1QGcdtLFJi2EBozHhwDRlcmaXPkQt9GA1aVLhCArm67D3
20Ao2mp/ahSMQahchDx5WSHG+t+YZUHSCqCSIBxO5tgI7Sp+7K7LKtQALHGkpBZ6bg017vQ1jdjL
PTuUPgVr0BhZ3gAwF7IW++xKlebp4gakiDN6fUDXzIY4cGHdePLaG32roFBwmREOaIVCix0Q5yVx
Mis7s+gWCTlSF3NrlxU6m4Ko1/4rDqm1eCsYt5lxB8mMAUO+fb4dbsQKbbe+gnOo+PvvgY05ln4p
i+nqcJ647HLs0NRPu8IoT9zOuArUx3851CZbV4BZ310CAcxihgmP7ZOCyoV004GBVRGuwPj7H4Fw
rxE6pNMQkbBPGpcnaRGbwX4KnURoXqnmc8Yrns2Z1EsZ1hp9y5VcmxfdMc1o+6m8bAEvckTNI1uN
a2s5LgsD21z0OfQ18puC1Vc0J2tU+vCMfYSYxkxpU0dHVfr1mbt/Jqkn1yIQkeKkK7MWZGZwKlze
nIvD7L9uQ2sBVQaofKpFZrNf/zmaVGC5QBktgVJa1nZXzGnt0pC7G3n7WNOXikGkQQ2/1dYB/6JQ
z2K60pQq+RuxfAHC6TateCwqi7GTPv2YoBpTEZCSKEWXSwX6ipqYAlkjhRayVggNBwkQNv3HtteU
ThZh2cWjaUywDLMsIwM4mSKisTs30AijJV23koS1YV4QzSO/sLpT/bDelbl/IlmUrMMsq2M9b2P1
TjhY4MKJ+kD19RfKV3KGO7GIEbCbuLhUC34ZXPy2IMbjRO6uHqQZI0ueLHHiAVfopmLDlTIgV1IR
iP8NKVQ57Ws4VTuc1ZzUPD6JGiwe+4TO/mYaHh3YpX5PxAtODddATmhKlYycUyyu9NLFt6VK72SA
rn3uduj9fPXdZRI80N9dwV1ZqNXI3jld5dCovaQQ+pQVEjxM6dV7s0q4MivjISfQ9j9gIrtiBheh
qRxBM2kIZ748RlVjY2haMowx1XusKdF9cxnuH3vKL6MSoqkdPPPr4soH/81rAqRAkKHmlQQcTJRK
WeVQsQrcFp7PLRwhdHNkeyPDG2QzxvMlu7aUIopccsCUEm73yAAkn/qRZFL+yml232rDwTxCr9jM
0sMjnKoJmrwLI3VbR8IHQW4QaXIBK7bS0kNC5gWMtAE5zMMP7fe9VM8/d4lDZhAHkQmEEN1A8/Wy
6oj6MjO5DlnDY3qZy5q1GkuYOm376AYuUvKaTnD3zqqcCGJmAiCmithqb/96SUSTuOHUniKrtVJT
FndQnXYjBcNMGxlhtQaXNJgrA2mTP1/o6HS82oS2Ss7QvTkL2dz38ooMcBqYyJaCmh5DQE++yZDE
damLO9s3w1gmBF5bZ6GFiJh0Opnf3fwdzMqe+aSHaBIhPHoyp7oT5oJmVVn39W3cJt3eNCSt7tLR
+TQM1PbEEFUe+WvCsIVcD9BSKZIm8cHtd/cPOTGEzpzy/MGKtyNG9N+3NdWwyUD6j0edPlhbhSyB
2xzRPyaO6ga+Bq0uFse0sKYVHAmhjkA9yBSlMLWSa0uut//d4VkxcreANUSbjFB9Bvd1r6qRPZXe
eljyKnxsAIkwGxB+B39uQyHV+a42H+vEUhD5qO3qLI8GRkdwYfRYR5ESmRnlebeRRWVQvmP7V0Yy
T+JxO6VXPhG+xi+4aM4soXlE4QmvZPMlSGfoZTXpyuiNwSdlFeh0bMT4BqNxhZWYFu5FQPQm8ttQ
b7NkCmtQT1CKuwdJQ/IPgEs+r4ugLB1daBMEtg6xaPhNeZFClZ3w85zlKpSDeCdLLgnGcL5Gzw58
2hqHxBhnfNabkZGOAv7igk1DHA3ejrcPRxMSDIJKXbVJ20+d6qmtNJXO4RXAV7FyB5Yia7afvz+z
644wAsDr3lAVHwY3buAByj15D8R2muazlFFqy856alWKWuwTIMPEd9ZjqOqh5DxgbppuDMt79NGx
b5+PG+lQx8oGf7fRBLCoX2ECI1szAXo4r8MSv3aw3r1x+W6qYz28lyBD+f88+pB2xIN/zAAKi2FG
rfbqpxJIfXdkinf/nv57E1zaItj9DhCZ0DMuggqZrQ2cHMLuiYgVVgFhkhtp3g6XMewXDJWHkmyI
0cUvbwTEgjsd/gnNDxID2i/zh9IN6NTTmpReaAJ3RhGMjP3RkGOkSzg4w13zwcncEXr7g81gMzrt
YhMnZPJ+QmnAL8Sb6RFnwL328pOLaUYrWvt6tEzeGZmhtQsQ815Jw7KkQa8pegmgpMX5rN/9tY6O
LHDJSqQgi0Aik9AgNVh3au6/3/j/8SHhLnZ4c3kvEEF2ralzjz+JDD86b4ZpMCX9fRQfnX9CrWna
8OeUkiIlmAsG4rA9GJqkShBNTdlUEz5FbxMMQrFKqSCyqwCGX/na92mOzAIjF8hdsx+RMt0RF2pm
nuhoBauBlVm6+CA17vciIjESZ5suJP/Y0RYbiykeT5P4yuBwK3PdNuagiH+J1pO0/jqJjWTpDezm
jGzsLGvonZ325jpSni6W/8o22cCAdmxtff9LSfhfTWKZo9YrQZxzQw7hMfnbnoiMcuPQgUwFJaWH
piMoZy3vfClwoN/XYSGua6UuWHxoIpY5k6OkyBiCKeUyrJPLMbVsJyqXqeKE12je0uE6WskqB37W
97OMvTUbSdorg1knjorhNNM4gWYLBCAFbluxYm501dZz/NbpGbW69T90e6kthkAiPOOzGlMqyYww
lf8vNRXm9cGZeegZr2Y7CofQt3rzRoad12ErSuN4zDQ7KwRxRxKThBKscX2g4S28pSdPLKrAcBvy
eZKa94skDxqvF6QTi+36AhkICqKr7loMoCqlntKvcuuTLeIK++eulJaCcSBA+plGw727LdmGCIFM
La+ZCHFhNLUvq1AXLmMEyPKJHKJoIGs5LlhmZ6th7Me/F93AD0jBm6j2aFN8hM11z4l4eerZbv78
QxfnF0sQ9e+j0dPnQvhLUkqvFJq4J8sLVxU5lj091hyGcH6Xl0rJqqruXV0/4i2wqosuZ2tOhQeo
nhLyhqJWV61ikdRPyQZDX3lXz/SQbBazwo1fkkLRTP2pLUIiqqG3HIOYw8JuMrkTaaBkY9AmPN/R
MLOSxgb8j+0/dwDzTLCjue4Nk4CSSF+ugD4C0aJutPNBBOgD5XkQekjnF9Gq1CY8YyjD80umI8gX
Ie0iKo+HIPOag9NfryE895NlSa+/8waYHD0jvr7s5gTlSYBuf0HhjpNPhdk11ISjHW0WeCvuGV8R
8Z9YvOs0JJCsVtajYUe4k02AzLVGF562tiiAuc4m8S9f43k/lkjeNP89uNMu52A0HGvmR64gJ91S
3n5DDtHREHA9VIdIpqSp9YL4XlhvGgLtlSqhG/JKKmzBHnm4yvKBfY6le99MEjUjZhaNuuNjnwwp
WOrqPGcWLL3EsMtsGH0n8M185Z6XYut+Ji8rz6pt2TVH8HOGuBBcBtJuEEeRjJsqYJrPR/IsaYqH
LWW7O50JFZVmh+B6eC7aDp9npm0D7oNPkvW5X45+whPy/v8xbfnYh336/efriDWbfQhgT2SzFlTV
ok4VIqnOWEHIyckjMX2Z0Rn88ueaMGKH85w16jmMhvSuXqFmvneZoaiQJlzrmOtxB6oX+Fx1+EHN
3KrnR4GRkszqRfuwA4DhvAFeqmZ0RytV6nx7LopRvOUBJL8PRMuIorPOuuzoYkarnhvqnODAOX/I
mQDttGQCxBEzT+TpBXQ/b/daXv4flQjWk6w5bDlLF1FSBsv3ehanzAbgWUKQtNp8WG99yG3/XS8g
x0aJilreG2CSbmXQHJpVxf9xaNcRsHfYvgG9e/C7OuZhcaelvMKfuoSMpEBuiL5B1JhSl+LwfsCr
DgdUY6xxEnt8spNSYy77vu3zXXtI3XRB0T0oZsZWlzpagJu83ol9orC1dW7Cacz1KqsB+dD2aEfc
gRCoJw2929HbSU7C1fOTZ9CoWPOoOEFPWi3HpCM+8sh1NH3vimo17LBa/PB9GANrFdCCcb+vJ7LZ
8/LWrRRMo2h33LRxv4AoVVo15Cw2S2BBWKTfh5TtHNSYsAzBu/z6x7d935yVv5CBBr2U9uq3OiDY
BHM8i+JaqLu8kkAwZi28tUznYD6OGzylxu4UHefVXHrIRUPWSdy/2/62ZRb3hyX1XnHvJSw5QmYp
TUfQduOUQ+Zph9/VOKFj0QRaHB6/RSc4VtLBK0c8tzKeO4YuQd6V59gTppXU1uBB1RloLFnkD/Zy
btrjtRuE7WIkhCNo/1dkN5Ntk6PePTP9PGfP8yvVYFllFbxRoekqR8DGdTBkjKfqsyrnJ0okRxfk
rwA8Gu7s+wa/N2i5tif8a4XRY/LAFxktz3MPd029+l6sDq6MsKlmy3m1UKjOPYEZuETRjW+FWMZ3
+8Spu+6g+4aYODh+EY76tDHDY/Tv1q58bEuMYSbhxlaTQC9Y3d/6W/O7t0aQ5AeWOVLow0AorKnj
lrw3iMw6cZPKA87d6jE6SaVeyRJdu3XKjSxRIkRubgPMZMl06kWE7F40/p/ceXUlQGpYKO15qeDO
aOjvlgyP7wPJnEpv+P5h9R37c9tRwuWtm3Ike/zmLa6Tt0iwZadKPfhd6K+cRseZTiHkNs4jatal
JBgWnEb4MpY3tbQt4LTcPyQnXNjdvuJuB3SkEqCVv5CcmoFEVHrUQhjyKqTWlFC9rMMLxrjci71x
sIPW5KfORPLgUAAN76rqovEkFAotjdUWamlQ6BlpEzSfkKAWKvekAAlMt5GZm4drQd99oHSX1khQ
UD6KKCnVUW1M+a0gqpig7TwsAXOUA0ud0kVPr1ARq/FhTFdbxxm25++HW20jjfUD9JRZ8XQlFcpA
mZ1YxG4UdWJyfQBo1+ztslhUMhw4OwvUfzyX7ARqTONUmS50HHL9OTstKfivyT5QtuCG/nmGyF3v
DAc9qy/DDSUalGF9RekQOPh12VH6q71DvF263LIKSdMGJn5RtaWbDt+Ss0Q/WicQia0vGevbIXbZ
YIsxBlrkaXJZUx1iKeMI3YA+TeBt2ZuSI5elqy5h9eBKcCEWuo3g81VDo8HnOot/nT/pnoBHvciU
9JzUG290W4EmNbEavs3E+DJvF77odzpB2ZprNRPonydUcqz9XTiy7aaZx1hZIOXZD4hvDAs8m9qQ
UoWwerhq6EV98TeEwCPGGcKkkTiRCqf2ZZXDAVpqx7Ii5mv7EoFRgoiZBxljXOAx0HleueB3awWg
EkNA65PsJwBuADCnT9rW/x9M7JTNsFm7GZEnyMzf4Lg6514F7jZxzVMsYFp0SxsuVez5RfhY7gc8
2JrfppSzZe44i6oWtqES4/Rw6P1c7fGXwivVftrpSzL2qioPffYv4f5rP+CYT/eSUBsYJBJfYkR0
pdV8s9mxsSV7pyVFX1Ino26DR4uuxTJnvR0GVZE1fBQYCXE+PcccDlq/RU8ls0a9cHMmyufYWUf1
/itx4wFJpVezN5awFQFlRKxVA4D3QcDEOcCRkYvuNyQISfQretzE8/lUkzF0BEYUchqrnQ2U9pu8
VvsHc2ECioPpVvUq0bBpk9TuB8afrS93MybcqJqjXg//+fmtiKFkzRPANGkUim1Z8tzgLlO90EC7
j1j6FmTK7f/8DQmkkDf0KjukRTYqHlUydJ0Vdw3AJN2RX27UyqsRBqblLqlad8BmjE7fqb2eaO/z
Yl0nM22tp9IEyVaJ30taA5DY9IE/evSBkVLmo5VpNUoGXH81dNg7WOaaxF/7o+zMGfgoch072YjV
TlV8VFlKzYEeiNxiBgA1Q3lVd9EC0mc56UlyVLSTjNLLgQuETKJNh/4aBJh1a9n93CjUjuz65jOa
CKfxiiuJE6EsGA1HySqfVXhwDjLl+JtI9sxc4RDyukOXlPNoKHxPXMGp/draMcBJMmOiLFTmKPzk
LBjEXhtL0F5HkPtlFHThsbQdXE+tK/KW//3zwgeWtA90toQCJ9GKchm1PiAbMhmzNsfDj8K7rsW6
KCYJBSqd6av+knoq6lLGPfVe9yfdUoNTmgt6mInCI1H7kN68WDY367J+CncNDVi7Wy1KNRILyoMW
2kX6gT9dHLNO8BRbuNH4KbJbSzmGDpUiEsG2Xnf/A6WnJq6wMKAMWNevgjjo18+7GnUxPjnxbC1m
xtFuo7EKRHCZRTwY4Qk61VDrQ5EctmkpTLgxmhs98ftoZvYiLQd1CWuNPQ5LsnVS4wuv79xx8IAX
0Esle9+WQSLk8NQ8DZQmbkQAdcQIo7epgByvelML/F5jTLP7xvjYMF2ePOCRADX4bi2ff5h4YSbA
Jfi10tQSOWclsJpAZ2yqh07GGtQGA74mkbLjhc5V53fL8n4wT2aZfEYqO1kfUrNMuXPCS9hash4A
GtJMg2SYls6oGme6N4UQccqMUR9pTmvhN8nBI7kl6YfkMfRsU6/Pux9NIGQ6DvAZ/OT7M+jDS6p0
/1t3Lwv5IHmQ2G3QoK38Y5ooxjvczxb97C6mmQ6I9GDEb7A6H15ZpaUuKWGqetbK5ogBcWazGu7k
s8SNIfco92JYYglMrtORB8DDCzV+uYp8+DJNjPZUvajF2xdqPPJOQ5GooRRTU7WvSBU5LiM9bDHB
BvxgKxv9zW+FaN0AAOXsWj+0A85bp59VS3CyBTjz7+g921Gbs2FhhtMdNdju0rzF2m+lwSMcI1vy
nwv9BvqMUQTytwootij9zv2AqWLiGyNaBviuc8PpI6W04bFexbOWBpKyWzFnk1wd4XBm9ytreVHm
dgveRyj2qQcLAnLHzaoY+tBqSnPMm5Hs8vJcVtppN0ueQ+Zyq0bdHqqyqIfhcnVrapdfMe7FAuDc
D/hWTPtmF/rBf2X1MiC3kOSiYGr5b0YneYP51FN17OQaxyf8GkrUFi2q5QPw7tbT/FQewFDdGcww
5kqJKNvkwxi7OeMcg4Br7aQDdiPKsTW6Uhw/mEYCW4VW2+qDsC7+W9oee7Oz/flTejl6kZqJHcKZ
oZ+orslvLA77aM6d1kYFP+WEtsxV3yzVqYCKP8xpVGf2wVFZJyBL1px/+JpciDrgly6PpgZN/jDh
gEZXHSaGl6LXobf27HlJymo+D1juF5yNx7X1iSZDNY1croDVaIvWcPvnT8o/ZF0AYN3veWCWkWxU
9/KokQxMBbYmqtFbja+knP37RDQ3m+npidlqH//Kw3goNBW7qN3mnARa7T4WvTSq3XT2B566EOA4
7CBoJwAoOOtkfb+kZ66Dm9NVsthMyoUsobgSRZwI/sYdqB4iEC3B3CZXw3RiuaWdVYKClbocxDdn
SxDWapTWOGDRVIT0A76XC3ICE8UFqudag8q/18M1RS4vs554G5JEyDUrETl7CRWYPNz5hFkayZq5
zgG6p9F6HQmHNuJ9bzLqnBB5oYIUBT+ykTZt51dIqBZG6A1fZT85rzbxhW2wvaxMzBf/E/YRakJv
t06ytKWOzyaK6ndV4D1TdwOT85dw9AfPGOp4d7+sUf7KZl6gOO5+2dQ/fzemsjp3qUN4j7ke6/zx
UY5yyxDS/l6Lym64jkQP/3WKnSVfWZngka2X5yj4o38mkIIMGs+jGLdKTgiNliB1tsmSItYQM3E0
GhZXQzM7NcTjliKd+EeUMjeszxrG/p6x6EfGtfVthkzaQH9fGoYeSEZ2Cx1oisgw7NbRPYgeP58L
diiwPvDMLqBLMQJxvZMKCvgifkLfnt887Eu7LDqqBObWgNyNp2lraMSoYnNnf9Zp3/ImvjLJBx06
m+8LHrS8zQOgxnipI7RdGRTWrG6W3IYPoONOFPXIvvDSXb6BpNtCtanYkBYPnB7KhTEzBWzAtHc6
GhH6AGRo0viWhmkd/AeNP7Y8NTVW2jscu5ikoThK9zIFgUh3n4I0Z7QN4Ye++9ctTVgWyPVVEW+V
cbgsrdfeYTfJyi4kULBXNgGkZGfEbFtPvNTxknEA7afkTrlOyWesECMiJ0PvGQpedf+TezQkOr99
EyhDwdIUjFEoGYP7f/BBXM6T7PVrRrCB8PyQHJNgj8PCkOws/3Oq+YHO122ACEfpLR5uzqgqkaIz
QPkMez5Upu1zmlVzPpeaDizMjIOVm26b1A5JFGyT+XaNSCdfJ6almnjJCdKVAZhwqgA7wAM4BPWf
eKdHwzqgvEKhgGJrW2AYf1BmedAA2UrnorLvn2jzKjhedQWZHjan1M+SMV46DpnHvpzDnSmfIWPM
WpyoieOhKCEDpYO8unraKZB9lYV1HJHN51JD8XgIvgOBKlYLefghbe8Fe9xHFwyMo739M9yW14Wt
0UflxSuLZi4pm9oBCULR+5vR5WKJKaZUMqhBSMKv6IOAokQURujocoVQNR14gNF/rAPHBkYmcpZb
uHCjaWF9/piZ54lqwDUMAyipeSl0eBgmgyFnt2XBgT2S73DHSWina3RQ1W0G5mC8tb3svfNNX4i3
aVhvgreNE8qstBme4ZrtNOYqfuuIyfV5AYbw74vILr3/Cl0okqL2F1cuuSoZOSstDBL2Be9NPg9F
yuuYKAlEfPB1PsrgAgQmlTmMBht87dz7by8RVXNrf7F9KpILPx+ALCX2bNXH35ZC0cAouAayvmBi
vMM3VWaik/GKNu/yigBrsHfNYsqhNX/sXYtajoLXLbk2sjX0zB1JgVN4L0yoiVK94EAYmMmf0+5u
UsfaZ9mwx0sDutP2tAHw4/8LaK3Rp99Ri0+WwEuufrTzLvEaIlifB/PTkaxD2Vx2nhtHNKW06TGq
IYdcgtmgcrJlswnwoefZlcQhFwmOhvxxcGh5GIv+pmRx2zWrbkB5iOqqa1OlFIPYL5U6nUVWaMON
i4Kb0G6bgvH6ltabjH9w4Jt51UQxwv/IiejDTPxFBNlqlqaV3Mt+M+DPCixJvTW/Kie2Rm0QG4l+
q97ucyJsv0VmhYsnDutbVd/U02mwwIaJwlZh8gBOyiB6GTgJAE6z3oRZDNnm1qSssrX2cKzp6M7U
17g7yMGYwNb6Anz8ejKgaMqDhaf16lZL4bSTh8YxFRpbx/yir2PzMTOUe5oZ5PFPLGZPr63HO7V4
w7xSqUZid5GmqHZeCz00elX4+2NGY2jt4xtEY6PJxa/iOMJ35E6fSM6mwRqZ/fywy5spm+Yyt42g
kCYQomcgDkx+0t38vW0pP15VVigKyAlT7eI+othY1mZR4lxFs9NELwEpQM/eALbq+GRBvzwpNb8I
4snQ3kPZZkYjs4TdglRj+GgAGqNBde7e1TSoiyURBbXQIW+ZsJwzIgsbABRDp9rk/RFDaL6zOQWV
BePLmJBbbGXkukzGm0XA4EUO4ZweC20eKs84o5kxzTlqfqhJ9Xq7p/esqS+4yIV9dRAHzKJ0nAMa
3IZlHoQIwPrT4N9IzJr9MM0rPcqf1+rhU6276eQN3ZIgVBWbsXCO4Jf+d6LEcveo04txfxEsfMhb
DgC8yZF/A7L3KRMSpGPtTgAxFkuT2KpRIHwi73BND5CZoJy9D1mnZAmG8AW8RUcrGWDDPPYe7c25
nrCTVw/5FdsqlgsKt9e70w6BiWUEywqqCAgy2+bXWcXdgxV38pRR9EogLzmrv34cnBrHZgEpxuAM
wIAegxeSPqnTecNO2suVo0t0tZpSmActkw85KPYQAm/Cq/wKFKp1bcltxn7s3hskfTmqeADkkQnH
HaH7cqgrNHB/XJUHayxVYWR8RsIUmVu5nvlfZ1Npk0a8kjnSWuuevcxR4vVusawpKnhcRsB/QI2B
9PZjWrppmtmFpe3+6kWxtKXkBb1BDlUERA1C4ocnwXFP5QKcVRFLWyg4YEzYJ6L7j+fkN+nOVuzJ
r/r+OO2xXuPEaeplgfjML5RFYB55RACUzomNM9owurm9H85m3E5Np3wghsLM17U688GxpdAtfvBI
dUc+mqxT4WjhG6rondYM5diQi6EDMgu8vRToD+YeAPX/iQ8neI5/ncUQZPPWlGPeT0LuZax1tGT2
yOc5LBjf/6/FIwc1qNuWPG955MjoUPkalOjBHhlLwe92ZQV65uR3JywxlW1/S4wowvpcsXJ2iJlN
yOeslqUPIs09GNFVNacyqr8VXbxLK1aneeF9yImdjSPcAwAs9g1zX7aZ0eOqaziWS6yC8GjTtgRG
OrXnanqeTVDCBCbHWnjlYYfT9nJYjXwbXEuUDkkLUhnWuoOGYj2YUklbNStXxX90PD/lxhBq1bs4
dViJta6XGv6I9ZzxwwlZ1PvYBWC8pM6U5gt4exymV/cxU5vwruSxzSW08H7pPrf8B/IFlr4YJjWe
+PU6Sn6cAaXXCpLexrIozsuKR5yJ5U2rwBxabY7bexFZX5wWtJ7RQrx5fCPKdgU0wQJwNH4nYk8S
Cy58E2jST95IXWdWhTjbwASVKgZ82b9IPsPEUYWHUV9u/SGQposcmkmfSu7nG30FnvpQnVO+oxdU
B32erSR6trLF5L4P8HQ1ROFMo/G1bAbzQPkvS6nSSC5Ey2ZP6kE0/bEYpaN6NnRhA5/ruhaM6Jnz
6aWN0LqiYNH6ZBNm40NZQARla1eqJTf8LM2H2/lLbh/vbrnADb9JibOwgM10HfEuc5ZwENI5Gl0b
ihZXlfueRHrpJhDuvI0y7Sc9I82+c5CAsC8MgSgXol8dynCwna5C2vII2gKaGlxzwztqfKXhan+Q
zQVpfFlqNhCDS0kTWK8j5nEk8tonhQ+12F8ZdRWCIYZU/aWaCL8AKKmujYr4RnO9tvf0gk/7Hc2y
MK0xmX0bdtcKOYKWHUMXoyyX4rbw391nQ03k6400UxK0cC3Pz4TaT7zwe2IExhzq7fcCWgBfqu3p
CRkQBAMp+C8W0HTH8Shug0NKzYPnE1RDXP/7xbTMTCP27Rjml1eIu+bW+EGd0kEq7JSXOzUzlnvo
5dP3Oxi8LQnsRcP51k1TOUO8KbSO1iNl4Xm9fue13Op6KG5xvz0dVB25JBevMkuOwXK7wntiE9Ir
+Astvj+JZGxu5rFYiGVPiRTp1uDhNNJfhl8f1gmdA4sh8V6WfphXNMGc3QkFSvER3nur1VXuWzzW
D4xlOyBA66QPTfs/apbZO4SRJxXTjey4camjFLG91TZlAhi6X9W8OOIM76VHBDaMJXbFsPXTtnm4
WRMpyTndUcjSih0ncZZ+28pwprZMecKJ4cdD+fJQ7ac5/s35j0KckE5gyNrk2cy99BkXfoV+nKvB
bQsgFctAABvSqLBAI8PgRwu4uUmTNaDj7JsWNCCBruqjtdy8jr2AXjYPhq/f7j6gQmSHVLSZ2457
CN4o7GvWl1ikqSOQ7I25yv03wiZkqArlJqSq6iYjQDICfMTIjzy29oM5eT6AQ9aXxtto85TQ8zm5
+iGT5bnWF92sN2rvjfVJBj6Dly7q4KV/rqpcpbojQSmhV38J0/Iqjz+pu5BIitCCTAzgMNrAeq9n
xyXNIysjOF0+tJOQ4xIEaiPI6lCO0BJJCjv+x9ruLaCqlaUIGHuRr3EJg4IxLnZ06L+Lz+m66pEI
s3iLveN0LLifZJi6ac8WrTlw+cFAoAbXRiSMwMjWrtlZNISEFezMcT028vYFfgSAKqqV4m5gfsKL
D3YXbm8l0wV7Q/En37EEb/hWH57IVPgl7GwsJxSafMzS+DLTcgI35ypIIlIxJHiW08GuSXZGoo5t
oz3ckB0TRE9hm0jTIFADaAXnj/4ZB7v97YjPjZ9v4NUZmqL8EtSDPrCzMdubOTmwcy1hXV0iZAO7
+KIOpuXv1fjBvyGLLqwO6F4tUsm16dobBoYMMCNsJkH3ctPAtWOt1cPk40oP1iix/19B8DJTTcGq
tLsbkeGgBqwEDbjZwj7UHQjAbKwJmIT5RCUgNWBXSnzfYmsEzoDsszri6wC5BhR8xPB40PykAAjJ
XgGY2xtIlahZdNVZjupK0t+y0z7OEYhQICPRiky0FAVYJjNxwumvTbfiKRWLax6riC/91qLPTVac
MvjQu0RGo3/K5qrlWgpC9UwJdf6JkQogWjuDlacCOR/9PCQiuMneEJhRD1ZBNNcHrlrE3TQyfiIY
i+OlHCxtbgXZAVLZiS2FpC6lQVBkFFzb9jPhcdeARZWOGV/cnK8kWPtSrPtoaT+hj2qgIxx4bNxr
YzVEre93V+cQdalI1CDHgB+sTQ+YLRZ4CcZOnoVQGqrZuacGCI8tYEHN5J9+E8gRNA2GdMK9VNs8
JJjvFGH95wb1ArBJIIm6SNyDV3zm/cVqyOBk2KDICcs9qBQwH/hWPdbSHbTiTGfwjZzWIaxq8qOq
RQgyIWJukmRQBre5qvvojamAzYCboIZwkAYsmDLpIxj4UBHNJ1enkbgE12uT13mOJb49HVoiDb5g
3pCOk7JWckuAwkftuJ5UvT1wYKBGQT8vCkQdFFnb92h8bnSOIexwgyEkMFMsnn8Lmh9mzv+Q6XxE
1vSN28rB/C09OcKgwKFj0sSs5jBahlZ/P+BN1y04CKE2it8IibZPlU6RtF5xHMn3Xu7afY/aiujK
C+tAre+IWoePfU6b+4/IdS6UGP5qBmehVrkl74WxsYNUiNIRvBrx76CjgLLo2X6T8H/s6mS+OtrI
9EbVdj08Mnw+7/lRNvPBkksBY9dz2EY+fcOKjL0FQs9XOXhDdfbV4+l/kHwafqDL6MgJYns9vld/
9Yx8E81OCyphfffZXHQTDzc8hc7XP0vHTWOYRl9L6bEioLrdF8pH6ONPlnDHRvQ15C0DajAwScIg
N3nBIyqT1uqXhH3w8K5wuxcuTQyaKqCehRsj0fcbQMyQYztuz45qbgHj9AEGpgsUD+hqh1wrl0UC
JPd5X+gSlEkpU+bP7e0AsCJVaMVRZdJQdSLPPNgZeNQUkftvy8YTiK2U3nZkEmMt728W8AHMGXUz
kCHLVS8phel9j4hbBzdemvlL1VCbZmN2JSCImkaThw01Kt4H2XYGh7ktll8cz5irSc5Kt9hptMpD
QN5hfF4YGcjvjURvIS+gbjR8Kx9ODQecIWy7NdM8goiC9qEOAw1gAmexrvOiRLDGsYSpP1ZYTQIE
1hDtK1M/bW7Mt+iA5aOQrA2Evxmp/MUXmBv3UleGGiRHHq+yYTlz1c4t2RpxS6N+x6B5tIxt4H2K
ryUHeEyT0vhmRmCgNeKBl3Zbuxfq3Idtt27TLs2ID0NjmpXtqqUSUP9IP88vvYiLAmDOfeN437/7
atcmi4NYI87HTANrfHwxSrAADqLykbGXx1MNshFgKscoq6U8cHkS0NcxkW8EH4ZR80fmVCu5LCLa
3wbe/OYKrSgtbnChgQm9Bsi0fGpYKBJ/JKcx7nFH1qIUudGFBAzygm03xd5zBe1zAo/F2oaWoec3
igI/rChkVW+cVn0n4k4ha6vWKRGSvkUpqNEkW0o3UoMrYO+/bTV8zPc5uycoxTDPxh6OepWPjcPr
hBhLpSMR7S97jsRIInZ/WJ3W6mnUKffffCqiWmphfUv3QU9dDtBVid1Y7bmHcuZwKdROA1JipqFW
TfS9JouAGSCzmfhI2JFA6Hj4UjGxAsVMX45rk60xA++P2IbNIcTpUFM1vWf5JECrAhqiG31N59WR
q+C+I+YsOnnYDJaP4tcX3VP9+mT0z7Ibb07NIKyk92UHKnhuO+MVPCeFNdF9C/rgPDAdbVizHwS+
mD6XH1S68Xsw4lYBO5/Gc+onuSaUa0xFOWGo3aEmPvoDppEENR6HqVIh+2DnST/5VEwiEpn0dpuJ
t2ue8hdVE2kdoIvXpChODd2YQ3c8HZw1ft0otCVIrF14ln9Eu88AHD4ULl5UBEMlVxlToOf1f/8z
s4uC0ve1b8yDYYcg6GmoJJiwKk0D4AugfeoaE7KY3vwF3i5J5E2KsfDaE9k5IMN1q+PFF0r412oo
gjcsrLm6ZXiRH7hpxxiJNYmhrOYg7j7p9oVbRfUcIOnLFzLWwWASRolhueR2Ar7EsmD+OSDKDDwO
vO443YRT/N/JE+gCTIDG/P8TRNC6AP4ZyTk/IiGTrQzkZ8mtqYYVqDtlnwePyYvAw/RdO6P+WhXE
csGoiAaP3FtDDzPtO4u72A7c9B7tEq/+9wWdOHCVtR9KPlzJIzH9M3+WKDElzY4o/I9nmSnHtdy0
PkFTAUtCqj9MIx1IbRreuJLPTNZXHS1uxJsS/zg2du3uR4Glx6aS44iRuFdNnI+16nmerhrG7bfR
6XbcL/kh/cjW7pLt0MqETmlDHqip8ypYgLGOq2Aoin+M4RF7I0DHVo15jWTYBJo+0gd1JgYBqb00
emL9xS8nGdLwY1C9pGSnk6AyabCHDcEMnY7r4d3BxU5xaQbxy+gqFFaNWMmYTgBh10O+7GJ0eQvA
AopF6MK/+ZLCbI0K6tO4WM6ScduGO9AbQbrPeIK1Y2dRgz/swPDMXEZSoP3qXowqmDnyUNwnJfNY
Jl7P8RdXme+jJnyZ3JxNZpa5zT+rcCE66/Edd8k7xyCAtEPB8bNR/cLOd/mIqp5SrslNl3rYxjbs
sNQWzzvQhNmUywDix4yfP2ea0wyIHgYHvbd1g9+pqeCBDAf7HLV83N6OWtRN686E3OS1c6A2k8Rc
kKyB56IJ0usOB7l4cQWXVcjpfJk5/CK413aqK2bLFkwbOXHI/iViEtrOni56O1e6yjqy5V39mQYF
2PydgmahNFTdaOdB4VTjlHiSU6u7r4+bEQFBrrhgGuTQsYv2Nl2C8GotO6z2IVQ7r8cKPZD6krEK
MSlMIpB3eh9kh+ZnDsGiOxdFGJj04apteaamHq4ZAYFJJMf6oFXSef5Hywq7WH+RrkaRFXUHWp65
tgVaZ+ZM0dHVBHhfkdoRpJ6ZPxvwDsdVf/qJWla1viRM7k2KOK3wNPNucmy6L7f0gA3YYJtf5DID
YkGdSkXpkL7GA2XBWi/ZZYdfHIQDCG1tjujIrWRUZO0Av+4VFKmA/CgvyEa6KQAzCvRZi+CwXutU
jPm6V5cJeMZg/hhGwEhf4Xhj4pscenbeca4gUPYd38nuRC7n1N0HP3c6TjiBgPWFte9QlgAcozLs
3SE0FNam8VEwdnbmTCSXwFyjygOlFXHnmBFnmckQ5sEyitNrvn/09GjpLCuZuK0sR6jc5F9+VB0z
WdlBvfXrETMoCAQCJ7+gUER7y+zSAOQyYPUMkNZ0ukG/zt0FOKs65vmEpgmu5Pbgxmef+OtZr08s
qJ3rIGQtCScCVeTWfapx/tggJDGJcNVRnN95zTtTIifhpSRKJLyUUH2pVEJIHIejwZ8Fk8ben0j1
QOlo6dfhVG7c3OGScbQx7Yz+WX+HUJZxMf+v4ELn3edBFRRQFYDs0BqIH0fFu8f2roc1jcn3L6ss
mEem+yUqt5Jd+1LJf1yvfIjGsMzQne52JBkuDdPimfWi55c3p1aM3C6Gqz8B4ym2bqBhF6pBVHde
HNHW+fI1AUb91q0TzvGixJQc6sQNZ/jkpBhyl9ASvop7ve22vlBp0l2xVyVtqeJDJeBjWx8iKAwy
f9j/No3uJ4cGnlJIzgcH+zgMfy9qIVTQ8h8p7b8Y0e8VRKzO2vNSlo4XyDAp1eh1m7RalaNpnnis
mnjp1Tz2dkj2U3JkcYRo8ynO20zyFDDRCOeqs0ZvzcYD60r4YjYhh4sh+RuwkFJk5Achly/gj6qs
4yuZCr29ORnbt14jbEEFGM1z2OUTAP5T+3ptBc1WEAuPXOohHfN4u7Q8j7FgtAzI0SVSUcBEOjKL
oMBric5JeJw071OkHGVW2ohl9Oawz7beKL6N3dpttfu8iWYNqWccs5LTn6RYt2BEwGwz7bIARNz/
Z6wq7iF2gm5Y2NuoYlHFCWEK7DGgkYmUQxV8qYzjpwDc1Iv0WdejVHPdoDTo+4G90tWErZmLPd51
oo+FL3P9m0okFSzOZsLwqg8CC3zO2So0/57I4SJBY2RzOPtGK75RgMyJBuyKxkTsDdI72Gndsvdx
UkJCinuQNI4Jm/LFGe33WrjMphijgOluV8WpRL4uHMMH0Sk8wh/IKjlRdV5aUch9QsJH6Dm3XpSQ
Oe/JpxuotyIG3SiH9T0LDFOr2Q9OU3qEcDSEIjZB1Ud7g95+EYvtbNUyQPU4UtTd5g69yTB3Wnk3
unnWvCjfmTEl3cHP+vtB2nLi39WwGO0tB4TnpyNpZI3CUkT2GINohBDtXSAdtBCGPHct7SKcEm5X
m0dGcLSqYOfzpPyS0Wi+p6MalGQPFC5iX8tbMTpIR6ITqhdeM5rcV96b4OkbwJF+PJUnIkCE91dk
eZgdBogqXzYB4NthxWg9re2gV7UdxR1RFmK3ZJBThq1PTe2O8dz08FJ9QkzcGDO9MEDVAVlRdUdD
sU55bME6omd9mQrcWinQOmGz0ZHwMvlwIjoed9o9mJZkS+DuSpwXDKtAYnXUmgTJzrj7oNErxJ9m
JuzYveVVDEpe9rC5H4oXTh1L2+deDThAN4fvbu9ccZ9XlhduzrQknATH5z8Btf9AA+9VnE9HLj1a
WyGwEt+VAnk8Y2ZoF4QfEa+apW/OrqLgbIEUPT0rp3ydpHw4naNwxdNtIYqTHFZ1OrdorhqXcCS4
nVmIr9lJpYUFj2CCFRKHSLGSU4jwDG47FbvZzSF/3ueuPbjRhoRmFPyETnX6p6oxDn92S/bw/Inr
pXFjlxPK57bg9hEEMzRPcHr8jrs6+2a9fmXE88t3MPcqsW1S31Z4/pFt7My28AN+YygEJi27s5IR
hscUWXHJS1bNKh7lO5Vt8Lmtu1jTTw7qf9TdZlh6kLK4A1tIRsAGcEptSZcc63ta917E2PRPCJ2W
UPRbhD3gA+shoeIXh8Gz3VnBo324lge9ny0AOCFkqxAD9fy8UV9AbQ2k7altMwK7g3augQNlbvng
sRuH00YkAVHwOnqq9ODOckOXdIPcOw2x2cs/6uJyY74T1htwQQ0tZPQeef2c0oGyG81XPqHUFfE4
5NVeI4+PlI/Rb5R3pRhtYNqeHBKzkJlUZnNp8qXv1eUwDHaIQTGSAUu1dIvLiMXiqAuvPEahUW05
POSXVgwwltrAu2vwVCXK6i9NblRmyObazOfEqnnvG5qGvF2o8zlSXt0BWVH4dAfzlS5RpNdsFzFT
ssTAId+czUF8XtE0HcKdOCbcGZhsqsYVmo+t1k3N1bgmlKNSex62oNt6HYrVUQ3DyHADK3EevsOx
HT4VdHIP13PA1Ve5ttV0mdqm+QtEcF61fmWyteSP7QQt6QnE+oE8hs09fLJJhABpRdJaitdn4/2I
uh9EZEkgB+rybCoKGjokdpR/1ibZo8ssV9BZuPgNcoYflV9juAT4SC/5cxW9LqZwtllO+U8ylCwk
s4nZ8Fywqkdhwi7uh/GIOGwPbMvouR4rm2v8Gz8plrw9lAlt2posSHUxX1FOdWU/FRJmgMgSFQLC
oxInbCZMJBNIjXfpWo371cT3nx8Js/kVWr9yTXW702WU6Wq4yuxjTlM/G9XgMNysj+bAGznEcTkd
r7n8KxqA/9EijG6yqafyIAXPsZux2sUE/9wf0s+zMmmBXZX4rqaP8v/v3p2irVpdX4VpLRXFc+kR
iGVjc/eSc2rQVYo3SOQRA8koE3ZkfTKyfuG0nALgTzh2uaXk+cNeNIwJ5GozWWBBqKGSpyS6mmMw
Iy4cVV5/QL+0oqaWr8w698xh6/N+/WIXswAUSNPHcBBpMFCs1i1elEXHWJCqqznxdL5fljv6mdik
4KeVKovkpOaxiebHr8/F5F50OYPyz4cxGiqXEjktzTidN9d1qre5RK590XPaWIh04wpiGStgIY7l
rRODj5VlWW6dIAMzMIGMcLDMFROmS7yykKigJKqhcFOf7b4P2Hv7yaBKpZXFfbfA3KQKtSrD8Cg5
UUMkgkezvXEIpxEhz+FVMd/nwHXXni4H9yzt6LdhG50qGsKSWeHKy0EU8l8u1KBpA5FHJs17sXYn
lotlD+PWriAtXqz2CqusChJBZxWToSRgj9dduTP3A8EuA6tPLgeWM4yTlHXUyAp8iTLDhLEs1nPk
prK++k0aociYBda98e1vU9PKh2yyUU4XI2x9+/40rwu7wG7eLjuaCPF/uZn1/yBPaotFsEdqn6X0
Myn0RCmKsLOXELl4E/2bSimZ7nCJJxwK3Z/9fLV7qg+T1Ilcf2lpXxpUy1JgcxVmdo/G7a28wL6Q
k/PVmGV1kiGeFrO5pwe64vaCgkfhBg6v+OBB0V4TBenY3RDvW2fvyB12rql8prhBdqVUO7P3KOp/
Ze61UwZCJux5tarZWIo8mkO3ztxb5UuVNMfgvdR5f6JOTIGL8BDq7d3bLBY9OINofj8PUnXPZwr1
pLguplrb3g9k+v6/gGb1g/BryjlqiAmjIvUW736YBJaCCWkKpGUKZeF0ucPWa+WL3P+NmYWOC2GP
SKEwftMOEmHksbbT4n26xzunvAtK74BA3V6I+Hf5ytDon3iB8MZS7EDLycypTNO/K68ik02gBpYq
a509b6T4/srVTch3hl2FEKFjc6vH6J9RMCf65AbOb7bPVtNKr65+QuBLXEChH5caWFKaQ883ccML
nZwcy69QH/C2mCYEvOYKMntezuz2uOWt30TUf1wjDxPqO11CB/2Ii7EP/0aQKFor+LQOnqDgv4aj
KShqf9xg16zhapNv0XrkG3p79jlEbB/fi/gFCNeck5fUjyOiCkxn0euDTK8RI7HS/Zj0VUPAc5Bn
oaQx5X8Ut+CjvPQPefTtTK8uyuZdKZgc7i+PT3wsYDDbV/53sZXcSQ8AJp2TsLl0m+r9MRYedAwT
rekyBkvkOABiydhfyypMLswIGg57cns6CAM5QNHfehNWWxcrKscve65YzpYGZxT1nQ9osJ8pycmi
INJSi2t+Uy/tfFNoXsvWoz8rBUf1C85R8KOqrs9PCbCqcDFpKKRgdrYwvC/W9Etpv0Ze7/hT/0L3
Pc6kH0xnYJIy+0QDn75zUxgLMDYodXDNyFnS60jEo3xQ7CRUZ90/ZXmve/2hK0NdKBMcLWQ4HKLY
7Tl5H10vVYdscKyoOVb/LOA18eLJxwJg7aYS0nqgQXp4RgryOTdt20Cs2FDdM6GK6mURyaW+Ab7D
msxhMzO6yTjy0XhG4zTR61pLPkXl7uyroJNohOKnYrjGbf4XCTFg3hutM3O7Z/d0d/LmgHbzXPM3
PmMyfIiw6GUymzstFc9QWqxaAPF8S7qnWi9RPMpa0ITKrfmyDKAsQfZo2Qs5mToJuLVOEDG3rcxD
brWLRjkBbM53RlHNeL0KBaM+dhvsAjTQGWjdeIUSvOaUsMHEmQvt2j4bYME1nvQygh9VZ++21uyN
BnywQ94mMUE1p2KqnQRBta61G4MmjSFMFNOGD5F5gsgUiovJ/3ba60503FI4u/Ms2MC4YATh6dky
nVL2unpw3UPoFnWxgIUID/ySH7o6aVvrKggKf93LRk5BBnJOwFDQs9pSOP6DUFhvEC2eYeCQkTnA
1nbUvQn7XYLsnbkOULe84PKQ1Scpf77SptkhKm0eNi8T+42hmKce4R/hqiEHMl9A8uZbampa5+Av
MQS9EXNokpMGl5FU6M0YySXfSI07Ng8Elmb1Bxf2LN8OPWQsYOUXAN6D+chA0VZ9OHyGPn5Xp6Qe
zrVvnHeRnxtcRWU4axv/89rTeKk+LZg9kCfat/K0fQ02/X/vvCS5fhIJ9Dm8YrVJ+9kCEBUEmWlb
ERy+HS2wEszbcWS1X4H7UqA0SmY6mLKHylz2/u2N/PtHSZNn435Tep6nQoCsc4Q68BUd4nonpHll
tL2bHcOEK1TOEFnc9wX3ImMyQ+ascTYSxGNH2fv48lq2f0rm8U7gbSKJthEscFBEr19TBJ23Ct7m
4Ke0eJZ83SzvPkW9gWY6cVuwyAGDlXAvSx3Uz/HmI4YW9sL2nSAaspEaleGoAJVfaUVJxT8RirzN
0j8QYbZs80XQxlYSkaXyVIbMNyERwLAREvQfcGIC/x7lJVPDvMRAoqRAgBRNu9yDVdvz8/tr/Fz5
EbdmEOJjxGgt9N1QhSjVtdevBa8WmcXJLtRtDyZbyTTpIY2EdM4aCyjzSvp4u05OYy30y6eS91uN
XAoMAbxzWMPXzqS6qN7f0sbM/3o8hH/Yl/YTrba1ZC3rJfOmLKZ+gFlADOtCktiVlD4VsijPeguq
MDiWzXqDa9a5RcW75CelKkFEtVxcpeygJNcjYackaH1f6OC0HYJfEJRU14gCFYd0/HKwlaFCTFt7
ICWPOB1VzGO4gbGur+Q64I+B/r1CbNza44agJGtw7TL0Z3QIUbuBKyubKGW8aiyxVCvLjs8QKBUy
Yklstu8Eq7Nf2dNHp0f6VSX6JCuX3c7b/tnruWAMEyb8E45Pb2/9/PFnb543ueA4HibNmagO5vNq
QAzB+vv2Kkwvu7t+E75dnrzuiaD1qwAv+MM5o/PfsPriCEwoJEznbuamY3QZS2jgwQ+RIut6vl1+
6VzydI6eF54OXi8+G2EaYWmNoBZ/tdKrrqzLzJhW6EgAwX3wAf6vdUCO/lGHxjogJ/FF8YRMZsa/
IcIehAr0My2cmoalAtNW7ymLkzha95ojZ2GQbGdhTyPRMEC0NVW86jKQLuTcbdwVOfN5OZMx9UVA
QQtjEuQDm/xzm5j1G5X4kyEDnLLaerrHlph93Ak79BRWVKViMSKKH8rsNB6ZrRjVDOm+G5fI86pA
bu898Yq6nU7ThM0fvTSOpTRo3XmMXLaezTG4dZBlTpJX01G4ZQbYhsCfWJU1F3dGcTfPYioLSEL/
VYi1PvROi/6WF0nTlLY91JftSxqcq1c8DnGKO/08gyVbMy+aFtUrQAk+n8GnAKKBGzfUuY7ZPCoq
fso+Ft0EFckrB5DwXjIIKkbVlt+5uj+xyGEvKR9IGkffBmKLXwAXtnrG9nISlv12mRezNW5GUx7A
2PMq1jiHBY+xtrJzGRAkt9yboGJOfCltLI0Kw7UzC5PAR/Npu3YthkIP89pyQ68V7VVNpzYsJAqC
vpHWi7s5sb9L/Pyy7CRCCs/usV2bymTUd4RiYisifI9qx3YZ90Fi52X6QFU6yJVgzhF3ohxbpkDN
WQAWJZo6rz+fonSKH7sdYjb7j6lmgnMs8/66lO8lZ+WKAPogoWnben37c8sczwkCjNpGoeUV0noT
9KaR8ceeP5bKyKH717UP8l5kdfZ+aA1ZG4Tfz+wFBRXJpCBCt5db+RvLapiKFapONCHVbD4/P1Zg
+iDN5iB1nQdNW5NA6Dfmj6tuq5TC1kmK1o08iGIIdGgPm/Icz/5/2RkP8ox/w8jm6JtHE9R+qcy5
TB23dCOCYTwAsIBE7Yc/8hnz5+xxLLzbI3+BAbC6WLcuZ17WbiHoBTpIcq0WROLqj5VP3RTokiJt
mySYAhARnHEEWrBAPYNHcBZ8ovtdqGeMIOQ3d7idAz+bK5tA73+jh7+fHivkPoW/DRiOmj5uktWk
1ywlbFrCQCPge0KveXHI4nOXZYhiKZ32hZ6OhP1WzhKv5H10PM+QHHUlXCvll60VW3aM5WCes0zY
Bdl8RKVpmPpRO9VNorlF88EVUr0JUkI89F9Lpg5SM6w55b6lNAf6zQ+6mrIJLe6+QxAbpkcm86eM
BaQwqW0hQGTTKfepdup2gbB6vCgFxkS7FvnpUybYHsICKdXrrbUAg+1FMhy65k1SLi1EhdvwZct8
sTSTxV4ZXY07OQ1W/lE1mp7lKiqgL2oj/VeHD0q4aoYRShLVnAyEM/hGdMlI6lY8QVgqvFyJwZPV
7m80QzRR8TUZU9Kv2lzc5drW8jO2y2eTW8JxTkOHE5Y4ix62zboHn3+Y0qTtpmhvk9LORQFdjLKS
zUbxO+dQyUAnQoI9gDTLom7aSTICz2wJ0a3wePFFt3Nm4Dad/p932Z5WRqQZMtQeZGev/+x17tuZ
JSSSiRWvndZwTq5wbWixLGhGeJZ3c689083qOYvyOj8np+hQxYYfISTf0JA0NRtcXg+6oXTCKXFO
V2jVm7BFX65sXAHOUZtnJs97dsXRVY6ExBqI9miRcKSJlvlaEKEqtV/kINUQkeNJ+Hd6HBJaqWKy
DaLpWXCWMqgDwiQ8WIS2xRHfm4S7AKKvO7+W9Hog5Mzz4cykVfhrxNIv4XMnvrzqrc75G904MrCs
ZqqoKpZh2cWs84BEmiXkAQsOEN10Zv+SJxM1eyfVBASA6A6xcPDQhCG0PuoCfjwCPaSrLOfGE46+
nrUGF8ayv6RmdEdJKGMqGbyNFrqYme4M61ytpjff02Tih3aY5cuRtxdNzYPBmvtpl5GPP8v4GHgx
voxn3kP2vG4L0+MZVVe1NpvxtUWEEI6nJ2yYgfiyoIjJK7+G8oVj4Nwe+PfUKd9qUDbEvfLWQ2io
kfoZ1mcm9UenxbseBpzxEKWZ51xO5xYZ9SgCJ6ygPp7KxaNm1vU9WRwUoCyBkZBhjRlxbdRu3IGp
K4I4sjGSYRlBneXfwqHaxIPETFcrfEpcv5eop+JSmmvjCSf5TCdDO1Fr+VvacYN1xpGewt7euJwt
MfAA67fhTA7BbEnwJAm4cq53866bILpW8t1Vd0hIDaF3YRSkivolcWxG5PvSJTCJ+59+1vTpvZ6+
xgYxEqmrv129RCJhTrDC7BR+Tq34zTl3kfw5WyPD683mNJbY0UoDYfStkP9NvRfUKJa/UiKsxWa8
QboJlv45hF4wIFCVi2HZCQiRl+nH2Cp+fzJAyBGjDq0th4EJCfCPdTJ39B8aQmGHwov4Z/Fs6/vY
O2J9HpPmcpxIw38JbhmbdmrT70khDIhWXkLtkZ90dp39ja9giTi+++k3c2Zt9XG3RqLw5V55Z/hD
qxc1Vci+lcpn98GvDdkEzXZUWImDDG3krBFTQCo6SqJmy+f8bc/Bf1sQsr1fU/TtVjYwz1YEhiTq
wLQQq9Lse01X0W7yGPhl7nJXyS/hSZG0at9x1OXJnOsQ67G9+pDJmQR8NCCw88ry+pGSPlreG4Rt
jOBEn0ACWjWVpQyTDQas3FngiccyPtoj+OY/hHW3uOaregMv5IGkORqbkwup8Kf8CPwgEW1zkEeA
rqHBOqnK0IiwXYcLvZC1NUDObCQMbCa7Uz58EGtx/Qeg0j72OiybFgHSVTis06EQ/sc61gScB6Vq
51XzsPUU01NGJhu/CZO8uonsx4SrmDOOQThTzEf8F+kbVhl2A58/+/XJFKlg6djPq+0LTyZlXxAK
uU9pc1ANGIoHMfWvpjfu6W9IxZZT0/8L88RnGYmmsWSsTp9AsgpS1ZxGJDiBOgPJNs9lpW4nS0c9
Z1GdM/lOuuzJ9hc5Fk38S1eQxolL3q7Zz1j7/ehmVbrC7IrZazxnxUwU11r9nFx7feNefLXUiNP5
SkpaoJj4/Mzlmea4ggKRvT1T5+To5HYOGIPZzexJuNLqXJsNEJa234zGLz06XT133sFKNJrTkAD7
oiU/6XbkTssUTVBZimhwbPOINBIHMOu7dl7982uts6O1vXUdL3zObgMyHrXPS8Eob7n6BR1ZxxsD
FZ+OaekLLSQWQvdJugxbEBm/I17JPVM/pdbAx9/8+9agmSuItuSLxGVw95v30WWDGpMt6f0IV2cG
Vq6eHah+MBieLUadGfcAVAOHkBLikjHm8KH7ZF+gYAlYki2mYt2z9dBYAXUpOsS8sIPa0Awzpoa3
0QNnoi18sCc2Hyv9fBoR6wS8xKfosYPqS1C2lHvPDa3g437iw3LwaAeFLhFnTpq0H70es7p1mMw/
H+x0RdpSfvDpD3Cp424a0wQeiEIqSEU8a2AxSd6bHJND8kF3jFeIgPrRhGKK67aw/uxDik6WJEaw
Y0Py/2l/t0xSVCHSbf1AVz/E1CkQLc0q36fggJdlNqKY3FilOQgg2egrosYpnlUxWBQVtsS3pkwo
bxUsORQlFpgI2mLyGGzJAsNHqjVwGlgerLDhf4VVTorkVaplWb0Ig97k3dXPbm66hsN2UA32fGD4
uQ58bj1qJglz7YjiPuU8izatocFE4jjYp4fMDY4LF/z77MjFbjrYwzXR2u1tCY62PR7UgsQE1XPJ
Rpmxi/YC+AcE2ACAXm+yJ6HYAv1OzeXEUFMJUYo7TiKfQFEhA84SWgc04P27ayXySh66LQzGyYE3
rPa1zeFqhr4yvL1UcmvVbqsCyttYozhsW7P/67YMDUcMbWwcBKrUAve8dyZyIUu7Oi29G/5zTHbe
bITqYCzuydyF6tqrYtKsbHuM9u+Qnm5Yg1iYgx44ASDvVB0VFTnAN0VAVHRm9ZmwYBedCkmVcM7C
LqGmBE1yT9ufsd3IwKqn998HTOkWeHnI4Qen/mjHhtad1DCalMkNVvFSWUMejOlgxU6m26byGeMm
3fbFqTxffsCaAH5tKimWDTpIuK8RdNShY2h11D9zJpBnTelmfGGp+JhWip9GC4pmk7BQbCyjZvdZ
jNCdYKSDkIdZLMWeaJVJoR1I6qCIUV5OI2ZuEF3UfOQ1q29qnMAxN/Kre0W2f43iSg95AMMqxulF
vRakSJNXk/cYZUxfkgJFdtES//YBlzKvsYtZKjJ65HC1jWbv3kv4UuBeG+tss23taYZCSr73mYqn
54p5AtX/SV3K+QlTSB+TQdvdtbi2HuKwCXD2qcovNi+d8T/AOa3rlTZ4Nz1rtEDnFXubBr406Xu7
S/bplF9i88goM7miEOfr/OJ4XsNxSnKvKaFQOhhObBhW+8wiuwbdZ716qcuyVhUsenJUsuluHZaL
Uo2puD+SQyGPaAsbDtJmNF0M6RRUTR3iruh8vjtGmwzeVRgcwgNRIsPz6ZvmuaF1O2T7MH2OECjU
xmXi9P6VtMQpzTIXE8sTQjZm4oPq+Z7B2hQUwV+FULda3bf0xV1Eiyv53hxFVKSJh9eRgfO88Rag
cXMmylgaKCAlVaf6QKrzd3S1XE6SY4pwO+qvD8oEJyHiBacauQt7avQpHCQDPNMrhYUepHzSBQrY
ZgNfiztKK52Hh4puFkErw8wEs+4nkl1rhhyFw1Bh3uw2e1mamUz9+C8tEHf0oR6/ce23vySus7CC
gIdbVDq36g39OtsTzmzRixFV2zTkaaFjlqPd1BvjimhZpZs8SCAHN79UwUoM5ZRtkEBwNO/UE1p9
u1yyYN6xZZMXUi1qaBQmpxMqMMORXkLfQN6ViJVKdmegfQKDKZkzNEQ9SiXNwPVAnbnrX/mbAEMR
PAb2FX8amYrHaRHuwuWHQM0YX8cM3q6EqdHkXNo/z0W9yj5TTrwMDLItRUdjx0bT01vJed//kAo+
IxoS9GmRYwrZvfF/uMXe4wUkEKBOQqj7YB++eumXX9FUtYTiva3Tb0yjNZeutgpmMsHHm5BGZo3m
Y/dSWAlkFuQEA4I0nFLso62t9zVwGME2ge2HyfuEOHIfEBcxS43um/sIaJrlHalPqMGoKloPpLRl
UihUG7KGUCEMxIkXiNQl/qV3AvABsie0Wn+FRw681l75673Ayo1HSphpKwE/TlVtLYzrOXIB6tAH
QiqjsBt2B1Uv+vIwCSnXF2dQKYUpkM8m2FgOZkBx0mjM/MnQqtAZDhxkJGVPyzxtMoRD2PHlr8Z0
QC9sw3/yhaEWqX0eQQHKtSYLk49+Eu+JLi1lunYsxJziPubv69VtQYjcqWvBHiRWzY1+0+oXWr0h
Bl6IxK3Al004nCAbUH/DXpXuAm/55n3xPsS65zHHt+XsQd7THbN72ncgtoor06Xw6T1FMohH+Ydo
FlTIlBehzkLR8DTDkRXS5GcdAAYGGZ3E0vIs5CTfcqgzzk25QASh1XyFaG38t/OJrIRTWX+QoNqB
5u20WYRAGXVjPKqxKe8MKaF3sFxz+epwmRp4iG93lreywApcKPEOeu+XioZLAmy5xFSvdCwz/voI
k9ai0TtiursdU6m22viory3905O4YqzRZELcHbTwECekTmGzHKN+qZHV0LIl6zxP1QQwRJtZj0uu
YtclszmyTDauUNha2ByYWbPuC1CS1wGkscihCYkKfM/fq6tZ6Bu348HnYfWFU02nVZau6g4OxbBy
H3cgI/poMt5TK8hELnBwzH8GU6saFS75hQg2ra1WYuOvfOwJ3f46wBNpPHP4Yq9DXFl6cftk4DWp
Y2hY/792Z0lCKeTAC8QwCXgH/oacS1La4bg1rD6bmKuuAOI3K2WrumAqtiNkjV0m/we2ItXBSY2b
cIBubroUhfikYiyegDy3xkz3mixBXCG0dgbHIxQCZTFYMtrSduVgUQI9y8yaOSpB5P233qSrUvye
wKa/Z2IQKapg3tw0qe67mHOp0X95WU3lRTq3cJt2AwzceHbywErdNIbkDEzXEXK1eB5xrqRXgMQH
yAJzfZJAuL4MEFg6WnamgzAHmyEyam4iJANnObGEi5xdDnA4V0GloyAbmU8/PYIdk+yU/hZRO24k
Muvo0YuvuDfLNOUnhTAyiMnD+6BEdcudWwTFjhYfx6+zQKHiYEVABm4u3a6+Gk6BLwu0LmDGWrhx
ECpPBlbWgUqiA18elphFUz+p9vdCE3kdb6TeOzBDIe+aksWR+WCfSeJbfrz6/NyHXVTzJqiCoIxi
jWvncblKJZ14/uwPVyYFYYdiTKYw/hVPms2eQT2fQNipgU64Lx2PlHqeJuW5b1wqy6e66kz/SsNf
N0YJFWGSMtjlqiODtdrKAqLbHz3D9STVOU+wW9KipRWw7FbypDbeVJz6lqlhFCMRgSh6pmeE3SLn
cBO4xWqk9OX6yAuj8I8aMsU3gx/ees+M6RVrX1PEiKPAf5g+Be0r7wPfG2F6ZjpcZEsId1piJFEU
eqpx/Ot2gAiLqm3ybgijqgDrclbdXOZLZrYVaMb87cZb1cICyrH83Bxi0ipZ5LwrWs62o2YRZhQa
aukQVpzKt1SVbxNki/Fal4p7wP75+9bcld0HBBFX9R32VRuE2oB+JumviU1HwfqNioj4Yitf9KFn
wUuIqyULqk9FsUMRc9aLLzH5VpYkhVGx4wfbZBR8+2mEGVdiPRV78DPs6UpV/v4oAMXKzdEqK26p
ajDyrAaMActmzETEPMxdkhN4syMJjmmomFWcwR1BtRJHFkLtEZL5KsC4khTXgsnQPt5WyRKkG7MP
ibpYmsdr7I8tsraIOZh9ncXlwsAf0sChs896VajHMfaesu3V1C/ihY1Bb60NnDVVKLRhR9yYs68X
S2bh+LWxT8WwbxPpMCaG8aJspit29Fd+LLpd1vCNRDNRTafMvuiQhzaryY2bS3xI402+HubZYkRV
U5vbwunlAaP2o6WVRfjtJ6qkdLgT/XE1bzaCBOOPsBRvPPLCV31KC8QeMq+98mlvDwEIDGwni+gs
MAJXLcd3deW1Qz3lKVczLw9DNP0cRfetBZ6lNr9q1hart75UmepXei/Ac0zlhGiEdz0JmBVO5oFc
SKijK7i7xbYjs0rOn+NpXUbCmunBQhz7qvb58ShzU3sHEOGXVeaIEEuTZ7A57FR+CgmqETPI+DxC
3LKURtwjx+Yrz8w9uG53S5JtTkE+GMhdyjyG4UDTmips+Dlu0BuaPjqy2PcmO06JDvIOKlPAchEQ
F1yh6UEgo6XPWyO0gmWteTC0GnBT5OCewaJxzIrClCg/WhCntHhLeEonICGxqwO02CnS4iAzRgUf
ZP4hR6XHRdeqS6h0vkanuq3sk+HwAHzdfMusVpNA8lDfsMtAFBHeqRdasaVTPdDAPbxpVKE0nLAQ
4L/3e8qoOdSHyWYz19WO6DcJELd3NAe5l+htztgMnsF2F2xBqf8A0R9nh1gPWVDMK7C/r8C1fS+W
s1WtiFTa/KQDgnyljhqkSZq80JPB/XMp9sPJSoRz97Id8KmlPEvZY4V8B4sNDxTTRHyMRxd49kNT
qfq7tJCVbK7xFXgJP2pMemmNw1Ifmcoh0Js4Fzq19Zw/4XSJ7zkQR4bo4OOBo4E24CTDtXLpE/g5
RdMLvsbmNT6lGEMaApTET8QjXhIdbbrOg6aqQJx4K8GeJWoOhKqLwKiq8Ugf0NktbwN98Y2bRL9b
Vuqbed77D92HXGf4lz8kuN0pSHkqY3yarqVH4kaK6ae4mmsSzY/z4/Ibwef8X+rASlo/Rm3LoJAM
9quxGqfubslVhnEEpK33wzaoDo8t23h79QXRV4pDrJbOMjs3Uq2J8MMaLDz6vTK0XI5aDgWAiuiR
PvC3fOuYRrYZOxjpH4MAC9vmUW9oDTLL925C5d2nkT4IdzStmy8PPu0kjvLy/+Hek7iYAjOBF9Vl
EeiQskuPPRClbBa16lWjZ5s+RLFKPibLUaZErcynuurUZ9UtEwQHn9l1x2Me2aHak1NyCm2Y4MSH
tziRsO2dIozLosMQXTbKkB5c4ZVLgKhea09x4bFf/K1TFG9nH8fFCTM41iUoKPfs8VZfeg+H7uba
NCtpVzKwHXkuJaaJVKTdz4hgfsY9mwxAKEw++uLB2o+sFxfMxQ/YEhkUBqUr/Pdn0IXpEeGhZ+u0
yjdXuZTTT+n68R6CRhG5qsUTi/a87/5eubDAhHbB9FWDTJIru06TeWgKV2baRUrYlE7dOWhb00m5
WMJhEDs+HGT7/hwX/nf/RjS5bEOlYWAvkDOpNS7apRBcgcnWM32vdCa84KnUrry6CQmwJAL3t8UA
wsmWaA6WzEcg0PyK2HCuE5xiY4DRG5CYaaTnYDhjZczPNjbIV4JjjskBfs4i0TYr583f0ilsLoEy
h9uvn5KX5HPShEUiO+f2gl4IFC82uSoWe7MMFHLZMKJSf17lAqoDumpTD6lcOzETrz7xkl1Ruk4e
mEdCfmK4DpSo4P8+JdHY5hGCMshfov6EjvRJKFhhCQKJGFYppJEm8inlcNFIitOMpd6xiF1IbZLd
Xr4+43Qaf0W74jTGoRMLMXghHp3Pyd18Wor5fvtHWsYhfY35i3zx6Sh8g4eKDxBx7SAa+lBTB7Lj
NN9xFA5F06wrG+dXUdU0nwI2WjrDwyhjpiL5zEAy8rwwV9xzRi6/kc9mzQv6Ll6LXllNNtwJDeqD
zVjjDOo9ZPl0ktIM/sGQRTwxCH3bxWtIN2RCi8YVQDTq6mSxMu/bRE+OB+gD8Yq1sP1BNLSoHlfG
eD6W+wGjC8oAoe5IXl4zQDDpULjqtWnqv5yTj9i74oMM1Sb/oRb/WLO+GxjyWK735Wd2C9vX6b1o
tSc8htCHKzZeT/NpFYt5pXM0zUDQdOxX+OkfTPYdIikLqU6ISkVp7+m7BV8Hy/CAlrUYSe0GxuWw
dFJ4Eut/b+iiKU0EU6HVNRnmcfIUlPclHzmhPc7b+MVSzaPKDKH9yGWWrm5HQNFGetOVCmp4LCmf
QscIiifOvtdMId3chy8Kf16SOnvDdKuWihF4igbQWv+Qs3Wwn23i8gSCGWtl4P7Hga/rDkD5MiUs
hl1zHnX3FBCh6fW8tE+dIdlk7VB2+HxzMvq/6DdSsFnlz0kkNwpxZakBDjFyaIJSqAI9ZzwXc6nx
6dXAHnajMErzWKGwfzBu+TyzaORPf+h6E4wn7bTa/NCbQh/EAdaHEqAhg9A6lynBskJnb4eCq5hn
0UoUhG8pZObvEcMq2WNxsv9MZ+NsUHTiJ/Phh9Q9TCXoIFQfVn1N/mdbqG7KISGy94XCqT5XCL0Z
+dD7yW1eB5GLuSbLtGlGfWOJurTVpgLKYPJmTdJVyRwB2yE2nwPi0ErFfgf3Go9+H/j71HhYBRRk
JQXTrFw53J7Wfip7ul3q7p7rJRzebSifeIHxub5ZeYk16LV5rVDkmdn1EAdHcHKqS06KFL0JDH/o
UtVV41l695bj4NjsoaoAfIfO85T85fvAFRHtCTe496iKh4gnVMOU4hun/MN9wwduYHlZmeRH8e14
Z9wDdB/HwXPyY1o3LlAhBCoMTetxwcDocavdsZjovr4uX5B7gFddCX/orKUwRBNd9I+F8nMrEmM6
Pt+oBbDdX2z08HC4chyyZ34QbW3bE2NMv42vcbiZd9oUIidel9a5xjeA9b4r8ntXFa9S1B4GrDcV
+HEpB3y0rgwmZiNioyMAAeeRFk491fQZJFuMGJV7i4doq5mwZL/cbDb0889jfU4JJ7mqTkgVA9zf
KGW1t1R5vnSiM0ochcaFOJ0Q1DgRBW5sFwXJX9iQuCGsOs310fjYJsKHz4DCDuQSvlHBGU4BdJav
jcSoB52gMMp0f5BfxeKznMQuwfmgR9PwQxouE61s54Fb7tAzDsP5PYeeFYxXLWHnUt4Jtw4yLrkx
oeyP6PB3alez0T9Hx/dl7/nSjySuOtiEe7BOdYV0mFYqYoCYqFx/7urbrS6gnt7BJbQ5RJZsY4QM
Kft6rsgV5RJGulXSdngyaGHCY++uveP8l7RK9OfPhZUynjw2t31VtTTAwiOsrgvErF/2RVsrxF5J
D6j8Deq+JWhq7WGiGO7dxe8+ExfD6BxCF8bSfDX7oLEKX3NXfL6oGH7Y/kaANXs02UVSaFrMOMzQ
G6dhGMBueIXq1xKd99+GrrZTPtWteuy2tLKRKvxcxRyfKC8XijAdVJFMyJg1RFP/WF9YsKFPeaT7
mWzgnv4EBDYZ79CyHmgD8BHr2zJJ+XoVc52aSpQYQ2UKPoBZex1O5e302kAO4WgVtQAIcEYTbU12
vysJPx7GXY45oAIY6eVWPv4piWNndRYxRhQJEeC1x7DEvK3GHnxjC2SLWAEubhovSOgiKEMl53ox
l3cU3kwvwxEnt9314Wj6acqG4vSe4gKwGJodQ4V2jbcnwwTYU81NDo7F2sT8R+sDzbBzO9M8jclr
ukg7xgfQg/l2Qft5v98CL/jJTv4uSk4QNm+e+lsnH/HRBFBikpMfv9bIUlAkL3Mnd4qJvIvDp1pH
NFWE5hUAR8oRkyL7FM2xhvqPKInlexnJntrJhr5NuOw6Yi33hZMLuJtjdRRtrBINwnMKf4yd+AjZ
hVE2ULxeNd3VBBNM115r7uXKXYmXulO6+9badbxvMloIYQc26XoVgrNKQU6FVI53/B5j2H/rwFcX
/s0NvzS4/B/tVBc3WwGsuYo6hqqW8OzASCFq5+u6+CciCYVpj2jBPuHbc3vm+EwhBPegDFnfCL8a
IjO7kll35huCkMO12l2NTWNFExFqXmZeCQaa32tEoYlnUKne9Wws0Zsq2YIfUhWx3JK5yQs0HMin
kH8DZaBhXEf9zI7oKcY++nO49pcWvNxkWeEvMfKLN3cUiEy2hdJu1ijdFKTL6AqNQBSZAbYcHTaS
vhzALvVM3o7vBCmfGH3q3o3x+woVYp6bqDTHzYHFu12p+fK7Jsq7DZL6pel5f6dsLl+bIOfpJOw3
kBmFtxd2BgFOFVxv8mLcfgybOha8YlKUl/gNjY4/jI9HnmLMzx6vmyolKiLr98BI0ZQC0WoodX2Q
c30OSn76kVSg15GTYuvlGaD4C/R8vFZqUwOrFgt5jv41+VATkC1lVX99qn43bQAY+7Yo9dz/gxDw
4Fq8Gg0R3/Zn+TFGfJeTmIRi7esHbFsuXJA6T2J49/OfH8XtYRyUuuDjblA1w2mCE7E+azTN6fIG
EUZsrGBQmKpMgjtp582gF/V4P6ji5H5vykzdoztk1KtLlqz8y8g0S/8RFG3oB45RVwxlLeIjKb2/
zVtT5ifNsKsCQZZdhj3WVcMRb6I70cIDOF/9xuG13BGthkWI4JX9VwjsdC98tZmmxaPjplTIAAS6
g+4EyCc8cpIwMLUbbuQ1qX2UUHMA+Nx7KjwR+l0egBbWQPTmaP6uiTfqfJHPjW2GjzFNd5Km9cHT
SCh2zVIl3OCCfvEgxeTAQn85vW8EwDfbSN9Ir/B3UzbMpU3P+DmRqR2hhKhLgLaXFCcvGVdYwoAM
EHQK1Kejsa+KL8+T7XuODf3qDiOVoT7NZROhFkCNW5h5xtYG0Nwmv65Obkj7SYBaPGCsnep6FieJ
Al2sALe6O9iLLUTjnHEvvnMlVqZcEeF2eAVmi0e3yfiuxinhONADoeeXNp04APkXUUI/JdzjtvFh
H4FcgHRCgze41wxD+ivpQU00wj0mluHfmED35IV0n1rhZRFQsTqYmOEnXTIdKjyQ/H3DKhCDL7Wm
ynWHJ/6CgM3ZgkOGp6VVdkTGNA+ja0p++HNai9FPSBQoZa7AMfHYa59yKDNy+c3zhonMRtsq+/wj
ungyv7GRjP0dWEsyUlwQrPqJkzb39Nl1LvvZcpAEjdK1sj11omB3vrt7ZkLPP+sq6rupWl53phVE
1s/Oz9FN9ugmraS0emrs0F5b9KNBrRRKTe7gHqxIKtLosP7o8JY2Mn6i9J9cVKX9U/xbIYRYJYXx
7ow3XBKLHcVZ47FNaj0R2pFTpAbl75QrJNWnIbeRPJsgOaeIKnrZuS1bfFDdM56s1VbAms7Rs6Z/
ljEzen+CzOYAXUqSyL+9z5tik90HW3oECtoccevKMrgcJJnAxEPoUkz/IhlF1vOm4RDLiKhARsHS
PL1CgDvN+uYNe/uNabd8hAzOVGSJ1BNiF8ycYzfLUc36EAYAq41NCnGWYr2HBy/iRGjdJyqEtWL5
68oLRTXJkoQzNNfa/TPVdwOv8KPG2FRDVBdArxB1tlQ6wtdhgESCUI9Q5KP6+CBti5lwA8tDN+L2
soBhmiTEacBcA5eFgo5Uwq/tJbkqpFaaV7JaTc0ecMOqIKQNVKHgIVAMJ3P8zhwQYUD8ZpYbmmeq
DOvcWIrf1oOpnOe0UOhiZpZL6M1O8wKSfYDEnWpyuWalTz+SAk/09QveUKHWzeqcY1zhtgG7tgbd
Mo+hwjBb8M8BIPakka7Ygnew6uRM4xXORBBNjzsqdNDq47JaoYCn4itFbYeotIOeRu+m6Dz/LYa9
3BKpHRgizoqFZ06o8e6USafP2YFONGYzLxJaaOtE3y3Edu2ql265dtRBIUBXklW79YhYgrKtjP09
IvNnfdT7lf14iVZfRmO5jXtg2w0NhBqc5OkuRhjoIj/9VDrPu5MuGpxEoh63WkZPsMolg4EhMZXp
5906K0w1O8ECvFsTP5iL/3/o7X5EsjgB1vIed70RbcrV1vi1fxq1ZrDDBGkCzAyyqhqqAiJROrIE
av79jZKaEjJjP59fCK1kGMl7RCAr/TGDkgqWgEfb6pvePTaxGgmKdk1Et6oiOn8gHuDzSgRV+WPm
vJHSbDflgEzoDxxjZld6I3pJIJj3EAB5LOORgwqByIwSVoKd5f00thLnfjW9WETXcbrTgUaSYmo+
uz0wYfEctcrsSFDdrtBn48CLPak5eP6ZROlSH+Xdy64/kteMZlPlK3LmbvAFpjYRhKj6mfzmY5H8
UOyNDP+Z6cuAhqVAR3xph8Y2FU+LQeim+j7nbJbzn3hMhlM+zRiZzBTF8RH8DspEJyfZIGv1QXhh
PQUA/vuVRPGsjTqvBT4LcxYs1GU+UICLjOivjn3eOIpdwTnQUg2p9is0rDZjeCyIIGOtMyzIEhtW
UigzLfs90wyfUPbq2IF7KXcbi9e567FEAwxJ1/YANPTTZal/0X/8QpfmotiptufDR7ODAkb+BS8e
tbJGxoAcxaP2FEvFLhmrco2qMdyNSz6SNdPmafdeqNkId6B/MRciwcZebS0daXnWQfjjA7Xt66WQ
TyMTlLFte/eYo5J3+JJy4ZfNNjBSjXClzSC3cswd2Wo3JrEFRJa26G2DTAL2bbPwcMO/g5vDM4Lm
oYSSE4p3l93yX3jHS6l0emsbBRp1/+3ILR0+SKOpeB8DoFYOWpnj50h8F8jRl7EB+UulsgR+eiXT
pS6Vt12HdiPOH2lBXx5c29b/2rzkO1iUpZZSh7cxZ7+rmR6SsLivDfZ7+GJy4YwD2JcycArLU31Z
8ZHkdwfKpaTvAZ1SNI8E9pkHy1oNLFUh8ifDCTXZPXYOXusUZppNtwWgY1GsD6zTyFO8W4KKgKyj
y4Te5mOOuArLra3LcEy6RQ7eGISnttPzXUuy6REdE3OXYQ92CrWHWA6VDVdLewpl4YThChwpx8cq
JRCMd1qp2lmg+GexwxWw1ftJoekyYu9bLtgXycu6SPFbcTvTpuOyRjCF2G5eP/IWxY4fF9nhodWW
aTivmTA0hlw/Q5+vDCQCoir4MsnifylkvHeg8tWLcTPRzScc+jBkxB4fkJYc2gazx5hBzunndyvG
ynJPK+ZJFd1hvlA6fJm6ORfcRwloRQBRa9NpZgEoM3SexCcpXLMNk1LO9yF79RPG2s1n5bAGE2B0
0uU0gvtA4bqLej/t7sMWOKl+EUWfrzINw1bhgOFxDQ1Nu8OJeRhfr9XDo33glstbJprFdnBQSaEK
EYtmtGN+v/Bx1lPN4zKGy9LFLMScYQwsyzDO/Y0Xu0h4KZeaDBvRysIkERdV84IVvTYIi2avKZ2M
X1+5wNxfT0zemUnI71b1JWF/U1YIlTR5wQM7BAWS0nR0dyQGGrkCeuYIu8sFE+YebJJ8dwhoPCrg
AYi3L0jsLGecwv921pSZJG6RtIPbgTDUtgx9rcFoLWB66ZF7VZW2MycEXf1X85g84RKflO5nK0bP
f0H1ifgWO3Wej6yEKpymqvFDDYFWZltbb0+yWz2LwXB3yIDXt3z+uhLcfeI9XVxXyoNywskqqxQp
0NCLOhaAtQJuB5pauqkOtRN4a/PsKE/v1TEKbI6v2SDnV1HMj+N5RKflPift//gfrPm40JRB05p7
mo9vNQdBz2FNvwptXPiCFvCgZWihMg1/doXBoBptYDcxJrfk1XWkZ7YCl76yEFWzEw6VsmBoUipu
zCffKCMP+mlxJqiY2QKZSFUZ6tbA41nc6HRVk0vNyK74L22JYceAsRlyJjdlczCGNH7ISGHMQCV/
1icXplaUTYRi4e8Tv/Be96Av+3H9JprypwGYZDFMQRfeRXfchW2KmsSgIdO7a4R9XiF/CZ5prQO7
4cApxtMIypWU7dPAwb5xVo6IMNm9TfBxXgSk0FQttjZyDm30LTjh34ouns9ZrEJ2gkeh79OM06Hj
UHqzIRjSCSKil8qeP7oljI62GAC/dYDJLBQTCYgfn/oKtbzujUKbuR1XMAjnvvxkPKXBem1xKB9r
m0Q5SqhXkAa8xpozA1BiGBsMiGzDTMfY0vz08n7LCOSB/MUhpotp6mUCy41u+l/2af/LZbRDx+4g
uInKyqCjAk+NOtj29YsmCbjaQdDXbqL7Hi4/uLSBIb1FsVLKdVvGcke64fO772Wv4JfnDgFubaur
4Kb07KmUpsafhlDF883fsrnGBXqUlDFHIxPShfJP2CCu/kyn9ZhCpGt2JvphFtmq8ui0IuuCaaRF
iHoEMrAC9jcweIQiE3ZRo1YT7M/ycs5dMD2dpWpDy2E958nShvDcPBJ8yBQh+G7n11FfQ1VuJRln
ETugd47VoVJoV3xg3dRxG6x6OkTBS4YvXyZHSkM862GSs/FVudpU+4N8ay956MBI2FsuLNr92DV/
PxYAxovfbMN/UkVhv0s54F6TzE44ATj9YZEJU2qoAW6ELgmtsJ432rCJej4PUsnRQgQ73Mj+fGLx
uW8PTCyGHX2XVNIJRlfabbW+RdjhwZc+U+GBsqAhlS4STxhzN8ujI4qO4NGSSo1KaV+B4j6uURE5
LPbf6TslbCkC9Z2/XlDxO83Yr/R4SHY86krBDXdqVvvoqShjvH1wy7Ed31bjnQw/5CFfvTyLeIqL
xHo7NFYwP6zF19fPKBmfMxyJ+dktXfhX5Y78lbVFAu97CR7cuLIGmCAH3LokjycpvXRY6jCvsRLq
2xHSE4A+HSWFzVk3tZXzA/FiZIdaqUUgB2CFlOYcHQ35q/zwMmLHFttVfyOmnUHzREu3jTk7F69u
2ArxQ+aUc9oYf4sdtE/Dc5Yk2RoGpD3BKmqjGUDRQ6hlTfiCj6lhCxRzxPEniq8Iqou0X7tdPGOb
dbWLWFl2SMHopVl+vtxatwEZDxZAMOEELJbiDQPbDzbq5KDdmU2pLaHPb+wI2s4qjqMoiwemUxTr
PHgyOquAV+lVrztJX1wKS8xMXdzWrXqeLQmF+U/3rOXulhoPWw+lcDZ/brEsBGGMrTKQ3N5fHK3l
eXDusImf8N2TrUp7KDeD0XcgP00C0m58RvLDTkWpLgt433lSllRLIuINnpPOScLI1D6GWdnLkj43
v5UhNK+jb4zMCWj+pJU3oXoE/Wm1DRklLdjtNJZGqUTnMlxNcMAlDxCd/UPbVfG2O7dmGv4YSDOS
uU7QE1Pkyl+lpithE0+yMT28+ROf9vAkVKSXjqNKFZiaKEr/wvwfETBFVz2bny3ISBL7nYdzyO/s
JncSL3EZBLHudSpXuaU78X3FR0rXcpJQwtiSE2/Gar430qKTb0gYKifIfQKrOdU7d8ySqf8N1ibi
LXiFV0/RE0MysBjwf7N+3BmXC62U2qKCmTYsde/bgEOIU3DA9S1mFWRPpWbmn+CvEMxbaJIDQA6S
/E+tddpZ46+nd7BI7pJbCCeQOWw9HJihT1RDzBE8eoAXM7kBCumDEmprPkejA85jPFsSoy4ZhyoW
0p4S58eITP035OGgTloChFRgoqXPT9f/BDpaoSTexlNSXKh80M1DFMdFjei8UOc8pUyMBNqzuogE
0HsmygsLOi4NZTRwgxiR5WtnoC8Iuza+IUrs/wazVmO+R9phHg0mL/ACA0y3weLJnUX+R2aw1uM9
EeJFixVkIArZN0xrk0/gPoVgEKzHJI5E8fioD0H+YlW1HxhTXWbVynfGO5ppn7qd8bjxOFJEfgnx
ieQEL+5ioeNDbFIk+P+/XTeY0MZbMcW0SFYDb5awpehjt0yjNN2KPJULOVVhSo8cAsp0kw+gZeM4
vm/YGBJMv/cVFLBSq4+77NXUD/JOsHuYuIrNRvMaaJfCV8mZ6iO+Ix8I3bfx7RY+y/nnm6PocM+M
byNEsrJyjTGJMaB4shLJQaC0bABmRX55LVzEYMIax/Fm3kUMgrYsu44J5UMmOI6IUGjFm8t7L2mM
wXqvy5XvgC9T9FiYnGzq1Gvbhi4i0RcmW72XfIiJKOAP3ud3V+9ODNuMeHWNMCgp2y3h7ruwYKU0
6n3tzr7sHSD8CKCIXkPIlM5Y7ZhOkYNu3M8aVsDdW+XI/9+qvmZyKbUt8E6rPeyorYqVThv12ARF
RRIjvPPij8D2owbBeCUcChSnxp8p2u7Xe5CW9yGktSszptZ+GLu1yfScOGALBfXSI0CirFTRRrNd
1q+pCCSI2HRY6lFgcvHJVRbEqA9hBPhCUsmHXKqfABU8hHIvU3FQd8zOoHGzdPsZewjwDSLXF4ex
kYO5tKdPNegs5tB9OTUkIrej17XI5YPzV3sHP9Ov5FEmFHuKmy6SNf5TKPeaFPlLNEp4+E1uHc5c
A1SwpToOCdde21IVE4MyMjCmlhGgYvWqEGLigPhuNH1kG2MBX9Hq8Vq0NACOUKA3irBXWNzUXfR9
YbygcNVtfQ6EmYlurDFgTO/3fkLJHbpv4fiT0auZ18EMeH9+LLrvXEz3R1ID0qAXXDbLXX1zVMHh
iv1b336lL62GuC/I2oAeF2iaAxYkf9fCF6Dwoe6W8CJnOHF6ssQ5FBEIyP2lA7vayAPXmKFTQBgS
6nN8tfvc479WkjM7vNYyio1Kp1SZPdr1wOexrOe4Ey7eu0z64rnqCHWlomSG1DnPQKVMwGY44UF2
ZqcqZ0S1g+Mf62XU+HX6JWWSUuEuo9BMze98Ghi2XP1AAnmDsTUrSYhssB+8YXrL8Yb7fKBaUUBc
NKr3WjVB3vvgoCXe/Mymo/m65XAwnaHR7/hk/fhQgrkd3wkn0hQYjDEHHcqWAF3OOLQrsVlLT8bt
KnxikV7uNVKPYOohe+emwOaE3Bp/Zy6Fl53Z5FDncxMYhRAuaDKViqwoX4/k3iOcPFquNZ205ETB
Q4yIxG4vvmtJSUot464BAe4C0f5GIT6vfGi6ermost8pqXTlMFb0hpzxH3cGAqHPaeA9gVt422I7
x8p9eTa4HxoHg67NDJ2iroBRBWnwJUNDM+jRvzqphQLHQ+uVfy4BR4RdXXr/2KJN4UjQsgHUGIsI
qL1fo9PJEk23d+WFkILr/7bDsg8LJzxKbjxFPF7+Yd7j8Icc1jW5isQl3p8zb64CX4M/MSMKLo/L
Sf4cUWsBkuJ8qKIwsTd0Dx7gKibyrq3RB7VFIRhyqPV6dkAZL0fbSYYXESSnV6NA2vs+mJjngqXx
7CLeDwEQEjOX3SolmW5AlpQJ3Z9YkIFsx1yY024ivljYRHMl0XFS9FKUJykZuQb2cnPo69F4UUjD
mNt0rr6/sARXk/BvxRPbxcWvHGRbMwZ+KPZqGKTGjGbGSRnYG4I3F6DmA1hTZh1z4IxlEBDrARL8
1y7KuUDbFUEE1HUNTCPDs145CaQEWmUoVC+Zc06oCeg9JjjG9zItFkMJe2Um78ks1vCeFmgVNzda
S1wZ3AmJisG6NE0h4XgHnW0MNvt+7QYiGvMGnFXXn3EdG4D4KbmAZCDtFevJShJSIyFQ/+gz/7AM
muw4WxwYslyHlTzTY5BcKmAKNR1Q+ZAsh6piYKo+eY+6sCIbXnpxdWtpTeYJ9htF3LVV91XcD+Xo
/VhKy0enwm8gxVLEKFy/Jd61FChgp03ToHDnSwVOVAQPLsVJ6Wc7io00shaw/dYL1AIFw/gkeut1
B9jyiu4rhUxk5ENTX4YGfES/eg5fusu98uqbfrHjaPbcvWl0OL4dcI6nUvOvTlSpVw2YLMwtZ7Rq
An8uahruzaOmJc4w4blUS2QCdQ3DZJdvxkEL0Mgapp//4/QNzoMJT+heW6yR1To0Jci/aLQNqKwG
WsUOyy6u+vD3twooOdpsfj1fjqcBaJIzu+izFrwfkTGJdX91XNvIKZKFxpUA54cBHpXEm9ycRVps
ZHp+pVen351i0j3H8a2p+UJGv7YQu1shcrdF1HPsZ3KEBlQgdEbuoEsot1nwG3OslEgY7zQ1Yt6K
gpzIf2HqD4SxUGxFl77IcK56CFlxQgnTdHMIIGESRR/wyMOPvbEx6sE6GyyUUYq4xfB+LCLpaGJ3
qWMjQgZkB5jI3SVDAfGOuKCfJfs5KvhEONHxIAaOPQqYFotLkVLLjCZS7yDTWGWrmhuTMfGDbX7E
z2Qj8EcBj3BQr/AQAk7eBXzOYNxbdFiCQv4PAwV/iXYuHQBXIlsiFqTcTikhpFglIS+uH2AyOyaC
gK0WRFZs4hXf2hdEJDRqM9DVh76rkGkx9yPZcCDY2RgGsKRDNz+RjDX4OKk4u7hLSW82k3PKFW3s
Ra5fKuYo4EhXpCvx6NDTwOIMW7a2BYy5w99mSeocSNoytZ5gm2I0urLNWPsWC2sc6noQVPxz/Mqf
sniJc3rzVpn5/vgfU0GpcIA1GgDRs65+qrGIn8qrDEAJli/tBmzKhaXHApuP4IfwUSdKswZ/2hLB
GQyykbLEhgYcPZLTNblSR1hkKwFRuqdNbo5tjXrCnHi6kk6VzLge/cWRTaRdkOgmPFibkm/ZoYhe
0eruS976MzCTne9IcUZMcYhVr1Lt9+Vrcj0+I+vdllykKhWeqSuwe3+pljxjtWjvnlBrADBG8lS4
9jyooQuXeQfYIhe+DITQlLzXBvEkJIo+T5AW21evVkOb5A5U7n7uAeGvb/vY3R2OYSNdVv5vjGOJ
FI6YbAiCNxVOg/R7BdMRBlVInR7nMnlbNFQie1aIhV5AJPMeT1D6fS+7FiVylu7xCtUvI51e0OPj
2K16POo/p/tssmmsHTOQmLzrilrijao0dWCRSw8e3KpCduwMa4xnHlVMzprLNBzLuItfOjuwvwrU
wQCia0V3wZa6t3gYwPDo1Kcmh75VL8MKA02c+1p6jLHH8puJKW9Nh/aGX4Mp8FCCa65Vqm2fLdFi
qkcXLJFQdXLrx+E0M6wHNQ7y3oLYnivYHwfvPZmhde/e/gxLn1VLpS8AiL4RzxVPyAGlVMy1m+43
VAe4LJdxCauvA8eXj5wR3uJlVA88EWdZDhvyufe/kbnY/TiYSZCiIdj5HVGIlt4l5tVbN3nMu7X9
jXWIuBd1n/x/XLEGW/n6CxVE76URy+JzGGZaeygMbmwk/4qGlgTve0Pfnu+I+3xFhH2u/uzgJmwG
ty9aNYJeKOMbgGGJjV67fh8ifRqDVN9H96Qb2aEN/pdzefJclP54AQvt3LslLjk64BEjiChx/KxN
IUT7F03Y4XEbXub7irnLksL1HCsdjO9AZHTMizz9dG98/9OeQ94+EcZMMHAsfoRT0c3TM6nj9IAx
bDMvPRqPl53069IQM6BKe6l5lolBQeTpBGm+5N1/4KBmeJP1ocBCfvZfMdaFMZI9uhwp05nXG+mI
xxOV9yNZIDAc8Fd+UrV7loLI8iATj4HKFwLs1DV5VXZeuY0sYt0rNpiIrDhRoInp9gjBKbaykwtP
L/sdENJy6xyMBbXM60d7kRAnL+WUuv+iXw+7RSRC0no6YMUefTWMhPr5OuAtr47j7+rQt8rgZWUC
jEj1PlT4iafg01QRMUqBcNfsbnG7d9CwxhU/AiSS54clffMk6ryM3hfl9bJx2PCfwf0gL+by+l/1
xBWnePfVFe5NhCCdVXfbhYDooSoSzi9C9ZvpzJJe/a5+V2GmHYTvgYXbpFW7kiBd6fsBDc92sZA6
NyNRMwNNW6mT/OmMThnl67C3vDwud4tF5A77nNzJHCRy7TLKC9KXAE31FZfKoT+7UNUK3C4Y76wo
GGT7rHiJ2b9f7ttiArnDMvzYt9V4vSlvPqupSXkC4T8rS1YrzRrNhlKRkCfT275PD9NP9z3emBEw
2eHsz0lj9/LSy8G4KlyStfA2WO8swgkbZMH6w4+fRH/wlwQgf6hZGHK1XFjPQ4TApnY6BVmpGeLH
HWgDtNpPtD8P0DcabbC7Z/P6Whip1XXx6eK9CEXQjfJZphHIN8ieuK9mvg031QjzAevQGrdAnJ7C
jeYFFT4QTtyirgZ6xDSsYmbviItIaNl4lEl1VawbuATxYAV+aH09+Z5EusS7gmwcJ7H4s67pgIkW
peky8ni+4cyzbaL/lxkBb8vMHPhNMVmbuE44P7a49KfC9MGlTJx5elSKURXNqSS1eHuvcYKYjE6h
JyfGuU8I25SJK6hsP8b0+6IwmhDHMLgcPBN9OVSIULkKQekTcWr4pD8uOGGnjsKXdDSpp1T4/p1M
AvpppYcq2YhnBrseEjH0m5wzC/01mx84Lj18CVTUL2+PP7CwgXZvy+Mp0OLWsPGnKUsi+1kORhHR
ZpJNEj44dkLJk0exXSkShKDF6S8QpSNGKfSy1cOoK6JFPiDVri4U3mAqA1b7qZ/s+UmrJI1T86i/
lx0msefrQitydJBXGmVYQmUIrrdNXyPy/YncsDyiYhIe16fAkyWHB/Wn+t0P+/PTrX3cdZTqHNP6
7XDRJ1i3u/JrZa7z1ztPBUXx3U0r/MGI0iNEPqJ8+Ifeb/j9HEgz54iz/bCCRyvSmlNGCabO/Ca4
9/TMXq58OapPX/mb6bgXZFxiCH5uxuunIurDT/VzT6Zv6UzXbpO7nBBVVq18xAGi73NuWnX0Zx6Q
nn/yPAMxHmMWuaiS9wkG5V803W2hDANTPHyR7xtcL+rK9d4uno0dgyrU0KpkBk1M8brZaKm0VQZF
vGB1NgqzVuJs8E5XbWG7hcWbny9f/vhZYhCtHkx36a7k9bynef8iPv0hUhSWWqgoEfkNtoSNJfgb
h79Kzfj3ftbWIdDdmfyMOctncrq/0MajjCPZ05//NmR/eAUmKHopH4cXkjIc/TvMCDmXJE55dAu1
Zsjy7e5STr4V8kC1/ZBK65ddBw2cXu/fbH2juP/E4LDvuR/RMCx+N9yJ1HYX/cNMKyLBQj0sjvIt
Wkt2+ZWNnTb+lMqvv61XjpPokbuPhwzwDjnmDbNTceGHQZFboigNfoD4BGVjaDWiZeiWKitg6gfp
QA8IwQBiPl6pDxM3jNmz4CfPh1zZDjBuKXuuMlIqVbMPWjkCe2ss2tq/6nV5sUDk/e4B94KtMWQz
NOqI7c2BjIP5uM1dWv+/dbgMu5ueToi6JXFD+16VQ2iHO5u0Z3WNps6upZqQBrndP5aN1ML7hLmC
4HdVQnfRY6bBZfLqJkVSc0MRAYbKwgkcr/vY9vPBvdeko9LsmwbK3zniQxPNmEPzgWpuG4qGtd3g
+idAhRqF7sMfOzK+sxw/3WugrQbwSCKOm4MmcYqQBShaMCTTa1EkaC+YXi3ZZJqGt5/g5LEhHmTE
NzfOKfDi1Rev8+1FQjyItFGk4yBRXNIr3ooq3fRRu/5oG6Ntso+6bttIdGVPbN//r3nmHTCwScRt
MlbLCFomp8skQXkUSnr9iMc8I0VWthtkL7u06+019MBKItrEOBvoKDc+7gcK5Hw6yGJ/gtjaeoCQ
F+65q6GAyoVHjHbR3jA2wZNx+5nLX4F6yVkQmOyCaZjQKXph3iD7TqsVeWf8uHyvN4a+amkJNNwM
IHz4iUeDheI1+WfsZjgx1rHUnn+pGaWXBcYaO++G2opBZLmUjZz3yZWjBb2QhTdFj3LMM2USABR7
er0JF2mXCc+1Y71c0NOAxx+QVtrzEuGy1AtAO8iW5imrKpaYpfgvDzcpzKg3pmcfoC1RY45vEMgl
uWqZcfSNC3iQmHceLKNrcTSO1smLwWsBzALxXTzrm+Cl/p/CEoGEkFzEhbsNpmqIggP8Y0ySwAdX
bbup7mXk2I8oGg9kl52UJcxolK/GXZdK4SP5vcUS58KyJIwBOVOMH8pX8Gj431+tnWFhWJrZ4JO7
lBNaG/oyjiKwwt7gNYR4CbpDxTHzDma/lYgFxhoxQO9S9dz5Y3VRtxCJ6fq0MfsZemlmb/mxl9Wc
rH2LM17eYf9mT/8LLE/wbpt4lYDavn7Pwya6SxjbVC2EvclX7QT5XUQ5sUMIehyWZPQy5KkI8plo
7/krQUkgclUrFR73M4Wtm7xhGTvrw1ELP6T2DSE7UCk3EwRe6Gt313zBB0Ty89VabbF3CnNfDNJM
092DVIf8ELoEuYlSz5S74pU9ajYWfE+OF5EraVyC3TJ69/hlbMCniNOvTM6JSe2pcXlZjdA+78+v
M0gcStPMHBzvLugZK4ycMcC6Ta434kG0u7hPMiskaGu0yp9cv24ql5w+P5fS2BEPlGNEIVqvniwX
IqMSXK94YlSM/71pq2D6lEVDwzJKRn2eaz0kn2Hp4pmA5uYGMa2kHc0Wcy+pxBdbxJD1Efnds9C/
I27ucKdBBsIRzgM6674C4rjTI01IBiMdMuwTOpv92tUfiQcCtFfXwGnEVqT09jEqOB4YV1zGjVvN
GFR1hU7cJT5gSHZZMU1RAzrMOchDiMbgqBo6ZIVeBszLcdXEnAM7qA4DBY76srftU/9lsaK5/cd2
gfaq+EffZZRyq3x7jY+aBFAhMnoLZNJ0hoU7N/p60YQ+7E0BQanVWCDQPvfSwrzEKKJHqBTJ+c54
lTVVMLz/1KMO5gu9dtQ5+Q6U156/IpbHT9DhQxkFgrGIMbaxBIFFXoFe4yF5UQiB6p77ixMDF7V/
F9bkZObs8JH9VW+pgEmwY/PsGy7VEbb7JOz02qMriUQjdic2vFLZQ6pxKfmKrdRjFvreBHPBbdtl
iLwWiwUpr00Y9uzwI8s1H5i6MLC3KhIb5wCfLR/igLiILWjL2WzbpiYdW8lDoMgLkpmQuMWUBhNb
0JQvRBY/LxP2lF93r808wHZ7lKDZEscmkt9BBts6Sq1Nzr7GNF2sPPdxA8kWe/W0tsojqpD0GchU
2O2qrfAGGruNucrA9lksGkPxEkRJnXChny9Wvd8c1jA1TBkuUzk/CatP2URUS3LXz0mRDazi6N5q
5bjRJhZn3DvZZdnxW5paq3PCeuj9PG3An/rpnTFfm7teKkAEVg0Zh/GEGK26RIHLUyzaO8YpkdLz
a2JvN6Bq6zfBJhECva+TGiPgpJqpYYlbZP741kNigOiDBtmM6q+YvtmXQOSGu+Zrkml8CwrI/4jo
tHPUBIkhz0EpSlMEQ5hkwkPnb4hdnCljTiUASvTX5Un9pQSziYjIIsIBu+pQMG3/UglMx5GuWmcO
tvYspyv4RVM2W2sPlMaWXrmpEMaODNGt/GgsJUD+MXnfiSL9C84OdnHUZpuWUJ2P+OAJRTxr+6r9
1FZvgVqY1d1Wq7dER5oh954deErBBHpEywvYuTJmJNjZgO9e8nAAoWAFlBIxAMpy9Op1hGvvx4NE
p03oTNIhb+j9Q7JevkcTuuGTqVZhe/ePK3ynmhDFcDPsVKwjnMLC25yMYm7cn8m1vFkjp/2Gbr8d
iGnvmezWi2tI1NguIlNYKw4Ynm4BMQD4gmiLiAKQfPm5VYrzfzcTVOQlzKlCZcUWQsjq17CcfAaY
abbtUyQFpbiRCkOAZfNEISTT7mikL9avPXZ8KduENuTuuPW7GxDKA8xZs/1AEVRgzLdh9/R0t9TE
CD8IRvbqS35dMpHuKWs/P7/ovKZSloTXqD2OxkYzARUoGstztWFX87SLembvgzjyeaFgnqRcuceH
rNcsk5rr/9x9xtxDqWyjhkH38chF9bvdGsx/h4IC/SktMS8qbeu4nJMeiV+UPG7k+R/WJBjqt13K
ig9Aquoi3e3ctKDjyMwokKVx7J79Ih6vQaylp0d8t9jHab9LNuyRaTKHrO2Ko06N+y5FR50feeHd
m9NVPxDX+t/PrB3iADPwP9awsiQiYZl/3rkLquydHK/rv3aFLI9AcfPIs0RGPor4uJ8fZ242qylo
ZkDfnGaGwdbuYbUQriOORtgb79qgDe0V38tFL0aCiXIsYIF0isV/jRAekmJU8FD13zFpx2OOlq/T
H0Hd3hW3zwHbgTPqonUK0KTAluECwX9qu0tCE+rpO6/dvcq/VMjrt9MBWApURE2H1NcqQQ9XLeRd
fpuocm24FMSVGXiVjSv4Ux+boS4/mDksbPZS0yfsbE7ryOwSgyDauSq7qChNBDEcEnKg9YZUgL3p
D5TQfVu8Rm3QLZR6cLX81o0DVp6/kr+QBa4adGTpf+fLfRJtrH+r+l3nKLdJOlpTUdJFSZd+PdIW
l/KPio2Z9MqJclVIXUDjW4edB5UEmtWgRS+d8MxxqGl8yo4nyzsGBEkqYMCwaTMPfvYA2s1cN16P
E7eHU8nTk/gyuQ4ygrMOF9p9Cb07IPlTiWXPQczMps0kUFA99LBPjXsKWs3vG/Q7VBnAX7bIT3Z9
TrqlFcKV1nKJgjEr+YkXs1XlEG+672xKAjpvy/dc4VkHMVAZJov7iyDRZo5c8o1WLxMAucgQRmqS
1uNjVqlN4fX0hQvhSnThpzqq8T/m3q6XUzYSALhtPIcQYyYtF4BWgz76l4dnoeCxBMTnaHnx4k+V
2xRtoeMGBubeilMYCdZSJ2BRwmk1zPU3H8V3hWB9c2J0xzrNrU2BKh0ypVootdlC5B+yXp8UVewc
ZEi+kkR5DYLXFT/XiDwMdwuJPKiFwRr949EGw3R7dPLIz6cm8P5YvNUhwO87I4VAda7gXdtMjcWZ
jxayL7SiQgl2spPBh73QTjlwexBe2mWNbz7RSD26MII3nbdX358OGsRpnEsQxqTWcmbv9RYrp1jB
Z7x71bepqeon8yVmAlY36g7D8ijuDbSO0YhWwxjs2JIyOgPGGeRKNbmk8mbf6v0I21o4IJ2cQi1k
aIQ51lrGP3Xgl3yQH2VYwBR/TtP1r3Nm5VpcrE3+zyTajpINc02EKKinTx2RXoStlk2rjcBvTMG4
VjChKW9tNtQHXG92w9bxjrSlxaE1NJG/4tbvqRwwipv2SUUR4aCpOLG0GymSF5q8U+wT1Qti96aE
uOKbEkJ5QkKHm8KfcN/c8cpGF6nS2hof2jD7P2FGIeYzHw0QGofzqF/ZTR8Y3TxOgYngoNIRp6e/
wBqk4cbrec+tSTx24W3FPSU9/rI7vVuTHumVf56x6c+gxVD6LDjGnC7zF1xjOIyCS9/nUSf/0fdx
3YLr3S07NA4uMAKr5g2MB2pYiQZGIKCzbR4vv/5CI/yIN++gCCLeIVdcv10wKnnF4moNtj/OVkl0
t33c+wJV5tlKyv/lL8xoCW0jdJ7k8PKz+Eku5OjmrfTMltIFs8HmtB52P+knjWKVcNgqq1OSB4K7
jihH0wghIWDuJ9kraYZv4Oaz1S0SGOJIRK/l5PEtHqyVyVZ4nVtQXdSoYTOZC6/hs2QFGI+ixyja
+GtZgSTuRzUYvuoFa1M1rbubw3ZbovZQRtOEuv/9ZpqeKcFut3sM7Cz1ZrQNDAm3cmCRKBKySOAW
tkY+CpXL5e7rqI7opkk8+/Q2ouKqHAK5dH+bkJ2jAsY2OXDrK1/PdJGytrav/MqcAvtvrCkj2+jG
c1hxFfwWg3lr7XADIPTBo2c0x6aMqG9EzWMj8YKs55PGp9j31N7eXwew0ycyJw0yWkLv/e/s88ap
m1hftsx5eQr3CRME7vf/HDk7haGIOynabO49P7rKi5XQAgOuP2g9r7+TZqdsjsURt16eXCXgnE+r
FWhri/gy3ypNz/ModYJ5DZJ/v+gKzS+fczAfdFNZHodiCLK5jXeLFl8WY6FdEAt3wO5Rv8a/4EC0
S75x8SWgC9fBbcPv5toh22JBNVckkLPHcsUYNVxXUghG+CjFL2IuUBOpWmcE0PePFXr/4dzCUDjO
AXioKW/clXPSdYj4/7Dc3E4H19cn+F8q0guUXCCxCfYRsknfcswQng4qwPM4Giz7Ol1xL+/QZiL3
ZwQVDjc/LvDlPcrRfm1FIbLLrdCqlrrhvtPFAMydyLE3ZByAL/vOxQY6WhmOqgF/kmMi4FsQcbTM
FjcmJKA1qBf2GGUTqx3uGP/o21pSOZiEVHZqC6T0DhpltG+5mlDQU4QaELo5cGqF+uZ9Wv6G7XVI
RXGQ+2h3IgiKfYyoGMu5ydAJx38WSQzH6v6QVolKvSHKVSuJ9MK1u4h5QgnLhjHRp7+0Q/+8lPy+
c9SfGPfeYcaOvj8YVlXPWAtom4S5pzIuMU7QiAkKNUL0MeC3U2FjtYqMUGFuOQdHJcj9wdnalGU1
8OKpOkEpEgY7Cr0IYUW9Ylj8LN7DqAcnjpPDl7g/BgQU3TkHrF2vM9rBMTrxNmgWSTyDnhWUDYNg
Pg0eKNDmwP+6KCRxdjiV4UtiYMIyXPRd5FtWA90v4bXGsgoGvkL6bKZPM0eDIpPHQmU3JUfdGWsd
LKsT7itVAuQRS7IWCWfiPUUsOdkqv/k7d3WGADuIrjQliQjm9j5UphW5qFrRrXzu7QXkbDWiKWbj
F4bGACH3soG434ir7376PfWbjLI/7exVx6/scaKZUflvkz/XeHCopw+8DYjAH7z07sW5G7eNW8yL
/fTiasnPjCmqy5EJ1xU7z+aIca0lzZ6L1cN9Pwwvh/ckbN37j39eXDzYsYFxXjR6uxZE1nuWpm9T
DJFf0MiOWwaoGSwuU/sXwKX4tp4IkWHtEW+HzXMza1Z7SURZokSM18p2S6LZuBfUwuwGTftmI4pI
wEdKDHuK3GwCKGgVXz0AGiswAKIFKeVDymkZ1ndY1z4FFsiA13gSJSuKA7miUADoc8QwZqk3i+QB
TgyS6l7N9W5/v6eucK/vR1WBpbANfK0r0TLd7mQ8mLmSMjzlQp/zcWr5z4Yy6OO3kfxIxCsTMHnx
d0H0ofh7RCm88FRuIwm6LVlDrRTwMHeoRnPHl+Q3K+0Ll946XBJ6ueRYePGJkU6VQhnXsDgeE7nR
wIngsx0yFNPZrpltQSLEYorU3l0miAQe3pWBy3dTOjSYN0eCX2JOGV2Y8IUpag2Dq5/dZvCPnheE
Kng9d9LPX4qnlWIlmzZGqXqa5tYZPbYKBdyZo8WOBZ0Q2tunPu8xi2AI4UOnRWTlHLFTbPuLrUh8
5kLPFtyGvo8f5qSSo33WiDZKPLgSFId6Y1r6MJK82rzrKpl2oQs1VdU6Y2qSXum7WeovUNI8iset
LDNpuX38bTOC+FpVZI/CHUF6HwdVONsrzun6ZnNsGp16BrIls+DhPBqtp/LRWMi5qMG/jGlGaCIL
3juwM2ShTNaf/frF5VAO7K5aax4kvGcCV0U34vYpwp44cQXO78YiaMVm6XiB57x6PwduhP8+1ofA
Yk3hceVZy6R8NkxLnB14ETWylZYwu6Ko5m+2GTUilXqFZlbZU7PvHgpsW1t99MOEQux9MHciD6e3
PDIglmh3JUfI5L2+2IYXIFRWWxBzpI09KzwiA5TSf2PqpSxZfJHmadWrPjlrusiKFs+GQL7cNIA+
Y2g0YVj1gcNYSLvGZkCQetY91dtLpBDKUeJzcrtMBQ2nWOrQF7ghTFjLa7hSmmIR8cIA2vGe/qng
ljpi73o+cow7BRfvzLolzOLXX8eh6U7LVw+zI9vTaIuDKSbkYpAdgYhREqycvOST3F+H8lUFKd6X
WmTwsAFY/rfgdnc1JxQ2aT0tQh6VQFBN4lZewLDg1GUVrqy1nElcwJLp4rtMiIW8+wV2HgOMWGrL
MHqQX906nSrXDp6zMQrYAjGpR54eK3yJ+12CYFWtEhJFAbuW+PFjPN0M56QOCCE0HLekukiNr8Wm
wYeBwudu7mgAF+fyL8Yl4MrBIR0R8EmR3XP0RZNGQRpuWgYv32PExsiUn7+GNJniY84t3UXPCknH
3HwRXHZmgjbn3zLskB4d9Uxu2OSwbM2I1zasNJY2tB/qGc6aMX2Y4Lz28EgPTT+PGHT8PFRtyLev
NABvSKfh6pWFYENtmCe/YF7VhgfMSDDCa9bg0t70PkkMYueWWMqLn0GVEYyvOBK5cMS2F21ql/Ja
c5zqS2uhhMJ1NmyyASUwkYnPQEYd4JdyTF9zdgpdLA6psC1wlqzKUB6ZSGUsFn0w2kZdGxrJ3gxc
gdKTbOcVKPSAlmH4iyAnbSjZqelaRTK3azAdgpSO/I7lRJC5ou4j2R+DxlSH38VkLIbMiMLBx2gj
ZdPPjPchmv9MHCSB/4nqkGw1I+tnweEEJZKEQ6IVRwLFIzb5Q3U8g3QBaJlaLPX+JIAuQZMiGrjH
Bi50wRE+edC+p63rwn/C/T3JSRKsoBp5NWZOYaeGJIR570AsP4ej7okG01fPOqVoWydwUKX7mvzm
q2fF0VaQS/mVbDaPVchtX1ZJw485XAULmzaq4j37ZAWnagcIl/CpBHCgsuzG23WpWnuKoJfY4N4o
c0nlJ7mH1oXFshmMwQPoMGTxsD2vMjLUY8ta7MuC24jV3vvTbz6eVvh8PtNOsPSjrxLlGXtVrN6d
uzrP5DQtrhmE+zPDHC0IVgiAhyF5DLr15XBVBOYMqs0FhJR4tJ3Zv7/hHyRhXyMJcLcFmChYFEUZ
fD8kFgOsjz6lljq4EA06WJZeo/uPaDNPSJTd0gCiUX2H53RRCsLs6xO3hgt1RUSfESi3GQy/y2YI
mf1jvShLhMNBuOXGDiVjQOEKtqc2t4HL2AjY0b1DkYpTIwmY2ut1a+4Eduz9eak7Y4YgZkrjnOGX
JgKH3LpG1k8Zt8nA8TwGBodZ/hRMJNxRG+fAQtPhu7knC5J2PoeKkMyhGeZcHG3ydSKzqtHyqXzF
OQsPhZakab22aHwv1gHbK0PVbThQh+vJLHa0vMKtqHSgQOQjdbByuxrMk6M2HlzH+jz8ZHySvGuY
74yT2y5ilEETnir9WZw/Zuv0ckiW6H/sGMmnBLKbfHNPyw1kc1ssTUlHuOT+yj9mwu0ggWJZ9qns
mvEge+qbk0U4T0+91GAVLO3/BaobpOEFlt99OjwoskJXyXqJbTrBQ+vVcHtfEBcyuwVg4ULIP4ZK
rWAVDTWxFBx0q1pLSxEPW7pnsNNtpPNf2pSH5gMEvkYIBHr37ruWgdJ3J3VlTOo/sb1lqWuZsv0C
+cMuL58GrjjZJY4i1oMIWAM+pMW4/reIoZj0kPz/VAVN2alPvpqrYYsuOcOnPrv71mp33w4yjndh
58iEM72P7ti5WhnwyDSh7zmFR8lQFRN/i91KirOW5Ede0UAVAzzSop8A0S96dTWDDpr5v5bDSinz
KO0QvONg76b3jTOGouptUdfMK2AGgkkEH22u056yFt0xQYaay948X75kxazs6UMwJMJE/5PyeqO2
nlK1GDnHzJPS51zmzLdD07ToV7O8pViLLS4UR2ylG0V1EOPZk7JiebkW5KZzb5mwOTq91NVWmzxv
AY9JyG+lq85oKbfxy6umzeVoHKc4/+pkLApm2SBb3r3H3qzJ51qjWBzaQchDVjJKtNkd3pPXCgIK
3eKQIVj3+T6U080ieBmW1rDYqTtvKmgRhnGdzu+vKuq4C5/RZwEfZckcMCZuHhpxA4qJqqCQRNRv
nW2IjuTeeF78fZTygzSF+BlAaHgluE04w23+ny/GccyaYK4lZLoJIaF0HE1NCJV0K1lUgeN90+pG
ywgx/47WhMsc6cNw8W9hAYUcHcHBgp7KA4Abvz49qNGYoZN5+eWKQV5TWM7zwrBg0kSVstCDSAAE
S1kaiOdegDp1mlkEmxNy5m51OguoJHgHUAp5ti6ecoG6RZ1kMgRzYDf4yddpXhA5b27xTdlxFBCo
HVOMHSv+ZYDScEJeREVjGY+m4SbZJhIiG5stdpLquLRL1H8glDoxaiJaJW9hDaYUP5SZSZjqkv5c
fo3htdylvLBa0f+eAx3Q/55hUKZXt2PZnOhLs+QG5yRNgySh4KKq1a+o51Dn/BngBMSN7b4wTLTw
SRVorfdODjuCw1DxIW37E23SHcXZvlq289PZKwBoPeb/kmuEdq/G7QhMl5Hj50kyHS/hl23ybq0i
wYBCYOo5Fa9q4X3UchkOQnXd8YQIdCzXpuBzN98EKwuJ+XTwEb/4RthLxId2BVy400jNhcKbhEZU
efYLZaqa1886/nViQ3UEetVk5Z/yCiA1Z/hHZnJX2760FjXKuJKQ4NGz5NbOrn0aIuHENG256CVY
OYJjApq98PDmYlPLvFt2eUA95o0+wuFlRBVTEXiq8r7xcBe8VCs5xSKICx2Oer4p+YMIyx1r42X4
ZuBYrlYojfeAstYLoSCYKnxD4f3sN+goFvaLAATskGb/rUpo5n9eBSkBBjZ4qHq3WQoZiF/45HUw
dJJrmyjKT5RVEG9TFd5wC5sXMzTSoz+BYmARk8sW5++CfjPKyc6riNoWOVir3rcv946d20tBmO2L
wnzOG5CK73NB8F7hFVsQOn5337h3FswDxKswHKB4njWsnFtiutnRW6b56QUbw2emZuk8tw/bcMp0
0/rmPx71O1B+DFrjCLlyzyqIEnRYFzSKXgQRcFC8hicBH4BNqwjq87iRWIRj7W1PjWB2QZsx/D/+
rQjlo/l/mrYva5R27YkkQ1hTPm76kqpfqYxMrf2H4uK2sn/2abslTIRCD8mZTGVVX34Q/GqTF0Be
NVirZ3d7XH2xGhixr16/+6pnfsqQvIylxhy7FH7mqN+fDPvFXu6+GGyDTPfJNvnHY7B+CkqNJB82
jm6lmV9dl0hxgcTBYdiZAqayZIG4nIHd+9EI47AQ/o4U+Y2sSMx7Ff1weUAjFmgVQz0POxj5QQ8J
u20LPKHfeBg8dHVoiuwQjuERyirRywCvNGAja65cDHaM1tCustg/KtbbXpV3jHXv0RpFizvPSNI0
A5lMkrU3WSnE1U7QZTwVtRyFmFshcXUmnrzBmN6m3JjvhlW5UYPJ3LegQoTMSS737iUYGHh4ft/Z
V66i106m8mTwVWw+5uVdNXEPgq+B62vt/BmNx3zsvhE0qjnb/0YFr+NMKoXAeFgwp56SNTDYAtUo
c7bAi1ikljsgzn1My5MBkcjmZkA6+wTjy7XAWIc5M9Lh+8eSLDHs4/svifW4aWD/xuF855P53vbu
wfFQDR24nN+Atl8rEZ8CeUy2wkEP7XL/+uk26pdMgT8VxO0tpU+4I7cpUiMvy1VKOqFCqscEBtNO
0/+aeG7ODFCC/aTJuw6ni2MF+3VzSN2blzgj6rrtBcIK8ziDcQKEd9rK33C0UszFFfn4VyY52ST1
/doaYdX7E6LXLqPTtTrl0o2jCkIG0G+TiM2/+8/7UQc0Rq3koe49251OU50aO68jc1Il4D16xHEg
CJWYH7cJYnNpFvPC8RJfwzFleyvcbmmQpNdEm3fgSfCQHyBlAsP5eO8gJ0rK9HNPBFsCDFo5ZiL0
xN/qmVx548Dqwe36Q1Hfh0Q4HnHV6Sq4+yh1aPTaeVEZr8wk88Bs8lBwiTh8bHDM0gt1EmZjKoKz
a6pryksDbniy3MASdFP4x3ZJkPaO+js92tDWtxALWEVYWjwTMgAuwL7kK8eDXHBdwD3q9ym47WHU
/UsUcKxJLtPLOsYMQY6AvSOcaIC+RSN0gk1XLSPwU8SZMskJpHtoZ/rA0kI4GzZyWIdUaQQVb4LU
R09lcZZuX0QRkUCzofjOWRm7xDM1ZMU0vka6BxUTHCDTkiCYYtXjIJiG+EsDN0cQOs+RdU16nxwu
2OjHF/wCllCNfg8PxGCBeIN6jaT4hTDB4FkZU+6YcBKX98ASC0+0v9ed/NQotea1s5DWemujNuTv
+geh4AR97HzpJVocG6n86f+XmES2H8AkzUFo/VpMadLRM/MlhhoblAdVIVtoG/g+2poLQxSQHW14
OlnGeWC/KJOeHuRdHImD5cTCcIHkuW8BfVPLHQFaCq6cOl4jrVPku/6Js7ea8X56UEHLKdjZotx4
LLQMVXQ+DjyJWO+r7V0CIIHWKIi+BN6wOkgJO3RwTNlKhrB1M3lrGfXZurZshYMbANwiNQr4+dB9
gM9K5xX895SZZibN/8n7kQigsa59gttPe7V7e42j2G5+BTP3ky1mtg2Jye93s7X6/ERvku+GebKP
JlLtD/LxP2UW5OLBJ+wUkKZxP7G5DHrn3DMSRN/+3SJzbzON5tBgcomw6NAWqIYFS3Z3T7g5//vK
WGYAtGXNNX9n76BBNVy8Z08S2eoNhGR5jDSZCI2/gBmhTwOJiUXmdIhp/r0O9VnqW6Kpe4BqK6Ym
fhdELPfXRWZ3Gc/2fdFS5n9aCn2Ai+KnTzCZ7DoBTauXLPnp3f7ppQ8+jai9k3ioPsw6RYpuxgAR
BKUPUGkxK/WAYZdACc8l3p1VRe3W3h3uxMwYaQgXdym+4t1bvZ9tu8QEzaGJcnaqFF0fjqIZnl7a
d6wM5f1S2BIy61/X7P4iDIXvg8EO/QmzTmVQGZUa5IMMiINv9+uyxWA57tOOTIjLeTPIU//kDmQx
ciV2LKO2b2gJpdn+Ib+YhgUBJ3FXhdRx+hf/3hs1UnQ9BbE9ujIe0xogrbq6sAtyye4InW4LKqjK
V4nVWwFfLwhCzST6DLEH7VyUM9rqgMEI3tkDZjdcaA7PMmKXa1JY6jq86SQqUMi4jE/1fr9zuB/L
cglI6YEjwhrbiWMQyJgtba8A2o7XZMW/HyTP7gQXf6EUiKkyflQhldXouH4JZqMuRiBOPuo44t4f
b2nmwA7kRH5S8ldKQfJmg7P6YJdtmJp6cbh9W6CAM3ji5rxViqbXgJHrdg1zyRbIbsdAS5t66FRZ
Q4xNf2hnxm4oKSrg0rZHKZG+r9LBK26ihaHft0RVpklEyl3xJGN46Z8Ws00CzPt2pkpdgEzUMlUL
uIeMEbs5/FcdDn26Js0C6I0HJB/voR86LN6XWDyKUbECWhlSDqqk9i9u6nyrBmgzdfBs+H20GeWR
VF838Jd/ODryIQB4jQFoJnvjaZCV2Xa+Ny9agH8F96Thsqxug7I261SL/zijtEuQn2oCjBlfhpn+
kBvZNJJDKlo5xTcUdwHp1l/YbX4iYUvQTHLD/8iIXB7PUItFa4zi5cxW6KmXb6u/S5jGQaC5fCV0
mB64nvm8MJ8n766cxqgI1EloIiVXZRB2mHzeXB76+CNtiB6QG4jwrP9BilfTrcxM/4cDhwubUl9v
uDEIoFkccyepvMCuXhw0Bmg2JENFnAQZLjUmc057n5cJPqLI2mPyTJpLEXDiAnZLKfr7Nfll92SN
G1I2QkqZJij8jSqYpdhJUE5hidtddOfTut0ZX1uTWC0IEh08gZeXL6Lors+gmRKyGo81ucMLdrdA
/DsKb3s79oU2qVkJ+dwJt4N68D2YlrysZH1DRTXRRg1prTreExrFg1W84+I/Kb/Ahe7zKWtY3pPF
OPbVnt7q6dqfxjiwftM/6iVUyhK+wZBBre5CBsy+xfPGFh7T1CzZbkEHiiNpyzCtMq+kAVU02ZNI
DWpf9ODYc8DmwikIjN38zzqJHD6y+zjt0RYVYwNbi2BilnxfCHFdKRwzxDz7eKr1zU4AzOTa8qJQ
JqPQ6NKAi4uzEeX0dr57Mcio/S0gM+WQB89qVJo0GnneSrNbGcn7Pyrl10nRvY1YqYba6jfyxx/E
37WdGSXggRGGV7cDZ3gGicHOETTx7GCLx9A9l6VB90y59FWPpfGzTg9AbVsTBfeLNCbgig1w5x9Y
lToesWPyD6SS94ozRdIjFdIAgVdwLuW7486UIvvu9OOYYrkuqD5QndKIs6DTEIzRcHlL7QJKYCFf
3Mar+PFSBcXPxnlMzGnd+UInR9AfEWjCOifnvVQcvBLl0bJW8jG/mm49JH5wkaSOX9x3itBiVxwI
uaLQeX9uhw+LbJ/6XCM7SSBIurLk2/yeLg9Mgt3Tijs3OBzhesmawV0lLRefDPZXQDFW0jPPwJm9
4fbks37ZZz/DXhD+ubuy9qtFO5DqjOOSQq8kXj2D+CpBVKrnEhWKkJgEcbYHK9SKOdSllAGm4LQK
r20QZ1kEC/qAfuHyjgWgJy1Ks4InQwVsbVoKxiKI0Z2PcbpSiPsvrMz5yOezAj6EN5JTJjKZHRBy
LgJw30poHkEELiOCPaW3mIwPgBAFu/Z7+eQCvflJg32mFQQSQKVBHo/HxEi4aYExiYqFWWPXham9
SuxC12bQmdtoRcS1ayL/+1U4UVAOsPMzWYMk73AqtgL2GaTALYU6U21QE9A5mhdl+wP7E2vO6L89
lDnbHvs5TKiAXxsMZEsb36IGX0bfvPZoiqLbsOci116Sy446XzBobZOS5DvUItf5jUa+9Jvrk/6g
AnfEPKKv1FxzYYvLjmwIVexGFdGYKIpD3MmCcBgZK18A2VXKmyvvhar7uMkrvac6Pf1XUKO56brP
W8yOA9PTjPPBsdnSmCvWiUs2LXOXwaJ/bwAehVPwmVxGRpWfxH8Jm+CSDa5mjWy2sr559S7sxtDF
YLDZ+/co3+OSQNAyC3cM7gncTBq2/Svmw1TXksVwBkhEPoYy0EUdYto1TcrX8/nDt5kPvGoFPikq
244qrA8FftfYiGvALQ/BSxonRsvp46El9yVR2pdaPgxwZTdZDKpDqwSFqk/lnhe3rpXKRz2F4L9L
UtqoNLx5osNMd/aMCr0NyRDiE2FHohHS4EgiCUbGpcc7uO1PyXkWJVrIpKf/dLC1OYbPU9KM4NV2
CIFhK+UrfBtRMd6dZQ8l9yAQVK6VpKCkkmz77S2cRVsekFTpIEm2l6bvVi959Hb1Z+lIAymSxQjJ
wTo6ERKsptO+xGYhaQE39rsTMe9q1v3VuJ6MCDhvoxPcSANesZ43yeglIVFcd/68Xqcf1hmlw/v1
bYddtFWGQLZnRy9wKepSCFYqZmUhYP+NxSmS6Sn6X2vVlamddrsmSz1VT7vnfwjzXo+3S/2vsJEZ
inCiQqOqNg4upGbgcJwKfrUucfbmxtKFieJjwRxHNpJ0hARnWa+3Zf2h3QBYMpWhLuvhf+Br+eq4
lyZ6aLcqlp4WEEkAZelBeXJalsFGpAE2Hm4kUrMYD2Dn+YJOSKgEze/emOrkk9SmnDU82b2GrI6j
3NVF1CS2U8ZHeJsXFT8DwdPW1LUuvcfwO3ZwALM78rzX2nKJXiD2E7DXuuQBG5YlEhHFHV9A/ruy
6Qv4WGLcit20BG3mEXBA2FXPK98MSeR+nmXvDQsscK8PnGaHWkGDCQVxEIBmHc9NuYyLjOYJ6ZL3
gFCCeFdzkRTx6y4YvhWe+WFoWnkWd1tGOwbloCOmwhbWxvl9obdUqyMPwSFfR62CqtzXek+6rBE8
ILierALk2N02SYT8I0QmYs2CYC860NP0STBglC1elbyUtjXoBVkZPK+vr1HOEW6Yp6Fn+ajMNWmD
rXqF/YqJus2U1Zv5fnGJ7GMjpmCKnW7jDqDpVwHJw0eO3ris1WjdYtG8PP4oVVcSB0S+qRlmVq8y
T2iwqnozpBqpCLKdYAHxLjT9xgZMZaiTpyJV2n4z7dHA8mOSUqaLznW5r6mvD3A/ll8K95h4TPlF
XGJ0yKffjUVS7WZftfp8lk1PQgut4n1Y9KleWZguHsvV4oUyWy3ENQz/BeTzNVzhL9zRQGFTexwP
cdlx+dDN4fG69a1+l/Y1kAiMe9x1jRU6DhxcXmIrFv68YvKB4TsVEpHpQIlOHgXKzDDl7sYraUvs
1jmi9MlOwVZheMzCC1Dczh7VF0dXt9OaiOoHqZBertaGKs3MPi+LyhGn730futsiKoQNl8P0+N20
hanJgOJiJP80hy4Em7Xtf8atxWVnnxvPGJAq/1rQ8gttrYCrcwKVwSUlCuL19LcfsGVKccT3v7T4
R23kvNpxE+wMxfAUUGAWjQSC9/X7ePfLKS1zirCCkr9OgzC9W1BDO95Vw5IC3qEN4+sV7N1ngoog
qPLcvlOeV9D3bbiEdUOHZUchtF5kEvvAH4aUoK6vqpqoD7Z6Vx6QBtDXIApkHI50VReBdfiEnNYB
f9V90zu4uuB2O8T0IW7KyeUOXOczpxailY82LHH2NOwkngMIlk7vN/dtgjHwG9NMxea8MQTUY97y
0G7RoB0RVe3/jwT5zBnDa7yCONMhA98VerjvI4pRZ68qk+ZcpVKoUEohtMisdn+pqWzoAlnhD5dU
L6k1bNBREGg/YipKCB5SFxvgmwJpIUeNJUAco/bZHFbTN+jYS5L1wTvhIoQ5Yb4o+hgAwj9dt4jJ
akiDoBthl3kuOCUJObhZIT898Fk0VC4tfTcEWNDE1mm53wfoGQXLR7Z3VqYk3/FHerrfLxEizIFL
vTzmlkn0SwvL7I9IaOnVIp0uQBDujl5LwWb83a/WiktTC9HMfTn6YEEQHtRByAvdYCGLQsbX7kab
Wp7Pv5OtsnpPuKwybCHeEVqMqHzY/HNlTknJll50eDU31Num8Rqw4L9eZvtLi8uDL8/Jb8kvPL51
JvQaqtCdJNsUsh3hZXQOgATseggCZcbP997/03L1WyRmDpqlx7C/n6GUESYhe6LHaLZ9H4YcWCfm
LLGc8qZdg8Z0V2JjpaOh+N1CaxwMq0mjJJFIAmTImy3usqeklis6a/HrOejj8635Cd8ybn0gqDW7
nGqHVoLFIvEkuC8bop0EE4VR9xArTGtBDPko3JwBQ//ndju8kG8P5O240lcqYpRnmfB9yuUf3IsW
zfXLHqvgWaSHgwkaARhpxeLXLemomsuteCHZ1QTq2Lgt1yffr/EilKargU1pyJZI53TSZG008C4+
GMmt7me36ZshWRp4dCwxN+BvQHDlm3GXDCwm9RcAWZMKDZ40MVEtCow8n7zHkMBVTRXNZ64AXrKu
4YZE5b57hBizojUSAe/KtAHOMwP1ZaFLVd/GJFwpnu1+IbgDTbZk762mALbTY7UTvLZFjUaVs4VD
sDmlkEbl95SN6+VwDHU5c5NyHtA1HiC3wj59a32Tuu+BEoeDBgvEyy6Mzy5+a5bwkhk/aECzfOxV
vMcC4LmHMCL1PZj3Et7sYn4D0YEa0U8xNOFpK7NASIVfnK1+aCLO46qElBxNfInvKp8oPLyOuy9p
1/qfQtwUijg/Y7ZagHy51mBEBYm6yNRDm3iLoik1UmpUOt50Yuna1KX8+bptFhdpEpdWdb5+ZcSn
/tD0d6LPtQVncAButAfTanCRw4Pg1k6SFDCl7FCqa7xk/FZmxBoOxxiaiFOihS7zEjsYv66JdkM2
hQNq5yCUtN8ev6huiTX7HLEDFpf0nHRe+6Z3UfXMkeEJDb4a60KydpEYwic+929CM2cPGv3eg5Z8
V3BKiAgeRfbbyqBhrG5egPnsh2a0GiUdkPMfjARrcG0c23P43AIK6TRPYhY8KA7LCX+3Ulw4zhPF
TP0t4c5d6IDp8rVhpF1Kr5f6uP9SEX/o7q5Sqo65JpFu7skdzGY9Vq5lswsfm5tdP8TYrU0UM4gk
tDeu2n4G/Jz+fo1Gkww/2xByOu3NoIlIuI0jT1hCkOW/7uluRTBRFeWeEZ861DvBNYbHx1iAEuWu
WnbWE+kNqG74yLRXe3iS1fX5GdJbF93bkRvFZeZKWGO0DW34pVqDyiyRDFPnM/7DfvOKhiQMYwNt
qNDK4PKzs0hH2Dxf9rWgvDBhL32L2SlKs8LDk6Hfhywy5p18bk6iywyQ4ZY4E1VYICe0uR6a3AdU
CzAoRnyjtc5uj6isQJ8/pOkl30CO/tIiaNl0XPaZvQEl2Q+PBzJnPI8D2tbgvgIS5Hx4Izhcipzi
NtGYziVetI91xk21GUm/FVxo9MJ1pS4phFeU7P++IULI354mDTDnmsQG2WFOOi4ekU+VxwoKHpaw
Wn/Fu85zBwHiMvtOMIGrgQiCj/KZ/QpDLDVyyhvVPqs77KmMniGuPwKwZFkMXlcB1EGAuoBi3W+I
H+HzMo8h44VCyL0bBt7M8/3Nn56+DOw80Hno6qzh3XIYIg139YGKUgQ4kEoDSSK3Ku9gOmGd0FRj
BTtGck+LxIjWDQG9KS32GMAvgoGMnUn7gjY7A2YWhOv+ohwYwbgRKh8zGmvrhFXXGZWqut3cGdGt
bxkQ4LjwYOWazyibggfawQYJtiBQiWl2jBWHQv31554xvlevNmq9LAFy5oGLBvmrUFRe+2ob1Rtk
c9VizCvYCb4IpEGQJs6Qa/3uzSMOnZhLzijLzFOOxYu+JnWcDv4fcI9gJ8kGss0AzvDn99FymVcD
aogsqHRdUHXMvPoeruCTl45vpujbcySlJ9hCMMUQeVsRFqWmR7Lx/CfxKxrZqdL8E8dgt/nVmKiz
gvurTomR9dSaeioURuUSSXHVxTMPEQ6Zu7Xb0r8WIeTppQLNp6lWzAHZuAPZXxsyPne2UelHyGTy
lj1HM957oqpEmJWmUae6GdciNW22H5uuLrTizzuJ5d+c5gm0yVcAXj/7o7AB991bF04BZchIPUoB
/J3lUaauBuI+mOwiivAVPUE+Q5X4NmzCzSEXf3YGmIAJzo77V1OvgdTUlFSeMYvgxl14rCPjJLdo
oRcIW7UyQwK3blKQ3Gxj40FGepKpuk4RngJYNwFNOdnmF2xMARCf4d5p2nMgFOy7x75Uf6zxTg4R
Bt7FSxFPNniwvg/c3OV+YzUSfvlu+MEGbhY1YGv6yT1fOLhL9MxtvR2hIcrvM4EBKEYpcHHaU34c
Wg7hUQx4P5ce1ywIisBA7Tu1WACi2jIrtplJJObs66DeERhQaR1srRg9j4/KveAPL4DU2djC6ugj
oiTVVaAeoSchZY5KkNVM43GconynbNWB8dx0tW6+OxG3pCqNCWn57+KGGwl7Yv98VnRfg4ROx+Ph
34GQTyrdpDjdP102UdGfDFKVeCmIBCNWsA9wHNouV1wBlIBJEDnNPwDQcXdKH57Sxirs0A4dHpc/
vv9vF9niHiZqVC0v/izhZlFO3lr1FZSkYCI5bLtee8cR514pqp69mTTXAi6/6glZrCiF70Geqypw
dBNxIPyCwdBVgohdC+/2UTGxr5xkxpvgTM/2Yj/XSyWDs8DJEC50/C3Cdo18P9WfeRZu8LWiwnmf
NqwRbWUXHNuAApQSuoVFb5HeVCXA4ldfnLb5skblrVTdxvbu9kl/xNfacjxbLHn47eVZ59XXSea9
owjb6J0jMqJkUybw9O5ydjivM2r/0D/RmLroT8roGRiA7Gfmk4GAE44bKzr/pVW5ZgQdJR97icBl
P32+VohNpDT5GPnTUK5A8IOvHxaTptosdFaD01JWInNb1pAydbrr3BNXeioOmQtcvm6b4guE+fjd
ieWYBxT2J98F2++XyY2L2yBCxFKuPjVY5uu3dNnSpK4hMR/8oLBiFYsPtHXdZZ82byDV+ayNRQiu
VKYnyYLW7GwU33nvQRjJEsbvVlGNoyNFl32Ez6Wfiq0Rw/LA8+V4CpFvlzxrX67I9nPf6idNs7Hj
w97NgcQwMRLM5MHoSZ3haVJKcXCd102SfHYU4u6h9/XgXfcH7COrBmPJblRKOW+vnDV7P9p71Hea
jl5Sh4vzwx3q4NeWDBjLvC7AwhnKHi5DP/lkLiUQ9irahF8DK6lz+M/3RtW956dnsZU/VoHG6rKr
NtG+gWZxkf46a9hG4bYtTbXFVkbnsU9a1L5mJjeUOY9DyeTNRjm6lLn7KosllRB4jHCGHq2qgHJg
AQwM5KHQH2qmBflFnRpPeRCPbrQp5uVVsqVhXc04ugBrKSwUVgnyIuXOjKKYp67+p7JobJ/F+7tX
hC9BfRpNQO6HNuSyozbnc9h/V3e8d7FdhZpeQEYBn1my92/jCB2+YIsrJkTaTDKpt9deHk/hASL9
kHlvoHF+87wOjRV5fRJVP974D50zwwfLF6puGE7c0OzgFcRzQIrIWITMfMPPa86evw615iZKqMKj
7wF3V91oAMuTjgeB8TPEutkK3hgB+LvIaSSW+Smur7gtXPWeS4ypGxj6ecuHWB6s4BNntQ4SflpG
dKCuyOYINmeM0nScnsMnYybxNFXAklWHVEKTRmg6k8L0LEAVVi5M71scVDP3bwq6R7YNXSsVAzex
TzpknPsX8FNftDaOby6BZvu+h/z+zysxxlNOe9fzXBvQOP4fthuv8xCHFsx04vyJGOJ0N5js8AI1
XDbOHprhu3RLeyZgFrPV+wYfB7EXlHpGNvfA7MagL2SS2ZVXsRl9ZrIJfE4vYXkmS+5g6aiMnUvz
Hwc0SM87yiuEzDiFXbzIMBxtGW5KEdeIDP1SbSD9IXIgbR6ap0qbE5ddckbfwCuxEB8sYoEKKuzn
KLrBfeB0P+UFiU5nVFQf2IJTi1eafkS0hWA0Zl72xYXs32SqmUiv7WujJCMiQbq5YFPxWxU/2smF
j24+nAm4fhI2+jLLcidmeEZ6r9iYuaDve6UtNJFQ53tMwNX904XCznVT4tjln4cbRYoOsd7FWTyA
V6tXSnNG+RPrD7KgiEu6krwQ2PNJqF26uhojtaXvi7UHsdlOGUacPfFb93C2EfLrcXhRtn4ZQ2Ct
YzEL9BTaIPAILVUKUZdhkdMzNRx0SaZ+JpUjC80IpZj4PLMhp60VGDc0kb38ozxEvkiTIpCdST4Z
k76cysMNIHZqvbVDqbfuFyf0Hxg5OO4XC8rLX1NbuhEGpZQDhPF5bvTGXItehbCFzyFz4/lpSLjb
yiVNZTY6hDlSB8iDUPhjmyUhiSeaAsmXbkP9sYTMrZt9ZOSShsZx2QGTANNWzIBGF2g3tHdk+tmM
ykLK6aWiqMzAeQb8/PjobGWM77navjOOP38mrEVBUfau2ZNRWPHXzRE43P/8J3qjR5u/A1zVBu0E
HSqDzbD3xwd0ph8uR/0yo0xcvJI+puf6eEUJp1yzZFzEUlS/z8LK2HHR4qKvwIw5obPsq0VMSRXa
Ukbr6mZam3+XRHFC2tnSXHCdgujvNiML/OYe8kpbhC8V0kZJIH2pQ9LuGmFLESmPlUuBSz92KWbZ
h0LdqzzHOKYyKeRpY1XpECIXUHorEvN6oQYI5KRz3DZPWQtfSmdPM9xe7Cu36/yvL/gQ73DB/fK3
dcimf9st7DJLahKQuiTQZ4Kz+DYjbpYLCAoGKpXsOdgvE3iXO4+fGVQPWq1NQ7fvHRbigEbHozUs
pJFJ11g2TVnsvQ6NPZgHArTqcY/r3Qb3jHZwwZsaTCJXI4p3cs254KANb99ZOWq1tsopy4M5Mgye
ANk4siKYnyIOIQokynxgPkqfwVFaXT9DQ+d6/oSOGyfKHq9mZwmGubPtvJ+swRyKsAJVQlgQT5Qb
0qBEXWc2g0JJ0WLyc6H9kkRVAj+jqeuoLeSRe4qUqvQA8kGiCxXufRNEpoBvSHj0iySEQmirDks0
Hcn37685xNhT3mA1rfLD+8Hn1FvGUU8EtpyGgU7O7TcHt2U7E7Fw3uJ4sYnf68tqPn3PLAga6mbN
i5AWsInPnuFRABEVv6IAfnV0TZj4nLnDy9E/sp4HbJ43cSmzuLKoSA0QVpheto9qNfT5g6pigHFr
QnjgIFPMCG2wPPfpoAnIxDjM+7l2zHaYAipWm0MNDXOJb80+PjgCGxZZv2BbmSLyMoohwpEVaMDG
bO/xa4sp3klUdGJ8Bb+gmmhwVmcJJKNSDXKEmhz0IZ6FYvQ4iP8ELzGM2NKMMX21ZqDH/nMkOJG1
8f8P9BD4ZDsmUKAekEnQnw8FIHjq5js3A/Tcr5VozKN3Ec7RiKhKwZyns8Npeb6H6upOwtAbZooD
pnTYmEUCHnmyxXY1yoi8RqmtJdDEU1LnAC1qvJed3oOabcz44FOV40Oaexy/5/YnoBzwZKXL3PTf
aHPYnIdf/6rwjdd3y5iA+EMlqPAsu6SWSljz2mvLqp8bnlnJmCv+8AyYKRdraKcm9Xhddvcrpn4c
zFY9zL3ep0zFj8cE8ULAZIL342S8OjakG+tkoZdqaEWvhstGZhPXSKk9yX4JNQMhFjllCT74fCq5
bizlTazqLMbfYVOGxUIxEgQ3OZN7C3YWrXCOFXM9joOXpwtAc+5i2Tmo9MxVvHq0ld80eXwIPrpV
m7q8u0XRJ9un3bPbvu9ou9GDzLBY/OPt7NYegzuMfdQa06PmEbSbBwBi9YUdg+MWZkU3lceibgog
U8XpQeI9MMdm/4QN5kpTj0AMK8ct2hDVUlNv0wNf0iuANtZYA4I4fnWAtGEjZfJU5ORdFIB79/2L
Hg9i6fo/LzYN2ZHkXoTGDZhPdnqMeV7iC7JA9MvjkTGp+wqSJHDt8H8g09RV1rPQA0AOoQ1qh/Zv
I/A1YZrUM5WK09AUU4aZeoKxIgUuz43ZLrwCDND5BhsxsNbkou/+xbAMFgcsk/4O0l/uVMtasxFL
vQUbBB6do54viiCJ59Ik74s7xrp9yUMPZf/JrXkx6tucIqi6TWkyIqZgfLRrFcId34Uwu4xqiKKs
d1QYFSr8jgPxA/TNB/3B+/0FzuZXRSzNx8kIIgDyzSE6+P8ykbOavf+aw7qu+FFWCkwOBfyO+dMf
RNNo9twcT73HSh2Jew78gwLS2AAYwc/RCU+xUg3SDZWAt4vI7hLXpNcPdZKuYaEKn8Q5Nf5r7hUc
rcig8YRq6TYZ6xpC8h9cSCnUDPdslj40K8UCZ5xT6FxnVpMnWeeujXy0QiJ+VfUvEfwFa0BN4GJt
gDrA8CrX4qosjvlegcTkrYBpy/GX42wfN0RrU0fZ91kTSaDjHE2aKeZqJJBqvuLvOUqMW/eo/SEZ
ORZTSYPcn5Eyb06bB0CBl1F6JAIWJaTWoDDhXbsNVZ68zogVlKfRpi6BeUgzbAPEmtfbGXjfCrQT
GaOuXO5IQv6kzQt52u0GcuxEsZd/Bu5Iql6AmNxIITXyGj9BVtVsnmxION3dfdZrLSnd5wnSEIWs
hlMPco910ebUo0fsR6KO3q7i0djW8SpkAinVL9EX8DqCzYemb/Tg6/vCuqOXi6DklEmhQW84FTLQ
8rue7OiT8u4w0cceU3SgGWdptr6+zduMRL4GEuBl/oeiBBows/RnjgBzbggAvkWAwNZJa2Q0FTyc
ONEfulJ3oFivx9X8gGTT2w1Iv41hT/pC702ca7aztlWpMLLjyu9gvIsOHmyvXy+huzRAeMVBY1j/
cDUkSCED3wjPwWCsrcJCi5tpnNfy5VXmfgg7BLww1RHpg5Ks/3eyJaQSLrCNAfHNJjYyBUG/N2kk
7yt+43/cgMvHhhDOZc1DNOB0CfjBUM2HHMsqJbvOOingDM6vfPWjwZmWvz9VI+V+HshS74ApVvQK
KNeqozMqJV0E6G4mq11XpRWFbx+KDbl4ikxDVJz7w/XdObM1ELGrxDOXLr7cXaji9ITNCJjKkK/u
hNu+7d+Qi6e3hS/vTe9EWsbaKtI71TIKINHjI3zm2VlZ5fMbY0fftY/ADn8SUGlofnwW8OdFDiMA
BmBwoGcFK58ZrltJlvQ5Down8eC8fMV2BSn7C4O/TEUoXXn8TIMYYIkhpzwMdG/NiwJkPEL8jDaZ
gs+kqg7tNBBMZp6IFPp7W4FcVr1h5NkXfzOI13JSiMjjv6dneIl7G0Sb5A+H/zXi8g4FG+al6pHf
q54buuLVwSlG3ShU3mNaJruOzYdgDbxhyq7qxT44d206sNesPm4V3dZSxQxowMSKa3CXlCvEKeLH
2XpI4lO89ICfpAOPpNHo6cjCEJqee7XL3Drg2OsbI4UyjgB4ZW+lnDfADOPwS47NkQ/JWm0h9xnZ
LUV4Ilb+X7QiPxzpHy5AN74tRq+ZsPvKYaCLycLp6xx66XS5eHaVnDxkxtT7yVbOvdhcoqIKLIvg
4AGJmPLYwCcciHjTQKXwIKUCML8FHLKdXVLfwnXW0F1JQhyV9ZckL6214xFXBbzi1RPzUDQlarLH
NZo5ur3pODv/V/hyrW+L6sguausAL3ucy1HwebZfhQeEsRQ194QvZDq8m5RkaKZx2R+pLWBYzkJd
XYriu719tNozsGYZAg9DYHngtKeY5th64JF7fR7t1As/MPAafXZLbb96YEVI3VKlW9yUM2AMFxR2
04+bX5ZskFnNWKz9SXOmDoDOJYsBjoBl14L7QRXm0GG+QUxllC48gH+P4w2A4sS3TfNxALk4EyKp
JnCp97n49tZHFhcBVnAIy5VCdO1Fsblmkg2WVgYoKKZ3G1OtfU90H7A9dIpQ8Swbv8SdxnaScDDG
twag4MmFcn/oCdXZopyAKs02zF9L33zIs9DeTdJLEV7W9aDHgfKazOuD8y4QYM6iNFI/8e4iaugQ
e62nTD5D4gtpu3xMO0u3wckb0WJB9MT4pukRc6DGCBuUMAFfMFhtbfQ0knTcSLBEt9e+lesT4Zjz
AyaT5StDWk9ubM72oq1awXrFgecKrXNXuDKHHfgWt8B3Gt7xxAWIcWwA//8zQ3798OkSanDx7PBZ
wIq7RzDV8Mmm83Ng7EJIqnrqjhLuxSqo9Pq2G/p3PyCTHVYHMtOP246PCGtbnveTefXeeUckH4D9
M7WaOL39rUx1qnOyDZhF3uQ+yMNRQCgH3ndsCwb1WGtVwXzBx49Yf6rDF4nHc3tkX5u0rygfkrY5
Wv3RAkoBWUBY2Ur+inpN+JmPnqyaRIT3wYTq3d1YZUiK/jdwkogZ9KmrtE3XOOHA+eWgYNqcUThR
apGsWTyEgS9V2HOtgO1XHHiEON3G4sPrrDqoaoW2RuZabPOs3H8pXzGKGU1qPALv84qLi7F9qgXb
5I5APjml/1MAIfjunmZBqNnM32QdgwELPP45X4BHdee0CIWep769fwZtRKggG6qh8sut4LPQ7hZU
wrRnMVSO8bHxJyP9zxrhZ4inWKaa8Re3Nq+Uol2gkhRwBZRo+6xpZwFbmaVAUuOGXGSNeMPrKfej
aTaVwewuX16HzmjQ+NB/YzGUfk3qOcu7QkphttXd0V7iFal8zkczbxsSY6jOpFondTH+aSf++rdK
toJpcYyno6wjh/Gjj7AW0dVr5rkDnTMJ96xn2EswQnZxS7E/7aF2kCciY2a4Y79q3+A40ilUr+2j
l8stCm/n8sQL3iWd/RyOS4cZY5AvPXnctCW5c+BVBrfhihCbGNI5E8kMI8libxXizUIq37vQT3up
ET3mK1jZhroDNHdnocCJe6eYGaraqs94omSIKcnGxI8x6FXqjLWnqiUOZPYY2CPoHFbWZ+dYFo3F
hSbVkCUVqwxdyPy7oo1qrjdhyNXebHCrEzfFVvFFR7R9uVZgBRmoK6r4vlYIwHu6tpth7AvwBMwD
detjfdLqldzdyyGkQI2LWTeYOZiWZu3LJI7CC5D2MkrNa0Mx9Zp+F6OLLwdpIQLQqh+HPZJrA1jY
jDzjhd2if2jferKvjUDZLXDDMVolrl1idmCweo6PPCXEMmVblui28ikbzIop77jXMh0ZWnQwqsdg
cXxTGrO4eWn/WW/Sq3MU/FILkoZ86MPx+n4U4jE44xkaCKb6sSs06r2qwSsviLet34lFH1ZFp4Mf
XSwE2KlK+f0dTrPlEWU9ILtrjFYT7snkgQEjMCSbgrDkncghrOCYOkS8AloP/xd7YKsD89b4o0AC
asgZGuXNy7s0/GwcDw/YhYoJ3RetZyrukylwUAqki0ZRMiMq0wDzN8opMhEF1CeHB7sulOCc3MpG
TaTLTfJnHhVJPztuMSp15sVNCm7YNCgwnhVajUEtrUzlnWkVJmkHsCbyns33YXcAan2WppqTGqC9
05gBpbQKidQUtMCJHTCG66HMLLmYDj2b5vbnboGSJtxFLJDwcKMsXruQ/r5oq+TOZq9Dd7l/PoDw
0vod7494NUv0PNR4y9OpDEp3m133NQiUlwwnw3ng71cPzq2xvaAByuxa39Os/NSyw0yczb/RQR5f
9yITZh0FC7kXM4EalozSQbIGqs9D84FmybU8haUktku9jR3o5zPgmC/VsEQT7dtb+CIk45GJg5vi
T76dujf5oUVyHCivpqruWKG+yNsWuNUoCzRTET1xeFZM28Y3Af4fy0SbMf08IlscnxkOIwuSOn8A
a3JelTRHi5N7x4TgzSJR+IjlzX0tlWplMz5IDRqghNXVkTpetPLmlWnzVXJwALx7EkIW4Xipg0Kg
7LStpXiaKs5osDmjSv3meJDCvzz/TsKAMiLGmAWjUOdZ0d6WI32ilUV3jwYBnuugxk8s1djR72LF
EHbizqRDgW2696Q2FkYS09FDx3vd7uXbqYPK8jenN46fc/bKQ5vrGwhNf8VBnAU0EpKPxb/aHFJ2
ZHODf+9Drhs1z+BFerKQS+3Ho1oNRuA07yAlxFYBVksEaUOtO8ynoTQkqlKn+IsC3Om/fYqNUcgw
thrKi+1ZbnOdjNunm30mbF7WsVP7i1axvH+Kevfe2m18/M40oVTnqj8O3gfdzxHcDJoKP7lmIPI5
/rfyyEp5NTNcb6LIIsgxdKNQNO+cdOemRyEVHgGD9wy+rF7fMQKel+KH6gdZehLjYkKuENGse19u
/QOCCam1J8wNScOSzSmpD9BLy8FjU+u5wNz53IPv5NO2Vn3jwCB79B85dwwStD7UC0lbyKPaJW5k
UlIgug5jH8fYF6tzr1qOGqSq1lHCfQRoq4wGqXGtRDah+rmzb5odUmjZeB+kq7QGJFyhh+pzt8+2
6SFlfP7/hGiWZE5H2izn/MKAvNJAMUWL9/vXxKb+Ei4iIlZAt/WlS7oxlj5XI7e0Fkahg5Vf+ADf
6lEvO5hcZnOni5yS99OIEe9vzkCF8RErBI5OyMUxM5LO1Y6qGr404a6BNrwnl3olcgerpzabTo5h
oYupH75C6jt/mDxwVea3Fq/fzdI231b6Uxe+J4Y14Hsa1BcQ5LMEB18Sf5IrxqiiJ8vfFVQImTlr
+K+CFyBYdwtq/T+VvfsHPjDAh1LCoHvmY/V/am+b622z/h+1Nzuz6Po9b/j9jE+jsxUOcyRh2kWt
PP6Hs/HI9HOiw74xZxZA8xOpxChfM0Hi5E+49GysO5vkZGKqDOsAXsqtJEPVQ6pcRyM1vWVI7ZQf
YnTiMJ7pVcilAfK7r1/euvWiSJL3xNz9/O26XiDd+ZkDccWzdZ1jDtdHeb8KR4r6snrn2KQdo0g0
ToXe1Hf90sF9Iiv4GkrZuS225R5Q2fxqlDoFxAGI3vIXbBOmCpC/KloNEBPzsB8BdcOWZm+JRCCr
W1wOnlprWnViuG+kjM1w8YVRoWNSLmwbodvv5RnMZNkk0G5wnRw9FGLnMCuYkRqGV+Px6qafp1z4
bVjcoVCd+RFvkX+RmVyVxqiSut/TaxSc81am9L5lypS5g65zGZW40TiRugwPwi6eu9nqN0vXx9uW
gDTME29ikjMvJPoQlueCei+7KADf16G/PRxCnYKNIHwKpetZSo9O0yflaE/X5cH6NlZrc9Vvf1rg
9bL+n8axVFaTmXeiYuc45aXbmHhqqhAzlxcbiNY6ATPeJfIEYIJNDxCCWWeCjXmhzRK8W2mKWSuF
yvhq/2aG4g+8XAB/U6VPLtazserAKBxVH6dEZbzmuEz/KHF5SZTkQ4nDw2sZbISliQG0j2rInuo1
N16COJIhx3WoUeY0RA2PI1RoIk0HGeVGrE+FGJ5mm3Cw5SE2BxlVJaHkELswQdYNRnzGgrqstfS+
1y9lfXoHBzzDh5EWsG+c9RYXzA58s0//R5/3BU19NU4shAACG/oOq4tT3hvj/hHJ6WseybID2jy8
/zthggc1KFN6vMwJZ3m/F9/QhdXy/V/mqgh6SeRL7RMbNm+BfTbz5JtKYvqDvW1xR6SgJEt3INHP
Z21x9QDXQLwZGiugAT0HrXRsh/5Wbr5uQkCpt2fCtwsnA9fLWIBc+ofkY2sqWySv8ZVU77ou5OE0
clwePcQ4FceJv21B5ri6LKqkHV4IgVKoW0j5klBcNUlRfiL+S9xWZd61031laxRwwyOoXViGENWw
5+SrY5RD3oQ8BcYk8AN9uIje+Tnd7xEG2YfS/cHEen+ICOs/rFBuedP/56wy0BCftccP4aIlg02N
V1x7xEKptK/HWlB1FmIhkSTFd6frvpGGOQiU6ksqRjuwyH8+V7oR/EoxLR9RG8GerjHjRndd9J6w
tuL7xGlHZqV7dWO1ljofTg1ZwkZ1YKBmaNQGOcwJU5NTKOyYUWuvPvDU6JrRnA0Lt1qKHzDDIEKS
g5vAStEWpWBRNSmnx3soNlgU1AKvxyWbpyEIwkdQ9J0saaf+7C6KUjayFe58mBE6gfma2IFjE2T0
QQLQsPcK4zOh6PV/8tZlYBr8DNMYD1G4EvkHyniI6z+zQ6O87SCJt53dCmJGicZBmaHxeh7AqZag
cWFwTOxvtdpHO4kk7qTGtanmMOas5OS+OKNbQ/D1f9wfMVMNPtBH+M3Ho4Gzdhaau8U8o1EkehlX
lwtcmejHUjY3fThbcwlkO2tmBR6+a1jU6yDZsiawfJhQkpmsbsC9J4LTlHUbropcu0ZBRT/9JA28
9IUUcDSq4LumS4N9D7hu7/s8Qe+7E8psXKU2oHg2HxHGV5rPDh9hKgpb6kPTFLNO3M2ELgCwzPxb
zSpULBm8gQwpIrJ5gbVeuIBsLYuBjtBViWpZ1jc/SCEUClGLrsKeC6UvQs9rlDcrhEYEqguPWnAd
0+u350sclART/RXXPjtI8+QQvMeH3EnFz/7Ok49K4Zy2SM8WUn3v5/1zPluZp3CaaSB91RxOfLhE
Qt9u5iYJiQeIzmu2qzU4jsB0IwbbIA8+qb65Vymu3UZONoiCKwjbODcUEcdt3Nad9qA5JX6KPJZO
GeKGR2QUjrZ9xKMZSOqh5j+rYA8j95hb9vYT/jxSkTYMaXkoSGW0HkU/miwRZF57sC+VSQ5jFFba
49/+es6RrzwKrVnWN0e03R4hI52j2oprjPJUuZpUYf8VNZyisj4bNlfZDnCqKzautRpAlXl+j8ki
/v8EU8zmS2otgTFhSfKjuLabur+AixdUhQwG4OBKRcGXh6MvAbAbiVJT+7bI4avQns0kQgVTM7D5
6DmJuHRgh1Trg8vjLQ/FdOIq8Hbb84hVipkhVg9fmrcmgyqOGzvMUWljyeSaDwyyuqCZAf+CsJHt
q5yLJtrmFNdJvqxYDaT9ur9FXWb1RfFivB57yqEsPdp2JPDPBsr3Pt2HEuKQwVH/9Q3RaWQ8ySDO
oF9e7EC+vSpOL9tM01RrFixudUS+gWoHbZslKZKChBRf5+ndAkQCi7IfwATve5y+G38rYrrzlmTi
MyEsmmbu3RJaiFdSLlsbFBUfv+ZLkzXUvjTXcss+gDr0c2YT2D3saVbf+qQdRTI3sKPZRFg+p2ig
XBadQYES0ZycdovCishGiBmqXqT0A2L5ln8sKe2VKH0mazWGUyMOiFB8WXevjNTkFBfBqze87iW4
tJBGP/B5t1wziRe8YhETmHzogjLv/2mixgzhTxx+m+rcZjelElkNCTy5MBBTwa1sS/uAt64pZVR5
nQ0B9ZYZTA2fuWXBxZ3cmw0u9vcGgRGXdbWrcct4L5aRCooZIQj+VuAGAG5ubAmtqVqkmkioeXle
xrL1G/zjDKYCbwKONciUmKx5iQFi6zXVcbpok/2Xw5lydb/KQTsbL785V8NrwTF+DYPNuH3UQnTK
qKJmDTBVDS9VeAjScGTTZqitcyIlQ1dJO7NWXaCB/ACOrnLQQtKxG7NHrAupHAlKKdacOQUd+nni
Q+qDUrX7bzGJmfDdLgeAGuIiUJn6ufdmZwvhogCuef9fg9jrsR/ZjZkMuU2HfGM02rHpT/NGekKY
/ls6yaofaJGu1B3IDVDWFI8opLiL+tVgfOXhcFCVX6LglCwp4mlytUw4MQpSakn0CTPe+2ogdNjx
BvdSG0SgTyc3OJ03lA9DwFYHAuhMSNPUTPoC6XC3kk8apC8td9asal2EaCEdL/9GSLw37uh1uTIx
5srPhfM5BuIxW4XV+wfMsaM/ENvn5BnrzjM+WmowpZ7/k8Pp7porX2jGCi3eo1ucSliKKy26mtbi
A+AuZeiC1fAF5oFMhkt8Iz/V1EgB/oS+ZDlEJWauOQfItilVgMgO7bEY1BvD16qAZlbxwG3BcVkB
BwVV8XzSKAE+B9xCSWBvkPWaDLkPfTtFSMfO4VJbZ8q+V0QljhiEF/+Z2YjVugSRI1dGmhOQcl00
6NonKX58uCJh16ERlJ1h+nDZUkDH51zxe7/IJBxkK7P+i2NVNKXUkUkqgi/wZ3HuQNjch8PfiPbY
CIxicUzexyvQ+4j3aO9JG98nwli7gKc4Hq4oJrCi6N43vwpsF9KYrtzrAlTIDoHQ2auSsGzjsXyq
AOOaijuDqO8+nkkknMLfHRiYGRhqrfmYBkzAlh621+UYd6ox+wl87qzOCErCV7PRGyV9k3amfQGs
Cop5LZ5+1npNAx5tlwrxXxNzWSBiDpaEGECKPKXDoC+IbNhpCko9qg+BHW8ZnVUtufdsHm/WNFYh
OwuSVtaLNiVvPNrNMuuliM6gk1insZMp7+lxUYnumQ8//PLByL88CuMOcNE5HCSwH9s2bW8vhGZT
D4RAwwDezvH9VXY6XtgMF2fGaQLlgeqrAelF3gFUXddUq7QZZC3AVm2YIEdDAoav7I4npMeexrGr
WApStuUovvAzVpnsH5QGWmaYRnKVSF9U1j3MPDleRxhc879Ezx43sV5q+U2BFybM4dhRNlEOsKa+
/IrJ1xc2oDx4ZPzFTjv7cE93LCvSUw0kexQ6nRwhCI6dcs0FvBDIdilt4QtpUTuU1cnqbNaSOGy/
ZgB+6LUICkHD5mQLMctQvV18NqAFa+UxiLoIfzmnvHjgqJqnVwNjZqifAFR4jNnq7tv9n1qi360r
Y0ou61tCU48xHbXt/r16ZXpZohLgYJLAaunoz1QMP92Q+qk9brwDVlcVhT4PzMQ8VcMyiB48izNX
FESc/obAseJdVD9ogC7vnjDU6N1bmF66D2CU4uu1qMA0xxpwCzUMtHU8kM0gc9+I16tZ2AjVyi8C
Ap1aKIVOa4GPNPHYQSc1AxseoeRklPmKxedoJYnL5KTtOX/Fpoq33QgUwgI5Zqym/2cP1tLOkBuK
qgvmIw1eeeKc+fVeeKpOQXjFS17yr7a/e+LVcgwliq+zyghepAlWkvb/5+wVxwLIkdFqePi6JRDn
t89qMDyxx1iGKwaQk16bglVMmPE89mRjSZ2uVrvprO2P4JA4ariTr+7jBQdld3aOVCaQI/YF91Qy
rTnbe49xuFS8KhNfUhekBoEeb3P8+8BpSif4HZu1sXHSteaHozHlnmOlOBsBWb7RAQE0QEuWnEU6
VDMsjSm0JZ7NNAaOVbyKOwFBMqk2I9tvr4pgQg84dRDBT9jj31DNPgb8aGAnePpw1O4Y3fCiYyOn
KGETPrIP+s8R9yGb/4NZkzBOlZ6fmdtBsZFlVN59gfxqCfnOOqqxmRa+ZRUXzbAKmBI9A+QWaKHP
uu8gar0J1sgrczdLlirZzxtUtzc5Ak2yPyR7gw+8uo7hOVgoJRxqC7ufzm3frgdZfTyuxlGzi5xA
nIZEXXjxlwlOFXvPKQeZT5OppEN5Isql12DjUCZHMXeXFiUFn95K5XtjjfWQowtHASW0mfFEEFI5
a4ABZhTVg+VEPPbRaxBihRcYrFjZ1aEOErrzy3lpqmsPzfioVT9H/g0vZT1SsqihRbKfjp9gMUs7
5EieEAVcapop+EiQipQXqJBrDo/uKnmWdF7QGhRYNch/J911qusCuUA23WxuDk9dR2yyaoFMI6Zn
/XsuWt6nbXvZ+bUGDhvbX/tiYyjwIJZH6aPbTpoKKVCET8iYjEX1BuI1bQkmT/v+oAZrQn0wJCLo
+mdStu7Hhs2dQtom7APtitRtzZ9f+oGzjqZZ33vzxlYRUkPujOcJVK6qN1n+LsK+KdgVJP0P7yss
/GXGuviloDr52Tko2S7aUQ1L1FSOsR6TBsJ4wPplpinBuL0+xUUqAAV6Ub8UBfo8Bo+0zqLosmhD
KGfaeEYkAyaI9tvPNrdimyHbFst/tjyNYpsnCU0xr/0R5nM/9F4lz+uiV77jaemM3WVO2AYVSW65
Vun8Crh36BW7XATxYd7gMImDm7VpsCillNfrpe+mD429t+VM/MDT5URlE6IiQ0M+lCfHNWL8xaM8
1iUhJOrx8Bx/QW9pjsx7/XkHlvoUiCiYpieX1mIGxAYxaqYEkDRhs7dZtHMw642yQw8toNsnzGBT
eOd2t3nmmIsAJhgGXYXnV9OTeG+c9Q6rRwPr5LOP/y8vLA2eDGT+sY/eHKTtb9dCX6xbL1O5Z9mE
OyeF6zdFCUjBU3p6FoD+Bv2v+6yCeCGq9tVqrzIgtR1WFY96eUIhDkG6hnvDTQDUbC1Ln7XK24IE
XYVblLJzt5L3uzevcJhnTkGhAFRP6SuXV9J8qEUE7awSw6Fzz/hIGX1ykFaIfRfs06pxjeyCLhb4
RZN7RamWs6wWPUKohd1/PQpbemw5eYJBVNS5TjD9324mHej2uDIA9yKMfIu7XbF0t/+HAhoYqIKI
OlKd8DWYuni5WX31OGNM8hMesXK0gGw8q/5blLmyqXogDqcuzi477csE/t7Z6OFmbTpdmLkvxFMQ
/qo8JUL6hgmkouVf4Y/0OwL+0kzID314MilRe5W0yumw7SRMePnMYu2Nkt7BZtnQYXzyQjUTuTRm
0mRrTPRpbbmF84HkshsyfMFdWMs0zBTZKSaD7lCCulltdrDW7Xr56aod+SwpQ6Wogge4o8c68qBV
x5RJOQzEwy9MTF2waZFYMOxWxzAVvJEbAYjm4da2bqx7+aXwKW++2S4rk9GYFdmnrAX3+Z/urPEC
jDVDXVFDh1loobtVU9r8wTvJ+0TArCJMQnK7AIJhVk1tQcgmEMU6M4NPzOxvCMnMjflCIHTO+CTb
s+Pf0UvzUpM2kp3VJUPjDvetCmqo44qfsSd2nkt17aRbrbetmKhTbn5P6ewtMzgTGo2+EB3NmFah
pjzv4VeuA1filhpeI527UbDRssrQt2LoZ7RSp6tZ/qw/26SZlbaPA+NwZ2g1EwAbLSMQWzpD1xBK
VyzneeA9j1VAC9Az8PCLBZenk4Q1U/ifuLgUHyzDX+OKstc7MPABAZeUydUvyvdEloaSay2PRQDo
2BWObPKFZknFRB73sSHNTcd66zjZL+8x4k4GIcZ4JVO7I+h6EmWL2AQ0Yw57rBz1u0kBYQgZQawB
gh0J3LT/H6WF+awtJ5x2pmJZFWJmaQEvy4bek535eXwQiZ2RxMFqE7lZ/ikBpoSe1MM6/EYmiNP4
Q8nKY1wC4yBX/+ZNkNTdIRkN5pSBfvo3KM9jlvwbwrsh3QKgXffHSpNC0TcHM2D/RgyPzVbANRSp
4N6ScaCgBPwdH0dgpgsf5zG1yzsn44bYIlShvgp77LyR0c1i+Lq4i4F7wMZhpAVxxWQQQaD9Tgm/
QZB1kyVXQ7aRjtlh0Fa5S7VnefhuCfoTS2HicgKtkIuwdsDiP4EDy/BNjnQqp7BBNA5nUhLZEYUA
lJQg8nIbY2rdxCfSipcNyCpOPdKzThREATAFPBS0iKd8lhVhEh3H+fXHWi9fN4uiTkEAZ+/Y3W1p
VhvoJCcLHkv8IEPYgVR4lLzap622WBcDTzUKdFiV3Gx8ZDLPlS956ldEabUphy+wLy5xY5lvg3hq
90bpoMjKc4TezAQBPww8LhbJkEPRqQFL/w9sD16RDvNowmvvMgIhfgC57iBp5iTlrgl/35d1SyeS
3IBkspP8n7JIrcMarUTd/8eHDyT6f+r5zaKNfJWZhNTwM8enTB60GAdccR9D7kCpgqadM7nWgjQr
eGSfkaI3JSdIDZpaZmUwWRhDmpxYiIb5lXqQz9t/TY0rYICLqxsNRZ5Ce6MNL5mibcnQJeBLs2dd
UFEM/kbJURfsj7oGGqdrRFDv1Ef0tapL4n0a4QxGi7b3tNUunQwhgu+b1sn1TaaNuW6aa6WEiQlG
3ep1/vkMwxYIDgGFFeEa84I8MCLHwntbRFCG1xItg8QKQa7UIDNPdCqM8vVawK//blh0MP5IzpFa
CsAQf2kxu2gQ8SeFzVoovWTIItcUV7NEae7KOmQ7AsSibqzgZ4VWoWSeS7rX3+x1/WVlzbhWqiNo
kiOTLXE/o88K5ZjAY7j36dPaPbTtOOwQdnPnDL0hICezt7dJ+sgBq0cxu8hvuzjiy+1o0T7O9NfM
i1BbrjIKb0FjwcEeNPtkrUG5NTaBWIdDlzbeRsAVb1kbjflvr9T+CAPfd1VPZLYs46bCsau1jcse
EBx/kfa5QXsib3eHB0yMOPWSXT5PmZRizOQPFTwM1U3rymjybdiswMzchSJjq8EIYrEk3kdcBRHa
WH7rksKMtVFIwpKzcVcInOymSduXheveN746W6f2LiT4BwVYsYqZ4HBm95hM9Rl2uS1oNhgg439P
r8LQer3sdItGcDPLMbyqCZLRUfvLuvdCxJxlUBDp+bTyzxSFqnKvWwcb0+OX6jVZi5IYRXgYa5p7
L199RSZSkj7uj9WEIGwSqOVKg+lFSaciaEWRNhnJvdf8D6e4LiMQz1dSSSlWf+4Bnz43p4T0odWs
nRMpUohv+fBwWNX6D67RDSobV2/RtPCGVF6KLOjcEd73nExRwEKVjEpxhvC/WxsipAudjEW7KLw5
ZVQOA3BvHIrXlxHpuDbWxn091xoFbAqJ5LfV93WeBahnktjE+Qeeb0j1hEpXQB92tcR5bqqqbzSt
lQgzLFpPKj50IwK13Z/IBE6LE3IFEZgUTpcv0xEJhmqQaZ/YPqhHTsvRtzJ3YIjXQn3cyeMEQcFI
hhWqWnaq66azvRG41nWD6dyMVzABRp7YA5rnBDsYxvpiSTx3LqMbmd6LNffdIfxXqETX6elRY9M9
7Ggd+0FCTZ/4e9iK8thnEVDOAbflD9dTRyQ8rerr4ppTiGTjQ/GmonhTSvehNwCzH2weIzdaPjcm
qKttqeFnsgU7gAyTB4PLP1eiq0GpOby2QIStV0bMskRGw1KU9Qwzb6KgIM9vq0eRbXqnS3OxBIuP
Ncs8h76eLXumyd0DUmV2FJYbIp7ij1UuJzAWijpkk7bzKGkHOOi2ypiKdHwSM/+X/H2r1aXAxbxz
dhcw7nqfewHvGAKNzyjVWmFDky8W9xYVDo3VTKclsy8lRtVTb3TBj1Pe/gnq+Tl/S1UM+1ybMX+U
VY+nFuTnUOg/z6DyQXDOKrV04xUXlq2JkUbhlt1+V8hgh337wEyz71Hcrl8wqq5Sl4MddYnYDscK
l7pryOtFetemZQXGYmUjy/5h6yDzwJdU2wxhgtq5Gf//GwHLywNJv1H1WlgM4BhtqzuQDNkspHW1
8gRa79RjB1o9VOEaI3Ci/lnwBWE4gw4H4J61EYO7le+lr+ULLIw2zo93joLtxpoVW5leIaYW4yul
085641YZDa73pFlfO5+WAaDZmimUeQJEi+PEEiSEvU+HxnvOIlZ5XdUypegnU9nYhj8qme9pt+Dy
xmyb2h0UqMPy7bklqDJgPuyLXt32JtBstY1DVqOMaFHOzfaDlLl+po2LB4oRoMTQsgkFwEO89UWL
bu1lq7kMkBXD8OL8kIMn+1XFoiM37Vp8roIS889Chtu/BEyLN2YZg5DSCXV1J/cUg4pLCt1qy94S
xR0KClKZpztCcfEQ3VCLJpCZe2/OtXV3cL/WRwMx6q1AVD5wyTWlthHArUcWCLGENxyIG9CSrVbl
Y2tyGM3gCZhzPNAjINLM+I2Rst+TwJ/23/xvumv/DyjTVTrRT/gZXM+eXP5FEHaFrDJi/2AjKFoo
+uU0lBpprC11Yfmtek8axHgiouvA1mz8qnw58D5QnPYMU7y+erdESHC+MniyjzTBdYaszTIWYhtD
cu4nmCwfcKJCiGTcGnG5p+sb+ckdmfNKrohDo0P9QFjqUAVVZtOBfKlswDmgyDplmKlYZJaSeJOU
n6QusjyGPsBERIc3fg0yatUCIpavnCwMgjts4B9z7czzTkGeiEdYbi9ajlsfCJ1VPGgOM+LK/y2p
mgeKMuVQQgxC/7p2SKdQv7uDL8D2RMH4LaySMrCIA4SJ84iYtn6hOTYX7dO0gkW4XFwr1kofELm2
wBedHPzuHtJobh7+vJ0exz4OZcXRqvgMgT/l+h56tg3YwA9qub6wa4IpPW8eLP4JGCPp0Lr/oMhn
UWcV71Fc8mNlqgh1yi2EaP6lxlEr548wDeafYvYcDd2DuonIj4LPaXRY5o631C0Tf5moZNxhO2AD
wODo7Nolk4ERzJXZWR77XhdWHRmsImnZsbxKW+7h5GUaZCHOHrYZ8WXvUqiGtsvrNcHoZoOOtrbL
Yy4NfR6awLEWJnl/wBH5gbHb5CqFPuHDCGGEuWM0Hlqr+5+FNhyckdSNa0MmWDIJ4j5QIJHScJYd
LfNzono5AgDV+aZiqf7o5c8WqRLdF3QgNmt56iHecD0j53mB8t9I+yM40IFF64vmx8tmOMt58seF
dKnyDRXrxROLz63Kyx/LOdnvgzbQCRZSC9n0KOvEkI88IAZP094Q6wh34opfH4WUsLE+ne0OHM2r
FT23AR+Fmd4B9edRtxTLX6jHSoHQyVIT6agGvPCZEY/5aCGGT52OI7iwB1WRNHqkVWK/httZ0V6z
mUuist7BdH0dDLXexwn2KXeNwDnaBefFSgV8ZlyN9FeOhRkKB5OUUOE7wPU7oHQYL4XrPDPzCXAJ
RkH0dncF7xmsxFE7cEZF92yd/h6vgNR6WDN0pNb4yjMP2V4B/F+40xubnxcJLnrcfzl35TyHTwcM
B4cDpe4VOyqkM5oQDXymOLZQSHkqS3oulklr9EiwNFMZlNUpb//EX+oLVXs+9+ET9IRGDQX7Vp/H
cOWKFkXlhtYeo7A7shBoQ2XFYHYT4eVuocCSwR9Ci9m0y1dHi2p6szuK1C0v8OPDSqfeU5JsMo7s
CtF9fcf2U9u6PQyy0IJB8LU3jJEKBNanX5CndxIzPYNPWhiPc2Bg1kd2VMd7lP3WqZfMNkYzC0m5
v4WXH3OKPON0A22/a6uozsBgGG01Yc6qFEp8fyuQIDA0Fb22tg4AZHvFIq8AFGNPNKN9145nqAL/
snKhP1UMCmjDvNk2yGg4Q0WBf17ccIsYucpFZ106/I2NGnar00C1THJMw8EdZspJVpcE/kKf5wM4
yZ/mtt3d0st8pt2S8OV5uqEx0FB3B5cZ9rRzcZt4MsSUlmiKGGk1jRziTcoGlbUIixARuofKGUra
4VKiIXpQdSZqcvOuVr+TMdyPCFB6NAb7GZaYcMJMvbMS83+OwqiSNFg9dBnmOtoc1k+6wV6K7wPT
tbHkQewCOrUwJueAEndj/aaO1D8CkKQ/nK08voX2yzvC6pOiut8obkLfqoEuUVVqWyuBmgYfkdu/
QZdC3+qmBMXo5VisbaMDxY27DR62x98IaaG2gKDOHPH+mm2IGLwtvxAQafY13RS9KPh0WEhuLzSi
pPo5+lhM0YBfFtFqmkFrSKOjSlKFNVHnqnmeiWHu2/73K4h1IMPtnuDpPBxFB9o99e3G4cxPl8r0
8PXcwpiK38OQqxk8FL0OlL4IJxUyWcBYCxFvlW1HANP7KdyneMul0+OFj0mc4b4za1Zd6EPdJoQW
HEwxBAkR3Pm+wFRpAWAzwjHaf7xLbXB1lJM0jomMn/ZHzSyGH5Wx+WNE0Fog10S3o79EumNQrf6s
Ao66fLqY4jj3pPcGwLYuoWdvVCIiwLx7t6wGnQfe8ID8bGw9feChGVYTDysK5RlfgsYSw7UPSHl8
Wffc6NtAt/c5okwx1mF5mCgpHg14MIPM1uAO+aeEEj7eFAWqiXeDkuYSh8dgL0I11ewIAXfhG4OK
zM0XqmCV3+Gjh9v+A1b5sN3EQegapSsV/hJLGitBtQLUGk6ccBR8qYFzIsl3y40OrGnrSgSE0zMw
fM+oYxalDH7CAH2v8o6fuusOKlJb0SLRwcYkPHidyNa+4PWM2vmBlYZbMIj+rh8gAzwGyBkfSrlr
pAfdJdKCIt0g0UL9pLk4PBVzOOTbtWh2v249DDwN1uO+7lCPhcVf+6dxdXpuVW6PvjLl5vuRaLKM
3YHyqggxuwl4p475kYXcLZTa6YWC4ORCFa9cE65sdk9xtR+pWOLtagoVTCXxNP8ugZWj5CyHu11l
OwoDMtc91NSNDAhtnAvl1Yc2+T8BMjHBP/+OFcSVO4CCh2XcfeIg+D5IJb3JTcucrXKubOjQUpB/
99jjue/DgCcufCm4izbPC4Kue4q3uYAHMABX+SKhshaj6W+IeOahQWo1IGAx44UIByzynSFaAc8D
tP+6mPUdRPbKRABfrPKtZKDv2B5y5vUSiaCp0+Zi0CiiwkLqlJINYu6Vtv+DbFT2wrs2smGIVY6w
3zY3h2jIox1FWpgL7I0YaUfVxoCmPWJB22siRxKPDbdpztskG2toY9hTnPhXiiiQn3RLTVmoq7I+
WMrNpv+HQReP3xKBRWAqrQ6/n8yT7hvQW1esnC0wfGUvzH9FnyZsfgGJLXg6zF8VneSBS3zOv7re
d5h5k9xj2o4brI/YkPrdkeAHvKZXhLu1eWLIVKFxvtWbwRnRSuvWZoxD8nMgP2xPJsucrpG2/fHQ
IQIVGg4PwLEbxePLF02My4+itWiq0t9X64hDYIUeu8iMPxZmvfoVaVQZeQgLnzm97C4hYKg1/vru
uGd7lotn/O87oCjcFUCvCZY31Oog81F/A+sm2tKdFWD52KOyhEWg02gDwfnjCoxfcRHU2znpLq5T
mc/kOCpW+bJxoadRXNGwRPfNaGsvTkSkJnoiu8CektL2QhZ1lv1DwTKHmtq7GhiLZHQ6tUJNx/Cs
TfuNiSF8/5215qsM21OtDXAREKGloC8RmkTfSqrkzaD8t4q5TphIAZ8C5GcP7dkRg/xxHyhTicIB
ZBaVO8tIv9m7X8gbnkaaXfYxu13UIXJtk9/1JJaAFIJmAZsHa9nqaGnizP3bHIsSWv4F+7Sr4eNW
VIVxwac3YRa2E2/AqauwxBjLS25Kq2UhmV/L9K9GkmOjNgr0sm4oWc2cZlu3oOvpvyspckN3iktH
LE8Vf/P/YuGvQ3W9HqWSRc4QTwuX6b/JCrMgg5v8cB858iIvQciFyuDV8hoOYx1nhs/QR1A+Gb9A
tOSsPOegcG5PRD8z6BLtD82L8/1L5DJaPbcCov6NqLXSu34Cg/UnA0qx5zePTb/L6chWIV2kBr+4
AyNsWeaPDwhBa8Ri47V6LfojMrmExal4a7Sa4m+dZIu/pRCCV1gqDoVFcKOQ7K95mfQLWqiT+6Fj
tm6vxhI28ehet1qUHE501oI5xUY/ucI3Bl6Z8FyTqjtaARkjvaNrHvy0G2gtDLO0hbse3b9uYVjZ
SlnlM5gD6YPXZ6+1rMG53xjvtG4vsHL75yNYwcNqo/8UxwfHXccgfxdJrycXFBA8Bof8cOSMs3Rq
Anux1lhWGuO83T3dfbp5hehXOOc9TMjohxIgWPgzHb3w7t2ww4DVXfEh8myTLrQ+Q+pdTRdCvWe7
VQrdoldrsYvZEWpKqBJlGq3BMXdo5sNZQgndAPViPWPzkC2XrO/S2r+pkrnl3yFwDySrJEb/cHrQ
cXspnRGKuqqOdQKhXUKyhzaI2Jo4Zwe2yfpCQ8tkbifmnhIwoNKK5nAUM5Tlkx6P8yxd284Z/MMC
7oGv/GrUdQ9OkwJAfMZxzTCe6g0VSt18BL41iGTpBPUP7/+jDMJGPu0MClIWh8SPZWIZWO3SU7Qb
3/OATnNvvlet86U0NxfI4JwPei+UdgiM8ALrtoy91p8hQMpQTQesbBZhMnv+6r5bHpJsg6lekCW+
B7JDNKqoqfSUZe1Dq6Rf5e8KRkM9RxMrAS/qKvZK/TABEEYQRD7rzjotFPPtH/KUD8p82k7V2lc2
sDY+D5rVjoLxRaIpnN0nMytX3pAHbarR/1yxFVaAjvN7SAXGh/2rgCdXZJRXmy66TIrpDLMoV/DW
PHzVtpcK81qzCwgkvnhvXSsNhdTYMIkW53JyzJG20iCiu68joSm5vYQAWbF8XugHAbggp3jf4/Wb
nVX1W3hfGZ/7lyjBD3N80T79ACzKLUjW6pfBHYRuv2pRbOh5tssi7x0sg32jS4167KW8MDG5uZPt
zZbpC2Oa3ZsAdHqH/DNZLBtlARxarbs8iHUKtSSQxsfZhYK0Z9tVp2Q7k9Hr6XmO2YTNtTtGil8w
PPVoh94c1itXUyni46L68JIR+OsapSL/GFQnplxrXVl+jtDmmc2RsLZVnsmNaAWrfOa2Kp4ri3tI
AmlLRaMMz8r52dTynmudLkn1vIyw2sXsihCxFhss/L/tgDanWbrS6UXoln3Y8nes9flX7oW91x2A
2Eq81k7/nDQxc/cSv2I83tE50kyGGCVuI5v3vzdl6YAmLtCFIILXr5ZO0LGt17PFrRv0SQMiNSC9
v2BSQ5UZ5rAisZBnmw+rSirFDhkNOlN+KnoPd/i0+gru7t0IH99as8/kSvwRi6QlSI1ZCW24hboJ
EKyGLuaEfyizjxOQWYC1RV4aSRQQW1e3kBjHptG7RCcpfv0LTBR5d4rND0oiDXi+LsVzHag3fg1X
tjHj+d9HdDYt/M5uyvJscQXTCtxZUlAONeJwpa/Ah6UU49hZ5l/TYBw7MOatJgjAk/bMyol5ya43
lUoVtqQAGWTFkC+onS0GnI9uUxS8C0imilgVyH+nRTX25MrP4LHjkV5bknD84ABjaG+tKu0GE32f
AQAqiJCD1MvsRuOUVqJjVSjwjY+V2YwSvkTyFXKj5NxEzUNQmbZ4xNL6ozZqlO1aA6dRcDT8WCu5
MWGQofcGUqz3SWJ0psYU2N8IqzLP1Oa6cc4qf/27rumf1Wc8qJ3b94Cg9lwRLiBdVZ9G3m7vpAGp
f5lCNHV0EFy02jH92JgSWuqt0Aicds/YpgCypivVa0SGOqx8C0a7ZDb0eogFvfAUQFkeyRPVZtBy
TXXr3WnMA4kNontDG39ObKD9SFhNTqv8agIYvavYbeFLEujMgMKYwfvmOQVmapru1hCVthpsfIea
zKr7KPJwRXM2mUD0y9NzsYQXv+ZxjhEGmNQrjlAJ5d9pZouhr+VqExqg7LO89xNtXcpAqf2U3aRO
SomHQPZG/6PjiS8z2EGjeHVcKIcBlsBJwbRiKD0p4Cio9vVFXoP8HbY+dc1rLE2qbXr2R4nK+K1K
C9fkMPJNxKzsYUQy66cPHjmOpYk6HRjXEmfFm+8geBfWTvNmiuSSU6Dx0BrQyxHwNvFJM4HwBQhS
AA1k0R+A/WaaZ2dwaV571Ls2e7h6LlGrMDsKCBo7+1EdmTQ7UMmOvAkZd7FW2CXW2yUTaWLBhgck
kdC1OPAbe7dIib9SOTorPyWxbCYFcV14jChemoffuI9vM4EZ61NLs20lFSsOZRq13IqseIKvHmeL
qGPi6iCPY9eR8rayUV2wRjY7lcPkAuRymGy5tszbDcnalXwNzWtGVJhMW+6LHLdfZceEe0kNeHoy
IULFAoUA4WVVoU+DeacrkQlcK7VfVye0nqKSWyzs/kEzjKjsL3QjtF2RXdRKOlPfz2S+Jqf7xzZt
pGXTDXoLS2lLIgbKWLYjOUnJDJIr/XYxfk5pW5dRK95w/STBMUml+0gMKivA1PQXXUGHW+KyZIpw
u1fsyc3zCeIVVPsc5ub5p5U7aAII8HKAnJFX/vITT91VXbbZdYauvCxb5stjYYgWgTTZjdrn2ZnK
znRFun7qtru9V5RXXa+OmiUNEcqGuyYMk+2ptd3tyTh+V8CUnfIQc/SpoNC8mDUf+367NdBjy7GV
qwGAqJBYzqOp/QN5DF+gShERv9vP5Ocq/GcouLRf3215yDXp0/bR1/VxmTMOYcQ/3PueWPj/s4Y5
nfVQ2/L29RT5EAqt743E9ZgcvVlPXv3vaW26v9+9BLpdu9USdPB85PlSODJKhoks9l21CkBXyfKu
hpI2i86evnTAeblxPTpGryh5LttGtT3IRzGFRHSFdjiR1xn5Gd91DCUcvzOZrDiy5ytqMqOq0t0N
/REVTSfsRybI7tPTGKLxILErqeHq66Dgru6t0ZVSSxgPNQgKUq1yrVuIJzVej9ziSb0YUn2CRuPI
pJow5bjD+S6LcP8BiCp11gF0i5+rC+G7nblNG1+LXuiKs8nEKvg8/H9Mp1uKDlzEQEQ3oNInRcCY
Bo4O1/9iodCLWWjYMQmPrV9ub8yA4ehA7V6ntSbIJEPQBNbzixxyIiUBKraaCZCm3kOjvpBsU6kE
14HHiOrTT62gWRHn7BnNcuh0OaddRxJ5I2fK57w3D/r9mhjONDZR91Vgpu/+uK2RXwijNNNOSlMf
6qLmgRrjQmC/KrFo846M9+uxIWvx0HAqTCJiVaFLl1f4JjsD7SFJyy4zoGXGutddZfXwcqpWx2qQ
cAOMO0q0nEjsmRHlx2wmHex9H6b4FuRO7IT8cVWEzm8fmjQsrR/SFSWo6EKf1wiAZg0tRA25un46
FSAQqFJH4Hj5elt0+0PpuTWPfFQoqsLYHopUakHefgOOns72smsCk27TkGDyHOW0p3AN8RefX7Qh
neLJknhrMym2W48I48+/1fcyL5D2oUS8f+jnhugqfC+Jdb8fwLz8YVAwZb6iARJb8T+83pimQvMo
VWsAeAIFQSNHdzGTWoqSyfZuGbSTDw8GlpIgMSIkupqijeOJI71y+j0Oc3Tq1D1WYq5PMNjcPOxS
0FjPOXI+EmfNGWVoqLR/oD0+PxUe5nr2CKCA9CQs/mvjDWYHcdMyrj3gWe/m/mBYn2142P0X6qx0
bpUPvkhSKyeQ4C2TDVKEUJ2fU7bzN3u5zRD5ws4bGkX83zBtQl6TTfQCoH7OFMAFn1Sl4uI23uy8
ZBU0FwbKLcVKjYlGNdQffhiIy86qY4An8yzqb2lfG3naP6xjT6Yn5RwWodtdAp5J7Tzc7pqP2APO
uteN/sypQxJrbZYI+ZbfEupyIx7emXexnhxIx0UCmNv43r36M1ErVvQVGUxynm21WHPL/R38rcyD
2g+rmgtbloHXdLcVkZwTp7eEaXmgNPFHLXwoGJYaN7Lb37RQIHAbs6ZrqE/w1T3YtCvKsFH5tvx0
xHnfa1KOh9cRCq3klaMOQMkAen5bZloI8sfHI933aghvCD3S1qGi5ZQYMrArX2f4CtojtyuL2eQf
4Rwc0PGs8v68hv2OfbEMv60gaQMPoGH66LoIJIR+iJyMHedvz/HaZD8XJW7f621pWE0Co0QEhALU
5E9Ws62ZcoVPt6E4VV4LSIhsXbcp06uf2bzAgnFWkaN+UGx0mtoYX6Oh+ITDJVumF6mH9F4SSwe4
Dl53AdEujmZl1UimwFMAVIeC+dUQGkUXHk+ARyxYGa1IqB3thjiJyo1l2nKkRTXHiHbSAYMyvIxj
RLYiCp/QvTwC1xGbO/OxDM0Lrc9FcGzhePR++T34M90n11miEMiFV2kY3t4c1MgtNWFMFhOP5M09
oxKUo7fZ71HG8nVneJL05Zw3znObOTJphxO1dITLy8+e03Y3qT0ypAcLisGi0puqeWX/Y683ew5F
5qruUbdanJZZo1fhSgXXfucXA5RMHx4O47gZtXASifWRr/5YFkB6UwG7vTxUhIoMwtew8L+8Ges2
SpN7Zj+jOTP+mmaHpk47I1K/akGab15wS4eK2Vk6zewlBlLTm+MHVEVREmvkjSY3KyZ8ZoIsneTI
UUPxcW9OGDJOygHYW3Bfx1+aks/ONaUKmQRsSonUrMUapdUGkjqTYGIE11dUbGfqtrITlZgPrPBC
vZ/pCNSuGasK07xPkKBw7jbOWk3qXWCFTJrU3WETkVpdHdJ+uP9vvrtxRlwUmuRM1tLK2Bz9YzQN
nkhrF4d4D4scdELcYVTs4Y1pO4Zs/XaeTz1yrPKP9RCEALTJ4xMfgsCCdmAJtiLc4/1dqiKHCLcg
ikdQSviXNnaJZiBHR5KYI02m+UFgra8MNlcHRTnaiOTwrZkblrWHZ0bH1B/3pTv9MRVuMAVjZb2V
0RU5H2X9ddX7aEzesF3KZ08N6h8inlzHg7IiHszC5qMM6sGGgJeZFyqj5HFa9LzPJYfWaPBKIp54
u8Ljk4l5FBs+RoF4azQLc9S3RcqMI8v/pxlvl5Sd+qEedJVT5KJoh8imsrSMdMrW5W0Frc1oc7TK
1DuWmQyK9K0Hk9JnEnmgYqfdvMt/DIjUw4x4SoVcpawNA4w4pVxRSr250xSbnHeMv6vFJSaBChY6
iVzCbquH+0UreUucFfOYeThcsyrOADM+e2d9T0IzHcF1PY2CQfrzSYtlhGpa5nccHK0cs52s5y21
H/M4hk8XAWJ9Jtap2c+kjw7mmrdys9kVJokNZHrivHgMcEgB//M3SDVHe6bVC8FioIGtg4jKqGZT
+dsdYvLopA6ZXwutatmrBMRHAeRYHr5PrT2cmeNULGzCaKIezDGQfY+k8mlh4aYcYhf7x14Wfpvq
YAYsXTENqPhqjQBNmDu9vQ8oqAw7EBBz0YE9+OgNR09Kwa6HXq3PH7BkBf/5+yeuzfsv++RMhXep
c9tbqNqbToyUbfKD446q9cCLTddOvWeZ79lLXp4jk36aLh5FJBQksWVZY+cAd8gVUyT7T8tL8LTm
tH8DnKzcyQ+DA2fIe8XcWCmPgl/UDxxmr9B+0JyBZWbI+ZQCUBrepj1Mk9BJt1MBkA2QieOjDNZG
UYBSExAj7iM+yCDLYazJSr4vawM2aZKqL10umaEMMNcoD0TdX8fRlvmbxjGEC9BhNw9vyv3GFMfz
RKiV2rbWQTV95Q43F3mZUg1rPh8qvtgkj8mQg6DjkZfg6fjCPvYjHB5BsVfdcmB9nBOTtpgHEyt7
WVVHWKMwnCQJWkw3W2tQVgFswWfh3MrZJkkMrWpUnA375DcM+hNjxlEnIgn2vhM6AxB2IczsHkTe
5y2PqzQmxywNwPuATNqSw8HWqAUr7K7SI7VWogawAuL4puBM8O5CDF9KpyVz2DeSRN1ZVbnJGD2z
OzgH9A3KwZf/XsU9tnUmOi4Capzw1byZH0YP2FVIgbLeA9tog4R11nJQmprbic6ZwdE2NnLW3SjJ
fgqxanmzGH0eC9k8IEDnZP49qaQ+5TjkkOHKAJLj+TaDiNSEDGshqI1sYDCoR5YtIndIs0YKJ2DY
Wnyzh8SaptuQ5kTBIev/zmG/SVg9Q1INZ9mBrbo7ovtbp3z2lx+aIk3QPNWS3tYstBUQrjXfpxVO
2OXWkjrCNCYqOFXpyX9J0vHbZa4FdbpzESdaN/Cg5aWtsiK+sZH6ibveW1agjooYdnOm6+R0v569
8HIxKXdFIueBafV+jGf8s0NnsLI0rCpIGIAHi5ZGwMpK5bLAVW2iQuZYfWwUKyjNDiOVzpTGXXZm
x/ygQjDBXscXeo60fH+bahZW1xuJDXPjdx/VhLc9tJ4Wl4bjg38cYXKFhCNkgVGWjab1P+qZjklb
LZh4Kpca8M9vZ1CgcTkfypQYq5KkCO9gZN8eM311Kab1Xmk3+fzUUjfUwfDNjNhyBWo0etgLpKvU
PjsmNRgMc5PW0hDN5T8UeHlCMuMe9f4GOEI3swk9/M4POypGvRS5HxuPj3qnsp9wJeUzLZJVLiOo
Ce8rrIpzL9bNNexU21+jDRwT0fUfzbVNkY2hKUjt7KPOkKh8OuOK/VdvMAOYPrHYnfT3hsM+7lcJ
P7XXiRGy/WYiA1Sp1vztfo8oqWPmnxm4dA3LkXlvQI3KPOo3c3kBTE1nfDF2rgRIYr7BF0gQTau/
/xIX8/3hQZWkoAX07J9WmsDkjqxZQFefK5Qxqw9i+dsV6mq5Cm/4gpd2ZJJYzK3QpRZM6ccd2gGU
7XLb7JT5rsOtftcu0Tr3e8TC1U5isREHnzyWWJf2K01RRnrroYs/0bwcEyJaAl2YBhWIljn+EV0T
s/77dool5uJBEDZyGyXG2pNNUKmRH1EBae00UEmuhQdJNJyfMVXt4HLFg024rWdzNHKMcT4bUFmh
PRZjPhQ23UzilAS6zg58rb1PXPzWlmXpPgI93IKNPIi1Ag0H2CbYMHtgWL3NC/q48eHyrqoACIFN
4SqXK22uHVFCMxDIeEdM8P9qwnBegGpC3H8vogsvs3xou0Uv+JozJy+uw4IzD6FFuzKqazdlOQ3/
w7xiLp3JaR5YVgar9X4joVN2l+QNP0l45Fl19m7nolSua0Z//Egj/fGmG6xD3cL4fSAmHPe99oOJ
7/FU/UbSHsZykd7AtwX+RfPLufGAOToodDYl/SReZ8CE1ceAl1XEuVwPMXdKfxbJZYqgvQIB/8VF
gbwFjeJ3W4Oyu7FFDUeDM75CqAyEnFKZjSwbwz7hjGM0XAE6BtQp2uEyPXzX3QniWf61SxLJ4jn6
xQx7hsZaD2JmgilXeJLfnVBG1U/A8qkkJqit7tOhPUU9xPWDB4aA8O+HvzaOeV8nXmcd5WaeHaZQ
/nnjdQtR38etb7k344DPWxdUj7+SVJqOM+zebk69bZ8IEqERbIYSI5q3uTfyCakNFTA/C+SNx6Ox
ebAgAzEVT5YlEO1449BeaFGmzda5Wc8o/EGzGy4gYPjp/gHb1UQrrl/UdR1QE41yuKxhAqRDiHW/
1zMnLZFurjRaDhFPNlWDwFJfYIhAOOa/cIL1rh4t9jDcSbEFcfqav2ktpg98QZId80XSePIMAZkG
9kf+dSaGXOxKLtdE6PIw7CiumL+HJ+0+7lFfoTonirBUH+HY4J8Gul9ADCQDhMflTm8hJcjRpjjN
1WhLJL5aKADvr7cPoJKZncGHrXRQxm1+5Hpoiy2trDqv9+Q9X+xL4re3dVtIp+CJpjUG8kjklukG
8bcPhxU2FjLeKeUtuO59sJCmBZOAxOt4FtbCdAmL3gBMXHKxzcLreUTavrSLYLqpGARy9mkjuEJs
qECw9A4Td9LUdOQwvsHvEKd/uEwydC71KSOGmr9Uhuh+AQA8ktbV0uWnvJtKcst8p90qoO/ii+Cm
iRrenM+LX1l9PozCD1d04BSQmTwwNt/+3P+4m/oQrXa7Yk9e4Rm5g/Bf1gTKHlE8j8OgcsiMrNPU
0FHjblgX+noBLp2BEJGzv73qT4Y04Fe4Zm5bOu/UmF/JPusiMXLfpU96N8wKNJrAv4w4qYv2q9rq
NrNpDZDP+bvYgoK7Ib+teA9lTYVCAz5GJgSu8VazecKDtRWf2VpoJsp9976vTxI5fGygiV1+pvWT
aChD+4m/803ZlXf6uRBDG9zbYyag87ocBF1j175lheVgvz+RLGW5XkkzipaCkKN334/pqSp2IOMr
1gfSezrhAMDGYNbqSx0yqZxRz5Kz1516KgjEPVxR7mnm2AR15ByDk2/jh6d0MFxjEFBpPa3lhSlo
enaIf5OXRASPdlNadNRZ+jjFhV/6aIp47fUmB+jF35SIoVeTeicRnSPzBRYYe5zvssiRdAolOLPb
pgraLl/zGEsRm4XnLDO4GcpWFVHcxmYuoJZvcnR6AJx6Arms5RWIBXnuH3/MzZobqE5kN7T5gAmn
7Aj8l0N+p1Jj3DIQFgON6QqNhwE/cl0cqooiWlVytmNmiNogaVHbJDF+WJlVlfytycdNp0+jk0Xn
5lBShATaMQBwb8ZqkloZzALCsZ+2qZi632bXLqDOs5Hh3XLQ2GTJk04nnoO47kvAYkDvyfYL4rXA
XZAz7lY4jnRRQADiKXZxgnoyy3icP/e+JPVUV6CD+7fsucr2avFnGhEUSvFk7+tqoXjeEU+8U196
FtyYEFDPdt/aOxGqW6lzUuCAek+XbXdf6Ra2y96znOvKHMksCflqEhn5m3VRW8v3+8ffe/VL+DpO
NVUTOSnX8CXks/C/e/WaOlrkbIJ1fW890tXF5MoEmCVTxFKbgtaso/EFzducW9q3jLc3Rbr/V5MO
OdEuAAlvbxtEcpCWM5XR6KG1QWGHUbtAl8fpQeB4VvpD+G319hKHme5Y+h2AbgJxgbXL++7+2AVv
hjkViTjtqT2oxseFSMqZLADF+WNx3+FEky+PmCNxxoflbCDqBWibJRbLyiz421l487WhNM6hz1xk
078x6At5TyAAm+wIFyEkIj9zwvN3zuUlt4fYFcw0rR9Du70yvXrduHQvCVd5X8gjbUwAUHbVDXPL
iJ9SwWyE0te6OlhimYqW13TLQ/I/4YaRLyUF8+15qESbOEt0hrtXRL/lTWBXiSWffyGsdAqN4rXG
KnnuAqVBt0stQQEDr5LeS63VZceH7PMI6heGDtk1Qo450gRMD5GQnpcpvkl8c3vE0aWlT8gAREAP
4EFFuuBncjv6p8o6N0yKavJhPfoAe0Qrnjmx/34po26DhD7Qfnsk2h7dyfasRBsT9WjoL/+uUnUE
Wu0+wIb3OCz6ECsTh85vv1G3nmVk7/CVTslsFkV11/dUAA/CQkexwITHPLBhqcm38fnXClLdQYgN
W4R37bYyIjIkdjvF3QtQB2Xji8H6bem7YIMWgu8y2ypRCYrfHYHFrqsunPQgd0wn/zn2OvlvP5A1
P+z+UApHcbjJkfjd7D60whO9NFauvcenyBoZ3nZu7tbpKEBTpIqGQx3BS9aPFcdKx1c3gCsSLYvw
C015mR0JTozRHy6Om8O6jvZvfeyhWjepyGDExlqX54+yW98apaxEpVKsOGBZy+J0DOkc+9Kv5h9f
3JVNFFZGamDh0umlPE2m+qIMPIB70aKcDQPn+O6+/sKuP7z7CAsd2bjPXAJSTv+qiJBuIx2d6hBL
g/gy5w1nKDj6O/gwyG2lt3BHXdpBmPqGKCNkaBA55diuHuQAR9vPi0gKY3sj72vfQpm4lv/5SNn/
11Z/qdO0K1zh3MfiWfkiP+v+sX4tROO0Dp4YOBVvQmgOGeI7BgvhYrVfis7aohuhqptKUJUEdncG
GYo8r261yRvjbtYomy+oCNbqcpZsoLQTn4KkgU5GLhasZpQXT0ftrkPlqM2DvVBk7UQKxkHzzDsr
18JNkhV9Eb4z1TRiLE3K0OLozYufm2bSGHQbLU6C0QxZBI9yoqUVowgiTAH88SaMUborm8xDuaXj
YV2JujV4EK1h7Clo5E4E3vvpmHaom2lcejPiqZFEeOZi1xayVSXEu7SA1p/bNCCTdv07/YvcidCB
0XqeLkfdYVpjGLzqYU2BxVPujzexlFLhF0UM27ZtCbKWVT4YHE5irr5Im7jUmOEKGb/iBfviBGzv
3Mf3Xcgxvc+Uq9izaE4V87hCz6hmohtrVyfswoiwJJFw/1h2Ul6L6p7LQ1EC/wghnZbadzCGWDLs
WkHQfmRfjfKGB58jo7p9IKkseQlf+G6cxUG2gdszMez+tZwp4JF9TQxbluAnhQ42hFjn/5Is7HYB
XAgyPt57j4RLAnXQJsfb5DXm/oJ6QhoQQ1TqLvlGUIDgpbUouX1h9EgGNnWRhSd3pIw+1h+MAc4F
tZ6796bmF87STj7e+sklRyeZLjwVlJjQlQDczBzbZIZ7Sx1GLIQE5jRRcGn3DCct9t0uNgQq366T
KuEXMHl6RtQvwCgbftUE246WCMHlWGGHglm63Z8j0mHJZ3OJelTqemG0ns7yQ4ccQ7Nd1zfOzRuY
6D3kRrIpCs1ourB/TvQB1PtzOF8apKrZxvmesxcMHmo7VhNZFRo0JfzptmzJKg+Rcr8JWbjYfZC3
M0nBv274KzudUcSzGDcQVW37wmHdkbsQ7ODvCQkU6Yotqe5/pM/I0vczF/sqpXX+wipJl3tpA/ys
ovF+BAgTNeYmGmMxxfNhnApfkM0YWoyA/nkwpC8pLjJwKUmAZu42454nFuU7Z8ghdl8P5/x6HmPA
XBU4fj627fHW9zzf1qinNA2CF9O/nj3HYZlCMnaQi9a6yIpZzdrYL4MI6pstcRqw85fjKW2+59r/
kzNX3JO28SrkFnj1jq9fCzxrOe4/XwEYBIY1+KVbEbOAD+ymBYDFwgNImCaY72DEZP7SaGo9GCwW
npSM1T87+/b3SiyEGcS5V/0O6CfK/7qoiX8TForWGW1ISC66InddE71Udz6rPsU6RJ4GYHgp5hYd
/kc1HDfVc1hJUNfPPAZp4I9cX0x/hxcBDHfGhbG0/+S8gOaFJef66HAxvbCUQExOFo4aYELc7ncS
UDy+MMpVMOPtjSgqxxkKgRNP575Oa3T/w33kX8Xjlmdal/L03VY3TfV9J5lSdmsJMRRFYfaTbpVS
2BMkogxzQVqnS5JUemmCE8l0yz1OT/horuqvSpJTYrcdo7M0NCzBVUre77ZKKnHlRHiOZ3f41G6q
663hIXrKzB7KA+pYhvMEpToN0e2VNLm+e6fPOfFnNhJvyFRglXCgY0YuWFxlSaGI5v7qKGPZu5kC
vvItT29WkRd3dDnLYt96l13nUoRS7GYMdRSP13y8biDo+GbNhaaNEzyOLGjdOfyLjAL0yzzgXi2+
s96gyMxyQiXi1hCMf2v5FHgvAf0bGt1T5ZatbiJAgpwXS2avOQZ0Emmg7GF/J4vMi4OLU7CyTWdA
CsWn871UNrT8v/FhfDWJHnmCgJvmXkOcTUy9qDstxJJb+K77+jORVnuS1sU3zbkPGRyI4LMCIek3
KjVV8ZP6b+JTTfMLHcaTXG5bTMhJ+yapYvZ7YDKpMOFb6GfbGTDCkqyi2lKWJmrxawkJVS2Uqxg1
ByfP/l8ZPWzKM4nvQ6BhhYgv5K1EcXZuayROQuoDR4NedtdHXz4tLXeso0KSKjNYc4wZpsKzx7YU
QqJD8HvBCLjEswHCbdG2CTwfJHHxFkr7zfrNOKG0r1i/Vetong3VAjWobUpAVuyLCv09IQlPcvRH
dVkTLpSaKCl5mPblA6B9EqFMxVPMI8AziqDZo4kTXsfVKw2G5HPvSeM+yWBLMjE8mZPsXC+ZXjm8
V2HjwYZlm587YMv+QSg1lCj/bIpv9/hhLCP8ghxqJDnJsrV+xJ2q73kZAZQid3Tx/5/QoemvKTvN
bW3PT6RJyQrAjuwkC4kzp5Lwh7nF4M+so6cld2ASj3It2khlagLeagjSf3NpJ+YqeVvbi09Pm8Os
oHPvIVLsDqKmbZqD2v45bAQPVqp4GtAy0gLq2TxeQAxFy6aUSEkKTlGT0PROopIoRuIStusWPBuT
uyoqpdEzCgcj1rCjjgiJowGnMlZO8AU5ShHRPASQdNKHXKKZfTjYQi0huHCFTRocDSBC1zrf4ymo
7n3aBWOGGGlBpkqxTx+7hlXzwblLCM1hE0Eyc72fSkvAxGouzUmdOSSBXNImOc3iSWBQz8r3fZNy
wPvcG3pgnQ88o5sDw9EJcd884jPXIZODmIT0v0Vq0OE+HfPJI+AOlOCfGK6Vk40jtvLhZ8AhdGjb
YNQcorbYqjgN4dfDQDLPtvsF7TvvnSGz3I9jRP+NU3CpUYoiS5x76Mr4h7ck6VOfSBFs22RUO86V
wpFVwIiYhnCw1RSNLIGreawXmo1eOLDvSMcmmAsk7AGkP1X11BK0NW5xQR5IpfJ5HDfhG9z8gzgT
iHTFwJyOWI7fUUykZnWFZ9x8THQtXZbTGQ6ANjVJdXKQPnAID952SmZQ9cgYXJkYXNTwlo2BHGlD
512Ey2T7phx1XVpZRf1TlAzLtdvecLieI8kI9RWCQHfXl84lCdDMVEVLK0Z3yxPbb2z+0k1D0GTW
gBcWd6Ob66emvExBFo9Tkg/BZyrCmP7nvFxJORIVqDaf6RRN4U+AFIt4YguLfMPf0dFSK3KxsHx/
n3AfdXGdkD74zFXrtVCGjuIvaetKwqMwYE7wmK5EAc15UgkUluMFKVGsMYWfqdhomdDzcn43f7+n
31xa1DZ7W1Yr9IFCZ9yOiPS7Le31OG25MJX+sJDFkm3nIh+rlIsInqndwniaUChLdTfzRvVjq2Lh
LsIXmu0NPFeuU17c5YrdLRRO92O2BpVR4Getv5swnEl+suSP3ilXo/NOByQZL/MdTqJ3/oJPCxIT
lR7WcV983LS3cD2nX9vAeDVtruxl3abMrOzOA2hvuzisDOSdeXrhaOkmqaWPb6873DS/h3eP58zM
hIfMsEkOViRzRGzwQEF5jW5bBCebuXx0+SZutwDuRnonh2QlksDgln00IyACexQGg8GB46NcDMyZ
Lzii/sc7t9wmDXungKv4Jvyqs/0xRs8GkAVad6ClQk65h0gnYbjfV2+3rVQAeV3ioMrX3Drk2Lgl
0y9Zog7WJSVbqRVPyv8f6o/yFvloj/X5SiFOarSaRvxelPJdvbKci+Iqx+YleO9SznMQ7CJ8JpdW
4uZTVANZpW9wiFHQBZhuBgqTG2EspYnbYXS9mLTJNiO+UTKJ/tMlqmyXgN7KcpDlS0cAKABZAMUq
KvC2EliaS5bha3TDouTbJw8DSifujDQDzUxrj12+S9s6WEC0PWi1skAQi3NTD8VwRfDzUBi6vaDj
oQ9E2AConH9TGG+ym/m0JxrT8uy8IFSBahlwWvf8cNREU3E5uIN0z6OjEs04aLywHJVPGVoUMoBC
fSrMYfD/UonXjD5IKQgG9rzHOogFwqUgtagnnG2q9dkjdqeqTbdoEeRsvM5Ti4K8nm67vRhSKcW0
HFTtrXcEkt+/82CG6jn1F1sfDq2uu9Dc3++qT2u4Okqy9oGZ6bvS6+PIZGSGUoXPObOpo00ZklwG
sOkJN841hcsmn8cHG12kv+bQLdqTKmSIEqzNBVp3xDGjMLNs3J0AH80NZuK7lTy45fj3OVLtMuwm
/Yf0e3YA2sdmTK9ZDk6+feREII9ZPvtCLj35Lnc0mALyB48XY7GFdALhbOtmtlQ4EIRu5QEVK7XD
w+Q6GY4UnmiIPJ8KjWjJzM1ClmpfekOLw66pNPSVWlXuLUPMDHiBL9pjebPpCJHc1Wdw/2CVnM45
k6BmzWDPCL/RdS1Z1SP/ZG4uLMyFSgf4/chkexctOot2GFFkva3Ap3+Os/hfKPVqNOsEt6O+5mZ4
qWVXTup/ZBGtCm+qQtt22I4janNS/+nX9v1/+7uqNBQmkiGiEwmWU6JrfZujWK4bhJBy54vBxVz5
zslqwavuct2ll9w7pYiuQ+maUkUnmauH0URTRqSb6DGULqQuLM7QZs+zzSIEQE+1Ree/Hdlrwo52
gvBxkENt4c8+MFQXHFUNdHuWb367CL1fa8f5FMcnmGzyOEayEOF0P2HXfQMVm1xvhp5FP7niBFA7
sU59kxDJmSA/GYlP+wCNpNYZ6unX95CrY+Jt9esWMJ7VlC0uDLCfmGNci3IXJHBCKAgm4R51Gs7u
wUc27MVCtKahJLwLlHVjS0XzvG2H5UP4Qt2Hmf7yww8tlXfR5Da0nVGfmuDnV4zjlk2GY2DwIf2W
DX7NX9hPwMPsWr4yVwa/ntnscd6oe9Cq2bCYHBBT30SYizKsjWvBZ1YGMTAgVEL/ZIlqMj7DzaIJ
by8DnDNjBkdMuVYUVvnx8IxT9kcSYWjAI03Vjnbu8qu0AcwMj+DK70vfh0A4cubYMFw98+YH/kjt
/Ibg5KmpinSN0RWqu7Y+c/9mBdp6N/4PUL5Vl2UaOdNBpPQAc74yg06sqKXpx6ZHG/ZILreGjyb3
5mO3c5xc7ekoLG7QtGTE6f+/5dvNrzcn0t2HNAYxfi6EdgYHOTpgvlltAvEuW6XUZJnI5OHTnFwq
/DdB56tTvCeBeqbcG6tWDF2x65kQp/EyvdZoX6lpUSAc/6CJK8qXNcUj7BOlnVJ2KoE+vmippDsT
LbCfD6IKW25hW9NikHn+gG+yiFuOpIDgr8NuiwIhW0bXkZgx2aIRXtwQphYT03fhJE4APLM74Gu5
DdKtd5LhOEXepHHwsR8hB5MDTSJi5lKlYc2dWB3xuGQ49vKhpaXyz8+id6OSF113g8ZfDvXXGlm1
QJeSvUz8qFts3/ITicGi9zNgT4fQejpFTnwlAqK+9H9SGTPBJX5TZcZHETQs3hhC/H0ENEKMie+/
Y5zlcUsYUp11IRsx0uG0C4y1jbE0naCmuzBdv2nFETdFh5Dq8lvYNimBSmU0H9h/xK1U88H+FQ2w
e7ZFdzEEFnbrqzNNF4gxnXZ9OiqCQSoKWJB40eQ4g9JQG5kAkULCZy9neA/1o5wVImTALFgN00g1
ko2bBqE8/uSgEpciQY/Euz6gk4xBt2EhavKdTH/Kw5h8E4Zu8NBPhdI5oTeCff/beW2l2lJvzvRH
gAiVqGA2qaHrPfBk38CIMk5a+AajxVPj9QM47teH/PyOYQxygdEV5xujhflzAN7JEod4NZGvLgOy
wFMd7AgFRI8qJXoQBOB2m7FotrceazxsgDYaH3s4wZhsl6fhkt9otfUcXYyESMQCkf3WfBeXDXsn
9EMsNGO+LuwADBkuWZ8qzGVlTVIvalrRx+AUg5N9rmCvcx8JsbtnQvTYP5xB6F+BBbD/xjuJJYtV
WsOlBYiQXd/loRc95pd3+sE6OPiq89eRX3LfoVPpdZt6S3cohut4eWWOH3o1a0rmnOGLbp5aFL0D
2wUi2HeX2/nL3gR+tjTsh/4BXbnp2NFm6gacI1YIxNHNcNrZxjfHlI8R24I05VGXwqcSvGGUMBnY
w6GkaxEgkma536aeRSst+V+0IiMtpj6guapvkwMKB9bgUwecHCt3jeAabJbno+2N8no5/yd7mpTA
JCzpWiATyVNOufW3wsnQ9GvDr0Vn45fgXSajiQwzFoxBrjUHx/0j3PtJ536MQM0Lpa3SXXLmYzG1
+mnDv5Db/G4qOpT6xXAg4MDu29Zn9bJAE20USyU0aDb4XOBvnPVzkLMvPgzJ1m1vV517CaAQRX7Z
UFBvJaXKkQNrEsU8Wie1Aaw+1Xq8BVu9BcBTRo2GJzUGmyN1N6g7zHzZwzx5mwTVIzLQdaxTxrNK
Erfd+i60I5VIvwAhep1gxSh+XwxrEx8+Fwa4PHMMOSrueo2hiklnLUGcfZ3yM4OMNvhIsUSmzk3m
8RtVxeUnz9IYSnsnJi1eO7VpIFLzRuYqN7e6qOFFz67s5Skm0Zg+M/NcWaa/4l3bLEjLypZrVLKE
zecBvCsUIkHdaFvfxCXRhIDfecb8AObzhSc17w4HBurUZ7tM7CtPT6MgVCTvXkG5tTt068i4/e9k
raSpcwbTF8l4CMaMq5MkHFAntyPV68AHRLTT8c/2FVh1sHTuZsRuCYVy1HWUDHZ0ewvzYgK7zY2/
Np5igfwb/PHuVsqc000RGDDXjEoifWt1tcroFS1tOn2v5lbmXLWmL57hyu2jfkzK/GSgyMw1T5bm
BjMbE5+rYnCOs6xrkcQTwuA9Z+uXZrpjQSbcrNXRF8oIazKQaEJGCl3JmUT/C+VFWLr68EEf1ZvN
ulDN1RZDfI/RJ/9SbmoXMjXzt6pZtsrqgZFYsKZIKJwk8/npyoTWdMRWS+WIxAPdrJXPwvj3qdsp
lkffxXKSrhLu45C0lF68DpSGbHID+1Lk5JWu2UqcAkju0s2EiEihmPLONFOdzQgpnPYDqt8ZYz43
JKh4Ak67pZcJgHWUkz3iojsXoPTzuRZ+jcT6bYhJhex3dGC1vVHLGT7zkQMeHcS5EvauVPBK+thq
QkP4m6nqRXMN8Oc5O2d6iKwXnN0oZ5SO2ekDPoQ+zjHY2jqY0dTHfuH8oIMN07Ey0auZwQt0n+6l
fiM4QG45AeAIt3n/Z6ixJDpHlX/7NwBbkcWNHd0PeEfQcn8MdSRW+V5aW8GG7i5RQoL25HkG48uK
9lvJzCNH3hgycQDV3uQW2syg3OOjVZkRa3fEhZxIs/fjuH9qMEMsIZuoN4iYWsAKnPNIhn2Xr5iK
VeOX7WlmacGVx16GhbhZrGTpIovE/hF9ZAUkqJ4l+eq10SELoHP2RfjTZaFwarvgO/P6c3ILv9xP
9o38uFxMfsyuggZkN7BcEnbTWm6bZStyjaw7jZAot4NdeHEnX9eIBMvY7Tsbgd+tHFkVQ0rRS4GO
Mczcj3R62vyXbGLubcdcdybU1uyG6Os3noRSvMQzJcEUH3S31kyJqh4TdlJ5K5yUBzC0ornNAc6E
5maHbKR6S2xrWTUgRvOtD/xPXifqvxu1lOzNH8y/kTfDgTVV2czjrVystrFK3GqUy2YmWQKT8/lo
03oZLTrXBCY2SsufqNaFWe5w7LKkQemqgJTpBHM0/F9rLCcUD+bDGhggYqdvXM/b9Ll0I0BIh/ST
AHcLrNaGAljpyrDq8rhBbpwC7sEi/twQf22YZD8Mhx9qHykwB3g51paqQdbRMGR6tNtzZdDLbxEt
5iTPjeqXZZkruBoA8dtIbW+Q6EVxzyAhWuYwXzj9NLtW1Zuw7+gySLE9n3wJSKV75B2fdAaYAhdz
K+W7+ZnZKOx2HfH8/4XZ0JmNSDKsTPUWvlwynzWdo2AWqh9Pp0yUH8GdUiwDi1SYGWWz3nCm2B4K
mFfsc7XGPbJYgLxNYNbyQP5s3Y7X/UifXn9Cy2pjs9WJyqhL8/VrZNdHVb8Qu13ZUprCgnZH1Slw
QgeV1Jqexb7IvwoKS/aWCdMo1CrTIUAeRxoKLbbJLlOWiWUDCx5r2gOomMoE9TM3tr1hTPdamc12
+2L21c91EMWke95acgnBn7b4lhO6ZAh29Ni6EdaUjwg2UaFwJZFk+jIWzl9h4yo5Qr6z/7/iWYR2
axplJQnl7S+bL9hFzaX5RrvkcC0vJOyycGYD8WiBZ7zpQN0J2gmmmkMjL6Kys0+QcX9KUEGVtSk+
Mt00tNL+epMDsUi0/ooyB+LdWAQz8/llQQG2QJxbzphD5R6GABxvY4DF4qEBj8oLTfW0VE2SeLQn
idF3z0BJTMcdT3B2Grc1WjCnU5aWD0cxl1DB6/riDCEVMbEMAuNurXDn0DsvWP3t/jsnqA9ezDoc
uE1bQhh20nDOwTqTWsmxGTanwh6a+4wRm7z05xBDR7E5TcCwXxFC2uYI0bH9RHnZZqVzJI3JeOZE
9cEsXYEm60XO7DwcFGoGRgeHdQq0WwZF5TO0H2RZgLeHEIA7+crp65t+FxEbLtIwmGIkvD96HWDD
swfU2PSiZ44Axoq8Yur8QbYAGAE1KXOYSu2iZN3V0JK4R//uUS/fDbA8fyOhmFJEeaRZwYRBaMcU
DXB+/qD5ngvCqqkJ71atEY3l1mXv6JkmKxkoWLERfWeD9VXLZRfz3D6aoAVJHlmOZSsLea+/27bx
GKPLlH46Jeco4dM+WFGOeTYhhTIYkAwKpp0FVdc/qvniMeHcS5d5b4Q+N53LSOzAHIpYnIP69D6E
WkhKoZR+ym08o2RO/lMW3rd+noMpiWLDz9YB8butgzFD+VecUMREhxcARpDvEiI1EtGQWPGdiyqX
uBu2KcyDqqOsbHK6z4gw4S2jG7anGvJlgcR4N9l46R5lljF5qCAhx6wkx/tgx+mfjC4sFrsgWPbl
rDG5ib/czoFYvKyq432IT47AnKprg776332kxZAweItUQCYQkvURj+tN+iEJ0muJuJN5WXYfZ0l8
33Oi9F5aNRaa+4EuUYuYHd3wPgQYuyNKxwb/PmPS5tSB40ueeacSwyyAESclqaGYsT72T/4iMHvl
Bog4LzR19oF2dnldQlnVG/8w0Zs1CiaD9SYUo7WcNDS7u45Rioa6efmdPIlHgR8vQ9SALzc0V3e9
nTY1o2lPTWLZhEC2O4p//nqdapamAmL1domOButJ2NK5KpygDqxPoT/pXEi54AXUHhxqSzK+ScJM
PhbJCP8uJUJFdqf06Bks2diINTmQOURFNOsmj/2OS33omwtF4o05LDDh4G1ewReA0A65VoK2qfVE
cm/HGlkpYtbZISGy7KKZ+0rpXKvosnS3G0P/w+1907N6DZz8/U11yOilPVyYjFtVmRcodmqPFwsH
RtutiOBQr9bbODFFtWq9NS7ZyHJLF1AsPYzn6HfU9SK398mV1NqpRjjlDVe0BCa55hLpRKwI9Q6u
CL3Yr3BPLYCzsja8fLhxjUqEBvrIf9KfsKHwO1V9qJnlUz5GIgY4JRU1KodOaUGflHlMz1xi9DFo
kr32rltAwPvfYiKef0ZCEYgTExXWhCKKkEUSgqI0HX9sL4OPm5fA+tSRwqQq9j5QYHu7AJKdWZU2
UULmrAo93XVO001z0euBvlMcL5XATEFu81KFhdOAGWIRaUSHwonrFpNw8ErBNNWAr0WrO7PHpZ/q
fBzoYbmVySRXd/MQUl3hw4s5+KWqJG/eZ3mB0N71Pb2bIRzGNMD9CrsRNdd65iB1h6uGULftxj2e
lXZNARLdR+4rsDhKy6B/5lhyNSQ5k101fuIM+XfvXFIUuVuS8HVwNzOtMgFxyYcT/+18x5MNswEz
3so98DqvOFYLOLJIDHEjVHigYO074FJWrxcltO//Cd5lh+Rqgho1U65pQDXup1vPwanLg97TRtD4
i81iAFx5KAcziiiwWnqVOtHgKPF665Cs2mKktSo3YSMhI4GLWWoQTf9scvLpeOy89Kjgn5d+cl/X
XI+NvLDdzlSWTjbN/D9wZx84B0Sk8UJdRQzihNAbc1msGWOisuVYpWQLKpKbp7Ag3DqluY5tWr5V
LeKwv2WjYAmVNHcugfm9aGgNgBfpOJloKxDSJjAXKhF1Dy9YyilzeYTFABBNjl0WFoOlAWmfEsji
81QL+tvWGWRM4gttSsZmXIb58DiC+g6u62uHBnvk8DIj2QMEKMJkflo/h9LHDm41s/jS0TEf3Sr7
UqguCRMkwrmNbGtcdMVVVbVpBL8AAX1QNkzn0JwBpO7QOpvkhqPrCyogSzkvlXDYi3hGMZGV1q7Q
3bgbpN3Slwt8FzVRVwmxaK3BgV/R/KkmsNyl69WGLVDdWUnNnx6v6T0IhaB6T+A6lphnp8C5iK4f
Ss9mB5ujK8uT848yTmnxvFkyUl7y/qifsg/xPbdGfXRdwBa+5xHOqjhGiEMrADrR5vuxYPZdsOGc
MaZkleie5somaMJ2yTex/pGsyWwUKghSG6wgewQ/AKf3Irm7iAQljt/B02xUqoQ0LzBJirsN06Bp
vDhMNhbBWkS/0P9EjiD2yCww7q4YUdF4BlMuIFxwG/ugitIgfyliaiAlfVCdZYZfpnNgAGob4rVw
AmwVr6+I0QRE4yEzPQKJcFM8f0YmI02ND6yJyAqS+389L6NEtO6Oo3+79HJLI3Cgo2hqBjqfLAV0
psO3RoSYYda40VodCZNM6rSn/0k1UZE5DGOalsi32aKnzMa3hQq6yPrzPyb0KJVEeWVId1M6t8r/
GST9VD11tlmiRnBczDNAjBuEZ2Z76Qv0vUlTSXeNp/DiiXmvDLWocuMHdw4O3sv7hb0Vg519juVC
HTG82MjiLIVjhno6zTltNV4JBHe+nPvB+qwGef3gEeb9HLZIo5itVnbIm9iwiRganhYRcEq6Flbh
SA/YaWLqU2MVF7jE0A2YQQDAW5cqPHFfSQEPLeXVD1wGP6/A7QuxSfEjRJDpX/G3NQYXL7/9nGui
/PJHbBMyLzB0R1jHT1nKvk7IyHc9XRnuSrirGipGNsUjwUDJdl46ra0UNu4ZimBsQtVpxyjgfnu8
Byj4+RZibdB112wAYiARHMI0/wPHGy9m8Qm3dmKAzLOOzPFqI4wuDoaL95CEMohtYrODeBPcNH7v
LNqSmijzenAYSQS75ux9r3C0PkRfnf+jCJjuHKLpbuuwypsJCgV2PO7HUAVKb4qYOHeCFTNeCKqT
qYw2Oq/HcXd0uYoWlyeUFo6jimNiZLZmF+I1nuM8/n0V4XQq9bB2ZAgH/JWqQT4at6udIvHtWqRt
LTv3c7twqwYXpDtXCq3VcWJCqsrdSm/qAVJCVmIhWjHRGbC0zaPAnPcVeSwPBgcU/M+8msm04GS0
Gwf5TIJx+YVK8p4ozNNC2RNmrTfAIiPIbrITD2le0eo/fkycJmo2hB7Rq4ssdn23ib/XYAim/ZY7
JIWTQUQco352liXjH9+fwv0Fi/ENyb+DaSpuK8Oe5+7f7JqAJKOnY3dSZBODP1qZS+Usp1bGnv+Y
N4qSEfUVKANHf/xO7vXBHy0FkwI/59+pALK6Hbg+hO9RFI2Bkq1aSa6Gcd5KfDjF98B4rcSP9Lnm
VjeOoTT+uaaIqeM8QJQ7AO2Ux4tlEYsfOdN6kfPF3N9kPk5aRnXYSNQiThPtt+pABxB21cuvlY3k
zvLZtRi/Ddk47Ek1ccrRE5c6y37O0Mosc3zO2DoZnct4lQc3GZtwSHaQv8tFOePgwmF2FxxS/LdF
7zuN8O2tNDVU9b/+UrHaUtLXD/wpEIXsk2Z/GxtcvvIdcs2b74dOoAKj8HNWqbxMooJJFy1r4Ist
IGCgLXyiOEt8yDttj+iQVR8tU4QutpanpZT2E+Rrkxzb98cSGvhJl4o9wY2w+KN4nW+IPiGWgaSu
8gTnnRz2fenu+3tZaPMGzzyNIanmoev1rQrjZPife1G22g92qo+79hhfRRvvbu4DcpqQwBtfEXs7
CftdLzILDYdbIJhipJFy9sG6kcSO/BBvnkLgXiwezcNYzFu10vvD9c6cBOFnYRLUWboH7I8LkWEx
Gp3Oo81pGDOL47dUg40oOYXH6jafoQlz06yGN6vl2HqVCiJF0mCg97+E71jEAXZr7rLwfiVI3JTv
tgFCigDKrSY15ksJOqpGIZjGp9rlkJuTin5GfRaD9SyMue9qRQPwIUtPWUD2uAgdEAsqZTLTuTWJ
XxgNmCc8if6IFAEar8byvdF99nA1qekrzXkNEx0iHKf6kWnYnABF5lI5oMcX/xJjGOuTtcfodbn9
JdUff3imSebrQ7EadTyFrhIdwDa3rrH4j08K9VOhqKva6WoxCSYMxe6942PejB3u3krZG8/UFPCF
/mS0hron94LYVvkgjg8TwE+zDefItPJBIpEhqOthwir9Z19Xe5znGjA+7rUSE5+JylOZzqIAr2wv
8kXyNLrFf82l0mLjWqlZ1zmOPimb+pOntPBME8PonAUcvSHWQBmQN+27XAg+gUi+ts2k0eTvisaD
uykEIWYXYJO9BO0rGgSDQpwuLeWIQz/7yAqLrODtRrpsZ0XpQ1OASQ/qZP5dOw31Ptc2L4QR+pUo
Mqf2HuzLzP0pzoFmAUicdZfoaG/SP5EPS7F84IS53t7ldUrQDzTBdB0vdanTF1GE2mpL8K5vCiT2
2MJ0exOZa/l+mjSTUOluhD8WT9fUQIrEdKDn8QmqYRbUS55x0r4gZp+ZEnKXVR7anNwGrmxpmq93
v63xwjl8qZ8B0z55JEIELR+sPWNL4a/48klL1Os4VMF2rwk7IdR9efLBWPcuVYb3R4+rj+yKy5sQ
ipvJXtKFSlEXSWiwJ1WZ+QvR2IMUscYWMNp7SmPlqSPPS3sZXAUulBvmSt/7UIYKHXMFkTxGgWwx
j9nQFfPpnD8K+axcYyZS5a1OgzPRb6MSf45syyWH4DuPgE4IcW/DpyHakgkcOb4/f3GVehQR1pCQ
Aos51xIiaH+AV3NmN5+YePdX+BsDQsRq3Sxlt2AdoRnIZsfs9fLrMKyS7FD14BBNhEsZA0dyuuK7
67Zbmjh7OClFTcDV9idnwSIsgWHvk5e+OXTooI/1oSGcvPeBFUgojcDSOxmpRBzUt8MXyYrAX1TM
+ytfDHxLwJTYEc6jwwkKAMKQE07QRO4iS8zYpapBUM2CS8xGZ9TrjEp1omN3PDQN6enUzJIORD8S
2ajNfXMgvN0VXwJ91A0IzBEYSOzVCrLQosn8oSRb2MVmpKO5/xScwD8UzIX7RORdyy7c5stJ52AO
Si/2Aqaa8/rxBnJRXhpWzAOJt18Pa/w9lR3PQ1pnmSKI6MJObZKALNvk+zqrBfT3nBP+qQ1HfhJu
d27f4LtJVgcRTcqBeP8Nzgb0r/s7PpbzyQgZzCHR85LSTFiMKS4ymKcxLp5c8DyIOtZcgYdx446r
XDaZE5X2GOpsIPOEow4hYnpuJOXYh9spn/Fj9UXTW7BMZsL2qNYXspJHdam4VGqjTElm+sze2E2R
8/ZDFOob1b99ck4CE/rPn2szguqC2RUqMISPUzItWtdTTu4vS8G+ruV12YE+OQmp7eDe+Os0r4YA
A6pa8ZcmBVPXqpKdEyxWGQAuiAx6MtVo61KMdGHhCU27L72KjU/ak/FacxbI8P5EL17pxZU9e2RK
xx5+8T1AY15xi+H143QJf6Xr2QqyKOXQYw31GVBsxHjDUqCMAtGQXInOy09pJuxFcTunW5r/N+GA
FDS98iLY6VDfsFmqXvBfiujUwhgRWjDoCNZaL7AYp7f5XmUz0eZQSZyoye11Zq34Jh2am7f3dwkG
PijZ09C8PA9WGK13lY4TNPW7YKpHfR4wLS22pgcqzllyqV7ugp9THNSLrLfRnwbO8T/QoKJz1EI0
AEY4ui3putP6/blCxAbKGG4JS5WoAjG675QPNtsXVFgXft6SZI77aAfRZfT51sgZ3l9tzCbk/ryl
hDRbNzDla0uKO003tIqzko45m4DZoNUsml434g74K0wOVr94k9Nys9DqsTlrtWEzuirB6gUFeWYQ
4QXjdI2sqy7wIM8GF+solCxByAHk24D1lTTbjPXlSj5n87H5p7+XVraQKo7YUzovFIdQMAdUG+Kk
pd0xWDMo5CjIC10Vi/7EeSKIlqkxxLsT9vvhGND/Y8Xm12lOeaJgjUkswIWfLPK7j9yCjQ8f2piB
EYPgXfl+bPPGOnhrKK01P4aKNk6A6qdhjelSaf7zMvg1cZ9W5kFr1kf5NX+ylUfxtd6SOj68b5og
6DseUGm3To0+J1SXZ6uM4A/DjxCg92ZuihXFMDiIJQoQQTR8GbhcKJpYyBfnT1NLpqHmFB2C36qw
JQ2xKX35aai1yQtbsDZM8rsNudZPUwpz7VTu9rrjkOlb3IMChKMFZuRqfXSB18XFczPzUVttUgZp
+vc7kqp69Jy6vgjCLg1CdxNfODQESBOTu4hYoLrJdghnE22NRUsTTc7PeEzWD5CuO8IavWItUVcr
GtCSVRy7zMUYc5y3mPnXGpUeIrnl8AhBjj9vqBkPCBDp0en2uLJ3BLJS+yC0y98IfPHCZrwH4v/e
HfvEWxCSdUTwSGG9H7OgN9E02DMKiCWJzQKyd3iD5NMmjc6CQiSoQP8vIfny5qR2CKUCn6AG/ndJ
OxHlQkczDGgMKBwL3qAb3AlGQBWC8edkmmnql8yF0n4OisqQjA5dVoUnfvssZqy/WUSAnSFYMGnc
QPXvNJpt33WzLliwx0JnZ8pWbhZc5V5DV6tKjrqZmZKO0h+xpsGXujldEY88+Y/Z00QEEcCbxUQy
XirLA0e2Y3/Jg8j4MNonwuLTMLq5dt+s5WhRl7VZjlg2nxWGfDVoiazAX7s+RabfzxyUrVBxOFtT
RlodB5O0AEkrR83ProtuDBrB5qRRBEAPt6VOweFXTxsRKj93YL+Q/sBUeppVMSb/dWTKTfCHS8y+
QK1x5Mbkg9ryDVxfoQQr9nniVlNA+A/OUIOtwLM8ob8T3qlOP7bMULUv4QApQfECIlkeoD5Bxk7C
hdTyyrLdHVezfRg3hAfOEnqZ/aE87qXGY259meWi/gltF6R1vWlSt8IPbTz41fTxfKv5UDwahxCb
Ags7CvaTVRBnoEXx7fGhuiSaHtDwb3Ao3v8KoHaty2w7A7/lr0E7ufD9v5xTTv78z/sQkAZ+6thu
2kY3dAnxZebUxroa2sExxVYos02mvOnctAGyysaDzjKqLS4kC80jGsIY8MClJiOS9WT0MYbEm+ar
g/9g0m5GGVZzdrbs2vpNiV8ZbMKxPblfjxVhNbRR7HbchAPvGZ0AwkJEwmv9F6Ithm2WK7eUANtU
f+XtLCELGGez1nCZOkBaGWDSM4nOABSe5UWwu6P7udZj+nlhhHAid0G3EZyR8XqJsCPI2fJ+cx1d
5Mt6nS+C490R7HR6VPE5MAvqZzHhZB2zc6yLB4kh8pVko5R9SH4M5/k3SWJuPgSspTdsL8DN094c
l68MchnVmbSh2LX7EflWf8MGlrXjbn1hGNlT+ObqgeytCArqFTVwgjY74wKRwGo2sYNkcp/i1S3q
gDU47wYE0Qzhy08kvG2sgaBv0aC6WwexV4ERIoNre33QtGVY6O1UAtHC5PY6KrVchr1WY6uT2RKY
monBOKHMy28vmAPjViF1TcfCoFavR2ue+6ibncx/sHFw3WXyDYmu/owjQXMJDa4YT56c0TUxAd2n
UGskaMOh1xeFv9156bTj0YAB11HfBqAYk4lQzwaJ1eEP5dEAhbosYEiS1lEL/hgeGE9v7o4qtlcc
1fACjfyjdYzFobszYcMr1BofgBpH5QsMTp+PH1Iw3a9b4WfO4gl1A1etz27LiiC9ysBDFmr0thO2
nyN3zxdOHKui2Uvuy+9dmzAyKALir+WDT6ygxM3Eq1nZQW0YPfJdF9pBHMVT6xoDiB5awkayaegK
hBUEuBs9vvS8YHxd5C/Hi8zSHHieYAX1gzY0u6sjanM2ztNGF/8kxRt8VyIhaLdTU6NZrA1Ik4FM
9JuKvZmEzbtJb72kUvA52ErzFxySF0i0vU/ahRx6PwpabTkbNahea2dPYZH+djXCNlt9BxfIOvrj
xoxRh2VyKUa9kbQOQOf/A7CWBrOJfJrh0rP7Eq4ZgZ9Sifi0RW4YDcHznh4I2sITxhzZE7VHxqeL
6IVeBOTY8ALvL/O63IxpGDv7DQDVr8DQSqZfAuXOGvCZYKKxG5P6ElhHJFUuM5lTP0vn2WAw0saL
alX3b6aRXcOUPuUQPKjUTA2C/Xi8s/zTkeJW8M9bBtLeln1gJlhBo5qiNIHov0mkmvhA+m95B5P/
AWUkmWEZ3TiDusz3kIHcqLrcpT9OLxWTqt7mnRlBSIIjB3Af7hmABnS9QI5pOhr7v3Em43bDfl/3
liDKeAfQBhx63h3/d8JOUYKYS1rmeheoSZQ1tUCfYgMB5FrPurFaBLMWNCaLiJIUYlTPRzGVlVg2
K9cKEpQxipKBeOj8maKh3K8TPT0CQCmjqvHA7kjD2ufHjRKBMZAfLq6DOcrrMau6eDPF68ezXgOD
dSM2QILpSnwuD3rbeuPfdhL89QZkJpM2S2K3J42ytTixZ5IXNNrNqBRDlTS7LJUGSlQRG+Ds1oXQ
/WcH12NRbLhoWZv1XaW+tCTUji9yw5dl9OhY2XkxgYtRcyTYVLdY/v4CEWxf5GzU0v6AasK7/dN4
Msgn6MO1jAmcPJd8Jh3f8Op1UlL9VAumeOtYQHJna+RYn+hM0MC2PH+oADqFCViU+g2P3X7BH+dv
tVmnqMvO0F6zjpTdyDwRsGXXYKrHGdUVUBg28I0ggijLn29yOWOVUxeEUr+2Nx/7PJGbLl8rqA9n
a22Bxh23BSD+9cBuCqZt4qFUlCbqfwXGTzJHONl1NP9Rje43vMw6zhZjlINBOajtHWN1bUP0+Qaz
6uaHhxcLKuBrRnfD1rWiI1KmXEAfV0+RAe2JkT4fQPJCtSirehtzollJ9Q8vVq32VCo+mD/MtdCn
eD8RsY9IP5wClEIfUYyWl+fvCzncjElZzjIIjof5ALOGoEbgU8rXmzFW9xLBAngvMA8r+2hGQ7Od
upa9jw8CWrbmH/ZVaUF5kzyivMlbb7fCnMTKA5yrfxxu/dWYZUv2KlsNi6bqwhvis7WAAfxg5tSW
Y+3Vnut4LVZQvUKwPFr7P3Ykvm5O/MeHFDyW3xKRZFmRwiGqlLuE/UcV1nxyMCVgBFShaWV/EXwl
oxJWnTmZv9wzb6KxIwFxfTF1Wkqn3HdPMQBoXJB4U6y6IgitSxezzuPm0J3qXo3l04/3SvKNJCX5
hESHb5AuTLwKQruAVOAw6iNz3NMxI3GBIFYrLBJwxLiRcRYeg0gNkyZ62nQc8PZXoCM2hIXebYXS
l3JrxqEJqN03BmcKrwRXGqgomFe3jrysuHrICXYu0rzkHE2OmAdwFA4vRHx9B7jhcKM4X4bsK7Wm
QFytJRusEUC2/49dIj59/MpmuKNx1EpWULqw56qSEVrWVPydpsQ4PLynhdEXPSp10CC8pBxD8Mvt
U9VVsYSChHb9YkTXISdacCinfO8FvQKfBxo1KIvKW9m8lLpzQS/hWIRRa7/Lg3pAWnS7matCFno2
7ky+20kKuBfrihAubteC7BjKpk1zRx8BLVXUfFFpOua3W2UQQYKCK99u46aIK1YPmlsaSd7ReK2C
i6mdLmuIuUJJLWgJuQFSvFGOwoRtaRSt6LoBGMF+/mOcPTRhqHhGWv/x78ibngT7HtFsXLw2Jyje
Wdcz7OKi5yM48asGiUvwi8R1t44bXnf4scjupFIRJACE8G2yFNZaC8QF/HNvNgpzD/SnEzDhFfES
8J+tzPLIYg5rADChERiP7fOAn4gsHuKkp5H48tumHMbe4ByetdC8zR7Vm4HpPS2/uFYkSeM5iffN
9K8o79fEKLvRBuWGrwpWdcNvYLKA4R1tGTVCl+wieIFBRkPGjhI+hmvFmxlVX2f63OPRI99cf81p
1AlAWvIVY66G+kGRtU9Q4eQIRZjqgWfblRFRpRLP+sDJGXxqFbmVN/mZkqpk1LlfJGK573RliOL2
XxW41KD7PNaBzBmNNAZh5jTzDVs7Be65A5nyomZE0+cMp6x9VGb7M3aMOV+wXr50a8B6qa+bRrwp
LE5ME8kGFzK0+cniQyDzTQsdp2CewzXtfKM6hY6cBqnVkgbNFPjxUGAZHD1xGZ4Ix/S53mz+OqSh
BEvdP6wFA89Du+ve3lEP9CROLvz0kvvNZcA8IPYMblpKAAiXyMMvGAFFgx4f8SMNkOvf/WJLBY09
KjieSfNZaPZxAXqmxbFW49bVUESgpiiQB2vDD+7whqRluEf1P/ClXkOnBdv8ns8xMjvu8MUXYXwL
rrJaPp6B0feXGS7cT3Vq59ELCgElG5BUSYn0QSFHYvm5xq1rN81Aa62wKc9CrQ871iYPapDlVMW8
Zc7b4mjKxXpNDEmheAHhhQ/+aIUhWXfX4jLotxNYC+yyuqeaCx6WFFqqpdAYIU6FOY/Wz1Yy/JHe
V+XXcZjBegVskj3jb53lKJvDt3nqBhUkG8+qkSeV4q4qW8XDnyWfpe1v5DhfNthGn5koAz/AX275
k68xJuOcKGOE71jdA7Nq5shJdxWwN5bgriTwnOddePxfkNnNxkKnzaYbFMS1FEy7dhforZw6UWvI
VrjL4bniZ+GSsa99DahnyD70vBEv0OHWusqKKCioms+ryYKo/60tLHLLXxbPdF9AIEgauM9CbV0g
1fPzKEkjR9PTg7psndwtJRyPFG9ZWdFy00f4qoz4ZiaJxJSyoTbNm7XKC2lwjXFJ4m1P6O7V/6xl
Lo9o3Vng7qANgUEYLHBjSHCN3A/duCuW6ZgEJrCfl3L3Kxscmy0JrT7XUdse3wFwtSyjMz6CJAvn
7NLjVrqb7nTVog5JxqJPD9ka3zFbmSNQVS/AgpYCFJpzHf8AS/t01HWlays/eMSAFWxHagVTWnEz
X5uJ9xAHPSojeqaAhh39KVZJDUjVoDyzm9zxmijdVI1CEyEiOfajQYib4IN371Y01+sBH7Qs4JO1
VughN2t24uq3KPTXVOp3+D50dBIGiJObuzrkSxcmYVBTv4qD6R2A6CBptM59D3idx/IVvR6PQN9h
yosZzX6Ey2l/XdVZKnihWtGZ+2CgLHssY9nff6OAfB32N0f2+bkUT9sku0IoLq8BUYLVbaQQ5daR
enSxwDr5QIKIUMxHxG9nZ0jozQuzKI69CuDVHpH+a5rNKg5NXDrZ/dMU9Mn0huXgHO8BS/WBkdAe
p/B15Thf6rd++Prcc8VrysbJEkwQhmCCEloA4EfE2RHBegf/BTtZCsePvWR0Lx8Ncptwaaq3RFQj
398pH+s6EaxMNHQaTCPJCR2zSzDi6891qX8jN+Fn+sLfSjwD5Xz2yuOBr3PnvVy883PD8ZtaElIV
uYJOesV5FNh1vUtsmyAeBxs+hDx2//39qd/kF/W1Krg359p5ctt6lOKuQQg7ARRjz08K9nSj3LXj
PwU8ul63xHB1QptRhbLvpRPcpcMCz6jG1GsOKjyZJhgjP+cnH1xH5Y8uAtGkYRH8C9Aq87h17qcT
pBV1/KzlqBsiDsrkI5n0IzcsxJmmCpoTM9ukJBBbMhGb3Tw+sPOa08Xd7fc5Rebr4WYe62PD1EIf
r8TKbzWvW1R7KmrHD5jkpsFEBAqIcuVqsze8MzS/eyEnZwr5HgMqRGgH5upPDoxPbWWEF0nUsNkQ
8m/z7NHx0MVdbe/f1rr3tCRRgWndONopsXFPBORNN+KceJUCE3hRn7wqQ1zkO6MrYz1xbDHMZGAm
cgI7knzL6EYcHZn86mC0dIV6ELQdgusILeIBv1XuSOqezd86lI7uG/7OReI8THZMaUpFQegvPinE
HFJ6vM5CExnFPQd9hg1CXw3+W2aLDtkE4M4lhNH8qJ6jYsqdgTak/mOOAZc6rB/W6b36Ioj8sITC
yZmsPuu+uQHQoPfakpO1TAkFRJqNd6pCqOZPHvxqI3JkBcOoZke5+vQni0PXCS5TS0SckWUGAeKL
Ha2NJsAmO63Ds/8Tde7EfMVNDM3duWVjTrZ9ogNOXnVCf68cRPgCer7rLktmOZ/tJGuDgfmsySdg
aMsnjTv53DH9uXYHyK6eJbafMWAkn/OBg1AknE5Lb+ejMn+xjoCKOcqRf7iwsv5vtLnYPiBVDDI7
9v2ZGJxt3psEAipeVNeuRk7V4ogtTzqM9e71hiJPv/xjqKUH5mOxd91oU5bPeQrqL/3IWqlcaX7o
Hwie+AUmCnVqxKOQjb0r5JLmvgfVNQZHpfWAa5nlbHqrvvMR2mTM0xIVbpdTLGsy7tp3L3J0EpXi
msWwLii/w/pVxd0l+OpNHizCz0hpy1QNHgHN/XDIMF/hSRC0Y7SaVlISt5w2tUKgyqg21i3N+7Om
cWltvF5PaTj1aRvZGKD8gYi4kgIPNJP4XmZw9ALueEvNTVdkFBG/sdEMOCFJuvLWzk0Svy11JD9a
z6qImuTtqa6jUHZcEMiZfLDRSbD1WHM9IdkIUcxALIZpXoBAu2fIiR/wZWPpqolS8Iek7XEBp3yW
+SJpKuQ8SNYhR5R3oNhg7SSRNGb+URAskjGKnog++cp2uaOvvACmMmSXX/26ouEx4Vik4Ae9pQ43
6ckC+sHZURtEdXuqYBngRDvk0QEHL9CtUchRJIVwB4ETdxtDPI187z0/WlYG0Zg2SCq4teWs72tX
Vnr2S+VIy8zUm44K4JQJGPco4uZug+nxwiOVxqdOfktBYfc9oZeCPU4n6ksCLJDrKR7AK4qCfGSC
69E/B1urV6C19fJiAx7kr6stZ9IoErMJ8okNKq+yHKf9CYOCd2HraJoizR8B1pNGclH7hYcIRcXp
b+IIxWPusdn1l5bk8rsIgo9RtFxVcaoFsaDwyNLqV3tYN0npWiUBLBs1WICxokGWKZTnGkJXWVO8
KKCx7xW547vR0OJPDs1z7bw8RSjK4cart2bJsmuYcdz7MOt7osZD+nFu/99Cm0FwNqVWgfjIK1de
emTn4baK5SEPT9NC7gDCDAen3eFMdE9RDSk2j0/U7K/H93vi8dgE9gnk5v0fFkjvq+/v7P5bjv+9
jyT4lmMP+PoFIxP/ZHF9r6ZKJDpo8b8S1v0UOeQXF2SO9SYBmo2+95ErCe6T2861m/dzBIt+ufbN
kGSpT1r40INEBtE6x0s1a7J9q8ipJ/bRuM3SvbsoeLTI6haNDd4uBbEcCJkzDCO7Gg5fi4vAvwZt
gnuLrT9zadIsOkd8CtojQthW0S5Qha5ehLvOCanTMF1pZYkgAt5lUg+nq58zstijWda4yxAyAtFC
7MYXTJlDRure3Du4aan3VhJ1/St5sliGmxPxxve6ls51qoHIjAJ1Bic6VCYsXhRnKcG07YE6K6ZW
I6wlvV2bGuF7IHY/3nWEIq2oPONquoGNzI29qcvDzTtM7yp0jPgEd7Mjddy6TwV8ZiDzYeL49xH0
VVgjer0F+JsAuLrZJQOcrY62qu942WKtruxk/R9JgP1cY31wnqSlwuIxrjNCskap8SSL2PmekA1n
3No74U3a5MNkzG1m1UyStL4WqW6MPGF8QLEJ243yqzq/N4cF9zJwKl1ZfibLt+QO/TTR5LDn25iq
R8g0t2GfSuN6GBCimGnTRtiwKbTL/z5yg8KEQU+2Z76K7c3YPyzRpele1ROrhGJfOCanRMukRhk7
FxKk1OS1XU/1mwEkAWiPuvmDynZGQZGdYeIfODEq1DOb+vnFdy0XLLe70M5ipLX7Yy30pJvNJt3c
6FLF1b6oxsBll7iofcu0nEujHRhPaRroMusc4TDEAkTKGaOHKD5XIFW7hkjjMuJRn3M5VyA2+ftE
lqUS9PtWfAxWE2pDmutrIMLFOqYNTRvPRKwFygqNIHBcYf9//xwPyVqYrzf8NvVZwKuEBqayIPU+
f4fzVHH6Ju6XpoB2tlD6PuYRviFeo5DTa8rq2c/BFFraBPyIO90blNAZlCJfaNp0b2rZuf0Yryu4
k9x8co1ZkuyxpxgiBYjszBpsBKl5eBXctm/VdcMHrvKP+TdnRdWr8qCmXt80u0s5j3uaJG2uLvJ6
72xjthDmOFOktlH7wBhcbLhyddPvXa047gjGCHCIWQXiXAbkSmmTQ8zsW7e/dniy7Q8qqUvxnoTX
spw/qk0ma0M35FFZXl7CfDiKwuVb6q94x9ytXu3uY4OeotwdpHINCon3RiHT6I6n2Fn079KJ79WO
SyjqWI7bP+8rQ2UgiyVneyoEACt2KYLMmLhn06KDaUn6J1leFwc/oaatYUQ9JUVleF14ETI3o1Tx
QzEp+XOpcpLB1ff+LwHQ+trCTZCgabO5WjDpKBPZls2DTYioHBVp9HoFGkKo8EJiD/z2lq4xTTYb
mbHNoegq7pbn/AUZwZLRQFvoFQz0jQloe6Fo2Bmli9eKyqsFe+lekSdTGKEqGGwdfO4dfq26TIUe
L0VpmT+ALx/aIB/EcGKGfhFJA8greO1TlGU3V73EbHo3/YVMAWD28ecGoFICvJ/nMgoCM8q+7qlm
mRT2atLg7NvZiam9zcmzXV4Ndf6i/JCzzHyloRj90J0eW7y6sr8WOHWFt4JbDU5iKhCkRgFcl81d
/WpkmWc9bZJCy5iQJVk4u2wPsX3i1JRUy4i/BaA748i8ucKJKDvrWu7HviQ45TvmYh/f0gQUw/FE
WB24JaJq47U7Cv0Vc+wZ5Fg3R5ifTb19RP4YcerOaLNJtwY9qZNdAWYbp03/NdBT11vkU4E/51MF
DUuFx4TL5dxatmfaXLRm1x15QxGv1ykfTV5bM0MYtnXF5UYugo+BpMnIfUKnhHRivX9McKHVh0Ri
zhlL4WiUh18D6G2glnjoCrbcsJYiHStJU+Oi63PJa8XqKuXl1VJfKggJsomSyeU1vigtaxmWH3lT
3ac27d0gi6jGP3RXzayIbz3HO9ci9EUs/ybXxJqR9Oh63zbK6kUb6A04XcWYY6OFtYarIWs4Leue
IHkN/pYfSGkDdxgDiG8nnBIU/bwNGXnr+zNP8d4707DO/JGroZSCli9xqAHgHyGVosb1HVoGOQ5X
WYJnispV/t0t6yqzahOPI+4PZs0YW1p54aIpHHRUZYf58XRRF3rMPPIB6uI+WirsempriAN/K0Vw
7P6kPxK9DU7Loq+bP4/CqmWBFNx2X9OYCjJMIJReOhC2GJNnUSGi1HovwCv2OMb9Np576y3QWoKU
x2q4TWSIi/MgrwN2jEwr7JkL6EHS/06ZEn2BI3UBnwvl6/SRo2L8D91B4vUktnQoqqux211IP6Cu
r/fsKLa6XuvlWDtDjjZOA2MRx3nQhFg6JAjdIy4GvcZJeXIG8lvUAGOJFmnu+CnaKUTe1msLn/pE
kPqEo3tX39tQZzcV/cpPLXLVLC5j2z/Jno9+/nPS+kRJ2aFyg/adriXh18kDJ+D8tnDgiuLiBccW
qjjQBNT3RT16aXpKGu8gawGDJPK/r96alJA0+xvhF5Qw++GYGWqpSDf1fYdrCBTNb7H5rcu3VxYP
qsXXq8FC4+QLUWysCUzD2b3iXZ9kNSXMdZuNXJAW8+OERp8c0A/9AA8zyShXE50S1zcbblhW2VHt
tYHh1OgpDdoyanehotUEguy7plVS3SKGCIECUtYKbLqUcNxeStSEyDwMgoh1HdVYUPeLKV+9SXqK
TMp30U4b7lxNQpoWS1G9n00W3vySQ4vovNF0DBu8+Ii9vPI0porO6RimkL/fRMojVmi4bUnwaaAB
qpifZCcT1o/6IMr5k3aspwDJDG2LIrVqzAvIH26vYQPfZAtrGED0dRBcaGkNR/VfTXwHvOg6vSyI
2IpV72SZPcL8p4GJykpI5N8EqGda2FnS9i4QTuF2ii034Ml9Xk75NnYAbzydnIzJEJP0H8hDU9xs
3hfruMOly3HCJpheo6FMUrWTUwFFdQwUJZMfqxSCUKm1XHhaWfUR21W67mYZCbFhsR05xKtZXQmF
OdQSBOx3Kjlc14TQrZXSDgGWnt5Qib6L7KQR8rTTuN0nAWShmC31PQ0qIja1uiZa9SyLb3Fyuz1L
HyV9UsXBnQha74e5gassPxHAg6gMZxxiNhF01TbuOGN7Lhi2L1jLRyhXIFfYOL9jFJSQsSLH9XlT
i7Vq348utBuErAqk21hnmPKb3EMuGu55Xi45fVvg/IPkrGOP1sWupUMlAhhQrymXhKj4zKj4GZna
dZHGmKgHgvq8TM6bk3DenRiL5XLvm3Gn7D2mD7YF/BlfzbYBpdugjzpoBQDIC71alfbCrXrrZeKT
/eORp45ODLbFWdbHUUl75XLT+qAWJjT+fKYIz+Wv/4jx3r4Q6trHDfQW7dVpV4iUcd2n3x4njwMB
R8DqetectztZys2APtV5XqlKTO0HFSnh+Xbcxh1sri+dVwyDjmWZqrxkePYnEoKIg3PoV9LNear+
O5fV1qoZpZHejVDtVVqMnuDCQ49AZqhXYK4lADPQYXn2e0Np61WiaCkixsXof2FNSlINqpZoLtOt
IxJg6BY8+NbGuFnj8IzxddOWmF596jH7UU2VosIuLrmadjcxfgoUHr3xgqtxe3VxmySd8ii0shQk
JqxgrM6J1Muj7A612oIW9deBPhyr8Dd/rKkhGep0gQMpfdtZcB+QY3G7f5i8UyOKXcxdpmbLIvrT
3sgXG5UAvNX5ypwMRxi9MvfLV0BNIQOIiXFugG44Mi8ZVOVDcVSIbw4LAg9G+p4Otym/NWbBFQtw
8M0ob6bF4xSIHJg8B3ejkmn8SDQ9Dw1VkUSu0Z/tUSjcQFht3lSlkWfm1PKlsw+itkCDNaBS+9td
nR2+ib1T1gvzJsibHwE/AMqlO5z3i3dAtcNn/MVYp/WiFugN9cNUufRWRC7a4BwCIacmV0lb+WaW
RoKUi3PU2OVtNmyecK+LTDD2+GXV9PNT4pv5K3at25nVMJ7Y7Zvq1dC8iVFsFIKZAmx28DQUqfyj
SUuWbyZ6Yw4H/vAEAqarGa2+UbaQ56JKek4a3wlApgJZZEjF/I8X6GtydzaxFqJ7xoKyxHz4/AEr
TJxUcCkdSKhrNR7E9bA+qzrOV3ABQSWpauPteTgcSG9sh1ssVp0BGZ/HUclK4t6k/lj2mpFTqiQU
LTLActRrcyviK6SBFh9+865r3aj2A58v52Pbj4fcrDvRySPTndXLr349w2kL8tK8eQp9FpDcmeLI
PeRjNjYTyrQrocrdIqfwHrELtYC2jOHl1DrFfnCCFUzEC5mwx7BHlJ4lz6iVKIxpLXqhqAmVgAHJ
zBBNIoMhxJ5mVku+vpDHPiqhdUWe8p6Mk8Pv8if5T44HfqpIbOSeCJOFBSo/ImYxtsEEgAixhiC/
OkK4qcTgV5fWNXc/lNJ4IapIQSqRy7btMMMeGge6EDvu++Faaygt5XE7XHvdEU5VtMui8A47stQc
3V/3Mzg+MiqeYlp7+ZMynDRxPRbNoCNXP18xulDuD/2hI/2COizphkTnczNeRTHxu0H5mdE8nFLl
PGLX0uz7nVvcO7IIZ8FXvWjmHTKNkA9WXqlwcdiuO3ymByZL6ToaXWAUsmBlgvNotbfSCCUk29bn
rXqLtBSrkVRBojBCrlS8r84IoRAgWOASy8ScqmD+/9XW6G451R0mcK+3uQwluOEPHaelBQ+3Ye1T
Aj2ypDdY/pamFkMJ90JtvPuilTAO4V1LilvAC7vmWXQCVRoWy1x+ybdNPh9YNexiE/qDSzdwDbyX
2P73erY9VBUmxr4v5qFvBLAqHO0LH7AG3gV611muu1Jj8n7PObEIWD2hY6z6m8jMaNaYkDXEWGQ1
Li7W3VYFlVX+WqcaDOdl4M6y42GWM/CoimLN0RP6R5cYJan0Sxz+E4KmxsJdKIE1538OiF8mpV8O
fPBJ+3cpNs24ykeIlPJdnEgCTaomH0oPBAYWC/dogwctXLqthL58/IjfrEUpBFlE+y1fp0vaRUAB
T7sfiossJ1AmHSrPV6wr3z3rv+B2pvLdxof638PeWp0vD1JprSTDa9xybfkmGw4UHSw2EV15Pcgr
nAf2eRtnRa+BGxEgy4U7z0NwxXgFErbIuoKfBAdJmhhTaEaiMRpWJD5l5Y0CE2eSaCisI8QSnMeQ
SbA/s0LUQBgCHQ7YRyJiSA7gLPSbg2ps2XCoI12vt4y8FQnlovedRSxNpLwwQiFnAOyOFP9uTrPv
ZAR0shVJSKEv6gPpgGh2p8+WRxFVBqINq+7nLDFYXuhQ7r37SVUHrHQEwCjZel51jP+mV3zeWYbl
v1j4pvxBhRC0tQhhzyenUf8Hn2p8RuZt1DdRkyLbC4OSGDT1Fa05uu40DFZu3FDdKQPS5o2fS4/E
mJskzaqdUODqvLy0B0SmO00/Py+JQ5IrAzG0AXyw/rwbp8fyRUVvZq/8tUU7Ex1ITe8zD1F3x/49
KPgPBxjRxvyEdnGd6HV0N2ozz/ZRdTJbK1Bqk1/ieD0rMhPPqp8pW/OVqnP+tNmy5mlWNVR7ZbuH
boQgODl892TE2pK2wq1X70gdqKS2wBj6NzaIEjvZwktMYddxKXgXM6ZROaxCxa2mHhBRjb/P6bnJ
GUc3zqoi4QS9HTYrA7uVCcjjLmldIRfDdiKwO7zdBjH1pCs1feB0dUHL3TY+ONPXhPHPo2tBnmGA
kA1bWCByC9S87RJocmR0hlHzgdJRkjaXDT1hHAYMSSzw9QxrMw68bAd5TXkKoqoUMs6agdseIvkR
tAccUMqX7atA8x8RBHEUR9npGznBkq7knRxXQZZAkqyHJ+EVKSQ6ixqC2B1Ny+VFRKD9UD7VdHtk
bsezEWLYcNjHzv+Fxi8JHPlSapkbMGs20Jkw+0RYtJjagXdVQ6XcaB98Hf1of2n8nrwhvxcEUtvW
RMxbOqj4MaFQ9oCxHq9E8UAejXTY0+BmFz25L+kRDlxS9WiaaIvjwqXBs5N4dSUmfO6fk74z5V2O
bgCBEPaJqU550/+8j/516BPumTmh3ToBCuNxbdmnTIipU6MSqpDT4jeG3h39ln+fgCvrWKrfTLuB
zXozTraVg/qY9rYdCZeVyXNouPSls+2+4gAhlM+qcgY72l2wF2HE+UNyOccqW0udLDREeHj3H9Dd
qkQtLUxNuzlm1x4QDSEZlAR0GxoRM+Y4D9tQEm8KcX7NxmHBEwOeAcyWrmApooDftogIAwOB/gG2
P1ji4vsuLERPNIAZ7gPVRuUiSIPeyDbAcCLAek558iSt4DudLfVlOLR5eLD8K02sJ2YRpmU252os
lWekvW2AAI/dggXHw85yXxf7N75D6YLRi1V4Sy1S/IiRt5PzDPVh9SfXd/Za6g4DRQnDVqjUlveH
QeNNwgt0YtKOs7n7Dc/8aWaLfihtJxKAG/k5GvfX3lYfjGGt2np3LtsGYOIEzsE9gfagy8ASJUjR
canwzdHwHw/AtiO6O90clRoVydRKPs8h05IYEOgYwlipPdjPD+5wrgRPrTkUCITx7ghSac6mICJC
rYms+crBVlm79K6tKIuLw24xSFCTWb3AOv/sQfzckc66wTDcxIV8ga5FhVsAA4RykmOi7HIhevIb
k/pRokcMoNH3f+EndkxCWBDx6VtaLv+kJk3RfRkZiXg+BC1zAjrnnCPvKVy7hMQ0dvKH2/aNq7Lp
mOUBF5FTpz+y9okJnD+sbkl+FSUr08P8ZsR3Ihvyw9TtY8BdzTDqvCa6W2NeZYXYfT2JUQuXVjJp
R2VUP6DrBNuV8JNvA1pA/u3GrmQ04fT/o4rU+tPfKIr9RFpOPoIYgOfd88Ohb55TfF/C5u4m7vdE
TH8FlFW2p9qWEYytjuy/rFBV1GxLVCOHhA7ILVIxG1oFS0c9BpFo3U0wup6UbQ75cd4HySDcHRnL
HOpj7+yZQz67GOnDlybGPWlOYKyGUmGI1t6npMAnUgHrl9whfZCqfhAZrbSBlHc2YF+kEZKmApZw
qy/e0BShSI5ulXW9UxVy4YQoJiJRtyfHTlInb/Dvm0pubY3SiDIufscXv3xjrBOTIP6Q+IguureE
GjeeAI5+gD+rLX7OTznjOdEEzaM4FWfJIB7Sb4nRxjS3fngvlmi9UWOq9k12b0Q9PllwEa6JJQsw
DsnCwvG3HM7/DlnqD2LP2btyeer+gf1XHk1tX6rvEmVlLGZhlTK5LZc/k7ufX2aDG2fkcPC8Rxvc
fqMZv5YnocORbxHW7z8OSzWWKIOjQ+3Sfa8qHKnGEI6Rn8XNrEWjv8YADudvJQmiHsqIPk7R72Z6
jBnXkkcNrR2yPXvbFM30vlUCO8Ci6mDGaPBX1SNBeBgkFp19QKhIEypmj0HVRIrBEI4sczPyQq70
3N2jTsnugE7IkCM+FNh/ildbPW+cVnUZFO02dla2tOJMI6UV2z/mepYR6LTkmH49JQV9dtEl03qU
1d7m+rXE4pbJU18gsChRXc/cN4g1u/umaUQ+6ciuCLrU6X7ZGmuW1FvjB55XDvWHFWPNL/h6Bkjn
ze1TZWC2EQWQ2TGLfcLw4MYaA34JM2iWOQzzbRmNRYTOBvt9E9RE0bQyH9WbXagQK+tSyiDtjfOW
uMcPQIfJotrvUwnzEmn8HfMVOVeMg5qN+kAQWjvC8FZQwFDYgnskaDxW79QAWJYvWWE7N20UlpVW
gdBaFyO0/VsVVKVEjJBHLfPaTQLCS4/ZuUYj9glHzRyD2nfvx6rKTFQPKZGB4YJwdOSsvN+SXrjv
9Q8Obr2pChUhIfZ6Iclg/3CdDyql1syMtv3m129VBv1ZVO2CgOd9HjfY2ZZk8Am+y6demgVeQX9I
OzSJe9kkNycnMIiOm1CaIfJpB1oPrDHt0RBTjIYWBtJATv3aOgeqMquI1ck8JxxiHLYEL25+HsJX
1U7/0r4+Cac45FomXhoEhFXiW9/r2YRyXEU28NyiJAz63tk84MlCR6BQ1OEZuOC9V1xMEATZFCfn
WYK95TJ1f7+CA7A9OFCjgokkH1Kmc22jEh183m/n+3EjZShcKXFacjlQqi0nyfXGYNgPnVWlOedv
6/FnVEZaGj3E3yNtn2Yz6xSE8E9hdKTuTVaWnZ40IhDa7TiB6hqgRui7ILqIcYsOn2MU2dE4zO9V
rcLRcyhOZxL/qh/b4xTlZwp0WqHi8mxeUQgYSxexU4hbNOBHQhDDwgBQZKMewyYJxabngwllYR7c
WPSN+ye4LWTCpaCrfh/YPjkCezvTOsARruAxgdz6yJdv7Ui7UnBJuissL+qGw++MTzhtFI9BzGVc
Ymlc394H2WLu3GSF4WzfUTMDH9NRWE9i0lgMbiwT9YE330u7VT9LUf5xEK6viW7+Mxjo3z+9TNOQ
baOakRueH14Sv+bHSYjD/iX/Vj6eP9G4CgFomxWhunWMlPTRUDrWGmj9vbmsm7GvRkvlQ1mg/7B4
kR6Pq0img4qmFtCqnOrw3p8a1nMJaZpvrq0xwsuv42FDokWBCINm1JiHmEuBzUj2svu4hUL0B96v
ud/pJedp+NBXFNpJ6StqGyXjSk4D2j2WDI4hoQjhK+zvlts6zRL3Mnj9tBVpBj5lzsUYIO9NPMmT
Dm/QkSzqTcgPUiGVO1gB4PyDiZAITGla4D1ojSUASb5cbNLv94QNKnqNYLmdRvaHHbT9x9sLYdSa
ffgXeSgJ7vpcCkh/bPZOaZnSmIV898qMoEuymFPBo0Xvuq7ZwNzvjg7PkSQk5qGrQx4KidWbYT/W
kV2DSyqfz3Ep9bAYYq78qGYXHUT3S/+RfSZ6zK06nm6todBRaEjjjp5f6sKvB4u5o97SwOjnbkEK
SO9tmsbRB/lPeVHIesAQdHslcaffRilTIJ8VZHmINWxfKfVR/3H+0hbkFAJwzFrgMqyV6CxTZtRi
BJ/oMQvbhcciVTg3l57s2c2Nmuq66+eUVFpkpmLa+Ti5A8SolhAd4ewv27VrpmIhMMvWBk1/uf11
eTLrLw3zxWvkb3r9EOLUo3HFQMyUN9CinRIwiWWEbRX2RTrh8I2g3HnuC7D51ajjQU81jmJkUvMY
oghGdaYOK1GLSU2BnNW0gzccmqtOJT7M1KknvoYPePXupz7x3k3VVweQN+GyeI1OrKtiyiS5Yulg
IOfpD25TrpAsQFy9icQk7EMGkCLcG8KqJSiSbQPpnxza6ewOr6+KKS4ic/nqlNdR13/CQsCTF/ls
zMXP6/t0SQSqT4NcpudrVaeG0olm2Th76CevjE622SFi5kjS7wdUiYvjWM39mwiMGzA+9OFQ30+8
coMkixUCpUwQ0ZWbkUgElsESajHUa4fjAWMc7H8P0twPcyrWmr57QhBcDm0IgniI6ZQRZT6xgy4l
i89M0S8nhkX+nkOkjx7jcgoy16s0LsCVdcTZW7krAq6UfA8/arHF8x4VV+nX9HyFwxuS5gWfm5Hd
qH7yKioa2q5W+YjM8kniq9x0sr0EqoH4GhRKhWOQpiFU217C8utCUgaMqCPY6P99fGldeBLXB4Cp
4YEK8Gf1ZwPHM2xgLOeqLa/r+XqTKaaBvxZItaU0dpVPNNxzDW6uma3H46fp2N2ZQqB9TOaCxXfQ
EcmoCBCRu4Bn1ZRgCs0BNgG0KfScx/iBvFtSrpdVV0EfxjtmjPTZl/Zu75zCX2C3KIzGNz60gsjd
rz7Db8Nz09qVE7+rZ4PAIR00CL0B6WusXWdnCcNJElaewe4gamogSRvx7kbhFFteHp72uRa2NFHf
qHXvA95fUXton7voLklHiCxSJSyWFi3vz0R3bToItAvUR6+Rwql6CRmImF/H3s9maHY4gukwwb/t
6U3/bFFx3aj4KTz5loc7fvSBlD4/qv82PXOy4rpar0MKb6JldiNr5N6b8iru9+iOr0kS2b7go4u/
GRfcU7PwgAgUtKq4c5RWGedLPdNCtpwalwsJJcoto9hT4uriWBfgaZWi9wRIWxqv1sVOzs20uUBi
wz6wx71kvKM7oHgQ3VxxojgOLjDwJjhb5FS2/p9iQQ0KYKNDsNpb+ocYQuaGS4djHSGstldWdqg5
u4mU3QcJAbhoGqFNKPFjsbBs19HmWMcG7+aOyxufgk3RFprMid4JOyxh+7l6heiFy1nSgKIfDBjs
GiMbxC3pYvo+XjIaFevTncwrRUtexXepFL+Ly5wVQ295LyolajYVrdFmxKzoq+qKkk5MzfjefbHr
Xf2svbd7YbssPGKMO0lSt9dMRKMITWqtQGPGbcpl4kLvOT/4X4Y0hr/fw5JDofpQnP1h5byZ7atB
sk68sA510sfkAi8UpxASJ30haLWfuC/ELOBk0k17ff4hIPENwnC6kC2LFFZi30O0TT2N+66g01IN
0GCl7bQAjei5uPHZwyxFpL0rpFSANAVFnMr/HhGXjNjFY8V42Q3pIh97JDRljKY5GOQAQmy1KTrr
Vi1tDXwv76deJHUnMcH769evEm9XnKFstf9iXl+APnDUWUGK+UDdBJoYqDqjh4culQDXca64+FQb
VTnMXVjzQIzIWzAKaFcGGGQo2YC/Gjh8fbj9zjFeLKHK4anBEewUVUs6jP5gzQIy5qRRIf/q+dzl
KJwqJJJhg0Y8XjQ06B1lcD6ASBB4SHU7T0qQ74+2yCHEplUGsd3s7Plvb2WFSxpJ5snbhXVYoFP7
cYH1GZibmsrF1Z6SyA/LoER+QgZtntKawtnYn2nis2ip5bOUnGh4xi0M9Ct9E9d4DStMkTIgww6K
jKPb74n2gFsOKNbstDmNEate0cgBjWS/RXvRVFqIoxv59cbe57Ov9iWRFo8kY8J426arSxA5fUqN
iQIe904aOgMVexHU5k5MveubIVbebB6XBj/LcqWvS7jqYHKXsO5ymb3RQez2SUguOeD//3xwFYq3
fV3KXCLvMaXc2ShHhB0VhyRVI0ym0GCxhNdt8e6cG5hTvhnRtrZqaO0zKUbNQ+xu9qWqzDPSdJ42
L9mG1svTmRzh0QiWGShQQbtLIc8pTagonGsoOrdhP8BzGN400wbVcXES81SrjlvZICuWf9Nlr4Y7
XbDKSkaQMewNjFmzh1ZoFnDi+ZDCLlcSUiXrSRve2uUPr0oBhL2NIUI40s8pA1p3QV6Pe7OYkr9Y
lnJNhZIZ01C7tDYWKJwIk9O1F+ALB3B7+cDMETWtHYu0o+jbT9fYjoS3eR1LcPot/DCl5EUx37hg
5Lx+nuVgnfHSnC7LpOg9u8csPYgVguHYepUAteeau+dLJHeCQ2LzijKGyZPYoO2qbVzt0BJoHu97
lQqw9hGj7fbywF4XmNPHYD0jWzDj0TZU92jDAA//RNrfCWMfW+GhipHo/rBMKb71DKVxf3oB1H6c
E+1Gr22FvjCIVUEaDHuicEzapnVArCQc9/5E5/fAFUsvTq5Fgb6MnlecyHDLgawLo33i0shL/801
zNReRVWtSbX6AI8cyy5EFqWvmbo6ex2jW2aIqu07bCzl9srFiA9+xpTlSHuBainNUsxj2NlFYlMq
oPYNal735DGPgZX0a7kd1q74MvR4vEgVY0iGIyC5hzfYb08nj4BysFLPwUCsxmiYcBxNnWsM8vVP
Hl7RJLjwkAY5iDOcSKeGOQOMs/R0vmQgHv1widjxnxIPiFGByR9Wzw3IAPWHw+TjppPnZzgiLaKV
lelfz7xAonm+0qyHricPDl96dhJwiG/HMRDjL2eEN9t3V9E2hHABcIg4s0mzXmU4z4+H11awJo6f
H45LxFj8Lc7tMIxhA62KZSsFU6oOtAt/NQ2jsXgg/sM1g4zy6yNoew3CJh/rHAPY5UhvWM0KeM2F
h8XtaK0DOZXP4uRrcb9oHiGd5cBV+rdZHI2Um21vvHWUbcBT5XnoYgT5vpz4xqvnEX+GBjXOOhGw
31+D1oi2vd6mBvCFW2UHRf4N4Bd1Pm3b+uQxLm9IeZuDV8+cAhdNTEoWs8Giz2FUmO+PcCkC2TWI
1t1tmsdgmp9qZTIK02a9pfv4Kr3lcbhK8fji6V595NNs3NtxNFloJsyVzXfOuP6pwOt/zepYeutR
sejJWZI4hpivrIIG9zK1eDoKpm2PcKAZaE0/P33Y9U9JKJXifLUj8os6+uW0xt9GLf8AxyZzLvUY
eheW0tnQbJB0M55CiMt+LeTq/b0DLHWz1RPHSw+PZf6UOPdPzyy11cvS/a60upy644F9uFvvhMp/
Dvj7YX410sMqscg4jcPK4gvIC11eQC67RS7b8Wgu5AS3Rw202KFdBuSy3V2ccksoKbYerGY/Ukb8
tE6Heawscd3ZowBMDCbTphFVM8sOayJtNoKE67wS4/JgyWGxHVRkuXcrgxEu8pnpAHMq/0xvG64f
6QbHnsmFgK+ddIjP3KBSordBOzqHwZo8no1jbnxNOb98ftVry8vSFjxQyqZPnthQyUF1w+laFwcj
STt6pr2baDKhM/9hoDodPbBCG1bz1Ex6EDEJPzpfKoMRPRM/ERyHAow2OnwhflvxYmkMPgXPmz8p
nLiazglpQbf72DbOh5XqIDlKZhnpuyIqy2O2Ay9MgKvfdvJ1n6oRnDnpbH/wYvXDdlXMCVJSCSAc
6/B3MPaeQpt86a0xItfBl6oaIikWoTeK/s0rG1VwcxbVtAOpp2ROlFXBNZt41RJ00Drp2NhwIuAW
gt7YNcSEc8T64bvbE0G2iKMKhILqY5VmJ8qFZHNgJnRWaKV26tBOFtvYpTpK4Z6oFf10Roqg6h0G
LhawrGuybahKCvuxFNZ5xXMhbBZnvDk/M5uTjeEHqmVSRC2i5i4dOlf7tv6ItUdBI2TJMpBOo5xP
DghEPNkpTnc51uTQDgDM4cDpRScqhohaatkJhPTq8f6kTxbMHVU6jysriDHtkaT+yAmJp6Hy6gCZ
aYDWv4Gt06os6gZYWDEDfv/dssmdZkFtVZYVb+2sqBzyVEz/xZ7DzvnZFXGM36ciznt1SMmXmSwX
7N0DwL8A+aJIN3WMZhMEnHL/vcOSQD777T24hohJK0SbB0B1wj12ApV/s4iqM/3f+bI7/fzntSH9
q1lm3MRVfeT4Lu/5Rc35E2iijKzy0jwi51uW/m1CYyLge1LdA7FWVcaBdFhfm5EM/ExESeF1qcRM
JSob/aqUk0WBDBq0TnBEDMH7ryamXkVlGIEPnS6dKO587xUJR4U6fD7QXeWRddzfqeVLxdUHneJ7
segKeEauLCb+P27oniaW71HDgOZX24CdN3cRA8o+LweuSQoPCZ7yQ8upk41P09eItvMhEDbKTY7D
6/+kVHyHKXZI0zQNPeCOoYM2AEKd41TEvQcvp4xO8wKsWH8NhoyCvbtF+s2/0ERF4AuOpFJ0/MVw
F6sano2Itd0x//bXVs8yUKKgZE6z4txygA1ykFjgYk7nWrh8DD0mFCgIKRaVk8VM/gvBB4w3O5oF
FYX9OSPqcb3TAbc71wp7AVSG+ptF2AbhOMRmHd9fVBNxb7iB9ydVAHRA1v6QGnbZmx3Elm4vQq9L
tHCcMRWG1Dv0ncRKDjdTPampQS3zSPXKLnl713LhbomMtQOG2QBcx1udBvMY1dZ9/DBWCq44tvED
FU/NyBlrYSyfpDyOAkm95GUxzLrfhOVilDHM5Dcfb7rEkvUVCf/XkMBCCUygNM1SLC3fGPPy+q3z
NyDmBCTxZ2nzpAdH6S6JpOdP9bkCLiLHG+kcRryDJ8KijPwCY/F079xgJGE68o59ELfNHJZDCx+u
sGT2ShlJaiw1GD1UgpG+yl9hjtEZFaBOmJKXfx5jydbYFz0ebYyfc+RrS6QuAZUky4Onlf+ZZQ7S
0pdYZ0eJ+3gqc8Kw/+zA9OOtV/dB8nxb37T6eWm6MKC+o9grb6SlEwGah9Va6H4RYl0C68ugdsv0
UCbXXEjqD4L8dDcTpnUhExhsSqf8USDVumU314XDCD0VYfPD7DYZlBSUiXL7hvu/uU7GZVqBUfv5
C+O0IgUwwk9e/jma9xi94Ym4vRkA5l/liPZ6pcuuRG0o0pyHUJVL+pMpZwZQjSvugFo3bN95gseT
cRCVB0ire4TmbpvIPxAsxurau04qfIDjd1KvnQ/v9a9+HodT3NZ2gK1FauzIIVw7NWTRY3uRCW29
nAVEUAu2efX8hBZp4I0woPCUURQnXt+oaXmLjGkkNqfZsXhWygMdqBQIRC5suRAh4gzu3Tx8y5h7
77akxLavEPFdBzOY7CluDQNP2zqwdQ7M162OzRizQwntmmTowCh/bxhxMLokvCLjbPpsj5EaZW+R
ztpWIA50oG3jZmtRG2ZGT+e35bvdjIrO63VacvX1la9jMxfwHMn+/vzUzu8KM5soNuYTdVlooael
lFWZN81FX1T1lHSeywuHzanLSLTWINqedtYU6YiXhVKL0UmckizW6xTxH8d7bqMzX85/sXvUso6h
xiLJcwXHk/evNs09DEknb6YW41JKIF0CIYO/AUD17OGvtkSofDQlF7JxCfRvLV6Uwkatodj2A0a2
SK8ozAKEZalS0xxBV9YXI7W0GgOYAMmmv/EvhGsmcsOLczs37StFZXFHoc6N7pr0F4XRIdk78Hs4
DlZ+n2es8OBtBggChC8eY4lvynZO9X38yG899pJBpxKOkDpapJ7JvnDZICzRVTZsJ+FDAqufMuLM
84+2jDiT8rIXxpfKlNdKO4W8FLOW7jV0oqWr6BmWJlHE1T2uSuoLFWhg2C0k4AQH6H9R5TmsR2Up
OF1cmuWEBt8KTx9GhOptHghsP6g63ip+xF3Dg0S3BXJ4T2VIevZ5t0VtM8LY4KvpyvAdJJOEeWOz
3ScJKsL2i4MBzcvpiGiWQpRPUfWXaV/3sAx0ZbM6WRLAj7gz7tBmqqyT0OzhYzMy66G+puXWIZpv
JSFvjO9N7LkeB6lNAAJqHZ0zhn87RluAMQuUnhw/WEGxSbNelueAoAYIhEnNlNTuzDzEB/XqGMeq
p0WT0sJIwm4RyEq3+kkcFko1n31QAAjhNVG0EYVT6lvkI9Co9Z04yyCKeMp1CBrLgPomJCNuOhx7
SviS0ffHHI8Ej80/afLY87MXMsliwoh9dEviBNvNiuZWNIOyoRUnqu4/wvnnAhnsz9eUWSx/OMnO
q+zU9b2dAHALFwQs7v9k52ntVSs5PIvdb1jGDcrwOj4arDSfec1FCMXLdWmqdgP17N97yFlTPw+h
67kGYqc29sYqbDAcw7p6W/jHceN0DhlyQobmPrYf9dOY7XzUZtANPMg52KCMWRTjhZGvlpajjLd6
Vx4fVVbmy6pkf4LczFgETDrEEIbo+FgIFSxH7/6QxFvS6vU1HqftkNZK9C+qZgUrvHt5gp0SzUSO
pb6XkVtOzjd1oAiN0gCM7ajKjjzf9u0Zh2DsD5w3AOx+axfax/4owF3brlwbst4M0/H6qjuPWXrq
PwnwAQ+jpeDDmYLypax9aTLXjMwRnwvde8kTUMjVmgywQPGtxRTj9Trg5tzB/NvekI1wuzYIcchY
iwm3utPes+KQIcyOoW1npv6ecnCPLNyAW6sEr558fKxklWCVJyh79Bf/u0SA96FQg9NdY90SzBx6
NlwIkTVzw7cO2//yvLZQhOv+5YQWElQkOzxyjd98yLC3I+d6zRkQrmuNwGpQzB22uKFaACqrudAm
exeU9c6EEmMyPljjj9YofRYgNJTTlLvTd6xcFSJ3WG5S5CLfZNziDQXQJ4dGJFxYPdnmEkwG4RYG
pqXxv4GZDObGNd3lWr5rLXcpHN5RZDfY/VZZDpPo7k1gzDdRNHbOWBuHGFuOhddKg20TAZDuXAPI
g5ZD4ZgQ7JPxzRMNTMTRUcvyY6o0xvnnqkkauNu6F4TlxGaiXRdUt502c/W8ro9wtol/Uit8JuWd
iaJ80qIAO7lWAI9KP2dZl/QNy9hy59xnT6MWqvU6zV3tj5u7uymoRQHhuiL5uq7vYEcgKI5a6YT+
9HJ3LXDMzAGD4e1gGnDW8WBKS9z5m0RlQCPAu6Tgs5lIV1CtylBkNKBWtkqOmUe9M/KYnZuM0rYH
ZyC42sq16k4vewNyM0PcTJlaOiuP3JNSruUjHQTCu8cOZdYXEDfT3kNSFemdO2vtElnHK6aNuxIb
UF/diLUAOqQOnl676mCo1LATZDZQ1UptUdFM+dHR9BB0V8SwK5pTBGVdlLYcxbXL0K2YAyP6Jit5
g5NhIdo++YCQAwgHolVy5Rm0DRfu0/bhNfx4TBwC8G3f+YMx5/KET9q8KyemLMmSv8R0tL4WuNh2
Md2GD73ZMDOYViNJqKb1/Aycg9c+XZjzytBtjJbQSTgFYaiTtTh8teQjcZhMxpUCUZXfnGNyGdst
lUh6DRbjBnsGUuWOvOXfpYx9roCCgihJ4ngWCLjp/u07CqJvdsnC1z7lopRCQzcl6hQ5i26xRsFx
cOqhXEcpWVvGOO02FlrZMukOe9jcK/WCL29a5EjYeCPDjP4A9+6HQt2iYFFoTqejhtZCQhmXZyhf
xSSreBoQEyVT2OXIFe68xJSMdjw5acawDf+/PovL/N+QW7LXeOvHDL890isDf0D6mPi2SI+Yobu7
aHMq8JT0Mo6sTybovzNmzrufUhTegtfiVxb/pKQN6fdmq8afsQCR3X1iFMBANNkyyX/ZB/A0hFAY
m+7v5wX//PWgGzo4cbOtc7JxDIj4I9F51B9HlDa7vWcmN1J44uw5hXd1826kUeTdBmmS2jFys0fO
Bv0pzYiyFNLiAxKtRdAulBbJwHwGff2a8qmGjYVd6qyVp1nxtQ2UKVkNub81E6k80Xe88SdIBSXx
xQwvHhh0v+MywWetKFBuirVYwRO7e4G0AhupaFKEk/oZORdwM7FaIX8mjTZc0zFnWVUNk1Wagp1n
QF+wLmatr0P92KcQz6e8UqCjIopOQj9Scz3S0bvXtRRIzh2A3lMSGYzdqkUuq+CIlDOdL6YMnvK6
C8k5+hcnN+PWcsQIfB5BGmThMnahjoPU4gzExF4sweYCFHyn3iUjIvcYCRNUYpnYBe5kYM4g4jJp
VIAI6cIE722sR4L21UVzlPM9YtIEprvXkxJ1iG3ffxiNOqVPoxLiyWxonYks2+uezRxf1wSdsJHb
NEiy143q3sB2Ppv8bHZ4sppdCRjk6IyqTpKLl969PzDba81hKv1hcs7eimbOpiBoj003aHWM5AzM
yt3XbJtqSmwLHpyVAGLMzipYbTIsSnAbrQPe4pi2YmD0TkHx0lA08yzX7ljszG2nu3bVHuvRQpqS
kFLxWJduzoYGBKt/nl94ox7qzYFx8fM/Rf8XCSrR45iGWUzb0jZJxugksAC3CuATRYIMkTqHN/Lf
No9jhMPNEh7qtkQIorJgFDrH9KFOfDtshamY1yp3Rk5BHsi5tcn2Vk1B2kuyW1zlGpQU8Qq7Zw7a
4wh68nHumzQLEJTI0UZpQaWf3GggtyneJMxyl+G7c7sYfk9agDKPKHbPVuxmIgbU2vAslgzXRU2z
fRAxHWbgyz6BWQlCWWgs83vwEM5aLBAk3wndipg53CqwxIkl/godU4OJ0DIN/Ph6rg/aGv1VIV/g
5L3Q0FDyh8Z0NOvgBNyUDKUT9jb9W+fbFqI7Ss7FAK3UqDqbEG38oyqJ88AYxpDgJ8mf4iZk0w2t
M2EdedSlj/UGhSwwpOLCRVf3tW9x6hYts3i/45hy0RgHqHUTco96AQcEmgY+B7y68Bjn6yWoCUzu
EfbcUgvsjb/gdM8cMO4q/XdvVHAzWxr0MGunFk205WP3DBALVtvlwAfxJxWAmR687x806fqSY3e6
OI9ZI0Pfq72Fw/aHT2ZCxtREczOimTfUU0Cvm30IfBM00/u11LC8Hx/HCUIFAyVj6RALQ2tGizr7
a6Nd6oJICHqMTFrUXlcuxUbgU1BLsQsDwdKJ7xstdwqN99XAjkhTlf9C7PoJQ8T4jIcpbHQ+0JMk
f5GgNUxqMhz3PbzZx2S+VPdVKAPvkz2HmgTJ6uBz0i24fSym9O+fGk9CVqnTnY4ECjhnhd99QW2y
vK6hzh3dN4kB+WJfawQJJpto6doC1A959UXe2PiMeF8WZ8YQmnuS8ZYQWah8EMoJ/Qk0oWfyIa7B
SFFvtJaSkxh6q5oCEVDjYMtzXdm+Z/VK74HgRuhyv3kXz1WTYC550TK1gDEeQ1zDBEoL63p/LrN+
d4HeqO65fZWUbRXS/pcApUK3zOSu/Fwc8VZdpAWVLs7V9kkQmZXCFL47iE0I76r9CcxYOggWCeE/
dqK9oUyhCudT/GFkRT6xpJOAo4wngZM8PJ+vPV/twDImR852NBA9v2y/pdYX9cYCle0pHJaNtyeL
pbjWucLG5c/5eRxocalGtVOvU4zhujf2o01U0LBIaMyOu41jcMDjNmqt+I7wQQbBJRZn9pYW1Hlr
j0rZKpvDSb093VF9Ku2PnSZAWzvZTFJVfDJ1xW0qbjBEQ5rIGACoSl1AtkfJGlxDDwSQ93MV52Az
O3KXeqfw5jp+JG5VKKhB1jl7BbCMx6cgooP6lFN6X3FTy6mnEAlz33IMPM7jUaD9RzE8DIsEORcL
NsUvIIk7k/L+msZWHVzSAwO9BrIIp+FOR5UK4i6oK/Cbl2CXmw35JJWbRezaSZCkESr1sSRVJlp6
5+1JZkorP/Or8N/VGG5z5a8XoG+MwSwqybXgE+sqZfCAkOdp4s3eF7APr8+jreNd41O6OeaJssh/
Mi2V9nNL64Rx3teMIEeSrmLi72Lzqgg2SIBRAZXWbEyi7asP+pDox5F/4PQcj4byDueWX1RSWZhZ
wpL6jt7tYuUFKHnG0Tf1fXI3tiIDIjLmOFR/Ivd/5YwW1r605zOxH4+tZuWp/qjeJMtE4qPMTfHi
Bill7+pksfCLOqwdZYDFsWVgn4A9X6KWTMELemJjHe4BWy5jmCAd+AGZtY9GAqoSNYz0XBRnztB6
tHbwmTiGQLRD0golGgag5HZ78Lp1vDB/AWq+LMG5yCbjp8ElmdNihWetOacNltzGS39u0PaB9nJP
Ob3kgk5A4tJ++ORd0g3KjlK38GE83lggNrbDldbzhSW/gLeL/QD/uUhAgu/pKE33bW6BkrVY6zoW
JRICioa4njgXwiYDd9KnOzv3LRTfh2aHoFJwQdAnX40YECSV1SwYb/h+q7KdxKrHNKZmLnB6TQMx
12UIb8IoPY/0YUIwxXCQl/8yqQ8tiupZIYkoSs6Irun9xuXEQy/PdtvNIRKH4kuNHByaNgLywwsv
3tQm4EyPPGGhebLiaVlyW9xKsXy8D9Qx/xwGLwBOdGfQ62cJ2Cp/RdjPrhpk/HuZHakk/tl3n9dk
E5UGjqms13/6o5DnXL1kOH8KLTL4yrcyx1x4QQlGd6cMx+i4bwvo/JDO2Ew7Xm/Z4BUEV7R/y9Em
dTE9MU0ZREfDvn9wzHX3iZCQjOq0Dyp55T2PjevNBOK04tOfLu6NdB6t0ji6rDtJNn+lowI7Fumq
4P8Rx22bkR9H/qh5iaN2H40/MCZmErkxxMtRAo6tMJsvd8RYoSoA0FH8ZSw9rnFgYnEFhqytVD98
MaYbu6PtrZMpOKPcM3g+eHx1Ye6wU5ziEt4N+vhLleLUdoSUs2zTwQgCZcwRDzAes0Qovwc9xyMD
J8DzzAEKSqed3ymkK41X3SFGVmzBBMNTaPSomfhBUw+4Ucvkwnsr6cg8iCZoNxMCIJr2lHdgesGe
oxGGt7S7HVgoVQs8OAV1n7zZ3ZY3FyBzU2rxiXGo32yOna+gu7rpV836xdfNeAdKEKBVSJbsLZek
BcWGv2QJkFAS44g67Xa44eHPRi2D2fzHlEPdxVM95+Wx45Y/FNWZ/xAasZxfKdEpQcL/bkhH9FV1
6pBy2tj5Pajrc3tl4izO2wlVHhGmMwP+kv90SzeCGJKXyBIIlb7+04sKn6ja8pHKbYx3LFh9hHHj
r/f4DXcYuLD9OGybx++ylisVplZje+X/uOm6FeNPBOAkhCbr04gPdgPWcHKO1yGXr8Qs2vUVCGx9
Yus9nFtx45UDkFzWm0oknwVX2qUEKW+EaVBslwC7o5ID6i4lKxAhgZk7Sxu7Iu1wwdiBRg9zNvUu
x2zdGZfOIwy1/riLl0n/4E1tvs+IlrBPj0ZGCu+yj9cjnnko73KCR+A7U32Wowv3gg6yuuLsU6ix
Tpkhn9yLEjNOudVaZGHRvSs3Oj821BI/Sz5+IvbMy31IVJlkp6Y4zcVp63Tg/QASwq4/QM1KGBun
qdAvlcet6QE1BexCsKvL4Nxu2W9GYIr1ukN2yMKja9CsgARVlZjFuQkQdCt3ONWetyNL1+i9rknW
1kKe3beXAMqzM146uEpsq800/z6V0KgqEE22ct1ZRzStg4k38sFKH8CfyHB1bYxPHrSeLHbVRmqK
o+yeKDtPrOqfjG30YyTSnwFSg6PKqlapgAt2Jfh4KnQ5XaEu4eVhwEOUDu8jsnChKFKZES0rsMTB
XV0P9fs11ovEHFn7ziZrrrmeaZLG1llEPheGui7/1nCJ2Q1JOEffqeHjevQa/tE9i9VEUltB2/yw
q69zfgENtesWYfx8kdEOezysxXUBzSkL4rkd2P2dgERuPNV2p31xLlq8NdGduVoWfrhchRk8pz26
K+4MxsggiIhvfCzZaKI4YpuRO7VjNQb7cI3our8yG/5ryaDKa311EeN6r/22mc2LreQibIlxowSm
+1Zn1c8gUtkBxwy3RCR6B7ZEmuLq6ami9IHGlQs9ZUiLH5/7MM/z3JSqZ9gkCd7FaoyaWA4yiD6W
OORgVMn0WgRzOkoxlYK/IeraOe+jv6KQMspSm/53pN4vtKwwZTG6fNq1Bx0y0GoJBHSlinBlQhEi
ZpXlh3AzPfIN0BOT7zyfaz8xo4meooUM4K4PzLscy0ZJqFYGUj+qZW/3PTci24sLRooSNgVckxgr
FIt/O9o92FuSDfrXbhvMabTgfmyLLGaD1M6HxudpxCvsKhONOJo8neLGWv825ErIOLk5+e3wZaMa
zLG9uccLFlc1dR00efCdlwgs81nza1LxLoYj8QMyAhrr+iaC48wLf5otcANErBVdbQx8JkB+N3Oa
5lfTxgMhJdg6QL1zjsbj0ALSktQKjrLWy7G/eRJ2zFvCP0782r6vsJbO7QNonLAVhuOIZ47C5jPp
iMoyia/D4rkTqrIbqV2QN+f4jzX8cBkgJRx+T+mRdl6NiuSLJ+lakAG3K+9Xs/ykUwZF8Yw9VN4I
a3vah8r7ac/ei12vATpQgX7BB9FxfFnCanb9INYWNgbHnkngpWN4JSIUELLS8Pd3WIb7kF0JGEO+
DAZxPJxQkbRVqlj8lzLjwNkjPkbLEZUviUYtXV7HA9gK+02IR3vNy5tGbyOjtSS7jYTlcouel3bM
Nrjs50Oy5canfACVHl2391BXT52RZMXTSnX20MANzzrWjDJ6J6n7fwWxk+KxaPYHeq/WBg7CV1F5
BplajT1232TxcgwoHN+OzpNbtFrIGpKXTYNtKzv0v56KSBkp4oY3CyFJWzP32pHQVGQU0S2AZWEp
kVy8I+MI1FOtQOa1J/c2KMHhlI0ILEuqOlQUvQ7wHpYAiUC9EK1kXb2iPdT32d2555lB+W8PU0my
+zaV88Bvp/QeaHdJJQIqvordp92gmRFK4vbRPiye6rlUa22y10MU3TNWvaphYjl4e0pc86Xu+M4M
0P/3ih4+Tt2AqiVoT979tGKuPrm7RzRDgKuZLNxklSJ8tXv6r3cEWHruO8LpWWSywhNR268jVJyb
anKRKXUh7WEkJNOcXErtkefv6J7/dVDOz8dIuqMOxI38svAClr8RYrDELmwtbe/s1sz7AZp7Q+Dj
hae/BH8PHK3RfAyVPA4ImoZ+A7GoIS6w4YK3T2aVRM7oV0gNjVJqO8SwUaITQ5zHu5Z3+7Xf5WVv
T+soBRe647ros4tPVIcs+sWO4QBz05PZeBxgqKcQqvFNqLVKdDpel4pTnblAZdXqDo0IaP6Uwjkj
7WJiopCX1RwV7JA+4h1pYP2oUvXAJ+K8eyc9gmn40LRKqkEj+/RUDlnrW3M2ARHEIO7eyehlkctB
MXVvItLLlVULOVktBkhdvG0x8k5Enb7DWivYg5YzsBHCF6+LOvVhWrq0P8nFqrbDsDShSQ2g/WET
egiLKAUjpXBGMvCqrztwAwdzO3KtbzLshMiXxwqSGyCwmWToWLwnJrcYAgRQy9FNMl/7V/OE2m6g
O+7m+HnhgUnQaIDUkqGFlUoTG5eqR7KT95sdxICevw4ePF8MmEoqQ/Ew/KtWkr8822Bixn6O+uWF
cizpbHZNVZrT3Uyj1JhMnfUNdrVbSOuwMrc3W2qdKjD3+y45fpCbGHEiCAlPUHS0j1cwmoqgTLuv
Lr5Vx3g5LW1BTcjgO0jTvyl8Zw4yk3/IrluIEzrSfgzIP06rDRRwQ0OlZmeSIWNNG4U8KHxBLE1g
4Qj61SeRZqBaP0dxhvZvVhzF1WxumjD/pQVUtlakMY31Bhtha6zWV8HnwGCCKCoMVrnnhbDKs92S
CVuCk5rfOfDjq9g5l+XXgobERq2p2C4nvyi6qI/IhpXZAchqo2pYtBOdqP72uNVmYfpVF5NRVtrS
n9PVXx72Jmfzg/90pD+HsVkZCwOQdBwmn/15RLOsGNruILf63TDk0E/zbMZBQzQJUWHwxXSOTZ5k
0YEkRtZ2nGXAeYdGhYCXqH0Hojv/jS5oZJVAocErIQi1AIZew7/tf6GEllxEyThiAvyTm8Tuwk9C
hu5x8NcVZyXlb0dWTtf5vAai0w5axqnuEcsuoxbXDhWmF0oGxU1O8XmeVi0MPt7cqyltWBjK/205
7oQ8k/D/bNEW2ioz4JId2rZbWHBkZ5UAbeCEuBmgFjmr6SsELYJ1n/jiS8Uf4weYsN+CdG+FTRQS
SJmXpBawT8stvMIWHuPB/QJVK8YIIOunCiM+CdTZcnEsiRRkg1jS/Wi/VsLb/ipTC6yHuNpFz1uA
U19+G1nHyndhEW/uYEd9pbvJ5yprE0VVwPH7rAfzKD9zVP4P/Slfi3wsMLlRwQwKtDR/c/4kK28/
3iYJ+iIvav2khN3OtJNIBeWn+1mohQqV4QYEr8xzogWIarp6jIccMiqyaPFAjXCih9rBaGOlYU52
F/lGDv3VVGpJkOBrTIeVwscpxEL39V4sf0lnL+KUl0Rh2bRSgfSzjnvCEWTVJKIDZ2dqUMYtOt0K
ZRzRm20/QjTvVToDziSd5pWP/bX6LsYRnNhssae83v3/HAEae+Je3DP8WvWhI6kFBBs83ZBBjSWM
OdwVDHZ02QFTstUtSRmkH8ZV02Y+BaJzWq+vyfzXJtjNGdS91p443dQRr26KIWJv+jfohia1N4Wo
wcyf00KjE3spn1WD5fpZ1lBCRl8SM+EeDY1Gi/YYPmH6OMDaE6YXbnO1DM5rcdP1Z/Qm7SJ2FFCU
K2TiBqQWwx5eVVgcRpafbTNoXUpwBjhRO3L+QeBwNuUNbrvkj0zgZt02SCWmgHigciu5SjyUoz1i
O+f7zVI1GgYIMB/JrCQzAORxjWQ3d/74xbpQQe2iMpWMhS9K/SBxaFV331RsdpEBZQmSAKQY6rxO
WyOTZzdxi6JjanwpPMgqNstuf+uR0bUszgNtxVBmq6aaPrqjGiZVjpmaZBtTb3NPlxQU4HmUWDsK
VjTAYjZCyprkkxbbFb2CJBk68AxNMWvKNURXydlrJWbAGjdrGjgs/SsV8CWazvFf9KxG7134YqvV
gj3C0cUaiJx/FsF500AkyYJAFhf5YBURly/G7Y9PugI9auWiq8CCCJyzwW3LVXHpBYwbqvG+pJVe
4H9GukUHSJN3kdreHd37yjGGaFD7y0FS0M5e7bkDqUNFc8YKrDEeFgTrtTfw+M9NeOm069PhBXSB
nisBEqRe8I/ZYd6QJEFpxdixZGfWrh8uuk16QazNZPgBLrOgv07LYtjiiNqnnybqZ1Yc8GNOd5as
7ZY4KZCgHzhSIvjbELSQVTkf5c/qas8WKPn+yZ7RiOS808lVDSRYkW8grlL8Tj23TYydWwdDSXOT
4QxB672FGhZI/xdBC/2OeemU+0BflOhwMNkQorRLuWl5np3nHOi81dtX1T7qGIns1QNOI6TtQvmG
lJ7jqttCW5fmS9bT6d/qgcpOoluq8xUUZ3vFjhkA6V7QB1712XsZVldP7dtDmMatgjk2lAIyc/kX
TpOjPX0AYkOayGDd2U6SlV1X/14hZVqG7m//oeZqM/NC+bBKt/FwNi56VgKHknqKXQAhAR1Sw+6s
m1VfuT3gNW8vgb0GdQybOmTADvXWXcebXHM0QC3ujupP73oF91yheoyyml3C9qbMd0bohkdkr5MB
BRMHF01c6Ed1zwNmUxJjJllC+U/DkXCcMMUCG7ap3JKHQTfV6sZeWmzq9pZbnorcZcBAWUAVBqfX
iNmOKJ+IQSkB45UPqw8Ylf8LbuQ9QtLY2OqAbwOqZLINmtS00FgHRhHNYM+yiwI52yAk28hyon09
5vB2odDJGCw8x9nCdOhVfG5e4Efn7t1XinN15ZKBoOsA2E8JCKonBhjE6D0rVejaPJxiJBzSw+0q
iGf1IejXu6SiWK88KXL2KKba0em0sp4VwUsTqQ9r7yM50KfvLs7O9TtnY8iCsI0DSEOYya4moyJ5
7wVseFzz9az3eqElwJnn73BTyUDsODP/8fKpvAOZKAKlFkyXCcEpHETMvRrF1gYgksDjJ46Afvu5
wBT1an4/V8BaCM80Zxklzx+AdTEQjmNcH4ffD4aHN5SPgcIyOO84x08rilAIgJ9I0qE7BuCeSCsu
kfI34LDBLEMxsMVR9Zsf3dqPKW9Pj5rEDOhjBJMJFqvpIUoXOQD37IpQ8FJxDVqnxwuwF0c51xTx
jbhnidE+Mq/9gBsS9EbQWQE+jd6FYGSDkn/bvbg5pBni3Dz9hCxnfblII0VP34owl+7H553gdUyZ
1BBz1yaFXK8xixk+/+GC8l2tfFTlPvp9t4BIlmThDeYWnfcTUDj5EdjvXayPNTsGPpIZEiSbf5bX
+R88D79abQPwRCZECEJ2cXcOeZ299DHU/aravesvRMMo54kn/Ey1ed1x3izWNmkMXiRGy2sOEgg7
9zo2XlNjsskVkwmwUOE1qwpPhTQdDxwLYKcaxDsQ2zfoStDcpgo9w7ITzT5tcHGu8nl9Z4bqZNTm
ezJOm65H8fhEH48x8yLS03sZzUokB5o6OO5YwKXgmX9s2nJ982CKxva8VLj8SiNp0+cHeCU0Dntd
OxZpTFa5ET2vCi6mQtBMeQP0fFOfntVoJmeIfvXG+R6T2GvuobVdHp00+oGtdyaq2J5V6rRK4btP
eYJzX9mK7SpCd89QH0erZNcQlSkDcYsuP+qRHlLtMoEYs0ySFLIK16m/Z6nj500pFKHR2hrDBDCa
dAXIu+J2TVM48OkkU2HG5IpeFooMNssyB/l1LQjMo6XMC/kUdUOcSUrCQaLGW0PA1rt2K0OIkAZx
honHcSeS2Ia1hO7QInfLv7Q20WgXO3aaZEQed0J+awEpLwDwvfOZ2j1Dv9iKlrjaBf+LyVOVcMbq
cPKfyl7hs2XLskB2nci5lAvreohluFpIhf5bzVu8LRkeFTF9IHz66eKqI/G3Zx4aWV2GzxaIkhe1
49bau6SkaVUWtlKkn76FEU0ND64a2HytsIgPoTbTIgHLiuX0fmrUR6iQmP0HaNMWrAQiYhC+2Mlf
3L4JJ3xg8bbo2RzG/XeoQbBMZqQ9R3hzR2ZeMHgOb/vust1MUNaABtFHRCJ4uPv6jA0GhUDxqfW/
zB16CpRujsvP2eowH3zM+8UO0Y2Nmie/Lm/95ev6dAjk4wQq105We9gZKSfT+8yA3nxipxj2gpKX
Jl0FrFaL+buKyC5MMpA9cx9QmEy6XCjlUYIM4dw2QNoNS5OW+1oqXAVwfQ/CS7IQ7HTOt6/tj0KG
2QHQCITpnqzfBM3bj5rRtdseJnVxe1VtuxnwHQ8GccYJsNePHH8Cm4UbsO9bSxoScalfAz7s3ii7
2rHsCJlOR1etPrh0l8k8JDUcxMr3wDb/L8O4CrngflNRoEs5QBuDIFZ+RN98VW+wR6B9n4Lzf74H
jXLQ4sOpIUFi9xsTmyDoSTjwjQbNyibjVcZH8ODFavwZqo5wwc/26JO3yt2/JrBG4Pi1fnpZQJNL
HZ5hVaAXazAzOfJV1zLKzhyqTUMgyPv+7WqCm4FxSUp3QK/GNlqjwvdrfY1TGqzRC5XFi3Sm6pP1
b+BymIhtfXtuPQCD7ygswZuFlMsp1eYUtnBM9OUzWcZ6sR879LUkHfY3rXx+udMN6J1XJ14wxCoS
GQZUvVU2fpJBXobCDbOJDY0EPuPk2PMZv3i1oYULN/4sTba4xr2gzQ5j3iU8fSQ87G7+oLC5OOth
4iBo+bgB/wS0MoYJfBT8MN8a20H3JMNg+So+ipm9bENRc+2UmbaSD79T5Nb6kz83ABnaC1fLoI3/
B9ho1GTmGaerYyOIbDC68nq9nJRzRbh3otHxzK9pHPmJEzmvXhplTSgcpamglb+tHcE+vSI0KpJM
sjIf8cCBLwfvy5oWi7gEONU9ORaZWgOQa8PxWIj2oVhx/vp2LygekarbntmWGChW+uop6WO+ZWrD
znqRsnUtALyaYN8qYmWD41Dy+sAkBVbiI+ZJGaahQPuioluFhpTlTDd6RaBthNLEmPuTXuIciauB
wR7RX/ZyJYVXrJukJCTme3tYwJw0brdDCyE36scKiS8x7tzDTVI0iW912gGa5NPbnEf+JWqALKw+
kWZySpPXACcb0NskCxXqUK3b7JIPxi5vuGrRBciu9SSoWXxDFL/hziBknXV4Xxs6g19i5TJtCia4
Ig8SImYSRkAcqvnWomH0r5lTrYUUdqnb+wJu4PQ480Q1lKlBSDrvN9bZZ4maBKGC/CpaOZPm3eHJ
bYwJxlEVKdkO9QBN1Axby0Qi8JjXTMTH4DyYkUU3Kva4yJoVl9xpaL/VK2rQC8KIwgy2kJ/YeGRU
trXZ3AG3AmzE3GJ+tm2gNk1JuVarCBDYzq/H8BlEmWwmVWbOSeDfqRmZX9bmUnS/Ap/ziKVObO4x
HvOzlcb6Xs1zBSOFzmRfWQKDFykoLPwb7SRNOLBKsO9JOEOIPkks38TFtFuu7EXLVXQhq7fLMxRj
or063oBMXl2DTvGjQTkhcPGHFP1Hh17ug51YbFSdFz7+bivPDECxXekwXkFLPo+OtAxT7iUsUPFb
mNkUq/wzzmusUJfTewcGXKEhojhcgQh0m6IAQXCxEXkk30TwPGP1Vjo9X7aZBGLDiU1UuQsmERq9
nYoTA7xm+eo9/9BOASS4I2mTNsSejFCm8YoI3b+Sc0S1HSms2C/ZBEhuJUG1GoVA7lHCUY1Ztvn2
wU53iPqMhmF+SzZBiM2nkJQyumvlif9xJjGEBIbh2tfW3NGk1QrfH4EzecA+gIjI6uzwNNOEjqx6
lM5dTYJBCVq+YCjRk6kgI+UHO4a/mOPZGtCl2DPr42AISKNh3nDmZ3AIkX7NAHJysXHkAvHUoRo5
ZEYkRC6f8e9Q84D3bRdZab5lnFYjaxpF2TIL6JL3LmE5JqhgWL4ktpkCO8zUHxCE8QO1vFa95Tq2
8U1JMxhbsxea7UUNzSPoAitKZfDFyiG0vTno1PHNwAxZKS2xwkX+YJ7b4nS2NHq02EWZewYcHDXP
SFgiJVBEeBmWrJSC0ucZ1xrZEIyMDlVpDfy4moOTAJyjOKEOtsA7SePXNtFTw5gdv0vGYSJt4qKp
VnBqnNNr/dhFwzfaxOw/xrE+GJYaYJn4z3paXjP1+sU6grbIrz5K2B4S2DJGHXOfp/UBJ+fFgdqE
GF6t2vaQwAymmYkSqQtbpBuhG9sIFde3lH1aXIY0jKnXRoFn05M0P/hOuKpTe7PzOMqcxOmLp0rx
ZWpuerr8KWGyJJJNRo9+3cWDYwHiyNa1zHkW9A7WjxkluMvHTtyUKEafsVS0pw9AlRQ/KLbu4j4Q
h/Stk7Etq+LapGoB1mZZ1fzaI14d6NoDV3mioEXnV4kRqHSnwBbOJgob9/T2PXgrYKAYmXvf+xGm
xYKtVfzPFEZ5v29hE7JQX0dyuuKVoPbSp1c6O4HVmzYRnAIYVnMB/2qhWgaGkizbxEv46r/n8Pqn
UaHL3JbbmyOWFAlkDQf+/rn++b81gTo5T9OZjofSO+x+ul5I2acvfuUe8deHF74cLkqODr0Lza09
z82WO9Oku3UhKlBCiYsBWS/GVk4jvhxTxqzrmJkKFoLdnXv7qomy27FLgTPoKjKt/jdnlT1KOL6m
xm2zt8iUdG7BnDmcq42lGJhYOPkVvRutxSwl/kUNyhzfYYa1/F4cYMnNgsWvEIvAMho/RYkGkGGx
0ufqLolvKUpNbptLZGPKNrQccQdNUSwos7NNuMfiW57SVDg/3wdDGFugntVlH6vlcfhEPrJCpn3k
pAyfMVqJ6NE8BCYEkQit9IL7JHV+HckoIZ5zUk2jGVL635HO8av2Lf933IQagvwoNcfVYG6cwiCB
81Rwgn3tWj5qkENPagzABL008M1Kln82mVHjzbe6j96x8Rxvno1wr8/JaSALfxhMQvhClG8hEL74
Oi5vuJTi78oZm5ZXgjDZ5dz+vqXRkDWRMhkVxzxlGToOxQ7KMWFHpGDwwURuf7RhZ9CSTjnK68hC
tkoxujNN7dc0h7HOSGZfzJHE3l6c9VIF3GP39EgsOUBPchJ57IIg0zTCtMMOqX7W0MUiId+caA33
zy1lrnLEhhoFpeq9IH3XGBMQ0LxmGk7pguDUIpH00sIqf1lPI0Bdg/D3zNY/FZ2KSpswv+0hlu/i
Sxvbo2cFQhhQefeSeDzPrKtPeop26Kt7gSyiC+a0BSuB2zeWVWwE3lNkDsO9DZvKEVL6v2PF7mTe
kJESvUqkDT5acojL6BKHt0Rz/br9csGIF7Dogy6vIlmeeHrvGW9y/V5u4VXC07vosedk1780KQl3
dnRSzeRVozXuatLdguMNgHYrQF/AkHRQVRjJPdaCtJ1GSK2JgSudk4pLLNEk8NJdHrGIHJEGjsIa
NH2R0/2CsDa2/CuX1eAs6suNjVHG/54PkPHaoursKOih0u0WiF26gMvH5rcSyw63KXajT432qmyP
3adpMQFYPo8K458Thm7TjjxhfnBCa/xuEowEe7s9WYLn55POK58JQ+2U6rYEo6DsAS5DFthwfffh
oUX+3/BBc7OO1N84aasdnktkHgKbwb0o/24fRAbJzS1BnU0NkoBbAP9hRHVKGbLeusA2XffoMfDR
6f0p3X4YTms1OsxhCxg/1drXw3EoS9iL1378TcVT9GBflSGwkETDyaqx9fSCc0x/09LAp74nT2Rh
l9Ke3BRnwzW7MLj8ui0wgmBYYHcxExCQ3KeokTBTW+ElmdAOK2WLJx8dQzKMKoi/KrFTER3AKeVH
8+WUBCkS273GSR5tXHOJHCi05eYCf9lxrYY8sL4a61PB3F/FWKrh6to5PuCS1u/zdlgxjZaCfCb0
K05AHBGKr4kk9fw9vLCYNtNjdFkJNi5ZdAVjifowZqEoIbybguvl4goqtotOYudDKrBkbbmr0Qyl
KKbH1Mo54d2EPKP2nZ4FqFYNrpX95jmSHng2eQDF5M8ae/qTXV1c4hBalnToUiJUXtOYPRLtEZuR
N1e+/0a4/IsmJQ7ZIdrQ5EvdBEBwtHgO1dA8Hw+wq6yDSfSnYoXTF5XWhfwfOy0Bp4tlqoEGjvQD
Y0oOtcnOneL2Xn4u7T6X56HE9jckcFhrtIbluqqNwPyzxK06k6ieJaPFQUKn7/A5aNnc/eFKATx6
8srDYnZEKRFH4g9xwjm2eXGnM18VQxmSTVgvOOI/KHJ0+S1DcpEjzM2/z03EKHN1Adm+wraFmpLj
sytxdh6OUuIK4+jSSdX6pPLKfH4g5rXIueAafwbaY1ZAxELa6qlFg70WJJwkbRHXdJ1DZbHLZZ/1
Zt0ZrZpLEtyIfx4zAbfvfI+hCB1LmZ6uvlvF36Q2lKilDtFJeYQfabPuvZKg8SLBcI5y4nWwq+13
IcBGORMWARe0PoDwX99SMdHJX9k2uBV+7vTQ/kM5oTjNUyF2axLqUq0y6xEDjHhV2TjJaZgH2W+u
7RB7XCpkmS0o/P9Sv37u2H6IUtcD3BEa3Q5Z/Zqu7R2GpgD93C3vjHmBfuEkAZXFSeErO+SUXPAa
ko2rvj8d65UPLKYbZS10oI/HOE35NMKKiUkJEUlVnvtqcDyOPgTfwTYF18zXM7LGMb+SFfQ+y7f3
OKwuF7QDsVy/7Wj4i9ZLh7q/n0NDJOpgt/UB5vxTwZyUxQ5FsMQvxe+aIirCAS56Ie5G00MhMY4Z
U63OmQm8gTFchbLa5IH0px/Q0Rftr30dsyvMLMaJE02wWJCUdUKyJ8XQzTZAqrNSB/u/USav4KZe
dFBOvRSAhvGOYtsRoz5FlZLspBoc87cRd4xgW8LWY/sUpD8Ptil4MWA/K03F+OXPaTRk5ifzMldY
ElQL6ATggyKFGaPjWi9mvhWCwXUBLcLCp9wfR+qtH0WvG1MdzwXUa/40aAnTJh/n7T3gBDWmmlaa
hmewfVwUh/ZaoAaRmeFMsUzatWUVGe5nW9SZkxH0q2box8QAlULs2Y5NXOH0FxHY/XwWZsbk7fEh
6r1zn6auMwCm1pyqnOJXu3bTKNGwmBSxZ14VYidR0c5EJH0TyUqXg4rFIsYk0GAYiQi+lsD7FuNf
Gd6HTP+NKpYnvhJ3zEDsy970zAD6TGaeBVlbl0HZZhaGI17bAkiSKqJyv+LouVbhfDayG9Zsc6Ai
rMRLoSPwb+WJdZ2Gv/l0NCqRfpS5V+EimbcvhTO3BZZO346ymGAf00xU9q/2iXi2xm2QTNLEN7nt
9lVyI8jhDAEH0keM66q2JiiHVwUmoB2FXYdQ2qI5QMNblmQd2PHRwUYw8U5kRC95GVqUlEVsLjsK
VAqItc545a7hg/7caN8Nxm8YzxomMutteF3j8lYszoqW2APX5TEitpmzSCvuiT+c6XA1aWbEZgpU
GBFEJZuWoh+TZPtsRn2Yg5bJ36ku/K7claSXYRSsIE4w0iBpT4dhVnNkCGW2kJyG6qzuAL+iecQd
8WGkf0IC+Mh27dNye0WDxj+n2sflvV9ou2WW9eea/KY8zpL6EKYEdxKgLqNlUb0Jc/iJ99iXlu56
tp263W595nGo8RuwfUjoXRI9xMvloUwSNbgkai99XdZvnDGTrIBItj5SqXyi8nghWSoYMFOiNYGk
Cs52GWTkM/CIrPnZlt9wsSlgprKh/zeZErfKpAjyFkvqg2W8oOkMbC6rtEYAdVuOt/yZG5YdKlSq
99of8Gq8kSpeDzZq2Z602lf+CUK72wymZH9YZAziVMSC2MnHSHPqs8tb+DQ/ol5RafdDqGjG8MNV
mwoPIc3gJbXD660950hqEOij4l1muQWHCZJfx9pvcwjcRBHyT6SwuRHkvc5Z48sFfi4lTmkW8QGi
XgIJlDhEiENhwbxgLINd5nfS6ZQbxVX9hSNG/QgYTrscwc6GzR3oNbteZsMS0kCT9GumPfyZ5E9S
dOt70pQ1emwd2AAuH4mLlwQ40n+MhUQQh+/c7nzBTfQrsLXY+ANVFVlRmRu2tS4Iwel58/+1qQV1
NmjHLrUKw4UjxzaooxeamoNg40ec4W4mppN1eauoSRPgZ3r6HqlTPgtUrZVtiyOYrQf6L7jmEYd8
ZhxURQdZRs8Ru/QY26F4RhRvGgDRihcSizU2KnssNGkui4IcAdKKnYZa72FV0z174qHcGWSrS+dm
FtgdUsdG1MWWL7j8LqqVVFgNYPS9ukxt1qDxlyiTpK+Ec30IzY6SnQz8pYUaGCk8vRWAvo95rlZe
M1HqASH89Pd1ybhyfTk/V2BLgqhwxZZusQwJJiarn+tija8uTsnghw91usR7HF3tM5s/ka3VdNI5
K1Jiu9DwKBcQpftv8V1VFuYUCY4sIS4kzlO/KoX5q2sF346w8hYLkYcfIigS/V/xkucCcX+qfZqC
eF85doG/1/9y3T5U3sCpQaNwbfACPqfh8K7HPgnF/jfBm3dVNxrjrFUtr/oIMtlSC+1ifWqjwe1g
1D584YJl6RQzSllDisi/s/0/o6fbENDQT+CiQ9lgsx90ulXbBnlRXGp6EJKTMCvey4fKSBxpDz2I
3tPx757idRoj7DMz1ESZPsnGiIJkq3cfdLA3Zp68ix6epgYRTGfQOpwTrm6dTqXKTbXGdpnZUFg8
rqHORI6NJ5WcMJdyYWoMuI71efVWnQi0Wmt7u5Ug8vtGXISmMWFyGn4R/8tKrmUZKdCHwqbrUDmE
A6CxDZ1sNQjYNvWfGpPV5ikxVLvDZe19KsPd8wgoXGvuTjkmnespylvJBgCD7vbE/zD6xnjtmleR
6UXaKuMJpUFGofu8V41iCvFVE6lvvBojz0FvL04izE2TKzA/539xWmuEFzHoArvQxuP+oqE2yLbW
WUT169CVdDfh2UCP0NrRrJ7Sz/Ca8DsbQo/9eqCs/7CqWNxsaYF/1ediWDD/u+HVAKNFLIlrjCya
xsS/uOx34a4miugm/4q5Vtu4iSnE/2WgpVbj8nYRJRtKO/Nghli8upZMH+DoyG6/w1i9iMCDeWKl
RcSDKqTay6xcugpqM21jcs+/eI9Tr2x99TT3IeVHavNAGwSTtXwSicOwUzyUNa0j4NzDmMv1n41Y
v4bqIou1ogtz/wMhKV/FDfcbkWtMcWUcMBqdYXYMYY7qTNFlG/8WsUdIwimuU9ZfolSyVQLjfqBp
RsEEHDUAg0aDZ/xav60G5TCB4ZXpdeLAKX4Toocih4NF4eKRydUSzuUZueeSe9fSh8kPt/FmH8on
WwwIg/hOh9yTJTDTGSedF+S0LlMkbo0gdPbk3txxgAtM4W/C3vDAoJVQgagCS+j0JqrrIOT5wVsD
g5Qv8dhN1/vjiGtBghu2sCH4zwpczxnqFrDIxwxyr2hfa1wdi9dLK2ieUE6vSVdiCSlGh36kdNmn
+rCeajGYe695yeRlBqCeo9Wp+UXI6TQo7EUKce0g0rA9nArQfLtJcyoKhjWUZanctMQFgZkwiaf5
VmotgBdg2/GY3GhbolMWI3YhcMks+OWmCzXWtBFEhhZ+KtT7/XXVw0jGgU9xBUM7dFhubaaaD9kF
a1cX7nEhMyGot+tUpNewN3kh3KhzjF1im10zLIXyRH+LQaf5Tq+vT58NofPUIsQo5djceDWJVYzU
M6sAw2IcncWx1m4IH52Ls2/aSP9Oxc9+e3phS8UADSdNQUlWuw+QN2wW7lR9ak2lfHpJY4x/cgiV
X7KCzgqRWNJzIawJqTAdlGrnVC4iNB0VeRfFfjFn+5ueWMYnCjmXAV78EUHWdI0ICGAvlb1s2Ivk
pb6Q8/seinw/p04F8/uXnAb0i2h4VKqdT+NxB7/ISVtr+f5MrKL0NHDKQJCf6cc5WH5mr5EVvtxr
pONTRTJkuGdrh9yS/7Ij+rrv3UjEVt6cRT9AoKPCairev7fDIWpUhCq5h8WiXdE1nPAK1straTQs
tsZCa3OGVlFt8r64z00CjPH0dLk9iiZoSg+QkTZIYcbLA6kDq8TqBKZBpU2lYAbGE1aY4gZEtJjW
DcV6hv2JtCVO3oBV354DenWqk9VEHLPBKNg5qMoOMHjUqynPTcb8kt41hItZ05C/JwA5BssAzRjB
YeaHPn9Y4pyA7jUgrBNwknR/BxOmYScd8H1PaE38u5ObTVF3jXfaQHajOgCUxGpOwQj1kLGqHlHs
SJjuQOp8lbpsyXAK+XTuXiM6+ELLR/YsCZJnbUjZP+s50zef2Gh1CQidRbB0I7uSPXUcdyQkqrKm
Ch6kuejT5XZP9mfReK/BGw+cgn/sZyeCzbq7PkbDh1RUguTKv6MZaAmpidywz9XsKLsSimSiyGqP
/hMpGFHN9BzGuV5sySz5vyjmPjV/zKmxqgfhEGbvCAYcpleRTou+63fS+moTvf21aEwPKBZR1rAr
X64xFeP8BpKERLvaMGRn/rcEs8CaN4m0tNAxnDxutHD69LPTepT19NB1GCv6vxZomiExrE1I3Wvn
lJu4E0BfD5Mpvyq48tDIFofSf0xvJK5pj9k+KcFKSpdpT4w9lH3zGR8lWDauF8u13VzQoWHQGW0E
dE0HBDsq7rdRIl1ksp7hXh9Z0S4jWWx1pCs8b9NkGduPdCqlkkmSNMNF773ucIPvUt+ua+Ov/mqj
/8PxuFJgvw1/lIhBkWKrFmGzL37k6Vlm/+54d6ef7eNGSqWlndvVxJI8vSj62YoolhBygdj8VmJn
dKGrGgF0xANHVyX4S55LdzgHUsDhF75PBmdwqQGl6SEu0R2qC3Oe5ozs1kMIdFTVPhqo5Mpy831F
LtLhXxPiTsGmhgJFGy6XcIQLUrQ01vbT4bI+pO5qOGiwgqZV7Dm10DWaOH9r+rxV0oCEvzrzwl7h
gF3ov02GeLRwZsP69cJviC8jw7LgAfSTpvjip6UT77/SZHCBWFfhbJFhrtuOxZI5Z6kuBEo1HNbx
K5LIJUTnETNQlEPy4+NHlm8cem+X3bc6qUTReysUmxcn0vv+9Pumc1Ew/RUSxNSn4d7bqnb4peIb
e0YSfUQGxSt6zgi5s1ycsTlasZzlNCs4M9M+kPs08MEg2ECeqSSzx4hRoUsgHFqzl6ddvuumNft9
awrOUT0X7Azvr6jcGic83dzi7S+G5yQW7l87Z9m4GOTZrAkLNI4hZge9cVODmmP4uGLtCNq3El7L
ycw5VOYUE39d1xcsNc7F7NVkAK0NvwddVJkeGICzdUWdZrV7aPEAiGe3l2qqRH0jYQXl8SAoRs3r
TuOAmw/sCyBs6N/S47lhEpIPRHqlh+uLAYQDpnPWtDmAHq7ZbAqadnCpMuKSP+YzHKEuCE/2vbiu
yU4LByiShLgCh5Yh4XLJzEnZYzSIOB2Upcrx8wr4y0l3JlRZwIkQ9RdNaKQD/rXo83YwZbsYAZuh
KqK48Xu83D666sOlZPBPrlvUOQBoXNk2gHSEqZ/XwKb/vuHfq+tBHclJfXbzXd+QyLcMRBvCiaky
cA2qLrSyhoGSWxr325ZOjVQ+MFpWfNlUukbld1m/yWh5MFurjg9W06geSRmeZ1P2HNizX7ZPwfm2
JC+8NT/nH5h7+YLPiP0ENc3Ife0uIVNp9y6QFFSUF9VyWgqRgbHkAz0i+/5l54gvEEW3qRgnDuPj
AQdpOgRDSc7ii23+O/0TrGq4Gjpi0jVoziXYf4W1Of8zWk+Cq1ksx+fLlQrnZN3Jtyj5Mbmq+TlQ
d3jOjxIu697YUhOnXzSDLpt6cm5DrA8FAtG3LJexwTTolTOCLCBxzh5KzTi41IDaLICDfa5Jj74X
ZRm2N99FJhmusWH6tWUivzrLujf6oHd4nKeB8Q8HSaVkDa0nF9T5VeVfLhUL0TWkedKsM6mUD/Ew
vvc8J+DikV5/JiajXOwEab2JKCBEUPSp/AaW1C/vZiSPG5M2w9PJjbUMPL81i/ZaiWi2ZmHoLUK6
Ob2uXDie48Zvo6ZllTl8mhdQZ1i+kICtlDygsHlJoKLOTclr6pkdC/9nxCDQYtKEo5epWT5x+4tA
9/pABMxejdGxPANhCkGxUCZi1tHRSfzW5ooO/5vyjvIGjsXQOXa2rEu9yskiD6RUqVyGHTguxxWJ
otL0BaN4zzdsjVM9Q926lkx2O+jZ1nYD05Fs878ZMAnUmc6cN8GRqsV4EZ0OjCUDqIOAwMIQa3UB
M8qQj7n18sH5B0TqWWYYNleGpwclti+U0pHGjI60yBYo/+kgPqZeZv3JvK1BCiRbpG84H9hKx51V
/g5p9lRDE6JNAb4KhBWEvQlexP0NJ2CXOb8zJhEA1BWl0htAM9NSfPxXv9S+/Y4ochfA0MQqrhsf
2x5no29XOdLkv2UluKwEFRRHt8clsxCnqZPXyDWPeAxKCJI3eNbu/zap6mrHc79cGdCt/rPkr4sn
bSCQ+SRqcmLxqZ8wudWZLY79WgiNpE+lCCw8mqbPKvM3o923J3tcH8MXFuHXJv4gI18smwBGTbkx
j7IAQYqSL7VgtLTTB7vET0yhMNGPKxFCx5Z2ezN+pe6rEqxF2dOCsfFp/YMhkFfUL52lrbCkztEg
TfoKCzgMatZSorW8UXatR9zRBWilizaZkqvxZp+Pc5+kI+QK+2Y6Sr1jwhZ1U5zmPtNsYSy4Ufy8
Q1zfT7hkbbk2ariIX01PzXicQB2Idd2altMqoDNU/zJXcldnsPICDmtq3miwTxvD9xjgJ5UxhmzT
ICvS6FKg2YX0a9Lb2jOHBcrJH8Kjsg5aWXHOUtUZ4TILC+/sPQVJUqqMjG0+9iaVaaRG/a+KlsJR
Y0806bBT4g22jGl0wLLROCr5woHFMCCVzcbCkg8gmv+yrMRmnhnnspMn5PwFbG00zXs7Kas0Gb4s
AqWw2zgtfAI/kvjQCa7riaJj2voRACRqw7PaVvvtH8VkcZfAJjVDuoYk+esBe8VB8vmFn/bFK3QM
zqVZHsTyU+bltO/g4EnKSb6F3LmC75b3GtJzaJGxJz+iktVejsM1Yz+0zXA2qSfDB8IWfq0wv0k0
sWQvlNcvDWDdhSWf3nTxLlnskNzn5fE4qZOTGN8ghf/O4iwYRTbPh19gs65lI0xtiQzQc90Gg0tZ
zYG9on/1LqIuTcr+2zdeAsdB2L06CFnXCWxYQjX19h5znMfgHomG2ltxqcZ3jeXzQ0uf4+EvCxRp
uCl5Drhslcrg6gnY2ljYueiiAK1yJ3ez5fgR+azXKerDgqAUfSQDIOO8QIUIMckhpVl2gtrqGJnH
znRfZPNvhTg0Eb9RSDYhD4dB2Wwj3KXnVZ37IBdyIkpRfaF58FBUtYl1NW5mYTfSCyxlyLcfj/al
Nz2R6J5HMxoK3XDxDPa2zx7nTYdvbem0lPEN7qV0hXDWICsd6Hzr8Je5gjvxkxHW+GeUB90N8s2W
g0uP8Iy+uCtYjvTUNxDKKWrvqd9dcm9JDefAx5/HlooVFUZqJoQHWKQuSK3oy5y/LTi9NcygTnYB
vwAeoNDBG8gpw87M7fwpgsGGd+3ieI9yop1Dcd4JLE72ZQMVUO1+OKPaG097XNhySuUlnWOAoms9
Y1osHZQduYjbtlITToKHM+pe6htcb7eiFVsaHq+U/i6LeKaNqqY4WSrKfV0nxeCqxskg0ZgAs/ir
wkwoS38JWYYHdDnPCB8DQ6rPcBY2V+ah1airV+2PlBHdM6Z3HDDtXSA7BCSUi6V6Qv0Csp6kS1iJ
/04Q2B0t9ovhRRSSrs22EPsp5R9L+Ale/8+A5krtnUHi2xrQ0lz1LmgFbGZgmbmYRLN6pJIGw15+
gs+zYe5olxBGG4jNe1ypDR7m5gTl6dyPYFGMV0Od6mVbqF/R+emfDSi11BnwPdS19r0QF4gigMce
b0ovDe/Q6PAnNqIPjzjxS4GMQmHrXrhAsJKEuXZ8tMSCBtU0CoBYHz0WX0uqdD3iFwMkCk6o2PwF
T7sDT/re7t23mPRRdsfkefZbpGtL2uUp9IqKXbaYlUSYzYF23S+0DU9cSOLoFIXz0IhBMuQ4Z6ye
1Z2Eh4x+Wen+SqjDPVDcR2pwVUwGRh8l8GeGCyzn8Fduo6TTUiG3meXUKDClbCmjNwjCet/xrDMm
38U3GL2GWB1c/tI7tAcJ2guyhc6r7TjSgJ3UCxW4WMCUQdTPoSHvpv1f9/yi/laHBKboPLyqio/5
/Pruz9mL8nWDT2/FzAj7opFwXEeVmAK2LFUTyTSpa9p3J+u2pdfpQDfZT0FywzeBo3zuCXdKQrGs
FJCOpA0va8LY+UCnR4mfSf9XRgAb6kCFBXoKhOSyuDmMupgZ46Tt4YEtlFRubt3IEQiEKlSthDlT
abId1bfGCieokkKfZPPceO7BdjJCygw8dhWzglNx4Sh2mRGZ+/nufWd7eiA7ckyqB4ru5wFpFNMa
5SA7ccmxF22seNqQjjeecuTlGJQpkqch79vjZwil6lX/P7j/W8nK5x1Qm0JbLTUNjKQNA1fn2bip
eXhi94XYblvK8gLLqMSFKcM08wz3o3WA2LVtq5APXAiDarkzFQ8NutJMPxX7bynSnId4lR/SnoK2
DdT2IO1pOUSaeaX6edG10UffuMnuBXeDlE5XHGD82F7xI7iFAnuoNdsKi6KOtrOJekAxsPFVeLim
Kwk7o0S7HZSCkNQq/oUKNGJkuI21bqR5GDYZjlvBe3n0MT513RtgabpBh5Tx7sIIm2CbYCAIVALd
IUEJAlQYSvuxv7Aje3nwbkSYeRfH+FfqAtzuxljU9pupQEtA+YKakh5EIaqkpnJDBkCadgGmyLDo
2VL358NF+pdr/uzGlC9BVolgngEfDSOmBJTjiZUgARtowGIjZ9+HBGzXLwOJyRKSz8z6Mc65lxbp
r2LNiajlgSRa87CNnT/AighwWB2yCAEmr9K2N1FfiqJNhtoK/CK8PR7PSfgjrkdo9BRdkTMoXRG8
VQtUsYtl4Io3nFrBMJFzSAMfzq6bF7WsyjFRnK7v2mjx3BsYIhIuqFxRv1R9+VDcC8JiQ7XeMyzK
tsqgSRlrqOd45Q3DsJYIJd2LaYasUp1DhbV6Jjp7q2mEa0w42mDj7IbruFHS1mC73aMvrjnsQ7zQ
SfzBsahvQENMeks0qgUq5hj4cAuRm1274JvCSuPxYZMLgN+3Sg1Op7lPn99cVnjll412G6sQy0pJ
bvqRYqidHLzydL4Kk4whJHqeqAacGKefubVGFi3ZYRTFY8Q6ib4DkRvXt41c/XYawk8aKE6jnn54
RTk1BK3uClP7SdZKDvbamIfKwo4XxJ26wF+voyz5RnFsoZK0kY/sAXw1To5KAG+/7m0FLsDn1nBG
U7vf9ZvNouSGDvJGKlY3ErU9yRJH+RcSQeUoQBtTzQiSxHVq/WPaarN12i8BsRVHjZbQVlk0Cwk/
JXxTFm7p9g8gdvgPmpGL94MfsbB2dqOF5xT5rm/r9pUiMuNRFku4ZIMoOVOhtcQlc39kpOoUQSDO
LBSQuUChc7llguwKVcbgcJPigpIMy2PCqIifLStvGe1ul+KrWgHVO4fcgWuWLx1QtmNzEUEOghLq
A/nMexkCf2fNDee/mHtGtyEujzKeKmDsAxowwaNGoHrvZ4HXXWLA4e8oeIgI2E5zJeMYlVKG20v3
L90PLUAvzAbcD65e3rtrKHzuRBY24jSd4QqJduoLlKs8yE4EE3VAF7ZwpT0GvDqGqycHA0C8PD/3
6qigROrlBbIEEsUSNoiZH5+lQQOTFE3LhQc/bZ5csh4nBKqAMVbj9notaG6M/M7bN4Vp972G0WzR
XHGc0R1Oe8VbLIHf/K+HoZ+MRggy80AwkOBjcvZoE2f70ArXpM0/eIf/QOp4DiNiTYTGWikuJR8k
dFGZSlc9zDqFdD6ukqCwtq8rKNtxaHVLy4weyDV0H+JFzro8Jd+dphwsjcgehp8sMnQXBE7UCY6Y
6MqmrTbdQVmCh8dyxSm0t+H59ojD0x6BCk+MChPUZEsFfemIJ2OJeNh8dOYl1xAxld0knZJzCbyx
Rk1kCLm+deBvEuGhIaiT9SWxlKr/A5fEz2JyMkALtxPakZ+fJuLPhs0RUmAGHpuZdNhumsvUEDhK
1Th8Yi+YjaCjZ6cPDrVkvsq5c6XYSShESYJrIy8tovjbKrnwFLpfNaHlFgV+4QvTb9hsY0ifhpMT
xCeL/dB9hk1Fozh5C2ZP9+7aGZ9sWSjO/rcGXxpjUaFH0yswk+uvQlDpxZkiJNeNCJzo8WtPjDlo
wjtUtVOy6atVSfSR85tlYTaV503X/iUykaAPYBmzb9TGODgAgXmKe+umO6UtARlMaWylWMClpuA4
Wrdds4lb6LLRbvH8iWJCjqt1hCKf3zXcTpSdsIgGbRDqmp4EwMdEXZcmmbmPKvGdG/UzK3ja7fgx
DFfW4lgekipeRpXOhsyR036GDXqk2GqwJ7qsbvsCJZrjs3yoHYbL6Xeg9USYafi0cxUvvlURb1Ec
ZhBHDkkLvK/jurucCx0tJbY9hc3YhtoWIp3lx/H5bsjdiNF6sSLUJgRx+ncoYR4SIxCY26H8UyFO
n1Q+fHAZiaq3R2iCleUxL+8bmcaUyh0dIOXu8Bwc1ZGVe6kDqjVN4OFHUcEuPwTsXbmpP7i687my
fn+8CLM98CuGqBLsoiKd3pvhYQjCJwZMlhpugnzeFs6jvSMG4O/xJ79AEsua1Cs2DJwXfhap5s1+
FHrtlZ9erERXbnuOzePl1nSe6oUv3ztUqQB4EK5/qcPj2qeYBjTtdymJieWZZra1SedWFe9pk3QR
R06jgx5gCoCQiLVTJ6KlSVdHV7b8Z6+m3MeyhTOzAeqLmxlaqJudldthps6AcRi4kN7bzqF79FAi
G0Wp8YC0++koF+KTy44OUFGSuAR5NY0+77KQjGCQ0rkEVOmMbcuIZKZ5jOX0Utc0R+8O/JHowGYl
kTuzoLWppJQJAnBHdvBUonuWTNhXHa3d3peVFofkNE9Q1xiQQ6VBptLnLXW1/5i6nVp2PktuKbBu
sajV8XxzdTIQ2UUjjiKs/JjJAtpRv4SZ/ITw7al9QCYcq7vDH6ycnLCU3yhGlJuuSEFH4TjWmVvj
s+jK2tjzGYYNFAIP5hig8eCBGR6yk2zv8dWoYosIgtdVFCjQfjWOW74MSMLqCABGXnWIT/XF9Xil
bxzHAYwVK1eGR7kv5GxKagosycklXaLl1pJVhYe2Q+OuBYvx1CZk6IimyObmhyqP3fhVE4uMuZnk
UqNdtfuuoXufDHOuMfS11NgB82sPIhFPxEkIR4rZg+BMsm8cSi26CAyhCx8g4U3h9QQUcW7mqLvM
aMpNa0d9d3cBVoG7EDic/cR7SXirb9iQuseWcO/osPFGVRHWiQDu5TJ8bs64CdbSUZx0IKZePSka
GbQHDyQ92/cP/c1bb0PFPBWnlNuukyPVpVRx2IqWisj+6VsgZLoUcXSF7Xu3YyemHuy1d7tlhFUa
I0ED2rH+oepyDtrs1YrEbpjD4sOz7dcSA8SiH0LErYpZTVCLkx4cb4hmSFyTFVTW5EVDxfXuBtnj
C5SuvQpM7sz9aAKPIMy55csFiBXbuZu8S9mTWGGl0hokgR0H1fWIKdJ76Ni+G3DQhELaQRe4l9aY
ieVeeSGlTCuZfoLdUekOnPPK4QwTO1VRi0OK8oQeVNTTYpRXoVS922VP75UeWj8rSMEI5bmVDtHH
9SlxZeqSuAFII8ivs4sWoXo6AEYkwXh4AgpTP8Yxf5E6pApFdsL6w1jkMiQ4tpq7+9+C0EdPjSJO
JfLNn0pkLAvDbkH/YfGCCiH5a5aBMZE/lFIbau2AFnajiFy97+oKGRQWf4bDt5QciFWX/3jLxyaB
qKzojDixYC2ZjaZwqTdxoIyXQmzngRI9sA9dTCBV5dkeeUJw+oZ5AkEWAF3M5dSdXlbjgddOjs19
bSu89f5wp2WHeMcYFQ/3nZy5rt1F3RIS0+mPquNNc0o+kfzKEHTHukFJyQ3rdM+wudO/bNFU/cOL
Bq62QkaREFGlEcmWl29hDz+nhF65CWTK3NuKHSn63jjsYt9NMfPnPk2XKel/i29hrJXyr7JRYBsw
rTRHWZfh5i/Qb83ifDLhlWR+dCIN5n45pZXAQ2zJLEZ/heup2JLoLoXrYBBtSWT7uQ8IYNFgWWFT
jqySTUZp+q0WDjitgqNvM6C8bFQ569JWLvHVVZiWKipcGkx+6ZZg9AvNfobKjvat6QVEBtXD9i3K
N0TUsRxqNmfI0GeykcTpcabPmpQEXvlOr0oT3kK8hChc2b52yV3iavA4MXpWrAuJdBfvtqdzJjzD
9Yv9Vj0v3cLrG7EYdYpU2QxHikD4KsDdXZCcUTGoc9g+8YT69UPkQ8BZj0aXfeY0AM6vuHHJCJvz
TGfsh2p849cvka5C2gietj0mjqC5LGHtYJVpf9XhzolF6LtVciyJY+u0nriJhfiXXapIpeXblZyB
QfefDS4g9NXdG+/lUnBHME2WgXUS3KjZxd9z0GX9SBAtKx6d7b/HTLPnCC3NRPmXJM6t55N+GcEH
PW596i2/GO0crKXcn9FW/4JI6J3vjKPGHku3ZfV8sXXhOAEg3CrCIzYZDR3OI3i3ANZFB1bxzfeO
nraBTU66GMmbfs4VFlCurfhCV8KNyO//dGaILoC5K7kR6HtcQIgZaiZs1LARsRHTkqOxcrpt2rVJ
y+B4Sk3M3qTakEcjj3H42ghi/+5QP1Wt+G0AnGK7OJHMSk7ogAsVUMzlz0u9ci4XaQ5dGf+34bIU
ugGLYGcGEeHDlbfWTLzKzyB1OqZ3WXAL7zyvsOpeg8q1iHP8NEQnqAaMRIhD8p1omUHYqTRRU7Od
6N1ZMiJ2KVb3ZZcltHpM61tvODJSTx8VjeW6cFvhkO1NcDzMP4g6SdNVTovHEGi35vmFSauMF0vn
RWF2P64OZvodeGtuNS3JC5X9gw/kEhanAyjGNKVMIptbK9KY4KhAfLik4SVdHg7kS1oclOPcBiVe
KKVQ2fmof/o0YH0+Bvd8G+anWHE9TrM5kkXk9FlIRGkTO0zQKoZ1pd3+RDekVbFkReJWsyhKS0S0
wo1t0ZFk9LgUdZl0HXH0uKrxAlGJqGrLfUq4kcTCKlK4MOVxleKI4B10jwd29FKaYGYupTS2nPtK
VIpW/iVvLjbDw9hs3XUi+/ZCWhTM4k4p78o/ZsFX2iMmbvTeisDrVzUm4yUQ0GYSHT1Ia3sSH0Mb
6uPlTxo0QiZNOBUcMItIzKcO6MAc4wJ0+Jm+wvs5KGulOWO/KuTVYrsGm92Angkc3YM6YPleL1sB
39Fb2SwKC1U3wTESzbjZdSLjWXpbCUlwPAoUjblWwaRsYqnzbbbWSzwEZnP4kwcQZ42tIVtOZBSY
EqEnjs+oBuoAJNapyFxCZx8hBciBHg5fqmg86Gfafnny+J/TZgI2gLh+Nod44ofMKCbAfBRIS27A
euPRbpBfpeIgffUsAV4oIZUWOyaWHfCyAWW3m5kcg5snV75N1qYWr8y9n0veVWHRSopSgjk63611
bMyEuoeJigl/zckjqYFuh0D/p9K6JHsQR9txTNfXtGuMfOosS9q0dbnzb1gLRM/EXTmCbVF3exsf
oxO2LVThEWk+Q02AjpDt8hBMwsc0XwEZtXRyvL2rKcfQ3oOWW3t88VPbGyklMVvm46oCQphTJOIG
zo0NjX1m8Ltn8HCpxGJHSQhIW8fDg6wNRNLb0qnyFppH9w/hRkii1QSy+zsohWiaRmeeFXt8D1px
HMvfB8wAydEzGdkGFmWSjP5ADq9Z4fyEhP5Fhrgw3WxMA6kj09nRBHC9U9BQBw5rW5fLSlfbTqbM
c5W7sYxETtI67IlX42l8yVkU34VhnOMSQAjtqyKcw/sc+Cin+DuXRVzAMKmp/y1pVIXWdS6yIhCU
WHdXO+P3AFMh6ciJAqeENSTy1pqZDR3+8hC1SycH79cb0KPXbf2lRCajI4EgqNAg6dPR2lfBrK9/
9/cddKYQmTyP/ZS8npbbZrZ7y4eQaf4TAt3X5uolWxIiaR8sBtZiwjeyewD6yukbX+YH7A984DxT
KjGMLSlp+rJv0wYYbWUg+Y3jypVxuc+4ljVRUsAna90rroDkybf0/ocOVSRug0nWSRJM+HUtNqDV
1jtwOwPcVBEK5Nk9QF6xi3xLNSXepn8ncnv6x388k9HOWln44Y1h/hsJl5Lr3xgdai/ZCpdRsIVZ
5zVxjUG2E1EIzFsGRPgHVtbU3oJz5ITxERVKERy17ZoRVcUklkmmuXPvbuWpP6WjmMMk2d0u8jbj
qv3NvwWgTUJDdvgetHS1+r2iyYbb0wyX/ZKGMLBOtxZyfNCVS3JiufgCEttmyht8MZ0KJjGoOydE
hMTmi0Iwo5NE4g9ZrasC0Jh65DgXW8babxFXIeBA2sB00vTrebjL88HODvjq1qFQvEyAso4oiZKX
zCbjSd45VxzyVtShAPeUmm9MrQnA1yKyqYYxiCcb68KrqZONzTIyaMTZREzBFgIDIT/z4RoM01lg
OXA8v8Gi5x0EivRCFZPXap0eZj6lS8e0jtlRCs09Fxu6E8Pc0kI8bFWC60lr3mvqScqaUr65elvh
wbRnmg6lK2xP6EJ+AZ7EkplD5nrw04ZLavfprhZkPrDc/+P2bB/pePz4GAxUdUsdwz09h/HyNnT/
90iKUTYeSgA0ECy3kimcw66u2h7WZULIYVaReF0sqUHdy9FRcsnqPaMVqdjVjNHcIyk2lS1YgClA
whM7vkECimVqMjUXzx6lujDOGpiGOgzLNQCQFpSbzudrdAuk1kMQl84+UPbWLSBClRD9thRwZMdp
dsqQURvwLTbOgI4aaJBYMiyYkz2LS393q+fjRENBkRjlcAA6o9GbVbenOVlKucizqwlTH4A2H5bI
+n0RQxlgjgi78PqJmiRaVUvAbzGw1fK2sLssC5neqaEYecAjx2s0QhkwxDVGQF1Uto+IFn5nBiGa
7vdARqLFg4cDVbxNe9y2ZGMIcBEWNIb/M4hnQcu3/zDnX1GNFVDHkY8CnOI9G/vWOfB1ZGjPP0cK
elG1KUxwgkj/oC/V3orboPD4RjtDLIALil3UK2jM5tCFNYsDwl8pa5ARAQ93BLXQIUTNUuL+BirW
FjVv+qM8JN6128y6StrIQVHwzuXf+CKpkyl9w498piV962JVO3yVV47dw74DMLnsDnUo8kYRRN1Y
S6icesPQ9Ge9qkTdpAX953mLMvo7rh3rALd3X3qBKZprOZQRgOsktdZ2WC883G2jLrdV0YQ8FHTj
P7ne8xj5CUyRcNhN8Lbg/Iddht9UQf6OTKBS9hrGtHc+6f/1nOL3DttxU0RWapFyWrYoYqQCSUto
T0mVlyn9gdAjr2E7tRNBCMve5fqVGuPODjUcXkmZt3u14+bdXnst1vqPR7ZdCFAmeBpekfT8HDBq
dOJx0BXJjZVYNmBKDAxYdNaWxSU0xgO85DvzJ4B1lJqES6/5J5OA9Nlww9vetm9e85tssUg8YsMh
khCTWart4UxbEjS2SSVQwNask+frn4z+m0fwQ+9RMsj3pu4w2JXAWs9m0QyKpp0ImiMtzdghFdQ0
NdXxWCh5CJzjX1much/0g0k4PrlBDx2IQTlPVjRM7QiHXrB+8s7TpxNQ48liDP9IbJlSeofuJ7XA
a0Tv9MGNdet3kf5j+DB2TGhnFM8Kd53xvkC1xgpbovSVH/8bWLrokUsmVv/Hku1PAIHqigK1LOgG
owk30yQ3ZaK28jJ7EYORW1P75y5HtGFf4FZE7koceU4vC/yOQYeZ7ofJAIuhFKw1jD80PV21XE3a
YIN/HWwRHrT3Gxn1TeBJLT59PXl75HcSQnG7m64hMAN/CV0g/NZdiAcv7/N2QKbnws+Or2x93yK2
oTR5ZJbARFSHGYbwcbBFmz3HY4MZMxgx598nnz2bEUnO1J3a41lVyAkLy0Le2PhGxdku26T0lR/Y
X5CKQ8TX3xPUQHL+7Et8WP6kN+YTHp8EHV2TfK/2nIL9nPTK3SWU8sVzSsCHrXWFo84TMAvpr6Lz
68kT3z4KqkHNAG1S614XzUe9Pf+GmOgofwUw4xcFIwjQaKjhQ8uyp8/zkI1WyJj4xRLxp43bnnl+
9Mx22gwl0mkWhPkJfCzC3cwX3TVczfk1moY/6fLnMydTpXd+IPwGwfdLgkX/98JOTpMZAhrUM7sN
pRHe0ZpXrfvvX3r/DwmaxRDne+v8x/Kxquo1sgJ9DrtoVVn7eSHyMXSkHzngzZ2K5TYSRaygTBNv
Vio9ftn4C5Dwo36Apdn7qtJQVFWOzRaACC3MwzGSThDxCQhQ6qvFjaXZ+oZPcB9vTbZ3UAFUKR9B
zvWp5mUZGZ34PG23vMCpO0JLx7/8be5NzoMDHM5u8HaA4QqTCqXg8q/bb932EKl8eUB5vstHYZaT
1L/ViYZV7jea6xUrshZdxztLaJsPfT+ke+j4S6AWdf/99zZMukdoJOuJC+i//Mf9nJVDPhXUsXkc
TjDUzppitQ66Ovu7SoGTIQARLyYAD8IAXcDQidt73vaXwR9xsrnEuDtqpAXnxL2KU9Ssq4/FiMfW
2w0mE1Ssq0SHT2fWleczwcRYOguMCRLqltfcLWBeeNs0RjCJ6UmRRPFkdvPCuxfINyEnGD/4jCuz
1NmLb1PnSL6tgPACYblSA49eiBsFDT63UQ2fTSs4luKxv73KieU+BbYnUDUYCoFyTK8obw2pL6Kn
Q/7k9BimJbdTQJe0s1/4gHkvAKOtwG/lyOKukm1+MlW2eJw5etWZoSrruSTX840XwZtbcjGEhieX
1lu4TN88uUonTCJJ6qMcC0hCdKS1lEZYelg4Do99WrLpG0lXeoi15pkEIs93oL9CEUwzRWFFBoth
VTye6flT2visY7vnJ7qWSfw2PXTXA9Zju1wkOZWuB7YSNgiKXlOZsYVO/hrOuUroSzkk576p1LLv
+FdbUaMAlTg5n+RMLS2Pp58WWxAbVSg0wjk2+cg4+LrJkrz/cGJL7dgHDCp6xPKIbmUAg3QH1P5H
UfXznpanhopavQEI0FfkUbqDtknatXkhbOO4pc+I5JvE0tOcupXry3gPA8Ewu4YbBbVZ0vf7E7e+
KUEQOQHpdeEnAFXEl1EBgBlZDtmjE2Q4zoJ43YkwjaXuox6vdOuto9fUw2jKqfGmZgdtIrVb3R0W
z4EU2HtNr6rPOjNKDg2e/OwZM8/yMK55Rfxbi7bRAx4OJwcAnb+y1aU+MTSPWEvw/JlNHjhPI5CH
2slKrU62k9n6cmjM8PIS1El5EUjwhnmcGvwLTMP2Rv9xjTB2OMNIYHTSxIv9MpSyUZJ3CWt8Wh3+
BreLvTlDOv+m3JyplIvIyiYuqxZVpviYSDfXzA6JPrUylqFq46pLESIuSJaPnWtaKV2XVkcv7ffo
UNGeakTk/Wn84UJgclr3QvN6ttm2/ZXhecD2lQxE0ZdHLl2xTZfkWrM2JFZRL/VcYMmR+vyt+d1p
TNgiDWpdpDT2SjH0pE/M3NGTmEJb7mhU5raTKxvOdHgYxb5qvtErAzxdN0PyrjY2OYnbWeG2Cybb
aH8IWWHG4A6lpmqWI4v1QLYfbLCJS2OdDZKy6SR0wlPoebhDJ+7ZSqA+l1a8A9TQ6kaqghM8pz+L
t6JkJ/gYj8BknE4a5Rmu1A97NgoSYvSKsK6/HQlAKfXccSbmi0bErqWAotnhp9Wsm5+t7JVEcKeW
wNd0iJIFMCz1xVer0QL5lI8+rMOu6fhlo7wE1Y+3vWqkzu3ITs8WFXMgtuU48Obhj6084V+Jw+SA
agQRiEuob3nGHVefB3i6+QDurI+zV45y+SugDrbUJgGpgQrXKjDYEyPEsTfT87szLLbIKW0hiSOP
UzVeX1OoOcV8EgW+7NVwmcJ2903SjL3Paw1GC6IojLHvTzRWfRi+0lDy5iA/4Pz8DpX5MsPFnBVG
+XKTU4dnKnFkDe9osjRi44sO+FvEeX/+fnBpW/098B5yuWTB+RZxNE4uHp3PpqWP3jDoVvccbPPG
iH9dNwTyODhIU4T03z8FNJRTSATe0j9zH2P42qUPIyaquKqvjA/RA/efg8hsA5XlJvx6CJ2f3zKf
nxAZlglvLhfEuMch5WuU2XIut0O9XZyYpYMw7rLqOW+tv6eRT4bm2ukVw6kXd6vjrsq868n5Ld6e
UwyyBV6UV7SDUzJfNCWZ5DcymDFlYu0EEo6uGYC9kVg5yDFHLiaIBoJ7Dh2ML1VBdWOnyXlTBgiA
Pk+iooQ2Th+9U0oZg+gv/rHO9zU7aY6CAJfpdDnHjBNmE67ZTfmiof0817O7l1v+XbGi91YpvUvj
5i5727lGWvT7p9bbMvEoXCJ49OQJTf+EbZWZ8F42NEJv1ctiRfTPMd6YF6rxvqzQV4rVbathCRY/
22CHfUI6OWB85VrWx2OiYAUUEr3kliJGsFXaxYqiod0V57t91XWF+Jz+5XmQswRrKM7CvqtTDGPe
4n6oOB8OV/Mgj58/m2DfOYOqV6xmR4VDg321Jh5HOPnf8Hgp5KJz7o/pqn+J80uHdwuJlaWHtwmi
qLfEUF/BYOcWi+udrQlrM0MPj0VudOKj031dAhh2JNY0CxEH88UwL3ECEyUxmRCKsNsTASlTPon6
I5DVl7QUJRlK0CfuaZL8fgoufOPYWUbFzJXTQ44FPQf39I1JvJElPdLAAJaR1bCIQYvC1sVjW9d2
IskEXhjEdHGNJAzkLyoZWm6UN0qH6lUOdygAzhFMoZqpdPeuhe4tAJz/9Z4WdGTsGOoKFW1xQtCV
1+q5R91sT2Vp3oklO7K0TFvTJgdSlLbqciHurxw+tkaCaF7qM9Dw0EykYlGNHzmB4um3ACh/bcox
EVJytY3avUznbJgXue1NuhhWBCQsQF0N2bSe9SakiQ1KMacpk9BF5cPCQ+3r2VRm3OlP7+wuyNEk
LhteIIoVbXJXTNAisB+mpSq3A8sT83Cdphc3tO2bwbma4pa/5WSR7rZphBXwOxjsvpjYP5+t1F66
DdKEcLeimN7LtmAHkegInXdpyKKm9Q+vTxG1FlRw012MxjIRyeJProK5AERKZxUOSmtebF1kH2mu
5+H5epQn+xptiTB3LNnvAlvuTqJxgq59Nh+U3c5xbIjhWSFAb7c2mN5ngOmDtMU41Z2aAQyIX8Am
dN9AeHfneDJw6pCeJ6yK7XY9N3cGRufSHLWK14j8Oe68Dt7Xg5r3RfxdYc6KuvcR2Wm0z3nrKO82
2YYxKaWPBxoy/7xuZGAAtE21ocaymOJ90EaP1scVcS/kdP3xqIomSuNQgMG2h0ZAN06Exk5xGy0j
4HNPBUGJvChujLw+XX6s3fh+WQ/u4kMTvSEJ1QoLmFFjGaOZ7WocdxCOB4J8TgCVnUNZnJQlUiU/
k/0AVNKTvStZWk3Et9gUyylZd5CJVddMOhMivuw/jrwHUGQrov/H1hkYdVqFBcaAxvhK92YN1HBp
Pnomj0fz5OY1C98eUqJt89db1EY0obyrnW/cpRQnhwHBSyoizD99XLSptA+Tb70LqT8pjpLUAdPT
Lfhs+BKXxKQFPsqYy6gjuxHNkXSJZMP28vARea7BxtqjtTyH3fuumIRzL2P2NSs8hwqsawNh3PGV
mVMQnF2RWYUBpXJswzEyfKbcezEXh3rttM/WusdUq5bJISzyJgJdJDgbdLrvdLy5WPWK64aWo8Cj
xU73/LlCJYanE6SwJrQXyxR+ENdlDvtq6mVnjQZzez1Bj/c2lcLa237zpCtFA9cD62dHBraORANo
cUqqtxFVQ093CLj0hOv3Ru/GL008FXx3N6jXDaY3sINOvw0JMObCNFt6/T5D+QSSI34EQNltmFBZ
ZfM6V1FofEuURqsq9K2kRs4EzNfcuJgfb5cLEZu8GfywLVREY2LQel5xPqlrMvjjPlPXM7MR0Ugy
Ajx77PyUKHSnZdL5Fme2nG1NPapJzoQF8g4cPq723yoEULNHWYIgB3Y0h5hO2jzaJXt2qmcpSnKh
acTHYgBrN+Q/gwkVhePBq8+mxzK4/Kk0AmUC6Dm/O4ZR1MtBZx5oHKs+vaiYgiCT11/WfXes+J37
djCwVvP8oyYssAgqk7ysMmlvy6IFtr1W7IV6RmH+uqG2MaNPRv2AgujWY+XEbMK/WHZKI/3yHrxe
07VAxTnGYB3hrzCsf/CPBSqxGJTFOaxs+q5rXpO6BrrSS4AmclWP26H0UedXvAwbLaJhkL+M9OZ+
T6EGWA7/svNn5/WEk6CDOby2j9ftKHaNiRWyAEs/vaIP+79UmL+en2T6qNK0KMYtEw0fhA7PrEV+
WI/heF7apx/P3e7F8E83S019B1kSne0y0q8ni9eq2b6XajdFgp75ZMNsLvXHRx8g9xbywLGuHk8R
akfhPdK5JNvUUGJ/GM71R38wHFxgZZZfgJv/epGm9yzT0G5n5n1Yr084alpiGw416siwOeqVLpjp
gSuErrNCPaQdr0c2wnpe2ybPXjY3+S04x/vPpFjBBqnsoLu7jxzatgPLykCSOIvcQVhjZExaFIp1
o9kNtpHRsRwTjkJn2vXgpYIkz+WOnLQWfL5LfJn+WAFXz2HbX88bSLV9PE+BJlAxD0MXiOGVy4Dt
CbqxRvAnnYHrn7PrxUZpz+89vo6qaq2OiXhy802g1QhXxtIen64R5p0l62kAhYSMvXmQp5hJzrdD
D7IMSRxMbENb6VErA+4NzI9H5jZlhJaf3UFJVUxBAlPqfFpihGuxgvLnG2zCC+2SEozqPkMiLwNA
SsmILiuvzKCY6XxslCbzeu5E/9zBCzpHRpa6uV2/HESBkrkqzThZ+bkf+UtuKQloKI9uY7ZPNwIO
PdkRGAAgKrefdsQShzjQpnpK2V5oMvsdBiuKbFzL3TlvG4lCy8adUP0/5G6qd2WfjYJSY+6+hisJ
BY9/ZcVfU5/uZB/4eXzc5AKzul4+Y5uszywrz4umZq353c0kP15hO5FEZ3EFAAw390HYTta2+cHt
tG5XlEcsTpLwa9OIn233xa0irG03ShRaluXlSA30VGHjbw72rAAuZDG0PXSuF7y6HdKVK2c2V8rI
j3R6gX3deHqiYjRTSnszlzzMB1cd4idTaooWHKRHHbiFdeXcBgKmXUiT13raNTlX5GA7VWm8BYe0
2JApH1lxvKbfaM/Tf7SmgSblTw7paDGSr+jrsp5UndWpb7S5doZhaGljuP6heALNLvo9bwlsVPzj
g7aTeAwHO9Nw4eyxZ1XKHskw42Lo7Zk32HKYhYtlvjpajzDGcGQii33DbJtnfUTCV7+GLUWzNOOo
EQYpj+0JzhiPZ1aSXTN5t/ebzjvKq6GZjilUWoMFvOqdOCosSMGgRB0SoOGlOQQJ79gl4r2c51zG
wXTnvidEX7ywmFjHIE1sWYK42aatwW70erXyUORaTeJ/mm/0QUoMkflAL6LCiDYaSdAiJZ6s82P+
lqb3TIjzJcGJRe8ywuw/031jyRp2rnHa7BpRUD8EWns2TAOJVS2ptdJds+4iy1VMFgcHTM+5MbnS
ewj7+IDXUzHYAtwijF0S1AjQrp0osykuG/1dLQ/u69qxiGp3j6FBX/QhVn4DCMQBxIHKFqNtfJEH
R5ANXQcR1H+m2C1nr7QhYN17yySra8nzLaENXJdMU+Dl/dLTTpoSEmiX/QUYcVETX9lqm96MlOfo
7QPUBIA5LCD/FKy0Y6dYDDaT1o+zWbsbuME0Z8t30XFYNZS61o8gKOwnwjP1fG2NOOqrRBMmgp4T
UFOQWJs+ApoMZRwEIg9bNq+poxNH/qJzYtQnuCcDDFY3Ou66zFVEqzbas3K55bOLmyIGqoGQ+XNi
q5bamNVWY38bhhkNufMriFZTj0+VnhpP0Emi4EcpdMQcLO45APXCgfQ3WtLxE/bLtqguCfr+PRWW
UGIjjwqvJw69u6YLqqrc1qh1lPiPbvB+3lf2Pyr2yFLSBrj/ptfm/SIdFcaWSka+XhLPpr/bOmbR
zCRTEpMfNTDUKc7wHw9CW0H1fCBlW2HXhprJsYmGWE/hC6Wf2zOMEq+ja2u5B87fzWrPdo+Yybeo
UfXahdBOyScDr+ZpMXB3u7a05dz621WF9lzuowWEpLt/MfO2YLIqYD4KqZVUClGMXMqPCBSW0Yl5
wqLH48nYRlA0ZD369Y6M0YdyknBqAiLWxdB83d7cfDTmQEvJ0CuF8QzelvSae4Ljq/9OFBbAEQhl
fkg0kHQlE1G4vULPjhSXkJw+4PRXC0XqobH8/1i3YUChgE04mIlBQaYmuze0mTTpHXi3zP/xBkz+
kXY8jNEE99vdYrXnjr2Ag9pBWXfy4pYq8blwY1kdz9u4HaQMyxPlU2HjPTRIJ3kOR0MzaKXCZrtG
xY7AIRcR7wT4ORuOlnLxvZuahSorzOXC4ctxr30m/QA6O+jbuXNq8AQ4aMRDlQ/7eyNTXSwE7k8W
5edllIoh6KiI6NpKAjNrejoJhxfchXk3/tjJDtuQZ2vpOmQ/8C0rUVheCDE4W2Tl4WYjObVzAf1h
m2YEJ6XxXbWKHdWuspIOyZLmNNyRbb59LxtFCWL1O25Tk/76GJs7OtM/d5UElZulfy5ggMhN2f/d
21t/DDEFWwUY6G5288flks1cpjdg4RYhodOzEs7F8igngkpV41HMcCwBIcRKm7Dj8H4B2mTYUu/W
8+LgQQ6DDc5c3sBQyhmXS+7GhFSyLjXoI7Qcrxxxvmvh9lc6VDXuwmuS1A0JQgTvyufrjRGFZ4Hq
DDhrNmMdBlgkjzdxnCdhTeWI6fD+K85616BYqPxjEHeB+999F/STUM9fS4IqKlhUBPzOJjPjXcdx
XDft4lK5Tg5MpVP6vOpUcNIKewCG3ay+HFvW1Wd1FtPiOPqqKvGQIgxgM+9IKO2mlBFSWpnebEgP
+BxiqaLrkOiA+iUdeif0epebRTfgTaNxip93vaEGptHl/Bhs2qfpwCg4ZMd0Wod5olW9RsRVm78Q
Qu3eSK6RAkm5Hr7s7ADDzKQzbnUKLBIyXfC11Pk/f+ckwk6dDd2ibMk5+UBbKwEc5XuJo4kCNiVn
o7DtxUJjgmM+Ash0m2tT0FSsuVGVwfLMkr5bNC/MbmbBSM+iLxYCJWTe0j2AoBE0pPcr8RnJC9Mp
N+R5LntCcmxOW2aowdC1MdaBoPjW1B2c7wJW3HLDVh5ssaoN6HknZRZ8MULTcUKSKNruWCm2lRwY
lKC2FLGFNqBleQkjJgkgBs5/987F20p/BorRjvY/w8GlxQuxi9ci+czExdb4+8H9c4QH+6wJfN7X
LnnElSpDrHoiad/f1mmtInj7p0oOoG0BL4/t1ZSIaocaKqDT2LMGQgJg4cvurh2ZDC5krSmNJ+xx
hboHqmp+xh0G2DHYjezWBG9MF3SAUaIsZggrbzYDG10czym1HYmKZl+9Y76nP5O95karM9VrWd4L
YqeaB/aJypfrKhVWH03nIAo8Tt7GeNU7fYReilnTt0zbh1gxd/en17ZeCaHtrsx/xIaLdW5zdu1N
0xhE004Z/9SBNgE+c7JHONu7uIlr+jxCY2v8YMGIaAnAWL043Zpxuw94IPkTcOaMe/WnmUEVAR2g
CSe75l+Rr4OBFwiB0/lT6sPpgRpsm9u6mhd53qKg1YTFhKArGxbAjEMEohQrS3Q7MxskeT7KkC59
mPq5UfO6O3XMl/61s9EJLh+sxsC8DN/KKZhE2sVupYsP7NUsE3SM0d91BZH6jtOBmBq4K63tp6eX
Kvu0pqcrKtMAHKL5F9VDmG+4CHlCWpI/EULvFr+S63F8XEI3RJ14n87eVaDoy6+H5TVCu1oH8o5J
XxYXOFKhoZxUtICKMcn8hqvvKmUlp/SxtjNQ84RCw1Ndqao42sioHsh8KrK0vqQLA3zEOQTYpRzh
X3FS+RtMHUUgauAkoojd+pd3s5fcKn5zOJ910lL4T9GdqitcFH7s7XH8HJRpEsTPDb0gkPnjeVUp
9DnvRCQ7pxmuRTJbCxpmezEHNpASVVggKhdhGYWOCdDKcy0EhoM3FLWAc5goqiGc+1lA5TgMS8vX
RuZjmOZzaXzmpKo0HC1q1AGQz0tvddRsTNZsdsaZB+WvoE37+HH8udaRuNQh3qLCwC9pu5ljdwjY
887XkEvmwm1BZgK384q5o9YxAAVRKvdiVyhjqyQf+YKEnkmK0wOV+2tRIyi0tmu/bDVjx0afYlPA
giDx3I1AuDGbbc20auX0ySJP6B6qIWzDGOy/T09t5WHTA8Vqoze3pYmZYV4zXS2Nd169iQ32bLE5
iW3FVJLzlKYG0w+JCqsEKwtZrA7jZl7iKLhrVbyV5It0iyV07n6WPnIDolkL9hqWHQfECp7AzEK5
sVCkgtrlTMZTxBXbyXx+ahZ7NMrD0vEOcgGWuDpneoAtapBeFVxjWutxZNv8AGS7YjOm3uaUuZdV
3FsXAbP/4CM3yOVA5F7MpB/2/uBswWJFlPgoDwv2tdm36iiSUo70xwcEXVAN6la2l4szp5Jnm5xB
tdNSV3RJw61vmlgppVaCTHuE+mVSpdJ3DP+mqtK6puttT+G2V8MeB73VZtLXGrj17gngQ0b1DfsD
ZQo4s64Vb0RVFxIIcDsjhyREk9ZKCI4hIS+mIUdOYZqQlmE8PVWmVnMGtnJFWj+SAiemZoHdH7QY
rY8iyth0MX6UP3Cp92bOCm94b2vilrYNaet5nd9ChBcdwaYbXCP5NlMVmWFjR1iFrWRMfRGxoBNj
G5rKXPMayL3PMOk9GW751jgjA3kiWBoOZTV4USDzufTeHPoyQEYdpvufDO5Wh/iAollV7SnlBrZ6
+knIujJM0fU5wy/6N8I+3oWmT5h9S5/0c8Pm5Y6oO2WO0Klo/mb7b6F3bcnSH9PUReAfWk5rRXtb
hYuc+UWHa9o9vhN8gE5o3oqM7JxbvefAxICKXFFBpV83+6+2v30nZmmQdlechBClwCyJ8NCIpEK0
HmtsouupoxIiMPbyEox3g3mFsvBaq/PjlP19yq7Y877ccqiXK33SgPA5QLqKzVbJzjQLBi4QvUT2
yx9laaWF/ZzSsGvOXfKnahFJhr0Nc7WaKREPSCs7PrrRRfXfO/CPJbBOjYq8n8E7cdruHVG9Xm8s
LH+qrYCau5U7B7u7koFVcUGhSewozvSGSvHMy7Ki50IQeyIVRHf7sh1rht0tcQFoqT037W365p53
cumRb4mtZjRIvlIZp2E0Pi+N7lMblodHPOl72PrQJJoIYd8AoWgi8V3pPIonlefQHH55cTi6WT9z
u4fneTquNDBPXbeaAdz38C0uLlpzDNn3txNfFVWGLyBz1ZTjcNB3DYdv4GsAEtPt53ImrdA4gt42
13qy8rZFM+gIbHcOqBmJxTXU99AvcoDsYlyu2xttbzFY+pxEViWMM8FHDHr/3RqsOYRhRC77MFn1
Lj6HAudiKcC43yQUjORtyYdNn67T8EiSHLi6kKFmwHHdcclR91tvHYoSd9YJocmNSaeYWx8i94lc
hQFDObWiP5dS+5HT+OEzjRafiAK3QOiLEK99rb397FP+Bh/W+nTlSi7jZ/Caz2g5Duaw+KN6dJqJ
VZ1AGTXxyk9M7qs9sSS0dNnzssF554ubN38cR9I5bChrinB+Eux94oo32CHHil5U/f0IZZoNK05d
VSv4IpeHBCz3P6vziN/Eqw/RGMo+My0XOs9xuk4yLkmIW7uWXo9x9rnvCIFPev3wy+TShvGUjN4z
aB8ysOx0PW0/1TVfgnosmyo+ZH2v16deK/i5OW72qfmYVpJ2lrzNudTwpeLKYJZ1gyOd12ofPDKq
ljIqcblw7bIkEd6GIkf4Yv93fF5oHqhVSbxkgLVEaNQao73eS/kw/OII4ToNs0U64PkdHvv9jPex
4cCkbIWoPB5fOfSh3dj2OdqESdfkA6DsHnMrQgTw4dzVuSNp6k7ZRT5nteHH+RtSgvWbe4UDI9Sl
4vsjBUyj3m2l5PyuwvLm/HzUwSkuFQrQQBy57BMOV13scl+WYLMKLm2JZcO2r4vm6ccMKoBUmhoN
CYBy+bLjMWyfxYzKieBaBlgzV8q+caVG34rqHmZXCbWy6grAgzxRXud4cPEgOvMwxLHJa4lIub+L
wapNqmYAcikL1VDkzgwkWuJujgi8dSAacuH1Vz3oHSFn0Ws0mjdT5I2KP21WSgACcBlwycKjC8iH
fubmzXwr67c/Fjp6LoZdKqmj1nLJVxy+EcJ6lD3F/mZ/ttjVxC5Q7EcCZBHzE0o4qAq0LK7s+i9H
/QMOCqdN+6hEi2RsCnPY7MAK3ovIGlZMCizcvbYyI+60XeRLOm6wSN2r82AFXabhZaCWPs3aACuu
KcW1XqKruoUE+4bmgmlEkP5AWHywFph088OHlToJ5MbbzfNjXuEqoXbv+aGySUNXjKzzhJmRgiGB
n5Rlp1zjGkeGz1W6vbYwtMk0Gr0OFltV97VB4f5/c5dkjS+gWHt7zUFVr5RZKXoR8e0MtSX5M6Ie
6YYCIZe+jA3wDqsQGSdd5rYiynDXgg2XNSKNHUi2SmbLwucEYKqvh/H+7K8wFLjbWp/+YJH5Bj85
G06OHIXi4V+hGFg1NaPvFZGH2zUSUHWbiIpQDvxsU6g4aLANEgmyqhMuM1KnPzAvW1KDjiqXMUL/
49bTD6FBLQ4AFA57RIZKS4xBZJdvfeNMCuI8fnhQqmHA0BcjuU1dCF9qkZmkJw6g8DHzqClE3AUn
wQ+BnDFkpu6FsOYAx459GRpC5M0mvmIB0vuRkpiXCL/Jr4lpRINEiVYVckettMjAeZjZlTbPo2kI
5aMYh2N8TUvRHVzU2mT7IrBjg+cz7HylF6gDziW1n5Xb4s9yT2e+g5tULMTZUCdpGwL1zAL3LNkF
QsQTpY9L5vy1qmI2Y4zxFnQX9pD8mGuHnnrQ/XV/K07Eqr/Qnso7XHbf1y2/2/NxDg4hn41RYMxm
6tPkErm4ek6oPhpvOes0TzpYyLlgTgAmBWT/c7oEsk8/02Cq7pYI7UfT60RWJYzkrubehTp2903l
gpOdCcD79CxWgxehi1xFXPR/L5LhM1rGwo2WR8o9/QL9yEktyDB2JJIghm9Ye/0xSjRbQfZDl0G/
PtOWIGmwf5Vba/LRmx0p32bhOOJijDlYa/f9wCCuoKRg5q5b5TfWPQn3/AhG0VXso9QGrOU/4i8/
LXDW7wbZMdnuCDm3lyeC+zjxR/qzM42PJ502kMiCsSImtck+zjetUOknFNkf1VNDWnYoFfberlC2
WQyG2jFfs8FoUX7UpCU5m6TZ4Iljdm407jdevqv4eNwVW8Ti/CtZgllnZGZ1HYCTyUnyNrDoevKO
O84sJYKOO2HAEOoJdVpQXpwAzHisQBDG4B0RtIXiLBP4ztWFRElMLn+JC9gvHpIqGxdd9/mc4rF7
k4KOJrhHlWZUVaDU1E3HrgtH7JkT2B74zRvdAuuXLgyeu8OPFPZPCSP1A9luD1r77/vfZnk7WC/k
g3OPc9P1g2F9nA15g8u76JYS1A5lO7yawyUli53kvoQEonPEUGPR44Wrdj4n+R71FTQ8CFDy8Ogt
CmvD0L4lodxfm7jVDr46lVazCtna8519mYlF9e1sYW1d6IBgocxgXA796X+F+bUu4Cx7jlQRVLI9
CF4W4DfhsimXaQHy6JbVCtSyqVpbrCo6Xc8hb1ixcbJagVLmCsru+SoyZfBqPeGFbIiSXYeTYQPc
dkM7iKoD0X+KdoqYt5RdqHb8910oBLxKWbmCyJhTEjaiwHaLgPjXBER04CqNwSAPL1om6vMWghpG
p88iLkIlZt5BKOhWttdtrcFQ1B6tqYz4kKhx8qSfd0hEYMoSyRxjMXjxUurFddkeZ5vlRSdCQZy6
3JV8sHXHn0GJcaxsdpRfEeaqI+0ndV2i0KfSy794hHXICOifFTXTz4kKsEV3uSxvv/O+1htIpzEW
4yrsFWkfC7O2CdXqVkBFO+MVeKeUFYouZHmXi1mHQUgz13sR1dMMDP5xK0rGeoOujGF6hWhG50Ql
3Y9b2Fe9L2MnskbmXFh0379yKAKI2Ew3M3XoOCsC5pPfc0PzGZKuQG5GKktMzxY1X+KZL7juq1cn
WaNw1fOIXBL7kBy8zT1r6DOKPemcoNZYCWGQFbjPI2LlsMxKd2UJsQgsuKKyw4LIhquNga+BwmgN
pj+RPovqM2SNVDb/mHM8YmRb+AkU6FfR2rtkfXp1/qZGGeKawYuf43MTE9qiSgnsOCAbQdvHg3q2
UDKixmEoecqDuo1P7GJzsWlNXdZjSr5RycN7FSScqL7+y/PbqWPTYNdusRS5X/6bkJ6l4ygQ1Xe5
HvzSmHdP0D5bs2oubmF8Hpn4f0V2e71mTWF+gS+qTVAUO2Jdkd1CKa8KaPV2ZnC5R479nXZ/yltN
+rV7NGq8x8dixTMDrHiAckdJgY00vXulPM5XUdehIMn0tkuGTDzBoqyCukknESm6LYRBwjiyoKhC
0T/brmtDX+LHOkQN+B1btzc8g+Qzb2/LMx7HmT/qr8pSEpDMdzc7T+dqF+zInt0ktJhidGSSC9yF
5f5DHdIiKn5uYPs0rUuyD8jDk14NVb80pxp5ZLMqyBPEbpoXrdQGrpsBVaDe9MMvcp9MfSKaolDP
LGIThsjydVXu4Of+JApRfsT4afr+jxgShFBmVWu14T1U8h0SLf6bKBq0DpT7BSz8cbG2NpVC9O1I
uVvPMLbji4VGsA5QVLBb3Km5bZJp6OEtpMyBoTQd9qo2Gh2uNGK1Hr2WzWaha8CszdKnSvtVsrIQ
QSDZ0i4vWMJPdpb3pmo6q7CCRNF7fjkGg93GnJummrn+7QyLewQ/P62XaiiJfaacumceETsM5SKF
iIaB7HlapXZMeITnWp38zu6hl04W0F5C+w5Y9u+28ek5zb1YeQfkKCqGI1S8K39ldXDuU3rqUVZW
uoySPvM7AoRYtLmwKoRQt5PlhDv28+0bXjuaIvvsa09j41/uRHNN3zioAQKz/IsNn/2xlETx2qj4
UqslNmg9FMWzOzMGUbS3DALMUv74xTdmXb6i+bfVJeI+5EK2/2FCf07wgMfJ5y3dvTzHDoBwiAwN
MjbyRRl0ksDvsLAZiNp2WncBX6fpT0DmxiHvyXr0o/WeDL3Zbaq4gcSE4ULzJNZzzGqvdvl77Cb7
mTCHFeqqcEONLFJ4hNCcoxMzrbyjBL6CQHz42axhF+7WW12ti0PQSjE4rgh3R6pUi6L+K+yItvfk
3j2k96kT508S2h0rPL1dF0cd0tQRgbuo1vzJDcfd4pmKzVcEsRdd9gcjmlhUZxuWwHSooForIrpV
93/pPxS4PNpwgSaDHbuxMVcCXJyz4lrRGWNACVigKMHgO0QMXZX/UUNbWBwvVhBLKmrtFCTEU6Iz
M0hd7y1INCz3YKdgL0CKXEW8W+qRfUpwjfglWbdiSVDnBup9UQh7seGoK+YSWvc661mTN81WLogp
jh90guGybzO6iIbd9osHMVgwBx645XiMvl+NSLNT8jZMZHvO0nDCCG1TRpfywqDH6nK578FGJwkb
ZzmU70X7i6Rrrtle7kkxGmW5AeWsc1Ru7kjaKrpsCgte6uK9vjSALXLUR2xVEegdAKIaFH0Kl92H
PZ8sPM2KjRCHV4sIxRRWq04mpLUfbXIsqeZatR3sEsYunphgIa71lkX7/7xehbx6/JKUlL50YQas
dvo1sJFtm8XWBQYkPd+hVXz6aAkJFPBMctNlijiFiQe4Td6WJAfG/Wbvz7gIuzNDN3J/DOc6S7aj
kaIBW7VGzvyVT0qqBbvjCYBSYmDdpOoz2qdfJxUu1kC2JqSwQ7HQ/4eI+bvtSe9VdqSqhtko5fiR
ensRzTv6Z0dfAcOQKIpuC9gfLZFQbAy9rAqt5y9nMGgQolCBhGxZbMS7tiZzZfZ9ny13XXi8YylS
A5qrx+T1lcNoB9ch7oEeGEAN+5Z7TU2Mv4ZN0peSETeBOBXHDPRh8hJEAyRUHiXnDi82X/pG+JMx
yuwHhyNgTmwgLbi7TUHWGKk7/WSrCkvGdL/kWPw7OMEKDkawENLb5r5vbhwTBI/FofTy57MVcK03
s57CfiBQASdvWuWNNrcuyxq44vwtk1tDwPFDy0E54bvqfu27nF3NbKwH0gHc6XSvytP+TPLgYVT7
q3YHlBWnrxVBAIxkE1J2uoshOiGVT8vfXJhhNNXwHhlj/pV9fCLltexyByhpVo8mvVsnMrnYl7W3
oddKsV6T+FOQQpH1KXbw+t1mvxn/4XyRqk4T1YApgchxv0LEr32kVt82Lv31Qdjy38N6NJdH6OyR
L8pWUWU2FGeGk7/QIZpn4o3hpxA0Uw4eCjJKbuRxrBwdYoeTNs+3tpsQncU0i6WqDfgkj7+1zjnH
Xiu1WMM1vHqmPBQbm/W58yUhPPNnkW36wpelY24A1sDSd8gQRHNOIvGrJ1YuqqxX9sIuouW88cmU
i2JF6gf44BmR0thGDpDjDKnJlec/Y/LGvqMSEYy399iavh++V5Rt4LoG9gujv7bFD+Wz5qg8ZzF0
paZVjDPe8ap2V78v9QhjOp3bNnhReBilG/HjAozEEnwPjfONU/VLNDqzcs20nqzaPjGAxqgkSnwv
I/Vkor3V/RO0jE99/dk5fdOVgWpPOL5zYISrmY8NPygA63tfpQ4VRwqal8rXHrLUjtGjM+abrfyg
wner932GpOKv//izyBKwH95xJCxZ5wrSvgNOVLJW/G2nrVlMXVdU3evCIqpxkpGKsE4UIVQgWeIG
v62fY5/pC5Hjwg1meifiJb68RIrvJq0L+wDycKF/r5G/vhR1t7WaczMkWXJPsRAKWaDJzdTImoC7
M2D76Xy0X/Ot6NsE0pXjKHk3sqGAs9mhPVdD79A4vKkmH8Lw5T09kmyp7zqOEp0JqBh12WuArHze
xkJdES3REP/XE23zLra8jvFLIdu6wg0ywuoqToZV6MGhKQgTMoY9OQl6uKUAvvEl08QH9Zm2iGq8
E+WFe6skE94M9d7xO+dHpWUOiftzDnOBUIVomR0DxCTAW+Jl3haLvm0w2T6GhxoRCopWGDfbRvQy
27LOaG2MqcaQgxVkawZ/vG2NGMRdRHsG3SL1U9UgHHIBh6AYMjtw4XwC3048M7X/M1crOuSvGCR/
nB8Efl/+HgcrUO7NgRsIiNYtl9LDyVkytuldyokhYOtxUkKo4urA8U+6lp+ZoZ1gKiSVfPwKCL7+
iDA2yWb/fURjI9OIfRtbaohxL/LvLT0uVwsBFU6UNTbVKWtLAjIDo/PnJkwXACbYzjXk80M5A4Da
xNKlJ4wOwTLoifRGxd4OjstRv4z5N9NoBa0/+2Xm88ktx0p7zDC0L4EYoRnGVE/74XqZo+5LbEXK
aKW8I3rUiQqNJyG7RvapCQTV6msMrBTW3MDkNSQzM9UttDHkAp/70tDzUY8UJHt6kSEE7RHh1mG0
eO0do0mkD/HhkGpOE1w1bJjzhbiiS25iPPDJQQ8vFLs67N/AUdfMiWBrZICX6zT4lUTjkhigMT1W
UXe8jTXsO6dGisCl/Cxn1/v3qH0lb3TIFpNbjA3xym0hT1iLFTKAHHYzFn9a3jirQvKPaWcSTjWo
v3ejcm+XQrVnsysbJPCLPakfFgy9YMqu+47bxdRzAgn2jxhuRkES0cdxPkK25Jxewt9o57a9jpPR
LnkRnjif2Y+u942jzkf4NryV928HToiq0Etb+1xIISXY6HIX1FeyoRYnjOm8V2zCN+9pN1ztowXr
MOuIfsp5k8YgFIvtogjqlgMjpx4cjGJbh78DMUq7WCZCHRdYke660oPfutsI9G0B2eHCreFaYgVI
qSLgJqI9UoS3HlqJi514TMP9BMmAjGZYGfi8Dg74/xv9Xj6YxMPcNdJwS2enST+XNK/RueoXdXFe
DEENq0JtDOSFLSuACctJap7vw02CJvyBiBYfjP3HUB7GYIGk1/nBlJhiAeBWhECjmyTLb00WphMT
ctlD+7UiWmnKKXFy0185fTyv0wubXFt8e4eH+22ZpSOna0d+dYqyOIPpsSb4VY8zJNXObhNZpy5C
A7q2Byqw18iQ9ucI5UfpGO0Ex40vb3UjBTEAkYWyBRiMB7a/5ybFUfDYeh80T2ftBQvNBSuLjYZw
G0cER/VeZnmxUNh0JVcfx74zdnHP6Ie1zt1Jh3oV1ju5rv3UaeDfHurJPc1/po+Pm+eBbeDcxgBg
zWdxRbLdvZbMzkakZD4859nSe9LCyvy5hgbDixG9LSaZX9NvVJEQcMgqZ2jA8phlxhqqYExAcO01
FWfSwC/Tl0h+s8trCIe+EbAhFx59V275eADHUp+ghS62fYr65bxTwOz4ndqhtYcXO/MYsjb15DyF
8bzWt4KHOrCvimYT2U0pT1B2SWOxetCdHeD2Rr+5HG1qqYzzIAi8xNG7jSHDRnsMFpX2VaCRxo2W
QTIM+D6ykAZW2mE/PyvEz6FR6BokKjf85IWp9eOSLcwhNFbgIWCq8E1Fyr06qPLZHXdl+9+3lbi9
N83tJZczBwY68lwPVll0+5DkJAUE0+7aPZTVp6qkIeawxeDgFia19I8HPryEt0dGHxuNg3tEaoXp
N6dzjl2vtLsqFRK9FxkD5I/Dw0h39YdsyGcDLVqufBUmcOnNYhwid2mV8WaJCqhL55ELBPNSaDb8
Sib0TWLfZUB8kRnf6LwF0b5pvXAPe0tsCN63zBvns5dP1y7DhGuFLpzFw4R4gm7+qh3hd3+iTjQR
+LKKBx+9ImVmaME8vk5rdwUDu7AoC6doiXFljW4ryt5IFfRWmrulXprIvj2a4ZCS7AFoVH7aYrQ4
hC2eEYbYcqdBjb7ul0tYkyiLA/oP1NpE0+3iAHwDlgFCzwC+jOA/C623feOMoWPmXkbd6W2s9sHT
tCL7/qa9pb3+QhhZ0jZQfS6SLtaQZmz5IvmifdtUMTGW37S2W7KR5dI0hurNVELxJp/hma4Xu5FS
T77sFzTtwRBRgKd/a2x6A1S5dS8QgThoFWuYJeCLGvUwZfCB+vQO8y7NyA9hoX1J4i5cQODmIuHq
FkjIiMEJUnGGKCELqtr51fnGuo+h8Z9kWynfhJmAl2YMJzq3Yu7wwkLr0gyyxMOAoN8q47SNUcAr
VSu2KG52LUSlkTjpHEvpdm8rvy6Dr+INne+eNaG3SDHh8cVkWgVM/pxFMu8aKr8Trvja/Agknnep
9g1QxZqK/MC4Q0kKRP8JbHL+wybGAOlMNqJCSh4AuELi+CaITLC/0zs47pLrrGzlK5aZa2aS6Nlg
gQed/+zwroHp3YYfxN/j0S/prWjOCB1cdbFwJgYG9Dr5QGvXiumj6xeoVZ/hdIYhnCLMDWN9Gd8r
YwthE2Hy1Hbxq1FIVs4stYRcis2V42X3RlFSYixr2xIqBmhHwFBBZBqReZ4a3nDjakyuaAVTey8E
jeYr/WncFVt/F9QwjikdomMHxNnaoFvY/2HasUsTWLIhDcEqiHrCcfFrPXfLG8AO/voFdIVC9ESG
ethkVMnWZRuJE3m/NUMI4lffHkNLhk5ojw5lmZvg479slbcQz+d6zDX1qK8nWvLp++ptPYJGs75m
n402RNT+sUZzipNuz7hh1Xbt2gZ0AQgyWha2neS5ZbECDSQAQNmgEvZkwUj96CeBZm89iaP1IkBv
9F0zaNEnLaUAKjmIcf/BqBUdmFnDZIgTEnlVJNIX1jPl/gTGdIaKeyayxue0L1AbgzWZZx4AL+9e
XP4vu9N+42JhGOxrm6pIc0aZ3Aq49y9rIwNI9frUAu4AQl+5zyJWpUdGcLg262/OacYchmvVK7qu
/097zt0fxamXOBjpqqVWmripRbuTVXAKBPd+DakaEDHN2VKGifC7YPan8gZgDG2VJqpsCB+7fPcI
TUc8lc6sqgngn3rkCfJ3mCH7DPWnlvfusOuQLXryqfejC/m0P06i3I9/5wJjJbdFLlamrqFlQ9h/
6uHJmAuG6TnUGbgmAv5PH68XXJjJJmqDUq5BT/3Mrs1ASvX/j7zqJM2owARgxU29BsAUs0ZAaKff
y+ohfz6nUtwAlU1qbqfW3yf/6au8iGySeTFcc1CsBV8PCdKetjz9gULCh2Gw7eidzos9wjWd013I
D1wHofg+g7y8FCeKnaXqlcQMWPRtIVA5VEBXr21UX9BwTbEThTMr4BDM1si3nBeJt5/Dy5ItDKW4
C5GCd/SJBSn9QbdT6JS/Mzg+u30AfMqTnEKL35AXIynKaIGicCc3GSoHt7VT9L5KITCiO81gI9wD
ThYYwxm9Aj7uJ6//JWhCkW/mmanAkf+hqfrf2+HljrpiDCHrpwgFyvX6SXU57Iv/HDSyJ6oOTIDl
p6By1dWxin9PYcMkRZ5xsaSOZ6TAUX8K8LudUXS7T899kkuAHT5RLHUb+pUTQDsUtwuTMuc0Gwol
vUxFPXBYls7i9NQZMYAbPl5P8wgH3YuPyGdxVxDun5xMMnGHSSOOoBo2JJQoJ73EkAC9CPN/i7ch
aCawPIqhXZskJJlyr+bbbRLZibF/NOLjamwdzkjWGbi6hZ+AarFFlzwwtPLogjnjEa971bTK7Mep
tI480LcmZg7sXx5pSW/iYrgmt0gEuFbBsyJ3ZzAAFv3IVe4ZQdbJrYKEl3pf9U6pDnC7PWa2ER6q
gmTpANRl+z8j31ubeieW4RXTX5n4y1nkFQWsNLNVAZfRmPJ9m60EEUIV16+PDR84Cf/wof/QXqkE
6vgoQBTEoCapF9YB4+vs7+BO3XXsWgigDV4uxcjB4blqdi5HkMYu11zV35aPduqXC2AYVeVPaHfV
Hmf1NnVwhMUn4ahzUSK4nd5H1S0ZlV7h13TfNU97XrPvCnFsIerRmYMgBBYF1vAnas0F65rhAzYq
2HNsKTcsM/I1+yPsNaEqtnBwsTSdDDT+JX8tJmdegerDUrN66ufQvJSeEcxp8rW6CD6tg4KV8UuD
3wLT0JtCD2oZomVTSlitgpLYWZeb54G3JofatCp265iDdw6jOUfFzBrJYzBEGWxAxzKtt0Gfffpp
qXV6KZDltTWoyWbMKI/26wniACl0JdIlFICJ1OQ3k80/fYatwx3VdJHKdd3B+7VhquLdzPnJUfkH
uTRhT4+Rz7RCs+ETu5Ix21/wdfkfca5GTAxCDD4XxJn/+PQKYQjYh+x1eHVjNyP+7yk9CJEYE3YW
yPzS4IvLstE0Cl/iJnKVuF3BfeOyfdbEa3ekjO1jVB2iAVBExLPgoC4CiMZWI0yCzQpAtxGCQxCw
5r1GrFB5y8xNT3j+gD1PlS05wWkN3+Tl6FMWmwcSFGB81DBDe68Z/heD5SRUHcSdV2sYZ7lbaB/5
tIBuhO1QH+9dWPHej7xvlgOwHjUXrBv6geReO2XoSw8gagwqHH1qU+4NDQczwI8ws4NU6bJnLdMq
Z6e3EIvipzIGsunW2iyHNz6fapBpG6yVQ3XIxKWxXhzohWh84KglkOmlxzbZL8o0snsqSSad+/Vu
Wc0EacwaEi01xuWVR5FcFCdGEexd9/vZoLN6V4IAWj884O2mL+abhcxkx5DTS2bLWcBQAiGYwmoE
etixiBdzo2/iUSF+okYkMhkhWgYA99cUIClf/UX5K9qzDMyfks6XqU14Ha9+z7k4ldVQovpRQybu
eTmvksxD3GLwmr4gaFbz/1JuXDNsOzKgbtptqEAK2xwAxUERB9j/cg909FPMbnt7+lHHwmNXr3yh
A/O9aVhGeC4X40FKXlwk52hilfdm4SZa7NHGMCLEZYHMIvpphLuHodn8iJ+ZdOTAHF0fGHes1f9+
TQJjRiqJMUbBCGQB1u4xs6K8XUS1bTkoKqccO/GCemQD83H+62GXjUmTxxlHk86BO/BFMOkzFKEw
s9go7ofPxEK/gqM9hAIUNkWaZpFY0oR6cjHA2bcjzRAEyQaWgWKH8LVoiCtMc/D7w7efV7nfg5iE
w4xg9OvJgFUO6K6/XCqCCW7lyMm9DcgxceB4cLKgbDbn3X2MuN7t0M0e2HqLAGWf4ndRvvJg62tV
LtM8MpUbLFGz+XWfZvjDpiSMsjloVNfp0sC8ClZncdAbm1HjQsl+hLFWzRfoxJwu4XfSEqR6s4JZ
DMAeoIzTE6D9vnp2Dpq3hI6OtxGaZzo9YWY4DIILemmOn5NzQODul5a4vro6oHmHxlkGhUP4YA+S
eg6513RUsa4yxF/ukfXgs5IUeaNBwpexKYyyPvx4xYEdPx0PnAkK8LmxToXuTz4IkjcGS6wfEVQz
nD3ldTJYIUs2w5UHMJNZSmRnKK3AL6dgTFtKqjyY9iuQwuRmg/AbjPDN20wfm5NPNsdpIreq2vNt
kTrxZwd9dAEAgsiiGyyauJImRlAhlKhTykaEZMTnQB17bOg2cM0rdTzF7CRi+CDjcmDObMYv2Aw7
P05YRNm5JwRw3a4CM/Z1dWgfc+l6XpHF2f/An0XQNjC7E9UcZB0ToUek4IRDk58jkUIlaOMTQgvm
Z7saOzWakeYjmqQv/15eLKFmfznX5Tt56h2ndlWLrZfRQDXSFKlBqbjf23pZKrQRhd6r6IphRTJ9
dsjw9VZruOyXQH/EeSQsziQrlYrHJqrSV7BYKPPcEkQoFZFyysL3CY/Lzr2vxbdXTHs6v1rWGfCn
gWc176mwPjhifjdOkWuNoeFkzC11Yx7Q5pTZRIZ+97WjwcryVf67P5erlKPzPPnRd59vOELk428e
kH1mrbOaCzRF9oO6AZNZ5HVSAAdKvc3dPx5oshuJvnh9xlTzP9auSxLE6ecu/eXBvl1qOr5W3rUF
CeLG+iDqSxMScrpGxU47AjQWInc/HjAMcWnNvmtm5zfCBpda2XXUyUkuD3OcJe0y0Rm4h5jQNbVm
DnzU/UpbWyF/wR/mIHegDITAsPOV6PXm4cIwpfv3UJME9yDZEWsorrqFLQQBCZyxJGOuCnHK90hf
YjdHHfOM1uBKwyJ1RdY204rvQMZmBnZiW5N4KkpVO/oLktEEY8aPA042oLhnA/OlWZwc+SW5JeFy
250KEr4AALf6l/kXXekU6lMtkkQVGiTzPXmx6eOgLMYCBq1RuWRkZK5VRjE4/IDp0jJwSQo/+gkb
RHw8OM7NWdfgvtXm2+O6DJGDJg1Au6FSo0WDaS1tchOxP733+aVY1zHDHriwa+rvM2ATAolVWKP1
5liyOGXh2TzbVeea3E0hQVUfzYW8LfD0fCvjR1TIFV6HkVY0WFOt5svpd497Gj24lcS3hLZqmRdE
+rPWrsh4eBv6XT9fVLNKcPV2sZ/5YVt+C1DkUWTk8iH6ZmxLkHH8C9a6JzD68adCYg9qrP3G3luI
q7lVQMlRjvlZhzy8p1MNFnMWuJ75c5osj91qvcSF0Z1GDddP2Y+ALk5LYaE/jcrVyLmZvLstMbgE
JLrWIbC1T6zaMMt6D2ojoBZe5QR422M65pO0HVO9Ta2dPcP0g8kKbRjeMTaOVU1geAHu0OgQcyb6
Bzxby4LXP8DEHp0DTTpkdfuYKkbuPEDls7k/NJpvtiYRcBChBJvrHIgeq0cZLh0iotwgmPCw6wF7
dPieuzfGkXMpvFrHFK8RA3JiWFXWcIp1V/UWkgKDbs9FmKsHCYablMHEeiprlaXPqhNOx6G7cjQ8
ur4rSNA69kgV9/tZw/RYKe8VrWhHeZ1h0EUJFb8cmO3mPMHaPftjWQvadaKv3o3uUq2hiGCjg9BS
3qSdfPP6UgRAmwu9q9FeWy3LvM7UvV4ZDE9XnAN5HHpVGTahjm+NNvk6poM7OT3rUdx0fhL9YEbP
8Cfqz27Qdg5lVWKAZHVJMkvWCc6F0vJMtTEksxd+L85kP/GRkqjXJvzPd3OtiYYF48aYSInyLq4L
5vIhgxHWD32wrnD1Bf66D+CtnHHq51u3B7goE/zl446wKDLcRWzP4kNrQIVx7cw0R34klb7Z1nVQ
VUksKrhDMawu+wTgoq4xPUezsuGysZAbrMMBVEUTSuYsGFP3Atwvy2buH0P5NDdi930efIKWYpNB
SGJoNQKcxvUIfBw7MWVANH454cFYhA2MXhWKQsSoJW2ZBM0q1fTk0yXWkE71yF58Qrz9bcKI8x4H
/Jjq86XilcRqfFgSyj0/lB82eMFaJkzS531HtIYCZikmcT0dAdNSFDBf6DQf3iI+oa8xZ2YmOxw4
56kQoFWPngI8pU26DWP2rTJceXxfdEhOuARlMhQCYTDZ1Uz92UhuuhODb+8tuXN+uUsD3pYVI/nd
up9amqlOv3PZH+QbonhWg03IYDYjb7PUzG7a4ydwFxyrpt2c3KLplR06DScADALtJcSgnl2+jgID
xn+aSrUnWpeqncbpTKEgKtAGxOa8Ltm7I6co4Jz9IX52REJfHp5XfzcE3qi/9lKG4e2mbRM8Wq3k
Fro5gdWS8X5hqGdyWq8SbMM2WCb5OJJFoCR8PLkixJdolcpSY8CWVowu35lybbLF+kdsKqwbNhyx
SkvkF0pf6pYrAG9dnmfmHQFrmudSz2RF6hYsG/CKd6w0FC8VjtrYoYMAm31UgKeMFVY01jzSTK5v
qakNJyJVtUSA+BPuTzbFVJ5Q5Did/9h/ul1M4koOK+nl3TMUdf2v/b+/rbkhIMkzUCNdleNpgQC7
Ygyi0sgruBfUp107n5A40xi9VH5rrIOAsISsOnjpSmd6OTwVrJBCp14qE5W61wm4rD0dDq6V66q6
YLL9mEwlxQdNr/zDkgA6pRH0BrQsvZEP/jFO/nuXMy7jyUxAlBsvblwA0cy9LrVFtgDnSkNUsNw6
e12TrFP2vcd0l9jVcw3U87IFfd1a0U0C6hrcEMcZpbn+WMXMOCYb3Jzv4mMtUyeYTaswpbNsVBnW
4L+GXQijphvhoeYJds9hIqMAQlDZQLHq1S05HCHlMhuYwAGZeF271s4z8k7ELxKLse4M2WvM4E/+
uZwq1/zxffCXv+QhOg24uGOa5lp5UIjf4FXG5Ui9KitpkU5CQHKoRcPOxG2YhrfS7+HxmCgP+6kA
AtXujHnn1JAb0607OdGwX2wC+/0JcPvr7Ke2NmSzaCtGmQ+VmDwMm0BY58Qvhuh2jGZkvGW3Y6Lx
54a+wfJvQwQIHemJ3qsMppvf/L9p2g4hpCnQ6XYWS9gamsWWe1DzzA3UF7Z84HTO8RNoZAUZuAG5
oPrEuMsw4q4U+KkgOfA0vb5kbnEFxbCx8IeT4afUOCga4QHDOq2TVJHrSJ11gM/5p9uSHYISi6N5
rSARHHmmkuQIkJ+StF8wWJLABwnSD3tFMFdUbkBssVPTTazKMPY6yIwt2+6EqoicpOCyja32fXJB
6VKfH9nmhzoBCv05X9VUsN8GlEp7EBbXiv1vz29W+lZr/cvHIUgIzmMDZGBeOL004euhtrXn2e1M
5/4lGyBddxxNY9y2nk9m02HcaRbWwB1haR7t/72R8Pt7s6lStm1jcizSynaWzfY6soRZenaUrN8d
dJroQ0pEP7WT6l2wkSez+XL3HZOa0q3gX1asmvlY0u9G/A8zQg3fbvLXEwGdFPuwS06w1O+s3R7C
WhSTuITR4b82UXbCnNu4Zqgm7ru3s6Y4mItGhTxHercnAa9/MehuqdRx/mryRX1fnurGNrx0BxWt
L2Lz0EZmXIy/SqAOOKWrsiULMzh+TX9MZa6mMFFxowcKqgHSfu/f+8ya55hnGdEfmJEQ56PYIZNW
CVlMpBmhyIAXYTqRWjVEfqgW8nOBUEQOiuu+Hm7t8V/6fgNJxRXmcR1kGvbo1mJC/P5e9cp4IYxV
J0MEUs9iBO643jdh5oShWu4yxfs0FQgsq6FthAMMEnK/Vli4vzE9exmYa4o15Rlmj8tsmgWibwRA
oNRUczg/fqncJ++PLsUX+CZ4FE5OyawW1dYrXPZhZH989iZu5JSAbTcwoBbfOCRHtL3HYFQV1pyg
405r0aYks1sS47FBxHH22QuPIqqcv8F8xiP0QzjowOlW61iSWItxUrr3lDoV2cK883j6IMT2RewQ
YMlIrFm8nbki2UEbww/S1H7DD4ie3miQczDhK4YxxhTfto72HKVy5o4MLgfD/txnR4c6+45YAF3F
bEGuPUYrztSjOAD5wxGKXEiNobdl14rdAlXOmVhP49OIo9AaKvl6oepnzWU14XCu0MYNz3fIok0g
/mS+AmcR68Ur90BZc3R9kwFgLe/NdawrA29DG77lcB1BQ3+4rOevK458N0ppHA4KX7FwqRQg8ew+
1XBZkMjKVA6WHFz9F+KjrLWunBzA6FQzGe59sUN1mdbB0J/57P06nTF0/5bz5YVtR3yeIRo8Brr8
Ac1qWp5dvx4dAJiUIiN24e7pUyGtUry3CEGAwuZV9YadtNOBMT9N+3jTeYM9Si7SvdOnwu32vuLg
Oo24ilyv1XBaOXjUUdejFwSor6q52a1wZVmagYH1cKqhkNp03tqxPSuAeuj6vADJoRTRdUCl1NwL
hWZlsTq7SGeySa+0VtshSlhtitiGpTI+tg779sUK/8OlTsakkB2oJEtrC4pspj/PXqBmH8NngcVe
1+suK6XE9QBzYZOeooVn1rtOAArqnZUdc3adufcOPJBLcZhBtFC7F3nBEUq1oA3P9bdZYEnbyXKp
N1Mon1IFNLB/Zh0NzCmJlHqAA3R4quMHzSrfSrBX0sj+BFMTj91NCjfnryMgb0ZJEwbF3HbexJxT
jWI7UI9HslwH+p/qQAYxNl8YEHsRmM3HRpw9Dhjb+oiunRUNGQAbkOuIPlS8UaV1kgE5cs+l9yd+
YWdx0xpe5Zo1mjnXh7JDu7cJ/WOoJej5nZDNibUKb3RfBpd8fCOUS7NVkblfpqYoQOVXry2A4d8K
xmZ34uqPWYGcYhuBWeigHAKpYvVu5yuR2Doyv6Q9zrwExXisdDm71dpgEv/a6JBBNWv+49YYTrTF
KaGEpOtYslkBz2YuA01ReiOfmexUcGnErVg9IFmtxkv9SuDK9bBokcUmRDAKj0LCSTekMvNObNjT
IJ2sglzPlr/qz3ag+UpVAQsTPOocVWIJD83IaJvIRe5u7ggnLrcZZ0N8tsPEbIC7fDPJgTtybkRG
bmk85HRLVE8HY+O1FEoTIP+rsUr7RPeVRpH24CBq/HlmRBiD+7h/lhuxaug1YznlepoT+nMjPIQV
ayP0CJljnZhwYYUVSUAK1fwDH3i+t5vVQmCYtsFcL+WmpSPMsbvN6drQw5ZPAG6/6TaPtoXnJxLg
WxSRVKe1bFK2r07UQCap/oFeGTM0mqBSl2GUjucro3ou5mu88o+d51+PYhVbd6vtNCRnqXvBx1w+
2bc2gBvfYRzeahqkNFgxjZr007x8JavXxYiwbZkWjUUhmQgTfw8KPh/YhSqhRA0i0T81pj5vCDKK
6stF8F/ypGsF5vDnY50LP5IhxDBwaXL9SGAhZLYy/IcYjK339x4OX5IwuKjd71CCsDjOwsEak/KX
sQGpLn/zZbnSUMzSaeccl7v94cXwyO8GXsJEArnzFp6wAR9bXMYmdD/CynyxkhmJbEjFgFxS71nY
kPQH4pi/UW4+24KGbzCacd2M2UMcOtQhJI6KSRAysle/884FGyUAMfsTE9WlWfGguTLvlbWuUBt7
1ntpLXXxvsdDYYNci8OFB+H59Cp69JMWcscco37W76c6CQodhLEUkjbOxP1hxSaqcAfm753YB6Ba
bsl2xV8wlxQFb0bWcESDHCuePGlj5ma6pErvwYFqSU9AZwKDtUoZISiV/r6OlQv1T8l3HjVNmQ42
VdQJ/bIV2/kPozt2fTwdlx5ZExoWpW6Tui5gDBEvbOqRTY99X3iPl7Lnt62E+2bPNJw9W4FiFd3p
sddjcf2kQVhbhfS2BomBA9vD7QzPQ4tYsPd+ZAicNJ2CIW6lZyPWonB2dA8hwgfjjhLtJVeV/his
TSZVZ/T9rU9R+wno+1jam2HwyiffU9mpN0F4yKo5cTqbk/nFeQFOr85NtBwiRv9HyRa301H77RBV
T63/YV1Weqt9GofjE/92nfkY+qoTT9Ey6pPQ0xZnBZaONgQVDsUlJElnHqm5nxrwZm9ylJ+rwqxr
VoaQllZ6demS0oeHo0Li5pbYMwk8ObiU3qWUvhLfGUCPD51HN//2N0uPSI9L4QY56pLBqOzikgCd
Wp/u4BtNjOmuhNBv2jYc4HxRQ1ZeDNyljJcYjrh+EFlDVM1VmTmX38wvIjzhFbt14ZUXIVSed5m1
lQ7uZ9tmbOkM28YAZNyCRf03CM0E5WOCFcAbS3Q2kEfRJf8z7Rq4iHCRJj3lkVeo8VM79Pf9YfGb
/XhLmA7DK9rKxeiFFTCxXM4LlG32hV/wZCMch9dvtQ07fg4QibhE8ADSwGNsTqH2auyOMJukUXJQ
hF9acFd9aNVvNdXaptlDcGZt4oCU7Bl9AJcTfTq63AtgW1MwRJWRr3Tl+bLfO/PM64C5xfAK3/rd
VJYhh3qAsusluyOU1zrOoRrNdE/jpVxXOThNLeVIwDq1c5sbCZFhNjGBUN/GT8WTMsaFI2ntG7wg
TYz2a2jM8nDHMv+p1mmRueIBkF7CHQXwpmZX14tdc2vFvUZUVj2Z9Ry6OnFY/SGRblgJGApSTxLI
xZaOqWykNa5EjOyXyMLC4MIfuBZvHK6QcOxyLCHPKPUDmpPisQcLLQsOH7pXXl4Kt5xz9qeqizl0
KTVYU1/gqmf5gPqz5GGMlMwRf7PHIuk1wMgjuNBEAduIlo+yDGco5Sj21OC/EIyNffppJeKMJoGT
tLd0C20joWhZAacl5yMmrfxYHTG9/KrC81ybS94NdRX9LgCEEvQxevqdyg/aBoZfsKYtLWLlGjOQ
1CZOK6+Q6ugSePD58VvRSs5X+h03Bwps9inWc4BX/caoQtnbYSxl7qUjTKCD0UpLb1CLo2DqODN3
R3WOlG30Vdf77D/z8xpTOjZa1UldfrCiXdxt0B3ZMoQz9+FS1G/p32BagD1iZop0nOAna0ZpxQ6E
rOKPcPEdE9+MgUkwzrOabdv53Sd+6akQ3Bvb6E9GtBsBZMiaE3h0A7vJXgjG0i9s9G07lavuQ572
zIUPxW0wGjHUqzw8PwFTrH2ydSvHw6ZaUlUN/lJQ9uCmX60kD5aEIcrSRSCEsbenAZ4Q8oBFerp1
7Z+NYePH7Y7b0LFpDeBShdO7TBksNUjffsqasfV+fe8sIQ0pnA+yvtumi7MqIH67p68Pq5wQXqSe
XHC99CATKorkqXNQnPrejLJlYF05yTI6zSc6BRWBMNRoxBebbQ748R20N9a8D6+SgHcMlBo9mOMu
laAFtxzGEOhKsfNIAUy4LSaYbpKfqxmxLoCa/sOjF/4NsYvYAP+KWbLpLT35PA1icBsjwJ+t+S2b
j/pG1cJETIOFFcaZ/QqvNgRYew1qZ+ugWgytKYBXUPowHsHAyKTS0ilHFKCkFrhRJDICnvnER0tA
yBxaOcaPMUu4dfvO16l9kAamORlI8TG/p0Avq6WTAf4wl5Z3ugJ0uITXeLJkxGXBNlZ0QwSD3YAJ
D7UsJ2LthE8GyYW8F4CFyifsbswQt2+ooJwIfo0zYi6Pil7T9YojoWSAVRVOpe6qTADP2e94mGxG
MDDhgvdtF+z0HozcpHcTWBpw7wzA/N3G9ZpH0arKpEeVz/GCeR50dieWT3pIZix92WmvxPaO1Q73
aNWENuiqCECYHL/STmtpsrGhrI4nCblfvJVlhECJ7VBI9VcXs8dkOpnY66dlQT9hP9hZZUE12mRI
Fxihm4g2PLIVDN25nPwPcJ92vX1gPliIWrMzOvbNC+jFlw+UdVFJ4e2gFvnlOOMv0UXZBK3E4uX9
i+qyq1Tex57LrYR6JuwlauJdAaoTbEWv5hQaSM5bF2g3aoy7g3e0nwWiwDKCYvuxIwPut13Ja5NW
Pu2whotoqCMoqa4x7APN+8LE3lmLnIsYdgx+RqkXxuLT9BYGfYFw+c2vmPCiJTc+bFFJHlVVULeg
uxF3vx7aiMmo6Dai2lPXnjg9DWPZwU6vyQCtwYlicAppN9eqrcYP0PjU6qJ2CdkUO+XxHHSvrVmz
VYcbPBLcnKf2ioG25SK2rQPv3PPlLn2TPsk7/JfLQly76QV1+PE329B9jdKsKz2AEnmc3d95qOMZ
ensZpG+mLtVf3jx+od3q0Gphjo4cpFzoT52Ujt6X+a1e5hiFomvRRs7AkRxaqfQc61p26BUrgkmk
nB2DbFfT/6UzKd23m8HJ/iEfILl+eXq9rZvT2bNdXI79YI5GYt+YRvGNad0HwJ+gLv25gQzcZ3HZ
mIS8FoFPC7pikCIGDmAm/jOi+Upv4VXpYL0Xq6hoJX7VUo7om2abm00TFAvsRjI0F0FxtQyBsiRv
bWEW/IUCR/kLuFZbLcfoN8jz/X/tqOeg6gILFrP3/1NZGvR9kWb8RweTUIQmdBhAf92lrLAzw42l
FIDbDyfn8LPhzHtF7wQcORTftbdSH4TisDTazIT5oSLhP6rS8GFpXJ8ijJWtYKaATGjMRRHxZDZU
vqfs1dDtnIfkhtpuGcGiAjqsoKBUjBNdjamdwM773MmWoN+gbmwXe4s6GUmYiS1n9B/GJTIDzghv
S4WCGxzFBwOQH8ToayOS1MfwQHTxd72xQFRpKSI7L3Brk/N/bxHnzQey/lAX8V+lQx7D82Kq7MEq
/GD8D9BAoq7OBRH5gOCtJY9EnK3CSxDXKAKjhWQ72OEfco3e+5kEx9/HcfRWQFBw4zFJ9MxsiBwX
cmpqiXqxR1m3tkAinJpO5NNzjoLBwSjfDy3QVaR5iuAEpj/K/O9DzBtCT/CONOx2THR1Y4TQ16dP
9Hei8SMrw47ScD13FVEwJ0GubW0pchtBNt5LVDEymVTO1zOMsJoAlH46pMtEznqFdy6zPFL05RZo
0Ys9rp8lKPLXzNbXX+hpVHNedeaiXu/Imk+BNkZqSX9cPCuJTuAXjbZQyIf2C3owrZT85HmX+x2Q
WmT03TXkMdgPs9JiTuPypNJifzremyuxi1B6kNtZKyPS0EEX0BwP3k/uWeVSvT5/yBffN4MAlGO8
wlv3xylCx9CBjCqN4AWZ0vAFwyfdQ3C+T8mWvLIj0u1CgsQppRJUbOCZ23iF9wiPUWYkhI4hLLEc
i9VZz1RXUCGYDEPQWDmXv7dWsABI9QxBMRDuGfu0judVjp8TYSbi1TNd84zdJYjC/+Tj2pbXm0Nf
OYEfe/Sdssi3k415v6heWJzv6a/xTfPps6N/wiMkvK0kYknZ73dhjKaeU7RDwad1+Yju/z7zhb/e
3Dd3QuRx763NAuE8SZmyInQjom0V3nam7XnupIjmY7UYKeova7U3JKDTLOY0AEB4aHTCba2YC+TQ
eNBg8ZApqizTW03CIh0ADCOZF7kj1/00fR/dhQFLNIVNMeEB5cfLTy6NPl2TWvck4r8/te3TLb0t
peqEGM92ftkTcKJyge4GO439myugSpVGVhs06d2MUt+lkODrCslhyt778y9wWM7Fo3m6qOIuDWiY
6CH8MBLJR0q+39lCPel0Dk82hQDd00h4REIM3hxvw5CU43YoyMVpERlmOSWL7hCk0eppmlM7Mz8+
ZGzrzPLYd030NwnmUtgdzZKFqL5SyLBaPDMzY6nP9PudpffW4iK0lAJ0FNzYcK5cAldHjm8QX3GS
gWeducQg5FrBKXwAgAHCz4e7wuPqTWHQvIhv3g47j2xsPwTfX7akPhJs3kLaBl4beZC0zFxF47/B
/3XsgMZH1zamh+Re/sV0ktkCG+pE0zg7/AyzuyaYeJVkdCqdsjxQt1v6t4bZ9WYsdrx9OlXDz7Vc
zhoOEBI3FM71SAjAyh3ZYZczkJcEMuoQjw+C2WYEiE3Rz6j7b76YJvj1ihWDtN1KxRpye6iAZO8q
2weyISk/RoZeRTnsZRwdzM9179ztx1GmGW32unEGsTn/KXTaHvGpQHmXyXwKfokZwJJ/pfvEsPZs
23vlEr6FmU9tpNDHDqDjnPU6SZDSFTJ2UmVOnso0ZTBMeW7Jkr+Mp6CXp4Q3frKABS2Mk3p+3gCL
rlH12ZKzEnIr4gehkUH9hp2RXQQl7tRBjn3vFK8rKO0kPWpFHDD1ML3CQV0DFD6Bd+aV+1/zC1Nh
xWvaPzP04GRyGCMvEq/jQn0iuV1egwMOkap28u9KWtFy8435HNTXcEwd38Oo0wLgIBYeKviS/Une
yHPHSIixwkCgQdfWUHXvmxgD+ICTRX/tqLghKImA0++QeU+O363+NNvOusD0fGK3ohNn4BrLao7A
n8WkjGFFk7MBftJ19l+LUl2r7MA/ri+8h4gDTFO/8UK7m5AsqLpKhrxp3mVSdFZYi9ndgeZioLZ1
yoUdXvxZQcKuitzmO5DiZtqXSQO979t38E/Pj2ji9jvU6G+N+AsaXXO1tTqZS6cyFjtHoAJUWsPa
pyNRQh4OMnyqINHQSxgeVZSsG3hbiyvdxDknnCYa0KbfGt1XdADW96ITDyeYQGSX+RxRNLUTZsAj
08am6oZfGHFM7CEZHO2SPTH7l/EAA4MXggli+1X5hklRdqm5kJhYSO9VGewwCae9ZrLCG6C3W+c6
oc+dhnE2RUs4CHvPGW/H3jwpRh1URb/x4CgW0QxtrMQ8LXJqe/67DLkl2nrZ4wgQ8RRZT453Vkzj
SCu63Wx7vft7vyAD4z3J0TjG8SF+O5ECwjfVegm2gjDypGAJPLpQeGsUMljA/qAJ09b6OSndq98d
cT8mPfvzfIMR+Z/xPUNfGLPYn5XUsSkXUpmH/H/bySllfevWARXd0TbmT0T9urkPXLpL+bpR3Quv
pN4YtRZbDs21Mug+MdzT4K64IbOumXJWoCo1PeX2bhA0WQP9J+WUnUQyYtk5SeowcN4JKdr35sTm
wstLyisn0sIpaJvlx1EMWJs5OjxMgjTD902PIObuo2RsLOuOkVms9FNrPidkyu0Y0X7KlPF0W3rx
eAJLGI3b8vklcVapu+NJFl1y7Htgy/IvKTbJmUtE0Rnwcc1cL/lHA5aqEn1vKp5DHNAiQ1vMCwTC
yha9zEd+R94rAEIO0XMoPwYQGNYFv3AnVxDLSjywucBcXVsB3yAy9Dx4ouU0VD26WK7Y+oC6UYo5
VGr9j4QwtdZPxwqU9pSckErLB7esDQws9cKOXdSWKiUuZOLA4gPVzvAtUu1GxCqK3gLfsgGp534D
qe7AMTRk9C3JNgmU7CocEpDoYLki7suUWT6lPPwkozakorbAuCYOdw0eDv/PUJsixBORmM/JR4kW
6LorAo3shga3FSpDvYoMGrGoyiv5fg+Ad5iK75fclUm8PgfGFczw6j5jy1SiojICgW/xF2DgOn1I
6Xca8XZ2gCjDduVVdnmkrQl9t5n1K7cMsKcV3qJ75QUy2vnvM7lP9ydMUisOt4hq+JrVUQhtsAYS
+TrLpqRKnJYiayC3tgxiCxdwswgiWiRQ3/7B17wZD/3lg4RZa8gT8Plrj614yt9ll09JV9Jxwjv5
P/hv6TXfPmC8TT7cQYxwhFfUVtpSw68TY8lkph9SaQQ34RXo76tk2zReG8e/Q7iYOW2hOfWxUyPo
ABxf4ra5DLTMXSAlk01lZtH/2wRMkEYOYKEySMRRB0DPFZHQctz3cdfiLw5Pqq1Uf1zsK2BBQkVq
Aknu4YmpCeTkHvambSX3eJXMrmXkg7f0uF+qK2QouKVYS86OvOhHHl+4qHqRqNsbur7qacYTcRcC
6Cd8SYQPJgmsa/a3PgsPawgXPIHSAk7rofhZ0IDJf71fTHcDS9tl1bsVEonC4o69digoY+WjwfDa
7dGZDQoMchDlO1zBoJ3rw26er36e3FyDSUdU8CJI3sLpe9yKAbBdR1rKPdBbBfs9AzxfRdVkAJwM
SnJD3yXTG2i5RGulXHy6BVkSfgnxz+ukEyxb0FwHNaZON+oFU6DgsCP74VgikNIpk3hltiGsFtL0
OZYpkrsLO84Be79w0KiVSq/cUsi+sBO9daCoXk1jFVe8y24VxLwiZuSu5gjcCS39xwPrVK/a3gxt
6slNX7HIQoa1xXxkUj4Nn8sXMrJMhM2K/PDfk/sxbIos6Keh+ZTUc3dCn8dZBqxH9Mp5LHnFEAxN
G2xneKAg/Y4RTlslPgyf7hOJeeLCmVu6oamKO/j/0mcBalE2G+OmFUM+C4GuHdtSi7oafWEQjc1O
C7V8whTFdI00Qcgif/kjR3M3gpAGUl1IiVZmW5MY2PQkiSo/RVC7q0YDg3f7gn2wbYrMd/bYyvka
pUDfTSplrUir/W5/9YKeRU3UkV5LjzqXiS/qJPNshsJixFwpMuRrKqCPlCuQkpn56spNfTGPFVlH
Yj42VqyS4sciGN/XmDUCnutXH1AwvABDhL42nBqKhjZlb4OJlydeJ7QTAwvJVobxkqHFABZ3Tri0
5IoG0OnHsmDwg+LXGYaiyhU0P3zADHgJUR1DeZEx5sigcTQKcSd2whusfC1mOjHio5l3J9O3GmHU
HRVghaJGczl1KXdUaoiA5CNL4uCKiJHzuofoJl+rr0gBmUjB4Jh1hlcG++xptfIhmdzIOuJZnsrk
/B587wF6WEQZF5D1txmjLWICouN0O5c4LVN1FviDonvR4Nn92EuvxAaFguRynq9fsEXlZmiALFBI
3JauEr0APji4iTSWIXFUVndR/0qVDybVhzzz/Lrh+ozFvNU0qhz8+yVcE5J3/PmD4N1nq1Dselhl
Y54rsqovndT/CrIef8EXvXherUVtRy+sXdS9NnutowgulQK4wf5tJxzfNXZXqQ+z5DBbtx6mGt+5
my5HrQ19vHhQ9TJZG+KH32qArJAe7cggK8zHBJ929gFK1I0bQ/hJjLO6e1XcLlEozi4m/lBuEAmI
KyK1DgqK8WZeqilnWqa/P3SFS4TKTGYwwssGdpX4mglQhb1XqzsSuMuAVyB/QGHT+GxqtFWTNjkn
BbNnQ+0Q63Iv/+QaU0UN+b24fNPtWLrYF9f8BiDpyzkHtZp79qVzAB5WjfIrtfG/ULG+eDgDg0mo
eoD2F1l4etMlXkRxhZRXPcbyAc/crVCn3cM1W4bnJmhV2eRtyAH9tOOj1IBSZKSSVwZBYGxY7ppk
gJY5hYqM4qYIZ6dkshLfcyAoUuSlZXknaTckOC6wx6htufMh+77yTNzKfmRiEA3HpIeJQURupPyq
mTnu8l/thKYqbaS4yvjrv3GIy+/FhL581S721f7I7fDWHuCD36UhiKXYQ2LgzTKLN+naVm4iswGw
T0MIKVWr7BRVHPCR2KROqqNFVFy3NaAmFgomtPLWEJM2W43e4uElywf5sp8Q+t3a0PD0XyAuznLS
TOB73P9WD+5cqeSzxRkp/BIcvACF1b/7mMKt4ktJg6+RUktJ3RXJYqZxtNtOdVeq49PJDt8UxGbw
m48bf86LR4y97EBAPD1Bq06TTq3h57gRzO/CiJO7FH+jGMRP9NigyUySrrMP0CybZYWY6/celmtv
yM7XYs8I0SE12NNsRZrMxt0568twjXSvca3Yd/2Zb12xsjmi8N5IbkxDOeI9Eu5/G8cF6JRBU7Mg
ouSBIxo5wdcHh5sW16LscYgmionrncJjUfcC41s2ZBvT9IHWV1Kq37q9r3xkwzsUPGxfuarWdVgH
s3oLCVgWcBlWgU4MWt51F75QJZJyo0nO/rY7WFz8/YEriRqB6P3DlnIfMIH3gfpci0Z8d0HmFVNb
frZJISAYmFWemDypLR4DQLbKZ02VPsTx4mHhx6vL69bfbSeSK8ZgUjQUDYj5U6F4XkpO8aBGlwfD
LV8ZMi0PTf/S7DdhddoQdpI5Wf+EnfPcsarvrMAGKbo25kUoqAOjgsS4zuCLqFEXdenIRjwQ//wS
tmL9xlcccaQ7tlhx9pUT8/uTl9iPraMlbMIfac/hWs+20nDtDGfiyiGUJmeiLF+B2ODJFc4aFM86
jC1f893X7GxMhDf8zVnAgAkVK8Zv71m/9CrF9gDXIiw5NqWhbsStIpsQdY6byRdgFSJHZUDBEKYJ
6PqCzpkvZNzIbEQcC34obz6A4ySrO4xo5gdR6LF38mFbWE1MXIXFeL/kFKXdFQhrZj98/owHLeUz
SCkhcXAFOWvB7fJcAwdX/DEAOtE6Lpc6ThWNnPyTVLMP2lqa1WCzyGLy5FA8oRpEZ2Nfgb8wGPUh
0qRk910J/vxd76wOFfNqmFsYO6OR+ZRZ54gETmXTXDDdn7Bl7cR7LpdrArtDCk37PLOp7mDC9UG6
ixU1ep9HM57pFq9UZpFCkd5aIRq9mNkpwJGMmEAIyK2dANFIcVi897nbmKsX80fre9IP5ga64ORt
IeIoNGsjx5AjmEC/okW4V2306zo8nD3VB72Jvq7ZtQCwAUip5/DkgOG1Z/Mzh7uNSqYxOo+8Bkqy
i3oq6j0JBw6Jr2vBfNq1vde9Xqx82ur+eHhH0v7uUvnch27VBlVodmwE0VnLFoY1cxOEf0v8CLcc
rOF9tD2NN5IcGET1iSvw9ekxbRBMBzXw1KxT6aiGe1D9X/IEEk8jrqDORD3T8DHLLk2/eBzUL0Bn
r//dEmanOga+0VBHQTdyj5i01MWAkzv7E7krbGIE7EKB6SIWJ1A+6IJGW6l9jYIgFzl4WNTORWGL
TIhM2LNXfy53Pqf59Jqq32NzXuWNQUIDH2tiwapoUYyQezs94TDx/JKy/9s7is1pE3WQAc0erBwE
pv9KLMjDgSzRTpq49DcXMHlK8l/nNbOdaslgHNdGHYrL0dcEOZWmyOQRrh259n6CTa7GwAvU6/eG
8v8p98QsTVwDnlKpfFYUmpRdh2MErN/M0u/uGZ+S0S/svbtdOtYowkBCL+7Y7vL3r9stU13tGYf3
XvxA8grZfhidAU9g1TFSS4EzHe/fzkgUfVPDJ6fnvNma5MqRYsp67BOBhTGiy2ZuoKrmJxhDisas
jyEcIyU0abCmZQFqC8KFNi6RiPD0BPYoC7K/w9U5Bidi5v/AzntSHB6+IrBVPiBCV4++YxQlByTz
zNNthxp1s+A9mtZ/QoKYfqfOgSpT8ewqzaJHqYCyWuUtAucXsivDnGMrkyTAZzNX4OulibEx8s27
WiZvdjkWNiGoYqmN31lwy5LHMB/3hZjtP1yX3tof2HzAK5AdlSae7OIvwvrs9FHf6fiwNPSN2WdD
Kz1OhusSWemb0m4f9qRb2/Sz2tLotx/OTTT/CepyuGrucI9PkK7NSUUTOL8tkok9WTRWSU+koy0z
RvXR61h1O2fxF+jouYODYgWagQ9TiCHwZDLTRxPulOxMXCvHKzxptlzzdvFwHQ4q/p+h3jOaSaYo
JcrOVP05VRBA5OtYKsEm51FmorNKGj9w2Ul4yelQlnDhe0nJQctVj4FmbUENnthS77gYmrjJk1jR
lPBlXtRWRXT0UZ/VysKSO76Ur704f+R6asV48g5hWxktV9wvCsx3oi46nVQT2Qpt3dJZ5LEiq6T7
/uN7tdBcUKmC6f67RbJVmuQuQKhwEovIh9iD7YqRfBrZm0LxfQ+nGQODPFqLFDwLHibDqaAqJ5BQ
QthBWyQLI/sPt91SdN+92WotLNwdM/XJ4RmaBO7IsXeuSlaiJZuBvuW1Fp/kyHI9GEjm+vk4vOC4
JlcOEpeWDjQVte9fYDdW7WIgrzN1CCUtUa0ynWwMob57stfBXgEx4GNS1XfjWlX2kTqnGdmOehTP
kHGGGyduqemZS7MsSToSvP7XXNFml4uXALweVZiap8mK0dYd/V9xveZuRakmUN/2m5wWXSfO2Trz
6Y9QY32d1QsxqiKLj6pxn1CsrnXfJ2y1pT64+DJpW2uGrvg+stKI1VsQlNAXPU+CG8bfyhyA1AZV
5ShnEA76soDIfpvPc0AvyTWJcoz4zxSNhAFSxEQE7e74Q9Dyd1xj79q9lhaALemfQr2q+SSqL17A
D1VcPjVcyu5BjaHXVxOCNpGRzengq6LiY2SxEeTHI1Rhb7JrOeP8zuMVqGOaVqZ/BXP1la5n8eXi
rJf0m5sMXVlQdLcGN9nOHw/njIDlZzl7daTKIPC/1RijRbpFKO77Ew9hkqn4q3fsEJu2cFw7cINT
ZDO5R/Kj1rhDjUIJjEod+pHlagZsM9aYE3Z+6nqNW8DTvoS9g8odGw6Ye/wBjxvqPDFXM7Txkxds
bNF/ShVuyAwpwno3iihOtAS9v65E1t98d7/wnoXEfvRY+llDQ03gHt2yG42KvCfWfi+E76pgv90C
LXgD5ikMJrtWsYnfUJJKK8eu/rGmUE7NEkJ39UpePDWsbhJV3dHqir30kIX4XUq9o289OCbW3Ozc
LLQKLLc7vZaHG66v/u6md+PfDoqJsRLAPe2GzygBl8qp/LnHSpVx+/SKgg6OxPuUpy1hhtGHq7Dn
VnwmY/GnjpL4/PlCjm4IHFuOmJVF1j+AVr62xnceWWenttMLE1OM9N1xRh2W11ZzdXM18vrFs/Bu
3xKNTeBy5ztAthzTCxDcoSdXReyzFVrgZCofAfmHdAXC6Nws/XETBTW/lbTuVQijEmZAPkFZCxcG
c2K7nETnMFgY1J93V4fvQQW/Zbpy5HxvFVjk4oXEQ3olqWZmzZ3kkSaZQxj0zjLfPMeEp9mWLsqd
mhaDqjYpaiCusO6l5gBFO+fzaxbV2ieuW2zRpq3Y+jCgDFCtT9qnw4MFJKTSHs412QMMQ+YE8tUv
HdEi6Uix1STHRSDrpCwpKPZXI1ntftzjOvz8Ze4Ieh8UyvLqBVgwHh/KD3zRmTSvCqPICxC4rWfx
83olnMRrwUNEjifT1V2EAmeIagBeNH8nWrKPdg3Oj7OmGR32MsKadDOY9gUpimeizI0728j/WCvw
bfqA8+VhE63GfZmqiIKeQOstUs8Cu/Fr5bkYRg5Rqz9ejh3lJ/myVG62AT7XbR02ZAIQF5ZFxF5R
NYL72RkXyzaDSqeKWu1IKuUuenv0+JFnA6vC0/8pqjTndZNU3sNgqRPPOrCqHa/pmaIb8jD/GuyH
2BwFfBrC1E4NXANjz2vVUfFRiGgzbsZH0AEtOircFImkP8DGNkSQOBHMqG5WWGno9IWtmRo0lqwy
qRzFFuRu2hTwE56MG7VXwJkP5wCxmQ9geWgKXkODxPkfwohutnFZTzeHXn0uEZTAGTaJ/kcXiNek
S4rh8LVpkRovmqZxLDl1tc+Ep2hBtkSrI/4q1GoHhRGeAt7MdA8gNUgn93mm0RemIzM5Bv2YF9HN
PXfFGrC0TG25tv0SB/kAJ9MBzVoOnbDVpw+LTpn6KAoKZWQ52b5PE4Nj0brq1TF2zygm2Ab2MQnO
bvHMtfOikr8iFo6CFZY1SMt794o16vrYGVt31DNnYh4tLAfUeaSfJC5afIMrrI7952r/paaMbmGW
yaxvk6JRDvXguS1M4KkDigiguXssxnyqub+ZsW0XXowXgUP6XEli6px9bbtIwr+zWng1GRgMwk8i
WjoAbJGZWBfu3stvuWdki4WaX9uOWwVwK8VcRl6qgNbGpd7S1SxUJWmRrgPmDSNDNqZOZtFGSqQX
r4CIX/PHv8lk4ruM8zGNhGhlb/75OZzQSoXVDle/B+XVD5jNcXsc1NZvPvA9YJsWhxX4un8pffOC
byJ7lkRa+AXs8jg+Ub0HVvk3mHoP7PdUS6wTXoHp34T7yWBm+bnTopIx6MZtnSEItHyohLqHIKE9
Os0GFe897/9yni2m9QO99Mizspc/CxW5M4jmMh9/1heGk3wEO1/hIp9efItplphzVojjH7g8TvmA
ErGv302SB7TMBOQoKBDwVU+xjtWlvfwePPINeanXJaHV17Zrv0PDzHvKSx3RjSTWKrpGalt49+Ao
6laY6ob1/17k0MHH2OwVYozXSe+fm2KUnbcfm/T1kHQPSaBKxQi5iWWk/s5DA0TlYGQaiwNrOQq8
FfnWPTUSiYVw0wYrmeCuyXi2Nr2sNGjXufJzm8pS7KRE3TwZYzTeucA5N6S4xE2kjvT5I/CrHTuY
F7fDWaQPmwd//AN4vnG27KmeHiCpPDcmnzzfsh4LijcWGiqU1XoO/I/m/fCcECamePO3KIURwdjA
lG2+655r6KhIz9Zb02/Zvh16zUq8j8ADwChHXzE6Uv9hoijKaAeUiw6D1dsy4RfGGrEJdcFA1GbK
Vkc9Ow5hcMwfw1wnege4KGRC0DHSy0fDSAVT1ugQaZ/SCG2CSEr+IaXgKUXknAShP+ZH4vydCpmn
ncwH+SAstJp+JnT/5whIEMg2FcdZoCCe+WGvKKu1V110F54zNDldiRcTABYDbaYxCIdpcHlVKOvZ
Qbsbelp5CFxCTrRO95uYiBtj+Q+QVahCJ0LrieLCMrptkStwiIS0F/w+wAv5UqpX3oQd06ge8o2x
nQc0bu4yfVfpSsSRYHxiaiZbcXTgwBuqCgpxez1zAR7FIYpzkNumr9qgjXT4/gseBS+TXX5+KNQK
V++swCvfsml8WNsqmbd5Z+ZsfLPFCvj0egl5jCQn30OEH0rOgVFWGyDZPIjApznLa/vKMDNu8GBX
Owr0C5iZizF9motmlxvKzR22s6lCR45YEhty4xispXME97GtDn0Ol3NhYbBqDeWSkvj5YRN98iUm
C7PKDoBl5OaYjRUHbE/miP2qDxO3n2ypPGCtQGCyMYVDEEFxsm3zpJ6Jj3G0otkk8Y3DlFrG1JBh
TazbR+d8QDI+vr3iuPJpKQTA1GJPibHuyWSpr/wCQJYZRTVhTEqDe8oY8CSAzNxop6+PQyYSyl2H
ecNpDYjohs2Z0v5oYW9unlzjt43bZOgGV81PfikB77J/4oG2c3fVemwXAqk30QBNSCfP5m4mgiex
wVqaFBclIdD5cQ1cD6B1MgwTTaXBvGn66fjqr7ZBTPzplquC++uXCrFlO0i2fONsRKPXL4QHfteK
+qvo9xKISNO+TRfR8fBLUGfyZ8EzZvFbmuPeUzluUTIehfEjnZcM30lqy0rVdYkD/Mu+lso958lf
YY5mMFmUJpRfrqxbMsaozktPa+mW0tsFU2Advbnev3eX7+FyCfZ7HuLU26Z/3RbHqz78/7XdBf5v
DAtn9IDFCpA3ajmiJcXc6qsv3VIbP3ZqSeJIaEkhx2Kw5ymSfXXMvsz4s8Ft9U4AUWO3XeYPsKEe
4C+3Hrv1a4k4+L1DeI8PEdT1eCo0gwoA9WQZvxH/R52a6ZU42AJ/R6UeMS2ZS9jSTnuXtxAjrlWv
Cz1ofNpTvY0YNK0okJ8Vt+Jqa+CV4x9+a7EHBHaxtMjKiAyc+JUbM0vsJt2pgmFNE81jOPmJeS2N
svVUdzxMzBz8X4bvHjmf5QI7BBRUMd4ysw5hkY9JYfzBj2nmBhJ4sHiYtq981jrod4AD9CGB0/Vo
wZaCG5wNDNlewg0qoMYsJAnZtjhAnFOXc/rqwIBy7piJoKUY0zMIZiKH5eIm/ld7MlK7TX3lQYhs
g5HY0ka2+LFnHxtHOG047mAWEWCbsDVtXV5jeO3pb7PjmUNdiR/+69/jCTkGP/+xaewqqhL7vzdu
lgS1BAKo9RPwsSRPxmGQrOnMi7abX6snJbRBNQYUJpK7l2g7WTiWewy3I3jT9q3fFEUlIzGaTXrE
aESAR8qNcTsWUWvq5MZYcON01oqsT6VKy8BHtlJU+eI5z4i3VlvwiJWtrk2A/lyxcc8bc8QIBqlj
X7a+4ozCgRJAof3hsC9XbZYtcDIPLs8Pj/HAq7Ya73opyIgfSYsY/kHvIVYzvxxOXysX3NGYALwG
2qoViVjpWE07eUYrxbqYgyV4/tTwXmJYBe03Ykw7iibCI+3cktqMBLV9J9gTsAMK2joLWm1xmnbK
jplWx+vw+CfBoIqPYwGfbrYA5SdSn7fUNGPbtB/82zeV+G1OuzImsdbsRS40fkR6kGL0mj+PKtW0
NBUXpZe7q/EO9PGpoxyccekrvTIFM/vjIC6e50YH4M6swNsiDJBPF5M/xmb/BjJEatTswUOf/6Ug
1qv+OEIG9h0w8eWmQrnWL+nXyiyn4QYbotnaWq0aXOOPBiVWUS+J3FN7dqPZoXJhD1Qz1a/NRTVs
BRjiZWdSPhxirNacJYAjOkZAUxIEpAxHuSA27XQA6z8Zelz/6JL7+YmnsWbEvUU/ml9MbADhrAaH
IQTmfF8O8Jmy68SuOXUTeZsu202enbB6N3OjS9+xZZP4oTrVTZSaBnhZgFmstmSFlGUEleMs4EW0
9VxowSHnoowQXqVrkInoNozGcddfy4B4RH6VmBvIyXLGlLRda0cCDNTUSJh7RfaURohW5NUDNVz1
5TPbW66CPcGh8KCykFTUS7M4/OkeJqux9yVGXg4cf0BG5n+nmeFTf+KnMhpmXsu0Y5TGp7hw1/3c
/3mPIDWUEAU3Lmh0eruxJMRSPcy9Okp4GqOJKijUUU2e6/iGLfMGKTGR9Lf5wxb4LS2TguKWl97R
41wumXTPgSTHz6APHXzcvKczvImARgllmd8uX6wR0eZDlLLBhhjrHTyVOKxKeeuDEJ4oF/JP6Znu
Guw+XCRa1TfkSXKkzpBzWXzkddBKh7jCrc734/JYg6U0vVZZP4FMdxmXJbyxdXks/krggyNB07mW
jPIWI11PyeHSeaJ45Z2FNBp2xgJSsPWYWATykZgVfKx1csxoGzf+g5hdHOBcfMlWSXAWjBapOHvh
sZpUdIBhGy08NK+s47Catb4hVxOlIMxqRzut2y62Klt164buDmf92+G71xG6u95ET+38KaKpYyvp
0s8gc/2aYncd7ER1pzXOObHXP6mo1oFWy5Ay75DrsFMCFcsCucxHaIoFdlLJX0wYJD2FmaZTP+XB
Ilsbv1A4PwZF6lArK5jPvgt+jIKoNJYRb+oPp3Fh9FMT6CoOOgl05AoFVCKG+WhC1VdKMHobN1Vi
BIBeX2OW3eltKgPeEWA5OJUKpBvnq20ZgtY52XKo3on5UXTUpCm/BKvec172H4ovz3NpegNZ2Z6P
PN6vhuvk2T7wGZZRnuSw6smCgf8l9YHxlyuiHWUVIGeiKyeM3Fj5nantn0rqcU3AZqe1+seqGYks
A+gMfTIpmemnJ8xpB76Ww0TKME8JOlA8LAzxDRrtvGL5/vfJ57+gWLSsYRZGtuTwyIlbQZDbMwC/
sIzeT5axKakxPFHZrH3m+4y5wgkAbNTBZy9fTTg2MieG5h1WYwah8WVDBII0qHgrtYLNKqxSQDXU
0yXzkb3iVva0gwXCdFrcFjW2aRee6yPTENrDO6pXjCYsOGDrkylwnGrSjg9G0HVL3THoMXI7HIIR
8ZVHJuEr4cBBFwIZKzqvx4ajGIXP6Xpdv0aVSy0qr1Oag8qte8ZDLyQWVLZdtErr8ntT+NEznCEX
dZLVAbhPnRA6Z691RmHN6memsefbKpNgTJhNZ997or6VU2VN2uCeh4G58joUek7XzRliUi47s5fJ
puJpriOCEzxG8bPLyByh1IWppKVAkuPHOUfl0NOiT42siOTpzGiu+ihzSZfWTR6FoMJJKIAO34Zn
oXL18tNuiNxR2SZweFD9vSCHEz8rL+bYDqiXvpsWV9qfFVKwM/yFBPj2166jAI3DFdZGdLOW1bmp
QFzGWPaFI66orHagsG2tLphJFnB6AyVEL9Wk4gDEDj3euv07e7BVO3C8j91LhjZBf2fNswB+Fo/B
htQpef8aDVUQdeSu9rlYhymfUEkjyUWMJOt+KQZuLM2ZUF1AJnBDZ90gCnHkMdEEG+s5HNKdS0w2
dBuPB7P0LuGyV51rZaAfMogA7ODVTzKLUD8PCR9pbXQqkXjHBWVt/5/Zs7wf3J5VutOnKhmLSaSU
8JsFywQzvsYRH6Oi9uKB79NfKl6xi828GsMvVEj4QKz/7pFvqukXyJzIPhYBjtLDAMYsY9dFMK84
dDbVvB4U/zjO+BFvp+LfnMoZiN/yoR5gmfko3Psy22FhRyvn8+8oFuaFc+MCkBLsl8rnfW7ocSPD
zwJl6XyjgVrBExpXwu/AkU/XP92wTaKq5z2Mp6ZH/QB/LhGYvIq8dEML4KL4r5PcFscEtDELzsoc
TnmFbTghVRktCL2/1G96qk3nyq+XScQUve5Rl0pNcOl+gbv/jGF5TZzojlYpblXukQeJ4RLQEzaM
etwvCgudtSxr3oUWMZiGsO+s47qDj8WzLDfibx7GpN1LRH8ZeasGGcfP8jPHtCWqRajcH+47P0FG
OftNLhKsnIt5LACZaNiPtpSNVAnV8GWtzBk+XrliX8KBZtMV1jLlDsHCWhCQWIYeew7ZKi6JkRXC
6JxTegG9yIU33zYZ9giOJBL2oMpM7+q+BEmrDnbFOyT4S1g9FZbHjz68nUnXmf9X/I6b+y6eW8LA
pnl03swxnGJFchURyap9LPA1fkNBVP4zTKSMNdE2wszBVLBTjS+uwrIyi4uBq9d4YKUAxdlGOHUA
voYFN5idMr/osL00O3YFbtR0YjveksnCVYFLuKfsAQAiPSVmpgnZNUQSDGJ4MDblqlC6J6WXYywk
AFwWIsNQ2mp3JvDmTKdfgutixcT2B4NhaccF79nudTFpuTOiJvQ9WYmHdvh72+J6U0KRpXRGWPWk
TsbddVc3LlnsRk7tcj8DWVmzGDG/gZ/smqoXAQ6EumLKgvSuFYgfOC1YqG6IhEZ96r78iWj4On/G
UCOOgpl33rv0iNhaOiJ4PA3eY/DxMdYsqp9x4gxU06ZGCTa67Wo2IYv3dwmTn62r/kIoqthp3kii
DeUA2a5t/mSkbUp9XESViK38KMuGYMTkwGyMJpUamrzVeGB4JPyIPPcH20kwhKerzuOYGLrshPTe
x4glQ89Tf27WYRt5uO/YwEwYm1ne4d0xC1JpRJmluWCpXJtxMBmVq9D977+v5AwOQckRrWVVcGun
06RAK8XLjb2gQgTLKMuoEbXsNDnFVwvv0QDNIoGhy8gxC1fGYmrXxCIWkXRE04MAKtlixjSVN5+1
4FLdwOeVPTiNgLLb+MuoRiVdl8UQPnxRc7KRFXge1miU8hqtB1adVr3XZTpV8nMzA/eSyeoq9aAP
YEdGNGZEXjJnHxZ6AoR4FlSCm9iit2h5ySIwxeUEkZ/iL3jS9CQKEvzp4JkYGFdaKboDTerZ0N0z
sB35kdrdaNGEDc1/ipFv7tZNGTO2Xu4XmmWNQeEVmeepmFbkgyoUpMw59GNidkBcK65ZTlaqXWIL
wzhuXoret6hI3Jg6ZxCRB9jddY0a7lJQV8A8ugAe7Hsf5iOlvItI6QirxtljONckvRgUaWRf10qU
leUJiV9KPv6V9SX9W4SK+tdsIh7wz+mPKiCWV5XKcHgUBHdr3tNyJfa5EZIhpRB2FVAmJRW5tUdQ
DGFRowBQFOD4UCytHXBlXedAXJWpyRhIV+uzQsXe4whDHaNCSGMyqyMM/wyEl2MhpU1MB8bjes66
kKO57KJyLMzvxPS9tRP/y17ley+yusH8yrLKs/OMct06Rb08IZFgdLCyjpyux1hVA5fd4tyN/ZPN
a5+t9RIEsl8julsl4CKBWIF9Y+NvpsI8lEfy7V7tmtBCYNqfPnCHtJJyQZPTVV/FqsRlsq16LXFq
q3mdwAhbOp4dioiem1q2VVpRpwb5mjOuNzh1bRalWyB8nvHbcUkMJr9czH8tOmxTP6fjSAj8sNbW
UDdVlHsbLCEQuH48KN+B2dUsu7VHGSWcgggeyzpizqOcM/5BGanBvhIR6JJk+/RLH9YcBbZ9ijG+
v+AMh9YSQVROZmcKrJQQvwhahtyvUh2eLgpflMFf9e3jbIrhJ6IOKlTFn7WqT8mXIPJzd6gJ/OJk
khVjJLdr9RunesoLf4lixYXrSvP3LuXdAH+NBzNc2RR/Vbo9BugqpF8hNJ0/0jybvJiD4h1LSwae
PN1LGNk17h5h7M1lIWfHrkMLtuAiedy0q5RWH9iHMUow9Gp+4H+VCaIBYZHcMpSKgWaoDXtNKNhD
hmPI9exjR+yqKDWsgKPBBIl/h1XcJAIVxufB7z4OmAJydnDbYUE5bewyJqGYW/66DYDHgVBEZHVz
qqOO4hq8wkYWblaJy0NSPi9TKj3yK3fAkVJU1MYcwRGcNxNdknQWq2nflFL5W0K/YwThLQv99cv/
Ib4wTlyrbv9ypW81MkICPnPBC813CeVT5Vj+SYtPakNekU3IxEO8IIZEnDoryJnagfeIfnfHHSjb
yYX4O7B4vtfZcyeEjaLfugwzUCOic2EtHM6YY2+IJBYnr7PFEEWhEXoX2hWYCu6aff1OgAAbs3R0
pA+kRmWvt8rGieW6tCKUGaGPpzndMXJXeK978lh4Fw2kQ6sEImnJQo01ERclX376qinnC6LeIHsN
IUXNp/y2NJWoWfGBYiay6+yGiKLgOcXW5MS6JAbbpgHAGf0lg1V4ynfIxep6rqdNjtTX9lgwpa3y
+gkgIBrCkPuIW03uawzTJWqFDnlfQJHqKEkkI148MF5uMRqA4dBXjD7ELGeTBF1fK5IpzrpQ8RDv
Hz2/aau441d7VcHJzs1KSf6KKPCB1h0yLUiH6t1rHdsxKXkMPS0bwZIkwNsCoCYHDegZdtzf3GRD
AWvpO6A9mAkNYo7sl5impOwSiNHPuwkDPGdLT9cS+Q0j1VNMFYAndd/jNaohFUgNliYYDDWwgmsd
fs4vOqg/3S68xmyf5HYgaeYMuaabTz0ykjULOqJaDQ/o9E2mStTr4thRcI5/F9TBw0pmst3wIDja
305U89KQJf2bCfol5yulTb6T0w1R8a9KVnfuK4VTWjjsTYDtYzDwgGhHYb9JB2JnGxZNNmubN6TJ
rd5mAzJnBneJHn5w1eWoWY9zUD54qu4xMa2EPjz51HnKAOWLobkyC1QLXp5dvxFYt7W8LIXzXswx
PkF6Ob65QMtquRibcAWiwDtG+soohl9fL1lmNbsgWhQlf6V4C2B+fsHnlVGCYt9IIsI3NlgI5JuR
dhmjV6uWQBZtqFoyl8IcaGj6GQ8NxuEbeRSTiqDQq1S5T56KVM7cKimn7tH9UiNCev9qGIjc/cJG
C0i+md+y+bqnTdV7A2LQJ/8i2aRwD7DNPnGFVnT83gMDBz0blZ60qqQJEvjGXdzWapioXcdH9ayh
R71rI0zspJ5kJdomtBJEjIW/3bGuZCWkKykPY6rX1nTEnb2bbNQdVXx/ZmnXl/bICsI9/TJ4qMuV
QE8SL5NhzHjBJeh6DXxxtki7h+yxWagIA816+2uhOy2DYytEblpa8gFvLCKF/NHRmNpi2nqT8Rms
9aaGLl/+0i0pdZ7ob0tgWWz3XzI6k+UU0MKznIrlucvRVqYJaC8/8A+1cXm8/xAYjfynD++wxsmy
OWT+nD7PZu4oNaalpJ6Gq62aZoYxo51l4aIntKwmXXtkm1tsZ/qftR4WPYfH0Rb/hRfCHPFpcNYN
SzEu9vyF3oawRVyj72tRDtCjXLGC9e8bgfn+pQp0qhDRsjbwLcV0Fndknow/nODhzAQgUVC2awJR
eTTCu1QXrw6455Qn2Nht95pGkVTQSqKr9GyuuxxtJDrzug6RzcbWT1GbXPsnih+3EXomWlH21nnp
/krWhRVOLbChf5s3NcFoqd3lCUe8gBfnj8LXulExM6N2k0AuRd6Ado1i7otJ8xKk2RKDqGB7+j78
LN2XphpoNlmcMJn28saMtzuQgFeeKA0BwGQgn6H54FX1yM1pSaBMq8C9OEXIZm8l3o6j/S5u2fEb
4rNAo1Xr+kug3r2ODPYbr/8HzFgCgAntwhNXX52bkKRoG8V4KmZ2pEg8fgp5fVvCKezUUB7/PFu2
C2C/uT32jsNRVijkE0DgC4Wg+YxEt6l7xW7jtNv4dr0a/YZNpJroBTUnoUPb2zFHLlcuxnTueg2H
ZwWb3GBddz4ZXQZKPhqOEBv6Gz12fLonBG/15fPHFGoukF95WVuBz40p2TopSWoDlOHv/IJ6X0V1
j54lnNCNx+huiV9PJxZv5v7jIRev1WdgzLPruC6VG8yznfozu7sx/A1W1ZxMftFViIimdWRWY939
555mM3nrL2Eon/EPz5cwClY9GEa/lQD033cXiTczI1GvUU7jwIk3s7RyA6ihEbyvxpAJAOyy1qLQ
HsMlVekYbXYd1ooMrHK5h+tGAm0AcIxyJWoXAchb2GCquasGo5aHQRD15Ph+BlDDGGEMKS9UIF2d
S/1xy39Tjj1TImW4G/Y/460U77U1d4fguYJhqfNJuWhZ8Ha7pGgEaJ3vD4OrfEMtHsinoGgURbjV
/+FqAxGLT4RkOI1pK7h8q4nbkGPviC7GcGKSDy2KxwQBpV4QsOHRHmtyOFy/OJM2xOs4FdVwhpeT
PcV1bc8V0O9gY8aHR7+ZN1BBaQAZLA7HEbjulQUmOq28M5Zwp5W+3qTxwEFYZBqQAPx3D3Pvouei
SsR+VJDjoVu3BtOQfkrcwg4KnBzwKvTiIhaHxkC03/44Z4PILDCdSL5UjddgyZbb1RFZVdouAt/7
NHcl5vbi2/8jsEcVbTBzs32tfoBdO17UGYLPxk+6F5DLV+IUxilo6EXGaddj4UADPt/uLK9dV15Q
n8HhFNEFY2JwrvrtqEisE6d/32h9SP/WP6ttZp3NSoPeEdK1Mm0d1Xh5WLqpxnAjfuglzLPAC5ps
hc+lqh2cA9D4fShzayEE1b+lp6cQp9NwvhoV4H/c1n0SdUiP+GfJe1YIIodXeAecTUE36N6sn7tZ
XLNGKcmlUhix+1BA2Qn3HWlDE4H5HvHIM4q8CBCvxyjhvBORZEmqosSXdGoqAOD5HKBezopw9leH
stZMR9AIPywqOCO68/XuIMXnQEn1DGYgpvCosuo2MPXlrFuJ8r6u7vg08RaYr47N1buhz8wSifv2
Jd1Crc3M9RZJ98dhcHb+ZA6DnrHoXLl27Z3Rx3LjHT5q1yXb5HWpPHEltxqnW97DKTTnpfDdvddn
xTulnHG3dAC/zEekIWnyNFjKX04OlSnAnz8lTd0YJGhGAtiw+7oVAg/lxm0/ooXUN9c0rNUcV0aa
8aZWL+a7XITc78+NOXjTgcoc12QC7zszZvMvN/DSc+aOsC2uPLtvFDJhZZXPhH4V72UcE9FIih1Z
fEyYTHcoUWX2+gkSXKYgQvcSlVzOLAVmikBVS8ZGOkujn6ELIVHg1P4VN6RIHXDGjc1Wg8H6pYHu
la3zlZp3h47UzhUKaMQujCuM5JcXNAAnRlq/cdecvvT1cr9jfLy21r75x4KEHYCOxRlmOf4/+dj3
mqZ58Fg+x/A+NBvouf2x3QhrsvkpwrXAzHLv49CLOt8t9Gsw1y7Xr3gQPZKdZLMfXkH7wBp+FjrJ
41PngsNxBC0p3O+sbrFZZgxMTeKnAyWSzRw1O9FU0tR8FhPkp7lwEFNkt7flP9W8bVrEVu/I8aHL
MSqwXZrYOZua82Pmnr0ikbehSEFGFY3ssJebvjw99yj/OJx4uqpNL4tx8gvAw7PbnvDP0C1H2dtl
v73l8wGiJ7XO9SgJ1LAuCwhYzQZM7fr8Glq+7BykhWJvRPB+B8xP9vF4TYTnGg2klIZ5AmlYNMH4
8WY2FQoMq1MoLs4dRNaXvpj44tPoDBM/I+q6mAwBhpXlA5qVaXrzbi/7XtjqBEQP3R5/vSaLUkcG
Us2UEqWOsyfmkri93eIvoOODznjwRsQUzp/O7VBG5yBacCbH23snf95GrMeR4DMBrZrIFgGi7j3D
H6GT+4jKPoNt3R5YE+6qwiZtemvoaqrsSQvKOLAY8M++cJbko8/7aS/aE1TiigWDNd74GYPMQ8TD
Y+/YY1QAXhUhUmO+EdWqlkNulvupoNrBY4TcauXguQplc0NUVshrr6CfkNIV1sMH9MBo23Us5N+W
0+4yQkjjOaJPcaAAHTZcz3uqi9LLj3z5Rf5Ol9XsxSc5283a/PjKvUZEsjtK9aAoLoxNuEYstpTO
CCAt1ggd4gd9FcVpPHunkMLzvIhWqvIK+dr3Z1NC5H4ao3Fb7/qFY/ccm25AMJjovsyDyqY0bB2x
34qplA9mc8StdnbHyJSO4TmutqaL4YfjTIsGh/rFPfbpCbc1fBoKiIf1RfXO5IN16XhTZJsS/ams
2NphbDMZU8G5mljJdv5sldncEeegjXKNpf0KXSm5/oa0YlXygO1pnBtxJg9bmU0pl4c0CK2vAzjv
crjCEPGR208QBB0lYIdc99JFpd2ZFt24p+SRZ/YPxLpVL4sfeFR7gYsILDFFcY5QJ0LWfnbhedfE
b5KQG1LxfWqKR0SXi+0gckffStUw3u9Pbb3iv9jpPMswgl6FUxLAjH4T2s9pZ0VPRLqoM2fWzNf7
0ZGhrXVrbxDUiA+lEaMCh8mtNygyOzYFIV2qBgMRfe6I+SWd+9DkV/5kpCPRL72zedQID2f/mxZj
20eq8FERRZr81CwUIcIKiobYJMGIL/45SvsTdw39t1AirsBmbMKX5YvaHADtPH+4erE+Wt/0+uNb
LYZW6rV7YAQutsl7fr5XZdsV6Y9fJKLJLdJCbkrtTCI1Xy4bvF6mPsXcPLYLS29d/xAc0Yrz9m9t
UcabWTh/Wj/dtxkKcDQhRfVCQCOnx4AvSkiZlmXChFtKun5nYXEc23JZeas7N4hTb5W9uFGtgZhV
rGYw6BbVJbgpcAbwGZOq64XonN7igd2yDrPz6JFGP3UZfnjRNhIE0WGM4Iqb6g5p9YfM7so8kxyw
iFPN9Y+BPJZ6/h5rdCEDXV8ECWKAxRr4fiJ2fRkyz/23dOfsKFAR5Hs3NbU/fAHjEEDMBoPCGOV7
izsAxAri+xUEGzqTeXF/TpBBRGywpUMG/GLLUp18AU31fdoLeKGxlLNb6i5WvYEYJY89m+Dkccrh
d9DRfaIZvhCggyAR6Moq0Ubobyq9/OcaSN3j5z9dm++lhCv2OF35ZpgywYq+7cfNkVmNSdt6IAvI
erRSeqVGqpvCeRcX0NOHTOUnVxKqTD2422I+f6NzHoeMkTugZGalFvX/kDd1tiyR8/p4ff1lIlvI
j5ap9c6ATiMuoXBagynUcBl8qqMPiSD1jSCAFmi7mxfCaX3ifdc/XPMHjZF7fB5i0iYhD7UB6Ztj
ZbD5LVp/ShSn3OK4LZPxfH+8vN5gsk7v5ZOlVtFRtbGrRxtAVdSYRtwiWNM8EHsh9m/EKe555XHG
9M+n0sS1e/cd60KZw4kGo3H7JN/bbWevCwaCE54QC7T5iO/OgSVnNbfRH0G5q6/LfPWrfvBpFBVG
1Clv9QsEB/eEWxoEMVuVk1+11ivTUeaunoFQAUZGcpP8x/h3Emz5mwtWHoIcNFyWokgikbD9uKPU
L5VaW+BNWhXcNt24Zt54cVieQuK78izykqwpACWop7BQkgWZdpMRdjbJaEx0MKuGhpQXefwi7pnn
MVMIpGEh03oKOBMlLreMr4I7vJH0zapztneVEiz8CjUES2XkTWZ4eOY1mzjPzap4Ar5km4ARG7Ah
GIEKh5+oOlfR0qDyzzG9U4SW5YlUeymI7YnM7uLtN3zLCN7otHLGXhOgqcKo+H54aHxJIkNG1tWy
dZ0q31gEu35PzF/XjIldE+q5/0kDhuj2fmSDnmX9O9yRYzADbNw4T5G8ILOD1Ys5pyDI05VPjNKw
UAER66xTPqitAEqayQqAUREXkPztDXod3SbyY70oy61s2+7E6VoI7azZLWoxMMo0NTAukMkaTEPK
RxBLjxJKjEhH7si4Vxrfax8dtEdTqDmLTmOgfgfoPU5ekGZinBHxo7b0xuKEa7nmsSndsrXvgO48
H4ONobRSM6zi0h9QbN2+2PKk+Kqe0p1YdCZtiSKh9efsmqf0gqXNEWrCL6hmhWLlPbUtmcBB/HrQ
177tN1zUiIq0PVIT9zKqKcpKfCyvDOj6XQnZVaCf4rlJPUWBlDtg/ZER3GPa0yTwuachmJmFDmer
wv7ow9Pj3DxR3awmjUAtrRXoF7Zdt/1amx81/WzrerjcBLfNVflfWeQFVE72S2x61Ql9i4xUYtmL
RtfMkAKls4pxFLHk+4DNuL3FnQI80JlPqvQDNIYPhR3xf/ci7pZaoxdp7+FCkaO+ZihSrkq7KNyE
NxLjFaCw7MRV/xH3loM1JdJE3pEWPln+t2LJqRe7Ed9fhmDBZ8hqY1QG3Wasa/Uwo/ZHwLXtp7uE
7b+5MTUUy4BsT6+fDzdI/uSzuxE4zePK/dzR3kNHRICzy+k4zBcApCWbqe8eHSS3JhBAe1R1yAMB
sICVZU2oq7QL8pSz120i8o1P0HUjIkpz6Lbdq2D3I1H0M9xwek5/SvFUURwR/vUQDE5wxH+oNCSD
zQcgqzAex4l8DWjZHtQzxgmjUCYbyGTHukoEJKfT2FUK8sCYuZNkSsImRaXkw0UwdSKLkbgXh0Yi
AGFeSuBRvcxLOVgMlefunho1h5Wyr8qdkfdAtT3STmdVM1mW0E5xHP/BPFDzJIuaODYgRuwe/e0i
QgH3cE4dxwh++HucWmXarMRIJKugMX5hCm4y048GFuh5qb/1ZGX4pis5y1e3XyZ6lfaHH3MvGGyG
rF7Fxdf9+qO6d+y65jlmcFh6xsDFhQ0qsBqIZ+xlkmKHJg3UZS/p9HyMP4fLQopnQf6g9VRgvThC
DrQ/6H7qeaKPl9k4lgJb6l6PaoQDIMf4Qtw0YNwFHs5djO+GXMGCoN1qUI3KtQ+xDtz0DVOAC/Dr
cWrZVCNbOHhgTa/ogQ9AB2L92NsDvR75npgOZevswFyjBMWHT8L54mmteuiy21hF6E46xFX+34u+
lYGqZEIsITJYEejcW1M2fPLTvdufz94XL+wovHcyAnaryI2nBzbNUt8lsJe3iWx1/xnxjqvZkOkc
Eo1psk3I7QZbmlyvUKJ8QKnf9tQWMM7HopUSxMOlPVRJEZBd23LTjMe+U1UeUk3abwpTuThxij24
xA066IUkJ1mcxgM5bPJ27mP51UQl9NU9Vg6QdvYjkkORv51KnCe+us+5yhtD+seZ0WV1VWhPhhNc
SOl47NGeh5sW1UImLdPSV0UsCBR+rJr5geeBD/PpB2uj9WmSTvGtRKLw93w2JlEqTC6P8a3vUoTq
BYBWuC9AwWo2MKrAoSst7WuSYwHrfv3BVEXXf5nGO1wAowNcdKom2C9LRIBTYamebAwm/mUU3sFM
oS0k1swAyq5cqqkF0ATm2fCYKpHOvYcj1In5gIh5wcItnVOtLUh7HfdiL3ZUbdmFEYEvbyFJCzlj
gtq4Bazv3KJ4D9uEEOgvdE+3740h/mOUXUoCVH+ZEtZa8lf+7l+nPpsG+rI8gJKeJlcGF53b0Bgp
PQYsNbIxORQYkhG3+zCV18aZBvKbTvBZLxkDO3s55qh7lSMIR9hIu0oQ1KoxSEb/DnrVhZLSYB1h
GEWhG96STnbg46uzebdLSu3HtNRea0KsfZ4bLCfkkJ8X/dWvyf74NE/eSNL50XMqWySXuFN2Mike
H9ydUOO7AQUOfdcn3/61tfc+uS4OoYmrrBFixCNoQ5QJ0pS7za5TQ62Bss+NcS52oFv6FqJnN5em
qCRQdJa27rw1j28DyyxXwZGCXmssd0WlEFf9HBF+86gQPjbF8v5sH77M0qPB8G55Vj6OP3Si/OFK
RCnh0KdlbSechhqQtvltJVBTtAmqB08Qy8N+GfKw1UefTx9JaqEV6xyZFavb8U9ISIAxuDkHffY2
G6qHS+bvUBpeUKT+OcfFj29X0uU8hlk7oEYugC4/DlBd2wmZfXCTkUqwJz7WyLye+vG0gTuecoid
ZMHQdRG3VNLs2HktXZUBnlX9XyH1n4v8rSGRzR81rOYjloqZZwo/vafXKErPyBDm/lgwSWiIkEod
f1p3FpO6870qTwecIAXeFuzuyX6X7bDZojvbYJPGXI6LAzcwKcWDVIxmUHwC2OLy1zmGsT/09sqY
7WF5QHpvBDqjVpvQmSbiN1mVH4FF5c3Rpudu+KsfUscYbrSJ4DvS/qK7ZI4Ehs9rrxSFJr/eNgGd
PNhb3Lar0XLqbU6YX84+SeNQJZPYoFP8QKNftTPknT7vdqQqrhyO4lFfTcyKfNkYIK8lpssN0me5
+p0Do6BZgPuVzsvVtQCUxTt2eGu74wDSKRjgHuOFfDnuJMveHuj1MZpFlTOkADmWPjrr9Lb2hB9U
QbID9VSfbVSqjORAWsYKgQg8/4YDyIiL8JlfLclZMbWk36hqSxPrtk+GEdsEmj3M33+b2i4/Myuk
qOHe1wUXendMZOtmmBRsXbHWeZiVuK8Q9LF82F+k0i16kBVb4shpQekcITjNFjQwEPsNAUmYlvca
QHC277kbzc+YjT7+KpKIaSh3qtyjAqg9ucDFcTVfEM6TCn0pAJSE1EelPrAA57D/8/ia3wtO77n4
yNxB0mqAZXJpPIjmn/WAYfBAwVlr9lgYiF4oJo8mZuSMateDFjw5b0bSsEQcdE/DsG1dmaHQOCeJ
VeZZvcLTvi2AnNwlh8Bgdz5YSO5Tf6PZIMr92cDG5lBoAVhc+imZQU5pTTEf98MI8IbHNNtc/64d
FEA73fTMUbG2l+M5eZaBmaKHMkByGlDLJSCKDaJ4psoEZJUalujRY/PE29B5ILnKWci575YYoLK5
hIkDwForCOOFAKpwZUMkbTTgam1s/CkOSvIl+KOjwjV+SdJ9RJZ9SFDJOlI10OuGk07s2vx9pmTr
9Vo4AQlvvZWSa8Sb7SHkHP+S3NuiqWwqr9Y+E2VZV3Z8bUEyWNo9M0RpGyhuzEHXWaXIebuYFk7g
ly5bTWzlMuNV3B+dkAKJOleQM+fY9x/8WpukG4Z2nDNPQhMvixHPzQXGWGjIlatQjw6F0R/APX1M
CZqpOrS8Ki5gBfDrYzPZuwrDh5QvGuw0hxGwvSMqSdV/YkZBBVpIwueCY1imDMFDXeYgiZ+/eVBu
nsSVz3k4o7/4SIoN55k0SRkoZUkAi4uAS8cZEC+BNDTRb7nsuv0v1TRJqTvOoJamONri0GZT/PPs
2zK9GiC1dpdH8OS4E2FDhUMvFhm40PDGcbuyQuXKAStTH9Op19KwxllaButy10Zw35CoHnUSdcRK
AYqJTH+GxeB4x2f3XLFdN40PCEFBnXs+a+oYUAyXRa6zoflf4ZAGJOM09NiYeHKetPamjitO9dUX
UjY0ekRz2vkGqheaVQLuQi3K7DMY6s+wCqkceIJKs6KhwXKd7WilD/Ji8AD/PBk9d0CC4Goc/CK1
WlxxKhZjmgWuW+/lM+n8JOyuhVZ+M6ivv7FtMg1H17bZkBp7E70Mpc91qEzGCMJmkzXdqNLgIuCS
vHUKHgoR4e2pm5Pj4M4/tMzLNCFb74QAUfz9ctkEAlWwPzOPB1bNvaw+/m/9Wg4oWQ0Zl5rOmgHA
VyTbqgmEESho3oozQ4TsE8TaT9E7KE9T86n5d0pg7zdKHFDXjxkr0qoy9d+bnlYoAvElyTvNX7tf
dHcpw1byiLzvHT5E6NLKqbnEOe8QWEhbZSCItmBIJE3TAW5K+SPzQxonO00jX0qKb4CXD7uBAlap
NNwumuvpLMOLhx7jzIVs6VMrOJfR7d2v+Gmep1JiRv8mK957/ptl2g9VeSl4AmWGXsdPVJXj1Gtm
x1ws7SLvstM8bi0H9HSttuFRTQEskbXWcsHC/fRPazReMwXTdMh68GIrwc25PDcb5+LQTkmMVx2M
91HMcSZw7h6CpcZ+BdcaZbt8ba37mjp8DsuY8zvQmbxNsjNwyL++qNeg2C5EoNsu6tbhOklTAVfZ
+qjsOeVyKySQiuJa+W3M75CvVl4TEoRYVY7g7FyFfJGZUGo4ys3k4bQtPhNLEe7Q/ppol3jupNOp
SptLha4rmhMiYe3Lw/8Ike3GdWFT9yFJ4tHqNDgzJdZ2IhcP5tgeubJy3XVhIbbGRjE+8VKPNwOx
QjYHFwv/GA2uMTcd60w+eqGrbdqP74LzGonpmrR7Kx5XG/4xeyq1oW618eE4yCGH3sFWgJo67gPb
bF11OQhm/CtLDwYEtuYndZRZABDhWM0Y+IppbOkCes8lxip6lah4AS7SwwMQ4b1b7v53mXHTo2Wz
2jzotK44nogJG+a7SoSFZ9XXC5Qi2HHQw3wMwHGSD97ZmWfteJwjBo34usUmokbUQ5weeCvF5DhR
RRHs9upLXgLhKTTZNBrO1dNq7mujwgzkLxCUNGu5r7CsPQLjyuUS++cgtxFZY/xAEhxv3JQkcrnd
CQOXm+Gbz6S8G2T5XzKmUSC0wyEBzoGk95FYbMCh9WJPRIx3jnqehA6xvxqa+5lGUl43JCfDmYaG
vfSRkK0qZxEsPzzK/vBt4A7gCd8eLpyvAWcI7u7VlNj1O8K/v1QHwu6E/sZPy0gg79YsdmtwVKdJ
DMjeC9SuRSVYzCvSkO6t+RfrnCkBGA1Rvl0907yHB399sJZ7v+9++qEwhfiwJKYADmVIxgQFxSN2
wXEKKqfvGpDnlJ33+U6EUDNZtJigXr1MaM+DcFbPy6dD6Zw7Wz9UFMXIP91v938fp5/hWxquA2YV
QlLPmLTJ465Mv4qMccA3PCio+fHhW1PTr7zgi8qTChd0wGzm3kkhXZ3MmQ2rYebCYjXph5FXYAN7
hgDP7LlMhXyzUXaGLUKKs469/Swf+cyGwJrCT3s2egoURaQCWF38hh2gI4oRKsk8QGhq9n4OjSBg
aVro4Il7PQvmWJAamlwoDUe9asiJZSqaAHJ/hYMfIgmuV0zOowqctBbqBgCp4RMK7Gc9edFfrffF
gb8MvK0z/kGGbas6OadzxAqzqHrKE/2yogjuuu6bSnrMcv9GYVpjJmEYLfLnlQVvJLcbj16H8L4Z
GFRXb+f0lrKvi7vQkKmaghX5Er+UIgMnIz8JRayMhyWg/pPd1H9SZHJsT5zh/cVVicD4D7c15Uag
R2d2nrt2Iil/wVEUZoz6Yk0y2Gh9vTIrxHKHLtmSdx4Ld9j5G60JwY4tECQl3RfUcDTcUakPr+K/
eMKxubnNGVrsBuZWLcO5y2MQAEsUyMqcgIV9DJe5/2I1duGrSXeQVInSt/nJhCw+j0RTyaaRAP6i
ko4B8LvNLZbkxrxvkOWHJld7hmrhUbWVjCMh1wOTTx/xQWzTFVhw0SIrbZkhuIzbIJ40FQikYOVQ
fwMW95EgeeloT3D4YTCsFDHlekrkNA8mkGCa5gjm7c9wJrL8+ZdzDz5TOx9cZXcqEuZ8iSY4LmBZ
rz4dLCeNjOvd9x6zXHiejq2gjyKgAFahLRnlEe2aOR1pzSxrdVE3HdShD8lilmM0+LlvSz4TlvBY
8TFkzKT6UqiZZvGEmfAsr85rm2UUlxQyb1yb9WVbE41v9BKU/6aCuozKLEiOBJl+SYEGH6kQE52D
O4V1gImUYQARUwnMMih9A0BR6G1bjxAkJf1YXoVgQ/w5tyQaHrP1aLe0Nm/1LS6Zf35Bs8ovJRYj
OZEWuwU9+/D+oigbywfCB6o3GOZKLJoCbftZxBKhAmJ/FCN/RRCW77+rJLd6DxuCHK0T5kzK+dXi
YGAzqKzhgUeMooNsAq3f5If9NSRgI4lSpDs1YsIabJn0mJy7+QMBHl4jRUUTiw5iKhGNPBn7IwxA
bvJU/idY3PagxPC18o73V6wcac0YR681AAU3hxKBRZOIwD5BM1WGzDUiJgVcq2zAq+r55rg/KkC4
SYs74cFhgkvxzKCZjozsZKT47517RHmweHKeU3BdJiyaSrqOI8/cTLtCv+Bw5rMaeeSJew9jJxjt
d/xbEhmp4DYfX2CxMleR5YtNZchQYmD1hEg+9ImpO9K8QPhw4Z2gsUJ8N3tUEqxtuvhOg2W9wYZn
KjxrGc/ebfhfsuyuNYC2gLZSt2pIWe40PxUR52JeqyzUpcHZr4E0+2wGlWX4sSpkWhU075PdF1Dn
i9WGOd0bhA7nAYNT1PgPMPIuKS6vS5SMGV780krkxU4jS0JTYaLqpKO7DfCUFETt5CwH7jN7Ht92
qkp89KSkS/t4p85biu8TX1n9Hio0ya8J45X43zGBIb3cV+oMIz4QqV4K1dHB2JvyB69AECsdSWRK
jKVuOlT1syCjJcCX4p8snvtX26riT+R06NVtK1/On4jfP99CPXnLhkmC1F2DhpFpCjuu7r45amwO
UaETyyd2/6I9A20usqLSEl9T9u2gOEwyjNQsSf9olIPZ7l0GXPIMCjbHV77+QyjNbjsLvqA0+3Fu
UCVDr2R0HL0chA0fB9PUYPN8ParfgPABHOKrS6bimGia670dDOC3tmgb07Fkx59sjcSbiKleLJ/f
qRBBgTc/tja41uE6s5ytCv/p2qPO8S0/oKYPzDIpKSnL8zutT4wt4n4N3jrhelShFFJSyzrz2Cgb
Pd2uTZHGZ7AsSxMIUqE1oB4HxQoSRRYGLkR2JikoQpOyBQumgw1PDGtBUMppSPwAyt348VBNyyLs
hW/sMfaj4sW6bNgmsOrQfxJRaG9OfZ6Rn1OT5L6RkCeQ9rBj/S0WHZLyrdG+Y5Xln9v7Eqcf+mpk
aiya62u7GlYmEW24mFXrBInfustEPC8EHpPiVYR9Wha7zS0vYyv5JxBmXgBBUiYl1plnhl414XcC
GIzYtqukyf0g48Oxb10UFAywcLidM2/ZOjtg3M+b388EQNXA9iVE1DVNfWupcceMSyTDuiZnNcYE
7e42VMxTutoZLFoXT89eQSby2XqN2bCcA4GYUJbrinMy/sedh2hMhRsXXj7++GGxuJqqYZnHRxFZ
0+WQrAQfbC/5y1HfAHIbngrlQKyqAXFrchZ2LFlPSwc44FYb2FzvLe0up75/TMruj4CuEos67srQ
70BswCrE6mqFvp2xqEc9waIBKAk++bN1ge2UTPKMzAWH9+8FucDM8a5qpb9uayJ3RTjAbzQ8Twr7
xMMyQyqK3RyK63Zpk/8PTxwJJpKnZ24ACEN5Dd3Kk36zCSLtGmZhnS/1wxD14GuZVAU2zyVUafS0
WJkcqZo7b1kouF1ONZ9MOY7MDr061R0mphQj84Cq67IpX5hRUncSRbMiPkmvquHdLBkJlGYfSWoG
/Cex80lpJ2nBlD4EbA6Fp/SUm6RnhzF9hoozap75TDescPC7N3IKBqc5GznbCvuCaIDvXoZBxnuS
FzPSEf8moRQIKg+tox3cS0HmxFzVCodk+XwhI3nAJcoTMXE0yFGdEasTy3/kcW/6IejMVOWw4XP7
tehJmRPm1Y2genx75a3MxoZo1bGLYtxvolVoMb5cqzRqcQI6Atxi2vj0E44gQxRQTJDv/DHqPAw6
P9Qr+CRuHvRZVD0/d3NNdcwedhWalFB+4pnLam6uZAm65VKw3b+e8SMmKDFjx2tJKVSnxjLApML0
A0u55jc+pMgfV+ug1ltgdaQSXX3vyJcJFc241lMJ9zTgaaFNfBiLnmgIoMXLt7tUwgt1sKZAs1zY
sjVj7FiEL03R6SUePO6VHm7dnbtZYqohSVz0sZv97HL9VR2DEhnoY23WbWzh8QjSHwdT6+Kw/bsW
MclZNJPPKMjy09UrPrIh4GhdWs9t2va5Bo5fg9LYI3+7/Eiq2bSmiUG49kKbsbwOlOFv4JGOqY7I
KF9KBzLU84DqoipPz1rBYSFODzvSDYaH0Iy8NTPw7zmyjdItt+9qRtHYeo8a8VLD4gVh6NWwydMk
CKPUu7xpVlo09eTjmCpp917gvVge6dK3HiKJHlzLOVOXsCPuYK3aFyZ+1cOa0xj/Q1UkIaeoG2Rq
03MCORxoJrcmLy7hrpuXs4zJGBL2zqcxdxE3OM8BTipWcvCg9hpYa6px2GCLFdZVxX+JPCi+I1mZ
RI3CQN+44dBhSuLMvBbrDnPPsS/+897CKWPrs/iUwpCzJRRnqzmtK14cFpXNUc2J6M9AS0FSRRGi
EyzKgg74bBmu2/d3/HQOzoGjet0k+yagSTTC9QA5pJGHHW4Yy7uFUwcpAtBGKBkrDV8LB/UzHLCt
SSYDAtZPjEEUt+5tBtOTo5w6ocAQSnlWvI9ZbEtwqvLO7z0xs3jUzz+WrRi7du9gHXUMrIRoyHmr
HBylLJ/szhoN/S84Qh5TrtndTqzCjGvY1oPQNndiMqwb1Rmg8+9GbluB2+l4xOnAHja5sTNkceHw
IQ8UoNphdlhBd1iktjAh/9/FsSU6fZAVPY1Z3qy/zz2H0lz9pLferI175UKsGMwTHFoiHrdKvgdH
CMlIxTucBgWF5c3WuIoqscISHZPa5urHUeCdxJ6ZQmKCkopGXlF2phV0lM3F1/KU5dAUcdpZ0Que
FzNnklwpQkGcs8wJss2Zqdq00/VXCjBjlt3jTn2Zxo13q3cdYdYMr//ehwZVH467KxHaPAVKt2Wl
TkIRBZRtOs3imFCz4aS7o9hA8ZW8CEOjWIPaQiXTW9n/9JJfG6Fg/Jc9CsrHjmP8u2dlcq18ye9t
pTV0l4o4rFGtrtWpxiJNAES8CLzFnsVMo+Rmncbg8koHegtUC9LPda1D6Sesm3HALR82c91Kb4Mp
cI+ZlsT0v4bAympYvIwuFRTyHKpxcTBdR8P+JmDpSAQ7+kAfpv8GjEmCgLZ4JxL30wB7cethHLwk
tYdKp1fIMoq1cXXHqeDbR3zQv3E1DK/8QKbzKiynDBx+K2rkjgiOvfQbyCzE1MLBC6Xqqjv2EBxn
DGplso89I1j2XK/FuD2OB3jmxk0+guXOF5y3ZcUe/8RGa4FDQ1P82Vtr6pDIq2AKWCONnnCr9OzK
4gnTdyzodKH0ROXF0c04lL5PJHqZ1xcUlbWBac2Zt4kXYuNJmDTCevQu4iLPVx5pBejPWTcp+NkI
c1eKgLe+Earnhup4LfHu06wU2BQvN668p8XHY+87qMTqMChaNu7crmX0khceO9Q30kT8r5Kp7AxX
yc93HiutGeHU1hOtfSEhQAizzySP4/i3eJoM9W+8P1KnBqy3nmpj5S1t92Ov65UlMU9TLI6RdtF9
Y+TmrdEcZdbl/F+rN/9QUxq4C11ZoCXzWJAtnegfgZtIe+O3fzUkN9dZ0B35HSThK5IiSA+3ptUC
BMiaNdY5MqQx7evkJ2tWPMudL0etcHkGw63LlXPOdksHALkSwWmzpC82hKA5KGTDJW4uCawv/piI
xNaxrfKscZdSHq1YE8vOTSp2yFMnA1Pt17NcQ/3M1p4Mdd7Ffy+Mic5K4tB6R/U1ULmm3JJTAbh5
+GlE/qmow3DDO5+jj9YeTNRELU3/p2PAJX60lkhMG2VedlKKcM2bVdw3iHzIkwGf3imcoWVB1D4J
W3Fid2zaOQ4LM5P2n00IcRvjcHiVoY6PFZbBzOzgPQPaUOkmwoLNuOuuwCNIRsj5KZoYaI0mj33v
zVnTfzR8sWxiuoNPR7AzEkK2HqrMacKq0ZJmmmvcg0bJ6FZ1ulhuzwCD6zLi6GRP0c108G2HVkc8
+oiboz3yFwnWCZItT5C8UKxVapGkfQ9rXw4Vq/EaqMvvcF7NzLVVrFzkp6pwX7gKGNsZ1ViI1fe+
AokwXd4GXo3sIOZFkZPXfU2ulB+6VdPW2k1djxWO6u7YLcZZCYdbt/gtqbE4G6i5pWIMtQYR2sde
OgwtDw4k8CCDdNt/z5szgb/5GmIW9F+wjQwGlwMfjdJ/+KConaIo7uNiX8D2oFHtbU/57CS7C1ES
p36cC+uxA9lVHH7aK45QUYOtICA7V5mZvj+FTSbNIJZomZuCQmyU4stu41rwTVuwg/OGbdVXjfjs
AnfZwBagn+MWzB/nqju4nvSGsL3SGdwNLuDVmK3TPRxtku12BoE4IwBlN5J4A14IMZZeny/PETZY
fACqt9HROilun5i39d6ne4LKZdP953yYnS3C2wb2m20W8le2YsBuyjM292NaEWJdgyjgEsby1Dc2
G+OKjFBXjGnFcFw9jzf8Eqo4fuMp/Gb55Mx18Hdm6haNTn1uDdh4Y7rnXNxF1Wf395XX+3kMvdoS
a3ROMvuIiRt81C74lYHj50+RseuCl+8AADCgENVZhgiWrEsnHRch0TplrR0GoRoApthM5besz9qW
L/wjPMkIzEk3DDHgyY6O/NwHPwJILeppMgzSBhtzPiIgEudtpip3QN7lzLBINuWQ35zppw+/KfSZ
uprdxTdUnB7vtdps6Wj4ey0NYbHzCz+DcOler79fTaOPqUTwc+lXt5zhOEqY4+8rkv0+OEJ9O2Pb
It+NRbQRW81agQ2eI5KH+SDmdkfDsqlbIOWCAisf4XT0qfz/7dIuABRnKqrLoxLHUfJFI2yMbUql
iInjKJOg87dWh9JZ9xpqfg3fnWrrNZKCdWWuD96lk5v4QGnxxudZU2hGKr8KpnNA7oleAcsHcSH9
c2og6LMTM35n6yxl9csDZahrcPQKBhio244bZnoEJWVpP2oko/L4iX02Z8Pwv0rdB5Er4vOGwbYO
rZP8tN7MNxXxFRz1p8QKnsbwIYne+RGCk323rlMzLWxCBI7oLErhOIfYm6jaeACTq9hduS9OEYHz
R/KOmz6xcindFRRbzBQ0xrUznHyQHAe3MiggxrBnRqQkJjYiW81RZN31Jq4gA7YURouS/JW7w3jP
IEzIG3inkgzbfd0nZ1vfm/oIuIhoSS4Tsty99EzcWTKlL7vZSVOzcl5Dkh9L6ODGHdEMhVy8qijV
M6ELfiiyAsb9KKYXyBin/GdlIao17kkrZA22xvYX1QM+mIO375V8ngpLq/4dBb0ABMik/fzWQXgG
HCpjMVknePZzrxFB/gw7GwuwMe9vaZm0Mhhku0lDTEcbO+xhw330ntH+w8sY9mmkvUsLZgzjJrJm
Lw3GliUkGOYD9qQDFxNYABP2NriIXvNiNqDBVpaTWQHqsgPAAMbyRVZ0cC3KhMrVKEIL7ogZuFpH
jBREfmv/rCKaPx7OpAiptELT33mXnpCib5bjGDRde7vooII4xQwW6j8/qqbpZveJF6jgH89UEViv
mbx59qadEOdSlpnrqOWgnIbvy/vwSBdNLtd5tzvN6Hjwe48pbF+AEtvb7Jo8b708wQl3mQ1BR5qn
2kAI+5B5JDbQzdTOhYwWSbuySpdUl4XzNg2w7min9ZrouYUQpiTwHqSbDYJsvlKRWFQStEXT6AsN
2gLul3so8H+6mGYifiBkFJMLMdoZG63e7yL3iipXQ+WzTgTSv1tBdGHe85RQMTSeyeJvmpJCjl6i
PopRFoEAB1MrrjXdNF+MFVjjqFFzJczUK1o0cZZGpzdvYvWo5Mby+SU3mfwG6Knx7nI5bN+XDcM1
e00a5aiOkDiRr4EjVrNCEJsKk9vnqxgShH+AxfHT/SzTuK051uNe3ts/mucPrxgb2kCvLs4/d3uz
5OiBHvdE23sBa1Zf26vRIiQaW1llXiEvwXe9yMCQJUOeLv+PD33HGV8/m950OPPrMomC9K7L0ayS
UO8qN88JliUKQsAljKRXBoWioCKgYXM6ykZ9VlQKOWZh2RZUZKnefJzTbob5LoCRysk/VqYbwl8z
KwmkJNk207A9bpG5IzqQwuwAnoO0xVY3asWzEHD4hvF5xkIlblKBq2RyUs3LVCS13qFf9lgoDXcj
Ta47RtMXG1ykfKljWpmjGdvGc2nufl25/MlggiLtLJlUU1JnBegJVSFZwemlld8u4TrzzRgNWuzM
I0mqz2xQiMwMnU7I2qj1IdgSnQsQa7oHDz4bO7g6aI88mQsW2U8glCDxioA/60/eET9q5DxZW5xs
EBtJ3OqQIt0tnw3FemFpYhY2JD7UuEEfeLTLSRpuGy/h66njrwW6wEdZsDnJ2HkgoBaD/VjlkX18
CYX1eH446K5Y2blam8AftQxaxH1mmUzaJDQyyZ7MgFrfSZ1mh0b3NjMx5zjjdi0tjC4fviA8Iiyd
r5mEiU8gVpl+bbPtS6mBAPKct02rjpNfULWjGl/fICIHqA8fF1l0vlRRJQmngEAcZ7MNf8TdFLsT
iVPLNXjV4Qui6WskMnroMEuC8JUkXO8ylMaNO9tUVf414OfGl23Craaezq/qXUDv6NtSsHuh/KAY
G/vGdbabzPPNj46ba7fiXysp31bw3aV5X8vUJAmCDrnrCgYLL9xKw0VlhV2r9P4jo6pd5AOnOzby
81wD/sMJdlUpTaH7A+L+4pbNCOOgQE82b2iIXrxcF1lavg3MEW6qXZtoCpBaclZ2lj+EmfSRjfZG
/GvrqQMQ+e16Jqn4j8z/oJYjgjKYTBt5l7o5MjPZAiA0raCDeyBn3uC8t4bGZPo6c/5/dCDFQZO1
xWWnDfGBz+xjpHt9tCytNf7jVK/Vv9EUp9WWQ7t0tzNSH5HVfoZ+3JMndXmDt/9ZExVtdVEpOr6k
vDLXyt9k4clTGffePwYRyU6ipBeYom3jdTCD98hWjt8uRUTOyFDkbT2pDh1OV1SMmlKm8Oqy+ixA
fATvdweMukoWTQdP8fV9TH25Flsradj4DdLeX4j7QVCNupPo4wgEwn+ZhMJQnS/SyO2u2GHo6bfE
QPT2/0aA12uIY3QK9FkVX1u0Qhx4CJ0xMZ2gi6Aqa1CQxhoGLJWBQhLut4d+JUAYjNhwEOh8ARhQ
TsOJBgK8t9r9D/ha0NZ0noEmdRs68sth06Bm8Y2xONTgSt04XtyHkBuU8XGx0aPLHNCR8+9I9vzB
ZwGd5Y+C8vUSJ811Mi15Svx4FkNvV7bx69c5whxWUjgLvxcUw3zWmdDziX/CA6A+3EWFQdfW7duM
O7O9dvUMB1id2EswnFimKfyFrqWxUPKwjoPawveG4JkIo36dIj89b64DvpooDfnZ0M/OBqdUKq6C
XCyMyTThpkgmgllkQsaUNAstNwg9NMDEIOd6Qt1d2p1bACURnzz2GhUApvqRIWiwLW4UKH0CHsu9
1WuErxfJMaHhgzSocrMhyoaCQ93m00zYJQQwwuFs8PBmbXtZi2FX4mFzR810bR/D+Pzuo6afvI/6
dx6AOm4xizNE+MCUgT861Sp3yDokAXgCXgLXuGohoCghjVvhIHLWs+3j7MSVRCbqD9LZrdlcwNhz
GjBAP9rgQvE6OX9fT0u6KIN1zb95wSEpUCfSvQmHraZC2dhUfWs23NL+y5D158LczL/67dBkndXJ
lXa3z5uDDxkAGevQ+TLigDhbAmjx+kn4TbzWNJSxAedxkMTcbPDm9fHOrw3JuCJwlbc2ORiNjxGb
7Hz1SRX99mbIivv+kiKTstxKWjIwc9YNGzM/gtajn69npg5epDk79VUUOPWDqodToCn2/ZBHVNRB
e6XHEU8grVp8gZeaptgrB7DoE3IJer1AThiAVpvWT+lOq0IVqkljynkK4L//unJa7MBq9phkwKGE
Z5IYAEhhR241gPtdIZaoIxmQh4U6inAyzIxI9dnea8H9Ro1oyL0zILatD039Xf0mcnXm+uXSVB/r
Qd1dMmvpTyHRm0kzX5Fi1AAtBEwueW+GtjF8ETKVTqvsYhtkyahmWdEjF0ip6TaniE6janfclBKg
rF5cCx5w4VoT+cQ3UWu+vHIMC85DUOEhomZyJWqUiE6hbB/5P7+aMoeNCv+9QuFB2ZWMsc6/Y+fu
S+sNq2Ar1t/DW0HErmbvX2j2piXljzdDd44ebJ2QxkzMra0j1hVEuwPHDptLFN2sExs+W8q3YhfH
nd5ELqDvEcW5gvshU7TmzodiyFmc+NlrS7nm7e8O0RrhR56AROXJ5jYuFJWQl8HpKlyBMN+S10c4
AoNNjwJgMirotl6rPTOiE8DMnT4PlerutV1RjhajyuBTHELWlKHb/bTEmj07y0OOZD3i/XYA4IR+
bJDb+OGKcvmQ3cdes33X5yAThAOo2KKNuuj6T9/WIdMoUhKS/BMjX0QjP7VYJZbbxZro2ei2xBjE
IU1vomIEqItDa5kQbLXlJPWGCGz3kUJsqIV7OSVbFlyXImvdCCKg1jSANFgobtPIZSct8d1H+DLS
cO8T9ExfoUuEaAtlcooceMnAbOw7xbzrNV9hwQVPe87hQK3egYgy5QenOEb5s5D9ulQ7i18Tphq0
+ptiwht363W33wzfTn/V8jgVuvNfQ7ZW6vSuulQztlGNyFhXowZv7bGRzk8tejo/DkP0CmoQmCDl
aFeB5OB9OvGsnN6ULZoGZVTKOPawvvEsiUD88nYoOJxeSPwwUrs/ZTSmDaGxxarzzmOVDV5KM69z
62kbm3JPo8mK8m4Ir6N7QWXPQIzfMRpzTJaLN6/+wqqaSfPr4ASR+x4kIsfruPEm1ieGZYXz9LUU
qlGA1Q3uBOncvW0lSAIQAmv5qHQ+D4aTGDXKVczBioIdWbV6BYV+6xYiCtqKZvSqLLMEdTYgWYc+
umEmyp+OF/gkR+Jz2Utqf52hpn1A89tyzWJ1XPMnOUUiAcY7mdGx9DwjcT81JC6cGvlUmhpOrFR2
xd+4NYH1FkvW1FZeaD/+LSvvJAQlqFVjwgqpXFswG/UuY8q2BE2TNUHVvCm6+05ot42JXopbhrvh
JI9vzI6pEMFLfv9NFgYEVQZebxuTmm7t6nJlyuP6Vwhu7wIXWsnx0DxFaU40tO1cuHzfj4SOPMQi
e6gV6NHv6ulKmavULBbfRh6slqevi6q1FVnfJxRn0M/FoRJWXOEgqScAguuMTxa8OflMP7RDJqIl
Npw7B5S391wCtROHza7uGLyCC8SLfMplPtj1WR2I3yB776peuk8KEnuqf+fxQlTpgEjgqRfw3fwL
2wSD2Z+erttvhcdTcijqKcKSDOPj4DAet+9om6MC/QU7LxJCY0Q0SUYicWIplknkZ3nD4XUklI77
DDNqEBcT2xgObChET3J+WHFgxuKmGgNfbOloxDxhnrJJvgH5LktymjsDPuHtiB19nQFTK5UF9BAg
p+V9D2UwACURAZ2Xp2i5Xmkk9L7+AgZKhey2Wpx+XnwPlO0t/s0TIc1Bcmn4Q33/f9VwR3cM61fB
LyGMIjr4OiDD49QtBCYGiOqhdAoqUVTU1MwLKN+Kaa+JeLL9aT7bVVFyAsrU1qLQ1YHmu3RwT7VK
5ppvooFhIzRzfBLUGFz/5zx6cEP3R30+kY2weoDBq5DsLpvLr2e9Tgcn2FocrDDhbh54aPax6qj/
dAzR5QBbCNHn649VashG+noD7u6HQy8HbpiI564RC2l+KhsEbMRaT1Yk3zrrKh0IfaB4YCjdhFXv
cNREx1F3+MpQlRcfKAUnvC8F5lHXLFChPF0W2YkeYCbJT0Gv8JTmW2EuT5mInQKcwO1gMVnUf4C4
EFjYoyw4Me+3X8HCBgzaqQmoy1ymLcv7AnI43oZA1046c7vdbO8+StBPgXAPOxs0qmhdgR5q69B/
DcYG+UmmjzW0nqnxNKJMI2B2Jv4zzGULmaXiWp0uGX+YEzbIPjx4r2xQXWIVbWlZ7px5dY8kjJPb
4jJnwzfWYnLGicFeVV/dL1r0KbLJYTi+LB6ybvEGKnIuK34p/mKvXTB4hahkrFQPL9BLD84yq6c9
PoIw23d9DRgH3YkS14Axm52IrsaTshho9RQ8RhPZsvec4SYwp9YArXhPdyxLbZZX2nf9rd7eaeoe
Uv1LEjI42pN6qdHoA2Tf2xZIJZNpYwhSGhQ5wVevm/wB55NCanlON8sz47PcaA8rD7boTnSI01Y2
UtDqjVhbvIuOf4AMLOr9xRISknwu5aGBQy6InaRIc2oYMWhr6pwalbfxcpZEl6zwzUbae7gcQopg
zie162V/0jIUINwYw45LNANnl9Ey9ebwDpe1jbHKI2kTagHTB30llWEg6caL2n53U/jFGHgmm/Fz
VAgQokNAX9YQmhOiaqROqjacT8Ysiw3JMAoTFukz7eJMLLWhBte6vZTlFG+FCbYKLNW3yCXpJdlm
wFIb3hJx9lnx+GukY77y6SxK686YSMniyb0DCuL4wjlYCLjY9QfJ1BMxOOQ8ih1pkxn61NVWAS4D
NFy400+yDsEJweni0Yqq5pInuADO8Vr+JbISvqOKUigeKReMmmAe5CGuM8vKYP9hoAuPrgTep87I
BmawKkyTT3W/ZLgrsRm03BEFReQnsL763UWIMtTj9GMCPCZ1uSYH40LVvFh5GlFOjjjczghmlfoZ
2HIj8cr64lYn77ENjj0fg6dADfSUyiSFPN54j0YiXeh9nAXXkBYjqLS6HPIv4ENXJe+WeDYNh4Ja
uKfDDo+OS/02YtZW5TFloi7zyV7SoQ6CtrTqY06o96YQTtlnPd05rG5a3lt/Swd1khb3xXj8uOyw
dnUK2k/65eLO4VVNXFdIvIihcm/qdMc6NTvaoT4v+jrDpM4ETiyntj84XEuxtMiUi7tv/anGVG93
+4S4gvHJM81nPtG/sHW0uLh3+Lh1tpnQ7z3HuddmKbTMUCiNJPl3hdLQMhnRg4EyVHJy/HEtpgb4
M2U/57+j5GhuLA2iIy2vJWDbQBycuVPLAu51Pra6UFtX5GYojFZViPK0p6q8cR8xS8QzdIp2h6IV
188psy+rUX/s1M2Cn0oAqjSBO+OQJT1dpc0DRutnKBjWqdv7+nM+gw7DogQNONeOU8Jr8GAm+jey
4LXEEciILWY4v7RuDewdTs3v1yVA8UNCAdMjZe5lG5u6YTHOj9drwHFls6kU2tAsHV/mNtVp1kjL
7ILH0AGLFTwCYbH+lKm8AvM3sSYs+2MuuMJXdK06Dt8tH5LMek1eQbkCfAbR+/9J0pM7SzSVF4AL
CzXxV/X427n4+a2NjL3BgMF4CHDncr44KefRpPeK5lma14RdJDc823D2dmJtu6jTADvhRkA0+wFK
Yr87Tuo6Bz7lmhcCdP9qcI5dKiPdDMZmxNqn54WUBFdgNS8XsssBzovHnJIY5MetfE9Htl7x1JJA
LuH/457hHMWIX3WTzcBEnk/UbpfuroGgXXiYN1mRuWyRRLI3WZW3SmPthpZxpwv+jFYyaX3ahYC9
KfP3d4txtINcYbLUbXAjU5xjsGRO5/fJLPOo0rUWjOwYUAnIyZCIUKNng6cjVuhXr8dmNEyX7quZ
FSb0YulIEaO3SfLtMmEFG83roWYDGo7FLIF5WT559lv/FR2Ugu+4uyFIoxv6IQ910QYceW9Rjmrn
g5s81BOsSP9MVzBmbZ1RG4XKa6YEs/utB9jEMJrEz5VS0bwzNagVTIOxeDD6rB4eEnuScGJwXbHN
Lo2zXyyU/qGYEO8WCvra06PgkhcP2ns4wwMyM+j8k7HhSVolkbUbIv/eQHkvKrSwKpuYOA+KUOt1
DM6CNcKKKhso7BABUYUvCdLGmTzIA2WsfMGc/CMlrWJz/iehtl2/N9Ts6gubsuvPsZeR8qNhtGvu
dPgk4Mob12E7EC+yNBAzHhrKVL7BFDn+Mgc8Chjdu8mZ70YHxQTBJ2VxICQoUEPmEYS3eL7weO+b
QfUC+RsLbe3A6rRyc7uX/GLYV25lDWcaUWE4QAqw9LaEKsrqGno+VcboZX2aYJxnGjXW7lDgRsTa
boOKpt42piqXl4FwF/Z/4MPKNs7zL2sIjKVNbqyJMy2eqQuttouDTyRyMBt3qoP8ONJyETqiuP6p
HI+pewAOXmt3SaYsx/TjqkTNvUYLxGseQ7L23BRuQUvW1qdt/ltw7xb3tVxmh3JjUrMhhcQRCwD2
acqDb4+yZ61wZlLEJJzTHjJ1wIvEV065bqJl80pGGXNMg8OJ1KVAx2vppnMxAFFnuSfmaO7xW+wG
ymgvlrAxhn4tng0iV+dQPA3TUCmdz4WqzPUtIhG+1+fYMW2dO7ITRvd4a1ebKeVqB9im/kqw7TE9
T7rv7N5oP7vt8Z/qr0jxEedSbQosb+DnI4+YQEqzof5BBO9l9rRndS6iO+KfRXBqL6ERDd3qhnbX
+h1H+HQNR8DnNuLeR4Zokh/5p1WO1F9obIfbmBNIRey+l4x7DOogNO+XzLIOv+z5UslwHFOtk+vw
IJxBufRaeBWPWToWukeOw0ACF42mNpBakpTVhBev8zR10tohvQRptZDakq3Zrns5ZX+PBeHRjZjX
9lbnCo+XU3eSzYEOj26j3KwJEUpW/Vr9KVd+yQkFBkGpdmhSUNp8AvOhz43epQAlPaY8RRd5dTmS
BXTIwvxfWgzsMg54TF+kdLY+CE/n+e9Sjc3C+p6SAnU5YTRndZm7FMlMaSnam1kDQRM8x1/wD5uk
SoZf5K+xa0ZfiuD3m1iUMYRClKk4SHbBSD+eYb4r6jmHaq2ddQzr73wqokDBLCGjhEvdvQzB2rq+
2mtS8tB3dQA+KKHDL67x5FhZz5W6wPgkqZ6xK5m0DRn1tC5zrbQAU+YwzmeLMWMi/pyuqeYHffvu
uAl0G4ZQY9gd61ugC7GRLGNNaIO8CYeRRWSQ8nrpFV7/aZCECRtzJMkiX+TFGJJaqfujfDo4FR49
0UeI9PjhFQ67vDRHc8dyetNQi4KmDcDbc6V0kD7A+7JbhK80Z5YYTHcofTpk+/nMHy+WGwCRwfj9
W/R3ChS74CG+rOgxsNUbkPmF/6Iq/yNkNVoF4noL8nRtTN4GUIEKztO1rfRaL7U5GVq6A6kJkZsL
5RTK1Hhg5L53QcKfBXDD+5XOU1YfMJTQqfIt0AsaVTPcEnmx6w5iUPrVnUxSy4sqcdUQocJMKM6Z
AsxdZCIy6HV++5EHF5CtBN6Kopx3At0GCjqNzQZN4apImxEZtXz4DMILKPR5chOodkEWFexRkIAR
dmWxgiG6hASz0kq8xKgFW19S4mGv3SklpeV6DpFbZK5lTFOf+olazT6ZW9ujkBDD85B4nNJz4XRR
T15Rzdh9ROckVBNDjvSyTIZVeZuKpB2m0WknUmBAt8DejeUNiQzn+Rx7eWnZno2LgSYtC6ZpKk+A
Tr+KNsOfZjuGR0wLzOZVpJGU4WTKljRrTucfcsb3nv87MxPz5d+NDICwQn27Ntq9uOeC3K+QoZpF
9lrTzf9rDF2pt1xxXE4zX/2NbtU07VsbfP3kGYs9Gy77QOwSMfr+Xq3oFeV8LE9+0xlkYijgGZ5S
1y3574EqTiAvlOMAxD37yjZeMlNmcFfqFa4HjpuMmvEJkDw52/smc9MIG9S1vvvVe8CleCWqK4OG
btFqGv3KhoaQyfO/aDC7RJYv3WIdsGACBEBOzq9VOLQzJWShDABmEQCypXIUr8UnFlPUm8xF9R0R
96jFFf5YkQPU9mw4Dc0jdQS9TTl3kFDazPRCswQt8wK6UG8j8xGFWWqxBfikF4zlO/UIOnih54f4
43lK+m6XrHNVU/SiKWvps0u76ocm2MX4ZZYm0Sx0gOpEOFrro4Ldfnmjic3mrOFHZlOuNLThVQOI
/3iq8Y/bSBFDKQj2UVtNtKcKtJctpK34wAWC8DbszlDQvHN0XrB9hXZocTv1IvLNspIbsriUVGy7
BcbDNW3aUTlAdwO/Te7UPSnJmnIvsZbKQAthtkMPZb9Yb31Ckn5sR4iuYG5+pLu/TULqgC6pPXdZ
p6+EYOuShtxmqpz+qVhcwc0Pan70zYIigIaVSh0YnbHMhYbQ6BmAUI/wBLUmWk2cDPDwLyvXnUk0
9+xsyZXeKySfIepj2q2RuT960RslLyWwNiFTnbHF2ruHGy0x6gV0WLUqs6NEFIx4fNJ9eYvljDEn
iNQFoeMe88oZbUDpw1mLX/oL/aBbc4/oX201TPivaSFFE24TOzIXsUYm9WXRhBNBB2HElKsUj6Pg
NI3axJ4v6aFM6VrcqHC5IE04UQlCKp8aakJEqgAOvW++a4VyyDSe+2Odpv7jHfwvXGN6qto+Om6I
3mCVLnAXd+z8oHbzoyut7mED+SIqZGBAQZqm8znkKTPJr9sEG1TzfJCtvr8yy6uQ3aMm+bgurDjG
LsrSSUhazsF3/agRV4HwCxzfgBtGHZn2a09qhaqspswmEnyM9dLU4TktOzuoCCGQKBwo5wO9D7YH
mg7cXkC0HnGy4RA2gWeqJ/Q+WRj6ViYetxCFcxaU1cN7qj08KG5ntHbvq8mSrXlT16vH+pZVbA57
IlkOHtGWEXQCIQTdMjlSPbxuwhPDaC6BoEPyeh3pcOqloR3ONj8JsHEdwywtRS6QjEjrLHJEgCRr
B3dqqAl5OxR7dfGEe+QwGhM9gWk9HdzCUgDfzawzJcFcIfS5axwRtrXgJeotWulv5Xn378TFwwWC
4uW5z2w8kgxyvLxxdS7lcuE6GeUvT57aRKCxmgF3YErj1aakDJiH2NLzKznrlmVCTbakTusjncXB
21vKfnuwY9o284LGSE6V0pzTXnkegutYTBdKMuPhoNfBDAWuoaI1BqKGRf9T1wx5Lw4YpgAqkhLN
zcHw3Pi4AOfWV2yCcSR6EHb3/wNT/OLpW2RLc+WU7D5hRz+m6hkvNqs7P+9yCi+oE3jY4id67Mv/
NhMDOskzW6rBXlS5lUtkLeo3MuRI8qme7o2911V5Db1BdhVo4J2aPYRMSmoBpjgS/Yo6vLvmS2v3
C5awSYiO1P1Z3EAmiKSmiPTcbO0AjFEj0077cI+5rKYr+V89W20ebwbrx7cNVnecFQ0kWm5ByMUp
CfYd5yjpF7iryrfNzpIL4/QVeYowsJkBLem9g2JtoLEQuUMabheoLmbUYprn9ESRYELLCBz9IAyX
hSkLZh82NApNpNzGk+B6LGj/9JBDkxj7QO/TxvxaGWuuRGxKVC5noC0jg968lleMxLoIitSOpfbN
RB0AAkdFIyBhKHSRsGp+TIj0EXe6OOOUrRZK/aORuouu3dAOmoM09nrSvd6xmG0WaPkTSi/bVDkc
AFX7LtsxAzBoeURYH2hHkdNNdI1qpsAOSZV4RJFKwwPJmZRTLpVbeS4w7u1iyTLlleIlQaA+MvIJ
HIAf/13pxZAbwWxlIB2qHiVirgfbwc/GkKX0xbpPKVegIpMjIIl1BgHkS0E7DeMW0Y0sCMlMfs0p
sBZxGMF4X3B2Ic813nx1yHReV2G0S/M0U6xc2GLxTK4D90JK9MrDbE4aK4Jvxr2PMuqYDSonr+SN
WasyTMK1bhyKUVuGlAItsjTzOU6nEfqvu6UVd0y+oAboUp2Yopbkwj5OXJz0iS6iZqZn6Uluruzy
vH4uS8btzY4M6O/l+ki5Lb7046ZsSLrLhaPC0Zq+zTGJLnVb6E7xOsdusbZnCE1rJ6cacHYWz947
lxud7YBiN2OKgg+Cc61uKVXsAoZ/Ak0KocaFG/0FJhmwOR0spgNi1JAEOzRm9fIPZcU2ZqoUNO6Y
YIOjH529m/ZHEoMvAZkjo91PMypuWrAVF9AIeH+Clr77zANRjXJrS2uuqjQo5Cpe2fj4XMht+ikw
msKptaariR3IzMZm2/ptHnbOJ3TreWtpngvkwaKimh9qGdgPa0373+Wa0kJYNunPgcijR0fniKNS
SjGZjSxRnQ19Cq08gRigRbfntPjsyRHb6r2/jNYNK8Rhi7QQMngeuxZoIKfKKU6K3W+Wn5n7CCYL
yP5k6uRlJXGEQ8vmHryU9I89ia7RNAID2oosn1l8RaLGXm9JFj6U9jbYKcKI5MM0BmNJw9aAm4Jg
hnFnpkUX9HLl9sO2b8+GgeHzENjyGAPwfA/26XTeg/fEKOdr1HiZjbbv3NuPkqztAJqPqr1OXROO
huWveQ2Pzbijon42LXjqSRwOA5yXxoc4Q+WLVxhl73ZCtu8ihaXcWWx8boc+qQ/PbJrD0/qDRYCg
Y/ZR80B8SAfHVW5D3e/0uCzxh77xEQRbVfrZeyhIUTMo7o+5tMym6Sco4CPp57aRNPss55T9vio+
iw0L1Z6qHK7seIR4VXwd6mbTjg2xoXp07nvfgCk0jUAExG+MnlnJhKiBZdmb8DIIN2k0BOcWytAh
0bKsENLuCEFFzPswjNQYJOPvicWs5jPrIZUGZvh+oj5mX6HoOEVlRCYnEccVLAgOc8bFg/2oNVzQ
Bw9bxlaXOFX1jndpuQx0LhZLQG0GKJybL6RZLdEzLYJbBZeEgdBFPqFIsfR8BbKj67pRzyA37Ed/
N7WN+WQ/ZnW7oRLGdzjCKOhU21BCogNeIrrtqYbRUQhagGt0i9s0285iZwSy28W3h6PJ8C+xZcG+
DfZ3saRZz/Ttv3dEUdkB4n8dg4K5T9uEdW7/+q2rHRcj90j0hP/J52DqM0H8LCoMq9Kr4lnCuLkR
BzGzQ6UdercgPEHMBk8O++nHwlwZtLYdkrADQS3aQH0sglfnLeUdYSqaHXG4+ySM3N8qQUHp23RU
KzRmNYepxAV++n/SKbXC+rlfSR0wBeLsMZ1cMDUWJHc6jQiwrJPee0c2c/WZaxFQKBNdtTn2Eemv
JYdKjK1s2baVfOEJBCwkeQT1dRfDMf1KZukEiWLVsfA6owZ2flR3GGwA8DZluBkPtvx9rsgvBXJk
88y78GpAkKsXHIej80eSqCBFdXcUaNud/sE1iv95hI1j3fyiSiIvkBpoW2fW55Q6z98IDRMXmkQq
JDrz4zKik7cNlHkSIwlDicT39uuV40m9G23/xK+8JNAVMyIL41XayDPujQE33RI/hqH6kILz32pN
OaNIAp+AK1FxOi73iw04CpIJbW2+4JwQg7UHVwONwxY/LgsVA9Ygax/qegBdbpMtbCTY0QYgWaiZ
pXwkoL6YPYd83mNTApAz1FcmLknxo2cEngt2raMk8sGHuBOiZLJI0pDl5HuBL5dk5h60aw6jgy6r
IKjn+iv+nVDE64yFkGqs0Knispoq4V1gub9ujeJk9cLmRbvF/IHgQQh+5OEwbThPMlwQWb4hxlkv
MFf5VPISwecougUBn0J8X4nUijzB63ZgL9RlLZgWyjS0roTgJkP7QY94PBwNPTQqF6sGKxy6F+PN
ZnOXaeVwz4+77jDazWIg/rtnXYi5pRpFU8flIuG2BQndtgK7xEKJEUr1v4ulylmXs3LhJCxAebpH
+4h30hV78UQbgY0E0zEtt8GZlAYjPM4rVvWGDThMuWCfx51R5yLsdssWa+SThhBib4QYQd0q6dRH
KM7RA1nOypcPEekxuBsuDo0YDJSdYnkfKVVEqPYGxXXU4Hf5DuwM3xLHKRe1megOnCW6YyaLtIVc
hmpnSfLQPK5fEjiikjnLfoHWgAJMx315W7Rl3jAIk/av8XjSEWKs+XPIpbbAeLr9MlWKXyPF/KNV
4w4zBRUmzclI7pjd/53yex+8gVmtC4HEcVDPiXM5U7Iw324sQKqMDHJN/hT6IEf/gxALXlpLh57u
SI1J+ST3iywX85X7mw/FRx2Q+5x9VVZvfaUujh+y7Hd4iclr+nPRTJrtpeGh8lM04/s5vX/MYN7E
pHs3sDuiwj/xDSU0wTR65zLfdjKyCYswL2CA6tBFOwtqnstJSDwDxdpPWlwAOSqPDjJZDP02Y/nG
M2QK2KcJa8BMwVSc/jtyuSX9SQU5A+8R791W1DDRq4q9M4KeUkRhqhRmt7PFWKakZzTIpQX7JIJ7
f1T6P1t5H3j/nczLBkdk2N6aHiKlt2KDszOnt4Oj6VVv+8cB3CKxfZUAUm/U1+C6oagNHVM7Byjh
2JkVzSNLYOLSgQ/qcv1geeyz5vzghILLypgaObvS7PYwb1RKcFbJ64adgBkwIS4Sff6i12CMv1a2
toYThsiagsotT7QEwBUCLJY1K4ZpemaZ7GNdr/YJYdH0z1V819uRf4iHTUhVr0HB0pax0CPHG/fL
8wjK5Ja0tXPDCnAF4pJw4mifHPvr1I0WjVKLCKUrh5G0uGrHbnTQ/fmMyAZXYIEdJnjDDi/z2Oy4
LmyD1cs3nq1lD61mZfUOw8WQ5St5sJlBdJc6nAI5XRDYH+kcmr0Gyy2xIuTkehRmcFRWjIQELdSr
DJa0g996tGIXEWkFpqRnYgg1LhM9lgVqRDeSvQTK/gY9RYmuVJtI3tqW1WMYOYgvZnM+WLGyNB59
gaBMw4MQrHlM4Dx8J7rrxGYe3BvhvA4PgwZVmxFYacuE6laDd+DJ0cEX8xfoqe7vdQrK6F4zorvT
rTezEnirZs7OVadlURdPBXpTVcXdeWvrUD+1fBhXaeWpTXWsGBXhuOTnM65/xMic8R+vNVmHRpsp
DgdJzTk+eTFCgG5AhtWh9fOf7x8RqMwN9KaAUGF+r+X/1OsMCxRAyGwGaZQnNhr9QSGVSys9WU+f
uDWz5/SVmGV4cfY0rs7CG7HnTiAMtiX7uF6mtsAPqw3NXrGAvpgta989M2HkuLGQkfXYFM4Tswp/
CwLbkVorNC+fPVUIWw+iCBjDptIAJtqmzS0lPHP++ZY6gGkkWMVUM1RZqRpaQ92kc7ndSwpxKsE3
9RyvfFYno4LKHR7cgi1VhbGPIcAMAxln3jxCHJz952tVa9wRgWdncXfDW3M4c9EJ83nO33dLL0Wm
6JAIysI1/JvMX3VGowsiAlq8J1WtYu2XQP9nB6p0JdGiD/4VmXy8KbpRLS1q80HrviM/AF7IYo+W
MqIWMX29Irr2FTR1T84a0MuFhgbd7mcuRaPVI/OPlreMFt3zniR7WRGUOmvQnYpvTKkiluP01MRq
nV4D7fPy74vYSqB/xhLlS7NknPAFUCrC+Tnv7MH7cGjgxLtvOID6mBvnWkM+F84FzJ1q2oTlOSVh
8RBQMCL2UvoR3yuqrkRMOFT+bN1Wmz6axpqKnF48C5ORWR9lcF9KKWAM0TYIM51r4fI+LBLZNO9n
XBxw/75xG3ePZLb2lwgaSt2zN0g+VSACRmkPiwjBlTuCxg9juE5JR6UTkUpqS2CwNhb0+Ma8BHi5
rzEyWhoSiRKnFdmljBf5ru9K+2KIYuLNaiRVPOGQftjssCfgtYVSQENFwyQ0buzJvFMwrz5iknLa
39/gAHFaIgpMazRr6Vz81ng7DvOZzFVhTJgRKK7jMc0H0CfuuYLkap087kzQJJf/fFdZ8rB2muvD
nJGmRIiiXzVHzj/EYlvl1f4ybF241aOrlE0Ox/LuCeO94rvA0QNTO+CHtqa184d9sdYh1b9FXd/C
n+kR4CROnGJVI1nI8ZJvev+6RU3gGiMrzuorc9a2S2V1c1t7uZBryQ5VxPs12zOTJYh4NEVmIiuM
by7g4uT7j9No83yUwDSXk5wKIEQUK2rb1lepUKWCo9XlpEVoCi2jhfI7UwxD3kbk7WlzEuuLoUoo
mEdW9WPmF8vjIH1U8RuuwCW5EYzXrWrBKpWa7KyAL6YbtgAyTN8mHzWO3dgOwkzQjXL4rj8zY4uS
0AB+xyUmj9ghTaHetitDwatE5Uvqh+onJYWM9KfeYMM4ooyB7GUhsybF31SKiB72K8doyDao9T/0
TsBjwRkdyiqWGtwoeFeHfybk0Du8AvR0BaUoJZjJNoqYt6XVbqp9GvaJsI5sldkUjxF4oM1nuzZm
IiEowl/t2LSDjFbnhLKzRPM/VInNLnezNBd/7dwAHMV0E3JjrU1AeELedBhit7lwKXN3Cb3tLp6A
QZIJJ5qF4MQCxjZbJ2e5wDCwBpcMb96YykV+8LnmUj/vilZxvTMQTKntVm1tAFvFCk1RlgG6gD98
PuUS7qExNvctVceWxzSmK4+vvWASEeHNCdtDmlP8Os3Z350Zl00bpmL3XbE9xq/fZ8cmMohCm0Jd
4upXWcl70AH7nErHUBYBa+kOdiSf5FDm7J+C5rnQBQT0r+Hw/vVplFjnfWVlV4qlmshp2l2aYPZh
PFCagVS2ojUNZ9WQunLcjCvrj7gr9eUtJeMj7WZ27/A7k5Jn1t0HgX4pXAvkdsgmd++t1ZklxH3Y
0FYR3lBLSkXPJuiMUK7T3Bt3rlT9rWcrsKv7mkmcAkseYE6zJfuHaUNOHpiHzSzYvm04znNlUM9I
+ezcy7iRON/n8RCFajye7xNh/FtYk3Tp/yoUBZLRjBe/vw9lq7XqSzH0ZjFfWI6Zqae2TSSLdgT4
2ZfV25f1Jg7LQcjYLh/wpFdjr4DlQczWTGWWW3MEw09ISZBls193OiQ+gr+H11jdcetU/wpk36m/
kaF6cKnixabek2ASsYYFjXYYdcId8gea0+tpBH/XdPPKO+4DyVvfLqvpDeYfyCIae/5vo3KKJ59d
GYGFhNYe0ZrFOMyfn8IuktRF1m6U0XN6jbFbR3lI1d/9Dq6uPqc+6DgbUlcfh47bRvBr+l7hOh3I
ZEFAX5Ie8DA81i5tE/U+mhXJyAkenyMpiVroZDYrW4sC9tMvH08yIISyEvcm4DfC/qZbG6plRQDY
JYnpBCgnZ5BTSX6DSAdF9LfHh64NhoFpgOQMX+I0yXmT7ae9Mp1SPUSN3/aR5xfkfOyAhvYylQ0F
X1NQ1RhtGZdUAHfIRHYE2sJbW0nIbOjDTuZCozxRd1OhmbCWrE/BB+M5EYcHkAo9FXcYCmSKOSzD
X+DexKdLlKr2Q1isdJRYQgYeNKvYH5UB/i2Wu+FKpK5e2pDSvB4hnXQQWc8evD8Y1QXROmUAYZNy
9gpFnYP0YBA28hH/oaC7BoR67PBtOF7QStSZlMHrEk7g8iroc0A6YcOKiiKwBczuqX4yz3ON/5Yb
KlR/tKoNqMs78burgKOBsCUa37xldSLXCVvFPkNJ7XKB038CVdGzcXKSvUcDjMG1FRQmidqrvgz2
I62AoPv9EKlhJEE/PB+oVksG41H8ldfqVsbZmarNTyToUmhedQMd6GjIWzRTnAdP7v0J+HSX122H
6HnhFU0tlVDfifVICKxbTgCxkcYQxWjovAgLS2hQRmNNHLuYpu0u0+e2ih2JEvC+7ETMk5Mtd6hR
Q6nmTz8lQ8Qp8baDdUgwMQwqNKW4c9PUfnVryzMng0P/O4lIe+ual+5SDsae40wjG+vOUiqaini0
O+e7O7NeK7SDdzCFTkFPSWPMd4Qcl7FF0AeRQzTteUge9YUgZQMdv2qO2o1VA6isNk7qQ0thxV1g
hqAlBQ5C6yGTLIsG+l2BH4WvshKosI+1pnnOqYiF9ZrMWf1roWwKOq3ba2iDtjJUwwylruJMrKd4
C1L8JYiFCelvsV6C1Y7kaome9WukEdbZhu6/V5RU0aJ1uF2Hvjt2t0bVqsdazPQzm1hiqWzyn/so
Fz4xxGSxZwUq81I2TAHOYdaBdr0x0kD5H8CnYVt4TZf8lYhVhx6fM9Ncoby3mIijNaV9FFTbPWQP
GyZK2QyCZvBBAloIlLfRMJo1yDeaXxbUplRmJ3mMMuU3k2i73Ro1JM7Y/ErHCQi3sCYclEiqMmLa
kz7lOyf1izXheCbw4v79ff6IIyk3+702KUiHaEqif9AxLBq5getxHnMc2idWQ6A0//Moa1muq0QR
HZYbLoouk3UpYkcjW4cBLVLkdT63TrrGae3r7msHtwueyE/VeDeA430p2FyOg6gIzNrOcXMKL4Bl
Hlvih3hHhWBTDDQJZinhXUPf6qlWDk6tcbHeGNeeNPLf6IxVKTupcXWpV9d2erDSVPQI0Yc/AQO4
7ERsUEYJPqhEWl4ADE4ascyoi8gUk5tFa23r4Aq5NjClk7oJTtOJgmy56WgtE1v0zyGV7eg6RI3h
Ov+ETD+vjmvfC9b/fR7F45ot52PcjSZQGoB+MWK0Eu52x384nzm29OWf+Aqr3OyxVTuTh5zoHd/7
jeYmwKI3iIwmJ0hn6ozgx0+lKV+SJmcx5iNRKUTlEmvntpS80eH5x153B4S7uaLgTPpm/FFOf0o7
mNBrviLjrPnQcoF9xucq8J/m7hoVu4+s0cI4qpp4NF3/u2aSAab44DH5ALOaPVRW4Vp5oS3XXK7w
ZTy/gZD9pqSePJLPYts6Y6F9mv+JTpqVIFNaitEkCRiO0jukHBAeN5AsMmFi1qDOhuJhyCe2r4vU
BlzYaBVDhuqC6NK17cNGmuIBurhvGSnx49NilB9PhlKioZmC83WqHhMvuZaugzW/8rbajrw7M20E
qZ23S0lX3cCdduepT9MxBFwTT4fWTRKMpH5JCdGjSOpkAoyMmOekDxHtICeNsoi5gD8UY2Rmn2z5
IBBXoCs+VyJfAs6XJXvWfXkHJNvlb+4hYqgovopnPfHnTxwVmr3GqDM0qaq/C/ygBCvr1kgseH34
p3XH6pfB6eMEX7cHvXliHWzd72FuJ+/Ombvo7dA9Xbw/mC+LMYtYlm2PQajZrCdzWk6ixIS2JwTV
UIgv57+2eKP4aT0la5mT4eVHX1Xj2TjTMpEpycL0E+u/GMhEdBn9pLQUC8FzrLRhv/kr2vlIAsa9
6zSOPVZTYdGbBrDCZz3Q+BphTyfHHB/qitfqg2h0OqdLbmO/kh8TqNS7FxOnaPNbcbq3Wolo+293
xL+QA3Wq14L/vdV5Zj+ElxKAHp4C7lolHPJo/LRXkGY1VWfgJ21R9MyG5LExNgW1FADisagTHDb8
2v4Q4QNI0sg5XYTRzZ7Uj+w7zZNv7/vnzR0nwyMHVFugzuRdxrJLyZbPqcmtGFR+u4OMbw4DoVvx
MJoSVl+PudNp5R3VD9LIxU7DJwxYrkSJESsxIF6bK2l9xy6mrlsxZJu3O4GYnR4+u078e8blJIRw
keRClbcf66lDLpWEbDByeTiL5h0aF56Q2SuwqxSTbOriPRQvFSPtlT4lHPw096KIsJx+HMZEHI93
MN4ii2AWIw57oHY8srdAp4cyyoVlzKh9ID6e0uD5jp0pTR4VzaH0lZLy19qEoLBox+94wXddTFa/
u/2yvcvhg8QBbQ2XfhG5q/foZrQ+Fs+8FAx0H+/pCAwZV1wuxt1e5rZ2LPH1nFti6e8VsT7JIgfi
iByQ6eowVRPMJkeHIxxIdCsfKs9hunc7+fu+GcKIw2TQERNAmsmb+xLXN4OQmJq4A+ocJe16fgn8
l9RPr/eRspDBEDwMhEez2vx5b8dqFwZQSrMfAT5/7tg4ybDsV9X/SzQUFZi1CcQ/Nr8jrf3JbmO+
kacKwggn7kszQ2iexPHs6wQAsIjxbb7wzmUxD0xwWun1UuyWhco+BZS0Dy+HrhPG6DOsK6kAprdf
jsxz/DX0sJ6dHKaf9d/YnxGvK12RGrTxC7JUiwISG4soOubW14OaphEgyxCAHEVjk36jAvgN3e3X
eLxBd4DZQ5KrcC/KA1VCW3sIbrw+i4PZo9O213USVwdkKizpN49LCsyUZlscX3SlToJ9NFZwJ1s2
aSC8DZb8K//8dlCZLeYsGN8/5etLsuPmOfBH3A0hnX/2jWfgmvwElnmvBHKO0Ko14L3Le8nKF3fd
frxdHhzeMh1Op8BpoO3s9QIEdMlH6rxn1ouvk5C9EGb8PgfTPsXptCQ+lmEtbMAKkBt4wHRPjYtX
zjQ4ti5jzxvzz7dVtCq2IZiQnU8pKzlxzWYGytgsZxYCauq5zuF8lryoHDWEZsArnGyVu2tLE4UT
dQ90OTXwp+ojQZALDCR9lfBH6cb1TLx7n4iEnvXwA152qylUBndePw+BRfpCIWRUAXf2qaq53j/8
XBK8lcAvw6MqJ/q1Ajci5sedn1+9rU59bgSmmIKdBVpbrpKwf8dl60swVuiadcaQKYjGsyf5wohp
58MkRXD3ITOrQ0neNaq/We1Ei7p5KHNAFTCUKUOfUIEk6qU5r9rh6JDqpdjcQj4nUSOD5XMBUFUo
LcMI1Z7sATifhs/qD/DfkgwKT3g9xZ8Q5QkXDb3jj4EMAkRKwmCoMlhfM8VvWyksburA2gAyXEbj
2mGrcc76duJgfkAS857AF7nY7jhTV2y6FCnmtMs9f6doAR1OmFqkkEdV2wJyZHRmRWlCCDCFu183
7mzDg8WYx97zIM9qRYU9Qa6rwJrhE0X/0AJk3uYZK+9GEkG6XhTFw3Yg1liJ7/KmnCjkUwQKh1JO
xnzNvkUc0B6H2wxmdWI+tTsk1CQmUtthI1V+cj5lh8g6LrEiX27zgtpjXmF5LuJU6P1p2PR9P4Az
UwofJaVAcjzHVI3lrjGn6KUiIjWf5S/U0P2KYIG9T8HvsKzL630j6coA9eYbsKtfDLZWm3J3w2+c
8eivJhhGlrzMLV2nVKq5ZIZ6OJScL3nqxaOj67nZvD91C2uuY1WmppZSc9yktQTxpri4ndm8iU42
QS2cz7qXY+By3p8bX2zLXbz6rt5/EyyXLzTkOedyVJQojKrGlqnqxLRg236qGO+DZRGf4hhQR0l8
cNKLx02zdOtg6fysMlWYalaqeOzKbvTXEO3Np5Z87muL07LbdttiHFi4pufBp99pXHrDZyz1KubW
YfNgU2jS8+kINHu32xFoFVATM7JfUYmelC9N56U2ubwBazUFAM5/6dByctLqzX4I2APQBeqgK0V8
d+muvuo5fw64aZSpKteJ2hxnysC9vMxXQD5uX8s0c37iTIe9h8kd3RDrM6ub670x2QR7b48I0YSf
HTLWyJkju2un094dNcG9kABhjQjCW+NVGMR3kzxO1lk8dNqccb3cFAWhBIVfZ/du+SUcSvbqWpQq
9z9aO151Jwq9p2AvC/OJPOIDf/qW+4cv4At7B1nTXp+VsA7IY5iwfe4n1igS8Fabup7tawpe4V/q
HgtflH0DzrvYMI2aBfdAGgAFFW/1IBsB0eDbivg+DC5hvRQskfy1n9NDvuVU1W/8l5d3TBMzyqxs
TkEv/w059R7pYLAxQHMxoOwK23wQrK+0PRZWnqhir1fIMQTVqvaYJKr2B4lIOcuRKyKahd9xCd3U
HMObRwIBpqRZtNv/ihFwOD5obykXYYKiKTHovkT+l28apuK/24KH/DZfGyJgQvrpI7/Cb3A3ombH
BCQeVNLToNTdSz1R7+xBIiurAflpXdCJB/tYx2dgUoFY1YBiROI/1k6q+FUgT5aRWqE4k73Qt6uJ
PXovf7ccqy+jl/TQgFRu3g8d+i96HkKcfpIjyi7ywzi35kPEFzMfRSaT5ZmnSIBmdhHWAPURZk0T
0VndmyndddMrdBZwmAiBOmOqHVNNbDydQ5V+IoK469grhE9ywzCeWUhMzUcjSqXWCpcrPDC75aqk
fFWcRsGHVZeRLR4PXFmcZQ6hHlHhHsSP2E98ha89BnNb1+uSRNaecf5iqH/afk9hJQw/QWq3nALh
7HNo+DwMBibV5UwMVCzqZeDhQ4WfswkwBx/dmpeWpDXGFQmNG0ebaIvGHUNUlJpon8UpvrfZglFE
6y87Wob3kwKijDAOgAdSaazg0xhC4vMDBtUZNr2WK+z7Drd+1n76AlxibNAwchkxemEuPFNp5F3e
9sCL7xRMFQnMwAQDbWoi3CiRuWWnY/JLT9d0/lvTu37+ZqhEKEP4hDauF2e3MSwlK6jQnzaxAp9k
pC5iq2Q3DHy26gq5fmrah/+OXxMpihYfeDLzdATQ2HkiTOsm6bTw5JcOt4IeI9yqfkmkESdtmGfk
HrV27FDNEXlXMA9zqOAsvKU1q9kCp/U+YFBYlcDgyv+PmENY+PS5/FPiqkxTmsTO78XJZY09w8C/
7d+yZjRPVlbi/k6KV9/Z+N6Kc/IGuIYC8YR2MmZ51efCSnEgP0FqIaWZa8SxqVsRcP06PgIsjquQ
U3l8SED9PW7cJ6VVI+qrSyQiJZwTiE2PXLlTRRdHd9p1AVXHipPKEYBilaEs0JTTIH8oImrt9TBi
7jSIE0hIKXh+7AzX2wPC4D+6jXmIa6qy1/X5TZju+T958hniXwI1W72VVzBn+gkz2eqHxSgHWtLU
8zzQvV5Nz0vDuJhch253MmR3E50dxbnyUzbXch2cezcLMEilGsW1D2A7W7rSZu7XQVmk4e/DFSHw
VuLui/HAVVtZ63db5FVWrb/rP6tyCGnFwe7wz/W3l/vyQ7eWmKzrVkJFj6HAftKsK42dB1s97TGU
Z3sYhiFbHcd+T4k0/YwOJsxm9cGCOg9kNkeVvE9twnhRGxToZvfk2/M2edl9E+e4aC4xmINwrmOJ
7saVwD4DgZDu9X9/U1OyRldmuTiucRUHNaXmWwx7EGkW0pJX4NTcJvvfYIOHbyKJQcanoAr801aY
0N7Z21QEUpG+mcF/8BSX6WCKqyTUiPdKxnbit9gQThafTHIs62Gs2dA9o7Ua6huO+gn1uhqwKUw9
FWg1hFOkCu5EE7nBPhO0OUk2gmAyHmXkqPsaFyAKfegdDo+N17t7HzPs6wID+JE26+pMtI50xiZS
BX0SVapdoCgluY6XolzA1BNM7wKcQuL7vDyBykgvoxR4xoUFytgeIPNIKtKM67I2VLdrcWql04ZJ
1bG20owJ3mZ4dlXvAkI4trFqcTIu6mSDp4jKCx7lCMXSdEVNWQYTY9c7/kEEgrDFWopXPQ2LG+aO
Iuc8pA+iJtSimuQansf3GUrRerS+rQwc0quIW/0QKzEDIWeEJWqwIlyE4MFtRLoriAzxIrdLVSdQ
Ks7hDJKQ6QpNTlHTlDlAry+7yk91GD3CqYv9mqMIRYRUS3JFm/YKLZ4UzaDlZzvtrreZnBaDWwE7
v7hGQs5QVZuiQttd4CULFdDxbz5+LUJE8nX4TT8SXGJZJq203JlS4tXGLPGY0OB9asxUuag0f49h
R8+W/NdbXhYPWbr/4ByB1b54bFiQHbEfe6EUdZ6P1Bz3oTQ/3Oa5AAKjVxGcFAqgUIIQAIRyyVik
vxCKdVB8YOGJ2Jfs/oF7BJ3Ds2LfJowwimzJKFdIxUW+p6Zt0JWE1JUZINpsx4Gf/yR6BUuznCCK
PYkEk7uhu4+j8/KUTWCuIOwP0tBmAsxSrqX93wVnq5sSFtN7mFBhLRD0wnULzQBElfxJKr2Cu9z9
rwuI0F5BGQl0A91wv38YqBj1UxIgMLw32bR+pA2zo/4cftCbhxaHvvrkXCiD4pZbRk788w81t3Ol
Y8WuIzzjW0fEc62GcCQ0CVBPcc3SYz1T39y/6SbTkktdc+BlqzfYm4I9YTdW20SVqShdAHhBQO7T
vi5VaYzqGEllolOs2CUV+wpJgdoK8kdqBar65WuawauPCU4jwTgBjSzi0Eswmwp/jYsnGxNEmNjl
R6+o2e70rOZBYJZFiILvYHRqUCGlb6IHpAWt4XQu/YpYAKE8B356ocpQA354djS8sjCa5OAibK+f
Io4+cRg3iUN8xyVLNH6CpgiDxTXKr81kTgpyEdB/fJoC5gvoSV1g/alcsUQ2tBkaR5nU2IK0XBln
/Pe6S9+Z0jvvhysJJCgB0Hbol7njZZd7qljgEjZ1wv5Bh14neKn/zPhslPnN2a5B94zyr9YNZCvy
w/GDX2NTqE9yyMWbbbLven0Z35AQMpUCbqNg3jDvVDJEiKO7Hh6wwom9uvFVrlTBJpqb/ST/hdWG
Efn6YuiVNvALpwiddskG9ZkAB/aJIr0r5y83ilDr/5PDUOeQzRlTwg5qpByfTSHrSV0ZyK0SNo43
p8wVkOZW3kXeQ8u7ECGnfnPYT3UJrvOa3yKzAusgEP6X6p69iOuwnp/oaXedJTQgC6Y7uVAU81us
GGY8SuDiWKaw4o8BAQzVXiYrdwPHBb7BC9fZyXlk9Kc4xLgV6nYcuGuRwtHwbBkjal7v8c2+lsQS
3NquHmoHSh0pS01j3uUsbjnEOK4xwISc7nWHLeF3Cs/Rq6ltyPIuZr9Fc3ByTMH535Us7dcmzlQY
5lO3LOG0/WIb3Tr5j/QpZllTLLtbY907QibzhaSsSp6RFZfskJjnAldxBX/HpFCNQDVbsa2SASvd
nZOh0BnxSz4RFPxWyxSWlGM9ToahZmtsrKw+i9gVTbF60VpfpkiBwCBaKZa7PSKBhxmBHtA43jrZ
RdNqgaTLl0xMypFaiyg2OL+Cy43/TTe1MJIfjg6IxNXwYQvtS2WUVe8EvF3kofmn6lz6bw+SP6Bi
Gs92obr/EX1fXeHoLpGaSnSWNAv3o7nCdICEsFwIxcCRiYw2P+I4zHc4tJ6ndd+L82mx8Y9cmJ5N
7/Uc8lJhNe5Xmghqzff32kFy5BHKi/cfVEwLro2vCRfejGneyBTWyFuVLACBOIIWBYvjqb6LM6HT
EKk3XeInAY3dmzznDnzoIY83Iu9WDR8PlrwAdfyWuyEa0Y6rVznhlwXOZvD8dwoOczVEyJWemkv8
Zy2nLfSa4lTJr8SUCKcXD+6BMaqMTF9WXfESVuPt9ynXKwNzjYa+zsaIR9aJlYQc+UBPEeICzUy2
KXppXWIgwJ6czyNq+dUjOlXwaz+6mTLJ1Me/+bGmCnhLU5x9qb1LzoK5ADvZ0KP00uZ4rlPuIXH6
HmBnu+H4hcnTzeDfT8q9DGPKay+ZFDVrXqS6KkQIoM1fDyfonLCMkbj7jo31lHDJ3NMHD0+LLQg2
N7lnsgidjC6k7auBM4Xt/Dlye6/YI73+vwNYwqe2PNSDPpmIAwGoTVZVQG0O1sFDazTUBgoAq8f/
aBtC1ODoVKPGdJmktgoZ8TtkvhoxZgDEcKgNW+XgzzKTfZhXgXQUK9OxV0zntsHlVMqW7QW+DT87
0X5e2PYd5Zn4E5dsQM9sgWRWy1at5gemGABzzStAo1PXyH4ngdzmyO7WyopC0I//2MGiu1BrlGWZ
dzcr3w6dkVwMvdOiIHxF4vSXByLyDttMC/Mzfn4kb9TNc5zxtTDyUBYTOEJ+Mk6KUOLQsKyoTk2d
pC4F3ILSMjgwfIbuSj8Fm/tfRuUhZ3sAkOiiz2jhvj+S2Dx+j+VTkZEcdZiVi0Rp7pdwdjZolYuy
Gjrfh5Bs2tA5yTPaB5ROyZaP4EtejzhR8YBbK9R5SQLWFjDLW/0HipmyVHILE6eWTxWUYQMLWspI
QZJ7Mikj7Pv30K4YlEanfGUVOwWfkKhstJLBNlceljcs1MkHp1ZIEeMOWS2dlXk/WEJnodzgfksM
ftB42BBFH9NuIMx6sR4RG14wSewn130FwhaRWT7W6qeis53ktrloLNQWpGwBqlGw5UjHJzIxXuXY
U+RQUEihv/APprGNuMBzW0Zsh1Yk/HbuSTftDTVgFSvES0+JRJzQ1T20KQhCJ8s8FVhFruF9JnvB
QxFFCR4xpFBiNozRhI7Ay74R4vmV+S+Nc2kK7Vpq5NoHCh/FiImCXOBkStPYcNT18CGythx+fon3
YRrdfEvaKYVxfXDJXXC5XfHqUpeDTRAGgC2wi7lj76VKmEd2BADdMO+Ggs4OsTwqPW0D8crUVDnF
pJqSYdReEdOdk3kmIg1axwdGGQ0zUKWLBLrSZZjtBjrLkgeP8zmNbKilA6e33pZlmawQQh7NvFKG
wFshJzulXiwzkZistTcCqU08/z6JxoNtTNYMia5RJr3XeMWF6dc4eRdeoa+ZRG0EV29q/CKUfE4h
McEZa0tA/ppKyC/zGWNCEdGTCB/rkCQq55fTjsxJD25R5SVNrMwmJMGOu+g8Bita+4eDAnda+Cw0
ket7QwPfLv0j6QPkIgjskMimKGHQVQHIF+0vg6nFqsNy5GvQ4wIcQ8TwnrwXEMYqInX8k/3Yy5BX
udMzQ1zzgwf0INoJwwnQ7G7W33AFM9WBNH5WSe+VISlxfrbHEoEWtZfl338WDTNJ8BUw6hUuIZ/+
AyuoK3caczSOYWDgY5eP6+1FVgZp5evcFAKr6Q9KDYWI3l1wr/tzLG70wC1FG9bn7ANDpnQd1I6Q
SVBGGGtZZZV6HZso87cm0bF5rLnKyesnabFpeHVuorKVQB9COvR4+6UF7B6vpHJrhFMtJfhmgya7
uGiKBf2rpTl+YyZXjUopA0YEq4VcSzOUtmjSxPCR2rndv8PTuHFBCAfG7LxKaR+IvshiedCML7ft
u2LNFoMxjYitWBJlfSwBBtW5uBS6HE18a607V7KZtQnMiyVzyvYl231zwP1g/+YuY9skcWH9Taxz
ZxFktyy77BVnsQAMHs+s9ZUdqFQgOMIfow8XrkbnwRyhainoZCdA+gKW8dCak7xiv/qGsWvV/PLq
7cxX8MG0ga4U8qFfUFc65H6hYFsqlLuffRuvAnQrl4vHhgPsP+EyMZSKh5ASvBHbqh3yTBp7R/pI
RKNCRLv76hch5I3wSLTPD0mpNG87+JAZvO5/mhWCdxbi0AsUgCRjH0pbQ67rB0KvvOMdiwzMV4dd
d19FcW+ayscvIKXKGcsrNa5I/B5Ej8kqLmM7Q9gYMwPRWXNMEDawroYW9AJDBQbrQzz8i+KpeGU/
9YVQChoFM3vyy/pzNmpo3hzZLdsrXClxDE7YhTwN6b3DZXeAOsGUGndw3lNEXJxB9S97oWuZGpi7
PXdZzibtEZc0LbhJEK5bfQqqaqztMjRqWYCbu/LU3Eq1gRckeJB3pU8DvQj54LzRpvNm1Obc/Ok/
6W5gIlfI0nEzRR5YNW4WMC3CgqCKKOJP9xSpu7VSJYS1DzVhq7Ync+U7RNCpO2DNJLzsK7l4S8Lb
srcnMmeEVQNZhjUs83YI4xnoculQMhTUgUY399O/JtP0Box70AjCCTL/0NIIEgJC5Q18jhRZgQQX
ZjvGNnDqMEWHUwZ1R+z9Q+2pTfPXG3lYGf72+UPRKOmrTMRCDLfl+dvA7chXmeNdD6YAsvIkNWs/
G9CLhcLFBsfCCMDCgEWn3ofZzW3bzbq1sFzy7fFlpQqOpl8YPCd5yxFAxASICpIOzrtzrk6lUMtj
+bjOcDLX77nuZD7XoaCBnjN7nVGEA0hY5hL0/V74UqzRbkJkz+Rj7l5zal6Z722JnKHzKELzoFKJ
akSeA5TxrCYsUmg1Rx/rCh1dbJFo8SaP5+R5pp/glcpBm5cKGKbF0Lq2JJx14fNUb4e0RGsyiq+z
8jWlMd8/RLdIo3UIRd/9wQcH0xW2QnrOYL7XPIpIvaQHVPVroQR8yZFKlw1LU16RTdBbGD2i0vTw
DH3fhqFb2n6y+tXBSoSMdm9llDgJBApeEpH1PS7FAs2X7DPjuawHZmWaMbfBa8e37S1XuAGI+xvK
hZmffeNiRCWruX5T4KYCx7yBFQ39PleSffb9O0A2vCqll5Whva7NKPRG9U2qlqqE312Ut/hWhDSV
Axgmm4AvRw1grHL1uzgYQ8NHzmvMMPzFxk3Yx9WJU/ifVVA0hrFyzQM0pqhHGWa8XfCRsGgXVj94
SUrIM197BOQVut/1MIMRL2XMCu0RqUHF0NZdzS4UeZRU4q2UCzhCy7gdp0JjFQGgIz/jT+HkabPz
MtXxbaRHjhG1u0eoYynFYz3XcrKWlBp+aSiPsCecMVPCQKLpRbqseZ950SZVG5DAm4aqT9385egh
NFtAVp1Do9i6TP6HoIo6a3tVQ5l1S5CQnNA/gFdtvfT1G4usMLpKko/Zgnj0mxU/sAAK0+uZCFK4
rJH1CNd0RmbIju5J9HI0J8XcxgWVstC9Bz0uA0VeVtNm2BOuWshVmzzSipFx1SA+wtqXTv+FOlBP
3pc89Mmu4d1f3cYx9P9iB3qx+8p2wQ3Z9lVPNni48Ws2/iwYUpFvLOeI4Mn2K9t9b8eUGjBnXxuc
nn4kE9I22yW6f0Ql9/IVNL6iDEcTWJeyHGy3lRHBIdpX4VvmAnSdrrBIaiA4IW5WX7zOtGoye05F
JRkhR5JbZ5w/TtnGrRtp2MwI0fFc6M9JFXu+3mi4B7pnEWBY3vmL6zfuy9bA7XmsPRrH7J31/OHt
BiuD6ye6bL48liwoHmjGT0E+lxLjKFxVOtrE2TauMVFTBum0/p05gec8axjNexQdcKqiIP1RMbgz
vvF/a7Eo4feqLtjM6D6+Epnv8peMO6GS17UlzgiM1Q/q1++CniSca/OXLKDlJ7+dZX1GPnAvtRJP
54v7iOFdTZRusR0tndfZCcjHmd/UDft1CZ6A+dYY8is4fBvi9DhS4gKlkrFNmeFsYsQZUCg0WE+M
tDOp87j7VXU8D502HyMbs+VRVHwtOZsRtf9PrCq9pJmRPOstmaZy3f2S79t5htWWcmPGGken5JAz
lB74qhzaa9YImBfpmGDLK4SNX/XurS3+3ZgdrwtxPx5S/MOOhj6XMa7nl8P26pWprFoUNDH2g7Ts
6VCtE60SS1xfPlpZke8O1CihrFsH+im15lAhyT1aBmXJqe73LBHRav2BTc38yi2c6soQRMGO/Un3
HF+hyDrNcqjl7SgYYl7yDB6QuQ+diCoQQNAkpOcYOdJL7lPpr76K8O/ApFH+NddSzi/ioUSz0GmJ
Dp6CpfKxmyDHictQD+rHGdfuXjUQFcbIKfwhPsdg4+iwO3kFWgXm4nEXyhyFpDYWUKkzJ+kRBu2P
RegjP3wHQsjiFiQkmTXT+nNVOyAOq7T+FHpKE8sIHM71lro4Nq1CgJxrVJxdLgcktPfO2SmH3GL8
tsTLj+AL9wGv9IDBMEW9YPMpIMPqCDvL/qq/3kcPFmnJszsW9/mFyXImaqK3eUVGeObfuXtKFAe9
Z69EDTKHgC03/L/x4Tngh4isUAj5xdDZl9AbT+nhMKbMGckDCiXurcYGYuAGUloLey4+cZiXBAlO
kpVKvBrd+va5uLAeiUPEq8qOf6egBl/Yj6UN/bivTL4vFLyhhqzM9IlGcsUB1ucTt+ZkKH5YgwWH
3BbIQuTVnFMAmOfeeNG2SgmnS3XPGWxQMGrAvQnl1x7G2A0J4PbRz8zBh/u+CjA4XgAu/s+1m5PK
M+EAyRrOOL1gRNiCl3CDcMxuMGzuSiDfpmTVEaY9/Xs4hrm0MBDsafRZobPRzZ0nwatFTm2JmU73
Cg24esuZyqz27zYzH5tG3pQ7RS49EuKF8HmHhXnVVGCOXVTHdKHuv9aKI3Zn5KfWWFpwfYqkui8/
RTel7qNSi1zK5uuif6SEUgdLzrdH60+Gyh4IsoyGUFZJ3b5YwT1128OoFoXwiL9lCLoMhI+BVbmU
uhcenBVbNy/3rwaHqY6wUkd4LHvPGbotw1pG95ig0vccPwtFo10ZgVh/QsnS57iHt0aGG0DxDCid
M/9ESNBrAVHHA0ETRi9bRvfcE76VXn2690Nw+YYGhBwZPHv9TwVwjhSHAnfQBlNf5mnLJZU4ilB0
I+jcKybW/KfB2Qn4BU4TGtKYQaNU2DVDjbshVMr8Wgn0XQfcpojsgZAv592a3RecNkAxuAKcEVT6
0VnjeF57hdH+CUzwFV0NC4fVFMU/e/ClG26EDSvfyZC1P3j1cShPNcPo2Y5SWj5xNkz6fVYizknf
bt/bei8RXc+MFPYfTZq7lvbB7R/JyrKB+Kb52v+NbWZWOKX/VoFcsOd3EgR0BgDkLHkJq9Q4QnLz
tfiAUf4bpfY1FvUdC0mR5p10UPa/XhxOn0IM5zQAwDXtz0DaNrQ5iFc0cwVrEuh4eVDv4r3f1XSy
Jpikc9fgQK4gAfVqv1jpGAev7RPVQpRGeumWinT+FoIH/KKxlXcqysTSuD1JnuS+qMHAf0uk/3n3
ITmDhGOy+lcKxVxXuE4Clb4Z0D4TW2TX61Jf2OTax1PCCK3fgUSGHDhyOqjBU2GkAoRzSjFfCz8j
ke2Fp9f1ZzqQly3flqnLVhv00yj+mMrhQSX3OorKn5wk+/pNueXS142WbwfrjYU3BM/lAY6fdHuw
QpAAWs+lozM1jxJj1fSBN57v4hSi6ccLeWAMUi3VYL3qiSacpL4QMTspgHkUYVPPOrQevtGlLcnk
kVvS8r8nY8SrzOyT/5lSFj0jWAli+8zVIRlALlAj+kFJRLU2EtRIk2UYu/dtQg0LZDIT4mOg0/Bg
Yxm5kn0WLI4Y9tusOxSW1dsyYNdt3AUHrbpHEazZXw4k1LT6cRwMtLi6DEjR/3Yb1lCzZlf3X5uE
rLPE5YerwgLnIZ2hHc5Apc+YJm+gf6pe22h0ACx670aS7RGPcsss2gGBUiLfCznFH/JQ0F1nGRsQ
TZe3CT1TyxyCB/HVckfdwp1K0F4PqCrFnCZgUX0vJ/BpJJFRm/+jD/H0zcqH3XF7FXtGOsaNSniD
y+6qGs9uU6eZ4V27/KFwdZgr9LjHek+g3AKJNyPZL98R/crCmHNuTK6mnlJvpeb7qkU22uy+hvGu
9PIF3tSEMAVNMe/Cp0O/b8iXzPl4T/Ye66LQAzc7D1zjmmCEvBWiP263FONJhLX9CF+SWBHuglTq
bFO1sZu3V80j7CkUGZOndNRzhMSPi22E+bDQCCKMsr9CSehjAVeSYZpu04sTgwD+lgozqFdnERiR
UPQAGvR1JewaM6O3/489S2WYL2xvk4r5Iy2HfZrDPvFp4hrsAEKseruqQGxvhWKOx2YbuQyYCExl
TcXrENethQywaCQEqvcoBNi8TPl8LrlYg/mupVUqPFNGjF/Ft2D4zUcwBFVwmT/LeYpNJOEP75AM
EO92oXo2bFJKLatfrnMQeFvd8F+9QA0hafzh+gYmOIdpNuQAqAjCbDh7s2HoItHi0XwfMPZ1b+4y
7C3LULNDuUBzIXPrWVX7/C65xyc/FTIIZtPh6SXa6WPlKgFl3145HUypJL4A16Mq5qdQ/pgMYsn2
GfotE5cJ0zZ7GMbA/0+rsTMIH4k6nfmO9HktaDwfe/FQNHoa42ts9qG7fQr7ciMD9alpppBbVPQ3
k8DcToeqedCi4cU1G8E8Irw/71l2tVVVr51M6PP9zYQSQK/pCj4URed9e3DsxpnlDQPm1c9xQ1dh
bNQsMRAAAaRxrp6wn0O3LhwiFGMZu+d04Yp7jo70lBu9vr/vCowo5TGpHW/CcjjK9QVY07NuHAB0
7QM864WTD9P30vqagNmdE7WnZIyJCGGUe8wJoF9/68LcTYbzaZCMPBYn+6wtZWUk4lT2GHV2J2lT
GRrgIhRnYFoC/kaGfBAx/O5TmySoxtU4/nUtvFiRYrnrfFnmTqNehRia6mOkWCthj7SMjuR2AqLB
tgdKIEOyMkB1T/WkIQpNK958/gSrXjN+dj40O8dV7XtrKpxxiJ/Grs7OSLurhCrqP7C2KmhKn/A4
5dECgI078ZlNVS1PwfqtQzXUAAZYY1yxd7M0dQK4lr0qfGUQwjapmqD+yqcifHZNZ1IVsdebY0Ky
rBFQDsrnpKvTxkGClgh/yNreuoXuA7fdFgFR/XUiKsoVh8ZWmjXjplj2mMlBgJwLFVphKn8mjRoJ
sPkcWKT3uHGy+lg4SCmJSisAIDrMMm/FEJFkihmp0h1Mu3ogPeZMPq1dWISH4ozEwxZK+zoD5SAM
MGnja5gTLfrW5X6l064PvwkdWM9skWdjvL/hXXZ1/gSgx7kW1v6dSCpL2+5FfvJlVkmJBUJSme6W
eApn2RJ04IiwefEKbGEu2VeMOkmXOQlm4COdLEtubvQL98d17HlddCP46UN/yEvrA9yYXhQQMNdT
4BcaM5BHUcfwhV2xM9kxxJ6eBGgQPLU1wsw17QEOx18omGx5uDtz6f3mWKDin9Udg//2XEvdQQsp
zDRM6ukja7mpjaEROwRkKRIxW/anagqSw4LZKlohS68ZSQiYBNVoGiJo4MFlga0JfFZPzaQ1hBwR
teIZQzCtiugMhchKWV0x7/M1VcfehF2q09dDlQoswe2IV0rlbZPOxPVIiDicmO4Ewds9YdLigmoE
cDvDmbJNeF65Md8jS6WXHpQZgfNC8l/BYwE2/XAndIptf0grAwm91EfDI6efU8VMealr/afl6sDw
Tg71dSkTqfqxvgktI246eSm5ieSC731YzXNNoNE1tYmVBhPR+HNoj1PNd3VAvIFeHBlH5C1m/dBz
Lj/oEaK2nDjnUt01n1X+nLnda9iYa09qDlrJBdDeSxBo6aLYYP1unhDxJNOtSBrJIyQsP7vPwr4h
VKnomKFCSfOuVjfIWbD3LRMhWS8b/wUkOHx2TnP1fGxcaaUqcTHaxlE03id4P0t7ZBuQQoEbmlPZ
QHkzrlmoJ7qOqNglWkB+p5uC5ARCusXq6jtW3Iz1eMy/4yvN+OUC1UNli6eQ7/SSXHj0kg1YULAS
tI9tSlBNyzFWbcymu0i3kaEI7ZGgBGfZ7HZ93J9aS/DCHjTTzlCn3gNZBGFqWkBiN/E7GjtXiZMR
w+IxXu5WacxRijjGPweDamMs4XxfbtQ3dWMA25NCW4n7yceul58Ojgk9An8hw1kiR8VahU6VkC9a
xK4FMfKo3uYIGkth81g5X9RrlLH4+f6inspB1Kn4xu94OpSvewzCiBMHzv7UTohPKccygRozhB3v
AHoDLSKnwHmE/ry5OSvAWwnvJKCzV4Fm9OFoh2jOwEvIVM4bQyobJnNhbBdNRBqTT/z+ZY7ZA7Pn
dtEdIzcDSq2N6WbtzWjlBDGnCLz6nti4EGeZukE61hgcMrXhkyzY83xJlwTxwl5vvTP9SkMt4yWM
cJKAdBVh5JITWsMCSdRO9i4dyJY/C1kJtBr8ptY1dfndxeDGxran7C9Jl6RlNDqhRbrXTT7c7ivu
y+5Ak64hhXjMTnYTQWfwtG/iloJE8q0N/7QH+Rkzt4c2XGS4HEyZaFEYO5iNZotFtiRkFHw+8zHR
2xYEtqhNPo3M5ySfbCARCJ4+tKcgSnoAnl/n5daHLHaA4ic8AptJECYZJzrLaTVSWNbobC+/Twm7
2MZnjBlcM4twxd02V9iuA1oVhh91E+qfQyFw4fu5BHNmzyZFlh4+dpBPZ8kVb3XACKn5BXcv9HVR
P3ngKy+/f5W+twnJVzg3kNi2V3KHzaeWTjYiYFV05/t3JS8QVyLgBhdGBTfj3VHG4Lre6tzyH4SE
UDypWooZ0Lx0rsXBE4I3gFe53MgvDuOfED/+Q5yBiA/fxgdxJHEqBTvGNFRDEq0dQaWz+P8BoGld
lHJLsX+hXk/y6zpsxWi3PHY6nIeBFdqgN98JDjXizFTqK8VuF6cXMYK2quPx7S970KPlDmSStwM8
whew3eF/RnfAzOAreSJJ4P1M6oURElNAHgUz4jMkToq0WjLpaF8ZRU8WZoDuf7CSrJ3vLrGeQGKC
0ie2HEiBEhkR5lZmJbzJMMeIGwWOGT2+MOJlWCo4WMIoDxABOIIBswoZKu6X+7T0qM936pc3lyV7
4a6AMPXXD8GwJDprqs3JrtoHa03NZHpC83sXAG2Q9BvqgZ1zMo+aSn7mLVnuuN+u26Jhqi4AHB9j
0W7SY2FNnFEDveo5O8J+0C6st84+Yti4hYEggWtdosj4PfAgcXsm0zVzhkMfjzwaroW8+ECwPsob
fXORTNcUT8LYZBSex0gP6ecbvmcT/ExjEnu1tpRNNE0Is1sLk87seS8bKZf48sqgaTWq8D2OY/3Y
VeIGx5wnQaR+WbP7EnGixLB+WEepRNNvPlYOu0au2lQWvrXIfPWlN+DtNht/CmBFgFGLnhGcrdgs
yTGnWNyo53gS7CXN26Kwqd2OUdd9uUJuoV3ukb48O+uMJk4iZs7lSV3w/sU6Yl1eruvCRWNGfQku
I1TO3bUVxxb0xoyNfEC9RaStVq0tEH9mNOC2ppVi7/EJ6jhvCaGK+n4LH6BIeQ6/CK5z2gPzi/5F
tEcO6CFCSiMOD6LrVIxCr0nUn9dt3iR+R0UMSACSlQqDxzcPv+90XGcw6NTgYAYL+7BaOrXUaQ+E
1ejZZHuQO17DwA6LO072ETNKgYU1Lnx2vLQnD6kIv6NP/gvAfVi4wE5cgPbi08Z43vQqvw3yB8uk
UCYS40r0Myk00rGYcIBuoIJu3E72d8iPbNN9lpGQz9FZiW+amx7RyXFOJZ7tcAZbtiHBUx4BBEyX
VtkTbdBwHhkcWlqC0hivNt6tX66Ad3LdYkOukdH6/KpYDXrL7gNhi2NylgOWW67t5Sj8DjJuWWNa
gZpjmhM0MvcBl70RGOmP0iD3ogut0QzacMIfdEeIUlKWP5T6bnkv3ooch3sqTEc2xIG0OSYGaQFq
C3ytvw5p9S3JE46r5Je/BU3SE5DcLraEmM6GGP9hPUApDgAkNTDvaAtQA0BCAKsoq4c+wgR8w1uU
Khe2gmgccY6sVgYqIlCosMNcJ3+auf86xJT7+IZKPEUZf9YxVVHOcdeKpXLbmwRX+SxM6V1mFvC2
Rp0F3qgTWtPPpo9FdWQFSy0IPm6VwBJ62MuG22NYOLYLVnuGkntvzPOmn82EBEDhddrhVyY5sfvd
kg/cmRnTdqkYwpWSdW9nzTwTS45SZEa90nxQ4z1V1GOi5tJFIaiHIBrtMnF8aXp7dpNpiWk7kj53
Hjs/vfc/zkvIDHeOM24Bqg0jT6Gomi/U4qIKFnk+ydKWCiqrUbKJ8S+VIuqKvejpl56Mq8nh+3Tz
l5Vo3xkipfjGjogClXPifeg2wQ0E4L4tuX++vjCcXkfIVaku9BUlv9cJWcdb9ki0kPnrrYOFVS/s
ASXB4W+QY72PadNQXazNuY6VI06322QgW9W767RRF5Gjob1cz6PlcIpRat+iq1w7L0V3W1yXaibp
X04WiFq30wvJH1PdaOcizP8IMzttuoMVYJSUTCIQoMHaWihXeDcRYKfK3/ReKOB0LmdLeas8FLjv
fIFZxHK0s3axNVqu6U2BePYWi5syEnvTqe3w56W5I/rMuxxf5FFuMZvlAZGXu6U9tF/IQmldIXn3
i8D2Rc9QNhapYzb4Q2XoKEfZPe06RLID7HHENLLFLknovxxE1V69roit0W54UIgCj52TJu3Qrh5s
fLMJAOOf/nTQvdXDJkpxfqLDj/eZZVvVcE8yv714wNnVp8VOpzHWGWYZuGjDKxJf62WPmHUizbQF
S+QI6IhvY1slHV8y7s3ZVKQ2/y6Goc9TPqqyQe93kyXOOeCr4T3QxWes6xZKMOJGy1bo6mTDtdyx
qvyJCQKWuxr9noQTvXSZ+o20LjFuwRkjHrh70kUoBGVUfhQZnNZrIZhc3BZBH184HCthQHXUXzkT
NQoZOTMGYKkuB9+qywRBibXJU3fq8P/PO3eLRrXY9ped9/UuRUs0B48okz4AwWNNx99vyT1hC477
1dffLJmDoeepLILKG5T1B3eXIs4pznUr3c8RHe5zN2eXSJ77m1qDGJ0sxBVdpY/H53huxY5FFNMR
/KWMG/CYwobgqiJfWusYN9f6XjVIRacOqVSWSeNJl5wDn5uV8uzLZwBxu+4dOeyy5viQzTi79arT
pA9SMRF0XdRNFZAgfydYnK148CXycaFNH+nTvQoidhAiTIaX8We9ru6BR8y3+iWS1zuIvxUvjWkZ
r8tO6FFjROuwMldeLpbKiG3t7omjBOunStRq7eKGVixSBJj53MevjWCX3KZiapclP84gCZ7qZCJe
j3qLURab2HPjMZUPh/sfH7jKfHAMFDOB9otKa7wIexc4RcYtR3fjC2PqOpVB0EEx/5xBUY3M6tdC
dpS9R370MembszdNFeGcxXBlSteZiSWt4KP3gJBekek5koKQ4QE4Dpe6+Yfozo7GkgD4IwoyoO1d
HDfpegzm9lrS5mEuI1YtQ2ocFuPWsBCoI/mykIFbU7yoda6oarMX0c44AvUPxVimrhadGgUI/Dau
eHFCMVvo6ume/qwRksYZx4QJaaHuia5RT4yuO5F8Di5ZSMN3dHjRoNr5BG2g9z8L7xq8Kx+AlUad
QrqpjwgxfdYyTlGPfd6I+Enw/9+2G85wJ4Szj13XpI2R//I7yRGeFuzMjsmp4akmz2T7TjcPmR7F
+4B4PGfyQp5YwIZ1+9ORfFE8HK+UimcOiEYE2bmDdRBqqdIxe3sqGXOqhdfz8sYagoVKhwtOwPCQ
TCxKsQpYcrQFnKZJfguc5wSr4DT+LZ4FvwOFhRXmbhPVPcigwnIdeSwocTytAoFIlsw6qssG0pv3
XmVFym9IhxxjYGDCMBP4FSjpCWTmt54iSOPv1QR456JDR2en0NSMKC7MkeImm5pepSdLDqFsIhbU
tYuu98F2uHQCZP7Dn3cH8c4dYIRadWs88YFOmmSKIzydyh1drmRb1esQmY8N22iSqT2KW4kKjJjF
bUmN+7jpDa5/OMhj7qEgvgkjcrzxP/OVvcFsWl7vqjYbjqsex6EsSoK/rxDtcXUq5xoQG6KBGd7V
Tr0U40laqJ93NWORE+xz29SQQExKLIcYEocok0YJa2wzGX5081fmPUSfiFjzlnFBegr8XE3NNuBC
bb/gVg+Xw3hVIHl5ciYf0XDqe1l6zrLG8nhjrIymPvLqnRjWAawlD88zij2dDmnJquxy9EF3lEx8
9tP0lHWkRc0lOWQGbzukWTNrfHrd8elhppMVjRc8PmT+Q7IlbeNo5Z+gfs59ZswL4642qDbsY5cd
GkB3xBwUTHBb+zA4LkewhX47IiBl4XfoQrKIS4jUGhy1reNUAyc1DtO9API1LspcPl+rcl5XUL32
Jrlx/TSyA/bEjcmK3pUi+QhcYx8ylvlwRiqPEhnNKvEWEPmfh9P6cD0XJnpswjV/qdjxii/g4kVK
noLki2uH+k/Ln0amgvZPnTTWcj2l6ZnGYY94yrw+HiAfppI2/Ot/Z+Qoe/xhx13KJdM0RfqrL78k
mZHnOMguR0XbfE4HQ/43P6rtRcW0wGkE069K3hDdae1dPsNVKlckvuR0NnCAIIH7UWtDu/IFCQcO
sv+/HIb8J4bBEa8xOQ/z/3dz2350z4mxuu9Etd7Iu2PU0yy8V6UtlGA3YxzqcKinsV7ZBuVahCsw
4oJJD0RkQxMijiI/xGawfY2Q2oleJDmMP+YFOTmX/y48mSxodelzVH4eGvX9wtOa095+dqB0aBKc
XPO4M1Twjhq5SR/QebUWxuNNvIE50ZM8+4MbC84u7RWrX87oQabcNlm52qnC3vvQYQ/XZFVGuHA4
l3uQYSN0BIqH1iXMouLGjR0MOSsUkzwH262DmnIfw5ZvvSNPb1Cp75JerTiqB8O52HjIld6VW9xB
OereALa0tVrfOhRDRP6pYiUBf1Q7mPB/F6RF1TqiM4fSyErK1cDaNm2wpOfYBov3SYuL6XkxcQn0
nvUc7fLvzaM+v7MIBpqTHQxyRRBs8/f9hWAdyPP9b24T3nJJbh1gWZA/h+D0g6HLJ+yui2xrpig3
IfZdPWbQeDzTxnAuEiAVogwLJjPxJpBpLyO4qhkj+bw1A3WIMXF/c8ko2jBK7T3GGj642xNYexNM
w/4bfCf+59H6YLF87QfiMBOOL4W8qVLZczBBNBzp2qxL4CtlbreOOxFel+07IDniSrgkFp0J4G8n
7XCo7NPF1arebs+v0cRL2vnynPqoOaM1fXtoQl6yCx4pRMQVn1b9GCUxT61NAJdkO7/emLar+/bD
TH6wJpTXR7t54lRggdxDk6PTwHhJxSV2JolQ7e3mS2qcyShM7/ae5HHYvvFKqjnGSXtBL9yLPIAs
Uzl8ktgkEJOcynj0Ibq+ZBJwWTRIa2U6QWZJIPb1adBpBU3nVhl3q5YbfwAD8ZYaCT9rLvBIcb1/
y4i/GMlo4t1Q5lbcPYJwm0W01weCc+Fx73uH/eJmfzNBvNiHIZfhWPRCcF0TZpnX8nf8B08OCljT
NmXgj+Enh0rUtjKlaDYf3AgW3N36mwup1eg9EOSOZzRwCsA9LjWzcZZ1ESdQ0doLUXQbSSJ5VpRs
VDcpZe/UybC+0fKLjxJVdTfQnAKPjVyccsrL9nEt0aKReBkKK4h4yhnS25KMpHwqF2Pzp9W/CaUW
kacFV8+6D+0okpISEuvJNVg6Ma/mC2DbebSBFP5cVFVgOwvxpB/1CDRvCiMgT/cqYilbuXSvlsTd
8aVp1fLQWOr5Gl8XylMrOJCgobVeKswQzYMwM+R/24WqhlugYEzM3BkRhCK/yOPQwG9gngu4WKqY
TX1vleDwEPUIvJRqyin3XE/QSIWjLYCu2U7Lmm2WnnYQ08Hr6BGmaCqEW5yqX7w3ww+MMdk8BTye
1stmoy0i1qkfEKw18RwJJ4bPl14h+VQVIUfrwL76NK/4Dmz5Yh0QX9yLTuoD/6OhWEyX28HlxSNG
TMOhoWr3m9GIlOAmRCtGn5WZ1klAmwYe2gTEBOLo0Sj0G22mI0yP3Tgs0aGQR38KI8l4AgVDHZSH
WRB7PK2ajDTENany7Dz4tn96PwEjhB0mZxbnFzQYzNJzPiYAruk3+/5qffs+QVNg7Q9KBftYDKE+
+ZdXSxXgZJ5muqFQWlKI82cZ8eA0rNOKiW2ik4U2MtpKAQ12zJgls3BW0s+cqDQQ6l7S+nIE7vjt
JGI9sbic1a854Sfw/HpxQXBqdPK+FxsHx+bDcQ6yee7+Rxdyd07kpHtERXcui0W9fg0EUF1ETL4v
sTBMajp2m3lGzGjx/VyxHHOAc2ppz28o9o40giGbnvDq1pbWYhExlDhiPRLcaB264qPfuAsO5ges
D9sYaZudRuqmW5QhS+I6q/B7YIDruwpUWkLpUgvSOvjcsuhtAsP1oFqM3MFNglrvVPWPZRb18wcK
MgQKlYNw2i/9UFB/fcUNoNsYKgNWg4NoYXrV3288hyJactrbJRr/A+sabXx/BIWthHlyAD83oZWp
3r39rF6AVZM2AhMj328KBJFbmAdcodhCBk2DH8tV3Z54Yw1Rvtz9zGyhxbhIrKoHN/ZwNHKvRzpM
gErcKxsR74dQ9cgJO7JSVhI1xu/ngnH8OHFpTt15DtY1rv8dN8EfOYKqEoS8050zsidQsv83Iy/C
Kq2UdIEpa+4FIDKC4ixR5vlLb/MCacei+Wt0bk29cZiKq/s8fEqbKq0nX//Rzbbx2VP1x8yhid3I
D1+0v+wWcJeqDW/3Lajo+EVKUITiBCJRu6LZgHW2akpPJMdYWiZYFNPS56Fd4QN3T9FkzPUVUpw9
Qoi3PVG3XZSu/FEufGQlDou/IUKBRaQBU5Fri4fVhRheM9LsigLJXPz9LGhC9GgF31u6bQ9880el
yEu5y4a5jnv2E2RauQJC01ps/g4aY+6nERtYTKvjqoAwGnEzGG4Elv0xm1X9mOZ3XjlM7ipZCtUT
CSKOyMk6vgz6nQz2BL2VeQX+20dgMWmnvXal6yIjjFQnzWA7zHO2QjsVzR2LO8GFejPG4sOfJIQN
UiutfX/z5YguINw88gnpAkvMnbG3wbK/fS3Hm1rRVMOYqUCGm/JPGw96Ky76DjeHKkJ92KqsdwIq
/sN7DF2OooWbX+JhoRsRZp7azMQdDmip2R3JryJZXmSE0V/ts9vFkp4e5qyJ0/wLOcyLyhNbJYtZ
y5noUBAdO7QRZr6IL6B6E5UpJuxIFxH7EbE97fAMaIm7s+nhvKqfbBn2R4YNmrWtzN2+2WRvPJSM
zsJW3/wYvvYFA9vQD0OmtG8dMNlM/QvVfcEPwsRo16sqjF5z4A76qtDWLLHQQZu+Sgm/HeQNR5Xz
cClGBbOlixBvXcfs1hfIwvV+RFdIyamhWkWMGJx5R2JABHDt6GcubOKpoeJLJSCP0cGZLEwqJfDR
uTO8VyKtP1uEL6bdtWxb/BrJxCKaVT0I1xtHC06ZGYxFWXRzOhCmoQn4fO6YxX6lpDXEXscjUYao
KYEfWgcm4tY4c3NILrz2IpQ/3mM0zHLPs7GxLEP667xzWyP+05CpmyDUummzN/n1FedDC53/nehH
+r0F8HBvs6J+u4TaPYGPNx7hzwO5c7grS0q2ACA2pmIReO36seexG7GwQyspEH0zvYWPU+y2PcRp
EYVnQsZvMhkXNKbHggibb6I3k2s3Vg5aYqVcBDmwWRKJEzuWBC4+AFNzUd8LMRUhT/Qk6hBWXkCx
A+8CdnatkK+bGeH4t992sWK21oyv3Ku8yBG+zzXidxLxbifGBsMXKu+GZVZ2MsZg3F5p+aLholzD
XW+i13CRY430zsvKascJotLqkYZqpQXh+H2Urgd2xV3rSGqEOHwhIXzRUfbt7PkwAITIM/rUS9tt
Jc/6OOeQyUfdV3dfNlXqtASGQvtG+AUcTJBuWP1uI6/Dnz8hbqTpsJsWpH9TId1ATPJ+Z9K1YjV8
u+u/apmmtUaTg66ZfMPadXVIHHJP8t6+DFpbCbNAg9tINy9iYEzsa+gTHODyp60WEhJf0Rg4jvfh
mnX00RjQwpkonnP3oLsfk4yikGE44dV32BF8PbHLR17r5DNpLb+tHlf4QDDBhVG0ygi3wF0UtmLH
Zjf6PnYY4HfV1Ix/YDh8VC1TnevYdZJ3Sn+Ulaxnw8rsNqJGttMXbm5jy3+8oerro35C71/yZJKi
D4z9kuv5CDIh8iG32zdt+/PmgwmVKU/oPSvBjiZMF39DU/wXnZhhIOchWA5ayisVojIfkemYvhl5
GIcJSlV66NIbv1pIIExf3thoMB/CIF34NiaqnIDdN3TkWrN4ZKvEzyFfUb5DcxcnVcoN0pvWr/N5
oHiG+j2BF4izcp9ymU3mmgdTR1+B1D//kM4V+84oHM0aUDQC6X6AF8DYe84nB8EtzGUvjDnWlJiy
YUt8wsGfRzJsGk0vucpxvNtJMoE8yMVAYeOmR5eumoEL6X6U1rRihLMdzukX28BdwZesbOPFYDsv
udi5evUg372RPHAEHYMCn5uJFKYY1j7rUwn8otYibGzo0xNVD13QowQgYKpnvMC/59Ydogbt4f9q
O+wc2cbGEeM40JfBn0KaTO0IuMTrIJJeCmmLotpfUjqDKCBJXtN4Kz7Dkqt+HTktNRy9g5dD02LX
GU3qZLnHmAAucYH6zSKY3s1ZnNTn1Ry6VfnOlFV/OPexwa8ACOVjLW2WKh/8tseSji8S4EN/jZ6E
oHKIQn/1/x8BaRrC0n+DLk0RzFvdqPNL+pyTtQ7tzN81bN1akTSx5/pQ7Y7j/w5NhYSY9qV6Y9M0
uo2fW7QrcqUqLrLHzXVBXGRxxozJuWktiTphNr+1aXZ1Z7H5H2/lzbfTsAYFjWumUXHEL+gNThfa
iL4rPdFA51IoPlOA6DzLI1ruN/llANzNbnMlAW4beg2siF/F/Ler0Hgbgqhgu8aDbtHitqIZBmNC
MWiB0pyJbpDaRvFKG/D78ufN2BPvEP9c/cmyB7xcD0MpZF7hycC77dPrbxTqqTCxRmEZuZVU+KHB
EqhX4J6hzNkijHxzVdS7w4p1Bix6NOX0QBv0/YVLiKAPZieDQIxGoyQAoNEXqezOPDQrhRXRC0hC
TQmv2bde9IU5myRdNPmLSAOg/TdbXLdt0LbawOwBrI2pmKVADswFYMoSudIM9s2+4uB2rxntr9wZ
QSsc4Zpc2Ei6M6o8n9jsP4HuGTAyOoGR0V3eXNTYktK36d6DPupBcn4j5Com/8U6bmQGdb8dl0Ih
4LWkF7ou+4jsYKTSNu5GweoQNSYbC+Bu/HdsdsMHgvbZMmJ76k8hRadho1x5+cQr68vaCOyZOQv/
BudjdwZxyGSenWJUEuAv3ZeRtTZc1BYB/yX2ybtFg827shRPxcLI14Crprc+wouBeLTUrmXNQB8N
hLST3wunTyJa9Sqm9XS4C+fW9huJKf9j29Df64W3nQ196nMzQOgwR2JE1J6KuE97w0KOd1QDY0GO
suzNje61n3HbNDbHJ+FAvM58tTcRDvb8jRRj7oU1PwQ4gdXcSU6IV1Kn0u9ihhmCn5zMeTthFWC5
1LIsBuXYQ0WXSUvSv7NSPgB25GqwWr0yxsZkQDaJM8Wmr2vHJy9zOzuAZQa2aoyd6f3ztyOSg9Bt
uem24bJjKVEOATrgv5mPzH/UaWBE8z/oKoTwTFwSIrJH0xOEzqO7NdzAiEo2tlidxftL3Y6O2HBV
B//wWR53kDf2UPKu6E/xTVLArRIAGhCXtdr0YgrAX21RnPWqIa5WAzQBi22DvtrN0mttll8QCn/J
qZw7bynkWUR4WR8+5DZbhdbmh/IuC/57n682talVgawa9rAvFKSkvLFo/kPjS/yHh4ktXuOQyXAj
VMll6W4ntikTZoMIgRJ491FNOAnyMliZPAZtkWFm7HhaK+4VYbE7UUb0wwObCxhGGGi1LkTUnXXw
MvKLcJxFfK9j0iaDV6FQ9dKpD77tp2bh/SY+3I3M2RhlAPONoIDsr95TOEh8nPP2ffL4L77vWKhm
2b9gFXe0fAQo3DjW1SIYsRdFUqE5xhUCaRVljNtctr/ePdmPeonfirtBB22sJO0KbpSb0f6EwX+g
2XxeWuexQ+Lc6TorFDvILrEHd9GzOIuZEmZ6szyqdDkWLGGLijEWZoynh93maUxiIuKMvnDu/Cdk
ZnS/sKbUKnfOniBlph6lILAPRBO1CbAI6Bt+KWzX5DMwlN2CWzin7XYfB3fhQ6TjizGBfQH8U8bo
IOF3AS2LPHccwYNK4aBBLv/37D5hy1ui7SFMfMFZ6BAEEdoKFgGCWF174CVHcUsYb1Oyu9JesDV0
WlUvzfgItEyoTopwSZT8EoyaOeO6jgftTgpPoFFmmN/gDtkSnX+yRiErlD1Ua0lwiPBlpwG74+2B
ra6097MgPg3z735DldRRn8+4Z0S61P38msESAqS1iwTRlXM4plblDKHllo9QoZBj8Y9lHtoueyqd
cCgo3vDn5x0UKL3xf7VdFxhe775P+N9EnpBe/ctt+BblquaBIwfIUftZLaAJrPftcA19C3pFgXFG
Xh0Js7+puPmp+GHPUzhvQoJcFtNSVxS5D+UjCaCaHkzE4DjUdR6a1hKpQrjDcAb5u1TnrciOhMDT
NiQyaG4rSwmPHa+wEYZf3SSkkVgayHVMy+Lpcg/lX90v5nUzcKL8Kgz8nQJ4GN8ojDbX4QjEHMRW
BuP6DVEGAdV44R4qmgByla+R6fn8MbL3OgIF/s+oEvori6eC5ylGBu7OkwAVIL97bF8CgEhksH90
ThKPFI1wL59x4BwDahXe2S3SNiSDTcqEu+MLr6rBsq7D/V4MTpJLDZuFcjWOpZ6dHPScUJ+PD7HD
TPkrR0f0SvukwXdAkj3qGmYc74Uk+K1YaYRxmnq+516wedZpVUCkKliOUXWxCEtG3G9xAmueHvK6
lT0j5jwm65gr6S3fsZ3lzvo3NizXQVp8FHJKRyzKkMaQT42iXqY2jx6oGyWBIDCrEQsEBSPiY6So
AX/R3UoLcgRzWdi2Y/ajqk4Hdpaiy8qMjs6Kr1STytJtMwZHnEmT3ZLtWRTuJSxFqPZKZsPoeXgQ
LsJicnQIMB6oh+hI6KqwKJSdvMWDCE4E7bbtVDmWGMQ5abi33EJf4k2BhjvCqRKhASmtJaOY1EHi
eq8FaPbbGHekPr0B/6qfEHYflkAxbMv7x08PKECq3fC0t7my10WcH8jt/tIolim+k6vNrw3yNWjg
6ltoSN0Gl9qBKOfVqIwIzmhKol162UoJJZ20mC/NNTiTv8pRHo+D/3sB+QzzWly32z9bGCS+2Ni5
9uLwCVF3m8sYH8AQPRL0PHzYRUTC6bzx9uB+d1XzS6Ejugg6VhyehYroJTemG1LqHDeEEHuPNL+n
76mgysWvF2qd3dzm/jwMdrVvYr14aaU8XWE46h+Zb22bDkbKBKkWFsO3BDF3rSg2l/J+6tADUwIl
9uiJZe90e0UOEoCog5XpQqvAPRTvP1wymaD7/WQloiRC9HFRinhH8C9cgl9s43nxh3Aa62c+UOZN
xOAfDUou6c+FvbL9qXqKRiISXJ4MIT2pv0mrIlG3LH/U+gZlCEYee2m8GNxfc3SFpR3BHMGJ4KlB
IBA1IRFYazV8cK/Pi7DJFyIrKT0oVARzU5nBgHY1agA/6iWqYcrVKUwLHTIIYCKabm5ETlJMzjWP
wmyBHYqy/Ggo+OiK3JRzSmajTSzn+vzm5dSwpT3E5UWfPs/Lt3XyiuTUyycu0Szmgw++9Vj5vv1/
fxMh+XEmq6ApE7Ccm1xvi11DlqGZ/cGj02RmPLe/ZsLNgA5/nlyS7JbkEffLVts8qXqBEgEWxJjt
abdSkjNTBfQF0XliU6nR0mseyfC1ThG1HvEkq/E/TEMXDZ/4tfZLxqDm2FGE86ZJtlRqv0TN4DVs
16TgSzbiio3vFapITLIVmqABlVEl8xcZb+kt5qguj2F1OIuzC4aWPCzsqZY59C/xhbtwUy6bBbpl
i3R8Z2l8w420UW50A61LYMyFqp5OLugmviBXUcuYbYbuqdWldMhcp1RcB1pKU26wh+MRL3Emgjce
bm/EvNib1HN4DpXyzWUPnbGPk19HGXfpXTA8NdTb0sk9ryovtCNGERq9u9Y3nN6rAh5b6lGPqXBd
nv1ckc4td8faEEwJ0i95zlcleVVk5YE8Ha7xqo1+DA2iqz/Rguz4tKqgYa42jVSTqcQRTG6D5Mk0
dg1ekDrToniTdOEqH72jAlBMmVvCcYJeJfg/esd/LDoOThOEe1uuvR1dypv/dOxciFeyC/A230jQ
XidR1QiBFcwtP2mRlb5wQwGw9YXUlFFjk5vvPsSsiWcXR9fNXGuB5kwNKV+sJr2aGVpFJgHcaZwC
YTAQhyEkmx45vB2x7ICQu4r0QQRKjcL+9iVueZ9nt30UepAb76HlkJuXtHmfv57st9gjXJloW0B/
plfW7RbIFzM0ueqdo3l6JyO6vPSHJiTwkZcgSrNK/vU3LgD2bl9uc30TNtrZE+iGcslQcO6JEcgs
4USgSBI2ZX2sWlyY1TJhwEUkmLuj2bNZT2qZ9ul3cQh+OB/ygUpy6AgqHxk4FshrGj4BeMGXxKSd
RiBCXffRSgTS9jZDc5uufnYOzavR9Boek2T4Jgp7KvMrcOd68nHcPRvDie3onlgarAhTQjphQ7d2
0AXL4gxrzJPn9S88VHznc2YXi2HYc5Pe9LVqfexElm//aKPFr7/J2frsTRFd6nKOBc6NNys5MJvN
X869nv7zrUFGb9uuEbruUXkonv6tcc27JTM12FTxIAcCE96lFcyt6v3xftexZJij1qSnCbuZ6tNT
qynbxg60j6m2e4Uwj1YN4iXI2OCCleNvlFOy5dCRbUPGCYm+7zItcBDRdDiPvahfOoZy4SrPQBxI
SDnkMbTmJVaiVyBNkID9BqokoTu+9D8PeTofPtH9RHj/biKFKKukvcuTuPJSQ9SgrUUzUnS4Xcgu
Prf58OaYoLjblKqhetIoQBRkbQfXRarhngEgWA870zmX6AjnKA3zESzsBPa8otl1Y7jnwLzz9s44
Yc7WPDm7hrk22pNykjrt5vpmou5I0KkIGM89A30cEa05fAiAW5e3FBD1/urALV0IaIQdDZ71gNPc
LIozqGKxIgKdnY8Xr6xONQoG/EK6/Lkf18iuHPegVnnlWg0brHQQY61qGjIUpB4PKJjTuOHGl/zM
PBmZqbTCWgx3oEKyLkqGjxQnW0HAddFKTda2rc38ay/nNbLNNNE1JUh43icKTZymZuQYScCzvOHP
xC4PjjVwxXf7mTv78Y6e/M8dRSQhv6OEciUnDrvcVIh/0KUHK2a/Z+5OadIkHopxLkNJkp0QTNoV
15ucwfAf11qpj8jeFm7yAH6syzskSYk15fzu1hKsNYV82O5ba1nZhbd7xGtjXDnCkl5PXJD1DD7m
9zT5RfYZ8UuCFLDPPlTOH2XeCfOBPCECfvDiFRDL3TdSM2cC/e5+cUgyqYPyngJw30hVujs0XJ12
oAkDzWbQtajuBkI66v21JZZV6rG1nr6ojK5HO0esQZWdSRvcQtrmZAGnEjuzlZzcENirFxVJmwGY
BpygNEsrsu4xC+wh3io38/8gNo7CwW2peUNqmBLMuX7icJ+fSWXhr3QoTLyTwkQ7xrfyETcFIjLY
o3rhnqz5Pngd5gLCQWy679DuHSbGpPiPH9veLnfkTokzy21swfl2jFsk4pp2XJTVrLH1PbJ+NI6n
91f7rJuz7XkBJD5+qOJLt/H18n1BFrIgCdjgut36WcGheroOHHXxh0YZPXcGSdZNJ4CG2lJRwCwl
NFKSuTow5GCby0NZul9ughpDoas/Nwsy24GwaJBru7BKjv3Ic0fxISxMolkT3PDLGvlEgf4gkG7u
ERWQ4jbcvpEep2FVlgZzlmTXTxiNeBbijj+3ITwtFdYhpyK0kxjDhdZUmE39CNEYHog9cK5kyCwD
w5i0wXSF1E/y8VriemYOeCS4jLCQZmfbPrC105vFmDhRzxaRr952fsvqMabiGNdeloXyBEIXMeEj
K80FhmGSMPnQquggfxHscs95oWgbupE0DTD1PymeAc/fVUpozXmUyTzgyxcnzt4FM82yHuh4wMgx
IpgqCFJ0a7eDGnQQ+gGcUwchjBvJBRfO4MY91+hEExPi/rar5tgv5CAvh7eVBAEKVw6T19Ajywda
5gfgj3RZMkokA0HRjUsPylx6/tdaRQ6KnlcHORfbYIHcZ0bF2XrR5xFFOSJiGutP2IOnT/v+lPH2
N7ylLdmLCbg1A5RNUW679ik/+FrtI45Jzw/I5HHqLycEItsOJpOZ3WTHqiyhCxpJhemIOhReMrvW
tSDUzs7Ly3wQcjWV7zn1x0QIgTd+W84xWKsWE8KZFAbFto/ZgBDeMSNtBwOTt2FJRTCBU8ns+sV+
c9uZbyHg5T2GdRe3lfeKV7PJzBdi08ZQzkgO+/OAWlB8y3AlltFSozUr7DLDAaYdjuTprvrxbRXb
LZP3J8pgEAmN1z1DcxplszoABORg2jVR6bUiHLgPhywXNVVwR+25RorLQiWaBlUFF9QR9KI+esXb
PebpShaRR4Q/Z2xyWIq51migpansxyWqKFQ8hm17Qws1WxeYZ5Okh4EKxjdqTz/eJ1DFlvnQX92w
WpybpmI3yRyofsOH9UcyI4U+qbw9eGRSUX22RotcgPi5Pt9nMPzCtpWBhfN+6BaeNzS9c92BU/EG
vKNhi0Ie11enZrKvqGoVHIDsxCIkJnVyu/s7v4gqHdKZHzRrO5adYYpEyqKl4OAwrbW2uOdacPSs
WDwJ1JcqBJm5CptOepvSmL4SqeDCgxT/vBphWifYq5sckmeeJAfuRoMQalzbNxlLeJOEowtlVBN2
WJj1Rp2hXCI5ILM3uSAMpgA1s7A71cMkNWmoEm63Nr3t5rapT9LYacBYYQedV7evJgAL8ieqG4FV
epJjV+65rDE3r37BcXsbzs7obLrPocZ8KpK77IluHyvc+GD0pWh7DKNxawdx3DKSJlKNKCb61v+A
pfbywnba0nkjxW9Dk177gSgTY+H+zV3MdgwoiPg1hYq5ez5KewB/oxWE7F3TC3ml9cYIXT8+IEXn
9Q67VT0vM6/OdXW7YiIAfPWy/F3j7vS3PKscCMfzPlWkjA7ZLutUn9mVDmYhCUeilFw5EhoDQK1E
4JGHINdPpUaFHTC/v62bfTOvfDOcckZAPqJlC+jwhdAk2l6L6mt6cnOKMSoZmR6CqD6SB2R5L++T
76D5oe+5IYrUcobHsaA+p6m+Icj+Md43Ap4npYssaDUGsF8CI5PJhwwbz/Vcs+ELtnxla0weo5+7
tUTeAs8L3jriy7+cKvFOK2nxmrRW5FbFyrV1zozaMuITP150Ddfi/mlk3XkIWw5rOH9S0crUzgHI
ZFRgStw1chFZa1jD7CBOPS3/XEEJK40M7ADZkryZUUnybLNzeoQRzD+E0BDUYjH13NDTpY52S46k
CYDj0XpCzeCQIxsX77A094GiITTRUPJCbp7G3T+wCAlqAPG4zn4ypERqk082zz2jZyUx+to0tipF
rWn+8YffGxwmT4ZaFOlu5m+cePbG4fIUR9Ff+QGLFhr5E/iBjrrOjXMDoXNqRl4Ek3FRcu5hRjpB
EOzmcHTPLHUzDcE1CLpBmqwoquMddGjk1oL9LrrlVpfRB/1utREWY0GzGfZ/V6FXxHjBNWegyUQo
CekpRHi7niyvM5w7Dnr/LtTsulO7Z+oIBEqDDv3B9a80kiMqh2zE9/knvL4tsGh4riKRT3t5InXa
pBfMi0d7HSxQRf4vmX0zYRQCfkS4ra9aLkA1Nt3Wg3jotG84nK97yGYH+PGVEmJzQ+nX7tyGw5Ru
WSRKcTwRscQz3ZhKPGUUfIlnUnDF6MlSUlwcWEaOaMCZdCO1wAUpaBUpN8d4Q4NOGyvtByek19xH
PWsK9BvuY/HU4zDWcN1WBBpd/K33RhP9UTf/I4yBg53QZkHFopomT5PJ3/7g3ti7PJOa2wEwlQd8
ck9BGX7HfCbps0WyHjDN4JpPdGVhtTQLb9xU9+teq93WcV0n0gu6OphYwyN74IwHnwGjq1vxFDd1
Ui3mrYB3oedEsbSMToaG95kMf5phQy3AOpsZo58GGYVBKav3V5itJnquHx8UO5cqdgO7OJrojUe5
EUrthbcptY7Z+26QNHwbdcnLqFq78GvJjfJiRp3qMfEDvlc8KjfIHsVaIwSOh9JrWdJqZ/8xvttA
wYISqG4lGNK2mOa/Um2GG+Of0tds7dMXGKtjkfKKpNTDCQ/bjB2xIceo3BMJgJv9xEIe1gSiMLnU
KXwcQ0WQmefh7EHpBR1Bsb8XaVhYRrSwjBVpBPnTtOyPQR8ihSui1plqOofy12rFa9A1sWLikVbM
YCrUfYkT9ZOEq0nAX0fXXKN4C4ixm5IXQLXfzmCGAJV30m9N+6bmCiUJLg7KQ5Jgk1syrg7xb4Df
i1o/1ymM/CF4BJ/Vv98c8XBoMgGjJIsij/BnOx+W8yLsBpAXq4sQbstPhpi3lKu/HEzop0fzSiSc
mipk8AcjkXwzVz0Vh0Gs8dFA7Sn6joeeKarANiB1qnNkOnE0fY1l9VnEryzEKvqEum8qLHMklYWy
ebcOr94D2yIN45DfiZNYCpWNt6uv2etWBspXOL34c4WpxH+A4XGB1M+8s/uAEZgBFasjulYkl6gf
yxl+K/+3o5z8JN0dmOanwMrcn+Hu6WaE4Gy1ukMlR1IVBircosgWeu9xg3e8lBmD9ZRWJr790i4u
mJbdQf1g1kXDlQYKYVaBfh47mmBXr38bq0qNQhUKY568vo/pSYh5QH7W/yC76VjPpdX0CnSEO3kv
4tMwZWGoZ7xHlEForIDnE/fyY2zrsUCTnzW9ZDmFtm8h8HqL1hlzJPBe5stZ6JPh46FUAAHPsoLL
YciwfJbLROZFBOpoUWYNnJFi5c/hConBBSskq9Oj+dAsLTiL5Iz4knjNmvbg74tKT4IKDBjtd2fH
cFPKZNEwlH9bVtlE5ypKEzH89bs5qq1Tlq71MXULdeoZ29e1/A9snZA6kiQfhy7Iyt2m9Z5eRXLe
5kaI786dh11A9LXMmxZidUVDJVTjfSRb7MWKfwByWKEc2k9kJ9n7Kbb/9/bMLBN+Msmblm4UTSRQ
YQo8OLp/zTBNlhE1EBCLAwxygr6YUtN1tc4RsgkH1qDS6ciDQEVg5OtFqtcAMqeHqcoSFBNnDgQW
MiVK+apMnPD19dbRnai9/2ipQXHWmLNoTSO/uRSu8rCHfWQwbSpMCcpF771sH6OO+u9383WXuWFf
mnmXpZqI6m33N0KO5Z25te8CMC44YFfonUaqjqUVr5uMZlHtJThBOSSL6rgO93yVtk6Ajn+zmiA+
kRW9Ss0Yh0ZBBkIxRsSRDYYmtDhAY5rpvcmJSNGhqG43qx/mkcFIRrSKh+IAd/RQxIxK5uw2lZGL
LcxBexF6aNQcdmXNAFfTOPeBZHQjG4acNeIZ44VSEgYTda4OwhPGGDq9NVVLJJfVB5aToJ9nzXuy
9tXqNFWgsLUAcvG5eLrGAcQClYHnudEWqnhpjl3tPw5+PTzmld0xEWctgjni7jWFR5lVIJmu2kcu
mztcqlaFhLy5bd1MzYj+oTqZPAEDofaLNQuwWO5La/NyFOYgl8+5H/V36Qm02WAJZH4Lw4qaW6Q9
MbAAT9SoUOCa56Y1B43nnEeBJeHIxrpJSCvrTrW6n2O4SO0axKoYYevxhyE7tl3Sa8Uv05eMbq9o
IsYV/b5bu6l+P+sbP10Q21VM173kU0U51pbvwuN3Ecq0cs5tFOyKpukDXMDxsjBNQSpl0e0gWgAl
+KZHMWqTeWPGBfTD3YJZAnqSsyjduYqb9Ib+Jaokfa6e91Gwz4/YI2C4kVnu0rvVtEv19eDyU79I
90M0RpJfSDzjQxsgPhaIGwbpRlKVhLW+D0FrXSh7yHJaVQMrdfQ0TTtIhSLf/+LIFS/2yJ3F7eZv
JFUhk7Fkt03kGvsnVLW1ajpacnTGUFJl24U87yK5SBSnnvDxStc7Oes6DrIVYXOqT217PhJ/7FeT
gN0NZK21I6SlSKLV0LdZ/Jo9ycG3Gs1Hwu/O/FHa06JxzXa2081CRzSraJj9IblILW4GSNw9wjvg
JsnEyttrEfYB8wxy09pgr+t7dsZkl0VsPsizuhY+v4fRlgusyVWndf1RcVUjY7FJbO2I22eRgUkO
lgnoCs5p8ZhlR6R8S0pkdolaScMpeWy53IRde2Sh1cm/yKn+GzDgAoMML8CgppNLalMEmct71bkV
E1c/4B6Uz4JAON//pr0aqrA/iY9Hz4Bq+zG0uDAAlfcU9dlZ+HrK4DYteiq9hnhE+y76MnnIt5hg
1dwjKQwtnlRNtePBqX5fGlquEyhMSxLmO1a1QpOKd4LUyekZwD6/ZlZsTMPbV+a35t10rete+KV4
Q2uUpjjkI97kglkJ9/1cZjRgyNZr0FbMTFty33Bfnb3yGQkvl1FrhKRkcoG0UVKTpxmoi+H6dsFU
p2TiJJHZ4uctNh8sEayFer0KR3emVjw19f+jheNygCVwAWJ8GjC6n5GfMkAllgddN+RYz9rSl6nn
zHMO7/XtI2GSmSUxv/X0Xx3AjPDS5FQQbSV/knaCXnIuXitE4VE/8wATOitlE/paaEGWx+6kufwi
plnfSls9BxxaPBLXl90u0UQXhq2aoRkhkeNEaANCnV9R2a2Cb03Z59Eha1hklwMXZaW5dXWTARIC
DwOHbJr36O/tbqAPcICG0b3fjhEzyD+n2GI/99WU4684jkUi4scLDbJz8P3dq4kqwPIzWI40PGFO
3q3qvjs7sIL6Qd8hFYe6kgoOYi4Zy057HKmEloOefJEvguBXGdSFUd6ebvwcxhVa03pxWvOA9KIx
TX5GPHQsWUghPw5May7QIkZMhjI63N1sJH7HNIvHIIoAi9mdyRNerYAby0ZbJgMb7bHUy6m8JS2/
ftVKVlZFTbL0uegBJ6bk3M0k3GwXCj3mBya1h/O6S3EaGhc2isEtOeGXvywkuEmygZ9Fdq0y8PPR
L07yQlhGNNSXE+QaDJlE93eOHR6KX8H6rKJacFqpzDea1RdHCIu8AuiGxqQ1t7kH073Efjq636Pk
PanHqJFA3osOJtu+k3BxSGYI5czzMMXWE0kHrEgFP+9e/qFL8xSBtv9ZTJ49xwsNRujoKC9yZGpk
a9Ck8Rc7QmakAKAlc3zdFE6flEBy09d+yBRy/bk21idM4BSm51uRrzy/zWbHYo6z4lw4+oUH0eCD
MW9JpyMFuog9rmhqwMcW5Z+y7mbMDdvHNLK0RAL1mzpiSw/C3GZO5WsHpH0XnjyaKbIf9YClk/OJ
5MCK1PFreCz7WGZBYQzCZ0lQiz6jiTi3jY+KpDgliJs8iMtLqphZibzlWm2UVzyNI/fllG11YQbm
JYO7WMca8AGwvPtV20RIusxtMHGjqV32gQnppP/5vuL4DlOhwRrgjrHyLWvKgoQ9UjmwWKdnG3gr
JrdUR36w4N/a+i7BVDjuPN/osSabD06Sp3brtKxsXYJY2YJHH/OgBClSYaMxSpks9L+AZnuPDtlb
HHxdq78DnF3pjGEfNBd9FEtrGccUlg/wD5a+jJ5LL6tjkXTjMArslG9qTx2zLC9HdlZKa8i8gh4W
xlHzPs/XwJBfncLjzV6h1xeCYG58+jH8neLdoOhrha5Eewl/J69NKSuQNQz1whNlr/dFrmS6zcHk
Vjp86gL7WaLqskeEpYAARz6HEY52bCPICRD4FOIj+QEJ3f6AnYUrk3TDrSgveNI99FM7uuLSJMb6
7Nz21hRtQyZ6UhMu49ThzDC1+/ohYUwLAUTQcK4tj0e58HoSXhlSdQHFa6rd85u6fH9fv1xdziG4
RLDC9kX8pYqel82zsQ0yRyHpBaBas30H14ApvNLmjUyJMoviRIVXOoFsD1oY42mQamTyc4mULjhO
ZBQcSntcXbqrF3RxIMwC7pbj8FEWtnICJ3jFPLiDMztNEotuYvKtqD5uk5rOFzdEGsRJrdvBKGdi
6DJiMOkV2WpJaqQrjqPfWE3cGaBDwVrG+dWSVNG2F6mQJ0T8o3GUEsuJLk1DVig2G4tdun0kEjGO
cM8oaAmW9NN+jUgyD6H2cPn2zGC6Xkq3oCHxmEAU9HmrOESAK6ruVy6WQbxBZevVUbOj/7/iY4g1
oldQ0fL8dfAjPgV8A362bKChZW4ZI3OE/fRQ96WMX2fpktV0/F05t+yLkU4c8ABjY5A4uRtQjeev
1/SUijVzNs18Z5s0fdLgPhDkbxv0TZ8crsrEBTyDCDxyjxkSEckLTpg9O3gZaWD71j0xWFISsUd1
rDErL/lAHpNLtoA9xEeHGmcO5r0dwizFfV6ENN2CgEDXXdh0FRHJz0osSgKII5B70qTsfVikFsH1
jsttdQTVS9e1bLbbKBveaS5Jikrb75kaVjZK5xqoEJz5En934gT1guh6t8kg5vSem/8sCeOB3w6C
gNWbaSuCDn0F1fkzYNVAvcamYKsTMcjgcHA8r8boQs3ksM6ooeMfRJ2Nsyh/T+P8ttOkKto/8Ren
+4dPvgofGX+eA+iFtA2v1YVprYSvo6X6g0j9SzixzXCNsqir5ajxd8W0FGuxovZNF8idnAWfdCYM
wgsuVb1LIf3oSUm3N7F97LTxC/ZnMENedXoP0G6sRkzkTlEAt0P8fHN+BW7AMdraVa1OGqMcsanN
hJ3XpZPJEZgo3fz11TWzFC4GIR/v8ZcI8/VOlEjLVg9fTppJj43TcrusuAa7IeuAGPJzUal+f8ed
37dYMsl40FbtJG8FvVSBVl520Lb37qrlyDkY2REwTShBpF2nQ1meSdoTaL7N9JIftbEOPOEw0Csk
K+RSxEgW9pshQggeYtuydyM8oXWfNK/+9rAy16+My5kp0qvaIAU0Eyhl5ybZmieIZP32IKNYyFCH
j2CD+hGfJsK5PW7lAdtElo2aDEA2fRjc0+X+WsC8tY/PSvX7SR7BqmLh3JRh9WqQ4hhGRzbgF8sd
WCjtufUpwgnreErCK7n/3e9MrwuwbXs8iFZdW10QepDrI2eqOWTHEjmtVXDpuarOYZRKjf2E4Fi+
L8rKepXTzj3Lv1dWk+rMmcaoanZ+5VmsVGDPq61d7VDqGLNJdVDiEm983nX/egLSCo/ElQCZ2P2H
bq3pNCEmF5/t+EYhf1XiJDVdITEBL72X8TEVb8VN5VZ0X5HEGVB/QQmDKCKf5o8SS+9UxoanCW+/
77M/dGeDSeLJLJaZn+ExBRsC5Funsycmf1XvOr0NGmroCyZzYAD30EbFt+YWpaB6w6e9Wnk3fqH5
NNVm/jEmi70VXX/2XVBYA8fcVXdYosLJEJ4/6iTXQcpaOGOoxW9cfa6AkEzrZAhMFbOh7naLV6LN
O1+IBPegMSPBP/K2kt3A0J9g4TauZ4yGcTeV7J2NO0Rx92ftvajF15WbQWHSc2JUSC1UvgTmx8X5
RsfF91QRU/i0iBl2BG2gjrpf9gQqAw0YM0c98ssA2REG5lnAanySJcqknAaHiDhE2lzPRZ1w8Bbk
SnSvSmMX8rRGDaIZhKIg2OCDxzDayCipce0kwY7Giox3fKzAZdhe3k+mAVgqD3c2zBIXDFsjTloU
wvo2lalM5tdJITEMgldBdlBhMdwO/3Xm+uUdsHDgH3ZV5iVpHV/N0MnQSbkxesls502TwanO5QVA
PZicaCTikGVaXE3ov5KSy+whXo7AEVwnV/kw9/nboWb4UyS2eVoX8+HIh2d7mwclxuZgPR5kXYt3
r/YCRUZeYm2zfqRqY1aGoQK+C9v7EcMGUvFfWJmTNcNsYqOlqK0SAAAOs8kDgYv0ykUU7PwIE3xP
KV0JrwsrA763uLp2peYJuE1ww+lNTIDD66mc2/Z3R9TIeGI4eh0CUDKhcMxm47mO2okhhE1qBnLu
xmExn070qcF4uWjqN00LyxMODOe95mfs9T0VPHCVgVBfnx1SgJYu6DMX9qgmxaBfeJcfV6smS/M7
YNSywd2xl6+BekXE1A8IfimODWKT4xgeqUTH05u6+FE8IltqaSHFox1RV5JNyDOTJDmzF0/IFBc4
+WwTIlaXKm4A7xnkWRunZxZ/+V6wMc510HNnClC0p3cMST2JEEWn1luzaWwZDnRs4hFTOt9hNK9+
WqGf/X9Iijwm4j90XMqQ7cPpOtGdF5ymqp8sDQ3fjnNy/uenIr61BAwNqtya9k4bQ0Qp85rV0Zdw
t7QgoaJLtV2LVqVroEZDUp/pR7q3uFeSwszRDmWj/1uyZuLWEyQcoIOBMx8dgwmA0+D+/PktqQy0
QkygJwNlnGFvCa525Vw+1ESQPcyHI777389jUMVYcszLAUbUf1s1J72O74J2g9fZU8zYixuks0ug
YmdAcBJijJXgz4b0X2trm3wYMMBOaoy4V9PYAf2w/4M4139MGJ2Fi+DCp4oABUG8rf5L+rjBy0dU
mKFA/BNW2wwrNVteRFMirG53QxEHZc3KhdMEsyEu9JXCbkdT4q72J5KLr0bW+C6t4aO2JlqmnY3E
1zFQIXDw5UQzuh8ONqkL9HNBj7ooCBCQEPAr1qa/YcrHbXrHheglVP1hlKVEjwczhRNUhGd7hylF
HNeVM37r5/TwE0jklKovjOQQ0g8DZosnLVHZhDysjwjoMrmjeZVbMcFB+avPvbJ3uyWVD4LyAGTj
hDt1DWXl7m9ufKprzPPptugZgRkAE0ZBG3mbzEAlVfQmf87zA2iLAVlDABhGDp+1Itm++v+4Zq35
NAxzVOjzs7vkwTLsVFsTfWkLV6ELmZbOtgqZO9exc5Pqi8hpA4BJXaB5GQAUYNNdKTiZZNM7Cv77
MdlZNEC5isHtP4qJTEmTlalRbJFpg2Wge14R07KUJ75tZsE+nRYKJrO/1GAR3svPYYCiP901tOwi
w5r4OcEP5UwqdyEWlxlUa9m5yEfYWhUqfE7RK1e/DsgMJZKyU/nSRz1ifNQPqW7SkMJ23hkGc1TD
dHylqP7TtOsazMwYC+eoX2t+bAbEdEfHUIvdXdIxEgnMH/sBENNijxYK0VjRYMn4BE+awj2dosc+
x5S0la8bYk2dR7HZHCN/OYYd64r+CX35alrySuPkoebT+ixKCU5tSEHL1wDThS1MGw9nS+fOgwOT
EQ32yA9hzpdBZXtOPeySZJz9Sf3/wUMQdHGnCn/LxO1pi55j0GhbPP+Vsw5KhuYnyuz3lATH5u+J
DWFmP0obiIg1uYrEhmRs9DesRo64ivPZf0Zx+wDSBypUIMfukrVxPxN5B6ruZN+imUBSqE+ZPkB0
00qm5Z+CA+/hTl5ypIfj6CZ0wcEiQn11YRYv9hyc6FfEkB3XoUCRXYzc2N2YYyCVKMXzLyyzvkju
B1wRGxbLH3Lp5vhptotGX4m6IwB5pMqf45t8NCFEJaingADBe5IkMSbRRZT/yoAotA+E/7EpDR5/
EQe/ZRrHJYNXnMQQLORgCJZVyeLclPtbeq+iRFeIuCNxViNYeo/0tZtcCEesvKb3x54sUvmNecTh
19kus2FrUhD7IgEQyIawxdTCp0xLOXEhPO3Ai6uTebdm5iHE+wV9LuhABaVH5t3MP5N1geZvrW+0
BrAZgj4hxtzLYDDRepBQ19XBt1b0aydpTGQKmsYkFgxX19wPIc52MG9JhocWgwkX8+JUKcabQ78i
A7ZErjzeA/9j/SY0Dla0yWXHRNboFgPK1k83KqVkscCf9XaEKD85r+wLuHaLTka5Y/OID7zsH65y
2uoKdB60YEB/oZVpQKIR+0hiI5AHlXitDr3A4h/SZXiFlFzNmvTRfFwQvOEje1i8q4Ybj6q7XqGt
9OSAV5PjSYxbI/DlY9lwmhSsB1qBSRas4Mh9cAQQKngP8ve/5e3BHOciXKp4wbTT41V/XeS6Yt/W
hKdI8t1RnPsklifIkUjtYQhrf4TO649wt8L9qxsrT/P+SGsify0MlGdGz+K2ykRgEcQ0n8jwF5fH
zNU4SIupY8QQ8R/f3/HeDX/LoyYqof/DeXei5SeGHUsn213yJ2kWqjyM7GWqzML0aKT608XAOip+
uJxoLYQxUE3q4PdwsOGFckkjgVbO0+uiy5NStb+F9/mQywMKzTn/bo5fU65CfSnSUuqsVxcgHwVu
s+dnErO7TGTE+i7FSg8+8JLHZZps1NM7RY5DJMirM9qTetZdUsgXmTdcZRMXr2E85MXFfPqeLsKX
SxCiwQJ8lENvw/MJCKmi4/sX8jLeAtCG0KwnmVAVBPIOgMMkttWZrtTg1hfesDI0kxmj6D+npaSo
ZDk9+kbCgrKrUGo9nw8P1d59v73o/wgsUqoYYJZ5zVLfdTwCAKpeNtMbr83/emYGdKHBTy/IKvLP
pzhMxQMFgIlQd76b+tUH9S+Om38xg2nWFwrYWfFwL2KTuiNfbYTbfRa3vCcl4Ns3xxpIOb14Dzk1
quzWYHTQCqmLq3t5v30dOZ9ijD8CBxomLqRk7RyobW+5+atMz6f+bZEfs7prYNVSmvz7sKs1J/6L
FU3H/VH42BjdcR/Pkaw4+2tJW3oq6J9TkCVYevYSZaLhk2zN21M6WBOZwgdtXVBBHg6ajO20kETA
NRt/Yj5ssCAExXXkc0xmheSlnTf6/4LhrsNl36Bhz8vbZyq6BDWYyT8/xfIJl018PUgBQ7ANM/kU
2wVztmayIDmeo2Dc+0RVd6lR8TBRXfs2t8pSff7KfgSf3RP3xO/0GcRi2zMmfdfcpBSRrHc2tWDP
/hmlSxSN3Jr4Wx0JCcvbjJRaaLp4qCo1+4CPKvNo1OPKcPbzVRuvImmEViKwv24yS9VPCHEu3AF+
mLwcuaHyeTh13PC8xWoZkBPIPht5zXHVzmbeyK60Y/4xcLCDc6Nd2eSjnvBrK/LHU8Gaa1EwnKKD
M9W/fuRSBz0oByyl9/U8gWtT4h3Nu8PyOMGIGc6WudQzY77l1uOKJe7hi6ZWHtSDtC2gmS5e+wOm
NSA6SpHCkhX4j4vdv1lR8O5gATblOBzTjFgTjUf4pfMACTcvs/9PE7TKntJiPhj7kA5iaEtUfyKJ
ZOLNwldLLIxS5EI+/MrF2gpjAwlc6jMEj5LBAprAth3j5kCaPx68vpZ3NV/cDk4+aYm0S77bPZe/
CGwaH+h63H4XhKZlgtu4b9oboMEe4qhDtpsl2DKC7PddBLAx+RvvN1Qm27Lba76gnPNHaIXq6oLA
NQN84WLCPc36ZUkRurNGCnNxCXOSS0atzyogCPwNo0SWsRWvQW23+425NhbKCMb5jB3+40RcoCTT
NH5DAV9DKoGOuioZssFDgH368P6UL3K7f1UhbYlTqpYyg3AMrY2W9EFUzc3gC8R8k1itDmq4PwIx
2wZ1eYRraEFur5H/zf7l9sg7M2pRnSNAQ6+oOV+3X3RPOCpIw+LDPSbKXhHyNz4kZsze3Cx7+Fou
/dfKjf0giSBCrOtpkVL0Eg8B56T0GSiMRBUHNKIK8Bn5ChQFj2tAihztdJVNm0/EH+U/8ZW6m3/I
wHA8g16qvJGLv2/hVW9mNwtdoRdkN/0nBVPVoI0rt3WVcXSMOAU7SZ/eRCnwm/GLjUqh1K8X7jP8
Zrznw25wHsrU00OkGISxuyS3LZb4uXikXeOzra3fQcyCoVagkXdFcu/CE04sB49qEf/9XQrKgKUx
68r0dW37lH2Pp7c22Bh18SkuM+Q+Dwn411WMsHzfgIsD73KC//V1qd0Xn3KkPhiaPDMRHXIsfEas
1zlmWZD25/WxzMqPHENgUmTEhJfCb4VDo+Lth4zGoR/u3ANpY0GhMDY6FTeKW1GqwU32vCMFT4Nq
wvxhkR5izwQyqAsaIgEXgla83eLzGQc3MVYLi+6UCRFc/tJozOtlMIgCpN+ExPCiQFxDJgHCkoda
yhrYdLQ/yVJwa6NRA/lMvlO3wMwt9WdDTUay/v4ueZwrjgMmf8ADwmGN9KhW1YvtO+sVdn6t8uMJ
5wm3LVHVzZ4AnyCEiqO1h5iztT1ZLEkm3m3ZScAKfq26eoMdqxTOwSln6qWBJCNoeEAL16ZLLlkd
ecdOm6woCgxIT5nZZGbkB7ikXvy1eTKleLvdis+sTTmWREpPkeE84Rm+L/5jJeuBDeAFqBLczzcw
6dLZ89/LG/7kgZfCVw30ko2495rcHlUSbl8VKPNeI12HVjDraMIf4dfMrU/hXs9J6r5XoKH/NfYx
2QMKYmKQHqiWMpyqIQMJk5iXNuhI86kLMD4hQ8Nf4i7VvXEub91nX1I4Y7DURbceDvRd9VZUuPKF
1XH5wNlbmcv1NHVt9DYa6Cg2QkonjhnKVNmyP3xMzQQ0iP4kgTSRVhd7Vd1GH3BhgJwww7zWtA4/
48Zl1ZBlOQfssMxomPfvEK301XgzOqZYVQdPtRXliRAH/wyQr0Xa42xBldES5Cvk9bhx5vJtzmvG
TygNFvDTQE4YJM4mzgfskbg0FU2L+7SiUOOPvg+zGtL3JmVZnbtWed2r3z5KPxkbpfioW1Ff9uFt
y63vD2WOJbvkl85RhqGRFjl5Uc+p9FoP96eGV20LUEk1UAmRSPdWcE3sT3XnsCOoH+GhHVfYKSH5
N8KV5jk0tYKf9CHlOqyaSNGWISVWeDLVQjkU6nLZJXNkAXKantTJMlWuLpbTJtgljooVTANfU0xF
++U6vl+ANFQ+YgJngoVM7da18H7jStbNDzSYLQWz+nV0fMbwqlVE1mOUoiYhkoBEw6C9aa6yZ0ny
/h7+ZWl3nhpBUdmsLJWFpCJJwEFD5zV2xbxP/fWsKl8WCS7DRbKrTpbPlXssDACq8WKMtgUCx5mm
yDFI/f771vW5PdwUIThIcj7y/6iud4HKcFEvA9FTKwj4kjI4AdjdGei7WNkmfnOcbTzpZDsGhJRT
nltaBpvUZIlzo7eig81VhMaRf6/WZD5ruebNmuYXeegW1JhO90VSWuuKqwKCzfLLbBu8MVP+JIMR
IfGQC7ZkwVwmZx1QlHVdnagvqx+JyA2jR+SL/NC6iaFwiuXQJPbW3eUozwz2rgAX15tmqLjevl9a
rFjE1QqaalfkhAXdJNkI4pFWvJCIwxmpefwq6Mhu7ARWwtZ2QghZww+q2aVFXA5o0+juOYMMXIlm
6JEjZ2m9vjoviBimLWH5FBJ5r37I6ye3dXj1dUJukJbFeb0ju1VutnpXnBoKxEhI3l/EmfSKiCL0
R+VR1f5rfx2QiFirE7ocJFV50Vc9kChIofYLI7BvixiT3s7j0EpBoO+XfYYJRVV88vi04WFdLhHL
ldvVvvuWnJhCjfRYuIYaVF+jKxTjBYJsw7EpRo8lBhF8Wy47pH8y8VqdjoJu9CFQyJAQC+wQlCyp
5wMtc2Ycu1Zb50VZdNVjZgsD4lU9mAyzc+w0zPLbgMgPWviVLxXmk/lSKtLP8A5R6oSXEidsjHqk
s17E8J2J+m11haVxbjKoELYKPrTZUVvMid1Uud6KEOFw61XO6SeiqFDWiA5RnztPV6gjFFLgTesX
cwgj/RzxpsNJV85yD7JbtQ50opo7LtOtzSZryE8nxu9mXZMzw2JCUj4JFc+nPIhde1DIjpEhvezk
RBMywf85pVFb6QKtK3FWMdkKwGJpOd+6Z59Okp5QP5YRo55G+u8ejP5Y2s+65/Q4cCLoSlMpSIuI
mgN4b5u3Lgb8xObUzbNWlV5D095BCEErryzuRukLs+ld7Lil9FSWvLc5ABj0WJPChYKHAdEz/lq5
TxNrwwzdMTzGZ07NVDDjliK+/KEyDP+Z27REQHFJLptZ4ml2g+PjoawLFrR7GG6zZfcQa/EHJGnt
jreB4grI/Vzl45oXoXzSKsp7HjHrklQ1Mypd6UN8uDQOoWA7/PeZgMp/U+JYVweDJEay3uHOUivW
vFOej5WpvSom4QQ3l5oGlTK6ivQ7/i4xPGF4Ntz8xeoxoYkjc0E/02TUvdwUU1IwsGiK/MXKncL/
0X1BkpkmF22hUMZtDRZKO4K3q1Wf0nyYn+jfC7pqaGh/QvO3JiQQbJAWeudInfiRE+KddZypOtsW
xhuHeCFcrI1n86Agnah7MocdiUq6ObkedM7B56Upip96wNElOUG0kJyh6LXhO06gTBPf+/m3w+HV
X79lcbsr4fzb4d4nbg1bAC5uv3dg3WA6njfmsgvoUdevawrlpw13mTMXznN1EsyEnlYDhwdmsLq0
e8V+bj7dWcddU8xFBhUJ7sT9smuKtaohSQlwgKme/1ZPQcT8HWCZHknGOAsaWXuPpApfK+aUIha6
Pwk66HOnRgURPMEebue2GkM2pHk1lC4kETRBu9Fsv28j4liYOAS2GpMF5Qwj2FVoocTdppSOBD4+
SHE+RxBfJOk//7zv6ZD/txm15IKCrolE4dFs1HNBJ38c6N3KO10kiRPka871VriKSuYB7f33B9rv
xw9Kx9K7zALicZ2wtIoo3HJ6QTx7wKkvXRSkCRhAlgXH4dfCv+Tleg4hGlhAYVdZXxpQ2QF4zcDH
xC4mF8eeF1NJDuO1WoRPXidIqKEG1AdB0WLaPDHFhwzqf07u88sGbUrmFkDBdiyGV624z2dO3KYK
mwGto5e1pc1OyOFWt9riHM/WiaDMubwJs4gGz39Ul18mTnu4UPYS/mBP9eSkz7sckEQtvLoPiUcF
ahi+G3rb9QVs1MY3FOJyC9nafjK4z81RfoRwe8L0RLzRL/NfEcSwhStT/+lMrXWCdBkrguhDkXn6
qWRjAAxvapeCmvJ1l1y+Np5f6cf5y7oKVLdoD70DTX7k5c7NlFFRXl5CMI7KgEG/emIiuWVdkO+1
Xe1IK8laadKEnSjqSAGa3m1bpvHrNYgZqhForjiuDMNDVQ78wgNUuQxjZvXAhupMZV6bWXogbeyu
AXa4qslATI/MShA6mlt+H+8LdZMekjJUT0MNGHH8STpm2hESDzkKGDVsL90e1/9YU2EVxGPg8cMr
9SrUWLGBYl4VrnF+6rH2IcdPvIjnZ2aq+hEeYFuJGILTJuk8NmrRASDdV02za+hQj6XmvOOuJU5e
OsHhbkUfFJqfJtqDif3JhMuGMgAc8wLxJW6ldBcfXECHszOfxl4n306Y5/o8/6P3sZi4tXewRaSn
a0ZnW5+JK0m/GHrLXiJsRzg1rE3aN7Q1fWTVoRGYZeEFmg5uONCGrAp2lYACXJ+Yojl8+HeU2/8U
ylaJe3CLzklGPIFRzhnNHx5mmYOGz2JStvDDuYEm1yLma6loEeR2CUVNY6kFmcKBSdZQ0q0kda3H
kDvuS3NDdpFJ5oceWZcY1SiGBSb/oaE9nJpzxxW/CIwIqAvRA7T9kRaCp5w1zoYZjnpyyZ3l/ztV
gTxlZQIofezcKsmX0Dc4AXYpVhlGqI3N1BvI6Bh4yHUhF4U2qUKqgHql4FyFycMnLq40zhhAGFG1
Q18QRqKz4u4H9Dsj1sX/ikA411SIWU6mM0vHJiRhGqQIQ4xjdKr7IyA2JutoMszHF5B0zGNkNAQM
sENV3+olnznfBs0D0oBdjOYO+vNyY6teXDh6/UiXu6plYaQTPD/SsaVr3yyZgOM7F4EhVU633noy
bP24mEkVBWqCno9GOTt65UqyWIaExwUvAGRF5fjZl5OTQno94U0BLkgCWqiE2DBtBHDVm0ygIPGz
623o9e8BCwg9rNSPKfxcB8FKNEhxNn2Q59qn7GHJENL3Aj0Yt8dtkvVWYrQK5kVoGpPZJzODPnUn
1t+ZTg1uJVzb6fuvM1hMnsRwh6b5YIFbuYcnLl8j2rjC3rWLrNfqqZxDm0MQRaWTmtpN6oy0HNPh
1yBuBUYwBHYwuJb3KRRttVoAk7mTkuCYSqV/9gJs2PmvbSuyoYEOmzwZuPOF7KnZ3S7yf4I7Eh4q
VhEFTX3Ao0g2efRPfgLENtn9Gm/UL3UvHEd3EQnH/VS8/Ktzrj4uzB3NswpsB71xn5Cdw2ViFs44
l9B8bD60jnrftw02uRwUPwuqltIoPrUmlO/WiwcmJin2GPQFggmKlOPEHH2g7Mx1M60+DnLlKiQC
gJKHDUFmw+oHEcs3lP+v8FdWLbexQoElnOqHXyTo2DcGhoVqY+BmavbRSDeNOi9IiZGa77MZENvO
RZXrkxHWN78k0CGcq1a5FE3oTFTv6oaW8UqI4uzABNaIx5MIgLn+h/lSzq7vUHlkCe3LRm2YeYMu
Cm+o/MF/aS0ky1FwdeLD/Jz6KeUvLJLklh6/XhNIonArcnKisqStWR2pGofnRgnR+oRhZJ9SDs58
XJBqQj+AExbkYW67z2RfjvC+TCfX/kM3e7/swCRsBEgBxzJhTWYLbHf5emaJFv0kQADy1nZ26otV
aGyqaQSXQf0PNaj92iuylSD2dv0YSvlv+zw9CvO8sDupajbE6lPVjj0dtL9ffIl+7+foMLe1DMn/
N6fJaIzJafHuIJfXeeXaQJl2gxtrNSRZyKuSTHQbpVoVi0ILLbuLfbLXl32qUkfh+7SGpTGq5gPj
ufeFlKPZktPbqZuckgprVavU27tBUqoWNxewVSdMa7Rz84Ebad+ZXKuTe1O0We7lYmemvXm/Mgs/
GxZyLwVnk0ToPgHgM361RgwVBXqsWCwRZBqQ++8U0m3gIVSQ6bqC9s8SvuPlQD1ixHcRqGupERWs
Xxu1VawUwcg1bv3J6S5p2OjsgGWasS14u9YnlCsRUccSa5nEKiZWPdNTFzObn5lR9Zo43f/mUY+x
OaHzIwEbHjvSDBKT1WxBPB8lYYxIjLabpkL8xVr7qfxt+s5frc6JGsBjkrwWhuVJ0uUQGV8jZGwl
0dVU3MOvLr1DLFc4G29NkWzMm9SaSmR/CxGLfAlUuZ/58WXxq18mavPUOIIoJSODkCzSp70biUD/
r/byciqhkSUhHcBfIymsG+mJH3FtLC0C9+CzmOluxvw2lLyh0etAiS38VywtkxVxPGfqtCgrOSh8
s3pnfdGo4w0elD8IUhMeckcnHsB7Wkwstcv9n0XT5lSUbPciQ2c8ORVADIKq6b0U1bCyD2K9kYdS
C7XB/84Evoq6C/xYh4yWvQ9Sqb5jilxAlPkl5ewbCUM9m0KvaHGpYqwNP4p87Zn/fdKNopwiKMTl
705B0DxGEwfZbl8Gd/SwhIJ3Q7C7huJJv+yrwLjAhO1ZjdVEM9JkbKEMLGIRrl1gujw48n6enwNG
MKH7llx0kvXPdIG+i3NRUGTZEUxewEY9kYyyA/iedw16xxAdnY6Npbz3n0hG9eYyWhi47zBxNn4T
Mnqn3YSuYwKbDwYgtDH2/P7cR09l4yofRi2Ej8x2JoWaOZjAn92DoDvCV0qOk8YAsX05M5mqdWA3
a4IGCJUx5KxZis1kU77POIDZq2S7pZMFDC9hp70VM4jdfpu+p5l4gpQkGVmzgyqz4uu2LVx2F2dR
p+FH9so4e7K2JoP1R6Dr4CrFZfI3Nv7K+y0V9HzdJeMRhBD3AaX6B9Q8aK9piDVsZU/yE2LZqmw9
9VzZcknBm01Gh34rKssvYRw7j01W0CupAp1a7s1/w+S6fJpexJ5ZP+bxDAjQxr8BEvaZziFao9Pv
5ZrISfBybh4/HQ2nyXUASUrudyQ39ArmwkO0+3jG0N8L06G7flBcluf8UENPpPYZN2WiKI0M5H9Y
Xszj818o9kLcJxdrnbgfOTaxD3EycGGo9MXA0jC6UCbgr3t5viquWa013ixwOVPklG7UGG3MWnKX
UkfZyhEz85T+EMFRzOMb9Tjkj9PvKS70Na4haTbG8KXz1KhxFRkdL193LcTk8lQOJljjEzfVff2o
EP54KrEeR9xyUKMeoNd8YVjBuwgdAxiK28GGHLgDoy8ytdxaPSGdEpU6i2HhIu5A0vQyhfoNnZQN
INzno9wFyyPkw2sTzkVI/Z1LL4pnRqQE2QwVdJnksI0vsikfZrJw/XQ73QrzuVqCV8MRLONsM7z2
S5M/Ah6Sm+v1x1qzguPKSKOQ0PDJnq1kTJLjXCOImq2zd27oSZ1CldDdOckMb6lW72Q0nsRP/1fE
W6Aig+kkqhH/eneV4cZLoSdlpACAzPYQbXG0r/tB3EuWAxYLH6Ji3PynBBp2bmAVnjAKmNqiIMUA
IPmzzILVQEtVdI1RtB/CT/qJjzH9WhGg8y8YSdu4OiVrycJSEZ3B2+DArU5CfvkZFE1ArK2+gJSN
NOlWc8fXJi2VEKI8IMWTHMPvd/S0jcrP/4DUJi9q7mTrRC4Z72kWptJuNcFr++nly954F92vSSh4
hLbhmuSWQFm+7h5Y0N7Lg5cMABoEDAyH+vmPYR2MBlYCwK8V6+ayQkgyx0PJPpdN0GxK2YYT4ILK
mT6k5myY1cJjsGEWNDsh3UYr+YO9l484xxpoNaVE+u8mS/u3EA0Vlobu21ZkWv3H+ZlZboe0030a
tfJf+HfoSawzrN/DHW2KzzVZyKbnc3uXGBlQWv7PmgMLlm/za8cuAIxxWCb0QcFlmdsEGFSoTclM
8XzDzdcxJX8EiTEc4uRYD0edRpHdedkG5ZgYWXStxvd9GGN4hTYwwGUsbh5b94nWTYEX392LxZu6
fF+hAmgwjDyhU7vnflMlS8Bzuz1TAeDs5VqJ9SuR9UGwB959fgcNF77snp+ioOcOlf/Acw1kaEUs
TBaLv7ApGJ/OMR7tHSB4xDv8D/+s9ZIVlOyC9Q6dDiFtqlLK/75eaBCwNVV72U3UOPLmWPXO2UTe
I16er3ralexZNCQDTe5C0qF2NTM8KIqhjITDmWZz4aCtEzDPcm16US5LrlMn5e9pNOgRZ2k14HRS
+ZOk2FtGiyxJ+NPEHG7E4NS5rWEjazLyJqXg3y5zdp6jWAeI/tivbx28Oo00omwV9krj3ITzvsUd
RnNr8nxAg4fjOQMsO0FaBWu+skDkDYGQfC07CN3ieZgSfv+kVHC8rQr1xn7KX5rQt+Znn/NrTIo7
RGnl3hhV5prHBhX3AXj7gKmP0qr/YUd3f894wGj0aN4k/WPLF6cjE+xNp6nioud5WSJ5CThjWnzI
NJRYR5kieKzSeT5SowN9XAmgXzKDGPrjVjnr/pVo3A6kXpAJ2y+9LEey9MDeWbT07W4XzEnh1lnO
guiJ0Jo8eHXchygMuW0cuoudZq3MQpITyL7wRXcFDPioT+/fNo6jRWn1RRqHS4X2qjLYo8HUXmMY
imdDUE2MtGT0jXnTDS3MoNOuMma6zP9hnYm+4YZ/HlzvZDMtCRAkCBuVOP/TlJ9HleaDdjtd9ATj
gQD6pyxN+43vrAsdI0VLXWJKedUZ3qDs+uX2glMRJxVPUCoShKQMIJxa171m7z7W9RancyVVxD3N
KZyWseh0zvdvj/yA9EXI1s5haTILc0PYTvhm16q9L7gPz4OgQq9LZ6e6RV3yfSi06qJuwGyaxKQq
/L+6zffSjYaukFI25r1tytBon+Cy4t3qzvDcUlCisZycXdH1UcOaYdRJISV6x845+XlBWdJCkBz8
1IbnLl9HY+6JVrzS6Pa2XYDcgW1fNs67LgeZTwE7KdDfUkh9zNr+LF2c2jQW9fb+Er+YHP2RSLSU
1A4i58et7utR+fDTJnPl3tnVcohuLgGqs7PTRHDgBgqANhbrL1TDY3ifxFh0+9R5ielzFYQ/lZm2
lzNMXJGBakuOHDigbzqYyuI3eKR5BHKHDRCPmGaeKdKcoGVhxUklRsiaX1+fEx3Y27rajdaias1Z
vJE6GFFV1MS1uB6EYeJDjMSRYoGutPcwMHrmyIdgpYd7zFtHfG8+HNo1XPr5hunBteXXhjBWVb+N
DhADvT8h8f6yqzRLgMO8jVlmkMqxAEk3zRkbCZiqcbHw/uD0R6AaLVzlM8iDKmcBCd61Z5234KZD
TZGcIrzlVg6lm4gwWae1RNQMhxWTaI7CIuCs8xfwhPuxh8QBqSb8GMn5jVBmrJJ2P25vYOG6buw0
bTtXiDyty++HGSWn0ZlPlbKwZd5Ki5bLl5NoZRoVgNF4ki0skwTBHuSpBdB/xqyAUUpgt7A0UAve
WKub0EDFCBEjszvhzcV7RMmoHxD2kc5vLowfMzaHRSRhLStWaeDzzeRJ/d0mdpQNE+f9bTCqBzzI
5gtaWqxzz487lxgcXkjYCH/r7pkn8wQ4ZJPRjTavQXNgUwhHr3PG7uAzUrUcAUFIPw4K0xWwK1kE
PoxBglsTeoz9MnlBPvUWEhnKMae1JAjuJFyBSaKufma9eECMW+JNyJCkUXZiCmTMQI2ywId8ETol
zE9ya7oBUlMAmMF2kIdGWkDhHckgCA48g/FDmYYTBqnjoitK0H8ubdjwdjyIVv7ekOI2lRNbEt4b
P/4yJve0o/bV6kdHrpAlZuxWg5kOynSqlJWxKTR32aXqtqUZb3Ia2ZVhkiJwyXKPw3LTdy4wwH3O
lpITKj2H/NtTV7rn4R1zs2gVc3afNZ85Xtmwj+Rkm7xhVqGd/sAjc4G4DpfrkIhJzXUTDeXkrWam
qLhjZmAoa8FOTLUrPIZaj3WRoLBBmHvVYUmgjppoHFK0Bqy/WdMjzrXvwv0B/JVvegcaPS0t9Bqy
tjbyKK5vW5kTdQuNPbXUuIbv6tbW9rMI7z0s8s/ewztpf8gkD9kHqVLJbtHLfksMfXL2B5CYw0V9
6/lJsvz7LvUf5z9S/qMDoOFfzX8O4QOkyM+ETKqV7GASv+wKCRA5D6/AuzAWVapdkOQkZG0rTWVU
OvHZAryoXNap6+pr105x+8rXpq5iuomnAdsMMs4jWX1qohiVIaq9pVJltceQ32jl+/qaTz++cXR4
wdiorPbQR/r8KtndFrbXBYhIEm47zse0FPCLBK/AmH4lebtB3Win/7cw+I3wNXQi6dv57VCfvIxK
2NZpD+Q6Gv0DKnF/LOrzMgiz8mIeJYlPDXxOPu/hljxwEo6z/5pMdNRY3xfUsUHC3otvnJAGG22s
8lV++An63Xa5DK34KOS3KdxE4iazRNpWXJWUZd1Fn32QFrMUqY/iHeTROPh9gSwZ6P32zgot5vwT
Y+O0h4GLjXTqYp3RJwFLt+nwfCSqoWz6AKZf7LWl6J+MgtBycOcgqiDG1b2NFlTTL+m8OrvmzjhO
Cad1+70cn3ab9FJLc6vxpTh7Ru85ow4x7E+BEceZYo5gH/D/gWBLASRUfpkKNXbT8jp0ah4jmnc9
8OGQk2E5t9gfU5b3tJIuJ1Qqf1nh2fVs2YFw6b8kTejL+MpZPwCGdLFHbiRJNTUNrjJplncd0/Hu
8YV5N7yC482Z2pQXLzdCA3JhirdamCsEL9hbqws1QwiN2DWzap8v4bAYNN5J1krmUBULe0YzMFRv
N/aFtwR6/GIB0DU/zhGTYCnS1vZ3+CtABtc9HlojddX69yL7kDiu0yBdnJbwg9uKuZmgikS9UjzB
/WCmHDWa+mK4AEvPUHVx4A4HdKWBEfboqDRsGApRxC9IKAPS3aD6igOoRUGC8p7YpqoZCsqUvqu+
7htzqnxB3To3lPpj70VTvVnfy/SxFlFRXiQERaSn9W0bbOsx4v056f0LOoLYYuw2lisWvv2t2g00
8ilpMXMXQDDRnznEE0KlMYJEHRI4Du4Iew0A4U6dzXBVeiNzwo4pUYupkVPakjjdkULzXYfieH3h
KtyqdaylnKjugDKed9AONSeXOIkhbH5obrdx4g/nNzrtvpKVJM7tfZ1xR/p4s9n8QRdgzyLDXn71
7gda8A8q6Xg3tTtf0kcc/c0Qn/su/u7JJf/GLHz3bH0FyQH+P+PWTBPu/T6OzJ42sOz3zfRysSFf
86ZiDDeui44N9OldMpgKIjBVZ8KafEZAAO7HI0Eib9D0LjM3+oMOEWB2cWsa9xubNKuWYqSsBDTI
dvHBUUWGNjDRpI7A97X6/Pw8zCcxsZMt/gTIGEQx/8f68tM0arafCmyWoVl23tX8XWPveI8Q/GCQ
Pd2yBYsnoLUpqWQtEyBgvv/4VvoF2/u4E2U4TosmMKjedujgtbKTab0tol8s3Xjg86Addc9MxdU+
LJxFj/YR316S4wicX5CLg9VYNNPdohqeBNxSctVlBhXVHXrpYV605YQjvR97vN3yQIYN+u+vqqXv
gVdCDP9O9Lu382lN/t8hun7N9+Ee0gyPq+RbJHaduD3BySbnTeymv822mOq11/l3i4M9W4GWCEA1
dddj2BdQlKm+iQOmVgKnPtoFzm7AGRH0Qi2m9SWlivUIfjaPCRB9JY2JNqf5WnFI04rlKTrGRol8
8y9SxZgVk6XHeLg1vpV5Eu6f3uW9/uc85T3sQCUOtwxOuzPR34gE5EYcN9vGj0agmhSa3TuHvBha
TGj/lEY3ZwyE0tlDwETvBvRqBB0pzx2Dz8LAq0gXDFhtwrJ9IEcUw6v6pS0qHaGvPOOUe98kklUN
xQMNeLJioj7gBKWMBSOgX7hnrsHCzWRsv0YQh1w/8p7d7/JCtxLwuIeNI/HR7HQnDJdf/Oh4SNfJ
enH230+TfgGAnIuIEfYTT8ojaoh9aTuNBZevHp2XyI3t1s3cMDiYqya/U7L1VmCWe0StpOfpLF9+
tzymaRn+rN/LA0R8IOz1bWypsCk+y8LYnIqpyrxCQM9ov9ER1lSfitutsFa6GKEV9kAVES+SyKj3
q7/YBTnUu2xvyjGXd1GS5FRpbiN9fP9DnNyF0k/aVnQzJv0+9QsrDzNFtR9f6lXqh92yLwj1+TUi
zTlLgfxK8GmzUoqbxNPm/crNuuJpNO2OLvxZcaONqaBsc7Zk13+7+CYUY3n+REMSvbREEUDBhOSi
6XZ2w7XIq71Py+uwMI8Gd48WZky8t4YA4jtEfCCyUl8tnNw3Kgj3PUMhdYS2VsWQkC54swYCXanw
uxuXCyLicwo5YQD2G4i8L+agSkIIu+Cy9gGZ7pkl5s+L2pqZp7zv4RztuigGJ1iOwpRFJQPqg1z+
fX9NmCev3vJkNJdDGUPLVXqjZXt6kfACjSF7aL/qNKVJgmZtrC+daNmzRkZBxGRi+zoqGJtCcsga
SRnHw/7KiagCpMrPQT7XNa9Pm3PDYkwYBvF3wjokoZMpOcm0JyOSaW3ZPiVr+P6B33zOiXHcNmeT
N3HAtJkzFAhFncXh8hgYR9uPe1ProIGAKoG6vtpmuBoxO9Jdx8pQt+EloDy3G/TAONmlDPi6Uqc3
/gCOv2aT8cPJAr+zFl0CXimcGRZF4u9yEYhMY+jaUfqtGwIjskr7vWnbj7U1/qLOd3F8xnGCFKE9
L8yq9rni5or5QJbyeRO/peYKV5Dg42EsRN0jMq40CbAOkd0lWHVYFQLUWvWj4u4r/bHjANjVuVOP
qYu91QRgvkyNxAzsxpvwwJvplPYio8A2P1SWySmdCmn1KfR55m/Lfo55KkuK86Efh9JuWG3Dxol+
tL1wNZa0hX/Y78MH59udE6SsQ2YSn+nfIK8OqGzcQuTvDsOyQpg6ZsTKcz260Z6r6Do0j1V8w86+
HF1Dkhoe5hEEZFtAS9Oq50Ev+rav9FnyHTg/L1yK+v/kEO32/5iSyi1qPzzaEH59klAA7D2tmmWs
tKq47x2GNOptsBdEdOv/oosuvPprOIMa8xrtiEwh5uvoEVFXg1r51fujFnqOqSfQNLhnv+fk9NM9
u/3gopcBaYDfLlT80cRfeajyxGyx1J18Ko1G9nYQac0TAD8MVXMflaGOAvpuF3eZpm8eUfPB92+m
80/jKE51Sl78FjnV5kbNpal+/Q9Y/K2yGcfpvB0kpr6DG0K05HP8jik2ceQVUuO8pHz0YWnCzO/D
2cOC7vwhrJ+N9G+kJopwa+hHftlu2Lj76yWMAOH5SvyBFEuBb1oRihu/mtXR28dodj13Lsto3g7q
TcS3thmB1syhcwKq4gf386yyYTDFrduVFUbdmVcjzZ51QHyp0Jj9g6piERqgtBItZHyvUtqj8nqd
sitpumLGGL3+OEqAFmcWx+NQt5E9rKKtx06wfn8lykXo7DYCXaLnR+n3nlEmIrIt87qtfkGWJR0p
P1BscoHhBUN0Ph5bVQv7ORCqBJnwvUJQqV0E+9yseaqlBvDU+6wxxBch5vFev5uWI5IiE92PANAw
/VFothc1qB0p4Grw1tPkppN6jKzE1QvqtmYmucoRP38M+UEtI63ISOcwGd2yvHTvCbTJupapQezq
OrEWiMFDPobjZkS3On3zym+7GIZ7bIdnYWlgN81InzdY//bbvAgUdsLbc9doez4drxXUUZFT2/RD
POHVVu1nPc5aT3EsL5rP+TmjYcp9ifdBShG6tHyVbz0p2Ayzy1bmD2xUGX5oHMt2DfU/u5LNUKmV
6W3IDlvONJrrLW9opnEXBia9ApDLBqh1aChVVnXIBuRm2fny9xoZtq/pWr7VRrqZo5ohPKuupC+w
LftWI/7h0jcYPvXlxw/C3ZZ69aDszBCb6xI6A1NkFo0Ufd0BTjYwVdtz6bpMl+BzCUVNRCnDsRha
9C8ejUx8ATq+AOjR7mT+lcUmRAH3DhhDefm9P1dZTpnCEdI0AiigyPeSfBFcbv8hRM+ijMH8/8Aj
HMA7NoCWeqy7NcRvDyemIDMn9DY+wYEpw4EiHTOARkkC8BQgLqhc6ytYuUhxtcNNIQPoPyy7MQuY
ciyvRDPYoZLSprHEpYEgwhms8aD9ndwotWIKYy2lnOb9+yJLJe29KzxQ43r+336Y7TwM9bRtIZJO
nvu6LGKdV9E+g3c4W2pYD5rYiVltC14X/S4EXqECCzEq+yQH1XMaPna9h/Cisuv0JiYDREbv7SH2
LFfBj0Ltkn5faeFkhMRqun338v62tZ6W7bNJr74k+F6TLFRZuw+STt0t19AQWeFF3Rr0pmfQ27pl
lYZbvPmL1mArpXZwkJoC59cT9HCV7Ycv1h6sZlBya+92G/CRMrsrAGegs+oLy+E9nFXnu0vI/y3Z
TzGONeKDjVcRDjary4v5RFz/kdclTC4hMylX40X5NyOk4/WpgmHVvKNAVMuk33e4pyJrXLZoMvZi
ANUv/j6nLya8hTb0MlsKwDm0yiGdlKAFmR213vVMqXrBiRQhsTxqkpKj3jI9twmHTo/ploVtC4Z8
SuTfoH0mvtU8dgJVQWSf+3AYVq/NIS9NfNSWm1gJ5PABhpS4cyQNv1aNbGZonYsTdW+cn04oPfJj
s1kmxEvGjLLAExvs+7Ui9sEkODXGLNEewWyMlZoC5DyDbV5ADCPp0k6OdQrE5vf1Q3+4EIVOnfQj
AxHKe95k+vCYj9euf7fiwfv89dWucL8GD/W8xrWGGp+EKUPzPe0b1+lk7HI+e98hNo8QRVFOsi6y
s/W9NpJsS7TDWxjMQXZQi3rjGLnPAzxqodU5PrjTUFu3Y+SqFz2e+XsuF4U0jhVIQLA/z4eJCZwE
kvLJd6beQqNhwvOjy80WRl0kH0ozCus9HD57zBtKkZUoXFEOx8VIBXeq8ZrYaQ9LPAqwA49WUF5Z
6duzcTaYlAREBMi1rhjRRp0ujS2U3lzzMPHvZ7FjGuqWcRvFQVMWUKhEGHAcFTFzdFCHBLMhnDlO
wCEwhkvDpzpilEvKxOuUenqnVd9w5xKQtHKVoI+w7iQywyb5HR9yS8TfLsMkS6oZgc2QuufbVZf0
GtVxMZw8OEAg7RSIPmFhhp86psQhKKThHmP6XcqCXZ++2iIF3hYlGsqo6gQuUbFvcU7PtEzdPQ+w
jgCvkOlVAfx0dCG5A0UvwYozn2dBqQZZHOkwHdros6Kh2gj8hikP7QVA55pCetbJzeHbjAQBMdy4
UWQy98iW3na46tSqWXTj9JRTesvNKd8J2x97gMg4cnjxY8R/IL9XnVrB8XcT7/gJTpxUz8lPVSpQ
+fVk0syLHBg6q9P1/gluEORjj4VAZokX42BUWMUBb1mwciMFLT07PIXaofY6Cd61hijQINCLHvsA
cz7OlZQQh0/zbA41IGb3M7i6kZPM3Hs364w4CkoZpyrAvQYhthhBRzapDpUMcptozEy3V2DNSDmo
hS6yg/lyO5XpZAABZiXOAgpCNkKBk8XjhfwhKZKeJhQWgJuyAZ0PIfwJ/X61SGgbMTANLv8Uidvx
YfynLZ4cNmHmf5udf5mh0wpv/ess03I0/C7GE8KAoH3NpCccmObVf0oTQSifaxAceeLju6iqk0c6
myk5hxNIhwZdGBRBci3gVJ4w9WhKRLH0LwjLzaYutbBcPf5VED8KCxxBcsFZqMXbjDXs6rbcVYQJ
wuhe/9HKWbZgDGxAt7iAqHuWloLdsieN3KxWlgaE6vJgReGcIbhvinWwN2v9lPUXsic4By3EIYhw
st+KlZ/BI0dmVcVLeCkCRVKI7UGRVGR5iKfYqt5ps6mKgpnt/yRE53IlDhzQDk+eu8bBoEKei19x
XNM6D/r/2mKH01n2RaVRFCFKoxXY69QbzkLvUuUvRo7iLpfSzK6/b/P/1S2EgKIsyDDDo4IZE0M3
khBdJcGfjZhjyVKH2Zlvjj+2foCE2pKHnypyzDKemsRNdt8DpDGgKcG6vCev4I3ulU/AXm0VlLD1
BohtyHcF58xD8zuTvM29sxzfB90AZhdK+GptNnuMK9KF3Ay7SZhx9oOBHwS4AHkSlR9OITcQl2ce
16GvCbgor7UZlACX4iHlbMTS01Kluwj64VpqyRQyYUnO5odqMNJZfb4Xirrfk1C/9wq6ep7hSmvk
8EgVWeIgaSbUyaSs+Lq94/wywpTg6cp21W4UpSpNDpHho3tQxyPTECpIvLg60ZPpAnp1YH+lwVgb
D78fmIW++3dL9SnOdCEjzJcqFeoBQENJHkRVhEW7Qlbhe/a68O664PBrPcGFGoJfE0kjivskoJNi
/fTCXfKXQVmIVqhw3rUlWUpzLE3L7RUgqdoncT7mPaOsdr3WLuSWxC0hSEpMQbAoDvfXfqWW5rrC
Q/HF2mkL855dsN1bgFO+xjbsOt8STQcmoiPod64juQOvhkU2+wKdSwEn3ClRjJbzHQZMREYS4BRk
b4sL5B1yKqYdahAlJYBSXYQoyyDUVcak5ZRvxOCaYcspKoGHdEe83MgUeYiiJ5WJr5+cBjXA712V
/b2pJb9UeiuLs15sWMmU5P78aNA7BP4Spj4QmiUmU3lVTD/38ftqv3HQ2uLHoGW2rN+R4xkEaiwM
Y2lb786ED2hQ2GkeBddmdLWJtr8vjC4fsZ3RlyAACGaY/RUsQW3NZl/yTx0/YhpNOd+sUHerp/IX
l2I1SqRi/yre62xakWAVMVhIrZNo7XVhJ60uBwqevcpWzPCi699ZJyQdKNJyHNhdZznSmWUXazhq
QMbij2K8Seau87HghGki+4KCguRxksDkSZJFUk+hv571K041xMSAnrEtOU1ohsWJP/p1kuOa2yTu
kCoY5Xn3JyBG0LLwbabdXELbLtyKQ7CJ1xkaEBKAHxcmHfzhAELB12gz5aLSIvrAKzOe14vcPTi4
Ol/pzmgjwNpU0aeXTKgcSPiUcveV8AOjFhF5OhuEtT3YqwilVrGcfUlVHQ38smfdyd24aNCWyiEb
LF9GsKzB3e0Am7LQoOKImtQafp3kAtQfjQAKjK0551H15Ia+CSVfC9putYqZKkuFxPZkTKX2Y0FQ
7VYoI5/FDWXAyRqQIGG8ByczsYU3OE4EptK17JMWOnQW89qqHjUKEZPJoO3pXeKANX+QRboxW167
b/3/WeBZdDbwFb6kOLXylAI/F9U/g1mItoE/xjBEjvo04aIOraxITEqoaFjpih2EzyerLGUBODnq
T+XT9wUL1PT0a+kR854OyP42n9UyAFp5fNEc4HOZnAmEO/oGCwIiSzM71f6qtq8l/prIOu1fugYo
gX+FqogdnLOJGn1VPgGGLz1tjr6cJrm5y0rtfCc/mqxdNywePyNc46xbgIcISlPuWEj1loHGprzV
qgiNT8Y6iDar9jmHzNuHZiKD3z4DOTrkrFEdcP+Aj3BhtqZLf+LnvT9IRQZSOOVZCxntuPgY6CY3
oFJh6i0XpzoolO1xQv0pXJpobM3hW7zm9VpviPt2mCzjWQWf4nfrO6XJ5ku8RfWMVcAnpykGl2Yd
bfRNF6OgBKN9vjZWqduu+zonTCyvQXoQVXouTjITUdrR7aFRtAAEEi1WPK8QDqY17MyTAU0zuCp5
rWyk8whdvuyYpvoyXapm4SStOWmO6a78PDdOiBDDdyRc1p/axZV3Db0D5X97KN7bdTUzHLbNn1Qc
yOAFiGgVLZTAZe/E4U73HLCLQ6spXom1FTYdByOYjfpoI2dItSYE4uJtOAKqFM/x+ZsSgcg8LWd3
5gvAV9JY6KETKegdktnipXS31TeywXT9q/nI9tyK6idrgpFzSEch0wwiovgQnOiPxozeTHlDy8Qc
HJ3AK18An3T7mbq6wWtdus+2kQJs4VCCYO/8mBc0rOqp2ppt6UIBEtCLkx+Yk5mgdF0M27CfMIFf
sN3FVrEJ669k+YiEYNb8Zk9bvLPskqUmj41sczV18rCmdAx132+FBwhwHFc3Ch8PYvivemNsL4qb
Ano4JrqjGeCocp5qgA+dNoyrqwJw2foK8gmFteJVHcoIyDgpb/OnV8/AUUQU6wz2TjxRftCHgK2p
hYDOJIwmAe8gvx/a9IIFeqKTkkj+zwx0IxsMZRj7Rbn9D6N5Ws2oRsvNL0sEFnTAThKizzb35WHT
VJBTFrGeoJC+q+6HVPUaaKw4YSFqeQTESFOClNXkS39KGgbC+m7hJ4Wf322m15ymg191MBYTB1E3
u+qf+necOetVYroro7EA4wYu4cBGvEH/nuAjutPcyY/sNIHvXjuOOcBMmuHBlQI1spp0TAvuC56b
UB1P7/ZBWYRqFK4TCug4VOUkeZ35H8zUfyGHCz0i6Srkebb8ZVGfEBMMAXXEW/daaTm0zPNALTOG
oiO21Mq+KbNqwCy5QBQSiUAPWmmyazzC2l2JhZ5sWSwml+7TAjyMw6uzgu1ZR7AN4Wmzs132o9hO
B5Ju4nFSdOW+yW6piROo5QANMyQ3BzKSsZOuHf5gLoverHKt7JPP2/sfKywKLJfjALQ13rlwu1Pz
kFvFCB3DWtLCrygAEzad1hZLgsD68L8iL4twJYRili+wfHaww1LIXUo+2fouT75mQmeIiBmVe+V0
/bs8Hc1nMfIvA9T8J14Jy+c4OOuVIePIpOxk9Te2P1Q67p5mJ+lpn3I4b6QcYLqQzJKw3hV0SXTp
dn7KfW8jWLuBW24UzX1Z9joEpDR8sqE27LMvLu3AObJKIhCSltxasOwdoO5uykPYDwvp1cmXvb2F
z4t+e4sA2ieE0LCaGY3d9uHmw1MKrRJ0P0M5pD+4BIraJ2sSlQ15SqDV4270ZtFhnDF0oy4VYe2h
ZdwgskWyucTDFu917sq0o4zXunTkU2lXo5vPE07ntymF7mZSgHWYzEzv9xtU9is6ei9hAfrmhrLA
+dn6lKiXKENjeXirqSAOhMdL+UCYuQvEIaaA+kUi5mYGL/uitN0yrJ71ISozaHPl7TxJH9ABrU05
AgwgGxZhPo60D82t3tPwrR4rndbtiCuhKiWbxF++07ZMaGcb4b6Pf8ark7LFZsG9GjOS5hufrwBa
MjpBEu+seetO8idAImIxVa6PDCr5bR8PUC+A/teaxifN98ATAWELXHmb516fjv9a6kc21q5KSgrJ
/PyZisVpjZd517q+ZKS7s352aLREP40+96lH8wMC4ak0Z33zFboCxmk3bpz7gHBNKdOU285ARhRa
8M2UZ1wkq4/Fb66gQcruok2SSFen7i5oxFwRdqQOBw2yuKeRyYkdr+6QeknB4QLPmgyj0pxS50us
90Rte/Nof7LaKoSBZBk36zRwqQqpyPNqpRgpKW3pvBY8Ry9mn/oeJCNLKLtuEW34KHbrChdRvFdO
0Roa6vF6WKBqiQDiLlP68cjsmydOLwaiZhgBCp8EePFNmCIi4uDhcUthh7o8nj5FFPE9ozbCR3om
rrFmsZx54k4BGmFGRz8JVgrJQ0GyU+azVfvSFUWFMzssXNLXfaiPrU8QuX/SssWimfdg4mlvSoVU
/Anax+yQeBsF49eKLDM+IvKvzQIxTJu56wLk2WXhl7nvQjg/Y/j+rCqPlNXpLe1wMaQGE+uKRxGy
2ixYKO9Aq8T6jx2Ok6J9Q1R1ewWj68PR1Da6zaqIB6pj2Jzxv41GdZ6tw4s7hZI8ksFZeD3tU7Sh
HeAUBCq2YqgL3yEhF7ze5SX7d0VvN8Hg6yt6XKgOhOPJixSSnNpNGe1kaTm90N/CbTS8f+bdP3S7
bX410nzphlzlvjm2p56vuTaIhBPFh5E4NKeZ341t+JZPYSaqkYgf6uSb3B2c5pdr4VYNWgoc50ii
q+R0j7bzB9vfrbANDievtofIPFWP+WsVVBTSsbtK1LEbWr1S+J/E8G5KYOgL3taYPHNwWEj5If/7
RcQwqEsMcvpvrPBc9lfUdUYnKuL80Qgkffn4u/7jjfdmBKiUvNp7pDw2iaQeyflmGNiE6d201Dzx
GxCvkzLPf370eL8nLPzG+VUMosMnIKvviIF5Oyhq5pV9ajJCvr0/1+DgwSA/De95PjZPi0H8V/7M
STM+1Wicw/CIWV3q9nG9sBwCeJyDs0IQmf8M3MIA67utOcM0RMa011hUGZfIZ14Jwp/IWsmpnKcM
QGzgIfUPuhj3styYsj+SHSI17Fh790R8gQ2wnsm2DBlnEMPKrtySYHoyG0fkPW9QDdaGXy0EZ/hK
Wd2I17tPJt9doBwnYuC30k3gst9vLkw3TXSFXXVZgE5fj46YxEBnhgsjVSHwr2FBz3psjH5sXcYU
IB8r7MClHmVNCgONz7VSR+wcdWmP4c1T6FuZ1hCwzcRR8xDCXo9puWi8OpmnIwKfywudlmFXjBFr
QaxYXt5uXzdqFMHvQsloJrNey3FwCY2m53WD1nEFiCTfXXJKphKgLBnr5vV0hCPuz7NjdW+i7/QB
07q8rA6nZRQ6Dy2b69jyWIOPveK+j7aWsVrZ24eDu8oU2cCUHuXqo36R30JgAf6Fpla/31F7EiJd
3BvCJyPLFpHPe3t0Nl63TyHA9na1Nt2Co8E3J15KkdmJ7VJ3J9gNq64jO4Zeaq+jLm41ktSzCUQJ
Kd/bv3NAMlL/Oysh0CtbG60hFT5cuY3trxENshpJF/N0E1ehcQF/AZGzbpO9Z/S8djYFyjjMnXzk
fmi+lJkzzDfPwXWtx5Qipqfp9+sSmnbFjaTeW0H1ycwGLDGQZ/kPNWq8EFwgL0VPNPrytso1JlwD
6cYFAxjaOiI0OLagJVzCi861+R/JJEW7iKVzNgYk4fJxmlgiqzKMQbiZ6KhL/S4+yhKxnt8AIBbw
CCguem1XfxU77JSaUzkPEct1gzcoxAwy2GZrVMqyc8rW8h6eCjRZt6JZxTUyTVFlUi6ZzFAh9eVJ
8USRuOpCSmQSvWZkccQOh4WID9tC/97cKFjEbV1r1BbBPLiYX0T8avScnxVkV5cw1gAGjl5pMA9x
cw1hSZLFRRv1c/iQg+DVAePs+iRHU9HM6vDDJtYUOrtfaB/EvNgz+10n2dUOgsbBSiP/6GG9EH01
wO0krOTVphnK1SqtrZtB5wi3vqtOgGH5y+PzgSIp1Ba7+6fbZYahcClde1IECtdMQMbIU6CMSOus
KDLedex/0WYRT8Wbfjg0FmT6dbURbM9yQzeTzBwvo62RjuT0s7KxqdMH8SUPkcOFRBMVfQdBsdnn
Z4kYye1Kw7BpwQYJhD1pX5YbWjdEDac3pYbQtXNT7xKxu9UK9hB64BzTYrmWO0tZX2yoBfKN7UzX
8ot74sY49yMiRzy/Aa6O1h7NeWPiGCXRcuya3+0ggOoJnbh02NNZeySV6+Io6ELKbQFd43NhEZcw
w3nsfjAjisHc3ZdtHZGsdSw23GwlnUQ9dFc8ASd1ihKroEZP4/Lq+sa55qHGJsOS30rLWe4ZgsNa
h+hcaNwHhi4v61lxGBQ80D3zasfm81mcDK6XTKMhg4onv1XVZ3CsV6asdNP2ExVWOWAVI8Z1K19r
jbkiBDhQzprU3H2Hhs66JDhPyfYg+4ki43rqe82Pc59mWJGx1OYs+AVAtBHVHL9f3+jMUxB3DeLV
rB9ZYnlMtODK3YpbvPrLrJ1bqd8LIlvcCEb/NfL4ym4VFlmQmGHwbmefTQ1lsnhi2pGPeFYew5pe
sLT196XV5z3X/H4RcgPR4o73CrN5EShOrtCKVcA9YH2Id62QFyDvSQGnJClx8jFDuOU0RfFQAo2j
M7noov81w/Bj6Fvs8FFpW9Z5xz2NLhr1Hcjy20N2F66dN9ixy2YJI+xPn6iaSRBlpL23wsfyT7dn
7kjmb5jqbR3ckYINyrHeZYNzMOhz107tG/oWaUSdWA0XS88ZxcJ/pB6kGBHURdidoQXUyPxIOvHf
AMG8ch6lgPu9nGuEVwbzjLSwp93h9zD0CxPX8CdTtGv4PbtZrj1mzhKuR8qex4VtAnQl0Rlryyts
Kz17/+N76EulPijVc2ThheaZiuoX6V/WBSfBZTmIma7CB1rr7IEd/Ig793Lea1Q4L1bqE5xqfkN4
FSDJOtz3bh4JTnBiGQ0YqB5zDC1RDTTt4bCO/lf+C8KdSabIgPsYLkAeC6+fCvOTmHDOPvRamJ1J
mC+VugaKc+vlgP7hjJ2lH/yqwvmnEDmPhqKQh13rIc/7TgW9Xu0WPpOWVh4J55tXUkcx3TuV4sgY
T4Pw0ok2lnKR2C/MlzAVQKYKQHT4WZE128y0lNsjkhufhTE4Pqab+Q2mxvMzLc3f0hzcWE+Or8vz
VztRWvEnUX+HO6ULSHWVrgEnbHP+Zry7LTwI5eLQeTjKB7Dz01YuOzQE3R+h/qi18qc8XBOoYpmT
qjGn9fTRiiCnMf56o2FHXzP5LDxQgX+Y3QXVUFWsTv44vnqv17S54JP3idONfLgAHn6tU9lTczpd
pHqHcXvQSDo1hADaaN7wmuMzGlJl6ri/t74Nbj1pt+3IMrirlYxIKGdcuGLXNv2EJ1UX07QkQoAp
/pO8vNV+jG5+Ojf36tYYl7hkNiU51dtLTFVWGWD7BlgZ7xtRBDVMxih26ZYh41zVnxw8RZjtJ5I4
0psOeGEHpS5wxAz+i9kFXBOVS/SuvDk9hyWmV8x/hSba9RK7N1KV5hUbsokpUCWDWmFMdyzh6HSh
FEQ/9/D1hSywDPXQf6txywu3J6CcPM3E/Mdn7TCroM4epNXmE9TroJd+j786MNvd8qadyHZN4Se2
uD4FC16fWhWB41B2+qtTmZZtYIRnsTTxccKsj76LMvgR+vhV+XrNrt0sIQyd8G2Y5kfYlZNc6Ax3
EfKa6WvHJ0ICtbydtXDNKDdBrBknyZhydQQbF0w0Xxk0bn1dG2YbKAgzSXcCTYPvpLwjnJLsnoow
yVgmcGfM9zE2Gr8laQ70XKkdn+uYYV6JQFue7X8K/rxWAnUJI76Yxm2W9BHt6TIfzcLnU+FGqStV
68n7LwCfLn+X4ecKEmkbEnJPDLnAojy3Pt9APvo8JATxzE8eDPp1di31jWqo3dOx0XGpeYyRrRVp
Zmuh4PN3Aq6VzVX07iiRmrHuLL93xc749QzW3U/QGlaZrqCqgqv6x9eEhBIzTSfgSBEWGbhZn7Td
noMrsojU2NE7cie7M6xwzMGkmCeOIdKi6SYveby7yQ87f44cHvID/AcX/h+jU67K2B/uLNtpFXPj
iwGsFSUcVMAFdMGVGc10D149nFPj2SJT2JxxPWzlGdeP++K/1KE1lVPWxWiFN3vYh8BZ761xNvhi
PUmRIXdNGWzHuzGMuKz/vsi7WQvagGXeUCl5CzMg6JoPZO8eLvc+FwMKho13tNTK64Co2DY/fBHQ
vg1vcGs4v1YyVSpJfZPnIJPTXWINAwaN/07x6j7dGRBOl0+zj+VctzTepAUd2stwnExUOqwozycc
+42jFmrBa0A8krKg3FiquvdytnryklQqrOi8qgwphopaJZ+MFwTdElFA4LLd8jG2PVYkr57lQjp5
/P7x6sn2jG3flccAnunvGbWlhtiHh9JN2OjAaCEmDe7m4T7NBRZ3kkZr81DWSpCBI1OATBAfinwC
tDbccIvgZtKjg8ehIsDZGeYQmIaSdiYxJ5tmR4XotLXS9yf6q/jAOcM+Bw6KH/Tu9pYqVVUnviTb
8YPzEOh3YDos2bQHXZvhupAaldEgKa9Prhh9w/CRNgxiY3RjaeidMAxzXcvohIZfuqrN8qEYYelQ
8/Qru6x8f4N+JcC32WYzJypCgffLDtDFx3UVAK7D7uRBARXCwh3jOSTu4EUzXvcTGOdvQU9POd6F
mWWNOeZGdlhZiYmrsTwD77XSsiaBUGKzdr/9pYsfRt5CBNzDvstqFzePNND+ei1RWhoCh9qYWaEf
Ham63aJSaetXh1lb+rfrf/lcsYwbP9ZS5AR1K288IWcQg/EOujnvTynn9EjXDXFNeMVZGffVDVe5
1p6WUlS44gl6sbDiZRM1u3r7Gj4uWCnYWuM/L/+Oqhl037KibXk+LOiMdyqVi+BS+SqfBdrHS6zI
Lxevxsr+afIideGNOFdfzi2/l6ouHKiOPRbodu78o2vqwSfbZZCsRsb/17FILMkpHRLFY3CYcz81
7POEuyN9OQ/Qg2jY8+dJr7ZPYvKEl9hrFoTiQ3ct0Rtauvzvje+vSyB1cBCXjChuZOYzdGkrRPMh
a6NfunH51wr824OqPjyXQuiQiIcKsgB/nn7K8YMBvfWbrA108NSavjn6ucEMKH785abBD2A6+i/E
R89v/t1VVyn5yc/ingeKHxdS2DbpaUmkXhpbHwJEyVEvo78lIXj5Nd95aHzQ16sQ/oPXey5WgZUe
p5UEx0GbWYVhv6MrtgLdh9BoYsTGQUOANQPppBkbs6JyosDvjCYOxypN8eTVWL3eO6TxYcLCpXYV
Dzb0vcdXK/+IK+Xa/rJfcdNRAyzoGG4H6jtuCXQOWVMOtBgpmyQZhMZr2pyxNEUSanSDDDVHpcgp
j1Vr5kDyTwv0YzSf+3JLBHHiKyDTvjxhJvfb44iIou9FbiZKTjpw9+gvct36Qn9LD8/9IKuB0Cqj
w/sWSPEUB+w0potRRGsZZRNptzAsuXcmxq70a2LO9dNSHISz6kwgk1sCj2gZjStSuyKXZcrEqlmZ
44XWK9vjDnrPwO+OO28b4yt50D71B4hE0doxhk0Pz8aMV0SUNBj3GGEf2bBlMyjc0B2BIcKm2JIm
XhT2fOS5f+pr1cjnMlE1XLD4mYLaykFNK29++bovQWS6jrXD3Bz+sYlWL1wdDb9zNWxYYigR5HgN
RV113zOfAMpfPjG+8AiAq1+Xh/phQ5yvHL8vC2YAPnhoVy9THpKQLZD001tV3IDMBLa7ZW92qU2G
VCVzQ3T2uy9tFMvQGmbgBQ+P+ntSWbWWDZVeIYOkMFMDHEnaeXBqyw7zoJnVX9GyfK0/yVA5jasi
KsuKQ+0D/5oKaGfvRr15B5LT4d0OzqbNqWG8mgY5aSzoANmZ2LDS0UCh9SFv3RdGwG+9D0S8VQxg
/14YmO0O0IQy3+4jeWeOK99FAqAZj06LQGLVPY//EVmkUn7tVwByI/BLNSH+BohtIJA1SMHbTbiu
nJa9cczpHgn6sekeaZIWtn5h44LkgDitx6GGfYpp8ABTpvDRlZGFI6BgZf9iWoZFlSoWC4cBWRlS
OdWQcSn8NMAagazkaL+bW2fAYcX8LAbrbhvV62FGsb6wp6tZIghV086Le7mLBj/5/Rc2xsCVlV1B
5asctmdjLCgpF863QJGPfgwpkNpYsPsaGvwukPiCVpoqAQUlsEG5+PHgQlW070QpOclTo1F3UWQ/
rkn/h6KPJeOM750C82rwsgLPX1IpZf+xGv1zxm5sTM5ZBgEE7XTIBCY5hRGlSLhtTzLeSvdgaUyn
mEF6h5f0jqKkhcdoA20c8uNVu/qfPHY7UMBF8mC9zX/6oD2e+Uu0vNT6lxM3F02MXdPfpGWenkw5
ZjT718Wp9VhSbZz7fxSg3m6tYD/y5OO/qfdkTauI5LaS9Glkajds4xdFSz1axAsgXDA5WjV6yBGj
5aCbsbQDHKy+pd8hJmqtikmClRkscSSbp4mlq+i+3Cx+Z7D16N9FzNtjaejIzIdj09u0YlUZSwqG
4Pr9fluCJG+hIt21+rAtnkOivAI+KF+z0b6Ud9SlSLlz1YRTDhpYQfB4swhqn7KMGdFWcdaX82Fv
JYY37osOQseFZ5SPybzxMqhtCq3fFmPUyCBfx73bEY6wrRnI+dHOObSW0A2SlvEobBimL6ZAdcPz
1vbSG5kh5/4cDH61R+6laB+uHx8JQs2bqwF9NwQiYDj9ZKc0P2piFKlLxSDMUUE1RBQrND/yLMGJ
sQYYQoPp0fjvhtWKo4PfuK30zf2zt2H9zsmdp4snE+lQvNouF8rP9MSCkHK6o1DvEJMh9vbgQf1Q
aHHLze3GVyKaX+OFOQIMlyEpjcR3eTn2JcZ3C8i6J/saA0OxSaxms8GUdvrKoboNc6/fPpschr9/
yPb3G6WU/NbsZJrK5/6vAeEsuT7L4yPO+3rOxAJn/sztgrVOxgxaiPdKiMSkoqeS4eKD5eZifkz5
nzvzrnf6Q4sIYScvGCNUkY6hWZalt0xcIYLuMDmlx17IKueDD3CPvPnT5tnCePB1uNULWKC8lu0U
9CBcvtlxgRiiK5yULGk6sI8LTFzZvG1IuOIuIUvraqDDVIBrkaX/jhI8ShqsJQyW93TJdpq9HjcL
uD0WIswZAPd4a53BkptoXPPcNAAx7uZkx11jvvdd6a2yFoSm7JQIw/alGijfGvxra0aOQtx8dRUZ
boYOe0ZX/jU5M29q5YXDKchiA+8M62zKwcS5JN7m2docJDnnFAkyMXZjx5OWaF2NR5SLNL6OcrnE
6enVpXizKkaC4PPJJuHgLhyxW0BXUqvDcXIZGs9snehONO+9vPqmkG2Ay6tw3Y+maWleV0iBz24n
GRPlXPYNIoGWFc35QhplRewzZ9KQ4w45wJ7L2IfbmQUHd4NweQuFdxqgEyKv8mMNbmMFoE2ZsnaW
rLji2Hz5gcDC5xuU4BhofPvqtlNIy9Thg5mMnZrXtAmD4J/itv+lJUXMD4w/fVMQ7NXSv4UYxrxu
AjXg3XprIOl9piQrnEH0iLPZwty4uTkQ94P11MNurFl/pbgHR5AxEDirlQ5DgMK075+hWPcPij9U
RdjG/yTBRqcCFH5BQRUf2QSkyP2t89FMXcncCNUvD59UD/9DsQDylPHSMWuYhiBZUWheGcjrX6r7
PdusNsqrVQgaYBe6PB8Dsqj9TjWhljyifGEpiUpfd8foR6G2ebJ+Hd80hUNshji2sGVQ1xDEpRjG
ob6LNpTMZXJ55jVDwf7vaI6gR/je8o/8lf8AXK++D6/wunevY1Mw3Ypa9YQvFQCy4hZZWQeDZHxA
480C/mwrTw67xcKyytAs5mvwqF8TNfMqsWAATmi2dP9TP2qVba57ZX+eISCjCEJMUh8IsZQO/1B9
MoKFESODuPC21UyuUefzywY9DesZt1I5IQMAokam5mg15zFgoSSv3rIy/eNn/+CknR5XOcT6u7xQ
CUjoxICkBOQGxQUxbHnQHbGxvzWELVwaw53QZNUTzZ0jaqxnYCjHtEB5tZ6/gYmuzLKJpFEVQOXD
IL3++3X+LdxMfKYiOxqLD2bG2cgSQ2qAEXQ/D4psf9pd+TSE+Kux8ueIb+YtDskVdabqN8j+iNgE
Jy2rJK86nYgndAfPuZ9tOjpZAd+8PyvxVSlL74W6m1uGNxkuUeSJXr0NqDQD1tEprwTa67bDxDes
xgb9RISFDd4CKkU+pvJySc9ZoGyR3UnIdArTqK8fH2p7ZpvqRl866HmDNGen4j81McSvdkxEQQ6s
Nkn1ZlsSl3HM6sdF/vJhqVyz/SaY7Bp+4efis8spXhFt41CGW/rVySTKZkxzjjJAinHgLckg2J6k
48Fypq5V1669S6jjKWoGTI8BL34Xsmh8A9cWrXRYvQwJFrSU2rILERdyBfBapKhj/XLqasKgxHL8
R0D8DfFwUGoE6YB/ddePvn6mUTz0eSZ2JJq6HV5ledd5AjIEaQvSoXhIOcLzSdAXUIu5zy458mVt
SskzuN8ZPmQ6YC+QkIHE7/CwJJXSokN8ypkXqka4IaktvGQoLrvrP+zgd9AlZT58NffF1/SdvgY1
Lj6FIjj/r/v0W3z5DKFjvYChJx/sv5xBxTVEF6UqkWDoZHvvf2pvbA5EW5rfLN2/3yOEzRifzTQh
lTHNn4gG7a2QepAOK8df/68ozGj6PXlhx5V338bBdiZga7M1MUidLu+Nma6pDIO4Qvcd5KD5pac4
68tnpgKF2YA65RG+Z8qHdDW71Iql/LNDSk4Dksqi0RABkGJwxv8B0HHgKd3iYbZzK8FEV6HZnfBP
evDwoNVqXdZOrWAlbqylcaxP2G0ANIDabMpZJZUPP18vTTJs7llYDPhaX+j7DXfK8Hob7soDTYA+
146SFo87N4JVfYL/EWe4vzTbZYcMcGsrvvBqKGlWyM8H1hfJcbl/jynduTuZeFhGzKN9TDYeuFN7
j5i+A24pysB9+wH+exx/TcJbYG1j2lxbX2To+sO1K10BvGfBy53tgZJ/jua8209AcdKnkaGAEbAe
mkogCXlmWXrsKz2z1OYRL0fcybehbYk5hVBwRPmPHs6XktatSbIP+cqklg6e35q/jk4csMuOsQu+
SCSOdCQBtK0cEPbPRqmh3L8ZWX08sQCUPD70TTn7rdA5WAWx9hjtje3IadiATm+FX4HIJgYPlY8a
V5S3TeZd1U/W7VLzEUVWdnkVumrAZNsW+bWdJwZdx/aP5XCn/4sOBb8Fn8qYnkB+qo034HE8ol9q
y8VRSWaCIp+XaiyTMvQMMqBTrgCyGf8RQnKxMeNsutY0bHZWztI05wBrh4zlsFLmMT1iQshEfgZe
tj4PB5mOAyL84NBqdmQ5tWog+EluCJBioslCtKA2d5RtSUNZw0T2trbpPCM9i3RwDvSj2lF1PlpE
V8P1/1/roz8pWm+3GzwR48oJdxx2oW5/aBLTanJyzaK8yKXUSZTIx86KZHHapyLurzkzWEtRiKxZ
vDEaKSdr+MN+SX8oSBgZWAncf0AIis4a8qNMtCmeQvvXxxlfTQ1IAKGxsZuHjLGx8o3oTrXPkkqk
ace69nmvO/qnbQ3/Q4mKZ+YXf1eLUbfdyHXQXS/pl0nDvQvUW9+tJtuxHjmULVNvfvP+lMvwL+LI
t0uB2Ku6V80p4bNpO6ViPCxdhMFe7ZWEVpYINfolEUn/cUgAlbAuskk2ZHZ38yZwoU14bJe3JjuV
3ymxb0OQlWg/dAxV/5MIW1O4i2M6bqL79qis7TluVFkjN9+IaB4QKNpIRrzJYV48GZozRjYYPrM4
noKcdc46tHdjJPegtXQeRVbxcQzpfWl76LMxo7QiAL1kRSOzX46RyN6tbI1qTD3tNSnHfumnTLkc
WhBAQeyNWBNFTcu6CJS4/pJvYQCiMVUS9hfXYQ081StWoVZ3lYeZ99SvwHGjYkZVXM6MsTFRLtsk
4rIsD/RQQ+1/ZC8/HHECom5fKSRw7iiHeZu21dsNy0YMQzabB3YR8vVqpu7ObJaXXUXqwwxxK4gm
l1i1ypDOng7QhV146whfProt5YoCa4zWYeGvLnFJNUB8tIOmL/k8Yvk6No5znBTlG2e1pwB11/Dy
/CVdtx351c9Fxwtb8mty/AvspmHKU5rHXf2bSGdsXMyYxy9iW+CjfPdklPtmH/5GB6RZMgKl1aVn
0cqVNoXLKMUnuJX79aVr1lTZ6/mEfBgFGuC/FZA3+73GeU4DCG8wqKbR0vl8i5p7hs+5JfDRT1rI
b5uc2+L0fHFJGCUGbU32ZyEmtUYMky6UKyeg1rIeYuFAoQl12qhSKJH6ojH5d36scy6CJR5Nswfz
YfEEP0yD9hcZG++YiP7/RQn7DkYjPB3RV0l9VlFFQ65L8GPpuqZ/XHvUmW7+PlTDIFSgXxJ1BLuH
1WYJylOXLi1VfS5vRPdijcdH9ggvlxAXMUnLI2GdYPBvf+Ja+oEo8T07f3yRsareN63EJN5MaWgc
lIValvGdxHPwijg6/PeVlspJWqKRNM//jJuskPKvU9pzy0TInh9zJUPzgmu7jMP9pLadasD11nsS
cBwkZQ6GnBd0mI9mKAjch437IBAmfDeUqKeh0wA9q/7s1skiEarl6199F39/Eeg/vMY2mjfAHSzI
1XD23IkEnQ4dQJZuIMC85l6EIUiJoPzYFtcSJckRWsEmrMiAAlrE2Ofgr10SDq+zqNbrGiY476Yx
iRX72jjaDY5DHtRaFZ9puPPKTgK0Tir1JAvyb6rvxigVbcQT6VddoFf+cE0siZGQYYfE+fyciBxI
DZ5UQLKCCjyerXMr9E3wkk81uJdJR0AO0X9h3zKiomCdWtOb+ceW4+3izKJXJrJTw1rhJNEK69CR
Jg+9toZ++cWaQ2Mj38oMjyQYCXn18u8wKRXxpTxids4y2CP0rjHrvatG2spF7exJlnM01ktzEaQK
doHGWt4t/2w+gWNt7SOS9SIttLDD49JEc+lR3DxpYdjx96ZtItskO8vW1c/tkgy6x5fzD8530pf6
rEnFDJV1PybuFN7a7Ci/XNzeEtl+k67brf2ZV0lp3Qp+OwsIHAp8lJ56QRXrD8wiOlIQbdRyM+Gb
d7OPTejPgfa2Ow5MQhnOvq/luqXcqLyAY0v1OpmWW4cYdVaRY4GIxOUzMMKsalERWCoxWfIhc11t
VyHUAbdWo/nsaBwoDo4g2p9zyS8TxPz6cJK78+26KieKgaq5tX7GnP+sPkV+qiJJt3XV24iVOqcu
qFWibgqhMadc9Mpk/BIlVgnlqWq8tNE+UBDuHEaTMpJQVSSTEdKyq1Z8r+r8JKYj/Jzy0wlApsYO
TnxQNXPaakQf4fGahLvypc2K4U0IjFML2JF4X2XfKhMHG8sSWTXugJmFvtsSVXZA8ThgtvQRT0yj
xSOiFJMow4ybqcBzJai1a9WCezpyJCjw1FgLgjp3HU84iEwYcRldLCWr8Vt7LTifGH+ZxQZQcJap
pMMSvYpGXtSmVOMG2xqL4zBbgVrUJGL/QZani3wwwooLjbzg+oA1hpu4NgVMCrB+EmLdNfpN9klB
XlcQM/nadVQAgHVEWoudsNI6S8yfO3u+8rOnqOZnCd1KdMPF6dQI2Kg5QThclu7Avp3MoCODOp8r
tl68vS1X9v4FSnAAOKzuSqjMUlqEwi34cRDTEf3TdXPGNbA5hemWYxDbXQcz+iHhQEcuCf+AW1EV
gz34qNvrFQ7CyrZ9eLVJ2i9JEDmRiuPpmyjaW8EdyS1Xy6Ki2iwLomgV6bwKuaaUL+ZNLgdcMzGV
1p1UMmKtRA4pbGUFgWHWpWBHno8w5cQEoK0wsphtHjLPk/fP9ifIo7TS0xHEF7YtbMi6zi6G6EOk
oOhzN34x34M99yYKj5bJP9Qez7EgoenrXHgZ+zT7dYrQCq8J9JzO75DuyAjSrO34Y3n0L8/ji2li
yuDhuzNgu0l7/TUQ9qWA/m134WXbPu7XRL8aeGpUV68vSdYnvwYia0tmdrQbiQov0qBE4HAAITl3
tnCFfDrbJ5GZuOuBF6uyiNMXPWP7ylr7hmxNTuudE0E1GKgWeuursvACATsX3YaYqrnvOW9TsJ/1
KT/1yFQJ7dgj9VgfQMldFfBiUNrOljrcn5SCbZB7nW25KAZ5jbRUN5GvFQdUOXF5xt+ww7HQbjJs
jzC9E7dCHTpoRIZb4A6YHodFeLqCt02cYgGBrK8dmVun2UhR8kqBaO7X97Zio4KhhFjmTM7YIc3q
0Mrm8gUNzHbvOZXhNoX1jv32Pi5VCk/KdqfoWu09xFn/lzJI3owwT4VJ3F6KF6xEB3T+9CMNPN/A
p3WnWm/0dY+beoNl/4TDvAJuv9aJljnRJXdVnEQS9JgyWgvgDOPOhCZd1DKpM44Db4stG5B+OUOM
1JmC86Tr3IM6tBZnWnmGtaoYhph6D/JolvdFndRSHA7NB4Lr4WT/eia9qhWosYOPmvj05M91GNia
sUKpKvhMcIghr60zt6kx4U4vihyOpefmPPnQCOSVqISCd8+lima/6wd7MtQWXJaDsJD67O7S0iEx
vGJHIsAqBMgpETFgPfOYJVLISbxf/Ga906MgTkSVezeS2VtUXmd8hHVTY0h8UqJSrJtB2hQqYNN6
wrvtSUi/FgqhgPPTiVX8NI7YoXYhQYRwzyl4VDry7yYCj+whiciEL6VigB/tF+l8GXZ4Ascfnp/1
RO8fUHwILJ1USwyZ5wcfCJxToiyt8ChkIR2tf8KPW+NqK0fhMvVsV01W+1RGvnVO48VqlxWQmdsA
4JLMvBYULKz+RpD9nnOqPfYbyrC+MyBiKgUCjUFa5dyRQ5ilBxEtdHKJYgD+FX+5I9pYf2ZkJDTb
l3hRspF0/6xIA++dCX7oRqcvIbUbabEJN3vSskA/3WNxSG5gfzeeRNLqEGtSpL6ue1UhloM8qf35
uMHnU1JAXw9MERCqbLk+JcAR5E4FfW1g/0SXdrIzuzm5OwbuzFBwQALTleII7ff4ABCFmgugAT/B
rxcAo7gm6ek+okbqMJyZj92LpL3wDOg36eBcj/TBtO7nZNQ9/iAiay8DkxfhjlyZuMXvcBmp5EXu
DscgFv2ctJ4G7FlEk4qvSiaFlXCnLtYoErUYQ6HeGmZUd1G7T7PgC/BsbTEtrj+n33489gseuvfQ
UrSMDN1skp84bLSt43XjHS2b6sbPO1VTISKHGqyOEyugGzHdHI7UNAtq6ps0lFW7SaqYZw/VghPP
Tc4vCCeCJl7A59UOU05CQ5t6qwR6vY2gKb5jEBjv5tPdxFnnZyVYSjEeJ2Tid9Z49aXyzLELmuXf
CiFMlCUFDMr5t5kt/6prLk4yWRM7iTR+nWzdG2ELxbKPznka4nPvaHasyQJQWlchnQhVH87gHePk
7OBjk09I/jf0A0xI7AYW39R/Tnv/etvPDstW/3c+mDgWhFnxDXCjbfj/oqtGoCCL9tnyXpxn+kIQ
PAYDIKiT+IwG1j0KJ1PvcNwxzeVuh5H/8P8ltlnqdH/TcqWCCb3IqfMJ3GEUFRzeaDEM8YCLip66
rzTH36QcvTeP7wpGsV+lAQuz/pjMTinCDmfxFshFmkQ9YHKuwpqdL3MbZdbOcGodR+eVwezkDMVC
YLje38jOMXFdTXI7mVNz1uGV11dJe3M8X9Qwo2vIjhTUu6KZEIUI3qS1wn6NjeiQN3zlStdpp9ZR
uUEEHQwaynryRzgbG2YSLy8zot6ZgBfvsCHXhRuSTRMm+GBiTU1zwoGIEzIv5J24Aam2n/KIPZHX
LJhew5lKH9Rd6lyCWXhz6Z51xVkNVCnGL1BCzn0iDR7Qy6jJKwgqV94nuHhEixDBVLg//h863F8R
Nmgom33EXjPGrbzThEJdqSeYiCt9CgRAOuf9i4w4WT0UfQre5nXlpmyV1tfi8u2SuJ39+6Fh9s1N
f8Fh4+k4WObIwUtuCI+qOsnqt4k3J8ew3UiunwtGWOy9TUATn14ggIagjk9cOd7n71ObUTpgcN6b
queRV26CQYA+un2s+DWkQtshj2BdXEubMxwMcdZPsRhzHlMDMkJCna2EDIZlxeED9KhDCpdkcHuI
9l+siCMn3AbYSLAy/qiepJwlZN0hnU0GgGDeIRGkkuq/VUDklKhoiyUIhO/FWQLYHvZ5aHgF46na
gxD0M63TdagOy1fSdi9EY9jkzAn4XjDy0QMN8YKLE+kc3WECtON70BJrBzFgGpQOVzKBcgnml4o/
1FeGRy8O56LgUDeRoFE68kbhBLDIvOxDOhhUZd65qXDAmjPoYfoJhYYufeRbt94MHJzqcFFk7yEZ
1PDL4nX5z2hINanIKDTwSYkqC7AIKIaMObPI6Ba4quzpKCjKATYv88ktAb0MMosVb1/uxGMfrSmK
8mHycDsgBQ+PG5jAXY3cImrUM21cIE8STHiowEtYg54nf6xXyuYk0JvGk5DXbG6vp+7Pi0QI6tmS
93Od16nr6R5iws9/e7TqsxJb0HZx3ZphbCmXaSkZ6sONlvoVvzsJD+49M4yATyyrjk+FZb2OPMGl
sq51hCM5j5siQDg4Jd/H322C/Onj4minCbwq3mozyKPFXmztsfh6bNEEZuId1s8AoemXS+yZbBIn
TS+2LOtIeZFPk9P+LvFHEY2k/lfZHo6WPCpvFeVoD/bG3uOXt3zRYTMRFFqTP7zqCXXwJ2/Shbkq
fLi28I5PpSXpchawvhP7I6gsopXItr4pbTlFkqIrYec+en3mqqakAAHV91PCZKJdcxhNjV/p7dLP
LGZSc481FgsjNf3SUA/qFHKnV639cH55l6RacNVJxmTKO3dq7wz83JuhHQDIWy2wtTddP18oZLsQ
McC7UDi/J88zAmJ1DXclsK4zEmRxwKwEWZ3Pk7bTIpn8ZhYm2X/8gGVgiOwBiON+ihyA9bxwT8qV
fT+w5+bsmv05PdBu2vOtlwZEY+ULWTOsF0eIkIEzLDVQcaCe2MjyuuuEaNP9ph3Nz43OdiWSWflg
zIUB+FtPdnCfbqHasSirG3N/TMoyHu6F8ppbSwVjDQYUzsjfk2mYfBbjDBMmJ5M0vjyaNiCl9/7W
JxF+3G1dA5i5YONy+EJABpvfX1RzPp2JH+h/QUh53srxdN8OT2p4p1yePb9tJrtiZOLzCq3V2qCm
Haofw/WJokS1rXBw0vXu3LsMoUgaT6SbrYurBRPZSTJop2CPoENTbOYj2yQmw0oxvZTTYMBuWZb+
NNu2FtBJtMT1nAwNuYqEsLxUc2qD6+7gP7N1AFhAcJb9BjikDiyqeR0+fK5P6bLMK0EF/qoFngm0
tuxMRwLXZWoEGIbuQJs3RgX2XHdyB+lk70Qz1o1BXsBVvTVdLa2eiiPqvrAY1Je1vnS51VqQbfDH
djDXXWiLGiiOebufGVA06BwW5LM1H2MdC33ZqYczkgISaAJ0yIpId+hAvP8Rot3Plk23hy+efOLz
wKbgkuGYS3wSxGcFsrEo6mAbEUyzz7IdcstNTcsk5jzc/YQCqO3GuKSjB6+84LuLDymfdBUxh88P
ufX7MWQa1TOwr+tn60sbBUE4mMJ0HszfEQKABfY3WrkXZhFo4zx4VPkCch+TUPG+dP8gTdiO6lhQ
/kNzRbxcY+Ml9/WDXvHsscyfzV7zCim0py8VAjg7WZLLGWWh6EcbFuXhOB2Tpvf6XjwdAu6wkwq/
oxvuxJjNdw7siMRTcXlBZHYjgrP9ynbvg906eebQLJDsidvSY6g2Glyk/tV4BeBhqGyCS3NRD+Ww
58Wylrh01YZP52ZgCDZvQUtBuSb/9IExmfSmxvIsBuD7y1lKn/wnO+/Zcr+QKo4fOrgtC1hBSR1i
w6cWdqDoqHidC95wsaDCMegFcrj5dFXiyG3d8TU2pBFBXtrX2x3Fo2q0GvOLljGz1skutlVJKymf
AVHOx3RRs2uuF3prylHVDVj/Us1Uy9Pcsvz01lhUuQ/N3ohuhM/vnkV4Y4M9sQ7daOUCUv3e/fBE
+PeX/8+jY878ROyPUSvfeDXaj+HtteXs9zGfFEa70b/np9Fq3a3QDnx9Ab/hu4HbBFKMnDIfx0Zf
PAZhpegMPc8FgFgt9xKym2s+p3dRxX7T6F26HV4LT2MJVaurR+xgdQdB4MhkxnihRSw6JNlmP5mO
mlsEQjbiVJmwbPK6BNiCh9Ej4uq7dcywn6FFscNaweiypyOQKMfBUxavYWOt9Suc9iA4Bq9T6UK5
dCP9GFbL7tmcetzYn22ECQUe0Khjku8is8S7uMc+kpwBFu12qm8+64oR13ofqrF88IjPn/wi827s
3SiGqUI3oIO8P9Xp2OpLcH4nb2ZAPRZoEgueHj2yBPFhRyJh+PqDvo7kV4rCB6V4iUooSk3GyNXI
+PCOoJXUcE4pDrNm0fRQL5lI8/uOvUFGyuliGWIqlRMEDYHyu55IRK8mat96z67Pb4Sms0faLFU7
1rAUcJs003C62P5lr79suzw1H06LzFqyS72+oeXxK/ejiFrpr6V4aWjv/2/hjms7fmxlhCd2IUpG
g/wF1P1zgNz57fYjdk/yjHw7ajCQEo+yu6fqEqbFZ6ixQ7YBPuxSdHt4d6NELLJweWdjj76YgQ46
0dqp/VvrpbXCdUiYnokK4UC+JIVZ+bGA9b0XvAbLdbyABDAcy3Xif6Q9jEwnWBru0WvXO+jZFg3+
KzJ+KveTzVFfRkIRLE/Gp1EARrJBP5DhEfC0U5IM21EHPgHrmJDam2593ZuT6AWPjIqyMCRO8lDU
8UldYrU3IY1WHZLhUvyJNxF8N1gWZtQzXZzkSXVpi4vuD2QjmS+yl91fDC+JNFsap/lTrKahahQ2
BPaWad++xElzd3Q7bzSWtTYKk+heo0Dypxq0HjAH6fA72guvufiTfMFenWAnS8sOZUXdU4YQkbFC
FIM9fPGDIkg4z9oPefb1gdO+oM3wz2Z8rulXve3/3h9UMBN62z/USVMV48HN/HG9QFTFk7HVLE47
zF16GxCfg0ARpEYfnZtjo20NUBV868TsIZkAZ1Q3h7CmmlG98J9tV48J8NAOTq4ilNwcKz6oZBUO
Os2uBnFTKjc8wf3M6vopaIs5T/aUa2upfqtgi6aE6CnCzdMTJNueILGgXBFXd1Mj5BrYG90z2at8
qQlBwZwi+j3b4A7W3h/nysF6xav0gLdyLLtABg53Y4lbUNFqs30npFbZu66HOTR8VbBhgK1TQDOJ
pG4s1MyxyMcW0z+vcuHGe8fOVKKKItxt0Xj7+rJkfEQZF3yZFnqfiRF0ZoSF0v18WOPzXE85jP0W
FK8RDnjuaohpPsvMfpnB6r1PBJZ1Oi3uJFnbGrjUsBzXaBpSI39MnGcWXwqa/Cyt1lL608EWwmiC
FHiwp7u8xbwZh5jqEiw3NYwfZoXRdwY9jal7OpJr6K86x9AKATaXAKh0TnducRNcAhEZJJFb6oxL
qZkdm4+qxTBQFugjzPV4kRwUYI0S4fVD5z+q9W3ETVq/V1sGZdfq65D/b2vcrYFLABTJtBCe8De7
xyJqV9mJ9Au8kPtMGvDdyaCpQfyBQPyCEXj8j2GqE6g7u+5gTtrhE5JBmciY3gMk02TXv9WNNwkH
t3mjusMwgHb3klJ9HZAoOvUOKQouOouf1FyIywO5zrY2nf/9HzIVRFQgP8EiXzfftA+dnxWykFRt
6VrZFfSNQSTHPuQNR9iGO+PTVMibgvL5pDpKNTGzkz+5Brtyl+DsU4u+a7Qx0hTe4BPwbIZmjVbq
TIxucgLDSfUsfv4zYxiB8La5tXO3b2uaB4MrK3txdN1rH0FoYRVgR89aVa1e5YUU8jaiMORgd6pp
5n22M36btGTpXIBWFmuSWYm9Ex1N3FFYsDN4fhTWl70av1O1FHrVBazhcviPzCdixbWgyQZ1Fz8y
dRwksKvT54tYghwHWheZGbK61PAEKwubz55bEK0yZROaTZVD/mmPh5AvpT8HLDNm3qB/BIbLBgMI
XUQvnBDlUEZZAdmNZ/ZBehJ3PFgtO9Y3ma26RVA5OnC/7AtYjhiWNjsBExrcdCsuvHZgJOrZVegk
PD3n1QMohwuu1uMKhtLTLzOAGbzNw3wOOnVh1gCMzpg4ZQv/vNAZ6d40j4E/k+7zyPnXNkCyUWF2
9JUCS8cgFZ7otxBSyKPZBMpaxq/5dewJZ2ghCPNGjoljoHd3qpurj48gysyMcLeabwqWiOqmXYuE
Mf+5k4oEHk+nDpMOLiC0S2m1nUsjXEx78pzUH9udSmio6DOaKw+/HHESui92q3Y9M+zktej4KDlX
YNkaRStJY1jUj1iI7mKgUL/0EP3x1RmkKX19W9XvvDlSLX5fKqzQdc4NP15fIaykn+iQF9AGo8gq
xxLb5FkJEKEPz8q1r4hwzxIW2GcnkRfORnq+auvMg51o2G6VUtjOFaKSskc89kZvflRH55qWyneK
0rrYZ3jzLzQsDdgaGhSVRfttGodjvAY6Pu2KVnZcvP2TuBf6drcAXSIL+PD4uzESMKyzXPziPvsg
2eqD8qlHnEzmgWgvguxHBGGy0cwMdQN4ULudD7dye/+dV/ho16wTXccwxQr4joKSFiQo01GTUz0m
m309lgM6JK3sJHyQOiqYElrS42MqQDgywS352lq5x2bU4+Q0mp6iMUwCxe9hjnGXc5RF/Y7arY34
duYRMHK/QIO9ZLFMh6ILPDQzegB6+3PMFCBFyjDmyduCN3yEYo0EYF/ohNWbAJVq1kqCoq2VBCiw
9anCk9YHpQGqw55JdWef0yDlp0yWesf1rSVeg7NRn0chVOqYLO7x22SIiIDyTpmwECY+4PLJW03D
HFRQ+TxTqa3UL5m0Fi1AP1Y78rzgpkk05Sx8ztC41Z0fSLobryM7tgsdYD0aqupty9KjwoXCqIRZ
3TpO+CQ4SF59Q3I2tp9SGFVX38pwQud6QsXO6fz05QIC9YUcqwLmTEv9KklTGqlpOmGWMZMTaywg
JfQW2rpVcVvV9qfH+a2aEy+L8ESS9ZITrW9ClwN2TOzkLdMzYHfzKADiHXNPV5Nq02rOeHPg5aQh
0rtezLyrac0XztvQaC62CC7OJMgymZfv5oW/YGaPVXDixBIYpcihBfu++3qnezdSGj0db1f8DXdR
JXZQKE93G00OaO+tndrKwnc3H0peYnefTplBJ/T5iYR3+YFKLUfPUSZlfA+W0MS37ZmXczYL1OvR
meGuGQ4IqVd37u4Lwq82Niii8FGC73Fpbo4qGlG75AACeNhTNwSKCAlNPkh1BTk5+oJ41IaM7LBu
60dZ8FB0QdQG8c4TPQotKhof/nj1wHCe40EIWB7MJhLiwIxREJdiV0w+KVZ3n9KKQug3Tw2CzfCw
LY3yURE1qfyEMlO4bxrhx1O3/0Dh6SWXgYkAbedhO/2G20jPdVSIQ/fdTWI2oKFv/rlFgtkGf7Mg
STDbzCCF9m6b0gA+EKsVse3fSdp8AdI+10nzA7t8+DqzA+/qII6Ai8JJYRt73Jd+2NDxbz7HcH0f
3VwUc7rEkFYczTlF+bTgnyO+4Q//rQ+AdefWID5IXajrQuFpugtPea7UuXDMDk14wx3MK6U9/CbS
lSQZEHfI7OZCy4n+G4L/vVbrITpJmsMKQp02rmrJ3etY56oW1yqe1kwgl1eIK2NX7GhTRxJe5flt
NTezTJED92DrbqLH8qRiuO4siUUMjZkm8l+dWU//A6hvss5Z5H1cahDxvJGnhjxPs0a0hR3Mh22j
mYRoi/FjGmNAK19+rRFlvfW+XPwfb08vVrdJJhyJrO1XKcLhi6MwykXt+tVUVwgmwNwtAdw/EQiG
4OOgCHV76GI7VhOqfp2/XJUuABefHU0ZgEFiCYAgNvf7Y8MAcVh4EFWSgPNXJZ921cVP9AHyXrdv
B3Fwwgle/HdVQUSoz7ckWCNfhqS16FI0Nq0UsWRZ+inWSVZSQ2JZWb0hEdf8FLzMTd6ArLE6AKM6
vkbwS9LEYyHtMuzhTGmM3fB/ni7WPssFdIhUEwDbDuK+i29rLp0ZAdoKk5Tcw+FyFl2YIFqMrNXr
Rjgv0Aog0I3g5hCTEVvZ3JSaQ/IkW0GmvGBb4Gm+AmkDerNsZyQA+WhFscd2r4lBrIdv38sAHTph
S0vn1Lxsg8dStjsZQlL0LkEdag8yZf1RBTvgzQwxWNCEUJhNtvwwzHVvTkKMNTUWWuB9jY7dMWkR
WFbiqMRjvMc9LYWQQbu20hJpcv22RLSTB7jtScDrhODM2a5tRCJU6j2miG2kSz2CMl1iR4OsCap3
LKHFTBGeYrQ8ges+7zcI9wX1L5ft5ex1ridufNnXm1Y/RrzjILh7vRvjs5T7CaEZ6a1BrHQ5k/l5
Wp75sqVqEWSeQoZ52Qhjb0S6BYmA3sb32kZ5d2D5zZFj/VitAZhR4j12MEI9AdV0spCbQC1EqfSt
0v663LG7PHvZXFtHAq014Hk1tjzkqYdwruF3Z+oUHQZ5iqx81/PASjCqdkzJi3JGkPWbStbqbtrl
SUa5O6FHsPKKb9TcmD1RTHVX8RVMmJENWkjTPDCr0kgta7bUXNyZBh6nTCaIfIL9ks6nR16MgMOR
QTeRT5rn/hZEi1UeLIdTPFuy5YYCrIuASSb9PnnFWfOOAsibduBTwLALYBoSniyurVTtjNX6rP6d
+XS8pCH7lxHgGpCZcqLC9qBWy3S5v7MxaVLqnQAQw2bUGYpc05xxOW/TcVG8YEE/7CMTQyhNaZkN
2cMelE7t849YC8m4xmrh2ETLyHw47ttSXAhptxLBNkDtS0n3GY7SXABu0iCcJ4/q0sFlj5kP7vgh
zv0KhGIYIx0CAGHHr3tdJTpIP17/kdBntHPAwpI5JEHZa0E1Ue90bc1TVyqGlQi6H0RUm3918l9p
O+y8EUF+RUzRbArfAUj+yOVVMRN8lHyJyTktu809HXoddMFHwjPS5ZQYrpbcjXLBcObd7ia7jOEl
+IkoM5DP7p0JAzDLI3s+vB1ri0MZic8sNAeIsiGRDcnMww86C2xG2ckmG5bPFJ37jkEtNN0IiLtm
goKCFZ+gIEyXixe2HlHcXUN4wnT6oLPxCat0+SmJLtwB5oT4zWzXlJky0Y8Rj6rHvAzKPNWY1jja
lT2ppX3SoBsXEDZsRPjDcihhbLVbOcQQCVMJ2xRwyiYFpHyKfE64rUumoxPEejCQMeA4zZGkp656
c5XdjQ7FgbBBoGP1aIhpcin1/w7Ip97AKwuwntA/ALtElLWHvI+H/KMmmUMY9BzYYrw+c3ddgwEH
S6o6BAYuJGCGlB/CmzNQIJM9jC+X8oRSovoSCMWvDcYD+1pf2ZCfO87h+WbaCabkfBek2JB85dF9
YOeawIZg5xcV1zvmf/G93qN5hp62pYd8nJreChdsS+j3PLqHigbnz9iXYuY05N3k1fdTCFN0VPTB
L5oA71+770qiZhCrpZkkwtfBsl9WqpXzD6/xBwB0OLs43v1oSlKKJIGEnEmZQokW+DWgnosWhOJW
shXWJYdTYu3ZDKho//jOasFAqILtY8owiqknIqdxbQlu39/pWCMGg//9iSPfz8+q12exKJbrqA4u
g+aSkdkQDv95ziHybfPDBL4RuL2Ha2ATsuMGqixDltY6igdvLi3rh0PZ1jIgsVtFx+RPan0YpA2o
jqikU+prKzJPrYx2rtlBpAP/mZ+66Qy+RuTunhA4nB8US8rMT/eMBXW03hF28MlHJ6azpkPJuFod
ouMmmTR5IIUTQ22R2Qh7XNcMYauNgBepx0YWGZ+HRBd4W5HSR4evYrAswEAQdcyMel516LrqLSm8
z9GTlMAmEhAVtapi/XQG55peHAXfvpgcj2WFw6Dlku59qiCWyKtiHMA0DAQnE7epS9WcKqqi4vkI
Qk6TTZnuTDm8DbqV6OfO70Md4gsWRxWimE2bfx5Y06lsCMW734DYMxTAW6fra/tbmTBudM2+3w1O
F9Y6g1sbDFhriU6CWi2qMNMWftrcqMi+Vlc+O78oIE5B5uYOB2YyBHPFV67iMcBjru4q3sz/bKm3
ug6bmeuzZwAdhFgDRH2rZ/zpMrwN8AcRiIUmQoXTcF71qPcCobz9VPofnNqj62ONYY+nSm/z5ag6
P2/tCafvYB/2jlR70LEavqL+2LF2aA1hnugikLxS7L0hjYkGIwY/24Y4PM9U0q7PIPC9eum/VCO1
e+fmHh1bTcxs5+nl/HHRV/6rHWoFVUlWjLmvNkKC0XVjyz0kgToH5I228KQh4djVBb2TD9kqkYwX
E7dAiDcLPW3sD/9ykGXoFHykStEM5sPbdrj3JcDtmz4XWf36vDZyE78xZDdaEAX2rDmpWjIhlbW1
p1ZKHscWxtPqg8OLbZf6rL5rT7HT8v4R/n//KEDL5cJc5398p+6j4QoZWJtcvt/foucVX2MNjUWz
YX9L0i0sOKRP9f0It+tQQ+nLLXby9ZcMqxxYa6AyurgLsaTjDwTL6Io32B29lOGhmmpaR5Hu4wCX
4+e8qvPQqw7dL5uADSa0g2J2JlnuD0nDU3C49z7FB5MvBs0JlrJLkpRRaElqxi+xpj4Xi0nrC69P
qiZzmkLaWEtKE88FX5g5iF46GVtnB7Y2945gvgo4RLLawIO4Ju+1qiTfxRQSRFYwpYag2+mj52Y3
dk28o0ofGrAIPEQ3PYzDWnQQPDUpWO+IaBgWqooZXdS2BLtSmQGNxcPdqiTFKRfllEUj6AfdTeKI
NBBy09sQTNFoBhL7lcNBgR1l1SwoqV3iHpaleSypMW8PUuEYwHnPB3aZLSd+k7/yA9an8sMYqNl7
ph3NaQqxCW9akZt2ciIxpxmDLOB0WpunMfFMXTnYjXJ/mUVUGoHqHAawhF4BbTZCN6OTkj3JsbeE
wwsY8lEBcmApgTLR1VfG8l2xObzHLMp0mECQWvl8LTkhbtBcl6dHu1GRAyyT/AFpEDNIIEiS+SIb
1gEuWSQ8KUB9V2CPAfjs1nd+KyFw7uT1kLyQ4pg4ROu9gTSPecoDZotQmi5KuD9sOYXpUT4LVdwk
XxhVnWHeMOISu4EaS0oQ6IneuMgnP2C7RhoK7bfgbI+xyJBOZB1PQGGuNmwE9XHXGN5aPw7cjb5b
t/NfJik50c8h5l095ioKnykSYBEeVY3NfuvmfcmXF1BvBQNmPaA4AM7ZAewdHI52PTr7+jGXFFhw
5+dlKNjiEMBnymfafgYJMJQS2oYwryo4ygK8ppadx4RZp4obz2mvuS5gvVRELK03rjDDJ00W1jNa
VO4JEgpDanyMuVGKFRl96vIH8x9aIy2Jzbk/l0qDvWsj//ftKazE6kkOrbbtH9hdVpI/yZzM8PVy
cgJ120YfeCwah/kY7IlqO5SZnO0qUAxMdFKSVM+hjajw7E0OBn8oR2a0PSVdKzJYiVvd+AONW2XN
hIlBH/nfEwvctPx4EPlzzBQnw7Sc6MedbaEmXWUTGRwOpoJQoT9uMb6N8I/3RLwvmQAOIz40VY00
4ZGcV05gh340SWfMrLpA2VKdIEeKk5IHTI1uxR0CUuWYzL1Nh6BK/BI5I50R+406BiH92H9z5re/
ieDYx3KVf/FJo5N5jiZgz/6sEb2GaJGWsikWo1ugLbP9tNVY5/vZW4zDdOPzlmEyRHgp+Z0kMD5U
ZF5UXNTprbdh7xINivC/Uzx0lKJaei/iMJSkK0xqAY5a6Df2JW/JQNi7tloXdfLf33tDXOBGUSxZ
D/hBs7AVVeE03zFJwJSzH8u5CjYAmUQvA8pYYxNxOEJZfwKuzpveJBQgfXI/oG8nZRc623k1/Kxv
RZGjxiewML5MhJ7ACzd+oO0UFiy2UWPmv9pZtR8C71PnUtWIrGkJ9HD4NA8bU77zMvB/uFkmUC+X
1DwH3Nq87p460u1zW7sn6Vfix8OJP2ecVqz/ESsh1vY+6dS5J4FiZgTsf8fuBFBGn8HUFJVaFa5J
UIGqSuKVF7HE2HL9SwT5Y1xoLkT7EBs2O/znn4ofMnS4xZwS3YvZtIXrmDaPyjkW9dGRWkuhXssd
FEedT7rtWKUJjJcGLPC+pJC1Hsm8SCM3rauLBrEz8VUVRLkas3pKllOqUK1ORQ+L8wILkairqeDy
td55czXZUHtFtxoVvkMY9pX4dXiVOCfNdD2m+RToeE9RcI3FlmMqmmOzqhn+IytdDeGwhTre5rsD
sgGDdmsLklILh375aWgAQcbagH4Oa114G7nBO0iN1K1v1zB9TnIGBmHQOnP+L6umAUPboIxasgSP
ysYeJhhD5seIvI2jO1HTTo3oe6m+cCMyjfmOWsec3lmW/RImFLW3ttPRnTC2bf2bOXXTSIyA8pUZ
mD/06QZH6mLgitQYkLsoAi41OuMAurr3MmHR1o1Aqjb1psCzjGY80MhK79xJauFu6+aDIJ+jwHZ/
jDgy94iTIKcPmW1QBk0CxXkwmcCY+OiIbf1VDoVBYlPcmAp4LcyDCAzwwseqAKtFQsDHHuNc0e94
5Y9MOS6KHfgHrt2Ykxqjd33D0CdQ0GQDbAUGX54rrvwfti1TPTaw8+H6Q3RcMVqPcXYkkovn9+7x
E/bn7uKdP5uPK269c9c4ha1RlaGaqbJOPSXBNA0NOttKJLw/DZZ+X0nLxN1DLYFTlpGuqGX8eV4E
yOKBhV0LPEwNtvoMFjX8zXRlbIEwAMHgdLWN+K5xrEjT3drc5zwNraiOwqRmWfEidkcWIQf9I8o/
XgxqbPi6HJCZlmR2Hsm+9l1bQ6xAghw2TlD2wqpS9E5J9ACBZaI2UZCx5Q2L6iB+TEg8W/cwexBM
FjcbIUO7KiyDsCyCY6SRIGe2hQ6TxJ48O8OuZxlaF1NGG+bWbkmhUXDW2TIJFFsEXo6iSVRu71pC
jhBwmsHPerADl1vCNJ5MrToaEl75GDbTtpn3tSqlCBngxjQph3x+hcrgw77sQp7oVqht+Qi6ssCZ
/23tVELA/wEpdOsX6sRDIRsE/6c4KAHpj9wpc6IPzXnDX2Q0fVaOdaApJcAGe6U9amKbUCzSQjVP
CUaciMmpNHZXVo1SEYPmmbxVI/ml0VkeM8pHp4IIjo4ZtOq2Se+T+iUuz8pvlqvM2OhWHqtjgFs/
nvBbrsMO3rdYkP1hQljxJZwnm2NJf88zEUAFXrKZS/EZccZ+b/TX8l/SFfDLozmWAd2XkL6AVI0F
7MxgjoTiT9xZZG84v1FTwbd/LB23N9OEMgjAZmorS67Z2Pt1NrlLb/j3UFfiHesf8rp5/kRNILRf
K6FMpP0WsFVKrwZ3wtDNdzElOa7+AtBIM1e5A58XuEx9BVUTP3ZN7oxRQznTm5bU0ad3sf9+5u65
R42zPjhMWG/FRzB0TyQJHPiDv6Gdz/evq/APYDVe8BjjN5Su0uTqLZgRPTC6107ljq/UHV3svJBn
bSWCHMrqziDbte4+mSWjYiN/t7n3qzI4Xy6zCDV8WAtBnVb0dhfdyUhwdS//L88o7I50PHEhGepd
sBzpC5GWmvzWz23bNHO6992IWtZTjjKFcPBvQKzBxY36n9SxKSgEKX/IYz5OepEdLKKl1JY/mzWR
mswn8pBuu3kIC4iw2MUySSc4nwHU22VDFRMI1xJDpefF6iu5ZQ27eJJ4eZRd7xRS7Blui6Pqdwv0
8cWgs9bLeH4PFJMLOWeGGJaVfDK2tsuA2yeNO6ejMIWDHV/zPqGVsu0gZwL0NngLQhb2Ug3xnI7n
9C40fzmlDGN2xJxGooAjd1gdO4SvP0ScXexKJSVDfCIsp/o6qshC6ibm6LganYCcZ234FS/Rcvxq
xnlFn5G+hJO/FRFqF5w8cKeFwI9j8QliVkTD30K2dGdFOloBzft9GiTAsF3JzwPl04HCuWJVTcLG
SpuEm5SGlDG2m6R/IQNpwRETovahPkg9YqV+BKpVG2XMG9k4ulu3PO7v/ni03pvdPhBCyZzQZe0A
PBwnz4z92lgaFzOaaUVlj6pjUbOnKRlsb2vi7yBV5ps2VSotmUzSlTNXTbk3tMPTvl93BjHImLIA
9x4cGS0iSCbBV1edIcIyqPGMNHoVZ90KRG7b8hL6HLPThjtSnlf/eQuv3+yXfOTw9QRJscmVT9RC
oPgCrkyFtewTQNduBo8LktJDIQRGe34f/rQL7jmZsHYLcgeDK/O+59VzQm70r/WmhCK+hKwFmGlV
3fMKAuusaLewfaZESLOgTtlQl+xOGATlLhi0fePMcoA25IKu4wGSFC0vMRFetRbkPmeMEl6p84an
lrb7vRKUZEbgN385hA6C1LVLck3Fs4Jh61l4SDOX0neEeShz1iHzyV6zMYu3X8ykp8ZQ/RyqKhRz
mrtp7e2nOfLszK4PhOfy4HYmsBGpQFDLMxXbPyTlazxaV+B35nigRwucsSdiHSpjGqtTD4W89iEb
buyXCWViTS9EereP79tSPcHU/hpYQEm03TkqDFHxkqHw1gesI3wCMuwHoj4VMi/a8zi6QCWnbf/j
Z/p8Ljr54QR+DRfT0HPlVDa9psyoz7+naMV3bYQNkAFO7WVzBF6EQ9hjBWpezMrXBvGaXMIFfxN1
3cLg1W/Wtp4SyYU5de+8YFZ99TTgIeNOKZ7vibsQt0ybRnM1wEO3xB6G6SU87Gf+nj2sQxycZK8W
c3XoFs+pFoXBP+G+QLv7SzvfPz0Bt3YpukGoA/0Ewqv82aqk1xXHoVTSKAfKHAst3vMcfXQjRaL6
FXSAFwUasyyoJ8pV3PHI4lSIV5s7oMPiKOxCZwRbNuCJDaGtsBhRW3GLAryKAZKRGQ5fy7PCoYqI
Yi47ycUVT7iyukD+6OWFfKDw4igsaOQLj1J6J7bfYGMxJUBXwsG3ugLROzv/iKnDQcXyMB6myyTv
Och9Z0XybxoE8R2za39vQHGGB4dRl7CHx4Ycguyu+WtGykF5oG6tqxsV4oPd/v6f9wIIKjSBXFjl
rrjqQch8N/agGvpJwHqCesYvbs7eCGYYGYq4s0HA61xT6zwZJCnOM2SpSmNiNnhEuILTwFcBhHf4
PqtZOpMcgySIa+9OVB8EfJku0s2QNwIc5cgcsG9jya1txfKhb7dAEXRxWxoiDMeSnMtp0P3CbByx
Pbh3OS2iSr0RXJAxF7jfQBGoLVn+nl0kcDyvlD2dLkNvcyn2UO+v5XdfypiKwwVrj4CLVWEoXaJu
zXxSOShLuEAc+bYSzm/6efsbV5gWv+89rODnzSnofw6EAfQmjKeKhzXM/b491COKMtN5+Dn0DCFH
HPgZPJv066RnB1RznvGVucHOEZLSqbUdGR6ehIKyAcckYjgmAO4S0Nr0K1ZE6n16r/nV4wpFkVmI
2ZiD7eh4+I8qJXirAFz2Yk6eq9eRZ5POh+hd2qB1aBEG/trUIy2SsweD1jeyFPxQchZTWKJWhhgB
5B1I6CxbcdRo4/8DtArHZgZFzKOC9/sFZH3WTMzTUs8dE23h1ZcSGNfeVQYH+vi4MXZ1DbUf+nBQ
219Lmo3deTHh71etHRoAL13iLkLa32t3fl8Y7JCabDvs2RQeZ+2GO23sEKOyds4P7RFgQ3SRx/DU
wh60wbOkm47khi5ZMnmJi8E8elfjRjxv1ouz3SfLToZAly61btEvX29s/6VqJ+TRntYE7QuIQLp1
SKtOdgsvxDTGUTbHVshS5+e1usFIyyr2/1XmdV9/WeHe/ZOQ9FHcvMQ9Uy2wMkgKmNXKfBerpU6H
vpbwPuYvFWwevxTe+X5xR+eL9VoENSB4Uu1jrR9clx2qZ/TKQPYdPnFMseMPecW2l/LZam5SKQb5
fAzAsVL/IKdfyFSojlejfOO6pf4mQeql/AATg4CZVOdY/ckkouG/nIAvyhDEutxTYBRGbEwcnGjy
Q0UnyQpwTRBEXasGodYwYXncB5ER8tfKzVpRXO6R4QmwoDYKJATq2JMI1e6xUM1FhhVSaD358Vrm
CCTrF7TByi5L6U27h4E/2TPsw23nK4lKO1JnwM25AHeL47v1wbPj4NMgq6brlhM3xKxljjRjCr2S
iuf2Qoc4OCxxjKNaF02H3kQFAXqzwQZxrkLALm0PMGYZEgGAqKzBZtF/sc4uvCgVA+CDIWVGuD3K
TNuxEeKrS94ZS1MeCcBAYWNndvOSSpjrR/GUdBbdMdQPDJDVHwvGIoH/uPnP+QWS2aW4qIaXvXx6
Z3aTYj2A5/m05u4dHx1OCy27mKA1YbEL0vbGwopgMdZ0kTMNrmhiEtDPPXgyuwhjh/kU+SLFJLz/
O8AXxcSh50c3nbNuADHuf1AaeBtLpAuQlt3+zRQ5UsL/xISNseSTxF6PMoHoq/t4y8KhPAd+rWb7
TzhH/BiIpESC5N7Mp2ldt4qaz5jwJWcNtPqZZQiDxT6SGEOHLwNtzES4bEO8ADh2p/EtqAduYlT+
VzD7g81NjLFi+02xdMTLnic1xIejSE11WK5rfcmK1sse+P9l17NcQXPETgGQkeC+w58NxYnjNDZ7
+vLGsLDtw7hYEKOs6fTt/kz9pftgRtTIeVEcRrNXUJ+LnjGMTw2rlFKCYohSd2E55Rk8KPnx7+zL
9WWgW1A8p4RqIB6H4fidSPHO7/pGa/24fqAuardTF5ewZKQ0RDiqe2UUkQfHyhJGSdYKV7tLN6dM
MG+748l4Sq4/336+JxBoOuS1mlJCriSM5tLk9NFoAxSfWMGIFZQrO45PHkZucM3TMtmoz7jjkERc
IOep7vAdgaViWhbOJz5VFKTPk2ov3sOVu4geKuDHkwZbS+nP6lfQ9rwuJ2BrL90mfO4kp2VI6z20
L+74UGK37Gmm0aVTmL15PqFnZmwih9RLj7bmizFXAfWEFLWk0ZiixFOADBXr7uV7ysWrdWTRs5Va
RecQmaWAI9SttM8XzsPV/rI+Qkhijn58gl8YMAuxfol0K76iAUa1RAxo3vSP5OnORh3PDk6cBrx2
ca2Wa/72rEsm37xbKbkDDgHPlYXEixNzC534UTSqHsHs27LSrMjWVO+46c8ntf1OSpclTEm04hdg
+QwCQ2oYfs0xUBDzyjblVXhDebZi/TKFC4K5hMyWddhpHmI80VeQdoqfJm7Da3bF3nLFK7TfzZTY
yOI49C14ZGPN8vLsbCdTFG4E76EFAkMPIceYDWfjgVg5T/u5IRz853Dx9bb/w/vxRJhuNzPkY2x1
rzho1vaT7f9JjoYs+WL3V8dZln3qQUzeuRoZMHDNKMiZTXVrWm36tChwPBleA1oc5Ap2WMtogZuH
fuZ32NHuyoWuVkKMoimW3iBfYsIL8XFMbUiOs7QJiAhEJ+i4gSNQXz6skP7m3dItnwvwey8WKRix
/iIqmfkoymLf+e+FLayIRf/cefQYBI6i9V+/yHm6zGrKAW34ISJ/fh37VRPIIp6IU13e8S69H5FR
kkiDFt6j2ox8MPv/ifUq3ykyRK7W9xHjPlXwjfi9Id6QOxTQgtYQeS48LZ+pWuEVMzTLePAD+T1/
+yq3O3tjZcUvzjH3iZUauzx9gbaCQjONNHdSiqiGRZ6i3hjH+sCyPLptgugV1wNIuscjj0I4zyFq
+BQReR5pHMXy1YlUe7UwzBE/g7z5W+AAg4q2B9NA0vpa2MHTGMUCfpGEnP4A0i0bHFPWQqS029My
D8zSDHbxUkeYAIldqQBB+dXZBfJYaYoUjw2BLQf8pRbHOnRFF7O16KDYxykKjdbVlj7B+WsNMcHc
QnyYILxjzZJ4/BmvC6GpampHvhAe2Ep+UGXFsAXEAg2haCJKr765myv7v9h2H+QG2jwMto2LP/wa
808Zq+yEuw6wGTO6aw2ahPh7aNxwOGgIiKofTWrAjfhadk/uKnoizjDsqTi67EkyJxr9cfpUd3UK
sWxNIHHDheSICZtdcZcR2bux44KZqkpqdkN6QzzoHZqTjxg9qQIcFqqz0dZyCBriav26nbcwIR7t
0PAycoXjkedkl9y8jFMZ0VkQWd0JSxAnyTIwuh9sx/bKdrK57HmBVc8n+kEa9ITyIPLybnVKE8Qu
hJuB4kDJHsBYPD5WTTA9lrU8XLA4h5/RA/pZlnyblhy7sr/xqlit48caAB3JSBLHCbAzi0Tf7BiA
eVA/CZ0oMG7Vf+it5bTuEdcDdv4+tLCjaaqckVzb5TqAFu2LIxWJdiBxYzjox/RSxJoSQfObW1A/
EKgq4xo0mkZpcO9022D4yR69xG93gq/WicyDu3fbMeVf2yUezOS8x/E2j+EUJpwUoXdbYca3LoSw
PlzPpUq1xJD3iCtGXBux4aXGXw1mypgKASWXyxcuayvhER6b2H1cX5MouWqOUH0vZuZa/ZgmIT38
8ArP162sZdtmBTy1B66cp0pSb9LxxHFP+BpQ5rEKNR0L5iprbxESGX6mNoE1oEWRfN2Ex7OOWlwo
dZcBsNj9V+n8LCfLiMYg/UmO8+cTtg66pilU3upXCgyPTQu+tcVav6NVBmUqAI1vL4cVeFIdkPMY
WwxnuPnlqwIk54lyEn2omtE6CoVGj1oEsoE19erbkpRP98GAaRfastGSFK271nDFVCaChnQM7TvE
wU4H8BbE41a6QVy6PAX2me/94qgV5j2M7i5Tj93beJ42PgzIT5kNknHxcpypr1x9mfF/TLgCUT+W
S/mHxUXwaa4WfLz1Zubz7kl0Tb0q+vleD949+UUPlNkMFoGrCR2DG3onbO0Dl+GaF79bi7Ol+kQk
csG/lezM5l6KcG8jLsWgEnZctIa9qyBoZY0ShKYXXHOCYAIU0sygEr8tETVVj7p3EBJXKkYKURWY
kY2Un3pvwxik63ccafQPprHWGvrxge/jnKCfQwhflKvw5TlsiNKEbpPTBUzFzGqw3ObFMjOuwCXX
rr+0ZjqKdLJE1rAg5to3im+2m2n/uj4Kjq+nVmJLPDPaPLoozYDJQ8Xa1gANjcV5bV0qSS4jHZyM
l0nOK+FweRaFmGFfSbNBWzRZOunnSAmstFpfVs41pzSkPS2mOR+2QSEeSX7OV41E9aThY0NJKMxz
my/0OULsNxqZrk49oClMS1Ls88J192VhTMN5+kn7uIqdPjJaGMzhtMr2O1V+wCDosb8d2QeQLHEj
SnD5fJ3chCSwfrTSyMG2DS0QLS2CxiOUIbdHWGphJlucIXPm3r7OxIB5DG91J2jJQqFuasKAWw4y
7qS60eQ7XKvLcqYiZ2qhfVlbjDJW/uBqTBAUUeeiau0Eh4e8UugJf19KoDLWLNLwBJ3gCon6jYEe
z9fkTbN9E6W/si5xEcnG/0wN4JfB+k9UUI1RhrjwO55bhndW9sIEEarTdVUv5/6a2Ho7x6PDf2Qc
W/v0ijFFbM4eMMh9IQyIqL7+VjJ3Jlaglq3LO0GJ94HdPdi9BivKUVMfnRm6TcZa9yoRm6e8MtJW
nRkP9ZDTRhY5PBD4ECZM4b9HRdKaA1Kd7e1O/d+j7+qpe+McOM6Rflaj5JTLvnZwDhEHYqBB0SD+
ccql+1cBU8fGfy6c6u5aQkyQu2tERtXU8rO8STRpkjijPodYlm/y4aHs6axYxR4/yCxQm9RgKoOE
/h7vc7sDNGMTwd5VBBeKxgg08niU/0mr3NETgoyOKemB2Wsu8UZthF/E7EkQGhoNY7enPrT8VVp2
Xuy9umSefT1h+9L8CDGfZa+Kftd1TICR+qfUNLYCgdtWGOoO5V35GfLUHHP9/Amqzhb0e5TTm+u5
58Y2EGgWzYVic9A4TDodCpHbtS1LeHQwzxIr9iexL91jyQMXHSZHQS0RiQ0o5GYJQGyi9V6/poIX
DC8ff2IEdM+Fd0Aa8W/AXXjGA/vS1ujDJwdVDzp16e1vJ6eaP5y39GLGhuYIs9pucshXcSBGpyEz
VoDrJbdb4kxRGifUjhQ+EI94qKIaaTOxBEkMtHnP131mJtypO/r8wvbYgnrK0ta42eMrYMilelN8
QxYhC+YZvWteLiC3FC6FBHFy72QctepUC9SdV+rL7TclnAajA1Y+J7f+RjLtIKhfLoglsLEqu4OA
d9LRYyPAfNPk99Bm4Ys5mh5gIPrb4EmYVa47+aqcz2M+jesyWFE42NP1IxEHs/r6Pw7MAAA1YKwj
MeAiLGX7GzSmN7k+qJGr+WacC4HzlPyz6CqzP2DIAHwROdSRdydByH0KkTP3wLmSfePrsSQbam1J
3IqT2USMR/j4oK2+SHdSyGJyE/10OdoczBg4gfYF69Tqj61WzK8zZZbXCkHN+vMBgzA0zrbJ4mNP
YDJJJ0ofBYSMRaKtXb6tYI9Z1+zU61xm7eNl8g2PZAkrhZivns5r2H9k30q3gOzPCzOM/o6abD7/
LQdvP/wRw2Vz6dZfEW4C66R2f9FcAgXNkG0FW56VL3m4mkeZkms8zEqVftOXYerjV/Ie/hqq5eYA
C/iyqcTCnkqah0DfIdJDZ9/sycWW5MxnGBxFeHTgtSfxidJgpGh2qm02x9G/V5UedGGJvJ/kGzkm
B//pu1/LsMXF9yU9KBbw7j/xlPqjPpJEoex8UC1k5oYWgeP7E7puf6IToSzqflGksqyCsvKRHQ1Y
ZNCN3XjYL6hPoxEM0mCnazMCTRews2f5hu4PPYhXLvf4yJLToiKfBAPPxnYGYPa1aNR68bKQ7/3F
ltkm3mXzniqoWyetm1hWSAAfD8vAY3Ghs+SaDPotupOwGYQ22iVsgYeme8QDhRCx0QILwI2MOz76
UvRZOg1IeuYT3qqsd2eQX9ajRJxHw46QEBu9L4DI+6FS2535YWFuCY/6TkNFbnowdUqLUzEWxB35
nvfgOFdi0BpPifzVMzj+VzDDzVCkVb/rzLd9D2uqqUw1qzvwgZhbST8gGYakRRkORAq3rUd+6cLI
wQRD/Tq3y5NbOcp5DtAS6xEH4M8kpL2mP9p+saRnuiEvWKnvucY+0gIDHASK1c+XExI/thmwm6Bd
8MambMOLqYfTEBg4tsNeQAbTPy1sOhP82rTAi2LH789PwXfcA3LblGOJOVk6FlBQT6u5mBG5/qyL
PJBlXYI9RDhUTwSIBs4rC5J23R8t3+TU4Y3NuvMtoI9V9NUIjXfwHyg+LkcGgZWRTgtaRU4v4RB7
NqSIBF1vsoppdCj9WYix4K2nuvlcle67yuw32YvLDhWy9Xr2um615nP/Il1SxYlkcDwBYH/kwVZY
EWUilB5mfkFNlvwC9NIdOpVwk0iILJUBn7cFlscwJJPwBG+wCxpEYgSMgeQntxvGf3hRISLdoiml
rwpZv+m3C02PCfdUXM6MA1IyPf0s7GgyVfPMhwscE3MkTWlWQPbnzui5SW0kCL4zO99Ui49CAsmJ
O9qjF/7ekXrcOjcCy2pbnfYZhxw/9YJLV9nkCbfuczpgAqlioMU4u0GGr3mGCZ+VkUtOY77Aaxzd
7hOiJm9B6yOpHgV6nsg72zs1ETybRK5VIcOOgOzsKyfkuMqzEpsJIyyKS0f1vAD5D507G7z2SCCA
2VXAw7JjIIRbk/93OWVzzAfK7MB0wDJ9y2IObxRp3QRyrP+ttJvH1Htdu5iYZeUj+9HXJlowgxoc
Rw4nrcijsUpTjmI57xGxJ+Ra78e/APtZhMz2ApzkdSIVzQiH3pdEq6qAoHvR1VnJJk2z+FuPBndV
9jthx7H+XfeZF79OhtulLBtto+B7/GBnjNgfVLsojJB15gKTyaUrGMOyrHd3rbeQ5W7Bcpt8svhk
QVWHkM5i5RjbYEl5ZZmsIqwqxxSxJNdzaCauDWxNKXWr0SMJaUC3ALh9f5S6g48dRxUu+h2OeD4N
LPJVJXwU+k9DKJc2BOIc1Fgi58Xl66pCNNzwvbpYMZswD/vPtMLbPfPxn76CMa3CfkfElfGRXVhb
dMXIZD2wEiczDko6839pHApEbSIal0lSELkTrvCKaPCiq29ceTPMGwF7uXG9d6tPDJ25QNAHvW5+
d1nQ8yf0wgGtSOWmkLV2rnzjwrt1ErluIZg8PPgwJwKe59T1j32Fv0IRs0peGavg+LnqRcYBA2ow
LIR+FCLJ5ZGJY+IwPRWvT0R9clMiQxf7DIHuAgQezm9VcTXE8/bsP2diIJ/prvWYAXnAUQQ3ntnJ
4nZ2nFZ8i3q/1EwMLFhaZgHDdp3Fn2E1B5N5/KmTDaKjg5PASii7B7GZ1Zjo1tHUr/B+kxMIRx8Z
GQpdT9rcplJ5rn+710DlrE8146BGnUSG+LdB1jQRQmgfXRND64LR01b7dR6/3AFeCINnk9+2Yo5b
8FeA8QzP43PSIJHkjBOFIAD0M6YSvdv4eK1fEKFJvmD0VFe8a5q77Gk1eapxRyonfKtAcKrY3vkX
OVYXYezpizxRxdrGnOky1KUUldKvGSxQ6JV3cGYs1DejkhbCFZ+yGGU+17sMiFL+jzelxBVUkhVj
La/sVwWv1P+HEDm9iTg0VEPR54NqriJcW9viSGAlwFRYZ1VnxBCvmRYHeemz31QQDuVzJ4p2ar/1
0THOSgpODUa+ikOfX+QSoz+HIRgOma04aiyUgqfu7UXZ2Pi/4KnhpqFspa77d6KGtzD8p8pXCQC1
tKtozwC5TqRyStzAN0IXkq9kl68x7Y2UzOhmn6EDKoOHmfUf0AYdS7oh2JcsvYNA+UdX+1wDcOM2
cfFIIPTfxVblxZfct6Z5oqin+o5lrvqND6EgGeAqgAWrFx7IVSz+X+hNoXfCzRxSBW4pPu80cipu
ir+TsUt3EI7jIpEsoa5n254Smg25f8FcNba9PIeSZUU165PrrOAW5h68/vOcxRGoPwNQWHhPw/BZ
kZ3LqjRwQeAAZ5t8fYt/O4zsViLUYAry7Zd80Fiql45/dteKvAldzJHEDj5ddObssTjMyGRdv3+W
e/Zv9o+dNykLOptPX2nWdG8drWGFb6JeeaTCZIMx9EBoIXmvk04QRfaXf7vm553LDItyTEeU8F7O
vmDLk4CUop/6uvAawJcmI2nREBlw9GPvzKj71L32kVyzcAH48Ll/GPXWw2dsQY/mIJ/aoQNfDNVR
Ya4AJpKzwQ6bNkcNNIiVOoCNoiBVjyYlPJaoCVFQlJnvR6N+KfvZHpT+oAdXnlPqJ+qUjO0iMyy3
TfyusoYkmRQWKYwEFpyQjnBSZRu7hgHJpNCF2Sbmiu650KAyZ/7kjRLOULfL5F4YCCKK2b+Ayrfx
jNBhsO7/FFeKCJxoMDE12C7sbpdIhvpjDD+TMWATqC2PyUpgYj/S9ENtSgmDos0aWpkYXdskL7hR
MhslcFw/kixWTnQrk+wzrIjsNhFyo1n7Yc96r0ZCZ5r8uJo4iBH1N7qKmR4UCflc8v1JN1E79aAz
UTsukljQIEKTWKcK85R7OLZOszfn6Q88b12x8pmlgT3c8H8fEeGml2mrow3YpKKUllzKvgk3vfv8
+/H7AwNHohVO9JhKe8bTSuwASsCUpWSLJHLYxtKXKWMTpgbF+CIqKc3UL6A7iHXHf3XBwOLQIEYQ
pcUVDBsfuTNGF3gAqQ70MGHAU+JMdwYpkp0vyDT1/bJDfnVp7LrURHV5/VaotjnmNbfiRfWA417/
mDFaCIJn9J1TV8IOO2EUVsRrQFXNpiQG0zZjp5EZ02vNntMG64VIuDWd+74+thybPwWMdKRHSsfh
Jp0VlmFjx2fAgTFhZ/Vk4/O8pQgS3MoUWBBUmoTQDwsu4kcFFo+LkNlzjhRI+iXDzz+ttHKv/XJN
LXidoxHuqLmpy3kvvRrK4RbshJVxUyP3Xs9Jmi2JOnu8oodWbtpZNwCz2Sp3PJ/ma/dhq8xOyocL
KCFy6c4/OBNEkT8xVJ5mpmh2rWeJfnbvcYuL0iaCd4Pp5vk5SLz3JoqQHuMXp+NLMOd4uR20lkrH
QPvcCqd1PgcWZ7sWf68kg9s2MnKRkF6ptlCfWnPZEyvFbdDUSa2xthTwPs8PW3EgISPX0d31UM36
Kt6iXzO8zaw2H7Q2+2Op4nNBesaYPS4PD2NpGHpivKiDvxSYyWp9ijFTz48TtMrJxfSbyVc9KJtj
zCwp96mea/Jfnvl1tnehwjMZLcqFqQyrGKQgcg4TcAB5K2LYS/E9kSbnjvggCvbdJ4D9rE2wAYDz
xQF++g8IPtnJfjByQYNijYREJhqwKbSW7OPSaNmQ6wr1yLx4TXzX0z1yGtYMqrCO5KNFL55bCUou
SShGRaSPvofHY6LlmB/4lebmBXDe5UyM9XV2VnzyEQtgeU0PP4IeLc00QcClxnDFQZHyx6npzuSP
S6sUUGCwzUu1E45kO5nLO/Vx1T4S8mzBCC7SJlLVARvnqofnttEOf4JdbVoKa2IdQYnucf4pLnB0
sfKgiaSTN1KhKi+/RQA3BAResuhNzJgIGKjVX+aaBrCLEghialYFTJKOE4VUuASDDY3a25M0wTaT
oaNMqBulYjxhiybBW2p/wJKbzRAj7B8Rx0n19sSfqncIy//MeQbXSuEgRzfWbm/RO7dT/B9Iw377
TR173DljAOt/LIVjhdV2dzSYHUJTQVfMhPxBm2E2s9H/V/6vUKzM5g7Be3ta92NBBuOw9KMKzTvU
eQz1kCXAZLhhtiLFdWUhYg4p0qszsavnZ4Y+528EFe3upaEKvqAgFPe4gDyLLI9Co9PoN5Cim+hs
wKMnBomdXja0WpzL5NttCu8VB6Z1oXvmokW7c96UQrNhlrSrDeuONVmtWahVWFeEnKZvd4VfNcJP
YoJktZKoBN3bu10psTp4SHxqp8Xp2t/Z9fJP23Cd4oujsdAK+oZiGGdmmzuzVA7+CNa2Fs+ruEc+
9nbTN48D8hcRzUuXYtXhUVTYm2cGWBPoJ0BqtVJuYDXYoAzDwBKpduwqx4wB3alRKNDPLVkkcEDZ
Q1A4SB2Kgx2h95TnzoWHU3Ku2cciM1eKyR0bAKrGawMZckziP31acMAawzds9cYHvZYVTV9hF7rd
ssBo6W2kpN6p2WWIclI8/MUMHfr31Xn9iZFkwhErfDJ61hhHV4yPauyOhLOgSkNZBh5kqy/xAY0W
uBphg1V/96jxSrV+WarIoh4n5Q4HLH6OVd113EibAg5eON5UGAllaReI3QbXyepg/w3bEKmVXchD
i6iy1cggOV4gLGZZQ4bGH+tE1Luu+VBwiL0TgBs8nWIjjBFhBHiz13zyH9aFcxbxMLtc+cOtbyWR
DNn8hZTTq5Bhb/Lns7D3hLG423t8DpWbbKcFgIS4rXLwe10zL9n0jeLt6hvqdozdZah4vzRC5/9D
Y4lCKYrepKu/1zPHvMjGph1jh29fZjBcqy7uW7s/w0n4lkSRakW47KeJWpV/N9mTewNw9NAw6IQh
tNA1YJq+2uLa2q1AvalgudUTuvWdjRK8WbGl/Ku4xd3uonJrqk73pdzVaagdNVG9sfFnkkgLdFyN
nXiVGlGojHZoOItGUrn6PxlxobPYn8eWBd6Df6UWMA3s6QrE0HXoE5TfzASdsvPofhdFD4GhHprt
5uslHlWam3Uk2GXthpPxrJ3gf04C4n19utVuWieVHTolNrBnkYjFs79GhJ4X/C2ZAdFltv6Naii2
ndMHBR/loKyb1QxQCamYAWz+kvWP2MlRa3gkw3DDowyU5EPQ/y9xl5BCTo29vKNgLeVijCLLAKSu
J23i0pK0brQnr3ryFbAD9ti8HuPlSEXitw2x4oV5l2GDZveE2p6fppbTMjgKaXDv9wvqrRONjCQN
prOqfALV1kyLGKtxkNfLyHzhBEeZ0ZW8JTBVEtf5MNMf1f1KaEo4oeQPzMm6/irA6eGFgAlMXQrL
YtsPLHqHK0IkuR/S89pRR5tuZa3kuXjXzPxrLA1JVTXu1wl3weptBaWaSSi4erT5i1YNlTALYSdH
n3gDWXtAXSp9XJc0GIZ/AZnqxIMepBz1qFy9ZJT1zPKbTIvOoOsj8WqluGnDi/Fvl95N5FuuJPVh
A2sy8pKJRraoaCLStUA/tysswu+utQUqkj3WpdyIDcYWM5euE3xN0Bp5IoySFyY2+DCxgwRVbeTc
LT9dpPhzgWkofpDTtW7wc01yFRDmLsg7I5iOhUPtnoUlMcNwh9VHKQoG75IMArkfVU4uVLSYHoAr
959t/YUXUruXm7LwxF2suOQGpSr1qTgFjhTawkkFtPp5029kiN9CsbFhTCe6z5d9NrIKLqO4MsPJ
Kvl8LSw9w5Pd/ZR0X3L+14OZV64XNHh6CWA/9Djx8K13v0h99C16+1mKIO46qaal5Tq2tPd57158
AWg/8rn+6CG73WursdI9rs+luukCQBisZgCUKANnAV+nanJHsRl48qMUGxz7n1TJD8JF3fJYvQLw
KxJeha5ADZLHI70GnIPv8VucwkBr0GNReIt+6qLTiEMtHveJwZ7eE3KcHf/Yl3+EDDMXyDI3/UHg
sjiCOpkXzFReQLro+6iXFkki17i7PlKenmJIQAHUMM7CuhfDhGluph7ZG1HhMSntSdsrFrJ8FSqF
sIxTnwM0c2N7sA/aRN3XKO3en3xNwNyn6JMSZ3Ei24QfxGh8Q8hDmULAm+ej+pTftb5IASsXIOyq
azvS3BZuBh1Nykq3H1yN6kWm5yeussL7zjtEWECXiqrJS5MHVCPp/Iu0NaZEXBOkPF6bi5fBNfhS
1BLe4GncQqjyNahvb5hmhBgC0c61SgkxIlVSrGB8TFRJVyHOYyMvJc20QOTKckkWbkghK7GNR61F
TTX8ej+Syxue9fFxZc4gNuwlsaP7Anv6cn+yBwuidWeA9tmDoe5FTp6qNsruCIRohxw0DwpKAmwa
05WyW1XBi+8E5LaxsFjEB1YV+ccavt5qdVond5NQJMVIvH8xKIaLKwu9LiTbSa9bjZMZpz75dnpY
ktPIHfcLWEFWLRAFgJqiZGmRuZGbSR9afdcQ4rw494mTjEjwL+KiAY2Wm47K7iH8el/5kGQmquCC
puiOimd+i50NivOK0s904XNZ0Pe+DU+iuyn5zrU3yWTwcv7akGW16YnVjeAJsEJYswZVc7m8lv+8
2wbua3L///x7jU1LYwmmt1309bW4jcj61PN7DAeta/UxVQNR6Az6Ttg/GeqVAWhtO1bs/qlocozt
XOeqY7mdCT0X7Jg0k0Pl8FABqtGWoa296+J9RYynEdlOdKJa8YroIEpsxRYeaL1I7LPTX9VRASZ1
504ot1np6/KsmuX+AgmFSJF9fs+8sc/ZFYNL7H/xW5HEp11nBBeFvj9ZzajreyGBh8QtqxtNgP/V
qA9/JcfSHFbzgNJUlXVA2YmeiVJH1Urnv3eU/Lhnv8zl/ajPrGQJvQeoux7QsaRjFa9IJKpLmJg7
u7m1EHO7iYKKwKV4mDG7hXIzZRktgzayC9txu1uGvZCL+FOQzNtkvvte5vuD7lWLCnuh0nSFS/xx
LMmLsWebiBqJPAe3qWRnv8c7Z0MTfi56tK3ulNSkJ05JSpJiCrF+cJL5l6Bi3Eanon7kIS0J4ANK
D9p9pcWYLQgRCj0vgxYi7F5XJBoAw2PSGdW0i5CILKOc83YW6W+Zo08xEtl4Xp4zH5xZQAV8wqe6
i4lBhwveila5v2eDKR9nY0DpQsvKPsOtU5vBs1tWYyAeBnnNLle3uCaIr/ADRhP+w/25G067DAAk
/3PvS26zBQFO8YPKlxFjRO2aQ51mL79Yxj+0pVkm40G0ypKoHXgm9OZ1N8+gmVld8znY7cT5wM9K
4RtCWctBQ68j94zC8gKOSL84mtQIPhEl0p+s4BMsOHG8cJLZnM2jUM6hw0nuHkcY+LHP0sfA6zQG
YnYUL9XfjYFNqSUJsykYbwyGVimks6cwHAKSe0czeRRwoJRbTUlxqzijlM102xGpOmrYFjx+Hjpe
J73algTiio5XpgHvv/oEOGL02VasDSLsotDNYEGS4OLl0jNBDpx/VGoAAvcDNswtmrESTlnc+kLS
TNE5Vv0vRYisficjL7MjBoL4+kMxrL/WcsIMhoNUjrA1o2x2JItQThX+zUbOThNqt86o30XFnzW6
3WXVfDFaq/RFDOXfU3yzj7Tp74uE4/vc7BH1rX+xZ6NcUSZr41Kz8iKlJyIVH9hVrIGKpOsigeD9
cwhkkUz0ggDDjwXy2L7EQWtbZgbao68aOBcwkvNoNQSHOZEW1hnaNCgeV6bfcwhpLQzoMdEierLp
g9aaJ0fRk+fm+su8yvWZceHvBvQx+j9ym6qQdsjIAzRT2zQQulV4Cg3iB7+UZzKdFYG2B2feeO+P
Ao0hKekoqHX5jrVNk1qwr9Y2e1pIfP/qf9LtU9a5k2n8MWJlhc9PQLKwnNFyi7CLzBScRpKEQLdm
4VBZpoyaB7Yb8hFSRmqoP8oFRpOH4yb6IseLbzFvnA3n/xCciLNth6roQA3bPur8QMJYA1tEO1cx
m5C3GLfxkoa1dp3cqAEfvHxTSGAkU6hojJE6S8so9dNz+lzxjwuLUZmntc0bPlfLyZkwGCs30WI1
zyYlA3egLIeIUjrzXdd1l8HrkvubhbHyeTG44iyEwl73JlkrE8QoDX0Z2bw0JAqGwb5+exXagu6H
5CGuZ9X/03fWQ4tizWz1yvMrMmaPUUzLl3FGbJd4nM/pwCZj9U82B7ipGWi7Adc5jBn0XnCoyeRk
4WkRlQyPkmtsYphlxGFC5YDiztpMdFMf7dtikjiMzz0yra3YhIuvWe30AA+HUA/x0wablzsvqUcl
btun6z+edRrJI69oLNJO1aKSsBN87gQdgBJSKVA6wsEtT4exu4hBsB7UgBAcxO1ZyRxPFNOkAxXX
nnHRGGU5O3d0oIVtxzaQPBPc3MGcuPPo2Pq63AXy7XwqBAMFXIGfxhwKSxp7oJ7I7N0nhF4hv6vl
0Ky/NB3qQgcPDg1JV2FuPsM0wyTmB+gIKpWfH9KeEZpiPL5ue4aEESyTafH3akZnCu9M5de49XXK
NB9VcZBepNRwlJutEgIqAqv3m4zzEXhWMTQMA37/xoAvoVeO26GsJ+PKLdUJdCmU11Zm3Dw80fkR
Rmi9MIGBOZo7LqWm/MDVVW79nAqnTxYilvFR+f8UVT90kq7iSZACZuvlOdE+hooHOFHEsDm0Z/RJ
rQhcmjWRsfO6qH9lqXf2IOTMR3I03sWPf2bMm0LzM0nk83ndjQqvGjGPREHDPrHIKu60Pg8JYIY/
VX/G3YePUqxlUpzdaP9od/6cKAPCdn7WGhDVtDebWFKe7ggPQQTmgTo1NUU+d0HygJztDxbb+SEm
rjJoIjf5p106y+U4YVPlG6CqZSbvqvPIz/klpFtbhKl0y0x/Vw2n+t87+YJj3iDT7mOFiGs2BFdc
I7b+4j6gaKBw6BTlhXpzuWoe1dex7Q5ok5zitJ6dHVKDqEQlg63ysEEL2sqxKGpRcVZObPPTKRlW
y83uRsv/YjGQCEAzanUMSwda0OmMujDTw7Xkd8an1YdVxcXuxbgiaZw+rI3abIKz5OS5MP5lY9R8
jkt9PZfLa7k7Y1ZrhUQlik0R4alnUuLnhqQZJDSC/bvq90h0Cgy4ieQQ5YXdmRxtbX1sV7xHWI5S
7ViBUZxa0B/yoIcS0YL2ries+188peQSseOoZtTZ55HYYDTVxA94IN17FGHVWFk1ab5WMyrgkOEP
nI5LGuhW16RJGZms8b0UFN49F5t0hpJG/BUa+16c9WI0boVBpMk50ORmBD0A5YF2PymTJ22Jd3PL
F8xPAjuRG0TC11VI4gW0PiRmtGNGDKI5Pg5DN9JfmgvVZD4hsQOBonBmy7y6H3MKoUOHawzCgcP7
413/xAAlJfy1DsPbVbkrW7NF4TNhKIks4mzJKHJuLuB029jDoskPffTzJiWFsFNMK1oH/X0DVrqm
xliglpdSxBZxAGDEJCKy73oH7ogmUCewNnO6KAKRLpWDnj5xZHt9y2m95QBow4089p38K4mgio29
NipalJSdLTqrjZ4oLk7Gp9rtMGE0iLdxRRQfl6mPKofAqrZ+omu22WKdSHxTT5LM/1FTbI9DSKV2
tt7gkKfPwYB5kusH4i0jsejrXTSoGZPG1+cK2alrehSzNg30F8gMvxOi+NgID+u0aYTOYbqi7zv5
MR/0Aj8TYhBlz6dfXfdBPiZpuTDtlsXEXPcsMcuGUlAv+u1NKyAwXg1B6HbYIKl3MzcAsgK295NT
zTpwl9qJi9JKLoeeUTyVtu0glmWFLyKJsmfhaNxBwA66lb/uwjYY8+nYNwxXsp2VlcznEPIL3DjR
z+w2RFQs8AXr/+M3S645Kc1Rlzd3ZwGnp4c61sDy9fx18E5bV73dTVHCfDvQIGTKI3m0B1eAu0Qg
td5hF1SCrPGY6L63KRG9+9JCgafHHYPI71F9lwyHUIKZaa1pPtYY0VyPrdhMoCwYNupLg6uGbDS4
RcvWzKLthOizou5U0I9QHf0YV0gEl8ulW55cbWK0NNRaGdIoGn+cAPEx0G/P7y1Y4LpkZ2i0Yx+X
6SZa/Wz4nylH8RuZShs7FDAHzQzWCXRBahFRkzSpHZROehGq30xKebAOobIZRfG+M0aHqeg8IBIV
QfNlL43sJuB4KwB+Xq4n7Jh3O50bq1/qS6+8IMvsAnqfPJ6vf7pWHjwUjBTripP1h3ekrRhGZ1G5
8dyQEEq9ckEndvacrGkMukaa+bjS3dC+GX/BqcoOb0HfNKqRa9y6BNFd07FVShoUekzvrYe19Vsf
cGfDJuT7M/q/QnLzdgBX/2i7PAERPRLGpRQ6SQdDu9yqEgEfY8gfkR4f5dx2XU87U0VgeghPLn/+
/saRinoEPfwtSXYZB1oL2xTtP1r5lY9SJwsz+DCdCFX4vBu0tuAqjW7/h+fIwrQs8nl3ph5IVUAy
D5pjrzLta0DZGg41gJ0Zii1up/YK2cK7lonb4lTC+yAA0MkoEbnzZwOiY7miQfhGb1xvKIIlMgwO
Lr0ojDOkxwPJ4LQ7cU2c31RTIli7APcut6dys/e/k069OFmkUpvcyVk/+FJ/na4Ph80xhj4T7+Gj
09KY3CTcOsf+beoNz4cz+vuo/cyIPoBR5BVFeIS31NagRvCkxVVaR32ntYA2N6dxBym9fzHzUvuP
2E6qdTOMMjNoQpc+o5hoejO/tDS3LaPxOLS4IEE/S/TOcnjT2vaK/uJnmoliCVaXlhDT9xb7Rw+/
o6W9T2aooJraGy9UNM3hI+5vegbHN9O0r60pVYKDxMRuR5KOKvprEfL6wLCdin+vUDUJ3ZCz10zx
wy2e03VpITUHFpgOaESoah28ezmWtnVMLP8wmTO1fjBT1sU7IIZlGDD7i/at8hQxyu/j9s0x7sT2
zs3lsP1T1JBAoJQ0ipmtylI52ikjDmQfVtBIMWmFuobGQBuZCXs0aCBAv36X7Z+lyH3G+Cxq/4dq
raKLX05tz+vdbc7ycFzt1TYjVIEwUNTmRpNUv+K3oGBcKRh3ElXkEJt2LrXmw2HbTNiC+EvkTo6s
NlmnSeT3qAwbKKwjH8rvE/v/Ib7tqImWYnIO2JNR1perVjU11LPIgnqY+aRQCDfIML6ghcSYkaUq
rJJiPcobt8MWB7eoQW127ITpdJ/8dfXIEEG6BYnfVqUHqgJlhmCZcLEbAaMY4zFlSVaaGNDWfPaE
hU2lXgdQTAV9is/fWjjDh1/DZSzmlVADGvUFcsKiPF1m3ofrca//MPoZWJQgEPoYmHmc2NhH0cui
otV9rmutbuM0BEuwIUz8jJ+7KUkepcFyACjytS/u22mWikRhW30jWxq4RcraMPmNgPclFi0Q74fv
Z9vbh6ZH9hSdDf6v967ehbjuHPgwVjkgEnRaHCUry00bVAcYBwAJs0lpePq3QStg9fU+3IbgUKtg
v69LkiWjjLSbA057ubW67MghhoYQU7mfQtutbEPUCREw1mZhcRAejxmvcn6r6BCq3ALK1Y4Zt+UB
0p0HYEzGav2SzES9fwqg5R4w/WuVlZjY3eBOzw4YrJBLl0PjO0EhUtMN5egvIO2zh8qLxHWHZe3j
2Bfykhm/wjQ6+HU94hwWgwFYVOj4v9nplL7BPVB/hELFNHlH2sckiPfn7UaNNi4UC2SnknnsYJN9
B5Rvprr1x+SjwRD0BM0+HRefxV7e9AgT1Fjeq21CJLIJPs12ghYph3ZnPldxNFwme2ZYnPMjGA7n
9i82pUsqRxffLsul5SD+ORcnqN9UNBAV0XEqnF7ckK4L6ZLAifqTatI3UKLF4yO2ZX8nKjCf53QD
IogU90oNDp+/BoZWc7+RsIiQhQpv+aBrzQcUdZOUslYC+Z885f0oAdiF04pD8OOl5HAP4p+S42yg
CvbZZWzwA3Gjx7JpBXoPXHoNMmp5hQmQN1bdHG7ibZ/ChIuFnDjD++e8i6BpeJz3+luEjoyTMbwF
Ka2aI5/8fbUv8yamW/tP1yatGqFMvOMIJ8pqfNB857BlvcXPCxpnzdNkfMeY1t27LAYjiONcSs14
8xhqEQWgGDFKZsEYAmgiD72td/nRyLdwT6dujPaiMqalR0U2HpEBP/9GvpxNn3KWi6t0bB0QHLKd
m0nHBjjfGu4hGSCq0D1cQ1D9IjN5pTKnX+mED6TgLGoXXaNEM4wGiJ40c2c4Eo274rwQYJJVwOa1
HyzLReS0qBo/H6ZXD3XwaEaL0JgD65oYqXNHYKa0akwuiu+npXqkn3LclOQZ/uRmm89K97R5uOi8
3BImx8Wjb00BRtA7PUtU/pM6Bt+WlZt6OJd+HIqYzCbe5/j/Fw0bXJFAawGClFjc+I9SgzOA3jK+
/Ytrez8tKOg5tWjIMpK+aRtfEBkwIFd1dPq4ZkxFKQj2FBfvINeRCQtiNkE1tHw1dGslEYSNY1jR
/GHuSN8rRkEtHrcsrw5Er8zsZhIK9svPP3hLVVb/kPae+is5jADvJ8rviQNQGqdWpQQs80xROsfN
z1J/g3L4h3A5Ecapkkkmz8NUxgg6CTqJ9VbZy5zhXLGkz54mfcxAQNy4psIpPgVjSVJ+l+BhwJwd
jz0ojgJ8/a1P5JoSx5ZpFOuYoXiMuyAgX9ldZv8/YenVA11kFYOhMYlswopLYlTBWQS9OqiN+j1I
DR3ZQfP4tUfQ19+0+CIuHTMqrlhyDb3RjejUhRJFS3KFJTAwMc/UmNebxUd3ylHffgfmB3WczkOt
IhL7MTFxFtVbm3NH6G0Vnu/JaCYfHok3zeCYDNDH7KfIxiJrWSrJ9U6K2PYSBrqV9NqVFlY96che
YKJmOecwXyrlD9wHFxan6g91z+cojKRGRDPPUrZt3Yhyxx257k/oI3qOq0Pcwo8jGmvO/sysuKV6
Aw7kBNU34MTkTdw9cvR1ZHDanQnXX+HmdJxAJl/qU0iH7+QnSjIR1ydXfMVJOzXWw57OlPhl7S7F
ltkQgpir/WcPIIABh+SBfSBvT+rHH0qqSW0ljCtQ0VVnywQ0E3wkHMocMswkU0PMGhe2pLLfIung
MeoAI7LLAWmbp0EWn0kNGqZQ4L7xHU9q7XNDx7TOl3F+B6GBlqS1g2t+iE6QIBzSBLHwpdIX8GlR
UfKZXzdG6iFsk7SppjEOi0HPgn26lWRNr7R9zTaSU/CY0NLPbhhz38SqWFXYEYHfmif0BWHlMtSm
uam9kVrTZcIwv3ArqeAofZDdFnoY8+geDtMMlWBIVyivi8z/PChaz/OdZdTpiNQ0L7UtZj/wuC8F
GREsOrp3XzEck/OYHA2RmiIM7JjpwmLFv7MpVfsLcgqbSO1SWqbbzw4PeWU0PPUQxsiwbXaYJh9g
hCp96jpdKn3AaxOMEt8OoUU9x335kfqFbuZOXXRCYN50ApljbYYs2w43dg4euqWumisG9rAmeN4H
Z3sCXWtVy1LhXWUtJ4k7bHOzRXPyw3O3QnwCoIjH1QPcmlCw+1x4iy8Jv6TVgI4wpQcw2BlrpQXF
jXAgGqlmkiHKrEpTUrK/cF0e8OZBC5awhSOhgqlzW6ezuyi81ZGEekdhdCcJdBiQYtPHblYXstHS
MdHYPNpqPIyCtp8hHPyJFAzEc0W1IvAmDNrUNfkG8wTQltWdy7Z/gd6UAf/uKe7wxc24L9RC4rjg
/5Kwu2edxiv3INqCc79XEflPQ0J789/ImFgFa0ds0+vvPSh1bLpFQeVsWVlzAMXy1o4iOk/Ufy3Y
oFikcSSflixYv1arV+KGGVxaC0vwVcPTxS5E6aH3eqL9QH9lpDqGGF93R3JDHoXt2d3VHj0DB+6B
ZtftrRxq8JdjPMYuNFUmx6M0mhdAnL6Xt+8Nr8jA8gGml+IOPv9nHhtGF96DDiYXb6G9E2IolvAL
mfagHr6ZhDM2dcOViIHMxxZ1SnGo1Z8iHWk1g8KFgI5xsJOheCCh7HBCzEjTm2/6ZUS5pgJDH40G
REChi7mQ/QMkPFJyY0ihx0B/X2GDEfRica6mlXnNTct16Bz9SFSCHSYOX4jY0L+S8wtUBTVNAbFX
OuzgsKiSYS1wPFHDDpN/D0T9JMhi5FOBXU0cFjwd7goizrx31Rc7z//NoQEO+qn+sjvhZJFJxB/O
PRGD+bfDhgfQfaWbIv/ZxaRMTvMIeG3pB5bt3TSFe45Ov/zydAhjwwTB6XHeLRt0fHkQTXb5xchv
B/2tXWI1JPV2dkgzzE5fnnHxc+qsm30FFGBJlxN/1VIix+xl3sqVHl7JRwrqhYiRaV0NIO5t/8gt
qDqAapiduh2nJt1CscDSrzAXki4944LZsEhjmx4KpU80WiMFGXDM42o6KvZFEf5488fd4WaZNQjX
Fz64cODQI0SVMiLZH2SmSAqQtz0K4TOce8yXuQplRhZ0BTnF/ehVP2uPjSQQ0apKHsea62hfZ2Ov
WPsFiGEznPC2HITt0zVVsu52DwgENyCSfl/iNLIaM29uL6ulnINmhWfSAPavQQfz1NTbKCV5nUi3
MSj2Uw05j2udLhdNc/OueAaw0a2X6MzmSaCxRO2nOM1GD3sC0XSPNauLcETXtA7/VanjPICU1wB3
A/E6/89h1FbKtwesT5C7aTj6QdySvUKX5NveJ6wGAYl+LKPHq2PPqz41uTN6RcYSvDsibe5E/AsR
jN54dkyJCHCUquuZc7dCHBtqEP4PniFkIowGKsca5Nv7pC1/oBkwdLMb6uslvPWP4Awy0BH2Lwce
oFTo7upToFbSGXRAq5rjtd/bZAdI2It0I8ZNBmh97BSQuUWvfeS17N0w5QEflRh5ZI62R7OMYPQV
t+vq0MSkdp9hoO+SmfKRZC/DLj+dL/KWXrv01vx0RgjhU/5pHpPCYTEidScAL7/xYVbTnWjZLWQi
Pl9sebE5eIxvV7rXfEjK5Dykh1r59ZW9sn7I5yQ0LmaGWF5ifoW4tbF6dceW6qq0C9y/QRRxq0e8
Roewkil7t+zb2TUh14WA+Nm7EcjQgiZlYmo3S9TZcOyuUmVzppxlPmlJADc3mJBnhhMA01cn3K2A
yWWCjLrbpRYynsN/Ge24SMKmRS1mCwGFrpJjSAWjp/ChWwH1Ck9DDNd25jvrccgYzbUZ0TcCf8Aq
kma/tuo5CP+PQyGPM/7uYEOlopthARDDHSsRfuzZcoofI0FYaU3pKjq4w7DLiBDrhgx3k793B6x3
ZwwkmCtZjMwBeeVyPlUMplSgxLZ12O+StImCaoJkY3dCj87z4OfN0UvuC8wT9nLYtkKfQJTTFSun
8dpQLEEW8s1RSZUpyyGyvn/F7Qs2LsPUM7pRdD8gE+5vjcOLGKkjw9Zm8Xwuyb3w54JGkJJYrbEn
cMb84onlannvx7ExPX0eQzR2KydfBu2kvjHgez78CbUNo5QDbupZeqf4OvmbwRlzbMBNYcb4dPTE
dzv56dOa/4QbFSdum8W+1MYJAre1XsO7yZkSNvg+rBFuwoEv6jVWvhwDzUCrK9TMs2BDmvVqvHue
7SQWLQCWSsMT+tdaZxUkKdtAOO5B1EG+2oQbNDv2/KAjIm3JNl945WsOB8xTHA0vIx2QS1LF5Rp2
Or7PAMCrrhm0xWNVHouQG7jjwXhzkPMpPsi3vQMFy7LCWu2UWYswA/sugB77m1sLpY/jOXkDRvt4
sR0ICKlZG+Qh0HB+BZ0FLyiqbDKxOt+VRInURDl5EfgzlR1ylU42XvkMAjyke2cBGAe535u5OP1u
VohlcGNaDZrAhRCCJNyHdj8VzwH+wKYBUDBJXhmTTyGb6Cm1xx6UhNjm2F12+xlJYsRqTKj/DZm3
DSbSqBBemQYJYB+hgzyNpCAixsYBMfxmvOPfiZrCol02u3HVPOGo1ySvo0EVZUJ7uj2mdAPj9HgB
/g1wTCjyKQNfXgO2Lo1teYMIoENOQ26h39iHZFRcRsBtj9E/NRWMo5eWcxKNAJK9rUVxSrIdUJwE
taSR+TgF9yMXBu3IUbz6gs+IQS6jwSWMfUunMdD9IBZF5pwgiFYYkdAQJbHX0Lgn9snGlVvB1wVs
8+DpifXWem7K5gLCj2lCiXRlh4WjFAVWDcdCr7v8VBt3sTVwKOdYccbmJD99IkcBXWluGJAfmMAq
MBUTEYFK1uRWhd2RbCRoxV2jiUEsQrD5c0vm9zJ0lZevzd4C2c5Q+RjA2zg8chUnZoX2LVDh2x7P
Zhb/m8v3HJU9tkOafupTxQfIXNMba/bueZMFqAiMTw6Uj951Y4Jzn6mjzMyGGBz5wd36oVNAy5IO
dFZTqLw920SZvNnU5MfGT96MDqfvPUoqCX6OBgExSfB1o53N4aLRIcWmF2bSCvu6t0ofI1ND70EU
qqR5B2UlwjynWIC/cgLjvwI75AwpTFishKGO+Ua/9Et29tKuTcTZdt9/mHh7Kr6Q3RfEWYolP4r0
VMSrrM/GtvfgQNld0AxgaMuD3MfX6DJ7RCGKW2TWhCS5c+KnJNm/2aINwwuZcqt4DfvQCdnkHSlQ
hSwggSRoTbu3rJDoVpqz6yNPzkqYlxKwfreQlJx3pQBg2zV8+qJVWA2wWhVbeyzQZXmZhuoB4tQa
hjXoxKQm/XR5KS4pGtC/PmqMYsrFfeXfBufzu68j0E5Lh8gXa6Z6oLEJ4TINbjKYeOc8HfTKat8E
cGyhb3n9EmiTHDV3KgGpvchtCnuGSCqRVN5dfPg3HGEh6LYCb2W08znxG5fkGuF1g2heTiVl/44o
n67SbJbyrvV7lGJzDfcwsOXp5GZnI0QtOXn4dbzanxaDkZnp9UAaTSgvT5RPQ5a5nAr2goxOl22f
szlOwTudbcWRgK9iulhSQLye/1jcQ9BHOO5nh+OW1f/Z+x2QLBecMcBiTy3ESSAJoQajFRs3fRCP
yiYxW+7nhYs6JgJ6bOxBMWjAwNb9PGQMnz6n32g5M04U29v+G0flgTUaszE8BICyH4JPJoq/cg6D
YbIKJIZC4s+mTrrygdo9SHHi5wxrNKJGjBoWvJSCI2v0wTj7q5nJy6fq0KkoQTcnpXNAVuEeR2Zg
H6Hc85x9fkt5GWlF2iE2L4JOgD7gx1GM7S8aMK0dWV3nlMnpzVQEfybMCfgyKuwWrINWdcBMC+Tb
r6hQUxfKUNB2Irs62jHEjZDIAgMUMcEOLstrfHbw5+YziqZNtRo8/Fz+4R6dypjTVhBJxOTWnb4G
7zrwm0Eyh5mGxUqkxvpDpJnuVi/0UQisE+3oi6ISCBfKgat8n9dKd7bRJazKecVIn7in3hPd0dBc
Yh52St3rZommdsRKHO5eSSYh0thSU8urhLOsBqpZQag1SYEfatqOcz9wF4S5+YJym1SG2VBjfLPM
5tCjERWQ+/Zg2cazMY391Stmx/v4NPAhR+A2ReY1SpD3zvTkIlF0h7mbjswuh+v6+a94+zRdIw5y
69S5azBuvLmsEDixzEhY3/QrW6b6/qJUegJ+A6d0yw0diCn/b57oxN9PhIKyPOPAJ/WRDTlE1Aim
cn+vpDo3TgC5tPBI7lk88si0OygPYPimhu/KPv2h0X99pRGsx73UyWcWU5qtyJCIkDrryHYMQNxB
sQK6C+g3b0Dn7r4bJVW9rkbFdWMay1SlkC0ZDF6TphhM9s584ynV4qNxsyxZchOLYF5atbSAXt3h
cLXWmxjDMM3T/FdHjaTN183EYdOVvKBOOj1OJxRt9ps05Ox6mHq6ic9J8jaPoRzKXIZBZwEMOlCO
RbGsZah7R/n1BJYFZV30FndtKTKDSgbqzQZoViRyZ1TmpdAQ3tpu3l+Ed8gmYp8BecYIeN2MIUvu
82lYMcKnd9ajp4FKKWRnX5kuy5kBBbYAbBBkLCf9igbQyLxpf/AyIC3zgbgIg/HTCVcy3anH9bDh
ms0hwt130o/xXi5QVyjBYNvbLvlQQhiC2wgSGnPFZq10JbTR2l8fPUwiEWk11/kYrLih1drj9vk1
1coBV/5gteuwEPl83xY7asPk1Omxnpkgyya575kS7xufJ6+TSSyfkxVfIi6Qjrv+xrCr/yWBCdWW
1AjZQKtvCUidSVXS3s2q4wVPjsZ/ug7kdXsZLrcexSc8Or/2qL+stFAujC1tNAf4bs3l1TbjkPcP
rX/609FA2+SL2WpE79t7oazzqvZgBoTCPe0cq+wz9WNSnm+bvPHbUTnpztnLq9Xh6W9WiOdrPpgu
Ro1nmrpgUSo6GfG9WzmHYBSNEGyDvfxZ+/S1rND+Ye7L2+3SO2c1VNSY8pUzDctz8BGrN50bfH1t
DZQGaWHvphGX9VDP+2TecD5zt0ZrK4dVzeJQSp9JEoVYtxITjEWuR84bR0IjkIm21hhFhoMFEJLD
KfGf6mtSp2BFgOsb0FyaYe8bjBYrUQg9mG+UX01+Egbo8lyk1Js5rd4aeF3EcfdxT8uji6aLhVHU
BMrpLQIdJ2DMCOpeq72Uhh7sH8dpDhPcC/vfA1CkrNpVKtS9SJp9WNGbbbFY43J8LSZZcWOnZ6zU
BtRmIEqOJjyrrgwjeIgiid6zgbUzSn6mhIwSKt0X4GOlJR9KAq0dhKA/2tmkLXtYNbDduxJi+Hf+
Yc4U0/RQx/v+b8VsFQCNobNuXRNvtfKiZSt7iU2+Otk//3TBoViEl7nM+JsIqbaFyJFX/bp2ojEa
0wbMUVaTir3RnpulGv4aGxKCdGrUQpehDjFOWbTFswn6hjDzgIYnRMQEBo9BYvNft93AoIjhbhJg
ZcwCjE1rWN/FAr79dwSaPudOllv8ndH4/aTRKVeOWj74grwgKJYQTO0mDXygvf1ILGGEMqEihpsr
UG3d3DfracZ4/Hy32EqOkShDN3YVEa4PZ7KIjKhn+sw04nPQ/a7EWInxu6J9DC7ii8QYJp4w0Jx+
xwVvc+WSQmSQ0ByqxRqPn1dhVnfq2Dcj5wqMdKKHeETv9GdDF3E12d4yLihyH8BF3a3z7KvOlMtK
HUPBj7QLj43KIt34orIdCloJWfKo5Dex2lg+pyp3WpHJrkc6UufaspmEgeqENGAkOk3ep6vxpXvp
mOZT93hVm331aAzq/YcMgSQ7wsyhj4tmXsO8T1vyuDO0DkZrsNztLNSXoQYRMVGnH6buHYDUoghl
39vehUXwInqA3RUmWr01iGG0Pn0d8F9OrYBnLE3srF70itL/FjYzvczAukjQQwHnurE6xOv1ToY8
apMnxJCWCimxrny1eoFX3s+bfSI6TNyqcR/G3CcvGrDRi6gW3fO9oF3V+n7qK+WkIOZ11SCsp57/
AfzKCPDNjq0GUEjztKpeY3yF3V94pkX/Gzp8JkVcx9+C94d3TsCqC7hTRLalFXi2rVvGKuM6TERB
LlpErfpnvodEUME9mSUVt7+JVy/I/sFUnAA+vUhx6DxhbLfOyfNuN/OkUxW3U971ZqSJfnOm0oIR
crcktvXxGCA8PPxzZirCnPe6HKjak5ivCIfvZXn3BXpA1KxwXbi6FlWpO/2J+MGS/41h2RVgRw8B
ukS73gKtu8OcBwuqKJ82cskngAg9ZZhf/CAqZK+xi8pcikNn5yE1UvftdBRglI9FRUcOZHlRu0mQ
orQOOlETv0/QEZiVASnmlTT8XoToBhzeuBWdwOL3IqFGJi2Kl5brRViAQzdcfDft6/T69HengzBE
JJ7nHcltUGIXlX6UpuiJYCGbFspgmSTBpKGawHdBfwr4xk3AaClV9hLKYWv4MBwuOimGC3jlOTBq
SN7QkqQpQby94akqPrUvlA8Yf5IKqaVGdfLu95QB1wyzchwQP+ea9pzSarPXWjHPb74U+D3BT3p+
0dluBhnm+KG/dEJbBnMKKiwo/DixYQRBpW6TJvc55GYi8qpJVKCRZW1H8bxdgh4K1alaqVHssBzf
6XkVCbPHrc87n49sMl052wb1Bp/ViREz5Fny8DdWrTcbVJxwIaix9AIgEott6U0VSTIxr7kCP2fo
KmEX9tHV7BD4mp/CNA1DOdQtirddbcGUOe8z4fchult3RkQ8qGAKrRluzAyZ4vfplUz7cfQrSIzB
eKUQtQYD4YcEf44foe+cLa54Uv9Mtnx2AaiobDHs7hyx81PygFjsQfVBroZvaj+3alrcnDOCXEI3
io1yCJ/MlIGmm/JNTLhZeRC/10Pl9rClfvYI/TOJsP63ZZ9ampcs59U0Y21COmYsqont3JAsihHQ
phStVO/yVRpYmlDoEdtnLf+x1e1MuQnxozyHC6ekyjd9k20bq53FBF9qvk88OSV+Hkditnz17ZtM
Q/k8iYJavRtYcRz3sFSZ10s3EwH9PfmSnfyFk7zjbmw2rwkkc9WnbyWwIwbFfvYrKjAbIcdBmHs9
8/7sX5QJQH6tUDyi2wp0Qz0K638JwFUnGX7xRnsjFBmsFAgpLMZbq5sUYQy7UK3rx8+n0f6ltFwN
6YJiN6Yhzzrg9HtsXKoxcX4ATlkMCiL6VhEsbNTyle5rmvoXG86O8oMSx8/Ic1UJfos+/6GpIecM
V4c+5ANKVZGPUg/bgDfV2qhWl0kwx0AKAUt6SZg5knqHKzcn1K/4ARcUgyH+B2cT/LxJG+TsO6s5
EDVNCmQ+foY5grJYBnt86Ts2BEwL6r03wuN/mbqwEmbQzhJvuqx/71ad5BsiIqTExshLEEcrawuu
+P04yucLkay1oguf5+x+rbZBjd542pehKbOOMTXVJZ8IhQuyFUlPvd6ENmlyy7Mwq87kqx85DgHF
fe5jiZELcedRR/nfdRA6JtZRb63XTLpgb+SV+W4Agjfjqq2hus37fTp2cW5ZAqdeYETezZrKI3pk
wfyhOF6yCkXk5OsVnvG25WxJDZph9jnqhbwGETbSFijWMU/84UAIwdyEqbR3CuWAPWmw0IaHr0V4
quRIgOlvI8w2TVT0WXmbP8dghuvdGUuUaPlpY5H0HET1dwVzU65mm6a2ADIJoVZ8lkRKFJcgKwby
5mQNnA0S/t2Kje77JiVMQD/2Qljzk7YLQUHzTkMRXbW2w4MRcv7VhQiAAsBDgfhrhARHRAp6QYdW
N6zP3JM6n24pXEhmMaZ1lTDhoE0tbGXY4EvZfJ/+hke58bYZKnV5S1m6W2LMaJync3ef1Vfi3d1y
fRBxg8OCFZIBrmz34R0mK5+K3aW5Uw/OAgRX/b2ZD6lkS5032kXQrSQkx0GIWiy78uTVdnTWjPV0
XhoJHpx/sraOipWOTuzHGmhKrYVPC0c4GlhDdLtwX0SVnSN+6/QpsGTDhfh7iG1xNqoVVR8T82uh
PWTNdADFOYuspBJjgRGHRjOYcHfwRB+oCKH5vn6YVLtOMm/LKAg7LQQXkUYqN1/KVgTOeklaNdu4
MmYTTVNTgKvWBfa8MAuShM5yUBlZMUW/aHsHrNrk2TE+FZfimpjL56Ok/8XzZNO6efaOqa2ss+Yh
nz9bLrUcucKXzV33hMymn7KtzVJTUV14uCajzDaQxLZvL9EMcPe0qgxX+QA0rAPRT+VIxjoEw/gf
hritVuTRv9hW/Y6fFX+BIGL8eH466tw2//yJPXXjSMlo0AfUhbO5iaYF60DlW+J1OvRw0QohMCsi
1vEUeeRxR82LEfSrrLGv7mV4qx7AFJmExBFnkRdiTqix+UdBIFKd4y/C20xk6/xkQDuOSBv69f1y
MVwndzqtmt87jwaqsjzlPiT4Ub/m+gKh3XhTaKVKEfRFSku3Nd/XGy9gHxMO4mjnrfbqkNZfj/kt
j0/uXhzGeAagEfSfwkxAO4T3sa8RGFvsF35/jE4XE8vSk1LVrF1HMZNgDPWytyv0Yc8rS9Vhza0s
T6qrjS/BkZFQFRQLfbVZQHg+5gPwhDINZAOFcAtbjcOm27fAfkPiT7Ew8N0yP+0898oyFN+ouOlh
J9GVhMQKXH3d7A7QIiOit2pSBUz1wHbnU2HA8EtPmwOWd//Bgas285n67tihfNGDfeKqUYBwx3EF
zKk57R6Mt9ymimUNe8N5ja4iuMF44heFx+WkUN2Vl2ztyxp5PRuPLOFy9USwYWVt7AThJV5xNiBJ
UBVc0ikY+NQwltLp5aF0rWkdTT0Q93NMEyxyvHn1HWgt8S9xaY6dzLP96Sn3YXhdeZOi/D1xJdoC
5RXUMgytyKPJsfyKI07tG6Vd1zB3dmIrQFG1kVooQ3SXXZOACpPl2RY+24MbQFidHVcr/+RCpMxY
oWHuSVzTWd95J7xdffzxSFTSwp6NUrf+gCR61HiwgqLtuM5YN4unHNnZXW0AXrtYB5unL53+jBzb
EpGMvEnkanUTPTzGkVMZiIdKZ3MvU5foRNKqTtTJTDmd6Yco38ZIGLp8BL4pM4aE29T3nSKEEADA
MW0n8ZsWlNOcp5e62NNpmL26Q4Thx1PePBrqvv/AnzK1oDjGZyjxGhDLYmbIAC8/0IJJzKY/Q7oc
JYhwYLgWUZmrjOm7y0qeLGGoV8JLzY5Ykb4iH6MsLE/VpgRJ5lNvT6fQjPSDESusLCvyZIoNFsU9
1XLlUlRTXleLIbjwViFFiS6TpG4Bu4atEuIbAJZVpM618z3Mh9DJwzX99tQGlanMzHxeAu2UmrMO
9k8xYbluEfg3KV1fWPxRuH7WbvVwYp23je7ixKMvIzrPatVI9nA3KGK17kr84c8n7AAlP4wxbU+K
/nHDtTAZ614Xw49URSRfX+3RUPyryVkkJoQXpPko/pDE5MKdtlGwlxPrOXPKTaI01LgKBi//hu0D
LHV4RPqYCg6Tcz7rbe1DhJ+J2QFNMe8LV0LuG4G5LH10oAHhxdB0p9Fhs7TGLjRbAFALP+SU2I0y
h5PSMoGDM8EQKj/NRe10XLmcFQBiybmas6hTrRtoBjwROFsbo4gJSP1ei/3uf8EehZgDf9frL8ln
OcDxcJbcYypZluwOFWcR4fBowxJcU02sj1EONYIlGoVNPDk8gOlYHD/YTZbUWPX5ISDkDuktE9n6
mXfWNoQ0T8TzWvwHg0N2IYkSTJfcFRgHpiXHhCO3cM3/A2IjcmB6OrVlv6cU3+Yiq5GlGywf6lq+
Jwt/uSKD9F0Vuv6vm9OAmwkAFBGB2kdCqmK0gTe02GsGuXUGyfQwVOAHlmygbNUUCcZC3QyHQsM9
htaxyHLnlq2LGZ35HGXFTb3h7gmrpF1CIHVXPY50gIPz1PuVSu5izLGqjQizYpclM1dnSwKDcrDh
bjpE96kyD6lpvUsnYcIgkTw9hZyUFuTPH5Q1fIMSyKbmeHmYDrz80SqlAYAoxsxQBmO44S2FCbHY
XcA02SfskzAYpQwZm4lcw69/6JgvwGZGnfa6dgzEs0uSKnYplrvGiMiBZo1zqbQPvnNbtYT99P+b
OcEWMynGm46td8fxecJDgmANclCYzJ7ZQk2NBgW9a3fhFlbcIPXSZePyjG/CiSKYJITfcv+ydztb
ad+lXPB6+R3xS6JrTfx0DmRURjU0ANgK64uYu7OTsFnE0j6zum4tsaLWc3+oGDSH7VfzbRz/p+6J
NhrPdAZdAOT5QQo7qYuCwoKCjFZJ41qpZbbnFUM711NCoLGXc37md/LfnhxCaFcIVej6VYxt54wF
JwCxuWMdkbh6fzqQvAK3G42eJIbk5vpfyF+tATOzyx5nW/2/DS0ehPX+UJTQMWnuaXoPpJvhxBVO
4p53wRopUpVKgLfboxS3FYcNDftCknBbDDpYrfeQgKbJyI3OnoZKl+CVyJ1iAKXmRVar4nXEdYir
zhar/jOPd8Dxrrrjf7x10DGVsp2j325UsArGGaFJUAbI5j76paC/HK+p72JiWjL2cH6x4GalLMiw
0ioHjnSPMguVHfH3Z6be5VjBjDfGJF1XAAMlLZWyu8YxWWo6Lh6u/6gV1PV/iJOQUuK9L0nb8bOo
Qs1uD9HZtSCMGF0riwqYWzYejWr4sFs+yhvSKgqJfPTB4CBXNs15LdynTwTwkWmagehQyYjpJKmK
8I+3kYioNWSGCtp03rzezUjZEYGE8NZ0zM0sksqjksLyRuOMQfbjcSea8uk6QzOtm77XrxBS/S0e
zPCEQqCy36zVjAPqr+b8OuKX6QcH/ThmVa+koRyPujl9WlG+9xLRajLoja+s5OqiRLpTFHg9ydn+
n1EyqXNm300LdBLzHnO/1CbGsPV08jnW/jtyMF7Krqz0QHfbwfP+v5vdFUbaJBv8ioARcyGFiYL4
kAinE88XADBxgHfiK8owAQ0Fc5N9BYrD/QbIgaTKEseM72qyoaWiSiJSWFgssKvMPcnUthVh7kr/
cza9e/E7vbDviUh5AQTLZzBREEtw4tAPxCg7KHbPP3NYoY/PDKguFMu75MJpw77PZnTZxnsP+FNJ
9RqnvtdedRR8U9k6w9TXtB24CGty7GFwLuhv26Xn0knDr+HReACMXYdEikmLBcGWJeYXihjFSAw4
RvU0tJstLhKO0DlX67ARmekAX3PzEX5oHdxsLaa1aaW2d10VSHpJHhQg/L1hQyd/g2/HCMevtsO/
bkw/j+Qr8ewfHzkoE/qrW8IH5IyzanMXbC7k5ulyJ+0ot0zDKUOQKlOdeem5yW2lO6uck4xnD4oZ
Qk2ziUDGLHIqUQsFE3ym9U6nNdYxWPey2VcTwimjXjq+e1WlJztFdl6F1PJQS+6gKQ7xHsRiBcrZ
smudg8nrF2/8v34cr1CuW/LGJH06V8DcnAAZazVph1H3b0DtFYt0E5xMtfSfq8cGhDdooqa8KcMh
GRXfqn4CkW3D5HH4ksXkuzdfHSzHEmHJGNummBPQytWhysCsuuOp6Hu1vqj8AQMBBU4fMqog6iuG
CRTjffqt4cX7VQSi12eAudDHRJv2dJoNzoBx6ng7+oj0Als5u+QG3Z7wM1BQ6DGR4wlzEpyyNPXo
mC9E+f64l5Go8RD6fd+owuUg7xMH9uRFDxflUgpMcB2EoVcCvBKuYpwD2PN7r1wbhtr+BwhVis7m
/dkXQO+k65HaUYhotI0XrsQ0JkQrVPsgGrinShd1yid1eF+DcfnYrmLuz3eJHhUjUeEF7u1zBDy+
YRF+OzkD0MqmwK8ldaNbLLoz+Qz8LWAY39cOkMj5Ul9eLGL9P/YQZ5E+cY/pCtqCwzv9myVPZ9nC
48YdsyH6UOQij3+XfuHviysip412RY+shWtq2IdlGjRPZ9/EBF99KSbd0jd1Fg6cln4by28hXhmb
HWwJvS0vPgkbt23bibEFxqAScl7GSyhJH55uO/EMYNM5Rn+8qHg2tt1ifHfhLOWAs2Jc9BCWwRna
TUii8zfak6GcwZm5mZ5jRdvwIKWcAhynFwXS/HdTcp4HTQXwGHecaKft2QxxfRShWrU50LxsFRlz
jZV3Q0VooT66xW4WGUS17akNv2aqUAZWTB2uvGEmU2gY83cn4vVisS4BdM78/rDa35Sp/c2lXnTx
9Tkgw0cvYmQqd0Xs70qVJTRGGfI6KNWrAH1C1MvBcAJ2NaX3P3+yE2+8jS9VKMxwQQAMniVBxB9I
p425zaYHw9Y08wNwBRLt4K2b4qYMt/ALMwcG26vn9Te7skma0JewItU2QWEJerv/qujTDt23FtOU
zALZvKDVCGSESj1rnfJiXasOMgIIlCAXsoSX+FWSucddNKSTH3Z2Zuu917pXxGXBBsP7ZDzRoZ4K
DROCR1uT2P/YIa89jMcW8AUZ/liRpLb8pT2rUYqwWlfovvWE90YSxZ2kcrucNh3wIcfHhbEvUe6m
CoxKDBHt5E7saM+r7L9mEMRxWLt5Ll3tvF7bGvRAD3fXmcuI5lHv+8PRCTTMjMzNktkuqGKkOwtA
cTIBAKVydkwDNiK9jeMrHf5N0kI3vNArARbMjK7OUgj54xK+feiz59HSV+PE2rKDfGE/LjECQWxE
fPrRTn0xjvADBur21Xxao7Y1gyggxcRfPOl+E3SWUoOzPZOEuQby/RPJfttgWqtT+bKczfqmuOeJ
zh3yL8XC9ybOxA4VoBsYK3ch+ZRrKkMqo4ONANyhapYIGtCbmWR22F9MXqOm3FtZ/7kOtkCyctsw
+9rVu5YNgkS+4FfiNZjnst2GIrN0tgGuogCH/zDzVV7wzCPQe+se83nBvIbYn+Uag3aS2tcSlwmF
zkjANTK4++wX0X53EJMHLpfdsPeI6RbhHGCYn548Jv9L1LaeBK51YzDotWYDpCgIsQ5pLGWrs5l/
xEcwRYUnHhKDmVHjurlGFpZpwGbFlMtKVBkPuITmqC7pAA6fg+Xyci3nmvIeJpVlFNDPk0QD6V/D
i2e4V5v6S92mBlOlUEnBnbr08mb1CujMeUCVXpTOhtWgujNEtJPUlITD8FXAxAo83O1eqdxkuvMN
HFKhAIOi1BcIIOe+Hb7ND4RndJ0udQ7SacMTr6+cZHX2LemxBlaS2bnuyQnCa7slf0zV4cmB6HN5
8IWyxUqvyjV3+ClTeGyRBNTlesflhG4s+dLZ1aUITj7PXqeIcLFBARNWZisx5q+pb93Rvq5PObV3
yjIYMqjJt3kmd06cM92LLxvETukF0SugbxufMAMk2r4teMqs0YCjFTcEGApBGdtqPhd1FcyRx0sx
pj/fCVOj+tiQA96PySIfOP6NcYA/rHRx116uBeISYHR6d25tJ0wOBFsrJ/iQ5WACXXeQAoA8o7h9
euA5lpsutAupenAZPhX/sVuIPKqVkBjKX9qh7SM8yH579CZG2QffAVEv2/ZXo4vZ1y1hG5x7S1Ca
dZHMtq46ugjDczrrJ2ld8A8MGELTxip9SDJH0vmJpPvGdKACj26UWh9hOaqrMMsWNAM3ACJQnpSa
5sgUXPAbMk3v3WHRfS9+8r+c6PvZz2/qVv3fxNsg7sH6Ms4skyXL6ZdEeM7/QJQZEzjeonWcrPqZ
kJ59s+hWJnWCgjRsf73hwAt3zgBo6VbAq+rfKFOS+hiMAPmVwS45uNQQZX9Tt4gU3h0D0IZ2beCD
NoSne6NjwWEaRF+BhJo2E1cuA6xa5JMQrjhXKX2W6E1/iAOqaQYL3Vj/XqUGlfRSeJj54rZTXRBm
oOAw3Pl/hDLqok7j5uqYHpvVK/eTmuTEDKjhYlyG8k9ajDgf34/nVHohcavHBMnac1guVtuLEDQn
gTAeAquOCF6fVNkltA2EFHPb26kvDJvEjxxLLpO+KU50zbMPSPY0AUsMQvdBjtfvi4ZtJ4Zf1cAe
BGmxsRyHq74veQUX6dOLE6W66r3Q/eWdUeqqM4Z0s9PR+bURCOP0ejZEElEzrHjgSKKMrgSLMKoJ
oYOQ1uw92zacoLtbGCYngg/WUt0xbLqgcGIWm4gZesXmd2jqR22ubMggQ/n7DsCHSG5FDwLfLVT5
hRGaYwWAyKjm4ZtpQBg4qlv8+Q/p23VTcOsa8Ts1p7qF2NpRq/LsA8zCKTn6ny7gwGhHH+sawWVd
jfgNYiyEu2H2k9fjFRjDmxFGK1eh/iFhzr5EjUj9bhhVSgHREEz2HAsFFMaxKgxbFi8/Fc4Y65Gm
Tic6tM9/u7sC0yDvhpxZ9NegNdzjX4fmiZG+oM9CYzVsAwRw71qs8RMqeI9qk8Wh239LZIlsfoHC
c/dRo9Xmr+5xgjK1J626OoPu+azWCHpTow0Ib8mGwQ4rMomaVydW2pkRoVpVcbCtWArln8qcfqf7
xd/R0W/9VlWJNoz7JtQaeA8loLg8KOYictJgZWy0Zad13Ebs5pnyquH8F7tVzgPxyJz16K8T4Hkq
5Be6DzbfwS9B4no0CeD1OM+Gg+4CdsjAYss76WHEeS26RInxPTFokInhASg2J11LNtaWIVmeh/Xa
W5qk42JdkuLbgAxCZX4+4NZ1hVXUk3yT8Vvk3OPCuYVRP6mKSpxJyUNZOkwWAL6nTbyFTKXvwCR1
5ObkB6IRPIv0y9hct5cXxUI1JSZCcjHKyM3Qpukr2InygpsFE3cWprIaYWrnSG496jeVDmTYJLpz
bU0sdZ/p7ALAeDrxJjs4XpfxRZDmhClB3njnXRV88Pq6LXwF2ezBEbChiYRm/jOWXbP+9zsU9sFt
PSZ+MGQkU8HOpABcv5PWjV36/6tFeQn9qzbCIjNFG489YvxNuhP9cp9ySDX9eI5GYz6RyVC0cUpQ
Bw0dwBGPnUEbuLfIq1gGQvecmXpg00Idi8fRjkLGjjaVcT3ab/IZ7MUd5plKtjyaje4/wxcSA428
tJuz0mhTDNYD+DceFzc5QlcfAo7wpL6+VKnoG1qObuUePFDOli/CEKzny18HqpCNsvK7SIWb8QrS
/yw7+SaEaVk9aLOb4WTJRlXVthavIq2YOHLtZIOg0NrxZ4vy/w8Y8VD39l+BXnVAu3a58QajxS7+
GzTOJWcO8af5CPiKWoYPp3eBcT613S97z5eMQ/BOKnwLPIS10RdpgFES3sZmM1iGd2l+23Pjz6Om
l/WS3PCaWWGK7mwqDFQr1QirXMsXxjLDxeY1mBT+yQeJ81BZY+0xtS1absD9cXUke4NoIfnVoryw
IW/1LwkgZuYEbQQRNB9rYJ+LDldGTSwzfT7JDrO9d/APSoDUr0Pc85mRtqbxV2R7Yg6r2VNGOLPb
41h5AI3NsI247zFid69xgWkfUyciwvrncJUZuZaytw+NH6Ikcn47Ni2xeixligTT6GfCOrJnnDB5
IoPdt4EsjzUcxV0nc+pfKmTv/DxXR3wntqdI98DngdKjA1e1NTGkRj1tVHcleVBAoxiQeHjGLZY9
JU0ZeZNNnIZmYIF8JGsZlntNuQpUQ4ILkTt8+7gJpHbtS/D6toFSHlpZhOcyJlDookNiHRkxTv5g
oztmLwiVGGzGkPtQMnhuDuNO+uD8jFXN9DYfWARaLQiofm8EtYzNF7I5l7EVnzIiGdPI70+lbm2i
tYVmK6G1jplTy0/KBjNh9HC5nIWaRqKQ87Y/YNrU4GR4VlTxo1/e5OxXO3w/EHRcGVOl3lY/chSJ
bvQicrEHXkxS7e3WHOgr0wmyrHAYYKy5b2VpsCH64WDOQQpvr7aLGAFJDKUocXK8t9upNqWvJLnU
GfYUpjltXvnKG1EAkLqbtouapmTGloWAZnNCnBQdYuNiZ5L+mJi/N88cvjzNXT25EiF0F7gt8z+8
/Gj3BW6t/fF1268wjs27ufiG5v06w21LzDrk3UA+iCxuY/9sQaHT4C1lonX6NOdAx8bnhUpua58e
59gPUS2sP2pALx5d1FNL6nZ3tFL+ut60db/EFVuqdGf/jejSO/A/CGfvevde2B/+SAecYsjRN0Lb
C+jnqJ7GXPLZyCuJghU1VR1Q1xy+WXRjvgyWCr7Wlaqs2pkbPxqNkS7Kp/RpgbanvcCi8BcphNbl
bH35yL1MXHKXgSemMSqW+xX1EHJRVUyX2yYYI0Fn3t3ABm4b8CxmXLMwQNdEUnoVLvFdgpyZHrJe
8alUWRoE6xq6xO0eG7XAw6Ia89BHfxI2lGjAzuDI6I1OtPe/9jSOHDoB6xaSKV0f4r/L2uAb+3wh
rgS8Lp48ZtEAlHi12WzxiK7BlgxOUKfavBrWE/kxYHPMjyhkrFshJZICs4b9FSogLCzNqZ3dqtGd
y2Ah6Na8Hk+hh7rH1pNCtt0dsawFyo+fztXEJnDVEe6yZ4N/80LllYeKazjU80S54Be8KmVtxF+v
8dsxYVkeFlAekEGqU//N2Vn7Z52ZqPx+LRPUn+Mre9ligCtRxMJu3z88JDLq8WUcpbdz+1YpBssm
5+r+N49EAVSc3HaU0bSLGPrXBtktfrNhHd+vL4DVGyt73+GuCKtuT5fqOEoh5E39Y2aMvxstGuCh
pPYvPb70ZnNCwZgUcXweERH3Fkwuyb73XLMY0URRIuVVToXqDlRz3M3iHWUr3vfuT1IRooW+dzvB
8I43i+sWyv9ENpGG4diM7SDDXZ6oV+Ub9A3Qo4ueofPZ1u6S1jRY+TSj5Ri6fAuQvTyvrfoJUYZq
1bxbJprwE0WV6ZvdAR+zXCb9iF6zJmfROc+lxRq0cKDgf21uAa6whFK8biz23OdpYDV2eyuO1l86
TqNTErGBoqNa9b1ypS0TRA6Rp3i0e6aRieJmTsYaBBzCYYhHbQBFse3G1IGvXfUBA0WswHjZJSMp
6vu1l4ae0mGH9CXBsYK7/Ds2jvhYJuRaQN+B7Pz/v2DIDOpSMapUX/QN3jS+DijOdA6/CwBPrsVO
3QKfRRqaKxWtcCkwYB1LACT0uKqhH/xtRWY5ApYRq2jWpxY09XWd7HFbOir253BHx2t3x/O+cd10
ClfCFIKcjQw2rvuuWkU9nJdjlLrXJkUui3jf3bNDQ1T6v8mVk+YsOUAG60BodveSqjxiHJ8qKjx6
8ZMrZRaaTRGZ0tBmro8G30N944Hzpzx/zG0TMBsin9sZK7KZcjm9k/SbryOzZm8sT0XgpnRqtHFI
3GdvvIcH6t0IKAjD/UmGCAIosYycE+GR07sID/LsaMLpB7rVibB7WffO0aohd6OQDiYeBRLXcNwH
6fNYOt+XYfKEAC2wU4KenDykLrujjb8qQg6VVhCzRkrSk7PwZTwQt/irq4WfrvJH+lA3KXLP0yK1
WCoN6xbQqYtSpnstPf8BLPW9qZ70cBRtsRAgk41BiBPFv2Q/i8luH9WHALI7dYiLksSv2nPn76kV
2m7IqKza8Wm+rTI3+BYZ9iyKCZsKSe6ILD6HC5c1cOS6fJscpft7wI3jKoAnktAk/OJ9kXZTUvPe
lC7QovVIV1aK1rBthSmKMAO37/5XFa565wQjWadvfOUZZlVhArQVkKudepRWaB/Xq7NQ3GmEtQWn
BKd1976MqtDG4NX+fklj/tFm9D5+eUvbof6Sv1uQEdzlBcyS4k0OxtycTWZ4MAMiwbZ+r64w6TRo
IWIL3uM2LZQlHrNRg2+d8d3D2Gox/jLlj8NJdx9Ym9ENYAlGseHYdGHsuWg5Tq4181q0+DPKd3DU
T3ybuEWaPo5PGKt7/IJap47Xv7g4JY92gX667RtPGTR220a9huH9pjmMWwU4Iewzdkv5qDOV/hu8
75pT7iDlYxsw2p1hRvWBtyw/0mJIn0NQ9Fs6zY1ilWFxz11TROAtoAQk3aYqY4MRlJknAiEHaKYC
ScAaK238/oA97Vtf+rYDBON88ozLCIwT36zb4PJjDcRNpvaFwBgyMP+LC9TLVXqMzpVjX08+XIy/
pkfJW71fJI8dMx+OiT5L9BmofDgRlxq2gvTWZ4T5dYU1r7jImhg0NtRTNYkbPiEKNWsLtXkfpihe
MVnD7xSuNTClrFVSNZ/TNhZmKOXu9fvBA9ZCf0lDp5NvMKy3NKAa5SeG4+/qO7oQMoDMqaqHeP8z
8MhJkmLRidx5GJMwdDTME4XdUajIrN9TKH8gDbALyU/FSEFsoMXreQcRofQiJhtk4/5Ryde2UEoH
iH58nu2WDkfEKxP7DMv/PFtT4zF6MyLbkQ8Cn7KwFbnKrvxwP2O8WwLLDDU8G7LVtoRK+CURs95c
DHt7M5jD17idqXMTuJoxglasfEFQZ6QSxBz9k06Prv4pRAfZN/rp0ATbofr3rYKpSz3W2BzkMffQ
AD9kExp7pOEDAzrodVRf4iu6nQQA7+nqSeTDJEzJ1YFE6F4SWanZA9vh5MMc4joJ6WErxucsijyf
EQ1MBRtZvpoUoBP4PFDf3QOxTOoYeiyexoCpatPnZHZCmkbfvXOElO2uRwKKrQvi5WfrE8eIVgfP
iics6PKxlj1ZjL11uq4wBOrpHllVn/3hAV6dxYuJ1b4noB6sw5MtBZL0ejew189Zmd1Ru1EIq/6q
h9WbgvnnoNZadnpn/m8vqid9URjn6mPXIiiO/UgkuPSTpz7R+sRDkAO92wlDD/M8noDIL4PnV21P
3yvo2uPMnF8D72iFz7ZtMr13vcEYKfAf5DF9BedsCeomrhx6GxjdlNbtUOsqcPiQKl9Bn1iJ1VKt
AJQbQpQ9zLXLPCVXxvHM0B/L4X6CzM+kalvEtiwiDSjULR21mVWInVdeeTHBeD4T73WEUfFZ6+0N
VRqP5IyCxU24s55NEAwH8jHEjusQL1cWkvJVRYe+ACOBUSERxlEuDicRWKSEHyfFCFs2I+Qh5mIB
y9SzcZOrwIfR0C7iPCTZeIjKMhrA2QwvEm7ryD2+ioo94tIq5eccCRQQdJLeOXhi2dx51T5IYJZW
XM6tW7ySWwQ0cUDJa6j4QR2ETsbVur9x6yxtQaH3QEetJFyD0UrRVBi6xheHHnkVKy3ZSzZuXyst
FpfxE2naUvx0Qrzuz2kaiK4hYqv4maijlrhmsEZjNGwAhVMS84atDfY+FXMS2EH2w/iOsyOmoz45
I+OBAu04QX6IgI5GmmJ3g6D0BtQBj4Y9Puex+2rCbI0LDUW6rW1W0TBU2NvWmRnEzvZpDm3dKawe
rlARHzG/156BOAtV/1ceZk2dNn8sFokeCi1ZSD7XJfRgGI9Av6Ax7P3OKCWU4Gfuo6oQNjul3GGS
sAbPkM+NWI5mk8GIjM1/kpRrKvWHpo8ucIaIPd365rt4qIUrKFDiMTCvcsNTUB41AlYwlMZ/j/DZ
M71JZrpNTYLcKIA/LuS83VgGqfAlXl4tqDDr+7uuO1bSJiCcf5zB+p1Mh0SMEWsRtW9kVpoLpT6c
hmrS/++HY3iDhXUwJ/24eDaFEEisYd9FrVnpXQr0XK8LQrzDbwxYzdQESPzYdpXNMyFV3aehxqiw
3eERqLOM8nDVLA4Sbjed/OTntVRCw6wl/k8hKIyopH+KNoR3l1MD81eShU/RXTBtdPHBCqaMfyCx
3qsriMC2tbMj5QmJPUnoiub72xwPC5Z1rZ/nNyLPO+kxwzQKIaJh1bino1Y7tom7fCMIB8+zUrOJ
hLZnCsuGTI9hknRufG5BTtXB5IY+4+9M+kGNQe+SSKNanD39nT4aj23dUitKmIvY+wb0Tudakmo8
SrVQKVl2nMBNUnVkpXe/TYDtDRlg6Wfll30fDIcpqwGdok9jQmatwE3LCrUMRkWUyik1JAbF35sj
IZwrN2209D07zEPZ3WlTf4q26T1Q0tWMcWdN/ziRC30zXYrLwvEthYKslhlOEpWQTKkOseFYP5rv
cDi2OoBBc2rQwNBbWos8rnojzQLpmIiOn+Kxt1BWmJmj6A/dwCZO0cAQ8FGa3wZ4PsdMaX/WBbIW
DGuXc7QDNIKu3mhDGpR+4RB4XnrJScknhbbEv91yB5KX41QKQUy4ekM8RLuMDNvquuF/AIJN7m4i
WWptKk1Gn7g7DVhSqG3bxDvm2Znw83g+qwK3mfxG5wsYNk98RkSXqcnvTeiJb+ojTisoQvR7Dv+h
ovQeXAWra5k8ICQNMN1IRDIw/pQlmuOjJ/+t1FpR2Pn5mMPlN8+MSw5TO8R1NueVYvP964IPkPaq
+jmNDUXbqurdKCDp4Xu47+iF0WcszoYnvbMsJIvOrEM/eHIQggOPp0EupaHNXxhyYoYJ7jE41ThN
LFzYPGouTIty4Z3AvuclcW5FRuBtXED321DWzSvwWuaO4tbVGhpTbB51HeTDg9e68S/ZNKrL5YXP
N1qp9WDghjTQhDXTISCZ3rF4OqG5kmtoegVf1rNLHu8z7n/1DeZYwuq44lEcykjrtXY65TJty09n
Skpwn/IZLjTUF003VJttNQETcZTn5WChiAPMzZXRDvWPcNrj+0EvLL50QhJ/fRHVNShrDCBTWWM1
NtgiOPbPb8fCk/TvrwjzYwNNEDOOBZxKTFSDwB7fx7HiDxEGCHbJzZyg7P2b+20j4MbP3Eww8uQD
I/hIPNkPOlvdckmF30J8p1Y6Oys1lpWFmmPFClO3OEM/nNs7ZKb2ReJV9qSc/4MNPChqqaCePiY4
rVU8K4WFd13E/sxe3NK4qPzkl1JudiSlBgmj2RG4kvasXrMBOB7di00z4zEPfN8CRBqaG1PA8F2g
I7rfTbJRRUegrtLwLDPAXMVnx2aflR/JSyXGNl1l/bdLVJbLDAQiuxkkZrsdxVrfT27ccqf9P32b
CRwTSmKLepD+AOo67G3RKnxq9mBxH4wXnQV14MKrlNJUNyN0w+fkoEEH1JlVB0bKFGPEo0mmG6sW
MlZgDZZVma4nIh0ytpatZuG031ah67zscK3MQk/j9m8E303WxyXezdQ99wvGJIS9bJKQkygrQ/X5
enOzbJIriU1RDD6a34z40Gv39IJGJ995xV0xVxwLKmaRpHYkVcZxPap4bvFMKXLrDjjJyIfvFEcS
06CcUSNpDeVdW/B4Hi+dQgCjOWnLuMh0879QIsGy+NmInLIufHSNTVYcuMJB4AZpT1yOcUlIGM0V
Fn1dqPrHEZeFebLXLe+fbHL8ByBrnUltM9KpKdyM5X7UmHIqahzEpst0+QToXxcQ9yn2PBB00C0+
/eboDyGS7ACLMedM9J3i0TN17rbXdBOHeKQ6QG0/Z0mUMiWRSfwpQs8UjBJS24KMCkAFFsa5YmIj
QqJq0vnyPpp+MF12z5aqv+BFFiHey929+0wIJ2Yc7n/hXzNcg8IA2dUV8cRMDeVaZVnid1oDy+1l
SiOQpOAM0rDaoxVV0XgaXal4lpZ6ynfB9JFO6Bye5iFFS9BwArAor55KT/JbS1/cEy9tRacntOue
gjTQrnnk1l8E2Dr80Pl4Plsd7+VNrwIGAGthWLfmbDQINDWcupj1jx+uCy3tyWZPYwWo6h7jbxeA
jIgCqKS6w/GtIWSlIjNaHsnFaQD+ZqgdK/2SnkUo/dsXN9q44jz7wF5LHNGcyNEv1ozVeLE2bKFx
M+5wVzPJJfyuU+5tss1+7JLGWluL2qGbZtf++ykHqlkyZdbCsWdVB8eUNYF9vN/ajXU5Fi1A5Uyb
hzzoIf+glWrESfYtYWBfbuY4rJmCExc2Ee+5swZxds0fDRpUGFlqHVWIM2KAiyxVupjRLofSFKV+
5fCJaObXlsLt6ODkYefDQFWSwefMshlN5SGmm/UTAL3R/VwCcLskfmUzEsLqXpOl+bya5zy0TW8C
bsvDC5G9UWDjrnsjDte/TRLgA1J7deYjlnpXoJtEqXwx+XYY9oWAFm2mQTmFLIhm4u4D4vnIkbRc
r0a58DXf4Tlggu1V69uE7IW8PwLI40Ck7WiaN7B/jKfQ47sNwITMvrjOdKant20NjKIvhBvgMJAX
6QOSsVTQBylNmAws0V4fREuS4Aa4aomzjS6AEx50L6UO5VW50fF+c9NpCxP6zwu9B5qaJp//XeBU
tlVWr7MDa9iVhYQKM8qr+wC+LfjifSJ0nh4GSJaDRJitdXRg3/birJQHLnQQCXsIgpyf8pyWEDKJ
ccTQpset9rN5gXABSaQ0KHoNLPdqoHl77FYz17QFPUpNjT9zxacVlDUdC86A9z8ZS6Aj7EA5xpYp
5WyUJ8BB/sUZ8NFbuydhalkHDZDnzMJSooZGBvi35tCx8csi63qQN+QW2oYK826r7eiK0EvTitLv
czWJO6U/5FExUfXI06n0ByOXqtFKd/sUZDph9ghdOqinqMCHYnCmBJqifhClnWdEeQJC/BWE6jWD
6ytKkgrR/x4r9cOoE3vujGIxmDRCDhuqSOsVZSp/4RMyjyqeJLrarH8QDT7lzKo/bS+jV+gOFqW7
Do2zU2Q9tWYQkT4agJ5grBOj8ieOgkAtrx5wl4AY2JXKpRaPmOJvOjoYjZBz7kKy6QZ8frqRWsy9
3dhrSVO5UXRIxBoLgFmsu8O7tygsg/0MjBZs+aFdaREITd0wtXRqbL//VaXwGp7Wjc+g7VJ8wPEy
s9Q3N9qdPONaO8RQMMaLHC5XeV9UyIqU2M8i9gcpse1AV2BVo7eS4zR7rtSUQzQAEKmUzHWwWpQS
cnMiPB5hGzV97rrJy5iuCCqWn62Dw0ctspaAeHDP7DHGa8C6XSB1JpJ3cnf2+SX7/LEds6L8pdaZ
PBFcuOnr9lrJSOpEozY+5PfsHS9FcpjjAk8s2u4lxmVVqVgTKmgGRpAENmFIFE5xofOL/CYhP6IZ
wT0ia2Ra0PUa/YQjUmj5GTipZ45IhVbKQAo+4XY3ycoysFJV0ajZUMH8P/bFGZq9ziZPhCpMDOy4
o49+5hQgVADeSvqW9v62ZSaEW1fjNM2w108iTyLneSvJhs1QmYf1FfyvXLY61aneX0zbmvPW89/v
5xJAq0zbWqYeCiEUTNjkacomze35fWligFyFyN7zHFnWH1cLo3ggputSXIJVzdGdMWKj/1Qbgogc
aq9YhQYytoCDHaDdyIUT6PEdwxaUufT2jM+4oe22m5QUJI59HV9lnNH8oJS/PCSNyFNeUl7hal8J
AsOZscsZCWeguxldsry0ZJ7hDAXKK5Bs1BH52ODuVb8EBATK0NSOGBU9AIOWl6cTevWbYVEXyE/R
bISyXSDCovmvWjl1wJR8ykA4jasaAQ6hZqfrUAoH0Qkh/sy3MbkGYG6ggdpqG8THJn0hgvtD7JyW
QvYBrRSUQhb4q06UaKVBbRxqizSeHMQBrcVgLp0wz4HoQvDzUGp7T5SXSJenbEiApdmaXZ4gWx9m
AYXzz+hp8m/y81z8L4jPoJAraouGMT6wWdJPyX1rUPn77IX0UnQ911I7reEzC/C/QpL9i4OUzRq/
SGLNs/N/JkU13nKhoBMkE1y5fagfe5jP0ICu4zdHv0MPHRSTzfnsp3+UcdDagzymUQsjlQ9eDGmE
HA+FXwthdUq4GpzPc2nNDf36aHWTTxspE/Sej5hYJY/pk7zlZQDJJVuRh2bWzNg2EUeoMNczCR9G
fPBalvVzhlX7z0tDyytoqUiAc8Fko9zoZjQQiXofhDL3FbcGaGt7zvMjsGzCtqzJse21+QRHAqTY
vv1IkFG0wm6djKeC4mv9mjuyy+a04CG/5ybu2r23OqGUpCzjPD9n4nJSg3M49rJg4IXPVF1qF2wN
fkLrXB/xbzdZPxVfD66HiZ480IFoXGYefA2+/lgolwK/Ndptm2R9lwnD0BYMrWvb0Ebr8TxcGzeP
9+ug1idajzmTuDas3MmLoM11YJ/RkA6kKXJw4uzsIWdBkpOpKL0GmZ3mqzR6qN3RLCrmtITU2T4Z
M28KW1FC8+ogzn8DP/doJFqPBYRPHpFB20X/rCAyQc3yYFvaqjZPWeiRjs4n1ELiwwL0EVkEVtzS
2DjXQ1NB8I6H/F5in9MTV3dYGJN1P+LrtAMDZX/4DccjckbiftlAtoJpsp92Ul2HuE3REHEC7dhW
DybLybW7Hfn0P/LOEsIvBp2/BYbHq3O41AC2irba6pxPLYAHLk7LhIukvZN7iQVhuRv9qnN2C0Mf
4oyvrczdgL/ENgIIL1L4Mby4xfFsV/+HdtiCbEwHHsZztrLWEuvBpCqiHe8y1EYEKYjtypG+Faaz
s/BcMEfmqR6tDd6bEhwdGH6uFzx8zboY+cSHaYEhJKiXSGqfRqImwLJMbeWHwoaz6wc7/g8Uz3di
V4qXDtub6peKxb005ZK8H30l878A9unLlABSjxapGe6pUcoqEqa7NOXbXODCmkPhIbf5ehPhzkzT
N3MJDbL61E68gnI3RZt+Gvm5EfR08Yioibzb6ssu9HvQDLjXZJbbhLyK4WqFpUaBnPzKv8GcnoA6
zQyLwIT9F2SBNz8hQLZ6oWQoAR9Gpz2P2mj7qhrnjbaFkDxSuBomuvobv+bkos1wXpKzn/gQTt52
GhhIgXancHQKaymdkeAORf5LlnrC/Rbaiqs3Zp5LlftLptIV1aqpMQdwx2FeyNt/KGga9/E2skGN
kUXp9RGoQEu8FFcG0zsDR2J2qyxp42Dm0ZR1Jadr//xZlV9soYLqTwE1f+KPLWyJHnxsKzs3WNXy
/3Pz1CMnWY1+VpcfIol0nhlfaF07QByAuRTgRLMEFATlLpcsvqXJd9ckK37DMas2DdLiA0emwz4s
c5zppH/dh/NQmLgzRrzzCKs1HK2fHZB7WcMWd3ylcJRKDjQvQ9n2B4KJoU0OqX91ifa4xq9S7y9L
FGwtGW1E5IKzEj6h/rIV1AQQfTQBxMX4upF1DNwYWJSSBcZLgECwLEnX6/T1Ib5/LWhw3fPoWyvt
LFw+gu6YCFVBdvB5nIjSlR3HX4YhVDhmNXRRDqjXnK1eCXqMeYunZg53GlykuamIxoBcVbuSy/g2
MEbSc882jgJaHjnWhAqoLEbfN5qQF8qcTZbftlJj+Sp14zdnstH3zSrFmxUqi3bzO17a3LbMjplG
0cUIt0DQyok+TwNw1f7kASCa5ccsKZ9a9DcNoNqNkU5F+AseQV29K9s+rhTJ64xz32xriDJxm72r
Zwl7t0v4nkcvlAGurwyCoVDewJm6rH6lqAtdNZ50PLhf9VlKp/rVrKfYAI8GLhgalmgcTxRXq381
qLmYloyYT0rVzqDDH+g/RjUX1mfCC7L8yymO90Cv2YmUC+jjGpJK3m4S1W0vInxXm2TUJzULZJGn
Ndg6S+wkfDY00Q/3iboOvkBqumrYBDLl53qZ/dOwvry7l/JsTK0ppeIo6gZp4jdFRqVICDcA+fcD
ZNrEHJNdjbczmLmrJCtix/3XDRYpx3y79YorBNGVll0SEGsgdFxbjpJmuQ0CAV6dPVJc09UJ37HM
2Ik2fMQgbdlAYRD7E5jPhC4qus6/tIV0EFli85iFsyRQVVULioWjirSt67AT8WL0KHUe9anl7Jbi
tcLXda3zfMNfykXVkGk9qTFmx3GVObilyI1BTzi++hpocHDwy2Gd7c0AEQqbibU0bJThgjgB/GlW
D0NduypcjHkxIUElakIjj754We/UvzYXv8ESg2cHVucX7AgRO/K0HV0Sb67K1miOBUOXYU+r6JyZ
Zh5KA4zPO4s5HpWoX3XT0TdfYnKVyarmBMkc62ZZrqm2ArtCSBj7vJvw5AxPk9NJ442G+qoDtvRc
44ku7UynBNekZkh60aG7jGUwCCHF12WmALgXNMaIUeQWm3+jzb7BWBUm0ZJzaOvmMNKtfXePK0yp
ce1Gotgr+kUJJk4opv+P3qGBYyeLpY/0mq3x8E/7uIvWBqhFUBoI4VQ2+DmD7xC+yybLRTcNN2uR
7asFISxuuy6Uf0T6cY7rpRKDaJ8ooM+WP/22F7O9Lf/VlYBDyOuIds/VxMOQoR39BkWa6KtBEnHH
FdPPSdTa4/M68JzdKHhkZT+f7i8Lo19hZQ3uaTxBo1kMJFVXbS7UjrHerd3qQRgy2/Ewoi2DD5P7
KS5LjOps2uWMLscyhfrAdFMwmWnprvziM2NUl8vDmP/Y3s6OeHosf/r0kVPMzzsX1W3E1iKii7sq
5sI5Kj2rjhhOvg8tA+nDtIsIP0ysETqnz5GXI0iuBeoBSMTGrfLmaivOQmdYgS5OVpOL0QD7eyj7
wgUj+7DYs0HUoFeRfSpS86pEH20B8pXthvoFvI2pdvfHyezk5p0vOu2vG/TWPXG3cOoJoq3Gx8/5
3YgAB3ziMGgtZyaNwcqHxXBBhih9Xk/MiPZMGBYcR3HHr8TGrcZg+64+uyyjyZ0bKcDIQBqm884V
AGQi36Xfn7zJUODkgd8HxOr0eikq2hG8zqqfu3L3yhRIBxy/VjpcQMJNXnsgyaIgNzVXSuQzV1Ad
8TBZ89tOiUmEKXytirOT89qs56/sQv+/n9fmqKzaLnXy2m2qWUqRJcyI/Mj7AXpVnkbS/NJupsCw
70rZMQNtkVIQ/++t5mdiWD5P6+ih0RUpMwnFN675x85FXmfw2EgENbrA/icrJYY1JI5E6GOv5pPd
V5GfCkPs+KMh/uLHFob9WTOSePiNcftGNG2tRlWfFCM/x39h2s+q68tJbH1cGLwxR6Uid0pfQ/lK
oq3slBit3Vp3neCBKo4YjaIv49zDHlq6Q3Vkf3k8w3TkKs82fgymy92TgtoJn0zr5+1SFGM3mVFd
nrGK1AtpH0t4ZaCbkc5/NQFOquMphKqQ34oxCq1GuHZHuyX4UfWHyGkdUb5WDfyEwl7vWyh6IlgW
hhOvL6jIO1OrLo0k2SpouSbkFKbKJU/VKsLs3a9o2X1L8e8jpzw/PtVmu+sG4WaK4nFq/1NM7SrA
MUAONJfiSLoZM7oQFLtYbcdDd1eqqyChGlRk51TUEvoZX65IzWWzE54kciDlR7SUDtQ3Y+Gm3gWr
W+bsSVFtN2/+3hNFNXdA9atxIGEIfXIP6OnQY82Z883QjKyuQ6IZn/Zh29PRy7oETVmmN7tCTt9J
xOpzfiPa3UZt+LekTLEWTu1nw6fBgyncWPOiDKUkdL3WLVdeYinE7DCj6T3J5z6qdiqe1nZSPYK4
gvxfE3RuieNjr0By9+NJGy9Y38QCqnwGOAujYrHIfxoamsGqZw4EYlO923JL4WjjR++l3pBBGs4c
vDFTWBF4rfycvPXKxUacX9/5MLlOdagfdyOZknLQHqIegyiomxb+vtGfBX6gUcn1z3yZ1hIxVW2a
XnIYUQPeTyMXR8yqGO9tNDrrofDPF/3jik2bYVRpnGuuGrKS7292Adhk9zQooLZr4A6jB070DFst
d+0ZqzQ8TipbtLq1whFrH4HMiEgcz0AEv6Vq59mTSlscGz7bhuHOf7iCuP7h9QMdS7uKTqQJ2XAF
+HuFLMe3q/i121DGTB7IQ/+4IdmAkRMv1il4vBf3uW/3e+YWdMUGNiUXq3R77ZsVG0ws3hKh+U2H
saQBmjG+UU4CWk5vrIVrJskT0g5r/XH351HKxWcZ5nNjkKZub0CLURw/Fi4bjzyG+zlCc4P6Orp6
cZmSuJABRpcGdF38n69nQ15X8ixjw2V1ucI2rhpsxzs1v+uoPH6f3p/Im4uSbbA04ZE9WF/H284p
Rpq3a9esVz6cJKRAE4uJbHtNLDpctUjlhnxlQYHyJAWldnDjQkJ+r2aVqJ3jkrxjzssHaJ2tSlqs
XVMc9fvGE/5+5NAbO04gslnrfAHihgsgZMFTidoKU3OFxBR6Cs1gn+XjIKpD0MDD9iuQM9CHQ+sQ
4RX5xIcxoRqEQy3Tnr7bbUwXCvhCx2i84LzhzvaUvAQqW76mytxoLZsmQhevVBXuRYVKZYhmUK9p
76Ox+MLTOIOROKdGyxrRfg0ycyBWmsbt1ymvgbuUxM76BMNaMql4Sjq/exXoyADUeA2y90iM0+ED
i5anMXvigw5OIHFTfOToxg4en1qcMh6fLFQyq9fvHVyLucIO+IfVWzAobAaXgwYhiJLPq/Eql6MQ
Gv5/ssv7A/CfA6cKzv+5apxGTMeSsRDnGdkZN0FfzKNdYAXZ6HbW3n8cKRiXonO6d3msKiJiztS+
O7qbN3S6We8PaU4HSaPLkB0XEu7U9MqFjAbejygGMNMFpI1tASqiyygjM5ZvQ/3m0Q1pqc7X5+lT
55cBAKOTiXFIWX0fK4UStiq6DuqR8IFB1zjzNelxk+6Ey9CCA+lamfyTDh9J+Eg47kbw88g6k/Ur
SOA59BqrvLA3yQdo55WH97UlVv/wXQVt2LlHtpbafYoerDrW4zd+HDwc+yvSAlp2LLFG8fgYD/pL
i1Bfpy6M6o7HgYiEetGz6LmEXjx8nEjPPZUiDiGMueVeFBJvQVORnCWOU6pG2C+KQ3nCIwGQDf5L
91uGnWs0opBwvvKJn2jSMbXz2iEHyKnc2/F4Wm5yjBAZ059s7I8z76ZGBise3HDxg8msdkka474u
x/uSkPvPChNRlMAh6NVr/OZAeD5x6yWT3TUUdVdzZdfvcZ0PmIqJws7x+r9R3OLNGWHdZaOAerIv
/6+w7BlkSjvkcsRzc7Ly6MV2rkKtEXN1jCEj1+Y5oy5fjpe+ccoGgtjlnWOWM5v9ktqhZtafxXRB
kgj1RuMXcpd2SX3iFzSi+Flw5imW/7z3GjArZSLK0QdntQ2PzW/BP5xvsMcC2bgzeHFmfGx9if/6
zAn44GUjmejWQDLwmtXRUpVw6jUrA291Cn9p1ZGWVxlXhnT0XdMe8N4s0trgAi2FgFwjCRkRfyMm
Zpznd0d0mU0ZaXgHiR8RfvpDJ9q/dCs9/WeoybMwl5Pnp9br7hoYqSJ1eTpC/Lrpef0cFOlPvsw1
LEjzFMnH7d+MgNK2+edy3orkoozvtwBnSYB+hUrBJGYZiGeA+adArBjhuZPvmyk+Twpz/Kw30OpD
sDmK2NRf0pbHvNwOPR46sFBbobe7wDjGfT0rZH+31Sp8DxehxuWhlAOmuBhVF2M8b+O62uh37KJz
kZEfXx1a1s439wxvj9o2j3zSEt7UmYvVFcH+exDDFD8GeGATzGzcvEVJg9hJIQs5WC1my40BpqjN
Qd+m0DNU+w++fNfWZDcXZmKUDytQOJlFCYP2je4V1ktV1h6Afgyqu3sXCBb2gm9J6n4uiA3KYfTa
EpnU4rZMR3RwUgnsy0bhuhhDbISI0xRRetPC/HIv2ZNEDsTpWQnwEQ3MQjOn+A0j1cHDXgaNACCt
zCSrRKJbqfKKR99DbCwT73VyEyGFB2B/mQkxDTVY8iDqn2dPKY7iJvQVJci11K5ZSxF8cVcIkK3W
R9IObsAvOeAZ27TcV/NlhxX9p91XXE94L+saImjM3j7XPrCzvCXJ4earBORV2n/GpcZ4BWRiBCrL
fCL1SoWRf7Y0jQMrHu90208lDK5Me4zd2+KbqPGmGBkJnTwlajpmr7E+O2qU9LJ+rpi65xDNGfd4
RfoTbj/DnYmGylcrS/xNvUS0XBLdhG/Wsb8krw+li+imdyILFr+JVF+qnbBdVPXjf8C88uCNMtUL
TfQKopsvOauNEV336Z5hnXQgDz7+eGUPOgnNobn1QBSUSAK3IPAp5regFIIx9GgtbZAXdpJMq4E2
Inpn8TtrBdtcgvyOKryvnsPyyxNHbVvfhgA0n9kAHA6+7V+qS4dU+HzDZgWTFRlepO+Z9Hxl67JB
jJt4cVap6Og68+z5P8TR/O45yvhFGsc0ReiqQBe3+jUKV3w3x8W5Gs7Hqyn0MYV6Oo5LP1OBrlmG
LDjcAQkHA+otXz2skEkUs5+vnzMpOlPrE43inofC7dJiPkqGpk+uT/ZjbVX427VFKhcftILIKhRC
YffBJv0vlZgHAbJ5AuMAfiBAnImzNbIm/6yrBEKXFlA0aj+KpouSHJ/pwEusOqMV+RZgK6p9sh1M
2Ak7KTLnpNcKAF4NNAXn6MgHDh2zAr5VBWs8T2khtIIN0GcaMz0Khrsvvs/k+z9DZli2f2KT67tS
lmhF+3c+gBoU/uSCqMummCaNWJkcG5HFojl/sR38A3bKQd7soKnjbpfwCQd+u5vvYH5p4VWkdUDr
JxdcHZKNZuUetmByN4lCaEqXjOAyp4l0Crv2V7McW4Woy8b7XbL4KLuouKcsBKQ1B+8y/xLkeeCn
NgtCoy3KbSaY2HsrJtuCxVN3KJH6SEHxFCTwLdu/6dKI7fplrTJx8ZbVeFuXiFqTIMJI5WGycfgF
QaUBaR+FHl9i9q3SMkNFNU+O6JSHJp8gB7Uqxs05XuVdQEqguo/CDIVFZDABmhCRSe34RUldzQ5n
ypnN0p0uvFULprHDuItXZwoPcFfcFLLuoOEbU+QFrPCoKFt/UdUJG+gOw2KjPFo+mP1hObDibxU6
9sLnzrI1XkMHLkrrSNz+r/+1XWdl+wZxpYN9zWJOtJuveXlUdxgCwQIi/sOkO3ywhfGgLQ29xeeR
54gL4sXXqnlYsHkgo/PVsB95TwJE76HWDglMQEg6PIfjNXm7CPnwGKVpxBzZYmpH6B6+YdSCl5Tj
GU4ACdQDX94HOSojiJg9iGr29xE4ij/ZuynDtm37R4VECJmHO9B2UxUjJjlzLjD4hk25JquTiAZW
H0nf4o9Fej7WAYJsYr/z9Ob4/DlYQpQp2ebP8wDzFe/B5CczS4VZ5Be6FU5dHn/ZuKQ8WL+jyW/8
dIWP7PwEgNZ6HcsJ8qUbqg+eZlV6VqUcrCgGy+jftNt59EizPInmmQ2fCy0YJERTP+5oqb+0HMPl
mL+Nkq6s2rkKOnvyi/K76BAZC6SbX1ntuX1WnrbxDpdribzHtLo2rmTYXcBHDav8k83b6uHZpaoB
IF7C4dY8ywTBFHC3BHEo+vAZ68ZmxFIgfkjP2dO9Octdr9zFyQJ3Ck7bHJZBOw6xwg6zH1QWMxaA
I4SWju5W47q92OIn+WwZtXNaJZbRaCrlEug6MGVl0eh7vu56PDplN7wxOjNs9CSEsfHgaLWm94Se
k7X2xKqnMrNLzontESavF0ENY9VNY+4ee0mc4w5S9lzw4KGA9uaHoGQ1iwcwpVs+6GlHMmOtSi4n
86Tdajy7ynTjT86ybBEKtDFEpOAXkW+itGOIbVwmZtMXE2tIHqGJplW0N9IMej0j4WWB2QmaN3Oe
78YpldxVGrpDClZFkDvC8OL5prNWurRglRk5ezO7TxQ1NCCieVkkSU3tpkYVjZO8Jbmvjh2oOBYl
z4NtbhotxrUE1MyKM9kvQ4g6MiKRHo4enUQV9awY9swbiEjpva2qHhj2VCM+tlXvL23a44ssZntp
BSa9jVYs76vcLBshEfMPXsaPDE6Ks1du8osk5kSf7H4SblzYbrRLN+1rr/bzNnT6vRZkmhIVPfGa
mCLffoglX0O0s+XTizbQEQ/qBiiPlTKzmY1bdkUcfIetUF5ASjBmTbzFfkqqjjFJUTS8zUA5hpE9
PBxS7ZIGn94G6M95RdxTN4D2KfFBmfktOT9fOF9aG5iQUgSB+fUElqmlGTACbR2t4jcUif/SBa8u
L5lViRzHJM6a57gniyPDIhWbqqi9PkDkQDOBAgv5GMGdEUETMGasf8OCrGOHfEffkJICO4Tu+vm+
cPV7g06RF5QgSpteyDy9k79jYj+0kJq3hotptcUrx9v43WpxYwEE8MXBg+qV05hIy+VOXKsAcGXs
00epsn8Lk0OGBWCfM+QEUqotIjH8wmSnorFKbznhQYdzyqGbirlQ/Hs15PK6+R0AKZRp++r9q4Cf
6GdMG4ziPYyfDbfvdmJxuNj/LhfIA5p2Bs18cFNxf8XyWloa6LDqmJECmAHmmgq9GD/oH2Dmt9lG
X4A2YD6odRDzlNjI+qiUcl554TiszFCRX/nf7nwYySiLOLHS7ynyowaY8pw0rQ4nq5KvgpwPuceZ
6IqHxIxw65GpPO9eAMSgdnwoWnFR1Lmfme04h7iDN3MY3Gr13H3P7j5LRwPzUO730+lgbJ8gXQ2n
053ZL60EiZ/KbVTQj/2yJ7xxbUlDamZBPuEeFY0x2zC88fJI1g2W2b/L63+B3V6cW/B0Y6PKbfaJ
6nHlyvXtjXfidMd4HWOJLbYI9XFPkBy2tINbB3sKnm8ky923yK/uZ+akRImlLySD5cTB8t+Irbbs
zRtQceawrnKWqI0VePTwJ/7DC0a6yKjXhAbmKY2do2wF1XpiaCdLxEnSzC3JniyA/XI1Znzk9Ny1
IOBARGaJKywaDGSoiSzHsK2yGwlKDje7j2hJS47+t/mV3fveXgK6RoBK90ZjtsiBJfzcgGjJy1Ol
H+n4sKXeLsqfDzOWNRMJCCb3EDKYZVyqqwpvwy3CVBzksLGqW2ejE5HIGZn7bzw/DDKEum5UCtXQ
ciP1jltdvXLpQbKSQHfAWzk9WKQ2ZpbN/q8OaNYoispARymeuaH+JcEhpEZ+gy7XZBk1hW4sS9r7
aYuW9DdEynBgsPB3aBmFerw7NVfpZBJd79I9BhVE6ibuXxHI5J0bx29P/dcYK394500Tdmu7/SU2
EN7EFaCtYdbSmIPJEo3ZYEXGDqINPEQsLhfZmQVg0RRrPZX3vEYvX3bx/yf+2Vd6pDb0bxXxsqcB
jjkkUPEZ3AA9ZajxVI0g9p2zue3/LP12bWtDZR5Ke6Go3rgaNTsESeplOlPRpz/TSN3OShid3gjg
rukOV3pX2vQtL37Pc59k8llC43NptX06nhf4hl1Q5oYC0A8RS3Zg7J1/jJPwfanPcIXWN4Hq6Ai1
TTgzDzXFLbEGShr1xTTSGpxX2EBYFNTSCq4wr+BhdiRKyz93XnFRipVD08mY9AC4w+6B3a5cCS34
vzb87hN1NDZ9DxGaAMbXPI3H4TqxZe1BtKlkxntBb48DkoUMgbaXYtGblYFI7dcy8C8TdtdNQ85Z
IED3b1TlV7E4wjN25b0Q45zhVGNBsXPjP7zSzsEN+03+TMhtjbJUItEnYzAtUzLOnLuvF7oK73FB
ZHBZQTKGsfrPsGl1lta2eb3OonX2ON9ZCmTTcCFFwAyxf8P/uJqTVBZeAOCvl+Ko07bUxlHWJqXv
QHIxdoP59qkFNLTc8cy3DNiW/+eQZIW5/FJr+0x0EIdbONbLJTBGn+q0B6cz2q+sDcC9IZZLQQXD
0OLYiVvRUOvAtQc0FHp1hqzc7UUcNMMA30Sv6O638xoF7cJPi8QNbcF5R2nwIpCXKOJZ02AG5uL4
R3gM9Ek3dWA6l1r3INJ4TTJvDLP8h+KwfA4skxjmvhT6l0QY3aL5HDC2LxGMrni7RkNZFcniDQPm
cCJ/541NtMMFoFCtyfOQ7ZKaKYhCwEpP0QwHnPPnWPugJgvlCfgfczdcDdV/0rckc5BtkljG5Tyz
aHuwLMDt9QeILv4Zdj8bNOrwHQmGxM/1jDkAWmWgyoRGTyJjwqgVDt4AlKXexczWrmyts2Uor3pz
bZwOHHo1Xp33ERlvwVJo1vHw44C5kdbQEFedq/TCg56d4SoT89EdowPxCGLL3KHEKudMbYbFX5oR
wcWvoqyK+J0O+wfWU8IUNQC4sYDX/tWMXN3ra8ph4P05fEM13hdJn1rrCDLneHyg/b7gC6mbKlme
zRmLjpVU2wfe4nROfcYTV1MUQv51neLDwodWZSk864UqLaDqq25i4ob5sPu4yWKsryGP3YRpq9Bs
Vgx72JZ3fsrQTQpE951LVCS25k433GEUsWeTqNMtRVf5cHaJvKMhoKFq9cTrZ5yC9oaj7W9Xxo5U
7TqhBxqoYVf9feJHZ/5r/gCiNIm2UZcSlvfrfWu3O10C442REg0qcEg/V+7/ueTUz503VJ/5R9L/
zYXjvX+Du6GCJXqAvowbwRGVP2L3ipqUYJion1Tp0rJu9FIvh9YlLIr6yHtCN4EXjkzm815t1tX/
CLNzgMgQ28eg81mnG1D9c1VC9fSSMGPpFMhi8nF13RhJc6tK5PclEGjG71hNlVY+er1bHSedWnBb
mz4AYSyBgA6u5mMcmP9E5Dzz6X+sLa4n59e1VW7Ajyy9gUtf8HEW4xjVHLoUdPxkXEvPxeVXzQL9
6jgeHl30VI9M0UN5f9ovuL/Bhglv6PEr8h/0iPGCbH9+6ZEf4Sn0zY0e8j8k8rzOlbNRATQaFwi+
vuyD7iGOqjyp1yEXcfGhTC8KWHaIORs5IFbgYkiyLmQ1RIVQro1CGp/dMILSLQOoolG4F9ZmcI4K
pTSCa/QYO3tRzhEcrOLnp3In1n8CX0uBJSLwV/9wa+jtCu25PluoOJ4CCQ4nKX55HvNr1oyvvK1d
/Hu+ZhgZIcYuwE//VgZ6aAwsgTOdMYx3le6CLMF8wq1C1vPGthMbXr+sPW6QNf2gzxkl/8++MiYj
WGU01SCTWXosjc0IVofMmPg54nkYZAgGC9wzjt2Yi9K7zi4zDicdeCMYgFouRqu/AFuefrB8I0FL
XrM1sjzphxT2fuajL2YkhyfD1VZUTlBFi01qNvtcmPIV/U+xm470mo/Q/2GY/E5k1A+Vc8DioQ9q
J2pqoot83vC2y4mvtBVzTcH0OAvqimS574X/e38BHQFljYQejC6wjJ6f5cETeyhOC/APiihrDRmr
D9Phtg84VpaJhJ9vFuUYighlBbQrYwTcwPYKRrU690E8D5xnFT1n8aG0MZI/B5sf6b8lUSG7DYze
z58CHV8PgITo0rbffvsQQchU1RM0zR88tIMOLJBiIem9lDI/IY0Ump/aOESjoCs7O3tuRKTIL7kL
4fCUvvj422yVJRm5HCzY5Qyy7ruToInq98BVGoOmhAdQOf+mlk5cZIdc2pKwJpSKA8Olj+BKvFpx
Dl+qHBv3KD4qSubKmHkmD6EGksn2Lf+B1BGFT3afyhd//uyyMgZEZWNwkJpAowrUycnQv17TCk9e
WsCmK5C4eHa0J75Jetch4mrA4UU+/Go1uS1X07txiWDA8YT/Io7saBC7oaHEszfR1VGJHO6jk5UI
07glRnZCTS0Idljn2/7CsJVvNvR5sWhImWu5P3gddZli0VfsbtFlsvRB4cTHDTpmuJFts5LnOI3V
tZ0cMu6/lGGYDuxoUlxQRpU24H/updU92Zmz0NQt+h+gmvqpKI+l6RyyjdGrMR822+XvDnpZDRDY
ijFt2UeplQE1XpGNlcjGscYl66UKOfQLoACdyM33rjdAIeulATgHfjVWTUj+aQe2GVcH00QfOorA
o2jTyGVrWb/7/DVbtGSZc5kxI3caAAMnxw2Ucrh42pAQoOwR5JkfqqpfGTQi4C6rTnWZIEgzLNG6
hLz/DEXlWm949JXxj9BjCMU+LnaKcJyPw/i3Dk3joPME1YLJH03w0Qdo8JKgV1A/QVUwWiZsbwM4
M2cuXiKvzmOERAYy5KnnFLFWZjuqbLm5cuZKXrvUwn6+/v14UFr57J20K5Zp0O/kH0Ojfw5Wa4ST
Jx6W1lFLhgjKqh/9Dc87Cgsev0n67tnkDiF/53T0B6fJhovMpyFcwfwQIxLxrfqn8v2ZZkWnEOfN
RySCllkCIMFYVND/2W0ffH9vuRgYiod28t1aFXAqqJbLgIR51I4RDlgDwpKrYSRO4m9TvJCDwQF3
78EoHyWMlxS0AmvhKgtRj3bX3jGL72MSXLgjQBmjEP5WP3XBBt2bNqOkRkuILvi8/QQcIxEcy/gK
WdCOEJRuwoE2SK2bqTAETQsoFhFhepPbsZQbLyR6oQHqxSC/5rJQl8xGhEWer+A7rGgvt4txzBtC
JyafXOmpTTCT4Csf357jJM5WU298gzMYCPLBQEh+ctqmuGszO6P2DrmEYFTn3msPEVYnyjejmarH
+ccQe9BfbkrWCcr5bzh36N1kjKag+vz5PIZEp8MQDh4WNAtkvwpVQON7EoyZ+f9nD1k5MSvkjNP2
o32hcBvA6QRASXz2kY2o1/zTFH1mcSJQ1IyH1bkclWRraHcbehHGiJDgcn9I73zrc+gp35iQWLAL
TLvxMvRl8i6cY85+mlxp3F4DAg+JGDCD6/GWebos7Dh9ynFvfxxiUwoxkna0L1Y67KhKULzACzn1
sJPsuJVmMOzHg2oOISshzZK/ATa0OEmIFOlJzdbxlG9k7RC/pHlp5kdtMF9xrOcm5vmIFX0FIVQ7
9HLQa0aXyJOrieIMeTKAYTYyaPawQbxGteS97wdMPWoF1tU0JjlxM8B5U5dQhkG6+LweeAcRue5w
WK5WE80QQfgwQ9Y1xLrdNoeY4/YEuGbysqLn2jUiHXNJAS7zWGbiSCh57/jGoRHnV8F/18poSmpH
igoUUn/xw9pr/7rMF6aF+scyv/z9wU6uvf3ZrcGPPj4el9wOA9Bsd4SmiGj+h2UG/D1Tjn+sndPZ
HrRAWZPdNIdrCovWDWgL5V+VAZkiBq6HDkh3GlNKW09rr7ozbEuqfCNRTaLRhPc2QZUiL3ZW1oBq
hlPF0lSt7ba2KQUUI6YBsVQpkD3rLIuPCqbFpRmW/uZDlXP/z9Jl3MdL8v9uYNcwsVDXFKvZocim
F6Zk6DxRiyjTUmGnJabjct3y/Uxce2GqiiyYJm7Xq+NLv2wzq7C5AY9HrOcn1rkElzthC6o0sbNe
OVduPwiRoOZ+oiFJXHfCS4Earny9eqtVToTko6/LnNGQKi7n8A424FMaWcnNMDThElQ/dzIbwe0a
Q8ZynJipfYF3Oe1Wj44tTjfN/Ae+OvNdY0Q4Hn3jNII5x/PmNHN02qNVkx7I3feni0XFdXlJfkDE
YVpK60KiGXt6VJoMNflxfMxWIE6sKkZxf5S5bLvoPoUDGP5F4RwgqF79C/i5w/lIinXv94tj8urq
CUAImlXSgs/XTo67IFasiFDtPwiuRDOU9lmE5Lkjzm3YqMc/yJGRqmi9bauuw9eng0qNcWztOHP4
9FItQgRqJWBHyrW9tB/CFva/caO3LZrgpNR4IcPf759jdVUiN1XKepFbw9tx+CwPJmw/NMgm1izE
NlblXjt1a5TQxfC0j4+n71ICuYw1kyHW+oU3dh1EAdBs9DHK9bexLQlZ7W1XMWTGJNIoPO4QMrBg
BYdfe+rWliLWKcgNbQZu/kk/WKa7xKTBE999oO5Wlp9gajikpJWkb91PZc7iD04ofMOmH7jxq17N
UNc0SgudKT+OE5VKQ9os4Xmid+gdllawll+lqs1UNLcOoBDdz9eCTuSpcNaCT9nNO7tF7DxKHCPP
5SoBobewCCdFxFh7YTqzgKkIRO5rDEQe20NCfyXHe0wTDfcU4fROCBIrKvaXWm5v5gjyg6uBJkSt
3An1dD2bMtPAlUtwUQ53iRQ0qTgNQCjY5FTOAe8owgZgzKiPrstFLPXLPMNQnyB4mAp9s9nq+t6+
4S6rne5LqYQLo5/5yT/WlEEybRb4UqVKGg71XDDeEoY+IobP+xdlwAkKUqGKeYS0MZSST2Tg/v9S
vX3Z5Ql3RDavIdfGy1ONUPGGLFMuSGVToI2MMyJadXLkFQc4IKZE50PFkboj7ZqJCQq0xWk5ocJ8
GIYYiNhnxuFgMl6FbpTiDj+NlOO6Ajh0mKhiF5aa5ErJgNb4wy/NNFsuRVjIM71QqIpfDwxADgeV
mgDdi5fOZqVGKp9MDKTrbcEBhOQtPTWXgy/6C+vsL/xTBy9vzRkR4pd7Yxp+oi8o2L12/+m5jOEC
c0A9wHW+LP8BZ7MMyrky1yVyEGa4+RuN5WIDRpVaIh9FNa9GpWTVq1kUU8pgnolrZaFY2ndhE8zN
U3RErgzv9YSjwea59slJQ8dd8RpGI3Ol6P78wx4If6gG+l9q31ZJHE9Wc1y2w1kLVQ261gXr6KqU
j5/5yBVC8wjWo4E2qLZcqTdjkJS6NA9bFmlFdG4TKO7SSnAUhjJnzJ8StOjP0NkX3Wu4wLesGcKl
dmyQsm2QBkdUmXMUxk3SZtiHddSaZ3saMboHM0a0lkjyBPL9fW4vw/bbiggtIgzF+A0ZYH+7gWNT
1AFey2vdVXPlbzqsQmz1RP2AQekFKErIS5StXNl5UL4fkO7C1DYOSXMq9+mNlxrsNS0deGSK/rVo
FWj6Fx37k8g7BlxucqeUfrJL5QMf+83pRS30tAW+BVfRZCoekkEV/ypBn0z/kNHMkfGz5kTXLErD
ToTArZB8VR8TXcvHPH8Tth1STqQNXffhW2GUU+RAglcumny6cueR+4gf6U8n9ue3bdJEQT/tPYbL
dBmbt9/ODxJK9bPwCG8QKKZUlRWK72WsvTrhvfDX6KwHyDySsmqXOpXytCVarhLIbDoDDfPGtWyk
kEQZ1iSIwoqqHmhKxdWJDKz+g9tXmhAduWTYqjsCMe7icRlRpt7GUYeltk+UPZELD1pPNnIdMUID
yVRFOwf9Niq4NTv6Kz1zOebdmjrh0azskHPRpO39Jy9g4molnSMpcNscJsUwuushNWgu6fA9hSwG
CZgtfz6t7WenxiJwHw2gNMpJpUqHmVQm1Iyyqx7Iu2E2QEZOKI2GB4aez+Gb5Dv2OUlsng7OuUnK
coEwCVZVfhFqUuoezwfFPkrjpktZrHTwYGIjPpTmqg8f1iBBbOx8dmc2VWRmcf1QnytA6BKmFZVE
MczxDv4U3OqAIKEPrQEWpQrELPMx3Pyx9wye3HjOgkfXtdl5dMKYO8s/cfUo9rG0vWb9B5xR/KMM
1+3xDH108eXREZURguchY5eCTSGFlJ7zARDjs1n4wSNFYBW3lp3sZniOB3Jzhc8Azn2EAoM60N83
9eqIRMPULnKM4cd3Fam5xbpzVmPzLuZePZoAClqUJaRvIRLQqgAi4hKQK6nASIgISLYwtHj1P5EM
q2u3gH5liFm03UAZhIeKWotqunkChitDY7spCAn+4jOBNgnMth3mBRGc4hVDgHXin6WmfhNPns7/
WwITGOW81THfwjfpKKnuK/IovezDjkcw5VsxrF3TsWNHrBdrhOGtNV8l5eKtSg5OUlsg2Y3WXkU0
3YfY8raNK14DdQhQnTTHGsU+/isD9bRhqrv6g9onNNpfgnq/qv90ZRVPhr+WCVVyc95uS7/rCmGs
e1EPHFCbjB8O8497MhF9Pa8iacFhXkPNUcgWRqZ1tvy6zrOVXxWcmweEX4dF5juSFutjYyiNgaqu
TFvsFF2y/Q53xbpJ0RsjPEJd39DwI+4VyKt0DQrUnT+JD8JvdsM1eli2RKAY60ezNMIc2J+4aqzG
zTd2hfWwV4fRaJ3vz9qjiVLKRvgLRbMTww3YMpc8Jjszq85wZ3mzupBK2Fc6IgShMEP36gEVRUeb
BZfvWisriqMIog66CueNuwtiMQiJi/wK/maN7MAW02HL148M8jeiYQnGtXZPW301vyNoH9okP7ju
pFYnx9WSEwuXGA0U/ItH2JPyPUz89NJC4pAqdsyBPCxPImpy68XEV/dW1JgraOMQ7omwiknTt6p9
R4CWxFdl8rf1G3tW8Vey0pqqQgBUrBVaTgjmW53b9CzSv0GLocr/Xc0h6Q5Y5YHxo3/hgkOzmMys
jk/UdzW46vEOwc5B9QR2eV7rHqdvNi4uz3vNZfVD7pOue32cipFhwQ9nEw++y/3iNKeokavfLuLt
knD7In1qgT90rcDj27wui8QrjTAhhbxSXWY5VLbWFEtA6YrhAWSA5tGcgCEGK3fsGG1hKFkPWGCd
2/Hq1VJau47pHJhS94OOve/OhRAvu7WPI/8fFjMS17TTDg2nZOBMr9ctErGNhmcT3Tju38DKMAVs
/LFQQKyhvz2PWg96fHcnGkYoyQDPkLGUe6a+SsRK8uxYIHJdA5YKh06hVUkTTh3ORxsmOu++qp8r
R8QvBZ1ZH2P9F6aS9FXwCS84Bxw58nmu/Ody0kzoqsIQoFdRxATxrSeqCw1EWAxtn60S/berp2NK
HDGMlmOuC4aemIWUT8pi4btF0n8d0UhqyGFFLNCq4uF3L54CfEWEmANsYLIxjZLObryBuUvPHk1K
P0qvJ+YfQGSOEdAcY4pSv2eXK2Q9mYTCmvJm/ExPMj1FzNjzwMTXonWm1sjejF90hEBtdxW1Cl95
XDyGiaCGt2fBoes0aqklPR3j0IY1PwTJi1TseOQfPj65OpZ+6COJSMDhISWwkIyMn8Om4dwYz1AF
Oy69ccOJgY9v6qIGUrUy1pwMDu/AKUkrIPVUr8AnbVyxKU5recOq+evVbAmNCi88TZ9RIetlN3SV
WSn6+2v/crmkcepjzcW5mA/CrAk8Bq+qcL+S3/TOr2NTWKUWl1t4n2w6fLX0QszgDOna++UxXWu2
Stdp5qDo6tWTdZ9xC/Re3e0zm74s260hJeSOPbv9KalopZinxscmiK73XgMhuvM9bkAWppGsxddc
uS4LZNfdFqbuDCdx5KPhz7B8Fcbe5CAZrOVLfAKEcr6A7neO5VU+018L24roqKnwVKe5LYwP43DC
NAmr6dR5yuRjiJF5PM/Tev9+x0kfHapjmk0gsb/8++hhB6K7I72ChqiX73kzZaloEDijBW8N5vts
Ihpv5/YAwm10da/Ec8sd/YIPhxzM7TtQz9jw9uWXZ+TUgEb+uC7oY28VAZrfBZKiBfvTAm+oMw0A
u5DJXPA3MQP70tRlOKVWVfGyLbruKeLGuxP98hjxxGjI1k5OkZerd97objSXXpg1Dr7S/9CHp6BX
cY38S6WI6ZKqZy5hNY74kU8xH09noXA0Gef+4gwfXFx2n/mF9JzpsgNC7G4JsNRjjdo1PEzbOCFI
8LxiY+W2WDB/xWCtlBiYNwaTSYToTMH+cZ/IlBEif7QO2ultlhBgPS/CjVx/3/T+5eQJ1ZN0PFeQ
7PzUIguSHtBUXrmFq7lBKhMpnx3t69BU2ofusXBH9eSH9OB+I3zWX8V/8/5oHAOL93OpHx40aYNA
DWy29jwloekkmoNq2HtZ/XGcLK3l+DbiCLAWxEswMigm2qMA9F+ULfIqEOmCLzVmNyCq2CV3MEwO
2mWktbzyJxt9aMSMYPiPe05NPh6akyC5uLK/E/eytmZoEgTLW2XDYKPiOOZlOny/fzm8p8mhIhs9
VDEm7AHK0ALzxCneMgokrUlzBrTq0OQOZ+dsBTI5aLxd2CJIUFw0dTwblXYiuQ4Y1/uxtqqBmI0z
L2pvZc4gVajHgEtzFQ0NifG9ZD9VQKW2xUhpPSGE7fGI5rQEjPEzBqtchjFQmTPKFpLBq0lSVKJF
Yy8fDhAgJfAi37qBE5qq/zmSr7RJrOCk68W1RezEVIGIwE0MuJCLHOmEDLUN1fF9zIJV0pB4GrWg
oQKDgdYAbJJM2y2sWzNrP3K8cSxjXmwBSbCfXqDkJDNf85LuOXzbMcJEcU+OT9ZLCE0Eic4bmy2/
aZwXGWCig7NTR1cSAMmtq1ZKosOFt5JcJQBJq9R+9rzQX+I/AU3S7PdM63LTPlxRdAVAF+WfdKl7
cOYg++J5F11UsFOUJf08Azv6tIB43TTRh+SNvgUIBcwLixe4Uj9F3akcpbo01EaeoiD11E723sc7
Oocy/b9kLwVM8yeSn74bKysZjhk3x86RkuUUe7cWJ3dR88/Vt3nFwdS0hOo9msRFKA1WUQp8bsQ6
+Tvhn/nS8e5qg66ajo2WgEC9po+PHVwQ5a9AOXG6QC+kjOZIzMijgbDZSARbuqjQNc98li0PA07y
sTijFm6J+RL09boxQ7ukd8hEiogJ9FwhY260t//SwyHsABgU0AL11qJyVFk8pZapkufnftYXQ+M5
UYsCjQTqYM04N/JipxuCQ8zpCyicx07Qc5S09s9Y+Uv3Z1mLPGGZyyiLCYkwbd7Oz27afNqrU3YB
t5aWsoEfTSzuzJsGYYg6115aIiwmlWATpItf83/TBgAiZeBkRkCwYwwGRGcVIeS/IWj3uKM6Artq
UCnsBSDhSJe9M7ipFUrr356NzH6IbcnmOfkH3ygbf0G0vPVdrr+mq98wRvSvMlt5AECAVEn83T/0
HXpMzHdrM+WCGydsorf5Y3/g8suwgcWCTemXUgyz8810q4hK+wS+e4CcWx0kqYYBiGuIxu68Ldd3
nyJYE0kfbunLZrXyB4E7Smk6CBwIYrYnp/RLuaRzv6bwLvXDGdHRto08sVJWvMj9PSWECgvZaW5p
ErvlTa5UZjU+bPzvoS426KovyITZHTym1bmXhHV8P+mDswoRJ/xZoMGr3CXGQHW51df+0eRt8sDG
d4WwyVH/ZDeuf3OaBM50TX7mdDEZayQu79qdO+5BLNiit7AIewpx4YUDXkLWBufYu+fARnSVIkJ9
F3PaOZ43Yttr/vsHsTewBF29ziqdE1HU2LnO+/lLeaKzLw0WbINCVrA1Lxhwq55g4sUSdPBlTp5c
Z5M3sN7NVdUpsdbAwkE+/gZ6sxh+rH80ix8nUoWwqeo/TO8efDlOJuthPyyiiOHhyJHGT/Zg9PDG
mcG75ULES1s8KaVGb9yKXvanx9zrJ9vJ7+N8BNdlaJ8rpjhSkdOxIl+JPBwWvUt3UOXX+UwthPZL
QcfLqqMTavywTSbN/u5d4pRSPaZd3Ls+6F5dwq4rUug1btHKz7uzq63b6HMjCGnZ+TRlx5vHOTDt
r5VkCuEqSyX4PWbehLJdrvLoHjDNNvxlywNQK/9lrrlnqRzbhuiT6ZFlJlYPGLYd/6NqdwOC0+Wb
1Obp7R5cNWoJNsvE1JCkblZ9cmUHGdS5UbkaDzIRCwHrP6arLaSq6tIgMJrfVQ7XwuTJ1tFVZ6VH
hnCzHyuMXmmFvaFgdlelP4lUOR5NTOmQO643j3V2TU288sMisTjMu67HHHpA0FGi5ohta+I3wWnA
r0B+F7PETf9ik7FNy0okDtXKZDwmx5FTNBVP5NPB8WY7yoP2dpeWiSe19G6SS7mOj/kXycrbuKqk
IY1NJ8luzT644JMbXFkthrml8F/l0aUi6g2ktP164Weuii3m08xEotNPsc6vEe18cm0XdTaR0MUY
47q4dfpmxdYN97HXb9GKMZfPolYr5hXybRjcM2BaBVNgtI3qQm3nWDHkZskVa6o90sw2JzYoH9bC
6NdSckqGNSrV6jzkMmAo8F2RHVRG9wSsv6A/OiXIbf3mx7Ld+azh+6lsW5OVz/hwrbKlzubNLbhT
sus6vkuSQlp+hCcbGWWdQGEIbWgg7biSaVZi2eBCKD7YQcBkt5MJ6ZtkK0XU9yctG343KUC6uDR+
UjiZoRj/JcM2ZT48f8DfgJT1gqMnFDeeVE4N9LFUPhXDrK17jLcy3OKhmNKBJszrRWr8oCQDR0LX
k4jTwSG2UmF/sA8kVXsUb0On+eCsmbi3Y4U8pQQeFyeS8IXkTJ9JbWgCtyzD/SdffY48j8SE8/pS
8klLg1UioWpQhI5w/kvkUVE/D0VROiB7CiTUxNsP+GFe807r5CDyxRqXh5drnAk+8zmdbuKPBqcO
0kPyPWGvBK/InRT+xyvA6E9JCcVVAgyAJkjykU5R+NrqYNPpZq1dibbBDmNZE2IqWnJpUqvDq3D0
0kF5V6x+ucng+iRPtz7Vm+iiIfaVmgBsSDlCMaNnJxKbLoNL0IwPTx62phsLYwP84DAuXDOSP5EO
W6WwCMsKB0ZJnKDD0+gIaEIwlwBr35ze1dAihAA5+ie8BWLu+lCSl4nF85SIh1Su+WDGNy5u8ljE
bsizVeYY2Pp1O+2EeFQ/cwavlVs5+EpqN9G635S09K79tz8A0G7R3M35/2IEe0FaR4V69zjwj1X2
6m6ZzMtnJz7TIIvRJSvuQJ7W4rWCI4UCdp8mdiV8S0vwb7CEgxUIBt3ARSQy8kTBCn2CnD+oPwAf
JNI23RiMN5XHNBFZdc5GaacZKOKOFSGy0F66gitfLONcj/OxbAnlAJokN/JU7+KAt5EDwlcQxIHo
ASCp17s3tEG7c7LJiuW5lLvnRUx5TR2/FDw7L1NXvhbj9xUF4INtLOKpz7SmA6U0w03D9gasfxRk
9lVNQLJLkuqdRQ0PtMWoISWHAvuT2uSOCgtDLbSl5w7yVJHqJ7B6CmAhzWRRPv+iinAmkpYGthQx
qvHX3Qf2M5u0wqTWLGutHFHl1zLTTEDgLuhTg1dvD12xDRlinU533fgkgRNn5n5ufuGnNQYWtudg
v5mPD6IcjSSc0ESr12bDIpm+t/RQU1MoxTdkyf2qC6PjrciFxd16vFmy/5MsdhxIhkr5xZOrhlve
lJP5VdzLtUgIQi3H1HSAG+YSYPLxvQeZ9aEIRlXXFZgBJCMbXBYaD+26spQH3FY3hXlY8bffdaGX
Z04Ff4g+AlKdWA6gkCmaiMXUBerohv/52QtomYBOcCrbzVod/iLfrWqJRbsq2xOyf6baE6Ib87dB
tJ2CCXIkVRQTROiQ68FOBuCxjb1TPkwQN+fCDU96LHUcxPJq4V2tWI0fL3mHRX1Im63iWPiv8YWL
lCs5tX5kJCxjXDJ3oG4mcziST2ibXr66xOMXqSV8lZU1kxsC+BwvTvFEHB/SsRYynMpEP/SpZiq7
tW1bpprIMAXlFPM+VFZqFXhRBwEiC1Q3db1kCHEAzsRRg3myBoEAtE6Hknjh+sik60y71IuMHe3Q
X2FzTDPy72oTUeAyk3Ex/xjI66lBptPTO4871EPrO0+soXh7XLg5V9TCtosQH1GelVKQmOnLFRnl
B7iqqOxj4xVBypmNrSEBDkmfMKzlPez0k5fQZ2dRE4sjdf3hSkTy+USITKXq31DGERqCzwaXMklt
pdbqLTplGh0azJ3YEBskhjDa2Q79iUOdPEuaotzwvV0Nmc3PCfVO2SxtBBqCXk++scrY5GwvpLa0
9sBNNdJ6LDmxOcCwF/nEYpFR+W/CbDVnnapJcRKBVlO7O9PAm2Fg9S8i+RlgtuEnBtQASeBeCVp3
YajDDHcBprX1U6JuLrETFUIRnB5pRVkxNnXixYZg9PovaQds60FrzqWwc4NpfdviIhDCUFQs+PtU
3GebJ1IpbYAaaH+um7lwPcJbeBlOiYSOnMH9fmxpHRt+cyUGbf2I/nARyTviRQ6OGTqi6+YD31r5
Of3QQU/a6aFjfWPYhbToj6Jp2Pi5wCm5yRtFB4v8ibhPq9+OuOW7poF14uDPPU51OEYz6fKlzbZc
uLVp3CoxvXuUCBiTLXDAf5mo0abWhVhlobPIDZtN15mrUgirk+VaLFyPQnVR8okMbc5Qe51jzE5a
iSHV1eGMtxJC2vOgfc+cIdkeuPQmfovxNgEfMc0UjOR8zvmjfFj+9IbzKNS4Fbv8od7Zu/9biRqx
jK2bIeM7soFA/mbgkH+VEIouSDOJHaFGEAmPxTtTrrBU64AmgzDZOqFFwNEoK1IYoGA9Sm/sY5Le
T74xiARtXgmI6Y+ybikS96pLxf2uWfrczVm8D5wT8/CJ0luPi3fe1lbK6YviEu52nrL7iRZouWxY
5DdgHvtUP3tL7t0BKLhKvP697ayUJFEUX9D0GEnTiwtBth+xqT8vmXh2MkJem+M4vBGFOG2HuyHB
P6VUGLPXpVvwREkWXTzz8Aosmgtk9tq/WHjox46mU6zCbLONPt7joRYFKEcGLkvHnjZH+ItxoVml
MuzJorWMM4Sx6j2Fc65o7GzHLZX2m5GjnbP+jSoG8HCyteJa58A5AaIuLLK/iTXJwV08Mk20mCs8
xby9kDzNym9gCSGZgJVceUZnPNZbVRfMf0GUUPi/gFREhBAQ17JCeYcB6sKYIaqKCidQVC3r71Cy
31wtWsuzFV1VaGX4gJcb6j8Xpg3DrASSvfyQKDOpONvIR+ZpdmSraHkwcEUVCnQ1cj2mnND8xPFU
uHcMufAaX05IGq6iDk30cTcw8cVsDbyTAtTLGqOVcd5aojvPU494AaOYy5mr8a+53fz27Iaktkoc
26BTwRkdOEOYhYn4LDEQ7VjAz9hki/aaq0/AoB1xkpLF2x6w7gpxz0ILl5mnYOlx9w0Dia9tJr6C
+Ob+wxE25Ar8+7btaPpnzmgjumS75ZjG4hx4OqxVX70PB2C/1LeZfVoX6CppxLSJJ3Rc/SRqHvsh
yrZxeDHPoXwGYc/d+7raNwYOmQhO9HRrFrjgh0MGj7p++skI4PLfWIPMxMmCqG4WFDHP0iAPOEmU
tcZRXZDENiaXN2brKMdKAfnfuUH6wixFnGM2HlmU07Z5OzWdcqenFCXh2s4QxJ0DUOhwZmfGzsFp
IY1RwTzsMzbOoX7FpVfP/Zj76finP31J9fPAhT40B0iMSyzwAtv0z1PqQAXqd6NPEK0QU3VXbEvV
n0lMmrmuM0xok1HkFiax2dSKTphtcVCKrQ/mVP5i8Cx+umkG+d8oJqIZMWck2cxokG70G0KORPLV
4MDU1sne1P+vt7cUHdiPb1nXvOCaUWnORK1Q+LtFvgBiSvZKPhweMS0Z+4SXFLV3ayBxBdMnNJJ0
aJr/cyN3EnINChXobaU7nHnw6NQol0o1fNWdRfU9C6SwJcrjm+X76S1wfyw+x9TbIQqn3H1oPpYq
XPPvR8TdgxrFtmkeUruCAFYW3aX9MyDElV+LS/PuYOgJgqq19UVcPS3VXjUYLWhL0yg/mOa/8R5e
mGqDbrc7KGkK/TA0bZz62d/2oilNiilKyfcP4i/c5Yj+Vj8QZhh4Hch9NlfHF4rKxG8dN9EGkvcs
NZ36cG2wiA8g7Q16K/QwYj96n3j/hmFPiSpwCFRwIZFU3XMH3GJjMAZmvRrJXeVq2sc0Qiwm2Q9Y
3iBYy28miMpLaU6FbZ0rYuBc/wmDK2nbrsTCROQ415yJR3yMZ2k/ntI2osdW0tXIuQEjoLhJYaWy
vo51L1/1i/6rWX5FChBzC+tQMbWIoDC+UTM3pPP3z+0NLLt6IsldTZPo8aFTkiPT5vgWN/WZ2x8Q
emA82p1i15G8+wKSw+IgGrL10Mh8hyXDMs7csgLtuBouilnv02aLNd/17DJiDZv8SJA/PYFrfm7G
aze09r1dXaqazzKtpuQWij0y1z4T4qOQ8uOG548sQp8QrajePqMaJWAppSiv7jqENyw/6N4Gk86N
hCKlfJZF3MOJPAZugMjqgA4M45Iem9ZRj53C/pfWOGp48VY8DUlpK4xaLX8Bd1+OQoTDN7ZrX/Mq
HoQvbY0uffvLD1qPjk+lInPeWe5wvfOJ9YoWeS6cwMuCP6+G9Ckn9OjqtUg5EuGWPlN6Ly6s+N7o
lYX/yt9WrkXLRTVDYtld/Mter53veNAWZqe447ER7IudN+U7R9fYLUo5xFkIifbXjWl/OgeJjhSR
sSrJccejQBiWCW5rFiH5T6XA4rWebBhnWMSVmkUm4NfkeeKEGZf1NtPqDdsaIu6OlYGa5KKa8ZWG
/Q4XT/Ez9Y599x1wGF0ibr4T1DBaQ5dOsA4S83ejUyPHmYgyLYV9XpRlE77gQ4f4hQXJNwroBxZy
Qt6Ks+X/WjsYXCBgwCHWg5DVUAhJl5i4JdZzs9nW+x1ha9zM4MDi9fVJBwGH1t1YdFHtsxZ7onNR
sqLnKA1BIKOGLDYiqV8MnytiIAgda4eQw04iEhJcs9tYarptQwpDrT27JLZuCj6VnhoCeoh0ynQ2
+sx9K/Hu0vYV6hP+sijGMZQqUkc5cs8MIYsBNMNmxopbnM+10abkrmaicnKpRLcTKA7yBCx9cMMQ
3vZNQZWS1kybIx0y9a9x3Vt2aZVBI8jnLrKGQHDXBkeBGR4MMogNVFMBKAAPI/TCA98FbkxNFKnY
zvejhGG3I2BukxpDIBBSJcKz4jGCa05ScWP/2ZWeV8phlOInZfRxE0gpFyl9tQwiCPNy5efYRIRu
fMy3sTLHDSQxSy6mH1XoC8haQiCmBSwKzvHjnx0pFxD1n1DoQ7VqPnW2DLPbjlULrQymhjwQnW7o
n4k2HXV3cGaXYLTJxYoH9upL7xH7XySgofhBDNty4UptlL4R7QaM4ds19Z4EkzV4GfoL0yOvXoh2
VlcnbiRfsQo869KVhKF2j9GVMLSJ3W9RkhTmuz5B2MQr8fYJYNemV8EYizvPStMLQXARJZqReMFL
OCOZiJxFxHECWovWNUbdlF14JuqvQBvmZjz4K73Hm6mj28D4FQsYn5fkU5oaA2YPJtapbvrKYJpo
b6Hh2PBB/MVS1KAwWX4uTbUHoyGKcIOs4XiU/iKryAv/9pEYc4Qe73mWV/lwNoofqrF/Ziz/flop
EeonNvucF2Yco5A2S5skKGQWpMaPniM0/dgGs3NKyz1oT3zMDhnUVk2l1rFT1nIfl5oZhqk/94JA
Fz8rQKuUsOvnRXVWHd1GS1KoPoGy9HjBrsAqgvgVifNDmwzOlrsWPN+/5kAjZmL0N5KoA8Tm+zGD
MsxmqJOQEbHOfnNDDpS9e9j6RQGnv6TlUh78L9wG8aJHIHKpCBSe1pBE9ZLeumeLqTBCh5BTCDCR
HNgJ3NCWdeuCotX7VrPerT76ucUPn6NT/uVRiIkZnKrwgMvv1WzSHpE+daMg1Ablc4+H4jMOQmyx
b1t15XstTQbmtZKP1+BIVrX83BmbpCTsDKTg7eSlV/RtvrHdMK84xY5yElVnqsDdpHU986GKP8vc
qNKdOUcWr4UP2DkpeHL+NRmSGEyAbruJ/v+oiiMUzVa9Ph8ADbHXehIq3+3KMrJHjaiy1d/4EcN3
yAoKlkvTAyC9zpiwiE1iHYaRPqGy7GsyCuR+42EtlkVlGx0D+rr4f70UORuYUqYRZjQnTpHzGPtD
gYErj9fFVWhotT5c4BgOtUa1NbtQVuuJVp591duOLrzblN4mv9LmU2AvzuxG7hN1qOnoWr131FwL
rbu/Ox/syU6sEA0x4pQZElqI4OMPLxakKsShOhkeyg6rnk80SaLRRmPq1D2WIkn9U+UM7nDqqbxQ
gLkWv8v5Wr5AePG6GcSYve84aw7hp0iDlbuPLnHoI3bu34+sNzVMlHLPyoWvLLQmyevfQbY3smAF
gZkBRqsR4aOP63D6en6oT5ir9iYBQn2h7Ml93RCGAEMSFXTNc0MwyDc2H3epfHCVz7PPIIc69sLB
+McJdn9HUPcU/PT3hNChA1XH9rZWS4zPB2LLbXLWsHzLYYUwqnKqPanP/ML3MJ/LekS/IpRQpNX1
fhsJ9j23+B6A3LjnkR5VdmzCLzIkivY7jpQJRFuS4xoDEB1TlvMoIbPsTpDDlitZatvEpRyvoGhs
wGZOtkDIDMKZTkNFMRl3JSKxo96QPdT3nsqQTul+9G6CP7a2srqxA8eWfjgSEqB1Icz8cybCtbFc
f52m5oE6BIZVDqq261zVC9f0D9bAfRi36s/CCuVdCWWUPsH6E/51riH5iafRSK1Q1Vfql0bzwp50
PeoCzGVvtwSPycczcmoMAdVpELcNOksiZs/vbyK0qxZ9afiWEzajaSz7NlnWwAKHvK5klDrLYILS
3kTOn72GuEW/9d2P3gxpHae+kB5LVl1DSvJC9uQm2+mW0Mq7MSJbVqAEOnyBoeVmnVNyDYfduH0m
iHc3yZdAtXYOfpY8vKfU5Q7kV8Fov4ROBFEI6xaVqaANowLKC+DgQlCfizsLbo80TJzYD4mJn8hD
uEflUxFQtlEkQezEnafYgbuA0tdH39scq/1uCYocPuZZ1CLPS8fgQUW6cPKhsN+eQGBk+3HZXoBJ
j2wkS1N3J/HGhrBs+f0jujOs/g+ySYUtoLwnYeosUzVQ3fHolxA06n0UFpfr06qDpAqs3loJpJeo
iksyUP8/zLWWL8vcFfF6DbANZOXzHvOZuGa9IAa2Evg5pJDU4LUptscYTV83zaOAvxCtn03GmvRF
BlrqkgVZ9OfN7jijls9DjQV69doxnie2xvf6AyMXWiT8QTyd0HI/G1+bgBRJmPGwTyTcdYoXqyOa
dgcrqamKfNdyWt3av2fX4tWrS5/WTqkKw94G7bDEbjqIEvlJj/X4SOD2XsX3bVOkSAVUCXlqicc0
BzbqdTlGdQTozekE3h5OdYSa+A5tNgiS6IQcDe/QkbaH7C8WOTgOvPOhUVMald7/G22ZhyGEP1je
Cb79AOdxoH4Yxjw+ym9itM6/ZE4sfF9QsM1cIzKMrG1GwQEY8i94dfXDo7CG3mbslZ8rc6cgRrVQ
aFwsoPqZXqRYp0JcNJHNSU1oKM1zZjf833SppbWGaTAobq8fsObsC4nYDrEHy0py4vWRbS6UCJK5
DDIF7epd4GBE8P2mSUWQHM+35fRppMD1r4FsoGfu7W9MQBKZV+VRgw6wZyjOQmVziOnSwzJ/zhYZ
kuTNH+Femm1NTyKZmD6mN82bNRUKOYAh3R+BI7wSlxP4w487DjQ6Gniu+uG7DGYVJlJCwfdk38Jn
UDG6uY91EBmze1gFrk/b901hC4txi5baGKQ/6wx6i7UlW+agMJTRV2mvAVUGwdWHSy4XFNJmQLN4
7xSsi1m1m5e+2RKjjzzxfCmtRpeawFVUDmWH5LaWX4HgbQDqZzwP2lj9OmGuUPFrcGHwpr5r90Vw
ui13s7mkksoJvMhGBAwkHw1p2SEEYB09Q0b9toQCQ2+1A1XZSceZ5BBOz3sI1Z8NCygFcZM8tR1R
3EV6BJSUPaV7+C714gBKwGKkx+jH507DTx2jHw2o/GlybVSg7BuvCD+RbMD8ImjVtl4C5W94tHeK
6prv4x9Wk2IvlmxNriq/A1GXBcAz0zcryPv7dt2TjQgbWF9O5qLNax5hOkyRcFuOSWWYM+U1kOSs
8kRTSNe4xO2L+mS/N+cHJj9mpLoN89eYoat7MYQ7Mq1wH8mkdeU4ktg1xv6sRivVf9fLYphptXIJ
H3Tf5SpGY60S6S8YMvQeIEoN/v/VrAzwdozUpBpZdJutJE9S47f5eSiPFtwxtrDfmlClbS03pVKh
jU88F5OpqBtMkIENk9czOca0HB56Q/chu9sHvp0V44y3m8uIiQig/wl+r/EgFU9QtZ2f5mEtHKPJ
AldnUewfkz9FDvsUHErU7xcyQ5B9EpP4QhG7oBk7lLs+nv2P2j+4wvSev6o9aXnuGBJUoaOjmlWR
980ZEh3UYXyHTfI6rmYaC5AYOAn24ba0HzECsjphbjfozS99bGY/1VV1KdFEUfJE37GgPpyhZF7x
AXYYvZWZl1YaypNRNPNhNEBC/g+h6126Gs8hEaZvT9R4XmIRo12R+VwKkH9iFdEaCcYTEeP9Rfi1
S++27tpkdawxXhyqKxq+0s+wnnZBgj3sEO9gnIF55UB2NGWa1A9mXfk7lSS9A/zBI8MzY+EWJ07K
n1NzgUEcLs5thZxJiOPftlAmWX+39hEh4abP2vg8Bq/NyTFDJT1DuIIvfmLOHhrxr936+zzdVF+U
zvxQ6gp/Y3jgY/Dfgvnxwsp++AIA+hWBINox/6RfJTTy3soyNuuIiVsvrHWOLKF0gNUW7X9lYNa0
T16WGqy1oNALJNqIqSB+mhbj3YqEoa0MR5nVH7q+TF4kFvG9ONDQPZV90QB73+GNnvA3IRoraHjx
d1WOHbs3bQuMn4PXEt8nJtBLHxL48XxI03RBzX3A/xfvL9uVpdLaq54reyStpvVoK3urA4S687Ay
rz1vtLN2sa98ofshkJ4cUnHX08HSiFJ66N3n5rCf0P3k0ng8uspJOxsCxQrLQvCIFZVvdruIAkrB
U0CZlJdSyK48w9Wf6KvKnwMvsLHePUEhsHka3GeJdfdXIcz8GJ06PQmkwUhw2XeqcF67fN8mz4PA
kn7Cgzot8DHJxsCFDRL1jOxxQ06kuoqjPPv2j/3el1iueafQoYL53Pq4usUOnM5qDVq6dOFGxlaw
iVX/nfZ//cYjN3W0Kz9Qaz2fMVx/5w8Na9V+SUXsBJFxvoZcmcibVvC41rqZhXBaSkKfwhIrGjs/
2gPAuTipg/jMSC0LqqXQdZ6MkbMwkTFkUIGsR2SG1OLRHurhbRdOF6FB3vxVkpe5MTAIq+p7txdW
hha20Iuyp392M9QIQoKkJ34ZHvY+w06yHMUnONp9MyGyrbdsowVWrePtZk0541Mrr7uRqePIXRl4
zkqAE0lSREsla3EDuhvKpUqaM30QUwLODbn4wSv/8A9UoRK+Itt7DcUNx88vr/gvharcDVw4xbUz
was7SlXXdCn+RehbimqLUaEvvRQNwxahgziHoNXzFTJSa1nOQTydX+auYDIyDLNQSPcaROkA44QN
1iEOfyeeWC3AhvGtIEYd8vMq7THAQSz0SweOlLAzZH2WcoDA60KV0RB1JPRFUsMG24xDr+V8uztU
JbPN09IMiAKziHot4Z6G8OBIi8nhgr/+5q3H20XH0TWrdYwQvtRTqel8XuRWJlUFc+/jGuC+sfKV
GkmENvKOwrNLotRkkoHoOSCP4BRjXweKx9k96nJuLz7kdELPKmx1jXhQepSqMGLE3fF2l/RlGoFi
epKtOpX7JV2l0PDmcgCkvIMJLr71AFfzz4/0wMC5kbRA68m8Ahw2TqP/tujYb3qMg7IbeTHm/K0h
1x5bWU0/3f1JjMZEIhPx3MVD+4SOiXjfOrJvn727vFR7H10W17DolqQo7hl4TDz/G8QJKAqTLQXN
ex2hRmmLgFastL52UxMTVupayCcwOz2NMknCLxzTAFTCDOiDA8nlQMvEtoWu+Xc1vpsAlU/lnNL0
X6wixuAP9+ZqRgjkX4o5QtM/atjhp8riucEPzH20LDAGFxUE7zGq2BgKUNKRMLuZDvqQxlUb1MSF
Mwii4DsGQ4QkioiawQntBnR7OFsaRTHfUVQPR405gQToYFq7wsaEbU/xPVse9SKtZW3WGum4s3iY
xGWTL+MltFnFEiKGXUVZhKjNn10O+WfvEWaoQ5MUiZK/i6ZVJ/wOR9fxRLbmSMI7z2R0HtdCxlWA
dTiSJ1NDEmzJzvSk0bOOyuuMKQLBsPjUXYBz9HMnISuPjx6N2l3S+N8RAGEWYBgjpil997B1+RMo
cRgooVG0o9NOV75n7PSbsUeouLkr+8n0YTFdaojJSlYjvW6TomFNbakFC1ABQAGbuRP8330y9wEl
5TEq2+XhK4Y+/wwup5LJPCw24vfrIIfzMfZshuKHURNFczSyMCadlBlsLrZuAehwA7AtZ7QRAEgU
w0YP524VEdJsUc99mj8xbfOhzN+4lE/ZidLaaLJNAjzAKww7IyNXkKQWvkf7hxJsNLCZrP5Z8C3f
9cgYnVdgtoimNxBBWP1Qh5VIICdqzsxFDR1zAG32dY7krU1HhypFG7ksIW1aCo3oQ/10WrhASbtR
Dg+rQ5DqW/t8pczocahxMzozWKW7zECBd22Wi38f4TYV85VxkraXUGRl+oWFC2muCvxrqZZ39Emg
a+1oBFcrNsvWxQBLt+Sn5t6BwK0Ze7UuUuUTO0IYv/+en3e23PdgjgGu8eq10QgONUHjeR3NgVIB
NUEYnN5fPup2/RZICYp+Jjpe8pwiuOMcOJ7MVpfNl+R/iGA9c8PXP7b2AsSEIs4Ph4YN6iRMicac
LXWQHJNzr1Ayp+3YzL7GN5ga7qP+9kVBuCmTzQ5CtW1BkMgeFaPEbT5vi9u6FFI81CfdWYim38lo
LwZdIvIVfgnCu3ShAS3w1jPtXYyZgNoB+u+TytgnrZoKEqvKjNnuSpR+tYZ8Ikot3wSv1HRWcLLd
hrWingNw8RcvCOB113j4lHgLzlfmMmQ5sVqrNvfrD9AjKn+ETe9yntkBZGkB9vBGMMfxdrSP/w+a
RvxndimKrE+HW7rnQ+29iF6Bb0BIwRSGfRGAFnCCkdNRr4kszvLh7y/dtHTRg/qrqnjGKSwwwFDQ
zayALGEPn6lIdwgycYzinBqjKAlPqGKeU6A9uodsP/7dGEull8vdVx5+Y8bh3zQa7drzoIHpsMLO
7HwI0iKAggZ8XmcY2bVbJjfpiEG5QWBq15hPqqP9wmm60A3uS2Qv7RqhcN77m0PMR1+ZMRFdRlTn
3vMegMOGaL7kEst5Uf+kvgINBfInnGX2vL2UySVaNcgx/bLuBhODfDUFYZ0UZf7Clm9VhG3NkmTa
o73MHYeLRyLP5KdX65KHDr+lkrPZ2qAItPsrC5wPjhPNsBmXYdjpSNeoMA2get/qpXUonouPvzVX
lpQyE/bR+ZtosSdZvdQJpEOg9o7SLUQmaSgxcXe2nHyTfXurMEU6YySaz3D8A+7LNJO3Xy1uvA+q
787vpmnD8TEcDP4Q6PDtoG/WNmwkFID76c/Cb8m+rtR9qsAox9wdy8ha9ECamwSP+UAeLoRt3Ek8
mcZTBn25pwGQ9YJ0DdEi4Sr7/i02YvsOOz18QkPlvnNpRupPK3GOk7b5+64mh/2HXcl5vpFBOhfZ
Cujpz4+UN9zLcn0ISkCS1pZaPPhrWNyLRSKkLDKRqFte98X3DYVh/fs0NaHM40n988/McW5ptwAZ
QWNxmoktDexRYeK8yUg/SihZT31PmROCX9VAtOGOjLSgYVt/jmPyu5y4ay14JSy4AJVzCxS6jeOJ
kfMBJEGzIN0YcW6k7vjcJVNPF2TgHX/h18REmmUdKx8pevwSVpSsiS3QwKZQk6DxY1qb/7Ce0MMK
OAVjdheW+LESvnNfqkY+MLp4LxJKmejPgy++QM4wuyXkPLxqn0n6weZApggEpmVsbH8FUT0dfQNe
zt79BQ1dpSkjvD7j/iJK8e2BvKoXlXZHzikAYxwkJ5bsfdFvS+vQAcxm5OhaqI21CZ+RdPr0cK44
ZFFnG2PzLoqWrweXWNDM2odOYU0meKsEnb1irrP4aBueFQVRUGCh/rxbKVbcR/1GtOfpj4vbC6za
Oo8MuGZmDU50zdVCezreUB3V3VFFyfNBOsYGfJfY1WhTGd4wZw5YaTqoGs0mUMTOekXbWH+qbqru
kzinpkrvTA6x4X0Biiy4FBspaG3xYjZm94VH8Qv0NG2QYfUxtheOQZlN6FNGVumgRDqndp9lSHHQ
twffEhb2vPMzZkGA2jEZmwWZlfGu4pSM8UUt1Mx3Rd6b358mZAZt5PP1U35dMOdYvznCCwRi0FYj
MVEVq4ZdB2lCpPOHQzxHP73wZpy85oj0/EDxFjzBhza4RWxDxI/DU2nBS72Nu/EeyaLLV2fj5lhh
h/nxc0g/uIIp7gCYjBnDtdQTHrGccfVFtWDaTIS+CWJ7vJATFL5AyIteF9QM8EbnEjRHK8LPg2sk
NhqJoS1FsGmEWKlXhrTYKh/3/AK4h6/ZX40QulIRBRbf/ANIwLOQQfcTmX4+ZVoIc8jIr4/D6mt8
ZxjaR4fldTg4GwzCI88aY2yM76QjGG+tLIaD5nAWePkK7kxmjWbO5w3U8raM/ubsrbK+M4zbULye
jk/rmlE1wG4gtpOaOMopxaKPaKPI87Zb0cePsiJm9hmHukJREtLL/FEvugFg2f4Rg8wkIr+FWSEJ
e5fnsw+A8CRH6oeqYY3nswGDAuZRAwoQhzFZAUULoyxljS+zSnh8SD8XT3gl7tKrOuGQl90XUv3R
feCAeYBQvGzCyJ1PgMk4SQ5InBb/cmQAyJb64W0FYIA6VSOE8jQteir6d7nbjM++LOOzATkKc2Nh
oKjQBziBJeaO8H3TRjuvayqNZs+nBml4XR0OWuKrVUlpbhGZolnaxF7l9OYbRpYkuMYoFOYg4Hdw
8Qpo0mSa2I2XZpFdh+GUbrSkcms/VFcZpyQUA+VrxDqZ4OWl26dw9e9MTNLZoL5H6eZSbQ0gGU1M
g7inz+aIV4emdEW8CMHHyXKcQKmaj5OsHFhBCf1u1z668+60JtXfHqy5LJj32qIaS33AdNVm5hev
GGlHMenZHg7ZueLS39AwMm6bw+P67jl6UuQJul5jwfSe7WAfU4QOqrc72U7Ah74w87LTReByWaCf
P4rlcpJxFZaDMd+D1RpGRizPf2W+uau7KhPpp/1Gyp+AMKRD7lrLuG+MFVYT8Vye5oHsG/FTtZA3
uZPJbd/sZopjwdDc8kPjpmtRhnRoOdYos0vC9a5aCPmODG6bKCxdt0fCgYt/bQ5jN/J+6oeNOoXu
DAW0NHBhrXCtcVyvo5qexgockqrcmcJXOuKhy1eRh9Kcd863QktHRLatPqAV6A7MJHLPEcQDMd1v
wU26njqGSzsxiyzl/uzTeo8jQ0xKeQ+g/2bolYoo6ugf5nj8sfJz0jW5BfH6hkrVhkZ2QBRjG3Wu
HPxyp2x7KwyFXo5FvCSz9Jb/dCPlWM9YH1ZkFjry6elyPfAu15WGxu0yAHkvhH7pKZwsSD5CYZq6
Ul2O9ewCMOjkPZ9XHTR41mDCozu+LqIGKCOO/X+FnkatX31Wo+exXTglHLpy157CJxdp6KPlMQFM
G6sZatq4qdUhZsLzftFG13Q17wCpxYcR3PIP54QjL0O1+7C+HbTYQdjRKBm7S9HRCnHy62+vtxdQ
5dn3qWG+asw1rq4EkyeqmHvZMn52rklQEQLnSoBt1pJyqOER+5zCxJy/7xIk9yWKlDWH54CHahkQ
/bapVewcwyKbImpvIC0o9EeMXy3JxjCifI/Uw5Sb4J3npCH9YjCCGExOAoh0bWz9EMke+KKuQhsr
bsOAoMwr72UylMjBJ7Sznz6QuGhbrw221y5SzSUr42q3ygwW+SYhPFUjfK/c+7uLa+x1Uv78OOpw
BN/0GJphoCOHFwcxX2ZAHst4+/nMcHpKE++ke+PxQzkbNGVImHDAr+uPXZ1X+bnOdb1djCciHoLe
+WF0pkhMxT9NuZBLRPIHeJVdsOv4gKvzpvP7rDEEUEbKbX8MGjxYArFjJykpVEstt/OwwgMoWHq7
jVrmLsw7BgSISXonJ1W0jOgrgTj3GMSW/u/7s1vhGHU5aaMRkco2CfzVU3IRrTN/LQzuL+cpsuo2
HDOvNaMcCpZd1PHbWnPYSBp6Jw2PNhbxy9+Eu+S+vRzgR3h7pIn+23C13iRsdpPNbZZwMcZ4TeDw
DfqRcOfMRxEcWaL3mDpdvxjQ9f94x8FQeINgkPAIpiaQZvCtwVm+2DRNIap9z64TP7q92PzkoS/j
8e5v2I4a8MPjf7WUaNEB02fj6rKG3P82Iwk8Yfkce7NzyJDQBlDX3Yqd0zp63qwhLM7Hq0/e9i6l
E9Zzt0BDHV3uJZfSoaTvfVX58O2U6BfF9dnLlYpGVfa9KWA0knkRpNNFp1AySrHK0i/RywldZCB2
OfHxBSBhtVEFIEIunkGIi8bos5DvorIixXHTX1N1xWbOgrTERMAJCe6JK5mWOUkVILDS3Kace+ap
fxDzCMH+GNLqURnj7qpDD7sUjqOokrAazOMKC8BSquXjkil+Zc95R8HbuISzbT/Dxe8w8sUlCxBG
aCHl6sC+7OqehMYyFpYkhv9LddlWDAH0H8SX8C9ISA/NoKnfWtwX0weMTRJ51EYW+xHZ6DXe4KZg
nj7MmZUY9vGGIHsoNrsFnbjr2yesht4+qqmDY/E0RdbtNKDEDWVHqoOK1EJa27L3yeHtGennwDoL
XVBaieK47et9/SUtGd4xT8iMbqxeGZZplYVKLz3taso5CyPp97y8xQkR/9tqrLgzg/u3HewEiMiY
Ijw2thY0r0PZxj8PLyVqGpYD5tU+pyQ4auXAZlfwN7BGy1ThUUgyvdxyLpF++CdjS1dJVXTXbpw7
LdiZ88kRtQuvKG0VBuoetF0GSODG6bN2ZiUyOtw4iS1+TRULFFU0+1szMsNmRYbD7RnHl6+bHrzq
n137/hFJuEvPVzvodxvE8bLnQptTcpF4mPbr3Zydyd0897GYYSRor/WSyKTjRpu2U+eY9kBWGyeh
7yZ+1jV0QqDujy5DYop/mlB+dM8wbE6KaEjORLTMVgd742W3CvJybRwZon9o4ecMBPLSYDlRB4Xi
+PsCAcBOXXc7g1lGbdq2f983KwAc43gwRHIQ/4lq6KOPfr8dodrA7jdOl8RR9g3w8YK/D+6C7YHh
v+XPNOONFaytjZ2a29zqnP5VAvP/s8iyp1u/AnSTHK7+LsQMrhqPhEJ3beqVsr5T4BQ4TXi7ExSH
Xq2dShYG1O26eu5SSgBddRZ0Svgtflaggb0JB6EaFXko2qhjKIiRhOVBcazKqcK6ZfwQf3ZGmcHy
3mqXylI4yB0gZd7zebm54SC4fTsRZzcyYX0Nq+slRGFbaqn3Py4mVS8m6VhTg3U6jx5cW5oAxq6z
oQK+zUJ/RQhkaSWpMc4yDwVuINlsFE+/wrJpT6uq+LHka7SESDebRa8iV41xMKDUXZzfLsu4h6uz
EWq9PqfDAh8jkFc3/f6KaYzLFujZyqHMdNoZdJvzpbYYdKoNUm3GDHi7rPczP+zm8vgKoCISsf57
WCIYr3UeOKBw8m2LSmYmZDM34wnWyoMuXXAS6ItH/el/21rtHxlVHym/AH1BRYceOTh2Ow26iM5D
RFWc4eZiySjMwLNzYAL09f3JHJP2h+EX65Qbx7A54FjmKVh2+1zDGz1UGPOPf69cSdCGXd3ZgZ/f
D9eTTaA1XzBn1xmjC5TSpHr1k4ssMmvYz/NKTLF8rGawkqZNA72hQl6DdrvqXmH9dJgPkZqE4CpH
DOPCP0oqG8yuAaMwDIEXMSYV6m18j3KKV/kmT19GwBB7yqAEzCsqj/TfORPRvcvDeBKwbIF0QxwC
rG+W3wc/SS9YRogB/LaG4Zlj0GwxOEcFpQ1ww5HNibrfQhjWvmQGWgmQV586Jxyh9MYE/Ura8r9n
Yb3XsGBMvz0UBeTrzxxKVEPOzCKBwpnrBxWwC6e3b2FdoxOvxLDgxw1a8KaTvMantKSZlhJ7m+xG
R9KDKdrAhKRQYBu2OKxw7k2RNoELoeUb4wz3oyZdYVXG0cIkJ1OXVozibvdu0HB0Lh5sR1pbXVny
rew8dtHZy6RhWDv8uCHMLp0f/nD2r2+btO1ytsfnskKjAy2A8EphreIM71JgkdcfA3VOXCTlFAsK
BZSnxX990x+laGBBI7vSVtoILYWFXZCgxLzYYcuKBrWDK6Yz2tumS3aB2GFmmG/OgzTQ6r4LE7/c
3WxvlbRHTfamBtSVBbzUX4/HwVi5wzvHL+LiJ+FV1AQ1Y+e7tHCbGM/rpjLDTT18N3uA+Q+0FdD5
SxDRkUQRhnDxDNmPTqLKPjHmPKFvof//RcznDrDQH8Xw0Ce6wo0j/mQhFSdftXTI7IAIqzeQsRZh
hStwIxiZOW+SQ+QOy88qIqrzHk66regqHMxNYqlNVuVfZZYR/o6OHrWLX7lUwkizfkKjgT2SE/dY
IcpSNWuSctph99B/L9MgZBQkGkZhZejVCv1NiMkRn51/HKt2WmFBPgxhzj91R2JCBxX2eS3wyTNW
bGwlm0LpzoOsJDQsvhGqA+vsoc/gf+pcJmmlZgy+XhIuhyIwng5fUSR0hjLQ3e2PBNI14vafyUO3
sIxp9j0xUw1chWtF5/S3+s+AWwlFwaAG/lP2P4rCmLVDGm+KALcE3xueSdSX7HWiouov24KUIXFR
+IdtQyCf2XxbZFQu4NusVvwb8B17oxXLYKvUZohfipXbOixIPOL3MAPZGy5WW5FWrFukvpG27bKn
+sIEN00vmjpCmy0iJAWvH4p0PxQJ7cfIQSxDgkEsc8GbUGHduWTZFEGu6TPuIwea/tsgjfsgCbMo
u58ovly2i15kbs0kYZPw6DvBNLFrwYgmyK0L32aLHW9nYqHNmoGRVzBkznIupEvKCwQhejMMaH3S
QcadJwv3lN6EveBGrCtejSa/gsefOHynzv1WYCZbpKQwAO2uAX3oyh+hcmEzfSIHArdVGOZWfreq
RBFfkHHXxQvwrs97eFPeNSQ7qzNYWKPRhUioRFVW9MZdCUAb84ZIjGddehoR5YV00u5ZbcvXIBHL
zw0rFFs8zi+gLbdJ3zVI24FZnYD53vfNTGfwW1Bwl3DyCwq4U7Af7rrkiaLNYMOB8XtI0oX/Tc2l
8kcAwagyVdMhrmOXsFy5Vx62D/4qee71K472gqBnfnTAeqwjw9yRepQ4eOScEI1QkO6cwtaiP372
0dcQ6Cd5CtR0c4doJ8daCdJegkvokVgvvO4J7G2e8ONB57UAjiNuRZxUnF7AhJAR9wdo5eu3UNoX
a2CRJk9w7iuEb7BvJIcakG5yZI5amw+AqNOW7ZPN6IEBtPc7HaOAHi4QeRBWPyXc2hHQ1o+EWALa
Aqjp/ipRilTeVYJa0tq+LzQk8vw7ST0FPwZUrU1J3dYWE6QzTOeO/KloyQhFzSvSFBVMQIIxmSbp
1Q8C5sq1+x2ikiIbnT2MFaP1gnne+R/6w/hleqELnlOEVRzSdIKVFYgi8xlqi/PbqQwjh71DSW0o
S+vEcyhxC5lsqqyxvzBK5zmRCjK22nOd/MafpDEV48BWqGHkAkL20Litui0HpL1cQpC3QRW1lxN3
QGEyLp6H+HeuCPwafIaqz8G8/nmcrtyraJLT8k0wwlUZIQXKrqwQsINuLb/05LQ65lTXZks2ENh+
cOdsDUaOJUHWcnk6yZnpLo7Yw+/FOTngVbqy5w6JviBOGhdsg6hv2T8wC3TWHngXGGUMot0RbILy
QEsN3NVjnBZ5dTBFe0QbMzeyghWKByyxU32SNPppXYovJHwVfy0xD2MzsjERR/w/VgQs1/EHqPhl
OhHRMMVj7sg542q0QG2ysnrg4AJUv3CtTnQUJau/ujyffNjU0dS7138MPJ9MfDXVLNlelLcKY0MP
mmq/BCYrgmJmgsJIh7aIH94KW32lr3JQDRY1RT3KtlNd9LwuUJuOfrIcPB4ZPXefaLFG7No5fTUy
CGVflFLXlIaFbaz4tDc6qiDUpAylgbcvRRrovrM5ftifcdxAVpuV2u/goAq0lSZBTHnsGEmppDGR
Src2X8kpXov+RCNmryQZZ6sgLtwOq+X7QoE3cz5oWfi0ZvFMdXTZWyn0phJzYdtHP3mxiigHIH4+
AVkwM1ANoP9cfRujopwt01uSioqC79KjuCTXnnc1027vRn7J4MfQZycfI/v8Fg4f2eTHJRxZGA4L
DNnFSAoFJVE1jszNIJwbmKxORRR/WAAoI5R0tjexI2j0f2O7wteABalH2/0KuE1faAMiLqgrvwmo
hLQ7TgWCGJzvfDhCZxx64pU4VI3IrS8URVauWR2HNxdpYi2Lm9IprUz2Fe4qzgOkTDRmoyD6ERTC
73GNbGPqv5FPeqAdTWfE1030KFVGyqm5Jdnr3PpaRvE57A7xB7XmSsAZYhI/vKxmkYAM4F4wSoTq
MEBrq8VEy1hok1S/UTp3bsNeMtTGL0ebmcdNB37XJHNYvr2wecWTXj+S2NEYYq5tkny45+FJAXub
KhfWkNzvnVymGWX2aoLVshZryTx2aAzQUIoeydsFcQME8usQvkG4ZMlr/Sv/F3k301EsXRc1hMG2
TZxd3jKX1wD6Vbpqfz1FV9oU0cxMyIK/DeYKpO1/7CTVhVU4n2dwc3emijr3X3cMn82o4dwrmqzV
tlUqAenxxcbn58tMT3yNzEs4rT7hCoobtjxixN3JRVUjoRJRrKF2sZExkO1itqqRFekmJ1HQdtWA
njcVZRIAtUMxR0iq4FNRwO9ux2XXOMbDBOGyIkpwVAA/P5q2xds7tOAzaEafdyKxtxmBntjdkEfO
px5fZSagzzzkc0UOQGf64zPKK7wQZvmxsgO+L0NcI/VBr11C3CZH3Gp4bszGWTJnzJxccEmbsSRa
YkBtLq/mv+CE46or7knndcPFNrWmIH+ncsM2u1Mmk12gcobAAdsuc4iGAy6walJcYOLco2QQL3vY
GqfhyN10gOiKPF5ubKskcJmomINrmhD5a9ZWf+gSIkGo5C2qpzasI27T0yz9PZXHT6cUFb90rkSH
qvClvryl/oyCIezx27BFIC3WERphl41MuM0rPXbCnMfh6jta2YjqzjcoVOgcKKeBV3fsDxuCenj0
xANqwDT2/BkA6MsVwa4YRBRI/HwyK9WsOIQxDMW6UOamQ2RYmBqekcp9jyR0Ks6krrCvTcxK/YiV
YMhMtXSddhhP15yhOvbWnl0zTcbjpof31/SzGmIRfSQj6pNAt79CPhxNL5r+ZHqQwom58iBarYvj
ezxQSlbnrdmfD9CGEtpamb8HxjwJAuUCtsec5MVmLljGbJeSzltBJAPygMkF0eF3PAeHmRvIt3G+
BM8K1eOikYc3TKJhtwis+xGJqUJClDq3iPoBV8yNkLNm2Ifen3unmZwhR2+LW6QDxA5gYl16b6Qu
OhhOylMO3lQfrScHmMLnzn3XuLJYCr4gAtXhT6REKcpe83NMD5cDjiEm3jLYPdpoOkLfMSci9D6r
b9nXWB0GeIXx57QjZManItO1Lo+B/DmKGNNEck/giH3lDyZyN+Pnlwo5P77O0z09DQwQONbqAR9C
y0v0B13pbbNK0S6jHIgafQmm69ykmm2ZkzgxabCFp+ADB4JDptx5/WF+hyv1v4KC9szfd8rWxHHt
jNpWlXGP4BcGzlSIlBUUuLQ8CJcnkwCyCt1WSmjznXrE0BJfA2L9xYcGSpuVHparuDc/JMOSnlak
yxQOIIXtn5baUhmrBN+JtNTnrfHipY4Gxeiu7Xt/E9WfhwQPSf6EARc2rmOCLz0R0MBDRTkOq5OT
QAueHMZlfxqOT+rrVGQznUkEhT1gd5PbA6e1DKdjQXwWWrMg18l3COUNK5XsFIMKx0Vu3ha1QfB0
+yPGE/rXIbR/OnxHoXBJBzX7JSUvDAgn/cnXcPSQsOk/r7fNwDHOVuDPCR4spUmzfmzbneF4AVyN
z9kpcDL1tv5Y2EcrMonlnWAvphKz9+fYqVzUgf5JaEUDkF/l+e2lN+FN2pZCkedEf5Xi8FfdnSts
Z4+7ATGau2b73lTa1vSrBzICVR5b08QZmerRPf0fGAObkL+7GWKqWQrnOGS8mw4bbWVEf89CGJ4D
wudqm7fELvmj2H1qGF2rEitTARgX2w/H3IPplYORayFcIWp05syU8xud35JA1uYTMHMJKFSGx7h8
WvyvUqSokUs5DDyRhaCxkEjQJwK4U3aGqJJD5fr4eEKqmQ7jxcm8kxKtpbmckDn/FRuBCgMb78Ev
1TvqkfjFrQ6wjfghDDQOFPMNvOVwhlI4PRFjw+MnITB1SO4CCDew6iArznfQt7PscZMlE7NF85SG
AxS/qXq0RJ0RP3e5tL/kdWXkMHC8fOJH5xkOg7eyKVnIg5bdH1ObdhltZWEjCW47ID/AX2Bm15/1
WmRq/JN27v+Rz5XMtJ7sZ6ALqP3q76jaggo/zeCLj7O5amI21RyPAOsPmWTmEsHgyxJbXts60mgs
lRrsSJVouyXAtpwtxsIrQxkIDQ3Fw4FZbiHCGErr/FYneWttNw4ycVhpP+y6RXrorr2cY3fPAXf2
+mI8AvxnkpTiplRixt547knJJ7ChJ8N3Fk3IPG+7KKjWYyHexxmQPvP/E4953r4agW8EKbQMP2Rm
8k0EJWgZHGQAu94XDXLcirrQN3YlAbObsCy/s7yEv8T/WMsZWoaPegwPITnV3GvRmJJpsTksHDYE
sVg83aooofHSit1wKmAFdL2wcIaiDHKNaUWDCRgd2AxgG1sgTvdVvlZ62ODTbqBxUhJdYdAlKgbV
SPzrRiEBvGkam36A6tQjgDjKBFuK6uMm6UK8dCiFYj9uaqDFoBMSFT0g8ByssSkLJ7vMYdsHctIu
E5FMnxVSEDyLLtpKlmSQtruPRnxQMerLZvwbAio7GILhMUWXHzspFxR/kfSXx/4sa5iToTpNseQ3
1uJWjztTm/9RqW9mGsGVcFImd3JBB0UiXErAuJdLfy+ucna/YsypVZxc5p0EwNwqsF8W/vdBzdIL
DeEmWVdNJuzMa2y2Yh8b7/CXVekMXLQTbpgLSEUzVux+atIddMHMlf7JGFtjFhULydETINkUuZkQ
f06qU2IQVHJquJ4BdLKjuhncHKT49+g/hH841tYdHhbLgpA0yXbToAJqWdu0PXShSpXc06AP/VtC
EgsDXrwUoPfk3GXmneEuCkxDgo5Fa/pyO5E26vG+nPz9C1DbggEAbodeXf2jtTv/Z8oh+yl9UdyY
WC8K2E0Gc76BF1xkQi6axX5z4fzQeL8B4fT0EcaCnrklEz9XjRImWMUhoPCOW5YtdQfELIAe4U7i
S7g8aXOGTTSYb3KYq/zSlh5Hc7TVQbOcK7pcu0RHAOO9XTBj+cxzfl2wu74m+8XS2Auux9m+BY6y
U6PccNITapfnEu97UFHmwF2k+ZXXrnBr/C0P71yMAyzUC1Aa/czqZnvdkcBBDNSnafgRSEm3MEAP
G3FweWWdtU0nX7G+mcA6sDUQNVCxPcOZ2/x79gi/PKIu6nKnMr1tgqTsThVsmR/Ncmc6kGLlnWxh
ZpIdMCLHpOM8suPF8s59d1coF7AaUY400XW3ZPC7RVx6gH6LHBQc0npMGUQc7dAcX+d/l3mWyky5
gMgz/WJaJJ27b1Zd1OBgz8nh2AcIA5DgEJV960DvRwuhLATqCMnD9nFmpIHkhMDwajNUlsZ+eWTv
lmTRQRwha5QBCnusx2hcSG4gw+K+T5+nga4LGeaStaae1YESGf/onxbEuFJk9Bp3T7X6U4h65Rcb
oyAKw1CFQv/VJsUUlsfuoqd27e1vHa37SprD+bCdeC8IJM7Fadcegl8eusyNDWj56teuXn2j2I7C
MjNkKQseLi/5itbuWK38xLlxSJorgE6ARsnn3eSdbTbcI33Qjy1raQZtwFvWWxiAi8Bf7E7aeTgv
H/Wiq/KEl5KoN6SjHmEEw0T8OPhFls6Bg/r2klD4NO2Mwuo1qFIo0ocylhnvb1O3O/mbuLSmYL2N
l9yvjZxkBG9fh2K1HW30p6BSvVwTCZeO+37UlRdPS0Hqlxl1j2lvu+J+IRaDJD+k1qbpZjjvZbQg
mYxnrdFNc34fZtHwi3+SgYnq7dxzt0InSheOWI02iE+Of16Ucbzp9+Zqg/A/7A1fCg81s0CLGTuP
9GxhGLVg9OQm8OSXtGyIXTNNoFz0aNZ8YGO2/g13djJGb0A76dia5DCjzFqxMjEmWIJe+37fNOy4
KaLuhofXw1/H4CJD9BNPhtG+YaGCMqvRQAII47EbB7TKFgF7OW6arTp2dH9xwzYia7KgKRGw1jWJ
Y//emIFfFSr1W1tMMyi6myZ2wDkjCbt3zbIv+1iiGOXkaUuJ34jG2LifQ57SjaiK/8iBVat9h5Wj
J3Ve0St2DoW253IojE7duXvroYEskKe6tQF1U+Ievg0EReuUS5oRywihXmMwkRCKyD2Pz4oe9MnS
byABjKO7Dn39V8vxI4FvWR8nAJcOuTNFzMvofAQ3cdBX6Lr2jwJxVbr75NfgVFilCFC+S60xoVAh
jjSeai0Db7NGwYQSIbwrHq+Ivx7KAJuIsg1SyEKTMtEbTpRaQpintME3H+xPwhliIe5D3iqHPDeK
T5hGpaFHxJqk3zceA7lHVvYje6uwYVnCkvb5XiCnu1GT9pU/IV/MBpvyH17WVgEG/zZ0P0TL7Ito
M99MT6r3RSEcbt4gsStKXkW8A0xoopqB2FfAe/d4wA1Rb9N40r2TYS+R/5iqKtLwPdWF/39JLjrj
5bt9hcvciS1lHVSw2na3w77+buEQknom5SbhZE0nAWhffFyjO3ygk3+6ie5RHJRdypbGY3gL2dxS
IKPmtWPw9VPAqX0y8L1lmUpCu95ewfy1rv3Ahuu4GwZklLtSHiWbLXO62AErkhtFtauEb51tPs7n
3NbRK1BuB8y1vLntIEuok6ueEYORTVFaPwrcJssClsiX0g2KKJV1LKr6TQ3pGZlqHg1HSZyKnRzN
MerkXjnbCEjh7fqDFCtBAKQW4oWQOD5kK245p7sccxllEcMEOOS4kizIav1sJSBA+jFjtmuGnZSZ
ASbeqFGvfmqpxDD+J4+cCrO18w7WNUtm4lLXN9mcKPYKaPRzsqCbL5N5KYslRzPr4r/Xo4XYgsok
lYPfsBineD9jtCZc0zAERqe+loxv0AIzFupr2JIIjak2PNulmNUMIku3H21GPmbpiimGXUzXwG1N
BjGZYYDnGnXbf+KmHYwBzkEqrksVHwYodCJ8Y4ozOKy7/BPt45HGABT8Fh6JxfUO725pDWQXHDU6
wgYSyWW96U753zjSK+9/7G2eUtn1alQw79qEmQKUO9bDwe3c/26DNK0zYAE0z0nwZadX0dr/aqjk
PskIwi6ApRYw17bFCf2a1PBV9PlqjRUZv3ayzzFtnrOmRoLp4LL+yTdTm7dhl5QUPJzjWHf+efNT
U4tItLkRWUgQLD2wujmQEPJZaov+YIw2qGHYkV67cxTc+aGAyMO//pvDmORCfJQ3DIlAAz8fqxhg
x7uf9lbZG2k0qAdfGGN9kA+etV6ZG/r3PFRuM3Dcw/EL+lLhr4gotzNCSKyg1n9m0p9I3VJosFIR
gHCfV2QlubM5JbFgADUJ8rNBwqkOAGxgWYuoma6LkRuv2EZ12Lp9qj1pxxxpXaAJ85I8PPZ1yjA6
hol97N+sfIyoadFUH7EgY07YFJvjDEhRIbxPVdoOAx9FuwRuv14iGaJCUr1TxSAvCizev3L9sakD
7aAY+MjOBiLnCkEnpHc80D31nuAOku0Kgi/n9u0cKdSXJeq+A+KyYM56/3zErG42wtO6PU+AnRSh
t3OsK+EstCLwY9ZfCjenxWHmF9sOCTanGIPLXj/rOMt0T2fGfej7e1uKNQ2+DkDngS9kmciQMdUr
dLtGXwmWFEJCLENvVm4lDaur6m+wOZ9Ma602aihsBj3iTW6Cp6DWvTaf+XZ+pIe6Uu3jw93WrBdW
Y1s+ZiCvI3L+x/zdO00iSIFjSbVLRigm7CWsUHWjYkwprtOsG/ZxdC49CeKMPXq8p8mQA6Gy6O2P
cmOT/BVsWyJ/mXCIv7ZLt7GKfVnC8W3Kvw1DXkiyU9Osg8JpgcJwM3oXKHWQQRP/NJ/0I5cWc1GR
bD2tWdOz6kj4KvhDXFFNbl+28PWgmkg///0ApI3PnaNP1tVIts0nUFTXDzqSKVIl3YahQKsLRieB
DG4ex1pbLcON+TRYoNYUBssoN60SYAtTIsdzkBd7/7LLvaB6mBK5nxYuqQnIVHfL82dm/Jg8ODjp
1Ou702FL70jw0lrna1wy4wprlY/lmTtjaA//pvZ1yTy7etBhM34bPla8jEcZgZAEkAV6vufsvMcP
u8VmwfeUr05kPfEtIpuy9npm9Xo4LE7ms1GFSfHaKkryXsRtlWpLnqpM/4oPUhcbOa7G8dqwaq+j
22vuCqoBDV+vuz4JB0f9BIdWqESUp6uw86jZPgUFFYG9Yili3/tQTnvYeUzWQCvQ6kKTdPO6uIZN
QMKkI/DQkgMfJS3bMNOxkW2AUiiSEiX1THCrv9zYJ6tEn4CGj7cwwosXHlcGzEdYZK4KdgeXDng1
yv1YiD+VWRf+i3cQS5o/N6hpsJxK5i+l4d0Mzh6bKdxq7kyCYIZVTw3oFEFnHjegxu9XmHrfzcT4
d21e9cu1GZb2ygOeNxMPEcMQb4/guAhBr2adFJ9ug/DpTC/9Cu53U5aKf8pVmrgiuKYeheMO6DfP
UpvXoORQtObLED3VUqX6kiD8IxrLeTBNzr4xi7NBodtPF2luqiDJNLx4TIeGC8gnps5ZCE7XxLt3
cCcmgh9MZYcODwtt9gDidf0td7P+yQALPZ0nHJhnYh+JvYn/CjvDSQlSkNlo2gycuWkIiyi1b8YY
4SZd/Qi7hIwu8yW6DfluZaAqsSHFRvAvpHRRItC0tyjBxfY2mqJOK49IoNaoU+p03x2urgGtOVSm
DKWj1DJJ0Cqeaw1aOMQvc55OQjD6g83Vp1DOKJ+c1j25hsaAKURh+s8ZEIA1wiA3v2GXrabETbwd
AN9TKuJfua6TW0nL9luTSK20ckzBe5UQB5Phcy+FUa0D4dXFLIFdQ11XaZgGtfOYKv7RGYsOaOxV
a1EAdVtXNDavdHUXHsVjmD/VF2JX/3hspw8sj9pe2aZeEQJSxAxs00RI6lP8jkS4h6LhbeQkVgZU
Y4Fgl4ndP7Rn69lBHvTb+UW6APV/Q6mWo0gGy5iPu/ljYGtHZoscjbYkNDzXtWwl0oRFMkCKheGp
/3eCSQgM+3ibs1U5SiEgZUEwcOSYUhDqbTS8CRi5O/TuL6FXnBjnPt6nOsGNgXaKja7NAjbBiP+K
GBFneKgjIuR2HisLPpoIQoXw5dCu5z2MLpSkBmB9gEHAQeUcYITGqLlewnYwQ7aVrhAvrXEVAGbt
vphrRJbXrD2/LCioGhw7KwET0wxY6wmuUOZKS3qoqWNPZd6oq85yp2M32LessM//X5rfyKaTkicE
z5aM+yd6Kz5Nc8Xyu/+3IZ0KDQrRlp+93AGHFAzbuhSlwwexG5yBrNjmpqTZJrP/qYOfx/+g0Esp
E4vpuCopFdpCmGG1Tu0OI8yRL3IKGdkJxfeFs+8/o8YpewwRYheIJ46oCDdvKhw0ylquMketLDny
RjqbXGrcB6LMZUw7/0yAL8Ah1cVG3ufBa3TtO9WJ8uIV5buVd7K/o3/mtfDSY7HeaUlUAG2iXSyj
49XMvzd3OuBjYTPFfKpamip0Py16dBc/sdRlSD034bC+RMHQG0Azy6JLBxGBfdjMus8fehdcnhJI
itXJlHWwkGtr4ntkRr1vzRdJ04MbwHa12j77xhbqNzTm7Y5Uvk1aYpERFqFjvNBr8/2EsjXQO3ke
ZpeMr/2T6xK1rGTToqi3JFhbKqWz+9ypZ5a07GiHb2lXxcdikbd64+/EBjlimrDZNyPfo/6eQ0HL
XELhN4SVjQWTJwsppJhgJPGzHvzScUGvPxJUWBQOz4VlahSwWOZP0TsQaGPJYlyGU2Zx4yfOzuc8
hkz2MSOm4L6X1PKXj+8H5PKwCave8CzZRDr8kpjRXMdelKsfiBd1OhaDDQ2ZtCjh63BBnEo6ZVdv
7BIT3QmLr7ufE7w6dzDT1HDH36JO7wmgNI4mJNUmnXpekYVL+tCwzuhG/bXAqJGC5Q+qfH+/tKXi
YQ1gNuB7HrI1QYA1r9GkJeda/iHsVuntnOj3v1T7gc2XRm+TR5WaD3h3JIjEYyp+wPdxTVm0rU7n
LeK5/ulGb/NNRwTZbIlsUkTainguxwK7F5OmDM+gxWKF1xXAMqKBIYiHVwLTUWUP1aRSR4fryVOG
7PnHUjXPi0lP1+XsvqLNMF2KZnadB/GM380abALD1TZW7+i7tEIB376PCPcuPFj0LqiNX7mHARDS
JKZ/MbR5MIHWdaEhONGztxBFj2oq/yQbHeMu4w+F7eza+bISAjvP2kdXsIu7Z80FOxsIKML7RbGY
NUja0ojqDd9UsEoqkfWJmJdVvHJVD7+Oi+JL4xNn5nOI7prKIZdZcsugwTpr7Xg/NCSZq0UXTH8k
BCEsqwzp9Bv/TclWrcmM7mrwUsW2CCbXFXvbet9a39O4AYHLSiym8ZMzKMRR7ctHqa5WERYWhkuj
tCO6yFeelHeiTJOYnQZM7dRXUvfVaNXPRcbNaYcKaTqz2PpR5djyDTvriqC8kr6SkGF5KHtT8JsY
uvQD+wZAkJZN1qJKTRjdxWwfiX5PoNTkfc1zD3JyP4DUjiHX4ZZ58h6XbyqR+Qti8RsCXuFuVAhv
BQh0acqVMhKFKcxkGwZ88seYYJ67I/mGS6UKWWIaGEN9y/xqOBNdBBcgLcvyoLqXVuTQSOjcJW74
/O9fKRy/sUXmWZd2NAK2jIu6MlhZAyeNo7bQf2TrzqEuZU9pIFth3WR8zO93a4CdIeTR5X9LnFQe
GNspPPvJDWGjfH+I+GnNL+oJYT1ByXWzNZg1qQGfvowaX1OKyCqzf8N2/QCBaRp6VmFhkKhHLDQ0
/FODi4BPW5xqhS3VKJy1zUiG0XA0MfrAsfRwzSMF7p3fI7nNOyhxrC8C3VDapwzCc9oYLS13GDJr
XlPg53krr0DpERnNwCg/lVx7CRumiH5vw9gfPN8OmiroU6AZkCtwsXYLnndWoNh4G8vSIMGQ8aJv
mqsZKSVjbUlhseM5TQFIXoKfqQqdcUgoi+TWQKWkjxaZ0+J5rOXhxBTexXStNHmuA+4up3ieGofn
piYr+vz1pgpbdoknALltWxCY+CbQCCjZ7g9TwtS6O9qkWne4V9DqeoukEXF8CWEQ3L6N3S4iozE5
Lgl3CaidIwUbRahO0HzkQuwnspy98YbZQ8+B/rYTmqyTqyoCfx4F1kgNLLijMPx96TQCMKj6J8nd
1WDUg3QTTeIKxqHlNhqFE/JLIt6oZlhicaH88Fj6gV/3/E2+sMDiHSuBR+TRzUAEuKCqBHco60ms
Udb0NdP8Ry9MF0+OdsFtWqkesT2end5lN47k6AUS/CI9aAstIU/UbnJ6zgkyOcS6O5LJggnEMNOV
fbmiYFnQG94esAap1iy6QKZuXc9qnlCRYmwNc5CLzumcI+gIBqEBhCjh6FiOGi3UVjPZxAkiNslp
0AsIfYNvpYNqgcxy3sq6vgwv+MWibR/Pt0wIxCWefMOAfPv107ok4XhLUH4E8QE7qfoWoN/toHqo
zYmruCCdChMtKZdoClHYXOMhOeciJWqtKh9DPw7e75tafiBxQZWOJaqAyEaR5NLN39XyPxTs9osY
8tfIg4W/EVnuvEpaihhNvmkFrQtByYU+1Mph4hHY1O8BdO/Cu3GgW6WwZF52HyC5JN8uhe0jrFa6
PEvhQlyatNTBNf6vI7+khWQfFU2SumuAYOdvru4TFZWMNselSIPENCzTYPObxTqvTEfH6BJjIuuV
bcBUV+fgzXFLsDVJhFBFlUbIyByJFmgD7UXMQm2AhJRSYBk6WAtLDi65qHX9RQ0av6dL4Shdrq1s
7bVJ8BDGJlSMloix6fSoW4c8fbaDNPTcUoF1jm3mp1LXXu5ZPaEvw6k37PV2q2saek6wgjNyVgh3
iqZmecgKMeQsTDGSRaxBHi2VfpPI9vvrWmk0q1YbUovn/GEun1IU01Go9AzsD6bxhwp054IYZx9M
enaGpZZH8jRhKV8fygxvx3nZCGQJUQU8GjvG0YUirq1yixytrFwuKoDdcpyd3uZoAy7AWVT9Xp7i
+lLbjOe4FRPrdrxn9iqQfuwJqwUh/sLTjUB1z9uqLFix83UIsafItcGACAXBcMqYv4CopSfqdzdf
TGH3O66GTyY8qhSEMx7PdIlaqs2GI8RrjQ8mhX5YyuYy1AHZ/BY7ZBxf/aQumO/fU5XGDe/N098n
ucMfRRVKmSMaLuaNOYycVKh3sK0XtRiRyUDDDF65hATrk/4OkP65qlQhdL8/lausY99DisxYZfNX
aJWbos4e/N6kkBot5QCMZlqxQTghoMFElbQnKmetrCTDc/fFKkMQl/lwiuI/LlDq0e027uFBWvLQ
8d3cjIZoD3hMtVtrOassnIfkaVguZDXVq33169DNxDzJGMc4aSex9swg72l7c4IHg4hTNsLNZwO4
Qixek606G68wTOHGAtLspA+xpYmxexMCQGedotowb+hpfrv+mvhbYS/IKCPUKiHaeisL9ehJrqAi
80mKYdIIW1XV7n6utcjKa+QhgfKLTVYeRwMbeJ07E2tcRbx3oYS+7fv6de4+13HQg42E1PEZ6DIL
KqSt2D4DBB+FWYc/uYIQU3ujU9HOs4DmMY9NQQ+73TsjWKP1LaZQ5fNO3vmTm6Q5oBna3JOb3aVK
6QhTDEWpsVcN6xx+uYTqzK1ERdiX84iGohsfKScS4Q10qBkCP9uoMHhmiOzvkkOEO0RtBOPFFePB
r31VS51/sBHVADkY/GGzlVL1KBF3NY1UD1/yKw5/FiniJmGLkQ10UPLoE7IhPr5oOEFgWJF39jjh
+2EZaKsmbaFa5FM9EE+ZbwLKbIBCXeOR3Wk+BT0Vc6GoDR3CH66suOVyKHucsOJNklJzTSTPXO+3
zh5w7xxOtPP6c2aRJs4ZSbQVJcbfoKr5Lor7/gmdpw5aQIPRdV9G7gkAfpJtChq4ovCqJcqeUBgU
DV2YTX7CkQ44QNTxbUoPf6OUHUdMZMQ/jldrIZmAB27/r06pcSPBVjh2eQ5WhRV9WrQTBgGzi4OV
dIRiyPkI+Hclx+Q5kxK0cULiEdy+4Zo5qA367PEKH2LvqhvpEep45cjg3MAHv3EUW72dEV1M61rH
MypsOBe7XQzY2x4W/XT8klS7uSM1SSNTqM3l3RDEFBKsfGLLHXBzf6Bg9W9N6VwmmmJErTkDYG8o
lPix4KcK0fllBp+23UafEHRb+n1aNjXjHpnyTWD/jsxQEJF1y7B4Mea7mrq3c9/60ksodxAuItqI
4ZhvNKCs7SEpbqm8GKqhzsRAmTqyCW4yT1ObgOAnM1UF0pGxXelBrGl2iZKpFcV0zgUHllAvzFbT
4pzwE8f1WHmjADTUxuTzCS0iMMbddcaVvE/ZVaEny1efhvJQB1fkKh0sRapG6kUvpedFCV906IOw
KRr4uyBpLx7VoOgcTkYjcjol46PBvmWADz8vZjAxTBQJsptQVxlyXW6wVY4YUjUjETwFPSL1MxYL
6/kf1YUx/1fnqVxtUK0v5v9J6q1bNQf49NQZrwl3+AHPNTpFo2JIVz7ePDvXINMfv8gmDNdO26H8
Xi+xFZXF/G4aSMPz6YtAy+QSVXs6mUmJ2sU2gfLyUW4eG1ypWVJqIVMujpEeoX9XK5b945Kp2wdI
K5pT+7DobacB5kuFKZEnjmpXIfZGiYibeAhixDoI6yy+VHKeAbwXf5HKqs3Pnn0lhrmIm4oWwcoe
c32CxQ6PNkKi9L6967kIp6hCzAiX0eM0Kek/ZdT1ClqKjjsuDOvLaZjStEp4bIm64fpYja0qg6dj
HVuYBRB1S/l5+AXUQSdpfExhhVa+y/opgRYlP3bsYaZb329ucv90V08jPieKs7e4YjchX3Vd+CoB
W5aDn99bvG0ggUeNJPrVq5KPzxxmkSihJXSVXIyf2YPR3KQJrvX25HaAJrHg/cfaCbH1COYavI96
9fAbfvoEy6sQ18H9IzCkeceWPT78z8krxkMwCwRaOsZsFLwj0wV569l2by0a0aFLapHgcjzlcRaY
rXs4yh18EhbQY2U7vKZJ5PuYLxhxTQKBppDJYK34ILKIKUK4w5uV9sb5rmoU4SE5plAVeZ3kMdiS
kC+HbhCs4MOIubAUiEl+qXRQ+P0raGgdhnZR++pXb0bIWjcQDRll+RHkVCgNPaaz7GpW93SGEopD
lS69NebbfkcwTSZBJN0Lc501oKU1kuN3Y3dUUXawAX7i5+KwMF4ZwlSx8mybbUzlmn5lTdgokcnl
MpBXbPlEWUHq5eJ7cT+PS2oPpiunSDWvNz42cd6Q68hn2naOa+cjxD9cX+DQqX91B5LwBKJtj6RN
0/QldTKsfn5LAMKbsEWL51diaA3jfTLqWnZwaEhK1Y0G6qhNp48A2dXCY8jcTGxUu87DpipXHDly
3TjOA0tA1WTIerZ00bzMzinF/Rwy3bZqHJhx8FcvVmV/HUWXXb8Wqkn3ktziwOlDauZQdM6mAtRB
HrAMoTl6oMyAI1oNsXMRrhhr4XbQida1sdHq5Ug8vg2i0SkLO+NeF9Huy8Q9QM8fn20AbPuMEEsT
6RlxyX/pySHogwCDBSY3FrTK302juXxe1N81FMG25D5u+Vj97sQec1AlOmMT5ND7cCneVC55tiT+
s23ABCtvJVRz+N83RTHkZWx/lJEl1gY1UjTxzn34BDRGZJMLTzNsLqJjy3eogz3R0w2lalhxj3aE
yw5vn1WZAecpPH9pyGDxr82eEXbWfYXtDdcMcQ+J3YxCZ+b2De1AqkwF07stYVptL0xB3JlCuQb+
IilqeE8FHVJ7NeICfwwK2imWlRTYB5aQ00tiwcjrchjBv5o7PX2suXj73oxinCtLqf4/z3LwcO5E
KdKOa/JzPxuYlkMWRxjd8zuJkEkNtJmEGpG1gI/OAwfJ/n4t6eFJU7Ns7P4pRq2pt34OlKAFwLFZ
xsyR6roulnP8xt6Xn7+W6YETtn4TV0D1FbRZ35tXHZQIorru5E3NK2VNIr56maK55qHLiUIUgjwe
htDJDrbbTZ9rJbl1ggDGAyp6qz5G6lVfsKgCNbigBKqvhM/7tLQBL0s1FBv9qonWNaZZnj0MLk82
zcDH+MW1iYIj3lvggI555ydMnk8+tgj+fwlb7zAwBkbe52OaFFti3lO/joH4YXSKLHhBKnPfNgOd
LChY5DfwOxXNAywbW8GvJ7JsXz1u29KZVVLsrTrpWZ3FaXfeWZngCvymwE9zQhslqZuLuQCgWZD+
1SW93fspuIBEq1YqP2VsgGlD23no3IdR6QxLtB4mqOdGwzm3nGdChto4uDgejZFyT6bM0sNCwxII
T3n2/I/P5iZYVKpDe1ZAxjidr55qmUuhw95SQb2oXr3COq2YmlZ5hbfgDYdhEnkROOxMwza0GdWl
UXnYNha+2zDFRgpmk7PBhr23FN+/CF+iH/ynxz+e2fx8PHNRcaO7M+pOYE67TXuuyBfBEVLEYYA+
lvmNdHdHzGty9m1vmS2yYgc556sC/1G51PpV6xkPzILGU+nPpRTZNtPqm2YxVrS0nuM78EyBKwRX
l1j3+phbjrap6End+e6rAsToUkG79cssoIjzA7tppyiLUGz1rAxSaZQckULLhsL4mPM2HqbzHXVh
rHswmzapU+o0H0hY8D32s0ubx4cFBWoLUiEpfpqnoZiESpeJ53ctV9cezX9T8rqY8GJZbyltm41L
C0a+34X9UFmTzOofzErK7EZ4r9hejUzaOQrtnW9urQnUfeqXjCTeZlZPhbb0635EFwz6XhB8Lt2F
cCqCcC9nXiFsuhtwz8pkmju9Rh/guRdaegzy0tB3eAZt2ggorbtrSIQh4816CDXLhi/gPCjbP0pY
Ocahkrq1MgpRd36MlgfQ1+iJcUuoJMql5uD+CNKFNnn33pJzd46J3TyuYla2Sr/NTua6Gac2jC9o
NjmjyEDUxBr6kVqAldxedvDS8EInMUzkXuYbUm2TJBQBjDQAdA0i0fKcyeoICecRN4+thMBweItd
VU1e6v00Hc3SXGQp5CMW2WFpwkKFbpoOmKD27ejL9hKJ9yvzLnmo/Bjzweh0u57GJXqP1NaKJl0Y
eOMc3yV8SE8Qy0EsZvls7N8Pf7D6R9UMK5xuTzBprl1vhFzJuRjFNH0OJ8+ze296S4v7WQCjtTJf
FmtrpKwh3FvXSuPVjswCu3C4nC45+8NURcxE/t3fkC+QHfz50VQ9djBWYCuX7AGT0NHYBrPWIY/0
xzxV+W+nl7v3o3GLn+73a7iRTrAgKns+Fm47RHxZxbjjPN4ORwLd4tYo8DtnXnM7Sqwvy+gyfDbd
CNmMMfNdELQP0dMnZecSeHYdSsHSM+O/8Y3ZUwpY41nkBV0u58gSiZ1K49+IYtMcbtJjLYVcvIVG
nmSzxmj380bUiLpRcgaD7ddgcZML+PIYU/Gu5R27Gu8vtktDYxL4VqGKYO++imYAC3LPnPrmmdKU
Y+qnvoLGthJROBLHPS9PZzuEobMXFQBcvvPBYBIiztXSE3se4DUd/mkQciZVenRLRmHnYixVwwYO
M+F0IqLB/u3kiqjs06i+PjtLL0wIsRAg82eXxOzFWaIwslxywnLGj+MdYVgqVtDFr2f2rDcM6sCp
yFXd27p10Ed5OWBq/qUdUqXwPm9NL9TsK2c2t+IFh7kcHR9tC+dfr9+hlARxaoiDw9odoecW0TNn
r55XkcEYgqNzahVTuHIo0jLtTsJismunWAE2gafPJJSQjGgWlQPekEyAul6+kXhFwMBAsy5KlgRp
jxh17JXB+a0e8bh4Osx7AjKN1p2TaSjFQGnZrMRuaWcFQag17lck7JV7uiP6qcbic7CGa/CGt/l8
XOLgQojIYvv6eoUUvz7+dbaN8TAx6nzoPC5ONnyD9VQ6zkO98QfCMCOGqHIjHgihsLCPX9zFFTxE
P3IIT9ldHsLHhb6BCQ3wM9B0u72X1a/2IHQee8Ry1skZ7dX6HLAjCPQBEDsHtlsRCkoGw++f48fb
AaQb1kvlAXPpmgEJci+Y9GDKHrd3wPafGwPSzrUZmYF39VglOYSbTP+zUJ8uTPhYAcMjlDyD9he0
eB+6sWtjGDMXpTvvk4xNaif8arOtgSAD00MfORqgF0+pk0jrn6oJFF+XNYjrjwPToY9ode0jX8By
Cx/Oj95URSywKQUtEgqxn+hBfmCff1bneCAyTlQdLWLoWg5C7bLBtCjbmkML3d3BE4XCOtNgxGDp
IoOghi7NnZljcOg6Pclc6lGOXwB70UXgwNcaniWujn8RK9LAFre1KMpNryEsBjpPOVa7sP5GR+r9
B2dq+aDYCsdQky+eQbrPwmhADWNLpn1Ho++yEQ2BcQou8zelt7QH1AQ+PXUH+aSTZi5wT1x9esfH
6ojrxw6ZayC3oqCtKkQ9tQqMzD6Q/hnnN/cOaMnB+0RcUNrWUuxDIHATPJ6DEX6/Four/3JDU65p
GANkWglxWfStlHETVwuWz5OBvEZzf/pDyfh+3Pq7s3yj8sT2VRn08pVPjOWT4Mxy5Bd8+mslDXpi
djNS2qP1A06ygETQxWBo0z1OkTvnvnNes20VOi3vzDIFj3ykfYr+3qdt0385cZ4MNhkYgzABn2Mk
ig828laU0KFD0js1gs+uBaNFz3sWWe6hQWisX22gdtLWLDExN7loq0sAktRyjifH6EyM3sG8L75w
S9PhHv/SQf0Knp4q6vJYiHjY9UMo2fSqcDsntu62Io8cRsAuvtyAaz0VZakU6I7aG9CFUgD9jFXl
JdOy+aF0g2Vt3s7wpfCzBBmooBKF0/wbSE+Yl4XXjjHVIJy3H+Nan/lkB1VbLtA2QiKoiBcGcd1P
XgJEJN4onpHi0w7hFiQOaKC7anyPaEzHlT32Bw7JQfKDzB0/WiZFt+UjvI3cN5j/Zg8UzSQuBC/k
WATSrGuxKXewVE4WVjy+P/lww0LRWseQaaVUncM+iz0pK4vgrozSf6fZUmgqRcWcu9UbHok3BAdc
UDp6fTce+ZUfK7JZNJ7Mir5qxdMM8utS29XGrkAlgBBfusfmgviYLCazn9BfA7oP1ASHJkPaX9eA
4L6adss8Lqy+/5QIb//dVe+sPyb6gyYQen1OhiGSlgP7jVBy+HqPn2mHOEGYXBrHvtziR4ajF208
GB/HevIlNkeYio6bklIZjU45TI9HCbFn8m1Q4FkSFYPIomaioHLccG50vViJuCNYzAFA7uMmEy/4
sfKGTq5cZUTy1pOV5p/t/HklpbafK8KU/RkWye1GbUDvx29ZQb8maJ2i0CjMKkPOPiAQUS4V7Hku
5Yrq4362mT93oN8qwPEfFu+FIDUH4tZG2XBm9csO4gcTmxRSe7tAS07+Ya4HwJ5l1iKKHH2NJL6q
P5NQBcsHTgSUmIbi2FmZGsNkm/yjNR/TNTNTB1qo5qu5Yh7gXLoVyp08z0HjciqGcMWW/Wxd+0tJ
me90dXj1fhpYIx4mH8o21hOdGdceC9Z+R+SdsaB6UcnQDc/ZgxYlRZnn1XCiq5snvBY2pveVJxyQ
nlJ5rMXkjxFysrZxb4JsS2fp95CQ2NfRycIogIHSXPI+Qz8ovCKLRP5vnROAc0HoSL2+wikNMXs+
oseraBUXi3O3IaKHosGxYjkz0xyDOEeMvunMQ5MHEFbQX0V6Ns1RmG2nwtbUJ26Fz4dQNgjUuYp0
0q7u3siz7m2BmpknsCjRL5OmoENKIxB4foF4PlsUkM8+YWM/gN9/L3PN1R2ZQlUtgGZLUvw5fgDp
/kKEhX7YT/SV0NuznHWPgsC/FGZPz1tj7m7YkBq8j/Wgw88QgzUkYFgj9ORKzb4ZeXcA07FAdvq6
B7QuEOsWPH6JTn/whIH3B4UcWCPbd/V57GI253wIVfvGwEbgzRue0NLo81aC6LV8zCWoPkC3SwWS
aOVTeEIaLrJ1GCGC5rzqTFOARt8jrvSm3c3gnvSIaL+Xg80RSQkVixtM5Ta9qIA1CjyBhdSZGHGT
n5BItbRnJlHLA2S/+OSSBb25NOu6pwSkUaeR6EzeeiOKW6ILxvsrTQVCBNUlF0wqZ4iXPLusSIsp
IZyGVq8G3MSZ+22HGdh4XFa6dZcupaQ9P4ad3aGnPlnK6CNE54z9GOWwfcw+lSaynGWT8DFS0wzi
fm6UtMYQLlgjt7ULOwgiEC+CQD8hX0C/CIFxYxte2Y9Xjv93Jz6Sd5AOiR+X+MO3YJFEFsRCegtU
WVOxU/77w0j0ua9wTYS4MX6HZRfnXJaK5n88OYMW4OzvOzszD7QO1Z8BXnz/fGFEWFiNQlE/j90r
ag5d7W+FzHlhQTL1A7EksLUxx18kd/h8a5qtY3Ai4R96jAZxf9p+64gVuEJxQLJxdpR0w6ZL/z4s
DlXs1bnzweRCeBKRh8hnnU1pAwJhRJZ8iI9XKJP7uYq2YkPeDdcGOxjErWvae+XQOaVyshA/xb7P
4K1H1U5hrLMG0UoBAL+bJfUh7z4z3U0TGOlAoRGwNSXi90eBRcjAdgDJ9S/sX7yzziDR3KZSBrZP
ZDxrUwJ+rGvHCMyqDgYnoO/icrzciBZgKTkyeUdFo8JpKCGnGlTtoz1FVF+dAOm8OsQ1XjMCBoDa
SorVrTxXKw8JlQ7j+QcnxEgybDXbbWOor8o4PIDipr3XRUoMYkDucnpuflkMF3rXURkzWb9UoaUe
1TTjSYxZi3Emno7AijHLErMQYPSP+wtrVraitSK6j6p6xPjVUH7yV+QGMXM9XWbDpfdNmYXuYldq
TbqMRGSMthOX9ImQyxablAnEl3ib1TDwjV2pM5n9op+wGacHYbhSv1xjmt+PUkGOaLj3YBb3x4m7
2yp1HKNF2a9dBoziDzq0Wrgq9uTSWmf6mQPJ6MphSQ5cPteyFTLvl0eY6g3KuUonHUeyzi/l4ATq
Wj1k+g+/tIfNqOX0oj8TJdjVsEYsLMFC87uIiwACUlYxHxM4FzCgA7K6KywicxcnoUdaryWWd3tI
S82AbUx9gKvtRbp1mvL0TpKLN7BLGXHTM0vum7tSaoIqvRwblOcIqKPv+i3Wmn2F3CITPRv5Rx6F
9dhXUifF4h35kTTtZV0Zq44lAPbNOIbSmCKfM53LcQQ4YkdkLLywYQ3Dfg8iayiTqHEqZONDrWKQ
oOt4OWvSa++ryK90RvaiCwar66CnsugO45h9HeOR5XfxE8NfuJfqJxq18XMGESuIkxnznNxjy6Zz
J6bE9bTzgrGeBfi+t26GDcspKxvhqNWcjKJzP8NnJkLMJlTsvOh1LBN90nSRx19IQV8LHNpcRIC1
SBq/Q/1qesTHLwdVbEefpko525D75MeEGTu+SWGpq7ZAvPDwJwlnlDSXgXFqcBEe4X07DNtEtWqR
rjCwEpjsB5urwFrtXd9wBvf6o3KppYtLDfMeZed2RuBUSUNdtPRdrcLr9mOeuGnhds7dC++I8cjQ
0VJjAB1PXUu4R8Xk/EmlJ3Mks7/HbGjBeOyAZsAZEa2cAocmYBWbr2jU/nd2hZ8GEBnFaY2Pv4Pd
6jir7zTRQKWo4l8CHp0qN0R2kDrtaIE5yszE9g/o8dzUU/HBsBxGjjDcgRWytBr8kbaJtWFniR9P
7CXe6rcdJyS27756UTLqBYki9KzoBzwysc+AXwZFu+qmEVDKkJoq+j9xTv8BYEiZ+2OrC8E6Hi66
/VvCqgQ9Ajefi/2uerrfdQSoKb16AmEpJkFeh/CbfHGjlxKuz7rJc79kRDwmC2B212FijWUMORf/
9mrCNiMLeeUZbAHiEj7PztPauxJKNXd9+/hQKKP+fjCIMXwpuws7yVbQSIqjpXJ94F1sApsGGpXo
Ysn10D/gFIbkNSMPgN2tzSJDkgH7uXZl12JFpKfAXOoIUykcwOpJtgClT6YmbEaMPd55L0RK5HC7
6i/Hfylw38SbN6JgilyvQ33eyizBDL5sJjE1xXO+c364DX8UgQicL+aE1XYaquMUaluI/nG8fjNh
ye4hEUwnoUMkTkKQrKyMUKFj7emgqjUoMn4hurG4rcaUAuPL5YWkrgk0Ts41qEkI0LBV0+KgJ9Un
vbRjFJPQSITJmM7x0eUkLleTorPVRxFFcyTkaYTEbf7igv5hM9Jrt2sV7C6zQ8Y4+89MuD/hfxKl
mHA1AzW2uxHUfGYvHxXyhrSLjGS4fyEGgMbo3WLvom71LQMiInJO6QSFmTNYdm7SXYk9NfcMn313
oE9NLEPKH0HHo4uofs7WSIxe694Kz7Qv9AweI1kUvq0ZJFcCXO08JZCh8WoE0IP6wHhadM5WRLpF
nuKMy7Gqt4CA64PsItv/Jsbdo8I5Jc29hzchIEL59/PHeC73lTxtiOI/dcmdbzdmwHxEhVtKARKq
lDucsI8HnDDklRnsnia8tTsg4hDJ0S0plykFT6Xz09opvRU7ejvaS3OK/r/eHkCr8ygiGXLLGG7E
a4Y4+qONmG79ZvzRwwWqwSpRBufUh0IB/U/8eG75SqKN7unZidegAARjMjcz+B8bCETbJe0JiEip
fg6rtyQH6Ozw8LAx7GOhFuwosZImIpJII2PU43BFUtJ/3PNYD7bGpLS/UZB2FHZi6s7DCnMRHwvw
/3Bi9PHEGkfGtl6IeMN29gN8aTp/45gmsHKPCI7o+JyWx5qpj3zCsoptj83Tu3g6se6PSVc0mBFj
SvbHg2qldfB/W35f4Z/s3vHLg/lqbFD3BC55HFc7O4GlcgjG2T0F21P4OWKFcwuttMPtl8+QJKHR
pTbWa+ThaFWJCVeBxL9KQLhwnJ6VnKSKHhgdPzo8VxYd3XxwHB2GeoNXwm256jnXiKPHIaEUsb8s
ymiXZ8gVl3JiWFqJ6f+QipV9mZ9rKzHDc8eFSeEkmGyiWBy+4UyENlA1CirrjgzxsO3b5wRo5c5v
3Zas9LMvHWM7z1lqD76OEZhxO7jdT4xkbFP+e42bwdLQGb5TBP2COhp5qMXMpa9ui0S0HJE1a4l2
ovYZ7/7zKun8s6Con1hUt+3tvTgzLPJd7+/F0SN1IDZ6xhz71sweqCWPyT4NxsKAaFy+MZiyulAT
TnUMEUy+ReMwkbo2DGVJs0Wt6Z3S2G0z2aoXmDJPV891RXPkuVumaFrHoibbFzkPYvGcWYl1+fQu
nNzHytxLxsgyDNLDFZ9/MPYVsv3FoNIT1sJbe/oB9E8t7e5i1LM5jdHtooQ0hQQwBuRU8GgFiK6n
6L9YA3mXnABkRm113SnXHp1V4H04vgxxNMY5Rbm2tLo2WiXjowIr2K0LxUkcSXDCdHq36ARXIRvF
Z5o8TAQMveCW2wA39oqiB6BR52S/3iApZFF4+yHlW6L+KaAF+40QukNb4wmf7MmAZmxo+6uP3mf+
JfZBPIaQeiMTYzIShwnkLqGhUqI15diqUroa3v9O5FPZiZJzxDGmAnohXK88DzJT8poh7PLln2Vp
ln0pHrFLcpvECezufBSilEtRzxgw1Y8veFMo+wjDBjLL8GpSvD/YUi1eQft1ahbjPOgC7+selBmw
pa8HVI4Ku0acCfZCUw0eek0VJiObPTLPbyosVEKYpQS/m9V7Jqz3gnJ09yWK1OyX4kfCX4w9cdgt
IPtPqaVpkCTAtluYZpchVWUvWal+kul9aRaPXpxsg29L5op2FNqQLHk+kLnkLIo4Cm40BHI1dv4r
rLQozBSSupIYTTJ6Y/9a2BC2vjEm+jAl9+g0IXQz/L4dpcQf2n49Rzg54NTRTLE8ufo1UV8djD41
uOYnvV0TtsKkm/5+V+0On+sUY7LPb9Yt/eHYLJLBgRovVJcRDCIwczby77aC2CtzrnjmLj/QifQE
x4Kr0dPsDLnOwikaq9RJOqWkpxeRwSFY30JFG5knxL08ttjaZto2PBlGHK+sCD1dgwTv6phBzEfN
gD3T6SP8n8g8NcgiiRRQn3oRAji/RNjqXC0DwbEQG6yOzYGUWLUBsKx4HkZw9Hb9EOThIWX5IHVB
xBA9zAMeQmBFOIAZLkx1Z0KMdvd4NPcE/HuKDCCyGtckoyWVB4KfwI28Y13zo4NIT+OzHtbwHFXT
VDY5httMlUCDLc6zWyvs9zR1WwKGherIjDief5no2W8WbkFAFxonEOb7px23GlyzFpXOJo6KcvhI
iUyHSVnLaFsJSxwjKPa+aQZpaFC50DgfLgkO8Nf6mlX485FPsV4qk65MNcII9dwcZWbbd8B05iYe
G+19Kmf1yfgxpdNdyIpBplpQHvERa7YD3vNPWY+VPcc3kkbz1AFJ61M+NEVmpFMVJ8vBFdD5krRg
MlOhZQbb7g0rK1uTTEZit4nU1jP5Z3klQi9H5MY4lUHsCaEHDUj4sp1ufKRuAPVtZNfoYd3qZ8cT
xVMa82vKomPtup+z2FateAozD2JednzdMyo63JSHvw+b9pETnRAlWMEY/BZuVBnx2jcloWCOWRzQ
k+rOuVeb6ScLVAmMJud4k3quBHYwngtE4CgOKNXIz6hsX1wJRIwXCQWK+RmS1vZir4iJLGBJoo8I
yJwqvV/wAcdFWp3VjV2maawBwsAJsiW0psTzEPWJIkfgYihSIH1DZDE1qG2mnJPK5iXJfJSQUi5I
4OJB4azCRhWwE71VjvtR1sgMqSQvFIyRDRa2ZrXM6Dxj9fNSUZRlDHnqUnvLLOAevstz9Jr/c4T7
tBVKROB2nSTWTd9fGimL2taqRT30Rl7j0nSapvQXbs+kGdgg9heyBFAvcodKVNa27e6brUoTGK82
8Kd4dZEURKxYwW/0l+CIKEz75eUb0uqzlRNmluVHy/8yDyolAwNuHGUgK+M4aTcMXGZ4fUrrH/YN
VTrnFyxT39nzizylxH69U/UZqs+kkum9yM5NhJjrfMAt7PrO/tMGrifJC4t4L9vcX8UwGVZcyUNa
HBlULWqhsH8tl/vHH1/4cKbxaZ4DSNejTMczC7BUcWMteJMo66slGhAuy58NKxIR8iRqx+lJ5P5Y
G3iAAknFMMv6dEXjrPZdDq7IwKS808WN9aaxU4a9HjE6l9cvaAF9QD1+WarSywdgA+hMRm/cKIOW
5x4CEyzZMhDQLpyEmgYA3jTXe77v3RvRylrFWKna3ovNJ5bzVBa1VcER1/PeEGrJTjoPJXDBCjdN
xFWMSspiB01DFrikCqiBgc7FtSKPpTskHusAR8+N0zFo0bAI0ucca1+ct7ITkkAen/reQYiD/+6j
bO7uBjLn/Xo2/MVv7+/yFz2jfEbwy/VP/Q8k+INhDSjSuqgsV5z9knd3jdnWjLAvGPtzD+Re52Nj
0Y+amOSQ1xCA7c6MNok3ZwvBbnDDi4m+MdwRdxYuoItFWbdREmJ/PQ4JVRipQngrYrJMyFoPVlms
cuVjkrLM+R2wxZtAOzqDlf4Um+mRMuN1Ow+f9gJKLxywHFp195yKlP9kdG+nbntZ73fRp48nlmJN
sJvOyXS8MPwnJhJk0v1y2sHcCRDqt4EtCf6NwqiquQ+emrLDOdoPaXhQ3y74YVMTtfSsqn7TYbtt
r/3lT66N/PpVgV1QrTBfAGUKsU6t8UYJLu4ueYHTDdSiNIqaCM+Kto+tLSJZdgdLv8nbxRVS1tjt
MKmNXwxV9C+0HXmqmQSzEmTWxGU+XwW0YKR5OW3VKZqojikZV1ZhQiBT/3QAUf0LoJRWlM1Id7JI
mI/fFhTbfOE31vpkAs147QkwYXu2fGnPHiBJ4ujlqqaHrkhErjhgm3+9X6WVAY0KjkbPvWtveHf+
BIH2uwKJlmWkgU0qIlOKCLJxawHUC0TFjs0H/tGCZAdEK54uvCdumVyTXomZaTKd2SK5si7gyorE
EZhCILdyp9hHOZDSgKPTbIQan0Hc1iS9ADuJHQQn1dhLQGDuH7CsNEyngAWTkYrT8Jr3Am65KhnD
44Nt1KCNd6AFL0w8hTUZd8rqKps8Ex8Ro9IJ8BNITt0Fix6lYhIwwcjvOZvWorjpL07vBuS+VhCx
PFpeUEd2RX1Q0+kJqf6e9zzo5BE1vTLzRYsa2MA8gHz2+eGWRcJJBOF4VHZq7tZeHM4HJQYHvcze
x9kGUOu1e3vw6N83O7cAeZNkaMHxR/GRtIsg+ZK88VWoYAfEkmEu08cY4j/Sp2/XHs5khikd0nna
wW2TChBHTGJxRTVQOJcgXnMGwOC+eMpBD4mpgluzpFsWK26K77ad7DSXGP7XmbOv23xPdwfFRqYG
lnfk/6iK1Wzzhvw3M7mcWFFrWvQdoFihVEYhupI/RYxFQ677c5sYVTWF6UJSSV4KoKaRjS+P22HA
mokx5VIRrKjv0xaCM+i7SNq2D/b0oYcCGqzWxNBG4NwjmVhWcFRGtmRe3oYL4+rf4InFjno+g0Bv
iiQ6UvQBDEQ8fX1npDzPyJvFqsnRyIMqrWRRfpkXpLJdgex4I5S2ULdnLFDo+hO8N3hYJPdi+yEc
eloW8jFGRvXbV4/si9Tm3ev+qlz/KF4PZzvV7IDTyJ+VrudvRyihaIDe7KRq4TgP7TgL85lxCjHN
VoI1tzJQORB05llM1DHAQHt07BJ/ndHySQ4CtXcMbKlMTkfKFyyn0GbOBAT1IYtvyYO97sZGPDLs
rt5Ce73jSrR2V7rbTg+CBZ3gGw1fj72aDm3IZp3K99dM4UmPQUI1P0YM2DMj33Rxtr7qaPTyTgbQ
dVJB+zl8Rt+TtgOyY6JQ4fLcP0X9KDoqlOGkqH/kPMOMrwVqOQuA7ifuUaDF5YwrV1s38PHkmdhW
sTAgEusNCBBJv1HSOWkksGMgqmNDK1UVHcbppy6qxIlKa8DQsIzrOJ65kQdP8q5AyWN4s3GNrC7a
nTySiZLWeE2sAiTVBy7BByNqXbnpQ/EVZdls+S4ki6QyVBJB5ls2oLluIzTr0eZp4ihF/UjBVt1n
kmV6pfBYSykXTG3Ofx3DwvRcqEUwmbQ/hso6fH+ks0smn1od3jFqtnRkM3PS1sMCloq2RJFU0W7X
4TBpIGsmh2kO4j32eyl5ZEtQznkmtKMoayobzHarEF9I7f9koX2+p67svPNXZ/sx9uZGAjqlW3Nf
WufsYFbyvFOjIV+3PpqW9YiLMb8rt1OtWIsi7oA2eYTnGfA7gt0wR6KwHF7GLWxCGCJNS4oTLVa2
ZmftyAxxunEOABhRkV+nqyAMQaNNDhArATOlB66sx3b5d4Kp8Lmpq+1W2TuEs0YpNE/s3s1bVxIk
I28t8d8QmKhOLmowhCzbo+gmsMIOXr54A3csN4OR82u7RAycZ/wdNQ/s++JOrDa8bnlsbJspqOw6
qh4cUtxVF0EwAdraWkyKQCpH0I7VNGdnBAOaRcbTiHbwtwPZRuE2ZEuFimwvjkVXGVj7P71NHcus
VjBmXFM1bJycBrABglPh54JGWgZ9n5oZlFiMCWBO/BsMZSSJAdCEb7Mh7kIWns1bMlzrFNiQ2Pky
xKlwrRnqUPsyYEQrvfB7Di1RtvFirfvkPttvQw7a6oFjeP9J0qLKv6kjoOQw82SH6ZhjQQKHS2fm
PMCathsDlyLOTOdbAhHfosi/fttleDIBeAKs9tYbQrcJ0GdI2gU9sykSb2wiC0AjhmhOH0UTrrW5
IIejGirTma/O8KrLBO/9Mi/kAv82c/bZRFzCXmI4r4tLPyvnlYzyN+vsl/sKa8RfWZb2pmEG3EYC
D0xKYgGsUV13YdH1cal31g4M/hKE2j9Ctp0isPMLaf8M1uaLmmxbuFE92Wxowrl1a4X2JQ0qjeYm
6rMzBkrdbE5/mziwLQ3OiZEWhxmL8pBldamhJ6FtAHx1hqDDRYuWdt1W6yzvlWAdiIjwneFtOkDt
nYESkTnduO3FXkLOqlMYjjNME91jEadsPeG4zcA9eEAQ5YCxomAmgI//HZQc1l3l2+WMINwz2Ya5
zXCgYeP2u2+p+i9i6T82fKPejhNu/Z3Q7qviZ784EJkH559E/1ICaDyDMTqMg74tCfGP7vdhzX7E
SnKt7bEVBgOkEh61WsPzaCAC8wspkKFs16SL//grOyn/aeZpeFxCwDwwhgzyjwDmAhLFfPN91sa+
ISayN9hNIDa3ie0Grc9wSsGGDKSYbi/2C7irYgNK6yiRrjbHSvp+G9r9oRjKRCq34XHxj/R8YA5i
lwPfHtX3+1teSNobxA2rdQwJswctQn2xSvHcaEATpKkzVcc0qzm3L70b3Lcf6Z7NUqUvKNCwuMHZ
fOlC1k7/YzupXnxbOtsSRihKIwmCLdpKoYKldczsKd94R+F9kjlVsYzvHltv/82rPx7k3BEWq4IL
+1Dl6ZTJVlbwTrJ+DFgEppKu8W6AWYpXKrZ8hqRK1r/Cw9vQ/O1yEOJW1/7Flh+8UsdF91Z71aTn
5n4v88P0JzHweU2QUtNJHeXzYBSbQLThbAoy5cIwr8e2DobQfdHrfVvs4ZR95WR9YkKggsapmfXf
kqhkxPnVACzBWLVarFNU9R25UoF9BwUvlQYpYA+Dv2gustW1rbDLrSuZC10CYryjTawkkzA9fo5V
763X343Yz/TYqkctclHnibsYpWzdJH//Pw8H2l80cEtAFy60kZzgSWt+OrhiZN7TO/1fq7cUeOv/
+v4v8t5tlgs+nfQsBb/skkZlan2svITQhJNRawynE9u49SPIIdVSvyLVLEk5cTOCfK679vUXzVIr
4qiXfWqFwSABcpBJawDcNRIVa0nCLKuDdMb0twyBCL2Z7J5oK3ki4wP0K60C6UfpO8itQezGmDpM
6M9U1Y0BU2guMRvW+jLGunpAyxrZCmaZzqCRcN7DYzQ/u+8cz/m/RK+xmO+x58tdUA2xJjbPurZH
kIPrTxgWct1dgJKSSXMjAc9mHznsZqJmFckWQx2V4t9u9Vi+nrt7iDcoEXHTqgTBr5HeATupHedH
ml8YMeiIAOiKTy1NyaqlubiikOALSEYwAWS1PEe7nT/5E2D0t4DoHns7ffSVL95OJeo1NZSoIVow
k+yIEYNnutQUn2eE3a/e8uoitHSto4j6BoOjuC0S8pEmDOJj94bTXb16ZUaN3vz0ByU6nGIlrXlH
mxfudeq699nWeNTEczASNmR1NRXEXVLVCyZQtuApzzba6NQlnlNmmVUDNhq/Zi4qVxnKf/gVOpp+
2HixUB+cmPEuSBfYlH+xJSWEayZ/Fi+r0oWBtSxxsjGARtWhvdcjzeotu/08W3ZKE5804n8WuyUd
4S5NEam1z0bpZMvKj1ldVP8/vwVcEkINgn1yxnz/ZyWiNhMilN8XZcQaSysBORgoR0lKL4A9Q2YV
h490O70bCovZXsW1QG+lhDvwqLMW8eJ+DL/G2hIz0MearW4FF6CcrnAI5FbWU7QkZ0m8X5j+v/f6
aKN5uFI4qSgyBr7CHqxrrw9GE+ocMh+IrN4E4sf+GFl573LYFpzlnwrNUtnUrn9P0jRUe5TncqR5
JrVm4GHWcQ2EdaxnxbiihJV1aM1arA55MIEuIO1S7M7tVeUlofmT0SFuTmx0tHZcsF0lci1fkQzy
h9nONmcFrUXx9CR5sFGmKPVZ4Ha1/7d1mEX+0GDYchsIt8DqyuC5QCul6JQ22STx/FFlK+Cs/cdz
bMa1DqUah7s3BZaaIH67a2mK7OPVJQ37TetLsDzPwLEmv+ZJ2AKB3iDMy60UNwbNhjXk/GAtYvhL
v2uvH3cSXvi12HGvgCiR/FLsp9FZ1/3CAGUFXetAGHsP+CQhu9sAqb1/fTURrqJiz5KQ/uKUc2cf
eZExJBvXEOJXSk+YIS0zxO5XiMRyQLLrnRp2U96oY5utVgjIPIZgdWeYTf0aB9TMO+TQuwmwdIu+
KDLGuiZHB9ih5tmqrxmnxL31d3NINj2ioAVyn1+1ICwkq4lyJV7oEoek6mw9jOXtSc6Io04wJEH8
a1nCnw0BFhdWBvmzVKY5xgs0XDRVfcbRrcmYUCpVbBWfqq7AqrUsYdIZhyUnepvQDXrzWJTfk0dc
5gdmz28Xvqho9elnUYRMo8ZzIByqZMPgy0iLSXaDKNzIZh0iHR+1YAux6TkR0X0Jo7cgWsLTmgL7
QrI+TeB9uttHfn3G/PBNlpcodGsVSOEl+bzN7/vWKGcQg7CBp8oir5HqyFI2uvj9FPMJjt6GCM5S
CQmqreWCJPn57HqG+0pWaHNdXoosPpRfZ+xTllI6zAfA3EWSeHGPRARlyAOfmy0O35E1C6n8oX6s
gEKBYQn9byJLiyznl65o42oNQlq8rg+HDoQJkq3sm0zPIwNcAGiB7Bai01ymyrGsuyBM9fBiRe8I
1JFU20YG1FalM7HUMuGLH2SqdlYw6/nBjF7Dlh9v19Ik+NFr6IsGmpEeDGZ7MUZQQGAwqaU/gBg/
DPBD9fffftaX1xJMuwJRRNTj+tPYXvfymkldl4VyBPF8ZKQXR3MxgOtBVykF1OHv45Z9lGRkzh8D
nlSYJAGuxdUx8xFKqk6EQu9mgYgJKSgYxW8FxPExY5qlCh3TsBuJOVNVu1qL31no4tCzX+polifI
B8xAsDsqcWMLyP4fyqKOjWuHUGUVrNVt4pAXhDg29/W3wlLKdQ8zdpplt0NjnVxdpHnCUrP2fMWv
+3/3EH04wGKn7iRDKK4i6g1GzLK3l8AazEWkTmdpI4vBwDbe7ZpZL2MdKiYFkN/guFvzqEh83Bex
XgcN0s6DiRa/DcVF15jxUT+eyamnjS1dgY53qIos2/80h6KC3ZVwmaKkoag3qHD6vcb02ulXPPHP
pH0Mm+S9/t499kNssyf14VBCi9pwyMzbFGX93iE1qlq0BNrnW733DX/iR3HQP5L+tnQx/el1VioB
88D2rnacb2JETRDsIppLzUlHPFuvyWO0MTJmndLeZ3JoFvzCn11mtvxO2HGPW/IfT0F8ebBlPou6
ouNZRVRIROm0/r362WcTkyKjQmOSwTzUY60CiUOHuM83/NuG6cfvwCY+D3t4I4nYvq94P1tk3jbx
IbR2xoxHZ8vqniraaMX8Dko641Tc4ohAp9/VnLmTzOltNZC+WwIrMfz+xtPbeeVYqs6D49mepZY1
uP50cJ2ExH4TAvXpLLinknPM8+vLadpOvzThWC8p18HTcEdHtoMyQErKOMb7AWxqOMhl7Mk0VlJV
mcbr6IaTVAxPFAGu7LKEfvxZIkCvHly6OXhCyQc060wpkYpYLGyuWP3sJDk2qHqaHAKGZqex2QPN
NQUszsqWFGqxX8fdRrvS384b4ITy/LQolJAh3zLjqsDDEdWxZds+iJP5nIqIsWHATKcCfZVtTbnt
zoAvGnDa0gd58HkGZ2+G1A4z73uDptMcNQjAvaLIlO0SnnyRWuqLc+rrfc4l/eT+8FFl9eJu1Hx/
+tASg2vJeEgju8dtqKDZVgmzCO2zb+Xwy1/CBZcjstKOU3a+fNEC0TrUsiWRQ8N3+nNTEXXLN1XZ
ykzv1Nzitt1d2GZU5XYJchJ6CkPriB3ir6WhhSeFMfMmBUFvqDg/NqwudMb7MfZEZ81kRmhmcyiu
J1hkIdkVXfKntgm3wa2Dg9152zOm3IXldPHCcky0VIYfwL0xTGxByXUzTIBMIBfhEAn7gVHvC8fp
xddE4hjwnkdjzO8ScKHA3v04aGfhYy5NTeRv0v0h4AxC/WNtdRcTnpQd2IE+bdxNNl5WGQ0KAYym
tZutRitr046MoNKKK1n3fDdDH3FdIgtpN8WY64DngCnhlHQ6YPdFL0N6hWn6lVRzDFDOTMg/k0Mc
OFX94QUktTHadqAe9G+tGn4SOqLnav97dvRJnE4wcNaMSOIwCc0Is47VEOPafptUrrR4u1tEwKQ6
LKaVQstOxCycDh63GMn+xmm8tRn2XtaandXxjmoq7gngldF+e9OSUx/cgm8Mt2qFv0awAZt0zZ2l
TQZhao+iq379DsRZYo7oianh4zPJLkuA/n1uJaAM8ieT34IHGU96JFOmhsZjoNz8FOwyjpJnsQoX
7YCAPW5zJLRerkBnwHprXhmxZjyr0Sp2dXNop7c7lboQOldPtVn4OBVf2koIQeDGjdyRoxN9w9NN
tn3FDLut29YexALnQmtuvNXEJjyJP+aRLl+zF2mhYg/ev1caP56MKK+adTg4xsmhORg8FY5UJhSE
KBi7uiutNnxiFBw4aZkskA3j0bq+cxv72sQXhSAnKFQnhrGWxi3b2qOo4h1jcF4baE8hL85/aUWt
Z5HlZYDyyThtlx1+uKnrbBuGwpz4by75GYWaM1qxCZyip17BsjBA52t5cpwgXK3CIrZToHgkBBrj
XrjxGFIZt/yNZMhXKWYjjp84wG0KIcdxbnNHdT/s8UgwJykMdk/db9ojEO9KXh3WVQ0XVqDDLWEO
xocCagK6ZIxWl9leKbUVT78RieBsUn2uajxQs7L3Sfb3bfN+yfAXT7lpWNDWlddICKFmbtHBiQbE
MmqMP30xdpQZN8qoFuUiq7YoL+Cd+6PJT5KdXLqxabKwtsLpDjrPchzEtXxSbbmnPYr+KptPVTlP
XzQmo7mJ7FCq+8XwQXwzda1b6r4WtluglM2glMniQUHKVLclICjvVN4mFJlDViTilpIvy/hr0pcl
c8qT7cqv5DjH8am3EbY1zOisREeictfdX9erYoZ2dncnXJo99/h+fZhbbS3/dm6ZEbwHQY/nQTDU
ORb6vspiOEhXrGdOmFZOj5o1EKyfP/CeXaYlhR2n6EI+jW0mRq8iikCOEJ/lsREywebetLk9i6No
4aRpxcB8goZ/CtAxMQiWP7SyG6J0wKkzb8KFhc+iUIh/2paLAm/tGbAM8/TODrSvd1QpwL4j6oij
djjg7ipZRBCIFzd+NDA0E7xemPx+ShamXg04XxojRTbiLj+qfzWOUiOKzH6buD+f+S+hiUp6JC5E
Rh1SGcdBvBEqu1b6Fh3Ns1cYGia/xZbHV+xGRmde/o2r2O62QOH1Xbpd4ksKgUSBC8/hVpMxc0In
xH8kSKDQ2hu+UkmleqRXLdq/nfeaaCz8Oo0av932r5rQfoB9pQjs2YIG87UjjEHfJ2RVNjKu1oCZ
yyuaWJCgygxDmkqnOkL4dOzr6YvD2MJFN5ziHvDAPxaq4Jbky87mA+D/eFIIautRtmawjrxXaEOn
T9yvPmhpb09fvV81novYXA0dNaHg6AXyEnjFCV+aED3GjkoSwoO6G/kHoJLDUJQ6chTRGXLNEbuj
fsB0jQE1yJs+0ADprKdYyBkafL80JePdmnTT7S9bYlYcFu7I9ilmoEo6HfwTlKh6qYq2yaeZMUso
L+6HkBYPv5oxRHVsDVJ+KL5xwrVnrutXWLMPJ/LjQAk+U7qEHJhmtcPrOKmDmwVtv/mA7Y4pVjB2
paiyffcPzq6KRgHuUGMwjD+yfc9DacezpoodnotUaS7/hpsOsClOJ1H2HwsLmTeynoIBQ9TCYEOR
QE37/X8RHxy5s7NBnvZHZc1nfo/zuT8RGoAf/JoOsHheJos56n/BdIdfN+fvsvtEaTq840x+DLSd
P3GMu4ytK9tsMOtQL1jJvmKA1zh0E7PtdRQX7FJ9/hv+7Jtbjb0R5ibNyWskWQmkOu8IpL72xSt+
GDKhr+kYfC5FDLlEpI2eiETuyhqNA4N/xxcjVU9TFQFmpgHyXP9hblmyE1qfchnsk4xbCS/akevR
KDMHmWssA+7vfXgX97KQRO7F9aV+mrcIAwanXCOtahgEcCJSH+Tg68yn7sHSf1ME1z81CXFtgcdo
iMstxxR05WWftI2qV3m+U5jXerbYkUafuCOuvxA6tq+aim0wF5OliZntOEomDqj3a+gP0wGfMGYk
euvFYgHbUFKq5rHwHbpi0TOT1ChaI4H534AYIkvPAatUytyFwf62ZdqKL1muif6iROdOVbtAWW9i
wYnYZCVqYu/rBmjnx8SThVTTtnEP5qQzJMNRwS6khfUngQlDwyC1z3lr9ksk2bfyAOpKNF8dMTc2
NeiTiLgdIgb410pTY4nTz9MLCRRMxaPe7r3mOn2uWQVQGhHlA15f8bz6YaxpA0bL4yAr/9Tjw+dv
Km8ZpWpa+y3RHm/dJC82Ar0JEbtUSSbIsNgWhHrJBjz1ct66dpBHYWmBeu2wOe27hy8xSoRDhKel
brjNTFEJLTom6d8y/tv13AsjK5l99BxO3ukV8+b/0w68azxuII+nBKDNU8lIhFUBYokUh4EEVSmb
0+hCSKMTC7hL510YGFtYanP4AiUOcZwDj+cwy8Aohlr4hk//7YYOMhHllu+S81mg5mbczy0h+ZQb
A1ne06VoRmvIBPSkC8NMm3+mfvLmg2WcqLpetKGfF6KbFDYx4pge3AFeE/kraNvSO3syflON7gl5
HwLw0Z8EDYMvqmNLpHIobzEeqUx7NDxVmYOPdyKhd1dfO0RPZdv3XcPDfyqfznyX1854fVsksgAG
PxIwWtjInt3ZXR45pQffR27PffhvvktiPeWBbg1JyN/P8NkOg7V7scjB9feRlgQq4mplo4u4Uq2x
7Puk3JW6OPr3pPlwi9MQU/4zMSt3ts+l+AP3gOElHrb+Tf1tlGbpFuskIgd+BfqD16herAtJBLMR
yoTX43KboQJY/QIGKvJaiEpHeSbmONPheu0nTwRtOFu9zTwj+kR1yJqPI/kW+5SQ2/HXpE/KPTLF
zMd5oZpU8J/GaCjxbCPFJBKqIOLiA1Njtg+EJGOv227RQN/lvysaO2K/q148zgFypxzVsDSSMGQV
sOnvAT2VeeII59atY6Rq8kkm20n58PFMtRnfsuPehBm9/4qm+31601A43rgo838Vo7V/bU9Ul4f5
Ss/2POP/tZxOX5OKvFIDHffd9BxzQaQcobdkeJ4bjRyQlGv2l/ZNvhbD/oulaE22CSZowdtAu4VS
30ciQsSwCy+xyKp5796QwMZEN2vFHBbKDDHLUmocteuhRQbBI7gO4i/1QpgmSV7wqtqhaPm4GYiX
5k+98nE/3Tc9acWG50TJzEBiOwhfSLMJSeUrgbli1QQBqnwBhgaH5jW0dmzHTsChIp3aAoGi05XH
hFFV9fvewvKk+3n4eHOJ+V2zS64r+P3ny5VFQ+sMcG5RqXMBDVYsImmkpyNeeDYeK0oip4Si9sSx
DmifnGuuuLF3BP5Kifm+B8ZaRrUHuHQtNn3dPWX+4K7dOLCB24laasVjshLIaDz8BSE/L2Zh1/Hk
OJLZFLQhVtJFaa0QqfjcnaKfugMdMrP2UHbKgPiriaszrPwIpwmOxqPwukFSWgFRgFtOx1xJ+kDf
1pvyeffVcAD2b9Oeo1DX48177Z4O75nKno9TgFBFqcdA68G9J7VbVsnWnSM4EDO1Vakgx/nQ9+k1
Yk+ShHbIb/HEArT2DCTS0IJcONFPzp+txwOnSxjBhe+arrmwOyfxGpzoiPJdM02g6J/dY8gzG9LM
Y4RcCu4OqH4DLBqD+PWuPL3sAF9swCOE20b3qnAEFawhFmVqhdMO8oDXXZE6CiSiWT1AC0y2T0DX
YUjjoCbDO1g+9/ni2QFRG5aUy2ka/NdfDX7u38TN9pesMcXylFdfxlCtsEt2DDJUqXaMVjCZ+Ne+
fBdvBCOvzzX+xOJMBFmCVRwwHmGCOkgfdxK8eYX/27+YEjVWFYNVT2Bg/LzCDCgr+3uAS0kF2ioH
2vMCkv5E0pnPHSyBrKzgfVTfELCe3+MNDxR79PcQF+dw1oB+e5jjGdRDw7ZlkGxtY/QjK9B8eJlB
ZBahkNMlIhzm1BQnsH1Ehc96lAkdiwnDCh1Vq/+kJbmKJ1t6nbZptvJNpM3sxxrcUlz2O1oPaCAt
7Wqel+kRDEiS4y+StnTsd1zWqgBg03HNUHu8FWAJbIt/exZ6jUBmnyQIiLfcJ5pgOBI/wKiWxrkR
uOFeFZO38n7ms4vgWmG2RyLZR8vN87SdbqeQGDN3tbL5Va7s11oWdnT+kL0609Nq1YMge3sC3coF
DN9x5HAQvDqEbw3yozNi9j7WvP1kL2N42SWAeNJVcIBG7aM0PsZ2coFcIG4WQGdAsmcq7R1/Cnfu
LIQFcm2rgEptwZtpVP5AXlx0xM1nAoIXpG8HGykNBM/3vhC4bDlLTlb3SMgIiIcQkiBC/OxMYNRC
XRabdAoitRwvskYP8+jMnbS5jpWuJ4NdWQYODBAfc0zWpSDRGkWZLOx/fQa7T8omL1W3+dCBRugO
6J6cyLEp+iEB+vXAlIcLF08zgSGx+A3j+t8Rb9RzAl75hsPL401RtxE6s6l4hf5bOyrCvTGc2L2C
FxaE2Fo4ejjnYXZsR7zutERz1hjcTzOJkao7UC3sZw+i0r8f9t0Y2gTxbp2xRc0TGy/ILJrrcM5p
OlRaobUjp/qtbdr6TlqvjO685qu3uDeNDL7eGLqgilJLVMO+P15rcDgyAroRGaxBrSjdYoM6QMft
ktJNuay7yZc4hAagjz0++j/mN88v6SUBar6JdBwNjqhMUiI4d5eycxaLZWg+jaDEa7QC6fOzmqEM
iZBBw+Qojb1IatLxoZa4lrIxmeRGvapU0/iep6rWR2thHNn+wNUuT+Svupc7Efnr5VtAzi77U01R
0bWpe5olrwDu72q058H652Bq4Pg4eBd7vnzZ1eWV6FHN/78ocdKHyCs7z5Gw7hVPTmFK3aDDjwrr
npe9cKAaqICNGK6SRMpoOu9LwT6zZoSASfGRTUIFmfWEve4SGBFAjdKSgW6ngo3B0XgROCCvE1YH
fdMo4tf1N2stTquAQ4SlBJGdo3o4LS3jBEenrIDlguZ/l3W2lWrgiibRKbX0w90i4jeRARR9vEjW
WnWNDVr7q/3DeIWf7aFPjPKGLnZobqNKZ7omhTWZyqR2E2gMS5KuD2ux5BlqGEG9IKGuDrukcBJa
9AiXMX33vyehJRqSzwZRVIf/3A6e0DXuJdD7RgFZXWaIMrdqcX3mTwadB+2Wyqm1si0/q1t5J8c5
6/v8rvrHU46R9OrkDrDcG9eNfFtNIKDWkYtvhvC8bYbFbcXfzqLilG7n7T55zyvuhcpLGFiuwFVe
3Bwc6Kd1rMKpZRaa6VXUWZW8JYfkJylb4KNxBVQnSZLor9U1U9iD75XV/entTkl+JhZHAT0BOEc0
fCIe2E03YdcL+XK7M9EAUrVWzwgzTxrO7XLInlavfjU1C3yMMmvnsxSc6J0LWtE6jcRICTSJSbNQ
JIJRpPYktpJWISS1O6/OEYvXLEv440i3eBBl0p2ByDo4/Pi2NlcRNjtAdWu8OWY46F8KP2denHoO
NSfOg1lSBsIcv3+MUbM0YtWkknPcNIQW4cpwRJnaA9RHlxBO2OTGMgw3fCxwuhPjE5IMShYSqbxO
Q0TrKlWdGCTEzwghPhA4dCUnJdjLXh8HLctPCI24jUGaCfYm9zZ/7bxT8gQrdcpgNb9wRkxwfarN
U+VxoQjw8zy4M9Zjfq1k9LcQOePNg/v5xD9wGKBFKEZQcKAvlxfEDn33WC+H30sKOSTmoDZ+0tdy
FTI76HmZOkWubmPec6PX91ooqArWIrY4kbC14yoLWGhudMto0dVvBJdUXsIUo81bbikbk0aMOk1Z
FSMOUfIRPyRdL+6M69XoM24BDlXK4amqHtv1ZOH8R2NGeLzk47f19BpHolbnmKb6t3yY0l7OJUEW
Y52Tu80jpBbv2XRI1tPoTAhxfNRBiQ6stjHWPGXhRgAPe+hN5Abc7BP2F7z3sYjxNNPoR3y4bJji
ISxJNBCM0ISlGej+q/z+8b/Pze5dQCd4M7nRyLRN5lRGFcrw0vJ4VtaL8SMSITs1lfSqPGXbqY+n
8uwFv+O598iMrv1A6pm7/TZjkW+j+xcE0NU7I965bNsEslv3amde+Njt4I61sA1/blWE3+UAouYS
Ttybicm3F/AAT5Ia1WOjDUiWjuufTPwJjTbADlk3L4zlmilb1trJaoM9SJZojHKViPQDgA5J1RCK
zeHo5DJdclwlK99L7WgZQsrf7wieqJ5le2MLCr6HjScgCFZ5hjTvwLIrWzHw8vOnvEiS0aA2AALP
9LGb3B/WaUmOdrUpzQXhS1e+ThXw3GTn1jQOrbQgFihcmQR2hkl8bT0YVKOg2xm01iUz1qKUg1YR
8ulVVbkAIMzl57sw69f/hWi04fBQNSl2sPGvUiRxoieVe8yJwA/8UdTXnvcXKmL2u+mkkOpmj3Uh
AZ+OwBCb8I9s+1RFv/HvuAEABjT1sCTi2YXPI4wlg7dGUChPWo4dXEvK31ZSrx9JSZxL1XRmU4Dy
mNF7MgWyuKaVbIN3jEc/ZfBkSkpQOAU7xfpmLSq05NK8BmSsluw01iKwFNn0eKePhyHqZQb3PdaO
J6YuRsBR4JU53BuE0mEryyF2N8Z/AsdV6THICL/Dwtks2oMCwD+9t83iH83aFVNECLovGObjEnWe
BW56yUbp9uFueOK1Z+KqfeibC3nasa8Hlxewa7KTT+4xRPGOwnWUhWweR4nptNidOu/o1n3+nPT6
7SWp2gREdrqGN0Lg/fpivXNrd/NsoIfYNtOG2jGfWtO9JFqwkyn039qj3aHCUOKP9IvNBvhVvnhw
DVfRub9JtNLSyD97ZUr3U917ZkNU0ZO0dmA/OChR3ZR6yenGEEQoGaVn2H0NGw/jkCAahOogghK5
eOyXBgUkICHXK85WZ6lKwAXcLVpW78y42h9sbKyKzI8egBqkm/nc2WgWFcXM0YQDXbPn1aN6tADN
Tmk0+eVIVXX3VLbZlGl+GmX+xBF3HehBFVhVIE7HdYkAK2U1EIEvtOXs1Lis5xT0Kkj3yoE7Reph
4Lj3zQO6aRqYNkoRecNYwXS38KVMINt48EmY/3ffz4GGkh42MqCRl1Nr/ZHwKfcWVhh8DbPAUkwh
kUm1FKR8G87L6TBMP1o8n3DVuUg5IGiXeEem/Q/ZoAlf0LKorq7lVRxxj11jNAOkHC/fN/wiiIoi
iV4ho0I+ZARvbtPQqvHw9N7Uc+8jsQh7T3hCkYoPTfeHbnWG+3XbDD6jnb35jKKUNI6+MpeglwX7
sHZzU8p3iA4GUwMf84DIzHy+EtifM1rrTiQC+DYqzEbe5kXyEABz4ZrjwMDO+gk57cvOqZuk5ijF
5QHcvJCC2qtisbDLvmF8sI4wZBPtCIQQMn4Bm7hIFg+JA5NsyCYVbdgoh07pya23Y3lQSk/dG+J3
OvrlztBqPm8J5KDm8rKWlhb8oi3o5mii9NMPg8PZnCNywSd/kFGj0vzqggCHz64Rj4JrhSkOwljW
MWJY5OoPjBFKqC+XiTiX+DfXCauEFP1JJFS+W7uN6X9INstoxSILXngTdjtfQGEFVCM0ohwgZ6gz
Fh1CKarED4+RUNac37Q+lUePwcg4CmsUxeLWwQVUZPavdoNue2vh5yWlSqs/cDDMNF3SwGXw4jx+
1mvuJoxqIR06/twdhPiNMl8M0pU0vQ3hDpexfA4O/7PjvwAJG5QHKP9MB6ykc3IzkVv6j82vHkRT
bSafC+k/A/djpXeVimLlc6FfRSoVLLzYKO2Q/QRKXjCsG99FXfg0IdI129QV81AWRUfmLJ0W6szx
wjdDp7497DtAFRId4hLoHwfUxxqiK7+bS67roexqwD+hFGRvFvH3DApekGF69NDOetVFz4DCiuAf
S5cr5DUyNJfwe3PSdg3y9Jkb2q7TqLxCrHFBpSNjzfQbUgXXjYwXUcrXFvqr7tsNI7TbQdmzD0et
LL0yc1/OqIw4iVouEW/7Vf7GYifBrLgMiZSP30d5WoKbndw3KLlVhMHPeKZ/fFzboHpu0ztR2fBj
Brm570KGSpsSKMKrfKC+d/cwFqes6eXAb75Suk7AmLFyt5ZofszL/X4buBJ9UZhnyf98G8ONnTuA
1/94K5a+kLesM+QFH8muNqfRDx53RDx66M/mqBkVw4Apk+7CgjsQMWvTLGo45a6FPcI3pemSIBVH
+DeFYq3RG0f+ZCKmWLDS4GC96W2ysZhYptE6z3rtB8uK7WT6AY2fTxw8iMwzFrIeH38ie1uTStNt
F3Le1jA8itzQEbSrmQb0p+RSBVTo2aWY4IflpCRvdrzHlTCtrle2cuvEADR6IG2oaFkniEoY8nUX
RBip4SiGsjus6pLrtYGRi8G431XYZ5//up/6EXcaRHVKm8vVslooQUTneMWPJN4k5nwBqCJ4fdzi
YpDzYB6mu+cJvxrxUfsN7B1rh/FUzxveMUqXCwoaefKJ5adA3q3xpEfjR3cMfiWQU3uw4jjgibcC
ICX+kGEj13ZUjq9lExRpzqML4Vnav8F4VdL5r1MWne/9wzC/vNn0AcN5FjlbwAzCH71EOnyxyO7a
eLGvYv68JtTBROqidbAdObvJe48c1z6jLGW4LS9+U75u3EKtNC4WjtLdwqGHBPmj+j7bqVFDczAJ
IL9B+QKHVvK/TDvkoodhoqlfqCATfhj7TTqYCfCORHOzCznAZUDBTR5AILjhInXsqQaa4R6c8XMf
voo94cK7RAgz3rCSfU6DDVeIHSUII1UNvVkkVBFYmmS/qkrxrbAv6+ZiZcD6lNLjbvIvC0L+/kpj
4l/WnMwLDHqCDkvDI6m4atp5lgnsqFjBuetlsTki7CSvM1adJAKevqIPhEg2Cs+dpxcg2g3+/+yy
k3hBJdlARgGvfwSsKKxxuy+BrGjR2qkBNkGGqKwg2TelWxqmbjcLwN0aYltYMZ0Ll48ac/dlKDhz
r54PcKAAfzQiS5ylwokstXpDLjMIuzkbzIAolvTnpnTKxcN+/rYu5HVCzDrN/HC/msqZUmKqt8Mg
EtduGeDuP/zHaR21lXA++DjxPvWRNx6tKpUa84zhk/kj4B7Up1Z150i2AaWeUgbB1KxRFWANPDPL
kwHrXtE+ucgIqbmKl513WJufpEKIbV39SjjoWS6SLI0KpyCSUe48++a2Dbai3Dn5yxfy/hFgbfxY
A3f7iClTDm1jgNr7e/M3MzAw1aFbnYkZVgnupLWGvwSupH8wv3OELh+cGJivg8g7z7Xs7VAnlc1o
Afx55ygt+m3I7vF288EQ3KN6ib+6ZIgdBI9Hk733jv7J5I9j8Xk5lR0lDpPSjjjmlDdrt1Hw+IFH
qeVW/zI2NZAXJu2X6jgpSaUL9GIbrC8YZZijsDdlmLjBaWself9lYmxVnLJukTOLT/ElKGhDbtk5
QgSzyJo3wnRoZBbLQK4DUoya+6qYrQc7LpefMKzeRDtYcP6CAbi/uuxCy/2ctRS+7InaH+XKFXzY
uAWMdJY4GRS9JabhDQAcf1aYpXbqzU+Dw4QbQdDYX2YiPdAUQDRyWC3B8gTXsmpgpmhSOPxA8UOd
Xj1yBE5EmLJaauh3wFK0GVrsCAXYcD+JXpOZbipS7aYkHFsGIFQ8OlLkT4RcYZjrnu2G4PbylH+0
/+vSj/Q2BOFvHkUKrVD26l//lXopXyfcf6EO9HIWxCvGsfSwZTTFUSiJxEk20qSCZPjAMN/gw9AE
K5WE2IxYwlfXXtkDkpPn/xWO1oPJgcBL76zPd8WEYHvjsrJ6+qqC2S4vkX5+wwtqRPB/WEceUDOd
V0IrrDazhuFkEcNZ6DxI8fuypQRgafq3bGlb4cwSAajGTZLI/rzPhOn03F7eHjrWQHbO9yenpBOo
ivAutBM2n0ft0bgMrij9o9Pz0n/GjyFym5Sd5ujcQ/aUAe/ChkDEiXZDgJekNY9KwJNsnr9UrP8W
pO4M0M18r0H3h0JVaNuGgDEd5hNuWHTs6kEhzibMZJCfbODLfjJDQt31LNT0TY4ESrMpHMmEi/5U
FJ0Ce5dczKsI24ZkBTTtETsMvAa1wMwU3yASOh+9RxNE5nIHN0t9Hwg+Vckrfeu58C7ztDEhXR8l
OTh5AH/T7f0zPRlPrrRJUFA1yVL1SWi1gfl/ahrISH3YaJAd3Kz0tJ7siO+eSbpccMlp3Abpt94r
8qeDfuw57rmhBBDNkq0xkuXR/3j3AiO8x52V2JEHfZoWBhz0y1wwMnq1IfatCnZQgzP7SaVaBX6k
JMQfdnzUEj+SnhOVm5/8nidvxH5UVPWYhbpIgFvMFg9NTqaAmIyCDW/rA2eVIvDiOjE0bjBFksIi
vn9P6HO2YA6JBAWGggRaHQyNlJuY3LGR3INLhnrGxvodq2uhcSVc0u3/GxQ/Nqx7zk8jR2R++V3O
XHkyk1MtgWKjmD15o+jYo8kqbyAYlBUh6ZGa/cyALqmM2pnkWGLetyVYSVJHYY3opwKrQ3+qqaNd
kHzLjWC0C3oNMtm7LvR8Bh48wGru4r0VOhgQTrQ/UVuRUimoZoCzuC5X4jkL4uI6+oQ8eVxPRi/I
Zdh75lt8OKe4SUo5Zy83qHvj5W4I4bWi4x9Wb9UsrwuaDFl4VNfwKYaTn/81gGZYs24xe1GHHOTK
7SLvpVjtvGhJyLF5UT+bSePfiJYh7CdrYqUvW4IQmlNVfHB8Jcl/owfJ7duQfFw4o+GkrqJQoTkn
feSLmIy0Ija+wA4FPU7NlYUyv2x9crsC4KGXFCxfeoIaBToRg48W5xg6RAXuHEvHHU8Y6VMZ47xh
J6BtUV0F9k3T+6DZHUU5T3Er9wT02fb/ZzeKQdAts23riHtfjD/cdcmz5dFHEywqec1BReiTKnmx
9lkeff9vSr4UIeK2/2HX9hWiMzeCMfnp6YYLIlfD2CMr0i38PfxjIQCIe/Fs+6DicM2IWA1ec8JI
I3tM+uDgqz6llUY8/LHzSFkvcQ9N5QW9H2D4wNgM5892yby3y8G6jq3WUx6gvLWfO3HosdiMYLGm
qo3wDs5aQRehJkdc5KCRxYxKY9DozeeyARyTSYeu4w1wiCvd7Jm+K8etWYiX1phSqqhmVaF8gqR2
PGokdJX7fPtComJiyjB+nlpUSwsuKWNcCIdhSyKrpsZIq6VCjy44dwwaLptVBUxb0jPYI2iENSub
3Yw7PIJFYPK6lvJCCjPflCvopIajt+CO0TvMUbgQczwUnEnVNWbnyaTBYz6lZsLwlIJ34pM71b6B
/7O7egYVfRYlmKSDj23NtNoERMfUo9uMNartJOJWosN5eqMkZI28ZJX1cIJygkt/CeoDuexdpYJI
jl3vnOTdb1tzP4CJ/N3vt9/fUueVoXAs8wd6Uzs16tBGlf4VH3KtE7jNQEae7eWNAfdzmjm0WJId
GXRFaLoygKcvErgq7yJp+tfpqtyorATMHuthOfDt64nQ6qDSOX/uvAqoakN8v8MbbxdUi2L+a1cY
kGSbFUyqtWFPQqfcsc02KE+q7+iCHUHBLW/WtWV5hnxentk6Zd4m5G1i6vxeNCTFBYMJbJVGSJgk
7wF8LhY3MFegcLcd2TpJJ+kNILSWs2+k/3JQ3+ilFCbuQf5JPN8QvocdbsMEIm/aRHsx/QJOmDHi
nbBvEfZ4byyk1pT0PoX0NazKlP4wGtGy5dFXwkwY4S3MuFSsFvYmb9yCJSmHMkyCXiGG4MxhhLTW
tz6+KZpAmfpLp87XRIS55eDZRJgLNeRv/4fXE4MgLaxvEC+2oBR4vCLUKhdWJZsJy1NH7t7kzPZI
LssiMI7dDq9ozfif3fmUGnUU0swt604DwOTI5vQEf+nx9byonaFbbmE/vE45O9i+Rja1rtqsBNTx
qaP4pkn8TBweyGpsYT/wO3vGk9XzHlT9a+Om6TdK8ft/c/DuXldwIxlHy6HLXm6YG2bYD01fqYcI
hEfyezHqZIt728jogqzTPFNbOOpnTN3B9G3MTn+SEpdtXAd2MD9nGzQ62Q71JAHRfOcAw6+aR8hJ
XcW8oOBNplgmyLSKIGS8MUs3p+uY3icdXuSBLxot27i/lIuSm2hoxEFkwawuIhQZFIZQ2T9jk4h3
xW/LhbPsp9DuE6QZ+iGe+q9Q2w3P3K4i5B3/kExosRTlF8FHLTuqGQqvu+R+OcFeGI4eGAGC60jU
AuuXLcrilO6Pf2M7EkzqYZWnWpAdD/VXANG74nunb1HLr0UdCYG39GDv+rMHHDSixQ1i5z/aRXJT
I4Jp4CdjW7LGlGyUfOHby1PSqHqfmXi98/omDHClbCRi8oqENJ0B73uJnLAHhkO6baLtyXP8kK57
v/mWYku1xJezOVWCVai2iYmi2rQpKgXEIgcwJ7WqtNCYIBNLc5S1/FDVlS4xNQYakfyUvNBkx2ba
ugneAqKLbeor75xPpJtfnIBuRchtc+V6jTkGyng4IQ6adFnjAiC3KNd0bodBev2hllgI/IB0kyC2
DmtgZ0ehkKKah1dTfARUXFwW4pXBVIYXNSG28oRb14uYe7h0+2/AeTq0aFjowYEoTtTaD62IGzUV
yTh+TSAeKfre0OL2VarcGjat1zfXJvxtyloAJBeMvOViT/QhLJe+VucZ8Lvs/3dKfXCIF4uzCl+3
UEl5jBD1jkZ7bdP0tSIHs0BqKCnaePSzSFlK7jg99B3hkoSHA8TIGO/BXTYu9gruSs8mKG9tcQMy
AGiam3+wi1ASpdfZaxENoLO2aSucDHsVtM3GxGJn4z0+q5kk85PAm6Wex7Bp6PFYRTai/kiUNc2b
FbFBdLkpba/nJSHqqpFnM3jfQIyUEWkg1xVbIz2O6m7WycwjUvphce9MQg6l4GtcwshrZiU5/9dc
TlR1QflRrEkShmI8RguV5C1bubFLsHFcKDc8LNYrJSIrPB2Z3ym4L9/aWeWCmdTdETejdluHu/Yt
HrsLQfXF3wq8wdVnSreLW/TzBXZYlDE+CLTRudw6MiiJRU9Qm/5eV9ZiU1trZvk4Fsy92DG7BoiB
7WZnpsAk/OGyIUlX0MYHFKix1TRRgWRVmlppLLlSAdIoUyzh9kGCfzI4fplnH67YTGwO+lrA1KuF
FSbDQ+3hxfN5I1TzRCMKMcsii5bGoFBdrv3UOd2+pbvV9osFWEzpZh2rNNo0j8lzjnJlD22deGzt
/Eg/pZqSU8jdozoYiDbAMvWbjhWoEsGB4kE1EC68llQjFqlxpU730Qs3q62VNqp7Duo7iKeElZIC
TgdMfBFIPUG9or5I5TWQ1GOyRO0nx/xB9o6Y7Ttbk0nUabpiot86qKzzKgkUl7rUMdYFdqxlBs+O
94WvDdQxnsmJJSYSM/5a833vnA+C9Sm6M/AwoF95g2PBQBaP8SFWbSLxzNf/VPLL++GqP7r4Ija7
MNd/g3AphJ7njXxuX4HAoC06r5FLMmm2dGEG31WxpBLNE7PVz1MV3uDTN1bko0CQDc99AhLSXUfF
M9RlD0jk7KNR21RLrPr14KcNUOOWSlOacBruJodkfDInaO1VDdtXqyoQWkjPHVgTGHyjidTX+Yhj
Dyw1ZCFOZwu5neeAdCIonQWjb+MZmzE9zoFrFehKCPVcw+edrjRW3Xanct3C+B3Wcb2ch3Agj9wx
M2Xj6ozyp5OYGSvO8AZFFDQ25+ArDw==
`protect end_protected

