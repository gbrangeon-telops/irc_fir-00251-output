

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qCd+mYB+5ZYTiHGVPy4TJGVU+1xhFKOwciEzku8LKPbRfJOghBFppfv5cFbq1oB+i1BSYIHhjBHe
eBlHNZ1Z7Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U42W2uzowOkwk+UQGZB3li5Wu+ZZMdyVhWtZ56tkrk6iW89qDlhJBbms676mTh2iLt20rMAIN2QI
nrgBsluV4yEsobcfFOejzkUO7m425YrH0cSwookeI2lEA6QsTIAcBHaB/5shcOjOwrXurevqKKI1
D75XL20Mu1iceA3triU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Nn+1VEi9KmQsJsZi+aKtcGLlFmSquXhfukwVLZNoicIm0aMjF4ddZCMvsg6rFcVwB/qfiEbWhQta
pSDRK+xrjxFlcTBesAmRjUBiW3/wICtAFebLqkLpSTW2uzkYDkrpfNE5IjiANv3SGir2AFafH3k0
HfjDFe0WiziIlRflhOF0bV/y0LPPvcdBpjP9raAJY0w7hoeg+e9PIbHp/PMxlJRxsOwGTLR7XK0o
em6r0lXpVib2l0JQy4vnsZ8th3GiX0bt/UuR0caCktJupeOBsRztdB3gkPhiKQLg0696Wa/3XX9l
8h+H5UXqQy9EN5D0ZK0mIS8tAdwDRw6O0hbAiA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2LRSSTguNLx2WvUvcdH5BTmA+6dHxBZj3mWZxmBysCd90ElOkYpPTP1RgJPbqjpN9tofDDFDarkq
+qbG4SV9hnaX8iB79Zk1+LwdXefyq97462WHnxaG3I/Bff3hJd5X0rJVBnbVgHIqHzt/V8g0jC8o
7m7eoWRXpC5NpNek3W8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MM8YGg7IvNumb+k802doh47T9OSqo/qSgWEpWTgYva1SqSP4phIChk0ewsR6o7XTxZAD05syyzDH
Qfzl5t+Blxw1Jl5F2WrihR2G4uVbXDgvFSouhPopV4gzzwlFtcYs8jnovuVf94AiRDosYHN8WPZW
68LlNRF7Ti2drGO+AuUCHhYE6L1qXzzHwb4c9QJYmemT5/44a67UOyG5CnTiIpfQTpVHSTGdVMr6
z6vPgkB/8JeX7+R+UD1AQWqiV2w63od+aHRP7gt7KRL+kgJ6qCMGiaLr3Wj2C9mfPy61ebJocomY
5wy3s56g63xqQQnm665jsZbjTUelVxQyQI2r1g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9984)
`protect data_block
eR2+Z2EOGYmrPdJlOg4PiPNI/09I9EpaCDBSZkFdTjPI2jz86SMFOSM/xuXQffnHizN9nWiET1Np
cmeSU6CtBJg+127bw23eANtXcw1958EJ7xm4dsLj758Fn0abnXLug6UO225nBekqEZ30QH6hN154
MtusNp7AqpdJ6cd2wUgZ+shHaca2dksDpE34Ci7Z7dhQU4w9UwC7Je/cOwW6NCnvTQRG0Q6prFt8
vc7lgzL//KVCXz711bGU5mon29SlRCMHWPodfxIg1Hf+Tlr3g42gvPDi/hjkGzN/Hugzb/2Gy8Xw
KBwgC6KCuYWMb/ojmUJHnNl3g/KWWsqu+0gVr7msfFARYjQch7mpO7z0Q7f1QYQsLZqwH7lrvvZb
eUZVDUwL5y47Bau77rA7ZTnGs1qJmsurhZNRKKModCvobDnmhA6DCU1xUb7D5NyTHEsz6ZYAaCVB
aYFzwy4t2hI+Cvcrm7mDqnvCDoC/OFEHkea5PeBhqjtmzr47NH+e6NUEQV6n/gjMUgzzbvNmrtc1
cbfAO5dOCmQfYtSnO6wHAQORG1/E6HIu3ya2AM3iOJFYqrnv/slM7/9QwlHras9lek8cW5hqF2On
rXmc/SL9lRRNFOeZe6GvezrBzXIj8T+e6JUHLHn+NItG8IJ7mydn/wIHUrwi3DehaZiMVA8hMmRW
x9Jow9lO3OQaxc1ALH0PiO1JHJkGdVmy2me64XZoE2RfjNbRBGonoIe1QXWd0EVPyNvgQfRXKs35
lP12xcS7nSYpttdzwryBvqdPd2QizW3MZt+agR9XrqlvxRz5VgJBvRkVgrTbgNVH1Z5Zcs587qbW
YrY/z08+hmJSmEZH0XNjHAPK59JbgJeMLqdY2JEvPRAI9SrZdQUX0oRUvM5X5SmwxmUpzpaAxmkm
KBBVhQy4HlGi+AxMBzaKGYXCBzlC2OgeP/R+MBISSvpoQ03RPwydL7Sb1+rvS2zo3kkZGNr+KhMT
zU2Pn4/FkU6cNcukOgYQexB5EkFWdDxJ+UXafr40LS4Lakit4My43Xec746z0qjuML5QATFOF4O1
XcA4VU7yayax/oJW1wQI7hIDa3UArpufnmNKW87u9R5vDUJ3zAvy4q825B8wOKYmH15yNPejYmKt
32SqOxXpbRRalLNQhHTsAy+hwDcaFtYjN74r9C+gBCtwS+YKbPpo0Vdh1cJP9O3D7PtGciZDtBSX
eYaS5D3MgwK4j/wrHlBQdtV+HqZLz4O5lFEbLJYY9pt56fhDNS1wDFyy10mQaRN51Z5K2lOEjwZ8
dGbLO10teV6EGjKplxGZk9RE/6JMq72cujV7lwH0FPWfPqYdjFSWnoJyowouL1WxQQR2d/7tXd0x
9MdmwmlDcx3nKEdf47LE4UaE8jgv5vmdY+dgbmXK1O53aos0512zE3uZgHffWhTwD+3N70RcTK72
a3pwTZ7QKtW0eaU0zDsrHgqLAuQwUyHBcgTiy5QmiHu5tmUqAxKX0uyJMDE5a+vlm3DOU9kigZXR
O1ag2PInAZRVsr1V8K+YzPHJnXBbQpM/gXB3hndbTqafCPZKNHhRxlwQfBBt8oeqYCKmoe0ZmJKc
X3iX6db+Z11P1AO0hQQ4vrRZRDs1V0m63xr+DGJZ5nTovhg9mHpvlFBmI8AZvLXaWg8P622FMTtw
ZQMxhE7Z0iqfNaG4I3pTc3GzsjOZdGm8KpOOnzn3M9dnPYIRKlcSk1c8I2dxAdwpJEJPCYIIKhKP
Om3H7uFcluIKGtqjEmh6hwYEx1Pb8Suen3G3QtA9WzhV5HzChh8dqVP1AzcA0QVhaNAwfvKP4faC
Vx+v/RaaSLVlQ14XH+AKM1oTZA20rDxK5rY6QJgQ7q5yx8XOd1929Rg+fRiuZps4pzASZBl7LXd4
tshCzdY7i8GcNTPgWrtWSkCzMHGgtiorfUHJ2wgY2lLupsA8uxGNhvzEDnhDzBMkahKP3LDqnAt7
MiQT2EbccpE70BA5hMfo64OriOX6DnYLYndAJ15YsJaZ//Xqh8jjEtxd9C9AidgbDPn7bFTDFtqB
5Y4M2dq3frP7NqEjplsA0mL7VU4tzV3Q7MOV3B3FKvpOuSZlqC5a2THENcEdZfV9NPP5cTCotIWp
h/1f8kWxvILDLLhu8wV1QTLSxy4BWCUHoW9bpJUkBB/G4h4fOZpb9kEhNTi1eGqbZ8F9n/shl4sN
bOnsnk5Sht2aiXrFcMAoEZQWqVKK3TuhDXrp4VcbGcmcRnPXNqkSV4U5V7lrImqOlq7Z8tgFs0rU
a3NCgBazwUyXIOoIsb6JU0OZ08SlYwjPn4YSn9Q80URRAHXDh1Hn9ptUURO6Qu7K42ATcB05CA7Z
U0zC3vfuzEb4T3yRn4q6lXqBp8hmKZ044MwiR3oSLxfyphtOKYNSNXizs7GJCSVRxPFyIyhipkIG
/O2K0h8lftqH1v8HDC8CyS1g01MoHfA018UbzDbU30HeftTV7/LZVFwraKG/+i4r5/w9Gl82jy/B
ly/xQvVnZSOgd1Lll+NpwE8PhezzqFiVna8znKOpQYAx9VQ3VHzuQY4RoI92NKmCpJbmBBTvwLTX
UQQB333PnzDsMy/cpiT6TR06fNY/n0oEWQKMbm5QtGslUavGpE9Ep+KufKZ8NCVK8x6hdTbUhKBy
0cJtk7FoUE5tO0cKB8nKRrc+p8K7yGQBFvEJfoVWqcTF/9NRsnG0QC5DDwCOgI9n/Aw/G3hEyj6e
AdLNsuIltYpkuzWDrrSpGZXy+xiKjsrBO5racG1JreuDOKf0m/cMnO8180Wjc2k+RIWgIUv6lVkM
gMQLfvNl8zvs8H1p2FlAT+7dUZzvn4419x4gqtLH1A9EPVnxC7R6Pm4dvcq5DdxA5ddFAj4LVI8z
OwcZjGGhh7B3iuTG7jJIYzYY7xCM7O4Y+Z3Mn5M2U8Rxk1mbWMcPiftDWh2vyfQ1wrB2jQ8Sjo2M
OH+Jb58Y+4mOWdgB/7j9Lrufd4P0TF8dB6a3fuDtV0Xdv916vFJbyQ4Ko0OKVNhlQ4PJh63TIFkS
s6/+czwEUw4v3+hGZ5b1YPMdGMK4aQSETfv5v8flOGwZj5EM2uLvUxj9pTyIuPa0je9mbowPqiZQ
MBdEp7jAXi9Dk5Rn5W4gLHPruRbVSovxrXSz/1B2Q4X3N/woBYpHU1NlPlQNagIoAnKasEszgOyJ
3ZmErmeGoSEX6htJDjqctpmTILO66xjq3X11jjxUHUMryreuizEJls+7aSvtdCKxY8T4uzyuqFRO
3OqVOwGWA/cf4HeFAgIO5+geaSJoq1Bb2tTf3WhOyphDccsZgg4ZihGLxLC0oOllDS6ytVAqZjZV
eoFFnv4Ork2quPLyF+bu9j3Ve1ARkdr0F8Ohg3dn7U916f3HSOjQtVM/QUhdetkQoRHY81fq2jqU
DtN1mZMaiTFQumwTobiN7FZ6+XAg3nR1qDR7pmxQne5tE2eV1KEanC5xJIy6aS42kTKGaKql7iWa
B9oc8nruhuAksAvUmkcP8KSEss774LIG8SW9w2uxTIfhZpLwnJPtdwUjNFIbopqUu7gq1lg2iPNV
mWPNoYIue+rpDrF+qzFs4TGxYpCwR6tj6Q7lh6OV5PRjAaH00h7Pcf5T+5USiuustokgIFWwOCdw
y82LvQgCZ6dFN6mq1NSin9CLnAz65XC4wOHPrhCn0z3h+smpjOjB69NCrjKtov87cUhge5mVuqj0
qXuhZR5/1P6Ov0Cb1/I5EKoDlEw60c1/eMaiUbirsznPMqqEBdgzKKc/TeCcgrKU9Sr510vz8Yaw
bR7EVb0SRbUimh1SdRs0gvb1TRSHlL2BARD/geqo2gGetjiucVuJU2diOEX3HZL17ioLqYfvbBC3
W0OQBDJx5mLCxgy0hcDVYQTuO1I94myi5nbwb/TIEtgN55mcfJuy5ppK8YFYSSQ8he+NwVgWUVxx
lW7+QuZ/x2nxO2Wa4xzE415Dull8j3+GAMViZhiwjLKAtpFyWjU5CsQ4P5XsGhJ3eG0vAn0L/Ehc
kx8HR7wry1WjLIt03p673RssRinvO+M+T3us5eu3OvOwkvXny3f9HmcrBndvxRPaa7xbaO6fgKHk
JLv1bJXPSHEzLebRISPN3K3TIAMY1KOypSi/U8SEopKvIyMujp217EydXUqX8SYUgpy0CYaVKwnc
HWXh701dqp2x/O2VUzj8kOK6wrNPIpTUcILt8j9FtLggTmm0k4ofg9awGDQ/kc9cHL1+DQ3A6XmJ
jA9dZ2Qnb4R1szEWg6Un/XEK+Y6LkVQdXJRoE2OpmBX9EP4iSSuUBXht14O85dHIFUHY6rh9UWRu
EClFYLsa4JYl8VbdwPnyZeP8C9FqBFqCJeS0RKhYX2Y/plO9XH//IxBjL9LYZ/RDBYUWWkBrVEW6
byBtoT7LFyAOFurMvRpSpJ7aL6gX3BPJ/7CDgJAjyQ3RftUosIdNYjPaqFOKJwtf2PeLlymsBqJF
xdVaKvBOPU9Kd2b8h/Fk0oPfZpgDIK+bXhEB5ZY1/NtSw83SQ8INpgq8RYLCZ3HTmvjhk/deB4yg
X1b0Pm34Y123B1OpThDM6dR+7YgSbQmqYi78Nup/vSHmDFWTcd8cYgUc92pDMSH1eBUzToVfTyZS
eNOX+3MucGO0027MXRCnGVr3aqZdZidIAaXmG/cO9aO2h4Q9WAbal0NhzfaWAP7QJbAMVh+lGQ1j
izpZ2jzM4r1mEIEbNLBRo2ZsYoLb8Q/AITl6MFjVSEiFBEuGiG69V8QhSkLXpk/eXC0T6fZ/g/oq
1B7YbsoV9h8LBmQhZvN03PrFDbZ2Gr3Ek5WZXnZod4dGE/cgJjIhOR31iv/WggagJ7nLV85Wyq88
pvJVEcCsckwa9uUYGyRhVckl+aJXBuEvuCG11oO6o/v9me/XItcE4jm3BMnH+1XkdaXOWwCYLgbq
qyIBkg0DcdqO8fbOXVU3WNt7JOBJXZxqgUdgwLn6TiAoiDGad47RRxs1Nury1Z1SKDVhw+1S/0oF
BLiKVKjbB60mkVOXxcMyCFQsu3hsj9bwBrC0KvPMyWbfg6PZO6AqSetAHgvuxwICXZUAxWmMRtAK
pXU0fXtDzdroBIFkTL2lTsE47EePKpbW55s7DcS97g4p1cKV/rZy4+Km9IsN/pvKxsq97AiASRT1
M7/JLG8th4zzAEdKlDyAnw+ktF5uf+XU1XW6Ft+E2461fMLFgos9iPe3xK13FG8nfnVPY4LN8uUY
xrJAk49ewr6hjMtgihMxfhuZX1LiYMvRfq8r4nzusoT5nbue1qY5tMUBrBr4dhFOJGOi9S5Crzb5
saKg2/+wU2s+Ft2CF+ogonJrcFzI0Eyqg5QckthvpC9aHiEV5nuGMaQIhAOHR8Kp0By8YNWxG95L
1heorR9qXYZNExixxu1lHJ8wZ82EA9sffkZlqiDgaIpDnmR+UXL7eOE0W+OS+fDb1CKAJWXWiTqC
hplrQiren3nYpkDu1h+eey8hKIshNXhtermdp92OIgw7cyd8U5ULIUakQrudKKfl1HLqVhS2E5lp
/sAlQ9KEqDe7VQYSlYglN0bWNYr5T+yb7Kk/0M4C36pq6Bpb+Zy/OOsmU+bNPwqDC4ASoN56zyKo
NtXHIOcjtPt1V7LvoBsrFrrEVTFdRPQNFZQ3Uaq0Hp0iAZDOdGpJD1ZtoHwAZklGVeM9m5BlZqfg
KTo2XyWF2lkWu+72eehFm7/clndUqH1Q+25dXNBd6Fx85az3e41DPQnlHTOPV3nZEy7EAYw+Vp+B
X2svoca8FCUEtbfOQw3rUodIK4R+EOfvCvcH/2aGmE8x9B125LNYX/cMh6dSfxGJAbZQ2HKasD9v
yMTafvjZ1ODYpadVaNvp8simhmzwNRPnKgMECH/4YK/YkK9OcGrPHKLeoF7HdQ96tlMsfRH0Q/Ic
Rj0Z2tPsPcXoPi73zk0P5CrY469zleQi1UAANzvH5l2j+ViKu1moOJoUdz4Y8MmScbRxkkRGGpQz
UZRwMUD6vWJLIlBULGb9hqNrz0dQmzGxtxOqUPfRf/3YVgqwfF+Y8qg5Ep81R4/p4LG2+vfh2+q3
T415lb2igIY+ytD2ahzXp+g6UKaziouAbxNFLdWv1akUCnFc4rh6NgUpR+9qNydWgF5XsdIScmPl
H0tEEsAoUiyufvUVh0QJnsqSMh7FvHkvGE9W62vZcznDkfHczF7tN1mRDbPt1P1FDEvgjWnt6mJE
PPhZrjog9jFqCEZZGfjC80su1hnrzjjF5/Fji2Q+vsD6KRQOCmUzl+eOmVz2F6OHjWXduXbEHHqx
CLXT0pdOkSvDfkf1J0VVLRpuKVa9ds6uY9I6whsZJ/pwZmQAZLjCq6NI7xcQCF92G1TA5t+9SGx+
ZiX5tePTHZJffYJSGF6sV9LwhSkLiOgDvOtbTeGGNce8lPbI7hz7ghTgTeUBHskxPinriYoQAIez
YafDLh8fncnvZf9a+2ASvarZuzPWtSYPMgPQ+arsaAGRk9C3IHNHlVa4ABysZqCuyQQrDsQRFcvf
eVMXjA3sVp96e5SoaR/3hU2/0SrZnQPhA1MXc1xxHTCOJvqAke4erivmZWbu41Hwi6ocnw2qr3hp
XHoHceZ9YE7dG7tJt76Nl7AlOg3303Fp2HZ0Vlu2AtkwtcWO4MK7kF3gWRjqwB+y2fkOjhAoIric
YP6oRSR7C0kQVoFQ/t/X77wKcvmYu2QLL3yx5n0Y2phi8Zy8mz/4O013OymMWCS+9Ikz0YfKd2kg
jpXgfTspvAK3DBBeyy97zKREh1sZV06HVGX5iMLoeKX1RDdzf+3vuIVUOvY0zsEL/hrfzqjPURz4
8QQ0hktoL5OsxmJNUz1I3gGnPTTHHH566K779No7P2p7eCNQluUmBX8d3vFn6ktduVtrcrWQHHfV
dqaBZWDy3nyVOLBlZE5Ql/reioo1xBNmCUKJ6TG5Tbwr3Thba1CHgycKHYBwPD6YqMb3r+z7Fgvz
Jv7ntKXL24tYZ6LLr3d0liqhWbSqWibOwkBuZKlspYT3FdyMH7L2TPhGz3dM4viXsZjZlUnnsZCb
JBW6rLjZPnvekf46adJyPGu1DCHqpDNk3DRDRs8ZoJt9zGmNK4OwwG8AGtukVTudRVhpcp6o3vaA
czE16RXtqGx8t/nWJ/L27XJ9BhsxcHdiHKl4BZ8sGJzIJYieV7hVBmyddUvBKfV6xbV9Ug5HXhH4
HNrW56werB1kTdwsRLmaV3PyQsNdVs059gAwNW1nLXp00Hu5wIPvgt1jCMNIoh1GKtsfNCwexwWP
blOLAtHjI22Wzow4Xkp/fXBvdAWEUeE0RQpmZ5WkErJkDsT9qkbxsbBiCsttu+StaeO3n0EwIooV
y8fGgUjTD7i4kX7E0WVkliFBKQThb9nazH4+s7Y5jc7YqI/2kEdzhMGoBtma7QtNFlVcDsoy2WES
7vMTe2R3xCd9rrdkxUmQrYI+0XKt3zra0byrJxsVyXDjqFUxc7pn0UW9lOpXARzbl5YZqwmIXPH6
Lg9eCnzICs2qwruhZdfXXDFXnEhPFglnqQZRHJQIO3wXCC7nJ1bx3D7NPZjoaeM9meb6P7PPQ/px
eHvldESya35EbW60JzLWEzDRgPBL5pKnw3qmJlXZqXtTcwbd8x646tAtihtU3bAL2DuC8xmkCTmt
pBH+Sltoz7mepvGRdm4VMBr7D6gquBTagzsvTGmeSb5awLALJd5FO8EtFGhQULFKuH1KVlxv72TW
zfoRJt0c/P90vov8gIolzqm4/sgJBHCtjGIq/lEsuGEg+xUXB7k388nd/A9KIOt/7ywuGK9sB/VT
rN12nswOFQMiQKm70IzIKyexKzCDClyfOqzHHLC+ye94ydZV9Ms1vJp6g4QC+EK3uReSbQJJ1cGt
q4e46qFDPr+bTSSzW6hgEMKsSaPa7RlxJgKDwakew+FdHm92klil5TQDvlRnTCw0zW3GZzKwjMqr
fPjPlnFB5J2TnfFQZsENN28OWjLAlXPq4Qn42fY+HaXmbouzrbfn22dlwnDWPVtyivCggOKwihTN
gj+6Reyvq2uBMwzM4Xbq1U2wFNIYMtgKVBer3BjAUY5fp4B4gQS5Wt89EUHGxFwMozmtjh6sdxBb
P8X5XUdJC3qj6fVWbL0iHo0cUY1CfysegGe5LsSxgf/LzKGd1Me6qic6UKaNKC/qTxME6m3S/XGM
fONzwMB3L8KHQbtbjYQGHzKalxPF5lJyGspT/OmSUKrFQxEwltCJlNI/LLfmrciIhGxvCvhf+TYt
rquFK5PnGLN954SFpd/TPOSaoMgvBPIH7gM24W6VpATXw78JdrXa+Az3FUUMHa9mgFaPOt9p9+yV
pVyfC2QY6phK1Ugy6KGMS/KkmGQ176+3nvUo4YUuWUzkC+D+iqbC0P/7wQ8JB93byuOyRzTfw7LB
yzjfVrruFgljbz/0dm3ThFwXILBzlngVjUEceP5LBUVVOf6nG8xGwOox69YOysq9esPsOQry4Nrm
ZAqv38Mf5hK0MMe25CUaa3G/7KsC553L8iLux+Gx2SQ1D0clfyXmi6j0C0YpGfKFiV9/8yaYGnvI
AyN9J3N67cj+Qd+4fbmDOHcIEzccnmwaFRpaaTSYyindJnk0EThhj0ZnHWEH+e+GxwMtDfayOnio
f2ylLoEJGOtHgGAiQAMhgb4hg2MPL9OyLlP/7mP54mNmo1vxf3dCsqTxiZ9d6BQe9x9DXrhsfgsw
JTnFHDbNUZFMd/6IW+78SgvTi7q+5EEtAQShCN2iLUw8pVQT2VLeZ3PWl/j/i8mhlPEZsN7EbbL/
SMOYsATsQ5ygryyF2yZA1K2nUfgF86p1NGSRvUhbwq6TCJ17QpFdMXKkTS9ukQf4hESdOK5kFwkR
o2/+6Jw+ObUOrflnEgfF9bMTX9SJbkW03Zd3YMWSEmeuFZpRgDP9E/9J4DYLRu0t1Ah+NNSJ4isf
//5NNsqLCHKaQQv2s0FOOJZ969EymzR1Ocv6PKLw/Sue6wNCUlEmZ9Ph3z7KMdy1+KdZCUAS1DEv
nSL4qxy7Ufwak4wax5anoLtUYJAhkqSxPGaer1coOFC5d/OTGR+g2PWMCHTO/snj3eZpZ5iegvca
PKi1c40w4gv6i9C5V6j8VL3XxMLEkyXfsrezZj3zeiPIcJay5sHiNgfVXTTqzNipDJHdmuVgwhwc
ld9daQa2YVpsNnbzrlrgh2uDDtqp839d0JDYQ39CFUVKnA3pxqbBCMDbFovhgKEf+tugK93l9Hnx
yZUFG9pY/6vOC3rjExXml3jOtOqRDRVCWMxDhEwvHQkC+/8pHn2jmbnuuArgyOEADmLh4qNDbWAC
amYxwIx57BY6VheEOepzWYs7r3auFmAHJ6qIzgMFLsMF+9Vm+3i2SIRiy0MK/kLutCBxi1WSS9u4
H2bDWJYEZt71FaflCAUAqntO32AliysYeVzxbmRr6NfxAKHb3JNgD+b6KsL+cot2GPB33UR/72Tk
ZdIjhI7YTG7IqNrHxBWpEySOzQe6Vi3KHAWoBjNTlZoWy15gLYqZVSleIIPG1RxmOtr3MdQMsXhM
k/984cE46yOAw0MU4+Z0ElQs3dxAqJuaho5ovNvER+p2bpQKW4UVp9IAGewXWoGAgr5ZXuInUp0F
uBYGsXcFz0oGiWdvgf2YQWtjPzx+P+gANNAaCfZ9NTA0A1F12EBromePIMID/DSVZEWjK2cFLyp1
f3PctK0z8R9cplZpmLKeg0AqfuNdCP+mIrlhIPbUIaCFkNYX5htivIJyOpV62U97CPj55hAE0K30
5Ja0PC98EwD9as0+sKYIREvtZdJat2kR5YwdUzlVXxMr/g2xXQEyxUg9qA1GtPxiVIAL1Z6hK/mn
XlHvOAs7g+WMZ2V8z6kMtEmZEDBZGHPQXSDnD9MmBZcyNP/mBc3k7jcc7oP8uintWQj0dA3jNDEv
Wr3tZh9iNtuMiQmcWgiF2dd0uZhGwGGSzD5lwDMgP7+Zb+zeAxV9d9Lc+duOGqoRIdqcDWzO2YVr
TBFLSCPKeGOCkZg6lRNlWillnMguhl9ucYHrDUd30QWAYaAzkRTZ842Xg3wVgpfNDbELwNDvZqGA
ofUTM3drP1ao1Qu/0trCjA0ubpH940nS7/jW+92eJi4C8SUwaxRWBE6HNMYAw8VyurELlJ0IbYHS
RgxNrCfpGdLZV9EhIT+tsR6Uqiq/FOy7ZQLE6sYxVNfKCzJgB1BRLXUFsU5neR8Er88o0VbnMZ2k
di8JFznuH1jof0vQqqhRxevvUIXhVXH82XXExkcJh/ppv8kQ+lGId7BIP5KGYYE9TpGxEW36nEJz
iNuBhD0KN0iDdAI8K6MH1Fu4IylIiyXK6sElmtYlGRbkdzRrh9Y8AoGMlr7C7xHtxFlTpi6XvKY1
CUP5letoqe0Gvyhr6+TzxkiMbPwsNW6KS7E/PJtK3TK45alFWsuDLgkdHkY6tYD75OgDAs+etdKW
XWYzhRZ/pTFdG+h+1LoHXEeMLDeR/0Hg93ubw1UpUOBWO0GBXdEmZCOhb89IOMiyLo7s4cMGsLad
xaN8SBd1xTF762D1rIoNd8Gdu7rpDt2HPjf/XzAfcfIp5pXyWNKdBXjzWIzGNw7Z2Fsv+ZeZ9fO0
RvdWX4ntyrdJATgjIyxmSPnMFDs7DGLBEn62hCU5m3mQ6AWPIWu534tGNshcVM/zlMSdZRQ/zKIN
vSGJfdVejwP6eBfkILH5PbA5QPr5Sa1Fc1SkDXJ++S9NQ+2I6l4KBKgJw0i0HR3uiwNVOY0Hl5WC
UFl9UuCz268Y9Rnr/r6bZYMByuYNh+5688w9PcH9JBYo6qC77WehgMaLS9+ssr/Q7JI1d1KNWwsa
juX+88CnFf0nZcO6KHIXgX18vzhf9FtTd+anyC8hwa5b0bypv6+5Yl+IKmXfIZgPi7sBiFOQbZgi
CuXWr2mJMfqDGsY9tVvxJ27jUmXxnQRAe3yqOxHuTrq2kIc+3F2V5YfjwO2pOnLRSqLHnm7Gkfbd
Ha0t37k2sktJ5aA7yyFgayiuIpP1YZSb7umNQTL5Ht2UV814Kw1L1NdXaDe+DBuDkX+i7Axr0KSs
WDc5qHl91FI5ep3KR64CbrNDnhguK2t3QZgG4675X5wX3m4y7g+YqSa2bDteScy+4Pnat5ZbhvwD
jIsgKM1rhoahQ3jQPa6gwdt/YWFtidlcabGHlTWtRbkmqdkfsFiQuDX6BLqUxQKFtfTwmd/S5lpz
vRM8WpCFUpO+Mmt1ndXi5dLJf5slYQQr++r3vDpBiZ041rj3hgp43he5ym7fBiDN/koUMlMBdWeI
gAMt+JqKlweNtUiuvsSu3lhzcX77oP8hJbUd7bep9Geq7kM75b4bxeEoqbOZRCWadezUbl7Ivx4f
GKnNuLI/0iRnqwcyVJy1Hp4ee5fsPWJPiKUbxYcRlO0K8xx5YMTOpPG8/iauGAW3AhSl2NSA5uQt
/H0daQztUFJeuwbt8dNR+stDk1c8DchLC7uHcqbtuv1xK855SkHMtdFW3aGYY4rpws26CDpxkNel
jiNrAt2qiye7aamOPxmVphZln4pv8jfAyjlUFapQYEZMetZTcyrr8MI3zcTykVIz8qwSVxfeHgff
qVy7hehjSvW/jdCLXIJSzKKtHHbboCy3vKZBzYXuX3LIDwm4ko5S0+d++8jfuMo8Gg9iSmUcQae8
/UIPc7Tp/nzKD9uZeiuCMYLM2B/GZoXWjeMQcI5OUwFO5nQHFPgGd6sZHwXnPYsGtiGlR7WgArr9
xKE1/egUSZcoJKAbjCQEy1YWjU+88/U62yBjNCvVI55Y6Upui2sd6gvumO9wNyaqG84fyVqe4o/i
2p+8JD+wsPmU3QqbBQq1MGlDGCokG5EYXVzdFDbi2pLn1H4xZ+5EiRm226Z6jvlac2GHVmQvVHB7
MSNqSMf9aajllyENfZjqqILZgQS0W2Dw/+FAUCgJ0WeRq5RJe2h3xN6lVj+Z8H29eyGTDNKd0woB
kgZu966N98cjPxZAHUzpyIRsQNdAeZBmoAVBQ49XVYIm4LFGQpz6/iNNMYpNm5wHj2X41+eoaYCX
76QhC8HlGAjarmqetluxuqxKUTA8F4UrkhIseIIAwR25xRA/6zMK3CbGKu0lWqmZHRYmq6wg9Klo
H7EkqQ/2su+m9MMc2+xtHbJdwGZC5qxTK6saXxl8FEpj6TR8ZSowSOsoFO68CzQdtNgkBGv1XUzK
t4E1Iiec/ILLBqX0xWqziME31GCWY0iXMrRy+Gu5lpLPbC75cwkm1G/EAQ3Be9Bfpo1XT95p5FI1
+pHCAquPzdM6TJpb2eJamEZpJOWWlV4yLuaeKgX2QctihT4iNEi6r4rDqpWdlWlnVgWLUlJISmuD
1wEJxgc7HiakbBceTJmxYfHjFJkaEd5ZkZgkel2uu1HTd3VXBqEng2M551mRBVxwWETWbin17e4g
tI/dhT8Vh6yn9s4DLp8haCoBFXnm0VwrOfMI1R/VzKbjYJpctUp746V9UbbEMK0qZS6FBqzpkEej
+uj98HBgQwhACJRFtg3Wg8zrgS/9mzRv6y2BKPtfXLzg+QGOcV1zH70HRDIJ5AcvteptFAKPiO2Y
flW1NbENQTxBx/d/1HyHajPhF6d4ss/J3VwvsBS1I7+Pi27Guqusi4Z5qyj8QUTocVHpj18xSA83
4WTxtOdoXLWFocQMwgE0OYWuBi9t601RhUtTfO2MqIUc8eZmLPlJtWqQ3cCWueGfW4N9Q2652xWT
BKmERDodb2puBCBfRoNfIxkZxn9UB+3oqnjHYt1Cj2v+PiRAY/NRqZ22GRjc2W0TPYcaEYyHUKnQ
uAE9De3/cMfxuKcfoUVQasf+h5QSgq6ntNMrSOGuIU2dK+NvyhBxzInUMw7jvaA/31ceKT+wXg63
9eHtxnwKAb9FyqeGLtHAvApuHFVSGug4LRbHnIIiWpF1697GyrSgCCPOyFVpAET5tCD/adNu2cjq
YD1K3AzuXJsL/CDHYvk3+ljBes8nSOfBI8rD0gzMs25UwjPpiLSJn0RpC0RhkmuEpHSW3x7EaZN/
TpnGEiQ80YQNfy+wRK5YdC/Q5SI7YDJGNiGHNZ9FgyvsuasDanHdqdDICcUtD+K5D20BNxxi0g0i
p1AEzOmwkbPjOcV6sNuT2JVbDdI8Q6hCBr0LgChMGBfKfMqEtPXc5LfUdD0vSnBFo4TTHIlIqXp6
yz8HkuoMD5vQRvzUrSawd+zz/uQgUFMtJOVTrOQu+voqPYVKEhWT4NkuNPhotGBxS5Oo43+IO5gl
VWAhtKXXR69J
`protect end_protected

