

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T6wVkTPpNtKFC5HWYRGz1pDJeqROUhDmQQB0XOtYU+hhB43DLNvsfjC5KYqU6Qt1lGAhH0laXWbY
sFGsB/1X/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Bo87Ik/z3ZMfvsxWdQ0fNuP7YOCyp4j/ygqxg4KH1VshQEFmP82QDe0umsG5l9IQ7WJ1x44Z7hUv
b2TxMUXo+JqxKnlgUE5S7j3ulzSH7GuiH1ZZMyENkBX9PvYGPAoxkfBZKwYBwge7dC+ekfgtgSTi
JmblFBaQfl2z3igDjdI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OS69EpuOCXkwKDIJ7c3PBFNFMJbX4CiEZKRiPCWgGoIatev0sXIZ8vRiD53mj0pSkbBqScW3T3bf
nStSylNR1BolV0YoJstQyT1+2pFYhZ1LLXaZugJ/oBE6vqGV5u6J3W5eW2CILy6xHulOJT7cesIj
cRuZgsZzN/xmRcR/wqC0vFpdgeypXB6mda8Kpubf32Dxwqfu3L7BPiBg+o1IuskbZi2Weoc3I0l0
OeBzQzAzru491AqXGKlZ7sf8bs7SXbbzXRpVODRt7n1NjaKD5f39RasUxEkDN/Mf2io8pxFG53sn
wj8Vha0LEKNulGqvG45lCg9sffq+6YoB/PA6pA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0V7+weIw8dZ+BPWec3DOIbteiwGwG6dN9psrs14jYpdIBALSrfKIpNuQOkhxmutTucD037ovCmPT
7tzlCJSh8b8Ydyh2TEeIpJfXn05PGHs6Bho7YXv+uAmzXPPeMsLwL0Zdj9PYL8wHeM9h3s3oFmE0
whlOV2wA/y6g8Y9g2X8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LrKyoRzDm4cxDmM9WZQaVOeA1DZCMC2sBI/JOp2hUeVDZFMUfjL+9ejUV+oaV3PC9kYwU9gS2N4x
T5QckNj/uBm/MDZii4ZX6FRa6E86JES6LqHqCKy4pn+VjDJ9xeobjj2ApHw2GympzRIfTHfg3BzS
Zkqs9Cmo3/2Uv3zdNyaGnk9f0Ojhxe+EEq2njDvi1AWk3nuKPvaX2PFiQqvWXWef/JYb4HJ0Tjlo
v5y52n4XeymzBXqfaj2Y0hccYVFZ6YVhMnGGV06K68vVbtdbUuaSPRKXNa9qJHwvtspPluLhH5Xd
ujRGgNTtTMlfDYr0Fh/3k9HYg9NPc+b+y85sOQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4096)
`protect data_block
YaG5dq5HvTLS1MNsiDRvGqaMHWDRm9WUkWBjU63IeOaB84+NXPBMjwDpHeAGmK7bhhfrd4D+lOei
oNdbaDlCPfp8Kaejzc8hUY1T4BwipKkI7Y+K0YaRRW0d92TtrlO6WNul21MNkchYsnV60b5ZXDR5
HdyJ38TZmGYQKCoLOTU4PeSvQpEihm9R6JnO6xzA20iApQZ2bH7ammTkXtD2PxUf7eAetryu3Pbn
YNfrJyRO2HGqRmXqrdMZ0apdS7tMCmo93L+Pl9yuSxNebD/i4WsDJX67XigUuISJSp755uCUzlWd
Pv+U+iQhvuIVP/waWlhdbSdRbvC4RS1NPoCVBlG9QLshP7n/dFZU45i5Ug6kQdEGLH+LnvzHpjlk
h2e0gBjDdoAHJ+RQCLDAyBFN/s23PTRRCx3ldmkfE3QYpeQgcr3hDqoU/1+WE0UdhoGS+Y5yiX4O
MiXHYzC/sA1u9yutyILr26hYFppCm7UM/y/KXteKWgbf2OsKI62MxJoVX5+x3ZVNN/fv8Pse3PAM
K3aaJKVbwYUQUD+LqMejpGXvyuKlNDwGbr2ELfuzUqRV/FMdZ0dMIkjurLzT8Ygl/WCZa2qC+9c1
hjIpwmIfJ9lNKcfs6KMKQu5c3mfJ3jwysfgEySJZIa5IuWI1Dy6oXy8yvuHT8d694yqfKkCbj3IZ
tkXroAm+8Lo0GVBtvL9sEgsHhlWljIIEVfQ4U71+OlF26M1YNHnberYlo9BYV/mAwv0dwPWhVz6v
4JddCXFv8OBmIUeA4zvw9u4SrCU19QPkALSmWqqd28t9geRChyRK1VS+VEavlAqMvsEacoOHXh8f
lCsfRFL5XoHCVYfn6P/jofFUzXGAH8uJ0MF0CmnTIBjzaaGbvs8P/OCDt2Aq9ktFkNhGDoMs1P3M
kjMqp+EGkrLow3BPLtDXzHRMVDGcQPm9TtNGVSPUyXrWHbSU6SETqrh67CUT0ZLG78qK4U5tOY6A
aMe69eS14QbXiZ0xKtactldVNpFM5pR8DKAC0EL0ZIb9ax54vERZL+U1H4yEIt4EAlj+PzPSMNvx
Qbrv/yo11jplZGl4ZATb1yCwtQTglIQtf+eMfGwEPLhwSAV4iDZO7idsg1E1Rp/Gcjj1jKGpgPkx
xTaaDkGXDu+TTPDYO7rCpg3eAdRO6G9XamzsR/zCHhyzLUdEaf4BZqzimqF9WVYLa9Q92L7sAS7g
aQBbxUv3cHWA/VfqZJZDMXP3p5z6osgzw95HPZFxL6zMcOuQU/WtzXtjdzZZH9k/z/dJDDL9lx7j
470/GaJ9zJg3fn56ydToibmsKwiPyvlvAL95G5Emsj8OSNwHNazczdR8fkohNN0zm+AjfqzUpdqu
3OS3YYZNHbANBlf7+x7Ivb7UoYXSnJETvJkrdghXQNgk1iYU7f/fhEy9ZkcZyoF48p6NTEARjbz/
zLbnHgBFOvFqEdj01QkzvYKyn5ljQdedOQufdVGtXGw7Z2w8XJDxP6V230Iqzuow5vTIVcwOvycO
BgIrR8Jb8Bg1JmN38CZXYHcshmp4eJ77laQMEjwIZg13kJb+pzuOqGgiPLSkAt+PGWKqCdaXrwgS
lJ77qO+iGoD0X+f7njCToh0suxL7UOASO2N1HcNd+/Pk1dmiQLbX0FZ75eS9ZOMdatpSJNJgr9w0
utM5tX50bJD1LpksGzRatD2I9rNFcFOK9IGlC0/k72eI/2OAh21yJrrNwJN1ugEginryAbZ4Dhdc
0IqoHZ+BgeCumL3G8hDLXXaKtz/0nTC0e69y9cao2ZSU/jIJwOwSptsCfusatLoU1k5t2bRw7jcj
iTeqqt0Vtrbb7ebNjoX3y6Ksnxw873B+64NV497pPMy1PZd8vm4XJSUeWZrD8vlrNHGTH32EZ2oK
oWVNY+Imq0OI3v1Cnb0owxZKJMtzC6BKm225Z50zePrkK7XgTHLNpIqvPN0UpmDvnInbJgUPZ+3X
zFu0hb0LaOAEEbMuL0iAfrX/Ub3P2UVUiy2AtwN0jVOgLCk+RgkMsgFHdGGaeVFy2v+5wE497x79
9rZuHjnnRVcfBMlZ68MD0N5OLkWb/swJbvC1xsHY/TF4fJV8+qbTW5DG2TfrkzSbN1isoMuKw7Pn
N3iOPpr5HndqjmT6ybsM+vhZz45pOJGEggXMzxXjrlUcque0tKKADpTDM69j/Z+eCjfggb9kzk7j
nNkT8RgHNLDjbodBnkc3RNeIreL9iLl2rPnYjiRIwt+q6bTz5YB59Ug8Sb7za/HbB6Gj5gzG6qdv
9joc63mELncNl7V4298Uvu9O2vQa9w3I3vggUDsHwxRDSaVl/i/PcSu532uRJiQKWKkTNKd9ov9F
1gmRk8nivAQhmrDSEXsv2Wa/JTYc4YqTcHgXdgDhFczwV3ftMjqgAOe3kO+I3UzzCmfEL/BYfQMB
fsWRwuvJThj+OnoqvleRHvOYSpCSwYiIUDlYTIN+DO5mMrYX1zLtsS/YVUrhDBAQcbRqZqlDe96w
Sm5d/1UuHRNzwp4zWMcu7FFoQ/+YwKjo5tFrdk0LLJqchIewnmpWXHlSZhC88RXi/DZahZrwYAMA
RNR/zKkloIJJC2+vse7+V/EnFJzSWodQSNFBC6jm2Gs+ZDSEdeF7qFJAbv5OXL9SltjoSWGf9prb
Vij70Y/Y561WEude8AB5OnpD+6yn5zt0COLz80YeFj/stjKCNVQ8q4ZTqk/0kHZpXUIigmJiU172
SjNbrrEVBn6LWupnMJrngxtrSsDH6BRGq4fE04gkVwbnUBpTeMaNWPeU3xVjV7X/AmdQTFrrPQea
McpxyQX3opvARnLv4hC5cyIDiSPthjnqqZQIcPatR7SXqxIU6feBGTP8EzMKRolgJOHE9uBpTKXh
vle1vmcx5GEYt8jO6tu2NB9IzwlbxNZ4Azh4Bd/EmsnhzJCon/ePFutqODthsQsoDkBl/wj5U8Ap
PmWl8zfJ1sE4CR2QYsdEieSHVoPbvkejO0xMw8eGie9NbccqhCANq/LjsKLhROvcVh2ppA0b6esJ
SofDAMdyoqKmbqpSCjp/rzcpnzJX1bN/ZUFBq5ERNujEVoAeDePGl97ohp7zztXJm/7URFaEQtDK
r505bVA8VJbwEh7irc0SGaLOfUWQAez8MCMOiJu+0p5YIDzeLxRs/h0xfRtfMzfiYNhqS/4LQOw6
2xcoBuSkQQcTMBavqyGuIgpwc024DQPhlxdHqvKQEu2niQrLJ1yTURvX6YFjAce3UVpgxJkv/f8t
z6tthfbWH4seZapTmk0AC/RZTUXeTe7a/2gg0uq1NGeTFHrxJqnq5RBiWEhTZGZOxxwoNjfPnrQK
biHO+c+oOOYeZk+jo0HFb4TpKbSNQ8LvBSvxZys0xiJyB8wVRj6SDFobgzPHGVoTWQfy/fiVpr1R
rwaYswrHFMcrpcGcZFzXAhg2PdibkSTmR0A9XL1lV1QgZWYNPRZOlcx7Z9gtGHzR+RGrrhFjHcAH
PH9mn1CyQ+U1W8dCd6L6vj61OKOFIB2n4pVG9qD046xICg9k0aYEImBtVPg4oWYPSgODxijl2+zi
wR4/SHzWyD84Cj1HgNcmm8ziNfDhBPqAd9WRNo18X/P7WsgObrqigmoNpsLx7SuzQqdoq33k4i6X
2xLptLHnl53gHT0K+PKgRN2tFeFr7Sw40hcK+HChEh0rSYWPE+MCMy2313a6kBt/vJgH5JljGhR5
ud3977Io2VKJPc7grr2wbl+aJwEIWuNF2yxc4uTr1exz4vuPh3dHY4cnPDNoHTiWlqC9sFwoodrY
Gzz/hUKD3uW0YYMVkMtNqR25LYMZm3JWv/Bh9BFANbpqCbdt4k0JDGN/pDoOLkVtcWVtVY3fIu7u
DiqaCoUEo9eVPJWYJTzHvKl2qIixhAZ6Ex1UMFIE9PkXg59rm29Neqw5BPUkVWtpPaoyTJH+ijzI
UGT/YO7ldnQqptD/S8P+FY6eB2pFP1BCwjx1REChXcmD3GVdJ3nauiruxErHbssTmLqtSfgj4JuA
rw7Owc9xA+UN4yWFsI1DCH6DEdfSfn/3d1cn+EFG1knP7GN+Xp3M7BZvPviCxK2Wbq8Zepozu5EX
d9uQnZ5H95qN+dLrUtRvqwoZ+Nv3beNdnQEkRS8gGYqtiVg/mJaB7WgQ4yvPYHvxxhvgyc0s1c0L
JIKHoxNg1h9UIFmMQoRGIEMuu02qn7kaUF/SYSNoZ2SPkqxT9Bu2RmrEqrERaPO//KT/nHoByLJU
oJdDbNRbnIJW+DooKWiKjK5Q3dg6b6cFCNVGr8dqUuBknc9HokroGuxq1qQGhc/M+Oa4njlRDxMz
74zoxKuFg0eBVBbx/rB1dDbKXYLb8UUT4uBZqlq7mpLGE1Dy1E/7eNfWFzockmcm2M/zm4bBUFfw
DB69swEX4+Kj3SWc9NV4B6MIHREF7qBBnNVQTeXSoGopopW3Boxf9S2kAQtQKcBYHvzYj+QkygJ1
v/iQVlKuTxIQ7ceeUYJe+usFtqyqnb2BnJ7WWy8/0epe8jbjy3UO42lkGKxbPVQmOrNRdVYEzvTB
4KjAD798KH1SHpavXZb44Lq9hNlSQkcx7HdKptoSHjGsX2OXYcS+PYMtCe1rPfXMEqLbsBG8GF6V
OE+b0IHzVkMfTClZ8Y5fex6kZZZm43oXWcUkNDLiRDDXGIwywG6DOfkD1ucrjVCp2dVLMWSQkm/k
NRTIihrvvG+hyeAPYmAgRPdoTQZ4FdGpR5jCoS8YYoTIqAvG2dl+iD7JIGWNV/0K804PDXiymzYj
la6yx44aihF1pGoT9jYaC0xRozdDsPgNoZpoc3cGH1k5My4aNCRY1nXyp4qi77rXWG13vZ4luG1V
rL8SpK371opXUyrT6h+FF6ONjHeUKjlr8QCo3O0Dn/sKv+u48heQ0Ss6AMIgVZP14Rm2gZgZgZKW
YEupxTwPJebqhIJt8Ii/IK0yzH3/NiufsqExXTRykTvFhmldFerVdIeBLrOVS/nvD/SE4JFDsg57
qvrWkH8R+RFJHG9uTI6BQit9Ets/ibjuo0T462lsCuQ6mSo4pC9jp6Yv12LlRb1+7Mc51oGdAuV/
60it8ufbczOY6NR47PJ0zYSKY1kshnQdhhSvq7psKEgXUB96Uj4esYKeTNYl9JOLmG7OkfEYW2yV
cbqcFwkX7tPgCwGBR+qsyN7NA6mFk9orzXjk7T9Tk8U7hgJMCpSV/jxqu0PssbL5uB25F31zBgk9
khqrmbO9NFceG0vxePooxXAH9vW02IUIjycGy6/t3ZAMeMnfvLqdp9WU3e3x6AJ/ih2OWcGfzFdD
rH2Oihf2nHUj1Lkz9S7tEfHOgZPvdkh8MIchJzdKVWHDt7bBuJAZoQOZIr02AeX5eEeH7/tPqDlh
WCW3LONLlgzkUJe+gqLl+4zoif68bFn+RKZYUE0DCXQrkdxscCuGCKcvR+sBki/QBg==
`protect end_protected

