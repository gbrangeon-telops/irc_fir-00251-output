

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ya253+37kdInKtzN3pd3f0ykMvIJsSTHE2tRr5TaFzMStJPqyqbq8G0/aCj9umOixPoTbod1oPEi
NM8lNQufqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZnAl3olUb+r5fzAKtbT+P9BDg9y9NfOiCUm1R2Jcpt91ydHcXeu+pZ8D0lxHNM0CXXGhs5RFFeCB
fQNmyCQv4qniT4fHHC3wrH5hPwmAH8kqSEyGt3c0SvSsHCYTeXhpF8Chp2XvC1WNZGYymRNjehFn
t70d4j3zNeEsu5WAW84=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iKnL/TA899sfLGiFOsNtfsGv8lNgBNaSxC78jj2+skMz/TodvgTxrRQVQ/h/L38N/D5FIkKYR4II
+olODWgmPzea4VBkBMLQ7z2XenA/M8Uvin39meT5Qbx7/ksgG2EdpyOtsmAvmeXZQgf/A59DevU7
Mrm0rcVFwLpmjNvbnBOl5iGpGgx6v231GzIUzFEiOeCx1PkRai2IOZKE9lG2BMKHN7Bhsm6JH1NF
XhuV8OyupD6h/Fr6EDMMNZqriSBB1MM7btJKN6VC9jmTT/Bega2BSYjqAkfYdUTeyup0UqEM3znP
2BL1mUmUOgL1/UMAmExO5qz/A5ddH+Ai46kqhA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bwfblhQfYU7J4v01pOh0vYth2hZJ6Xlf2qmEYdxkErcnbM5+VpJUpwU8+A/bDOJB4gUPbJHCeAw+
tmj2AabGe4D0Pf/UukkjTsO8eFOUvoPbwDwH6UV1AKQFszUSN+Z4NTgaKs8pxWumW0juNgJujhCL
2ChBu6ddPnHdB5HG8uQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UTW+eKUNnZFWLDMo9paR505jK3kaKnyoN1JMPNm5SlY5iSmlguqsHIHMaqSHkHrYg25dIfFqsLa+
ygBhaN4bDhxyus3QZ9m0sw/aVS4ly/5bNlw+8ePaK1evrFFnRWDzqTt8U+H1O06G7NfpkTmeK+am
Q1esOyihSrmjwIiD3aw5SiSY1J84QcBDQl5D2DAd5uRtMADgrmEFzx9Y7yHel0j2iF6Z2vom7g5G
7K31eIbiTPvCntdYde5+aN/nl/kdiT8a+6o8fslm8ZFdkfMYbKE6CsL8CG+5F82TWbIzOMfxbILY
sXfUaKwgi3ZDGoeeudit9zXCRYxReIG0hfQ27Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64272)
`protect data_block
89kteF7qmSf9vb/ZM9yT0qaOyEQ4SLmvZbEl6YyFclxc5ZSTdkHSjA4qiA5Y3Jh4FqvNEemxdqsP
YgYh3wdQEgNj42+thGMx4YZkYy03hHjUq4pSbiMd1UfquOKC0vIhGlgLX36ukANHWeoNmCMk+y70
j2R3tS9W2PfWI7hI2Ly78tWcOQCIYM75yLaPs0B0SDxCfbEtcQcBLnRCg0ZZGD1Q4q9h/VSSHgVM
FisribOrHjIw4SV7q1moLvP2SLMfCxhkXkuBOYOAZvzBVFVFAWC/y0oG0DWxkMZ/FGFgJx3jthej
+L1LoHsCO6CX6VlWhix5u/UAElIru0swf9uFm58M26lFlgHpf5ybCwql0btczgPBJ5DDrRyN8Ou4
nmq4Qq1bcoNVaIBQ4R379NaPAecVvk9x7TAZBhy84b+FavkdcO84G1ZezukiEuvbUDLKx9RgZS00
3kTifUFsQy77JLBIrF2HbYiw7hnqHULpF6LSYqnWrrlXUkGVvETtRWLu8jNCAsZV9rwyZBEOEasa
+b9n2zGSuCgCVZiSTh0FMk+AZV8N4RbLnC+frgMTRKs3IMo70B4UJJsTlC1Fa6zliP+Z2JmJ5KLV
1zioH4BdlYyB5dawTM/Ynnkvsr6/8W9jtTKAlg2fybVv7J/SYqFobzLZJvOaH891+xOym7aTvmzd
faZ7T0AGLc6As2cUqW91Ap04BXL8gkfsoL3BTO0McW1hwpwD1gUhXmjxNBG4wZiIXdWxAR0K40aG
1MutE45Cy/5nbD3oEHH5xgIZ33EhYeKnZXWjlB8xBAEuwmo/bHCYghkM4Zt8xE0wfzvOHGfub9Lj
Mgm1EyusZH9jDtGHf935ZeNISGygxrHx1PPyI5BMPUgJN6EnxSG8tHvI1zhQfPv8csUbU5q5KhWY
WgY4af8jdSK4t/+yKkOQn3EVqAz/l2FZxMtJTgnOtu+tQVVwMUErdKMGLLed1whrMSrH+QMKKTgP
3Cr/AbOpji8bccBPNOOBsa6lYZF/7rPbl7dLkEG4KeLNS+yR6/IAUPx9sLjnEfXhnfuAVI8RFqxk
n5feFYjjbAeqskzPlkZr/1dEhdhZK86finunIJ2s1qKiLXTNDYz3d3qMslqS9lGnYSt7LbHT9B/5
L3uxpq7yGU7J6ru38VvSlkDN+NsD46bddc59Z3cVeFDF6hcHFB5KDQwZ+t24Br/0af0X9daf1CGR
OZ9kNLzu3Xyw5/BirdA/QXO8bCxa8dtAVwXU0q7XtBUq40cX9S6A/JFerj9TakIb31WPoszpQbsj
dKz1ge2Xa7vTLA3eFCb8AprBTMpJmVKURollLhV/E1rNBGQECdYiyZUFh2kM2szttfrtVZh7K83y
7ajThzuHiDbFLWK7E9HGagRVNc286i/7GN5X5YSiZfOJq3EnkWGHG5j8K+egNFE6+5y4wOfuKuI/
v8dkZXyWv+7c7imZsgluhxuqSAOeVh7UwrROx+vBCdKY4qdlWMHB3z2gUU+BYhrKhGzm+9KInkIQ
4Jb+WA1r6D4SZ+wbTE4ebKNMpjQEh33vgz2SaoGYwe2+f1YwTTehCLLYZP69xQDxWxpMZUpasv+v
Vgvw/P6cm1T241SUx9HORlUfVZWEcFldtVuloggLc2YTADvJuHR+LdTPZPop4xADpJ7BMS0HXxk2
xQt/YSUBrIKGZHhANSVBuXChBk3jieZ2krOhHSaXz3YfUegJr553W/zfSA4pMLIRniquwpCjXdwu
o6ELOgRvd/ABghOR/Ukhul7dYnWPBdHI6F2pOYaL9HEDBUotndEofYa4taWUINSgW9xbpuCOYZS7
JPSGcmsHHDezOj0zstibbw3TQaAHjXogYcjVSE0206OIHalRT1CMgZlEAgMisfH4WnfdjATUfUHV
JoekQoKFeRqBkITbi/XBoOpFXv2hTbCcanqtYeN39DeS3QR8mYheGHihcRdIAp5v7Jq9MWTjKqn3
o2HISa5N6gkmcxSSwqYmcQZr9cvbGPvKO3+UesdnP54aXD2LC1o2+HpOyxBDImAbHuyXAC7g06kL
xFx6QbwVBpOm9IiUcr5KDf8PXTuz1TUsP3ABaA+b0V9ERWMmuB/Rfx7RqndOYNVOCTbnqBkBvziM
feXLlgdwCnu1Yuosn7YgmtMGxmCsgT8meuSIoR0JLzw6Fkg3Jz2vqHQxSrc7RARs7fw3B6H+BMr0
GN0I4jyBFpAjrjDdi9FV6AEmPCsAOypfiZfNfpw4Hs6Cbw5Om7G5nFqrzKiqyjLK55sY6nTx78VU
gOlgz8DGza1J92qLeTpDuA7colp+/tP1zygai+4ybwNNdShTc1r6Lxbyu8gGlRh+JV9N2wdxfmSP
hy2Ji5y5HOumiWwan9y+FtWVKDPPMOJH05t6KSWpMREf5bNJJ76wPjItFmNQBp+ryDepm6QytIJ1
dSn8hRL072ul+9NOTFQ0Z/ilVJWoPvQw4SO+z1ERcCOUmaE/jZfzRTTWOAoXs+AtmNLBayEiC1DX
SlG6+Z0XSvBTPBSN+YeLDuNVg6iSb2w0PGqSLT8Am9yUyikZ6C+DxNnHrEd63e2xAmd1ORsJlHPG
jjSTZXrE21HlXthr61hwDebXlrFEZOI0jVK+yM+d4TpBHks62Ria/hzj/sNthZC35iCV7TA1gyfK
A84q4GSs/9XX47IzmscenFT13pp4I6eR40iK0yXzMfqKIrY3AaBadQFq701uagWJDN3d3uLXjA4f
nFrLM5sGZ8SJN+voEY9wvXLS6CiavoxFyf+SW3T5wzUQ/1e1pGZaqEGq/RT8HNWngQqkUTY8qZjo
L/s813GHGZhDEQYx5h0tCmYUMAGQd1/akzaML6/Fa6B80G8tqo8BWp8Bf/iEjgXRHysS+KMQe9zk
0uyOa/NBFGfaMICP+DLfTjcw5udTdwljYFThtKGspvByE91lSsCcavuSS9u4HYInmnqQNiUR6LdD
G3ozMds7kjNGWGVcz+phnVInODoihjKyiRmWVO/06bMsfj3IqpACOosxetB7nMDLw7Z5GIXQQe15
a2KAUbDt3TYChhmQbVNre1Jm0tR3BGqG1FBz8o61FDmgQlXtzMScJ9Ux5q4dB6er3PO5Y1XWwMn3
9zQxBAyky5dPBtrgCAi8WBKlMkOQUH5lQkasTYSGU/fgd2LUG4y/MK7fXBS5zdqlY23cEbH0BYfU
T9Ght3qKnXjCF3IkauRPpb1HaMLpFy8f4smBLGoGP/OMgustq3RqUC1TzcDVRDLQDDZBswWIMKXK
fPg3yYmYuC0KYOixOXA6rFIgROUmLaXxssXLop3N22tFlsWoqNVYccVWGgeASdhXKi19QpSNXMrJ
V4WEmeLpcwiB5G5xxSNV/ZI+sAht/72hk+RHXvIkRs2OJicL1n4Zvf4Pjr2+IBFG6MgwXgOlgn/C
8DMlHYzlELkInBNPgFx77dXpOEEQBQOy6jwos+2s0y9C8G9mPycmR8aH/rwXPLES8dkv5qPGpT27
AYIy507OnIQh4llE2i8yDFqYGzcqeL1WkiGMUNxcdYOlNdcgD7mvlio1+lwiFMlAtxRTYq+FDWk/
qEV/ux5hupVICqkErQDyBkWZ7/ubdtOLlf7oPpL4ZhdtPPncl7WYEHkciEZrNVeUKYxpgTq/0jma
WNzKHUlNNkp4tNqAFwJGAU1paca0KM4QCOepPK9oO3H/zCVUlB8lfubzDDEhXNY29+zGxpzEJFCL
syONMD+5J4cEWBv+KJelDwLP0aRZPFi4oNPL574DYEWeKSM7qMOMhBsYcLucyjTX3KPISjs5N/rn
n0HOcXfZMBVgyiOXsobo8Tj1tiqa454vuTGXc4IL3m4LPFN9PEbyvoFeSxWhPTvLFianX+PTRpwm
gC4gsCCbtgKBMqvbqyog1g1gr6JpFeJWEl9PKYL8sOcbie5xnTaXAdZzP7aVlHheuLe8XM8vqxUY
/GFOjwBKhWI17xVXrYBcQgqdBE3fYz8QL4rZiKFXrOJE+EHBYJvhqfwenB6sz2braHlsm9u9lon7
t0NWEYcZOGdPUvaR4GCg7F5dVcIOdVnU7N1Jf5azURAnadZKkiAuSevMCNZrWhhESXfkXST8us+p
GyJOopIXznt/GHWqqkLuhrlLLyBFE/ZYVOTAgJH1kKHHEtke1T/3z8J9O9mxt6m5HU+lhOmB6Pnd
G3d/apPiSr5dNxKf0KUorAF3Aq8Xq0gNhzRChKBO/Y+dsWCr1fNVDdG5OK3JJ4o0tOws+P9mgMVJ
oNVaBTBhZuKX9ycQlYyN7WC2jwHHQh86E0EZIs1W3IuhGvZXUH0PtnA07TQz2I3CfED7v/p5LLuS
OTnsvrUoQd2luH6P268EScM9fhNZoEZeTfcgtiopwlLWv5ao8QVOlSp+R13VcDHp++sDXmwmTXsn
ppA4332h6N9/ANE0aMUbhl3277zKNeXrUoxJPIh1BNIXbbnSwEhXxvsHW6OvDt3C6SfLeFUoPWS3
x/FYBbKFg+O1uU4Ck7wtB0TtwccOdQIqJtDshDDkbT/apW/rAjefU8J2z3jDEQ8rDwGB0geBE2nU
HMhkwAnfdVEY4EUlwuGtv/MuJDZ1m50V8EnGRZSPohJXlzeDDPtabVhLkcH0AQMFSDDgDy6d94rp
3xPZesmdq1qiE2ALcQep6MhPyZeEX2fcVd88xz0/+uxMWb943fUaXo+F20lj6BqqJuSbH+Z5isHb
m9OtapV8wk94MzT+aInexA/zLUdQFdN1/HS6vnrPQ9+XPjqSf66UqwlH5v0XRrSJ+5hMViAc3mfT
/RkNZC2IK6zGSNmkNKc3jc0/eG8QiCDrMSgjEwgbvJwxppjRP+QokfGxUZzP3GqHSkp9V9AojECB
7n3rImDZnE9LBcrrXZwVTnHIgBtK+gbT4XNI3yIDlJZ6wfVHXp2EnfmlA3Op/+sM9rN6Xmqirk83
Wu4xZlMWEW8TWKt2yn8I8G33PbZtORZalaq+oNuiw+fTob/2Egf+AV9wjABd+kx8p+EdfHz+UTQo
VJmjKGR9JGGZt+W4CU5OZnrwGHwZDpqSw0Vf6/Jycy3WGQQaZePWB5yZdUBXqMoNOA9RSfYF1cgK
SNH6ah7978y2nsCxMA9oumWjVKRraKE3Yw1QfIUpk4EVOCxJb8BzDqGXeM8yCRyVCnxlDFaI1AnM
uImuCHpUQi6NlqoNmykjJtzEU+U5KFJJOU1Gkmz1u2MVxwq7WRB7inplOiZm/WTZYhNtaqx8C7Dt
VF5PYv/4t3eGA3mxdi49NYDV8AM5hjO9hwQ3WEq+1NbYwhRFA4zBRAcpJtQ9Nclxht+T0ojlswdM
ggIqkEr4X+kYhjI4V+wRw6Gpw09venpiTzDGm90K2D/J8kriWL8oECf0ezYlksCzG/1ZKh8KZ1nA
z8AWdg34iJDtG09BkNPhQf16T9nEs8+VIkcEyoaSBng+oesUValYAatfogDw3L2nf2fj6eIvKrWO
+nhwrrxRpTEQJUL9Ga9VDOZnbs1O7+TQ++RXavgkv8qy57OmkrWGWDhOhHBhPnfVWyRmFezDk1Uh
UtZcJEN+ZIBYmEvhJ+TCN+SKvbo60mLkGSoZlIN7fIPtbwFQqtmJW+VRzndop9TJomUs9CMMDyj3
ofDgkqUMwD6ln5dknPUI9xfA1dCgl+a8JAvNr6DZfzxj4O+TNM+qnEXAeVjkwG+dRgmev1VgJhq/
Hq/OEjcWuKV7P2XYjUAjstJxqBPYUooDZzb5OMsd79zNBXH+zLRvDYrx1GiLyW7Uv4UZyJxeAG0O
Qem2cmc1UnpDWheJcRg5OohK+Yfo1xikm9dFsvAuTLsiM72slFSoVKS2/elnn6VJZJbtPTrMHECL
qqFB2sJ0glPgemrxT8K0OM9EemUSQVL8iiuSY9R1yVIqU8wMZKQEJ480MQQG5PVpLADkHc7qvY4C
X46zbjYz+6KX59DznJCkcj1DDm4lqQAMJp+FSt8Ii7xEDrSKvsAPNc4wnK/wWSPzIJljw/Qouj2s
28rSQIDALIwVFLzORd1T9+sp0BgTEfAWkk0g/uIlsyz5bID8X4NcawFB+3cuA/AvU2y/HawkBaZ3
yDOmYtmiiT+GrQhap3bUyybEt61dYbO4LpiSAnNkClrgt0shBH/TGlHXdtjCRrLTT0fULBSVkgKa
v6CNcC6hcIrleH1HLGBEvAouRJRpT/n5PBVnzqy1cAEA4bnARSlNzG7Yza5gwKJhozVW10FWLPKg
UPl3ftfpSkowSeWEm7RBzMVbiXyluYOENRww2RQFIvZMYWFn2gMm9OYJdHwQVU2WKWojIcSqoZ9t
P+4wNuS7rvDxSLWOzYZhlN/4EVCuSGjGYngjR0DhR+6zyG944PE5BF+qqM0+oLjl3CaRSFXMsTp8
0kZXGHeAKqVFPRw/AVxQ7O0ktRT01vCuQDr7Ha8ZlKCAo66VddvFYgRjzUJjHyyB1eF5bD9piYsx
CIZGuAcQ2DghIDopQLgHJhfnyIFyaAZ+8z0S4XndsnA+C8y2lP115K7FR6d5UX0XDBWCPCH7eRq0
41XjXD0mdSTYzZnqIwITtPSux8PTfXc8an0LHBSayJmRMlNA6ru41XYlx1kvjFnDwtvoyIN1+ijT
MfTqomNVBep9HvWJsHkeze0AMBO4Kg+Ro0o6yILCIU3ajnBOR9Keu4BcdwaHQNxpBd3d95cM9wTM
WPR4Zqkgy6ETwrR/YMxHpBTUkgQ35qnYvVUyoEmN4WXaUD5dInOn3AQINDLD8a8Z7NPGFX8js3LA
tnzjSbZYwt9w8ikuXJCl0uaiu7OkVFneoj7TYnjotGTSnoyO66mveicbTMqBpAEAM3JIxCOzEnum
7n+rd/YFBKVGbXelxJc4C5fn6t5YBYB+K7EC6/UfqYJaF6oUQCU+TnMiT3gb9dE5b9olp+OHo7CS
cJ2BoCHD6rDiw05d8AYUJTmqRta4GFRZ2Pi9ybmFw/tEU1MLqFWZYR4iwHEuqSXahAoQwuAy+RkM
2S9U3KyIbkCOXftW3eJLEmWzDBDSrhsgKExCmP1Wi8pSMtaTdKcDDA14QAA49dQ7dOqJkUcTMUny
fAKq3G/+sbg0F36p3Egf5m5XHhVBVRS25h0XLNNXSHcEh9vzC105CP8b1LfmD8+iXjkpyLNxfhOu
jfSFeLeM0ludTGp5RSHoJpUsIcvPeB/ljGA0Ma/ZQqelSwuyBMRvk/Om5q/87WDjMNIK0vvASyhh
HFhU4VoI2Tja4dKNH4+1J1U2JlR78duRLUZAauPQB90VcYG8neY8iih/fQ1cGRROhZAw/XgswRvN
ktJFjcEQcmCzLjGTz9k5N2YI6PyApTMZFQXevX0/bGpDlApAybSuNcsbCUGIFpH6aDacPk0MHwpS
tPLjb3rdSpzeOTADgmg5OeQV5ldJxV7GcrGpzoAvQh5apVZqkxvaY3rBJqi5MihNBtDZuh8KUoNq
8uxBsom011QYcI0+cA5x81ZpAe83eA/apDCnZwK7ffvPQLj683P5vS+zwuYayuiKVrkO3LSG2qeA
eohtEGWtdNgMKx0rf0TJzh1eDvbx4sQVb1RAnxL5SOP+BctQzDtbiUKqB6LRLyboq3wwK5liHgqo
QEu/VyFxuU0KjBKrBRnXikmJprSztisDMiGFZCvbcuEJZD29n3E8SJJoRIgV3jNRWy45KELodz5Y
FeccRr5vZqdIymMJoSv9f/jXljneK3x3389tocCwlxSFrFAzh/0dmoxup1eL32LhfUbZ8sFRlrYJ
+o93X2ZRhoReTSFYPa4JrQfRDEaaB9Yr8fj6S7VzosZi6bK3wg4S0PO3UVyNkIeHDMRuRB7zTAHD
K333BATxM/t2DCQOX3+6CHDP44op8w43/eQEcgGbgm0jfix9z/ARxRogAhlR3bJV8LRVGhTEyK6W
Td3bmyTPHezHfqZ1kHtBLETQX4fipk5HjRnNEiUOiwaLVFApYdJN7spHM/DajW3901/ULeAsp2/j
AypHquHR5zjhQ99B/6HrM/UtOrx12RF4jbxSM/f44K/0P2pinjAndJE1yLoVpCteLEjCONr1pQmd
uPShyd2BOy1RbXEzq3Ed5qiLGyVWpTG+l3/RR7K/f/bNd+GqOCCi5fwZ3tKpNVGS3RYQCELe1f4K
VL7b6nvrTk2yfSEzXjT5AYw55DHzw8DGTds79DtEIarStpdT77X0AgG+zIVZO32c33RENbnwElHk
5oHIYubzi2f/xVJDyZL0cQjaBS++4ZeztvXOXJUIjcCiM42Gk83wtp6S/aI9daOk53Oq3axITZjq
kzbuNdQasN1WHXfRXsEDkfD7bJRfDtomnk0rp3XJto1ci8gNXmTsH28yy2IQjdIJwql39OOzBfcM
OdU90L/UqxT32pEPse590YKmr9/53eMDMyYUhyG0zQJoF2fkKmkU9A+9OUzCk+K5ISK23Q/F94oN
ddDfThNSTsu8uIQDXwfdubSbpWO7lEbPxqVcLqI8Fob82RZhJYXV37bGhsN+ef5lYHLEBtzpUANV
rs1fWL9Dfmh2tEcUGFzYOmKGeEMeUeGvcKGAEhWutlWBrA2x0VFZqu85APxW0Z1Dnxr+w+0TPRd2
KG97SD8WO/zH04DowBA2h2XGr4eaNWee9OjLHhOhzdYUaWXjOqRuBzdfs3gZJ3ULvTESF51MGtv1
8EocLWZ+wPkspoXqGoIbyBSaQOh1uBmxll6/Rl9Vh33CdK9UJyBu/xbazEM90d7WCVsc6tlPa6of
xKcaWjdkF2cUNzsNE9F0ugq6EtU0m4VSdBMkrOppnPT3JhTHwqRBZ9Ga35q7gOaU7zeuuxF8XAAY
vDlv2MRE4lgHKtyWnlUNN5r0riuKHm+nR5vy1420/7sxBEvyoq85vpkWDEWU71POwuiZUfqqs03+
g+8Uy+/StbsHmLQm+F986he4xRcc8Gdg5uIoWv0P9I6UBdk093SA5Vx6Y3vG71Ak84fLKzVonUVD
38B6Xot8q0s0FpZQPl+Cva7vTCfJuCdk7+ukHDsSPhib5eV6Bb/KbGvKEI9FfdHtXXzfyyJZuHtF
Mbaf1rkFe43Xq2YFALZmKMogZwvlt91qXpLXql9LsfZHeaX1MTnoOkMzkUjmQK/5yk30trmAVVcT
KDAUUxYBt4Iv3UuZZiOIm/K5PoXXkBrn/7BgklCrZJM4tJZXsipftghigUsFG4iVIuRaBNvcYa1s
HCtCQndic5Z2sBHD2qIhuA452Zvp+PC8N/fbAtFama04syx+xMwXMJQ8Joyjt4FO0fIW1ZedBSjI
XbR+t4jFMVfMDcMHLs68c7hGRf/Qz21U4W6jScKm8oLdad85PPOHNmA74Kdn2mo3ZjUwcimziHdZ
sxurXSuaJIRwYXTQtxwOvG7MlZ25ZXX9X9SSkCyIZ/kZSQIPTSVAMMbuibKDxDhcVG+jCaJq2KQa
MSl2bdAqg6hQfp8SXyCszhzdsykBMZtmRhctmPzX3vZqoeSISbcfrzFA6PNyIOd3XYkJlEAfenlI
dCEwxgm+fMdTB9I5kCZtL953860KFGDL6l07qtZG6y7NvehrVwNeetkO8FMwD59rCpcO8Rrv0AlY
tyIhVM6hK9RrurtIkkvXlIgemt+QBfipVCFNgV0AvTDxotqpu/JYgmA9F2kBXBlmHGOzeEfI2rG+
7ztStruUdbuLpa1/izGvJAL73W+L5Ve/MRcKxffsJcdtR+cU38/OvIQEqD4fdq3NUK4scXAKdfS+
IDKi8mlYn6C4G1Hy+vap+91+OgsPPKZXR9Jg4SjYbhtfLv9MtiBAosUefAbAmGxJTKie/nXq68lF
UFqSoDuC7WklG7dhJEOnaMegUrBZ6JfQ7Fw4gvbfdpgXm3UlOHQPIzbrprphaCEgR7NxXxeZQl2Z
PtHoa08R3jbi2tXV6fdwK0+Wn7WBmzJ/hDIyMDNw1gGXXMElRqBuuey8LRSlTvh3JQavfHuQIYlY
kKUVmGivBezWzzD+oQe4O6eytN4dwX6asz/c4ULjuaxIEnlICyckMO7Td3GGXcm8qGlg3fFm3Y3K
vtIYq1b9xUSz9jxTqqWP9WU6gHr8pelzQRC19ywMWR7IF9YhTiyXkob8k0jtAjRaG1hUvj1DOm+N
+dNDLiaiC2UWMcvLd1r9U+rj59++AbNoJpLdR7OVJucQzI3wXLMcJ4kOcDcKOmZBiqAciQIJR8+f
FbsUgDF1L2spG43dgTaEWi3bXyuSSzVrph4P+p4iTNUAgGCce0nmnC1aij/9vCA3I2aCGZ45aSg+
dyJmLy4Wj9V5NOGn7O63NvS0XrsSiEM0MQr5HQG1b6rQhN2PkGPWx2QCO50W2Sh6DviDwDCfJc1J
NOJ2310eOjxLrB01tVEiSBowpe/NuZu1VbVYjcYKOGv2ExrDEpNOV+L8Tni2bpnVpFtOlGcb4Q+Y
aOaB6cLl6jTgbrftdA1iIkp6BjZrunQtMhGaWeHeZfA6CKYnjT4oPkIH/+2C31qAN8c/vnc5jjad
N6lhNVJnVvgoKa5kWM9EAoVZeaMmHi5wUd0Icht96b4Zk1ku1O2e/n8eOASEYfXy0Sja2I+91ySz
EUuGjwyMsDXJbd5t+gzwZH8Ud13kaFBFXfm3mWsUOcNs2m800WgZHGD4mGiT2SsemvkyyFvE3ikJ
TgXToCH+aKZ8GvqRMD98de5+t0ejAN8b6h9Kw8ZhueiruaBkHl6Kr3WRl7EWJZikq12ufg1izQlJ
OsUfasLVgsIYfNdp1Fe7Lo4Hq3Fj43/G18lcGFC3X6CSlBVzv8V3MZJrRV2lA/FQTVDEEWzptWDz
9NNNbLLhpsnZ04J989sAv6kTU/+OIKeieRwvB2Cq8X/r9ttjXxi8GOeGmHvGisGUZ48LdEU2vowV
oO+e1bLWV881WYK8imJOF5UYppRi2Y53/qOTZ4ts2By/fKsB2WY54pFTVJGtvqi++wpOMeXdZ5mF
y8DmgZd/WsyOEFaLWvAlj8MMfb07sBpCb21EV4afD+aq0A4mMsLl+GMCEvdMOsBa0Nv027icZQGh
RnylYLmBOL73mJnAQfK8q+RT7SMgwI1CsA7FPGmhfn1V6iBaMTXYEiwgBrTOyinBxAIZXRI3DjRW
MbNWksodqNtleekJq2zv5dp0rHvIRCu6Df2AhAsNfr3KHWXL50RERfZ39E8peLG0pZiWeESKn2eN
vubZevfQj0nxpIG5lHP6R0rZQ9dRBOF2+gMFhKHqIsLhad7UXR24zeP54uBztF1t9upiHTtTFPCv
CWqPUSzShPuarPlE6m6Hj9ew4okf3U7ykEdZ9g79y7f7C3ffAAdcl31NGnUl/7U3cNsZdwqWERjo
UUgfJ/F8OdwdJSVmtgiMbVjh7i7eUCBTJobR8TfJmFPiidrwoaTF5m91P+J7r2h+EeG8pcaZ7Zq+
NVHfBntgXS33UoO5b17AWaTruRx6Spn2v9ttEfdAnzwkekkBf5FdhlwLrwtf+UV5X6v1+7hJEsep
mNukl0FzbdgTY3MWHjYQ1sPdZytd21//JDujAavsBJ2Z3y2Ies0codGlDzTc2h2aM4E1yVHPqhKo
HDIRzQCnXcRSpR0yAfjLpxzl9rXCBy5xDSj8BMCQYrE7YRHwhJe0WbkBjDMl1fHftJNSP8hPTOoH
o3zZHct+kVmvq7Es2Z8mFNHxR13/T2o4vE1BZygOk+1WOv/L43FgLOLLLXRLIdsLT/WcJ5rsmhw0
2+B5u0zbR/NZcmLVtdNnNLRxCwJA7bg4J/JHTayvItJxY3htYzbZPatyZDJZk7llKM9Nqm2E+yS3
nLZTeirRbYHTo/8X8NipjB4Thf2y7T56P2C0NBZu8WBDCbQfdyCU9Bcb8vHXCadojNpYHlWMbAVU
kQb1DdKVj73lTS/MB0+P0iTesWW3+QO8OHpK6AN7EfnD+0cxRArpE/r/sLDeFGhA762WxFdfgl9d
yZvj1a9U9HtVX53nCXiEE53TZCMHiOvP3igDG6Y4Dw0E4nWFxbwcsN0l1A37HUHOREybNQLw6M60
kSqf+bLebRi+gDmUneutc32R1e2lqZpTUZ5QNl+b1g+s+d0DgPr0KEcThNW0usCm+dvVGnrqcTJq
5npG6tl7sAKYrnjJ40K+LvtC+axqEIHMpYi7/8vuWeI/3W9475BleJl4howhNPyKXr5jz5wY7HZK
oVkHxbO3asy6DYI1eswTjbEqiNoEuS5H4FSEv2deMxAozFJW5JZXQZl1m/Qe5pW5YrugiQrepcSQ
y5gSntN3a/bPmFsdVNkOKzxp2z8SGTFUhpo9Wu1iKr/AeKQnbnBH4hDJwarCnIIj9giNVJggpkEX
gDTBGtyPmInvAM7kvYxeRvmjUflP4pBEIG1ihHbMOPltP/iaw7GyDI9RlnkxATnlGdgg1BDti2/A
iBXWJ6XH69nW2VlACxypL7dbfQ2jqpwPBxsXbO2AP1+Xy692IbUE9NXs3hFzncgU6t3dsUDxhMXr
cWS63LcOL1WNfqbFWtHEzBd56xR4lairFvTqWdusR5X3sihJ2Ch+ylyFBVgAdI26xF3SINABBa/z
5X5i9NWrjUKwcJ6+R+Zxrb/2qq8PtsMsPUpnx3uvizM8a8L8M6Cfzq7mjVjzgUDasMPCAYCwrMBW
1bqYYX9zu/LU1XcTd6AuAy5JHNbPkU4YxndkwH5mJpycBHYaHA5S+D50p6r5T8aZJN9JduOFTp2g
b0nBP6O/rShDbuEzMqaV8lxpWEtbCEptgeAPWn9/Chvs4FEj88J8x3QKqfYdMYWmQmTTCyQYwOJr
pMwVpIyi+nMvYR5LaELknBjLEPXvCB+P6QukSqoRrZqfj7MKD6oMzUKbYhKJQNjcM6NhKgB3Av6+
muAuLcsryNIM7MZq2Jwdsa+KrNHS7B+fmbCQ1dFNgRHBYTsx/JPMti3OepH9s5w8X4O7yhKd9xC1
o/DF5TupU+36KD/wDqIBHcTW3+f9VqoOTmdRrYWbLT+boxjdWqbXVaentZ5MwrpE8egFqLA06wfL
tYz4k+yU0/Tb5gJKbCWtc+dM6c85rPdFr1YX8KRRctpqjVuzOYCX4IhREZ2NkgQ2p/iDmTJaiFFw
e5mVLFJO7kwCXHLVScvMOhjGFPCO2Bm4lij6tx1ila38WAUNIfwkEEZnWOEhUBt9mZkAqOHLB26q
+saKZx7bA0rXnxmQrboAIMQHu4Q/fU1m//nwQ+iOhxqQAM82pr8gqUdkpkpS7GGtqYy7gKCdFQjq
qtD6uLcq/O1s67zSqsEtmnVAa6iVLuzgANTtShbtwsuWDQQhrMFTGA6oVDUfznr0c1aj9kbfqSQZ
djxVjvqTZNUcKW/sw85+coYl1MbFmztsJU6FOhBrTkqtHezkvGUTi2IXvraLr93xvpd1X8JAQ5YY
rOynMqEj5XVm17C2Nf8hUQXK1gmCFk4AKkCpeeYDgBVxTVntaxn3V5H1PlZd+SDDJXUR2XNFN3Uv
gni00VY9Q4w0bhsw3Te371yAJvDCDiy74D9mFj8mn38JwJ9B/gfLK9d3YZCIFJ5UC1yaBSaE5380
Lo5mCkW88pKyF9KIHjuzZFj/n5x3f9gA4wjWIiPp3n13N/ogaLzBVcyWN0al7rVl9XDl/DMtepR6
iTljq3kCgY3GLFTst7/3JYq9K9jp2lmEAYPrRUY4PbvfgtpZ3rCsV6j2s8AanGFb4xBPvivLj78S
KyNe3x2LK12YOmqmd/oWcftawpMpzZcz6hoLByPS/+StrxkjALttq36t+JAm0LGu9PJtWY60rZgO
gBpK0XA52bNxm75rR4cyanjp5Nesbb1cQiZpVnwZvzS1zKmgKDEK69q6grm/iAOF0bzK//ssom3E
wtWv2DM1iHyvFqKTaEZnsP72Qqp0iPdbXnGPCs/SslOvDjUidN5qqrXPP5bUVNc/xes2AuCM3a26
HRKjQAe+DKF+3I+pYF/zlLbnvnXuWhfg8uxN7vUtl1EOvVOJAZ+tW9OK7++/BRlCRbJ75yxsZKhl
bWgCaIDr5x2s6Vqb3bSBftC/Wgg80PSehxW+Ye+ebuDAtZEP9xI/GyVx656CtKspeMh5hes6cZKe
fv1piBm3nxx9XWbcbdDjVjipQti5zXgwAHvY+YmynI0BZCJSV+Oql0o0slsoIjVEvvY8WN60Niq+
N4p18m68SayTjB0IFcw7Ctrj9+Gftin/IDGwsi/qBGYB1WdwnHo3Jss0O5EoyVwxKXp2gFWSBXFV
cToQ1Yai4jYwgubQscKZpG0HjjuzMEJWZUpHNOP3BQqLY+bvlBIWa3ws7/bstCjzn+W3WZVJi1vA
twqoELyLKHLgxI2urOetbp96REe2xV0AAeNtZH+Wl45EYIaFQHMb77WsSXd1mCGlx3LDaSs6uqzP
/2xo9J2f5T71jmdLT8vy7vdAgBkIiEJ45Nak25AVW1oCDYk2Eyn/aJU+vfcHXQ9jqBWWtgv0QBk4
ZEnKviGpUcz/VVHsNEGg4G3EhDsZWuTn0Vr5Osy2UnXqbqQ4w4IgGFi0qOVAfhELkJXtQjPi2ODj
SvjSK2XIqEyR90Th1TC7DB3QX8M5hPd5jz7YdeI4xb4z5BjFAGWtGwoKmghAhj5LC4NNOW7loBoA
0U5vzxzt3Tvh/xdu5gliKcYwzeJHHOD0zpsp0FrV5GHTZ5pUrlOjtmYc5Ysr4sUkyGXJnxZY8unl
Tkg4plLy6Y8queX8BnW1IB+sTETjNf//KPdkPQPcabVEeB9RIVXEHMf42QBHwqYiKF+2w39mZFLv
QDPWgx2jwxaBugNjg00ZtWK58NYVjERDdVUeYZiRUDCK4HBwsTu1R7WpqvuMNWvJfdQtw/zQa+W+
z9wrRhPL9BqW61HKvUoaB0ak5/e8GarMuu1s4qnHZR95+Qh5QHa8DVJky1AERQLXss1umeTGLGzF
CsQYed5Zf4Kx1bEYwOx0oniViPPqhCj3vLttObSUbmxO+XWbw86R6IjifTbeP0McpvJyEBOXA4S7
qHtP4XNvYn4A/SR0paFpCZ0Tepz38KDX+rJ70DAYOqRaito/AJB0LVGDahpN85zZmbsCbxIytIXu
6q5HPjZewLuNlGcLo5WeDvhsnwhj96d6nB8cdiLyD4CSrIJHNJmlnAE+acmA344JMfcpfbaehc+B
BPZQc9wEtLIHDwRCyr7gMpjEwphzieuZUqbMjyxc7ct3HxgtPOu6pEBs/g8ES73OQmEvwnRF5AFg
b1Ub60MflNkE2q5KHFHgTN4ihFs14uYWUSAvK0+DLN2W1gQruavVwd2ODzr0OM781ItLrw0CXetR
xD/+am38hikj/+Tx+qp2+uXsgadIJIY4n69lb7AWGQ/zmrp8ZqBWaLePr6RhMovoRAMkUyLPFiuU
DBzvbjfEIg+VSj9Mx1zOwQvEwn8WWQXtFX7bmSDWYyAhdNQtImAbJANLpAioehFniBmPW2blmVW5
/DzWMRrQF4Q77GIGc2RqIBal+O0wuJfa+lEhWsVZuOwajxo2T8LEv+m7r/2SVwfXnCfv2uiOSDHE
6harsTEk3IDPqZ1IP5OWnljkL2QgIrVKlWVIn5f7NZLTJatJxhJQF4woZi4E1TfHV0FafNITc2LP
Yhga2zrEiYIgnEB2M/V42X+Nhl8JkDkt+3lA8txAB7z2auXk1OG17jEK+KmjtTmmFKAktPyPu3O4
hV+nICs7SZPMetsEiC5hWEnSTIp8qQxAILidmC3kPbiyNu+kYnpCM1pwzYW1ZmeRZmompADsWFLJ
JCGApn+jOs+9/d+zd8g/9ry8A20YFzs/cueqwVNv600cLPynSGa+7RlTetdsKpEzvFNgRkMKRnn+
hr/pfy2W8d+HWn+o1pQkh0ebaM6tmtRRzb9yx8SVSk8Js0aLmjYUrw22xNeVly173CU/A2Y90ZuB
oOHpoeMToWnLlD91g3o4S7W60nvE9/pA4cSjccnXIEwKbEW/0zTerH5MBsC5LOhdNR1FK6RNxPn9
mvgGXwJHK214bG3bL89PdVcl20phA4mMH7rKHVnOGA5PE62WHXcTKVr1jCKKRyQw1j8UfV9ZOjhN
wFZt2YQyIpudBMDKt4RU6Fee/WqX1kK2upV01ixLJjR5hojruKyeNjv5CIXI++WpDl3bEM3K1yhC
g/XyZW+g5d9v4VSqnXjocRsKc7vETyzJEarhjeIb9DCdjlRTecvjcfsShJERg2TCjX4FxfQ2wIPZ
WFnG27UWBcJyhMlGmzdDbhh6FOydNuoL1f/3LFcPnCCbs5+s6PWKflhdjI4nR9JbVXasVbpydYdP
4IGL0rf11d2HfZbSvK52KA7vwcWh0WJdafpXLRhMYDsD5KiM8JkPldr19JeF6l/cPJx17WmR02km
TWOjNllV83ezYNnigE3vuy5Gbo1zMmnX+NZziAwImrvT6iIkq+hijmmb5JkplEQYZ6RJvaJDyKPF
a10RH9Gp/LqfeTsovf37rNXBwdQg1+CYkXFpusToxZoJ5GBiVay3Cf1i6bFu7/j2vI1kBfArDyP3
Llfp4NqKN4RsOjGFhnJnegAUrpE4tTGEmrEjjwGFYWNuP9jVBAI128u2+XGUvBaFIFSo+prCDLqu
mhMbEiI5nZFnP10ZNu/jLLgQp5htvp99TGvl5edMZcNrAB7wuGXUv4ImcKqzj7ZmcDJJQHbjHHUW
cbvR7ZCoBujOp2VBDgS1wv/f8KlzLnChTUkHnGfOmGNv8RcJkyHreblswad8ek39QlAhxgrWCPeV
ilSU6x+774Xjr7jWznzGZhJpDg+cFACVFVYaflMIE3a2uf4QcTzVvHfTtjAfctghr1v8n5aP384H
mGFA0pi6IIoBIlZhGTa70nYC4CTp9nLiREbenKuY+K5Rf3keiI6a2aKErJTAFott/wThU5GqRjxu
3ucALLdF+u1w+yXjn+3Mg1gm10lxim6zwIHvkwXZu1U446wff9Y9eXLFbcdX+t6tDa+0yj96dOSx
d0JMW8ZzOY+MuroCnURx1Vc4r/RcjLxLvaC3Plab6yXeMssasQ06CqakhEQSu2cDVtx3UC0pTy6V
28QQaS5XBCsCxYtTFCn0KJfdpTDXFvlxiiSQZqrlRWIy/TxTVqS0jsgMrtk40hZQcx+CCLdRb9lA
43CJ4yAO+8kEMLz1ZBa9ybyFe7RAIPEnr0u0S7nGZgjvMSrDVSRoMC3uQliQgoJmC3L+7ApewB9J
iWvKKGQwVk/dIbqVp0cEcoQeaPWhgWdJkoaaRmiTHbzNTmiWJJD0ClOCNRfLmIxblTTCD+ggd0XL
WIiVyMNdpFX4lO0iAjD6oIb3Zs831L7N6UL6e0n61dofTXpRSVsWSXIyw0QC5gn5WwQbRvuWWpZM
NNYZY3zGMRkgPOFylAKcuXCpd0zS75aVukzdwkPPCH4dD/LClfMDH+tswywsE9d5bTL0N4Ofb76j
7zUu9DpU75l7bwauJ/LBb8w75rIczBrkY1JQ28iqW/Pqz5L9BcU7gcXTSTXQk94yWT+ArM6CUkMh
FDwL6+rNN7mXBbHhY9TT/0KoC2FXvpAdksZxew1AxK2ptY2ey94cErxFizotqQ27202Dyvmg6mHe
XjVoWWUWLvz1GIVmmFPbd5+Q5GDBP/4e6OZ87HJrWcVv9ovJhnpgqqwnEq6G/O7oKKkfhjvrlM8W
W1E07gUzObY7A7wWfPiHNXJKeUH9McyV4/TRem4RSMNzybacD6RRULNM71KsmgCu30wER6xAmH1V
Dh+yajgiU8c1eyKtyGOTcP9inGgt320serA1xuL7peS0euPEwyXF6yYy0+M+KQRqA3h214LDYowT
2wvXLB21B/KWvDA+kr/i7wOUuycsYrwXuXdR8FjVk1OpTwfrSvDV86WpAEufqCHoGCGwmdulGGB9
VufSXnnNW66+u/OxARlYW+1TBQTARxok9gwNtNPORnzudnZRTaYVNAl8VZDLZx05tSHOQZ33F+Q/
YdU4C13/WhJi0NxKyxiA52OtKd/ogUiu2LHdT9w0JtJPt95syyKqHLZ9IyeZ7Mj3mSjpRexzpzGb
qn1M7+StOfdH4fWRU4St4tlJroJf2V3GDSsUX2JQzx/vdCdEKBeXNeT33pzg6CBF09ufLQTfJ9TE
cVDCt7dz88x2gWCZN76E/+Q+suuA/6toznAMPsscA4VL9uzL7iz+ScC8/L6HV+xGreFCkfLTMpUV
jpFfArq8zj4LPktDVw8ma08/yShDIIkBx6SEmfT/m+G6hOpsfBjqew7aBi50D3IwaCIedMY0NMTY
vPnUrUSu0v7GI7xkf8YChpFAQeGazTT9YOMoFY4787Cauh4jTSAmsuSbdnfZCvRZHuiAWXz2E17W
zTBg71c2nhnrEMRbcu6yw9DYyXt/ct66SZl73bs3kkXoyIFNRIzbKo9NhTSBrT2n4fbT1P3CRlXR
uaaogFUTFP7JREz23gJlOTuncpbSZOcKqmUjsvv+m8kvRxzy8LswkCDAMdmBw8pNCZlcxHa+yJxJ
g+UfgM5FPePlfJ1gEQV/FtyJlQH6hN8PXQ9uv5LnLd8VouopgfNCnsATXK8wYwDCZAryXZtevpV8
99TUZFkO6F5QTSWnkVXujUZbWVF9J/9Ft2Xg2FyGtCG7VJL+0SMkUUaaxm/IrOQ2dlIXdw3XwlhQ
ztgZprYZ7UE25zyyLx/ljp9rsJhCY6LoWbNs0e4FcPgmUEH9PuwjrVFAA9JOkylPppRVvk1UFDP6
HE+0PCeiGEJjDMOweGIg9G9xK8NBQl3qHhsZKkg8+xTejyiUKiranbrdXsaZzwALirMKPh3NDPXf
J2r6dOtM86bw+jnZCjy3PA8KRdr6MoFH3gxLI/X5eYtw+2EN/Rb81GeP1Y6kCBAJs7NykUqy0Xza
F/30Txqw2N6N7OXMb8/BNJsavGOhcOn/IegMRJHMDX9zA9nyD4I10EN6hH71tujMr+NbJmhK6Eqe
lHPvpkmi3+MFNpee6Sq/hg1ehnJVqaH3slZo/uGp6momrHjJNH663mozZ1l00uzDVB0LV1k5/jK7
3UalKY9hIhMXBZVQazh4T7sFgk92IRmD0c6U1+KzRJC6UKa4RBgY6/XSKyISPFxZTLPK5gtn7zJD
ZAVwZW81ZAgan77Rkz2dmvK/XGJ5SS/B6TuyrHgS7IW7XmstR4cmao6klMwymi/sCxiMOarmdYlg
enA1P+Nt0YCemmd67UluWg2F6sa8rolhFfQJg4BRYnY3hBlCaOSRZIjr4eXf4qa7aKDwYyV8PsMr
jGU6MkeUewFTUj4lWivhYsj09M7978dEou/uMyCBmdjPg4jf00UaTsg8SWZ26uYbyDyklyGjLiQq
K5w3RhFXXJXIYxyUpKPrI/ngztaGPNpnuYMvG8z73qp303jpHf3pfeKRNncLPATYqv5eLRaXFoeM
H2Xy07iL6LFgK+jJ+8lZ5AHdql2VBAxQVQLV/sVuYau4ONHg60nAA5PVpfZKQ5d0NqaZHxb3JGln
pvUC/W4wG2cLpODGR6CuigtzCpvgFKn/80rxhi1TzZA7aQs24dtcjgVSUtjxGGPPQcZa6jBgPJu3
7HGUUHVe6ZNDFohz6PRPwV+yK/JciQC/v1RBXfmTPOkLa/Ijr3z4OX4HdauT+sWArN/1K1RaIumC
xDTaPCyWYZ/3qtFjg0TpCgN+BWFLDhr/T8x9T4I4dqg2JVC5yjYqvL7QTnkoWQZv4ajWxlTM/VuK
VYSiuiElU9EUWF4mL2h9P6z9BwuRKB7KxszjDVhZGEYH3HPe9EMUiYVSmc1/APuJ9uc+diobWlBI
yLKtUKWUezsO2M+gpi5iu0ei0d9q7WttWScMqVjEQswZ/frSWcTv62NDijx/V8woGMe7pDYP455i
GMzOfOg078iaeyC2QQ4cidIV9yuu0wrZj+K8aX47i/gXCzjimOtA8rddPxgpJlcWUDdyryeVWsWT
oiupzSEBee/MSHEkRVQuKxGBOJr1pKhuRgXXTzt33feoO7Kvl3Nu4HNZVJsUiTYSTDwpIIe+0zmb
z06UEfqGA8R0tIUhNXRCm0ZCo4GHd+Gt5gfYKItTWtNZE9LF5bB0PLJR1qNPrCxAN1Bdb5RJNNYR
9Ku2eTXXKVd2hc5ITNCwOjQw7bBBCy6nvh/vxxFb9ebEd+J0A3dWsvl35mIqyx5OHielk5210TJF
ar814V0PsLwbnZqOHpXlThWoaGlSZvG5KyDgZ45JNvjDI1W6dJpOP5xllCw1hpCMSR30tA0EXVxb
gCp1hRxAxmLb3gozpkOXNRsQemfePphuvXfRCZDs0r0U+NarKE50tpXiJlIZrwXToHdFrkPkeb8o
AoSV9suG5zq9VoeLJ9osuQC5IhUddv+mxFzmDSFVPBtlRWKVynPzpANQtk1fHLGw7ghD/gKuaKy3
3CWckf+7gZKwQ9MCZlmb/mXRpxcJf6gmH6i9qIRlSn0uyAL5flIqNP8H3XSMmb9G+zrwDhvd9IYs
P5BEcWJ9chl+nPqH2CdAp7IAAmJctSdP3DAhsZtv1MMEMXGE/1Un4pHoq/Nv1sB0Mt+Bwg5XC+Y/
SbhjEnZ5RM4tbcn/kSn9NwaGCLQJ0ILzxUXjAeGtN+22W1kXQtYoT7kPK2C3fwCDB64URADYjDC6
oIco4dCSKtXfOhHjGd3sKAqGSQ5U5U7MCFrdQwZtJFCm1U//XW9O1eb1o6BQcMetsz8yEDqIoNjN
qef1dJYiGtIEqpppBbMa3B1gRF+ayF9hvhm2VgiyW5ZUrFViKXJJdqT81wGCF/iJYQufW8ErbaFS
diNy75ENa4jJuqUktAt6H4tOnckmXeFHALVsZjrjZ/Lcdabz1QmpA0kuUcc+H71ItuCXxmBwEWJR
xVX9RN/Rz7Bxsw8I0MCLMoRfYN2Ourh2dvst/we1IMnY4wevesknTydWCDyJ/xULsXcuPhU7bbfN
pQMAU95PMrrWyXZ9FPDmCkhywP/CYQQVqQhsHz8nnF571quPdadql+KrOuBwuozphs3eiHj5sU7j
Qku5XeB+KyNwRyk6rFt6MoJdsRY8CO4v5M8pmBYUiSFAYkqE9IoayD1DF/z+tG6R2ogP91RT81bL
2WgUboEG98S7+ItaVxcOqYp5BIC28GEocenkphdFEJ9a6wELQEdxcpTeQQGk6dnOHcepQhZOB2uX
O9UZMzVzzPt7jfwob+L7EdwPggWxXVIxJDBu3Nx8A5KX9pxI1kFEQZjXivgfSqCtyNFlunl4BoLS
dm4afB0ipblzf50ImJGk915uobBDR3EptLpNGsmO9CHqrFFA0vkS/yye+9YderPb3fwthx35jXwr
9hhbsf9eKqtQMZwa3h8vbbpwavEc9ROVhWKFwwREB2vz3q+y7cAlOh5HvEZaUIB4EGKfYEyjVDZ+
IaNB0d03/YA7GqFTDbHQgPPOSQaaYJINN/gq/66ltKZk1HmCC+bszShV0wyZc/1Iyk4LlJxBwktF
Vd0xQRoSXIk5Hgjlf8rSn6UIndumS+XolHswROfYqAqA4Fi7/621ddigQ3GESOGGHXQYymKRvIvI
0y0QxmXXKkHXvzXIQ9fvo6XMeXaGNKJ3aCHBLg/QnGivh5OTdgSRsaWAGVkATo7RbVtjTWRmnfec
19QDLjq4bh4TAO/C8WSnXq500p9jOvqHmYd7vNkTou66qxvMYI7as6L2xMN3LSHrIPcFyiRsV6wi
Y4FxHFPo0jCQsCMpeVJnpkE+4UONMyIozhiuyW/5Y98Gw/apyHesCI7Qs9IKRNyTX9mSzzN+L0HE
jcflv5ya+EvFDTzr7+Q8TlpgQx3YGrSm2CBOALuopzBiODMCQSwdQ8Y2jMk3UdaYy3fA2BH6lhC7
bh6iSEBRk1zRqxbbZfvKutsjq6NuGs6fKxQZnQrOmvyUh9IORIg72iwrfYV9HAVs3bL13d1vkOUH
jZGXh4Y3xwU+BeDDmXtdzHy+jYtME5ffXT+btquHoTd5ilGCN49rh/1AOOJ6YSxDMU8Jc65BXcCU
c/GGSPbPl3uonu6Qx5spCuueEgVHKpXRRsjiLG2xMHlsZ46cIse3eYODQM3oE7dhAFJl+t1O7QGv
yvItN0Rxk0n4VVrQxVj/piXY4vvd8PbjEotp+mq4Okz8g378jecR3KH8EtHLwxwLu/TChOfPoSRH
9sSJUgzty3lLZYBzJVH+qnWZyNFTjuseFPkwcxhraswZXveFiJVmPQN02XP2IB4sCEaspzNrfSv3
bmR76Cb9jAEgpra48y2P/4nInLWVuXqonwIe6BiRwHezMHiR1XAA0FJTT8nbDF+jeNUDYlSOePnq
rWnuGGMCq+nrjjmGAwvCqEghuvGrMlN21PeVzR06yBl43/oT6XEZN3vySYqAYxpk+3bp609vvdpC
xfuUPdz8b2brUi1OctzVMkdaFRK58RoZMIMxFrSLUclDP5NsMYJggjr1weKNLDSY0ZL41UQ13Dc9
xQcwgvTubxkddywnOgc2KqIdhSlEZfCqllAf9AoQltLfLalQhxC8w3k1sFvIohHChH5tl6ddKGv3
4CVQbBqpphFaykIGIWOnJ25uYQJaHaL37n75BlzTcZUSUxBxSxR471fu/TlRGxf4Ht/F9HxwDZEt
rnDjdcuY2/Lvl0GrvzBOxZdHqmpL508+z4bOulktnOj4DOBqfUQJjhrzDTHu9XtyRzFpqTF8dZeJ
2t7vw0sNE4wY8j8tzwt8MFNqRDDlOR7CZ0xCFiHWZ6qcQmCj+b9cW3++QLh6j/B/CQsul3ZULZzf
gTVSDRGhwdzZZStgA5ym6eFS/yGONWxezcJZM9/pvmpIzsmPsSrrqZ4PgnXfFzXN6oX2x83axzve
sIPzzmFGHGEY9fCvMBqUT4U4Ih+28YbeY0Xu821wLY9hQWR8O2NXZEp9xYXEcRjLc0bCgPCTm4+y
UVCW/RvnXX4K1ncz9eR4HubPoH2H4ccbmIx/3fG/pZn2tBL969UOs4MeX4xGzuPJwlbLIwsKwG06
lcczDMtiK6dI0/qKvpW+aASXaegPcx095oe1xY4D1kROi/pHM/fgireVuewb3bzqwloGbk7RYHnr
5sxRx77qgVAB0TUIjoAZQQ9o0tMk5VF+ytKBh4Q/wqKgWZT+daOGHPv+ZtWjsLcgzorbhhRXXP8n
nzNKnUOv2CAiY6Eq17pEzDteNLo4OMUyjwGG5f0vx/qD6Q+YLWdNFKW95QSZoJAg0xYkUNOm4HW1
PEX4oFFJOlCzWzGvE2KAYqKB+RFpuS4Hs7cWbJQfuiYY9A75IcdP3tlGOvQyjBX6vrn2Fj9KmfCE
aGAExg+CyVb1Ln1m93zikyvs4dnVBsvqFwEFng3GsGelfX+390UnXDeVamULEnVg1WzalXlEp+7x
0Vj6AfZnlCLPeAJjLcwcHw22NNU2H4NQivarBSFq92kEvhe18K64IARJhCWA9hwMwf4cxWPyswl/
yeV2xUFQoN9KqV/4/3C1RD4ish7o8/CecxhcvaE99cL3b1xCI25cTXXwVWP6cKpPQOGc6zYUQxJr
jWSGe4Ge3vC6Q5vt8bbXySZer+AIib8uk3KN4mrBbMOtI0wn6t0T4oMSKHYKWb66sKnCnBfBBRf4
vCPpV5WEb2e3eR1wHSt5ykYgxIjs5hFNPXyN+HH1aNWrq9d2IeXLxnTlk4J/9S9JRnp5VWSv3BNP
ukToTaAWpfetzIF3s2i288hliUZL98VynuOTM8l+s7RuIXYPTdjbao1bK/sYp+Ed1E9i29cA5BGP
W9DsQ2ybZbEoT/a+lam9/TmkTxM57itduax5xPgvukwPRUeLkKildKpX8F8NK66LWAzmjjLigtxU
QkwgYT+YblYBTtnwe1ta1ufUhNOCoEYp2mkyaGfKFeUkOUcw6Z+ZRIS6hAcZ+51XkttSIjL6WjXE
7km+pMLOP4rN8LVD+moJZtcGUncE9ReQGwmwfsECFHze0TMaBN53obzbgSSpKiGVHrcdqCLLwMOr
VJTUClBhpKcPfOnTU9Dv8I2GwDFzZM8kDLLFDVxH2eifeq40QhsY574xQHOJJWEmGZ/f5TsuIMKN
zBui12YK0HtScLF/9gbmWvvj5yE2ZOuEFRgvm2QebF2IQfd22Z8VtzTcAvSJEEHB0VoKJv4TuVbA
S6QHmxPdBA1wvUHjSa6gMWGmpwPHdxCmbcoGXxmaj8j4wVgkN5LVkwxN5WYR5svgQ2g7QChtw+ZD
TebRf3/LDvXJ588qEeYFm39hyvzt6vaisMCYyLMvazt+0yQkSb+CrDQQcnuTBNwYm/5SXJk7UOtY
7M7xQwhmXV1KITAx9uqX5j/GgP234K6OXGrGOGebS4UCno9wZQI2RimZ88kNSH3jWF571PgD+lVv
R/guz/y5oyqn/EMidSkTPSOmnA8ezNueccf6FAoofBzKETiyAEGZcv47+z+uYiLVKI8+HdfcJAy/
RZlBDZBeCoPxn5LSK7jpeagINlkCZDwHfhHrxMu2s+IbDxNKEitlv76O+kQIUaMATNE67PXyG6Ii
hDIsEKUb8ohXk///FiCRmwgGc5J35QbhaeiEceEwpdWzJpTt7YNBDWkf6xSIhq2WLooJSK9uHc+a
xuHfU+2X2VDAqMxKbSvpcSCZ7PMYezPWlG7K2it6myZCxaZj1Ait24yIvbWLA1jJoBVTTacIhX+I
i/Z3pNI6CdYsF5VcZlqafF6AzJj6ld6gu87SXPCxETHlnyIaudkf6tqKsVLgmuCXxK+WYL+XD1hq
un9jB0eoheNeNmuU9ecCXy3ESOvnwX5ZblIc2sfGnRJwO3yu0tpv85y5WJjzL63Iz9eQyTE1hC/N
zlsxej+Bgougd3blt91jPVwGcYLfAx71rH/Y2QkAcPCL7hL6HhJafsz1nF56GjiEUsU1gDaHESlu
/B7t8KBw5E1QleMsv8XtAR8PXECk/vUNiMsRbhGlq4MMTOzEGWGCxn9M6rM1mLc8bIfJJ8OkZenX
znYD1iDDkJ5pXGA1Cl2gj76Ce1MBE48eejjQxpabtWX/uQLjVwhsGw9kHYHfKcP0pNn36ogo3s6I
ZDEBtLV9yC2uncvPrIjIzpbYPlSsJfH3SVB/mrKHfJntSoENOJSa0Jvrq8z6j8v/SyV4wr8GWABN
HEuScgL7JhGXe2cwGlG1BOwur5hkPi30UBnI0Dv/oMe1K+JHb8FBZdqrz0orNMXiLKDdA/eaj7LZ
C8mlw3O9LMfVK1Cy6ORkiDCBhbyVlnIn45oOW/GjaZX3OkOKXUwtSk+13zBx8ZRWRLtGi7Buz6+4
pnJQlrO4eucnxVKosVs0Z8MN3riWWP7IHrGzkWrF2dGwbBuR/kqDDt9vRyP/MeDasKg10hKW8kyv
p1xMDTfC9//k4xoY0pHudhTG3hGzkDYUQz/Su9OMFz1x6/2AJPM/rOhT4O8gO5lBgI+dkrEQVedW
wM9OqUv31k1gsLPLPij46kqtgIGSByMTuuXweJQNjyQxcHBRdEjIaF2ML/iVvALCFly9bXG9KT5b
anzkxBTT6gPeMAx2VBPH3lMcQsvYqGnn/VaUP5u5xSrmbUMtXm3awK6PoBMF/pBufbFf3TC8q9Zj
A/GAaQH8gTYdQHmZ1pLA7eeZuQ2mSBUexMexMm6vTSTDUaOLaOlB94GDyZS75BrH/OkG5E7kzbJ+
ROvgPXIrKmJHen4G+QpwtD5j+QCX+3xW/yViDL8+bIewwtRKyWavWDgKAaPXj6b2idNAhelFelwj
MMbUk5NX8VTrBbIIe0jV1rfq55BzCi4r7OwT09gAgLiRwKCiVYVLkvtAp496q2MP8YNqzv5cZHkM
KJbURDlKJfBIzPePLzsMQfIl5GL0he2Yztu2bw3KpCDAaXdE+e7DrT0eghBLJcBxnuxP8BK24esW
iu4tRvHUuXVtbit3Cr5IdBSVv4L4V66IzHFwdLFlDHfnXAcrcdUq4zF/M2ehsVu8XFKUxa85/dia
XJEzvHLbdzJXMa9m4RhsuSj2Te0Vuv4Y7K5Xw303NOeOHqhNo6ehOnHpIwNC4BvaT4AOL8IC/Uaz
LL9aKt9mFOoycDDmBmwJHELAxMQ3iC5OBIdZCHm7cI/touzJWSYzxkBxjBlj4S+Vm4eH/wr4Wdhb
Oxog9+gHd3hCV1npOGJ3DF2G61GU8eDFesgBYgOQIXehJFXx5CMWN9GVDhesUfzrvUqivmLtbjS9
tmuWxzgtWRLcLOKq7va0P+BZQ4CLaL8Dngty3kKiC08L8qOnLQ9Ad4csZtFaCMRuIhCSCSQUEAsz
IMQzT+sCDzWo0eQ3/CFGpu/+eVmY/cs90OUEgj3OaElWQg/Fh6rPt7ZzWGbh+20rYjfghixp4iHw
xi7xlo2KlTNC92xgkPIYaPTQXPIg8RBhBr5edNGCE+6a3VWA69S+Uvv4Kk5BXYTPEIjlP5wruWl6
qSjTZeiAr4oIVjHIiVUaOt4fr2RIGZUXfKMtFF4Q0GHi5k64Cx3GJ4trh3mMzQQK2VeGnvC4ZctV
ieGHFmVyu4MCD+qTEqIuANHNWWYIcUU9p5f5jHQBFsBpJ5n6vrLjxhG26PGRhsmGlCiOYdB3m9RI
s4vJOidXUQw3yVmEr3M+uVQzygPYI0cLbYnMIH2BSCSsJqYIXhVBEZ3z+sIoCbp45iPxp9QPb/Qs
V6ix4shHKwM5K7ciM1c5hPuvvu/dBzy3wXkbrnw99OqymUv8dDj0eBAFTTZPb9TILN99UnSUjAWa
7bNbS1hqoN1+ztPhbX9UoCFTZcphW4Ib62GTtCnMq+2JF9wZD6xqJ6gF+/PDFhhEOHgT9hIKSTd4
WEgxYmFzGWTbnwOUNmViDDTcPyg0ZX+e7uOKASLGH3QJ6AMyn3L7Cm6AfjetHHLbpfmacNS3POXp
4PeUHWmler3CqPe6XwB8ZSLmaIhgoJRFdcvOUVwfP5WJczgO/W6iXBVHdGLGhKVLMiS+Iz1cu+c4
RBx1iUUpnQE18fAYPeeUy/ku2xdUFm/HFA1hrh4O27u3GPUnZVtN/PY1n/jwRG2WFO08PISHTSZI
wwu0r5RwJb0usQKVePn6ZivFQhNl2sB4C8h0zlKRDGtHjoMm8u3XGQP5PDBufi8eqsv74cYCX73e
bVi175Q4pv+cHoSs5xBpX4kzUoyXuqztRl+nJrAYEcmQfjge+LALdSOXYhef5KbnP4V8Qd2PSZHH
qvojBq8SbmQg9Oe08yRxH+6AZsLV1NmUr2fu9gnOoxqA+QWl9QSpKHVX3Orf4tR6lRLkZd5k+/L+
rCjB1it6hO8vTOqJwDB6on+AoS+gEfng4rJMAVgOTABFeKXbxiSwecjCc8gsWY4lrtWwxBBwUamg
qHujZeTGv6czAbVvoH7kqHSYQBfWqe1Btw+OpnAltVm5PejBwwGyWHgrkKQljj69l9IqNxlvuYCA
FKCL8IP7wa7FIy5ZkAeyy5GaqMcwl/C3GTb+KipGCxknOOluTHiZzw4bJuV7b9gMyldRFIEcv6So
xf2xNjKayGg4lba4pM736ZijMUyT6CrYSCsXi1z/h+ogR5RtYJrwFEYM4Ua3CPnDStciaFH7sez2
uc/22m7MqOCnRnwzbob3Y0Nkot1D9VJR0Xg8tdzlyLi+F6tXnMndtFkFfql13uyxrqdmaFsV92//
NkWSToIMOVrncuo5iLE5Da8eyEq7WVk2U8gYS1MSjBkcFmZAPi23JFmPnaJtDx7QXFKtHGzi7vVO
y8swtzE8fO3eRj7pw5rWL2/QncsgPPpCdDNb2evoH/NqT6vxecXC9vJpdsos4nFEPvO54ps0nByv
03E5SCcBFPu4PZjS/F1Zcuq0HzykHCOWpFTMeOp1cJVGBlf6gRrsO8VEaZOc0G4QFL11ZNE1lCkA
2krqahAmkWanESx60iD6/+yTV6caHkwPyR0mcxo6HUhOvqmfvw6zkbV/PHcTbEEVoUuA1nkXC6m1
G2tAIfm2OvXNhbS3Bbq6xYNd+EK4Mwy8WBSRvLb9tmfsWnMX0/FHjXWzDbt6i3FYz84uZ6giS5xq
1WcTT2DuUVtaCR5c4soGOl1ydm6ll+2Vz6A3/fiq+pTlT7vYHCwZjJ2vnEL9N0kZat+/0IVSOyPd
LhGf86ASGUzdPRPL0KUfb90plZvtaBst3yN3MQXQVbyxI3Q4k3h7uLoVT5pDwnDdgX60Cj52fTng
ZzUs4eEnLmTxk66OmD6PidWkSZNPaGQJ7zzdqmKvhFwrDCVOYszZ2VqV0mmhq21LY7g2vfrqbWTU
6dy9d3EhogIfA9sBXRq6akyT/gHAIEAtNX5qqB6kAKJDdTVoDrg9Ih/ht24wYpfW3pQyF79OuDKn
PV7WCg3bTFlLAYBbVYo8QO2gQDF3djzSmzpG5Q6uGGDeFAGLvUgABz9tR6wx/MUdIh98VZz0Ha3U
DPIWjLJFAyF+1uS9O8MubUd9YXY0dAmPBqIEtyhIzGB8+reJHtrNqSAVkUwHz8v8RmbqnCgRb2mS
2vlPy7BnOzAbTCFGqednUeuHpGodEmHpdRpILK73+JXU1QCBJCwKpD4vcQz8LHn5NSSJyrJKvsiw
7CcvYmvXBGgz/v83q/ef5zsRDeP5N96cppd+An2s/i4d/iq4WhORuMuxw7dUWy5lwZAPpIS7kzDk
NoMLHGF7j598ehG2zJ+rfUlf7af1ucws7U1tw5f7qVXz/bFguHqaRE2+lfQk6H/ROP+/ZU/9hdSP
XlvU2BTLsfOx39/fyCCTU32GVgTXz/Jh1DvJ/WXQf0qtRRgBRGjSGWgSpL00ER0h49GEN3LTFPed
hmCPZR4XTV0o4nkUbWlOCxwttvGr+fAUzEiZPG/xNKtaugkgBl7bhrRAAGyJUighkFE+Q8rhmj+Q
qLVR+P8qr9fWlOJijyBoEuw7QyRAIJsxSSolMx23u4JHxzYWcAf1NWQd+NcokafDo+VwQJxV37ga
Y4oJVN82FTEjPaF5c4plHk//FcFazPnXfkIlTTtZWOBJKe8d2wZ8UgASgWn4tuUO3ry6ytO0RcgC
+dRhkS9O5LoQHmZN4hmGNGVD31/lTapHnb0RyWa8UCET6ui2Mr/SzxkKMFG2xgCRBVH1QWfv01Ey
Eubra4MGiPBCsRa1I/W2fs3oCpTOHA03q+h1BAXGLLYsfabF0zyZp+hK38sFXx65uCtveOEuQbQe
luX0awQ3l0hU0WMnUIzN2qYYo1adLGh7TBjp6cik54ou37QWit5lJhOsuq0iptTFnzMkdZd9Mv4+
FipfGpyYUslg/Le4MVPuHOo4CkJzk/xPh2jEABUUq4iXTdCsMyefOhRM4dSxoDc/ZmOR3/CY2K3l
nyn+I9cIUkJq/yX0dDsHhgl3jGlKG+xJg0RuyJr3bWxYkVtzKzWQ/Kdvhqctty86dsOzY/fELiaF
RKiztxiPmaimJLTlCdCcHVY+GSJaMoW0wwjJum0xDemuNmDF8lyZ9xUQ+4lGPWyjGWVFFsx4T8Of
xMhiBHvCsq6bMB/1nNZBJ4sFBWDEQyqZ+Zl3+iE3iuov30o28m/vySUVS9Hl2d2ReBxZpb+exVEl
so3h5S+AXLQEf9/IKxdyQGUjMgurGltE1f4bb+TItMksPoMmqt5nV55Oam7z8fhnEjXt/UgO6XnC
ZZLhTA7WX7jNMT6SwHe3qP9XpbKQmTZlcFQvgTwP38dNnMl5I2Mb1J1UEPHK3oq6UYBY4TiJXWLD
WwQz9+IYtnRKfAl4DavlNxhMU9GUEscIt0I/FwkRsKXLRkaojAoQV4qiCmZts/XeLQjpb7Pz9APD
OYAcljXSAgOC/xlWKNL5Ye0GTe0V6Z/wpSGsDPl1jRkLnicWQOhfn05SSaqQ8gxjpTDuth74zlHY
muOdiClQ1jvrxiRMYZNl1XHkdRVPMACCdsgRVjPXClUB6lJhUpLuGvWezL4PyeWJi4XoTo/KVf81
49AhfiYFH5+zgfeyOSU3nbeAv/o4cStlMA/YDI2QX/VEkPiY3RhivkgkaunjXBXodBPpSJMp212R
epNh12SdJ0F6WF/31h9+d53JqNR1sdN6bT9OITtvwXjAPi6h6ouJzN/aE14r+vIR4xD/fxsBqcAr
5tg6gYB5LPgPbLCAxueBVbGdSYNzYZsqmNslItbpCoQduT1wz9sWUteOkHQxvr1pR3o0wRTCnqQV
QuD8RFvR4BDwWun/BwxrkvotxoEWZDDXXVm8HdkC9KMTQYgyKXi+1JCwt0UdV/l6TkqDViwcPvL+
DklopTE4Wt/nNsiNtAvJRgZBrruio1ybtvMOnoNjcLldGvZPHx/0cxyGlZSgdzw70vNEsSsW0oRL
DKTqW3S5SAfKYgQ+nL+C3RbF/38qTRM3nz/obMeyvJl1U8rQUJkgw27m8I//UQoKGcLD2k52u+7n
4GKnL4Do2/KLgxmrgQh0PwgAt2+7Q6n27WkxRsydETKw9cafp3XHi6e1Ls+pYVvMFDTjUzJKLwD5
SO6tqN6311jRXcHlPRueOC7vIKC8tW3P4wi482q/kzRInVHKBmSUUdG42Or7te5ejfJc/+DuoB+p
KiXPdx0mGbEG4OxlMtkh3oPEY8YauhLzFvvsidFYuGWVzOV58W8Z95gorSfAoMq7JwgmlOr0yXUb
EO75lP0s3X+ABX0aoFInlxcHlZ80qbmKFZql/6t0NAaWJxtQP54SGknBbEaf40nDsm08QKCplQI8
zTkS2PAhheZBOf3w3PNybNJevyaLDPIN2o7CaJxacP/drs/kzmDdKhXBiBB/4Ua4d0z0HA6mb4yP
UwMknGvKcrVgbZj0t1GKNZD8ij9Ar1ydK8ZGSNahSO6huZvhjuIu7Eu99TmqeqdxJRVEMdE0256q
R0alsZwckLELcH+J124ClC3dnDcyi5rSy6S3S4hqQTBDh787SFkysLlqQD3gJBz0aSJllNdysVct
1YHr4/H0+1KJJas+xHHsM8c2no6vUlT6Q4E+Dv1tZmsr6QEQUBmmwX8LOLpFFX0xuM3JgEz0vA+z
dC3d3Z0+EVLtjd6vhKT8EBRFyY3nLft8sUzO0en9rDHvSHT4cQCK4Tsy/7/lXuu36ChzlqawlqPU
49xjmje+c7waicnSttwBProeYqMf6iXlglN09eEZ2t0zqAoUl3PjdhATphvEpZ5N6OgruVeaDn0X
xhQF5VnsYavzZbEA2yg6jsCzgJZrEn+SoR2QwRUXvhKZJcl2UNF6JRxdThcAzPl3JO+8AmjE5Aci
P25KecjY9qMe6u3A6xY/sk6X7/kyEol6APMFTG5ALj47EETQqPZj4yAujxdwC5LDG1kIXF7oyD8L
BTCOZmVSNe1yxXFI0YdtVVSXTQW/VOTS/JifSe2ysqX3MvQ/y8FYARbdtHlYLon+io6X+AMWsbSi
h55gkFvwRfC1CzYkmbpdTywhs4heC99x0hGOFDOUkwBFHhxMk9B+HJIe0bYLIQlqkn72oA8Kzu86
JmRdoYNdrwBNiH/wwyJXF4ufTj/exgXIXnifTENHtijJ58MlOhMB/U62Fb/yld0VZKxrD00O0e06
ZoTP7X3Wpkb4z6diptt+erUXSLmPvEMpiyxJYI9gxnUWuDnnHO1bf025/1z/pEDrlBhaXXOFPsmA
gR60mg2NU3uPgyglJ3ibRcaKT6GrpCKE3YJIhmJhdPeE1IW+nK8iJ2K5gILZWWisf5ZVeE53HP5c
5ha4Lqfaqk9J6F+Xl5qXsJFza2i+nFA9WFyfFG/5AKoFT3Pge+RHHCwsjoWXKtcrtzlfCdGl8NCJ
agTUEnFE0cIEI7qf5zc/W8IlK0pZpUkghh4nooEELSyiQ7+LoJD9ndWdy0650nnMmE+hdtkLEGgs
diWVICWXhMyffqu6zGp3ER5ub2IMHx3B+KL9tc0T7IcCO6tt08CoXizsvd2oMOo9SR8mIGuJuxrB
fok4anHhUMDivhw6WwWmIY+xPHqrGfBJM3FI/+Rzkj7z14Ucl7MagHdZsd2vXisF/QaHobNlJZIN
yHOsjvje3cp1BI4R8F/50HbGYrgSX2eTovosWgBGQqSxtoR42RriG96CkQfwpJcsIGpkDVKk6IOi
+jcAtCQKBEIhQrlr5gLRsdEWkXidbG2bW177zR0mmuiW8hzSYBNKNb1Lxb2ru5FNSo8mifEl4+qf
lQTojXFBFkg9cOSUD1Kz7YHoB1U2uF3Cl/y0t08ZQ1H/m7dM9PPJgX+5pOkXnRX7TO4Fp8y7Oz9R
cdRW1vEKOeK+U+jNanPtQUtlFxrPt7/lciKjLxFVThQG8DcZXN9UIjlh9GJN3s70GQ8K19c/DyXU
2DBpp3qH1OhzxfTTJsaK32RlPRT82jkE6RJjMsdTCjpiSH230qTuDsfCCCbLYlbW18d2fwfFpqRe
JYawia5Srw7FTB19jAGYIr4CIZshzxXHKXPZgUDcZLshx78i8nbluW7prJ/i34HJc3rFZyoGHcO7
7GsITnB0vkjcGF/4ETXS5uzQGGS4P9pmHjuj4uNLcD3oq15lca/Wl3dDKwkIRs4FFutjKiUL5mxd
aOxC2VjTMBWyNlUIuXZXePVIjL0e6WiR6rEJnUv0ApuKS2Evf1bWmPRgG1b83e25huhiQ+w389pg
wKKEBFRTUG/e0TLggoE/WF3xqusl7r6DBhuM2/zSboQM5WBxmH4uf6nOhvjfgSVoATW3g0bxXJxN
ao1FGpqRDaCrrz4gSNayrO33NlsI1EMk8uudBbJObazaDHdSj5OdeM/hHI1eQZIou2EfTZowlnEK
IPI+iBbCjOnvup7XQ2JeDoXSQZppsfP0ZQLsXKEsi+55+wRCuSTGwEUvna6EJ0xEzAp/j83DjHvM
Ia8JslKFxB6dkNHBnDNMO1EsiB8iyiU698z89i7drNypltrIGR1Pz0Ust0o0k77F1SpnBUB63TwS
qCaRtF86OSfodayJF1btzG6cjN5hZMf+hVvsBDdew4KjFZVrLetIpJyDyG/P1miPojJtdXuXOikM
+ZVDFCaNmQsDTJH+v9j91Rd/9HseSfCaEgRyl9ztv9Cj1iYwt0aWefdkmulNtexjotpVRacwP8Kp
U+oloL5QY1/26pqv8mhzbPf7roY+k/AyWOn6aTFtK0PleATJJbfpvtXN0hLXyNz18Rj5/Gfk1jAM
OpCUz45SnoMd3ItZAlw4QRfQdNcM2q8YCvTxAZU2zXzp1sMpvfdEzep1Buc1fR+vnboxcgXubl+r
vCaqdfEpeBwV46KSvGk0TBm4yfgmeXLwCRSKVkpjgGA3gC52xzjrwIYQMY6ga5G9IaRDS34Dg7U0
+gkhpqZTMMB6CidhmwIJzlKPMfd6wSH+9WlZOBwINzdyYPA0tKghYBGefYFNX1BQGZMCDslUov5f
t/9p0ks78RqhWDgcroKqQJcUg24uxqIGCTQMIn1bP24mifErAPql2bj4BZ8/6EP4UJOzD98CPFo3
Istenfb5ci7epvA2S07HtgrYErSEC9YXDeTtZxSFeSWkkbNGwgvsuEmcIkc7wsHcrWX3R6yf8cvS
s4A9NVBZZAitZJC41JflOzBqcdw3ftF15EOHz17FKTFRtQ5GUyyIRQ8M5QnC9Ero8vvg4YxYwBuV
uqA39ILSD7ZqmTw9PCXw7pg7vKCcWbBWrtcyDJa0at+PMjHXlv8CEzrWZKzdQVuhkSCd3+S2X08R
N5+sKkpgc0Qnbrbgrbb5MAsOwuE7bvAyUgflWOzOLwrVb3ZkVi3a7QqKKFKfWm0t6t2RAdSSmwnR
Wmk6hMP8rLGxHPQiWu2UkVpxn4p3lx5MhEM2ZamJWentPQf2RqpxonA0bGOv/gIfZdRKaiVruPIh
l1L8y1IfY+n7UU4sChu4/7BXdN/9UYHPZjBIFnddfPlgA5+uwvMECh9b5OYvj30EC1HRGZXXId79
kJLR+24hx9Aeo/5RLX1CtzNb3VEKLfLZndGDcK6tzlnBwf4geq3WTdknssSvv5iuIZ5levzihvJ/
eAK5J0PG6OGUFdUy4YCzN/FTSoXTTjUJe6XVobHFxnWZxlQnySqxYejKrH7Y7l2ZXg78nIjI9/1R
O3wDNJUeeERcQeq258rtR0xjTpdp5H9PiyUtPHQR1B3m8/nso+BcV8DnIrUVTPU08leU/omHkH3/
UwFscnYDKpQ/tbGEDmnzW56RzNVSeLv4opRn6p5tfRMUSqwtEbvxGRJ9cRvmipaPzQL1kt6QGDSp
BP9DkvYHVCaY9g2EL1xM+abcwIPK4Aw1tCizqOb4t/PmvOxJiJpRcnRDC/A6aEerjYYfPIiVA8Qg
WReWKXCZDyU2FtF2gVDWQJnzhhT0dsqTNoKxSkZEMXVL9i3fL90GRsfriILND+m6Jfy01FMpZbyQ
idGXr5uq/EGs7f6IacIsOqBoeBHStvItlBRCKfXHhD0zaEEMdbPjv5URAs2S+xHs+T1pU6vi4wbQ
RsaMdAVyQLHEXFAs//ZQJmTin9W9HYz2iL75zOYObXt0yZ6XvCOg/ddbaaWw9ksUUy0rPNPMPm80
IwsRRHYVWFSxFqeVP4qp+35FbMstI7DUuSs2P3n4Bd6/szvvCOaQLen8866IC6XJcRGPHsi91hXf
fdeiYutvIDeXXeUKuBgYyZVB3LH7ssZfb7W1ZpBFNS5o80Mzl9qrejjSkVFp1oMSqcYus6ZRdRUw
cW1Ou0wPZ4jFdsL/fdA35Y34qjjOeQSUms/vKnV/uCIBmTWgF03JdczF1Xr2YsSl7A0nD3oAFHpl
2q0qCO3XZzG7Rf+ykZY0PEtcYOLMoebZRoyLpL9VLc03rcaYTaJ7FgzwEDhntoLJcoROKvX3+LJh
b5lcvaB6gcdufGzeeyDTuvHBP1Yr7+QAij4k7kQ+eHdhQ7GJX8QeTyIjqph/QZoFLVMXWKEkSgsQ
b9AOMkGrdCU9HiEYWqTTo2wW1Y2Zf5PUFn2O1sACqUlZYvpLGpDnGPcKqLxZZZDjbV042eo8XBfw
RHa9mQNpp/hFCtnXlbdpUPwlphzyYBxPe4Htvvf85NkpYuiFyB4FuUsKe8vfZ3L1ZpQzjWOzSOYd
mMH0bB6H29M8dGyhvtDSQV7R5CPP2k3WM+2oTGHxfIicMRjyznaViY1yQmASBbE8oB21W2iIJRkY
Wt8q2iiKSHdLi/zamHosWwMKxYXJfMGV1ajTW5X7o4CYQEijICvJgXGl7HfnXA0LHhxqjiQbP6iV
uTrgsiuNOc2lMnSXiPvZ606oUilbLCWtB45Zfb+pZ9hlVKMGzz+sR+GgfuChqinD0wUB0hvI+KrI
8Xa6LKIiNUKabdCoKcY/5V62tPENkFoVwLV34HOHlt7VhMxPC8XGbUM9Qudaa5cchJIB0dn3e6fY
BGPgwNKNAMZ6pjjLot/2geay5zFkTHSzYOjae9I6NzwM1Y3WWo1YH4g3gC61mmLer9IdFJiHdVvI
2zVYlKl9ax4PjCdkP7jbYfiLs6639JPdcbghslrcU+5DCJ20LfadzvWXvkk2pmb4yR8tLSFxofsq
YtADz2rHUtAPoAVY5gJODLEspo1jMuYtcQ0NwvS7nB2LgTa+16vgnoxKyPvExrM0ooKu6IcGvgXj
JluTtE/JRUI/mgCaqhT+R6H8kBWdsyLfslYAzKp5faBJ65FanD0J5gCZnftL68l1oRji0Ng8b9mz
twJoHRCJ4zl4laL1dFCwRBQeSlm8ZvlVA7XBHUVgpZqn5rkvaCizLgMUuL0HxAL7NaXsOUNoXoiP
ASxQFBBluARN28g7qZVwug+9aVCVL6MlEPl+1V3nf3TYR6Em+DeW5rBvl/AOsxgVi3MEChWaq7T8
23J4rlDSZzQ3gQwCZ0qMqhNHxWaV6fi0Roqh8wHQfs3MDz5OgeZw9c1+t6Jp1PT90rWrgjDYRYPG
yfmx7wUyG6Y9MA+WT8A53dReaTpzyNuVonhKio+3oqKHVS7gdXM3m3YTBO3cPSh2FzQFBLMdYZq0
1bkGj1pKv3H5gnun5ENIWKHStpx3JrBcW1XYRatKuyaYQYtsJiwALuCHL6THoZlqjn9HSzJpXPey
xIAlX0OLcYcwTb4eEkOpxh5UVew47mwoKcwXE79zY6Kvy6Ee6blGAs15bGHEGv7kpiTntveVH8qB
mVOkBNUsm3qEiNeOfbvhkXtPhuYEYtwYTzlTTn0gTd+//MCsRX/itw0aRcwITWLz/eMdeiHz5BbF
EBiAaFxj+pv5/bnFgcWnBmA8hK55EdfJc4u2c2LKwEPjWlrQmo+5nibm9mLj5WqHYrFBhf68rW8+
RgAxGaSCy5gFFJ3db+5gfWkNgJCM5sPmLhZjuQEXwTEeC3yRYVT1/IchePaidds0eiJibQdqX5i6
RetiTWelD4x9wyMlo/v04x4KPmS944Uflyh5wY/zHoevPeDId/OE88y8FJMddq/EYQw7QD97jgJw
Rla2Pa5zS3OIGPLQQtZXq+IKHP26ysnVuFiYW16TAnJtsj9nDy9gfnmDlJQ1iyg7dp9M/M/Z1MPx
E+eX/NcnyMhN45ZBEP3v1OswLWxgPoWekecFNwxNpRmSDdWDNenoXuZ0suQa1Lke8gxC/bfEkC9Y
EW+8/LC6LQLaMbQLVtKI7tj/Qj10l7a6F81pmU2A64MgDf4VxDb/dEcw/cFqA9K8zJkLlf5foQdj
pmU9v10GUfeXqghhDkUongB5cHskHwQhz99KKfAJ5NEFIBrHEsspL7lLZaTgvll8GaGYjh04rYhw
3O69NKCL6nNBb/NT2Sxm//aPqns3jMt7g/54szVugzJlC8Elx6ThKSr/NCTExY6gtunMu1Ed/VZ2
5E+1slU6soYKGe6T0AR6pz7nI4zzNnevNjZEFtz6+3EtUnG2FePMbigRNKiLQ8YbeWnbE4/+NTLl
USDqgNczSuHhEg8ItyJZw0Foyar1oshxjCjt3BlAxUXrNuUIXbJOc16b8lQrt2SoWA0jELOcA5Xf
x0ePjhEW14MQfQ1jXbi3wynaxDTCec1m3izcDi9xdrkhc0bv6KUMDl/k6/B3UEqT/ievbhmWonic
s2NisRXVEWb6I7kcjZ9tzvEckaKHFSokUOsZ4IK3q9uPmqFRe4zFuQpH7uWkiC/f3nbzv56YYjvK
TV7IE7uNRO5uZe1ka0IT11e2lAuYVUndyJKbvpG2DjqzFDYjztSv+J3EvPnaGw9P9EZHpSP2IefS
A+cVmO0Dg9WT4JNs8/9P07iiyqG5rV8UB4Xcr67ZvTKctRPW2z0GMfH9DblfpoE1TT3z9a9QVlnZ
RhVhpS6TN11Tm/037tvEUGnPbE6XfAp7zAHJNYhhfcw3cwDTo+hkWKJf19Eb2N2IRZOmmfLT/orY
aST2JAhYMCLn1qWEiuOIYyC0Ib9cc9RbLEMEn0NmYQBItr+Q3gajCJcN9CrorIpzsUBMLktv/AG/
4odQMa24rEGA+onvNjrIN77MMC4tghWEftb+F0Njrez+g9BvLzyAJuugbUWfAt1ckQJ3qZaKq2nW
NkwMFlGcFHY0p6fr8NV7VmHkD6Oh1cZx/oy6veshhIsfzaOSG9/HjvEvNUkECLL+Eph12G15/7Qz
mKQFaK5LUXdx4Jdr/IVEwsmiZG8WJ8J8v8xJlgWhA9vzyEu84pm4HW3rJ0f7Ke69urD1iPKcLr00
94BpqqO/r5NKC0LA1uvjsS2A3So3Jp/k0nJSAWJPODZdEfjAdwyDrd3E9gkg7gspnHFVK360Rigx
sI2bziGn+IaOIdy81N0N4q+xHNIr84J6+EMFG8hTXlTNmWqlkp6sKrj+xjBdwzFeoOLg2L79ok1r
VDofWN+Qm638ChLtdmsPF13xGRKxA5rwRBqWR68+5g36R1R2c11TTG8JB4FfQmEE4s/+981520l1
aFX8pYlesqykl1BdnvwEDGpHC4KM26CKhKEkKwDFmqOn91J1pT+C4XlXjri92AztfREYmbd0r2+1
EL5W5eVbZJADCGXCt7rh0Dv4fn8rWfn3oWSBYEbIbLoQOenyVxQWGu8bKvoAUsTLVyEccq8P8NZ3
QcmtujEm6ShGoFQFNfDiCuaxw+wgEN9eaixy8ipdsn6YSN0GOBpqLOBulq2+Wdbvg1EAUmmBkCt6
qeORfZNV60CqnKLPBkzqcUZZiVg/BAYch01cjk0YEcUi/6pURFI7NpQEUyWOpz2r33KNSjZ0b6d4
3rKTLjHIy3rYlxfdX8PqBF2f/aaB73syFp+v1gBA6l81eV08lU318FNvOUuabb5b5VYsEb27pE76
Dy4upiXs9oL+f96NG/+0a6X35Yt4Eo7k8mXe+8Pcjx3mZMl1rOgA8Cf/c8EUbHlckUV9ECLQlwL3
OOZ9eHSkKi1lVtIcLZvikgMAm/qbfqSjVRY2Y2oeeqK9gI4jNP0Y8CxxEunVpD9KH/qkW3MsygG+
q1N8MuYKpO7rLTF4k2l0Ui2zBZcpslFdCKRL5nEuDwUrojU1m+9vJVhWFtUgix+U4CV/iHHxU7Lc
+NjnKBkAtqzDfLfYdZov0Reg19q6Stw9P+hsIDkJzOhfn4wQWiOoMvkaFVnhwvdXfb9Jc3ktiiKD
CVpc+rX2osCDDqYPWBJ6SMdAs3sDlqBJKIitG0kLw2DxxXPRc7IZjEVxT61DbRYB9rI6A4BNrTce
oW7YEm0N8OmnltM5CI3di+P1kpT5se0wEfUrgwjpNZ6bdycea1mUIDFsFInbQ4RHeWKcsJhr2oVp
79gRsSsJ9l/xu4fMLB6fJysg6s8+oiNKU3x2X5tH4nbQTaZ34IT/15L9Vy/u1Aa3xAv1zd1AGH7U
mU87v9PIBOpAU2Nxfa4ABeKGxZr3lDXywqPkzHyi4PljEwKdYe4dW9Y6VTckXPTFiS3xsPaUXaxH
Ju/7g4b1WabtHR1FaipeQKKxwq5nJ58Svl6OlG7EqvHErCACkN1GmlIDAANnkTcidA1M3tuCx4Q4
XwGQHRytZhQph3wi/68/OvqkeNXAWcyPWsPw49LSQ9o2FDn2aLE3TQnVxURTwBnybIAhswE0bhC8
V54uKalJeNS+8K3keCzfIGDlBblIfiu1SWW6EMNTwV89kpTXBQfMzgGoDYRKp7n4h6Euff9H27PD
ArViha4xngc4Kmad9g5rHa8big6j+BNW93qY7sdK8MoyQgcyuUpE0a7Tr+0knSJkw+50I88ZPtBr
iysJglZZgtD22SDNbbGyOUeNfJSsI746nWloQenuvGlMG6b000gPCqOGLet186fLlvzfF9/VIdkB
DrZz05wTUGEcc97jB7RhPO741o/tm5QJKUDwgCK13MIWTbXtKn8pzdfZiDFuQUmmbpp36qXodiVw
VJSze4mb6fQOE+7WTAwU6Wjso3r073dT7fyL7fiKHcRqcTY5sEdqijFUa8IF3x4lxNEFFLZ4p5t5
otRB6e+tWxSsfSidErQaZCFX/n1PeVdLtqevRNNCjq3YEBy5p35Kbvv9RJbxcEYAn4WIdqiYRm9v
HVK9zegVhLoRBBomYMRgPyeo7ZgmOmVZKVILBkOf10N56X6XfighrkwWrULq3oPGv54h+13EYgiW
T8Jx/6/WKmj8Dnz0XF1IEk9/+6uSdHYFrrwToUSy6Kje8pPllWv1lu/CR1q36mTcK1yjXFuXd3Fb
oSBhe0fdSxHqAVQ3zLKrU+5ZnhTa001BG0xXonBRjnmSQ/VVDAvbYxi8piiSU6nkl6sNOiInXPel
EoyygzmCDETyk6NWevCr4ZemmjQOKFjfNFdPZTbUIrdzJQOgCQfgR/9N4N+eLd+ZcvRkI7Z0+8/Y
D3et77SOCC2lDptmBA+iagX0p26L1Mo9LPf+Eq27LwrUzMTteqWCfW2VZAg7G4MwSgMYeqi+MVGh
41w22Whp12ojhqgzoRoU69wYPzpJlcxlscJGHyMPHBsY5zhCugtwNhvVJl9D/uq3sW1wnFDDPevT
g5Ek/14Kfu/DiSgAhCBv6HuJx8VdrB7le687Tvv+lDLXd9j88aRyjXhSpRMypSv5Nya15DHC/xvS
bQVzH5tnfgR0HpJJwe/ExDbAkoFTOpfpkZIKQXoXzOqTHcFDz1n0NBXpSn9sUGXYScob68E1V6bs
axyQfnuQcKenEFJAiASAZd52GGAGdXcJWsgjIRykQd891beNHb9AejFLsfqNUS1VIyLeFJ7HCXt1
LWN+e0BciJBaGj8nmg/2AjC7qGRYN/SP/bt7nxIIWIU/sM5PvpCQgzv/hmDzVSxYr+NmvUmcsdYc
snKMbbsJ0IZ7yfiPvHJeJBAxdC8hT7G+EIwyca49vjIlfnV/5CYMvtEuD7thl/gg4uAq6G45xUNC
aTpOkAtTX3MwIeJmNOx5VWTMagqTvq3aAK9RTU4wClI7/J05TrJqeZ+GMlzNIBbBCYd7JLmA72+3
77mqvzgqmbVwubkq0Y1KGzqbGTT7EwbL+daS8VraRHmoyYWmNuDnjbDHEEh+csQrlFIb/0phKmKn
aej7bqMjw5XKsJ/t3ZHQlyC99GwHILL2mcJ/RXm54+Z3imPDirNSJ24ntrl1+pZwojn5ixNB+2ca
cKVPpH37yR6WRHYjUMB4N9gKuOE/3aQhQxaq/YJOyp31prLZld8MGnGtlDa2iDqY2DcJoscYpJKN
Urqqec9TwNeNdkwKf8aRjK5fZ6klDxGUA06HJzvB2HYB5gAenOwd757suNmP2OQEDB7MGX8EoGwb
0FUWmS19GmTKlIKguQsjNJDccaDDwx96kiOgzCvJjNrl6A+g/QylPWWJKrQSn1o/v55xzuLWGvQM
7pzxP7mkVjqLWB52Tr8h1wWjF6vnZqjhhVwFzr10Xc8GatE1yTyWk2m/qZDhfB7gQr0hspk8RKbZ
s9Cm+DPJgDa/hbCPKXbuGizONk0Am31WYpUGoLBdHIxtwcN9HQ/CaZO4FG9j4dK9+Tb7d7/I56Am
YX/hiwv6dn4A7hS68FrYSnQdUfltZD4lP/es/EZwQP/oyPFxE+lPdws9njj3awcVadQDZtY9bOVW
gZpITEnNB/h1m1fJoODec14rh1QaZQ69lFow5TdqMoe+HWpUYyMcmgpDhByqf7b2XHW1fvmhSQ3g
Isl8QLlp7jXyWDyrgoXwGyuoYBGCj53tuqCSF5p0nDkWOdU17wGaLUqCmN/0N3fK9YOPe+VMDKNR
d9HgJz51s7HRj0j5ms/+cGcZ9VjXnR9ER7toQppmXlzvgk1GuELXg//Oa6MApfboJPm4I2aiy2RI
h8g8jv6m88nSWIOr/ITPFsTwpKP/Rt8wN1PVUDc0A9frUVIrGYbdOFIHr2wz3vxSZ1Xqw/LXA44P
i5+SYImVMl5JhXjyq4Lq7erX5Q50ATlNCAQ0AubUEjAjc6iI5oFzYzkjSNJ12ZiNwhe5IRK081pQ
kAtDrlNLwd3rELXr++Qo5/sShkFOC+gaiOVmyUPc4dGw9++kVR5GcFEubnEwZP5ZYy64VVC712Rq
8SLkISx6G6ezSySsIpMWG1n0q73pfNs/aVzIIAfzdQ8MRlNBUq/LTqvEVvTjTLs6zoRZfBJxGUDE
9FzS6nE/MHMM3FxRrGdwlLI3fyrGx1kuG5IiX502y/R3ywzsMrCnzm/Geys1JY83fPuCS60oSVsm
GH34AN5VuCMP0UnxJ1Gtwi7EqcVreTeEWttPQTPTyZxdoCJwX5fF+/OFHTxnp3vbC5qO1JEL2liu
R/tsxf3pTV93SIAXucPvajMIyzHSQbpOxiNFikJgPtcjV6sesEeOMsY1FE6LBeDOUAIxMFRA/IGh
9WoaPI4SUXMOmlKUwLHfX3ykA9bOXkvuywtPhgNmARCd1nKwQUChXDWJZoOoCe4w5jNyFCCiuCVr
LeqfHk78UQ+A+p1qBl5xVDt+e/WMmyTyoO9PrVOB+N3WlZBdvuRwRsBXfazrlGtil5dJES7hddGZ
nCaNZb7+Qtvegjn6iATwKADcBFDJHcX1yx2VP+x+8z514G30ugrwIwsrvX2B1WBbpoHbMb5Tzd3+
RZmB0mhMv5p+UIj/7ZoOoKf7aAaZoHLU3d1uJTuaByGL/EAYSCfZ7s/X/UgXXnJg0DvWpEA6JKu9
vXyryR+bwNXmDvEEvalvLfbfM9mlRUfBvJHdrmMIb1p5Z7OKJXkynSGciaHB7V605A96mFkvA1DB
dmzGMCyvm6cI8j4O9JqjkcBkwpWeGddp4Rg8fxFNc8jEmaM40gjVDWSYKY/n4hcy0UA1oFVMdjoO
oXVY+r21AbiaM6ZIr9NpkBfLzf2cLsb0cK6HLh1HsMv/KMT0QppxSA8S9LVA41p9u11gLgrmDHR8
M1tV9EGqfuSxUmIMtktH5Hdq3Yz8B4THCU/QVrDE++aR8Vhii0JZLy0QcpqWNmtZrnv0npkspOWO
loZMDFk5dSSZApdcj1H2Um+lJ2ROtMogKeFj7YWlFrImKnFzuzjzkTHDu97RxZpN4rwAKJqwwBo5
OwvXmkv7M+7HqSfephwyAvK8lf5YQajKMsK/9rbHXjMVENk+teGinrRmOQnyVz6iwaGkgvxKZCTJ
oDEsGSOb5H8bhZzWKi42EPLwWW/OYLLLbSscutWvnE8XDiEGbh+7+RAupTrIRLTNNSHX5td+8PBL
rwxxnqf1GXddbDfqBZW3V9tdxe1HSiUHxJ/K3j1dl6Ed+UWL02uS8sHCmEAiN5raLTe07bEl0HnA
E/U+v5VBgv+yktLvT44XIoB8Utk+sBVbbujJspqTp1wOYqe58lW1yIVaa6n1JapAAPEC2eqYEIXT
tz7eqm/UFIC0qNrL8RGtfcjm4iQQ8/wSK3Q4G+igge0tN3+BuJ3f7q0NT5dFXC9UfiUfBcA8gqrk
GOotVjfclslBekcvlnt1DUbQ3raypXrEJntOd/DtThAIvmtio0jDh/65AL3zZnAcKWXn8/vP2KJQ
AaBaZS5dDjyVnSmerxlqmHMA0dZLm0iYb3ks5yt5xUQNHdBh16ZjgW+940j747Gj0BKD1BX1kVSH
EtgpzNvX0vTlN1K6h2oO8juTePedCrDOczdUXCFCDnaaCN5F0dbdVsbWHfIjmI9BMB+GkxKvpY7/
iFso698pzroO/T+DmlL8JRfzTajtC+1e/AqjVFkkM/DJR8kPjwwvW8xwuPi2TK5ZqkomwC9pT0iK
ecZIIzeswSV/Udf87WMVK5VDeaBQ9xuSKYawu8IzSNhr3Bbz1xHsxCE1oZg6r2Z80arlCNRtPajH
eHedtaAyjinrcdI9GbgfHZPge05H8cO6UjjxFOXMfLwYgDgTCj7x2jFGEFFxRfy2EhigfNtDf97N
H3Ji1H9TZdmHoRyNFo4971vMoAq95sJJDkFq9D7JLHUthhefcWO/N7EVisbd4FEffPS/6VxXIYoz
sV43BdIxKkn9oqzf2Pl9hMc34CSc+DzOo88F6AySYYf4NiCR0vyGq8vvDn/FPAUapRRIOsWrdxKF
NqWv2cYPLi3jaSMsZv5WB5CgAUYZQE9WvwWBaxd4aRT4+FbCzAMCQoD9ItwjCPjn+vvl9TkZlFHk
ryZI/LTuHbvJ0w51WNhP1eFrKn2s7NlYfkypf795oRx1DTif39YHW+7PK00ypP0bzdyfQgeRUFZm
VRIJsIKc9ECD6/7yBv/KI5C2zxdL2XGRmu0/Q5G57KpCbLdVAgfYZt5rH4hAiqID0dop7qQYPHHh
9sw3OMoPbPVWx2xYyL8dAXe96vuNwomx4o6+5mobAAsXDj1/QwfvGPW1iuuem8afVFWKr0QN0Y9Y
8UHLVRNkfVp0PauqIXd0SykH5MY1ftj4mrUnJAh4rN/HewHWCGzeEUGYe5NX8W4EPeU+UOgUQjDf
dWTmDScHedBcM+p7w0YxMISumT9x1puqJHIhDUREtspgdbvus3/pAM/tcHjbWMPyMeSImH1mw+jm
kLkYhvPf4+wGYT1jTN+l34NwZjqhJZye3R3H+7YSF4XsiJ0hWrUnSciE4mlNzChMnTWMINPJlNYH
UEEdKqV8Qw0hDUzcEGAyZggL9aM+tSWharjFQ5LhZQn5PYCkMoYDSAo/L1YukekyBYO24KxF/1ez
e6Sxv/CWNsNf6ogDtIx6hL+8h++bRgUUPK65s4YirwCcGMyCkBDqgij1H70ipkhSsrDZMaHxmgz8
IPr0yJx9YEWWlIo2vHuLn18smXGPgsPP9IfEYj4A+U1QU+F4RJ7rii1sOL/wFT7LzTk5KxPAT0pH
3ucxW8HiAtevbGj9RWCunWPeMe7FNUvNsyxPsxM6GF9Xw4vhWVxt6v7GpW5JlkeFbh7uNOaTpGIa
LlWASFd3hdl7yafnoj7VqCwwtRwmiUxue51DxhAvZjYuEWA+j7oKSo48Ro0l9jYY9RD3Jt9BA6QK
rv6pQC27hoT6w0fw+gY5hZ2d9mK1qNsxk+AC7WBSIhf2r6vfU5eBTcak5kU+Oh+G3mImEfWfpNsT
tj5Z8pJYjCaihZaN909lljXMeAuUuusKi4rG5l0/cXvcZf4YrTUX1rR2ayQKnLBtWOPajChUCsbm
N14db8bv4l9MYSBtDmTBUL2YTJbbMQ0l1uuWtGSULuPhbBO2QcRIvx/7WOFUfjJjYcCzK4SX2W4D
BhF14xm1Xy9zPVH7/jhSgXTT7qpcZOdZY7bJBV2zZD8LRIjtl98rm4jBubvvYp2YCjTQtSFELEhl
ZQFu88NB9Ouq8k7v8sQuKXnsUAowpQaySQeAzozvameLcY3bxPfSNaM9f40k1LkW7cIKKjDJjqrF
ZN2ebXvR/MsqVdzKXmgRK06DXyFirhFLKFrm5sgvA+neD8uAQbim5GtAbDbO77P40zEd9Lhznajp
1efBnzATA3wBIBlBcAr4bwkRXRVRJcdeS0yx1mKo4bGyYZ7MIN2FO2Pk9YftjbjbfFhW8cYk/KAe
GSkJA5MsZXhjCqAxqQ6JLk/r7khkzI7cE7R9H0M5zSk00uSpxiHa76Zqq583mBCj8qsEW5Nq9v3Y
BnQ8RRz7iCvs6BvZCY3k3Lmn+XBTE3+BhOvYjljcZLPH+K8+Hg2GvF94+D2XF2kc0rYR+NQuVwHQ
XYbwkZ1KwgOUf6jx1rv/R8FGLdXZN7/3U48At4xotoI9F49iphmwDllRdIr06U6I3EVDW+9xy/M4
WFBru346uFOnF+YUbDsMuGPfAb+lXx50i6g11ffEOmLhO9Wzn1gYaPIovMW5Kuqufhkv99pzS42B
/S7MUgxQvuZPZFAaTemm0+MVXHENTth5naEiU83x9wPYI1eE6b5Wzb6XrZcWZeA1WjB5h6PB5/Rq
mTG6aNvhMzPMIXt1p7CsXS2MJxzq78GJpWdPjW5h+LSEIyXRfBOinupOpuXW+WPFPEyjSGQZZzHO
c3d0RFCATWm+mVsVW/A8ue1Phhg9s6PGOQPOjhSITUDhOqEbRCpo95ZivBRS7Z+4ImzL14X7EAdT
E2tO+fXTBQRmZdx7wm8+zwZ9dK1EEyxoaTosNJl7oITsWdYLjFwO9SfywnmExaiw/RtjuStMNKjc
JjnCcxJ/KG3/NzQEjVuOi2MbTeXubX/+pb10fofbSGL6RXMzzRbmpeI19oHdnOLGyrvawNGV/Egw
YRL1SGOp07e+E8aqly/3PiOIEz5IlEwKfMacaQr4uLSJj6E7scAuIZo2jMn1ds3nSJdFskLnliT6
EQ6DwJEJvKrd0tz7Bjq6GsAKliOmf4z0uxY+wWAPOdzeIqDiyVGmjQyRT4GKrhUoml29kfHyxntx
ZSj4bNJdmVyNSuS/iRm1WZONCMxmPbL7XzEHohc6SaJgqYuKynucIU5xEB6VNB92fBE4OjqUmFU0
5+pnSMB7nlO1D+qJnqhdH9SQwvMciMziip3galEUwqOn/9AG6xRMaBqYlVcKIU6iU7mdfWO/Vx1g
wmftdQlptJTfAvGqqaKPebRqZsv7/ftSElwlQGsFpirL85UA5vGupAj3iIjHH8mkyHiOCRFWZaP5
n+hSx9C+XBMzGQz0uITVbxx5/MYX7LdWuFk/Uba5QAY3JCtMTdGF2qiEZntVEu0okBOPtIPQ8py0
7hIUuQlAYNemhUy22oTH2L7uKA2SaURfOKfTbXE3NTU/JP+0RQdSu64cfAzsTvIj0v6yTqzRomWV
WFA9hk81/Nr24MtS6nzuA+VUZbyr1DRYZ7fpZXh4Y0KFVLsKnRQO3b+u6xDLbdSoT9QhasUohBud
7SkHrKf9rnUE69uIRdfkGM7y7fpRrdkcWkIb0sEmZ7sGohMi6HVv/fM1taXebjhC7lsKREq6vgXH
TgJ6sDuPv/A15+5QcwPS27y1RBWO0qon+8GepqdsQJ8S+pQ7CIOXRf2YOad+vhndKF46vnidCDUe
cFHFklFxeErfZzKCmSD/HY8g85LfT/L5CIrNb0Kdec2yYdjsUy3zrrZGjwT/5kffBygRkeWTdQbj
72zadlUR0r19ygS+rfwtjmUtmeCk5jsWeAfnPk1mpO8gr+3BwtznTamJ47186nDIj0Qipqpc5qWf
p9q2icfcdXZRw+Z1+mUeNqQ0tP+9d4MSqW05F5cuCAp0Zhx6TsTJraYeuSNGV/qlLjb59A2qDBwQ
6UJkJ8yXSn8w87u+BqJ39wqCric807yKmo+B7BD9fNyDIJeakFHpguSPhh05oDbX3io54Bk+Jj5J
bBanzc6TQJgKpCkiNNbshR+1U1eAKZH/RSYbX8W9dNt9g+jd9DIpdujooE5Bjs4TGYdoyNxFRkEG
C4k/PWPaiCWfu2ZwjLYhCpr9MV6WlxI0om+HAQmdXHw8WpBY0dFIHGwtzhGzfVtN1l5WWKVCV1s6
jZdAJUxsz9mpI/HWmKwj1WmB7Q60AsdREAz8pFa/79h8AI5WuICSdH5ogIsKgqAigCjIxmF6Zg+H
Q01lKMsNVECBiY//iAaw9fnUR1LqlgOazmK6F2n+BuD1N/SeDrbQ0iIamWL2eeMXswFoltam0jOV
Lno2N5Xbhl3HSXTwOtpyMjvioOpT8hk11QGJ4xr+bN7NL3JbS+nI3YQ7yaZ/JldMGr3bq1earmdr
3uF1w0srEXwdeVJnpwVCxqfgT/kcXxYykreIDB/suZcxwNsj7h6yfYyC/Qpv9fyG5Kznkncc60I0
ftwW7BX38sDL+qgDcpKnmu110Od0Lv1B+BhChW5z1jcY4PpCQh9SNqmaRh/Xnb3asTtXVF1Uod5m
Izs9sIixEyBEhcu99F9QlZvBcg9uzDWaHjzEjUp1zmbTRaPHxUD5Q7wq0FjheVJq3X5Byi54VKy8
9VtO6eJuLKWs4PFk1L6uSBh6xLg9M1hoZekj8sYRumD93h8P8WKTIJC5DI05NTN4RCz8xo6TEHLY
RkhMbQYfZoKQ0e+u5aUBUgYp6OLeU/aD4rTBM89ui6gkizLXJ65Y3fRHv6q+6pPvLNOe8RJLHQAh
mBDe/d84eBs+h1wIBijRzO7FzNDH6pZrwYd3/tlcpe/XF1I8SxS3/aMyJcSlxqsZcJQjiPJqmnSG
nOW/BHakQ0H4u3zpmCIv35n0TSMclbNs+ws1rJTkYjh1RWpwhZOiEFzm+9VP/k5scCaRwtUme7Sg
3jMIEqFzqrQkGUUrTqSs463criyNEzu4zVwa8ZHHEkJT1D9d3NXTvxYyrmJauELoifBrWJMcMC2h
KK56qTGz4j0XceebHsXRpu0HF4p8MoVyorBqbT0oAWxDpIBmZbEN/NHGlaPWFmuBEEDkjPUS1evZ
ZzPaEI22yP90BqSnBWaI4f71WkTqM/1Y/uj9FWw4mU8kZ4/JudHNRtIQPANlD3MFPUMIgUOi3IBZ
bEPbbnWrotSoL84IQsXcLfJwD6P/+L8/gRc2k0t/71zP82WGAGi5/KmyW7mVN5u23uyaibsIHtZK
Z2/JiMZz8PFM0bL1yMQXyy7rRRmLtEjPsJZD94V3oSXSXdK1XwV85+hx7fTZeU3j3kLbjmaK35H0
g4PnVB4DvMdyEiAn42J5L6wiT7Ww9rhUX+BEl1C6pl8hWbav9EoukHEzOgyKbN8EGJZJt51MWksw
WeOUOQETLK4SKsZ7MGNz6YbHzb3fAY7F2U4Fy94qVLyT3KnAGYCKwv4GFy5Mkyc6Q46exmTtl8n0
83zg7YXn9wo1M0QJ9qcJaNyFmjj4PgbNo1CzEW3K9+vQlgnb9L2AzIDVM5v9PFF8nnvS54BGZFwA
JDA/HT/KJGVxfHxfwjM0FCDOmGjMZ9shUz4FgCKX2298vGRSqZfm64h05ep3/uwdmOa6GE1/Vbyg
QNu/BID8DLA+AzBxPP4EMU85vBANVlAm/B8uD2BhJXq+uno53M7s8qav13m0WQMEFgwmvuB/xQ1y
Uukq7z3NY6LH84rnT5yF1nN0GgHMZpLVDhcsNEjdQui0M+l9Cnj/Su/YltROUf5UdwzvSpWivPab
l3vHX2vBs6tAsEbIoS/s13y91Lm8KgZtgrfJvzYw70V7dl4jU3pMd9z3BOq4IYsQO2XhLtIe4wnS
F2lGylaIwakfkLtFkxuGH/ixIrkRrtfN9Wk4DTtPW0wP62FDCTQvp7hzRM1TBSy9ZHN5hCYl4tEk
rz/ZHytHNJ3zOM14GzbWiDVgOV7+MlojwbujtlS3o1zvc7FYWHf0RCyG3kWOMwK30a9MDbISnPYM
gXZHPcW+C8AIzi6y6VzxVlL3cs3pYVppK4zja/TEpXKX2/CZNVUTG5tL0qsE0CojNPfHNleJj/NC
OC4M1IaieBpiR2DZRerx8wTaBanfwDndCdHB+aV2RUgyQVkwhwnxckRJ1ekwCbtVXvSISmLUp9Kg
8Itw4V8drcjspiILLEBCI6LItg2Atj+PcibQsT/xgHGzkhvhBXQh1TxxR6NBcxDpyOrVQhIYfWri
AvVJjLsGwCUVe7ZTnpN+pABS/h0mCU94lGyYQ67k7ff7SojGcSstArQ72MqS6BS/uBn+giqU+V+K
Yvct/huNEDVAi5ng/AX249SeSsyWoh2CgJNqMIyFZFqlBW63PlE5Olsr3dlHNbmVmLsjGDv2vgVa
/rlr1TTjyxFqtXe3ltm1pkBPyWa3/0PmnsynwePOmWtJbKx+eN+kAzuDFJ9/EMsNDjUsgOOUFsf7
KTu16GB5tSEImT5JJ7cpLkd3SLX88eXgp9nKZbUW0McfYPZu4GsPJITWfvTS4qKyQ/rGNRf4rveM
twr9FFAWmuoD6e4pehp2ZL3oeJyAjD+wwAcYcklsSpprxXo/bPTbnUqFEgTE5nqxcx/hUoXGviDS
4k3ca+Xfh8w9VjowzhLmuEDEAjg99nEe8z2bkczb9gC+VDw9yeVUcNzPbn/FcOH8B+rRBq3v4YJ3
HnxhAPTsNVPuY2B/4yW1QOFctro/rHITELfQ2IdaxfWaHR+7m0HwxSossV31/lZHeE2cvSYEBPTE
RkJG9phIgawJUk1gmHMfCv+07h+gRqJV72WLga+hzzMOju9P9hek3XUjy+gvjGEZz0Tp73lAU9ha
rK3bRapH0xP1AFJqvmTvuHMEHS/mCNOdxaVu0KrUqReOJHm8fuTQJjVgm4zzpG+zEMnjSFB8p63i
EQGOtus1G6AEwRFMHNoB1nTq1m91mbPqd+9hWa79uXPINuavqRYUPQZrXWwM3KOzxKaB6H7xstE6
RagvatIezDknjVdo3/iek7tirRLkWV7cn4pIWRjKLa9qHX5AvvDhsKb6JtFRdVc0GyrFBViXHUfw
s3rr1rAI3wHGkJZi65ufqWJSVUmQ7yDzmdvWv5Pq65bXsQdPTWHF3fSKrx/HvL9/w/UR8DOzshz6
1rPkR7YLjap19A5s8yrpSb+6pnfAUyzxrEtmYlrQMM1vkBGLaG7GKYEj+kFOg+eSteMMucDE3Beq
Z7iQvrECOYRiCGWgyO0SV0ZiaHccmV4GzCU2yPKuaU0h715cgC96AC4YFTn+gIlvM3ckpY9y3kcH
RN6hqPfB9TWcJbudOWvi7QiXZ7Tklkc5tc6DfZ1SV3JKyZCg/CtRs+hneAgt2vvi5dC7VMQ3Og06
D33P8lZ2t5qCj2FvAZUXn/pwXUISm2lbm31zBw54ij89hltGDyZ72zWQ39WcEThXNw5jJB9uSb3a
BT4GbU9gDSmAlJEO4cumpEEeSAfFrUMlk9DFwwY/4V1hhwz8fVJJ7Mhx0i7TyugJ16TnS2zz5ceL
RqRWKOCDKULMs23L2SansHF9S4ZZqeEjIPxxDF4eEnjWpTuI5tlLIJC3Fb5SvOz6FbQd2YeBAwwE
RdsOpBXjlEPOUrlBUcpBkizUhHY3rzKRdNnIkRcoatVs6M4nlifZVb8KUXYUWZdcn8Bl0PVmfmi4
rvY8hkMiL3c/NgzABA7vdp58pNrVTTjqPCabujaFvj7a8Md7BIk6rayajfq3L2ocWThbT6Cwvb5w
JizsVPE0Ic1wpH0UxkF8w4jBCrdtX9/PPnhe+Jso7MSLhNHfMPCYbY4odj8hdYYCVXJcjymqF+Ye
p4EopJ2guKsXvc+xH3Fbw3C86ySD9kAr7KTuWmnOjiqb0sQvaDyAU9huz2KUHGlkC4dMWreY0W8y
VyfV/nvWW+1CM4bHvI5xwG+9un+R5Yh7R9+fNRUEemI2H3zZ/HKZxCcN81jtUyiXejlv+fo1vouV
Fvt4sq4YaNlTsmVMR9FXu8qgWeTC1O0SiYAvH7yaanrzZL4V0jO3CUQkICJajD+rprdEqnVtGz2D
DOXI989K+cHvMyeCtlNSXYjOuuEEFBce62H+ErtUkciRifvl+KIMcyS/TXsf+7tvSHGkGVKB302I
k+lv2BLaTxMX1cMKG+78ulV65rYrYyaMpLQZGgxxHFJDNJh60yiUZr66jgCXxp3BH2jzuJ5LTKgg
CQg1vY3/Abdx1zKVf102NOqRskSezfFxUPqWtXzrnil/IpYfLC/ArdcWIZh3GxHUYrKy/rR/VGXx
cwQe9qHSPfxX6yPxafegwS2GDYEMNXEZfqudpnEHRuRNETw0WXK4jG2eOc9PJlnzOoLxXuj2J3nu
yCL9aiXHcbrrfFB7XgW/TEidHJOYjAWfDfy4hSqUl8lxXGlgZAaDddTHf7pY8SJyww/sh+wzfALz
kCdrLVzV4FBbt4SMzb6DgEEzyNn5jHtxWX2UwZj+WG11SBqS9dVvHfKLHbv/IGXEuq35nn7rOMF3
dD7G46wA0/37SKtchS3/8pjaO7tNo8+XLrABgVD5KvHPxDkwG1YZg2qTLlDP1iNb9Au0/lk7w5Zy
av47kR1ZkaZmEALcnCqX6RR8nYG0MpOGZwI18N1lsSgp2WKGbuWIo+DlQz1hszbsu4DVUfj17r05
VP6bbS0e7znkHf1W/mIidDUKGeTybHQ50nlN0vl2b4SHDFCrkzecL1PrEmA71AEPXRryIdTcToR4
RbAIun/JMgWoso9CdH6miFzgpS3yRNmCm4ldDqSKmjHyKs4mIv0Sq5mlp8qL5KX3r0q3Q68CeW3e
IGZ4WNydvTKvp+Vwcw1zaIKOGwUoyozNSKaMr1XWGrAcZ2phkkk6yBzSwmZ7iXjwljg1ICgbinTp
ugNlfYE+kaxo2GAJBd63bEBzhYd888quvTNy5M+SAKHEtD2c0gnojefNbU1lI751YWv8q7UDSvgK
bk4k7AxWej2y3Q8JngYiipfmbmWUAOwJy/RPD8VsA4somlQ3eZvl50n65dGAB+94kp7G5gRu6leG
LfyjpNt8OaORnUfYwug4k/9GGOINoDI4B2PtpDnN5vI6+1ZbWGVw2GDBEJTX0+h8E+wqwTGds/wD
z71yz6bYdJ4aSpNsTcVLtsRzZ5lsxu9/6tqWjPh2cMdq+d7aQXaZchQsmJP8RziaRhFbALVApm0H
D8mEuXQJeiMoYdNOElnzDTciLz7xTS7vcqMC1dQwl3MBdCifMe5I7rr6L0yC8R9C4IxHxuNMNoDt
n9W1I2fdpg1WqJJAHicicjFJXFWIZR1BIvm4Qg7Ke4b4OijXTrY7HIdfwwoDbFkEzHwFfHJXKHOR
CaITejWrlFYuFJAt3nbiE5vlA9x2vBQ9HdzAF9VihkH/IETc5hAOHXzHBqYL5KQt7bHmhodU79QQ
6Qfni2h+1mbDBOLBMI13xDlq8wYYOTZxrDxJoA1qzdBRcBtVWKn5Z1adGRDdCFkd+yHZrUOixJaO
oICufgzXgTHyGxXCFT16t8Ou2yqaVB9mRDqcUOZm0sDNSViZfsMpcZB8dPzl638C7mVSXGAca64v
a3HWqoIv9i7RuxDCA27QuRZoSzM3veBwmhhUhWrpNm+4qk/frWtzR8d8flc7qqjQGCvx72qC6jv4
xMF93BHfdgH0vCN7weqOc8MDryH8GhYUcftAs+8alU48F7Epo5uyAMy6FU2m3Y2VUkkW3Ow6P8Ms
ygj5iWOt7fk/pGwcKYWAOR92XCqvdaj9ggnaiZUQZF1K2XUyJegJjcaC5pSqNANILrRq7jr/1DN3
XAjNIzYsolLcy1yLXW6mGrPnkEYwEn/NRYCIbKqiqf7oagZHuwA5hcfzWLCUZ+m6YVyCpUdffY+8
FBDycM7o6SLPOiROjT2GKQ8aaZqOmolBHmtFuzLkSnACZ5LYqlZhuGnZ2j+IbC7UaK+pgE5EU8fZ
9sgaTmZd+yIuhlF1h0vtdNebXs8oVpLhfN0yZGAcyaSrG11yFxrnSjhPBTRZvsKeHRHhHMVC2zPN
pxUWa7jQgc8qI+cpQITn1M0PoEAGsray51WJhwOf7a56ncH20P9jyOXYEnpR5nrmI0uBwKLtkDhU
ZJfwgfr0V4YJU6Eq6hq/qpMwf673+kDkx5vl+XQYRIYhZFqrWpsqGVGpEOxFoPFYnRJdWNDIRTv9
grqq/xhi7ixTY1kFVXaDWz0fmsB4pPXD3yizWnQN7K8MlZ4U1Lt1vGXZLEVjQBYLApOe4qPoYmFy
YJKj+ou3ToTzfXyJbdPPVU5rpnE771udb3jI9eIckg3nSe9BAfQhXIAAiH34Bk8dyDFHMVo/vB5O
IIeu2GjP0w68lJbyMEV+MNqVTRzPSprawDJqWnltyfhUE7pWeud6eiuVwTQHhZ0ltxxfRxlI6aj1
oCwGO1d6RwY7j0C3/BUEkGVQ+CRwTLL1TfMdfBs7oH+ZGCX+Eu8+soqBGTOKUlUTK59jnQc06c6R
FEPENHR/ILu6RrYOCV8GzjFWFZ0XHHgP70zsGQ4D8ZQuixGUEFAhJRGwX7x94OKGryqbJHMD6DnD
VmVYQxd5DDqhB6s4w1RgY8yv2WFxGqQFkJr9Ifbi+fBjPY+bTmMoHCAM+fIzd/648qiYe2S4UVbL
3O4vAZad0BrZFQO+clhtf9lFqbN2hiYa3IjG1TYzlx9PuoOUwAta4V9OwjE1MmJ+hnjhJQY6JgdV
KBoxcX8mXrCpRwbW5QqJBijp2QL5/p7BRN9M5LD8/GhtDilEe+ZyvdVY6sXu4PE8JPR4vZDK2NAB
5S2t/kVigoRCfPGMMdcsu0N+QNTibj+Og/Q6DAAevkGu3rZQtZ4oyfYDXgCv4JoEzJ4CqBRvFSFn
uRc1v8MwNeH4l1FWVBZmS3vbBVopHNVBc0cCVaaLyGdabiOUqqnaWdx3kOLEgzqVnE8ojjBH3Nnb
kqeqYd17We80IzeTDg/GJm2h8OMi99aZJFXDa4OGdLiBJ/uxOhQQhN+cvZpJDGk2W4koZFL+XAhZ
tRqkve/uSjGABGxDDmKxc4cEaoVaV7yvRA5iZvzNwTnso1gHlPLO9khfptEtuMY/cc4WK6vk/yJu
r0/5TMFKGW93Wyk8N/1XpQulOp0FJ8LA5ggEAgNaofbPqmCbrtCNujAUIih7zy3ttkp1vBLZRT9I
jUT9ZXJuX65FUhD08f/04uehaayI1meozJAKMrXzRpRK2Z0/mJLXcNVlE5o0OniNpbISePDdETx0
j6jbUyY/44mISDf9kZhBkC5rRyzb91ng4MFjSwZtPae3c0xgkboHC4OtbbfsvVMqJ2/IjZIpa9R6
of4tyigd9yCo9P6yX4DRSfZ3odo/U7Rq7TCSBiiffirfvsf+nEnKCOe4IVTnPCOVvehLJK8v0z4F
I8qQcd8vqNDuHqJo3Okcom9RZSvKkvHoXUP80R2EHFyglx3Y2crs0LGChCuxvZ/qBInsIcYmkNdZ
X6lToW5s3HSyYWRcipS7k4Xd61OsQpVG3tizWLpCw29mm8CwnVHM8AAMh05lMlObmkZ18isJN+7R
F006P/n1ecytGk41leG70wqbP0vl9H5PhDoFkcE1LCYlCu4brWO/8NrotMRre3kWiIJe85zGHSy3
CQoR0XeFBW14Y86fxuaIA3YzUWejLB44gZC2R9qOYxB07lMHBcPpXzQjVOg5DLKNN71m1efSSBFD
nJZIg7Od7nQ90DBVQDwigxkuh+QQx3TafPMYWARq/ZRlcrNlfocwBqKvRRwPXj045j9NEpaU6U6j
C0BAT0xUhhaDBErrLL2kze212Pd09yGoZF0mrZrCeOFVvGWwYB2yUp7Z1cVOAv5o+p0pu/R2PrA/
/Hz8C7lRbp1G3Ua3KzV3KeE3OVxfdijm5F1otwtm/MsoN/XEzPK+WJA7XbeKre2bq84vTfumqlmd
mMJsKAGOGpbSK7RviycLd8yydOmRlmpikZq4k+Dyk6b0MkrhAfPjXLqUfCqMUnetir/TY5/5sOJp
gIaB+7dTHNN/rV75j0luKdqf2lqSkn8nR5XYX5EX3pegkH2hSyAFhBNuPC8Vi2B7+RrJWVL/i++2
7PwsGEMGssTXVGQD1a/OslZazEofmUKO8kBNyzibSyUffonomO96Fn3Ab7kQTCtofBcJDXKZgTjl
e87EFNuo0OR7zL6QyDwMhidCmqpQwkptMNGigtBUT3sAs0rSs/ogUsQD9x2HUw978lUBKfTMc8ym
kquKA0iPLNKqGqTpnscA1459Zv/UHR/oymFwmdNF580s8ZqKwCATG/pbCV84t8rsxvSNRcmN4rO4
DP2lAr7He/jYoRgeYmdhSTm/x7GHhYZvul599f8wtEOS8Xf/XPIv120RbybjaKZrDEetAZ7xhPZw
N19qGJPaWNG8ILkykHS7KSFR6e/7/I5uNliyU3/FMUcL0CLs3VAQHs7n7DhGWoN9QxQcFYJIYnv0
d/vK/FgenfJadXRZAvZYQ9Tr2/mq5ToFjBOYlvQ5kEBiVmQF6lDJgn/nfGuHIE6ARpytBVaid4Be
M7UHYwdWKha+1V3dsTGo9RSSUtfHuNKexr4w3VSNpOf9fGH2xIta123tI6fsbKxbZ2BN0rzB7sEz
MwVJv26nXV1dCNxDWTdLRNkI8xKuDGdIhKyUAxYGC0XIn59QUpLkQthkFxBMFY3ACDIA3pjAvHnf
rSckJ9+xSW1c4VuFfM36yX3wdMUf/6GtAxZbDfZzT7dcI6oF5XDiAnchnfgHMW0zzOtXv9L3JfaC
8AO402hNEfV19n+LEG8/o4hLKhuXXT7Rzw9iVPSeoATw5D0o9eDoaQ3cErMhBmuXfPoY3uekLIv/
lz7ORyhJfCMJy0jMc6wi64AcMbfWd/wnRFYtLqUG2oaE+oo2JcjMhEvfEp8JHRIGxqbkZDFfLGm8
/GNr6THlMgqRy3yXYxAwuWQdHK3yNNEb5wBdL97ldj6DBw80i+qg2pZ5CrqmtYqJCsYVg8vsVf4s
BLVeEzpd4SYPy6azOgenjwTVr27n9amSQy5rUKLNJ/aKkn8BNyy2PFe0o8I5vjjuxJUfYyzyj3BJ
fpwf5dA+2cd+lm6vv7XKDx8LojUzRIgV3pOZUN8R0Ctf3ukpcQfR60PAmpV/EOYlckZe7rnqAXK7
y5EjFPk3RlW8/qusD0K4FAnYt0XsIXOMcf7vgww89Fo/VxCU+yQY6DjZbgzsyTLTuh2jWUPvjMDv
gdeRGoHiDtID0EMi8YIzPc4QIv18yQOcQ50jKcvwFNyluDemEhP0lKUEXI+sLPmFl/888z9JSeaA
mHK2QkZtRYjvVIjgq6MbpnerJQPSPdukvk6GbdHY90T2BDzTlK2phBFDi3XzQwc7Yr/+mJ+HiohF
BeUB9qo6vuwI3Aczm7Wr7espsfImvbtX8EgAyCJoqmsUzjZntJYI+UFI16/ttreAisWbTkcfcMnP
XrA05H/I3ic81xcRVOs1XQB2R2iOJRzb+sIaMloiTKvEcnxGoSOpxeeVHaCb5uu9chjcaslSP1Xu
GcppPsZtRT8jmFWPtfG8keR+mAE/Y6ApmaFPRL0KiAI8OYUiigF2Ilzni5bDD3iyasufU9CDQ7oZ
R1jtPUIvCXxqH1zAV0Mcqf4eSJvi1ym+zMprmx+OGFEFHUrVx1O3SBVyu/B33YFPLrM6pY+ynlTh
I62xaiHyzM7SiPeDCEsxnHme6qu+ZOR4rOpMG1FzbO3vQMiqX0In6h7d8TnsyugGz9lYrTGUe1Y5
lUDZOXsjb5dVaQOhq7FYZZJu0JDht5zENOSGOsJasRUV/AViEY0tl4U/2YcAbi/FGlOlQNeTMoQk
RCeQ1ILSGqxezu4eA0lU/y7SKzTPpIaxBY8+TdZ3YvI/zQ8ca2V0xsi0Mn+DFWCZqg3QL2V4Bdt3
eXOsgLHdiXB1C6luelLLgokM8+4z64nYH3QzKvUXfZSAChzRwaSybwPSJea4v4x7dtJciCpTf08f
AanX1e6ybYF83Dp46QhYgG6E+0ZtYBjBJ7yYb07s0v8TLIbzLpw4FNbFN8FIXqV9lbvGqUgLp64W
1YWD5BN3ekBE96gI1QgJJL7NbU7hv3tuy5Rb5JIRiVzWlP6RUUQWOCuWynQMv2l28DmvmptbB+7z
WJABLJfKyPyo83gSXhZidhsNguzHclA1EbDUZtWJ2TWVccLvVEXga1itgbMdQR5+XbzW93lgYMI3
pQUPxVwgcqb5ixcMKWNR2DPi4DvAYOMlnxQ80LI2FvJqf/PowfMcJyDuu2lvhlH75pkYCuZwv2Nk
E6ZDIvGpad06JkEej2ONqayFTk24BoComebt+ziRjG2uIwHqRX8uhdWrtEcbBjgSwOTm9TW6zNwt
l/v2tecovAO6BtyQKyOaa0+OXrrQPjpV0k6GFqktVxwCJWXJrlRvMtWGXckpczxYWs0RwTWMt1/S
dIZuiAGkofhMKqnz0q5tg+WEMwKuzyqeKATEdscXdL6BzSqE9f4uKILL2ceH22P56p69bjcaeLJ3
EDT5BuhqQCT2sDdmqmRJ/rISgqYCb8nB8oRJY0QP83l0IsJYP87BCaBBx1WmNM7BTdKpdnhvKjuR
9dGSR8ZBzLCwCOxnTr1cXYYMgs2xqaXk5DTpVxX0otNTpX6TNPsOXiczvF13XuqrrKqP/8Kp/i3Q
IZYUq2FSn4M8gj81IfPl0P9fqOGc6npV6YS42k3DXcwJSxa5dREUbz08zwQ8DKh6XD7iWC221bnR
MaeqfhTZq1RRbL6j40H0iz1D3BsABFF5NkzTr8J+NNztyJVbhzqr9GMTBmuKCmMFOBA5WAJ3C+nv
CFnslmYnCju6qQyJbomXPZ5WZZf48A2+estBmj2IGcK9P5roUO8dJB9/2rAumdqW73ZX+kkAYRjH
Tayo4bTpoSA0fpq6cDGILLBFrWAdTOg8qYXZ58r4K5pGikXev4KiHVH2zCg7QQCjGWTjA+1tF8LM
UNgLt9UHB5odzQjEy8LwWDjdIqCGwyK7/+zCrAUyIDSCLE65zuQI+DlwcgqLwM8RGrHAW64KD3mh
kEylK7aVdYfOPngcnMw798RGTYbaFS0vSxtJS+/m3Iazqq1Bdeh2v3CuQ+weReG3uBsIK0WrZUyU
4lvK7fxgGDhGvobG8AwCMUDcldD+AGU5NHstPQfRlSSRBoXdvkf8UQBTbmsSA58ktfRVBNPzP/fd
pnAcqJtCMPkdWH3yr+eongjJlUldT1uMOLpmq+UOMcBfuvBoRBYcLaQGF1VcUEK/5GsFa484SLd1
QNnBTELqHCwGpN2FQGkTkHqW14FmZbOn8YSP4LaRrZ4OwBwIpz/jR+pbsKmeWe+PfsWUwD7sFFBs
W8dSD01EJZAw97+WPZVT2KRcpNkNHoPXrKeHEZiWcQ9sHIBqmmS6FcrEKHxsI71wqyR7Btouq0k/
3/5Z5TyKiYm8zYeKiqkWVO0BaHCDbO6YuFI+Y10eVhEu4oj1LpLQzcmDijlR/raoXRvAM6bB6aM+
B0d2q4ZJgM3DFDJLmMPW7BZHN48orBJt5WsnClofVYfUnPGRH9Zj9q/7f/lKExYp1wYocLSEgO8q
Bjrv8W4wxYJQy0VZeEvo2JsPKnnEaODRAGTvFJpGx85eOmT7Puze52+ToJ4zDQxetpbnc3Pf9roG
xovUKMDzxHxevEmP4n2fv/hjw35vGq2xAbNDIQoqX2jSK6NQ1uHWv77bv+FvXdEs/XqFhlj2a42P
stBTTjBwsNMmhAnkZnWV2WNY7AB7dzszlF2i0NPN2XgBt0HJn4C1L0NXGB2M7I9VBHw3DkBVHvd7
UikBP1X/czH1NYsn3AiVCRfjVfWWlcK2Ee8bBVDHgrR1n+aCBGbqrQuOZ8wDu6LrxDIdGa3N9Smj
ZX8RMTm92/ppoWhS2PBoceSBWUY16xrBJ9M0FYRygc2fcJ71rDcisFTl6KUQwZx23TzZyfATIoQT
Sd+QwU8qCWl3NKGTXXilmawBiP3Z2Dq70TKCgPTIdLLQ7oWbrNA5qu4xSWcEejALtwYl73E5dcSO
aHvuvGZivVpT9vXvjAkCh6uAQpkDvacrYRV0a9+qQxM6Nrmg6zjKwIufiqUXtn5791GUA5s3GniD
9fbxnQ5n+TfI5PtH4dRp8Gk/U3o4pqzJWiKlgv+ThxXC4xr8My8B1ovY7DCx+8FIDWSm5sOCTUny
FitPktLXfqGK2OtPbmQyubTegGRkeUvpmceu3AoTETvJb3wT7AuA7sDlVQbK9EBfo3bmrFIqNTml
3p/dazMpDCSh7hvdQnM/XblnhhnLWXmEzyWzX3uQhvzN4c8r3fjoU7Lcq+tNaerNWGmGeqATLVzO
7DXAiTMCR/fl7HYfHakteq3Ysh/If0DLGwskYWCWmCTn/lJ0X1WUIQeHGLbUR08TwvCmKQgkmSHF
UnvFwGRwHyeqgTSP8VvBoV/DSKKNsI5T0sWwPF3spMusWGm1C4daWUm/IdkI743jo6dHmMWQv0sg
cJfQfkSDwsPAd7GUERjHFAspQFIo78LOLoBAUIQhWAfn8aJ0j0/Kox45tJ290MFGjnabyaIljYnw
mnmNc97/nJxD4eKT5t/Sm7mSj1vaGRpc3yWJxsxxM7Z210/0/MjLv4/S4W4HimLPHPiT51ieNGcq
izGzrP/WKOqTED7y/TYOkvdxrZAyAZR0g0TH5uiV6gVqVT/uHLq9W5bqo7LpSQPQrInoReMw57N+
98I+tBBUNZ0/56Ay4RzQPE0uBTUcX3gVHiD2nA5xQ6ZsU+2+HIyyJWjLtBNQBy6fjziW+vH6JjqQ
n5tz/3MuZ9uX7BlQAu3Xhaq+OoalHIQVMTiZqDbAILOuPCBtJvLzwRV4WOlKssLB0LCm0JlGSbHH
kp+RlKVyCnn3Wf7u5dnO7er3sRCn2mY4/J5slBhx6VpYCKiu8gNSzvaTrGi+f+C6rTcS+pt2tOga
h3aYlXpVFSGJ2cm7HNaqa70044zm2w6PjX2IAUK4EMmyy/qKNCtzhDegm1bt7W8x9OSz2xcO7SKt
RaSDpkAt/N2qURIsVHFdcqRaRqt3eHCLvjM1qMDo1Sw2CeV6eS/WwWOCIu1QpkPCBN7umpSDIjXS
JQlxO1AimUoeY1hHfF/2TVmjk2Ss8vpIQm5E67jI9CJ41qquGxOtqSXczQuDJ8o1ncXhi3xofIba
N4aaPqJOFS1Dck1kL7iadcAGfjfGxgHwvp0epN8gYrVmxfdPuF/FPBtNftR7pvmUYt60Qh9ifmDB
OU3fRKqKGK49cUXJwipAgzE4n7qkZU7F77nsHf3w947P4+PZD+UOkz/dW5SozB1Nf/8YseFpxubz
gvIB+KebYnevn69oMo0EUgFQQ9dsPTg0xjQ5Mtdi4gETYgvutjAzb90Knk1D5LJ9zCWSf/7XOEHH
j5BnGUoRyeaKHcd3hxfMEQ386dOYeR6bgIpgixT449gMeN4NVoDZ3SDQGvadzlfwt8Um8fYLVNy7
GF9wQtZnkzHiKm4H0oKeoXPylPDKHJ0E5k6iwkSnp0ICt+IqJ0R/JEpBz2mELLNUzSe7UepL+k2D
YSzHypsHAv8Q6nlKq5i8O8V0NIsRjawxXQSmatSCQHNgzgxeeK2wMNzudDiIFNEfCqTC8vnUcdMn
Ld+CU1XzYzS7g1QmhCko4dLT6tL8rbZJSHRdo4LrSPdlNICk4UfPE+vZ2UVQoJWoqdllhGNnviEc
ILku38xEioDzBq65LQh0XmwJKuiyGkYmrLi9CEtthClrO+QArgI4gliOj0PiOB5lBBGmlqLWRuB/
n3C6emr4s1An+3sv70W3Q3Cp3dsu+a17365bE4uI8jf7YeOY8MQvdzgh0oNYfRfAkMVvjP1pll2c
+LxZqvSg40uOs0d18hWmxVFhCX+XvJHw8boZVhPQHCzV/M4KWx6mBh90vn1h3VqCfQ82SIq83rEf
Ml+v3ghCClW0dvZitpg3c8+3T+r2H9EPhTpI43bcIeC/djS4ITv7kVVTW+poOB6hoCL5zMZLOk8d
21BnB7X3L0KW/ofSp7nVg9ERev86ehW6OgadfRoHBa0fVNAomTxFM4GwqYmBBA3dXlS7nenJq+pi
nGgqlwSFjO4UU7XpEg9QJPo8OoANzaow9iUe2YhcZgQnG4l6kVjyy05mHTqfkPI3GcGfU849ygjF
M7z9TpHPYonRt8vNyFnIW/FDYPXJpBZOpy5a7jDiFF3A6YWqIsmrVuYXhkpZ/2gplbdVecotpgAt
u6skJHiC5z+3OYzUO2N6K5gGyTnWRzNGOAuJfjU62LEj0hroANhPXLtchj9jcysL5HK/3fMe6aaJ
BmUdDvaY3rCFdvZ0XP+dJ3HkH+BWWaOLK5yr5dv83oOZ5m2ekr1W6eLwFIRKUp98C20kGPpa9g5x
nnTUGhvOchH6i9gQtdoacgnLOzPuSvy1oNZLeWqSop3Rme45JthgHv4/9wjmBWGfTO4jb8Y5e3sM
5I+uXqept0KAv7hzQNhbV694K/mOWqyDm1bhqayfvE7wHTZbC8SDOSrSPOLxjh+juJVC8HcKNpyl
A3WBQtw8AZANZxOQc3eNEjYOBauN7HMxnMAF8vpj+suogcUQ0NDkwFFB87eWV0+7Q8OS/ZWVXn+e
2gSxzZbDHSQj6DgHT8yTj4pBTe2/kAQUFSC1/Qd3cDtZa4zYi4L975fLNEQ/bTUcnXol6qN1ckP4
xjsx6gv3p0mwAx1/a8k7fTQsaQeqwfyQlNmnC/Kt42J3cPCSjfcI/4F8BGOjbRjksDvKI7A38yzd
h9QsOEqm+Oy84ZTrOaHbQu/ZYog1gkXMXchJF7SfnWR5nVB8EwVVTeAEARLPJSTXONIMEvResBVP
ZrDUVEni4cPANhwwCmTYEPY66a97eWwbcgOWdDA96Dhd06Sp6T6v2maTWvE6q2j1S7IcBIbXr3UQ
aCE6G9XhoUgC9hLACr/jcuwaYPtwt/yaLzYd6QTT554HDguU6CN7Xo/TlWtx69CvDuKWyqhIM9l7
xJDAHQGCpfdRfD1JeeXeimse77zY5lH7NxUpFAsMcftSOMqBPhn6b1dkO3HE/segGFwC4xFn4ZkM
RC5XDo6HqrQAQIrgnOpQbdTZjsNqmwiWtNZKwBiVUJlNdZ1F6kF5Pzrzz7Y7ne9manQxqSBxcRGM
6jluoN7cGI6w3dfXp92gOw1cIFzoXVKdlwkwTh57RRH9o3F8ruAzFRRoLe8F2UAuZzDXEteihajS
XMhxfSzVD4JoLAJQ2GVVhDgNmiQrAbz5l3JOiTnwoNBSbAUNm6922aAcplWJE9bk/qrsqa43F4zs
w4dGBnO+CqQKuqWO9W+dbQQmK3zyjkWRTDZepCyZZF2t8W9iC4frmGAtL2xS0MsNfYigciirxCCj
HoHNGWZMal+/JRt+ejAJ+hAOtZb7a4s5+pvgXukdXlm85HTV9G7xGHXs42LE3c5JMOK0WInoD//O
yg14Ymtv0XDKcUzSlU2eMa9AhB+3AYswZr84zDbZj0b5JDBo1NNnNi36rAfqbmiheqMSHrehUhfO
un0Sps74AiUSBFSHfDzE8Ro9aSHutZHo49Do0nXV2ly5n/nbxueEAibI3v5e70ffUNOs3FT7dHvF
NSKbEIKHneXx5CMg7OExtmD+Uqrsjj+ouXtHL80VaeF9swasC7Y3IsEVYTluDYbkoMvTvGeBu8G0
wiEvi2LV7RJx49h7cHwQiqHuv0JewsvnG2UY3XfTMegPYIuZq0uzNrWCcrrkFi141Qv3UI8AhM4r
SD5qf98nCcY86r0OmHMY7T+uX++ZuNGih2207ByVTXzPdZrIlIlSbCicFqycUM5DwHI2jFSh6EH2
ZmD6yTDLodssWPNPaLfeeiPD0jdrThDRPJ7C7wBvAUujxUdJr+ZTWTURW96W1pzVxSMF5b3qQjPe
sIYqdDSAWrRWk7BWz60xUL+YoQWU72w8hQNOjJ4TzLeOjEcSr9TG9OQb2egpKxY//7zoDOJJfxrE
R5cWVqytLPi7zVYWeHvVYiStcl44iCTWifSj7lkuc5xJegMp6xOchNekM/5sbSiYRO2x0nAbrMWV
a8X/Tf4eXaJhUUN510q5XNHhL+P1fc/wl7lf0GRfVaYW+D4EEdjdVV8q+Tp5/+sGAsWMmgskYR7G
DkANswHKqB7aOuILdKDX4TsWNVTNhq/JnXwKPzS5kkDVFO/TBgS1SGk0iw+R3qaoYPMpGBghODat
D/hELdZOXGjmFEMviTGV6tZXMlcZdW+FtCThV19M8pD8faz146V7trGe/ujc4YRlS9RobkpBgs7z
js0y+jbDiUugN6cbEw0msowTVehUMaNyHvzUP7FTniFICACn/O1t9CNqnpjUGgS7eOzzNVoz7m+o
X1Je6rnOzWbvkJtAAT4e2XGNZ1/AVEgOO0ZIEXO+3ND8u5ftJDtQsgfqyQjJjDV2qAzA2C5oVmOq
MBUzxapY0nwqdYxN3v2bk6Gw8H3TpgT2DoAXTNWiuGD4PJQfqrUGkWCh3RZVQZBcRnIWlkILJLa8
oN+H3Fcu6tSQAL2PTGUYPa31T6J0Kl4AOTyZT0RdK/gzfvYg/r+D16ESBCwO5tLBkraXLTL16LEI
lWOjxAWcct6AL+OOaa5MDfOc0nInK8e6qRiJ5236xJKgSBrzKqeTIXaXZD4VyuhC2AZAvu4vJ2PF
sI03kvzLXcbMUczQ7ZHhcBJxV82eexdTLI8TczHSZwxe/KTEXrj7KdxHgsTW514K1Prboi+1qBG0
zN1tedNnpvw+DV9DCv53yOnqVX+A2WY/dhKFYg3H8+fjNbgb0MChWPfn3ddsajgM103Hz7zcYomb
7OzvdbzJbnzSdVrT3EjIjRIsSTwd326YP1UHJW15Zxz+zacJ6hYUuH7TL50A/jHJadOvPXRuWBgC
59ZaSQtMtRHOKBx/GIXWOiNlDm5pY/z2TrJdD2S9/pexR93xW4NxVFXRMNBsvTgNpHPt7rPTEPqC
9xgL6UJ2H0haOEk8RLxJ32rn1CjEUvHepJWawOm2R0oaOj6SuvC40t2VAf7Z3OopinwGMM0eLHdz
WVKr5NkyyU2JeLJW3lQlOGQH3PxBVQp8l8C7KLTBuLBV4EGMi+kvSkBFPxxAmk7jnuc+T9nIgX8i
4lteHKab7BoPL/zvO1m8c652sLrs9nzFxmDwr9MEM9HKMrFICpacFAC27tIL7olfNlDp0/hPanrU
NEeXKdEOA7b7AjddzKrEnOV9FuswpT141ifcQO3Bm5n9BLmcsrcW4F/KRQtkQVjMMbLPm8/R/g+o
NWQCVMufUOensiWvjcynDbFZCvCrDNef9WJUOeYgYznunsDHz8JLYArfit8mV2enIgU+LOayJaQ7
+2JkHnqZTm7ktAuBmQ50yu3cPg/kop10m6HwjnjA/T/v5Ae8ISOHmEqPi0IkwRoQ62pIUPzMhu+y
UUNV82yMGLv5QmXWTDdKgP9Cg/OBtWW9Rc++kUu/p+DJJFhmUJayDnn59lYNZsfILykfA/g7Lb7p
T5Hnr/du3sFaZAWabiPfvYKtORDoPEoPdQz9307DwQE4DxeZP8HQTXas9VQSdyqQ5yTyyCOR4WLm
9QnrhT9QjNkvexzCYxstc3+xZiMt0VfWzFt3deNHTRo8DFruFHqYN82CdMsBUQOcvaJZVqDXHIZ5
JRoodL8R19ERwlaNIiBTauBQUA0CXwzhPBFc5EinZB+nFvdB9q0BjWE7OvlGSUiN98uckk2LY4au
YHsY2mPE99sW65Pm9WyDMNYqz2Voy7tbQK2+h1CmmI1mG1qosgSlyhqSyTpYvClpa0ysQbFKmP9J
8UTW//jgJaUWCyuWye8l+FLqPWtUadE8jIYK30AK+UzxpLMPd47i021iSAgwQZCYJlo0NZ60Adw+
Im482x21bgXLANepix8TvYXaFL5Z7ZXi/TJaXtFxBmdPGKcbg8nkqVLOpFY4RBNytnrFga3OSvbD
2OEkn9AeZ1ifIGcKzgeDuKdP9Mur5HdK81kXl5DcbgE8EW8YlstArl1uKMTyIOxj5YMTovnPZn3A
HJAYxS5uC3+dyRObhFuFb6Eys5HBj1d5q44/58v530hWryvi7bSZh1eSFfozw/ozS1MZhua7gs/p
p8MI2W02n0jWNQxl3PHTSWq7foIZXnt8q9aZKqw6q5JXodt8hWw76bikR27HLtnKIQZc2r7aQqGm
yIVAYPVfVL4hlcs5GnLrna5HL3ajgS1LFrnB5RI+Oq0iutf+Ah4kyMd5Up02Ut3PfF8Bb0vytkBo
8iQ31TZ1QpE3DcN/mhJurKJXIaeBvKZP9MhudZxSi0UlqgkEnzTk6OROvX7nEP3OLMkX3PsxAfmL
e+wB2H/+F1pZf8D26yv6INc4x+/b8B7/EmPpuV7d5YS1gWEBy1t2Nrl4r8uDDHcaFw4WAsoU3mlf
jCqBz6dow7x35Wia+j4CQxvOjz3eZgAE+DooUhZzKRu0XJoYm+KOElw19tOvE1hcH4AHPXhtmr1p
Jmrf3s8q/yire02fE5kMqtz0vJmshZaDlor7PlG8G5trQChSzITwjUHkeebUnIDKZHHB39rd8cNd
nt9AKOxWYcgeClXWTUjGuCDQuh8FnDXNBcu0wL8wC3PCRDAoi0uNo1Mvh0zEtaLz/USaH7OZRt8T
RYsIEu+bnJTTZMCIczND7Xr3dYs7yCv6IVP+6+8obATpQ2cJCuna8X7Fy7HHZKW6skTFmlg3cD8W
vPBoEHSJGRDDlzQTsO6G/wUC9ciX3au5Lts7Pa1I72wzqGWdUJgY3kDHB90wNqAknh8hRIQyFjxk
C7KNzS++2JB/dsxGzh0rlzymQ344avRq4gD9Ao1RyGNWKRj1fpb5AsSlsSBFNVQ8blZPuPMLHJg+
XjjQKok6bVbUsBBGYLopqF3076LeEbxhE8wKV4i37y5pSiI9kdqDBHMzpznH8sdAXXhMAXzfsieV
YJcmFW644OrwacUKAvRekvE04hEDLuE2znryDjTx1HJFqO1/GVAXamKGkgI2C/aergNs2s1c+FoP
2gAe2o1BXPdoPpmHBBAQMmbTMqrVoQ/RBhG0Y8h3q+OJTk8NpVtoZI3tEEUjlUfJXhJJLoyadrPj
rOvNNwJvn3Xs/f/N9Doliq1Ws6Tb3IUvnwR9hrwPkmCUBwEsdklJK4oK1YRD5CiVcqDFcQs8fDm4
cc9Qm/RxP10hYCj+nAhmuu+390bG6w8kLAijYbPfp+eHcYghnlMp35yr4OY+qB+NACdqbEMXKTYd
B9Gx9gPlzcAs+Xt4OMuycEWLy7S+ivMNdwZxWmaaNAmNWvQoWHBbT1F0zoo7cNPZNoOPa3W+kEqa
dIXRpDtOdtppPPiND8dUfDolOSgZnz9/aQftSAUb8kmrg6tzSYH0Bb4p2nlsnWNmZKZ67YM4RBcO
jA3yvcxvrkkSIW4FvSeSls185TSHpWY8RXny/U5Hkn3wWMGLzvaE2hfgd1WtJTNgU7s52x38ozJD
YOEMrdUrmB1aruv8TN4X/KOx815LmOa2penBe5mnGWMRdhSYRBju0Xvs11Dp4WpBUrgVAFM43ydI
5cKvUlusv3GHE8vwKrGAgIxHIg7OoFs5hMmzry3aOVxyPhBAzJGOCgA0ekZseX49oZJuKhoEWLh5
OgfK1EzYIhtHddxflzZFBySi/99iPKrczQ6PVQ5XLdwc6JJsHDAel8GQjrNohU6PBGuQBouPuWDV
/QGUf14LFNmT4Gg7J2fj5pEd28g1YpQgslkpcPob3EJuvCb+2Q6C++IjYvLfGZyR10pxI886/dzF
zv6r9jfSPrDyD/FyK8dNYHmWDPe73rSMldhDbabH2SUHBpBLtTwA2eJlu0Jx0f9Gipx4gnvMltUk
dDTe7f2bH8AVUkwOH0Mcr7/QVXx34KYcz2l92dD9YHle6AOLyIzU+ouepYYCzTMLJBA+eWT+3hk5
T0PvYjP+xYOh27k+ZDnRuBjWfUR+Ip8GI+cJvT7gW/ITXN6fyNezG4Jhdg1gDbCtej/95L4FIeRb
ROKgyce3Q3Oi/YG2ukwiyZvN3Taew++KPuoFxypExPRlDs1q7BPwIsVDyCtDarqP/z3AjLYz2PsF
RY8PjKLwmbeP2tqi9VZOUQazoWE9xIqXqbtnw3As2EE4F11p8FH5rBNgDWbFcQdHEwu36TB5SOQq
aAEa14q072WBOmULMJ3iXonCTzFechTHQSL0ZB/U+yGY/2e8tZ5hWjwhQcFMaQnUqofKgiYeSwoz
jZOILpflExVxjsBCJQ+lmZTlU9894lG50/E7m4AM2hh96EPxoXhnKVzGktoYX9UnO8GgWaaXzkQl
mUm2apmkHsrRctLKBBUAuv2nDil7fw/qX7UDIbdmoGO6g/HiUYJM4tPVZQucyhTlfYHaSUcqbtYO
WCeYRVJ0do7Tdbbs8mOIH45vSpIfpHIMmGH6ZWYzb0wqQR7UYAteJmM/FaNQtdQzOKGEe0O6bto/
tgDEvJkBHGlg6YdhMKqdqXT219Nq5oHUnRXQAYbRyDkmQE2ZGWbUnaMryDjiCxwkaPJChAQWRSnX
8m9XQPU1S5SLgknopR/Pdy1YYVP0WnqihRBWCTKfMJAg5vdK511DSbqH8i+fmlyIV6ErvYhjUcln
iLFf4ZDvzdOxLVyV5hHt8fMjj6MBYKQqZNLuM/qhBhHU8a5z9ob0aCxdbrE3GZNHYoawBeDTqEvW
XXHTGlVNyHJQtNY2aeZ5KFre9ZzWVlbJZvPTvU6PjIaqm1Y/OjzP/St1IyP2sEfEoncdYIBqmWVe
sGDCWE0oD3JQ2vEtlZ4PQ2/pNJar3oyjaP2eIZ1CPY8W0LiE9t3VTgQBaeqMBKCDJvu8QumVIRsG
CXs8Lse6dSjLfi14tDdQaUozl/gPf94qk7f8shSr97yJObkJH24LTr0GU6cIiidotXqC33cxDMTN
4shJHCTUiX1QZVpV0LvvHsNyTUVkdnEaolcoe5yJ45mmqNiOM5wCyCbYNWWyUScmSyWjb45g/xqD
ZzU/LhP4KldnjLyW1dwLTXG9hT1htMbGF5oWXAcaRDTaAffMJN93qxLWqUS6Jfh9BI6+jEpgDstf
oaCtLch57bGYVV0vbZqRiMuDVI2hgDp87mYxkQoc5J9Jk3jwhFkVPI/1EDhtrKZvrDunDoXBWPS1
MudRRGu4PLXJGUbZfiJCwWmz7v5J+6YdsJIbPaHheR6wjVScn+eY0CGHCXGrf6wft5aZwR/DH48z
+2s0Is+JAYc5uPvtGi7o8hNiAR6t+jfp1iHzsjwUms1r8/CMoQGhiQEvyKxjmgiNFx7T/b75OZEW
UQIJf11ufmuiXwCDLHtccglOuiFz/dWIXsilEYsAF8Yjfbq6fxstxMUcQSwAjvWNYYldAVb9sTzY
cOoeu89/VYrWVRNkMz6Kjfky4oiygUFzMV9de+rqM5OguGT0KVgCT5AvoPFxBTQfJ4CdBbI2Nw9+
JLuMls0RY5/ZbClaqGNQTUL/B69AbfMbSiyctDfLailjy2QDjWwslIEDpZ4PqoW5neNWDUkNAJAF
629VNCtbp1A9xCNxwdcymX6W6PZHn4XQRjJPEPdyjeI7mTy/oOhUAzyiBAwy2AgCLKwKdbWOvIId
Qym1pKHBtgxz+XulfgoX4EbzowKncVI65qUKErsMZ5nIQwtekxJQ4qrukgMG0O2/hHvG6yYW/Vho
QodZiRKY62vVX38UfLz7NS4ZcaX2u/eIHfExstwb5gGphQWvIRFWymlbXR1teqDJ0J6w9ycwpRSy
upOfKW9T/IgwnmCM4F3ZiFbQGWXDmgTPEtffOREEIqX5yKXqWpXXZY8eBfKM8z5CYDJ82+adsa5j
ATU00bdha2jOtWNHB4YxwyQFu/kEmQHsCp6oo/W3v7cX4oSUaEX+89kWz0zFKnk/ximgsTbEGAIn
MfPoqMpsV245k0DtBrJoDXQ1LtynDgCtrAOuvs+e8KLnZusEmyZl2hg/wk6ZkkdYUSFQ2G0KeUXy
2E/IvQkgBUzgeDY3Ub7xSwioFuuZVCWeUMzvj3Tsfe265vtxTtd4pIIZD8POAoiuaYqe+GCYdxCh
8i+W6ksRIbvojH75P1a0Sb+FW0dkzZmBJxo1I9mBS8J+fdrNd8uOGTIWPx/QlZYeuVHdN6uVSfpC
0mhpAkdBi1bEIDs0q2sEAYLpepRSg//pqZFl7vHGiB2axkbOhit+TmJpi40veHQ5ge18SKRrlpAY
wm4TIXptGc8D5sGi/pUT3W9BUGeXarGO7X92Eh2c5rPzDv1p8RpgBwb+xPDaA1W1Wryny/NG1e2H
ibDcsEr/S3YwQf9aMNgrdkiX94yvqMMlIlE9BLWpTO7KZx2Vv94foKHoDNM3ZYDYgZxF2Ej4c0lY
kwYgiAMzgFe6C4CVU335QKHihHVtnsmJzeTv5CgQCAaYj8czgol98me0HvprrWdll1OL252Vqy6r
pH3E5LIXLblszyk/fkt9E/9iGkeqa/4IjL1ra7ZTPrbqHaPIEtXOBDUQGj8EJSKALfOFCaYvViaC
VKytLcXDLiShhad2btEHzvdDLv1BKlMcpUikBh+MNoDZKS4Eh27v+qtuKOVV1y9RopyZqRs5icrU
DH1ED1eWbbOMwjKJYXyvOXVxFrWMY7MpEkneba2HPtHVB69LTn8sdYdtZCLL3qT6qvzr/wVhpoPK
X71MnbwP3svSGNZ62BWulkL7QdLOnc3g8IAKLX3ID0BzGZ5Fk46OcLthB0M2hNuFVN4/J9g+ScR9
OBftdgZvv+LwsVrevdmh2aX9W2WrDWN/cx2bXXq/v+jYtxnUB+xLjLiE+DcSxuhTWxmlSgT0biS3
g7lAUpFyqniEovsNyHeEhF5ZeAzkHG+ghM56OD3gSnCpN6ZZSMVxnekNdhlMJCoLp8HKGNmn02mo
tK2o5182hfu5jlw1xE0L6Vrz9T35bK3DgFC5w4PynsODhUdRsDSBop8k4bXPZqtILkRg5UjR2cuR
uhhdaRdpNDWZU+a8dKujVpgtQoVqeq0Myb4t929ZvKJRuWNumN4ID9VIKhTiBPD67Acgd9U9eKjz
vvjaaL5t4kDe3ws59ffZCjp333mwv/HuLgVH3/xjqhA0Zv3IDqbWG51biSFMBlJDP78PW/iTqfg4
DiM0TMSZtu2G08LeJGnBTsa6I3a4IqAhDHtpI6mX+H9B+v6YdbxiUqOX0I0G0QHIn5siAyhv+38H
miOLN2VK6oaiVRnKmkF5qgFy096JhszEbmsV2qLKvOU3dgQw+enjxI3XCIdUVF85E0Lj1fmIz42n
2qiMeV67B/4h0W+WlDa/qtbNF/S3k0sccjHnOzAFmrcGzRQ84yL1MmirKoJ4/3opzjnHPedJlJ17
8Ked15/FjpRv2iLe6PApJTNnUNsadjXfxlsQ1kIrj/QWdVnGMmR1Lu4fDQ1QwuyK34r+rwqseAB9
TaVGmojnltWtFRX/mZ6hCPwCqDuZBSljmXKOiMbAwf72dzHARum9h/HAZ/g3yQS0BtoIkb4jGlzK
u/KU/4JP87MewztP7TFqbIH8rYffSk6xZlwxxLHfa6+HZH68edgJwrt9ksKW6ldyO6LL5NzveN9R
+rhA45jciRXVDsSsmw+hhp9SWmph8tkzJPTIvwdwKaZQleec2slShor1w/U8dD4wZ1PS4adZ0ZWc
3tziBl1rmk+xAy3PYVGfTp0bIdvHd70jvJs0IP83Cx+NAR59cXtsJ/Qq5yUU0lZes0/7/Z8s9TsN
aOW0ccoLNESOyxwgXH7bflPK9ZVhRoX9E/pmvBAckOXwzjrZ8f4GbjNVCI84t1+sl+zfEunYihjw
JV/uJH8bYbO6Pv9c6Bj9OawctODgOPO0bCr835MdkAon7acNc3T9ewNLNesPlQpsnG5htrvyP2LS
ObcBVQX6EgcFd7KGRe844A48IUhFzAOsRvKgFMh87H6bLQ/vqfZ+oUmw0pOW4fAKBur6bAe4pvHh
kMiE3mN+Rqzv0MM5qvcLoBbefSYZDTX7U9oxaQNiRikKOiEJ+N89MUWybQrq8jT/WNCOfhBkbCUQ
7g/T5vZ+BG4I0T75+B5SGIY2SVLNXfX/meL6nd3Wh3lL66LHqFngE6pJLexzyce1iXh+HyNYyrYa
T+921tFOI/pYnMixxofPWK6gmx2VmOI9i3MpwuhvR7u0461DIf0qEMFVpYvu8kOXJWSH1TAz8yNc
biQdZsnuBbykBVG/CgveYirv0zffzU7QGi9cspLtydEieLz2MxkOBPUbG5TMp7m097Fe4KtfJcwd
gCTnZuaL0pchUtkXVVcGu3STLulKPh5RmFaSyOBdz7eripYSFEsKJhIVHdxv0NZfZ+x1YsWBQc3h
MNLk12qL6FFRdk5f01CVghzpJZXxlZl2tvf2j9e/3v4vUUESoWwIrFajzBLNmjsOamam57VTENqG
JqB0vALa2Lf73SJmHOlF/SXjaDJEebxACO7xGMNChlHMcT0nR0qDKITepv9+DoywU4OdiFUQ3yeu
rhFPmcxjyAWZL5WvmJGmExWJPhwxkanCeICmvmVv3CyUCdkmm3TvO9fY6KI6Dp0ciYBHbdhYHQZC
M2N3LMMEC2XzsN3XNEUr3mbQOm6LVt8MEbwNxpEBAd/c0Rh4Pg9u+mwu4QCguof+QS2hag9cG9Mq
gKkLmDu8usYkXkVV+mPMqgztrxVrV9C4Y/KraR0Jxi6CaM9zuz7bgoNaY/WrdXN8IklIXEfVosaJ
e39fGZUmMUk4rWTlmnMRnptaTMYQebQ6bIn7841cFA8+ysTmmXCHm4Hqv9N0TLko6lL0SU+Kh6BB
zOq4cbiVpgIWoBshJLF7TAjt3261veu4o6QbYuNkvNZsAqqFN1xlNGwCavOoEge+s7u52GGmtSOH
0MVQSeKXq/LvO0JydC5hu4XXmZdVAmgEkIuvyvRSc9lKaaCjM5Ycrfk/xI/YdvBuTrQBy5mNfoZQ
+VBo/XoGkmYqIuWI4+tO9j6gyxSMT9N15FX4ZOyneSdu6T+Q+CgBAyL/n8hQJx5jdDdJAzrHrLxm
dxtUkAMTjdJGl2NIHGNm6GcOJUfgqOYfH0zDADCG/TRir5+KMBri7bhV0Hz7UIdmON5nlxMyK5s0
Ru/qZCT3t5Ylu0tEReeKeOy2ccf+0DN3QOir5r8jNq5IVx1zGbaJUweZ6ZP5m1ZT7GqrBJWj9din
SmQr91N+WRNaBgQTPhyt9nNdv+6Yw28vH2jaBRGuKXakuLkQ/b4IkppNiK6i/7w/slO/4CPraHPS
oImI3dzhNIOwMZowELFhSmLVWwI8G82q4WmLRYbfcC9GcUGAJMnKGHyHXkV9kqrlqgTZwov30w3p
UvXWwQR9xLFUX/3Whik06gMw63W4aIT5cz6rP4WOlfD2XRXrf8j3fA2LsK0W3MWt3WMTG7lqdgVP
15Ya7xhr6OA744EMnx5ajyWbg3Me0AcvSEzeUDuq85Hcl0ZdHWyzfZSHM3joxcvQGfgHYNpp4R9Y
1dNa+8+eyjVYx1tJRZkGRsMHorrBIwDB0PEq2wzrRurQeDYuH35nsK+EHIv+9PsrF/7LZdKKSqUV
MSMBw3Uz7nDgqqIB72caFCVqoos58Lz4lCR6K+04lwfkMIGNRsiov9gss3bKR/fa9TK9OpU4aMAu
KtwKpHvk6/REnGir7s8WBvH5nsD8fqWJDtnK2woQWC8wj+Nkr9LEP94+NKz4GItn6DWSc9U+KquS
2ew/R8gvpBTg1fsozlFBvUoYB3f19BofF1xdedIyNrPjQh3RsJSouOK2krCzDdlXnJN18bBuqABP
VuHyje/37tyG8wBY7BPvmsqcZVT2c60KapAKW9vacmqmF7pVaZMdZCs4YgxfV6I6OEZtSrlL5KKj
9N1XB/6QGFZ4QxmRDMhKbRjEuaUar+nZgdckn+aVy5WdXTirFRrPIQcQPuncnmaLclrX8X/CJ/wP
Va1qdAi+YgWefaKcQ1feJlVIYF+OBWUF0PwmJj4vvsHLICv5P9UtC0x34oovPzydca6h+EDAAw7g
XcD0m7+z41R91KuzrzWE7Nb1xyhdiXKwvnR6aRiAV2X+q+KLuZTUv2dlq32A/5wwgCzxU0oqsv0B
YGTOUafH98oZAH/wFgAbdwB0Iv73uuLPLNnLkv7L5lYv3WteTcj6tMAepSO2wLBXCu7R5/XhyX0h
CG9GsRlN/Nv4QDEU9HMbFBu8VVZ0ZvyZz6BjwGaMjU2G2t9181LcZg4eLtRGCWtnv13hxLU56HYm
wfTiMBy+u8OrR5Vdx73svglZMdezNtLkTE54risLGjWSBZOQsa4ZyDRZdfhVeVWvLR5dNHkOhI/7
SWe0ewqRaaF5LxJ3guYtxfZ4dJv5WuhJ9fbIir5CJ2HZhWdqtLvY7Kz6gJmTabylL+U03kbVNK+j
ZAjWVQS1F2a98LcKa68BfL2zTqWsTdIgdUlIXH7DOVJ+3lvQC12CLxsL9x862EC8QOM1DouEGObK
e2qoHMtMnZHohvuf/8s3beO37R6EJwmSJYsyRs3vBSsUQeFLzRSUh+W5uBbhmfsggF2dNrMQMrj2
t0FwSqx8a+j+WnW5/d/8KQMfgWAJs0JfydJCf2dmXNnubM0EZ+KjMkfi163Tw6eKG+vrbKmO/bEb
DCShtubjSIKbTtNm0MlAhg609kxxZGuUdMP4ttH6oMrLNYQJoaikY5UyEgAn0ZGCXul/uy3CnF0O
FOmCH/1deWCNULXL+xBOTqxOInJmcFe5lNJlP20i/ujbKR/N+5GIsQLMNxXLl0Oa8zs5oof2cHC7
vgYl++9U/n6lVvX/yl0uK1oF7uVcv9oJMAxtQd8EutGVo4ouISGq3zD7UDWk2mOOKAiGdUepGlvj
Gr6F1sIgXv+QlG6HzBqRaTxCGcZQn2Ir7xCSX/grXo3kHfAb3ANrmOtNAB38BAW5UOBmeNRbXuV5
10+j2ZAXzUPuDEgZjaLAJsnQ6W3eMqUoO0ma7db5nohtttHGYVBvfvqaZYEc94sY6a/N7t7CbzwC
nx8k//ZNAF7S3d91H5aGVZhO+JHgCb7QMAP5AWbTq+wLwZ++QUL+BYiQ4wKcQUpuhO5GhdG7SVdj
SwtxgIrPCNB+oGpfMbPD70zewWVktsSdYJ560ePaV6PQS1E2PP8zDanvN42vAy0E4NK0cn5CHvbK
jv0ScOBRs4iasPQavjCXY24+LxwoVf1etrC5VeLhdNgvtk8H0PX7JDdoqlAG5h7uUHFI0R4nWdTw
D8qV1kIwfgFvEKSEsj5wHLLFcvFxK27eH5/1xk/fOXzXXpUirgNPMU+lEDVBAimSl1yGgQzLcbgd
APsD1C+qYdmRQP3yKOG247Ewc254jurijitRvS5R7cFGqLasukAj7PlkQUi8fN+Ydx5W8D+hKZpz
I6XpsQbO5/LvRTocqgTYghOFIN7fgw9wwifbtrQj+XSUBzzc4OSGquqYw0AlNVjgGKOjPThBt/wI
W/8/vdxSiUs1Nvk8FXVwFXl5T6299hOLEh6B0xA4tZavTdii7e+U4bD9gVXdESaro9A7AmfuK2hg
oHfKek+j/yJFEMXmiIqPe++XgtJB9v9LVvFupysDvF2FDHfzcHBFoWtaLyCLW9vFCE76Zu0Pofcb
w9NA2qjV5lK2IX5krUryjNV6nT99EH1m1XAGldRj/JnSqaYr91xeZ6uYkjlEPTAf5ehg76/3FifO
I8M1MPTJ8biDXrKSZOPO/yioeHdjqJdsRGhMiXJBdu5eExqtU1FZczP6186XHee0zqt0cgyfhefT
UbLNwBSup9nPvd2mtlUuBjPLWcFkvn+FABppOcQyaZoi9fmTuIm5ReF9j88QsLAOtx7/umcrThya
MmTq47GzN90b5NK6loOuHR69fpwJEkJ0oenY1MXFlpCh/jVNHZ1YZvykathafIl0Gd5sOTKFDyNZ
mCocTgaKPRuN3qUnfKy9Wr776W/uHE83xG3HuTct7F7ofo9oEpvRaBNiZlCTTKN1VDEtyIQXkUd1
xwnvXchOwDqI2XMX2a/CvZ/RiY9E5+q+wUsPkHerBD23L7Wuzr65BTstwLpd56YcgsZy9NqtjWUr
ABYixzzBzCDvziEly4ARpBmA4xl4p6B0SXHTiEcWtznZx3xSfkhWJ8wMwAFVLgHggAc+co71Bnb+
7/d1YVF+YYUcb2yvxQTvpDPJIxXJ8ULj59MYqCSy6E9hl2FkSZ4zI0rqIIrUmAEBC0AHiA0YPjUv
VKhPXm+sQ7vMMwPmPmo4ufqsyaGEVkB4mWMYY/TrC2qvxQN5E4+Mf0S23qp71tOPnHwDySciWGgh
OIfafNpsrjaGH+vRUxCxkJ2zw6eyQOZj3KnDIEVQRAun1KlYep4Ynjp5MF8VquveIK1LY2+nSc6j
y+lS9ZvnpHkGF+7I04Go+j4bOpdeEy+mYwvuWCW2zWixe7ypQ3BrvjKRUJw540aLDLSpjKaaVwik
6z/8aTbP7/q7z4bQu+RJ68wPJ8pK+Bx17wB2rRj3HKLVKoXC24EA9bpq7lR+tAft5so2duuhqOrD
H8B5ECM1NQAGmic4vlpo3JHjkPULcPJUbPBSZgmFH2SGBZm3SIYKEBckVzE9oIiH96BKZSTGKiu/
XYmT+aeUiwe1ETMg6+mwb6vWasaWmoA9eujEgchfDMT+mQMKbnYdE9f8rypDESZO2XFp7ZqjHO9l
P2gB/D4hzPY0MM43u2TjzKTbMX9WmTuqdQLq0a57ms8a4fHuXFykfXKcaROYFlrkKNYqZ6If0DzP
KtosFYE0crcWnwwz/huOyo70hK9ni7sdk+/2hZKWi80yO0MD2jtL85aasuoM85q6A6EpZNA0ssq7
ABtX/gAsCw/XnYp2j+uCCPJ3E2BW//meRc7hQtd3PY+ttN83+ezsBHYJhrBpAOl+4qUzFKRuCcmP
cXe9+GpMFJRVeABhCIzHU2FaWHrrfh/krBWdXkRTYkNlbz+r5DeFM5wUgLaP/eW/dKJ+2FVlFDtl
n+NTO9xpVnB0/XTDpupRALNzaDcu6o9hhDm6xhouS7xS/nnK1n6MOAR+ym6hEJmj8bPZ+4kONKNu
RqmORFItT/Qlpv6bNmYZw15wloUmGmxqdSVMbEjHZmmp/ST6SE0+U2Rg9LfcDUm6ZhpRyEXAswds
mPQKAkuLQnDkWTgKYRP5bYfaE+JX6a1WAfIg0nMcKEgf4g4wxDjVzqMG304hYxkZ4hYpUPEPrr6U
iuAvNcL9wlX93J0kGudCgsaYIZls08zIMT/Uh18/4eAPeW/sb+TYwwjPzjjf6MvqiPGVB+gH+BKb
p2aUQyizIh8hkyIiyRswH97dgzQm9M/uKH3KEpN2yh0SkVyeo11YpzrQpg3Qqy1fXnwqDBM7BOOn
Jjwcu1Pu8bzQAklUVTxJvRJyjOwzav6CVFe56Mxw9mxVlEVQdYMGqeNKDg7ZuA/SVZqq5DIYgPVK
VKqy+Og5FgJBx8hcT+rqx6U7pMzCWHlb3llu1VesQe7fobEGOfljELaA6KG5wCzwaNsMZMZdZWBW
sKuUnITI4Vt0TIV7/GCGIjRpMn6gnlJh7Seo5p6sQ12RUwriKBEFt2XgLhSjCOur/gpcxdqwE0sf
MkpLBELTag4SQEWGEtCD1tcH+wEUDuQxwyGot71BhcA3tZEkSssOy5qtitXQ8vTa+LjLyGLEvKKA
5eObL+yScLltCBni7+7myD1C0eLXf7Fp9ksqXVmlhTpD4MjBFNhmnTk79NQ7kvOPms7yDOa5msso
HjGZpkApHfOHJKsrP7ldvxoiht/qvxGuxBT/YGU0hq2ULx1v/pIY9TNUtTsvsagshOoB116RmWAq
FYQz5VVG/X3jcl+eb1CLdL5qHQuYWOqpPlGoov5israH8qGaYGuYAKIhhbkziNfbKitDGTbMdN/S
+GAxE5RT62tsrznpdSqbZW4ShQSs/kqcBpooHGt2ppUjpqkqRkhVqwIDEcKsLOrwA6eJ+nreE1ZQ
qC1ZryaWME9F5uW61aRQbTxhj4GjjhYrBNr1vpz6oi2WU/9cDzdS2iqyRTGxNcip2luOk+tEN89T
Hrjq4iokiZQf88COHXvJmn7JlY28txuTmgbTtKQrcD1Js0S0jY8MAk1htlJA/FhJQk3o4qgH4iDM
x8U35LPRdTkqrNIN/DZw3YjORmFLhL0ClqbxXy7FlGqz+Li403pn4MMXUCm/KXwE+mq9YjM+EEMm
Yz8KouY6CV5FJ9lNJdrVjUUnFQ8s53cBk+mu9gc5s5pdBprgCyLakwVeF4D6/E63sNqPi3kjdtGp
gwB1U3/dEE3nellwOCUhVb03zBddPqhfyTiqJUTFekeMdcWIkaOECSm2Y3uBnGd2IUIMUJCwfC1R
oy3Ar+kYJdJVps6xFSq+GLsAHZZju7DjPLxnQyDPfdhHTgOroqQ7KRNYlMTpLWLNjGrPZGMVYMxM
gTdNaH461NjYt5mOSW479p9MUr50WIuGuXzfgDmNIRobF3zUEXkqcA7tUxw3dU5HEdfU/Z4vG/H9
N7oCxpVQiOWeBH8u9vgPZN6ldEyYDYGecuW6CCU7LwafmEcJ50LpGMXgWpURIoyhS6Hm5pnMC1xq
Dnu9PMTCcnEHmbaWFtXo+hK/Cvv9h88xB9MgQTpPsGV1CURN7pS+m83tiXYtFB9maCi7El26uy4h
pjdeAtueRODte5ROyZyub3qrNdgZJdyUFoIHuQeJ6ppZFxxwqAr3Cf4QS/OyJVgOWlhf0sK310MI
hwUeMY86A6JGKVDVJLa09PUj4LkYA0Vqm9EFmyj/zD4yW389YciZsRK2p3KSLqi3fsUWVOL4WzSX
M6b1fWF64NlsMFIZEO861V5ruWgVog4WXhAnzFeABrOBaQ69Nq/v4pop9hpi2AVcaFNuXauGBo6l
6sAxIeGsU3rhgS8TUHH3j29+zIOiGV5yTSqrk1uwPvd+iz3YqN1YpaYvqWum0kNj2U28RguXQtEQ
+0nO6OjmLPHU8QLC75Xq602859Dbi5txhmR7yeHcRbcZX+lIn2at0zQfW1v4l7te8zkFJmVRoPG0
0/mjHKUjhTANfo3N38g7LAmsFdGVvRhfbF3m5cWZn3tHdNdr3byIxsSCEbXYdcUF+NbYuYW6IM0o
7pgyFlkWYdulKs/jh4ZQ+eH834pM80OEmuMwXl1VdUfb2UsBYUiFT06xnhtTA7XOV+SH8DmuKNLj
U8imDk0tKxYsFrzaXBydjHcb0+a9Z9f9C9PjdlLNuSopLmMce3SKN2D7GvZAt4E5xaVwmXxsBpgZ
O4UT1GJ6Vl0bqhu0keLz8R0BfjB6ROwqVAyghOl3O6Vcr4O8+6fopUATwC27WPl6YIqW0P5GMJhV
l6vcbaDgDJFtC4pb5RV67bghd9oBMOQo7TjmnH+me37NHH3IfugttfLFurOwQNuAJSK0QRhzezpY
8mqu136HQmcF6w5E8nssiQn9YlX0K8iRu1sMly1OnfJpgseTpOxfwb6MaNg0P/GItg8S+fxklrrg
wgxpgFWB/wpHEVJv+SCmdOT3iiDPfRcMoWhM20tcbeiA6M/4snx7GxmA8+NLqRNyjUIH2JLhSzZw
Wo9QV5fciaXAETaMlkekVmMG34FygQj7uhEZYSM4/rj5z4NyUfvcTTBn1ic3bDuRXS/dv+PPWO/t
9ccvunpk97J2gQPnlA7w6xdqsUSAsPTxltbLndsUHPYNaFaN4q7WdDY/LLFZP8cZ5Es42mPuMZmZ
AfajH6lSmTL4gq4SFLBqawueFICQHpIIbGP/QmDaaTyAduTSzoWwXYrhicJL2sECbqr/FbdJ3/wk
9qPTs6z1s/767elgzs8JrCb4JMXgDGRIY/aUgHXgi4sciIvjjImUM2BDbb9LcYQMrvcbgBiyNVYH
JQzRMu1kzsQhXNI3z3KzNcx8xtCwXHyekDQTDfmkl9HNPYnTLPiqvHpzuKBmiBY7p3MJGIKeq/Q/
iLUor1wENJVuB08n+TRgfN7irNW66hUSNdQdkiFPfPgqI5bF8pygXLiRwrqJskTbEfnvTUMA2RXK
HvFrywkTwVvCrrDeYLRMolZXft7Gg/F3mpmAuBky5yhRQGPHn+KVYr9FfCev05S6t1O3T2fHB2f2
34DZ+PYoWyMGVQPCK5jl4SkPiCXq6ns0iXOPMuspAqPaakY2BH8AkYchTlo+P9FPqMPKsBIpZK3M
F1QgXmznPUxPcCdUAxYV2AhiLzyDM/w/UUNNG4f7zvZfpOchaa0zKF6dAJLroq8lRPEmxCWeFVS5
tP4wBLX8HZ3hXqcB+YjIuHpgpiJhYFWtq6VTtlOmy7w8bMidpSs/3uuCSc8MYccxEz2kdpLpO1n6
VRpKp4TPBVnsFD/v4Wbsh3tqkXOBRQFPkYD7yhIAIa0pMR768HRlTJvx7KW11qJnVBV58Yjlf/ph
Irr1Zt4tP8wikJc4vq3jarD9EL58+Wn0Dm2brXgUYT2Sqsdu6J+yBWjB18snIN5Z8lC8SY8Ufw6k
o681/CH2X3IwCr/5O71smT9AlWVrB0mmNNUVj59a2DPok1Q+BivUZWDJjgt6y6mLkd4RN7FEqpYi
yBot/2xKq7spdCDjJTaXRz9rLspZkEDLZYDUQsfdXVJypZAwUbMHiPV/eiS8PujIAe6UOJQ29s8m
Bv2bVkGCznakaC7JZIu3g11A0W0NnjX1EFaaw/nMAxIN9ezajKlJGo1+vF+4x866fMpM3cEowGGb
BDi7Or7sukxCNv+BX8LOeZxIXT2PZaT1aoss5tVUGlTZUXdt6HVhADyVb6FnN2dvV/KhfYWc+HIY
5nJgrGR20kcX0Ex4Iy9OBihtMsaiivWShX9G76CSXJIyZE1ZnkyB71fw7Cs6cCXcrnEbg05sllL4
mVeGKgNyweyRvDyS6LOHsvHHZwX+MS6bl8fXNrLFJLNVvMlPCH+fSsY9OQg1SNyDuuLrFudLLEyi
kAsdd3lP+gRh0bGlwKWTsWwmMrae7Pko3sVj1mdFqLD1FKd5HDekRQtZY4n/5MhrMJjv+pq5qVGw
3+gJEKjHg4mJq+b9cDe94GQnPW6w4NACIEnl9P2x+a6lwLf5iouqPPNJ/yU4ByVKDfZCEtp8DYFW
cuEBcoe/Qw+22TiCHi5KUinww2qOg2HenyT+j9l/ZKXg7zH9P2UoR1NVdDk+bgebb9mXuwXJg6Dc
lVbUbLVflAMpgqhVZdYLhAiy/ZIzuOgEPj9vT/8hOU31RyjiGm6vL5dO3cgCfhfykTNdk8cpHqJT
lSv/NqmDlpiweRcqFWKrMdKehMTPsKw+GqLiYtnUxymucOhZ3jDg4sKa7etafVTrcdseEghl9waq
nf/K0eJJ6rq/GMXoqU09FDS69WwSR++9H2S6A2ZPEg7SCYnk2FU10zNLUuuS+xvVP5HW/noNwTnB
UI31ZU2Ma1O+CbSTiagyTsOZ16olXeLC5n67QnHf1KX+5dX+9u5HZUOCQ+UccOGoYVYeGT+3/Vpa
Yw9w029pssNHg52dQ9/nrBEnWwbpzLXm4ELu7VYtd9+cR5WZzOZGRNvdmrYj0GEmhN2Xqu/hFc/K
QPG8oheSioPOp9dBK1zBND6jY1C/jPzWNX+CgCxAZbNUQKdPNiujW1bRxwmUpn7+BUdgvHgS0QmB
/GlnF9HesPtRc1cdlkatildtTf6rqoi5ToHpUd/B1qiAEJtwupaBjS4CYZfU7rr7wIPDKdGT/zvr
0jn4XeXzrVY5lyLdhmIZmqsSRhcUqu1fHPBWds693aZS4ICr2YaDkodfK8bP02/DhqG6iXOh2s0s
8/Y7P1/A0yzCs3Ty76xZNcxZkimlYn+y0ayfqhgB+k3yvwvW84BKJleXPUuIIzovK/hV55uqASXe
KuV4mlZZ4eLmUwjTjPr2ruObepTYo78dSHHXC3u/4Atj+d1FktG627VWRqRPLUQzxck/i0VwqQou
Q++FWQ80IF6GMoZLmW1FakZMUWgidndMEyPWZYjoOF6qNZEnCagOuWAGDPrpMfMtvvKDkZQ4Tdbb
4+t6+U1/s+0Qwb9WZMlZXMXxK/T5l/LrGzwXPtzivfnsZo3LYComM/h/7RCj7lnGd7e93u++BxPK
L0m5wmJ5PjtjYpvjXrJGeej4VvBINlplmWB2nQd26qzI1NKQdwowIIm/WDfJ6aBFyBQQai+wt5GJ
+PsDsaZ3CRH2JFliysPWdzVqOXoJSr3k3oNbYru/45qx97bJ8oh/rrEUSK2VofPqQbnKviKZMYQj
1XljjrhQSmI+ZnW7QI6IrKMVkHyeULVoBbBZlZm0mebf+9FpJwBFZs5EPYCdPm2ZXBfogu3k8/vC
uFuzrG191OtG8ZViLUNEUI7gXEYpnzRHAxwvu3Pb2ZQ7CLrafaYq9JXnjNztR5nUKopJ75ykmZ/3
ymoWgz51uZDBqycKEjMCq4jxUmJ4UWhm2UalP9ATViGXG1XAu3M+PpIipxGBNAhlFzxKNXtaauCj
9EseYG5SpT7WRr7KXhY+WrpBGpB80xn3iADXADsvaXf/rVODIL1Ptg0UIJlDPbDSx18qFPRyiv0q
5uy8neGWfF6OgXy/2Iau65cvUgR+CERgvG9RW5VTLGaQxmD8+lTo04Nsxo8+8XwCBIhpPhDmmBJ5
DpKd9EjormXxlRPELRFAX6UvVrq/nxrpE8JxqfFMIHsqP5bg7WukBp/+cm/JjRh/Pi9mOCCLGE95
3oImUf0Q29IzmrC0tCRvSDqB8G6wCVn8NC+pA+u0s/6xPE7d7FdsboGKoXXrIyd3wSVaJZEScCmh
5VIIUxD1DIh4YRV7lIVMBUpukUWr8Lol59TuH6LxnSW068r2qxWSEl3F0z4MZcLJH0L6MBIXc+dy
zY2r1o3OSn0vPa9yG67VijnMjNsebXbhHO44YzKWMH0rFywsUmBPjT1/sUvpdCBtC5rXkJD7FGOA
CpRdL3vVUjQVaV5FxI7Ewc4dtIkpGfc99cXeXhBTYJOfP9snHXk5lTm8VBodV49y32j6YLC//wXQ
3uN7IIAVx3Z19DDeCpPJCeTgRW/8KS6sNWh+vVgeKe/cGXl28bvLURb6o2NO9+W7iJdD0FER27hO
BsSd7jAA7fgjwxW+y5WaWd8ZFz5UmUvfsbKgqlYBh/p7wFdgNlvi/LiMpE4Aykatf0o34E9Bk84e
IBYZMTM7Rd6rFWhmrcBSWIvflf2IjaE22RVibMkZRZ+Mxn8Hj3dS7IkSdIjS+W5kjPpIRy1x4X/n
PZ4KTLmtLms4Zb/lWeX+CXilx5JlJBEbgNwwez9+Q9QBRr91LGnEI2xWXzdNA2ifIKqNpVH8bTzL
h/PthHKn6RmFukFsl6BXJGFtjwWJLZeJiGmMxMqLDSQTnp8tAH45SUqayCnxVtxaw7AyyiPKRjei
vA437UVAoDvooYK2KrcdcpUIVcBferLWyaXt5tLhKlRQsZQk3V52VvEoPKhGXMjSOaiw7xZVla78
IQ6CyIQxA3D+Qf4xnO1X74UUTSGiFJWvA76eDFfl7SWMla7LZqMVARzYQzPo/LHueXTQOB1Wht08
ribXb6OcIn9moFrRp8ZX7bDDvH3n9ZD/SelDvMvKEIJsYPGG5X6muOozMm6bw56JVFbP2N+TGf+f
mgD55ssz2YoMxvcLqZqVsJBBaYUa80sdrg3EMtQahGV1FaDsxO+JGv9ZrNgjI1o+t8Onb8qbEq5r
ymCgsFUsQ4SFOqYSJdF9uH+ccTMtZmKQASGRnD8mfpxMoIXH7Gh4V3HogxLkm/TiEXa2mBpy94i5
0jSysycdQw2OFGMk11FT3EFWB1FxswTb6YfuWzA1jkJPMdXjMnF65slAt869IC6F0/KSstp/1SYK
eZhBAKU5Mda4GsAVZi0ESZZqG6vYa31QYtU7gFzmbdJm93+B/3znOjd+uAX9kAfprAOm9cWg76xg
PG0B5Sr8spoYF45SilLQmz/cRDDR12toqgLblLIxVjXCWjf51B+1SmZhjQyNx9FmbTaKf3VAsIJd
a7Cth/RakhidwYbK5bKJ7XQv/lNEQHScYVpLVmnktSvFxIftEdvchDRR3pWSBtzXjbl+lY8Dbl57
uifQK8Q1PJ1jpcIlEqJ2zU8LUCd7Da3fyEL4sqtShn/YFRyGrJz+TuYoOMVCXvg4yT0c8eLCq9ht
Sjlp+Vn8L5lxiMpCFyzz7vGrygEuAtsNwEFBoidNJu/GPIlCHjGx8mSRBBK7h/l2E0Ubxqi/Og1M
2YczcSfVuM8NdvzLYxrzWZe0q+GHraKK+MX7IvuNREGHQ5d1i1p2+MMlZ7ns5nNkDIrjeY60RWO0
G5XO237pPpfmXVGLXcEsdeOyoz3dWCcgtrXi6MHQgVuG63Vux+/TXp6w2zyj+L5z/oWfABnOtO2b
jlPxIL1uU0a4NqMSvYM1erkt1G+sPztsf8mp/5Ru29jSEOon8gvJDUmSoj3Q61Rb1NfaFbXxojPH
JGOC54Ycl4mFprCxjZRuQGrYjtzWWH/wLC77P3sdgC0E46L2NtMBKYPN2isJ76UqW5fxjOOp6CEc
/lA+vurD9+9Nyko6E/0DJrLavjmLmfRZGqd+H88tG4EUEZF7J5mofTU6Na3h7sY18lSFbFllVol+
ZGEbPO8oodRpFZgU7e9PYNHYuC/CpKCQGoISeQC1cd/2He+StxNpbGgCb4bjGT4kA1WZHeu//ppa
S2VpYuIoFY013dlcfOqF8Npg8C7PSXgUBkLQrzfzi8KaooOIh5ORLBIrvIbg5C32cwWimeAR1ihw
mZEbzbnhl7JRlwGxqroeIFBGOIc4gk8GfBrkV1aZ8MTMFPRM+Ci3IuUrA+6vLetR7ZBT+XWQ03rt
UpQXP63HBpn8fgcRhQcpKsNGl4RiJ1sirKCEfc3Is4PFAhFS7OfPdUQEoD9jAl7wecmnJqIXyB75
ddXVs0+Uv4YjhohKVw7KeZFEk4J/HRhQ65u0ouqHPcJ7esbQwfb6sJ47dYkzOCLcFlLQqQvlXcfp
CyDl2ABZ0j/F3yIlabXQeVl7aupqrTShTF3o/RJlT3losvkKzQeFSSm/sy/u8DzjDAhLRMdiaGpe
rKWxjFTQjB3K0VujITV1idpc9J5qkaZCWgEdZAoobtxQS/MktXC7x5fZCRYl5cnNwQRF+TTXyFzQ
dx7HMcbaqiclqLyq+VQrwlSh6Lup/iwu2wEWoPXMcnJDPzuURCWPSjZva/kdQMnDE7xO2Wg+7Dq3
znzseg17i33m4AzwJeqQVWaXCNQZ913sDOjRK093NLt9c1IuOvSG1qis5CfODh95xO2C95F5VJn2
HanLlrWoRNJMzZs5Gxmj2ahCqE5wRAV/uyNZfyOqvv0tiR25nlCscv+gYbingLh2YKuM18eK3LKi
13Micx9OJiTa3gwjTW63ix84zHjhUJv0JFoikqssmgeVkMFu/97CFSHiVbW4dIF1wuxst13ZTPjA
l9Y8TzkIPP0Gi5PyVlY92xB0Vr4h8P+TtQ6JGHjbfcTd3rPrDeXU4v2BRekdovVpDlfoz+V3BoDV
7BcjjIVIndvZUggyT4tUN0nIuYtnKnnp/4QOiw+I93H61rOwCOvc1PcFC3zFGN13WAYvo9A3EgHC
xio7MVPMxqGZnYXrN2oEbixU53MBkc/PREm4wPMdzkwEXL39JSQskbvGGkjRFfaF6GY2jX6Tvw5w
j19syqDJjbDPupwKZ8NEQjMHrs9s6pWqFBCVX0h1p5KGVicPJBFvG/rcKC3kWQTMERGRMAYvBhrC
dA1NNUUUPPGKzqIOz2b6RXStwzn35iDvEmX47hAH9QAQ22cdn0EWRPvI0IBnUB1esiemUwSc8rIz
Dd7j7hNf+e8eXkiAmY0QHd9Pxj/pVEdyX/XY/uyws5tTtPUpfdfBRey44k3GhKWXd27k99qaC64F
xDpsUbiDwh26r6VE/a5yZ3JyIFQYLMcmEdai5O+zlEy//RFgopoJ39nSScZB0MKFVcYSYINSLqZs
ahcHXpHcvzNARwhNQWztnGdcvW4swjyOWBVz/+oG284oVvuRPSOUFd6IN12hptTUwwmtgGAj11+a
8JEh7y66ftgQTRNAKDSdffqkMIJ2vaR9bliVO1y9KwrmTl51M3MM4Xp/qP/mVpcrM/TPJ/OcKJGU
RJoIjghcOG4YZf0rDFtMsNo/BTNYpdkCoNgIYb4hOFxGkjAHZreJxwTXAVaKR+L91uFvdeFjMb2B
ECSBXMJEuPf1Tge6hQxKSnCtXi2EWWmlCIn8Xw/iec4ecTklhEr9fmDjd69r4+pvmwzvTg3pLb6j
HnIsQ39aqM2MiLh4p6MftfK8GDPiaZ9/rIdLiHNvWmcHutqB+uKFWQjZTvoyiFnkR6UYNa4j3aAh
8U5ZCWljfBQ+zBOcvRsHOOgLQWqIqGbq0ce/el492uUn3IOYuWeACybMtGxGG3YxcEo7k0Z2P81t
lHs//7AtEYJ6cCIbkDA2OJAY0Icoawm2O6lRkFi8onb6L/Pmy1WAAG7MYtKQ8O+FvLS0g60S9LR7
Tcp8oa/Kz5nP89KHL0pb1p8aBCQ5VSQIL+3+Shm7Q6jYTbeiCjg+mDeEIVvazBZbJ/n1gE1cMK03
nMMzICoef+LR5fZ1OEcMHffvpZkNQrayNrTTDZkaWVucRaTeCGHGUHVIP2YsTK754reshhQKpsU2
dg4or69EFOESnVL7rAaI/Hl3WJ2vXzvq6+AOt77bJgn44xa1BFvEAnmgSzZPUOT+43IRVhH9twxf
245xisB76GLa66R7UYU5UFLoVhypS0PRn2QQdO9d3yRq+LCSfkUFROWFNCertJYbKHGUm+yh2tGo
ruY9hAsT5jFsmCC5wOof7tVsYYXYSZHvDwYuAOR/vM9OGK0t3wJ1Bv50eI8+rtA3Dx2eiW6gtrIF
xPA/GyEZJp6H1wjFnPFPeTCN3UB1S186sfE6Zvt3/KLKhNxxVnzz3NAuV69ATWv7PvsEvtpDMVCZ
8upQoBr4Lps8M5OgqeQmb5DpWMxQhZn4K7GsMac5sFMaD1mAWtDO+UHrZNqYb9/BRkrC9ld68p7D
PnlFx2wmaeOaGBKQAIwTeRXo1ED8eSzdT/j0ixEh7DobbFw/Xf5qGYuw0MI00hvMDu3QwQHerCLW
f14LkiuWiPbLpWQan7xR+Sfho0/lNFk5dNZk+0XMFN7U840wqRWrdmmymxhj4zPVm3mXyubxLr17
P6T6yw8Hj/FT+GWJ7Z4UuNfkZceUlZJePhlcCaPfjh0o
`protect end_protected

