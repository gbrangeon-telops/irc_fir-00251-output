

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mCyyeqqjg5/0TkdJEsEEwiyDfrhah9gG0fpTMwUWGOKZ3he/dpUva8HsS4xtl5XP9zdNgeOXA7QE
z8wIFX99RA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X35C+3C9De7vC0qODnacg9gsvk+3IzrNpqQYzh787Czr0LrIg4SN4n42C6CPfkCBLDXSXwC/eOXr
yWqN/Hj/SYBmrS5kjeF37AKShalo68kYRaZgUNEiNvBgjtaJt6WRpWYojbh+ogFdK3xIXCNq+Qxl
K0+QDwwSCDU/YMofxGE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n73jcH3HYbuczKsWgG6ox7VZK1YnHzJQ1B4KxEg4B/kZylbLOe/lb0i8/kn+CjmMlUuMK0WQWfed
hITAZaScEDQ3B6jcHH/bNliHMpa5PCxNetq1i73KuqIUSMzdaxGWTSuFoXR94e0GNel9SANUqOYF
vTOS9qeLaefJfWuMi23yYpmliTIg3f3fAbSdeAfef4vuNm+0XcFw60RpJQs3nrsFq9KW/GfqXw4u
TZNQUQbt6cL25X91FZ9ygQq3zmgha+CzhVMH2888hx1Tg3YKoHcpCHNpnuDfIIlbv8c/WTDMb67v
IK74ph/GlcH+s638TtetKCgz1jniP6o8owuM0w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lgEz+Sb20/Syw0As3tLsdRmvucviIYGeDJylwgde+NWKzNiVP+by1Maor4kKAxxHjnI5lkH0wLYs
PhqSC4UmzjejXWlU17tjRxtRz6BbrpAi6gmDH8SRbE1L1vIa3LM6opScw2kIKRT06DZ3npJLvb1L
GQYpSvbMBpeOoeXBKyg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cuBsFlva1Z5u1UA+GZT5hw/3RJ+t4o7i70J4gtLUlv3Ik7QI7QGdbqQ4mg46AQCjs/XyJI5tDPDQ
SIWqonbFU6W95Sa+82Fm2FOLny1XsFw2bfUdFeJCVtBal0R28pkG/kXPwJRvcecEIrS2a1k5PBE5
sZrJ66qcp7DI4wbfzpv3ic5F22QlsAxZqXZEB6lBkhSRHmx8sxDYGL3gz3qyqFuTzoFlxGj0D2l1
7IJKcs+gQikUKNCj4QKZQHmP0x55BD7tR2tDFNHuJwLQeErQDiAmIcwGhliqTf1RxwWpWFh5JUyZ
nisNHaWXl8SFhFbWbHjUNb33VdqRqkyTz+gZkw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49408)
`protect data_block
HDBfIqsMKfNDtsfduPd/Ofw5SEUd8gfztnwYojBqcF7m2lmhoPCIivzLcdAPb6CwILMQZBYiQPDr
iwuB9LtWhZCKCxNGb36OflFOt1BxczLfGlfFj27F3w9GuLIfwpzwY2w81jZ67Pitgkh7NDFA3Oat
pZFedpxT/XXOFvWiohv2VrGymFih5buMt3Tu2meEK4+JOQSZLAYH/3p2YYdrhqB4dh4PNzwWJ+41
SFEgiK+F19fOU32V5RhDIlaimdDcuKETdtKdfc45k6FiC0Waz97A1Z0aD67tSfE7Z5445riylsAG
Dee4PJby/keYqN9VG2KGG9UPOJjvggn+K44YE1ryKqXuT+BL8BSr5y4rDdBhv8wkzlEOD6YWf3Xq
7QLsVuVeMr14WIGi/sHaui4Ws60EG45BMuiS3XwyE2gqa1tHTDVnxlfM3mkkriIzUVWAzg8ZeilF
HoYTtBsgUI1lDTpqxUfM9S3cxF74esTNR01Jm2OVqmyt5hVIb0MweGbt87FrGSZzhwtM8lI4chDk
lRJCS7EiX/cxnUgJds0s4YssdakmjDwfgTjmaiak+AbAp8OLaGb02k7KjJaNyT6nxugz5JWSUukU
wDrvMHoYQ+vuGh465Z/V6xnbdf3RFVfPlJJdipYvzQx/ZkEqPES34P6TTpTpJWSVAP91vJV2ik+A
zV6mpcp1Rm50z0zCzq7Yhc5ztZo5yHkL5phRSAJJURdXyxtpMEVKx2QDFWzBdzNEfDhJKc4qRGEk
OsJvSXRxKsNJK4JsHLbIOohFXcJlLfoE1mRjYStOOStjS5Nvyvqn5pQvf+NHjd+ffUN1BMB58H1d
iXwzNjTRwHgMOxcIBXAj2HBptvcKg6z2yxMt9a9UxE4qXyelbKgI0c1yBQgORt9mVU3QF9BqK4Jm
a1bL5cFtIoqD3dofSWVCDKfIFc2Q2ccn/ukeobFb/+ifgNwjdj6TVGTz5rU0jG9IN52TPFLnvovg
QaeOih9SmsDyy2id/btMIkjtEUszeKO1QSdpW6pHqVpV8ul3v7gH+j1OUcQmJ5mOTLskm9mzcyEh
NM7XHn07v4TtDc6vXFAXI8dOOGZJVC0g5aGxdtymT6F626+wrw8o/kdHy6hCTjwoC0As7nHO3x+Y
IEcUeXLAj06d3i+ADEFV8LTrVtmh+MvBXoXcggbbT2FGZn0n62X+DmmLos3QcqDpfcWB0qSBLVRE
QUkJqnOVgIFd/suZBcMnsPpdW6tn7nf1dknGK/fkqobgsGhEg3e1H2SQtaR7lSM1dRW0qTMANDYU
+8UkxwI2Q+74tCk3Ra60CAy9oLxFHiMnyUVokdsGkmyzA4oeeimB2RYSArF5ugE7MstvmzImJfFm
zCvR1OJQx8bfuu3q8O5fJ12pSb+L25FrCHLil2lSAo19DUEVFv1PHX/gFKCz2wFkQIjo6FuMkkA0
HaWF6bYYKIZco5jVNHbwO0/gBi7kGt8vpVtZziq9iAZmvhfxJNWxjTKmRXhzVFAREJgBtMGYEKcs
TmhYkHBgbGFHDUrUWcEMeh7/JB9n1U0nn821gXEjTP4q+3VBtiMUGfZKFrcsQQzGu/Kn2icfyI0G
HjDYlnhu3vr0M50Ajt8pHHPvKE+yYnQ9ZwM1N/TEK7bVWwKnGIRrLdmb1/qgx+3esaxVN3Lu5f6K
qn5Y6svArVNZY060XdAgeRlJ+COnr5o6/16ptp7zw/u3tqbJBacmrTvdY1NRh3uHhJImsJziYsok
fPgmdoWaszt+Kwo55/PQ37sW7wMbCGMVwbSHp+DBjDHUmACeTbuZs48tut0II4n9wwN9AyrwA03m
zOvrUEx+ojr7JouvNso2HwkcXycjy+LQ/pS4YQ165fhHNG5gJWjeJXqytcVgYMksHkm+kydRGKjn
1TK72OdN4iWUQ04ghwj8JAnDJ553NGV/3OwSj8zTf7RMyMF15z7nbWChv56JuSv2y3+tF0eMKm3/
U5ZNofxb2AwI0xxIPSlKK8aMGUaqFb0VFvV6EZKycRUMD6hli/o859Ws5POdf61Q7T9VCHt4Qg9c
okvGt8eOQsBBoEiGc46JtdMyBiJOvSHXsDSTBDhASUWPc66svQ7vEWkC3PMjdg669OnM5mMR8AeT
DfFIDMiUc0vn5oybpF4Iwn4clExOnaGbFeRU1nfQW3S+BgcW3VpkjLeGzFn/aFxBLwUuRoWyfTIZ
vJ5A5nrEnMrZ1REfHKCbvH4iakirwEL8oTgnMeImw/lXafNy4gh2/3UQ47Z27N5+FocoyCltdq/c
tRbf7Wz7qJP3Ath5J0rgsGBjdsm3iXzJNARfx4ByINGY43JxMvvdDNvj+Z4OdgVenDTMoo4zWOwG
InSGSmrV4XsRYLdE8YCqJkrSygfz00M9C3yoXJGJZeRUCAVx7Ccywl/6/NikIRcACeH6VFbxP381
cLMzPJ1xBALPaXbJgS+eKR8YD5gV0pD+lq2WDxbdKlRQnPrEok6AiLZ81zGNYN/1jK/YEcqE23jw
Sqh++VRUamdSCwVR8ZfJ5LRJGGwulZBJ2fnieaMQOBFK3Cp2Iuu7630hPOKYEv1JJMaw5QEMiJiA
JMSYdgygTq4+7rOU8+HLN1VXA1FVooaPnkV72BCnv0IP6K77qsF+Sw44z07IyS+B1xws+q2dNJGC
hbki7v2XU/dC5FyIkKdtaEqT2CZmFgOIMils+re75Tw2WUsvDXNajl+pD8FkyWI349qryxp6X4If
gJHD15BNNb4tKVQym3VScy68BIaFLu5q5ELxOSRKG4wGtrBorXDeiO63vur0yB0nXKbgzi4u3/yj
TSFQOW08JhXJ79bMuP4Vb4kUxJpFmeOL/LApA4J6wjmgUy0thFPSEDXXYLowYP4IY5KqilGGnebU
BjdSVHd1LQXF7wzbXVRa8zA4X159H7j16+XCA6EnMX9Ysn5zh3aNYDYS3TK/U4dM6SXKNKgT2ynW
wOrtU/JPEuTC+qHu99/SpLKnsir0/WR/Yht2yLbajCoIw2fBcxSrfkscN79wnFyPE3zn7mz3H1Td
fiQRM+I3GeIxxwfDkqN0vep3SM1LSfU8DmirSRw1USMCyv1t1ce1/H42+rh6W6Etw681XND3PW7S
cHQeopQNafQS6sMa9TZ3Fu0RBcE/vXmN46s+9oMvLSOoeQYSn34Z/bkm2nUXuxVKWBcBMQl1O8By
+QYsYMWKEfrzM7M1eUU3l00a0csXXUuGJ9/ntGcPbSMusq/Knf57fBmQ8wdaOHS8t/3QXB8Ai6Db
jgvu0sMx1ueo/IF5g9lfuhZVIOyeW+87DFFQmcVLz+NpDEqOtOai7B19cWcB89VM5nbro03aSxIa
toNa3RqmIuFXN67boYP9lnZ83OgLqiAM0J1Rp+AxkSJU8bxBc1PqxPuYWn/w45sX4KRyk3j37dAF
drYV3tD2aS/5JfuHmDLwvuMykWI6a2U2uKhEsCRlrmgMdvTmglVfkbDhF0qmRQwjiCCzDGl8p4er
JC1VoGvy6miqTqvqtOJafNmO7JIxVtNDPs4HFKPrMH/eHoQ/10Ww2pxJzgH/FzRX3/Rp3YGhry6s
GHIBFsfKegEVBRw83PQDI6aOUkPfFXxvmufQSDXbf4UtmA3qtKiPclR3Sd+cnq8u3cWGrW/wwnzP
InvOUApOjqM0E3juFmGTL0ZvenmE0pQrlp3SxAaRM5SJao9vnFLYAj0A7SpUO214mEsufy1HHeru
PILZ7ryLFg0jzFq8GvOOKSTxHwAJTNGZ5A81q4qIZxSznHnUZRuGivojAurMsjj6n3YGOgFODCAh
t2pLLUbam0c/TIv+b91ebUnF0xlc316jswImAhwFjj9ZvB+wJ/YCrxfFCqeCs3khnrkWnOS4BEyA
jhvjVHSkO2E68xzIDbq3IWAeMCECpOYt9E2ix+2GAemkIxCjwPvVgmHVhOluJOJFpjt2U1Z++Y8X
QYaIuI+KZWuQBfrwO8r9mRDMSHznaN/QA7kk+i2elg7qwpn+AwVIWDNvTrkPciMa8ErBCjKxqdsl
Cqos/Ysa7Rapzewv7TPMujPkGQtfAGRc/jXZngnSsAirM+h9eq73sSaJKtMXtKO99RTEtOm1eh3V
AdnwzeXWk7HqLl6y3ZZZdZcbDNcptFFaPoK8IJsM97ZjgTH8b9XwcVfBqhdH7bDGGVqLyuZwwEqL
vvtc6ks5X4FxXew04ut1kiRe35jcIMWsqTZChXyl5QuDHxAZPe3BX/eQYABDZtyKK8GAh1nsjLvC
l5ycHKk8/IMIZDdckVV/1B7jo1tNk+ci6JlSPqZCZUEW0wbiWdE6bMNtxfitveM0XwPATUUsiCHe
TDo0PhwaoFbdY/dQ9pwSsbpmEEjN/JOg6IXdkb/QuM4xNlQ6DJM1KDBm4dkDMdTWwn8nJ4CRnojy
drRkb51jVSQO/drExYrIjmlV4DXd2vmhjxrYFaokF/loCky5nvhgEj2TH15n07ReQ41IezJ/HMe9
dTJ7QRmVrwL5OvGYkwCN543ElEIrGSh3inor4rGuEFh+rgHNJlNMYUVkWAtNInsL0hABRVDJ4XMe
YekxTsbBoMp52174+Q7gpZ+Hdoj87EHGs/SaasHNOepWzF/PNc9dLsZ2eH/OucHknjSHnePMD+YQ
MJHHDJ6YQkp5Bxba72ldGwcB11cWyq9PUGPidGvTAg4TMsgY2rqM1ADayJ9myBKAPaFq/f/Q7+mB
VEr8jJH79zm0/EJfp2MuxUQheWIey2zxJHUc3Mk+hATBR3sfua9eXSA6D/HvtFdDdcantUcZlWMZ
ilLapwpktTbkFQeeoA8c+fnvjK6F/x8yvuOB8O5qc1euYrvZ5Og4eme/z9IIkvwrqgVOl9MTIVfz
PrxSxWfCgzI5PF/frD89wIm96UpN6vw5PkEg4jQWPjimR+vid9wnAuwnKNLdeL1GehurB6PNbucr
vyl/YNF2XhHgtfYF/cxoumc88iayq9O0RTa3zfNdPuXwJ7Y9Bm9CotmI9SO5WfLZIHZ7LfqynSPj
Mx4kRngUswRWkoCDxJa1fdP2jSF8VhGE3lYkk0pCQ6ikPACYoeA5KLEZUQshLJ9NCWhTVmKIjEG7
p8PRpDYX5u+svmDGqkrsLTaEqWDXzTXG/BPcOjHQn/43i12/XKHWkHfWl7gfk+TNqTbuyrkJoatY
C8k0Zzq8v6rSWGj36PIlZJofrP7cuDovA8OHK4lY5USEh8X6bn2Fy8OaOWh377aBOrQxTQcorLEM
dfUW7zELN59PPGHCV4lP2AaDGnxKfh1OoYUthroj7whK/LyRVJtfZHecPVdvRdmYS465YqiHnZxM
5TSu+Zk1ZtzBe8+pXBp9gmImpKLNjGy8nI6b321LZisMrU2pez3vozPYNPRjuDJLkKpwxRLtNjHQ
+xSxIL+x/vBQz/yRtTQJlUgzEzapeYb05N3MmbcvB3XWqk1qnSuwlPEGgyv693Xt/8iuVAz9nHE7
4xzpsgJCpqGGP+BY7CbqkiEK1GfNcinjIISTTSa4g8/dY3wr92xP7c46nSudwpFrLxQNiEUyaHU6
h4S83/Oc7SaI7xKzT6t8Gq5n6/oI8G0dhi1vD1D7YlAHqpjkMpIgYst9QpiQ2Jg480cKMKjTIInd
vij+ANxCt6g8PGazFxBL7auE4mMKeawWp1hStfm6aAgvYr4f09zw4UZ9OCFzseK6D6FuId4Vr+UL
uO2bbYH8yb9pxcmrS18wEbO15VLpcGLs/j4bvTckd4XsPi3QOc9hhuKzkQ3r2kKw/GReyki70Ia5
UIHQcloOfj6Ce10hm06a7MsZygFJI2k8z6O+kNcwQXmR6cCA+PyFw+9ZPFQXRLjtCdjZdTyos495
90ZS4qaZPjwgB4myWbAVLKGfTJioCCGKA4iUkx59lVn1BiDAUVFNeY6yzZsqhPB522F5iRN2oV/L
zfopuf5l460Ic7UtC9PHh1RjLLnTa4PodhSijOZjKyR6dOlzQ5nho9i1RvaUBlsPhqauFbtAaE7N
mABY+wqZ9JjohJvBgvV+huBDtrix6d+azAno1q2HU7vZzpzN4x6RFW9Qfl33WZ8PuUG2zqfg4/lv
SGsHf/TL5vbk8ulmF7WnLGedkn7nCznVoexNZAJu2jzz1X9eVqs0g39XIO2vDNI0K48VwVhDERNi
DTv1uG7V5WJSioh3KrqV2fDf07zNi0f6dhjxsIHrlCbxuimU1iupXeiooVExctGXZ8aqastcqjjM
52RM6LCqchjO4ajl3hCw9NgG14TXl2S4Ze+LWCq71gZXZHkD2e7G7L4BAJrw5RQBofYUdFTVjpxk
YZyYwABqzVpIrSGI4xCWuEmV+Wyvl6eTgtJgGhGC6T/JAxVJZWlSHzO7+SERetqtac05JtZtcj1i
fVlAEhAAgJT1uTN0R6OJTs6CsFEwcBGBMWfh2czwHHQ5apgCwlMc5IqYnZHhbg94fZ6Ap1pdxfAM
sxZCzD2JEbrTk3suzYP0CaH7R3oEbyTsmp7g74WlVF2mCVIFFn8oAu1YOUeFln+QeKW79A3yyvfb
HnBrPuvDL1V6A1Z/PCbzjh8P/WCAqnGbyVOHZN5Yom0NlAm7jCFcv0fbc/pWyOlSApBkyMqxdcjw
aekoxsTt9NxmZGx/CVnlMnpp1bE+TbuRfhjE2THrlQ9r1KTRmG3aJgu6yI31wCqogdAV1ykoBfAC
qqtWqzS5fQgXAKOczmxNyHiO8ostgdemU2CCeF2XhVvTm3DN49DH3r/4SkvU465v/q/RDzVrdMIH
yZJDj9tDEBEP+WuAOPk1Ism3CUDpMD+DaAzjq+qJ0FewxcfAfZIVZc1+EQOQbzNvc5Hl+WomkWTA
nOB8BbPn/+sqvA3kV86AGxmSclN5wMF8V8PzFzI4xxBryDMdMq4UM/1TGRO/6zK5DXfXJIO9+a//
aLvU6AghQFR2k/a7kb92NWDnqsFjQ2rc2zBlIvSCr7gYXk23zQWrakn6G6EwLVyJF1y0yxmPfgtQ
mb/5+/aCEdvnA4Gd1jv+pgrG+oZGgyUCpVG6emsp1C1iTt80yjaLvxFWfk+vy4j1H7XzSvugAr65
dhn9fD6nlb68syiXftru+yDZhoLOAnpWKftzS5moc7ZAJ+LTmrdS4VdzXV9eKqaLKAUe0XbQ/7Yw
XYy1XYR7JhC+7KQdJNM1LpZDDmTsiFPfwI38xb5wBG08Rhm8ofcYr9N8RI4BEoK0AmMZa7xD1NWF
BJQefK0DfRUhZTbidLb/PS9wtNxxcydkpI3CU1HSdVcxj9b1T9JvJ2vmPyWgi4Q9pUks1n2OMxC6
Te8c79QfPYZ4E8vhk3aWIBJQ9uTnSI+H+yGXWW3oAWYsCCFJgc7iXgyD6EYMvPpo1N4lVBEK6pGT
U5qxbhSD05lofYESccqn5WBXr26lgFNoY7pIC3PO3ZYLgBACTRqPaN+qgIEMj13G+G0SGBMc3pv6
dnnpwKH5yqw+eW83t0s53aQA7WDH0pEAaDqBPlYOBnlrFljtzoV+TOu+zbRF/lvYXT7wkp9btocj
ASUwzjzVujIjLRa8X/nZJjiFo/BbxsVOc3Tog/XWJkW5ydQN+ULPFJDPLqzYuVqnu//AZVxpZUB5
6v2K/s86g16ELwTSG2LW9oRAMqRzzXKey+SEZUBcdQTkvPjGRwvdH9iOVqRWYZY/KqpuDtPFPbyE
ySofu9kl8Bnr0rV5L83noZLSOXodYk/IEJvTIXmVoil4btkPmHQ/1bqV9xx9zkC4tNiyxngO+xtN
3cDdvwPcRnQs8Gqp8nyJBK+9FM80zs8R9qYpUKS4/zvJ8aBR+7cXGYX9x831zIKYVgLTMYcWsiuI
dehtGr+k1O8uZsOsfSdVb6GiP05hUApvjxd8BimvXA3qoOmEGi+87oVjL+bSBrA0gl/4PEdBB4qO
ht0lUThn9rS9eELYVsssqyS237jPG7riWBj71Uz0zzbbIKL8d3h19lNA6f/aESpQAU1qmqfIkWTA
raEQ1cY1ddoMEa4qDGVnFuZWckfetG2ZRr9T8wfqjgJBbIdUwg2HA1wKS+G6OPp6YdqC1/v3kDNB
EbGgqXAy6yaTx8C9pNrb7JCjyP6NwhZeRCyv4WtM5IEAM0P8QTv5Dv6Hv5jRn0MnDMdIaRYNihmV
iF6ZtCfctv79SZzKaW4+tRrKNk1sfAEMWWeLUHAlmzbihQbTy6OrTlZd5tzwwCqgx+IHNtfysbyc
IPuXARGY33P9pwR6qQ/VE7B9YmSwNdpTXQsA8jZd68APCfEedxfd6fMr/wMmw2R4NMxmH94o2KSw
RcTbxBosj2v0MMAJt+U9v1MA7r5ZT9AKzsyRDLTXFge7FmYZH0OmBgyWA5NrIvwC5wUmwy8jOoVI
0Cw2qyrvmGbqTT91VDz0rV23sTtz6iZOO2oq8SA21X2+PueeTsDiwzwMwzE99Z32bRhL0QUdR3Vx
QbdhGYAhADL9WB08YQl2u4zyVDiAP27UDM316WxbRTXY+C7McW9UEZdtDhda1c0EkkoxD2hNZMxy
2bg/Lr2HpplnYskqbClboFQp0VmzmWKS8TdcSci6PRcty7dYIOmNuh9Y4FdWw15r7AsTn4IEfjwG
1PeGLq9GqSkrBq7loo9bdA8FlGoGVQ3uhW5Tm0JvIj+rjBzu1vV5BrbQ0ynyrmq4Ov1F6lsxl7d0
d9lf7nv3JKSNQB8+B7GYQvEbvJtb0nHIVuco7ESrTcyE6x48a8uERrpzVC74dP1KZpy5phcCDHvj
FVyMePAb7QUTPu7fqRUUEnlEI56pgSI4w+fkANTfZ83Kw5Jilx4vch38J/QXmD06KNu+KL5RgCLZ
8Kx+OQS3g3RnMu++xWyQBcbMt6y+BJlV1C4CTGSV6NbKnu0I2hLrZNEVe7nLvq/Akegd1HfCJFAc
ozGgomZieTFKsJLiA7IN43zJ26tHHMA4IGGJ8jlL9HXApLj1v80OGCdTm62HfEVFW7vYp8fEfcue
tCfR33/EAptiYNhgM/AiSe1hRR2KbxOU/sFE8DFEhEz6Hy6SEswWUadrkoXxqep/kG8qP1HWfV4Y
eTaxAyZbCoG8VcaD568ED9MxR9pYFd4TYF3vdvg8LHmwIWdyaqL1uxLp7e518AJbGv7rRb8gybiX
dSgg21d68dUMde4M1yGxriFGSAEWB3oEJSoSb9XUwaqtf0WvMInxw0hJO6sIaYUm4qaVybGZQXZg
H4mGk3aQSH+8CM9Q501JBK+HcJPjxq+6ExyjE6nBUijuvrCJ/NEE+vzRKKqvHHTO0PHp3G3OvjDN
PoxVeHC0m9X/DsIYdLPrGPRYuYgJYjZ/a87XXga3fholkhNfvVXaSDuBdkdCcIZfDLx/aVZ/U8Yg
ehtUI8zGgj5UIochv0uzUSks6v6NgpFyfX5xaVnQYJWVrK9+fkwHFKIH31MtCnZnx9W3Glf5LJ/c
DYB49LicX1gBb5f0PSNcS0oZZZ7djPfMS6+jiDNWwjyWXMgltz1ChmL9TlC4Xmd5N54l7g44wK9A
Sw3GzTMzUfX3YdkMLMQ6CzfWNCIIBczRbqHxBuCZQ7sVWpXm200NZF0BdV/cacYAEeBP4dRb0B3G
k8Gi/i+yF2CfviQJ34iI9B8qIbYHOKiJjgX6Xo2b+3ELbpf/AcMr9EANRT7diykT7r0pBcWjiR3L
q0+1lwcvSbrTQP2/x0Pu1dorl0xAC6fqVPgG9zHmo/qUjWGm37sywEnXrIvwaIZdJLWZS3S7vOcr
eX1YQC1OzV+2Bhjud7BaOL38CpSHb65WVpQqcDoC9zoqzCd9RxHFO31inSBaaW4v7CrM0YhQ1GiG
1MDx2/sdojVEk5qnh1MC5vmPKogDK5dSjgZRyzRRqFgLtrLQnLgN3TNxJJdXUn71WNKlCG0aB/zJ
7pvqagpmclgAj03kecQV1x2Yc75gIWoZarUXiDvrwNdAjnOL1m9APzKgeNF9nnqW0ReBmO1Eyzv+
eJOUj6ReaQhF3AwR6ugg833zoW3ytZz8eRBrkpNqycFB1UtX++VzR7fgmM/xOY7y3d6iHkxn56tY
imop12JoT/Lq39YmtooItllLu2YUpCaJ1qcyiRK/Oq+sqlzozUq5zzc17VJJ7uRQ1tQ2ZFRD0nzx
lssBvMNAVIJbggb1LWbEaK+f3/Y6ExqwZaKyuBGtcF5ouLwaFSJhAE1P7rFoCBpj2neH1V2Dy0Bl
w5fDhoQHVpuSXK79PawzTr5he8A98OZmXEir5NR+9tC4q3JVUiP16LU9VrPJqCbAHtHa1/9BNOXf
DHcvYmrEfwBpYOysrsmkl97asAWTCvcD80OtJSJdVGsBJ76Xwvyj6H/GvQ6GdNAWin4WemnUUFkv
tjIED5hPIn0xP0VL2KjYaIhAKQuU0KinEbsqpTivJYKV3QljELMErna7fzLeu9MN2bmhCNERJivG
QBLvdACDB5aNJqOQGRR2aHtTUNHsiPGwhddJaOpWhYsuk5NDtl8cgsE132/0oZegUJrfR0NvhtFc
zFLr2O+d0ostMP+zeFMJ5zDl12xSSGYe1kbOVcxm5UKu7PsqVFsJPV2d17zWkJxOu/9Vd5264vCT
qZgzTZeSJDqblRipA+mw9HAu/BfhltK5VlUinjH46bxVC9yImNtAsn335wa6VM0Q1VPPi0xx7cov
YaPXqMMUqpnNs+qw19bEOm7vcqlvPfFO10gTd25wJaq3WlBX7R3zldpX4j9Mt4cIzvRfgunggURG
IPvil68ugodnG+6odE+GpfUGbT/kag7y0igGODglzkRo05QvY2WLB9eCk7Yf0QjXdsEEnVLtCG/j
5Soc28bPZLajeQO7l3r1/4gH2Yi33qnkAsGZmxdXjZ6ssGGKlP++q0Nt8Cqyx/GNLpZNXOSfGdL/
/+WExlhehig2x7ubvew292SVfwOXwaWHn7vafTqiuRW80WMPsHF8CG1QyQ+peoa6EJ/H5HXGllLm
sgZYxBpquLTHQEyyuZJvGbNU+UUKRr2ZTdoqklom1OBHt6m/VW516zM8Fx+Jo98brkP5vuHF0QLC
hewT1zs3IPSkN4D5gh8EY6trt6u93ZJPYEXYYnC6M3727jYtXpPK9kCmJvsYPM4bc9Zuv46VfqLL
MHXI9U6fd2NVtr120WqoZuX89YDopp6skJcyeIeQrfr3z2uDQlMah2NRrbJngre6/8vmtKNpFzO/
NWzFwxbnh5JJAEGrDGFDmDGxmCoYCcmxNfnJXJHATaavOFv8OksOqD+15FD061GAtEukEBQOZLe4
FJV9nqh9b1ViG1X4DMJwHoRvPby72N1+fczrLgYy+wdW8UeUR8P5bPecACeVaRBjVyJKB10FN+LA
kF0aLRmuSi9Okl5aRVHih7GhkV99xWDAJzQAPoVW5qzjglMd6DtQssdEGVaoNQk8BcPZfoz2PV8X
QKODQ+EhGVx8Bd9vLUo1EkvlnrYuw2gydOdFFabcQGrNjpn8t1hBHPMcXVMzbhe+T2y4DtxB0nKP
y+Wz0KPs7iAQK6qlBodBmPcvAqP/kI6vP+N4QJTy8cjJ7bYaBLeDwBZe1Pvu+qUQJkQMg3yTL28V
EUo4dTYTwrw1vp2SJfIvxFzPloPW2uJpy6A11lrqWvqxWAierFz+mW1somF/p84hb5tx+eB0yQzb
XKSORcTdzwSfqDWE3qgniQlwnYvOnMF3BS9V5DJup7NA/iirwvoiviA/VF8lIMNI+Mjd4nC+eInB
A0TH7RJUJPmO91J3+MgsiBbcvYqh5MDfTnp2Dt0g+fl1/lUl++3F6wVp5sFymBQJdsO4Ivm0Msm8
EzsbJK5ltrBeRNozEMCkSxD/yy0cqpanO0TdOdBLk1AdPrzNlyed0PedE+ixOnByPcvTm+XLamjo
hxSDlLK2/FSRBdFV5cFaB35OQOGjtuoFff7Q7MHKYSqm6g1gD8mm+80c1rFeBDI5OPUAfVBTFrSl
7sIhpGqzxtvD/ezv4izgbkhnXb5wIXePFOo+AuK2QH4rwBsQuDtkThbskwkILzfxuiE9Y6jPtCwe
Fu7T2LXuWbLeoL2ndLSTtSM8M7ZetknN+rOqMXbtGJwlyAk4qJFqeX2f2gg1KF9HUx3IgUr17rmT
j+nX3hk+gtqFjhdQz/IL0zwWZDmzXalOaCABOIw92xTxhIT+OJHDOwuWSN6IGkIEdc3OOcBrfCYT
xPKUab9/YuPvEMht48Cq93UtNk6/8B65GA+f8VZUX49kKJLsXNYTvQHCmgNZHSu5Myg35aq5Qm8F
/YSwkoaXptIR2Snt3whHsMt8uklJtWMPVa6CDuv5ddh1Sn2pcTKurj33F3G30aGQcz3YhxFGx7sy
ZG2pBzWN27pLfOkwbUWTw1WNsK0SCixTXJXq/ceg8qjaDD6ZxNZ/a4woPaFhfEfgfZHBP9I47G6h
L+BIFn00McvGjBL/FgmbOJkl/9/ZLGxavdkslaXTZueG2Ou4aq4JqWAVQFd6hMSZnZ07DAHlM8wL
lBMSeu4LqFv1r3RixkM6WFElXdstZqJNV4fxd0GMonl1pPZuYzamB9oi7Dtl2q1/TSV+/PjeGERk
y2WuruMdCtpBX7O12LzEW6abceKwL7BtGgH3LynPIZ8Wi3AHM7VDRg5bWaAZUc5svrtJt8u1Qsqx
avlCM+xnHHYhaZR1dFaFXiEambaXo1JZdSidIdze5Mt5DioaGRY/HfoYD3kbAR8aC1Jp4B2Zf+YF
5Jb5ibwn8CYdUDWLyzTgX5mx70O+i3sAgFitBnpqBl6cqSqC9GjVBBGpyb0C/bO0hLcP8l6sf4FL
0htnWUwnzAXivZ8xcqsnXxJyiClzhSGNfHvThDN/By6zLOx6gCv065wj0vNj+oKvOspkQNBejf3E
924T2ccbhZWltT2Eoy0V8NqWNaYfTYMCFhUeWjWu6QC40yH+lXhovzgg49Is2WPkxkCCQNvMnnKT
V+AzS7/WVPt7YpsknANHTcR2ZNdxbr3DOn/X+kxnLs9xxhXihdqNypBb+lim1T04Vbh4Es81WO2I
wKjM3p03lu1N8gYqpcNlvKGGWcAIzFV+TWSXlBrW1NKXfWyciSZhNEp5btsnGMk+ac7hVXgPRsPJ
pdHEW8mFFPvQzutKYclDgvyLpwco1YHGombxpF/mZespvTImmUOatLQDB8WxMHyew7UvFHgVp8Lv
4dm+oHyNWsPbQJTs/h2WuK3a9gVtonn3ZXeM6VvDjfgeNekhzdK2daMFtLjQwqRjSiX3EJmnLP8T
K9vQuI4J20iDkHueH3lgFRHn6qnQJOnohGz2ObiQgBZnRsfGYbQLX88at/n4fXJ+Ii6bhGyX01ZX
VyPLpLt3kdjp4Cb4yE7NJUzI6RpA9CzW9aIOYiscQVTrum+NelOjF/rzOPNXY9x0OOE68Ie0TmWw
4/jJAnbeklchmsy1d4m5c1LOKue7rMW/7IT9RJGWnCGUDk451lwlYUCqmubzz9cqDFN2XVMVfMcj
e677NimgoeT4TVe5IWQRyqRvNrjmE55pL8ommKUUEWxHBb9vBq6V962Lko/blfLAqNrnHB6GCLwC
05sgKUx7lYx8Xa9KU/mR0tUbXW9UIVfS5e8MK8ZrG2izLb+jyf/57dF2jFyiT54n2ri/FWJrbKCw
tICU3rFjUBhjlJK1Xrd0i6PCavNOOoBVWvgoEgc4D9gF+OlfhxNRhDD+GvT77lNXhkLpku6mc3bB
ecaifA1SMR/8OFnEEpSizUH1fbnz9CWH72FkgM74aJ9rH2+b6JW5jMyu+PPCWg3TMd0dqzLleI/m
stR5L+sn4ih8oAGcApr1YHcPrKCHwLEqAiDqfe5HmzkKeIqNZgWt+YEdCYIzgqnfNisDy0gJTI/f
y/nFfCU2cxP/MJv8YYVEXLZh8R9YHFaCfC2TLHA5sca2Gkwz+ObD/uXN2wv7qLEmMH+5uXYnUR1y
DU+Zxl5MArMaF0hxiILnX2XtkhWF9FV1u0DFRFli67PQrHRP5YqbMgMDm7tCRsHXNhkLBHh1KBRR
1R8XUjeTfzbSBy/suZC2LoEWnZ5dOw4zTu8hj72MOKkqehMFcnVQzILTRgSOPFPc+cQfcyJRgvqY
E17jVnHl1u3L7OPKz1EZHY3cfl3xoGmNyQaydCiHpaBp5JMvqTMiADea87p6CGYbhHSLKX2veKgG
DgCdPpjw4c1qYJ52dqXohTT5YlBuXg5ZNIUjEJsexabVhV5n7kPco5KWX8DenXo+1qJPlOxMTruT
W6uVyDK5scRfWZOhK/igLu1nGG7t3fPwLwIoLog6VaRNdcI9CKNinW+ydJxgONJ6Uawu6iSryvd7
r8nCK5zUcE1VJDSwdcrqCXmr5rgfQwWb2hyZzf57gPBRA5wSN5XQyckgbMGj9LbjPR8nBZu1kDal
fvyg/OpuJFWZAV0WLSCjw7KPvP1SoOtG873HHD3d7TdQD1KmZaUPIQej3M8tyKvPKKC1Tjpcj948
q49SddwYqARgnr7XaWH3N5TeEyZIpicE1w4/agB2NEDP52sq1fXbAEUOyWz4UJx2VSUGG/avVipA
wL18c2BDbEv0Mo6f7jgPPzGVa/+9Z+ef6HtW7UE9/m/X3PaN8oCIbI1+012ZVjGY4AWPBzuBj128
GQqpdvY367MNoADP/5dztXDe8uUp/zDBqhESTo72LS7BRg3u90X5aBbfwie4wASCYDGvqOOYbqs9
huQDZ8aTiS4+L6t9k7nEDLdTlJosF5SCdTgd4XcksBLfUzaaF4lHMhvPqefICS7XxuuKahwD4tXc
UMrddiwnJnTGRg187JZ3UTbUhb4JTKZaqac/zvPDGP7T6C17M71csX52jCGxx6r1gzvZcoXFohRq
PXL4j/fU67s/TcXEEmTZdjL7JgizX7u+T9LJoUYw39J8Fz3f5IaAyQzs+D2vTNskqIXwqyZmYwUA
95/owGLRqR1EW/wNgvHtJ35MmA24TNg+Aq1sdETPG6WG5OAVxnMY8+2jLSonzCthJMTG7dp9Cky0
9voxGUuBKxlj8YGecnX1DMF/f0q5yul68vJYo4r1fif689qhsipE9giXCtqfooDMpQc1QiisdN1g
zEm0RCNs+MW9Lyc7ljT/hEBrRO6Qyoj4QSaCD/80O8ofjKc2Oc+ZZG1w36ET6IBI7cwN8DyGPD7J
oEN8uGotSKHHrrIht7O1wKf6DHc6DAfYt0WlXOzhzdB4bM7g2iVhGpeVccz7psofTBPoaYum0Mpw
WYj+nm5vIoY6qn1e3GypM1CxLtLkU/qj3c+P9sovExi7iItJ4ozOwRsbTM5xupz4lKcfk44ESLZ0
eUUx4L4Zd13hAlZYFue1O0kJvFYUDQKeCDq3l0HZkV6593m1DJLmmKjEcy/zciybCgpv2scTb1Vm
oDHstidjaVqI85v4riSN17dAk+zhB3exiraElURjwIINgxy+n5GK8fgWKTorA0C+4TmRsfyV8sAc
i6gc8EinIABl8ZcrsUI8oBH1d8LurNGgPYaERssDCHR3ZJuvfYNPJQPfVO78BAtdv/C3lOC4n8VX
V/2ZbCErcBmsV8+KN9R915Scm0z1OA5Av8+ca7LbNSrmraDctcMnKxNQoNeQJ45nL1HZyPSF6r9Y
Liy2e58VhybX6gaOpoW1fk9qrGXl0o83sLs5ghakErdnNRP6qkvl32jjBbvaS5X4ckNC77xv/YWi
hXmOHKD2gNmSdwA+7cxnIOhnBAQ7Jy45kV8VwK1HGRknMKvN+E5bl+ZEwxdxirLHWxG/1TL1ZAKG
TJT1U3qs/7EYlb1juISfJFrlIUysfdJjfK2fqIgP0WE+QLW5VMV2u6NjUf7xYfyx1qEeHhhZYO08
WtNK+cEaBZBlAFT4dJmlyW9AenKtXRJafY38mCzVnIzUNOkksViV5LljYP6WwE+FO6ZPQOPm/bwc
7K1b+eRf3/K/6BPFjXlBDcyqW9OShI7XZ6hjR9znvwlzWOgSaK0qHmCnjBIYHWKLcqlhI0w1LlDo
DB89MuJsttrlQWT4gmAObldqsoLhxC7t797B893wsYdfxsg66R6Wn1dHOWPkQ9fSoPUB3jIPtCNo
Vs0Vv2DbmOUPb8EqkRzG83SamNp45Wl2T85cE+1oLO6+3F1H4F0FFRvIpC/ltaDGgkkPm8rshKjn
63FvFAWEpRn4gjmgXkEhTK0f0P0q7LrMTzXz7juGaGek1Cplmcsz3MjyVXXmrWx04odTwcfQJrhm
W2solsmnnDI5LDROJaPc+TQcuJLG68RNRMWGTi/gTpmvIVeNPxcKS0PndtzEYsp9H6NL5VavzG7v
HsS9Wp3BePckNFObn/Kw/b/DZ7g1kvTmY3F39SNF9zIdN/z4x3FyFhwrxi/da044ZxpowMkvvLwQ
HCbHN0CIpvA6QyInxWUiQ8nnlYh3TpqvJHj7Np6Pf+kdGIYW+yNAUtYdXsX7p3o+SOKdPuwCYfoo
wePcVs5IOZijBa+KXhqHXdCSyr+l7Qh2+o955+jQJKpGM1zQ2vHbC2/zH77tZtkYe60/UFnVkCTt
scRgAmOJxKOoYtqWwfMGGbXd2oTOwc6u2W3LYXzA6pRJzg4HsalltCvIoJEdU0tZNkWkSHctlIbn
KR3U1gnIxKYS4cxIerqfqU0RagIwXkS8WKA68/YOkj5fDCGTa88Aqa1XXuUlyGAjQhzSnhPqhc8Q
dlJlMcREK0lJidOwLuhi0hOIcZeRoxIeP/enFosvA2qZyduxE5nIgBPtXFoAn0NEblPTgoM+lDJB
PBDpxLfMAbIFK0/Hb319jPpmVHvLmZeCWB6w29l7G0P19BpQrP/9qR7CtkKTj438yhv2pRJU5Vk7
CBPEsgV1MWVs7VVatPuSkdGGQvvWWAW+TPh8UpDIGduMpFNiI6u2el169y3YJh49Duq45qrRMUUZ
liQZfNWg43pWaG1EPOCtIuM/2aHUi0P5+jvmqGWoEKcXwNlNcastervvNci7xw59vHEW/DvXxjCv
Nt80VdxEK1al4uXGR0eHiySRSNqIba89QECLhP7Oko9lz43w6WCCOwECsULQfqZTfM5wsgebSJZg
ughk4VcdhCuSJUbm1kefdASxLdbzWluastnpp51N7zodqrdfaYiFOAzpIhaAK1A7P2QJ1c7/Lqdm
XprvxGunz4ktLoIFKiVonRDM+EesvnZij2+kneTGike/eJfg87+mn3aevJ1zMJ6fnTpSW3a5F/5F
W309hdW2UeSKqAGkwWjuPC/wMQezrwSA5qJiMDEqhPgfSqX5qrIip6bTmaEydSYr4IMAvVxkTrhe
TUO0raXKwId7yUBaerkkzBtmoic3gK/KjwPd9LJLNJ+nXyNLxTM+jU7+22EIZElkb6FJHICTjbuC
vLmJk0HS3Setmx+WKQkiLcl9+arsHv7Go/SVN4s2oSJRpHOEC9GVsKwxyXr43HvsRLEwDxAEMewJ
uFXcpqfcOgFXzRccW+py52CQw+fsBUtJzfPZ5IKBomyJ9kcSe++/43JUrUx3+wHEDYBEa4AKaTeI
UsA54sJzaQ3zhW+BmRfaavbIFStBKWJE/zxIEBRU5ewQlDFc0fyS4XMu8nO83kOU9FGLGRBEoJ43
IHCqq3bMuIaOm0idAmKrlUKtwt1X1snxdOwRwQUHY//Y4ezvQ/Ihkc6sQB2UfzdH8WvnW2rnTsq3
oqb7vebX+5FAr4jTIAlVK5cCyhZ5BAhRp6scy/9xr9ajyxBE9xCw+Waz+Y4W0bKwCrL5dQDww60Q
O94ZkDAaHDQTminUUkL8iuN7lJd5UJPSFUsZMO40UtHAQEtEm/eVEYPV7+xsZh8F9xP4YxBVrpol
eYoM29cvdAZ1lUQtxPdl8MYWPwOI8hofzwsUG7BaoF9V4jvcIW8280Bgf2pkMFZ9tURW2yvLAhbk
DI0k6E45yZLJ76Um+X1H/k6g+EFcnRgLrqqO4K3qE0AHNBrS7wUcpC1mbOsX/mAikLD5W4i5B/Bn
FscTN4GJ27aZWbGRyZKFQJzYqI84Io7d95BsjU+FA3c5aqUB5PvjSdkVGwQTZxSt6Z9UJPy54m+y
PwFw4g3avTQT0EO7iKf3BkE1Ddi48pihyZqBYM+u+JIvAET8pZwAashlfZfVaEZhXsv+ksnFPv+M
Z7pz743FkQNVtjJdxMMLRwKOQogSSHk93Evl8JgxsAMhrhpzHUXM98cmPnXI3TzXAOFJaWCbWDeH
AQgXLfdfimwBFY7B34YpLHwf5cUr/61UBb3x/JqhopkzPTVZsGumaKGgY0UsjZ17IMSPuOpajAX5
/HaPeS7TAuUDH0k+ILtCfTeUoQ8Od+7M8iq7p5WhTB7YpmJ0lVXHeG1U+3sBs/t+DeAicu4tSG8j
EkzmszZQQzTxgnISPtBxJgtbVFjIaOaI9zPIATPdCO13znyIe5gVTMrjDasWyd7MOijG5Mh2TlP9
K/DVE+Grwc/couPc5rxEi5a67YAtl9/b7xdFBAWBuglFIEq+jaE6EdFKmGw1S4hEQoAoDCFRLxmd
1Svo28Fa/Es7/896Eu9kA43xNHhHuMjolycNZqgkGqzFiFwMOKwjrsQpnYrDMjcOSziJAe78FXpd
7W2L9bkmRapNKLS/LjeEThhuFL0TfGudFqYMYOywGox4QLELiCVPLFq1Z/kJBIqo2D7Nldfz63hI
T+yWzFPlid4kdQchDDZc/AqMfI96iT03s56mcZxJlpxuKFohrqkgN/2WCtMKqsb8Bhum4A7RByuu
BqxP9gc6IDJg5g/40FXaomp7aJ5PkyXLr9OFxv4NNOhMG8T55a8ouebu3/45XHkIf8fLh7Dyu2vr
JFw3Pv6xIg+YUf3JMIWVL/WELaNw2UdfFBCFb9VVWXwQ9hTHZ60jVdD0bN4qdSwcqRgTN0YXdJ9L
djCKrsDo87J549ZiogjsH80Nyofz4fPe1FTZmEZQg4qxnx4KjFxKQXxPSdLT0pS/2C7LHcRPrFWe
VRC4dmWAl9eF1+KyvdWAKuiXlN87OoMtHxE1gPjVDX61QSQ2aIKMI97g1fCkXoncif9JzD/zPRrK
rwYGTO0ctpXfF/bTO8sPF2iWa0O+WBUJzH+tDt2FSCK11Eyt0JoMVUUK53VCNky1xpuM1nYDns59
BgTKqtfE4fMEDOuGBtzl+XzrGNAC21CnvZj6CP/m04gnsQuRhPYUZuWWWhN2LQUoHsrgpwMagKqI
RsqJR2wzHUyxE8+RT2BLp4BVC9cPtgIK8WD5CwK0O4+h63ZLtE2jmlXInQyaYAlmWExYZDnQQQHR
d3O0ZFn7znqkgVNGpPSE85g9fXikuZ40xDt1M4hJb/SXVIXHb6Y+qWlScM99wXJlWpupMT83Pi15
R/+41sbw/NPdVNSe9j67Sw877U19V4D7Ot2zDG/hFm+iJNYnNt1OgRG39oAF14oCzyItflZFo1WB
Y670+EHXBuy0iFm8HCag0X/J7gM+vfnIEd6xRCH88hjm4zVYE83kij22EmvGRXCrArFsXYmpCIxb
aZ3esDiuM1jLEizRNoD2QBwzw7TmzUHleU1N2fSzn6DVIJcQOzxQmR/OKNTaa7pQad9wkymNgUps
5QdxnQK1h/9sy2jrNcOUKb96nU+11u2kHBxwdELH8kfIU/djRbhApGWXeid+IRssx9bPIl+Ejv04
n09yLrk+OUSHa/O0F3Ms9AgnHBOJ7495diUeHT4pqjLy653Th7hpckFgjWlpgtLA4EGSuJ+RLBqm
kqE6YXQ/VfF3ZPsDU8/iqYRSLxnVPwcDYyGKadcUpRIDXIBH+4WeF927sMCJxmjzjdvUbSxFF9zS
Y3deiKKyMsxxQ2JY0yGB9bpQCvqW0CAv5efcEFSfcd8zhfY13knBeCMuD31SdzWCFP3+L9hQmrj7
VncMnPeYYRsYWV4Ogm75Vxz3DQAiRVmRGGZvy2lBaHwSd5fStn4ImzlAk7RUQc+9wxw60ntckLwp
J2uiEeJOcvLxPdPNz64ETPhnWjpxXsc/eAMWg2KpFBzCytjznpjAKFM3WjLpjiD94m+yt+x8HUrb
RlQJ/AqJtLnADLihoTq+3lNxBr4OK5EZPPquit5+oRn6RV1eW0TSpA9GieuQpDlnN6Ae21VNOfcy
l5mmkBYqkNs8GO2n890DGeret22LOGr0iQVRQEJxKuTm7cqH/Tovh8+uhTdKb1udxjNOKNwTp+Ub
yufwxyPbZBC7Uqt05bpgQezTqulcjV4WvoP+lSUG/XUFElyBsqoYsca+YzjRAz/a2nvYRbct8sXh
BHRQXi1QMnP6tuRrVVerzLZhEN2dbQu1bsiIyFDijPQrxVLx03AS/9Hlrb1Rv622yVHV54kyRgX1
tUG+HXHHQTAsn/5tlwg/SB6LDCKo8KNv/s9VWUICYWkdwvpfYc3/DGbT/oiA7n7sBj7Dc4EhFhVK
y1IpG/IONqYIxng8BqyDarURjdHEWR8dXqA9dE1H1vmVwpIgb0NilTiXNBoMVr3VGNVaWj4tVcXQ
KRrQeY66qOCAj/8VCteO+E/CoWZ3lUNAV1nPLx2dAQ6E4fQ1z10bULH4pWT4mfpk/LMRuU9IetHV
v8/9SNW6OlYRSPiD10MzxGOyd5807RGqNA8DZCaR5BIOmrabNRqI5SHjhSv5uzxMWuEhBop+hwlo
0oIRYcKMM9n75gAAhsAdyT45qz3QgcWF9C4PqBm+asaJ026woqaH4zeDT4UG8yIUnVDC3T+gUBLk
6pd2hOjkiuanhil3IodUN6hW5QK3Uy0hGHH2LquICn+TYOXqTaVgcLwNw9eOyP4ZrEBON4y8nCBn
/He+e4EeJwcI5UN2SnEYy8TLF1QJjyHpJJua9Kt3I4WGe+KUASndQflIf8bpgk1Tu+OSZcDCyWOE
X13Y5eQPhGoVucMg/1BxJo80FLDD9lkXBQRm+/bA3wbm+rR8HoXrTtvkaP5rDb3qXJ6BmiNpajn5
YCraWriWZJySJ2Ki99hTD28j/bpRLpmMCgutTbkJEH5HVpFfTGQtYqqczlLHA9lKp3hzX+v0Q2d+
Yomatv2WZ9PQBqOl6dGMCPIg7SwtK3XspD4q5o/UPzmNEaO+EaEqpKvZNQu9dpzRs+NZc+otCSac
lET2seJXbByg1U1j0xslcY4G3h6BrwQxs946w/Kg9G5qrLOHb+d6ZJ/Uyccv8pM7Jl+Nu58rpSkx
ea0wNf2iRrtYDGbsxMS9cD7Ddl9IvI7vtrCit/KvkMei0eukwEAfuy62J92gG3nWeXyIBg9Rf6yM
hbXCBG1yjjQrAg7jUSURDLfV/iHa1gJdaGt9gFVUn5wr80W2DVWDk7lh2eXZrOVUCpUWcB6nOa3x
D5C5lvtRq0MTn1Cf5PrDTSA7CV7YrGFfXKZmo8XkdwCqe8Y3LZdFpKE1d6JK1OVE/dTOWz58cjGK
o1QrnbAUdI44frNj2WFxoFYTBDCRsIBTRHaNWdu7jkbJlpIarfAaXzvtUcboZVFsAtQW6vdJKqkT
2aivcSyxGucfUpr8V9nBCCXjUGuSF7aLWeJYyXYNTl1gZfv46TjUFWuJ36tx9lp8RIfB7RYQ5gUa
oqXtWrUv6Qi9F5w/l8OsDhKEKzEDKsJnZyb6YDNCKsf3lCm292/v3fw/dRGTR7HmSo3VBbNcGXfJ
x6tSySJaiaukFSvyXBxlJxEOJW7gekFogTyij7OL8Ng9BhvB0ajaUFzw6mJMYATrcOZ4P3sZ7R++
37IWsccipfBbcqqIHlLgSut4X3Lfdr38di/Sm132HXOPf7tcMCzu+mXSBorh/N3us2FGoaXBKZKl
dY0CiDmmViDVh0QG8LrPicjkc59VOHyiChkiRKooZn4QtQLMWvArQnm1rbDh+s6GPSKRhUKgR1Fo
WaM74vld78OM3NwoaFINbQxWOwCtV4zg4kMGvxIyJ+xj6YR4Gf1gi7sTtxoIM4Fb4/ExCGkV+45z
wVLPPkxxsh3+T8KFrro07loZ6xo3xVhD0jyWQsBbqW/XHYD8pms1JAngtKteXg+RoSzQtAMiUCNR
3IBRncNbhz6wO49+md+5FlFspGliCgz/JZxMzk9A3P41IH62ArHntCYL5IN+CK18UuYe3POs0wqk
djBZ8p+SjjiD04drwhfYPvI/Gcy+lZ18yw+BMwLTdu2ppuDurj8rAFptSeVZGhZBoW6PltpcuLyd
/EnQ4LDVfacfLXUbMU9c8sste8Z1I00gBrLmiRIUfIhBi83UfsxDvV6bmEBEVAl/wFGDsXKTwPlL
oKRxn6xNGYkVCEKojZ50Y556EtmpW8rVaRJWKz2cX98nLxSIdELW+p0oJqn0AwO9Q5bvz3Qp0zkC
CR6ZHr5nw+qCxoMxk2K7cvqHn2HsnXX13BWAjrdgK6bzYmr4tSWmnvZpDpZp7Y/hSIJZkd60tF1s
txE28QB0/8sXDrbwBAWoYNw2nunyOCZaCabc21y417c0YqawXHEUId4IFwSY0PtG4/IMESwr+AM0
XwqgiFAU/Aw2hVwQnM/vpVPWs4+92uOEDwQBTi1K5lYv5QJq467dE1zrfMoUGaPgEHjshRBc6fHJ
k4sVTz9yqh9BpNadHjXvYyw/PRCYHXk/H5xxA3HBGa6ICMok0Bqz2h0dC/Y3VB13zg7WX98Ng5jB
L2JTWbkbfxRIjztOPQqxU38iFQUqxBAmaNjXG8UPKH3WzX4IMFoBPBH2QNEZ53okX3RqA/KmpTQG
ynTRg2YFZDRHMQB8xorpG/dI8pWmGFMmH2R+uzEU2z7yl8ebZbi2ZWAS9tJyFL9pM/C6ljNEqUR/
0vc0nwei4vCik3+UY5qEZsHJti+vfb6+sJFLD8PGYWUgoepNEG1sJbbWdhFFuI7KeX0pseAs0Uxh
8kWIXi3PB6vD4CnzyIo41OkgWLHWZWHi7hptNutK9ijX9s06K24ksDtY1/2vWFX/SX2gwmWk6MPI
tfAYLDel+SMXW3hSXHjdGFg/nfzpq1arHDnOhQyrHx0ozpYhJAObEMNtbAGZsMU8h7MPBBtzh5JK
kwVw30Gb0UNBmtP6H7KLVP2ZyF59O6v/35Zdy1ISQw8hQkfPkF2J3nMbHMvfLV0P0qmsE3VNjWsM
/FpK9G9ytiZGePuTwRVtlumSnXVh0N4f8NXXP3U4TL16ljHrvXc/tPnCuQ+N43cNCiclR6it471u
xt24vk8e1S49yOqZsgrLgcw9KIhScveNuabIg9AIDHXuJqSREQ91m3RQfAyTnmEcn8tgHE3UJRKe
xODw6kP4szhdJ9eB144qJrIZYdy0qMkWoHXobG7Zl6G12YV425Hrrhgj9nR33aVEWzYauYrqTRG5
xNu2E29NMG6qmy3gsFgLUbM88kspkPA17KIIgs1xh6GqlSqVfSGA/mevvdmWCmxrQrAMz3bdLQIf
yjrEBf93fvna+1t/Big920DE46S0UOgdNzn0aQNp2o+onC20eb8/uI2YALjZUqAek7CbbYQ9rGZ2
smAEgOeFLYvCg5Aqd8BirHYqytjla1vbCEY6hQ/HMGCxiIAb2I1no8riSq3W1OgXSIEWoeFNLlDn
4D5P2/uVlM3juuETYwSvDEoUqDRX6GXpSs9EOUGZddC9kIS8VvLXKXdCV94cXk/KiY4haZvmS4Ey
AuZYpNQfTVOdOcv4doeHMfWQniJ3XMpX6qbCbFrLNl9TvJIBpbuNnGc/iw00hTXhU3KK0cXjfalU
uoLPw42Syd39+IgvArib6jTpMxXCkgZABHg1FDOb1T72+fdDwuC7sVfLI4ERluRbTcbCSXy2MzwZ
YgfIqYLcCBlfjtZfLNJUa48mSBmWHBpJBXgslTWbyi4zEWvI5MUmukk6JZ6R+8b0R6OKZ080DTEk
RKtZ9JLK6DqgW8Fn2hXuCqdr9JNR8izLH4syE/XNPeyV6hLVpM9c3utNBOQ/n4b/T5aaGTmwBMY7
1i3NPn+eZvW99somk3WmfTLRk16Bp7rMQt8dH33BhOSbfumO8yJRu/agAfk25gm23224cf3fyTRe
3iEAYr/QhShpWW15jplgTIIzKsmQz1Ezu45RONMqzwmt4c1rS2GN72LNE4ByrvzPTjORdhWOtS6M
OIjnoWnVC9YGNenJpQlrR4bfUnrtOphRqCvf14cYUWmsSnviJ1Qu3qFsutG3IcX8jGIkKSdQOS05
iRTg7jkDmBAxc+OUSiv0OXlM5TSRDusCnmZDPzkRTph7nADNcapoTtZJNwA9ssbSwnDB7xgh4kTi
PspuGYd6TtzVh8dBhlKW6yEEh44iD67MSf4LuHirLckd6TIubD8mz8RErx7pYHDjkY1ZjT1Voxah
kBlFDwlBixuws5YBLoXqscl7+W0mxkOyFiCsHhg9ngbHIm0ND+VC9fFoeSQOtEl0sEcgBUGLrSrv
FETZvHoytEole3a45bLkchzupjyi7FKc5YWyZeaBHW8uf8XyeyDY+5P/YoTfDt0ZPGpMpRgqY2LO
sL81kQQ3HnFRfnKATQfx3EeoOZM+WdFyAhdf1uNVIDDN8WK9u2Nm3QQL0ki0oNNNwg9P992oxrh5
43TAj1BffkFcJi3FbGccWrD1dBkEn2Li/Yg0dQNGd5tak8r1ZXsTUxqIZPMWHmHPm9OWtKCGRQkU
1U+gt3F870cP1r+V4HqxFIXJa8t0rwYYwt4bHwPWHRIQZO8+MsSjBbZpsfJEwPF1c6vz8G/bs8VT
qXF8uMzj+BtiVtMLj+P4PM/o2PI1VVOBZo7b7W9iwcbpwW68EOOEKE2eg99cbW4ITOaDtpWEpeuu
/00I0HOP7bDUSP+aLbk3inuoB+2kv3riApvrrnkle/4vqzbZ19dCohNxGe/KsO6LQe3NRI1CLyfL
iMG4KXTWAhDay4zzIuNiGJ11q5ArCX68sieRTnlRU5UnDD7fRkzvbSFTCei9xtz7OOneI60CAZsc
70UJ624js2aVRKIvKz/HlujQiAjFViaYZBZT3ArRzs1U+HAe0W3/5BdXxmnaHxzsacXeeVLMm/TR
9fSfqqjmueiyN8dJONCdWY5273RPGFT7TJRUZNuDGM+NO/F0wvg/uB8Aa2yuxXZ2jrWxKKmF0Kwk
uQmfucBLPbBtkpmwzbr3zapjlRVoqA6wBB5iZIsLltK5EOfQ32VUK1pPNqQZnEqv+/Q6L/iXM/TB
XUZrQvKDp2dnsxWBtJdOMQ6srlIkMyclnj5gxDPUQ1lwnGBUWBtaxoaTJX4SIUddRGoUCYauDEY7
CFnOw43mn6+okpbuvoxfP+S09XHCCr1lBN7TcziCMvYUH/TC/qCHOuTUYsv42eoyq0MuS70uHMUk
2tqSE5P/y7qQNKTHbP0PClEmiT8Z06jSPDxkwfP0Tr5qAsYcCbX8fj/4sH3yFSWL9QELhZDz6uL+
iKVOEocTVDb2pBBL1UGJBPjjh+iA0TMMc4iVD/YReN5K4UfMxRKn+AtxeDFF4zvqfP8tZ5OmdRzB
TU01HsxeYMow8F8OKxC7pp7ySZbCOaTHET0e751zsH7C2dElLenQUOeTm43e3dMSZKsVswTD0V0w
5VhIJTjHpNNSibd/YNBbtqVuWcCbzVyo1ZGLlGHz1ecNe0ZLMVZ1bcdKYFBIWLFD+ybwGYf9BXNn
oRGb1XfLIsITiPUZmrf09D3vixNA88OOf9S3R2lQSXcLNeCKUnG98CiYCq4H60hmnz44MYvJQsHE
eCGD8ukoAJ9Z8SMgEvIVwNQiI2mLewO4hUZL3jarFagwddLaC6bX5jSfkqGhfjmvLv459tx2r9Ek
rzZRDQrv/HxBZY4raKNeBGwYkueCynydyYH4KpHlrEzgYZGd/jQ2zLPeNkTxCGCH1qiEkCPqzkA/
9EoW4/hKIWJklATl9tcDLeZ4YoZiz/Z1hkQocn/3QfVStLzqmMrnBOo9lCxH+xvCAauuDpLnliyy
47nPyRPry3kYOfF7+2m0XeRQ5QUCWel5oDZ/bJ4hzDkI9I/1FVj6CjAVLNFs3QGJBXLHcZTCTj7X
M9endTxV2pctAC1JlpRpEJf7nwwvEe2z8Y0R1C+WhdYuP1x9WqxxfgvWPWTlLKKR4UtSyF3F/qkI
6mUEGHoJQUx/ALZxHmaWr1XCyhQS3y212hRR2dMBYko99olCnBuSpgemstFoB7kSnTjfLEgvDKeY
B3neb/YQQVq1F8BzyHdF+Smge2c1slVZRPqnXHfqQhJ8XEd6kZv1Ek923QXvuLdPXXX3p17zt2hT
9cCCXD7Y+cb9Owcbyg6l7q37It8UDJQKs89f2LMRC5jWZ3XM9LLlxgo/NMIgcgS+SxP57RdOvgfS
kP9kgXJoET2IS+kpJY5hIne60oXqeL/l9Fk9VgZHWFtKo9L+gOGwS8lo2cKEVyLZn5As7Tu42U0I
ktE2ruLpNi+hQhsClNyUNtvF04fpzzufc5PCzElRhSpOy2uf9poe/snWYzmuVUUWARysjeH1v1Nt
2Kmmu91/eZvUdCtsYMn99QYzni2P6Cm8RmgdtOqKk02nMxeunm8c3g/RxsCmPmeah/pvB4TL0t4S
nkdUzHcejo89ElEB7z8bK7/Bd8F+uYLDnJRfdzFngnillq1BGABW0CIeBK8Z/VMouSxb4Q2WcB72
+aa1k1vVe4D/XJsJjQ6oXJ6Am6IsbDAIvVst9+cr8uMCZgYD/L3oErhhYpJygUopLfILjLZjt5aa
TK8Kw232I4gj/CAI+HTlNq7yAbEcF74txxbmqCWAISTQp9Nqx1rMWUecNdnj7vKSk3RTVy+mw1rp
Kz7duhuPGAc9XXe7/Ln8eyLSCjpMDcCfYGeog66wuxzGA2lCC1xpTRSEsEhCfnf4xMv5fgJ0ZmAE
fLU7xXPQ901wFWnR5+Laas9NxhDQtaClKoadBTIF0UVub0jGylCavC1ZtAYhSVKUJMYLLqJSSold
YXKgsjl7Nx72/EaUxdvk9HKne2idhRnNDX/T3KtQWt+x0f/Pm10x2NX9r5EA56Aw0GoOF8Uao1jt
UXdXoLF8/SfiqZu0SnIdyaQfWrSY+f/cFSkr9IeIEp7QsdcGDKW12U5aLt331mMLa7U+KT3CJkc1
nTVqLBcxJV8unKCdbPc+qLAI2qGWkKVKBMO5BTADOvKysIXN/zGNJ6FYYjhKOBgN8BdxfHIOF9/Q
V1vfRPUO/E6qxGN6QTZXu0v0KE0VvepicbLqeFGMyS90etJgSQUIHCfguKp3TZgZSJykyn0tLSHF
OIMmvJKz/LFxYD/87A8aOiQuwRh/6X4XqQB+nDa3iqIaFw6QLeWOGMyr9tqzv/ClwgRZg9QdgkSk
jEeNWbmnMWV04kOpK++/AJkVUBNbuAOB/xvLqT3B/X7xUYXi8xz5X8MaTf+TcOwd8QWHCJPFvaQR
dDOLt8pEjSVvBFMTnp4JwBrINtSDhvaWIIvJFymSQmHNXEDxKHtI6CSW/bFP9Byf0PNjQhqxZRZA
zKiZE1uMERdPYCDAjWo+/DShiR0wMFhejgnSfr6JhxzJseMe1Uw1kMRp4JpAflELsMlydBOzpnqu
+vVBtZtNC92MtySKy9TxqX7Qoc6jPWNhhB+rOYVo20qKl+z+CMtxwjiND9v9UKVGWOYB1Qd9mN2u
rJdTu6EQkdMTAbp1qrwJHTUXOiPL1aAWZXxozbuw72L32gVFfNQwIcU3Xdd1qGF+fvF1FgoiRbOt
RM4tZln2kB9F4eRJdsaJC8hbe4qToZ8Ag8R5ANzL/uoAmhb71IbZmc6Z4ttAWTAAEZytXIRqRpBw
eC2CvEEhdqFQz+HDDLoY3IcTKcnUj3ny94wzXWmTFAi34SP3pVb4+KZDCrx/udod0IsmXZTgbiLD
ZiHzPycnQ/oRHtWMNqnTKbwSkOTpu5ZPg23Um/I3buAj5nubQ7zJi/MDdoBKAEefymwah+/10+5c
eDS157hO38zmPFHR5vLStSPAycYu5znKfJVdf9xLmQC5feCMdwXFY6pCk7/0LVbEbmEg2szx01J8
7dm4i1WyI7jTyDqYOcZ8zlC1d3043I+/qbRsCHTx+7pteQIl0qDO2rBPiiZC7TMjJa1oYhK95ClI
3N3699Mv2dZs6hv/UJYbGuC4mPKzPq6SL70oT7kBNTQPc1LdsPd8ZC3aXRQJ4yoGBoXJ3Ml9ti3h
S3NqeUEIbynPSXXTgMRe0AiR6yiCHsmDVVRkQyZ2Wzw05rkEezOErMLSGgw4Sr31MMFMBcdjTf8Y
SI9OJmwW3aLABglgGj8CBjSYJcpiAB7J/4sUUFB1ZYOe/FZ5WOBLUUjHR2Irhgxyi/74ONgou1YT
/wQENuOji7mIR4SIpXel4QGTSKi0EuyyrYCUjE1GnKNQvfrKvkKq719YSJHeuVuI3lMWDAi9eBil
PYBudSkUgCfzzD7wS7QCjW+ZgYmFN4DQPwE4MdMyGcjTDiF68Qbh85xs0NcGMc49CjjF2Q8+xAdb
pc5XvJV7jqnrcTj8zJFQHbeX8QH+SLgRy3qVtEsZrn9TrtEZQp0qLNbzOUADyNxFgd8/YZ0uHY4g
nIOR/cCybNnGzOYaT3uVJJ5yyHq+9y2dyy4mwXbiTMAhSfevloUG3JId/zzPBvhpQgDJyfX2Wuf8
Gs/doitVtuChWp1rOzdZphSlSNrS91CddL7AQtl6REfg3Yi85vP1tf70l72lwnD5c3a0q0TpdXTu
WyulW1zLsIECyKDObyr6wq9J9Gqov+2OVPjzkH8B1NMDmcdBKXmQ/grkMqkqUxv85HX3uHAUk5w9
HP20znPi6ZbGIbe0ndOVk7SKN/LD22ayBiYnTH1E1hf2GWwhtjvgCMNO6BcE1ljzZD36Lu9+gXUj
5xwmuOu2Vh7gkrS1XtYmY7mY6GIAp3Rqb4Pu2iWpkALFEFRpOaXYkZXVT5QuqUhkNAN2OpVYJroO
YD4x5Jq4G0RxX5S7rHRZxBZg5DceOLudiK+XTB83kPpiNPfo+WjvESBM88BxG5eFA1FZ9/uJRUnj
xo7kczJyu63kBOySMgBLXEkzLq4qGGs5jz5Cg359iHABLPbddyAfCXjtF5En9DPuD5545NNgjp7U
fcXhPgv7TNfT5XKBUt4XmfBrIm3XIj6DcOkBOvTlYozyW6yLOYZY9WMeo+xfnBzwBmlZvvVH9Pf3
IKmMzsu2OlRXKEHBtJViHPXzZZX1+VeiA4yXRA/WnJsPKKXA130J+QZi7jSIgN2M5mVDhosXQOir
9J5L8s7b/vCFkS4iE2FxvcUzPIkzS3LfIBN+M6WwBzjjcR7ZHdeFrtVvHRaiEqJT2byWZEqyzHaU
jdjEfc3xbRIk+JFviabuEbYnc1xUW1oQEuMi5fwkPrMTmZDJUl4scbHTrkbWxt1964ZBopWEqOco
s2VZqO1xnU+lm1s41ewsnl19jTmm9IiAGNM9U8WsD3MvDkbvgFxtji63EOjUm1EwrUaFbj8rZfGW
SpreSKJZQXWrQ1GODVQBKww+nPGBphv9CDM16HHsVx46trnGF2g+NzxMjg4DmsaHItlyx34FQ2+t
tT4t4VR6aMgFgvrk0EvwPEpz2ZjkEYYmYtQ1T84h0IGt79VWCNPSyEYzMwD7C6hCkQEZCAQwCEuy
tJb+dbaDkVHDzwSUv0COQarVkTiF244ZLWU5mDP6bRUZ/lInVV4wjDWQWj08itljmk67Wz7dd5kN
xrYjj+oYaL9cUt4noLUwv0WV6SgMMHsg7uzMCMHcEaPJHFpG0X0fqnNWXc5zNCFydIAHOkPptM9U
Ad6ZZ8MLWWEpjOgdaf5f4leTfQT5uZotwLe3r+yUHUHiwcZsfUlhyl0E14gkrZfpeGrC5j4ykv3I
7X0CUgStYZW+cn/sB1xuSPF6sqxB11qveh4pZrsRLvKmNhYjr+wj9ML7vQ/YyoiIQeNfH7utFpAP
eB/cL5bYvv35HSwIKTNDQCrVosE7en7ZbFPVqiZWQ0Khc3FWZb8CjtveXaAOGb76pmJpuWoWPXpF
XRHPODlrDayxrPNfMvGUePlFqx+Zrm41nYZxfb6YacLlJGmkXzZNsgW+87uibRLSOfUlNd+NUTvs
YdKjIUgmv3kuQxLQgy3rp8XwWSD52wssWJk7kIYIlZeK4JE6oo1K+2Xi+mIS9H7hypOR/CdyBXB7
UqvciFZbvIQHu8L0YMTTuGxTaEJZLdtyotwHVjeMc2eUcnBK1bQlmgwHuj43esQ2Q2Etfa1YuqeJ
uDNEc+voZBpgmfTz0QkZtGprJSfWt9I+fgLrZ5/VYJXDaNDvqLhqfR0RIDGlv7nikSNzP+7nYFUE
SrGh/NsdYTdXksTJP0zY/O7BBwVEWbiXeZ+iIHqZnHrLfBwUO16oiQh6hsDkyvSSl9vlrTC8+LSq
EMJJav779kchclDSQPjwXmBXqsJ4dgOcQZUcVWrgxkg3c6zdSncrTFLiqe13Udr1kWNb9CP0YqAr
jaBZbZynT1UN+EkRlYFSNx3rHM2xJjecuLzGLU0sAls0SGND+dE+XzHg2PqW7y/TBOF0XIy4TGO+
hlpIEkdqKdC5L0ulXolpxORr6OYtsu6+UYy0nheUHIoQ8b2kRoYWwiK6dRWaLxT0LEpffVh/h9TQ
YGGnw5vZa46qq569L+onIVzdea1cNQuluJgdY3MZzVyIH/0twHyBVIpqSIboFfIswLVGGZAbLm0q
WKyqEp8/O5s3DRzkKlzDQKzLt0zJBaLSMn/DV49mzatH1UHy6g5zncl24dbvH8h6yqHi0tFel/tX
EvcmgAK9sed5ZGnYyYDugyybw3eOJFNnza6v8Dw3BzcasTIt4M332qffqoizkx6MJjKJOZGUCUm0
cwREC1YZMElII8GVtmZXoVlM2b6nF0s4X/MCVhfgqBNu399AvjF6F/lSFjNsL8qn90EkzLVmJmsQ
k4IZ6OMLJtgJJ5OQ56MQXfRJZuxMldRCxITab2mBNUI2EJ/XnvfliYNIpp/ioLnkopKTroR71+uT
KDkltJwNFXX1AA2i31FmTfWhw1gxsM+6ZEZ6dBw7a8RNRxN09oDNB/knT78LoZSoHdas4KsUOYjD
1rBvab+KvWYpdPuYp2OEmqfjWyAltlsddy1o+g4A//NyDXQjnAIQ0XQk3bmA8KNd2LQcArmxguTx
wR1tjFGrizTJNAULxpvTD6gBCBb/22VslbkpJS5UC9F4dkFDxnjHc997thyWaWCVTwVLY7wQeS9M
UQHtPWqCZ08Rsr13uApXebJMK9kI75Ifq4gbEqtgbJQOwH18rJ5aFVfM5RqrMGwTY4R4LgWv0xJX
9gf+hbBE832pL2QPbNcBNGfPLDGm3wE5mfciksH6Z4uJV7Csc4/BzCK69HGbQFMB1F3OXRbQYxuQ
WIhrd1hKWMCAvY5OBkTa2fUluzzGR+2fNEUL0a6zb2t/Zd3uZh/qE6UQAf531RRQ+G2BJXaEjtZW
9sfOgcVWFFbB3PctdGdH/76JZ62KmIcQswwBX7wyA89TKj3RqyeOpDtGe0rHSTzFQrvAIvNRhsju
Ln7SNBa1wCbQyexdaiQRxm2ev/4cwXnkyAARINVD19AVBdEnIqIwdQfqWIEDy3Hq4LVfu9OkC9yA
rrkSkhv8oW72tRpv7VadAmBJkM4q0BrKCE7f3z1j/I7av3QLWpDqrhFARUN9S+FCqrU1HW1JkGzj
2Zej1jHhAOyI9ERhyZAomN4H5idII5gLPWEt3uzk/oBzxhdLxQoq2OZodb0ESvU5P92A1PNPwTNK
t5CwWBPL4K4LQe27nzamp32jTUd2DHKSq7KXdNN5urDrrqR0Z/WTVJmjQvYn9irrFAA8anIZbfYR
DBIzUxA0T2XhsKzpPNFTON4PYw7nvAymnv3osxGtZ/fZIaM9k6OBXXx+qwJYhJODOSE5NpybW5JQ
CRt/JHLFn1XAqXNIry8AMrlKoY+BX6962yk+Xpd3l6WwrDOXS9ZddanBvJHnpJsB9Ck0TuRz3jI1
OowGWOOToMUIrWKnH9y148EGaGTyVPOP0NEr0Qcnw0K2SWGuzQdKrBlJMRr1av0LtDTdg2H2C7+X
rAFr1gJ7rKboc9ggdUg1upN9S+KXWAqiF9rGsbaNYPqfh1JpTrEDiAD6vV2MSuaobUH3+WACt9US
W1Dz9RueEbwkbAkGiBXhBI30sOFp7Kl2/66fcOFqr4W/hjgJnajLI+lvzRIfSTNjJ07Sy9QqTL8T
yuyKTcEkeQgsxoLFhxBpsIEiGkg3pvLV8nVJtIY1Z0jTGsXniqQXGzcpCwz81O3iXf16+sEy5Bsa
jn3YdZTN3pwyw3/PfyTaSHxLDU6prUjVTlUsUtOGXjJj9a9OCVj5q7O5RdxuhoXzMNy1n2gSZCSH
chq7jC5N+/6hIMvDNBcAOoec3d3S0d6dIPYTRrDQJhLLYDn6gsMN0pjXAPmAXHk7v1MNRDzkhV/G
yadwcBAoSEv/kDEM2NaFubZb1cpJSkqw6gOKx4iDihdbIvHVgm5mSPf57wPRKmPpBuJp11Fc7g1R
c/7cIsAxH3N4IJiX0c/1gMbUhaSujFObVL8d3nPYKybALQJkuAY/MXvjtsSSsf+v30RSdTVdYlp2
dR3+jvWvzptLcfM6IXpa80PqP/vv5jFJXXy64tIE+CG8TVD3Trdk4sUv00JtHoK5oVZHP2liuw35
JDo0iyDKDE1r0FTs2sm6FMXqI752tIIL+sEj4VL3NlVe+banCVxTD479vnkQEoZWS/Ev+PuZWFWG
2SPGEqjY2WoWjxEmQPC+e/eCX9tghBFLXjtXdrLQUxhDRNnbPSO/S/OQPYm5XEUi0CSv0fO3ykcB
L4+iDmNpf3igXtCJRb8RoGrZtbIXzkwxkiP6V3OPEz0oNkkANwOkCUVGC+EQFcUdkn6kWVP7EwJ/
cvfqMv6g/mlLgf7tn+cVWInsQtxbIMKU6FjpXjNn1qstrXnZ35/dpgacQKlFEydhYL3GdLKkm6mJ
dUEvQ2lM/F1U5EKpRouRlNsT+vR8e9G0QwYQ/tISEd2mAA/fd1Lb+nl542VV3woh3xhBXqwcuedP
tkV9dY9/4fZD57ALgoB05xAcbMiB5Ce4FVo4+ktQ8h41wiAIPSEeVYtsghjFvI9R0mzncEF1tZPZ
2OFAjuHGSyUxpbtO9CkUOWdEW/zrOLqlnGyC8IgA25LgmGSV4VrhVJihikDIdaYS2gOEk2SspE3Y
aEr7EfjOSTJGZE7TAj+D5OAxgsWxT7Nnia/gfFp3CZnwYSSq5YnMaVFKeqc8bJoPV+opAnnt+0eN
1IW/TNsSc3TVGVQckOw6CPLRgLIv/iRficwUZQHYJtnFkTCAywtrWg7jfXfaNnyj0gbSm9b9Crbg
o584YxbBSAxvXEqrR/5yDNPzAn5IH9wPU9gnUGDXGzzrN+i7dAEOF7SogWdbDmmuYszk7juvO1FP
iSJVvxJy40sY0e4cDZ2iDWZlIM7+5IvtO6d2OHlkM3VtBoF6aZ/Cvnfd3Ar7p5vXyEa3e+0rdi6H
bWsconwUwmLExYLO7uxu42lnzNAIOZgEt7sstdoI08atXfPCc1OEXKuPLUULHLQ2QBFCAKuwO7Qq
UDC+ub6j+dNfiiRs2Rp2ekBAH33Y0yVh/6QJ74Kdqs/agTBVNFhHTYXM2ZOpbiA4vExwSqNSMMKC
dgrpchXQh4cMNCNRE6FhmeUDpNzngb5PfhhjcL72+5T+yDxBFf8fAueHToiZL25M2pSujDpRRGXs
PjaG0sJozxCUXyLBfGLvqQfFInDw9/aA8WR0+W6jYrYSa9CX9hHz6OarKz02dmC6T4Tl9+nBIf6M
aIgOr1yPjUGEpIH8KfHBqdVvswxAbhQj+8Bmd/LZ/iNCOZ//LE7KqETYHnrR0PMraIM18c1E2jS8
93aU/zZ1NO1p544nM56+3YCZUGrIsTuANjCA9tMrojk7h+nQW1GpKivDbajc0/CbBXUCw0ccJcA1
vM/pgqaATCK7IhwyQV9KM30MAUx+djEPN2N8g2PNRDO9Ioi8l+K5yz9pVq5AA6cZ6wR4qUJv24I+
1iy4MHAk5RBFSBw62XVK/VaxG8e5cmWedY8GzjfzzIBSS9OxqrYtQZUW99eTnFuNtnjN/e3FNfXA
hihe78fVte3qz06cyYDs0Bjc6bT73ZId9Xi5G8z1m+RfmYYttkMok/yC+WuKJKH6EXrUU9XRwkk4
LDxxxl8n7HajBWmeBIHgSzDFu9Vu7rXlP+4VvlFPCkPqNayoEsthkW3ErUwy0br5qvlxgDgtH8DD
/6Wr3NxIhoaccOBu387ey+JfOgIv80ZKXGaRFL6XC6BesJsiWRzApjYUGRjC5e2YvCO7n5kWSEwg
D03Z/3kU8c1Ot0bMSwa+1T23lLIVcVi4h1BgPtZTyiztYcCEVKufHIG2gtTRXNNdIyojfp9tp3VY
VLiG6eJqfJE86uee20/HigTNxMbPrbVuBoqtqDipfKoOSAgaA26uvseYm3uaHE1NhJIrggznzR1j
PoInXFpYTxqP/IEc8BJxO/pA24ZGnLH3CkzRhIH86xEXUeaOx+uyYfEUVneshsxoDAvpBjxPKEfN
JbYhm69+smo7lqRbBqnruI9zNETVcmLE2dogmstBhqSj4Wr9NlPtNQsLa0Kptso0g3IEkcuUCSab
hQT4WKsrxNufqitLyObLiG18RcB5C/s7CrmYlohfoeXYGT9PyBpYE+cTYPQHWTuYHO2bxOgUDssc
3QzNH2h6QtkpWm6vg/XxvIBD2x8QhbOiI60PxSbmDZKSGul1RlH2D5/X1FJBCFsGyV92nocxtLu9
ZuZqUDQpk1UbTl3v2jJCqjUBLiCXtihx5w4U0MQzhKNDySpPwsEdTAkclNCPCixaIVWn6rClvvnT
Mmj4JZXnQt8ena/aoiZo52uQD0eiO5D8cR8FQsfqwfscvudRY6oSC7fZCkw9VpOFb3QtRvR3z72K
mFyfq/VKSSN+5eSbyVbSvOoxQRBHVwpBtaM/qW61I5nvL3lGxP18ORLula3YS5HlBIlvCC9BTsoz
csGz2FWXl6HAMuZLSMs9zVVr9oVcmyeFJFQJ3xlo/Dn5DxZdEew8KLBdYf2sH8pcxR4SlXmtFK69
RYYjBqa5h+upjjofN8XIe1DX/CQm71Q7ZYyVyyZtsFbGuurpBcp0w37Mh0lBwekwRCF/jad2G0gZ
/df2k/zucq3QhjtCKxy0o/9w1P+Vw+aBtVOJLBYjCW74vn/L3od7DZlgxaiqOj4Hvb6URDnmRYYx
2jwwtDN0E+50sHrRyEFG8LSy1l88ytmt8Akl8UEENZeQLFUIwoXD430Bhe6PwwIztEIUIO/b5Ynp
H60/u0iTStxM45pT3s9NG/5JGbelCzJ0tBzLYEqvZn6KK0mmECIy6uJDJdiiK910j8JI6xIRjhXC
g4/GW8+Ku2l8C56GzqZQ9UrkWWxddV6sa+s/7T54dcse6kwnFvISVs9JkxE92p1RdVCXYNnvoGMU
Ivy5jNDctgSTKq13XFqjubAxS76QUfMnM60+jLnTgPoVXviBDnwTlDm8PONw2cJIc/MYE0qvjzwN
GQKqd57qC/gtBCg6bt0m8FE+2GIGW2Wlw+3OkOcwiAsjyA26xXOn1IGkHI2VFyx7iaPiWjM1JZer
ibuUSREvb4Z/7+a7BFFh2e9cKKleUpOZ/QyJfvPuVbsyA/5+J+N4663nS4mUb5VWd4/b/MWe9gKs
wWFet7l2pgzb4yCzkd26GpZs1uJ+ykYh4IFc3d6VZAP4VLlYBHfuVqPU15xLQrS/WDMW4boKq/aI
y7OO0eFM4o6jElD73bTAFEF2bl8XUbq16vz2fR+Vv8FePe3CrKRdpxUaQsUSZrFPOfpPCMKH7Jlg
FL2CloLZaWUZZAyAaC975dBYfdDOXYNJ8falYu1NkVz/yuvJsEIuNB9vJ3WQf1xy/enahVvVopqQ
pc2uO8frdHkDJ73hehXcreTQPr8BKB0IIcHuUBy8knKd8FDGGCBnEzK7GAGA6AnMPDLTxYFy/2jY
YQAKOtuT7q8cOJfiYeott8MnYNpci7e5DmNWiz5AwkGNukEUJyy2D7MWgsWB9PuMxSXoGqh3hqMC
bZVFaOOx/QceoqGTWlIi5WaaAU9CYIc21SiJhD6MswFGJ1GnShUbJbD+t7iiyKsg7FdXnHrvvi5a
jcXvuvXRyKoAvBNoP1zg1LtHuH1nOrB3CS1s0CcqTNHI5shV3d6wMc48n4jvgZSHqWctwcxznKsv
tBlvFbPpKcGOfR7g3o2Sgwt3yUMnmWmp+kUA2f9yAiy/4FLnbAPq9QLtTBbriTgNrNlNQsF93Jmv
mbPZiw20gLa3NMoVG/Ez6HL+glFmQoLiDqr5Icq7032fX1ZXov42D7dI/iwXE7yILhiod+W/dkYd
0XAXPvAdBdsHyRTy4FreRWx+m/ngWDRvsSRWp5Jk4Pj+YBWbrxRH+fqNV55ZXCghV3UgXXrZNxV+
tATqViVuizkrwT6rNoigLy55Lvi7k7HgFSxjbsaG4GhX1kXgHvZAF4Mi5WH2542mkfq2nAcmAfCN
ftO7kq2dqpRancbuJNYqW9ZI7vuoOBxQFXZ59ZJGTelL0tDxQBZtFEryoeNv/qgFlxMT63UnZEPt
QIr0KdqDJYcFOA+YMGaDQO6sc5EotSyCz5zr+14HgXlI/F5Pr1h7qJTvRt6jcG2RE1feu2Aaa+aE
QkU3adg0snSQ56Qwwc/BMr8u9iXDVDwmkCWt+s6G6RyoLsA3Oyz0pf2/ME5f+TIVzHePc2hgl48T
FMyOqxEhdGlBvhmf6GCVX7EDhgzXkHSGi+1XLQompZdUgOCvHJbyRgYQFtcmLmGuuiELZhwVyDsK
DRxlQ3iRginVZqqclgHdg4mAc+MlKlwrXkjY9CUUDyZpNMAV2CO6B7e+PYalGELW5u4Vxx5Wgu0w
Ss2fmQnayKyUQgo7wIHz97xpNJsDF0rfXYXXioSmNiy7i+rEfDQGf+AZK4OKO68oy6Hg3eXPMA2y
UXrXRS9XR2zx3bd1TaMU3tB9i+yHIwk+EAf+p78CDdo103wwcQkKEIokPanwprDKUcE8kYR27fuQ
U5RZxstsnpxZWr7ipNwHmr2v7YxZg8ljX8Poe2wzHURIyQ/RRpYs1LD9dRdeeeUB6PZo5fWIP/DS
WZuSttnjW3JylYJGap/dDFKR9gjGPgnvX+hQSeuYb43d2PfjlPXIcwyVdpGPITAC3JmKxXc/0Bqo
KhlDmFX5JoiBXUXR7I+1QDaJP+0/Lnam2mC0WdVRdYrgENk9hWkvEN8awioxIL2ydqovPvF4rN+f
zRLtyP6sORQv/YQECgXQCbLaGNRi2iGottsmCCrSYSoWmQ0BMYsG05y3E5eUBKv8GB5R+IebXxDe
7lJkjJVV5ZgfpQBXkzAqN6tEhOlaZzOEOZVYNnW1WPup6NsxZoqESoa8AdmwVWDksDWMXo4ZCjfk
tTG6B/uqbAfKs3EWRMKJdLwXXbwN0+IMRZkrmw+zcspLCh0VcilY2NlsYejW9sVETmI+9GxyHWIx
tC2gP85vt0rCG1BjFuQ8HC2ooccyKTmKZ7d+zqr+OCNDeAZ0g/WRGVdug6hxgSo713mdbZidljYn
W5MAiBvWvgmymgQSlM1NeEmHqZbOX4J235wtiycxs5S6RA2RU2gdB1hNERGlWycwuxy7kqf/d5rx
6+mDV1cLaMRBSa+2utNOESKS1SktkVBPrBiKKMgcmletdaH5xF1nr9iFFVUkBK/ctWY2S+C+0gOx
5OJkIknNuq6yoIW261IfZaa4rJWehwkG7JVuNZYGDCqX1NR1y1Q7wP0F4lZbt37X0KYLgpTE/Jhs
JSqa2Pv2PHEkrHv+WGCaBKBUxzQamB+QOKT97rDe4SFvpCQpT2o6za3RV69gnv/Mdu67DfIwp97Q
m8/Qc2r9FYFA/burKPuSifYwNper32YE9yIDdugRZc1gql+E+h2IER8NfVeC0yQQmPgMfGoiAlS+
Qi71xFwPQSoMrUMgBM596vMMMyHmyR6VnMOGdcDuXtfUGMWzzyYZgYHXHHsq396shegi3hLpdrS5
tS8VNYYf7LclTN5I38PZXUuh118l/baSBrePRlSBVLSDI0RU0EWolWAwbEJL4IFERQziMcEaNFfh
XYfA1FFUh+A45xE3WdQMynAJv1aDbUeZYZgb6dpcD9oAsDQBWhwcRHJqw16eAoKuis56pB3S2sKg
/nc4tq6iTepfRpl02RIyisgmAcJApWc7yuilqYBTRVu/YzDiEbGokzXMU8LHLA/YqkjHOf+z3mOp
Gxx3leXTUayBHD+kJmQhBg5ETeQtADCyqYUyR6Re08GJ4d5RJp9BHGmajpomFd4HB4yrWl+5tV4D
vV0LAD2wQmgFv9WvaY/BNRy3xfT4mFkyTckLDG0SZeUO0dmZ5G4/Di9P3w2rsEs7xP0YkBYvdOpK
nCx1zYRubIS6tJBSwzsuVU0571jriR/HahYhe3GkFOSqdqnIv8S3af3L4a6bvrfb62JbZ8KF2CRi
kqmVXfsUFqKjS1XcCwHsZ2lPnSjwfJe9FfmxNKh2LVTN7T8QiQNeRiuLC0GFw4EAsZLIaktbukZt
L1lwiX//GOT/YuJVCgbYuqUT/BKLyl1NokJuMI+KIweJ9cH47USuMmvW9stnSJPLdZn4yDp3KjdD
idnMFJJPJaQLsqTUxBG7jLBhA55/g10tGARqHiS4DIJXr1YJUePXRujN74UPefzRVlB7k0DAMO3z
/1sV7RyTqnDk3oLZZPKDrVx1kJbZaSu6Bt4S3QRbfokMnjeiQ3qBJpj8dfbJ+xBQp7EqSIp4B3rd
K15R0S7GP7aSc1I+AvxRbeGGvDTU42mf4JhGQdg+AvccaVluHF67QFqd9TIrKm83JVLaRz04h8J1
zBHsE3rhSFro8r14cfbk2RzWMvsvBPGOfGpY1LngmeTzFp3+Mke6PQL/zC6HgIq0sXSXPRuKN4ha
85/PomXf4TVXRGdvC1CMUd1X7PZUtDkMaOgsFroJex2W3fHwU1SIYLyF9Gw+HD5HLSyyXxH582l3
LnqhFPHWi65Vf8VF6H5J5z5jgOKyU9g+YlrvEimhh4frOlTZV1dwGsx+sDBugwtDrxUkYgyLlxfQ
XJYnWarmxnXmpcYODuK0wuLZKQZ5RPZOmTNii+CHpGXd60nL6P37gG6k11Qa36Ep/gS9xHCNY6rj
3mep3DCIpNDLPysJK7Mb777/qo69FVOcLAFatSIHI3NPit8O2Coq5dXOsYDf4ZdoeczioMUf02DW
Idt7vQVrCaRxULxyfE4qnIW4DTTTVmERLnI6LwARo4g+Gm44GTCiYMVpq+vSCtMY8E1BTNbzcptE
iM6Umng62/Xhc5tgOE+sihwyvTIxFSxyw2QZJNnYGivAP+S2IXNj8OZsPfcATwJ23R+/Z8vUSC+I
i2BYswmP4N5z6R4iq2pQYZT7OY1070U3NFm1CC1YLZpERtx8UP2w8dcQtQGKxUekvsJJlCtrGSQY
623UbXdxLr3qswIBtyMom1cpmYnMyu6yBVv+DP2Fa5FFMnRyioAi58eei837cEkcTSS5hvSDRO6A
rdC2CxmEhZE92AtPGocEdIIdqUjzZtIs/qqCnmQynhBiMBJGu8taxqjEDdsL/GgHU+wPv04/4XYI
zj9KtNNgMVWULCHsXx3iwrFae3ehkbE7CxFfaTuqkr1QpTmtaVkeE8M+HRNASqEwYg3rVfvy3WDi
l4G3ewjnG8OtFJ45V3OTxlKFb2GjTqdQfkwDXQ4zKzhniqiYbl5nkNVfIA1OB5QstqHYZFkg1PnO
DbN6Hfl477JN9Ewk1+VwpQousAURK3caEl1ZF+1IT+Lae4go3Oo7heLhS4cI2X+NrY+F/emyHiwM
Me1knPH3WTDsiCOpEbHHd0RC0buUr/RmaCrrvwloHRjKUypqssn8FoZV1CXxyyOTl12xvDw/zh28
LkAQ0knDDj78+X19EKDMLdstFDO1yvJNTFd0FIprRIs4EeWJjWB/dxxdTp/pr47HZ1VvwziM0Stg
fOgOWXu1poi7KOx9TXv437tVnr0BQaZMss4Y6JEIlTloM50Px0npyc7mAP4p/v6Juc1ZmdIIlbLD
8TfyRZTSbbwHwP+WpsP+RsB0nlp4gRXZ8iZVK1P/fsH+HBDZZDLxffZSqeoeCvOjS9FbSakLt1ad
IaLSP3Tyhj55xljgg82G503ovJ6sMVIr5PHQvnqQXcsWD129nN+WHkWuD/XMB9HWb6SpC5ghCtiA
bG2M/VrqW+Iec2gx1W7O+zzhjzD5zbs+r6ERiNkuYWvyAqLqhlFHyrLmlgvCMPmerqkVuMmm25Cx
EFMjtaU00dtgS41RZLH16ewgI+IEPCQjbUbXg0x53PeT6Pxgr0wmk0rwAxv+K+oustfVN10TsKd+
HVgmNV8ry6EjO7xSLhdt6/lUDP7Y2Gwb7xKGppwcAophIatI0dC0lsfLVuRUHPwE3veUEbCoU3Hj
jY0S21+mX8yyxtSShjlaaOW8iVYYOVaR7NQYzet1nrUT+5900A9JRTpJqoNYcUVBMzig8xpoQ8Dd
SDmoo8ApglQLYYdW8x/qKme2DzzVJSSIQToWeGzvehoKiQ0gn6kYgTrmcTreMb+5QSNMVpF2IhsM
F65Lx3DODkKKalFPMyEyE93wpu1G43vrBrSPBcvapkPfe70YbCgsVmV99LluF3O1LqnqeZrgiDRv
aQqcKAXONUUTNeZgJ372rjXhLCIre56WWbbbXKXjf7XY64gsE5DlwC6tCMzB556XNCkGfH4ZxiOR
7TlXOZqR1unTq44Zw223433arH6texcN/Z9VVvMcubUmmC7U0Lxmy7ueEHhOI563QeaPt7VBasmS
5WyPXe29ojb6W1138XTPlKsBxQE5xyAqNEdGQ5WZcaj7DXS7aJG16f+J2uudl9CVI+QTReMLtCuP
UcKC/V7IMTsqeo0iKXRKFXho9rsS/OQIlWdEOYjyApOdUvBNYnVhEySX/LeHC7CDUl4LDu7a5n4E
+TZkICoFixSG0fpHFATkfzuuHDi9DXhdyx0l+3919GBiU/4O7pL5kQIPKU64mmROYrkKbV7qpwZx
yYW0fuX3BwCnZ3wLLfw2aXIt83FIvWNYlueEpBelOM7tw1lylD3g49jOnKcGxFoRbmQyGiNfRn/J
VjpM9Y71H2v0yGKf5N4g982KZ8sig0RIwAQ8xbfEKSOrHJeNXh8yEsGAHYpyvXCye1GUr2AqGayO
8thfk/6uR3LDfXxlM3EUfcyoy9hDVlmaaANJHJc3shUmN2ZlNxl62gFONQWvrKsw0o8Nm6Y22Dge
+q1re1ivt3GsSVCWTLbHlpgE67gOi7A19j3PcZAUrQAbCr6z28Y8qOMelvsIZ8uDESQWwUh8CY9y
STAq1ksncIb8nDODC9SNLkpI1H2VtRxkmcJ9M1XlwJkCPKBtXpIor7C136zsud5FbWU/57VY7Hxg
aXyYPJHeqBr2Nc6KqaN1areJ98w+gdkLzA5t1wKyDKXnLppNeZkYkF66hjLc9o4Y2+oBVq23WIYb
wO3545vWP5KQDzYjDFsAqF61z5WI8T4kfSC/Y9BcsdpGAIkH76YLYELPZqlFv+F9lbQne76xjC2A
90EZRF2o1kUmqvdePxgJ1mvZBj7j4ShJNFRx5M3UcbdIbBcAs2H1DtsD+PrCKg1oWWmfU0sUN7ZG
ME+nuqK23T4kVuQ793UjmPFWj2Jz+W+OQdKTosT1HX7jdGzwc91uVTk4YckoHYRiaJSOcXwpMNi7
Jy5xNCUyq6fu/6r10YFVNL/UaodqmJeKJa5ZZ6hZP3xHT1UD1Fn9cMr6UCd15YwxDidkJpJF3V5m
HKsXcnnN8L6nn5Snr+1nCGwpMZ0C73ITAUtN53eJnjRRQl2GeR7xcNDq4V+q+RXQRjCIyGd+/uK2
X5KYvQZdQ78fgORV3GVB9Ui7JZ4Vn97hL8M10NwJmd95A+jQVGHD7qkve7nNNaXIa295WPhARh2y
HC6bNHKS813JXjIfv3tsufRzTQk5Gn+F1tMNvXvj8UdzyAC046UaqGGpfzy5J0xev0l1c/pp37pZ
agNdawnJR32PJ9HcF/+TGDzSuOAir+iavRmfanG3TzMovdGrOKRuLafX9J068235T3xYvnuMsNkR
OWAM8YHUNIPpX6JkeeBygafj7ah9INRNeFtcSfHkrWz8rbBx8madQ9RRrqFscbDYS9RDhRzt8Hg3
mn2TLUzIc7B/gHKRc4NEJzXCZusURR165RZeAuEvTR/SnULCmjSbpbOXeRGcYyCkcVV8OnxuuYRK
BPeQDr834f4mq8uH6YwGzvcDBANP8nK6AcpYo2zQ9QLw7vklCAyCapx4vwVzD7vrkjTqmf1KzEHK
L5vtuwqKmF9suM2WVw/8VWjdyP6nBvX7xz5vAoeNtulLqcGBhxI3tqcRgMeBHqaehqHu93M5iF0/
z6IPvCfF1l8N0/U+w8incI8fW8NFlGCMqwm7YOHRyVCGJz5e6oI2DxvA2cgru+p/u7/EJbtx3E4R
WK4fwQAsBtops1r3EFxmnXD0Ycg4E5J+DDl4vK0R/cGaeSHC5OQvdJzTZ8ETKsvYL7kotgNID/7v
uj8v1C+tKucwvlqvG7nf0arifBKihwZChc+jQFJOFk2atb9/mWqUn4h5Ldq/2ZPs5Pe2itL/Y3vN
IhuAMN5GAuJ6x4vkHtLS0/kyuTi4DTYW1NlBrYRRCHLYPfgNr8TWqtrWHReS609QeRjldFeb2xek
TLgOI5I9wVoVxC56aNhOU7hPxucnzZgYLvp8iX0wbR/zac43ZIjNXPUvpiiho5xBsFP756p/reBD
X2gVIXVZUtGzuteatZ31BOs9T4/WVYs7/ymHQp8vA85IY/g60PLDJXbFsMnTgogJptONJhsYbaMy
8fc9NUpcInI8iT/158HZFtoiV1COAEW7+x2RUANen9NnkoYDA/0G3wv2Bfe+P2acLNSz2nx+vSY8
qGDtVdxvQ412eVkq3GnkpLpAlv7pdQS6R7YwF92WDQZJQ/vAp+qnm+tMqUnd25I9FJB85sungEDl
YF3fuqEFOzfEdLnVjZDaTqLpNSNmhOYVCUsQwwXEnp4F/xya4Il7bexf1PCVyNxGPMSu1CQm+Zv6
oWfKj/hEKBl0f7lun3pb9w1VSdOysbgQgI6X3Q+SFarHOAIYHd6g3YOkQ/LD2zqvwIWL4E50IZWK
Oz7vW5SRrRV59KAk38nNNFoGZogJHYjh19dilb/7Y2XHaFouZ9gT/pL39K9030rpN0VQIKcEKN+a
0uIRYAf8uSVZQfQJoKsvFQCZdMSFmN2k5Pxh8yquh3Mg1Za3ogg8xF5jpVi519/uIIKcJinMlAlK
hYi1xsHGxNRAbmQr1PhUnI/68y7oXU0KuSJ+xk4o348M8QWZxXOAqgpN6SRjA4GEJ2q8jF3hkoSi
nP8Dk0cnVejy6N0xzVD/HeCGfWM40bt6+Zj90s8r8vLGGjSU7dAS+YQuG8KMyYrEJ+AIC1MDGnLH
Kj68AMA5zKAS1YxXUx2id+0Ce3VWxbjKbVJLR3I7DFlX9I99dw2W8Ij/PYTjRu6fl6J1RIKpzyEJ
8w2EM7PuMtkdiN9LXVVJauJPIcl2EX6FgUpwF8lLSUajLwdgk0iaCe2hDJAnMgy7HE0fJc4/r93p
1k31SjCv/yPDzYASfNOyNwFA+cAUoe87NK8AOiJq+K2rbtoyO8jozIY4WzVeLx+0Qpwb/QwTDRz8
hBOjOqjBE+34ayJunpLlTqyzyxp68IQmbUAJ2Z0tNfVb8JJo0dzpFgkHe4H5XS1Kefe8GOTYGeyu
Op4Rsau2gseMcmPUXHQgmP5T4D95WDtuYdNH/pFG0dakKOwOjSGeBI/nD/p/MKIfZEXMsRBy9Bzv
e6CxElzVxokOkcFmKl8owkAKPMZZHeB8obSFo74WjqTikl5hv9ncXycOT+qNJsLgRb2RP8WiWXKM
cD4Be6FoEYyIuCNfl8uI482rU/8XpmhL9wCmNelucl/qD/HEHmGb+pAIEO1o4fa1VMA0rgJycFQZ
JVXfOpMoww+LV/qnGzah7u2EN/zcgvVpYrVT8nyR28VDNprhOPWhRqfptFZAd4D0h+yH7Tc7WDdZ
agJ4uJpvhKnSaLeoCoadhgYSSRPv41Ak5qpSYm9wt8mI1fUsS3X05rxAXg9A4eInbt2xjCvu3Fjp
fZy7nAV8dJGLX3UkGf3VFvVbfGUN1Qnei6x89dC8vc5oCTGpA5I7snopkPpglzxGZuwWwxIQ7M+1
P2G+3SWy9jgaWwIsXCb+doLafvqj8NqcNn6oyL+c9StAMEjgbuDOQXXenvVm3cs1Fk81UrG20Fmj
tIf0Je9zVRvNcA35WE/pf8fYhUvVcfXtmMq7ek3P/Z3LZ97KH7BwhW/MwFb5dFEOyKPY+Q2RnD2h
Ro13zM9rrOjD46dztjLwZl28T9iK24O0uIRcx0q3vhzM5v1eDPbJcA1bhUIWF9INiZMnuMoXPKao
bbzJBspKxyby+LveQTvRb8k5mOOT34l/eTRG0kYFLmfE1qq6p9MBqPHHcTbt9P/Q4HsXV++x68KD
LrxDVsE4DR3tx1pGWbK/O8/j1N+Do9urQOeknbx4zFqzVOT0FAQIIAfioDL+EqeWSQE+yJ3SQVnG
MphuRY/9F5ks2Xtq3m5rc8Pn/K3WAa1PBCS05+SfW37t0wtzrRqjqzp0nHbhf5sN4CWzdpVEU+ua
CDb3ILuw4B01vTAHd9nHkMkEbRPGiPg++C6r+GTcK+DPo5OxGKR3XYxAsTirlxy5t+i1+VuP799c
cr/5Mi1DtNaakJ+6w8X6nEGAxjkrq21q36S7Bn5Nb9Xs5DdUGEtQkWSeEF2HDLEHhw6OFUUgIrcA
aKfMnJKihd+WVe6iz+rtYJ6GqEZNEI41feQK9DM6OQHrYShZbYign9DgewzLwBIXKIf9zWCCmS87
Qcv+x3Ww5SVTQPXZgDtGZCRsX+eUURU9+Fjfuywhkw6u6aUL1pdoD+YUEuO3DvKhmiPBpeOPim4v
E8SUVgKWnONVIWDmlCvnJI6lGIm1Jw1Ba2aOEKqIIBKLtD83bLJ9wDtzmqa3Gj90Pxu0Vt0u0TJQ
75x8w8YKEk+iol4WSUaR2iMzFdf4JdmVfwXOzT3Ji7jaRAL48PSBzKjBXIra8pyciD3BKrv7AebN
uADkqlTxeWDQC0RKp4/UuY/iKe4rDBA7BbTe4/z/CBTGWcERQBYPsFCZ0wSeKMvcQVPys0AbCJGF
7HTjXjSa3GDd5HVagfGonbga4OSHBlsOnak0/Z4yBQURBeNG30m0ONpAW0XMtMS7EKpOn9zcVb6t
rjqxAERYY1zIdv2f2H70msGg6ybAPFBTXkBic9aQIZoZlcuKi8FJBJibjZTmtjZurGmYBDBud+nh
SrW55qJtVP6LWpWHhvIX3CQOhcQlI8tkxh5e36dR+s9Pg87zC98WHhukJfaDjWn2MABm4mEUC6Xa
AH52KsI697P1R7CJm/TcpNOptnXemSYjtdamaigz8tBzKLd73odolKAKlvfg8G+aWljokWtOMqoV
3t5nIOBTBMTiJuKZXrJ5eHqWOdJie022kTwTUNO3mUk+VWZF/Tvyp3Pi7dGTX20kZ5V3CnKy8oQa
9ouGbaMxCWpC9Jsv3mpHbQfEAEaf97CEVkpYwN/Ccx0Bg8ECr76W2QdwyvHwG89q6YExBhCp4il7
fxI41Dz5dlFpapeDl7ssJxgizS2KeysMQ80MxzeAqSE+ao1NB0VLoSEJK/o7SY5LHIzO568/CNoy
xTecS3+DzSRLyueltf5LN3rpd0H9tCGigJ/dy9rSuguqb1FKCp55V1t9VEwpnfaFo20BrPIUW3XV
AhK62MNgIVijf3KJtUmIsOMAC6K6ZLlWT9hqvjUlxVxUphbRomker05KPUsMfMaki+wXIbgKa5tM
ruNXQXblzo9U5nZU2mNAiiw7qMRSElTHxLd/W/6jBU0Fawr35C2vhHsCiHjg8FHR+aNQFnkIP9Ce
+R2j3N2GizhdpSlenVqyCp/HiRR6SDhiLCURcFFiUTdGIv+YP5xqI862PgHYVEfG5NuDFo3oUUH8
zq7s7uqnbAairpY74Hoot/K1Gl6NLldeqsZ+arPqdNk6FM59WNiOHuE9MZrDKLSfjuh6MTRn4C0Z
lg4cnCmqyVXSp3+VaoEOwr69/hdyphfzvQPumgObu8yIkmmtDQl8hl8Xxl1QGGMmyspOP/wcGpWX
gpGyB2mSCOsChD4nVK2uK44CBO1QVzFBt2klXmHpoeFOMc9k+YhZSVw+sosG2XsDFRAkYcANbZUJ
ODu9WfCX7Z2Jjv5mli/DoMismR/wV0NgoC7tQmNmDr+Qm9baa76gNA3xmdm7oAvKyo8kwHoarUmp
cHg/tS9AEnk7/du7iNbfRQ63chPjcEj/S6XLeJF5MHRhr7MHiWh61pD9Y2rJwq4oSjRcr6zxq8oo
dNaA3JQVG4ZLLkDjhuMyCo/Syv4UgL2TWa6HXuRieB9IkdqnDsQo2uWBiWFSRSp+W7orHOZ5Hg09
s0E8rtE7ay3u8IhxVrMx6ruT2E4sqzJP40CuPabxMmGNPh0Xv0blLu3YBsjz7jA84exmaXjvDJ96
If+mbsMujESyjL2UYpLkd4hP2HT3NF42xKf3X2D/zLtDtuSkGLYXs5c4HpCNYniSAnZocm8sAGKc
hw270F4MoJb3Q0cb8Ek+GtevcFy0QkAQy1l4KsZSb7xp0VQr6YPdFNm4awEohCBhJXz9GuRIqjN7
VSRuzs13X232fJ0FXAJVohrthQH8M2oIyCpI4PrWpY3JHGQCoPEMm0iWLYuuXrNWH9UZkprcAvBj
kfDT1gE4sOSV7e+rcgT4UekagJhWe5INTms5kTJJGFMesVxBJ4f6o8rM4cerHbBcCbssxN/h0tfd
clQidas/aRVYVooWkE+I8Vz34CqKc9NktU8eZde7tjFqZnwdjE5E5nBOZQ8oWJ8X5LLMO9OLsLCI
ntbWYQPqXd/DZxMZetk7LXPtnIMfcBI3UT8wpMsiKkJhob62ESrtUO5VQXpRnsGRYLnx4A+glvTM
VgwHSVkN3/o0x7YInPUnSz5dvAstaleAymEYMw5llDhkLsjAon2JJPt2q2oDfv27QlKK0RxVlg52
CZPkftHxK/cNBpCQBWbHX0a57aFQlmifey88HqKIfLM9ori5/Ca+dEAyBYD3c9pvWHmSE5Emo6ov
5+I4FKythYlPtJ54z2EC9Xlsat4UFQan4bQIMdZ2z4H2JJZ1RcxYPYPVA4To0b5FUyDVTlOLZmZc
IryybTMkyuzGX5QJug2SWf7EAqbSdnhaySvRj7G5Eq+0drXRwFaTg5I93UycuOMwGezsYFbkV9lg
NPo+fYS/ca++pT+u79l1pyMxYaIGqYQLqXhFHiDqrD4EeME7RqLph1KRdBv0XYbcWXidEh6v6bUL
4QJJcmOjD5yZ3YM1BP83RGcfaAuVGjJpaT1hva5jROlT5FuxhBm63rcIYEVWIzFMv0anXgQv5Gn4
8iOssMIzPeETMbDbcvYenfhZ7qqCPqvi/fN6xfUFrOLVGCImb6n857UJnlAGAIZu16J7QtS6BWoP
1fiHzgzNT9Sd1sPthvJwI3YZxtCGeRqAt5CccY0bOO9soWfTno1v287YkNQqsOhzdEA6N7b3nTKE
FCfQi4XhwDS7h+wAk2mogwHPkq24Z9Xkzo+zmGxhmYLzqSVU5EnxyVwQ25MnbTln2wjso59g0kql
7hSBB/Tsn+yI2afCpyJkhhGgxHDH9UPZvKeHzKKOgtIHLzQRBF4Haw0+bKwW+sGZxOII+6BDV1+a
hxm2nB7cZSUjELI12ZqoVVTrc6DFAqojcuNMBY+3EF923+liR7+go611fu7hZmdRwkpKyNDqPMWj
p3o9n0s09+cBeke4y44W3SLgVChVfpc+kaxXXA6KjS+S/XmVHPndEkw6wH4N9N2tS/+U/y0usoLj
GysmIOb0ZDyc/xSit84MTe0qPAZqeqMGMGptQniKzz3XEpsMa7meGuJ35ogrq8cPNvqzg8uTzkTg
ehiepgh1b5+rp5NPgE926CpAbczl+hD1eYRiX9K1oPGa+lgMW/m851YL50vskwSZSiUDqJLzSpYp
quu3yw/bOO1HAZQrJ9iJ9uayNv1WWpch6Y3ihzMSWg7Q+r/Hjq52Dv6dHcGsIPOp+37lANz2IrN7
jqz3OXddNV7ZMWioupfP+myC4jZTjBPplxjmWTGk9KLNMFi0X5MtIssrnUlOBzJgeT0VRdBFxijO
IZOvRuYBFy/io3VykfKw3pT3N+v8YCXAxUcaY7TyuFmj+jqVWTe8hQy0H+RzCKnOffGAWFYk7kvL
jtpe7fs4dNON+y6SkdllH43PyULqMnEDLmTPhVZuJRs0cE9jtQaa9doHPlefdIYcY6qKBcoo/teN
xNo7sp6R47gdWXl/luvs8nna1IrflX1xMB2zHa661aYs+uFl/S2E5qGAlzDGPCUBWEcu0GAt1kLj
l4h9LyY2AaEPzMGKsDPcmGaDNtcRKL8rGFU7XP22y3IQIBklpXLtemP9skiWu66LxbNmNZP1x0Cm
EbKgp8FNrlRZrVTZ2CGhbSGFOjE4f9HBIHi8Fti2jWZHTuxQ2qJGOU+q/bG381Dj8nEHWf5jQI8r
aIxZH0XCjYP0aVbTWzS2UmOuF6yQxYQlq5154DhsuG05u37GiTv5YI4orw06+Q0LQd5Fp8UyxDE9
nrBr0xIiVq76ChmE9McDq+rrL+dW1pMymJ5t/OGdg2RRocHKhwOEl7PxtNGTOf73tvaOnH67HA4p
koOyxUFtRArC8A9H+R8O1IRP9X/OgUASIBeeqYBk5wzQ+QNeeFm3LH0I09MGGqNtDNQFJ8Sdy+9Z
utL0dpJeQabnI2+6nh1EfhYLTd5rTRIzXHzOYqMKwcVOZRteZ+zUixyBODe0hj31yK081WtIC6B4
sad86PhZfXBkfCYPKbo0J+sKwNnx4QVi3FdQoWHHt6TcGxfp5nsbRVAqxReNWbOuCp6ujBqzZUB5
/wZfSvcK0t/l0523e0JVWW6yAuzBe4Q/yT0kzyM2tFaWd9bY5ZUNvfdrK7zPaHQCqo2Vl2Rwy/E6
C21KRofKqDEu+pRxBoO4e8zeosrYy4MPRZSWbFRqSCnM0ahOLEIdgEPI5qgeEORVMrHYpgGfpgzA
wuJ0HFABGyugCQ/ENFXvIFzfsLDmCj4TGOZ84cRogw8/tR8Qiq2TWA5kC+G5QUpIhv2Cb7gwPxZa
iTidEQxljimh6JhsI03huHtzThl+F05qOuVDfh3rLUOfEiy4JUda9RKJg9X2aMJK2DqbqaPbdNDz
bUZsJHlM++LpSxSDmum/pCq9EVgvdBhVY2RzX6RxftXDUGp23pU50tqXOhyEwImDtG+LwWYCbUAG
WfCo1/uNLjwxMcTF0rZP4iN1go2njsFBtzgHMho3plJ87Q2uHDdOxzJl9AZx1tYRfYCrpH3aRbWG
fqNB4fXhO+5cvzThBY/njI4rJuulN9ITYwmV4ByqZ8WYm8W6EUrEdx6x1zquZ4E/S8/fMAed4fw5
JejZEqU60ekaspcY8XHhMGmc6w1LLYG4W6WLdy0k7jn/ATwCtDCgQOuvmG3u0hb2/X/8kQZwqI5+
RaJcwX1d5T+2kZ6ivT6NFEZUBpz8R4aei2KCWqoxKq9a7OwLrBfqkgHUuG8hPEg/Kmynp6hobiii
waclm2v6GmnwSgg+IK9zkjy1gj8hKtg3I8PwLIir+SEn2glm6sE9NkvcbBweeXizm0/5UIni7yE/
V1tpCRLIrZ1cfZ+GyGTHiRq4RJNab2IpJAKkMtby20v+K4EsQc0quuZnrhspJV42B927NuIYLd7N
yTNWcMAQ89PGtW1F3Lc+A97nfQ2VtDN419yVeg4ogs/zqehEG6eenrwBkilPb5zl+jdVevlI2GNm
yoyHCt/prnyD8qfRKnc1Bw+AkLU/4gzKs8ol2v/XJzvvsvWWkN3L2GNhqyxT6UaO5rRif0EpY4UC
tD8eNJNBsV73+1MhaT3+Z3Wk0D1t9c/g7a7wdtMhyrzgL+ZaCVNkZaj1OButpelQuk6wQdgfxb9g
L5jTQaQct7hsqXKLap/iJCaKfETmPUkP4KFNDC0CT6ozZowHH1aNo2+XBnyOhj/FURzFHlLphFOk
kjdU6A5Zj3keNG/0/d/dHY/2Y+RqO19L9uW3BzkftroI+BVNrDSyPFkPeIYm6RQHYN7kgcncG3TY
ZDitA1sHIb8fbW1cl7y8escTIHNtjVfvn9kUJ5FGCDWVQ22PtCp/95/k2xbfVhzD7y/DQ91rlTwy
BZbfvR9E+JQdKHIQs6qHBZ25vL57h2BQ0uGwts4xxleSkvOjonAr2dKtqF8S6mDMEKzgs5v+kvXv
3ui1oYc5HOsx4Gw1gokZFE7fB8tR3NLdFlNoB7u9HYUUXPK3JMcorPWRizOWrT5WdW5Fha9E5gqr
igDOsVnKxFGtLF6Mz38xZRUOATYRtwcZeJ6jCTVCT8zyKy1R0NuxOMV+A7AqeYQCJEFvFj4DCY39
Mj3SHNGTkrz/mwRKxi9VRmRWX9EGX8E907f4sSdw67mns5S+kF8tcbx1526fTIjji48SrM306ExE
u/FGPJnmhgn6ZZ/KVHYzPuFspmK1T3iq5SbUXNNsYe6heAgOHUs2kKR+E0JrJWxTlk9xwDp/UxnN
oeauOAD48/tKckheX8p5iRCIiH3T7Zbuce/psacdKkrpXmHGcUQzZqxCqYDCGlhBhMnyC1EjIRUS
7MlqgxGpUt20RMmSXk+LKJ2VAnJna5CH0nqb+iefYHyw8fa/xkho7M6kPZr8bperdFNHAM7xTG9d
9d7d6EP/dD1fUtlwKhx5hPd+da01qCmrfBypGw459gkgFWRIyrmYCLalXHDo+DKGudfc/VQQwmbY
pdrrlcVKxfrmd+XUd0lA4f8r9gd1u6TXG9nKB8MQ8BE3PKMiqk50j5cLLNmp44j4Bqgkf6DSkOph
I+8G13PtPpkkqoGWjXYgMYhbwYtIsApspHBQ0Vg8F5LbKZeS8CSSQoFuKYQDIjfTBMmsvS7g6kDE
tdR5ct0sEmoYo521+HWR02aphMKD9DnBr2Mj1Z1cdlimsVZmfgZ/luM4qC3mPySbxeAv6lYUr/ti
Db4N/YNB5VGdUrtzWgzD956gyyIBU9BsWElIE1fV7MFCzO0Ydaj9P4xvbTa5PhFqoDJ3+htKRpX5
ZqUr53dtJo01IiEsFUP+iOG2T0Il88qxbCq3iiEgTH3VoHe2nbFa94RRTUSyRiL0bDXbP+r3SpXP
fMit/hANk2pR91CavAovv8P4XmkP+MmQFlnQChPPQW98OkTsi8YgngQ6MOfjNq6qIPwQP3k3+dRi
Y0GpjTrpQbTBVsPFBXJ/HCxtLrVbjmaJ2fXJzc2Egq9LACLl00mqNtcmclHUAZtaYfM0t4KB66gf
f0xyLdlnOuyrfqnJJQnlfKGHRe4ETyK134ybIk5ZyqsVETq/zZZBaFYJa/uYOw3Ub/TapzvKqsFw
w7sZNafzoZI7KwrZ0ZHfng6XO7kA/x9hmWzuI872pacJZPKpWQJBTYhJ+7TbfLEYCeIRKrcxrUHu
LtN59qHn3PqVI5ahsh+5yFjNyyx3/Tw0ivZCy9MBQgSQRUOaFw7zYWOociEuTLXKYcprfHKA2mmJ
OsiBkhQjb4UJ42+HkfyNELXvP1/DERAUmHhlYItNIDdoMPSABl68hrLcu/mTNtZvZyWfmqfWGpQK
OaQoekcAzhGXuoqz0EZCwSjN32i85MaOE36jonfugUjRu6gmkqnUKpXHkwRNXEe8suCbA2L9ycvH
/OTHiRdtSsmPEiGdPn8VeybydcTonJwrT01fqwgdruwDBcR5v3Vdajk3SobNeprlA573KeQRJKgx
URA62a/1gBj8HTYh1v1wd6KOB2F0Nff8ee4jbQM1y0UANPyW7CnAgf7rZ+VC7Sp8yYr4c1bn8Z6R
Cl1/5QMwsEDluAUVoyeTGmFplXZjDv1I8IDE0wj/gqGGMfZLsuy5fQLoNPayvUu0BJCexwuqZVQE
CJZIQyzw9mWIJ1lVBJn7BwHcCF1YYHNxVKo1+9hJdsbL+K3RhrSHj+bmJoDXOVRiPArXg3pkswcX
iP4XizO/RK/iMX79jokgn3/h59tUw+pwXplyxm9vWZuGqRE95GRRYw0lvcBaXO1xyisiYgQtvcsc
FywQOhDuijvqrTHiCYQEAzIqAUnBDX+jUsdk+U99iOqZRuoJJ/cQBSNRYZatKU3owEPbYPxdp+50
HskUdGzkhX2JEQY8JLuaz+ZIFzkIUJ82I8+ZpHr+uk33JQHMTMP4R+nrtebESdFAZLQiG5FffbHj
ZfJk9r+ATrYdIu+DogedDiH1YTi5DXmLEjEbQ0XGEId0isyJfpCe0bF3zIr46coEx+l/azQZDFpl
ersPGABa/VhxWhaESuy1hMEGmgi49B7j1A92rWKhCXiyHSphvnMbPt0YG66O+zDt8I2ysBB1kxDI
J3N/wdiUGDldgJngWI21TnsERqncTCst2VWL0VkmQF29n17V9ESclnSDKwJmCXiGERlqAzl18U4T
ntViyahwBIDhqLxzHldkka5objvHROJ290gLdowx757GPYMlf3lFZch9aS/4BLrAeMke0895+Twm
YeHknwFDgPGnzb2DxuJMaiTCbdSGRdztsVMK5FLIsZhwSo2bu8ZVjaTu9u/pkha52e/ZO8T6QaNS
sPdvGtDSG6O+bO/i1bll0KjCxaldEi75Wwuw8nfBPR7VI3Ghup/0zwjLJ2YakzaGYaSBVKZ/FUx0
Q1jGf9ZTvypeELOsjVURFE5JFcjL1g2KMsZ2/FoZZE9Y+5l5NH5lejpuCV5uNJ2g0SOayflcMSJK
fAZCl9aPEG9KHt/eQB4FtvYvwlhtk11y9tAPGKcYis0ZIDE7oManxq/v7MjNDtWuxUgQvFz1d9pe
Hup4nDbGxYE5UKNnoFbuUdhIUMyepwjwO2M6lpFw59Kd29cEJ91LgtTFTm6xt524GXMWZLABtQct
4U3eU07gPM5sq9AJ6W2e3JBM7s5+cVcu1cS1f3olSuywd8StIgQDX5W4qdfbdbBZu2qUW4ODt2jc
0qShgPE+L1lXiBZY0MqFcSHCSBtjg+LT2b7dFK8Hpp/JRPsTgNLmrANF7S424CEGsL/fZb28iI9a
yaLvRvMBBpTq6iE0DVctTsQOgxzyRrfg4MLllRC6gjEnxwza1TmqfimpOnMkoFHQWzZwKSvHTNsA
dg51FxTybK24GuV1LxZzycIev3ROgYEJaPmFeXt7cJFM+0cBQJWlZj3RXrZgjXJmzn2nU2s7+IRm
fq0WAhRbDqvAbPEK7IJRsPTxN4FSzbVigSdiy9a8IY0I/Bz2poKRzgGfzyxpUliJsztAwsNNoOyY
A08aaRa/5DIj11jYkCGd4uvujgcyW6EPx7fOUFVIFWtQPVNytowrdhrT0QzwtCFSL/NMxteylGmh
pYaFklWRD1RjUpDJ47i6q0T/KzA/pSbti5uryWxk/CgHd9Qdl/uQYtkKGYG2/NUgS+lF8D0ljJ3x
GDYaua5mwOtHyrgLZJdppJ6L80JI1xQzdpdsvIjd9kgSyPxzAfDlJBRjaxBaGEBWnxBUAUkMrbKT
i+4eG/NG/XmLxQoDN2CC3ZmwRpqaVCTYutWrxOaZOi63l8FAdgxS0VAeL2WSqQT5ckzzj/vEjm8k
WNth1PAYYX66VXgu5oWJ1BfhGuF4w64yr59u8imNgXjKDinH0oUqPBxKcN/jNT9jrI9E3XrvinK6
SvuQhSWH4orwHOv2BzCzUugsx24suxPTazdu9dIEx7lcdO1UE0TRJx8KKHkyg4jSbx6i+LTMoPjG
yat5Ntg0VQRC/kZvqe4OvzvESLLfKsKwmnu3Z1LOeXIUk1QzQU1mmRabLn9nZxz+Pu2imamiqEZh
ma0VXM5lYKX4WASsw7acTUtTa3B7KCLxcqc61eFiT4gogVJ4D+03JLov33SvFqTpbi1k6ZsEEYe6
OmIQTulDtqSMYA+sduwzXETj7iDIw9puk4VWr1X4r5lVCVqhQMpcGRQqZOh1CTN4lZT/LoC/NguI
5YfisBfUqDh991Rce2VUyPFXOovYsGOlYBXcXlD/QIv4HBUBcIDBWTY0XnYcJFPGV06UX7MEzVGJ
z4L39Rt4fYJyhC7AXxwBZZ1X/Ys3hXiKzxbFfdvVtSUQY271TUzTHILYX2kZrKMlrYm6lDeH0XM/
mZoxOMkJ7em+USAE86rOrBQ211TZ0lnYUIxeM1f7y8MJVtFchI3eM5SXGfv/Df7SnyGQ9+KVGBzk
YSrayrZUGQpzOkOcGIlmmi9U1De6XwR6qjE/qx5j/9TfAK8WrrNxIAsfsJPvUPJ0lWSFGZO4NJ3d
flZ3qdASzL2H/T7eoAuNGB+hclNbGpBbezXjt6y7q+2eKTe2oJUy3XOviPLEMLnV/siOC8t5Lizd
UpJZBX2R4h8alovMnlzqtbsefTg4zcRl27DQdXdRLzyqfbYUgCwxt4fG20uvV/E4Ji4837lR0sLG
gKrkE2/yR8LeNTMD2RgO3/VOpuZooViW3UsKf0SvBW0Gw1TsdP/uTavz+Zo+6Giq8tHIg9Fz4Gl/
urUlFgU+fnCnAgA3nFAJ4LdoXI4Ie44J0a8ml/k6WbyerIahpaljXJzLsQMp8UkeTZefrrkj6ZGF
VEzKfuWVQ2oy//fJfS0BEco+WWGs3YSFN4dTD8XjflY61mqlTSPpbkt6e1ROAYWaViPEmz2+9D18
IGUR8CaKwNvzpRCyKpe6Myo6RUcSILXSwuONrTwfOQsqDgpOulPMrcyeOQ3CJHrXOebhzEmnzq5L
Jp4sYnjWpY6pDf7KbENSCauozt9nQCQy0NB+RbIjPeXG/dKARzP2NPGan/rVmJoFPSUIhngMEyQD
GzpiOvs0CasQ+lbCU0wV4BrqpI/5dFIb7PVFv18qpVONRB8RuVlDe5RNAzCyePmMozffO9QJLbwO
Tyi13FQGIbh4R/KCYU+JlWOE7jNhgS8QsXYO3bGirpj9o1y/MAo0pUb0S1HLk2pXviHq8SfQRpzr
7fqMvbpT5L1RuSxaFuV4n3Decvg5idXm4ATTnB0eJPPkZsv4uA/JpzL5D85yjFyDs6C/IzYIgO3f
L7qKgftdGVlIRX1jzpseDY7lYl63XRf5g7VYu/gTCzHuPXhS2cMO3BI+/fT8FG+aCF/uEhdSOrLy
sDJfsspIWL31YnnwRkX3XS8e4QHtZgJcU1La3kWdulb2sQXKztHz0MaycXtUOd5NYSWkKxJgdjeo
JCaYnx3+1To7oDXYJjAPV52oAMlsHcuZCQgSVjX98YwnaUjTWirpRp88BvP7C2IDD9vGJdKOrskc
d41Gc+PHl3rSH7I2kN06ByqTKt9x6xoS91+UZCMN1V93sc/d9KteUIZcYJyYR1Q+zVx6Os5g0Zh8
UAoFFQiqjuJDI5B8UUY7HSgeoXsnaOCSLLEbUS4o3/WgfQ7Rj7WCw3dfT+X39DG+ikdkmbUAbqww
+3Y1Ngor7nQQYsMTc20E/Iq3oP/VyOkbG9ewQK9dZZstIxKd/L2yrzzEap8ARc31cD2gFVMO7dXg
rPsAz9Bk4b0allT+oiteNOajNvTlY/GYltBfXWgxbnQUqEgVnUN9HqU+yUG/jRbOnnezlAScGOPa
28grjL0+qYNULWqo4B0dYeL9LIyZYEuuxuX1HcIYUxJjgG+2VjO7zdg19HVsG8fD7/Ew45ZeTjOy
myuknn8Iqn8IxRLHPUByOTDAjk1EE8Lfnpi/wF2oEeGzv2G9QM5pQijMVm2iMg6Lead5U42D5Zo6
0YgXVzKlPlVrG7mJEF1pCAWZH0/x+3zcvoGqZfx1Ptx58Jqn6WLi7F2WzQRaoLHaxkwfH5F4AJrG
lEAq5hD86BH5gkQDUTWRCEY7Jau7VJavTUAgDCjG/02sELt8MmNtEQlJgBmW/i6pPRl0B9vo4ZGi
tJfipgxvAqnfOfQjPnVtPuLUoGYA0EHPj0mS/t6Lf/n3bPNhlKwtkWu5GfbdqP6Li3DTsj7KAG1E
Sfm4CmVaZpkoCbkB8ODjv7b3pDndnPzfLWJDVAcmNiDnuM2QHVklEbENtmuEQtuRPj4S04XhHZT4
LzjuS7X9vt9yqVeamvx/GEmqDP7aT89gApJg/Sr13p2uv6OHlNqXWC2QhxqUCXPWeAbgwsLHeBbS
9TQ3DtRwHcSuTO4XYEx6CTDLAV3hqCAPJprNaA/VdvQPzoADFL8joCv/Q1znrS3TY4yoM2eid2cy
21OBTKvnPp5/U3Et2G5u9I8rEgx5rZ/Yl6A+cmFN/yGyjGbRdE0RB920tYPy8poN1LRMoN1aQIC1
zm+qQRuv+QgpB0SKTHHUsWPGPPIEpJp0Hd+Xs6RBh7/BZULMWZttc/oEa7ECbwwJusT4z9KtWVMW
irrlbsm1ueKR+1q9/uJHosXBI15HI7hqpZ5Lrh4Io8rLMqvb/IB4yM23pcHLuWduefnucxtsi4Dv
ljlJ3iC9ND2jl6P2YofIiIbv7H+jTeYLZxUfT4J6aqaNNz1P+JjRMH56jq8buqLlonYn0vZFiupC
p5LwYFE354bR5h1rH6mOzcmO8sIpMRJ8IxXfRbGZk2+fxb7YeV5hAWKP2SiPFLFbnLHeXfX1EW0I
Er/ZsCEYA85VjN8gAXjPC7oiBkZwp4Xx6XrutQg19+DdAyWsrjw2/WPzUPxanvsR+BO5/IivDO7k
sd4fV88VCicyS7g2ra4MP55bkT81bevrvX/SJxFIQ68OmuIgpqNm6Vaz2o1TWaAcHvxzroIHkYm4
LCLpuWbY3Pqm2DMzx081D3xVc55Iqv6jW//DgiKc23HsdAliD8o5qzKTX9yvXIog3LHCsGhH+FmL
2HuCnAPf6zBQ7eWtWQm1sYTgAAS8yq+NipvsuJSizqUCaa3IfOIr0QXpSE12R5lvGJNEm4vC+HWH
rNlG1ffOEu4eqiy19omZfgKKBg22KI6kdIz9Ib3gUEECpBamM0hs3y3elurPVgMB448qTcPqjGIh
mRWgoAbTsgpBDogSDnoMotZXM/u99GVe2yq+nsID5Umcw4sSKz3AIFCnRXfmwjB+mVCXATorZxaZ
+VZCEJppzSFqySCzAGh4ZWxG4lQnOiA3I99GFDVskQBUUnLxI3EHZRD0HP4oORPVM6NtNlLsRIw+
RTh4y0MxGivbdw5LL6Lq3QpBoF78re/uGKQINYQvlCpC5vellcuX9s2+F8I+s3X05aIjoM330HDr
mmITSBbyu0NUG5OH0KW/qcXZVw7AiliosXy1Cbbxqzq+a/u+x2u1oNcARXS+GZzb84ed1YrjeChI
ECLiGsdZr/Ct6eHE6uSSHcSNlvOb3owbTff3f4QHfnC27Ur34jw5na2cJ/uoGK41Ry5SXEVevnWF
SjFWNgXpSameMmIFad1HkXxJWC/3s+Vsc45nmSNdSauZNhMJ3SHGEzyLoD8GTim7HOFRl3sKPsrF
pxFkjSYuAtlj1TTnNNtlTDRwIbeeJ8aWjJz656aLK6FXO0JYeqt/AlDhqTXpKtZwrshLxHNl9LOB
cFC8Y8J7UG/NsYn4R2Ldwxpmo4LTbL67j4QELF5fxG1VElFtDXAisdSkrfnhZwlqc/H8iuKOuaaU
T/GHXjL52UBvCoH7yuav2rf0ZOcvirGr8msWYQyPJkRsxQgQK0+kVFTUN4LmLDEd3EcuNXlrl8ee
7I28sy9kFlYYZCoRiAb7h5YkcXFJmC0+rILHZvCBE4lcJT4imywYL4XXqJqn0VZAIDR/ypDp+i4S
Xvi/lAiNrmtnvdSUOrLftvd1na8W1nXNiGNUViPQlqlH/V8yz+p4viLIGTGXAcnZ5fbvR1P9siT0
867GE87FdQqzgiaNgCJYefMJwxVaKG0o8SyU9lvgqtlbCrtDifcUzaaEuKPzcBidEb15zWm4mVgD
VlFRgwSMRLHd3k8rKavwWZ0m/vMuGlRljazKwcCldbuNBnBldP80QoGHZC155yOPH0fyMCwkfXC2
xWDt7xQAmUlonKOjNpCIZyIkL4OX28RTmCvwDxxiYKLpBPLJDL702BnctO0b3kkagaAooe3ORPBH
kwslKSt/HM9Sb/2CkkDTHRh9M4/b3Hfniwm2Mg4NBMhkWzDjflFQAmsg+DkSWtSuEvv8kzV97rQ2
mZwZZ71YclXQqLT9IZQfEZRmTO84AqTd0D0rPgP5po2f/mONwdfhdfI/qaZbkgNx33UdzR+T+mgT
4qsKppD2F1WGyWL7QOKHBdJKge0KZJ1i9tiCrM5dCIYySFXUUU2OVPb8TTmhpHqTFm53ejVw9qSQ
Y9KLeKuG+3aojUTdtIyQ44wk0rviq0P3l42CtU2pAmGQJ3wgAhox7+VE3RdPPYnPs1Emk1MmajfF
HnknJmLhH4Q3VLevbqDgdieTzxDFIGrhLyVyrvh6xpROVgiUwjQ4xPY0lbcNRV4KiaBhimszKAek
8rMpb9rdzFYxSoUj6IE9QBeSXQ3xDEsSBTE6Zoqp+FLQGGsvFmJN9OqLiQGTWRLMh9D0DiHrJ0om
n0aONV94q6F+orbPXqX+BAjz+3UMohrxi/FY3kVzBfh2vVamldBd7rIaJKBU1yvPPq5dmtPx0GaJ
1DLZ0uCUIVOTLqMOMHxzYctPxptQr5RFk8Mz9HaPNk1UJl64AVRH4l4cxZTGiUJmKznxd1slTR96
Pvg3/nVkBusGRcmrWckMDu0mi6eEiPjB9Oly0kYpyZzFNlYkGQaQ3mpG4Drpz2XI8SoLBL2UB1Dz
NcoKTv5olgsepG6LmmHM5YWQ6CZ8mrdI6GE/3pefTZepPguOD2nseGNJifodSg6xR5y3e/4aza0Y
cWjTsvH1vjHfc9TsvvNVrurS7uPge6VShDJCNeMZ4Tn3lf7w8Pysm8U4H1gQ0LFQjT42OAewxJjw
p0oXi9bWSkf5G6dFJmTxIp6WWhh3KEs5qPTgkiJV+AQpJiA14Rblwlq4xXECaemgxBY4Qn8GccE+
yi3Hiwx41giJEYFj9SGyEEAdDhK/T4Gqlw95UcDGGrecs8egyeqq2QGPe63F10O5+IVs8IAq+p2f
dYXGxo2YlrJ89ci5XYwidWcJCcBlTg7sj/PZF0ArIJhPy6crDn6pagz3JWfJ1Siopc5KOKTfMOMT
UHd8L0NbEwPfM9ZmghDJzxVS31Rj3rvoj9qgfTDT+/pa8UE46L8newKqBULvGCq/KjnElbRJVONy
aXYTeSYaCGgNtOyrs5c9EaSHTu8Utkg/D2vKbzpO2VzeYtXxrsQ8+eCjnPK8O5c2LdUJArNm9/2J
JCuxcmjD9kGfBmILPlJVkrAoth+Wbu3/4kt0uKznW0VCaPoo87MOr9iARgCs3j9YtccYkR4QVfBb
Z3Nb62QprynSWQKXzgh7NsXnn0+AoYFwL5gALIuB3AQr2jPlOmnwg5fNPpEAEOMml/ifRMooDqFB
86jGUCwWmMZfgqo5aKW0Ma/C1WSZdxlcjwOafexPQlPcgEQ8wf0lW2JdhOk9NfN2RuRR12xg0XQV
m7+ZEmcvaEAh7ZJprVnA2PFs7p8h11euBHXfrBi82pOVzNtjiYAHIRixWJ5IhpGSowzcQVJQD8cX
syq97fr6NeUZUzm5+ocgZ2gOBBxCyqrEID5q2DAU5bmKXZ4ACy6K3hfzfGJAXyTV0VObX8ihd1ib
qaPU9ycs/WnuYaOtxIkW9JsmOVsJHAsf0wAdupHAzEs6m2GIH2F3frjb4OH3WNO44YHacynWQ/SC
iye0RWqKzCdsvTo3nPHPcUEqN8Ns+5UQieEFvuqSt2nE5Z2cjZWUEplSozjusqzojsq+QfuYwmgM
xWWTGWSKm/15qWQ0ysLFa9wfHlrME3lISBSl5ytV73uKOOPqo4YALbe7m6pIdzmhV+AxMBe6NGYY
Pype1UQSJEPLX+tHV7N9FgQvkJuxAopqwZkHSIGDIYwsDhfhvLkRtly5n+IXXJUhXHDVsW5QbXqx
EDbDF83ani9TyCXYBl6aHQxvuYFgN2ueD7QfIAXTa6UOFSmR8RMObmu407hLnM36QQNfkL/zMDez
/e2F/zMuyKfKSbrKVU7OclGHlAiDJriunGsQyuvqZhi/Jk4F0+2u8T9lOhh62qr3kEWgIJxSjFRa
eBkw6/+7/NGGMI96iNUVs4BjsOvB01qOXmdeBBv7Kg9vAlzuhqcCHTQuFCEHGvwUDJgHSU+YVN0u
CwhDMbVnpAnslzMOWy15Cb06Oeldboj3PAwJWnlOLhH4JVa18SZhxMhsdTVVnM1w2qY6Yd3URldn
pMZrp67sH5p57rhSByoVLVbgYQDPgV3YJqJrtazp5Jb88FxD1th5BCpWo9bHCYqAQIAi98Lt4YEq
KTCokqmKW78t0FjNUn8Oglmmz5wg/X2oUzKvABtrx+9KTC5w5gVz9CFz5BwWccNp8FxopjfLPdkA
ZOjkF4wyrDkxFrVW1wpf0+LOo/5wv7373gxHlyZuuYCCfuSBU2D+mOo52udFJrRYzeqDxEaufy58
gGmn7+XWj+6Oo/GYXB7jYofDaMZjVNj834dUAPP7DQGAijjzDM7yQg22T9ND2iYtVsi1MAnNE9Fp
1p+HgbNZJ9i+2H7C1lggoj9gvtv6P36f5DvIfQtAEtWqhcII4/4//myAfvK/DV2l0E687wIgfkiG
Y5Luk7OeupFalbt8OuYI5w+1DOX3KZI5nrXUjddtpM8tQZl2bcr7vExZ5cNHoPcsfXuGcA9BetO1
C+nNuuNs6SYIgy/tNihbnAihTBva7njLY4wcn3g6yP825xtb3JcWcaI0Dy7VRXSSTSXFV5tyAQ4y
ir0pKNdxbQPjTo6IN+yMqq1ZyBSh8WEtbO7BvqAd8riy/rosB1be59PMI82DWaMIMYoSe946UEt0
x1ZWb6KGoTiu0Ch5Xk+NsVQPgGb9YLuCGXLgY7yt46aaDyFY3PWlQGzT2JTJ6Csrkqyts6B167Ts
cB0L8drXzn6u2J+G075KCsiEVWjaEJWoM4JzsoJ9c8J4lD+F/70Rm+EY9W+cawy76KaB0dJlrXMn
2TvO/0T3ZbS+7j1l37NkLMTVCb/Ai3n1OjsDeBSYQGFH4jY2YPP31AguAdfJ3ckdXLWnA8SVzq3r
lKTM6ePf7fhGoBKSN8dOn1D1Z5B+3RLvo6iWu5cvGgkCOVq0LarIBdNaQZwybedrj8I0nDQloAyp
SjfjfBdYqhmgHyHDRcqaYJym0YvTZHmp5TP/rwQfCrSJB4F7zNDXRI4S0rH+nObXwvIBl52ej3AR
RqlkFWFn/78xiT0hKHHYLJgeUP0mxvq2NcoPtjuLUtRajhwnFTjKqazgJYC3a+plq21oti1bLdrQ
gDInl8r7m2dpOH6/gQd/D5a8/rrohX5snN2LT5E9SBb7GO8GOTDoyrOs48XV9yEJyvVKucyvpcKU
yygn3AUhVsh+eEcUseuKfMgTSiH2BRjzrKvaxOsB2uVE8W7oD12PsbHqQOsTMSJNSQWqhCGTzhXe
U+zDmLece+aUj69W+nYkzuNa+iiv4ygPpWnCpfMj+P7lyiLXL0AFMw6U7I4aicp7carw26qL6cDw
gK4aThZDAofFwH1j5CuJ6/9RKVIzjtV4EBgFmR9dMk0hnXLIepxY4wV4wn3Pcpsf3Yv+y3nFKye/
AL1oMnB1N6KWcCEb6VEZ93eH4HES0ZRB42NOFPB9tPlyP2Ii6q1SQWZaGn6HaVJaQDIJrv9MSWKJ
Qq9kcJUoybKJ1oO8uAEez9IpdGg1u68faNHexiJa7oYv1EFXtVrt0Vo3V1Jb8h/67H66A4gUPlK/
GE+bZp032hsArPYeT8UR2y4GB3/eEaOr+cbDyBJd6Hgzklec+TvbeC8w3M8HZVaRRV6BhXPDbSsm
6PgUB+RnR7xSgrucFGB3s9bppvKSZ67yzoWaWTMTVrxUTgPhNlw5DeaHcQhqzgei2RaseaZ7RFYU
BqodnWm/ZwRRqiKHbKJiSvf1TZlzf/0KMrtesBjO6jbxZgj9pF/iFPaeT8Qjt0t6Y4f0S4ZYEHu9
U4P1NJ902oPzUA7/+d6S5wiMpjE+lf/r2Ke8b7DnpXwg+SbqZL1TniT5Wv062RKFEGMd0o6rYWPk
pnsTjsrKkhDx3bVS3DO5bGiM5LxjeIe9z8/JKTJzdJjPqLFboWJlbAxxcOS30wYJpcEwpqIr+0Dc
kIvDt1O3AzBLsHAUFljGG6VKXWImrfSH7zFGKluu/uVO9YiaeGrzYiJdphwDNourudn/wXw84bsy
HdvoXsIZ6oRpTa+MeERc89FWSY5jAIfwO78dwIx7Rbty+mKO2RgqFdg5UoU7golDAXXGJsKdPA9c
fPoN9EL66Tot/1yI+ch7afP44g/5lFJfdfbF65HDe4rfzlkJR08cHIguqq+EGdDs254qAEvY9dQt
zddUSmuGJBgOZ58EmRotS0UxMWH6oOcbYzovDAUws9ewzEGVxwANX6rPzA7XemU6Nu+hNBWRmW4O
23GRaTtK75sYsP5zeG23cUvUk/xKpmHSB0DdEHJRkP544txI56ehBEj6F202kIx+nshJNaYU/YiQ
VvRFfsM2EdcJMJJ+MqRuPpbdK5Hbn1hODfRuVMBMSi+IxgKkZWDF2YaNNfaMPkKm7/8pmvf72T4E
2fm7qr1Cuw4o+cj2xMbXWKc5psp1NYul1zFaSzAd+Pfnlv64YjLQqpT1FVNTHats0XLcYJMPD//R
C76Aw9mQ5wmoR7GyxHVV4WE0FDrXZCgdlnudrEa2/535LU5GW+OUAHQndSjAh+TBzTyG4bSRaHQh
njj3lyk7qt9Ev2PIuYB0hdiyfEWHCG1XRkLZ24nX91MLwP58fAAwLpxrcPVbaLZbZuxY6nj0pCMB
xNev3F1HqfVnZwN53WIGagVa+zQDH8zSshpRRUyvSeR+QEdgQgi2GM9xpZs84Zak8p4qYvkZHYoN
ZFY3UyMBWYytkVqtTdWPqyMaCBvWVuz6BgPzo9AhmxWTT3JH2mucIuoDznsw+Stc/dMEy8NnpNaT
JQCXxbvJTKdHyNmEBUF1vVY7e/dO8pMcFO6GDCpOTdhobIymFqpSfrt2vPv5j+ft7O312BTair41
PB0a4+aFxcf9gagdHxbbbgc0tip+qLv8hzSWk4gXHaDmEXQ9hKaU77odCo7SK2Cj4yuoncnCuyvV
qej5/2PjdWWHYdQ1BIwRHTeTmX5WZIB0njyWY+vg3Ge3+ChEGVGmrc+f4unNaxxyrv43rHyoAYOg
zjguGKaLIyD482WivnByGRKkl27oGDncnrdZmnqq0cXjn+1+7duuC2YdKauDUJ17e43oooxjku6h
e0extdiviDslKs/poyyZ0XwlcCHdMXxj7u4gFY0oFaAL3smysGBNKE+fWKsmlVAK3aN1D8fWERcI
J8Sjr02pU/Z1lzR8By3uZb/Tnl/Cgo58vUMUKju2RB28nwPo8uSoeNxXXPt9GjTVqTDoG/+6fH4x
m8nV+O0JYyXc1es723RPdESb9q92In1Jwc86t0pYJ/I7ER9kCEHh5sqOg0X8yEqJyUeKgp4Xjy9O
wXlTJ1xVOaNLJ3Ypanhsqq97ITURzwiXHbp5PFXtt+ts/z0M2VYHLLdqZOfB8V23J3uFtQkUxOp+
XgqYbmCJNP93WWfV8cui6oz6a1Sr+09CyPfua3Tw95//c1r8XCUuHRvPGHtBDKMAQpAbMIP5QeXv
Zt3fxeXb8mnILVgHWlsitgr7U1I1DJZ2TY6kvVQ/WJecApWOzwN42hwttzZ5ldjWc6/u/bJHUQ/4
q1tU4+Z5l7U5wp4jYJYADG31uy+P2d1vEinSS8q0e1DmsKhlIiG2LVYqEr8PqRd7Cb0U0PTYtUoC
epykAd+9yw6PjlzSxxzLo7mt5a2lE9SVHZ3sppDlLR+nKcGfCr9lkVPKHkpb/KgI6udwg0T+s/zi
2F94pF+An/wbLueq4inAn4QYk5IhB//Zep368EDsc0rZxAedGSCPnpnrAol9xIdQFJihaM6aRKJO
DXN1aytmeR6hx4h/D15QRHQOt84RqPUi9XlfQGOjF+WGf+CKU/T1qkyzutsLpuXQ6GRQecoepRTj
ldTP61/ow7f/RQFDaYX/Huc0CiCrcNVgWbuVTE7qgEBMTcORJUztkR3l97XviZL8MFWpi/KKMcWO
tOiQ75o/RCLw2/0lvCxbeVGQ5oGD0BCFdIc8DhGQ2NSnW8aMj4r5Aeg7XyRrYGlYXsW9v34+DQpC
djjaAbCIvq2CWrK5oGSHFMngQB9tEZehXFOO1MacdA6RHdhsaTpuWsGu1LeUIYmv4WV/58LhTNHD
wdRYht5m03gzi2k7n0zBxwNoUuxSzKtMV1BF0UKbj0Vv9veb67MeF9J+cp0rn7rS098dKBQyPG/t
sK1lQPXg+gSBcG0bmFN8K32QwDYs8X+GEnUivZq/oWMQZjVz56Fmpfn/AkP20dRqICR1eKVi/B1/
9t//eveMhReEqxAd6PzawLxw/hl1MeMKqBDf4o8oNgLw5UWynmhgYz88imDe+3kQ+thDmvO+L08D
O1KZL6+5BGA850yKzJi/Q2RCkczQRBm+fizB4M8pIZ9sTtqlaV6qbRUj0EKRm26p9gAJ0zVkSm3w
bKb+gV5aMLjK6RQFfZVnFg2iBU9UW0rU1db5tDzv+PjblcOW0fFchEbZvTNk2+L3ab7Bpe6CnK+6
Yp1u+/eV9dLVh7Ldc4GO+8N4culpQ5NESIPXs8caDOxgJ2TGmCJJ3xCvdPneYdRAfqdy0EHr2mwd
sPmZXq0JJCGZPZhKtRj27X886bFc8dcQfbpPI44qKEs96uocujXAk5XAjHW9w6jwK9ECoIzz9jzJ
w13eVFuRqtPWUQTLdx+RAmIp0KLuhds21wk2xWqfE4ziOkGsWkY70IA8Z23sA4e2PUeyL/oWYWN0
/KbuuCP4npcpWinYoy9UBoE4yOXrakW4sZdWsnGIiCVWHMxIXwlRJRm7MAb6v7jhpGqB9OUwnjDI
w6DGcCHWzxnr5sPxH7zosKNF5kFFKChRGL6ivWpLh4gtOD215hx7MO0QRTtYNa++XHxV0w8BwknN
7sZJPT9NlZ7NOi4/5rgPfvuSvaOx8M8HRbBbmhgxQfRsgWrp1t4cLl5DsGhH4VGnXG6Jle3SGVbE
LUD4/8+zLrOElCshSZ2pJ0Y4t/3cRBuIngq/P3F3aPFffDXiaoiUyFBuJKtEA1zrRl9ezrKUAd4V
apM5Lm1JvbViLENSkJ/TiUJp/tKjxtPk8IkKYU9+9j06ooADcG7IIlmdUoXBHbYaKFXna3BHJlhd
/nvxFMu7+yiltent873MG9yvaZla2K90NgJ3Pq9hxOBtVivka7Ps4gCJIPcRnQ3cOBVxQXD4TlPE
9K6bsTimhOEY4qKw/iCRXoGkzVzIoiEbcw9Ba2GnyQQc99HjGvfXoPXIcKhRKu3NnYChiEVRKu9K
dmuSZ/hFyZ43QmRXjsZwAxNDZU2R9PyKmOi0X9Kk+VVOKB58dtklzlY1pfL1wcdvZzHauiB10Ue7
T0AlxjkfE67nzHhK50+kAZtTba03zV12A4f2of9jHJhTi+3jDAsggkSIf2+Lu8FunfJMijasA/nd
Z0+rCWqfuCs38CQF+Hdo2fZ7QRLwzECCUYbEztXrP3jruKW/NsWpk1eqkSN4qsXuHkC0xzJbTl5H
7XROQIlLczMzGux53rqQ4ZYaVEfDtVitNR50HOWuyocPIPBUYJXMDo73w/FTzD/em6hudFa+WkG6
B2+Em0BGNDPrRQZxfwxQ7DUCwoVUm2FCVq9zINAdRsviZi1d2VRi5JBZ9tk72f8sSgLM8ZFRD2tN
3w9hOUsb6MizwefJJFzogjuaXCaxmQqTU0c4rQgMIzln2uszzbv10Owl12F/RQ==
`protect end_protected

