

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VqgplFNkI2rH3rP35CdiLJAesBBzx3ahYCWVov2QY8pnSpbbPHZzKXALTXuf8Lg9RV/60SesvL5+
Tx0kf3Xi2A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YpVJ/AkbT/7j7nP1FpW0u/1drBu1Ym0xSQcZVVNR2BH9CeGHgikyUixQxXpCsKnhOEb3pzk2wV6b
2udOCqgzaZfDIjjaxTt9/C6XIY+oMyWDycOTnGwR4Bf/A6rFEzTLA91kxNt5/tS1PVy+wjb7FCsa
mgkYj9eNUdtmSsLezko=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pSdvSF3+OBx+pmFIuKYX+lTRtc2CK1xqA/WmTxOA/9c1xuF8tv0giSEc/96tBGsFFqc25YHyYiXZ
gYsCabVJMk2jc2XaKW+XFrRUGrQYLd+QPrzsIggnGqpN1i2vEJ2/57QIQEt4pR4jX78IzCIP9B1I
Mief83M338G9aIgdzONBxsD1Z3XK2M1fqZBI+UT4b8E2guDKnWsCC9f6WqxH/+ijAu2o7kXfkz/w
wH4eaCjn38eBIq4U5maYpwbVxvzCRoB69hlCwEEVDievRmXHouMD407mzOTwKaIkf/tAbFyB6i0D
s5Boa+TiBtHShhLBGBRqGoq+2UpGEaVgj8o3hg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HVe+dxCY+VHrZ/rUbzyWsz5ix04KcDyyUrFaCcS4yZ4GTBKi9GYUFVfTsXMpSX8pxXieZIsbIrAR
8ATsmu7QwmViHDzOMuS6sHzr6e8dC4A3UKQC6xKKwbJdSWPz/il1AOb6t1CcrpGMLBXMZTBj00R6
KptQtwRx2C4sHo/bHEs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gr9tWfnRHlUz7X9jwun0huNacy2IvVfab84T3X/BBntsyGpCEQL6hR0/eLuvmgsVt+peH9UtRKIo
Mx38RlMVlftuoIDUnixeoGaAc4c+4+tb16q3/5V7og6YvplXdBH8LQEEDNM3+H5ouvTLLeMul2Yk
sNNMGtkGcvzxpzj7QTVn+eSHg5B5sba+LhJuLxq02/5r329tzFZy8dtsa4HltD5DQbMsj44UHU8g
J84rl4f5z2tzAq3mdpwIqfhK2vn+BHZu8UlcbrIJKEkQpY9EPDhgx0vX44IIfHNFCmG2MgNy3yn4
3WNmBdtLjzwOjBTyBBtqdvJWbuTYLVDhGJrWQQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4656)
`protect data_block
1Ec3fwLeQvXnLrI3I5TGWaC7JjZP0OfBiDOcqHyPmbs0rfO+bijCIE7SIpws+EJwl8bIzzAX3XEm
RpOFcEg/PAlZqa98jcQ6DYVgOo1H59OLrGNloD+oQIcNmYJSEtn3ftFC7cAqr00twINtsg6Vccce
/JwCtDQVJBmUqh8CO7SG2b5InXyl+MiPfEJXtkiPD0gUbqra6k2qvdduqWg8pM9RfboJuL//Kif5
F6cYYP/3Sw4NuKQSTP3HtlF9vh19XG4EAJeveVV5P70NtaBp3pMlLpBSuXhkx9I3ELGxJoAm/6SX
WS2xfi47Wbm6x78n9V11kiOsnPfOELr7YkR5ahPWRFgkYRT4OE7miClYrmUxJEU+VUtKJGmo017m
WlcmcxweXMavfOBh5+PGVIxydTuN+YYoeEW40XQMBaIxxWWSlYiecTikLdZmgS/Htr6SJ2i/RPWB
9EbldiUZTvI8Iu/MGhGarAEwrbksynu5HLp5zzEqAdIINKWjP8v8GzwmKVM/G19BaHOriAtmdHqT
7Mc6iU4WqKZu5ffG6BDtNqeXaPbrWVMTrOkm25EG3OmYcFmzoVBztod+mJ7OE4xAyq8xFs6rV+/v
KFIdaFVKRJ3ZCRarGqrv6O9RUE7s2n6F319Dzc9rKsUH7HvwkFTbbJC3Tq4unQ/Yh0aefhzJcbnK
vkdZxOcAvKe7ytVxUUkowZ6eYcAqquTniSloawhp781CKhlXfaAHHR1J2bHVIQuwFiEtqFE6Ro4o
ZFVjfZr4cz4DEdZQDjqQMKTvZsRln1fWntaIAOZEkYW2PZFMGHGE9UwQpOhblCIi+cRQc4KWS4sA
wcFsVrcp4Ka638+aEwXPQU23TokYRVdDFMkFwqfeNMYAwZt8GhfBQRo9LFhwdOraM+BY/uaoSSfV
8REs9mNzMLSE0dQz/yF0N5dhUvOCVIZ0MQL+l9RM4hl6Hno5mLg8hq/26ZfXaGCzRKdMzP02L7TV
lwhKBsIXcFqliaJFcQLA7IfhJ9iH3bB6uRY/9M6VOfF2FlE8zAvAMBEzwDJTe1QZnspJ9zD52CW+
hpW3lytpgLNbN6NMrqe3iOOPGG3tIWWJ0A31SrnnzthxZDq9gwJKMYTSfXqOcNlqA3Ii2t7IADR5
zY1TdLa34fjtFdMqxgLjdUmHFSeZWHdux1M6FDnGEm9GTAkXFqPkleg+is6ppM3+yc9+WfNjxiOx
nKm3GueI4K0+q7Se8y8ThwYUuSVGJJ1QH8QmeDyChuHAA86Mggch1ZOmahzNcj3PoFa6CgM9bWYT
5vYPsfvswVKdfG9baQCknJDid5JP4V1ebIaNSbM6Gy7Qgb5pQT4sFeAST4lFI1XvN2b8eA1OEbV4
ioABVdclV9+QjFpQkItb+VHo0DKAlgcDcM6soUdQGokVkLRLjR8G9vKQs5N5myi4OsH5964YvpAN
4DjIoXFMcEqV2UGM0u2AsIkz/65Iy2YmGGpDUbbwMXjlYiMyTtWROcpwmyeejGXIJPimqztqZDUC
dHQ90Bb8cJ0RMNbAD/hE51ijjgDOv6htX+3DIRwjYF3LBfiNQLv221TrMHZKcadO+F1//RgAWSw6
jDpOLzbWxVXIino4wNOuI+UeH7V3eh//cLYBIuesYc0XDmz94O6qx5HDLevufwAZfToDe9PHfYH4
2cBzymbcg++RR0rPnECdTGQRBCMRCgp/iR6WdjIVayA07sX17SErNjDnfeao8tb+M5PSHqYhPErE
gQuqxvo1Z1iZq5rXS6Ber9ateXLNq+mN11J3ERrnoqQo33pO/al9WfE23ZWvP3BjpeyMxcdfMq2t
pUx5RRCA9SNJIUmOnzD5jCRs0El73f+R8+ZacLNsZDV8IWLJtBz1NaDcTib2cAvvILRGB0UzS0b0
TppnYuJeS6lkY7SxsKyQUC7o9iCGUBPAIFMgIb90O8HR4JdZnwYkzOCFgj3lE8ji/U1OtU93RJc7
RUgjrrQSHxNbkxqVwNFS4ZfEvDeUfYdzOB6GzQ59b+JO9UU21CcDNOJzYAKunG/PXQXaXnNDVqVa
lxLwtHrfRj1u27bz0n+9h0fSxUruVIF6rSX+0XadsAk6v06cQJ2jtyaFLgGI/AQUqoZCN91wyZxJ
gMubvY6c4CbGQDWCe/xzokZjh7dkg+jfpTR6e1Zqn41mGRN5CEAJU8Cf3GJpDnIl6M1IeUAJsVLT
zJ1Wo2LeR3jYXCnadzFo7eZ5fLXCpdZbnpOB0WNpx977X0QfejlS2MKjGAjVKM/GqveEFsbKAJky
xoXIExdoMREHx3Qx4vBu6AbRSSFnUyYYtiYK3CKYdpGgyZ4eoQrYDUmfSPIThOyk3hTtHrx87UPG
2z0qW6CCCIjma7Gn1jjY+6iOCedXjnD23iUqCH8VSi+/1N2Xq4i7+XtNLhACqzjlItU/kRx4CbQX
I9Uob3eTJ4Ww2EDC7l/2eHqFRJHSqyoZqcdR7z6oEqdED1Vu4l6qtn0zcBVGfPOiFVbIvGpoDCoL
ASPyF0ekEg7DR8AUP5Su2p0n+UZdIlzOdIwuCFsBh8i1TcFocHB4+2Fx5dnbiVJNRXjQUuN/VTwB
pxuZrnjMnnkJNHo15TwoXROIsbWoSu9NYa3xS2FBKNuJAOqCtT+7G4wvkUC5xDnKCXjX+FGBZdCb
wfehpkdTj9A+3ew8WKKbP20IRDX++Lso4qQgsyr8BofAbsVKiIOu6XZ4hc/5UtHndE45qSX3khtk
svx9+HaEnS8gLgX276NiwiSABJatEIBxIbxuNROGXevuzdkcNu+7U54vTmuPjwZhZDBJvH8znVYs
4fyvRao55CCLYQYZvBQrpEFlDGamWLIuNj/4MHui4AtBHVKknv5OTXKaj7y864DAitNEWNeeOwqR
85KAOmvpjXROw/wDCcROTIxmjltK149AyMsyKJgU6Bbi/8N42BZkxh2W46ob+N/aaeWCTH9DTE6g
0H1p3krT5yIebe07Yc5hOHMerDTJWTrcCraBtNhoNReK2nn89TdFsEIij0sULUbHlRMqtZcGoKuc
onGAMsi8iiK+Z5zwjWb0foslegloy7DoFzogmOr5DXflg0yeQsrDK0pjtkgOAnE1PuJPaNoJOB+m
PxQ8eAZPyCo3m4P9zUejdhs+LJnU4e8ewvSqu7AKqtEPjGkujRDgQh8EzKnV1Xsbjd3O0l7sXHud
oWl7rCS+GHO+qO3Xr51DUbW3FjpGL6NKx6ZmrFWAWj23yQz4mLhwFH+iGINR91BfX9798fIHr/OU
xeWrJPUL0JK3mV28Ix0P3BSQytJMXBVFuBSQupjKOR5AWfINcpmoGH1qM+DvKjoHoMWpbscM09Da
fL9P9DKYF2JKgpkUrG2FjVyuX0mVDABi4tJBIPMlRZLAy04bUCrxxAULCBL31l+G2z+a3o9FuUBr
sTlKeOH5YfnUgGqNO+9bjDdJUPVzeHDFusiHX9fW1IZ10VrGMVrchakgJ90cEqMfsJoasa2OnYr1
6ok3H+Nf0RAelziwEfBjjdv7QUFbHRTypnAjnuQ0pz7rjJKXoXZy7+dKlrwVWOjJXXcY90uy8QRh
S74+Pk8+LYiik/SO3Oa+Fu3dsk8L9wQtOcT6onfs18CtYaLTcQIFFaim3qLWbxdXAqyZBzEl52SY
Sp8M2FwhWm5AbnEYGZFnvDaRpn/eKUZlpk9OdS1jfsWkyKRHbl6B9JH80cisNYr7RCHqtOftUZ7D
UaHCr/jg9rXIkVWn7V56KqCY1X+xEmEDo3A/y37sdwGEJi55gUPRFfW1vV4RpWGSRb/JJH5WSnp2
fAagmrjP0U/WbShkkyMuXeGpHLIx67BDlGd264mVzCsLoSFgrdRQqb6R0wnzJYGoAGLdkkEAIPF8
NsQotnhg/d+DsgdGlh77ILcmAlPBSE99uNpYx9NGeomJmly6sd/wWoTQJAjcOt61C1lSIdffuOfV
J7GXzLyIo0o7vCFWMlNyTYwsBDFeOSn1Tbvo05iVmKdolUK7RafbZjnXK9aj+6ueLGg/6GlbfSxV
wCgDEg5NmwciDTb9AWOI69WMgSqN4Zfgd+Lwu3wdUlRpAJHckmFmnmt/yb3onBvwLRSk9QUhALGT
PGp7e9zP3LuPxOpr9VEcx8X0d3ylhxp4BVrNBueUrh9SqFMEeR/qIwYJub8lbL4A2N2zld3+2N9Z
vJX/vm3LrngdMLMkjfcGhrzQh16sQu/npRaLNnfXGrSaLFeAfx0wYbHaamdsa2L1Gq/MbBBsrPeQ
4Ev9efvUWTxn38m7Ems0B7vI+F9HH3VCDKRqMp+2UKGRqVvFz2dcMT/mPj2jYYIEHA9Fuw9lt7oV
V5wp47Zso0OQ+yp4JtCQkLtDo6vsR25jYTwQXlp0WCoFCE0afVkcLBK4KE9/7PA91w1+ZjPV9Oll
Jeda0TTls9D09dcuduhPlQMSfaE/8loXC+JSEFzaYKXxNjPSQXYcrfy6T+Nx6Z3RUC53iqG60Rdg
nJw3lKr6P/ik4MFD6RxhaeXkrcXTCpQBd/P9TMIAkp/tPXeYPnQpAwsOt8jOaI6b9WxNZeVxW0pt
k8oAgS3Uj+EbQjn+wKVBYMD9xEN9hePowUPK0YRXBaVW8tw++ER/72Y+bvkrhVD3zV/S8RNCxMEs
23sSMSpb5QytpEO+LpBGkxgx/ZB6+FrUrJcnquritb/wNu5a2DRV5AJAh6qvMFUOq0xhc0jnobT3
h5LexPcpmhCnVGhZYDJoWGs1HECcRlbwCgR0nW5Qtn4r0ZuPxsXDNUx3vIuSachh5ktAzBsBl42y
LwruAfzIUhcyM3sd0XEx/FzNCi/cNheVJLkGpen255+VeW9qMwYWrc51fZ84jDgFZz5Ui69Xgfzb
R1oTXC2d5Iy5MPqZ0W1rE5xLTOsVfSFd5ROj+RHMEYCrB9MLM2z9OYShTrKgxsgTk4dCQQd6k6dB
NOw2/7aKNdo3uPEL/QhJr2XGzwVRrsm9bR5/E4a3u1hQATnuVuPiVrorEbbq5TlKwlQ9sPZimEfN
XKY7wnWkMvIoI9f60Wl6/SV5H5eWsMkyF7qNgmGO+nxLsBLHh4m9iiB0CQ+m7bWliXVLL3CGZUF5
iHeROljY9IId/tEcgsdbKip/dAMz0nVsaqFX/aWCwE8AvouFats6ffRTi8wTAf3AJT8UE/2cBKJD
F+badqnQbDjBux9G5XPkWHv4wOYqXI0/hcM34aBp7I9nMNOol3QjqCxYLjCneaTHoBaF6SPC6syE
HaCmKr68bDYyQOStp71DkMQl9D/DYP2jWooXlRMPYLq9DtF/L0wNkouOlDsvvHmomvMEmJNUCid+
ecWMLN6Lgn5nfilI5LhjX7CNxooIrs+rdxvZ3IlG1lg9y20N6ZY17D9t6YpTlMRziSeVlKCUCCa9
Hsxvmm/Gb6GDpY+wxPvEG52zeXa5qeUDwIClNaZ0iVLPRGj0utMuJ3iSkgSveAn4/mTYnLe2iXrs
aG5np4OFyZcTQ2SsjtGVzueKJE7iWE6VHTQ2jzgMm23Sj6fVxCMONQJzkd4F/4RRHPPbrjsEIwHZ
GDxaHbgSel4ZglG9dk0mfjRqPuU67Hxj1xml2lhuMGGoJYpt85lRHz2t697gso/Ujglr3/twTN+i
8AM4f71EEPQtnFXo9dj1cbahmU7o/AhhPOO+i6r4wjOhA0mt0wBcq8tKNVO+GuMqFF1nx2e2x1nn
MEur/otOXYwOu0qp6U0dPHuMn4YFFBOAZeyZMpmlr/4UfAuHEDpbVeE5L6KlN8V0Y7r703BZJYYp
Zi34hcHAbEhzd+G55AGZTqsTc6rTxaSzwt2jvLAKke00N2ReUOpJxfX6ncP+2Z7HX5vpFhiD3VU6
ictuOMWJdoa8RdfBPSlV5aJvMyBX7ahrhU1xFdXmAwFdB1Tg1WIEeNQtscm1e7qO4eBmMUWvnk5u
kHNDbkZ9a4fP+sWkrhKWEILDy+0EobynM6dehvmxUXKrtUPKhjhDoPb+QLQHsxhXd5DEBiwzCQR/
5Q/LSVAZxqwygn89QSiQJE3FuamzKCoEy6CfEVQVSM3X0rGXx+1F6AJ4q7YDe1oMTyZdfVh4Be7X
vZ68HI2m8ItUjJTILG1Xwi2PMd+jgcIPxexINdMQCR2DhOemscy5S/DE2hr2fJ9ANJUvzum0+iaa
Yrd8jOzs2k74f/aAhCK+8iFUuaZ1WrtyiHkWGQWdlRMGNrfj/hhV
`protect end_protected

