

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Syf21YU5JnKptD7LOLtaHZM+q1VIhUFTxsmS2r0ofwQ3ushsF40KxXOCQsGAnXjGfc9kVb3Bn0ME
1qO92hlu9w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dY69aEX8OSz52Pib+7B1y1Wvr7162ZPVuHYqEcMQ/oCfJJrpwF+oy+zQI55NVyz5aWKsTxE6uM7J
HbTWuphJFeGo7mzwyRD7dy/8IFTp8OHV9aN/fKWepd3R1nKJ/+bdmSsliOOw+inM7pfx0a3YODTn
FRAbVAMQuwe+OVuT0dQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q+4W/1zvXVAi9QMds0GLwNMATdnR+yvz4Aqge4tYro137XvQ9NhFGdF/mXOn40o0ijOuTLANSGZq
Y1fe5IvAhv/BzIqGLvvBSGadUyLWCe23JTco14xHGh+EcGpkQzSMsD+MtFlsKB5Lh4Pk7Fki+zjY
CYS3IH1yrExDySGaxaJ/xIpVmbcDUIB29ts6Ape06rDNuWSEZkqi5ATlUPCMrVpXs0LgVRBipzor
Mr/lCisQJrroeVDmbpQGOxCT0USTTIePtqKzCRURmGOM39JzikVR3QvCxX3V9zs6LEiHJnsAr/WX
JYHo8e0tsbF+S86/2TJe/j8LJK3VvghHADCdOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jFetHSEk8pl36rsszcvK1lxgvI24/D3eeWIqqx4SgMWK5zMch2RGKDJVjZdo+SXrQZtG4vIfoNJ/
M9NL/crW7IJ+pa4Cb2wH+GD2pA66Yo3aRE1Ld7EknU3x42o8aAXlhcPIjcxq9tmSO5RxnhMKlfjh
dMPsoD+Mezyol/EwGPo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Jgq62sziWqkTYcR9/y/ZRFUy8fWL8zR/UZTwiK9JRpmOKe++dsuUuVffmjjAGJoOkGM1fnXZqKj9
LDnUvlqAYGJAQrwT7QRdCNBN9eBMyr6WJUCOkpNRo5aWbRqVpwZihLgqtvesSbzoaKe4eDRdiEe1
xKR9vPyfNmAnPN1pwf+2YDUftVl5x4CmlqRUCO2c3iETzT+xwYzxqYKolk4Qa8DTTYe9PvjYqn2/
dj/jpAwnTcOKUqpa/3FaAU1zgLKWphnnTU+MOfKNP/ow3ZLVrmyiraKTGZlBmdJF18AzYgHb4rrc
8Z8DuRLa762hnT0qbzjf0vtKn06WBHgWqansQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19248)
`protect data_block
I6G12XftaevrI9TMwMIKSAGNl2XgDm7mTdVGkecFMa0Zu9ZFyi/k9OAVEuN8R8GZEYGl63ISsA/1
KvkhHwpLO1P5j77gSokXj3z1KoKtaz6tH2NIeLHFwp7Q1cDdMA+ZTc6I60AjBBuLF4cpdpGXRcmL
POg3ILta80hxXlhcT5lFkOzD8gyFXi1DT2z/MMf33Dwy0+kJI4L5EBiKvx1X3FxD11CbZt66kZF1
nDGq+mJzU9EorO0Sx9Bu36aAef+mR/zuZj7fGkGAKLesX3gdOR1GjSa4BzJBZjETPIUDJIr42UyS
9OSvnSYhAoEqqivPN2vNwULxQjBoDvhVyNPTkRXIesulure+p84LmsE+GkZWNRinEmn+6XYtov1I
5PNLmEHIgzriYzP+48RCIRBrveqMjVako79066RiJOtKgjRN/XVP7UxQyxS+iA4QDVFbnG8ViJSB
fILdKq2sg+eX/9DfrZuIfWFeDcofvaV+vw+ZW9h4HuMBnCtpP8TmMgo0f0iBF2YAi7mMRozWu2OI
EtqwBpv/nV+qJv69Jqaidzku4tTnVGL3RgBOKpc9dZnKBkhEG9MGEQCt/HbKL8pZohdECki83n1A
eajyH2OLwEy6iUiuToWuZcAHSY4HD+2IkYxRXmOsgdftkNeceN5nVC/H2TOS+j2sB46V+xcTNUm3
53eBc+z24F9osfiR0n+JD/k4i1TMWyRiCW+tZr338dEdC5UN7S8cwEo7035UtguxGXBWp2LC1pbP
g90ygIH9eEFh6EPWKjZxwuRNhB1Ank2CYa45hWgJOvLtAaE1w/8PjGVChR/NREQaGX8o9bKYrQZp
ATIkEqLj247L4BUbtraH9ecCvEX2LROShkTRb4JOKBs8vr6CyxYJbAHI2lEMr478N2jzN68VbA1Y
wvYnsFbx3ywR68SXloOrQYUaz9N0zgIVB968Ni6mJdI0B17nOCX9vXLpjNSmGM0Hp88FzLlJ7jDH
zhNK3+tCprqfFtYAKjCJ1nqMzQxbM8c2B2er0fTVgx6Ezrf9ueuKPP+kgp4hFiaDzCaKlZAy41+7
keUtuMGDWtPfgkEdCow82wtv4JfpmrWFoyV/Sj8bw7l4ODljAutBpTCK4mdYn0JyNRBMwfpKfSy4
9U/R9n3RMMlKadAGK9lRLU+aoTq7BwFt3/MeJFT1Iu6bfqNTu41n/fjVXDiQ1L/UyDrF21Wwf0uC
kJq+wSMDnlI3Bygm+n6UspgScPZfF9JzD41XYpFVXEw6gAX9akf8WGMOkwyQzXHozsu+mrsT0gUK
yvpuViRbxKqEZBFIwD+LdX8BrXLAO+7KiSe4+LH9nuhvDKVXM3J3opXFZrb0TKK2WiALm73WjxQE
hsLnUD/Qz9Y2xNtMqsd88KlEDm1v9T0oTmTX5k9hrNTkJOqcqaRfhnTNs/Kpl8sNFU3m4Kb00Zfm
X6uFVeftrrAh0TDLoCFSCz5YCnxO0dkLyZQPqw/LLHrvU1lRLMsiezZMIGZAdZOyAXfHPRH2Coqx
MLIybdxFUpYv1JbouFjBY6ghHRB0MsItYieMSq7291wa2hahcEshuZI1stqygp8JU9v7i/eqTNNH
KA5fgQsEvy2/a3vMSzLTOfu+MYHfplW11SNnZxgPmaKkCHfHUgRnI42O3WvE/bts22mdezFS9bve
VgBQr5YZJfs4LKO2j8TXwh/BSc/Me/yKbL2XBKgTIP090JlwcGZZjq9slJq+LM7wAztZOxFdiDcA
mJ83A99y14Q3a3u6w2wtr1F5EOUJ+9wshMuOim/AUzPpu8NuabUpPDbfP8XksCEsgtPglyMTIb0X
7fSAmBNQaTlJ7cVtOgABUnYjIuWG3aTuSomNrZOoXojhBkWBllKF1Sn63mgjXwBDolE570vUo8rD
ZAoaehbKYJkkwbrGKsLUKvbybf0omWAYojJXTyzzea14RYHQQI4ZESuXdyNjF3r1jGjQDZkgNXJ5
e/K1eCIF88MG7yh0IkfWSAmgz4kN1vJfWWKaRuPuDqOsqW7fFwSmuwasFyCS1vjzUxq5UDZHiTnL
129qlGgZ9EZfccU93+eOg2sr5h1gewLO2qPBDVbmEV5A1iXyjle2EoY/RNaHf32bzwyGzUV0cNrq
9VQEXTw5GuPPFAXUuKW9NH1hdqlCoqz6w0tl/i93m4U02f+Y2y0EBiclh/46lGlhkauhHZJKJ3iK
ZQLabFMeC1xfMogB2X/Uf+8eKojSNOjG94mFEh5/X9M/LCHewEoYOhW+HSF3KZUQ7JPsr5rLSHKZ
9gy/3ic+9ASsLooTjhG+Bvzee+Z/sMId8hChCu9IiO0zm0/MMFr3y4MEaKM+jWdDRAabgh78lu9L
iat9U8MeWjNI3C8zdx0cdMRW+PcF+2A4u17s8rYP0XMk7RPnrUDXekQT9V4VETpHh6pGShzHCj9W
5rLet1leDC9PgJla4sfrEE8PH6AtOtQD66MkUz7muYeSiItjxeEmLVNQw8VCdfKcH5DCJrurbXt4
kgY49uD+x/1jyzXHlefXaGv+5PS+lpxFj06kQ3/egIS43Un6UYQfGWgsNOHS9OiGN0SLoos4Wx5s
xxwsyztQiaEhrdscT3Nwbd6BrOwpUAlFRgy3TU8Wc9Nh/8XkmOQvmwk/FIX8nSOjqaOsCSwOPm02
zUD8bgJ4ivxlQCSEEordJrdqXiAckCx5dvrVFmS63yg90/XGFlwGOXjp52RThtc3AboQkgJJmbmL
Ai+QQ8bAyL648sda1v1SlZgpNFQ+M1AURvJLR10n37fnUWLFflDWYuRsDFAkjoQndSUdgdJEtj97
tm/ec5KKepMT4WRa1SC11VOmKxO7M4fbxUge/yiuP6bYXL2yQ7KLjyziW7mymeASvWVmZDkBtf+N
5WBF/JS7Ig3hq4L2vf5Xi7el4n1S2LOd6gCO5JPWHZtND7IziFUkJats47Oav2oyU6kl2/fiB/dN
TTeLRCu3OwlliFzi91BPOnnqhGhqQElNGe3KRYLwlTg8KplEVBTPeS/mJ8tpBxjg1qK2IkcW02e3
Fn2K0TVk5SoaDq9gXBjlONambcwDfxFQha+PBfj1j23tm50fznA98lR9Sl6RiHFhgFpOnf6Rz6iM
Y2i3jtMj0hdPcnDR0J1oaQjyOblKd12qOxSvrd93s/TzfOI6haYlax4utOwwkh23va8dRwghCYql
kyd9M+XxW9cmKQNOMMJmxvmOPev85qAqvRBsbf2Sf62wroY2aaRDKSsoIXU/1nOLdVltD6s+J9zh
OsyIRn6trtHIXyzyFiWsvdyrJTcXecCTvNJuukHOS3U0Jg4eDgVXwmlhrz+blpmXt/3Wzy13pTkE
ofQgHcPb0wpw5niICvhmselLNi/wv/5sFYXQBVHA6+nEpdu3nGJo3FQPl/jqp6IiPq/Tnh/hdK/0
Ob/CXfBRdISYIJzqCCaPyLT7SSqsQvuhMl1gVssWl9VxzJE1igDTHlSEdOwUD2xTqCH8LQ0Z6LhV
SiLRPDV6OzwyctDSdQg9OIrUe0YpUMFgUR9q/Gd6SZRGpAigGgE7DCp8q9kA/tqof0lbtw5T8Rxb
Fk/R1a0UZi92f+Tdlszy4+qvKg301DBt9GFU17fGpIIu2NQlZ4XANb9GFwv4iVKwpR/ef6KFE2Ae
S5X7rB8LGf+WkLYtWXBtAM+hnzr6pnPsYHurmXEwjfiaAsLmRrs2kPyK0qOuG8mMKVR7RiMQlby+
+adz9wZlaLmNwpf6E/Gs2Yjw4kd+wTcTeryR1BzVDB0Vn7ZLbZIIuWa/SzktBaTalAiak4u6sVCU
tH3wTPqllX7zIWeMB6ZWIZdxp6EqmolozTovC6qPWOciS8rcJ4BOWhaJIIQUg4DfYBINnFwKZ2H5
gDWEvWYIbRb6LxfXLxPU+W7BJIxAunNfEFFuz0XOi9kqsSOQEAPRfEOj4hJlH7OOZ8n47EB0RwXB
eTF0iYGLvkiwOGYWzTNDYLnv/B6A2gVzaU0M3xb32fB4sOiwJLbPEVq14kZhqYxNx6T/NxiXTXvH
34rd/0Pc+SCQYekmWZyCZ3M5KfPWH7yPFgus7eDbhDmdZ4LK1a93hRATBhJh8JTK2vTEcbGSmlfJ
tajY/RhxHdBGzisZlGxYwPzcZkLMbz+FveYLP6d8F18Jrf8kDcedOsVuPuVt5ZVSjcKmG9bY9/MD
hM+JtdTEz8J0L81N8VKDb3I8ZStThuh7UsOk3pNxpPPOTp5d81nxGsbT8qxiIgrNUCUXtwTII305
l6GtDgYy8TpUT03Rbk4XNsmxGLfx6Ot0OioZ4p2o+3wiEZZTfz1i6p89mnMDkzJ/beTbTf9Gh7ZP
Q43sj1Y2Gnh+XZVOCUQYddffTeYECM82u3Rds/x4M2HIK5euucwql2TL/0L+/12kzP4pl/uqiSBS
7GrnFs//GtWs6XBvDPf3X8ovVi2LayGn3LqM94+kAV2p+8FpKvc+geRuGy2mQQMSkmHb7dJYD7FC
uGUXkQwmMmz7+x9QoZyPM56ptgpwjGA5pUCR/HvxVesgQISry4QEM7D4dFtNKp/lzOqIGLdole2s
iaViwqGO9DFTY2+ZQXnodyGYbU5yIgju/GByuBR3iHBcyDdhA23Zdx73zWsBcOzIK/samWC7m6Eg
mu5EfhQTp8QxaPMJSDQp9Q/j2I4/BHBhCRS0OXvxC7aVoNktdVz3cuBuP5Hh5lnpD8oKGcOVnM8j
+0Vb0r5YuMKfaX3I0Xi9PqsPwvizploGcYFgdUz+vIbFIBr6BvUeusQUd+1iyqQjjzpy8vLVsa1D
2bFiKrcEmj542VfwUx6owW2XlI3pwLObhJh7VX/jdbxuM4U1ARwzQli/gvUyDdesnqsZWYSAwYYj
HeFESC3FFXc7IDhxxrG2EkMyogISV+/O+PJqSy9rfEXY8n6pdYzdGIWDDwppjRzpWbZKpmiWhjtz
BLu3ORs5cgwilzRH6qjK1T7vtnuXy6ziABYWub4oofJfk2tR9oluYsLV/5s6ttZBH0roaWfhZ8W8
VdrZ6q3i7xjwSx+vwrvXNGcc7RAPlBiNwoKDw0EuhqqZU28LccXKmCfgRQkfVXr1QBu8tg8xFseJ
IYeaeQFo7xMTTDK2rpijRxMFP9Y6CWrlJRG73apHves1sp3W5CfwbiL7hx/oaD+TdLS+hz5RJWvD
Qga9s1+WEsnRM8FOSWwZls1d0kg34VKnrIsBPK/yUXoAuCSMBezrD7ZKI15p5TR0MPyEhgrmu+Ja
uSR/A5/Brln352elrQ07PnOpWNCjI0y6tzUJPgOL4Ldojs34nwQFM3P8pSTNEn58sYBQitruZdwq
CSYJD93eIU2E73xbR5e78zRymBXxIO5L9zKTIX7+UJHdy7eWO612qCrrCI4pY0waPFBZc9IWeqVE
dkA4zYGSp+YW2+0vNg60X6pNt4LO8PfvI1BXbLXpRgPluSyunGBxI9OZOT9dmQLaE8UXnsavVoPQ
w6JlqqlrfBMyCuWSQFdcr+DerKQDJgziHOrRN9x0cyePiiTAs02Dw3nJVXf3PJhbOMpYQx3k58CV
ECASkx/UnIl+DJpygJsm5fW2vp55Usjb6G2G+22CvV/VhSNSi+6tD1ZJsJDLLmUlD76xQ6+8GvQz
7MezAxrI7iRaNR8cx8htogMPRxzCZv+cSn0/XnneHKlt9C/1Iz0ODGSXvXeg6AlVVrB0WpG2sCCv
/Y7A9yLHIHUQIHe5Bq8BiimGv4vrImI57H9pxCKjd9fzOoFPaY70IH3Bsyn5vdUc0GpKUM4ZPrxJ
2GGtS63DgGDMlZz/uEGd71JXkWnRbldnDPj/YmHksGAcMrLnlytTf+8MO0Xe92f4kK/hlCXj5TlZ
GlvEMuZutafzrGJffNbPHrtF5/pQUFK/g7CXj5SLMY+eeInW11ssGgONCXn/FB9eWalzvOfmnnqZ
75GVJSOY4NgOHoDWEpLlxgt8lM8rkV+iL0LhKJPLqJG+hI7qMJxa6P5p/qbpaf+RYHYeDCp9Jy9q
SqPSLTsaxbmFT8b8T6JtFr096hI3sYM1zjNT3W/rV4E52M5ez2W8bgghbq7YFejGY/T1ckopTCSP
4DYSNyHuPIexPUro9q2Xj31nJikStSNZG6NYMS2zOJERnEVzgRwSlLw/VOTgCmyEHjxkeYCic354
0SFEzraUpYIFsZI/PDC/CM2GoKBJwVy90QdBbIEo7zGfCBXs9HchyrnVKh3N0AWis3edYcCgWWtF
FntyqklvKGBJC0RTn4KnodJOkI81vwEGpYuSKQSYTe974SKPgXnI2usqDDAA+DfYse5ycbNYkkkC
JhwUq6J6MLXItky8RBEtPUbK7PObZwhjQZ0DYTVzW1YTEWZuU5++peRnlTO8BDWXpmpmplHQ70Bd
BfkcSGdK06TwQDT9nHz7tugjNCDNZbcwtTE0stRlK4yQmpHOwk0aatZqh9TcatP8GIV9lHYYwuCY
fr4OCYd7hyMcXJ4qb6fsdxrwzydJ+Wd8uIfa8J7phOZdF0SArzFrbf3FIdIakfQ6jOkh2XxrKlro
nPOG4OwdLeRvIjBcfzkLvfdh02fSH29b30eb3OpZVzQg+vc3OvhxdJeBaaXQ54ixE8yJ3nh+QY2r
8lp9Na3Hdees+FZEjfQPzutUNCh1AyCb6f7yNP3Ygh4pOV6lkGsR19LU3K7Q7jwI+pBhm12Z+sHX
yr6aor8f54gkWMmcNBt03KIfzqTUC4m6pF+Vl8LCeNG+QhYjSjx4jDacA5Gwr1GWuGOAnIo8aDIr
OZFJOO6pNsTv1KzDFC9BS5BgdZf7yca47H69QSCawo2WibfgwcokZGrYyWIEEabV8v8Fdk/OmdQ6
nCn6+diWbRYvCOjhdFEtE8dnIcMLLt/zZWI+9Li8VC3faGn9t086iszsRAg5N4+6MdkD2v4PFHPY
MAE+gUBecTtz07tup0ojb6DNBY2MX2wM7G56wD0vTjPKS2RulfohFxXdoT29O7fULvoc+xB66ggI
D6CHCL+WXZWUqPlurGx2nCO8LWQvgB1w+R+2G/28lIlL37EKZTqu+IawqLqLadoauhppchlSCZ5l
Q4HDijewJ3fWTRYwJBhIWcpjvDmb/5HAOSFDu1EuTxMPrb1IrmUJnZyeSuv+bOB8JhY1XjnHb6Ia
Qg0Zu76PC3eRbUHF7c1QflCPEWI+nJ10b8tTmDBLu7KgeZJ//77YdYoyXRR9a6LdlDwdQqv/pvvZ
+k3rlE1hjylPdUfSQc/YaIt96cIiKrmPbIZk3CuajoVm/OVkfPb47wa7kOq6avejlFt+ZMq9KBJr
PL7gS7NuLKnr6FR+HVUzTv/0SJs5Dx6UfjX+KHUf6lKHZ30hwmhLWr7dupkyunfnjcSJPKJb9cbI
H1Hpzr0SZftqaerUNjhcXJMbAm0SBhfHhSda4VGfBbTWBPiRQomv3u8k2ey5+Wp1khOCn/HtBhXp
9FB/MQ1vr5ZPtYjC3JeVcpbH7VAJOwhl5bgjeM1QXvk7Dh+tgePujrNY+R4uBNx6bpmo3PRiYb8Q
QLxxj8IEAeBsfdSAO6DQI9Fm3DB/ib975OiloswH9E7hglR7JFRVhjchWnvVnnbNiL5fqBlevINX
3w1sFgdst6c4JS2oALIDlwqtbdqD4mj4U3J4jvS+HEUO8GHczp8HCuZ8kJKv6vlAIP6Hy4t8N2w1
hKCNGuuphbHSxlvPQ/yhROr0IazDjK/yS9UQdPnh0nsbjZuPk58OKt8cBP4MpiX4T8T5ZSqPozXX
zOeKc7Lze7hZoPBp9CfWCNKyzJMlt+UsIzE+tDZ+Qfxny+SDk7L/h/Il5hS8NvQmaT9cWGmkzXUS
lmXaUnAEHNHd5k7UAcL7bjDm2nIPeqGx4AD5OPQw61yOKfhgAKTbiNKLDmLSg8fsKo8yqXZ+tyPd
82aaWRPORv202HHJIPIVbylsKObQZ39DYwNTS/TY0x2S0LH7mtVFk2pVV3Fju/Fh9hm0+K7ZAqBd
BOCKk40U3GvDn5IKTiXJTV4tT6sGxk7Ig3Aq1W9c1oGUYEfHzjF6bylVY2OBaGq59jtEynGpxxps
3DTI+fz7xQhL9x/nnpgNkQ7RGLoYdCevdmpWt9HW4ZFVz42/nkYDDq61/myj2pyBf4pbt5qai5b2
OKH3s3eULU3+Kbn4di22Kd9P1S4CMQxwGNxx0E4WhrZH7DyDyaPx7/WPoFZfWpUo5C6MG4pOglB0
UINWa+5t5Wje0ganZ10724sVnSScvwMqOzXFUZZeBQT7ylLsJ5SPMHY3Y+T3V9CUlELrVJPeTsnr
I4hvNs+7Pxq4yHwpZP73APN9LWgtIDjoZ8Qxd1D7qJhT1aa321QZg7kKSQwKExsKOWnaPWbpETWB
8p6n1S18J85oQoWd9MXn76DPGbjsDg+P11w/WJuBlpjawDb9woyp0TL9NyDVscayYxKpdSsLXJSU
/9CKwPc0WoWZQdtR0CwmVpqskSVMUzdVXymZMqrZgTgrKCPMR1w/OWfkUj1625nhTHQDbEYS/boS
t8op/4fpK8kxZVSjSY0FIT1qkw7PWwErW5SM9jHPBUj1zXL7uAD7Cykved5M8BM1bmQ2cX88eVhU
Y9jTp13z0gkL4sIvxrox/lZkUGzA6LJwyM77hrWAPLu/3JNJ9YNbrBJEg2gsZAV5xtcZbrV2IAcZ
1iJbWZo26hNmJiWB+2uGBW1bAQpZjyYqD9vUR14Eli58uHEzb844siGDVg//BWOUmS1HEeTPmI6b
rYVQSfnzxDD1rv6QbTv1C/iTNGR3Gg8Wa8UsQcFV/yo71cISONWw66YwLnXGGWlOUgpzOzHFyANR
mSEZWSXS8mL6ro6HKAL2DXuoth3nO4SvYlXq4Rf4zeyeeHeUjieMYOdk5Gp2YVi4ep70OBenUHaQ
+Aa+K6eZg5S1+LEA3JT9CS1FmSN5V7r4//Mk5WhX0MVje7dVpPZyrZ+CWfj6ElfyluWAcpylEOwD
XwQdm7vmxFATEp4zoqe8ma+EATODKcdqaK6839nwQR/mXYIr3pIfHGTp88rKZ3MA7bnKJofWWPj9
GjowUwW/XwMstNF5V0Opf4a37MUwhj/cQJOQfQVcOyI/mxjVD7RUchSE8TyHhuOP5S1bTr9O/SaG
o32feolSkarX66QKMAD/nfjSppA8GrC0l4tcdUkylfqzNV1Y/ZqLmPd7hRDPFxxAHTbGBnIyy/Qi
9w1RHyH+kkMayRGWTg+3lNGMca/MDMWeNudbM9NjyddTxWdoJBddAtxICzoiJfDAUfG+RFlgkbz3
GaXSjkS3WC12q+w08qqAM3q0hfRH9kEjS+JnuVharhTTwDgOIHuWvZJPeHWGxNcndR40wRJVr5iJ
2N1wHgEP3gjIGUdw9N0RJFrr6Qrj2qBwb9q4hQcRjN55nkdlKozW2+dh3lYNpZGq/LLz3K9zWzKL
ahSTbRvOjecWtPbwLzAKT62vKbJ5u8oOrfLy+2+TgnwyXPkhYvhQ4j3kN+dsy/1hMQdqEdljnJ7/
47ChFUyWV3751xWDAVuqKZz20eLzoZbGU5XY4tCh41dh91d1rK/gbmBFWNhX5dwwAqzhntLx/jQ+
JtCVL3cwdgn4y07ovwLXcpLW/DmBa8LgfBjmjXv4W0HoIGwj/F6CnuP2bGaSEhZ6jLi0cAPEeKgE
UYGg8zrZcni4kTsf9Inzd7YrK05n3cctFZt45CL3IVOwnX3gx3ztcSbToiJ+m9Cs04ce/BKO/ODJ
26mMvjmRkj1/pg/1XtDrCHxfgfWgPMlytgZhgaCk6eRpNOcxlSVnt4p0kvTxQK9+W9dk6vpk4IeA
RuppVLxnzbTpdLsxt/PZN95oEHkWdoz8pWhM5sc1BB4Fo+fUoQkDKBOSZC06Gwa++QCLhj4vcSFi
CmyGNnzDWz+zRvfgYI75cQhxFJaUFSzbS8T/Bwzqv6U9JncPSEcEzRuD0YyhA1fuRvwgxQVpaU5m
rBBmIDv6tEHDWLLtid4fOhPVx9ydS2brq9jtb59ngABkUJ0yVv0ghH8yCAsNXClw+hTJluD0v2n4
9RybTAxd421RpRVb7b8ngtuoRTXPSD5hpZJrLWU7ZeEqk/VTsu43OOsaMRx1jZr9hVsuaE2XtGG7
Rgcq3PA32WqjavGX9oVbR7y4SxjjI2kv6WvK/HJLGy4hmjQUma6InR3xGA4A+gvxGyUY7vi9lwp4
gzPUSRBhBi+DH6zf+nOPA3PEjMsRt2vA8rZQRtmdn+l7TISdrLuQ0c5KgiN65sosqVmKJbIzA3uB
bbhtJPRA5tUMgPEXKymw1JhHYkPguGRA1K1pRKVSrbLV2vElxVacdbPNjkOF8ITGVfzOoEOarjgX
gUishf8JFrbwG+Uqw45xdRKFdUq1jw56SHwAgbWm1U/TuTSKc14Bgq59s6WnLXlv6hCP0BGjByff
4seug+ADmHurCI1X7w3vchwITwPCfjU6x50EXYgyluo1HAbDuVDGGrfnrUsFZxlA4UHzAJv2ZH6Q
zfGZZ5oV2yI28m3vNTrgcztw8AUmfW6KGlEggPq+0/tJNw0wIBAgF+Afl8au2NzYOun8RveGd1XP
T09b4SsZDZ5yrMGML1BnonXIoEbZ/vdlLHSf43Y7UvS0pAJQzaqEXH9QmTLaHRvcL9rOZaRX7L8C
0xA5xdHWHXNPG97DGg7tl6Bvd3kHQThIISLN7i+xAEC1+GgHUaWMpOnHGVdSADbyNg4c3ZzK9J3e
/0boNcRcc/w2P1pB9W00qDlH3vRltdlDyFfiPaGyKtAJLXmvWeMxniLIjXamv6+HjN4ddZv/hlPL
F4puAMGJhX0qPSML7qLxunPxLjB1BshAGKAqUv+TeI8W+dr3UTf/ozh8vObKjIjj0BJjG6s74GOC
5Z+U715grscNL+zBvGPBUUvyCBUSdz9sJbZoYfg1iv3z2A2nDqH0XLsHnfLcV5x9bTm1nCfBUCSP
SY/DV03NzIAioZh3afMKrv81QxohcvWXjtgS/Bo8SkjJK9yBeiJQ3Q6/oUU89PYegAWaBu2Pcgny
wd8hNkoonrJzKvsJtRODKlWsjuKaD55Bc66+2ly1Dv0e0mG/Z3IfpxS4Mdk5D/0/pMUHC8UpDZAO
CWDeIfA+cFA3XFKpGZ0eMbbONwJRfjPjEnqOLAqEfFo7t5t6eySH4ECKUPszUkfj8b2WwH3CobzF
wWpPQyd+Xb3BWOd8lJAARNNf/n1D46twXsLbzHJYeRV9cOOwRwEeFahcXinv55VaSvi/6yXSm3BF
TMIQeQ3hBxo2X/mnIxL9TrBzUEjVmBZ2W+areT8V4ZaqtrLPC61E65r05sqa5hDPd2lehQp/uguw
tbq7aRys969RVoGeBe7QoMuxO1YTXOqa4aq1RFvIxrDjg2rj4cOoVr4JyHZ/YmIXPYLnUvVpcoOU
51QwWSMjSHueatrv1GnxyBJ367oKPLrRtmrLNf+aryKSW/+spl5ucnJGuFaMdQ7b0GL5VAtQ/Z46
vAtVBUH7+Y1oV92pb3xjR7aGs5DNrGjwXqzz3A2IkcVNmRHoebcUBmRMqutECnL77V41txNYm4ZI
w/2v2HfExOfVyzv9dOSZzaCwxsKXAan8h/O1pMCIyQ9XO4SjuciphLlqeSMGiHZXiNyrrDlwM8tc
cNVwnFm5TpgVwGnihfHYrL5c0kHrj2A0XZjqoWIAXbWh3Hz6n5ktHhVpvv4ws2Oe/w6AAgdoQ1pk
fntC+jADgtEixBOsRrymJiaLTG4LUsO/DPPSli7jNy+NM+d8gIQz4q9lupC/aGM3dU6rP71bMcaL
mZ7sc/0BDigmFmG6N1h1B35naXf6bwHTzb1KPNjol6G60RBjPDtcG4XlUJqUIvqrqtjXFicuZlWQ
9/t/eh1tv/6/cmoWOzQrs5P8ffVDhUTjl9agYZ3o63DLO/88yKaPo8AO6F5sKM3Dq+CexsFbayNt
ONrqUTIvPy5xgjDgLSeP911pUdO1CoSXQAyWHRhkww/tvMTaTsBwdHZ8paiQM87VHl/oxXfeKEhQ
j/QNMGvIVaSv6r/Qs99uyUE3zN2xMYl1l96JOSdvQSQ57PM4jluITiT2QdlvW4G0slS2bmLYzaiC
6ie1TH4FlTSv4qq6uA6QzjTg5J8diJ2HcyK/0rKG3KbvZ3unHKxRTy8JubyH7IHfhkldw54q5+D6
kxDq5LXB0C1Cbw5B6CtA3wH4VqqbJmc/2DiizHjkUby9e21AUHDDLomqi8o8A11k57TYCY318/a3
8zeLHPb8XP1gM6ttxRomw+AiNLUxV5c+r89EIYKD3Xq66KX5/FjLE14vH8uEEwKi6RGiISGfWE84
hriVLps+7K2EUq2mV99+7f6MRfuih6xiPPe9ntLOehTNFaFDxkM0nQDBuTK8ykUuAc63xuOi3pmf
MZPhHY4G2sFGN6xk7MRWGluh6yfvlEqf1Qcqc6nrzqZiBnF1qaS9JAKLxG1lqnimhAjpkNr1f7Zb
t1O3zSpG54Hm5uXy+WCp3WfFiM/T0zGeZnI9gKSOPgFhmLx+pHFdBrK/QA6Mqujpkg6oBPpKjOR+
hmNC7vwce2QX+ycQDDpJymE0gKFMp1XTEgjN7z3WIY7iDAqZjF1QdZmdegFcZdj9Q3IilQSYSurr
R9X7Nz9k18wlbdYk7/GZBVKuk54+ycx53CBWeX2TwBJwGii61NHUEO1xYZzHzm4AGXmXMOlyPs1h
bDffTmMWWy914rg9wH4onPjjJHJzogqKlACxVrMfC7WxhAtyyOtvn2fI9MS8oizU9Y0oDwqPzZsI
psdOEXGkMtMcfIPx0i3Q6HF97b99d9i0oeTExWKfmSeKN//uQ++kafm30qIr+3uBrnIkZ8eyUhJd
ZbJ9EEFxZyxT+/hW8oAUPkZxhYYY0SDvfUHs64Vs2tJ+6OtlHUnvY/EuMRLUWrr/j6+2ea34lCF4
T5wf5B2fgOdvvQ0L8nDNU8aTSJngaVb8AGeEb2Y0r6D2P78w1Dh3T9A4hulfP44qxdaB7V58sqqn
/cnTmptx2AZRcynNnJftap/FYhNnTqeNKx6B2KcDaRfEwFxFZcul6o8YChH8P3xe26qOvBjhqJ4F
0vo7ogw+uAcEl8359g+zPdVy7BO2GNIPdganzkWMK8H2N/RR15LQZylhL3SzNLocNn+v3vOM+bic
P4twmqJlsp3zU9g/l7eBkVTOuCieUe1zIdNCYol5kdg2FgYPHOvPevX0XUFb/xyqgBQ3e1EfFtEs
JmYf3byly0KGLgrIKxx+nEmMpC3zKoShnAAbR/LLdVQ2dJ4ukaxdUpZeWEdQxraFCS27EEx1rl5s
i2J2lo5Pj1Sz1x9AJ45NwT6hHzjsT7tjXk4FPg7SG0kE12fcIjTD0+MEeTMb/T/a/1HRe6Pq+zXG
vpXf4gLYQHfFSk/KH14d5Y3D0xlaFysNS9BNG6Jza6G9cJjUzmKKL/UiVpIiEEWic5r5vD4la8vl
e8KU0McoW4KCBumE5oc4Gkk9XmsWHY8ATAVRvqE9jQDRqmS4l2AwRBGzTr1Ts4MHFRM3PtQFpij0
N1tMLM2LHQV1HkKRC8V0c5uT0YaRKCgxfRh6RN1eualRBiZ9TgSwhAPTq6RhdoudGpq5xygMwHaE
3GRr5e5B4Bm0vxU6vf7XfZ/b2jYuHvByad2WWY2PU0ZDsyRGVDiqtcDHKFovufmY8tVUZR9G30Tb
+HwQjLS2/lypq+tJHayPAMjg7if3jeXw3EEr8zAWT6SGvq2MkNoq+zgfQo3546DBbzsrmrFtCIEk
q5BjFxsDWn4QlSnq6NZVlV9j4xBNpM9Q72htsPx78TrbJjm6KNulgiGvPXQ/7i5rEsX7xqxYpFAY
jI3UunAXLllUR1TLLmy58RhMkut0Ew1DeIn43kAkFgEkBAMy9lLhvSGDMEUsBk4LdmlLDFbLye2t
ZRYXcP8HuGMGNJW6wFSkAND3sUcuy9Y4elSGJyO13VFCo+6huEaQgt4iX2T7+kbT2/2rPaKjISrL
PoyZPm9lIKDjLY9+ThXC4ZL66wv67JUklFO7KQXd3FGkASs0ZX9wh8d46wYfvrO46DByoyuRLaXm
Vkm6GE/NYDJrzNxevqRab59j2OeM/1NTXda86os4GndFMCxuyP0In9t44GusBZ/Na7UmgEBvUAm6
B4A1LwDNjEpCNQoVQJ6DyL2wpq4kvTrzcreLSklP8l91nUrrscYMxGo8tJu5wNaaN/WL1BakiWzv
X01prcBCXYEnhwkk0emanJOB+LKrDdvAZkgHbrwndDvTLNFmiTmZOdhvHw2Z53N9aQVxXVUW45xq
0Ile107lOp2WIl9nNNPb+R8W5lLA6o/yNaKHJ7gYfOBJPxe+0GVcinrFWJF8K2fDC12mLJlFbMuA
kWdjruhM+CHAxWf5Ibybym73DrvEQlyQMTSczJZ/FWZBCqC3CAQsrej23UFIDcFpTGvJ2/PQlyFg
qSKFgRgu5u2w/QqSmm1KcfbWcthA4Wu84dlsMhOEyNYIpJ6k4oNLuxS8VfDsOVzP1GURXc+yvCgL
yl77KFY6GOPe7m37Dw+i8TQlSzbj7K0oCFLsPdm7wI4xhVLnVM0lHdw/6mHdfBzM1MuS24f3nThj
r8tRepfZ8zBXzQIDeoQbQ3YViwREMR/2N1ED/9N0Q9clymX1ZJcaq6i4Rt87zIQnxRKjz68Fd/Zg
H9QcBmEBFUWcAnCaqyxdB/dtw5Pj2cL7j2kDs4djQb/UxIoJ0IIGDelzMPXYau3LEw6X31FG4pxU
XcmzrDSqJVzFCb448KjmzErI+KD/jPJuwlI7Hwx6Cj6NkJLNN6roQmH0qTEPVajlI/wm6tvK+JEu
xZkNk8N8tMW3rg8LlKQBIlk4COp832jtsYSQIGoNqkFM1QBB1J9YGpPlN+9ADoYPAB+S/4cfxJlL
Enx4aFdZQqVCHs4sbsB6Ylw9RIl8cMtmG5TT3a7rs5cLTl8s4rxxyLWFkrXK7qej9zDqwtsEKdG+
HX6xwbR9xoRiCh0IIMmctMjBnABvTI51lxqsqopHvae13v1QNUtS1Wy9/eRes17q1pCF9MuWKuP3
PExBcm6C3JdebC/iYhKgzF5G4lGrOvZdzLxFYiCdbOA/T74XkK8r9vzWl3RwFm2WlgBw+Qt7KCiH
Mv+meoXSl/Q0dXekSWILkND+RwX8fEW0U5LksAg8XsK44TX4Juz3q1OXOz6XSRKmnEruMOcboLR9
IFH/Mhiu4/wFeMYIewBHWJv9+vFh8qkLBaDY87CgvdcWEpLbRxNa7ERrofb33DMIpluMl+0sizzb
65EB0jaw+gUOIqFybrcPjv4Ro5oMFQve9BxiTCX382aE1RVVzrgBqatSUhup15uldeKZCkRCFyMf
bfYtSRVXWvW3cBhaFikwntgkcKcXg/jBBZtZLaNaaIDiFmf5V9AdlqeIDpdkrB9haaYxOGcAsbwK
mD37eThz83xtZNPo6BU29oXSN/Cj54cakJzYll8jEEuFtgAgGszTOeqnul3lP2GKAUYvbZd00kmq
UHgquokTY0gbbeOq5DZUIGe+X773qwdq3pq/r2736gCzFe/R/S1wRcpZD9zYgOG7jtyg+e0FMN0z
Z0zPHqbhwzwgqmXbNyn+QaYvmpvWhHVxLC6RSni9kbBgG0oLn8VH12PdmI0Ta5g9xUx7Lta8gLH2
g+lzwcfD2AVr/0QlrmJJ3QECOZH6Df7/kmdCsAJxku0wADKHDT55dZnLtV/QjfN5XP5b8dnU+xI2
HbZQ4CmezetCQOtxbqLKoqChLGf4bWR3+5W5eMHsTc6HnafMVF6h5rVFE44oRjnn+ydKE5PKpMVQ
rLmydLZfedxkMiBOlG3DWciuV88ugJ3jzfgglWlHlABsyPNpD/5NVvsX1FT3wyiCFUgf7bNZNs4J
xnNCab6Iy/kuwOsvFWGI1vLSVzg6vPeska7QKqyRO/9hDxYhLXPt0zcBXCeCO9jK7cZmCulxutIz
sWhuIcGNzSGXZZ/E9n/xRZGL5l3kDNJ5VaJD//s93kuQKlddV8SBi5393nPQHTQvahUTyk0whM7N
CS67yXbvT6Pb+rV3E1ywtJPyF9ap/OR/lkFQYkbCB67Tc4yqDDzJVL3lA+4mRG91xhUXIgFJRZg4
EIvSXxttFXbGZyQ17G3H4z92FXo/YENq+16h5HiAl+mZyFkZ+Vvb39gbWP5u9UTdtz1JIDnjnQf4
zubbTqhIn94og1o3AsLAgHfCD/nBvgvdiWOM6cSw8wQWl89M/9NkPhDdhuRpnpXpTEzG2oUfr6PE
u1Y1L46H+kiCRMCYWfNheuEWWrzQIbaV40m2YaoBji9yf7XGFZHgwRWpp6KahIm8xTHQF7WwpsjM
602lL95Ss7M+8Y3v9v/8TYzzqq9YZebeDrDPO7CjmLJyDEvZCYco68czcHPjLZbdohqzqci90gyT
CjnHJhl1FhGggfXQZuDp9kmOHDYWYK8MVnyE5841Cm5BRJ28Mr6BYP8bwlpE8IfPQ7LjwyWPkVts
fU0hRtluKRNLZcTehpNqI6s2wk+W2h2rpPkYWWkmdtH3BrzOVr3KHwB5kb8SARyhDZv8KT0uvmj7
eWvlfL7w+h4+a2wBaV0gLUEV+GVcsTSAmNXMuxWdA98ms0n639yb66MwU5cd0G3BKSE3i4ji/kKm
jh+a5gRUPttvOhR957klFDGLuKwSLSZ/QS6N4unQSYpl1hbAL6pkooiLcglK3Nb4uRt596uQEJp7
eM8rbhQzlZErHzPGAiskpskLmOi5ZzURdDFyaJLBqCD9y1khIZhlVqr37aJnJMTJj1h+lJW96m1y
mf/0IEzRqeGm6b5iEIUqc1oYOLxhiWB0lXu+qbsI0Iypf6rEvojmVO+rd1VaAX74uP7M0wsVXJ2B
grum+QWAylgK1k0OOl8AKk4egvCeHs/XHuI/rSMQEhg3Dcb/hqaU6QRzfsKIqC5JrWaQqou2m8ef
58Jc2juXIsfSWzsoPZOz+gXrcnRjQx5Rax2eVeDaWA13LJL4c0R0PU4Psqznpwnzc7oqmQR8XPFV
lZsi9WVeG8+TOkBE/fTVdVFEiP7xOkvgYb7VBuYZgdidTRpEdd9mNdvf2Xhib0M7+aQv3+2NbW9l
IB/VCfKnG++xhfq1+eLTJn4armicZ6c7D0qoSi6aN1bXzN8O/LK9OwL1HxSSxaK1w/FFUkGoYfme
Tvpd/dFISyIzOy/nzqDv3oOeytwfiiYDxnn+e39riF5U8Y1UzABza9hnpUhlz8qr99a7CaGDPzSe
iE2rAmYgcq/PzFBbLOjtJhiXq6KTASBAyarZPA4G+W4d92958gOLAuT4NiHX6tjsOGmqh7s+g5Ez
QpMMq3vJxUWwmFUdpkKn3jitSMJmvH3TtRMFMS9m6Zhjo4OMwowsfLNhlcNG5chvVJQn+UuBwsuG
tgiX/h8sHAPUnJgD3jJN7YT0MPayHX8zwDUPGMxfq/l6NbSYxcwYRtYkGfQigBntP7lR9rXuaFhK
49WXlh6HABT1BsHO+As/wJfJrdrNzE/51u9UPQah+Sx8Wi0oV7MaAn+AMAomlSwZRmIwrtTJi7On
ntuarAZMzvFPkU2EQFpWEnqtYvTew7vJ6NWSWXUvIphJG0A1jleM+M69TOV5u9W14oj4uXCVteOC
eQJfKygXmX2obZA7LX5qIkpqaubRmE0Nkg72M2JRvJ7jAttLkSxeqEItaCYeuiImvo6T59RdIRSY
EYGpmoZUyLWdw6CqnHNcX0Zqmavx+7vYKgsM48sZRxTp0JYJxIcAGAHdeNNsX6oIoSAmBvLl715l
d64iTPetIYBwmAe9e56W3p3XddvFMKJYLFiezVA7b74nhEXGOVWrUDSgC+2fsBq5qzXWYgpREn75
cnQ2WqInHRiEKLaH501dk0irh+kGBI4dk4Qs4SZdVWUTwRS8u+2bTBPmoon1wxGrmqUzj9jNed/N
tXxwQP4fmnyF72/77wuhUkBIBZ+vD0jL5MC2J5NfJ0uR4oSrAASjCoaMDOx07hLI2/BrZ/yL1DWT
ZzLKz70EeTkjAZpNJNwyZNCgvUx4Axrxds+EMyh4xYoBEUXs/rrIwX2Y4GFAOiaLoMvFDVJ0LJkw
nvszgKJyfjpSyePxhbk2ZY6S1PY6Ov2AIFMjm/GVtcguh6/OFaoZdciS9TdOXFiEduiNbXJpp6F8
ncUGxzqqezfvQt/KA6Bg75AIehlZVPl058eziB39hihXFRak0vPdDCSm0lga68SmOp1Im4UcbRBT
e0oz1C2gQYHBLyfMwxhRMygsa7er49WGZIGCNRZTj9U8nQig3WEVZL7sV4sGgXrVSRBVb9iTXvAT
W35h8fqEm2eCdNh6+yshmqYrQsSpAA4KFejbhOiFtcPKlcma/pfy4IVcxCqeuwFzxLET7SN//f2j
ldN+nj2x0BsLqAXszpNZKgVA/S1KRgq8PyQUHU3nR2NnAMYO/wgQrrrduPj1Ozd7r74Az8EtaH5v
WsVMzRQTDyONcEd7xI6+V+YdUb1UQmNFBj1Zu1z9fLob4bS/rnkIaysXgP4juvl784XC73RPVYxi
uk/NgyfAfeTD4pLhWWR6dbWyCrmIh8O0O3R20s8oYULnU1UVBfsfomh5GXclZZ6ZqtStVt+68F9g
+d6UauhzqNLAt9+48c+dQIOLmEYpm8O8Ixhvfc5F8uSd15O5KuX4J5kR9h5ykyeuCwnXbucjLQ22
4rCBPDP+DtTuJuuDehQrqbNauRlMmL2BMPLrMzn41TgRcrHs1zvqnUbC0kWIXhm0g1ZQXhum/JAY
Xq2qKuZDUWMCEY6sOnLczppRztV1N+03/sG6TpPqmAxGYi1edXTz6XMn3ilvX38gVgQEFJIlvedk
iXDcwbHqWxnqeEIqP5O1PDxHIr49mXesd/GUxhllsTLumrrObRMzG4O3qCEQ1jXSMl3a6sWlPAqT
uon5RPrmz9O0OGu6fJybIs1DrnQMwf4kq4wMsBYtuZGE/L6mfzbZECf08EluSOI7TIEKY4EGdQz2
l0yJHNXylnJhD1wYHaZul/TTS6b8DLMAAQg2D5OaPlAhCirc+hdPuRSFRPeM3yYBlp8iKHTO2vr7
uHcqdZQYnYn/l73V2HyQ1wB8inIuC4YsseZEGkaPtP0IsEiFAB/kzzH6Ze2fiT57NSsh74MyPyK+
yno07JReXyLlaWWusAQBDfswpIdFUlSsmQXRVOUvWzRmjdCW4Ck3QZitx2f7GVtFGw2ON4Twqa36
BtZ3lnrmSGaC8KRvneSkyqgPhOH+/+LizhnMSLOI9Yz/VE84n/zqj4PbMW094votKzl4TbRRyZVi
oXhRirVqEhrDUJFFfSkhqP31RFuUFaa2jLqFcWfLHzdQxI4cVkYkQN6JuwQZXqF4nOrCMhhioRcv
twkcXAauBjMi8a3/oRfAAlziarYiRKOR1bfh2h8x4vEf8LxiPP6GMtIwOlS2igNYDOMCSWbHhFoH
oW6prdBSJ15mRxjVZ/4tT4yJ1aBCVe2q+ED6b6A3/oOq7n4PahcBuRpc7LjUAe1fQaEeveHlTsaX
wdOON0ZfQEEqVGOEW4qookUNOlzFKVf+PksoJUuQtN2j7cz3mxHSLejh/j3XfkoTKnnYAnfPSj4l
3NzYo038kra2hX3hGACT7g+om9xml8ynuwfZC+GB0ZyYTBNYe51Oy4pHaAkJolDB8zUabwXUFkXR
YB9jKg+o08LzXGa2uLbT/kbBosa7inGjXXyyGE5NIl/Zoujot0jlR8drstm7NUnbPOlQOKWew3ag
oxH+InQT1w3M451NApRHdt8iVDcG00ePN4Vmm+Pj4L7x1ZxhxzRMP+7qlPBHnsamI5/2vox40uo4
qsvUJ/ST4oF3VyqHAo3kXMnUPgRNQ2DoKKs9NIpmven8m3IK4V9M2Fb405wFRAmkpkVow1wAu74g
xqvsEIafyQkjdXiM8CPHmOfwmmLVDUZAaq7RD9m/bX5PekNtlFs7OKggs2P/9iTc+u9UUazY+X0e
Vkx9UhmdlEsy8mD8xE9ueO2J6Ou6+jYt8o9gjmV7uPXfjfjrkH780Ob3Uah/kH4ylJt4UKoCsvBv
NDk0kQJinR7CUz7HXSYBDND2Kl308IXTWcjo3dsSp8eo/bTkE/cWcPWUkRFIhJKt93oADC7B9WpO
hu8RyQscOqRnAYVHm9WwAbsk75Ow8uqlAKfPeOHGYiugzZBluJo1aPKX+dLMc5IAml7CMFtv3O2D
fNukgFlyNZtAe+wa+sERZ7Byo+OQo7GURvlKX28uBPluOGiXmqh4SmFSaCDAJzHbx9wycpCnIpnI
h4VZYzwwe/7rOj7qH5+vSgLwp9VCC1/zZm6zpW6DK5Ii39Q1UzwMBlAu80DCmTJsJqJHpDr71hwM
Phn4yRLcnfuQuWgxuzZe0JOw6Ij0ugustpZ//mABpG4hPAKrl9mWDM5gvd0l+Po5ljrsoLcIdS6m
qeHSCEh16DRtOonrT3IJKPoFAHaiTLarswf48VZwaNzrpXKoZEXzpbMj1C/i4cjZgEGXk6L6wt8r
t1kKJBrR2MCHBMnai8YK5FIGwE8dln+fIeWwHCu4mgR+PUFo+8pTxAZ98I+vQWDazNebIIYO74Wf
9uf2TsjR0H1BW5HzCJfXDxkse5P0DaNPky7KwU3HFxclJ4umo1dzXvGTV7fDSkYOMhKbApjkaS4R
QeUKz3x/a7hiA4bktfqtuSZnee+3yKH7L10zR7tfr0YuGIrJn+1Sjs49elXIi15MjM7Qr6nQ+UZX
M7BUGTmnkoGYY0jyKuZhYTv0GDnuk4huWrpeaUyf5FXPkrCeQ69N66gp+UrrlM3kN+nx6QSOTHKE
5txJWSMzj2QOI+PdnWA5yFuZKTZIE1rIyllgiXNSBYel0L5R/N+560yGSWksE0J0WqA/ssbZtoZv
6LD8eiYgnmEGfR7io3aNdPPLIRAkKhMKdOLa0P/Z4ROiAGVIPlWIS8SK5zzBfX7AuIHbjX32C+oj
iKajUz0GzASIMsVhde2sCA0uAT5nghfqndsCodoElTf4r5HVU8UbIuQZUeTa9C9XVrSzfrvwynJn
kGUah2Ar27e1ki3VKiaWJgmbde4XYdmVRKZKy8NGOZ2p1KmHg+50683vgKk2Gwrax320wC/Z95GD
A/gx/cJPC6T35V08mxAvEOjiPUmgLfTKqOTG841XVi749hao7mSq0RE1HwgjVpeWB/5o8YbZQeJH
m+ZIXQggwTyok475939JNxrzj9APr3Grtfqyjv6nN3EiWg1ti9ZkAubPAkpnC75T9prVUOr3yf8d
Xddh37nmHO0zz5nwAbiqIqBURCtKbVWfbiLSyq4i1G/Aa/RiJNMCzZ3DQA2naXgBejFmodbAzslx
M1Wfb8/a5uz5nQbgmDCqgcJzhlMbGN8Vu8t1WPdFFQvIr6IXYmotRQtwzOKq6oQicYHTvVR+OOxB
iEcbxKQtcx0ztGcOyxo286DoSuvJOmlvbawpgJFca5KzwGQQTppZwS9eZgkulHM9CAoZfzTU7Iyl
Z6aR25ctX4d6s/eQ7rpQqvxACwOKcLEEIynagNJMEPBwVfaydINLjR2uI9v+xBBuUR9NI+s8Ilde
axuE6knA8sRuzbrgAvYQXmzrD3TiNwM3/BSAKS9HBO4wUaQEINemfHHR11eZvr3xO+55dhNdOtYb
72lmv4HparaeDE9S6JqWtXVLLPsJR+qlIO3QpXi7SszWdTIlD9CBk6yoyIFv2MiQ4l8Lyn7B0P0h
yeYCdvsaAlQWbyPxmnWgq3CScjGSoSq/C7tc/Xu2SQCqdfvZ1HT4bcVG0U5GkVyffflo1M87kzPd
xTdWFgc+fF9FmhPqPL+KWkMaw//2r+TIS8br5+L/5VZ0XeDvqQ2zpj/XXtFXeBkBuNQpM80c2oyv
XYtYGyXlMs6GIkbDm5q0YqPJ6sEanoRwzFRq/fUOGOIK+wsA2ad9gVTtvn223nGSnIWAJ+mHgsRd
fTIaixKBtnqJIgfASpio3VLqDN+Ltx7KmULAGm1hQnNfg1VoBOFeM0eFCUQydcMqNT7WoJWNP/4h
3ldnKk2DBN0Ka1ogIGvtYTXWAWho7MwumoA2ctFlVFqCDvOxd4+Gxm1hx4M5/WfopNew3WLVmUkp
KDAWxYALyoRIBhh8wr2zweVwLBf0TBVi5qTByxtYHfLQdmPEhv584opBUpP3TiQiORSQkHn3UGiK
7zGMVV66Dhe028jb9WMwTJ5fOSCFaXEzaoCQKjMZOtlqul9Q1m9qcXQkWbR5RYugCN+WwrAbO6lR
/l2jITLEVZvQ8lF5qz+9wElesfHTqo8R0kKV88AlKUyagmQA3HUNjpRAcrftakTN6OAkU3aEaBOg
6qPMzUV1DOHceGFi98MDX6b49LpR+J1k12oQiuMtOzvxeJ1T84G6JueTLEUoSxQ2B3Scd7C4eyy3
xn+mjXWJzTzhgi8gBwok/LPSNLEw6P8XHb7bJUMMvZvrkyOAhOeXqZg+NA8pa+WFEfZ1qtThUp1I
4CPPNR1CcFNGRowQUPSm/PKunNUC+8SNFThDNr1DORAjTVZM5vUUemtsEbS6iOlwgGTNkOU03J4j
MXie0AgftbtM0yGOyV7ToIzFWjS6UtaIj3B8r1ROfkTS0nYbKaB4DAPM+yRDUfRpxWzKdlecwyTE
3AJwsIUtbgMG8eDsH0aDHkQU6k9/HTlFeI9sga5lLjN88SyX6sGKm4pYjMD4XZF9GBpY5h3ckspL
IrTl7PcCudMJVaQxAViSdOMOu6BrULdq2aw8Tjh3P9NMkhePa9wFuIgEqoYibh9cMQtk/mhV50E4
kbTDArxNkI5dpxUcm15H8NjswhxyPntDs/zTZr/33jhZnm+vU2lwhD4RGMdZ0+sFJoSyXxnJTtGx
zpdXKrv7atW18FKdgD/RGzwwc27nPoxulQfMX+vixbFbbPR/oRpUnpGsR9L/6QHrZ5r2DBYHwjm8
wyR5TF00JGHd7oduvbx+fBEcffYAT9Lcrxb4gda+k90juvEGl1VKE64AOIK5J0ShVy3K5p0BVKCg
uMMZ02kgbdlF9F3UZKgJuzJNwKnGHFGNbVhSD4LwACZnwXwyB1fXxEBHPtNWCT9rWjbZDiZBo2eu
lawG+XiyfxGLhEBbfkKVkcn8h3h2+mckEg2fbt7y57RGJbbB2/qYrgVjhBOOJvPrJZ/YTBXMEK8Y
1WS1l/27VznDlfggOT9IcGwms580ElRg2h5W8vUnXSS1ncapjK5bB3N5bkGu4bQmNS9ajXgvi+nG
OJBLF4k+RsYEnuEhEx6TZOPx+uuhcxO/Ek+mkTENfkrUPvBeguPWET30AXEp6OUSMZqWs9FiOuPd
/FGS0wgt1m23SO7rjvO34zMiCFBqy0CThWekW3LxHL6crCyvanFOepvMFJRASpowEPedmTbN/wpE
IFyjhaXaESX0YAgkEDQHg3oJgJw5Xnkzp756Nd3PDKA3AwduB0NBhkN36RE3ZS1lkTLl4HMpCip2
y95/upV7Q/9B39WvrUsGG1kJ13rzEwjI5QgFaWvG6wIneN+L5Tgm0lHe8qPccJNP4bnhhZ030c/K
29XFckQ/0CqtytAuoVYen0TuqCW/1pQXNAe0fmrXcDGC0QfCrBOuCGBrkO5oArTF9zuu7FpiPpZ+
DsnE8NL8VSI0C1GdZqoioLG1aHzp4vfWA4CLj6ExxW8bZYVDQ2guPyYa3LjVlcBT7BCD+RnYoq1G
P4LnUjZ2CkEy6CR4u+tBhX43ZPBeMOJbLwtwNzBYuiaKwH7zEE1ncPtIGzhxe7jBOU/wr3/8YSa5
S6QWjyADh1Ukbc4jE8q2zLzrSs//DFRu2bdrAlpiLlxnqnN+Hcl7YfxuBwmw/eR/5urKXsfS2v99
KBmZCrt3XTq+WdaiaNbhhpinimUJGZXcQDcBpmia+jEnhv41gDXRPm6WwmXTeYcaR4Cl2H0FWHQQ
nhfM7UTWltHfAyKnleTxAS4qDOI7OYeyx1+e+Ikh2uHe2IWF11rR+IVYGWMcOWTbfD6/f/WAW40H
hTh81QCF+7sXpRVoIQ0uQvgH1eozOwFYCr4Tr5Xqkg943YbUN0qJ7fSw9gr7Wcol82rB3efWTKgk
COoGEJVKmBz6wfQSk2Ir3fP0II0KI5rOgo2oqzFMcNyOuYzFpuGmAxSWih9SwLuKExzI/IBVgxIR
nLU00PV8bQdsYImtM4vq4ziqbLdmxVwXGD/YTzkDE8Ul5b75MCXm5/qzpoJ3MitDNrWWIYrNg6Er
QRU8TnJaNgzCuo7cA8QQ7BvybyMfCHPD/c73GaZQkLMHEbMRKhVowUIoGWa5K70NKZEa7MzDqQb8
A+qxHW/y7OPt+H+qR+oaL4j1KZ/er3jf+fzFsVG9jCP0vM9J25d11No2CS4Gg4zM7mFqOuWbocvA
kZY9vWLGGwrSuJc6hYm/oL+F4Zxn7xw1m3v2R3TnaK5QE0weSTv495hXtq8mGzVRtstlNUTjUoIV
wsyunQnK7F2zm/ozFMdCj3s1uHS4+XM1qeebhfBs+ecXDHWRl6lMgWQU9KclyNC3BHg8w0p+Tka1
9B6stAeWNRSmcv9MvL0zNlX6jD6weO4G6W2IglZbxC5GTqy2YYsa4fwgVUXjuUHaYFr4y2assvfM
nYNfRPmDwv5Xy8xpCOyn5jLOogZpdOCMQmed7qUehldsk2Ys3ijkNTO56gKf/pXNc6OH5utrMiwz
/jYfuvjafT3+UJL2MnVv7OM7q2DaEaFVxaD5ebYEnVZTWAxAvgBRc0Lq7C3FjRmwZRS+jaeJ5818
BCQXzUyrZaNZL/dwZCuod9NN7PJwSiwvTSZIywUotlRzAoJeUifXz7k/+4T68CgRwb6Sc9tqkObh
LpAIM3esgF4ONIa80dIMuJ6YHKZWl9qgRVn81S17c5fXmZ/gltX5zGuOFv06bDMiT8kQkXNtPtGv
EUus6XMTLu/YiCRVHt2yoMc2eAAapgK5Ek/HeY6L1Ea4fkvIRkJl6BkOmgg8ekp9T/HD18fh9mxx
cKzd18UhGS7lWpmfr/R752XPnTvmyiD5LbnTXH6GxcLiFt2U0w/YuxkfbCmId69xBc6TWna8vxG4
POCjmzwf7X63eZVoVz+zyAsFRVmdEVkJGCujvU4osttb3ixlOFR9OB4rh85x4biYSDJcAE0afe/R
AzmjvA7sgzoioDDKnhQM8gPDMY+MSuC62HyIUYHWRrfYBgXCLxelN9SD6LMyHGPPrAp/xMFHXQBu
3BkeKoXSqY0/Frj+xxMxgW/CGqnVf4eXcvMKOtBQ3DGrUxKyyD9ispNr0ZPUXSU/rC4ldJvmh//r
dvcGxPWA4ncGAqDc8072yoG82vBVl4NfH4Nh4iJxToCr1QtNskYVjoJzxdX9l/DiXsz0DQWsqzxo
zvSwNwhgo4HoKOn62hfvRUiVVSqtB7n31CpKUHhEGi8N7kH1b520Nke/KkRe1QlwknP5q2v2LwQs
Fs+gDm3EWuT2R9ye36SujClHcbvIaGc0V7QUTy2Rs1u398HRmQ0p965VWUUvOZ3tKflUU5edA8Iv
nl9FG5ql1bg6iEx9CHlLe4qGj8OTte+dNhufz7t7mkk9YO+/ZKvCiso+LT106rMu5YZG5YmD9MZj
C03kBi9qy7YtWDikM8Zdsx0/RrQkTmgum/NSM7Kau98M1OmiqlwW
`protect end_protected

