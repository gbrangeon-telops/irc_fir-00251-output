

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lHZAv/MVAAt3F19GG6CyO2D9ozHTHXUyHUqVqPhHJ9Up8V3v4BMtL2rZCdPHvvrLl9m3lxdPLeMd
yZjuwpNKug==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V11pDh2GdTX922gInHRdE4PGQC5LocLJP7s9hbeXjPbTiX/dPLHGusbEN2B0toY0K8U4vuWNSniM
1aH2SNR2JV5BnhJYTc5D8l2e07TnA0V6ktY1z+NOBfbsIHPai5FO4rlYQdX0gfNxjRiE4WpTGufJ
+8B9yaPmasK5qJ0hmyc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0akrUk3wQb4EqzKkib7F59nSOOeoy+q3qc0fQDYykXO49Ll/FgY0ewL69TWySlFx1Cac/+BCy6vf
iumuPLpTjOS55mFm1JTMxYzM9NsagXEQHLi1lEkcr65/dw7cjFH/RPICXrv18S5beJM408VyZvsr
NCAeZ9gbVAaeGzkHq6VNPIh/P5GGGWEK3241GOn4p1v1t2GkteaDbOSjGK7wX7a4kTfRzrAH+xYH
86BcPdOp3oyEseFdQgL0BZboHxt4zJr0bXL7Ln+oOm7kGCKk4PXPdudDDSsXKQUPtDHqr2MHJwZk
LDVjKe6pX7e2DnCF/lojAxyhWqtc4aJmRRvYWw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P2FMFi4MUNbCcmQEmOw8kkGKpCf5liEfyrVflbrNDPfCQyQhrfO1z3elwJF/eYuRk4Q8ng49IhJM
QbJUTOajY+rTGsCSJpmNj13e1oNpCtCwEA2TBzHdzEyAxDwQ0hUh3ZqnFSNQ0MMnavo9wEIKRylK
MAHL5TjDsmLJG1Zi4ZQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GFuz3jjDcNus13vZfabnTsKTQz9Q9tOYpUUTv0v99miJHiWg9X4Bm37tDSsBPgge2ZWYV/fIZNhM
o9RFowO2ZPIK8CdMOp5y1r9QlxbgxiEVYj1tH56LRgvbv2A1ghGFDDY3Qvyz5G2dmEuSZ/58uAtK
A8Mm1zy2Ln16qChURWHrjkDuCcIOuGQ1GysEn2sqg3E/XWxojTbAmy+LaQrAOqIwoDTGFZ/Ek5fe
49U6fyDbugt8sjMOq32EEkOAQwWmc5uVOZWv3KIDCD6tRxPMIg8J9cwcCTEoanlasaaRs9KqN5go
7g24OWiCSjQz8Pf4KXR9USnCWt9Xh2mPsrZAPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20576)
`protect data_block
g0PUNryVn62xHXvwuxX3GqwZFAWw0o8uR2+QmsKUKKh2LMC1ln3izCyNaRbavn+6DLpG7XGBI2kO
G0qtxRws93q0YHimuAv86zf0UxCdkDx8nbifR/6rPs42xWB2Wf8gfq9KyOKzA9zv3DfAyiZjUR6v
/KGsfQ9JPwj3cf9oJ2VvyVtmOVAuk6gCWbcF8d17J2T0swJLsdGS/iuMNCIcqcyEgGo7NjXkI1s/
wXpRLll7Mr1+LCWvNHo3avspqP0esjhkoz2oRcBp/SiW23xP2sk1YOqhyUwsRmPCjFELSg3qqKvo
FJvmhDtXZ2SalQNXnHd560YpQT0cSoenE2RCDZq0Sw2PuOfKoMUBr787urwr04MlUV8vRdTmVKn/
dORONChQCWg+wo/osL4Hn5mFcilmGyFwQCUZLDm1qi/z52Fi8l8yqik/dDRcFoVmLpDBuVBDU4ty
Hg65K7jerpH48NYFMIbg2amaciIRxCwrkfNT7rCBE/ydeLw0y7Bb0M15h5QhfH1diqLRTD1fbDWD
cHzLExvBQ092hQMC9GLiPhmQULmhzYYyD0Es+9MQNZqnubg1Trs0zypDp04yYTWLIAhfhXyN5G+h
lYzFrU1ekNSAnuc7OxHsHyH6pyHdbDjVPM2SqKqkrZJ5e0tFbMcu1L8JdvgUztqWOAEGlmChbOBS
dy1uqVguBnkZVarnVSbJ/Nbu6KTzI8gg+nxVHjB3vrZT5wdUWgfgjOc4bCda63583RUlunbqqO5I
xERCwU5D/3p+zV61hefmGV0KR92kz/Lli+KTIL26ReazvE0y4AylkIeu/chUoK8xWIceoiC4z9qt
bbHgEUxZFaTI1zHjmorqpfAkWRvulrc9RjMEFAI+4+2fQadryfvjKhyrWMPnQ0TgjYsoJox+qFR+
B5fut+4lPsarFgKBSHgRMBxiE0K5PsyjkjXnEq45DG/7Jd1krZstUVBKgxvQKAYensaJHAY1/ryi
Yt5+qt1OYG7lFimLh2TBDXuHD167Tgrpnx49pz/scuH5c8gRhf/QLFGQs0Aqds7bLkkUZL82RlIs
seKNGDUYp32gxbzCuJgkXn1cP+BlUR6uMMt3EqdHdzk0DBqPRRUo8oQ1m0WhIm1HMFKvMrYi95mi
IBsr7kDSUCo413uanbpbaYC5AgFUYwPpWlwrlJaTS/4oC0pfgFoAYLExaNZuYjkTlMClk6NgIGPk
uutKZV0QxS/8MTJX4vK7NKyGASt+qMhchc4zZjliFZOdG5+e/HVSTf8Orr+W4gXP+we2nYgFD34p
WvtOReiJHtnHyyf1nz9edlKDyFR2xWcRBMDNx57Ou4jq/6Ur9bLTvqpB25fBjbYqVBqwAhPfv20Q
S60Ivcupim1TrsYpERVkEYaAxCjiCEUZNnzvuBX3yHlFKQRt9ftdYHrWxcwvyA9SkPwG/FAIW+mA
VyG/EnHl0bpJsGFuBxj208F4VmkpO0ESM+Z2gfFS81Indivb3HcsvxNl+sO1NH1VE4HoN3kFXfWU
6Dt+dv7iwyzQbb3yzWYguNABBLkTywl2wBYuFp8/6cOSeUwdsbmpng5BhnkeFGDG/bi2jVk3GKJh
Y2NeqzGcrLtJVjulEtDkYFNeSQaHhAZQKhD1Rl6le9WeU1UDY0ZTghECj4WNoKnzoyZX1ZQnT0f5
vxt3KaPbf/kAemW1XHwYbH7M8QNGN8fhj7PdNiBcZANoMXS6raDfvyRygLvcLwYcKS5tSruyLqkV
EtSDLktBvsx/1ALFiCwXvsgWoPF3ym4enHJLPV/y1mVPvbpPhXoMsOQ0+zpw0L16upvbzRMIFc/M
UEHqOMx69JcLSQ1Y6gZyBzxXP7dGEP3jtdff/Tv+eY04sPqTKwf/rMsxtWzPMqbgNREfwZJaHPXi
+N2Um/nxkU4hfKq7uZ4BkQv6GDTlFTjFKuDCfXCquSvBJzeAJEogPhWeQhSWcbY3HLD02o7VLNGl
fw5pMMJS90Hft3pvKYhEFs7JXrIKRgPMvVHdXmtI/U0mKHCEWdTyXVGIMCqUK9fzssn4DGBL+tda
gLxY4/80TpgI9Bex0bK70fiT0Nb8PTt1NDyzqchFg9inSutjJKN/H3v6HwQBoKn8PNlolgydRxxR
4+qwvzCPo/ChO6taaVi27xVOhvBLJVv0QqfFinf5dFw8ryKudl3bxgfKvsEuJWvNnjXBtczDHKxE
m8no/Py1i7ToSHT72LneiX0tq2dUcGuSfkIW9apDAwyOJVwBQm4ZFwRkJx96SxVY8aBRL17PS9mj
2wVaxouv/5oyAQOhtfPkRPTtaTUbcXXD4cf75aDginn4fxe+KBQ26SrWACaVfrYjfk5xWvlAtij5
VqhmTZyPqVmsIBroh30REPMxek5H4of+cytloKD3RHrUoeZ5KSZPHed1zY8QjA3/Ha6j/zq0NrW1
YJFSn7Y9o6blzvTN6NMAmb8dVVeZPNqjtsoFT2UxQmclYnACC4t5Ut0W8b6Ttp5kRR5aDThKwaIv
mS3K8deLsjk4lFfFNc/IRTDFNTtCrIHGQfbJm1OFPlOdJsSjA/eiWmdtFgv/rs+hm8ftF15EPtBp
lpXr0W6QvFUV64ZncJnpBwFgcf3jNpVrk1L9Qceek5siElzGbUybAgof6cspH7PAGQDmvO4SLe/M
jIGyzleh5dmrlG9AgkUxKt3A1+9bxUDXYVeVNs1WYDvSYNwzyTVnWNXLTVbttJd51QxJ3Dioo87+
0cWWdCw59ac5NRH9NmfA708MvE7h7M2MD8X3q4LF4WBPZasOUYJNggMuu+hoGVLYb3dQM392RJXx
fEFNhAhQJdjIczt7xOoTQofBN0f2OUG6EaK0FAgr6eJYkm+RLOKdqqk3fy2pz9WvX/AGlbN6ZrdR
mVYqubcBKoDCSvEIkKjKk2ykRZoiDAjpT3S51vxLtm1orFdp+wJsYRRjCef2rYLHBJAca/6Ki0E6
XtvTdJKlqACfxLhgGwCzFlQOpsAWbM4A8Z8YpdHgK5tumYdXjONDx8o2IeSSWRvSixFqg5PyR2hn
797+CFD6m03QJYIvU/lRuhs0K5tYG0fKzzMGewdik+cJHh1qWOWaUna2WI1yvF11lZY731sQ4Xj6
Gw7k1YrWHo8+afX7rcFxzLWP5vQo346Qhqapuey5kAENsgZxSvSTiWxH6+Eq/jMafyy4XwaCr0g/
reZphKI/ROtul/AQMpIIsqM6vmta5byT3zX+CVoeLXdIuHz4uGvo8EbdGit03W63PBIelyBhW5mJ
2Z9TwdIeb9GgWNgIO2F6VI/ZXL4hI29PWPzN65XPW9HiqHFWOgQJCdwJKBL0elHl8b7+a5w1qg6w
2B/47Fa/yLJH1dtqWMCfdG73ozMkEIBkOAD3SFToBPG/CJkojMtQhWZdgx0MEZ+EcdrIMo6xgo8p
8Cci7J/RSLpETp7yam0oIlGcHRU/w2O0OuyQkF+L/tctlQ236SBRU/J4vEkAYPrwm8rkHbwtlSDX
Bcv4trR/yC5idzQdYC53bp0VpoxVBriKk4LjzPQGaI1mWrkO3viFWmIjpLf2+xRJtSUwJNDvLTBa
0ODDNMFDoETd3Q4sGVjlrlFFJeKnTn7n3kk0cE97EKRsWPXHEtNpXImwR8hPzPx6O6UJqosB80Ix
/1A51JSh5nJZkoa9/nSu8iK6qexcqSoZxGgmTb4sjAeoZjnWky1CTjt0WBHIOCJKuncNKricZgiX
o5EmaaWTswsMsYChz0Y6awweeaw2kkVLJj70aVGEGTlLkzjYpeiRna53CIUWfVEl/Y3w6eAGY0oO
QUlsTM96B/+hDGo6j+CpFS847i0YAd3F7h+bJdK7/w5KzDSbQLqPzDpcJblToLWfu45N3lzE6JBb
b3qxGRN6L+GHF5Xc69V3RI/TlLz6fEBUBUiyuHhImhtrcCdgfnmO1jH10cXnW2ELtJmCBiLrCnrb
+uw17z926dnWOjE/qmAkEcEFculVMVffKdKuCkJOPGhPJ2bYffLsOALgmlFeSZYdWtF3H1+mtA0J
anfmS5KC7udMEWIQfsoT3gVD4fKzpBe88IgAERvOmceVoIJCXGGtmA5j4IhrIkTfqYV63i6hnmmk
bE2vPKn0kAJ8cBGFoA3ZyS5lqt8as2ubx6RzqqxpYFwbF0WX0y3ht5yMy44KCIKkQuP8+5E77mm8
177aqCkUtMQBwASPVNa2e3TgzzZ54fk5SGQ5h/tMdV/jlwQvyfceHCgq7cynEnsh5kusrHoL43ry
IejEZOWH2xF2aJulmycMz6ldgg4LyO1nvBxXIGA5dZwpS45ui6OJV6v92Kf6I18yuW81IuN7SudV
N3NMyPV4gmz1ntcw2qauQXhqUGWw2FEpFxlbeRxabHBP5UeTzPfis/dVyrcp/2o44UuN/Ivfyayc
m0QlVa/9HDGvVCFeYUJHEKD/mW6Uq3CRUwqjp/+mR65dgsoLYfaHfITxlDR7/JSaoWbPVAFxx7mu
dYWY+FvlUHHvOjGXPuP62RO38Rt7av4dqybPD/wkNDDKioicsh26OlBhZdmGOoUnf5t1dSehAHpf
vwPN6qUq6TXy1ShVmabMqRNxW2FKVsClawI3Z8d8wWJn/xjLgiVg6vjSgkeCJC+5VCrAGUyQTZ+N
0sOmgzXDzpMgRee5Njay8f8p2ilMxvy2HOqWlMM2+/iJc2n0qOCaYvC0SZxT7YvWN5y7bPuS0j8V
1rlpvHDDHlTgpc5r8a3iB42CkIvU6Wn2X928UVnLKVpNYctve2ncuhBodASKSVomQ7bcWB5ODZY6
4BfrM8u+EY+nk+iSpzuuu7gAOD5MsC+HXkJfoNwszk+Z6nzf0OInlReI/rpqyl9syfo+oUxJNMEX
l/yvlRy5BTwxo1fxO5rKPaTm6m9rZlloXVWtNGmVxDcqjHrjLeWiac5Uz5f4v2J2t0zeaW5NeKRK
Wpk6MRkBs/8ZtzWfrpqDoQWr/0UF26OP++y9IonKBu4czku/33lfq0AYxfiLJqY/QjJdWr6E5EAG
0qz1J/eBZmBQ46PwejDBYcSRvMGrRUwztDMod7njfY1yH8eHLxk/3HskB4l4LjxCuvR5u0DVdKXw
h1iVLGUHoVqxqQwWns8SV5bwSSnieykCbYeR5ibsdeMhoySNWgFQF1fqzOsRBPMWYRM5v1Bi65e7
m01erqAoQG/dnC5T9ncG+VPNZg7pGdPEtbN5qBXTWa+lrKeb+VwW+xJNe5gGk+tIdDppM9XGOm7D
o4QgoJZ9hS7O4tBmjkjyp3QP+drzf+Gu/PyQGlIFXShHKrGZvmsOcOUm1p5pfEBfYETFo2bT4LQe
XI4IyYiQRARWPACydjeRS4Cu18YH3vY4yhuD0Ioht/UhvrD5h7r8IFa4FCCqicriQcVHdqJ7L3eJ
fpfbDCcSycLXrYfowT46eRvtJMPWDcUJNcB3FTWC7bAaP4vUHegurprSsNVXBx7CG/P5wu1H54SA
E9dMChJwt3TBMYFSgc4yKZ/ORVSP+d2c0qmjAJN0DvkTPFUVJQidt7aNNaTzxcU1z0H5WzkSEqbO
orfaryxj1DKh4J+i12lFfED6O9B75wnBjCW0yayMY9L/x2VZY14Pa00O3oe3idGasbt2sQtEBc0x
tjX7hbQzxgWqNvxDTlu0qnfPZR+uUUginkqVX2II6wi0CzMZiDc930iz3GJMMDH8z5xvgSdnEssP
fINf4o6liCvRe8mjuVZhuRbFyPIbmmn6yWNTsqcQFPpNUjhR/61Rn7EwrdOeurpsDLecWs9Bf+RM
NAqCw3we6eFmkyP2IiGG5NhexMOlwpwxFnIN45y6+Wx3RXBGCJrP4LOmuE1itbA9jYVRTU8XiVF4
I7CCtkWo3tHKP976naHDVb7nildff8E8W0vo+Q+Pctlt5B0rLn8aHi5c2A686lte0mqyLjwHtmYn
Pj9EK1amVrkptSAnEMsQk7exFqxGwT8p6EFXuft25feGhrrcEh8tGzlonLZerOqHqRT1y4x1l4k2
W2LteYGAcfm+/2+ATHYQ4MlurvuKyzcIRCWYRpolqeGiVG28Wiq2FiH8P1N6NNRc2dzcizXzbTdC
UgGx7vHv9j7y8M/0dSoxCc6Q+FhDtlR1eoHaEAOpUIu+zwrmNQtWSuR50alAxvtiy3w8oshb145b
YeoTw+yXdFijfEHQHqg46XIhRwSX1F5KRALIUYH6GTm/C9d4+IcppXx4o+y9/XfOZB67RkmLr0rg
lQhUZnuyVmYYCumPVy+ZeURpvHhU5V5tFx9xMQeq5RGRIL/k1y8Sr2iv0mcstC1KhAEtNgnXgAyJ
hZrWl0lXblEntimirxNGHEGkSOUpaUJlFRPEegUMPmXGRxba3y5IBCe+MS986MKl5En2K5P/D8NX
Hi1IxLZ2cNzCtL8qzBtMmcG56rcIkaszoQdjqEvMOqRkfCo5bWem3j/1/zjCHzcXc4k/qVNgEFo7
v3Nbhz6m/M4FBbGvpUKt7hnYYwtRy8mBpBSYPMGpmVoOLN4Ip/NDdsczOSS3N0USktjnuAVhr0ho
Fw17IFfmSgltjRLTovJngdnHMN0fFscMbGX3urOIkSuXkktkAwxAF24CdLjD6DO6FWymn3K4BQzU
AU4HonpbvfiQ1RqBc0vfqpbSrt3kulqP2WQ5SSRIFWEE7Jgv22tBt7DDzwW4+oDJo9O5vV6wqa4k
k6V5pHBPS3TvEMBVb+ObcdC4+118L+MA2dMk0+lqNEpmNg5eIZu7+xglKvA9tgwtZDr/JbOBBsQy
rmfTQdfnS+YTmvFxTjJ5WOPtdyaQHg17TPnhGsw/GIfK0fHjopxTyfgo2JCX0KPGrpb+NDZcV6MD
8TP5tYCswjDI8KOSUgMDMykRAY0gwGnOo7AdmlR4ukNkCN8EJGtNrjVhGtX91l0JVp+cm5c+Vz/Z
5BWIYfYIAVe+V23xpMiSqFwLZbgp1Gky1KRfzOssiZRhHJQfeGGiMyjQRW/dwpcXH7kEjY1kmptX
Q6BdhZQcedHoXJE4F0xQbpfzmtGG6524AhlRAWNG2G0oRINuz/p3B9ZoGOKxSf2pBU0/r6XGVo8n
v8tvm7zbfzcQweiEJwXQB1cbvS8qIGU5B/D5lcJnHh10IrPa1/mIUJdluSGGhD0Xw/LHQXBMR8UG
Nxx0NRu4vUfhLEYxXTbDBEV08HTVYKuRukhvf0Zci1nU9ZLtBHy0RkaGy8vdgDMStW6fyt4i7S5V
gb5J9JkF+J5Lxy/rNuMWIt2lMRwmq+2q/tMbhDGHvQWk8t1YvspMSIpQcfvr/PqOGVgGlOUHpm3/
5XcTTglI74YsztG837b3U2wx+lNNinT88iDB94SGcYoS+H/kZ45UpkO9w1TdHBkNiggRCOY3SpiG
LolAzxE3BDe4fj5r8GqrWs6ZIru8sRYtKBHZfjiQlu5brvguk6+qu/5QEq42Zra3SfCeNNdmeuk9
7TeFeSX69SRHgcLfQMJhAyLcSzWseWzSwEytIgmAc5ElfQAGvxLCuhdlhEAxq7mLoGvX8tv6t96V
BHpOnNfnMminm6D++mDVeiWSrWJ+IBU/ho9eKFbNGdF1fnzE7XphT8wthWuPBQVCtv7wbxZZykpq
d2UFA1unqoNDIlqzLKqIbzpFqMXnSnr8WNXiY/vs02kgBzsdd0OvcnEWQEIOcKvA+3Yp0K5hmolv
xjO/ZuYhhStjfltDVKWsyD8JmB5zXfKNLOkhw0vZ5aaTHBNFlu2bYIWkhFbweIX1xa25PbIhgZdU
2diaINWDanDvzc+sayCjk00O7FS2rGRZ3SKjOu55dXYaPHw8gt9ea2GtCzHoPFb9+v9//Qu6BZLL
7sjPVMFwaYEn/8yu1826MvAOxnC97jY3h8e2BC0ieSVOQcTXPexId6vfn7wfJ59jF1bNcyiACeP4
zFJBqOKRGki0Dm/IYmiUPoOTFf3lkGKswHNsunSx4n68qKV5waM+SMu56XpDlQVJ2LBdgvIueiuP
U7NFk0tvup3KLdgJOUjJwMA/hpIKQhM3Jj1jiGU+J2S5eh2Tt8+ZFaVEDQvnFTdF2gVUyyioD13n
yY3rcMoHztKz0PM4DZM3fgBkrfo41eLPU56eTdf3Opir+vpDg0TbbIf5XeKeK+fAU4aI5FKJrasv
15MCErOno+8IrO4fHPmF5/uPzkG5FomuJ7zlJ9ljNNeANJzQAcSJD3kvvPfgCmdb/lstik6Z5QB7
S8yaCVvQwEKK8eA85dAKMZImMGKEw3ah1t+hd6QNWBtbV0SXPAduJaEFeXmW0t1rSGO/Rz2DbeYw
+IxdsOTNBcpwTdpNpZtEerfjqYgHeho/AY3ejOimP6e+VQo+BkeKSvZzCVdeFw1wpkt5+m0dxoS8
HQTc20It7MwerGU6xlrmIUPvijYtzGXROuFDPGpb6E4aQKY7sNDUmzYFUN03/ZzFLDyFyshqjc7G
KC3UsHTo9inxgKY2kLBsx9w2JgVQtMYVNlqXSEl7iPhMLIkBAkHIakG+2nrEVJM4EqvzGW2nmdqj
pgs0bUPZIsSmPoh38ZP8qJmbO5uMrKWuVEWD2pLcCMUophhdf/GBL/44ucMI6GFYO1tkR0favJou
iszYG6saTNc/x31KrPO0lN4H5CC+oeYzWeQ2iuBdkvW3fj/TTgaleDUvD+jilHoau56LFM+n8sjN
z1kZV1o6mo2wO//8oWApOJnYLu2tXQYrdT82BvUr7CWhCKFD91OgXMgrU4cnksuIZ0hWA9DcMoFx
yHk+T0UA7tchId/DXuN7KESqWW+FK423sOXR0oXgzeVrNM2B1xcUbt18xWMWZruu6K2NdUipqhZg
mn5iXOoNMSFfQ+HDgJGSeWWxx62xewJ9HcdJUmknmkC7QRoGderL88V8a11S02tgG/LaQQYaLcGw
suhF0vCxbKDpGYspq8G5hcnLCPqXQvQ7U0xSPQDfC2/aVXr80QhIKgFgTT/zlcQuJTzqJO0dWSxC
xr9jQ2DR+dwL2loJ2zQUtwOHZeBX2onwbr1cSlqPSer36xeFVtFIKsK2j0jdqdtNZin2kDBnh8TM
1IAtJeYU0jpJFoC3SGwmhA9hMn6fWii2vLt71WkctLIjOFygJGFGwjRLm+LV8IEwsjUj42pHm2Q6
SvxhUAtL4rzshrIToC6wiXDgvySQ9SJlsgLwCkZ7bsRDWznMZZ6AjY+dR9ArYOJTuNRlTasKf78E
qW5A6wIQTR26Nl/sGXv4jakT5P+2BXmcCjftQyFuckMmQdM1Xe528WmgIlVuNzT7/vDwZds654Ts
EoLHKYtPWqc62hGaaGKfFdRFpT+Rf2h3Q+UF8VddGtH/8LvXERBOKJ140tv+ypDiLBwUYMsQ/Gag
LZ6UNFA3t5DHfN6d2vqwypDGtfYliW612POtRyqgo3xkDjxsxq9dbZxkgGgx5WBp3gNQmOn1iVXu
1c04EilGGf15P4jYu7x/ynQWmbMM07LXRBbMyahqNuWvrksvZ9krQI3NmtMydGVvFGZnoiElCGRK
hY72A9H/caopgIYvAX9rfnXJKedo3ybFUXb/BabLxJWpLSMvO8swxqsQIAr+r0UlZeHR+XkMaUjW
ZDCxsvEcsBXHs0GbM/FxXn+ISy3rMEjYUO27rtHOn/iOHb69ts0GRnxazUqgGivgBvxY2k4dybmv
s01K0efaoh9fSk3ECYVG0hy05CGdyAXwr6FwK8d/772pNfx0d40eHdostkQa04exe/BnjP9vDxQE
VZuImwQqBNLcD6sXiH0Xg5x112mwkv9xma7RlNMAdnIJ2HpkgEcXPXJYai9W4K+ksuI/Cx5gSJjh
vswogz1QJ15drfXaQBeps6lGg8JqSpcpUdekEKhb7r3F9j/V2fjJk4hzVwrXzHEZviUcoycdnASE
6XLaDrxgZnmQVLla4W4ZZx0JBNzgq/zuGpmpOjV/2t3hAaDAAaBXp9hTqRc7zK4iXJS75itWeFoX
Yxs6ovn5MVdrqOZ4j5H+cFQk7458mBObrFMOFj76ep8/PGQEzHSPrB9skvBSZqipNkuuLAxaUNYf
tW/yytV7nz/F5rLw2SZpTOuzQOcI0iRNJXsP48dkUzClKjh/+81KN3jpVGMFM+Giw8u4llzGq2qA
MsqqMm9tJZab4tUQyaY7grg8JBVAUU8f0uyqCIV6TnEo+/zveRyH4ELp7kr7ic/r/bcMmyGbAJnV
5Te3U9G67qGio8jFOjHD4jtvM93d8jqiR4GnZvQjO0J6tA2u6aI9GAQdiC1NcflO6vDOroQqKE9/
lVbwbt9AqgHojElhRKtD6q04jQ+TOTdY9I3SY2Wr+zTsGER2SWO/a6lcrLCltukDOhilfIUcataH
l07o7WlBJ5OKKSP7dBFscfuQIPE2K/K0X05OTNttPiXB6Ezo7O2D5VST5fDRj3oaiFzXsN/E+JbS
ehAXUqIZdk9XQl6bOx4gh9OWMwDk4o8OoXHAdEMpIloB6DOL14/EMnUqFQ+AMTtPDv0Zx7h34fpp
lxmSugwKmN19tuExJ4nly0LHy1p+DyIHEH/zkhhHI7XXD/oDAVib+3nOwbgDT30KUCP8MAeLXPJ1
EZcklEWg3EJXsTPgXXuz6HijPN7RErmILu9dRXyO5AI7StGqYV2sIBLvT8esyB+zJHtlmtSz220v
IGDO2uIcBjJBDIbnwgY/EdFBDGSP0knACpIowzMsswibBlKqBfpUOcmIzAVuFEZpNmi8rHstKuxg
G8Ojtb5ocK0HaOWSl/lchnabwzl3N99BSS19c/paA+EzqELmP5SVTJ9/H9H+EiHl2hpCXf0ykQx2
JzILYuTL53qTvNgrVWPhU+8Cvr2/cuk+mj0qZfjisN1EbzQO/qhOHQLsP54esVqpFLfagf4Te/t5
xskHKtCmwc0q9TFFrsWzkqHdrwPbxmB/lN23zUOmZO6eKabAL4LCmckvwSugC4mMSX3PQOTsuH85
YsxpTW8787N6RR2AMSxvXTY9VY96Wbb6gxlm+bxfftv5x3uZUe2dt1zshkKFzU5oVfxCYfz1G15C
HnVY5VIzlGtm+lKNla2aaWFbxYY00d0tagMEULuni1rzI3jDjrvn+CnuH+2YxxOuCVAKYUNMx59F
MR9vyDbplE8KfXRhcTRijW3pJ0HU1TihfdfUZfn86UFdzoBX6PjfxZtcLFlpFtD3vjKzTo2TkNd/
0uMNK50me3JcQRpjtWw/DpfsgJ4avzBSdWzVb+nroqRpgaSPpoiwJfpwUq9sMAZ8LoQLPPL6wfA7
Fcdhe2+hciVSY6tYZTdCbqdSp6yzoW4knXZttb5+oLjywM+jrbEQ3fDNktubV7PRt5Z/mOqNdJM+
Re6tpXvhNjDUpmKuIooQwLj+PdLYPLzqXrnEk3KyJ3vVaBeVuwIWLTxgw7o4mB8t8DyUhQpoWazp
UFwzY8y+pq1+ErBL42udEvm9MHT9AhcrJxR9yVS6Hcg65VIm0T9QRzuEtLOr2D36Xrx6qibKVGeK
aAz/OrWSby8RxQ6MLWr+SCGNcodgi2cpRzWzGc67sJnW1vdVfPxZYTGZoXfFIL9T0Kz+e4RsPlLG
rqRtmeQEZ6P3PONoLFUjPKYHsxzwfppOEA4wpHANo+5ZE3e3jBj/FMvRHovwH7XKXFkTIW6vPLCC
E8dVCOWf0qyThlISfaxtCcbILRJK3kLipF13Q4p/MRrBXEVbnBnwYLsdUVUOcfXWwedv/vpOp71Y
osY2CFXrGpnSTofAbZC3l3ERG3oeqiXO20nDxvwMb/AuxeoL+93J6b2meenrtlKyL1WgTdWHZQFX
OEkneIcwc49Ik5/nZXjcKI3tnoxNW9vEcYBlQpUCOQrR7cw3Blwdz11V+3CyYcGP5XYFvaTLIv5A
+nKlizpLbNaF0U/Ah41a7yIP/YU7XBIG/YBICeVDm4NJZwkkQrWHem4J99VCaEb8wLtQ+663LNlk
A27k2edbNQW5iaQwNN/wuqkAJEl+bLJxhUKWa8lqser4UmceDrpSbNsnyTf/zokNhvajjLEawaiN
+wjLi6QFeaBSR6hWGKZDwvHBVzSV7uhzpQ4iM5MmsjtqOtF4NDH7r+2imutY5jmZokp0HXev9qUG
XOnZQRFGzjHXU8bmCpG238ngGnydVGy/IESjAEHvBnM1Mrz4QR2g4OuoZKGek1fbBqXV/PewN3ox
YzlUDVMTYMZBnichPBTyfIySZQ/uC8qN1NmBWjyEYeYjvNEbvfr5csj0+U2qZVMXKbnf+FNXRnx6
xG8pjsL9w1wY8KVsZtdXWLxU+gqg4jroLdp8Hyzquf5FH7xzFzMkEoENkPkBW+VO+zRjRkY9l8wv
5V/+JzPTGd6I8JPEALBizi5jwhC0jN2X0hK56TZO/Tv24DpHh6/5CgG3KFx8slzwSG1pwyAvEGcn
9wAZ57WpCcfnr1uPB+j5PmOoxQfxtty4pMIJPWANHyqgmbDkcqPx9XOIk3uyYMy6rbD37vGzKVQS
j3sfV7H9o2nsuu2D2TbdUNll5oNQHxcOwZP2nWwZVjh7Ru7/jnnhHYu7/DMCkzJUoCU82S3/iSPx
CVkhM1nl+VtRP0NVO6wlnpph3PuP9BsBVhvOjkk8QAuDOpLmKkw/Zdu6jA4QABVrOB3n5MlSsOJB
E2Y5luN0BdeXwDwAuCKRfLVgJAsjIr39QzZFvgs+4MHUkE/XKtMZp6kEH5mxBgub7g84HDoG6rMS
5y9I3RDsOHg4pbJRii9Ojxa5khwn1yWS+lZPQzR3tKpk740+UsyNl+35Vh8QLN8v6DMZDcrdxQ4n
TqSiYCKlyGEFRALaslEK/tzZN8HBO87j79ru98Zv5SJWo7fcO/weDfrsgJlDntH34wvIKPpJREEr
FfFYGn5FCX557JyR6jlD68stCLl/RnbbuGDGdgXe520oF873bHmoWDd9bnUdpnKR1xKl7jBzn/8P
UUu64SNXRGDuYAPFl7xIP19ObxurKWNStpI3Ue44Uy79wPiubc3/Ac/ij8qd/LK1NOQZVqHHl97g
nCOeKrpxNXQzDHjotHTRM9Wj4/fTpVDLbeBn/ZnFfrZz92O76CPS1P0BXL6l7Dw21CiFYd03Bby1
/HWXadRbk2iHkQoMfPQwlZV4hLOTBoN+cJnNLMbPDqpdAB+x9aWfX54kCG9zyul3wzR1O13neKJD
jDceaoc0UDAsJ71FfA48D4fJhBs3WqCaR6pYv2G01UUSvz+68e0JDi3Ab2yt3jPxI4fcpxNK1oDt
FHa2SZ94XGTHbp0UQNDloRJbcKljRZkfojIEzCI6ajF7axZuhea3DcFdrA79FQnu3at63uC5EXek
zR0AuOeLesgh4VkewKKitTnS7HN3KOHCizPoIM5a48JSIgTqMuzBrKgwsi2CbBOMoMWre1Gevxyx
Z95XWy35efE3OyTS8V2l29GnVsoiBbl/p3ZJ6aw0u/4sdzNuZJhxvSBN/uNw1Zxe08YMETT8o+zb
+/Sj0J/PMGfJS7lH7FLcQbMfYGjaNgYvE4wcaOjWja0OLEz9C+nmuiV+jQL98DB2NE27uuUnppVW
z4MtpXVjCvORvaFfO0o3FXCaueVdY5b+1E7DeS0C6BbUaI982nvyIskZZfxxSFcUug8Rc++DVaaE
w83vGVrtW27SkOGWrplxCKPKSlpPaMuKyS2XIhwPfUIn3PttdqQASbZeh055mIXTXOLQaPGRDh1u
nwLGrO09MRuPBa88FHS7kanWxmpWg4nfF+PUaxjrmcYKwswmT4pp85AMQPzD/WsgOFt69uGUg4qn
Y4tSr6ZZieNhHGhGglK/7Xs+boxAM+DcphI2TiU1G0SWttp1nBgUWUofh71YmtREoDPxJFfEan40
xa75/1nqDF/+QkIfNZj5oJ7p+B5605mFeYCQdIzUwikC8snmrD5p+gP5xnuhLyPwBepykMLS72zl
FBQocxc3V39CyI9KfBk9QoeFF2Mts9DBzWdK5/VzKTu7s/ylT11AY6bdyVInn+WJlUOHcWbzR6ia
CxKkIi9ihz6CaXzu9G/tuxwL1hdB6M7xxwyzFafvCPYvJu/iIcPbK/9GqBLMByefk4U9ESagWst0
7w+qSEPxDfqzQiVQr8U91OJcAN0361VlpmqfJ5CfH/OxpdzNCvPkZiFGnPIhGZUuLd97HRwLuljj
dVNrL2gA8+zT6tHSz1wrWtXaCZ4QRP3cdpjtDK9f4p9m9gkbV847F3PZUclMYRwOqxwe2ZgNjuax
NvXoBt9b1TtvVAsHz2vT5d7qpEkgQ/wfScnate7ZTCWW1oZVEo6dH0P0IhstdV8grbWOvBpaZ7fl
OKkV6MioU7GMI4te0WCngGwJQr/Ibd55IQCpinDVajMt1dAmXP1F0rStDREut5ZFHVmQkK9rQRwE
v2c0dylC/Du7NivTtLShGJXp7Mw0la3YCNhqJ6dsurDmVZphLi/gkiZ7PbRzjZznDy7vM4AuZjZk
3ba/MJ0qwBC3JP1cRedTAlahnm1DKivSJdYj71BnLjhD4vZIMtXc111aG/wOYXEUb1U/UpXJFmcv
lGwxaCF1jrPeg87728jDTVQsdzuyI4A3icZEa9p3HMIy1Fubyq9qf5h9/4/sriXac0eeh4yEDSy2
4xV+MvtFYvrUqIqpB7uVy/SU6jVO9YUNcYPaDEqBvCFmqwNb24zkXI+r8uFLlwsdzzI+gm09hefd
skHi+VHFtXnUrRUacSRH9PMejk2bdLF2d/IUPaRbneWYP7Q0XxJQRrrOyBEsQJvEoZZGpjkczCTv
YEIocz8QrUwrbVBCYrGvp25qQuDDRa/76PJzJmfELVN5DeL0Vn/sK1Ntg11CONfmfNhKA0Zk9diC
NXJSLSZRw3OttKKRBlmQ6vadGAL8dtjWnTiyIjj3veRev4Dyum8iVKMfBNQ88ieQn9Q6vArnMDf3
28WIzTsOkbkiaQRYZadWmN19ND80nk+d5i55VvuVUaulLvjwyeKU9Oh/jaAvBggIjgHvUU0Eo6KM
KXIOtswrshYWFxOUVkhmdDrbIWxCofi5r7ZQD04ZTabgu8Aeia2Nlb8jMqVI3rfihcFXeGpp+bYS
d0tWo6hBT6q3hRFGIHuWf6hQT9y68CJSWsZx6F47GGw7ScF5PIsSNnIy4ZCN11WzBMvWMjtyqkm+
GmwhAsUGjsBYCwVpIb4z8ZRv82UBdDyCczVwiCl/W4PGl3rjvU3ZnmV6e8eOtucXFZlcVhw39ICv
9HjlZTTp6gnRPn7i0pCGSWpjVH4LNNFBrblyhEdsHAbwqGxULLfvv/nNh94efwe/Cn5o0yAdti1b
EkcrPheyYk+cDKcxpc1AWvMKXOiC1SFEqDKB1D2/i+DuzJ+BgdfxxH3R7Aq8wWtBOIDzfB/PJAc1
1T1cIRDr+zCEkX1JR8dxbROxv7tyjTT6id2bNEHW2oQk7Tsbl8epU3gtTKFIKowuLH5QIiQpjTQS
nevOlARS/1RbWAl8e3Fpr5ZmuLS2LklMZ6+WVhqsEpKOJdZkOBoOSLshMiv0Dj9EQ7I+DXDnofb+
nVzDer748H9THhXGJOKrnVCyxEOze+sC7uqtQ+xr5q/ze9+UiRFJG40vF3o2kt1ShyqHERL9nPXQ
zrpi/vJB56LVq6cEQOGVF88uUG/IXw7YQE712FwxL5cZONrFGehuIZGip99kiiqeakkYoHoDpFSt
Q9RfoWjH6QuWTZhMLYwEimb3lHQS247eXuZCSk2Ee2+r1QawdGYoRgLFmVe/hbWWtTacJiCf4ODn
RhlTIOg/qxm3Z/8CDvqKOD7lYsZQ61Bd8PvwdfenVBXBmrUdenVxIN7OUwT4mb/E/eQwT9+xyozX
6pySjlK1XbZ7GVuUGyrF901zTiG9cofQDjxetyTRWxSSdIF2fo2BPwyKDJOn5AgMPLitMiFbWUgN
w34/23PYyK6/2fatPWBKgig0rvFqx/sZmXOfRzfESWacMt0W/bUnHXd4mx4mOBcJH0jbYtfmd2MQ
u4vobJ7qqyHAeq0hoop9FOYK/C3XNcTDiEuhg9aIYsBCNgZWjTjUtV9SrHwPKoLygrwKpkKrLzE0
jbqiEJhfz8jMk7YOye6J2p2SH9s7rBfM3F2IZJ4H+TgQt3bitCZfAUxuOFzFK99srANXuRpkX8PU
aS/sgdfCZxjAeW9ZrvqlAHR3HPkNX4A9Gs/8J6NBcRHdPRjLSBaSk+DswSnPVPh1T2TT4rqyEkmg
78zaOh8UW24burUnB1SVo2n7HSS1LbY3Lf/baYOj25PffK5dnkw0YWnHOgbJ/OGHN3juP+53MFMK
gzQSyQfk+MEiW6aRnnZnJEyEkyyv63nYa3rGh0EdVNV+GzkylihCQ1JC+zXjDqJA39bdzpAaC4o5
t/EcHFaz1ETlj988vU5DJP7z+wKNhglohkI1cWafcNMbRUeFma8BVOxKL4pKbbpn0ybMPAJMlOnr
PSacIyep7EznEcAXPUkVvoKVKDERbVKCBA70Hbc9d8YDDhehOcOz8N5Ch8Q1y2aVQUHZ9gy3Igdx
IP0mBe9BsM3u4jF+0oBH2dSqUF8/G0n9SmfxkWht5ODqog1SJCLx1osjhGwV8Tu0D/20rRU40TVF
81x5oqzDgW4QtINisyN3Lgc/KaOPRdf4IWbpQgpXroaRFEfL43YmZEny9eHkZZ5rXHTE6wfJP2WA
Hqjy8RgSoIjbbawHRHlsQZwfi0cQXRQGBGFTxkai5c60+D/6V9VaxojDm30DfJNfaJXC4ub7rCHI
UtZdD063xc+6J5EO5o779ZwvTJzw3/2FeQK+dUEK/0la/EGwk9Rzpkwh4b1uzpemZPKddFGOQf4D
FRBDFbq/ii6IFCuR/4yr3hIqfZc4iFyPeqVLvtC+QYUde8EshwfC3UdjnaHs+wp1jsV05MfHZjmQ
ALxpfMGGvE6HMLdYWO4E+bKWe8tQADS42Kl/3ab3CcroQ+9AnKBWL/1iArlmPtur6eemFJ4xb68g
pUL1VYxar62RyGx/wJ3N3U+en3BQgMdDBHvFXrsp1kSsRkEyrv3Z+Yw+M6yFMx2sZ9qgXbskszsh
JXhHtP/5TLrRCAoN2TJ1dxzyIzLiU3P3TiCpPngZuNkabZVtnXsCRBx7UXCzmu1YhLyWlWuAoXrK
BmdmbHwirOZ8oSEM5Pd04djMQUNz01/OVCiZFdu8RJuNuHsqmySTeesLMwF+DJ2GW69I2DKQ4gHe
WdQ045EWwjnHr7Li/ae6A8ek3xQ0UiK5X4J0Fx8/mb1hAPoXX7+J28bIYCBarlifxF0U6DP0Sq5D
uN3LXDKexu1NuoTyuV/9HYrfJ1WxVZm1MwPiohrcljNDg+z4qpPTWc8becNGbqunhz9DEoPxRwuS
0JeuHmNNCnupZa8cz0lqmZ37Vcan37NB1Vqnm96BP0Dbr0U0nkA+5P84E7VND5OraIyA9/iT6MHJ
uODkaw3efXQUcgsB4jn2xePL4Kx9340vYIl4r+isCgLhoUc0fVyM6E7VCht2WG0x1R1vBe40q8nX
tJfhFLeVmhaM59xHY47NcmdRpnPmjMniMi9VyCGyq7VRhCw13THOlKbQMOU5OgT3C6ue0fInZ8Qb
WtIMD+Xi++Hq/n3cDQqdsUgmKWH4/Y+R54zs7O0tPBpyLiSxEfDlVsxHS+z/SdeKtnH7IoKHF/6J
RTjZq1ugw68GODUS06SLg5aOFZ8FN6ZeVsqwwRipR/wH1EHi9lFjU9Ht1jzLdvBH8avZWPQtBt3E
qtZUOrQKvpp35bY/TGTp0PzQ5it2MtLwmILP7Igk/MMhwJpKDxJD5W3frb32AnZ1KNdEx2h0R4O4
gNY7K0/Hd3WromzhWX4lfU4jguLAvP9KLXOWS5d8kvgju2ORVXQyChE4cAMHTjXsu24iyjY1fim5
VfMpDLTE2cTKY5R9mCBKzFiEFY6E6InekJ8ir+Vj94xU7cnlJxe+Y1c+x88cSrW+YsN4fyFP1MHW
8dYGiw7t+FMZVEp7UhSSjJTYNFPVLGY568J5AGJk5hE8st8d6jsCUvcHWHMVDD96AkddBweZ48y0
lcsOaxB6JyvMuc+u4wyi0nRnzHZy61gXm8rdwxI4xzP1JcFwpZinE+ipKcr0NEyAhL5pnd01qL9r
CHvAuC5DuKbiN6DNfLTnjvnJ0zPnDClwLIKa4CzirhqktTHL5ARwoVkd/HO4ChZNvFclgJmFv2hq
KMpW4Kz8+llbMTg2wTv9SQ4/RMKsm1CzQDTXMWU4GYuZTrPBlDOQc5jM01w4/gEvyBMrBaSrDuzZ
g58WkltmMmwpMhwSwUXEPXdhFRYvA68WjQfg3wU6t3ocyOCSSIk5ASKLOf/SS+GFsZKw2dTFtL5N
p1Ap+AcBlVBmmprKqXY1m1j5LNV2HIUl9fPq0ZnaMpZ7in5zVyiy97mAFNfSs6Gf7XDKKIMeXjx7
QQHndHv/V6q/nRuYuS4IP2pGq1TRl8f0c0+mWDnM1fIAXPHk1tnlhVeyp25SDqU4csL3/X7xrxnU
+ytXahBrf0CeMdB1RzfhtFF8ECs436v9+2/4gt1mvkJvmvTSn4BJSm498E1VG22y/3nc4PD8U4jE
e9aRF6t/pdfGYTSRljE8AlyIV4ypmgrPEO1i7XezAeXNLSTfivvLpUNpyw1yxM4IAXP4g8rV1C9y
Kjdxs3b8MxQaOBM0IrVLcqNdwP3/Y3r1ZwcbXJqVLDHc2HV0t+L77mRFW1x0Qw1cmpDdOG6KJzfD
YIghyEw+iTfbOLW7cUg+8KzDRJLH9gvKTFSmDp4LfB2rmvYbygKVT3XTKKgdBDDCO6FZwL/v7H+A
Cy1AtuX0SV0/QMUfF/qKVgctk8fUj9ntLrKZHVqXXGC3GkAd0LI2mov0xfg/0TbX/AbyoVRGcFbV
XxQF6okNwSCpjupd+qTLGx0t868crAodsDrBvi2+i0jWh4PulOoKbO6unOMsfAtJ/eYP6bD/x45v
kTg6gUsL+vIhKsqgxbC6ydbSbvgk/IuOzoGJoQs2H8Iuqcn8I5/44h8H1Exk40pZPl7kVP+Gqr5Y
lVyUQvG0oCKCr0yKxiHYQZlpBzBDddYIoiIS1Rn4hFiQsV4S74ZCLLIVyHxoDqDZjEtoGhFAKBlv
0hzpkLp59Kt+pD6AaBIjg7V78ZZUl1STmvrhxNAWnKKAkCSX0dUFFoPq8GusIXAo5BT+C6U3jXbd
x3oPQVmql2c9wOITPsMuoCPfs7Q41AgXkqvuYURcJN3ew7lxlZo6YFlfzuS2iMjnKq10boTGBGno
zfKREXCVdl3Pz5q3F3cB+XOZUUIRF1t8nGfFPb3Md4tOEG/jLNghf2ZsFAjrKP9bRbnbU9GjNIfs
AEveSwJ8pAEO5gqhWEbZw3eqI9q5okBwW4AzWUjB+Zy47fSVxTdGuudtoM01C9OZ0PQdWAUf2O2X
d3tT1mse+Pv73y+abnCoiZA/3/14ms7mT9ofi8JjTj3Su4Omin7UNyfxgnnM28dupmII5KNpVEe/
+6T5XEspG0yqJGtndcLtM0XT+lpUnbjMU5Q7EZXEr4aXV04Bt4IYoXTjR82rBidm3QzVcaY3btcI
CA+7fRBOF2Im5zFbjvpuxUX2/7kg+2BOA69g0ki+GDf/xmcke3RVd2a1oXt7sOp2szXWFrFQIWBo
rMZdFWTL1ZtzgPDTzsKmeU8FTr6/K+fUTqXL63jdUNUJ2iMV3cAOL+S8KXPu0NRGyI3sp2WcP2Qs
JmucRpY9j/21QCJH0Kv4BbPk5xpIcp1xx6FkEYzLb3LLGf96PQ6+/UcR7D3i0ZrBcUGPg+kpziZE
/H+SfRJTaMTm9H4KgJz45lLBFuMmA3w7PaFGdPxvtoGYhG9lIYlh0HnL83+8VrA2AIz8u90Hpp4s
4x+1mHZA9puugRvoQmstFfJM9ivPlfDQnqV2Nv0oUxfTlxf9JzrRFC3djBk8De09iYK8xhVs7WAZ
h25AupLnXA6TeDRqrie9e4tb4TTEWY8usIcUxUY0pvPDDqD0bVMrP/lS96V81horpZywzPk8yHNI
zXQ46V6UEkDMy+WOAelhD3J0hrV9GASNGOSxPMjQTDHP/jxeLWPEnL8nDCfT8K1ptL6nTskfTU9N
cU/v6J3bFuoV1F0Z6nHwJ6wz+pIx0NUL67tKe6OysuG1rb+s3SMuICgsqDdtxLAkhcZS3+w3HYK7
0Eag0s3bDEhF4e6JaWRJ9md8Mh54vlOgXU3KUYyOl0oarBma5rs4nC4OkPGynXYSixOCI9Lkbr02
o8Nvgqkywetw/XpVcBXd41vAxzHLgZ4EgYxaBzv4aocCe3JGWh6aAOM3PEqjl7ISgKZNoK3kQ1Kr
HUMK/Zl43x/hgfuqAKzTyMa4iu24+BbOwTReUsc6vy1zVVcUwYbuR7a7cX6M4n0EdEKLllqBX2Nf
WLEbgvOC9TNKoi1Rozo2STN/BxBnHIZdk3aifQTD8RWaz0w5qaGLWA/tn03IlBlR7wYkN+aWkKJs
b64KAXatFCo1P+wXOFTP3qmAbOE8KGrVCZIZiWnaCvSqIsP9LFzl1weK3VG1AG/YCwOxcsa9BhKl
UaH6SlATp5tuYBwl1v261LlFXFBvFUIdUDa1+Us1HLiXreaPu+2ogYiRACBPXIxTJs93w3XlmInS
qHYEk1wIBrgSSsSoY2vo4n5R0gpDdwSSPeuVspg915gRRtQa2n2KFl/E2DbZ9BG0ftSN+pPa7duV
3lexvjrtm2Wjd45opqLWqv9D1nHY+Bt/YazbHeS3VJBR2rRRdtvLn7RVvYLkenEUS4V5Qy863ZQV
U9UZ0h758EJPtP7KjILAa7+DkvAUAggMNB5zedJF8KnqHtEeyrgoiYSOIJC5wqJNMKrl+ZcZ0eUe
FuRzaK13ayV6mo2UYW2XuJPmpuj01D9rqQyl6nAqxs3PUFC29l43MO2s76sqfZo5jhH+tMz/YBQb
rVIl2IJ3QmGCpvb+yrkJXSLxhWYCfogH5AfZGQ3ajqStjzdrI6VuQLUdX5WON7ZShznFS4Te2ios
M+QbL6zivuw7GWXdevLcVs9c7fEEY8fbG9wBRooL0SoWX3Jmr2X5Iwq1CmS1KBlb6yX+Xs3p8R/1
rsqdOhkcBrNjHrnIX4Z85mD2XpXaYEcgTikvTjo5Bn/mU1fm6EOou9wfQYJnvBvO6pREnNPaZ8N7
d8qBGX4RjmzE39DT7xIMgl69MgXmFQLPjIp37WpHiADujDDo9J6LCmpA/n9d9Xy90T1LSNcDROvz
8wgNF4VKdpMhSL9c70YDtWwZTosF/SWoRdvYj7jxkRMW9h/kvZroA481T6JkyOJdlfUH3Jfe40Zy
WbTtxVFCzUWKDZ57WKRhi/8DzJSe9vtIoi3p+wCmjhRNr8YzrKFGn+QJRnFiqqPVFRsG63KdrjKN
QGWNvZADlX/ZYfG52nsGfR6zLMD1CCzxWq/l6mdwy09AaQf8IrdEiZ9XkNR/1L4g/HAf5E8A+ZaT
gjFztrKseqn2nAcBrd1pvBtS7G+qT+oS9SIvyNv2OqBfmxw1j1trU4+PQ6aztZ3X4unCuaNl+vPO
Df3OwhezpVGvj27WPlp7iNjJ4N68wAo104MiWo/crb2Rww1XvBhgFEmSOndPL69R12zTCWqg3Qn1
DoAc/RFmWx1rt2y94RRxvJmPbOQkFk0+RGozgnDFInRxIej4VCUVXIxbbaZOQtnaenEnUgyyuOLz
oT8/eGVX8vvm6aMM7OYpsStrf85dK84tnC5suhPeDPTGJZ5JGqozd43L8xyxzunOWQ0/CxUEBUaF
MkE/IRdppUBUquAGyqroA6df/KJhNKlQ5aBeHtITXnr27yM4Gy9gcd9LjND0LUkUczZDRbzau/JU
3w7HQ7V82eEoqsw7L63rdPSt/lfAK+SZzZSppcEh+vmAh4Zyg9oL7e9of0PZYlxby41y4Z6EdIi/
EyYtOclxaACmApaWrm9uqvtaOWCz1VuNmVCjcA+R8O2qAoeoujUA8WlK2qly9nZn1bgG6PsBd5V+
HQYS3VndTaliCcnHDaSUYY4IhNRCq5gw3vld7waccx8GpMLaxXEL43gUF31EewUgfgG5LqRuDNqE
6MF/C3804lzYjNwC7hVOX9pBVBGTy+MtR/urNbiylyrvvTbr+WLm3Tk9ZpPE03yKaWVE+mlXFrHq
iI4lmdeqbbnWo2Sj7lpIlC3FIRYsUU1A2xFn+kOFxEBQ7dMLDf+YVe79MVs93snMA2lQzzX+Kom7
6MhHbqDfadURo4J4Q7lHs2g3NrdxaFy7BNM465z8le+D75+V3xa0lw4pBpmCeTVCg2VSvEesBXzI
Vo6qUn6DZwQSpaDlVQBakgadMeguvSk3HZhlNG42yeeV51HX1GOSDcBWYPbTx8fwkiH0eme/8L+P
C3GH/lTtp+KelWhiu03G3yr43vq6UN3tswRKIK4he3bCjPAzeECi0RTo5l1A4WCrK/c01UKPTP+8
YYTVbCS7q/98na+pQBFMLorH8gEiA4NG3XEWA3a61hj1LJtsNSbvA77k1UO7FJA/nabAWNxnIfda
2uC0Dql+6iRB4oe29vH51Yc+C4X6+ZvTyA5XlXkabuF1wFF48Bq1mJgfQ/eyuHWrsYkK2UhadeFw
9zlZJiqi1rZJJ881THN+xom2pRvjPkK3xbj17pqnOUJs6ecH3+i3j/h4YbCn/gF+l//yfdHRXKnf
JtLrsuQC7sioJztdPJOPQesmgOOE5KYZhuWZ2eViqDUzorsM60MzUZsLP1RoVaFL2FcqLX/UWJju
bMl2vIiLsCqIp+pVggmMikqT4AFyJAOTviXtkOAtuykXCfgffDydKoPd127hQfGgUaPstOvEb5GC
ZXr2El6AJA13ZtbWcVVybi2MM3KetWUXpR9c4wjOcDsCdYnipoEUEDa7BSBfVcvTuod9cWLWtFk/
Q2A7nagKhB/FCknLvbeOuXCxOcAhwd3d1vH2LezJ49gIZb0PFzEa5YoAnQeDmZuZupQHOQaq1Vmz
w32dQCYVdPFrOg8cTg4oEEdmRduHfHTZ9yIdhbgpKlGsRZyr33C4aNNTRFOR1+d/+lgvtn4F+NFT
xE7KeX1ZXOgrP4Uf55GhlMquLVDRVzNrkM8wzXEigFKI6iR2fMLo3SjETwy1UDUgRB//j54QVkFs
ZohTgomUAMRJSjfxX0UCycjXNLYXo369QFkijHuy0o0Ja24vVsiqSRJZnMBpuF06rKWzCdqKUXjs
2zVyYlFomQCC/SN2jHJ4FMtqniyaaSbMiNa4PrFO2AfCe3uWldnzkePrKXXPoqM8el9fHdqOXGi3
HqKYu1qR84U/KQxusXXqjnkpntXiV6FKexjIP5STrt4WTNFK57XKaJQeDGJq/SNrTJhZqduRUDyp
CdwPc5+89YVzCbgt8ABpGmpTP7sHxtGN6NxbtAZbnhVNn0R+jibb7bOpdV6VRSgtot3M37p8ewHM
41jLOVAJnQS1DIdiXwLJhf9/+IpMHUSmahZns3XeI5FQnCBAWsoxyP7IHmkx+oVJCXtbGp4AoYpJ
Qq+xDse6o5Or9YS1wqrnQGDpN443uVbH8P9gi0T+IlsKWKPakxzKYCs25AmbmJL/msHENoPbYxFD
takpu2WTHec9z224fbUsa27cHaVdaTteO7JdsxpAVtbWY0HMZsY/zdLhw6r6DwRwYrQd6sCHZ56y
3nYmV7lDt9I+T2BGLBRd2LfkVRcbSJpJxsY8pgF/AFssIjAXd0e4sC8Aee9SfaThqtoHT74lfJhV
ySsaOPTVgv48BlGN43QpwwIcaOlqk1/XYW99ktGAJgjyBUHR2ixYpeOuJUazFZEmPAy2drsuAwQ3
iHsQicpiuUK1RdGwrRk4TNykARH8cNOtiVyZskt5+M+vwf1E6emhEzC24AV0X83+cWE9e5ugNC+U
on2wI00zRqVr9RWmEuN1Q5/o5XNv7DbCln8hcrytQv5uFbfz3qFTClhJl3fHrUMXXiNfu2aW7yvy
1JfdIC1shtDovDu3CuuHEuVyRkn0TEGE7qj/klBOD4I/9FURvo7eROlTDDdoM7R7vWDXX1RrywHb
jXz3cFqzbROBH2pd/JurzfzgiW0fF8orAEr4Zlq++mvGd0DhYe1QnHTw/WH5AO+HqjV8qDhDg/U9
Jy5xRBOkTg5xHXRPoAosDMR/XzQPXeZLIrN2cMu8sPCB1+KLp0ZSs/WzgiFT/+Y2rjoSSF++2D5u
UVToWLFKEUQKnOfMdok9TgPH96zduwTcWZDcwbBxeATtvKWrL59yoNB3nMRgegcc2tExBIIGhksC
tlxGj+1774M+KsNw/AbidZfS+1/Uswm12HetPDGkwF/oL975aiMFllD/UmRTOapIj/KPrP2E57l6
fLP1+PxKjRD4kixVJd+RH0PoatJN5stqiUwdBTlMr7xhuLIyTKh9Kzb95szyGs53HRXukE7tXED6
G3e7MAWsro+jSO4m/LbQC5CjnXpcmUiCVboBpT7hspTHdECDerB0KFq7950IWXEUvEO5oPq+Y9Oz
wHcbZmPBGlVuZB8T/OI1Om7L4KmNdKAcIh5sLKC3pYaQUngbKkD8jQZO7ao455V8V+raSEW4JArG
Q149Ggca90qoEmq6TirecM8h/4dGyPYRjZfTHaCAkgfivuCTagB2WlelZzAcdZF95Dx+rE/PFGbW
k0SqxeXM7/ONWr49LLfT5kLQ85E4hUus7MNgviHxB+m05hQgep/fds4aqybtyMBhFWkOEUFhEogk
QAU/tcEff1oYqsznmzg6UvH6dPkJb8sAgswHtNJw5quljvT0+Rrx1IkzqfUoRnnnzazXuBUZ5gUW
Xcr+apjgU7BQECHt4T3DEyiPlGE5a8dzMa1xr287YdBR8/diwKpTCoOK3uOQQOwMv0vF5IJkhj4X
h9zSiEBwpoRMR3c7Z8eISh64I3FwjQ6gQJdsChSDpqoAGJS6A+wKuybThKWp/Xf27LsYpuAnEkWp
0JK1jnKNNTQqfplAz7Qn8MM9F9ZKGSLyojp3O68yJXewBViSWqcOz6+am0rBtbF4XxFfC+Axe3u2
1+AspU2EzaXkIS4cNyVwJVecBNYl0JvkBmVU8Ty4XnFL+BGlDWmHdR/ggBDIiGJVKNXXVr8CZF04
iwf8s214F/pU19JmxfKe4Lde3ZSaaC4tsfiXs8r4x9ples3joQiGHUJ35P6uwtQ69KLRWGheGUKB
L7+BF0DCD7yYEn6ld70DV4cJo3D3d6NhWtsCf1Z3AhWvmCB9+AyHP6nGDdTmhXl+AzA3og9GZnoF
19jIs9wxXIZ+VTeNSxMiBWXr61khcesg51866eCGn/FoWhGgHaZbZzPoEVYhHOcHJlaobKeJ58QZ
dXSilIReJBR8LhMq1yxSExR6Cp16ZpOTW8FGzu9tqmOtEhxQSH4anqPYNSkGg77H6MRhrRRobkBo
Cm1iV9JjmUPhfs315nx0EJ07Rw7F5UFP91pqT8GIrWWXRmhwwenEdPvl+IvC8tNg8S8ZjA4HIq9M
FFJmRMYzY0p+HKwrmqUNofyWJ5ZDf4rL/+OR5npUTFQywDecEiKatwzE/7MT0JeT3btX5LSgsiqJ
go3tyUgb5U2IwLWOYY2Q3rWKhVXa7IUNMGHAy+ult1wcZh45QyTyKpnObbhN6Rc2wi9M0R5QzYrU
bEsZi6DggkCFK1oa8yB9HnISj6IcJkIcYHFserf5KCQdSuBVMfuMQroJJNhPMUojnVpdBNLpqMCM
My8+XN1xnoyzuQKTl3lLQyDiiYzEu8gR6UmIiDfAayKcuBQyc+94gLsimZa5STYEMst28YgRxkfj
+AuFIJV6CmBR8XQ3rJdXTsG4VIGVn8bqzW31HU+brtn87HMkA0eHzL8x1NbEUMwO3e/DVe+bhJGc
TV97BaABC/LxEaoeUV++Nsw7dBCfGSSNLCs/c2cfkgotivrPP5Lk1F5uA3QXh0BsfsrU7te4mWTx
MPN5av30dCT+vrtSCEYmI8KaxOsHfZf1EKPbfZ7v/0HZZYRpp9TNTYa60/iYFI9ByvPbFqLSWWgf
oNEdw/Vf/9EjOIIkOX9YOizT2URCub5YBNJd+IvfO0nSdnbTIkGaG84gJVR7tToaeU6qnpLOTlYo
p40WsUr89kYJUVsW2StNRXEuIEGZ5XznKy/NdBnFf0K/zCd/6Htbb0LwiUCiQ1OoZ5REakLYKgQN
ygxBiM0PKyBkcIYgO+vGeXCQ5Pl1BIXOX7DIvYFcpNIYx7cYh/f5OLAkEgGxrbEc2T2seOS2itqV
5hf3PyX1wxzCLwjbbBH/4KWK/9rKrgbyo5MbWX4+ZDGzbpuyW1HKWe/z0ZQtnbpVRM/hTkpQqaE8
3PNxbP/VkACU73JFSbdRViMhT5Nh9w1PqxXCV1xwe0+zxAuZK1MJeQsOyVEqhNA9uxAxeYhJdJcb
7GE/4vOqQ8zWkS56113cA/k9gjCMjocEdEHBubK4GBvrsks2FhGLIid4sxuf/GsgaMof6mOZKYEU
1ERCMTzL4gbEwRv+uUkllxl1gWNEoYdJpgJxKvyjAU4ZhHdPds3ElHsNz2LlVVHQZn6+9LLEl6qU
K5w1VawUdo7cwbSUx+mmQbUz068HTYj/zjP+KrZe7kYL5iwmHRxf13rLAKdgDHlPaXTXd6qg/k1V
oEJ52Xv1+jITnVnmhWVQxgaBasIRAc6PaLPAj6TKFEwt93iUCm0X7gFH4brT/jw+d6L6L+7S3hU0
Ud5+Njz0sQXBS54s1it5cEwbknASmhuL9l7Mj7GT4uiL3wMHcRValA9dfmVZypwnasmjnCqKrNPj
3DxOabnwrgWwS92iG/yzivQnTfD7iYXSoP9S6ZmBM0XRqFz5bGrN6eJhsYIYCJR3vfbSxgydt4lY
SV8dTPlNAQUMZuX0eZWophLRkqFcGE5U2hf/3QY/AfNH4mtC83I1XQnrqgqVw+6bMImljKJzqOnn
ByLvXCkFr1XKVtdx9Mt2+A86qwjAks5Cr8dlMUV4ha7ixu4b3mwHsqh0Dhw40xJ+tcqpQjGQb8a2
6yf0X4ltqQlffkclwbpPXgz88PnQOBqZlkD4EEGmMEaLcNaQlZoTVpPV1wtP4YRrqNB/D+hTLD78
IkSsCUIxAXCCGiQ8QOSwrer2asVCE72K8r9lg+DmErUy3iuFbJVXOtRtBz/mfwuo68KUykh1GOSP
CfzO0LQgKgtw+x36zMETqCTPrYEtPNWmEc4LAeWh03Qj1rjBIO9gnvZTshN96rSEpbbET/tv85SH
4+Go6aRht1Kv9jMsvlwEgCQQSjPYZ55Hu3WKi3Ql9akYPyZaijzTuqbm5XEwpkN45ycWINlMkVAS
GeLEGXWuIGtdJGI7jqFKoZsLZ8iknzv7OSBylC8quW4lVYBc7vNrroZmGxXbagc+O5ainOwn9XFU
pSzMarCr5M1T1Xu2aVUSqIq5/KK88i7q9bI3X9dtiFyuh8jV3UN6Ym9bEBKV0b9KDWUeWSYGRBk=
`protect end_protected

