

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eRz+leRSRPpou0Iyb6bnhB8hg9kPbBirrzFUAdKqw/be3+N8ZrhDizYaLfXqnwxlgZsSWJCzRfM7
HvMw/rTLhw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rl74r1iJC/bnSjzA+Rx4NZe56NnmjoVRFzUux12uAkwgT++rVuZ0cWQxVSY31Gff9TGn02lNxavo
U1xWF81U2u/Zi0XY7ZHmbpbdUEdpSv9huiEIrpuLuTgWjBSUwsGYqRxHLx1vq4vioRXFlAhPk9JA
iYodwxjKI7YbbZElfVA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lO1ylq105LQ/xiJNZcB3fPTy1RngsQ3yQ/KJ6FM1qs+SoXmUQjQaEb6hJLPAypYN8r4VdJAzSC/U
5nFe27DWNjEKmiIleROkH20okne+9N7+PhPIZQnib521U3SV/ecBImKKPYRpHhAeqE7OE/DzQFWx
10ISqR1I6WBii4R8gkz5k4dkFHhiTU6fgkIHLUXXclJrpQ6fHHlk7MPcpQDjK7bXjIiQ81qfpVmp
P5Kh8wiY7VppUj33GlIcYsNio8GAIV3e0kBKLoX73uDqdvJ/2zBzKOZoDd0As7C4AHF8YSixL0MC
djalIDRCSOBX8Rd9h057rIe8ZIXNMu/BHoKk/g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aJoUzTg4Ju9hNY+ZPcuNUmGg+rCD8aivgSTst8VRB5/g9QHuzghA24ad2z08gxWDFeIOT/HFgT6H
g4nDsyLlbHK2gxUijkJ6ORkRfGOxb8UwHTzLEIRJ5zmkHtJXYM250JOsiukrgEDT40HqdtSgre6O
kXXliGFm9MU0LwRby+I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ca/+TaSll/KHF7mIE37XMZRKDQpSdluwuJA9x/CRPHNmOrubSxRKoPtbXlxVM6ehE2hXp6yB6qBf
Fup9ZI873BFwgulDsuQHuOSUPGo4bBHwDnNbSi/4G2je8uxqj4KeP/bv0RKunNMT/FTascQdDh6n
SVSARZi75+ElUvhBfAjPHB+yugMvSxDk7TRPn1RomvNtW1CJTL51/PQt26FoAtnxmwYDcU5wo8WT
ATzZmP4jq9ClSvjXHkf/VnlLenBFunDj22Ef6vdvxByXWMZrDdZyqqIvDvktra69BBPdtD2LNyW1
FCI6v17qDRdmShLAB1bJHs4PPkDtQbDOwcgx6g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5040)
`protect data_block
/ck9Sd95TYG8VDgNIx6en3Ydm53MnEFasy4NdpHziXfkZltvDLrn9d7RTpd80juQaz8mK+H8VDxw
KJjtDTDhFgDzxp++nL3NDDkDytiRFWy7AW3YB9yQKiLkvhV9DTKOIVnBZc2bNNwY5Zt7uxSLl/Fd
YPRKq2dsK1nmpme2+gqJN3vOGYE8f1FM8mmmfsUyL2LyzqF/3ndN2ki/7nl+T6Riq1zPsAfwy0UY
iH6E5tRJTSkL1V/Xhb6+i4CT9pTHwqghVNeSnjfpgaK5oem9/75qOJjYkGq8zZgTnH7jbYZk+NvJ
7Tk7XeIWpDQCzKlKHhcbw4Y9W2KYwPrTRnkHgvHwXHccxtMhzv6U6h8Q0RQzMfys4suvpvISjgSk
WJRdOMys1G9jmRZqWx7OsqYWglGvxdW1uK462q7sf+RI7cozVR2aM2ENFHRL/750PE/fSuSjrJlS
poYCGEVn3SyS7I5hOXN85BfOBB+j7b1kKWz2yLBhsnfu8bYfdGtbBdt/4av5yqHABkrvK3aoiTwK
nh4Z7mKA3gmfLUbx7UkeLrFo7/27KiRA5+515HPpRsfuMKdSC3ycIGJ1qcCR8k3B4nz8EhELTaTj
f2GBxjJxVnmz07bDuD9LwIO6Y6bmRH/n3fAfCpYeWu/oj/yS7lrKYtoEkUbTQrZtOF4ZYdXdohhp
2bxkOwVBMkN+2Z41+6q2ok5VMl+P2tzgGZGh4u6t65s/JzSlhaYKO6NabjlMj9x6dsjBilF5A/8h
hcDpU4hCzLqY/5vLZtYV+QaqHgwc0CAbn5td5hO1oB9y8OT5LYOz3mcdmeU2bjUWbDQKqaM3vtIm
bIRRVA6NxrUwXalMwcLkMQTpFDSRfTyzUc/4d0ZA7Lew87/RAeRUS6HGQiRisaGLswVi0BKyQsGp
1sCpzvk1Lceiv2+FT/zml53yQJW7OGAJbpKu7BU9ZNZhhAwJe1ssrk/cg3Nvi6q6zEqZ7QpQ9DS5
zjHYh07Asj960YAkc4vPQAMBFrn7LHYRqbmq3n5xQg1qDGO++6UkrUMu2XH7oD/E2xNj/BIM9hzM
18U5V6QvhRsY/6XGwtKphCD9VYyVSPClSrDcJ6ipARe3ZG+IbVeQH4UNtqEAxzkwB8f3GbR2JHDx
iCpoTttisgJRnXpLMkLCYGc1ONw06/R2Xldvy9wi365X4b9JnwXPrw7H3Zp8DVFW8dJ/IcfjJI8x
7ssH4nmH7gX25HKQcM0WasTF5jw642egRNcCBnPbLgzTe2VwXOwili27lwkxQN5ZTxBW0+lY9Ok3
JceYVuVJ0KtA1VichTisdu1anrp/AV86HYhc7JwwI4i/ARMjF+3Bu+kqlYNt0gfYIbsdOHjCw/5m
HPOEK9t4mFMr15p8dZvJUtNQ/ZjFchIWYK/bnkVBYW/9N4pKfTlWnTlAMGhcpgTnT3jQlcvOvUEg
ufAHE0bgc7g0+XKv8LVilsiui8NLFFN++vzVv3/BMcdHpHt6Z6sA34odQMHUIhjOZE7ag9E/B/jP
6/U0f6mTqD7t7M9MggYcVZQm5epVWIAMyOg75vQgifzNiQoLoiZTK8SyY40sxsXiInIDYbcE66Ho
ENWW2k1q38Jfra+NqxXB7izYeEGTFCz+YEsDqRfvGV1gieJNYwyG34cAx+x74KUp4QsIOe+F9Hhr
9xaf4MhKlsSLu0xjvk4pY9sMBnAe0g9QJMlC6IOWjMIpcUW3dXJUn1M7eYSPVhH48e1rjhOmppX/
gXyINcmq+34z5MEzBzhWU38omqMeQHkuE4WkhDPT0lwQ8n8JfvjtDNjK7DdxHkWtIRW0AqUrl6JW
BlOqtDdy4sGLPia5h2gGD2wtZFhoE4YB55CrQxfpq0wwVML9ht584Ny6aAZynvI5RRTXO3be3zrO
1Me8ZTz+xyDGzdFtJWijlT5algQdKlhAcGznRC9Tw4VTj2mc9k4D4Y9dz2YhcnfvAVmVrzoC9rju
50/AxXGlS6rMeEGTnOetuh5WpBp/oIH4RUwaE2Xg6JIMVXSpllGdDHPKST4NDPbohUNLKDIQniZJ
mH4JzZnbRuHcgL2rtjPzZ5j7OJefBueKcm9aakxxIAKR5wVifd6WcTPNVpg6gzdcu1Re4XwONiIO
T2rjGkMk9Mwwd8aCduTnT4OsuevRj5pAcR2pGUkk8VYit7IVUbeaYEptFX32803oQ2EdCFgIU9Uj
QKo3WYx6a6u4Eg2XitMpHciNsA96kwHB0tsoWsS8ZbT2z99sROjFBA+F2EW8u0ASNI1QrQ8hvery
JvJ7+w2fUgv3j0FtiLA+J5/jZprAMUCwse369YZmNaCNKFItgpw33Bsjbkhy+WaDuJVAOfaUoCt7
PXiwJeHsyM/BRDlBxyR5y+5LCjqlFotZh/pgTsCuBKlHQgbT6Hk/eh8Ke7jafbCoDFHuu/71Q2KX
9WkI26tJIlXxZN4H5fkPyV04570fnCpzHGM/S7fDVJ6sdZbiiu2WiDPYjIFCIt6vyZvy/ZxilABZ
3OaLv9vnJ2hjlKQPf+zSTAhV/5OK8N2FEBhGbXvYl/iKDlig2HeJKAJLddrIZD6/w+xG/DgKMoB+
duqhNujc+77vneNEl3GcXbvzNFbuQu0fcoYnvdJ0bosNVWB4AutlJZuI7toKAbgPdfYpE7K3E6rn
PX8VaWWoE0UnaqyirU8KMtAEK0w7Yg/fWk/VCmovhDm7dEK1rASMMCPX575e1mo9HwIh+avMJs/f
82xQXwZqNa6pDrD9CVv/ahkbY3e6viDeSuqkKcDfFV7iKatJ46UYhpGjBMZGmtMay4MBDJufn0sx
UZdQMkIo25XPNx54houxkf/fa9+ro5O9W1EIbkSvKVvZ6psY6d+FVw5VRIb8foJsVoDza6sienDk
gxWtwiVByIwghO8srJh2nKf2pEuCyAUGTwmra9Yr3VC0Sn8KcsBA+FVs6JYVNe3GekasXwIQSAPT
d4QvTj7K2MyY0RMD3ZUI4abqDoL+tiwDjXjLeEqN9wIzKu/jEPLdN50z7vnLMeLHfY4FUkNSrR1F
dp1jWSaIzg0am08EXH5pyftPBEGs/tDnek/LfprWRcFXFUyDlUNzSTOr+pjVBi6gI/maKc+Nvlh5
snJSE4aRqtAKtYPEAxy2dP4zMOjx1rwIA18CyP0gD82RMYBH1GSTkr7qfOmrkEjlzdv1FbQCa+vz
y0sZSrjyrbaYqvDNO4q1icdj5mSu30VWd3p9hiw1b6LXUCakt/XadJaPasErS2mbp19VQL7u532w
hXvCVsDxObYl5MjnDZtsvjAtFTPNzmzHNKkj6dwiPzGE5KsfFleROyOEd9xZe64bpNF9cTLvEYGS
VX/XnxGrt2kJAfQXyhgwy3pTXzbL0PqSGKCOqZ1cHGjW1hkqvL88RESnE9vlC2UUq6X3SXxBUkWA
UMJhhz3VOt1bBSKMLRRMhgTaqpbRulJdckl9o5PfW4YOvhnuLvHTH/AZ3nmbFl1f6wGA/aMNhvQL
FCuOpKbe8pZobs9x/2XetMEHGTDdDw760JBTRHBZgFLzjkoHMdjqJVx5LSc0Jc1QRgfKIiuKb8Ao
770S9b0ACo+WHXHEh3eMcVSV8jejrsM6VaKjuAERwTAuuesp3TeZBV6eGsDMiXjLA3GGdiauKK3+
Rpo5Avck1hUyz9cRWf6lOlowHdFhv1NSk5Q31c2FOGWrtehxQDBZyQmQK3wrNmjPT4G3MP+Pf8Nm
heJ8FwfBsdEuqrzCKllXEgyq6pIURWhJWQ837LjlLQnQjRBh98P4ldatMTx7VQI7diFq01LrMGzU
llFDBKnNMRZEWhQi0semNegOiz1OH1sfDAqxKWeQR8pd14TVmyf8Ld3P5Qnts6Sk8A8IzVv/b7bH
5tfwv85birYGmG5jSuKCPOhs48cyJVzZPslvmiwo7/Yjyd5ZutkToFDGYZ82MuwzvWdE0UFKV9ts
WXKaLvc2EkX9Y91T8dPhQIERYC3cjud15v/AI0KhWgOf/qXUBDWatfutHyTG8dG1CGrlfwGX3W1f
i6UGg4dwAt+BQ8FNa/WHCqXEcoTmyxOT33SOWo3wdB9+ZUi7z88HKjy6hy4gKuaRXFAdA6zk7I0c
QMn9HCoJ/3XebeTMvoXHSfuS/rYUa8ApEBEOxrB1Dl7cpp7FvbBv4mnF4yWBdnz8Hb5FQmohzJN/
XHpHd+WercTjfx/Di2IiqAZWxjlHvgSmXKdJq//KLOp8Pk7kOnFoNqWbLRLEwsiXYSsXbvYHCTpS
KCiCbvEevRBhhVtNZtLPvgZFblxxvPbWgMr1wvgXkHRK8Tr384RBJoNJrWNjfjkdDBaM1iBPjtxX
/Mh+DOGmLIhhuUmDXudBZ052WKOkpbhm7IwiYjzjO/iZEf77+XfM1mvBthgB6WbO8KTSdygVtbBQ
XjJVn6++hF9VuJrR1mO5PBfYXuaIpp6jmeCb5m3hWI+mQ4Kpv5FD9WWniOIP/985x9x/c4rjCT5Q
cYmF4ErUEQ0Lpk7MdKYPYUcuh0J5hvsMnigS/Y5a0bY82BOnfxrlbLyN74FQaF1vqxEcC83tThpV
70pIOtQQZv0zDR0bxrqRJ2dzPxSHMnB7cIXbF3L0Cf0a5+IJX4JsToWzwg2oNw0w9GidFkIm/wc0
sYp6VF/26p6IINCrPXGS71LPltZKZnRtoS3pAhu8PipjWtDMgT2lvwpocNlGJcpmTmwQYxHFg8k8
14BqtWtQawnVBXbynCO5zQY36Hwjz705Tvf85RBCV92Np/zW1GmqL1Mcs+X7ntExYy5hdw0HCLVF
Xo/kE9ozItBppFQUDeWuigKn+svJkt6POLxZ+xZc4t5OwiPrIUMBnTWtoianyDjAslwrGONpVsl2
JfDYnR2gztQCYTpTSgLzUm2rm5sy5PsSZ3/EntBKXLewkDTsmhbGEXyEub7kf7KX5TX+nPwWet32
xULsbz4O9c4F7ZgEtpYnT9OprF6Mg2glYmEGdIvL8hmKscpa/gSkOlDIQtFtdhuOJ1mHDsbAg0hN
6E8BAhClaa1yGJ2upc+JYVjpY4pp4yi9Ku3Le6H+I6o9SUt24rmdGYcfcUymrfl8+dQhC6r+1Z7q
+HBVZ8mYL9LhI2CKI0NE4BYU0GAKtPiF61DCFAXlQfDFZtWZu8llTdvXNUGPJPipitpOdmKA2azc
mdVreWQqXSMCOrh0ukXpPULnx0spubKHA8Vzeg90eoYxYzUnFHSDNTIOQwRILvaKxfgaUioilhD7
19aiuOLR5rqqxylOlc7n5GMja8gSJhdIdVnDzTNLfEgS4TPXXtSMzsQxE25JLNJFEr0O3dAzk3h9
vLcLOKegWfXA8zO0TFNt78GYhPrWiFLdXrcOxphCBdQKy1QXAlRfU1LCZt+jh0HYW61TXKNVwSRb
q1hzqh45yXr4DuKKDC1JvfDni4dCpFw2DkzUiCEF2FyDCi0uE3XgguwRPo4UM67pagAFT6Otxo3i
O4PYP3OSgNyh+ZvAa3THETGW/p7S3PV1lVLml8F+HV4/N43Mn/ubyQxWCLwbuZhhCqUk5rMaOPqJ
1FzNck4/z2NJsUzF72UX8Foq+EKRwgt0JrQYi3yH8wWIh0fXxlm9h9fepJ89QjYtM7MNtmCA/zAt
02u+fG7uKYJCSReJx9XgUKfHZk6HIIQX8ytgVQd84lEwNnhqh3YzlKlVu5rtctXaa5LZps+9l74n
ne/j5TqICzOqKMMd4EYwUKK2/rKqtrhb3mSImf/IPtgcSZ/Blojhl/uycA+R5E13stx5APtgb6Jw
tomIG2cViW5MMQ+C1hccj7LmkkvVH+9+5WAGTeQiNCzepEskWX3qUwfI8PSvXOvy+yYVbSL9Hqds
MvGYTJQS09hAyQY8G4gn/p6D4TbQEEKNMIi6XkGWyWMkd/ZjzMscyrgETM4DCGNQlnYJ7Jqw+uOq
JChyZ9opU2CEPNABvy2ePYe4oKECECnqi9kEhFmaCiaLLOI1+BW0vffdXkjrUj8dvCxOiiAFmlkS
DebXdiiq8pYP3zAeBkgyDjyffwN3TvetZrpBLH6mfOHpeRQWwQhwQm+y4bf6SyTbkAUqNUdCEln8
Lw7iKWAk5V45YTobDt65WRZNhlgJK+d+cztbJZvMnIzEvgaax9xnGH44Onpqf/IX31izKXZaVDql
BfiZu8COjzWhWHD3TcuCg1h+YwhKHrHmLQ7dAEHsnZCG8UIiR9lqOWuozzD8DVT/KyRHa0Bim21h
312Wcs5rmOhMTIZFMLpa79lFFvNHXLCBWLgTTi5QAqQ6bLvCJXpD5GR0zCIITDeyTYwMN2wBfEVP
fUuA9/tTiSIQenAgyEvyViLpWdvSkeSsjvl5KXC+tG8ChSICozmvOrGKTOhPI4jaNjaWe3IH7h8g
wtsVAqHS1yMJD1T1YRcTMevdt6IzvS0BnYaSEDG+q9rau00fHI35MadolM1IFlwezZ7Nm0bqE+9t
FepcrCAo5MIjMxc9FJ1SIs3sV5gulmbqEJrQHmDQFoLn9H0Y2nxiGYtqkdGs3DqX3IWhksnut3ss
qALDnKGA85D7rFDxaZ9OSbN1PazQlnDrEb3C5nN3/3M6KG3SRsXBzEGnAnS2KjDPK8/1T+UV9pHN
CKI2UCSYExDCaUiSF/N6+t/0yEfxziOHRzIerlvCAkGMc34qj/MeE92V2DTVzPUmEuAJ9adth9VG
biY+NZhI/71sf92eCUyDU90PuzRurAaw
`protect end_protected

