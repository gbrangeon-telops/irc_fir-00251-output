

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VInMykl1cb/eyCcstyHEIOqfXLtsMYAK+iioa3bPNZdsHyKysw1sMYrwKEQhbdDvFZxexFV/BuR3
E2V10xNsGQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cUXIMbq/fNZtj1t37ez/ki7n1ShEuWgIH8yPxJTOO6Au2Dmq6/c17dbZtzNOPZ13Y79JsIBKn47t
AJMl7N429e8DmdtbuhhwCbJ38cBiFdxfH1AfVZI7GGjMAdNcJoTCbcfH0JfWJ/S9l4OVfdRveiIb
dXW5fh7twSl61WcUJpk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WHbKIifiSnVyh9VOrHbsAOJaiYfa+g3aWjT672CoQFGtZoHYX7lHrwPeDjn9R48BpRkqqMyy5V1E
kZ30rvMKCifKQNzf0TevcVrl3t6QqBIPZj7dsFAaWjY+3fu0RTcnya994wdnAwJ92k/2t3MWJiFL
8UCO8DDPNY0Xt40qfK/53oP7zxzhOh1lPvsgCruLCaYCAr7BplNWzKtgMfwt5ZUX5jp0hTpI0y3m
TFH3zhFRvsKAbe3q2U7sLVIx7P0al79lRmHpf3nBQ8JKs1WigNl/h+LWFmAr0nyU052Sl4nQmc1V
27CTe4+On+Y4xMsv2u/myTqMuXN6bcLrIAsu0Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xu9pS63o1o+cY63azBQM+vsKaznHACPUqoNT6W0vN2jhydQX/sdcqaY0W4LMPjU8g+1LDfLNYA4a
7f9gcYfJbb3zaKr5Y84jP97vWDuvkp0JSopB7FwosaQhgC9ZFFZSHrzYGBzwuhbZMni9A5RqvV2b
bQteOe3Z+NH5ROjD29Y=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rwUkytz4o3nSG3lKXYNGBGGd6NQin1yD4vxAFncd1x1HAH4uRN/6Csj8O1eFBSdgBZrbzYpSigyS
irdheULjGWq2hoVKG79mqHugwoJaQ+RWNnILZnDjYUeFGEu0ddu39e4LQ3yMfBCfQxRQcGTVly4Y
EDooxEh83Mu9Wm4Uvi2+2y26u2oEwtbjgdJCVoicm+J7JrH1l744lVTCHFaZPWdZupXmaLsbDTF1
IZL005EF99uQ8TMXRMkzqTgTLlajCuwvHoYLTNcLy8P1f7qEEvcak6Aw3luT9m7/agpHKsss3X26
y4VegtaqqF/A90Z7VEb2715YgMpxzFEM2FzMyA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15264)
`protect data_block
VujVyW2x9SvQonwoKWUty7uFyqN5jrQY5cD28rPAonxCSZIdUjdruh+OXFNN+Vi4AruWzZRiYM+V
VF3sHvx7DQTKPbzc4ZB1Cl1xFT/r5LGWV2jWRBOqKXT7koPWhvLjh36H5VEEJZCeriu2ENu5H+GG
DlhExbpKTfAf9+3xMGoPa4lKQuK5ba/kRubEBnc+ASXLUF0t32pHtUxCv0tNyP0ymLzTTdAmbanX
yNkmHGDCtmjXP2gp8amS7bKbg6Vd04m2QISZWTBs7kKq9EZqXPjcC5S+3jJEb9wjXncWz/G+Kym4
egQso+wEPmBvFnD9yGW567scteEuIEFuf2rxuDzW+nZg2r++Vp32haILUPlNLnCHSN9ccN53tiWV
JdycCo5dxqPrlXsxKWMruzq1pnHdiKCGsQkUYrnUc8go2Wg/JN/HPuEU7OqUXe8GtyPt6rrFI6aM
7TXzusvT0pWChsiE2Uuyb3xGp33/E3vipXsQzz1xubmymlsEEQyDDr7c+8Q8LUYAJgzqr+UPCNLG
ZynCHdP4ugEfZyB6hpHwmbcIqySOe3lkLl1wFv1vNV6LIWASEWzGJ3IS0E3nHpDU7YYP0JCfGq2v
8Hk6ENXL+ZyEF0gMZWnCxNwiDlyuIFtZb+cqnyQl9eglzcW0L7Ap+m1ON8DOjr2W7V/daM5oeR9Z
CNa33aH1lmbXeryswIbFkxd8hTFnt5jk5V1j7o/gItxWHsCCrSTfA4m5n7Fn2XoTeeX7W0F6OXjI
6RDv1S9KCJlgBmnSiTnAaMPDWl5hVC3tCH4KbvOaZ6202/iMFQ0tPVqFuF4NpzpJ2VWLfpFe5qtW
Yug6O6J+ni6KjSOkPXn0JWDuvrNlTWNpKo10iYrZVGfVVfIi0MgFrKanbETycevQf7bBp1Bt6NWq
xcEqWHbuavlTKOfFiNoehVNJ6Ad6Si9iJ3WT/k81LYvNhQgVcIHtk5MWxwdXVUxR2F4VX3gqg5W/
QEe4D2cGoSZeL5F8IgVIYHp+OoED3powvpzo2JJcagc3Upg4wY20lK4lnPK3+fyMoxbbNnIANa/x
NQMyMMMQ8HZAfxvZ/Aajc2VXhfn7Hz7SD9IfjZRzp5tfBiCWSVCZiCP5md3g4B6yDOt8r147tizq
n4KrpP7LpKcLkwrjp2/MpSbes3HJh3zdC+r7kGF20jnW8wXWHVjsl1I8M7cWC12R83dIP8w4viSu
McVXEcZsjqBBFiZZj3ixOcJJShwIVqtQJLP8AmIW7ZoPlHnKO7MPLbAUPm5aYGdGhLzGsMs9BXFs
ASDSqZw30+luSIFmqRuHLZhHV/6nSp8UH341xz0eSRKkmUXRw7q+luiH3HWgzgk2ZZ5ZwmRZytKU
m/0kPJdd61MWTlFHWkZvQWsNbgSci9e7rWR7xlDHwNkVHChFFXXXdRyBgKlWSrcTFszOCx8HeQ71
Dy6ZPIwRFlfBKPqUcrA8wPtWpE1C1eI/MOihEkiRj+oRMSUIwY+5DkclHmGGFFCSSKOBizELpT/D
3y4cO4Z/Ew9HAK3oroE1QPygth1wsPvcOkuDc919o/SuuhYROmXC1PDzO3r5+btX82MRg2P+2ilH
zzEm7ea+FjIdOeTcStytZ0edvBOrU8m3a4fK8OiEuE75NCypRQ2ogLVuwkqv2UMrKEpjxDIrVbIe
HOjiO6O8Sd74h7EwrLFkWUYIZX7sd7+lp5K0d6ZjT6K5j5C0v4tjzvW039JfAnJibEpc4OjpYVTS
imIZ8fDEk2OA2iNVuLOLGXtfKqPBX8WQD9oz4t+ePztXT4Np9E7vlIGy+L4LLajP1QNKncPhFo93
Bf1nXIicvkHeYorrYbvJy7RWtEE3gLnRuSR68EzZnfBHLvXh7AGxMGJtxTv/jdFAhiGVE/UfuGgR
eHGfJU09XXzYAxFpDKeJvMqFuJ99Prc0TU2kEMt6Ma9h3LOOl7M5ZsicPNWF153QIYuEJWB3MAbQ
3NHYapcSAnEkXraG6HzLaKGNP2CvZZmnbNyIDDsFUSgSpepuaG3Hsws0I4rF4zdEMSDv3tUkUO3+
YtwugTGTzbI+uDaQm+pOvMGfuyryevXGsvow70SnJEt8G+KtOOtRxe9f1YdRlXp6L7n1q5KP8nUs
y86hV+EppZLFlF4YHfAfe//gE+lbOmKecJlEjkENjP23Zad0Tnibyg4RdXme4v28KG+PRqVYrQXe
cdwjXDLTBjqivPLdj7mIFXY1xaGw4mE0dLLaRKMPIWAEXRa3lbXg3urfr9vcyIRF5sTDiUv/KeQw
2ClvEzJIVDbSZOGk614MNeK8LIIQ6eNqXSQdfIPqdNu9hCPfOXobH8qjFsrv+RWGpGC2onidyfOw
CWMwsTPoBZG/J4OtZu2svWOteTzgOzl5ElAmEgxgv1xhn4B0qsKaR/OoIypi17JxZubjIsdeoXzF
hqDuRUIj6RNflXLTnKFjJ4eNsgZE+rTpqYtccv/mdrvadCEW6Or3d7xQGZzILUOXfVwDM2Akngry
Vth8AGKEd+CzEiZtzHyMi/jTJBzB4TLP9eHhbUqvJbUaIjS6ckcFaRZuJ6i4IxPkTwAB3dmxQRo7
dkgmRJpDiH1EXNj8sRPON/3opexTkRHNmB6zOi8fw+KmTNjA0Mr4hm4jJVOjs8WeoMiSRzftA7fM
W4TRo1NATyJG9DqA/rgCoJ8tcbLEFqJdwGbZgMT7kK8aVy0dJzlul8cAwQQu+v/0CLdVu7FVUZkf
6s1oxpxHy7pRTEMwDOkRIoVy1k9qDSIK4El2DY90tpmP6UgdC5lNUDsfyimK40GrFfS+jf541+lQ
8+tzZF/PNGOAe+vAAHgPJanpVhU8+uIhlBBcwGHLQXzlsgzK3aMMr/Nn4O21IZwpbsD915qJMbzG
gu5z11BWr0i7HHJnnSGZqrLm/mwJ6lFEV8XNl6n20ITXut9mtf46TOpy2IwAURDtSVV4YRO4VMXk
JkXneehQYMHmj64gnk/1FPgoW3VxLi+hjavCTu4PDvZQWi8qGdpgqobX5gYsfuElDXEORj61SuQA
Os2zYJHrlmzHLJZnVf9f8hi5RfNRDErswkfG8m/0kXTZGm3JTT/QcgE585KJOgcnrrrStNt/XQ0I
tbfRWh0tJsqxxpC224Q9DLdzSOPd7zvAnj4SSrAd0/sTXNpoKCCbPVOpUAWSd2mFxA5MjZQbcVVn
JjASmPwpo/qZY26DN9S1J8R2qREt9rc0iI9WROV6dU/rg6XJ4WNf1iXSKshJyMOjgOf4hE1Oay/C
rQmjYlOGmivA+v4nfJ2IGtFA9yzBrnnqkeTQZRXZnO0JaLK9YEf+PlfLOZZBeZUARcwmQl1nw/Jj
cClSntnoqBJ37d0Es9u9ItNaIkDex67ALrtfJFKt2JHWy4rz1YbIsgl7CBaEmV+SPRZt5lcV2sbN
EcVOJBgO6KsedbqykH2Rg7j5I8EFu99Wp9j0zDCFLE94i1QQkrPIt3hLK3fl/vC2dL/emXcwDj+o
nwHVNQ5uf1GHbDVBrV0SyY26d7BuvhdEtfSSEaKVgWW7q2bHr3BWMbVG0z+TmsMstfOUps0MU2Y6
yeQQPPcUfm1oajHn/LRwaQDbt8kBM+aNq1cLd5clKnkh1mpodgdWHxg7YxK7GouDmajjOYQxc76m
WJvq/0lpDXq/Q0loDlRC5NgGG0f/ZLg440XoW+Vwfa4as2mptO0O3bapUztwYO1jsuynIvOK7Phq
u1TAuk+13xdFylZbcZqMY0Hv3N+TXCZROud4Z3fTwnCv9XriAZR4/MF8/PHyX4DCFsVvO49+0n07
K23vvchGQciV9EhEJ4ystk4Tnn/UNQtdylfCMkNJ9SYOyrrMsgR2rnA8FPmQSp9y4ts4kbtn/koL
RuRMi6oFEfhRwhuMxVvoBmGu1FOPyPP6UAgv9nl1bkDxI/7q+IPp3XLzWSKCoQCC5zdrc8Z/go3a
F6hsOHOYUXIGJJaG4D2zSbifP8iW4GPmlF/9yiJ8JF5NY2OjgpBagrtzUDk+AHm4MM3EJGKKXI4n
6S7HkAgigYndf8MEEUb4cbhDNd7eu7+ZI1KKm7T9J9+vDevBlf4wUd6vNbqSQbo534eaHrjgoIf4
JMqxgD11XtDSzxFnlcrzcvrnaSwrxwYa93mtpvYa8N0JriaCDes2Qs+Z9qkjnTYCTm701jWe+ynE
Oq63Y3dRqjtDI5Y6tMIv97WjHQ8f5jCiphL0TVJUrCsicb9O5WG9ZnUgrsCxO4yzPU/9mfpQKFUF
+5L9EqQtDeOPIuLNTdfiBXjUIA2TwAVMGNBRwrpzq9fVWy6sZ/BTI1DaK8cufvz2MmCS0ilnldhz
AtCj3kZ2+MaLkyXC6iVU9KYMkCXhlRdem8sBnI0fw8hg2yj/KE4HE/ZWWnP1moe+ery0STDKYJOs
o+1rISiGBw9O94ESIrS7NALGLeQ2Yf3IQvIFWzSykuukllkB2xqC4AMxaG3Mt8iS4f2gzDpmjvSg
aSOp8mS49Xvl7pDXILpc8uKZXOlVyL5jLFRdS0R6I2V18dfWASBNX2453m8bQAMb/2siILgxp10M
MrG4ZQsjBUzRUapkOW29bU2DS510c3ntN7KdU0CbPbIZ8u9NK9PqmQZnwOLOkDmqesOSH1feyEYG
XCAd6fpQ1kekSOu9Zy+gxnnuOhSRC8Mu3UlNKqgPWd37i6jNoHsVScXbdGwxw0EJERvn/HIAjRDC
1IXsvCiR96Oglb5m3Ww0ovTcVouKsggjbATqaUOesGiu+T/XyMrPaSG0oFCjlkNXTVSRyHhm4VOl
Rc8/Dwz/cMqA7PuxvrXkGdInUsdYV75m6rMaZl3MCUVNZhWxVtLYqqgKkw1gCzWEYmtuhDQal3h0
Nz2vVDp822QWyLqhy10BKKYeXbjwt72Jocr/DUciZ8heV4gEnt2AnMAKDp4nsgjKTjFYjnDjc4RG
B44D3CxjEexUtYxuflRa1dDXUil4ln7Z+VnAEnDLb8uu5R43mJOsRxZVU1b8igCB44zqLSEb4tIw
GQOILi9QepE9FzmSCHPn1H8MsgCBNy60hjH6XHmDAxmHAlk5wOzf/++VDW9WmpU2ajKXxJo5yEqw
UIi1I8U22TIhI8s0lrN3RJcdxe8CAdNWvkHnz8ZIrWY5q48+xCOfgjkyDDi58HLdpcxYKRceSRj4
frREvYaZIqsyuD1/vnsdJAiKezdaSmmBA69eX3s1zF2+0Ymq94QcIQc9sD0xvKq7oMv8rin0Q2Sj
mbQU9WnNzGUESlm7eZUxiz0efCUSplpTkfBwCwK470lm3IeNN8xPIQEcEjO6BUyINukSxoeo4oHc
jgQarFAIwg7V1uXqFDkBqkXgZ93tswZZTLdxxWi+hthfk9ZRgZ7rLMPs3j1JqwjTll0ebtY4EPtT
/DhUlltRUjg8eqZbtcM9GQ40y3dI1EKnNCn8lLNhyAYeaweuOl8lxl1jIZwyZlNxUPlopk3wfPCp
a+fpB7x+Ag59iJgGmfvugvKQh1Q6JvKhBA98WrsrtGIieCaWke/odd1cq6H0nBJovhUQlrvhdmMf
5IzZtWy4/xrRf+Jd7hP+PIVX2fF1qs7U0ezuw5oLsK8ziL7sdCFEqmHc/D1aZns78YjHHMG7AzyU
HxN4zcP8m+/xoejwpl2pMLBmPVTYHLM2u2N/WRQAXDr7x0snNHZkbHPKTxo5jmXebvEUXkmr37be
OcHZQ2o4X8IxfhBL0WpnbX9hSaXSYbmA9u72LqT+kE8Aknep0nqQQXlVkFouXOZ0VjTc0spz70e6
O7IObwyMXVkFGa8zf5QM2GgiSJZ8PQFwClVcaHO7cqIvGkyQaXkVApVII57HfB6u88qm4Bicfm0T
l9CniT+tfbaGudobj1vxQL9nusZQMsF2ONV65aR1b1SnMZWG2sB0ZmGUgZIei0RLVb1rBfrMs7PF
nloqlD8b6Hs6TSdJmVPVqxq1ZAaTgVOFLz5esveuWr56XSSiLdMNxiR6Sj5tK3s+zq1Me+zlHRyp
u5XsqE110LDYxLGibccAJO+sanxGn2rMdjPGAWwG8f1WcdA3qcf/mr3SxUQovY4Uc5v3VvGAq0DB
qcIckeHwpOov0eUBVNStxWMZxrf5gRje5CI3/sVS64Py9GI6Gjsh1MvWG3FRk5s14SUYE66UNTrA
Z6RkBKsziwPk5Oqhugv6nas6qxx6/1PpnJlp1pP+7Peol4gcK4NNtEjjAJkwYhVUhFomkOCb8ZlH
tb9jxZmOqml5IeH8Gh5e1Oa9d64bmY/Z8rxseB+KW9M2px5hyEbL/kZz+d0hnTX29NptKGc41ZcA
4zx379BHMwKqTh+u9w171Ih94XpoExSuZw60m0e0JunSIsGZ/RQ8F6dAOqCOXTt09ARB3zFEekrd
SMj1TaWQ3G2ZTyhWgzzpLX9AIjkk4Eh6FWoo9OHgVRgBZP3xKf4u7hro1WlsIhUnqpU8/ORkO9so
kUcmYf5E//B/J7k/pe8AgvJn0Hpe0X9pV3hfJpJxLF+vXYseqLc1CEVgQ6XXkwElgc1JL3VyOEUW
qtPlQ8PWwa0V5lTKwPpqtNs5UwQwz0wDl8ax0VSJoiOxPC++dWsOFfpse1VlISx5vRF2cPQR77ay
HnMGPBTMPjy+ID6y5aD+QK8VjzTkhHfLpyT3/WjnIJzJa7zHN0ptDhn9Yl1dOYgf7WgIabOCj7PD
JGvbe8zPbGPqFRlha4BVNaAxT01aziqI6fnemvsLX2CQPpEL/NKr2hxRGIpxT5Nk+EremNr+GWoh
+HsxL3acrrYkcc54d327O5YcpVFRVbExzHGMnQrLW4iOchw78tChFU4dsjkJ9oYBQCrkK0RCFalw
8+AH2+RUP0/31o5mEWTvD9FU+NCT4V04uU2L/dKT4KgXQHbpveZxBfibjn8Bz2hKoLK1ejylnwyf
1QO2y88UisVJlfzQXnz8DPlUYCl0KLaYVFF5RwBolXHrccn+QsjT4eqbfwTpUckO3iaRHK7WDt4m
L63jJzsiHjaLCMd/59xcpfqmDoDTFOgZZswNEJKSxremkXY6AytcrvrK6xaymMaJiX0Sk+h1nY5M
8KT0BR5YDQGwq1TD4LnAWAivA3nx5KDPR0+kv6S3guo/IzTI+SYCEbEDI8piElfty28iMb5/WIoS
RxMFNTwNJNi149CgTOVAkkYx9OPDltDTaNHXmSCuTWHMQWE6oBxlfxMOFCJMR1Ftof2X7Ys6ZmdA
tBvYRdrf5pErD8Km2nfX/rrI+k/8wJZD0PNpzJMclSkTzjqdPV4MPLWXET71h5d+O70ULa845uVR
QPMJn1wijAM3qyZ0cZk9luT7tflzUwPXXRyww5W6ekxIDYh8qU+qbinD2kETrQP2t6dcytG8zgws
u57boqlPxYq3B6mW4/G1520I8OcxJZqthBWcnTP1f8JhqeKZW0OTYrEbbtd68pWd+6mv3jfoOM5E
7eIby/JeP+teX8QMAoPa9+tjTXWFW8SJgTTJ6vUOdn5Z0JVe9W2AUKUHBSJuFriACj/bkG1+cEzk
KJCeDkFgaIi9T9cfwTPybPOz29otV42lW9KBIdwHzdTZKceaF5l+eLnQoDRK0lFP4vOmBgQsuG0O
AwjhJmA0IXBTCXkkStq6HbQT1uCJ9z6mRfpRONKb49YOnCA6fvLpxdpLMwAPuKh7Gkt93JqBx6Fn
owCmhHuA9Cfk0+yJbksPLn4CujkSOUqP1JhiJddw7d0aHgqmdcORuVKNuFPeZ6OaWmS8aqew5G53
zqXi7zHsudh1DuonzbzMZK9ZfocQmAUPpLH3YR3VAbWQwM8un5Pejxa8GEiATRym9cEQITEnuITT
0FptIlZThOuYRwtMJWLTd1iQinG6km+SqwYc0hi/snSWiU1lxgNg3RetVwf/XlOOdCOSlAOEFYSQ
RWJLc8a+KWf6GM22DA0o6Tmyblug1Mp5uu17XGSL4WT4vc7I+HNfoBURDSKAfQZGPlzDfHdQLID7
AIYIlwJIEAgVlHKGHx1FLuCUarO6Vhrf8xPeC7ZjHxmXnVBk8+HIGslFpxRrm6qOdk80hWX00PhA
dtR9m1ruWEU300oosQrcpTdLkYTLHXgby0FvCq4vakxjp+E04LCMag3d8l32gFFp2xRbUHETv4IN
M3KTGNODy3xyHSpASBJd3buD1gMo/2ebMnB6bQdXhCC3YL3EDPY0rY/EBjbxfyU5I/G1DZe1mIaP
IUQi+XLx2QKIR1R5D8iTBghnL+HPPwulxLgKDx7cJEaRBvMCb6SedFKCAeRPzRz29pfWv9m8jogt
VrPF0vQW6w88XEtZ6Fwt8B1XYbdHVfUn8kncMhi8nZGKGdadbfGOz5fhmPIw/ThUKE0B4h6aJKpz
AxwBPi+QUZTL8pgCsD3zq9EMlW1SFC+ZHi70LQ6DtbWCdquH+7qOOozv4giZZ6Un3FUSEm0TD/+e
6uO07gaxhDXFBLk+ZFNozAAFBkjWAochfRthWsDhH6pDsb/O4aSJ6WNoadiLL3GXg/flVcHsx4Ug
j3pVHQZr6MZKCjQX7n/tGzOd1bXEEA9y7CId8KI/JeL3tceqSizsyg51hARaln/GK7ohgTtK5Hs8
09PvrhO1zl7p9Ch8t0EX6JYGea4ZoiltBFlABY6IrSaJ+H7F3gRVm70O2qvcTrZKdjBXFaqt/hRO
cWdKVDPOk5wpSJgiE5LcJ7Vu5aMQoPGjkuZX3o/v6cK+/IedMZuMC8INBgxeTslRa2fJ4Ldd9da9
9iDVZC723qMnUxC/vU+VeSnJl2r1VnciSKZu9xT4XMv5XuoeJxCXIomCS/hcBQ8VwD/3TM4NTelt
BHRWhWGhLZ5LtijrSrLfgGzv0iiB0CYtbWPMvmUY6I4XqxPgNV/oKM+IIg3WVavohkRfvXPFjEVt
UxGPI2Vqx4fAhTO8fBQwdQKBShChDTBV/FDNvfiJgsTgbPesDg++L9pofKsEDggbplYXmcdPOkbm
tJBtFJpTbrHvHctwLHpU52BBxTztu2YnB88ak1dZRHO7rPn0JuMsEIJJPR9dBCVwSGeOOhHtW+k+
P+ATOyz7GB2o2JoslUixGnAQfQg4vEws1GraXzU2gJGPqSZ/Zk7ha4yqelTdR8U38IT/epXd8BwT
BAb6nYT9ORCkrZofsaEUdLzQwVqr1iYju3nkJioh6f85y/9izwP0oxrd4Qb5uUx0b/fTn44oHLwF
wYLw3gYA7kkd+gotncl5GptQdzX2AZC6OikWD750iBI0kXHO5lgDLFH+9cQvAcp4fJKvzQk+yFew
B/qqmrd6yKNgMM2AIvyyWUIzW2/deX3XFum2xr4pRqty5m4KeMq8LqLoCYoM1rkpiNaXUm7zZxbV
d9L6siakC6ytB1yL1/BaucVyJ+rDtH5yJGc5xs97hNWYMN1yB7W40+U7R5Eb5/UkgsSp3zS1vQ5Y
G8EKCP7MNFPwVBpmqLzFkSY7eBgkkTtqJeCuYdTtybTRyzsWE/rVyM/wxojIAXkkJPLGZXqNZxTF
u3RehMSUz4Af0zr+LxlFV9fhQItxb01dnvB4JGLH8BKDX36QKcIu6woIYP6L3kiWwTb7rx4Llyy+
j1yU6IpUfJFNGvHrcn2nQxb1+v4bQ8KzQ1IX3pRZ7LOHG/bkrw6m1caRAvv2f0hXdA/g8Zb7lajD
iT9KjJgXYLnBDspIASK/ZR4bXqL1rM8zYWdTHw3bKObayzFUjZqqDNCYbB0f6oVFmaXSnqL0Sd8I
+PtCBrxK3TJKpkDNVpx7LXcI9ubutAKQ5wqn7VcpnhKnp3WbhbyoJ3RLwoXcMYmyB2C8XDMJm12a
kuWJWjBiM+3Je3dxcOVvJQqRmua84SN1rz1+KzLxcI9TqgyBx1xlHTABvzpz9snbHdZxP1Ao9y3O
RA3AQuP8W+SdWnHiy3oah/wzizc0DyrX/O4TqXP811ppYvrh5QSPPCCcywEXmruI7V0/heElVQ2z
r0n+LVPBJTsZ8l7v1Si08Iy1TOl4Q4+sXO9xmp4ZpEIScaF2YYk153aKoDVhQu8h62pPT1MAV4LZ
pPUx+quiq+ckWNDQ9vUxzL8jH7BtnY+hGguAhDCtwinxmThRWmzzHfGV13UwSOrqlYVBnwrTOjrm
ujEXEjLwo2qpL2AEOCX+630gJqMVEJLyuTPxM4DAZeeRjpcc/UvYH/4bZuULXXwRW3fKIKGZxyYr
tb+jMohYnZJjKdiwpFRtjbcqgNrYlPTwW1v7UAQChTyhHeB39p/0ULCC+dX8YMmGimdccjQKZiia
GfpH8wEKjHYoRcuKw3p+OSAYOMI89RKBJv0v0gBEeK25Yaz8GK8pnmEdiMBXzDlIgXUtIGBxCFQ7
NApEAFVwdBJpQGaakWB5/rTW5YgRdHv+dezFhLfoqCBWaVE9mJ8RbHwSBFFW/qY3giZ9QnQv11aw
ELXp4utjyNK2moOuu1dXBz9YiqN4qmWLXdjBfoQdWWXxUZwoTmtZJc2PnDPQHQ+Tgr7sZVvRQN/f
Q2BmMEPowVk37aSZQC//IHNrYhKeIL2Jr8LWYLUS/CXcQbD4pBwRw/V3uQ4qTNC3xMfE3aV37rKU
1WDMKrCC4lvfEi0q+woyBRTGhJhCZWfgK9IpzqY8I60kMrZUMBcqy4tGkBtRPVwyhucDK/37GyF8
4BCdseQyRJX8q2dolYyVwxTUAgkiu9xnMpZr7qRZ0zAhuSKLDGl0LxpLhRWrAiGoz3fShMfCNZuh
tDzVVq0qiOwg/oKwaE4c6z6ttH/H/O42ae39m88uoST2BC8z/dOkcCOilNgov1qZ2C5yIBt0S7KP
XQMu/fCsQYeo3zXos5c0lbZ2OWL71Ds2xxFkVYBFB4/bXqNKVR78KyFdUYs0gzxDziFZo5+X8Cm3
D68aUgyiK/IU8Ya4oxL76TN7n1TBbxCvS5Iz/eG0Gl08OgV1CwZTxQBtZsulsB0HEnIUpwvVmI3Y
16n6XHy4rCzKYRVdBgr3z95nsCkFCAF4sG2xtpu5dA5NPVTawp7yZBjFdtmvo49Up4Qw2peuxM3U
b4YKO9g4HEZBy2yyjK9Y7bWHq143JVJvyiqXBmpgkp4sJ3mwyrWYNZWmFRK81Aw5a2uTjB/9HbVI
LuQhxegwfjoLItnbjouHap5sQH0ExJp2dfaAslavVexPaxCBM3JyRWFcVExo3Ytu0Ppvo+prxkXY
oJIBRhQ53j60PAeGZ/H2lBCy9UPjh+FCtJ42gJHPqoDb0/m7lXMOimQyJw6lS/tsoVOL11/U9kvW
wAvlZLSzQuwj/VL4SS6rgox5hItpIXID4MCOHt1d1lTg8QGueCKAKZJWrdoFyfmEP+lCwqiV1BK8
R2goRbU5YJg7m2ZdXGP7ijIYOuD7d6DKWLaQ3l37b4wHS6XkWhUyg+bhE60ir9u2zvwsI40TWMat
N1FJmHKeqH8Se2N+7Vn3gEKsIwDFik2LjYjEamIjwxdOvP4AgMcQ3mM3bjfVNrgRok/cCNTV47Ot
A/bpOKNooshCIjxkg+Ip6zli4H2eG4RIqSBTBiKaqm8LkS4XM0EAqnVcfUSuBQ2DATb6DyA+rzas
yz0xeVIsGFEHelREMq/6VnZjHxt80Wa5onXK/azBmdqmudZGy2OSHulnwNzKXIEMdeA/IdPqptZg
09zrb8jRe72vnqPgq5rK/asbKlyQ1FVdWd0ZthrVf61xRLOCRUa73BrmEOpvOKzJS1pmOjPWL8hu
JR8YRIKMPPjkjduIVA+V/n9vCJSdqgp3hWFVfTF6naW2I5GaTMq3EfX1AlGC0aeEY2rF55ILAVPs
o2N8u5T26ol7jsPIUR+WD7dbk5v7/HMXLc7NJfbxE/cU2l2tMGJ4ETD623NhbZG5H400XXBLqLKd
dQaKnqdV+6gLRTAMiVa2kPcpQb2RV6NRXFCe2M+LDLukCIDIcIcWmX6aM/394Lb702Jqs8sKAhlw
2m52xT4IO3Ngdr1H9oaFJW2L+JZ8Y/V6RnsIoKuo0B4Ze7BGlHPV/OkHbXNSf/zkUTTzgW81rw+k
Gxj3aECCGsCq8e2DjcvgO2RzqSPPpG+quxpvyX4jjGpEPt2yRwi8kI8mvrp+W+LTVL1w8YL+RMNg
tDPyNXT22uyJ8bAq/Iwcn0Mt7GSilx/4nw2RMGPlTZ43YQAEh7gnDXGdGYVRLhMPueGPYhMx/S5t
P8wTvs2lEdl0tW+VDWlU78VNqOnJE2OcPRsv5N7kHG2oTsNUL5WhrlvrjmQQOVebcPWrBASFvx1b
J3wYDWmgETfv8xAUfMcl3Wc+DCtQWd/QbKvsSZoeqUdtsyvM3uTGO+NT6belaR5OsrDf82F0OPwE
TZ6ie+UB8fGfMDJCtpakuEJaq4BtBgPhFnfehY05WSs+E+NXVrG4ZqDmL8aCAQ4SXYEoopOsEFnv
WSk6hRg29LC1LsybuG2Dy+l4mY/TuM1Ir2aa6aOGE5t00GHnxzZylWYme6XcUvVeKN5NtMUOiPcd
zUEXDM273cuuy2y9g1Ub5/SU623S2fS+bkFWcPUk+3RxFcOTrXtlkKy3e1Q1rElABS5GR0paatcA
25rG3GjNKg51jC9R7ZSZwHgFmOirTLv0OsMIO/4ShRYgGpDQ1+eRbDVNB24315+f2eKNpfKM1NTj
ZeKBZfX3xjnWZ69SXfag5Wg0Bag5G38s1Pfy0+BhZ38Gf8u7snRIg12/b8cLttffeFcub9cpUcYY
2WtEvPNZkZkvRSUMAF8R1vM1j6hV48Q5JwfQRCsv7o+dzPVMxQASHc15LzqxWXSfLIF/eHW+JaM5
EOczhLcbqYVf8QX7gjW3sA3XlUzRUWwpvQMhNih/RYLyac5QAM0/RkO348eFx8F9bdokzhovuALT
Y4nMGFZUpBxxWi5neVIYH+dA1xgWNhrRSiZzo5oanXxIe+VTmZnqoepUADlbGFKXxYIB+Z0o5c+4
F8mRysVl6Wf4DasPBYmplyWg5O8ZcD/Os6gkTbHLJGLyC18d0gzaTzdaGKYdeISVnNPuUXHuEQEm
1/rciLX9L2vnNLfiHWXhVLHk2W7zA03W6v4c9FDXTVx4nzIQ704K5gNar3s9vsVAmmbdzItG5Uvx
tf1YUiCTUfrD88KkEgrY/PCcdcEtHEvbNetpAgcnaFpqaG2x02u8bO2mFdSkO21lHIde6l7wKJaZ
zzNNszEwlfqrvkJFr3vfwYZvXJsvb7JvVrsH2HHbKQDivRyivUSwVoymmZKLkoFXo5TGiCCfvKCV
xfO2C3+KuF9d4EvX675olfl7gqUh4HjKtxPmezJdM/PR/cRZpqKkpG8XnmM96NjvKmnAFzLUXV3w
tM4MfD1Qv9g/AvO2IWmsVy5urNafPZr7vxan0fTi/IslZ6C9oKIh9xUG/jFxzFJc6qdRgk1w8DDL
tv2GI0oxAi2SP6ML2LOa/7pmF2FujSWTm1XJgL9FDmXYcn3x2J8oH+Uv3/rdnK79Ru+2hI7ziHrg
w7PIOZjDLJfhgHOtthvzG3BbugSuAMMzgYiTBOo7HpTerASrmEr4147BOzAaGXAZQCahJowSVrO7
XvEXmPQGpbP1+KQ+OVTocuoe2AnT+8VzBKxF00sYmnMwCzmnD+m5IDi/q0TzOQXXMFAVuouW4gbv
fD/V3jNoKeQzDPj5EMKJgrMVp02CdgjF2Ro2BZ7aWVJlSbXmShtp7qbHK85SW4I0XF8yIxx13aPZ
zJJXaBlo1Odi7OANqNruL+Nsf6HWPv/rVc1eyqX8/EHcj8yOru7nIJdI2vQ6e9DSkf/ntfoW2CTt
8CQgGz/iNpyi0l/LFG+0HPiZHe+G3NZlvavzjV/KHd3KQ3fiePHkPmFgHyIozKypTsrhtCgk4p11
aQlWb1DODlx3kUXkEcvNQjDFn8/UXZ6htR4kuw2RUKG9oG6q4mTfM/6hdABlprI6kEByNZcdKY8T
xvdw2i/1tULEsOd89nGQN52L4bCq17P4sth0MyOJyOqvamPJFl+vtpv4inln+yJHqk8SZVWrswxS
1jxmlakkJxgdfpTNVcIJgT6FEl7A+PoJu1WYyX1lDtpSUAML77k70xF0Cczq38heIFlWiD44IZrU
NlLXOLcn489EHvAmq0ITyLIAprhFZBNEF/NT1V/4xyrAp8zdqyQyR8M3QpwnQ+zTuz627nvE0JZF
HFhg+YVqyK3w/3lMGD822r8y34bq3dOAe9nkjgWYmiOU0Bg/Z41sgH5PW/ZMlRjP0hXcAoTUregW
Is7SR3T+R00Tfm3YyqWEhg5a23bZcv63EaFIYt4Ghn157XAg6WceJiYUi840r8750Vin1tUc9Hc9
ii3OPwMlKwDwAGxGrU8iyqqwY06VmYRHxxcDZr07yFdWrKB/B7mxe+n7tRAMgMemry+lQ8OzmcsQ
A7YIX3PMY6cfvjyez+msvbbBflCMxTXdlkcvbA11tHkJMtt2JPHTw717LKF/5IvsIz45EGCRxZSM
LlobMGOgJuXNjvxhaWodzogpgYW7ZT9tMg6ggdsm0hrZlnbSc9osroffeKll7IMu1hBGAKjJXdkz
xXPnukHvsfX3ZnrKoq7btpfzpcQK70PCbmImkkri5hmq4Xgu4p/XXmIw0sm6d+7ckUSIoZAof9vH
QT/tCh0Ed3yN0nS/hw1qEENyz5Qp06hN4BAsFppsVm49OouFiqS3D+DdB44iAhNQHsTE2fj2zkrA
3WfF7EuhpF66wTw2NarUAnEz//l8jev7iMjAMyUKWCh1ez+QINv8FbMhteo3f8OgYDoJskY5CmZR
HZifR82+plxB3SXV5ZKPKAMTMMUAM7ErWfhHUI9QGb4lMkWx74lMqG1aktnp2GhNG+PtN6bQhy/c
S3+nCiSBn+8QpritdOPAb4uZNwbULelmzkRbHKzBVGSD6Hk0c915djwGcZ2hy3ce8F3CqFPdj5T/
JFbBYDWGt5MYt/600PIxNQFsM9gUt1xhYmSsEfjadSnQWJrKLIFWrezuCcPbGsxwakaRBjho8Bws
Dob14ef9tM/Av3aygYvuCTrvwx3xUoetjZ6VqQA/j5G2+xXlZM/nDCugUjdpVjg5RrwlPgzgIsu/
H6pYozsU5Fks9XAokQIubIitFGjE9NgiwQrWwvWMx5z7XVTMaqIwTRtvyzIo3+CwsYNn4VYFOPXl
SwlnM0sRSllmwIyCS8SS19CCx03an83V3xwKlVY9PNlR3sa7farxaJ5ihz89ZbcnGnoilu11HnSY
63YlnAwwFv6QJtalfEp8sybs2SXyfisHaKVV0+VrJH1GXWvgl3uBdOfxrDdm8wFZoxkT7SX1R1TE
RCZGIA90XBK7z7SP4fA5PHP5jmkQOMwuQsZHF0TSW7mHBNTeK+tlG3XESpHrjj8Y9eL0CHH6MxHc
RmPiRaNJOPnNnGU9J2aOVBX1AhyWsMpjAokxuEfDpj9DTlJL7Om3nuRe69yK2eO9dNcZ18TFE4Fp
G+Cu3mX7UBkieDo7n71rAwHCWO5CnnEXK+x6KEIcGyYOR6kFqakdGcPuhYXsgEqsF38vdVkEGad9
tPZjRV9iL2BQVWogL4IlmiULMGXp5ZSaQwDyPmu2PzoqqqlaECErTVXGh9sSp1+I5ILP1gK324B4
OJSfx/7ctu6gbFlEwE+47GDPbycBGj7VAKmSkFPUtZnETRvGDl1Goth5i15TCT9TPDjqfp7bjq5S
SsDi09f+eDxhqg/pNzUuNxS+cfdb/qzVwxqb1l5VjCIZ/lbeKSyVsO6/5SsXdD34l/rB3fuENK5X
nEuwPfjn4evJIPc31pSbOq9u1YxcGcinCRxBXKQLGyWc6ViJwRTykFPHALI7IelbB04Dbk+++jEj
LHt1N6iBglWePHhqBZ9g3dH7FdHCDNfAs7XfIA3aXIE/M4DPRE/tUedyekDHpA01RdNVvBMfYDhC
tVimh0jZ7ok6axC5qozonfENVTrIHWcPFK+N0i8sn4X5ZhBUY0mQFtNdUH6YHf2izJ0Etj/H4w38
+5eZU8iMOASvpnsYu838VbP9P/pt5ipwrNa+ZCnmThisIqw9gruvKJd2aPO2NIwpVJI69ACXeO5n
iluBE/xmVTa9fsu/GU3B4oWxDLQZrZ92uym5TEYgUA5TTD9lN3cYrb4ActhT0KHRC8d6X0pQ7XJi
FmxBeu5pPBsVKF8pgDFsRVituy2gkyfn8+vpZHFiVH67GGansemhpqHn66lVBFnBEhC/OwG84E9P
N3gySXpMcFM9Y0JsME2ZA8sZWuIkZNyiWg09DCpH3kqt2ZpfaH9SSDhHPlC/fKv16Rn8U3gzRQ9q
QyaWwzkNN9LQu4sXdkuz6vzZzzPmwWYsRRrqc8ZkiCU+wrGPmifkNQp1oPUCZLRhiAnuL45xOGks
ZUU/XXHmlnjG1+t5rr4blm7RGHamcRrWjuKAv9WJuhQ1NzaBqXr42UgrK/aBrikCl9EpqGVAg1OZ
EtHVHaccnpDC2iTaL0bfk16z/OfglHWXGU4cMGNoqM/L+foUqITJMME903Ngi0ClgZTo61Otczj4
qHDQJgAxxcuAYM7of5rAFh0GN+o+DoMXSoq26dBWkIxkANK+8arwpfllSstAMEEwm0SvWfBcGX6j
ereId4J6u3JkNmpllwvTt5DAIX5RSbMigGvt4M9lFEDd/2uz6x5H1YDgY25NAXSmqNHrd9UdFFYJ
tPtsSnXqw3VEYMvc3sKatFejyiugh5yy73LqREboJag/c53cMXgdc/QlJ0aSln7tLtCAf9Q3K66H
52HTaPyF+1w/ARD7fh8e3mTX4yPQdQRNYph+DjJUB23eZhThvVQ9ffD/xUnuN4LwHCpN/sucdaoR
K0PjoGRu+2fB6fS4pyw6+z/WTtDqk55sH/rvXI8HFAt5YAM5I+bf2KeLKRESjXE8B8n7Z5biyuPS
cx/0JiEQbV7VhU9Hn5tWWDzv0M4TH91FXaguKXktHZfkfruyhciuGQMXT75WD9RhRz8DHhFaYkfr
TKzSXSgFP8Nb3574plQ/SNa8CvM9VxogOGJg2WqXbuE5tMsEzm18CPNlwPuamxdsIPNDE9X+XdBx
/CDrZj2etvGppaTKPCCFgNaWGqeAf2VB6zAtVQC6VZcE54H2dQqVzGinbi9EmHYfrxHRiojNGTD2
2A/aPs5zSIwf17yMeAYMeOTpgGZLet//7jaEDIS97NoKFqJdEAuriy1ohYcpVFs6+GZVuP/LwXzN
tSQD5jV8koC4M2Bf8YHkZCDGD3rukN0y5lJiwld3xaf4C7MQXuc2XHEXkWoRwxhpDlrbQPhPhsPJ
aD9QatLWl34HRikGU/VHm1VXTjyNkGZ70D3iZ84kypmmYMvY81qWfTPcrECaGvCo478/zLlkIJIU
3bmzQWeo4OllgdG8hKz2EQKZ9p+gjzau8/znTwBp8RTTWaFyG6p2STkcscg51fXhVOkZomf3Hsxb
tV7CVtZObSLybHSh/qx6jwX803BLqUWf46jJUtBQU1/mPvpaMuBp5iqS1XXSvpBtN9/ON+w38bdc
eHoeNsHCW8gaCpoo8mXeGklit0/SSyGqHApx2lu1ok5xhs7sU1wDcI5wtqXMZLlz7Mh9o/0f5pLN
gRz/5FMjq06boJ8IONc4RPLstDlu12hOk5M78hVhL4GlP1OPHlBDs2TUwFfI2YnozOSY856ADXWS
cIUcQI3owAIVHpJCFJA4UhriUDdIb3zfiqC7sftww461rJVZowVDIzQScWLE7V3yr6wcmGtbCeRV
R0bnziMPF1cyskGbMXf09qSDHp2/biDKB6lsh64TUK5gpA7kU5OghsyEDbrXkASVTGLeBluOza6T
DE84MwvU/e7GJqnp2SUcgjwZxAzP7k7Gg5kxxsgD8IuckyroIkaDIojux6jJ63bImOdoQ/Wx69Ct
+Dh+1lZtawQpHZq3J7g8JWaRrPdCHsfb/psj07TCd8DVYHvWj2t6IiA63XWiiOsrd3SLsH5/NslZ
v8JSgGcfyU7vRwY7V9qHValugMBqs2/AiIW28BBZoBJpPqBOYsIq6KUsU49pzpb+bzqmfpyNkMxr
a4vclGaf8Fbrj8HLluFQjdAqb/h/MJB9kpxLz5ji+nwuvIPJswcgH96nw/U4CqKN1XbCfFvwYYj1
VLEZ57RbOMQdppZZrDm3VhZJz0LxIyFRPOkR6062WQnxq2/67adxWWWsqdnHoksyfPve0+9Z6Ka0
t9q5vGkUoC8/EADPQC1JtjWJFy38q4xPplWi9TLP5Q/nK7PRzufBqHS3c/TSoiQskso/Twtc3YfU
xkvvUEUpioWzCUgzStVoa3v6wh0QXF2Z7a+/VtxBBbxWqDj+L9ZSIOF5IgPBJX7CD8Cmz8C8ZTMn
QQzVPGAVSeQ0791ZD7RSCxshOAHcKWTy3R0QY9HSV2ATKJ7fiwOAiOyi1noayrPMb7y2DstIPu8k
fQ1ADJIAlcc/+NQwHszBCnjvULKXhyHNBBRwMKN49Oc9PdNgmPRrMjWmO2RQvwDjQV9jGMdpNzmd
O7kuL72qtKZjvxXdO6YKxTprktLuY9fB1M3CZz11rKSfXifbOuaCCWoDnJMvM8LXeFG+iAPrNyvt
0i+AS4VR4yD6yMX00m42ijOdUzI4iWY0ubduwMbfFb6uhhy0D92mnuwv5mnbvxUfC3cE7LMxj+hk
Gz89MmZRt/+zvaMweWOt2qflaoWqTsApzCjzyen/sBQrEanp48aqzmShLBK1kVCLw3xtAWss+DzZ
E+GwGLP5hLttB3GkJNFg89na1780hOHqhJas3szL3w0ZWzIEXFrSdJaYZyik3LNbCRxLK1WIKcdk
mZGA7Pqp04ZWdl+hQSjo9FVpIwbakHVy/nXiAaX4DQlbtSVKqRCqWpdtvyeVqPTnngoWK4PATwYP
/Y/sn9UpxuGh6aZi26TLGLF66TIGRTlGaZ4I9DM4l5RmjDO3hOF/DKGxRFwitMpEVkgSVk6Ao/vw
ip0tt9yt9lAt+DLGhdsRzAm6iy3EN38uIRcCrhrMHLgSUkNWF/hNVxSbOJo5i68iAoR39oP1Zasi
JIhzWwMaQo8OybrFAbE7p02/kEhIUPIJPbcBz7UA1kKOcl00skoGUVm/Wg7baNIcHp6cO2v6Sfl+
6saDUPQjLmDqcAZDi3gPpx+LI5xclRRe3hxuCP44HfA0NAXTEA6ieu1qd5snBlSpwO/JY2Un4yWB
anTzTBJOW/BFLlL7zFIFJU+PqTl5M428Q0sU4I5ubjyLEJgi+AJGK0PJ9/pyuM3v+0DJETWCWs7c
HVweHXFiKYe6coEnfvddd6PbT4pt+ESbUzBafsEe4zgIxbKgVRq6b7p7CUZcYsCwDBz8pPSiPTRC
0/yM4R+C29tMTPPtCgufHY66sTQAW8/hGEITcZ7NHuYU9hVIzIdYonpteMM+Z6fDBQc+oRprShYc
Wmpb+fnkPaSEDZVz/m+c4tMrzzSkuj7opjnXaLPbAI5YDZ1BsM80NgrW7t+jDXGS5A6E28dwXTFU
pdELPvK8t+OkRh9HtP2TMLalyRQb8CwscOQTs+svvce2s4kZzTWq9MSszvtg880wICmUkpYAZZ/Y
8V6B9yJjjC2PlzEI9G/2YXH2hZgnVXcvquf6UAWHFcD1o6NyzHKNNzX59MNyQegeHN5Zd4Otwxoa
kDdrT85EBGWP4gc3IhH7M8zGtTSYV1jPPi6ZpBDzBPqqpilQ6GmzVOYtZMgF5ImpldRV2d60E97q
1FrGWZ12F3vghef22caLZXZ3kSWJQRJsYmrlIKQ4kSnRrLcxE3jyke7FOLTOtjgHhSRN+S2o7HWv
k/cQ2Mm8LBpg7i9Fz43z26rPsA0xpfixcT4ZkCvGUmDL1CN1LkmwTBYfJKiSRWgPiK9FQokG/maq
teP/Bsm7f00Mipy7RCzZx66cb+wkX8R9HFoafD3+7DXlFk9ECLkt8q6oizJ9BNGAuqS5DUUvVqv2
0b+XX0PaFQRn7VSLw92Jlxsh2jhrNCgAZfBRPJtVdskvVtNc8LVFFxqjzDaUofYSziaWxbBE1Oss
C1h++TnFQtj+tEGl9ylkUX9nn3L6zb3pSoXD+fsTW8kmE3ExjtONUVvzuMmnaIyARirDHsMygO0R
XDe3WsNyKGik6gxv2oGv24x4ygtEexcQ02TECR2yp6rFJW6w/wcv1jLksIwH2MUviYvn7/GB9QGy
KWSYmDl9Iz/WmyVmAdnDvkH+VFiCOOXLe1CMXM2PxiDEGLwRw/yWZsY9sbSjtmZwSojlkzS+cq0u
PiyoJQXI6vM1wzVn5fYwBzCJQrLZUCrA4u5O25pqcGP+j5MzX3Gmdr6wMJKnVflme2RHSifsd4Ye
IN3btT+NEx6Uwyp/D3AppCwsRMUe4BXabDvgdxXIDNsY7azeBLge9kd1eNEg
`protect end_protected

