

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
J8nZtW1Q/IGk5bZ13EIEEDntauAKqOlRji4Tz7aOFZMrRrl3qAAP4lw8839dxHbOPehATkI5mWRu
O3oQzXKv+Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PO3vY49rlamMYJ9pWAsIelQmo4roKT2hFecsbIIwc9Ce9j1Gil9MEDKbHqn/9XWL2CZb1+nggmfu
MhGokjjD0xhuA7bkrZ61EFG47AtPbrzrGJmyawEAJ1PNLVKIspuVYNxaD9rI6pyGoENRti8P0hyl
/TLRO8J/SzWO1wVCE+o=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lek8GlHbeyFgFk70bzers4fkqEzZWIlCFJLfSucq9OzFI+lvPoCv9lLJF6jbu+G/Gu5TV4ZuNXdu
mi0r5LAo17AD7VicMD+MhRKb3DE2N3pAEqyDrMS1jasKAHiVpH3eXVPN2AI+lDAVZoDhvjSuQjfy
us+5QMijcCxvAveyXwnL06kT9i9dtQ6hie8/MMqHXkiG7OYqxKm0Iia9+F6bzSI9YxeA8Doz1sM1
HWlzlbYLDBCHp8//PX7kMS2bPsw5C6UPaQ+TKox3agXXgpP4ea6EVU3GCBe7nIo37nZIVwI8YFKU
1lK2hwoX/DoWAQ9zzkBtnp8rOkj66EFG574xNw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H24CFb/lxJKnebrcZ74EB0cwdvz2M6JUcau88JBt2iuFL0aDDA6OprhhTeP6OvCciaaGRsBEok+U
cbANkg9G0zLP53/WvEkpdYtezlQI3mkakzT3UxyQr7e+pL5MFVi19R/4mD0m4WBOiVFQ4vPfnILO
XObce3WQbGcK+NGRsMw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RFnK9ETQkPWYtdMW+yKQ1MaijPhYXOMfuPVBKnsFVaRScaR6M3W3RRHlGeNOaiw0ukl3q+66K1rC
RHUWrifpwoSOSO54nuXmCv6joF0+cR+UF1LUkBtOigSpmJUx9SscdsvDcBNzrLmtogpoKRScYdGy
LrKeBNVoMEblduWARlt0XQCFRD4X03OLybCK5/hlbwAJA/OXY8QP1rB1MFXLkjS4zFm16T1j7dVB
psuynNAT4Rwsqrw26xpeXem+8Ft+gBzXVIL10rNKj0y4I07ITYInhk/p/CsNH9FgAhYM9jsWml7/
R3A8DckKe32XlGviTUqdr3zXyrsrjZFSJ1kTGQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 107936)
`protect data_block
K4vqjRW9vQw8/PCxbLd3pcenOl54ZvcDXcyBLEkytfva25GhkvdsSdHMGFuXX3zdzFcdQSU2CTtb
0nOkN4Yh2fPszv/p2v6seI9X4o3emh0KCYhClBNzSq5IGmbsK/f45mdv7kD2/pkuiQ3Z0DDVb99J
gdDZ6lfYI5myS4Y3x5mPH0z0hYWfeCh1LLlYHMaaCfD6xgK7zQz9lm1grQOoH7zj5ZPu/IoFBMUQ
ifrH9bxlUa/wTRfdH2YZkmc+oYk5f+Xw3Ter103iYE4wlO4POJmzwP/dUqs66TtzqkHcgI/dFJda
Yc+BI5golNOszcmLb017zq9sCpD5W6mHAIqtO7J8/8ZS5n1eZxw7eVB3/l5gQRLEySocoKs6sFQJ
BTH8Wdw++Q+ivC/QsWNFsJCbjBZr7kSuaFIntZKdAn/4VYkTCh91v2+f9s/zskNBY0IWkZst2yQl
7/yY1h+3GGK/GFlOo+Eu/1VWfEWC79V8Bk5TLAMgl1ea+UIuiVFTKJXBqfbqNv7fQ86sDk/1q7vi
iLL6mzyUQxN/7337AFSy5HObGsuJJZtYWhZusHZ6lCVnkRQUdB1XDqz1pJ7Z/bD2kU9jG1HUmmWl
7ayd5oW86HuZG6L0j79OVhvnjfwKU0U+weZ1JTrxDiD2sHmJGCxjgsoMvYv/AyfozPMXWTqcgQn4
fXsT9K0WVc4lx7r9iqJevJYOrBO1nWLWGuUm15kg3n0aSEgc2PxkvWIlaLTgK5XR5qgEs4kWPgZW
B8ESS5UoGBLOm/JSazKeYF0lFm51Pb03K7xbrSPE0yTXPrilVAXKYh/gNQucuJ3arHfzU/i6bFbl
AilT5LdRVcEjozRothEDApPWrm4l4KMM80jcX2ShpW0DPJ5+JH7oyfv4b8C4cZ6vJSnRj5pAkvfq
vR5IrwlauRt2ZvSLDlbsKTvX7UE8ZsZFkKedKW0HRd8odLT9Tn5gV2HvyTHVPUgrEDRQVmN7K7iM
lLliEB/vxlJnlo+gYR2Dl96JafFhefHGHadkpwA17kJWCp1gcnWgRHxcCuImcd5oGaPrVnvbleax
BYN2LjxuUkxWzXPBpO0vQPEr5kGvQLj1/WJcnyAUv3ZdeIjk2VlAAuV8dGoMswyvY7VFLvtVMLRY
4ucaNFvzgqLUIu6kEDVgTp31Hkt2KgBNB3A13SuKFo764TA49GaZcYcPq0ZPw7TI/jeGRSLr7yxt
wSdL9rhCOeWN4N3q1N6UJ6UKfeZoD+Gc+wXTOp1TtwvHybe1lBVqHx1oDDs7MYfz4yVsPR0RJEXW
Y1MiBXETMMa3fRjwqjipjgBVlZDdBz+MMb3kg9t6DSvNl48Te+kPiwUctCnT+5SynKpMhK38nTEn
tcrQqU5bdrhbhpkLmXC5V9Z68Fnz1Plo2Gm1XMjm1EdlFtaK2hPCMeQLZDWjJpExkCofn6g8bX1L
QcC0biqN5NeZoAithhNh80iJAJbVOxUFh8iNdd2bwa87hzVsgMxz0Wp1ioPWEWgrIou5bermdwdP
iy/k/FgKKj/qs3/BWteb7sEqKMGBj1NoH1XQsP4Fdgtf3lZ8qNiikWjE84rWOvhIXBdyh40PnbzE
vm5qR/vtTNUCmK6vH/zhAzrGkKQNBTSp2tZPFuvxmCZlVWL6IeMJuBValzrBgpRCyoyicBttkc48
0vVeE1G472tG5skyDgxc7HHwikQxhZQUUCxw53GwTTM/SQG3jCsOiXoSoHFXuaCowixaGPonqgWj
Cvl9nMK4l69kO04P3k2BPu1Z1W4I2KmujeyTB63NDyV88Xr2ufM2s2V/yZV6/P5jx8MqxbS16XFQ
RVkgy5xnL7CBPjjzX2tIFd3IUsfW6UojpOCQDGkuFHYwjcaHLhlLo8CG51VZzO2ZJaQoaM4Y1dVE
AutlhrGyEpW4NT/8zS3oKGtfzhNBl1cPsi+FsjbVECFrRh7M7F7OSfWN4mUQu9sZOrz+pCA3mjKx
IxL30d0MvX8nHKkdDGn/I5ACkfK+kbMeUC1D/skwqHPSSK0mO+L0hgn429EqU6XDo7HXtpet63um
eSh4IpxoEiJBxWu6b7KYaMvuTTF8c876qoSU8siCXSlSfIQXXAoWb69MKrh0T7DkqOE015pQSRDv
v55Ewo0rEsGk87hU1LnPyqSjNWhpGhFCz0R3ldOodKMiJ5KinvjTCbipwcqj0XtxyW5oDLlEVtpi
10l94dIOMmHI0tzeEKhEheI/arHwriUl813BHZjrhkAVrdWxcSjpBalFfk/tTXiRPbSAY/2irmsv
FarihjEDt2cKrlbD6e45qd2yul84jnplRH2Q3B09p3176Nbenp89PKLT7pNCRgxY4DRGqu/9xGw5
0m/70rOxc4ejtYV8iYR3fjtemHDb+qMVPPw+0ndIARX2B4QJRhP4PQcHwwIJlwdxurNNjo+tCWZW
U2n1nEZZ4WHsa/3tTgD4BBseUf+YYsXYEZ3WIyODWt0QN5vaWmH5viLnJ2e7vcz/PzS4Pn2ERzHh
0wre/rATAchrCYUvJhyT/yPzd4gxJYePimx1q8t7AW6vNTkIf1V20QR1OV6w8KlE0qbBaGa9xJL7
g9TMDWUfQmC31uE+Ug5CSik89hF7+C9ORSMMQy7hHBhtA+xU56X/xVIiWVuag0DNo1vWAMrjNPm2
8hrwsrlZI7uf5i6SvvY/u7j9cOs9OEl7dvUoozxk8zXEyJBwB6Tdwjj7VCpPDtiDSvlMNA3R5o0v
o+WpHP+Ju7FRQQuxk7i4VY77Bx9wr+CPXTsFlap5274N18O39r8+yCek+2vpP0jbSzX6yeEXBxZd
CMOv51i5LeifcFTjvrYeSxY7pnIlp2dwsxaMI0tJxSPBZazdyet5OlO0hvdGVoIo75Fre7rSw+cW
jaCjESUe52k2jxJhlvowee/RoL+T6+0tZVCpOOA0o0TAtcpgwnkgPAl5o6paeKoCubSvYINHWxeU
A/Xk4rsaNSdj/+jwRwc/F3y2iDy0m3M/QGrSZmkLd+ATIxJEkOVkSYug9PksjejdLwtPHLECAPuF
IV66l6FrU5cgbea4Dfw5SqZzHRtlmrS5cnBe1GCRwUEUkXD18ni9Chv1RURAXTEy6U7jhngIDLAt
IEIILSMkotggEA15d7PYpWx0Q0iCm5q9OFj/QaCMnQB2wtriXYKOtVUuP5joDQu/sBgDwBn6ZSTv
7e0oiZRfxZXQqZ2txUl0i7C6m9DKzWBrI1LqChhHMs/bjjGtModUIdjMhup4FiCOz9A4EQBbFPF0
g6ajxrcKAvaULJesHt5pdAfybNb2H50Doa+EK+hIRTkKUcqHYkhdJHZrDZPHfSsaurgNnbaWP11I
PN3K0skH/xn46oGB6yR/MJjVYMpDklZXA75T+OI3GUpkX9U0BlfVNwJr0INCpQjgk3alIFYAISSc
txnkoPqJ5fczcrIuZ6tHVi6rvnRNoantiojbVjN7vKnPcjdrYsZRX+xNHBjRLYJYy4wUjESaYpYQ
IicWfA0ns4gUSowNxZi92T5dmvdCaS2+cW2MdfRxdskula3zE+LYmXXtwHbv3FiI4n3GC0Tn2pWq
La+2WmcHWaNPa/V7AG17Do+vxRX59ogt/lIYfJnw+lEB4UIYVaDbMyJNj67nyt+UQ+yINzQHzNRI
nwUMXB6DWp0aLXjjlqTaPQm6ZYVKzIKdqulobvNHwzlYlSX1Omid7cHGiVSlXPWjLTSKaepkpQDR
0zPZjCb/vu7qtIMFQ6Ahb45W6EyNtmd57YLosWu1ZQKNyQv7Mw7DhK/sp6Yp6oiTx296xMsE2bkQ
QAzszDYc/65edPeH1X7CePAJCzi7V+26ArVKV4HAEhgdGKEoYs8qOZJlNV3qEHoX5NX7I9FvqYwQ
8ajNks2L8R22cD3tnHiXOgu6BKwUGdG1vt4JlguCdMk/ypNbRTNhcRLe2YoQU2fqmi8Zoali8W1i
0SjJA11nIB7KaaYb8TW2sk+qOsVrRymuzF3arKufewVCbowxl96e3CULKx5KL9v/mgkQgFhy8zPY
epJIMjOM4qracOx4S0volixK5nOQnqNB0jZKlk3Vri99Im6Iop97ZtLEnqpHJjr0ysUSoYc2QkT+
zZtA24qTJfFMJazGkfcgIHW3adPYZLIodE5xwpwLmSg1qDbN+4dh+SNhdpwnLB1iBQJG8Q3NF+tm
9VuQGE/o4za1E9zlarwIWVK0xoY431GokhwEnyswQJxTXDgbPVoP46cloY5Kag4UX0/2/AhYjjeV
LpIgPQrPOi1rNUN4h71VoiPSopIafuW0yffDqht53CEq84tp4zwGSpmXE/2NgUtoygbHWqaAcoAM
JEZKmLYV0d0i4EgHKyLMRjL+DjLmlF3W5OT44ClZlxSOsLZFSvta+Ek3Yj2l86upiZDBjMorixA5
pOnuWtVLshG5wRKOJfLzagZ1KV6Y2i+HTZ3MgrHpXClTs90bfQxwNwTpLCLnRJvmwBwuZs7c/U3q
S759NizwoUTKIqQyoCLFXSakfQJR4Z6l743i/Qol7UV9SEoBtak7CkWnkqaaxcUf7xwADVSlk36D
1pLjTRWRSHtr02oeZWkJODvR4B4hb93ENwNZmBUnk9KYVsREo3iviXspixvT4sRzKNkxD5iBqE3N
r2r7U3V+8ZMcObyL8nOxarRSYUfadn/xsCU3z3K69wgKdp+mZmvG7Z90cQEQ/CE1F4uYuvjbbXue
/3X5R1MO5UrZNP2XPzMntS62Wgd8E3XSuNlGSPqdHAN8CEGGjHpo2iHoV8XFPjTlZQZwSD+yQNei
MLN+MfRyWIsAuPiEMAuK32rYvfIlSugujh9tx21frgFiIoYu+WZkBlPVyJCzNtDwa+0OyQZJBaPg
0nPTTsPyLqI3bVtlGta+GFQgdgwkIXqV5kwRdCwuJFtEIkK7RZpokQScuxCXm+pS8oV3JXS+aRKI
XXbbzwF4tL4AvgEeUzIaFZrmgOtyq89P3H40wcFHl2yNVKO1NiHuVJfrx31DAolL177w32zf6sX3
PMJANtZUinodXd96VSDfTHWStsq8aUfVJXq2LGMbzC5yy5enknAEsmlhf/8jetZ0k4tv/gGvoROa
TJ5aG/P5se83mMzSLawlpVJvBxVXIVvCI7QVAqtKRqti7usBkJYDZFbepTAa3je/XHSxE7WEjeiQ
PiLsUpocrUDmmjmxuNFZA1Vt9mtjA3O9N4qU2rcSZxcth83rGVGqUPz6XNdjOWu5WgPxZWe/XFo1
UnHgZ2E3qf9c9m/8zdBlFTvM/Dz2YOlwuH0p6j1k9l5RttsP9coVfdBdbXcYzAsWCESDgr89EzWY
rAPXlCIMIKouzkPJ7cbXTHS8t6jAFCbZlaoOxOXR8IsAQoNdXx069MmeCeWl/LMZ/h1qlxPhpMOY
xkfoC776TT8gZiIQHgdzD7TbkgOuOP1XEKsbJRw6EtwM1goYaS3wHQgtHpGPTOuD9rHGKwZ2FAh8
YMjaX0Y1UlJMNW2HholLM9xV9p+JQydE/syc59lXnAhwp/Vk3EGkQaE2dp//+J2Eu3Ads2BNVNF5
pFTHUFvFABKyRUdEMa9UE+5ZKIXWPC6rb5GCPUQ53u4wQ/36oPt+aKdDRGkZkndW4toUstXHKLlS
vraR5ttb2RjxsoP2vAkUhX/EpzGVQ7yCN4dRbMWmQgS9HAChuiFh0k3vuc9RC7M7DV6OQGjuV9A4
JwpfCu4gDCOTqhqapp5t7QoJc/cQt0+Qn1Tn1LWyNxm3ry7v2amyLwOn7o51daxECOzfS3yGbwOh
37FBzHmSb97dhbCSEihOeyFJK4/NVKV0kBeBVuZBC5az0ncUrUnspWAuRNlyy79+VfTO8rIKc3b2
qJdaeqdC/1qjB8i24oiP3m37mCRX1DiGCj/jRathGmX0poF4akYJ7TMhvdiFd8bjuzmR2CqigVTy
vkHlwoyB9tEbRTazz0plJAf5jZ/ou5nD+jNfJRsAWQyzPALUe6EWAY+K+nsM+nCmTw5aWr3wptQV
XLJoTSZm0f8ZzxswM/RUnvG5Yx8TMeiV0GGV9GJzQjm14P9WPPu1abXc3m5I51rL9FkewS+SIC53
VFWlXqNyyS7rYdxb7r6oFinwHlZDjy2ck9tzwy+RW4LAR8j9/9S9lpRYb6Wfol3pps/PpHE28wKI
01zvLtuBhgnsxQfxOwc3yHROnYdEAAEX/IPL93ZEcatw2YjZqt+NTTtQ7wf5mTSigb4+oTH5zOlk
GaS3l0lHd2jvM4n+Z25tJZlX+4lppGo2m9UTy0/K+QIMlD2wzlWs7p77WM0D6CfPNjLJsFv4MQsF
3cpT4Bi9Qr0WZDPW0qX5m5VZGicQ6jQJ4VwpZIFLa1Y3nPvklOLqcPv2v6oriIRtW6sE77b9Hba3
/LJcTdE+ULgT3CbHUBSeC1Z4hXCVHT5PWurXvI6V+C6H9rKLYn7DIaVsZcv7tp1j7+TEOi11LZGq
7hP4fCRRFLeyyR7QXEhBERK9cNlb68rV7H6W/fETZh9VBgR681XoeOg5Y4ajHeYeL67aSZorIggI
YV5c8/o63A+ltSEDLxh0lBevYL4vJVzXF5CMwku7OWZd/UOxqCzHjrtLajSsmkc5JErRtsi7D0zn
p32O3Pe/7X8XzhuveFtiujhF/ceTtc3sWWrnnTem3s29X2/7UNdq6uMhVxBK0WX76R88wXEXT0zp
4ZuRJWqLytYioTM1wqCJ5c1W5B23eGEFhRUU9M4Tv1B6/IQbuX7ldJNZn1AgIZCNCHVlt2lYOx6d
ShzaxWQzj/4eiKC1Qltt3rjgCdsCWNaSvV0KFEYpNdHd3pxP3JNm2xHT0XoxsPuKD82x3RJzq7YA
2CRomt5JfJ2rwwZKEuiY+H5yYFiQdIdVH6J4xdXB3xJfOUxuiYvzOoA5EkCrvFMeKCMBYRhKl3L2
jjNktHA3DGpRrRIW8DlS+XXAu9M0ldavKikdY84BND47AAChtDrNwp4ToUvb6gOXd4qTDFBNedaH
SfdIPAocCY/W8/XhQTgN+lPRw41NUH8T0j5pqRWXhig6Q9WXGCn5+f/VLuT0Lo4K8Qna133Iu+6P
9auKB7EmIyC/pxc3HfASvZ0aIKGVsEYdsTZEyD1LmvYL39LwTPl8EZWaCHk6sz5bdhzqhL/SRK6K
GPOT6vNmjpNH6fPT9P9fpllZXUSSpn091+qJMBwHHCdfO++faeWBJJDRrAIn3hzda37U8Dtf5ZWn
uqaPGPebkburP7pEJwGbF0ndbsmvbv3A63I3THEq4oqtKV6bs4tqLqh+Svch03En7r0VMilzMitU
0Wj0Cv4wy3YgKZyvAYT3h1aJb7lc6XtdwOAx6LtypP2A7JApS1dGidqWiEcInyZlUBjPa5zvz0kn
Wi+7LhsH2+L+NqqmfQ+GsjWVmIGncy06GXHY4zBrY77fL4reIgrGbVVuWNtCAWuoXPJg/Xr/9KxM
EVJwZqMG6HL6NKyXPGbLBtfViKRsuwHVhJVccqofmbNQILZFj0BFuB/r0853Z6pBI+F6QovPkMBA
URLANdidej7PDPpQvfwmzWxRgPv3Q/KwFfntf/8lOwjdcQlQ8PcPrSbSeOG7egJCymQPhbIJXcB0
cJHxrPynAFQ3tshDHYW//IE+4oZQc4XEeWvaicXYHFQXHNg3IicUKh9JdRDFAxy7PC9QPqbNEC1C
9q9p3HcQYCnofA8kd6HfRvetZ6AGBm32tX1/13tdfVnMtC1YDCiqj65lwivq6WM/dJaI8v0Vxilw
R7U2mgtjQHEZfCr5MS18qxILQQOW2nP19fLChy0KFNuxRruduvL2g7bBRFQzj46idpN/gJSbU7kL
HgMUFMx/2Xyk0tV1r9IOMYEpR/SZl2JjXOq8q3jmHV6Pqsp5Cp6UORy9wkt23Y+RV+nSw1IeW6ys
sMy5UM4fQLHxZXKonhywwy7jCTQz52b4GNT9Vx7tu21R+yWxWVKELaqZ0vauImSttYCA+bPXX0JN
4ae7Fog9Og6fcVTTjzJAfnVHZqWrWwIPBvB66zVLZHblNDW/2nACFmJXT4/oVkKoMkXWVPhT0Yb3
NF4gcN4KMbFKxIwE+QBgl6Lx+3mW6IGQlaelIyAIJhIW1J5AyOnp6DPXBhcvOQU8gP0RF1/3wRS5
CZESG7YuApyOUld0AZYG73Asg1qJnncYExb6SrU3Da53Um+dB9G9s/Hnat7+m3vFkzWnVnSpG61I
u7N8dr4Rg23N/RD5wsBTiYTSq9l0SQftxwJe6GNG/Bt3dLE/T8tYRSupmUfiGnKLE0FO/GUtXnzt
IS7VHMFH9uR4xJqZrxgRBHHp/3hnfIHroqcHnmBSEPiTdq3Rd7+QeaIOPX6pH+wGu+oE2Rl9ozBF
kzGV5wpBMFQwZPruV/zhZY/Avk9d515UflSYaOH2b42ITXm0h3rLlUganyHl9jxJO5+B2QDJu3lC
lySkqjRDuMgntzDeF0RFFuJgIDJmmTU//ZQy7PG0nM4sVCnrRvK4loHuVraQ4YPMs0SlGObP8Tyj
xE7U47PT6YXOYBaWAIfeJA2qZoofKbY7t/rRDcA2SVIIzhKeVHcrHjet6VgTWyiDRMrfh4pHGlqm
5fY0cCfcI/nbOXb0upQteSXKBroRLMcmE78mrKSXgTB1lUhSi7iR8lTHQOJTa+SJ1k165GgoYer2
BPyCJgBMoVBEeQN4VMeX1p/CYfbqZk+6FGdJ7Ok/nTxhPqWBtmFYhp/UjiGbvpfzpzj7TB3bSJWX
eVj81a8D6M37+QZQgm1lYaWc1hLt2ux33iv/OLj6bWLI7Vb8+N5EoCOOtG7TcKXwOBxotjFj1T1E
pveYwF/xpk0wcYFPm854G3ZEYGbwzyrixQCw28nd37DdDh7kikBAPNi1GYrsbomtaYLrteIb936E
/ti9AXqHWLfi+TT6ADapU1LxuN3LrIzwj3ax5vhT7ovXw07tzkhrhoDHQHQDcbBMxazUG4vLqPWi
3MJUfAKyFpc3nFGztBNFiloA68vc7W1Mggt9l+68mbDjlDLIzL7Zfjm+u6omm3tFnbuZjiU1rti7
6YpaF6BgfQYKB0sBLXIi/EPSMQ5Lgt2R727p3Wj0ZgRJ0nlLvy4UNcBswcAxYYyzJC6uIDfqPm1b
mL6FKrN8lX/LDGxXmOF5QQGIov93VAtBYPvG4z9BaOfY9eujIbdfmf+7BTThOOcktefehCiCqGBk
4DyKwIOI+x1lrzfgfuaw0bm6ChuCTtIACEhZxFQyp+6wfEwdxd5x0jKonpiswLVpMvhJraFGXmzC
NBly9UuMG0wdhmXcR7mlC1i4EPSnR4wHf93iehbSvQ9qsO59/R8jkGKfFDB8CJpNIDfkcHAhVpbh
nJuwvqLhO4+WZ6eLNu59Pur6FdO9Xw9heoqzkquyYU4xrm4OGPN2KPjykmCVWkFEb2pj9HD4cnXc
ZV7gneOl1hl948xbVPySNo9L3jIOLCe/n3rFH9pATsGv81snyAK+AHP3ZT0GLG2eM0cr06QQ0kIW
Md4ZqAh80FpcqxwuoYQtpMNx7BUMYVKytLHiEz7CCqNlts5jXI7HSFiWkradYisQnlv+JouqaeOr
lQLgpFMTdtOOX8B0s1R6Io3KJAivNaPEV1itjOEz6xuc0eycVhlysvwBAvZTVj9ynvbuJLCHXzAp
YFBcYtYQPBQSZD1keONuSKKq+rQ0wcTbE7Y50Ird42/2l0oWOIMrAKdNlxHy/Ia6DAK8GiPYwrCl
MmLHbbGJTuAOOV9FCmUCSUWhgMyGbB+2uuuc66euhfRpQr2XFXurA20CK3O4qv1iV/Cob5kbBBVG
BKzldCR0Ef4UWP914brgNRyP7tPSyBepFSJ7fS1PClnHAWCPU0x2OulORGZX9hjH1A20HFJM3X65
L/h73nU7KHy5y0UnZ8Ks7IGAGlGBIb4MxMoeyaAiph0TXC+ktyOp+MFl6xX3rcV6ecg8TVyPv+7s
ikqHWkZ7Iiq/zrmioClMPA3IRnEc+eMm/1dC5lGd4w1Sx4sGLlnSa/5vKKmQ9xv9X2/Z46/OM62w
Kfk84WL34MApWP85zBAwSI4UohrU46tOEELaBqE0X7eAVp0yEVonIllAnuMtHdI4L5TOq0iWRIsH
CZDmaKkRyaAyAZlv7o0ZwaUWZ9wG/BJU0KBV0pMOzNgyrJKgl9J/f/AhWpZUgyYzOwT120KOeh5x
DRMfiTcPO6aRYuUslvBJaP5im7OGDGJ1vKoUpdkrhq64VkoS8t6e9Ou49oVis8ctEKAY5D0RQd25
U6pRzIcNCqr0FBK2vDLPT5mKixIpqFk3zZXH7O2Jjb8XrPlZfvZGNLGlDTmpUHNX9/gZ0fTi1es5
J/CPVQyKhzzb1JzVvAOwybjJ933RUBgN0IxN65skUm9qZ2U/1PoOi7l4/oHRjj2MLRg9wec3wtgu
jnQ/wg6lxBQX96ZjsrXmt0ZQgzxAys7TC3H7ayHWqnP+Ryhk41zjvzYgpiA1gDmGIhlLup9RoeVJ
fXFm2sP5RU2GvCFJ4ia/1XMXGLHhNKS5q9r5GrI4KQ2hh1JXqx+cQGC+mR05DeYzdNcrSCfj37TS
nPiq7+KoOMQhhYA7TudCCoLTcpeV/fDFtwI033BJDETwDn86vHTts7wPN1NB0irtwkxbDqFo19rT
2CGRb26KAcFuwKaSHPZykMADADmrey2oQsXHJcimMbNXwW9zeWAgXCGwvVCk6DLslscelc5xJ8V/
3pEKuSiOCqxEeNABI4Kj0QenP1OC5dIaN75oQ+2JjJhSXM9DvFVnB235e8CseXLbT8Z9YU1Playi
ntd+ISsRrtrB5gH23uwXbZwWJ3NsNzUXYClSPCNyLDat6g7WTKee1fn6c6OAA3Y8QVDrhZwr/NZI
yfH1HyLvkqS4qptQGkR7ZutZczPwkkTCt3GDTb3g+LV6nxf71nKJzT4bvlZlr1tgPOl8fJ5D+e3g
ztR1ycn5WWm7ak4KDoS5bL/fOdGczQMNJ5vTt2ukACD5I0fqd9baep18An3p6dIbtUBBhs+pOngu
NBdNnmpg5l3s72XU2XsRHtF0aVEeLXdyrE/NRw7Hiq33M1KXRZTqrQwLc/0yeLJW730CnC6pyaqQ
uxFt1RHR23CE38lSn2QTLCcdbsezBfihVvEuDaa6RSYycxeEoTFXb6pXvKnGEmQQljac91s+buqZ
U1sqacw2BpotBim9oCVG1sOF91X8qJo7WRkVNcUxB3J0CsLIlTJ3RDVsR36uhCAp66ofyWEPA4/A
io/QoCk0UMQVoHQ0EhV2U4evrC95GxA8RqeCeIRvphVs5HbGGaTu9Hq0rw9ChyGFZ2apVLF1wSLw
0n1sVqmhUgR4IoIMLPCiUVEdb1lB+EbIphQh4CYggoAn++sbngd6tw+O4ufbueXu+77sHFFs6SEW
xX/C7UKG5AvzFW6tdXH7BtkWwFujpCTRJKW9jiwoyXzOXhU7gW6FljKHA+ZTSer7cN3khwNzwEKW
IxVCYj46Jha9nuXBnKQnwGuVH9fnMNTXBf4Hk0maY22Tlk+vWx4fvkOajViJSZ/KdmS9T+Lhlbk/
sFO329tXgEcMcMGvaURlEd8RUK1KHS/6zWq6vyEYriNcX7Jix1XKXRbJpt8vke7LqxjQz/2zGsvz
/Fi9CxbmFnQnrUCrtn5mgevUihzV8GG2v8Wv9e4wunPtPzA8kQK2/zZOejxZYmm1DBhQpMIfooTk
1ugWZbcyobzuopdXn24/lz10tIEyzRylPfHTQrYGe/Htw+HffYcOrDHDf/PYWpF3TuwiPGi8dG05
W0gE/hjtEQZGIdKFuPUgoKXZancJfErakZ1M+9mNStcjrPySfN3oJgKcbT5eNTPy7VJ9siRiOdXL
84TSiFcQ7IQtKPlLoJG/jhUozIkbhGIjzFxjWS5llGsemakVmpM+rdNGy2pmkn7X2gbFhoVUs+7p
JaWUHp0bJCHqnoHFhFqZuCIMSDeWw8BD/rOpLNPn2CxftQmZ7KNrkSpPvaMTJrYQJ29ucOhOWT8s
RPBxZUD6bhYzuaI31etHanVxoOlUDwj+VXOpN4JFYMwQW0HeuCwsYEqh3ECUFyCN5q72Mu9t5qUx
nDNdKvTTd7laHnCr6qGHQbkOZwitNpM6s2u+2tHQAitwBFQclbkra9L21PGdoD6vysPzZgdPyFXR
Y1QLIyKMCl6fcEc6IeYu0WyWkkX9K/UPV6OALlp2xxw0m0PDRfLZgMtb+gOLtvzV6W5xFpiwQXW7
UsBeTFXJ8iQG2YdYcvjo3noCGA9T7YdzouA18o+NCUd+87/audXY/idVS1hcP20/hur6bNK0lrST
vMIWGXYHXK6CmAyLaWWZKgjo+cZtQWTxxWwgtt7H2ydd9SeaK5LSHBUW0GgTzAIhE956mTSDiJL7
pyf+QTHX08+9ztbTteyok1pgQkp59r07I4SHd1lqWhHDyMbCm6fLHxBhc1hprRRPakqoGRPmrA4N
445I6gZDaOuE8ArTxS+SpROvsWjKUA9wzkEQd0cX74cQuFVU7rYlgjJqySlDQGylQZMjqDfUlrrZ
6BXQePPnOXy9+5op4QFNyvK5CISv4cptLicH4f1E0ZGd97xqXNO2K3niAL2RPt/U+vavcZ+z6rvC
uGpSsO74NDOr/ZAzvQsWeoPAEFzZVu/LpGBqj4RrQX9JEg5xfzNuqen0aqv9peg4OuP29Q9OQtyH
8ziFhhGvzlVXWuQ8tY3CZfLC52I8ARcUmvhJsPVe6LNSF27PFQf5A4pP0duDC4H2NwvLXyIA02Wn
r7HzMcQTPn1u9v2E0D7WV0t+ZPpu1DXuOzlBZujNArpJ2k+KiFMG6GV1lwquE/SEDZ2ILmNQzg9m
/mh865GulLwb9Opkm1DUkudBKZBvhzeCskL3z2DcwvzD4ppCGqgg7br6b/6T8UmobC2mN1CIEIVL
DHVlYqnyJt5BAzGmc9GINpJCoKFY2S7ujYfy1PZc9gjXfdCCRFh2GgoJsT3ak7kXRoNqoKZ3ilgI
CW3Oq07K1VL/nU8NIAuhWzaGvPWuTTg8NmJF/fcRqprFQHaLPNJqQkR1SyNZ2s7siuwYi/bBzyXP
3mvtn3E/Lhs9WiqBFGbvlP0UNw1j2OQe8FqFUem4jcfHumDoZUr0SO70aJRgwg8rKbgvaIFuZcKm
uher4MfUnH/Gthtc/fheWhbs8g8l2b++oF5UYFQ0hS0qw+7HlkMP32m0udSWxTCkbq16cUJVf1bU
UUtuJ6OQzlQMcndG3vOGCyl5zHO4El0rgnywCs7gLGATJ+DRllrRdXSqoXxq52Y2l4/eaui6XbqN
RjK+cIvdeuQ5EE/wewx3o6KV6uAsTthflr8caaaHYapY1e6b1sxtLoLIQ1TJRjHICx/au6yNq2nU
1zjLFlulecTyYUFpgfj2eHKhod/VxakKhx6q/HQUThbfRTG6Or3iMkJXE4NOonwp/3lTU3W5ehwi
RVwO3ON6uzAhr8iGwDNYHM1Fd4HE/sf30mCV8ViDEbOuplOrMHz9AQnGNA9ZjOdDzy1t4eMjv5U8
oTyyWev6WzRAMh5dEzj9OAa0uG1p4N6e+4jwKSNzLYVyGqWoyKgc+4FFR9WG7nv3xOfUPXu4q9vt
XCgvAhRWk0CgbWXlICTNhi0RhO3nN3JNayzkvJkTmggX5Owu2Fdmb8/Z+2Of1DIEK714dbVQH9Cp
8nlXFo2YgDAWP6GHJP7NqZ5Lc4E85VsgaRsPbwSMDrj7VOFbdJzjAB6qKSHS9BoQ2BhQH6LDJaJk
TN3qhtNHnwsu7NRrZPFlF+HGY59ogUyhfUU/O0d0MwmPbP6NSMsCsaimw0AiUDeegjaYx+gajEB5
19Vt2eisJj40Le9BZZRUH1bIbiZo7h7eeRCJDof5wSqTMoAfj9eI2wo/lEiwiQRaZ7ztfhrCjZyg
sYZYUkSlhq29UWZaFCmMaO1KUJtrRTNnIGXmm9+4XRJm4rGHI3+AR8XDcKQIZobmBeE94+K7xViT
tRdODLuzxFJaVBlIuUcsBHa37dRPK/1wBp5FHTiEfxCvXspblpiY9r8bIQSRICWZ42h7Ajjwz+b1
GrFUo+lis1VzKuPhUcvZPDlHYFL+6YAEzVw6U/j/543T9y+QhjJ/skG7436cuOYKqmBTLcz12VsI
W/ucrnXZ9qKayFaFEnowcjdlyJ7o9wqSgfmEQbVghRHHAMgFOP8T++lZF6CaYzRrLnWK//hn4JuM
ijRZp+OleFKSMpyQV/Lf1P2K/1MPNvg9j0EeKfEr03r2tGLpLW70cs/DuEk0IDvb+GLXNGB6xQ0f
NVdV5N/hEWf5mPMaC8q+kbJB3fOVMkVkfz793T1RXhAR/g6eLsqhrPtTPOTf3p02fdldj9qZu/P8
SzAhIadPVfJAsFGf0XxmVu+mVXNNiaiWDi8uGZqnLmVmLER07hi5BqZmgUaeZ57vo+eCmUbgMajn
x82weoz9AYP4JyDCKQdixz/nmVoZGKmE3mJ0OxSXOdIBPtfbHjrSH4rRGNq7ey/6wDqjU2ApnYvX
5RSd/6KZU6j+RpVK7U1qYRHYQ3soC9hS+vdmWFDS28FDvWyJ9CppLlCfk/oYQ/t3Gu0zyj150p9H
1LXpU1DL1t6ciwmO29ZA7+vBgURujMawLnplJLkbfWa/GwTqgL0AhsfLJwPDOZbdw2oHwM7TFdCW
xzegXaBNopzwfN9T27FjcIkrgu15g9WBY0ikDP92KiMHoz7uuSCaaRJD3hfmwh5WQK+7NYicr83G
EpiU8uob5PJBA8XIKQTAr9akTVvP8uyNh4NkbT7rrvMoleSGqhggKBaK1q0Nvg9JAuYgc3G+mRHB
J2BU2xQJ6AzpoWRn24U9fcBO6aNdfBsnejNaMl4J8ik/19DMcwAjENYJ1+swHsg+vqnq+uYqHsRO
6QmkRbSY1756ndO6sHadfe4iSXQcfLC5S4s7B4LXdwyhnrp5HeGto/5pJPCo6gEBh5X7NdVMcoVg
vI1EYArLvmiAZJT3ZWhSmucWq97LC4nzkR1Z/A91jmJo5VVtnO7732ZGlmlghSMR2U29hlqDDwlq
WPYYXOLM7MTLS9+rSaxaAN/AfdpYE2M/hSI/wr8TA7PixnHNE8gVNt/4DIaRNwBzEXjg8t5nXiWW
9ae7+NsctOLiD1xhwHMihMpV/zZkLkMg4LdD75E7/YlNe1BRAOANL4p5C/j6JfSAIlZIGWRtoB+q
hFUA+dN9dyPukYUO8jnCAq26K5GlO5gZg0J2whqLNJC8ERND9mk6Fnu05B24gcFI1iqBhCatz0jz
STSKhJZGtwVJtUqbPLsPqNpfcO8vAppGLJGV5e/9IZgVKZLXEbWRgFi6Quj/LO0SHCCHbYBpospp
pdkpcS9313WHkenjjSTif+UUiQmq74wU+NiIv0L4fNvzbhFd7gXdD1nzEQUSLEyuRSqKOPFXSZdo
SkfiXVXPwldrpc33Iy6e0+UzsT9gPtp7z5DSUjUR3d0bS1qqam2G4hNSzgNvD/xAnj3gixr2JAKf
e1acj1VhOiwsezIfE9Vb/8XfHUoPEk3my2sGqlaDFYZxEaNiEbBAvOhDWqLR5pSVObIMG1z8Z71F
76sg9sM4uRwQJKiMDMVnCfM+GFtHkCxMHrO+LpKSjwxukAph4ff1WuoyO+8Y/NUP8yJcbYcUT5nb
sx3zTZb2AfPZbmpiiexZaEI+3OffK3e6uk5lyJzZx4RKja4/hUnvEE0MU3ZflhRQxjAwwV2KlL2n
aC8yyYqiDayT2BMaiif+TVrlwCgN1qD2wj3E9ztcHWBF1/DvhcseP0VIsCssv1EbhXTqBdjh31tk
r3vRqO+4II3zb1vRROa5nB8t3UGFDu6uBxgLGdL1pYdK2Z/BHSBjfi816uNdZaudCY2p6FMxMUBa
6FLAKYVs2W1KbdKDyRx0czy5biKVfirSz+1fxZMl5to5WU56Di18DuWvUQ3NKGDJIMOSKx5ZfstD
GjQRmGSME01M7uKShu4D/IRiYmXr/BQ2TFxb6zaaxygnhhQ5CnRuVObAG5IltKgoCER1mqRm3Q8U
DgRmiseIqbNLdlnuG8kx8I5BXJDbGhXcqZEIL+nv6A5Vv4s9RkhRvYZyruykIJbI4Cr+muxDT0Z+
SIvGL0no6rBOG5IuRN5B0DOgI+sZa1AxZWQCYkgw92EWuVNLKRqIIq1T42cTZFSJx8JCcpeNK2bb
umYLUMhTHIHJ9mrXgmvD9M87luDK4b9TwWqUwth5nxhujIoRPHZ/BoL3vT22J9ayCtVIZFeMhW3d
5RJB+K7Yl1cUTkbnPf9jDNm1CCCs4ixT59L3GqCzs0bxpnYK8eZRB1XmhNotu7MarLrvlr5Y4Tbu
74QXlTWt19UUgVMipC89tj2YV/WDXL8JskHOBDy+F7rzxvmFeAUGEuUsEjKLx3+BqR9NrQ1yltMX
9sBbwgH5F4c2NUtLs/1cIrcMVKpcHsj0sA14G5FwsWegugAQx27M1Kj8mNh2JnpR//tyA2xTT1uN
JTUGY5N7edGdYn93J57z5dHeyE3ghNwoWaeD7ZPuOsTZHd2/5h97hzGNHQNuaQsB0CszbMo09bIi
FMWr1kdyKFoidSmlMyZ23QpfBLTNR+2dOkjMOwrklAGW5CeoeGoJU+LILF+17n/MRLJD2X4nY4C6
8ZSWVMMqN7TWNaInJYWZIVI2RKuFbMQGnx4tOmLNrqISeJNncfN+wMfOTuwZqyd3I5USzxxqUC6p
cnU4/WCw2nOKOCP3ITxbDRoYy0BQ6qDJYFQbUYSuiJl7Q3Ih9Xa5R2tGd6134b+VJW9himV8r4zl
cYq9eGfax0pEiGa7aEckT6EGGW+suItfAKGNKQsmLUl9D3UyVIdYQOIHRiuAYFMHNKW2tMC/9Qg2
S9jK6SgTCv7GVbzXiByIBJBXEl6raSJW99yUpH/48XQ6sEFD2+Z5E/ck39dZ5KgWQ5K2bBA+v+WH
zZHHvUpGDEqRX4foNeaI8DGkNOYpGTl2XY3K+6RuvCTf40r0eX2e3l++IIvX3Sqh8kGs/K7vAfKW
w5NeQiUzDTEugFpAWMmYqQpxpXilLBqvulKwo1ysXxaS11x93qnsecuIpgun19ZL4sy5cmBmuGtw
wyBUiJCsizL9I7f/gI6ZUmLXnhY1HJxElGij9lOyPdF3AwrXVnFDS+V6rfUsiNgXCKRQ9/bBl9YC
Sdf8UW5xSDP+Qu1WOWkEVmzeyy6AXv9nhcqwAeImiEaSMZ4kmORjhhQ5J4/aD+stLCwXPRpqlAIx
zpZs4KRAiE+pWLDvxWNizu55cIN3hFhL+kYq5/prri2a/6hzCcVlLVFxq+O0OtnUZxuvCK5s53Td
Tu8B7Kxhd32NS2gT5LhK0v0Guf0P6s1VzskLQ6mfPdbGHwqTxOhSV9DmKo5JxPFqzud4nWR8N1/S
BrbQV6q/vPII2cjdqrbNQPYAq4xFAWTO+/86yC610eLNOQLb61UG03P7iRLYku+ru3XGDVHyz0NV
9r1GxPULsIefc58qUUZEM7V+PY3WH4ZysN8w4CGu85JRw1dcdOcevvkpcYw5EU4er+i+KK1Fmd91
lPathD8OEGUXyEgDzTMACNdQuDRFzPvjWcDS3G8czypvyX2g/Wkb32rXmYIDl4Fzf5ve14Tgp8v7
dci9TbyqWRk3QdqkHQGlaKlhCwMQL4945OTPniVKHS8eOZ/Md73KOaJf25nYq+vQp9WnMla6XEfh
z2s1qzVHEcLCTkFUBWN7VmdWrp3j1iJvIEKtkhggPm74jM0yTLSX0Vx3RmG6u3Wz8/qORJ94USPp
vlP7Pgtl2Kdhs8GDhcIpjssdMdlRwFXl+BIxUdryW61Fp6JXUkctbfjVl94pqY7eO2H5goeEZo9M
lu/n8K5ejI74j/OryhjBE9wji6VlnDxr867A3cORmXmaTwoUv8d3RKl2Vmo9TVWbmvNLtu1mXcok
qB9K4r5/+X0+FPv9j3XtNilJmaA25TgOn2cDW9buCrzqcffYJfWTqoGn8N4a1tk+KJtwZbkC/q+5
8PkVfO9MOYhoE7VXgL9NUBm7YaHuKwYvBydTCmzqIPJXo658j1EVvWTv17UOIrXM/ZksSJha76KT
vkE3w302/inkD7Y3Ek2uvn650eOShnMjDd/iinD/4bsR4StIE6hKd7aXyUnzcXJEHN4Z3jMgo4T9
7Tdr0VRZtZ4AOMyAJZwdn7TF2naRiKiSwA4bWTVciUHQCy2NU8jW6fJdwrd+gNHlPmdGL7wEf6oP
6d5cqZSOf1JnXRu6G0ujNnUqxQv4N61rh2jm8FmCphXPqH57kqWQruF+DhPlCBP9QQLJUXTosHxU
QQOP4mLxiFZJq+MyNEDVO79xh8jcCZ+vfE2+9TLjKF0VFXKZ1HbR5aRBF0aUQVx00HXIVeaLqLFO
xZ7FovxTHLC8zYXyfkCzsbE/XMP2xZQuzyN8cwJL5FOrAP18hikwd7hdYAt78QXxrI2c7YqHnHc9
5Br7RzQk6sHvWDf5FVyR9oqQiHTTCBwk62jp5S5QgXqzNv4HFa/RfHRQP50cPPiKdxL2b7AMLlNO
73JyO1QF1UmmNtujanmxLfM+g1x3NP4dYUveBd75SRU54xRSJol/eMg43Dyts4zDOq3zjO93EDe7
cNo9WzKuQdVHjzao+KN5cGdQuJ4l1F+0Y0S9XYQILC4vsrranyYm4TymPLSLsI4BmHTQFXCnZsDJ
SDUeh0xgirG1nQPF1OTkoejUE+uxPeOIcrcuSUWBF+lkEHYxthOLxpy7U9Ba/YvjKVQ5/anUeSe+
GqcX/6m5NWG5sv292UZVTMwap4Cv55+fBVb9nlVlqLMe9yKzfjryQUcS7sT0rSLRnWqTm9NUkvbM
9PB19CQ/kQrvZFPzoUZDjJ+NxAD47BniLFUAWNW6lMPQQOxe6AQ/sTJklze7fySG9sX2nJ8NN3F1
8qHQH2I2TU3QV276tgLYeVRluw8PxZU1YBLVSXFzXiR9mX4mQ1HsKAPOz65b5Oaznh0dB0FjGVsG
wlsk4EFm9X9SaB5LK/+rGBXet/j3QOhqzcJvKktwMm8QouRT946YikIr8DTTDahPMH7Jkp0Pda3h
T7nipqGlnW4U5nYuM7ev8CA1HOiX5T44X10unAHWirur2TJrM+KdV3d+n458Hn0S4n35pDWp1Up+
qnj/rXe+uk6lG8swJyCkKGzi0Dh4gZBLRkdWJS3k/2cucUq6Nrj44qYqEaD6JTvFzZxusjkLKDl4
feFWQLlOoRWdL0pPOd87E4y9MDqqQ84Nh79qtnnWu/8xtrpa1pietemE/abYBLSvRgBN3E1T69MG
Ip1DXIHg47+MK+gehietFEdhQ4GaPM5EaEMB2WiXWi2Dd6Rb4VymB11Om9mPSrxACcYCaPCR4cAo
NzkTdCPmiVOtcWU0JIZp0ER1jCwMG7tm8N5agcQ+w0yBNjt5DnnJVmhsM2JjUACq0D52z7uqqtmn
uxmEtSQibPUsiMGWP/1/JMPyXvDK4r9dfP+OXL7okhGHyci6n8u2gswq2PS1VxQINAsYS2MzcNeW
BlZdvX/kXSlrXco3kysrLpjMLvvb7SQqmztsbDom9fMftDrhJ5SIp9NToDHvhg0/iY5GeVCpRoGw
IpIXBQlhXc8rUi1bCWKq75enR9LuzGlIkvvKfNGXYuZz3ERuEv04utidcvXr5MR1DI8z9ISwsdyZ
Z3TknywiUeSx6lHr1IpZLRwwkd9WLR8Mg/aVNKdVpDzy6THvM4NEwNvgehfO+CLJxfRhb7QwzqfZ
oL5ZnglEzxr6ZMQLiCFhn8012PLIN3wXxwW1b8NY09vrm0V81h0UeV2fjq49zTRt0vSI1fQ4VmXx
KCoWHpfD1waJgNV1VZWQ5UtmKTGQnv4p/EnVd7vGYgdsQL3a9FqilGvIAsyirM0bPc0xbow2vTKo
lqWRNCSxHbtv4KmNu7L+f6p5q8tx7wm1ZiD7svxqmV4+/aboD8cI27BAtOX+WRkqtUw6b1h2AgNh
D6T6pQD43oTlj5rzJIMrFN6GTZdFoFns2htrE/H2n+wXHUtPwxjAB/fCZATXalSlNoOmHazWLAnG
i0TeUFqH6+kuFHrQD1i2Nza4oEXx5/vmIryXkJtwAO08TCOTaqmmM7rcKCCVAJEomu5GVI0uE+cD
6OMqYW75FEEyO3g3rC0BwNm8E20+/+HY2Sl2OJdpvVwqFeebTSSq16+OnFcz7VWsNKVn6CO4RROY
0HoPWxCb3rHmtLBd/nfM56KSe6ZVMU17Ve0p7VqLSPNIpocUiopbm37k1vYAylB2da9sYrWTV0/t
pBytKomCOXj1wdAMdn6NasWsiNCRsVxaNF2t373SBpMTltuOQxogtCh2liIwIZzXgo6e/LjkGEPI
cUsQLkLUU9Tu6LWl8Wd7Ct3rLME0wtmHrinDWHDd0+VvJKOhzrFqxcdyCKyPQK+cfQFoKyC4qYT/
ndDAewsGv/jYWVQXefWKG6t21eCOXIu88yEk0ggKMTG115lIJbBdI6fQHXyHMHOYDQ9YjObVIPAF
YuB8vLp2jhjNMIWTuqqX6Ws+/nkEDiTm/EPKyYylY2Mo7X/LDvI8v4BC6AXiOL8jFU9u3B6bwmPQ
BcbE2Dl/0gJlRYzS4gm41dSUT5Lq/OYjgntX7bHwWtnJtL/KGuN0YkdHzxz8C66BgzNrG+nlWdFl
uXLrFHuFfF98HlcddCpf2pjpwcte6heYOjEeMJIPiFMIpncEe06DQejLVuVjQBQo/4ZICVo32uf5
G6axhjRc51KnzDtyiq6RYGVAy062poDHl47a0uZ3B5P569ShJU5ziL0hdezcM2Wjk4pJctJm+EHO
yEKgC8q01UULivOVLzs0hwlBdlTm/cuii+T/mj1ykaDWtezNAhG+o3vrnnQ6nlDetuCTMuE6hQj8
Ut59IsNvCl4dBb62P0RUfyRaHuz7Lyc+slX1mQ08eIy9l5SvQDfReufj1YfEnvuD+h6AsWpsDLAB
XG2vnckBEvMDlj6T+s6mmW05BJDlCOkTrtNAl+QG+ze2ipfsFv3x8NV7XuF6EmuyqgycbtX+ld34
KG18Sc1b/BK6q0HnYQmgLxGaSRQQtTBcA+ifqpH7Gf3TnBeU7pxBMbi1RYxzQa9zVl8Mj3zsyXqq
WITPmD3ktTfEwq5a/HqPfsuxf1lT2Su5K+H2OQsPlzFO3fTBU6wiWfPUkf0ZOFj2s6RSMLe4RGd6
kZU72cdjsDFZ+OF89RBwHHNFQeFn4/CMIY75KyCdoeeBUIp/UFqesVUJX5ZHGdlMI0c00bFC6dMS
s6oJ7+8J7/xKAmyGHm8D/rXzk/EvKGtoH5kRk74QUDxpZ604BfHiFAeRJtU26Kwq+OQnren19OH2
hv+V9eS6UkpX3gJZuH052EIWieRtaXmTegM8puubFRTiJ8OfZyoW7iuEXCdyHRclLnwpw0uGR4R0
qsKXebP9XJ6Trwp0h7bzay7/xEHwqbgrKdKh7vfBV08NzaUkUafn7B41B2W3bCyEKqDBz+U4kF5q
JWCyxXXtZ3V+uZv0LdwkJlv9CFjp2zxMn/NKpyCnXtmsT0EZcjrHPxP1OoxrhAtOzfGq3/0zwCIy
qg+a/jpXjysWgwNyTai2o8d5mFWmhoGJIPPHh0AzdfAU1AGSIQfxTlZ6E3wnhG1HrIJDhkQNkhTL
hBvA2AHjlg5mOZ1qIo/SbkerNuHAM+mWbE4GKnrerrfhyA0XkoYzEzZ8TrU/ULDilCvcIheI18RX
uqTpawVQUbuAnwUkSJT85iZqJ1eqXwl9MGrni3UDIwj1f+1puKgwUhga3k5FGRpwLqQSdjXiaOuT
CjEJ9taaOglcImcG0OgmL9b4ggfZmidza3oZMUXOA+bXpyddiUha7sfxWvgElBaCwNUiIOruFok5
O6el/ERJbYI5lxdoSPuR58BMPobpAWW0+tUGGNyjhZqEbRsq4NKtkl+fimMW/hMyEFx5gDVMWGEQ
JX+6JsCTFwKPWoxEI8ySLnvMNLLA+BuHxFIdoRFTWaUUN+e2LVH0CcXIcmGZfm+wJWQ0V/JI7SNF
JRY09rM13H+rY9TVzULbH3dNNxkxx4Qa2O+7PwUQ+JzubNEuoU7sYWsNoHc73rcOsayA+OsUa/gD
+ruINpONW8cf0kxE+Xdp+Doar8di2Ai6C5Syx1KAD7eNm18f2rq1DP2B8Mjtob7Yd65/vm3syi5p
qwobllkoeYlWxEnpyZtDh9/GNbceUTWgc+OZYEQoAmjnNUCpIFa6Xot11NqEPsdgeDiYAGzwuLJS
ZA1ID+0VLTFD5qLnjX5JspBbfrpNvWjvjXYjL14HKhjHXZ/VAcH8oNSFoY+7lDO/w27gb6eQjU79
tvCu8Cf9Dx3921opeSi9jE5npJ6h1gFMm0d+9hLFrwdYGVWgb9GbJVMz1y3E7dnVqseiwfddSHfD
Fd5Nrp+op2pViat6TMPxIA8MoFvye1RSF1e86zvX1j4AxJqJ4znRdhXZ0xliV9IvJ/klD7znPp/k
GvCWlaEL1DSb4iuNaownTtnVFSdzRCMJUSSkyrrsNlLFPG8UpOB0jLxLqt3d9Sf0LL0YV2R/clRC
GfX1T6ZihlLyAtNoBkxt27SSy55nV5YWVxng3kSxjlApvN38EghdBjtOra+SFrrCuTrvkKYX2Whm
Eoxkdva6HLwajVI/bZ2acJnF5mVTzTITWuLStgOKPe47YlBvwIimUR8B1AqhaT9s0Hvn3+BhZfGF
7X6fH8ck76B4F2IiSDNekalOA92sZ+UVRGiROsh4YZXOTI0rJ8MVtwarbC0xCul/ctwy+P64xXEh
DcNGmqR0WT/Kei2K/1cmr+uHfLLyGTGWOqunDwmm2FRS8Vt0NG8eW6oSVnTQjCLR0Z0C6LMbO70B
Pl4qoyDgBtTPlqiO76Tm7T6f9aNHlC+TT9tOlkE+NjMWXGh/83pUrZ28X5CaAe4PXcSPiDkUEo+Y
omHYBBIXDxh0A7i3dGUaJUoh+hr5RH0ts+CvFtqefEAW6C53UslwsUkUuYx3Lg4Y+1dZPAtY0Mzd
c3w944ICn92jNSfCt2FiDDl0drj2USI5t1Txeg1BdeCiEXOO5aSv2X0TRjmym5k9QWRKpRrpCNtJ
37QDbx2OdW+YfQC/27nytj6Md0bixvUaC1NgqK6Ott7AI/aZZ74Yo77q5IXMWyAdCi1qzefuE/iE
CSZEOlfhwQ9yqoqDCfQIZ7SwcZWqXzC3rXrEtsJjaizFHiGPHxvWFJP2At1c1d3Sjt41QfzH/ZPJ
omfwN19pdqWcuLuLLwTYkzErK3O8bY5wqYO0OiD8lFAyGbUDqiSgcvwWf3QR8vHDu/cRjD7keBYL
02G0lshIQ84F2Vk3Bk9KsRAlcrmj7Ra3luG51bYPqJrCrPZlWf8ZN/DG/7zxOCKmpbHJxrZau7fx
6fpRTmKQa6e4Ew7SDJX/1Vlt/PbjAOtmg9bfdMlVajowWdRhv7kb2He07S6m6vAe0THRUS34i7WN
NJpQOFV/jV9lEpRkj2sBhK0xSlHTdz5//G7FgEQHbCMgIsUsduRnUaInx/q8MTsxIUtsu0b2llvj
HNPXMaPiXIO2JBjrvxDSU1zRGU38ZlA2pI0cZCtXR9tUaD6C3JvYd1GALfGekOIRZFrcbBTuKo5e
pSiikKrd15jFzoKY066bC+S1Q6scK6ISmfcEsNidmaCqEOolq4BZTMrUUoFBVZWcK1w9WLzw8bON
NPJmcOUKkQcnlHN/61dNaJH4F3ugFHoMZxDCnOV4YFahvZHkdF+F3JNKEGH4wigGH/Y3YhBZJSgW
MhMPiH6wD3ENTjWofi/OFSw2zpkqQ2wZ6cJOAbesgLHW2Xj6bXYmfo5rwCxOMHF7krzhe15NYAEP
dJv4Jolgh6ArObiw03XWpYzej7ItU+ZrnbYnh5T4T4VNVr77hfrwC/6vdkOoCh02XfZiwTG5gXQG
YcNiEiXMZoyVzGVIgGpswlzJyGZkTcX+awoTVKGuvWKZFxZOn5/gi5cEbTFw8godLGChQd7tCmDu
20MAMLtfHM0xGMBYLpOELFXw47A2O46UEimkFjX0EtvcjHXUStRJbRJxsLqqlRhTPxMH/WZL6QJ7
9+5h9yG490RIszZXWHkDwoU+GhETfOJjmQAeT/mCXzSyyr5VdV26ghlZeYFHCVQLPFx6AnUpITaW
dLZ0B9OtGAdiPIyxlUNvAlyiboQosCBZUIq+mBsirJ3tHyHSmVmwQXJ60G4RkROMdOzsnYENXw15
SoND4SG5JHpi7sUiQcK9ToEBOm1oW5apdMK9g2bw+jbFpvA0+Z+F5d8OICmuCh+yjjwhGaoBc3Ef
2ERNwhTDbWu0yvnGzOz7uBxWAZZ4w5XyigoryVUV8XKRlb1wBpKIj4uYD4C438Unsmu1fAFhxGMu
8EvIPcoBHkuSAvnitD+sClKdKNWhbY9+0HewVGLFJUAdpgMELkbUfw0wWZ928erwvmNkl+2JYPYW
1o0cHNDSgu1ubWOaXOf0+zo1ubWgYLHZnCUaEE0VWj0JWPU/Tl6OVHiIaI4wYg3ry76RnVeBp3ey
J80L8tsSCOo942HHynDMPv4jfB0PObXxX48dO/ojAwxZzyVg0F9H4qRPlMiChPJbyyySs/j/S/J9
t6kOMd+r+dhANIc6EA7shwG1Nu7UmnWb6rlgDbV2QWjjAdEEOsnyUaJ8tz48ec3TPeBAwCdZxTi+
MyRocPBv6t2rFyqsZhcU9ImLTXxCrCWVw8bBZ8UtbMWfhkvDAPW5vUsVQ+KTHlmTSTk64n6r8ZRZ
55uV9I25StC1nlnPIGiyGKvB3+dIT059cbOXsBO7m/K5ztCysM2Wa6/ttL8nnLPXxVrHoa+wk9Yj
BJpgq1eY4zbmpSsSo9UvHTfr5PkG2Q2IbzSkJKpB2bnbXl10pF58fL1fTbajPeu5e9mAs3iNjPWU
MGm/FzwLe89e5yD3I2ep5g2jrcSaLWWXuWEd8sIXdou1CXR3k1QvaxtkJyKQ4s6HrPpZvLPEg+yO
tEZvtwVCMKdi+VCBLnUIqsbCDcv0QjQjUpL3ApCKyYssamZMCCPHDGC8WN3tKrWJ8UINWkqxHvzq
259NULYsRmLYC68ap7WqSYdgC47tVWzRJZLpoSVMU2avQzQKrxf+VshHVCvIsuCw31ga+m8wTsHA
2QOmPzCpVOswJb398ZOHCZN7oMH95aSHjvP4ky4CScq33NL/ius6Re7pMOL2XgWPbp9gSoU9Ekic
WlKYC0W5fVbTNJpWIRZHrHGZuOGp4tb0Ftt221QUKvNTxMcZFzJ2BzsD4hgHP9HSxFsxLo9TzTXs
Q/o5P8rT/1uRcjdRh+VemR4sJVNq7hKC56KzUTsCBrKyVqJ276ph+P3QaNaKDsXp03uJDeMPdTF4
yx/KUjQLPrxTDuNH1ZL6D9OoC3JE05rKqsXAU5s2KbUsmwmhuIAfarx0LCS7dGkFqbcvgnlim9wj
n/XfcH4oN33rXxHuzfOO9C8E5Kyf61bVAAmFvCEW2X26Fdukvdycv0KzZDXIOe1UyerMMY0XJcjg
RlOyir6NzmDbVVNLGOqsBPpuEXpTyLVSHYvMMyCzv516mZHVjBkrtmlwtyFh0fpVhGiOSX8B51Cw
OI5e5EmkP5dTFk0z3nRhDSt7Yf323Y7OTNGHAJ8USSVjOKBUXACzaEZivA2+iwvNSXL4+6Pdr/gr
Krb3gp9satsG37cGpQA4b/TebAfOshVk6GXxof/rknXw67WgFVNLm+g+M5bphhl0K61LI5Ps5F7P
xUEslNl57TPE8AtrnScz6AEQJHewIAWqMj59xXNXejimvM++QgvfyfKVnM6SWGkBzAORjVwhG0Li
Np1ZMkCBbwAp0yKLXJ7HXr0Uc/Ch7PmxDeIQ7Zu4FhDhqYYHzyQ9ZdPnc4ivfi0a3g/O1fHnQsss
5sMNclrMwIFhhIpPtNwfxbmNCisVbx+D9nSioQ3D1qkGqhXM+4k2dlJ9CUUWK0sfQv7bEZnLTzdc
ARDlr9MBQon4nbNqJ1r2FySZa1A8CffXi2GeCL+sd/oEDM5V3WOC5kS199dpNFkxJbXRtNnqf5MK
HbWZNQQOO/eVWbke5RhU6MhmrFG/awbAR1TrYgvnsMONqwelgQKkTelzPAUE+IoCOpaG5lVDCtEU
0mcp9JhU171S+oKokPPgS8rFDCf+cN1hhgKxMGnayDKh/Woy7UFI6qsS/KAfmCrjbJ60qmQfyx7B
sP35tLNnKgDpMRBsPDUMYv6DsEk41ohm7bhkxP613GrjFLL1XagQzk5HNMbpFPPfLfIcJz5BYUQQ
b89CBi/Fd+NGmyJXyRbWrFEhANJZG1qHBYAZVbB+miumITM5paE+ScsraVPruT0nPJ4hxOqOjayk
iNPdBGQIJICnaC/7XzEz82PA0FrDggv1TuGvS63DGDyjW4PiHpA5BVRhEKK9CMYGdf3DykZ4FG3G
ViO+TKNrS3EFBhI6T1TjSa76zXeHnRPzTgc8bni75b99nHVNu7M8nD0g/vdqScnZ5v5YjcVDBkG/
NjNSanMU3GNqE1GAXKCTzo5aH9rzWl8ZEo5uMqJEamEQQ1fJNyxGz9JbvcxiNnEaupFFBmje/zLe
RB+3qkuxhWxOPBYbXQHqmrS0hn18q9ugnFdw3EP2FNLp6YcqSsCw4qLoEAz1IFWnCVcUYeVvwHfL
dF1W2nDSX0aKyitAWbZyrJy40CkS9CmRvsbTdUwdLHJ/xAeQXQnHhPdsuVs15nM30M6SOZw3JwIr
GdjOT++2hNA0DOJ/V3t3osV4R/kK6SU9fsb2tRMX86MeGLrYK0sy2Fuvp5q1iShyOUPp1HBDT7sd
t6zArRlFju8vbPPcvUeBTksrzdgT1zXalnJY0dzf6UHkfU8yo2a8gE+0N16VFSV+b1n4ntIl6w0R
KMzHT2KsReAW2iwhLZ9xythb5GYRlIJZIINeMFKBW5bYfrMhDT8NmyLFmp+HuvaGoQPvzwjin7pm
DSVBhzp0WJEyh0SqRdB10QwZl53ep0tKJcSAhOdwdUPT3uT8s9AqU7lOaeAlARKa4WPIq5MUotrE
F8iAi/SPMPJJoIc6faGTbsC+F8zP4/l3swcLt29nKUjPo6BXajyZGGQ1ZNy9apiPJrVgRF/TVdVS
BR7t+grUuSD/wN8I7NFW+iBAH6LGz8uSlVoH+sPweLPW9P1p3itPm3e36AAc5atXHyotzk1HtQsT
8gSJCwa54BrJNX6iLLFMZQgiHPubfI53NpUtGXlJzEJmL5mt0C2ykIxnyG9vSL4XhEhfozeZLZXu
By/PnTK79Vnv2NiLPFqoygmoOW/aGSHrtLpmEhkdNPynd9XJa2IxZncnUE9GatsbRHSKlXi7TOo2
5XWjsTe2l4DBaeOpebyR7g/7/3bVYsqAE6EeK8qyQf32mclaGrHGPBw6MEjRL4IZRANTvyzkCDA2
x9h7EEPBa/Cx7q7ekglwGjLN02W0PCNyoDEnu6HsxWinpVOsJmAuNfmggQNBckU0biRu4NRjll5y
Kemf01fNPJdqlhv60xey/spY3fjQLJQc+D4+jzZwbBLEz8t9r4i21C9ZZjE5f7heJbOsbm+aaX2E
ex56qQ5tidkeVlZspR7hcY14bABpUI9qRm55qvsBPqNrBzthjfS2racbVz/1aMeNr9pBSsFLBxp1
76zNCzR1ueE0OPXzbNd/eAiG/GUlCXDnYrqdXiYrEXAgFNvxsOsSg6MtIBHc0Bj2QChC15v06Q52
1VtJjEkIHx2JmTh2YSSSE730CP5ZPrLNRIw+ENi3CjOiRuM1sUhLzf24SFnfj4hYJY/S6gj/F8jO
non5PF82pSrDDwtIWPkK75osZ2OlQ5RuZI8DRytfnUDq/YOYKvWwuNnOfG4Hs5YE2MZEho+54j3G
ns5Z/W0iXF2lihmGH/RUgPKpB5tw7fetgcp/FVdyT4KZfpsk3FsmewOUp1kl5kgYHrR8m9+tqRgP
uarjTNW+vI9dQ2XlX8tSHA2+1hbIpZ/YRU4k6KX4bEiyGJlVEGmI9cBn1gt3P33za61OViXOLqaL
Bj0yxu/1jA/cOVS9Oc7Bny3RQZqen6AXtvUTQOiBEUb5gDgTuUJzkPxU8L5KUAi6gmPr89xIehzN
6RDCOHybci6Dn5p+FXtTL+x3iQNBSocpA7Eu2eGiYIO+cyuCtXTpPUGcUxo6IUB2fYc42TiXB7yo
9GwrxHytQJNJgStazoch+iZGJPfx/7D+228Xu+qpNgYVMuJsA7LtMiM9wcwHeJFRatAq5tQwxtIN
CtIj6YACQg8uplQ42FWQpzXBP6mgRqrMXSFI7DJCuTB168C/ROXOrqJ54ZsddsKUDFS8g0HHwk3p
uZl6l5DKkfy4/h+FlaIynofgZIQeREXgPTBDpzxY3KX8oESAbPwKG+CiEJ4jq1lLAvlPlAu53i5h
ZkbUz3lUK28OLvuFL8OqLdxgAwMnedinv6lyls/gHV/LBwwnB8lpcTXVZ/deFTNeOF4VkGlv5BPQ
L6QbdCvS/sT6+n911XT217liYJRbg481VMP0SmlYwSYjU2B8IuAr4/GcXrpepEYMkutMdvLm6ANd
oxdrDoF/w7tIEt7DlCJSfPP4DH8Ekdf4dUu/nrGtX+l5sNqViDJEqpc4AEmszBy9Si/OPg33lSql
tz2HB7Alv1tEDwyomkecJrl34KTsShpsb/T5ZH+qbMK8VMroQU47v/fGqxP2gK1pGPeM6IABwdiT
aTE+ChV+J4xl4RfojoZ2OtuhvPyHwAx/uJJRczC8kmF6tC87Bq4BdxILO4qJ7L/040JdxUeL/NOz
LJ1DaETrTHd3fzB6CsEqMtC757zHw+vqHMIzenG+M1j0UmswpN2Pyv6JBS21j/2M6k+Vm/W9Tgvi
CaP1Hvo648uYSO+nnT51lswFiQDbyJ0ctvkusIJdLwPu8FjqqbxUsVGSzUrUJbvERMni/xIVtnSv
Oyptw93NAAAKuO86mJ+9oSI0dek3FbZgkVbeHAPpPnCoVQBCcuWt9EIr9Z/pWMNdQ3sr1kxNyWZo
fP8jHvu5tvGPBpj/mOpjkSMvQYK2oTobHuHB9nYobVUeBxlWQmbKsXGEYz1g0l85OWOP/fKYS3TZ
Lp1svzYHspmezxJ0qjtpl27uOU985zpynJ/O+JstauzBEW47MVOeqsEOHCF6EmVcq9pavg3htpmm
t65AptNjUjzExbk+50ADigGTjEEM0rukHfm3nSbhZAkWu1qum5QtzlhWDREJZSCHI/c3mB9Fjo1S
CXVcwQtHfb7/IutiO6RvezGFcuHTWF61Rk9iw7W0pSF0RGNSRnrhtv6jHJFPAsxwUMyfapCrfvcQ
d8+LI3oiTB62nnl4NCtOY9Zd7UOWtpw1doIgBIvEFz4xDRXrcJvu0sKC5YjxUcoLEop2SaznTuVG
Bi/7mo2fS6ks11vzsOBD1UUjoEf/GAmpd+Asf2cTGot1vGodjL0cblAxRFrNAF35NAZFleVUoUAb
1am1q4Y+Zqckqt+y3LkDDClEBzw5w8AAiII7rZTVAdeL+64ubhDuXPDT+kc6XmXEkEIT38FdaWCC
dNyEEElAAp301Wmto2xR62HwTMdS6iNmb41bb7unWsEerFnyTy6HLfPMmlhfBs5rtOvkZDw1kJqW
qsewbgyyvynk+KddXjle06cesnYSgQDDHyGm2x9lemILAqUW+yXgxMeFwS6ke/lULWBefo5d3G15
bYfpp35fx8+kBUKaf9koiobEdNwY966T3043De9HMSpvhv2JDGrS7cXbm3GbJItXdHbhrEpR7nQZ
fLGCC4D5QL1zFNP1xZ+OTtgB4WCos4cQKd40qsLUxWiop8taQcE/WaJL1H7OvwyzlDBdBTiI/+lb
AnGFnc4ThTS5JZMlkngGLJ63ue5b8H6mi8LzUcYxnT1Gxv+NGupsC7ZRmyct4pvpBzIBhQmzgXbP
lY9/hVm4Wl4Bykw2rDOrfXqiM8NrbRmqcMoD/PjIeRv4XbVH4r0oBgVXt9KI8VYkqxRZBsgnitml
mTOWtZmRAuZxquQH7qOWiVg0h/PpcVYmlhaRHxoSGbNviYqo7UtQ2RdjqS9SxrPKOacrHfaFNTG/
TPDakfAaaGl7BTcRm6gFv/B2fVj7b6qV4Eh6nk5Pm54K92a3wS8UxVCsgzxPZDXJgfJmDiKmZ0HE
AtHVOuU6F4ESFpO9+1ivx/GwM7VrVS337A3XMVVMc0e8h4OzzxTCH5nt5GF/b0b7GSaisUDH5qd6
bRDlKgBph+wZDuS76b+RS83OS7iHFo4WtbXFVpIUB5iT9OOxqcH8MQzuvFnGQJ0hG+9SWtxY97UR
uhR72D6KHgou4OFSlYjCbxq0Arrv3J88zLtfC8yIlD4whpgCmVb0tym/see/EiNnW8ETEJLNw0RE
1RVP3B9ooEPpop9bS+/Io74n6GOGjPTvjsAiSyjLtGeZV5XnHrm92iotehUsJ4CnhtyrUENdAoZX
AqQVmWmUUORr6gOm3rC4DIZgccbBOCB0XVXDnwuehl6cbpQWZrJqacUj17x5lG0eyx0yZjjIe0Om
lM7iQH1JZtkTbYX2JA7PU4TP1S/7H4K7yqy0b0asRtwLaxWqmowrzCPFQq+MWb938/VnrHKbokQa
5LRJt3AimW+AKnZ9nwXb48vfSaSgqIm9nkD+Q9F5dYUVMpeEelchyU7CoKxLb7PDy3zDK/eJ0d3x
n3gzjexjcRu3eWyVSIDY8M3Gc8YCSOvOYdNvM8BhiJzQNkUxfFaapos86sy3noBpokXKcK0CirPF
3COZDDqVmAdd2h8/loCtETxguhHJaM/67M/wOGtpTEOgqpiXjbycs5fjdEcqtRqAWkAD0CMnjEgz
WpSb9/lQPXqfi3xyZ1VLE3cVfeaIoCvz/tmfbI146QDjRYcsC3d4FbqCHR3DFA+cdqujqAgMdDSm
O28Y7oPywizrGK/jJ2Oxkgu1wfoKLGcQfIuL01xktgylN15B5jZXS1QVSmRZh2wRQRNMbyb5PyWS
OzCf8t04l15tT8kIf4inPPBQccRlQmj8aB9G6EoICAZlOzMShMuSU1DdI+aj0G46SzLWm6zPwPr8
ClRd/Ix1oUn8Xaasrnwc6LvMaHLKKJn4oe5USeoSWv9yZ9jhmTQ73iV7YI2NE0GhgPvnE2kheVoe
aanjnx2m4lZR7nINj2mdhGGdnmUVzHj81c0tbkVyFjXUwOZyAL6P3ZSl93zp9MU9Tc9zf5wi/9J6
LbJQnahJdWsQl5iikya+E93XeQrk/LFxF6IvVPgB2+zboCWfUchHOCuHKj72wo+4gQtx4BtKjy7X
nvkPZqoMsPzMRSMLmbnA0nljuoGLeTc4Trihmfoph6EyJhxVfnnxInavO2n1hUFDuzSadGQENgMD
Uj0juitkgrqHogbXJnjM6o4LmzFIt+NMJB5m+6NOucJuyA+mSr3fII42Gp/MR1eECoB4hkjS5j5C
EvvTl7sZgyIWuOQAbk9H4KSHDcnuDBMmmL9irPBuGkqxKitQA8vKhnN8NoUWc+U4ntX9gDaXtt48
nKULkRst0/lBEK7QqXZe7+reUDOEOvElFc3vYyFX8fZSESJw1BYxYDDuYFH15R8bkrRIoSGDdndd
yQbY5KOAJKkohBKSkPbYr52Di1J+feK+X6TDzUYjA6a0tSRDLwtW1to004iSl2YYIgJIzGexTDH8
oQUlEuR0Rl+Em+sYUz588zp7Y5fVuHn91Dl0wCK4xSthqybpLJO03zcuEclmCzdYKN3nCX7r3HAY
mzDdfYPgiGFwAkbehsL/ieGtMNIPymCnKlg7QznYQZPw1s8VZ8BxWib3ONK4bC9KWnxzPa5f/Qc5
HgmgylGuAFRHGRnc++YDPI8rhhYOs/lTdNo4xOOjDPCKX1GEEP4jMNWqHYhK7+tftJxQnwPmmrSQ
FHTXIJrk0EswBYGVshS3cZAiabJCwC/L0wCEfipNP0M5dyaGk2RYFszSBRExQDqx0HhAVzOX+FIT
cEurc64e1ul4rRJrdBJyPnPxG+1EFnwng2d6E5yQtV67hMSQ+T3NdL7cCFOTxn1KS28LpElYTmCK
P5qOuEMmSdbCYtJoNHp2HPvPZAOt4SwYe5uTdZjJc1K9RUuKXrOv2RMcp91UpcnBmSt8UVlIzQvV
FVU6qAgwsFsZiwqaVR6fde61MPk6Y+YqbrMjPRKRK5+6pM5aUzg11DRZ+E+97T/Wst9XCe1h6gsR
7XBycwQ0TacG1cqOqngQhl6iv7V86yCnZ6k1rLNhgL63BGRqHPWf9YMgzsW0mYKhut/Yh58c8Mkt
wek3sU6wgVv+TcjOsmxhxATGlkmLQKVF7DQrgZLciYSK2BRmMT5TPONKTdHYZ7QTtfh5GzifqUiG
Yiu8gskLR8gUK7MwB1m6AuCWRDwhmZpyKNRYzWfBUWd6zMiz8WqVuuoc5BYYBXZaMzS3Wc0RnGg7
ELcZNbL4mcGFi0WckietWQwj1mvEDIhJcjdXko9YRPn33/FjOO/lkq63rhSExP6EyBwi9NFsNnnJ
NOZ13uNjuy7emYd//yrMB1fXnapsamuR6Ju4C30FOeVN3Cn9R9J0lm2+wWRPGG2Xuu7iEV3WDGNw
g5JrpnwuE80+LjnMi0UxMnZBbjt6pXPUkMwIpXGkqwt49nXSru8gZZQS204O08FOE87vqKMjtEpG
QKjYPHdFj7tT7/mqupluxFgLtibjXiCkIwHrUWA0a9UdsKTue+11LiuMIpvqjptm/vEBbZ47nsNi
yXwEjVBdvdP619P0iVyZInxbj0xrNGGAfDodmDFFrgQpUJ5WjKBdPFmh8/F5GlfdnO57DlpIG7aA
/fV2UuSh3+CY7aEimTBbLLXYV6GhQIvksbj+E9rddejcfC664A+bgu71iChtfHk3lIBM4vTJQtq9
sXOiJkDjNLctCUWB8FHd7YA67o8Off5PoTzx3GcfDuYZstEPckB/WLqszgNBAm3TJQmLR0mLI8hE
kcd48ouqKviU4FHNN8inYZxJaOFsgwl+WgAZVunc77EArIm0nBhnMXZNq+7s0gn4C72XxFpcqPNg
AB1UyJ5JHGMvP694zAn+UnfDlI+eT9M1JTbd6YDVpg6PSdOmHEz2cZL8vHVOA55HxcLLmmRC/4JQ
E8yoVIQlR3Vw6trrACYdwzoteJq2MEK/UVtn5DQ5j68uzxBrQMC9E6OAoHmbR7KnPg8CXeEkUx8F
Vc9LVrGjXEbLyqIBVPzVFyqyg7VvagjosiSbIoZQDQ8aIAC1TtC5ZHc6f1OcGa6q1lmNtejrhSak
08MR8uMFVkFrs8n8IOKCAV/sIwljcDGCtmRqk6jGDHpWr5pBZMP+zws75CbpXsH8cvVPvoPF4wIp
bOJ3jNHhqR1U6FQyRbLnWURVlM8mTIvtJgTADVvf/wCZBNNsgSPcqPDmWHYKMWJRBwr1nDYnp2zu
ZIgysxl0zIvoShm1d7yNKpmYmjdn77S5r3hH14gr+XA/4p0d2lYRCEvctU6CWn/XPXC9wdH92fGk
n3UsfWJ6Ew2TBCbCDfAFJfn7Kq24ggHXuPuNxq7DR+cLU+zkkj+CwPjEZyuPsCY+Cjxd3+GtG1ON
Wzf++//hpzPMQxg+uZWJXddr3oITXSzaRNpkJdhc3T0BgMU6sf4eF+ksKDUurV1PyeSe+xU2mtQh
RO/Ig5/vlwt8FjWUJSiNSQ2CvFtzCcl9xCMpLrFI9iWEj7vaHsCp93w6IIny5+F6TPy79WnOCF15
B+SkURr/i07ESlGta4Be6MDfpXZfGN1oCAXFnOufZ17/3pFdpXjdHmwQiUyUb1anx6HT/akFaABP
b+BT8EVC0K4XwYLr9VTrD26yKscDoHBpbA4QyQpw1n4/XEoXPS58QhbT8s0UX2R4gFEsIMeg5fvl
0/zFjRjntPNGpH0CEF7Gs/gl1d9nJzTeQ9yzZAF23ZalgKOSfnCooj6qm/Asizy3x9ucEl65aMAy
8QBPCnL1KnRvMxVubJl0GyhP7fPJ30DiVb/z6P9OuAGka8KSpqAY77dKXa53cUJ2fYuULgiMeQ0h
52+gXclaRjZj9PC+fJk1VFizziM1nt2OHUorW43gn/CJqFnjldTlRZP0Uj5T/wtzYHQB50iZh5xf
0UPcZAu8mYk+yzP5hnl3hqyu1PLz4+c1QYuXzBa0gyAWsgcUnJlMmFGhuzY2TWP0rljGZHYKpOPS
BbWuT4B82mfcIVS29Go5wabywAwlnQZsyS/UqUy6P5riJFm65wlkTYxcAov4eYNOqcw3PVa/8/5h
jL9cIvbzL/Jnkp5Jq3V15QMaEYrE3z0TE38Wdl3gUq1udRwk9rNEnnJfhmY5FVZftqLIvuspwnRm
SHGDGErt+XxeJaayMG3BbpUfO9/Llj/o02k598lxaTNcH0wv0doxAg1kjva3+T3kXlNMxmieb25d
cIvfxnsNpQNqXmG2hyzulRe3H6shrTEXLSfZunSte344A8TEGTAQ7GYaRqNSW0TqzhrwFnYFSnwm
U29e5I5BIwNshh8L4qcSJ+x6lGMZ8qknMZVwVBN/LR0wWWlQ1TeczQWbD3Ox6hcU7W/RVE3zi+Vp
PLDVCZE2leC9qfa/NKZKadNQYtcSkg9xXip7HATP6LRz1CbBIAVjvjeYyd/X5e0mrqON6JBDjakB
9f8Z+1GDPzoeV23TGreUebAYjnXFZnKigiWtMB0gwgl5L9bJ0qOrdr/7CadPnBdVMvoahYhZP/92
Oo1BV9W+szb/Og+oO2YmdfeFBYvyxulchnns76Y6/yj/OnWjCbgFulvg5LXcVui071nheK68WZ7u
856usmWw0kIRIhx1DFgt/zeVNOYY0SxEZRFAXrcV7K4xkbjHm8VC9bHe0Tw/qj+ZljMJBJGGeVU7
aiALlacoR07W+MdUETrnmMPboxIKIuEjNhKri3ZrS7YYCNgfiM3yHAi7bFMD5g96Kxl44A4eM6Rr
EEgw5TWWzAyR76ljtoA0TZfMAja58apnh7p+lQrdSMqqOo0tURduqjCXqT/1ZRHjfN1uPJcsCozV
ZUqugAKgW4QAdNHbspXeLwYst9qXRAVKOALuByDecQy/0UdqAI0eFvCySDdfRAsuwR4pJCtCa+Sm
SERULcdED7UgR4KaGewBMSdnMsuO7Kot6FY1i0qEGf7UteST8qJoEF//iUXXIrUufhxKmt+NDbGR
6ywJpDh13Ozu4hMcYBKAxMJTUeBcX4EYTI9XXYYwjW7BTzfP5GlHljxwQNKuDg7o7rdjvyLCErrs
NbqYiYwYqTOqjF3ZdrSRa/LJxGlGN/0nPc3Qt3Ukr7m7RpPBRQMETMl1CldfXp4BKe+euEPDG4Bn
jg52qsP5jx/3P8z74Rrz4XBYMwM4fLpDBMfFP45Fo+BTxalC3SkYv+TuUYZD/qdia0emITYMHikx
+F7u4vDSLBRFj8kcLM0p/UBZpKckIQxNljrpAaUGvcjCkhGY3c65zMPLTeCngie73aH+Hw02Pujm
aeYDztO0Xiqz7lnibvqkQZsG23jcTGVpZCa1r0eORJcvTS8RAgV+dy2UiTOOccqmL76q8ZVAunm6
6eph0lx+JVGN/DMbkGhtH5RnjL8pOQeXj1T0tcgtHc6zlGcegMWk7+P2D8lif6JlN/+l3YvtK9OZ
iynZwV65SAS7gFiPk43rN0iCjhKQG1PivYMWGRpBB7+VbUfA7LsIUcEemIG+5+hkFKOfoJT+h6SE
VXzd3YP5FDffvd6dDPBnrR4D2T4FIZFM6si+d2LylNq+gcycaJpBKR71uX0PqOvYThZacKbCOSnR
yFEVLJ+pkRyEPer93b+QuwhcPR00sCFdpMTQso0Pj0+95Cb00WPC3P0pykJacsmX3gHU5ZnBH/GH
yc5Iynym60Iq4uGt9sjLprEFAohtbCV1PyuQ5SXlHRgo7hlg9gaypZMn7FKu2nlCDn03l3oRTzSq
5RvxVWbSZ2E/X4GZZSO1BpjGB/F9dAE5G4CuQnXzfvzJ5rMQ/VNjwlYSjso3On7R/tQRgHtmsgtY
1IiNC2hvj+Xxus9ailxDUsdmSwiO7I1sagn8kpbEoLY/A7XaNYHSw4c1vNT0P7VgofY4pMDz2V5T
xRsDn/MXHLp9986yeujq1fuzjvOx9496/eSg9ifh/FDaHaShGHw/h5FWb+Vov6CVYSdEBuRXsgxw
3XVci1MGeDNyznylCrXEbm2LUuuNUf9b8JOPxjJm7YbgqmRNcBS2Ercw8N1jiyJZ9IvHsCqQhOjU
CzmwiCY6rBFmYGJE3aouVqUWEUaxjDDaBODjfxRtQQEBbyVqoHS5uYEJQBw6UW44hTfnqN8fcHXh
y/MGi2cLaYIxRoY7pRQ99TyQJyQErLzsDcUuBjhwuk5TgHP7eZD34sNbtxMDDb1EE7S/KzddzMRp
MXd1EIsoGUK6mJ5YzyloXy4E5UflxeYNUJtn43wAspk+44ts9kBGJ+3zum9x3wTVGfMBxPipLOjB
iruyKuEwvsTiCJI3gegyUWSN7mC9Hv2RJRyoGlnjjGNqi7cbxS8fYigcWss1vhUcL1H+maVmd1Yd
6WNrH0MlGzDMl+8hv8kvYo0oyLK3FwZvnPl2wEoKRIjMX+6TFx3JCKJerqcX6d2Oxp6cJQkDT4i8
cshIc4Fy1If85Dh57fG4BvoCnhefa12yzvIG3lStVahivk6ugJEvo72/Dp/cljH/rp7UfwzhFxsU
lVQ/kUgLubYH98PW/BBZtujjr58dO1ZjTCMHWWHay8MF0D3niGfAdx4eG+GdmNaw2eLv5hxxWimE
5MPx9IC2KdOJRaHTdRngjYX+aLeDFrsOEprSiROUWF5aQrI4lyOU7IOomPPwzBdQGfL2fBrsMxQp
Wknwavh8R0iMir2PF+cb0MASAuKPUThJql0zn87EhJBrYgof5tnUHvI8qTJUQFEtDk9Zvl0R3h5P
eAzDrfswKw6Cfi93Arkka5tWt7YEZ6grJbOFB+CAMF0NcLOp6ZV3QsFu7G/eTuaYxTAKcsYuFMWL
FiLFRokXyYyYnobB9iBDiXS5xu+KUUjcDiwm9/+levNCW5rIa5RjMLNvokp1luXZGt65F6v39dBu
6lLU0rtKFz/QnmSd4Hr4r/aZ+U+lw8zvnPFa33Ddgu0FSTa9yAxAO+bshJD/6rwTzHH3SsyK/BXE
2HaZSsXJA4zaVScXdqs5EERpYdAeDP77X2IJXtO/EV6R70byMfoR0h9I79cTJbY21/GNobuXe1lu
LcoZsiTwe5fdIOkTgl97d518ziHMmWBaNHmwAe6OiMEe4kdJ6WOR7Ta4MY5rvkWn7XEYawpuNrXs
mN34TFRQfG51zoWYcTJYSc4CLfAbRDCYW3BmpuzvNpKcujgFMMBF9/yLPFTfN9rv/4jTTdAr0Ghr
8XXDTUYzGRI35dLtp7Cg0HSfXzYiWr1pPaXpZlvA8Rpi7UDL820RxSc5FN/AcqcP1hlXP/0zSFCO
Mu9KcSesX4C9MBTqVNvkh8nojwMHndeONn7PAD8RQpih6m4m2T/H86LqPT4/esQNZacjOZK/PEL5
9l0XKkP261DOk+Di+3hGkqgmA0Jf/eqWl9BMqQGCdKX4HqnvsFiwv4o2EM7/tM9FMVVskvSlfaup
hhrhAkEnkeQ2lBjeCOaahOybHu38eAk/W3elA3lPAn9g/sxqRE1Bw48fa94QhyqKj0tNjvv5Ac+S
Q4+o19kIciGPSnMXN5qnOmseoWM6apZ48CamTBZRJUEX/nVSKNDEJNG3NNTtD37I0FuT6MjKHbzl
DdLcOE7zdELIzkrdmD/zfVTJ9TdHw6os/r2aWeU2XzzhznGKW7yhItlKXZY4ucmlHegKkIxkRgfr
MfK4pc3FVlXjOioQh8Pv1wyQpXrKfisuLyPOiBPCxFGoGoHH+FCAp6VgUFQsrGK38eTx+/g8UXt7
kDAd7rSC+T9WGWsQC6k8rOMFSAyusLijpZHKbqX1MkJ4OACH1I1gCQ5zjKiF8gxLdt9iD7H6Osbq
uBngP7wvEIcBFAZRZ/HgPJH9Dp9VJ0gzcsE8x2ptphF89dV2ewH4fERW49/sM6CT9oESF7lkvypH
Tc0Vm2nkvRpf9ImLLCc2PnjnIKqCBj3SOGefydWMHhljFTKj4K/71YJkN0rFK4KfQvfkY+ksfg2t
+hxfEBj2LZz9fAjF1apCH7dwUbRj0+ALlAJHHZAhLYfnCeiDy0kDxiCCJKbb8Kkn+N41qzTf9TTj
oFaH3ffB0/lRhu7gdnfycvQYdeS4fc+Lk6ipP6Ctatb72uy3HoDOlH9UKpo/i8xPuk7UKkQbqSCV
dm8YqJ6PAsycaSgL+/ZtopMHISVheJLo/lbSg4UQHKFcgtupoC11PW2SQ/yCtUkbB3DXWPc0LWjP
YzDrwwZ2+UZ29XwzEb9qAaUOoIAziOTrmE7XS4y3bhioRIiRVuzFwAqMi797eiwpSkouyM9An58A
q272+/pq1KmrNI43j79HkfXVPvwgiFH9gsVXwepyWX0hdCvXeD89SkLG761trT9nzc2Yegm+s4pS
fIs8YF835OcT7twPD8+JzzS+3yO0/Jy+lQysfTmWvb/r7do1Sab7N325GGCg84IBC2xYJII7qpxc
tH5Jbl0/OBcBRFLyexuwvNjrYURRlwObJN1NA5mA+OzyYjg2gPmiId6fsgmLqDYN+2DxSFZjUfFp
7FuxiLUIRnQJ1W3aT8vnpmy35aX9sls3cKH5d+IeVrKRD2uM4iqG/6+bHZg4pMqx7z/45PKISxf9
RAzsfmgu/oqvaVvchKiolBBpUY3NfvLBWBpA8NyLhgozeGctG/0SZBOc0PfbesDCBDSy0DekIIT/
ORYwzDofsjpb1Kovt/yXSDM2hJH4kj+dUMev0T+TMb4xWDARKlaiSYU7+RR+Tkki6r2F4q6fIZ8t
El3XMsH4fMR4NO531Iy7fQKPzr0kAKXKS92LJdPKelN9+y6XURnLcklp+a3UkPME/lvIe/QiBRS1
RQCG0uaF+L9DvddG3BtRMd4RKOXN7Ro4h8zTVZwfYJebvEzn4Cv6VXvj/SMxzVTWFtOPnlCW42Ul
+CGVxS4w+mzs9MWJ7zftImItCfO7tQ2M3Lgp7bAiVpgMJlMuKMJzCp1d+ibnwL1GzlL5cWcboBFJ
lg8991xbHM2fIiTFtpkJnMr8XYXCD8lwOCDiZtO9xcaJn9C8qzcUIVL/ygPZtnLS5Rfm2AvnOu0N
IssAM7BGdKS+tmZ3qrVv4NIY0pPqjHBTnUEMO6BEFFei0WJ4P342iz76cKDRUcWd+3XRbXm6ui5R
HujgcrnaO9exUncs4BMgLSTFj5mXW/mRoumqd/tOE+SFFHCxL9uL5nzA9ZNSlCSqtszvgfKg2wlk
0dTfN0H67YINMlkVr0VRcD4BLN1D//VlAMg5FcrX42oZpOpTh+hUahEzkiH2TIkqr6DqmWYZhfum
e6GxH6p0dNDUGQ92X1kanMSfoAgdhiPuVPC7DLIfSiOCoCsHtnXxpeI/Gm4CZO+JZiNVD3p6LTvg
NfE5breqR8B1LqT7tXHCq9uFDqHk/ebPXqvCT8zo5Sc1g/KlEV11I6QZGehgtZ83QfCZ5gwFTs8n
fKo7eHllf6yml+HEYYQRBs9tcPIkk5gLOrX0b7FAFHRG4ULEvo0xNLGW/bE0LmIVpRN3vsvP3mc8
aKmMaMyXmIwnOehEoX8+8EIpQgLcbNunljLp2fzqgewWGRB+3UzwLNZ7GYbZk11KNlbjtaRKbuZJ
UJFtjU1agcIiVfcUwJDiWGRrC7MjfZPgiIpgltR6l3nJ4A0DkkmTJDqfQvpIPXErxfvQQOZQq0uW
8uxWidG+VMXqrTKzCMbhMQ210DvBKN2YBpYPWFn7XKPMtxjfzLrPnEiG6odWI9+E3TBjASPW82U1
I3ILw6I3cxjUIlObpBsx+98rlttr2NACg0/vtS81NsJVx2cfqnxyaTrho332voMbxiYwIU8fa0QP
77iO4f25SRrNcP9+UuzwCXAu4ZUO7RFviiI96TZBmEk4VNGsffdMMhSyB6IEPWd8HO6KdHjxH1zi
/qTal6B3fB+W7LAHwBAS+eKQHqI9nFrU7rzk3cIYIQmFs4gE4s3E5uFP3azCTEgX1hAX0gpjkPZI
ozSgjb8O124TZtHnEJna1VnXpTAcOykvmdE0eAJyY0y0LbsaNNxnMtyHhC6buJih1CgkuUzlxZ/j
bs6O2UxDLJJ2k7w9o0K/fLGhnGE1Qzh0k3mtWb8juKFx9bZdLn07Ctd5lqaM2oXJYMhc+M6IBBzK
Px6wgHgVnvE0ezRUswmRX0tIIlrZLQwfF0cOQFS2c2HVadDTH6dkFHEmIs/ml7VrJm8w0FF5a2K0
BX9Oq2wZ7imHJjSGvwWYbdg6Ece65C/Q2PMlFu+TIin1UX6VjRr/N33HfuCCO/wiN0h3pkJNyath
1uVRa9RYFuAoM20daM3f0oNU6onlT70aHC4o4Qm8ApnrgXPGH1UPzGhTVmcl/PLyBfNL8yLhVE99
K2q55AHEj7Ev77QeAyHeTByQ2CvEnhJIFzvvW/CSwWZQINle+Dyc0pmDspyhOqooRS6NM7anc1EM
rqbzU1RHNtXr7VO40UO4USveT0WxM01irSsNeb0u7CKaEH3t/lTDdrOdKy7ALQ9/JU3kU93tWuP2
u1YCiJm4ZDcnymeZueD0m12aYp5jF9Hru0PPCWIGbp9ZA2yv++pugM2CvWPffkqH+wI1n0A9YEk/
s/iU8W086/AKFDBi/tKe23RpY9vm4IyalArRmdkxVh3BslQFgFqkt2gGYRfNEx0XrSLJzf8KN3p2
7Ng/WnsUffw2pQY//1bf7XQE/HFKT5JSen25H3CaYHsYh8BEEa/lyFLI4phaig/HrO6doXM8SHsQ
WBf3Uiygm4U4yiqXm+zk1iu3MOWhNfFaB0oLME80+WLpQ5HC70Et6aq07y19nJR1ywO2zY0eSTIA
tu5WLhyQ8zKl4V+A2pagPVwsfa4BoNN4M7yEB69147u5wyzfQjPrARum3tPTyXU6xyWTE47krt9h
9+99rOPnrOloYeitOQ17CLBPyZitwMD4KSZivqKAl6UBGcMF1TfauErs0he8gs1dTNsxVl4DTTPg
heq7Us6PqKa6UrlxbqweK3dNZ4uyyNFFRq+H239yV1NIdgUGGPVU9GSlqTkmqkj4F5G+XK9tTtXD
emcsMz6Yoms0/UGF7Xok2fwC7PpXhYi75oR0XPesnii2wnlGnk7oBzxl4lA6Eo1bb78TdxQAciCi
n7e9jrs5gjQuFYfNswUSMExXZqz/8HbcjVyNKQQQNqkpgow9V9i8FoAn8XT5bgV1PRCr8i3HOa3F
GhefPtqW6t3dzCwEl2tMcCrAPKSEKZRX4bbQP2ZUHbe3T5r71uQvhDRYQqFXcinLpUbs2iGOjEsF
hmu5tNVPqbyqY31m/bPnYmTgb9X2mduxB221zqiDKKqCtfNeaUhbBjCvQOQSGTs/9Lm3COd7pSna
jZDNROPg5MUk5N0JCy9Itu4wxcIoGI3FUHMWXsW9sIKguyqylPeONY/x/uoa5XJrb+CtdaLcRQqK
WA3IKrDtdyIv+F1puewQtT44bxIxtVW5jy0a9/9gIiwud4Y7mNF2BNwV7Z69pJRJJcd2XioeQ8oA
gAxxAD9ZpnzFF32ijYWVj5JB//+Y26CaIl+oRQ+KfCWyDD9jPQtUpXqRaMrnY8HOWliYarpobItm
nrzEajZ59FCJVwVu0dc5Wk0bqKa2fjQBRl3Ks4gvEHesFiQqLH68F36sHPzHRaQnMHkOEVuDuAOS
0ZQvoTUBxiOQkBLe7MB9qGQr4ERyNF2siVwlGbiVX+DDYchb7ETRPrpUEnEtoPGEuI1GjhkR/hVh
8BLKo2B0JWbk/aAGfkv3OidfpjPa8aBmhTHpJh27msyjaf0EVZ1Kt+KV2+HiAxTzjcRysyQ0j3/q
ic6Zaqmpszq/SuKUK8eAflzawcYL6X9wpjrTji8ZSIwZKM0GdTvzJ9d0yqD5mzcDPnBxKaKz4j9o
kQa0jpWHMc8hioUPTMsGVbu4WIwW+xbet+ZS1Xzd1sbcUz71F0w/+Awr1MnxmUnwW0WHolMgjTTa
siojubHHW3l26C37KNHWgKQlnG7BiVLEr3XsqjNzRff8FH2CFTjDzEB3tEcLtjTHhRr0yI34s2Vm
qleNvc5UNem1zBqjNPTVX+pJuYvQ2+s/E91W0roq0gFrXS5B5lWNSZhmsXt3YmzVev1P9mvgz3NP
ZQX/Zp6xmTGXyvZOPaWkSduUv+I2uKcWaChCOcPnn572bMpmG2odBQquJinyDvpjZS/A6/GfFIfN
GbmUiK66ucdxGlS3o8Nk+3bhKePSGGkBeB8uf0fKOwe/KUlXUUs0z34jfcj384jrTwsfAsrl6Re0
q1uM+AYQytBN72cgBEQVUoCaBB4KW4qxTd+hG39LZKtCNwVdFiMXhkaWcg40gMJimieDHyVo4cm9
t2BLN5Fic20VO07BstoLSW/5c+7tJ1R3AhyVGIWvG1WUBxHsQNKut1t7WHHP6Ez/d1sWLo2kGfwN
qd0Dc0T1loEnj8fSvcJ2cWJLbQGvEHkERfw6J0QsBIN1GQgHt1nwoppfLy/KUxh0syxDyzdPsndb
2waxrfnemQbxaU+79UNfhQeRu+ed2cQvaedYunaS7kolB6MUTmIm0LqSLi9Ao7tgJCWO5Ha5uUCJ
ClX/00tJ5lqfAyt8YpTkvCNpcNEh2Vouv+xcxbqszQsTO7ADxXdCmgACG4LfYukWL39NJCbLdS5l
L2kmcfxE5b6k8kAvFLgUewO2XIksrnOOjHQgDqH1Ou51TgOHkR05+84xJLcOM5WveTmDUQjoOYoR
Yh3hF+kaMxgzbYdz33XAkvxcY72M5SYOm4JMt3bIxBTfOCAYxZQTfZMRkN+alzbtuY0EjGmyDPC8
WzH9OUpbkQht69tHbzvvnNNc3/FmARqnR1EQ0RbD+lX/0HQ46ul59aqhDzmnKbrn31FqzOuy6hy0
RSnu3QFIE5Lk3Xiu3udPSHDNj/IwO2rMMLOKGaSDP4rJ4o5lN/r+OiaRI3DE0mNHPrgU4HuSSKG8
BQOlDhX9kQsdER6+qp5eJAx4HNcNUk46nON2piTgIdjzAZiXst8SbewuvaH1Ie2EJFObBu77K+eg
lNRW0xHr8/UO3HSTWLe9WRjK5tpfD0e+dnAIl6qKHvam79uar03sPi84BFRJ2BB9GuzzveTHndZG
lHQcn3j1iY2mJssAeXH6vordc1r/Px14ch/v8+VtAWRfNtRtrSXYAK/HgKTnJFaKiairU/1DveDH
1UR51KdihjglJB/CemlSZMXWEVpRT+mzDSRccB/LwFu9AfsKttPUr5IbXEFndDZJyUB24lxX0lmD
EMGhSCXNC404BB81A+LOgQTwMVki26LgsAJyWuSj7SpCGZ8nF3mUHoemvqqnj7k2rIXmEjcbMC1t
25bT5KzuEGuB/IuFJ/SGAtTyuTHl72QRSprZAp3naBbe8kr65fapVf491FM2fnlpYwQb2P9dynvI
hFHiHmhotxe/yHltHq4xzS0MT9qifzDstitcVBRs81ofRokAtcyuVRwCkSsrk4o36JL5nK5O8AEp
+S0wlpRovUPAdiTUVN9N8Gm8wUwEyET0USd141dT2uKCrG55IO3dzE/CVPNeaXiYaUn3XltKmgmp
016SW+hIEiSwHOwNP8CNmfm224PtSiH6RIgKOFY1tlaV+a2qQ12za5cVLVTS297nwV59CwCHurC9
TskwTtjqCLaAD25bQTbKe+LHjEzkifAxfFuv4cRtzBtqZQ3ElJV4fJo9KRi6cNeqrmRcAT770KmL
Hoy8CffL3RNFJj92kZ5e5fc87JH+Alhy1lTD8Jmon3Hx8HZIVpYfFfUA1B4G0cMdCAc97j54UJbt
zc+U323rOpszphCZWLFufo1vzXj0tKBK/FFqZ0bjnfzFTQa6OpjBYKr5t974cz7s5ld+gB1Nz9BE
yWtR8KhfXpkW05QCromFeVWzQnDhGvLBpjYg4dhSbjzqPXVIqiEWWSywZp1Fmd5i9M6JypoT/t6y
D8d6c6E2UagcsrfUpxq3bKHU7VM1RUuqeJz38nahHfO9a3MirriTXi273OTskNCF6fVs2kdPTKvY
JwkOXdEsx/Xes1EOiFJ4Puzwjh2tSWJsZLdQJumhnfGMT5Bh8eIVVLYrMuBD54JNlcUZ3pf9F9F4
NoFyevyyAm0smS5sDnVYzK1iU9Ef+GcijI2XEQ92sgKatzYSC6CETGH4u1Ho1oPgGp9KuCwtymKT
tZFLVqT1kOfKt3q7gQHVRuNygiywvuCGtCN+xkTzsxbRZ+a8sAZf43Ke51zyIf0UYJ3KJ0+7rQ9o
+neDlfjZjyiBq4O/Z+DJvoqk3kMj3bpAp7arygKAivtCF+wMQ37wNOBvR9HFuPXp061fgUZK0Mio
XK5B2eANnqKQz9MXAHI02CR65/4FizSXLPVeCzi39ywr2z/LB1q/sRQX5gB8CH8NUC8DsZ5yzz4a
JwDGc39koPZtMj4yMtZDXVBc7yW/Z8u0Ur8Tn18EkCKI+XIzZMG2T93FeoqtXwOiDKuz4wpVzFSQ
k5jszKDoNSFz57vYTB93W1xJOwqC6UcRgBpBwTFQF0680YYKZVpBgL4nB5p4yPPnn87/gSKKZKr0
teql3M43Zerj+fYBf6Ucac2DlNU4eDpb4keiUMDLAJksve7xqoA7aJtMGRF/oqu/b1BuVQKI+QS1
DvmXrtAMOnI5sG7+PM+3pwWnK/8h5GcbomZQpw2NDALyUSEtDOxZ7ck4oQukpkoY7dUKv4UvPeax
xd5GHc+xb9sFhmgL4P/x7Eqzq68SKNFwZ5sIbQ6Fpqy323w4XeVuNG4TPjQGxaNheblW5RkEYfWN
WEAEdGus0Zo+AlOi0EU4C1gsvwhkFjVLzEdZwt+5R6tUggRfz3HN1dKjAqAd0T7RNTDJsU9/FaEc
JK4BXsaDmgV3PmlBPXp/sYlK1saIjw/XpkjJzeNyPYu2tnKzlxpo95+mFgozsdNN7JYP15OZSxYf
rYVAQ1SVOjCq39oa8Ak+Znl31/4C4YYyVOprK0qeC0FHREfIyiPMjKQTmsP3clLwt6lGZ8p8mvMy
eqERdmOq/16csRj1oxyVCgYrPBGB7b22/bnZBRuZI1EUGWYGoKYQaM6/DYvQZSgcoYMKDYX27glz
HJlOaAhLPvNoFAciFHhLm41FrA+83yUi/iX31pKxE7JkQtxmdbOrgspt7LLc5RFCv4x4SyULtK2Z
kBDLz5cW5L3CP+NFMB7NFBXIt6x4xGNw+VfsihDAGavbJeXygCbrNASp6Ujijao5bFaWGrqqsl+K
S9R1JLMKAVxSObWWRQsQ6nDAbmvbdt90qhQFneh9G3hlyMtMAAIrQA5GJTdIpIGPZ2LEtc7hgqMW
4H/Gy3LSjpKZ/9+tWcpxT3oKYKCQTxw+YqLAMjtSVlXDkAJb2PvjkGXA3FZe81madrigUw1gIA/O
sOnE7t7VhVFQc/sOo4eARDYrB5XAEJ+oMbdysi0fGlfptq5tQaarPQjE5w+e6x967uPk2Aisl4S5
95c3B3rh1loE9fry/J8DGsY40cqCKvufSBHSCvHt7xl2I5N4roKaKJAUs0voh9YKYRGFhlwt0Jhl
Hrr4pOkuXSjUL44Pku90KkNoXN5ea+0sozWqxr+/kAHQhKH4aNc807gQ60JBCOrFPUFI+V89AL+n
ghw/dtg5IHQbzZltdKNIg6HLylE8A6h6e4p0PbmMOhqg8Z3ZfggsLYdLOoEsQAb8QRHcSTYkUUJe
SJdJeNapYovgEdoUrS9haPYyBXeFTTm2HzRQ355AxRKrRRMr1qjvsK7MwEcGp6NWK1+9WVeo5Zex
p5qWRv+rEiZ5BQjxFDThPmxJSewTkOCSd0RCyh49Yimif+kyiHWKHe6mlSj6/JcSe1rreFpcnZt5
3f8ick/eFV5yxhfCS7rJH++nkzhrVfpn5K/M5vBWCaQE5VDVhynbFOdSTD+stRxScp0if5AOnmEq
/eO4+fM3NsilZfOjpKP+X2DJ+idZo3AeeSVEDidL0txHDVrK6c/7W7g1COHWxuJglH/d8Z5Lwmtk
x5x0FUqUk50UxLF56lmy00kx43htZHFBOOTiKVXvjDKTY31TSYK/s/BlfymMfE/nAnhNB9ZhpolC
enb9Sie0IlHpMuMNVCs32j6cwq9uT1r8Gl98DNlX7XWjyY6WwU2IQHNnkNfFQiYeyc2RdQNsmK6x
co2DazsuO+nepx482Hd4+z28JK91qCPPAAxzCqdhtn9azZrkEmYJpyswbpYPDweJCnxeKM0lZFU5
073i7ksOiJ8x50iOaZLhcQtheSiy/ABbZoNFn+f4sHEi70AhRrHmyGK+cgWTqV35jI2eULbo1/j3
0FiUA0EOCZNKzBfspAHJtSXavZJ/uiv6s5retQ4Uj6z1PQnsJnARjATN0qD60QyeYEdjZ3Fn/aaR
DPq4xn7rD41P4zznyLAVsaWHTw8nsvUvNG2437KiY7vwLMu0fWnrLo1pnBS+RFoY7g10rzDqdHOn
Qlkt+Mh4MvxhZOSswQGMHu2AlW17yR6wtosBcROO8vh34jXsl7/z4UWK0Qfh1pRsuiWfxuYzS4SC
mQ64Gjqggk7T5WhAkbdTZPI/ev5HYH1zXZ3xUUSGanHGdQO7m+hj/b3+agdBwYfZdGs5C3XArgfS
qeDP91IThbpLsuQ4wEDpOz9kEnImIMwtgPIf7gVoRtfkFHEPpVoyPM6ckvYzcG26uoKmSESgWT9r
XxYWAySLOtx8LBs5TNvAMWTGCJu9jvQQp88SCVjyhralDKLSkvuM6WP3lB2XOuFK3EdPmeKRdPBD
YjK+NDmzs+ksStbqpCJKLlf2xlqssBiAzlUSDwNO4xUfx2GHDUx6DAKW7XOEGi5FhWL8B5IZjBWF
rHuke75MzpiMWZ0O+IUcCwdahEhR0A3oFM4j+/jHqF2b91UOvYxZ/9D5/ROcQjeuxP7e8li4H4l9
del3KR6hWa5jE933zSById9UdSaYq19099IJn0W0gpSpLmwufYjFSLbV+sKmwdmP2r+amYgcqPPm
3GrqmmbG1mQe7ShXmWuIw4GLuMKQ8w4g7pT/suLAm3lPpc7XY7WfqNr91mXzphVmMdUlYK99Vp4K
n+Ytu/07/9agVn2FWIiP6LjcMTLVAsM5v6AIhwMxcRxG51035xBT0D28nB8F+zIJd/96PSuTt9MK
VT1mEh2c+F+o/N0gKqj2iZ4w5r/jIkZjq2rVfeMKJ+S+unbwL/OhEmNEUVL3KmNmUC1RYNsJRgrh
CisikhtuDOplA48BlkI1Yf/tZC/s4n6vMdYFNtzOZnL3k47NahFB09CIUXIVNPPtQGv89c4h/mFj
7Zs9Glu2oY2O1B+m3IENayhLcQXD8bijRxrFu39zwglKYQ00WOJtcLOxRi03faGF4Ci3AZdJpcLE
8Nnt2E8dffGV178M0O9mEf5PKh9dy7IDwXWhwN4jmWGnwwLXo2UvWIhqVZhB8N/OiCMeBK/3EU96
lDudDcy7qpJfAl45lm915Sy5bKh6GDkkwe3YBpTeoKY4jri/pbM7NtOCLyqimrOUW350IvivVVpR
N+wkg/3CWqEgCBwE6lRSGiqlIpZ+ji1BfNVHtrteLyyN3b0bsvY+S3FDYXKTrHI6rhRzBcaD9AqV
l3SlYXhy412Zxwnb3kVmeyUAufv0MwIZzo3dUe19mbKoL2SecpxQe06xwm4hkt8RKkWlZaVjsRes
77IN3RsogYVxZJ7JDR4/KR7b6F08fUkhNMAEqWRGaq3/VxQdHJFXFwu1ucvhKSAYI/cX45nIILAE
+4PtpeHBwyo3tLmuDvAfxz3rEnwHy6EhWc0ZWQaM2KJ1Ntnd2d64TU3MJ/12cCEEEhoq2UCQXkZK
KONa1eGAYp1N59lr691adrtahgt7TT5iamlBW7RJRKnem9OqJNJVZjL9Eu5BPX611DMRKl9dhVRc
Jmz8J/Q4vf5Ils07Mcc3T67qKFqUNn0h7KHG5BfWMs/EnBrCLPA12kNVdhwfR16aMrKrVK02Cn9m
F5jk5NIW37K0rkK7kXnUkG3q8/TUK0Z8BSXmLckdrSdd+MfwTs09Wl4sEDzwS9IfvYH/i6k+Ul2/
l3QOEqr6VSHvJcY58tO8yK1DNGTalliYQg33aKYEsMM/kV/YG621ll3rC7pLnsvZftI93oDoM3P2
8tTCQIZKppO783HAtCE+Xf8lMCAYHgGH8RWiaNjA4IsBuiQINlacYQ36lsa+2uqh5n4exIZ+yUE4
7uiKfsrsXYWt1V8wLBCMbYx6gI56OQoya3SdO+bysi+kXO2Pw05saXqqku7ISeGXimtve+a35R5t
LKDfcknAhZaRrHMNS0PxdQKvuJV0KtCp7UIqdQws6akU9J086rDcNLXULbMSxElGWJu7uXNSuPPk
EeBA9WfolhSPIVWqNPrO1SKBJQijhh4g4Zt+mWhrpN6Uf4bqCQ4fD2nM0ibv9rCdkaR8sOqlCutY
QLXtB9jDiNRz+DeCQL1L24FNUQEzxj3VQcCCnMfCEcuH75Qnnp0tJVnB5gnsuqhVxVNrhjw947zW
YNeaE9Lu1X0Wg3BIMBgr0hktlD00TPCWKacPIDlePJCRGhGSIZoJWg/+uLZ7E+jBkkr25Gxj3yjd
iKS2uFy0EjTB/86C7VpUTtgIbJNe2kBZm8xNktkujYmR+2r7orqukR97XV83PYAOYeCLBdAVEaRO
8aHhZZ2WLRo1obusvZ6l3+G+mnK2/oC4NdL+MkH1IT5PcgMV6BIm++WUjtsZQxXKaA1srhS8SoQF
3obnLAvODy9ZgLHdnQUbCCWccPHuUV3uzPX7IlPImb1c0TbpKdJ2xm/2LaMCW/yHrDYaNVuqGsgS
NT94zps1NNGPzY+pHMdzsTNdBZCjOMA731Mbm+eNGt9qDC+tGOBIk4ghB5cqfjkmvpO5CBLAF69W
NhllxaQ85KrHxi9ndwAZWXSBAPRZqhkUlWQ056dNvbeAlTyUgo3jmt7sKwHtQeOIAhmS4x+fwhbi
lU9/04GSa3ae7roF22xJl6wYaUNLw0faQ6utLvAH45asmXbhvBsQq+lN7KQ2uidNcsvWCJDVADnq
7n331RRBPZlI2198V3LTjsRg5Q6M8eFICj4WZo9QxlwqOXru4q6pJuR4cHFJoAqWngsawwGvdChe
Yf+McXtjE4ePWvuWNX5a1ut+sk61tP89ZRW2OFvde3iEF8ed95GDYulxkmaUHVr8F9n0vrHtk0Ou
XQYl0u5EcsGGiK5N4MG66kMDYgeJ0LqP2Yjv5oWtNzYNYURNH+K+J7gvy41Cdl1F4r9toPDhqkq/
URdaARd9Sg0kbm4c98rOPoSp7UX4NUIzUIvQZyFvjU/251t9mxqZX4aq2HU45K/izcHcKgHe/M8M
bIonOJK5KUHHQqagtTKmZJh75T1PRiTtJ9Wxx78oMWw/Ytc10L1LHE41YPbwBZ+FWPzNiO4JdrQI
eY99Qi3xmuQGycuda5HceVi+rRnal+JQF0yacetT7VIo95/ZHPiH536MmGVeJ+ayKfINvRdGNs3c
H/cw6iO0vN7ALDLMah/dCt2fTTUbkUWoaj8o1ETaV+Mk0kHtMMfh+omPwOfT5B1C9mQzQLM13ygo
E5PrFcHFUx5J8zSCyRic43I6T/6L/+XOBwDOk0ENPsiTuNCNBzEX4EE7xGZEUodzTWmmY9BVq8Mx
4PtRfdi8TUagdqvdUWYB05vS3ac5rfdagp0f2BaEVNsUarEO++NOEjRsmxvOcc6lvYb03GVh/PeW
qdmjy74+siZBjMP9xn2nA7K3+j2JFGxDGkyzJ87A5kJliq/omxhZ30ulm72nT5q+vYSGU/PzpqHY
uROG2TCrHDFJbLPYJCFP9gvZ+VsXmXuOlNzWp/ohtSrLhtQnp8GcAe3PzkG22Zt1Ems8sd/UA/pM
tMhBK7u+EFT9+NslFcLYOJzCf8WCrcwPVCv7zuuGMKYWDx8VjCEUskjM+OOySW7ewx7qVHQ6+MfP
Ud4uJ0+YhErZeKv3/UIKH53ps53VheApL0nn/Or17ftP3OI/hLhiDWO7NJsxGsat09/EpmfVue4y
hyhy8X4LlCIR8q72aLBzE7QQfeVp+CuZPy9buc8faVWFmqMzQkPaByzFqhn9WoBo6eITJKi4x734
qY01ZMWXlNNPa5t/rRWJztlA7zIDOlVSQxfuWe4U2y4atRGBM3H9f04iYcPb3e+vTBcIYb0Ae+OR
GXNIIa04pbMsQIg04NZiEjMn00Bt8vOiMvZfIXFWQSsTao+qRHlXZ+6f8zj8NxukHZkNfz/ui34V
l/NS4eQ7ncnSuXvETYYd2uHgwjDIMPprgAqYtCzLYHOxVGIy6BiqwEgkp8pgrWB26ZXFNB9Yz/BX
9nvYAw1r0wxyAZKs3O4HuHDTPnoZyFXq0VtVvrjrioxpRABlf9h7lkiYZTTGf8S+tPcxOVHnIGnM
bNuyzos5LXZTY+XsvqPi+OCh5xDwWynLkxI/E4DriyliOgbahAoLBdT3Fcd462Wz5apHJf6qUuG2
3RixRCF4FO8cJXxBAXsdjelPLNxVawrX6vaNBwqoJlIoOYy/O8ch2XlhdEY517IjVCEXO7VUf6fd
Awq3H1obDJtsc/K3H3hqu3VWnT1HOCLu4AxXljPxqlnOkTAyWeGrhIyrUdeMJHGXhMbEcaOOst4n
PVt9TYs71JfsK38zE8dcwJnobgguRCdXTLWg0qkImh920Lp25noSjdKvmr0kaQ5ixnNrFU6RPvq4
iifX7MofibHeHGgNlIa8kFS35T3G4UEatA7XAgbAmSLBQq9aNiUOzxe0LF/j8KbLIALnA6GfQz0o
jZjwp6Sq9gzYLI1Mmyjn2lTGIN0ZmsEaWZBRKRKwTG/sLMouaLFGwqewv2ZG68UVY9dUUiHT+/jX
W4jsYrVvuJ1hQxdQ2qPOBC4UVYdblp0hAmWMZu1fLNARTOn0IzfiVYWJf8RIOIgLAo7pEVxpW0//
9JO5i3JGmqjiDwn+vStrH/W2GJ5PtOcx/aHXxn0VKhS2EqCV0XCWM9mz+LNHKuOLATEtfOPHps+i
daQbSSECDurGQvWMuliYA9od12qxtC58++rP64mR794qZXat7hym3FaK+j59fBsBUQBJJN5ucVSo
sxLzwv74Wzxq7pGhARaKm/5UQuY5RtHMrb5pqm/e6CKtyZ0ZekAwzo0hWd4fkyCzssBTEopRKdqj
LgLSw1HwH0y0RRVwL7LPZE1qeYvmF0Zj0YQbROS0R8wudtTK/2s5Eb60uwgv/MmytXPMT2UIHDkJ
B4TLKMKGt8ANt2zGcsoo80bAFWj0bC9rY649mKWrUNbL6n83WYb5ovLQwvlZ5tfa2ma3zPczyEjK
2jxwlTcQb3ohDtXCLil7OzZ0Sw0m7+gtoC6MzcF5jdtgVOvEx+SrGDQ05tw9YHTxm9fDQKmFL2ET
RSMdUoP6fSHFcxXeEYlN5woqcSLRpCnsrzAkjGZy1TpBQsoxX4ucEiiir6lqdGowoK71nbkZGhXc
MVURe89WaxiCFYdtuERg/7zdlhoDuu1cPdT3yyN++V2TsU1xFVZG6SZhaEVdbNGSqRXZFq/7cEjk
6p1fHBEslJcgS2ExXvIoRfurxP8HsBuNJ7AR+p0AYsVt99UAeHJKuaRa8QjFVg2BhbokcHr+s/AI
Xzwty3CQXVkejkb3Mv+r89OTMjwnp3/G6OBWa9nu44fwcCHTOrMSiGp7mitJXAgA+GOuXxlPcJ63
oIPZUuiooiB9KfEzZGeKgmYUfyr4f/ICNa19c562S2CUabSua2RmVmFdv/898cJ1rYwRwv3LTZIQ
KWMqD29ZrHdGlDA3CCWlvUFEQxa9KT8bk9BBFoS9De0e/TrtHqNW2yXCLywE3Z0zBHItPTuOOivX
IlKY+Bsn1jBSiyLRcrdsfnjilUUvKrRyBpOeswNcs8mpvdaJ/QnwBzxN+kW52Z8mml0IZwShEznG
6J42uu/xbj4B8tTAS+WJYrjc9mTv4GKKrZKGLzHwljbsjtCY2ysWE+wzRsAtO0hvrf0qA4DGdi9+
4bsFqhhyC742KpvuuuwDG2AIQC9YXvK5zf5bmaxEDcWGpe4ZTBxGcQB+wLETn8RFbcp2Fu1WyJjX
qc0Nkee8NGJON8uJeZh12l9XfcxBGIqsECsaSQpbTaJba4uSkGVVv6pxnCIZxdo9mDMilIZYKs9m
oNtWuHlA8wbRuL0cRgs0qrr1zTYd+9X8Py4hiDlgEeJHjKZIn2IObRARWd9fbae/auREtOcJPGhm
fPgxmMQ1HU1hlNgG/n156p5YmIXyoNTz6vQh3wZADE2Lc2pt1snbS2xwEdJwSt3WasPEM3S6mW1X
imDMPkCLl7rKH4gY/5l3v0xJUCn8d9+Mui70tmC4mqwjeByVDzqCfUiJtBWpsBuaHvh2Af8Lh69x
QbQ81dUSTmC1vngeEmFSGW3pqn22UEsmB+Ph566JlSyiCAlh0tvDxuA+jH9wPGxijZvdcjGvcqLu
xYFDTOjrjV0nWkjiE054Rifbuf0Yuqp0NnlCoDG2J3w8F/LJXYlL7kV3UrEbadPpvQFshd2oU5uq
NmangCnyMQ2nj1+oUKJIahzMhDNF3gp6P1SkqqTHk0dXfAeEK7hH2fmmPH08hHHrVo/Wi9pRTTta
Fm/3pi0bLbeHk6aspGqP1POUzZxTKS9jCSmDSIofh58AmEsOiv5nwKNZ8VBTPiPxgujbfqza1bIS
YtXG/pSgKFK/354SVcA308OTVI/G5w6lG386KoXyYgOnhMJrLHjSizvDx606xgviKjY9r/fAMqC/
mE/VZYS/Zwuu6EdzFeOAmwCO8YG30uRWOqOiIqlF5+SOHTqxYS0ChyCihMcCo1F1YFLqGOEQgWmu
FT7izMDdnILhAj6bWY/bbq91F25Bu0Wsu/xfOLbmkRpS8Rj9ajhVKyKApPH40yHOa4mjEoIrNK42
gNzwhpXu+v9T/PezTaYF5w9I1ZrwM8hEb1SV8OvcOVeVSiLkiqS9SGYWuVgkvJBwKZ2/XsqojRGe
6PsFpcU4K8TdaCKd1C74qJPs2SLeJe+sEjNXQ1GL6hRj7l3PR4km8p63nIfmAI7UlbYqEaxTuXj8
IdIh9E8Xah7qkHxOSlqNpV+GXnTrYbA2WJAilfxNc0zstTNHhmxrUa26EHjDs6qoY2860/Z0pVKI
AYKgpiHHbm9xaodw3k2INQPpily2UROLUwzVZ3VfQKq5nrRhub9Yq/ehOnjuZ1iG0CKw55/cDv+X
vwq0MuuVpXffRL+4UCQMp4xqcI0p69t5UtZTmmNH8R8NTStF8wqhFy60tyZPQxV7VHefjET2q8cn
8dOOeCwsFHfOjaSWcL3SYkHIr7+hOqbv6eFLHvdwvLkn+ZFtzFVZkv6biGpcVR/xd+N7UXjDcZGa
aiOo066mQDGiWvt5eL6SDQaUVRUGHX2aUxoDPOw8h7a4kWaZ17vMX0G5hhFQgr2ha9UkGNJGJUNc
G7+xoT/QbtufczixeDoGltK/S8B4JNVq9OlZsjkCQxdq22PlGNv/c14EsaLkTI9gh2sHKVBEtevz
s3WqGV6cdyv/PqsDGNwSJfSOeSBFbpp80/U2cK/MbZQuYBSWg4dCb5fwflXMYoL645T7B/aJzVGH
RY1Ju0pHnw0HQrqkRLTkseFyzvb7PQwKdCf+q5kFd9BK1dxeWJURCbL78PuAbYNQ+2pilS80gp6E
DeMWMOzcnwZUkXMCOVjVO71Bo6EzKa0xu5BOvoWbyqlvcWPDvtCmvG2yFeeq9MpnekdWXPgm4zfU
RLaVVZLDIMY8//o4xyW90PoKbUjqBS5b8YG/1fMs72RVlKLTgeYnczB0XMmubRhqgOhDrlWopJ1C
CZf9T1ow/X9P7WZ1/G6Z/C5h0dCUt/EYrt5hH9k8ONILKOI7uyNOmc2yhROUvWR6ZxzL7vi1WilH
9myoYcGINibX/tgi2pdVKxw777nD8t+QZJLf3ks5ygLA2nMpqWiHOwutgaJr6sUKRgZqNE1WDdpU
THh1O/ggwexlfUAE83W46hACD5wVy265QjC4VIfMz+q0eB91Tm1oPDCNb85apY/6zcjlESk/3mYY
FRFc3zHYFdT5EPYbX3J94HaDMmSaBi5u3Hlcxs1s+/a2R8/cr+/isvao1p17iPREprpmz7W0w6Jt
HBXXmTnY3IFrJtP1Y62v39ghRu9TgrDok9Hn/PUSFpQD6WH0/20926ukgMA8IbpT/8Cj0Npr0UMO
NjbsEf0N/H4UpvtKQCk+U+cbMkk1YKSikcC0JQXcCAK9fp4puWUziyvy/MFIQZ4HkhF5Eart2sWG
wDYf8F80lmuqu9sV4aGv0yIAwMdeBnFjRKPNPVabEXifYuAg9QsOrlFIntYLQ/twxQs3j9/qRu86
egnr3olK1dNQL0hojeRLmwr1EhojVJTLeZrgvNQo64atFj8Qd/xnAnJGjlIC+2wd5HsSxlx4mh9j
/Vg7VmMJJdEjYgV74REEWL7aZ2ugVmlTR0jbA4RtGOWUvTTJVe1Yg+FdmVQ6WF9RT1ApKNvA44He
vrmjifbwxV/Wmpb+M1Dnyy/zmpE4k4VHR6sKOSMLJwN403twNLNjVDrNyFn1SbgZEBDF3twq2FgR
smVJc6lbBapw03Ppvd4cWXOehh6UErpH1bWkZBn6K/GRErsPLf33QycayUGflExlk6Fsbaj3N1Am
5MSp3QyLmztVotWOHNuQunvFPTl3nqjdz2FS1MnGhyC61jnQsWycUTRSMVhyucgKmiRrZVD3CotQ
3TGb5VqLdJYV6u2LAE3Tgu2rO0BHoKjc9L/OS00vfNFccPvtnxZ8K5ll51pBRBU1e8tpIEa+pcEO
JE7V/liAU1HRdCO2xvFQSUqW/Dd3TpbdbZkppGF5eGhb13fkkOpRWadlIbE8bBNvrhxHCWpa/1n8
/svbdeiOImg9Us7PuCTwzTwGU0Yg3GLoMshv894RQ4LOZwXWVZRBDvWHeDKlLYM7iDdlItPuBOap
eCdjVP8th1mDLfp29azIO8oJrQE0qr3wMPLBIpfk46HTmZa6FO/MwHt8PqDQmDkCCCcTftzegJQH
1n+taNedSkCW7fJy3oyYkr7rjwUSnzqAN+f0dILPnQirVEx8MOr+B4cGoqdsPUpgfQWQfVr8Cn9B
mayip50ia5m6juPeposVKj7lZIcGSYm5nN1HjHCz2nK0wiQtEsRXMl+tlMLdX47D0gVBROxEWGWu
zfexzj+Vub/9TXcGRFbmwcxwj4HXu9dKHEKHfY26eyq7cBdRYtkYhDLUy/kXZ+GXFoyPEqwhJxM+
QCpH5dwtXNglWdOVq2d+h46S/RFNlQ7q53ZCQrAOX4oDgGCjKdD42pVNU4DrfBk2YilpB8ksJn8Y
BkkdbJRW1YvnikM52sYkxGR3Oexr5CJe3fa71JjX2RyJIcaLI+6p408M84gaZm5L9jgVNPWoGAnS
/AIGZtMARWvMUXb2O/wXufMxp42kRgm3NwYKW4LNSEO/4nk81KqvxCQCYB3y9O+BmnHbulgBOZd/
/zYAf78KAgfh1iplsKjffn/w6WPxip9J0LrlA+X4AVCvzUNlTSh/Zdtl/CZBy60fTXHmOywkGVwO
cVXUluAYCLReJ+bGZkmnxxWHk2vxOFOg8aTDgi9/L2YOtQQvMglOlLjIWFKcM2ceG1fyhS23OxVG
/39P+SsV3m38aCfZrLCaBzXafKTcZWCOeYNposN/3Nip4jbVccr37yG22Zfd6QCMMbI33EjkYVuw
YvWaYA2unE13vOHJQKOmG1fTtHW0wfzN9nWP9m1JmfGN5HKeH65wsjx81k/oWUDNrHteGmqMc+tY
y1kAK6KN1bGxkNTxRvr0v72GLbmUhJeiunCPNKoIhcD/iSwPgctk+fEx3l85kBulg4ii3/YzV0sh
XQPhDnB6EkvV4AzyGygFrOFZ1RznGvy26f8w1FNylsZsIQv74z1w08pwYGhFbhwo4WnAKcx1lcou
PW4ufTVLCOrrMqh13MwQoRKZ9Pok4ijAd28QipXHb4wlSI72xKTIhKn7/MbVf4sHMx2hz7aDXBQq
OEyOmtOFj6m/YnQ3hMTF5VDBEdVlC2WCTlDwICVOI3AdEvaZDDqKS4xQxRWVTpZVbJKu24VCoqDL
+i47eXdYd/giROJCnyu503aBWwFXh9Fou5xAVcsNozsAQCTWl2HMsPy3OtTaRhOCGysfWAUCHwii
YZFUx+0a6T2kXzdOc22MtlrX7c2r1rcnPuJsHgaiDUvxm67MzI1hmPqilI6Xkxn4dzXBaIjSXJeH
eSngjHkqdhngb+y150qSjGKit2GLCPaQvbuj7Kh5JpR8bM5qbMKA+9SzgNCUBHdqjLmc89xqtsTZ
hmFBu+fisO9dUnE2pjIlageu9ZpMrDicqUtJxwvGzzHlxewSIWozNVd37vrW+DTeDmsPJv/zm6m1
ZKKfZeVQwQ2L2fxELtZpd85/dC4s0OmGnEvEBb9PDympgeQrF7IBis7ysSMK1M5heWT9/P6af7Sq
WPk0Ls7AsbVAdXolNNnig8V06I8dzmS8BnUWzrU0luhOvtMsxwkCx55XegrUD2c44PKCr9/kcMYG
eKKazpQvnTwRIwDQ1AWkGFyioNZgtaoHSpp3fNwR7MPmTeGUGOgQPgrPBXYqwSOOOlK3sQGwtbWr
wgPK5OvFOdaVxbXw8p4OMdU6rhXov6r/TC2uZwMBdzZAjWeyflQrXQ9DHaDL5NXkeU0/7xdANcMN
lNZGlDE8g1DTOapFuYzBbdIMrVlqEEmPXQm2ubTI0N62qe7q1ckVfvijkf5hfin4TkpCScpgRGyL
N+yG4BGoQFnOubfkKdaEw8FPdqrY/zU2YmNXaYPOfhgM2rDE4wr1h2+M5XHEvp6tRP0nV6edHx9N
Z2yVRD4WgRgb6u+S36yvrTkUEmqjzGHIqtpOZBuB2L5z6U0gE+FDN/YV8KRnRHFkuPxN+Yu0EX/i
sHeZYfNOJDnvzlhnxI0letyHmBBnXXAskwXlQiMfYNmtGWBWdVsjf0uZfuQIYFK4Xk+ocCg5hwzC
8XwH81HPTT0W+RfZhX7CL8s91wDTu+cgSTFfhUGsAnncaf1elasftl891fCb57fFWteMkacLVbre
JY03Un89ljxWLVae9unlstLB1RYMzPxYWIQQgWdzmvn7OaWCpdxsLqipJczenP4AghCeKzMCDjeC
ehL4CT5WA306+7+ZOuHqNYlH4Q9JKV1bp+1xGFQLeWGqbSHnllXdc3Hu5Spn9e2P5V7/DBmYNzle
GkpN97bVI6VqdeosyJ6sv5kyfWUz2Iers/B098lb6M2b77VscIhtQWJjXvKB7aslW0fJac5qhCFC
bGc75S4gLrW1FvolkHGzp3EsyZW4cvPyEo7ccamCuVkXVm2ltyTmZ203btDXBODjb2vyE5O9UTTQ
5/rL7/JoySTrkMOLi+fqFojHxf4JLZeSBISsAPXTbNQAZu7Hi7wOQg/AOPEVAZWL0wryGXn61fYM
wWNRplyImvOLd4b0WfpawNeHzkE8qM/85mwZMk68T3t67HGGXsFvFJNr3xXwjpcr9msEDEEvHC1u
bNToAOpxQBhdaLVaj30esowl+ODW/99HLXKRnuZo2rYzqJxFtBlR4fM0XsNvDuEZNUT8mxYEViT9
zpgsaIg/WuMfF+tH+UrSqNqPDF6//ry/dfZ9xKPkQ2qhWAkyrIs+LRWad4tnbBNrAWr76b2OQc9Q
J3fqc18k/BQWPew2fLD5cwvbwgjYT67n986wrScGKTt/eaMQFpyPkJnkZUEy4bhY/F5HTyM4p5Pc
swfWl3OdPEFdlLQzntBb6tWr436/mEJ9qbYsajhP7p2eMSS/giKuKtIhYrtJSFBs3zrjezfonokm
O3KlP1xcVYknjo+JWXV93NWWlOafJeghvhIvhATPeMx06K3BBWwvpf2wzeCur+bsCJlQxML01epo
TpuFSpbCMTuFtsXjX4redm0jAkeFJQRATIpwE5JT5t0dlfVhIVDWMed1w6oC4cuI/RirXr5ZU/cl
CLsOiPSjwM70bjPqKLnYtTi01LoYeHLn1lyiFp9k9pDLK6IdHQvw7rhLRskIvhgXaZAv0/vQSMUn
A0k45Q0kKNUuVEq2mKvhVWDeYi1/VP84wuvuQIW4K428ahHyBms83xopG9tP6c3R4E+Le30hiU8d
Dmg+btXivWW9mzK7TL1irCD5K2zZ7Ip6R0lforsEN/EgfQCW6mg8lmSoEnUFoADJ84YKazvzTYos
BWj2ErxMxLha0ldFcPD9EQoVmxqbBEbtPaOth+A41xlQA5NcZzhyjDLZQujTFqTPbkih4rH8vRXa
tdDUZW44gVJ5kHJhsR8g/Z3+qQBu70cTF40Gf04PVeks+JtwVR6433TS3hDz8ssG25qMvI6YPduv
BjuDHbM2cawRv2qHCdz8sH2lexAORyfpRPtdmZJYhb0B5K1+Ow+fS/khBGq0ehgM+dZWygLJ8yVG
EsuYXMBsoOLMESl0+ITdavmF+4TO1nx3dLQFiqZrwCq+cjWNmteCS6bPnj59a0oH4OWBF2zpK4tM
NXtje5xaY5pUzkP5eqgQ4e3qVdFFsFQCSQ4wN17po3zoAjNnDJvTEKrERv3YhvDk4FkslcxsBKVl
wGDRGqdz9qRxS+7diuX22IpGg6HqRUGzSnsnf02xOK4T+a+6N9osB9nq+HrTdTDjSeHW+IHqhV7B
iT0tM6mjsCDZUXr3Eb0pFKsJc4914zQla4hTd364Gk3Xu8sF5ChO8sV9HVLP/P51b6vWrYjKM3qB
YWB6ANHaRqkmtc9EWCB4oot1zCtXp/buzvL8vdLMkgE7FnDaQ7lgXIbp7GEaE7aW7Cty4G48sqop
oSfaonvEUFVq34z5hGE+4/1m8/ZvkLnI26uXBpz+RJQuwovTSGNJS6qOvlyCpP9btE0j017TEB19
07hI1JBPjmsqmh2qjNFt1SjOiWethI7LjFGAdx1yEHGUxdy7h2Ld+k/QknAutiKERAOmVU8xNIp5
6hwBROAA1xnn9LCSREvKYiuB5Wztot0r9f+ytrn/WjF5MeEQ7dra3k6VVNqMTy6RDW5Y0/BuwWG7
kyWG2IcNSENNf/KjRpTuyK9WspSWPuyPxw8YxB5YMjJ+jhpmwroSsmxA/HB8mfUkUaXSnKRXHbjD
KGZhLwvjKm8szXKBxEHt8LDBHYlvxccELt2IN52VeAacva1YkxFAs3Hz67jz64AD/onZMdL0/AqC
wiSXXLttTN8yq0yIseJqWowK5z0tgAQr/xJ27M1J22/Xlc6zp+zP4oTVql/U480QBEw7A1dsw9v3
ARhRL00SoSSUqeTTYWjweu1HVpTEeRzG48zgIqM9jJ+KhizOjCujF/rfWa5rs7oL1tVfepv2Mi64
T0FkFn+IrGTWGH1qYYr++RdEFAIJeu8jXDpv3iRqODr+BCB67xcCNDVFdwRG/0+KqAZcZbaZpGDV
UBdmOBPd6xA3AfN8K+B6N3s+iHV2iZ+kWpca1u+qH4us8JeP7EVepw0Snp3UCyFQbDLlWq9S4hih
OOIWt+UecrNBw8Jqn6PB6QNsvdpKET3eSwQQwTQ8jC03oUzq3NIEcooSrJkTI+Q9AaInlStC92pA
JOPzF4jpmfmWHrQyG+xVtYmRK1Gr1TJzAikaz0GqxvL1Is8+p4tbkLz3dg/DHhyt1lmJSg5FWBHh
w32U2mypR2sFBW+hTQZYnD76a/ENy5oAdG2zfKwpdiVf+BbbO6I2UFAr5S5Esv7uSpLAkgMFu/wB
9KpdEQqjQAOtk0YilqhtaaIV6fVJ1YdJVRHVlYzLKDy6YNpKxcyDwvVgq9JjUHcuskjMJzr8NI0Q
hg7L3k1p6NftHxB/UFHqdB44edSBvby3j+AffEsuySBtytdhsZDaxfbK3cgofdKQ2T+vNjNOqOQC
oweVVGasD5WND9I3sV/My6LWEJY9UuOt3rMFsHfD2vTBg2Yv93QUqa1U1HA9WKXfFtT8pdWeRyjB
TIoqTw/+eB5bpqVn91kfRBFuccTn84cLhQf/2VURT+U2obIxcAqRr+owleZsslMFs5jDZp1jYmWS
x+cwUVEBuShHDcjhCvoUiswfpYG59wl8WCimBeAOUeFzVHbFqs3KPJim/TijWXWmEISi77AHC4RB
nhVBUq1ocPVmFg62U/cbRAMY3Q5BnpuNusHb+II0EHSBr3xZ52el3Z3jAwWUtVcDIDZCCUpgG7I9
/pACY8zMm7pqZfGBERaomTDbayNmKVnI/fJvpLNg2Zyy8ruJ7NBHY1sfI7KY7/Ryc7BsTj0nkDJx
yGHI5mlI+WTbTNYp0z+g8tWjTCdi3phcFinuifmwbkvis9CA0ZcQ1Pl7qevc44SLddWjQaJ61NX6
CICMCX+yhAvD2RU6DXvWr154w/1bg7IRdSjd1X8EdgIi1cWWZzoxHlborzuw74Xmx7gbjJ4Zk6zX
xMrAolKbaewFcfIfq/SWq658iJeyu+9YflpsdP2Sx7JB8WKi3E9KUCltoa8j2fk8yQA0IxPSI0Yn
BXaIZRN5vAXB/oJ1dy3dXyjiod3FWZRHhJsTbHT487A0YjxyWYyQ0dzVUfGZAuKpRjcti26qZeqv
9Ix1sSEoF90KdtYsc/boXLvut0E5PYj/aGDoocPFQURz8e9Pzk4c06Fkomiq4Kz7dQK7/5sb61ki
1kTOlw/kiWapXTBz+/H8kT4fUueu/ED7Idmoy4CYghjxY8U9Mwn7ctKNcnvM8F+EubfgTX4CnPrT
tYEBufOkeTvb2I/Gef9IGDeFLfwkXyruscNDJEQwBMen3dut3gNxRNtZsRPrQ6XWyXhbE9CuFbBD
uMrIGhfc8EJqMI4c8twSqghxUpXw7Aut8ObWAKoOsihcLzK920plejnNt7kaYa4h7ABf5sDWWm6H
Q3KlywzLKC2/2SDOCAtPhgLXvXeU3lozhgQTaHWZFk7X4t3QEh63cIsz0ITA8dtPJcdqifUZeKYq
Iil+rqWMuEXjB92I3KAmp6ueDlydlnLXA8P6R39Lz9T3OjR3Takf1HBRg1CUJ2gZUXifSp/Q5TYE
N6dGwD3LL/MYnXWx0oKDSIH8BOyfpeX4bw9y9vhWrKVkVYP5E3DXUflwiwk0OoO9q/x7rT9iHjHd
9PQgTjgHXH2TYWWd8JFW4wm4oAHHIUcdB8J+GjsHkDbxolpGiNw7x6s0nnp+e6wyhCDymbnKt4xE
LI5VY1R7IIqr+tDj2XvFI8fAeynvVfG3ot6S4dqjIdeyedg5gl//oXLv+7TjNv1LMjBFq3eRAXhy
pro8tQJV7DnBdY4YXu/2TUcVwTgdpcv5jUKqlaidzEkcUoESQ4A3NGTIDzBOfXK75rHCRZJc5fub
g9BAuJZubNsuvuni8X/9Cdq7xrCNzxKidmvFdnt72pfbauAe0iVKZuoD7qTmbuLdwTHuEOQ1UZU6
JIB9rK5Lwt5M/F+vPQe6zs1NykZBj2oB/GskVUVqk/OuJicoDO8GU3ru9BKUcC1Nvkb4LfhmMuWH
Aet6ATybK+RBypDKF/VPogTACvgUFFOw4QbHDs+sAW5Q3aKxxvSh7IS5hzvv0rdu49PsY3ObGpGo
p9k834TtfKxwMOa8dtjEAV1TbKv3dV9PUP1cw4tgYlrsRyEDxsyy4opwT7Cplar92JURl0srPrrF
ihG01ajq6VkqlFKLLRjzUfvDDGlnftYgrYWCuf2Lt93XmitAgAxHO7NHcFaomJDCKLEyPU0kjlYY
yh4eHqt9JZxJ7dpnQw6t9n2En+6+AzkbvhgE71qr0mvCfrLZNv+qA5Xw2popq6huzcGVQEehaqEH
Y4N2oGDSosZsjsxR/OUhKSMZiiwA0LHEEKEqQkEeFHj1MlSCAbAmRd4PsCykqYlXxm/i8xGns34H
rH7pGCIRAge3vGmGEvQpRIwcGjf0Xn55pb561LjitLxjxv1YTtdunAqgYQ4xpAJAX4w7wRBWL4K8
phQpcHiAmvQRDr8+1XmaoMf3Pm5t6TOxJi4NiDi5Z2fUj3EfI2/1UIYTW24N2XDuSWA1MKtzgEiE
RkhyY7RC67CfQMef9+3ea51BeDCtkL0jk+bkJraxgW+P5MkaXTfJTqgeynL9zlQRuq7t3I+Zz/tO
UnH2IztHKOGSLdy3bmhZvq///VZn3yAMzm3k4Ke/cojlimBmUjdxPlj0Vev0nl9lA0TZ4WBigpaV
xAySBr+y2H27R68Y9uSSduLlQX3Mq956ONgKYGc25hPzdyeClw9VAOPvbcOzrZGk15Mhx8lQcMEq
G4NumD5PnPkYsay4DgHS5YqSAVn/Mye0S5zfha/g4vBM3E1aDHbBsDz2vD+4/WyyVpPXbmPA6MPv
vHU1hJbG2XGl4Iipt160+P3UE2TSx+S+IAdq/Avb0k3WV0VyBzAaxgvlsd75wkvR8fHhMdk8hNfd
Xv0EI83WA5uHq+GBmI/cG1utJQSGYx+QmMiZF6h48/nF8++jwDwWBnOjOm1phf3XgL9dVZ12cil6
S4t9VhF7T7nD93L5ApqtSSKyi+1TiErBckLxvPLrsINkpSFnJtM54dJmW6PM4GCzRIc0yEGpu2jB
i1f0E87W3yerMUsCmyznqPEpX6bdvIe07WFkc0p46fPfdklJ+mHX2ob6iS8BOIo1sSx63odFr+3S
YHKuz/Z0yxkk1qSMYeHEH6h8qXcBQI6jDn3E/5iXD6hg4FaWz1SbPQc7k5rXDabxwTHMinfM7XJD
2yWjIi1JmJrZoqCslS1ZXwGXfhyU+w7V/HIi+zI97GMDLa3L4pPV38ffF+OLn60Xhl0uLE+yNULk
f3ooFxLSHZE5QGROdGeay7VcWU2rh9h8ISkPFvKksRKKl9tW5/JkIKUZ+AXDh1RfkqnWrh2+jO5g
Iw4ReVM5mIuSQIZTe5bcqUA13HFvVdfeJah3dbgsNx/7Y8pYCFiKaNZEtEw5JRYizUWrA1HKGLu1
HjFthLR1TBU88bhUwTg7KRIZFEhvt5Vy5gf0RGhpSZIxsOrmRnXWBXQ04Yfw5OfwZCE7hy3cOuyT
NrslIQ7tUTFjXwlTz//yW1S7BXtOLnQ5tG4ymCHfbjDXZxxzy1+r+74oCq5A5hYsdrvvv8RkxS8P
eBxm4qq4rR/1NwZNRzQNP/jew7C8+zscqINQwgKJY4KHCRFTX4McgqMuz9wGWjDqtk04VbPnODYQ
pSuQDHM5sfoZNwZxggpsiWjvDwvkoXllGzFRUqlh1h4PFQlHa++bvzBj9eyy9IEWVqm1xRXeRPx5
pQm+mBr8HSnDmQuBLFDmsQyg+pBRAsijZzibUUNdcVqlk7vF5vmNl3/wFHQYSmL58Iu9DS5Xt4pb
a0X7q4K0PRg6f9+I1KHMcfHwP5DWtSnIkbTplGlnIO1Ho/Kzp/S8ZLOBpT8xV/QU/pm6K5hSxMX6
I9y4rehrxz3clyGCZ6AsxSb/liGsdbUIc7OdCBBVc5bN05DzFB2kjROPoJbTsC1CGCzwRobooe78
Oe2UQEP+dACXg1WxT0s74lv7s/iOsrOsaCfZ3dqSf29wmqgUh0XyIog8YB4lJpEeMOK4I08WTcDH
P1W0N93HJLC3MA6tqXkzu/xjzNETL9YfxIRCEo3NbVOBJoyskt8InCV745GkPDwSXY1zfwFri1sy
jTH0Z0ORLlrykTdvD8c2NvUpgD84dteKfoK0SRQe1OVc5E6Vy9nOhVB5ZLYBgfoqOe0+t9aMR6uq
w+CvaVkbOWzdGt9GeU+y7ND9PosB59HvkjzwESoeOYNzngpbg2fg7tPI7udR/0UHae9sgSnsZBH2
CgPmt6C2nOOK/TMLPGGAPihXEnErQw+eqPmZz5qM/64G5zb5DIsfL/zfKt++1k0knL9Xb4/K5etZ
0mZAEkluCy3rb7ycyunLHW5o0M8PsljSe7gzwPYFv79ZiNuiLqBl8fdfb0I7rdUoLNnfzwekZbZF
Rs2+Ia0x/0GmH16IffFrqkL1+FWNEF3VoUFZNF6ttv1ffpb2CYcZmj1+JXhInZruHGJgud4q0dk9
qIIiNVDoFZDRcl0nm4AGVDWUB0FYz4rT1gs4/6eUrd5KijuYr9st12gVLNWlH8ln0OQyjE3TBLOx
tK5x7G5UiL+6uXCZK/wKIFxIRHFjfNU1qUpCYNJKLvBfJDVtRqcej++WBFMkkLXz3SKE+hFCq5SJ
rUg/vWZlR/yxIdvRYRL1RK8QcgZsXDR+3dt6frkmzivIRRl2yEGSGSDjq3w4MYbiZ/yoj7xGitQm
POAemZxmT0untM+92DFUrgr4XAga608lNoAYvzzeMXmLv4TbDQsswSLnvO5Ghm5thehsBOn5YpjB
pviG6ztBRwnaNDwbD9w3E9j11hpWjJZnj9i1zLF6wYORltn5EiOo5wGB/EElfMpgh6C9AzDPUkAZ
8PjMalsTKur+6Lrme+lL/pKX11Ljz319cK6aHYStiOE6kGiE8PgT4To0oMc0xSRjubKj9s9YhGub
THgVgk+jkAbGbdGKxlgDkahhvM5Aei1v87Y3SpwzycGLTgPsVzgGeui3ToehDaAqASLtCB8RB+hl
mVzpznY0Mt8La8g+AwR5aJsRzBfoM5krcNig2BtXh59Dq7CCdXOkcMzSTV8VaVpZ7StAX4HKz3Cl
ZpcLEVsaTluH+pIbbKoBFmkPhJ9eC6WDICgwKth3PlyugzQ7az85iepF97VkwvEt19i3b+jzyvda
eTiwMIA1dOzXD5JFcrfT37T+FCW94h3tb/8eE6kKRU8ih3D0c9+jadecL/bGwiyzIMWAHDIXTxBg
tZ5fdrLfQY/GI5EEydxrZopH5s3ApnVOdbgEK4vLtFlbnxoOrgBwW+kskq0voca5kp4sx6JcYBog
KHkjBKPuNazGJDZduIJmBWu9EprUpGWZFP1mhGxP9Dn3501TJ70wJ8mBJBjdQDRsCfOwb+J2uVGX
BuklYCR970fP+choE51uxaz6hbjk8igAdLLS3eY3KJhWSOLwD68ep84E7Hmr5si/ZnK+9lD+lLnn
bT2vxSJF5jGsItlyWQUFxlQOBCOs1iw90+vIvfOKqdsh8YQYAYPOJ8Pnhdde97VNu1pa1PbByudj
+RY9iacABX4SNbR41gV+vYXEJZzzTlEPF9iQmPD2X66ZCT/WixhOsY5u6k/Xm+juyGss9m85Sr6o
kZUsG0G23fn/F9vjLotKOhibhxnwPunHsqDTEPUGR6vOydRe1h6ASETzJwjpFnPh4WNazpdQ4mBE
JsD5/3z1VFIb7xp5phZsWABACHQednRSjjvB3Ua6mIg68VFrIcz2rJFJZfNTOR/DdYCdn7qm5trW
aB7DqDzqZxWSZJ8wfRUUIykThO7d2tIXFPuVVGpESJbk2u2kd9cNJ0gVGcAdR6pRh6QU0xjW5ztY
NM65QG08Yy8mxYsMik71HgYFsGbPBwaDFaPa9RYpfb6qp8SVkMCbNiRinTriJ83gImGDtLSMm3Hl
ECRC5uLHznQz7wK3Os/cR7wUDt02YEypdxKn4mg++NiO9JRmeDU4rNkKYZWIZ/RTtOoeVshM/ec0
aniHSG8mXjvup4xAyGjHTsuui+wFSC8KraKp8bRhcDLXytLJ+8Pgt6EADh/XuNeCkzauQeDfPiM0
5B6p15HehGD8EfG8X4YTs4djCj75Y0asKvwEsyWbOJwuRdd6nSnq2N2nJCwpEtkvm6I70leL8tm3
1L0nWJjb5CoLR6crHIEJ5d9v0bhit8c3DyN6vuJhV2DNyPB/K5eir6hoxRJCfOHwZlqeXdL8p+pl
ZUeS7RwDJkMpMu89aAXJqW/kunzIJYmbWeOScx8FvCLemkQ3qmzRA93My/n2Zc+9ppPjOQpIHi6f
6RfX2F2hTbnXMR4OTMOZexI3nbN2Z4cIJ58rkniP2b1sMwEC+atmfNm2LnWG4XCYZRDfR+ryPtsG
XALDwJmD8drLC4j4zCQNLcuycEJ2HlCH1Av1hkdmYE7MzJBwXOTy3qsLtlo3RH4JrR3blkqY1Dam
DjWvBjm9o926OirevYdCCdngVE1ALtk8q8WIbR0R0fcBgVStHqaEnIe0UVTiA5iFTgAVQta/qqyD
o2kYZa9RgXngeHUoxuvyNPkn4MEr6jghHgkwdgFXN0/+wYMdD0JOxFmKvHKxgm6RANe3n9cbChlF
tJvpDH9I9Q41MFz7XLqsszg46dSEkEyZbO1EbTyt3zdluV4Y+Tjb4SGoAS9jOCvOdp2OANVAa0qs
Yr1UFlTKL1flUCgQjOy8ikhGQxQzNDjHkKjQ+3dJLRRthiJmC4CExpEN9OaSaJm8spBd8/Sd/h0b
HDnad/VZi3W1iQYTOCgOYCm4C4vvgzvSU1wSZafDsnbjTgFOgQ5+vkX1zL9H97KvHPE8/DpOEgBs
Ny4l6tdDjF4HJsn3f0m31g2z3QE8VgUnwKDucp9hzrZLQhfQTaO+lODsL8Vpsen0XuVWrpbUZFxo
fo3QBVq7UfU/HW3C9Vri6Wldb7PYcf3wppiRzeGvT1/mRb8FOQnR5gnSUL7ILzWJJel3ynCNN1ws
5vjUKnKyClTSXLKc61zTcCQ9uoL5/6VlhMMmqx+dGzGu2xI1To5UXo35eBxd3qbAxPE6lyBLpO6Q
hgwkyIXjqCBp/yegXyVpZ2xMZHFoM1lgOWRQELw2BP9NPOEaoZ2Tf/Saqk/6XqdvJjZhodp3hzuE
MzYSKadYd6GcbrR6x4NxpDaPUPosLkM+jPHxzAI6+D6cjrVwi0HId7OE+HDuvOnmZ2J92FNUVAjr
jhW9JP9bBcOqjSNFYGJtuoLZImPBySP59NqCgKJMfVzlkVM1ACGW8o79QqfdkLwE1aRZoC+l3lCZ
ZWislNPJmbe1BY2/myRSS9Bl4UAfB4vFjeOwNI3DYWUXJpreCrjbtCcJvk1T15UjDi+HHW8oGm99
SKgIXIiIbZmTn77JanH9ENpaG+xH+ayGGVTB3sr9lkDaW79LlZzp1xGzmEcJ+jLf6sz1/CxTWfjE
iU6IqmVYrsn7dIeS6uSR4pk28stfvrgvv/fJ/XDnShHTmIsl/WxcaONBATQd2zte7zZvrITbAyGE
ZBlvmlZkCJfep5sHBrv9f4a36uojzfOLuxK1u3EdgXftZkXpFs4urnWSFZJVMut8Lu5d5jF65ZTz
Pq5shWwtD8wVi1oIt8tx1QeS5G8TY+uRafehmt2KiyDPVSEgh6U+0kidb57OVg/QLH9z+4B6Tjdz
RhYS/GC3RgreRq1s+vxcFDEgsDH0/WEc90k9ePCE+2Yd3rkZC8lGo4y0Nm+Kg4QhiRZdlCF7VmG6
LT7sLh4hkbARVp3GFsItEgap7lynKS0GazfhrUYwiDuCceIQa9GfXikTF40OhrXhlAvdSxM9QKaf
vCTc2ZgHDWwvYtX8Bi/sSncop98zUOlfjTVSuxwQlHtW6fkl0IcAtaT+G+PTxRh+PYEA+tvEMovu
KAVcgAgYxe90OxZtzuTdOAEnh7juAAfOkWdZVhgz8NILml1+BWz1X7i2pfZgCAmASynAHxjtlJgF
VxsbLmtUyJeQ10bytTNmIlUWxvRmjaEi4YfoPr5u+SfnWrPOOyzgyOsi2c0okA3rV7tHBrr8KTOx
kAFSeHAVXYYFN0U5p1+Vs6WJk9MU4WFynZ5QhbBMCi2XlZJlwSgi/HuzsTawXDAXPRK4ksP8I/4I
FG0i3u58p+ADrSluD2IvyJ21rsgP+g97r135vsFFLZWVmSfU9LnTN98fiqhTyXWuq3WxS47dLZwk
UoDkBtifp7Kz/LT9umLOJW5PxmERON9c916gZ/9VuHsa6u+o4886jg8NCt96BQ3+S+PMBP0LJW35
e9r6KfPaqUIWS7yZuxPgK0Qd7GaZFAsmcm5heJyzX39q3/BtAnQ9YPxG/a5RWA/crIeNiPY6Jo4v
NEleURcDotZ3Ini8g4wRPX7Y0LhkASRGY6pRWAJR3wkP3Czch9QfTQ/XAHC1rU14kBTVe7x3sMIq
xBZ/7S1jcHrzd5A3FfPGOpFEvoYaj98sSPaT1l9XTIM91IFwv4Q+vKyJcEUT0OKOxzBfSyAUKryg
97RP8Hdw6RT8Y7hE08chO+nBIXdKWobMFUZACQKGv4UKryKIvRTLh2q3hxSMZmroFaD+HaKhHMRd
bJSU4sCsrW9NHMID8yfqusIZ1VOxWqlnA/uBE9C1vReX0ZtaOKq6zA9L/YIl8vQqhOWMBfx7ErQz
Qu/ooKVNDQjD9M4xQOYdm3Pf/XHU5P9v8kMusO3xa8ekmRU4ATf+P+DS+JWQWJeppCuT5M6TX7ti
9t4w4HbU/WZFI6TzxRtnzMHcGdnbpnPzfi4GEvnM+RgTWtr5XyHqCpaR46gUKUssYZD5Lrj5CNye
Lle1m0F0HwYUDsTurtorjnoruyc5RIZ5ciyAjfeteANOUIf59kOmjW+myXdlYa+lRqINi+k1yL6m
iOtlEuYRhEyMd/TEH0sgGQph4lIzMYlqdxatCSpUNSPaziDc9O0Ix5z4lkWvKvcPB1I/pwVpmWfD
Oz8FXkv80d7MOch1O/evstcKI39tUfM4i5hTqlJUADCGBdk5U1ms3odX4F0wYxlcXgFy3+FDr1Mm
cW7uqBMWhJZHKytA5dw9yrI9WUUTOUBFLMB/9tyATXYohtAMoer7/EyWV7lKneLAeUrxDwrs5Jqv
9X8SKkANMvhdnmak5OUGxaHqrlRWI9eFvfK9+Fi3nhrzMUz98TSlnW18D3EOD/LU+zM7pLuXgjDC
og0S6q7IJwgIIJn09NoxLIq0E2cRmKxKIMA/N5+olNxj4Qim1g01IZurdqTpbSL6c4jO2NSQ38kl
hkqISRHI4Czz8FP+Mu+rYMwbgRUx9ZrcH9rovJ8/Rc2kpcR/s/PTB6PYj1l+80qRa4a1pW9FSOmz
lECo+4kzpfLG0ZatND98zKzhArJEtQit2lpcYcm6gnDUQyJ0L/ODPZJdDvtPOPvs/IkONOwlK953
Ium9Eo9YtcJjdiMlmCLrhapfuLU1KLH2Lb1xAyi4KtzQ/DB4QL20Zx0WhqZzi7zh87sxZL14QuJV
PDGSrO2V/Q0ixwHvsA+vhmwJB3VXAKmVU1BpRiQy8ihSRezeKpNS9C2lp7ooDhuWrLK5sWOwyYto
x8N8Lg6YCUwBnBrOQTenAa18dNzSl3wQgGDWH0g389jMmjhbgo658NGXD9BJtqaZJ44XxiZbw6ti
2SHB9n6pg6NBzsRB8Ap6vpkzz36WyZV4//MJk+EOz/sbknGhAaE2KDxNFjanOEhh4/ecSbUZntwb
SxSEqueqK4THGFd1VxgVsbMijQJUGffCZVCeoecfVzKU8Q3jEB3MTO3bc2hBg1JM3EaMEVm9Hi22
tbV64/HmbPTtxpcq54wIUpHchDuw8EN1fApyqbxwDUYMCqgpOmYSLfFg2R3nGNlVr6CRPJiaYWW/
6g7YEMFKN06a1HtcP193w6zGA0fhzl9cmiLEVA3LY0PzvqeiyUQXJOAiXnb+uaZktd1TMmwkvL2y
7eQ43tjjaaGiI3dmwglDGz2SYfhFvUr+PbMDwPjko0deNBaWDXYwz8PMPtsmCt2xWt6vduDDcBJm
cNmMgURaU/a9u2n5QwsNUmpy4ngghsFi9kvmJyhafezgC8KSgyXwEAzQFtjcrlOtBBuew2OkyECu
iAstBaoelu4F8I7Ci2OQj6JvjQWGnSWjrIWfd9EIlwu0jMD/z6wSiBYeXsfIEjfhL9umst7vJc8m
hi04lNZ7YCPYNTiIEhgcc1ObBIeBtCOUIaGOuwGzahkJQkTYDkuobfPIkWkkL0FigpLweEaCfUd/
ymUtYwFn+pONglgDkH/aB7+LUquH7u8iSupGbk3MqLz75Fnh8bOMAicMIV/oedMCQZhoEsXeZnyH
lBkezEmd3qMrlUkXV6gzDi+iC4c2tDnv8R7YfBqEIRTcEXx4xeLeHoo6gpHcZa8PwxbWE/Azn51l
IQ2e2UDvMBNzkawnqSTnlzK3rlR6O3k2pOeMpnDa017+G1zgXw1PGKcjhTyysKZ0gtnbTy+mPVve
jCCelT+pUXJPXwgy2wo9kMbGF37fR72o7GZ//fFlJGoX8kESTPBqYCjfZhtOHPFIwDyOD3Z6KkXQ
ts/C6/12/KrIKtTZjdLj8UZxWIhlkZ2AaTR6JC8A6WDZHHsvGKz0GknCLMQEWSrXG36zxsWL/Jpm
AUvXs/T+/Cwnr6O7Sh8n9wS5bUVz6wqIf7+f8Hj9uu9LNOCWCGkc8scOX0oBW+zIfbjHZRvhXrdB
vUnJ1zVN1CBFWEwXfRIDB2CcJUFxzIpYP14YKmce2Y9M04830PA2Lz/juNQAo3ZiMlwf5Af/JvxL
p4xkoBVTFJ8VhivkmrtYA59mXWI9p6UikREDG+/Kpmk75pmfnKAaauaLT8SP2PCtVylmpZ0R0koA
ZA2NFMJCAPbLBAKK52iRjsB1K98T1X1UxZWt907cRyrgWWaEzFemZ7KJCcPo2CKL+++hQVkqE0IP
pEozubMElbzSruMbXYTHTnU03h+wWh5+0NB6MSpTvfSSMGLI1PV3CL9aG4q4vxqcS9c8mYH1oY2W
zYWivW1uxjEGq2CM+pQyMtlqacuQAQcco+qLDmX7jEkeXJsc3ph5KYmxt67AJurYzMFXs07I+Woa
FWSPVpM43XsFqOU1Gm1fvhdYJ7qsbJi9CZpzbGBGEtf8TDnRQIIDEeX9N/RJwHwx+ZaXe/VMw29F
Y6eN5xMEvyTm0fSFQDOiU3C8B0/0PFWARc2E9r7ERhLB9nsrtUBAV12tHNflSgahZI8dp1gWOpyB
ozXv9CRaIycld3Lf7gQgHB8StLMV/q6f3bFaoQsPx9wU3l4eLoXfbcFJO08/bwaRnCu85v1OAVh0
Hm4gTNEDUjENEWAXnsRrcGXsqMLod+oj9ky/lnSZefCtmKdx0Mdudz9uOznFgbVU/hKEtKzgo0TP
nAeN1X/yvjgKqA5KkRpg1YdxbxPRn6bmM8iTLdgJcvPGX982OzC9Eas30Djgr8KWPb6oNfJInJx6
qP/Info2xOXYrlTtPJLd5ft8jtMuFLuUmsHaDQo7egHl7pYvD8aaqrMI3BEQfeDNBceH4aErSGnk
h2sIN8Tuka+t7VxiPZz04Io3fDCHpo+INNKNGmxk6tVDFML+ogvX52LL5FBcLNvA7/YvzjcoKbHf
q7YToeiqyDUj6e/jxCdnHEn37+8AfI88Fx7TO//o2Bj8niWGUNHTd51z2OzNaitAb4HSGtvbnSPN
3sQX6Sa6+yhuxKhKxHn4wWm0LezLZyTtR06cB18qqhMnLt/a8XV/XYaYjWfI3oeUh/0lPAN/ZgSC
RYhbgoDBPPyPMqbr48cqVN4sOkZSS29b7+MIvMJ98eg8jx+RMNXvfICRopqJqSYTNHqhVrjEzZ4p
h7Oqn/krUVF+PLOlUC0QQd5LfJtOna+QhWtp1uuswM6iF81s7L9d+Z4gZDj7fX7sTsD4ieKH0Qxk
gpBkRDQOB+Jq9v+oU5s2Kg5JD6sEUfWn1jdctXpRuvo4TaEPMyReC+kyxfnxBIOxG0dDBJ3YELRP
mNCC6A/umgBxEu96T6y776LV/D6kIVGu6fbS5+HK7mcaGKDZ/xpLCgTWf5s/qx9Mhnpiw7NnP6RU
y1GaaxlA8MI/wpNgQOW8BuvEOAzQ0EqJ0pc0sbHW+8XxE13MWfn7T48h+WLbkTP7LlXxCgPKORpY
4Yr0a1PO9NJyeSq52j/HhgJ9senjRmZ9lW9HYnWCv735n6cS4YgMjb9vN+84nLQBpTS7SuDSnmKD
XheW9EZboc/q1OxP8RZi2P69cMtflDCWe2hV3+fbOWnvpj84o0j/sx5NlAu9d4XQIsOsufKdY05I
afYJEaLGvHp89u3uxrhwQc84Uat0NwxRNKDXJ3s6MT1IZ/w1TDXWDxktf+VrNG5W3sisDiNkeR5O
lloQo+4fvyOPgdi3yKoyHKO7EHoBMi6HN0jiLH6fa4ZqRftd1lM0lK2kjl38sWy3z93autEdZaTP
jKC+eGXA26veAUBx7+HUELljW6Gqc15r3B5cnEEsBIr5eEBwff81LzApA2g2gJqGFkHm900Y5z4L
aA+jMnHP+enJ4nm/fDnij0U2W0tVnfoJFtSnzyrXY1sdYUaed2nDeMYDcJ3zB5u9x2Ghsuxq/4UT
i963Cyd7o1LPNkbvERcIECwT0rf3BfcLqugYgcXEdC8lNPno8TB2y4iU/uRQ9ANEFe2GLFmEbkRM
848ytI99dSAdpvGA9jsj2w5IE27wmAbE6CNOsIetzpyPd/lIoFFdXVW24llU9dlHo30sU2MyLHz6
TpzDNKrDcPbZt5SzR67vURo26ZG4BpERGHzyO8OqTb6TNRLwk5FLmEJro2BN7m/WY1CxF5JKtd9k
+OSxtk75DHhhHn2sHEuLAlV4ozALANVWsELCBJDEyw4mb35/jdFtU7i63Q60CbAiI0RJVshd17iA
JveHO4EMWjnrE9hoh0FBnJT0TnuhonNPiDaq/ib1buqgJcndlj6dY1Gq+diQ9/MoXcKASdgXyYv5
ChxVU92fml5bfDyfS7whrgc8uF4WbqiF9CEBlj9nnEl41GUHpxUSF8u/gquPbUL02pPuxiJxqiEa
iYbf2uIe329NG9VKu24tNll7KSwyyQeTwpllUZQhX7nIi3w34+njWn9mVI+prLuoHMFvyjUOBUh1
+9jVV0Jrw5kLOdu7nIV/oatQw/0s86v6AKfXibgLnEDy0Sbo8MjmM+Eeq/isRntoGSHNUCyY2iJp
1jLqV17MM873L103PuQeTYfdkKAeRGYjnijL7AjOcUgjt8ZBXlRQZZK7mpI5A39e3KHQtjvzkpO7
JCiSaNoGE7B8ZhtvU5i9sw1GcXGPkmFlNjac/xzZVBCCeFBmjXGmrnv+QnYkg77BCy9Uxxyfh6Ag
t9w6Jpsa5y6O5THcrCvtw9Z3Q5oWNWWPn4BaQ7zAqBOyyhdwtAZmrq7qdEXP5KVfWuC5pjAgT1P8
2lcqcx/A+DDyWR6h5wZRVoHAnJEq7qxK5v1Db+nDhNQE4NXnDqw7bLaI/qAtdC7KDDLEbDJykMPP
R9t0VKDA/N7Ifq8vaEmbyqRmnDfYx1UmaCn2aUkZrt5Qd3LpjM16tRJUTSf//aihbcCm8ANJ2SlQ
rh1OchmI5uF/bQcuM8WrXTVjfE5AvmaODYZls4RxlxEzqVR3grqVpfE2RG1vSY6sReo4/FeonXCH
L4AM8ql7Q3Va++YV2ciBmEhbx2RsN4YR09euK+GE0ljfOKXI/JSMwnFJ9lMmWhyz0aTxT4q4Acqa
nB6My/Yn84O2T8ZfYtR2RhTfALuuKXwqkG//CxdwlKizLGiX951cMzNwEK1BTf4m2jb71+h+ikr4
LlG99sO7HVco+J3zcDUHKJV/AaAETOIXz4z24do39b/4OhCugbr3kbA2U5s+k51bcb9svuDbBRFv
F5K7jT5E8xliilOmXELvR1/KblOnDu0LP7LtsVaHq4QkPPLi1TXd956Km715c+8pvx8jLrWYCr9E
I85INh00I7/O7kWEmQLcYVe56k63tUxziHF1HD7b39ArLOBXD8ah7zo46nqb7CBfZ72rL+5hiZB5
Lk3cpFw5tvDl/5i362mhDgXBTFIFMi9xokQITAaKeJ5rlKHmwZ8EFs/Jnv6Hbrb9S7DSlwix52+R
+Q9djtwgl24BuVOYBn8DfESJ3gOYXOZdsOt1dLqRRZQsBRSiGupvC+3DEBr7spMV0oT1zXWk5BdS
31k6V9n8iefIrcq+266/7CuUbWVcbYhtKjrcZ92osc1WPNa3ZpjndbnOtmbUV4HGabFKvpreTJhK
DfFdb4stQEuywnwhcmZqdval8DyxaqnNfXvh6ZGkbRZcYiJd2F+f6oMfIzfSWNWp355RgRA7d3Ms
cgmdfu0FgSpBABWM3RyTLaOGoQ41eYHApFYsKJJ7FMlBvjKZO9tpbj+CqGJOo7Ra7TKZAt7iqPy2
J+y3meGtASHhRUhFfXw3y2CMUiTu4apw8xMOraftcyYDb/WGt0waDcEEt+i6n81O60X/0UU6sAv8
C3OOH0ZjF4w2/+ZmIZUwBsudf3X6ANK5DSEpDjNlOcU7SJB3H8xtigCTnZ5krT8DohnV/icMjH8F
vh6EgYTjDCqIucpNNsEVnudbmqlYIUwdCJ06SgtqfuxSdypXEf09VLn2rzXEQF8LGrOYAGsobsg5
Iswl5uMtqgxuKOXG4bMBaUxMTBtyczEHQgVZlWMd70NElDgTNQA3pt3NsH5PSANBPqd2DS5Ac4q2
zGTZBbdsCr62FFxWadjZKeTIyh4jESlFv8RNFu5696np4f0N9XgyJQssMqC+8bLIubRtdVpBmhz8
R4pJs+5GE63WwED4MAXQ2TTR6O+9FdNmyu/tHOoaYtXPemOxxCzB902oEIQzbJWKApJJIrhlxeOJ
X1UgPQtqcZJdjRKqHnvflWTj3J7I40nTARVVc7RNYJgR4L5107axW9l8VeGx9qD9BA2q4Vhwp8y9
tKt+Yy/2pj1Ld/WxRMvaMzHF1ssYPzOFek1oBttYtBYD71SgqEjZxzHZqg6J9ajDIhDbhmR47jPA
yt73+GCkbVBCB4ROr/5tCjlgXTuof0ycNkF6M92XqUK5a+Caf8KJ2AksmIBCAAgAQ8MksGuMbqah
jVSgJ05uI98EaM3PLP8oL1c0ow+b1CvQcfDXSa14DOd2QvxHKFR7r6FBoIMyt9nBhYpGzOe7lUNK
tWQrEbDrxm1l7nX/ea5ZslTSXOWMAi4TeNonuIVhJ2PsxQna7rn/JPexr0kJ6yvkrOsNZcvbZW0P
nSjjJW2uock1GDCaeB3GqLIj4OPNyuuLhLPLWuXyz6x0jtVCSXnoflv7SN5PgG5/aAXi/5rXZL+g
yvTDxXdaTz/rGD5Y2aYsx7a9l/1oJIqWsrL1U+ClWsPMMPvSFqnfUZQ9ov9H/ti9uDUziQk0tbg1
qeIl4XlTJT+ycI48ZXJ/mcQX6yIBj8XYjcnNcwFwsAKvX+p1VAvP/xXN/PA7lB705HKoK17dBoDC
/UsXVOQV3Lt84Ac6E5WPKPinqk0WZxpbT9PbCHgmSwrRnvGurkyfp3MPQoqgHTwSuPZe5SJ1S00V
KkibZ0ad9kf2/7OVCxqtHI0Vb+1ggkr+Vy5QYosmAZE8lCP8G+xJSrbmbl2Pipl0RdgF9u9EnObI
JLm4eiJwigPW17mH3h8ABi39XaB0z/TSPKkS2keOmRevT8CUvOKzqUdDxqEA3vCvxhleeQOnvk86
sWUBADNXxc7/hVFNVYPdZCUPMAFP7r9tYOGTuH5YVbqqzELwkJQOzKHZbjEvT7xNp0Ig6c+Taw53
kzmaTxqjO8SNEH1NUU7/MEwBWOuMgimuydj+Qmpa+3dQlG35QXFwJb3MIomb2EAJcFbPU0SzrGHG
WIqghA8EXk8qkN3vqrzUZvbZZ5N0FLo7jhHEHNy4dexZEVYy3d9xXOD1Xb2/3Hg0Pnnw3iHp3Xow
SdTBr3puc1WCmbRM8FR9V4QnCiDvUiKBDqKxWA530RynzA5t20lgk0ABq1tl2g830NpbPQiSpUrh
+xmljEwuCGYhPTYROef9RNrXlQOxWVJD7MiAViqcwmLmbLmaMwyIVXd7fKHB2KneDW/NwQrUIYKX
eAkLl1wh3rrWCYU5rfUrd8NM0YxUQw16k//8HrtpzQJ208KliVSd1IKgaLacojMkw+6oNWbEOVdX
1EQYobeIh/z7+EvBsSkrdTZ84KiDv47WY3lcpdEnpbk4OpRYFK201t2iR3lyUSTEDt/xwvG1Wj8A
7TGrJuaq8PLHGA0cYUnpBjJVS7NutDVO7vlKfp8p4Gh7VHiMTSObyYgaptdLaslgnWBW3ugZU0Fc
3j/OysXc5SHI449Wcc1MqYvR1L49qHcvn8qxEDSnW56pkPWO2/RTgIyugnIu+NOUr5EtoVVgo086
PL75NU3plzZfg9I7S15+Qnj9nnwFEPmAkq5F0rSCRIyfnO2NdWN2aYwy6zesl3gMJxyS41l3psJn
rFYzWeC/0tQXpUDIRTJxuRzyL8N1fIup9aiwSk8lK4UfWVg9NxnG6d89aR0oC0uLR+ZDEOLCgaS3
XIvNWq57EG3UrUO6Fo5E85KCOddHxZRHLSFQ8/sGRi+X4DJOSCLFvY9OjQjBW0KnVyjlTqQr9G9W
/cBoDcNBua5/Unh7iDucHxfN7+3lP/Wr0DvWaiQAnJ2BDai+jSlcLZK3/QQ63ouT8VgzkujnEI5m
lUgINTbbcsX0aZmPA44KCZzPN8Punoj5cYVwxz49Xd2JEHAuMk5rD2KDYeseqW8Cn3KZMWpPrUdu
DE8MUQYumiWVXoeVdNu12Ekmi5fy8LGhK8PnlXN2Bc6mpE32U92/OAxKEeojh6Py0HzLoyh4aPk5
REUvNEzTjwSjmG12/7ZVpbXpa0XWm7LWz6ZOdFSncEnHOPH6YJR5t7UNebxp4wh80EStRP9Hmpr5
z9Ljf/FaVDn4naZLTPm+JXFIFWzyHD76ltIgMx/JZQk2EzPhc+prw+SquhMPXBoyAHLGpIW5eRYe
huZbPYFyevf+8ptL8PkKo3pTkjI12OzmRVVnusexUUv+FqCMXlhay8abql/hPLvsH8PoIn8Q7qoP
V358Ut5AH7sWHj+lBVCeXkCebR8DuuAkGhVOsOUsy9eVPK+b9borowAzBSr8gUClUFuWbXTCaKaj
Zz4szs+SeCPOWC1qLrsyg72W2k7+rocHh5hhZyFOtWvOP8jkZ2IWB2/epvB6p/Gk+p/wBZE4Eij3
9ybmjsbGNMzkyVXio1xYCi5rgDRkGy9LOdiz/zCeU3bz8P4vd2i9MgBXtZdfFez7VZ6FfmCngPUN
XMN4HmfKQr+lH/tvUabCEd36vn2QA6vh21usmxXrgqzP6e8rNv6cA/hYOlJ+t+mhiVahpImXTBJv
s5bwkr+bpmi3MBo1tSqtSmjhpj0wNmiTmZhvQ4owo4sjca5vaTuc8Bo+U4nx+kX6MjgAu9gReJal
EKkYTjpwOksfqL5eVcfoeOxel1cGcL79bKZGBQqstlK91CTIE5Mlxwrq5mdUQxB+xZhlDXePjijt
0xzOoV1B7moPa/mZjvtWXhoep9y8VKyfPAgnN3qI2Td8vj/OJoIyW4HFyzapiZPhfPJNtVEQ5elJ
dpS59VaEbh65u7g9WT4eHIJfEGK0aysuO8B0i+GYxMssuerTSHiHYdlanVoXcRJ/TzDjs1jf1HBT
Qgoq1WJSvr5mB3DTqFbEI8vJhuCaehCMwKoFEHVXAkSkfwUD2Vv94bIayE2IFkVjtNAoAV8M251q
K6Wg1Hd5iiK2HyIuKJRbgl9l/tdUIenzFPVk3iGY35nb8DO0cFQGAhGfMJC2dXSAFWGGLJ7U+6SQ
+1SivJbGeKpFRnPWqQJGZhXOYrDao5Y5zDps+nvFiZr2nFlmYzpKEgzbpX8TWEKJBPtlq+DoiCXR
oAJgJXOfsycTlRSFc9v976qkQbh/6kvjykjmK3S64Kue1Ft2ZmN9StA3b8XPECmaJ3XQswNXpYIw
jseuhqlW9MzOuyYCn8zC5gWaxRZ0Vfx2Ic1W7MpL5s0P0rsrFH7W2A2ajHSGZEord7C7RLOrfeQ6
fCX5+1QcC2+i5XG4u0llWnHy1bZ2xU1GTDLaPo6rQCAiUt1c4eEnDQYplPCEuB8NGV7nMJcPebUL
Jv4HWFm1igqFVq3TIQKsOKnKzC3la7fvJocKtCxtqpDGFrVYQTIEesk1hROTJox9kDR3YyPaxDt4
fOvc1aXE0Z6wThLUyeUVQKfNRIs2Gz0CvFjbylxs15AtrVd4pWO4aHET3hyhrzqCH/NClWe5LlTt
pftNMSu5Ahhaf4o57Fzw25dDRJeJKrzKvjUaD+HNnYZQUidOk/v6OyWHLI9Kd61uxqIrY0MDwvdH
QS8N4xX/5FnuuqXIKv2S/E/ffEZqSXQNO1aa8XqeZ0Ziy4ZSNgrzArROYyfpud9T/mq5DO3FnEvl
LzKQ4BtI+88gEZq7P3yRhY/e2/B9UGB4PSmi073tR7ldwjpGZDGCnh6siy1rYqMAY1ie91yXdovo
A+MDPtkEL9AkewuJuXlMQ/UOrASj+eh+OfuIPznA1zd89BDCXnmTLVjroRv39C2V5bw22plMTZnr
2js8+MTF3YJx7deci0WVzO0FAe/frvzEqxXsTCv5ffLAw8moVeoEuzs97wYW1d0A582g/FadK31Y
1iIMm1mP4hl8ixDdBx65N/yhOGdyv4Ogmgcg7R+fHLF4PqnPOXqL2x0ECLK2cGbKaRyzq8oXq8EJ
WlSJv1KyRZVdJjvYETLgr7BFREyGnF4gxbyT7L5ALyEpvXGNdXwMzAVrmFxmQB16BCPBV0aehNIC
1naiGY4MtIsQSFw8PSHkFYy9fWfrpeeXK2BybOs59cslpixxYSPk/bXbiMVgqkrnMxsFRhgg1say
hSkLGpBrdKzrcEU6j9EJCxqXHyylf4tamp6SzqHtIIjLRk2uIYooAlgw79FucmtKRjz1/k0xJRTE
SIuuCkcksj48Vuu4rRcs5yqOsxWeWxmD94yW2BIkvmRjtzFXCUx/kgADzlky4xZhinOn82/ixYr5
MRfseSgi/bIIqEsnjJXz/xUi7z+pR0WTQLGRm74uiOEnN962o85V1OgEksB/RlCzHa7LwoZMf8xT
YIUnk4pStGqXMG4ndzmTtVTRIuW2CUKt6+Da2k2e7TyJJCb2tsia1og9LS3OHabyk59R372lv4IE
vJOm6W/YxjpH1xGMleBmFErgBjd+X+kWToOWzljGgmtF4RSgTAcujQJwkhz258svEw3Qn6I3e14Q
KETPzGvLPeHSmw19gDYRjJHHdo72A5qDQQCweqhXYd/B2F5k+m2tTKs7JhW5nu/Q27wBwG+PSiG4
4jNMvWZgzKX/Yg7L0WiKWvJGt+XrIELyh9RT604z1uHh+AbOMlVfU2ym7AxloppyVzNekZc/EpS9
/RvYxNNP7pX/CMrmZJNL7uGzT3o9dNy/wR5W9M6TBzNa5qExrW3VqQNN0NJuOQl1ugFjU3XIij3D
O8BEvlXGSMSrW8o7IgrLGprw3HJfHbAAXp2CiCTwhiJZQXQG12SCwyYj4fqGJ/1wP/bihycsgNVJ
siOVeJ4QSN2r9WtrF5nFPRA3Jd7CKo7XEG7Xg+JlxTwGK6VUhmF3vDT5U2AumxmU/Hy9EAgwml8h
LBMIefiWMzr1eXO1iY7/tOhq+L+a9i1dVM5cJhlx6B7/8p6Vnoy0R3llDxE4D6B51Cibcqf6sz6c
+f38/WuDMWLuGidh1621fMLGiC14bGjoxLgUnfZZSHQ1ivDh1f5RG4fgrVyrCC3C8xyYnE6ovQ1u
898eYZXiCQVh4OuZbfMb3GvLCQVohAXlk6y1GOUz2/GOwE2o4aXeh1yyW/FYu+eCUuqD7Bj9rG3n
uJodJXK2ndlvJaW9ZUnWmolV1OX52kfYckY/XZpF/KwyKPhPEeJdAQpW6D9OgSBWYDqjbLAZcLXN
10bPKubfmExKqJVMzk+YcAR35EFoZdtbOBi65tP5UtFg0ZN9ocLx81NJkD1NVPFL8/ZbLXo2n+y8
KTBwHjT2vDYyI5eA5HUoPTJQIP7rWQFVyANdwxzut4a8jyJhndYDhAy0cSskGUEmy0UPz8bKwoNq
lIV2V7wcblT3NV74bYlp1SM/ocj31yu6r/986uY+w0A7sUxVwi75b2Ar+fq5mosEd1cARkJBS+oJ
dtYWJwSeIfNAIxXOcuqwFGgv3b37mWsr5MrFPMEuxQ1QsAA5SI0ZOJa5vmvwlZG5LlnnSIOsKVho
ll3KszTDYciyZkmHgE014lP9xStF0SSwxy2cSLPVvOteyTzS6mFATDydV0urCtvAOG3sGpVs+Zga
8qgtmnQEbYcovAREw/nqewXwOqmz6KboPJ0PcBBp7ATfM0DgWxdCvedodvQXRFz3He+PvnRzEkcd
ljr7jhMh8H4ZrAMgVbis3MEE5mGp/JB9+z64PZKo50JpRfFkYGMZAPlCAzWzJYwYKNgh7QDHgPGy
1ztO0u02L+JiOlqSRTf3c+j63ZViyQUzlVfp5YPM82IW563X3wSehHITD6RYWC/c4z3z2AmH2der
UNJ+51Oj7SQspUj2Cp0daZo8lVDFSUZlUzwPZ/WccQoUNJJzV2eAmIDA99ZvsnJG5OS8qdx0DoYp
mGZz+0I1JBrG7VA8HoIu+HyhFeuH7fiwlcCXFXjTMPYEBAGXYlZCYDtTcNRZ74X6ymcMAuzgHHq+
K5LzO1w4/U19tke+Kpwf0YRGPovKDgQ8DpAf4+Qvu5Kpt3dKOTiRPu5CBKiNX+8Vu7Nql3Oz4tHV
vAZRGM+62ROWHL0qgmBua6qaonzBvgXXTlyUPngNxa8xNpdhP37kFoNjenqgVrnn3TvE7ZkRufYZ
hS1dwkvHffS/dGPSIIhTIEvbmXFGmQUBDQ2IGVoTAv+wOVaDF/6iqPESsT2oxTEDU1XkFKghkRRC
YCL5m2Tx+IzpISECai3xi8KEz72MkXZIIzLWbh95CFFrzOE4d8NI70mqH3Qj210BdSLzraMwa6dG
yP5CXPMCGOcJRdromhCtHmmNFp4m2AajmbUiw1DLR5KnId0nsWbbE9uDBqZtrMQ50ZsSyzUPwhvG
9uba/4wM4tP91TtU89d9cl43tzcK9ipDZ5oLSRY4LBhdCE8Y1vxIWk/T5InakUDLTMCgX3v71GQV
vR6DwiaV3s+K40SvZKYpbby94B2AfNtwSr7a5h3VAHkiVKJUKADkkXJOSUhkF5pUYjRcj0fQu6Yg
mQ21/zgwaKZtOxgjiiDSEOcQUV0l9ulIpZmCxe7RsuuS/gtrErw1u1eeuVWUowBrcL4FNznGgQP3
q4dxvaKmZcvuhPkVRy3n5zH5MrQ+rJu8BcnUJVu+p/qtWm6bOeCcOEgafzu/Iz/j1OBttU2imVcN
O/+XgBKEH1s8Uxeh41R+aAKrp+x8Todk60MSzYDr36dCpCL8KmAaf9jlNBz/X6uSmNtJkwGlHQoG
GTrSLKktELd3d6V8q/AJ3x8vJQMteP4V8c2XKcSWEHLw3/emBMn8unis3VTqhohG+sFYtQRems1W
gxEdhnTgfbHHUm7EV3b0IyqoyMp0eayE3fT2PWdYMmtINNWfED8FDRTlMb3vR68o8SckIK468r4F
FNsnypshcXGsQ+700MFGTwY8dTAevQ2iLvZHjiaA1CMxIN39sB0QPJmY5NKTAIbI+ytfpc5F5SKT
FKB45r6kbPK//eEinqOcgBqdc9lWPaniZWtwq1lsXZdgNc2+KICzOWaYfnr5L6iN04JzcfeKFKz+
R9/KoHbChX+5fvo3InWQL7tABX65Axkq5Dqa3XGkQ2SQc0HpfoqDIHWOSwhq+3HEFUyXm7mgkk9Q
MuR2DFXIKEHzt+ZYTLXoKmnMzWr+1bOfu9+632rX6vlRg0UDAlpPVTJbQyW6QLBnO6lf+0E3QOeg
8cqz6Cp/SR9gJa6B+xYzLuClZ9k6nj8yKASmA1xnCC1KNsKxH7CYyvtZea+/sJWiWJVKdVWARTlB
UhCx8EtRZIcoTwNSNKilZV9aU75hQNU6U0ICyprXWIpLWUt+hjQixa4ezsMqkX+hUrqZgJLqw3ac
JPfwdNOLep99HjJpZTJhCUUUFXjUyJ/UXUWITqIsQwHqYNfu39GybNF1uV/XLvpbL9t6W5vr69xU
DMZ1KlsdjR+UTKAmLB+4lHeCERMLk6kEBhTYtjSID8pJL2f/3PJfLFyzKQRjLZTAmtdKTY9aRa0Y
GKdqHm41BQsa6iOLUFm7xswVNRXGVlXeHAaTM0EM5o7Vsn+GEnMPkzxsK0M0dCJYiguOowt5xgc4
rUIaLslUvBuYu/vWqoVv4ty2yyWRgwtO6P3QINbAZNxSc63sntTZICBRRL+5QB43/e0V8QA3SNQm
WI7IUF2qNmM8YIZl5oExfI7faq7KJ6mRFGj4Azm6MF08Pex7LqUgIZHyUkNATpZdBdl+vG8MyNpZ
HH9MAJKxJRO/OarbFRRFti79xtNjP3AmVtPTlxo5pQMFPtjH3W3+oay1BXgWMKMqytpZHHDKMXTr
Fyk5zo0qupPgjNY7TQ1wyNfR1ROg+9bPJXnF8eSGgX+wD6X6G2M3x+MCwjHEAGR7HtNiBlp16vSD
wb5abqW8cs4nihn6I9vbIbWnj2fmVBcCA7UfZnr1ICA+KMzM3RZ6Pnuu2UHygW3/8rrZ9FU+JoZn
NxtiCidTT+vMcHI3ZN4j7pLLJZ5R/O7B+vcbD2UakgsLTzav819Yg8ayO6P931F9Gvpf7gfJ4tDz
DMArD1jU9V+EEUnDiP/sytNciX5czCNbW8EnkzvAnfkpP/aSPvoPQ89hHZbzufHz409NPAygM+uf
KMnwXW+YOH5Nc1lpkUucLwoUoRBTnqDHaeoRKtO+DBt1wNW/7Nszoy+/9DImn1906AGmryDqTRIi
7RmvqgOyFMJVWLvThJOrdWrIybu1VlDIEleIBmxoxQC4P+LIPu0580ldWfPX40qeH2pFyXWpP04U
UWM7PoxSowAnFKtvesH3Pd1qU1vYVW7MNTdDfKIR/iMyos5t9lT2YQw1TvvyzMudGkPsx1N19sFo
Gv4/cYTtm/sEBvaGpaBxacoOgQdnPHT8oSd5qIgVVKSfxhDSXQBPajnb5f32OMrnmjtJy4Thyung
TYLO0ESgvEafqx5uhTSTNpboRDeNVK6sBU2pN7DNqfklYehO284SoeAy6Hcj1DiwWbJWhXWUGawm
oPWbmGGx1JwjDh/O3tAu3HVrnatejgeYjPrZgSpFSK5UyyGZZ1S58h43C5G7aP9Y+mgluNzluS/6
lyuGaPeOAvfkWrSGmLSabL9S7MxVQ0MN8wKjsMvEwaVmHX5W1o+9NLXjcI5/GildQHE4q1eH3l4k
OBRojWM5+BmsgUopvtF6JgLKGw1rC9tb0gkgmKmn97iUXX6aS10VNGcEQs7YOdzsq2JbK7CKi6as
GWmFMRx31dP0WaIfwd11aGAa0aK/R1MWvnfAGH31kn3sCOUsA+kcAe2SQ5FfYBprupn14YcmET0t
TKIjCbWEhZcC/KYd/5hTfEpmjHyw2u8bCH5dUt4SZa1uQKSOsjvPatC6ZsPGMZS3yX/p2477BPGH
5F1c0AO3iU5i53MVoAM0ntVMRiAW9cRxGs+t5sJzYo2UtkeZSit/BIv+HPZeXEcxZIhp8G4YCpJB
x8cma8/zHp97nz9MqpK6T9ZsVina/BeTRdhg+sZgY4+3sQfojG8CTHTy8uqIHFG2tcNdUOacwTXW
HXOI2p9hPsKGIIk40gX3VkYltwKewJ/fff7MkKfOQn0YjKiFQGAA1hKS6bdKfGFys+5hCX0TLogt
PGavRG3kMjamVhvIGPvKGQIjMY3uJn0Js2uAbmdH5wYX0oCqBYn1Biq9QyVPU0aMx0R1AI77VAgP
sxMZQY8tXmqPzFkTGOFutj2KiLMIHz/8alY2zoFdRW2t6yQX7+ipfBuVi9JpeHvswjH/kNtsj8en
WGqvrJbhac7TdA+6KLYeMHC6g+9PRGQ+yU4HD5Hpx82bI+oUDT5aMf9m9bwVn9FFHwFDAE/B7wo8
fzCjdfUzqSwoeKVVC+qzJ/d/DTfPD+Fb+EZcV7/Q/Mq0TS4dSm8G5h3TtvRQWrk8oDU5+8HiIftn
1B85cS84SpACG3idozsic4AVa9MXZ4gaL8MjoDuGl1Si3c1IYZdv0yj+peInsyk1eh3TQykkVXm2
JMwpjHY00dvosBO6lA0D6sPq760FJ1dFLtP/+T5GXZG80xaVT5psRMeqY2bGOigiPccgyITZHYDa
SRDhRXViBGJ/RDouabxcAb9rbwQ91+Y9rgSu4MN9Dp3e+Ja9XxlZ5l3GDtdmyfxjA7Q/hxZCeUrs
WfcB/Wma+nhnzelNmlw/fFammo5lxne2c9VD4nW9hYsxfJs0ahoOqOmPt+4WgYYxstvwcbdBjt8a
XFslq8dcTD8FEbHjEtJZbN0VvI9zUnPPuJMytVP4Z+lMLQiJtY2nvGZ7FL2veQp+CfAsoej1x34+
So7LW+e63aaXVjR5mDLo/XfwcBS+KjeHtmiUrRSp7WaPXmvtmB70sgMwiu9bTENoAVHN0aw9n+qo
0zQpW7uVPEMAn9pVKMJDJphHfEKi+xDsdlrgAfDbvQBM34fIOOWlIb31uxdHn8OHB0ZwFUkMLHRA
qU04DYBzC2CS8Zjq+d9xsQUkhDj3my/b/+WYAwW4cANplyo8jxqSeAW8NZCTmnzCsyXeL4Qu3JE0
F3PuV6na3rU98JqwedS8BWB2fviQ9GFfhWtGz3MGZrzvxTwY4ZRoNm/aiCMdOuJ6hulgGJtxtJuO
gfy++PKwfA66Vq62QQOixtLzdw4wjnxxSH/iaP1Scf06WGp2Q43v2GJMiDY4bQCWGUWSceMb48R/
mexE5eyOq4AQ3Bf/POs2OOcJ4WGUTsZjIF3aotgra36gYrORFiL2M99TyJAnFQ9+pSDr00bbQRu7
qRviDV53Mt4LODGGqIXqt8GUevRPgAJLpSOa/QR2sxmmR8IOmXjdDufWIfK1r2zwVOu80fRel5hg
sxbcbBhTfcLpEEHBsmu/zOzrpuiS4+vGIAunLJbvCfYL+R1gUcG2KPRijMdyOc2vkMGR3ok71C98
8NmDizymV7/0wt3CJ3MGo0R3/2K/PXkuq7si58FyshkOrlFlsBpgLSwy34nQnwjsvgNVFhPwC7d2
I7kU76tW/7ZpQaDDy6Yy7AE6wCUmvGshAreUK6mrh15Q4/ytfod3sCKJJB06dA8ASxfZi/p2SBPI
urPRmlOZ+L0muQavDQHlrn9QkIFEti3NGejJdZ05x9BHgHnvvenOiRzlOjPWfg8vjN/s+ICUuDqh
msYgmYDXvHQj3s3vcgKZWYuuqR3ro2CQ3cKOvkTuqAaDhC1GRprecE9ShEIZoVMfZSiHX10cJeo7
ylLnd9KIkLZr+jh3AVP6wvapfG3G3T5ptZiagI5yZmtH6o99pynoJlcuShc5tNmJK80wkfGNSrHS
D/JCRDoCadIORnWnFWIBi8+udOO8DgBTDLxaHYkIEkB2yhHwVhYY/OJ7ns0Laf/WP30Rz2Ke+drg
/ytGK2fJaDQBrHtJQS5r0Cn7Zc68J490svJ5OeA8F9kR3FrF996VDzD8/TQsqrAa/DcZ1qF9yFc5
yPAjJ29kI5s+uq7BRS4hRttQQxjByeIGvOaSbMDrYpLvIP5L/yyH+AkeKAS8uscOBz72YkfMGp++
QwqPPUl0jawWCUE07sEf7TkcV1qSgHKibSraFFROV6RsQ1Tv7rEe7/XgWjC+hJnf+w8s7ybdqaTa
zzD6YwsrZaDz4YQpudL7p8UEfVnCGp3Gjw+dkIAeEFRXcCLnitK/U2gV3mL8g1jKXSvpIDBtJM3W
SJ9sd+ctFVGjMH1Do70AjEdRDjeH93DE7/zwYgHhpogqBsp+E/v5nD5plfg96zQA8y/mcxq3/VfC
PjcWSt7QLKDE2MLNPbqf5irKqc6JOfHfDjhDMP/JU/oqgyUTpdO6R9AQkFyVk/y+EO9+9mco/fa/
TXSHP0YBHWC96vunWX8m8k2LwZHj0ArrnhRiNN4ujtELbAjljIhRHm54OA3GzJEy9TkeG1AROEG2
k+EPdBBmSSkTQiYLRRSuFCCyGqd1795vPH9V1IXp+Vo8HpNkr7RgkHqh0yCKiLo3kjRGo1lYPA19
qSfe0s23O/dCHBnsoU0j75lcJWoW+tU/6F1zcXSd6V4yCGYKRUC5MBkRaLtmIbAmyJF0Vw++wco7
WdzTLNXhUQHKg1Fc4bvTTN/6GFyQBvk1y2GoQe5CMInMEGV0IJZQP3QlmmxkGEEI5rOytgk8crR0
ZJQB/2LIi+kAO3nmctlaRgtc/Lxp4fLmvgb602pNdmez8hQ2Dpk3poG/6wWcaPllM7b8pMR0b+BM
fMsNi370uAdcsZKLB8C6jf1YKSZmYF6n6k+W20uRWlv99bynlgtKXc+ZDT1rLnEsRX3zU35n7z1y
CIC2QU4/Syt3Ul3J0UYwKTA79KQeDNdL1gUgBHuNDoTkHzY8v7xIueXI7tXa8lhpizE72M4YQEAa
gNkWDe3Q19/La6oJ/ms9RGW2lwOJp/LRNA0gK2DdoH+QobdGf5DrAIy3WS0D7+OC/ssZx3sFDu3j
Mv2VUQFgFe+Y9z/TYMXsR99HZz3Kpy8UhGlamZIx0++1FMdgWKYCJp6HxMZfN7LBoEm6T9sntJq2
FVV7/FTC5kRiXfmI906XJ/REAZb960WzUoccos4XGMjh9ch+JKtunawOQ2EoEZaLIw0q2p8g/7IY
OpfGGNQOkP0Vna2HmVpvBc7lyfEhh1IVwd8BN13oxoO0T0ZytJ/Er4B4TidzLep5gnOlYWcYIVLS
SuTIVyIjMCQnCZyPZg8qmipC6Vc9K76kj5g+MOf+xd/C/5RSiL3mQoABssfSNc+1xxi8UHDrerB3
RDX9VQCaAmzH6dORhrwQE6kcPsxy0d8Bl8ZtifNh88fNzt4vHqjNHHnI7hLWqzIpiF9OjNP/XRpM
sjyt+MFX7oGtIx9ULsiRZ705zyOASTAoX/70Kcbgoe61DP5uwjCzjazZE5T4jZhbRk4t95Cl78mr
0BILr8cXQUxP9DuRow1VSnoVTDm/h1N2f7thT/t7tpPrR8fOS5yKiH1U4276FdnqqRXldUaC3RFU
CFbzY8saeaf39QYOrGXv4Ow2lhjzvWDZEoaGDDrpYreUkiCXTbyHvpvYh82nAv26ija3p60MQPb6
h+ti5ClFJ5n1B8s6DIbUt9xH8oOubO7yG6ELIOCjt2DvkYxcRLswecSeQ08oX8cXVATYfqyvq6Fg
DxbElVY8e5jdo9yHkvxtdvIZN33CmSABMIjnL42017vT2i7yzBe/OQz3PWnzt203HiCVODE6J1m0
hu25PvwSm+AI6JvAAxqtnfiIN0xOraq20YZMSsEIQCMkNP2Kf1/lKbIX4915bnK5W7w6IN4PsTbm
XO2OQiuoES7dT7IMXGsHzvf9Do3tEd+1RMYKAeHClG4II38zZiAoBmhRENNsTtiAny8gQOgI+Etf
uuL0GDwgcjUM4AYymFHlfjRukldRqbJzRI34bue5WWJZyCrc4JSh8VfjwN0H0Ffq2c8uauqILrWX
jR8aLd6p88E6et0JSqFpRvRbuv/rd/Ql8qF9rMH+wZy7GXW89rt3XAn3UYbVmoWd7ZFEzqRnw1KC
C/KF+Qt9DS1JLrQ4zc+aaD614Tyj1aG/Rjxv7InLlqtzgiMQpEAYgoMsFFJ7LvXord7i912OolCC
ArBJRupv4P1VORkT38CD4762DiWGl5DNwlIp67Z2zkhqHrt1XHof8YnPZsjyKZShsp42/EOV9TS0
qHQNCeHhZXjKBa4Q5ZuZyI3k1RdEOALzSmPWgZjgj1JhmiB5IJKnWEt+yJ/Bv95K9F3Pc0jC2liB
c5pG7OA6KrXVVHMU/EHanrL4bkqITzM/+B4GA3o30Pqdk231Qh7kZOaw6XqSpa36BcP2STGqq8JN
cijptiU3fynczeXIQMDCGtyvWXk63x1sHZHP0d6dZzweNNoeSMMdW9QKRLXETlb7bcxKPRbBzgpW
3gy1JGCvUSZTRJAaG3j5Jrr+CLI6/KkV5PSMiFh65A8a+PmsClX0mhgKe9G26jbSAAo1ecc9Xkab
VBv6Qzk8xYZOQpVH9tx53FTA9EHkGa0yvTYOUwY5KxXqfaEJK4s2d9OYZFgFGZ881FgGBH9T2cgX
Xahcj5oF3Z6mi18ELjuK/yYRrbOwg/kKnnEZhzy9K5uNX8X0puzj9GVR10ZuF40LaShUUBDc6wMd
IXNcMufuwBZ4j7MqKldCeSZKijyz7CRA9AaTJ+DI4dlKPBpcGcH+CWTXszs79H8gGKEjqSiR/DmE
zz1J7KUdrYP28Qh9KIbUQ6RnWqTkrvTWY2uLBJyKyRNBJp9VsvzUgbLBl5vOY/yDDw2BAhKd4ZLn
+yledgQQhJAALVeirTIfMS9jpRQo+g/C9WoGpyP9owgAdrsJGZBVRA6rJbvy1LbACggGXdN9yhkt
WeBEdJ4uWROILDnso1KcyDM1G5I9Cyx6IxL6ro1BPD5qIx+MLl7LvVVksr8kjeLWTqld0nubFgnM
jQPN9m4B5ZEYOBTzO1oyhlJFnqDyFFb9mbLLv47syA4czV+NFRfsfSGEP3zXFwbro+QxHJuDt9E8
kVxCst+VTOfeKsabcRTHVNFM7aJoxdrrEWLaK3Q4CsD2UaStCnSHrjtnNsMk66wyWZPO4uCO+9zT
+c0KY8QwRfcKW5su2Jqxas3OaxoiW+Jm23RKu9WWzn3T+D7if78J1DfZc91ocNem/nTxFRIVsb39
XVWKDV4QZ/G72/mkJY96lX96eQd4Eg18L6LG3xC7NSynYqJg6+WhcZGaEqHjSF1dBnSR7ACkjysj
J6LfydNhTdBqYT/Kv3V2Bjp5YbDv7XSKw3Vzyipt63oy3G81200aH6BNeyP+Ch1yrZq15YEswoIs
FGQTYlmW9WGIbTh8S4L2Ka9wLx2aaFXXjsRvW6V5sBdWkbdQMGfkiNAhIkN/ZZnbxI+AFE6jZ/Xq
hDUaBNgefq+GhmAjXfBTw5aUZB3mVrzDwTxrJMCrXWlIusJtQ6x/PVGTctR8Rn7ACsKdFFoT/aRj
c99dISjQos3zW2G6iZFZzlqZDtmS75KJaSgl4Tj6/hdI+HeVg34042FT1FEbDtIR+Ss7TPQr0v3D
r0mjC0OSYSg84thDfwMGqBeXTu7QHrDzot7HVrX75Hzb+RVvXN7DKuKkDaIurPXOIwuc1ZqYNNY+
kbp57K6w+v0vtIPL28nsLV+zgB7zaU24FTb/q/T0rKBUoCX9/+JKqo4KsTnB98WbkQ5Hb9c6IT11
PTONFuLP1PBDQxkD3TCUm+IR8sUDa/OprJ4U55xHChwsXyq96w7AEUlCAi7s1jI6A5i/J/lohfGd
UJ41crRShHIUEZW0awdN6gkmZajTlPB7kPNAveJrw0bPfOb0lOhvooA/quGphcUkdsn/tuNnkbIA
S9qLSofbcQJSCedixtAuKuOeK2IBySxnmzEM4ZfA5iJ4VIggVia1FliZPWu3pvqkJ9Pq7sW+dRU0
aeE9d5SLJRMKYhizmjZRXW77MyKCfdwdEG//VOnjWWaBY+btMUjD10ZlDcAOPLqBwFHne0lv0zIk
GuwZqFOTMEDazz2Yk7bDKbU/JhjEWLqMLq1qqStnfbyqXJTdh7nVqu+Rybf98auWNZVPxG221IC6
xMiUHnnatwunqVRt6ULC5wqbposhyiXRiffNA9M/kh0+qvcoDKikuqmwmUCVHRqpMk7N+G8AVYIi
HfPkaM8AU8aR9SLcnu6HMoXSVf0jJ6OrdJALbeoS6p+gFD9AapsdkDsRoMEfPQD2iiYqZIpMsVM3
+e4tiUwKyLYM9BGJ+Wv9BV/BWiNBRQkU2yoSwMNibXcfHok5xZ+urkn/tB0Yu9ukFwSiEkOCJ/qR
Y6/zRkPmrHoUMUNklBoZ4KgTWnPX92Wz3tXC95QJITyhx66hUKpwj4p9fOcujmerUNGgzE6jvirA
/UlD7DBHW+VAiYkm1IgjBmuk1xUjAji8e6LfTYnVqvxED2hFZsbMXPiGmBgZdVbatqGyLECSEb8o
XyVLTokzRB0gsrnbJ49dLjqXYihDmXYWoqnRzxq+Lx6hFuHXgVlnNmpoFin4JLA0Y7b8CVOcKG9I
091USuLSLGJqCwV7+H7Dn4+mj43Xg+zwPxuAeUJzXwBvhFeznA/nwMVmZUVJUpqZChd79HAVDo2Y
+QGRMx9blVdqtoObhE5xIScPPo48fvFQChzhJAkkdz8im/C4ms5vUBdctsqzRGAB95vsxsj6+DU9
UN31p4NgLQ9ZkfALpee3EHZaxhXBvThvt2t17nR+6PAKOYtdcgKZp1rLwqHSxO6n4zgUQ1BXzJfF
9IxL4n+AxOdqbqgp8839V8iBQ22Hdehf3Z85PKCAZ80kMoFvCzJpSQEB/JeqJ8ckprhGLgU8b+XU
UZ6Y3UYo2Crrsv6qsC5dv40rPs8Z7eHXSCRuzzsNMPZx+OFXi3/jqZjru0rvZGE9vM7naGBROUYy
yzGi52+fcLjDiqJx7UBHrzdETCHA444u4nGpYNhkQrgbvcBqxZUdKrWXaElbf57BJpd0TJdfD23C
meMVqQSpXuPU/vWgsAe52hC6xwoPVf/QDtwloWfhznYGpzP2CAqB5AKz+0AVG4lTbT3d3pxV+T7x
QwFmfD61ZJiwWEbbXU7o4fEaB+458XwAaVh6HOkccRRsB+FTWuS+0e03iWKuZNWrgmPGNpNRVijR
dVBc3GLqKKZFe60RqsfGfMZ+N/J5BpINctWNI0OTLCE1DJ87SMCJecDy/rIma5R5YgeZc8mwHnj6
9MWLaibYwDIsxJuwJLttZpTxbo1swswLiFhxLhBJZCwaSPH2zFTf8mXZx4g422ExDAnHiZ0Ivf3w
Frn/upzCT5odM0XVwfLkgzGe38rMlElh8JZQSeIe1TEw5L4hHGI/MfT8ZrCz0mFJfojeqMFfI1Sz
mWJiiN33l3hcZMn2UoPCD0ra/YkLVKvyGkfmSwO3/s4v8lWy1htPAGg7bXFZ/QdryW8A2cPIG6IB
RpYyXNUH4WTEZHgEVShMfJCwucbSJAuIxAl853tSUIPJjxNuhGzXpEzZHbYKYO1moridmOwAWyHU
rggQxN+wlqrZjhQDNV8Gorw46Xn1E9uyAgYo6XeSZRq9WzWalel/KY7Cs11EmYJ3Qr4C+g/VNwDx
XOBINzod6r6prq8tTE6Kt9wzGfr9QwGAMDGFNs1Fe95vQry2z4ZtXMZRydqcWm2Jw8SDnnjYcgvf
8ukmyO78K20VkDtO6u9MW7IHeAyyeP0f4I0bT8+VzgoY+x+LCHI4bI6qalByMTjls7mRhWkHj8Be
1HJ/NjEMjdHhJhb1bosUXEZABZXFKVoLmlpMAlAyXfq1vBoqXXJFYFWZsr7NQ2aK3ox+TRI9vJ8z
u9TVqB5CYm6fX5WHJ5+kfpRl7mBWsTGRV7x35PdZgmuj+sbn0pnpeKmm1Zr2N+qD9TnTJmzoUI2V
T1S28soFzvDJxDZz3Et/h+jjBmJorAbwERQoVB76YSeORQzm44TVjJWEnqOE8kCCSf1szTK4492T
hbbdx3Q/HbeWPA6SLakRYljYZaM/09eIkaonVfS7w1YrsEmfVV0oG5at3tqrmHUDxX1EyJH+qHtx
vdZiVgM6DRrPgGtHUrHbyHHvwSZDMvssAkK6jiORSgkIF7IaL3VhtZQsu2AOwfX+1RGzBCKu5lAG
QqRN6KMQ+7Hb8biBMThYXNhm3nZ4+lzaEshYM7NQUc72/P7N0KgPqqiAs05juY2N1LVs7gdK6lrw
bhqAdlwjPg7vu+JRvsVgfJa+xUAYt931YM5xhmIDN//JTsdbN64TUhacHt0jYg72l49aHpnCFdaJ
hihzAnV8GgvglP82H8p2YWegn3uD94zCBsqhWToPbSZNUPLYbRwx0aryyFR0pACYvtwOrJicXCgJ
SHuPD68mauFSYJ6NPaax0bJ5+KTJUsaPoM5lF226JldYYSHgoIkvNUg7UJ2D03yKyUBq4ATS3H4A
kB154G74m0nLzE4rmlat6Pkvmk241RWok1VcNzyBQ7QP+lc9aMmTWah4M3BmkPnnYG8OX82NcG7K
QgPo7Cmu1wJfr6BHAlXb/pJSHvsj98U5kUhkRNzgtJ5Fl3kHqyJLOdJIymEhApdIJ2crQ0gA78Ud
q5lX8vtYOsOYhxVRI9bZk15kllLc/B4Fvtrnm0QFG1bHAwHBuW5W6bF5sVk8gqDzH6WVCydLqj23
YqHe/HFsr4MlBct3xZuMgIZSAluy4AwiamdWjEQDEGa71UixNFowxdNhytuTgNkCJySR0xDDJmZe
FbPPuSna3k/RfjstWpJ4j0IFhDmd2pCiDxxCngSLEWW1JOaBJ1xFeFK5W8JG9gOM3iKMu8ylmbXW
gKtUR7HB+cT9YDXdLVyqO4Fw3Ixw2XGSBXHRXYxzbTl5xyDBxuYIKVg+OTppzhnTl3Q3liXzCcUr
8nsVxXM2GcmD0mprXt6sVkdfeuXcPx0MnxaagXu5kWYyOhp9AWUq+ZN6P+VE5+xWP/ELJ+5qyRtm
IywBAlaYGsTqraWdwEqoATEjCOll6mtHJz3rAAPG6wkbLfzaQCiURrMVWtR3PpXtVFKnLBt7lwxP
teVvbDU8/N0AKrxTCK/IeL3wZiiqqjHYnfYvlxZzfzzfV3XwUCIeVY3KY6qvMqnS2QEdieHeQljn
4fuB6a9t3+NAkpU126xQnH8cEbrzrYhtrd+XTuLHN6CVTi4ZoA3HPwHgtmzgocuvgWdaWawC4u4E
6BX5OGDrWUAYy8L+wAlKvbbtuV3L0ZWCV6F56y3f824xbbJzV+TnDPcYbHcRLXKjaCNkpWseB6+n
CazQfW+1SsDbCgh8IpHXgVDTVcP4OplNOxtcNLGvacnoZXieqd9wVwxs4Gjtx7ZQp262Y8GWovOo
do4aszH/z93CbtPn88zqg+o1nejYuNWU7afR4NzZ6ImsjvmQO650x3Fh29BsZYIVb9ODE2XzIMX0
cv5/3zTkdqWNWAdbgVgbUWWdzTDPMZ90W7jlFzymQuadjGpqgghofYpiEMMykU+r6beJD/ta1Jy7
2AA36gJJUSxzLZOZK6H6oldg2f9hTF9QqUUxuPk4Fbg2aiDQHitT87kuXMmjV94vDrC9tjFZJou8
usLQRlLAZDdo2nSQnpXQ7X3/pwe9W+dcKOByC9PUA00wiYlokRtMxGFa31eFj4UiF/8E/W6lzK5N
/K7ZdMMh7wM1n60RJ6bUEhH7zkStKLyStgZUbhzdLvyhPXIDegCjzcYK8lALV1EZH+kctDlow6x3
h8ypToChw0QbsDhlpHm3Q3ZoPoPtvz0woZtMU/pkiEaUtZvoq9kCFYJhtcqAbKCPaUevNcsAc9NP
4r9oTlR+ZADe5qxZBuFtCwqcmR37Cy+fNmy1Wot7GqE1BweXDRTs8xok1KfGikgowFXbTjRKCP4j
Hkw+YjL4kziN7vQS4VBUW6hlIWF+tKrYBtKylZmVelDgvTvM4yn3qm/wkNsuHbH7WfVVEYjvIHf+
lHrCRqRQRYMKSyfzCQpiXn6yThQLQfLDIXTMadNPIQt7fOSg0egyeJfwcAYBwC11LoZaZCI4aU+9
Lnvwt1Nt67lI0qz5eGtnN+zMOtuV0M9RCy+n0VaXV2Yez7g39ni9zdwdEJYpU6XmoF9XLR0VxRzQ
kivLmsiWoSVwhv7R3Z0Bl+Z88gOkH0906wfHZ0hyAqY3XLYSXpUu9fV6ZLLADo2cOahwH5wu2Pxt
puaLx3lexFLuu1qQW7K8XGWEp0/AtIKvaGqqf0rj2aFbNeU8ceOwfN6F6M8/rzEQqv+ITC6hhQ0a
Ydk3G8cQxu2pXK0YMNTpY7Wix8qql0a5RgnkPQ3dQYaXnadlcdUp8I0oeijgr7jmzGp4z11s6Pni
boTEr5+GBsogF9mJGEiBx0fXaXDV/N1zmmOgrnG1UPlCBSHLwGCpggadgkDl/u6K1hEZKP0tUeOZ
eVzZO1Qg4GyRD8/6QrVJBhl/TSt+UcxiXJ2YIqOwpMz78MPYpLfpXlhdbVLCswCjz2PspXmgyHU0
nWSHeyG3QXLj0rBh4vy5B82hFvzBvdIJSiRnQSfL/7WGWawQIPv5MJgFHfXIbp/qHhb6ysAFhr6w
vuNY28k/gufDrfkH7Mbu/5g7E7ZBIUWxu0HTszfrk8TWM+TIj1O2kfOmQbTVqx1N+N9AmE/ELFiz
R17KZ/glEay39igzRCUp61J5w+zwMDuGG7emMdeCFG8M3H3C8Iv+insF5JWK6Ttwi66MCDMtheph
Lj05z3UuqY4LRyWACbyUgCUsyKVNLpzCAfh2FFQULfc8lhogthnqim84CMHuxJPLrtr89qs+OdKI
9FYCvgMP8XMKVbg1q7GMNRNFmSw/3AwCW6VVUV/uqaZS3au0I733pzsx5/dX3SvpqcM1ijVzTMcK
Plhm31C4pipqsl7n+d1Ujh/BiswSTPjei3dKWtqyJ3LlrZkRYVDoQM7d9Lz6a7VAFGK/4luu/J3P
NeDIovh7053pz8Ox4nWL9VMvmg/GHemhx4ujXYOirNs0OEyRZv6vevsCl4Iweq6PP7z2xBRn+jAY
UOS/VINhTfVcqAJbKKwjim3h5fZVtE5i8ZdvyeryG+EWFcudJXldzeXYH49Zoqg3d2GeVt3PLAT/
Xg6vHCKcSkTHKDwLraKMPx+JS99mYd8fzdSWMgsgpCc34vT6MY6lgk+Fncje0wuACcNOw9qNqwzV
TEm+EN2GbmOEjWDNozlgJ2QcN0mP8VQb79vL7uTdKnb5SuDg3Iz96c8f1VClV8FMTQDSTeY+d2oq
IqtCMSAetFw7g/fxBq0tKbMtm3kUfI1++OOlsE+8fleh9bgfWq1qrVDSsVvpEDrWfqPEtgryeRDL
nGYwzIBGaEx85WiO+xdVsMtquPr2TxYO+8pplEgof0w0Lsvn8TiwRRdlU/yUvlVA7InN/kZLf0c2
Sglknjb7wevdfIul1nVm+BUQn7vPPZRahfLwR3xB2UgrJVL0nw/9kqKmU+13jkXz2ftZf/t+mg2I
+dOw8MNFksRGiz0F671cF5NWCk6uyCk3ewwNMIMx2VQcN1lrbTx7hFMOovTI8RQmOxA+V5WXzGDJ
NHDn0GwFIF42vVSQddOex45jMZLLxRpHODFPBB02zPzWHOfYwDCJLpW5Ew6sKBHbjblf2XfRlylR
j8RieaOL0wFryk0q5cyl1OFGHkPH3ZWru/MwYUyBC1Ika4w+qGOeFKM4nNiom3UBqa7OElhWmQwv
q9vwBJWAS1Ung+HZsRDFvGYh+7tsgOIDl4sJLSEcy2U5M4WrK/RSe08xSNBXDxnWAfY07B9YiFQf
Du1UXWn0KqsGKMXmn2glpLJPYgKsZSI7KBuJtxpbOaw15kE/2l1DDm3i0GFizmBQcQx/MxO3vtPt
eePldamUwLoNYUY/8VW4/IkuajrIK6SElD8VddGS1AshN8R8DaJteEkfuifMQkdvikAstiPb5dws
+DS/Cvo+dtXnrTh94B52uAM2sR5e71MhKoMSXo4vLzGAbGzYFfhKWQGoMbqT/EfSs8u/OYWjw/iq
mfMAy5GXow/k/x0/8o4YbBfJFyzJe00HqCYXlIQ6GzwfyUk5BFI2R6qovp3sgryxULeWAJ/ie10a
btF80khPjL6YvccqNI4rtZjQ4oIf9GZL6UP2GJLlGcwrRIyeroKssCqb9xnRhSWuKZinTwPovS+V
C2cGyut/uNgDkdDf0kMlAzg7A+XgL+6qdDBr/KNwMZyv2sAADPbYyrKtJhVWukju8bPav/LVp3Yh
jjj9VMH/SkaaF9dazN4KU0rojk3CDnwUHVssM93njcgSoVYWpQbGsiR8JNUyNqW9WLL2/5bt4xWh
gHruh6QqjpSf1qOPkec/n7Tjfq84VaNCmwchE/YJD1pivWnqrfMW6msz10/BVetaNq0NEiQSFWDJ
VCMMRkIob+gFOkrDumm0KlJWoU8BjdZaIXd9WSDihTMF9er7Bg8K3oyWi9p5fcRzkbe2/JH8a1P0
u3Iutv69+KzjGmekE6bOt1uX58GQhPcDS0uRMh3oD0n7N7i6B+dOhqn3B6DdYFY3Vrs6iPyX7K8z
kovAspR4JGf1BPOKmzEqMDKzYzMRkw+8uvcwTnEIUUXVaIW7TIdoS+X6ez19dM0A0j+FPvi6B8+w
hEHiQl2V6skIOfJp13P0M2asaneHqvHIMKCGUloulCxaWww6PHvOW1ljVtmOgZqdfCShYQjEqAZm
OE0HFUKwi5LVU+AwvPlr+HA4PsPmnaaUAZTERlWi1xpcb6wCCfv6qcAo1GpGzP+HHlCttm4f/B6H
BFDrlfpKKs24G0PTiix4LbZKh2LsgjtG+oqgzY46QTx9PcQjDoTA38q4uCz+sszMrs8tzZV3yHiu
TS6fYU4xpTXVr9/Q1APMghw8T+6AHBZYO8ddmPgJ8M1zCS6nIl7RZJqQ6/sKgK0CpW6PqsgMU+9y
eZ8aZwMVierIsljbuE3sEG5/0sfNeSVTpTrHzZfNCfeKG6L/cjlokIIntwzN+a16Lk2pAyw90z/w
Lc+rsIWj33G2JbeXqR9ZVaQ4+XKkL65eNswOBpVgU6BI31s2IGz4kV0q6jYUo1y+iPJwT6EJzCpH
dYi3KQEdi61UXEx7p3Vz/IRnT5VG6SKcre0G2RlQvFQ/C5k9CKfNqpLVcV9e0QRMwtJaSlvs2zsn
RZW4EGiMJ1/A8rOzUCvnnpg8/jzPHnqsqTV7XQ1ejS7ieka/VUamf6LKg8GWQ1R76bGfiaNUx9Ps
xIPXwKe/AEdobkYulP7CvGxiMXQmXEF0d9lGxR4YoeBS3C7YOEWJIFyzdmNPGy/OKGuNDXmD4jf5
gnAd4G0Y7pr2MJ0HCQgX95BqtKuZJglVhZgnsONWG25JE9u8z6Rt1RRJnjbIxE+FR+zKYw8HRgsL
YFUlzqckTx+wq698c7DWhpUY3o15LKRel/VzTKHggivDTcuE9ezdStx9q0j2bBqLW81bGm2ARBcA
3eecm2ppq7UZMJdPwbzPnH1kjelOSHoZ4jHgLpZn2yOCShX1zCt6Ps1tIdaiPFa4PKDLlNmx/zEJ
Pjggprna33S7NXYJ2hJ3GTFGJ/BqGzzakB70tfJkR6DDFbKdZulEatp4TbXZ6w766+xUeytSGioI
ppJ/haHzqKsl28g28Lvx1OqdG9wGvutGPdpu2i4duW5CkFu7kex9zWL1BYCnb38j2VKKdNJFomhH
vbMjf/d2dJJuFN6fbnuV1nGSKt4mtMQ6gkcOiEd5mwBBOrL/N08NCWkvT16hi0PWNx4DDZiNeSdW
cUpaJK+pO/1jQxnNFDMdm9A9sf8yg7q7mj+X7VZtVHhZQZ/krCsiS4A3dzmYp3qvKidpe0XvXAcp
3OhTHHUjaU4uhG5yXESFDfgYPp4IzwSI59dLP3LWa81l3wd9s3C8qUUDUw7X+WLkuljcawpEr5j1
c28FK8wlnu/U8K++IWckkAp8/Td50hM+c4PZSdbcBGb4VXAR9hxZD2ehF2OXj2TJutDH2QK36LpM
nfZAWqIQrFNmTLDtdLEs9CkkjgdmU39e+cUfheE9UI/82u4p3MTHLv8QAgEV7ozdBkjw7/zmtoFu
VznqWwUINewj5cJomJ5VoiNOWGv8h720M4/R5DE+xnG4seD5V9gfvtt7gE04K8t4bexoiTKqqAsi
c/fuUcGqXaE9Zg6xkPJgzlBaGyo29nVTT/A7gp42TVg7UeGe+piE+frb/XSQFfk8sHEz1QJ5GS8T
eLKhwtzSUFYl+5NM+6fQcRLFm3+tQ3Exe6vOd9E/9JjIlAO4hvaUV5wgXgEJ+y8aJNkNuRKf6Bm/
rb0fEnk7HKdPyCmeMtGZtARPTPOmfsUr7ib9XnXeE4V4iP4+a0LO0MdpSfORK3FfeASM9U+m2RGI
q8cMGAHq9C3/p9tAsS2lq62t07i9v90fle5ri+d3j9IV4mNN1/U6v3DqDzCzCtrVT2pc+I7/qdwz
17qiJEpcAMissQP0u7B+aep908jiD4jaC/VVVBoBZKGKUvblosaYvO9G2sOf1YyGP302zoT6aKCz
/z9lkGJ4AAhISy56F1DMjY3E4tPiZUbhQfzhcR60dvoJqao2LlVRmIisSBpA/+6Uttr7WKwffDTr
IUjLzDVYHQu03odoiH9v4GhcxgecFY/CJhQ1u/JdmF3Jd0K1jRuSDhzCB42UQP9OFhbG+7AxjKyR
aGia/vv/+tCW47k1Lbd9Ou+JOgVO9puetrzHbnXnJdQo5mdMBA0VKdZn0cwi0L0ZYs/9EtfnGd3X
boiqH5nrINj95YBaK/5o9r6KBWAgYD5T+g7Cq4xxwvlnDDcK4FbfBLldzhOhayvUsoQHCKWwTqG5
kNWATiCc0Nacz0N58LKExtTWBMQl99YI74CHblqMxSCbolU+YPfqki8NJbcgEZY5JWIae98hq4ZM
bU185ygqVoNU4SoG059xek1ogIdYvkl/rE55nrrUNPG/C2VXqh/fx5VN9Psu2jmJLpdaUehStAqQ
Ko1WRSk4qHIBCMhRyyF/BATsKJ5aKXizG9Q33vGGbPw4ewFZbNXW11MDOpivqRdEpCFvUsU6ISLq
mLEFCC1dqH2lYDF30zyejXFnHCbrW7/hc7/1qyfhGRSUMrTxS6PPY4iAZw+Vhlq36hcdqphwhrM7
QxbSLu3xeJuBStN4iqLOX37ZYxF8WRspV0Bfq3gVVpo5ZYKEoFYh6yP81HEVpfsEMEF0x2x6d2R/
bx8sdVVRxonFwwwzGXSeyHeq72hqsKQuGBUy5DVutLHbPWfvGz0XAhYMHQ67DktFUZKC78GDt5xt
W1ROpHxvvwtovqLNHNGa68UoOm443Tb3n4EZ3JISw0UCZ/sBZh0jboRaKD/a6FDOHxI4E06DNSwM
E8AxLYro4dYzzOjQz7JRi99mw4NT9ydR/INgomsRIxftJQTBYEqtfeV+1cU01DcpzpevCna2JtIG
pHJjcVkn6RlrgyDuvvYhPAp2YMreNOVYfNFLWw9HOOboIWTJZX7mwIZwZ47EMJICNNQjDOHfRVz5
gxL1eJ70xRG3Z/xKSp6CbBkPyEM4bp9Po7dEJYcSBpgVQOdtBQHLYAHpaVWzWC9DBAhuJh5OV2Zz
Y0gYVywammPeGMnHT7Lv9Cc0t9pSkOu3FssSkfOdFCxsxdwAacmzhyLyuI6mcx4V+Gx5Ip+VaTbX
B/YKfQYG/i6hWAVufdOSBBXy+Wp/3yWoyzn89vT9cd6Y1BqJZqXtJjE3tMITeHQe7fEwKaqoY9xh
Cqwcu5AuNRUrzE0+osuQBTmnTeOmDY1FxcriXLMLIt6j4+S1zTONfNfnLkfIGmgKhYttj1mjcB7R
QXXBpATxBwmmHRTSxfa8qvYWDRs+2DfxNx/TAmdXucwz21ywBGvwXeN88DI0N6gAozjyM+7eOBvP
uTLhhOsF6KQpciZBXMzhNMWzBCZ1yVK+AZ45EOJi5RBMhL4763yY3U870DFJPbaw86hNRDawMNqf
rG1SosYK44PHhUVQJR7364VyeoVLgUNqLgsIMMVW2biN6urermN4DBCxYcUw1Q+2FwA3z20Z3kVi
X1a/OXlSITM9ET6+5KnRg+oI4WPOz8HEGx89ktSTxmeTN/HdfhMvw3yRcPYiIu930TrRzbvogQde
W17p4QuO5GycKRGcoEILdFJPCtKvLyHcK37603Cg2vwxPp39KiDnOtryKBZvewoRGe2w06xLkWz6
5oKdE6800rO1IWOOKKe/0QAJmjQZZNFvGxpKXkmlqwdYUDjf54UL0h46wDii+BQt33+i/Nycdiky
ERNIaFQyxM0JQCPJDSm5ywSUo0NR2I7d8lah13FiR2w554zs22jaVVca59NV8dr35zovuwuV7d/C
4AvLfgDLZM9ojgNbts8EEe7yrQ69IRDQ07CLX5NSluX+MNa2gFa6MhDpk5mpeB+7NCwzDpar5rBL
PVZBI60t+29qK/J1Kq8x0/POF4ixpWkSGY0IFjZ4EGlSajVAjRwOPCZSmKped6QJAq+qvTcbPnK0
UoJNdF/9xLxXebfWpGnaEXuQaLJiFGSqdM8/4Kg59WiGG6t11XGs1+1pjpX4A1o6kIhNQ/3JXBBP
4CpHdy4Pp3sEuw/dg5rX+xNLiqHRl/AwjIPCtUAZ0fK6y4YKkWLO6zjD/tJ6dqs6uWY/+XdLp9H5
GXPPm+fpHw8VlsL8ZR6cuNGDSCGXKtPkCw2nI7vatOna7EC87Bw7CdLtRTl6pXpdIUlP5cUcgJag
yJunjTUrTj2rR24Yr3HBLaIcd97g0zoID5e+xKaAaTEKtZbu6GPjVFZPhHQws2MhSaiLpxRNYnUe
k7Zg68ToUJjfbJBjoiPs+CE7sAAmN3QyLAPx91MBvqQMAtHVUNbLNAXHH4lD1xKZVqsZ5W+iVF4E
ANAPSZzFuqBN8HJ/zOrQEg8lXLMgZILcO4839w3HE0wPYTtG3OnT3QsaEiSiF4l1gk8UYSJlNS3L
tAKVMNOgFLaJcPOeVQC13DFrNZsswgT1f0WKHWDCudWwDfbsp0wkBLOmli3+ClCQrMNM8qaNghIc
ele5XySIRg0v+DQHU0FFJ0e/4k/COzAepC+QhRjyCTIYJYtd0BuUW4+cNlQOT2GpPU+GoueRyrzY
qZA4mQqYuZ/pvNiXciNE6Gh0LkhGgX6SuXguYW3ONEq6qXkoWJuH5LamNQHEmd+3KyFjHeDhEZ8x
rTf5AWpFmf9stlLD50eCTy1+1U14z/3FuwxIRNkVQc6Jf04qSGxZc+ZyV+QcIkA7a0snxjhUi56x
YZThZO6AQqwR0/oGHDOfQ2taEFInJgupFksuS34XuQRT3LqhdIvytLZxQZYQH+MbHbmVJmgXyII0
0h1Dvs7vMwinkyH6T1WMeVmyuLdCxCtpCkGpCWFFSsOE2SE923TC4fwjSh6C1e4eDzBhn1x+c4Pt
u8p+9SAN/4lFV/0cb9gOC41IlMDhH35EGwz0F8nOJ/b8djV2erIyisOZOvn2m8do2pdHxg0FI+gw
ockZFIdBU062d7k0BPtGnRDFmt5swyI6joW2x7ijRHI+t+l+YAC4gHZGUARxlR1er5zRgUoKX4T5
2p5TPRVf1CWiM9uMlM03rYwwZDu2E29HWKwDash5uUDrgOAtszL8C3s325cAh59zUkiN3qeFbWmk
z/FdQ7arQHyWHMuwvYq+RI9D3S7kv9k51pTfiEWbsnMH+WFRvQsSDwhuPg27A3FxYLYJ9Vj1fXeA
voH7/r0brv2yyRGNo0G75vaFbB0OxJ1gX891qGfehqesfJZCzQ0n1cFD+nIkalPonwLy11Z0rBx7
H9dBj6Mr7D9PhRPazulUHKwCyW+GngL+WC/8LMCqjB80ssABPvN/C/aVYwTmOiogW0M2pEZIqkCB
12fUOf/NHKmIcBvOosU8Ipxilg0rZB9iI7MRNOuYq8EBFV8x8hu+I8i1e91bYTOT5YXf62uaTmAY
vmWMFtHX0ucFd7nh8T4MuaqjRXAD/3nl76pSOWgca6C5SP28extLNf0LlXBp0ZI+QDC1EeX6ImDS
LbWr2wDpp6tT1I/2m4i6OTQih3+lwz7yIiS8nCT/9C8reQEmoOafXXrRQiTDDtEroMhGA7CwuDvI
+Kf6XlharWblc8fO2G2YoYN0fUOkc0lyFvp8JUfgqy+s20Jvr8U3cHiCSZm2xTGKA3M9AuF2DBvs
dPMSdQawyCCUEO8DrnDeCd3fFtaFiuppJ2zGiCh9KPoWFV22HqVs1j/nG1x8EAUlt0gXEB0B6Ww8
a6DTYlVmDm2QpI0g5f/RwgivvaGQjxN30Qm5f/+8zC7J7bMshaYVerzfKmNwbTzf3E0Zi+JDVNLK
ykrRhaL+TFtiYDzQEQ5mUXcKjc0D+3qHhKAE3KbQz836Ug4uBzhI/bfnEV2HHsTvgwJ3g8vkDf1M
5Rpw2fUblFtMhae6aqaPSc/nd+D63LAR0T4CegTFiklKDWrQ7nh0sLnCz0ACn76zdJXdEE0TApIC
1M1lpTZqWJaMB3ae4qjdl0uMOMDBbCbDh4TbRmTBcwJpUD0P9zhDWVuf9NY7aEkxc+CEb0sEIV39
hTWxLL8n98yYv1WQ9XPdQS2cvuQ8l23fIDLKeBGJDSK8o0AjFOV4AiB1Nzyqe1v8Ma3UgrruDdMJ
SodJWW9ojy6aNSoi5kI05/GgqLKIMgD7v8yLaH0hIupM030YKTt7drGVVlly3K+jU91CL5bx7tnY
VYW67b7/FjVqxrQQN0vfHA6LGuvftF8W8QHgfljAat1C7VQx8HVKrJziTPfbEhHXcQZUNTSQR4sp
Z6IJSUT67blLrbYTJggOnNoY1jvo10ysH0PWpbqlFFyFOWHOC2O9wP5ONvAFIuLqz/XQ7wFgNJGK
DA4WBmjYPpjY0j5VzL7F2+kVHR0tw/Bh2NPIwU1prfqUsVg5O4hGGb+Lvlfvv2XqmI1Lec5PIUz3
OlFagBwZ9vQdL8Y5r0fxrZGluecKCkZUdj1OoQIiqWX4fbFRvJ3c1xi4NmgZsufXzLw50M+qgWTc
KU7h6Budz6qRLMBF6bcRGkZtmQ2Lq2YVueHTV5iZD8RY1SzEqIJsI49F8ceUyO1BqQuo4LYbza7v
Ogjd2QHJQw9Gca24RZzWip247HzhZ1tOpU67nCwvLw/WpcqhibTRVTGWjHU8ONFf7IRIpIcJCvlh
Loofssq+3Mkhusb72iGO7hWElZu8rvTN90MBYoM3E/CR8/Wa2Z35Pvgq/7U9ae6KmZxIcb8p+bGU
/+hvMKurPFyLclJsYqEnw/KHkzHRvWyTK2QHNH+R6gQbctvaJNZZRgNa4evKKOSiafQubObyKzJX
KN0b5zURO0wNwz+/AKVRawY1gdup5/cMiDP/1WIedEhlcgWzndM+Ou86/3qlY4Cvg5WuDTe3MmHr
ggi9luhVTFG6YnTacj+QZf3olsfRZ92dyf3SZcGOUQ6Vfm+a8WdPQBOPbg9E5g2E5MhApcBlF/Tf
mKjumAOnhCYHJn51DSSWPhSatxrmxvlfO0gDyGgC2lWqTvgvxkse/4Oyh1uMhz5bcC5Sv9ypP0rq
g2AVJ4/fikpM0gI/xx2oY7eRvaqvBs+4SnIGt0Po7OwGuUFdLF0Kug6vsp42+kbMhGAu5FQKK82f
eaDHnITyjlIAhFV8bl/i6WQdL+k+H6Y8e6T3QAbjPqtEuiQ7gZU7Nns+q9YnyFwPeb+9IB1AAy8f
Ki2uKg2Ji2LEMjAvPpDEaLFNhrgvAAKekFRBwnPpVmqLyIVOc8/D2O2DmQpva8/PiT3R1kxyCluA
x+Eo3zP2WrbAGr7uALe1C0M0/mc0RkEerNyVAtZ5tktWyGzI7OXb0Bu+7o6fBUQb0N6msJQ+cxP7
9BDMyvM/uTL/5mfWR3ElPGF3zNkQNOD/LubWw+Sn9AD0GLydCN1r32b/5ZGUUvU+ObBkw0JKn7cz
MBVgmXgbb0we45hRcCmGS4bTJ0AToFkr5ARcLL2a2rtaCzinVyLbpsyC+QbTVxut7nqdqdfQEdt1
lC+fxMnuX5z/lBR9UdG3FgjDVyksERYd8X8KpsTG72P/5DdHQPHAIJmIyQoktGBB+xny6ySPdDQh
O/U0kKJ2B5xwkeIgrD/+H/Bj+TqInmMG3eOfmLayfMJ3Uo1iklBF18AVkCaX7KSMVf8Hhj1m0EDS
WWK9qIHjstg+OdDhih96YRdO6Ql5LUAEg2i1vr5vefU33NjJK5ykCi1YddMmKluY/7lgaV5v0aYm
wAt1gvEKGB//2DAR02O5eNjwCjdStuBVp01Db7yUhoJivFZypNRKxSNdfqIRN5/hqPWehNqATQuk
H1/mprzGuXWY8+/KydnEiUqgrm0Ic19YYe5g62cMZcmaUHVn9CPl7D47OMgs4ul5iz9uOJX1pwD/
awPzCx+W4hoQ50GgftpxFVMEqnRUZ18IBubBNQ2DdYgXcibQjrEiQOmiIDGTH4DnPUN3lp1P8B9x
4F953apbfEyMwkT6FJqxoIA8HhOrOmfgMiJ+rD97br8uAcSeB158oBBPYBNCZYboUGWCuCEAzxSh
oqAPHNUe7nt4Nll8kBPRZt1dyhi2Nb3EYb+CGXbDruuScjmjGAv8svl4E/bCkEDhfw9SECyBRdFT
9cnWAPySqdMpfnL6J1WB3yET59ltJoyF+AVtCb+/eREodE6nlEUPoMU0vgBYAyki++Lk1+DOsmrq
0twXq5rxV17Oeisfko3/Wwb+owSsLL5vunObgUpoqHOYAl+03yHsQaFFSXS4pOTaQVwdIXvMJlPj
LQiNGZgixUY3xIX2NZeaw4IrrH6KN0M8Ruu+38vstiq4KG5gRHEsyanv6+lcVPIA9f3lqY8ZH8Ra
lG26hKuBHZ5w+LUBZKoVL1CcgPu9qQ1yZ2EAW2z03VYPLke7U3pSDzk4Oub5/AUlEoAZNopbL4CF
uWVQrvN+M0DfyYAhSz00GrCAbEr37L5eGRTqJQtB4bycPPvAtRla1u/paCF4NeIuyKn7M4gR41tY
blph5Kuxo1qrGpUgxWnYEbv3Pt7bcQs6PLlOTzDUaD6YzeMB9/WVi2fuUeF1KbQFL2HgdTOoPDs2
q50QShhi5o1QLvN6tgcQbeX5+xmbPeWHQTM6oAN8iJHlqJw/Os7q6m69/pTecZ+IbhDU88Zqt1o5
YwNkI15gaHWR1vHXczWxHxTijbuONTY5wuSVhP0JJvdHUpHGHyPyxvHnBWET0KyGkJ3vsPzkAc9y
Sv781sMwcmb4v6ldbMYkuKP4yS3fL2eP3RGD82SH7Vf+NxRlPVBD4GlXAcKQfTpN5UGzeJs9vQ4b
r16aspEg4bsqFEa6Xbg699693mP7FAYk3hunIg5QpO9XTylQjtXPuJWNQOJRP2ihTCNvFCeeMTMP
sQFSVgq3WTcnQ7WaoZ7AF4HwT4z5GWTdE/GsbM1E+X12PaKMecFx4tPs5yhGHSHGptqI0v2/SCMB
WG61NI80nZaZEWjkwOXu9G7DpyxjW/wD7luKG05pk2edL1/pYJfO8PPdFYA5XHAt+2CBF2yoFYzl
dVPO0nBRusjyBEc5sciT85R93kqc1fe+NC0YebKCUk4K49dE0sqwyJkCBhbRGefhc0Acyy6iGIQ5
wTg/uWQI2TfWTM/lv5GK0SYa0B5BAsG8DzI33Orb25ELKaFz0/hREU5S44vmiK2Ml742nkJ2ED+7
4gk8aLfoJynGBJRGaGITvPO0iq8enOFZQ7lYPtqqXT1ZSbOyQQAD92xydzS7xrWYlMfm+DVFGp8W
egGw4rXwCYvDdzB2igVIfFvy4NLQBFi6KXEqXmbLv7JrVGwHp2ahpjssjk2aO/+Im4ggebQQU55u
TgL9tnMn8eu136WHkLBLM07TXO1YCdbn8uN2qBjvROXhjw3OJJ/fPNvaQ2qJAwtuo42I/mdLgwwo
nyBhDDoOeGAn2w+6uuDuhg/lKdz5rkFkDctniYjLPzYNI1r+8ZcNPTeJdw5oR2CrhdlQSC0M3OGR
mX+cYyruzYAv/yMV7sgPAFT2qPkf3F3aIQi39OKyGTxB6Pqv1IQt6vNHicQlXxozdAoWoBV14FiC
lkaq3vvlS9r5yVmWP0obCO+6jreIwnxYvg/krQ8L893SlrLRvrL9jjTCfcnTKNQS/OSxgYbAWzx5
uVOrZcbFznI817pE2wdF62buHf5ud1fopxcgSg22NwrCYtXISnE4AyyhGfTnQ/uuxQI96nkSIbSr
RpKJTCUeQGDN4vUps/L1jyzX1nD6cODW+Os/MRD+8DC3DxJvZ/jK1F0BeU4Gp+PdQz85OviBRpFX
U0CjQTnd/McR3tVLK9mtqqMjrNZp/0NV1LXInvOCxfLr2KtLh4jJ3kxe3Abtjf1D5Y5rQPJUCCQL
tJBiPxnjZjv1PTLwNqt5jwOEDdLo+9mMsuZLdzDEhOtFdG56HLhC4W1Y4qsVmcTVUVHn2cx64dWU
VwFzFoTXhChqq1dSTdwCMC81A2ByPsWiB26+t34/fNiXfKHspO/XiSxYAi8j2pYbn8K5HVqctEoE
XU+tjJ4FJQIgfgTI8/cQsR6AhizCxFL8dKVX9KfeF6rB27JSSstxegZs60InIzOwqxtMUVVg86x4
3c1LY2OA59hwvkf28c0N7K3xIJmU0W6EvtmCc5g+jgFI74EMjndNP0I930KrVTcUK86aiA1YN98Q
KOO3uP/uFwhPqQKXT6igFCtVePVCjta5aQEaVzszI5T2Btz1XlgS0QMkzHQXT70COUNztRZ3ggcD
6EtNhxIP4SpUtmFNl23eA4PKw4HgF0sixRJXYabO2t+TPynp5ABQEjMCgaTw2xAa/FGOXeGE/1eg
nvc+n8XbOJUItgNoC5NWo5ObxerEiODC3iwwkklZRmZEdaQsvenaL/HaYMGnq/JDNp17FnHIfCMz
RfalBXiNMBrwQ/gPRBPYuxB4C2lk/V5J0mkv5ybEKqlSOl4wNhkeTVSCooMdxz9wX+Ugi5AlyfJD
4ZGhGxG4Xy7KYUE/MOfkwExYCPH4DwIzaHNx6CUl25kGkM9M8KOfm5DVHRtFhj7BrnV7ydk2ByZ8
Yft+NTHIZIdSx+l3DhpQ0La4zCO44/QxNgOOgdLkggnzjtSWCD3kCos1/3Ngps8erY/DxJC0H6Z2
NtvImtXLYVyhxl7OUpAkUdafeyIO8pFjIhlrzkbLq191ySK1nygFe80pUhVLMTMgjQ7cqjsaPqO6
5o37NBbgLrEoZGHuwDmWoYxfVHjIEVk6VI8Ir1J2XFuizGeytEzwI7HWOWqhoOVRkiMsenxMJCGy
l2LauwtcfvAEuh4GUzmTnc1gRF0mMINEKUf4aY2EVzVNPJlefDz4UtgxMY9usl+eAYvEnbLKNiz5
0/8+/Zw+dg9BrmzjrEBW29RaEaOt45zT2U2ux1Tk3z9PL5dN0oCpE5ko31eULxrL7QrMl4AP1H/Z
lNFOXEflFTXOyOaQ2S0GzKIUs9fR+fxY6gANf61KmffCp27yJbRrW+hBr+xBXCf8+k4tsIxPbSwC
1BbGax1SXLEshW2MPXuHliUdzv/Vvajsy5OligI9KmQ1e1J5LCPbQRW1ze3RAJiNq6CKMnlbiTjq
lPeTlHPz+ZzySGfq2rQ7Y4qt32CbaaZ3YEqxXfXRQ4AXg+zjKkIQ1XsSw2SOaiyrjzy1XWEb+S3H
7ZPs6B2gtA9/royGU7AHcmi66TcEkfmIyxJTzGc/a01+iWu029I11yq7tSPhQ/LX870xc7lyO6Pj
au2z6kQ0OCHstXYoSjU05hxoWuJzip0lTelUvndiVMegOPPH5hRMp99830HyER5Rx8KqjdzYuo8C
3WaNeMfV3d0V2ibjKg5e4Idu35Z64+gVH84EFPsvLqm9uT7JGUNeJyHPMtGX+FAyKvW4iRNI1nuV
quJW3VnqeHXHaQlezRy4zmL1ef3KERIdOtmL6S2u5aWKWu0yJxsU5jbgJz+2Wl0WTVS8rdBDGdmC
S48fC0/SzRTe7ZpFSzHnI07PqiK4pwSu5w6ePyEjaLgLua4J3tVxUFGTcVvxtJZPOmoU63hZ48en
QzhTYZybSLEcha7StsO7iUvSiSarMGyI+JI1SHQP+KNY8KlhkID7ZRI0m6mqxpEL4n1j+qmJSIyh
yZLV6GdVeCmKSoqH5GWMaA2OeZsbYOBUmkFHNbnXzgiouPDEF6jma2fn4sS0t7UeLD9+5frLm6lJ
X89wPNgUmjeumiFWVZUT7zTuJ1aC4G7Sr6lnAcl9XQ5PgoMqV7UnZUBCPz/J5I/q1TadpSJ/euBa
dV48GHtugEBAqc3WXgAu3363DSItH4MTGDUyKaGIImlp6Oj82UxE9du5xyapIuOLovt20gBqfr2a
LDhfNrCF8fO7bWiaIguUp6+fmZ1DgNzMd8ZflthKYPZWkYK5iYefAhXpPzSwV6blPVNdljI60o+A
5l/HQEbNQ68/ZTSBKO0RMVZkJiKmwUbeiYMBDDq76P6O/lhMpZyhl9juqcFuFlVI5DkG/2rW7ths
d/mpMsflcGTc+/uV3xU7ypq6/GDzNNqqKuYNfsdHnOLGfqspOGkVOjIGlX6QhDrYfwpdZDzn0gMj
6LJEwCCO22l0YDhW2RNDjx6DzPAyVvRtucdhYSMHJR96i1EeqWdAqJGOzc2bnwBtmyic5irHrmv3
cVx2RZPrAJVU5m6oonV8tzuC1NHoCIf9oLy5qOgy9+NYNYv6maq45Qdew/KOXEua6+RoJ6EauByu
VxXq0sY8OM5a81THALvgpFME0iLfzIqTKoxks2+Aibl/adkUIhalWC3V7Eqw06Yh22SwUeoa45UF
peTYAhB0PzIJtutYvi722O0PwbG1upb1Zy0hxZBbqtJHSZ7TydlxcUL2slrvUQQPl/ocWpUB3aYs
m7MT0or7m0av5NwZwhmc1aP5e8h3n6/UOX/cXBjt6Y1bHpqePOUWAuq0ww+TcDxcS5mI9OWFUrTv
AtlBNv4zYM4y1SaNN4SId9NtaH0x4oE5+mSvcfDk2UnR1AvCjM3ow0EWlsAsLcEiMKE090k3LEjb
mUSM1pph9sK90ldCGa54KJablGHr4v+gXzD+E2VrNPjtSDsRONbGJcNk4mNU9LtPotBUkbGWlg0k
ZBMtb4kFsOpDD/EsWZRO0iqpr9jqWISbCescJshlwOfIGeT1CK+QGIbLHsfOF5t1jjMcZKFdqHEM
GQNP2RkXqdgR9RPq1RfqWcZkhV8DUDwGvyxrQHAYdXq8uzDRN5W/j39CVPbIKc4UGsrLOzrnF4Ff
Q9ptqlkU/VlflXiGsoGBpL1bV51oPiB+c7J7k5//Mnp8qsaE+jlFeuF8wQXVRS8kE/icQuFiAH5n
fgn+7CqLYfEwsOrupd5CNaYBzq77JRC9Wer51MshQUI45Och+iEEIl0cOF3LxBqvSn4yz9aP9HO6
C6EE3RY2bAYX7A1NC8vntbikoFmhXaZCM1FqfMMgmp7sQpASbvCq0z4yDy2Zl099r7Qgw47zZF6A
Kd6nh2SBlh5eGHgt+tMk7g9l35gguV4j6/QU68N0MbaMGb2uS+ZZRVIXR3PAb/br4D7X7HvXu59O
KDyxqTxS9rN52qQ3QIGrGP5XPcJrwKjkpr6A+F4fgo7mmwXpoIcUcAdUHjHnPFRlc9NLaNO9LV47
mBFqBipZtO5dxxB6QpnVzYu4U1coNWZZt1HYVlvbiPorZoFZPVMl/m6hmttzMWZoY3wXrjSRe4kY
+XRxYlK5lGbUJ8p9P6gwSGJNXkyJz/AROL5ezi6zCWVlCJ9KRje1YwgFR78KoHKpEpI8UB+VtUEE
+8HtBpMxn8a+PIJsiMpF1Y4hXbsx6lLbn1qK7Qzqe02dk4QJ4X/lJHXDjmyQIVdckpJmpbgsgwTc
RA5lQb2uhuWkx7fXz+IiAZ2Gz158kr76uC1VCW4/GpI3FbIzL8dwsSicOYVm7O7U2MLHI5ucxLFS
HD9K/DIS7L1woTzELD+Qvqq49NdXP70caeq2Sonimjwp+3QBVxnwKkuSA/0PoQE8bWhql2JHdE/L
vquOLE4SGWZQXqvRQ69FUhgpInVe0U3exBpP5SocPPvajJjcAxpyJWY9hgAGv/1qvQaJQWWXf4r5
hiMlQvOww/BCes2lEykmokDlGsOYxVeGcXg9kb0SmiqmlW9jIq2JfN8ICOWo9MEBC142/3g1pULD
F+Petz+DkepJMZMAxYbx8zoGcDqmOLwL4+/ZtO2xiQX9ObAJfZ5h6HTQMHtNw5ISjWzxeeayce03
k+6K+sIE+D9i2OWgjEJ/+u9s2Mr82KmqJVoysD7oA24sqNRTMeeryZqbDEo5wamp4kgseA/OdNPQ
ZlmChl+YLq5WqeuGoDI4fBgdR2Fp2JibS1HZiBguLva2OrBoiw42Nylyw03uj2mMvz0Fw8Axfwak
No47n8g43OtRKGAA8i1gcTLkyxOAMK1uPXmCI1B8BDeB/UMTTeWDpf3bpE6gHZLcxbbADRyx0U9p
DC+ibkVr5+sBr2Fm3lG+Aiy1fJOmkBBHBMnHosKszSUSuEb113H66wfFUtAo+kpjZ1mhmRyn7nbM
sVd6iC8HdZcw2jeq7kUgSnFKDhCgxno1Wdl+1ntcUl7Cb6yvQrHCQuZGs+HwS3nMTz0xxof40nok
e7rlSPApQUAaF3LJQtVRcn0aF6vU4cXem+MbiWYJA/Nuzy3GWFxpZI3Ws4N7OcL91mD6Qtu7CiQR
M638tazBRHjSxBZIKXLmD2azqJostsVu0kq7a7GvK/70ErQdC+ycId4Pvn9Smn9P29w2KN1KnbB7
lY1SEmInfU/enVw19aRTZaAnY63/lCzfu08nKNlG0c1Ri15oFu0sj9FIsubHO0gooyIcR5KwT3mt
HoLz0A4l4KuUDy6oyht+xIYHsmfjEZGzEmlmgYkuOQQdQDip3oJGQepf7yXLGfyTgvsucj+VgtM0
4E5ZR0/zASzMAn7G3nougyfLN6k1l/Na+R9JbtaM12iRqZIJUyS1GIS+VCf4bOVainYVR83QibMl
GAa/hi09wIx6ASEgyLmmW1mvLnkgnmA8C8LCVFffTWgIX8IDCXeHAAmYo09Oqj6D5b+RHvk8TbZF
n0yTotBPlocR9LjpJYNEjlNlvTdMRUpwH2r9eXYFp5c/zuYNT744wMnF5PjowbgyVVcyf9pIiFvM
PuvqAMnt9FckrvVwag+6yZXuL8+88ZLrl0aaAe6fu7SNelCZy2HLXHcv3Ai4t813asAArATRrekc
7HXIy17HArxCEfT4VMszHUNZn2mhiflzfB8OHo7r4KdRHE7N9GstoIYIfKWi0WZl6zUOeia+iB2R
7BqCS8JfhF+4IBabRM0kkgYZ+R/teSP4MagODUkNVcZn1p8YsbFHBHhX6y4ZO7YyhhAnGwVqGl0i
pVlJq5UImm6ffwa1eLLs3cLYXf+wLJp1K8z4M/XCUDZXzLU2R4CK9zTlhdVNscWRDQ/lxkIC5GLC
HtqisA3L4/Zao6Hxsax4ens+WI4+Zrrvv2nBSbiGd4OcS3RGSS7T6oO/nHun+T7KEW6NVk19buvo
cjveto34YOpfT3ZNLtz/Fg3zklIU1RfXqlRWV/cetqev4xwBGxMw4FhaLPhXaZCG3X+DJdq89raf
du9CNwSP2F2hOr4FWeMMLr/3pIq4nzeKH6cT6FTIsfAtgasVIFAOjoH0/MHcZRa6g7oRoIkVyNyU
6PA67xE3asLw6J/8cUWI3bhjciMqpNmpJcpzE3ZybXSdfWdc2QOiyXT9caxs7vEWP8e3GxGgUSoo
ygTtSoOvg3ENEDk4oWkoQZ2y7Hz4SbCXxCEHT29vwyPxtySYA7JAa3CtdhXlrYdr4m5sdMwyZJex
9SXCogTVLdrTteNKvLpkENTI1TJzW7H9U+6sB9WdqSjOL7piOCrvZIMdumYJcRgA+EB1CRoy7nRu
6CT8UHKOPZiGvQuvAWInfx6Kw7Yj1WuN38bTyouy6giiP3/f+7n6uMBDdtp8BBJkzF2jdK4e5BbG
dQKbD+R65ZxxvNQct7/DVjw38JD4fff/Z47ElDMdd5NQrkxy+SznavFz7BfVQZm4HmiCyNNW+Aez
lYzvyP0rB3Ogb0jzDn2MVhcWuZHHl10hTjfqKJSbjqfk1/xMlHCIMiSdDPAsPPRrfQAkJcvP1xe5
Ifa+dOZsSs+eeJenlOScBUD+J/xiRnT2Gw+QX7bsM5VRhiWd31n0eQslqkpzmwQoccvZ4m3LQQRc
ua7m+4lvU4hOyP4Fu3Di4OQPWfO1MLdkvxpWOuBalngVBLE4QfwhGP8NIKMc8CvP0cyHTktYoECw
DWGqRSF8n/cZHn+z4yMOId10yts8XXCrLS+XVVngVXP6VcBneS/N5RjnIBXrzWlUe2XS3/ggVa49
1VVbuy5XCMEMZoNCi5MPO7PQI/Svofu0eKipbgMuB+rASSLZIx41n61CqhdduK40611ROKkCg+3d
AdDaSe4W3/NSITHH0YeIk3fiJd2RqSribS5/H7nsRCW6+pJ7sFogOrbiO1y1H/kglwxjgaOIiss7
fQhmArZ9ZePvlvw1lPMcUuTWevu0eu8VdfH3TP9H8jLEYyZtB19cvRyq/P7iLx+N9Nh8S3egnUHR
ReJ39YbsXt3lI6tujDuDCuL4j1oYsaXPtHtzzcmlHPQJs92xVHRpBRin+VeaApaL92aHWbwp5Dxx
odOjvbtmsIyxFoHqoYh0RIT5SVtro0PayzgY9Nt82YJ4rIJZFo/qbKzhcACGl18Dy1x2KCIeu286
mvTuvaongQUUnBKspwz1llww6TlX7KQ2aLRtb4Gbx688zJLHaix9TMizEmykdXGBcKipIjcAeFnW
Ts8wfqoe7IltfLbuqJlRjAnuIEODdEH1WcLn8/Vv/SJpj0uUJE7yStFUqzOTS/Y8mqYVk4nhJOU0
XrefSwy5eotT3cf42w+rF81w2ZGXxrKfyJVRSl2loyqfRnfGqQxqicehYf+LZoutFHSGNwNtdFwO
DPsFEtcVwZKeTcxDj2yFHX660VEccS6DSvjqUpJe6awbfudszsbe7eWMhjAMv0K+lrVnCV9v4AAB
r/cvoWeyp9eZAJoS725uvSERgDl+veOgbBKmJ7Z6SisAnSAD5INeDykBY8IXjlIydxaKOY/B+cPX
qwjgx7VO1eN8NlqSRyrEzcQc/BtgPNUTQRnB6u1VrLd27tu0Bz+47Dry2sKsC5DbdiHyxdLbRs7F
TX0+2jSAGPEZLV6hu00cNGnVqVDEP+mY4I/7cCpOrpCr0yEiFNr+kqBDQEKus2KJH73GG0fXsZxb
ySoxxYzHZNtipCFpE7+OdlFYIZb/DIEhAKSc1Mj2Q6w80i0CXpuhuSiSZrkVc6QLVg9BUEXX0wfk
WTwUJyE7EUpGrHk7dmoibpUPRAG4Q5kSQCPjhNMekKv+lxCx6EBQcc7gfSpovCexojUybrzXg0E3
AYTU7XPLswEhFaspzBbXoSOtmZ2+rXZCJ+grZ/2pFOZvY9VnNewOrfJzOgbC+MRW31IxFBBJWFBJ
V+yXCGldbGx08iioEzPhuY0m5Q9rPntOjQ2+J0JaSDIX7i2j+sWLOj8nP0nM88zMwtqZlSK9Ddm2
UKM13sN/Jdlkfomd1BVeEs9xEvWE6990DN49FA6pdP7CdcY/eDtbf/NOkPO09NBlLDysL3fZn0Vb
TgVscsBRAueRH3kbCcrjxdKS1RMJ2xmfxR9DZGxHPfiU/1mM++c01ozL2NDwUO/yimjx6gdgsfhJ
PE02hqDcGpLgG4uNdTOLPForQUZgK/zGG9j6lUGcDZbp42MncEgHG4AXzOCCFh6TD2p+pfm8jNnD
svY9gMSPbU2yOux6aIZrv958/4zs70u4iJo1pZpWyBLWfAIruCqerLQ6AthGUeIhm0gaLU7jhMCa
15IREnkRlg7+At4SnPiM0l31gmj9xaBQsuo0OPNA3zEL2iBXjGID1fypphclL2+xgyJ68H8TlzEb
f5Frt1yzLqvFIN0bj9FR0d65igoV5NQWC61C/DDzwMU2olK27BPp9EjNjyAEYeZhwUTtBAY54qSN
zXQvN0UA6ZIt4aEv0QRHuXtABaC19TdGGSrEUpSfXhd21MEQlSI9mMZBgL/ZY+60wAnd3VXN9bFK
GJf9U837iwy9cbIizkxjI5zz0CdRZEGiRJkjdRip0xG0TQm0sJlO4BVdSPqDYK66l4/09+4KWY41
kmAlytoykqX8GyWhr/j2g6AaWDywhzIuTpLGufvZ+Bn8TApBNS3korqv4stFFFZeAXmP58xGxmMd
iaLRHxi82dnRAlrC8lh1pYgFGrbhzBqHaU4iT7iEFDwwtVlRIbS2/YTeC+VWf3bqMDOxO9uLk8Iv
RxqIuo1RfqkFYj2OPnjn1oXAxHOIhR4zgDyaPjXONwI4mIP+U73NHvxhk39/cUP2QLNEDmysY8Fk
Dl7axjzPdzjZ4++MVVQa6GsFv8VKAn4JRCsUL575FSn0V7Dp32EDYkYeHzZKHibxUkI6MH4ZHPH6
o4b3PkcFpqdhdKCl6Q6WMQ1U/UTHqOsDPow0WR6vvh+m/ElbuXi8UYeZ/N6Ys6Zwz9teOxFGWeS9
v16rugM0qaPLmXPrET84WGQ+rJsr4s93Q63un35v4u8Lpkk0hpjqoyjxuW8VybCBptI2UM3K//85
bnLX4MEuIc9XE8E4pJ/GAJ6fNVYh/M8mDeCkx9J9BTv8fu7GgFymi4HhwCgXex9IZUkzIvn1zqrF
9nnpEGBRMp1FmKWtbcPT6uG5ds54bXnB1xZTju28ulXQZusQVn8SIwrC5PlUsC/CwZcO7SOrkSaZ
noUYCbR75jgLIumhY9e9NxkW/7IVpXVf8Pt0voXovgMavbwFRRkb5G7im63TV0MdGY6QfbAYHBEz
6YcP+RSMYJn3ZQUeIiIvApz1mihmAB1HUzFXlJiYHKW4Kedsw5bR7+DwdG9altKsNSRN/4pWwzZR
4uz8z84c3VYiOvgxyJhUaIXHyGaXMBRLH/ucTljuX07c4hRlYpVOdkHwjqlWIgdktuwVchUU/uPI
N6Vn1Sepo+9RqCbLm5iN+Eh/r5PEbDErOhb/oc3q4RErS46VU2HX9i+U3odl1JwYHUT9IgFTwS39
aeD/UKwsoDe8H6to1ySwuLwUBur7GcjyUnpIg9knB65pQDtAUXVzZmOGsi5zVfiiGhOzIl9yhyYW
zqJaK5ITFh56wv7TrbA2VW9lzOBKHVSPm2ckDSxbUhU+4VMm12Hzd/gHP6QK6iXg2XjCz0XyB7cC
vyGiBiU/AZwJZZ1r2lHunlkh1AwM87NBWRHhaeQtjLOF+CP2YjyKn6TtgPcf7LRr28HKp9+l2ITl
LjxOlVZLw8tSbfIZaF+exLFPd7KU5ENIrGqfgOUv+o++wWicD8egx8CK2QInrQVVkjAslgd5RLfL
AM+SoEJLQUASLubzJp1u0ZAW2qNT1e+TNMMKlcEpOVRjT5VdFIHcKW4r0hRXOIhlKq/GgbyCZLQ/
149IuQ6nV6SA4WHmJQGCl9NiL89rKccQ34OuBbF9oVDLZOuo2DQIvDGR4Os8qEz+G7Dz2cG1VYXv
llLJ2/K4pICqeZM9hjaCeii8fJJXSQWA0jOJ3rQaNNJO/cAn6fWYAQqjqGX8uN+OQ+XhLZwvMKcB
XUjqCji4DzuLvMBvRLjzrkHf77Vre1ggxXMO932NHX2Te97XEvKqK7yW07K3bSNmAUxjqyuYYUB0
MkC57ZG+ea9G7iT6+z01654rJ95ODcGROCfuhoNtae2Y2CYxqtBNO8Km6HBteWPUOlsugoromP3y
DsSosrd1y781oqzAMpC87hDNm76OQ4cdjwjpCuYmq24lG/T4yW+4Hpm4FMuU3drqJ8WffmT0CgQJ
94jPySmVtZGqHGotfS4WWtvyCmiY/T0cWyrmSdX5gNp+FgT178t6VpoyanFnZEoxzjctiZML06tn
L/vkixvmXiO64aAKuImbDlsBbW819mD4y9JwijfUgi6wCddRaDfVNfU7eat4Ae+yiDHzNZZkaWQl
cByt/KtK8MABNLJEIjFxdSqOvNqH/cQslR3ViRisI/lUDPn+pA0YlSUGmW0CYP60d3tQ2y3JFf8r
5mLK4xFuWO39iyH12Jkz2ULx8PNGj3KU+4uw/MyQtz2FrdNhf2uN4toPCclysDhTAljxIhwKusVw
wU98vWqyfc+DtwhfuXHFSs2ETbq4plKWuMTRhCWSw17VFDgmdLWP8pwwtOrF4a04vUekH7xHqEyB
j8vqemaROGj2X5I5Bp2H0PCygyrdMOSXEQBaNKMN+6VQooJbF8KawKn2bm4JujaZ9UKB5DyTopWd
2yNuqwcyLWOBg3CuwnbzbgwtOC+ZlnX3rt6TtqL0/sHQKUrnOR3Bp4n3SIhiSbkaY4lVl8r2rLK2
svv6DC3J9DrKpP/bEtROw+j1FUuFtAeXzquqLDb76yAmIB2AX6OFJv0QhHpov796QcyDPEdSxhvc
poR28pLPkd3RtaPOQkh1fr68dXXCUEeZRWeEH/l2EAbWApQUYCBg+clpEOvTIbixeraEXQrgu6/Q
b1vFpqUtfBKLHVxwptGu8qqXuVcgVWV8y+oNAehWTgN6etT3ggM8Te2nGWVp7X0CQs2p96O0eNf5
Rrbig/awSDV1ByxqfWF0V6tSBND5kDJivPGNtacdV0KTk0oK9JimNQpnnVEONFNucRL0OBN9RsMQ
8Rj2MTO/dbrgb4djiB7SCZ5VlNwGtk6PJ130wTpZiXKIjjGbmFFdgCEIxGDto7AaybGzZ5dyaOIn
zTTom+6ziNHBaNweHGRZYEdgjoghZh8CwZuLNefejL8IW96X98MoKW0zz/Tpe9zadvLFaZQfkyvE
gOdCBZjsYWtvP0+POJn92poiOH31JSLAWjmVRdanuuf1s4NvjZ01bvFwxSzdSZur26sjtoK0Mu3X
8KnH5GtHuLdnxfzHCqTwrV1FryW3iNCqIfj5qlxWVLAf4a4NN+UdT/OT6eQU4WTuTabWyrF87I9h
pbRWVjFBP4Y91NtroHI6acJZgy1fRm6CXO+6nlfiOxlms+ZIZIe+ww6L88lCkywgqDNAgTwI5LON
mZYJ3qbDJDhMliaZCt8sPhpSKT2uCjipzwygbgEVCUROMPXXXAxc2upP+SJFFJJLIveeo0Xtsk+i
ZMkJsEy0q0cH9Adbq4rJST3PkiNnfEE+h6DNMrvRODHoR+D0bhWOKrBdfaiOvIAsM+sX+7lH510s
0HrT3bctWXtilU5tyccwNt18A2XUl/BDnPjaHRtX245+HmoT4DzS4GiflnBRnJX7nG3xDxkKbKlT
rV1LH0uMAd9vry7VU/0KNfSpWuqZeARfo7b/+qfeKsyFUbPhtWgil2ZMqCAopXa28ozVX+P3I6Iy
rqCQ6SqlQYh9RwH684QUITyq5x77V95e8Im43woF7pSV2c9QAWwT+qtG4zYPKdppPM51wJFowkGx
NUt9HqEmPr4ks/+KPkTryHakHAH3voWO5Pzj1q85JX42PaPHVF212Fi9GbaScTWiD1yTKmu/vPSL
de8T5lMDUqm5qRf75ONc+42iDSM8BJyj34fWBwMoRjVLbZ5JVo/JoAQYW3WCW4nNsEHCljus/XL5
6zptwyukiEyYQ9pcIiABaCcYMX4b4JnqgYvCP0tyutE+y44T6cdtNwhdKyu8HQvGIVd64vd58whW
W71ntwAbVl7hHVcPZFjZEWnRqDLc9FzafSl7tqvlB58PLo0RbAIwM+QSxWEloMPfGs757J5pDr20
YDm8gW7JtmrYbZCP3p6ulnwAEEuKAyk6IRt3BCxthrh5sArydmH42ikzgMpOD9mcA/lmTctXWeBk
DKAXYRDD35cQTREiau5pidDTgJim4yI+08HCZfT7XFdKr9ntHYfxrgmQiHSEI+JHMLBeACbzAaA9
0iOXGL8nvgWbG59sA8wHVSiREwX11OouHc6stlhhZgT9iyK7bOGc1xVj4s3g7oFmVtn/h0dpkpWq
kvPGIp+5rv32ANDkTN8MA8sQZfYRJiDiihytZiS8neW+c6RM/7cUQIqh6L5VqCNBa5brSkjbFNWH
E2mzPU5JNuXzjMJTEW/keFFMJO0QtbA8KpmQZPGJ7r8vzVitIzsF50n2hpU3tqTwPJdLVuFNovTC
NLBY2KZtMQ2M4LeGY8QYrPMFibMvjpRy17fqgML3KBNj16GX6PoeAvTeokuPaQVy3tmeCpGEsUX3
JvRwj2IFjVPA1mtHySlf5TB6a5ShIG7LUobr1DRoJrG6kDsRKhANRZrilSoC3RJZGNPO3NJpjgbL
O4Esaw4qdNjQrfVWul+z3Y9wIi15PbCcUBHAmNBYIbEBkoyb0R7rVFDntQKfMQ2aJeEc0JLA/Bwo
D8/W8B8JYnbEosgFLitMFd70Yz+lkCB9kCgNkqB1i/VNCYnLOMNwXgn33x34Vq22ERX9JbQ/rH6X
2EFhrWZ/AsXV9O9t9r36he3NfxJCoUOjEj3NQhXEUzARbJS8ecMAliibxEOTG+xjdEWZ6djs1aAL
MFVwzEThdP2Slgqw0qs68uOltbbyU+yHZjR+gca8INvE4h1zw+rGktIj+P+jcBF25mpjJi4qDKvY
5nsYCsqCb5RnRtnnKPcWtbJuVjcFEgJPTXA+8WfQ4e0l15bk9/tTAffrCR1O2v2rM+F9R2YbsIli
XcNvzA2UdzerqWa0ZE0Xh+V8hJdFpm1LIhb4zIl9HSYn4Bi2ovzNGgCK1XWGpf2H/+jrGZB5saag
tfxWnTntzTe8rNGVRNqkK6gFEOr65v3rYRGHJgU8vNSpoxHEOsEPg8y/9BNPLeGUeEqq9vRp/GkM
6+lUnPipH+Fj5V0qSfO22EAel5BZepClbs0DtwrQOOKJG6KgNCxYXUPKTZKT/T9tCyf1M5CAWyx/
2wTMDeCHJB/WRisetfsCwGcs7daEqAmYyiUoImbeRRXqkoDjVTql1UWrBuoscwPg+clnY/b6s65J
EoBT5ydVuLYJwxvQcavB+Gk5kGy+OX/LS2+rdP1cRr2E2P6lkWwUKa9eSttyn1iwtE/V4EHRJLhW
V+JTZoRKrVQ6jOfISjUzS3YC8ET2WfrQRdOvvEHzpSqtHU3+UEX7l++BRkCg9XVNODpeWuq+v6jR
qaPtbs57c9gTmqfJc6/PnklelVnpD5gK4sWJQXdpkxn65aGgp/mEQAK3lV+M3EodmP+PdBxJhs2S
8WcxnSYinw+HPcIZoZWHL+qxiwgvVd/MP6SYHAYLN7G6FffFOphPlhPOYJgtPvyY9HM+z6bPsPuQ
DkWbfjjYpTcABJI4wwo8wQHgOnQkqLzWoL+q0ChB8c+rExSDCDEvQRmsqU+XJq25jteAv9fYVAsL
EXPy+EJ28Qa1n89bZfD4GqdXA+XT+iNK76d5swvgn3ftE3B7edJ9oRYtTt17DKEMQyt/ZnbOrego
ckVjqyyLoXDB4vfcv9kv1z0Pz0yreArdhX76Bv5cThCH+tfQNI7T2M4mkfSbL0126R/mayUKug62
2zFSXJX+4DwQNmHKgSm77Knba6rM5eyCqitJ8Lt85vZ0yGQHSOYpmACAHNdUBHotXvUL9iEui8nx
jFwnoGepc/YmHRI34ZHQpYN3JicA+6m1xoqZtXmj/jQpxJyZqMlLJjOabuwMYRUbSZMC5buvYlhu
+nNPRx/AJgqJY4+VJC8atuisHQ1+DIYSRpoviA/Hp5+9QD6mkNTaxGb/16Kzz5YAiQ76FUOw8NjO
COkmjCFvkPwwQs4tJL1/FL/JLRkPAuu/RHAneEuJiGTzn4vE+hxbvmWWphzkiHSIq8/D1kLn+BC5
VPHMGfI6vG7a6XgnCS2lK6Znrt+UqPT9pHAsfOxxjxW+p5NntyIrHJtO02nH8eq22CzG7wEHtsq3
fqHulBiggaB/nbpguYMyH5HuVfGzDT6kTnIH4RAefg5eQs8rcG/WeR4KrH4koRQKAJVIXJ4NCWpo
4M3liWUx8k0YjJfnR8CRKW1VUHDqchDCT32EPf7ENG6NlLAe/CeRrhNF8aKF0NNUb6faUHwbjvmF
dwirDLtQy4RA1FZgEb2tASN/whai4ER92K+iCxYhdpe0uDBz9eOJfqVQT21L/ZqclZ7Mab5UiudA
M4Mk1RrYlp7J0UTaDGb1b7MitJzN9SdRwIhIgEi8QpQzjAsJfFScjYR7FwzNsnIjdluotODNWmyE
FwYkXa2Z9moIGnpZSHD32N3Ale6hPJgBBuy0YAaInrvuUGLecOB54LA23tOQ3DFo82BC2CPsbgjG
NvwdqBaTdItpgoeE0fYElvDq/Em1QUe0r91IlTwBkA5yuUCnKCX4cxF5Gurko4NbricpNKnIsSRn
rWELsQ999w9nJCVCfGCtudlWtRx7hswxwpjboe3hmeOCcPpI6Pa1w9frvC5INv1kn3Y+Baupo2LX
HrBYYjdOtJehKP6K9RLcWGCWwXy9Gw2dQ9fdXvVfV+0G5E6cgUYu+opCYBemsxZ2IEYKWPeoP+nE
LufXxQfIL4ao8EJEHjw76E6qy1ANbF+V/K40TcAaw5lYomPBWOeAJDIlygv94EJ6r+KBcw6EzS1v
B1uWJSeWHLCYkXvlt4jKqNF6P99hsN6UuNS5DDCRuzd9oDyvWO5CMAQJVJttt5Z30vsdjYKxYJ2C
H0KXEjJNn/eXeWnijgNrpgbv6a+xyjYUtA9cOG6M11tWQoTeirIct2zlaPwEo7TUR4ZZ4AxIi78O
snoEz3G9Uaw7N/+1NaN+N++zHvjIqdPqWIb3srhYhmT81VoDj5tBv1K+5Xz4l/Zo4G4At1P5fdca
+mnp1Mrfu/8tPuxl69Ro6DHu3EHVh0DzV22e86SJ/rZRmZZRSK+fK+OpuXEeT6F/eq0d8oX7ybPV
pvN3+Y4C9PuLf4HNRqLOXMD+W6ouirT63HbvRzaLxLckqmiHjflI64gDx683JDXcR1qm8GotAmO9
CAxXhrYElxzUh5BgHa/4FHhSDX3BHuzjjM38eRBaFpj3ossYkeNu2Zrp0j5gApake5iDFljasDdr
avixKTNPjxIwQkpe3xfXygMQ5i6Mg+p9II32B2CUhm9kjdOj93Tj4RLWAjAkyRts4mJFNsod4ceK
oHwHKuE+PbMO99/0lTyEQ4GefSVAkw/spMWf+YBzfYksQQLCKtzYhQe2QTXn4PBpg2QzDINmwsqr
JAy3DjQaI7Fboz7iVuhw8IKxtYa6IUKgWzeonoU1DpBUcMgTXDlytKExKdy4ssqKxOZwlxTpNOkb
38zEYVZ2TJOcISSavAfDblp0bPtZ8RsPpH62mWXUiA5oD8V8KfyzwDqyHh/KeJlHG3bTFnLFCl5w
PzecOGEKDZnqRSuPs/3k6zeleihzsWgg9RAaz8WTlhdMwmeQf8X/SRCHyqgp618k/W5BVsuM9YhH
uGdKpFWDgd+RAEHmqjoxISzQKH9sEeIW7RlYOfpeLkWjjNyhJYGqGIpMfSeXGoZOFgAnWj0E8OHA
df/QvhxOnt5F9Ovt3SxPIlbzS38bSax2STIb8CroW/8rlPBJVKZhwiB8vMGKmvp4zh5G4Ci2CYNp
NgIqt7wEASpOkfDwyoDfPUPnxUJo3idti/YpTsXvSFzmtlH0lfsnLP4jz2sC7oOXOD+JXXXsrLvp
TK+TqWQ7N7e3yupcMD2PX2BEKS68tVUuwQLe0zG1OsyJKN115PDKcKxsb2KUDLYXaYzpNE0oe91m
mfiTV1hqKQQJWjwRB1A/2kEMdn3E9CVb9SOrgGIKIJdGHgXnUXRxaCEC5b/lcQWdra8WRN0RFwP0
O/9BKRsu5FkkyE51G8pgtaOMMpR1gnGxF/z7gR1ENXI1dw1653BhMm4yCIwgJyvv8O46x4AJxJ6Z
SZ7q34/qzt61RVUtLVvSqW9ehF6EHsL9CdmQftfiNpwfJpf0XDjXuBv1XrBB+mJGPJK+rlM13Lr7
Mqh7FqDvEBTp95kaUC8JMop4wCRSULmIOihKAiEPXx8vz9O580DFb30yugkISPht2VVnGhOuwA7B
x0bxYje1KlpnaNyebPjmqJik9NKwW/yCOuebbDftu2ydiznGaRRJh8wnJKrJvHUS/wOo0RBTK7FS
dux671JsAlz0Oc7mnaedqW2EGIptoV+INd/2d3Yt0QIgpRLCz59UmhEVmETQizr0Q3acloq/HZT5
uWYoE6Ha+qgjhpYcriBesTA2RYO8Vp9IXH9KH6Wc/JbTIW0s05ZYMPcIk8SiRM9pzSlWvs1Dwv7s
bjhogJ5tV9hibRDtjKWADdURoS3Fe8l32OYY+GmqMmtLtX+VLUjus6IeMaYy/PJCCj7rRjj7922Z
O6o+slrOMe9sthNIM3VX7sHgf3AGIanTMVFZ7/7ZBNkzPJqv1YL+2qNq2WzTDfF0QmQXkqACkKef
NuzCUQaYJ/6jfjX0/jIZWLgBW9Etx7PAEyG7XSXwpK542qCrvroPqR/xLvh1Q/Ouyr7sSKbDzbku
8WIfure0zSPPpwuqFU1bfHYTpQZ7Shs2OB1Gs9OJs4DBg6JiYjjzWYLVwTKlwT5hyeerULnDAXFB
rTOfdrMCGTpl6WQQX/dGiB4+ycl+IhTiyEpeCnVhkq8/0MS8wczfDW0g+jQLfQAtDEJD9Gqzl+RW
QTQXzl15/t/K+gAyqg2900d9ZenOYiQQrwJcuRmC+CjGT15Vascn4VA21ZgaS5UOSFkjqhQmEVOr
8mABGv9Xp+M/SnWwMs8tB+wH7t+bm1akko8YUEnu3zYsFE5G1x/WIa/GiVwXeEOVIW9qPpp0033t
SGVRy1GfzFo4TUrDwkt7iO2eOfSmLUk68y0+gyGgjucNLVoOtG5A6nMcTAOa0SKIR6lZTS/ewssR
S5Fj/o26wIRoBTT2+5iYdEv/6G82otwnZw0PR9XzJMQNBIffhRVrLtiyxgVxGAjIJCWb3NHfx4CW
NATTIzaCLHtdG5POKb3axxFqJw2ZSp+hdS5uTeU/saeS8TfT6gUHtTd3tF6SpLC0t3LUi3q9We5Y
/oqsCZkHuyA44Rg7Rt4paPjSt1L4r0T7dkBwWX4xYHEBZPjMx7Z5CFi/db13pd8VhtOwdMDYi6DB
anwYHVpUWmo+7bErSGAhwhx5ImPxyVT3Fv9z4xwmpaOfiWKJouV3cGna54USYG15KlNLynu53U2u
/spHNyt6NXZ4UpdSqFTkOPTTUMNOypuQj3jT1SvhiLdVqSLU9co8yRM9f3t5hFFOW8x4Yj4G02V8
WywihAmJf3iGutVCNtdOJQljfqAIZIcF3PMXNZMP4X9LGuLxHZ72VcrP9S6uRu/OW230e65rB3wq
NGG2TR5DPKRSGn09YmmkfKnLdxcwVBpHObqWOBYrc9GQGrRWfYigWNdnOlAwHkWGomL50ZlIqi5w
72hM5Ecc09KD8fZWKZ6GblsHwi8OV4e/DJ2I34HT4R/scFjTN2TGug7WwjDLHgD5IPU5h7Hgv6yf
nYkPViotoz2NMGnTWYyqOaxrfLjNhw6mAPOepkJN3J8+9VzXzxDiwMIKseJGP3mcmPpPUrHBTVs4
l5/32B4ur68tZRZrI/hX75yZOyQOIZh9ZPWTKrWqoV5hzxSHv8kM0/rqOIpJZtv/2b2k8FaGeogM
/rfMcheE+Aa22M4sNbo7DxfAI5IukXLaGD2cI6Pr00aw/aNXVxcTAkpqnG9MobKYrcG+T7HoI8qc
d5kAvBFLJUE1zZ4SSJIuTkHDuJr72M/Gp0gkefBcN8bwwl/+ZjJDKgJOVR99cqCpVPxxmBMVqA//
HrBeOa5rcmqImzdnwu9U6EuX0Xzdf8ezUJW2bxc9SWAqhqjf/71R37rA4kWMOfmMC0mwoDpTu+tx
DWy21mY75e4gwxCoTaJUneKTC66V+/uHX/lH6++XhRizA2CZRuUjzc5nRdJKFf6UoXBs2vdkQefE
P99LQuBbgKxaHLgs8naNQkZ5nN+ob+Pg9MOz4kFyaf5V8TAPdgR4UCx40P7s+KIKTp+uhzVDpMO+
pT924llkMTqj5qFIYYxksNm86Ksi21YWSnMqYr9nkZP/y31gaOMmgK5DNMkZnCs+JUdmegtaNK7/
dYETjMLYS2569GOJzAPjXgq6ftldkQosafgn7lpjzgr9ou7rXKyNPXMqv1b6dAQGWKbezT9w5FnQ
hdhPj4jSAL1uvD6SjfBpiIK37trp/+e7Bs8eKd5JbSu6pVWFjfQ/B9xFdj1TWmu9HuLqj1QU9hHo
W5tfTav9/XLBDvN3S7EOlpqZrv9ymgl0VPhKXlBg1mzk6nr4BLy+40Gb/KsM58t83cOM/ONFHeqC
NPWn4hef9g0rZD96nlYQJVIGia7NcNpvfA5WA3tpKvPIPQ5wyZVPAnuzk+Bfxp8HRPQXRrpKV206
W4JqHl2qhWsxsf+tjVzlKVCPwWrhrFZluHzXDn7Kl5UOjvkftTDL8rnxFquuLVY49x7qsZ2NbaDS
5ZAdGzLHJNIjmRncaKUz3jLRwBMNGSzw5fsqdUOnHchl7EbMsDFSKiVZiObt94j/9PiE/wEzoA82
rdmwa1q0G5QsrUImZsLyAgKEdJMTWuwbSUSfVM8xD2+IoF7XKa5ujHcLgvfVACuOIFNyxVLwqoV0
MallfE92YJsXhbB1yF2OwFIAW6+w6p0FopZRM6aRa5skybw28Ugfx0P1J3QFr7VrD3IwiefOU1Em
4VjJN3id8bbjQywWDJsZKpGvVTmn9hZGIho5Tk8NRBUgV5q9RYaT963nfFENIbS6b+sUtdbvcZZa
9ZorPhPmJM15AxC7wOX8XARyoei10TPQXT8OcEDGESqs/cdaTv0Q6fCrMYWaXy561QyuoIdpBpLa
DXrAowZvTuBiWoWEwVLtxI83mPujhyf0rL2T4G0QQUzQRhISY/6hIavJIzRr3nnZ+fce+eckdyJe
NOI3Uw6iWlr7AvC76V8XfXuF82bEqdxaToBXqjw/e1IcObvVwTJPEd2mFygIDb/Byeoh34UXlPij
U8uO6TI+OUxmir48NJPxvvSZXa3WA31590zGy93boOdOoCwXoae0EPNfGCZ5qQyKr/i4aehEZa81
FBwIqU2HF/QXh1NPzehIOuOLy+l1ZISHZIvB+wFdP123pkWBaHmWJLnTdGhjaj94yge1+Xqo+pmw
sL/bt3gm5d3AhgEyj3xi1cyfTjKCkHnaj/4kctnSpn4jRs1Tmdbh5Wi6aBWERQAhhE8rZw1YUxkV
zyA9lWd3uuJ9j0ClkQ2UFNps5vgRDRhzvKbSXUy0UO4NhdmViKbKMM5bijq2wliRT9HwAyayZqSn
W8k+VygeDlbYKyOggsiTlVPZR7F5wDN2Dbn/9mPZjjg6B+luEVodXxDr5/X8XwKx8I3u7q39ndll
o4CK5CHkcTj88npwMHsAhcBM6thOE8iG57Vhym+HRlAYqCe4NAba2h/h5/8EHFMeHepQ1xauaqCK
ZgAA/lwLuxJVt/hiiDa3JkmEU6GX3gNJ+dBAMX9uQCtYOzrZF2485ut44yg2KUubrnJ1yfjX6dP4
Tg7vu7ZPNU1E9ddcBSJJ60PcMLdNrI0JT6itKW0HC4hOGiWUaGN4o5gCeKwIoK1sHqurEKjodkUp
BdaG0UFAy0pRlwTZuK/GosL9+ewNH9/Laim+5tHq+o9hEWbO0e5u9dFQedU96hg2uhbYaP8Y3OXn
n36hdFRSQUQvEuX9NgjWBjtfSgTK2AoLx/V07dbnyh3B0h5y/wGauvDkciJul/t7D64WZNYKuzLr
otYLyEd1GCHMQpq/2S7PG40TcgcNOBw41K6eS9dsoBgi5glVQUiS5gTdiWadPcyuMQ6YOTqF1nAY
9mPLNi0ypk9jJY7vUUMBQ8EoU2KBlYq3zXjxZGLvz76iXq8gt4fqfMjJoi32wzLKLRYFT0G8ntba
vI11s+TzRbtXLG5xHQPbuVZUHXotKmO0JFzOlvMNLKaHxx/PMqFgFKrE31S1fT0SMFkLEGwDro4y
BXMdoiY9Jo9t+xn6t6BV9uZJ4gPjlDpNn2AUF53HvOOLpfRc4M6FeHJZdgND7ydAZ/ckhp3PSQBL
pbSXC5+2K3me8q8ZMQ1++OzLs7YZI7pRo3OkZFmHKXRHwAA29jQeGAr4qnLkWIatQflf0DhQi7tc
532/63uv64ObI2oFswayBLmrVTMl9SN9yAZ3cSejeU+caoLqDVFJ5bGOchlxJhxsnb/9Jn5P4NEk
RdBb21HCfN9AbDPaz4o73xXyX/qqaPMlXWDckdzUpl49lPIISumHlAC0sTZEB/lqbZDxME3jzSZI
RFV1gonSB8FTQCaSo96fwPqxioH3+MBuHK3iN8FfZt4+OIdEgVyikpYIodUL7ZGF91xCKHiKLbQH
qoWGkWd0jegfkwJVuviNSJbPFOdhaElpBROSUcgPRLmfJoyYohlLhKImFxmdz4XP0mx7u3Dmh7Ca
6TRMfeJAcjLDres2crOAMSs7iWLxeTe6N1l8iaWFojbSd3xtqSU7rn6Kt0s1qW7b8PGIIV2hS7sJ
uWmO8zDAAfl3ZM7RyO+i6eoMMewZPBKifYcuHIAazDxBJZEyFK5qNxmTUCWe5itDYnh/WcBYkozn
6BWwXD7xV+rHm7d9yrelZC/lU8GaPChNDElgUoFp/lPznOEyfYighZmf5Zfm7sHTqSEogXnJv+3g
sIoKHMQRXCKp0apD2GAoJHrGn4g8Di1kh8FjnOvr5ZGPNfIh0LB5uJ7a8YSKi11VbLpcUExG3HJ3
OX98d2Ue69rLUeonKEbPJTXMq2qaVfSe1gONziqVzxn6reVvRuv03dUP+qRtrXVzQ9Hr1S1fBh65
gL0N6vonwlJf24uj+lBU7/SmPcjqtqFcLRIFpFJ09TzL6OV6jH/hHCRH041kpTB81mg3cwcexcyF
OnDB0+JVxCN0qebLN0yFUSfNiPDZU9+V8zDJ+vGnl1w7KKQSYGtRmKRMIbyBo0njpFTnQR7sJ0By
8JSFSsqOT26yQASyWfp8chN2Ph2hDFnOf6gM31cdAp4/YmjCoXgmoKAQJPlZOUKcIKcXoNXAIyCi
N/oay/dypCWAKn3MjyisJiqxG2OY81+rwkaU8ll/x+Gt7iZOyisGoQb8+qv71Kt3/HOKi8y2PNq7
/H8JO+VsU7l+VNZhrEldmM139CV5ZayYvwR6bbPfCPelig3UatYOWs/LOxkY05mzL9xmTHHQWWKN
W1wAtyunyW+KTwKInOfZi8UYDskKT0GWlFAxxTwPH/E7r9qb2h0QOVbIpbyMDd3JREY8hFVOi9c6
8viFo2EkMp7YHMu9+BPEQD979jnTz6H1HIjnj8HrlYJkSEZBDVVh1LlrVzLZ9x/3oEH7Vdb1Zo/j
E/rR/l1JkYgsLMGAfMJtI43YpNWqiFdJRJYxxsgxup26KeJkK2FNiEi5xoC9XZqlbkM3+U2szVFE
lVXDDr3JxvOhi8KK7btZspYAZIQXCocHylZOqskxqVLsxjwDX4R6+epjnyQIwp8TQetTX2Epb/Vj
DNv046/KkPc5IyS0gWMv1XNDXWZYvA27Ee74B/3JPnZlsAZ7FXyzJbwO4zTpYh8PWidetxtwwcVK
at6mI9jUigU4aGP+tCoGOQ77jKuGBEcOx85SRH5r5c5/Dq6CF+7gMl1jBbpCdwUJ2Vd+jnSxdjea
IMm+3DNTBQwsxMyvSTk4xcGchnVHnBzggglId41CI0EJrVjTU8knYfacuJsRPY6+A16T38fsxgyo
3SIQ995Hn9xA0xd/2lleYGxm2TsEmVMNfcIQ/AISj1ytituJFMBcoaJ63Ec6x4G4IuHvUokGBr1s
HkGxNniAMBHHQcjxsmzJ1eeS9yQ4e+AYIh/ZYt32FXNs9fTI6DfEf2RuyMKi6TpRnTWkn+HDJ/b5
nAzB9Zo1QqP+J1kryAHiP40iBMUqL/M9WtUS0W4HvvQXgdoHeLjlkZGT1s7nFvVkEFREe5f0k3O1
1GmG1wPsnjxR3eD3NyXdbKjRGg9M8/e0V9+jly579KfOJkgXnRGatVrHadg8CHjHDZjpmCg8+iJx
9VWZCRpESnr4SeNXF+OlN2SM7pdDJiJXA4sVPYSrRuKxmUXi6IDV/bugnMyMINFoyRxndbCSq8tN
tChI6hnIt3oHF8n3k7k/QyJku9gl27lCC+daGR+RCjQedDwB8pYrMbJV+QoEDXrZfqwX6YarZcWB
WuO1JObm+GMGLJhRUY/iWqLP/NBke0fhxzhdc4jCHoU8RI6w2Tp/jNq24eAVOlrvZXunuyGXIgWA
UeP/OlF0rmx82fw7BUZQ3+rK9niK78KWrXjquzvH8I9BO1ZbqSevvGvvMoGLVQMJY1I3Xgg/3v01
PT73XsRfWtq46VZ2RngH8ipij5b6VIo+/aahO8BCegFU3Nq5CrSyB42iDYaivANKbM0Uj1AV4d70
xx1qXklDFVo491GV4370JZgKqNFw1KbQ0EQAaN43Rsp1u31THKtSTljUHTk0CvbHS4Rw/3lgQF0v
pM7xIcMZPW9Kpv+oQTrNShjdXW5QDn3yLGtBb/pPUyr2XyKdP8ydI8C9HNbhLWDpBcuJgPKfiqO+
nMV8rtU6iaoiHF2P3aNxcLjwDZ//gCUyAYCYgXl4zdRMcVjXlgNnVfvdBHUGG5mc01N/opJECF5+
+ESs1y5t2p1lLjmEK1fmCk6ovJZVU3YaSE0+yXiYNyZHLlH+8Owi3B02ICHyoU2ju+6m2V1BOOsD
RVguTVGhKYzVjmuHnK4mtEXicEA2Rsy+Ef4KiGHUtji1+OG352jCl0W8Wc5FyZizUknDYgYvJu8X
PJ1VJp0920UKgOzlGaLM8bpBK9qkngbp8sFUVJtqi1hv5gXukjdnEnCa5q1mLCu3GKCOKBpK+Z/v
ixzUu1PWe2PsMjgC24sE+O9EcfYlb3Tpsq6qT82MkXmGhY85VC/dM0aFncC+N2MniqVnuh6Pfz0W
phofz0MApZJQl7+xpIIr9117I6DlDrP23eBEuwWt1hnWHoRsSuLDml/04k1GB6sd+4exw291w7KV
aVEBrNGYaK+vTQQ1u4o9198fWM6R+RPEfBuImZo/n5ILPCD1z2wPv3sX+meRrajOp/GIGej4JRyN
4QV4RbKRzBJPtJoGhaSw9wB3hdgDpgcOVmDZHGQqQIMc4mtOTcZxAVwqtzQEqXqEEkcKtEQ4UKMJ
zjULZX0EqCpB5hPKl0GYKsuwbe13wVGzy56QFDdFD92ccyQTFl7P6LBVocD6T2WTU/W2fPKLNiKP
/kdmWRnkx5iZkjG2MQKMMDylayoOWp+dFLn/oEkUSJKHiRFSR18jWEVsO71bmf/rslOAJBKq7Mwr
J2OKd0YVUefu9dZIUVl6IrcVxsSWqest3iHcYQuV1Eg+ukuRj6qd3b0eEIY/lAy/rGDUMG9aRnPZ
gNUisulDXa3IioA0EDK1gzXPzKFtuHx5stqBv7hgt+QCg9uYBkSWMeMi23O7hzCpV0H1wmdB8fVk
dv2O6vgUkDtt5CzgIRQuU0PW/7P8dJqXDmAuxVoKsf8AkzlQOsgkOorXC/RbqvpprQxE8d9Qrgvp
925TZ03r25WJf0XDGCR61vS/Exbx2O7mSEsfddGe3e8s4DWJ4k3rozWGrWjnJcZXLUnb14EktNuJ
3jLyomyV+KkDZg5xehbhALg6BYnFYkc1Cha2k5gN5OSBdZx4vvH9WRIkT61TBRRYrnOWw5d+xeUS
ZD7f5UQy4v2bjyC3fVKWV6wFXdsjAAFcbKM8O3Wfk/J9Gs/6Y0zAybGAhZEYjdqTFfzPx9TS3xwk
RdzQesu0f7QGNQhLyetGNi1qppTomu3fCkMxAE0rwyAJ1hB5pjzUxJxxTXmq2qsRkX3Rd/7Lz8lW
uKvc7aAmFKVMjEBpUo+ydRMI28dOiujpnZWIufVa+oLk9wC2/sWSVfA3SYpz1hO7BobzH8WHuTYH
hkeYgFEbaiG7GNlU+EUE2oL5oH062YpePeSg/ieCXw61CPkTr4HGxerFkyfRMYbvwDN3lUg0A7mV
9sEG/2wdzvxtDDhn+kyPNISFqDCwctosVNqVsyf+CQmYo55WLjZNkhNutO4ka43TtGX9WhpxswB+
loFldXX/hU2P/1RRIVb54VD1Y8Z8oy2VOR1bQN4tMHUMMwcpyljibF5huWvpXWscs2K5T2OPKGn7
VU95PFcBxoyFGFbhsJRkULsH+gkaOFCvrENhLrcycTzu8kYL3JHq5gj4K+CcM8T7Otc/XadNTrKs
p8YzvNKrFjMg/UAYT4/XOeFsINhu84rhNBwSh7v8F+RsxlLK4qSnmmkEfZT12K3J/9eizfD0PJH7
sPWRbeuZvDFZal/2yQkOuqwwPu8/mE+Y9xHl+uN4vqagRGtwMt9Z1rW32/Q4VHVJM7kAcG4b2dk5
XxQyJP0ow0A69ngfXlyTQmGtKKesF6DYEcI682nEZMKCD/qa6bscR5QAPNhUpGhHB3+cqBymc3t8
540gWGpqz+CilylduGeKZhruinhe/Aie9QtPipuxvYIpNCT4pd+H7KQyXV0zCq0UV4z+UBlMqAdV
cpdjw/F7KhoYMaeXxaas8LZ9O83tYSXsulg3cMt2bzOOwkfe6B+PGIbr6bQQYZ6n7lEKjxhT+wwa
YfirPKXQIStzU/DG8CpZiCPcy/1JfZWIyG4vuwESDwtSHvwPw5gFr7RGGgHa7d6ApcnEjAzpCTTO
Wa7TKPuAz0J3XjSb+MbtjPncuNtZCEZ2/yJ9VeqiQHlrEDgpROfR8O/SYQ79PQLxhdX7ss8x91p+
cD+5sX25UmqaWoYigH2voHLmmWE5iNfLmZjHXjs3aFBwVk0GB7eR6F4APghFNPo4VgI0pV8qzPvn
w2Ylu4dCmmAltqm9P6UtIkrS2RaJF0vwZlyxEnJ7XqUAjYVT2wc23zKuiw/WoN2Ch3mXBvgebGaC
1NZHsVWhtQtn83uJ6hozoKzw2HytbFjbDycvjlXyxgCdthzItKbsX3oXzXPKq7cFXUovVYnm+/Ua
hpt6xFo4zMuwuyRndrC4cmaC+ymhhbE9Zt7VSgEwqdT//8SIVXsjf1ajp1X0ZEP0VXMnrlcMdDvI
c/MTP1c0z3yahiDmPVYkgwrhygh4Br1lx18iNk/9S8NPgylZurFVywPPUawJkr0240gTSHNdyzRq
o4DesYWLiKDqa7M3gCRW7v7qmHraWK7dxHxi+wObWVSHPi+5YVTWV8Ucf+Z5U9iu1JJB8fDh8n2F
Nj/MvwhN/sTg3WRKzcFm53aijqsxrkICp5E6E0V+YzdclDbQ69nIVLy6d2/TwqQiT+ktRdPj06RC
eFVaRQLJuDTx1VRHGMqa6cLI5bxzlTG05qXnaJUb03rc8OEzjRv6IFPtG+p9wnv2BoDD1qkRCvCD
rihp8gV7KmwdC6HSBKNbR1f5SPVoHkBd/jkQ2yGipqd+2gQqQw0gUgivUT6E/1QA1zVVUYKXxJ/D
AUiqRoIu886riA40CSpbEo7DL8oWUxkOGZZGOEY+0DTVgKMIgnuRIcu3dRrKA+i/jQTNxT9eFUvD
ywWESG8hIfolqPlmfI7HIgRmbkDhtJfbq2L8pohcHQLvfYWu0ydMrs9cWBOEbLCjc582Q+N3O0hz
SAW6X1lRnDlXStRGBZ+XISf7dTS26zhBQkibhYyKsdPiVtc38mfVVSoOEsSdnXGmfMOaeSSwPY80
Fkl9x1JRrX43iZLYpTz6YpJubjYxS6YXyoE8JN8XwxZa7pJNJ55yM7fop3+a/gnmPnZsY4I6LwFU
0OYwV61HaK/CiyMyjN4EKLIqOdiZwNxpCqlGqMItlWin6yH25VGxsbxsx8YdcGsbJCP6fitYk8Hu
UCdtd0ugpWqOuYxm6b3Kg/1Pg7uFK0mYQZv8XF3QDTT+Bv+6WI039gA7m49x46AFaTMIyYLKN6U1
f3CnLjfsTRCatJTKe92gYHlkhgahRoOVoi9djxmiYjJBvNoxMG8LyC0Gqfr8t0gq1Fa2X7gpQDrc
Aw10gjZGbByU9P+Jc5pi+COL7+bCB9JRV6Y681Hu17J94wDZyX5p0fVFigxFuHKiLYAbZT9ZYoGC
qqe/YLlRvVgnYdT9j08VKNwuwnr+NFydfY2h6JbcNqXey/EZB6YSsfQ3nJ83ETcnB+fYECsmYnV4
fgd8F1GlQtgkxynHPQmDsnFGnJZ0i8MC9QQDowYnCvlemhfPSKrxTXYXUWkXbxIvS7UNflJBaYbU
y5FQNV1yRnZkLEQN36ilMeqCXMqp61LVxQc6dy9xm11KTHJcPZBy/Xz6NxWBHgfwykZrltYGya6v
+z6AwLrEcu6REj09ByJddtIGks4xGKOSbKMk8qpQw1EYYoIN7J9hFNvPhCXfAcBJynwB3wZdDL1A
JBumJCyDFqWmGK3ZSQC0BIeY7pccnNDRnii8NCHTVP6iE7Y+Km5NQ/mS5QtXyrg7mWXZCoSChqE2
g9aEXJYCIPzQp45s8k9GMc+1HnYEU1I1E5qQM/4xySt/UQoVot98wRw+sZfSclkb63sQWH/nNz03
thhURdyobcCjFsjy7GM0JHLFJnD468U5fzvHvOlocqJuwC59GNOI1KwuoyJx51w45dl8ZOaIdx9/
l044OQ+UEAyrk7ftgeRoWhQimZPIuLMdlkMEVpDS58jlG7P4jabVb9ix0K/t61pYaevb87w5O4wt
Xh/tJUANwMEvmE5GB+9JVo2htiaiEuGGCrL4v1QjCcXUFBeKctVXCBDCqGpCowIFpOrKxMV7YoGE
pa8im2TbAS1lX2933pLc59gIfWLsrgtHB9Y9RMCvZJhzvaKaGrh4qj7m2Rz697byByVg2oVamM5F
4efqPl40+qIFstM2tcRayhIlq3Nr8fvkv0mIOyys10S/IMxmI8QBh1SY3AQ5s1ynjKHApLo8WVJ8
v+s6Ig6c0r8g0dq5NXGXl+FPHmMqp77pv4/QQiNk+4T7mq41l6PMvr+Uam9qXkM8nofF7qNSYV8H
tNs/FaVBCYeaedZj9Ip/O9y2PekoxOUbK5AlrXcEBwl23YXh1K2JQAgcBEojOcie/zniX7ChdWPK
6Spt/EISFfeBFNEhcXyChwl2FqQhkGfzRqSC94XwepfEv1JwfrE2Mv+c7t4sAzm9aCkD0xoA26y8
dFt1U6zxSsaTtZtYnN5dMRswg4rw9q8KnSQZjXXV/qUwEjjgS8UbvTJQP544deLwdtH9R/pD6xLF
4OSXo8vRAefLlqne9lmlPI0rJtli8LGXHMlDVvtaetmy5S/CubjnULT9chAPb8OSfOdqPtfIQJsq
YFu9+lL9bBhVex5JsSRH/iFjW+dH16NHwvlyF5nVmQKcq8b2eREDOYXFTP9hejDBBsNHypkDI7+6
03SWFGH0DgKkN3eJ3p/t/r5X6Nf+X4PXi3kJGZvlHjJz0GlsrzCwNVsfpUvsqGtVAX87I8rphBtt
lOmMKwULJJ0aHlRvaoSIpfIYK/VMrThPu87qJDWdU355cgXoy4w93KTgdKkN5M9x4l3UzVrGG25n
V8L1I5f6stcWXgy0t67DrjtIR+fsOGj+YUj0JUksPyYV5SPwy3pLCYWWMU1Uu00BeuuERgY4k1Tf
Q5SDyt/A7nYk7ZI6qy3w2alDN2srt3ZRFppM9NWzYt6Ul1BSfVOac0se5TGwMR8v8URjILxDmf9g
ciKp7cOeYPahRR3EoQ/GLo9YHVwm8K0K+D8fsqnwRlukb7O4hGbLADNAD9Gq/BOCinHE4IeWMSSQ
7vX8/ktdgstJLuzkKsD2xZUkKpe1ZVe5BMUa/m3xZZhfAanCcJgNTD/S6LjRYoV35s4KNjMuVdud
pRJEwbe1eDMf/pq8orUHujsiYh9a76QkafzlCoZpjgn25jeeHZLabvKp+pltkzLKptqSR/flBXyX
ByPs2kUiYDeti6J/CS92Esy51kj0VzKf48+9F+ygp0wSmDsJCj/VNqUP+IPh0LLupixkSLpBKnCs
erE82+rfg3E3aPcoe6tn156b/uqZcmpSC6vpZiZYpp61KG4urWYGIgqXVCSpEdR6bfV4Tc6G6Lay
YumvmLrZOLpNfNJXiSWw2VI6j1tv+/HvPOLJAxsBVeKlwwv94FkU8kYNJ8oPWhu+ocys+LtIAUww
5PikxjxY0jzepvqpxf5Yvg0h5iHlrqUuvrh5PiSiisfHQYbKz9ZLLM/nKwa4JnGPr/lbOH+OWkFx
4Sa7SQoQpqeUMk6CO9WU3SYqxfCgObLf8bzbCZ/5fanIWGjPobdljqZBG42BmL/AQR7Y0ph9LxCU
7RgzR53mxhrpaeMRxrEkdFtXFnzPAyPwwnhfMogBVxxf0BQjDc6WQBNZvlIzQJLBkKTQk+UsWJ7y
0eNL5hjWmioqkqvjEbM/bFi63QBXL+WH3b+yJegT7hpr4qpVksLjKqVNkc3Qh5cgKUDtvNPRlQAG
RPGjLKBL2sYeXy2B2NxzoX0z7PODaaOv3BYLSdokXY15MFkN38P+S9I5+rEnq038MWHR4UnsPrer
X52qDqKHnRB6SbB1N0rFrOO5Uw3LI0aWIc4lInenmaAK5L9/Nu+ZB3h0qWHNATvx7VvJV2yVDd5n
ZbhKeSThk3KTGT1uJDJoGIXFtx7Wy+oPD1u+dfGeiIb7uEaeZd8uneAyOJxCVyUrQ9fOya7MEd5l
W198BxHBss5fAFPJ9MTSNLQU4R0mzhcHzJjSDT7TNB54t1xu4S2RtEX6IZ09m+QmM/sQSdujKexk
zQfW0PqUn2m+OVme27mjTNJT7O17CrzpDxjdSNL1T3Is6mRte7bcEUlFjhF14qqsIhCcHqgmEb5h
6hkKEDVUnclWL49hbVLi5IwwuwShl8O7tvvgADx5djLy2m+mb80kh1Yd6rVISuFpWlN5uQNMtf1v
iQXCmorYlnqIdPoE25IhoiGpOh+CpUeT+/piZQlwBMZhXDYokuSNVWmWIN1xZ2TPM4MawpGNKKv7
mpixE2oQ8nMW0LLGiAZ2s/3J/anya+76YbKHwEZahUfmK2NC6Hp3USpsVWsEHDPuDnbznoyq2foF
AnX6iQBgBla1AcT81NBbBbYjYRpi0aVNVdtL3WpdW7aemSMr5HTN0x3SzCATs8k0HyZPlqpiONQG
vbGzmjVkBrzIJCicXjyH6T9JwL9nYkRPCAJw72Zdld6YFd1Y3OsXcsEYwZKvzb2z4b+OH4IpR0Pn
WYPj/MWLetRbehHvYs+4/twqKzD1LUTuhhUxoIyrq5kq6P9O+Pc8M7ZI2zGOww9ko8+lHO5Ko+Sf
/gkjucgxzivJORmkbOtlud+PS8PUwgw1trqFIehlrWMcQocxLigoIpKnUt9IcMiTgF9b9UY7prE5
ZcsiF52IVXyFpNQmJsWKNFhPnVW490jwNOPuz7VC5JpPbj184X02PgZ264buy50YEGvNTtCkGVy+
hOyuNxd4HoBZBltgDrF5RuzvS0nCuhLtYmbXDXs7zVVWtt8WaoweRQWcDCJltMDL4y9w14dtgUQU
MxWD3WPsSsawXlje1zc2nVFyGHT2pJFOATTY5fSpErm+P/zbj47S52saeb1iovfUls0POmXr5zED
A2RwfbNEchx3be9JMzKVpdn1jBRUgM0UXYa9ZPFLbW4HhyOErttlXjBeuqE1YIhbzV8vWk4DLH1y
LSuv2T99wTL59TJPRDPMFnKP14R9+QfOz8bWJ9Q1Mz9Qq/b+Za9HR/B5ePosbb9CkigfLhXT/3Pz
0wOEFPKcMsMgu+4UHDiUC6yvbBd/dgiG9BS2Zv6ycj6q2hWVC/zzLwckGSVNCdAtJTCsUyYYH6WG
Rxmm51bqPDUwNH/FPgiwPIZa18rrCMsEy9dz8DKnUaOdztZxToF4ryD9wclfVe5DYrKTY8ScbDUR
jXE3j8bxG08pspqxJyVy9luqBvPPGDGw4+t41VMtkGNUmoSaoukPAxQsU6djfAza7IUD+8b1qPYe
4qWlYyb44UWKHwiGjFYkBdJ6HGaBzhk2iDyJmBcNByeanBqZHCfhBRyIzR9w0opS1YWfEkLmyCbW
jyPz6bTYKd1qNLnHgeElNwrr+cJyKfDegS3EqoTtES+vMh/R/0xQYfD03DC5SQCsBVSoYp8R9Fzo
XdYHHwEeJNOCeU7F1L8d2WOjOWgS7irjG8NS/k3Tnvuzkc0N0WvQ3p9Fj2OTzUhSWj46WGEDKEgZ
/5Nq8PcZweIqdVfMQtjNGOn8hzFgq+381Q1a4aWnJTlS4A3eXAfyM30GwkASG4Y91SDPogRGlqGh
hvRHpm2h88139riQLgCQbDz6aBuh365TOH0fEvqjHOSGk2TeGr6ELw5sir0HpydCXFuZEnbHBWCM
6QE2S85lYUjRR/A5QFRfBK2MuqbnsunnN/8I8VTyvJMLjFGlGrivVpmsO5bGZByUKBahyaRwmiig
HBdBy2Rz0NemRkPrVc4aWx6desZ90n+In2RxzBEoepBAypIna9ZJ6Z/8rWLEe+N0bxC/urwyEDc6
/0a0nMOV3uu7GgtaiAOStWAlymN7qIBUlXOUx/0BuYqOr4Dj+AQPf+/FvqYodmaBkvatZ7oPAV9b
JPJ5lnAT0Tnt4xbQX+aVkK+VxVPHdL0hDoBSgO5U+QbVQPnPDVe1cMHIM7sjNBCjM17+sEhYg/GW
1V58wdhNvT+TL7Ekno5YfwmKq1MyEfKED2k1gPCePiPy+UaYg0B1s+Jax734yufO4N6tGg52mhav
5qIrr72T7wgy/0tYIdjA9BRRRRxXdhUk5c9ajmWaBeZOZYS+38ahKXBQiCdFzznJzm7OqTmZQjf2
1OMt8B3fxwTm2MAG7meC8jDW+x+woBGt7rcMNOFMq55Qs00d89zhH8+z5eW4GDZdSyvsMcU652aq
4Y+OZuNl2tne0kFhHIU0f4orZVqz46CsXuTuooPYAYMDVc1uOwe5VZpzdz8NXdU9XF7VP5xAaAKY
62dDqr5gjSWfF03iQUz/VNasfbjEXy5YMyD1UDXb8gJftGEYd7lCdmPsIOiX2x7pJjUsYfNxQjL0
c5VxRye9qPlW0Ly4DlQ4/yZi6fd6B4q6c7jTd0iCvwKoqsq7iWGVWcfXT5M7JfLVPr/4RZY8IFUu
ssgmpT/NKWF7Ye1IN1dZ1zCe3sAT5jVE44KPEbU13XEh0nYeBopMVPXki0S5nZdGiy5HTc1ttOvq
rHj5CwS37WhkXohe76gJgRUa+FTf0A/ssQo1G7M5/Fe0Tc0jDrPM8QD8QZBjPR2uflMywqm8Dopf
jSxgjRsSXunCc7yh6XhgV7Smk1BWgYPUfjwQYKRsh5gdRSFkpvT7aaGYGfP25ZpBeh58KboUdv5B
/r4d1WfCNehuBiG++pLlYCtGoWMu89XD93tu7gSElrrD46oAnW0Kzg+jaG/Y6kZTBMgVBBkuRDm9
TR6d1P7EWVUsPHPhDXG97H3elwuBJlwlGZggXpKxcigBC21PlTJLYXppMAfJDp5oO4G6Mx7kI33J
/ohsEjU0hjroM3N1te81Xooa7iZ8k9I9uvZRbjav/3R7+PYxcnpygSoGUA24CNBGYavNLht2MHIB
K7LxcDB/wExkCmu/WUEEI3zIWinOqzEi8NM6kxYv+fxBuqPR9RSaRFlYyeh3ycI99TL1h3jdKQU5
pfBh7qBn2Z2/u6yzbmpd8lin8XW2BLMMZ2tDteGPsVY5F2t3RPrRehJZrV9AZskv6SS/wvQTdTJx
beqhJvsbxwcPBjilvHCwLtE4fk42rwT8bltx3on+EIhgOM9pFNnb+4Fgz73tyUqGFLOf9JbPGWls
s51xciD5uQDfFSI2mBwjihwVTGwgYxjLOzCDhmHPJhp3ouD9GL1sNaSxnUtEUUQkGDiOx3qgmHXk
nlgjSuc9PpMaqpJ0BMRMdTTzu93V71BYZeEH8n00HeMAm8xUk32oXIa7WtvXIs6G+K61gagb036q
c/Da1Qkxb2K7CWsn1dupUo6uCp5e5CYFgeuyXB3res1de9l7HMIYHJqN3SBH57BuaeB0KWv54iOV
M3Izur9lZMgpjWQtkmedQgzT0zqyamOmN/GaeIecX2mgIe2pP0clhv98aj67ZzVoGsYbsIost7w+
UztbydVth0b7kkASUZ69FsdjmT9kkGcSzHv4MVGvbJHvhHcu0p8lDHBm+DvsqGU2x7+c02t3+hxh
rvO5zs9gu97UEnchJiNPvkEQBS59ZM9Wmv35bC+T4Ddb8PFKLdUwV+Lre9/gDaMog8V8Z6LUqHvo
Ihmxfflx5HEUWz7woOzUUWGm28qcLZRBwzqbQHT/j5uMHewqJlm09lkrQujVu0wD9tPV4FgciN+S
OW767bl6YSoHpR1WR7YWjst/QNd8iAYV2X0r6FTQxez3Kbi3thLEuFLHcFONohnjwK46jXn7xG4G
YtptZLwcNiPYCGuJqo7SZpnLEDWXhpuVS0CXAzrbBirGoVP3+xqaT1dW1nAOWMPpL913Ch7WD7HH
TcqmL4HmwFiC2kbyoP7Zs4B9aPATH/iwVI3nicLLzgJ7kuWSj3qVSg0jZJJdUw5uzbEQ0mKV9fcI
4f3k2ntfxRSmXYobRR18L7ncbfnp1bSkQHQCsRv6o49MzZLDbph+y7scbBga05Ddp89UUZ2KTpkd
Y0ZhS7Xu3PWvGyeywvoYPBS4Dk+XH3SxF4MzcRMcrFUdPPTuEB4zEGa00LdCiUmP6ap3pIcyGcy+
2FUnD566A7LcbjNL1eudZ/f9VP7GddzIg+XYqcXo2OoWa0v01r7vlsw1GAguLQ8PLRFDW5Z1KcGV
nHuGg4yveYKUU3BC1CJN0R8yOJT5Psbt0OoZktn7jkWOZ3LXig3G8oEq8zCjcDW09Eey6Nn+P0f8
pr2j5jHPUdgT8ObBVz5H6h0l7eQ0CGYopRpxfApxIEkZgVba+uKpfGZkhfprMNN175qcPEw/TtiU
f7YrMag6gtJ0wrUZi5/hptWQG4h0uuIer+roHieLc0i8Pxtrvv7+Zfx1bdL3gkOy2BQmalIKW7Ha
ZBQKSPROI/FIkrZ4ots855rQ7+wdu88r4gPK67AHh9fIdBGetZedk4fGbUyWL6l69jVy+7d/MqZl
8Fc9qLrhcBJ2C9iE3YnV1wemQ0hzaITJ5T2uUnoi5FXiIsNI3ARF+LluyCXcFdrUn9xCd2wt6QT7
HQI519S4vKhW+f5E7fDUqZbNoem8ealaa4VxZA3NWiwBYdO9rM+DMi2VbZIEYPkrgopSvEhDF8Az
JrBj63Y1do6wSL1wkrWXhQeAq66Ry1yo02CsLFRNiP3/S4D7bJ9mrwp9++6buT/7GSFLrFSmXFc6
jq4EFaSwJBj9pneybSzrsVV7DYTj1xlv26rys1C/tIhgn+jBdAS00t0/DSk/IC3txcGkf9fDB3YD
Vd2LDfdZyMpWv1GPXmtedMxWoUUJnErEX9e97U04FzuDmL06D/tdoXircSDc1yg4SPp3BWYeId/d
iPEXO9V9NymdiXUNG7aoocJms3m0afNERT4wgHBSmvLwkpBZDhopcCREewaLK9hvWUeCj6ajzcZu
c2cnrrny4oAHAnKnJJXJcVYhYI7JK1J+Cz2/CfoK5e6R6sTFtJ7rIH32Bg6ULyWsAFxtkOU93kkF
RkqWON8rt25NdFwEWkm94f+F4u7ThPnLCa/Y/SoFLvar9in2P09MrD3vaCrGPalhg7a3/H5fjnVO
4WnHiUJigV0HJqb7CT4DbfDADUbfrYGYOyjWAx2lj9lyVyNqw6Ka7EeXqePAX/cj1BCxUL0FIT7x
uT+hp5nFtI7BdZAKO+SFIg+sTAhqLuDGfyyoCKIZWiGIJtr4Q0l7WLsEyeVw/dbirulCR++Lo1NQ
hNFV2Ptb4N2azjep3bBKAhEkYvdl0T+7hMesy4fSDYe/gNRe17NEUiSuivo05VGz39KNooMJ5Rsk
DvglIH9HWc+Y54ii6Evsfx/G9fQDBBscM2dIplwdVmp5guLmjeMvqB62CYUlnUWxS6KLUHOp40zb
uktlpKzt5cMYVAsSseN/gnHd+rqJparcVie1IXn9wE0iJeYBbyTr+HB/KWBlHslqdSwEsiSbO4LP
90bNN6DnROa66/TrU/1gO6vRMG3b/h/fq/aCSF5h81SYCjnzx+2TsoytWvxqFoR+VRPLFNjdaQGd
uB1ydvbhBsWfjUwTeRvve9zS4HMhGQ1BAuFY9a1QOgslrw885d6JGHGnOn7DMQIs4SiT3ieh9lrb
GUbDFJGZqUgnWfvdMN2igoCjc0ONII1vg5pdymS93XbjXb3quyVbnq2uf8Yq2OJkf08zMWvxFldm
AHsOu5ZNI+BK5ZQbkqh/Sr8WHf441xmfmTe8Ey2neyLeuRBtYO/yM7TvrOVl5fVMgLflL8uP0dop
CPi42b5qqNeyYr2j2789gYvHIaZTZSZCZ1FeFazq84sD23e6FeEImMntdEM2t+Da57oRFDYHw8da
yHSZ9JZeZxTp8A+lEyJ5K3Er5c6kT6Sic2oBolxdvoYlj3Bz1XsnMB4z7LQTYDe58aArqlkPw934
Cd5DdeqOpXy7VLFBnasJ+T5JmEujI58OyGKjOVOcm+l2tvsjpm2WXfQjNTAaHzHUWizYcXpnW881
dyBIs3Mq/99g+P45xQqL3nAdMT3sDujOQbyTEys8PZG1OyoZ8XjMogAmzuQFk4LhnEI16dlfKp7R
LAVQF5FG8QLDlgRrILHLLGrut5PADKAzmYKgwbj588eklsL1xU9DB7InFMHqgwSf5qo6LumX4Dlx
MlILUqXPqKAZPEzC9PrJNHSz3287WyzNQBqKtUi+u99Li0l8H3/o6PIbh/JH2llFf9Syka44IPPC
MQHsdpMyqXjp70e2KmB4bFECXGcvj/7AqfNGzmC07cs2+AtOVfQ3/VyCl5b9VYPiazQfokiPxI3r
QVeGbQVpE8uCBYrWkV1xP3jsNxqtBV2cOW7SnBIzXnsvsiuI8lYir8KOCzXy1OeLacb9Kqi1ncwC
bm+uXASN+mqvCV3b6mNhlkuBP+ImQGOBLSF/8pzIYWXOTj5ZkFjMdpE+BVyFjeCA7PYAHVDs7pW+
pmCjgICVyklP54pzcfLw3TqQD4DGdtqUa+slh4JRCuYdOvwSQdnVhsMxUZvhIuByr/630kq5zFsC
ndyqsO5H1wRuJ4AplYDf1GHNRup9vmkzrNGIBTSfuHtpmBjBQrAcBxnBbWIuKT+qc7UIiKqS5dDT
/q1M3In0zlPTeinMlKsusKTSNbLEbRiWEt7LcoiEl/04Kai/qcDXjJ1CHkSr/3I2NTCSQvJmxciK
6nWpyQ9BpEiUsCk/T3kvz4XKHDmAceh36+UqHNu8F/vV+tG5EgeLgRgTJvLPt8UzeslZcG1uBJem
1gIZ/fB+3R7qNFwnDTSrMA37xat2u+pAfTvdjoDOqwfw9Yo6gAq4TJfNgnhOyJ4YUWk3laSmzLSn
IAGGquNZgTMcwSSdm4nLJNJl3ncvUFOf3fOrndFGch6CP6oPlzh+ScCh4NKcO4dNLsOFMBCcLT7R
63zCmt9vmIP7w68JGSKt6blbTk5IjCWiPeGs2WINGEvwRi3GnA+xyL+EKzXDzZJESubgnnNiLK4f
f1pf5M8aECO82HZUO8q8Qv5Q2/8bG7279DdvSVi2PTuMX9w1Pt4ff/VRfMtK3Si9ALTBv1+9kwiA
5nF9sMmXV4Qthv44ZsBi+nc+BWWe699L+vnhU7e1zMUbNrGG5YI+sdv8G5DaSazdP0jtScb28uz5
au9kIO4bvQZt/7N3D6999LTjL7GXTDeki508pbYPAwTpnVrWXX6CUtgli7755ZlQbttLcEFWh+Wu
JVbLlRvyJZ2RGW8DSvAkBqAPdjuR0Wpl9W9WvLe4r8VYWa3G2MD+QYJvqoP6e0KjLma9fomubgiz
4UqHKIfRktYoPJk62PnvuwxAzxLBP8O0ldpwCAm4j8aE0KjR1qNO/oj/g13uGNu5nN90Fk7d+Vqh
+8skjWMzo6X+fCfgZBD9LAXZEJg+m9KvCV7NlaHk6azLQB6RYq2jloepEaP24uEGBJlct6OeLAiN
A4cYsjaELSSyb7pyJ9hhafxl00tVplouRYr/z0mRxGBqX/umGSnMYmdFvmKu4dzWJKmscA8mdXKa
Z7MOoAKhMoD03TsGL0f3H3ASScJGWGz4GVI1/VhKo1mZkrotzEkb/ScPLDsv7+g1qb15SbNYBSuN
LjerFEzOrNi3hTwlkV1h9FqhFkPTnqaUv6f3ysBjzFK8khgkwkXSKiJIHFU1l8LldeVrP2o2h2bl
Rk9IxqFX5jr3zUtSKzQUrCyKP5dVSs8IB3Qu2gzuM8ns+fMmfMseN0Bvzeyg9grxF9/HXfqM9BTM
SbsNUE08wwoUXEfc0QAqvOORwOlbYaNdaEajIaFWIEahQUKeB9hIkh0QQJCeCwc8G8YXxjkhmjx3
mHFOmQlm13M+TwzSGit4NY6lmEyB0ooJ4xhdlH2uTQF8Whjtk024JjqAKllahemK7JGZ8+fjj4KG
geu5tt0zbSSkVgG6ReAxmub59zQdqGhAne/oWHtgYi0REmbwGBlzE5fax79WJ/FycIU6Dsxun6ou
MAljGaUZWC+yLb5ICFEqQDQQeP0yFAhXyReUh5Frxwzf8OyPLh71PCEbynxObJJt7R8SVu1GHTwY
ZKwDjS6xAZkBeMvp3Y1NvVtgWQhzmPA08sja6fAQGwVkkEhkzQ3MZpcb9fpyr5h/NDfAmzNgYQ+l
vPkGiL9pCSA+2hN+ycyr8y8iJMTwVwoXu5iETKYjVwzMxnrhjvit10YjiW1y/HkGPXUvKULzdTUm
ia+s5yHQ2lB6xqZgB8ny+U7euTJwm/TiWKIx0457nKWfGj3HavlGvcxgMvw70aGPGGAzftM4og9k
mhbn7cVc2cK5NlLH0NPe+jmsbS+Pt7hhf+G/06gHUJlJfJDZ3DLju3mNI5IBDvIxmmUZQ3ix6xLf
AUE4VQOz224HYxScjBIvKJWN5f333J3dAX+PpBsFGgEAfwx/H50QhogxiO68kECmKi72m4AgRYG4
kdKDwwIYx3cz2v0LQAfk3yX89uwx/AwLPaSLnQi1Z5cTpjGZi/1HTrhaQt6OwreuG05hUFxbbAF2
hNqBqerVRaxzosz2RPhj7SNAZLG76OVXL0KtlgN/dixdO1MyZYBbP/w/jTS6oioYkbCdAbWOHR0u
vhUcqSKLteMEIuAzbL3meSHTM4rZewNVMtVOHqWCv+KWQNgsrERYbNSVBcfL3/hajFXfGwxsd1Nt
4USwzy2ikM3XQxOugI3c4fCH+4rKqWzFHXKHuMv0y1RwPIej07N/ml75ag16ajSBwJ8RSmdCZ3x6
B0s5r9nGqTRIVGW1EX/CcZ/hDfFusc8XYe2vZNGtINgxKeZ5J0iCxqmzti1YcHvTGr5devdN17jG
a/+yxZfJ/YuLJOofIcHySkTJTQBR8/JjYXRE65v2FfTxVBKPdDZYamoiY51A+FzsfnX2ywCKj3pw
ZJm9377BQyfeeS/q93zRe3K902MuEgPcSiaQ0M2EDZwMDCwU4V3eMsbaOkKzEJzBfU2G6hjBeFdU
g71W043vRmoVs+agM01i1D031cYmUhs/TuUxEJLVF0vuYcBfk/ATdg7bgqHg2bOk4rWQMo7omAFC
SlISlI/HPNraorP58PLpDZWg/Z1ySn8e1fwW4yiYq7w+Q/yW+CHNPPqOVAKp0dFnoSDQz1trJM6v
ktJy7+PoyzS4RsQXAzrEUe3y+wICMsjfIK6HufqIkUJaFdu/QP/hvStonIc8xJ/HER64cpbD1y7A
bhUcYKxaj2D/4N6TsLsX/WV/0qXgYk3CyLAPWSOovAiArr/fokaKsj+fpDMIZlSPEEBWmb6sP0hg
F/iz6nVfk6WQtY6HcuEwor2qHGT4wEla7gwl8bT0rEdSkID0na4lk0Dv2RO9xfQ/LnPlb7WUnyFw
zw34MFwjaQMOGRpGPoTk+f4dxEgh5bcAZjFT2Az8BeEcx1kfOIjJy+wXZ4nzqqqcr9TPf0XxnJX+
zLHUfJD/d4cLwlf0K8t8Sn/pSxoxCBVmHkACUfzbVvUR7kFVaggfGuYmwrH1k8VdTD0Fnw+GPSbA
kmbNw4cmPEpMTNawfI8d/IkdqARYoed/66oNi/yo5appNVD3w3xKbsijK+IRM4q1uJyuumfAQdy0
rttU8VFJGQFXb4Smk4A5KT7hJ8s8XxpW5vY2yIiBh5Wf6ZTulNhXXmRSKyv46N97wrFspEtpLU7C
sZzLVdb1LzUeRX7zL3YuDNlTrhzplJJlq5CzCoYxwKSQ/GX6vj6b0zcrjq/mqUFt9FnlPdT+ymjZ
+7hA9MxP+F5HqqWcP9hLAhnAhUNnhnm+EkkbBnl7zokjyf3DVkVy/GmZxWrrsYNYsLaFRCX75bAR
V2+hGo49c7pvKDwZYwW1CU1DENRzxbbuqsXoiZNGLYdg8WTUC5a0yDWWRweF1Fts6Wqr4Zu+1uN1
bh6FENa4cK5p+imVK8Qi+mERc/eAOygvrO0jy/CRDJRRN0RattsyFvNOdb+QVl6Ztr7O+wJnlZ8q
R2Jbn6wl6MM6q1kb+RdobIWAoWip8845wAOeiXxpcIpqQIU=
`protect end_protected

