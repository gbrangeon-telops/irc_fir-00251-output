

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bvOwtDo+u1XQuHmmirIW0G1Eep8h4q1lu6sagQVNOpqoo1dUL25zlZCKWpryXBrbavlsSVZj+/Kj
u5U6Rqq3pA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R8VeuF45EN20zhkGmJksRGl35KTSV0YbXBmOJfN53AFOKNxf64co0R3kMl1KH48vuem/BXWPzNwW
17k9On+EP4ryAUZ6V1YvtlO9Er2xv4nZefuEO+pELxS67R6s3b0HhdPIKa2fxDF3e7AwjfjDxMiG
HOQbqK01rVOmqe+2yps=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qqYTedtVydnDu0uy4wgVS9xnI5W4e3CBu2tom9I4ji9x6Du0u8YzLw4sHBXlBjTr0CIBWi+453uv
6i+HBaHUw6WLmgP+uD0PvRoMp9iMm4rcTjCZCtUo+5bxaKDQQyKy3VozWJN9cYsOEXUyn41sbHk0
MfnFQ231FTzHKrD8+sW8iXzJhrvAxVZSOCQNc8FKSuvFHDKgrQOZi/Dde7fskgmy7Y+pQzZQUv6h
7xsxzMyVpdCwJjhjdow/xj17Fc+yTtNKSxkHMIxVK6RXkbOidb7jBkIw+8aEzlqsG5f5vpboGqLH
6uQ8IqqBeKv3BDowwIwUDotWgCgTdyFmv35LwA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xgoCG0tChkhv+ljdCxpV0I73D5nOgliZqF/G39R6pkQNEQixpt7jSEz4sP4s78dR6d8BiB9A3KNg
s8gNghB9SqKmhRG0Jvm/hSIBQCWAqWOwg26IvTnT3j3MalMVsj1r5WE9uyiqdJ+QCTo/Y58NBx8l
pM5ABblrTJM59LnIcqI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VTcA7V7opij8+vJ+tjjgJGiOJ+o6V1u444VHa/k01STvZB7T6/Ztq4KXHSVmD+driESiC+2EQRes
dfVcUifCMaPU4kNZrlpS+Cz6GGzKHuujVBDhNOZum+ncGM2VGmayYd6F9EbhwKFTOVOkQmEz/eFL
4IAryyIE59LghhLnEgKJ/yOFNS6XwipLZ1ztAAj7QDruS/h8wJcmBcjwC4vXftAO79YXKmVgRKly
SlrrXAPgfawAm5V0hj7SI23oHUFrT671NQiN+jfhZylivDC/aANQXHsoSuY7NkiKvHESuXKmJ3iX
cfk8aGjoqSspgWZUBuwV9vfaTHDt+AtBbt97TQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 174368)
`protect data_block
qoKBERgM6/CXtj8KoB6CiBcVMxmAjORk99mr5WoofRWEl03UlQer1dVBWq5TywWitkvAhHJ+iluL
y5CeTf8Xi9OPB1EmpM5EkJ7aVSNpnnH8gnJr7v8S8lmXpblaFU6p79RZ1xylO/XdOI5eC7qx4Tzc
gMBNv7hPVCV6QbhvL1eUl6ghmS2wvOiof0QitSm+BSCVhHGcKGp/+KexgHt0hMnhvFPolDmV0GBY
4ullELRmgdyAqsUF18MsZL6AMtVUst364r3wMa5Lb1KAMz2uCne06Cnc0UH0UpkUrCBIJthsAklC
dEzzt86cgfjNNctgRccsuFcG2BrZ/CFJisxtC+wFHH7hQR0HQ5Fdk8FOsUgXn+/53hLlNMSkwnLE
AQFWwv2vT+pUApudj7HuLQf1VSVkZho77XROK0TFHyL8b5ft7VANYbbPT6/QPMbn/Xvmedh63Ee7
8T6vfyRU540sI10mfBcjGFltVz2m+6J9LunCD3HYaxhqiP+/q7qkPWsUW+MVphQ0PL1YFCRQ7XVz
rwYHK2Xs58Iy4skSmlLupdHKII9+DkADEKmBQdXznQs1rMQALUjkxRtfSffjye/p8g72IiwAv2Qc
ArGOB1ldcEy30FIRIgdf92qhPb6ksIhJODthhJzDA+8xL5eLSrIuOhvo26++/Iw1mylgp1h+VOFA
N8R1fFe3YJ5E8qxH6tujOYujfyQwn8XjZuaS09754x/BSu7OstzJ9G7HQsoxPiwgHgcEhGXkGNcE
84Sy7AxAL8hSbFrCfMtCW34ecSNCu46FoMa73tw/68oxtpvMOzuafYPh7x0etuanuYXPosP9mAHj
yEQ2hojlheoyBVx8iV/gPCH/OF/3BS/Taz1nkDzF4FPOJ/o/Myu7Y+rUro1S1bKhQPaOq/ENvNuu
OKVeBG5jbqmpq9D3zXWfR+dmmA2v8HiGqY45U85HKk/5NS4RB5znblHpbZIfV633V61wRSUiw/z8
eF3eYQMqTjGiZ1GxKiaXTmyPMGseibtevcukjyNR+dc/LBW0IG+QuSMNY2hhR5ow44GNViNHJ9tM
TUlk6UMAUU+aXOD6+ff9SkKU0BfE60Flon/2GZG7eo+xgKBkpVihdWJuqGuMMyLSIrbgYKTum6M0
BrslxQWKhT6unVoE+YN9/To4IIm/NB/PMwGUNi8g9EPocTvZ+IdbMsKP4Kk/5e8cgaIP+Un16zx/
ilCn4n5iFHXUATw7sOyklFvUYGuEktr2LhDKWyoh8GjK2eKwMBk/Lt0QsvT0LGx4la+of0y08lzG
9nrDeENCG16WAPFlvjgS7X9zuHjalIdBGHTuSkcBTofrVXe5PQg2CL6YxCkfWsKPMvEEz/4+vKF8
KpWTSjyhdfT3UvY0hOrtbIkyUIRnpCrjSlmDdHJVHKpOrcx5vbzojuhBuQALF7eYxmq1quvH2Kad
xd0HT0zCbemlY8OArEHQ5FeKgTcLOhfd94gbMMtUf6d68pQwRUOUGuebLMjkUy6Kt8wGJSWYt1KW
uJKnrpphXtN8mksxVxO/c7bXvD4ZOvxqTsjAI9pQGoXuZC1+IIYEKviBfSXbLEo76y+Ozeofrd1d
v7J0GHaxiobGbqEwNRsc8oWsyXGXhWAUI57p553UPLTl7hcy+MSeHGU4N3jCwe6VakiJdDDt2AnE
1+dXSbK/s8hKIhkdg2U39XNOM6jGpFmqn18lZuVWw/HuM2l1seKdhUQUvXFMOts4q3vAz3OWIQJp
nANm6C1G/dxeQeqC4O+xRJPf31JuhlOk9eBsfS+ceLzIJhF4LOTGrlDKvbUVlzIc26yWKOwyrB3g
mHMRgY8RgdOxbdowBqzfa63NCEwgvpKbPo27cTicCyUoGTQCWIgJQjhpVaY3dGvPabNlZRYD1Z8o
cBGgNyb5D5qIWFcbe29F6BfFgMrdos1772JV7iVSyYHIGUM+bf3y0Aa1YImYyskJeO+9aeGvDaRx
yCCAgUhy0pqGFXjDEXT1wb/1A3/h7gqpY+8GlXYxqAsDn5jq9m5qfKoV8go68cXCVP0XpB0FcDQ0
nDxqHNnG5fOAuUMNnPUhypilVk/CCcoLd69J5vENsSW3ASvieMfM8iqoSCTA9D0GGmR1K5bahst3
s/IufZn6ZExBppCCRRwxCxgusu8cmv73SKs8YYqBCxBTj3d8aImP5zFuppRx80jgjYbHNS9CmA/v
hfDaSbdp02Ja6AxLpNUYfa7mr70Wq//DJZuCtEZv57p/v3MpNJvRn/hd3XOMMLdUR6jTKHCt+AGF
CKtAnxkGWn3E0Yu/nr6YcwMlAYoECFP4KVQAu4DLZ074ycCHmn/FEOc6/pgC44s6HT+7YL7FnDYo
dq5GFPdrql384Un0QhNnRqQ9LCl+vHioZ7tQyBX8KZIvxUMsBekHfQHMX27OHtYd3bgGNjsdxNbM
1cteQcnuo87KzlrClEZR58kC68j0b9lwXBEoWfpeciJghGJ4+Hb9TQK5i3V6naFpRdvJ+U6jOwOP
GDqnHTY6xKySGLRpLk4Fss8OzIR6oXbGMr4z3QMvFSlQWrq1pQQ5OxHtKbi6+awLqqhu79mK5i/+
EXegiK6IYn5GX/asCz+m7W+/OOHHaaq460gV1EX1P2jGFHT7oomorpGYRt5iAypk1ZAexilnELYV
qTxioSGzJaZCyF6hBJ4ftbB4Cie/OLy9NKe1VPxdJcBsZV8yPSNN8X1jiEm0XhTILBO0/RdQC2R6
0yFNFUQULP3CwMSpFv7i4NgJvdHc25kmxTUt5hzqS17LoZW+7AJuHPG/vyjG6+vQfEiDcxmVR+Qm
CqglS40gv8K1oesmtmD4ajMbwihQVKu7Mv01xr31zqKR8yS+vJgCD4cMs6mhyFZoUrsZee3/lNSv
WSZycs9txK97xNhQNs8D4alKBn83WRSZvIk0si6a7hKjNK3O1nsIS24RuNsgveCoORyg12VhODo4
Y2BSVS2GmGJ1wuQTlgzbstGLpEmW3ifYBj117ei0kjjq+yfzhThnSJ5bBrOiHlHlcvQJgkqSQuki
s8LWXz/u+IWbDzfb+s288hKdD7X7R+3uIzPje96Z84PhBrEIUbxkTkI2jCvfYigLnu/7BUaQMswC
AUCbA8NTFRC/oOlhkcibGmfk5O5YSYL36ulZGcmV2awDVT/Ds5Bf2Gi7j69tLTc+z/FMGW5TmPox
hhWemj0ZPKYlZ/I3dpcGAOMEhbuzQwLE21zX6jlhKZ6huHniAjRBe386hLpQjuftetay9QO598gO
OmdpC68wLJfuQug/haPjkXebThc2AvcMTM7Ju9AMSozyZvCzbWCsJfRSYYwHk60TkPK3QSGNWlgq
HNgILhJxaLJtqbbr/xfswatwI6DhUziI/Gk9NReFNwKftPiX4Yi7FP9dM/l5G65+kjjeabjmrngZ
1Rm3qnjYKboWh/drePeMAU4Y0VhsfzV4JlUM49gUi1GJmK5bO9fzOBfzYrGd8VB12qQIvrs/YFqB
pZJzH+1deTGzZs3ogoVcckQQGloTLY6NLG1iM3rhWb+DfmfWiMT9ezaottLpynH4gU9IshYzMumP
uHhxCo318qYLMYi6nN3wUUZy9EzbVpXKDYEXauDxzXtNT4DuqX3E+AzfHpebrsmmq61j73FWnBtt
ojd4JPiwzD5RbIk2JdHevgmHygot1Lq6y4yhSVgaYrjZcHhUW5oirNzOQRcJdL5+dJ4aS+4l3LV2
19+RbFvn3KGwEic5dOa76FwrYDjAxu0uI+qUyNTop9ShJ0+mQ2djWQ5MDPQSZlKivcRL1wXG9vw4
dy7Qy//lzpYKJNChO70ZSLp14PITEIwSkI5uPx6UnPW2eY25x46Oej5ZOwPi0zXXgBsqBMuleu8U
/T6cB4xB6X765sgF7AyHO91h4E81mWkvm80Cd03d5ZEmRDVLk4Xk4FJ9pdINQ6HK8fpsDGIb/yuZ
FNu+bYiE/QtIY+SyKW3A277HXcj4F32VmM0C7Q5aSPjbykJZQ5KZiMvzWjo0rrwNcR0efphg490k
/EeKlYZ7sOSedDBRzWaZasAV6RKz5iyj16kiZAtOkFNQSsDqR8atcRdlizDBt1My1qcTlM5GsxPy
mjADkPFSHm78pKjEXDxFRgTE7iOdkQ6lm6gYK1zMOHZasYAafvaqHLA7QgUoD69lC+mKgFwFN4iQ
eXte5NGAGoWmseas8ntC0tINYPpGkqUV6UOG6d9H4HpfDBQ3juwxfJy6tpKktSDYkegMAsES1Vvk
PmTcyh601dkS7CW684T2WbJskfH8weMbmrsEFkcxRwyzOwexKECweS4PINYPnxYzVESNqgFxcP2F
Fp23oCKHsLLBMlqdlFYKL7uB7hrhbb6onzuHB59leLB4gIOvhLx5I+uWMGqGJjr3rQEQf9bhyUsz
rwUdWAsMZMyj0Vt0OxZK8THnNGGEHHg/fKc/gR9Xh9N1l4+Tfs/cxi7Jl82bYD4gqwYhLDP8a0Ca
LH9bbHXkBPtwNdzrTe7wPilLb6voKfv1qIwdtQlJ6J+Z+8mFnSXNovQsmIlKfhAnieqo+aIeEWgz
aA6+jRSzZNjLd69fzuJfI+u4ZqL0Ycb2ua2Zw9J1f0hHymONQS22to5DxP0iWsVie/5FrMr2BGkm
JFTfVLEoK2Fvoju58rHT8g2Ot4zUvCEORysiTNfEgT8sWRXJ+ZZ82gckHlejzSsHoLBah7fut/Zm
TdHcfdZMiAfIfVAkW7CLADHubG7vtDa43i2IXYH6gWlbNq0fQeB125M43jpm2j1qUBXwDtPhyqFj
lIkmUwCWJSju85fFNmUlXsXe5EXLRhZJeLSO8Hj6O+KNoxWGDJhMyzxnKsiqdNPr/EdrG3HZvnaO
dRcmTuv7Xxdntru1u96FDwRs83DkyUKq4ag6QmzyURCxswNYh/+YzQAWAn7FHarYgmG5zWO8oQIe
I5910txBygipEPomFXojmVVNdBTvTTDFDxG9oghnRmcWYWaKS3Vbr7IFXZ2nonpOrrly53S6DxXq
r64Vqvf2GeC1p2eGAWmMShz5dOoBfQp7k4knZyWhE+UryJ9eS/dhbekAiVWqHrwbTBbtoc8cFIsQ
c38WUL3m98Wm9OcSmXBDbxmE1D6VBwNhztZKXB+7bNXayponOzz7xFCmhKln2ZpxplgKKZOqceuo
cYQY5OdTderkrH9kzIbdmDbUEW//DZ9cYWgfJQqwB4qQZiAfDxSEqG9d3xuuk7ko32dg/9rv8+xE
MLjh7Tfm3GqzV5ILBn6b2KYZ11ipUZRCIYQhSxH1Tfhl1KsWNt01CrTUiIa9cPWuwm+72s0LeZzX
FQ/Dy/qxmITIt0kNR+sRzypt5RnEoUhcsJVgui12A0KMSONsdCB/dhqT6zsMJbEHytKK8w9VQmzr
0Xf7nnoNWof7xiiNfgaSJWTDDIPGK5Ma8Lq4V0tUokoBPjtoaHQf8MWbsJkg5/nng/etyDTp1mKV
an4OmLtg89NqOGTE01wwu363lckXepPHJdxzf12lgrMR5ux0xA5y7ZZSmBXohVD+scejiSea1xiM
4+Y2NK5+DOqY5W59+vE48dxm3kgdjuGlRTYBPjWBf3Lt5Zc/Sz4W9I8NhZH//fUbDVJd51QKlK9E
TE0bZ7lCBgkZjEZjsblLIiU0CmozsI01hGiNhzbmLuYUfTPMbdhFnBfVNT5LR4rMVymcg3sKB9+Y
UhNnnRIG5pwUM7070d5nXN2kJ6O0jPog58UATpfjRm/I0ayQSZuUseq3uxhRpZlC8njIegjE2H5c
HNQqdT3TsDHtprLvCpDE07b9k1f8YXXFGfIXRrbStScn8tT/qpZfnD2lDmtf26WZ7HJAUsqaRRrb
37LcSUe/DELkvDjpalkChDO3Xi3cS09a2ie7e1czqt6kqkknFceKz5ZQVNtGqOifGgLy6yZOoTqh
uq9oSIuLxllz/RD8RgQSoBDms6DshAls4HZi5hGQpq/k7InIOrzYSOlVFrZAETWJkP7JL2VpNyzR
EQo6n7P9GOwL6AA8aXHFYZFvab+pgP/2WOUyJFT//XQp7cobXYLBDuZVkYKw7eAdY/IJrSicO8JL
oqU7abJdWjS7zS7v4jcAP+YsE944kfa/sTOiktfYssEWi++oIG6nB1puCtsGvo6cRaByUj3Ujccv
s2xe0bAi+PJXCR/EH/XuQtkQEsFMBwhYW5TQ5XVLvkzXQCWkEFG0i0MFZ/QQlTBtK2wOmL6KipxV
PI6xgds0CkKbHQN8HCnVuOk3ilzftqbUnJTLM5lQs5Q8oGX5tm09Xr6ZB5FhODsok6BWyfVJU79a
s9Jyg28AhGjiuIMBvVCx+K+tJ9qSqK9IKfHWuTHuf8qfk2++C/xzc8hDdBbfZ1u59O7r3qbeEC+r
oDsedZltf3Y8n6+2me+yzD6wiMlqbRsiZ+ImfLfwhmn4YPQ14YyrDEfpv0K/g6MPwwoM0FGP2sl8
nUzbxYg4wIgUh5+AHW39l8uGC6cO+1xbfHKGHahdHIe8S4f+nvjt51NuKoy4KUIs/mSvW7/cJl+W
nHlm2nn8BDT35W5mRrTCX9cVz0GB+e17+9ec+j3jcWcwSvQd1IfB0EJfyLncemQpxoHmqTu9QONz
giPXc8pCbnUGiqHgglcwOai9N6BVmzKua3hbbVi693Sv/t4vAfOPDPA78geU0d90e7OJjOhLAm5L
Pl9bP2NGieAAp97OLUJe9iVrEmqxJi76Jn7paBh3HOvzWj/fyNCK08N5mNNlsmVK4nt5j+LUXSvt
nrKZbOAtWfJ6un6Ex7dCsnR66GOPaCHl5Joo+t7yp3sFGwxOlxERe9CXeFCSTY+Fg12QGuPfR/Vf
FCEC7IngreEyMGzWgcW0mnW1RY357Td62Fyv70EJiWseumi3/KKLJmA3dQwiUZCw2f1q2XNiRPeq
6KJkZJARgC87roPtl2BEAF17ye0mOiji/eDTKbcvmKlc02nSuaWDQFVd1rpxIcCB74n9HWOhuK1f
PwwdGyBtONnuGULClo7ggYOQ3fxIiFerANz8nAmvu02D5X7vZACRZCYgcwlMcZmcHk6uy5FLIqk9
o/S8LFG4GzW6vGAF7iBmIfsz9+MaDEI3oaa6O6Ki2uVmS4odKjh3Rv0U+Orsso7Ip00DsuZ3PFXR
qDz9t97hHnP5g1mCvhvfbPsXN6u6OBw907OpNjI5n4rNZLTylecZjWg2ju2j4EUEcLB93iyfY8BK
auEZ3blREBL7vZuoOwYa8GwtwPBP3XXgWDCrykI53AsceV/XO9Bwq7aaPBOZ9jPebCPDNTedTCtx
aFC7BcmbqyUi4KglBy0K5GIGLz7+/nYMVuh7bSjOQPX5QtAWpHzvYvpvx4Qtzss+ggEOwfjYqo0r
hJnRXPcgY4eu+XT3LhXrd+60dNnMObTOn4Zqb0toIboQcSCmK8yNo0923XT3F3Yd+mDckfM3rveI
sbfhwgXzeYNg7R6aKiaBzboqgO5xraJfgz2lNp9Ut34zcuOZt1kANtncWYIaV3jDz+UiL5lobPad
Y2BntxBjyKXOuLUau50Prk/ds2VPASuI6Rpy7ALD2qHMSEESrn7AOzzOYtn2qgtdxo8UPSFXIIec
Ov3sYXL+Vi+ycyoDSrJs8KYjkJ/EttkMViDJY39KHZ/Azm3TIBjy+TO43qcSLoDrsKqMewmQEBTT
7gPvT/F87YcQW4Fuj9uOf9ToJuuZgM6rM+X8DLCr32FYF8qLXk3ZRnjB+VEUNH+7op4m1SEd2Tug
EF2TFnGVk+xDNEyn0LOmMgHV2APwExZC9sQrtL4+HA1ZMW6KbMrExtJGViuNrSxFI4BCKrHWTejz
Z342Ica+qBGCZCD9hBxebvFoyLjueMlp+pCcrLGuwkvElW1GKJ6Nvcwe6+GJeT8kXwLYfg4TKu/k
3mXTBBuhcoRng/20YWDk6D9dLXi1xwAwKArJA4eT+nwCioD00+vpKa3t6ZKYzQuJaIGF0JNo9uax
ZQ9pwbGGv1v1PSMRlY4/P2LeEuS//XoI3N9ZtGlLuPC8zyn/eVrNCzt5UVAykdyFaEoQt+8X+zpm
3BtQookc+FQmq/91b7MR/c4bs/i5GlNL7peR0Qz33mkf8XgmP8Efq4iOB6F+8H/oDCpnKxkkKR8r
Oqkv/BGSIUXXvpWTwlguPtcX8akxUa0ZmCxbr6pxYlpwQVkqAGjsIRMDCgtalNFgD0UZJwOm6fWU
B20rXRyRNy0gKNGOIfC7kpvqg/kzP3MztAeu2GJ6p2mMKv1bk2PU1PmtkmNA68P48JZowMZ3mbKu
n8+X6Sid+MW3re1FszYPchvPiIV1s7K0unkO1kVAdwisxQLOYfVKpB9j4BzrGu4/kPkCV8Y+Z0nm
WzoyDfVjgom2K1csvjECCh8BKNsoNLo1U8sX+5qm8InSQfSHgaYEpRe0+uu30BK0x9Q7NZ4CHK86
esQaVnVSh9AkjxOGU69D53mtMqizSMAVQlXEdDUeiZpj2dop2xZqprvs/gIoqFGRCVCQHTmY8ac9
5rL17GD3xHm6gIRCIIPpl94jbqhZnVaQ3NxDuU7/JPfzseUlTQw3Y6GPq1LR5kghaDsstNzs6T24
ixH5IjlCpgeWVTwotXN+ZtDU1hr+xU0+vzV9DBaI0Wu5yNGlt1Inp5Bq4tBtM2A5MT/aZ3yMF+ou
pFkLAOKH/QAGq3nYHGue9GZex6/C7l32fMGF4nYG9opre84J+wRoL7vKspi5WAEKTPX/FaUhqgQN
4VMdKlidoJv4X6v+Mjq61jYOn+Rll/GoHmRYgAK577QZmwoBItJS12RH/kPnbU+7KCOSz0WCls9M
pqh1VWZ/o8DXjmOHrKIdKhZoYZNfwY9UavpZlQuK14/zZ9cztfuPJR7QHTCJckXokeeu10W24o/i
8IriARVQpEL/iQsoErTZblfASLkGDygIZkqWCdZxyLU0bY6yMmijhQtctI7vGzqKgXRqJpFHaeg6
J7y2KhIiBzrwB6L9yuH17CmQSDEdu/dRGzC536AoAtYKkCQZ25lf32x5daBxWSFXz5qZwZwkXGhc
lYcre+R4B4niRtZ9mg/sb65v/QQv4BJEc55okyu7WkpjAvlUFZsvBkqZ+jO66n1pMEVMfAKbMAfs
DwpBn75AFq1saG+9f3IXwyXDD37YurTbYs39a5vVH+kwNUXYbIQjlRv2PvhiXwxF8CPQZjNtVuwK
KDBbV8qyimV0tzcZfoZix1xFMDOfJAYTFjOuCuyavbyEbWYzhcFF0QTHfilf/MAMYCyadCkqUytl
IuoKqvJuyog6xS2YDeFejKrJamQVEwzFxbHuwJ6095vifHXLhchr7cVQQn5WH1CbypOIOw/bGagQ
1zyKEnJcW2f1nEaZO+b6Lg7RdRKwfg7nnoe2E3IHZ+mFtCUYMOiKux2Ssj18VORrIvT1cKAQizDF
aFDAjh8NDiPWOMTo4kOd1B9hCFHxxLYXVesjZfwkwtM7wdm3xrNjWWZ7w6Y+JCOueo/vTcP7LdCx
wnFXYkfVkkV5BjGbNeFDYbLq1iuXSa+VIT72T4+ECbTEJgaPzKQB/gCL8aWQ4razHBBtt5SxQh9T
HgRXCIjxIrSXwG7Ys/Bc4DVqkiv22vRYmKzX3T73vMyQjdB42lYCYM2MhFsK+Gu1HxH2KdvvIbG7
gAW5xFG/fnXaV+uNUMFn4Q7tMhOb9ejQd8mM9YIlvh56Zyr4OmjjTYqgNdfPdeh0+LqGi7S9Nnxb
BzUmWmVRR8/YhWEpORGP2AFhHqIZtdE2Wj3jDdzZ/5m6UdM0+L/skvwZRfrAb3g4Rr35L6TAQfJl
jUeVNSy+DgvwIy2YmcSEGI0S2k97XnIEcLIytXpRi2mxdTYWehd2hsz7URTBGlVR+bPBaM7szvpL
SwTDobUfCVI4lb/gpyqbW0K1N1lmVGyPoH+4bsBFdCFzdO08xvRei12OF72QL/DmwkbCfsHhp+O6
ys4uo1RIPufmnwxgKj1gOSpIs84tPgf3evLIZkU5L4NCWSxdtWVx9y+H9YAI/D+3t5zym34wswOd
yejuAzoxHGDI/ElVwm8nCkfhT+3FcdszrO6k0CByZVisXcOvSSnZV9zpBtn5mUD0xKJdu124GMzZ
hgM1KOS3hLuAc+nTbWksYxy3bBVRz+PdYS4FgQJHRu8Pr9hPfziWi59YAHPRlrmlkQORJdlL4/Cr
ORRJk5Dx+xRymf5JBIKK0BRgggNfifFNcvdtDrcfQigoCrFDeW7ELhvuT3eUfEG4N1/6BleeYwOB
0B8JuTVz/84YLjMNRQ1RSdusdpgHuGvAIz9HHx43cyS9JUGWrxEzAVEvTO7KqH+EcrPOUnzwo+9l
mBeE5QH3//u3bOyL027LN2mGrZ3+xSA/tXmRuvkh4bmuqM/8/3loC0i0/UOXjJZHeFOdgQaVBreO
zYcPHkNdrDNLSNahVQ7UnQjeHcYgJ/l8mI1iCuUJw3wXJKK2dIS8YeWxgxw99yFiRmkkrvFhZCb7
uEMgjOeO4LCILP2kL7dVPOH9LGzbT5iJXt6JEEsfdMAwPlNHQ+GQH9m7YmBnO7pL3zRuqqn5eaLs
pHNIEV9onuw3PKM6ThGzeavPl8idBRoJuG4l6JnG3lsxdGOfIeyCW6VYWi48cYcLMyqQ+d3j6NEE
nc8cDMYGJd3DoO37wAb5fw/wHISIli/JAJX/n8GkhObWs7st1mfiUt15qHXPClzJ2G4464rjpbqi
t6NvGOzE4j87nPd53DiVvkHn0usNTAHXfeRKc+yyepgwbIWwgmKzPBH6tUbvUgfsz9Vad2KExNfR
Q642/IZswd8vcj62IWWhNXzbbU2xIQsSkwvSC4BSybHB1Vje/oT6lBJpKjRB4Es1FEdoFzckff+k
ePIkoOOfRKnuLKFCNLrpzlqSR2EjeYGrAOjhJRjnjoSFUcIDNPixrteQP/Fos/2h03SwFnXXy56Z
G/jwt/IDkTI86/YqabFyZ3Rp6nB2ondjR7t5haCPq0K57q8tRoUiNONzius/EQHwhiKIA7Vtn7S2
HkKSmwoChdBMcihcAAyDQD+cEqvPm7QypiPNID4HhtYJsSjEvVq4j2MgZSiy9LNCtrLkj7sO0y9q
Py1eXeHTnRZ2nqrK+3HMU30+6J/vChlhkV7gGSpN283OC/oiF9ZgmlOlSNLcJr/rzeAx+ZXVSB4d
b2X+a9I/65Z9cdAx4F8l9iGCN8483GA29zk+EBIxWc2e86Ak0LT+cYm2JHWOo7f2O6gfoiG4I0DW
H3b9lZDvh/70/Dg0XKmUW2twSQkJFyuhxTf5AlOndupYt6tWuTee+s2EwEr69asB2gYnuOqW0NDs
pCirm64ESvcd8/c6dGB85d9kqlk6JVkdtzkvMGptjP5XNNwCnV9rkJeRGOgdVR4a8IULoTy1rG9Z
8BtoVpswggAQ5B9BA7D1VD7ESA8fVvG0RFMkpWZq03R06LNg5Nm6cc811BFQK3IPSjtkk8FZNPYf
lg8hAHCay5Xcc2iZUIWKQBgeHFozfsxSr+2s+/TW31DHDHbgADsgmapb1NcWA1sDEvV0DOH/BMWA
fWN61fXrZeorqCjnrf+//5Qy7LSsLwiEyxyYyve+FIsL/QLY9q8bA9RnXIB1rinNDKhVgJROyqZB
psp3ltczUBhHClRolA6bwLMKyyZDbZtYoVbb7EFBv4zmR8VRC3GmpS0psNOP/5pv6RG4WKSQLQGc
UXCknEqnUfVpYkKYh/mbS9KTYVMN7wqjGR5IS9aQfs0hmeQLLqbWwPg2Z/8Xd4zYz/L2b23qljTb
Nw/zLF+vHJavk/S0abjpVxSMco1gmE6oKyn+/tZoLS/ekvZZprCd49Chir7Hq1JqGLiyre+DVSBd
7xrmwjhXXSrJ+GiNW+6uEH5/coYGjYh1M4CBXH0uDItNYqSCXEeYn/LdcCiY0WhHzL0nrzefh1H4
5Qh6am17MhvZ+DUIUg+XxXrReJPHNoG5bdcO0zxwwZZeEq516uQMukXamzWesPx2KNsdPtUxJnJc
W9zop7AeDEDUmu2aiNEdptf1R4FmUzwD6px5ZJ//RY/sus7up+hP4YqEXFXy9ryeRpeUx0vCMgaE
FR4d+9AlYq7Nfeutd2CRsA3H3w5cvfdUUjJ/MD+BNaQTgYUTGN4jlxPpbFPtC/2PcRa/IiRS/LG3
W/WZoOoo46e1zf16GtHQM0jcUwDBlZolexKMbqlfS9Ne1nZ3BrUJhVwVGoOT5vdveG6jg/JhRj1a
4Mbb0uEB1Qhw+Ri0kn8oKBarAYpAWbBFMz2puR7brVYBwihlHFRbMDTDublaRzXN6QAkMTYu4bwM
9cdY/k+CWAFgQQUWqeqUlC7/Ep+jvJREW5yucLpd306mBqdi502OgSaJ7LhYgtClpFvDvcAMrmBh
nXaaq4RXICszBeqfuMcnM6PGfoSymywY2UU9QyhaT61EMB+Q/90oBLoSrsE9vCB0XgPspI+9suf+
stV51SXHZ/nScS+b8gWy46PhbTYoW0lRndgftPOIduOBGin/KtkWe45UIiv0A4lFUNYG5FtntoNp
NL1SspQ5vqkjCcRmycTyjHB5ysTqZC7ERpqfXLJkICmEjpNoOkHLvSSGHj88YW3jhEIJ8JuFDwYE
TWcVDsBkGR/Ue9Izqe4O08Ae/PXFduFS+PmfQMB6VFtoRLD1Nlsy3h3eyhxZTFsZ2C07mAEL2XGw
6v9ojfU4mHkmziCRIW/XWrNDdiNjnH7sp+nHtE0kJKRsWDj/8mf5lDrvZQkUv3vjSHk9dp65NR9p
VDmLbxOkUUkItOU2wg0XMUCv7h/zzKE4660KmVJpF1G0K3guf/qnlHE4byfAVJ6VI8yc15cD8zO8
qX8Ko2JxlvpKO1dzvzINxC+MuuoATNQYE6zmGZLojIhppb1vC/9cQ8tQjuUE4dpD913K133YUCVs
bnB8tiSb4uaAPgSDz9EQ1k6Xlh7rz4tzMXH00sN8mVK5p3sHTJHDXEHKbhwmkw7pHWgZ3+1ay4y9
I3cO734KepDCD352abDnth+mDI1Mlq8QsCuK5YP9S2ZRK2Ctpyel6qP306bqWaJ6UcFtc0c8dfNf
/JMMwouXXw9Ly/0lBh9aEsmrbSOXprGLL2jZIBtv4ToS1CSgW+1+Mv8fa7SpF3YgmXo5g3dgdH2W
9BF1sYuZVWZtUxWY7J7ncU5Gk/WXLKtp6AR9wJXxb4cyON8kJcrC4zMD/covs0HN+xiIztajwtjy
EwlUr3Wyyx3KmlBJFZtG2jUkM8SK5d1hoRyYN0Ba2jLQ0fbAeJIk6W3e3dkq1YDhh3q2K+yekVQG
vPi4/aI3DwXRZjZ+zAODcSEFb4+S5yOFE0aiNkP0XzteN4n06RCqYyX+Vll4XnlOAFR8HBZEI3pN
PbmI6Th2f5P6J2zG1aqJEZnGseKD9GT/3S02/sq1yfJsQQ67KK96OZ5cJcuC/cJTWvaKPXVI93w/
YHTkJOog6jFczYaLtlDAQPw9jft+I09yZiLpjd31pYwImLYHfAR58FTtI1fmyKf7v+Yl4miQjjBc
z7G6wzwBflHDecvOc1JS6hxR8CO6eDaT6zS6+jYM4El0IHR7ouSQc2/SengKW0a/lftPxHKpdK38
Kk6fEUsW90ubR59BjKEJz47NDxUYdQhlrnvi8LnDDesWlkt1mDHaCS/inrk/3+yxa7WpW6FHDpie
LhXMn3wkFQyESb21jvuVL5Z1l9MWm6YW5XCThn0e7Szie6HbCj6AKbYjcCPmCzcEtB1RnRZc80oy
ugYITP4tVwicW0TjdjXckZgLSsg6mq4m0jrZRCqgXxee9vGhRW1cJKhhc66HpRZeA+WUetdxU+8E
nRO0t2H1wWzBaAMBPobPy4TUG5psj8YnCJh9dIVVNhLUHU2zhGFt5xewGtjm1WxAzOptyyf/brZA
DLcNNWQARASuA1DtmBzqUw4Gd1hXYhgNleY1x2tUeg24cQ4wG/wSI2rzEnQHhcF5WHJwCDfMuGp6
f+G2AYZgtUuZkZsRH5rjjm2FzCgbsb8wZkehI6sCzihMYkkxyAB/ArWJqrhDn1xaQvJYCtq+qZZG
zADr5qV89e2pvlCbrLnvwbICaWbYQLYRPLdkUKrShAlXqxuooPRGWKctwzWebi4aXdJ7x0Ixmo3p
yq/KLrh0pDlQxvqCN8omNhg7i+GhfSMdP3yNp7CKARV19zCcY47wzekp3RQbZ7jhpJLvKE1N/q7m
dTAsZld36ZjzjnNnSpL8mDexHutvrGR0wkz0qVj9pmexfX8yOQ6kIgZD4iBsgXWyhiRJBHrND1vb
mRJH8O2mMCgrjQEEGYIZGV5+dXo301J9Z5w4Udjq+4hCpAYDinC+EbbKxVPdgo82nWQg+vCdf+hp
rIvYcCA6tKfExCH3MUhmDSg6DXSrownWdKfpmsjJ4yTWfX4PoOaiLBsn19dRj/lMtX75LDExDcyp
tA+8zNrWz/q+vY9luEkROOOFMpwttbKUKyhwE07tdM1EIZTXT1eyYbVkG1B8GGmZA4ByNwwNKoiT
z8c600upJ7fmSFWvHin8ikHR7GEXsXv1a6wguUu+MZtUxi8cUhdMm1mOg2y7qF+p/E4PcqbVJC06
SX/v9vSfoxzRgBfiKnN7y/3QsNAL78JejGl89T+K95RRU2ol7AfFjaKfFEtF1SSec4SEwL7hVsoz
tNCY2b0uJZNAgyQL8bzj0hM8Z0sLs8WKyHZ/+Qi+Q38XptQLDM/D0Y0FMW9O3xpL2geMoMblZQjK
G8Jyzc6ZHCCjBGpmNy+3jFGgCNtgxXuobPxOjpbQrzUCg8G3QuZ+bwV1QaP/DRqP2Iox/q7r2C1g
+3UjgSUzjSPg+vKS9Ok70ty0RJx65HTNbPPt1JgickSxvmTXDpNSLax8vtEEYIRNYg7pCZ1xy+Cl
nGbez7qCIakWQuR1ekoJtvrgA88hY5HiPSNUukBD/OGl2SVTuSrqXzMJ6BH6syH/44ZUjc6A/OZy
JoKXZQ7uopa7Hof4vA66JADzsIkd4jkvknccTsapW9ih0unlG8JFowOg2pzC/MSYJhi8Pjpw7Bn1
YPcvGDp9S+ByKigk1iLRgWtnXczVDgqwheNYNF09zeFSaUCbeMrspYlPnSVVesXwYnm5/nGl3Gp2
2xOWrwux7m5L3f7WKoMBB6/rfwnWlNDmJ7bxY9VlKk47t0jRu62ptswzpSsQGmUBTix7oTwww9jc
wgITzbSQ3ZbAIdyHhDMJFHMQKzlAJ5+1jjtSs8lhw8M6Ssmu+WRYpTvgOHQC7V1reDAj1sMtja6K
dG+WfhjCH7iUi8OU8Rh9s9ti/ZLsCjXnrpkh/0n2+ZPUpozee4n1/qBMydYsWyCm1Z72nqNfuuCe
9OtdsiphZdmhPD4dzdjzIHTDYmOqZrkvkxEA9Sk052Kjbh1MpWGme1oCwtlXYA0sKJXv2IoVlOwa
7HkzjNgASd9jfyBSe4Bgd5Y6uwaY3heAH7YzVjcij+9zLx2N9QFt+asWvsK1iREWez9LU0Fr1Ky5
wPOV51PlGVMGcpX13qoKLJ99S0QV7XHusrSNUh7YYqawoirZP+CxsXEkFxGYzQdJfgqXy/BBijKj
2qwUZVVIUcDxKTGtoZsWM0750hQlStSFf8SC8QaePLdjSBjvHZh0L38m5NELR090E+hY9oXuldUo
pBV6DwSYTARWXgN91mCQnTF+9gyL8LfyHQZrWzyvXJdeHoKz1aeS22iIdcuelv/485DgS+qr26Dz
cjlSQDAZEzHrnlo7dsdtyLrh7wcvlfhS8AYDSaKy6NDJMIgN/lmBaMgjSm/Ux3uj8yHSU/Y/92PY
P33E1uBCMGEO6foa2Z96W8Y+87oCFrDz/WrerEosG3yEc4Jxe/g7wqlHh6YzkxfdGawt4s8FVsg2
JjC1JvlgeKt4AF/SObU3lAtm8rWtT2BAnLj2mXA2HeMszhY1SFeox1RikuQN3tq4Uo0ki829MylZ
wrzhllZCNF30bc/0jEkMLk+7w+A5f6IYKbv7qcDKsR4ykskrKvc+Y6HFwJspya62lAliHOu0vXsX
3ZYP5/ex1i/EuYQdABRVZH6Wu7SXO88/n6tScruCq28eqdM9nwlbHvdE8AXuaPac0VgDX1IgZECQ
9aW1CraI3WSAntN98GGBILr1an4Jix7JwICXbD9Tx/BzIaWdFWVr44XMl8JnDIwM0agRtFE8XWFm
MQFTPVerYDXBKOPbu4ZJF0Dbkr09vAky2+iA9mXhb4ZFxCw+SD1guRi09vBROtsxl2LIVJEgw/jb
gKwH2UCdVPgWibHsIwRr+Sw/pqhLiK0hTZjouv/ZNZnifExpJcIrJQU0ZyiYWcErTGfqTXOuke2a
fdQByOUtbucKQ6lRrCBmpzlYQDSIAokqIax5+kd4XWsAWzuJpg3vCV9pXqROTHPbELlmariE5FSR
UohWfBlkM3R0uVYV3adUWbppo2bkFSberbJdVxmsAK89VVmWTdFOAyItV9XFc3eXvYt9bTVcAmXq
L3Ym0Zj1Hrm3fY5TzAGsyc3VmgyHQYdaFA+1Ls65HJ4JcXu433M0v6sxur8zzeGwGgU3a+hE7Q14
3W2KvnpAINOtfVOaIFhn93uKxOTsNPw8lhWePKO7IRr5tLDPrgbif4mVMgKgo0anSykhHBI+oqmk
POVWApBCkWQ8Eajpzts9zthdWib1jRBuYH4uJZG/BMv02IprnyPS5GiquojYvAl352mlBhdNI7vL
+L4elkI0qWQcOT3Cz0xChb5mZ2EGb2Hb0rNzxE1jPIPJ73ne7XwKARNgeNWNHbxtKXVrT+mcm62D
FEjRt0f5DpeVqEEI4OCPoY32sMbrhMHNA8p33nTjkU244B7iPgOfEs9OBZ+oAADpHFGH+aSuX/kO
1+jB2qELZIsKf/vNxu94Uid0t0kA3GMgtQp0UARManxEgYUmcYi+kw+gnPILa02A2zrdl1Zw97M0
g0tQ5Nna2hT3WJJ8OtjoHx+ENXF49NL/IPMpRihRgpc/8C5mLXdYSdEnbEF2b+0ZwmNDMVbQOdR2
+CETLQawi6g8By+tn0qn+w/4u1p1kaR0j4whqr/cqiZYAkfxgfeFKxu9j458e0q8dyGj4gBsQOzY
HsnDozAGyU/iGqRzmKvs7tDPFJR4UaMce3kfSLqNS/oEhhGMgCDpdOLTIj6sesHN2kF00BfeINEq
kcwgxPZfLEGA4eRP6HLebR+NDQHVKKZaClANS6Ni8c34ocksERfQRFlkMjbwNJDv33n+H+MX1jnS
E1YviwQrm2hRyaFfyzWpPZ1uiWketxD6Zt2GgrY7yzZmQHqLKfglRFBPOVVwS3Qy3UEtvrkR51Qr
CERuxdrnll0qXXNwcWRyGzKXN4mu5RjSgOjXJmfe8/umhI8O0ty6GfVv9rOAfZnSsr29kfg0pIiB
TRRVVPKtuJQx0ZsDBvifd09QipxaEueY1OQl5EJXGab1kWn1kH+EhAV8Zrl1yJQtx6bI4kDtK3bs
X8q9pqcQE3rHOz0XLOJEragKKmjTJT4nXVPWbI9YQ7eW/TZiedWZDoCc/IsdgMoYfVJDUKK7sgXe
U/qUHjOfdHAghZYlWJ8w5F6i81+NYs5Bna6FQN4048o5R/ebMaRBMIV5d5bXDB/cWo4LikVMrD5m
HqzKf0q5kdLeE/VhRBeqpScfNqRfzvM0QRHtM5SbszAyJvmk4MtaXwe6Lo6/FcXT1AAOc79SFuoK
K/G4tpJo0LdzL90M+ST5IzjKQlune2CAlLB9YdG2/Prj0PULuE/P77hCRIgotLKSWWSXG0L+jYOB
W6sEA+UmgnCgqWc0E9M/JaWyoxdtvXzFeRg5x/4kVLOuA6RxV4RctWh/uzVo+QwEVPiA347ZmKjB
K6h3PAiOSjOgz2icnH+frUWM+pq/EbKqFVGk9f2REU4s1mNqgrOOApm1InvdyoWeLPs6+SvGElYH
ISX0+2znGGaoSMiTIpdtaFebtwIH+jHsNbiZvN29cbsgK0wjLv1TM6+WcPGo8kyyYyHs4HHcctI1
BeIBxA+YK3XEhPKFEr1VPnJ+9TZ60eKWY4a/om+BPYYIW1/QPMini+/1hLssYrZVyKrCEIXhH5gm
3jvU2PkjQs+wpzjNZPcAfoZoo5GqGssFxG4utgiUNX/+goTBQtdWVDpX07BQpu/kzudSPbr9Hpml
U2cu1ro0S6yu2zYgWWk0tJV2qpl/gX0bj5zx18gpBkjvYMS/OdrEHp0SNg2Rq7AFmCUbQ5N01O+U
MGl2ORY7NCSG/U0FAaRZCjn3rX8IJc5Stt7oVtoWELy1p1/JOLNp0VwagnOxn8UVUIyfxEYRJO4w
UNt3NHeYt1Y/lLMALaGURXopb5fZJ3u5k6RaOK2W3Vh6LqABHWSmGhOhGLuoW+NbzcY9uNiKrgyX
YOP/CwSIt+66TxDwVdK2APlGH4y3NnunNBRhjtBB43ouotyK0tMpQEl0K2HEXV9bNtOvy7E2Ce5w
SaPXDhiQoxzbIidrIZnkCqXPoOG4hTwCnFp6ahVnyZvWH8FXRdJAOv10lKcOJJ+nCTG//oBB5Als
/7j2QmXB+hHzBEzXTweJIj/B0MLTiT6AfmOFxwo04FfUCbaBNF83MCtVUm372CrnI+zmxSeWWBv8
P/8rvpiK0x3o1jrbVvrSo3BfJy+Ivg1YE2nCf2Ud8yD7SXB0LdVYHv7s6YLw/7IFKy3Qn0ebzbKt
Z+82p3THUetKUb3+LawDa3kcWk0+tBADh+0IkDFMgsR6Rin0N6EsD0GYB9TsUpmvCTp14p15XpEI
DhgMJMjYPkUcuZrIQ9rkQAts9dHUMffmSVoJgqgmIlcshmvGDK/fkpqkjJtWpO46oxxDs9We+J34
qDHZfeF1HCzDp41hviRIQYqJB7x6CT0gfRb3Wl+dT/COnZDEGDVDoUdjd4WhPyUSWIJ2ccKBIFmr
G7BXFPIdMNovgaEpGJJMUlemd9Kndmtk0zdCBpq9SRXfCmwy27525844q8xIeTN5YOqrj9eVebv+
QQvUMTByQBGMIeFIOIo4U4lqhJuxHNJVF4d3Lb8zVgBmwWvwAMbTaSqkSOl6G5T7l2gmBkf9wRnc
24q4C6MOjCaEkkZ2l4denoGaDa3HjcKLJHVO0WvCX0bIFjjdVO2O56sxG7FNW8gQVMkNBB/AOgdY
eHunUIeIm7GYvdJyDwGbTAzKroaKDMvDOJxhfxqsToOg4WzhjaZiARTaxXKlEhSIIJ4IAKRl7mQy
hY9HsRxBSqm/Y4no/h2PvtApHfWOoijrT2noLNP3iX9cQ7Ec5lAGPcoU1yebQPqTC64Ofi/JkkdY
eealKrUIPExGJCQiHVfBTWtWxanY+1Ftk3OSGOQe/eLgvKoSGnt973b41ZFCf5D949Ne9UPwjPdx
50nBiW78ahqSY4zYzd5GerU6SvHLl+vvhKW5W8fwjQXKkUL/FMLqeCihR05yyOIFYUVzGRgsJUvh
BVuI07zbOIRpbbk5ICDZVAh84JTmZfYKhXD1uilRyxQJ77A/0+7EWb42rbkyNKXsFG9+XPTQ/txE
WjMgOdlCo9Y5hXw1cUGzz3NIY1oH32PQ9aydYhUo2MaxcZBk+KeS02+ER/aDxvsponFefcP8Fppt
Fxk8ktHf4WgZlKfVoaKJvki2vD0hyV+WZ7pOI1GmBoB8gTAZ+br98irHW2BAH/LmVrExkSeapcRx
LPLhYBcPCAq4b4cwKCQ4P4wMU/XmNZcbeIiRRl/4CrL+eX54+tvhfKYhN4U+Tyy4ILBGZDpqFnwb
9UgQJWKheGVTjz3RzogfahYaBzv11OV2SNJxnEpzQnq4JwTBKLJDsRLv69tGbN3p0680ZFqBy7A9
JAYp54pdxbgkeHXMQJ7lKzHd+5s4BBYuLDKQe+hdr9D0e5cbyiyi7ai5rdw52E+AGQ+k/gR2ti71
uzc/0BWvh0pHu2HObjc1cbDthdMDh6QNSYLSA0StEdScYBcaYjPOk0gZu3fdVeo5ZFTx6wu9biTM
7U5QGN1MGXmBQUzhK5wW7JZ8XMuQ5CjDt52Vv8XaIry89oTx6BnTKoJ8vWfyaqLIb3rVg1kboJgr
nSKDc9fXIxWeZXZVT4rBaZXMnA5bDWj8cHq6kYxOWZmhbVk0kJITbl0ZRHeYK0hKCcAL//zoKQ7P
JmAO+gpgNz0WTEeoHJ2z/E1E5gXTBLyWDpgNPqHvRDBWMdtmltT2THiGGTD2M5wLFaEa2PDAfdza
udev/QuvbWCkC6W+fXjVSFv9u2adCf489g7mdK9PLBHvrGJMpC/QZBdXwdBXPBd/5+U+MXglB2lz
qhn57llBKxH4Suq3wxci9TWGtB7fDM0u5F65EJ1CGYGgDYcE+jPi+OcaycXnoMJVk9iKOloTs9oX
AGNBlNl/f3S7DzpXKFxpi6nkdDPuRgZK+TvHFBSWvtr2E1DZrqm7iyQvqZbzVYAAKFsATxHeXor8
lnDdcliajwpZcgZTm3bkzSkGv8cIO5+3d4u2dIRfTRKnL0xKOrEqMMogKTZ5sTL2hl0r1+mrWe+m
dA6DD/GGzlsQ1olkE/cHmmxCpPALwovqG2kkLtyE1qH/KOfNrDCqidKGX+/WNMRjbxYNYhg5U7o9
UEuHWSZMIRrj9yRo3yPOnIdtwfrsOh3VcFZwR42YiLcwBc3oTxACi1UUarishqrpGxiwFWaIgnBX
ypCMbmC839vrTGgTACy7hr2CGMDhIdKZAlvtrmVC8w371/ITwjvuzoidLHlCkz2hkqzVvMhxd0AB
OpMp8vWwAcX2xD0JlOGAifXF/C3tw64jvqAL3Hx+lY3fbH0mkWQUTrqdA4woowC9NUK3/4esFeNc
2+RsHvn1rvC2NYATcq/PVUOzdTX8YrQXX4NOJs6Q8blORM6MVBvscsbfm8FszT/S/SKshT5J/YER
fEP6NAUFwbSQDm3yOkDjFSadO2+z6e5i5NaxTxnmvVjcwA/yM+ChlVtiw7gB3BEcRnrkEA2mxKZC
JYuFhLvwDZqAFakrZkqWqXuBLwLg/sgqjSK4IvDrRgK0rromAxJIS5Q+fRqXLASNXjyEyyUiog8T
L8dJaPfjNeP6uJlBZdNcnX3e4ksbOquQLyVBkR6IKQXM21dLz+f3FYoQiDCz7WkRfvmY6tnjfwUD
au9QeE8ZsKXl3759w0uHrwzTHEWuOD4p150QjP6C5eeNOy5sAEYQiNezvM4rARVl3QSzR/Ej6UsG
TqaQa7gC/pm09k3KkLH9Vv7a6o4QELpciMcQuYawI5Es9P6Rajg5JP0MdEbspMLcF1aUS0/oHCtA
SfUrxCZncONtAgjp/DuJWDwAyvw7BxuR6ag4pgt3Px9SuJJdg/1Gk9p0vfYvJIm/CI7v5WnADWAz
2xaPTuymGoF75qr+DW4MlgAQRoL9cUnmWBw6BbVrCu4/yGI5wrH3/wVU74fugvspNXvOh2wNLhH0
XxOoITHLkQEDG/PHfGbw1/23GuBdC4SoQpiee0ZdGguvNS2pzdmjLIEZ0gzW05WN29cgJOcdrpf2
36fnOfbQCQCjXiG+kqhiiRwBKaSmVV2pWZUUTv8DFNL8Tsx2yV8EHs5HGD0mX0xKYfZgvOnVxQ+2
yJHqdGr4ywkglIdNzZrP7P2eLE2YbFyQ6gL8BF3UTBOwu2HieCmxKhT17Pnez1/luXEBkGqZvc5E
cWmjEx9FPH3NN2/YDBjdSjphtXbE6epOKXl9oQZM03SGpnQ/SrQ0Z1j1db2EGV8WsQIzmXHP8P2U
H80n4ijUyx+EUARocvB8rVNVSQe//QrEDppzYQ521i8eeUXi+lg2gSSVdHHfxscYqXJQBAuyBzAR
SdHbaRSf+r5aqEt4hm/S34YsKCOddWhR+qa7i+3Q6pVD6MRNHC0lsBMAhOr44WUSEYb7F6QzhUdO
w8OOEqPcER8H2tw3MxXl2O9OZz2HpAxSQZdaP7Ox34Hb/LGyVOqVc8sdRK6RNezHEcu6tKoQoQaZ
NqonAnVJums9OrowJfzPMW5pSf8T8gP73tYGdmuwBqm0FyR6iNT39hLT6gUSAARHZWd9XC8s2yu6
pDyokG6exvYgXr7JjI17xSdYZFtLRdoTbK+9qKFVIfa98dz/xtK7IG30TkSKSMeLLmd+moU/pkDF
FzHg3Z2TCkJCW38eEoo4NpKIHsSG48Le1GiY6s/c9vWtjjPGDHh7pc39OzmLngsarJt/mnJsLqDP
eTUQELk3EvsFhZb8YFDODtJwcLwLuKDuElq9BbHmUPLqOLPvnGRr9gh5yjtZJuldfcnJBve0IIbI
VavMu5qa9RDs9R+2+w4MEt7QIATkWeHvmNjU1q6eVkrpNdesGto9fvFCpzStkdgTY2DpmQL50nby
Wjjqra8mlgXwY3aAVAJA3LM6S/v0vEAkPadzx9YdEnAzotJ1bLnhQ8xAl+iJNUT64z2XwBvhIm5E
uTZ7YMbUvo+M5HgIY38J6UfNZ/BV+rBe9a74PyeWYU8IlcYqnkpwwVaxjR22w+cHwZ7pFzI16am6
9ndm/rZ2an4U8md7bJmOTEe7G+TdN3jNryP8BO2bTK2MM0adiQiui0Y86CPKm3XP+8wqAqHDq0sJ
t7M3PjUM6dbm3DXoLbmWdzxyB+GxA/DoBbdza4/P/+AX68YwicY4gKBHhHVkbGUxeLNpPyyfXrv3
JbxzZ3MEHfbX76o5TWI8t0aXw00XEH2OFD5RnL4g3E0dxyJ9UrQyuZwkYQmsqLiK78cOFfpKkwKu
GDk9W4eo9PUk6xexdJn/kmu4z4bzKHg92nF15OfHGhxquaryAZ1pdqlua4r1DwZRu2/9WqWCo8Lo
gGdwieNwYoE0yIMAiAQM9GmzRwFaLvfkLOYPjJpi3AZOXwWriF+foQe2zpvB8Re26PLv+ocGFGRM
QgPDvmKTSnCfJlvXNil3SCRcM+lrAOttW5nWeknvPU4wtQX/3IJk+fGDfH1NkJ1GNhlFeJCgARES
ETHL1QmG531RbZzAbFI7/DcC3BNk2pO8F4xYcf/JYPygaJwD2VUOhSbJeWDgKw/cQIdOWal0Pfy+
1lwRfWlOkAK3fK4GRftRajAdF0qzMA+bF9y02k27XpGPJSZE9lBVSQVbkPNC7JJZbHBPYTKVR65O
udYraPT5IXCVp2BzG0ypfdY/W6WmcgGLnA9i5xrRJetFTmMuQ3cO0Z73O3SE6clKK3GsTQqJOwmP
OUhOEBVkdlABDd9EddzCWVdxLoV/5oXdkNyrCg5CDwNizFivQwiokBiduErtDwVS/xdU66blscTj
vHKecx8f7gdYA9EHQutGKgc1o42s2ygdVRKTTQXlCHAWQs+9vIHBo6R7MgPBh6v6Z7A/xOTceAk0
1d9h9xGuHukA9UM1MdpL1sts2iE8r8wLuXm8V1n9CCYi7ZVrvjzItyVICqFw1zyRd4JithlfeWs6
73CgyrZI5B6PaTsAhpeHwGy+7+G0x59zhGZwtClk77DiuIJT4XdOHZGz+FM1Qf17EEEDrld/smpA
clRQE+9ruHNN/uTpk96SIDtiwZvxFl9VgFdkjHHhonNLIbmRtKaUVaqC9jTOEoviwHIdwpvhgJIR
6OJk8QaTtctTqVwUKCNYIjTFktVNHDEFyG3ez4Rnak8MecJTbqjzgQ6/fvBOpGMqT6o2LQj9MnA8
RJIiWDQjx0q3wANK657jncfPAkYYGbpsZEqLLqreCL0zmR6LQ0hGBQSAuQnp4VnxmbYnEQnrWsvo
rSZCCwcpqxDjffflj8j6rtKiIfmzSZ69tydrrykeXhg0h7HVvTTWEinx5OmWZyY+yv/mWWE1ygNq
Az0fxHM58bfkpSaff4IFI0w1dO6ylQuxKhH96yAkwFj6Gq3WW8MzFL8aKmLLDZNUVBh11lDsrOtP
D59y/+Zqehf2jcmNq0GFh5leu6u3a1rRuuKDwr7zzi5D55xz69LBHxGk0E0ZyaOJNI9a25XUvT64
eKVqwolyBFlUfDbFg0UNpPppxlMmq02DxOGGT5xHwuQs4qQc4m7UiCdwjE8qDtEivDb0e2uWlRoW
oXjzAg8kvo9mDjIpZ0ZWLysv7levBxe3o46xeoVh02jQpBKU3ldA7/vxFe0gDRJDZ5xLQwfc+QvB
VgwG2S08YjkuiHn8q4S+TXrAIj47yWp/NkdQtJQfuw15LJYc1lXu0Ldtq6F6MLgDJh1/wLM7TfUu
fOTwMAX2HXgrghnJUqmOyXxOWIaiZ2i9fzsqFUEBeeee23g2nCtocre6ZqIJOe+M1bBfUsRrkfEf
gbfyK/fZ7JQ/mZC9IfAWu8yGCKfJTZPDbgI9VP0/kIJKE8/QqfqYM1U9LYbxbUUuvasqI9ccsdGN
WldOQcrqT8Tv/0hf7IZMr8m1u1xIAUmlfMaq43JVgDPRqHG4y1QG9BIXN37bX6BytnFxEjdqUAbW
g5h72NjMsKwg/QdhTLkgGRrkwxIhF/JZbiDigXDsAn6tKvWIrcofLk7P8o2ppYHpqEaFKqt9diyl
6o5wqKRCz4mAnIj5FWGbvAD1w4Zpo5Tla5xV0ctbXCVf62/F+jJU7HBA7g0ejExhxqJ2MoJuhsjx
fWLf/7KGQWu6xmjoLdOQVLiG62zYDYFqRgn5sW7rrAbh6bO9KkCeZaqYOs/0q7tfzqUmUCqJOUpf
Np1cYJJtzY5FUmPaMSUsHKIHsV8zv+ociv+uh0TDnQwLFsCXmBdELR0TT5/k81yXKpOXTHkQ+IE3
71z03ZWCvCC36b59h/Td7FfLr5A0i/PIPwfzlW4mfLWtTfJn7Tfercbrzy8D/1vznEJ37SWWK7JW
/ttokgNhUxCV4HB8swHoT3I5j4t/MOrhIsvzY3QqDzGfCI3WccFks1NBDtZiS0KCCRLJYYM3NNdY
9tTi47HTNmEH/r6JvTZ6zgcQW0paclqx9TCq4+WXqLYwT+5kNmIjT080C+DoUtkbtN5SHV9SiP4I
5oA9CVibVXXbnwmJ2y8RBr60n8dcgRolcZzPeiVaXjL1yPM5E8QAloctlMJ7VPUDfZyJ2XfkdgmJ
66baU9v8pXpsHwILJ8ZZyetrssNGlGVbmFUuygYIs/FshCdyAa78ptsONFz8GIZTP20Dg3S8l2N5
NroroM++kVHz5zkRntGr5QstbRPCsXIH76AgdYM4OE8zXflMGGBzOg6ppldjDz4O4rcuzV7mjzaI
j/JKZJwoAHJ7tOd3KxL0nBN+E/PPkCZWoq8i/7QCZkWzKH0IERqMByFumAghW1zvc1KIzGwXiN4S
88E8hlIrHjT8wcOG7fNtt04myKZpd/ByWUQQ0lPOykj53yQgUoKl7Fu0xvHMmZgaGDEMtuXcGwRj
kxpYfIVP+g2wP67mW5okwnfAMtu671dEpCts2ksY2QVrte7ZMRB8BcnkCyiv6QYsta+shPtR1gW+
IsIChd4m2AU5H64a8iW5xz/OHMZc/GBQtxVQbEWRnXR0P4fxlUC8B3/BvLW8imKev/MpKQgliy36
/JZfeG3Pvw0xk73dj9dQfI9uKAV8bIRinEr/kdUBWRvsVaQ/PfVzwHy4jRhGpWW3rQ3ftWoewZF0
l8zW19zfqtEzZlQzfdLqYqIMLosNYz7K9G6isKgF3fmWBPTvl7MAuSXNJGoxrFpvBbWDC3Xq/L87
sXTdb++EjLnLF4n+zqz0EVsv79AW1c8YFjH2ymHe/DERMKOdjXBgY6qf4Hr4hWY/7n/ddAn7i8eT
00lg5FJ4hgTNC7D/Hkm0ZscoRf6VIwZdKT+doyyHO7PKsM/tEs3mv/x314a1HG0Hbblu8OMTYFWd
r+HfzSL6SECKrqBAsLJRBDRUc6hoAQ17YWPXGr/Q8Fi0O7U45cMxqG/cQiTQ1qIPd0a166T9CqXY
D6aNGdjh0Q8X0o/PNJ4cA8gbnUS3V98RcwRXmQG3KKRu4YtgcdRiLdeCzgMdwoxJStjdyiAq2lvd
3J4jNFBah1ffzRO8j3VEk8S8NECb17Si4V3yRAhwadnlsKyk8cF90FVi32lLvBhUDS/VjyfXrPZG
Zl0NIANvOpJdQhbIlQHDiTQleHRbcSbSAHWfKhPnAdRqPcviM+4+VN+bbyv8MbxfqcTFMQ3kB6R8
8V8ClUqzCcmWp3SkQzb1PVc7AsAJ7kTrCw9IGEJWehiYuZ/fDDnyaK8FulUENtR9BbZdGpw/pU8i
bOnoW4Q6qokydQf3uxCJYMn+Qy5IdGOUciZBjFfDR1t7dL4PcghxTQjib93+71cQ1ULQ4wWnuLGO
2KyyQ1tqGycjSKqQ3avmDh8Mjln9PKZSJKgaTPqZBkrXnJR5yZ3eIouZvSgxmn2YLhWIld2p6G6m
DrTlA4SvXCuATtw1l496uN7bwgpmm96tglVOCx5PbY6X9mKY9g+jEtARmJpsuTk7I15O8DA5maKI
//Dfx/cWhWYX2jyQscw2eySzfC6WS0/0X/8n99VxxvvF/+RJckXfUirUIpX3w+PICbaZYH8giCzO
GSywdK/VbaMIiZ+d4Gfh/JySUyhN7i9Tt6RFozAAOJ1E7YhacdknNFcmYnYb3U0yDnJPYEMbg77s
8qZBw5J+W9BzvQT3P9DWX2mSGYFX07Fcqtobwsyick+iUrmb3x1HyF8SEq+FTgFzVZfJ6VzqTz1s
cqG0uCbc61rQ5sVx15Sox+og0dDI1b3R97F2cZDPIdmpkYDNZJo+bWa3JAzXXT9tKQ318uz+nmJV
hv/CmiDOVo4rb2HMOrT1bF3cKBMrMQxM+W7ldVbDFZToDOJ4OWau1iq+7dLiBp3oblYxE/jxbF1f
eRwU7aem++sihb6iQRafd1TxL8sEyVYjX4Iz3pQGY5yTL7TPV4cCkZnk9+y+UgvvziET/sKut6YW
YlMHIRj99rACvNQs9UkPjsdNOrom7QWQsP+w1W3wwDAgOyYsSTCOxc/FDuKCN4exXawNjqPA/auU
kRLIYfQln0kSsnjdjiORHHPE9P9OaKD4adhx9JsQ5y8PhajHtslBxj5bQiN0jj1nSqg9PQXJhlu6
bnIX+AGBy/KcYfRa5MgGOXOlQW9ztdpjv0TH4DDGPZ3r/MlE0G7/xQCdbDyhsDYazxPW3TRk5PkY
y1XAyxPEtwJkmGquCyT/KkR2bU787zNbk2O2G8TYriBuKWx++dDj1cdn3m6r94QLj9135y8xaZvh
PtAqzfisjGFucgT9roz+AM0uvpNETPiGo2nY7qa3hQ4vjfBB4aEyKazrNhlcrLJTz06y3pEoPqU/
TO9pjyefgtQ7KfH9F3tcpr/8Sq7oyBZ8mjAswvOHYi/cBfFp+0Ki/ww6nRQd9O/aXHRUjHTOHASx
8KbdFY0jBwHmSle8gMWATP1VbdP/vwtG3GRNaUtjwFDK/mWQZPdovrHfcSpOZTR9gnrDbP9CieR9
sNlweW6XlACI8H7/O+badZh08f5FzH6Eik4ChT0YekKJ0IxEB1RrrtqUPlkx4HbGHZjfK5gIXXXv
eM8nlHpFqx+DuyOzT4rp8694igRnoe9OuqZkTmcPr4fRe+uDH4rRoTvmE9r0dGUUrnjAqG2v3SF2
sAIVcLYwFSzTNiC2h9EqZQH+TFy/ceruUogR8V4115pVWtJM61o3/YUw4j8Of9T4w+YsvYxSBv0+
YTIPegmpy7Eb5l7cIHJ73CsUZ9fHfzFhvnL4xHATmaOYSgXrrVxvRxv4DHn//lB5ip955CcxFD/c
gZluT+7sBOejM83gV14GyLp0hU394yKNP/kxSzCusj+d6hEZflCneun8lxoz2A3hKo8Z7euDzTnu
+LaLezd/Z9zh90RUzb1bc8ELlfutTPj2E8ZGBrgoctNFc5rEbMZfkL69p4i33bUsKqsOLI1h5GFd
EHUYw1X/VLWlyVsNpA0CK53nsh3EIKpVFtFQwFbIYuwlhcCio7o1bctWYMwYq0HZcC+U35rl0M79
/2N2z9ZaSZei6k7GEmDhn1B+gc5lQfWlThgdw9QRULmo7syLRDLVIuWYLHYAkvd9yJOYeunNNNaJ
XOmVZ/yE6ELfS4Auhc4dcFTalkbQS6gEjoMMOrpXZxZdW9rx5lp3Xr9xCCYTxvJVFdOTzFvWpGvO
V2Qn4aOyZimgpyhJoU/99p4yjfRkY1ad7QoTu3qcU43g7f9gCrbUn67iSE7I0nw41mOxIX1dPETP
KQKkYHJ79MccTMoQBmYlbiI6MVXDuqo8mCgdu9WVpT77thijnrHa1oc1D9IcIDdLdIGB9/hx54Z3
Uquv9DJa2aDQ1UExgE4CUyMAI3R3ZwcTb+DvfX8lRT7Xk3pZRPBJ7e1WxQxsNOAm5T+JWPBAsrLF
557IRoQ5s3IEFScBEPJE7NCpeoweHjiQjnYZwb5vrhSuUbQDEXhj3TcFnGi2rTZ8BuxW1EIFVtkS
ug2wbiINhXUBxPM05cn5jIXDkJMV/dG5Lhm69+jTJXuWYcWUT02lwI2qVUGFaIjnkK4UQLsGDFQl
1n6EHKxprdykddXAivIH5FGu4Lx0xvoVoc2Uq7L0hN5NL/ET1+Fq6xaSwUiSrHNsH8XeYQCHla/s
c6mbaP1jBoda2iJbkVMSXMInB5UCKKN0E3RjJj+NSSJuHK2kSk97DkWv0cGGxftrZYbAFKAbtkLG
tPg8ax/f18XvKdBVpN6rpWFWTdGtNmKUbRMZOfW2M3PZY54iIBaYyjD3U3wjsj+KbqZLWphb34bD
7bjWauwtI1GVSJMBBSM5lGG2uxzRfcuQ0Zavk3XdDacc6MHphqFxN0YrgpuNxhuklW+dGoDhc4Ne
rymJsFwN8bpT0Z3ZTZQh7Yeu43rtwN4vZYdrvQHKGMvoMVqlMF0eosKZjpvuKuCqfRFBmjqT1zdE
o2GHjovr33LohjCFgYuUrLa+PLrf0hHK3+fpn24ESiggIP5NhiZR+W8l7b0YMOAdw5saYygpglcV
AZNelg93/xeRt+UgC5wySp6mBFOjQGNb30hAHto0VghoJnGjMcaQ5EJ1wAgd1L+/EksJwrw56Iy4
sDE4p9wjxUay4ZELJKZ8zFPngh3nH2fQSmhbY51obk6z9VYolzw3tzBtlF3uH/Wk11+MDA5ytzrt
0Ns9on9hLaeWMPsNXkEWyckkE65l/mlYCsyalzHmve4Kisyu4BI88uIFoK+Q89mNIHxLe21+yR93
h65eyf41AxpuvTo+EQEfoStuAUkg8FRHARCP04k/54PmZvXafwS1WvHhJ8kKFJbOhhnG/1dB/CNx
3qx1ekWmdS6UEmkLla9Jg7TmHu1n/vwCsQLZ8R7DouKXwowEJLWZNvVbDP2EpEHZOT/ghrAbaFLO
p5rE9sCvzM7FW1Qwga0ZAQNC/cxpOfsLa8vMjYDMAWDTJr5D6K11EfbSG2nv2DfPmWVaGAVLBSB7
U2hYpKnoX8sdlpPvuxoBv+jHo0SnL2KObazPUH23JYOpx5vA54NHCsRBVU9VJYC/8Su4ovTY/3Rg
le6xPNi9DwxC23obl8T1rMn6JyhWf77k164n4InwER4dzefp/6QRW/bKQHAyuc0BZMy/Ib4kt2gy
0tUlPRE2CjwwlGpiY8i82O6U4atC7LfPq0j4zqnLiVZX8C43SmxgebnbtncY24If5FkgA/vIFJV2
beOA6WqGZzrcB70xaEwmj/1tEZ2heVKGD4yXZKULHmE8KKSt4wCZ13khc3YnLcILbsZ58MK3JDhu
1P1j+ZgLcJR9bJtmUm2DM/PvthPf5CSfQL56Ik3nmBPlly07a+g0HfkmKwUJ94vFE5g1MYW8tTxa
l4ZGan85ni8BiuhsVrDtPD+4E357D4tyUtBkieMQf06d1h1aKQVL8dRsPXL+LvOhwnftWry1RpfR
JRKRTdVPOAVZtaB1bLMRhykm/zmNabcflqVCiB2yjvgzJY1wf3RW6jTurY3G/kvzUJ+BDKjhH/IL
xG9Q8mFBoy7Jmuv6UrPr+/NwtFtiLGk8BeMx+51qvvxpleKnDLyNHCMQ738JUmDVJgbvlP+PJzP3
7IMcPp5/Ee+7O1fvL63jj5hWdv7qDiZL2DJHvRUsap5a3Zso4GesIl0Qa2qKsoJyB66uRmWytGEo
Eh6691VyoIbzy3DJ6XXnZj2UQecY6fUbTJHDiUj18MeisKA2OC846ELu36S6DumhilEMkk+tTXAZ
vdRq9+Yf+4+OidXZVuurMBimxg1bYBZEJipwIlDv75L7PPBOBqJ4ClwUe3oy3Y43+T+LTddI3l5C
UuSvyb2+YPox7M7SA9NWm4aXpKmMKM0we8JDDvjCdRXpKjM6969gCUo7ZFQ/lkfk4ZjISzjmdx5W
T/P/us3qH62D2QAOEeDUsNBcZuuJEYjNjJM2UMNxK4Jl+mwqXYlQ2cSnpgZspLoAXPQuVbvPTQrv
qLesRlm/IU77fpEKbEqG2szl4yePOAZL837FGFgymnKPlt8PGvI3P/Hlj6jeyX6oCXJzjQYMttOe
LogV/C+RpKO81cnzqei9SODNe1YVdwyOYsDnF13vsmsSOatq2VT9Hj49cQmhGteDTvWe9Uw1akmc
KHEUJ56iFVhlI5q2pZrhKnY3kZ5ZQZ1boGbHG6AuIsWhnvwFMH7bh8rW8LJwGUxbTc5wXHSRF1j5
LniNvomiVocEueNSv/Klq28bHip4rzlJnDj8cS/tU4G+BbFA1NeXBPfHdzsEbMldF1dGtfOT2r4W
jKHgyS7QETHEknBFUWlQlsU5tONpRgTURRpaeNOjBHDMi1fExvqV0picEYsGXY1/u6rcwI5WBPdk
e8mxBpUXUXJeOoXkKT/T0eq+SvuOtTPYRakcFAVUpxn39o5Fnepp4CieEY1C0+xbGMd70h+7bsz8
pb3T5adoThyfnusKlr9lzOucIkacpY4kZT7ipvTu08NKU4GJK0pHWiNLqMfq80UL8U4C2dahlNML
Y06iIoGUwvk+YwUHw5DOhZoraDpyCS2+qlW09neS2qR4ahtnEiuAPH3SxV9eyoyXoz7eWuhBT+U2
SC6vZtbvR1cfU/3+Astr/LefpiU0SuNyugJx/tSWmxpVyVAcu55rDweodSA2ADaHANqEt25cMXsK
cXZkcBO8Wrevd2ribhJMj9ZyTFmDIWMDHg8RYkmoNO4iDMYr7R/MOB0pdIQvXB66x5nFzPdkwSC0
z168NE1Z28aaKrsh5kJCMHpnqqoMnnBj8NZ0okoSwgAKZdqw6J5w5wLzTUrXjEIKgvdHjN97F0ha
9Vw6jdhILUePSxkDeoGemM8bNITnoYeOPSgRuT8YzCPBq8kSzrOfMaVDV86Uu2Vcwl06v1GvMMoT
019CoLLT4FJbt7BgW5VOahsPXe9uQ0QLDMbQEMTRdsJO6d93ZIDivRY5eHB80Hfp11r9TDzrCZaE
wqdaw2KELYmRBAWMsVJApVb+P4JZDk5Zr2eQCRIBfg1zbJDYdvFkSFIwzUBgUvmWvSM4NpzobYdB
9gxHq3mPokxk0IcKK91+gGi066GxwjRT+7ZjD4LDJgnXGaZwJlKibiSkpS4hemojhy8Me9Jemhix
O2eZTJVzJuynW+EfUSpfmjCjkLJlW0Ouh6I8Aqogsk72IftQoUX4H12amE/ycedjsbFgPJUjmDiY
bwPGg/PbxPLyjlsF9vxF8lAC95tlcJWNWfqBIklD6ElxgZq+OTpD7DVRbzDGJ3Az6RuxWhUm7Mhu
/ZbcMs7UlOq4O5iofF55SUflMEZfspI/oBD/NQcidKSYZJsAQQUKrOns99ossSXelBPj3JRI2RPs
LJRkxmRQlCyaja0k3Ahyqg/8eMf9zGMj4tZQz6ukJLyzxVwoLbWfWDdtTO8VHn9QKmesykgUffYV
AbzJb1/7SgydFbxADM9hDYyR9lzpWuP+e6hLdyguUHQSw9pM1tpEB3SP/YS5moJuQHng2nB2ovtB
UjR/EsGl6cTRLG2QE1eA3+2CWanB+9LM7S2IZ+pqM1DxQhXX3y8hJ+yZ9k2TjerUk7wSdaM1s1JL
AplgdT3zcRB3nKX/cFbV4MObjmDLghw10jp1MLBXGL3IDNYoGVnp9bB5orPPTgYbaDOnDcg+8fyW
0uhIVB+Q38aIAHAiZuq7yjtRAJO84UeuCxJOWFPZbdT52/0ulcsf4sfwdz8rGNHYVmmc8T6o2BJW
055evWWGot0A85jbC9mpbYJ3d1LtqMnq8sQoyICseNUrKOxPbAh3rb/KO2/QASbwkgIkZ8t+05A5
T4uFnPtGmq1lQSd0h82CIHgJiBuSYG/gdYdrKgG6JvSAGeWitAxquKEST751mgqDMxeWvi4/3vSI
eiNAVQjewum+TgfFS3RMLyZB9pXIL7RXd7RwXL3VFPBz76FpH7A/lEQ9WS0ZJ9Z9vvWACWSgkocy
bJ8QXiyneItHvLD0LFzvH/gmSKTyMg9bhSMjBX8DB1NPJZH7BtUtdGMB7wnDkKXv9wbH3huBCzLB
POo1n7uvWgt7xO1rWXaP2v97vGouGZipwCQoAA1kfo9w88EWIs3ztHQB1b1dOcVE+dfkYF0TTHW3
WrA4MrhRYSACMKEvW1W2CH+xfmT/nS2GPmpNil+B+eJyd2i/xmpz9znx1o3BU9nZ7912SRt146oY
5yMlihE6htCph1WQgRv8hVAWVuFhSYI2BKVlx9ll3D3yw+R6jCZ0uOUakolmeCMsHna86VzmtYjL
eCULqEfzr893G2u9YwIFliPwMJCZQ2IC3eoz2x1MjPk/6aAiJCaZ3/t0J97sXwAyFAmzmmLZyIf8
FMxOSRyQNRv/r8G4ZnhCQmubIX5H7ZFzHulgdE9Vp38tz2gHfyDy9Qszj/fy6H9D2YNtNa3QrdZK
4bqBS2tmj3n+4ztQoEe4UEGfkG8N4MI83FNJEkPF4bu1Id2yhjE3yuFjNhWJSBo1XGrSHoTlgrkN
oBYDD+JUxC+LQrUbH5cJaRnpCMUh79fP7Bw113Hg10ymdaY4UNrhPoVFL5A35jMVWbiKMOU9uEEn
fcc16mc7lTcP61jH36NWKybvj3WWcTCvWx80mQ69kBk2KpGN+sUgiRqDymDLhHLSrxs9Mi4HKFJP
hcP33MKZudQmQXCrDKAzPfs+32CyI+4LoE1C69JmJu/DC/zFoQtbAA1L8sbwbfBbKbe4W0kgNd5l
1/rhhXgi/+53s2f58Nes7FhIO4ICU5XfzJcj/5FqORdX0nQZCmUFkSNIDj4BDiXNzVfGVo5ivSCk
Y/6/nxdEpyEq0q4BgX6AtB5giBz++bZKRxM5Mc6M2D+HN3NsG8ZZ5drHU6wSKvqnaxTEXh2d0c5O
r2UmQVp+9yN57KNQOGXQ5u33X50bDNOw33sFBMGpMkvCvqmhRdhS+4DMCPw9kJ4oKzDnl5rpD53z
H4rVHUKNyW/AYR/TXAExBic1IqQNkVO/P2ZgUDGrW/kySj4pSHZUqADe7WgvrOByoCoc/iRLw5Wz
eXY1wB9CubaspXwccK9o1vVkpVxv9gqOcZEWUsKPFhfA2yQUnc0miWwq7ggl4JNvmAUQ1ZjKKG6/
7jgV3y1yKdnQBQzsBBeALMOKPlJLFD3IB64F6eS3gm8Tg+FSJawKNV7mSG+asbbglXhug+C5hFTA
dcMpwfTWQ6MWqjQDmI7HC5/AfC3i5zPWX/tO2rTBYZQkAzhmxMeG1FzIJawQGj54oTCtnR60F5ju
ryQGG5mlohGcnTpuuq8Qh5eB1eK6fce2XNhOioOZJdnji3BMoZPulHRZggfTzua73m+xlWSVsfh5
5OliM8Z8yXfIAqOKYDS9a85JJ5Ryv63Cm3Q3IjowpsOvrEtGU8RorCSWFk7V1QF+908VqK7IyIV5
e0WCkOk9c5cOvblcHltKyqrJdBxPq7ZQlpnHvz3eOxRL7m8ZkDleLmWXatgVq+e6qkktr/b3sDya
QBPrU4rUgt3FoPtM5s2+OzEnp+ZrEAL9q3JGFAndXz05ULP074hlyyle6fmX8xhpaDAA413W4dES
BG6e8ypbGKmACZOwun99qiyx6i17KXjeqtdxM890vq0NXUzEmL8RZ2kqS4FyZQhjnYbCntcYbCQY
H2jG9l+hJozXc9hAsrhAN0IDCyvY/IzCPHItZEk95GLYTMMlrXncMs8zlIQxedG2xkv3Y3a7R8Om
aajEBR85bx37/+9FI7D94+Sd4TbxEcvUBt1vyDneBeJz5LxlAGyp05hBqU6iz+xCeUbIbZ0YGdLk
z4D3fmyTalt3qI2ovgrq364SB41o9S2L33N27IhBu4CQ0Sz5S8JCZgxBCJH8lvwjAYOQmSZgxDxJ
hjAUKQ3v2ns6WckHrmfKXThpvEVWHn9qmmgMNlTAUK5hVvq12DYq140sS6QOzPUgRw46v8ktdYXy
e+KLQm/DzLNt/o9NRTdF4s8A/xbvhnHghmgJF5azdyzA8Yh6a2vw6HFd74HPcZs6As/9rciIwRYv
ti5QA8sBOa6rqJ+nSkYA9MkwldZfhtKu58i1tayurEVTOW2BtjiH8j9pB1ANd4d+WR83ZvzEAJRe
ZIYq2JhLp60dPuzxOsawiMdwiuXriQJCKUEj2mJFJh4/ELaXUOwbibz+L8p+4+8NVLfMqP5EjIXU
+Mdjj1qbUicpVAP2I4GfJwVMEFu1qgIP68LsES3WwRQ+fXbi7QbHY9R2vK4D0RwqLIYcf+9TUV3Q
mQmK1PlOmBJgmtVF8Hv3TKVOmUg3203IoqweAP4fOV8RxL1Uwpnx858lTYXdWHU0WXbxs4T9mHcO
88JAtMuuVxUN6rsskGLdm4iPOa32Zpw8MoP8U3Y+SMowsBOtMlZworNlXT08gTuyLGgwwDMNrLiW
A5O9dtRJLiaSbSoBzxWQFSH1JcF1waL8iwCQq2BUf/ZzyyL2atBttNqnZDROtHPMnSsLiSftVjQv
Q56KA4U+r+6gCyY0wqTziwYb489RVKlvr3k7zNxyywrHj563vH1Cqcls4qmKXOBTJ+41dkfPNU9d
Uw6nCFe/I5Ct10EhKsBDCKQdact7xGiikdrxuEjAR+mmqRJP7jzYVVUiGyqiSzps/DmDcgTrhiV9
sBbLyVMq4tXgw3DDhDhytlblfPJiCdfUwZ0qNRZxBYGGIRdQqv2pnu4hBsgkzFgLCGxi+fZ72E5J
ml5X4J1DaxrO3GO++yUhU63r7x62/9ynHirTjJIIkg3bwcQ1UpvslRKK85dgHXKo2gqGLxu9ih2z
oVuvo6cVgsP2ry+0FnDOgSq50c6IUZQoHPeKQJHCnpAYGx1dqckOEJdsbjDUz7NWWQ3CHUz+MkLJ
UZ5I90S4uEksSIwPoIdkAWdx1dwdRmbjdT2a0XNTwkQWd+kA4AeJLBeNgCJFotXMk9n7nA8/BZqZ
BEOICSAQZGEG3I8iG5qcGiVis+QqEldeVK/fTHg0x2Sq5Hoyf9XxjH5lY6IKi+zYPBz0KiJnd9Aa
VHXsHrCS+PfAYos5P7kWxeQnyGrcBgH3/Dj6YgnlHD3JX0msbvT+Tv6c8QlmuDgvcSrblXm6CapI
+CeiDAh6Kv5AdV5NSa10f+94nEgDziyZXD7nqkndoqy+UGJ5euICeFGgt/y2k5XFmpF+jGMOmrO4
ncLgyehPuQA25dmu16WrIFjr2GxRqW0pIrly6bh5b6LdFH7cqTa3dj/2CATFgLWdFWHBNbMbBo/X
C2Jtj65NCDMD4c+QGLXqBAOeEWkk1WEtGC8fI8Sc2Ug3XKFaBdGtYE3cSiWleYKSxjb8KWpIfJvw
aC897e4rDrEsnSuAn/8D76tk+Yc60fJurjoaVTv8QBHBRgm8cmRSiRs79BfE+zsI7mc+dD1IM68v
xjU/V3qk6LeX/URA0l86IZpisktDNpPbPgKP7Qxpupt+8Vo/BWF+IpxgOndGkI7l+bv4ASHhaRZk
uoJtvocYuL4VFsoEgtpib2WFnnqU2BXkPfeDex7xiZlgjiVo8zC0rTowjubO1y6x2Z/EQGrxrdcF
aB9SUYw/QNi3LQ7Lt3P2xLsQyQvPM/KftBpzniX+uhR93hqTaqiaqFo3VIDQZBg0B0zpQ2CQ3wZp
ZvAHpr00GYV7/Beubqwh6u8IxKdT6KX7Wm15x9zxrminbGN5L0EYXB0G4kRmHViNeEinoTXE2Pvp
9ISFZXkxvGVi57NPzcxuSJiZ1kjOm2kQX6Us8fYcBmR7D9PnwEdttcOZn3UCG3+h2CbU+NjOEx0a
pWqoTov019qjD9cY60FLDSXu4v6OgpxGnGmAj34M4KlE2cqSlA1wb8pUUaasLuJW169dsHO789x1
nWUQXL++2BCOxFAbajIDwsDilu0/rYhOFOzh6dPQjJpk9iq60iGQqwZhlYfMVElW4folhTyrtv1i
QVm6bdPJUc9lQYFgJKuJind+fOaH5lqZECtGXPTE4D3zBDiqvlIkXhTP47uXUarUZEU2qKCGN4pJ
LCwFnYYfs6mX5K53Na7vcGS95WYgmD/I/gAGW+Z93BMS4cFnDYdDrsezIF129rHFL2Osge+YAs5N
W3CvlFchilaCObuaH3kB8Uh2vU1AGkhWTc+majK/I+KPWljK4HSUDmdwS4vyr+dBWZRvtDEFnaFV
FoDglGtX9RMQf4aWIAjL34ka1AVPm6ECPgK7FWUma+/CbW2hRhyfMGHq39bnKy5nA4F5pspOITO8
XzR2bAGH1iG0JzCt1qLg/PLoBQCwFChxLlEbN2UEcgkroS+YnE617ikn+814nEHPVzyVehWh+eGE
/r2VVs8ZbcVaXh2uyk5ouCKBqaFFg+fS4mQAmkO472CVq5kQude0qWoPOVUXJL+u9ehngcRZPl3d
MEUcH4OsMzK3XvjdutEx1NcxRP1IeEKpSuiw1CjvTcGEGsiZ93joTNu1ecEKFoomNQO4iwMtzbhc
fXkOA7rt6RqpVT8FZwhGPI01deodPLWgT1/J8qvC42gXrmeUIkolIH5IXka/PKHKhtdA+0iRQMTN
NHr5NjtT/mY44gamXB7EHQ2xF9seSe2rBM6ZGiyb18Cm1L7w6EwkH7uGr8xiXfnsADJmVjxhWLNt
JyMQB5szlIKW5RuBrslPQOK4e21KSiPEwZXBBGFeCwMj8sp02kmQMSw5UbM3vWJiKLXzWHzYnQzG
PYbYws0XJDCymBbjnyw23MbytdqjJf/RgVgwSMOAX0syWTkPmZPCqdPGMOm83V/OVG0nOYFJlqv5
TNewD0mPXAcra5G86BFtzCLfRoJ37ZfJQLD+wOLM2Z36aE+Zzvd4J7EoZZ9PEItuw/mae5cQL8ES
T97SZS4qHCLJ4yJBBKYINOjeOnD9fscMid5bRRYNRyB4P5XLDKVSq6T1H/BPUlsmeZmWhQSM8zue
LnP30lUgBjTgrmHpMUdMT8NOM4xBx57gvmjxhi9yl/jgzY9SfjoAP2fz7fsJZUD9My8ocJDRk9re
B2wmXcACTqtu25ngpMmAI7AFHC5UbD1KKtOwdFYcUQXaFXJm3nJcdxFX3a2PkBWGtSkg3e/fu/Rz
1BSS6mZhwh2DZ1oACMmtNUdUdhFHiiENVWH/qUseBanRiYWY1AO1KO3bckOXxQWjYYj7Zn7ZGjXc
OIFoiem3meWPqwsrlgz3Wm9Ch6ZmfKhrWO+USAUmC4sg83T/h2Vt1TYWa441K/Zguj/bBApZKREo
G/PBdPdWhzm04qi33oL5jnBIQMW2/UoaW/76IS3m0BUTwG0wGfy7jZvNY+w13joXZXVmF/qd42pr
gWay6ZTFEHTM9tZQnzSR2WtfTSebc4NfMRaW83tQqVBJ0ZkCD8SQ86juE6SBPGB6l/yDjiTQS6gk
NGa9tx5Ra9OmGVeYDyRGnOPtO1TbTGHAHDRcS50k5C3KSD4nUQBE0X9YmJ+nY+IbQdiOpLX1GoGi
zjI9VxerSE2Cr1thm+6o8nT1CQckwHlzTwL63OGQ26ZV8n9WzJrnFP1j83BBoy+6CON9v/2Y7MlC
OH0HYM+7tmVhDJSOrI/7F73uYlPXQ1BhL69036cLY0Ch2sjxGPQvvMAN3rrWkLbNaILcrOCjzZQf
/2bxr2dAkJRlkMdJSmyu0oi0aH0zaF8Zk5nwIWUFCJo9/Z6HvPuk9YEUWCzbF2xZ+NbqoGQVvo2I
WNqbuq43oTWgD1Wo97HnVD0icebhB+DpM7jDuZ80Ra0GjAK+CAWym44fz+1wDRgceKM8lp/mLeWf
U1cIjk0MR5muJSgiMSu2cFRkuyHPFzltdotklGCMZ7hZDZDrm2NNWqXLlhwC0ngReC3zm3SgDg9X
GATO/J++dVLvJwz+g4WipO0Xc5fgWbEyLR0yUvASFrptPRjoHx/TvojHbwx7ygnbLMhx3jJTCMQq
3oV4mipzS2Ygx7DnOVI5OZJ45HNTOGPT8ILKB1ldqjX7P+z3H9M1IVxM/0KyZHIpmFyNrTjYnhDq
Ft1hT2TEe05Wd5YoIh9/HPdWLPwbBRdtG6JkM5EMFCUawmqyTp5JxPEMWruwm52k0lzcDNDw7EGM
/VJIdSOFE+DC0evr8S5zHrX6dLcEANtm9Yrnuv9bBs/gtTuTJg0IIzW5Vccg0TeY4Dc1Lrk9GT3z
nXGQwnwgIu/V1M0MkDO0b8tFyVx0o2cOW9Zvi3hiVL8GMoviEIbdLcixyJ6TJcWhbrqhYsST+QCv
7KrIxmTognuSEh+BjIAE75mnj0GYtXwL+YuNvaWSVVc+2m9xXYvoQ5uTr3eP+m6CbW45AMkeLqvy
0aG7kjLMFs6r7TghygtOVd0umQaP7nYcQheWHO5krElS6+0Sumfie7K5MCkPKHfaupbazvJ7mvxB
Mlr5SQYAiGmh64daJrIjrTGrKlOFcG6AMsl/IoX6XQpP7mFKu9sNV/AGxzOezdkJAo64C1oJloX9
HcRiL8PV4sd9Xt8L6oMeGMK9NouHBBONTeP7DUnlCVgHtsBNbxg+oUbb6lwxYVkCkTeQnWIuemoO
nwviKz6nrA+0zjfa78SZmZhHnpOWfDVGY0/8tK6GJEu2rRSE2txN6B+vrRCVj4+Z4pHGzN1jA2xT
AzEE/5YOGjffijFFgj6BboB6taE5rptP/1s6yY7NaMVmwf8OvnxTpYWMOzGb8YlX0mbJKVoUYRpd
SbhJT2G/TP6geKqfI1/93lTW9SZmd9G8xvltAIf15jVQE5m/Mi2qIFxGH99jANfjaQd7QnqCNiIf
tFdhxKBpHmDT/46QJFuNgpYSGRHCdQXUUS7Gz7hjPuYn7RAiiseu5/atOH11mquUUCKBqXUEf8jH
x3l2xoMUPp9AdYjEbKi9/3PcliLJ1iBiY+Nd9V7mC8ySz1LbpUY8ZAEAnzD1VmEvPza82+vLC4l+
6K3UpU+geror9GquF15Jq3l808dGHJ02CEYqzeR0cmNshpERTTzYhM4uv3ofvM36E9nL9sb2kIMb
XarQI36ZnW0b/zi6PZelC0419k3hxMuN8rmVh19LeKeP/9o4BETcSPjXvxQ/slvF5G6iWipEsuJj
25N5Is9nDYnot6TOgcK07Cse/1/CjjV7KKd4zi1VHS4MAlH04T/IDIqhRc6P4qwfnVFH9njM+bJI
amH+4jsmPZhy6KLop5xEWy8eUdohAykPmJ/lsZh0h9xrB9m8WV4WGtON6s8ndgopLM4oHHfGhnRa
ZApx3fcfYo+e0FN7PEaiI9MkF2Snyz/SYtF0/taxJCCUDN/on97dQ0yED/TxKat9EjSKbpmvinda
tM0okooqVNUFpL/O2BQj6sM/iyDoZZIZHo/1r4viYDHqGhx9QYeqkzq4wXyp+gJVrihgIQogqW+E
Mc+IM06yp0mofTA4NZ5SCcdDkGa/4k2WJDjfQjA0Zclp0BhBmWdWarwpGh7N40oV7GISrOpGrozn
dqKXhnxot3nDSVPinVRJICaq4u7GRsmGOXi7etONxp44uVxHjpgAY5LP77oDO3nV4TMMX11NGMyQ
ZPolUk7V9YlhqoXFRDwEN5F8pWXInOAFPraBAr8Gr/abNjaV2ns/liweAA0ZIJstAiDZ+fqmFFLl
1pdisYDI0jcVMS/N/LOwheLUSqdw6YT8wQ1w4ZIdU/uLXmS62j3VTScHzjHaFohRzlKu4uEb1OLY
wBRu+XL5dEOrkZJUcIHgDesVsNWPNYbAxfma3v+cfqXTM7bYMZLIIuzI3Us4Mbalnd4H/hIr9O4k
WKx5opUssgd362LXAAkRSZvDFJ/iT1kLdEMlGcvSdkdIeytUZU/EBdtYlVxb7lSM4OZh44QG+psV
gjPCanDTk6wFAKlkuPLZS8xD0cjHq75j1UMipVYZZUnDgw6bMRJcSGgKagWbVfphqILsJ4cYQOK4
4Fcdr6mcIqlTwLC7sQEoisvbi3cjYWYmt7lb59gm58WwFqVYLROmC9wbpTLzvQL1vMewL0WGizWA
4xZaWxnN3EM/b4kPvSlPJ4Xvl+teRLsVb1f2A9wMLEM07a0y8UMej5g+qLeFoeCjvaPEr6i710FE
jU1Vyvgsqu35UNGj9PQ4atlP1EDLSpz9Bp25v7g9+cjjC6Omv11AhAVEtvLHSzKWDmGcK5PRB7Dd
QgOOKyg7v3vdc7VTmQ5ZX4YO31z0HPLWe0bfMPt+8+N6q0bLs2YIyXyO0v8lsTZ/t7qMeb8qsSx1
pMRZzu7KhWGAk4WNQ/ggHPQCNG9JH/OTzCC50ShJO3d0y87o98zbsJQVSjoV71MrqAE779wSNNv8
owiE5RSEb5UC2NcGkoqiiQM9V8SksuGunsvSbUAsyE4TgctsWLKHVBhzOiidQicny7dmi7Lpco3l
/2s7cfj2OhjMMrWL/WNfPJJ/WaIHIhgUO2XAa7vs6FkghN3anpVgachsLfARyjGhN9Hd+24HRpqe
iRZDSQ4tpshFDnIiIhFlxjlZmlXNMAhatK6zleU1/C404FH7safvKMTcq3vt7a5P+eSrzMX46cLl
I7xhj/81mRJOueo/RJzdm013W3DOgmyW2q1D8ajp3qnhyWYrbFJNXT9JSFfLHoez7AU/Spm7gx6L
oTYCz0eJWAuUsBKX709Zjw+85D3O8VQl17HCp2xxnCyuuI2T+A7USuhrAYb1HtEkbKXsGwOe986n
iXs8353VBzAukUHFGNuvICd8xoew0f8JBwzkEdE+S6KtmtBnudwcSOEPSNyOeGGn9YluI/jE0JWQ
Prq+6m2uo8lYfUxohoJPfOMaUbZ4DpJXH/hWSUWEtz+QwXwcNtxiICGAG9CULYG3ETj7zZ4BdHqQ
k59snwLYRIEKLgxx2Btjj+5urSZ3Cc7C5o1YLdXIKHrcUKZ9tC2ALM2K4DUC8VmB4ahfJpeHwx4A
f45TUN6V7X5YOBI7XTtT3qgzrGPndcYj653pz0Epi70iop99KZoDut3Sjr/gAEYUNyt2MLP9YeBF
sbd3fZgEPwOgJjnqeXE0Jujc76k06K//2wgt3eOQNiK14YFJNLwxnFqoAVNSEsFsc5vsPEW8tbfu
aGHu/vObTtdEL6RPY8TXkqlGP5rdPa2Nd6L53MCCND68qzKJzT5soia35an8dhFSYRC9l7uaNnRP
evEubEaknzB2IIkDpE58cCJSKoAIuN74Gb/rRn0Pckj9QS+HCIEvjkoF/ybgaml/aOKrqu6RGKLP
wu/xGVXAq7wHKfuQgyfAsNQqJVdQTGj48O6PsrP/xLG5DAFGKqZn1zIyPpef+CiQWWHsEWYX3gZ7
0SX/SvfnkUX8ruOc1m7ea42Rfy48hJHUyi1JcIJNJmhYumKAmweu8b+HjAqDgEojjHMzFRSplyR2
IhhCVsdSUtsOLVdkSvrhpJgfjS7watiJyvI5vh2ZxveGjsITL9QcDGNw5LUtEFD/dW/FO7d/ZqkW
JS7JIwZoZ6bwIo4IztWQacSzLlsN0IF4Y2qWe6zZ612IWe5/trwnjMuqgExq5SH4YlOrRqPtaPzU
B5W7bntYOMpqmoD39pG8Frok5eGhS3MXAb+Hmv7rf4m8dfk90oGKqchZy2J3/EFMeT8adyvuVS58
9laQk25qiQsf++i8imksgBI1ZFDIe80ykGxIj/GVLMSQpGkiB5S7JrOvjBxkTvXNmsRZkOu5pDjc
KnqM6pbpB2nBV+4j1xr7Nyb9jz/qwqVfVtzrf4J6E1MBzbokl0yQ47pu/bFcP2khLU4jPv+UeGht
HllTXP+81650BEYQenx27S850f0y4FQwEpxEzTmokNSUFm3TXFO/eBIaP08JRrldR5JYFCXmXMI1
JhRvHpnL7RKoojK6WxdiSiOnzajDRytPG7Gax4xY/93vPMzpvgtq72XRJai+yfPz5vz1qDLG5ws+
0MMkN1Bv+ZcsDP25u9IRB9cgZJTr48X/BeD6rN+FYDdlmxwpohvYQSmZKgtBUq0Wm5Q8HNbDDR/j
c232KYfLIQ3g49dunL5F3b4RN+pkNkB5w+hF2UVhOBF59Ok4WawFH7zkoZhpao/o5n0zWmklIEEJ
AFqRmZnhR7lsfbqoDjUIqfHCJ76Cji24NMJ2UqxxYEquyIK5CDjKB6q2WX+ixncqNVzhr6ji1F5H
DUk5Cxg5Hzv3/FcJpwjRjXoGMmBYNCrqTgLNY9urbssN/1JYWsrgq1yaGrYz8rP65Hsw1GmBxELA
BNo+tYJAvp0bYLqdwW/Z6PJJDDHNvg+vqfAwAm92FLqyO9Tb02Ll1dz6HX213S6iihOw8Hgq/A5H
EFAsRcg71gVbfqAVKNuVo99b78u9InuCLNEC463YlGw0CaqWmQaSWC3/E0T/JUU+F1SC40Vir6Ti
Xs/cBstFe09tesd+7qnxLhzBQe8vfIFthlVY1OjBXkTAZZanE5FMIcz4W5BuPzb6vx3mMH43c3zM
gRn8pmXd5qhGIWZjcJcSTNRRyK+VETLIJqxCjiSye3o+SQqO360VEkY7DUzUbOdyiSdvw532mO8z
Rw1PYTxtAZfcDhumO7b8PVbtlS8EMDJO8LZbvK+Ypz5HsOM5iJQM4aH6o3M2JWYzM+lt8uJBBiCH
oSxaTboP2wh/C4papVmJP77y6MJfgGiEQjvP2tMqWsuveMClnRJrN9H9WoZ118fumP9XbHhhdXu5
ledziZ245pF53Y4bAH/C5ofhIpzHQp9y0Sq0PtGiX7UpPBQLRPkc72sAT8DqLJHELIMWzsS3tntI
HGk0dvptCl0VQP1I8/AIcJz2adXT8lEPiq77d5Xc/GpZ9SbRFvz+vpZ2ZXwj43slxBrVXqAFdNIH
2zpJOCZl6xom8LW7fqCWh4SUz4spam7Y/ec9ZRccWYZfeZjUVkJk2YCnXnKOHqRDI8bYviVh4Rcn
NGfQ45ztMI81tVkhiNloej6+S7OgrYbw0vDZNDIxRsW4etYl9cLYoYQvA1HoQQc11dDBj2yO4bYv
UVbC4ogFX3ZZ065Z6zliuxDtDTkqMdbvkyEFe5tF9N/diWYkAQHXXf85evFAnC5AQfbKXdIXfUzi
+0eTNNoaq4pYlpT0FTYOG0bLupj1dKEWx8YJHNihr3UJ7gfgqgf5eY2XgJXFw8X6o1jl7tCvY7ml
BBdnC1MqUCKqr3Wm5DhvyPi/4OFtvE1IWRR80VAKaggyGvSlRdqk+DpNvBDq9g9wFETRHq/RYpyD
Xpbc/ZLCykojzAT3mBF/lT+lYAF6rj+gW5ZyR274vSZ/E3wzwG5/K4Dqm7AsO89x8qszLMe93ZDD
7b+VY3oi67/o8QJiVBhkVVFQzCxhOVl1XOQDiliTMwwYmtN3/mfuoPxTFYBGICS8DrdGVjhCBdjN
nkKn4WrYRRVIMFQrs8Iu0O9D/I3lXOpEbkiFVZqFNKHUetuTLw/3ASj00nEIkkVGczS9HGjfxLp2
SGa77jJohSwYQU9/e+rAxO+Br/aRotkRXKsL9Xg6NcqqdKoGFPLU/68WHWkx/Dvo7V0zB1rCMQGB
HzXhhBHg8dqggFHkQrjtWgsGFWyn8l3Qouw1Bj4P0Yi6T4cIbHzVSDTQw5MAnASnoAaqfjF60Mfo
z1xLjkz6d0QsqCe/azNZbeeFDru0S5pmsovsA7cau5QEex8sOVBwACkrLpEtlbJZRxZx84eworJp
ccs/nuJwYOMkjhdKlSKbOSB1Ybku1W6TjWXyQvrJBIDVdQNrPtLh8BKUJc5JWRl3KL4F8Q8Jyqoe
/6HRzyUt8gBqxceMh/H+Rv+OvhTk4m9s5uRKlvk8kVxin8a1+97C7pHuDCSXfq/1QnCZKcYsFeyt
oQDV7Olw2U0K92+QAzSy2rC/+LYzY0DIPhZuLoX5LHu1tvYFdwn4GAN+pdPn6gjSSTpS1PBxbsLu
x02kOMRNlazGrf6VYenCbWLCUCrg1XXd3ROa13eWANKTZAMcHXY9XsPTRxmF16MWO1BEEr9SI/iX
Wk6YaCLhm/HkQLJY97XpmTmRDIEA6L9J/eLp1FLk6BJvK7Cp8fiq7tg5pA9qHODhSEnIezvf/3Uh
c0yy70Wywfkox7qSDDi8L+ncK44HJ8xfXziz/5glGTItnyUq8wAJ+YQvt2kT2mqf+sTqdwNTwGht
ko7WTyuG/89zZv8MC3hyP+zhRJ9UMjJ0YieGPAu6zkeMbmzwPfj9ON+FAxY1JuhELG9lNJd2c4IX
KNveckZRWCIK/OxBIsEsLGnl2HxxBlygML2Q/X5GY2L3uD2wrQu9zmZAMN1K7E1iXGegaD5FpsTv
MoyxW/SxYCo4iq1BpHnYIUi8MwIYDkSbtSSUJ1sACOv0eidINRemZq3mCkLbww0WQOx92u8MZu5l
gdEYN2P1ABYtZ3fex96vCdWM+Y8wfuXiba+doZxe8yFQtgAk9GzR1pEAq0aNmfOFnzPOZttRRoG6
lMNq2VuNQctsHidir0K3jfmOtrsltZCwpdTTgabqu08JNmT/ULe1/KgCpP+1LJIJmDEbL3LyVamW
gs1pEs1pu1J8wZ9p6SeWz1hjurTedfej41djp6gBdbg6oV5j6kk4VZxAxitX890r7JFWIg3IwU7t
y7DBC3UW6B0x9bcDsamKcsmkT40uB2S/vklUrt+dsCObHSAW1h35+/oDLJmSfjwS+8A0c3zH9YUS
tnxcZQe+SAmYpagH6+zPM4O3S5gfgSbcer336MAWjykYjVuFInSlu0fCveJpQkKISGF8YEvEL3pK
yw1QZ/d1PTVV5JVors+7A4vP/6pRnGzgDBE1j5rvBqQWcWqeqcx5gWvq3M03/nDkp7rTElnhAxYN
3rBKJ0rm502lsnkZWQTNYnRLcD5Bkogg7MKYIilzXPfPeC0SgLzYO93+yuoY7+DMiIplL0rsTfsS
bgVB4iP9id6/SSXIjEvu3/tPMrMxFK4Aw4RXoLevFIFpLUUaspzcorpXfhbuSA015ZlbxRFWP6na
86ATUBKCn4yQUik4sTvJCTxsbZbRRum2NIHyIyhI5ZnW0fBkn5NIkvRGYeO7sBvmknPOK1Ujt7GV
do9s0EGujqn4wxFHZNuDbQ4VHW1G+Y9DLxXvU9m09d24E6bPR4f0YBqPCIpkDWqJ4hpg/FGSj2XH
ooHJeeRAtE2Jz48GVm1V6OLDMJxXfoaw9L5JDEt3Z1hA4gyFPTFzBZ/c/sOBm2sDWu2S4qinbqQh
iB/7v0h412svrErooWoaZJlSCRKmtr1vIddD2FBv5YPoRzY4EwCbxbx+tlhP1hOeNoTooSsZfpC1
z/SZ/nHCsMYVhlLxUIqOi1V1celKuanf3e40JnJoO4Q/+zY3uHU1JmCuzbm/fyGLJG7zrbEJ8TM0
BYYYYcoHQDaiiz6uZqARv1cTRQfbvHI0Uox0w8AJ86pEtM9WAOOqRnZTFvwocNzkBw16itzlMxmI
CxSNtWLvqERqDkEb2dZwTSBt5SbJx0Q1xiOYb+5MtoSaln4eeUPbvydKLPs8iO4EsblCvurXpWaC
5rc6Ru+GUWaqADYFLOFzMj69k01UZZy3dlXq6Wy8FtRwkELqyy9OwGemx59oEjlfVIAeMvI8Uha2
AGS4kSaCszwD5MUdUw9xTrKElf88UiANePXx4VsJVSXA0x0ygM4N3Hyx7HkgV5p4EG4vyIhMWIwZ
Ws95rfZkw05+IuAQ1CtkoJEY1fRt4BsQwo2/dFtAuoQSzIFV81JVlBB/uBKYR2YAPu2bS+7+ciRR
8m306tUxMJAYi6PYwhs1evlHZeF8TosvxRaxKcaqNrD1ZbXG3zFhn/ZzGdSHt1HQZbddvzM9wRK2
+D1NNNlgjCcq4aY7qjiNR5wUsBe84dBt1AMgJtgxOcInm0xuwiFuFjoW3thvjHbHHtmdxQmf+c34
mj530RoBfX09cCIMWU208AZyoeEYLqWngVEBwF/FR489m+oH1qSMv5m47ZTUoyTTzlNTOC2+2025
s2jCcFghFHG85V5oRzLTSa/Rq4LQ6Pu+QiBK4JxQ040zAWRVP8xDGd3JriBADHIBuN8HCBOQwWvG
azAvQu7WgnVa1lEQcljBqmLqCS9IqRa98XqUmxEm0JJo1TlP5idZ87oi8T/g4qRSKiROE/cMX25F
ixslivH2kJVSaPlgiWvhgj/lplE+zXrBmmJH8v8Ou75tX3YY8W3vz+NNz9aTLkgTKfgiYjOsgnN7
s12CCPB5AzMwUlr+tLFtgylb9mTuLknJ/gEqfoTpiwNOTE9KU7yvLP5JDUd/BQLf/JMcHj6ptRxI
GWzxTmsQu23yutTJHxtnBIYG/fQaCFLVX3H4m6lDcZv3D7LQRoRBw3ESrUo8JlRXlH1j2UofWFtw
jphudIqmXuqOfOpwZWGIRAfsOh5pj8NxMYvj+x3N0zAI6GEna52gV6Infw6qURq5lC65EIyErdKk
YxcWP+Kd45hkOJ3WDfUEF0u3R7nse3RbpY3keDYEV2UxHdUlPNc+ggJAiXftfTkQ39haC1/uPByN
+fsrPmvwiIc8Q+r5Hz0vRvT6Vn636/B9d35C7Jz592nMt2zTvnO+f8K2/zdYIeBjGN7TC3lmu84X
vOSNLrgn6uzVOpILsVCBz+e3HNZeTzJCGxbwtoVkY9fo1tr5VkI/5ef5lZIIez1nLGG1pZQPy4JM
1eV1cwqW1doOybWRKaLaxOYNpoaSeKRKVkntetN5UpRGTHJ4tMX7H851FHMzmLUYA7rspCfnMulC
QAVcs2BE623hXCRWXq5eBh8DnyAY3b/wsX0oY7yvhW4Do0l/vYcWX5lVSQxP8wyHn7sLNlqtQ5Uk
sMDxLqImcRgs3z52iLwA8H6qKgjd2l2wFG6S2rvSRS4fOsN2AaO3FweyOm8foXE4K7QU2Y6el6Vz
HD2q3uTNToBY1p+uTcLnlP6yo6RF/l82DwJs1BrjIVzWLcgVf+6+SPpCH1p8WdLDOhumeHpcNvD2
nJ3HyOOInExGgJB1deKEKAeIpG+nuv94BTsjG01xwVqth1c0sOgjrBb5W3eF4iVsNXgBuIfbF1yf
Wy8/d9tRI+jB/co9zrYcr6EAeLQsfPrCX2Bl8vvRfdQqJLNoAoJ7coGrnQk1L4uyWW6uwjBFAAHP
kBfOX5s2DH+GA5rCnU5V17n9vR1DWoZ+0IpevRGMeO2mBEqY9XHihUtFiJ1N/0xneatziQGKPOpS
9V9RmR0xvoWVKuoGugJOmrtD6fVy855uwpkQhXTadLFR1gtF4585+f8Rzll7L8xOz3sQwby3D8CR
1wSmRmx5urg+Rfvh8st+mVQ4Iwno8UYO77y+WDlEHmunEqw8eWwR4eeTRRa1bhWVQjRyWNBM8vMu
a+RYvAzhzKGx+ttV5C2VHQvpoYePKBXlW236leJmN6RagRIF0K3PyYm1T7n4aEXUSGDqWFQUNNPD
6rvcO1zEf3vpJfo0HmEkCsJ405Vn9IDnQJqDwmmPoJQ9UW6prFm2ufxN7R4CrwOIDqR5Uyddoq1a
rlhIQdDqg9ivXo2mCdKmWyKNOClLuXv7YDkv0Lf/ASQbXzkt/ZDhCKrb/wcc0GtvtMn+39m+aNvR
XAedRpTUcvkiNYohF6ePW2lkBly61YwJh1SFeSW47aAGihfXmX5sGUa49pOXXcrsoJ/d9S3cCI8L
+cVOBHD2kG0xV0SQ988a4QdJaMkJt7jXQKej5OiQijl654+RAmibQvuP/mQpkk65AwB28ce2PbLQ
zxu7r5hLJ1GztbLK/aqJ18yelDoH0w4CDoPaCg00Eokg3Yo4aHLl2pESSURZdd6Qhn3Xqi0ifonF
QM03j5MT1aN14Ee2yUrb0bY2UZdiMSmS7OZ6E8oov4ktMhzuqVjtIOmdwDsjyw6rwBV4HfWsptWK
OpyVCFIIlFZBheN8djQ+mjOgxGGw1WYZd6SlEnVup3F/LAWF9Z3Fy7LazhnkPwoGJqowm7DSQjCz
we1goB8klzPpJrWT0s4yIfW2Ph0w33Oso+V3nY91rf+kpJYfrqqAfNVpXC+vfy3uUKRfJD9LfPwK
TBCpdSedAJ3WyA0nvtwkGRg4IXPy6XrcELBeGXqS/0CNdIsaoKrgAa7Ucqi0nGPJ1ZSlX5ZUUqcP
vVWS9UDgQny3b5YIARRQPEIj1yJfb1U+yyDhxJcYRgxM/LfeigwPRG5NQMHpxky47Shs5O3djEoO
cZVCMLxkfagNF3ONLigNCiW53V3vZOPlPkgXdFU7h6iuX21vkhKQUOa6KwEFNzLvxKjXxHS5XWAz
iS3aJxf//e8y5eVs2TiuI62CLuvYIPhZvVAFH+vh+Hma7LYjuvh+OGfCuBKaf65oJc3cN0V2Nrax
tcNML8oUQn7eWEAWOG+8He0b/6UYjyATWH8Swdgl6ONuFPu3qxf+fpARynGXxVgVdNtMAq67cTnT
fLTJdLpLVoNIeFSOqf13nafpVEx9Bsm3G3CwX689SoqlV8XvVKW8FaB+zOFyY4XkSWQlGsLWaUcP
1UdlmG+JOJm13lMuoFh9L4cy2wATuMI3fZ+QqZCGUbyVPQqsJu/UsJLiTGXltyvjUNYV628nSK7Z
5ZCjRdw72/02HFcKD7U3YGONlJ/348qfDEXcjOP30b9u/MNJI26JI7Igo8GZqWGeuLNVyVeKAkYM
LS5lI/GelKzBg/AjGl32hzUtrTVmYiIT3l8bgST2OPwLbhU5XreY6zhBVEB01RQ2ZslMjg2/WtFh
PLRlY2n5d19dhAh6Osmy8fNVeBoun2nZfrgZH76BkAuL77q39x5Y1+zNw5Bvu2KT53cKv/btsf0H
uFfvX2CiQc0ghmUBvfH3g5BJf8MDMzIvd+A29wcnmd2Hq9NkrxCVeXtPOHa8VqqKM/ICIEGCqSp+
jf/oJYUzs5IPHFSNO+35iiK+uYyduuH/mxYFY39ZiHkyClej+6l2wRKLMNz4yhxu66RNpH5WRlVt
SYi9K2y332M7PQ7ZT4FHm3Ms/WmSa/9IKb4/WuUZKQiPXGUa0qVBYSme5GKtl2TlnlsL89cYPE6F
T1HMrsGwnMH0AyfoE/6M05cuz4GTjRO2bA3+5mqewhT8sFN/jKyXSEKGMzHIkZh5SlY58R/ozpDS
0VQ2dat642IH+hoMshCzWeqF4bs3TcVNpAJ8lsPcx0yxsZ0cMrVuHtDwsDO/X9uHAPjW4zYnzYfx
UUMTVcMiL+x22dkhAU2ds5w+/qMEq0Ae2d1yS1kFWle9s3Eo/w/agM/qm5iARQYj88LFFaFt+QnS
rbXGXfqUpVwCaFRYR1koHEwEvHMY8V+wtTniqY/sug7AB9jkS0/aJ5SgLqM4LzSDJihg0YfAtTNP
j1YLV1Mp8xIVe70Do/KbKnjNT+o8dLFDwbvKaf4bxEoppqGgBwvQFyhhVexZ1UkYdGuG49h0k7F8
Nf8qGDD67psnXQl+/aSNjfxHkR82RnOZWRZAvzueJRxOey49mkEBTQaCpfK7+ZeeddhKJ4Anvg1s
0YVv8WS5S0wY+veL3f10RbBCg5pDxYfhgOWzQ+76VrRDzTw7h0qvZFrLd8gnMvWNe/P9tuuz4KNw
IVgBDi58wwBh8tCBtRK1m1Vuv+DvZx/hZf0UFZ+VmxSV9vrHPbX+Bx7KHT+aCV9WYv+c7KyOmtTc
Yjt28kuEvwn1LQotHyXDK8bZfj5LuOVI3FOz+p1ec7ZZN+mZTU9V0kUL34Bw7g+l2m6mcY298uCK
/9eshIa1rViEVD2vbx8yMtFGuMrWax0SdqkOdGS8tJygWAW0R+v75rqfCjH8epB3Y3GBqbrr0G5a
MCIO819bXRAm5Z1Sqxka3vsLNRpML8v55zuCw8F1cLt782eXiGbBUL+K3FVOLF1zVeJmlzZKpFMz
wJ2bOz+i7ihXddMuNj3NtbPr3EMtPY4LBUZilY2M7bzJIP5P8VbXFQ2gd4DHooM3/eFNCTH5OkMB
aTnvTpNK1zA5jhwNkW+s0OEWHneHjiQa8+sMsgCNB39eyiULx6TaO6WX7WNdbTQ3OlrO8Mt/ecGI
79bUR9a2aq2sEvPBVtIMSk2sMwf1O172UDBVvEfaadTHbM5tf5o7Y2gEF/Ti2bMYe6xilxPMs8zR
4esDVV1YNo7qGBuYqJGYbU3S9Tvxr2GtWd7tl0pXWgVWr83RK8oFjTd0wK5d8bLjA0XxVYynKw6j
SfgGnw1GdOQDm7cW5o6VXoaUZIyq6uSQ2PTcpnZhA37+dvvMcg1ihvcuDmn9eo7q9lnfoHGgvtHX
bd8TnO+VuONo0w40Cw4tJiPkVLFSg1Orv/R/8Qaso6DbCrfQ5oXD2yz4/EHIJZAO54LAIHhGnWIY
EvNd1HH4rx+x73+GnoQ8Ce3nhNEN/d9Q1tS8G1/JlFRmT8d/BaPVyeN9/MsZq3tuzflIhDTi//ot
MFw8DuqK6YTVn6nNVphObJt9/a+3ULnjYuMB5QyvN25QFX7zPOv0gmbAk60rd48/nGA2lZbpnczG
kOZe4c0ofc5xuACp2YmGO8L8hdqRPhaR9fBwgGWqJgqdKbTUbee7iXkpk5h9QB/WQKF0NVItJ3T3
n8aQRgTP5ve5VUg7xh56kn7nmORuv543jTkmZrAlH7hhQKBrVE6Xpsa60STVKhShkifgAACFV5Tg
+KBUrTE4ltTpQ0bKWV+0gC+XP3bWUIBTE0tH4YRQFbjQcwBE3xibddDzOphg9cy5ln7DBCrXBn/p
FtnP9r7V5O5ws6ubH0iCoripv/RKbNJ5e50XA/FL/GrOcnblLI41vExlT/1QgZq0RVR0UcPePWu3
taAAqWj0WH1lBnq4R1Hfjm768NDErMjwMvp+10i58YfYA6eNo1QqCe8/fXBA7ED39Jqqd53SZQCA
omSBfbMu620IwJbXtz1r0aTBlCRteRX+8e22t8XN77LbCPqXit9PQmrAaDdIAnGxSu5C0NInwcyc
Suds9L8Hqn0oMzrtwBjeljmct1QuiO4DKEHkH0hqAj0PooO5bq96eONbB0yjWM07yEFhdN3ysbFG
TKvw75uXtyx2TSdlh5NJV2LoVMf7fskDn04JJZdfgoIxlNd0E3I9ihFkM2B9cGntc+gljqkQ3IQn
hfk4mjlo7U5WcOJEXrIii3hXchoEpmqVfIJwu/g8Hll8mzuF/1x814EDkpMA7nyy6RGnA9mzWLL9
TOX+4lavEZZddt2aSoP1+N6ABQzDkOsw3rtmWVQfX3eFkHAny/End0wDVPl+CkdGmgBqfnQXZl0V
ppDyf/7fM3/bmjbtZqS58f8fZ6fP7SPwY1ftswQduXDE3ZOqDUp+c86NiZwfa3nuAurZCnLqyJLh
qjWdXwUD+KxKpHIGk8pkjiClicmZ/Tn36ebw0aUa7sVC5Xi0uMqZOBuB+/tz0/6Ctf+DHE1qBN3c
ROE873UTDXX/hFzaRFm5xjELNZn/zCx3HPkXWqo4NdeKVQiYeCWk1MtyXsYHtCgFKPJsvFfPR111
RHqV80gPLdtaBvlNs2TmUmTNH3Z7ahiAhHEcKPaqmaJxdDfY/buMxkS6BS7C0iQOFr3hKnHjjaME
U85TWUCKgMS4cHRsvVQ8QP2oR5WQ4LqM78V3kaiBLMMUR6H2qYQlpHPC3Djhj8ScQ1D6Tmrqa+nC
NK6tn8GexdQBNYDx/8HDgCB00mV3CcK8T7/h5e5BZj9MqWfdmyK+Vwy5RCUIaCmT63nt0zM6ayEd
ARcxB10SQcNGE3SDY+He5NlLxoD5CZUTmlHMGclRciu0yqPtRHLzK4R0ty/6ZO6q7YJob1riubxH
XJ1+Qpi1OSKI8RL2YJfrsAkr+EFmZPzs0BMeQQfg9ptjwmjCc68SANWox/0ge4JJ5x256HGFz/RV
NYVh5qbsKvhPPIz+Y/PGDROq6NW+mD2z8NHQXrGqAnPRkccbVbMNsWqrxOAh9/ViqmIrAOACCfzq
sW/nERux8Di4SyhMAEVKLJ25PneHDzisImr/SOdS8IEoCtoxBZJN2xb32zOHl7vrXBCh94Hlelms
grz/KflxpHuVTcWys/OIXChiOQyTrCKCWStB8JYMbj5NUKr7HGdZJUbkoaf2hNEzSW2wf90YOQLu
bUS1AKuHA9njx+M4rHeXt/X0U06AheCdpuhA/J370uxBWDaOCETFWWojHBrlysUPA3IH1RjDuo4Q
3HR56P01KbFzODFXvLpxuD+l2rTWeD4D+8Pyl3CGaE0OFW4lNvroBdgU/OhLSs88k5MpbuRme/3A
PnycmQjUIA31kl5q98GPi1BSu4BzcgFDNklhW7oztQYNQ3u1KsYXX9dLOuZI23g2dOrLHDLzg2hM
BJFpcrk8XmrJiNN3GFHjfEHkluLh8ntU9rXvLBIWeEumRXa2D3Ag/dthvscB0Q81RzQVXd0h5+zy
zWsJ9ntUYTrHN+ytxhQtkES9chvHxhekY2rP6020FKRGk7NWdjH6W1a0eNpRUk6Jb3ev0oBpe2q7
If9ipKU1tDD9zA0teSC9UDTiRmEeXBl1PXk+oZ1oZcVdi1lcvqL+mYmSAXrd6uoPZatU2xIo+3tP
xvzpw2uT4yaOzvSMbiwXjeisZLU47FKoKfhobNonA/gA281OxlRYc6N/uY3SNW+dwuSJ05fhQE3E
nI+vhB0w9ezI2Qs/1iie45HvZ02O/Dke3ocjD2/EBaLennSsX9VghzMESili9hlkR4996oZiVvRP
Xv5bUbClDMaXkBIoiBOoPCCT6ao3Ob4HAZUNo65uFu9KZ5rioQLqGzFtnGmd2LAWb+9Ib1hnQCzl
yRGEhfDnCnwks/yOLMWdcuOLOTELRPZSg2O7NV0+uGB+1V9HCodSp1J1T34FjBqdtxvH1X1llhYs
3u00kgJcWYT9p87FqlPHn/3x+zyoeVmd2a2D8/n1p+oaC9Iz7RrayH0fzognDFRNVFbiF6EgNq7O
F9YLSizKRESM0EtP0EyHyG+nzD+Ab7Mo7lOsZLMJ7NPiaGKGZSOkPfbNhWQsrf6qsWlmfeGuVoIs
KFyWD36AQwlvyI3swIXCeXLCS5ufR08mQ9tADhv2M65SAAxs22trEqDsLehlOP9v9lcnY4YN5fVQ
RWrZ7IyVWWYB5rAD2LmyR5CbgkIXfu+g10hanEuw6LCHpBTyhADsTPECrvuU4AiFO9rZQobQemiF
M6iob0nxIvgT72q4mvyw6DOidqB+49SuGEORVmV5AqCh3TKPLrYXQxegd96O/zTXZiQe63cTBueP
x6V+inoMzuUkG4myxIhrcaQKo+eiu9pqvewapUpub9rOFts1d49jbP0oSlFHXV+NR6PjIifVDQB9
sUz5pl2T8R2UbPtT5oLQjoqhOXFETXvL/Gjd/OWAY0j7SFY2PnuIqCduXimcOYPOXXFS8fjOi6bs
nNvg3PSuRXg37kTyAouxUUoof9abmQ2we/TkATSBp4she0E2okvsaDl5wHWmQtDDWsZSpP1/O/uK
r2JyNSetE0n+d+ImGAxB+34rbG0whPYYRmFMPcpQtf5SHXjkki3IQtlI6NsROkwLXG+p9hZpIgfY
bEg6JoOKSs6W3xrJOVR3iFaofhb7UXvHrBQlqzIr4GIbKLAb9/G4vz/APY2yfjlkK1CPmNll7i9m
zBf2R6isp9xIzswEdDY46pct0mFaeXmC6WobNj8SwK+iDIHHDg9NFbQzKSpVat3o2m7T7acAodoQ
j853v/vljJ/NBtSEVbOmCZr7BPTkWCGoSbfGMQnFwyf6A67HeGdEhhCihfK4NLDyO146v4+Qie9D
0qCvEpTS4cEie3RfVQIpjbJ8ebl0w7L8oiwyurvayK4MF7wF5kUuVBWCsFe99tLRaxKS1Y06b9DV
sgSKKCvLwzSlu7nVyCefZHQpebkCYzGYIUqqg87VAIJy9NPj3yhbemlzCyPjG+9ZbQTGGcI3lFD7
jSjefxWcfMFmyhsRo1R9eCNDqKf8dKrSg8gqFmuZWZjwoW7UnGItF3LKZD96kdB+u803c/yUtQXL
YhJnGRPB8jb1rnyOaBLh+LxpmUpyn+QwD/fuRM2cRglCxaZrjd20UZlxWlIkSy5KWb5YIN4AyWbW
9R4ZXFz2C0RAe6sFooJTRW4QTYHGiKJ6viK1w4fvsLKEKm8MzDKUDF3L6lrmyB7+tBWCYKLC+LbT
mXdtJGsVewekVo5LJPsF7K7YfVPn1u13+R0fvQLexGG3lj+9VFIPgyEQcYqjYVQwOFWKRUxbmCc8
5zG8q7AFh5dcGaz8vA1SGNaJCBn7XaoFi5aOuPV+B0UBD4MlBKYGSyzCiJgfpmT99g8STAiXafvA
EvMoKYgPvHYNz4SuaewaeQXOaOqT195f9cFbWoybfL/leDklPEaBfrx85Tj6v9ejUUnjddq88hu9
uH9kTY89YNAPhJluwJ2iwCE98nhtBGipWLsh3YJWwjBgBI06938LU5wDIprdZfAhMn8prE1/s07e
sYxDS+Y/3XcmBW9vSokybaNPIVgImqVqhLb1EJyZVWnxVf1cXOCnuFyArfUGwLUCJmWc/e53Yx0f
ugqY2/zJdXsotsgmHtokpFmiftaHniGeE1Jv5Ym3leE2Cn4Ox9I/HI85B5XR7DBa+qYoQ2masAO5
pzROS1kgwwmQaWrKvtNl6lrpqgpcms89qE7qT3oynkngLPWgOkciq4z09lxyZ2ZBogOoxm/WUf1J
JcJZMFMKKcK4zVsMqzMWGHwyHi9DqGR4Kb1Yk+325qJGe3B7DDIb4ucQP8jBvYJs13xYxQ2CuS3I
gLk4U6DH5MqQteddo0KKRl0xkPwfQNPhkJyAM4Vch283H2/RNTLHzqoYjoxePLRQpgVzSzSXpiwZ
0eT2z0GTlWic0l3b51SrY6xBmGweTp+y8BfGzfNt6wtXfw1afZWosBjdQVl2vScpEHnGAbCmVUPC
/yMqoBdaGnOlK551PQ/2tk8EACnCZP194TBluY5cKna7YJgtHDOaPf+enBZyzZXMiX0vfAp1pBxv
wTTPl/M3tXdS2C/2XxoCkaDlrNiuMvjj8SwrDp35aVxQwmAXnV6T7YfSNQhKBHGbz+dSnRavfT8G
bUFx5nMCnRxwxc6JMN5GD2jedjtI/+yp4nNlhnl/wc+xQi3qvdGudhgNuRjjQoT5OgYkos8prM1y
B1RIjfBXk7LD4a8FfYfb0VGLk451emqIWbI3/jlTc5HSJOI1xGxGbqjodoFZBVRxBfQMNRmkyn25
cDk8jBRqVY5lgAg53Wx+5U2H8ayBA1+TjgFVyvu/vUyAr/hdfbwC7DjB7yKqhhjOaVkECh1sDVK5
QMdQgjN5r5sUG1Wztf/cPLlUadS5iy7ZeuUhn7fQh/RPXDJ1sEpYqrDgyJ5zY/ueQ6vvShpNd1hZ
+7U9z1Gpn3Zi0Dkl8jHsRT8UwLZOGXoIYnEZj5GY630qFoqbfuEnfYpd1PyNz6lV0hOf5PqekxM1
FsZs0+vUOGqOoD+NDUCkEzl2ufvVgjxKGI+SMRTOeYD3RKbYWArI3MAcZ+2nCzkCruTkDFBjJmWA
nbFmKAg5leiMctx+KmY7oEN2vsFR/QYaqAsXsjX9jshsq4UUIFNpz1dWYMY9U9UEgPYBGLlITDOo
gnwxjKzMDLvcGqDvJ/Ps+jyi2ACKB9basq5bOhZ+K1MxmTrF4rba7VbCSaz1P+YdDpylgL0Ay8Fq
YJG2HuS8waagt9CyslP2/Tlx1k1QzzFUEM/j9ySZjskKMBlwsmKRnsf3vo7U9eI0oGaUu1hhGXEc
QRgF+Osn28NJfj5osBrU3JSzCB4VollwJVtYUgJihDYLgbUH8IzDglCuxLkOdG3BXvTJ/1am4mri
ayTOhHcZ1/vfAoGv1kmMjlQu7nbdzFn4b0BQQkWvJZeAiQx3s5aWTXMklYUWoIDWG0LXEY7cFNOj
wHzEUfBRuPFESnJjCmjVy6S5kkVLA2BAQJ4ftue4CenxfmEcqs38ce+RAJ3p8AdpxnsofudHCiyE
RLDhm4fSjhKCajDHCIUapgMZur5018xq4DZFFnChoXMLage2OpNH7LBJejVA/tB69abB+r8aazBi
1AjjMzOLhX5odkVXfhroUPoP3t84dikmAQ+Vl+b5nrhO6dY2iolK94JO/eY0CaL6eCXvXr4cGg4b
0rgt+uy5irxlmLWKaRI50FAkiTRflATxWEZOmcQltsD/xmPcObK2XA3Dr8raujq8LdZmGQba59jS
EG3L+aCxbZ8oD+nvStDZ5qYe36/Y3q8asl0/DZHGtWaY1T7aAB79CEZ9ao7f/8a2JU0Nhw18GTwE
sucf6RhhyXT3dWvFeAeuilc6z+rfonazhuRIMS3z59/DOSXsl3KtOlG06H8/GRaxe6CwQDJIwTIR
b/GZa4/1bY65y5CGvFuECBSNK1+mxRL2xH9O3BtwExM1iAtKYValmx8VezgQ8vZrPzfJkJ1Ufxmg
jihyTkGREOXXuBKlZ8ob7KY3ScDhwXkJE68pV147BArTDnWvkxZoXUyU0QNTSwFlYQA3v/UGomsG
BBoEPuNPhVqWd28P0MTW8QgXuV7p/jRRlTfZjK67YPQOL4NWdmMn3SxG2l6mJa7f3g8AiSj8vXQT
TaJgrSJlbtmzi0ZPqNHLLbEZcAtFoZxjr7sd1QDtTG1y0S9gy33Ycu50NuOy5Cfcuia9e3yjRAj4
t89heg/2CC8SmKC3FWsk4EX2VpYlcHUjXe0SpN5LrBkWNu3GRsy7vwX0n4t9elDCGK21yg+CFLj+
H4TWvlNJpRfeprMXtnYljr4fArtN7rxLBvQATsKOo3hEqAJ1iFxH7rss2d8zkyJL7RdV0Sl11WW1
owhkcFtu42fAp8FiTBWMfXrAWsMIS5m3Vtkp9lSd8iNynx3foeiuMlmmLzUYaKCi7SrF4JP5vct1
6VScgZTeazoBmyp0fwAkTbRaXf9cP5dsjUgkzwyMGWRh47IC3Q4rWi7Wrr0Vbx+58uvZVW0QuCxq
mNvlXJVd4uffG7TDDhDRqeIJythBR0ZEMr010q5lYmv8iAPuKvPDJLaN/6AhBnsg04YKLe9+jX3s
52fuFVb2b2LEF8V4X+YV8MVrFpsXUgDgnlmO7D71bsZWN+i/soSdi4fcEGJuVGX6XeqJuDAFzwdc
fBqaJnS3aXLmjN29wjDW/VasUsdpxxwSVtVj8XW74lpVzZV8PLD3HEBD7dIbwBvkaN6LY7WNaaJP
R4TVMxrZ7B/Oimr4w9z/W6ET42XuiP9cU3HLXuIb1/enMXJIpvXEDG79xq4fdhGrdr9vkeR2kB5v
9nnHZlTsHga+SMa3IrZXD/ZKqw2MlNSOPI9DwxvjUjDKEoI38kE0q+Mt1j/keSd2q4Y/fEKJZOEo
JbaYTdPW7lmdtO/WkrdsJMxkmFw4aKE4VqNblslAITmmVevqEx3OkjQnEWev198ugX2W+knzZrzw
NEHUJIelyfjLJpmVo1v/IYcmwM79jOX9sQhmWO44HHg0PlhRJYdXL7Kkp8VucAbmloQlmoIBeYgo
9/76m+hONIlam54urKDpD/8AqeaeFoE1U4uR9ZWkPQrH9n90Tn/UMaPlwaeiWYJykcsolwtbF2VP
dK/a8gMlqA+UImMkDZKcY08k7gu52zXbBsml28QrPIy8dmomfXH604ZxfzfQsMoMmkVAVbNjCiLi
xIacKa5Dr8pV/S/xrof+qOvWLcJ7NObYkrMPc2UaI3pceo32K/Mz3VfeZI0e/D0tXBizCg3opYag
ch3cXPnmKfXtUv0wjl888HqTSAYlby4Y9e7VZCTR+uO+hFF3NOCPyo373dmYpxPUE5S0iDZyXN2Y
8+qKRv4Q5s+gFgAaSWbG1wg5idGqZDMs8YWweb6IefSOMCs3JcGlbyRDz4JRIuZ/Wh1KFAounIoW
ZNkmpWSwUtUdvM44cBk/tZOK9y+uWGMQT18FF3LErQwArz6B5z7CBF02GOkmdqvzB8CbeIUfsdhX
hzcUR1hf4J7Qy1Z/NNDytk2dsYMOp4+Rneh1HAADEDrvMWSNvFr7ngD/LoJYAM1agdPeovNr0sqK
kD6ewuJSWxmoBeGigB2OBnW6R8odfN4FJjW4oMNyw8oDsPfFBn91SkRbarZdE1EKqpwcsJU8X90N
uXKpiovAx3hdOiUYFrpAOsdd47QEwril0WEx2F3Y7KlBAbrwlt2su0Crtp/bif9HOcV03BDYDyrF
H2VKOnG0mwcT24HjeltouLAC0DNPFAMKbRP3SgMoswTT/2FsMaB3EuohpZGCoJtOC+Uw+1dv0JLV
jWgzqOWAyx4xiDX4FxOrwk5UUlg/fs5rHnecXFidbDrZ/hq3HvvxFYNv1ybkFQZ76vpWAmvLvAOY
6NuOI61u0Zb4G1HxHomaoyO/7XM1mJFbPyselKJXfXi999CNnGkzFXlmwiuDwUlicrXPWMzIHuN9
zTnInwyAhgyiezFJewTMR3Sz2zfNyHfSsYxpLi2fJI+W+1M1rkvud9beqfZUtMHB30ZtkjC5h2vA
ZbrSM1RMM1Nxb55bB8ns99O+iIF0ByBuHxwB0Q3t90K3NGyZka36/deGW+k6gSh89N+SF1Q/ZmUq
dl+mLknBgUy2lfG2aIBMcAqU7Mn6YCuXA35EowTq9migGGmrVJ/uEW4eIcP63CGZnvQ9gv6F3Vmm
PNjX6VuWX1VTmmTwHH9GPXcR/YNJjYnhrXqVVhvLnqc6MCDuBTnrzOGfCXBSh4+uMtr1ZZPQnGtM
AgQcfSNEeuLRIHkd4dwaMpBKV66EFpWkht+vMWYrxsuuM/Spj4xblkiJ30IpS1roR4IMHC/FaqQ/
2A2cSUAM7KEmYt5Oycy87vHnHXOUWm1JUp2Mz/glDfhSi7xcg8sBZVGuWTXkMCX1DQiCFywMntEb
6UtNfOgfJ2oWUqfFH8nxdozjVp8TOdr1fRKvSwCcloM43zxBlnl2lqLzTgKMoGC5Q7166xlRD2GG
wOk47k/5yMwjnDQLTJTg/T8kn5J3pioWHa81lgbv0dplZ932n7oCX7yF494xmTqqeTKdIR7acSVE
zhWOdo3dvoy+eQoxVJKPDy8Rm2Kf527m+GN+0kSeJ/jlD7jHERk9268nfilIK1GIcoqKl9MfRL7h
HNzYzOAcPpjLwtLCZ8nqwnNWMeEXjhiubF1/IPEM+OAzqTPOk/ZC9ihQxcA/I5Zo2eXaZjignhsF
0EpWyGgdFnH+CpnBOPacLm+EYhA4DJwwgtuOdqgSv5HHwzl+Rg1v01M6BuQBxbcTJQKY6fGmJK8V
s2BL6ktL/Hhsun/rlbeO4hmKmmECIpa074XQxNO29IA5hG82HfZcWaIEt4axWFohZ5iGHC0B3baf
5n61ZhypLAVNvrx+lqcWiYbg6IWEmljrkXEMif5ZOfnAgUtRT3WWcktJrotIqquVl+lgEJrZFFCi
cJXAvmimj774c5ifUxNFfcj4iZ+JKzrIELkVgEff8VgTlm/2XxwCu/II56bqMGY2okQTeCGdeqHQ
c6Zw+jSQT1AiOxfw9r/4eEP/U1VuhjCPQoa4esYDbYe98OOZvEqffJq6WstY0h317LT/+ybAwhfZ
5NuOE3F8KEdyrLD8vyk0/MalmuBDgbTUpzEAm9K2gi1C7YFHnYyFXGATQW5rg2wZY1PqxrkWcQaO
BrSnWZy1v31iNiiIKc1UCkzhiCLaOQsTTvBbfn1zx8yVI+/Pdosis6jHh5hbWT5AOq78VvFFD6lD
m39S+xIOasGImLf/hA6cI+de03txeS3HT2nIZGtayuIvU+ytl0on8pqr8MnRYSbEmnHqHcfTkaJq
n0S5wNAz2sYs+RIckyOvuk6CYCOK/ZvZpDW8JEfWYr4mLZlcUPjsRYowqpCMt/X5p3AqvoqGr8Wz
fEWtLTbwCcgFRhrY1b4vpBwBqOPnWmij5hO6w1hA3OGwxEQnr6Dd+IJE1K84eiyMK5AAAFPfJ1Yj
YZL2Gl6gC4wgbB+PlP4DJGl6mMJsLowGCifXHmTpLRZvGIyessVZg9rbW/ETk9HFwIQoV1Wq6moe
MS8e8TKwEWI50e3fz2g3rNOhfDzsPoLvfqCurRWh6yYL2gTegyJq7ABrfwgkmi7WppneDr7Lcd/W
IGZxKp/zTo1KPRqwBJt8/vtZO2hzVwHcuJG8MJ5atob3y5BrsrHPzya9rRU0DnWR5+IYc6RFd2qx
Sr8vQDo/6QLaxywx60vlGT5PzTgWHAlhUadrV8Usp+xcFNecra+s3NmMlDYRmByzhqPFGJZ8vwyw
p+nYYMevSPJwPQzlK5+gV4vy3ot6GGhhbiquiuNzCoCgMVIjus9HMCcnWodAEYf+zVphJBMbEn4s
AB+XrjZ4Vvqm8ffF/w05wV2/DZr1jpVY6mMOx9nP5Ib1jmVhvwIW2yKw//lr/cXExUjYQJVRk1S5
ZGJE0bkv8690GFmuhkPtw1kSp3Ltgi3Jbxn/PVnyeLKYNcFCoJvyoq6f7KXXtxr3CdANoxaUJBM+
5DgbIFfO1uiQEcXCTHyzqZQWDtNmkowkpdSVmhBCWolhwFtquTL38hlmn+3ZLxn9Bczte1L69YZZ
EYC68x748OypXEn/q+yIkrkL8CjJ7qEKRg1aZuz1RNaPnXNjmCpMkYoLbGltPHrvshNaO0yI21s1
aUoL9dtv2y0/+SJHf5JW6zPt6irBzVo1L4c52WGXhouzSeS0MZtsTGbFdY2565g0XiZfVdwKi2Jj
I6J5HbRurabgB65i2QVGUYQpS2JwvZEz8iuOyxwd2aPNuIF7bnwTLhtJmUcVW9floTXXtVbw4Es+
0AVldGmyX/W7gSmsXigPFHsNShFcxIjxHJPMBsfILTRyvnVVVLbyK9KA0QdzrVmFpc6YOPpCc/Iu
8t+xxxs3qf89biayGMq9viFa2+qGKkp7gL9Dt61+EjHZJ2f2YsvcNmqMX016J+FT/I5Xbbln9EdW
03ASZTWJBdgiqffYvIQvpZwCsX9hj/vHRpjUUDi+pBtp1iJdBCNUdLpTGJJlWcrV8rg4rQ2j22fU
TuxWiGbeSwh/p8mNOaFsOUm577QjxiKjXS8zZ8392j6O7hIE2kJUDNjO6ewQ8JrmgCKIANaqonrp
ew10FXT2YnkERzyXq1EGV12oeZCrAXtyHh/feta+Rlvt7aQ1RL8PYVVUUwO4f7DLZyo11KDF9iar
8dsLhchrAAu8PYzEKuUdOoSopIfriFnZOMrUioCCzgPXcFg8VILD3JkLQZXJ5nBwIKWPpcZ4iqMr
XVOAmIreLWsYOjDzaS+z/q2zvY5MpTBUMwzG5LzlZgLamtUShMFWcMOcsTKSzh0jysRjSwCMNXig
faQgnvhG8cbaKKkSY3+j1YdNHgE83iqbew2KmDWTOIg6GmYxFhoXS1JyZ8TbwiAyBPUsvB+m+yAh
u6G0guSUV+mqbJL7sx1MI7KFA0G3WOUrDHBRbZz6rPEHsVO01vgPCdoiPGboIPN/x1ub0x12sUY0
s6gdat8/5oXCYeOokr8y7oQkvjY1R0dDM//LD4q0pgLOWmIbMx4cKk73LzJZ+mAHdw01r2oJffzj
3XQbP0yq2Ya8TBci7WoTrPB+fcKlJEPlwrbL+NIB37xG5BVvvZWgrOgVuYQb4o16VnyJVTAvVyD9
vDy2Z1kHY20SdGWeGGi5xcpiouoDqxclnK3WtfVM1YMHjGzsolsfz4EV54YrDtcoHfZzayQEErtX
PxdIO/nHZlN8UmsloRi5Xd7RTVltSf3Jg2leJvltbCNPtX+DN5hnOslyHonrBTKOQaDRpTZxlHOd
dkN9hLeHDP3eekCf9cKup5qwANwDzsvWyiqAqXEwjmuMN2u4kgRlkFfZX4rXwkRR83RWQf2x28cA
cBLLEWmm51VQyA2YgVG6OLx6Aui4WSmxL90MJ7enwUk1518/DxMjXfNM8IpoF5pW+TsRJTdiHLL0
VHADQkC0qGeAVYW9yY4rcj14sA7JQ6GaQwRgP0Bnq7hQ7YOWj1at3tY6TyZw7esQ8ZHl3rLZf0tM
0bIiqGMaZE5z97qn6uoJsvnjzHeAtlFOqLM0Nt0TeFXHHjn0Yy/Rjd2Rpqiay4xrupWEbmbTZ0bA
XddxgiKn8DHCY0nhO7tMngYanp6vHpg257j+CJjQjT81zRvCcvOfF3SAEgmn65YPM64MTqsAozzI
6DRDVsm3ecpMt2wDAIPZ/FcnuIP+6b/xcNS36x2hMlcf5Ss5LC4OD8RnpA1Kq88ntifWk0ZgzxF1
yRbWM1Kyt3cQAHN/gxDcEUw1gDV0RdlSrm7sAB23B0a74HgSKI47A/XPCEbxm8AwOZ1apCTdoQZT
dPBuT1lyeXX9YqsPwXqHmOPE5Es8uYbwCZeIyEe6qo7TcGaCUAQQlN1Jbqn6cdXLY4K4GoRbdzg+
jRIbs7w33wARtffD1lg7DMlwC3qadX/TOTU2jZDOSn4RnZ4IGhLEAFvFvVdFv5xVixG/mO/r5/0H
fwBRl+I6mCGH3PNsf82DkN+S9u9N9IzEOQGmx/NBvnB1Ja4veLCobwnZPyoDxH4P6KZRHh/IaMfc
U0ZCOnWkaHc67RdnLoABkKcmCCd0k8gb287Gxc3bTsAO/7uwTRnc94vsrPEjj9yTI9Hc7OfjOWcX
nV8qwXKRB0VbyOxZD2VptB2nh0gZoNF8g1ZkaR/9cyNWhZvcy52MhK2tioIqmjpGPFVW5sLZlcTL
jOHRYE8VgIwpYze10GWrIaPY1uLXM7Gek2STEt/BNFAA6dj7X5+26yhC2Pl03SZ95SL9K6zP55va
igjSiMCHO1G5hm6pbEo2hqaE9qcQyWOb2gqlVbS+qj75/P0AK8465h+HARM19l5PvfWMA/X2chlO
46lFiTswwmM7WxBJxvLESAN5O+VJUUsnsZbq61udGgsn9w7XkYtKf2648QuTa7TvxKxgz2J/AiHZ
SNmJapgqBEDowvSov2kW1JX+I3J+WBaDe50aw5ya5wvzOjfVoO0KS6MvbEhPO+/tzjRGnsJNFGct
I7Ah47SRXjBOLrw7qYj6NYbqNoStxDifCic1MJI+CGk4+ThjACN8zMQ4wkfMRoZAQkMbQxAQ35tH
xUCGUAjdbTsx7vF7BewzDhpAcEm5EWB50fRPwHawr4+3h3r/xQqKUKN+ykrmd/e2Z0KDzhIVE8iV
coVqnHgdbYIuY4tuvL8u9+Ye7dzNn+mNxgX8ohL6iyAn4bkPb0QdZ/6Ij6b+c2bZG0pfkr/VGwmj
/VD8qOyBh1u6iEiJMuczD8K7KsZNuVcbceUxvGEbnl57bpLcFkD2mlDHDk0282H/Hdu8QcU4CXA3
aQdeB21NWirb5iPI0bFBuSljvIXhiUMyglxMDh8G3wzYHiP2ZQHAkX/05z2LOqDebHXWd+cJoHrb
5kA2URSnTXm/iMRePSo2FKF+kL82SK0y4v8k1nmdscIOtqW2Hs+lwlpH+r4QT/5I08LfH50v0kyN
GWi9RkoQM3oFauOtFLsYtS3NqQiMRsdbg/d0oUg+jiNlw5hwhjRXk4eu/PeKLepLEzANnc6iyPnO
gwxRn/ZTiuuAqVog92lVzjVNzO/QWyIM7I1w2DnxqrxHslTon4klRubr+zTfuhJGxyaA7BxMzhq5
cdkbcFSbNePodwLo2pIfk76V6KngdGtOp9v/ceqhbNVXKpBV+WOhZWqd2yItbyQxiPYG8l8Ca/xu
BMNxzMkm/iCc4Ihtqza7vPp6fvqdB/LZPV/GWPNlRzpv1NWUkC0VHZ5G8hugYvjk51PXmm/hW2z9
PUBxxfG6zAw0SD6n8vNnxSAShcj+66KWIKKac8XQeR62mVpbtcXp3jbW2UT+OX2NceuMr7cEjd11
fa5qjU7FBvXgxwPplYxIGm2l4vgGDvOYpTcIzL+CuMVmoXT/2VT8U95lN9WTSTmZifoa4FcwaJDn
QcjjA1az6MZRu01t7QJ5/SSe4cfnZAeHiZa6NoLx+er4Gx1RzZL65xX9sKGcjBxgLWsgJazTGkne
TcbvTImIIn8b8ZNB96UOGeb/PYXmZ7DjeMjgerOdzB/pSHBa8xWTXbDC2NmfDuRt+CCIk9aKhPRA
qEBShYXrfKzjG3Y37z95z/6fqLXCSbmZ1WGSk6hoWd9NtEjLuroYSyQriwTqDHLof5JmJvqZ6trN
toALPp9VjtUThI5+cP4WFOhHHN8g/Z/gZtDQXYcowUpsGOuIvdqmM6EmrRrWhIOtl40xPF2ZHHeI
c2+/Y3kHD6zncSAsyAgBwaxWLiDP9gSTSRu0oxMnRxxPxOWM+UpbANZtvVOg6ds+x+AeNnlps4KT
5MAvBxx8pKjo22hv8AYcNd2aZ7xI5fPQPE5/CMV+dXzZlJz/PlWlLABujccrbHgcNOHTyPAIrHH6
Y3m6s5Cbm5AHRLQNXtBagbg0b+b/rOBdwgF4+fjUfl0ZR58VKMGaj5cD2/DtIEP1Lcc+y10EFVkU
9AuL+iiMGiSZC24ejzbIfNwjhIMaORY7fc0OP3zmLsrOAz/4zAvx6XZ6SMaQYU4dpeYelatqB2CV
+8JE//Tr6ebZ9GTIWxBCBUwPnlENBC77pxSn/oi0vkmDueMw06sHPZdMPj4IEPfDdngRk6Houkwc
tielffc8kAenHHMGJaxfCVKSdrfotrDa6BWSKVE6H98jACbkQKlzSSxW8O5EeJ7HD94eThu1kBOh
r4vWVcjb+78cq+maMf/oEeEvBkUXhKDnSpxd8MsHz7y+62zOAhfxoHyDaCE0FD4ZReqIcAg9nVnz
PcPTnO8Wtlhx7dVS3JZ6VeGHnHUUaXB581WxF3AC1n1p56+3bRIQVui2iXFBmHbN7tfQnYa0We1J
8su7567ANqdCD62g5LZu218z4kTFjTvKZH6usU4CxH1OZtYxKD5KCNohWaDicnW3AjQy+VksYWC3
EIX54wexNb/VpdiHWGnaN704SOE8LmUROVCyk2EyMKNqc1n3i4W/SIEYZQ/4bHeEFNJ8nXkxzU+S
N1uwgkXaAk5DlGleNlRdmoJzxYQ4upMghdI/mXp7ZwwDxfMc9+LPDkUgQ8ULpUkgWc23QMEN9ZLW
q9LeTMH42/qU6PmeI5Y49Y9o+i9r7WEtVu7qR0r1du3xt2usAy2UrPQUwjB97hZiSbLMIo29FjiX
KOazSwj7vAtr2DswqikDXW3Xo+S5zoBGd1F5z+sxIMpSKIlJ19NX/na20aXmTr6efrdmLWbrz5wK
xHk+V1/RDDPjMifPEft0SowhwQR13l1fYA1kZys9r6TKCcxo6bv3KcbN9JtgIV0I+pZo7fO/C7Ms
pXkvyvDQncRhZgLXkewbn0CE+ofkwmcBOeI3Lmp8aWrad3s9tdWtqeAFl/uI4pRXTY7nIQqYDUef
wiqrCIJ+DlMdLGB5vnueHq0c0QrDT+uzkqT6c927FhcJ/xx/s2C5Y1NhF0fJ2cYJ0WzjqNF+itup
1OWQl1JlGHK5FsAscju4BLcjKKtZcPSj1ew8kdL1t68o4hqnBPgn8fJ84V0y9Tyj5Drsj5VvcyAd
ZiOZiwFaGTqixagNC8U9QUh78Wc/58DwGkBQdO4kwOkaDhQtXCFqnmK3tBnr86sJQf0b/wfQudaM
A7QFr8a0z4XWKFTySbaogp2ENqZ1dOc0cptEm8QaqoHXRNux642ksYxJB0/vOddLjMEXeBKkN0dv
oLByvMCYfkHO+JlWw+trZVIR8E250XUir/Y8yOuP7R+PvnbCM2Cpp3GizmGGWyBNZEhLDjBSnspu
f/2lrHvYcgxZCAlZgxolahZLXpJjz25ArFc3aPBmtsHvSDsBB7EHvOsLPv3cs35hdgNsgYg9C7y3
WAEJaFUlz/Gr79kEd3sgmy7VtoXk9Lq1dpfJH9iG8MH0iLybmp9khy5iTSmNEERZJdKdizicQfUZ
NIDR4jAQ5QbkW2akiEWQ07Ri2nShKIfQqBwOFgOFmH9Es1yh6qfJVCYSdgam0mFdrfmLf0dPg+yq
UojEsIf97QsbmmtBmrnZwXvF/3jXS+n+Ma7GnBAyJB3kQ3+kPfvcpz3VHd0Q7axbEqBENaP3cfZA
cz6a/80JsNOw+pUsonhQSSrp2U70BrdhfRN6vxwoMAH7UVh2xgt7r7ro/0PM5wTVCA57VjZxA6X3
PAUP0D5HqFMMhCktVeOCj8hZYuybiVgMpn2SMNhM08TwJwWT+eAPAXPOa6KZdoD8Krn979bcdCoJ
dKe5gejtG34Q/tACxzPuH2k9j4FrhmF2K1wqHC5eblDd3mNPO7TVD8DIGs2KX4arhb0KYi4ZNl8b
mj4gNhOlsFHSsWkn0qNsL1e8NN7mr7urYr3C9QujwxigWbA6zTfenvE8Z0t/s1fp8vx2ACthtXqE
m4srhGVhBpdEkMHDMWoZgaZMPvuSC8vcK9esgnUeD9exfF3dMj1KBs3LNDZaWypeKuMmaIEFAH2M
F3V5B7FxPXN1as88AA6sTJYjTsR6Fv+wL4Bq+iYDqG8ffe5sYLz1sJHNUlo+O3bZqQiwGQNSuJrJ
111Uw6kIN7/I3wSgGLlFIED4BE9DnVwLxM+PH9zbrb220oOuiNYQ5WoEPYA7PbliiNA/qT1Ew1lU
wOO0o1Jt37909QjNmdcKazxODGBBL6t9Asc99XbKVzviMOMYYIKKhBp5uPWOd+k9kTGqaJ5gp6lv
LOPaj0K1Ylr5EOkOGQU8fNy4ZQmCI/QyReCGGwKg7LeF7EeIwIQ23MFJsX5g+dIU+gR1DH1hE1QH
4GbaketG4d5CY5DAI6xay2hXywsc1FuqOZMVo9nhxh5D+cAp0kO1YEnpJKkbZ7E8+Z0XrTHNmzuP
NC+RTh37QCHYSkIcNLkMMuGXvzHyiiUZl37KD9dDdTJTgFOaPAW2ZQyRW1lPNkxOvLekSFQG4Mar
NSnPssdNMNyklcj2tWA3gWnkWOgWyQeK9H8ix+6YHvFKG4qHWrfXAjX1eQ73VY+sqyXocpyQy5Ls
SmrnssQvjr14v6hktkQNN2CWkOzE53CEd9ypGMEjXB4XOr96kLeneSdUYqFO37XdzxQ73mHNdiSZ
GewHRhgFlHcjaymbAuuXKdicv4oxtjUjzFhwyt4t2enMh8FBizMukbKfbeR+NIjHXXSUyj/pemeq
e+PxJo/V2pOYOvEBAOaFURnGhj7SpLpSSAQ7VH27+96v/B2ceh3xWH+tm1R+bcG+hT7OR2saAfAm
Q2RKtX2i0bTa5J4KDE7elIlIjssImY4B7mK96X7YIvphpvT/2Ec6SSWOVTM9ul2OuIFCkEWgsdsd
cRvimIBwa0cyO6UlrmiOqsFNmFCC68O7siWQi4Bjg8qQRqS/jIS1rk28ot02xtVL6rcqHWDBrjUm
VyUocau4mqizC+dtl1KzRRJ8AEpLO/hgqeuuIVhhV218ijfcbiSFUDvtRddCd+D8mo0BuzOf79fl
vzJ2Prmxf5tdstadv+IFmOEp5Y5GiW8hKy+tQsKnU4upx/NkIODiEY5arG4wgrDrVfMol/yaQLCL
OtHq3pjAzAO1HlsvuzFiivIP2ipuwPWFq15BGcqf8IHR5/VhoGwpXamYm9AyaPoYAe5pfON5WHyp
c2Y1jJC8rxCgCwv+80hnMjsrl04aVfhvmtNHhAWXtzlZ1kW/q8+irjZxA9JrGx+Rk1Ws76bU7UOK
NaI6FV6gqYyx1q+1uv83aVRQNE+8VeibyF8O1XC0SJE9mEO/8eSWNRrYRz2NS7pfe2JrjgK+YRoo
zAG/DQdqHSFUguI1BmuyDqeo3Vl+YPQIUCoVjYeUNYzl6BohWhUGfJacbBSaFrkEt8W275anfBqJ
F/e4ALrWzUdjPJlipQaWB2FE22sT8NX24HTzfDLBTFj+7smPsDKfRWKA/37/w10bJWLcEioblC8h
lxd0lSPq7eVTo6nX1hvZPoZpAYm4fuaXEenVmydq3KzJwRhfFRDEfBf7T4jlubLMP5aJnsOwDUoh
/mjafLAvjs9weOCtDWF0XDPz+d4mSc0UQkOimADH8OBzTLb+OehPfruvTBiSiOJVDvFXM+N7Xg7y
vPufuFDIcC+MbSqJ8zvpuDLt+KEBOnlAqLbqLbKhQ+hztWQv6eKBh1hh05OtWe1Tv0zws6B2PPHl
ATIO9Ie8jx1wKctTJX5PLGSVkKVFJf5+Q355TD4kJNxmuGf5jNuA/R30VPDNLkvQi8kOiysOA/6W
cFDBTGHeyHM84y6sYU8EdJFfj7UjFpXMROZoKTNO+Ur+xJQ42STH/4vs0ADfRl5zV6guP/dACnX4
KOtnrjXm0/+P5/LBMavKpd2Jw/d7ZxmlHaFNNFwfsLMuN3j/duj9IAaDJ33qx4+OOLvPraITTaJk
2t+qCRBK9VyVGTGygpHbeZBf4zKW2w7yurJVhfaXQq/G5SJaWIGhaI0KZD5BaRXjERRpLifYOdzU
AeSK37ZKLtvhHKOeHRtVz/ad+/f/sJnp74XxUJQBP4BZpFNHFA90Hs1qkENT7u9ZmweMOojZ0LcW
rq6aadgfZL9kQm+/E24DEDNAOap9ldqYgqoaz3lJ25G9HXcSinG2YXh2/Rp4WFVeduzfBIExJb7M
4FYiUYAibsd/GJH0fHiurc9BnpRCOT4KwoqW/fmUNa1uhWSne6yM5NjIP5K5iQfbabzNU3NHwTTM
wDvZzE1Eamwbg2P948jshnczrKjN8/CHcD352maePi7SWeqVRqERgfkTOhZ4EGdqPxd5qkx0+hbr
kU2dIsUg6Cmd8eS5hSnMOduG2lV/8PQZ5dWBFhGynxU2mTblYHQj20f0ylop/UlNYldWzaJJHKgX
GWscI7bjXLVvWeXdsBuIdm9yjtRDugTbKa4QBHKL003ZkGYj4z0+TAA6UK53HU8VHZ7Isq7//IFW
iXgXK8f26GBJ+KLhlvSm5nqAwRO3pCWHdGnyiYqJEIjpcSE9/aXsbISNvgKA4yZLuaEkObgOvLEj
s+Xzv8/SygEdcvy7AEamDcGbtvvztOz+Sbo1DCGpAfPSgRTXHy5CMsb8xKUd1j8v5kjRYDZTF3FY
200ij8nxzupAlnwz06y0t32D5oq447zMDh7BFVA7GOkeqXoFoi622mGr8QySg1Fnp71P6iHSCZI2
945ydjImwmYYL4OuPvbPFfpSrmFZwMcnowNqiv+JE9ONGNulQ4CMPukhgN12nD3DrYzpohtr8cNF
HnUgsoaaykYhlXDrmjzZxyw7RBUN/INp3ho69Lb4agUgNxu7HvcPLySWZRMU4+ZKScThFoiiW3aC
74lA9s8rSUukuVTLJQDCJHz4s4/9pBL3xAjKMJU11pDqB0PFNz/gpusY+0jTEi0WWJHJfnKy2TFz
J1AXdEBqz2Es7cZ1sMvUuNzDl2XBhJvEJ820w5Rg0xxcOH/Huq2E8tCEOrjlZVJV1eLp1/bMsj8u
+2CJGOxkM1jcv/lt1X0FqrSXcRl37VWiKdm1Cot9W0LtxBJBMES2+pO06LLECyP8JhEmhCOoA6qy
WHsEmsUugwiZS/uCMCYgFUyR15zrYr9tUPzkWXuFNv7iyEwwcb1J7+kMXERw9799+7ol80F/EH5d
DgQeFFZpveHgCA3IcMxacFqnBq5/pc8vhvCffBeKhxYSFRiGndXt1oQVaTte09ft/Man2a3XGNI+
aIqJ745dBuqRfy4IUXMr9Go065NiPzlmX+ljF+HDbXUC3F2AU7gIINMCIdgrXDrO0uRHkP0pQM8t
k7Bm+6UbppQfCzYOXj6dWQRljmEmhEdZBoe855kymlzAyR0q3IbrCeF1MTqy2mpf37DnKt9qKYwx
c1mBwvZPqwPcBtcI42Dh0/NSqeXXOsSzwz6gQHFYYEgf2LQ8ZxBKSvIzktD6PTwtkqk4uDL43u+t
ZseVgJv0fmhwdd529Wc/32s4AZvNbBnUkJTggZHPZxLV6FdAOzoJfUKduJEbLPXqT1gTpOK301iQ
vbtgnNt2mIIcSwD1jcaH+GGh2MsYc7ssH/x128eFxQFy2QCoWUVYrPQ+cSlPB8LdVkKzluOUTBSD
Q1AKSIN+g/cTUUUo360aGU0KB67eTuFydXeTq9G/zb7qvEbG2FQ/yZONTbKqoTsy5TjThu41EMNl
qDLnZ/kvNSoZxWsGmKUCrrIyABMXCnlQhdRPTJ6dADyhbmdFdmnicI/5gxeb2zn36MG88KUZ0/hJ
G/4c/XVHUb3lenX5UyLN9J0iULowmL9EhVO3utioZ5tTLSqjZ/gyOMp9FF8+3eXlD2Rin8q+zND0
Zzu3kj6BH5ElLN+nqYHzyk4LO0tUbiX0EgZ+JdvgiqFwOBK7YhKUJjwfGOt2gCLhSw6HQv9g8AwK
kCzxEJ9/Kp07aJNSwUt36zWK7FEY9yCLwzAzbeEE+9Cc+WmUhMi9yNpnpwHJPr2qXxnl1PnEmMH7
RAG6XFciz5GSs0X1FrA+XAAf7NrrDw/OkjX5Sn1QgKZVnBBQXbTZ2UWvnu6+hB+EOYBJOg2uIcxy
q8K+waec3D3j/oK6o7QEdPwS7MkPZd8XCfpA4n96Ry4Hsj0T9bVUMFQfGie8NI3+cfwo9IcN7ONH
zsodFz6E3soi3TfSdyzkMvWOVIA9B49leD30YKaIKfUw9Irnk+rxx8+UZgjj12ZhYQ+uVdcxtWZC
+hFCg/huCI0BabLGIRY1xmLXMyqOVlwhqnl62gMv98mt5LrzZE70+DGcb9+GMRKyozz8bkIkImnw
r2MhoACZNQDlv8MzpDFHnjvi0Cw4/h0nXPHaSzpujrHxUJriT5YuWVRevfxHEpMuY4bI4HaYJER3
hIPKZzHSUbKjQNDgYZvf2N/9axi8SsC9dKhy5lIf5dRgLc4pO5M0qZHYU/uBWMS5uDKtr7ubBEZ5
tQ5rYhf6ja6uyhR99P2hTXCG7xsN1OH4uZL+276TdfEPjM/W2ZFtUvoTZFWn/PCBTyIb8vk4LDO5
0ZT65htOpA3iTjI03qR6GxHBXqI8e+qOG9edG3mxYy0OjcV+59UHQdEO8Wld04L8C3wpEu2UCAnt
Lj2jHgHqgB8MZH8k4TnpNjrGOjcjGRsgXoteCq7FXAUcsL5rSPsK9qLRQiPjOsctwDybHV2bxFI5
DOQYG1bBcY7d1W+3doKPFkeRHOilAy37BbquOvBq+S+M1tMmWV158oh/zuA1RxBPPRz9aj1b7H+0
W8OzQRD44acN0M64KsT7sDggivKKeqmbGpc8JkHNXCI+amkDfiS3QfCaSOQMdW7Ct9tOEeMeq1GO
z4teFNF+0EgT3gsTotoHtXWJUj6HhtP1GEFouWkhtyZq2zS81aPEZ1z5ZMwUAl6WkzaSmNoe+oSm
KpRJ+LVVasridLFEJ1wcH4jT4w0+h1cHvDfZXp4nhL9/2sZrsnQq3NATk6CGY1RTLwJEfjT9NX2H
FC21yCcb+Iebrz3IysDes45VnrY2KvMq1xZToT4iIrTkp8dRSEEGp3G+66K7JSW3r5vmQcDqpten
SV9URx99BnRwnj3/dbrrf3wAUC27KsfmtMpe9xa/4UlVS6/r9KWmdU1Cf0zTFONPtiDG/MKVffrK
USmbt1t3izgap8WnMBNrmvTVhKBs/B71ee+wWX/QjhQ6n5pLtHZTt9OsgUjsrWgX9T9pwvq0aH/Q
sFhMEC1saUeZuIfKxOszk9Cyp7BGEI9iY9JT2XjnfA4aSlJGY+VKBTUh8AW2L5NRc6BCtQW6F/nb
QXq5kwBNGGun0x8JPfVGvTL3ExYwGUSVxU2BKG5NuAEYkI1ZA/A/I0fSJmoY95ryw71/VLpEX+CX
92AQMYWs58NFVq88huMIZhZm4yZZj77O7FztgHmiSaatm4lDsmU+H86vghtBbsjGb/9MOlLLUi07
y4Os9kWaVDdJqJPwi1QZJR53xD3pa9TEvjhU9FA5VUgqjbsFo+2CDREukfpe5PVs39vzY7rM057f
N/uNhUYo6S+e1ZPniSWSVuRK32wecaHRpfvephPpvjB9hzXNKIJE7J0PofVa2phgsOSBE1Rv08pJ
p9g+g9Nr+/0nZ2mn83mTBakWJPDpkAsS8t8XvOhVc/pH6kIIAs2gL9T3w9MYLlua5XKVISJno+Qr
V+OLSZLrhLCBHThOR9QWYRF7Qv0xVh+EfY5Wrl3d25j3eqBp+xrWP8L/z8xqIVxuhlcnQWcMVklc
Uq/8ihd3vRy9uEpLyh1GC/9zeF5D9T2AhTp1QXaqw+gBa7x7sP7QJtiXRheicjRknSkvmFKb8JMe
tcSs7Tde5cHR2wKO3pfQBjR7cxmLGHtXRnEA/m1JgGAjndlbcfVxEHZyuDZKSITCYXJB/5ZE/BiN
NoNK9tTEc9zqlWhSMd0Dktf+72+xTCuyG/LuucN+8wPMyr9qTrmywBd915+v34772X+62BwNFOq4
eXBMKG+ZDqMPZh067lbdSGPwvps/dwCNrybKdEUwK7z5rWiHaL7biboyHLz8sUw4iE1ufDjeW1rg
r8a/02IDkjMZIBxp+sucHWe+6TDJY84QqE3RHUELlatzNMxu9Ch2RVHxS5NTg9e8I7bx86Ak0pn+
RFpgBImNPg1T5usr5MJpMl8WuYzAI5JDP9E+1taU1P1q/ZRNRQZTgvVaIteFx2Wb2LtH8fqyMSyW
KaQi9s7PYQUQODCd7P197cCQFVpA/IiH1nlVuHZz/XJwqM5LsVUGh4D8S/9zUNOql9eqDWImQKgh
5/iZqsZ4brWvSeFFgPhdKIw2xIV0JD09qQgLUw/8ghiXnGUMc02BFKVMkz72N1fmdgX9moEqP0Br
WQOsQSPR1blZRvWsbXBYcx+lD4nLtnW0EmidNkO4IOa0siNuQHjys5cm0vOpeUgwmLGv22j5eLYP
ku0nPyIHg8zrra9DPshn5YfM+1ty449iZTmiiE6cYHs1I3lowB/5EWxEagrYHSpSfxTczuL9JubU
pa9PjaQpA1DTtG9qPxEZELG9wxt36aSRVrIMSx360dzqWf9dG2co3/S5IBeyWRpYYieoMRokKmqX
JJQ9rvV2FsW0cTvFfc/XzypK1TzaqLulTDHiFYcT5CCPSDaKshDmG6SdleAVmlyw4rxHKb+pdUT2
jiaCByo/OmaPTo1SsPzg7RmJp8sRLIuu5Ta8EYds9NpZMbeYyeASS7tmUKQTDw2I1GJl7mzyvn5q
2JnsbvZqe3Az6fxk33y16+9V1dsWgavuU8eG1HzpAcJM+XUybNMofpeZ5M47h/nVRtTGTQ9yvomT
erR5QdK+RMjVUOlpyYxmUq433Bw7CI4Khh2C0TGyQkHoxInxU3dIAY1DLtGNyNR1y2D5PEDYVnd6
2ibpiW4rE2CHGBjxAXNaTx64kTXwwBpTaPQXPxoj98rYApFP+OnsK7DvD1/1tQjNcSmPDzPmxG6X
N7GcoGghGaGy5bnq7+jRXZIpwaitIax8ID4N2nBhRYfbmxX2R3ncx4ei9PODTq6DHFSwNZd5Ml0L
XsFcUvroB9N0qodbmqbCygkvEmXCR/8OEEN4UVZP28YXPTzp3AVdeimdO0UzoqYqlmMX6GYyQa4S
jRfF3FvLylNHgrFeeSpN4wQ7Qu9xaQul3j5trWMsrqWXxNlEjme6BtTyKUym4QMfqAT2U0Tyf0we
8vPjrXl0yXxed/oslUPPZzDIoDkQfQjRddwLpr3XISBFyBrgxNBCJB/KnaeVxLJ9xbTmgtwvg6FG
vJkRwpm4wewMecguIlPIaC2qbgqDGgVAxfa5glpUYPbt1G5Q62tB5/3zWjlcx+grGibVemBEBYv1
QJGoRh5LTLCArG/RCh757QtosifmW7U4prZm/XVu6jwAMNgW1QU1IkjUdMhSM5RSP9ofaEJH2UDb
SMkvhXEgF3Uqu5Q6aakUqATU2c7519RSALwFuiq6xLYa2tJrR8OV18WAGPxFmbzJQF4qU71/SvzD
vrnEf5xxPGVcsi+cWfQdtTahinHKDr54Y5jUBjSRQpQQxNxQPltbMghEcR3Hb25RumVRJblzGB/c
ijmP9NUZtKudZRwJAEiR5hUNuXbmuF/7puDGXKRPAxO2M6/zAVzki+4HM9IjdCtyQ5hiTqHIL4NQ
amkfNM13u3oaH0fO2Bl6b1wLVvm7XIcc+J4pN8QVljFYYZ6HPt5JPYpduFwOZfN2UjFA+X71xdpB
/iNBT1shxissB9n6+8EBmXz3SVVOKnh1tRVOzPstPida1pI7GAbQGtk0nuDfb2gvwyh8wym6naDA
3N/CGXhHTbqkRQPD8iSJw6po5Z721WY4kXNXA5oJQdN9oj45IMPyfHgiKpxm+SPFC/1YLLbfNx4F
RO/0qYGLzMvvp2RYU8N9C+64b9Sl056MC3it0AyHWU0nt0LOHeYW6ub+0LmSKsgsvaZZjBroR/Dz
4OoVMxDBNpVG5NVqPcoRmOTnZ3AaDPajGyyoyMSatECiwNrb//DBAN/hJvjIwbdG3WA2d8zA2XCm
zbiXL3zM/mHZmljSdavILhWFNGknXDSxZaVH1heEIMcb7e5mdizBLnIA5EnbqJY/gS+nihRVfSu5
VCkl+3buwaWY9KvTNFC5LanBYSrnVDjN+zjZBTijc5Uz4IrhDqfGfI9zRz45AjFZskz28LL+PMGl
3TcvYCA8h0FGnrtgFcvCylOqH7kYrElTrG0OA0OMS8DtTKEpmKtBdYfQXpME15TGxHBEgygmQr5S
pL5k6re/ue/szqVsXjR5+IRgnmbDPsXnsntHenRSc6DeqXCU4mdCO4rWsB5Zy+q2tXzzTBB5Nism
PJt7UjKSwlDSofNVm/afEJhAY57Xxx9VlGTaW4PuVt+5CabDh5U0FCqHSGn2YDZjZinoWDR2nwVQ
/wIxwhabhvWYyriAVZO/OJhfNVp3+Br6xungrrRKQXZRG2HBJIcb7JyUQ3TtSG1fUxt70j4l6dK4
okLFS11KcBq8Kmi/xkCwCENQsWm5L83irCkos+cUPtlAsz9/WHHc7ueISzRM3UsQHA2GnNFo9axH
uOKRvUrBtXjuF0FUhRjUiHfGxqngHPe0AKJmChdofXsm1uIn8tQs451sPKF+XkwYeFqMA6x05pmo
D31j1R1Je3JeKZgsB4FToY8G88ICj7r3Iq5zrKrz+rHMiAwxI/VT6N9hYUQsMGj8XVFvVqYDAEta
u7b4rIwnp8ywAojGRpbkqIzryFsJPd9CgOlX4Khirkowl5OsMm8gnd1Sb2CtuClwoF4tGVw0H8E8
I7CVukBkAPhi6YkSfrQVpr7ooFVS8yNEfBBBDMm1VtNLyTH3ZZM+c7t1hKjmlWVS7C3Ij7uIdC5Q
kNrFkNZfehp46H6n9jPt0arS8OQLL9VVwfgK6RlTa93vh1zLzoVHjdgZIM45n+Bp93CbEcsSG5rP
r6nNuZNeGVjHZyG/XDDkgJq3IRxsoimPLYqW4PuXlFP7LqoQbRXLXeUVWTcMa2RpdjCiVTqYZjaH
dUBetg20a3Q7KAmPzUvdMO4Xx5de6QQU3LVL6xGIvZARLl8U9IEFta8Syko5Y73wuGtgIYkcSPEw
bTMAFFE9qtBsLMUNet2QBgsL4JktvtG5hQJpXWqh1jYeFa2BoMSjS0qLTvYRg+tMjhVNM0Am9vEZ
LHH0Eq+SHkkG2eH/e1bAmKc7F7qvAKOUInAsi5aZTDGTKSbnpinD2+tkfHbTdQDWSGIYbBDTTCCZ
CfqdMVejbaJobvPu4X8+iAgaYfgnnOblr3Z5NPdEAtqf/n3UBkbXmPmM/4ec9JcVSRLBXu/+vk+y
hF3+o4YoqBROqiFCDxenGcAyCFHOx5/6qKoyzlSipvu4pkXNCwodTkbIm/UIBF1odzuf1zAipFTb
K+uHtBEwc1MgRJ64EBBu/Bpt2jSj75/nJXq0NnB9/kFTilRcDQ8fSkeN+R5hhfUjXbxB4wUrrk7J
qtjwL0Fhw4w5iKN9ngA7uX3vExsedr9rqnEQ7BAXMWAH7CMXi4wDJcS4Ndd8MwyQ/vMOeG2pUPw4
tiINm2gK7Hhh+DbVp6PUtIswdboyjPP3m5zxx5SfaP9xTtlbS3X8LsSoMNUvYRFT12me5WcOF2Y6
Ki4rL9rldXAgXNcAWuXjTEuP09faPFbGvcfICq7CNRl7+Q85ZgJcHHWsleaeT39eU1bNGDuuMRF7
O6Rk3vRwmNeIY5ZZMjlDx7xX0UlrVOxW7Y2Yf5QL9Z8pMcchlPF/WseXhmbhYJ33WTyQa8234NTF
SzDak3Og25XAHpnKVsBFOwEPj/G9WmMUodE9eBpzE3ESj0je6vRwSN0tCIHvqkDHHu8UfDAkLQId
dLOCQUL65tIZVO0UKMYDH7zCY4hNL/eSlU0NzC/miR8ZDh9K80pKEzms6ed1+luBVIRhGPLWqx+M
qnrU49w7822nEcmY2mP2WYG70QMJGoV+s+eUHiHqFc8LczsK6yQHLY3KkscKt+/U+UufTIlLKw6Q
9AajaescZ48nKe/tr583EuAMTl59RZQGVKp3G2hjUS7U34NTr9gQ37bs1MpdLaMz/qJ95JP21Wrz
4oEYOmWWEA2V+UwXEraLY5SRZwkld1FXS4+WtoHST4VhOcniX8w8ZjIoaJ7tOCqYcM09/t1Jvbg9
xmB3513248wFu+bTtW1x9HAh73CCcUk2q5nHB/0YOXFKBliZrrEdMtfRDvEf+2KfM9oKkLMD1IFL
0y/BTewgL2PKnfVEiw0jQaZLkyjZojCXWLiIQHfgkw5A57CFB4xYbIjv+CY2FAsBMSUwJhcw4q+f
CARWItPQHXIsJkBR352tb5xqwet4W13iI4S+g8Bwfz3S2GoN5iOSYGUpWjWZ2Y32l1DyEWPHTi/z
CMzcXRAiJlaB8iiZ+avBM62wIZhX+cAcTSBfu4Aot5b24gz7aKa2oV6xi8RvQj+aZ3Few6bIoRSM
MnY9/guMWVEsQJqUf5m6t6J6EtVmklORf8g+3njGTwVbImWvJwqmWDlm75RDBUUIQxLr4oFH4vJu
9+OGiaWTxfgehV3pGsQJS++XaF8uQN4C7Z/S3pJZmYWWXxFlk72agPL9KGkjzENJL+sD5sJuD6zj
QfAAf9z2wSe9OUVGQxJ004ug+kkwrV/oPbtas0c/BtrUD7yRaM2VgKQci99BRrl0VMlYCura9yHc
57d2LNvG/HzCm0TZnqlb+V1Inydf3gM8V0hEQG/iDVQJOLirZeC9QrM/DNQFFaU42B2MrtnOhyxq
LZqmM+MWKG7iGMdZ2Q+HDzEnaiOlg6nTGrR3fnSUHANRRkbR0qgHmPE4Ox9bEdQefnHMjQaTTqgj
HeWfdX04zISkjhVWe43N1wSfW/FxG4sLZscNPufHylWjU320bC1wTr+5+vReCCLcnymy+tZiQruO
MQ3jD9R5nK/gK2nfiJfTKUD6z0rVOSXRtghVTMrhFpBTmvHA6PZs/RMqR7c4H05izihS8eJAdb1u
kGVNUdAte4nfHf8yrJDSzyUqqs6zi7QqwntzjTOpjOlxMX/zrV25fHvUHIOeYL+yYO6MaodRyT+Q
t65Kai8E5YG7l1PIyyGgqfDUS6g+6tSr129c5Qcrnc/o+yKFbrXM3obLIcTaJ8TbI21xxMXSsKrW
lQ8M/2B62EJeh4RELyW6wjlbsiGxGTriKU4yVifPsIRJAo+PtjHMa03pPDFnquCex3bC8dV8/B4F
yHmUKLm3jsbjYmtq6NNveqNCTrEjx4Ly07c5yH5RYXDJ+han0G6pyUvDPR7QiXC4n9DyFcyLPLSt
m3E1tyQCfVAjNg8BNEVSKCovYDfOpjKd9xbDvR5S3dJHgp6N7amxlRfD+smL7QBkqpE90YN0Plav
W7P54fKI1XhicUQML8fNMlWK0CJHQwLkbxoDq9eFXSzyI5pm1RPMyThwsNFX7Ce900U45zAQNOQ/
sHWkhDvvdrFsGObRdkicTv4xPdyt+MO9/QXLWk9y1eWNr9YPFg1hL2YFxfc4ETu7psk5JU0Eq1Qb
pRqT4Yzy4kJIhevtrdzgpAYkhgj+J/kqiaW/nP816hUrakxwgnX4LAEdvNzfGArCKbUUURdMFLQK
vgUWsIBiuWdSBqKMpu0s4F0+OOOccUYpC8EiU9aa/qVqTJ2KnpQn0OT0QXheUlFqCk/TlqSdNhf0
I3NM83NH6FEDO3ZSiwDte/n7uzMkhVJToP0VqifQRfhqvYLI7wL0B7phEhTDN10IGPTn1dJM4wwr
DAL9cA6RiMv1IpgoXcdtwLu1RwMCAtiHvPnR3G+Wb74Bws2EiUgnsYhMmkX/Uv5PlD8BrUzbFGVM
tNWdc408PyXiubDN5aESHACW4MxfoOCo2I279IGQPVpWPxjHmuCNHMma26uY1fCF1NipJFynuY9e
PYZWDlvQ3p84InXJqCu9zVYiJtu7Cn6KaC9dFS72cbZszkwsb7B7/zGmIx+l1stmcLKm23KCx7qm
CdlxVQucBKLWwgSN5KTqb4MuqMWwFriMkmHhsRW2UQOd+MKnP4hjWphpoQmwWe3SKQ+fqzIlDBoe
obNkOeP4PfXj9YMCwh4/19JYJnH9MdBC3WB28mnzlrPegUVXyX8B3gJY2KSqR7Wa2Mt+3tv2sAQ8
fQ5RJL3fELDsSs3RXnY38QWoKyxg7ApGtQp26HhXF+ALloPHCau00tp+djG/mMGydW0rvKqChEMB
WozfL50dfWBVhL+ewMCXatIYSv9UNV0u43lhgyR7AiGyZ/2XuABtSRBUVuvSuD46ylXmCEbeZE+J
Sm7mxrOdsNvUdDQN5b0V/y+EDku1fljSAHvESFpoLsQ3mVfrjhvGPnLLQhdJW8DmreQ4lsGzHPvS
z2TWaEHl9Qmr4DknI8zsqhQaGL4g9L7s9SZ1+BaSMqlgi4wQGmzWOZtflgGIQbRC5c6BOvc/dWBr
HHWwQtbhJNxlQ5fMCkYKQpElGxfAry5SKhq6g3Fz1/dP3uTOTcHz/4D5k9NMyiZEfgkCz4IH56ff
IJCtHnIVUaBF7cwgPYquzV3C45G94wmHRFYiI2szq2bNwMPEn5CQg7PnYMmWIlUYlWoiwtHboZoK
rGOcJjEmheQF2lbvCkpH4LY2xz+Mbx3BjgijdFSYdMkjvugp7YYaHP28C3pfd3f5plQX8qzBVt9J
zVCNgwkjt/MdJ41Nx4ZseWoXpfCmUtXDPLe1vLRV9HoTs6+U8h5vqjHWqui9Upl6dAJ5cIpRZv7Z
wJya44qdgM0CJqPNyKIu2L2/S3WitSzosS8WGIkYQ0aSoIh39K86o2UG3iQiQfHQVEY2lj/ObOKO
PH4scoaAWefYOBOhYJSSx+JMxYxaK1ukXkKQC8SbYxOx+7YUj7uCFqbesfE1ECi5dVoRSAcw04/p
lSADpLmngNc0N97Qu/B0w/VQv+8r/9iA6ZMelNkCL98hcH/VelAxJm9MhMxqfbLBtV7sDAoJY9yB
3C09NRnY0VAW95ZvlHe6+ZfvwuGoPEqBrjWwhaloN2yRR2H7DDhej1lr4Tka8YGosg9Z3zv53/Ie
IMoom5qYwuaGvhXpoD+Fy+YQZ3m4eHI2IGnVC//5Lq+XFxK+QDIIOQVCTaS3JbZuQoMR0213FLJO
sZkzYJYgza1ORD8iQZdGWRGMpvheII92SArsds6nm14D7ofBzAy8xQNXlxaAk85lwifzOUVt9JID
hYl6tVAD8rYqm93wJENBg4K5og0idIbWHqdukdktHe+78M4CAnP4NFYVqEP30WbNUWJPFzfhhJeO
r5Zfq3b0AWi/zRasKsrAkIQPTmjNCQWZaJufcktOUfPDbN1Ew+kl54OrPpLrNcMX14pumxVgX5oF
c5m/5Ze4nSYDlYc3jBYkTfa05da3phoPevhVz1yFn2PpEgtdYHODHzhxLOY4wLNSUlzAU50l7UQh
5MRoTqffDGb+vMQYBTZSzwcWNMxWrtQBQR3vlCvEGb3wU0MLgN4HOggGhG9oPUacPjnASBYCuAMU
5cHZkzWASHfKD3tKi+QUxiX/e/Je4R25o77l0mWEUMiUfL7zvx8nCfm5clxDUatAVplctw6c9m1I
Bx8YvVQoP2hzth+9eEbXaFDeugqJPMkkavgaaFtauVEv4g/7+PE4FHAN3rnQGVSGjeIefjsd14p2
nCrENueC1DuNUeB6/BwAuVE5trI+GdP1SiK7PT+smEyApuFSpdq9fCDrV1Muvl0hEsPIZC959W1C
fFqe3FTjvWhSVEPSjnhUrU+C4J1cf6IC5CImbkx5ft3xXKmIjMstw0T8oHbO1u/B1rClpbZ4Qnfy
ycD8EuV/7EWO3S9PkGBl/YypsIpVEHNuyi+bP1+QGEhveki/fVhI/53RHLwThPOkK8+oTniUlrYl
RgJwO7qz6nUrOff5dvZimaOQ5LPhv5Xtj6yM8uOtObu2hwAg3DtaB8DStXpBaYPrkgHOtEops9Lm
tzluegUNzHhpBcvtL4vhTbsNC6+Cv03eJ7JnvkoN3tU/DRD7QRFGXuSprUdkjDHXRGQgY3RclOkC
a4OrnDUJpjmFcDVtDHF/qhyna3NEM5UwKF3IwGhntPSRUeQhYXoiOTLiOS7RgCK/fw11IZ7Gqu83
wsA3rYR/gT1vggqYmfn3QZEijRS4+JKuiW5R8/mD5Y9v1Wahbf9jl/HVHF3hFWxodAfktl6HH/AP
KYWK5jCReyhpv2zAFUDNsXdiAiqCKxtVGV6tM8FoJLUAdm3Osuti1KctEitTRV+hx4/oYJWq17GD
UxpT40Cw/WR+pPvgweRnkWwDHikCDNq11oIYkg9X09BM60sAwLr/J0dRst8dHSDQAN3QbrUwL8ok
W15KykO9OMvHeCW/SyDinBP/R0CO05wtCArcFSdCKmY5vmLVPKdMTdNDd+0p71KGW/dldbeb9JKp
ori7ipo6Td7ULdekK2woi25TqPQVKHzBEt+RpXWMh73MrGPcdxI4LMkuNa2gDeYnFEC3SZlxVekJ
1EQac1g6DpU8sg4uO3jx1WrN6IIa5gom4pB5q3Ifb7oNFQcZDghs5tR27tIsdLamXZV2bsJWQObV
7Z9iFJxEzdQsWkMSS9voEy/JwVZEvtDeFXak3F2oVcdXggJBUmQrNtq8oXXurizvWp82eBdJur5a
PkTZklCpGTPl5uMFGmsugcwKdfpM7a5hAsUpNRz25avhRSJYesds0WNUkpAmkeiIbeFbNpSI7cyX
I4vLYf+qYXqpNeVOnMaYDCym2H4IzWWjF4I35O61eheYUkUsu+6lhSj5HdRQhmvXYsxE9az9v1ys
Rctg9NRi8T2LMDbRYYahkhWoEfU9bgDSS4aSZkHOJi9pRRFe7mqDZbqZMP2D5pYOwh7ns5WlBcp1
FRrwi1shtrqazl+jpgdFOhQJq2QaSItl3SA9mdJqXzOAGUoF9iRvlU2lrtW2snpOufkP0CF4iG1+
PRmIqdmWysv3dxBheRjuci19QPFOc8PJI328Myf0Xm8zkLyxTof+B0ub5yUhTqXfcoOZIaVx8YkH
3+clVD2faONabTpqYeiZdc7fW9tKWRKRajX0QYX/Aol1G++bHC71MXxDAHmQTqdry5LHLMgKlEeJ
qPZXVnYCRxpMKdusZtcQBLv8iUgSB8xA+OCsNVl6Hy4+/WmuTydVsV5E8Q/3CegpHV8VXjDGKhg7
j5wgMyO9HXVg3ywh1Has9X1GpFzbCTnikMr51OPk28EnNKa44afO8dIE0lB2D60yuPotdpvTRq3Y
wvNmaIXYTnUhketqf3HCanNca9q5N0jdzfCO00WPY7jMAGRw5ltchC8EgYdEHxXEMdhEMZUOSAlE
/oEGDbs3ddiJJ3rdE1hOQLEJA1hocroz+wANBseR7mSOso/ad/yzVMyJ/S+ZtkB3oGkf1NXyPfeG
1o7wBYp5Bhiaf6PBBEPO7dsAuOv2WGewgl3Au+exn06YVtMNJmtTt4AVyVvS47LwbqAJbsIDWC6j
qlkdLL0RKZvVnkRJx5SprZsR2AK2Yq146E2pVu4pW1t6Z9clIdHIhrv+cfdGNDl6oZSuRYbrxwRp
Iff7Di3kCfqAIvOSFjC75NWbiqbX5RJseey+UXNzxx03PjSnBZtuS6mNlvYUpc154nw+7tEK1Gg5
ugsfb40n4LdfzTMkA6Y4iZj4aiL7R0JB4XsnwuTdMzeqfURdlhjkLZfQiThRxBLwIbClMFwPeNcQ
x0Pr1M/AJmEfjtLtMKZgwzlOV66fmtkpdG38SPX74nbpkD9TqMQPxMNbV0dMGigo/xZRIQ9e8okK
aDHKDSz+4rV0jrZD1qZI6g2n2UczU+UzjRWMeW1z39r7K+PGiTmrJpRsnE4tfNjzWftJZoUMuwAM
7J9Q3ac2l5zSnpohEkr3l/plvGVdcqesIdvZFgRVieLTw0AhXlVyG2/I3MnOcY5JqozDVudewlfN
q2zQt167GdXmfjlTCz38F0CIEdxMSssOHLS9yANGVkqmRV418vAhGVy1//2zaGfqu30nNkiACK+X
jyiJGNfKSKhotpdwcZdaGkhdEG01O6i8BZ0h8sOBvAk2JUGJkf8sP+qKXYh3xMGdhNUhb1kGN1Ld
SP0zJ5Zz8BtHfryHdN4WdGOYUsw9To5YTSRMCl9JPGtlv2uHWun/AfBkFCVUZaEMBklknVgVoKZw
UoEnhbHbx40rJVr0yNkbasIQePfdmPRZGFfV339n8pK1qXroI9umkQf5E79JtzqVn/Uwhioel1Bu
Lz83gEotIvTLjPlkPrHLgNTJ7pLopO5++A6v6t1qNuWrsUKA4pcSgNlOMAgG6Wl2TpUzvWZwy4vd
iJQvZQ9dnZf0iCKgOcAqaIqfq8LeQSdjLU62QJiR+/cIupE3ta4/6JJV1uc842VrsXPV4oSXfZa0
wHG8ZNKUI2N2Rkthzd+aRYG1q4q8lJLQ2aONyyoLD3N3HNgalSd1EH6l5RyACcJkCdmNMwho2hed
7Di3ITXSjxvw/1YSvC9CwXow2z0NCXBwaGbcQNPj/CONsvYYmzuQN1kUUWQfnNlkBibyEs+qikFX
vUderxB0oRgejwlD4CO0Ty0mDHfZHglczPZKl4XiDiUWlve02FITuQ4EN1lrShsw9BliIDfdczhD
yIwEK9IgCnsJ1DgVXr+TwDPpFbxcs9QrAm+EMnhLR1BUkVPpZe4+9EnPUC3LVUjRs03IE1xLcmsN
q4jvo/tQZk4CHzpm81MdCjxrg2TBgMPigpcMioz890OqId1HmFFDemJwjXyZo2ptB6ubPxb9xyl4
/3H2pK3led3bdFQ0yLUE+gmGRk7fZm2RjzcCGcwU+fD+Lnp+3vGQhtFIxtNXJX6kdY9xs1xAxPv1
5P44/Tie7az9QTOcuXSncg9WLRWj6MfbEGlZjMpyz2W//99yp9YMGR6IcLZ1TxQXwDOqLNwZS1p1
JXPbH8RbKpC6/rI+8LZUAMv1PFZREfpwmCy493rJYDJlft0etzTNzaXdfieDo3++E5yP/pRkD1Jk
QyuRS7+sGzoraWVB9gBl/QQw1R+AkyeY5eJuIRsVWvnCUw2r8WmpFP+95uHPhfc7HrmbpDd3QfF3
naVQ41A/9kHo0JtaNdwlrR2IrLGHnqxIlLw7LEHkX4NJ4qlg1tGC9YWCdRnsvJt4yPNcqD1KQyMw
I4ghpNew9YMD3LmddJjJsNPBiIk5jqByZJxU8A9G0ZOwPBitH6iOKoE6QWGahOz8lfQCNC5hEDLX
VPLlRM8mtPqeDpSGWsAwMnE+SdnTfLCgkkXXJYLWMRrkJnJzL0t6v/Pcy851GHH73d2BJ+z0px3/
EsBq1tA3yKp7LOB4ws/bnEXGTsBsohrQlYG5ydFIhQ3lSkN878xHjVdvj1wB1f81KmOmUxUs1io6
NcxiaHQS3il5dDYzF7TiEe4yarQ2bwSkTEl592+W541o8l+k0Z8FGd6HCqhPSBWOrZdVrH5appT5
nklf/Q5mAS6bulT8TOiFbEKhgbdiCCD2Ne2yt36ZZxPcxE8oYYpEadaVHI9aCZZ9a8hRM9IEw5Xw
CSuP+NHP0ipmZ8KoIQ4ReVX6nUuOKgKAbzH1E5Tz+9HDumTAAkrAenyCCnsK8luzhIFucwksa/4g
ZfshDGJ1IruNQDKGDIXK7SGvIYIJ8FkqI+KqxLlO0xmRmRh8pg94+XiPLrHJWFDlnIHXJB8Owhad
Mgvt0t6Wz90Jo+Bm41+g6NpJVDw93nBzoMD72TOTsamsPjMU8wVSFxHL02o4ATvy6O16jrjciNkq
db5N4OD0qsz2funnV8wS6IO3hl7vA/qQDVJ0n+Z1aRedNrtF0SkIpSeEuslBaVHkwMh8BRZMVu98
0RWn9xGfLL1oaWiwFngLpKFuKFzHQ2yzgp9GT6DOyhXnuvUqOReoLUySW5iw/0aGOsst+jIkE8dB
53TGktPIm/a1oDhLXBCSWItUBFKFETiPnDP4SACe1hL/QP2VB28mHTz5UF7NAvWMKF6STuLR0u/h
VWTNdZOUxsAgLP+Jc1w8/1HT7B+xhVKo6l6zpIGWw+nu4+ULcoJd/SrQ4UlbOPWqhiJpVaU11KAE
HgzuJ8GDRhV8FBzugt/pI/OBzf+rlV6gKxg5QWCHNhHfkh+8heSb8Gcun9yjoiu26KlbW+BlpLUx
HVdlO9Vh1dA6s/djPFehkPBA4yP6zbqJxo7x7ETkMtoYzm+0gc7bOXbF8taoP/0bVBhZzVd59met
JvsDHCQf83AdSFPrulO19maq7BWl1Z3MRHZY4bwkILOvxfiy78oSPN7clcaHY42oHm8yQGzswlWA
ZN080qNAPglQ7v73vMh6CHgmJe2nqYh0TwZk8mB+Uf1nSFq+02muCqhLeEgRpZS4wdzRxFYGUmlk
CnhWHUKxkR/s3bX7IKKeNyJXQM1Dlw8YU5xXFnRXioBhtSI2LSCnPZoeATRVb5SMX/m1WSOM7as4
t4+Skp/pFXc4GAquvjvN2DGCwXDQHuKBs654vNZ5ii6O8XB4vvZ8KJVY1olFaybSJEzFGhtG9ADN
D3dnjXFDGMKxDu8T0xlCgV6LaDS13v9OZwZMKZDd55rxWNY5PXVe5T5zAuE7kBGu4CVAHU7kBswG
6wGFv8COg6JdyD6LS7mJCo7WnxW0PF1ZVE/fUNCGeRDePmAWAbU6o3C+vWxly7fhlFYiyo+37a9m
Sc+SRXEXSE9+CZYWj0I7ZVk0vcc19Qc/HYjb/9dTFAbe4NPJ2PgY1vpg3dRJamvR2IrY96deLBKe
3yjpVZFhjP5Y/ZOI8lJrJxwvdWw42SDBa9WqmWtHsbp0vn4SsVr0JzdxTQO70z4VSyZqNK9qhBVJ
tzQgMenwK46Jxru4xnY8uNduZZNb2VCUm7g+02NcWsoE4BCvzRAdZHzqn6S3LnFi8IFDcFfRDSVQ
iZaVNj1ZxhwXtDHxhlKmgoLKGThCD3PXM7C+mniW63PYPO5fpcouKBSU6FEHKpOo5odyokBIQDAD
+dNrY9EsAykmLT6b6ko+FzWQ7w6GhMV6hcdj2RRw3CAwKDdwFAEv+IGH4p+gfehU1XaIYdrgDs1l
z/cILBlT4sKyVwD5lkgdqXF1CQv5UcCEkksF2eTozDuuPv2VK7vQZmdUSdoz7BvgyInLczzSExIY
mkFsRl/eHsM1ab7zHP5yLI3HmXFItr4wJDZN/moa2icbgSpJneI0LAOeXkbXdeZ2zXziJcnXyLfL
XhGvBVjzna1GUcHknLEB8tp8YZfX9NR1ZJ7XADdphaYuUx9ircmu13nGgVXkP/ScKpDNkx4P8i8K
ahcIAACtBvnmmc/3vUa8ZuCeAjTviUEC4jEHDbqKuQzc9MNXoIJu9yXjyVUzDiNDIUQUtwsy65/B
fPKH70N6ijk3XFYk7rCyXUpuzKJu9qsD+WrRpCTE4WZGkoDedh9LVPvfugjHZ6OH+2bR4CmOrzdi
jRBjH71naV6pa12e4c6HIwTG8Fp4afDA50VjiULMJIMztNnMj4+dfcwuiD1DYmQVmIMZVrQbMmaw
gAdnLGyDtBiAP+TD57ZGnF2ZKBvDPW2CgYkXAA4YdRKogWcfXkyDonSCoxRZv8Ule/rgXFltD7Za
J/wumSlXzJVPyDdmjUzOrqIPoL83eXTE3PJ5O+lZEhOX0PMNf1i/uU/iv09+CAB/maS0/aSP6meE
8y0cuh1sjVBKOqLJi23Sce2JrPAB49p/2hAl7UGHoAzu1zERntZyqdN6tL9d5AvuRQf7D/M90IzT
jGfcDfv41XyEDon7RhngzkBdnWQcfbQtzjnHIebetGuzqUiA++dcKod/tozyc4mX3wKNId7dgThl
zL0JAIyoJymZzm2vzHyTBev1ITf7RQnTncb6POzQ/Whf6Hb25X41iSs6T5XT8RYyy80SqTXdtmxC
UIVv5TGQWxjSCZl8KjMqHLxFP9kTIEG8N+0o+j5zWK09+/l2n6GuaAlWNEay05YWPmv293KSUxQq
67N6isjmVJQ1mwRcMsSxqeHHBccOOIwmP+7vvH4FKsNdo5qCo2SBR1/+P1OkFluwetLVK2YnimpP
MH3n7zUrXrVPFc9d3yTRsPgSYMbHhZQLLB6OWiQwDgfU26R9CCIDkeBMA9XXmPG6mgKiyFMPYlLK
roQuQ7LJLe7yV/MNCBcoLfxIJO+Jx21DxkqhDmWS2fZROuL+KVmhVzE+CX9kXGGaDjguwgp54rCC
LMDT+nwSvi4OFVvdJjm6Iy3KjVIF4ncmXg+y/CbmB+erbRdQOQ1VhykiiPS2bsyXYdEaKdwUFMkr
9UXUDwiAyK2F+ZBBJQSEwcl9MBSzuSYGjqZl0OwwfN6iuDXRT6vwTeFNISE0plGTOgbj0qzsCa+B
CmCM11/bfJB1WPEphX3ytE7g2OSicmh/REk8wE7BiOWUIyL6mSYI1H7LXLVC+cmJj39oEv3EwLQ/
mrNytiQtT2WveV44l/Q5NTRl2U4cBM9bu1GCooF+yQQnCc2tTYMGjDCn3dJJLKGkgDwDDhdhm4Bd
AlbO//cJe5QcgbcyX5mbcxaOhWA3bQuEWdeUQ4da75wJ9Rzb7IPQxaptlXwpri8EUnQoUmzPfYEy
l4r1HpiL8isOkAaxSIijCY+sOxo/Se13CaWJgBY/SbxyQQ1eqHezAZvfc3gufDBCfmXyMnTDhSUd
lao1FaLTqg6pyVikBjWztJ6O93AH38OIBmRmqiyyKeDhQWBwSEpg8nGK35WtDqYlGE3Mmya8mg5U
VAnJ0Y+p1bylKSRKC+VRrCaozVJk7Lbakn+40MuXIhJvMXAO5qebRkLIqkV3k0goKy3c4d9j+S/e
5gM7FmxPqqHED+PKLXkW++v+h4inS4Gi4d+yeUGf1QZ1HM+EjFTTOQvGIuWoBu12bgq8XLdN7TdR
TgQo0exGvhUkrrGZyeWiKuC5VqO3lOfyhj1JEuAtfZubWaF89rBMYPtFTb0M9ktf+kEH1+sKhkp4
xFeblxYegmD4+4qTO0yhM4c9XrMGH03gODzBi6gOjoatwjsIjLEtaY7BlCukMAOEq9x+WXathFmt
7mJX0CEjXckQdZfKnOqJsePCHm/JIu6dmE5ZjB0xbcPJqlIrtpPtqHjEaXQU1/5GXp1UeHh11WCd
nME8iVtLxFo/4mWMrxvS9QEU5Ck9hl7d0Ok7XYAhqlhfAiZEO/NVOxs68Zxl0i82280jmzl20JpM
3oM/1IkeIcat4mJs6bDMeLH9CoNk7TwVo6hO0hxcKee4h5brMWynV/vdoNBxu92AUiWDOf6GLpXF
SZG2nlcGamJdy+m8P/NNgQ8uU5YTXOu/vq4iPd6Zd8fcdKDb7m3jy1SfDnnk5Ld5yQYGKz1GD4Jv
mpwMVu5O2m5eRET/x3QECFzbrKo7dFwWbFaXQAsMOBJC8qM2I2jLgiXmFkOyVeHvhZ98dipE0OHS
z/JBnG03Y6DKaERYXKhs/h1RfTal8hX4DotGd2BFk4QeEA3X7WiSZXvyW4z9/EfdcUCyuzlMHz3s
bYZNwuuN+oYIiqdl6NBPMLCVdwNKJDdUXqzN6N7dyiZ34qqB9Ayio0Nn8tsgkXyZuz9SarqIW8ji
tpzxxvGAysqTNQl7XFCfBHKl5JgCMEUOqwaMW15b1+bxTcG1XvS4TsN2ywXo8UPhAuPYMM75xfln
HRqgIsNS9YkzH4pvKcg7JeL8eM9cXymal60DosbWoOUX/IMN4SDANyAuy2Qz6Ja6qh++hqJfv74k
lFNAWxI/kOF/u3RYrRZtiTML/HpeqlWgfMWO1kAwJ/p2UH6djLp15Sjp9A25YKoIS6bJ8Ns13K19
6mE+d2mDLf8+sJbCQWzdbH/+RFvXOwxo6lsD2RIRaYFQqN7bu2oNGDZCzNPQcb92nkfZ97/BTzaK
29Wm4kH2ycKorACbYsea1tPVcgimfGoOiku6RnWaXwU/9loDvzP8cE7fg6n6wgOKwLRl8CakSvmq
8+7ib9rtiUmqiet99q6xY0BTofqN6pKJGH353w6NQ5Bs4Vxw2vh+5Aey/hiSvClW9wDCT3DBvFPY
yi3A2h12xYTWfXdM4ja/HY/kTxGxp2kCiGHat3BrnJvJ32gsa7M2EUxw0oohg5J95B/pvHFK92G1
P95fZ7y5k7VaTJ8PTsPu6MwR3DA27I7vMP/Ro6s6DXyUu05YAI9GCSXtufWMr8HTcAu0Wf9JfIxJ
QmKGaRnN5b6fMwV2u9XhSyMjFnr6nBomc73JIlYr6embiAE5Esyz833xBVKo5zWbcrehTwuqVLsj
2Albr/kuLsmpsoqgdyUtOmiuH/LUzzypJEVjT8sknJMgoW+leRTBroSK053SS0FWUPyWtxxBZDUx
yinzN6x2Nvwv7FijWOHrlj6+OGbJHgtecRF9W5pVNtAPi4wxvWZn/FoBsC6f6W5TU++ownbJjdtV
SKY8y38NAwj3WDVHlGyxLuR4QiTcq89FaplbbREaio6noNfpLqB9SGSpRlirdTVphsrJ3/STe2Lo
EF6xKlgpKTdDjPMUACqYHfadJW8PN5xDy+ykNxoW+879WKawUPU+cF4d9inK+RauvbcIdg1Xq8ZM
MW7IqSUJNWy4zOx1BMOUTHiiyCrBZx5lCTrJeuLKL2GeEFQVtXYPKuU+4tuhdeE/FcW7+NB6hkYh
KMQ/TSiVL6SeIpxUpDKyn7IRonxJu158yWBbuMD+86/TM8T5yuIdeb8Yk03u1HUM1S4pJa2NbMpc
5pxFcc0CzezZtbT//y1uCryKhtVmjwUHEZ72iu7mTmtneG0R+a84DCLZLUux+bi7KvN1qfVB3d5e
nCpBMhlvRiWJrzq0l5FAbnxzZ7VIqS8lQoZA3PqJ0HrzUmbXonCuKDcPsaB77Ly/+AHYPataH6s6
YW22yaVYl7/M/pShOlMr2slxWlxYmG5pX+xW8y4KgKUFR+icUENZ5yYNdnxFvLuecL9YcufBr4D5
bZwAfEfQ3aMrTP44imAiP0UIdI/xooSymAzvB7u14fnVRgZoGFFP5ojO8lyXM/CumOZ8f+1qyOBS
mclG6pTGtMLIfj5V64cZvr9ES1or2Iwwg4iZ1O8wJ/tSocT3HGwQvoWISSaVBIKbMkeANu0w98t4
y7YbNqZSPcJ1s9PNyLAv/G19lTDsh7pcwRPgu7saV+X/hnu5UgQSp8NTbaiigL56NQmCOFMTKBca
5zq+DFY/umMwNSDhdaYlzU/izZzev60tbTho1WP+4xabuk+EWwwgwn6f2FB/Yi7XBIFDHcpR7VI1
4IX3ghmrtRqXHZ5Rt2i4eBzr+lug4LbAfAkGOCvfsMzsqTSh5PdDS6l1PBqIBPhnnXsaN1DR4XX0
G4yUvSKFNUefyZxpmYsTL1ZxnGNTniQQBG6nDm6vqWEUfcbAD4VzxMfGBmrjOE5cCKX1P3BdYZR1
edSENYze56rcwvccoelY67GhefC1WVcJnbwQaioZIPOxp+eORR0pCdQCpJ0SYtp1Z6ABiCZJPsBr
/dFfJrtlPUq2+QUWjRf1h12og415aXso/fDt6nx51ki267Vdm/if97t44+dp7Q3Tu6d8yJ9+dEG7
dW6wJGog9lr6xRdvgDeLnQmgwP2AaElTpf5IwFAaeLJkFzPSmXNFIAYEqvSIT+9yCvhue3flUNx6
nCedzxr8p6arnsi+0Gjco5AuoeGjYL8MVTC0+EC/5BQHVw1cSviBZwGmDtjB65//oxpYa6st6yVw
GwDPjmZ8ewA9LGpgESWjRtnBxElt+x7jhmZ/38R2MdVwBkEk+/m1h+BRUWtphgiLsrKI12AFCYYL
dJ03b5fzaRpcnf7XAQNdoeeK3UASIrAjZe5iXFrPY0NamC6ZHHxBAcxhQm7pG0WY3yUCFmQUisTv
lyGwVwv30vWLV0hFnsyLQvW4+JrVDk6RRlMmAJlnEAr5xZYfVedOjPmq2oM/H65mYRdXGf4bvjby
7sCwCWICpUz8QgJjR0Qpl6+xQIRR0LzMKDUOseT2MIdmB41nSF0uMh1htGVYAaiyeXLa6vuG/Xmg
f1FMJ0jPFZZ6h06RV8xZRraEHYsqpVdRgtjECSZs/361EKGnqZJOHaXIUZ1CWe29JfaAlPZYEBaY
0Usy+cOFhMjsAK2JRVD7zdP8y2EVMzYGa6QxIUegM5a48GhQFTVKn9+QaQgrIzuKu9ZQ4eCrFaw1
/6XCKRRzpXBO6RcyVUklrrhszQE5MZOlCUE8BN5qRB61wffAeAtF8QtjPmF888Q6FM1DsoEdh9Ns
eEntO+Iiu3iJUoblIyDxrVppu4jfg8gRe6TMFVC9qEC8HUnxBLv80GzuNDPqsO2wgT7CdsrZR3GT
aM0t+kWwiB9svP74R2R/l+kzSXo2aZX3oBQ5s9RqPPAqdqlKzvAtAMpxeCdxZkLG2EJGh0ri9jHy
TNThqmWUZsf5R/dlh+o/sj6rctV5oqfzSzJS6Ds/wR+lkaVcloT48hfJwLZFepRCxgt3j7IWO1fh
hApVQ4k/caVMYh1YWtSOiYXQuVbLGH5PUWoJA9KTSSxVyZKLHTXPOUwyedGCpbmNlelFZtgSTn2q
zoqlDo+OGkxusUouzeWVUn7Kr+2dmwLt6yOLceTcCNdMpBNugMAE9FXLHZ2V+ge9sqdFFAcc1tDA
OzyNWZ8pShgumabYBTrtx4Obd0hCz7U+Z2gTDoRc/ZGxe1GQt+eCX4OYRWrr0+1u8xOL8tzmNRKU
wwWNQO8Hv7oEV4jtDNmIpbVtdG2wTkE5SF7nfwMsZ3vFFxcwG29d0I/g8NRto3IOZX7SsqKeRIVe
8+YbEkXBDyE2QYJLj7ZqyFhbscBcF4ltJeeSsLjQjfNOVsfTrCpr4Fi1x74YXRE68WmEJTa6F17p
QGlytSsqqphZQ5vlr2O6XYnFSze7WxvQnsCi9XNoFL9Ux52f3Y5yePHxOEZXImnn4FtvsPT+gF8j
PNkfK8cmueJqTdl48uAmp1YlgweEOXFG3IHy2c5uJuuYepsEJCLvZiCdwPVVvFLPxx9V2BVcd70U
h8lRbfQHN9+YOwjAXd6Jv30G6Cu510YSoYVY4IFPlFgNZ23YTJUGl6Z0nuE3zWfw1PfzBM3lcgDw
T/GWFdXBtD+rcPPbXwU+6KBGGubA/nLQG0CqgKJo40tSdcyzByNA+TWedXD57SMBQoepxNLqa9mf
b3k5nDTS2c5JY/TpWxbvn0TQo+2KxxNJEPn//mEnmu706jAp2MupGB06M35ggmCAd5I6T4KgSEC+
A8U06Moj8Z8BfQkk6OOUtef9UQcT+Fsz/Ayyk1cEWNPEUxUZsTYaolM2NIRtlOCg+yEdw0j6oyU2
AbYW1q40oq0Vqt1A/mvKjOg+aJliUfC/CZrwUbpw3vvibt+BetLxmNXS1PT/p5c0TJAHkdy4rYsU
Np1AL4BqJJCkQliI2Vzaz/0zSoENfl5wtUQgf9yeKOyy0zPdRF4taxSzqp4zpoEaQe9C7e6lExtI
IqMOWCFT3Q0ZdbNRRDW4MOX2kH+b8219C6YAhvV5xCIp1CHeeoux1oYqQ1UJaZgNqkaqVwUh31Kr
SEVnAm1Dz90acqo9D5AV5He2uOOPHVn9wT8VlUPqQIstNCLvvAg0nCisUz5C07oqQhStT2cTy9Su
YtMiuMdte8nHjRszRh8hnj5hl+CyC2vTaLcAUytmtSQZ8bOKzMHjrnRdVcAcZbOma8ICip6Y5BtC
BKzKkW/O+hd4dVD3LRx/9dYB0GYLC+YCRXKrAoUkTbjVF10fRtSJ7CS7QcPoE93YSf+Xn7WCRvbA
LsedrtUDFAC0P2lAdSWW5UbN3tj0ex8kE7ODn+u3jx2CW3xMtCI3qzymEC/suOnp9h2+Yjl9rpPu
wrALgBLPNqt2Jy5QQJjT2h3Jov5hpn7dsbjdfiGZBFL6Lv/pfe5Tq0X7qAP4vbqbkYwwP3mxTeLp
rJ8Xr0Z1sKGFPIO7RGCCbztlUeyGRto1YNmEnMK0ewY+EYIIACMkmiq8s8jTqUZpHjg+KVP8Ohpy
zne/diOcM/fu/7iyUnM0fGHGAr4+FrjWkPA0c89tI3rHTib1xV6Ro+uxPJrQiwh8eWOiTh3oXVAc
WWii349IDaeHzvJ3dBRmufYKTkgK328sBelrQdtVtmGdIJTSRih/aI9JqZPsOF17EqWBrn4zE6UA
cg7ljiPbpR7rKkEb4zYvaxXhLcANXDSYmczNAXLCtdn6ycT5d7RL8pdkyAu+R+C9SwGN9FkI1Rvu
rNWZwyJsXFUDE+TUjazg5pS9ByjmzlGrCoOZCkn0c7Oi65V/JzDN/16xi1mgXEzEVAYtpI+bxdaY
KWe+B9iOGbK5p+qORAnFLQtPfUTz9ClCmYjXme+JitbLBiTQBKetMkNar4Shbe9P/1gtlw+Zoutr
6tWdTNdQWIlCDxhofQ4wvlCedHda6+N4Vg4rbgeQoVmX5sCeyMAFFIh8oUWMT9up4JGvYUnIw+Wu
wXSqcp5NIgLyOioi5Vi0Wct6/VaL8+0eYwZpRsroFGm6ZC9ThHWDY0XMTt0ul8MZ3rdz36Lwtljf
d5xRBmYHDMYLFyAIeeBM46BnqXyuRWDzXhONzmtGCOMZtB4E4Zw/8PKCu/JVGvifnyaXR1jP7u86
i9GrzjWusu+2eT1U/xHoGB1PU41j21CGDqk9xProIRto4xBMkg1Bo8rqh7QHd/32oJe02h8eVQ1/
jSEM6ZW3n7/XqhN2CVnGkSQdv1ZIwAIfzC+Zkb+MAqM1YP9AqbzYsH7s+jVxoD/XJZLpYFnyyqcW
uMeV2O497ckeXHyQ2Z9J8t42ty+/yUVPQVVXlYJS0F5mwS3Zu3JYlnALGvfD2aHqqvYDZLUAz8jq
4b6O4joumA2G/DdSucSuxNqqYkMlZmaF+4Z/zhYNh6cZC6BN3EzV7Ij35wRy2+vgnI2dXpWU8X27
MImbYSMBCXM3SDNIoWOHU32pNomNx81P6T8FAbYyZ3WaJtDcv0XiTo5vt830jOBT7kSnsQDBDmME
4YFaQ1dOUTD5E78URXrrOZbDnYbadf/x3rGOBcByCmB94Ht0IhXNn2fY9JogLUmQ7i0Afqcjx/iD
FoDf+pmhu2t6DSQwYPt9TeGqRZ/mwEk2oFrs5cE5Idq2HRBwktFKXdLeaNc+In5X1AdcH0EjC0LZ
rEjnWbLdZm3ZHNIXAgfz1oR/tNkp8HC7mv1YU3gsZXxpnidtvlPqbkYbDYeeFl138AaLPJ/RlKsa
DaXTH4MVFHnE1J9GLXOmXNtGOs8Wof3FJCIWfBxrgqMo03UKtTgtzsH+RLpMGVRjN1YScgRotVq1
zreFA7/ARDgXoqFrN91iR93/p75FYPOFhV8CcNGI/r9tHNq1uKn5FPLrI8bEGtd+nUtcE3vHKPSt
RbpzSJ1aYHuVWU0Bwgt+fDflSjxaaKVvYh3EhXbyWsr/tCk7o2v+6hc4CEXlLEvnQm6bx/AuyurL
RbNrb5zTEL74itPy73NzAakM30Acd8GySTEeCspz0k45sIoZad5yxLJBybZP1O4H4GXYHFZpUpHD
R9uZk6a4fmY9aLycgCkrIVlLjHI0cYFEYvYpzljUNyZ0Y+D5Wknw6VO3swN1OvjchwuMbveiQy8H
I6++M0J+9toY0QQA6bwqcF0cZWjbB2/Lf5S1runHLyic2thSiQyrCE6FgRisIoZrEmhaweU7Z4IQ
NDB/agxfvZ6VtrRId6fr2j7NHllTan6BlDZLlnAUIpl3kU3XQ4Fh4xLbP2F04AtjWvyepoySf1oP
y/L3+N3wDFe/egCqIdSFvAAMC4AOgh35Lh8LB4YsvFfol3TcdwfEHiMVjl27AZy0maVW0XiUQ0zX
83lf2OEJcAL7VbypEonVczjKWK1R8m9xRlzOPoVcTufCtwdGZkljwo2WeH4o2ek+LFLkUONDkwzY
AeQaumxXN3PtvBZSyapJi18FMZpu8ZLNaYeZ51TrhBnfMuvORcuuim2hAlVsJOaVfEmEVAdlPByL
xIKSICsQwFhRDstwQzNoUe5zgChZ4tyHV1FmvNwF4dtLphbnm9r/e+i1RoAqhp9wbsRz5WzP3yDp
NTftIRimUS2XSxCEtPzmS7pUeh4vd1p3c2HjkXqCWFyExnMJPrUpt65h07zLp0ee2l9mRBQnRfDl
6ez4sb42QoKOTN57MzZ7iNDXO5QICRpV3cp39V6MibLGqtZsXxqvoAGZxxSX/KIO4bRZ2I9rimE5
K9eVyTp+H5NgIpOzJfq2glTnQGxkiZzXKRfdDMtbuGOyrPbvBpcZBHp1b+3JtcThwPcxlbTXIDFu
kB4hbYZDc3TKaB5EwSFNPcjFAoM4MTkeuedDv8ZOunEWOgic4p4azpIZX5cFT4UlBLd3SYtJBSmp
sqBf4JeTXsRq+6yUrN69uIFUNRjN/UcTCPMFBkFKtQKueAfO0l8ECN4epOApgsav73m5G2Wb9Fdk
G6iHp4J4XyfaVjgpajISjYPPNky4p7FyCz1cjtCSz8SujeD6gtg9BSPYDcXJpQ7eM2p6vk6KUTeV
pKyt6RFK/L37ZKIjYp1VVUxXArAW88flum3MEF93JSlyJM6IMdu9YEg46gTk1VxfM+VI546L/BS7
f1Rv9aotfMid1+5NacxVGEq0mMDbCWD2BdUy9MtY1xLxwN+HUD4NIRoMXXsHgAACvBmMTbexXT2S
V6NXJF60JpMDIOZErbVswdrIGkJrJXrpNK0/W3rA8KJMoswpUDu7L5xH4pKg8DlCKLY5KgAA3Kd5
KYH35fewdWt6j6bPFagwLdAkR3gUttwKoYvmVNJCjtd/PNafBPEPzckWXNJ/IkRYnBxv0lvoaTSR
zgKVD9uXk0aUhjv079iiy8Jlg89csKMQhKDOZ+mDTJUETxRtMh4uhVDgEVUopP28ipfRHszQZuGr
vBl3+4vzCT55izorbfxqEExD90dRamlIhHzeCUtlXxvauNhCBVam+XUDxwSlMgzgq6HIEzkajDcb
bIZdsZnRAQuK000jvs/Z3X1dwTNrX0+ru0n/Jbu7PZIGdKbH7uctPcqsgBN4THZi2sp2r6jsay0R
bjW2RElS+dCHagPTsjrsHtnuZofNfqxTgslF/EawqTMjcYDpZ5pV2/JJbpgmxM1fiZMzRSfOuWX3
2pluRIa5wzQA4ZZs55FpAeMxK46jO0KGuRPD+tb/CO0WfVcVukd6IrLShEuc2a4gKNxr6tagKGcx
2f6R3ebJPOjxgbqdsEkW4KD7xJqKqKbgK0V/T2VoLxvlcfMAYhI3NVnxWkkgYxVX5nr3+Z+w8Ivy
cTDaY/W6+zv+8kebeoTTo+5LkF0qpiSrCDm5Kc2REIT9j3Ottm8KZwlRMEdmu/pHFl95uljxdvlt
v0lm3sTCRk6VKUlr3zQEjr6xHKDiubD3H4tNbv4JBtdje1tGEqK0rafmt5zxz+d33SfCcVl8dxj3
Uz+sT+X7NADCK9yJMo4KuFxGdyJNkl9/58X9xPSFPGeMthnDJDXrj6cusOOzldUZLI9RfaWGjWN6
EELkFWboffxIm1phLrWW8xPCNIIfB5mx+SHME3kuDcDgihM0fn9iWSdRU0NqrNBZkRLQ7RQANe2W
7PVqAIAKVahwxyZI+pXiZyGRJP+rbCSBOBZW1JmcpOY6Lxv6DPomEQvTfvXqrfgSE0LwXhCah+d3
O2Y4E6jEf5gXmqLX93jZp19dSGfFvm+Pi4Fxvb/oE1Z6/RfyvIG7a4rSrVAf0XMwFdCuiv9hs6sR
UsA2tfUb0kiXu9f6c/J1IhyfY04FqlOfhvRIWOlvlHC7ur9wMNn2G6Ge36s8ESZQq6ASWBKtoH0H
hNc11/SbNEfHnCgtWlIJsCVGuzGOXzoM4utE0muSzZolGFX7PGitiiAJN3XCh009wSJXetw2ZMet
MFfUxCDiHKqPPOa8jiBcWYgKXQbNUy+pCBrQSPk5ZL0y1nQxyN9hbxEvd0xc2JwNrxang1/+4+y0
7Qt/MZvVuXkf5q+wg6Y3mhqbFQo+k6EoNOVbm0Eh4rsIUpp6zOWyC1293bumvBQ4JrVlkZ12SFS/
Po0qgnKcJjjVXDraO4p9HHKWySShd6FwqdC9NeDiOHSLyLUY2nUir0KiGG5LdyPxb3xatxFAivGe
gII5aXPXvtvOC2FB3/nQceHHpp6NY0z/VoKLG+r8nqRVXpsj0xkTnIB+9qPWZUAgSDG78jbWDns8
XBAJ6HMBnkSv5AspfXBneAjNAcztKMvunW+4K/GT/l+Gla9P/ZnyPAAoUOCMEs43u7d4+QpDaNOP
cSXT8s9EuxzhWIBPaShvPXabIwCOEm67QQfUeAVhyj7RkJ5XgiCBn/o4nyCdN0K2tBwB8XAhyeT4
YYwSR8j6Hoq08zszeAdbjUgyG0Sdnf479oG1fGT4c91BRuJuqrVcUaJvIsvg9YGOInq0vvqkIudd
m6efxoXfTtutXizbgwEUaOJqlQltif4naRK7S1Afd9HQHIqH4EXggrMqXOLmf4jQdme33eY6QHGN
NgBQxZWoONW0OoIt37x9wAcA9LE0Ollo00MmAzDtSyr0HndrPDRozMJfuXr9yECiJG76kMODr42u
tB4LoXhtgkmV8qnLwOR9TYViz4leqWHqE8okph2IHhiwCYJShj/wWyY2B9Y/6A5JxarAvKhK1GNB
FzhEDcqfDI6NdIA90lALUl5gPtOPXGN8m+J0iq3VTXVvpIv31zA04wkO81Ux7igSVIFB30bNM8sP
uLoIZwvJ/Hcnn/jKVGBIwqf5fljNSIN4Wef9oAmxslwMejpzcnqLl52/bJ/yH1zAcoPTOsr92bl2
l7wnJrUHPiZGaFFD/qMBmPgGz8GRotyWGQ1CLll5thZhLsqLwdeehHIL6HpBQpn2z7BOLRqg2kXW
eJW2K2p3EVGalfQ3wyb0K/uMHbfZrHn1Rp7zXilOcKz8pYUeHpivR9GkPgUpm/O7dMkOz8idJaae
LaYdgc1xtIh2CrFqkZUJATF0ODG0qOIxShd+ZplfEHGeyuc1Aylszrvc657iGuI1+HbPU0MaOBNv
31wtY0gnLVxl3SSbJRMU5o0AOZK+yEuXf6Adxz8eHq1xnQq9077rZO+krmotaIBQgTXYPQHYuL/Q
tkdJcv/eYPIxImhHaS3B6jU2myfJI9f0ScrSi6bE1DMYspJtgWwNtzJ9OqcCMKT49iNWdy52zM8g
ss6NwmjWegoWYrvRuRjLmBpA1NVWbHL5QQ1jEezF4KLtDLCi+e7AMQWMY/ldMMJV834jGcGqH4xx
NUGnq6X7sjnZL/yE/HRMU8IO38wU7wh9TfUmK+9feEigDiPAku+0DQMB84cWnA8yjpKEvuxbRCMa
2ctNLkiZPM0uxm5JGwiips+zmgb4RhIskfVFF5JePpR5B1j3B8AfkuboTVW8muZTCdGmKU4qk/ba
M04MeCvPv+PEM4h/EnW7XljZGa0nFWwq+Zh2STHM1K7HgcAgidcgPGeLNV5f61RJ60I9jWcBoXj2
1P+/ve0e8qdu+vSEFwTezDGQxPhmAV1ZFMQs6LFnQVu4nAq7mU0BTTdlgp9QjqLbhkBR1U+lxIcy
jA3TzN4D6sf2YWYOQOcceDRx7PqVfiCFY3ehbQ031YLLZwMqSF3Qb7N3ObLWHvpMBHrLHewD/qPH
ASxtdQu13dWe8zWnAOmCLtzkpk4iIGF8+/pwr+7ipSc1Oyqfzsht2A3xMyRnzmg/KcRF63D33RL8
vftL/6s9D/NwSi9PjURQ0inVCgFn9he40RCHjXEFadRgGs5B4gHHiwuDq2RSJy2X88B3ZFTnj4vX
o4RWY4FSwxwwfEt+kiT+s1GFSMJiLEWE1H7ytd4UDe7ScVR5fcFTxCmfJne0iBF+uM2bXNt/IzMn
SNZQW0bicEiO93fPbn4sXc4yNDW/eE/07bsbc42+prUSOppd70Rj14c0xpzAwfyapHuqGdT5Jw8x
ODDODIVY7oERh0EyUikuvfwJfLOsUQCigdhMEUlKN7YthaxC9gvXuo/LRyZMAqHlTYo1r+Myrwj6
J91Wc91dAlGxK5isZsorpvBnRjtXYVx+rr8iP0eP9ufd85J7EfTZtgKES23L9hGpkKAxIJRe0Q/p
4K8nNB+RoXy8uwWX0j9j7TbkiizRAAx41Vu211bCd2SXW8Yw8Q6sJ4a/palvMYkQWl+wy+3eRmvU
55nAlQzL+Rn1oJf6IFjFfAFtLHe0Q6zGr3/4IkH/b4V1U1ZYN9BLOo1pafooNuHXIO1Wgh8fLl/4
s72abh/4riHlHL4G97xiqBCp80noVnWvDQEAgTCjF9mpu3hOQLsoi0A70/5qYTzwjce0HVlqqRkO
ClRYn4nbsXsP3xsQT/zpEnO9BQZ+lfuH+8fjqo1vg3k3asL4hY6UMQ7t/aquD3nTR9fJ5jvj3twy
Qpkoj4vfBa64BcyokxpwVijxN160QMM4EXbR/NTNEj/4gwnWeKdu2jxRuk7fAdPd0JKvx5OCwp41
Kf29uF7ISapdSRFZFxuNY2fc8F8F/v7UjNRkbMsbwn59elksiuE18GGfJ30tY5CO0JnCLXABSttj
ubZPSBiQoglK7QEC8JZ7vix/anT3wBFL+b1zasG1I954+sJGRhyNpOL9KrbhXMA4p1Iq53NMQCCJ
36M7a73/BjphreHIhJvUTXUt6cVl/I4z8G3EjU/CfRnCFK7qiot44Nah7AlerbTpw+hPJbJlmfJu
dL6cS1sq+fUO2LJKds2drn7wIE6qbvaxSkHMJAsWVX2TILxDALu64ggxlCzOUpij98sACBnTV8XA
kIKydaqiknOkujCptEgz1aA/gOeVIpp2SYftYTNbp+qjqtLOZOyOTsTzewTqw5jWnHzSeGMwurYZ
PNQGOq4YWoAxVUecURp9A5d8AHTrST0nFr4PcEgav4fSArbYytHycw7B/8oJPLNGu7kaVeIiWLlW
mFTuFXx1kZ/pS4BVVXWrSO2l9OW8H20crPZ3+OBPGqONj2K3NM2QECgf2ts0vLwHW7g4Qrpd+QXs
NZi4ojf9Lz2jrh1d/w4BXKw2noS/pnW44vDMfP/5sCdkK5V45tRjgGbOfXJQ5W3p/xk/IMXNowN/
4numYCAqzFD4IjVZe7zaYDB2Jwc5fIRiif3vUcpydXqzfO8eOldT58XRzdVnQFa4nwyNsdz4NEuN
jsJJE9SLsLwVIm2589GYRQviwXzhy8gKbfm2XWv3VOT6hmnCpzr/dkySAKmk0oBzsRekfvO50FbA
zMYKf+E3cJp/rX8/6y6aaaCGWk/avi0zFdd3lJCWroOCMjqQgt0iEAIaIsYctNEDHf+GYWvIPF7o
63XIfE02AU13gqxbA0BlP6hz4WBqnn7IgeM/COSuaRXbrCaJOkwQWSwdq0VyiEAm96A+R8MV7eVC
eZSIhCTcAic1pNGGr+7Y3LfB58J0ARYr1YexlXzmepaGfxaxiTL6kdxLI/2e+9pWKQP8R3P4KTcM
NofIULYZ6KeksVVYQ6Nclh/cCb9uru2ArFQViGTamBEtHkZm7qITCstJnG7m8ryrJI0wfKGKKamK
Ac9h3K78FdJs1sVOnVHm6N1yoyZRRoNYeTPu01QAYnZRk/wY1pTdYHVr7tfa4D8AKTC5+dnTQ0Cz
KBe5++a+1x7zPtnCC3ZwzgKxKoGIKu6SpvK8AXn+n2qXRIXHjjCIUGltiMvVwQpZadH7aLP0g/Zx
irTmMR+mSGVFWmBXRhs1NEXPyhaWrFK8LNXFAoLh5GvlyL7MHvqCbWvFH7lMhTv8ILi7RoECP5UE
zpdjH7AtLpTh12/7yL5WvYCsDQedJunl8W4RPtG7KKnRER6YmfyrgqhwA7X/o9xNFzxOJWu/rY8D
gnECGFuf6VBkR7j3aFsYN5RzkPKC6+3zZMRUg0+FGtMxmJmwVmUt6XSfX3o/ua1qdfSvRFt7IQXG
ksU92xua3HK4K/w8RjGFPl190JXtqO49BbkbbuGnbqYQMfadaDz2LqwY+Pk9fyFUBhNnH56DXLht
2yfdzbZuYAX6cC6pWYXZewM96ZEw57Aci30sg6lK5Qu8fXm4AlgsK41RBr1uPZVNJ6NNsmQp3fPR
vHgPb+QBKx7wHs8erE2T4uiVqISPqdnpIIVEgBDVSgadW54rhyq5SVL2gHYdkartW8BNRqhVE2gR
pVk1PLc3EAMCbrljdYf3Gg6BUyF3bJi8K3jT9VA16FtbuuF5DEaZqKQU8733sFjBdvLeZqUST7An
dJiTUYN8ye8WlcJ9QExTUuEUOE9AydDy5SuCGbb6Ndb3knmm6SbjYS1TZsyeMCWCljM1P5XIcgDm
GCJaLLk90BQSLHcQfxyHZl9HC+9GooUUcveHDlW0QTh5ra7AwSxDWHEVI+g+XwoGR1oiwyaKfttS
BPH4WM3or19DjBdDPTZQnpF1GpQ4sS/uw9WfhGXqXvd4IynOST8/NLZ0QjVFw7iy2+0Rg28oN8rk
YqzQ5GoUhUyLURZGaWSrCMNH5MXHrtV9nmi9Pm90Z3MHbh5KIjH1CBnORb18tUoMVV/0wlUOoKOH
kVC9QVAr7zlyLJ8Pm0fQo+orPP4tbkiLqSj7pJExF7B3la4hOlvgvkKH9ZQaOqMK8Jsncqkx0IgO
B4dx8E3ghkT28fcVW7YSsF0NbXRENElRQfTesGEDjXf023OEz1t9KHvRZprb7OvLZNje+IGfC6TS
kNwYzaAOi/k5buP/2fz78+GQ8f96z8/jCo8r0Aic2KM4uvk0dzWZdpJUct4uMj4CaHmh1J45JuCm
yOfsjbP6fVWoqojMNkd+LfTP3B0Rlevs2BZfyKu7TdXnogNuNUsk7f9CKyLEM2U7BB2mWbt2o94w
2qGyAqzAZhpj/bGjCz8Plj5T3AjiW5iknBFc3xOJsMHkHxy9FiNnxXZxtkrOZbWRZnsHhtRXYBaO
YZIGbnqOaFEe6h5JyMzdGIJdtc4bIEOOVjyavSNzOiv8vWYeP91LOsxYA6RuctMel1g4+p2NKlP4
NWcWyGVv9Sur0PUNeFmNrS8Du87gyMvolUOBW1xU9NKIORV4gkw46zvKwNe4noc6x5tXCdmP7uc4
N97nC5I3tYf8LIakx88/2Mf1UoyS3XvXaunPKPg7fZb1FbqUq9SUr3ob3kaNtfuISuMshTBMsSG6
Ctxj9/4bnuOoJyHibmcP2ze6tDTUgq8B2jGI3m3JlCRBIlAxiPQfmqX1TUoSee6FPMYf1gUSYUSU
yYlwE4o4iFLQ7cdR5OAXu9UoUcYwVH+csbO7uYbk3b5CFyGeIgiqaJn+re04Ni6Xec5fJGO8LqGT
VtfP4ZHDumK/6nAidNgGRhahXlZ6dQUA8/tLrnuqxn5Y1HW+fIxd/wNVsEBhz8o4SsvvfSMaG3m0
iTaD9DK/lvvPBBw5C/3XCiS7DHaop4KS7CAEUIMOeuuC47yRJw+t2RuzenfQ6CRqzzBMjYz455pj
9nggSd06h5ZRvny3NYrcG00xbt6E4h0xKq8GZktgW8aQMZgOmDEpjPVrjYf34MkQTjVSUrUH8O6u
bNUU2tzOT6aQbysm3WWYkcy4mKdcKAKd/Ay5DZMX0iyV7RPYg+9sKxNMFc1kXTDvryrel7SgT2iJ
ocwanMVMWoEHYtjoXJW6kv8cH/3kdJL4dXfpAI01zSCKS8KT0Q0Q+BtJD2jb0qH+KlYyXSFstiLa
LWeoDKNmeLPoilZLoBgATSeCs8viXzxGXizHuH28K4QSHc96Xzp2bnK3X7dZ08f5Wlx9OlEQZlkb
4fVcpBLTwE5+m9O8CyFZ405eYC3Rwo/nfAMjF76v1BmsZJycpaLnwOujmw/gSI+6kBVkdyuyINJU
ZdIY4w4cHNkTe5ctgshGapaga+ht2+niY1gHYsfYaujPyFFRtLgLeB9BF1rDQWf+aXIypFjz5/9b
eaobgsrBeq4sg6kBisV9dlE7Oox3WizP9m+hCci5EkEQjXz/Stb/7mCtwWWsF5ZdC+ye2zVk3t/5
W/Olq5bLo04rnbXkmJhXjSsDY20FV/HEYd1ScwnoGgZOCFJh+Y4mwXWK28J/cwXakEiYgWTdTTsP
0L6SqAdH7R7IDNeCuDE7wr/K8iF7q9JGE0HYhzCnNQ/H5kEqMlfa6vUNDQxoq4Hn4DGUNXRs5MRz
fJBAzZwP9PLli+/EEoJJukgkB0g1iyIFPVFe7Cy6+3bMVCPMuG/1rFBYDenRTUQw2Mn0+aNNb9Y2
IqbDTGJBu0EwA6RwKABCMyXpM/jJU51noyRJ3dE1Q0NH4gdvBkzu/mKnFFpioKOKY+I1yp10rjQe
6tFQWjhehrO8DifB7VOcMkl/TqpI96HmOxUN3XzJ43f/oOYUiu0sw763K/lYxINmhGJJ5ghVKRoX
NfiuU/QBugpKrCzCIijI6lufVUXwpquIji6rdRur2kQiagOZl2lj2p/P22CbDkyR2vFW0B8+sdNZ
H06imugGQ3M9L/KPl2woK1iIQsYIjhwtE9TL0GwuxvWH73HtvpsNFhZLN4TnQk1Sh4+RvZFQNoqq
dCRZsP6aBZ17E1744Lh1MC0LqrAyiqqxtX25C03WGxV/RbCbgbXnzPVWJpW3WFeqrSWrnIzelChl
cw9G03OfYOnjMSv9OTgjiU7D9BR135m6Lux4MhyEmrDPRFnhKDuXCfapU0YKBE7cXfQctIG32gVx
dixrw4+Or8KsaOonxfREtZhqpslCtk9WUPjhh++0WXrJAkZ/z7TUrJqak8xLFB8VvACNgrZgIKJr
FTxLv51O5ju4T7FAjO5fElkwwIex6yc7J2ype7aGHR4lwOJxmEz5Q6c45ieDXnIBV2gThBUMuctK
jboKNrtG0YLEq5gIW1L3hCmp0AmcBoMXRIuQ+vhyB/IoudXaMQsUboVE7sgPFfHeQuKxTdw8PRIp
Du34PYAg2U7aaWB6NXu1lg3co2Y9di9xuil1z/Z7kHlXytzkYE3ss8rypTo1tUQ8h0gyDJLOXdHi
I4lQH1gn8/l8S62nNm9juqQfM9Acv63TB3Zj4w9R9D7HRUNhxV7CnoiLxbBHAKKYAae/VuMR6uqL
WI4Rm6GvvpAF8IhyyA8D/UMigkZoBSmpvAGBmYOFa1QeD7yateBexTMKXMnOWFELC/pFWrdtvJuv
yNEK5f8Q7dj4PtjAYXCTj1gbIf3+jcvEUQMtS3MK29hHRf66o/AlX9w+IW0RUeN9UTEEr8apCHEX
Q+VaFzxnCSxidPJEpBooMTbjGpvCZUw7IEddsE7fbXxI+K00oUetEYdYv8ij6nA08i6yhWCH/EPu
QXUh78pj8h51+7ZD3nzms4wQz9F36RBTldMf62KvKkwxAeh9wxf34yGWGcIbi7rCRv+Cl6jiI99L
g/u6yXw5AL77ErnEw1JtmUqwngR/u1P0rKZDUmz6J9OhsW3RmPtDqh91BoG0MU3s8SqIQx5W0IPI
ejHCY3mz0m0nir7yGJB7kkBPe56gOMRICOuIm6RFPqCNwo1420pWnyP4sqVo+0uNU+eHwDIzzfYk
HM5BhK/w9I6UjQXKm6e9MBLJNd+AHol5oOvTnnM4I4w1h6rmd07d71JU04otjqPn9ssIMJImcEdQ
EcWXjqDz0TvB8Q4s1UFFIvVq8Ik8JzX2oEV6VHM+7yo4/GomSJFJsls31MKUREjCURDCSdxX6T8D
6ehJK2RisZEqjyDBstnWl8VwObyjtsgJbW91zTQB6Ym8MgB8kKcKD9JiNIpj+BjqDYfZqpEzXbrM
R+RHbVB30/4XVqEmH4hi83IadrmD3bzfqoQpgyen7Q+T8X6N8OzrYrQtwWtp8HgdsMxGbV26MvJR
6gh2rn59b5zHHhPu0IKzzeM1cL/ki9AoYdvd8hnBKY+TDeP07STj8tCJCzcjOYj0gt1KHb4MHg7h
0qVWNupaOMH62+DBJFmJToYIE9WjA8PUKFWDXOSKKQ953IVI70Q+wZ7pT7/+SKv+0FKgPBMbCH1V
VxGc4HTrGN0W1vN6TJ3hNnL02ow+JGtQH7FKpCoVzHHjTIkGlYFGkGZnrhWHOfArnZAsRFmnQ9JB
wDeJNyVCBkETL4i1kdJNGhEw4apWJG4nojdXz4+oscJYoEd+jni4WceAqRnOCRCQ+TgyTouPpQ6O
qvjZMMvE6hpFJUH6mMcedVx4Fyz4pLsYJWTSfriSvtt5cqyuKQJy0lCTHZyp9hyCXpFGSe+fuS6v
m3WwavM2ijRYo4nQXJwlk/QdrZQahLI3SIt8ZYBYE/+ZoMLkWwqcByltzDIRgS2+eUc4xwYdTE/y
NoIFz4hIOMLm0lRFiJElM7X8KE5Ryi9enfG0JPW5nNuV2AtPa8tbTnbPksdhUmRvBABp0HgIIEdt
C26bN2uNdbmW8VwTESSBapxIbe8WzC1fW/ciqDFkgSMc2Ei/LnKPVOj5DckJY0dZG3LfwamXhI91
PZGJxHSC9/HvWVx8jFYHKRWVdthZRel3IWI+v4Csnx8YKHRWn8etLvcZivyNS/E92QmbCdo6s761
OCYIp65cFhOyG9pj0/yc38NjUPboJSy5yckop1GMAIoAmEfNOPfMlq2rCncubPDt3lWtobL0+SDy
EvUc1o1mSnKqn2RTToeIUWsUgBB5mRM5HVfY7vDHCY4nh/tFakHznZ4Ti/EBPgD3tnSdmllRfPU/
zFm2FuZptyDnLEjBBFoI+1C8626qzzDqK36R/48MLM3NN5H/l2BHSmF9RdlnsgZrgl+Bkks0T6lu
cD4O5/IeqPZTQAUOe53s1F+u06HfRnfxIC5F4M1/b/1zQjsRYNK1FNR0X+XgEZOn/0voXQ49277x
+qaOvQTdSZ+uuphYrLAefJ6cwAz5xwX+zKSDg8Roqa4tz91yGe8nkcHHwPpGpv0IsX6OP8VJqpaf
w54rha5xXP3VpbezK0ifuc4RXFhWg/yFWli1GFKuijEuDUZnxvvXwFx2PNzOZAAVB8yxOVOTVOR5
zb1dgg4YhmLPDQmZPBO9kZLOkb6Ck84tq6NHzMGkFDUmF87dbUnyjJIDdBA02FmBVChgvWxCjTq3
qti6fLcticOaD77UjjMq4wpm1+Isb60EMLKRJ1YLdIHCPJ63xGeUMxFYi3iAyEmeqSniC2WfWEQP
y+YbzITX4p44wgtzmZ1xyXDjQDEiiwao8cCdXIlhOKhznSizzwovjdt7IPPTnZGrUQtbvqaw42w0
ro565irY4vmOT8akmV701Q2RVF/VeFY60N+0EiMMgk5AzDCVt6VEBbyRXPELHiaAByiGmjqoTn66
2f2LijUtJDiNH1VXNT4wqfV97l0JPI6tim3e8GFgj1wCFp7+SYR1t6WuE0mnP0A0h7OsBPixPH9n
wSRvQ2L6U4DnIotMH3ffw2HRcZ/x08sC++D18zXAiq8BFjcRXeshtwNM9Z41+oulqBlyyaU8wTql
0SR4oPZjDKX4EP1HvOpqRmkmzVOMUPlx1dwuuXLFYCvfVp0ZY9ZsafkwSP34KsOcGbzFdQDz05f7
QPThDd6lCgCMLpAxGlcAucLlAmOD40Wo2qpXnL8iN0RzvsP9WrB5yQl0UxXS9VOfy8vw0lcLcVoK
1o2Xyqpsim44VfXniOZgPnwAVESZMG55OZc8H9Rc94IZvfIGgCnQ9X6LRlJT9emyKatAKDM8ZOHg
yZeOTdL7zWXj3l9Ey1duvHi3zCCNW6WCDKihnOL9gAu6bLufSjDe9srHtVp0Vm4a9ucV0s+GqtpN
W5r6LL4rLw9Ex0CA1xDAHMBuV1bjEtzGyecyhArDTeGn2CRZLNXKXU7m+Djc6vus+HZvgisJpwaL
k54AXfAFLXdJsD6Hb4mYxV+uulflaRbG8bap7IISlXYNf9PmbvGfMoKWvcpUWFwEE8JBpFeFX5nY
lS5Og/+70tRNJBMj1muLPa0RdnYl9ftRhmsrllQuv6nsDFz9tSYExzrdhaJZONsY6IOrpe6YdoZw
XhKqxIdFmE4LczxFEQJgObOhfJOk4CFtSlhajuIY4YY3Qz2EwvDithGQ+ERe4cNbiedVKGpOYvJN
8tZhnYWcN5oxiNXgrgReWH8a3kxPJ7zMoUtFzMFiDqcvOOIUSWJZsWWyPvo/+lLyoEfIOR0OtAif
OlUIgCWJ0wKtzXH/2tCkplRAjPQ7vwx+m8Bs78+HEOxEAbLPhF1fpYEs8mfglH76yAjh0Re+WyBr
AfuyVbyxdH1CtzVeR7ckOC6NtXcDWHh8AqHtJkDA5v8K5VdY/9VSZXHEGHyClBXZG5iYno0MtKoJ
ocsJ9uA5tJHRBr4HcsWCDnnv9/BMOhpVxfwWq9huwQe0z32RnjryCuOCa/KQCd/SfdUxTsE+DJny
H8iLjTa+NMTLIsoB2glTyAsEq5W0MX4kLQ+N4yJUOgjoUb6AbkSuZuLTu/t88lbbHp7eXmIgmkCb
F2V/Kz6/m01IG/7yR2hHCzGfH5jh1cNICtSLGneJJAXU8aBApxb0OVFb5SvQG/ctau6z45/jdjIu
Ya79HO4lfFpDaU25fKpS6+kcFVY75IY+7YCULRdnNbWDTfVPmPnsi5/mD+8dSd7FDXRbtX362FUj
xP3R18Mxf1RNlmvfdn2BomFf8Cs6pg3F6oW4jtq4UnZBx+/T9UD+TMTWQ9rafOZPU7Na1fvOV/Rk
zqx8/p1X0b30mJa13Y5Y6TSDctF2M1Dj3tcHgDI0DSC6cA7YV4ela6b50ABEBcYs7I09+N1/GBvS
eQyxz0/QJBwxFcO9JSYxuXCSP4lzRMGgzG4ZI2XnL5oMcx5a8cVEpBB8x7lQYuhvzaTmC3jGnb0E
UEM93iKOO1DMiPhnuSa+BQrr8IC1Z5Hm4zbW+YIZNsDpe07wUyuREadbRpRAjF4HqFmRaWJ+F2Hr
HvljsE47/LkUBz17lLP5nFpnJX9wcj4NlpAeGSabpvZ/zQ6o0nIx5/00ix0Drk2zJYKOuZnWWOjl
DGfJWLe6e/A9deftAwda0dxnIhoWukkKhjUxNL09+yC1Btwp6rt1u0IZc8R2iGj6gYQCJcMhbTJX
y/9Id7w77dUlpKeTym9oiP9cJMvxTxuclCJm+mABmPJz8Fln4cEQC13NJM3YFFQeTw2aJs3SV8nA
3lvbX97Kejl9gxd2w5KPOfobq/oxAsxh3u8RiwG8kYYOx6nyxnehczHlBikUjIkL/Yb1RQZUPlWL
ZmxICkNbNcdLvs6API+ufVWFYrcjJ78SMcukJlFSgSmcMGmoe/0qlngewDnCDZ87Y02rnG8cNUpz
bMaX4jmBFqtiGVXaeuvraEMIQEM2hGN2j+Fw3S0p4WJYyXcfJpchxdwiBlYPRGSOtUsKP/gpdFu+
jLJXsKbPFOmgx83CyVLf610khglZVAKu68vSFd4dTAqKvdx9PhwcEMqdPTBxZFVnM+MJNSlw4idj
OyJdnEn3jhwLNTPPII6xQLOUWpqGcvZUvYRiuHpPpSZPPNf74jxFBKuOxSEAkdRvsqPb4q7qdNfz
xxoB35fsfQcLTW+gDxE1MIFObCXCGIjVvDHkiTc5+A2zwA6s5N+UQzL+3j5b0BILzDMKhIPyHqgd
zqwf9E1LvIiwjfgaPsViru9/Zwxeuzy2jsosbuG7FO/g97x8SO+HXEsuFWW9F7Ynr+bxUv4je0oC
hIYmG/YUWdHV2YTiCMZJUPsqkvF0SAJglCsm5kT7LAQPkINiWjATgfXsrqVVOUh0sBYHaVtfRq+m
DueSs9yvJTArZGiHtcpoxnJfpMbaCn33rivqVT7lSAzo+8uF3RnmCTypFRON/W6wvEWFbfqjRYHC
XAVWQH96uABWrr5a+eeKFz/hD0w12Lw4cs9KkyxAuMf9moAV1iqCMqeCvJfuf++TR7CkOmPWA9rb
C/GkHgiXwAy68ybvprSi0GkyaV2PltTKrj4w1pM4wIGXj3E14/2HT4uN+jyzRKQ3yFlG6a2Kt163
N6Zg9bHl52Eo1lMgwn5vC5+JiNSUZYWsPXZxlZhbutbovgYN07TLmSA204yY/7q4AePFXK7Ce0sk
bicsnsA0Va9VbZnkdU/a10BKGPqUhG/+BTywO8DqZFjiHd0ZaLuxHkdQksrTL4TtLa0zGW/TVZuH
duL4PjctCj0u9Qmo99bANST1kkhmTd0WIPohUXrVvxQOyGKEON0utoik819sjOXu6FSA+oGcJUgG
+J3GBsbKxbuZyWWkRLdu9aCel14cNW32metUmd/m5Us7aqf8qs6/KclY4fjIA2uOtBRtcKjVISNA
C5O1WWpotdWPRx+oQhbywYzeszEnjGTSctgq+FuI3La2rzbfHB+ETSO4XMXy2TawWT2mE/uTw0Vy
0PdVD6OkJz2MpHTYISqWhF8sg9al84pB9NRocV+J3wNL07D70Wdi8APTMtPmdz7suwncz19Szleu
Nr8ervxe+PWVterh/RVjQVFfLr1/4jp3R+9g8KQyMAjLDhUGg4vKYo+nDjLaIyJmImqn94L1A2Bv
97e5xv1EGMW9BfbiAwmbXfW8V7Yd17CVQeMmo3HqTXUFOJjbI6w2yukcOr4SZ/UsB8NXH0rnGRC4
gwK5CAruCli2nBoGIHNI+8quxSBONrMh1811i1cIjH+PEINB86jC6OYbUWiNMwsttAgd3/yAfBLJ
lOa4FqVooqS3uaz3SHY5Bgykk3viT7oOpPjmL8oMqIMQ9DwLwb3iLf2X1s0aX7RcaU8Ret7EsMF2
7wVM4fCl2SkLUZF0Rarkp/RLbrnEiiqSAug9/mqd0lXaYLIGUBniF8r3S7jNtNzCxxOa95FuigMs
E2eFmfmyWCfASjGOXJDOq6t1urG4C9yi28xO71ihviriENWTW/p4VaJq3NMhaJdtQpz3ZB/XgnEs
H/M9QtJyjRBNVP2l3joC/rHOpsbd004QcXS3X7Gxcl3YQtF0sK+dxjUjDSfMNNDAnWccbG5RIYku
9sI9kAiCJtlaq+bVsU9N9/4Pv+QKF7agfuA/62SVLjZa2yJn1b5iCaEQhS3p9dL0R1hhwSlRkzw8
VDZklWPb6Hk3liqAyY2OqH9xhIoNWScYrnWKPAxJ8xZbQrm8vy4nI0ejVzLIxdtWpUIygTEVJ0dW
FzwnxeLyKZXVvBCEYJDtQlV7EgJNTJlbfbZSuyz8PS9XVKhrAFDlysuYr9wC0SVLSPKEQTUDcnbM
UD8piuHP+QrbSA5rFdeUZoUUN28T5iZoUqE/zx7iktubHJw/KXAyFsz2/uxoKqWvbUzoXYor/2rs
+mOnSGwVlsjZsF5eeDISEqYxtd08F1mvqpcgi63KJPgq7ff45IvWc8NW8Nt9N2PaXpOBkd9L7nSD
272jCqNGWo6gRxFsUo5Am2MlzS9ei3Gf7ScjPrmT33pK4hbw91b+SlAk3oJ9IGwz47nIjEpFTUw0
v4Ru7CG2tIIe1oqQ8vyJosus1p0/94/fSS9Lgm6k2ygqqZ5L/9zr7fpQbFdJuu9vuAdOCxjUmzu2
8lxiLBRN3C4ZyOaSK7eqM9+qYWrzwkrkh1CddZ/yQDMEgHvxE+E4Sac3Yqlj/FVztDyRoS+GoMjs
auf0XzPva5y6gU/8wFyTl6Na8nVsG2juIq5itplZ7tdqt77NvlJfTYTi+P9Fn0W1wsbQbqQuAcHw
XtoldWwTQbiSP2RNBELnS/l0Al5WRkitxfvGf2O8cBf7TSlUpWe3gAzHOn74MNev0qepUB83sd6D
/6pRPfT5z6FaERoUSzTPnzv0SZIK7dBHYSYrcPXQeEjvHvBg4PfPkgWbCUJ10J+THPG02wW0eGHs
Z8YNzGnuV2jsXUvu+vgX0IRt997tYoIRekKRRYejlkxqrzE7NZ1Jgc8wypHOI5abol3vTxGaAqWa
FLuTWr9iTJ447eZpeHQuvwOmMm1sToOnlGxVpz+3gQ5LhqORC8Vznpr6q3Gfbs1t/KUT5uEE6jqx
sPfeSmwOj4x4ccU+TqO6KfH6r1iO0+kLPoExv82rkfsGa3sQX6gvkXGAO4yvk0MMyl3ZP92gZF52
tq8JbMysl5jsH9PJAaey6fWu+boTpIpQs/eCswf0jOalJhB5T/FZcyUTrdW39yogYksLuyoX5Bdd
5EGJvnludG+rh7FiZl0Wb++RAjAB5ayB256EhDzURo1fsRWAkQgVBQfcTtVvc+4QHlxn3T7sjZcF
TEg2lk4+QjQcZTxcwzS0J0CBGdR9HZTd3NBky61LDWCXz/mgPYgPfsgOPSSHkaIIaNU2NDtexZKS
TTdDxlB/O1NEZNSwxsaRQkg5E+VhbP8wTiIB+yQHaYKu83FSgIRx1PKIFWxzl98X1A1IQdFuZSVy
rpSTr2s2PTzUW/0T+dWGk+jltOopfiOtfiQHxb2g50m4vWf06corIjW0ea2Yk38Sy4Sm350fXjwf
znvTFjW1h2qO4JCWgLPKSmkK/LUs+QUiBEaqWGK3BdgsYqfkWWQaXQ5IR0IC2DTh6LdptbY4M64w
XPTMUKU2xEFtzEDntuPpSwtcFQBrU5WfBmH7Wrh3r4RtGsF8iBc0ywRy7I4BAZCGJ0hhm4YwA7b3
r4PgVpUlTaE8CuHP8E3nHNW30fLMfTW4+lmHAyWpFLUV2O6Wpvde+9IZfiIYwPzz5zhHtBCxg3xw
PbektaLrtxsj7zfHuPeHj4sFJmLR16Wd+niS49mg/lPUdO1ZU06yF757azRA5f+YSsT6ugmnpwZH
2uRc3v3GPshDvAP3iS+eqghdxoalifAHeELiJ/BaXRVuA9xbFbvBsYVsC2E3JZQpEzhVrXKsyxSr
qYpd+A0TeMmgITUF640PhjUOGeRREjaCBzVReP5Ql2bw2degUutf3gQO45cqE2Lbfpeb2BTIwzCD
7KCx8I5ZGXucEMcsRSm1Uqtsm+qrL+33yELAIxc9YOQXeiM7sPBZbo9xYGHbc67tNbKrnptOrpXz
NfXbbcmY3BV+svrVwAkSncEbqZUTeWGMDkq8heM3q7DpHqY/1D8H1f7pXQqBURhRwfh954upL7x3
CdSSxP5secdr4EzmmaF8wNd4ECzgIuQ37+9cMPRqSpQrphvfWBbml52V6smT9kPFKlj6Aagn47Dj
A4bgTMbfaRXwcEVqeGjIl9h1ue/kDfg/YKSXF5Vm8uAkmUZw5OLxGkLndDZNFaPHModlIQ7PYTTj
4MEoKCLOksqNL2AjNtGNI5WJrrVNZ3VIjVlyfWQrBlY+55A25WjncVYbKe/9dliYlxNbk/Bys4g2
EFYUyPcOyxtD6gCo9m89JSLttcROsXYytmdpUaPcYjJDxZkx5lJrGlYGPw6mUNd6qTkCz7qAehK5
2XeTM1EfTwOqXYzFDJuCgY7kmf9WLzQZ1XazduaaRWX1zYtsb4FrOruAdVMThPstypDysMfZHb2u
tC3rpzdpJYOrD+6qxKImQ7sLYivC0ZOhn4fvAAzOF2ABTGa5iQBGeANuSHduKEKyQXvlgZJ4+3Cc
yZ8hxtnxpXM34cB7lLYUsErmrFnBcrcgvHIB8FvFugq0WgEQSuTBJEKm6VFL1Y+wfU7V1YukeOra
sAUBeCCRnZWaHPJjJXJFJpacUmi42JKvKyYu0TOYQ+Tvy/pvNCCkXs906HATruY3h1YftZ5qNc1J
4w288+BFH2yvhwp6QNaKBgacgCZdN7+ueiLaGrEivB0ksKmSx1bh9bn5YLibjbnUQ6I/XwpjEOlJ
mnGH4eOl7rkwjNPotIqDl4aRQdh3wS4djsUSBHcZYmKPEFXhGYlkd5I95T4Ky/s8ZgskwFgm5FCI
ZD4Nd9xXPSmt6o+Osdd6N6v6oKvXO40oLqsH48R0SeYOcyJXNnwO/StHEJAmRWVM1c+bO7fVs3lZ
kdwrFe+3Uoxb3lHLDvzWye+iWY7dEFxRDxa/FtHyURia1mU+k0yY+bBueQTK4F1xOLP/mAWgMXjR
cul0TElfdHVsA8fjyhHlCq1s+3c5AsSGKdZsZO88tcEWw84rC1oTV+iaGG9kkNJMHv8JpOYHQdg3
rBATsdkx8DbzRA1dWvX3KvsJfeY4cujM7qFY7HVw8k81q4bV3LjYjXfVLmEY2wNN75WGNlcYEO2s
KIkv2txQUXcCiMuzGXybqA9YTPUdjf2NBV3Q6nVizkS1WIj8kG2vVZP7Ns+qh13XzJ8IHkVWvWcW
B+FHj8livYGXGHihXJ9WYU1gbeeeUdlhUOVex1Eaby/r+CynuBviqwhdtfKMqHyPEDgpxpui7uMk
unTWCDxoyA8idxmsuHrmqQXJ3SPrcNFs73O0bIv7Z9AVoC8Uw9eK+6XmNXeT9/kOZjQyi4mUAcj1
xd9GTB7oEjVGgwx12a3TK0KoMm7FSAGA3OupgiY8ASNAEB7HdfkAFgT+oVp5SYo71sVWqYbkBkHY
YYJu6QoFw9C41N6k91pbdFEpSxDeYBXbiCzx/5lL2v+evSTjPIpGzkV0nMe8Pz93TUqjbDQGW5nO
zwh9FxJJytbD+YuFZcEn6B7HbxsZT1bhZZay7c0aesC3qyWCYTtqXFUqvga9f2ykJcwvzEekLwhC
oMno2ColLqhOgakP+TbOjFG4xs1oB6iduA7mbamWPaP1IQ/g85CGSIGdzEDSn8kcEw6YD2psyxR2
sPPOdKELfSGVtvEt/zHUc5JbDNpKFTW7jdh+MnIAybALH9077RqXp3cV3fLG+cD7mUOq6jeHffl4
a7pQX94o6g6slMF68QOKaJhTt2h3YOTY61k3IzZtS/htuOYl0M9+kvlfU6WdNyC3WScObg/x3wlL
btlGLIiRA2v9WX4rRj0GdR2XauPu/6zDe4SsXgRgITA+wADg/3b7zKKEQ9YGL+/+elB7Rhm8UEDJ
COI8qEtNeZvqkT9zlYbqZUfRMQZAAAlOG3slEt9SYPo6BdX8B7+krrR+Xo/BoPKp79xc5Ly+8y7b
QCCX7crX97J8UyPP3s/6mvDjzeK8FdSJdbpasBPxT/SqRkXp7xgEwa/eDqWREmD883xTQX1MeTdI
UKORGk0aXIAgT/Kk/NH9NpoNsoDBo01UvtJlxB7gh4QH8KVU9GghFoc3VVwe7+j7P/jB7LlLCf6s
2CX0M9tyPtfarQTDW6NDGZWQrDapFqtDCKgreNwRUJ3YJen0XGvp8RKRMXIkEWSvPgC8F5yeNRyK
xc88bhz35JgJs/n4JcOnyRmP8pjcsoWH19DVICKpvWkJULSNsKgeJeqCN4AMADung5aqj98vTYVS
64mckN8hZiJJLvv2JMz23fDGh2ooiNUec8pXR2rqS3XGlYKQfj5qnq7ApSR/z2X06i5FfFpg+bm5
Nc73s9cs982y1Tt4ohM0VrfN15E4G5AoWJIN6ilB8SbMuk/ss4MNb/ZRj9FyduVQQHrYKH2L8GLP
PpeJofnS2yaO20/lI00koUz3O+Tt4sXgJUAEjIskz4wkKLfHkPL6kqUjdf8C9uXtDWuwU5B2rhKL
uyL7Ez+s9oLIXQRtScfkUZtOQuMY3h+tqX+ecG1wA1WskFoxBhpsob488YG95x58Kc6PjJ4hc7JG
wDlbg8v1cHlj68b+AIbLZKBddxoGZGT0q3VEte5yFfLMYA0fC16l40iqqwpM3CASuE8FUp8imMcU
ocIoxXnb/LIoi6PHOl0JLajM2j4/Ykbeoz42Te5S3KQ4SE4RtH/T1WMApH0Ejpcdaq/imWObM2Tr
ze/7TxkI8zzMSGkKPgBprQwslsiVeJfknCGiw66eS8lKOSqOYxVBOU/Iyz6iioqj82EY04dbVKKm
U3LAKYpJ47yp9QHMQwAJBSj/K4GbbQ9zbDqPsprN+TOF9f7FPh4ISxOIeJoDqpPB8Is79vAFwn9n
uh2YaSAtBxQuNcHsYyFeogw2S5KSNa/anvBB7RKaqTW/Om6FS9jQ86TYZeu9Rl3dM4B1qZrz1xlE
BsTDYhOFP94yoIfe5Enhq43NokOFT4OxflqX1AHAli90xS9hDjpjVEe2lRTmlJ6a7gjZSjhnuxtV
V7HvSBmQW9cG4Hr5O6t/Q0XOrTjN6gRbMLAqNjkJL7aJDQrH6147IyR2f6WEl0AOBTIQ78FBfDph
32ohVHpDyk8CofXmEcaqHPmRPyHSpUntTBAu43O0PTPrJ7T3XLIUZhvldkDUwsWnv6PNE/QXnqfE
sEBPxZvcYU3As1FqJd21cIiONHoPZWwKFpvSY/AZvy+y8+5JdkkBZt7uOvK2I0WaD8srQJ3SmgaU
CVZbaNr94oNLq1shMsGn6geDThj+85My/2+KCKlB0YxeXF1/C/VkTsj8G7x1XS7r8Pz6ob0TZlyc
IvpPRuHeqt1jdIOYj+o6ThXspYkdnrFP16oFj8JT8X1ihnR3lEnnEEQmnkLwyXly4yY3sYFBt82U
W3o8/3Xradl9DmOoXDG78BBcyJCgrxT7h2kx3AYWap6WZXOJLDsw8aQxp2dew8GGMC1hIA6Erp3Y
gzzIX0qojMwIA2NJAD3z3nbOFf6Wc+UsBICZ8yXsvJezBoJLwzHdM5gk/umJt7tF+ThHxKkGnlgl
zDXsWZXi38Ze7IaXNwcKeqoUr1p9Z0LDAGtwg3Z5TMd8qGRMhTzDIdhLV4FwoT3knwZrFkIaufUW
Ux78MbAaO1/TuE5LDfNWpI8iZqZzhwpPnKl3ydRM4wZTqASiQzJ31z3hAwcriSzBKerLHnyne3Zz
n8ShIgOxO9CWqE5V8P2OaLWsqtS5kKuS+ZjAAqAwO106VSZJafMHLbFuzChRPDPlCUNW2FWMq0K2
6T0F+XQkZXI9v1MmrOx6oSonDG2jvjgsQMNGufxJYp6PIYpivwwqkH2SONr8HMhdWp0fsK6aDgfY
OYFSNGLeXWWo0a4A+YHlNXWHyCcIiSePmWhPohxrAMgtsCrQsFqPRn5eGfFSF/pCR/Col3rL1ZEv
hCQbKzXFrITsXbqd9gwJYzuiSIUMZ2uVaEy0+bSaqRXdz5inmoKZyuUoR1JlZX1uIRqpJgIbLydO
Y4X2EzkPhyDLGEz8tJMR+Ye6wfP6sKOGRT/WH4nOztrEUHniW5MvQdrN/XviEauipkiuMF9uhqWn
oBWeg1Qb+0gEwExgXep5ninTKkKmPQgj4KKtZAuVpYZ65sobgK2hlN22//MbtENSmIrYBFXkeV71
/eZYOBta+ebINdeWhRbWF3DksNz/phISd3RPyZf36Msls5UGGd77woAWPAlfv+mgibQEsK5E+8Zt
d+fzODksg6JU06t46RloPuSidKoxJ4TtbdkVRLbBTX/R5dKpTRdeTXzaUKubIaa6yriWazWMKqYo
lawaCiRnPw0LG2jh3dv4+eQhYckZLaV9qBiI0nEKITzp8u7p07vnTmZZMtUWGQWB03GbnLseBwLM
q4kOSarvgHnYfy0DaQL3AccZwJiCWR/xkK6NgY4ayVTSrg+GPXn+YAXiRUusTeFIz14Z3kLc40vY
4LXAbLlvgZCu4K6/OwUkZiUxQrZL5KEWWsFwiQtovNUkOSVU/H95VcYIrDN4vKnsuLq7LajRzpC4
wQvo3qh98mdF3SdMumwBtGjlRG+zjRaDqceLqhJLAXlUOqXj5HMh8UAwgJMzCrmrayLxKDoe4CKU
9Ke3taxpPHwaCg4DORmDgrXm7wbyZ+TROOAS5o0+vlKdj2SjsrxUCCDIMIb8yzg7NXZrWC4+eJct
f4X2kUGVShD3gxTDqYvKbGCEdZwNtI9UsJHtNGSe1AB45uDeD6Cl4xD1mo3zR9Ph5dbEwgXKKAnW
5qY4z0bcR0tV+I77QekK1EQY4TsRrmnljCwS0uEyE4tu9LTUhaBF2qVvF/lNDjChbb1okbvaLvTl
8025Mh0ObIVvL3qyOXyCDdJXmU61xFeNhJzBSYUyoqyaEWninpKqsCIgHZ3W8BMnl31aXGqYX/0p
TFmI0IpDR75aGT/vL6g1kFk1W9FaEKl6o4WOXzFQ8DES67hOwAQliEEo34jp5DNIZzzf34hfhJ48
DGp2vZ64SqVCzibUs66bKoEHOuy6XZ7jFLO1hX8RjT1BdWyPAXi2LDiwHGesfz8COq0JYolc4HHQ
gvJnxIc4e+Lth/nbbWZePbdS/IkF/FqE7D2Nvb+YYzEKKDScwRAe3VKDUY84ypzQrl3SFVPQDDbO
L2vw/BIts2pBGqwjBuFeFVO+7potUoZnJtHDXuLuDzHxEsS4UEpGRFW9dopLb42OqMylzQNQkv2w
mWC5APdOhYgs5lGNjNbPjGeQmu9HM849KiDQlb+BdUXyoeNmzAC2/7fYBQETgB/iF4W+wRaZQ5Yu
UuMU3vEUQYpzeJVYSJjpIeT0Gw8S9Cz0hMYIgWBVRjVJ/VAlNvcEw7Rgft3p1YwAHl5tkvOKli6/
SJR96Qm8M3fP7LZZwrzTRRmONw5bnA6uxF2HHL5edvfBkVtA4cTbVY8WSYkoIyILFMmt5onOQBG6
eilavTxOTY/KllplQD6nKln7Ska0sEiyGfjlPPMcKf0Py6tlpjszfvSNGMt1j/4mYyoM2c3Eq4mS
0mVI8qeEaHQt6jmWSQEIQDJsGmYmA5GkNYreYkb9GWJVhPHZrNZ9issJroeCelAyU3vOIopWZDwR
EEhtRs2K8sJ04bD0KlEUUS54FTX/tBlrBqBmOz/6JmgcJ2LupqwycY1BZLvnsLN2oxHhksHmROaa
+b8ge/65SwUU5QICXAVVDdryhuLBrFv6T3FiwE5TjIXKC3VjfneeYn/by/1/MPXFJnP15o0iVsIG
geyx3oJ5tCgww3BQUilAR27Be6ECfN16Sv21EXi8Kl5sTKIHycwGWaYb8WzztkwRCuQjfglRY5Rd
iGLPhWkBM1FUMxAWBoz6+HtXusJSbs6Io138BSJSYhM/PAesR7rY180Gl+//LEhmwxtpnOHP6JoO
KQ1X/7Bpzazyp+7Y1E20MAkk+xx9EJyaBXU3VGlkYeNYk1G1mnpZu+qaBl//te/TH0mNiqMQUpAH
AvbyeqeDnHJHFSdjHb5mg3bBza6wgMCQ0h6xPQxpdPMV3CWsExOdHJkSbz7b1VZuAQvGpIJqPtWP
WSSf3KDP+WF8gEIfY40JxD7/lwPpRAmzit/i1cUzXtAQVCX1HhlslZyuZOorba0CtYGQ47C9rR11
+gIyxMdxzDZZgKDQbFhTdEKLphtCM9SGsAY7VDWlax7swjGekTc3HuvwxwaaOCUJvG0FAGNdFREx
2h0UKo5ATgi8r9IZilLQXu0t++AFKGwNvq7/J+/zV04MrxgFWnNv6o+bcLnhOV4LxC77h6Ow91E8
kSF6nlXUQ19TWegb5HhK82XlZEAGkZh2TJoECDktlhoAadQVMWdtbe/scmj9mIhmJ6Q7wefDgenl
hxihd5PgnbrjVqwSS5zuPgZ0LGF8dQsoYJ1efgcNTrxpslS17VhJZE5v3268QBKrHzzSwAyKLCeN
3W8PfFoaWYpapsK6J990fzmwwErxd8xjVOgWB0Ov2cCY4AS2UV3pEmeBjXV7EhphSKerV6t9f0lo
1HVQtud5+ZFnBWqmIT79PLZ5v6g4fX6YSqSEGojrq5SIguWtSjCZmBjzBxnExKnl+w1Idky69uk7
7kgb0CGft48NkCJ6aZ+KJ6kJOjFReuQY6h2NfRDyjbrFZftusNkFxzWFo3c6p9WCYIVnuNKqPuv4
LeqdXbez4UgyWy5VKRs7Gda86mZn5nQRV1PEy3DLSGrr9HUjWrAub5eqlYkUK8EDCbc5y7rj9Zs/
tFhpCyHeLdY86Y26Bjr3un6bHGcUwqtupxHRFgCYoe4jGawxGdkrgghkWF0QSrMDN5lD6AUHUeWx
NN403a+gGbBarAYwdF9GE/GmK+BMmamTa4szGVEVzQrwty8fZvaK+0FPnmZBIDWN5ZAoCXtDH2yk
/Y2rvfjIR5IuqLcMuTlv42W6/MzlTxkdtPniOZJPDMLuWfHVP8yKM6bNIcjJgT8ZDkaG1wUCZEfh
0tuay8E72xlaC2IjTI3TylV2V+EJ/xAwcbuPqCO5oF/DGZJCe98tg+0Xzzn+ldqWFntL8GAR+I+K
MzzE/+TxhndrvLzfWR7oLNjIQELnukQJt+Ay0uk334O7XIzruKmnXBxgme7ccZcoH3TcHEGcWBs9
NewncVlhENvWLHV7areycVWWzvPgjkHCRXD8xKcmTTixWzr+f0j8LowyPXN0WxDABwgg1vU6nDss
OBx0vaax6mtToAxEuPVklvspfNhdXrU6PgXTriWYH0q9PxW2qtS/ps1cPVCE1dio2zSC1XzyrsMV
+AqISYIWFxHWU7NMw1G7Lyf6B57UsKgCvA1jFpjAalnhfIATEGkH2ETpq7D6TeFPFvH+MuBfxamt
Dp87eCWNDcuIIad6Hz4dnTYbDh3Tp/E83GmZGz4LeqBum4wIKzDe4aJSo2Ok+/cb84c9nLy9cB0c
SJ5I1Di5WM5+4wU5U730t1C1rjgH6cZQgaj/McAG880cezejNFnUCycXYzk6XAxSLRhrSTlPS/RC
NnKEtFH1emykmNcC0PkVK/ffjrFqJk76Nkl79VDVHhllJOmg2+pOGrLnhtInaS8AMbGb2nvnjSqh
DBHiEY6FMfLRzZGwDgJkZ92akZQwuI33dcDJ2pmoupUh0PxO5c5yYhZe+Dmi53rwjMlRn6XvEcoj
R+bdUslQTl7XbrEvhLnRM55wBlx9R4/ZmgNLpW1YuzwvCOQx1dg/E1KU2xRsduBql0FqYEYoLg8e
Tdy1L+9ZuHegXgdRwnbcqUqeYCGdF/f8D/g9eagv4MAffW9p10AmddYqbXthy3FlgThdTBgDaHMP
0/38CTMSZZRF8BnUaMKxCPrNAhhyBNHfF9m0CmZTNdKdWmsHW1BjjDgOF7wk1zXjVZ6/QLRD4Kuu
3vOBo0D3cOK1whn3y3NgVZWXwZophwOiPoVQSU2MLhjL/i061wJn1rn6+B3+AKB3Myn1eQuTlDi2
7m14gIlZ5j4pu22L/gijXjyCgcpkE6Hj/sBMXf9tYFRWXBVdgnL2CfC2/hfYI6xovMrY7TAe4YM7
s4IwOa9un2BgmBD4gd4eug0KKXZOqG96gIE8LG9K9sWDjxNvKoqPkRqgru1v6mvcgyUnyMhe+q73
8paTlAJMh6BI+GjfIVJIDgqPPd0IhLdhTX+MMENvFt048s+TrEMZ++0T0cq0rVEDXw0chDyuJE0i
4B5P3fiuG/CfkycYgWGsW8SphRslrHg75HfK7PFfZSmsJ3svTu7YqXIc5Qgfpz+MaS67clPy+tzd
hvluXOBhDQ5qul4hIqaK1GzTL6n73jYjMQvs4wQORupFTN/5U3BNvuAsYhFrrR676bd0j9DkQ75m
2IV8YIWcqDYMlkKCtLHUSOrM63d9GyvjIakiuBgtvRHrmXeahYxOrdUMh3ncSQwsculfzLMHRDDQ
G1oSecSlUaRSjnCAl2zWOL14PoU48TW9qffMabC4ya9Ig4IX4IQ1H2TdK3maov7bHgvKBqhPSbfx
qVW37JMAht9ulqIaqvHojEyBNAFn1WaQP7LPhDWkYFEFDCC5BRUK5wfsAEdZVkfQZrNtcqcYEoud
3SgpppIhUKhuPSIbWMyfAuLqPd8U+lXKKHOgObt7OKPuzKCxdchClU5jOZ65R3W7hda+Ii6cMUtN
NPwl0jEMGL6Ziq/yTiy6+tkByOuY/gOkT0ZWUOxn5gTjtbfdM4e/8f0ZarZOfLGWg0eLd3wT701y
f3ojNwJ1k68ZhfccKpmklaosziWWbLLO0uN+TiGqi8b8lsLWQfiQIQtOFaG2ygN8+gPoa9Ej2vHO
Hsq6nDdueaWk2LTdxyU/pad338Q/cxAEoXAGSEa3QpfgBH+yIEBoROgYKYkGJRF6i8d7hIegWwy5
ZrX+UejAP97/TKI6MKYiLDWLiVUTV8+W+L1Poi7p1nVBAtmBo/Jl1TrnJGKE5Q0NoDLxpCfExtOp
YcOwxe7jXTn4YJQ6V9j7x9wa6t+e2y35nA+RwjNfBkeedxXoRbU4DEeM6rtQ472FXViHPe9G4h0j
mkCg+1k5Y2WtAzQ7ioWf8fRMaNjaRvCCqu7ghahRy4i6z9tYHDuyi8WiXS5GrGZNlnQrSS8LezzU
9sWH4YaEzO/8WePCC1WVFqRcTxX0//m7/g1fJpzZTBEk06+3uS/L5AjFzSvgdSvN34BVASA8RzSp
DXrQMruL9FjK5fPdSWiSbF2swkU6oz/y6RmApQ8N2q7YIs5VGsU6y66fX6LHJYtHfW6l5mn0Vsj2
jZMjK7poQBDswqcmxdDy2EpApHJZUluTytWxdVruRx5AjZYeuQmqhjIUOtYB1ao6Ac2aPLBKkCZS
jFNHQo+zQV6cCyrRmlSItrvj3axSvV1XmCQeY3IT6JBJwSdCp2Rqh7wZ0SqLKIsf7MvNHy4AHFTM
qGBNT8fy9mPZWYAKeTaWAP5cuQlfk1Cqj1PFwj2NO0lA8RXSVeUlXMmfqBuaX0LYcsH54SeQcQ2t
v7xBBMPyJjr22gSVnIbzMZdVvfLcHVdFsblY2YKCcEf22baKjtI1iKeMQZSWIj259nYoSUZdHK2d
L2x0aLI+xi9GiWLR54g885P62r54ra+gZAWaWRfrJ/6TShPAXrtdT0Klb9na96/2uVkMcVg02Snd
RMRXOMcREJQMpgFfnqnAVoePK/wyMWUnPAoYFC1EUmjLXiLypxkomztVLVgyYgP4m12ungKHxy1h
31ejU5AZ51lNjovUH820hPvTPzaEJNbXPSwLg5AvxzNRO8xQJYtodC1U8YdkxjwgtdkZVWOdR/eg
F7ERho7FHEp1uFqNZDxW6Bq4W946dbi0JvS8wQaWrulRits7GQ2ts1wjZNMLflI4OpsXHaWBpVfB
rQWiYwxkQcJvmjY7SDaawAdWm0wg55mio2+uywutBlR6Yz8DhwXBPtBWkpjLYbHmoSOTk6OnUyFu
yBDb98PAiSiATWS3c9Rk7LEkZn8ORgiS3TVO9NTtB9x2SMdAlYvzKdwSlqSPGqMYLV3p8qT4mCu+
Qs0vQESbxfV0jPQYVsjgYx/XCFXlzeZiNxL++5i2QBR6FXXc5pI9zKrMDeWaCx3eOjl1xzo/4Kip
JVk11SaIPZX3Ejq0j6K2LrZSY3jyqY1P2Ghoyzo9wzs7+/v2TNyUhGCCcxDpI0aKHTaHtUXze6Nb
vB5eocyOU0YCrrnYEHYZowlV0QJ8zNZpJ5jmslSjaRdi7wj2WG5+CazGfJZWRRBkU14UuRQErCdE
eHo6s1i6qBnwg8sOSJsAW9tjBWhxOmEMA7BVS8y6lhqQtAk/mngCbJR38OV/+3GcO+Xg5GN2sMdM
QsQaEtEO0cwIy/bbNrUAmg1naYWbJsPJCjI10Od/aWbrPb3JkWd4M+NNDFVL0bej2gmHH9Y3YeLn
031szm6QqC/39qOsCQoU951UcfV94NthplwlVhf8f2aGK7R6ra+ZRr3ygrGoGyqbN5CaR9MxChJL
0U0BajMi+PIadbK45Vd+0Meu6DIyRWaoyTkincY3QPs8Ymog4Pq9nobVxQh+NeE0nL4Ns9YCoiLZ
OOVFf+LHBy4dEdqJId4u7fbB8YAJ1fpIa3wI2Q9NbuEJVr+HpSwjmZscCRjDD1L4AKUIlTfxxHxg
aU5ukVgFRALPmUw9qhlT16f7ncsHdSFsM/HthpfPYdVREB/qf5/+0BSTDp/NqssMiaSDdXhBaJSG
vADEoFA+Keri4EAAda/MR9asBut3pDWNrTcl6CjpFaD9RhtNAC1ruLp8lu2yHXqwW7AtbkCB20N2
Go0iuPlMFoW5rfT0Aa4Sz3xuyBUFDLXOTjzlKuMFsYGi94nu4L0SLgDSNr5rfqa3W/QOROARyctb
wV2Sw5F6nWRiyzj/R+IoK3idRPU/VQdP89jrV0sPm1Q/q6sZbNhFDDvuvlJyWY4k3BNA5vOo399h
7DqFVL9q77IbBup1kV8ufU29233mxfWtLu7eTe4Icb9mTO+6jn0N/7+8sPWSjM++XPSgXrJBFZfV
SZuzXvXcEA4c5rAOC0FYAE+LL0yXkYoxe7WIBpz9yhV+k5418Ewlj6i+hpXZg5sw3GE9okRlfsi7
R6RXKYnFKQtRvMvrmqmofCNSzTQZj3fnWgxZLLqaTQJ6wFftZWEJUrtZ+m9MUyp2CazE5lDZgsxp
Wcs7EtO8ZsszqxS7K4nN3X9NJoxavgnfODNd5qihjiLKaegybUHgSReHWXXWah2E+ISndZlYwLjQ
rj/7uiaUpmJNA+adhP2AHf5hND91Yw5acUZs6lsk7n77kPM9jDrGhp7Ku8lPcmpgpBR8oC3uFHPt
grTy1abXqMtC0/i4bDCyrIyxAZbDEONWbL1nZ+kRdSKi3Z6WXhcqQao5djqaoTZ3wX0YFxHAgfzZ
SRuhb6R1mzX3DIZlblwKWF3v2rSA/MW9e6GLzQh4ETEljoht7bu9DSZhqHxkWpk95nN7gq0nW1h+
Gc2IHDvdCocsb3Wkbt3tTSqeot8XxwkuOtxm5e69iUZGQk5ueXQnh1+zJpoA1/jrlCC1hLD5meJb
aQlp9l7gt3zEXuBCtS81XD9YAufHi5ItCYXNctceX/GlvBvNrNsDtDzZWILa4C8Ej6//PGYi5n+G
VpXtPuvKf6ylrBxc0+yqEleAQ1w7KVgIkLpbSwN2QE7F0JeQHJ4m7WK+TPe+fOa5ZZavHBWl7xGW
IQI+GmdrWoD4KDQDC6XLlvzFzN41yj4jTj/jQ/g8l+1v/5NsunSE9SKKs61asCp3ACmxkaX75dee
tRs4xDJg40/e8eAbdd3QLwmd+oQ/K0BkbYltYMFBW8uErAOucOHjRQEGs7S8wszQxFgoGxWk28kI
dXZFrXlzbVUr+kmW08obj8i69NYQ+lZiDdngdiNLHOGBg2Cnas/mW5VkoVYkqlUM+VG4inuOuw2P
AqbiSYAAoCtnrgz2o30ZfqAK5Mo5asF+vtc31XjKkmBjHIGmQKFotp/4s3b7WAlIJNWGoXjGGS6O
XffE3MuGr0U/OmaSPWmxEl9cpZO2VeDRQWzML1JQaeNFcKDD28ePeUCvTnNOpgwwwg0Cv6YoZ9qH
E9wD+ujEVxrg0M/WGiTj2EqVSAlcRrSpaNfdE0y+eq2F18KYQxNm9P8GCuJgTS/HQYdX9A0W4mXk
RBtXD+BHtx8oW8aPLJZlib2jpbDeg/0hG1zLGqA4yfKYwmx4HrY9pEe1keRv39ZPLzwKSDcF996a
N/jctvJ/mnDIokfURR1ob+CW7Z03/gtUZFSaocOPGyefnGme8ASghYrlKECLq0p/sTEzjXXJt2yj
FxD9bo5VEH9AuYFJW5wcGRv0+QC83DKCV9v0xm/wGTAfBIhH9++AmNS9PHVISHEK6WqdIShyhNr1
eoAmTjIS67y/qsGCLZbpG8ojk0xrCItZl+oGVl63zxtTIlaQHfWqbVydjcKK2sd0lGR3ap90+c5m
2V2Twt3ozGmZkiec5Ygx5MKWuypD3AgaX9w0yyUxLWoPwVW4GLoB8ZkrmG3uaz5QZUt91iE3wQ1k
AjaiDEmDLC/9jNTzPNrq+JxLwUIxpHmVsX+nFC1Hlr9M0F3f0sgZ0wVwTE1hYexHrTNcRzDGBpD9
TnEET00d3Q++xpBDLlvwxbEBoIC94kRS01y2j/aRAEJUtKDDvoeCnTv1UyuONS8kR/OKTQpiyi70
8yy6evk3ZWftF3hb7De/XtXDl5HUe34BDiIYJPeT7bLzqlcoOp8YrQapMrnn3m139OKDei7jZdsX
8Czu2YaHfFcULhLbw3xsChjVWXCV6wVcuf5pDFtcnDebioGVWdf5pRvVfHM90flaOkGv1Y/nQCp/
hObw3Mk02RjcuhsUAvoGuXgp9QFtGpNcm6DA/MunyfO7EA2fE6x4guS8jFXzAIhK/j8v7wmmA4EC
OOr/JMl8lD06u5meUzLtfcW+iman6VofCjbgCgJ1QC8sr2mhD8oHqz7KHBYcB7poyw6C5MTf4Q8Q
GOfWwwe0AIL5uP0ujyYiJe8oM/JNGgDIjy6vxfzff7VfJHRvOPDZmX052v9i/GaYTyhAprcxqaiT
LuHyQ5SrTq0yse4xhPCbfKRfayZAHQqyEAp1LM2bUcLwf8Wa4FjYjZ2QOWuMazVtgGE6RXlSunQE
54ZWLL/X3oPboNYeT3DgfzgSKdH0AaBJDZ/ffvr6UbhM+7OrrOJ2T6La5Yn5PrqdV1IWOIMoDxmB
pal8bRuOnilqG882HECOum5iczGqfGhsakOICEpVpBpMe3TBWZnkAxJ789nfS+pTWatYeqkQsTPp
K3OKDRohDt+Ff3Rn/kpjtb542O/sumgtCueHuDAFQVZDquVih0D8tjyTYZ0QdDla6z8OpWem8y8E
EyUcQAViz/TR46/yTk6gXQu+h8qlVcGZdcTxvACfgWMpN+pwn/iYDK0/Ha3TsE7wFBeIfOjP53Ns
0ZX+xHUYgjMrK4fC/2lHC+T16YxyQgqqcg+CraZx3eWtZKmaY/TX/+rK8NjmngVBj0bS9RHUZLxp
AJlg7geBJ1VfUl3mgHr+NjVUTZwJRbh2yq4Yq8ARNTy4dtkZD2+u1Irwn4IyevDtJkhjXzKNefwK
CXebNKnI4y7ezcYeDbtHCxekZqIuEUgDUN2MjRMZ8acPxy+Hw0vKIHlETGkneiNR1pNyXb2NNeie
NFvRTlA3HTa3r0t60ilehp2WLRAuMDepFRVMyqWc2UI2Z18tQ/Qj1+gc6Me6WAKJkqBjfLyCT4uT
zeXBDk8oQ7z5+qYWZKHzf66kpDO/mNcKXTDXTfFZ03ZnYDA61tnSDj5aoD6K8sgNuYtGkd8k92fU
y8T++fwM6CAEQFlX+ijvf/QcG/L/1t1d3UlVnMSVhp7BB7PAQ1TqdiTwMvX6dDf7XE87cZpnmBga
vRvl4HvH7q6Nol2u+HJNN2ZH5c2ZZ/3pOy1dDyYBMpbdsuHkxuOoiwHYyvkBfecJihlaoruJPYFf
u0A4+MNNVyhsCqQAVSkHwID3wrzOR+gumR9WJoyT+JiXT0LZYn7673wUXRJt2ltBmVytkHOifjml
CQYNsOVWm8YOgSXfAFb74J5dXHV/MNQbwBCLYr1MglzzOWi2ZHF5m8BMPA1ToRlwOe8WwMuDomMK
g8lE1VKyHBD9saU6gvycCljc4lvbhB8VcoumvQBBmOvVBtZ35ss6Prdv5HyOGDvi4lUSSGYn7+e5
0kl562T1q87bxHg7RriFOaOn4IiG+rhws2f0KUy/xCOwyGUqjxN1JuXpjcMlo+DqEBq+GaM5qGEO
BJ26Xw3shk65UYey0Q3YmAzSeB8nD+AY3dEpwi7+urBBDFVHgy88a0hR5Bucb8OmrCVpOs+T5ctC
+wKgy1LvEq+XqFJTy/xl40O2yhPm29CBcPoCWmm4zD4Nd5uykfQvZ07qv4LYGJ+bO93d6fugG6HZ
FoVeIsZl5g+hcnKY1qRj91/GDyDqlKMAPSD22EpoT7FlbDBklT5/TGRIinn3kefqywro9WiLz5d8
7AUbNtSNj68CmtcZNlJ0BJ8cBFYPPlSBr2AmdNJ4CvE2hfHoVazu9f7pxGhBVzKJQUQ1eMirzyeY
TnwGmGQfxEc/loIjzC5SI7YVhjeazdYgNqcOwHdJPAiM81XwIxzd0M4SPa6+0UPS/t1P58s5c18k
17aDxv7Nq7YQcSUmAHBTl/cle843aKzTfMoGZSUnUmz7hA3rKCd5ws5RQxR64xVih8jKOaluoWxY
/imRORL4gWUgqgpr7pbXanwL5IdvRfiiClb3+7cxp+iqzhoVerLnxaoV/9nn6OY2rMUDU/NVoOIq
1D/gTNZqQEIVQivqC7L1VHFZysWlHRTEEOx3rLmnQZDRq6ijNCnWpH8Cu/l7+fDZuLJdJAqYHpOw
bwZDQSHQROE10pMcLjRFxu5omZPNbME/PGgAY3CJoo7SzeD5Pby+uOwwI+sTy6V21yzG4WMVZUON
3S80VRbCuZcoh6sGaF2VPgM7BQsLMECkGeP9jb/BfPx1RwkkJfNt/DYrE7Yscc88o2DQFixhRrro
kfxsYEP84wSQ4WMrk4xpRKwc3h+6HrfRdORbZ9+/jDOcb3x/J/s9wyt4GlHOumBIpku6rnyar6PR
AE2Yh1NulBthK3GCmAu8bBIUc7exHGpegj+63a9V8SSwBDJJxxTk/U2oydraRFOi55JF48cXU9by
CouZN469nK3b54S1iJyWfL+z95e6fv4+OuF2Jk3D0P4aASh3hfUHvqzmlPu55Vv6FYUyR9bqM08R
Z81YMQBabZzqJ5O4bb6ZaJCPlk/WsfAEwA2sSpNDDDE21EKBMFTYNcrx/rETL9dc87RsGNWdblMk
hzAUy5xNxsvlKc0cJbYkGNmBUPYN/p8CsocSxVhhd+W6LzLLK2nO2PUVQ5Bean28+bTb11yilC1i
9sZLUO8BIev0czOgLyotUqUDFSO3qQkeVtZ0KbrI7QCy2QTwhLSLQJufrNyvEcDMsh68q6R+Meh1
OUAGUqCzOn2X0qc0DdPFVX3JWfekrKmzDV4/BtAthEufCL/wvku7g9SeYJBOqtjovBsy+KqkPg3y
aJ2JK00Bsy9Kdo3RhSnSToMbJjhA5kXbLvAe1QnWLkSu8BhV70By5AnbtztG07prPEoyJ/vEUQJf
ckJOGMMuQk9FWsrLdtDaI3X/ksHGYI2/sObVHK483MzaBYCfYGSx2BbzfNroUe8jaaJRMkdnavZK
5VQ4fRw0oZDNBpEinylyCUAgen+ReM96f/WViBRrGRb9VcZiAyJJ5yxswzok52npcYcOaxIG1LEh
Fj6JRIKocpE2aS6q5Xl0SdRunwgkIr/90BKjIN5lXsxVf0oYuykgxEjvzM39hoewKdt+FOsK7Hw/
SWnc7guhK41OohZVzI5M3NNK87Guc7HG076QWI0MLNOahO2DhEBb3mIBekyiCkxiRYo+l4rbHmN4
v2a0Z2u+aozMg2hy50osX8keNEcv1D3QXfrK7yF1nKDNmlv6l2iWEZJSqA9dkTV37rLMBSwyGSXF
dwCyH9LO6QONlUT1znfyuyIRQoeVPqDUPSAp89zUZuSnlBX8ogaiVwlpN2928GY81/Q1tkAF5XmX
+5lPHGoeDvkKwhO0bcyRvhmtonVA1CKhdeMeZspGBmqqBs0jS9qLNWf420p+lwXUl2RJalLIa+K7
9SvjtMfdhEficwwkw734wMnGp7KpAhPDDav/MdRKpy6MIcrMqXwblLRmTRO+6hifJ6H5PulsMu2P
jJU7qL+H4eAY/6PzJgVzzvLCyac487zwB4ESswIopTkhSrD04W1tj/xqEpNyUJLg0e7UzG5DJSXS
NtuqcDCgeWjGnzrCBcxO9MDtUtbFXE842pbKjfoI91Dkda4ICqmrFavOeomgUChS090gBJkUutyz
eA1r9Um7J+xYYrC2KO8bfaeDEoCHEQ9f9iZgxLCajgT3TJ5LCecSGPWPcUlA43o4/cdrwxQwZmpy
7xdK766Z/lp4n5meR2I5BphbEU1qy0WPwqyUee+IZVpicnUjqSKSK6IDVgfqSi8MXwRsu287hwxy
i6l0+Dugf517hc4a7AL2XWfPrerdQMSazqlGQsCQqdXjxAzJgAh71Z6aVJwkfPZp/iVVEu9PqVxI
evV1jQeXlGfiKZww9NZDRFgWyYQ1MjIsPy/uKtss/ZlipcyClYqwrUUYqTeLt97MafEvfTv1syoZ
jXVijWkeRMHVQfmNho1h2DkmQ171V/Y3gq5PixH3wItM4izSs6MbZ+GDst0BedQ9Ngo7UkNJe8V4
RXzUYWpXLwNmlysADsYIrneTikAD6sbzaCRRjZJPp2EGqiicG5uvQVkfELdJgI+aL13+YB17PSKF
JHk2xYZidJqkE671H+ewBRZpqwTCaCdya8A/U2XGE2fo63WN/Jq7knvWCNazJtpV06MVq8QIH2Ln
jp2945EIZeyrRZsjyPwkIBEbaly8rK6j+WEXU7qSVaOFrMLzkrPTdk+McdrFtmYykBl+rESOJ4Qi
kAAjMXRSyq5zl9oE1I5T+K9xobtB2Ha9M46BVvF8fyvX/1m+pCOHE/SJZfQqaIypAAgNRhZIYFjB
brETm6ce3gkrmWcjF1ayjWfFowqEdY82g7q10aNfPI6PXA9BnJtFIgGA4ncZ8jYg5mtuKH8X/Y77
xRLhH02fPauJTRp2xTmlvU1Nbp8ht/8habCAI16KFCNshnHjALrunOwMrQfstfIeT84wHJ3bAc2q
PZqyRrarNKZwfHu846yevz89IluSiUr9GuP/WsRJMkYwZURewu3i1vHrBO5jTQbJ02hbf+LWd7qC
s/YvY8DUo5CGXmZuHLpgxV2KTccPWzXvoPjLyS4Ed7a78p2/z9dDt3CseKS1VcUtFK8WQ4LqtSvo
nfr/WO98dd8QyWqO+3W9l5yRi2UmZnqw1VgMuyMESECk2QG1/WX8yj9BmLleZGXX0X4e+2cJACLp
7r3RxwNZtEmdFbZjtgHUAEwwLRA8mrHkVTuumUGlPEKc/1SfbR1f+ShiXV6FLIwRouw5dJhp7qo8
fIdvvOPCdIWwcld2cjtmSAWr+VIIOOPunPYGxlpqaOc4rErMTqVDKGEsyLF7gJ18k14+3woOuJq1
Het17fQROkDIZTjXb+qE4SHSpdbbp7v9mIBNor91P3ZzZQ0rvVzl87c7PUy6RcQnZGxIixFlRWc+
MfAjh/2Pir0sJBhzXa8n5D6ZNZq+85xRGip27Gkg7TLsLAomYyWQFZM7IhFpoXLTUKxDwGwPuhZA
/rXvwzRoHgG8kjamrz1JNBFfykxnhQIv0yCikpGjr6dIlIlAShlm/YDoGiWbX9etUlaR/Vvxyjee
FyxB/TIrIAmeWd8dwtnoM804g9lwQvuTt9G2BDrjrNHZymXe58TLLsANN1Nz9x2QrPAvarPidkLl
FoDjbX9uFuJvbWL3nTIyt3cDxZrF6kwTaFhRGPFd434oOpx4UoklCxJwlDiG77RMMqoDrWbGdXIk
L//zNglhPPDMpBP/DceC5xkJGqb/jFH8aHNS9DsT8wI884K9KW3YmGJCKvQUPj96GV4FS3YWJ6xK
Gho4yYHEo/0z6/O7zhlz5vElAxb2yjK4nDY7dqv+idVSzlA5aHQTzgABZ6ZanfbVq1UlCJBdisNz
ITfsElgkcIFzvV8iLT5AIUNCI1+4KeHiEpcxbQy3bdcmR2ZbHkG8UfK4OHkQsNvTAOw9Ls2ATPfL
/OTWydjh+Q7VRacsULA2aByXPbvpN07PB65arHB0blaQphZ4jEcVwmSHJwPt6dHsZtk8YYKov4Ra
XGyFPSc7uk7IMQuR9gXwhN8LkzuABK6preUVkV1qVwXCJB45syQn4R2AcRPBQGIGenHS83Hqz08v
nujuzXf/rsEN9WzGWww3eBHuAkS+DzuqwUpsILETTUIObDuP0fShwzfKtTAP40NJfXoDX8R15xe6
iXceYG5ZlB5C15ZjmhuwiV5m/2nvfM8k7FWIKP1qO3sUesGd4Y6vVQeKDqlqiq9wUIGR1Of5GCY6
bsy/FAOTnvaDGtQMf6VHWH9fNlyIumSSxCnRnRTBcSQE8PwjU/dd0ci167NLJSwUfAytoaAbMkgo
6usQwl5vvBrxT2TpSBZG7eMQNQDghMVOgePGAynKf5Xu1ngqLliCiNKahD4pJhkU/1To82lPfHBx
21aH3AS6aU73XyDlPH0Ylxyq7soAiB40CTzLM3noDH+HjagT0rjGbyxeib43SQP/j5rDPLvoUCGL
M82pj0zCMxA63esKkUD6neSG5FbJnH5Nmipmpiw/B6jwmkH6+pHOyavjdXsfIZ25Apa0dbpvZXlO
IzRU+XpQS9sD0vKgtmjeKvVJNR4ZklVfmQJx5IDhIkUttzwUKXLDeB5IVm2LqiC6y9BvnLrg4Cl/
D/f4Xll3S5pIBub2eclebwpmazHczwT32tGzzrP4lpEFzOyXwTBEkt8C2AjW0tr9bwBU1qUcqA6Q
biidUrilSk99pxEUV9/DY+c3AF+NPK24OvO5KTjIC/1BQeadDKFDdfM0XoXy22mr+ZoMoVwc4+zW
4wMtXms0iOfyEQz1iyTNmZcoVXYrWlt/s4xvu8/8itxdeTPw+rV9EDaMomgvqrcBMpyb+u52FbGa
xVhRNbKrYhOooMr5DEtDGQMWodTzuXKvZH3zJyXpnaeTMUzo3XuxQYYicZZzv4TCwHhIbf+lHi/x
MxfpUKmdNArsGtStsW8xAowzfqLWP8bMOmGEKN+CH985EWLKX1/7P9eO3KNT+sBTiIe2q/EzHsht
ARUHGeadRstT92OcZ6K/VDfKxlStxbXZzszNXcGSNcX1Df2dXK8/iRiE7xW4RElgvQ8647nJZgdk
/hAaDeiggXloOYTsK54icJzmdP6uI5CsVGbkdQV4Q9cLKC9S9MspIvknxXybjkaZ1ztvbAsM/Muu
apuJGgXB3wz2IJRUPQ9DcG680s5esE7Aij91zUuu1ZW1094aa5Z4hcKHWdH1lHkCfCBYTxNcprQE
2PV+u7m3yIYtSE9DnNbK1AV+WvgIIonmAQ8UA8mQ5/AiAb/OVBe1NwQuq0TAkuVtGgOos2tEsCFz
DdclPXAdcN7OdMkoTFIvhpNliK4E1mnXUsnEsUoySBTOZOA/wqLsQ4Dq78H1R54tz+AdAhASQ0V7
xlR43GFHTTcKRt9EVBfLH5vrOXM3y+R1KexP/lYBZm4QQnwsbOoE5EzBtSGA85oh0mpoqxi+clsL
3RH8Nt0gTX3IXwBbT90iwwaXsYspnuOwpyHID2BurOmhZFZzNw64AfHpI1jaGg5ZutpWby5djmMf
lL7oNBIPXfGxQ2B/xU10L53XRnWuFYr0vWU+ZRb2GHh6b6tuMGgyu2BI9VdVCNhJzZC4O9QkZVgL
Uh9YsGEXVkgeoY5DAj7qDoTf/khSqrQoAsrtVEzUmJTXEavB1WIkm3NGMlug/SuS4qJi+Y5mQlNd
A/T7TcjiLiWrtpnMduUOkWQE2QX3MqSa74HId5vSV5Sx0FpDPu4BZblWlz13sD1RrPO92dDpZ21x
t3tXek9gljV0pc+Yp8rNMme3iN/drIvGjJV0T9gEh1uFe0UZ7SQVfzuupletC1Ckd5g/oMWjDqC2
XG2aqUKVEoH4W/m62ET7jwdTJShRtV9Ux1YSidGskvaaI+OUObfaklf/S9tmUa+Qu/ZZTLYX611k
PubSGxOUMe3pwALg/lBfNBR5T7yMbk7okSnyqo3hOWFiMxca7T543vBavxbdVCK03t474ddslVS8
i4GsFgPGZmVUQYxtmyj9S+YFpjifoeVZXT3sMGIEaLN4wohhY5n5zrZHqWD9TDwQscXSxgJ1FTTC
m8wuPosBIp3Vc3yeL7j2KjCJ7agMqF2JHa/f6dftAnHrEqRfiGL+y87dGLheIVH7LIh0nFMEVcMZ
4WzJ6yBnZBkkx2WGn/O3W7a5f3tuNzQHFZNdfD9OM+bgjEb7Ahjq0xQOAc+uIxiCpxSrCbU3nDHj
2YRDFnzvstfOfwaqiWAhTQLj47+6y/UFBTE3FKFHDYnzGKFt/oye2goKG/eI7I3qgoS2zrA+JrwO
mbPYdwMGsbPr3y7a6aWb+3uUCSXnC0gvqBYO2LReJChykeEXXpdjN5zKmnqsIScdMHPtZ8uXw6wH
RJ45HoxUvCx/MW0ZJ5L2fnWiolgqVY7x0wEIxRGELJhTZil1SYZ+6Eke28lkBRd+gwGZMT5jATW6
vh4mi0cKwdpLiRCMjouP/EQnxOtLArrg7CSx4npgFwvGcl4MRCgt1lQMXZyUJsHbLizytZIzFjOi
mZ5C6nshJBApod1Kf7iFAgpSUhONKgDbuPiT5cnFFGLJTuKdEplk4d6VqVYROLmkk0PzBbfEM6XO
CuE3Ak76WCVjcXiPQZbOePCEywesSQPNVpnKWoPtN9iu3ZB/X8gDbTvPW7SvCBzTK9id1jVEzP9i
N5no2nSeJDsLikWb5xtlBDR4nYZg7tEKhjoLJeuJ4CenwUkOycGJ39UPRn2KMvcyxmsEz6P6TP0n
YQap+64w2BmiqOz17LPhfh2wkV3z/fpOPXTm9MKPeK2baXak8/W6iJjv3sV9Mai446Q1w9EcuVCa
tDoybsnK+1WFSA+PuRFYjgywDX/CXdm6C6qVbPy7qtN8LHKm7iRaeyAxgmL/vUNu9/d2PztiRAfU
NzfDWFAN2NeazDmFkaVi5QcuDrLybzWksr/YZ8DMrA1Mb9N/r4yqTfacWxyUPR4XzDvvzvaNKdLq
VC+4DNk/IzvuLoGK+0tV4b4oFTyQFVAEKuUTFimRL6ID7eFHwCmD2hQL40GnPOUz8SeUHnmO311Z
2HJVftJhU0sDT0iPXd6tGiKcng1+7FZCU9brAb44t5mb0VFHMtcdRkSs/62A6L4dScGW1M/its5/
RuMlR653JXwsS21+/ktxeviEX5MMshErhyXBZHsVTdw8aUSRl5dp8fOzNSTtq18TGe533BuKgDJm
NmSB0JlS71lKqwjQogeoXZ7aCvM6bXVGgTU7J6exBjwGsZoCvq3z+v+yZsvPa+a19YH5Fh+Xqj3p
or2ggaXlo5Fe+in7GS1GIr7b3i3v1YrwWgS3H1WNOUfNau4BcenHsvKXgXaKjHOrDkt0RssP0i4n
F5cSGvZovAV9ycmcDMOOHhXxW7VuWUMHA1d+lUdGCusY6XNRnUHHKO+E9sE5TKKsDv4exfOmeZ7R
UaFmNggoBsjhOpUEpHKKDhwWoNMohKBFN7e3XACyr89qlKhg3FQZtRXvn4YCATAXYweLy58H8Hy+
fm/YHhC+sxNjCjSbQfAo0GHSuzzdolT+MaQGljdZ1UoPsO/kZc+9hSq76ytol6jxTCkzFTetcv/y
g83vLdcx3kR1vnjMqDTIPI0fiSfzr0qh8u6q+L9yE4emTey01/DT0OT3OETAaXpeV85RTYQkIbdS
qpaIm2FSLtCCux/5+8wPk5xRlCaJewb2d0ANr9ME52MCNSc0AHWfbrF+0X0iQgs+wI75kETm2NnA
QrGPMwIrCEu8RpccAfYguIwo6gZHURhaGeg3bxeV9GM1Ou4FZA5MUlDYvVNBc6ONHEgN9zC5iLKy
8R7ZJbBIrLIxg3uI6ozuV6AWuNw1JoNIxIjiBdjQgSoYxR9DGZopbik8k3o90/233qNvQTAxrq3X
6MyaNvttPX7LZXhaUfgBizyO9l+/co9tmMc9LLGC7dtIphrDQ4asyEhLNEDX9Z8AwJ128FJdnuGs
+w/Spbl0ZVX4kVC19yVFGEnpMzAzP8B2Y72xVJy7ruPWpnb2Pimt8WaIHPr0rV1kjz8HD7LkhNtL
gycr/0u5inNRMQglayqNM407HZaUCzeXe+1RN9Cq2PpPFJA7+gmriGOz5e9Rm7XDrwQ7yGs+R2p8
iZyfsou4q6d8O3SCW1bZwLn+iN+UCo2osf5yzyUi5u6n/fKaQPbbTmRc5bTnzVnATHvPuy8fXUGD
gnYHwNzTh/24KjuZUMNq0tTk17fYxeWlJVoH4A/nIruW3NydQhnavjNMv7flMybHREwSWvkYf0eA
//njvakp1EPMOIyEeOKQVRNd12fCkunZI+UR03hv/hTGQXfxJ6Ij1no+VcE06Hck7LahST5oqN+q
FoVFlhQOzmM8OlzOZGxidodCvukIOR6UDIej3Al5YjY9MoN3HXCJ0PIC4KVc54i+EDMUhCr57ZES
aGEnZZOqRuSaUJVeDjXeAUXew45hiQG+RbQgONpuZ19KtQCUrcp5GifAxxCFEbb81DFcOdMAz+xQ
9i9W1F1Ckv1MmH90IJkJGdqdfApyfko/6hWFD2RDokNSzm4nMcx++8Bq+EsL79NgtAux5VYTdlnU
O8TjF8ZuvIAn3tAlJbbysjtHqcpaIusTlrUUM8VbesVKXiiFsy6Flo9yKwWprM87D2i0QlQOsXr3
xPGHUvlIjqhNAc13LGntiLian2HIks89kLNRD6yTgrYAcmM8c6RF7SWG0+ESJpBcIap2N5xCgT4g
yO3ZlKbKGh8wagNTzby9YSaoQlacAxcyLgL+DQ2BnNhaVPn7Gea0x9Kk3MDCpPgEoYHf3w+1UAnx
aYYoFet6nvG5bHHE+KW+8bBBCXuDnAKt7mwSOTo4CVOhOOXM9iyPBQl9pHoD5Yc0hWfHzVfYu5AV
GXgqcTFCswFfbjrhmxIzUcu/pVgBVbGPLtuqFv5GyAEy8F/tWfvfjY7HXqR0iJg2FVOlCQycR0I2
nDwm3lNvk5KcsCpcm36VzThTpv+VoaIXEw9XFerI7ZxMgMgwQA1DOSFvGb31WtSaG8ZdCWsypwoO
GY9WzGsH3g/XGHwnSBS8pnDwYviBgmtN28B0JcJsnYPXp3VydUTwC8IXe1q2iPqS0iffO7SxeTrt
s/e0Kqhcmma77JlfQ5m+A0VW0h/Nt02maWafrk3Mb+B6ojHyTfTSi6+YlgV/Pt3YjkPswzuNrE1e
IESEieWScTm54rYhQ8EjVVAVgXqfDaLOfPXEj+a8MeDK1LDaL6PA/iyXkq/DD726URx4aKimmuxH
z/bX3Cjaogy3w67klMCYDP02xoyyn6gmRFPcDxIoX+C3KprNexdBdj5OR+ynWLKmzFsRsARhKGjX
OhMcGiPkTp/ETQ5LAZGU2l5gL0xWJFH84+EKp3ZtQC7rDx1DVNTpnxku2nytWTHXN5qZl+Rbqo+N
QXi0RssXKJV/4CphTEa66pBov85Sw8MlcRAjyPhO3F04ZxxBvU0Kqc4I11qpXIXX+geLUyhQ4Z/U
+vxPK7LDIZcpshCmU5wDJBhxA8JMxQ9ylVw1UP+APOj/jtwmjS06TcyExepbnZ1yp1uXLXtxS9BM
cM8gOIMew3UsAJhtWQ2eHzSc3pPGDzWTR1sn2wjODXKgJ6FvswaVzBEXnA9rY/JY4qSQovxbkXKt
zu4tPh6xKfEZO70L43DuN13fBzv1M6YP5na6ZoThiarD815yEpcTe91aN1fk7wj5fGzB5+3HYiEx
fqA6WO/VBk9Vf0nJL0SBy0ETjQN+nt4eupVPU8801zM21rC4pMHXole9pWc0TmJPZZrAb+t837H2
EICJxFAEE9n0/G3TN8zzxJL7Bn9sRf99UUnwsDdUIRNgYAoW/AB9X/SWUJxNZoznEF+IhBVAS2Mp
IkUVSAiyIBYpPINM+vtXOMrBFQgtJbp5xKFPRQU1DxikNkavxdwKhEG16pB8JEEAmNMT5NVG3TYE
ONdErQ93sgpCJuu9/V67YsquyfqLb96rufB6lN07LIrhb5KfsBsP+78UwFjBIPni6brCkilWjqwP
s9B5ncRd3E2FFUzMbYUUV1QYYay6aFF4GpW1BFwbpKfpxNVdqM0pZSNDlKeWDxdLqtWV6Pscl+5J
3tLXT4odfEiMnAMoeA7fCPOzpyY95P5bmfTWM+F1qxNEFuxh25LrUc7RzOwodo9yIm/sZDw3zdPQ
1BBhuY2MjY+y9m2QHHOd8esamNq/k3H1Kmmw6cWNPE6uSlbExmVxnr7CmnSvkq0KqF4QNEXu++LT
8/BbWtAbcJPZYQ217WYkDYv5BF/8qEmoDCxXUpVPoQU4JkBImUHtVUSFcJ+rA6oDe0ZoVLRljWNA
9h+3AbP0R4RJZYqvo8IBOI8CuyjgQ/pr3hY1m7fiQ5DAo3Nt7/8IKO4TPjPLLuS6zsEAihC0XLW3
/eGqagx95jbA/dJ3eB+IaX1b5HqDlKvO+tIG79AKdjMS5zgI8p3RWBnOtMcpezxT9/9Pf1VufUuo
YCxlG26p2t/RTeh5NnDfQOuPI5rgSE2pQGLbK723mhLhz4VGImEaTUxWKTFlmJj+vC5pQxf/S2m7
3p4Sbg2j+uA8eZnAYil7FTgvZXpEg+y9gfXMptU3NCToJDNFtYM4407JKYIdTmmfLwgHnGAYjzcs
WngLtyaigCbOrqTXgCd1HRY3JAIw1xpH5j6mdUIXhSbDnt2GX/1xrqtwXCNvbxUrbrVzdLd7Y45l
HedbsYyUOAITIm26mCfI+d9xvZ6Qa0C9TukuJqAKZ/GaEq69oHU9K1M35uJo44NS1DvfX9VRQEig
rbHq7OAtaeOR5+8fZAuohMuHHcbbRi6WkRdH2otw+IKDKqXu1heyzMzC4eE+PeTaDd5BAofjSFGT
RW0S1+mcVI3PdxDQs3jpCDCib+hE3JCJCSC7z8xCZk66pFiKIH+Cg6crppwizJJ1ZjN6Qebz1FC1
Yg9BYCnuY9SdDW/hHIctYGRv04iYpp0qE09MOAoJpW1Fa1JKnnlOe9ButFngJ9FhP8JhL6Ocl6mj
/MonVXUbJHJf14O6419Mp47/tUCr952TXwFVZHiVAMfy3+Y3vn2ranOG7iaSJh9PECsKsMvn4whY
E7KmJ+obPJxk2Wqd5RI1GesXrn03ksF7hMui+JOtTSCpMAV3WbG1cSHTHtO9RrNAbb4KUBjdL+W1
h54TsMEDdg8FN39Ez/7YWkN58Igb5kTVDA27KNQmDn8kIcZ0K6Re6mREtnpHdcfzNRnQIKYK/kn2
JxUlHJG3vGfbbu7tlIB2FAbTkqYJ7UDLqqiLj8itRY5imZiJj1FMEjY/MG/6nXHdLLr1pGUbNzQU
UdZ2lGCiwqpWpNrqEA8rjkCiz6wmOu5R1lwTEEydcDZMOjmoctQfhCSTChqHSYOsoJLUaqRWblBR
jfpKMp9gupuHgYsb+d8RkMaN2meDKYKRVl7AjICGcpB3r120AwOjHPVedWy4cTGhdm2YlfzXfd/J
FB0iKgqFVbA/IlJNH3mams5KEF85qmhKQUGcr5f/1lvJlI0/5iaA2VyA/KyxIfl7GBHvw3q3hkdl
3scG3P3Mc8C6L0Nfa79CA2bKKT42zU5Q2QkPKFRm0ZkYkU8siN3Olubl5x7Dwv2iudv3SycVBVel
jNlQPqylQGmxTU+yW2HQYeujp7KtGVsOKUvKFMby9NwKtzBUiAsELbtzxFcxkAm5GAld3QK5n0qG
KRQaSkGgwD3KqZDCnPKqzRo77Icxi4MZtIXoDIoEzBAd+bVGaet2ohA9Pkbr+ZxSE2JmCevTuzMH
lYH+o1BpCzLCHyiNGndHs9q3xDPtdf9qkv6BvuktLN9XkXw/mCKN2DCwSqL1vtneRK/nKc6nzlis
63JVQl+C56Y60RNeIyBJyQ2kpGncytLhw4Dq0h2Q9oGTxoa4lu2rFVW+whY1thgsq4OYlD8s9Wrv
kbCTCw5aSxFoSaDU8QEfiW753zznDyK6zdaSm5Q/u9yQbmtI9taLCXrmoPm1cTM33bgqHwNP34L+
wll2lhBv3mOMstNujbGefRIi8t2nD7KKnwVlsyzxElm0YaP6DsL2rP1qFiTfq6DTZ9iS2YhT7kc0
CucpMxhHRyUzD4HSLLJ2/G2VXtZLMGF//o2ZpM0RWvnS7R170C86yXc1rg4cQ5L/4iVI1VIgZDJs
Qa5bAPSFdTy8rYn4YeWUznTfsPFwZXSuhhyhQCViMJQ3yaTbb3VUdbBR1SPaSwjKOqdyGQHn1ADE
gp5+6DO3GpahsKPKsU5GCJNkv3njqsL1j4zJMD8sTgaU0z+/EMSNhcMZSJO04xkS6nE+9OooM6Je
h+1D2WiQ24WtcIY3GKl7TtjOG5WpU63jMm9/nPcIU+je+wrz3Kjzj4pa2jLmDADrDh3za4uFogwP
2HGcLdj0XF7Ve1ksh8wjv4tKKJ8OXKoj4QyaOCDg45dLqGdE3nVSlgk1QUbYieoWdYl8ypbKMPEe
jHdVcAHF1LRWe9zZ01d/3NuQ6nJexbsmLmdZ7hgxILu05WXCqHu/3Ep2lfpapt5tPfvx0kxFiXjv
YPbKNdkOv6f90OZo9ds7I7qQRa9sy9A3UWLokjv5EVCpvfo4ze78S2kJ+PjtFwBs3EUxBZvc6UbL
GxA2UGNU2uJmFhq3kKv8JMB1CDbi/CAs3Rxh7Yiwck1zLBxg+7FN6qlHWbHLT3Xc9YelPxYWrpQg
FfeOZKXbzgr/omjHVucxhd7iRGGEHsDq+EzvN00vo3b/xEGSBY0784czMj6OuxaIWPYoPX215kOO
zXgKdEu414kQ/F5cRdr1pEiJtJql2rdM3k8pMPZdDzx7jgbWYLOLPnTVGddJLhMWJa4FgvOr2f3O
SI/cbiFx/1M83CyEBNfgI/q1bHuCORy1ROQHgawDrkA0los/6ce2u5ru7e4Io00/mDtNIJcg/OZZ
Q6QtxBMvD+nUyYA5A4SsmB9uZXhaModNPZYbH6HiC9YqAY4d1yZS0RHfuxIyP4uv6aItdltn+Xma
xqKpmqVPRvWGYgB76H/7BslbdDp8YKTn1J5b9gO3RYYDrPLbC4B+mKlt3MJuUoIFVhiPCtSuNnG4
sKIG527ku4wcE6zIpdem8/95z3+frA4Lq47dFPgI1oPdDBfCX61VR5yaMlO/5qerHN/+q43OcToN
Beod1M5b+MFoohkeI7tTrG6wQHfYWb8ElmlJtqhKyvAGsTs+lX7lHkK4XajtDUJ38et9vAmjHoY+
xYULi+io0mT8cFuZe62rQw4RfHL1aigXWVHLx/H95bpI/UEeQgmwXsjt4UbO01Rj+vFsBdQB8zUB
mE1JVH/FtKyZhxr5Bqm9eSzC/knlxvcYrm1Vs4qaiETj+GY5YDgA3O9pW8mhuQglRtFEE7TGIawQ
McPmoD2q5UXQpKLM9qbacmQnRPOrEl9z8boP8aYgDKZffbnSZdbAzhlbBzKmHg94yfYwWq2NGeuG
ej58vLBdBAtgiMhptylHITPbERARC3hcPboAi/0LBzumZkEsWXL/CA+lnTmuEcKJzcAM/FCdddCK
rhNqB142PP0VYtFplrg/uqdrBWkb0RlzXKFdUhcf4q1Vn66tSnRZ7CP2ZlGwgxLMNlA31ouhNBYj
+6W1Bs4UCav9F6JJvXXmf53HF7defFFsokjk//P3RrimWoz5J9XH8W3vm9zb8+N88Rhy+cuJvYST
b79xUtV87X65dPdYpg9yPGHbMa+0y3fPxwQqLbg0Dv6gH6dVKejMhZCFxJF6hEYKu7v/QMSgqFFt
SRlrJNgngkXo66Ki8bawaipthh3kXiTAgIsZ12rGh0t/rm0U5C74UGaRsMPU5xSX33YLffUcKUgl
xTTyghRNSW0aJI6/vVpuiYwHnZJxi5HpHyyq8xIOuuYLFBucaKQVxLCDcGb6+A9LkvWumvsbbLRI
tWH17ulumfngJTTrzEaB5rJlibTfqsrCyFdmGwa+VT9bYLOfRvx91tC/XgputT2TgTgFiazGGA5l
Vqs0SPa5PlUI6aqIrlWaHn+ELK5znIssg27zL320cnu8V6uObaTXPwWDDmPTfjE59+/zdS2tB1Cq
ylLEQVCsS/PFqocsIHZx8G9G70uPvSvRlTu8AhwCxuBbZVFupTnjifMH+ARDRUmKRxvLRYdAyyTq
/GPVINUV5ouUiAOzI7Oox1lPTeQiZcM8giUdgafn98QoRCqulSNAshzw5mGJF7IIZqwF2015IZJc
bbvbCdN68Dm33/35XDO2YF3cJdiJ4rRwhFyNvnp+50pRI+UBNo9BgBNyQFVFKjcLHzLaW3lXCOnA
XsqSm/l4kcj9Mac4Qm7p3jcqPazOXN7WT7TMPnsZIdL9Fe61XIfGWJY1j6aOsBXWThBU4yzhJ6lM
bbuPzMYw/vFLx58yCYWdQ+jeaQ3QrN6BSRqh1gXjubCroV4B1RTIIvfFSafqtD8vG6wgSIbnDWMk
KAy0NIzGrr+fJVA5qZDklnQvm1ZI7IsaT+GhmUTGbFLnPUY8o+2F/e2QB4/U8oBP6PEX5weKRTdO
yBHR2zvCnLsyy5lBY9earaLapN9Tk3occVYu+TI/bWIEpKfTrI3lng3iQZrRAVl2IzbuwjiO49mk
fswoS+RmEXiSDTt4VO3cMxodgrGsC6H1ec/uhHcVGjciF2AI42xSaUmtepUPD9JWfbwQlxlX3q5j
M1XeZU7KphbZ3hraDP1RAPXgT4fpP9ZEHplLxSYzybxQ+uXTDrRkHnhcErK0ZOXep7287ZU04TH6
mnFWmrGTgoJAa6NuRhdtCXxKLEozBan/jvUSxJn7gAMGO/FWp7AH8lLpbO92hEUMx8t4a+p8u9Fv
+x1zPIsvV6ddEBFafOfrQkTczry/0OvecbePQiuWFaJ153ye4h0/rhBMDsITNNEhQR+2UcjKNxC5
MR+hsbBwRbsQ5kag7OZ6d7VAHxYZVYMz4b9Bv6dIKjAVtVDsRD8ng0cqfTMLVnU4vlmiVJg9wgfK
IhiI3F267Z7eflLvkbjFVDYKTrry39Iv1f2mx/aXc5eNkEOFwrjgGnxbI0dlfawnlGWorlS8xyNm
oOMFg7+5AVFoWKKs0WHVq28vgq99EI5SigC774Bz6DdjECioMnsOfoDvKYVmYNNV+71ZA77ozZU2
zqddCzpya8CCHLmA7mmBkcCzsruNQGNCwp5fR+dwMCJkK7sbvc7ZYc+dMTiapP7CbDwJODF0R+nz
7N+/880xRQRmRbNlH5ehMPYGUH6GGvhWAGvIJm+lI47joLQp2Q8drvnjeARXHOjA+IWDaW7qHgqk
pJE8JliXNKdDHwrc8B8IK0plP/nfraEeapwoTdndGh6YS3I7E1VHqjxrieALwTHOGxYQehtRSPwW
kCXhDzJlLgl/5dhKEJcJnT7vdjCt4tbfB04w15mFas9yCoNEaHJMh/fUh2BTPqw2AWQB/njQ3dPj
dHxnFrV0hywKPfOnALltVGqvWeLk9U0nCrZHmm4sU8yaE3hi8n7iI1hCcnelu/wnwVMq13TGo8vd
JmNLGvYVxAc4/0RvYPqRi4oN7FM8PxBbntphrZ7Vbqkum9sPYtre23+32RDhqvo3CoIg3u4MHzEx
pdHHXCOGmQr+ZW6V3N7kGfTH/95CpFlgmZ95ieLZayx9qm/8JJHIxgpVT87pme8BxEoVHj3bCRBp
EIFkBRj0GE/pionpitRaNJaR9xkgMd9EEw50HFGdP+q5c2G76IBb4Xolgex6/cjdUovpx/PZ59gx
2srV5xEOcfDmRyY5hVAt0tMWfU5yBQZBLxKrV3Ds6ZoIN4Dh/C996O1ZpfeKTGIr6LwknbooeIjp
pkfJPvMuUfPAUEP0h1oZVmMTf+lCvyDjRAHhJVJi4Csz78jUZ3HT8VTCt+Bzs5H/ZQli+bLAYPQH
RThtxlMczkEVXfimWq1kRUdJjlejc0TIPIs3sUGIn8qcOpDZRaLRemYRqZWa1Wa0vkw+ZG/QVW1u
izH6JPA282WZg2+noIUYzWRkrbZmjimiHAsW91vS36wUUarCCD4k145HQ3ag0Kdc63oEHKLAz18G
I7+EScS0hJekmwCeCt26nDYbRvqhP0rahEKpm8SdDDcUyOkLzOAgP/EYg3Q4lu8YTtZ4g2M8Ykab
hnLf7dlt8l5kreUdNhuIVMmW+JEr//pjGdH2J/x5MnBzd+kKqqlK3cFxHb4Xb+2Zzrq6i61bfjpM
N87s/1LKj6JpchmZ+hXqNtUNqpGXDPa5Ww60fHAN4F7w2vzXRoiB7KWIFFMLbn3uL8qz8TmOdYh6
U/2NXPDD95iX5a+d+s9c54hIlikFoy4voQcJ7zGPBdLb3RflI5qNkr39WFVYthRLFWyjWKvV2Kgx
N1ElFDITikmAAhLfdt3lM4r3BVvOCMSS0p4uquWD7omLXQriiMSfmSkaW47tk+rY1Kef1P1z6wTV
J97nGH58674jBS/KutMD0Zzt9EisF168WPvOxL3UpKnldF4fCSdQarPNAyZOpU5aZksfDoLy8hq5
eGWVMyko3ssqaLZ/tst2OQvMTesLm1dMVfGyp4ao4o9Kr4L2iLftifRAcZVrPMfzj+LZSY6713UC
1kyYyygMGjoT9SiPUTmvaHZGOeBD9HUO7gMsuPpwmMaa9lhQqhdp+nuRmLisfrSh/ZuDFD3s9YeQ
Z0shCEpeKdhbxnA2QFFgQcdEAm16JS3n6UyxAeCUeWQEXLWEzvKd4CQYrRPzA2h6TR9VE1EvjXfL
pHf5t11dImVCiRSVFbtkGnKPbF21JIH+OXi346LR07Rglm+AkkThuU59NvGRLmE3fVEmRuCrMXNo
Zjv1G20CbWBx5TNPtyXwL+6NWsazpdVgthl/4GzkX2/JRJoDUQbJM2vp5BxDEgjhmhb8nZcFoHW3
NJrP9zWN8Rj/8cWrXduatKGdpLpq7AHDwBNlHjmTnqJIeH3B/MloNAKRPSLWSq9RhQWjvU1xZmW9
wVQjJZ3hMT7MXmSL2uEhEU0cl+p1Ah/RJtH9Z2MIuwwpWyb6x0DGSmxwtrE4XR3npDT+jzxskzDg
OixSPCEIwDBlYD/fYT1pjD8jFTUWgK/6uQLutbIVTvWuJUlD5/2r9OW7MC9/8bInPZ8gIXnNn/1H
Lw4K10vRf6/iTlCxTnwa8hA8zMRB+76OHlAHTp0z+jg+1D0Z8qakbKhFxiJO+zWf9jJ18TO6f42Y
RjO/4BTVPEk+4Q7+yVk/EyVFsWjcqEbfoIio9D0TzpVR1uIyt+SErwNmLpmuFQiu3XQA4tZfNqmP
J/7nQyeyzCHAjIGrFHs69Qlf0RVIruxDZXspN2IV1tUAkyioFgLJTi0tJ9E5Yi0MULeTN++JDoMl
/qmutocc3IHt/ThYFpeHt+73vpbarKCexZ6GpycxC7gYntjsTk8uuJR0TMbx/nJAcyVarOoXzs0W
nOTiGt5pPrXAF6TKvG/gWwUxpB4Ks8YIgjNdbO1pGb1pKEFFdMBLOuciNrBfcrOC6GC9HWh7sg1+
xK6/uVZ+hBg4OUCqQt04WfXi/UTAbLp0C87JWe43KAZ905hrdUlGD7amUOJhK59LIAmeVnVCeXYu
ypYfZRoid5d5VS3rubbmjHjdO45LxwkhLtPP8cdF+rR9Fjltg8xJvauMHDW9XNd7tmY75DJdfKFX
XOptE1o4OZ9iqNs9kgi1lr4oyklFcLOPw89gXM8la1HDTm3KPjtWwtjLuhd10jSQUGIo6mNeaC/b
oiRIdxpJwunxBp7xdoDz89c6fakO5Ta4fDbUZDm7Yr7pdDnpoqVgQhX8XNd8dQJ31Beh7p1jK6X8
e+S9b7TBIl3y0TR7qWENfgRgLwCqiYd/E6pton9G5D0YGEPxpLGBjqLqfbkLsq92EFaX3fcQGJPh
/V+nVHANVkz0WU9Wp9r9qCHfJlfW52hzbFDE7Jk0uuxVsdGYoggVtANXcaHN9qyKwSKW+bOaHx0D
rc3FHV0fKXfd0oK4yiOc7l4wrbLN7u8k2JUuvawmG2KXe+s9ByY7deoBr54h2aIaeCK+alffTAuA
Z5pA3tAvsy8L8h3B1diS8zQTTum6y8YrCuuAiU9Qj/CO1wQlWLG6ReIUC1xE70HFrKYD7KzuFL4I
UTLE2phjWfi5zpKC8oS87EcKKpHq+IcZLCQSty5xYLGtLWzXF8FoVO/Y4u7l9ZrVt9GYEa34VQYa
KW4VW7KPw1Ow4fhBW3abwqCDqaUI6Escy0MEY5YfR6P0dWZLSDqXNwFsKSV2DSkT5Yqv34dhNlrv
HgDGtco6a5jDnG/sR11SUxqeCiEzfGW9itAZrRejEyK58Rrr/+MAoCdflMolv2vBGM/toF/bGncx
j1qSUjNjg5teUjNZaQ/iVfribZ2FTL9Gk6v9Kv05l/As8HGlpyy93UDyscXIUaKVvlfXkG4V65n0
FFXy/fpypf3jP8rSoi6lyZWI1tZtiBE5HX+mTejI8yY+4O6gRaL4G6xFXWQxupSSme/0ekWmWIRv
5doFXvP+VoNUxHYLby3kn2vIaD39wr64G+Bzph0FeDvBBU5jMyMXlaPCwLOdiVMjzDec6IbCzCZ6
6fnIKnxkOz188Cm38ZEQqGXsHKV5Y43nHscSzCSEe789eQUu8bc40n8a5fUCRnDPIcSKnXp6sTh6
wiqTRhsYvedCoWwth9m0/7psmfq2Fy7FskhG2fVithdpUiKarYzCi29KPtXu1JGRDB4btSDyua6Z
UAK6McK5+0W1zBze1Ik7aTvYl8uGGnfQfrcJknUZxEsFOvD1nwMvRhbP1T9SctQGihgkAyEmM0W9
JXNB6t0CwJtbXLRMnaHEFbXPQTqlhpajG/XL9KUIHaBBWZztd5OYhsvXzU3F0rvt9KjU3fOjPdxr
Zr8FY93DHWE1Ge+XZrV6yuRe1aOR9Y+UxOWDeu1LLifDH0GXe23N2y0blTQIU7rUPgnyy4DjOlQQ
xInH2H1ohuzE0syvhmVL+N/RZbYq6r8iiC/AYcstTDB67zoxJFo4chG7AjPpMOEZJPVuU+TS3FmT
ycHkCPZJ4x5tLTp8eLI7Pe41E/iHLs8/K+ktLfgmmGgjusIg+oSN9p+udKoTMt8B5s7dpsSTBbFr
b6Xa4N1tmVUQBLX2X4GaKjsf0krHFE+IwnV1Z8Z9Z6RDg9UxXvFGMm63JEccOj3sM+yXejnSUVC1
b6+HhE87hn2o7zFPeyFsjMxpmjS+5m2D0C+D2yMoxeu3i/sS1V81hLNt5WO8go+7EpkBHyhM8rY4
gzMxabHAX+qS89Dg7fH2jtBfrTyFYrSF+EmARgADMW9ZJo2E9ou8QAl66aURCKSI7qxoJmGFPFwd
ZT4hvxGbvnM04yw2KDbNPKd6PxvCq1Gpm6WHEUWQdcc9YNk4KELxfsgM5Rqg1hJCsKiurUbZz+ch
/FAcwQ0MPVn/5ddaPUcC1HgxNfIkHWigRH+dsmr1FNXFPyHMgIdZOGDSU+1QidSuwQlnUxdZxO/2
oq8XA96y9il3/x0i15pifJytb8yVsPQhJ2IM2RKaiKzEhgGlRytmDbI4+KBPxlqWvvilGDsxav66
IOGef3rePMm+vS4R0KelHyXSmuBnnKwzqai1/FilfXdrI4hjsBd6o8yEq772YIU+GF+dhWngdNVo
9WEaAWRnlfwWg5SyQQg3P5/O+9RkRMEyw6LFQwfMLxfcDLKj4oZNgIL98LWF8nNoZe6vOjpMUGeO
U//0KsY5Q0QWUQu0PyojrTc2hhq3SW6k06l3eIGDSu5Le/BRFv/n79AGLdmhuAvd6fdgj39AfvqW
LTYm1MKtge44DT/6MB+ueiEwthBkfu5eAoJOAZqOoWXF9bmrK1DjFi3Vz6zGYGFyL5IXgCMDob33
h++L0G8JNiFRSwxvx9jkjInn5b1Iidhsc1Lf6qCmb+L1FKVwTQAchwla3mhtlsQ//BLqRQSjTo5M
300e+zYfHzbdFOLtYxwxvtsGWldBP8dDKhH5rXWR1J2QA7L8TcEB2EKtuq0Z6yEvdO1cCiMsMn7p
EH0QQRgXIvBvb7Ukd1eSZLX1YemyGOSNBvFkDPu7oyXXYN/vrLZZVIrjLaMBwsirzAIwTmElUa6O
x8rlyzvE7TIA8cX18XCTx1F6DZUPcSwl9gYFaw8F6oMzSaw9PrPcBnX8noFeTq5xcWXefaf6XZC1
43DDrHCLQ3YYyoNRZJ1bPdWglXQCh/bPYLUmJy+p1U06SDujKcwzv6yUJfZ3wDCe9Jt2RLKo1Un0
zEyOsD/SbwxWZyJlTzCbU9koSHb8STarRfaLjvM5qAngvMRCjSn6p84MiFr6R2tJeeY2lAwPwxvP
zVdvbUaKYjW4/zLxKKyv1xg9KPGtM7MtfnBahkeRK3TUm0SBooXZsCKTVBg3AthUOepOa6OtFt9O
I+fIUdm0kgpccgHOwbioEJVJc5NZl4A5Xr39IySV16a25/m3lIVPK8R/jHXvkKEGGuPQTMn+mTcv
TsBiG8xGwwvrrdOP1TAzpVw8AdQtQoKfVoyr+twlumXHZZYMo2esBWm6BPX2Xx7VUkfJ7UIQRn24
eTJ8nRmr18U3j0og4nKz3UTa9wuUZMl/x9V3KURr8pxSes2jG9KhtOtilVNTC1I7e0JQdWsVMW9Q
wgcUoP1hJFAfaQVsHd3PvQa6oqLOSYeXw2TZBjgEWqwYFnfd0+cmmOECIAd1GGu8o0x55Kg0F60F
YjhKWRj9vVcYbBcSBMjT8QrtjoGVQkuwgKpqozWGO4BYOTGHIpcKGgs+xjU9XcsdE/zTNgtwmuhr
SfFLzxF3bzkPkkVbrjkHbE7Fl8tWzemkg6I+InBPLHEHjvu6RCBJK1jt+MBY4SAaJoZQPBwOEAM9
0o9kQBd+YrydI7NOGZ30bZF9W9v4u2BptN9DpsmwMzEb5cumaTILITvL/bjCjTKD56foFtBN4jUG
h1aXf6Bh/+6uPu0hWsP9CbzaWV+wiCq9lVEMWVvAopbSENVwMKL66BX+nhps7z+vRiGlT+yAYb+u
ef6tJjz8Cm5tdA0J7qQyYaasqE6b3aXnfTash/kUZ/ReGHVDIcy6xIdQDn1qxQ4V9WddjoSKPTlE
j7lAZBNOAt8woY2Fk6UzJmyPKCGLTYYZfE2aMIe2RLAqVCQd1mtgUGIcj0m3b9/N7UeGSRjm7VM4
9Z3mTEhPPwYZ8pWQt3yCPxeOkO06YV+wGlYATWWH/+7BTAfF7oaTc8PU0GTZONkFGAzQs3hxYEOa
sVAtJq2pI11n+R0myZMkTWhvmRquC0tr8rlqobB2dvUdSmbki5HEv0tB5SmahS0uiuLZ/YyhQy4X
jXihkLy/0YU4ZfhGjZvrDSeUXl2Il2Smc2fEl3O1465ieSS35mX8uzA3ce72bNdYtuTyeoLp1SKK
bghV8ebS0+IYuPELpzhBbXFdYu/nDuQyDtLZIn/Zm6rB/gI634mdoo5UdgQYCdTcxOftK9TyY7g2
s4H9v8tiL4EcO75VkQ15koIUNanp+DusADVmah6Qq+eII92ebpqKKXdyksnaAXxpV9wTPz+gSc1z
iGEqjqhCL66ktFeagyLFQ8Eo7+9wp/6/++gizy3L49T/OpW5d3IlJPoyQQfU/qjUOoPpTp7+hBxh
EX8SQZlZ8PCO/R2TiqNhBb3OfQOY8udP2ps8s/k8yeRTwBd4SNhNvhgyJb2pxH/w15SAFV3F2QMu
Xq0YoTpJlSx/rjB+7Z8zqpjz7gwr+BdoTIfYIijyeVMcRoPb49H9Wsxj+HQbKjt8UsJNhCKbvNH9
rtKY7o0D4Y1Oi7WPuvBjk8EjxNVN2hbwE2KQ6lEHVM2a6t+Ux7XQsBuqP3TX61JrWO7qW7ezR4xC
j9M9eHS8ModNzazcj80sxOBesRtwB+v752X2K4z39qkJlkP5bj8OeVIpLu2lLQwf35TXFnNsCv+o
6m428FI3ZyyAjlzIa8O6CNI+c1jcGlI+Srqdk13HiFYRJ9rOv6B/dSdECXlPjVYueSYIC7fWWqy9
iyuyZtRCiUauhRdVjKLQL26dL7dfjuu/mw9To3+tRxPFM7BwkARqjwPygMhdzGBEQJf/6Jp4t5BD
K6LKXG/J2+CtolFz33sU2RhhMHcR9g6P8CTko/Qe7xYwqMW3Exam1DS0Y+zZOX6vDf+UBSeocGFi
y1kXvzuAaREEI9dfa+bahz9xKCD70osNowyhS2BkOP3m1tQHlEuNGX8yAkoKa6PvHHYM2WSp+l5Z
jtsGra+zJTaqVhmd+/FVox+2o7k2asABjHIScUSJJxCZbvnKpL01kTGz1bHLEv2V8QPqvgrOevjb
XfhWgALQtPqxbwl7Njek/19SkmsJ4UzLfUmtQxqy8o15hzMbAbbpDLfu9KUS4dV+G+K+48vO5kk+
UHDfeeBi5CxZF3WsNtLYDtSN2utCl+67Jv/s7t4vI9l9PDb5GzOR5G1bXw0X0BvF4qMrvOwTHnOE
qVcbgA9CQl+yw52qpmHGWKPCZ3M829othnTcbXiBSRWd6eRTr1hUhCWYj1npM/zCdMKBMBntbOYU
a1tmFDhCWD42eKRZnRazAQwAJJqZV6+XuV43NrsEkvJ7zBCf8lpZYjiHzs0lLDYB2trRwJ9QQiq8
5dhHPbsc6A0/99ZTE+hL+A3gLij70S7RsY2oH6PTcaj2yPnTLjV6sTk4+FgymJ7OasxgNdwmrLNK
ev+1haFgZoC7G/XCGiqZvhnUWdu2DuJKLG80DkAFxogkloJsX5W6Ub45+QAty8VVqkoYLAwRDSO8
RIQWyLAwTYYP18g3bEofcgAx8KQloIhc2KQEXfmVtgpvTresRzGyUSMLWJwWGUT5j43fP/uTQvt8
mtiyasEzSEhB8hhaY7lD5fmmfSYBanWwW516mLtdu59rfVQd+B0/foGlaAwRqt3PSuu5AK1co91v
BKdJRbjJ/zjPUj3XfP3/PZKXEPyEWrEnfvoQhFcZlw6tZvse8SJOobf7Gc4zGRuYLinnaIvn8CMy
tKcsGWF2ENR9ZuQbBiKdW1Ms2WnW5T86irU94W+wNmsNUeuNBSDWLkQMoZnDOm1pqkFMnoeVX97l
NbpMlpvl93JXN+lEJ22sLnenvjFGu5gpxrrLonNWsgELnY5G6uSgFoHYNK3kycAEcBrfZ1M2a5U3
O4TCgNpKftBwHq6UF8Cwujao3KgFcPEmyyODbIo5ZFIXGyGI/uk2R1LSanTbV9rMz73ySsHynZDC
Cqx9vlqHh7Zt6b/3tIlM4hJqF5Fma4KQZ6rxj9R1QoJRrmBcvBGa4X19nydsi0dNgBvM2VrkHZs8
4VOrh5ythumU/AU+tD0nS42u8n/UGuaelOdhUo4SpK7Y9oyNK5be2fWJD5lqedSMfb5pt5mVNYEg
RGfBP2JahmJyHIjZRma/2FZxunAoMznrPNYxV9lCa5sABYhx0B3Cfe0e0sL2hjl6+LOXMYy2prkO
tUPiAe3NG+Iix+TGkkV5PZ5envuh6Dw0o5hk4k7vat7sVbS6gYp0RCAYQQQcWGLKiRSNqVtguyAl
aQARMChQmJfj3bUKPTJJ0k218Pm+rfT0MN+na2mZs9ZfZjhIk4CZ/xhoK8gVbo9solzKoc+PKubd
E7WCQn1bivk3On38uZyzvA33BcBJWLuVS3VoHCW63rW71D7MDyhFc/MvfX9gXoDIMQ6lWXDg9kdI
EHKuo3Ofa2WSz4XSTlt77jG57d1auGen1ruo1I7wHdS0ulgZNHs9hoWYTkybRwPzCuCV1IYqJInO
W4jWLLxd5f0/22EGnynl0hpMjlyK4Do83Lnqi6kg1jWYTLW/kl5dxv1uLvD0wjImu5jSCooazRBx
BQBqLUPSR9Z2pukWbedFjE+AcGIbKu7t54QWoiECWVBJd2IpKlxoeLCl3hArIISrk2mDEP792e2X
Vo1bUkfPj8xnFzdTyM9A8rYdCBXcLnvQb6UHVcwb4N/VzZ+rLN5r6/O+kXMqArJTFDIJb4wgVMym
MNYDtedp56oFHXk7OBDM1ZciGG4ejNRyoYq9FcceQbTcwRx+uJ2U/FHZ8GUVvNFKLhtKDDk6gvPu
qeI8+e+ynj31qZc5Ggmh2lEXoxQvcw2ewU82/D2VsLHJ+l4TPs5lAzKG5MAPzEyLOD7W+LXLmK1Q
X7/i7EYvg6m56gC/nU4MMukInwwH8VvrPXhnLB7pCFF21vShnzHXE8V9RhUw0fDIt1f2300sGTw9
GjETtd+IHmmYtwocEJ/A1hQyNG27zeZ+h3nyQy3v93h5nklPLePenk4Epw2pRJlro0zB0Fhzm1p6
JBqG6LIXmOVYE0usU1TbeDfRxpHRJP1KOnJazZ9Q/U4eplOgF/yEcBMlMWR3i5tGkxtsjQMFCXPt
+6FUe2B5rqpi2IAZu+Ijxbly8BYYjL9BEULlrVykB0ggiaYznBVUY1/WRl5BID5OUQTFp3vt2vXs
goyRPOBk7XaSQ6NqZEc1vwoNgQWGmCWCI4GvulXtFeR4pxP7pxs7mB9isJZiNp08dhUIb4QZQz2t
3a/z08bLRgglevuS66dYh5NOpqbLA2u3aGOhwcs3uWNyz2I9SaC7Dpkz1UAJBQqaRA7PHIe2D5bg
Tt7Ye+6dcsWEwAelUQKJRWjer2ZmluZrjdiNq04mZtc52+c4Okt67XIRBlY5kT11+K64Gos19rNw
E61sSczDFVeyDYtxNih2+eZhEK2KxhrEGjwer8LkRNoa3fvP5lSyQUCs/HZJutrG2nqzEvQMWJjl
E4g3PCV9D9SnoxlZRzjSBrJDhBZrAxJ5tomrytatolTnGedc+6+uEEqD5RUzbxb/sCx0xKBcUU2J
M70Lv3hINaHHyVGxe9lxKdhkgKfYog5PmTRUokZy3jaswHxb6j3rR0zeDfGpxqddD0Gq1KdQi2/c
LcIvxCRgPjTwWVLmAKwOFjql1b1lMiCqSZ0NvGYVXpoMXENJ0TjoDBooG+EoB4bc+suBjuawYHVa
vXKfDkgIn0g+OBGjVgb4LfBW3BGo6/+DE63qOGiYXqRpASJpcqmvu9Ld5A6k3Nfiistgrz75jlPy
i87xilexCHbRhgT5uiEFCp9JHtY7RSLqi6q85oMXs80jxI9DpUZfyzEL6IIEFXFS9pnIuRLdPTQr
7QwO6hOB+Susm/ivcw6LkqeffB2LPVYH5IBH1YOC1wvIr8n01qGG4u8g7Li4AmPCIFWS0IjPdcTi
ni5WA6smb9ZRh3ErJCwsL8Th8GsS1TJERlzkqsSPO+lLYI8IJuCgzf+LgEfdqeFh1q6RzPyjK3Jp
SQwhCAfhpV6RktwxjdodD9l7OuxEbZMauTpe/Aes8wmm0eweZqq9YxbVFnsfqplREWQgDAmD04bB
WbxMcfnk/6/Xd0hUUL0oapRv8Fp/rVR4fKdVT640cKl6OphSzKZfqoxbLXptKrUcdWUv7Ixxb7Jv
pDFav5RARWPY7KlW58W3OHsd7UiQ4uKYFRyQYlsx+Y7tKoljd6G+BZKm3HGt+8qEEELOyAxp/gHU
HCIbdxn/whJwU1LfdKicqXwtXDB9fLkBZbFrGjf3xqc3zntSXAeuQyGLECvnlp9InJ/Zd380gzhy
0XHGPdA1F8PmjYrq1HyL17l/SxtknMx5DzWDVnwY2aGt5ffCVA0uA3SzO5+DmxDTbzFzPZV9sbpj
2eShXmwJ9SCwrsT0vfunjac63nqJ/d1b7PeICr/xj+zvsABu/koyvuzLNP6ey1/hHKBAmhiRL43J
bNweDzIdLB6Ek5Kjs5AEZd20DVpnlY3Vzjf4z7sHwY7WHlQbVlGoqdJn2pRX1hsgVgKuUsjbeuIH
hfbJCtHML9E2PgDQDJ3ytWJwQZg3CzAXaKuwzM8aSHQdW9LkE8m0ABttg2QMYaQh8ra4LoB7eYPM
SBYi9St6VDGA1RISyUHgsPawX3YJire4KERvBtnLxNXh3mVuxq99eNeCOjc8cmdDGpPcohPJwpLr
q58TNt7b1ZUQRF5CMtHRyPGG15wq47kT8jKYMqMMAzM7A84WWQqeUno1d1pP6lu3OVQVlcICPNB4
1Yb+IbisKrk/s1O2e/+eUTvRaqjXCWEmZ17qIfvEkQjMfbxzbxYx/qpnEFYe0msxq13fTD0/mj+T
tsa2nr1iKBqweSSHrPyNhLyJ8Y7rxc7sd4jv6t33rqhxnjIYukMkJY3QHF9T11BzXTC9eZpwp3dR
8zQl2qjP6T81qIXoBCTUOjdYECQeFYfbBaaBNjNefZpmvtVyx9Ewkx1EBt/N7Y+YVC6KOw7IIr69
80EgZft+eaFpmdszjA4phTqQGQp0ImqVQ/o4wKW1jKWWcOTGl7bL+SluvOxObVjBlnuLhhdNuOWy
kSRH3c7nC5K5jDGJ33xMU2ZrUESfqOMmyqfeNOLOr8jxwhd2OnsoGYAXCVxpNRo3qm0iuF+QGw3s
bWinKzkx80NiNFUPCCP+ES2O1aDfhcOUVeEZmQqW0W7VvVLInV2/VMkuJ3t7m7MFd0WorS3wtyQH
J3QgVvSLxjEUDCJepYXJW0g6qzoMAonY+qpOLs3QbWUZhSwzJsgxO1GeHjQtXD9+SsKWlHGVVDOU
Y8BEsbpFq1ZRJ9rHTRIeJfhaRqBEFtRUa57/Bpq3N0wAYHXM2/wJHIeU9Q/t30GIM9r0J5Uo/sgT
UwnkXWdocOPDlzSZ5ceGgd3895U1idZT+LijnRM7uSzYIInVFTFVFd1Akg4+qjg+VFyHObsakdU7
GP51DaTfq/Ngi/f1fM7JdTPGCL1uMeTZ2vUT6uBCq6IcUQEzdtMh7of+ELMsLHDPZDdq0TN74qpG
EU/XVqfYuHJ3fTpZB13Qm7cA2o88YYknjXjsIVZo5dRWFGXsUScBptWdOyPU0pjaUtDlPsFSAPK0
bD9YI93TFNDI1VrnKTU/m0W5hV94+1ksJfFCh2bAjuKOO0FOAWLYut0bJY4Hj5lKduZvLM7vwXEQ
C+nG6Nli79cKhpqUO/uSHMdRgTA5rTOIUux2Q/D9vraTZcH8KUsYzvghco/zxuhUOSv3KcnZAh4b
BH1Sn9TKyxDARIOT6i/fz4hTi/fC25KIgFpGIshbPzRiOQiGJ3zMEULV3LRwiEQzY77Sa2Z5QUr9
XRswpaMZYWNYGQKYzzeZQgesKmTGCEeSuchEmvtuFRbbzrWDgX+j6TbBpmsOq7RIOgUc99vaBLX7
RCbwz2JBbFT5v0mHp/M/JM+Wi2ZsMP4KBbwX+Hdva2UVv2N0o+UXWbRtmd6mmKwFlOhabDaD0ywv
LIDeXFLrOqCoT+MIQCWjlk9x+Aj+Z3klDhT2IXVB3LXJGn0So2u1mxC30yhIHJ2O0j5KUE1Pd9Sf
POhJsL5h71ZYKaQViQPcApxaO6IAV3OpTAdSqkOtPQ+dYW4Rs6pvlotg2TdgABGDQhjtqVHXpMv1
bPk6limQQggUZACtCDuYr8d8HosmihdXiqov1dyq9wh0W4HyY0cdsPN+EjaspdMNhWWIawHoZoVM
ND/XXTw/PzqPDkPHT8cnqxS6ymeUQYyjoW/M+iYgI9/gxbTtwOKUTLQyMdnJDjg1yHbZrmrAreO5
gDTfCbLaopMSR8ycwK0XgZNMIwgDOuDU+aG1q2D1nyJAu+cyMJUZJoSIJ++7Apnt7F0nJKWthQCa
dMEOsSJ+GwczcP5I9sO188LC8b3QBrmZtXnf4wpLomZ0h+agnBTHJNzhhFgb2YJo6gDVl0m2574G
tQmS5plz3R6+lFIIVSdyz7/E/G7NhF1mh+eaQgAxHhcfRdQCKwBisFYxSYPF3XoSFW1cLY8G8BYW
zPp5kVHtYoEGONQgU1rIO9PV/vcpXFID8/44JC7/Tuw/Uxjbwllm+wG82ZZz17CH9Snq3pQZM4mN
0F8oXk7mFD1eK5Fx1adZY2K7a+peyU9uIXAY8k6OB0DKWG8sJeIHb8UxmTJankh0OUGH+NmN0Uwy
vR5AR7+htBqSAstpOUZT8sm+SJJPRlEBKR6usZ44YmO9cUoq4hOYFQ4B5f3ItUFEv7HgENEsUmg9
Vbx0e45bWCeydKMUyUh9taPIECfixKsIXtrPKlX45uf8ec/3yK3qFAUnx9OyLc9qVgQZeE7+4c9J
LqsdkBvGaVLcnrDGnCfqIS63u0EXCbDL+6dDfKavJUobRRU5aNlGv+UmzDIdEFDNReA51VyEdJUr
ZdS/GhWs4Mo+25ht8o+XNKyxvfOeQ3iUO9uR3iRQOXhC+jADqNbLqDzkXAP0s/p1fjq8pJftdwue
fRxcyiDmzebYy+5PxdtSBGCik5PoGg2AYd0a/gLnRk/uyr9tIWkaN3zVfJKlNkbKHs7v3KbENWUG
Zd/U7GuDmmVR15LINBYo5anKLRcc7TnUc6shy2wIuFNGo8u7NHeY2FzOhtogycdcIRv6CW355agI
g65w4q5+1CFINXQZVnzmoCjfgffZ1zXZWcJihnu1q5Qrl+wJcgNQU1jsi/D+Sm0LZ0M0H2NnjW0O
W8u4SKq0HaN3NJX1tdxcmAqWnOD02gg+7IXh7LBVYSqMcIuHmIkqeYGU41+PTIARUnTdZ3EWnWzJ
fwMUk5MHAop3/jiOB696yTVrIngQBMWiym22PXCtXiUxy3auhACnIR4oTDd+mUWx2m/WHUCP5iHX
g/y0gNn5YQuuxxZWE4/75a3EbWGqjrdWvWL7L2kwPUpjK2/oGXsB69lDnd8pNdtn1O6/yJu6z36r
Wg2tPh9sJyhWFSefLULiPLNkbQ4M/ud2/7avppqGwFNV7gi3uyggayX5dWVHk804e0FsAyOjdb4B
UdDOe/OWXlwP79V19Ijwl835WVlfMslG+82XdB1A5ijNK1BuBS2e2iNUY5TaLVGiEGPQNModvGlp
MTIatFGbzYnqCTQGyuJCOD9cHLILgmBiZoRkh5fvKigoqr73fRWTJqYwOo+jLR4Fg3thRvCNEScb
zL/kK1rTLlZ11jqPcOz4Z+4ZwQ03coYcS3GQ93U17/8LTdssc9fojtK18woVoh/M9e9dHcDOBqTG
JSvuBV8h207QuqtDgdY8kd7qOUgLC8Ix969Z+HsXAe14L3Lzjn4Iy0moJPlrnHwobcB7HB4AVZKv
u9wemm6B2mVUE/GkMQowCYLRajGXOi0kWluKwVNmy8qsnkp05KWeyyrGxX6EtNiSyYlfyRSUsdwP
GIyKsjPoWsrlt6vC9SR8ap+/sORDOTkqaEJfObGDM59jgdUGCTrdY8eWGcy9+u4mauIvXrQiELyP
+lecFUtBCJIXFSIFSabS5jaZo3Bqh8LcIyv7LOTDBgM6Rms4rWMB9JKxCHOhAgd/dSIHn3GQl5WI
HyqDHQN931XaYvlbBnqGE25JH0lZfzTSo0QXPEGE2z67ONeAvXBg9BfKAAgfTPTGS0UTNHAKqZ6C
yNz9mQBMKTuV08W60DW/yJ7FQU9ehJl3AiPcIJAce3Jysz9gRVjdee3M2cokYejgAxSI1yhHvhNN
cdNlXyv+qptoitb/V3yRV8rase3Rzh/3xhsIyg+4GH8aPcP2VIZMBtIJEkI2sSDMVJbWDALlJLN7
zeBhFIwUbondRsJkpo//qNKd/QIW0UJi8kq8LDqb/aFTsqIYKjdzuECJFPOh1O1vUD9dg3f7EHep
+ZQXmloDGTHLUAEy5l9WOq4WCJbkptm7MbQrsW8KrV6jtiD+uTUMwiBFwc55MSxqZj8CvOy7qibR
4XPvrsZ/iygO9ofPyCKqWYw9IxNQTlN+9o8RZMkMtC/NXf61p3KjILUa5j2wuWfxATWmgbblwxIV
ttWkiB6gSBGlJNi21ez3PtECyvX9gWHMMogwCH1zXRagtQPi6LHwXiVaCxl4ZbU1A1Hd6q2Qm8xi
5fx58R0hOkafkCrq2n3ZES4SE2Xuhu3+ZZiQKD8UsfTkNTsF6jpDVkImjbmNLeW2kUx1uMUI/JBa
O0IdhWD+cdItvyzU1fz/4J7at7MJwLoK7jiyJT9mx7hsBX2BJ8Ov9bOhKzp4RtgcrpSoMqqP3+hQ
+63LzycHVHTROg6duw7FJpEoWDdJBVpPGw6IL0bhmOhrt/6FmDZ6c1JCTIGHB8iFgam5idtjzFfx
x7uP8umolVmxUc0LMieEmE0gykPtMRtgmzI0WlmXh1F/gt96vGImeeFWLkmicmF0Q7aXOZylIG2s
lkgoqmvnYXGJuBa5JPrY4qhhkOIMkglXyX4lhX0vhZDpYpdOFi0D8F93ETclNRR14f+xPZCM0hGr
aJRXZDwFGw4R4bjXkPyeCRLAEpVWeAzP31/kpng84ZdmJ8SxFq1SbPyzh7RL8lQJVqvsOAAF0P/7
DxUHKTN6A579xelEEEikLPSI7UI0eu56OejrxfPk4U7lYXR5LZKlj0dAFVLecjQsC1LkTFLU0tfC
utEgHsjqUZcrtykUfCNzQMo7wV+EyypOXwHql0HHTWP+EHqoln795lVBB/v5g1IPpQVuWD/3roIz
vpiQD3qwhB8Cb7CEgsIpFu+CnhevL9QR3JOxofPchKfyXF/ME82g+kysUs4L6fH3usCamEi3hiZU
EY6Bf17hjrJnDSfSNJTjfvTP3QiuXw4qzXoDIqTfCvsfQ76EACi1C//A0Ednu9Abf1ty9/aef2NQ
CRWOjnQ2prQBasOkzxZ20ghpqpoOxwdDgq55d+lpW97jDulwOMimZJXKErwBECLX+ucVIjxIJNSk
riWIR7u5+bvHNeLNgmEOyBrpa5tpl/993lsNPteF6bIxc5Uxz4u7r+I9Izuz8n1+ij4a+SwxZ4dk
QwpP7AwYTRyu1s2sM0PEliYypNJBKYN2xqQb+nu2BM/dGJ8iy9sSDstmEt9pHMKiBH57Sl4tz5aX
gH59Fm37Xu/54sYMGpIZdIx/8pELDwOYhoWqeRSCSrF2qXbTRuOuUFcTM+05zyy/zsYXlxPLxrer
Uf2p5MOmOFUvaU8V+k8BrwYx6m/AoyMjrAM8DmwBzszkiXNOabol6AVvWGGYIWlblbauzmyHeuJ4
Zpmmd2lWLO8moGOzXIZrZ1+4aslqdZ/GQeV3IPAYyugjL0Vh0ceN+inNjQ48vsTwFNa9TFBw8dTZ
xF0MvrRjtPV4+IyOFyy1V9zOH+loa1j499Q3GNalFKHblM+Qsf7xclObZrenmvlBbzroC2IGuXzg
9M2iy0VoBjO94Ls9vb050voH/r3jWwf5YXo06aKQjgLsM4KmdtNyCF7L77F7MI1gn86SeZBf+4lo
QclUXrYANFrUXIMsDkv1gnNAo/rH+AotIVw+ikTqrDqG674WRnwaeBtsmjYSIGnp9Yr/thKC9+zj
gkMy2d6h4GwPuMeWXHSLzEIceLZAY/ykoEWUVQk67AfoWr0BE8ehWPqT0uHwdw2pheGER2EjaDI7
LHIyrTIYWp4XQ+IW+A6ZfwCh8e8NoEgQt6Am/8uJRgx9bf4iKaoikAWU24947spD/UUkAIUGnE+T
HDyEn29CW+vS+7yBeEWR3KJOw/vvZg6S7b1+XMU8/QaQNIGuFklv+G5lsp236RCcmRYOvww3dNOW
wI13etEwfr0RdAaQABYQ1q2sDugcm4J224zmJKyGcBRIqx/GIolG3Laf+lnV1Y0KB0MrEotUPGko
xWbQHlEb7jiLVJcUBjHMdOj/dkVQbQYwz4cvs2LOkJ9aLB6CmOnM9p93srsSDvCMVuonakuz1J01
sgHWr4qgxviBJ1396GvYysr+zYGC7QO6665N/5pbFbo1i7tlWkzLwLfo9bPzAfYuqbeFW3l8n8Yj
rKTDyxmzEL9h/XrKeVtkDzlXM1gtK1ucIw5x/akShK0rzhYbdmPqrVRNVQ2c0iu4C2Rk6J0kIygW
CvSFeIpo/5EQWY0ZG6Ec8NneeWuXlH1M+ED3yl4CJuI/iI21eSohdknd9rxFzN24wqgmWaNjPkVm
yqmhKGDkN5hZAciI2blYZnL3DdvF3yTJyAKS0Q1W1lHjaoSCbUuAulNGtLwZpGKYtodpqrbfqF+d
d3c0YautKmG7a8d0dcxB1sbDmSVAqsmKruVPhy/d2EXFzUxcgAJkBnATukaCo5G5Bicjs2XBTjjs
dzwtZ6ivqggnICEAZergSqoDeAjXIM9rwIsgiFK2HWcT68oYxk7BHKf99qI6ANyMq9GvhTOA6maQ
PkxWniRoLwfYT6/uuqKJCRPjtMUHVsvJhe+bYqmUNB72HcUmeVLJFJlLnj7DSqi6NfG5uJAEZAbA
uTV5WQD2yeylpCjO9BYmmiYJJgGCn3nVdzqj3HFLisWEo3qUtKZGEwxkPdF7PmHPDgYqiM59mmCR
4/Rov4JW3UcJYMt8vylWU7BVSvKObRK7qzTil20nUCbTyMPVNMvkk5EqWmi01EjoN2HF0R8hiJF3
E94UJ3jtYz6t7ZLgdUNnK5UjBS9dIDq/mp+t2lmf1AIvoWsBuPPBcETan+bS9Kb6UhHA8sKB2Slo
FSZB08xBZqhhDwhoZt8A0z7xJOwImHPZtTr04Mqu/U8bWcI4UM2O9yWdICdKAR23oHkI4CyustnH
3Gp9IHMQ6UMKF7xE4UWTOLBg8vUssk7VV5A8P9srR/lXw/85oVuJ0IEMQEcmtJP8vZSyq42C0WIN
NrJA8iZoQU4SqSWnD+MTwqM5YpbpG//4KXAn34GBaMKJHcvQ+wOnYV2GXl9TCbJHI3ljghtyVOZA
2eDAtyo9hQHBM0QLhx3qcBVeJ+U5ZiLlZ1KSPlIX4OvISFTF4IZscDXM5olB/zuiJ2S/Pa8f9Jv8
Omh6PinOuPh4VDPOec0d2SDjCClsHxYhUvH+1OD57hY3iawv0XcsPw2TnUZrkfqGL5jO24ja6x/M
0brtc6HGhyztprmT9BVi/z1s8HZTAgzsmLhaO1z0grxwMkwMSjK4GK/44k8+vskNEryI3IFz71Pt
/VHlNz+uyXrhqd3KrUV5rn6BsxZRwNiZNuQCugIiXsTncoJ4GAEqZYEhyGO9mrCZf98YGmO3KZ89
K5lSKVyI/OgsO2H92QCQRE244ANiO9skiTsHJOQBGCrn4v4AVGvTM/Xy9uJa4Uq/9x70oiB2/gqK
SMR1/RvIxknyPjMhRA0+f7ZOBdFnXHdubnJhRA4sMZKA8KYkE5V1HUsVMX4vAjk9zmSReI/0wsWi
kCh5OPijayg2g15HaCw3fkAJo8GPwABGujTDDZ/9r4Q6J0LkQHjiaH6NUZoYMgzTf7alkfcSkO+I
8pLQebyWdDbeG8ka87NHts5+l0cH65zxGlH2UkMNILgIuVWQERJ7x4pik2WXiUVzkHgADOjVPd1d
/ESfbSvwWqiEkP8foJy2mBOej0F/VGPykk/WqoFpl5hnMszDwU2IyOIno8ccKMPKpsWv0Sa5nSRp
rSrOcKIF+c3LsFnaYKwJ7EKHoxIO4NOBTfUEQhrUhwf1EsU1rdWR7ojhqD2uU5frxt7XA3lTPbu2
XXd4TfaHg3nAFZQ2eEwZqZqMGlkSmeClKC1kfRIt/2Jp80Q1FDp6SkKOB5B9/ZJxKRzO3lZhBbtJ
kJw6J47XBg2J2X9Kp7VVYUn6nyJJTuEnCuyv63fXuQhMO6UeUaYyAkGIxfsN4m31aswP6nrxYp+V
+rnIZ+tRjVDgyz4lkdzXpRBvYClc76OX7pkUgA5T7EdY7shYhiG13ZxLm/sJIyqLKdvact0wM5wr
RzTRCXoOzAzNUI24cPLXGIny3JXTf3d6B0JDHKizSQj99AFHrD++nLheFjktVL8fJ4BZbRFr9xSi
iCuIpX/PXUgsdzRzjvN0MiF15s8+a0zRicqvF6rFv0StIa2Dx4khJLFtB3JV0IBiKRETS4Y2H2Z+
QH04hlqQU93beKspPAx5KYQ6xYMTX1aNR+nGORaP/yCVJgv3j/epJi0BZLhituYDLtXk4rJiF2+o
VkQmCXOUZLpgDz9gOMgr3Z/E/VV6WtJc6QTSF4j+Arwq9LEmYl2+X52BRlwQc34PpCqC9NdK9ZhY
hHNGv0p21feDqyhU10XODCccaUMWzKYA1eoz+R/gfS1+UwkxSH9JRxEyqaBTAxNStgZSr//prpkT
KHFgC+50opuZoCGzrqtrKnV+CJiZB6b7xfK/aOd6UR4cKdMpFJ3Nhu5/4wixTyWh4me1l0ZsizoE
v93QENp5khBr5g/RVKfz8jK6+bQC3AYyNqvTfKzcywIL3POLyYDlqrxmKO6wcoMv5NffZIN6LRaq
hI7JRwkJsKzH8p7B87xUflu7n2G+q9ml2ASNHRSY002ZnfLL5I+nbN1cijOgIlEVg/BGlyqUWuus
q+aw+E1H3Na3czi3H3dn7ECZjQUfzzHTH4WXEudR3E5PsHwbWEY2hg1jjZIelzswzsQ9JAzM3y94
lrcJ26Y8mdJzJZgGRzi15tXgWYHSDR+2pco2wFmPafKcWgNGnTyVKN/3MQz0r5b/rLwseLp6iiC0
M24CDavmhWL4qvSAjAvj7CigU7kuRikTV4l+jqIRaGL81omi1IqqpDntJ28m9GTxrh6RbsGcExH9
7EE0/uXUcv/pX92aC7Abb+FxjIrtAX3ymtoOWWMlT9C4nDAEg1WRauwT1lUePUgUxnU3rBZh4iqc
y358UbVDMBvulg65X8DLbTwomDuv1xWQq/1F97FD4rIHmh86+NQ/GoikCY/d+HB3lxgM9Vka6QD1
YZd1hfTkfXLjsx4sYNrViMlOQJlNO1sq5rhf9LrBtWFpKB1Ldmt20le0BJIKfbwY/SRWQpXbWi8H
9lh58BLtGBOMnH0tJ/fNWc3atSE8+PVM6XgEdjPajjA/9iKLTNWtwf9pUMNEuvv29vG0BD/W7+/C
1UIR/sNdJK+rCVCX6F8KoJtN4Ms9zymhkwUKD1BWJ00/X1hS7JQzRvzxLuNQNIUHO+rMrDG/JMJC
JMTl8JZ1wlz6KeX8WpRLTYuRfYRgggB8woz1Dg0H1sFGhCmA+9b1scvWMNqtTeGloaOC22JVFf7f
Ev5Rie/C9lMf4kt4WAUk0AGSQpJYhORxU7GjdMGdPhXPGko7c2udvoSAMR+9V31K9wbQOwsXMHaD
PIX/0TBJlt+UiZsFEIFWPHZdcIM4AHShxVC8PtrvX9Jh/x77b7tc0aDGA9h6vbZEIBcbtz9+5ApS
q1BNLumWNzOv919yZYsFzX2Z9dDAbnYQQKGEF3q5diD0wBOXW6pOW3miJ7NOCgJEILttsfBORpwv
YIggcGuLdgeoEfsySg2+Hx/vmEJgYP14+xynZRmMUOJCdzV2h31mSXrOjG3gnuSPa6f1KDaKemB7
PfgXRKhBJtTfSptKi3Wd8bYBCC3v9j4ozD66bUEFPkta6h17KfvgRSuwKaz5EYR6zdw9JDmd4uZV
HgeEcbZTTqndlPtFj4n/4yKq2KjwDQamOAAuz68/Wy93EvuJW164SK7I7H1Ts6yrR5TZmRLk0Xtp
LhG1Nx2U7efujVYi5TiNqtlyx6gyvKqNva5jP5v7hhhrNt8W4O0zHrBKYekwruEA++l9IsgwqwXb
WIOtIklgKz/2s0KNCp39E381nQUXfbFgDWm5ZjIFvjS4mMIAOyiEnUTHqtCYvmr8LX7HE2tvOvTs
UNWlblqNBpSb0oxOGl2O0aPz9FGhCAmNWyuQ7KBfxHUcgF2JUMdj8GUAhzk15UR/DVLEItU2t77/
9iNlMU3bczTibNyiKL9UNloAbILu3G9YyMHPzVqc9UbQfDhcL2f9Gei73oeAWHAhOIhPBMDHjCK/
N7V71PAXagWexiBeubgPFhgI/+nlCdZFmfilJgkyOR0Vh6gNUZHqrLZ9aehTkXUjpRpBa6Kyz3L2
AjQSb19tOf5wYpdd8Pqvjt19ebuYGh2WXqmf4SpyBnQjpjY+/LwIFxnLzJqaO9QQBd6ZeW70Ir1j
ffy18rXuvIq0XwPsVJABWF+r7ge1xUQhmqlC74EiHgF/hJWNVO5TLgwM0IMBbZQ/BJs/8HLliF2Q
AuM3wSfKviR3pPdlRHKAONlAK4i9KYzxV0Ix2Xvd/a2bK1p5fQjsf6R3ZFCiDDsZtQQGuTbZjgae
YI0duDkn2P6rnXhurvwC113kk7YurfaSlWCC7EKCn1zRtRHzhJ2L4HOo2PBK1X9LjPtmVhyr1Lme
Ux81DBE03EZM6VjiESgx7z2IM28C9yD5R2rZjleZMGsgsGfxxmOEBmh5Gwsq6X8vbeXyq48XmTpf
fZxBJNVeLoyLATtEL2LNmXVJwjAfSZKi2YgARjmret4l1gi20t0dOGok/jPH3S6pSA7h8q7Cm1V9
ex4paPe4gcKWqO0q5OlsNNsdW8c7CmaOwsTB/1ykKjfeti9MtaXWtsPfAYszu4oGD/Kf0R6pEzYl
T5Cdi0o4grJtwhozcghDleMqOHrPvLfWOepFVKfB9wl5w7H6KnJbIEvVELKmI28gc3KCDIYq+KXP
hqlxYMDK8xzLZ1GtJ/MujZd1zRJYzC2Vz+GT8Q3uX67yqa9sug9mvHB1bj6Nh122ZNvLowthOR8o
Gc80AfSE9d3nTFkqjiII64mBTCa9OpgBwV80vG4ip3DSebVA7nSwsoHXLds5tFDfqqrO+j6jIGhW
eRPbV/JhCjY4TWP/2IsQgd6CdL6kfY+aIQV4YSRVeoX8e4JJBuX3aaGz1+lR7C3TDolVjt94RLNZ
lIu5x3FRB3LAIwHXE0Sdl3TB3p0ex+PBCtMCqKZZ+Z/gnlxzcQIpeEyk2rWBMjFKSAp64iek79Sk
ry1GF4Ab/gzTGCQJpcGlcJYZVD4Fp6Gt/CM3fVuBr+5lP1pdPsUnTjUjM+g6uVIjVA62fJcRu4l2
abdWRJAszJPXieSFBSqADJ5EU9dqGIPTkTza85CMxgEViNvZBV6A1BCROPMABSt3HGlzC/87rRYl
ZhmddcD8zPQJ0StrTUvlDC4uNNzeHQQ4okG/vH75q0u79ZjTTMeaWTvAEql5PIoqAbBpxY1uAybb
72ZD3yrEQsd8IDkYeAgZM4FScv0Zwz87saOXeFsXSkX1nEYmEUoNJSqytretFyiWhofawJ1Gh/5R
OydLYmHSwMfYcxcdVHdHa5nkUo58qWNbCg8ijnUL9FWHnST/wol2YY+am6fLhhrym+rzDG4O75At
EaKGZFA5r+jONca3eOTLHgQnIu/hojWmCVIR4XHQrSJZXZ1hsQWAgHPBopvPwGSbEAza0ax2g9yt
n62FarkmVtY3x6MltDw8GPArzrLTja8BgDuDYP8eb0BRzgFwaPfZH/uxpz2RkpC34NO7v2Fb9gtP
VPgJZBG+77yVPY5WcQxBvwIbVDsTLAlhkB9kd0CAV6Vkpfmk4bU1Cfc4msSY6lhvtvNbqwcSisN0
xP3g+0qsEggNaDuOVYPvw893xqe+T0WNy3sY2g2+sgRMJD1sOq3mLMov5nzOl6sjeu5UVM7k+e31
bOmCXuwzsb6taCmIibAk7KbJFAz4CTqilbcWcZDPoREGCLfhs2VDgpItAnBmCdc/Fmmq2puI1LH2
nqtjhlOaUbLsJFgfabOiy85iTUPdwO636xDbytI4x/5O6m1y4OFfV8WVWhJ+WiwaQoxRCN9B4LVE
DJU7mV9BEo2k9OWCXlOaujRnPK4lUH+tVxwsiVKJLXLTiRmR6PGrC6OPR3kfZIH6XG0XVSxabfLN
3vIOBluhduvyPPy/HKVRKluq4Dve7i1PRt90clgHzjcU9bN8wuEXKT2VslbLcXg9jBljBZXPmL0a
YmlG05WXJlX78nxYVnBxVPVFtxcAJdtfpZ54+g3YDYOptNaiKrw/Z4QFGbWB2+WxNBIh43pyvzmQ
xGXfs+YWz7yyfAaWGUT1qqgiv0l6APgGcNGlnFk9cKl5hJYMBmgYZHsdWk2TsDL1GJJCDbw/DKFT
zjXNF26BCUH5coH42HYwM8vhuPwRMoT5aDD/xZwkbmYPMvTiZRfW9CDLCgMYv/idstqMbKi4iSoq
mqlOnq7J0Mc3Sta1WnKgSzIVRid+EQv0TqiHwP3S+8XgLSgPajdevMDYfa1vmOAWuVVGED+CCVlX
pfN3k4zzX9yCqa3NT2yS4CMBubRwvaVVhT6ibVAf9gqSYv9JF71bDSgT4DmFclsyXPE3wPYnnbcj
rzYgPwmkV9joeTdilEWuGLC99hN9m41ZEKtvm0h0jAthE3H1HCRcU5fYbJ52lQCQwFCEPj+TCJ5R
UNV8VbH++M0ILIRXHgmcGx7GCWi6nqO/IG9vfaLjRt5ZSI472nGP3skmfBn3tJmxwF2Ez9oQ6Bkx
emzYhXbIvseje3psdwSIeiR7Eh/ksXK3gT22EdhJxhUT/ya++ztrezdi7TT4wnU2SWRurQptgzZQ
yRNowbmeEIh+MaZwRBz7pKat4zs4sUOJLH+52a6zC5X63ah6S6cRldBL3/IkyC097CfKyGyve/kp
T6jzIk0tAratqxi8jcZyWxnrLAeBF1M0f4/JRSbIIgjFjugpvY1Q6yfzSktem1JE5kCs1V1p7VQb
YFwtR6mn0BnwjUCl7qkGOAczaFQxzZgfbcoGh0FK6cfy03zztjBQse91RdoGR4K5iDh47L248q/o
q6X7AD0V0eCwc6wgyvtIc0XXepyOGEQjUfzODkj2Y8t5J+65S3699IfoMgjUCvnY2D7K8fopU2GZ
OpImah0yxTdU6up0cuShg3QgIH/q72nwbH7/NVQHCR3oQVfhFi9uJ7EOxdD6f6LCYrxyANa5exnB
1BJzCCwJYACGM/erU5grzknq2UpsUQ/09Xiwv5kns9fQ3oCjZCVJsEQhTV0oizv/M/PW0O0HOrql
ezlyEGra1CtCdJP4Rgb+UR6f4eOoRfGP5uuUsaQ0xkKdC33TK5jEkKJI7i1Up3msJ1ptyGQirW5m
qIP124XROXgeM+lv5oixOt1LHBd0Xmry5KeVggz9AsAN6ancdci0BgS8xv8dkkzgL+PKSd/LL9xQ
T1FZmQjaAOemR5R9JWyZ4i9bXycGI06GnaZvtGGed1pOXMDagtoVyzqTp3llsHhuBHQZYt5sG5lr
zgfgC6tjN9/YyveaZS08p3hK/xdQZCm47uDdxuDPVAvghp9JKvcfjzy6/B7PVFZURDN3Qqld9ThM
SD7lKqRK20qQjiYpWhSv4GzLjECL6e0CguPk/mHr1S/Q5NXuXABkdjdic5ARAazr1DeQtt3KAgj0
WlmdKRm6+HOTWYkxVb3advqZcFqVa2v07whgzKbWD2gDepVFI/DCNg2xGN2eoOe1i0nYKBlErJST
LOXH0dCNwRHrmovSPyPqTgQ+4Bj9TuaMAeQZocjm8mfVC+B2SanaXIUK6YwY/aj7Ai7gbcdZX/TE
S5Lz6Blh3c5TomJxdXom6OMhg6ThNtA970aDROpLTfVgkaYXdJ2/xgFqjEG+IMcoBmS2M+erI2KQ
hbsepgFJdIYBpbn6GeZkbY0LOVv2f/BosGZy1KvS9ZRCEoizIE+kfjGlFLGsZQ0Y3+SXY/jzxD8G
lItrDsM+ordpQzy+LyrkFmOaFelPe/HbId3/1y7Zp2uGKQtUkdWxkLxQc1VK2WrLf9WVzuzeNInp
DAUVw55iICRBSNBA3JgoA+fvh71HqIEhk/2PiPbePJbwysbke3hhUsCx4gIc7gKCLbwtlsSDGXu4
4ikWLnobzWWIEdUNy6I8u44p4PwxWzRB3nuIOvPKU1J3yz9/hA65wTmyYjcdbTQQ398L5VyG7DFz
zr0hN4x/COsOuXow7TscRQStjkxFt/zon983LrLirUNnE3FQYKD3gePLAym7DoAxOPGVc0eEsl+6
RQmqV9yllrfLczWrIWDyVStq22DGbd9mf7dsVQpqvhxK07Bct/PCJ1DvWoSajyd83vSEk0t3rfjJ
ighLfFcHHhf1hD9+Fv/oDgYlvCbvTRffBJ1zIJYDAeZD4mavqCf9MZDt5CweAggc8Pfouou1l9nK
xmZfCzVSfu+nlbEe2/7Tv/kWznoEwvseS6LrrJhUh4HtYcSwD27j/W9RF+1j+uhSiWNNJ6orD11L
flyHLIAZ2vLvT2MyJ7MnQadj9iIJ/yK8N52nFOLJ1nFHp4tHRSIOagWX/f1LE7c8xcp+cK48I2YW
p1FckH1nyZAtjgVoZxkVQiffOZegVvIFa2fIMLgBfZ323PtIireAIbSYfqKFho+98RfIGIyewHsf
aIe6sU4IfdxNfztHUFk+reaHJ8FWarwueuzZK5x0C8sq7KYo9b3gy8t5bbSHk2OchHuzhdEnpseU
d25k61dRtmOsunXzYAjJq+npFkA60hJ/IEInntTvN1BJQLGwVGO6vz5RLgUaasOw2xtatnFarZs4
ZajFLpeGfvUFgrY0z2aZBV2o2VvZ3lzWlrGwNClaXD36IGFSLpvM8Ta58A5WqMQHwW7FMpGvrq1T
SV1LZp6ktiXGl6DLqMhMaR3Fdrsys7LMj/ZvWlFz/vj16mB2bh09ER5wR0B1di8LBRrUEVj2aSsr
ifydMU2/aJ8y58Xw7ptc/hYMTytBbEiC3PkwgHhUdFN99RcdVpyrqh5w2T2LrV8nZ63SAm1PMzbW
YmfFu6MiutWfmEiEHF5ZbF/MUpcoZ6OhDkqdkNUz5+yjSB4hT4UB7HjsoLFGDFGzHjAFn+cJh8uB
ageknZuGL+iwf4LvpcxhUs48Hq84aL5D889qBswHLY7y0Kq7/X+cHurLAEfjbAXoEb4EZelyWnDG
h+7Dk1qIq8AxE7IZL3etPBr0g/wxVNu22StKeiYrhkPrU5PRPaEwjFkA5LJa0Dcoolv5WcarZFUm
Kaskt6W3n2FzBEodXLbg/yZQeIm9863NOVl8Kr95kVjrFxx/0Yx1EI77X8GlFwK4Ku+toNZysDJ7
BiQODcjW6U/jV4RBjOEtVLUcs7bxs3vClWgEeHEEtxMK/8JVoTtrsPb5uM8cggfDlBU28IdcNOW+
/PIYFWRStv9IXUL6JDz+5nvbXQq1i4Jg9TYMEFpdwozRZ63xlYs0jISbif6MoRHhvCI+D0oD2h/a
Daio/oZUdk0+tYpUa2YLlUb4nYffD83L5CDNwe64erZEUrxndqRzqg5Cb+oT7GJCSWibPPkhlw4n
4Tp1VY8FZ0S3MTTyxrADw66ZKfxQevQo/my44GMgSDsjooAOJrByZFYx26IF+C9CMQm/H0lE49li
Jbm1wmcWIJ6y7fxCWPA25aRmGD0ccVhCDeyyC++pGaMUwlFB1qwN3r2OlknHszb6FKUbBYwvL4CV
Zdh/abbBr9/Zn6nBMpgRVAEx2Wa64HTXSsD+rZ2ReF36Vfitig+zulLmrS+0udwuAAnNKWq+SsTN
aVmPNhM08lmIHsB7qFGZYjL7PNGzcpYBZIwh2j/i+CywvK6OzrhHVoKNoEXsp9U1wNG+iHOkdCil
20K0g5gKx3g/aaDTrGmczhWGjvozzQ0CVle9fGiHr0DMX6Iw4eg5V/WYUeZ4dvICQMp66rxTh69U
z0M39OW9F6YqTjDzAjmYjNuFh2EMNlkBE6zG/9w16kpHmZsM1A+YG04EEIozXh0/5coHTcEMaF/q
PfESDW+kq93dG3hWw0tFLsm+7+mBO6QrNqXzFkO7mWDqo9mHckSdh68yrU9gw3smlYqmp83Qwf6H
g7rVbN3Ie7XFeSkzm/K2CJPmn7nGyBU4CZIKVBGT49I/V2GWDWuwnNgr/aj+m3bvaSNkl0xm1JNa
xKzHPPeaCbexB5RlcmyLivJ7xSLpk+S2daFGZX1pCS+ow0NO4rJAKXylYwdJpUo99v619B4GBxJf
Y1kbnMqrI1a4xMtiKUPOTwZXbTMD1xEk1zf/+mUBnJhZH9GExRb7gpgl9ogCA/7zbUPhpq41HXgu
AoBffHKxC1Du9EymGcPf6aFVNCObzleWF+eifcDSqxaCpnxh939RyxXPA6jIMFDBokUtDmp2/O7w
A8LoeOoSF2I7fFiX/WuGPRNJCY6XC3t20xzlR4GcV9nT9a/y7wSgQxxlbfBsR+S11QmxzZ/fNuCT
F6eNaMmgJTD4eeIhrqApulN9Y01NBhiGvi8SuWb/9H1lWCQiv0y4aVdHXxg7+mHDPSWUpWb4BP9P
BZxq8FIZjyKikDwOm+sz1BPIphXeu6pzm3l+6XphqLULwMuplNhDU4aF7mnqrwBwVcchq8e0axgK
gbmat9VbATSkIGVTy50D32Mc9HfH9yLX7JnsZ4SbjHqGyDjV7kBe/CGXy73xjkImGjZ9vJAD1fpJ
hcMlEftQu0KNpstnJT3/slOdlXOTb1EWNyreOkV2RmKM1x9BI60EHIid3e+JeJbqtXOi+tOEMYYX
/F91zjmZqHXDNGRyzIgTRpvAuMm5oLV+ctzE4siMDt5tkBABW39e6P1ZxDDt5LYPWcyvTYwlx73I
95ge7CMh2DIwZ89JavpnzKENBNqwX8ceBUtuJ1/MtqYpJR/zaB9HHFDjWZc033zKSXKjoQ1mZ85b
S/gtru/0W8s5zuMet4pYXvKKSwvkoCYaH5iWCW6M3cc41wS7RjCK/npo7CIPcMkp+qUAbvfSSHtg
H4T4FZp3CsHQE/AeovjD5W2P0/aDdzJUJsBz3fTJtph9UxmNSdQ4+v5YF1z8HZo92y+ycNq5er8p
YweIf2UZZ9NcRG1x2KVHDG/RJeimYoVognwoVzZBGPXn0LqaKkZdohVcl4RyJc+K50BYASY1fCty
5WPXCUQDO+yWeXtcBT646m52V3XXsXKrh7bh9elq3sWCkUEsVvBn3tMMja78Gnk2dC0ypT/shXeX
/FLgPAFx6GolDF1vXIFbqCe+2zAm8rfOU0bf1QaWRLpShwp4nmOsJezLsUV42KkiTltJqgLtuMMo
F5QPa4aNJgkp/GDivgJ/PQyVl9B+0kwbLpIkn96o3RsvBopA6nkBPOTVuOG0PtMj6U1t+6frLMeM
Xwuh89NHQKWrNNpO61Zi2yzgeesxIJEDHE8tAXL83lNPoiXCR4FTE85ldKjtrxQKCj4QJzASvRF7
AvLNibiCNMFrLWYLsK6VaFdZPbN/FHWoOV5t5Nbd37y52XYGpoexlIPks/LwQWAE+1ncnm2CuPZM
1vG0IK6xKi0U2tDKpJ2ZoBpBwTOTsK/KnvTX9wYg+75SyX4n6oenIsLsQo7UBK3mXzJxAgotv7BA
RVpJgwHSt4y3hCQmGM4xEdU9FMUFafvT8jKUeQ1YBzz5KsqH2W/jeT04lmSlJZ+D0mySlutO3TJ8
Z4hjbqZmIQP3L+aXoyetNCSyVZtBtSCQf0l0Ro/JNSXudviy1FNy/PYUKyiFDQ8ntj8suHTCF40X
ypBkvqkbaa6p8liYaSxDEa/VQ36R0t70iKudleLtGkvJzXED/54taX1ZJEA2qXmgAEAM/HkM4DK2
4yaAiR//aBqh4rm6hkqUk/HmxrqCoaGlE7l+S1m8eYFs1uHxz5pzAsY2X0wBgb9oIC/9/WUZTB+9
RXxoxkzii00r/gGqCjERTpa8zR6/SZF/C+eT4gGzWtm+NRRXVPGvSQo/kk8RVdOjKj46fVmzC6/A
ygPcAo4iNWe4eghMNfaP4O5kZCsxXEIr3QVSpORR919H/mDbFgddjAUuyxM0rEbJNW48SgCBRsnM
L8vHS8hDxcHqd02UEqdt54r7PzqBo0Uv95anlf78yQsCTTr5UsXROxNY+GLYavb/gk6PPeA0uaOC
rUBogYYbCjuLTU5vv8hPbc+waq65YxtZZxWKgECs4rWV6ZpEys+5R7dZIX+6HY0PG2tL7fpYIYLs
LnsuMc7/d44EfuwVdHguhnXpILdS0+21cgMtcTCI2JRPdMhDl6G+bjJH9+38BtUwFKoHxGZRzQh7
U3XqpLLrhpeLN7LBon5SphUdBOy+8/H4+JM2KuAieNPTXyaF1n1zBA25msi+b0OpwoDvot3iGEhO
VaacC47fZQpakkLrbU7aIdU+HabyF/T6r96Pvq1Oi3p/2UobbLJF8VjJhKbOmT5sh3kweiBAjdJ3
3IAMy53DCRQvpATtbBGl1vL/OrLDYt7iUZUQU30N8O+ce/YfFFPdBKpTrY4AJCadRrYp71+zhGrU
25Uc3vzT9oIV3A9RvU7WtbxAXWAZjNFJAIQbrSXZ8djFOCK+VBpW3iUmLdTsX7/3RqeJS0It6eGG
OfsoYC/U7YxzEwVOXO4DvNHjZa5oFMqbOBeYEl63OpNn7fcJjQBfblzrVDQsN7Pl2tbPvwLQ5pxb
Ej1ZcI+E55qp5oWpZ866cOcbqEDL7j9fvFfT5177KWbq6lpMimJ5RLkAF5qNF9c2NGqFM6S5y/oS
8xPpcyh3pFI70tCrGni6nN6lmUvW3TIBkDs6Onx/qiC2RcWD4HSu6j7fpme78tVXCk/05INTksYk
Afm5vjOIHXL9jk9PusRZ9Y3mLo/ERBHOX7v9yty+L2FwBErjbkIqvDV6SrbfZv4EOXYgJbmm6mAJ
ROHlJ2usvVmIQFHK15gATBUByRRJevLdRbbbglKH1lOcmKtVFVFfRvUqRQuml5E1ZZYZJJEjYCcL
saDbuq/1T0qSJKGKlJJI5DLR3Tf1wzBy5wLdaPKu1xDvQwTLzQNiZGKTKtVSesHxyUFYeBu5fKWq
M1gKuTNprkK3Ok8I+bZs2B1DeY5fsth/SpFnmWgnrXf4R9RIn7YpXZ2ugTe5fJhchvJrE+RFmNVS
n2ndsmrY9SrLM3st0TPwTxMGuxXwC5BsKDJNFT7KE2b/k0KQN7fEtUvWsmagaKFcNyRUI3hvcgaM
vBMDoeF4piZKkv7i2i78g5X3ycplhRl9znop/Iu1C5L5yB59C+yGviEH/UfCSlalJ8Y391hVhoQx
+pGObCcY50Ac5zpCAQmWGX17nSeoHbUtr8o4FxtY9nSnDJhjO7kZ0lSS/m/2n/5bGlqCQxsYwdmN
i24qGFX+lMl/+vGZc81YWMyjClSABarMor0UseM0q7snVQKoDarreoNqksaOvWI+I8Vt3ZKJUCqR
ru6M4XmhUrNHBY7rdvUSRDuE7MuEq0XpoKv2ccfGdBa/at2ImSLuSC5t5mB5ZhEH28/s6wEZEX1N
W5pX7DzUsW621EJy13lZVUBWXyS2b1CJMJeGgWOQpYge+rb5r6Swa+Vt6RTBsG25AGiiZKvrmhrZ
iUaJ93vF4TVFPCTNy9tTuZCzoeRA5xuoqmghW8+GetDFC52S5WFX2mXZQfMo6y8jne0b1+VCbkyK
YjX2k1ydhQi1riZwyc69/IDvT2D+MrMbjbdLa1HZZCeU5tGUprg+hUwSXxQtvlLG1iCV5+4L0z/4
OI51ivNwvIt1Cs4vo3GhM36FOkFxwTL6QPRjgMMQ2XkKAqg0jtstgHTLLqyIa7F3xp8/h28DgTD8
RIYKRk9u0FlC54q4zn7TXlkwBgFt6PQPPEEk38dMxW3fnsoUeT9ydRuoqzNllDYHiKNKinV0dUDF
Zc98uhCbmQXLXMdaRWPNEGd6m3oq24+EHTEeXdJ7ctFMZD5H9K64nQ7Ii3IUrCYtTvQkVgbgJn88
Kk/ViSQrphZp8RpG/PTBjxwGYdA76A1g4F00SquEU5j+YFZFyIhA0xyzrDA5a11BK5mtFPHjvbkd
xXCOBH98elisNvM33+a22udT6Gs0hWqlIyQzlxUYnosqnIJpEhZ8ZfuruazEwxxtlEHbBbOMmPKM
sNdtsxLRAAnzQ+cikafErao19aFO4ZFPCMcm4c6P/w7P8Z825CCK+AjMSPiC+YYJYEmoVl/but0Y
FvO0xdOeYh0BWAxTlwxaEEhDeTCbtYizQPmaet2bBZMVkgGc+nWk/tYHwSqea+SDMmWSVmosF1QP
h5ZuBiEMzy/Zr+3u8DzXNTj7eUHy+SBdPzIxorS/e2ebBZ/5MAti7929rWqhJwjwLRDjP6/HCJtC
2Yl6WTxcpaBJAvF/ywnMsz/W01lSUDAs99wnHdLzzcQ9y26xDbQZGyzwl+rJxxDb8qXrpgvgNQRR
l0J6wnMsqcnZU+QezY9K9zD783OmocZLCguQE7jTYlOFsRG4V0Nej1GIQzOBE2U8D4fRlUyiQkNu
5WULF23o4dLX53SxHmfy7+m8dUjVtTKGfBruJwsbfPof21tTjiDV1uatX+BApuaiHkA7FRVdE09u
Y/mFzSioirSyMU+zIwVZCNPuH6r85G7LM9bqkfSvjyAa7i7xFoS7SSmg1w1LqHBu3mdbr2+Zexge
M6LPcu0RLoVsuq4bg9ydaqrd8efRIyFxWA/as7FI2r/ycNgA0GjmSRynmCyjfSJlrJzCxoB9fcRK
BppFoXJq9hVKOS4aad4uJcC4G7ljzCjhkGMTHghMUe+YBG9wPGaiYzpIeLLKrL6JgJ89h4rrk988
00n048Oxy6hXtUABsclt5kTwdiXlCzfmL9LAttj2CQYQMdaPKxil0eRUzEV20D5tdD+lRR/9HNl9
TtPcqaS0LrZlphddFy1uQilwkzaNEFMPE3CTYt4RpwKUA5TTYU15I/G/pDvnqDqacGOKDxDv+tgW
z8EWLeICJw2mdlC49pFVK9LMxel/e7wlo1mM4xcneMTBvLiEnUS834JMCmtU9Yw0gzp9ZtACMlEF
iY2p+1MhAUrvxUa9w7Q7DkB+BePjQde4pAYCYKxQ7No0HAOPIcJUhzayD3xYYu+beQqxQ3XxpENV
rSnv2O8sKEqnaA0Tvsj7w8SXUX+Dl/LHP+9VEX8lX/9zJI90zkvtBHJm2xNcv4ivtlYvsGg63IxB
ylFc/dkoiS2mHzKQc+nBwyxRwhhkxjTKlleCG3sL0PqIl61sPlV6g2Gr2RbqRu8QJJIc1jsOna2I
U3eTuonVQXBJSWFPeFe+L1jUnLur/QKEcHYl2C9pA7EXMa/9/INhes3N8w7SyD2JgkOe04Iusiew
AHWoJEZDwfqHrAiNNIzYzTo/sRJgTpEodQiHrAXbYAYzemdBhc9xAoKsExTcuo9zrpOHg1jNT0Au
wURXMijM/XVJL9m4jyO1I4C3QoCphm7zdeA2ITXHEHGeG8/J28FEsH/aP7NlJrB9BWaePkcGh5su
PhSrLt3WEBYBxjLCiA4DZdpK5N3Nk2En4uEHel4x1873MPD8bD7jTJKAS7ujXSMlb4qvxtd5Va/Y
SbvHkVN2EJyC8n4ofQ6M9JoJdReaYqu+o0Kgou9P/BjAMf1kzF6pCb8+b/KZ9vhHtJKRpKcG+Pr9
0/2km+J8neXienncY3Uv+JFEFwKEro+Fmd6bUWezSTk+nT2I/YMzN6vw7JTyv7S04lsuDMon4GG7
pEfc4S8/CUGev1M1oIg/BtnmP9iiAUSsFoxQQU4uj75ClSrJfElV7XbgqfFRMnVR/Y3Wu8GoQExO
7vnacxw74bn5BgmA06MtO6W5v82XsRDsTgkmliR71cUgrL2D1XMJjaCQu1kOoPoiaUM6q4sy5OZa
Vm8DfWPFHtvPBNm2duqg6o/FqJg6Uspi9CUXPxCZmGTSqSynmKjyFTlMy/qmWkaFcbwrT+S+AIFU
KlIfVd5kv/C0D7ku7fUDlTp+XmX1z0eFeF3TuhpXJkicTUtQRT7ypXIwUqDNBI7r+oXs4JE7kjpE
PF+vcbUS8IfD4MizW5Zq3/gU0y5IAkfDZoHonB8IZ5/3a/57JIF8uTZCIb3HwbaQSeWDjf+TPDp9
KGC8FH3qw+RvjiRn0g9uZ/ZUukWyFQ2BsBFZGsWTfPvNMZn8hiM8kyyxhJM3tr2xdT3JuKgKEC2e
zUhrm4ocLjFL4DaLslyrmLOaYdGqjDNsLsKSaJwHBE5Lb58u0UIkXt192uSCilMIRH+dcviSN/nx
iA3mjasBM/yEWBiIKo4c/9HnpA6mVcVuUjHdc99DQkK4pVbj7Aj+EhQ9YRRDUl/7qj3fnTdi0J87
2oOyspXRGLb2xTSv3B0R+pATuup+CB76MBP75uOHozpNRDUcTtU4aJkCNsxvd032fbe6pqXy1gZ3
j3r2hUnbhBRrVMrqZL1QO1MqaVgggJ7PEjpoirfNH3EvKvwzuK6N3wnyy22obSgvTXJ748Om5CZu
oa10vLxXiTa6230j17u2snPIxSwPVttAPvzorPZ3n3i/UduMHbirRof4CjsrTRbo1Imc3RGY8HXX
MsG7/QMN5rqq4gdPjAslHeKwabI6kTrWMgJhvNJ9UXxXzKqrcOGHrk4kuiScFXHgB124HTQtwxjG
4lNBUVl2ffejS1us1VrP1lKTKgg/KHn8T11wXY42WgrzdSMzu+b4V9eD7lu05EAMbe2FRUBFTC/4
+8PuvHL/QDQVrU0E6EJqm8eeBSeP1/Z+OrnArihHOlJxZop2L4b1gjFfQ990D1uZu/P/+ceA+646
jsFtqyyoQh7i1djSFofxQvtT1JzM8EM2hi68sk04K683qpE7nHs5gEAJXYicrY65BfEmRdAwpkp9
/8qQroOkeo1Vaicmt93hpyqcfeDhe0LPv9JxgIyX3SV14GJXKL4j8RQ4zons8woi9XQ3u0Xvr4++
pO2LGonsy5mZMqx52aldpdohWQyAsHfY/yD7CpZzpZE/aLdQQB53MIcS8To5BrrgXQz1VP3ui3OH
7acwsVOr2bBoOiItD700Nv7aqIkkgMRjChXsjffqaDMr1fAl8aW4aVyS65oyMRqmcFidMJrAMoEW
PSV0dtzukuGLzXaGCWRUjWJDQufAtbbLy84EKLK9rqIIFWhr/PDgsJBY9iZJBIotMPnSlR3NEZAN
AHNGfmSmWT9Owrt16VCNLkH5vWNCznwqZeiZiOwx0Bp4LPUg76pvm9Q8jRC/ZA09pi+zEdrwbgmS
W7ckGTf6/QcJfa6WQ8e80GwCzrbXbVY50iEjwvSAwGXhrfUi0+PjmL1gp7WDDihE1sx+IgbXJUYm
PPXWaPHyGaAjyNqgw9zp0YpPKn8ydwgJUTT2mHDYmdvKVvQGKPKuoIGJ9tn71KL/3t2J3qVlBuyN
eij7Mf8zA6AwclIrYgAgIkt+BPu2iQrJETbeBi9oFEBfAh6Zck0AXbWFoppkPSQ8aQdtNZJGPEHN
3JiP3J96X/PRdpzDUdA05GxjVDVj9Pziyr8hjg/YweM0ZXC+JX3ELXE31dggKPM7LFMAXfLPL5Ce
MLlJzlmUsx5+rUhXk1mv2Ttq/NfgcMwzoKIcubvcsarEIqXpZtxI8zIK8vf13XwvSiJ4sxfOipss
GcIc1+JGXnTnMQ1xvnxwOyNXi0jQTIcQElT7nFszZ52wC1WaArfyDRcT5BVqSv7xHZQtdqXFzZtK
P4JUFK+CL5j/HGRvibI29CjRgHqaEpONYENka3tZ3uhVBh7hcCK3ZBi1rVuPOIT6YUxJnb66WyFv
P1WBs3nzZuynHGqzUIZ5hh3jgcq8Zn+O2OG2K++MkMWgfTfaGxo1Ru89RhxbSoAHZhlnqi0aQRAf
e9Q6VZkfEkLSn0L6hRcy3BT9GWEq/Zokm1MkZWm5oe+N+1skLZSia/MaicVJsECOM2lFMGdcXIfW
3P4b9T2IcRAq7a9edswt7ze7atL3tQr9qkf9C5Z1mhYkcWZDwL2sNzKiysfYRNq9NK44G9vdNEna
afEM3whAisLZ1dLMdfBl/2rvKLd251gDty7PQUT6rSKZmHlZeB/jWPQwTJZaEY29EZCeN7rQDWT0
JQ/skbYEHZnSoazgsYgWugkv9SKl5qXAKkxSLMSeVVFBosOSUeAOzVvLyInLxGsMBt81vBIqkDkx
r8FV98B8eATUa7rrA9Faf0XMK5kVarmCxQZpQmgt6zVrisNnsnUZsegqiUIZ6n6b31yD6HrFKevj
vKlViUzDmJWBBo7O/+1sZUYZUfnc2gN5OFhZYMWr0AP1yw5Yj/P8GBpO8OjFp+CzsOkPsYGAlGtJ
7/nFmIhhm7m4RpI+3V4B2PRCTZ7waszGmzrrlJzqO50RaoxaxvLfzQbNRLgrCTbgYaTcSjruIrkI
FVVo6wVvq1E4iwCpmI0MifJsFR4CgT9ObNHG146Ewj5ASp/iYag/XYinSXvF0X9yIJDpFQEsWWQj
5KUWQBnWkFgXMYhyMoFRvq3a1QMlusSRUwo63f3q9zG2GdlEtw0sK+F8ggpkcCC0VcUvJC7MFEj/
t0msxS+uwnm7psntvMB/qOo6aa2qHMprNS3v9TPrXGqN5Fkih87M51kFecjUyhDNFNzcHtg/GG/w
VMHcv7i7paNuHuh1U0AXHsCJUvFTzKscV/lRdXyX+dP9ULboY3VWnfOxiKKCxRCbYlmtYgtdKu3W
G4X7qmpU1h45oB9BcRFR2wLsi7xM+qhsNdXl8UD19Yx21rfmh7pINeaXqetdLybKq7BzHzPKmxyD
HrB2z1DQLESB5xiMAte87VcO40R5QmtIK8UG1KVPvfeu8/ykkyzYule4evhVgiJT7Gma12xrfcHW
at6x74zgX8gfFnd6N4KAGWITPGOEQjPzT+IjEM2lnSTh7krS9STKtEQdt05LGEYdDY5OTrV5JGg4
DTTLsHEyGRLpWaFptgCUJojikaMCtWW49kJzkbHxvDfT0O4NfUrq+TeRiU7fZFC1HQmbhK3pKjqP
NCXqIQQyJUIjSzj3Jco58jowzFFxQ9lbWXflKM4ZEvk3PdHEAgvNqW2LMyAmBZ/xK3tqDv9zAaWQ
vNXlAnvs/uWZ2C9IaW+1MYDrPMQSkTeys8pkTCsqoiwlykqfh2Cp1MyDIfdUsk/8gFkWDY+5fU64
OndRIAwOxDbwxLJQhkNbfkjofaHRDqPx/y8iAQ37MR2nDITzCnfOD8JywRG76RrA3waeZ1y3eTk3
iqkp5+D7MkHIAdNsTO97166HBWxJvzehBSz+9IYHI4rVTXqTg1ub0SFw1t9lz8nHuOVz7xbUQnF+
72KPNDtJb/Tfr22/xWQeqXVU1CknkNzf0fSr4j4YthFQaVyD/41g9Fx3YtSdc9a81cFaW2zfqs5z
P86q1lABJu0SsWf/rSchqgIoL9p41jQFLwxOos16B8EiYUVDZj0b4lH/AujlNwN1ElIjkXUNmWHC
UTFW4Q/iEsIohQQtKF8sNKN1VFFyyobnM/7bxFxAzkTgXOmn0UY2HbMw87dlmXH8gO1KL7oPlNct
vSVv94WJVWuoTBYbjB+T+9gl6hFwJFYJqHlU8/qb2YEZ+IaqZCUjnbRwLqpfWsGPlrZueS26i+6A
13rY2mj98L1KGdvxfShZaH7ReLxQAJhM9a8GfSObKgbjIqpYtewHoDYh8XfGlv4xBrYPuC7Tyq0t
0XcY+tgb0MO+ev7yVi45rMo+JuYIPtRDmZVU+DBSmxp+t5NdHtsB2IebsNtrdBHFFpp1+PM5dUHf
Bz319dnrU4UaEkeNib+c6Xdag+KxYrHTnrk+yXsRLyOOMpPr87eyVV3C0ONp/QTYXigoX7Y11ucV
fj/tHOwYohiAj5twdKcmliWtoCJr2W2ZjwF4ZsiFb/p1q/CpPsICSuFZdYotnffMrDNn5PCXpS97
dP/yGMFlxtOrxYSmmDvC10rTZ6PgzfUS+2/PMHYiXy7aesPf24QOpQRKUTUxStWfcZgqaXw1kNa1
AU9VAYu6GXpGHKKaGeD2EZI330fVvngGqRIZ+gsc5J1p3J9Cqqli9M9wleFoAIehSy8SBpB1RBy6
xmzE35Yuh/Q0UHbh4syRqNX70Ce/cOfL4OqpWyuUlTOYkuCuYwVGhdQj3l8F3hJf4GxMCiAi+Yd4
UrZFzk0VWbRFhtcxjdYX5J7t9QRQNUopaxr1MGoaKIeg96yMoLKAxMwlMs26tCAdzixOxmLrLGGc
H/HxeVp/8eqbgQvZdgAohSKK3ixkqPiEsR8zdoLAbgF31cwCAY8vMt2FY1QNBYiGd/O/Cuget08T
hAT3jxLYjzIRSmxrbtRh2Jw2w5mYnWR2XGapZr1vetTfzsqHtw57ADvKw9gW+hFQsma4MvvPkibE
9QD1DMkbpLP3AlmdsAKTg8W4LavwKKsXV7Efr9R6APAKNkcrQnPR4T5tS0BsgpvN22YGZNV5CjXc
iGCERFSdjuqRy/DhJELj2vcXK2XRpykI21KmzpGT58pImTMC8Ecqe7el3rwPW0ErohnrJJzArxLk
0hoD2QihwHFfC4DDj87OxOhPiBhS4uXUKfRSGUc1VQu68cEUy8FS1aSrY8Lst47vUXjVvjH5osgV
RvIs1Jb9kkXHUu11LNZdrQGu0kZmwuY3YHjcjc9AkSucMbkUeXElOomX8e18su6IW4PelblrjVkS
4vq6yUp1L936+o8b3pztJxe5fORLptLjOY/7rofPctJVI6x93g96ta6GLRzZgZpfEjA4T++gFhLE
9y2QWjbXSqA19oY1s5Ps8VUrXocso+xyfKLGn3w2Je2stscPdw18jF9rh8/2ItaoyGFKcDPWbXBI
l7GdW0/pA4g6M+gptTJ/toUIg+GHM4ypCTdDCN5SdsGPwOEeFsh/l4Mchvggl1z3po8dLE+NHHjZ
Cxdkh0KwrXMgZG9MTg+5V6vjPTuUgVCmT6wl1KPnGLMwh8IBDI/6rrjhwCUENFxVz7OV8Q90MEqY
EURrUNyiKzB1jfgLI4FS+QoScjD3r7iDWWLBGU+MdxvqnQkfQ69GiXBpD1UJeogeDCAe+G4G1y7P
CkWNuLx9fl2BBwhxFf5sROXL4dEDsgDs7hdl0iO4Fqn4eBz/6xqpTTRSTBXOYI29TNMn/pAZCf/P
jkXp9+zdYxS0uoBEv6ZW8u7jINbcpwBMU7ldimz7ef/mzcGCwP6tzNhr+LZ3jHxrpsqFb0VS+kor
2E5CvSSNYyW6zhl9GTUXmc6e5XrhpecrR4+aBc9JAuUiXNgGtuwJHIgx9px7LXAIe7/AegijF/xw
PMGas1dvhriOxPWNm/V7J86Z8is4tQFPzhjdxUGaZCk0/97kRfs66W/O8mOzmYTPaJoeBygScZtw
MQkk29miJr3ug9OhIEaIcnRuwk1FqBpGgKt/DQAPWd4D1Ep/tZRE0nopHAnreZDPcXX3y1U4uCTf
c6rNgB9P0f39X5+/S67d3NAXwLV4SND/m1LyNPiYMnpdsPXKwbfjP+D++4dVKPM61qy+ymzMzw+n
nguB5qrkf2A93IHhjf7TmZLozezpqENibW1KTeYC3hOPJ7knzo6EWJWQitcCKsqKcBebB5395a9V
tLOke0+MnWJaKm1qHGByqW4LOmu9lxLJfia0KZo+gPK89OyrLj4NGeYh7ixoihnIAS/GjjgowO74
Hoi3zNNP0bYKox27ZY2txULuwo706fRSHd6+bV7QXhRAoiY/iUENB4VSzW9QSYEkv8LATBUdQFK/
o9ZRLXtTz6Q8ItWgwlusjBrbIYR3oNCJnvJ3ky6MhJA/HIPwWtNKuZK5XJH0RRo0+QN74a6+VAzT
f+p98TI7tWRpNQ8AaPgdlHtjEXKm+4gspTC1klZCF/8VHivd31DNBo0/HQGmKMWGF3K97JP34krp
luVXHv+l5rk+mQoMUbA1P93hLGJyEJojGk3AHFw6UJsWC3/ehqCxanRgbTFm96qbbCUEQL+vsJAI
khqIyRylFOs4Pad03RS2Xk9z9vd6S3oatfPBbEbyJNQBrw1lYH8r+ch6rWm00jswU5Y+dtl1UT7m
CmElC88ZfZhfCCc7+FNR7dpPEcJMKCNmeFmIPg3DAL2zf2YnHnXMwmkK/qBV9Qm9sRo/wK/deUi8
mZZ8eMiJVuLqJ3TkrAa8mB93BfXQZkAWIBWmBtY0rayDNSMYrb1RB2ecaAQcOblUbvajMqUOEl3X
NG8Rm8I3eJa0Buz0EUsjZEuoVKdsuO74VLu6c5DDoAE759Ln3spTiOlIQH0HtcFuP/2ehvmc+G1E
oHmfpNqgHcx+rfhjobo58MJBQmbpfmRhMKPEaphaQXGjcAb8lRxNvM2mWLEqDGNwiGZlFYHkplFN
etlZggVdnl0NioCNO5imj6HdYQWQR+z+OITxjIjBh304QnYHOG9tI9YtRd3VnH1eIWuvQu3WuKDq
SLyvv4xFd9wy3vzh5YFjMYocILmPoiPYJzf6lqnYuKRMzO/hzTcRrAOXjXoxrqUr/9f8/VX1K3md
Qrv9SPml+Dw0vVowhN7DMjslZUWzGTPyskn428FPzlyNYWB4c0M0Z+E4JQP/vOkDgt3HpAN3lDyx
L17wW8xBEcrUfAjLJHC6YmLfQUcvvVzVo47GRtPsS9dv8WVYLPK3/BfoBFV+0HupXB4LL7sLmPyd
o6NE6ATex3afun2TjuDBYwBSng0O7JLBO2hS8Xm/r0se5k9ReXDL3PSnEjzVpZH4FH7CIu/XAhjC
rzffw8G5T9t6DY9SmQ0Z8jcQM7mPk+K4HHZN8cAfLBiwzUwfPqpelNvc5cYdnHBKXmjx8YyyzofU
NRnsDHEs3/eqyLLtZ19KGDzvSIUGO0MNdprv0SQC+ZSMr+2/7DIoF/BN+kB7k7RwxVGLoB4MU3aB
i2Qw88GaLhZ7IxMnSzqdsKkK+/OThx5g9ZgllpVGpkK7f41CxnYGw+haTQwz/jCc1Yp+wBYMWE9g
axVi3aIvTVYpGty4SeCT7A2HEembVFbVX2VE2uERN58k5EAiHhGIA/UXO/WD2ojgUBRuqNOiF1VW
BHzzBFt1MplLzQ9GENP/JOt8osZVozNIggFe1/GCq9dTRleMfsW2WLQSVExVZYif3zqLMgmhq+n5
bqSFd4XLTC3esOlV4eXfhHGqe8w3O/0mZYPeP238DpJyPVNhnTQqQ3cfOCvppYuevTGDqvJrcoUL
lWJcjtGavl1jVwIHYgZfJ9VkHvmrNC7oYJZLLxUVnliH4TxgMB52y8qAwHQv2VG7t5irTR5CWZAT
/FYooc0XxbLsduaWF9re29QNsSE2Rc6i0ZaL+Q5qtG5pRCJoTpna47Lyq4CV1ZWnPAtRaS8pzRsB
vXne2Wydh2OWZtm4fX26qiAQzBnb3kOhtuRPWQfGesFltLgIG3PxUKp4gvLXBINT2GUH3Wh3U3mq
SCuhNtUBxq7eKasx77RAHij5EQtKsZ/d9FPRwf77L7EnQUlibI9KCWKwnQGD+NttU8KoWrT/MDpK
ZQGPpCqr2vqizxVBHyAXkJXS8Okpk8EsqMkME9+nbL5Y9P75v0nA13it4Wqe7IxpLWcn1xBQfZBa
nWfunI1ZXJmVlF06ol+vdosNqN6hTG+QqsNtaoWY/eIvv2/u9d5R5sq5/hi6GGD8kDEVU2dCnw1h
H6f9TN7ALRFnLdphL++MvUrD6g7JGsts33H+B29qVFq8iUG5YzcQ9iJ7GLeP1LuTpmet22Qpt6yY
uqvb5SDXY1hB3hj9MPPMbLvfaXWNWgzAA777GUCJWdSHIt0bkKEDWotWj+QQaj5KxCsBGtXNdyhK
7v1VCrimM+sL9j9pbT6N2ZmZKMYlNBix2T4M3RVUcOpmHRa/VS3IO8EhjR4tx+auUxvu6aQmgIVZ
UKypGi8KWPRnn2Lc3t791qyadZooPnBW1tcchbbDlDNFe4pSHNQOJHXUgI2PwWj3D0V0uuRN2GKg
XJRjJMJqi7HX+nyrGnY2EuVwOcwp1PlC+cenizR6FwfgkLrk8VPj98aJ4wBfdtU6/gHwC1rQNjeR
mhQPWU/uoCrEtzj38tMlmtJtveAn7usl1u3DhDpwXO47LhGuc19jQTJMTJqknEt01GwJxO8upz2F
fBawu07L+TI257fTrU4c5KjlHgcKHtWEGW+CcReYZq4D/1Xxl2tX4QihWBk2dM9IyyCLNb7/nbj1
Iv5+OJo5VnWbTByP2Vu4XV40DMfLdovoRILXMYryZ2EXRzTUb9VYeqYQzPzmkpKe+TU1+BJJ90Mk
OtgtDDU0ygTw/jno6Z+mM7uVYWdMtvy64hEJrPqSldppy57SQKYVuWb7cssDZBafsYezYuXyOEyG
G6Ys429PFfFG90I1NGjAVid6c2rMLdL/VLA4tJutLWKsccSN8g1xE4Wo+OXQyKbrhT4hYSsSuYbR
sddWrBuWrtASqxJ83QY373+zlI1VIaebcYB6/vgtHX2D3ZQbMMCp5V0+zaDPRRC6INjy4XVvKScO
TMxMUaPUG6ud2oCZjAL23kRVSsN5+Bmvo81oXoTyZrWsI3Y6M9LDpsQW+QdHP+5J+gioWBPP6dQG
yHTBNp9tvnH33Dfk47IPt1cC7JjVOCRIIbQyV+iClA/4GSH3H1tkxB8z2fTBAYLlRwYClF8WZJq0
zwQGGLvYT4anTyVP9o8i9whquWujvOAh18M3tEXava+ntwbadxhsB2NONvsPmMnp3YRs6QxPyF8T
o8lXMbzm5qrPubP9VU3/z9aB8Kjwz41pkKxMnAEKmY3UMlDFSOZumN5MJu6XRDg5Q2z+z8F3t2Po
NcbWFTnrLMyK/GPcscsB32J3cGebzXAMCAj8DnlSTdNFVe+oxoHokIJ8c6fW/qrLWIBxxZsnIH0/
rqfJUaxKQghTtBtxUuaf2skNrNAX1gJ9YyvWcLEnBHLRjo+EfCjLcHorE0OHJ+Huq1a0J7eOywag
AQT7mimGP8EXAz0zW6wdXZjumXPiZNseigfNWmL3h5lYZJvI0jkpMdofZlzELAAVzM+/mOGqPgWX
9xHhwalJPBNW/Rx0vp6rdopBl+rSFNtX3rWnNR41c0RZgucZ2uLF2uvjvyZhEZzLcUguUfHwmrYq
2ntXfBZwXn4CMbANbJujQi7WAqUQmaCjNaYovq/hMZl5xoLRWeewC40Kj1dznnwqZD8+g9pWhSL/
r0PeQFpx0+/q2JIeKxvMa24ARrMPgueVF9rbOn3rw4mHM6NjmUg2ZKX8GzRAFCeN46uPGguzZNFT
BATssjoWqPHR+r5lULkFfgwwLEYJu91Q13cZbdL/AnC3KJ6BVKcQngh5k+B239WKcResrnJ03Glc
GJitKwNO/E0pXKyDZF3YfpnyKNwO7iUcq/BY8qKTvj51i2sgSsmrPCuH6fBTGcdf0McePJb1ShD6
h8DdHCm632F5N6lUpxpr//qBKzSEXUhqUFXp6lJCCuTvuGZdp+wKSzasrVigilTYy+owTuhe4x7A
lib12xxMfovim6x5R5YUye8TO6itAocYYA3Moym7HTiNAKxiCgAbjGxVA8tdnOfP7qly5pQ8KePr
1wESFztJINEvEnaqj77YmmGgFCxMzJqZV7bO+Pk1FxO1rFyiySLSmbLjfrbRCcTV0+PuthIAMNEl
Bs3jmdj5aPqYMHTgGp5hK0SYju1NjDHRvAYPca/0zqSiM2ThznRTOUC4DcuiE+KrHp3uw7LmTL4b
rJLBCLdp01cMby3s7VxcMovxFp7HEGP6gG3jq8w5+piZUCULIkQQHyEls6hPJJ4YbayhVA9SEyfE
L59OYmCUYR1D1eHZSNsaPF/f2imOJWntNqMymxB7CFJcUPzNh7bZRVa8OHHCGMEuYrdxS4qtXh9N
BXpDMy+63aDYsh8eMMaGW5J4ZEUKtiLKs/zqvZOp7Puyn/lUQAgNFMx9vioSoipeI1P0w+ZDf0t6
N1k1ktsLU5scdZkM3wUTXoqMphFdFLAMogRgQLcK6crPG6ZdRMb+rVP81Jmw6hCFpia0vH7C3dWD
TbhYCmHdnI/9FlRzb/PDOf7ig+lbfMjbEvCCQVjMBguTvAvDkkxWHxQLV26MlkOyb8GADAwGSvMy
TJO9npD5bgGRX2q62kFnmAsQOM6umf8eHrK7P8JVK02EYgcALjnncGOOjczkUvyUjCGJ8weMnWDw
x9Uvxoi5uXmxSSukA4T6gw1maDvuL9NBy5xRxrmNMUH8FYlFHZgbrOurIiNFUzCwuNDDJPRZwvop
Kj2h3mPHAI9fVpbZ3gg/u1gmkSi39vfApFJluyXokk+ns8qU1suLuyOXCHC4mRq2f6R635GtMFVs
c8drH5zK0V/7RR4NvCK+OI/gr9+HjXuSlKBjl9JqsZCSRnL9NIAK6wwRQGRYBGq+sPeKatOoof0g
DJZQ/A2Ih2eMKIh7Jinf+JBN++LMWE+O57y1+WhhO3bP7IIjOjSBr1ALOl/pLzfn4h/SPC/BOECX
HVPBjRNtBilv4D0cVpDbcJeoLx2p5A1nXCfy+nQBwnhHdVjeGX+H0C6JQtxkGH/pqkrsBBVoqKZm
7UTaNbH/VTAigfKRkiyP+2JsXcG3ask2PrNUFTdOiAvdGV2R6WG5GRrBFYufRIt7QxDDue3y7pZc
LLyFLEXMonMrAKUO4dExHfYuT+7dEQlIli9lPaKbdMeYtvZrJ9EZT0pOlCB7T4lh8z2tBdKGIJXw
YJXDka4IAlMXaliIIsIYrtv6ejv+EiaFb2PWpLp7DpuNxEWaL7EJUZwi4AwA1s4dPoLVB7K32VZZ
XtUwUSnyoNOF5tpUNdx1jyrsz8yUOpQK9+NgqBGf8HyL1bfHeeM2qjWabzVLhp8evaYXKphhVfT7
apd9FGeuIYxt922dRYyNVYPPAWGv+lwXD3LQXiKlmt69g9ByNjESOhmpgVFmoA7bAzqfivtQH4VX
E/sCjkOp3tvY2zNnneO0c2/+OnrCDX7atNfAKn8+OzE9/X3lFY8gw+KQXxHXtmp0ZbmVg05RJvFl
zxrcgWmtPqwOa/102y5pj/kxHCFboHvZnpuOUmgUQ5YIxrU5SHW2UB1pDv0sSYnQhzxrtQzpzmNz
kadM4qsVDJopXXqZo7bUBxzjjhUrJ5QV2DhIZPdIvHzg19/3QnE9avSllL+nfy4GUn0WlpaGPasT
7fHJhMAoUeL7NxT2RZB3ITqWRN+iyOiUeLhXShcd8LgXKGHkpBUTUCD51+evRRY8JTLg1GV50MYM
TZWA4hQlyx9JpHNSzQSC7OjIb2GbFmEDW+laFL9wTKGWQdeTTg1vQSsDYkebsesnHP/ogJUn1Lix
E0Z0PR2wv3beHiGAqYy8hRo9NlgKJsDly/PCvgUK94yilPn0XzluX8BLMk+VQOojXwJfuPzwb2g7
whQbi+RV9gqur4chY579mMg45Evc1Och0OW+oBxKFDNp60lzyfUcoswlMBINP3MNT6Ar4QBjBQ6Z
J+vxSM9qKKoElIlwBih6s3WnODKnOzn5wZ73v0QWvZY8swkxcKUxhmWD0Dwm6MxeOO7XY58nYKSM
mwjCMIzG7Oa3S+76SvvZ40jk79HHxD4iwOcRdMjAqsztJ29d1789/4do4ziuRv2hMV+Y7SZB+uKr
o8Uyrp6oSGW8wEzJGtXCnaWIESlxlBMwZfXRJo6ZzzKjNe70szn22kJIfyMF2WTJI4F/Ynosb9Ej
WV18avd01MbfiAKsD3yJS3jmFONurKJcN/CKfiWtr9NpI+uWK1RA6ypHCYuvvrRQdcnz9HXc2mFg
SexjwRTA3TQAwvzAWYIKR2d0VQ0Ah8q2pbKiRbwUecoEEQ5SYfq4sTUbN3BU86hZQG1eIcypRtti
yxuAmSfd801251muwjCOKsbtRBOl/VtB78aVy92Ye206UifnogDym4BeEevUjagEgPgBm/QREgVm
OCRBDEqdCLD7tP6bZY/5zvY2JJwoN9gH9+5+9TlZBRcwYZMbHT34tAI2+sxiG1ru4LMrBEr8Bdf8
eBoiZluuaJ6UgHVD8buFWm4H64dtyhJhuj7DB4srAB7ZoH14ejljKpC/nXToB1L/gbME/0B8hIlM
Bch4lrVrHsO5ObFpgj54aS+4JGNcDNdVrQT4yZouzQ8xvhCsu/RD4+1BJHhuOux4l3/6ySwHjMXc
gQYpC1vIeFSVbRouWBKxK6u02aFI6QyxZPG3vfavZ3ugpsXEYU29P01kxiJy9uXFR7+rjq4yyLGQ
NzBdzOl21JA/rSqTEia07bzXb5VsJeg3/LGVbZEqfq22ZaiPx1d/cCWodroPTSuyUbVqFUzK9tui
c9n9hGJwE8/hjyoJ8umUJb/+PRgFODudiVgBGGUVCcxAmVqUCwj+GES8dJ70O0zPD3LBKnuO6LEN
cTQUZN/jhHq5CHW8kHDEb9x20Mdbl5Q1nJjs2cyvR6H20hK6hkXUdVi+Y/f43IBl5EDhrEZ3LuRo
T2a70P09kynzUoIvrZRaUMzGZFEK7AeJGbJVIvT/Wg5KfJySddYc3Iu0KDo2rtM3K0838zXXQ1zf
c4Y4IE9s4SHZ2KM9EfeMgnfhNCNqIREGLzDIcr0HXU3rXKpRmsFer0LvnEQLyP1lnPz6TK4zG15F
PUkLabSLHY76uTM4XegP5knlWW5JjCeub4CnqVJBY0mT4r54p0OT1tAKOhxl99ElYkXWDa4cex3B
YGGl/KDb8jbYaerVUngstQGDzsSPI0UUeAC+E/Szpoyx5iyy4nOtzAnLd4VtmWkPYHAfV8IdpXkG
/e28Yr8sycc8SH1Tdjcb4GwBbORW9w6KQiUJcsUqHxaof0S1KQsTPiVQBuJ2PSpkrN9FPJvh3y5M
3QFypTxwKkMUY0VzIQXO0Wy5KU40VBZwJcDnPtM308kGftizY9VLMO5i0woFGl61kx2nNxbNMFvw
a6X1VSCwZXG0LlrKTED77y0fuQmeQxInRcVjMXt8YZPysnDtbkSJEM6olzGU65VRlWszqKnvuC4Z
PNVYI/Un3gwrIkQIaKVtFUsA33i8ZVfSGCKjtncL8hnGuUjD6Q7RcPmlTPhIICWB/5YS1byOS93i
jT/OudM5wHpvSepyhITb86PuqiftsGFe8l6YjAGZJznbXJXmdtz64HB06GjKCDlofuEcQRfzaeWl
L2gftE2UvAF8goyipz0IZSnr83XWZYCd4zqSgc0ZTUnL+YrfugZgtn5JReCehTBLYfw+HSHNGqfL
Xgj/fZnKNl664XgumnCLbedLj1EG+K9vcFBUr9Ml7Q+ngts9v7pbmSf+5mLPyKKJczU1yiPsF36m
dAPcdzhuDuZXKm3/wY1ff+C0C7M3JMSOTpMyKAkPT0drxYGYXe3cFVAYgmw6I+pocRkUAmoorhge
78KZgkZI8rKbDJnlWhfvauXDsk7VbAC7UODm5DRJN4AsNGzHUPH1UsdXC3L3DqFo4NaRnLe1TOq5
2AEAf4ICgqWkaRWjwH4lsAL0P1qVoTpMKR8uNonDPjxVLNXjUHH/PYQcQR1cdgPoJYyRujhOmLix
n/ouOfwKWlYX6FturdXwO4MYqOaltIiSeTZ4fU9x3pButk5U4ocNSNUCqFsnyKiV1/v4h7n87JHv
rtliJ6yUktY0GGn1VagcJ0BuOsJlHNaH5jZNKa4subPfAjcS3NncIqB/7+ETn6vgnbm4eV5OGW4p
Jb8VSdVw7X7+NkHPP/ZP0ncpugMqF+RnrtAqKQ8oeaA5WebLFzXy/CZUBKhKCpbO5UcHDYHpOq3f
Cv2wGjW3AB/5OFMkrUadjFjb/UaH6yTe5c1hC1lf5jXWi54rhgOUOHgl0OnaBTN2SdA51GxbU8OM
I+nguyx8MHhjUg1iehBZTgtrlKuLCxTPGxDDszyQ9fC306U3qONKOkxIqIYvGco9XUCC7puMlDxu
lOOOP6FISnJnwBiAbQtXJXQtCHPfUGJUdGFw/efiR5rkaEq0R2Ij3FIA/k4tYb96gTZVJqCfTZmk
BQfySiP3cSJH4PdoFYnVcKGxds0pKZar+8CUZOHF+lunrH4ctdt0sUMX0mopIkmmPHr0YNQTGywG
rahR+hArg76h68UkBufdttkU6saNBCsX2m2Xbn8GUIsB2S4ShcBXh77W5xwkLsxjKWD/w8c4ptzk
XtkKUeBqxpX4PvOWd7pElMuH2f4PPPSB1WZt2n2BHgbibOoKn4EjmRFKXR+bBorgR35GkMm0rdhw
ZzBo0smVv4pLNyRWosVS+r2K29Jfb4pIztMFBR014szZ7M30AmDuJXg7HLFm26n+5aOiyv/D5Eir
U9sWoEyhLmHA/80VZ87051+CvUQZyNWHNb6broNLkzJlQRZGmf0VIoWvuiPgxyhQhZ0O3K1jhIsU
9naPmPSnBm5jNeRzOMXMgZUkH8qVXiWT380sSETSowe8YuOWh+w1mlPHxcsQDhcMt/i4scZVOEup
mh6O3KY1mk432zpmgl3oAuiZBDZke3YrjnS5P8cpeSoKTzaAVld9khG72TflM0gejVSxUCyJPE71
bz8JLzzKG+PZ1MYJa+/KyoG0dCHyDhA6/nWZcq/VwutDBS+XjQxQaDmVINe70YskM6mmvA7tvDVK
Uk6U8OAV5WXzzzUKOu3Rmm3qWpUmLf2gwy9QhTqqrChY0PK9b32QNAfUcfsYOHlOXaI5oancsSqr
EtiBag56TdEh0CMjhVFDe1+c4RV4pHWZpu61vH5+wm/qtS0SYOGUwH1D0BdcqR9IRypFJ79EhpsK
fvZhkccUYaobUJ7g/1R16uRoar5ECwsvDe6aGU9PBAVHZjpjSS2I/aPwoPX/tgWXltssQKtcJgl2
1uTTAMJ9syOq4FbxgLLO1hUvREFFt3wkrRK+XYJTYyCvBpCijvx1NaCOtNJqADIshUa8wA6c6Xzv
QBNOZJxm5IK96kqMdUQ78LWvwWre2UHbFlwNfk86egV5jcwNiAc5n6NYG/stIDY6wIMinfv1figF
3yYCUkGzcnLNpxgtSZcLhdrRtjPulU+9UwslyBYzymE879OkYYJoS1rdfrKnVWzva+qBdMQ92eRf
qEoQB4armCtWq9gUXjyZGnGRuE/OiJgotJqDqxqFp9ecqWgq7FqcyvKSfco05uMOH2FuyuG3rLfl
P2LxRMS1SVyxZIhtAJ4ZGhv3LmRDLpwWDBKvkJmst7G5C4GqMs3FRrN9BTgsZtMWSY2mVotELXVO
jhhtOrM72KOpM5g9npdj+l6O+JWoLRU2J5qkr56sIUIy65736l2BdxbX/mEWGmgfxBIC6Gsv1lgf
L9GHvmH6QljgSBI9x6gZ5IFNDqaKxdhTpcHaKjEK8HtR94YGb9vtOFPDIHLB382ovsBwGTbF/DP5
gce0xA6Lbdgs+93GMU0ljqzBjLr2OVSUXSokEyRNIHu7DMopnzOXfUupZL5r6Lyp3LZoXrng7Qj8
W5OhiMCDrRz6J5OkcFQaVwaNWw/B4Hc9R1Qn/W07GUXBXSdtsH2Dks9NNr0BJG5SZLPUDwCG07od
6il50KAZXFs2NAyHSPI4xTHYG6EobPAGkIapAMIWDOp8YEHrYlGERYJthg7WuAzgZXy8MGhZeoTl
qtRZDS0Ax8F7dBckY0oDwyYX8Bbmm0c8ol5Jb7Lx7nZF1yil+ZfFnyZR2eKoO+OmOYrYI3iFtBx8
qUKYgA9oP+0dJ0zZl5cyq7d/1QicXrFthwVVUpnWJj6+e9foHl9SQ0l0eisfDGqqPEyhagoMZj8t
t9HtVyqmj1qqeVPeL3Qfof2SIOQ7/NG0pJMwgU/lV1hDIbyMwi+T7/Vq+BDPEhYl5QK7qMT0olNp
JBu1mlTPol4MY91BdSC+mTuWMtLbwUAtNTfjdaLbxBAcEmoJ7O1+yA5Zp76pj5/cdbFBo6WmoZtG
KxK7sUAZb5CafrtZSyVQi9RHWLjgtFVRW6BgdjIOj4vl+lzRhQtN8urztMNIa3Wv28u5gTs+4hTq
tcsLkmRjLUgFtVdzG+fSXJTCFDbM4fswlt9/O4SrSQmD69pTqbWDXDrtSpTVlyFziNak7P33yS9O
e8N5hg2/dP87cG0aTfGEGBkOhXOnlN63pg2lD4MZ2Q6ETz/VbyILeCMKZJFD8IRUfdw1RkNQt46/
TNG6+6J+77eb3JAOa0bJuI2o+c0hURECh1tj6ZGjN0o2GjBZkyuhB7LVvkenFLtspgF2AvEwKVpj
mXwW2b/8myB8PZe4COCiSPNzDBXL5c49pxpaAcjxguHs3otaOKzYSAWvoZl3aOvGdE7cFFeB0Hlx
GNI5AcojMi0HqVADyP05HadpQ+7LUQIseVh8LyMC51Ml/6opPuPEp+Rl74ZOyQ5af672TFHAH3Bk
Vj8Hen4JGtpAOUTL6Yj5gsftRcgCRxNk3/EAiO1rHRW0b6oh+/UqtOlUPMn5/TNIGsRkzJSJWy2N
+pD6AOefYMGBYwfkvaXSBNJpdAEjZ7C3UV6R/V0/GuBN41yYv01EhzAziBHk9RNGCQ3KVg0xYckY
fIND5AlYa3yo9nIUQNP0AoLC7lk8fXPCumoHl8iK9++OaG3vJbTsSwAVJIeqJ4xuVvbR5GhUpikY
MKx7iIkik1R8PyreFhRYL3UIAYCQBU58he8KWINm55fCZgT8WK6gkh9LA3Hx2i4To6K07dgiLX6O
YM9MtOjJtCSJabSppORwWxdcuj89L3IHm0DFKk7EinBin4FQP7CtweTCANBmCm9V7XdAZrRK50mv
T7p6lLKreD62JUqHw5R6eaDEtebxkFoWiniI0sedSZ3QfiKzG/blmZgGlCDL/MIzl9map2Jh0Poj
3M2aRaNS6AVpB8suYTrGnktvSbB5IQLXE2FXanRDKTXZF37o6G/u4iVy2CWHENOjZh7Oqfbc7G0+
j+XIaYrzYgqrq7CAo7xmN9N79P7ofFE88ILTZEs7Zh3VFo788wwGRTiVHdyA7ldAQlIO2YO7JNfT
2jbkDo2eMmPlN7DWk9n4tpVVfL7KucJsiJS+sCALuhZX465u7/ZMCMqJegZjSdDZy718NmzONh8o
OD58tL3JFz31rXXcZNNxq6wUcgMteyjL2mGuQBa7Wcfqef5RVEsYJq2SUMOas5IGESo+jnb0aVc3
lmNKr/FJQ28iBhR1PmqykXAgDaxoQZ7vShEjggmMJ25W78btYBlTgeKbqwhmpk56BVQaiDdyyO1C
9gsYXyJMSY5/kdeWecOiNmWB4XEqsQk8cqsBOkYK9VnkiOmuOmFaBhjsH7Yo5NDf31Vurg93L81G
6iKnyXwNwhOfkYb/Wt03Gh9ZPbDitOlW2VMLwBGIHj4i5NdrOdSFtRAe3iercKvGoGVsMBZZsea/
o64L3qKz/8DCnGe9dTT0KdRkR97pMzgJXW7IASvZRFYedwzmSEdL4pPy5Z7JcXI47biV3dOPMESB
9BUGP00JwZpuPjcZpTh0vTZLQ2SBwp1kB8btsYANHA3ZW47ueNvSJxXIlhaj6yGhIpLb5d1qQtyz
CqnY6FnVxR8J0A8ATUORdgv4Afz6MnyyQUkk4rA7FWCi4V9beaEEJNYjyaHH7i8+FUadnvVvonCH
DCGF7BujYQGeNdrd0FyRRsMh15eZg3DkN6AvU7qtIJM0neHmPQ0JNZ3zek5vxffsVHpshUiXhyhU
5qeYUPeoOF2t7T7u/mEz9fBvhXRLmLCf3At+vWoGDdcw39BAR7bT8Jiyl5Xk/ynsgCgzmfWjn7rl
JdvS9pFfWLwymZYlg/L30ifbOTeNpiSv23fZHjpITuwq7vWNfrGbngtZIyGiMtLtQQ99/cKnUbxJ
5bshmIqxFgA/BYUHNPfTUXnCYYWAVETQh4YPzbWCCvLghA2sub1e4+6Edloho89nShUleZgAMG8m
Q7O7yX6xwqSVuhBx02LARfI/RMOPXCXkpsAna7zI4hgIwLeYmNyAPkXxd/io8tYXalLRd7aS9/JF
YRgpa6PM+oYeMVGmvkJuqHmMLGR2De4FthgBXg7/IN3vJx2Q/0v8VeuBxYie70cdV+lJs3Fs36Ag
9HkSthrCpEHiL2Hfw9ezTFaeU76um/8I7yO3hl86e/NwkUGw6+zQjjsNO1EXXzz7RkfGDi9fgF5d
j+4uWQJ7iSqCm6zOPA02+MIaTJV4nbA6YoAgQu1e8kvBBVKIsTc9AG06bFEIwrYb/ezJACEGAv2q
e977mJJ7jgH6ly0pNAfbC1P76luJ4sLClAJEwCqYlBQuEY6QbDhH35OA4Zdcfw6T/3B/axDXKhJK
yAGZdub7NnSjCVjDDiB0OpV1PaSRQFaTCK7tXlnUBEAcan4UssCi+9RpAdr5bZVhJms0b4oWewdf
biQuNBCgu1gxg9WkhzGbdVtMq466xrkaT8Si99GZbXjUurvutBltw0VZR9H6bIC6PF1webfQI0E7
8T+7dTdsAZEBWI4T6QDnvLq12vobZLkq3kaGaOuLWkrZZ3YHDWr36oRHLjua40xZmMIyJOQIsXY0
XIDAvI7BE2dL//z/DgF3g47LOrHUaTT2jGI9mcj/h/ykRX2N8u/AUqbQyHPoCTB1yXTn0MCmln3g
D0EpLXYX+Mmnsxvk5pomZTHFB4utgypcqWYcmhdhxopRH3eYliArZg6pldyEUVXqvuRIvlv+SNn0
jYeBwxKRnOyZu506mKPJwPuqSqdw7mqj6erYrwpJ/IT2r7jruVZj6lc6uXWpVbb3t/u8Ql/CqbVg
AjDWpqPhK4NGOEygenIWxBVU4k1BEp7ScslL5+wHoYYzPo+kNMPLs67PVVweo+d0y+BUG/mdipm+
G3n33AfZKe38IVWtBy4ZZPU9OQbvIkctmj4LITjUeIg27obPZfoo/xQjHnBkPFRAge1rFlavcFIp
p6abp8/bBDQ9r4L1jOAUlKuvOBNk3SZLGjPgla5Zu5O7gaBuZh0wgc7zx8sIhvFaTkNeciRchfwk
h0/vM1Qh5Hr3wnvyVLvRJGqs0iuUC5rk20FCc1ZOcwc5Nmy88Q8PNITT/5/wZ9E+m8s+I4bF+X97
69ufW6Qz6wC5RcSDCXxhASZTItfgs9+suNw/R/6MqP9FdXRKtyI9QsiPf3LORzFGWYTtKjhZxDfZ
vDbxb4RA5D1U/Y3+kdTXASWmkxd7llg8zsDPMtGcOc3f7b7DAIglEz+dV/UCIKr2B9osCAiajedH
GvI7nNYlDEhNE/IAprf2tf3LgPF85sOG3XwJ2xpjwQ+fipVtWUMyur/XnsLD3TR51nBEiLoCTjOW
qoOc0Jx7Uzam5XdBOevDwBbJP1Solj5ug2aD0J7j4kurXl0lUkPzu8KEwN+map/ZSPGuUPNwCnev
uhVyYxVrpvUTpzqHtoWBx1ipONhhElRCyZ0ZZNNryJttienW+MneY9Y1KRNzCRq1fVCmD8Iirh8A
ZRUPAiDMQZDzsvpxG38iKD0HMMeRQZpvbKczlJtdp94iUgGnprQu2XsaG3TqSuoLLpVoGNl5NEZM
/VfA3lrkfbRRNaMyyQJVxuNDPxPvd1LTRGBnMPw3MdmbTglifUTnwl3jwbqLgeQMVzqzC/L0UuSU
VOlgB640XCrIKmipSShWZAhBXwR6mMeEmkeZbvoI3o1S+MCtd98pI9T/RaaAgy03kuLmlEW4gDNC
khd1ivBxFpfG9n/5EpQ2owVLQuKK130kT607lBFJ8YxmR+sO3TZ1BmJHNr7Bbom8rk/qk1JYMXEV
C6fvl8cZdToU/v8s/piOBixjWQPeWd0RCubXrGncOhL33diSrfGwQmfUhrkkjozY61CxIa8Kan8p
UE1O0yke8JtUw3I8LNAH8cnxwgsC9kkJypXlnpU3de7K1sjihu7wvO8VZgioAiACRtGazH/DcjBV
t/OPUmYa7KsP3BJiBnIADIM3WKjaPQ26SPaZ21quCIGV6pzmIdfkRgvL4Wse6NIMuF5iwKcZH98K
NQOVTNYu/iavOKbRfAHsuUKRMmNTXgVUQcyjjIVEoDCYNKmn9R3lnkgXs14IoEkUwM3Ay7btpzn5
H1svl0uZORlYaCRKGssFIvvJyf7GMKd9Php0UVtLG820D4oR4nvYUOF7aCBOc0afAqUlO5jc9FAq
tsitJJPMW4uvTF+shP2Rr9olz0ZNaf6yhDGsBBQhO92t+ai9K9jexoBnllKV3calpbinmnGHf03n
3C1C9HKbZdBTolxQpuj9vgsFAwHhgJMHTuXLE3xn9oi15mqFyY7eRnsIXJ5ahdzBGh5EXWBrMDE4
RiGTrO79Tk6tcDSJ7WxlPKNdUuKVj/J95b3kMDWBs6uldrjgelQMQIihgOQNffn8pmeqqbjcYOgR
AgeKBe9MojkkVMJLh2UHUk4hCVwqbhs3Snw+4OYRfpxj/I1Mq5s7/uNqLhIyHZNMBTcp7L5yzVvG
ntYP8ntz9NdNdJC6xptkGcCoqYrSaNqOU8Peu1yeBpH51xeS1HfIOruM5IZZG3JRI5JDYP5i+Cfh
Wv+0uo55poAfZH54Qu2KyOnYQeNvHUjSfnZL+PWPWyXleYvJhlQLHcV2N40/Cp/0UN7jQEi/azKr
5xyRAf22AHvIwBIn6c7r8ylq4RM/gAqtyYtlPifGKv2gug6etfeVMO2fMscHv6RjxsViucnrHDKD
InO5Mht6KT98yBjL9+FPy6MGFG5Vj4m9wu7oBRTZu1lLY0jvxZGUFAcQI6VKDUzjkRKg6+WrjSCt
+IrQ4grO0+fdOMm9CEsBPK/Hr1eD09z/5xlkzmadm8T9Usf3JJ6il0G6aKrE8rMo6ydZOGRPQyw3
Bonne56tAhBtsAgd96lXFsY6YG3m5Ut7UCRPpOZPYo2H5n7SacCviYkA5c4jwFdq41s2aa95vDno
CsxgfzQj+OABnlOj1t32nDYyZHwxE+n3fySJ4w9KpIxL0QMyhlCvqoAeqI2GOpA4BHzQgZadlY1m
Dpwe5wpbk/s+Bb1tVyxTlxZawoi80oNTkd8BD34gcXZWQtRJC8gxqR3vLp5VLM+JV5D7mmzVd+IZ
gO60DaCGDuYEF0hHN75ywPzWRIsbJL/IxrX1GXXaU+5BL2pG/cZyQbJckANF+QttnhjVev78u1lu
ICeQ3nAYCGGAZ3JCP1Ipw3hRCFhAJZuevDxN33kTusSOt0/fj5xuiFjod2e0ailLChFa0PIv9X7W
lKu6UFR/Lk9If5G9FOr7eJdg6hR8LbxeD3NL+hZWFavGpa8oj1UHg6XyhcLLHjHUgym9mnORXQ7Z
AK/4WBUMNr6Ld6B4Ollyxd7mxuskHVbCT44rWVBLLL/ZU1TXWQi9N5kqgUAzOOkqwK23jiePDKF8
RIiVRNHDyCFAxuHhx0tg99gCIxMI9lS+1IB9U8xsaGbaXf8Wf9/oGbP5Bs41KWBeIaYOn7psotz3
fXqSPQkedYIC8++CxZ8pTIY2PAIctJ3Ol3Oq80cxeU4bhamRPLDSQKPiNB4UYbtkU0/IH61LG24R
irqqBOpS67TT+Runc0jnNj8RsxqKbGVknuNC+COlSevL4V9LvSXOA2+XJxcwYv9Ant4a7dfVsguX
JpBu4aG641aDe2/fU72J/rYryWbHXhFJ/pBmcR8VeusjLE9IULWEttOUIPI/xWBUv0M5bg1khIBc
lS1eLseDqcSElPHJ8rjX3NoY7by9udCiDDKJlx1FDKeprtucpoangUdJ78v+RI9eCxWWUW3W7Q/p
YQxAAFKZqM6bw11LV/mD9Vnb0pjTUjyDFCgLU5V9o45eSzZNZ3tAd5fsFfrX6e5E46opfBT4LqYF
wXqlBE7dW2vze2IfoNhuxin5u3se+n90SH8sPRBOYxA0eHIDKerfaq2OTKbslNFRnviPhR6sQSWe
aDlzwc0buAM/WKnoGCv5k5SGSefYMIsrp3TBo7Xtaqawlk7c10b67chKx4MuMBgJh1VsyEhPy6rP
yyOyADUVQv5SFbEfnGvE+E015O/x0xVby1rZ+/4DbkDS8GNTpTpR8ZlGAZeGXom8mn2RiKt5oLp2
EiWyRG8lyN9qhTXO0obws/n1WA4iYdU36qXerWl7jDx/QS8cKOE+MePsV93N/LZ/W8W3ZBz1NkkT
ulo/j37axAb+1Sr7msMFw2PjU4jjnthxKpAeSMxxJ9uyhKZblzlpN+IH1XHpxrkJoZ1MZ8uRBGFY
x8rQ9IDfw3Rrt58a8k3/Ob88gYC0vu6hDL2+AImMzv+FIiU2SjpkIvHAvL4ewNDSwO885LqfTEeU
RBk0otcZr2vLgTgYqBsO3YdxATuhVdG35vgubQCcd1mSLI/u0QmWMEkANGwnxhtzkIbA8A9SG+BL
WccolopL32k/U/eNYU5rQUoIrfetGM8rW+Oc0yyG5SlSOgS16d73VY8zN25dlNUYENeRZ+G9/UU0
F0rR3eb7kHKgYASxkaYk2+k/8M5m/gYWwKuOSKY0zC0RI7egmaqkvMDBMhYlTx/U2epgRq0zcG6h
5V5oKivIrjTnG1SVJND9Lgkb6WsNi7CNRamSH0i44mWPxsU0FIDsvNZT37OYl7IF/435gCjonsHk
vKqDksM/eZF++NmF7khti+fejURV/uoJXmI9nEItEWXSe98FwarkKcCPQA/MVb6vEldXgeoS1lM+
xCDOIJJGG+OpEaM1RhnLDITv281oLTbrC9Z4v1UxW9hX5+9188j6Ko2ZxHHkx3mw99fo3J8KA8gl
S5j0dtCZU7MufeAmOa+Oh8Xaa8NkshKRegYgiAqMXDqNbauiRIGC3GgVaD1RKVtLu3EkcslQn0Gu
u4R44NhojHLHxIZSRwRiqH9IHK2ZfwKT7jcp6wgiwrsm0Fn+Zu+U83GVgORffi3dYkgY63NzYFLS
t+BBuBp1YiE8Xql8n1PK+u11xhKDfVJs8qiRKcw15YlLyq3lV2baZIiPMUEVMjGRfINnb207UJgO
bizBUTXdQXFYjW59mpyBLREzAm+NvXLHVnc+C7MjcumQAaoj7fP7UkaKtaShSW7dJ3NAyrTKhFfP
IObVxmUsEvJFGrLiPjb3vG5icN529frzAgwOuvJOrId7n/i2TmZ4E3TZzoUx47iI3VKLOfFK6ewv
vXmg20RcmvjO6xvk1ntPxKIowxg3SWk30YOaQggAeMheQJBE0COJnRmebCtdsCrOjjCCNf629PDL
szh/C6omJOuo9tl/jab4gqGMEYqXF2XhJHsxzvrZKtgptNtg88A+xkBT0OfTOdN0yrkoomJ4/Obf
ig3QgB53scDP0Lfjnukr+IjYb4ixnIywJyLP7ig+uAZpYEmrrSX0JQUeLT9EtThaUtkUEuj4ritq
3Vc9owoOwcT1U3N3aNzm0iGqcL5XPu35RGkbueecK/3MqVXqmMhk7kH9hrnXJ4j1ZC4oFYIRYLjb
1Ms5qZfuW0wPYlPaZnnEOej6oo0rscHRUcunlJtBe9STJMQjTgw5lpKk3LLiL8a4PznfC6LTyAFI
AjPamsypbKEZQvnItQWe+QVYBXexziaH36bozlyJcnV0MMCqU16L4Zv7K3K76PkkiTH3fd1qQd96
AI1xPxCft597y81vE0k8hsrN8HIiEsJ1i9neFIXQzWIOUBl7SVT06B9o6x0fvOxSriQLeDizQBm1
8NpiqB3txwm8YBSrwUxBaoXGtMi7+UG8BB/apcZ44vCW4eoWFiIoQkHIRD/wQ5wcO1izC0mycyDH
TRv0A4u39omw/G6tiGOO1Iu6FNNoBwu9U3rHVMcRF8ILpfBt+VFdXsF/rGLM9/dKGzjbQnnm2oWk
BAcGbcKyGggktvCvB4aNF34k7YoDCaxS09eQiuXXirU2Hq7am5DE2suyLosDQ85svUcfYuhYeoLH
6Njjrs2DHqIG+wYKJtZMKsdtf53XaPMldv6loTmJvsKHeWG/VJ13BaAn0pZHwX8PqxgrdoY1rg1M
3WAroQPFGu3JTcoeQ13hSnRvZL8Dr+FvRl0utba0OhAgvoeKfd50kjqBigjE5kKLexKyEU2DKDZs
0wicPBHW7gzaCgSZGoZOSvKnP/4RJ5U59YzK12qo3LlU6XRKf5hfeZKpnGgs4rAWxewKKUVoYwO+
biOjN0L0SDr3ky4XBGCwMC3MMenFTNIlxlnsftkpuagwGAHBMUrQoeoO98xr+VsrNuChjVK/qJ2+
tJGX1aP0vXpQF8cZwZF3L3EbSDGvwLaeKjjlEzEYDQHNSb8rDyHcAqnBm49IdIdqT/ObaJvH4Wmo
gjCdzkiLVaLj5beADeYFU4vwUZKGqC+aLMoZChLxEwno/kk3IZL9raZH/oQi2ymmexLESrWjCDuI
AGxdDCSVFiSnnGmbRxbS7CXlJOAjPqvGIFGEtfa8Nf/FyIIdY1AQvFugKD6//RxiotNYx9P5UjeZ
/3vpso+Lsso+BzcqKiPg5KFqXDSxmNgVjQkHFNZ2DR0dQ+O9HacGt4UfruSOvThb8tSM3bEYj1OW
SHqbd1vZqlJqGbdvbj6k9VQD2FdU/wpEHIObEpmQ+vKqIuBgunTZySRSxjcdR8DXv1if4/8eDzwM
SnJ9lgF5wRe/yJmHlgnZ4UrLnxyv6jVxSCNYSeXaAgAkne+FsGNbH8mNuX8clewYX+BMjHJ98JFl
iIUFHgiRLti+QjQLZaeut3hY+B4yJA3URATysgVlD9mYAnEHFpDSsOawHfX89YwpIWb8lrI/XYg0
g90a6WwbRJPPHdGsQEFp9IEyy4rkbMl1qGV63rcgp10feDIb+4qt3XI4Kq14jV+gHtrYxI1c7rfE
Rqh7QVQLZ/wTSEx+Syl6rs4u71zN2TOT0zR23Mou6Lm4rSXFXEt18MX3jXm9gudXDqvAPM9N5zp2
3ashIlg7LaGwgVuas7l8A1/K5liEUB3k4SLgmTReuited0wIzCoTFsblyPt9d6xZ4Uls0RRsF2Ce
5VR6LvBq+M5umOJofvzsh7c1XrgmTLgkwF1qdeQ9pGQp6ds8O1V2v39l5B02NEmYegTBe3tAeavr
tGV4VOr6NW2frPlLpNOFVVZzTVV/iDvSukrGbUVlJyEsz1qiASa8KFMY/BjX9du1PkKybL6vzNGe
BJyS68xxqnNQjMZQMEAZ/PEy5wfKFnDSgtJx1zxL+vfTURRIAjp0df5EPQmEmFHnI1+JN/b1yIE9
ZZUDOMzG1kLEy3zRvgJG7g4ZmM/1iZ5oQYJnIxmw+cxDjgOIlpMw4+OWUr+PPlh0RD8YScJLsp+9
H5SFTcb0sN46EJwwKVfiiS0Uuz91v8bIxGE5wd5SCtG8lOzcbR/Dn+5ukqJUk6MkN+ins19YOHWe
yG8n3hinWgDXmLjK9Id8zO6Dgs+ujGUsyxdLeNulYKh7cGOvG66dZFObnsjw1O0+DE9en4KPrNd1
3yGFHAV8CxoGeWlaSUucZ3dzHGfVkzmlYG4+xZz/C/QwLW1Jg/J9groebaj4r3yngyRvaQhk9nD1
0SbIZ6WlkUlppOrPJyu/vTb3gi9uQ19Fk8U7nBFBQdzM/NJDNmY8x7jkGCiCLLFyAHIEvuR8wCJD
D+YHk2pRi/rtSyMR1GkF7FmEpRV9qWFv97OL3CECntFBoHgyE0nP9CbSrgwz0LwRndt2UA/FGl8k
TcoN/xTSwCChccBP0jGSRTOgSoLtKz9rITr5GzONBWLPeGz16vZ0NaiIngFrweT5HVWKVg9o50gP
eLW1kA/XIRzvzVE62NDT8Em5xMUuMzMLsBEymWFhTel0kpScl+Z4oQBkup9/66lQHY0POKuDWF66
NiV0kq3Kn650ovqDt3LQU2VDlgqYJi6K6ipwP3siuvbvsMF1tb03Wg/LMOUhsR5rrOwkbPbpSqZg
VRChkyDbtkvvpk+HWrOzvclkOBvRThyprKPe3GIotF02U690vKpE6y9L+N9cwWzn/H1uzgR8xeTc
GdVStFqXosgkQiDtGOu3adTrfVGNsp8mYdHseM+NEYTMrzTEwzR3/xq9UUiB4O3OD47JN9TCNnVh
T7zaMcgjBanNjc0MDdq3bQ15LK6PKWGfF4VlON0gsuXEJKr5O1PsBjcZ87UQpjHa+ryfNqhefjFP
pI8HqDL9uKogkqRpPanpYSZ3idN0pQesC0UsU2TWByFXSymTILg08J81XJaTZYiFLVYgr51919oH
M8XWBKXPt+MR6jhwMBjmT2atV1zSyZ5NJg/uySlx6kZnwjbmJmkC97IAA9dfqPHertFuJ+nyxLvy
1AW0Syw8tOs7iErPASsUo04FzMXz36uK/hw1D4lS8cfoXlUxR3sDQM87LvWVjG+dqbNsDzlq4zsk
ZZaiVga2KHpNKNdunAlnwNw3DkiYME6romv9CZvtuD6pAn5D9TaMcHmfg6hD921k5LJw41ZCWwwR
UqyccT9vmKZnCD5FeFHUkbW2HPjUwp1/I6gVTzKStORoJRt1r/s8jsJKrhH6rNgLrWI6pa5uujgW
1Ra72Is1m24M2kRAde3Q9YK0cgZ0Mumbn6cDgPTdgUABb4jYUfzxrONkH6jvuKylMMmiafisVRdM
pBdZumc76qNoEcPr0nEJZWgE0qa81FMPLyJJ6bqQpnwEz7wtPxaiiDj6S1iDGXm4LNBU1uckXkSI
dz9kCGPI4CpO6x5tLzW8N1MsbX7a+1RUmJVgrWPpOc3bkygMdNXINuuQPkjIL7gpI+m5/6rSs8Zb
S7jTQwKjlbnfns9s3Z7gX1Yq0hiPj6u7szxr4m+nn9yFO3ZCyjcNBc5a9VqmT1hEO2X+VelkkOiO
nZTYKhPNrwf3pJdoTjla9PebZLHBaRZWNGCDMKITWCqenTTfPgtO7K8aC9taxLzZkfNGsVePDUZE
Hj/y0k2zI6KZL6gROdneqbmbNQkT/b7n9eL6c7Gdc/MemC0FXsKVH7FCQJD3R4hWWBUnbWBeZfF+
0xE0Ot7t04W1voapj2FCStwvsElBtGKgf8EZY/3SXYBHD+Y90P5Sov5cpa2SzfOsQimF7rT/VC20
DV63RNfYxeepSRoLw16FHnmOHzfqeNv0jOBTJKJvDBDC9TrrL5QNIaszFH8aoRSn6dc5bfZ+MAjQ
n7GFr0mFz9fFAoiGHaUoTyrmJKB/rFJxyecdY4Y7WKUTyEGPRR8uP+En5pbAMVPvqXXDD+TriZN7
o58Bkh1FWeCjGIIxXEpMoIYYevioCN/mGX7cX/nnmWxvL7hgt7ms6RKH7VZ+Sz9pFuBuLkHjNueq
jrfwhImIJK0z4CyQA+8hrsjEvZ0imvQeQdqmjGCJCpXjWku4i5dJ81zlp7qwxK7w/co5uVZ4wM/r
MxUFC10mPAFO2gCsbEDHbuaOHWNCLgcyhr5vF1QTbAWVoHhpwmpKmP9Hp0EFIZA0ecGwjbG+lfJN
B33vWcnfWoTVC9vazOs3qtOQ5D1t3V1Fs4JgeoVyYKb25hhPtw3Dveb8rDhVghNsxxq9VkB/wgwq
l5eNBn4gQXhg5XXqlIQClyn3aOJvrjEvJ3Wg/lV0XoUPWNF8yIx2roUjnwgh7Fc1xDYO4iF5dv8Z
gPnCWPVChYbcV+g/Qm4at/JjyUH/13+efkvylP24nvADZd9rQMzBeL7laV5z6JhqxpFq/UpTJqiE
wIhUu6bgx3NnVYYMhC2KoJ4bRGl2TAiaeYuyXc7VIjqLmitamR1EXMay1mYztnuug6DjWr6xfCZY
yjTakkrxR72DwCXPQAowCDUWEADKDN4oOId6HsBFu7L+xRtGOE6hQ/sEf0MExDjueCyGPSTqsuqZ
mNY7QkD+k9z4JY/KPswt5jRf4F/duhKnlX+9cd1UaaWO142+FQqrKi71OMjv9ARD04gRYnbv9OuK
1J+iQGTg2+CdtMLNspxygszQOWnPckJfFUK15aGGgu89k3X1Hhlojr0+j5mmwxgDFBO3bHq5+ok/
co63U/6pFJ6ARc+oKNXMNCYxjiLktRxqtdD3dXFdd1+0oStyS1qTS6ob/+k52Gn71DVrMnGuDrcW
7dyCplYKnt9mah4iGK6aEiJ2WWMpM/whj7ypbseaMJhorUi7QZxm0w3bpDIbosiCGZZD18F6iHNn
N4FPVE95LB7W7jcAyeOWL12oPN/28gD1PV1a72oxdtYFhEsOwCEKq2W6tPSjNZquI4lJAF0fzYCH
LXR5UmQXGO7n90eUHTbvMiYgrHaSkf/+yCrC3vdzAfY8CbhG9klqlFxHX4GYUAPuG/nzKUHebGHZ
a/TCfi6Omn4ZmQg6pGJBjAJUmkchtz+OJDCmE48NQsFJQGCwA+608pgtrJhCUmMdGWKYm8A0/lsi
GTPMw2TLYUHom4Bk6CQSOr5lwN0Fy3e6Kkmge57XA+/jPYbhbKRQMMI7QUW9xPbOk8adg1IlqUEf
rX2lCOxtzrI5yuN8pIGwe8qxL5XDTCPyVi6TWlprd/98/jC/e8PXs/AWJJ47EXcU2NnUTEZeaePU
8JF054BLfaswjkQFgxdXVkVE6CyMV0k6YNkfAaaO8sCMVr0SNNv9S+YjCrrtwcK++Ox7Hiny2xEf
AFSHC8BwfTEX4AJBLBKp3MWDp+K2y8AitwhL5podDm989oldv3Xa1PRVThfxMW/ZIOLQ+RzGMCBZ
77TUxNv0xZmBad2eVW16tIiJJfZjqQn67fp8kfaTGnKeYLa6xJ9hApbBNxa5eFyoXBfkXLStEuG1
DFkYFKoD+ytXvPZ2lJL6KpwFrVCTEtjXvGvgDTjKlOg41F5C2XuxA3R5zOm2n9S3OQ5slwreEF6E
WoGvMR/+N7Ii7IWpWDZKxlu4l+2fxn+AHH10l2POK84PpuKk2bvmFs+NTlMzu3wmUJCESQ7PRLIv
1IYOoSchkmZKNts5AkVmDBuT6PLbcUldWPyA9ds3pP+c4AJ5w6nVO3hmgZrHFgu5Ag8s92K7ygIK
oJLeBB29/wmL2jl0j4nQ1Ds1pwRcgtS4F4l9pMu7eoMYltUAzVDtnDnwfZt6Y4qYvjrATNdhLvya
vnqqFJtfEvNBH9KGOEtn46W7WxPvtyb3IpeZzB0cx/4znmRg0WOLcjXYoeSebNbyJQinmY6WTM+k
tFwlartI5ywLmqMCRDekHvThNQtgfQsFfsO2wEuR0KEl5zbNvOT1QkdLBUKTqWgHcFq9RVE8Llj3
qU8ocXFE/fthXtfX327kQTPL8+QB+7rNs8lPnTixKvrnL2OhCDVBXqDmvSs7TW6piMA65h5Iva5m
snttJSpcbih5wjDeHW9S3zG94XbdUq8O2Iq1cTVaRfAev+iMDtQaKB9fM06bKhOQnOWGoFLStObi
Uumg0nXE6AUQwisXKG6QvyaZu/wuk5YdU+XZAAKpSrrza55oHYvlUMDRCwXiK18JgBtYngv1nQia
HyamGCoS9865wznrWbgMuXqbtOTpAilLIoZs+iVT5u8kttDRS1t3XqyH94LZt+G+0h43/CiakdGk
V+ORUDec1ncxHgwO5NQMoqoe0I7hqNFScrLYxzxquPb0Zj456VJY8rAoyQnoCkYjVhQkn4k3G+Eu
f4AKLAAPuMGlsEEv7jKUyxCMkNDp8djBHInqpondInoPCxQWP69U8XThgMp9IHnVjqWNkD6QPfZx
5RphgssApF9D1eyv4v1c6/Mknu2xj9kehKxwKQ18HWVDwYF+fnUACtwYCQveqEI+FOUr1u85820J
wXHToKEwMwesNypO6A3YCs/a3yRcdyxSQNZaS8TShwv+Eg8cTvTY8XSmde/bAN7Rrk4Q9Dr0Xe0H
DOt0nUx6SHW9qw7XjMW/c4yvDTo2pSy7hOcJaB2CKoxJMzStvCD1+VTkqXTTKLC3wA4MeltRv2Nh
l+JRug8uk4jEEJsoIwAp3YuOQ4cFshG9CyDCVWuSSdSUsBhnq8pViJtgIjzcPkQ6LwdjREGdUzyc
jSSYJKIVxiwOX/3G2Or4pvFWO7oFPnms5RnIPP+RDC2ZpqWrLXzwXeSS1rLBDxkqjNOCxPRzE9JR
AIGM/yVbQRY0ZeNmh+XUldgDp2LKBoSlEN01BPPHXBVB37il3kTLAPk0UspkTv38qAiDghhYT8y2
ivtEbTyI6uPP1CfZbnd+szGcviggZ08/tqz3omct1LTFNoPSVmAmjZL93rsewBzZ+CewsQZqQKAY
418JdRbxxQJ6zLGjdLIPckMhNtsMaN88ZXv3OGduodba3Lpr4RcYkKuSB5aweW44lUQai0Ed1WpY
Ii7s1F2k1+49ICFUk8rQgtLEXjAEuTysbxic48otPP5/DmTqweWOEGrhtaohie0H2vL2GS0a8hJ8
xlMe62e9pXJ49wNOZ7biS/ik+PtOgh/hrtyKUKYyZOn0CS/0BxA5c7ZZ5LyvEOrVChNFNq6dcRuV
v5IstSfi4HpHQiTVLdEmKIk9za/MB2B7NhAkvWwDpaQLpfvvjFtcem2pXdyyXQ/bHPQUEGSNnLoT
V2aVrrG7YYn250FGY4XnL5y6kY8WOtBnYg/mgdPDwqQf6zPhjKb4I0cIJNrPpagZ4MBO5UN1wJkY
SsN+3Nmp4hHBownc8pWtN6sgUROclknyLF1T1Qrcz/dKLJF99zlWi5EKDpAe4Wuk7fwxCJkqerSM
KeTWPWxwLR3GHfD/G0t08IPOflKD7XofvAyhfoIaMKuU9TMaQvVYbh88x73Pl755fzg2pv2K/47U
95UzyOTUda+FOq76rAsBbnXeoWGZ7yNe/lUD2/eK7+eG2LzybrObyDs11M0Dtyjd8Adfo0mO1tfV
uP1IwsexTIBZ1x7HNqsC6wACHnN62zPL/LhhQPIcjL1majS6zue9YZvuhU6tAmcHHto8rh5DQTRd
0XfsvSi6LuatlrGTkB4DZUVXWkImysEI62aH1D03KomO0kDiBo8+Uj/bOQw172Kaj9XXNVo+xwWo
cRtsmgbYuDwD4CmjvvJCzUp0k6YpzAy1sKozV/zo9tLCSUliay2ee7S1vEiQzk6ttGothu64VgDY
TJQvVgXflEUjh1Jnti+14j4eyyulOdpuz7o/zo25QAxye+JqVvLzJf84c5H4yUs64B0NB+YDQd2f
3kH7NHLNXFfkWbVJpjqXeI4AAXh8MIyzMBcWCgEe2xyoJzbAD5wFMXr7ogWZZGcqLJaSruXCa/Nj
VF3kuM7wErs778fh+BLdul95r4PMW3IbWV7prHclEoI9kep6EPQ3W5gWS6g6WDdLnFSmlqWO4Ux3
WhItZo7R48fzSi8nGUDtlvL4SrmNFa25g7mUEp5qz2TpR5bjZbnacK4tYafrOcS1oXruJEU3oZP+
Nq7As8rkmJKi6+pE+lxDotCqcmcwVH/WModm7hFRmb5XtI7TlholeSzNiYuiSGERw9athdUnY4js
n7v9WzJnvEGvk7njs5eMrVDH0vMuI0zeVZmMpHQP21HOJqE48IguX5OFlAfPxzBCuJCUhjT01aFc
vagGlnJdDY3jF9TzvhPBL6mLmyFOAtjw1t9IxYzaIY1W/2490Cve+8P3nfvRu5IDNEZdHEkZ6Sqj
bm75M60NqlozZcHY7x/WMg3DVjdUDddDyGKfKRutzwaqY+JWE593qDejYkewehBszikuB/xfMGr9
3y1dLEqKcDS51y1vowEwRSOTg5I8FS9r1qvgs1TZLJK9pnKFUw5Wte9mNSMZsEW5Udzw3VbcF7js
NCA/cEJnCYjiVhD5m/FaE5fJbVtc/Mq5VZdHv7k4REMMhZ/mzbJzYdvNv4NutD5Jo3oddxuL0Uzw
4fubyEawP4Oy1vmS8fSc3XNByLuuv7WpMFCWM8nhSToz9fTy3S5GshOEdHEqnbqCp5LAoGys/sCN
fVo0gfm75pLv8A858kajbIiiGimvZAB4uBR9uVlv+OvE+5NQyKI0YQ1SJ6fBsQf6+6kp86rIaL9i
AKcjPWS1TyUbD6CjXmmWjD31NgudyJXlu1qyop4hXCk4paecKkWjUZ0wO6IvztJDrFtBTrvvA+DA
rJh+yOK0d4zGzA3eTaQUdHdlt8ln5h7U9jP6EfbB45YLH9qymtFZURdhUKKIFs4dmQeC6Nd40R6r
cKwwT4Oz46FRheUsBaUqTbLIP+5eJ68gqu0pIDGbI0AlulHEDoaH4eQ5r1cUclfK+zYAnI0qjQi8
iq4KHDthEn5/SCjaYgeVcqPm6MWXWJLFNa9JpsvnOl2ZfEjqxpBKtxP/ta5xghQ6ivCojxJWMo9d
cUztbt41F9zMTbOZbhZ5DJ94TT+t88IpX36K5TAm2xuiG0MinBJ57O3nn9xee47pxmydGH3/abmV
uw5CBObVKjNbyDtga9X/3mFb8MaVkxuc15VeaZSnJF4w6TI3LJbj4II9+TlqkXL31xppTGG7LgSG
yT5SWtdGnC8WZ/6i9dB1dmnSXFj0LpA+ybDFpOPztySArmBGYX50kkyi3Ut2gpUaQ01QtWzXAqoc
PwUBO59d2v1Vsy5BcqSYkVSDlRM2P6mNb5sLQJJ960Lue++z3yPQH/cRx10GfuLBLlDkJgcF+q66
oDed60VLGEOXhvc95by4MDTWXamBEDGI4dEbO9WMEQXr95h0jG5x8cSGKIHJ5UzlE+zt0+isz3nf
VD0720O0457O1y2AOTYRSrXFXXrDU+grloDCdNgS8QJsqafOB5cTh5z6jw3DL1K7g5pKWV0y8I3X
Ir1DbDS3fCFS41afo8DOoPOiwTLkfapL5xGCiyVh2fWqNadg0goPk0qf+u0C6afAn+uKAuHX42i+
wq7rS1Y3ykEuNFc/f0G12qIOJjhFdSkLFx2IVS87mbxM1rjCzToMxjueIsnhpaBF3xoN/GhkB2hr
ttV82RzyYCgzsvGfZh/MGHaLTU2VvvCHAr6oYWWMp/7Ps6uv98jfoSOt5sh7w3z+2sxQ1TIWSyPN
JC1hCRaIDQPXCcVepobmuSshG4fWDtot2voQjGAMiKj+FleUqStIAP7WZW2cxTgqEP/8daiF2btP
hW19sZoXFNBL52jJrVA4Ia1WjF0XCuHhjWWWftbXQrEhAoLZuiPM1ymH3mDWURA0jADQIak/OXMD
xzMGek2amUvAHIhqk25S4QpFMrntNnNvwDRc3rf/GZcPy7SZ+afHRRrvm4TINjaA1nbIlEBIBn53
1QdpkTlbEBKH4zpZhkeqM132pcJPiUkBphmseprZ6GwqBqwur1EhIDM97d9zzOh+JKSQitT5lHC3
CPWqUUEke1bVOJnIJE/+2j9cVIoxz/TdGcq8shpEddPGkxr4cTURu0R5jOH9ZFizJP+Heq+biTJC
gXAWSMIAavSub2gwniTehkN1E/ro0Mr551r/0G8C2CaPfYmisBAoTovcArIdpsHi62FjAmjnPDyR
LmubJk+OsmWHhR3xl0SuO7olZxe2BhlzYdCzVTBeY7ZalXaUW5oCDMCj7l3TbFdxuDUVI2e6hGMA
K4wVIjtaXmXufylufRKrfyCCnEiLjZjeHlYIFYKL5bj4edyWViX+ik6f6i2v6lxA1bYsaRimI6nr
gXcJxbVFdr10AQ0EArhrSi9cYtL1Om8pvmCTukjrahXRuCGHvhuvgRFxHv7VHztB8xxaugseuZEl
Nb8KD0W97fVuOgXlgOeJxfvA6OtCclh0JvaW0Wmr3qTR61GLDE9Wvxb9mblWCOeA685AgrLWdpIv
gZE9EhM42GHumeQXt70qs0bBkq3unFr53JTyj8MN8GC4bI7A/SJGCtShmxD4G1pP09l3jSuWyoPS
O0y22t46U/x74mnNPhC3uTckk3/9Xd3JrmzGAR5kUWloNAXx0WjGU4cWZIXRJBY2AoD5pdsPiFZ/
+tfAC3Ybmd6fLdoykhNXJ0rnci/ce40mrmFXB3Uo4v7gDSJ3nCgLkRO4sgjXYPs364NefDtl0a8e
oC7G8R44FeDMRF8o3NR8+NyE9wxj82E6DYM8GIyyvd5z6BKvcUGVriy3qS5k3fiU31NEsesHUnlh
DTgIlnAMEZzp+mHiBtmBoXk0orXhVZHu5RwK3emtDanVESb2SCWiAuJIO6X0XLFPYoUQC0FbJpsx
eXhVRPMd0a6TuEBXjzL7XwAYpZom3voiVUJMrpd2+jtSmy+xmFxDksGB3IjtceVQdDgf52xs9wXm
oSxFk5lQIFSbZ8ppGTnOoOcVuszYWihCgKuvZYdLiB9jJEKJk2Gs/PWJ6E8NFz0yHKSEYUzv4WAt
DPsPj3wGM92wN9P0dlBOt7IdW7BWzoi3ADd+9S1CY0u7XPWJihjxHpAB5Qm9i41+C4K03toEl9MC
Kh+/sTUt5BRk+4fuDA3X7b0g4gpUwwqFqpSzULq6U4wvXY4p6KgE9kolYk3aC5xOSButL/CG8PXe
Tj4ti10fl7NEB3vWAvorHlG3B1xx4+mRVp45s5HBnM2vbSb7EvzgqlnD9sb5JmlnQW5JIwFZD1MR
/RhryX3L+bSDxL9m4pIe91ggzAeOYtbmaWqVyu7aorO5qjoNInoIgGMKtT9atPM0eIOtrOOCtamv
EfsCBzh/DW/SP8C4Z62i2a5WumHTnLolJ4vHjq9xxIfLQxwrYQNt935bNhHia3C3NENDataLPqYJ
wucjvqeXBJJjwkYiSjgb0q/TGCNKFmvklWB6pi4Dq+rlcJRaTx9UtuIP9oJ6pfh88jnI9i32oN6D
abCUNNLcdoZeIf+VSzj1UcfS4CPHcwKNpziOJgeQJzTv5gr3ddiHXKm/Iquho8NXMCMVOGzKjR3C
6WqTatmPgl62SXMe9IKmzBanOBhUuRdEShwl2gpZy9TzY5IWg93zyAfAVbOPwoz8dM16+t6WpXDR
ErAFbzZBbDu1Hs+kAfmWlHjJ4XX1BEbFOUuYuq/9AIVwnf0iHOlXURUsvviP5bSzsch65xkZx/C/
uggKaC5rlMiLgENieIYKamPBMljBJHPjzu9SGHUwe/3Xs9Xar2NLQ1KSadcovl2mNLxBwxdzrDdC
AFrguLvlNAc+MsbO05SbgkJGzQuKzLtwteUCNy2A0t2ujjiu/vP9vRYp57zoR3jkqohnQ930nf/O
6gJCPSNWyusDHhe8D8gGe2/ItLRBpeUZrnKOU3zlAS82+LmqJouCmwLgVvDaohny3Fifqa27aONx
/c/lEswe4SlSiJKqP1FJE5JXivYq32V03uETp+mB5MkQWGwp6n9LEpKhbUsK2YDaDc/xiNMsziio
YeNX8DnRgaqhbjcYXMfJ1gY6rlWHbUygvKqpczcTnvGZMJuaRmxD743axuh76wFC7fp9O4KNV2qS
AmK2iD1xD7AnviDkH9CAoeEDs5Yr0aNTo+OpfurX/bRFMiNokSuFUsGZbpYDnwDtEVJFbNHh5Iwq
HBTHo01on2hxNjmZMI74bHt80Ese4H6wCKWmE1bNdPLvUlhwQl/xQyPHyRrg7LtDewyguMzSIHSQ
zjDdfFuHFjLIfFReLP4QnD/veGFvGmKggBxofbmI1i6rj1q4/yLDv3Ob6Xmszh7M3IyYzcAHxNd2
wmCQ9KzOzIZEJaabPSXQ0xJCshwYZMDeRaG9UwtbnkHoNnmNSkRCVuo9iapVL/eUBQ+4+L5+BuOZ
hERfOJkqzIvSGEMvL/q0J0NjtLjuqB+3BwNVxLirRCMhcibaCIaFV176FSr6IHRAgQeHpVIAcWYc
93RNp3+C3blXXGDBvpXeATvFL+VquFYQBaORY8RQUi16Xy1+gCxB1LbZxoaefw/rgU33H/2RzYhc
f/GLGxj655LptMd8r1OVYQ+dpOH1X58bWQSxccv99eMe9QcKl1Z8W0/kksPt1ACScgdDdulN09uL
q2p1dhfDQlzq0x3CRdj/evKXo3NOhW9+Ha1M1wTkyo3zj7fFB0HFDDtYe6nasZF+5kP06GosZbB2
qHwWRVQQ/lYTTsvnKIjYp0cTyYynK2NjtWn+/TIQa9XV0zAu70RhiNncabGmXmW+M/nQHqTHbhNZ
kdB62kKe54BVrBGPIIFkqmikDhSzTXA4M2Rl7zaVQ3ixHNl8oub6KhaeilOD5WcJAtFd7prTNJCf
on2Tx3sh6dXKtARg7Lq6dkWJ6iZj6w8UVBqXbDJCvdYjkPbYPkTnEy8jK+fTQXozrRIFucO7ofsz
7CZHhkBIeIqj9q7beeFrOcrWKfphGIRG+xHDcdtonEPqRk1V6v03k78EF/rqRBygDi2TF8DVdwcC
Xz5s3e4B9DzTra7A8GO+MPpHn032sGOcbxqH/FdQ2YK5s/1jsuL9iW9CqEraXYtTeXfblUr7a7M+
PZxqtz8Ke6WjfslK2Dt8w0t9T5OFW7YUadzzpOhqdJfczpbJYVVuVTEtM+waxBP9cenGX7fRvnFs
2D+ARIM4k51gmayFXohcdHhUDOl/cBb5Er3WXH/72+dU/2S72zw24IXpgCoKBIyGWanAyvXerjX8
2ukMmQslEAIbF80KbpLSqf/TkwuFlT47+v2Gefh3Q7ndsrkxRW1DW/gZhqeVSHbI0zYp7vuoLwZe
uRr8AUSlEiByszMLfaEnLoYt3NyseDWuHSkkmJuvXGVDPYENHqlFGR7IMs2stn0NxBA+deqX9Gyf
hUY8BfvS+QeBDxPE1jR9eEmFcjzzw47eXgySOxEKHfGw3dpDMAGDLmcmu8gJncImQP0Gzi214+V2
9gx6tDKaaMcMCRdxTuCl+FLnkhBhZO5XW4RKhHhzvPoLvfJBgp/YTNrB9PvnX/QrnyLdr9qob4fJ
5nqHF4XDHITip41L8UC9z3DbcagbK/6GX1l08MjcmMBGauLibcgcnZ/3+Wp++q4lIKF/k5kUT8UZ
mknmfPH6GQ1Et61e7rqiLRcMWsm69t19Q8xYdHC5ItJci6MgLt/Kk/pHTXlJtH5JBQrqMGnKWMwr
/3xKehtzVnQrP0DzQXg53yqUxDiJW4dbMUpxYT+MoJ9K2VwBRXSWnm2u0+dvRfYwG4TJd6GHokH/
6ZIlH+moeOi4RtlbOSxqzPEVOFMBt+owMCNcHmyWWw21ZU2P7YQc+aw6XHk8Ctd47kAUxew2bAJK
YndH0sHuEN7AoSmCclkGKZ7JAJgGHKqQPLFak9Cs0J+AvzcFM+UzV/F+KHZ+TEwVi5ONjsRyhYZw
A4CpiIBMt9pbp+3W2+uNRhwsMRfOW0rutQiLOQzGSq5g5e0ry986pCp3dZ7UMlZPJvrb64VhzrAE
FY57MqJ8E+96rwPcf+QXoYMD2c0VQ+JhGjK7vj3K+h7po/WUQokMNjp3HpqMVmdMCk9Z3x7cVKCW
DRy2VUZQJePiUpT/P7qTl6Pm/pi1Z5BxghqDE9K2Sgzdkd+Q/YsPx85rYiBLkGYldR50ImTT+bt1
GIyr2EfCzAXxGfGE7k7y0giO0t9JZY7mh4VH83qrBnnLgbi67wEHzHJ3umjyeOWIdmqUR0OFZmFY
vxQAdcbRoEKcQtxpFhQiT7R1elKW6VyGe6VEKucjss6sJylGCovDR5Wc1At8D0V7b6m3xD+3+9Am
W9Ejm+wgsQwHfs7EoEK1apJ8uXLpNeql2t1iZNKhsFW2gozxH0HKGmN+WvE0VKhY8rT/0IPIRb2+
nl7LpKTR7Nw8WelRs5eKppM3F5Kzmhgn1ezHa5CqwhMIn2qT+63lDP/btWZIuVyrhdQGUgq7BhGd
0gAj1oJWSHP6Pdqaw0gNVaRAC/3q/hDQ9AYGrdi9h4aMV9S62nMOfIub9t+BZcgS/oJnCENYs3zc
tSBvmJQs201k4mhBXWRqsBWaMa7f0Lx9Q9YKrARkZ+P5QlxqvCMpg5BhI8DOatIj0S2zkyKP2Zrh
0sceLyELkLm5x1LNous1eRN1/GKmJhrS/I964f4mE4ypSaHh10PGrpDPI6qSHq8vPJYbwmhCBdTv
mrxjAjch99LKVv1mmvcgtD93Q6b9sguU6hEL14RHkx/Mf4t0ZTgxwl1npSnbT69igAPWNe8eYn40
joDGEKcvEKs3BSKr18yFCUBuRVVzg2az5tTf/HpyFUK4InTMkxm7OfQo9iZrfRUVfcx4TZ2t9q+K
wB2kVWpkDTScqMQCe6Tk/kympIQYqvumsqNtkC/wcf3Alro+XqcWLx51Oz3oSY+YQKilZ/SnwPJp
aokyJ0yRdSLy28GwZkVG3XZT94NMK/BChSI5U0ixkeGmQ2mgPNKKHlGliXl5Nthy8KfLdnq95t0n
oct02W+Vih3UN5oT9jYg0Z2I5V2tmphzW2sqg2p6jhy63DNpgjLEBcf8oiDlj/P5BTVigq4jZqC3
qdoTd/ECDx0FAubFOdp+t1qPeQvG8w28R0jrAjXApmHsr33M5igHGkLW3zSjv1QLgTj6a0Hs+J6D
ch87TVVbhgQo6mCKDVwC2xDIeSVuERoKwEW3e+Zrj3u9XwTdbwMIJdfMNmRPcoM0L58DQnFlaoUf
M1lV9lGD1eD3ebfQ3k4ShCxionVMjq7QIZ0u6ptoUk4J6xiY2JH5K0QEXbUr8S9xZAg7Fywc5AHI
F0lJ4vgZ7oLjdIlNqWdP3rYLwDxEIiJDQiPMuB6NIG/XF8c4xgydB9G7meDYpSZVrXips0X8WP5i
R3fcBo3hSckg2hfAdk5m5dU+JuSn+qNIp5EjYq3WjuoTRxidrC3azRAOPwPvlwDY2MQ4SQroqOCx
pGlg99lRPepxOo7IWTdkvRGsnXriSktkR39ymFjB7nwrdKFdWQqLOGHZEnVlYqk9FBcX+q/6OInT
wjqbe6m+Iov0lwo2CjbI0G4qEf495Dzw6cbvs20ABmXEuzglMj4QtnTskSGLVxMEgmTlBCEcYKDy
8kKJSj0PLW8wby2DD2yVbMfYnsw/YNliqXsJRNhxxuAB8Od2a3idQWhN4DRkmaarRSVOoYnzGApH
nC/lT2j/CzObMmJufCdS8JHvrQQl+j+vEXZkrWGbVcyji6kFVSvHLU2THBjwIIiTq4R/r7hhkAfp
0qOtncJqwexWRFUM9Lcsj1w57O5a982IQwqmn8BfAu8dUPA8z4LXD0qZQW57UZwaNPOuE7ZvnwOH
tW7f7dMX93jDwGqdCRo1BpLBdmSbD3UepOZHfgsZ/kF/2gKm5RKxcUMLMxUH4jl29e1d7ILSdQzP
juFJl7rLao23mFlUfzi4Mwmk7xA4yUSLAdpBl9j2mfA5LE8mrScR5pt80l9ThQk33qSulmJcOdIT
sl+YntVczpOsHtSn6jfxStxuJMxHMRw9ru/MudL8byjkwTgU8r6zyI1fTgZgbtvEaIK6aKkiU5+s
ZeIpCKrah5vwGbnxHdPWuVtfBzJlMm4LAbMec5CzdmD2RXsKeLUWk/DxdLn/dZ9vQUSdg4x/zQRf
pKreM9GNlAeVdIusbhKvUDK2DMD+oF34smiU+K5xXKukkrUzmWjKBR9d62hUs30nyuAitvMO5N3I
ARHJ9+iejl6gJGa3H8t4Dfc+D3/AYHSbz1hIc9eso0vn5fUEhKH+5rwVXOgawrwjeJ0QqbBXphv+
/H/yJyMYE6fzG46nJvCAiHcPkjawjCXa8GwCZob+Ptziq6XZBnknpq6r0+rp3/9WXFeQ3LRa4Bjg
RIXOXOfiP10WnTOd+E0ZVVraP3fyK5tNl/L98lyyOhrnLiUvzWPLg9iOY+h6tn/C/V3EaAQ/ekdu
o5+J6thI75A5j/M4eSNjkiBIDagwZiltrLylN1ytAmHhB9m4Esh2eQGtHNrjYrgtd7RZcc0bvAZh
kBohiOcKeP/+wVWkR1yVNChL42czOaCtHkmZxFc6OfUF4SEp/wcraPXzpgDEOguNOUOR2vYxPlsz
NBKfRedTo4hGzXW1yg7Cs6lQoW+3dUn9T4Xa7wAE+C1229CalrwP643tHPzQym04oLqgeNjZgu91
aqzNvUuClwOvw7taS+erlvkMCFh2R9pahpq8pF0++pngj/3dZThs5SKBthbtiB2dJByF77nF4Ffo
3iX6rvRaejRwJAfuA0y5EWyxO4AZpWuJL2LAugqkH8nUDhDpAyLlo475hGv2cQWL69WjDo1egvDq
Kn1txuG7Rl18sarcdIIuChhuObAOVfOhtq3swaOcLOB/XVpamjijZl1LnfuKEekUvqS4yGLx7grC
x6x69plY+lNSAbGU+HINQdv5VrckbXbCOuMaDE00SLqM/cQfYb1vVZdrqfvcDAf05ZK9/5EN3Od2
CZ1X5qme2fOXNZXjTFAF70vX6j5NZtYJaWB2eBepIIZfNWaQKIFL3Y4dDHwGrp+hOE5SrPFSeX8R
xeYPqnA1k/vq+cgw+OMg0tMAP/gh4yVfKE5Eg7HpbXfncSb1NwtwMHhr4GweL+gsLwkH5olJzqrC
Ttraix7vonDIh76tvJuhNkM33XvWamRE66epzWOajsPeojWywvxW1DBk6HLaQV5oV5SS/h/iMooh
hhOpGt3zZ+BNnhYsFFwzoBDHJmGHbTyXj2aGpebRtaatlSsjA9FOu+Tbciq3YHxGt4g/sZSBa1wN
STF7fGgt54MsaBwjfNoLK+hImUpnpuYnVi/kplyxtEOQy7H36zkUssowLkntmVDALrNxy5UWygYk
qGNRsPiVlZUEAHFtD7l6mGwpNNzlu6uRLOr4L+dB0FFwuphh2W3f2ts9cYyDEflwkiT4M8KYqKDm
YCxHmeEerZoFKCOfn1hMwY2r3105czcpL+eVvDLDmtiNhfBzQ/jr+YcPO0hn07/sBpacy+sSlkPS
miyLZhfqEt6uhp23q+0Pne5UOk9JD7auNO9y6Z5wC075bt06VBztWdOEyFUkoU01J5WsJQWa7E54
emyks3W7CKqzr+cfqx2mMSKR0JB85yjFhRb2nzodZyODSNzifkvifE6Ckyr0FD26i/mPuYBfnXt0
CBOGXZTD9RH+sEjTnApWATP/qHTOf6e/XcS4cGEmWulgvvXlc3IaFinSEtmHjUh3jeBN2T6fhNHO
aDaJ88woAu7hj3KkEnfC7eliUIf2z9HeN7+E7TBRsOmVARMbU4zmSyjrX0NracnBYNBqyAFfEYTn
ItBC//K6KX8/nYJFzCurwYia02RHvHGN1nQHNr/EexNroVlRP8ign/RZdlVNJC8HZQaiNWCpZuZi
adXLoYgmuha5CReV7JxJtXureT2EeHOSW6viIw1HiKB+WL+/Eu2129Jk9bZJhIApLY1XQOuSVqVd
WcbAF9MLPbkC7LL2wtaN8aDc4N2WD3pex01El43xJBas6ucv3p2YVsgdBBqpNHBRPZ1/V5zzFgMC
86O9tNjZf+FUEOd2OCBTxbN+3/s+xUtNBB06xiMem0csBteQlU5Glpk64Zi9gr1oVwHl5JpS2+A6
s0oxhXlsl2fgg05cDzsfMQX8n3aq7QD/tqskeWQ0Gl2pQ8Ep5CMMJZsVgQBSDE5aZWfsPCe3GI/D
ux1ZnVxkNOtR1e5bWW2m+7oc4R38zbqVDZKtlD+40nbj2zQKB8OILaGmHDuudatSth6hm6fJabou
uEjwQp8HgAZl81grmY7928zTXRa3zBFQHRV13QDLgUlv65WbeiV/fwr108+gYk23fjYuUcBdjSkt
guv4eZqj+SjoSHeT6mcrXDSOvJZ8XeC6u1+TFDqu488gzOGrbOm1gNROkysvwYuyNel8mvKtaX3u
bc8KDTap+DU0T3pgHQeG7v1bAac1IlHbU5uZw3r4yNlxZEmdIagy0qIT1md9ualIK9ozAZGXsSek
EoQYCahnlqqaQM9+ljU+OVeBLRUrmjNgAA9pWrHGGhD2oGXu+TzLUSrKqS6RalfYMWqaj9MAddxl
K6DWFMmdsPqy0d/fsX1WGtWQSVFHUzyz18AQcUpBr8rjNETtDDLT5yWe9kGU3aV7kT0Tdxo5NiCO
Cs7jXrzCoKyN3AZ4rc47f0qJiSIRjSNOqU7iZVxXS03y45EtYO2n4H7+UsM8owielMLSyupTUiS+
cPbG4PVfBUIu67UObMYs+uOgBcp8abZArcdIYZqNz0A5IPzXQd6DUoNaeFUklxBbHziMNkVjAQX3
/jFWUPJzErMI5jcYYxdJWJ3UdTbgHlm+3Y4SvJOFaXTJc64sx8Di58MmVybm6SSoAiTEUUmEra3Z
/jFge9D+HE1WJ2stdjUIjXCMOAoYXJ6IebbNf2ngl+ID57BTT0oV7ALX2L5BytSfdQWrZH9ZdW78
VgnciuNGh19nX0ArcfjyWWvge9X0OkjhBEly2fLt4K8wfS9voN0ZD1XcH9jVhaaCtqkVWAy8YDer
hvaByX1Y28TaqYc0aMipNcfIfMqxelSWVvgyp54q2JXpWQenV2gLnBZW834X6GkgNUxJJQZwCinv
iM8nja6McM4dU3foQdzHeB4M9GFgrUtPzsP7LlTaMMvZr2TtmWoflMhsA2nVNlCNYML8vsHwRUot
JbQW/fw2eWnfQBjSFZfm/aByrLlHANbHEHSaMJ48GuvvX/s1J0B9W8zlx5VueSbdXC9RqlL5wWJB
XVGBnahSZgUzCnLkxVuQgeKN98rP60tU1RP4omTFgmFqvWEZnlPVjbIyiwpRS+WfSpYbbPyo7tDU
I/lMWmTPYHJGiUE3NgMPyEnBes1rEkim+hrNfeas1qFQ3XhvffQSEqrcDnPWgWvTTFQFN1o/gaF9
NPZPFiB/UFVnKQVjRcIqx/Af/5iDVbJY0/JSsDb7XyujrAaW3EbP1ml8nNWeSK/uTFQ58D9gwFV+
ejZFPNjXxkUmAlIoaHlHo8wGlEvIQZsXEf2XjCTH2eWgDNwIdN85QiGq8lbgsOi96VkJSFJ36Rg8
FbBN5fN6oahcTWT2XrLLgPZtSwyErqzJbp3V4B/gJCwgCWPpHpZivBKIh/JbsvJVwWuIJN369ckB
105Af50BsFFBoDvBqFc/QlXvDy+0sUez8Dgtoaz5mTpFUnKnTJDKE4R5P2Md2xFCP9GtDWHiwaJA
RUJgW+QYgvKbDIdHkQvDl1hdeKwWk+HGfZD3NruHjP0A2f71HTzru6lXCMuxtsbZs6w/Xl2xL9uM
Uz7BzAL9hcXjA7qvavA/UUJFRqe+ZmoieIgQBSTmN4m4kulBlMZ9UyBN3wlASgD4sJFfu1iG9RqT
ruNquICWcd7Tf9xF71EiOeKboI3nMs3RxJxYXjyANg98Cr80ulL57x5bZMZpAR7BLWOuYb6Q+HPB
EiYOCNc3leBrebSf/SDTXXZZMMy/fsYL2IYfh5YJzEERtn8vJ5rIhKfsRwOEhFpvBe2j2hP2ddWU
RWILjaIjvzmw/hTcse2qHk+O2QHCT7s/z8G5oDeHirKc5pzdtSxX1TzdzhMuhe6opEGfk+dNWygi
PlqHjH5cK85K1kVWMkAlrm1V/gU7T2I9UJyPEkIsrBuycDSQwgIWs7YUd5w1O8JNL5Q+VlSHOzR9
veLOS+QSJ+WlVLARcy9yuZyhojhkHR15pwhjLla/XrE4pNsrouAroa5XRGcTk1GIsYSE4dmlwdHw
lylENUyKG7VzmPY391icXpRvam0H9aH4joZiHGy+Q6WgtgBRQkbMU4P1CAzBuQRFZ91rZSW2uCm1
P2FnTD5HjKwEgJPCDac9L2YgUF+FLiL7BcnDuSl1e5tSRq5UWt2mI8JuXMC5wx4Eo7JkrH7mug0k
coabxmo2W6tIT0NVgU87ZSx0cjo7ZHfBibkCukVvHaleRHyLr/1/Z8LCtM3Fv+tbXXeBYnWHBWCd
xxqbpx/TVJeE2uYy+UPwwtR9GTjjPYXxuY507ytiheTrXQZmAefINSK7JZAiCErz2CtYtQVlfVdq
c1Lm824Dj7Hm7bqJEJTkCrKHp2xw/Q4+doySK4pDynJXMA6EwuARzhceX0IkItc0EJbTO8ayS5Pn
YDYeGyn0DKQEq5p8/RpqzPOn3QgGeUJvdUQ5JtKUTxL0nEnPRbPvxwsekP6oeQUh8JtORJ1xTlnI
+i9n7u2TzCS1MFrIotP/RLks4lJT7YLEvlomlF/A9s4xI7DHMPNPxHkkz/g4j1B+xn7wg936Iy7m
zJoUY3l3yj/Cino0nCe7h893GMnNfTbyhQ9HBd7NRKDf4NI45kx1YiVMKBNL4p/ev/lN5+OUqnbH
M9PuuPEzPDVPsnAi0JSwtz3fw0Jbr/DzYZftRKORySBUaDSXA2fjN7CyIFDZjiHJyECWH7e15dvC
VXAvY6TMJmT64a1Dw0EwLcWYtKE39ghT32vzxrj0DHT61Ib4qxmHJbUUZnMlxpcGVMxbD4VZImGZ
h4x7q4Mf9I7r1cYBAXbnYsNIacwkGC+1WxmWtTjznN7fYlIkNvFBLgvynW3RM3/5zFgnjhQDRBkB
RCx60HqEFC1HsRwqM+6xdjzXdnrO3xFPhJ4oYOSk4S9i5Rs8JSWBvzqyOT/RR088MfPzxyswgUBT
pWx/wGe63sCUbwOUFGjyKiKHs+to03FRkkCC5h6Id1VJ/mvN5BhcxzhyjtaXgjFwi5rIJ8BdRF2z
34qA1ip/xYRkfjork/nWPxfcDpsb6cpU8+EJ0TWFvjE0eT7LExBn3HOALStqSBfi4zO3NjgnlF3i
+IRMrl9YJrx16I7D2mBpnby/uEpZSTmrn7RDk1RHiuyEuMUFVyUNwlnxIxodGcXT33Tn0rspKmr4
viPt8FgjjUcipWfwJelsNhhsY5w0CGsLOVxR77z6Sweg0WvjkmseLLM13aknKk1JPlQMvnSG1ZCx
yLxDddFZhjCZtkcWmFEYn1ULh1comNa+JRgqNlpcGouGWZgU3sbRKLY+K08voVEtK2w+uptiHNNY
yEONK0YDBM2Ziw+MqEWV7ZJl6sOQaQodILJNL+Z05fwN/DKi/ziQWdpZlRaQb5SlsD8LG5zMKfpo
R/4wXbm7WdWjJq+IsAoNuj676sxa5pIargwVlZrYsNQzdohtmfD8ZH3gHlEXANjClEMEbV+zqamH
+ToC5CJ6MU1GHDm1DrP5LIPhr6PB7qvGJdiCqR9q4+BNZd6wabtGyI1D1pKAB13nGYSip41NNpXl
zvYUVm1Z7iU8z8DYSUQudK7tZTqsF5bwKw9/mwH7qQiyKfvO+CqXRWLsPd+0w09ten7p6I78e67v
Ga4cfJ/ZmmCJ0MhCVtO3FhYIBu5GYOI4FSW1EJHIUB/voz95at0FODbO8Op2GM5646ITKyLoJ+hT
pnbx9zhARZzzj++8hOWT4lW2jtqRLORnQjFnVP2ezUw0S4DB0YDAGhvf8JhYSJULTbGqa9UV3Xin
NVSmQfXsH9DqGz19zz3ZbAGYoE09OsGAlaNlCN4DISCXu1JInhYsaNCSFJPqUq7Q+fnmSuHCFiyN
5DVS2ekd5jng8eoE2rO2xybg8k447ItWPzJOGUD81bEYvHlTJ+0A7XdNAt+y36+FDh4crzchqTRD
73wNAC2YmYVyw8q+CTMdTDVL2FvtAGyKvfFs0jO2QG5EWJpTax0NGwFbTzv+l87F1CI5YgRfP6ZE
dqtgc972Gb2Qhqo4rku9wohWyBu4XaErnfrVfwqQ54qVhw4BEcJcJsqYUGzHHkaoL21scXknFPrv
V84+X5Ee3kcQXBOjB/StDdc69bnAg27tALFzhcQNDKX5vYmROp6HU8s9xi0pH55rQsQL2RjXfxW+
Fe7nI4X3xHJCthBUfJopaDQbvvs16zPqmcua7M7yQWbtH0ILqF4IktUPjCf8AHgj9Ae15FmFM4nf
My+pCoB4ywywwFS5PIXMdnlSKYovmyTsH6bQjoOdHqTqp6Iv0tJeDHvoV/W5aClM6xwF0GABLk5R
4ChKY9wigXkKK1vdaU/IMGXOPurJjvCcwnbwgJOPC9MT10JDvxPUBX2ndu1LFUJqPQKr19zbiVqq
DoQIw3vrdXTZ8hsghSSyouIXxgQjDLCF3o026Iy8+f7tVK7uHDzxoPb/u6H8oppZtT/XWruOB9Vx
mEu2X7e1WYqThWpnqzSSUQNk8zXYc5xNtNGkvl9ExGuEo3Tm/dMpjKhZ5ZlJgjg7u1lqFbOLV1OG
KcxoKGuqtS031ZLsIlch4/wMlNUa6Fm0TRjIDuCEhfuwLpXvkpb0NUvvBGbEVaiWqSJ12/jUZpWE
xjRfBSJDrAQAJlzzpPdCs0f/sl7tla2OYsUw1aj96Qp4SGwoPE1vHpEr1VjK4wor3A/YUGnJTgeF
fVbH8685suVoQiPBxWN6Y/GfE8/3prfu908VXRGpWICEM4tL+gl6oA60BsYQcb2JHKBnKhEC3wpJ
2FuMsXql6XxoVy/O1xFvsuV8/N4q3m9RE+Ud43Mm7gvutbnKPSpInvKUXrQQu6hs5nPWJKlHrZ0y
PZLaQYeIZWuUJoPmWn8kMe2mvF4hi6mKK7CkUliytDrrRFPqPL7MEUNGuAJpzH22reFG8VfqEGFT
q94R/EovO/9FTNvkLyR8KmV5lmVMxF7Tr3S21uNRYx4lXqylqVxiFeebk5Mlj59kTw2U5vRaZlzc
wJpaM6eIAaK8c9SlFB/Yst5y4Jawdu1KyD8fp1xosRw2NkKCt/phHWYLjt+B56yjU9eirDPC4Gkn
TDVkOJ84g/dmAjdMu+QsDTEGFCtn85zv+thzMOeBCbS89uh9WBaKci/+oFbK3AAeyOkXeJX5/Lue
Vrj5SV5A+KApkNT6c8ZgaukEWHp5EvQM2RhJ6143rkx22uNAE84srurn8gA85U1tjpRRp3dQv1D9
ccYCtJlKbHoddAEZFPeUPHD4rVvVFKWEhTjm2tAw+ic28/be0NVcMNlunPijsN8C6mKruG+p4b0M
8xwXs4F3RzMyBwiG0oC+T3LOs2b35bJJKFbzENtwxBDLe01DCyW41Kw3hnMlRXCS2Qisg6gTLc8Y
LUm5qXb6j4dtD2AAO0RtCfguQCjpT4Z+fKk6m+UUAvm5Wa/pDfyktGffbL6Je9XAKl1aFdK8Cz4c
Wa2ioyG2mU9s9W3C+tYo9Zfasm74ZRRHaHtAoVgExO4ktH78NJnmNl4kBE2gLDW4dPNGCDqadQfo
B9Ub0WPIZhRHCg/7q06uZf0XemBIT02/LhtQNCqhBS9/AW86ErdDKKJOhhb6/CF5zTJgb2IXBjbW
QPnbJCBcCWUzH7/kDokpgju6EgBhltBt4KrDHmOJzTZkNvgsuzbdk6JuwyR74HVWiy5Rumhnv7q8
/2AWJivCv3EZbFYcJ3ngEV6mDgaaNdZ4zW1SE8+4sGuDSdpVwgOY5cNT2vCoorFj09WaC6mZHBbA
NEq9c7PZvJFgaH6eVhTqVFGIKJqj8DbnzaOky+N3J3BhKk1Dw2DrLvIVL7dzId1r8YHAVBHkPNeX
r0sPT20djF851Z/OYT95EAZq4IBmlkE05bIoHPK0BynsUPAEknD0wmIylrKF8ybB1gI1CvWjuptc
cOT4+t9ea0OSnN1QtNl5Os0aAyi9EPVck6z5bFTNCnlaC/eHJIn3Q8lSPOC6Wpa1yXA1PkUi8mgZ
mICGGu7rmY3n4zw5MiEKkMpQCcQMAVCDLlPBxZ3q17x1PY8t0SoAMmhWHm3SCLs3cY8ES7vZNrFS
5i3j/3PjS52js533YMWLLG2EYHSEb4a92Pz5Mme3gfpjRp+twOPd45UX1O8E89z0nOBD1huaG4Ud
wdaGvWkZNwzWqh+1EwB0VmTCB1yF928a2MiPRphZeJXJUr9vQU8RzEjSXlUz/QDdRhQH4t7FVehA
9UjlflBg0YUMkNmSYeQgFcpJn9BOVdWfqSfADEXwP8ZgrTiuUD4aYUDu/mTncEary1wrjCMg6fS8
eIT3RSJG15GoXj/D1DkwFsyoZstB2i0CsQSaqphpYEndbn9P4o5AcHTabTz/Euy9jPwxSkfRNEnP
DaspJHcehx5r7piwmNmETVne1P3NgWakdGpn77Rk9hZLznKv7Evza18NnRQ+avumpAbSNc0ksqXN
kb/1EqSltHVT5vbkQ14O0dbLk3rBXkFU/oFpORp+DfoA+eB5i7LScV+6qu8p6lRuVTxbi030F4KR
0dNz8lMjtztbQzEHQs6PueUZFS0rLZYd1kVRJdrnJqistLgIr36AKklS0p9/DljfIeDVyG/Yhb51
SkUgVc8/V0mZLQ14lqFOOhUqCL/jxRX2v+TWULi9UKzmfF7UOgUeUwNsc2TupuSQqSVNp8nTR93c
4qbqZ9pTkibCw/GaCb++srgxE7t8y1QkpKYPiyu5jEcRkNNq3QXl49WVZq8hcDsZBFXs3ELaIbvW
VgxdZM0ThmTzdLmoqsYGqgbhYNSRMoJhpP0YHqF+77PLDyryW3qhyTYAKQnZFCaAJlfKCW1W8FZy
mkXb8eqqeWLewbcxu7cTqCU5hHXfYm9SlIaElx0NZqtbrDa44BdLAOeqVF2/07c0FiSL7rEOPUpp
5iKDMXnW7+/UVOk01O+29rqS5LEnOrp1Jdr4Jo/Lvj/0qFFJakhy/T0ukgoV1/a9pAwJWnVn+oXw
7H2gp79dV/ycxzd1Nh98WV9vrCOfWc14K0TWCIfVBfD2UIxL8TZjnBgm71HN1jRfP9nFNf89Ittj
nSZtofFWBPlgjLHZN7kD/c8V5yqCmrYpGnvZhr5YMSDvxrIaEhRbWmJI4DrDcGn07ZaWUbpo0Cm/
+p1MpohPnjCpWMzkN1U5X3EsVS6Ocv+RBOuY6O65OTZpWbr2omnqWfdRnrghFXFgWV4m9a17Dt5o
4z0GDMf0zI05tYfq9EEcYEuk7GX6oF4HO1SWHwWFOlyfQEglmjsbg2tvy+mde88rUBBmuOrQlLGF
ShM33WKAFyXzbR/XR5Dznzi5HQlx3ndY4YCwTtBvBsALcUZwaR7/OjN7dQId54cm9odDt5BhGHpJ
AESHS4j1M/ZJ7XYWPqX5bsjxIWyV7EtmHt95d3lSIN2bT5Qnz1Pex2a3btgV/hgmhEMsVhs5dUJC
GQSHsoeM9s4lDzf/DH42ZDMbly+6VvYPmjYAX7ZR/7GtZlYWaXU1KvVaOzKXeqOJ3UWbCkFjk4DT
ZFLEfYCJFsbxowLBD5Sdl8AkzTGxfA81gw8JYF0glkwQrcGVhMkYVHC6v6E/p32h5lvRR/Vy41HH
qnG3EGiD7/zUKWpQqitg8totw7O9XuYvuHydZfcv37aLysmQKnA1Nwo+RLCmpU40k4fMYsHP/HVu
lB3IrGNZRUqW3gFiA3o2gV1XDK/kfaLdetNjkHae2cdMLwRe/bLWBuAApuZ0WCknhtuFnDNQGu+t
I5uVNlZVkA6G919Q0YumGw8LRoXZYbxHz40rcDVDUY/D8x5Wtz3ynPj/YBRaVZkEqWnQeHMjNMlS
+ymHAEaOk/qLCW8I9XVC7OQEe1EGi//vas0IZwd3D1sNzdRoRxcW9YNCoN7LQBOBEzDAseuEbkw0
czukNW+PyP1x+8qF+NAAny4J3dmO3KPH3/giVOuJyRpjkR8k+A1XxP1tWM9URaub99b6cr2MOhad
/jD2aNZx9RoC0iBlILuKNCRlegja9uyLzEMK2icN0ObjBvuky41ZzMKUeTKfQfsolcNrnbdC2rLT
zNBtJJ2uqfmLjYts2GgpLAv6THChTO2xRVXMIVvCrqwszIIwW9sooL0TydlagQlOav8Oe8rko0G0
qcycPsv+2n7HuldiWPSuRrEmfzUpQabLHM/DIIr2RcUAva92Z/J9yxf5kD3M4VS+mPcVENIjXthL
G2JjVVY+EHN1mAj9t4lxZQC6rd8Qp+CTQHWvn41aqVnZpmc9t2Faz55Wezf9nblhBrFJ2kNxFEo+
Z+KCduUTEM+KvcXxjx723KFOsE+LqJAZx2cyRpCvNIvwjhhgi5PujlT7i7SUpL4jgQCyRTL0RA0z
hx3MNde0DEYgN99jeEWvKLOGJbzj3Bwj/gP2mkhi2aEYS4lv7NM94anfnyYvIWWE+jXfIfKJqjG+
6zTZ0JFkrys3pDAhU9z8q6Gu5cWyDVHGqceINWJ+zepGanFmT0Cncbg92LTsY36mXEkUVZfoYaWU
CrhvCfD7OQLPB8WKMRHu7MRLOU58DuU97zy0kDguE09Sdd065oE6jhhQIlRy7EFNHJshPTTZx1Ji
qWLsYdzPmRKnDH9xCQM/9R3PIuYUsf1bun/Afg30KGeo2vtFKnKMAW8oU7F/CHzoGXlPP1M2NV+j
xgT3HeGKy7fX14t0wKFgLTJt32c1QAMjDW6AY58oeDYrk59cIJPDoFa2vOP50iX/ZUcDp5U8lFvL
6bKe0X0wt7p4+Kzj4KYB4u7TQJYysxH0KqGF5ekde0L23nvpIUcYm8wbxXAe4YOAAfMc+mDHehXM
EwvOpbnAXQ+SnBYsbeF6EgG9uKAsMZYSpIbMarDSZV9gT4cxwkvWxDt5GH8DH3V/wTtRCib9VCva
Xy/IPR0ERu/3bsCCjLSeAOPDxIWMn4ryphFrXRjnL1PFoZUXNfNFf3WWWOpTwVxtKaxMNV/2GHFY
cRJdf7HQK5nxH0lO73kUhNlt+DyLrKSqzvkVv7sdVZTMyRfH0LiDDob0fQW4xEkRwgrxSf9o8P7b
PL1tasxM81pFBZCbmqCaAEs+2OooA8+T4dulsATZ4kqi+sw0xm1sJQhV03xvaRzk0EbHqDPP4GjY
Hc8B4EQ9v2MbFWzrgbf4i+IJ9gajLX0n9AnEp3G5ZDbWIwhIBIVKEpQVaofyOetfdGY6XoxUOCN6
obF+biVlL5YKBWb4/fDyTCbLhpMRbKyjlnxx1KWQzjWICMCyYM065zUdLTFelu606WyuAStxvrCY
vHn0FAzasOU18gnAd2k0cM6gItnEKRfCWmOhGVYbVvbQC26zhRUt0UnP9EIcQnUGqQ9zS+f+RnJj
8wkLjlAnrrqz88b1yiiKWSg9Zx4uOhlAJMTgmUksZcfiNNwqYcsMSG/C9mnJfHyZB4CxOy0Yr6yX
YOCgRmF/E83WW9A2PNQVaz7CFr/Y4ohd3m2zqEdcLzWv/v0/BYbDlpt1CTdyNeuXhyNyBZingXx4
I5j56cQLFTZlPeKn2aRiBPkU+8Rd4RD2hKJrQARILpZqQR65rJl8WObSGSc+JGf/xZqgNNDW93g7
FMqWb5aC/84MPJuVTOKeaPKfLOFhVcV8CmEb0FQ/OhX53mRbuCU+TXCSFarNUYXRNXiNxtX+XO5D
S1TH5GA6crgNJe7D4uq91cU21kUS8VFR7+SKGpjOSO+9keGma2oqniEGusA2IJ6G7uFqoSts0NZm
qJKDNkM+t9gR9GxCqdl6nSR07cF15lYPohpwGNSFs/0QgBK4iEJ0OcBpcd5aYPjvf0S4c1Mg2Gjy
pv12YKexQyyK4Du8xSDUrU41tUrUFlyJqf3vfqXEzWBRUyeYq91+FhiILqA9gYFhXRs0T7Fn4rp4
HFVe8bvuw/cAoj0LAe05nFTu0QfVIQFAZjmQmpM1wAMGDpPS4K0TcwrSMl3N8+DO2jaLIjaROCm6
Q/0IBBHMno9WgUoo5rRFnqOwG5kzzGVbbPjqnnYzZS+oiGZNZmjSXuxiaXyod/KPg/93wh0oNHT5
jWUKZ+GjrZvqyAgUZDxdLekMcLQBu0DhuSnvPnmCE+buu7LccrhwhN0fO1NyL8qqLkRXY3H6tqMj
veDR9WJN8sMEQGDugYH3zN77gtoDfJX3oVke9S8DJhn4ZR6R0475okY73bXjOKW6ekPGAz4yDNWi
r1+mTLW+ENd1MME+CXDOO6o5dx5ign+2H6FpDiWM/w0lmwodJpBNP7MoQyC7HBG9wSqEuMxkhDyE
x3iJpD+Oi/OP/SH3UQhqY0vFmQnwRUoYDU3Lxx+/bABz/Atx8ZHo6POIPRAEWh/Cs1SNfJw8F7+8
Mpn94bI9z421lLryVRsgyvcvQbVBrSkdarNci0HvZbmtsZR+7LOTiqLNezcldUVdkaj0RQX+Mcuy
VZpwdw1ZJ5Blr3ifL0y9bxbfwnk6QWQCbECrTGAksKD72EESlJbD+fX9svlhUMyV+8pU8l1OgBNo
NsB39+EE9JI5e1FI/7s/TF4bPlXXsrQjA2frAuIxev54HfD+t0/dniOGsSCucsiyQ+q+hYJUyNyB
cnLKeD9J0x1rCaJ+yNSWPxcftJgDKD3I6jmXNf1THSuEx0FRVTMD3nvdwIrZy8kejUVPYifKxTcZ
f0Hv2wJnnbGcx1ipyL2YN0TOb466cou0ahpJgm5qFY7tnyDjG5PF/BxZDYWW75dL17u4ARXJHOse
mCHKA/Y8BySnboJ/NeyOz1UZaynFsy3CfFC7xoZ1H0FnDi+TJqmTBqkxOyEPc6DiOV6oH9GttxQl
KaTQOrN5k/KRpAg8Gr7jXYfwvvM+HYuTh6CEEIUq0vyzATIqG6mfJPtg0H5ZnK4FWq6sjzv9m0AT
yfNA3vJXxay5sFDqAi/xg5C0OhyMhl1QY92nu5UOLIULscuaWsqiq1GIC7xRW4EkfdZ5n14LDjB+
Is6rH838WO6BCQqzhG4KwMujDnooYHYXxGl2DrMeafzSFgojS+xbjQNM2f6OqI3M8/iXX86gl+g1
cWiRjIYm8UzHpIU8HMJaaYL3w3FgqMNjaVWKB+Rv9kTWvuLt3SrEAOI5UEdTWK/nwBCBMBMvZ/9i
qAz/VTuCZ9JvqDidJGt+R4a64piZaiWoGvAEqQSFidE5iNLYrhXHEHdKETZVhiq1c7hcI1NwD8gM
dd+2C5rwI73rhOw6e55Um9EQJGAB9jdGexX6XVfIKbcQXh1d+595gSxkRNY6ggp7AKI39VtEnhZh
MbgKGSXKZxnNev5HMcoodV2YCcyin9xoxk5NvAqOvvNxu7Tb8an2jsRKW0YjeCL+7rKOqtdMGSaK
it/5P0ol0aktc3+OhFXfaqux4uCQ7z26iB1z9YUE+0n2D0H3ZgDSyLeNFSOGt+kvzrF1QTjdovxu
bq7bXCTI3HnWBTKrN5z4o6ggdeJTSu5hJW77qsaZ/H+D0NPOXw4dQMrHMWHb42xsD6TiKU8vmhhp
pIpfhX0r4kRanCTmB1FiXmfHO7jIj5kQEcCpUoSalEf19r74zykyoolUawBV/yQpCw6rzfKMDscZ
VCOz6fqFFMicX4cl7ng7TUoQZ7IEIfRw8RXolrJS1nJt+csX6T0s8WwAPZUJc5AQDsh1EEtAmmjk
yPbleEmcsz7IVGAG1zAYmhKwRpkOVj07fsIHebWzginb1BFT1z/sgyosaAQagEgGiHMynfDb0WYx
vFQWu4yvMez2Mcu4c62JxViQV4EqYcAokyl0ueuTLl881nJPF67Jym8YwdAZZiDtOpc5ugr++PKk
LAiL1T1TaV+PtcoAc7nUasqpCyG2vZ8GyWF8JRYEw6vFiLDKHT8GxbbwRyIruq3DEhRWjyoLrm28
bHto7wLRh6FxNAvpFPD6nVl8ZM+kIP07duiyRtg2ft8Kv1QwIX5gMzNVhKIqhxJ1dM4568N9bVV6
XT/V8/7i+ekt1nXCpxoKsG4lTIofyRwTc/+66NXvbpRR7+weH2i0uYmNI1Q7LwP2HgpE1+fHCt9w
KU9JOw+NNo73dD2MMwNVgKVZTJBqCghEn6ZtHZOZ8Di7FB8n3pxClEu/uxFUAIhAbNMhnHsboHcc
ZBnxuabEb3wkZ6P38zAEyzXT0MGPEFO6bWmFjJoZbF5kb9EL8vGqk19lXVRKU65tb1DFV4LJ7FLF
nfhKMMhAbOgeT3vuQrB1rTMLcZiQ8/u0naua8xR0dt3jQinmnwf8CRRoqoaVPDvw6P/jlMFlwF35
Ghs4BhU2mAhkRfDzltL1+qeRLmZFZB4RPRdunbMWdLmj+QQF1YwfsenOnRv7FLFB78Bf8qR4UMNE
QGcCjqaxpqN6hs3m3dt89WONuxOHFvfdIaOuVY2DiglDLbJSYPuqv/NVeAP6UfC3flCclUTj3wxo
3gWjvkHThJmbvFOsoeVRHDv8ac+GoMmCDkvbEyG1sTfp7FFDXukRXL/Omfu2ZCh4gCxE0W3JeEjo
hkTbzsIRInR7vfdqSAT7gi60O0n2B6hrJ98NumSPvCYIKmYBt8iyjltRDfScGDQj77SfLPHaYGC0
S8X+kzlWxmzbKe6EUNafCEmxcPQAqP/xFXj90nPPxntFDF2h4Ql1Is86NDC6d5Aycku601Yrp7Rw
GQ6dkYoOjnXTcULQXmpnaWhR59PJyx02rIuaO/9Q0OeQOp+hiVxorBIwih7ijumiZ5/TcbW41FkG
8ywgq47XoTdw0zzek3+gZ31FG/ssT8ZzqLDn3Qm/HWqS/fhK7Sa8D/2hWmYbg+GPzpLwwMoZyzc/
WXI+Arf90DSJKGmdGbY3bvBnqK27atTF+OcPtS+B5gmUUB/xZK35sdmYTJxLGDo2Fwmmf9bIYLmH
34q8Svio5V8Hq/6ohdJ7phOh2rBPoWhOg5fvvdvCz+yGnLXqpVL379ZbpgE9TlUZpq3+lAPcDywQ
FOkytwMMx8M5BV9CB/KcUIqUCdqW4Gn6YThDTpnQiMYg7npbhzaFER7cu1y6mXCFXEEFdDZIrjOq
+iRYVAh6BSiQdLP++ixqSkKnBjKmlvvDqjz7EFlcnvETTsroYdfYbyQboYZoe5R7zDLNN39Jtfl8
3Oij/GuGQfTjLlcmjj5s5eKLVEbrXVL0DVhy9sUOLmpCnLCn3qq/QsB2SNMyxsdWZe8HFTr2CYA2
VwAh8dtpXujcegVs81okRoi5ayDemQpTresFGdIcdREVV1bhSUNb1VJT/U1ptI97yYr8IQnAaGPB
IBQZt+qJlNxP1i1NQPN93bXXqqV9aDj5/5Zdztpkb9chsHnkhsPl7mMwIc95RA4SRaE+JsgoqEOj
hENKU0Dckc2k1N293TMOaUxUFrNsvM47GzI75PEMnpsn1EHCMElQ091aB3B/jCVth+js7edpnHvb
cmKAZ/qH8KB8g11dT3pd1YasBoe1dNThPAHWAS5sKUaXBurNikMOH5XzB+mjjN0HTDirRaxJ+FQG
mPQmdfQOYeYVgI77xZjopjjCAa9ULPjtayO+eTWMtq2GniOmjCQZ7hYkgIIWGf+6Xfb8RHFgm4wf
jrpfm0qj+C7+GvNpkdzL4Ys2UkAj3fFPfCVQBEa/jCUEHttK4O0ZNBF/jt+GtXDZZJKgLSRTkD2H
NtwQooxevjmvwZwAOxRKY6+wiVcJ+aaRXiYvGrolDxZEbpIOZAts0bO0DY15G272C5BEIe5SNdNF
lEn3kCqolvcFywEXdp4+bR7gRsplPMnVUpdS+YSYEBK4FrHkcI42SHWa5BO69jS8wZYieJ0/hXRN
Vf4PzNWH9q/KYVYX9xBXj/L6j6MHmnYXUXr4HUvMVAkXC3suF4DfqIHAXvNYamdf4Aym0VqZikVp
sUH3MAJZZBFJaM8db4ToFWOFjbh69qM5o8lV7S8/1vqpuHCq9UqOVSmgz9bHyLEACXb7U4+RKJOj
rba8RB88NbFktPPROyPdXLz/+s1Vyu8ETdhQMTKl80DneyCuSfzbO1s+k92x8Obm8kHKgczWOPHY
6wFZCwCpEgx8O0p5I76ccQ9I5rNVLdmqkM3ysu9fS7zGShqItF0CTXe67rV8ZdcMf9kuJYcs8Sug
ZuQr4Mtt9nKzcgc2LTAiPiOmtot7iFAWq8LcinoyNJiqhCsHCcUe1YAGMnr57KLhX9XOnJhbIiHK
bTrxQ1XoGjbhtZHad0PC6rgN7U1rAytu9TZjC2OtelQNIgww4x2dZJpu6Y5XXH7/ZGew1hMlZdjI
4zxNzADAIf7c33DmXiNjU1cNQoh/wXOy8lTNdwMq8DrrCsEG2gGcept1AttAuC+MLwn3H/J04pA0
+lQe1IXboeHpHTiHXI1vokiPgCoONGFAcdUumE4LSzv9ka4L6FSEBqQVruMKBx/u2rGpZ5CoXKk5
IE/ERQ57kz9doC1HC/ZL3MnnmlvxeJAiA9cmBcXlYUx3kF6diJ1linABgveJN3YM5CRVG3/eFclj
G3o2eCcL/z80PH7XpymiV/JgtlMpsBZxKjwyqoh29ccW61o7N7bKPx2kiD9Nm88pLmmZ6N8y/ghF
gjRq44qlO0yMmJ+9JZcuH6k+LiOOTeE9Guml4T9Zp2ydmXofzP0HnLr8f3Wj+CB42ljEyV7YMrHz
4YuYBZpjOmsUJlk1xx1GjJhyNMqFobwJn2urdGAm3eCpup68V4SeFUKpIZzvS64uXptyyiTaKu87
OhJ1oTXXzu39l5k1lFkBtHCzmIDfirle0yAj3dRrjIKDZfnXil0TukUt2n0mC2ymX1pZBuDN7fYD
ct9rSCXIprj1J4JkkKR6LsBdk+MjC03Q83v9NVob2e0q9VWJXvvwRUMeKYt+1k0bApQHEe0l9BIN
+hOvlpr7Yo9zmtuC0RPGKBIqUXBVq6RPQnpOF/3gGj6ChRq2XG85YH73qoIkWxuOMiJpKMmuKucL
trVE7762CaoKHMclYZZE4/hT/D6wZq3qTOywsS8a7sNE6Fi/IOkNhkcW5YbfR1yUXLc1de49xAO+
IfK+o4SGxoxtWjdITzJqHQHMolyeyoGM2/aXINq4S55VbZVPJdQhftCwrTWke7ZnoeL2YXQXRl+m
i7T+3d90InYc9MMiUCbDXkTZaGLU+MF1qZ1H7MUdsZUMLUeZH2D+9aEY3W0AWXhGAamXtwamovoO
eDMPmvrBYjh2rpkQ754ouM5bjjt8UdtzkmMAHLOO1DZKW2f1QwWxx5JrT/prdj+8+rePI4o9y5X9
YrB5dDy3McOJmQBYNTE6Wu8xoyowgmhJmCPZiIdIQpGKVjdskcrskwBIQYp6a+6aedXchT7v005N
09JvzIvznd2VGMFFzgrA86kV7YS/p1JelCk7HgK1NHMbIbunypB0YS34II+nCrVA8NXz23geThAu
/DV0DZjyHoA+r4jUQMzxS1emCbbaUOBGJ6ZmgnGlyxPnT0dNgXDr7Cy0wxe4Oy5GUUXvZ5ylkoS2
M40jr7frf53Bskujtnw7O6t3h+tIruSTZKbVu6n4aaWXhsZy8FcwThWWsD1aUSlhWJquai0QjfVc
JrX6G7hMMeW1g5pfEll8Egb+qH9RQRV6ZOJ0xO13gjs4lV7HvQ9dZbO7tF55re1HF3JEQ+13cmfR
WB3iKIvkAXiKyRg5Zfh5CHyCx7gNsYLXQ3vmSjtG8BxxQnqgbVvZgJq43XG7oxhxCUIC53rJgKzj
X+BYLwGoqxDz6q+c25z7quVlx+Rivp/jmtA4qNo204Y5BdrxZ5MWRR7KqdRp1ONtC4eyhTFXxQDD
2da9G5yyEAGX4F9WdQGUrAWYF63AbONSr6pjMfMeElRl/YUgU74hz7RSs4UE9/Sf/fiDTsTxeYfV
ILqOg7fsTqcr6TBAGY5WBSDnzPiBDLQlWW4y3ROcuL9Ds+2McPr8DfDvvBYNLiovt6bQ0tpEP1yz
xxyz4ZQhdxAKh76wNiesiQ7V5tEQYXm72nKRZ1wGLJLs+T9u6Ya7JKkhuLQFjo3tUXhZU2UkXWt5
ZPfCRZcWmzzJvtz7DzmQSbuUCMI9PD5YDd7cxpNjiA/4mKPEEDTjDo8K0lFOfCftlaSVS8j0KWgz
l6Xc+20RwdUCk+/FcpA5qVG7I8YzIZjpw3Ps0U06tBy8DL8VpzDPdgp3fS/1xUN+ERAphyoNyECf
fqiuRNVUogsYVOZFg2NmLxoCk98Ts7kDNpWvNsl3BvtCEQwhtjpBB8apVX5ED6wEGa8lR+hO9tpj
LRGrXtY1pwLki525EghwCMRLBpKsNMsB/IaVGKiaypfd5CiqPk2Psm4k0v2CzjQ9nUY0VpFzxfO5
56NuSswk0YEUUzz5okOy6PPzgZHuWrMFqB0bdXL2vv3bU/kHYxwKzDS7M4dYYjdBWM54TY9KJbMv
HdemmhWNQOCiLKop52Kyx6p4FTCJRbH5rWzFfo9hJmXWEOzkZbY36bCOb5MeUfK6EG6MHUoydnRh
ZZXbq3NUUvYNpweC5z5d+KB97E5lfQsl+xCosRaUUvcnFOu3i4SUx61Btr3fYQEmHZUHE5M3Mfyn
lruYv2RwnFmAx/O74umqxC4PFIq8f0r4nptGcx13ih4nFL9wKEhS0wPMElFY5jyG5jvB+h0bjqi4
qW5tQJYmtF1FVOgGnhku+lvcRuVc7aFuIPyXDMMv1uj/XwOSlnO4Ixw42VYU0QB3sOc1VQXNPpsh
mBXgmbe4GQ4PD2p8CKEjXbpA0bnsgFCMhuKGZOQTPUTOThO9LdyqcOWT1ulvod7nxEP0vssku6Cl
wJ7Z//tGqOf4gxQVG89TR+tDZVlihcsuirGvaKr0EnkPEZFiRlfPLSg5k1vZ18Rhx196JjKMsIzo
0WP4Kg+qHWpjt60TxJKgw9diY/J5OYXITvaEdXTD/F0/Vo0bK4QTPyxlQB1ZYJIIutzelFyUoAhx
qONVBrk/tOShqEj69rO/pIDMx14iEzRtnAzK5J0lClOoofUU/mF2ky+aDr+9y9BAO4Uj+y59USxa
zxdtyEFftse1HTXMeLYR+8NO1Vi1VFvtTLcHcvGVDKA821sOmmt673KzSdY3epBeCg2XamJZrVRE
aEdjMxUPzO/LK/iiCbG8evkuo2jTTgKrszmaxEzFi4N9jLu+VPPV7J1Aw8d/f7ynKqt5j2fX+J67
+2scKEmb7qcS4N4+FZ11e1a81eoVF6h/oc708dMWqATb9zMAJqF7PrGdJjoKwl4qwUQaYH0fBKaA
ZUflWcEDmzTC9s9C2cc2EwjraHWp8Wkga54DSpnvkUYLLSe2qWTlduxNkBsiRsxNYTAKtYK8LJyQ
uNo2/M0iBqeSvt3z/VbAHcvgpeDn1y32RriJn/8GF7mz99iwDPFbmM188ER1JDOiuL8Zr0lisv4J
uVxdLmXLVuMRWqipJv3sIzYvORsRcaEbH3p22TkoyTDPS8cICYuwp0PQBpQP77KUotPT6FGJWHGn
JbkSLldSs+T8H24ToLdJMQw5x2q6757femjZr2j8JD3W6sEcT02FsqSnhP/wu2GNVGXP3C7j84kS
Wt15pwjNDSLlzrHsA5V8gLmRDJOfliI4GvX2rNcbwaVzrwPPCnbYe65v2eVcVRoK1L4g58t2/52U
+hqPTOIqGhpU7Mrw+zhiBPiMvMcN1oCgquXofTM3Pp2DvSgc/NTRa6uORkp/ocaz1i2CgJ4NJ7PR
BmYlibpFgaStxEK0B6CGcH9bGy1ghhCRahrVsQ1eZ3W7f1z//5GTaPHKr6IXi/nCs6ubLcKQ1m1j
Ot1NQkH3bebe6bE/FBKdKYgfXKJmnwM7kzWHpdaCuElwVcb4lawKfdC2m/VA282KGTWKXMK3yfRe
prZUtgqt6lcCmF7g1fmFMuedIRGN5WYqewMSBPcdBAPJc0Th7YrQw5yXOsXjfBDV5WvFQftQ5nG9
Gkvq+Q2PcNFKTkW/NsTSMj9yWSRyiJDsRdbkkb5fyE4CFGHdmNkHWkUct8U1/QS3m8OtbmQiaDrk
fArFtmgPRzK2mMFv2x+HWkW9HkwTqsBlVgR2GUqhC3cI4/aNzY3KTbeM9S+Uyk/usbyYMU3t9jYO
83pv9CnqB6l+qgluTZQI3aalhgNOJ2ZvBXbYwqKNTwPO2p4Ax3C2Kq5JMof5am2a/Glm6l7YVRFC
chkoKGHFg43SUguYxDLZRUNhMRYZo1x8Y4869EUNyq4T5NpISJ18QRKVxNSugOpGy0yXkLpXznn4
vGoufN48FWtSpF7ToIOzXGtRfufkrLeeH1dTqpWKEP6hlXGdqWGQrRkeooCnvDdyemCF/FFOcPMY
o1jR8Botq4wgo1wTzuNWTeV/L4QCoSSlxpwgiI85qVJxXvZFm0QC9RnSd29VxQxPbN8XJQlSw6Ls
D0Uk0qo=
`protect end_protected

