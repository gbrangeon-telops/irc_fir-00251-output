

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lHZAv/MVAAt3F19GG6CyO2D9ozHTHXUyHUqVqPhHJ9Up8V3v4BMtL2rZCdPHvvrLl9m3lxdPLeMd
yZjuwpNKug==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V11pDh2GdTX922gInHRdE4PGQC5LocLJP7s9hbeXjPbTiX/dPLHGusbEN2B0toY0K8U4vuWNSniM
1aH2SNR2JV5BnhJYTc5D8l2e07TnA0V6ktY1z+NOBfbsIHPai5FO4rlYQdX0gfNxjRiE4WpTGufJ
+8B9yaPmasK5qJ0hmyc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0akrUk3wQb4EqzKkib7F59nSOOeoy+q3qc0fQDYykXO49Ll/FgY0ewL69TWySlFx1Cac/+BCy6vf
iumuPLpTjOS55mFm1JTMxYzM9NsagXEQHLi1lEkcr65/dw7cjFH/RPICXrv18S5beJM408VyZvsr
NCAeZ9gbVAaeGzkHq6VNPIh/P5GGGWEK3241GOn4p1v1t2GkteaDbOSjGK7wX7a4kTfRzrAH+xYH
86BcPdOp3oyEseFdQgL0BZboHxt4zJr0bXL7Ln+oOm7kGCKk4PXPdudDDSsXKQUPtDHqr2MHJwZk
LDVjKe6pX7e2DnCF/lojAxyhWqtc4aJmRRvYWw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P2FMFi4MUNbCcmQEmOw8kkGKpCf5liEfyrVflbrNDPfCQyQhrfO1z3elwJF/eYuRk4Q8ng49IhJM
QbJUTOajY+rTGsCSJpmNj13e1oNpCtCwEA2TBzHdzEyAxDwQ0hUh3ZqnFSNQ0MMnavo9wEIKRylK
MAHL5TjDsmLJG1Zi4ZQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GFuz3jjDcNus13vZfabnTsKTQz9Q9tOYpUUTv0v99miJHiWg9X4Bm37tDSsBPgge2ZWYV/fIZNhM
o9RFowO2ZPIK8CdMOp5y1r9QlxbgxiEVYj1tH56LRgvbv2A1ghGFDDY3Qvyz5G2dmEuSZ/58uAtK
A8Mm1zy2Ln16qChURWHrjkDuCcIOuGQ1GysEn2sqg3E/XWxojTbAmy+LaQrAOqIwoDTGFZ/Ek5fe
49U6fyDbugt8sjMOq32EEkOAQwWmc5uVOZWv3KIDCD6tRxPMIg8J9cwcCTEoanlasaaRs9KqN5go
7g24OWiCSjQz8Pf4KXR9USnCWt9Xh2mPsrZAPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20576)
`protect data_block
QQDut7d1tme+jz5RiB1Y3SFMnzpu2ETaDNItHZaEh5hl16YT3qVs8iRk9H1aBVvbBYiwM49RqXUn
U6o7QaNNG7mXV8aznvmMbrX7e7Vqe+uFQuIGEvMKUh2jqcVzjtaD86UXNlHFtNRY/flpRcX1eNIr
eYZKa0FIm86YHJHZs/3trLeyQlYAgvjNY7d6h+RSK+rEUeiCxi/R4g+cDe46svMJEjSMRJukFCXQ
XiZHZkvVC3g67iz0MM1QNlIeQyuclqlPREWcyRRfAr7EAy6yrP/oKPoIztJggaHupvbb+3Ze0NVH
TzDTm02g7WirpbqVb9KxeEMsJeyPU5THZC14HrS+Z+xJGV/CF+U7vvsBrCKkOvW4psioEC7NO/h7
5pL0vQjb97tKfWnr/tBjlkc2X37TiQumHe9vctI24RcOGNHskNkrTLbMBl9U6sWpZJQ0YVFyCryY
JuVnPIpTm7LUjiiJBCLIZooCy0EB1A5nnpo6y5XYKNF9a8PIQBNJgnM0UokeUjqM4BEbmoI9So5V
DHDT5jUr211nbH0kNPGsclhs1Ta8sAFYV1AQSyIrVwmHgMps30ul6rJEZkqhTYVDAYqPrtLECB6t
v8X7Zm7CF26w3n0x65Srqb/Re/ghntbL8zUWOOXJe+HRB22hmbVX3CGUK/eRREIAiBRkX8TICF+t
8BbKtND40iXw3bfysUnaecslH/Wq7MXbX3CUn/PKcgb6EVgENptknwVO+W4sQYkIvBkcvq7YSDOz
mld/cQGGXiGh9ceGuR1K3Tkhr+TBt+IVIPgdpZJE2aTALVkyAVd3BLk3z6UWq+1j06Ojk4SrafNr
WklSr4YazGWoszj2VKovJaGbHeXXkjzk6BhXs6/j/dWKo4Cfp64uMj9p+2sewfxziEm1okhvSLb3
VIcbUq1ENSJhShbFg8zKVnhyMO0y4Bu6h8IhW+hS0/rGWVG5WXaXlo/zwTfpa0bIZIBOakfME2Ce
WbMGtElgFhTzwy/IxehOMK4glEqVAJ7gEL8KlfJHQmst+ZHOiOkYlDPspq/x84GFyT03GjTdCwYB
BM5Q1Xd5xqVHftU1MR3RAHId1EB0X9pvRgk6RJh0eXUmrkzhXVGnuNjzk7ejfGU10wuk27QpA7cA
oZLFN+qbnV1iQa3gPSFGifN+7PnkZ9Hl6s9Ny4foACRkY8r5rq9j1ZxXuEuFwhTv2L29NQx6W88E
01pikROUxDPV9wyVvzqA35kjD+MgH/HvE6rUmYJ76vBH1nK8txGYcmGE8kHtAeEfrbNFBbv0trdt
+qOpoi0iA+t/Cu4VB6qQO9NmpKGBJi1K0Dk4Hpuzzdo52ZFCHk9LlWJ8XSWJFhWCb6n78vb08aNb
o356Tda1+eZOYhnPosLPZCyyYuM32ldt2umr0rOdFU7lf/h8DGn74nj1Odc5o6G0d8lc8m/kgiNo
kMdzT4lLUa+Ux8HHd5NMESOSxZ80rlIAp8fa3zMHUTmUOQ1ke8d/bjTmrZA8RdzzbjPdQJK2pRFv
3Ws+CCfMWVVwduyYsQHYsoKSHIDNxqNt5yvsD3f/u2LJhfh1leQOZ5biGPk4jM/K8v5shUHgWuBX
H1jESkrr/09fLAqxICQMFLOFe1wIJiEKy36OkZvJ7JJ3zC7ikrAOD5GCXBOEIGUxV7MrPun+19Y4
FIZltV+nneBvZ01iK7fQF5vlY1/A0+9aoqKtYCoMqo2osbm71cm0eRtpjMzxKm9xsTi/SB+VPztk
LOSv1SVy+8I6gTAW/RG4iFQXWRm70C5Psg1ViiIEe1F5Nun8Jpu/GXtIagglWkSPLS9lsIrAO3pO
/WfnxwRifgkTILngqaCYcRJkg9EBWYyjCCXiUypxrmpxaph7mQ6JQV112r/456Nc79ttthfEdC1s
gu/USF1HT+eQ2K8zejQpLHMhmPRW6fN4dKr8yOEKT3d6kqa1q249PKm0lwxgRwupSO56dTKfSovX
BvNocryvcVhlKbdAf8Qhz/zU0r416gCyH5pV9UxyQhme5Fn/LXaMecRlvH8HkiXcB/VLMFMTcPKW
+IKag5S0zEd12y18VrNV1tItPUvChyX71H2Oeqv/cYJ3T1p4wAxDTr7dxCZuU1RiGxgtaoZyhLIX
k7FES+AoP5pb27KtTcYNEi5d2eKjNJGl71urbvA1cdUuxc7d8Cm5kAK18XWNJqLjg09hyUJALbVf
+RSBZMni1orvN175g67JDiOU0Am+JpKHCUamPoteVDtDR4WxOlqnfMVR0LnD8d4OoPWT8RVOgTfg
q5qh2JaGpi2riR2xalAR1noL8cxcelw9NSIGLf5eUG5Uznz9uWRgSAcYUEYHFCA69lLKeZxZAfuH
vlgSReadXMEchBaE+e4fDy97tj6RUO7VyVNf+wo6P3pE5uNKMZGBuzfEKhbT6vNx6rAaodoowoQg
7o9z4iaonWKjyjqeGvF1esf58UBBvkqeg/1sns1gLeAFs8296nf5c+uDYjGBaMG6JzWlDaazDMWa
5Sbg1AActd8uMcTL7NgOizIimE6c06ZSNzDc6x4i7K6Rxaxf1tcya4Ipredi+4vK40jg+rGa805m
hlCg5bc548Qz9XMpnOQlKVTiax4yxcyBA8Xk+IVALl6tVHMK2p+QUrDv0aaxvBMNX8tOFqu4Annj
ZXPBspO52dTJeoZ6eeEvbp4trFvTD1d0+OEnLyjs8azXUiqw3NmI2ammo+c/0XCWM0GPgVN3i/6v
sSFL0soKPvMROYvXq8mzwPS3+dKJNrmPdicVNgu/SaNit4I+EptQbXh+gUV9GIRqVUT04PPppj/N
2TSefFf0WfIMvP1jSiNMiPcx1P80vKC+P6BOPL+ClqwYzx+GpRXwWGRChaeYNQLs42DYsOkMR5Mp
aHuiYKUaEIVvqv4v1F1rne7PU6U1tnw4gajrapZdlfdjSTch6qSvJHjwHgT0YYYAfrA5nhCNo18Q
YX2Tp9sd8D/QDTXVoFeSgJk2An21bDBo9gp5ozYGnNk1vA1I39fYlgjtTRpCBYu9GC5EKlgw8f2t
/57cWb+U+kS6ctsP2T3D3fdkzYFX57xky4wOSsblNA7zxWlL813IDI1cikDbNzD6vCs/WvlfwxFn
UuYx5a5otKbL4arYlyExpsvlyMH+dVdMdXBrUoWyT7R2VfUbHF4WA4pkWbbw8dGmO/iyX+NJYhP/
xD+SkwiqEyd+91fP3Mr1TsJZ8Luf/GZFG+YQiAluiSapqAgT/zt6fCf2CXvNN2IjMXvaq7cgII8u
oJM00TmoTRBIXkoUHxqs7/BcWU7dO9X2UyPmifUpbVFklnun8zysTD1ujxKy/dHQhfJ1WPrflBJM
O2RvItgB3KqGj1ZQoSnFpDqoRjfiKwytD6+hLTDioFbB4kdDkUus8wc70iiipJBvVtAKGv5uGlkd
1rtGcOFV0CIemu4TRMj4qpUnyfjbKSyKWIW0UhXSDi7uTlCrFwF/4DOZzlIac3GMubMiuM6b2nXz
7b8f81QBJM3Q1jL1XvPnHPGtjUe1H9AatvzGzTwrcCJDUbqyoigPStBy7svWPiUN0TsZj1dEu632
XcYOaAlzbEsVKq5FjxBkLK+1vc+MviLoQrhDxDP7aqPqcFvhxDDJfn4qEoe2rOIpF6BVz98c8aZn
NUVpcR01UW8qGHEPJTdjzp3L7jd6II3GWjWKuR1ITj8bq02l/7AsT7rTGq2Vdo7aMB/B26dpJUL3
YHusJzhuEtiInTV0li01vnrzjGtbdfDSpE2pAMwdJXnRyT3d2RA1gMCMR4tVi99OKF3Idn1BJAcv
wT2OZdIBqrhxxFXNXeSHWwQEus7mA+KIdrmhYx2EpoXRtOWvclD3EwY0SbH43QCgKzPK1O1vLRN6
HgCCbgqBR5JMHWq4Dt54uke372dS8Rla0zMfFUppymUN7Z3pmlhBF97a2UVikgisF4wLuH5xmYO/
iHoZZUe1+KR3W0FKQmnl0HHD65x2RljDmEEh8e9fTgTdwmY3Ra4hh3X4cV6+DTy3YJGB5jfYEhYc
7J32iLNSuKy4eVxWvjGakxdH6MHQ4yKtK8t2vpE5QZLS3K2QGqn/kkOmIzZgwKTU9MkEmzU1LKei
zAgaWNMfXXr5NOY0PMrQlXp7VSArI9ttIG5fJ5G0Q3+PyHhVS0o9pdRTf3vEUIhee3htK0lOvyOj
l9vYZm0CYoFxZKfGwZ00Zo7SzzkGJPbOCpXRcXJZLEcZtH44zPBDGyi12cl0xTEx2dV4enOmzHJy
TG66taaj1lEKYC2Sn9Yh5HA0Aq32h8kdKS8foViDeLF8DB26A8URvH+Z4emb79H8fSb6Ot4mO4NX
W+VzBvQvCLpY8c4/JWThbLUpzhkcp4+44O9vMAmRUEUjaM6DjVT6fmHl7YWZgb63lF2RtMFIiwu/
hOTWBBI0QR9f72Tpz1y5rBkBNjSz5QSdgH9iFH7019Xr1Eep4qrIWmv+XYcA80XYByWNgNB0CfRW
a6yc1+bbe6hE2Eq5Tr05SBkgigmdU/K0v5GWZ8PPorqZeYBxuCtXFuIOGZBIbBREDB8vLbrP+lmc
zmwrG/ZiB1Nb79W1lEkEZINWu6xs3axivHefxW8OohDwn6QyQD5oMOGIdYOfzQEbOlUFZ5kotsyb
AFJT28hJO21h2ZArvZ3jVCx8ZtaGUlN537QN3JpQpboVGVbgvc+E2sjVqRygBrQ+NP/eHFiWVg7y
s6ygIHL0U5lF2j27x6hs8ktQ2PVy27KIyF7NnzQJstYvusuki9yIqjfdP32LlnvUGyn02t2W2bui
jTv4XmQFlkmXlkJWTs+hp0ZBozWwL/SqwnuPXpZ3/z9PiRVUouRapJSp0X5Zq6KaDQqOkHAi0fxc
QlekwlPghwm3Gkmd4VRdciXq0RQ7cSY5WJm2N6ge9vbLM9fyp8gSEqWw+CL44FRfYus3dkX4cO+U
dFQDitTpMLQUv1Q/LMLBvdr9bpArFReX4oNwTsPp3gyj4k9Ts9LCkeySnwFj5jOIGgeHhAZggv4L
wOvUGIQivB4L/xrZDsMv48gBH+1M86vaPyzXvVafQ9WKgBkRndmz41TUOa7MOHon4roryOM870Hn
kz7qYu11lpOyu/cXvy4AuiPCa9NoThM5ufy/Gyco45LgSj7f7yJ8TVv8dDO8aYw27JS6hVnHe5Ql
CbiMymPU33/5luOEDwOmQZyox82zOIWihnclzB8ep0xl4HdgL2AKOB4cVykl5QMu3c8hEu6z4km3
e2IP8ldko468dMYLagssZjsEzp3KwjuqMFo/qPduA6/9WJa2Pa6T4N/C6Do9cwlbM/98+FVam39y
BC1jJ96vYcWGFDDWTZUnzakGt8AmV0UloGE2FxvykSzOUUpoXGABu6uyAiUlJRU9IWlQm6INBPzV
canmmwGPE2ZWqkRWFfbrTQU+wNUo+qbSVlnMt05YG+QH6XbDyc+5lHQoJMo683yjjI20RwlVHUoL
OIVrUjPpfryNcXAhmY8D7w4HUSaw9VTzm6MSwhbz8hS0k00qHa+ZtkOPJByod9OT+GkOX1Aqt1i4
ENs+gR8SovBdr4KtQ/EXFOMRT+ijLBnFwCDJTXLTr7pdf3UeIvU/Lc156TD7EQ8GZNj8+DTf6Q6W
l+E2Jlqrw0fTpcJignVHNoyzkpK06UqR/d3WoCvShyE/mZViOshrq/W1JrqofbxaXGS2ok6y7hQQ
deKdSYbVQy1T3cctTu/DL6q57i0z9oNKgIGgC+nvuJi0FBtsWuwlIEohQHPPZhgKxufZXBaVId9R
+Cf5odLwLU8HrAmcAryq8QIZbOqQ8Y9usyM2KuefiFWnTS3rKK39aOwT7s6/59Ki/c0qAT042lnQ
3DpCVmbCDzZmKqsYFAzrXepRxnPazW8NT38kHDpIqFaPkc3VYge5kZRm+VeamL/ml5UcslHkh8Yy
jky5ORNMe9OxP15QCwEHtE4z6sjf9qbdewdujyRJdnoM4GdCyifI/hRPvcHtm1olK8SefzQkL6vv
50V+JAAWAcCChA66v6/gMJwGbAm8thoNngklA1erNouKEMeKyXzhFo3/kEXwZanHrYySIWSG9EP2
2nYrRBTZ/5CGVpi6cq2NTD4UF1QSe/4nVX7kGXAyYg3+FNjQ1qGTi60L4t54xuuF026oemMI265O
fz/sVKqU/zq7bZswcAWXRhXT4LF/+E5OcZPmHQFU/h3Ac0tMdKVj2JoGzSfXCHwomN8jiv4Jk78J
y+ZBh+u2rS91V7l5vucYQikKDNmDAy7NSrfDnOHif/nh8u6xNRGfhbUzuWuNWx1tYa2xPnNSgFL5
iP4ibIbLx49sxCk4sW9TdAPOukHUDF8VweUiMgI/a01NUxRD14RECUkiDM88zih1ULNXRg/MM/jU
iSoWsDc3fWTfp9ABvwYo9x+E01waprT0gAN8+2YNj8Djam2dKvtI0ZU0aT6kgLyC9AbCxzMw0SQk
etzgK//GQA5+elGkNoXr6UpDsrvtEwxvC1njxWb31A+yEDIhs+h6mgryULQAd8AKd5ptolyYF86w
4cpQOT0DIWDt3BNYsF7Nw3NvtT6pdrayb2sMnqbhM3ajhJ+ZMykDIHbZEJIEjMXtRuVhCbR0xpdD
lCz1WQNY6rFf+p9EFu81dB8EKFm2zpzYx5TBAL/mwyOUmagqTE1j4Gslq49UJ9HJad7/Wzg6XTJZ
QSoRIbCxd9H0Bc2LWpPsNQZBBcYtdlnZ2ysK2g+w0ZLsPKcRV0Z741VP50DOhiC7/mVPJKINZpQF
5rC24+6VZHBB5N1xwuW7Q3HgHgkYHhWHUwO9o+7+UStZLoBSiVfHUDoIG8lG7vNQpHlTI1WMrbpO
iF/I06MIQ/mQ1VjXl+5FdZWaGMpK1L4eILZf87eGYTLGlwJ78eKLsrIbNRz74iRs4OXIuTnAlnph
bpWrZqW85BPUlSBqUo1izgjKjLOKNJYFTOKFzDgCeN8s9R4lma9zWKxIFIRKGTf8sjBKTDgbxuu0
wGjJobbzibRkgblMe3Wr0iEM4pa9G46EylV7OUV4solcVZm1dMqmciBEmxxbmyB/msu6Wwdyx0rG
VpA6rZ4ficfvwIoSSdrO0/JB8LnXDzmFEL87hO8bB888JLvjcUl0wP3x/EG6iNXyQ9mpv3XszFg9
5zvm3UdobcdHgIiwKZd988dkv2IWUYi/ifgbq9pK3BgFXrKybn9lKDNBxiRgIWXX5TtvwX9RQDtg
KIGOcBKBflNXI+UunkXEswnkYbV1qp2AXKjrxnT8hGGNvYNwmEL8PNZi9Hm5SqExQXKWNrJE3nDL
q6rhh27Hw2HuhOfHTP75of2v/zMxKdRyI18a+j0Ze4YuYz4jVE4oi/gkDN4Ik8LNztE3J77+j89j
D6TGHwWyGu1rNL9xSaP0uEjDRRuvezGv8u/1yojPyI3YilF20F6qg2VFp7oSZh9FEdFl23Wnt2Gj
AGydbvNFrBJXPzxZIhPpTE8LmerOoe4XrzeMWT6WzkLfFoSc2vLGtOx/3w1Xh0CsqySeMNgOqoGC
NokMCAq4iMLogX6RC2rnCV3m7eSqP4uqVFq4A0p8j2nx5Qj5K8T9djqGavCjFofnV4oyVbR0nbUJ
FdCrXp84zIKeKw9LNfebN3hDN0SVLdLrOUrPtxxB60dm9/JCdcz/hIk8Ut1k4/TPl4CyyHzAgevY
PV/dx+TQDRpQFqcyO7DvBq/MIkoOLoEUD9DwS71/w/j90AJeRvf5t9rLXLk/YB2ZqcOxtYysJVQ7
fa7UQPRnjPjCTiIEMaJEN/7v6UFrMwyCz6Fk8THpwEJNoAu5Eig91RgpDqYx/GvAVqI1Jq5999zZ
+ofmm4iR3W44hRGL6KXYRP6ZS4L+BeB8owr5ELiHDL1Tc84kxUqGDCXZWWruc/GvcwJp+1+g034/
FjVBQg7WXRQXZUtrZumM30lAfmIRyVyMNvKGqCA2HjkcjYntQ+araND9nhP9nhiegY4RJddP7jEc
H4uzWJYNmzyrpradW10fUHE2ytoO+S2g2Krs9zm21eVoNNizDvv2+OqNGckdtwrn5YdfXjrtN7/6
9/D8oNAygC6XvDYuHvMxlaQwhXGUTXfdd0A7zou2nmN7AHVbyH9qheY1LiAKlRlnZbdeYVzWPpvE
G2NzL1qeYn4Ije+K3Yl25/yLdHDsd6+iVo3CpparZCq/guDFOl2XZmf1x3hmqBQJvjtcS8T5miVN
48a/fboxNbUX8OYDmkK/tpxsc1GPEhi9IFfmJkM5K+aT54/qdsuzHsM9VviZtnPiLQZAhDEQKNt7
lvPGimvM8Wdva6mecZIN7x5JnOi4MI68cSBsurVCa/vLYFZJ+/kVORvkmdPJUGrypDrZ6JgOBiWm
R1eIaAZl7OidVRbo3A3+ly31xPobi8W48Avz9Qh0W4nb7ouFWuLfR1n2ExH0L+9IVKMODzz2T/Dd
XHANyZMQmGix7ato+AnDX6G4ha3KuZPoOqzpB2MwEbGOv065UzgayvyNNaIKtcBFlGuAAqnwMDCl
KoO2rf0pcltiEnwx/RX7cIyLG+4cPTHn8rD6/fFFr22ILkkLUUU/VaLe775pqoDnXg1QmW6Q2DvX
o/PY0DgAodzrEFLOleqLur4X1pl1vLWVoBdu9eZZrH220WjFOB/EEColZ6KxuxSxA//65tqeQmkH
zisOcdGbzON6qLG6RnTIwB8Cg7aLjbIubHcCcgkX5s/OoMU2oMFtGB2AK4voyiwyzsptyL7miqDY
9kMY7UuKgBFpbRg9AEWLn+YBr3/FPKdG6fBQFCD8UV4tCJ0IijyvSM/mEo8MLeFoBkUqdFeakdSn
2nlaJJm4QXzsp53QuhIFkd7VhGd54jPNCK6T5JKZ/B3GB3Mx57WKH6s3vkeoP5+rTrqrNwCVipow
rqLJBkWHVu3EUAB5HIW8UzZjZjDIFRbBWNaLqvCV0Obb+jZWdXUvc46G+pODREehBfePukOzDYkp
ZD+zn90dwTiuCbo8RM0Kg/doh+/eX7TnUL32CT+gJlyJj+z2xfz3FW2ZtNlzU1AmveHOskHzjMOw
J38mmOHujI8x4L9y69YzOSIXfqe73l3SKs1PtS+t8mkfdvSWD5MZh1ryVOuQot3TXiLIFYAfKGFi
fFyvPeCQRRPJ198XgpsuELnNMNtn8HK0VZnbF7yGL0akRh2SSheq2o4uU05zvxp4jpFtlaSyngsT
9UPq76/oybDeqDvI8WdBQSWm18TDuAWUJHbW9PHajcnYZKz59+XyBjrNqjGf4ACD+87TCKAj1H1j
VBX2ycw7y36KPdwUqGbRsqP4MqaL2X0WNeGcqXZCH8fLX8/rEGOw+eI86hCDteiGjlUZ5Uz+xiVA
Vfxb2JQKotVYYlx3jXjYtqrI9JnQwh2fd0PVXoxhD/DvUoMXU5wmjUxx3JZfvPi1xqOwirKsXalY
MTMH8QxKF44+DcKFESLAomn/syUpikXDC2rr49HbMScozQs6FwgA2XFG5xWAd3o7asAWvWzyWT5J
GCSgvE8SR/5jwV3MRiQ7aoeiU3IQULDZh9wVk8p9CQk5vuHxABslo9kARhqidLl25thd/e3iDnCq
2YxbLvOcnuIWHus56S0Vm+AeMTL3oeu8EtkjYVumF2IDStaIGH0zcDzpZTZQOfmhsOCk+ez23s4r
2f4dNuc+PaJFmpI+hXZxs3i8FVWny3vVNQ4ZRCyyFtMllQZ4BADIV7ROxUsuMEIRWUIK5o9DnVFq
IB1qNbxfonuXSH3ZbwX8NR+1kyvlpKUeIgNswnlYg2PWVPUaVHJjqgxFShFS0tmeZYDQl3SinuRk
YFVsdTwVhf5KW242KFyucDH8h704RAvrTvlnjU6CCv8jnKB7Z2s/RTgaV9PNFVLfvb5S0xKlv3ij
A1lIXzQQgivClJSSWc8SURUKIwA/XBhY7Z/yeQ4+z72rzIq7T0cNrlNom3F1gvvqg5ziirgtHDT8
xRgnuyGFJDACS3gtnUkhR8mW8bZ55X2J5sLq1Lr2iUfM7uWOlvVFrYDGYXBAXKt8vIlhXHvKJ9Y/
PjrKEGQmnyAE+hHG5p1uX2TiCvf3sGKpNUI6mYA/Fby6oBb1IN3qteWijsHKr0Csoec4AuMCdTNf
VuZWbmY/35rtlyyRk8UwXMN+966bSLCBvcar6BTY0d6FX5Wldgqe0lLXqgowjRfqDK1ZW7EJ9r3M
5hXUjymU5RIGDr1maHO/3X7R/YFH9U/l20vWioNNSY9LY+ddFUb7Rvr5JFOQecaGGoBXwJiiTTv6
xP559d4TxldPT9532PPtn7wPGFwXT/vNzagfh5LBYbvZCMvwmuzviGaP/Pnw7EpkBkVtatlO5w9P
lJMaGiRKpVQJab9VS5//FM8+4QgQD2201bo2QWl0TXC+MQ9cOrDEF7e4rXwyE2nXW+FbVdqPTTmg
pUX4cEtZqdS1FP4c177Z5Ycm7Qf8xkBWj4IWZv2Nqw3bsmKmbMU34Xf8s79IztAMlzcZTQZb5M9K
rJkMVGlOMg3z9VysHxn7+PHQ+Cvkrh8K/PiSTpnkTYqUIuL1bOYZsN/2Y8OiENFu4z883QZPYYDj
0GgDKoc1BPwMQHJK4FXRarnRd/Uh8OpXnKJYbsaThuKsgB6JL8apTN04pflHcUjifUI9knVBqF0C
nBc8YJ13MbzsF0xRXoC72xZ08zpeg0W883xIViqkBBrtrptLiodHs5DrZA56R3Dk2nVhFPrxqYWc
Ot02EnAjBHBBM0+jIZbmgmj7EvbBQXl13yAX+mxDevbpj22Pol8Qgub7ECR/q64mcypPoB7/HSZl
0pYy+8so0U1d/Xc99hMY03hlpyZcA1n0r932vm4DBx3kNE5i9P39ZB2EwCIce85flZqbmXYwlHFv
dPQAPKq8/v2Wx5pY56Qn7F5Hix/UgkpmYaZMVP6gWMY+w1ACOGaxhzZZdLB9rcr7Fwobr+L2ajtM
jE2XZ6QNMKChZJ9Rv6m23vrRQyXX/ysD/KucRNnPHi5N0t2FdRHxu2tWEa1khpoyNm/bG1U7qd6N
HA4jeHhfbN40PZcqx3498dI8EGswykB1q2bxXW448Kg3M5sN6o6z08vubVmPC8+4H66VxP4c9BvE
Wg8F6HDY4FL/w4ZKrAu+Bp6qlg/56MGQRad4Ewk8BtoIkjdDLSk0Xb7LR1RavbJA5ym+ZJKGAedI
iF7sJ8MGIgZ+FKLySKXoFq66up/iBN0pADGx6Mw5Tg0C1AsK+XOYT8akj/z74V90yXwDElXq16Ag
3aQrK19nfgcfVWB2l27ikexaZDAHJMNugdf4ZFLs3rskJJdSC7/BBY2gRxqlsTeoHNQm+sS0LrCW
S5u7q/YqYYg1ZQhnRXrJ52WqQz/NU2zrhULadkm03Jg4FNHpqv2TS+VoSaYkWmuT2c9t1VdzrgDh
cmF8bwqOn+VysUtOsl0G0OawQEVo1fBSCFUoGa/2XkgdI9KT6I2nvVLfbAcduXaIvPkiszqWXHUb
pWHqPoJgF4vNI1BS2dfJpoiFIoVcWoI56A66P4EMzXIFOu0UgehAIMFXfPJ37i78wYEn8uv5vv4l
Foj3wN9bztmj5uePsevmBXlFMEM79M1Y2/lIV7OSa91hBxlkneZNJV33oxMQTB2bPIUD9euT09Ij
jBzoYKyQglfFyO385rL92QKq11M09yLnh7yHf8Qz5I2ctL0Lj/Cnv9XLn8elvD3Nas7Bn4iXadjx
zhodezYnpF5QS3XCHpB2PlGS7AH13WEMohIplaJw16Dk0P85De/R5PRklfShkJnRxOD3R3Do5cQg
GL8rygz+p/gwhRdCWAEGcGSrTb1rFIZZlHiz6CJP6LWCsH3t/N7ZRqz6pi8pHM+Tj4tKsSiq83dl
rwN3HDFlTR3fPVzOjSbhfa5ubXu8tfuTV+Lg/JuWB/nCImcxMT0+BSbGmAXdnxsor1SvwKt7uFw5
upf87L1cOUxHHT/jXtPc/qI23DRXH3wzH9znissXBPHD0BAFVua3YhEC6GbbB09QMwsqzU9C7y8/
aIntWyyBIUXZTZhfqzX5J3t37B9CsUaBs42kDbButw37x1OAk4UZlwbY4Qan7Y8qJ22WG82eG40A
ja6eUbIflUCtx3cNUhY7ZPkcF2D6XLV6ECn6ilv/LIhmJVWg+a5n9CXw5APWiSFRIEm83IJsa5/J
wi02/Yh2e3Bt75iDkEguqijhdIZCgicasUlvKswkWBicqjyPLmYwTWKf7Hck7XREVuQN+KKh0VBV
s0eO1a6G6hWWQb+wHrGUMGyCWlU0nnBI8UnVWvOfx56lcPo1fMlt2O+SyQ980JazARCMFTEIfl1q
xbwBpKaqbXVMt2amTHSvSDQpPnfUAGlfLv0PL0ZkrbbiusjR2I725fyWD5LDmGrRqNkWpAVU/bOt
n1C15NewCnse3Bk/sIyZT1gqz+8nxNVoeuinGzlU7CfJWCli/g4ETfbVSuq1B0fRI1sO8bVjArf/
3i8Q4r383A7V6bbG/jkQeRZKfDMqxy+c2P4uSglRKIb7Ct9YRIWkB32xom5/hnwpXfsdMJ8chR4j
uxYbdk8usYuoy+o5ytPGpIPqG7XmfOF8lWbDhvDPGAD5YY/7syNOXvxJuRlEdhb0AHbSlzYNbV5m
CTkTVj/K629EU6W+nAhyRsdSRha4aXhbXmxhqChqPRA7WDFpSdRNQlux/znag9VlLfd7pB5u27Sv
yyLpOjyhQvFRrNFvtimlSZceHgUzkYNKLqj3BPrZXDxqVn5PNAl+BiVGWh/0pwlnIQLFf29wh1Zz
NRWZ7wfFQNhQU0II6Dcg7o7p7EWG2iCzL0dAdku+/2W/dSewntqxQaJjDEDocLcZ8+mH6jEGAC4W
9q4O4glTNRV/93v3MBcNl9L9ELKTD0S1zXnsxxZpsb+njgOS7T/+QVXMti4ehAp9fTxx/yBde1Ox
LSpojAo+GeUOQLJd42oPU8GUEFgNwbmv1zJxPqswfVrVKFqSQge2LWMQqYTlMPJLaY0dknKEdImI
fpxy7rjoc8WdBaism0p9F3MQ6woyjnpJwjnBk8AmuyTJzGCpyJ0NnVpjjI3V3wvRW8kZwDilPbEQ
RSOUOCIRVlOnGOZO/W+dxz7Uwo0AyxWvxQmxR+CCp9W+rgSHkJFmRUaCXJE4loOMZOafyI+4/MLt
XSPHNXNP2l9AqbbGQHiCynyym7x81sRaJxU3UU9ixkhNWR3Pzt1mclFZfyLctC7tCdTjVeNDlKB0
UFDcsHJK30NMSPr2wNrsRdI75YhwntgjNOl5AACss7j1a6aHZnR98CwWGwdSSRAHuvtl6P5LdJ9j
ycUSqdoxa2+YtVxTcaTDp6+xLA2mFWsHHSkgNhOMkseJZdpjT3A75RFRwV9a3EU3DPcad6Gh/+zB
vR/92qmILxHhw0Tda9okOR3yG5fJp9WOcfjsSKuqmop6jiNlqXi7JQL9QvJ1a6ulGDsqSGpEVMlo
iNub5YSrKDwyIfyzBmgZCmT2d0tkoNZvgzg43qsHIrg+6dtKCJ//w1wKVC9ue9mAQpZ6nlcahsF8
/qxufLG75BMCLgE8Kdbchx5KAAhikO5FPc8i/+sE29OqzFC3hqBNxmJisEXVRu3ZKqOhFCMisa5w
xcVm4eP4Dn6/bMuP035FkrYPYnQF33FqtJ4EKRWqBzgFN36Hk225QVUPeuBReojxmjlhGoFanbQ8
kJnWEP1SOnAw7YQGYSQTZob+0esQvx9Muusnhblj1Poapdxc8gZNnniDh+tnwm1WODsIzFnBdP8U
Kinvh/+qGFOKc/lWKIFDaG5N/bWKG2+DjjopLKGesY/jFjZpnQUd88MlCWtus7pEw7kVVlG13anR
IXKaOgWuX1PqRmzZ/rAmrw8NN+PNHYYjBTA2rFq1d2ytfDXin3r841WAu7bN3Q/a+52Rhmw2+npk
7amQgIgdG0HLM0zzPnAtKn3E1gDA/N11H4xd+lGjNh9wUorXsB9a6LKUfhNPFQS0R5AwrZbWkFxO
UMLZARadR+8oqSnn7FrSTlBmrMOgC4z8vk0V/TuMqshL4rM9e1zlmdfNT/x2YKu1DhjimX+3j71k
ZwAMlTzWx5F29ihEEzlNXLi9STNp9YUaRrxDIJn8PB+ZuPMuQD1kUiam93Lkxc3ItCfoW/JZ8Bdy
IDdbN+INALMPzqtHbzZ5pqGQUhHrqXZhHz1wYIdRf3JFGiakubAgw1j5Sus85WcBAkbPKLrTsfGO
yilV8QnIrD2Ev5JWvU6rrdkA0ddP9BbIVBirCqRJagQFkY8Q0/OgVgSbUaxdZhAsYS2F+1Oh6fV1
6AaifcHCLYXAhoMMUcfHZkcyw1GgT7hlZAPdAaUFS4cHrmBHwjMH3ie89AdBG1LrlzKT4vs67Z4R
yTQ7FaGcNmGXlvHJ6T/KLc/CUV+sd6r70gI7ysD7ENYKDSQ2aKFhYnZkmVReuoIj74xEiuVhbw9b
Wk6Yy3NwGvZlQhzshSi3BD93B8C41YnpPDgGmV5MNn58d2/kKH9kVdpjFDpl4vLMAOFRUzeiX7C7
28cXgscMAcXm82TKaPxq4Cji5wlaxfHvwb2b3pQv5lVu5QAVSyGCiVnf9IYiF55lmAdiJ97HkWaP
g0SA0Vb+fYh0SjKgMK1Mi5RD7DR3ZBftntJboyka7hVqdYml3/7f++ArWqa6nZ9ZKDI1FFAPzia6
AJcIamUd3BiwuAFWz02LWtlBrMMUDxif6OM9ZhujJM03sCLSl51Tz12+AESmkaNHYDWmMsOZEcUV
vTruZ7C1MSg6y2q0GtmD7Jp8lbhkp0Yv0Hxqre63WNEedjBYz/XStQ3ArGzxrra3ajp2T6n4MuVZ
KN08hKmgzuvngJPoCm1kSmBkottfShcvupn2CTPW47IsbUI4E/ULC8Inf94ERYwSjvSwt9SnIGBI
idmlNMmCbmx3Q8ye3s2UsfzvVLsanYFLkNTlu+YyFkuEehS5zHIP3tfrjaqVAXnZw9vi7ggFD8IW
8vsARxBTT0ISJnkcvBRI14sQ7wMJlPf6cUeeB1fdaBIuZAvZWhHnzBnH/DgMpClkT3pYq+2DQpl1
t/T1jJeGXfY1tVC+pRGXTIDwumZnpQ6/9wi40uPutH6fEVvBN+CDE8WLryAoS+RPYfRdv4mbinNt
zYPwJh2358UbwyX+ORO0M6Ulr2fK1EQz8WNTEBeqhLet29j5vpUl4zqeyP3bI3GihUmb8JJfawCK
R1fxmgLtu2N4CjabzU+BSYhgeEAF6S10H1NUE7LTypjxWOp8L4shRSM3nlk8UCAaNEFm26XKHgWf
0ALEw/PmRS3bBEFK/FoAVKTGVcrVBLjc08KXGnxHIFcHeW1p2YQL9qFPJInmZcNOqNcRtk7usUKh
j2hMQc4OUhIoaZbrl8vTkAH1v0V7Fs8cbHctcs3EFY3SRtZX7lwQOS+NgXIIuOWfkQM7oiViN5tL
jDh9wJLs7mCnQmN9n0B5Q8D0DGh4d1uskkoB/Vj9YC4ONhd4UbgsRkOXyJII5gnp8BsVth2N9vBs
ev9PldI7MM1WpAMOjBufd0HvbsCAq/fuAWr8xVB9NrRMpuaIYzDhPMvfFfgweZAfzMiN15D3TOWs
sBwx9EsBvZFfrIbITLSIy6ykLOSW8/I3DhxHWmJUiVJYt2eUqUxiCyDQBALGA6hJ/podPXsLq/yn
6WfyfFcAQk6+l0YVgrzwB8uHbq3BZkKbwu+g0hA5U/+uNlImicVqfN8b3rhSzcCdOLcqzSh/J+sg
HwM7yBE837uyDsTit63sh9KFV486xK5MwpTAqAJTPxXgrPK88NM4K2chC1VEPMDIKljplw/WWmG0
ZQ16x2n6QrX0qRI5nzkj9WBjbFedQCJ9xWeKmRCOgyxlpe/bOqk74bobJX1oBmQsoybZ9BOQu8w5
wYOUS8yylG/Oxmjk5MXY/nUS1KGsZF2O/cmIC3CA2Hma+Ep2djDJ2R+szqk/gWrrmvmeCrdvCs7q
NO+N3QzqpRQsC9rrKJl+b+tD42NOHG4nN1rMxj6Bd+/hSnkzhsv6uJgMg9+T+PInQjqjXTPQ2ORN
7uIsLh2xuKaoZoGHT2DlEwIriJd/LQuKVbZfwqWhTautU3uSAEkhhufZSDa6frAppdxJYmWs/Vk9
tul3fvbrPOVk1Nj2dgTe6za5FiyPWrU5SrVHy3a8wEO9j679udygm9G0XCyS9BwbIqhbuVCX7HQl
MFpu48AUALJgc7THRy+IpZexNFN9H8uAZhHNyb8EC7okIHDVx5o0WALxWQ2pinK8lhfhd64J+xrz
95UdXkM8TO6elQkJBkaX9CwwMvysTOCMKsZvHBvJZayPaFbD71S2N76bi0OCf737kB4RcKbn2dOd
6s/4qPJUXgZK4EZ4EMZegoxszDtGpwMGm93oy9ITstUbLjC0XixbJxabhtuBM2dzQv5p/UwUgVOZ
cOFacLfsc18wWODFoUoVelKTt3lBUssdPdYRGIEiLk+5k6yvLpjQcvbr3w0hYUMbMXaQF79eqC40
gtzLt01iupB1OsN0dBWgz/sK2zzFMDNdkgX0Sth79pCE7TKTX7cGX3bBy7ZvSg40A8UcdtJmd5yd
qCvlA6lDIWGlxdCuNR9dzPvdrP8jnG+cBJZQf2Tnm74rzNoj5j071VbNKSW3yg7kSgjnBG+PMF37
PfmOIsSZWTJRfVc/gRKrHJL8A7LiFsDy11rv3+U+nwBL7NM1tKEA3lFScKZX5olWIzXoJODaA4Y5
dOjkpdWpaScDKU63UvCh9epPAvCYXQq69jTGdPkL5HYVjzOPSOA83nvKgRqmym3rNyCRbPz6yuxl
4u00nOXjZ+/CBxWyqSyv9GDk+3KTLEfukGuiAdqhjPoNbSDXXtnf3Qg4jnBgDHk2v9YL1tmSCSuQ
UqDCnH/twbZMPMv+5iVg7xj25BufB9yuv/jw1SRJ/dNimfekNeBI0JG9QMVyusapa/d1YABAftE2
TNq57/5HZpM/mj/IQE3m16psXrQuh9alDFE/T7zEFvGorE0hIo3fNdvSGk4/Uv93tyfI/W38bWHm
uCfPnvHPtKjdmDncVR9jCQc8B/20oeaGwY5Mwoq/Vuv3W5SvnN+YCaLbH8ejvzEgFp/QZZ/HJMZC
ZGovQzVoav7uUSu+liYQ8/ndK2fFE+/p4zuyq/ZW37dqMJLjER72dnRhcDNnLXJ3RlogyGuSB1UY
NfLxAuFIaAjfsrSBmM0rmATJrDaoUkfydJVvsHYkq3oE18a0hJf5btHXR+G7yxnnbm24dhVDgaR6
7352yHc+vMiEikoXIYgF+UQ+GqyPZmVR+fRo5eOUEE/GUdw8ifAXEnXZX2qtIVcrjdCl7EzsK8BA
R0qtwvRaLXOfNtViPic6yu31Qw9r2TXrDDtX/XEVI218EsYU1mpOuWo7WYSiSqlm4lZSNb7xcToQ
+qqe3PZ/a8TRjnd8zWJU7bJ3VzIeGBzLtJyIoNPBFmNkXzSLWCjar2IgaE2en7OJXWbTnDshULb7
2iEHoUm4vZMBx8cB9vERdFDXLVJO3q3KsEmjyWndCUad3G7w8SwxSDSC8vhwzQ6gyrntX6O+PWpT
irarL18qlWfu6tTtn++hIu7xcJP8GS9ocO3+4BJX65bZ/xK0f/rtUHzytR3QW1zkfnm/87pPt5hn
IyNSwppoh4iEbRS7m1VjyYFf5VzOoztmcnapjkwvmmYt9/ZWLOIyJF28zscAgwaJsMiuN+nRAiSp
a5OKE+tR+kdGJ3CHfSv4jyVpT8M0OOZF4jZQQqhjzxbflXUIEe4EaJnWrlE3W6nzJV0c9iwiPwuF
x6JLOXUgOsM1dwd8kbore/zwahvKARC8oHOo0EBHcXxtXdu/2NCQ/jyQCgpBOi7J4jOt7I+ru53U
8nuTSnLDJIMJ2p8PvbkiHS71U3vKOAqRQG8ohT9uC3YWTRu5ZXn60mcU+6QCc7kZOKsaj96J3VXx
QC3PmUgiPAwSSnTU9Y0qR/XZJtBH2Gv7EShjWLo4CE6ED7IjJeFjyFHZmQ8fbbW6hz7PVMjAlTjC
OpYrwNF9S3ur0wJqaJmSaaM2RKDL7deFDTQBxjs7pYvvjKHIzuJoEq0cd34xlsId03aqlRk6quMZ
DsVQm3rkTA7wiG+z43z6pOa+LFspfCrkqAN8cMuXdew3WGeIN4eE3MjQaeLYOoh+vaCbG8TN6g/z
FhocTSS4h/zuxHMVtcaUbRPh/Jgis9+/wLUqPrkkXW4NzwSwP9HIgTOtnkLNYRRyaQJtdzRRlz0S
6L6/+3HKnibQhlzxT30Mqz1d9xx2YzVp6eN/MnlhMP7wtvkgEO6iupCrHJ/XfUg6fIrTfUmyNgrJ
pk0/U1JLoQo13nNNOrrFTMMOTrH6K59T2PR+mFAdi78yRqH6AlUM74jlefTTEt+Hko9kk8uB1HJ2
agBOuWLKNxSnUOA7/SI3ZteRjAUDUZB3SXBEn5tYwuX75xZ6FS8cR2fqg4479kJ4VHgEctjEXSLU
eonsBC5nI/EXDKbpaenxFT+aUNqfAcDsUTGCLLEXHJUqyhETOwFd5MqYIWjRZ2HNJyEnYPjUV7qI
9ahswHx1jhX3ytScTJY0lpT9QgNYi3Cz3XT68yqG7wW08nMmT3sJ3ryFbcdVeS2hCpGBWPPE3ILZ
H8kKmrGN8fk1aFOmmuZwJjAcKTUyV+P18xNHFmOxyeh4BQhDydA5QHn68S8qaW8v2DYx7Zv12upg
DkKfhy6OqxuocXMlXxyi/hsXWuDjfVV1UauixYlfuyulUslEcW4VIFknPd/qQLsaN1EMTdHYuzDT
u8rZwbdpPLmjlnjIdYBlPee8dBEJyXUSB1V7YSMzRj9FUGGRFCn/Fy8oT6tVifPwiNVsCFQ+XRM/
CoIl3HRj4p46ZaehtM/JtDvMRa5mQaHjVLS1ZjrFFsKim+pax5EGhvh9HvbjRyUCCrcvN/dyf1lT
zrE2huSP4/eFBgdsOEGm5+ELJfupCURztiC3MGsFz5xClRYNtnErpvDbUM82Pk0ynIKodnNOKXW3
eQQZv0P3PGbfZgZOjiLZxIl+VDeTtOZ59jASfVW5u7kdfCqU19Nnxb6Qu4fbVE0YLhKx4AMXg+8n
3iVWFhTKdOc/I6TeQmBZvCTuv/fVYnEX42nzfefFMtE4YlrpUSvcv6/l1dulu4e+fTDxeDt+9boK
uu8XwwwZV84fqg7K77d5SIawBqMxlB2bF0+pyy1C3PJeYebUZ5Gncm3fwWqQ5Pof1sXdfixK3a2o
cKsqeSsFaA5KO07siWb5Wr1HawccKbEmuNNT16B1TfzEfwHPP2/t7iL8QQGqyIixswDRpeB65DNC
e7mN7DoOJ0GZ5xbE+MfXWxE+6qh90v1++/rcoxm61tZ6W5aTyUZlaoyEkQleJyM/keDs6o4EVvqA
xSs/VfNv7lMJfwX1WHaRQEfFcFHj0SJ1P50s3ZUedYpIJrsXPiw4J4DEaJ5+13BmCnGIKPAE5x1x
ltWwoCSnzd7DKBB5U9uclMSJaZwff9MgIbCq0sqXHpXscMMIDehKBo7FYYJyNDCPOFG9UoAyU0oe
VulBoOLpuU9Iva0sF2dNOTsg0UWWwagI+s6axjAluQ0k1B/fpKRCv76wRzv8hJz9LpxaqUnXDV4E
FFuBAXI7Vt41vzj+a2dHKZGXzbxVH6faINKo8HvKFnSSalcKfcjay7vIpgWoOjiANkZG7ckRbEZC
/vUfMWLom5fmcdOcZeWddl/Hbf6kArn7SCCy8ewUWJcqdbbbAqnyUCQEhWX6aEvKpZ5PngQFBV4w
jgqV344GsHfTwHIazkroh/9Nja/RZfNQwHF2jT3KQX7ZmZCSAyz/q6AbxKi+bVuUjgQgQyi7cvR7
St5W1G69VuWHVeHFLz6CrG5MbdDRarBdRdooTRi0AqQAKPRPUlUSyuJlrM3pNjqej2WOcx5GNLrO
laDUf/VM93qAgn7oRvSRdrqgccFczHHyG4/toYWD14uNn974JWONbHBXYfUJ4BqVVLnuo5H28z0O
CJz9yM0Gx9O3jSson9PmA6aKeT3xBKmV6I8rpuiS5dZws0nAgzqRtSuejd3KPHnqaka0JC+LTsB9
QLAgXj3t57uvOHqYNZUZtPdu2lLy4fw8h8UjunyRzkOSw/SE87RPN3YdGGbvSfIUCJnm+H443jLV
YaBdPM9nXArBguWjsYyinbJdQzQWKSG1/rbEFRN0/Xwp0qSAqQ9AggrtqwV29tYs1vWOFRV1WhZW
unzH3xwc4sH1SRIoTwQVUnridH1lak4gPx3fbA1eSWzrAh3oTjLJS4fsUNBJzRbBUev9UYcMpnnn
Tru9Wr8JkCrZXtRgstC+0TSHNiYTcbPdXJBKVor6fFDZY2jtXp0ZIFbERoO9wJi1p+65/zh1XZqd
q6dDPR9hcSsdLXEGUerZZg9TfOvisDIrZqAXi18ssLwkEpcgAyJylZG4KYXveFo2rb9rHFZt7raB
r0T+5TCXagQaTdJkYZxEOalYah9RfSnEmjhN5bneV49STW2RmC+kbDtqg+UBciiVRizESYIu6pY7
zJU2aFRBj9FrHabsPG7zKABIHZdAMZJSoJSxwWx6tIk6YCvgz4UnifIPhQBc1iksiswTUqJOcblg
M00aOEj1y9xG1hH+xeXvI+Ncytbmtr+oI++w3dFdaEhDs27e62KcMYUWpzkf9BJvM9VSizpajkvg
Pr+Rkl/Muv/mWynmXphS18N8RK1JeXbV8TnrUV2kaYGrRQN5iuLnt+xOKFETLSZYpMFxjh4TGsx6
05rsZ0Xz7MOv2LZ/VOBbGPe4uNWtnbXpOCb4OmzR1F0cbRXI80cJG0q3EZ59kv2NCe7IR5hHIJ28
Ea8Uro1FdBh6Lgic4k05r/fbIm3Jj9ABHibQAE35TyihNGp1MjnA7+gGh33353xrj2aqPpAR9TbH
VkReIztvmRjGfhMq/f3R2zisGze9RqBJuzRkmdriazEg2A1e/vRkeHbNv0CE937KDdGAh5wX3WJH
5IB32kuUCwBHTHNzOeLw8vkmjSyEjx0VidXauASA/8jrX4/ERWe+ZklmRYcgAPOHTHAWO8rXwrzl
56i/s/U7dKTiPnX3q0aFUxnSIDiRROGMQHwEdYW10FgnZLcelp5xeWyAaY3DNALOu10kxWuUGE7y
QD2XaHGmbKrFbVWd9ao21Z4XkrurV1kXmFCl/r4PEuMDAr9I1qI2Ix9Eq0QC6FijQxyhR5ycz0jZ
gXXjOgd1oIr1j+xWHHDkDlaKMe7yAb0XfLHKooIFDUHBFRYfOLd6ZjqNSNWvKWcp4q2jBCpiCcEB
uxCitHOP0PugWbBZt9j4OlLDRMWqY3fC1eniWQmX1DBe/4hi07047Fvtk46yyTEtGGIfFjbaapoX
9X1Z6z4STAqus6aCtKUDfaVjPjgCkXcd+2aysJEIPujhKs5edQgPom/PXXnjkbyOLMDpvqMIEMWJ
H8l0sVsD5JHa8nHYfxBZNeVwlD2wc3yldxJefwnou8Bl1NnKC4xX5+0E7ya/q8PjCjvMlNNn07G/
1btkrc5mzx4VGTk00gTmlwIR3elQz758hw2VraLqilaJEmtt2KbGcGTntK4XOti/R+aAcDix70vk
M6iEJlbyUnkck6UfzIEHwM1bkK/urr1U0fAajXVCxtWKj83Hsqf7Kz70Oyr5S2c2bUiUeTjsnjq1
YrhCB375ZGrCUNqFsk/haATHQpAJjs/X5B8+WF+f5uWoqPc3AKWnBEkjeSX3R65A2DhDR68EGj7C
BYaxiCB8BuTh0gs+piCS7LAYxnLyreZoVb9fOEH5Mw+9RcGi8eDQsCLrFiniLf9TAFH+YEh3FrMp
mi7rEWztaga5+btkFDzH1clqwu90IoxvHSm0fzaJjMAriVUBxzG2Ts38o+Rlz0zgyp0AgflvleIm
NZEA+mtpcjzWhA5N3AUfDzvwdVBcgrnBXO38Dhpx71T0Logg1peVYQWLs5lX6n45CiRX5wqlrD6B
rtrg5d59dEIY5ecXmKSigjshQkMGXNxOuOtc9roNeEbhoPDTmZWu1aD5M4oENp69E8Vy/Rv5XKGA
uuDN9bt0ja5KzLX4pmLOvPlkf2ODRroqubx0+tniafrzGKLlSQXiDGJe8BMvXkA46MHiPgqtWgZl
Us7u3GVX1tPtEV3qaBhEth5NyBW0e8/8lR2W7hITw8rl4oB/3jsQnFRM2hlgRyYDnzl+f8bN1Piw
mRYfc82Q1Y+j9RZ5BlG62tV5FNv9HXxuw16c4Hx7CRmqgGU8eYDS6QWbWZ08WBJXrWFxi7AMfDSV
JHF/v1HV/W5BfmeGYbDGirUcEfgAbERQ8LVgDjOAKHJJ52yJ3QNRqRGZt5Y3FKefZtQT0lc10iGm
NEO0lVFP1PFYcG6HUib5CHh/u3Z7k7Vc9Ke4G5ofoxEuRwdgjOFHrkCc5BdVTHtsRrQfBQBPUTm0
FXXfPqW1HH8pYfrZTSqwQcb26+wTk896kay+8NEKbVN0HQ4he991/NH/w1JYDmZqdkOZHuzRxd64
yxA8of6eSuoHJZpu9ukWbtBUSYU/PHrVAz8p3BtvV1yioC1lWHepO4kAzB7FU/oTqDHkevimTn+/
q41QIsQJ8Z/MfeFkIJVAaktPHLubNdiuoeBJV0efYoH1bZcNGqRnk2dJkTZHbGHaasuHB+odjOrV
1U+Ty4bHkLqnLz1CVGRXn5gLho6Qmdv8rYfLfuHR+9/QIqyB+Z/ng4d7vbAN3r3vdMCi64nyZtoI
4BQAMKZmpyCOpSZWmeNipeA+AQ1LpsvKJ23+mYY/PnNcxgiP1gbS3xU98r3+TBoOJtMh/PNJ3+ut
FyWz73UcMK7Drbh2xnjPO/Rho9W6ZhG9iQNsjEjQytoUAc2xSAgo6tuN+ccwS3cANMMUN8ozyx1j
109SkY4Oh2+oNSvN7sn5dA8GF8TbsyRyMpGDACABcZwZroyNwxJrs9eBMEOtZ5VHN0l56QCu4+LG
M9Ohkfo3oq7Zba44JoLclKTymhVTIYVKoBMFADdYQkT2YLdA7OyEEgG+GbejRR9ahNONP22xa5WP
gFmZaYK2DD6Y3dU41FOf4ApsJfBQNoFq2wbmEiGUOwmZ4Szcq6xG+DSfAlaXdNNBvGxwUFjWdJUK
xp89PkrAoQs0w/aSVZkVPTHKGL3r2r0MUiNa/pZ/DEtAl7ZAjyY4HszaIBaClwknhBZLmztUeEWX
ez+i/rLb+KCCUnOO2NtJdeT6+kcIVInXqBxerIJlfdE9gJFrms8gK5WvkQj4q8wtQi6PJtxQgMNd
erHicNl3D73ElKSqpCXhrtuwTyCYFLJ6TVp7yHQJyWHqCTGWyOqUl0n8O7AxQSnc9A/Q9d9r51Sc
3mmmHJ6R5YfzDyVJHz/md6uFjchiqFRiPC9Sidxjdp/zn79HKocPQ9S1VHt+c98yxC3J7L4IurCX
zvk6DL0dxolWdEmFoG85uLNf52Zfyivuqixqs76SuCAmLWiZgrzvMKvknInvEDuVrpx6dEIQsjZ4
w/afqgmGMQRzWGHKfNC2rzUWeFx3s2erZojpJFLjCrrIBM47WB/HIdefRhKwONJ74V+ZstXLrvI7
2lvlxm+rkB9y14bVn6iVVq/jWGLh6b04bcLKuQSCGc4tTmKwKGFHxQyo+Rm6k2jPwDwbRx42T3zC
3ghbMebHuYWAjS8wnoQGJLVp/1+rJ8HxgJ67biUxGWp3t3QxNqZYq0a0o7K2JOZ0y6raxp3DgyA/
5BLh4eWp9OkyVk7wkWvg3GhISxqU3CCke7YuMCXBrkkZTdRjuZvjDgJJ310DDn4SGnMFNfuu+U+n
g7c/AAFstntRn86P6+WD0pC0A3dotwIhas7FKfmwnOEfO2MvxlpTYLj2dk6rYX3S1ZmAxDlZ5mbS
H67dEQY7nvC1Zbu5l6sBjhZ5/VJBP3ITnBAP0Dik8jjG0MYCHVrwKNSZ113s7ox8VRr2JXzf/own
sl0HYWoXpqX1K+s7sWltCxaadFmYeIBkzxaieBNjXFm+eWM5NHn4xGihHn4pYNFvjpLSQo9/E+h6
gZpxVzzqwgwUNstupU6jn9UxvN/H/3oqyGvwri3DOVXr+vVfmCDIrh4elFEtKj2CAkghIdet0IRx
/Q8nw6ZFAkSWyaKo9PUcvA9JYSlx8JX0RoDnQ0C4V0LEaH59NrCa3OqmmFmorHioy2mzvuYyK0lw
MUQC99NMAbEd97Y19x1YjlDgX2oDD6MNtgzSiOULUeI8PpVTJWJYT2cvG2hEZOAugmMBnBro+pm6
jOA1HTpQKtsVZsN+BSIhzXRQWZLTbX70EJtLHsOEtcX46fQzNhjxrdk8YJY6itAHMUW/czUPqnpi
lxOxnMjvHBEeCZPV+Rq66qsVj7ZNBFQO+ROCscFI70l2POOSvORbydgj+Ml3xXV7WCbba40yW6LV
fUeCSuLak74F146zFKAvf7K9mkY2MtN2UA2bdcaII/mSbup15RA1ZWmhy+NkBvHECiJjuouc+qge
C5mEqsCX+QfO1DlTlzmOKsKeLhG10Uh/tJHaVeN7zI4Ni9DBBUpJswrJ1N7zNTFQvUrBOPNyZ4Xm
Rb4kjvnHk2KEcQ6hDQJ3Cq04qBAJVeWrAEhrBCH+lxNAnxR3HGx95BXac5Nu9LusP4pz3Eiu56yZ
BmU7VCrTxl3nO0g+kIlEYHMzvL+juxBGAQOdZw7ooTp/gCRzNlt8Z4xJilNpsBZaoVEOFQ/Ly4/j
RnpKd6lQMAJYgmOO5FPK/8jLHVSmmSkY9Q/ivo0jEGnno3NAnAPdHfRiyRnU7nCGOpwZqnvda9d7
WIV/21hFMS39C9DeQ60eS02AfS1mMOoFJRXTgyrJDerFHSRV85gev5HOvQ8+OUVjuuDMzHYkOB+W
DgVlzOWt8o4ZbNNM3qzgSN/cDrIyI65XZHthGsw3Dol7f8DGPRpQ2fbtfOsCO1QU6lGWCR49i73s
2ByypNPGgkekNGoczc0hA9/dYFvAF5NOweqUcrd0gw2hfr1IXWmx1IAjZpvIUCcLiwAaCoBn8Zyu
kPweaCoWI2JjKy7r9gTeRugz6cFkkWMKxdLHfKHkHvR2Ah3mCjBN15Djc6JW5IVci4Ikxz2S8aK0
5nYtrapF8g+q60J6C9Uz6+/iYS04yA32i9mfepiALkk4UFJ3h1bQim422k8Z8Qw/mWMp2RCAP+tO
Vpeq0O4FeDgxTeh1v6dHCNxGI6JBIelQmAPUpLxfy91gQCh4tmJ8Zw8hrjXu1yBHAtRZ6Vvda6Mn
ayAFrpxx+HkYqkOd56m8OcX4aPw13G4zzEkSgKF1vNRYZpFBfo3gh+V5Jk1kx7U8VaP6bAg1744S
4k0g/z5SoIDDcFuSwlI9Vc9BSCX3Xx0O7XV5AkeJSY0PgMxodmNkrqawhoanRRa/hCDGaUDh8eGz
vcnpQwTbvT7AoqdSSPYlFk0e3QsmTI6hEsvzCksnFuZth+GWaV93mx+PqtT8JYCWWAodU8HnxnOX
yJE5FfViv+RBtVyYIZ3rnN55TTx2KuuP65USHkmdDCHSr18mysuWBWv8Qi7TEYE8Mik8fSD/g0+q
2MEeLyWNs7k6p4MOtAdBNa96QnB+YNqqbFAwweW5jyMCK80Q+gx4nzoon39b3bD4MUjT8scIpDL0
eDegbx2A+xnIAlrWdPnod/1fNWJJUXleveaYaK8BSIbHwU6mpgtE46vTNoS4uR9wCbUPIOAFwvwk
JpmYEkjp/4gzqFHnRCpAsUOQRsGbIPbSnQYE/nXHjZy9ArRbDX/8IlRa1b3XUDHlNBCpVfi456+N
Sov3DL95F/Z82VfpEEE8x3Ss1MXF1t2QFhjB4SwBHLatJtw0vg3aFesKkOqsq9E1Ok8sRdSO+p5q
AOzl5ZaWgKNO5qu5OwKLDmBYGydZ8HTuzyxbiGrsJdVnOfVVHQLchg049FQHHzw3Zs6F7QKQQ8D2
GlY2ULfgD2aHkTgeuERj53qvNC5v2MotmgMsL8jSEVKJlyEXN4oBtyfGJ/3qPGFr+hL5vW9caP9J
R/ED2MdMGbUxmgQKWY0lkRPzBNwEfJd/5P4eisuFmwE/8a6N4jA1LVGZERiAyEiAmjwBpHDy9kG2
kLBYEKnmsL+bIHqBmmNkX+NSuz225IIIjTE2bqXkQTTtffPqbM8s9IeIxcK5Tl0d2F2gJrLdpmgK
Jwtf+3l8LSCSD97Om99yey3HWQyYLzhg1R1ZZ8FtKgsntYiA0fb9XwM1H2iHegFyQ3/zFooEtc7j
HId2sctSRgrB/toJNn42k75mAAcGPR5Fi2vlTgah/vwSrkyfXsDNm2dBRnY2lfTcNs4LhiyuXFWH
XbPJ+sTmE/F+OoPtBfygCKB23U7fCXw9T0blNFxaBtZTh489Qqg5CJzHXHnEluZGRhd5pZSx1jqR
N3dYN/yjMIWxSQDeS8i9YLw0r0mVgHv1KT5eeNkjbdx+Pph9uXyRKxUA+NBeKguRfHZRre37YNx+
HtOsud3S7G+j+IA0IFGjA13KKlMltC3D8J2h4YMrSEl0BaAWmPCyYWw9d6RhZ3c2yS9t5OsHg7BB
erJngWPtRHbPopwdqKQO0gNZGuiQYyUbGu9eVenn3pi/dNZqCmtrp9ugXd2w0kBDGrEVcMbOD133
16WiidUIDmbF639n+RrYZ1Gqj0f7aTGd6HOd7fcceIPWmwBl86C0v4pEjl5ai1YdIMNQKNDrQTPu
a2WiweH2doDXO+JePtfrIl9P/NGLi1UbhvCVfn2ABCik50XyrYWNd+GB/nd0J/i82Dfmq8PEYKla
XFY32o50mP7f1LNHiIH4un4a8Y6/OJG5V5pMuh6DDPxgF1d3aTc6AMKuxotk63OaZuqpoD+L8af9
WvMACOCsSJRj7kZoMOxPSLb+3eVzZaRmUn/8otJkPtpSRs487ndPN1EaqZA+pIFNIghJXKo9IpUR
54PPoN0zMjBfaj9z5TFIDvmidLmDUnGdGg8s9OER8m1Ggek9RYJrXTZyF4g66bU7ZPopmVgTTaCG
E7wFy5COPTooI0iaQmvAri27+LhQN696kTA9pr8wPgDeOSeQWeL2bfS7HbcyKy+dETKx2oO4I7RO
wJLRNolkCdsQq2Ri8p7uVfEmPTy774o+KS1dn/pH/kG1l6bFLQDuZYBFDxpNkEyUfOLLnuvxjwpr
/rA/z/i2zkSGwR2RMAmyGSviiKsZVipkiO19NQLjF8wPiayQ+erd6bhpBFT4T89ieFyjgsQ7ut2i
RyBFCmg6lO1DYlGul3enubNkR6jB5OifUgkNp/+BIjpsFL7G2tAqIQvNsVTdlfJGPZ5/LieENshm
w4J1reh+sDQuU+VR5sdEWsd7vM3fTHar+Iq5APqkh0W0TnP/DhljTXzZ66LMCDcg30oQJDNl4xun
r3ycqSz0mMUo/QLCDWFCL1vKZB6kczxlmKp9j3aU2pb7tfkHljMXyi3v+5c5WBQZA7bTXZPjK3Y=
`protect end_protected

