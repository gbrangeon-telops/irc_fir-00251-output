

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VHfaMJ2jDU0R2eAkOntfC5B4/6MobpZ0NSnc7trviKzQU5KHakm896MNUQ/U/XUDUOQl1Ix9hEug
uFcdFGHOlA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jZ28dq+cqatvP/oWT0j+kbhevax+rcvgcOVET6FHORIxsClPAe5EiSXk6mDgtoieHOJgnr3iO4zI
pViSw9QXhHwC7nkjQzCL5GNnIAYREubhi50JKwxrsTofbyKzT/U5b+jDP0girnK+nPIjwrQv3vvD
PHropUlOeQU1eg5rEJo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wyTaR+5BBK3PMm+GuCvq0Bco7y5f/oiFqNMyoEJ+yA7qA21Rc24sV0Xv3v9W4doHSIdeeP0oUNh7
9I5Dbu7bsdY24p4a6rVQlpW5VOJjg7abnoTszev3jaBtBOpAM+FQDIkOj6hl9ZK+eUTOGH08ap1P
3rtu9S06fVXB15p5GUL4qJ+pbX9as7bXZJVw8JMDVFn1WsdJ/zMn5PNvL5qC5jZb/F7Sf9m7DkwY
x8I3vpZz7RsD6/RmMhT4lv1FkcH4MpJegB1J0hL5KoGG72FOKCqONCLsZdmnqz5BmJzgYmphlYZC
jJckdSX4yOLEg+jbosSObzMclIjrm9gORAOhKg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qekQcsRlt2+SE3/eW9XQwKmx/wWWvcG3c3jSLvuGiy4GIetXM6PaXqKAuGTMI8b+mux4A6dEdodI
mIX5ojnf5ZA1jyISA9q0jKtn/LDbiV/JtKzm0pK23fPqh9/IUaTz+oirXN82WQzZFKQ5TKpwrFn6
ZmImSJcOKVgUcM/iG2U=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tlEZl/v6lEdJp5aVMLYyANJmLh8DNrpNnDhyEkIUHbeTfiozIDqQ3eefGpJHd1yUjxDr+M7d69UI
c7u5loKJo9CP6qAEjMhB9NE50dWkO/cRVvdlBQSlpGD8Asrd28oTNAHTTge+6t1TRCmYfvMKOt+b
zBqmGPTyIDG3LI8DiLXNfUjWjl16n5IRikeD/e8FsFJjAF/a0Kjal/N8CzCmRiQPdsZhdMiruSdi
vpIRkNPRNpCK4J6asTfuTemt2JkEkG10IvEYhZ/qTCco9PECc5G9y0loOf9owc6R54o3iALi9D4Q
T0iTW1tROVF1jLbRTIe753z7r02QD4PyC+02yQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24176)
`protect data_block
XSN3mFPLRzmR3rQ03lBeW6aFXtlPCnuKtxKePLAmpvtNFlQamWepSCHa0QKpIosYLVqlE9VpoUk+
lCa3fu+0M6FvXRj4kx4mhUnu0/3BJqEFA4ikkVs9d2bFMctdu4ARExFdZha2vHzmd9GQfmWToFJU
1kY130mATn9GTSMWqLRTW1ES0TjjbX1YGuHhIjQOiigUnsxev3CEaqLViE4u7sZXAcM3lpyFP3bA
VcDOMYpaF2NU6c0DmVW9CBdJup7dCBWmSEgPdT9gzlYpiKueLecxYVuKh/cc3Yyt2nnEge1aDfCl
XX1pDn0EpYc1ZCCI7lOTBu7d4SuxmHrbck2Hcrjp702+fDBLRopBdPB/Jp3dAOYoJjTq1OMekciu
u5VGxY0aJucCnIvAL+RWbJY4exe7ubCQF7qsCsi8jh1C8NbWP3EEGcJYGigL8anBc9EtecjaO+2E
ZJWfBDly7XLoprzVwZhHyYe3k6j7On4lBM8+xX6/T6ejKdkuL9AcS9Wl2sKskDULQzO3mX1qNKrW
iQDlQlIQpBcP2tNmUU/ynSFbVOnt2+KrWNDHgmx1fYHoYPLaLzF43jVI5HTKJ0E4QwVC6l2ssSMf
IRVROZ/i7QGV88iuzNub3eXKp7xLcrev53rwveiJnDEM0CBQ+c90DCMFgbAOXcjKMexJCiDr7ziI
+nkd+FRQhVqlxAO1b8kjBi/Ak73UlZs/lsZdiXCDFeTQBhCaIXyOTchBtmalyOP7CAvj+nI8NSTp
BJfr9cftthZybmyZz2GiZBQOiAVZtg/4Y4C6WFZzHYuxc8p+gXDalOdsGqOKxgPk7W9y/qc43HUJ
NWVnFBz9sjNX0e2YYdb/vNESK+Nd7mqgqIJu8EYZqhqZIY8M29Lux1JAGlsICjQmiWFczrmgTu0x
EPfCe+HRhNuexBMEsG/H/6YvKF+67fk6h2RmKrO/5DqZ0S3ls0vthim+8bwH9Jic6cJvp6XuqITl
IJ7PA0CaA9gUzsoFbh6c9hx/ki7VvbZdgHyJCoZDZpU+DYABYgkH7EEzhZ9DxjHUPQB55kHh50VQ
NsuQChcQcpGl5gJHGEDto1SCIYmsy+wR8BnHXPRQiup8a3n4nLxyov2xWtvU3+ozwkF6wNk09yfV
Dd2716ryc+179npdm2MlkRsT0Ncd28SHkQ/jZPOiVkY85+z5nOfijztz+QWp6J95oPUdn61J0/Wj
4FrLpftgeiRRt4vrsJ+5PKmctzEIsvcRfs/u29UwsHKJiDBpZhNrESiWYib43TPFdIrIDPWtaDsi
ZF1Sldyp9XMwxMfgokvKfY3OLQ/QuC1l3lU/9rzDKNbZgPh6f3p8PHNPlswDL98e2CV53BC2l/ni
Rhm+/DEI/VeIkAKGHps3QNbYudUViOeRRdwMgIgywWJlC++UmpB13xDZKtZw+LvSqftVbp9znn3Q
D/5BvTnhnETdPFsPCunl91sJ2I9nD1XLnptzbhzzHlxJn+/p+Z4FbJ0xjR8698mz/tJxe7bTApda
m3OgiikBMy7e41o6902qN9/JSSAeIonO6dkgGD8Sw1ALcTSM8TjOby5+RTnemZG8SXl7uNG5GIEC
ZnI2Ln2YrGd1V7TY/HH0WCh67DpX1XlTSWOS141KGqWkEYDGuIeCPT5IKlagUmwnOEVi56fdiuSZ
8VsOZmeTl6XCbvS/BySFXRsecQ2FtEaVWk3uSTVxf2tDWebUKOn0jFOwV2lpG2rcXOTVjFXc7YqB
3OQ/jeDF6VQ55NW3Fg8L1hrsXp7PQteVry1GNa40K85pcbO0PeTeqmrwCeCgK8j9XBn4S1JmtoOE
Z1GUOXOe6739O+LA9mim/UP51HuvGFY+YGYxfTSqic23/OaYj7pniZyH/RL/ZD5ddS3Cx1UKvdNr
GUejf954UUzAMmkLpTkoYm/dB+h9eHgAy1C9SEQ/1WD7xko1WCDdUDGoJzGzG5dH1nBW+zynGMJ7
3I8FCJ3ys7iItFSSaFrGuCtvTTymMrMzqDOEsF0f5mO+pL6ExvOW+6zbK/ljOl9/WmUHCmj+cwM+
8XqKTpdY0attvI0XPDvejdziNiJaQ4QNC730ofP6gOLS3UE5Bw7a4DRJM1Qpe0lk3JPZOJ26e/ML
eOSBN6pR4ZFRaPBu7y0zLRLl3kumzW0Hflw8QxVku2voE1i9teEko8vSXBOAKhxEMiKNxFp266ci
FHzE8+wGsEHFWw7Fc/hQBNzasUI7K+dm/Fm313CmoiOlkklektnHkRPXIKtoOz/lHquXvw0idvRE
PW00pUkfO45H0GuvFe0nq327psqWCy6nccg411k0KGwolDwMH18Pb+/3VX9nxGugNTqRrZ090V4L
7sV7B5sdHU2wyl7UGqx6Lp57cPWS7yS7W3BNyzfSKcn+I8V74uvwNY6YlrnDshQBJAYhEcMIu5Gu
yqe4j2iRRmxEd5KLyU5LejstOMCzD7ruXEh/eJJFLT+pUad13SH8s4mBja5uB5/rrAdw1LiIrMnI
IAhvzsSSqkUkBe3Z+wOITJVBMePps98BI2a4COKDPEAATxvZaFZ1JaljgJU9dDnJjbYcHcuKjXVG
4P0VWgMOEXE4WsDLoTQdRo3eudJv2XiY/ZTXss10vcR98fvAL75BAJahRMSxGgefFIR63f3fbDPz
dI3hvpQ3KK3azSxU9Uu1HBBe932WKVpjkiHCA7Ars//g4XbBEpMuW8smWVhecsSbMnKjeOR8TJOr
h/vyFKeayOpZBMsc6EDNaYwCj9p7rsyC+xUOxf6yGPvsZGv09AR3DVuXxQag/1gvL3G+OAW9diTJ
5Fh0NfGZbbmA7gbUMROzqn0u51/1QNFD7hZvcOgZl1NgDQGNWcK8Dt/A35K/fEY4U2rYIL9npTGa
v9wASyEZOET4ljDXb2kqLdYyahDjuXFFueEoHupk7OhPabGs+abaJC+hBXa6rOZWJO8IX9hKhPRq
xNOJRt5N09KCd2VLFHv4jOyLAfesfkbVSq+MBL7jh3mX5iAxqiVmlyaalE4TwbjA2g9AnbrU5itJ
PLxNqQsw93vtA3fsSxXZNOJiWnv3n64TnOxCwgnnlN86AWiz3fUMFu3lFeZi3wGP5qtNt8zH+Raz
9i3feO6m0Z2drCBWkH4tvh0LFY95ngyYXFt5zpR7syV6zf+Lx4gjLULK5rLwQ62rg+/vNjUA9gRG
+AR3PsGZy0qOK2Lt+u4COgZeQsIEVplnoBBdS2W6ussWYFHeJ6eqkcCv+iHbzptY3YfabQZA8Wsl
bROxNDPK2DU8bC6bh2LFlizqnjHu3mi1mBcI4XCKIesrunSmS31vw3tl0464kZmjDy7fuARFXR78
Qr9llkcRvjh/R4nFtJwHbVWbz0uY7Pil5TmgWgh5fWahUymgYkqMe5+IV+W25emHFtRAF4Wt6/ig
kgWLs4OtooHOhZCFqBgHIi/2cek0lyCLfkhKpJhaj9uKm0SIuyhMBylMk9u7UR+ONW0sltGvLwJS
DCzQMMAFdRSx6Z4IjEtiewELLGLn8/Wrs5buhFR5NIueuT43UDKbslWJG3NAdSyDZRW58BX3n6y+
MiuW+VVux6/fe99pIdZBFu0v5QO607VnIbD5QisIgR5kFtsDO374JqGHDV9audhbsVc6bOIY7Qg7
v7iVr5icAkWIvbhvnA+wM+KEysTvvpwobRutVdgyGk2kuEWryoSWceZNyhZfMTrzCZaYO4UOGnrm
gvs9OdYgEij5/m9lsptnTw/hq/xzabh6Sc0WXyJARYuiGxWLMk2vI536mRDFZgxWFQVP6c9Tgs6W
viDqfZFE/ZGhGvCENgLb26ITRgZisoGUQtg9l4aPATTl0ZtNqDUcf5qnRXdZamswWSc1EKRK2/Sh
hUGOOnzbMGIBPttqIV4xluUftbziR6SkGQejcj5jACfNrmdqfsWYFs+Z1ztxlfNViuSg3hEdEtqL
PuvjgbMaQ4lZL13IO8DHFh5+Oz3hZQVHrr3G3HmUYOOO7dMR4nDp5lWOpMxvG+yks8NyzvrjguYb
z7JD0d7GpSo9EdkXtwGs+gtAtfK7gbIscEQOuCNmXl5jKMvCbF9XaoIwyOuvDn1ugL/KshzPdEwE
C+KTwSgdmsgSehXOPMsK1nuSCBwNgy+L/KDJF+Fiin214bZfNbJX4Oa/sicsY35oWfFT0xskNJl1
bJdLskn+kbXuneZLZoJcrqJrwcryoJhnki/IJpXcTuaTiCDidjPVy0sFDMaIx/L8M9uI7+JmLJwB
ECXfnCaw6xPE3yJqjAkwTgOzFGo5IH0I7uhdj31NfkDTB1y9Ls0gN1oYFFXHkAy/iSXfZVIv0fQO
PyKs30GAOco34mSWzQhC8YSsSAYmksTL1LudFnjsh042G3E8u4Yqw3oKNXW2kU8kH8u3RnAc4FZU
7qQ9JoY0wyJqm4c5oN5frNLSY7ASgZNZkXCv85fUsq1oxz+QhQQQf+j/j5OEgRLBrS6Ydgnb+ora
/qa1Zu7930hSUrtM9UQGyhCfspyY+c2z3guo4SLoXsQE+aag1f+4ZKB61Ayu5Mg34N61KbSl/6Rs
l5/99LJIH5xxiIya58CkeOBqhQLaGg5D8OUj8POBLUaUpZg1APPr4OzrQ9kkXjQwAJv2Bt6RXbEM
bDI184nQgpdiwdJmDN4qzwnybPttfoks/75tGc5Bwj8meaLoeQ+pcjLwur8wt7W95b/NzODQRcLM
oUq6JO0UZEMw2h4DGO6cTPcZWqHxYWFIWAyMNEtyXS2HAZKISKKx9wZDPi13Urauw6P4YrZwcsX1
Vd6HgP0IxwSAU/fqxLW0vU6KralAHlBUy96DtaHyoM6E3ihRawMTURspIa+ShsjkOpL/U6Mm0VZK
hFVCL7p8RSctWN/ieBvjlAh+XssuItafv5x4+sZT5LNxB1YS02i2TUa+JKIoE+Z1oHiQwH1CEQsz
c6CVz7ALzKbsL5wuLDsypftfmcbUtSVazfT+K32K0gEPuE9kn6f15jfN6zKdeLoyFqZAPBisaWV5
u0CKuPgk+6/QhrNB1UBoOSTiW/sUeu48TBQpvG3PICykUyRRzems/jdXwVI2MkWwsabiA6PEDFPS
SvxpJLc8ZpEL9+tvwrH6SXuBvufQ6wjaQcIF72MMxh4gryr7S8vbVhfkj1TE963/tgvgq5yBI1Q7
RhXPBqyFq0S+FyWEosi036B17+OVnWaXQN1Ef/OzmRf2M1oNjpnIRoUkWB5lIFNa5eGGyh1c90VD
XrP73gUc7k8GPFT8EyFigefGs0N+6lgw7EsFW5mrsfR7ENct0XpEAK0QgYxsrczC/BASQXmiC5Iv
fCIkX33v830JDFkyUnyOfXKBA2k/f7/fHJrX7lzIHZv2CibDcQ52fhBNnvztSD1KCluSFxD7dnxW
hPVp8visS0QNAGHswwdC9euiE2AqHHHNzDH/FwmWl8ODo/YpySn9HhzGuLcI0lb6uz3H8x/rBI4Y
RUWoIVrvMEvVNFo0P/Er+9JKAOJzYkXc/YQIuTG7mDqe06RJvws/ExNYBUqMKuIvyBLVNbJw7RlM
075VwpUjOUw3SbKjOxi7lGVRoSvD2fiAbpVWN1/EqFnzFKMIXVzSHwxkrJjBPw0MlsZ24muiPRT6
tih4IQi/CjNeXgHmD3Yaf/H+2Tx8X1aiXZ24dTSCMKl88aT1lqRul9Kmg/oolf2LcqRj//yUUMtG
YOvhY6LHtZFh6iUO7UvZn+Wep8dnNaU1e5/Xbe/qzbB4Oy1o+MGWkzEEgV/ZmwbWJc0nW5eFJiXY
rECx+lcyNdil0FYz/AUjFif85TmvZijZEnKtOjG/zXO4NibnOqhlHJJ86IQkIpXwiZfgcyluAqu/
rN16+CzHP8tzAE5W2loTPcrub2LJFxBULK2oFLdVzDu3o+vGRf8N9dSfxn3dep/BURkmci+OIW+c
tEH6El5iwBj/gEoVA5IqzBuEAXY0XP0AhxPWrvMocbR2/J2eIxh6zvdbhZZtusrTTU0bscbroKmp
nZF2zf8vS2oHZWoVfu/N9SXk4zWMGlMjw2dpB88dazLWlEPjKGMgNMhM2y2d8x3xVShThDxKxS/+
v6M7+sg+tHHQDOOL8xtnsxh8ryPdoujJgn8OvcSFxshc077vcmHwD7g+SpPESpbPEA96XCgwJLa1
kc0xg5XHQsfzSNBFdSH4S6rqAuTtUY5Xyc/h6GPnE7AlpgTHjD27dV3tpyoF/TESnhnZpt+x6/Ck
BDZbbXX4DGW/qAqMW9sqq+TdTXuJcQSHTxEv9/MZSrzReFT/bKtQii4e2kLsXGENdkw8dYkaXxdP
dlh3GOnuf4vX42NT1hKOupTs0jU1Ht46JOyjcYGkSViz7BXl+JHiM7E7spwwbUMdbAfN0MgL78yg
m22X4U1PO0Av4+Nbovqw0FgZM16VM+FLi6l4znz+o6yAnEbzyFydsQjBQNTBKbZ0MDapJ52kGjRc
Tc21QBCXE2oCXBDd9nu/KO4f/rcREgk63pVkZYuYhU0fHsBrngCWITYcxNM/Kr7BdvOXvb7Q1ukg
MpmJZN7D2spIeevANgYyX3HgXjcIHgFjRtic5gUl4AXeCdbHNvOsmXW/boyb0qq4J4Rpu1/vvpdh
jgc723x8gdvKjeo0YrGa2SFHw4J/PnloqnCW+9Tw7mf1EKXSEF0SkVy+AlS7pE/ZAXW8Ozjgwoiv
+5rhfd7kGW3YwWhN/cwY+GxGXoRgCxTMdsuXn1Setcd0Ezly7X6aAKQ7OPsupGYpF+HR2lwtToWT
1SVqjoJ24jyDfmA4c8sa45ExMC/xwmdrYSJ9TgChuZfXZtXiHy5qrBjePXX6hulRRR5O9nf2QTcl
o87J3/+FXS+HPmx+B5NLOBUAEjGH2xx4asYn783twp3tKzvCkGfuqgP88YT+IOVlCZzHFYGxe+qT
zq0A6F+fcLBAumS/aRZOs4fqkRpc4HICEBWdYvRXx9WmmRsvfNpr5QsWSCLNIV4IUPoXZ8jYrmlt
1oTIcFjUGuFRsWsrCVEPl0PORa+AOBnnz2H8kHrUklhaq3V95+JYLMVxtlbWE/w9Is719+1V37FQ
nfL5CxaJnn9Vc5C18KpclfU8azb5VjwoXUP8bXxqne6jnKMiAt4EEg/iTNb2t5rdvWo/VWixlkDl
ijh95Y9gY/X622wsjy7+FbeDD5Bq+mrZZx+YsJ3dzT2vSTaFG9v5jXQRExyYRUY9TI6jLd2pklXw
4cD4Ky2SXPGNPkqXB5ZdLQfD9QWGpc3mPpuJ/zTiaHoEcD9zSLu2rpXQzT9xR2pfVjz3E9Q7QMkZ
G5oYEG6MIbWLfG77Yc3HiwNml9sHJxc8yIBgc86RLv7SlZ8Td63EIktdGy5xATOenM3oC2I5DwB3
eEU4ZzfL25ULR6pwt+jqsRIqxuv9LV4flI7zVksEf2jKbWhBdjkiepQQBcshiGem7IR+3JFvcZOI
sPkXXIkypXcpyd86yI9UklcjhrR0dnim+8TtZ4uQYrd0bK7xB3xXe0BFicN7t6lcIvNRw1RQcR/e
Q2q95ZhJBQPyJjW6/mN8TtkpbIUzr8o1J+OmZ4YJ/olksr/YATy7//S9zJUPM9Gm8F8GQBLF3rNl
6Y+Ct9BQIotFA948RBKhlYjxS/i/ZGG4s7cIa234vjf6F4fPQnWM6BluRLTdD9l2vMdva1Y3kPYk
wwmf20MK/tguoSnDAXHUca+gPW/zkIsp5qkYOEnXLXI2rs3w0pQ2wK7gHFy9K5iDYYeyBik/UdXC
gL/PEl4N3dULLipX/WAwVxYmMzgvvQj6MqrP7VBrIsfLk7HZJacqgIvjL3S2QgT5F/I3+rzw/bbC
+Rq8duueJp2v/UinVpHhAq8pAmoUvkKizGfTSWJK85maLmM7YHN9ML5QfI8R7n33owgDgfnNTWgV
HHUXFu1xRU+JZAVgfmdQWqxbGzIU11mUhDR4R+1pF8413xE3jOKoxIvG5IQCy4c/0H97oBkYUnUr
bpcRBpFMbltNkTTPbCZgi9iIvn7PNJ/HHt7pwFhJ54amet7r8ilMtKA6GF+75gMRklJ6+xsafv8K
wF18xn1r2pZq2Gg8GgptwwpZZz3mkEZrU8axVM/jUiQH02LblvpMWL/EMxjl4dOZA+S9IKeNp3kv
d2nPfd+tMPxC8afwDcz37EtTD2/AH/BahFmbG1A9ErV7FylaLvPgDFl9pmg+BXYG7ASxOC/wMRuO
OZTVbx6WWA3eArD0DHAs+yuGw9eIAI3WFc1BkgsN0gWUgvlm3fug4PDtvKE0AWe3Ngtu+8QhpsOM
1jjpmbkBt5pMXOOvc/sULLQBy5FuyFqMLLVHyfbLlOX712dg25GKKgXOu1/DGkVogbIeUOUPIgT2
X1rPS+TzosgUDT68EhJTGnLnG3zsx3/t81hCZ7MlE1CRBoH4y5uipctkzCrUWgMV4qn1Jh51reGC
GToFeg90TrYqz7JCtIuHQuC9uRv7lYFDMoj4yY+NOGucMkTmNVEjJpXbOQW1oeYSVCkwpaf/kPlj
ICxrkyYaLDllSecWdZzfnha1hvAiQd1DpjQWFSWSsSkl/pMNvYo/XQqkEgP+GwclPJnPOAfOqeL1
a0QEt2TF+xlQT7F5hta2kgDb71g5u1LUOJGRHJFZThf7YKds9P8N4h5YqsC5EM578pbu0dzeImPp
aNDhpZ3Gf9kfOnCLGsRHbht514mJaauilpJbvbg0mer2icjvRqQd5vbSMdVl67SQjRSLcO3S0uiN
RoLFWF7i1tDbqnQdSE2lWgy+JJZkmgeEspHrcMJoSxKGi8C0BjDqsPmn+VcqKsaNR3d7YC+3qUgT
tKF3PDtGWub5x1k8frH+UfUSwqd1VdBQwCm3DXj55MgUMGQMhl9gdsKISAiKFpCrdCh0VSdxmCuT
UhzscbO9mqUfj3g5AOohLuU4XEJALzLMJ9zH2hvZ8YcFupITfVUAAB6gtv7q0uSSnRpxXcMopZxH
F7t/4jJpHPHh2aWE89vem63qWVUIPGnlrjGoQMvORvoVlvC8FiC/tqafJXN7j5Xb8uFG23UqUhom
VSRahfSSxDJZX0QRX92jseXRf5i2avIrRW+Zi7UdJF4Cp+BRP2NqOL41z0iq1pS2y/4XbAsMWCGt
HMBewvFefcxzH8Z1Unv6gQTHVIXsXa+HyQmSGiigKmTGQNSBShRGEdDVRP2kUaFwwinBLhPD4Dp6
sa4RDMlLem8A4fAe7WZgzM/5mF6sSwyQITuQJoD/VYjfBsrMrp3u6cqIerVppqzc7TPqjAGHvJMO
Z3/5rEl3Yzj37CHLRJCVcruxwBUVKhBrjlD5aRa0EpZgIegBFwA3xhktM1awwP7C/HDseqAbKBaR
9SmZ6G/WYHoS08WhGkqU9V8azUSrBhqKoJAxEuyXTglFwPXsNj3steFOI0McDkNQD1qHrAxYybpP
PDbHzoS8f12eA7V9FQV5PmSxzeuWFSbSvT2qFAjvQ9B3vaYxvxCnSHeUTMILdsZrmujBA9+yqaBi
LwAq7lTn2DDLyAIdpApi3Zu5rQ/RvsDcqy9ZZRAsxWs9QxAl+rgIFuj9H8tLEE0tfUYSI7WJxY3f
G0xGmZ1qwBZlKiE5vr1By2vccX6CZJ65ATl2DTXma75qJ5YAZmO1gm+wwLqJo9NiDPvMDYDxVVhw
n5HRDnC8zXq6xtdK8L6GiEfY7AKW6NnVA/dq73g2uigR4eNHupWxt3uxYS6fZ0JZyG00ck51SuOx
4KiHtaBJNI9weaU9euMw8+Yuc0+j31lSQIvW4T+FCN8Mp+BknFAM03ctAT3vKIQUyG2HwQlLov4i
uPs+j7xbZxNs4ByriDi3OdehHOrsflMrUYbn4wlkwL4SrasFpNQbOtDkTNJJNZtqf6geAkk4pj6V
5LupX+BNgFRw8fPYc4699J0LXMWci9Mf+ay3HxcTunZ/t0ybMs4eChZFGg9/MsLIO+2APhD/DyDi
cdkW2MrBnUlDXiaPLI9GWKI0y4Dpg2I7KhRq55o/sZ+aNXvPPSX/p5+mTZ0kcf7LkQL+V2oc9wXi
pmHVKeDPTDKFNU2S1yn661euMqy+vBrV6sag2gZlqBK2hE+ZOQXhBfMUTBvr8PqNwIA5lvhFk9yz
Xu7a5kAv606GzU4eRtWKk5achvk0mOW+ubZ0SpocpcvwgmAOKTkaK5QsZ7peGQZufgVd4mBg5SAY
u4Q3KTuerlW4O68A427ExRu75sARjLpZKDFFHvwcFJusR2VZcdP5h9ELtgSa/yx+pArNfdLDtFTO
lmzcapKWcMAIcn0EVJWmgYM9LVn5udXAKhSZLUOcsNdGoj2jCLtBDTwG+IP0JmIxVUfKE/6YOd/N
0LUzosZbj3cfKvgezfynos/xNSA4aR3mMSQSbXpcAopD6YnzyN0N+z/hwWKoqizARaCGuuCPDERA
Nu1rmxVr2w+lx2RDR9acSwVSr5LPh3jVrCOpy1uHV9ns9ZvYcDMOQbXWdIgYEqRQj+yTBYdnKrdP
6lRwXRsZwwqu5XXGkerVg8uzMBK0NDe1rZ/ipfuVSipnqxJtUNFj/6RvA3Bz+Be3Ex7mjE/3PgR9
BuQXuxAved7DD/Tyv+Exz57UTaeyy3eu4hP3NHsmUrLEqlecClO8ZFCvcMQoxyjJKfZdtlzER9OP
tT297E+s+fPQcmjBFkYAF0iPnZyr2gRcHGOQ4ykxODq2Br4UnothvXXwtt8f38DdWCJ135ME21wJ
8bLQFZQz/Dhozj/r6WKN7LXfWPcLBUfRhvOcyXIvUa9doBrBf8nyA0MWdUcsQW4Y6AjNQjs0ikHh
SFa23NlCg5xrEVcqU5J6H358CA3dKveHW9XvN8Mq0CC6BJK/tka9fwmxLh/G9n5eoF3K7qDhd0f1
kLck0wH4qthS/w8vBNMR9Tnx133MabGMdL4IFd12pa6XQ9YGtYZs7hHsneDiCGHh6MiQNzSgCRW8
p1xOmGpfwFMEuR7rcZJMuG4pM3QssiACFrTglqqbnkGO+XhxPQumv9cKxGx7dI86ZtM0fnzsN0wz
P4+Jw2U6c7vPKX4WBr43dLCuVbR36QisVQByoIoXXiG/PZKcnQXPflt/99St+Z4PdZYzVLEYwubh
3nVuRnmOm/9OuvxTczWhGPBj30tpjpKd6GNoLcuqImWVGJJGdu5DpDdrl7i+Uy5rS3Qz2b8+OFDS
Qq6dkb8ViGbdovRhHsgK+xouwHiCVi+/MK5MzzoQnc9er/rrW77CIHqVZkzAEF4xZqbP78wvmtb6
SJlBKWVqdhN6sFa8Vc+Ta4IiCYcHanFr1lYV5m0s9rQ5l4tphmgyDK5aUZZ5yECC8PVeTgoCQN6v
LOAjDKkwcs/NA01pmria8YB0uGvUOeFJXKHM9GDsuW6MOvGDQmYQGyOX5+AmHA0DRk1jxLji6k3q
Pf+Ha8QGUxOXL1T4tQ0WZwHXIewkP4bBGz2DTXpv5l0KktIEvJo0ahVYulSTTsD0L1KF3Y/Hp1qA
acgyaPMqsr41CM2RlIduKriSShRQ0k9nlnzAiRUFFsfkjQUIfqhbpNHbENumQ8gCHGdoKIgu5tMx
EqbGHDwwQg8xEE6sV2b1K3NUNNnJ39oeyYExSBpwOQR8UX4SNf93aNRrLCxZ+yon2PjycCUkntFe
evrAfkFb/91OC1OakENLWbCdI5fyOo1xrkzS26gzouw1RIlEUxxEKAPPGYHhxxmON+Stp+blnvtr
GEPl6qiF2erdhc+eVmdWaySHQ63M5bFrhucTib6Mjh0ELXCIBoxcX60V8l8HSy283fZOXNAfkT/K
MoUAKKKFAkrBY5Xogr7GlRhk3oQLXgToT5c8DeW6HNPMPg2ncAJyDVyfJvezxKSz9ydXWuV2eE1S
qV5qAbxnte0BDpD2yp9ybDtACuT0MB2GF4YFNOR/aGdQmQwqkoY7PhthPihDbTF00PQk83dOx+qg
4OxxVxYwLlKctIhLb7bvcLM5uyX911S2SJ6qLVFGu6yN3PCxyGBL7O+se2VOkcjkKofGfyPva4T6
aaaMq7USDlamhdr2x0zTnVw540qX7s+Ab5i95417Z4/Yd+cwgwnv1C99BeEZLxNzVio65JKaF2N8
VGDKLHBwbPZOsI5D6FIQ4xD2Eff9e9hI5m/2eweaTaUmsH/IK+KG6vwNQ+sWAzDAO2fzFZ1kyUwk
2gXBJAaIqFcLpQO7QGSatXfvjuunrMDVj5rXXCGq0XVTnzMvzCkgvGVK3dpDt3SF0cRThNqq2fAB
8a7fLqXQWSNyMcsqdnayJFgdUOz2LoeRMn65D2AWhDWq3l/M+ynZEUtk9H4VKESFrd96R2cgUgOI
idiT2IwHYcTquCHxjRBtJjx1A8n515NhnR6YLkbHxYQevxG7zRgu5BjuAATQLArtJSYG50OTVCWV
WNZ4OlNhY5Ly6hwY1KxS9QeuAcVjt+kQFHe+037RzeaoqkfEANyDuotFKpiNwgdVMv50AvzpIhz2
lZ8abKS6M3VkI5y3pyoQ+Gia7ICGjeY1cJrHEShv6TqEhmpfbdc6ZcCTnhiab3gdCN5HMCPVews5
xUBx1C7jNupmp3PZc1VlSXphV2IPa0gxHdtnY9/S92S2OyGsA6MTPqzMmCuFAKlcFaHV7yW+q56L
SSXI63vzYcL75MANX6EFnxhviOiZ3OVOwzDHdZcUW10SXNDOrw7oNgelWF8ezr4ubaAityfGyTqG
dkEUcyOlC83yswnJS/BWb/MWz6fI2VznoSiCqxtdJ/RIxc35UNStUqLbC55pdcyRwRXZoQiM8yHC
m0segeJY2nU077rd2/nbR6pFUiH4HUutnaTzqHZsklY55MTQNfbZGOIGzWkZZ/YzTExsni74dKgI
dhdY70kF48SiSGrRTmgzqq1mkc7mY9ttfaxwclRRIGEBxTqLfKKHM6cjdMlBMDW34jlNXbqR1IFJ
bqrdTKQ23ANBBMTwdNiArR1VKSWe8tA1BRe6QzLnJqMF7HdTZqbUhQpv/jS5ntWNfeUgbFxK0eEX
RqDdIwb2Dn7GCWii1GEi+NE7QGeWZHrHVy2tjp1uP+Wl0tAay0P6/JrV36iGWzAWummFqNGqppcw
SIPsEuNjU363ihy9kVFUX8JRGg9a8xbULwMIVsO9VwZCTZaobL5IjHxV/odzcDG1hpGUa5MsT5d6
1dQ27wTntX/A3Lvc2SgHDgb2uogxz+S1sqtuMyaRH6IITvGWdL4NSAP6RWVQmsZoFqxoTZXC60bL
u1JfcdWnlXCfDFBkQTquOssfk8fYQe+WXgqEuRjL+0BMDY0k4AGQk7CL8CZ6BJpL+mGy4GnTBBfQ
u5gGo2Jn1u85d+9n404P++qrOAT8awNOgAB29yj0lFiZ6Kz+7LCaBtNcRo6si+L2U/LDq86aQ8IM
n4ZkQsu9ErhMR+y5pxSqcSTPrWCpI5OlAEE+YtHPw+B/Tz1B7WEon0jZ5nwsl7zvs5uFSvArXTAb
FrQLWjbZYCZ7HOEL5v47xcsGvW/JW4qAoQ0O2oXDKm+b+rF+6cZzwAKohjwr9w3V4MtAXMg+HQNh
UY53YdL9UqcSxHFkm0wCf2rDof2xY8QeO/oXyaLNfPN5NougngXof4LlZivGFBKYH+gNrvuRShFt
udgY3dUMQzkAs5ggMRVMf2t+oeZN1Okv0m9Xfory29fEqYvZB+KT6Rp9K3eWycfbFJH4+KI1S1Uq
NE+csVygNldf2arit1AEU06aZfAuBREyg9gZa5Lm2VaBlpQVmA5x5NVG15vMhH0H0uLpoZioY3f3
GAmVGqWKPH17U1EWbTAWa2yFEf10kYcZ6alkLFhIdn2aGHyeFxINSPwCYooOSG2Ox3wtVaI422Bi
f4elWtVZ68Rj4RNRRALONKkDKTuG8cXmOu2QyheAZDHYlHgHLIGVUet0QNvy/rwpHrV5wpWSTTK6
izWQwgdqr+zbs9uH3qCRSNOhPCpYnGhOqWXkTWzA04wRx7+Yy12uibGnipa3iKhVi0zzR8cG9za3
1pxoWbqMfv0Q+NaMoA8fee1EOmlp/VDzT9qr7JJEUPyV7EpWf0jDHxMgN/WDLhyeVnOsqw/FO6Zk
qojIVowjccR2f7WSPN9ZflBwu3mjN126EpPq2PJrFG+1AHr73rrnAXdMOI50w38g9z5bQ1uWSYuf
N5BKebsLEeFa8DqhNhWnOOrnD6+4CQjfTQ4R+Y4Y9pn6L/zXyTe4odgzga7rJGKdK1+6jAjAGQ+5
BnRv3T/8ZYNUqFWpi09Xvyvy6r/M3047LK8xHI8+DvvKON+G/VDwQnHdKCJs/E9hje0CREiwb154
atLFVTGTBVyU5RoyjPPqS0tw2YowyDpdQ4XkCiarAphRiM9htXHjyLJJxlHgPhnSpNDjidr+fpQr
ciaghcbg9Ut8VQSgY76igw8a2b+5Mz1uhEmWMzM5QhKvWUxGeORtORiLHZoLoVYiNAhZNVuGiLqH
8D+Da+533A3/iuoSr1StNWgK9MvQIIKViaiPHsdaMiLAYbp4glQZwUlpPiYKZMinTEZIJlMLH7hA
cCHG/+Dd1k6kAJeou0pXJP9Znx+k7b/kKmIt40RQDxUuGD6v+K3j6fBJF+zTd9uLwiK5ri3aVwsk
Hs97wW0yMfUIx1qjYjbzIYBBdliYkba8kxzGmPU5Y9cYM/HaGaFKYNj/pzJxpoPPsSE8WF4i4gsA
N/wsfPnBkKys7De3T4dYjta0zqjcf9sKcywr2An96gidX70iT9/QgyePThGmT01v/zIU7dLUYQIl
ma5lCbu9zuDUNlA7eihstq7dwU/DQWl153YLTZATmUiLCRY4z5iwOYdb7oGvzfWFaeuAGacBDvSp
Vt2WQCRSerczMAY+h2CZxdsvWWc6jQZfqlwcDwo1DUVzPD784u60pWkEDsZwJLXIS7DRp05XBtOa
45o2qU/oXkQkLg+W0maGvQjDp2256fQzX7TM1IC836viN0Ye2qx103ypSnY/sl068SlVnFBPA/gT
4V22dJo99hEyDenvGGQ9NE9bsdcHw9HIsQ43AZ1ZeSWo2qBbUqYk+K8W7z3qsEP2U+7azu0ovfeu
Pg8oemGc6/q6pJFAcSaWz4ma40pKVQK10CxXzwLmizChFtAMG4Wzl/vfgzQ8lGfrHZZT9kkenaJX
734+nFjw0sxNm4eopQW10TDKa3I5UA/dAcOv6JNBcLm0sC/71/GMLnEzOan1VDDP4w0r4CIK3Gai
Kmmj9n3HWUIsvtaVJIV5virhawn3E/DKsLjjt0NbSXuRSh0koTVw0Q47/tKffNqUtnyeiv011dut
LwpFMNQ8YWokpMZ3nWiMExscI2oA1bPAzQKnGkLAxvJ+B0m57m64ft3hrBO8hbtjUV8eW7jWXS1d
2srYdQSoiY7BC3hOT5WOYPeSOZ9BYpEJqGwq53ZYjrOVcw4nzFdO/MF3a8EovKf2oP7AV9tf5aoZ
ExmhIjQAXrk+TPY1NYdAQDPM0hD/jPcPcZkBevirUtJulIx7Kc2bmgpbRWudCq+fLFmJzOhbhcHT
QDyKXnVYHZ92Fk5Yhyw8qxzVprmZO2pSIf0STsrMz5upZ25OtbMj/4MM3xV2bu1E9lVWSq8bm7eB
plsvzgnkEynhGupQPD/TEFuUbVRDLMfdffJsopSHKQjLchdzqy34Y3dcsY966wvIjGhqliAFA+bH
+r5aMDd+UjQXFpLw8lDyphlqbUkBNPtflSFzrveIMzSckrcSuICUhOf1cwkSBz28o/96LwTYB7JP
a3zhqXxs98fpqseorzuMlLyFOnO3n9Ky8FyURjC/2AKLdJXuNhMCtSHguUKWoxfneA5gyiMpF+Up
AIkNKWEO+LB8Z+9K0jw/iIt+vfQIZvY7YXUI1OnuUf1BMZ/92OCWM7WJZwocJ6q8H0CpoHFjMhb9
tswv/zoF86WdMnrk5MYBHUoMo1kkZt43SOrWho3vPq6xR3EMn03vkb17bavqzquR0ZjHm2/6aUGQ
JxOiiyy7WJZKSnNx8YrLhwzYwjhBC4rUgOoB0rJoWM3B9l0fBN/BqJozvhx8VpBx5sQoRzYMNo1y
xio9hNSrR3FyqeOaQJJ/37YKX/WDR5thUEfD6RCYOkV43GPJ5OAjgC714TBZH7VnXaUP2LSp13Nl
rZTpJDIFU/hDG+aiM+u4fcVrlxRxnr2WwFdM0/nwDZiih1pehie9UcfRET55NOpuj/l3y8WAGpPr
I4YLys/TMPYDGlygA/1CiImmcyizVqryX2AWydddukAzqPlSF2za+6o1vj6KZGgjf8NlPvJj9TOA
R1bQYMJi39WTJP5SKRdLz/x7TOfDqLsIIWxo0WSvIgKBUh1HAd91vXUYKi7Q9nAxZBsTu4OLm9zJ
gfePI4P65a7Q6Zg9N1OCLKYmM/Ium7WP7Z0JOcdtblp7OvcZD8H+EhNihCQqZLS4YpVthQRBbHcH
n5+qYcO2BpQTYDsYmxdTaEILczeUbOEm7MBmaLTwZ9w8OPRNkBYfpo/ojYp0OJu1Z541x+NJlBWy
II3IA+SH2NE6lpzujiTSTYP0eW/qlAa4G/08jglQfLBNMe3ZDQyzqJyymIG6W+ikz/IlCIQ0C9dw
lBZ7OQKXBmaEI4sh7BX+lmRyYegAzDRm/UMut9gspLHTmFl7wQ2R42pYDZIkO14cnL9j6knP3yWx
ptlGApCgYwFQwIgLUeEt+Oaej/9ZMmjOx0Akp6SS4yLrXTlD6uKOZFn6pt77WEIr3/BAvsjR8+/J
xng9iHFYlvYOnAwraPzZkAymgZoDwLG6K8FKJzZdUCz9fCbxJ1GOWvZbNC1J0rLgL1cKL+rPVuPJ
Ye0hFFd8+hZBJbip0kV+AVqykFIHuAqosegcuETkz2L2CphUSKfUct2Qko93YFh8Do0lBGJ+y8uZ
5ZC+C4cfMP1OgHNaHoQFyMAov4kcf4n5xgVxGWUsrZo4isxzifSHXR2vy9YPs1oKoQnjh7Hg0AHj
qlpGyQRxUuREBS47AfJfct+p6tsrU9I8Hor4WqF8uJ8HqzxS9CYbnD/mSBZyq1wAl0tsOlQG+YR+
M83rrU7m8l9dLo+UfdeO0QUHXIuafiOw2vzKNHv5DG/oJtN3y2TCatkcX53lCBLlbw7PiBEQ0oal
Rj6YbRD9u7xFgsNjtZT/aUBj+hWMocegveAjHu8nDF/At734dj3DmO+3GDA6hot/6mwrPEkaHixe
V5eLhGVDrACrpvrebLHIYMN556YFtKvt8Kyg/IniNhuEqyVEojF99slT851PB4LLZ2mGB50H5WFw
754ux96vpsxDYeHJso2KdiulKjE1bnORVvH3euMLmarncpxvSn0PXDlXDPoL7KllkHnkCZ1KYxYc
GKG48eh0Uz3xoYtcjEJdUijdXi2rgUSOzyL29bPKqlDK1cvARgGbZxstKg7ihCIEZFnE4PRRHnxo
AlO7vyoogVkxZTN3pM3cW3aklMUJYNnHzmyGIr7F6qs99D17+gJAyp7zB5TDEEyp3UjLRdpxyqOQ
ASldmloZp1QfoGVWtlfiH1hKaF0ygDFcVOPOAQF6HQ4k/Vo6FBp+q0n/jkbm0LopiQobKyEIs892
NFpMhQcrlEnBd3wTvQJEjSeUDqmDPZlV0eKcw6JFK9WR1PrhRI1tqAmDjRDBBcIyMxKDsj5oXsn2
DZTIX+ofK5WFS2IZIwXKfSrGi6sBcn6G9Sl7uCu436xRIe0ihLwqS6EmmAKuW730mhf4IKh+u5iR
QnCHDgNaYJqu25pK6K9xmTpMug2CEbaXoImVkhYyVAZZgNrlSy1vP65JeG6/KO18xE/xFk8BOhNf
IEIJGaD7dqimPvKnsX86I62PA57OykxTw3kdTZoD6FyeC+fBThEY8pKupjMoKk1fctdGfuJd52/a
oTM1Q6hnFLkyQvIckpDuHyvO39P1Se18qH4VX3xgOvpXlIFcbPGLJq9uEP6EFBV74qxQZtE4WxgT
g8L/kk7GD/fnelOEoe/ccDYis1LzABkY0TpCWc8vB/kfzfYhR0sWzaoXWg6saeLG+VgGlGtSyg7a
LOeQPo7mjLOJYGF4RnOrrOYo7G9i3Cc2q3idVgkNgSnIOX+NrBeCHJCWHtWv76S+Oemorgl8B293
WZxF4Ji8zeiL+mzniYECl8dqu3oCA/YUCYlnsqEn/XbBeeWOsj9BsCdgmEzRbr5yQs+5oZBqpQQP
t59sXj0OHj90mklEqfNbxjV8JYp7Jl5/gKBNdcPoCx4WhateEGVUiN+FVNe1Pc5MpaN/DAy8tK7Z
r4Gq/EnYU9c/X7Kkfg/mFGcDoBD79BrG3PJQJKlLmuQKK2x9urpbbfARNm8Po6K43Cq+385s3PHy
rN0L8NfYzX//1wriAfljBgkhyyAaBP1pZPmIr598wMwEh8ZUkG01AALuBj6aOxsC2odqEdAk1URe
ROEFB/nvW9wSrBucHkE1YI9UGJHFj9uLSOhZnMMDfvatVNj6jQ5mwl8bToe65RdmIIER7OdHls/0
+WSltjt1NmVwuto6pWl5wiWcXbHNJ7T4stg5Tiv2li0gm7HXUhvTgQMRTinQOB36esmVo2DxDWJ0
dlKa+1HiTx7hvyr7OXwTEth2VGvkYu0YrYX45+8INrawgHZ3a4Ej/nzQUjCyCRX/6DDa8fhoAGW2
maHcAwF0fT4FduZZIo/62jRRbrDSYB4+PfPlpkg2PuuELu7t/549fpLrB5puwLW+564ZRcX5Y2ie
dHREgV9A9PaNyFnIF91o3q7h5ypAL9Yh8GOX5iSEir388oIps9NmS0DfSsW6FxgJ0e7x5POkj7E6
fcmWvUMTUeP6RYJBxYzVNpr4N0MXT6GVT1mbo8Pd1uWjS6R1bIbFOAU/qWXFXal9sQ1NhYpe/c54
tmh4NVlq1GqGdB1ZBbHdHoK6HqO/11Qcxis6e5oYHXo3bzNcXJ5ztcdKsM6a3VxHgpYpzod1iMgF
/lO644eLn6bU/JFU/AxWx4EneCq58Hcaj17p/VV1a1a2tVJf2EiXOtnBgLcwiiIZ3sRRz92if6ou
M9qFpVVOSD4vt0zbLAHnRR/MDhn9Qd6bo4gq2hB9lwo3hGQtzgCqF6WSZS3jjNOwZrZySkMaocDv
USRXJwWObTpcV3NtVS5jw+sO+jXvv36RbeKHzUkmtkriYLPz1Aw/627He+Ss9116xsDEpRGxrdT4
vERb5GR3ORHD7wnTgPN4Lxg8/Kjn3xzbE5kR9eidCBVfqHCWqo4p/+qEP1aSujtadWI4F63aecc+
QE1+f1pHFXY6znX0a+4Ij6p5vMzCrIpsQv3d2kQhlUFmuRrMQ0QYDSUXy68OFSBGfurBQTVi3FFD
QmhYxCjTbOJEHnY8TeMHmMFUOSEnPZgtc/dNf5h0yTfp+92/dxaU+PLW1uX8oX3w5TdJvdBFFdde
rEaIdLAVjg5ia/jsSO/0gTDKeliBhJ0uOalD8PYcuIIgA0j8FAQmT/Eq1Bt3Y027xvqYDoxA0sql
DSL0abk7lqR+a1cwsMSitn9bAZ/Jh44QFLxVPIJoa6YQ6pjmssFaDJ8WrZu3aVtnijOu5n+1kbVK
FWldzjM4oNIl6Z1hX2SW8TGEI57iA8vMviBa3c1BJ4HOi2Q+rcXZyqowgBvOtPKxy5QWsPLNpQDd
mNvdqAkHz/K9aRpuJh5CeDUMMKZ62yeCJ7NQqDTqvqs4qyR1SYYMY/raWj8AxT4twNWHChpk03Ka
+39bRjjw7CN8cwzcsC9newpX73daqx6rc46ei0/e9EmF5b44dgu9PaDFx1aGyjl+qJNeCAWe2wq9
g7lnWk9zTC2RfSdpTcZS0KkWAE5lzmu/xRqvzsf1EwiqyXjIs8JqOS/C6+rwyUqM1LvcutpkQjim
fk1wZz17wf2XciEfe8xhj6Mdvzz1Y47zsV+x5xrnV9Gfi+eQf/Vypb3UDoD401zIrK42D2ikLY31
nAPqKzn+j2jZh1idD6bSrzFE/cGnRV6wP9CsazmhqsMJbZ8svPdSkYdnXd6spd3QTHPlJkiJwcgh
bGetSNvKCmu7IsnsEB5eppIfVs0ZaFxAqlDwOP1iI000+vy6afX0HdEZf6NX2VS2WTsj+6meYcej
tr8eHxoEm4QK64ZtnYkR3yXRgTnWmPc/qwvYH+Nk0W1kq57uOqyxq1SJCpBTAGDIKr49cA3m3tmR
kPYy4RGD337KL7u9ISJc6papQf78Z8qFCtyYmCR58XnGhrMqWL/5bAD9Nv/6hGKAApuV3CkTt6QD
V5JGAwGAtHttB8jziJOETf2cAwA57VN9v4As8ILoqGqJ9ft1AUoimizD8i+/loMqPiFudI7KrGwY
1e7n02/mL+OjaO6r5FZsVdWdfy0zd0Rq2E7lw+nhUWB9MC4mTfaMalXA1HOr4jjaIdLgPvHz4BYp
9TCI8fYPY9DA8KH03MIBb/RUvev8mDIqzAq0chXlMoKXPHovnbeSaAdGg71rUK3nCQPpffFFhNqU
14jaY8ofzzGQ8wahnsASo1EzlxdWv46JScJX7G1UEpxblbZDmK+Ulm3HqouIlYk66lpi7/Afgopy
DjEcDxwnwb0uSyY57GHmnP/TIyiZ+sNw/xO0Y7QCB749NmJnzkuei8NIrE0/HrFOgcteC6MV5VDf
BxoAXhkxeCdHw7PkdQHLwI4cmbZY8VMtwnKBQJv1WyUH2Y2ec6tKtkNMGMkgojd/Umha2WM0kI1w
mVQ2jxn7GnkQXYzI/wP5R+7jhZsP7mPl4ZW0HLJNeybTAuOWS30EefiAw5m8MGMDio1E9teSVDeU
+ZXmA6I5NfFeJvq4sIGpOzyjNK3+fgUQmgfPxfW4CisBZi4Zm9Xxq+AP7ADuTfO1YTGpLLIiaCxv
CSkYYLJxZY+xtgVhwW9iolD9XSR68LxRwRRJ3UULKOtRAuLp2BkzFiDKRdP03QJTBSWK7DNaD5Ng
S3ZQT0GBSlvicottHZDVFf3/LWBuWWB9nlgNBkkrEEL4t+EXPCB/VWV3WfwRE8iFjNAM22ANYMPd
V4vBLfydIZ5LZHLJYrnpFmXQ/FhHrYg4MRs8D5kGXPCUEQdcWYfJf6jsIE2xf6X4i5hW3FcEXJpR
x/nuq6FzKjVuLK1gO7Mnb9gpg0nzY5/tkOPPAYub8y7otXh4M0Tke3AvUe/zn8hqQtnaCzs9ms7v
kwHxl3GFpq5GYXAGGvqYvRfJvCfDH74jm3PYgFxjwjfe4K36F4OTfxCykKnrHNvcX8cWcQSZz6yR
q9MuEr/wYZBz186zSWwg9cyRT6lprL73Mqx/lUDgEQ1c9rly/m1boR0iPsVAEWSJvBvCE1AiLiU8
riBiXDBTeBuVQ6DOCHEEuRDHeMzFf3eiAEbvPyMRycHRL4KKMsSOQUTRBgqmFZT8aitD6DtUFeCG
MLk4I60ZGV8+coX5SsOrLoTG6k+jkzTtqQFGf9FOr+4GD8TfGJNXSv/WIXmjNXf1dvKGuTBA8DpE
XqchlGOaAh3getEuxjIVc/VGhCkt8+zZgwE5gzx0ZHtZvOOhsN4unfVhAEnQOSQn/hsnVEvYqtJ0
tne2S42c+a4LV3TQRBg9sl6PxauTHx1UR1Rd0PuUdQJGCGQvTi85J/E3MiVA5MKQf9hTKs/5AraS
INCgKvfpinJ2jhNoC6BpWaoWnM+gM5RikOXTTXbjmd72vkz3CE2UM1xFTcWJ0ckiZI8bFiSNTsUe
OhWrTPQz0N7e1cL1v7nT8Skdxhf8hpDE2lHnVV3GHdbF9bsyLmnYIS6sr6O0ebEwh+B+9lm6m7+k
pvvLENlDBc4z2HAXBbkm8y/V5EYsbxdVuwCO7oP/LAlUsS3acVqkYAy5UyqGT8IjbsGvwQ5qM3Pa
U3JoSgLoprS0PWxj7Yv5T+OCnTjJQ9+RfMjbAgNxOAlSSiH020m38IrA1nIm+bqGJVmn6Mq2uIO6
l9Ipv6jTRg02cVoNwoNhjqrqM7wUD9a6WOe5k/9qw1pEOnzD27N2572gFX8RcyKjlcCC4s8EGuQj
h1ePG24pREPVsg/Pmhz/9xd0+xOa9orO5nB/axbG/Ib/XQAK0LKS7BGo2hRq/1VK71K3TlI+uKQS
F8TFSnog0L2NJnoxmTCjjcVxGmvIeXrpyKoNaetAd1fcHOsyalhmhz4MpE6COqVONV3ep9SL6cFN
dIdvCIv0J35UFUYOq/FWOxQiphKqe53XpChINMSf+LiOOuoGWIMCRe3tEl61KjkB8aRZruCvt5RW
+NO63N92GfGzcZmGiN2Biy7F9jpouOe8I0nQRm8Rtov7IuISHl/B2zYn/xo4cBLFRtyFI04S9YO6
E2AFuhdVaSI9rmeVtgePyEg5WovETAlOqorTQiwMsbPMOucStmf1mcbDmz4pHrHhTblQh9vPJKdJ
hEA5Ikq4HbRSqp0DblhEzkYJDsWcfJ5ofRqVL7njDel+8+/DClZPNV2lIDrZT8PqGg2LW2IsBN7e
ZWjCtFGW2nor2LMGse4SB9crdMyFrogzCOATUGRMzLjvwzFeS/WaITRoAKsbg6bGDqRKIaeHBxK3
2ytROPzVQZSxDS56cdgXTvN1CAZBe9h5pLxhKXWjZEVyZZrBFyXTv2CKJm4Y7zozZjReChTK3VE1
i2/QtrUUcYk7cud3v1W7ZWQpBjCwguhjju1fx85PU+vvyIqcLV19oS1GDp2LtAgoVoqyy9P14iYr
g559NJdPUejlNjWPFS6WKzffxIRkItFEonucYiNz2azPO2oid7v4Vhm86uW17/2YYy1LKLUok6V4
2T84oo0y7ANtxLdqTmt2Z7+oK/AoQIIDE9eVqzQtg1tyV2PMNQHXLw0eI7AQjnMx2VAogV3VYOIZ
BHOsvCcyKLgQvrOkhcxJNdbflPEsKUoS5meT0LqOFfKWWd3WZGjUxkHmRI/H56gIzMptqJ+CcSGy
P/vIdchcl5jnpXCqK77hz4zV9O4RJAezARm3v9EuJwZuU8KnMfTcSP3H9ewu/INfcVVI4oxZHP7q
+SHhEOJHZT/lDYYbS8Qs7yhNycEN3tZgufqklTHvSnAkVV67sv5xRxZySBSRa9/2A6NtO6dsUmQB
rlidHHQ8hd1PLppdhmpREJgW9DtcT7uIkwvATqmoijVMGAB1FugUWP5R72TBeDhx4TSaAqt7R8Ty
TOsj/qJvBgORYyHIdSr632/o/bSaD6mhVJHCvIBAWSzeiLkJZXPVWduxFB99XD/QGSA6Wy1yqyzN
G5G7jJ9eWv3o3IBtxnZuYHR0HXh7uroSuHyAD8hpK/feUY4zMgzxXIlV7vbMXS0Qf6OMZghjprPW
fK7AIr7yoRplkjdQ9DX0iso6bkV+nTZ3MtefypXxRrf8z8S/ak0q6cEWjvazE/WxvrwBI5XWuk0y
NWeQwjfk+lba+zbaEWtbBSmHtA3nJYJJ6JGNW40arpmiv0AGTj128ZgCJxoieNj+MWB0G50pQkjk
A+URxW+dM7G0IUgCKjqUs+yTWEzhPZ+8nKRVHr5BBn8diz0XoKSHtyCO69GM77373ylCW53PkHi2
BXYwrZiao3+qM8QXbgZDACLikM/852RKhl7bCW5kUpgN9xzFNB6UqvBlurz7sYDdYxO46/FEfGTY
emdX0aZlP6MP0AqrYpBtYhgjRNqX1unMGAznekE19D0AmIP3SSgShKzxsK1Gq30JkWULgSPE2vGs
na5f/F/3TXzdZUUJ2iAz0SL9BqyS5JoQXaO/dNmWPTyNxznR1+MNkhPHLQBuR2l7EEw4taJVB/Mp
rBSN1E+ONG/qfINkFnJLpxnaHok+lB6FqKi6ukBZQWbCGsv4u420WrW2pwxND3wmI+ZRyIRUjnH3
1b5YkLOOYOvIgdSKB8FgCevfBW8Kz48Jq6xYeA+zSzyoN0BRV/REwFh0Z4nSp8/yWnp8L7Ip+1wZ
2Hb3aXpk7DiiTBmJu4lsWur7BOcrU7GZCTyW3Uj13pUfnmEbY4EL9nBFSI72pWLGFTnVPrBnfEOZ
Mtps82x7B3mhnlr5BrXN7MSHpWS9QMhS9CgrgQwDfeLug+zDJVybGXaKiqD/sW/dN/8N5g4g5qHY
VurV7ttXwOeyjIJndEHCuDGt+H14MHDYukev6/gkhsk2r+6bn6nMnTzN1CFGOgt1//6eqLr9xa9z
6gThFGxfI9EHdP5VsTT44RbLIA/nEdXYIOmgFJ/S/lQsp6QdSgF8kJOrxXCXO48y8bkHfjTEkQ8d
XYtt8qmwbtSypkWIEZYMTBwZ//xlC259h+7zxrjBKSZbGTl1O0Y1EsGu7Mr++7/XW5S6eV1b0ecl
m6BdS9ksPdL7Ei/cYPSGq0thQh4FfYBid2a/stvRpps5jNFOJcjzBG/hdI9iMvdzb+NtTEUBJhed
sNK7ePG/amBTorXaT2N/fh3sFcadtqEaLdeqxgoubAgXGzKa9J9eEEB3a6Yk69qf1KNxzU7l6Jfy
YnerQn4vWYivuI+7vy7ZIBmP44so8ZCobTsjMlmYpmbdTuKJohBZtDlG70x332al809PjJqvd5Kn
n8KqVlUbGD/b/E3EoD9viZ/CPxvKG4bJ9w6ik4eDy5M0KTXhvbpeNyo0+bYNbRo1eCmsGUj7CiEK
D3/P6pvF07szxcNA5OJJbwb+lcEvfFxLcvXUAEIIMqYREcMwsYPnGQvJlqZrgnBchVS86/4hA6+8
MyvCH/TUHgSrBVjDC/7kRmV1i2dUk45QMIYoA+Doc+pWKNj1n7Q8P0775UEJq2BAbkXiq+ca8mZS
n+xwfbHm2Q1ysPqtbkxEVDz1seqPfK1qxDWqfQ7aEkrTvAS3+6JSEIm9URaz6rHtsjlO2tZoAYjl
cGT3KN2CjbgjTdFOPeuBMUMRWpHqdKkWqTEZdbro4aggtcIIe2g1PaPlcdHypvE+PwcUFiEUM+ei
6gwVgQan0JF3monIK0KMcL3pHZiDwb9K2qhE/gVTUetbYC5VkHb76ksX1phUo/h0Nwth2qhQogZs
47KO4+NOJ1mXWCXjD80FGLH0FSKibvbNAyY23Et0KaVokmdUnqZLeZ/mprsYaIaUP1xEJIaJIClA
7M05ij9S6KcT0UAYoKclsCagSR067WUNHPW4f/TsdEtTCevdiMpLHa9btn0AddDT8D7Qx1HRVOyn
HVDpAQrR2ZzoO4JCL0c8JtA3SloFJJAyjl9JcK0LaJvdUcPlqw+q9wpRDjWuQaEtIfGE9Wcu0kpt
HxjE17uyqgns1164KxxrPGd6sLgEGCdOQxkrThXPAj+58QKqDdHT6hPla65IcIuVLkoB654+mfri
lsWntn7LHyLBiPhb/aADCRb6IkiC8rLiJ+0zD4Dkw6hYAvjY11i6X91HE9WxwOkugFe/zEBk+Wyt
p20PK4+pPYXcdEqlU1P7QPcvnR0Ue3MUk3T3Mr3nW+jR/snrRiAUdcZ8QFb/H+4mg4pgUVurjocE
H4Qd1No2fwWcuVIjRpiurcq6RnbQmCtUO2vPqKOIH2D5lXEr0TEqx2JZByAnnq7R2+fjzw4OwFmX
51ICLYvxrm7FsCuR4wcRbDXP81BXY1AHbnh0MGCaWlJPMOJFnjwmGmagstxNAs7Txco37GI1jqBi
yP0KBLP9VGxhMv8utzUcE0bR6/jokdFt1jZPS0jdVH+mRUWP/dqr1Ev7ggENEbmsbb6/T1zskNCL
Pm3m+hTKAX6dW3hLk7VKvvI0jm2oP4DmBogdBOu3+ZzgVmlF3LFCmfYSeQM2A/h9fDy5d8F6IYDy
7tuPblDxj0Y/IExi5tn+b1a6gHaFBSk1oI75Cf4E97al9U4ZYg2I0fGLsSOfk7RLo5sMCWhpYLed
q7Bwk429UGFmCUd0+5iSenhonH7M6qrl2hiHsWdfKvwqLxE/l3kvPCrjyn6NlowT22aAQyOVVJKf
Ndu+0E+qXtgxf+xqe42fManUE1F2BpxPYcOZN9bmgJa3jobVeEkUNoen3fwmSVUs0pjfc+npP8tn
2kn+ecgolR/3zduc/6f4zYg2C1KMSTmevs1lXri0HLn5jDiHqSC2HarYqeUA2hxFqotkQkEIqYGx
wD2dLd7HtGRdeIndnhq1AQm6wz9RIPfri/fIz4m09rJ1aGLAKuiHPz2LS0Q/cSjFM0EPJk42Enl7
xoLASCc/HXN2iXn13/5fDcNE5HF/b1jeFta6VIZxizza4boSoQPQ12vXhktFVASwDcnvjQuz6bar
kYWLQwhsegw/EZ94bZoi25TqUQQRhNcNMZK1Xly+dq88MUC9i1pvqkpUe/ac1WxiLahD9mP6j0z8
HpiNulBi/LgXJ2uan4tSPsE/GsAXTWnwa4fSfBEExTM1In+UJCQgTu3ApexUZfkVSEVg43S3Gws3
U+iSe6393xpsKzuV24zfwK9bFW86x7KXpglM2jGdk6QGwrDqsn030vUOSFWv2imooxf8XZIaZU4W
/k0H518uChaiB+3VGTEu6pA6OUx5vBrfsXtvShutE4NFQB7FbpCq3ox8j75zCE43zQUoj56AR4Vz
05lvnvnKgTBrYQSxq/zhH/51/VAt7/uPdj8ph1WtDvDKecIz8M8a+NvQib4U9POYNLuLFIGnKQlW
mJHWnMPVcSlVmwwXqqnwbvPUGN+qS7RQqCQMwwUbvSRcCz7VxggcMfvNL/jawYVYWEqVOpNMLk+M
cWOcgqPgY6pnEolJD1mKcY9asCJpQC4ik2r36CIYUFgV0x1yfXMTqMkzYSvZsvuL5p0t+lDXNa9C
qtq/fgbDxDmVVbvhVG7OHn2VrNYq4uR4LW4pF15cZIcbaicyMusTEiT6Dzjb0xUTVVhMuzqao/Bc
om03RYq/bpoqLpqjQcAgmg52PhIv4PdG9AUEzUKzcnFRnNKC1N3jRrB7m/lbFK//WuOrgeVEprlU
cInoWleDdtGDaab44rQQCLUzo7L6yzbz0d8wUYae2f/oxvDpGpurZLXUOzN0TBwO1GC8asDl3LGH
DemnjQZ6TINOoqZ+fYnsTnBBFFiANKd6RCdsS91+vo9dY+91mQUx6cP7zFrPS1l31nSqfosSxZXf
RPvWrXbQFU5potB66AwYmMPcH/Lo2OWXAroPHitB9+zfINndtH2wPIzwWohhgIrwXQjL7BfXmbol
9guO9KKSyfQHZHuFZwPpw45PWC5KF/ziMEPOTrGiJvzSOKs4TXUDjeIBaw9WbzKGes3PqBzYrke3
k8R5O/pzuO2IfWG3r5MInDOYR7Y71NZBU01khSNQltlAAtnAouT+mLEzyPFzEix3uBKR4rIXnzwK
Uw0s8bE3ffmCfyedXf/BDOUMShtm7wFQV5PLChy0skWLmjtWyAaQFwvCwtc9aZHM3fprpC/i568e
4KF+qUDHdbR0tta6mWhKc4r0rYudQEY+AUiaDDhlvwU2Ej3sMGDL6r3rFdhRPdVG40jNVL9IiWzp
rFYPEmfu/hEFI485YJ6gYyZfqjovA6aZySclLR6nJoHnqrXZFj2aFGLsA0Qf7RAvfzSylAbrwWIO
K8TvTtuP6od2It6v5gqgzA6NZb3+VNmfxk+aJISdTQn6ceBKoBddSyW72F7p1j9eL1aQmIe1S1IU
rJOPE/5/ZestW3wA83BeU+kkLSE6HpnnhuDZxkWtG0k2WSx41XbQmR8aTpYPJqCEaW4AoQDR4cxC
qIUu2VkFZLDhme+hn/mmRvUXIfAFMPHh9R+9tzZEKFIogf4n95WLXrDdSTM8/7wrYjgmAAKC4c3/
NrxL1kfH21bDJaoGr88TPlwkPjgtDCnA9sWNUWuHC0YuaNJxEaAm7j5kfAB7RL7VGcR3Apczp4Vh
3F7OG0UrDPxORkvq0F51w0g1ieLFEyzs4oFApW0O2MRGXTULHLnMEUmWlHkTvw0wMp+Quw3BlJqL
fvIeQkOJTPN/mqJ2FXCvhXoo6NxOUxS7PswlHVMH4zciLQ2bUwLYybRD8u2ZAG99173nMgwEJvqr
g9GwImdaGBhkkrls6pX7weB0WntNbi0f8IlJQ1tFp3SIA3g6R43ke9+dz3Ig5C+ss02XU6ch5Hi3
xbFsNcgIk8bVZhV8OH2X3cHNdUF9N4robSN/wH0GJ2RMtKzMvu3dMlX9QmEJIkacfDsV2zn0/3Xn
AVY2qMYDjoAAatZeMy/O3p8zhExnc83xV058ZcrykGBKs3NCHJ29vmAO+4YbkY9v+S/RmI2gBuFd
eUsff8UoT9iDJ8BPsY8DM3ZmOeYbx6Ow6MlIIDxL3BdTZOXDzGxFxt09s9be7uiiyP10WYIax7xY
vL15mzEi9OJ2K3ypXgI0gHagVs5qBQhgHjBDaT+1J3jq6Bptzwc+lrw7RrGQnQzWJSOwILRUzF1h
VaOJVJHSSv9ELyX1+6cS/2Awe3kv/C1G+9FccpAb6rUS0llIMw8Ai7rh3gm0dIxcLD5VYDt6u8Tj
ZU6lXiyjJeX7doQhlZNO1iylr3RXFvMXaU9f7C9INFrKJEPCatbuN4KKXE8Vwpa1zCLVdc5lQSbp
x8qQzYD3tfeEtcBGgOJ5V2Nk6K8nEsjfuMAuY1WqzZWIsNZk0qknIi2l2j4CN3Pd98SaXRqo8Eo7
WLQtg1QZ5G8TGmzVwBGy93irftvejuICmEiPJ4+d0XuZ9x+2uXZeM/IYSA6u13830D/ghRfXyCNs
vDH9nacyrpi0qNc+DDR3Xy7dRDojLVzlX51ZG2lW4U3FDoanhjyoiGKUQvpTajagED1j31gyYyzE
yfTN+6c2gLtyWBoX+Wd2Gp4w5Hs1v/bgBzJR7WPGXCh4qZKjZckLqZ7ZVYoDPqokZMKsTWcb1/Ay
64v/iQyELFcHnSI3dJqL8dCMVqxdOfxYqBH7Tn/hzyzcLDwR3R/51Gsb2siQifaPcJstVcftD3PV
SUdvn/fGhMcBGgKPg1ejUKqXhzFb9gXjRN1W5EMN+w9GFp9C452tzggWapRQe/DkIBKJzH2hjh5P
JHY/rO9rbErF/35NVo40hVhH52DT6Oj8P8co3mo6UnpyByk3VDrfoCfikp3lpWNf7P21APK+BCjf
oMQmjMpH1VvsQ38Ne9LgRP6eGJ9PkeZId2jbsbCrNZoVL8nucaHv8te9YDWL+PPZ+hU1V2eulPGu
IkclrkvtdWOksXd2YDJSVNKsJD5S6Mq1biD6yXgTE+Mj9W8R4OByyWL+hirtY8iK2recjza3Tofe
kYIRgSnNcnX95E8tfmsoSRC0COF4GB6qb3pHQb0WNdpel5RgUagOxbry796v9glfaDCXbQ0WEcPR
rRBCfefNo6A3MoQ1bGmnQ4elEgVlRyGjiwRaLWxijNhbHMxQw6jOteR9NKBVbhrFWVpOMlfCPMRY
66ERpWitKpE5CKctr2UTCJEagtFUbDTbN5b/ZuEgj5twqq5qWZK4nPEFF/UYzK/i2tYRM0B7n2xX
e/FhuruudTmQw6PdnRlh67j+Ai3D2qcEIuTNtucMHIzxuGcHkonkwoXX6y/dlGgV3DZvt5EhxbBb
9+WYc6GWWUVjJub89grF9fZnD1VQnDyRSMkdWZBGnkl3d3nfR2kPvmiKchTso2GL8J8YeQk4I3XJ
6urfvx6icNo8/306ZPE2wcHwxd0Zi4+WuOTPvRtDX2StYXlHeevaJjyMImENIojGmGbgVgX/6/zv
nccOGu/eMX82J2pbxibvtA69oqdkuwFU/j8aQfdj9gOW1IDN2fGmUBH538Vdvdh3lai3swCAmxV0
vw4/45RFxIqI2BjZrC5HC1cvVKl+EHtTLVb0dFWwy7VmmJWjlsHC41vd+kgJV4jA8YDiHgBmlxg0
XeKM0bvCZL18ZtPnvEx8bk4sIqqRor8qgcBw4nf2rMY/+AZBRHwgPsLBrCRmlN+1V9lP11tseG9J
VLCUTYLEGCPWa9utqdgdvOFOjslBe5jUIBLbKj4TFJj1iDSFKU94SmAPEdOtZWIeMgMbyJkAbrDh
RCVekzIE0pwyJNZ3oAkuZNORKoynuKfneSTjTQ0fRTn7GuEPF3aRL/ps38/e+O83ojaSR7rF7Ddz
WvZEmxQ99b1tr4aPMSWT0P8HKudis/hC4pZ4NYfy0lSLQjfTvCsLP+gcW58Ba0T3EqVHgpCcz0JY
Gpr7n07ynCNBYQZZ2KnAn0KQlQdrdRx+M6ztUZ5VEVtUEOP9VH1HAdx/17zthXJot/zxi/XqLDaP
/Hcbs9urQsrHA6vE43VyRUx0jxG7HwhJN+mwQfwwBVfVkQgTxUyg3+nM32VBls6kHmvk6hroWV42
plakC6ybjifrL47Ej85ZyMzBQjswvsVj7J5FE/BGCa1jP9dvzIp6cKyXU0yF2SZJo2pig7bVmnnK
7PYM9ItdfO3ai9NRFskq9aP456TTWwnrxf1dboVhbLhGJ9s0Wmk7JLvOxE3BF8EjqFumrVKKa2Wf
LBPjVr6t6MQXU7x6VPUmofJjPX/XNuakzvxjyEbNE5ddjchfyuADVInBKyZLqAC63wMEjO6gQQ13
xlQJfi9OG3g4KGFGKoFojWNBJ+mumiCIqAfPp6MtwQQyWqm/IXZSiurMCYJZfMCj11mVP24kDCJT
N/rOOuQEMjRXbu2ErA0lpa7owp4QTPnOWwmOyNFd5RoilcTpvRPtrnKx/p3nI91HwnKxQPyjnTuc
1l3hbwy4r5+c/xpaAkMBUr8q395d9Wy7jNURZAyaailTuH7nQEZIeatVlSHNZ+FrL3jcWKvqkS3d
/8sJ4zsgSrmp14ypNxZIwmyKpIA237QiO7uPp52UhblK+gHr2RnBN9JvKZMdiIfcstWQizf5hOSm
wdXMb+fwYlV8XfaMkdPgeVyPQgKggbtHJXAu5lxRu7TS4cF7/GCsfTUmUHDHVC1PNpaICisVKyMy
3v57epIWJIRuibQq3QgGD8W6IqJwQH+7I9FRmY+RFrZ0v3/yYSQOa86+GPFaaKFdV1EfsFTQWKh1
irvw4i4hMy5RuHivEaePxUDRJ1US48JhZ2oOZuGwLMdFu7BR4FjhJXKRJuCOp8WUYsw8JEFq/rxt
CFkfVKNCuQxebd7CETFcAyVj2ekGSTBPAxtpUlzDco4EdT+wQKIJbWcu2BYC8VTA0H18bAb+HYec
C0wm4DrZUgTkRM0Sx3M6kW4oq+dyAup1AyBNYY6Pq4rtees+SspblcOKtPhhy0LCBJ4rOFHffhJL
x53HzP5tseQwA4u2poHkshagVNoOnNdMVZlWltzwIRsFl2moMxmcLjlN/nKIUSrfcPwDiOYO8Zg2
/ykxnxIFyVCQin39LHh1dXxuK7H4AbrhTzUhq6TvvobZEri+rvqaw9QQaCZX1WrUMWoDZx4m4NSy
gysSht36tBJgLEoeTMGpEhQdIgkjoxq96TYPxvNiew985IHcvX/tP8KIWgi0wxoRwIu7YyzNbZtk
Nw1KNauW0qthBX5KQeDiF5JDZS5GoVx8LHeNnRAQqkNWEwr09k20P/D6wKUZrs5r4hIPeZsfgkNO
JC/5FmdwxGLEUxXy41l80+uwDSi7WnJ563VXBWUlDqU65pI7urgnxlH8apRy6KbLyEU/mMmbuI8H
NVtclgJqIRJI1XQR67021bgy3JDJkEXT6SRLPzL0CtShJgVmbesU84E7bT0RM1ky0LjV+InAQzBC
uV553qStHmfCNyuZPgfMxKvioOMY9De4dnPxotk0rfNsGx9BjYfX2HhfJC827rdI7MfxZTbldJTd
Cq7Bdu8TG/nOW5/YFGXw06SFJFL6Q1EBOEeK6o4RueCvjSGS5Dy4DDx224xIui8OyEdd34zps6rc
7oNGo7cFskju1psnMlZSCaDFFP9RnmiYdzjCce3g62qX2L1iQ28DuSzfSXR71jquWM6jjHAmTtlc
liCV2KNH39CRxD3c5yZHtbd32X5WzVbjURtVIvK3ZIRqHtW2BZdwjhKo8OGUPgjupMwPZtEycJcz
nLSXCu7bafkKHEKx1ibLm4epna7iJNIEsNfwRGq83v5yJXOcLybqDlxAdbEAAWUBTI/++1Ag/eDA
az8YOs1n3r7PSa+qBYLKqetEvie4hXTMII54i4b6k8W8yjDEHyqpZBevRxOqgJsP7dEElKg8n178
YEA8lvfU1sKDb0+lytiydxpODC9eVAPG0bvistyv55cY8d6WTV2PL82a5qQsLI6GDpSDnAGhbe59
C6sf9uSrvVbKbxyiPnGTWHWXbTJmC3q+Rue2iV9eIJOTsFENzOfnCO+n0WAiaOlVsoOgXYSdnBIq
HvHitjOU1Z84a5hkg5Iif6jvC5ecfXsL0ad5viWHtQO+5/IEwUzpDSvU/6Ufmg2U858bd26S+02x
/6BOip9bl/g=
`protect end_protected

