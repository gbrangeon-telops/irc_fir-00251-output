

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Cqo+FjfIOIw/0Kghh877RN5JtWmUPj/KfIaTRt94dXWp8zshF20HfBCWrK0/KjFcQ6xaC5bYfJZ4
kTgDE7VoLA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P76DAxdsqqBm7Dhm+Xv4UBWtxeM3n7VV0uwUkGrQnJyruFJEvMXWtTIk68wS1svCurmxJblglPTM
AUuHl8lZTHelg/xsbfqIjFFpkYurRbfQPaEBBncWEUkGXitk2MsCEJd1XKoy7X9zf5gkivM+Dtc/
HmQtcrnx7yMmBEFf0wU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TS87/wLvg3wp8BEZbJFwjKct5crsKQKmGgle2kFCdS51Fi9lA3booRtYf7PKimLYtiDNKzFnNmDB
yS/M5Wwp3OXdwvzTqi7m8nPDGJzv9CPlgJYl97xwwfb/xlITgLx+mE3FLNjQYh1k2fW/YeWIYcJ6
dHaLGRiPpSzATplaiEnfWr4z9y5Zgw529sAAgbJqopXb1oauD9xMSn+2U51TKQlk6QzJOyaBGs0Z
cYN8i3mMrSJtz9+1CorRnx9v0S2lY1WHtTTmGGV3GXP4WDMI7lTnhoLYTdqSlyv31x9qhFidZzgn
WXAPS6oNxDavoZXEycPxfYnQwSx2gi0tzG/NZw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NpAOviX6Xvaq+L0foSrleTOrW/NGnS56aJ5rqqn2Dmt6YUNEPYGn9LoXqfbnr2nu7OxEo+FueCzR
GTO3m2J9405e67h9qARcSi/hF0VUlC6bqx3PVbV+Lg35W+tGaz80NE2OUHws+A7UXDQk1Cp7m/EC
XxMS909JUlXKjJHNQPk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P7klUwNMTreRZK7TaA1WE7CMMEOTtEjomJfZ7pHl1XNp0UR69ZqgBrqFP7D39H55daou+YH1hnHn
RPI1HarNWCxtLMV4hOqf8NjoCFBgrnnB0U1fZ2Lr4Pjyi28WQhnjcgxXDHuFaQlXuyVOq9XUsvMJ
ssrZQdiUjtMyy3njm+Pnbmk63891Ob2bUkQGGCsGTzQYYho8qCUxVS8K3X2BjFQusmuscPspGR3O
NvboEcmhCLzlJh3n01BooLiI/MFAc4YbNKfLIovvQV4EihZ5noxjjP5wWP91DT3v8RKOECGo+vl0
XfgG1PKzgtiiXSw82pyP+WwelLF2xj1qh8+H/w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13728)
`protect data_block
3HyNHJy64jyQgf6OZzGcRHyj4dVcYsCdFgyWVHTiwfPUGpJicKLWMXSRosER5UfalkEplLWyMQuz
IUGcYyfTi6cIwXHCLqy7rFnVBKTEiJ2Z83hT4lN6JTTSTuKPvXVzslxwwxSkAR2ypJnj7AcwU03h
6lwjJGTMja/K77Z4vi/EiCfrNMIXdJZcNvsltyC/rbV8xOaRAHEOWODmw2+uHuNJvVIyPbvhuiOU
rmEhSTGUgznh7dQJrLayjBD7Kplvj4igPegbJkMjVNJQKwWvTteWp2x28QZHWuloNiUPEnBZTtLG
HOOYvGLW5lFdyzpOCMNMwhaDNG0KJh0n0iGsQrGJGojj471vA9B3apzYHF8DIJADMtvkvAwm0HCt
MhksQGJn0sRX8Z9uDLWE7tp5B3ljXpxt70qEpHAtOiRx0u99LzaAPQpCqFLJSqwyRpQZx7Xbr0bu
ZvBXJBOWZrO2Ku9JOPcyO780IoqKh2SJrlYAbzgiusKVft91frqIP64P7JmPMInR57cf9/z7463R
22aABehLBFA91zHEMFksgOT3zf+5U4zM4jHV7BabaYLs9+lfEk+EX4Klq8/PEQLQP2Oom68O4mMI
7TyUwi3Ra0bSst86bYGkQF158cPr5YgsfxifM4eYRtngIQmMeqMjyObDqpj2v+JOstt/R+qwsgro
sMZa5moEmbrrRzOxB8ypimKRAvcqgVaaWZAahx65KbXZkBn7bTtQTZgFX02hnyeE4qFlnZECyhBF
r49NQKrrKoqi4+DagD5X42DOdj1LWtZCp8LoQSBVi6Y2G/7iJV2UOr8mzzdPArHRpzcDkoFCWJ3C
pt2CM7wiWLMJdF9zkFhhWPhfWXhRWRJ8LLH37H870rX+IkCBhoJlD0kKmHcxH7nHT4fEE4fEP1ul
1dKpRqiGBzSuTSGV5wXU3A37ISvrVYNiUoo3vm2WX0M0A+d2xUHTCEHu/BFrwRauMU0J1ks0NXW7
I81S1/krEZ5iKIb6vgcPbiVPuAgXanDJj9n4Cp0rcVLEzYYUmf75cNI7Ik3VD6XN8Zyh69KI6cu0
B4HBia//cbY0L0JFvqJ+tpIyukumWHlH0g23jVSv1DYn2MM8nBnZCLLz1L1eexJwvfdOD8tUisKk
c4tJDLnIcLKNiYWVz8qYmj0HJUgs/ZM77yHDzdyT7MWRb84TvasGZBVb7nmFC7tsub3EuxBS3z8A
yn2atEz/jgxtPNkHm4u+5oQREwqO6lR/teWqrMgP3fEATYpMO53640RXXYddsszKfiiDNUUeDuiI
fEQqy2vYGjRHcHZdfQ0j3Ad2rUkNizl2rEuYAKsGO5nqTx3NFr4YUie6Q2Vze87PCQhhtI+Jx1Tp
kXo1WRTOOPcbeBs+YoJqdIfK+TIsaaMkqcqn80aE+sVhelg9uZKGaYXDiODNIxJ+aXvDD+E0+zvZ
WmOIDqQvqsG2LobHrq7xSSRRCTAW6Ijm4mkdwwCd1SS0IbNr5laUDCSGm431UEyLu1pEaNtk0Igq
DV8N0/8TGTtz5Yrz07JPW2MSsrnGOw4WjPgX1FKlW51OMa9izll9uQ00GfAwX/+IknaDUOMhe89z
qlyPAlb3gtdv0iJyZw29FM+YukfpDFpuCeOPFYe78foOQLEHv7lHGfwfOJXQM9HUAANENLFBsxH8
DkOxH2fBGmyi4iZRrJDtZDX6lUpvCU6swwkJx9QDZNfuu3xXkLdsOb9XcqPv4CkEiVfUx+nUUZ7Q
QRbYTHkyHdwkEx9mDa0lGRs09c7GRB28ovfLQjeYqZgIyDL32kCTKPyYgL0Ueuyz+DoZ0GRLbGBP
lcEa7HPGduRDUkzv/WDi3vXKxTIEvQyY3P85ej4+EfkOcz7kGN1BBiOhm15BS6GVA3tq6NUJSNHX
qZDqvEdQQLhSFJc3dBI6ltyTDCikhyIVdMxuHufJwrGVc8cQSvCrdlHKZTedvBXCB8gve+nFoe3K
wWvwOVoPw39aqNuIrxmfYdy1VudAMyvRred5gPlb9s53ut7NMoQQJ4Dwxc0u98JcFvDc+ukXKFu4
1HbO52lgWbG4uobBrNT5BEtK72jLTHaunernICM0VDRjNmm13TItMriUb71APTzfWw64m1TBgBGs
Z4sBt5qIb23gdREvf2eHHMf959y87AhlgXud//IMf2VRHdkZfxBSsJJe1ahrJs+OWt/5hfSuFu8f
dVYLZUCGnSKU151qcSuGTu/lF1sjweGq1BJHW8nFUV3Tftamm5H347p+vZNmvwhduRr1/f7Ik4iS
298iAYJsLPuQPEyZdLpmApl1D61FXkBSt4NMvZumY9xFEygMUjX7lNNJcg7/2h3GqEYP86luMTQL
1aaEln+m56r16QLZZ9A+xxjcQYB7OaP9i33g9XxDwUmqVKqh/zgQOr/kSKLtBBaTTv0fOEMe0qVM
KV0xb/njRqcpukDFrZmTnkCyQwz6QPvXwMjCxgRXZwbnNrA0XbYHM4AbKnTo1gTGSUpsAfRKZVXY
D9vd0OQoZ9ufDuVPUrIx6maQe8xYsvGA1xzqj2Zi5DR7xCO+Rw+oRBrpXXBT36HVZqkexJMOOmEr
DgN/H3UIo7o8C9Key5Ia1tA9onmsMNmKfbxXPTP31zPglaVRkhfbB6LAn9owFAuvqA1IaUlZd9vh
mjYwEYG/aAz2lUUFQGKwhb9mAJCY2QLjKWLS+SdWy69LGh2zzv07Ajm2qngDmS7VOEW+Pdw4Ttk+
+qlzKC/why9MR2wpDT+21r3bsD6geDjkbSJnikXOov50NEnsAFURN3qFqPrMKisnEElIrBSbFYGK
hvN9yY3Ir1KzxPuts4DKUqnntXBd8VYjCZVc/JQ14BN/FJBPqr9NkYbkYq0m2lw4Rh4fJBMdV+8H
0NpdVijWsITIx+Gr0K8dkNleuajbulb1pOpijUlBz7mfBRGscYh8vyU2Nn13ByJAbUCu3xeTvMfh
7cMpHiWhcFvxKR7Sv8fqd/ug2L8eV9EZrYndu4rUFhs6ENmETU2HjTkk9Dg+jrUSsjiEkjnBw20D
9AFHa7zXyen6h6pHmHtkC92wRc8ZxBVh4YnigVG1UQcnerv4o58H85o6ILQKNLeGZFKFjUnmPKOc
Ixk/9ybBIcIz+9tv5uJOVr+xx6TQfAMgNBUJa/X5OP1IgJ1qn0//134DpRD4NetwZ60SBX4M1Udg
gmYX1FPY4Y5dM9QhWK3mLjwcw6+0kEE6fKBHvCix4mH6zRXJODp+IZqxpqmDArZknjDtHvvuvQHC
p6JX/5gkfKHP5QW6pVNoQQ5oY97of0Frhq2UABp4fiCRPT/sRWooRPBZns+3VkKt6NCKXIp471so
8gie2quqO+hzjcurVM9eRal/ZCrDdtEJBGpdPuZ3Mb4MZ9blG0CkVPtGSiRFSIIEaR1MUkMjWrEB
qD1CfwFBkyQI+9+khlqE0UoeZY46/bUUB4aqw0Jtk803nflNb4U45aYTRR1NljsbD4fpwbR1VwaH
SWnwaI6bx0dCyqvS9AfwXfdWFLCY1P6SCyNdKbiraZXSkplMhyRtdxMsDUDo4VVbhfpAgHEvSbz6
wl4wflhIgtgUwfg2yD7rrYR1GFIiOyEar4mguOd4Pt2ySBhiC2HbatT0QPy3wxDbAfrYCiFMEvEO
MQ16cATLnjy9QmSQfChPIRQ4xSc0/Dc5gAdaxjDAZCdAtfGXEao8J6wkcDkltfONHDFumfo5awwZ
UFXJeToJStrqqntqg9Lg+An7a0xDC5/irWYjMqTt6+ivQriA0c0d6mpOBaqausfMgu6U0abVD1U+
dRAL2zKOXe5BzqU1A5eoXCN7XKaGZGsZGjv0dXMEQDoUw+1HGBGzFmusH0jp+xDDQ/TSF6ToirN/
k5JA31zvOLVUAIF1IjqVqM4wK4MNuZ46REOtgNO5fp5BCYUfJ7FQm0b3AdZnv1yJJGLrn16QD/uo
NW8RCDLNAeqQHgBUZ1IsntSupesYQ4z4PtGb4W4t7tIvUAFoRlIfbry3TVAfoYriHrkX+rpEe96F
6cckQbxfZDtRre7mpRsCD1B6enMBRUUSWl0GyLErTHNcyMXcCyyR8VEsg1nN32TsUQLUB/G9azEv
sWB5p4OcDkaFdUaP5V7uLnZdxw3PJf0AKoGT1kz9sZViWCNisl42vt5ngIKlsuMnFLIsDAWQ5Doo
pQqxL882zmzyYcqUT+usWhmgZlIDRdyAB6jqQdwjgI4WAi128eXheuFqW1HjdMKE/TM+1DjfHsET
NvmO8eyDlT/EqhkzatNQI9XIKjLM0mp6fvmXbCCKFkinHMYB3EUMJ1WObefx5VMyB61VPG5jXs7J
Psr0VnZvDzdFfxPtjSryCvMCHvCJ/I6Ku2nt1jBms02mdn+aObZKQs5WhsC4gDFFdn5QFJ58zWOm
p9sqfjPxcqWZcoMfVjG1BCFyiSYHHmRiEwdlUb44uldtjntxEZnEwE2pvUK6KGHZE6HyOk5MFJWe
2GGijdFOkQiCqld9cXdnEvJTnjDsBSdISfqKbpWZsNjSYHmaxRspfkTyr2mSBE7r3Q/f5AVnULF1
/ZVcymUXr9ozvHk02Qk8FISg0+SJeZTQ6NKLa/xkn0pfUk76iBwJdtUnul219rYzoUWqSXgid8qb
IeabBQ6fwMqdV48Ol6ngfyVUS2imBxE9WzvW6EYK2XtWbEYmdpQivKzuVZ6gLfHdbfHZNhcLQDWt
UwDtjdTZRIW0HtyhRQB50UWNhUtEbJ7uGjBdGg5A1Gn25DFwj1DrdR1IlmPnnm00YWK4DnJS9heC
4AtI5FqNpDlJh0n0wWS6x9Cxc5IG6NNX0FG0PjAcFP+JKy23O1/+d4UDfJRzwpeejqZrziVI/jPR
a2jkfH7VBivdmGvRqVgF31Twf0gwos9MlPzu5fyXU9hgXVrPt1bVZhAEsEDhYNAioTEUTAW42o42
OilewfxoEVZ02pi6R4mctUoFComL/LbiokkNfCyc1T0bzxCHpUQQsts4OaHlje25tndbodn/bEEV
EiDbLPVfmae46Vru/8VdolhYLb7dG7Wtb7CI4h2SlNHupjnCsFAGRWNUMkf8snCK1I1YbXVgyhNc
I+SGnvqTuOYqytxxnmddeDpbhe4pk4uPML+JrNy+YiF3HNWWutE3BGCdmpN3Ei8ocEq98MgP0Gti
FNMfnnRI7Yp1tmq6OPX+xB/nzy37645ieFWs0uUsr8Rn6OUZYRcNh0ixXoETDIYlNq3WfJLjlTQL
kw57FE70mGJM5x/gcHzIdJqhkbr3VJbTX/2nSI3aefxWtgxuCuGNJQCaRY6IDwkLAfshpb3Y5op6
5vDoFg8oPs4m5FOO8yt2BCV9utEM010ZkOrXTI1IpR0SGqA9E4khqQk6auSrDP/d9aY6K54xr/0t
mZfDr9UDv01OGnaXtIGE9QpCJU1Rz/5T0jB9Myj78FX2PUdOmkQiYgTumqfhl07ErDwh8UIci/fx
sUmyp5sCx/uQFa8qqRrpYh8p/G8RehaU+XgbPm64Anu4QIVE+7tMfaE2MoMcWeZuQUapOcM2pIiX
wBxNsh+N7pmPtVii1fLqeECLZPBzvTZlID7DuLHjEoSk3T75s/priAMMd+W34IzZEMfwWf30LasH
ahslkjXiB4+jZuG8i9jHL08yABnlDP2k/EArB/sTtieI6tzzK93S5uEZb+MBTf568BkVUaYs4RLv
00qqfFdVe2GTU4GKvG8sofqHvJTB0uEpyWgveam34Op4N6Uo3uQ2gCIDq3lejycAfGNd9KPG93AJ
xHhr9Y9uYpD2QcQg3jRpGmEv+xkjPks8U6y+RjORktmqBxSLp3LfWOwOKtfgs6+t5zrvUktXl7Aw
EQaAgcxrUyOMQ4O0LXcCNZin7uy4EV6YgtK8WnXF4imwCrNp0BwEbPXY2uo2E6FVSMoVuaRxff4V
cCi+/WkdO2lPONnBJQ6eF4BA6G5kIRH0V9bsf3+Z9+WjE5p3tqvG1e6Qfi/Tmk3AY+C4S88WvRzX
dbofWhScNoka5ReMwgLQjwLWoJYyGgY9PuprPrEoZOx9DdJ1gt6+xOzYIRBuAPmUdO2sWDJnRZhG
y0bWZChMUL+reA7ttC8h/IXn1p4n8/zPhQJbdjsu83KENRgOtDG3IT5viX5W1Tsj4ky9MOlfFSAa
UeLpGw9Q03Sy8dWsFRpDLa/9LfvJpAZId/ueHwUdLWt4viLmITwYIY60LDk4rijQlrOttxgSsL4w
E7ihKCV8nFG6Pr01tLcgS8kFoToT/aGzN2i08+oH6wFdOfI2rRI22+YG9Gz7eBWVA36sX38Y2sVk
/zYSsQRF/lZbdoYHFupWY8q31KQrXZL5ulSfAdK8n1H+rl2NQ3efdCwSxIaKyEv8czZcD6uxDVH0
7enNA6uGXcGT55WfdsBm0hmq6aKChgFvSmeNKJBVdnD+aaykP11CoGnJsG1JyM71sR0/hP60n07P
OdIjqiPBYbWR9wf+5DeTsj+ZzOQ2OQnaIAMueFE4uJdFUEOlroFU79ez0w7vDkkYWSdPX5h9NmAw
2oegCESqJPUDByfu/JnNPGCXvQSTfsaPQxAt2PhqqZfewPPlaEJpJM0hUGRJ5R9cLxQeVZ3udySF
s728b181K7vE+PPHMx9BSkaCeywq6ixED7dOZ2RQtZ1SZIkoTl8mS1voBSvEtPL8d7hBovqF9K/8
8rtl9mrqMzKWxd3bCnfZkTVgAYCabEgLOMtQ09qn36OMbXN4V4J8WHgTZbw20POINjQCLqwVgXVI
mA//Hxa+G9FzlRizZIj+/r9pkegaORW1/okgvXtOhqGAlJ4orHiUDQ7sv/e928PoIZzKLHRm8U4U
MEYsWxz6zI0J/tnBLQpuKW3rVSSft1lkDBvOXNOAf61DCahUmOOEb46uDH4YE6qcx3zqDqEJvP4S
C46RPDiFVnCHhYgPkgLG+tks3ddcKhIgyxSrycv0BOpqqzBBoXf+u6gTr/bk8GyRgzBjqNwPV//r
LIYZDAkQ7EL3AV/EERcOEy3MvdVJauekyj7mwVCvDh8TeHeCdaXoE5tVKELmkt9p161kQjt6g5/2
ZRwd8yKZKS2m1yo3R+dBRvpdfLom5oUfngcDgwIxSX9rw0p3QjUAjsKrWTjcCHAGaLqkV7HnRycs
8aKXQnEYV4KybQn2nt07a4oSOV+k7oO7uXOBEwuZL+JuFjriglO68s9r60F0dErzPrAKr1Zhcgvr
Zhz9a9zJSW0DsTtMpVtUS18E4ykeeLexyjMmwlxQp40cfbgIsUTBCi4Tdd+XNkGEQNwK1r+nEGat
9wC4qNEl2PQUC8akIrytD2QMDtsOKO0+JcT+3Y7ieeokx/ptmA3LV44PJkORmZWu9R/T5x1Xp0pU
72YoNOEZIcBvDi4fWBB+a81Cd1RdpfaNvq+l1jQqq1JiwQALiBWFA4cZSvmJkrkywdn8uZS2dp4A
Nkk3Ugjylcz+anmadZ7c/YP7NtsM2UA6qma0MHJ2cIZL4cvvqwHHZYb9zRGxO9IlcigStiapBACV
lkWLvl1nNZ9tUxqGb/VPkAy+htw9BqWO6N/NXmcMwnJOiERI7FrotwiDupbCuFWjtCxwhzg1YuKf
NQDhUuwszsekpOKjXgFa9FGd5U29RWtsoW3rKC6BUbtyPlBXD84DT9pS5VuHHTQA7VjUTP0SWT/P
eb65SHatPVtfj9DDb0htT463KdGJfr8Z/QM7foOb5pjZjqt6fgSB/UMA3vE34akIR/QbY1hN0Rq0
js64H1a8SfrRjZmT7ddJlVbNpq+WkQp54+J2WrB8TY5QXv/eHxGialhXJByX+YaloXd99pZ7zs+2
D6qz/eWV0ShehB/DYsm5S4NDygdTWwl0KovG1DhgH5UX5goHVjkOyzO/DyhtWj1dLiOHiKzkIswO
VEQvDXdKIhwP5MgvWnCzfYACL0h9baYQcmUd8ABx38oN4PMrUqCcmE+ngh5ObIIr/1/kDaO+sJZz
kBTlfU/R+PiukwxRP/O3koDehC0ZwUPMOMX5dq+SqP/1aJaCcfVvHmShv8c/p2AQugO6ogYkhM9G
0OFWqvaSznoKB6ufqkWCWpjQolb371kQgvGZypR59hwTVbO7Zfz0O/DjJy+8VdfiyrX25Y/zpYFI
NhwSz0fdHhEospckKv09Po4dJUJAUuLaSXvcMu1CysxySnEby6izt18VGaZNnK9U2IsfKpfVVMKX
PmArSnq8dZoyS0C7apSTqwxb8m6TQq58hsCXa5tOuYPTnTc5i0nibWXAFW/dAqakjv/CiXH/ebp1
uJo1iXUbsgS9eLKgSKaYbgG4cW0WPsbiIoKjotmIrQP5A6JxLgmrDeyu0PdNm4o9cmSSVh0fbyho
Jo/psvram53J0WNx4ZUbiQLgg85sjNI9AqFCp0VwBbipfwDITPVS3Fs4lbO3ENTsPojtIga7ZMGZ
peGviwwPNKP8P88r3xHZKUPHO9Ot73EVHc20bvwIkS8oBSP6zPOqZvCtMMMumm2CznAkrvO6PkC+
Q9dUBV1b713X75dqX/3IO+gbF4Aopm4nXGkb5J5wh6cjJOtHjTLxJdfWn2sMlg/8jJbRCEPJ7Y9A
JRUYhN6bVOPnGn0nx+Kjfj4CDiU/3jm1w+EIbGF4/D0UuDO+0hxw32KMMM6/8SfpypSeYWHR58bO
ko62DiQXFcolA9BQW39A02XM0DnUg/SJNbIkgrC1e/anmmEa2HY3jS9sNSnWVOqF/WXDL/OKJkdU
jNUw/qJ4WpgcWqG1/R4tCMWYRdn/PUL+qXdUgspUFF0z8iRw2sC6WUwa7r3RtOvjYN6aL+4yHkyx
MGeC5ZwmZ5pMOZUlYQnSGyli3CV7r85s8rQx73FiSZTklkogTjiJqGdOf1odfZWifmXHUO68js5K
Y9rboZc2iPsgLwXgXm4eVefWqWVqc5mjYGbP5ijfBpDXfdAslBVTkzltQ2O7jZ/pigpxmNd0wBuY
NNNXe2D+wAm/Ey0JiTx7Uu+NaRMFq1gVGUHrdbbnnBq9ZYDCCKPulPPppX+xMHDEMP2WV7/pXJQ+
KYlGpHMIHxUSR0JFCv7aZpRz5ODEbfYHhKpmTeapHzQilPT9gn+7mqMPHb3PkSxGYpr9wUJtiF9V
pQ6OUSzOSR/KgcVYR17wc7bqrCBnHdKK0rWRl+oirbR+zCTF2ZHAJxKn0HrOLLYW5YPMDfknZKhl
lqwYNXkwpDVFK+ugmyU7/AWl3dTs3c4i2cT+2F9Pn8/WANTfL9hBp7BpgzQfsxCt7QQdQc+HZF4e
HWViQo27/QmZp/VVuJnppwFCDdisylaZ3I5G2+hPxktgJe1tNVrPJ+Cj6HEt/19istXSZACKmvl2
ROGIFcuMdj7/J19OJ9YeP4B6aRYT+RMSE/ihDGGhexufMwtwBFvlMJf/AwuYttndhoz/j21VwRMT
4H8l/AWNe3+CAavckdAzPy+1dl7nDMB1HWiGdHbEPmvsP4CmSUjzCxDpCcXoZmP22grfoxroAZb/
5X95eg+Zzg0HyPjcakto/I2WyrFd439kWqK6I1F4DdLyNkr1gONd8rDCUwExOd5Sb4UU4xiQUBtq
X4Cb8esEX9IzfFSh1oNFId4J/yED/qMyRf+6+axmZwSX0cUra7nh3QAAF97ku6V2DzoEf2sS6qcY
1XXa+ycGE0nwHlIh6t/N1NsDsIdk3fXPP2hd2jpXjg8wM0erqAWE76A2CEixC/o+gpDsvhyrH2Ui
rVA/8/z0v8DYBr0bZGK0/cA7TxaBoxzyLIlLDlMbJZowJT30oEttRl3k7JLJPfeoTxl3c8dTiXRI
EaeLDlZNnjo3BoFfYnsHiGyRwxozHEiiFWunFS4azEoxtCkgyURU8Na+EJZYKZIxK9nltXaIawvc
QDFAU8TPc7YkCBFpcA/qRhi6ATXhtpBlKRi2g0HRu3GmtGJ64SOIpErpe+wxjDZpAXr2i/THJiTg
c/voIwbomh0sDmrNZD2aKXn/JCSDt7pIfVolPMZZcSg8krqR8bqRvRKBIuYYiVc8HpA5Nxwnb5ER
OYIdZFR13UQG7ym4OvF1DApMco3dff/hby0et1MIzc2t825dlNY/xcYGpBXRMqoHdJwLj9efdAPK
B/MhlWcX5oveRr7cgeu/WQkRx21VUtyM4BHAmRQIv5gzl7oOJ7mSQ42TVa+o6/HRtIZo7mHaPtSX
CDloEau+YR/7CdD/4ItSPxYBXgMEe1VwKSyErtvmHZpmph3KYuvwGOkz5iX765LwpYEImfuUKu+l
QPp+PD28587hUPwL5sDxNp0m12jgzter+4OW6RXBUA4v7tXIh/AVHxDGKbQ5rZZCsKrk5TcqTtju
SDrZKGt7mSwD1AmDXzeWCw3TcnNNPxJd9un4MUgyyqPlx3BWIQX/oTxdckev0IqI26NZKNEmWquj
uePnp2YTZqqA8K2M9JOUMd+jVs1EftGgahqdgQQ6L31CswKivms5Z3WzEkR978nE0Vk0qloE3Ebm
eKupq3j5DohozcqU8j18w8pXAf0fKiZfWJgRDUCUAHY3uURWxiO0fn4QK0DOGTIO8iabL0DsFicE
xGgt3V+1vN3Bpyya1ME+Iybtfczigl1+qhvD/thBuQM+qLChP8ll5zUPoFUjAGjLr6xvtuk/sagc
BAs11F/FC4C3dW5aWKaPughPjjZH51dy5j3SsoiBp78snPg5FTixY+t9Tg6t6SbX4E+mBPVDPsIG
qigZAZW+CZ55AySJ2tfw6l1nI94HUj4z4BMEpWVmk3oXiRy+SHktVVCX0pAV9ij/EJDsrcne7IMP
Yem9DpA0ioar1SQ8bJ8G01+7jBjNKeyhMN2oidtyWgP/cmTTCccIuZq572KJLg9tWtj/xKI34RlK
arkFEP9JR7z90MrdzIyuJ2yh0QhE2/j+clDrUMhWwICgkKDYC/C2tXexO6fOOh77zvtn6ndk1cWW
lsi8ZZGVWs30zwWhVvwD7NmfLOxewe8U3HjQfnNgaHvOUjpA+5LmD62Mqfz0ClK3p1dM8ByyjUlM
9bHq97PYP8INYt8ueblY0KZyV4bKghxuxDVWy6wwIELmjNz/aefg5UdXQGkIdcT8f5cDtVh+zfzX
7QbVWgeaoyhfc3v/goBRm53WCBdA4ejIYCETTN8de9edB0gwKvlC021T7KAVEA7u5kFPtljl/XIs
j82qTEt3++zu97wI8/HD4ldaCNcDQe+YxI9HMxHpi0ET75ZcWs69lYtI3wqkpmF5I8kDGvObLYtg
GfsbB5b5FXX60IziMo1tRprEuwQL1NsZHhog278MhXDJM3E9/VwqLfg22C2oDP/3NscpS1i8TE+O
rK8YA9oEbcx/reNuZL1sQ10RtzWqey7J4Mj23YRYySMHhOIiaq6Sf4jXVikWY182kDijhxRYMtcv
jaqnn0kPLivEICqzAbJ4CZryC9GECL+YZnTSCX894MsOHmvrryAw3MPpqAk0h4vZlFuFfpLLHynh
R18n/aTwNHHXmgOTdhR08touOHYw4IP9/w9ohBh2MxKScqk8+eV5aB20kT/HwXzy/5OP1EyFSm/a
QZqNvX0aYJVTuxQPPzYszuD1IC/eCWeNE/V+Bf3XXSiYGdUdqWJqqrKOVrE1bmrTz2bBPu+MHCjY
ng0gwBu4qx8x+KLi1unlJnRatWNDNU3qeVyH/3yaxhLrZBGnUXtIcHFRIUc4ckWCbyq3CaPBgxYF
kvVOk7/9x55AFLanvweorHXKbrLXWW91Cles7TrcQFxh4Ivsn27OlOKAkuw4JNX6yru9wrH0ONIt
E326hFHlQfyiqAYQ0c8Ls2wtPu6NYzaJJrxa/jZ3okOTusRG7E4AwmQsXm8WTbEZddGyAIg9VKgN
XA1hO41elX7bZ4a3KFVj/SfGyyjW+HAfzkQOsjHNYoacOOfINZWFWG9EF9rkNJ29jDpj8XQN++3d
PJG5MzOddnW+/16ka0E1ZN/7n8GHTyndI/yQuNyAhOxeSp+GM24TDIe59nWjcN/x43WKVwq8z0fg
lcbiCgJLpwujqtPMclicmYI7PdGdRf4txa1zO1fLj/1kc87n90I65Epg4WEt/F2e66Zk7jJT4pZx
ZOs6FpBuBFwiIyoDgj2yVjXXLK9fGw9duE2njCOyBmtWZ9dQCn9ZZIFz+MjJw1hdimO2ysqoceGg
u6YTOPJhA8Ot+8q92wGR9in5ZXl2GUhPngUFtTd1LN53MGFF3qSQiBL01i7IHdmbvDPJBwtCv7Ps
yyHHaVDQ7yez8/JtHB6F6IE86jO7JBIU5Dv+1kp+9GjHpVQUXsz11yvvjlH1zt3Aqtny+ZNMF4LC
0cl5Teap7bpTka93W8qmdiTYv/f2bl95LVQ+osngj7AEWjdnrsiCx+ipaPmdtsyll9OS8M9ttQ6P
75FXFyzlCHG1rsBB5dUB+KDdxJtGiDMrLvQoiaywki0y300j2hR8O82QxlYqqUDT1DDNdYrGcxLT
eqVGUuzH/fQV4xu8Lt7n6A3m/jtCw5SLLZ8b5P3y+9tg90UQy921xA7sF3oDYB+hKEb9XlcsOYPP
OlOm9uenFK62WRfyERi2uoHryp1tRxbtULC2fjffkwLtR4QrkLgF8q3d8RWZblue9uMJyqFfAE3r
/qBaqIZ2+KDfYpOuJ4ycXIYEQws/qYkfNZEZNmqrb4fznbxBWCirqhIbzMAZ+Uv7ZsGq3xj2hmUW
zaWOHPhauUknVEvrkJ3XtXT4IXh4NTjlWp0vGSje6tw7CYZ8Q+YIsQ3IqhNuCzWZyLLz8xXc8Rqd
13cC1L1dva+28MZGD5D0qtMVRinvLognxQyMnGuNCdW6J7oArj6uNPlBpxbKE2fmHwj9GafSaiNb
nhg1DGw2tGM9/FyF6BB84qvZ7uJWstF1ypRqoC47Ul+iYmTiaXHMsrG6ggZioWKi/vvMcvOZFQOw
Kg4mv4ztATNh1OlUZNJOEuImf/oKJQjGz8pwpicKP8CTHGn/hCi2W4EEJwHwV4+J7o7jXID84IvB
Uu3cmIP+igW47+rQYJSJd2fEDpEN9BPClvmxkJrE7dwnl7ZCJ3AkbQI4WcycrYCKKMynYKGs/zeY
FumAIngp5L4w/Wa7OJ639J7322fY0UFJVQQaK3UbNv5d6VLcyKJPAJYf/M2XkgFgM5VU6muUJHYb
2hyTOz7kPjjplfwRABgQFevEZGpC+X7qbi091P9TxN//NgHDwIrh7Prj9vbyx09VOzI2NRDcXzL2
Z6x0J78Wq+ySB1JQKSE4eMQcBKzIUqQljFX0MqELXX3hlm6nnSzkJYwhyCjX4FVEUsC2zGypcDzT
cOB5fHvyQ/qLqZgtChNYnRm5+1XC2VfKGoxHAJ/v1mrEDP3APjb0dzVHLNT8vAG6ZAcipwak7J5U
0ipZNuJbUNgK4RX9gxyDdoKNhcVNRn7QdGFGITpEH+li//5Wfe4vpXs6uZracA2tRAFvHx64aGTU
wFZbz25jOLqcrMpovAqI5NcstXqkdYREcze/U3KMz5JZeEp9ofaBdVkNgjtZRoI6tE4wFSMBMhok
T0fuAgVbBTvkbaGrL3CaDEqatgRIk7Ki+YhgITUBHG8hoRnnxwbWg3roKuYU0jJJbz4IstMdbYYU
1PnA2QHoAthbqG3pdCUIa4C/Ubhn1Am+QkmmVmHVTlBVZ4njvAciJrXz4/raB0RQRq7c7MVqXa7l
kddehDuMZiisZhBHhoYmfeXN4CWJxfko8/xKkrRsjbs5TDgjbzcFJPkiAqoBNrzrkRpExjJdbPA0
D8LzFplpLafH4zfg0hWG64XRrgFimXvsS/tKJvKIE3Th1YxUJK89hP17MQS5lsEhg3buUIk8DGAk
apFHi0SPmvzksDED0Ro+PV9Fj7PQDeCx1T6B74wTmR/cF/aOzOUY5zaxvKecfsRPgCj8A+smhzvV
Hp8Ap8Vu10Ep6o9wuXBeT0OmXkpEPRjYdwS37z/OX1u7GpmJOySIeb9ewUjPi292Qf6bQdVOWlbX
3yJl1wkzWPy7KDvx7A5Ohzeh9kVBL9Jr/r+d987v0biRRlRI7XqQumTBrQ/YSA/H1k5pinNbaGbo
iDN2THrzLCAGjEBEM8R3qSpmO7H2lPrD0MRYFXhYLC+rT5zFcxaJcxGNfYXOb3KFOF4UmP2hvJGd
1dbPJXZtBSlzoDi74XfZ7UJFZtmSdiNKgsrNhJw8bSllWgHtlSCZddb6mz5MGE7Mw2xdEJ4ZhTLx
bQm/crfL8lay5XJSujSQzier7kOP/KA0ny1Xwia91jFMsSqI0ji6afeWCtUWCxNrUxqH9+RMFwad
/fT9Z9FzzhQBpWqmrQ69UD7bfktrz2Autha3+43/Cdf+fhkmATH+j5D9DYw3cjbwCQ2dKjPiwt+T
rbg0i5kfWE1ue1VvXMnBTZnWiLXNghH+UYYdf0nTKK67xROGe9xj4ZgVC0lJgzNY8z5W6bWMftZb
lUEzWMxhoq1OL60KD/dUojbFpt38+C9Yf14ijznXZlPDB/RiZVFsH10tQxtUFtjnXKzF+8qZ0e17
A9wh2yOXgnVULfeOYVvNn82Uq0Bg8VKYDZteIn6sswPJxlLIUPLtImGFkO4t/DybStizWS1Oh3l6
NiUDsvGzX/v00R3flu+MQzab1LtLPDaioPIHVDLYztsa1IW/jGHNV/5F2bTC0fKL0Q/LvQo1ZfzK
EklANnevbIqJhRt+GQr3Vow0P+rPd6u+A4kAJSvdJ3VWP0jBD/ppbsAZGuzTiBhDw0kLbcxo6Dxe
iEiCbFgDda/D4RAknluqL+G2YED+wWesZE6WzV7Mtie5JVJtw183MBBZXFXDliJSQMvWZizVc5mb
zMTIcxlXWQ3SbXt+AaaBi9nhROxCahbIbOgEj2u+EXgRxfuPr5K3tyFPck5eeLL+AGcFcRyLJyKb
UXSK0CCEaBvU7p5gLmCnM+DgYeI2XrdHAFqzeKN8C+TjUdc5MDR5kWOhRh0CggIPWInYMpUA6a2L
LpRaZufMfCHpaMPZwZdRp8q3F6lDWOwKObentsgYE/p0zWu1k3efcXU3wM1Yl97q5U7d0SL7uvkR
zfne1aQwTekW2SC6jfO1QHgLYWv8sILREuFF9II/5kbRXk/cqWrBWqlaJ5/hX2J/H4la3M0pVIGh
d1DujskyRqW5UiNE0VE9+0U8Q6JWhc5+gqzK90BUn/XW5i6LxSCWdGgQBYiVerWRKC+Ohv8Itmgd
I6flT9THqb/WLerrY1QBVU+NNolbDjk28ZSLcPro6YKwXfABQgiN0m+w9LIqBFa6Yp4x8vRRKJlf
sjGGDE65/GVeO1fHobT8nbDUVpi6fWpLFOVLhaRfRe5mvS+OM7do65515ZwzldswUctMDT6KJPQv
KyfTxVM4eDjVqxttS8e/0DbrILKBFaxvXfRJUhzmYjA6oSJzSfzrFH2VbFbFlD/nhwZkiubQWVNO
aAo8AxvgUDOFBUWgE/YUMBeBB02EJkmeR8FwKm7GK1fYVV7U5pSnfqEUb2sUQJ/fiQnxF/TdzBM3
3BIQBBAIhJvUaD5dP5tqmUjcE4WbKDHvHVeYIiU7TaBPuJ3vjvGXPLVFufyI6htatVOf2E/RRkKx
Ny6H7fJDZmHjbf3Cn6Jp+Byr7SuJ1lxaq34hyP0ge6dlqsXALEYl3SscGZ6G+uIlCZOaBCmLUlSm
yosV/+0bMJOMpnePSJB7965/Hozc2jlAS0QFRpjdYIUR6XaDt1BczutEtvV7/IhpdB7D/xjj/2rF
0h3TKBELqUsvqSLKoUtYPNFX8LWQg/EXaY3g434gDIJ8yN+ni0rqr7/f/U1pxhm6DHeEektHN0JN
xwldwK3w7HyFj1cBQ2O/fTxXSfqpjXV0GBs6gpTcx+AfrrtTc4CmX7se8sjZ5vYNf+QXrrY7qRSN
Dd+WarGgDMSgzdfMARlQvM3DelV88EyFhWp4i9SwDW59CKlX4//OZE+8Ux+8CCGZuZcJPpWjToFU
o9493CBQDefqxny1+Ow616Ki149hPzuLhvaMgWq5N+lyuyq6q6ffntyMSs2bD0t2mLiegx90dsxT
MoovwIRLeiaEeQIz842MxY04SBkfMkV0DMZdUXMbmLISRIVZVkfHtgrHVBBvnfwJ97teIkdokcvi
HHvbTTvls/DhL5DBlawa9Uh+5vr/F44pPcKy0fbZnoJ0lgrsxnwX+8FlyMwASdwegw9KjvqowIQM
vxshPU0NT28FfSSo23uxcl+R3FYUzHTXH3nuRv2vH/uhPoAh1/1zu1QXtNH46v3KNgbUEYyormtq
aZ8P6GtcBilkez3BjOlMy20drHi1RFqGqI2Hu3Ym880XWvTzeGaH9vfPLe0QAwHdxDZg03LI1I1O
xdTSLipvGfeKgmsnDnzgAdPEHOaQ/eg2G6+XZATk4qYxHPvQTguH8zmOX7m15yqH7YtGDHoqGFbW
N9Yd91dTQ0kzC9TfL2TYFZLV2QzJ6GtgLW1vVz/jrZpGc1bQNsOh2PpCN1M05808OxlXTKk1uoPa
uceXUoGKl7RB38dV7E+MjegcW7IvDAeCVx34+IG0N0aEyqQoryLFw/IFh7RETW0MU2s4/HaSYgqZ
2vLLDQtfCIevEzUZR+tNlVaJglODJPWazSKZSyif0SANlObtndov/FJC2RFm+txK33U7rAfiRMfu
MYbwN5v2vo9t3KtE0KRcWMq96lZ6TruBExG56BCVPcNPQJmPufe8HS86EcsvHDez7iZ9+2MEf2gt
K7I6qovyzRVO0EZ9UGEYGwSSlFFFVk61t8kyX2W7mfRICgSTvO7svxmoC8zrYMVXWEGJP/i1oI+k
uodPVNDOJEzUlTYoWlKx5xz87UqnnRgC/5E8oPwYolumia1cdAZd0IdBly2LBXfgIuyJVgBpbCNI
flz2vwZ4CoEnJBALj0VHABRdu5IlzBs0DdNHZyGoFDfjfWGEv5kWlZVvEqLngV2VFUtoeRyogEdm
z0YdnJkH6emxOFR3yUmz3SnMsQEl184zbbmgbYUdmTWY+Y+HXQ/687neSdqEVc53DIlTttU8lq8V
Ldk1NGJOQN9JMT7coEQVjTkKphEy6AC9v3gNDFALH3qZ876bdtW0FBFfecGAxnzSIXLIwgqX3tCJ
MYJYYa1wGBd0z0Qoq3wXLdGydCge1IOqMcHuazlM1fyPe+vFQ9v2PSKBRHELlx8ne/W0h7vOfoCp
f5gnL63SDVZc2+Y+kDpuGt3sJjSRq905YVeC8ogMap4mfJbdM/kPWDu/cnxeTW9zLNIgHonVfx95
KC8Vc/adFv/shw7o9zcrzeDaq6bEYjiC/svWNLni7cV0g1hTr+OrAnFH1s/J/rfNRsB09SEr98uY
yFe9Rugb/xpVC/eKcKxMJVNOzD0v3TECnSFeFwupGVlEHgXA+8XHkXUm7aKZ0QistESj8i6FlNGA
1RvPPH3YwdVLBnumsZsJyrq9/rQvdtV9/Zj4tDC5unsysTpuzjhALx4qon7FOhhe6tz2AYwbovcj
sG8p/5DdvV705SRTI4vK4UiEArxDIw/Yvcb3IeRYalpKeGf/RokuxaRnDAx1WGLX5qmkdn1n4WHZ
PI5hjujo4lxpKN1OTB6pbAeGK8/O+uxDEmDnrxJQZ5Cn3EcWRsTUblYjCoj5LjSE2mpxiSLITdG8
dBMixki0sMRx58cnSWAMpujsqjwsEqNS0o4sOo7kKL0z55C+1Q3YhEmY3qYT46T4uq4fwZRim/ot
RLA6z2IAeBP+KxT47YDtXFdaBWt6a0KXtcDvpVvB05pFG5ylr0aLNIV3uZC3a3T8F3pEMKG5iEj+
ijtzZnrIJiKZ1PCL70Om9KQ+tZV4TBWix+Y/HANDFsmhAV5MGsMGNP/5loq81qgppBBdfpCx4zuR
uBpaBA7tiy1bvSD4R5MabCYp3922+xsE8+ceDtQrJUVvWIEPjmUMVBZtiBvuVDox/fZZqj4VW17r
qChfeyVlJTZiQfUQlRhBGos9EG3gImJqZqH2meMFzB3H5Ms/NjOGY1Ih9aTECwLq65hiYjNHMheP
hYUbv9wvX9cVDi9DbGI1lbiuPR5t9HeMl0ciixzgA3i9gD9vmeKzExzs/6voe+gq6yN31/8ExiSm
MeUelTf/KHS5KrMhwoCCTStPT35xyO8D/5CNMqZmcNzgGE0oyQ02xWSP3xzaM0ZRNRChd+Y6/F8d
dL6HGfgXWQXFHL8g4qn0qucqafgYZ51ckmZtNzZZzm914mSb7Aeg7fpUozBBZqdgpcdxDaequPwG
FZSDmJF4Rb51SWkbo/+epUXsTs3+A0DePhXIbSvc0ZMFqYUTTLfwBmdEbSKj8FIh
`protect end_protected

