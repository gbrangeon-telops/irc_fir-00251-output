

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rMj+x3ocDbJ+0HvlMPtFLLYN4V3iOWmu0i3VYcvwPU8r9dUqilqv5BoOperD1z/j12cu4ait0bNC
TvgieQY6qg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LiFkBwHJvbvIRsrs7TuS9x+hbpgzWqPRKAN+86jD7W/DWOy2HiTI+Pr3kejl0F7PQ/wd2Tf3u0hB
l5PFI7Uciy5uXiQA7fDmYLdPcNoMNQWm9hohp6Q8wB4H3kSwMFgjlrwYcv97jBF9K/DD+f6kjMEJ
pjxxREwM6oJfyPhyhBI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mlNr/JQ7BAznEw9Lq2hOb9T0FUxDG5TxOJH6VJoPGS12EjdrVMK5Jwy/CrH7dSOtWY2eUHhpsxFO
HZJnPHkoY6pnOp56kFqNAyiHJP+z5BexlWOYCHMzTTDXl5ecpknkEs/jFqX2DjV6R1MuxPdeXOjM
JpDfpA+rd8xFCgAvhOcvKEKjw2lJmNukB/NqmGdLZU9Yd/iDC6mJcVuTrR2gzFDMoFjQUitH7TCG
r1krtYbVQjkm691WyHmxufh/qSc3KdzrpZqycBevqxjmEqCq0nMXCiMyQRHMFNk9XLymhnx09LIk
8Ck9EeU7sTUKIMhZ7oB9NRbr0Jmue7w3V7zoXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jcrZIuGwyVPSe4eEqA3CjxEN8wKBf64m71qLvmqrllZ8mLFeyFjj3f796U4fol5LeUOSCUITklpk
5B0LZiT34IugfACCFG6eSa/KnYkpqdaiyFEJag2zBthAbQTJIoKzv4hrVDSwoJffRhWS6ZAZmMOH
9HJ1Z4KODhrBj2PMMOQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
He/hsXsp9htM4v1ezeHFxTi8NbCInK4GRCTZh00v46syUmSwf+mXhIjhLm4sHKCSUqmWt1TLUp0m
CWcpoGxiawBF6wEpl5GgUNyVTq+T/CrlV9Oykyiw8ESh1/7hqCFXSES7D6yS14KOyEm1cr2UmC+u
X/NTzDDvOd9e5R6zaiks/z3Qdqxiq6f6jnMuQiSiMBsAMCHxpq5kEezVTATURKXvDebBjGkSTomU
Wve9JRKQPSiMHuUURnaiqzi8t62PeJzIwk64jI0DQYpuyHeGDNIZt8qQokGYPimAYp9IilmsSuGG
FM6CnM5XioVenoNWDUkk1F8M0K5I/5eHgYEnkw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30400)
`protect data_block
THnI6V1UqYa1ePEXxtbd93Kf0ihOvvoTduiKDm+p6tJcoWj5VXoaGFrFV/PuPjFmArDsBGAABLBI
H7ybt/SrQhCn4B1PgdhEnkOjG3sjkWX7EKTeKlq+LOYbCko6kIXzyAMvc8UFxuUMlUIK6C6PqkRY
RplrwjO4ybUEnoyY9zq1K/5MQnw2//Ket1Kl7gdlMnlQQUOszmABXRrG/OobHVnOkW8bFuDefgb7
AHA+1wV7CJMOdB3ZirJqtplX+PEdDq0AcR0yIfdBVIbQ7+QVJQEy+VD1tyvdefqjjJh60fSdiVJn
GSuJmWOJcFUisb3xqUPIVTuvufubQV/DJe8xV/CYZgGCcyAVskc7xRcUFMj2bSXwRi4MVlLtucMn
s3GCCMI1l51eBdBJ+hiuY7MMrASR0Xo4A2PtZ16bB1aNdcf/jNxyoVLzpef/x20SKw1aMNGZ6H/Y
Sj6Pz4nrfsXd2OaaGZHSkPeJJgq65N4aKrwLVwlg569ueWpSEzKFboYx9z4/jRr3xOJzKdUx4DFF
oxnCKRsRVEUQMZ6dl4dOeclwasPlHh0b391PNZbBLGHnhe7BbtlH3btjvx9ixmGloTYvkJOQqWZ3
0+dTf1MUyucj7tpwomMo74lzJo3BEXAzGUxj1eyvh5Njmn3+IKoHMqYyDX0CL1bKU9H9SXVTA86G
+zV2HFSnlqBn5KGPIwfOLQFYLvkWjbQPDE8j9JmmoeaAyGMe8xpWfYW4jOuTtCRLYATHCMhscnNk
9vyvcPvlgQKJJ+OxduRfIv77E+lTgR3kY0uuyoxLTSsPQrsVFOmhOhwfwQwJ4LeQ6lT2lHyIm5/+
zAyMBqRUy4db3hSL4l2k+vEV/BKCrYoGxxz02sZEmovjTBh1FVYg+QqJx0diyTGBpT/qQ3Yjqnw8
7qOBfwMxSjteVUTFpE9whRA0QFByTzKZIksik+TAkhfCjaEfefRCtw6VoAnhipIwUiIJluGd3srj
NnUU2uWeGRnaLJeDryir5J32+1w5+IOXfVEF0LChuXZcH+J+w0njg1PGz/PHxGXrnb+itPxKUK+d
cowTRjcjW30EqTtCgdOqfVhTgv0od78e53g650B53cRnG5msNwI02G9Y+lWpQBnVZBU+XT7uyaii
kdpRvsu3p1px7zAOZdkC3NjhHOTTaQNK7PJi1UmAryrePnLliGFJRQ+S5JRofy1RRk5Q8Y+ePAtM
t+ixv9y4y11tit+MmSGLlcIUmGe1lTPOvA6iWjOxir8upVJIG1rvrntjYKR3vkCb7T6sBjErvRkz
adKonKKhNHQ2TiJzt9Nv5Pm3BNAkrqoQi5FdJ1+ISV6zdjtDtE0lAEOHYKcihEETz/B3OcmeL040
qBwunE35e2IROUOoGB1EXnARZ6zffIqFVJ1nvtR3b1hx7qMpKeosDyOjOYQRzXna1rdirDxsgKL9
PrkJqhJef4Vmw8+HomE8WXgLvmTKR/nQ9pjab4b6mh4vqVT2ZVjItDtiM78zmru+WeX0AdWJsCeA
HFQrzw89Of41hRoOfmp4CgCvCTOX4b/juFdWOeHaqbPPyN0tCk5Dwb4Xhj/d9+BJXX/7RsHuyu/V
pg3Zb25J6XJy+di+RFqU25U4fH4xBZ/nXMhl0ZQxccz1VXfRzAcHvxxbgkildoPd83ePhTiQIX1/
/LHAjROC1YG7RtsMPDzU1A34QaUi8paTIK/DUx8YQBSels3WCO30gAqauRvyDDS5dWuGJLnMbxDt
znIYpkjleDwkprlJUOMQdFlRNi6HG/21NiwtLw2kUfT9eWko6s4HF8rUNpbw6iTsxKkodkc65XPP
ZDmxRJEBsLVRqcUO6z5pxim0lG60KnSuPK2r57GbLg3mjhuU/EdqPYAuPK4A1mYj+RFFg1keHlB4
NAkY8ZsJFT/Yf6D8f1TNwq9YLfNWpF9WBCj8xCKEtYrhlcb7K4waZryl2AqfvbowoVjRPFP4KnTu
t0V/FJ3y2urB/sDhWIwE6c2uVzgZz533GMKKuvjcG/F13t0ClESZpqiJ4wGEXo7mszUpc6mcCLN1
57w4cxxQgmgCNQvUpwH/+bQA+Xl/2Iz8xEVvTSQxHWQL8yyzCz3wmpliHZbFpaBjBMbsvfVpzgLy
NALJATL11yJJqdSoNtKatvmNXCRzwKVHl4n6dolfeTPmKidaxL/usJhcOcNfiJIR0x3ItpCTmfDA
r6RA4tkZTl49VvPJB5dXWAUfWIE3v+XkFj9x7/Bt9x5ymp4PaP/4qi+DjFQYZS5WW3NYMEWzj1Xb
bX3pkCPtofQCbPk+u8D1IQQCwYUFxn2o0y1YgT2DjfsDltRHedROgqrgcqToMkDke68BefRLIHUP
HV26FZSQwHCF4ktCSFYHUgEGrjxRX2ioZVslG3QeOuFYJxnlBKYeGWbz3tMoo3wcOPe48aMOVfdo
PW/CXLiXvr2g4QxKnx3DN5wA4F9HNulmH34Fao+6HN5n0olU9WCwPvtS1eShKIItYM0vgDMJ0WnE
gH826SZO42AZxb9qTyHreSXIh0GsCt8U1c3INVxBhaIzuQdJv46tHvVC/r/efohsYdoCcjzlnmSc
xHqVPaF/975pyK6cs9ddp8iZkqvg8kbZhG3N6nln4LwJGAzCvtPgxzowUU61MwqroTq/qvJSvYr4
hAFZrVFQ//ON4KWwOLOzhlO06eDlhfWlsWP0tGSfdlIFsTafwYmHBAJ8UbqhBKsqy5K/bHkIg8hx
PFLSoMgqkTNYWjaUfeTuPiywkTc9iTqiMmn39iRO4Lp8ylSTj2YZQxKyDtRnt9ml1APN2kvtSGRH
zijJQp3uFgM3f6V4dP3UhO9J+s9FjF8M5gW+zU3tn4RrktCH2h1KtMbbP6rdptN0SBy/wWHCeCZ/
LISgPlRKz5zKuD5lpLIYYVxS1/Nf3DBcGdjmlongpHOAUvg2NOzG71svcfSLEE9u9YCThoukBNHQ
MA3wtR8ogAqmNq/i8eZaVNOOZk4RAPHeu8FAil93jmPehCbADC1NP5RoJcEA5mqRsDrnAU8OtF5X
08dV8MLieJ5PH8HEiU6hnnhoGC8i4jz8k9SEsk0dst95WDL23wRwxjuAAYpT35JCKejnGtlGaAxC
2jlnLcmZpRXwXuaBbeuD7nQkdFyBxuLQTQvMCF4AcMqxXeICsVAy18uDYZ+i09CgLR4Qeb2PGf+u
AhRjFSkoY/sRMZeVzpwTPpA+uGcJABjJz9G0NXgPT2BdR8ZVjnTKJG2UxcmDdW7LsfarD73kv1pg
oLOg/ajm6TJjYFj+2yZu/9/R0iLGL/7cjWcbgbzVS9ZcHyJaErvGlXJE1uEL5mIRAIQrHhytM6Rt
8QbFTfIRy97UKIt08weXSyh4txmIoikgr+IL3i8V6jooiTYBAjAWQmPuDxARDxEIXN9xVfxs6tYi
8Bkk2IJ8tnAcGKm6+SE+UTPQn3dKIyycshbSmnkeEcTtAt7qh4upud3oK6UBltxRN/9pk+A3Paio
AGTrZjLLUypHNCV9ONTn30Ni+DTUKtfU1IMLYHGeZNMTqNQkf7bNOA10OmJoKW6Xo8p+BiglqDVF
6u7eEDjgrPC/rkyNhsWh3N2ZF+d+1gKy1rB1W5L4Hzdj2d0a1JDK9Vm8AZvVOZLulaqPaBbnfy9d
K7+71GjolRtkDBRiFxml1pWgn+MeRgc9DnsPC3xdoAWKtuXDra+4Ehi8F0fsY6nBHi05Rs3atEJA
nFn/0TsMdqrff8QlZsG/gXY3w4S457F3NndZ7UakhY40wnYjQJnXhOl9wbw2yaVMkVKELuLNqBuF
a8Vc7AUL3bmOPyO5Rpcu9dQ+ZsER6Yd+IZNYvtsyFcx/YKf8TdqpVqUisb6zTVkO3PFlMahFunHX
lEpIw9OBzruBOq2caS2sqD0t5DOi2FMJSWOqRaznV1oSPHuDnAXouIPExOU4IgTozFjJuiRfQvi0
uBEZZx8SngWHpifH/Y9bfQwFer9/3PPjlkuG7bZZOAAtbg5aMiOhGZwoxmJ6UjiOaP6RniTrjz6L
3gkGvsualVZJkDUwT2Fq7CvDN+zjim+TrPQ5a951PfWYhUKeoD6VFpajjv6B/Gi7iU604qL0r3N3
YAWP8sqfT3oNJFDSqyTt9TLSjEqRJNWaYfqA689rUjZpMANOyJYazFxgxu0XrqO5/+jPLfqcD2CX
6O2MRw9vJGrpWved0YM53iwzU/gav1iTlFsKdsFhpl6UeNnbdYGsI7n3FEKnnOcEaDPpwXigDH9s
4/bfzZtmSihDGDd4kL3KzDyDvWodaBPbk04NH4rxPcrusAk2ZjGx9e2R7/JwPdkqbvLtJ6ktfXJE
cfcKTawYQvGIC2vOrsxo0yANU4q7+yx/wZsdW2cltVyK+ibLDS2AHtFTQq3JFrqsLlhYg7n45E0X
gC9e2MHDVgJ46udnxFmL7kgglXpwGL72nXhvwb6BuiTKlugzGtuL5yHl7knH3IvSuPGP7s+HhQXY
C5DHENmbeRa9Ay8JlVY2GzorsiIdyp6ORnVEMdMDyx05JRtuvniwvc2+hGR0XpFRYzQYA21RU++E
BDE1DcdevG2PamViXbQpvzyHe//lujJHDC/YvB6kTQ4NOdrh0J7FB6DVJ0O95MRzDir56PXhTa9x
jW5vJlfw2W4v3kvO1v/h014NzqBPYZFfBk43t8F6WszgA4gRenbcBZr1vDK9FIyxV6G0ybWu6U5Z
GdQrPM2EwErjuQ/gINZImJJjWlzW+Out/QlPiHK0xTP9GepbQGK7ERi/e8Y/wwwIKijUAgG0PLYS
lxaRX11JwdJ0Ic91xjJ6Cv4b5OJLlAw6YFZytJaxv9aq6GvgbM3dCF2iR7nprsOFD18P9u37fn1e
y/25nHqmppW0jKUr0Fxu+3J2QVGticS0uwfkxWcAL4YLspRd0bPwZiNVRXbVHWl26Ib8WuAQrIqZ
xYjUljnFqnojh3ETJhMoYUeZCz3i1MrkFRZXd0blf7gKEGk9OO6zoTYtQtsvRt3rlFQYbfwNaFr6
nsFqgR/z9Q6W27NZcunmXvTXRmbu3bDUc2KHKR2/cKnD5FoJhU4Wt+U26dUTC9xxh9fUoWt33swT
IeXndrzkGe5CkktNlKTlz1UfiOv4g3ASUHf5EL1/AgU8G7cFJlUAzTogq488B+fQ7s0xwNS65jG+
0IgPx203IIjqnkGJaiWD3VfTx99ts1iHD9suQH42MeUiVvTEFxf/8Spjhb0RosHlci4vPkfFtFpg
cOdVIZpdNO1s1ogyIRkSLN5WpWv39HFcsBQmqQpYs8mMpaNQ3BdE2Yv39vDI+WlcSNwJcBBjoP6v
vSdjDHD1H5NdzaCB3SoE5cI6RX9e9GpEePp80sCqPHgEAXTz4nCVHbvUSIiODZ1fPk5YG0TmHfhS
erM9scG5fudhCybG2ZSFSK4dP+P941NH7XBeg0MmACvYtxS2Np0y9lDkMZzHg+qi3Y5LXppiGVX8
GsYOYBjklVvG/h4sW+LRfLCl2rXXqAwxrC2IjGL6X36yqZN4g25Vs3kBJwZmqYe4sm3zWW9Yf9sA
Jyhov1Bf43QPf3F1t+5bwjruASH+nUTPwsU8qSA85JMmI7LT7mW3gfEYtuStZKUXyl/s+gHOu8yj
UgywyiTzVKX0XaYUoRyG9h9MSgjgWk2YwXY6nH38Xr1m/turUqY845T/cVB0NB/4fTkQqnZEIe1y
mvurVRUq3iSbWNyesVJRw3tDNwar3w+VGWpXbo2trpa+hvjsT6K8RDjh9liOoZGs0t2gN/EQZNHK
Z4V5XK1m3rF4Od9xgrOscM2JRivkvarh+An+FUCRJO2+K1aerU32k6eJdf70LwD1ivPpuim2D84i
bgj4RMuukriVMTF5Gqw+Hnvs+ZUjgmzTulXfcgHyi3Jt4W9iYyDyGtP+ubBtAunQxzxJjKhYjMEx
0DT+W2pa5HofrKu6q5QbCLaIOctM5P7mGibjq7cp5alKrdm9l8LpIJALtY7estVlgyZuMjFqk8NV
xSu8tDWP7PyLITR9DvvqyyoNdczhkajc1XXTd8oP+gq2JNxyC1GrIxaZKra1x/hLPVxQbNdeRMO3
a7ZwSL0s3TiREwr+fcriUG2WwzntYqrpwDkFekreqhofVWZB/CRJiCPfntBS57toQ9RURQ1VN/YC
D28vfgnerqUQrKlDdqUQLcf5Qnx+gtlj19LrO0Y8b2z17fzymMUbCpUZAlYQ/ZJx02Fe/bPJEysL
MbhEklQ0Sru4UIHiPXlB0b/PgbeiQ4cU4ziXl03DWQ9/xCKk9GkFscYEfOvjhgqj3fiGY8MPa9gn
cR3yw6TYUMYfEbTAmqe6GnbH/hHBAhvbJ/H8Y/vidn78utRlSYx1zRnyn/T29hRIWkQ6dI54Ysgg
gVyMtIW8ZjQyka0NsQoMKdYWOQTm6c2UaUzTRLSCi1P0qmWiF/Fz8GFb2aMLx3ewmgQ/38YRbB+k
YfUxPvC3Wo3jCt1kRt/0pY4+1UPfnLx6dPPSxEubWZrECdDDjvRmJlsHH+FWM08AGstyirNz8g37
exuZicAF9YjCH9b5AxCchoJACk/U+ueJtDJ+BADlMjaA0WjAIVc6UxO0J3prNJXhrZKLKwT65nVD
6A6rnY3hN74Vk15fiVqKZusGmL5kC3/+WZ65U7Fef8CSr2bS6uae7xX03CZpGHiX6MF8PM8xI0T9
sQdGYYSfdw9HkWH24umLHOFGjy1XbshWVZ30w86fFBCoMbmameA9x5pYXFrEEO7+EjLMsqzHf+gH
vgGA0A419UfCrcbuiUUeK3wkT1MTMugojvsNSb3bl+erjWbje151E6jW+lYRDIwKGpNMEa396pvr
udRLDrriGuwc7YUi+kEM9B1F2DpXB800t5bN4yelOOT4ZkTEOuTTsugZj5itPQ+atMuBjbuZujrB
h5589ascvTHF9VF5WNlXhv2Q1jovxXzwuXVjHyZtH4+s4YfkbNnrkhvzKgbyUKu7prsttRveN9Ox
Rv0BW6UeUZrbulSnq3/sFOiVMR3oZINYBguAQssSX/smvyjJMGgnQ3qHRIW+hlFhTxT1r3HDsKpe
ILh25xTLXGz5cAD1CI8MMJZYAS35d7Cv9PWY7HmmJWgePRcrchBnvVTSzGeejroxAchZiSmp+BVK
YKvYO1wg3vsB1vWS+JTzPNU7OtTl6hiTD7JkrkUycqjtNspfOjdZyQxPw4sFR3fsELaRvPSdilPS
5K4vQXYSTT4yt1mI2zcN4vGvlShnWYmHEYnZ0l3rdmZiYJB+NL277anprfThmEqG8Mk6opq251t2
oNQvXnvqssfIAW4XlXIuK3JIx98MDp+0PvrcqdfXueeSFxObl4HnTAjzatTpMUxEDL5/8lsPuCHF
xFth16b7X+WqoG67TG4qe3S3sEcUlVgmz9cB6AduP4WXrme8YJWAh9Ni2DyP6v7JEgQjAHeF1pT3
yepCkXo6Z97gbqyzORw5cKp0qRvVr0WW55ojEu2TA1lc9iLB/Q3qCqMZkqH9JDlUusrzc4ExX5d6
fL7veFDzfDfLPzS/PSbUAlxeLWM7M1b/bCaPuc0UEnOM9RzLfjAlb/dpScQ/XWc6Db7g3QMyhkYk
+F66Bsbc09tsHfJqnXT8aDEu8biS9BejdsDTpivHOk/CJaiM8GkNycidcyPclt9/81IU1yg/59Rj
Kh1PRGCel9kY/fBDbd5SR7xVJtfj+pxrJjPsfPJxhFEOr6uPfz+Q9FLWGRUkmER45rduj1hGM/Gu
F1ueza2eALDjLazNXo5j9K6WE/YI+Z2ylJs2VygBSzTHjfB4XD7a/bnQhqPPePfg7x8ss8wyVFfl
686jJTOr8YAkyX9EfvQkF78ISzrer/moUvj2mNyNdMvbo+L+VbWv4th28Kv/rDyO+fUYVjvbn9p4
3roAM5QPeDYMi+V7JmPFBf0Mo5iwfe068nb6nIEUhebdnoqXddTZdyTc7vlUj++mcz2zKu96aH2+
pjkQZqaX+89Nd2zFupGi4zgnX4t+WBmoYisXdfhGfEbFq/2ClmAz309ORdNrQaAxFE+o/PTh6AMQ
3zlo1YIUmxxkwbimdrKfgBdI69opkDWFZ1X/uZBat9K4/gFY0V8sknQ+oyFbgvXP9j3HjtPW/qB9
iAAe9qrGPEhR6Mb7p1TjA0uXc6p2WlKdm6Z4NkO5oNlEzENnKYCasWSJ4xsScwdK+AvSTEIp9Vyx
RbtaOJm1r8A8pW7QH03BfJdU8mLJhnmzBSZhmYYeOwE5x6uuKO5vNBrq2lOwCy+uq8pk52rMORh3
APyb6OufXV4qELk0VsMkURK1QbSzwKONfX4eM/mRMYIzu/a08tFCzR4L2/WKFHKpBBIog8akdyop
IeSA1r/N/fz7/lJxMEWwgArbD78Q7QHPUnaTg8P4Ub3BSx8NJ6Kxq9KlzJisbRZqoc49SV6Y0VZa
Dw7T6GEfne2vTmy5s/ikQelMfjc2aby1iA+gNXcEhWgamx8OlcGbrb3nXsOiSlgs/OY3cZ/ooErm
frTR5Lwocb/0dbhnsWr2JZA5zkEutVzoft0Lphv/EF0kuCPVNfEhxRc9EzRiXrnSjWH8kpTmiLvA
GOn7Kuz3fpc6wp72deO6kU3ZrOCk1adQHqv2mnPMtBTNvbElQyyjki9Mc/1OcEgRtUpU8zQWcmZk
oMUbLb3LlPFu0isRH0tZWtnLNSgFm8V0mOWm2mR00FBZZZ4KwpCxWEYMmsdMtfISOG7oj/Mebmlx
RGU/OIyqG//OCs21JgDufBJ4wTlkxy+LEralfeNlOgPLNVoQVzP5tbDM/kBdD4iD0+HdSyZt9A27
PjWpEEiba8FNe3LL6PeAfnH0NyXTB+A4sSyD33OiVbrfNqZdRwUd4+0fGnT/1Lgki6GF9a3voPMx
eUvQCWJXEIoVje048vUBZjUwW10Rq8zOZgclB4Lwj/ZBn7fX+fA9rhcTIFMLAUD4sxUxQTzaKtXs
wxWwtayZDfPwDsZUqgFBkouo71B866at+NAeEhqFZ4L+jfeQVMX+YQzhVY9uAVLfbzTxjjRXnXwC
osHQCbqlpzkQvSgpI5dr9iDyzoI43XTyvDPCioe0YKKg8ccJkd/dlER0kRK6WZJvFHtyGyCHR2vX
DiDIuteV85QBSElJPczuMz4CZ2DJMXbsgO7VxgH05SoudM16cvGHa061hUt5zRRTi+iIluhRGCP6
rXhaLiCvw6V4MyJqpScwLKueUIc75ZljC1nGGpUNSNC+7Fm/2iI/ySfU2EiAuzStk4nHa05gATXG
N92A291kmgn6cCYbRd1ZO2iKOrlKxZOruDpBMTA4j100oPOGxTyO15vntzl3N+MEFecZHEN694Ht
BqcS4fineXl641L3+bYw+GZicAy6PewqfMl0o2JuzV7Cwmna+JYcG/9ZOlqr30rc/Wh0Iu+fecbt
x2pQfhMczcuKVzQ07B4HiwBUdhpjJBESfBoLw86afFQs5V9PZ/Kp0JB5ODAWVdxVf/nWMk6S9+V3
kN/11z2kPkw6ryJy08+4RFI00Wtpq5Q8wWsbPIflTNfKkbjogijzX6hMQQ6PbBz3N3GV5nVt1Is4
OCxHGohbcMmPJJopHAZCG5jWVaUAHUVcDsZBMdrM5swBui6OMJoWWzi3CB7S0qAQjiMMj4nkXJRm
VIKLeCjymLaG3HbMGAKuCtnWnH9uQrnAgs3h+ndASa4lbF+clb4iBuVqSISgc0jiYbjyhMFo+qW0
cDexP4KvnWUfDGvZaBqIeh6eTzeg6QKuN21ZTJGs6tEonMe2gtwXSN4PpmfnNbPzpKEdxBuAITfN
dqjmp55uR//UrhoLqvRggCrUSlFNDLM8N3bqQMzSIe/SsgS5WGoXVRpooAwJEOMrF7avpLImvWSS
qwFmvKPHAPovj66CIjKDRPXF3cR6e7FZAUIKF7Jz37rzeb64fAqd5g16KnL+i0gHGtEupG+bFQ6e
XeZ1C74il7HTeYLt4bATPemWzpSX0Z8Aqyb06A4DffNA3qWZg38o5HRe8lrb1DZeTFIBQ000egdx
5L3qpq3tKMHOTFL2ONm6AbnlaP2aqo1R48p6wY88nC5txNd3cfqg9zYOxZPzj8OSktg5VxsrxglD
0JHy8Dk21TffOoxp+SeGmuIBZvLnGXbz3C0QEQlnTrxAbi/Jh7LxHFhkas5qRTsaM9conON82wYD
1nnYa82JsoGZJyxjSxaNn4kdVLs5yA9Z7c2USrPfx0Y/7Bm/h3AIUAIBJa9Xkxp2Eh4H3xh0A9VQ
6QF1a3bhiIf+Sy+jgsMq/BAnrfY0ohqK40B4p1fX/GUV3w3+TsEii4ziw8bNn4YG/c4yAZcuBGju
9Er8N5x/oicZBuKnf50Q7gsbxvRpyAZrSBb0xtc+WkIjTMJ2tBvmzOoJPwkXr9phaKOZzZ5qajKk
j7nhpO44fZEQQ9NifZbIF5qXAq2TlDHToDwDI3e3Wfwk6nu1MuSRRLRbLmmtUvX07Fzjn+psafKl
UgrjZPSUd8/NP2/BXoHgOW7C48SOezbL/wMAZ87S8C3/xaXYCRJHovhQitUZ+TnucuVlq996gvLM
PnRSkehe/XoZrESKhgjen+4Gttt0X43T4Ca4qBRzORFk/M7UnMLKlrRkifANlkO3zdrTx/ry0BUA
RVKVuWahXbuq2UACCGyZv0Xe0ofdzPahdjOHeg6GPM+Nr1OLkIcqLxJoEPPjj5k8Rh9Th0H4xz62
O7Ju4rUB+q23gZRXAOi8qCP3EpbduxMqIH2+Hq5IMBTy1BFAvvlzv8w9qYOuOgpjyHLnKiJaOR5e
PkD2kVpllHNlKCfeCvGIm7QrzJW9clXscZZFJM80CJMJ3R7A5cwiyKTOYoPa+yYRusvyJfGj/788
niHK4Bhv/dD1Ds1e6aKR6h7XXZZ+kWriRr+qfVoe4ecTMFQztIXRx+n98tXApaXzbnLvUSuEhNdg
op40dDcjIMkfTeVdU6/QdZ6cbNFiKxuG4fToEIKrJDZE9KXMVjKSV/WtdRJbmZf4cxaAZUFxPbiW
YzJEhBS7n+ZyRldBfpRnpwHBvVxsjkTsbVEV+YuPNVwWa2omfCwNbMFp3Gt1YyfS2fUdtJXcCq5g
T9EihYVsLSXwJloj7URQCiQIHv3LinssXjj5j4kdiJyDMpT9NO7JqTYYUpR1PnjwMxAEm7l5zdXi
lnyFNH5r2u4aUHQ1dbVBJBdAIzwdgizSv9/GPEdiuKY8Yf7B3tmIW/evMko6bsyT2a/XQGzK3apo
1OooxYXxAVhDLal1rw66KLdHuK4esBIa6hPMgMK8ZV8USSDgsWkUA1qpJSFP9azn+X/i+xK4YYmZ
n/vFb8+dA/VujRB3lp4CG23ll0uXTDVd2vZq8BwDhr0frYeOPla7S/khRrcNl0Oc8iibHAmgH1mX
WHVP+W2WQuzm8IB5xL3+uo0yU4Zs7tUZKPSGBzMqimcjvvZEUumbeLdyIHbsGn9rCH/cZ+5BOLMe
uJY0+hnQ0S/oELfXTYSdlM68CRZXHuPYzVj7JBMtBQGSvqA44j/S64+L2Lr7uuN+We0TPpaWN0wB
dY0YatrJLVA9o5fUgQfT6dAr3b9lNhyLEFQ29V51mw3aKlz3ikOn9CZhf+u20zhV4RUe/vuKNIaC
NMq0zEcYnujeugXdNWh2HIqtmMk2GYd4dn0hgTwgwXRizaanHOkWtUKCFD9WE2+w8a/3FVuMl8ti
cpAxnrS2TG8edejm7cJhlWI59ZbFOnmIZmzM43QUINuoTbyOYZ7QHaeVO+ez8Oj5jla/TmNP+jrd
01PDd7/gR5JSNU6rpZt7tFqTfhgC5SpaRKZrj3o/9w4gcx3dhvS0jyMeKY9iBXd+DmZvY3cYPAHK
T3JH2v+nrJ+VYaHLuHaBpg7gOjeR26tlBtd79/GvBzapYn79CUtrPmBpK8yKne73CTvJdMj1usD4
8NO3j1xPQg8TocJCfEXlVUsFTrEVVUXqriNLl2YIoQTNX9llLtKFjzUzU3CbxM3I63lAzgFiC0xb
L/JoUxcxQ7jvfo9omYWpxZnKcZPC44ojKw9UDFw6kTAqGxSVOERq1d8pjbM7yK/zkgf4TDy+cA5j
q2oiUu4lX3c8W04PJIA1Ty2zYrfx2mcw21LZKq47mo1iKkb8vnjKOsXDjRVcQ6kXmjG+yHt2y9RJ
QNQJY6s2igiPbJAn8aeXAhCW1vEh4MTfO6V8M9HJ9vx6ZylgH7u6VAPclOiKtFG6Dcr00lS0GY1l
FSnsqpIT7sqL+mh8+PdSsKi428fHy+RwJvn4WS4GShOuxiKJ2OjN9MwVeNE/fOP51FSPWXgvCEFs
1hEkBCc08eur/iYvvKENWc6M7zZKUuqLkyFnUquf2mIuOpQU9b9sC30q5GIDVRHuD1y3wVSpijBG
LDnWgrWxDavGFjjo/YPg+b5sN5I3tn4qe5dbZuUoqC4V0coV0qxE4/YKSy+dC96FdTDUpDTu2YOU
61HxsRlpLO7HJGvyzOJQxe5tb+B/efR3MKk+XSg/K9xzrf65XxSjIMQ7eG1TSRtujd0+OAQKirGP
evbq0Dy0wpPvvQ9uV30nioGesH19UlbMng2OjVrAvPBbsJAo31WMOyM4B3GOo6QwUH3HdxlhuXuk
UELCyB6i/EXHxceXwfBTMwbKO5tZcZ2wYgiAMGTUrdLP/TFTrvlkTBAIaHJ0YRKXMRvbXDmKd3f5
hCtaGkmcDNox7qDVoCM5X7+2a7VUF0/sTf5JI/mFsI0c6Hgqdqw2yEUmt8KsmBuk799cfZ1paC21
UIxBQIDst9XtPRyPr/4AjS2GVypfddAHfANZPt1QtxdMbkpKH+E59FktAc4WOZ7bC7Wqnhf4kuZH
PxAsi0ell4Uh/Z7mAj79HScekaBuTdXcqXA6t8PKUugnA1XrW3HTuRwGxqkGUeicpPsr9mIHwlrj
oHsi2kWmhuUYv8ULYx6XFmsSoO47v067FwU5DUsRi69wDj9pU/jCwqEIOzyiNMwARRyYa8JiMym0
s53Qi4RdOIMmpiNAwy6m7H+jEkrPlum9FROXUIJK/mw3Sck0hf1rPQGKM2EECNAceryXLBJt270c
65ibqIEhsa3gAky/bLrTGz2luMHARYnoaWotD9aEJyFkJTi51/WhOERTVPEnmvcesAPVJLeqpPXc
Ejl6dpDOAcrvhhJmNsEYAoS+bfvRJRngg1rPTdGqWMTrgwWAYEp1vUJSRDgZDhddSPQtWDOPvYjX
ERb3SxuB/D90Ickb4Hd9Cn9xdgoa/4XuC2ruBqv/Ebs9Cuua+pKMUxiWEcGnFlUxZ7mmp5DUncAO
6yYnfzvcel5RY24bXpb2RE5Dy3nXEKoT7Uu7VRjpVVrEXUjCRgJnxlvfk9P8tmoKaPfZ73yQrzat
dDNIR1EFLrrSwEY/EIfbulcdxL/Cbs8PXROwDjdcFe/wQSAB5mlUxFXqRHJsuj3yaAw4yjZ9rFUT
6TjXW7WygM9SY8t5H/bmuqWFDZ1vD+xvR1CowJ4lEkkUubT/hNmgfQHjzXTZFQ61VtK7Drsfz1R/
mkSm9mBhqyZKN6F5/Ja4nQLJlB/lejKrj541M7JZVy9sx167EbT/rkaAKhXlHL32pItSQ8NPIvIH
b0mdQUELXiQ50hnN+z3isaE2QsOrImKwO9NHX89OMleAZ/OvXGjvUjjwbjdY8cBm96SvhmnbniDN
JhOaJgtIYvKSpCg89pK03OM4ZHR1eJjUZLsuxQqonqNWilEt8Q19XPRs5HCQuQoX/h6NIgMPnffU
rhmkUmszTEWNTpYkvftF3GcsBv9iaCFFkepBjgxkyGqnxbxCskTmTRS3Biq+H5uSPv0xJBTTiiqV
m0H5EK98utrI4rAgdmA92E/Y/QrRgKjCwHFdh/1iEt6U9qlyU6vkPkBcp5OdsRcdqnHqReAqoeb7
h2FXrliRNu7uMXYsR16R8npZKVvY6TLx/bo8/8qAnhWoTeCT+baC3qkgPGEzWhxwbiY5nTNPvt5a
zMdnWwEegFsIvTYkprfXVG9IojHtFugvHq61IYgS2UM5jRNCsU9e/NDofvrkArVig9X0xFrRUDGH
uw/ETpvsLIG60ffgMGcKdHkUXt/756Z6RnuZX3ucNw/xleZTeIeDZBuzSmAW2z7+QFuf1wdYEV6D
DFyqI4L6MYkChb19otyqEx7paoAt/IVV+igrXf6N2iXb7zEWl0X0ql3CrDHnL0WVM7Uk7srnRll8
HDzU7h/Kvul4DUXP3n6QtT4GEl0Ov9TzXJFtOrbLw1n0RedzMKPiA54Og/b72DYnjgPY/60hb4xU
T/d7LbvuWb8Kx3TulkqfniX5gK5I5KewfhhiQXSm1+uG0pubTeCUlYrcVpHFyMq6fG8GdfcwtqAR
icaDLZYvFWlhvFH4VcbhnOeiG53jxyq+OBYQ1g64QMjHUQlqwI2eTCMj0VJkIZXiWMVMO+DapMhk
JBRLDYRtjph7idFxVQcp2BNUTIRDTLlOMtk9N0jWKN6Oc2oUBFgtGsG4bwFyY0tyfxydCkZh9qWt
xgrxG8YcEnxgpwN6KZ/HUR7wigBGuQdv8200j6GTZ1skxB+qQ3ADmf1vRfw1sWNRAmwdT/MFKTN6
z/LVtGDS5S8nhnz3qhwZ/srtQc4Z+PUTm3N6doU/Ltp+NN2CfcWqjhwcsf1VK5QalNLohfJmTL/f
5Sj/1QztjzQ9goEgyN1pYnETyHRmBnItd7jQ8vW7WMy/Nl48AvhtqhaocNUGJVJVWok3hqE36IvG
BjbH/AW05rpBIAJWQyfgpU51lwwMqFO7RkdJyl5d/9yZwfkWNauKXzqHdGPuYHDvdsOmY+EFb7kS
KI8OF1cmpD/3dYnfk72eruJI1eutXQdhI8qs0VnyLn2CBCvYiyXcUYeg+e+6g8H/lRze7VyvXGaN
giXcQIfhUSo81KAPJ7CEesz5kU6wE4qRgrgNFu/QOKsGtoeRzQle25kHJ3RjRRv3+/mQeLi36xQ4
8s69KiaFoTpp2c6prd9g+gpwz4zsbB3Udjbtuxdpui3HlMH1GFlSCu7kWad67d1SSfd7WsjvMbpj
reDgKSjvEpyRknYt/JE2+dzCx1c9CrNBTYnuL6DatxUuAMO42P1Zo56aVodY2vlLm3ajZHBXK9xI
ZQngH2EaAVJ5fWlT/mZ55GRLd0rrX2IJGp5UxOla3bICDs95QmOAsCqgT9RNstkZL7jzImw3Tv9M
+So0s6NXHoR7ZatpAs/Vjm+KTC/xZD9SJhCoKHt0634g9EitHm5FfGwmMb7PTNWFAIpY/fy5H1M8
tPZw0q5vF0Cs19PurIoa+QhkbkpXK8AWfmxEHwWGC/Edp96S9r8O581QfE36hp5W8zyoa9GZm+ZT
rCHtFB9De0L7ADAaIbrZkcIaTFgBiPMFKdi7OaJHy6HzpsHnwcAdFp4l3nVNeLpTEnimfnZcX7J/
TniFpyeu536Eu7ICfi3LItcpzJ5JazJmSVXgTem/iM1ICdguq/q8kU+FtsEj+6KyLmzEtdjSBK5p
/lB/EVT8FE5YyOprfsrrjUvZIMCXON9x+3tXL9/o76Muof5BmVpcGIJOVbpj+vGQ5ef61lNro2Xy
4+eEQ10k0OFr+cUjmFTq2mtWSlNkeQwpUJ+4qNTXNK6JpjU3R7/spTgiQTSJWYn1PReOjfdh+J+j
3PZoiuGa7riJgFVjA6Z+2OmwYodREgHT8UZDiUx9DsCn7Z2V9oKiuQvZjR3dSW+TRrf4iHXZKsKH
M3pXYSTzGZO90SjI7cMBB7E00aLMqNZ5YKfP7yVgxntsGx1EBCuJdKSsa1HHKHWBEr4012NawdQf
/CuITLsZgO2IAy7kk7dLZJr95nLldDh7Ab59a2hhbgm2FBpNzBW9HBA5saVN4Nw5cD8tNc4UUs5Z
8KYD2oc3MjXCBFC3Aw9FNlqwnGUtVROyYLImupltV8b4tHpL6UqHuF2ps76Mz5vpd6xhRN4l6eXi
HiuFoann9gnwt8WYBcDL+pLs3hG45IyYpCGmOlIojWsWm7R96aCIZtoqbzOqwBHloJmsQwCLQFtt
CYoqimjRVS2cyJtDfgm6Ju+Y3FNYf8aNSKR2af1beguCDkuPqF6GxBupreTYUC+nDamsHxQgYB8k
2R8GWdpGg6+RwkPu5QKOeXqHtIfG8GIobO/OEECO//wIxR7XemRGDdgHejl49205BmmjZqJGrXW4
nm7j2MEV/QMIB/+0Lp+zHLq7JIawywl6Fxrc+ZX0SnCsz5vGpZF/7TzqyyP30ipsUnCIVBdLLBOM
oIo7p4YDRR6lWpo/3M+uMSgUtH0TsbMwjzejJcd5gGcmJrVWlKTCDscTTiP2DmEychqq5tl+pcO6
zuvkLw4p3YuK/f4JZ9pDqr+F3YUluRrer+K56iUh7xf9IjJTPazSEvaQ2UMAwDLHMCuxGF/Hhpxe
Kpkuk2Pe6dtckimeU9eA8yFCKnLSFwse0UOeW0FouGUOY3Tlk+DzYO78xlIjLVO+DxgsppxUO26l
9sImgWbF32k5/Ob/VASBWnFxjLaYrkr1ufvTSyjb1vk0sa1GI1YJ9+9TkAZO4GYxfXSskM8B8DIy
nJyBQw8y18M5oRcBJGjJsEE9Hj8rT8YXqyvRdPPQ9FzsKGu6r/enmIYU2lV5sUwfowiijIg8b+um
+GVfeQo1ObD0FXzCB0A8IujeYG/Xss5r6PBrnBkpLVZUsf8cBpXplpg4h97Ysc4wnEgSMSysuTW3
fU/50NMzvBUe7yrDj/FYHJubaM8Y6AHif1n2W2+qDjIIhBt9il96EUH+rZFUxhnINdZ/ZQTTr5Is
17WHiTGKjFpvSWyga2LGTl4oMOiVZ2vjyRISiAB50whapsvJtY0pP2ou4Uw5MLRCp0S5Z0KOQqn+
HHHdkprUmCDu2XS3B3yg6gyIcm8mt6KnMl1/3Uq2pwKIQlF4/AISsbEdn8YLnGDTjtBEGEtFkrzs
tNFBjqsE/WV4YiXU6umjSVhKbKh0hH2hjTZUmQdl6TCEWj96Q6DuJhR5qMI2gwXapcIM8rkgfl0x
lfALs2iUuJB2sEvxDg5VSU5i7DtmbvJJaacOb+0ugcCGaUHlwXF6Xwyk6YYm0+u19BU5A6FWEtyF
m2KARiwnULI6TzGlqDZXqP59Ml2TvtZ9je6igUj7Ap2Hpx2jI1J+PGmgWzKCfAtCxNxMBmxT7oxn
9wvPZ+rP45deGbsDHaV67fY6P9viiYCmAl8WVCAnAVB2JgNp/TTViVJxjpXBxzgCgtNa1BK9z6hd
SYGRTiX7WBFoYNwuJr/6jNRelxZj8qB1wOWGPy21KnAPi+jEwAdehllXFXnA2bPk2Xoxd3NKfGoI
EfH482VkmN2KB9uVxj2HCrkjA1aMZF1n1aXCiLy5v3vrNE3hqmgsl7909IKYMTcsOrsv0esoqb3s
Q6W7pnFrXEX1H8mn7lWviwXI9BkUpoN2MDObmxtHemW05fE7/M7aQkUyUTnsL3VnS+uh0eiVelZv
5UW/YNI5cIdIBmTLWvc8ePJdeMqR4O/jXYmItQhScgTQdHPbqB1f6lp589WckBhmRGwhQOIMv81W
7DKM1UpAXq6LN9DqW9iGftEylST+rhOYmVKsjW8T+FxH8NADuHmimlB7NUuT48x5CfhOXduJIR/b
6lrhdpIXhMmBAeYfs9hTw8TubBSgKeAvHKLfRdlD58aJaEoc6uTEGgFkPshdwFLO3sgYt1I0RhJk
fiKUfxMsq50hAjOAeva/K6Px1mIZCjyanyuyID4aSDvm7C5qI+lvnx6ajZqdHb3OlMX39fByQHJL
aKWAg7iXQ9pPdvxKG7/qyaP3j7xjfJWaPXYSDfD1/00W3XnibvvgddUXj9b17m6dWpS6Hok8aV84
h7noA9oRzLRwlFqtLduGrtJmAZdmZv9ZZ22iD/csCf+MCHnU+tlc0ob281csbvJkKgeW60G4aKDh
Os/p1TL5eDqFHamBla3/M9hLF/Jy5f6z48L2oi52PM6X19ZmuUaulRky9+XB/4Ux79ZO1+ZIGTre
zlkL62AoXjUwtzjBm3y2giPIRIm+FQOoiYVGI6X753g70ADhxJ4r1998GuAhO8f3Bt/blEmtG2R4
OQGgOTG1wy0AXFfRdkAo3+EsY6W9KFiKDEs374tIkEU3yp/dRSn+2m26e0ICa/x15gmoEk9YIMVp
+/APMXvzS3y2C9eCg63EKfuDF4+8DXce8zpFiyx9TBKvIEEANyrJER9oO4kEq9jvUDMDOfDlcU/l
l1E+lUgmoXdcL7sjMGJK2P3xWkPtai1ZtQ7YFbLnt0MjgvfHbxD2j67BXpwgpK6a/nerjiC5uw1H
PmCWUTMu6SiEOZRiVwDhipz62Ocf3n92rXuDUNNEhI67C4ZA6HWWF1e6JxAMV6KmtYJLcIjbJxHj
C9Tudr/Yj9FHRQjV+QKdIWtGOQq68NzlIF8nEOE4fPZtXmVNl/e7gj5QmhW2fPuCDwUn7uPDLjmx
hllbK/DGdf6sxFhbsQZ4YVSOiDloRNl3Q3CoNaOQd3fHARZnXqqNwc55ob2d3gLYrP6S6GIjkXym
VPZySyBEjxE8xh7Zzd87Jw2Jx+eP/NvwOoaRIBZ18YKBQqeos7Rl+HfunYCSU1JFrcf5bdkeKNHS
1oI1QODg0fMCQI3Tq65JzOrtLXzxkpexvW0CJHFIoB83PeoxE8yFyvCypl7aF7M3sciW3gcGtd6z
kpFMsqpgfow/Z5XHaCMVw04cS/9Ac60kU1KcxwTvsurQeEDciJE8BC7pDRiv0h0E7WJl+G9khe3m
VAD6nz4JrRM/TMBkes2IVGpxR8nL3x0o7fxlfZXQNa4m9neUY2Qgiua+Me1erHoBTgfR7YvhT77j
zYKzIWaEe77qHZej5jpNRDPo+sgs+eDZ1xxnEQ5VtE223IFS/zS1QR71mbd+mIcBPe1WYknTgyf0
jY2x76E0c7+SK5FMLZizW+Kkzzk954dV77Kjwlhk4x1lRrka4X77r+91aSk3YBkSGxiMUvkV0Fms
NZqYZN2UwXvc3CIuSAEAXMlqEpBQ0cGgbrI1GWLYXD7P9oTVWJBgY6bLpadroedoUqmllEFmhCkk
hI3qAPPYY9pACfXllmaC2AcdnI131gyMhUv0V/+6X9SLne+Hmn8Fm+BZgo2Dvcq/zJss/2glxVZR
4Hy+NrJ3yJW0XML4twJQMOlNXZz4ds85x5ZyPHh2FrZMsiv3TRPmHfICQFsm6FfYWTqRaEe/xmWw
QG6WiPL/iNZpqmLOsZ9OlY5lAVobqvaFagV3K/7Iy8uqCVvE4g9N7EETmYY4J/LSoVRag5Db21u2
9hODKRgWCoVpJqb7D/QfOkjeNm6Nm/uDMuMSWtN7jdPYOrc3W02lVvoAB/UVHfk4VVKwLRWodg6L
m01Pyh1K+o1FMnMau9TxJPWizbszFAl5XUzRRRkt5tQZnYGhGKlEseDk6Jg4yhFcWjZRPBWTzvdM
gr+AzgA729t2E4Docp/S9qtqS/ZOYCb+4W9fphB6t2p/NsxUXvBDC0hvdvDT9TzLA8/dlrZITwwP
UZym3i2WJjghI1kEP1mL7yT3FP76zDbYVFBlzINnwDSejlirbsPjZEpRaOFLuc63zFh40Roaa7cR
OHgAkbk7YMahRcgJ0eK7WDtcVQhm88+cRJqkwlL7hYDKaSByQJb48a1ULwyTS9OTxIoMw3z7Ac15
G+kEw4wE3bUGFwq9241YIgx0wa2C0n24xJUCwmla3+wY+mauUhGYec8Uzz8lrMRRxt/BzSkSUfz8
PQMdWtuCsOXpzA3aft29M5JdBYSdjkbQmeXZblKIwXy42Gyshd2mXTaLxzIGDDVImWv1uKt4ZPAv
YNu4/KvNGRv/6gP1wMLo0mf9KFdRXH4Bxffc8DRYzYhuv5a3yER+j7+9FWF6rlrs07t5UzEWE0lW
qvyosUvr5GfEnUIEyueWDql9Hy8pjUNFS8xgT6vo5oUVCJ8LXZcUMDgi0HqrLaNX1Ym1ZXb+gOXp
ypuV+4gfEQT/mhyvqWUjV9LPnQsA6Y8ichNc+s56zL+clDNjK7nRtRm8Cw8mwx3QwJhCpadrj8gu
/8vAnsTAG5GjbeWNDkcQNf786iWRavPV5idE6spoxKMuPJ4B1jLtbLLi2zXDAhetaG5Svqz6F5lg
JxDm2PfgZkJhya9Wv7Mwuv536qQXmNOxB//QfmJPTcbjOtsRFCvnw8Qg44PC7S3DcqRAO/kzG9rQ
HUVgwpmEdVklaW44ujxqqBsz5OXsj2wGg2AYMZfvOSJpNOvpWFcnTgmVqJpgcQI+MHrG/li29wYA
2ZO3nUXJ3+q1fYCh0Y+HInW7d0N93NN6WTe64fif6W3fxhPYKDPaaJQMklngYzbjzU4HRDVge0Xy
IDsuLc9HlNvcoByMd6Pq5TAOUwWno9eB+oTreYUlyiPhmBTzIQDL/yyxjNupeVIoUJkYCD5ytKMX
/jhlZW6IiBpIGDqHE5832jcbt049QO1fbOjlmTBVdj41/moD16ts1sjcCkt+C0N+BfQcidXjV+DI
G9IRHDwJSpCwYa+bvwbzBltzcKnsVQUQs81SnVu1PrmzXusumsDVBsLm2V5y9PDd/JmjbKicvxVw
7x07ueI6E64InVQz+INTp5QEeLfAmrQU3OpnJu5n/J1/8MoR+4xQY9zLPgoMxxwZ2uZwPWNn1hXZ
m2h+pfRnuFCINEqWszEoMXa4v6r/jm9KCpASXJ4wAradvZ6XUCBQ8oriDh77ZNYa9uGpJ1m4VrUw
hd0oVDS/PUtNJJCjt900kJo3X8YtAhmzK74Ztqui5juysxnjb3BJ1xphJYTLeSH+i5ORmY+vtdUK
ZeAwA/eUCjmsgZmeFcZ9dUhqfmLhdui6GuOLDlii6yx6fsKZkuQmdM/TyL+y3/lm13Yb37USKwlt
ZQ4bFb1OKdt7T9ChFqaVDbDib/5My5cHac/scUp0wFWhbf87fg2+hEK1yK0bjLsDqRxxf3+Bi0mG
JbEkyV00gamv64wxPJctC1yLpA2i7JGfp9dIVPCBlDDmgf1NAT1uizFGEMq+N4DhYLAWsM4v77M3
KtR8lf1zQlSUxaxoYhwWspHoSnpbQgQ94+iQprLPa89ceb4k30/04wTs9GyzkGbwJabmWDNCdNxr
QEX6Pgp/zIBcZ9andzTJCclJc+gmDNi3vHIQNMmP1jMxeU9FdYWJ1THh5vxDJ6pjtN4JegM6blXC
Odu+qRK/LT8z/aLWHC+MELKwz+yO4gR0RmhS1pHGy++XansbL+auMB0W6FRKivagClGv8fySHq6M
64q3r97EeeKthTNXlJrI3gBk6CR7v2GEiyBF1O0EOzFXQCIi5Mu5hsbBNKelsATSXCzkOhHQZTfV
eaksUrSJgWlQZUKJP/2VpFaoecd+mh93yiTLH03CXNedt69BqB7Nz5m2mMrWdqy8n3uG2pnNRqPz
dhzpLqFxL0gqRRpI7aFaiskyxi0bjYaMi9JPWftHVRPGjUo+mQSyampYWIaHk7zbErkeniSCN8Ot
/D5iaSvSFi96wUTYuFl1wTnSGTmMX5aWi+jh7HT1oG0Z+BHkA93q6nSsh+T4Qzp1etBHqeNomLLZ
N2yy+D40erHZGSUv20VOdQ211Jiw4R2Qiqdw2VoWlpmh6K3z2esIYV1Kt+Jc/7H6xVdK4xuEj5ax
elK0uoYKoDEa5qhPQyU7KUAW9b3RJk+xXwUOGMjtKLEq6ONfAeDdVqkQg+kTPuiVOBasCQX07NtV
EU/Okiw22YZb9VNxACtQ/EAK5+eMmR6B5xdSk5EPOAcn1smcEnvGg7udVN98wevitbXeiQ/Qeu0i
V6Gfa4IRzrOfis2MoxxXNj0e6EoEAH4eIxtxGC6Da6IdHEB8zeUewmA/Sq1Uha7un7o25YK5Bxv/
TA9J4WBLjM4a+3hVBdhIa8Ep384A3KUkbm54nATp+jM8+px8OncKC7KlcOQjIgiQZmVRvZ4Gy8ma
9wbjqu9UcxIuK8+lh74B3fOPb/jd6ucd1QeW8qy7mgaSGKfP8rAiQ7agVkRV8yj/5iYLE8LJ8+OC
0Iv8cJ+EgdI2UsnNLpwEj0EfrukT+nYNKQLUzZipcI4d7A8TMCAr7dru4NKYl2HwvmNYWWc0/0A9
UwfXPNj9MGyJkSiUXRyg4d3ZS3EZ/w6SUa3JPTgKyeNmXLghyEDq0rI3jVJqzjLQC+L7Hs0k7f0u
inSaDBx6ujziL/b+cCHwqchPTdMf6rd1GAsYmLYYE1mGEEO+teTYn20Ga95MIVW6htmC/6/K4VA2
ZST7Kq+BYsXb6R3Q4I/JyxZ1R1M0tgPPesV1O/6F+6gmq1vqiYQjliXYrK6flt8vcp8EA4yOCe/O
ZuZIouDV8gN0uOr0osmSTx2aSsD+mTtZjEWOQKUbjekBU0GjE9lBpzMYK4j49gEi9V6DNnLaAWm8
S0pgjNv7OtJWBt7vqCzV1bOBlS/c+cUyQ0OC7o4ZrVLIRwR0C4/VBi0P/uUjAzr7IPbMObnUUIkI
QPKbNcc+0X3p5HfpHQ8+CEyBhyHoSCqv1ZoetHcJYlbzDBtEiUuDxv5VlYk52NIEIrG8Y/FBfqfF
2BfQXEfX2e0hjkHwN1JAtTGEKI8jTiCT4J6bx+0peiiu9Z/31UjNsyFaT5u4osYkL7SuZ/oHkm99
OI/ZU7hQ9dmeqQ9cOZ8NH95s2CCcq2Bq2Fo3vgtL7rqG5EYSg2yi7he3TJYy9H3QJmgrI0B/j4Tc
H5BIusZE/hQWUGWlTj8vCJk8OM7UsZFjw1ZNsFZoh31E0PjAaA2n97rTMZhk/S6bUFho5UdW3y7B
xsh+ASUDdXGbg8yy1TzXJe8xNwjjWq8iI5MhSoykc/3O2m9fDqHI8371QMDV0AoHqTctOLPnHOCI
ZaO5a6W5DMYsCIe0vkEuWJ5xPkZ3l5QFoMUR0/NTR1rQwOJwZdzeYUqbgyeekm9VYqFwbw0uFRS1
/6LQgzSXZarHsTb+OG3exa88ywAaVeP6j+MKmYt5b4nPXMTSXRrFFu1UsyN4pG197mp4nOlMxyWn
VW0R11WDCxACa2CwgDM4gazgSmDn4rgr75zyAbZwQuVWn76lkrOA8dKGb4G0/GUg8eP8Ec2rvAWA
HFWg4prR5zYFRNQO63HcLrxAp4jBzEy+AOAq8yLoa3yvQKSdQLm7TH7pjH+yfkLKJBxk2db086A2
NhFUOs9lkY+5OA4SFb6q69Wk5AFXbZh64VV/4RRuaN0McVsiKKijpxp3aejkls7AkS4GUXqTEYFG
8SJWtvC9rTKsBs95gmeLb0d25NhFXRjS93dcC+sPnm3EmCqLz6TCaJ7qdUqDyduNdH7/Umccm6Ua
2RWwp3gzWOZeDTqxIAAgMR3fJOpJgSv66vpGMgONSoHuycfbjPwusauKgnZ/3Zk09u4459QtM3ZM
QNWcnNbMa+rvPubsegD7vDsWNIG8ZFcA9t9ejKa8jv1Wer7K8MpXtIordJIXo4Wvd84WOjAK6YcI
CtmMMByoHkD5oqCD/CL24B1wRsgZZrb8Wq+z8ACO/SSee2jfjWq7YXygqeQZdNJHQlSwOMVFETJJ
ykjr2xaNq0cPP0c+07nJjihIhyHFEiWhUeVxATTnVdfOL7tgbgKvpiFahc0ItqBRxuMb8C4HZGEi
fxPLOx5D7lW1i2D89cFapN6o20irGY704RRJfwJLiomiDYNopftCMddR9DWJM2YrBYak/NKvZHDm
4rLChrmYA6xxxecZdsIxdlBbcXH53YRFvAfJ6t/k/HF3HbaL9vlHCKcXerKHMVyKqR82p7Xw3f4K
74keakhMq/jyoJlIzOq7i/HOvfLmlnJw5mWMQnfZzj4jufR92DbWeoWwyCwPHJ/WGKq/aAVGt5hi
m23O6zB3i+UcMe1dXuRDYmZLhar3L+AtF/Qn1pJP6iq4XhygVCifJt84gVj+eBVXVeHvmjg+zddb
CUHZmrpIYy1WKh9MDrTk1cc1PiHy9RUZFRgKtsFhLJC7vn4uoVWlzka+S9KB1YfGVxUX8gLjeF85
6st32sykmfHpViAgMaaahJVfZtCLS+6M/aTNLx9bd1gbee8mN6vFaCzo2bQ0llgO5F/cmA0JOCEC
djuWM2FaVg5hInu+3ZYXNpR6/OQnQJ3Rz81m/+IH+saoNzWfD4peMqwBjssfRxwCHor/+7PjT7/N
Pd7WBPQs+3H1vFBXAiznRy4zdYz1TBsmpExBs3KNpjdsjacpTbajbMa3agvJ/m5YYg6hEJCkLDr7
injFQ0u8XBMBM5xoaIq+eU6vczzd0C0uhMkPYEiXa91npCRnAjSGXrGf0e6yteVFmnc454Uvw+FI
Zi4NFxD241m/CITVupHHNAU1W20AnC4MyMx26myiaqXzBmezINm2I8/k4/upbeaaaNHRBGgEE269
QGfelurGKC6mrG/lK0PU2u5PORZVPUqmmspTQdEI9K3LJ0HrhJSLos1OC0usfOKYjlVYlaa8J4V0
vRyEWiv8Niyugur79wPgj7V7N6kn4wV45H1TCORuScZrG70gBGtzo+zw5GUUEUbb8kDrSWpGl+st
gPZ7CAbbmG5CDjhNy2RNSpE3MsCgN4vLbdCvwnnrJ5IsG9KL5rGM0xraAExmNjKj49LsTqjov8Qv
SC+HB4oQ7ZYaBaJsLSQf8qUmw39TvNQi3p+KYDbiC4U05lEIR7DZXjLrh5rpwvUZtiYGcVrxKACE
sPni8FvGIIafwOmlIqu0K7yWxJSRg6xtlCe6UluMyYhtwLEkWQOyOHGPqfA/pTU8YB+NF3eZ4Xrv
oxOyMTGXlvA4S9hMN91WL92Bp3kVMJ9TqSlTOguz2DQoc3zqSuGq+mfVT5ySQ4OAzCCEBBUACwos
bXaZV9KkmPo4AhP7/0y2Xokq2qv2FV/TKOdaNPOiJgfszq6XctU5JOXeHpaCHTddvVBtmBGnTuL1
3NgcI4cFWg8gR5vP4vyQcTlYZbShv34SSf69sPPVs31Bqb2jKJ467TNkyb7spVeaiLlL0HxVNVfi
TteaYoLIDEDJXTAFUTgBwCoBGy+yjRx1d8O6hocx3+EHqyPHCvcMIWKv3ZcQHK/nm36O1BSSytYy
HVNi4V45dXE5XgVNA/MCnNXe7ZEtH6hJJCJTm9zqgxhbhzLy3JCkzu008NrKm3ksTm43iBPo7oKP
6imNwVdCyQjWFDG2/lx0rlUvM6le7LnoDNwxfTRlsMLmltQDLZRcm4Ky+JIugzzTc6gM/MKmSYeo
22MotL9O6N9rSfYzuzZPWu+UWW2B4GFol9WiK4XXVOFSjeYjNKWdpbJC92YZvpE/cEanQc/YHeg7
7BViQ8HHXvB8q7OnZAdHTOPGQYcQawm3IJelHw/lJAJiOBZaBh87Y3Bo16838nlQqbXy8w4USwLM
ub4MIBZIPG9IOVr2O+oqLcweCI3ucDYjyRwDv26H740wQQgZRtPlExI+982jPdPaj8NrUlda4sZ3
T2t4xFJtLSLHtrZsa/uuC7Irpjkv+G1gPoYlFnJvpGbYRiMwUCd1EKvAJ7g1TVuhvIkgRhMWTV2V
vXSS2ys5xavmSqttq/VvSOBCc0Yu8LO3zKdPCy2fpfNh6L6PD1C2tM0iH8dw1fM/rU5QjzUTGoA3
OwKXS2M+Gigj/S7hTEI0Ki8Z1a3Rt6yDqT9+BOE8Qo2xLBwn/XZf8w5e64A0qdmKydCFmNmi39U6
pqgVP+zRqM4zTCCs/Z11YxJjblUBbFjtWkngb8jX5Ndqn4FcEtDxrOSwj9hg7Xji8bmurBtBtcF4
ZX95ctbdDTde2fvgTAr9IHYcYu/PxZ7WrL56J3TDTkQkVz+MRnONI85c6K6732lNXVRHrpMEqBcp
34Idb6rwMCRWrZcq7gldZe5NITmupZyoMCDvvFJ8ES7iI71vU+EVDmWCC6SEVtMylgBvnhfIv1T7
1FCxLhQ95Y7bCzuQynbiPjZ+JrTa3Npl0UGLRhwGpAKmwyB6YrC+a9C7AKXdrM2IqdL5uoyGxRvK
DnAcGl7bgrVlowRkLf/zh1hvGrGPVNBM2pCszXCIf3So4/FbdjSRqliR4tPq4GO29+PfgdOwvToe
KxT7/Pv8Zl4ck2J5ccVhOfQA1bSkW0LHelm8sFlI9m3/wNBNNVqjRUlyiInjbRO0iyNsW/f4h1c8
K84VZxne1rob/AXsME94VU16PG1XxNZOORasZRGkUk/J1FjQ3pktn9TLctUKgiZdqhHtDqn50s8i
lZ8jrphTUmPVcGUzk+CrdbN62ZZu5sD4+5pfCSCOtX1+TMdy/n0WUKi/AdOIQT20ciOVxu4Akqqr
I2xbOZaXV0jMKAQTFesfaTZ7/aqy26JtLA5I+9h5utUxtdlsgmvOjmovAolekCV9dXZmq2eYRltu
txIY1I1kB9vQgnhYpDbiQjS2972Rn31cwV9KhW2ELxEdGBu+/LiDnzlIDgwzlf5EZeyFTEpNCv0f
2LEnWe7CoJCYk4rQ0uWMBhbozU/TQOVh+T0jAVymCPG8lfafyl2rJAQYhqPmNmF81TIoXHgQjZjU
D8auK2//+jNBFeSzIhsXTvCumXePtTbBmf809Q9iEgCuglL8SHcb13AsLauOIKWiPWG4mOjc+RPm
HBJR1X6hrgFowtIvn+qaisnNCsVGrcycKW+hfRdk7UkLsKJBjAU3Br6nvN5MDkAP2SEoQoXtiF63
Sl1JIYqOpnjvPTFp2bL/oO9y6VaBC5SaKuluO5tjMV3+F7ufiMQLzKtvLlyZzeneOMgu4JLBAsfn
OpfwyB2Zf6V4tYlyO3EcZpMwuDMD8VBXEONHXesy4Bvy6WVivVzKR6m1mkQ39FncPgt2hXEIoChi
Z6NOu+ME2U0F03ssLjeAUirGcSA80YLA0ZWhT8R+AhqfKnIk0S1v3hPAP37hVOkql70S7pKtewLN
V1ly8eHthqhUDulzBBGa7DfgpZWfb7b9BjrGvbWc0MlfNBV303Tb3TxyO3yh6jhTdARTx8pQ/YDc
23rPmu0Ys13hPRPcibdi++m7F5vY/UnmQOP0NvuaRPv81rntXac57sc3lrWoWCQziym1vFRUS0yI
S0lzPM4ZABHptwRug6+9qzG3qOEg+A0shdzyjk11xcnSTs5c8vO8//VxlAYJaF0AJUiKozTBza01
tzRMu0QFmLJFbcsdrE4SZP+X8splFeY+1Uedx5ahqt/ly7uyGg02Zg/szkHX/7GFqpNZGiTF59rh
lU2c5GlpQtsaz/Z7PR1nh9SdLpc/IHTFWvnciHjkgHXrma815dDe5GJI1H89HdqPzMJcEiexSJiI
grpS4znkEQfNfG5pkKb/A1gugfoN5ETau/LEI9ef66SqBaAiDgoXiYNxSU/2Gm5d14sv5w7PkZiC
oBYv0MFza7CM9e26w2YAaPOuP91V8cZdFrBahupuPJBM9mkpL7aT5K6YaJQCMbfPPC4iwMBF7Ag7
4eQ5mF0JywvrzzjmGvmZoG9FT4njcipzdFuyMsfMA4Bka+4+Z4BUEiYvl0g5zoSJTTsVZM6V+tl8
c65YqtmH94HBMTzqIdrQbZeNBEc0IkFL4YXBY7iKU//1cH5eELW5ZdrzuYo6udGSd/BSdROzbMZl
zPtZimWjKLAT0lO68XxBPcrGOvcSbBLSI+ZwCiB8MLmRXSypahzzUSD1IwK3qil6ahYHFtPCNyR9
v6N8EQpMS2CXPZQqQDewX115Y5jBMfcyjSptDCOC5YRsxaqAjBk3t4X/DVDh/bR55h6YUfCenZ70
B956CJP9TSKXhy140iaXs4lRhd6XM6Oki2a+GIOdth7qxDl7gyPzXS0qTuVAdgg+jYNJNDBxe8HW
3JNnb/O7mscUYz+HP56c5m6CeQvmRVNAfkLXFRyjTZg2Tx8a5GbTdhWxBzFsCN1IVQEVrLGNSmPN
pNnObdHloS1n+2+2cj1a8rcwxaVWuyvWtCF2SfvW0nUthwtEzkZE/QX8/Vl8n75h6VB8h4DU1d7x
TKAx79Dc1PHjqH4QpSRDwPmm8QwbZD8Qp/Nl4TcWo0Ho5FfytFwmBKawbXlZTJWrExv5r4JQNgKG
dA3+1zgOLgjIQAcBKaJCNPKx86mxvuQPGXIyZHypGWkD0RgcvFckMU+U3rgV82mOFdyHlAMGI3AB
mw4LfNRSf5rUpqly1+nLn6kfQkd5AkL0oiFIuPHpgheVYn4oBw8nd/KaPV2JBnKnuoa89LhdYxVu
rlgK9WtvNjv2PG0UMHfZ/jgHVDLLyJDSx0h2KV941xz23CrRt0GRjQxvPQwKisLKtZL02EXGcgQ9
qY+JrkTmgAyP6c37A1vVxFAkI5dsgrU1XZlYlwrsSszjNx43FaqppH2tmTu9Hbw7+CBwMTnoodvL
Mg+nsg4LIz1j1SzL3rCRQq3dpN0AT3i+8fkGrqIuMu/Cy0BgND2A6lfmicLFlpMIhd1O3qAXQzCZ
5KUUwg2cA8dJ3dTe2ogskmtVzO6KFeAbSUnr/VsWpG8puI9nCqwUItwuRFk5NKRQarR8WudgGRku
qOFkk+dhElCdi8wob3OIXBIV9o/7eLdB2rSFi+384d4CB4CdaTJRka8Wyrk9sOu4TRi5RsiDJnxe
KdEjRmohlfHW8ZEGmenITEdj6CSpPRc+pgSwCMutt4SUxj0nBB2lH60STuGDOg+wey8hkwhaceg2
hegA/F2d4tYLUprXGd7fFuDYOFXAqiKL5WikyuNKQLrqW2B58JHPregAbI/boyLqv6OPXt3t8S/U
VFKiampvJ7SMKiJXXK7AdHbQnIsmCYsP1FPeXrS68HHWXggx07cjj3ZOjtMKeuiMmgahkCxUUHXQ
Hn6sW/5JEjAuJq5aRoEQpYOKrniIf9X0aSe8TuaKIK5Fkhfh0kQSlPn9U275IDvXIkDmdFiN8f6F
K7Myt0vhUfuGW/e4X8TtroS0VXxGX7c7uHeUUkCFO/sjerDAjE997kTPlpa3ICdNluQ1HfCBBudW
pesh6Vim046EkSHmi+cyACtGYMprJ/XT1fs9cSTAxdOXKgNHv+Cslv75/8i91bE16JEhVTE86rCP
xFfkVaol4lQQ1WGvmhQ4xYV8HY0j2dcYVj7aIm/PvTD/xXRjmHVBG12xW8ez5Sx9jDc3xFtoQNXr
iuhPqdr3edu2N07uDnFNKKi3kmqj91t42cNAQFuqPz33mLi/T8fl3ZeZ5Ue6KslM5zi8/sllSmIk
nWATFP+7y6Af970BfipzGgOw2tB1mXAHIB2KBLui6p8igvYnnMSoNqAHxKtEVjD8z733glkucAAs
w00TDcs3CGtsHMaHIBk8GnqpO6t4cEINdj1EZG1ZaFlZ+XeIFMia13Ox8r4DFzePHZ6mMC7lMdOC
oaCTIo8SduB9xJc4hDp5fd66PMmzB8/dmuMyprIydU1V3GBXw8UWhQu9jLenbK+Y2swIy24LiabY
MmjEk+YtoqeHRreOnuxZpT5maEe1GccwnQLW5QYH5cN9eQzpX0pyXl5w2qdZKXVDOPzg/USffxOC
Y4zP+B/DKxELvHREcQC8/+uLju7hfNZH8m3jjsfzyUAUXg2+ftzAyCS+HU3iuOFGfnhXL/9jz0gE
t+zDp+hCM2qxml/I+m19CbLrN+hy1X3cNFOnZH32bsPrAQ2IwqcUanE+BOngNeaewK0LQa6b/s4U
hTYcUgZRMQWwTa9ggC6IRJnHYDp/z4VujTO02tvPNh1DotiLJLw1gF7sJRh+ACf0HIHPMqm9g05d
WtVeK/L44J7ZAVKK3//r9cyj7bo6Pi3KJz9Yun7pW+ef6+EqH1w9eCnR7N1jycj/9jKAA53S6pOf
5EmG4r2Z8oiNiu5inTu3V3CrrNC/PlFqAbnYhrNFpvaOakxRo7xUhNZcat6I1rs9whT0Jyjcij7f
Rp+splt0z9OvISX3pNDuZBv2tfdS2YiVOwam2PgWjZUH9QM4vR5EgGCL2G+BOWnpKDa8PSSPskLE
IlUC9bMazIqJfEr4y1QVNjRgvX+GZMxU7gu2J9I2Ls1Nrj8tTAmkKwCILzjyE5qet9BeWS4lvI4q
dla5Xrr9oCnX699tIztG52L7QCUY8Xf5jPUuwbqEQTNw4d5oO0dGfXgwzTVl6TRg2clu03IZlizQ
Zz6cwUZeJrf8P6wYqmJAus8jK6WZpMZTuqa1OGVQonI0Z218ktRxfI87MefIPnPoiI0baVI70DI0
L3TeAZ+DmWh/quM+teBfmDCOLRQbua6YV/xUBPYEaxUyGJC5rm6yMoiPKD+OOSmRzg2xCPSDX6Ww
iTv8r7Du3xIu7SWQ8r4d/V+o1yj5yuT+Zsj7/h87+jP5mCMjoFCnXe6qtyXVDr1+2Ut0hv13WhOv
DDYLngrjLLxmT98i9rjISKrpE6KgXMge0nPrsqdN+UDOzsUqtGAIM8q4NjDKX6m5v7BWTm6wvmHN
mnuNV17N7DsTwAuvUWL+Sh2boNICLM3cBvXHI9oKT+Ym+dWu4/AAkuQpI9rxafev/SJbi4OqBlgq
SIkiNXvEBAnNhYnw6AhCbzY3bO7PRR+vpL49ye+6FH2C/KJ/HOuIykAlm0mY/LRyohHu9IkMmhT2
k4bEfYNDO8rUoXFRCSCdyyWKFGEWHh+FObCls7mjmRoWC5UpPjhjch145Kx+aHzd0eDSTnKo7M75
V1UXmF8n+ydZQXCQBIPee9I4DogT3ILifi+qxe3XSs6kXSTiu0wBI6GeLP2dfCIqGyaJdfoayEoR
+A6aHqwcP0gUtJ68WAtj2cBxHgv5Bvh4YjClTL4RGItbHwgs2LxtsX3mJgdQ2Fkjy9JAM4TqST6X
cmUq4KgrxylQUzXeMY5PGBIhWp3uhYypNhP2XpcJMfyWvw1JWkadQlyjPXbbvYxla+imz3p7ZuLP
QcugRgJKfEgQPZ3iLWMsL7bV/KkMzCFSl2usd9I+Vz8WTIkgKlonf6RTSnbsOiGAK8SvG1Kl3Hq7
/JpVvULuS9XFjESdwbfETIw29Rxsg2EYGqQsvvTaSUr0KUV9sVBAAkQK6JRArqz9gDH55ic/Y1Sk
0Xw2nQepUucnbfmPJgDlfKSZhWaPScwlMs7DiP82PJIGISLYbVOZmP95uRSRAXCniyalOO7WkOuW
xTeqGNQjRuLbb3AJKCUIUwcPznUu+3yKSepEh87kziVDTCOAB07BHOm8NWgBSUCEkMzkrQ55evbj
MdLQ8if/CyGJ7JeofXHglz43tgW/xuoe6UAbWZZlSvugGHGJSUEBhh8+PnSuXXPEeHqh3JhLBJKG
CiR/QDjgjqlkZ71hB6C6XGxrhYmBnkaOMnnEPuV2+yx0KmMMlFnIpz+ikRuzCuFb+mxETdGuMmaz
3wVyNIHdN98wgsD6qPufAfHE1gHfoLKhoHAunko4nXUHxPHXHKSirp2eRE3NL0F4fiMKTY/kyKzq
UtdXhUfTSUNaS+8v9e/LVmeH/ow9g85dAPd6Dyd4Exk2n08sB8Ors8CgHiUB2kC4U/lxy/0pD8x7
yAArRsHdNuAKjWgvozQqFKYaipomG2rbuXg19BCaY/oe6KWtKuNOX4a7kjU5b40TQ3uNwzcFcgzi
WppxHtLbjJhNSRvUUyenQp/vohavLhKKci2ZN325w2WsXGZFlhOnaQZ/fCv7CgFBu5ewWceyPYyv
B7l4qxZeC1SYp284b6nvyERriw8PmCFLibjk3mYPp9JhH14V5OB7wESMKCAwhPS7qel327YHsaSe
Y3LzhSa9VQWY0XUPIS/K4qB55lpIWPTj0myd9g5CeazhGk7PfA+KbRMOWFGxie8jrilPfXVK5Yw3
uOybmHydte6s9KLxGgptXT3S4kFVQcdgkuQidT285NU1e/zSEdRbKKxL5QRGpyQSZ0ty777LtNNz
Cs19Hz02ZuRlOsxvMwHE+WvnItTa0dAWX7xpbNOL1TPFBEBppEgbt7L7eBOoTbARyDRzjMi/Oaea
nusrAHpqzT3aY0YAZoRLveqCL+p1Z5Aqy0XgtYMwRnRbtDZd2XerGgzN/dVkEGRUU03K/TkqdYTo
4ZGK6q6eoZCTTPypbsD6EvPAWN7KaFVYOmtwgL0iKg2RMyNOJT481yOPrGECtd5zmruSUtqPFx4S
4euqOFbeF1fHKaJjQKxmJWVSFmxUqGVJF1iUdZ2Rjgyba5dN0WL+VuRVAyv0fnAZbCKug8tk/5Z8
THF2H4zfQl9HZYtI0mQU14lDTdDoGg3ztJ2jDG+2jza0L1y47eezc1Dum/9Rpy1pnXgByTxGZtn3
4pciTH2CaPXKDEQtuWAWn5B1PaUlsozqBRnUrfGZuuCur4YdzhV/02serViT7U2S/V/o4tGutg7u
0x7VBc8s0HzPodI7vwRZWaOP643MRkzuizD1G7kgGVIgs0HrdrKbD0KcSWVV9bcy+yIBq+O9DunF
rAbgKKCvHCLd0z/LQ18epGkOXbTU/HvpwMu/+VE2iy8uKm8GG9S5fOXVv0AX8tFwNehUw995HklM
B3EnQSm7SXArVUgrfUtt4auNLKymEN9A7b7DHIn8Wv8SQi4kK8SRMkF4k4RcbNfqCslCo2+ZXP+O
3a6bRHOWkiMvNyj2QfBhoToN+z6BEjkPU5HOvFfgb4ZBr4OraS17CSkw3pb7aeIEsKomBEak5P2v
VJ8fuElUwlvczwKAgeKyEmeXsRc6oPHYaZG+hzXDON+k7y6FG5itmI5hPQMGZPUU9QAyOPeZ9vOp
TDSbPIwbwp08Z1sxsWaNC28M/lIpd5/u6hU3tPH5wet5mb6KhiUXQH0orc8NTWRYujWX04TpA2nb
ozmws4ZcR2Bxn5OSd+z/5WqUM1I+5N9hYTSuHjK3OY3ey1Zx0MmtJPNzrS1COGWeYTFLecKmvgWa
pofyBYv2jmXP084TOdJgQp8O7B69LFIMCIyrVfhrQFDjsWNkvilFXuJo6jT4A9hAr5nVF07XftXo
ja+Zr3zCQBrAE//E3dIQAltkFUBNjDcUw6QThiJMj377UNqeiJR6JRf3jL7f2Xu3JdPgb473/iR7
9BHos3b1jo1Fb7VN9SXsMcHoodKP/FaDHoJPG5/vhsOp7OVdesIkyC8PuIRi2b/Peq2oQ7fxg8jV
nIUR3//BkmFIQFZrLu2SG4XNOIjU0FkzOuCG7kCSsQ9dq4VwCpx+JAA9WN+pKD3xh+BKrdkrEKR7
U4JSxYPYfflrMhVJcMZB65KCQ75zTwboI9IbCPbLH7l4ooJQ61zxQEImhk4tcbWu1o4N5D0pEdGy
YDtYHJ8Z/LO53DPm4M4jlvKFieu0WGXvad7Jw9ESPNCNjbycDXRle4MQU/GaBt1QU/bQL2ZQO///
opuIBIiJRWDgqsM2BErhj7QQHTm3v8GkDILfidLTWJiTcI/9e9dHOQhqMsnjelc2ph/P9oIZqRMD
rA1CKLNSGXlsUm/mS+dzOgEYIa05sP06O/hU+32YDtJVa6ivVrDE3nlCDz7kkCZ8huWocVHJdzTx
3VRMU4AiD0DQtWuzAUSecONA6OKZZ6KRTk9pWeu9DQHwQ7ZsM1zwN4exbzF4yzFEnQ5IFl8yvA1m
c/yCE30z2jOBSL6ht+J8NIFAov5UvIaCTKxbNvJgBFp9qP9qaopS1zN7Ai4XCelL3VKGHW/TT0in
uD+qj7gEZxETu2lCZsq7I7kKiYwfUX0SapdNPDDenBFO+nYFHKpSWxeMPiIz6s1gvku1JB5w3kKo
cS5suB8QO/c1PhQ0o+dkg0yPPoA4NCZLqlwmbXtVXw2rasjTE5fIiZIZef/vZBfTbF5DmXRS8Frc
wDdAVFUh58a4ub7rPG7bNaSpVgQ97Hqn17XrXGmEbL8vEIQeKN6bdv+0cF+4GTnbAE/tEHGii5OQ
oitnuvncs2+vCsfYj5rQ1JkiGpkYJE+GVPukGaJnxK0J8SlwLqHmgENGroh2+0roRAWd33whHJkf
2CSauQLMXbKe8ArJ4SYfGUNIZnC2j9AUQykUFIsoNqK07mHqaBYZKX6s+OZA/VeEKmL9Y7GG21yo
OwFOyX1nj5qxzXe3344NMS+LRuXvjgd/v0phZ8g0QDGgWugKFGG4tt+rpcnTjHr5ez/znPtpBpIE
s0UWtcLjYbpTzijxaNcfCclLGGjdZcLkNm1svV5tHHTpjeohedDqfz7AuziQV/Dx5hGHLUfFygrb
xJvJeZeuRqoryFHVWeS8hXHpmz0a3wlbFo1bkVjo5FRyqmpolg0YLVnrIphS3eRDvjaWjQk/EQ4F
15305KRU9Ln+bXymtVaYBZRNqe9tmvvzfmJUY+VRn4XykgOVl+wk7j10NokxKUjCxrVynakqyNfl
gIxQTXOtDMuxok+clNIDy0b6+I5kOHqopWEV6+i6bBQV537ily62qv9xnxWeqR0pDg7MlLaCF2ls
R6OUWAJ/L5QKlrNZ0FJg2InSc33j9rjojbWU6FzLc0Gk3VlCho46nqPtcQ1O72CtB1rbOFn1wefj
FrZ/tqAbqW2qA1+r19Z9qGqoOe5/7miNSSkydC+hH8S9My+4eAaxf3rkpsRzMUYur27TRi4GroqK
PRVhpceJ/n5/FPlesLphGYmpe79rJPiLXCGYgbHdv/P6s9dpGlvJ74uKBnlrRm5pCOGG63Xt7rAH
9P48Lx2OeYF4WEkxBbEhBF9puxC8W4qjELGwSPKuQ8h/IRQK/DtpBtgioZV1X7rMxHcscntR0hQH
mAfXmg79I55Y/LgTPk2EsSaOTwFMT2migaZuL/6yVmBLzxl5+qGuSKcTOzfAozbJbY7okbNvdChs
OJTF+6CJF4bqk8IvLTA26EPpmkRLlysDak9UXmR+d/b62CJn/sXiSkOV5Fh7/92oYelIV8vZDCIs
/pMtq63HoBWX6WeoBFALxzgOiYEdxd/6qwsy/eZnO/59JTPeFbfQxFwB8HXP3/PYwwEBX8InwBCc
xciD3G+foJGwI8hBX/QHxYcCwiteVr8W11NKsCbm74N0FMBxNCHCijwpqwuGH59XZ4zLlE41kC6J
J1D6wdRwWVrv78sDbnQhRQv58Ug2uxh17e2Db1VpmFpWOF05cIvOVbLybFlEHYgFmth4S6JLtY1t
CmLOF7c8ghttTIzz5oehTE8Ip0Hve3rAb6q8Qwyi37ecox0eZ8/HWJr3DgoLYbQE6xpiHYUfGnj6
lIAHTZrBomyYOPwzFkowiK0K9U/yNGOVsgPcyZVzrJZry7KdB8n6IERG3TRTXJKDv2/531V8Ac4I
VtLDG5CG4LaIN2NXXqOXbwolhKIvUK0mifjB5bZLIBNc2L81vSs02nBHqeRVXWQOShf8APVKXwSh
BiUOykuNnUbw2iDajCgvt9yY4aa8eWpIrh0J7eX7ovAlueCZLZGolSVWkxqiLkKgAKtpF17geQMY
Fif8XPCgVewm/JL81UFF0aNjseCKWGOPJEI0jehLHVIqsqKpavTOCbU4C6ICayLICarv3KCJ5hrx
82H827+mpN+edN9CWm3/JUb0VOYV2rFi4bzwOwt48jalqEVFFNF66KJ8+Fq6U/pi1amnt5BSsoZ/
vVkJFtk+8mDvSpgXtb+RCECiUB3CzK+5yaMdI6I8vB9H9pM0egwAY1ve1VMVAkjO7uzjMegH8KBR
WZxSN2M5FDVWj3Am42PtS3j6y+Crb0vAtiWwkw40xPUpJvGeZ4+AmX5MPHu57hS6zwsTneYm8y3t
0aWqr/hZhVtCjMyJbvvgQ94VSEhfJWuBhhgGYJQzGMiQB8qWhlROGHCseMaRtu12weujK2BVI1k7
HoBuRSFKb36IM0qnv896VMvYKX+CtKQ2EnjgsqNFaF7jFFMkPmXDlbpMKr//tfF83dhiZnRI6j2z
Z08cxJe2LW0DxZRCtvJLx0gef6CpDraxJOUBei5uJxLSx9r3v9KrH/bPSLOieopaRLhOQcac0wwZ
ZZWNCYvi39lU6BeAULLoOBZddfFvfZFOMn2LNvcuS2jrFCqAnx7RYLc1jkuDeHCiojdy7qE34EiD
k5MJG5Q5WqJMJq9+btr3fpKwnd3yokYlICBYQZzfqk4wi9kkwzcMxr5ibazOQxn186xKpt27rUXq
SvdnCcKJCE6x2je9T+afL9i1cvZKRuxYbmWw2rHRHQuTNe2YX1dY0D72O2aGDfvFyOxGYMgvFeej
8iw6i15qRcdfg9kzj2FjcAYzbURiO6V62Jj/79FrBiX+iEF/2ZoorH1MTsytRcwYBI/cM30uqD7j
ldBSDeZsPtJuFPtkG5eBPewvfRZNaXEPU1VgNWgz2lWOW0SSvZqIWvq/112WIC3K1tOpSv4EN1rz
cb4sZJdmI6P3EQGXcOhfY3mgFvKZDIw9/O8jJcxOEToMgy8j8nDqkR8oHqxurt5MK+jKrZuYjXj5
EMI5nfA9lL1JWK+bsNWeh5TJMEHa+RwhzL/rjdmpXGd//EB1ec5rtx7bV7fG3GlnYYkFa7igN4sI
C3x8Bd17zhQh0es7l1ZSUr/goGgMlzfS+F1kIBCo8N9z+WIoG1YW+KR/i1YgSrd54/cLR0VvC5c8
OmoclYo2j9C3DVYCelPHCAynn+eY/drIdp2/f7Od6U6uwg8ygfESymHw36OnljIV+mHcJV0CbygI
W6sBybyfNdjnxqoPpTnEIujP/mnjZIyI93WJmuy79MtWZHPn495jcCBew3/zYIUrFaxOVddnM/lx
kWVyV6QZPVs3XBRgShw7djVShg2FTkrCKwWvHgaYUMw6dBQftHn0jkIBeSEY+WUKZudDiD1XVB6F
i95YyWkIJU6EX3/TxSVt607sk/XYGireQtChQXuF+cVtn20NrWOWhBWkUGtDl2//yLL201TiOkwl
v3+QDxLUjNxjbi05ueFob5MPAUkOru5Zk1YAaZ3KwK3UivtH6BnZBKzheAhsWc0sBpgwul4M7mWV
EoLN7H5V1Dg0+BgyQJUYp4ZrYt/4fHAv0vM1wP3glKC+bggZmE2jzqUx3dgvmg6owpAtQLxhvWf2
zkrezUuc1nw/1IuVb8NJXsK42N8va2EHc4xHnnqyMOjAKAL+AtHzmYpqWjE8cljmMAUjY5MWUkn9
AFD96UDDPU11FFj+9gBSrvZq0oMhU9AgvNVSy/MbJLRYbYh5to3XrNPJGSnNvRTrEHFTt/pTwjcd
btGxJlp32ss0IhZpCYsRXMv7li5rw7zAAWy8h62LWhOZCCE/bh812Jq0Nt3qJbPZReZ9D6/Aqfbw
AhPmnJ4xbHYSQuyBkvlxmVdMxk27cBZw2G5FcQ8UBdtJeDdXHDuULGR0Ds9me1HyN4fbzsjJioxF
fr6u5idxG86EWJNxsjSJfCpVFY33ndpthP3m4hUj63w4tQnabYhPK8KWsXW8Wvo9zlk3uZQpRrn5
0Pa6x6W4DTlBtvFf+5vcXzIkxnopWZeZNeFctmkSJDBne5pWsxu6e4asLMTR7iTJJNxfsQMIpMIy
wnJ0ovXe+8Ysmeo7Y9SnGfJB9Aj+3OTqt585tD//OF1LEDHXicN8Vti7Deircl4L2b6mPKKs3zhv
RXAyNXSGzlJIbCRgQ3kljBsTKC6SyrJWcCrNdUvVRY+9rbo+IGMPeTs3kMDvZNVaSLzeTkRor12A
fhyi81/TlcpXe3kuBhXib6T6c3JS+eBFZODJZMm/hHLtwJiu+k7vS2jFcJdlGgHj//gl6wiokKkP
rrZC+yDjfj0BmQm5szyeRE5j9Y+2RT4JquU5P45fIRh60SM4LM5OXnDckFKutbtILEwKsyIKRL+8
P5OsvVKd9oXNJex1ugyzlWmLL5/fI53VbtbDtKs23OWF2rnRkn5D2zW3HASsr0LbMFJ57tf4++8U
dDOFBGpARFkAl7QBXLlqYuhWxuQv6GB7SBOTGiP2qRipUjmc7VjUF4Qhki2sdIIUzSxZFSfKTvKa
I5/S7+DqSSmDN0iuAGsDs4Aa69Ho+/O7fYyChuzKMrt080YjdA6P7LQ7E4KAkeSdzhN8B3Og8N5j
Uc9SXxcRBZqRhfZM8HgfQbFDds+6kcH8mgtBMybXprIEOGLWUTEwHiZeB5udu4nVVJYWv86mY6I7
o9PVYs4BR95M92FErAub92ICg0dpyK/hIYNiITqpLVgtDynYpZHKKleT0D+fKDu9klSNL1K6yoX7
P7bW7XL5uECtXybx+4+HqR/yi+G7rp9VE8Ep8+yNXy2bHS09jgI4puVNqJtxWtF1XLLpfTRc3sUq
bvP7efi/f+gCIkfgkNcwLpEIxgW2U3SFL4JjVFlO6Fppe85+JCvD51tRhAiFstKP+wdiR8HMwEA5
Hzqygi0NfgKV5YyNThpoDDHFviyEHJEkDVKEnqfNOvslt8j91A9zWwdHISADRSwQhKp98iSl4Z/s
VIhEDTIOSmhX6n3Khs56j7KBxL3ZC1aeFAm4F35mxInoEWCtHuEBo0uH4UpWJ6Q8xvcudHEetMkd
bw8LtxnCP05dws+z9nkphqYeKBmPG9c37jQm0UrJ31wGgIrpTo/OzCg+20xrX6zr8dLfU/yZM98P
Z8y5vT11+VFcGhy1lrIjKqU8p2iYx933opD97ntjB/iyrezifg7KSv7WnHK9K/vXieW0pe4Y2V2W
Vkv/Gl7ol1CsBsFB7I5V3uGVNpfQhjqq5wqzR5/mLyqhsH5+dwM4N04aXEAqvWEFn4c9xGICMOmb
SCAwPS48g/n6psBQjQQNPnGmUgGadGzx5gCbc0ZxIKAV7kMYHvqYTaIKqkywpRmOP+V8++9gIBBR
m46fsIUAknIHvg6Srns3WzL4LD25AycSvdXH0MVGxBMlJxuaoVqoSogh+RytL0jHesM8BKVbEhtL
F59vrP0BQkjOOo2OIPJPIggrdpfH5wSyArAljc+yeVqwFbclo/lOYruDCSRFSYCjEl+DtWEuMWgG
y0nsaHrZob0o0ni3eRNT9Lj9+yoxkjr6VW1NP1HSxVs1tMVFnkgddyXe/sU6YwooKHKxCsKaXgRO
a9bIpR9RpLPTm0W9B4JtHCzgnpi/wK/NUvXKHtJ5/DRhORMGfluvonc1rEPblq7mbi8eDq2ldgMe
gU7lxyY+UR9WDaO1iUUt+PuSOWiWz4EqwNIdnS1c/XbiXyDSQgMEh1qSPazL8PD3ClhQzR2vjT1g
evS3tbblmEFRs7Y8/c1q7EZ/uDLlrTuvrNmh5ATKLYnp6REXv/GVTJzSGsWfeprCET+zCLrKBqxg
oYkEnQz+4cEb9NthDSN+i5xhbnrNUacl6+CN4mqMBfa8QB2iTps1kGKm6QVIShllsT2R6oImuDfo
xM0XLNsABdu15hUJ/TKROmQ5gXW+TJhgfoA99u8cZ/yKFYihqrJkVehlX9jE2yf0LLq6Wz/xjUxK
/M+1Nb2VMcLi/d+gbJa4RGWWxDz0EJ26DDJ123hljalBgJ9aSSGsNNtOtiXat7NRf89XFnqLt3/s
N3BAFDxUXQzXF4NW3OlXqv6Qke7LfWE349/k4ig6hwTtB9VkbORGzpYtdXtIzTW2q7rV0WBAmhx5
rgksBeu8gBS9STqtu7Eah9p/+FzZaPBHq4iT7fP/apbJVkhD+9dkE6Hi3hHgEWGKs1ehn/GDlOtj
BcabyjEJRwbF+bGTycRdqXzSU/kujeOCqGyYzNl6jQCR9ekQQw/iQYVbpssIf2kQAVJrpWhHQYns
tt1MfkEhd55yQE0704x6RxyL3PfQPlmBs7DAlowUP+IU7Ld3WGUVvr5SKsxPNhKLghXN+9M9EU6p
LTG+MKmV7P/wDD2kh2+0yzpzV1JXFaDVX+vKRAkdF8ujlbC+15dazMvn2lNSxGlzqZ2IOHGUpraY
06nE8f31URuRu1rPoYcb6Y7I1QXMXFzoS97dTyJ3ND/cpNEO1KWBypW2tkMXxPgG9DoSYT7HyU1K
7HlE9mKTS8L68+Ncp5CL+tL18X/cagr1bpszzu5h/+p4OIpYTPoAsCJmPRpYcvuOBpSZ3hRiW3wG
w94N4nIrrLgZRt4y+KrqfrjOhOTHTUmsMsE14N7llpm0rYA9bdY0gVVe0q/5KaQxHnLNjSNBnB6m
8VsSrsZkXWE+cZxMqYHVD/Lwv+NRYxmM23g2UTDClOakx+qL6afagr0kmAn+zThQXK45zgSrF5kX
8zfZ5Hlqai39xtkc5icO9mVvXBSqTTfAyakxUxKu0ot2IcYeduGUZ2V9H5stId3D0n9kiFWb5Sa2
NzTBPzdGTRcZFf9opR9FyId5/K6DM2N3adZdt+/ePgWCvDD87ZfWDy2W1E0g+qh7pdthW06rExGh
2LAc8imzWBXruwwBR0TthjeJjUoOzU1HTWURnc6yvG4khy5wNp1eaF+31u/9RMtkidaMOlr101V2
23hDUUNwVAUw5sMd00+eoNPEZX3qFhh0h0TaiaPIfRO+JGuWbs16GBpNfpKxdODK0iMlc/fEKQhv
jaPBP8jmoRbrxxVlkpDyCJINn9OfYLBXdax7HLo2xV6iSLrYENWsdRgtr6eBDkvu0FMyJRNEkIqV
oy7pPSh8cwn7jQgl2Ik8bMZzlU166aDTEeOFTB7/Zl4Z77TWzSqdq6niUG7pqH6/GE0QiDHeralh
zghQYKNV9BdjV+QZv0eGp3H1bA==
`protect end_protected

