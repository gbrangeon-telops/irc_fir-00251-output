

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ccZ+VLNSpHtEulGuEKVDJLwcsmbh6zDXYYsSS4iGpirAhbXM3BP50jl4c3979n2YR8HDHLXE3QbX
SjQosk5Agw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b11dY0owYoWaWqrEwg1RlK8C89M14CAO8cS5xZSZiTQ60prhJpRDDBFmDC0asd3vpmdy6xip59nG
z+R5fGAzPFXPwL2mdZ9u5u2h5M7NuqWsd4/PSQwIb2Zc37lWRpOZZLKl9FzYzSgF2YNv5/jfYnLz
E/n1SJLECqBWTvKh2d4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NDjOIJz/ezAa2sanfwA4cBF4MUjfAWwRdI3fhKW6WomA0dTdlLUaUk3d7HHvjRwYAFZbgsshlvRP
BFUgnI13aIFlirt9v75NS6zbC9iHo4+u43o4DjI7erTR/V7n1KuL02bh7njjYqFW2TM9DCTV7yyk
HpE/bHTEqhTIUHhN3s21EIF7fvF256QO+AgjOS/tV7UeysPdiXp6gUoJ4fZfor+WTfQVkJeKE9LJ
0zpHP6pDYIRgknpLIxX5LP5O6x+a+epaip1DIHLGwD6CJeBzPxV1RVmuuHt0FXHAwR75O/YbsdQ3
OLvEz7nBONr7GpqlRI7TlZBuj6FdMW9zmU7ONA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
23D8eH9xZzeJ+Ojv/tdSxXVchNNJmk24MJAcRI99YbyO8+bv8JOBxvZhz4Qlt9qTY0ExdOGGGFmU
aQ35HO0+71woQEgUY5FOSxt7Z+X3DhAwHoCaoUzrhIzpo/Vibci8Aq5CktZeDbbFyKqw4AG3L+HI
gLdEde8Lyo1jpmEidTc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MgM0EI48WvFKRy0diETe4cjudrS6vIt7158toM9vdseTaMD0TZIog1UmAGNvdE72kJ9RDo475e8B
1F5FJia14jZNw9OSBZ6rrUB6Tjk4EmqoYQgrN7x0TfSl9ybfwnnJEUbiXZrL/obnsUVUxuBuPHw9
KwRIU7YdWp4ONQdRCD9vZVkexu3R144yonCk7ZQbQol5voGa98xXkFS5wJ9AioaVUGfDCcHlVgYv
dd/x2xkSx6aLm3qbkMFW3ZMl2N86VVdkP+mRZE7JGaPyJ93l/kjtm21dSkDxSaPAALmdawaPAmzL
9Uhkk9hs8yLNZbslAd/6iUfM8JK7nIIDO1E/WQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20464)
`protect data_block
dLOSomOb1oG6D4YlxzYa3QaKvbRaiirXUl2/LAhq3iDprFQt7XHz6kuWjhl8TRGdL8wq9L4MRA8Z
wRrqCFwalhwoAzQb4MuhoTmFlUm4i42dqMgrF9gZHx+LRktFTIRPY/v6lqHhaZmYE/ACLYWRdHXr
CaylkbltF4iKc4+i8rRA29iIReREf+lurL5tas2a/aSxWDMOY4usXwIdjkVukTTPaovbG6NtZKQw
F/g4FnHkjVEatBWmJislwJt44rFNvPEEDA4sClSqLRct9YEWkzGxGrwIC9zlVyXIvwBZW4KvAIIb
Jo47vpzdqtvITRm6/Iubj1eLKHmim32i4GXl0bnCzcShu8dETPv1FeY2W4DZ6NozFiEQ5yxvf64q
/psaDhyUBPbcnYOi98e+ipmjK79SZU28bgNSf8bsX6sOIv5ygR8sOliPn+qufs0cp8nHmv+aF7IV
fOESCP78xgiB8C8OPHd+aclWOpkNK9AIpAErCYj0i8wLv0m+9JeCALpaoudE5cXvmNJCJ6JTs/RG
l+BQ/HZLlBkBOTA1NfhjvnzQqKMSWi1FKBwTaoesN70BGXGNUvrLCJmZDgtZBZ6NiOgQmFFbqV2O
mz3QwNnBt7N6qVHX7CplMegxyRvntgFhtP73iyPUSNSJ2aiMWQgpNTU2CiTjpZi5HB1P8cEueZA0
H6yRzeQ2PFMLwpCY21E5qSxgCZKg1uOoHf6arAYeiLZmRR/X1npb8eOW1FCichV4zUJQROH4zhot
ejKa7N+c25J19HQhzNWicHY8llK/vyIsE/CznI5dx/Q/YYocdgDOMvvsjNycI0tqc9oSFpzlkc3X
5S4c2jRwrfrqv1BBohKGj68SlTX57bRFS3MQkz1BowaV+zYpbHGd6c02Rdm3MHj6paGx1A+Kbiqp
Xbjsr8VpClfi82qGBIQ9mGabNxLmDCQYJRnUfr53c/fbZnJFgTF4s2Fp0nWJeFnG5oM/dvW+DP2E
D4QTqEnGbphejVU8Mlr8eQvXjxNnPkKy8egXrrtt2UASkex8gYDD2lTOKQLZEvGiT8iEoKa4y+Sq
XTVrgZRYECBy7dNY+H0AMSNgXg/5Q9MjNfwEioNWe97jrljxTvu0dG+RpibEiwYtwlcU5WJyIKNt
o1FSdJzWQtBp3S+/7kcc2+YTpetgVB3XXGzXQe220NlkixmsoRLbMfQRZhqVk/kk6ICKNMG/+/Z4
s5kpe8maHpWtOys6W28sy2l2LJS3aBtc7lCxD+86MImgBaF+wzZ0B9SwpStUaqt4lNH6je7eMlIi
9wjvu4yajbBpU1f2fQPLIg4vnG5Y+XiZ62hqBfiBYjQXjEjXyXwDNVinpb6NISDHqvZJVttzeECY
v4WBmmaLieqqxFtpC+dvfLdZr0fEeAMNonDT91vyQoH5XshGJ5i884Sp/dcHcqdrzbbb1OFdE49r
1QMU0dtlqZ8F1vj6oS0Y/S/akJfCfizb/rxowGFLidJWtt1fSa4wAphIoSanP5DSY6UgKVJ3gRt4
QTmkTP0fiEOlES5q7KrY/jZm4LBsPouJrlY7z2Jl7+0VTxTIM3b6LzwM9crEzdm0QVVPOhckBXA5
nyecw+U1Zc76AnGQLau1MrwvggswOHG/5UQM0nY7ZSPteSrts/48/copOrQC8L3WpmYXi7LBp/pM
QUnStwq7XYC81LeV9AbgLgzk+LOYqaIIuMKhiVyL4QFr65TzlAxffx/u0zaLQ1hCNJNCf0xPNXPG
1dI/LKI1SHiEg8LeP3N8CJMZmNVBzN0wWGVHVa9rc88nN70yZLlhcSHooyRtzyst9xx3UEW+6e95
ahZ/Vq1RGBo2sV6algj1E+GmZzGA4q62X1aqCF7Z5mnE1+dDaRQk6WQCfVGuSzZY1eqCWLYo/Umm
3OppPlTtcN+5USPja+kJxndsuzZaIhy7d/SoVgs0bzz/n+S1DlXkJtB2hRdgGq7RonJrquGLhu5v
syeNSESaF7aMjW94Y3OJoarKP+eErD4VfWxvIryCEJPKid24Ok6kFqgR3e69B88gXfM2F75fzQIX
lKQBz5Qs1DzOggbzSFGF4RTqaGogMJk2FYwB36WfUEFZc6LGzV+fr/rtbolhae9peX+Nn0ap40rm
5/5rWmiM+z4XaNexz5n+CKiJ3pWYFLV2HllwapGyzW5fTnwKziOR8HzzSg27LGrxLiJWB03kT52P
yEHHdMIeVEBPbXXHbeoZPxib42YtedZFsiw+oqs89M2mZACME4WM0U30+VUTLxPoHyHV23WELrQ5
H05yEQSBcRMNaPN1aZDJz58SXva69fs8a03MHvhNpEGNHjXxzXQxFclwiv358cQDYl8L/5mPSVaw
kbwTMM1M2WzUfCrNda2u8tG2r8FicZ04U4o+LQGGO+nMfCn9Jw0D2sKUr2wrGuW4Ychm1lY6jTCh
OLLoI/wBG7+ivtlr5iFssNGS+P0latqE+YJ++6LZhZvLZiwHUvqZlDl/c4A9Ps6CKXJvT7j70QOU
W8ZbONivtRkNggwVlfQSnUKzRgJ3qqTQBQ8ADwXW2p/QhqLnKF8M1Nnb1m2Z4/I0MDhv6yIfwCUI
weDdgXOQbLXAdCL6HC5LTCQxqQWUI0RflPbjPc8GEXnk7+cKdT8VtbThotttTuVgdZdg3owr7bkf
aZfInV2nqF90h1NcS+Fih9sCKk1v3smTQUOC86YBjmvhEC8g54BV2B7+RbqKeOz+fcCYDZ/eywdK
7gSnK/Vne9CPWhe2gS2F/Uj2b1o4bagA63oNsbPZpWp2pFb6dh/RQgCWf78gXWW/tLd4k4hawBIL
9zGtyr0uksiGPiRsQbhXak41Cqh+9Bcn0txGvl2LTMSooUjEcV01yV0/jYyc7mVZOvd63H8aZiF4
OZaYPghcPYYlUa52SVQ9gze3IYO4ATAqD3s0gnyPUxi3C37ky4AbbWThBxxKVBt40s4RkjZLapiS
ZuCx1tGjPJ+hG8P14NwuqB6zH6AlX+qd20g95toGj31+VgRNfJaMaY6UCO3pE8U9FtVMARYz78mr
R3/ST/gfmQYTnh7SdTVLo1bQkOZnntMZV5RRqm253mIkiOzf7RO/aK42Qxbpva0bzZ2q1zPtR22T
6eoBpzRhsVPouCGdGQhjeT2MpvYS0/n4Dgzr/VpKB41Dm+79X0/xviafketjUtiNoa4M34OsMSIx
K0VSemTxZiRVlz8tL16Kn2CoNsav7DTZpa5tagFz5+q9WtfADKBpAZMpDzyHpr56MmCHvmD4s6iD
2eS5mKU6n4ZwgiA0mgb+qiwu4lzyxIkheRiXuGgvAk0BkZonYS7YM1Z/u0UrN2AxGvHp66/U1PwD
mRpYP6uW0fz9MyKQgg1qFOW3SIN52vePd7Tut7W0tjcynYylxC1UmbQ/38B1NY/Nf5rPJtahN8yq
kkMnpnIgI/KOf2701l92a++IFE1v9J7amVETL4noTlwcBNH9PYfcAqbBRbd4uUSaniTzKsNaROsa
O7dWtWeb5a/l/ubY/U7cby8AbEIub7Su87P4HXOaIzRt3tLZ1sZDrwpCsG1wIxO1sRHW4WOFCch+
25ajocROPeXiHwW1pnSroay4oMZbtrT6wnclOIl47oU6Vz9d50i+fSn2T7X58sHLBrchpQ/ltbk4
vUjJti+5ogz/0CS+e1bVBJcv65fLrSFL9PP+cR1xj2Wrjvr09lzFwF/b1+Lh0PcmH+pYEdvWH+SR
KLRgOfWS7odaXFnHlCHHuRfWCzpII0jW/uOsyj1DKXjYNbwDKaT2AeQBExGD/9LzSuk3E6luGfaQ
nc97uAXGECeTLY/kPrdD2S1pQPecnExx4WfY607ng1I05S9brGTsCd0h9Udizdwl1+zBTMSA3C+N
ctKvItxSS/EMlfSuzFVquLT+m4VmonVx62mQoucz4+Vo/AT1h188TIFE+4TchjEPuUvBScQRZpqQ
FA4NC9KtrRTO+OBeP/4z1HT9MlpXKai3Xw2p0nga7HLELFsWQ5e30m7+MbTfB20huGL3QcGIYTzq
bbFwjuNsGkIxkVMV5uVHuG/wk+0H7P+JeKSYKr/szkAIYNVYRRVPHu2OcoJeNM36fBGGVnH10X9N
fiIp+UnaR/+y+scGAqTVmxb9rWIX03kAJxqvmFQdSjYkLlT/eeX1LTUyJ6/xCIQYCgF80Vbo3Lmp
PnFYp0zynW6NI6Ys8tndQhAfXLCPMHfh3JqVtVoIDRizM+N1BFcOX6Za+Xu8zoe6B+39vO/GtmLc
ln6/EdyGSC/NQC/jfF2Ajkr80dEd/aD2ob1xAZ38rFX+cM6hDZE8soPaDUUTp5VhN4JbTsSvPIUG
sdcMl5f3B6j5aneLidc078e8bzd7Qzt2Xtu7ok9TcdiRazKFwRgmwf1K6F12bG5PSGAw0sP138p3
o0m5UrcVC3AYRROU+d4Uooe+jA8XzBmb274N+pFMSpx0j7q+eqjZRPlLZp2yWyQzAkOWs6sJ3sOT
kdWoADhirkIxhzirQdeQCXPRzEbpUv0VshPsglpH7AHviblqney4PmwjA8VjFMJqKS5h8HlDwLWp
kRhkmTpA/VTu3hGXudTBQ29SLLYMqEgCT2nXYIwEoEmeEv6cRib1izzzHvyeYn1JIgsvG4CoNB2f
WAFYoDJz3Uzv/Ss6ocY3e8a9Brcwa/KN+6HzibQiFoNjEKsVouIISJOX+eArGKhcb7H8xHjZ5PSD
mD0q+9aXZjDb/yuvESL81ojxHH5BaPLpbT+iZ/jJUj1C9y9M5V5FQf7K7DbPtQCL+ZqE/NbBMXqi
2DRmq4taEZSszEgh1g9fTS/ZBV9/M+7s6D/Mhf952+jIgVK5A54hhFgokp+f1+cnbWshYdPleaj+
YyMf9fuVuJToo4XBGrNfT0JRAz9mmjGqqQHldYWrapSp52ACTKy9Mygda79QOodyCPFpDtnEuqxO
ewdG/hS2EGGWqf5WdBWcCnrdik6q1O0b8PU/O0rdgA6i3w2spAJcqJ7R6ZrEhqn7n1WGNQqHgxgC
jqkZqbHBea0Y83sjD3VpIoCsKkaVkW7C5juLbePk3vW7f15JUAf4djSofdxKlt9HSypdoihj5a4m
a3fE/58nK7ePa2mySCM8Z3SYnuJHXGOII5Rr9WJ8sVDdxkeziiDBv5K6aGxhVwAVlmeMO7O0v6HZ
YVcz9oPj/JiXpJyvQeyGvM4ZI7hb/I1km9u/uXjNHfh88hCU70dp4w8vSS01AEw9vcsNzq28sA1v
UGDwWUauxbJnKvdqUbkhl3HPhG1h0QI76rtFctuM1nGr/P7A2s9MZMN2WHGJA68zs/pkboliY4Za
EVqIMov/ItUTPIA9poBjJooSRr16LcYkOYjIenBY3oe/dZRmfa3/W3kesSNim2n2fN6+H+L2kBOu
ba4GShkuVOt32HnBjSkQLB5CEg3dc8BLT3QNpfhfJxYG1xcDva9RtHFYocU1LSvLkhHxfZAcLS2d
CapA10MPkjvx00fj5qrr3YObXtSykZS7o71g7WcYsJ0u6hI55BaCUjmSsU5VTJonSKgMoeViy/Le
KywTw83l/mkbwu+q7kIMZzQDmM5/HOinlr99i5d1eWw68yKuLpNZwz4mpdsNZDlEGerBjJI+Ojdc
AU/Gx59ef3YDow76NeBYvA/T4zSumGeAa5JyHkD9LTfI7lPrLW0ksAFpXogoKabqhZeV7NcO/2DM
NWyfwoFLlXlQqFMzWCmREy3A3dBbpbBc/Esu5LfLMRETGMgVh6++jHU60Fq9mVNCawxqQe7N0d1R
9Yngzfwln5DBGBcrDwkLAD/Fh7QI/fUAy/ni2Nv9AZyPY57UlzxRDfAPNakN4GJyRCZGcUAGDPWH
ZcZBkRtRG4SD1q5vpohluoD+v/BB+XkfYfI6YZdrcWh8oqI+Fxmf8IlGCSYwZsElyAkg7V3wXTQ+
z511E/D9lzT9ZGfA/nlVy1Uk05pm87vVNsntRNGlvrOdx29ZHkcrUksefOXTKZw3YzK8ALz2S8NW
uVIVqh2OfsrjwMBqYcGZ72eedyHLAJHFFzL1FCRT3TklLtkNep9+tp9I1hap7eWz0og52Whu6mgu
KpFq7lu5IolKJPWY0kAxcnsza/b+4PAvtDGBlGqhwgHxX2K8xsUowGIzwIpdQcgNKpKUcNwc7N5N
BJfjcv90oBgeFY7vZ/Fx8W1FpZrLFJzDKwp+qGb7TfbDioNnAet1Jeq0b628PPQQftsbiXrdWoi5
PUcc8TbgsPIrqBm/y39RcbhWUngOUSx+Wef6/V2tYiBeYsaPLxpXlMpiqbPWpXyckAgXlOFpfr1Y
2Tt65ehnpvDQihE5J/mOeOHIHS+pBUzDxekkdxRlz/eEeOiSN5WTJ03B2IBCNGuZsiOBVeyhhlCy
+zEBmQiteFgQ9Ev3ru1bsSRP/dOZGCCQpYc0luAAPdjeK4G2wZ4UCVGsz7b02P1qZWHmPvvXrlOm
azRzBQVQdfuUrxprSah7xuWlxsBNhY30Offm4IXRlM0h/Fur0Xdub5WXCIBj/QT7KZsfVhjlpOma
xj2uD9WD3KI6+lQYsoroYslBeVKtcBZP6iw1epMR0lLLwPMDAuFoRpYjYDpdHblQNb8WdxKIQslP
ypnpctfgmKgtysXF5ZmtTF2JwaqR83uZEcyE0FDkQ/wrf6UhyNP0RT69f+CFIkNVAgCF1RdRjdVX
Zc8PMJoAWSBQFEwi3yxUNWR7mm+23VhC2lhTI/NDvLJ9r5p/BqgIDRiIVDUh4qt4iDsJqBBQKbol
FcZNdQS2yQILgtYmQn9nDFvxGSReGzRaCLh1oBh9v2Q/DMOn8nOld7jX3R2QVapH3l5owiaJM09A
RPQd5ztcPskyApj2iVchDcmDHMlAUWUojKomcq1LOyrqunI9jJzBn8FAVF1sHOwxJF3AZdB5dJiX
X6oDdLvj3feCDagMOIIOmDGZ4RA/jHXC5XfPqIk4JvVIrvi28EAKwCu+q8dakHd2JgRrik5NMvtX
NBDQKtXeuhGjA5L6vJO0lysJrcJMibdH68dRnH03w9gOYxOsdpducyiV5zbsF9+8VYTI9o5RwFUB
0KF0S8IfNTmDd+Z0Jt60Pk4qeeT0qiPgU9QHDFoJCxHg43/b3PRSoWnQu0ugVhRUJGulMFejK69A
ByDiqhv89byX20+jZOClRfKQWWvTy6d8p5OF+gc6XEzxxUcdBUc/jdsXb8R+SEJUVrGTQzwFWQaP
IwQku9GkMaSv0vIbZjxzmbqvrmD4UwwLOzBjV3kls3TsBcnQJLmeigphZosAKDh2Y7grE/gA8KaI
BW906gKWYkZ0E7y1jOJ4aYKilOP8WNaFzwtZAsZtdRYc6zPFobQupgShBwmqsz8ZAr0vgJ2UECje
UeRI1qOzLTsFuJurKT5ZaGrVy0HShES08YTLl872E/hLrFgMt0FDQ3oEVwG7C5kje18nJxrG9Fmu
i3ZJypS1VhAlVLcLj8/p26z5WsDFW9zcJVQXpxleiqQSnWpXEF9rIdjZ1maojRdmjGsX62/T00ML
dyMXLQSAemsdaTE2cgB1gZcRqVXd5rC8Y1U+HH5fy/7cKrzE1l2yX40Evr9ahXtYwjhDMg3Y/OI9
taLOkzS0eynwe89vshj7xP9wt+jfXoc/T/wvY4FaHe0SekbviBmCZQ0ejBbMP0E9pQlB313rsrwq
jG6ZoIXeoodpNoOTj5QeXsazeiMxEMlhDRiagSrHU3XwlKXmZ9DNP93NFb5goslCrOHhCD5VeUTh
ie9d6/7RGlj3EnHtlUkFXqM4GgpiG/pg2bDa1juCv6qsN45YOZwhGfT+eJMP3F0M5w4At9BJEvhl
TTBHKo5OhxeLNH/xd0GNbHKoN79H/BxUnbtpP2miPIcPVKZXOdqSCFF1Xkyl7zpaQaOxuTl375hE
BFqmvbuRZNXzgYdVkZIM3HmTlEyQ/n20tVvM3Vn3pcqpo9MnzD78/NU1QullbLu5m6BCnEXmWqGr
A/OF4g54OLs48ccEEDwehWwtx16ec0ar+7YNqHUQr9Bol/AULu26u+v0IMYXV8rBJeSENzHcoSUo
moI/0fw/59JyhBzS1UZOwoBohVDk7zu9Y0dp6X2dOmEzJ5V6eEd3VYYaIi1slAcqCvv1eMfyDf1m
8I3PdLe+j2p8tlvb4cIYEK9cRVNfpSBCoOaTIvWmvYZ3y0REgGOUCntqT94yzuAzQeEjUHihEzcQ
D72qF4O/XDrFb+Xm6hoZrDrWdSgyDwS2GAkaMavofqIeD/hcf9zxKi1vt12c+5AZGdrXsH4dgHyo
tMf20YSYGGKvSdSbcCAnGkdp9dlFUgf+gK9jKgX/NSr0ogn9zfm74QO1vqwlAMOPBWLeP5bJt4Py
hdGqEUeI1dTh5iovohLl/DhrHxczItcFf6dJsJq0BEMaNWA21IyTmIV58Bjg15n5gDb68xHFpBmy
OYVNyAx8LmvwY94O6dOeNUCszAwg/mYRY69JD62B5++MJKELO+ohkHOUStyrby2eb98uwpqj5Or9
akba5rmdan75uNJAAGzRcnvMZe2BJ5phLeXGoQKDblJHS7TAjNVcTMkPn014IWDYAPvz2M4s6v7u
f7mEP4d+oCPTHGWtkijKFKMydZQXoLS+1gjP+ZkZnrhxCeEG3xsKg9Oo+RGVYRkCGfCPKmRZAZSu
bTDIwrTYSzbUKpy55d1zA7hALFuwbcNUK6Mtj4Pp1esa04iCOyfN/ivlLgZYtqexc1qURvvv17Co
oNo25F4gWaU9V7ki3ohR6SoSiCqmCokYg1DdjJUKGFTaipXJWBPGH/kEOUdZXsI1ROSwC20yKymK
3ovX6J030zInpYb58m4yPkTnkFNj9Qp9Y4BCU6RPNGQkL/pCrwTQgwC7zC3kh6A/f1M+4Fq44SGz
QK2H4JaiAhvRJCWUze+XmcUwl5SXrIx55eY5b7FYgSGuhyZHKxfjFz+QYFTfqUbos8TN/gYQuDbd
+gUpAhqlKfgiCyiyPNr9O/ZVyv74yB7+cA5cj9Zzs5wvv0rX5HuMugIKODLrhStrCbgJTRjeh0aK
ruEDRKLjd4Q+YF8XfEQ1KktpIOShHy0EjnxlKuihqZPHVsIS8PchGsCrg2cuj3gTdbdxO1uTg9c7
moGoYsPoWkEijDZx8UdJqnjwdeloV4oD6HBr5yekpsh9HyUbx0d85iFXTJOkM45/a14KQxSVcyYo
Ad/UQUPSgh8MZhwu4+6AguKLnkOnSiSOwPtc6j0ra1thQ08VNMzdqVUfzIAWHtRNeWIf8e3AuKwg
mIcKab0u+ybqUrnel1w95uEuz47DVmBo+RUT4CncZ5Mlvv2LL4OJcH0tYlf5H9PDv3jQR4sU6/+n
Pr6JbNacyfJYF1URvpYuHS4p74L2D+C6bKDMCD+WYSIJKWQeXVbJEWCuU8r0tUkYag/pBKDLP8e/
Ce8JXQzMzXOvfjfRraItnzUEFG6tiF1/k+GFADLy3YmXExbt40WEB0t0Wob5FhdX3VQYu2KT7Y4s
bxeeXLNimRKpybihoy5GeHrRu98BhOLSEIVg2Xawk6fOa86zBFvIAUSOBc+TOBwZhvVxsynE4qbQ
VllrkRO3sBeM+vjrKq+HUW3wpPAjqwdiKljiKQNfZumRyzT2IoQZ7DPtKelKnWoLMB5ehJncTpaY
0gMwrNOH8IlycOo/1/OK1HCnMmh3HPL866j2IBjYpnuGOEXJt7FrqcItKW8Z/iqVaI+8iKsoUw6I
7IQ2MPAayQoXIua+FjEm2o92CoclfTlYRXpal9OEsK/0HnHnfsmCh/9FUWxjGeN8f4fudxmWdfX7
uN8vUadZL0QfpDRqMcYHS1CRfw7f1ei6tbGrIUY9aQPuSGg2kj3eKGPpEx4V7t0s5TkQ98XBdm7Z
7+fkBmHJ4yDzM35+89VcAVeRkTNbhy7fPe5OVBjDjky/cFNImlfEzJY8koAYWl1gxe8yjO9Iyr82
SaIdDYUZAWKJLimh7WkEw/FfCR63NSHrrTJ6QPqYm6dU/JZeildMlV+W46X1emrmhWQOMkLIshT2
4+Kmlx0Unm09MO7o2e8vINBE9sAJLJrQWuYppCdDGw1PUQ9wU7eMCjEokOjrpDTZiZgtUZriXjVO
tcfjycfMH34LfIH9ymxMhxVIUYZYx2PGlKwieFS/5YW6KELKq0URsXc6b77dtkFz+xgSHExl1NNW
mLwCdjUfG3EMI4dX8wmvLt8heDf/4Q2+eF0cDeUOLXdhLMq8+w+cXdiq+j6hk34bBbHakqZYzw16
jUQUw2U3RTpfJb/MB4dmwSrfMuYA8sHYvICqQ3cLv/M0SWsMVzanQPipOSJYGWvtegYO22Q0PRR3
Z5lTtL/NM4h4CBwMH6IXZ4EPFKXBvfC6GqqJmcBRhV14uzkbCX+uxLS6LQLMtyWfS9YsosF30Ih4
gyj8rD5PBAskGXc156EhDdAFi81iJOYjjieVLeHiIKBieo90jJA0V6dBxAGHBWPvVljNBRgxzDeU
7H/r+PJR/10sWtLCbQPq4uN8HhPfH/FeIJ03G3IfmjynP17DiY22pdsirBVDGBhtPELeB+kGBnI/
JUdz2vKLE0AfPeX7apKmeJMY3MyfLbftHfuJMgaXECBFvjk+gGqiaOlU3jj2kEFiFuYwUWsFaLDE
GBrzAiC/bkWCxN+wDxbzJPenR44TIFtRGW3eHc8Xm9YXsZ2Vpot9+r682RT2jRiI8safggNNvPiY
jgbgxn7qpy8e1rBw85RA5lkpBjuJnBG0p0kKcur3hzVKsFh7IMtOctTc8lhCwGnCT51Ekrl071tL
QJExHelbT/1OnZpsvNfrkkj2qY1/1Tb68LtGHGIrtN27B/UgO6NqhUrmIWmZ7l1QETqw6gDtqkhZ
SJ2Sd0IYL7olnVEXz2SCIFrHpTnVRxM+gGCeDB0yn7u2mmhTZPtTOeYZ3ozakITJrVTVvF3hPU5M
jQZ4KdxPzUuuOE6D3HqAwocH6X2vnnkFXEdqDLjG4SpTmfrAtSpNf/0o41VEyOI10/bYC5Nh5rG5
D/+dEo9w929RIIlPiNPPi5r/LQavqs5xLxELjLBqsHWHUL9jYhP1kQE//F1R9w2NS39jPaDhPG+b
rLPmQ0ovUYkn7MdoQppU9az4pZwuSZtmAYMphBfQfPCaGbHQL/LJ52pWZ3ijMHfxB2GUiZSZHTC6
KhgZvV+b9kIzIR6PG6tBauSrind3Nu0n0mg4aGCzUWR4N+LIeferexAgT8+rBm+HJINUvafyEvAV
cE7VJoULye+pzeYb0BTVjRldbnU89zbnM+V4RbzcH6sXZkENOu5z0QAZDhGujX0NF11aw8AOiLKg
s8Ly38G19uSOK+c5f6UWfZgyTLmgcY0cvTYpRfGtBsKCQo4hWpaXpG2gaavrPX8QODOnnsNQk9KQ
rZexbLdHkfcawsx0PtiRRS0amrABx8DlJ1OkLdirrPLZLjMv1rAkv6GANgpPvfnABSzeeBPRkNMs
QP70sC8u9XobkWc+QG3pql/grNF8GFdyA6934tvDlHO+QnyyhrGiYAPYW3WP1nxJIYv36/wwi+tA
38mGG+g+mrqTccVcW32AUH6IKnpa4fkLPGoer168YH5uw2jou+r4mtBP2A6l54seyK7POyPUxHSW
+POqGlkn3hbgmfATMOnvyRQ3ENYpbLv6TMs++SWo0PEN9kD7sKZ/xv89i+wEOOQEqedIurAhFnS1
Zsm6pJfE5bjsCFEk9nQjSWxDfMRe1XIEKIt43ZvRNJhcqSnQEwX/YKm2ZFYpGbR30q6FwhZbwkeu
+uON0BrslLx4ot4Pyke1vKFv1BCZPwFAgZkOPaSzFfj2FpKKqWOZvkk4Jk+/kcVoNH/Im2lAJQiF
pyyCXe64d/5N6R4qWV4sy5nLjms8UiviHTgKkFUotVqtuTWdbF8Iy+cwocEr03QZcUfEEbnmCmoG
8HV4FDw8Hp+IVI1LU2jcjSHKYf4LIF0QCLSAMeFMFR4+cEyyLKiFYS8TMxFGqDcVWek/rEobAr4q
0vFkw9nUeWh6BwGfLOG3snab7kANwR5iL4ph7O76Q3Bwt/iKiCWb8VnOqQqFkkAq7ct6w1YVfzkN
d1bKuWVAwmMOmVgG4ETfu7QA1JfiXSjQNC+RPPDS/+p2Lh/1EoqCTdg6VGgf8sFH3MY4/g8Y2etd
p81eEONsK7hvVKuXTDHG7jsnQUJMqWKUbzoOqfnju+o36OWFMJlVhXy2l621KzYUKMAYK3LCWzDu
98Las7t6qBxWRE1HgNZb9y+RvyNUNlltXZ3QZ2uTa/xzfRZ7XsWedcbMR7HZV7LSRW66JMJBtqLP
/7dSq/DMBLi+QeexoUl7ppD4rxPSVN201vZbfjJj/FX2fVxRlM989YgBdhqhwfbA6KlBQOipr+pe
2ZFtncGXcMhPOkpZ6yknEiMeTMRG8z3E5ou5Hr1IOP48TyXDoD81XaK32U1LSyLQ2AKBI6aJL7wh
gciqvsQa35lLL5u61Ao1g7JDNMuLC6luT/0tpt2dL6WaQyZ7730Zn0edZnm8Iu+RiwfIwhnoZA4R
bHxq3QzlxPdznjY1PWsVD7vqPLqoqe1F9loHqD/O3+sI0hQWM8GYmvRbl9JRxpfCVD8IQsFBZxXS
M6sdSTbEd2cOoUhwGNmOFWXiZY8a9NsMJNS4LmGsZaAB3Ob2SFusCEXrwRWSsSLS7dUhSZMGeS+5
jw8ZLcR7seu6XlyTYpIkIE6ltoJmBDayJh/0GJuixVtCuMkJN7+Gdg3lbTAuIbpeEie22XoQkHhU
qrjY4Gp/m2OExie5q8tMxqKPZKDMS9YowuMBJKAERNy2CGtXejtJ96ZeliJJoeST5OgBUSBbM7Bd
Com+0KQHHtCDdJqGly8MAzsYZhA9/VDFj2FFEOt1jQTcozC4jvpeJ+hozjnrGIPIR8qFH9+tPuW6
NcwtDuyZnsL9eOUdP8SszP2YkqxKi311yKgPeDskQFYed16s8ob1KsGQ/Trv7tKfd7MrR2s7sBja
Txnyo352Z19grNUM8WcAESOp3NWRladoMqwwjkUKy6+OyDr+3uTzV6TqinAvi6brEJm3Dutqwjxu
plKfKSzZVZjK7/kEqk/xXQa8A4kOE38jJkv37sixqg4Si60gofHiVinnybIEjFcrljTO32oqdffn
0y17L94HsNML1+lcGExW9Q+qmqKVJHh40Vur/cHZlFw47GznbFSV+Ny+JLgukCDr8AuhycnspoyN
d8l2o9LZ/Ur5EL1o7s4Ba0HibmvAxHlVUWOXwLO/14v3a/tqg0GLDc4lq9xmRuSna4w4Ws0u5Plm
fMOCUf6Y71ikXFWI52QgOKmi08rSN7wZ3n/DyIbPxbEZmP1G158I307pYuR3dQn/F5YZ9n5Nk9zL
ZU/8m5Z+V+Tq9rEPrIvSOrngNTHy3Fldg+ZhXgkAsxOnCTXOQl+kmzAgX5gbiYAsk1zXu9IdsTPG
fC60pcXe8UJOBUERUGDJB+t7pN43As1G2a/n8VGEL7NbOBvrr0D96rldPmZ7HBz4n9lPyb6GoVEs
YwZaD0GubrDxLrrIt5conIpLc070FjaCKwujMUPbySXsX6av8EbLgQiKaZF4opHCPvT2auwtI277
Ui2c8/RKfjmgKTMtLxCFywuRm9YXdA3Ai7Z0FJSye6r5RVVqwryOogCTvapb0tD74MEgWZKfQEoK
K1jeMRiq8CizchLVV4VFqrDYj33DjpXebgVfYDmZ6GAB6NG/NpNFM4xdfBbxu3VXTl9cWXcpBXZG
li0X1pap42POBdQoja3TZdZGO+q9XFW0hz5fKVG653i0sdaeLjjUHgVivbhvzSNolRss0H3qJwPw
TyUJ5Rzgpow5csH5VNAvyVXBj5jiFKKlRKJol4LU2uxa3AW5VaAZMpTKmx4LW6ta1mDJidX0r4z0
eUngfPQ6WB59ZWJYXxbjNsK3Lx8F9Y46/MfZykFLCfQnyAfUcMx93TynnYBZwDcPcyfV8tYbvRZP
VG6qY60HDFmsmchYYTnrUuMcB15AgMfin0kYzUK6wCEVzMpdk0/au6wnu8WIKGza+p4H/s0bVzyJ
7Z5aELfOCE01Lx6drsT8KVzOPSG6NbFp7NP5cqR0z7AVFLkQaMHEPeNoCa37JXjae5Ix2KJH2NJC
2uWvSl2Vyl0IxSyQGt/XPza0WkxapxhNX3EFb8t/A97OGqn6HV8autSP5pj+aEDBVVrEGkCNX8NH
2qBFMqGOutoqPer7dU32uhiHEr7Kl+4yj0o1U/qzb9znp8jeqrqnjrmC0DcZkkpgM791v1bL+dtD
umoZrMWysM2CKTj/zy2d3mlpsoh2WIUPAnEDblzjNsdO7+tX1FRyytLee43Iclq5D9n37btjLuge
UMKpHFq/DQNur8lEc688n4vei8dhhHPdvvPq9GeYYm6S+LrBHIOroHs+q8eon8mIdAD3rf0Wt5JT
NUWLuiNF6skCickDBnw0BtLIXTJNo8yir55BeeCM1Ro0cwzE4mu7mCiHaJHuO1UWfEI2rnl8yub5
9F6oRTYqNrWG9O46a2BHBPPBX2CKIEjM8EeIvbCkc1ZYTkrnRnT6yh+WLIlIKHYUWu5jDJmv26sV
IhJwXNp85rPqv4b3ow0eidK4fD/fDNVAlVPxBsbS3fxM7+QhsXVZj9qe++hNuyS5NgtB6gRf9127
44KPvkaogOkaiJBn8BhwKupzTkFdEcafYCftLoWZ6vtJiOyqOQ1y4+6ULUQLPYSwvr5wl4inAzJx
JO4DepQ3djhGvnDJtWfhqGEykXc8duUX81qg309crduW0nlP+QILFV1WU013lhQoacb2JSXoE3Vs
hDGyiiX4DPwz7sW+omMqEpGaoWYp82zDGeJfMf2pmt5BMN3jX+AVO1OTSIHUAR0pi0CubCTdmn8d
Yf480BZwLrsBja4mlscPEtsZ1J3wl8EE9CWWvkOqZPpZqZYT7trRq8scs2m/qqVRwL1MxcztaBjY
0VmA/7sfrdNaPqxEWzWkMQBDF/aycFI3i8DLhq7Jw9gLzAwaNdu/A4MqoPbFvXZaPx5iYB5qxzzx
zrnXbWqiF5N8RTh9Tuq1BdgYzusvc2JapCytWoAFZ6o/VKYgxRnC5jDo6Ab1MF4Ti+g1oxdIw+5P
sPbRwqNdZ8UxTfuDzlWCM1cJIRFxXwPWGtCb1FnvQORBvtPO5j4t/RGb05XYxXIxB9l/qW5iTwT9
aJJcpf5UdQaBIaPCVWezHM2E0LZi0fP+q3VkpBthaEZBxiMebNYprRSyT83hFJ74J5t2rWyY35Ut
BaqwpbcELIba9PzqA+cbysRYpM0+Fh7JQhyLU8h4tJa8G3HZHqp+MrQHmZJv0zfKSHtVIFPmj3ZA
IYKihVN0EiSvbobedCNEfjR+E50ZtYdbLicucQl/SfgjuHhCxu35OTeQpXqQ2arOJPLVDkAyfh1y
EXXl6Lz7xf+PbrClSF14S+stYqBBltgLexSPIAZN6JOJJMJEUt6uanjcsvp6q3mGZNv/2q5gsnf3
YJ+qCJmcR/X/Qm7DonGK/HK0x3e5hWdjcDtTnt/Y4JTQC2L/TZW+DrPqvl3rITNF9HijDyAzOEmZ
56kNseLfAkw0pFgpVDdaMrEUrTK/J8CcV6gPGPx6ic8gKgJEAIHH2+ggURPpYIdTsLzgEPwEQY64
HcSinSK+IEY+mM7udYblS5o3z3DqEDZA5Po1RvguFpDMhze9omdgeqgPGSkhBZPBfldxfeRgj6va
Cm+6m3w7vjwcrrLkvB3M0VozmvxCDpmv5qh46noRqfGl7x9MbRPOuwGdaCwBQpTcIGrVsCS3/UTU
3rbFPXnd2fiX2+BpSv8w0YaU2gM9JDQHhkfg0BAV3Vke7ht6GTSadOYdvoHPb71MMA8NeCGy6I14
usI2ZgFAelE7AS+HUo3RWcHwcbnxbj8XK5SRjMPyJypENyDNExJfXzgcb/Bq6zG8NWVU5o4ycBJF
gr0tE+1vNnkDTJV5A27MbDW6Ze3QvXlPKCv7IIaTkhYY3Gw4aMIQO5x3QiK52G1EpPS7UPMJ+RZC
YIZTG3MZur5HXritYFVmSXHtBDAWY3Myp01fTOvuPBVkhGbks0K2onjaUFk0Pi7MXE3PSQb7IpMj
opFPgM8tX56UY8UuYpKsrtSf+QRJC2O+uDwKtoHkaMenn9LONYrdlu/BLIFpZ2unQ119qM7EgB9p
8cPlYqYUBJyQymTmtXRzBMhja8sBAH5CY+EXYlC0pGfU0zlr3OV9G8Pzi3MCykTpYzYjeUyJfE5t
ZVqaV8lAgtVWY8GrTA2DvbsjpoyVSDc2VSEjcm0jeaVZTwA+RE8l3iBVHj8nBoEyD5woWamD5K+E
OKn7DBvnxqAzll0XoySJiJk3+ML6V65RxthSIpPTnw8IVjcREJkJseVe6CHJLaZlnQqT8qZWBc7i
Sgq1xxuIVvzcrzhoz2on4CtvlYmW90nBCq7bFcd7Ypl4YfDFjRJvX2bE+vsgDUiZr80HdEuhZf31
RaaL25gIOSlBsjuyrn1rmU+RRurGyWLRp1yLg5pyqshZVfjZHxNNGCmjis2Z745vDilyRGuLCcyT
u5a4jEmgy3//7GDhCI+3nxcC79eolgJmeOoR65wcTAO/uxMMR2NuNe3KxZCz0CcXrobvvn6Fnm0Q
YXbpRnFuAfoDTLpzv9UkIipRYFC1n9X1IwZOXN/vckfOieT/HO7Sq587be3+5mEwei8grR+FVdj0
VJ+Q4ezuCu6qp2aM4kYrZzld1QPO2lzQI09JJicY/IxatEQJmHkOMSUnG3VDDR/8vgfa3BDgLNUp
FyAgezVtE0eQ/LH0qW8osbHPerG37sno8CrkridQD7QXF1bd5cnSimjGnbKLwRaYBlO7GMum3eWA
JX8NbapWVnwy43zMXpzySRo8uCOM7leK1H7bWRRRgh3HmWNSYR7hksPatEa43uIcqu34GMURPMTB
4tLrqMyRCaSqpFNFP9QRLzQOeIkIPE+Li8HVfWCw4W9P6ypXLsPbZGYPLzr42lQJUvsCjjVN0wC6
iAELW3D6nBvFePOphS9hbRTcp8/1pYMxdGNfzUj3rg+h+OGGYPrD+o3+sw1exdzD7IA+2eF/4o7L
0w5GrBahF1ujLx+BCDDZfIRrrXJRSGsehKhhYK4NdNOOuGeHNtn8HOLIhVMueRC0cBTP47Xjh9I0
UN1MYJsZ8rcYHdNbR0JuCc7tXWj69GwQRg962Dulb/NmnirZ1Ka0TMi3xHokwvt+DWo13Q2v62GB
lVZYkTgm3ASonGu6icg16p2AfXRqr4Hlnka3mSFJRYzFtV7z4pg/NNNXXzOmsAdZUI/hVYYhdnBO
w242QZqLm1SEqtzbUWSxwm5kURdebncuFT72QjET3SMz24jZ5jgDTctd7/VB6cxZeYhK3HIR8i7k
EcO5BBlI4Ia2U/w5WW9rwbolzy4/4gS6THIDjw+V+1QRlFv1eeG0P+vV32/9IbmsaZV06U9VyrF+
syhEiV66dxvmpaEygCFd8o/m2VTx7APn2Ha7REX8tWKQ1IjkX09snIN7KvWosQRtSAMc+EJQWxdf
+H6dGmJCbt0mqJGGG3UXI+w4MNXS17aY7nk3Lh5n1XURUrUKOmSbjE/XHCKu2cQ8jNqrhkEOpDmr
J8JWgX69V9qfsBiHtSnHMWSDfpTuz08tH/+VlfQSYV5gZixkrlU7Uws0d5Zw8yW/C3MaOVlkG74t
+sVxnK5BOvldWbnh/DDGZBTWeY1IASiyauBzkoCih09plz6xPdFVn4DC8jBg9SX4KTiYRx7KhoLu
BdO6QH5mAMR/v8FVkBgJKKh4NXihPUneLKBzX4JWXiftwenaZS2O6M+R8KCN8786iQFW+IzQfEk1
9VuyG56iSY7IpoKUn/Rk4WzQlosJ4zqUO68SBDAbOqQNQB2HIyjUvCC+kaJ/cvh9/WKMN8odaupg
mkq26oVGQ4Cwc5ZEcqtInxhE3vaHe2d7efJ+CPAD3W2pcC/2tSahzyxxts6Pm004Ag4LMFB6d1ya
H5PDqjNVRuyR94G7o3Py/f4UcR0UAyj2wM7s0CJ3Fe/I+A7EjFOa4UfLz1peQhpxd6OH6B1a7Sxn
dkzw3yfb9mlRafoF5ASZLlBwfDIjJp5o90zazPZfEAEAMSa6d91v9GebvIpdNjOQfZg7V3uZYeE9
++7cTX+YXT9Sx/1bekohumaZA9vCpiDWjP1VeD0wJh8PrVab6o6lTP3a4I1xHi13WPZ0WaczGPgy
0dRapHpvOTIDPyR2ytECUfAvBrj8il1Rvk75z0HGOTjwLHzuyGASc8a6ekpE5Q8m8NoAlW5FqJoR
axMi+dqVfK27idgQ6fM4WzuT5/v0tBL0OB/Vk6LSsXn7M3NcMG/BaHkaXjUpE0mV6H0ZTjV+PQ5l
f/UPEmDPfq5rnyOnWOfqgn90KnE7+xUi6CAgZXq46f1aCleocBORuxNSiCKYQTtRNcawrwrd7Q5C
+mdqJoSdpFumSq1aO8awLamDdSRtTNTMj19ZO0S1nAeNlT+thT9RkGOIXsjRc6GNebehn649fOxg
gCogVkFo4O89CHGR/OGgjo4bIVxVcaLJnm7DC0pqiKyeu3sIpITHg6WQrOLWnhZbVz5coDPKHJyw
GYAz87S9fl+MqGw668qPLa0B4a9oq8qGzGVqkUV5WcKWmgsv3A6x2afH0F4WiEvxibj/G1sRgU+4
QiZ6oGH169vs2DAaTtWcnUR/LfvyQE9ESXcHLS/Rs268/Xfzk9OADJBWW2k82G4z8i0UB6y2p4Vl
/sxJAaQiGNfwtRO28WdqGRhBIBvA2zALl33mEMGNVhJSIJRFu6/PETMTTDpA0Mr4Br0+yhSA+x42
sUmkDWk998xWNp2ITkUHdkRPc7hkddnyRPxeIZ/8jQcv6zoSZFoDoXikGKQoXTgIRIqrUsdto3uD
VHiUkYrGqVgNcWR4xokfTZMeTkHTNlBZnom3bKvYXO8wutkilv1u9jPiDV2OKyRvpQ2YnkkMHdR5
mbtZb2e4ya38XHoOtZIyYc3sB0duTFQJ87ebTIZ1itUCddWnyejizEIc7xJkjpTiCbO5Wute4HZR
dbCrhX+AKhPKA6xcqKLIC7nGH4w3zNHBzicwMI1pICWMgMVnMIeR9Yu0LvQzmzmH3id6A2g9K3kN
L/CLBaAaNah6WHTdpj/1SDvmBZA1OUWghSQLOsJyDlW1xl2PRBXoEv9id6l0hDtUc1z9387Cfays
9Z/HGrukWk0RSahItWYeJO4/EuUNjFjbn+bK2ramvkY7Etszzs1XfOE6CO+tINwaOPyIyqFh8vIu
RZnBzFnNXoArY+2R+fj/wyc1ZPdHoVqj3eXyL/j4kUoUobNjGowSopyEY+l3Wwix2Do+e33aTdqr
+P7lrmCd/VcI7nWL5LJRiVLcLe3kOcX+GnOpHxyLmM+lfU9beAx7sDoFv2BLkcmG9ROD4Zl2dsCc
ZiE0+yZnuQidVY7Nz2sCAAKz6MiKTAiMVTIQRgwhLKmKx/YyWyDKDd3Iz62NGTm2EUL+muqn1HiN
l7P8cNnRvjm8GukeKn1Yywm/x3cN8qodsc0ebtRm+4DiIV+MMTijMcBIYVj5uIXyx3TApyZvgFdz
+5VClCfSWgoQRBN9xjHxJw1/j19Y6H6tglKiaOYoB8PFt6ig8YZI3kHZUT+3oeFa+eBd01x3MwzI
ZuLxPDXHrcissvMeegc1msF0T4z13VImTnoYNl1geSCyIyFjIfm0/4ej+v1+W1bSoXTwOBUekPvg
zquLuAkRYyXvjbbj889nNmeuTLyYycDbdkduSeXJAngfEmk0WSKpkL/yIHI+r8DfJxKmWyCFJXE3
T0+QB2qVg8F4O72+/ikE7Sd+zscAmIWhd6Q1HUn5YVAGkCIrDnfqizLVcCkHikN/G5pxYJ64cIoF
C2kkAYksnyItwAZt4YYCuyyk1eLgmick1Zl78nBSaRjAK0Je0a1cic476eBoVuWArL8R/1uo8Dra
yOfT6qMCyE7p+dHfsfbWCM0v44FF0xrSqjkONrTNqNS0GcsaIMia8JtSAnIXU2mZkk9SXaG7FmbF
JQagki7uP8/FfeJ5LGHRkCVt+8KGq6HTP+Z3hpFd7mlcts7Nl7SCbsBWcGNNdXRg2sHSFtnTMjMV
sVjXYmeBsKJsexU0LH61KDdaPDUHcg/Vxn4G1NNAV5EqOC83KNgKzd6P9HkUN5FI5izJ5DNOBLU3
D2cukqhcNxz0F41KZ9Mi6T7y4NJaf+DAuFT0v2oRXSMK0XfGRL1Nv4HGOlNVl/aX2+dKea18THN1
Cn8v+y6yX+jKNXSxeLG8t3zg1wIPOsoATUsuoQ3J9kk3zRyUvKxnYiNu0kawYcq5ww1V2W6FQApJ
u0eobIo28a16fmVHnAc5sz8PYWoO+AO+GUPUqoUtPt6GnT1bwQDtssE7BkVWmlCPJBHEqorn8DDh
gnDGKHITYZ0uFn3TnlO4AxFoQ8POzmPAyNl2yaZobdTzAPrCjEGOOWxxTPt2dwo6fG+nP2E4WbOj
8uiFYd+BSC0OGKowS2duWVboqqmHBfhxF9FIPPkLCNp8qzTOgzeLVq6Fz08vgN3Eq+8nHoIHXsdA
VPEq2GCPiQtdSRMktQJynJ/woTViqtvjeiH502NhHtoGYTPdLp9ePYKZM3h2/6UuaQTjVvrsYi8Y
9xahC7NywykZ7AxBEkWl4EswlgyLnEO0HsIJqcypj0EEGDHvP1riz3J+BbByuvvJKiazXFojEvCH
PxRVOLvxwG9v04yQWF5ZTX31eE3Z2pDbcegrhmghE6RUf+4W17nKlWJ5VKasZUVHO2FmrqaqABG/
zpN9OobgYLeX/oTZxCxbyX98rLTeJhx4/1AkbIbnd8uxzcmbaBWuSd7Q5QMNKE5769Rgu8VjFG/Y
xpHKLldQVA4DVTUzzGlJxG8tb9/WoQEik15T7aNnEMdTDrcFXGTFLDykmbRY6puT+4T2iXNtWrx0
gxS2AYDDdEmQBpTFqidIClooHdOnDVx35lZcgPgl5dxhaAQAx5Uv9K4uz9/zIDSjDSKYdSXHq10N
g2vdN7IttvP5O439hJq+WCNvil2v/w8H7RTn098YGwTNIwOhOh4kguThHpwzZlLmHZamfbjUGjOa
eugF4giH/bOB6+eMoVldiJLG4dPKTpBl+8PvmB+a/ijPifTOTVMxcd+2lT0okIT+SzhMXOlLtmjz
VnY+H906c4lR1cF1soyRQjd4PaHyJqX80D0tNtZ7Lce8LfOzdqGqPZdvZR6Swx7wfADqocSzlyJJ
9f/ENO5VcFQy7EIkeh7bwFURcrPxyuSOQeXh7LnCmw1aLBe+3eIF2S5L82FNSB0Z1Vbm+wuwhLio
VbWlsKCM8G9UliDvt1S2cXbgDKw+2mpUM9L6oHSLYZMQEB5XSCNEpJ7CM2KE9XFlO8kzyN2ssH69
d34KSfDExNruFFLz5qawANqu2OvEVgJlpFdbSYBUXTN4Fwf0r69OX9ZI/ZZbiDbfcw29z3Bi9gwr
hKO2Dex//15kqr2duGMD69rM0LTGPz4CzkuiiGCSCkIRUCCTp3afLxER2RUYI4pqaztBkzk5cvfY
L+zjo0/gi1A3P4moCC/1pwY3zNUq6cw7/5zYNxr421iqOOZcdTrGpHkJUjLtjo0cyjo22aEznAdx
2Si+IWK8UMSHXl1h8797+RTrgpf5McyhDzcwKaPf1d+7cA7M9xVeovTgconYbZKEYCKWqAdczCsR
sH/3QGaNkl2lH5IIcgsujykjj/rmI461vuYLBXUF5ahRmt6mYDGW8Tf0TlS97Zb0v1GHaHuql4nv
OHXGuBDqJAJQMHxjgjKOfXrymTraownUzqiCCcRMg2Yhn0Y1v3OLLmZsn39h1h2jTQtlAXv6s6fj
wnqYdIaWgMgosbH5oUR/drFnAUJYZHug3fchbIUXPYC4jo978TNYrMcGhh2ZqciinIr+UthNjECq
tSfTGeGVGg3/2Gir4a71dKFFJj2sOXb+jXf+yYNfGANnlJpkN/3XzkR7WaDaDzyOZZTkNpQF8WBn
4lljopZca8beFE/fzdJwGnwxFqWKg9gNrwMS8fzK1WD54wFsh9op+7fdlFQDALWoIqmiN6bpaj31
h3HC+8iwNYD4dm/fU7OYysOFb9CSM5srJmSbp1BQDA6kdhaUOv9HRsQJ0ycWENo+tasnhxl+6fw3
k17Svf+RczYH/fWZxk1HiMCUpzBa95QsxVtrhQM84d8nLBS0YBYkvAoM5AIHAT0HkDphGH3PVxZ/
Q1p6znjbTwMi28IbrnocgvTJVILQIwA2Ay5s2sE4dsl1+o27qT+g5iSq7bUe/EmsMOdwcqsmHgmL
0aPQnFXeYNvGmXDh2r1/wMeKxPmE6ckicCOCHV2LQ+tyOHqBCGXzSC0P6ftoW1sZUef74FZbEonz
GwvNYYBaBrpBKP+ahy9hs+4NAnFE4fJQogW7WPmWxqi4wsTCo6S6TT6khFdjLF3b2OkOd8hONhc9
MUaxRMm0CbR9HSSMDllyHsuc8DCowaeSsVjdw9DXVed7Ka/k6xoGAfHq9r3S3YapSsMNm7RTbEz+
sd65UsSiCTS72xgWK4XROOdufBfZtQ2GTYoVFLQKRw+HpmQgnKUs7cSnx20QpZdzC3EyLVKvY9tD
4K3q/ZSBSYPLm2a6/pv14nuEqMyBqz4OxpzjBOFz7f5RrBUiVCFovmsGEl61Cukw1waBJtM3OKeM
tIE/PUjx/bvYzfIHt6rq0WiBmwVk9hl5lSwSjqVkASggI0ouoiPi7u6ekVAc8ypCIkYpZTh1eurl
qqFcdINgH3JiAAS6jt0oJiMUyxywEZ9R3e0O3fEavoMsBlBLds4DKQX+YBV0/n1+uA0gKHPC8mAV
3c+2SYXiJ2RK+2fz/paqQuZp79tiCHri+2pitIFu835NGtDhbsadPzZopeV2RSO5Fb+j/GHE8lEA
Oix5L3VvfQflxCiVqD70qm5Bu/ldcgV7woPxM/W3XZdVGkaUpLzL0E0pAlkNYFd8MCbdjsEA6zu0
TSlEyx61yTQjQ3tFJLliHMrMnLp4L5zUPTOUVELPHvbmeY3yJ/8neTb3ticmG2aON8PHt02ASjML
GndfSBkP5Jzx7Bn5NpzuLbj61hp98tUaJcQ0TJrDVhxLhAzERl5sKygRTSVWnlVjc3V1lNcLGc+J
PnJp4FERvtw4EbDMUIbUwYlPmtopUj6uj7mXKLnx0WLi+FQJ9XhiJk6fomgwAeNKdKjk4CHUaH6x
OsjBm8oyAABQOhabeLauCQKcCMN50829XfVYT///k3SkStWBLrjy/e/2tZXxtHttA0XOZV5CEO4Z
ZNhKl9N68qyR4/JcnqkjYo18DCY6QbYeyiKwNSSxnWPKfT/iQsYnOPunZ9T27LU6h5yTgd5MFkyF
DXcEx/gFFtlutG0AEuULNrINP9fEvww7QhO6NDzWFB6Hf0fMlls7FpaQGDu54Y1psmGqoo7OtLer
v6WJZ2X2V+W8GdxgE42ecJnZteAc7220BlzoBBwY7Ego/HzTk7QqofQOlM5n2mIIzvIM2PYzyWl1
vwVe0PuY13Df9MxquR/LQThP4sy7EK0omzrBsXISpmpiaToRHQ5138SSFl3y9KTKmt4Qm4vQEnww
+l1QffZ9Fd6x6QJqOvhmTj+7LNotz/8hThEcF95bfz6rmkIDhWONVo4eNxNSyOQmfzra/2rGEh1E
HMoe8gkt7El/Wg6hBsTUfzAMuYWIvR+VsK8cMC/K5sjBPHCqYIjLt7oyjSeqdifMpDW63G0ev4kN
8K4gBRx0+hPd9Vf35Y/zi0WBw0edQO6awXXCEjfBb6Ut4Z/ApqVpKyfK2KsHN3slzTC27lesDDUa
YqAqfhODGjYA0Kzml9VwddH8dtp+wHfXxeYeAmnfySqYjXZDb9ssoxYOBoPavDHcxOeIHUWrV537
tNblsb3eJX0T2nCKTLKz2BNFinrqWNRn+EuvLie0V2973goRYMr/K1l6xO95oGO/NjPY00P9d4z5
K4tSTB4SsRFedQxLb19bO981Lqxh2fp4EIu4w8nEGRUq0vGkG/R8U2DE09Z4t2I4boWrbleIQmmP
DrlT+nFJntU0FPhk7OLCNIevKrMMssKgm+p9+Dz8HKA1nX4CjETGmRIDKQ1w46mEx7dJV0I6KWcB
4aLgfGMS0zTCcOYKOhwLnpcOmm8OXl6YdgtXIToHdaOsDSn/4CSkfgzuKXvxSNug4AEv62y+U/QS
p3p6A/OKqRrDaDLFKklS2L3hhdxqNt2kmTTCtCzP0zrBD8Ndzd0ggPowb156qVC+XnOAn1EObPG/
LEaNDTk78/cvHvtn4RapBmGIiotNJq9ToRCxF4+OuHFw+ZDAtbiuzWPCEQSTwFlKlFXhrH6qk6Ga
BYntOG+1dWkJARJtZ/pAGO4glSgIG4Ewy3kWWDfKBd5WKHrLPPNBCWj3B+c2Spln2UWI5E8WIf2m
ctEftSx7ZfZlgu+SnIQFe4wywiG4Ixgn8lIsXUUHevopMINE0sRHjCgGv6Au+9kXz1wMeWiT21dm
ndb2midVyqlxUeul7qVwAlB8BYD2LjF6tIIoc2B3nO2PvywqxN3BjqRuC8GCT6pWAzi6VBcEoeJ/
/dRg+YyiCvg3x3klNneR1H//WQ9yj3FbgwCYbnDXQ+60Jup1Ym+2YpQ6PPHW1ckaiPZfJ85042mi
sCb9T+FgxIXXtv9EE8ltEEsR1Rf31IBxj+c+5zD2zsv5sZLjzmAXpcdeTimMB4kPQHfe1/gKvDaT
IoYvjRPopdZsLhuZ33lRiVlEfs7OQFmV5gRwzd0n+DQrazrUfOnefdYzwXSygxm5Ubjia3C3zM/v
Tb5fBEh0W1D/tFshMmLzbmjz8zHJw/kwBa25vfP1xT2dxUZVa6v1CJkyVRPpIY4DMYWwMvgXAIcG
4h8xRe2hbKKW8eRWAvZSHh7JQz+oKSrnkGrA8LbF+GbNHxWQygBilw4sFbo4NpKc/JdSCjVcih73
frsafyRXsRpuOlmluShXQazVhW5euVlyqAyYMLLqFOkJWp+vtH4J7mlLoMBah4ViTYNUNQUyYg+v
M2GYWQCHo9l4fSJbdAnYQnF75qeNkqC14lKAebeWWgPBpBtnTB40ohBUxNUbJ2fmtycvyX+9QRyi
nNT867ewegZ+U3ggzFhTjGcT1p0qerHvgpJ1JH81epscJ5IrjG13WJnYZVtlyfCFO6lrzc2JGuym
jL4ls+kJIJenaZFPbwTSUvUJ+lB6/sHYcmwG/Hn52NEHwiDtfJF0loGmUtvIDesNR3L7mab64R4Q
IZZxhnx9n5u0EguzYN95QxhWV8Z4nGuKFXq2amHViAtNNRmun5+Xorl5gaBPfzHDX0df3CcZE1+9
6SRDBAFzOQW3ogSt2yezbjStNunJ2VVZy31Ckv07ofM7xUl5Sv1yRGHYV326UvdoDFAXuCJgwuIw
0G7PvvQtqFPa8osQDBwTN0zyBSTUmrcLKJ1ybM6sw1jvwjVNKRYBLdh5L5shpNCodUren6qEBTtj
3fSgv24FhgapPxjFYaUpJP7T6/DuG7zY9r0nvpovZr6rQ9z2W7GddSYfjMeeKvqcssG4DV+5ROEo
ew49LvH+Wv/Mn8byJyy38/ffGcHf8IQBlWT+hwBI/eTy/l5QLrn94cDWEeBLV3UZucAwljRI0x4b
VVRL+3MiCbfvIkZAUUvgw7q0tx7l7XMNWSeRO1QU2RkyRw6wkg17Na5ACsgtEWXHdz1VEdmk0swi
jgb6/utoYiqMwT862zEecaDc8UbvRJgb/zqGi6pb+1wKRhG64H70qGOy7zEaIvwJmYr6qaVdZkCt
s4bgKGDc2wg5QvGdjG0z6U5Yx2hpRb0KK93V0tkG+OLzmElkgf5vSP/UV418PEZD2ug760q9fKMl
p7e6x0AtyfXd2u0ANXaw4VnVfgWzPBn5/S1ylEzW1azhO7DXsUcC5PK0utqbIOox/Jatbihxv3Yk
KvrFqXHb1BOxmKaTXBlIBq8SQvG9UT5uxGXLxxjCkyIJ49CFVSvtne/X4v9cHH9veOeDJzhglslT
lbSp9oLdKkySo1aSFgVqZPD3IWk07ERPUrNStvbAhmHWA20rfK4DVjOFgdZmNe+bTU1hB9/lgNBl
byc4XJAqcVU/HsAoFcjH7EuKKSp+LofD/S3iGg+BWiGcHuUhOOlF4kKTgvTgNtz8JZNtD76+n5qS
ad3CwNlMKbQYTIPTR6N/uXV7BRjmVNgKinoQzhDonk0JiXvupJXOUSWQ/7rRusZTY/kWRDF76FkW
g/etF+58AhV1F9T54MMAxAV1bFOz33EJ6K7ZzuGbnLkvF7ttDGP+M5jQOFmDeCW23x0uxOA6w7Yj
qDxUXeq6watyaKPkUzfO69Yk/Y6dm2oNVMi/G2E5UPX7FgeNDtwlPEXopUW68o1edDMYOWRm42m5
LpCKqqP2tGZIA+MamaYZauh4iV5DFdr2VKuZPOf3ET7ztlaHUch6s86h5OA+zq59UsxNgaU7KTdt
tlaLGW+B72uknaHBM83xdVBSuPJKm2xsX4hR3f2+oJIM4Rnn3R4SXgEzLpZH5H4eqO+8Wyv8JKsV
eHLQ/SdFoq1rNVFKiiC+YmQzQwouai4hi1hklxLIB7j1PBZHfF3d0a+8JssJwHyg/PhOsmt8/XuO
eeW7G8EL1g8dIfhRLUpZ5HUM/U9MBkAIHq3MyAVojBoVjIXoHzStt2NGwQrX3KY3QngyDhnh64KS
uu6Q3By8y0OlKar5r9M3brkAWRSFJb7TGoyiu0Sxng9tcuCWG7u9HMWU3cPaN6j40NDgphIu+/m5
xOZwYS0BDpTjTr1EiWeWlCcAxVv6ZLonuRg1XagYUM+NQtsXrLYKKDjza9iewkdxgzFY9NJuEjIK
E4KGrnSs6scJ8enQ0XSvBP8FGN8+F8Lvx3sVhwoVkw7HhSF8E4Rn3a1r2WUYGzmAIcHScoK6oAVs
xAknb8lBObd539bu7uO9xB/YMWmZ3xeAAX4+GKmafgyCpGmpLZeqNRQ/yBYJfolzYApPcIDKuYla
N1WkGLPQBBRO9s9wo/Ot+LEwQJaej2e2n9FSuYSJwO4aVhUPrtBn+J3od4gmMzkQW/2HvTsW38nT
STVQaHiw+sNbeBP8Oqh/bzwrfTV+AgA5Do8kYfSKXHdf3+kwTZXCXalXadmaEX1vDHtKJKoQWDsd
Fpiv4h5xuHt+HBP5naKs+RN+3s3BCCwzj7m/DvE0SKMDtLWG09vySDS5CJTtx4yKraAQRHNPq7tR
2w==
`protect end_protected

