

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ccZ+VLNSpHtEulGuEKVDJLwcsmbh6zDXYYsSS4iGpirAhbXM3BP50jl4c3979n2YR8HDHLXE3QbX
SjQosk5Agw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b11dY0owYoWaWqrEwg1RlK8C89M14CAO8cS5xZSZiTQ60prhJpRDDBFmDC0asd3vpmdy6xip59nG
z+R5fGAzPFXPwL2mdZ9u5u2h5M7NuqWsd4/PSQwIb2Zc37lWRpOZZLKl9FzYzSgF2YNv5/jfYnLz
E/n1SJLECqBWTvKh2d4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NDjOIJz/ezAa2sanfwA4cBF4MUjfAWwRdI3fhKW6WomA0dTdlLUaUk3d7HHvjRwYAFZbgsshlvRP
BFUgnI13aIFlirt9v75NS6zbC9iHo4+u43o4DjI7erTR/V7n1KuL02bh7njjYqFW2TM9DCTV7yyk
HpE/bHTEqhTIUHhN3s21EIF7fvF256QO+AgjOS/tV7UeysPdiXp6gUoJ4fZfor+WTfQVkJeKE9LJ
0zpHP6pDYIRgknpLIxX5LP5O6x+a+epaip1DIHLGwD6CJeBzPxV1RVmuuHt0FXHAwR75O/YbsdQ3
OLvEz7nBONr7GpqlRI7TlZBuj6FdMW9zmU7ONA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
23D8eH9xZzeJ+Ojv/tdSxXVchNNJmk24MJAcRI99YbyO8+bv8JOBxvZhz4Qlt9qTY0ExdOGGGFmU
aQ35HO0+71woQEgUY5FOSxt7Z+X3DhAwHoCaoUzrhIzpo/Vibci8Aq5CktZeDbbFyKqw4AG3L+HI
gLdEde8Lyo1jpmEidTc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MgM0EI48WvFKRy0diETe4cjudrS6vIt7158toM9vdseTaMD0TZIog1UmAGNvdE72kJ9RDo475e8B
1F5FJia14jZNw9OSBZ6rrUB6Tjk4EmqoYQgrN7x0TfSl9ybfwnnJEUbiXZrL/obnsUVUxuBuPHw9
KwRIU7YdWp4ONQdRCD9vZVkexu3R144yonCk7ZQbQol5voGa98xXkFS5wJ9AioaVUGfDCcHlVgYv
dd/x2xkSx6aLm3qbkMFW3ZMl2N86VVdkP+mRZE7JGaPyJ93l/kjtm21dSkDxSaPAALmdawaPAmzL
9Uhkk9hs8yLNZbslAd/6iUfM8JK7nIIDO1E/WQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20464)
`protect data_block
Ctdn4hGe0WPfhQ/UKGCa3PlStrDhNOBHqQkf/3uaXIb+ZA/WJO7T9Fv59TyYueayuGLxODvAo5rE
hv6rBiTspoQc1H8aIbkOUfVArI0DzkXbf8u4/q8zz/ex1SX2j1t22kiaTX1No8boesVSCuYNRRPa
h5toInGNxX33Dc4hSpbaOntXP6VCNkHPadA0pXd4mESqgRJpAOa6ZKOdtHapA9s2Mm5MpUY+YNva
4LC3JFhxKP7DNnsaSEWI5eKtcCFek5vso1AARAeQjxITQ2qWvx+8efBpmiSKlsJQ+5cSTHGlSlxO
6u23A/r2ITzU96ukPZa9H0bxiON1jgAgzkG75Yg+NnthorSlv2zI7f2C3K/ghJkxToNlToyZI8fD
aPs9M5tYy/N3fKASGc9xUp+wCe1sRPqhYWju/lwF1azjw1/rXP2/VHATQX8W0jqQbJNehsy2ToSp
UhunnPgAyzexxR0SacI6z5IHd5jj0z13yoARuZYtDkm+k6AAd77Ay3tg3gbT1hDyywG3nadJ8Na+
cDtkDK41SNLs1z5OubrVbJoM8puKTmSrJ25uLJJOcEwdFs5nbb4KzCoZt6PaXFAvQAUR6F7Tkc0E
HL9OJAJ2o8tVmIQHQHM6d/x73O9/DSMas7RFZuftnRD/eL+Zzetgw1ChwpI3HSp8eei0LxDXxxG/
uE4GUKf7E1OzyjSOh0cPbzpZ67WnDLvNCZ9l/FTHYCw3PwJBum/GMx6QHOT0lcYfDJtcL8c5hjm+
UE+5P8zT4keM3CxHjuguoezD+AXxuhihfgOb+lqGTLcYvqheNZSlQxokIyZTY+o/NW55RCZA9P4W
i0MqgFT5h2ogaF6cuQGBWmCJT/cIBFdkZyMtPIRevdzecGsAxvMzPIlxx8HKhXPEk4mFab/z0htG
3FTWvr1UUnfxjeC7vl9JZ1eqkk8IYeFTqrBkrFTdZ8akvWrZ5lsBtM6YhPUd4XBWMPAL6k2HvY++
ZdosoNeCxNtkGT8deAqmJYz6/hEVJYdFPb47S0LV49Jk8dZT3Mw3TdcCXyPmx+7VZscq0vVhkva+
k+OmyKo3hxZ5/V8tri/ZnahYlQyhPuX1FEZbi9ISVfsIAVjJcxQW4bhMeR30bwkOQbnQ5BTn8AZT
e4/jpN1XcaVzNq/KQRr0O1Xoi/XfIbJEx6j/FOJysHtjD8TNYloK6nXjrkmdOlzl5O/E4PVP7Xh0
w+gEmDGAAqyv8+6IJ5YrD6MZeyj5+xc7G0U2AHNbvIfHl9EG6ZZ43gGJiiKSxp42hvIj9LzJs/W2
s3jT6CcuKtC9FJBmHU9ceH7PT/uo4TEUMEo1PdDCM7ZbmAauyCHHJfce0pdVNlxCcSX+fjqL8CNu
l1R/5auroIAPZZWcDSXe3A2YHU+/XFCP+iTi6Xg8uVdO2LMDkSbu52SlzK+iLOoVQTAYQUiBY0oo
+2WqqGoB7xHNlMKbDbFeLcivBk1CY+E0LbrKqxz8ByZQSJpBWe8YDq1CjytoFn3YdYZK9pUggXxT
hRJiyxs0xOyO2N66JedDS7bKvNNrmCRg5g7RsjVUFeHvlGMCx0tpepLsWUknzaNvCGc7580oqDPQ
8j3QksCAH3v6QRvXJj4ue3eb0EMz+7de+zTU3AOZMHbR4ZTWZrlhXZE/xV7uGIrSDXt6vjSPJPH8
di/UAvVoIz9AxkKGxoKzuLHiVhN3PeREuRbWuNyv2deKi0aHTE9/PL15MAT/jsA0W57En/t2wiIx
qEFCN44HSwLI9gt0hqlktIZvepfE5mO8Hhu/bq1g5yu8ZLCStSlpBgf5dOZX0bVa3RJ/sxN4WUvZ
P6Ce7o9Ch7UeEK+teBFKMT6TGU2K/lUq+s1Nqz0FO+n2WDF+qBFAOa0KJ/QlvqAyTMpFCs7AGg1R
RriPdfNaPCrzzxY7BgEMThRfdnKPh1NvYAGnIGeIHr+GLWAQROsGBDWa77gagAGtbuRJ0/I1peeW
FyyQHC2vIjpKgtFEbUNCgY5HSOKE+CliAqFDpSHV1VQ1YyRPuQbENcL6EV6+QXD0mkB3AZhlYn4j
d4LGe9jcEUXgdWg3Udc2p4unolcuQCFPoFNPeeDP0RCwHrn4ZsBNrze1VZDLY7wNZyMgEzCwzfbK
ZcyxHPeVS3+2ta8NAKGuV9wzanj1ofXjPMRj9lq9/i2NTgQ5UWhDvgz92yRC9KDXx3FrMyH8kGp9
fDMs/S4acdTAYdXqH/egyaRRIBruoLPsvMs7Z1InB23PqBWLnvPBDFX6L09FC9OI0t2uBj2WXg7b
/nYH8DWeiuzYfvkAED6jZHl9gaqTNo9+zDoqYWvSVqtBzNnPnl+LSA/CYgJO8ZtSBxRAbUyp9E/Y
T2LUL/L+kGbc1k2WjksnKUBXM7yMTy6bgFKGzYhhmexmcz5c8x+Onlj6pw5iX8Iwmusqev0bs3em
9/FeWG9i7VIe7r6/uMhwNhne9nO4UEXVYdYnSUctbArY88SVllUJphIG0WXTGhOUISM3UKG2pa3/
UzgLu2d+f9ExPoL9aD5I5ejOMSZPzrIgPDFN+D7bATLQVrtG/ITLYjp1uD8JvRR4USeVyZsQ2ALs
H+AlFfL7Y0MAKDvlojS/gECS2USoMCC4KpP7DWhDxgpiPubjO+vLxO6vdF2c+DChMf1Gx6b2fcvC
hRYoDwmveol7O9m/8fEjvFlfgQ+nHnuqts6MHUzpe0XN9JC3mGr/qb27L+S9czCwnRHmZWnP3//O
MWbKGB6nvhf7VJd/WtcmRLPON0RsbDRNQtoZkxp/HWCw3GsFZHZFwZriPBgGiQ09RAo5o5+BIQOL
5hJ+ynGLOCQYt2ikao1R4KVSwO0QeR7Q5RVvp+93nuCWv3nlN92mjvX5mQs6fJQ6VlRGpQRMJj8b
99B4Qyl7UbKZxHWHB26FSxSmJzVl0jghpQtqlxVkks4JbdbDSc3MDJoqyl8D5bfunKQA60PgTGKU
G18UR43jUNkJk0JQ3G5qKl3RSXo0Fij1qpVkXHpZ1vuFBkaqTIdEiOPyOJISM4bcDEl929104wTv
ovxPHqeUGTBRf4D6RRlcpI9JdxOFmSt8yLOmelRZ0d8M6QbyaO/R13mZl5bsX1/7+cAHiccaW6FA
dx4aQQ0Tm//5nuAQ2CFB+2c/V7JfqW+dDrIe8qjBr/kk9splAjLlWJM8EvhFIRkNtbj1AXfQmLq4
spvSmJU788lZm45M6WkZy9vwAhYcDx5lJ/8bGWqXjQh/oZaj+xrjjFr9D9s+gRw2B71Y28RaI1Xg
T3lVw8mr82VbvRz1G9LXqYtQBgdPGW6heouYIwN9/BULlaUHav1lLTm1w+v7LhnH6IDm+EcEOjUF
q7CknkyL4UNp1TVYiAWDEqVcIqS38hP0myDkbySD2f45DbypeKFv06IY1/M0J5R3fmZrEdFbC+8d
Yhl/PJx29e3iuPAxqRBS0ftJEKKlR2x7TEpctgp0L+rBYLolCv4z+dOUuW6bjAbzDg1Ty9+teK2J
KnY1PUIuaqLNelU/MduyjZw4hy9xBRyyTWvILnB5vpz367YjxoeSC92NILEtcJGKmn7Y5uXIhbXW
XQJZ/2mInXAtAa/S6M1cfX4N+1Coo8iQQTi/xIwceNEuiIROBtNwYrzor567w+22//5xUlMcBQd+
sHJBYEbhFUtOFDRMs/tSfB8UdEOlwBAg7QvLt/DxFPuaN6b+c9vvlyxAfql4YJbC3t/FeEca2kug
57RwknhcjfOlFeYybMSlpl8uJDqo+qx8KHSt/6+X0t4IAUIM4H4zsrSlV5rJ8cCV31k5HUQwVfbo
tcMZDNkPSnqt8nxU8EniJriKXOTxpQ5VmhlQFb9Peo6SVTO2LQKsRNPSeOiE6PLmtZyoNmIPJ2g9
C2qv6zFAHWTf4qfSqB1CDVf7CYyInQMaRdR0HfYpbpG9wgSEBG4JgxrSErZkB2gAjeRQsoeIgeYT
A3xjLa3kykkn5KwqqRPmqU8TfuA5LhpOFgDvbW+FSploqYPGHvCGy3v4kN38Xb6g3AHDiElm0+5e
vvKfoBVQOcmpWU+Ox/rdycA+52c70tVTWInTluvQPP9lLc7khAOJGpkcPgY/+ivuHygNIoVaTT+o
hY9SZBuBR2MrFJcx4c1m8XYSFfSYsb0xplpWx3re+Sua9yph434Qc3FXt/EG48vBUNvLaHxxTEx/
3AVYB6CuLORx8QmkuWJSM5mKFogL/Oo5C+Q2harrA4BTFzuAeG3CCNz6qoQlUcTnwjRhuGZr6zSg
izgXUWAhj7iE15g8eJXHaEMM/iDYdIZke2/qJ4Pp8It32D55fASsgtksZVNCupxRAm1Bt1KqRXBW
3MVCvBNE921mEu46HmroqtpcWHurtYaBeOBhQeq5CpRrHbj1NUiOzZ/8fJjyo8xr8buDPXM8T49f
F1gFS3RaStQIabt585GzUuzlmA0upc/ccQq9XIqE/qqbzaOB1GebQ4SIRSDyY2p0Mz4M0mHnzffD
4RghnQB+OJ7RLyDxjWYpOs1LapSsm0SukAUKR0kRNFoCokznTfV95iKBvoGtKmuLfbum/wY3ehEn
aFOIiz4nSJUQck4AiKxRjVh84cf143n0G9qzO9zAHUdViCf6O78ccZBuWWOg2+J/W9itiRdKs29i
tnbcE/NoSWxkh7/NFWtqKsc6Han/9OuuEpH77PLWeo/p8Ek6LyvcUl+qs69ONdKZE/gdC+jvfL2Q
kNJshmqfQyhObBEHDW2QKhTL6kD0mj9bMCVdMxX0tQNFajGfB/oOLCujph1UIZh+3CrNZ69F7bIM
GqKqmeECaQ10GewY+XEN/5EYJZ1y7NtLCt5UueIF9WD1lfrQ+Eiljz3tY0s3+vKDpL4Xzu+yLcDB
SWknyFlPhFpzYszAMyKjPHjdQJV+eDc+vXS50OxFibiwMAP/6GfxTEEmZnwhWNTak/OcOSV0wSea
/dil6Wl6rdKc3jPdOPnV86GGVUPQESyzvsmCcdmiGEd/RDqgAsUeo2D+U2Ro9E6TdqPXEy2RXpZr
ZSnysF19+yBW0GTYlH9CMUq0pdJwgHcdUMF0N975FrQfjTy0Z4Gadqtpsn5woq0IIq2WrpnjmPgx
VbV/Rl/mY9/J3wW69cjfoEmYQkepNtfd2ZRbnILtEb7T865B8O+ScgIMqKOLfDK0gHCDAtpS4wqv
BXpVLGe0wjUZjFiWZAZgEVZBYX1kFYYgWWbsOssDyLDMpQy7YY4RY0yLfAZ9CvENHkUKiaCGNsQk
uPiiFVLi7YJECLV8tPRBa6JQ7KJTB83meX5tyu3gsCzlyBuwOsESHS67SY+QpWtU37XWSrkd3IH7
TZYf8V/ijMI606AcIbBacGadAngFd+J6ehI7s1SUv425hHvG0eTk+HOvewwqviRLqQM8zF29MPlE
82WhveJQmsS8aJ67e9bdIs2MzakckM2rFpGwYXVS4LGFsY0e1mlAMmp3IhsgnYLe9Ruo0Y6nHaVg
ZNPlx6P0FEV8Xx66WkxPXW45pz+DEwkGALgHtYP3Q4YwarcBgNYg5DEIsUiUws+SpJJpfpX+s6pI
f0/zH5n5SRZLUn7VZgJjADxzNRaLvLa5eWYfoScnNDLuUQw0Y6Ks2YxYXZFYihTQ1FC8yI2NEne9
YXmOgTrLQyKLhdJmFrAlo8nQSilX67opoJLG1OhxgSVtPNqoffWoSwrWwbCJjyl4mwy6jopIyfFu
MPsq5YV0ES3oDUsQgSIlv0Evrwy9yEXowrGe6adkIysTz1jqXbDWmFfHEkmy+vh50aVYmSMNhApr
8xTNvCkRg4iuspWNuCU58ONN8GxdOMHEJlZXEazmLZeHrsT9YPTHot0Sn/KlMo8IJfZif/OMEz6Y
nJXJxvnyxSZ66nUj5HYpVSoHTiKOX2ViR/LvEazRoJLPeLdeLvFuMJm2fYgVuJjprKxzhv8M2kio
2sAX8Zl9T8ni9jaHbvoV1zEIt0O5CPS8LCPm6PH6KrXlWXzSVBeJnncb54FnBPsDajWuIBDM7NHn
4u9ZRysM7vqYn0Ii8JW8qqYyZsBHXtS7M41g2/DIf4qDIXyjuSr62nHDlv+djys8ulVS0pWsWAsg
zSJ0ZGtpjCECRJD9txNOOLYMvlT932HmFYhqCpTP63ck+OLyEtWOE+rmmiL1q4zYoDoKuR2l+Oou
CpICxj4wR8vKg/VEDe+upgQXk8skQzDpP5goRlQHVhT5D/CQr/ZjibKv8rKvSpbmq4nAUcbaLhJl
JyybIxfSlacQROioDY1zGdih2bY3VjC0I/Vc6uEzqSUIjizT17ssPv7tLag8FwCMI/1jZP2/hoTi
9SfmRtu65O3PNCdsJThi/B73ubSrICzGdY48zNUWUgn2zAnA2vEpTqNwG661mU5VOljq1twx77k/
JyedHOSC09nWbsyzlVgWA9V8bvpsRpGpR/saLkrjtQtrzILqORku80CfIbtjRPf4Ay2vG7P+kNXZ
OanZIcQx61gwkwcenfMuWU8MW78eMCFMspt16LAJqqwP/Em1JJ+j7BB+by6DWQRxwi8pwuWDgyaX
4rny2FXiTNeZFEnUgHgMCLLyGfVas+lVjCdSzCUcnCZsElDO3z83XSE7yqI/KQ5Lsba5/gbm+JKi
sUNLLX6M6lPZzyAhONYWEMqxQt8DkAvw1deZE0kTxJ739MUSfBmkr1rFPEC5spzBkf4fzWDjpq9g
3dQJZ6GDf8+T8i/gSjOytZ0tXno8FY7fvrurrD8rHcnx2nCkNzIgz8MWXFYM0LDxPAva8IICGuAR
eczpBSNtKSh+KKluj73Ldj+eN1JfBqwTZeF/PivH1ScmbXyi6QYYuOJnCSDliVk7DW97ti1pAhZC
Z67dlsg+OhkqWkqXVRoi6Eg6HnuT4faRSB+Ejnv0hRqSBAmhL0BU+p19oYS5IeInhROdiDVaqfxf
6O6KOcOAvmbryzUxYK8aE0vuaKc/grMfjjADGIEm9M4Z//7a2O+16FLgikzA3LXI/mugzSQzy1oi
JgfHfXErBHLwo67y92wE/fU/i7wpJqTsLLJMxCZjMMsrGKySH05/G/EKzQuywP05mllA8U7e4tpY
VISBz/2HQhirYDTqc+Mldx4Qr39MGI9PZfDtDxr2mQVXwha9x2NgyahFMalqNY7nlIi7dIVJbQh9
CLVucm1Y52ThUmHdP46QPyIeRJVc0YKgT9K17vsJKv0JmmE9emGFgA8nmC+C8iXXuw0Bc1vnNlkU
wMI0xYeQB5cljJphew7SYpnioD/ZxVzx3DvAcnq9LkclizNMaRLZKknpY48pI/JZBFIzgOQezI/u
ziftjC6cZ2HE5nqHyoQ9/Fdi9HML75YDKpvW+zBjMUahRpIO575CqxlW5aaPmLsEKACIkC5IV9Ah
QPaZfQLj7h68oSSKVwp9Wh4fbZR33xNFU0F+Det8PfKlrc6UAm7XTOzeVH/ncGwoqnjfQUE1I0UT
UuQGh03Esl9VNpQBDSNMYWnhgQYq7mJOpp9khwuiB5Jlqre0ObBg68pZKkukxogl2uSBa6yzfF7f
EawFiUrsuu5nsSIY5B/H8m2ojZ/2GduH4e3yOdW6QHT6h2uwdNDrOTntMPpLE9qBpWHHHgg4yplu
2xNxdGRLmnQQ9Lmm4MTWfri83SLxf/ZuJOZSW08r5xcAZTg89/DkfBnqYrGMbRl1JLswuiR5o+VQ
WHkYGFBEBnElxJwpEXIP7x6HTLS5d5KEulCgjuwKKk/4ugOUerY28fvUXAx892zVbGepxvKmIsNc
K4wKia11YB+cdQ8mMOC3doysZm9ncJUmwS3aPJNU9RiwXCbb5T48L3jOcKXg0R0bcX1Jcsr/dJZr
oyx78T0dSseMMSbqbN9mMMHWqLX3QSSK/3u4qFnNeNaZcbGdSSZftCCYFq3/r2P2AQMkMzD6tapX
LzTLd6mhjsxrtD4QjoMd/lH2pWvtBGKv9pyRo4mNupQhvdN1lJ5On3xfAdVhi5WchTFCj6Qdgn64
cKqJmTXuJ5QH8yS7sqLpHZsn55oxAP06exQKoGG8pC3O2O4csiymbBw1/V+jtx8mvv+GMnYlD95a
fqipLIdPGED4cQMLbp/QyHsvgiRDC+rkOKha2Dqkr63rTs4FtYdYSJbQhXtelDf0/1WtFQV6FVhk
UOZsa+qHk8OTa/ikls4pPK7m0CRfWg92bMtiwxmUn/gox3JLJUvyZaX21ZEL0TxO0B0/3TwIIuFB
BFmCQyclJCZTyjkH3B6y7X8FgUh3LoJepRF1x5J4P4rufYBe+r9uM/eC3Tu1x2K1u7Wxmd8ub4j1
osxzvU6cncnFWoDN9WMfek/LyqM7DpkrWIwkQ5mhMD4iviaf5LSywnUaSdrLgk0fz2WxKzIHwKy2
f0bP60IgaLSy3Jy7njz6yKECYuw3r/6u+gRy8sNait/zDYvFilIzPo1DRPWbU9XAS16D1aoO3gwj
XtlZ+uUyUk+zHDOcS9+oqpbYxVb9/xvn4FZ40HMqHsVxodlNBVoof6e1xtqLijq19h9+xy50IDmb
VCKLP6VruY3/BoLTqjxPBBwAXZnaM8qGtkZn8v8dlczhDCTL8aF8PSc5lu0GBWhkiGZEg+Q/WwM3
lJO2L/4yFHoMLnuPVD30Va9J5liRZDrrrYcR/l4qAUsvBn3phv7vuwqF1SYIgES/vXpv3usuQ8nf
rzBqMt8FcgnJq9GBOkFcnVDUcsum8/VZOlbtmoNV2LMUacvw3d4kkA+KJGYurk4OZg/AC8Krb+tZ
idZhitssi5Sw0cQYfaWCnHUong34sJBQKn6G+Z4+DfEzBKvtUooen6mzPFeLgR43KUWUmNFdHB7x
UzPvoSZUanTZbxxTS7obzXsvmzJVNhxVr2Wy7J9+pDwzsPX6CMqYL81WL0f9uDrVNZfFdo/NZ/De
I+G8PLEX1AzJLy71Ry6Ox2X4zae0w/C6UqI1d2BcOtJn9wR28jXJBxPJNgoDi0zGu7IGnPgEa/Xa
27KN/jbQPKxSqeWXzlwwmVCBfG3QNzX7HBMZ2SdGXm2Sbo31YQH00in4d7D92BtO+7EOqk4Nu14v
F2nk41wEDUPUyg3ny6724V+CAQv8Oo3bH1Pl9bnFXWngr3pYHPR39aJHG8BlX9TzfjTa0tw/9oEY
ML3SheZ1xqGM/Z5EDGLV8tFn97Wv33kJ6Ddo59MinvxO85Oq3nwVkxGQBNBizrz9soJqAQKE+93l
9xNUHmgVQMOPzNZTISylB++1nRYD074KfRGsvGhXmOoNxsMlG6pMCWrsNFWWAj5F/K6KHMgxx0/q
z8dS6a09KPj3Fcxktk/KONArmJJzKDQKlcNhqKXngYjqX1ZkOErnun5urDd8wJN5KLw/ubNWy5vS
uQSwAx3Q2kaCOYMj1soZN1zaIdWb82Q4jQgM1q8+9Wq2tvQfaeAppDFV9hN6zKoIXyUxBwxDcHi/
hMAIwjos1OvoXh+EFt6Hn4F1bo7X9jpLKWRdDJptVHww8blQethm/E/1TUU0hECUMl/JZx/I5fd8
LOqhAQOHL5HZtbba25Gro7fgaEZgxVTET/5pzv9OejByziQaKIihQWtZRV7nDwn9ThoeIQ0mthI1
W0xZTEkvHPXcoSowTRV/TeHhN6SpAReWejQ52ENqS99mD6AGGUZvXRtTw7lMwK9DjGrXEhxO5mj0
gl69R/MDW/snb4VfD6ItOg1EbZfYM1xDQ2aj70sbniha/d+25pD6lDqquEoRXASxH2TRfRre3KDf
No+HeDs58tKTjhMXoKDRf2zk5cgv3iuqvnuBAe4lM3sgghoQTuXY5KjWuYdHEV011wQiSCxEdXyN
JfYgQKkAdoBGQnCnNSF1y12t7tEYOFifyLjk7C5Qv7f5/F7U4nShx3l1PPRgtRUWIeIwmla79laT
Xb22cKze0CKTtjPYXf4Cyw1+w8SWFbR65PR8wULiqhg8TSoxfxIuw4nNHOLeJN2fQQjuSbYwCJB4
bU3owPMYd94w1/tkfvuILnb9XtPpsbj6FRKVGaYjJb0zW3IHJRYSMUj/t8xUIzDVWxk3DEPWoI5o
RGq04Vsd3SUrIxdn+iNBq5vo1tMMP79kpXsyeEpgI3Sc9wk+pIt6QT7ffMYNpMshLeeU/GQUAYsF
iuNRypjMk/gV3TVxKJOq4iytwzbNwKVdbKpYxiWlXnUm2jV3kR8b9k5vZn1zdSwkLsUBdsrHFr2C
DOWW2Nh237CaJg453X2Qr/TAU1XX21nDbPlUspeuj1K01xC3v3//mLqML/AIBi+L2UeSMnij2Thi
L1Ilk11MVVE7vdrgTP913rCjODTW+h8HU7hj2p0mlK7VAYCs+7/olb6Q4dVn2CSm95Cw7zrVQiQr
eZANRM1DF+WVt8ZvrcO2TwrREpTMJDoAk0Y1f5QEfxBsSG4ZWlUFPrdJ7N9Vy0ueQZN/249TchEg
RxaK/kY8ou9ELeUkS3dCl5MgcUuwxycHaO9ukAQTRa0ywd9002N7nO2oX6Nqyv+hL7HcsyGPYXqy
p2FtlRNqFszqJPoeZQID4+4iGAWpKI6Y+yjqk7A/4xIp5xGsLWrmP6SzYL9SE5rUqXhBAutQJiQu
Qve7KTo8GDfLJD4gWUnefMnHM+O8jIYBgfht+eAl63RFE9a6tHqVAUH4xjrW0/8TtnuWtMCduiAY
6cMrcXmdGlayTBKfBFK1hcQthAVPQ4nWI3SGfcKM+YePp511plTu4DcjfA+n9Vkp1dAARSiVw9X/
WS4VsAwcmho2+VLRigCsQoRvcwzgLPcCAjbLwOtvnHkaUzS4fsWCpTyFc20pFbtUlIrFXLMlCk/6
bIkEj9QMAvJpe5GCODpi6TMUNqJkEk/D0H//+X5M/JVSfaVtwbrR8YDwYvllSQ6Btm7sFKxWCfJi
2wJCSIqVGzgHSMGVKF3/BwekI76HnwNpQcl/rj9rz4dDIg10XRAwyudfhIhAboFUtC2n/0lyJs5G
7aL/t8RWrN+3raIbwFPUl8y+WG8RrHXBHBroUuyH7iObQJzJEovHunMWEO3FfX0n4dxeb2amzinO
2gImaPE6ycsRNKMrd7Y04Nx1P+NrSM0JCJSQ392dSa4QTyFQgcsdwkqMVfa9tyIp6aop3FAb9jlK
EdtB1dVgKgCE5sdQXAUS2ePRBH4d2DLe+gIpwYqKYiDOEIFkxrWXg8VnbpgqJENi7R4MksPRQSLh
BeszPfqlNSUf3sfZzkro9WifWuADlVXre8neBYTpAuIrMOhd43CXvseFGL4pYcA+BvnTcK2z+7K6
PLe7iTUTtNcgt9NmCIDAsx9CvdewR0hr78W1LFy6zsdDRXhqDvwbqALRSq4AFgVBiIgIZmAk8q85
fU2mn7voPdM2fOZMiFJ9wsoMYWEkS5/+M31RpPaFNKg4vs1+sqyYa8acw5Ldt7FWO1cb12G8Ne8x
a4Iy5ay3w+qH12ORx9mSifkafD90/ORtcX0dJ3pGO3AwXeikvATrPzoMO3Iflj2oG/tid7rMyRpU
QUdu7kTnC8enky5Ow/DJTmAjU/H+rtKs1/MeDztZf7yRvRwd9BVy4MBqec+GEF4A9qBG4sQUcfJ5
xxB2qUir8IPh4uwa8yYTh1q6vQlNNoG+PcoQqwCHTkwR+KhkBfpf/9wprOHpb+eE+/502EJI5IkW
33qCKLC4737QRJnL7HITtEw5aJBUHk/Ly9CAZPRcANsNyb+irxzxQHBkv4jVR+ftjmEaYygdLwZa
EEKjfaPKxjrRZf88Ox/4Lxe5BXAq7nGlP6lSYEfcv0U7IEmIon3k4tBhzNzQc3MGAlp5q+N7rdax
dDWeWSP3xZ9WQPIfKZf/+QjPdmRUbXRx8aiYXrclMw3RzBwQwj9mWLkoJoF/nk7/gTosCD0jODDZ
YR2hKP5bN9E/xja46Ea26GfR1cdxpzsW9uQiucifufq/GqoTqVxIzhdD4cg/zG2sgl3jlWZP8A58
pWdJBG73QXj3AuJ7h10iAtBipkITJRJ/zawRdmbqWQ1xF/Wbtl9TTwX1ulo229RoL8pz7NJzKlc2
gQHEd17N/ncMUI9PhxtcnAeEqCJmERfOKXrqhbSlkXiZ76+Jwsyt5GahI6zIgUJGl55fw/wsZe/w
K4cttQ9/0I2fFfVraXHEI9Fk22O6Upwubvajoch985+q1p2sIloTsoo5HeUdp36BGoNqXc7ghBoU
8rjqZKznRp3iCyvkxkXntNIersmh0WTMGfEL4gTmaps18L1qWsWTjGaoE/rKUjck8Lc45KMMY27W
nIGP2Vxs130BO9V0WInrpLgdpxq4Lyt+8tpXwYkMffV/TYxmXIx2snVVP79rwgNh5/zMFB58Uxj0
8iOJkNSTQTsv43E4Y3ix6BHYKiZ/wk2wJ7ZtSPlTRcKcPwCUCPMa06R3VipVeH04ceVnB+bOnhAK
X5P1RmF8WbY/cN4vwdhu6s20AC8fGWlg2uHfpQT46tlUglqOYtyQAxALhSO/M4zyjyX6FUO4uALU
De9LLGEVsKtckzrldgknSiFB2WvMQjkWHJUNgrs/xtjoO16G5cnquYWEogEGpZ61AlvdUqifaOGc
1dX+b5OxPVsYGq9YIY9fldb44QKcX90ykkuLgWV/LbjJXv0WipQ+FNSFpl3NCWbcmnrlAzeh2YVR
8wPlMyD7//8sb10M83hQO+9HijrLXCVzcHod0Hxn6Z7VJWmKX2kqKQUSyaIqAMDEKVjPFAGE5rJH
jCMWN+R4u0pXg/grV/rvU9nf3T5sHG+fbxv1jZhmSGmbe0NO0YIkcH2V+7O5zpNVHshGRIMeW8BG
fPJcCOYWjMKFmPbx/0uKqJ7s9qGA9DerRj8hr0ZfA7OFY5Wb7ysORoRRmtjNQPoRwx3IJgIqWX11
GxSORV0jm8XYprIazom7JDDjiBcgGmgygi7lEtMszqIcRzSKz9N6mCOkyghZlPR/RO3hMvPVERzB
7puS1FXRnD/eFrO+d3NjmWkdEDdWne2CeIPMP3lDd1oFWoOWUxLq7EKc+fC4QxhS5A6n0+MLOnYY
pmRwEkDYlWYeSqwDj/u3tE7JZgUWHAKC02Fp6qU81DzdcnEyMOWKJGlbTMUH1ynEUxQknmHVHq11
Uwd8AvEiB8I54zFmNcXjZXsSRK1UVh+qYYJ1ABQvvVUURJ81Ja03FqRoOK2cjW/s2LOW9kSuHvqo
VgnTUXAuZzPZnJxpetnW+baLEApx1wwKDob7iL9/8OYuFsx4K9rPYB8QnNZsxVTMK1dz1sLc2NDd
oY328k3WjYd1XJJLNI/+PSxudzZ/p1nxCfaim1gJBKTnmNOI10oFAPdtEIDowti1UQn75im2Zwmi
WwtBW1uYLjFQcGj2m0ye+z9g4Z57WtcJpvNwsde6Jkw8GBqpbvPYEnliqe5xAJ1eakY2cvPmiLvv
GK1MMioiIfp9CXVPdHtKl/8lWm9tv/GXIuGB0ZIV7BEcQhZvSxwSGuO+2SsVyMZL6/0r5bscOHFx
weSS1nRceaU2kChelhcpsib0Cqsf0tsegufAog+xfihftsd/X/M6i7M10vYiLBhvBupatqo++PN2
NwGPE35WoflGW0bu8bhCDiDZ0LMWHfjxmMdDn4BBXLb/KIi22lw3TjbLTvFwrxtHTELfmpAkkWyp
Igpla1KpVzEAeiDIc/oAK0n0zFxzl99pwl/y/xziR3pe48MUf7v3LFNOXSkBRC9RGvvYQo5Lzx8k
m8sL1rbHnGUSBt7sAJ6KT96B9KW9ikv0Fsj7sZOXTMQ8FpFYrbMgBfU2jTewb/iVIImq4A86KCzp
8Ex+o5aIlT6s70ugtgGLD5ekSa5hacvN4dC7JRwRFT0/6fsxzzWwAF9V+PLxcFQr346icQmXH0Ku
nx/vzYUoxyc6mSL7rpUVWqGTAZYdCHKPBD9WVRBD4pnpaVUjaFr7JxYswUZobSbizQXsGC8abfzY
76t0kRPlacx2vQ5taieHkteARmaIAgbR6b4cDw9NpAcmJa3MK6L5rVEpi9Y0SfG02xhg8Z+1hxss
n8kriVEEVYZgPpzGOmIZ7kfdZT/qA9llI8V94S0/ecn449q6B0dpuQmHBrL6h0KQT7U6nyM2Zsyu
E69Ci8hZRSnFAKMxgTCa0o4mP/l5L2qrWHR5GGvXULEJoLVaQK4YVqyujnfjyC43SaJryfGu8fVn
CtXsGtJHpWrYZPryHvYL2MaOAMgnvszp2hS0JsjMbEJPuZ6HgZN2g92xX/4nqYNdfJKO7Re5O+yh
pjnWBPAjGcEj6aItgYVKGMt8LEBuLj73r6IHswFq4+ssaTDgmsNv3wSr6TraB3NBtDPY7OuHVZUS
KPSNtcd9d3nhs4u873BZpJ95+JjML5/sgStx+5hdWtiScULlI7PqV0XXwJgiR33rkMeT1HXQAXgw
QjV16mLkJMyVJwmCFMPoNMpmE3mzZKQjDVh4kkLc2Wa51h2WkO7YRUMut+v5pvo8sISnE366FhZn
Hsu6pdT8NNg7w8aAL+PWSfWr11uzW35P5Qzs0fXBTKF+OZha0Dwr+k8p5v0JSQUvApE9k+DSRvcf
oyqvCfsprpU6hxxn8iBZ5mXTmnblxhUrlhFQCGHpgPbgFiL019w8G4Pi8mpuToXeeaRFZNJWs6Nc
Hu2k3IvCC2oPvXqOUCG+yjtvZdZ+444PfCTaQg+ZvWSNLwcL675CtFZBAukowqir5M9Rqduf22X2
oml7adfIJofv4QZq6oKSmvhq10zNmDbzVwo7502GdYQ3Qc/+7hzR6b60QnEKG43WtHGqzIt7nJwM
nWfFb/Ppy6h5b4arWRNn+sfgCGoUXLGegA4GLN/4/1rhByaBMGi7fpg1752X5fGa4xRAKaHdS9MY
vVjgBkPv3f/sq4IiQhn+DcAGlE8QXjbNcrs9NjlbDWccrQr4pfzTCBmkufO67KCl24xFC0LB0ya6
WkC6UK98YZ1N/+B+uMTgmZSPBYzWS9lhHYENxz2FkC2BPBv8X+0O3Hfdz6gbRSriGh9RLHwXDUni
017LRzUyMdNF8MPaaoM6sB/W92lt5In9WnkF5mmdaZNeS0hmtTrlE6yVF9kWIB2DECT3bPd/nBKc
l0MvrSY7CIvTTutv3a4xI0LFGk5JVyCjU1g/iHZqUOYKpubeqXTHtBNo5bT5fIZsX0eQRyFoJQoM
Q3B5fCX+l3ra+uafFPi46MrPs+oLI7R8lLP8Y/eb3K4rOubuA9uCHf4JZ88OdxFnmLPAc4bn8gq2
yHT2+dxIfEe8OSie9NfoQUyweFa7s1nJH7vtvivun41QSquGPgfOYWZ9BYolsKyaHSqAtJ6I4Ohd
q3ggzQ4WULBjjKDC+1j2Wk7gBTiNyaH8Kw3XCdGdDMn//DnyvsW9bMip/4T7yAJ/sX3FGuv4gyaD
M5EOFZW8vA9r+Bqpjll5G8BdcRYAhMlhX5EWiGY0Ht8FlSgV1nblxXko7AM/UqVOwy/mt09ZZIMH
bXrm1nsAaKbH5GDU11EV/Aezw2pHOA+awDo8/mixIqDFTcPwwFMpsPJwim4MUdIHs8/+5ya0EylK
KLy89pc22Hx2cChp/om7jcEViMnwm3geMpEXqnNEcu3zKIYkjn4CU6Zmjoq2HGQw8ix6rdL5Td1j
ffEQD0Qg4+y83PLYlKBj1vYANTfwTy9+vloOphq1H+0ou/kpXIRbfb77SBahnj/XvCvBs6p/VFwH
pM6AsDUK5CrNsxhSTNmARkayK76rSWJrp6Bnd2/kLvDUKe7iAKPl7Q3bVSKN53BLejXh6VTwfJ/i
WC8iuOrvwFadtpxZ5qigFz4b1j3A8HGT+7py03rYM1uLy1u3n6QHK2JAM4FiwfqstKOZiWmRbKXD
qjRiEEGUz/K3UDdUJjqmHGnfHiovjb/vQa7z1hqSyCN7p1WT8hOpW9D2U0Oar45/6qPfdhvxtbCD
QHU0LZZqAHHLl5hbKoJSjOgvDh6CJ9ubr1B2DPgT6nCu+BMY8eC2nfTBEzJrcp0Q1yKvEY0K+eIX
7cYL6XD0VV0HElQ1xGpkdaSfS9cg4PFC+31lZgGXL2bzm8cXRLRqqx8uRPEA6CsQrJQyD7RoqSc3
fQZPx0PssrWtAJTD//mc6TGIQolDx/cr/YsodEaPK22awnum/jKyRrnsv835JMLt/6WtBe1XvvgG
Kc7ZVrb7hiLNaSqVANoJsN3xvPo9wktr6Zq9aFefwMVjkKnb2YKSR92J/K8zzXiTUrIcVlMz3MWL
TAjPJZTGX6afT3nZPcjp7CqvS6NCbdKBuGYzkQL5S1LRmHZQEVGks2J3CG26qyKHedy/evIJWKPW
na8zAKlX7FVHN3j6F1MS/otYPrnsw76qhUMc5z5KbbxA5rdnBtXDFke4tgOgoba8ADJsERp5uddE
swhTNdhM9bsSucLI/x46aMOoI2HcQBw3T5jRsgjocwIQYSY5DKVP+CANm8z6dw6IMmEr145PswZd
W4QtMcdbdNU0aeXyOMccVDb7KpDA7IWbNEBu6udZLUVbSiOrVa+hz9iV4phKwqjZdThXX6Azj7+g
RM0yXRcetB3dJDteotUr1D4LgJJjxberp9KSHXKmPZbuO+VssLtR6Zpi2zcYBZELhgG0uVlFoymo
+j4HUsg4RoLVCUeySy+ZQ6g93i1G7iFPFHOEr49cJDE9QySs6GqhLMlngJG+pvU4cVaU48vWcX4n
Kaxkg0GJ5dh/RBjXfZe059LtX2mgBu/frN8MCV5zYO+ABaXLU+apn7IW8sXkPGhypBusunPk+SMN
xt5uAXj7c6hVP3wwUOu152Eg7ftiuHt8mgCQY6BKILFrj+7NJMu1Zhdxwt3uKN7Ci/zZMSPzf5wb
4rBlnNkZ7FLrYEOSI/i8CSjxMoCjdZCxw5n4zRhu/WLRA3P6LER6ej51XzNmMR9zZtW96Bq36U6Q
CMVwW1UA+a9LyZ70pHIDO/pKM2sbuJl9U9aCV4kGVkE2XpYO5Ngfc87U6z07Y698XsN8nt/0Q0NL
51gW+AxpDkKVRopdxSkfU9rFahAeiYpfEs8J3cegZV1QGQaQWuLFltB6ITCCQbsPdnL6AczGZ4Vt
lJbucpNCV/5z3hBDtFf4VBBJMEhlHAgYRPRkSVkZkwKqnePoSNeXuFSrqj8eF8RwN6TPaSvOT+zo
TFtfLcBlE8HaGF8mPXxyghpKsfraEEQ/lJFx2NYMcXjHNzY2WrEuOct+VmCGMimO4fs0mhtsOYNJ
HIYb+8QEvLNHgQsMXXTbhAZiYe5FYSnFlZiw/wzbCre9UuD4yQ4XjTCo5A6ZSDeu9UrC4b3AodUK
uFcJowjGeYoYkgwe9OYcutV3W1rie36gCXJOGrIDUm7r4YStp1frMCDDsWq//9otrrhleZ9a1iej
u9pvzMbdmQvV0p0Buv9QQChXQ0KaHgXWlm9t+x6z4qYgxo9PhpkJNahqBchyoSRnCc/exGJSZFGn
I/gYeIy5A4/N+Q7bs+YtxSTVKhYEAu1jRlsVbIV9oLqR4jSU7ygwNsx68nsOkP7LMwPug2gV/Asw
K62eC1+0u0hw0TH8Bl1VEK34sBmvTcfo0oSVNw9uhHA8jVnQOg1zoTBoNT5qoGEcdJnsvJFm7hM8
9S0AaZx6C1BQPiPs1MsYhcmDVQX2MEs2/m3pUkYmTJwYTLAOH0fxkK/MxykvYD+9m4PSIDpHW+YO
G4lmoJBNXR/BE194OevOvsTl8sKebSnIrKuxv3QrTt6C2SARQfUfKDOx59cZ+UiYMUyRjouhYm/S
zmidMRk6UScBT3ePBEktbsOqbPfW6XzZ+5hHzbYGdaZgwSYNDu97n6J/DMP++9xfI4fhT/bXqlBK
HHlmYutXoXjMGRtN9Frte8z+xk1hayEmiHKtgVZktG3WB0Dr3KUUhpix11YTQNIR56CrABthY79b
pqmCs5blw9bmRY2C+TXl96oHoqgQ5iAs/xWf4x426o3mn6Dna24wB+GAcBjkTW4PMQVAotx90eaE
OJSQjDoeTPC9jur+jBzQi/zbm87okIhWJ+QmWtOFQv+VrNAhwnL1Hggd0ChqTPmtgkbdXCkuU+kl
0NbPAbAe1MiEAWkSzynSrkQg5pfQWn5yrBG119rN4Ge2Q4ca+UkGGI6kkD1XVNoY6zhuocFN6CIK
rICdezF22uW6GZwe3eyKR4ekiWF4S2kmSJ6mpzN8SUMkIHcQ+eYJkamX2Z6SHa9dAZHUZ1OxnLj9
FrptDZdM6pXX+EhIq0hKuVYMFccNZBPmoaswJViIzKwPZ6S4Ceph9BySzYQCmAXpKdFPXlLWk1j3
CxIJjLNuAl4US8y5ecb9QncKQ+nriZT2P1vepC69azkSZqZPI6krXs+cjbSc0Ea1fhVWYamlfZQl
2PtqM0l3iWVoDQEN0MkWLUjtMV+oFp2Yv0zmu+6xBXGUFwz4WVJwjUMAskp1mA2mNBAn5vHEN72R
fNs+CyDGxUO+C/Wp1lOvR6cSCw+0LOfn6DO4NXtO35dRmFin67TEn5DRd3cXzW5GgzsmSq8jrkiO
Rovsx61+G0RWeb0HaaT5lWmRi3iRLIF22lIAmAJVkH23+f7qeBZhsVk5aCM12A3vl8fAY3b12TAj
oDI/VKspjNOWuKhn+LwQRhw5X8Jp3xIOZJYcLGZMhivSPygz9bXqGzDnXpipDIPt54OeoQrVKBxg
SzTjrWq0zp9kgs5v19EhdXMJHjvm0AvRcuM5u6apJvXr3hzUEnX3hGw2Hi5zsTur3mxCxi09DwKN
dVENtmDFuwjy97zeHrDNxEomArhskVOCNj2MuC/GyISIV17OJyda5mvbCmtJWuRV+OcX07YfwKtt
NpekbDVbTE9m3aKxip54gw2E//0+RWBroesylqzN6Z+rcbqYsJe3B+NJqfEVKihzcDEpxZPfGzWE
jbJCi0ivxvpv0fBcL4JhRu6DFxQO3o2sQgIFYDciz5xJKxr+izE6Jxb68gq0LW8WFuQm4ezuNrU/
78TwVAWGMTsUyziquYvPbj5vaPxOCbblEvfibOKy6abMdRj8HFrW5ZdY2zXe9oPHyPOIAY2DbPXn
f/sXa7RPn9bL2WwrMo8bdzS9kq4SZ9qMpOZkwyeTpyWPDf9KXaco+ucBm8fwhCD/stuc8kH/ZVB4
6eIsQ0XLdyj1RUPBAkmjsv+eSyt8zIMS4ML6/8Njh8J2KX2fvXbgZCX9nFF+ZfZIKi2mriNG3ZYW
cE9QqdYy7NhH236HCEkaXE8mGJgfw2JcUDbsdgXen3ylpgTpEITtzXkhB/eA7jXUKifDkjs7YxWF
+k2ozKV340ikhRVQy+SglNBXOr4RbBxH9L2WX8HgsuyYJIkEZW0c/+IsW5zciAuWMAuqU3lIByvw
MyR1Ke/69vp02GWQ/Rw5Vrea8oNaJOJ4fkeDXPQbp8FsdHaANk3ZhDo5Hsw4RXr3AVlNZLNQvRT+
8XI3SUKBDZ6jJPoRe1weiYi/RGeiv9r3W1+BhySgD4uCuuxm7+CgP8ODkeLPzDZr7OPLmzcKmywH
2iTWOcYvAtNx1XoSiUoRlFSBX/gT5euLCLEmAiSEHiehsfxXuYeULmYl+1zYoMQFm5dtQGEwIXDt
SDE0/L26GvdD4Og6OCauS0r+08CHIBklzcwgM4IoMIb0VrwYh78HrpgQ8LQDPFVx9h6Azkd9J3YG
K8eBkV2/dPAKMtkhFaPOTi8nrh71mQru171OEBwkT3Dtn6Pm9pNx5w0zPUYtrKn9UMln6/o/1/qT
8c0PZmvokGMoRuVgdha818bgO06USY5cSg3G8NKZlVII0K6M73fwX3FxLICK9DKcIYz/PIlZCmOW
kwCLbQb/v3/iP3nhs69OMoZDot5RJ0cjIahoVi3EmThTPuhB3+ysr+kQLYsH9j1dwDuRQvQOVcYx
/EgfmqlJbsUkRJ+E/0HOtFktqGEdMk2wIwFXnzWmVLNEA7nOF/vFSiNW4tn053B8cF22WpgsibR3
Ct0D1IFkor25TA2esmiQ8X7WQmert7S4aLY/CDHfN5ij7Cvb3lJdk7D1ApYsYO9JyIrs2IIoOK7O
Wpg87rNc7iH9smyVuMP30NZWckMVh82C7GCS5JqAzYYUyPfXWF97JOVkSKD+AzNGleDmTmCf5SoD
AheD6xHqV9PfhyoERrwN8lZn5p6/dO/zrCfmy/8Ppk2oxhqD4SjvYXmn4Hk4PdIcw2WTGDghS1pK
W840MhnFVx0vuzwpVdlt9DlaDwoIA1Az9qdqKCInQ5ccIxkfaStd4fieVFxufVX5S4aScieutzs3
hrseCfdIOHACyVrakbLUeMSmyncHPI4o9YbAWrCw4VDqNtlFxuHlvdaSOtpqnsZ4BsBLNIIeDeam
XNcY8b+CZf4LhGdr2Dw9DbsMHlWIQ7jPZ01lKIWeKNI6zDAp8DQ+41lVWJWDzsJMamv+Qood3ew4
FjTh8AvTBBLpMhAEYG8owpuL31nuR9f1mLLSlssuHQsb6M9nqP1fpvlmxfnR5jlzyB8L9tPcgw2D
+XvRWPabt2RoyqlXMNJW5vu+zJkmQ6BriDt/lDN4XbHQyo5NIklmGcUUwAj/0jB+5sMKJbUO6ZjG
6OhQyrFl5OIJk/QG38e1h2Y3q/0ktSLq9zz0p9OgxU9ZHBI0grsJJVu9F6JimZOu2EqLv0mjK08A
JmcwGNptnhbMu/Rc19DAOk4vbwuuBSDl0FlD5TImqXdk83vGMjVcQxKQ2mwtyl1xn0wcGxP7bTSK
ansYJAcIetJ9PerKyODVRxX58uz9d/vZF3He4maOd/kQHaaJXk3pd/FS/pFKeBf9NZUkigdlOsUB
f+5HLKwv5uZVnDA1vPsOIgPzQ16iCOAVauSp4kUvkLC1M/E96Ub+pzArMrHQr941JXcMjw8Waj1R
Ue8Y2Lk4Lzvcq7skSj9N5W9R+35X9USnwiYjeTU+XIlPdS1bFRL3qT77jG5p42i2kr1s+US6CDZs
SfQOWym/eKdfEMDXM/gzTf6rqELYgqkdZpwBJo6bEA/WzpG7wLXU7lMOZjb1aniKrT21G7Hre+j9
meLF61iEgnq0zdSxqwC/YdFcUAUUfTKXYCbIamhbEZrzeteP7NRCshUqHDwYINtqpN7RQugJKgZX
kXygYCVxC3NLZDafS7ZS9uB48xpUQg+l/533Un1om9tiqMBZ4/24t/tIhDGAu8E4Js/+iq4bTv/q
ihpnm48TME2G8Tb0yNGCJmOucMVsaR60GLmPYov76W2JrK24C/hECcrqmYvHeUCHQq3vQNO3I3gP
fzYd/nZs+Y3rxf9t1/y7EiDppiqqX2yofaf33dlgWf4f1dmnnt3aSDAkNKCuLY7oSh6lB9epQt7G
RghGZPMzeu/lPIpxA0eUev9CbM6ufBR+poilj86vAAp/m3DzSh4GSJep/lPDWifpI5FoTuse9wXJ
UWFPB6VIeu5TARWkJdbmAOyb01Vw+rTGpsIEB650AFr6Hs9uDah5W2bBNKkbvnreuet0+aJ3aU/d
ju88AEdnLzJn7zB1TTwuStNUoHm/NmoH2dSlh7g0Fs5yPOFPJbO83QjRyApD9B3iq6AUMxYTVAor
WdC19xYl1Cvf0Do7C0VZ++OR9lj2KT7kXhs9dU+PiDRrhff8XkBLVHE8fejlCzzgEO2AkC5bmNii
233zf+ib8fa/SVDcYZenVIyHb4GZnd1wZbQoGWx22GzzdEft9b9mmw5Rxd1pF2Q69CAA5Esv5Jk5
ZC9OtBbKe4Re9tNrYqLYZUjM+b1XvRTqPAHG11KTEA0awNoKZnQWQtls5jPqK8vftlDp/h2vBfc/
qW+cvbirjh71IJ+K5msxKM4WFVl3L1QhXxIMCQ2el5HC03w/Ih+NfGTSRpxHm6a5Wtmfx81ClQta
Lu86hrfOnthM5UO4+pb5ZhLRpVdkBmjutOHGC7MLGy9JlwnUq48yJX33f0/YEU3bOhwytWjNDD/G
u1ZuATBrDQwn2bO3/HirnHChueBzKI2Yr4njxTqNkCgBX9gU9Z9OlnVPC+wUkQm7nzMFEg+3MlIQ
9Ksp9kwc+oMotoI87qrO8v4fDFU4GrIVIut7F3k4RGcuLMW4DmUZoxvEIfr4Q9XmrrACDxVaChSj
Yu4oixZkruJ1bRF0ReXICGv6DX0/vw4ecU1DIqaxC5W2ImUOhZqLosvpzh3bdYse9kebqwX6AK1f
z5Ax8EwYEi76uS4QWaqigE6GyY7BRCKxKTe1P4m7dWIkrFA4dvq8fa3lapJAVZkOCyUYpIEf0O4+
OnmXV7nHhQ3LEP9DOyEi/5FiI97eD0ZSfPkCtm71OM2yTmuZT/s2u3wbt0JYds0QvWN0aQY5s9qx
elLtscgVKs9oQwteffr/Of9TkLEf0f8XTMSt8g+DHKx9xb34L61jxUXLf0RlTBVtwSlA8M6bsHtH
1czijk3lo3vbv/FfPVBysyjSMQkxfye+6ekvRYqZ09sHjJnBa8ALC4Fpxm0wLuM5WVpCgH+7mgdx
3t3nx8+Tdehpd/CM6bPz5PwomDiabjzKaSXW/+EGQHhr7rVJyjSxSFsFpcIXwo1QnZvBdr415naA
zAsLnfLOb9pbYTeQ0WN9jI+oppTo9T8eHQs7HYBt7fNoCFk2YywJzbhuvd/9a9Y0FIQQuaknZAn3
9jgdFRttjbIezbVsrV/Rgof06zJALfM6wpFQctmwoA/0HSydOrpmt/gSpLTfCJuCtzyP0QdvCsjn
XrARCGYjlJ74WeTAwSSHZ43e16/ORB7swJSCwceYMmwhVBxMKFDYfS2qjnsqQaqSweQmAFWmhnJo
rGk38+bBq+FJMT1jRH5vdTZXAELsRrUji0fRdzGcg/ORLqPo33vwwMO9P+ed1J4SByJj5Qc9FEq3
RbxoZk7gKb4c+zJiWmQanHfcB5e3If4Ly7Y+jT1WXn9HIdsGAJ8IQchz+ld4WTH2v3aWMz5J4fVJ
jksuw5SA3OJOR7bq/NHGdCnKoYQFqluxKkXiPVWhNofoGurN6JKLXfz7FvwLJ6StMA8LM4NsqDWE
BJcVKZqxACprFP+wfXIANonWHrxTg5aI/H1ab/OAr0Mv0pmsNFj2NP1GDPIeUtqhiTgUC3IxFu0i
4M7nx1Kt87/Pe3aWnSYzEy9DV3wuKu+j91Cn8qAHncVU4lRCjZMR3uNWA0ZqNb7RCF2OGgi6PmcA
6Lazf6EnnRvjN9yUxejKRWHCFPUSHav6xxT4g73/L6coCyi5o9CBPbO99X3UHNtnHUp654GmOiJT
HLRL+P4EgR3HZAPb4nH+xdWxUQUlbW8ywVXTM/TvN9N4nFKZvaYCdNdoDCPpMTqvO0770x3nuuyJ
X2DUwQ7DARcgPSL1zKxiVZFnTfkb6nlr0lBtb5xAI0JYRXVYEQMbtepJF+9xa9ghGH889W/eP6U/
NlvpjN3S8TBYcnv+byRX9dggumXeY93bblawLy8g9zhw+8I2838v/bJiNJTa/+KN/lcLIg6/fb//
DNkIaK7ruWpTsmcfeyaubc7m5jb1kG2lsUuLh3bsdv460QK3FhLQ2DSnXnj1+t2zmB81VvTmYLIJ
bb6PLbz811KAuKvdXO044vRmj24Ai3QcdjZOZL6IpxcBF86Jp8qapAtk/Msh7NlgenTmVjFuc/ES
GvEmwlAMzggRVvnNaoqzJDzUW1m9frTyREOCKIpPOEdN364/sRUEWp9+y9DbpijWg/tOTzmR8QUD
ztU+kmiFkGECCntchyEQJEsuVcmfC9InTju+cA4gDULYmt/Ht6uQoNPgzr9pttO5YyMtAdftkp+k
gE8/JFr3b6uxukR39pCsqUgumisgrVdOxO/I2C4jX6/glPINg9RpPZkQvzrXTiWpidRzkhl8ZXkX
tMUi5qP6mERjwhJX11f4vn8u5U/V3Ie++dc1OeKcVAPUSsgpg5fb66rOchqUV26KnoEIo4adprtw
OTmiBCv/C4wNOnKOuMNuQK4Fw81LkR+/9AsPQHKleh7OKwhGK2sYQCCz21c3AdbBiJ6KgLSpjHJi
cPwT9Ck4PS06l/0Ju3XVabIjevngTmk+WnP/kap4HUp96h/PyFXisq3huOSH4nIG7JfhKraYIhqJ
2HhZ6wIY1vhdPZXq6RPEdPiNyKWQUNqJ82tViVuDzlcC2SUOyG/MLLQNf4kFmwnpO1oK7Oz1EiJ9
M7nX/5hpz3KdUpIWeo+uNPFansF4gvgPJsHK2hSYRH85/nbaeU/Jipbx/uEpzJHNzRml6xY+PeOh
egpR9Nopq45O1DX264qLOvV23Sch8LYh4Wox9BAITKMdyuJ+NHHdKoDnxUj14UqBhU14DJ/O5ceK
F6We47Vh8GTiQK2mYhF5H4pFXJdLCcUW5KerM18g3JC4nHyyQCk4HJ0mzEjfMyPibWsn9g6rGrV9
GBndFMc619ckqxK5pt8ukmMRQvhNr14vH2ZfRN6c3sqMt7t6F0Pf/1DkmzeK0LGDUndOiDIL86kh
iaqmJwAqlmWUCuhfpgc8MX9y3+J7xVv8WPQ8wCIz9Gx3qB99iM3fvt9s4tSQsCuKSAhm0r+w80P8
VHgwNqizeruuDq83O0RAftfBiR8U9w7K396loCchkUAxnfmjri/Cw3CRnNI+l7pocw5IF3oEhTK1
CazsYuwHFyaEf64JK4/CknZA5ioT4FA7rlyEckyGC0wXRTqbWT6ug0cfGBtO2g/Wp+INC7gj4VfE
y6k61wtYj9hXLKEzME1B8v1G+aOaBzx8zJN94B9yW+i/K14Zryq21eu3ExtwhAywASz7LDNcmhz0
ib/F0oF5UV3h3Ob85hxJ6OgA7P7iitfsDzrL9zmy2NUAurGVDNHtw81l+FH8zeaz24rzd1SkEDgm
dDHthoWgGUeNw0ieeTmvAG/hAu0Eh+nPNEQpt1mqBMeMctcRIUbhrnPBYWvuzt6LJC8GXhx1N9Fh
cJ0+g+jqLfjJSCkbWRMxLpSFJpZD1iQrECIBtTPXJTVFO/Epzh5v4c9/WXhcbd/O16JDYCH5ZuvM
OF8wnJoks/+e6LfstMqzcdOqq9kcz4ScPS9hVP1VYf/SnzCNFfCTx4UaT3X2Rn/GXazojP8iQ0Rb
qo+cwe45/LWSjK+a+dxXJFmVh+F/R8zshUzxMHaCELQ7Uw3gSV8A/Udge4YJYs1d5E1LngDKbi5o
QmODej+XNSyVxVA2Q3A5NXCE2AsqEIz1NWQCnm7Y6jko3Q8bUS4flvnBIhHUKbPTA0OLquYZUGVe
+pJs5ny1husoPwBUaZpORzGge2/oka6JOhf3Wp+DsiepcvMxjc5nKaPKZshsuB6yJXyf84VUNCIn
AEPCX7LWIx5NKO5qYNb1dthkMMntSmbz2/uDkBbvIsRYDTPVXmEjFZtOT0P0eV+x3wTskY7U76aO
H+5o+s66LMJtbwbBSh1xqw7Ias5iEzinCDfwJ4XrFtZ1n/iUBXvq3u1z9wBZuqDMPf0ckhLWKEG4
4FRJVw/287FGjvWqrGqXu1gMAS3Gm5mKpWNba2FhDVr97IUO8NzyIxjDOejsD7uefcVJ+e/WH7NJ
EB2IIQYiFNCvqLgTkQpkycpcul7prZrcRmkGO3FKkxWp4DH+Dn17aONtq77BLpBPz+xf/LlmeerM
QhihF/jeazr0lkx1LGZ1po2aMq6/9UJiDHjEWuPDphwYEXXz6KnhGvSoOKAD12vfVr0Pei1KwSqm
QvUGGrV6m12HPX/kzeEEXskvYyI6EfMGYn1oOAah+Pi3ZepNMybOAF5O5to/gZsRTR7lQ5B+Eab6
/IvliwtPY1BeScW5jRHT8IFWFQfHz088VWiVRX8FlVHizn+5hJWIRykDpu7964BZtdT1cX6Hn4+M
ka/PEoaNRVWLAOm5Qa/krgb3fp5yZBHQvF7Hq/Inv3nx+W6Ma8WWmo/7/JByPi/KjeJcyxrn/YsT
XZHoX77u5gnC52qaBnsDtHfwbQcZhp3mAEH3+Wu8bHmsjQSSNIMET8AzT1GToQZsgRRlZgr0IeMF
3J9T+JRdtTbuAPbTTCEc4LMMnSLeLkTNRr0vJvELAJxtk1o2lW7t1250aQNewMH5geyHwQZa6BRA
Q8Uxkk4R03ZdVC5ynjetx9GHF/c6Xk8AHz/11+z0o2HvKNLN7LNAnfxSmP4a145nERaA2TrCy4Vk
iUe4MfhoB4cZE/wAahpL9wfRWk5edgKVxHZuoSieiS6+StJesRUM3X1hxlmU0vpC520KMVazLQ0t
eQCgeVnF0PCbvpKTbCaK710F/lkftlEDg0EOrBD4iGK3id7DGuthsoFvNK7BjFNctv704Y8omult
tUTLXGqV70dgQXXWQIxRpGMMLrN1jXSeUPp76D66O8axZeaCgFpVQP3pPPHVRq016OlkD03+6ZGf
zfjiMLFAWhd1fGbZ4+wXEiuwMqJTVEkdcmoD+C9QUlcVZc7EHQ1JVCz5yLbg2cuUeDVaiu6FX0j9
7dQMd8nd1LCHbDrgqVkANlDeSPfGPFRXx5UTmfV3T/O7Ed6pvTsAOcXDEtKQtljo4IWXNGW+6ykR
bcrpooyDhVIf0m/8MbtZz57vJWzehxFWRyz2W/8H2EqTVzeoO1FGKZrmajimtqFM6XGrQbQDYo6M
hQbn9PG5CDfYBW2rOhKc1v7xA4Ws2S3jgm+eZ6Yj93IcQZUFqFHYzTVLLhYpY79JA+leUXPQh9gP
rN2+QppSLyRiYL6fQLYrcKXLVHSJ41FLYnrxecKa51ucShFy1jNaJyf6zVVw2bfvlSUzmsOdYzHB
hJK6SX/NwqGBbqpGbsc916/EDnxa3I0vHvSphP+74apkbXNgSpYbbepo1HpJDoRObnROohzb7tFm
4P7tJgMi3oViCEjsHfhHhqY2J9FJ8LeH5dEKxBoGiLGxhoWwGmBFk9zqgjvovRuwcHpxX28a7uL1
g07z8jjB9azOpR1Mk50/nNUTKuboLhDKpW977Joko7hVRGz58SK3mrN1nWYf/7d2lPREgNYBuGoB
EQGFVM5pQnXPBYqmIQPxO1SVxQkP106mjHpEFhdY9j2rseWfiT68Soqq4TMniqZuxkqv9pGFMLo/
GIlUu6qPaoH6ZIfGH88iVNPdrOyg8kif0PIRPg1UvS5VW74GazSLZP0KcQstXeJhNCLXyoAhx9+j
fTKthHEczS7ofFVqM7v2+6K2/AwpKClumux2uf7qj8KMIAOnYcgliTEdWxlzWbRYA16qvtz/Jj4t
n5ouh/MY8/pOvh5Cb804K+nB5iom5ZoMIqlsmqn4pPRxvKShTA+TOCwggdP9ilVlqaqMeCVVUog5
aA2bh/Nhg37pPGDX0KhvNBxrpP2J0EpAXXazQg8X3LAmRRD69wQMS9MxKwQUUHg9aYFtWFBGPazQ
rQ==
`protect end_protected

