

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Syf21YU5JnKptD7LOLtaHZM+q1VIhUFTxsmS2r0ofwQ3ushsF40KxXOCQsGAnXjGfc9kVb3Bn0ME
1qO92hlu9w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dY69aEX8OSz52Pib+7B1y1Wvr7162ZPVuHYqEcMQ/oCfJJrpwF+oy+zQI55NVyz5aWKsTxE6uM7J
HbTWuphJFeGo7mzwyRD7dy/8IFTp8OHV9aN/fKWepd3R1nKJ/+bdmSsliOOw+inM7pfx0a3YODTn
FRAbVAMQuwe+OVuT0dQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q+4W/1zvXVAi9QMds0GLwNMATdnR+yvz4Aqge4tYro137XvQ9NhFGdF/mXOn40o0ijOuTLANSGZq
Y1fe5IvAhv/BzIqGLvvBSGadUyLWCe23JTco14xHGh+EcGpkQzSMsD+MtFlsKB5Lh4Pk7Fki+zjY
CYS3IH1yrExDySGaxaJ/xIpVmbcDUIB29ts6Ape06rDNuWSEZkqi5ATlUPCMrVpXs0LgVRBipzor
Mr/lCisQJrroeVDmbpQGOxCT0USTTIePtqKzCRURmGOM39JzikVR3QvCxX3V9zs6LEiHJnsAr/WX
JYHo8e0tsbF+S86/2TJe/j8LJK3VvghHADCdOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jFetHSEk8pl36rsszcvK1lxgvI24/D3eeWIqqx4SgMWK5zMch2RGKDJVjZdo+SXrQZtG4vIfoNJ/
M9NL/crW7IJ+pa4Cb2wH+GD2pA66Yo3aRE1Ld7EknU3x42o8aAXlhcPIjcxq9tmSO5RxnhMKlfjh
dMPsoD+Mezyol/EwGPo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Jgq62sziWqkTYcR9/y/ZRFUy8fWL8zR/UZTwiK9JRpmOKe++dsuUuVffmjjAGJoOkGM1fnXZqKj9
LDnUvlqAYGJAQrwT7QRdCNBN9eBMyr6WJUCOkpNRo5aWbRqVpwZihLgqtvesSbzoaKe4eDRdiEe1
xKR9vPyfNmAnPN1pwf+2YDUftVl5x4CmlqRUCO2c3iETzT+xwYzxqYKolk4Qa8DTTYe9PvjYqn2/
dj/jpAwnTcOKUqpa/3FaAU1zgLKWphnnTU+MOfKNP/ow3ZLVrmyiraKTGZlBmdJF18AzYgHb4rrc
8Z8DuRLa762hnT0qbzjf0vtKn06WBHgWqansQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19248)
`protect data_block
Jp3vRs9u7YOBVBur0YBY+oENuVcW3487Kq2ljwiNe23LpB7IHDytL8Mue8QVIMS4MPpGpBbRA38F
LHmavXWXLAvfDuWbXSLlGd1K7hZhTqy7tlULTZNOPFRY+7A/EuTn4SdvnQjLp0MPRKbX3MRpkk1h
Dod2xlkWLdPZSYTGDp82Ppq63xrKYjrLY/SdqjVbDCmk3Ns0EcJWV59Lbgp3s9MOUUp5ZsmbZqye
Z+NKa/d9jrM5Qsujw2I+utbJ3CMtDP8rhgwl8N+nBwZtFIQ98zFlKijnYtR2OlQp57ufAzeFjsur
4XW27MNo+oCcdZg8s1fBVsTQ+uy0tFWUutMjcFFMcUGnnpwrLBSxMCrGureJWsLrXStr0IK+5H5g
l/TeOXRnoCm4zm0v4ebiDdBzriD7UxF5locaCuhEQuTB2G9KfFSucYnlSko5l0fa26DuqUbT9hGO
IOJAwlwpo59cfMyZ0t1i0/nr+PtBwRToPZUrK86xlp2pnT9HtZ9D73f63RwA06SWeNWD3lb4q/hZ
+Lfq9KoLLf4n+UgYzaO6gjscbNblp2E1IoFwEPHO62OW8JdiNBSWdurtzibE32MRwcLCrfDC1JPU
M5bpLcVloVqk5CQXj8QzVJQz63Aw8rh81kBRfGTnumhoS7whixIak6Ji7E84sWWbGnRnaEBrm60C
SN6MRLIKLxBcmzzWtzxp2f4dadQaj7OOeCMxCfY3iG1af6onvSrjmgwu77Yf709OoNuHPkKm9e42
3zfMk+6Unsex+UUnP2GLKsirxMiM1jc+PzPbXzWxEHop7Zo21NklMHvffcPGxIFE8Bu4cZ44qbXZ
TwIK7VQRfsYDiruTWQHnujV9TcMwwLHmoS4znRFhbehtsux/lqxB7PBGvzMkJknVBEmxF7MFdkH0
cJikOxwc1qQc16DJZ98RxKDhYhI0QCFR42qmx1SlUqP1dU6UqLCrLIGYU5pzTYzTwM5CI44TAzhL
wTa4n1DnqvHQv0HdZV1G6Fj/PvrzYQyHBrXgkmpnJ4uvVF7Vtl/RXz9G+0/krtwDFuZJpHAn7L/F
kM9XI0dcAg+nGb+aFuTXZYI2ZXRLlgCTsz+T90obe36Fj8WYb/LVfAX++vgWTJZ52YWztRgAd55H
G8nf7vjRpAMmkc+zWisTjaNoFd3Ow4m2tQ0rIS1M8MXa7VCAkDM9sp0FX6f06VWz7wykb/PLzL+t
gLaj3b2SBGmBF14U79R7ZKV7dSGwgJbuyfHiJSpHwSvNCgwNwI/wgY4rrXCfWLiukDO89mo6ndby
zQjRXsPpKNjZ8lKFW0bmZLtXz78uzQk7aCWqYZ3CyMyhhMuOVSm7YRBDguYt0icTlVY86Hvxy2dk
t47Vi7t+NakRnuo9ySN/vG7BdvnxNZkxofA4UW08KJbgOlHLJQ4+1bjsZDEA0o+kyZPMZBncx/xO
veNaje6Vb+t4EISStzZo20inT4dJNBWMWjL3TMkyNlP75DNmA/A2C2EYyT9OcaQhmpmkllA1ymEj
CN3gaSbUaO6HhvAl0R6ZkMnn5HJg1egMfAGrT6s/iOZHfKvu7g28CxxkUdw4n0NlO+NGAq3uDqqt
mfWlht01UAKhzEjwco7kMcClpVhfxX0WcqxQkjD6QGPGn8kcq9jlTzf/Jmf4YZHR9wQeM33jYLjE
PzJQozQz5hVDVmCMc80IHK4YDV/EcX3uMvvTjWvCCAiQA549eaT2yLGYcewcAFjAMgkdtI03aRfP
xerKERENsHYXaGi+4zHhYZvzNzvFPuKchTHl0C3atJfadsFizkBdbnxYPu4Z/UIU3rg3Ia6N0iGg
3uoTAMx1DX6ATNeiASnWhkJXbQ0j23UJF725Xn3NP6ma3wtxKSFlF+KUH3XMNdO1KlnldOfBeELs
TvxAfZQQY059HRA/gxFmDttvLndJLROAjZvWjRLH4aA1tHS1bSlGUzPrzWDv4fWAm+UdqtiDqbEz
q7X51Qq56e8V8A3K9DTbe55kxxELYghwYwX5FtvNRGe9jggG+aSh4PtAJAsBrnNcDkuvN+EaQYDd
9AHuPD6bZY1eM3BCInZdAq1R4mNQlKMllGsDDRnUh4IcvUqXYg+snJnxflGdfwBGhO8zBZF4xO7C
DfXsUqICfawByX9NZQhWQwsbALjva1umfecFtLyE5ZJxOH8hU2PiiJW5Zx+CfkSpctYoCcZG8/JI
VWY6gZkkW8JNCbjLFpsUpY9jNGITyfT0UdGmg5yGjMKTXIhaoWTM52giI7P75ToojsbCNg+cId1o
j0UctwGqAA+Suce1fwx4ipKYwjEsoR3xDNSfpEHkLGWKP2bNucUSF31V4oXX/nWOm3SEQfgLQcDd
9ZQV9hVeqxSeT0pBoCkCEFkLhtUM1SUtnDpZ9VK1/RdgcBcnamaxmqd4RjJUHXNEUxV2kimMHdL1
K0gv/KR1WcEBuG2UF6h6w2wjEYMjav37cREIBNtyrPVK9tuu5wur2MuM+sxJLaqtEiJbykVH6vin
uzZx0kWjVE53K0gTn2lVv4W4wgvBJMAyEfFBN5nlhnyrlEUgndnrvcsfehYz6w7/90bjfHO+2QXT
rJICISDDPvsfvy2SqGdiiQ/AIiRyypMiQ+4xVb4opfdZ3HzcWBC0sIzl/SMVDNoZ6FkLTQ3f47ZX
nTWcTBm3TaKvcYrP3tSo3UxOBuO9l0Ob3DId7ZiykOtReztbmmFSaKUt7zZ9qX9Uz3iOE3h+UZ3J
ZIYgOCy+2f+pPVE95kEnlXH7vU9BvFa+PjCdqIyT4SY3o6nLgLO0yEAqBo6UKn7WgCCUR6ySBwus
Q9bDk+2ad03c0PtW9c+PCzbcAV06kZJ5VBzW1kEDGLCPGG0ap2gmIrWBGPCr1BrXZFpJxyAnGjte
m4/AsLksmNDDuRpuMQmb4RdsbZNsybkaKD4HdieCCey2Lv3e5dp1zWOqwyaTSvWQ5MTwSii8FUlF
K7HApWjtFOsOc/EDAQQ1pa97QIMeMl9OZ8pGwYpAXEkSm3c4wPRSl21B+YLDvNXRrra27wCTVn28
DxB+/YMzKZzotvNzjK+bfCowldyG3ndH15vP5jiZRcER3pUDl5ob8ykwr6miVTL2+lS8/gqeKPPa
4mdNdRc2TZZ3oqGXyOC31z6qnv4dx7BlgtC1tAEVdZf1Ul/IdnFoEpB2NgJmzXZqD3gyL4b6Jq1x
CegBufqNILIfP8L78ujhQGlGPh0AD+mKpv/8/NpMYh9SXiJWsONjyatDW7IMnrjwfIJ8AU5PFbmO
xO5PgX8eFzBCV+YYcCX2rQb+hVBneeWj1OTKjFvXOTrSWhMOLGjUdl4AtYgSMIWTEp5vK8c1Mkh2
XaQwDCgAaFAClPR9q9V1/ZVBkHpOYoNg8jYPyO/kx8N7BzgUr6+/GXEiPs5Gwo9IMrZ+S0cQL8BS
VN9xiehVReVDdS9jxHXoupIAv+4APVNZsKPz93KNevlN4B37M81HXKRq3je60WjBuKYQn2zHGQtK
fs0+JaEIDk4ktYKsLqolVJlONfyIaoCBfL50Q6yLU2pRAhK4jNOBu1q7ihxtobnJ3/X9vcS2j8Ra
kXPY0Nq++ZkVC6Wo8IlFYqUMKYlf5TMt+P9kJnhGYBBjx5R/qdxVIkmp5Ijcgswycm9rziZpymvE
nY1vYv6sDRhfKAkc3OlENYIoluuEfXcAxMpPA5htkMUas747OiuNZ9Cxr6x7YT3aZSVyMSBMS1QR
tcdoYIqMAE/iLKEom42SsHN6hUT6cI4gWLGeo9QsUC+sz7y801r0UUOxMBQD+iMW+oV/PYCRptqz
wWYP02z5kFZlEo4rzh0QrTPEzYVRmdRoQYVApmeNEuuF8Ks9cABt9ovad4BafKKOvm549XGyNJGk
aNdCsLWGDytiRWfphHVIMIdeYKnjdTQ8jLSiSjI5TZR5byl78bNWANFKmK+S/FRL4RmQFHJ3PgGl
G/qnrzhwCkBDSivEsK4Eux0Z9N8BTntQMn0W13irYEu5Bkna53xql8ktxqYrY+dnkgEh21WkFXV5
wzn4XWMsjUvO8qq60kJXpVjYKzIqt0T1rnMG9B5B4jn09Oztv261WRXAbjeGigOasl64DK/W5+c9
0sIbN7t8/847/gc2sZmqYos5EDOxKhwsDOEynL1DQChXqwGYj8Jxv/SuB5mx0hvOUN545qxGUtSs
5TC8Kry3SFE811i4zqHF9KyxjbDobEf9z8F4Mue8Y0QEX2gLRBJ0iUzr7FaXZArpiMGmxKuveL/7
qBVmwSw255j7Z8XsYP2mhqLiHG56698uuz5xx6qhgPijO5gXt0yUPTItZ16pjJpZauaZphquUZcg
DAr7zhh63FyY9dNizcCk3iOQmj/hGJlKQ51gQLE7t4991q8MS6yLtTTRZ55R5ELD7OTQZhyt6R8E
nLSq6L4CNiuxS6kUDYizy/eOEY7uheVL3uvF5HBJLcMO1cAY1lnm+GU80JbaHwhMPvyf19GemGPT
Cq9SmHMJeLnL+PdWrRMrY8Jkukqh7SqrGmEBc7fd8j82nYLX6MfKP1LcaHgZ0LxgITShW6twGfdn
em8ga39Sqb7AZR02AghvswuM0NpWZkViAwwJ1mBp2jNxj3jhumDhkl/7y1Sm0GDql5cOFIwvM6Wy
Dqtp9A3oQPiuIhPfRJfHk4U2fqZUjRvsHXObSVt5BpFMyGDVA7qiALnF8+BkYiIK3KQu2l4qxGn3
J7qe/xbq5ctY+ATvIfsEdVNVsezq/0dgt3AXk4aLp0iZSugrwk9tx/8YvdTWlF5p6abzx3lne3WG
qu3H+6cCvdK+NtquqbofotORMQrq12Y2KtIz3mF4nH2qI/AA08tyC1/oDkbTrQMBSSPE3OW65azU
+6R6VhhafpW6taRc2JFrIf5s72hItUsQVsqB+O4yWlymko07yswPbWzgSIKBb04QQc72777uIqZA
hRJfWvl6n5VayW+AL7Q+Ez9KViDeiYRSJ0m9GsEqbxCsS1uNRuVXyPsY1d0/2J8LKkKBSuxmS1Yt
oWHjN0AP/mIcl11LdtfZMDvePrDikzeHYH7aDnROJNltUOkmbBHWylJdE9TNtqGoy+Ymwy+oeZWP
nP8LScpeE13OpjxhcFYXjcEgnjx0QiVzezQTe5XGwFhNaeCoL7RQG9MJHCgDlfgZgBFx1zZc5GNk
JSVDsvL/KfcXxCD/tHOGhsbpghmoynddmw4cF89WAoH9/VgGYhZ3c3FO8C4WGbVpw07+OTqKc4Xz
JYJMQJ/tkE7NS/VJrMtozC+ueGEErea0M+7KfO2CTQxpOB6SwKVpqf6Gv5GIh4j2XUaoDE/BxFAt
3McEiNwvWN33pEK9cR6P+U3kmtmt4U255Wo0g4gpPYg24y3wL4N7VBgACzQLL1a9aJby+yVygEkW
k76MI/5yQzDcimim9YpcOl8Ga4vpn53ylWd84yyDfGiRuikruQqlNsHOEsw059g1E02XU7ZoTM/p
e+qRkFmCypU+38XBF9OgyhV2TeURGYsDQHPSsf4TpGdZ/UDJ/dHqabBjVEPbPaLjt3SygC/QtT1X
mW7Athau3AgbNKcuXv/Fy/NIyN928rTZ4EcSngPrnKDeACZWM2fKelXoimgMsxbrg/uGZeeQlpC3
ZBfTKCKH8LaEtRhIPM6Bp7tqEkfQ8rIK1UABtNXxx2Ka5/0o30FTKpz6Tt9P17EcJjqJUD8jGiDd
q0RR/Xk0owphPmBVSdH1Q9zrhrEnXACMsJCuklcIzF5UG2eh8yh118pTKq1LbaEgb8d8TQoH/Kpb
QuBTtLgkquOUTcQ8HaDP142HSxDVoC1JrM/8bcAwL+LRxR6iC5Nn+DIVVIx5wUhVzA8LIrN85CN4
D6i/8JucydwhjqzV+ruSsp2Aa48etzVtwC98izfsGFsDCBjo85c77H/ys1Itc1VfPDOouz9HcbcL
kEMgZUpmrCXOYtnCzEQ66T+rfK+pLSiyC9PhC3oU6FrTxQoQTZdZiX5MVV/rbVqrixdpz0r5/uMH
tMer7NqGnuYdSZkj/BJQfvd+5j723Tm2sHXe4YxaM2MJsP25beaSrg4sopTboX8NBN7++zwZt6TB
y0XaseQGT6z1QMsfT6nXHuQDZcptpOLzjsdRszMqhQ0KdZyvxeVhECjZMVbFChFjXZLkByg7mj32
OGs58SbfGWD9pPedwYSMM+ukU/QO+y1SP02gVdu3u82x9YzBMBErF0TKlqJcH/9GPJk1MP7kPjqg
8offpsEjfoFC1lpMh7YRra1NEFv890yA0qj8FJoB09kG1Ne7ac98vRNaPhaYnIXra9kYYJ8GgZot
Xxyz9YMUczJHSbVWOUcaQCpNR0pLYpVU/MqBBB7zXrDSLG5nnZIOX+Xe4/27SBJv8F73cmXIfw7Q
NtxJrFUv9qQBjQWStWnNAB5r9P/ua6Ri3oIHaBRsiTqyV+q23MVCR4fXWtCKKFoPuG8GETT4AUpP
rJyJyJIfBNRyNEP3Ou5z/PndTU/AJRWZaQ5CyGBZh1bpqc9d5pv/Wv1UpRX9TFvqzJlq9MitEHaF
ca3wlzvGpg3sbPmxSwzW3ZmBrYl3D8jJhKbdB1ZJS4XyQSn8aUEvGh8pZrowdE+3QyLc1yFqY7wV
eAQ7u96TXWVxt9E42W42hfbff1WMBN8qNOXgHW+1/FzRRq6u9nvHj6jGpLZLDzqExDHBRKXrBK+3
nX6QAb3vzecAoWY1Jx3XphPevb2NuB+s9xtT8mSrOa6XsEWuoH0CwuE2CTDm/I4FncgVnSPTso5m
c/KVXHfXzOgpOw3GmGavw/rgLKX3nnYrIsxuxfAtwHuoALk2kDUPUhdjy+hfMJE3oYDgVwggOYl9
OgKaVKzoxSazQryfT0Zl+Il3zJ7AjG9Db6p//Rg7VyP3k/lx/SfGB8561U3xyg/a74Lj3RKOKU28
65aJPjd5pKH5f1FO27muWklSxk+J/EGBACKIIlW7kYCMVdpaGMxMxwJ4cVNU/VOqfIOmvjBigNSz
kY13ddBoTv+X0HmXO2KeAlJuCmgk9bfO5yDAFumYJ42y7dne32y6Euv4MgYCYHdR6+MFhhTfqlxT
3eMUCMhKAWYsY/eS6y4eymItE8pSqajHcmgOz3dBm0RVuIneiFV4cJIYGdCBRZeMDUcm/1aoXNON
DkZXwq+t6QYocltZC63+ckBOqeUN+xhzZBk5Z8YJq9X45so6GpZotv+mjZQCzOfPWuWWNxPSFcBZ
gA27/hDjq9+NqxYDE8dhPJme/LeholtL1ocKal55YlAM32vmlSZt2NDILGUyIsbpyI2NO8/y0izr
OLMcIS4lDJVLV/rjzKav12yD02y1WSmKWOIQxo6D9LAskAb+7zDjm4mwxzFIpx6quUn5srgKXG89
GWIOS+ajpYhnUvKH7Xmo2OtzyEhCwcs5DHC3NE2ZDrKkpI2B2f980Hx/o726FqPPDNYglnJjLjVc
sI1AAnzlzIz6cpBu8KJhEgTdpbAnBViDn1ya4SjC2i7BuaL2X5cYVFozv3PLD1wFfYyPnV90fu+Z
HQyd5Nx+wZ/2ek3aPc08zeHcMcfOkmmG2Kh5QfKpqgKWY762nsShwYl9cUGvSajMB5GtvavO+bkb
Y5Ide2VTEsRZqu7aB69yIKwoIVImiTyWui6K1AkVn7YHLkYmTcHoJ7aHcOs8xyL2yxWHi7dn8cRm
1PBVNXYOmnRGqlTcLAkqjcYY2tBy9jwc1pRuEkI5eu6fGCHLzTYXrpfvdaeQKbUeyqcohPbOANE8
0ecpAL9V8iRWgxpKXR4QF6jiZ2ZxckCPaxqkiuYWxa7GTf3Bt7AWYmziMCOUovHnGfLa/x8caEQn
ywS0hzQnTr1D8c54J2ohnOsGGBXYko1piATpnytLuiElR9Mvyu3l0Wp41lPCs+UQX202QzGh2kI1
y86iQ9fZsaFivtOw9xDXm9Z1nUm0h7QouUlE/cXnckqG0lFRpgJBa+FN0i0b4knigJBNUg3xJ6LH
Nup+bZp1IWxfKVwvP2ho7B61wk/gRsXkcBibloB4g34046+E6NJY8MbyLymUpN0KzeHmdqkkJXzV
Cm2mBkIoY9gaQ5DJYcJjJwP5DhuiN0tJm14n+OK0ppU5jm2sMYQniIPpt5myYau6F8KKzkYUijka
g517KgXTgaZRlrjUtbcHg/Q6Vh9cIcizwjEa7qS3kEeKgpklSN35lV7BljMC2XKwJ20w1JWltiGB
VTw9geB01jrPOxQH+Ts4oWJTtV+o7jF8uSvL4csLk5bmUbgeinWf/ekxxBu8hQpdIdRmXMkyxgJe
42jxtTfp2ke0cVxVHk5qcee4FpeGHOFx3VuyPCExNyVsOCPXbUIhHsB3ngW7+Uk9Og96C6IOA8Ip
W06O+4Z0OJkwfcI1/gBgkmubkGGGR1J6jglO0YT5k1iggXhiB590y/WtbqczTMwj6QLGjk+rSe/Q
Q59/N9ZRmyvn1XfqFPtwsm07u9cIfs6P2ezon7r20YN6rXJ0oZFpVwSGfENF9IUzygONIiyewbXq
zdbmC52lf0rHrfg2sz7s9wYurvyP3qLKoXV+Hq+H0uNg6UNhnjw/u5eNEXm0i3u8AjuryD9uGg9Y
tCe0glANLQ5mg9Lf51jdBZaP53cAUKc0XyLOvGOTjsuCSBt1tRoI+N44Yc/llEF63S0cdpKz338K
lcxgqi0kAQ5GxMe1t2iVZziPL2eB4HDa1OhGvKovd1vUXudhl8ts5DWOB2K6NpBwbMRxC0dF+ybE
j234GIja8PwOfVnze//s/eGOCboxuNhJLuqs3wnDxDq1CBux+c2ALF5ZRuylDQpw/C5yxqenf5gm
vrMV1UYqNqYJZ6f95KqeKUx947sZ5nH3yDwI8Hg/t7qL6VeN05dzSLVGMSVRx1x8wwvZa1MTyjVX
E7QGQ4Z7UTsSi8uqTzRL4xdZssTkcezNiQ6RTxGf3By8PcoaJUyTxqEKDLITVzQtUmedRKyO2x4I
LPB3sdnKvEFz7iH4kNAs5ghw+RLmED+ld2nPGkC700vdXH3IUxeo+gMnRK82I7XUvqNEgPLJqWbA
RE2/r+FFqtzP+SSEQWX5NvXZ+o998IFdQ9HKsJj+VeE+xOI0eHbQUMJQnIvU1dduVrc96JWDc1Er
2arhzKSwyl/O2hgdEWQ9nXZKS0VN66eufNwEiMhtsQbmofbXDxeD/gvxcyVgj9hxvCrM1iVEmmam
4A4FUMnOZFw4oPkPnuF6SIOOIIew+tyyt8YCpytiHnkswb1oXPXB5sN3hwWRer/ExjSYCz5Ft7my
A1wKOSxmXGUyYyVwqlgNkX69WeajpkiGtBKhEp0z0lyqgHAZc3uS4Y40tNYQnVTZVP8SdefP5tZf
1SjU7aZBLkMvt1hfyIxv/B3YAXChlm3uAcNJ4hGGPNB4MFUL/Ji0mvXxaRkKOUnpEA6KzheFKKHl
x/Qpj10r9sml/SBLWsNR6taiQd+dj5FCjXF/Ol3rtU50zu/ZjpYCCypSlra6WHD/PZVIAn1KSSt4
FfzjELGZtTz7pIio7p/dnYSCj91Si6/HqwKS+MJbhWTMShUtZEOKtaT3mlBfh+in+w22/YLCKur/
VCPf0ujk29iGrYdso6sSVXkseKzvpChGO4m7UWu0sVl6tHdfwOxxiBbcjUVbylUSImr+uPAOvFSw
Rb80pZDSdgrpWI1rxhd/yZOmoKeBN/caBFmR0a1RBnpxoJaNK52xVc7fAxeKOIp5cKBGJAWhIjQy
IwzFzEdp51I2nuIJIIGfJlGMEQJhxpmsRJJ5BvvayQMmNBEo7d35bZ5/mYCe0IlpyPiX2zLAn5o/
l8gIZoS8b5I8chyoWO5CzR55yqEp3Bp+9MQNd0UIZBcwozn4XJORxP1YcpV0gUNo86slEwfnD5t8
vmtWS7Hoq4jddFOajUP5fsZnU8iYl4DdgdPRl5uHWQCmd4LKKXykSnTXv3EL9C0E9SaEeE3Fymjm
u5yi6Ht2AaJE09Iq9cBlaxRnBc0/ll3lKUgJ09c8ux/ttSnZbsVgJQGe9be2JRijYeWDq3Rclc0j
Ls7foxue+Grg0OFO62xATxPZUPejXsmxUqO5/3cVIuEuPIK1uV0/mQQkEOgE0o9yTMEN+eNDwIpO
NczbnXtIDmyIVIVtfv/Z/PPo2mJ5zyefUFv0kHAO4rDPvh/UIHlGBza/urepRQ3dp/dZZlvmA508
Yr3HcyLxJ4JXSV++E3zm4WQx2My/B6kpDcaHVAckW3hEGUzecp+TD7lahy0Jrz3iQEyrVW76TLdd
Ybe8THEHQPyhkdy+3pkvJW/Sjyh1xmcg41YpRzKlLlTXQWdaoz1SlqY2FnhKv7gdKrRR75YMVfne
5C2rV8+DAoU17vMRL3JsRyO2pIkvHVQRy4YWMRBgZIHrvvCb8BIWKBtE9FZdefwyJipvtxuMp3yJ
zOBIgjNghJORUepB0L4j0vmWkQYON+bRWWEVvJRLM2wy224A60+JP+jNgO9RgJzSsylMUwt0WlfG
gqYD8HJUub4hFUYOr2HatB9DFILMJhIHL+8sRv2S716VI0je1cF135HnfE4RmgrQLHYxMlkNHXrv
QA6rcFIhBorliJdLqa3di90yPirQVcZxrzwnVaZf0WOkEx2JNkqLROC9N+ukLExjP1nr1OJ4ldFH
JhMHQ7V1dicmQjVJYTJEnZSlFfxe4dTWL1xhFnPJY3r6E2IebRBtbnx4oPrpZAXdyfmqggXMI07o
vGqsJV4atYKSsEq6qJmn36IpGCRjA2CM0gB14+tl/APtz/ydBvSECknLM7G2ZGpWZiFFVGhmp2wX
VZhpqJ7EeL7j8nNJNcj+1rwMaguhm/u2TD+piWi058AgxwdVYlG+jBT+BhI9pigYJKTOcBc0Y7dn
OG+BG2bkwO5zjGV4wuh1XzUsW3JmsVbB2sCOou2/KOiL+g+S3qseMjfCCOF/TBRFIRwc3M3uDXub
x+PwiSYJuTFGXhm9ZK50tp7SoPFm4Mc4+18XYgWSrtjnJ3wJAXVjjWurXUT9yKgKtbN+DPsdc2L7
MeLgfi4H+TE6dgaz+iC73VI38BaMZjbMhBj5+jFGTSkjFL7DY+fVWGfA8BmPGpA/aff4h8aZuqgt
d9mup56JBR1KVe/TRKbAZFgbO63G5RYXeXIKfDCM4SKLXbNILWQ9n5HaTXC7CxQCH03l2tH7vY4R
gEbUEsRn54DY611Mo/TMjsIeMsXTiza0hUZJRUaWHu6BcWaRpUZLlzrTxN2iq+oW65N91CoAg1OH
+1r9NeFRuu2JPQmC32m6LgMCSIybBiyC2srqeADUQnLXaoHakb6CPp78QYhKlD1jOO8X00OWSLQS
/gaIQidVRUbKTuu+gNR6esVW0/oCqbQfqwGUxkx2+9LqLalDaUFzkhrom3zD7OFe2EfHIOIpuPIu
dyWIEPyTpXl3C0SRU+a8EtqhsilePgCY4IcQDRZ/vIZ8/RwdBnZbuq2Z6HYOL9VP/4TmZl+4VRNi
5glCgkA5QNrNDTORAzJrvB0yoAaICIVXsKhl5n30ci0Qvon2Nazr743HCXvio4LyxV2a8eUG/OT/
nqBP/hQMQejhsYIZwjsyaGi8hJfgi2Nl/1Idu03XWiR5jCpgQzwh9keYwU3IyMO3XnfsoEExkpIc
jIKUdQEkxV5dMRlWSrOOw+Gh1/md5S+wWS/I5YBvtSomusK5mTr56f3AC+KjdLNbaJB7F9fPO9M5
wMOERgH9wOUtrFJfexcn+cDCZZkr1d5WSfGjHMqnUI5ifX94p05b8jUtYsRj/zrGdK4Ba4CnZG2f
/CetgLiF3FkQ/PxBDjokCapMucFBjsqrl1iugwzNLxWd9Pl6EVua6uyOYTUa5j67dov696P4Clq8
pgD717mZvESefcbYYXItNvDbsH465oMulTFoMBo4tC1vaNReKdglaFjLxPBW5i9bxqzW0d5ANxNz
BBzC1hO07Fq2Bf6m0mTJX+GfuHesK+54NP4fMfx/3dDQmelCrWW5HNvzuxPqwsGaaQgn+BRCzk0s
TkjBtZMmwPTxHCAvdkP2cTXhx7w0QsYj8TQ74REqW6TiZIKiFc+AtWbPxgIdpYxJUifsA2sIRIUI
scupILsld9kmT7f2E4gFndsTXj3/K7MXG/kIMfal3No85NGoJGawIwAMwul6F6K1XTzO454clAG8
C4UZroHwTKIOp71BywQ1lAAhQMzY+yf+5bPuoEE2IAkePYHAMB19rrYhvkWWmVdVQakZ13RpiL33
QybFVn32ZuMFLysrb8+2kXwc5NXE6tRUCZ3zRdM2FUOF+6YEJThLQuLWFcZ4vj50+fARGChya9R7
NxE/v1ZseADrpSgrx4WnSdDGJSX3O/5ZBEd9qYpCe+knMEGXlzE3Ggqg1QgQqw5DewKhHjEfU/4V
esfJgSyzWV7w0W4eMnoJIizBgnqRRqEOtTyOhGRhZTYhEB9DB7CTcTYKiO9OsHdAjbQSZdYK/y/o
NcRXRnHVInSLQyDO1c+txjcLRSdxEkqiCEADLo5RcdM8PeqYUTDMMcwWZbSErNs7gOrbRlLAZHaA
f6bZ6rQHtujbkgnEgDSMYCU5c+GdKz9sQrR7f4xT0v6jOupmMT8FCsIzOj81JizpHG7oqGOzMVDI
Kam9xzAjppRfHEjgmexc3SelcchA1ovBdskjmHV4uTuE3rFUoqYkAMLATrkK0p/D8bMOKk+7iHeV
fOIusHWkgdSJuykJ15pBa9REcNhbKW5GfA2iBouM47ho+eGdaLUPGbte36P0SVqQORsjSJhcaYUJ
W6v10ljv/FPqTDwcRXHewM2EhMSr5lozjEAM+IUQJZXirtG1jkKGOnaXx2AgJ62BKBioQvsActhr
XME8q85b+IADas1EUXCj62nt0o30S1MzWi0HEORnTpOjeLj9vutIOQdXvgRu7MFyYDjW3dqcy5pq
5SJ63T/g+SBiS5QL2XMPTOjYLrg6eqHAqhmV5xziTv6EDcrSIqpJwcbzGZdwL7ek8vZSBzF4Dh0x
VKq0q9sj5TtqukeV9x2BaHedZ+V07/FPZtbKZmMwjpSBOk0BDiEhmBAm6XXG5ld9NcIMsYI+Bugu
wWzvZWI0jlSwPhLVA7ptXWEemBqdwpP5NK47P6oZJI3gnupUhLAjoE2P7iCVsu3l+4ZLXSk7g/Ki
Rq6Ba1Tsz1zVxfOju485OqtVp/chRE8GlK3dRtBRwlWJ5GVTEZrq7y0fHsy4SOBzARfY4S1/1wpm
sUWFu86a8C4v1gqrUh6IJMfWfEYzors7Jhd+w0UG7BDg8B/CgUz1TtT+pZXnLYbxt6ZZa8EwtQHA
bCqXQ51qW6RzWw40Cin89l0/RZjrojc0PMbwOTAZZuyZPxZi8t8XFx0jACPO06ZvceW+OInI86/x
1NpSliw/FuvaI5M5NJrprkNNGKpqsqVrAOuY7jFC8E1l/cbqATvyHrsQNd3txcSFxKo4iq3AnmbM
1ITdujH/DgfxFWVOa37C4Nrp5dbhLlW1yqUEXB4gpNX0qdGMQm8zrBPGTBp8CLfqvvP2I/KPteDv
o0hVdicP1978h7MSBvts33J19Sav8Hsb+G7cMIDb7X2EDP2n4KWFL/L2yBGaxqZPzsXH6jkZehg/
YkkL909FGyYDbtRLpDF1jFzQ6ofIelBATbaCZl8yTyAyCarg1X8fvjl/M45Ad5h/a2eQKfi0XVjw
Xsw6fM3OEAgMmPFSE/toUnwRAFahNfCvWUcdEar4CDZrhQVOS+RULVobWdFCVr8gdkWgJNd+/nTz
/hYWrfHvASAzHJ/bhqrm/WNYCMET1TFyLLMjNPlbIKotiAh482azIwdDIv2A4tqIlDoZ6RyQE3UO
yLpgV4DtutmcYCvh7GXsQW8nLJq8P8Lx3Hk6ubLtw0GnRsMY9PgCzERh3YIpXOY0VjPOtV5TrzoQ
07djqk40InYEHoLSl5xdpBuaH2XgyeuXcOknZHjz61Ngll3ps2LtFv39cn3rUlnNgUi10d9JNStV
e/LZyQxd+vUQq4Ip+4vSbfZGcghs7ZtdKOVxVHcoem6duOzxFuaIp6T3iSU9/BKNFdZ/FeRST2lL
CD8AMF0bsAiUxoQ9LI5ifXzdxbq9gZlFUHK8xWnt4K1pByIaf9W6VP8F1gfIJcpwZWOgv0wrQqqZ
tb8r+FnUWcURtdi8oOjwCbqOR59QyBvQURnRsR3+IsBZc2V0136w9Y4Rfe8Gnl11oYhQCMX6d5EW
U89OSmk2dHUkIPky497mEtXl/nG+G4c5pWmWlaI21L8eXeZbs1k9Pq9f5v4yckaScI+Z6Xz6YgY6
x1my5cM3NrY1y8SBZlRckUVlGKQuoCHTM9li9Y1P5UMNVxKGNEdhG0V4uEcfIoudp5OR4KfnclQz
bbeI4y3I6SOT4em2YhkCQx4yAHdk6tlMDHVrfBrGIZyP2xCByKM3MVIfnB0v9qE0Rl4vESQiWWG3
qRQmcObKTcwOq0ZfaFrNbvV7SU5jVYasKRcq77NFJFRrWmKmY7r9LK1rQb5dRAWwJLIPTU3QadLA
zHz4wS+Z/sTeH5SF3ls4URMFHBXGNDYJlTw0eM2TGch1lcXlXzToXtdU2LaYHFHoWicYVKqNHYb+
NMjMusTj7ITvctOGKrjdwKRBX/C0hFOdh9K+SholEaogAH6BZ4XxXJkZhS9/T3CturVMXV/EanV+
BYq4D0iBPFRclXK0v0QHxTczZjvKo6EAuVviZGDBdLhGUo1jRoy6Ka3e/PG6mbxnup4YKgzHSP8O
S7+5nNhmhme37t/LZeVMXVvMcXBwiBm7/7ScPtKQH8pkgjbQjxEjO6PL+mXok4rz3SYjfww1inMC
pPmnz3THsq3/L/Ro2FmJuSM2Fq3kyEWx4Fv89XbxMx1AwPXUGJor3MOMOVoYTwfDlK0f9Yt7tcP9
Fk57vgXLiBYoUmFQGtiDQaeZOd3qYFT6VOA7Ah63wEFRwbLwKv23S1IR9OezPCr6O8iyEVXIJSNI
nSkXGZpsLlSkrgZRSkET80e36n6CipX63Q7+aPTQQxVMUDrywpg8QlmbbVQ18qF3PnpZtTdPfqfk
/sDqXCD/W+QrXsmtN7BTkbE4PlMBblTAGKu1UE9j6VFwnvzsC8gWU9fx835csPsIjyN1rhaZtKLI
8Jvc6nTzs+SRqK9CQu+EVPFx4hYHNFiPmvw0GaSedp02N44RN2iqDUC0isjpXnIs+E/+v31zdRY5
4/R+eJXya0FWGNr+c8vGhrp1cP4HKYznQI2Oq2w72nbzB7yHDwPXXRT7FoofTVEZkydCB3iiG87d
/nORN4+rDX0rs+e6o7jR3ZZsmnnKQKWQHHp79z8Pt/9kT45oBejBZAfNWOn33GLFfOY15QpmKZNz
eBuP2Tnqi9YQAp/FZT3RpRaISyNWDS1TBedsbludIlf9kCBJaH9VTgpB/1H6lRUbW+40+NaOjJmv
9E8jTb5YxSS6AyujehXQ4Ro2NI0M+Ta/DpLHsmWQiY9azw0ekzI850G8gafmdMttF6CsreOazfli
wj0TndpyKuUIVRQQTqMUubhtzkUDAwR5ZYt2gEJOwI7CP8IBCexBw1DqvzWkLfRtbEiL7MeJbc2z
cG4MRf6zbr7LS34FQV+NF/1SpQX+rKQT2JdKHCZpjF+CxG2kLZh/57V6I8mZGrxJM3CDD+Sb44Qk
om0GmjjDqpEHKG8YIkTM3SoxHwcCQtT6xtiFAPALbfyjQHkuC/dyiUz85Zulefl/C9VSyA+Uv2f9
0YlWSFqMc4IcFty5Z487f2LZdKwe4HUKxZF1ii42QlclOAGC/brEEa89ap7xetguqGjHOjhUJYUf
oKeBmXNC/q6hQmT7lHyGMdg/K5v9K6D3ZyagZWJbPhB2Rkl+1FTG2xJsbfxgGe7TJ/PKaZmw2N4q
kqy/iwE3XIdBBLmWWPMBUmvSsMmpEleZoS7E9TcTP/5ruHEDFiOKUlYYEGx0orQSFsLkfYS3hF+f
XB3HsUdCIxacqhp0qAyBlSZxD0eUxZekwyzLHWNF2HCPOU6wQnVYejve/80UE/qht7IwC0MHlMJl
Y8c2f3U5CsxVtYl0LQhmO6gBmPq5sfniu//DwfqbpDcJzGTbBAbL8R9ta16NwQ39NCqFpR9UU+DZ
ed4ZysNqgXMvEqJBLSOp5AqVCdWeWiKJUwIlFjbqoVFIv1G5+EaCOLPsDoit2x6PqQpbtGdhFFB9
Gvc8PeoAnHvyJDLizqtwe2rgAycEu1I3PvY3AfWCFy6C011zHqKi/2k2exfjr0GlK3X72kA8YGqF
G362UIOa+IQ8K11Rk29ysPhbmre0DjRzI37fh0tUajgg8w7Hf7NBE6rShEDfATz12gACRDliUVzF
gCiMyMuEEFJ6guUZoI5CfHrlVYNqZk3D1AP+wDtxNiyiOlwuVU4COj0bOaKSisBT2SZCHvnb4o5c
wOnADLxdG8McYv2Tm1bqIYMxEVMed4spVElsdVsbxLL5OmM2e6rEhG113s2uEJNlrnd8an4ZaZvf
XXOsNhppYknnfzj1Qcs60sWyo9bSltOdlyBx7+ThOzvsUG6P80cY4uz/wTxpbSG5viwMq+U76QIl
UUVoqtdBRWLdi0uYZ3gMfMLJRZzE+ytyc3AaVosesjsfilH7T0oXKFeNO5OHyyTwnUAhIDBQJXof
tb+OM9Lcr86mmY0OBy1DBnVL6ig6Q4U62CXKnKOEhx1rqFEcD4SwJt0lM7ZNRZGlnCZE7nr9/jAg
WX+vulhrtDpnGaTklDxN8k4Te7njlOQsuJbEK1W675SYD8DgTxecRde1JCP6b9ixXhe24WDyw27X
KctuumvsvxWt3fhy+YZq/iGPZ4u08vPjo2Nq+bCNgMBTRURD11FCX/tyx+20ZJJSBlMEKz8E3PUA
zgSGVBUDFAj1QQ6k18j9BPhYZ1wI6YSMg7nxROMOKskbg6Qi5dL4LTA4vXLVho38zfIdaPP9lIx+
nyabVWGUr+NrOUX57LpDH5ypdAQoCiQtcCJdjX5pKCNQ72cj+ZIhJeBNc3vj62GonBCjurdWajrZ
gVXbnNHpqc3lwdS3elzJXMg2XzShdnWaHyYvLXWJujsTYMLDr+a9W7GSuM4tRbcWBlIKPyu/FuBA
BgpuMtzWze2EXcihVFZCNNvWJe4SqG3tmcMl57rdiOMxoI9RZxJOfnMiJslSEUDtNLkww+MAV3Qy
XwG0SlpxGJxuMEbSl5lM824OnYXIp5hoIZyPvMIjaX127mz2Xobv2aZOz1KjcxzGk6vbJkvabpB5
DqoSCXHnK7p0x9ZmsbGGk4P7jGJ9tRkCkKzqh13PC/QkaEwiOsXEwbSP0iLk81nh5BHQHUIchAIH
1MGyTh9+6Or7OQRjZkKZRZGToJcGDMXBa57WWrhKys0Jv4V3hg2sY5Rdv/rvM3YvcMmRrKJuXfGL
xjkkxhjYd4A0W1wcDbFpWQ3qJDsp4/mdQ3A1qg62LqKFYfLjl7him8o9EihvQKbdRtLGZHcqCxky
6gL9PwM6Z5YXiffKTK/H2ta3XkbYXQMq/yAl147DvZ3ElNzfn8+XMfGuufMrn6pjvAxbOa6GaqFp
Gj8C37mHO/0Fw37Fe0FcfISMx1Mar7hxYv6HQ9yC5F/n4JjoRghY2fEFc6Pfi11fXY3ypA+sS5rD
pc6PiVgkFRWC9OT5I76uOZcLPxnyrwwjV0NsyPZszUuunKCzxWKHxgbrEEA29WpUr8oco0hMXZ5+
P9b8FWufYsLsiOAuZs0CLXJZ+KqHeMVDVNQe/xWbqZKU3IYcPVrxuqLH83FFX75/hFh4P/z4c6oP
eypQM+9B3yWb7NGnvakegQh3OELoaaLS0RVJkQjcbZ40Wd3D4oLC50Ck0pM8h4PiASsHCU2jTi1Z
yx2UTj6mFINkffEPfejK6ehRFTi6GVAXgNxua1DUbLthvkvGU4G+W9g+VeSvMKQuPBiu3ruQEsM4
m5QU+hKNFSFAzPbyIJoyIhnmBFLjEs9Ny5mzySyNQ8CgiRNU6jRT+v1phbBvS0H+YSN66Sm/gtzs
zK3cS0MHdoz6SeAOfx7/Ta/RRhobV2KbHj13R2gwU+02/W6mesPxINQkkFfE/0FZ1MYr0jB6e0g6
uinxTDrg/7yaoqlHCiYWI+cYIrMQ9UupbOao9KwKANUJOjheWDuVBfeZnuqwDDtofcUatW+JnuV9
U77Iuwxo1/cxNbAMu5jYGm+Zk/IC3hsvb1BpMisJMnRsYLOZ2xjI3vu+qAcZ9JXHsu4ywaos2CIR
pQdWg1END2mP5v40UOn7XX2KW3c9VBY9fwqAZIAt1Mop7DmofB/Uir1GKzU9MQn+EOOs4zxoQwLp
zI7eD9z2zRlT92oPJNOAqHE459vBA7ZiOpG0EC5/gtkrxU7RVuMT1IUg9zJ0La1S95IddQ2Fm4yD
suRLOl56g065WTux54u7e1Kfi0+JfzT0dv9ZvqLbsZZGlCGM/yydP2bNAIM/BolFhOqhMMDjwi20
Yx9mBRnhIM2jtSVIGPwAHjelHPVoIDCTKh7pBWrHIKm15A+QZOVyNeLJoERbmWu+s1iwlXz8TVw4
cdsXB5VbLs6caQ/wo/X7y6K80dNJorNABp+1nnTIpW9Htc/CKnm+r9bo155bUPRqsgMI87hDKZgk
9GlhbVYXhkRRiXHgZn+KLzi4KQPr3utfiBUSzf4nfngtBZqUUHrIJd1Z/Qrtr3FaDOTR6Iq17DVV
vC+qnrUoNSWF79hYV+budoUoIMcNnpPB32wEiRmDKARW4T6uH0ZOM4MMUjtdRmJu7qq4LNhpM42n
ey+O7B4nFuqoKSLPS3VLlHQRMKF2bP3Ql740UYY3hdD2rjU7e/Kkpg8U25XpFNLxjE06W7np8CmK
r3NLmg7jzHhg7KutG1VLVHLV4yPUWLcYbxBEUaNhF8T3wx03Xj3G6Vv4SyCzMPJjryKWG30oQpSi
EaVgXaxxz8Exe595bC+nrnP69Uz2sjAVuxn8+Riyd7WzKpOUoChxHWpdyJxU3L3eoxZx2ZpWEhxe
maHjRh7RFGwzzTr/PlOP5+zkv1Z+dBySIbNAuAIRxiD6e01fOfv3p779UGsFinT569v1qTSmNPLQ
nGu6p1VE6vhYq95wVpAdJnUeDJ4sMbKZE8e1B3QyTFT6PMvyhanOST+n2/QUaIUdfzrPM4HRuZ1j
JIP1kFYL66ehVhMj4gZdA5l1XFnl9Ht9Br6fd3XOiqUTirwFECRYMMgMMFpHYhIfwJsvzzAXt6gF
w0Nwdx730ZCBQ/OuvCErmxzCejZRgNAasUk6MN1JISX7Jo+S2t9ta0UGQJrn6N78j8kWd+YIbB2T
ZX/TUSHC7tX12NY/W/r0tHgIHaEwY7S67g2cTPuz0YAzkUv5QHybo+DBfMbbZPwOwU/sLADdtFyl
Dooi3FLyziUEOLCXBfEZunIZodsqhtlOAWA+QI21z0bIcaaHIXclZlAhH/KKHCuntcX4Ue5mT3ML
V0WohnhTcYQQVyTbCtxJYi9F6P0yiO14EJcJPFz2o57GusYKNGFcSWpz8LhxB30yWRxEmohSqbGT
fWvp1Zm/wNn1D64mcxrayLVZBM47wotA0XKLGceMkkgk85gqHWwlyKw+Nd56cVof4zobtTR62PUW
MGwkzAxhVfPGreTZ3Y1M/KY0Iee5kBOB4RM9xayffjEjOigv6jpkwmEZ9tgz9+88k9vcmNi0I09R
bfeHf9Mx7MuWR+xoZZMiHvS/AjG5nsoEKQsUs36/D2XrpRPEijYujjp05TUyHLJZ1/9EFFfEwsbx
MZ7VG5UoJkrKqTYUmIzFIitVxoLtApNJZ1awc6wcbV4pgY03OprS5Fv5b70mVMP4Ubsu4XvDpU1q
lq3K25n9OyuH3eDvPHIgICBV8r7NtJONDFlpmGHdbyLc1k+dJimkPR/ZzPsWyNCLFpwAB/srouF8
VHX38SgN+VXuuxHjAdSLyoE+bmaBJNg/OsWebzBE4xTJRr+zFy5czx+z9xm8UZjX9YjPenQ1A0Sf
2xJMjtrx7l0viEhszsfnP8dIWhXvPdGZWoLAYxQEtTPrW/csw/dkLHwAg9BrvKld3IUa+v6gvbof
WMRNUoXfj/1Gb6jDSZEsrEGB4ZZOJnM8KsfIw1ksd/puPzaQJ0LXaImhzDpO9R+cmd7oI7AqGNKY
YdRiHGJ9yZLGe/w278N8t96r9v9T3gycDrjN4KN8nOkpuKl1Tm0V/ARQiXYekDB/giwkHl9cZ4Cw
H0Q/9YXEoQCJcjLFPzEllqhvRGyCwzKs+OMYEhzK9+OEvC3DbUdnkP4PA+GrXMis8ejbqlP14JKh
pEXKTtlylKTdwGkAz5/vSEbZvulnsJ+eJhOy8AcXVTXcUesXPRUMaZBjbgbA3bFptyD/66tJ2wh3
/z/moV4kfw42l5dV+cIUa9hubDDKn54Dnjh4GPurFv3OMMHSQww4Byw72R/Kr2EQy1f3bxMHoZnw
o81P0oJgMUqqQyeR0L8P1de7fhBBB1ftSBfvMKXTETO4cz4/tPRq3eGeq2fExgcoB0gCcOWTj7Xb
KsoYqgHGPd/FICu0pRBPb0JyzQXmqdMEznifQqrxPaf88HX0yl6NNuk20cip0IQfmcu42QVsN6za
pW00awc4EGVmvNvy9cQWBoMpZ1wmIHIKbtwufVX0UmY+z5KuYFovoZVhcxohL/du/eYCnGcVJqYQ
nKljqrOVCi3qIazgBnmIiotPfyb61CdpsC9YJWtbwwwIgBuHXMfNVzx0NV5By5SMZH59JFQfuLsd
YaQZzhOy5XNYrVK5f+z4QgiTz9+BTSfZHpsyHjNuy20d37cFl/UNtgTlYubV02ZKlqyqOtw8asIr
zBhvUnRBsca1Lu+Qz+2kDbMHccPM2f1kDaLP0VA5+58o6GHPcIz1Okz0F97gGf0tXeweezfya6Ge
oXK/PMuT2Tr834JortkkGMMOvsvjgLuT2djxQ1+bxRxMgKnu1rMiOmIv74cEz7q7dk7p2cz8a8W/
S4+AVgtGYMzTvAWihhPnxJj9E4jS2ENlIwEaS7Ot4FbBpcRaqd8CqjjwUcR5lQc0m1HEmYF19/QN
Xq4xh7TOShjmmr4YM2DOCCqC08qgtPfTzNJh81GTeNWKhPGTE0Et4t1wlHgbb7YvMnWhmKKG1vRP
KShz/5tpfu9Gig1quxM0WiJvM/TFC7BjvlyjTUKhAW9SGCWORICBdi8Zz2R1DCe+2nuUsHUWWq2f
il3rJNJsHFQCg+cL9BrXdjaPf5aUlZg2PilaD+OS+T7OaOJPaaz14Q6oFfmd3Qp7xMM08+nbAwGj
KuMB8N5vGhlv9c6GJ33ZDZTomRMWxV4j5XL2VRyr0gNSrGdNbqICl+GM+7lmYOBUW2dQ1WUVRH6z
08xA5T5xgwINU4/g3hqYBeNCMRCKmFTrz+ygzVbix4I4fRDim8QBBYLigXQCuQoOOkfH8Uf5m/J7
j/daw5U4WM5bXva3avop/QmO/ItaXENjCncJ50rhpgthr6UHqiq+m1zntQGYIxPYJJPbul4tqtau
/sFX/80KtCCSoo3MyG1whsk1QOQGumP3jcdIKCt+CJoixCRb2GxCJUn0rkboOB3P+4bQFuMc+i26
9Cx1yties1hxZ0YQINcErJ6uk4HXa8Z3i+zpD/rWBBHl+iOwmAkJz1ReyL8K3ciWlo/XXe3BsV1g
j4NqW9AU4OjBGD85YmbFg/SfvoWXDfYmettRZ44Mp87YD2VAU+9NcV1nkdi752vys8r1zzOgVCLt
PFnC41qeNXwTFNN20sytqVzll4jdr1mwUxReuX+DhjrTAQQGusr897OGvg90Pd+Mre50rmlKb/86
nvugbJ+1/k81r1OAHLcGKDgJkiIIo16rGbTXW5E7r6qeWeltTCj5wehY7vtS88niGevyYpfbRl+c
lTB+FhJctIwihXzatncU9ffztwwOiymbjXNrhJbenO+OGXt6trF7VrojmnEKJGHh9TlKdUt7BQ5f
K2j2vmJhCcz2I9gk9wZIF9Y+N/qof1QU1r+Gys6JF/LJ1k1w5FmnnwCpW3UASrPKoLDN8OplRT0W
rVvp2gg9h3k75eQac/MMkJG9M9Oi+CXOSwo5HZ3LujGEUU6ou9fZEEarR5VUfgJrvy0KupT7aB/G
7sh204tec3pXxfFUlaawiQCGh+gApCNcgCFtahKzSbll0/MeD93uBEM+B9Wqaf5quDm9wM1Kt2DX
ZhS521XWFXSUPXg+pS5DwkUGUGUm8g5VJWgvURoRMtau5Rsm9rA6rLMEYbfbj+e8UlUhbYhr5yJ9
/THQGvToUC6f5jyWDjyazAzjevqHhiXfEB2LUziKE96XPaY04Bj4/8fSFaH0n+V7eFI2/ebmptzM
5r8DanHasHIWle+rtqkXcilnkTqtOkNn0EsCd/l9nkbmZh651RhuQG6CO7b7ibHyaOB5XOLDjKLF
/JvWIK0QmY0rpafqzenTzYFUXBbCaugdf3mCxDZHmm5TRS3PcAPlqraDIwS4tXoZcL+T/1ppqqAg
h+HfyNA78xeLeBgN154BgVswCeThiiDDFzer+mA/TkReo8bDyipe8hFhJefn9YFf4jPoUrn6Fjn1
4zj41FL+Ve4oGykHod8y7rKe5c7plBM8yPQCYH8KuxuSOWYnvH9kIRsgfFZp5rn/ZlBTkInHGHVb
hENY6aN5f5szb2JQ0akUgDFCyulTw5qvPuVcxAs4RaqvZeM6ZjV12uMWn+0DUo1vJ6xpJXs+rU2m
qsj+BgyDwJ2GlxuQZoe/7st9K3YTw5z+klSj9x5GtAybTJ5VO7tpqa/W9Ny74nt/PhCFyeK8w4mV
tiE/15jadpmeIeOSPyY3rlytEn6x2syQQi+WDARIZP7+5qrFlShQS43zgSpBFE8F3PtZw2cm0jGj
7dab9OFUTigc4Pw1zo29kA7JlZwJaUXZYn7WYVFO0/hBVe8RyZBqSwQnrXfJmWjvLb4E6O3nE9S5
lfAAipuXv9euXT5hpZfdMqsnALTAEVFGmdkkyfji8Q/Uvf1kfTe/MWeIwZTJqNwy42GNoHfFyeaZ
+0KrhA70pAXd/YYb+fqO7dNtGjHVSntkzuWCjtuE/lXfS1NTDURr+vcKmCE3F5Fegsuozm4fkqLw
1kvjd8/6hUMoPDjPWo9K4HOcyCdebF2k9x+8Vdc2L865IwpCaQp3UEiCJ58kxGzqNn/l3qtxEYB9
0CAccYNOOfSoiDa1BFMKUBe01Py68YdyVld72i9MxNy8QYDVUPcVG1Kx0jbIgKjM8W9CioBs63Mr
FE+V1mGYFR2+jKf+F+v7Mz0W5higlkuf7tVEGIwAxK7L4+lo3c1cKL50Re51FY2EIloxmwfaeDnm
4JvlvFFMvhSCF8RLhBDdS/v1B1MOfSZ1gh13PMI3x1k03J7MHwRKxXmgwhOI8+WoiuiyVTpe/HPm
tuYvZ8PyODu3yWvDrjeOAeN19Cz+wsEN3AUiw/139aezn8DcAPbPAl9ym7Zi69rLOXm/MOcr6yv4
l+oW5XaeAnCoUElWpVM/KPFgzClqBOyRU0a8OY1xF/NJk4cTiDxGlVlrQgnOj92JQzE5RLsnXTWX
PSRpPz0eXuJKUVPcw5sE1/rHAtx3fwvoNaueJ8Uhh8vg3v1u+pWUMurCXpl5PDqpW0dggnE5bPWl
xbDLg/CV04yROjLDhHUY7Lx+3m0eUnmqWVkau+Y6+TNhqmiAsMKOzsTY3zRC9Ztmi+zDjGHybr82
+Zn15qYgkrDcddSBPzLhRqUHRxwk/z+5cW6dv3HISiuWHSpmnrJXh182W1ElN1HIbtj1wm2rH01A
PkDCbP5DIPchUHZoeCJtFBS7b6KYMGpywIlSAyHpzboBMmflzu4PDkVIZUY1IrXIhSswIAF5Z8tO
M2Zdgeo7KXMC6T0nCYxsmx7xV+3a9JXUW96FXeISpDZNhO+Yw6ZvxrkWDDbx1X/qT8QrmnTQorOb
+KeyR6DzpbaImKj4u/3qeb7SWvElYlCjTO+x2o/C/+BrOWMxdXqaina5i71+AClfM32RWGVca1az
3oZKMazRZLjmXfjFWg68vX0VMqJ1i5BPT04mcH9oRIz2Ei3uZgC6m4sVNOTgZ3pLRDBYOS00CmmS
lH6qAU9IoYHQjjNDmlvyNU78U7MYtwpu8JWPIKcNsJ31UQBdoiXg+F9nDDRxQdbF07lkVyHDevMI
kyo83EvA2gv9SInsgKUkz8D37AS9YfvYDXicxOGOa7xqJ/73BQ5NTOOrcOzb85YpQyK8ATIdk6Or
rgQU0WvEn0J0a7uHlCgcoiw+YtKS2+PvyAoOCpqLcMNMO3EWj8YpS2L78/1DdOIt0W94FBTvAy8k
RDNyofcIMDo1mYLq6Z77tVHok35leJ4NIL+yn7oAbLjjnCfwrAcvxsabS2uwCSqwQNQhpSrVWYYR
HJx94c26zcWCEknRdRnoa0HCy6yJmW762l2tTgc/pcPmj7zUWMUQh9wV9nJBrdm5EA6riw/YZnse
rnhs2nbmBueThQJx17vHqMEW7ODx55CDbb4Y4rxov2Sd4sf8rhhkqropxa2zfXLjpJAbj7/5LRGd
vEe7AtRn0C3YKzeNgBAAcL3jJtEwfUZqOkKjmSUg8lV23wc7GOe59t973MdeRGh9Lub2gDLiKZHo
Y/z89l6kxk605DyoWPswDK5UvhstgSlgRiN10nyNfqu1np9LzRxWy7kmcrx6KU9ATFIIru2LeaSD
2J1E1XKZe55W688omOTec/ooqI3+5cHoKBZmw07aQTtvTFFbxBWT9wtrB7PXivi1Ktdo7LPmJkY4
D5F+ann3YCZ4HzzTowNoTS13YpJc1kTTnlssty/WZd/s34ow0XgR1VP9i3psCmRgZW+QJ7pLqeBk
PUwZIdGQS96YpS1RBhNp3u6Jo3KxykKsKSpflR2F1Ua+aoK2uaa97uXAEOw5hzvC2in6EvdMsSpO
JSW6Bio1X/3FuSw0YekxMJDW37UsVhyHYgJu1LizoVtFQ6BChWbQgnmrSq56uO5pL5ADRxZ+fSvF
7XkvHqY/RPtEq9RYdsZeyzFDZAH7uwmFIFmp/ljGFVD/W3F7eypUs+l+xt9pLNmfolCY6/FVqrZm
/hU5YToUzPhbQGeLu2mQdMXmghtqQX8HpmRH4j/6YNPfw/U6Z2HwNgHtfPKUQsKLiTUIuAWvgszX
LpNZ8I8XzqXVIgMmAtW5XJgpSv0LpSlXwA8e4qwdjNvt+HqgFcieqoYtyrS9l/26v6gxGd5rjm4A
3foIaVueq3M6bHEriPIUXVwrnh8w5m3MiYYqJ7vLEAtBwuS+YJ+gScMRlvWTtKI6CgGq0gWEvKPB
vEwA425lS1dsDCwrqzYGGpeWCpp8fPyPImso6F3xrxvSC4l1a0+LIDRl8deUjXO/eaTBNJnuvUju
jBFmtWtpmraJlBPQ4WXnd8RXDV1B5CHi7G5dBGUrjX8GdjeCuk3I7hRk07K2MfNUqfLoqyiqcAhn
Y2WRIY2Pew8KbMb56wYAaL+0dfQmFF7qKuS1JGtx8TpRPJls2Bb4LZ44NMRjG7i/UPIduNH9WMiz
CdFmjhU654fhUUak7uoLviofYZPN9pKmIV7wwOkOBaMdMTH0P3Fz7b3YayJBeo6eLgQNLoou3Fku
yROCy3X/uEZYM0HTO4M+b8X2xA1j5OUPhoziHSDzicYaUuoEdgSc
`protect end_protected

