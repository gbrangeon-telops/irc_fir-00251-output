

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Qn7IteVsnZ/mdHCLR8tB/KgmTn8ijcYuBtDLGh2oUVKuF3qoFWhv7eC1IOCXLirwb60qousghfg7
0xqsSbRyrA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VgzxfdCZunpPyUwqbYGeC3ulpMsK7w2LNEgFOrFKGlFGTp9v30dyUA7MsiKFgCrzzKT+VrIPwMvw
QxU3GQIE0b38WJ5xx5bDenrFuj9fMfRnJLJFcG2V0iBV/hYdVoEecQkZyqCPVfkUdjfKW2nQQ9vE
YSgHM9qDx8fLqyQ6zAA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1ig4g7vOmzvtScDRtVb+tZEnSyg+feSk/Z8usEB/u9AljT40pDkFhR2JxLDYn3XXgfKo9dhNCFm0
whMJYjKNylxxgSFkNtQwR2XIg0BWg/XJdnzmvhE+MtmxAUvbHjuEhgVFiobIjRufLvFlBirtf174
Rb6IlMY8DFzGP8TNtNYlVuQtzXS4NvjPSDwmxdLLBUryIvh8XgTaS4XKcRx4c9SU8usSs2eZmKp1
PQzsFR6KYhbJsoU+KNdgC0qr7WxKSf9E11HFfNp3O241b9T36xgfVJMNzGcu/ZHXpRemcPttjJFK
GMln0o/DwR0gidlS+JLK6pgrPDgP5/6nmLlP6Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yE7rDdP/qWpLchJqOpJirpc1zOl8T978Yfk6G9kBcFGYD0r+ZC5agvccz99iMwduJEgIxwFmjnzG
7g7dI8mK6Rjj6eLbQ31Mhsmq+p5Y7KQTNM1pfCzFCw+oJzuBbgsBggo35NClB7Hfb8DM7OriNRWJ
U8K86UkzA2Prba4TIBs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BN9F+vWJYtgfrzbWbiAE08ecWOdWyzeeA+i0U6sGshkhExwtl0R/3hfy5ttqQZECat07SJZlP3jh
V4CCuSQw513kvIfiNR1n8KZK1ODiyg59gOwmz19wCVgWfDfnfDXmgYxf+0derYmc4F2n9+pXRhDQ
enznNCCvV1TM+SbAXbMWWC77ZJDkWposT7aeuix0KzNLkoMsiFOvzPJVJxWsxkGPtD/xLXraVjuo
/R9zbJjLpYz0T/O/R4G6FwuMiIZFlEBmhA8YI04Xnb8Of0h/udsHa/BIz80Zs9KgMYw1jOPT6P6u
7aYcNrAi7eu92a51ZSDtMllbDqQBzVGgrUZg9A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15376)
`protect data_block
EpH1xBquEY6WAyr25WgcVYyLjxHjjSo7j/0NeZBx5REAEsd0RsWSIqr6dJmW/Rui5J/NiVame95I
8iw7cK0Dyhq49wKX1cjmbjVcrYNzBq80/68ogyS0qY4FNkyOZ+DLz46x9wHFRtV3ZGc5aWEbJFhY
COL/WA1IOClJrj7W6SCutU+yXYFPCHMktMCYGq40WkTuYcd82/r/p03v0Zq+Cv9dkA9QPMdJARnZ
v7ZGTrF4UWAT75+dp051hw+lWR4h2olxbxH2hEBOGesexqRvxRqhbF5I4Zsu/a6JYuT70lny8TnF
Rk542W4+A81EXl5m9OE6UmDAn422sW6KGpFUMsghcKur5EGIsmOeP1HImZXDHLQgRy4lRAYOmobQ
u/67LPKJF2U9xB3KrgN3lUPyBr0/KuFPuD6K6Yh+/uSEx3IZqTvpMx2FSP+Ev9g+lhURKkesWbNu
c5RQ0iqFPjh/8+7KSLcq+bfaElkeGUmDO7bGOZPmF0peSogZNY83ztX3Lcdgc0R4jT7EK09OptC5
t09UsYi7Tx+s6VSXZQ2oMVbxKD8drnfV8jcfoebCWZGbPbzp5Ef29VYDPyL18YSR7SWo1H5Q7TEi
vzM/hbK95vxZrPlhYyfGTpXkrjdKrjYjBVo0v7J2pJ/2jntLoAMHJ3qXr77Fs7jkySKLpkOYT6bY
NOg9aUXQnuBqOFwB8a0QCtA5QGvKzukTWp6OeoG2xYWp/2cku3Qh8uwxnRZufpKvdvpxPOTIIIxi
AeP5mV8POZmu8WXrCF27WoenX4d74UFNrrjBI+DsaBdrP8KZQslWxefsLpilbUtBBafeoflDSR2E
OjDyXHwhGRVJqkY37nRbf+nMCyfL3LpffCUXfMpnwlyovUmp4S7uF9uPILgmGu7fcDpox8Jl0bLZ
z5lT29aOnqikvd6+5FaxJQe15N3tbphUU2h+nMQgW96itCcHYCzjmTRy+LD34Yla+xFzZQzAYgKj
i6SKFu09TbTWv6cERc5LdDGS/1YGJdT5PXSPHyZSvamQLXH2LjSJO7DdT+hHx2Mt/LLcmym3kFRv
YtZW3ubtLbavYSWayVW7Sw82uPpnth8rFhfbplmSmFPFGHQucJS7Eq2NDO9ibZbjQGZJAcjXV2XG
QsWu/MYhHpGBg3RQO9jVGv7ubjRdDPll3mM3RG//nz6um/7uAXTWiktGlVbLzs5ORxh8jYmwZjHx
cGFlbBdF/S8KPjB+MLxV9GOodDgDLY3c4ih0wNVO7H2SiQg7wZ8jRCp3e0Ja5+5kUDo+9WD8Gr5y
N4FXAKIb+hdGugBPKr5tLU3RO+htygEq9Gy9IjgFj+iB4PECzXMsf4g6qWmuusS20ZcvwIfl4mmn
G+mvjqC4TRbyCJVmsEdN1C2FRxaEwT01MjzNOE38fQgSGrvfRhAtKdF1m193DJEP/Ci+pHXyKhiT
i48xCoIFmlAaglUGEOOlUi2ezwYsrAf1WwHRluRYickeVvzbkgpIyJPU4HDViYo+0FuBSNAO97cz
dxQyGdjj+13VYgbRwQXmJRAyJRQruj3bLtWnTQc3Cg2VLzkkDTY5OUFdv7dO0F4bR5q2WzcsC84X
/Ug11SEvy3PCbjOSdPAP2O8I6OV2nsMaAL0zc5Uavfr+8Nky082fXW/OPNCg7sUL3OBpoMFaax7b
64oInZC8oXtJk+Ok9sdSTzLjNIE1QT/gfodFAAJzfdf+DLBfh1U5CgU8JHoO57zVS+3uoiI8QG1e
Y6o1vBd43+dsftwiMFo4TdYtzVhJgoFdjlI1iK95z+ayyMNrb8MJtNFBKRBWp4ZlTkYYwbit27XR
hIZ5ktSWTS/Hl0mdDTNxLAqUwnz0JRqo+UMlu4MN1RGOI5l3PGBu7Adf6W6/JjjzfeXLtPx54OUn
sqCUO01wT2DDwmvLIxeuRtDvBUwZX5mTAYs14lYMMvo0D+UUi59UkI1SLeiU7aTj8Ds2gXXQes29
qOvWZ+tnAEXwp2L9Ily/NfgjGZD7Kuy41TdwGqdWgAq+zkxOhEcOpdBB3fHRg5KppJ4fT/I7w53p
KOWXZyGPyvMjI2+X5fpye1pC0Z4+wZjZ7UQ+fSwV7QzDGzcfGPouti0YinPtG+NNouVoNLywzxoC
zHWbdtYBOKzPaOzFZ923N7LXNTcXK3gI5UtszUf03VDFNZOFoR1GNorRqEA/fWSpXbZ2iQlKdCLs
drI6tOHKkILlG9VFxhZfkw8hGKWkv2fmzmXTthm5tS1ZTtBtIOLyfkMbvGSXg9EvYtzwI21nMpEd
tkTAx0JoNncwsez4upm1bakFV1LxWb0Zx1eVew6zpEzQdU1XQG/Yye1FhJ6cRBEZCWR6Jkj9qJPK
l0wnyTjdIRT9aJX2wUE+DoZcdJhOpDxfijjj5wz9iMhQewtpvl+F63nnDAE4sMa+Y/sEWjPal6++
XKIrerijOQDydqQ+xQRoXYYrOeoTPN5r43sEepPjN7//tEYqnL1K4aPaCA4DqBLnUacAdIvAGVwY
OYUpjT/bZW1QAhsjxzZSvmWYC0aPp4AOPy/nX1EZNNv3l/Eue/TWimh5QvoniHfoRmw55LNzs6Zv
pgR8ZjIHLEX9QqyQOH0l5D9ioH1QpNajwtporechkHtJ8kKruES89ePvqT3B2nEhPx5xeWKSywqc
HqZILYosj65qA4juGTDgTzhCaG03XI1VbsPQ7xrcDloSMfmBWZsQNQKCdmx8QGlb8nhGaM7Ybu0m
AqMZ/oVr/Wn4QUHHZOlpu9cCJDjuJ+EQo7IsImI9kEg1sNcz+Mh0QE6RpE05wNKX+UMEJVIWgV8m
Cq3Dn5ZCoo9OG1sLq4opavDuxCctx1QnfuPF3L2TXWKWcWfSTkn1d+wB+ycvuSAYjUvBLCbKmaLv
X8YChEkDa2amVXnQEeNyZNniUCsz1Yib2F3ECk75LS436bY4yDRzw0Gs7AcGKXPrZ5u3EEgnfGlc
5EA3auD7OeV4WAe0NWopOt6mPf1FR618L5CuRt7hh5YRZd9ciXr9fjX1Sb22rKWEfSjJCgfV2VtJ
M1KTMnzVZY2auwhGnzpzQUKjECpa+8xYItMpF8iyelQlrsZhssTXsODLa/wg/PXMjjwM5aueDviA
MvLHlAxGjuhUzU7HySqV42kwAjCATS4ntklifwn5b/LAjubJJa7GMdrjXbcqsJfy6Nhq78CBlgFv
NDP2WK03Mv32OwhDKGNoAx5WqjUOurpY1pfA6R5GTvD9xvVuHAa2qvzfdv7W3vu9y4QVqyk8Upn5
1plUwb5+nUwTcFWuIplq2uf2sXgNI080hIsu5YQoyMdYm4GP5WFruoHfotZ7/czGAqMrznHRyE1v
LI/n5lEwonQdAZ+ErGYAeNsCr0PcWVvpT/zmvfsKfaAmGE0ccSMW6QHhh38jlI6M4wAEyPLXY0fX
xqwSslwoANomlkXbshrOPwxaV+2IZ+7Vd1BNQEy0qgBBpu3AC0GSM0ZMOiX1paYRODNfpbA4cYZg
iyCDdObzDEuLiq6xcpZT3MbZBXN08rgS5v5+eZGUNNpCBAi168x23Vgkmh3wYwswrnHF/NqhMXOc
JIE9TwbD9iGigVVqwYyK6aKxVv5Qxfgscp1t8YiDJAbWaMkdl3TVjinwb6I4IFCd4D2x/WHqPHnD
D2r1mraWUImpDnI0kb/7ZFYx/tjLcuyxRO4bYtVwzTXclCrqsgKjrLejEjHRP6Qs5RuvzzrSX0fM
FScNTr+6T9ZeXh3hRAak4Na5im9SU1DrUVsqdrNzGL0VRyhCY2j7LB+GjCEYOtrqMg4CFVH7sQLD
4kPZQ/lFPLjYxocPbxsPyQHuU50cw8PXOH6nJWjZVlLOnPimMSAVYwyukGKFoAB63nAKYUIbO2BE
Qq9Ot+qZkGEFEajfwEvq95WCvr3pTNhwLkCw4JOKu4YLknFMRuoiK7Wx/p/z84pXMwTbXCdqGddb
lqQT5mq1OB/xt/qMZsjPA0mSJZK+7sbjOijD3I8D8oHclQZUIKsNvZCL840Z4ZxIBPVfdmhfTpVj
/q8v5+gF4ZycL1v2+rLi04Cv7/zqw5Qg256XyrS4y0GlAMBpHk1KoFhv3y7O2SlA9JRykkk8ez9j
3jNi18MANDukRd3fwDOvk1W9RDbmjy7lpjlWXUJMdmNOtGBVsCW8TtNecCfEfb4arYpBLCEiPziG
zjNQRrmbxrqBFVqnk0YoLRG7GBU63UUmN+cViJy4HfE9n4mNLOmpXlCbio5fucZSPXOdmzJZRaGx
FFdl3UR0jrM2SNJLIiKA6sFPH8LWa0peopnF5O+cNvm2VPD6bJEpNDQTEZuAs5jbS+7EJ2Ys3MZC
uMIFS8cmihdSdLGOaUrr73OJOpTM2i8XeGXoWfU/I5THdyvfnz0DZ6Lk3XGzG3VbR3OUt4DJOlbf
mHvFXTVQcqc872jsFI+5kWyGS1tHUilPm0U1t5m9ZUTsToAYUgrFvjdoGOuw6O1+0Th4KjuehuM4
a70XwglFz5wbVukjWbnX2XxsEib5oozMNP/kRF4LAav0zDouyNavzYPan9Z9epWIGY+qTwqBeKbf
jkXI6QG+2Ks1PumlEFGSr9EbM5z6i39/zW3X6cA/hQGBLQcp12BDEaeysQVXoyMtfKbnUwf51ADg
XNARYtKzFOIrPPqNh9OYUM0gE7wFooRZilrKbdeANsT3zpuBcAn5CryBJVd+DPf9kH7po4olMrZn
BRb3peV29Is2kYQTtpgN/y0uAcwZlEwEneIGjzhaJ4O6wnzQ+t3dcF9LCum9/TS0OnhdK3rTDzBa
JUtzRSX9Mmt0XtuBfU6oEkFvgYoUI9PEKfd8nsqiruuq3symi56sg7YsdZ9GJFW2ACfHevUla9VH
H78IX8mXPqdnZKcv6Dt8Uv7CP6FgNawbzQbqz8XOoVQQVl/jjLEZNt0vskSjBP9wL+jsSWki/iij
k7CJAzGTD3Zik1sQaMGEGQwHtuSeYnJv4p/XtZmZAtRZJzVRM56po5ZHcy2+lAIjdN7YFJxHT3Nr
dA2/mD5xRBTZeih6lJGve5dzDNttGzlg0TKyLStO1ypUtP1cw1/fE7JVmdx0+XgJBFbnYudznEt8
GtlR2ETpXTmxWEz08dljmLWi9oYHihU+hTH3z9rpHl2uB6FC3pJYMej30kcxkGRAjEiNd/Y3gp8M
kUpQyXC+AZetjJDEiFY1pk0PgqPb3lAhn2Ft9uZLoIC4WdhaG70wgpwNVeokCkfLsyZsmzbnmPaX
PRkCb0GvJUKVlRFgkVKrM38HYmVibdnz6mEPWGI6U/ojdBIxw5Ln9lGBuAK1xOnXrjZxKqx+OS1m
nX3E5z6UtasQ/VQM1ebvoU6UJqvxk0blMl31AFMWYv3RIubjWLDIq3IJNlCyywOpRjzPYpzBQs60
AM0ydh8/inErRGrfO5Z7LC7asoUlAMdzzF1tfYqUnrhfUYSMWKTzS/m2fajP0jKLGmJgfWyMUonS
6jAba70+esCItFmuPod3bOO4q+S/nZPyinNzncSdvwqwTgsXVmBrytEo7E2QMXjIpb9KKg0tB5vV
xQI+Mi8PNyCJ+u/gwEl9rW82bJw//X7nRFz8+lupqBaXeK1sQt6OKLZQJoHkf/GbskGpE38tH6D6
tCr2WpxbwuvtJ1m7R9r8Oqk7BivIe3RiY5ebfKovlDODfHWlEIkvfA7OPBgl4MHtRk7lqZsJltX5
q9LmWorqGYRhCFpvN3G6fX+o5Vtv64Jd7bK8WG7/ycw1A3aD5AOTXBBi/yOrdzG/sW05giWFPiB+
JOm5gTVfrw+4p77vd4BJOM/73HuQC/SCDi1xUseqcQVVgTe6P4OPIQlK8FdFw0apaSpy6i9ikLYj
6/O9+sNGGaoyG5ak7HOUZKOzmtodlfFwMcVUpQfL0eCI7nIUUrnsXcEDtWf1sCkX3BXtrGpJoSX6
dg9CRxWVITdKKQBFvZvEssWk4FPZoD2GqtYUE7iYWPKkxF2MkfJtoiMqtQh9n55UcSlnEfSeoMvZ
91UmdeR3+poJ5+bFH0vawYrKIJhJWIHcAFjsN2/pzGbdC+jykyjVk6SoidT7H/1oTPSuaKgqdKAr
2DvlnKqohS+MB1yryeg/uplsIQmYeT6nBvcwodOKQbYT6KVnmqInr3mwFAUWIC2WrT4YWFMqzM1x
+9dR2agPidkR1RBf1svYGxpwhNNltb5pHZbqYAtLKrnbzhqDV+GT65zTBlq7Zw9C9hlhUhIvvEkQ
x9z1HcqCKM7NgIDFEoBrbQ7+R3X7XnQcyLZQUk9QhYaZgV7gnQBT5x8IP5MvmrhatQ3WrE/HbA1k
TKBjrnI5iou3VEx1iWn+kgqn9NVawFhzB5an+R4MgHX46587ea125dXusocpO2iO8Mz+QcPVA4ah
SKF8DlqPvMGMO4O04dB2pSg8MEpPUxlbDUoz5rCDlMGDGBoiOiQz8mz9O9+Sd1wCFMqoHyuNteFE
3s1PnbPGJWBMbsv4hnaS6j9Z0GpoxbjjHjiB6ri/Zmno8DUXYzPHuNB3r3QII4QD0MF+hgp1YicF
8bOMKrwspLWyGT7fPp0ZZUlrisgSOxKYVmheTNJep4D2siFDyXN4w48N7WcKCj3cyW4cDQ2da1dz
E8WKiLeh/aWgQaKQ5BHyzwfQKQEYvfISHZ+rT9ufjMJLaoyt7t0P7IK3hed1bNKWqd+SZ4E3J6t2
Iv4ed0Gtc5P4E3jG7Oa3c0WVDkl0Fh62W7R1DMYrHsZqfg8MMzW/xDPPuVNnuDlHJaVAKd6EsTbw
JKq2iSAVvtnZ0WZi+6eOuLBOUtd8pBMV95HvS49Z1u9qiTitrAvrC8LQzUAfStLcEaapQXufoZhf
AbzW8HjVRaTny/bbSHAp2Su03cqZYHDt6MkTNB9HZeGuXx2Vmj7YYR4mOii9nbuD8DrMNsksW2dI
bz3QaLDCDC1tz4B6A8ptmNjAO6X0HwBz2rBWCOpZKqKO2TPSpuUW6PFhlx6sikQn2eHSfftx6H1A
NtV7FB9pGDbqoTsKjaqYsUOXfmij/Bfr0yHhE8ABVpVd32NMcx4OwK26tOiU90meyzNFHcoDcoUr
X7VzXGMcWvL8fJH5OXUTKMO3mC4N+RGbo98NFfEOKIDvrvuM470P5O3TmIoiTnFj5tjfnRMS0ghw
aiqyaSCnemhYBkB0GRwm1sxFGeBtOGBgaQewYJ4fjXD7fr6Fn1znDrA212+cunUggWgwhc3gVmbH
ZbQqdbbRBtrIHZGjMjH9++5vff/1mpMTnP2SoqoYQ+Jf11zFyB9Gv9Bw4SACOfb32xusHhROsGfN
Dv1le36PvgppOfDeEVVlRtROqc683nv79Gs1eYFF86zUdLkLf484nZ2yU+QxrmkQGsI5OKGpeckC
EQkp7pTBQvq0NN1/cx07mXoG6v7H6CEDK/J249qeYw8o0e5RLulRhVjgAEOgehcGh6MOK+g05Zng
SuGlE+g9caMHxECXK/DOrFmz/aGT837usqJIFO4L2NDStXJpR6B84Iux/7uFU55cSS0lhb/Vh1Wh
AaYJeY0TdwiweBephnsHDrizeJGSBKMbujH9v2sy3UkQmJb9wGyBAvtYW0YyAKzSx/lLB1QlXhxJ
6oYPMvcoEONuuvQyfj9kR3wXAX3PSbjvA4O1vFThDZBNlXMAr4P6QcR4JvsccjK7vdY4Zymcxv50
RBqjwwd20Wm0c5OOrxZatQ0EQLbl00lsLNd6g5ocLhsTU6XuRIlsIKkxP8v8Tu+0Z/aN8uodMBtP
SO6AwgNxEI98REaQSxzfEXMSRhOvlx1CenkhJtNoof83x48KrL4ILh9ULrCWWLY8G1sdjmqzdXX7
YmfcSieo7e0MTwNtwdeT1esNhjSuMxhibWwI82ftD6oMzHokgqCKy8O6EEfNZFLGmVg+LpYnme4k
alMFVdue4hPJJeIpnwaEfS02bpD3iUUa58/bzxvIoDVOQfoRNL59Zd9uw1zocnIPfdCSCKvWUWXM
76FgvXkBYUpKazWlUpAhiEWxtu3BI8Eg9iDB2nnhcsk9Trd9eCVIRZjf3GkQW+rMxTFbZzwCdbr5
6z+xSwsmtvFQv4IZPcTIJI+8j9TcOFypnI1TCDmkdlTl+O/1hkB0/tqWhQUoEGiYyOP2i4804PWi
GetQ8PW3FUZ8ANguL4gmTw4AXe2E2Q1YSte4apyOvjZ78w2nPuRBrgevsLPWEaV2bgf5Q5/3cVvh
H8NlvYf7ZLbAbkyKtmkoUezgEPR8oJICnJnlCrZ/NNvJVul2nEfK1Y5faiNvDvqaJ8D7+CVIPzp2
R3rr+kyGK32uzDXUGZ2y/y/+qbfaT5hkl2CXYltvP7wHUd78KEiqfQhlmaJFS603d8BSmV92nmNb
B1cShoH0fNe1gRxPzrEl4uxgqoO0vJ8j/g3z+T+vl96vKjeOCzBrCuDT3eBUbpVgSZEWcQeziXuu
WUQdqPO82DxHzWqWiXtMFwY4jlSG1CHROwLDxliHdwrIcY/5Y8wfr8OltUXLzj4ZIhnl8jBz61dL
FvAVSQob1hJqb8mgErk2qKMSoexIaOE69RPirxm3Ayq2BrtAQ1Xjk5bfbW0LhVHYhsLAMHS5TUiC
Zhug+bHYzVzFYrt3aRTiQkz0ftmd0xM5mcRRZRrvWPHazWrkUsb44WvxfFQO/kSqICVyQ5swJDS0
O+uyT8kXipOczRe5oyHGNDB03JwwNkEyD+7vLH9//KvvT2hULqUwZxZJgJKc9uNPl4jBet8Hi/3a
KZ8QGTRl8GQ1zQm1r924W/phZLcGgk5BuYURb4YHvAmyYNt3qHwyi2JzAO6fP50YvJwHrkYY6Qor
FtNtH+IH16ZR+AAZsF5cV/uVkZpCjZpw67qW0r8rVUDwvhGw5QjAH2FxcpLJeCZVsPJBlxl1Sip1
JkORBPIwGd1zuboD0X4SiHp9HOJxDfz3cNd9C6mF3qDBAd8H1SjR2sO5CeBax1NER1pSMbz9UTMA
eoPZV7NHTjrG3Wee2ij0p2QWrOB6Gz+RExfxXQ0/sDcGCYQJWM6AwF7oo7dSZGn93+LF1CiD1cRh
tB2nGYr1krCIwOSYxR2eGoGS/xTeBINgQ4mGxy4GM5JqZPe/i4rJ/ykTuyijvpBUQpvb187SUJ8/
sbCHCix4t52NRLD4X9vI6lnCSkR+qmSLEE6/I0ElWpgdJPBOW4sphoc5EU9mx0lE1pwYeDBDq5Ie
4AoPwB0gl611KXTJ0Lv/JP29oWwu18oAbDBowyEk+3Gcza/z0W5w05IoEuqS7pb6jHphqf/xlfZ/
rUJWc2eXX4BgyGPwvF62mrxwRcan6aFwUyHqbgMGWS2S51iYnKVyY8vSIL9WmdyDFTjs/sEwwFyn
/yQagGp4GXJsdrYuiSMUIqFbnz+fchYXaWjvM72s4HgxFvedeCs+BnBLaf8dRmcdwg4hhRy+smgg
AbCM6S5LKUxwQnVWMQ8ERgMK9pdpaQjdRnIzt3CYh7WQqDKUt3CpL7gqqwygB/mlrjVT6b7zeSMj
rv6eOR50DWzpeqT13Yc8f+9J9CVxi5HECuvog+kz14loTffYVtxTEHKIFUL2QJUz438OOIH9G6Kz
e2tm5DEflfjdTDLFkZNNCn/ZX2MjoqZGhqxhUl0RCwjenejNCz/UiYkcAN2MZqaxs68sDpJSJSvG
+9T4awFwGao6TRUS4LZol4nWtTuR7X58j2kwPO5rbqwDkU9+Xuj5mtEM1eGU/4HR/gMaLAzRFjr/
YXO+V/ZIvLUiOjmM+/KakH1j8eMmIKS7c/227ihYZJF7vqqPRrs0EJYk3iY2BToZ8nfRwvILA2YG
OWZ4tTKA3wJfUpeoNzrzhj/uN6ONvOFrNce8ZGGNTo1mLpjrZ5N890SviDEOGBUgEv/AjEGZRmAR
6uSGgdkj8PwwLwFm7fZAupBmJktLDijkQPPmG1SQe+xMLkobcqJe7DUworVZDSr/Enerp2FYRs9+
oVQhchshe4AjWbzpKfLwpe3d3eoTVvnMsLus3+UnI56Xw73emWqsz7jQ6V0UESHpDFYdyuCOVPnL
H3tp+5xfKANaZvqSjmVhFNW9PFX1iHkm/RmdDbKtBlOLuynmMFE0tgwP1Z/WdVnO7mUtnxB/dniy
OR9XXX/UoCzKjHJP3mhN8s5QKsS/LZG5whjZhnyKsNsOWMF2w0QAwWZbvTfQOfCsiZuvPmiwAOS6
cMCv9/ZagkDGv9nLEav+5G0Kr9DsoPky+4ekS4bjlnXVTxNOADoLhUQdK/xxFPkhd0yo8eDzbcYe
WdN3XLEew4/764YfpkMT0hLKkwmkjzFEnEy/U9YnCmPOSKBPeyn/p7sKhV8K8DBGGxiDPXLTUo2j
LPq7rMwye9y3jfeDGRbXFYrzckKCmZNBD7Rgt1eGJ2GqBknKAuIWuFtJ+pbzVc1/jszXycIwlSEI
HPcI4lfUPtzJa7FWLgzyKiuyeOp3OiP12dnmtWhlW3nxbGYPy3buJWEXD9Cyjacr//RCPC4MkN84
RAnj74+8TWi/o2ds5o/SL7y6e7UToY30VrFyV1vzKkYh8EDE8gVc3CBVowW1CbydDM65U9l3PYmE
0Q5wIbBYFtFgm71wiqry+d6bLQarHN49LSSuou64ODRyE7RKOuVatXoG/HRKeohdEc1sZM0i/xTl
LHVeyyJxZ5hrMqRob3Os+2CbBn+ARlmjOpJsFIjjP6bD173Y2PbCCRUs5HpOZYsCaxzs9cm7PydE
1gHo2UqZSBiSUSV+C12ngp4Zs0vg+ZX+/aYRfV5beTfVJ6T6+BLt7Nl9wBZ7uBP1m33AFLc34zAC
UTmjuFOhJGrGMRDI3mFXd64q4aV1uEdsJ4/o90XdsP3MvlINAnRgKtnV26UkZ9J9maokYEYHBzFs
joBc0uZ88YJAtnFDiSTjkqSdUL957oZUh2pvVrXlRZe8kPVdzgyZ7BAuBfdj7Dz3ciVQif3Mf/fc
DoxyRHi3KAS0Nw+TsrcA69kBqNQl7BexpqhqjDLdak4ZUeL4ZVQxL8E3IgDCQId/znjNLYL+XX+p
6S31rs6S9NbyVU1XiAZLTDd7hpmOxyoqhkwtoSlS88UX6TlG3hvf6XCnZTtbpsBxydwh3bFalWbM
utM9ANMWIs92NwWO/cyAncWtqujqg+MTYnProMHOOgNm3J7HY4j6nDrgzDuBSmqwpzN9OtCyprPs
uJZqxAR4aG0+lq0BD7k6xvQQHSFnxd0Q/mWQYs55V/xVe3WICSqTGi59+Kv9BXu/OHH+wmgl7Lt/
lTalejfgNkKHGjkxBSSzly/RYSGoUTI8lA7afQjs/RgnjtzyemO9fe0tVN7tLDamcz4JVwLLef4s
B9Bu9kqRb3YJngeuhquxGWnfJFUczxt6cHoYpvrhDcPJ8ibkgn6xiekbzsAiUsgoi5emp0nCr8U+
jsBePQjOzs0XtjKN0E5omInox93LT+575ysHKBsWyLdWHMhSOOshDnNJpq+86+xU9KpybdgWOo5B
k7Niayi18+oAd8MWk7a6jGUnt1TlYa3pAvbKASZXLJbNuEGqun9ErVGgK8Mm7oZySEwo5KyBd8Oy
Ad4jXWq5GpKbL9ZBGFIdCNPYFJ2VwvU8WY88IZUG20KYo7m9Pq0UigD+GUz/8m+s76gi/+eudckP
IfqDyZW0Nc4aikiOyPqw0LBnQjuGh/K1I2DIdcyVHZZZ0X+3K6dP/hZar88KSDUpr2sPYqQgR8bb
TV/FDn3vIk8MF+B9zvFe5qHzDPf3xTBeyCGLIjVs6TuWC2m6A1/ZYt04hn67qB3b2Pko1lUMaZko
O9x1duNqRKa1RVQu+ifWVKIBO8hOun1mM/NmkCTzcu738Pdh+d42/90se/sxAo7iwVCB+2sZU+d1
d5JHxZxqXyAbRvW6M6KbA2Mgctiwi+hnzedADkCJNc6aBcXAhpPEVkHnvgg5ld+JowNyKX0mS25q
L39l4MDDvcG09CeDgxUG8QoAhUaZnyeLhXGEZOA+WKbc14Rv7GkDB88/EqwdHRmjGIUBCkSSeCP5
wPhO7a8zV0PF97cx184LsaHt0iEqwp3CncgR8fVwgIi1Wc0QKtAk70PRxvPaGLbKgRMwu/5UGFSh
2MvKyxGVJZKN53aa/mie8p2H5893qD2FGWHiGM+N+fV/WBVszU9Hu0wgDBVcfVgX8DZ/JVGBzAJC
h8RzmPBey5BVwi7dVaQXdD6nrJfHtNbQqx1pbnZgPeNSNeuLzSckS2HKivR7aj4b8JK21i1LXoZM
xsxHsq3U1Rut5IvJ1PCYdxJqLyDzIBWW4IwWkioP3aF4/TDv3f2jea91XsCXZlC0LCovR5nIGRr9
6RVdmjdIRBLe0eG4mm3bvfAzPfuEceN531nNU/TYq3OH3kfrefkexmSN3NGms9SX4TCUhGbIBJuu
qRfPjlI0HXqiKNhr9/DdTIzv2BjvKdpnJuwhD7vef9zztN8/YSDX5pKacqb/yWVdh5O9soSlIauG
wpvOMnTaSJCuajPsu7yAIUvNBjmnK6FJWaxawEDkg72zJsRyZLSImtVlMGxQQVyhByB01mM8EWoE
ijC6G4nJdJefkvEvLMnJaMF8SSBoxcg0t7LPIT98CyS5Ljpk33azGi/xH2IWl+E2aNPie1xuboKn
IPKOGeZ2tpP9kw/o6cqXTgeY0pqQ1tJcJOu/2suzEF7OeUGJdZ7RTSC66yjMKt4nTGnQhwXa5XoJ
MqX1g2uslh+EoZSLAWty5LfAo3TY14iBQ2rRAUtQg8hGU1UMa+KNe9WEJI+m5/pv7k4AVLU9lNoK
tueQjjdSW1+vZMD3JIAcDwsKf1zJRdFJKAI7f6h3PjQvztb8qIg668bmna6cyqEcra1d6wjGaxsx
t2XHDqJuqNgt3mRbwEiCCiYwy9Olz+2bdWYcF8y9I95qjl39YBFza3TV/uTefi21Q/AqQn737mOF
KrvW1vQ8sloXdrK6zB6Xwd/wwI0JZ/E3NCfQSthyvCFgBgpYJcLgQRlVLBXzFGzsolOPiEQYx2wj
YpcAovEbkHXAQ5Xi9u3HRly50E91z5SMLPJzmq6sQAXStgBPgdK3s31Yv/dwjLx9xnIulKxEAF1D
Z/JRV9Oe92553CRXws3O334IaX35LFpH5iFQKHeuDYUTAbR6K1JQKoCOVnDhmI6+mONZPfxM4K2K
1xzSud+jQebHcHoNJviP85Y5fYO2/XDDbYM5nBpSdXPPtOY/8ZhWYyP+bZqdgaQJ49y6SVk6EQca
Gyx+y5wvnAIxSu8vNNaqLQlW8qooyq1dYLzm9DQO93BbAjIoGAGkaIkicI3W83Gk03g0tJCV3ezv
uCtI5PrZgagceEXf04HTPVy5UbqKi4UCGDMKT/6SrXCN2UBVoFg54s5Sk1qqOTc2R0PlNvkQkG26
C2+FLk5kx94+E4zwGuWyTcT/BiyOZMNNWMBhBIZrSW8EoFSWP9i4GM9mzs/oOrDRWe+i80GjR38o
kooxniVYbkUKo0ljU4e3j+fKt/sP0zYGQs0PT4U/+7irFB8zNQiggH5yw/vTqgmFLfZo80XgOoWz
TL2Nf36Dlo7u15hsEPzISS+Rulnn0Dqz4KV/PSkt9rQ7goJcJk/wtxDdEImC+p7uckBLpyssxFSP
quY6YilOdiP2YcDfoyfg2d5J9nVH7JtU5bS+xBazaViDZPFHS3DTC7/h4txUPCRs8ZJ/0s/5wj09
FbfGzRaeXrfSeYbkzEAuI80R5CDFJ+nXGZf/VPIyOmEzp/UP54uZJvQb0Ed1It84dDjVHZZZtnmU
rQvRact8+2LzeL7ZMkc2Lb44QyF+ATbDlTksNnSwqg8VKpfZCUURGXC+w4VsXIdW1T0pO6GeCg2A
Z5AzfC5VPsd5edI4K46Gu7bWVeN0IgQM7sr5F9B1JRx/8htDs6nKxTF0W/BmILtc11o4NdklxfHm
87CoJcIJ40rXMaT2Phx4OInVYJkY3EuUkZeJ+vf5UG6s0yi0wnUk/jVNiH2EjFhtakM8hrQGLExi
SRsEfT5HJMKQBdIRfnYZ1qWe+J/E+giOnroBGP0dV1hhHV4MHt43z2TmBby5G7Q5iobw1GnHPphp
8TI+pTY/aKQUBfOiw6RYEqRbr/6gT1fgI/LJr2bSEbw7ERbvSwiPS1xscIh5McGsnk/dgrTDi5Km
H+dTvB0HpG79lUycLjpFyAWUCM1UhZ4Or2TgwYpirPt5qsiUgSPQOmVZFAXH+V0MhDS28E2INVsV
u1uDYSxbvKxH1oUCD+5CaTIKxdZQ8djsrZz0AzJX4tX+xHPb2nqsntJAQYoCJLeR2MW984RR6jZ7
orP6JR0jtk2bepJU9afZ/shrs3u6q2/GXQdVR9UGCKnQsjmrf47gqZz0j0uhIo/xqYFESpIQAvBL
IgQyMvrzu2wh5nX1mUf9e5Y9iKvcs4+r+DoGvWYTJfa+/YGSurlUeLxax/+shuhObq9HdlC+KGi3
pqvh3zCW4/xxfYuPis6ExSVya+Hk8dSGmB52BOWLUOKc9i1FCMP5RkE6fJfOboGaCxKlq+1UiRmz
oB7TyoDqy4cnUCYlWBwtt8yaM2yEgph2/DjtVZ5OcYy5mM+kcR6x9feft0T3TKKP+iha0dRsgRqG
2KEyP2Q/C/SOy3gvNuE8AdIDIiL54HyTMjmgwkObNiju102YeZ+wabdAdKPCP1nhpYN+NTdDoP5V
jYiJ7DQof3SnaOIHUMoD1zKZ/MuR1tBfGYYVl4aOGmB6cTqk2gnBX7SkCrkKIuz8Z6rif29t9pr5
Y38j++kNgGMHxzeG6RA8lKcI/fEEG02lfCmuTE9l97Qt5gIPg0YRSgagul2H0HOiON8LFUAdLh51
Mw6Nk0Vq0Ze+VyLoHlaOz2rnE5UodRAr38Fb8f5PXEla9i10f7U+RhIBsJyO0y8m5bVjy7slcbVo
KHuDXiiEfKoMm9xJBKR2xGXwoGnEP8795xaFq2IPEC6YtFPXyrbds7N2F+iN8UWG/g2uF62btKII
dYsCTNcoD+3nbAitXSXyMwQjUnsJu5pYlBpAx+7I/xPM/L2RcBlKVTDlmt8sbxEe11//gQcZYNft
aKgTcCHafBltf7v5n6lzAq6urknoTDHXI8qYXfqPXkUy2BYqoU6EQiHj7W0hOq79Ex32RIZNkThS
pfLbn+i4Qj9Bhda05BVB0WtvZdmqpRnfOQGXeKr7VN/PKe6Z8uUrdnE+l+Q3He6RcnjO9cQeb+E5
rt9oLQ/bo7xTLK90r4R6Tq1i9j5cyYkjLoufz9nx24QCBO6NHDiTAa3aKpbVKnG7Yy4jyqyZA/Gq
Pzv+XlOn6wG+oLAqWZdmqLTc8VGNrFrbOIsTf2Ce7NXF/W30ygrHWogjRYbTi5OCz0r9fbE4xCiN
DlWPhOIdmhM5PM6FP5bc2RUQdF8gnJPj1gVBJb8wFVUUupgYsyh9fTtdGZTpYWqY4abA5h5hALy9
NjrGgwQXyWSvnRRBdqVYYOuaQTB5Dqz/cPM3S2S/ZdvoNvSwiwOcm5KvyA3upDITQsZdplINHFgP
Cjqdv1yCAKXNsaG8bKkQmuyrdcjuiOxrjgQV7375K9sOg3Eoqu6Y0HICl1JrgJSLbe3U9HhtYPgE
Lpslxlb3mZsofsvjXGSPe+i0P0C3XEhE9dteCwH679lbfbxrEs3pP4r+cqRdKss5Zvd2y3jGqTJY
MW/EMQTA8VrT2bwlKFgXVkRBywIXgcw4xTEq6V3OsTmcaaMgAG7z0GpF+r3cLW3+FxyOz4TlVHSE
/EO2gODirvPFnFrLdcork0Y03BISyItYkJ++rmpnjmWGq+ISTRG3YV1d/tFM2iq2O/ZkN6GBCm2r
Xzl/n9DfXLxBIb4O7+jDIA7dpeppEXwgv6T8HwDh3t6IjMwD/xAN6mCvlvzBS4X3faQYzpJOxNoG
2PfLWoOrgr4vS7a9aJNpbsCt6He5bAi9Sjmo7MiGafSOVj0zNHdndRhUwYKQwcwnyk1PCekOKpJ2
LbueGGQnfArtHIAWvLDfcHQF0qWEPemCf19IAPvDfpiP+X8MpgENKkK1/P1TViKxwGoOBeLBa8Ho
YwgdZD2Z70ojl7ExNSDjh+aP/qgUXS5DJ1k6pFw359O0AJXi2rOuvZQv7FYxoGEwzxs65glRoxuA
OqLTwSPVJnUIVXJqq5u91notTu0fpER1jnDE6UOL+9p/KaO8muX8mexVhJMJyVHzbzLTJYIDZ7Ji
WxysmB8R6hLksAvSkpoIf7hNY0XL2RfXiarSlaRPR/65W3jN7RI2H6UXO8oYc9RzUNeKiIWLHker
OsVFuHWYfvQN2sY/6S+YdD4h5Gu1RhnJSKJTVoNvRmmk/4W8dycQId/dnaA5/1Pimz3B8/nTVmIb
VsDyWG7QwMY0bTvYR1OGouB1iU4FqCQ9Qy94Y2D/o9ZCOxEayi7yBs9Q5HN7RtuGfuKKLV3YXdkU
LdcvHtvekoD+PVkRbgrMjq1jUxSPEJ7opfS2vBWAlHzlaAeLTBNYu7lNIJ9UkhpizQfKVzf9TjgA
YXYysGtzVR69GJVVOpkdxcblZPCo4ONkl+DbomayUp09W0tHCi/frCH4zMeQsMy292/iNJPdjvLT
J1v15wEbxHaHGVgx283qakPM18tI67q6WiLraVMfPDEhd/IQ4mo/qTH6GzGr5l2QkHt60WFGad/r
pvwj8oLRPs4IEA97nEnwMh8ZBsTfcjBf9DoF/iFYdfib4qDdLghoEfsVp9FYKhVb0SXXI22L8bE4
z7fvOtywyU6+8gFoNXOZQ2uNnBISCWlwFQ3r60kGoGO+dJEhH2tCojQJgct743zlC5ZZijqx5bp1
X95mrAbKhgPYQgXmw5phPfGOP4szUiBGTfAVKJNuuGI8cK8rqn4oF+9+mrtIsCxJUsz0XncbWJJb
4WLAsM6IqPxIyJr62BR2q/r5MWxvCEPU5sZnohD8w1i87Vnq5ZVLaL+8LaAAeGsMCtZMWIIgbFI8
ECPHuryfd1i0LdOu0YngxJe+0gIi3Ud69CNkn4rDlBt6wQLQsTjVzN68sUjiK6mb6oboY1CKHC7p
/S+hnfmQ7Ka+rWcTQX17z1s9FCYd46HLQWrSo2CNV/STrzrmBsSy76/aDtSxJgF0Kr0q8NLiWqdx
YK3rMAYAuqHtt5AJYZ5nZUVBSS6QU2MeilZLW3JrYdTzO8EBjgBeHJ/MYrzzXF3b9i8/0J0ImAgy
hhk3JZaaeZS7lvBpmSDgHk2rPFfATd4ppLJaGHpXiN+R8ZLzS5ZGFhjycyWziiq8lt+KF12wlQI7
4pzM/bw5uOkfvUfc3QyxTeU9u5U0XKi5qHUb/wGJ4bvfakZGJqZl+n2IwaOsODPww3irr3O/Avqh
eCbInGJ09E125AcFT27C1OLXSput5yHAUJOabbNZw979bU+zPo3zfhj11tSjK50FL74QBaxcdBwA
IT0QqOkFFNUvU0ahb07abd02wwehLgbNsmuJ3QITZrg/VYqiJ7n3gRY2jRCF6v6SCQcSuJHerSfa
mbZAwL/EGQZ2WeYZID+IgB5aHNtpC+LydyQeqgqxkeAOQbVxCJP/VfYJ5Pj5ibWlIq8XszdsO/Yr
/vYRlDkM9HfX63sFDOriLPJTQJnw0EXRrvhAEk7M6M39t9N8Jth7j5/fOw2XDHu9j6aYWs+PVv01
3VlgWa/AW0zGbvgznxIdapYS9yNRjKKiL/Ww9oiJyIGBCvB8uRxpaFhyFefmZi6Mnxqngr0a+M7a
o0dBbQleedjcTQ+5/5TwYRGhL0NPf9+kt9p5d91qayt0ICrzE/OvSRXqcVOwvbFYWF5IJlGLIcNC
KVFHTg9Cj3h7sub1OfTwzNAf1F9R4sjV7iSgWbBYfO4rsY6lzf1JsxTBLCgLyefDY7pfADN4ybR5
5lx/i6Nyct6HvHAqKn92pocGMlmDWM+jblmSHx92SJzT02/GWnt327T6o7fGUKWOPkAuq5WGFO48
V2l+JMPPXAxppn6TagCwStcEsMdUnPuyg518WuTLZkJ0HQshIUI5nhi33WXfWhCsoMM1SnIITjH7
Zllc40pEtoHvVocemmfmJ6zBZQaBTwj8AXNBMDN/21+zvI8Bj3qLZo2R1RgtGGvS+Sk0HAQZPo7h
IE3GQNqkKVZeLy46PKkpgPccuH5sx0ez94b8f/Sa62m1DcpGS0hu5E1bz1nepGYV/fnrA3MZSiJR
oaekkaqJWOPhPizhR9QsngmESRbLav+1Xu2RD2zfDuke++TSJu0DMj0kT+6ujofmQs6KWVbiIrli
h+T9v2Kor2rtfqrO9ukL9xTb1RXd0TY+8+jz8pO8ovHxU3Stk4QaHbW6xcvUxTUd+l3EsyvlodIz
Rtl0wpyqnzp3tnt50wjVDBiZE2SG3Ja2Ybw4cDt4Fd6CNxVPdtH7PrmxtbfQiwxxBGfJ9MEEq2RG
mvFtgleJqmky4GCbvzm4cU57UXhXtzJbVmqaVPEH93O93v1f3XY0ZgD63YeEHGIGx00ufG4nzF++
Ew7quSImEDBo9qjC3Abo6TA4pcxFgum4U/zCXcVbZOY50+m42t3EO+UXk8gseYrQVL7oRN82/Er2
7QMcGMkQkf5vUqOmwHj8SWJPGWlG0VhhFjugn0booh6fYpK6YmPQAXRKUTiIuLCTbyqIv5pNHcCJ
APU/EvJj/WyRBTF20NzO1paXewq4mP2Z+XKWlXkCc37huiWUrBeALypkLSwZTLbLBH9gfFF7kYvS
2L3UqVsy4cPwABQPNKtWKG5Wrl2DZk+PvYc8l8si1yKjroIKNvvRlQOiGgEfvRANNGJFsDcBGTtW
oCOe4tJkAfXYll2y/rBB6qFCWJ2J9k2RFsta/LblFMIQz1bc9lPxFnZ0aQQLJmQScOZ9ywgJ9a76
27Ac6zqtwqo0Q+vxou4mwJRzJzMLQw14eDzHD5sqMKHxTtZHy4AfTPor+M7uxdJznEIYOK4/omC3
uwYX1/diejkADo3sliCBpfUtbrVN29a9mhlxaOxbvICcTM80mJyETLYKBLHfE0huo8Cye+c4XQsR
4ktzPQBnUpp6yJI33vU/UDyRWdSYZ0ssVxPB1oLvpL5xr1xsS/lxx6ZbJUL+NC7dNLWveLAy19Jj
mPpfOujH/Pt6/Hmo1WkRPnzAJC71FV97Yd0cNvBm3/oAFFjCopEup0QFiex/LnigB5zXFAI7qNCs
lQoa6grj1r838dBpzKahAhJrAix2X1UXsTY0LIAWFBHMae7hJEWTsN5OchAbu2NdfDcIUU4ev/qH
GodPdoXs5qB9qfE/OKii4DAZKTOFfjXXP2PR5FmqGHegMSFSBLldpV7b4Pkrn3C5zCUQ234dGP9h
vpSYL5yoe2wIA+LhWP1W8j1w9oKp8UOTBVfUUmMKUNR0+KvlgGzutKyDhb49WBQnbio/j9g2IG/J
bu26nt9GwnXH1CpPLVn6KYxEvydfzz3GeH+BYPtpKwcJXkm3Nn9nfB2XJayzFzvo1LVCKdeD2qR0
dVNe8VpTeZb8OdSVUG+VliTw+VoKn9z8KI3eJzlHqshIPwS4wtYbydbamqhveruzeL7XJM6y65Ti
BWlevotKdP5ruC+lbCZHmfotgqrkANRou9BLpg+uDXec7NN2eX+zz+IDGxjKXkF1Fd+ms4+diwWb
tHKpho91D2TnuHWLTzvwJDeFeGoWWD49mCUKAOH0kYbrHv2ttP1Zkkzr3/Wi+Nv0XU+J1IqqvYXU
YYJifImjfzu7kcOb+jLAh5gsrO5jav+y78Sx7Mpffc3zMviP061WMKNMlQWulzBnVrd+y5EWoDge
A6MdhJSGND+PxQD240eZZVbuJuKv9AyjxERZTrLEFecRKEXzYqxwq+cn56P0D32p8ic8DiB0ltzH
ZPxHzO9UWXkMlnXWtB7eLD53VkxtF2R7ByNZ/vPyB1jsOGyiBIYZshZRECjkDEtymZlWQG7qawEd
j87hNwOULCCEDRjOmI7/FA3sP9Lu8HY5YuBgc/jt73nDzWXLoWv1Jvd2X4AgpOM2hex57MbscsuE
inXvX3QZO7fMZgeTKzoRFbMOMtU6lQ4904pe4dbGa4xOraAho0S/IyrPUutfDolxX5BHrvyuIbN4
3xxR0a6zPcTqFlG2QNY/qAZ8xcNvICNN2KPrxy0uujm1933Ht7JPHAfPSZ8vEc1eK3VjdCuCf0jd
if9PYG+yoew7gQdmVW/CG5ZkdI8YTP7W7iZpsc6ISbOLuO3x7tZSw7VxPtFvC1hUMcIMiTRi9HyN
ZkumE3YbPcb9HJetrGasRVPSzkC0fpJuyNld2KnY20+mg+7KDHZLkYBTlZz63cvfIV9jw1U4Zxi5
BJDguY2jKqeOk7bABFim4hnpkaOOTVX/K4+ehWX2IYIry1mHP+N5Rw65ffDw5G4E9lQoLlVcy6+4
zlsN51o3pB5yBhVy7oG7Gj6W6B0qoBlfEjM/roEoo4Nt55YyaJJ/euw6N5J4tkZ29koIr1eWnGYO
6JldHVrOJx4L/xEW6F4GGJiD1lU1a5yGoFX4/nJWp6+bEawB5yCS7+oleg==
`protect end_protected

