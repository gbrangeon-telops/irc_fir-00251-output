

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JtfK/+1JKYw3I976gLBlwV2xqGRbyVsJ3RDvlPNJRewqWZOfwn5MuTyc+U7c7Y8NUZJKZ6RY1Q/g
uXt328ut4g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SKJFICLwrmXfYqYNdiUThnnX5tJzUEdqxXF+PdKpwSGA61whpH8w+itTbLnn6xyBye2kcWPZGi5e
86BY4EjHm7kmXxm6GHfc5MWAMFduB72GxoAF5LRKlUMCOdVsZag78zFjXdMU64ClBQ4zjB8EgXvA
zXBqthWa876wjTEo86w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ho0WiFevcJjvoEEaYGtHkcW737RD7c5clzugQBBm9an3ZkyNmpivYZbh5x9redNVt0HOAIz4unf2
BSVy7qVCwKIsJQlB2q0JzVYTIfuco8FlNbrUR7/BeLSPV7XOk/MTxR/0Dg6meFJjnWuC3OrBGp8S
Ul4C2x7zg4t68SLTuFe/LzPmogzBzDfD3+nozb8sS3jX7ZaQAm/T/7eoy3grLVkFjUg9uj1IhVTP
59FDPnvyx1zZ/V9kzMjvM4XKEW4i0DGLbDEkqT5cZNTgcxi+sBHO7OnQuIvFzoIoNFONwh8iJ8xI
jfha3bFVgIjIJWFL/KzL8e9Uwq67H4YDz6GAsg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tPUgwDCRFsMzMdJqCXSx12cw+CNwvndABCoiKOSYIqrjgxTgSZ1CAyY61ekJUz6cu1q3fnTmoaAx
Nh8wOKV+UbnkqjbXLltbzNbjSEawEnAI8RSn8gStXvDoHe7R6pRqYg2wbvEPk6N6UhaMjVC8JxUE
Nl+LL/ApnNDqgvTWrcs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EyCeFS/0OQO1er1RAmOJ0VIpIQN1auXP1dzcGUAOeSe9eyc/jA1mhBpZ1JPfDCNxALRFgLLGYZec
wCmtwGwTJ9NXiyrouRmXyaKsTpp21jNq9KLTxpWtw00JZFdcekT3NPcfNHa7nkycvsM6yWSUR/cD
frws/8FBuaG+siAqTh5qClTqkxCmbJ08Qh/l3c/D5bCXbr8wXY+SVe6EK7TiYFpV2oOMuwWw5VVW
3m3/ZK4knJ1G5Nn68ZhcGx6rqQE9ZbHMigIgQyt/y7vXemBfmAZ3xkMsYj2X3k1fFfReGPYzTOCE
6J8z+FWVfzx6XMFACHDbKayB8gE3RAvjSqIISg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7056)
`protect data_block
3hV/Qidq55IcFtzIGB79Vf6DEBi5yGf7j08ftxlN/vBAWPV59uIWe9DPgN/tCSldneQaftOuzH+u
ciLQrbOPOoL3Pt+106uVpdo0f1kDQQXuFZvBqRUvkwBMw4Yc6ahzrtEcbCGhFsU26daCzsZbejvN
I06skoR3LY4ns0QcUdHRrwY6mphuTbcrCvfHQBbAyfwiiFp2iK47y8ma166foTkznRuA6J+ann9g
xCCSxWVsnYg+QirvRHUmWxOD4R5dUtR0r7kQCOLXWCLmz0FsEzIIfs+6C95X8YHCMPm0F9okrOuY
bFfcS7tbMaKY2olPSNyNdwRk6vOlhxonQcVNZZoB93MRMEwAaFq/C6oXnw7dLziKsfIWeOZ0mfxp
mMl2IVj/nrtzXGzQuRgWAsVB4+x8P2okwYk8tofj+tN0hlsbzO50b63H+j4tnco+wiF8uXNhRg19
Yw5ez/C6LJslYuohRhs5KnqMqc5cGwwzJZBUMD7tCo3FmP3BmZH9e/3RXGIsI66Weif5HX39EUBV
5CbNi03MlXrIu31ZseN+2UFTJYdiX9SeD4zbgOVES2Ws5cr68OKR5WyeEA7G73O/Pqt9JWvO/ty0
u2lKYGTqPGpzqAwtbiZhip8MB2h/dbdaGssH6KFlKJVit7QpNN5r+SbI/M5cGHBii6N84ejeVmAd
ZvuZHJmyqYrquUo926T5o2gy+x1m390I1WcVC05l7+q6vBwOxc3fJZS7nvj2/02Yfra+8m1YtxN+
J72fEXeTWMvnhhoruCmWJAsHTFp/fA1OVnB08oiNr+J81ghSv0tLft42fNn4XGc/EoSIF5T+3NI3
fwFyX2YlEYi4RwQvxvII12iCd4VX77tcUOKKem6UlUQzYFfXhztqV3zpECK9/wE5zxjZdOTPLN+t
yHZitA4VZjMoWMSl72jQHlvvNvIjKJuQyasTF9FaaxNxwW3drOIklopQ7HjzR0QavaMJQ07LGq4Z
8rrWAg8NsYLDoJXswsw+aXUBYKwIYZZHn/hnmTT4T9CLd6H7NGCHMZHBBPK5tO4HzP3tadUUO9N3
erOkkLBuEW27Mr1/omEeaXawJIhI62wbxzhevw4Z+qWPGlH3qDEppFMKLMVhTpW/1C1out9d2SfK
V4PCOstEhwdmQkTC8YillC69H1G6y22JJjvAVpwZqJ7ztrDTBnS+ncTcdVSQzI6oUhzof0yMmtyG
AsCqAtYfsAzNNbWvBV3gFC2f1WEWQP03DGEXmt4QAjIfyq7HFUBoqBc8nP97p9Mml3cZvEZRWELi
7KFka4rTdzN4DFywMqWo9GU4xQAfeY2yJ7cpmtRGKEB3rrKLcjaG0I325tlskGhlOWXqm7s4WyRv
jEYMJYQSubJ2Imht0T8grqUquKwjY66RuSMYIiSMeSMlS5xZ9zMMIvr0DyaEdzwIaWW+azwFadHW
Xi40FOq/RHBQ4L+kU/djy4Sx6FetIohNmUPvpB+4+pi0J15Rg+zUAX/TpvOwfHbdtOtzNmRFiAGN
xkKcYdBWhmH4QzOsf/lClqwmAggt5MTzYF6UHm7wKsBaYobf0LVTcI7pHplXO1vld3UAs0eK9EIS
Vk1VJWan7fpyMDHMl07GIcwRQ1CvaMOxZ8V/nNjd/mmoN9FSxl+YIs53XnOkkUEx8sm07PPXQVir
ciXyDFxTA/H1Jj4ZAIelbng/qbft/h4GthQ7Rd1A4Qm0sWPyl30lZDE/Go21W1/iq1HneVmpdogE
aKsPJxnD2z3AuaKY5PPf0ym1vdR7sAi7nav0iHIDiKj9buvTeFEhZ2aYqwI+6SmRHUrM0MznaOlu
0kxsT+j7xizriYx+neM+IrrsDHnuIAy9BUZnlnLXhpRmAZOCudFF2Cw+qwGTqOAL7pUXnR0VQv7t
eBWA3wiDzoBZSwDzFWtrIVXzE1j5fIni48PeQuTAIos7dJaoUM9cbmk8Z+dKgO3v1H0ZPnQDPi0e
o58d2PpnKUHHRoNmMARSNnmbDbdJRzYZFOEzirdoyEpwlIMw3SfLkkKgRijuE6rfRVniuWKVr78Y
mvAo6BGJe/eIyRzMfWvfwqK6FX+CdnmmyeUJifyiAibsmvv6AidtaXfjWnIRRR7mvIf5TDTL/sgO
zKVWSqJt/w5NNFm0iAxzGLLYaT5GWYiIPwqmad/2r2tlO8Yo8n7WP1Hugm4/CfLPe+RZ0GZ3mEBg
PUsz1z7NRAOpw3dQcBXXKaWzB8/ICeBC7LkkbpZUWSq+667Ud/tJHufHtdqwxxWdkSbocXecw6tv
rBB6g2N4EGF5+W6YE+MiJUCsH0T1hbeUTvbrp4UcGCRcBufamb6qrJB7+L9GhZW6F4d7KpMvMzha
fua53kL2sHMHtrnlufUtdhJpRZXEslmMMQ0YGPFcQ+PFZvE6JJeuF0qkakS0ddBUKR8yZy4WNibf
pOI/pp5TguwDBy9SOskvrCTT3OvnYEhrhfWJCAmtUIjjqceXBySaBDNuilOe0h1aPl1IY9ExMSOY
aHaEzW3/TvZEkaF1ESYvTGpVLJnHsUm4U0RKIsW3oWZrJJucb/RaNYgUrJBPHQSqqRxETLISCOVH
yrW9/FukgTE3KTHtsD11m+18DVt/+u+FnnY32D9iSHf9RNOdJcbDBsc4pO2WmP78bnZHtsyASnXN
fRrZQ2buPfwJ/KiXkCN0zAlS4lR6gE+m+wTYOTAIa0Cx2yqrxWNBldw3+p+jsR8Xw02fAWoA5P1u
VIysnuy9VzhSQQ8H6VKIg3VoC0PTxOjwS9KB2IFx6mPXIUYGVlZoEGM3OtieFeQicQmfRGAUBo1Q
HQb/aeOTNNRncMQdJkXOebLPEalSgR4IL6uYB1MEWpMllwCQ5NaJEt9LK5yjZq4p1UUkH5Wlohvj
ZzAgzEbfzlEVoL61AKFsajUNoMTRlfqVN0LC3jZL9xOxOXuiE42BQrcYbsohoff/5Kk29UkaQzzo
YoQXkMJ2KlVrqpHMpRfKoNQDUT9X9VePyoWeXbBAkpVUo95PM2OnnDAIYGvW+B62wp22Z3r0XqPA
KTYDSQotXoeCPFgPwzzbEI/GHOm+KIb/ZiPrRR2zFzhpu+Xu9vuQGrcFg9xjB+nODJrXWzTLwiPj
2bsgjopmC+xX2Nyew/66XFZrawN/xnk7T0JtcOiz2vJMMsgyh1TOibGq3Nzjvl5iWFAKB2iBYTyI
LruoOmn9VK6RoCaZkipTj3vksJCgp7Vzwkpl+Et5/ua9da4hss8AH24bZUaAKQidmrDRTYxVk4GY
IMrY9oDjqxzbqoCQk+8xHT9tN/+FVNErEmtvE88h7b4rZggfTJYAvvIl5bmKzlLnEmgub+UDcWQk
+ygF+JLUKFarDHnLyXcWX6vAPLAgESusTudEzwsktxSlasrpjja5Nr4scjq6XJ1D7OllULhFg8l4
bmwqMMRbeW2sGeWugEMo0TjiqzGLfJmIC1H9aiW1fCCZVyFnJrRHDNKsdCI9uBYjaSdpnTta7ikT
ODdCaf2JNZP6P/TDQKplK5W8Dz58y7o2IZ6TjeQrhLbeQeo2OfjZA66TIiVkcAq1fwdZoD/SeLOR
4APBEExIbBu7kYmwBtbxUUkOi0lcmT7YESTH9EkWJ0SgpOwCXjrbCkwXM7MXZsely9T9oIQggUgz
P3Y3n+HB1ZzJghcY9fLwdTZgeO1wpA/mnrGWyMMrIZ1fs/XPykQSFomk61Tg/HNk9fkLxqfpOWoa
bNMfDg9jv6qlbI602KILhhaVVZwA17M2yo6hjoVerDPdkm4fmqWo8rHB5/jmyVJF2b6SttyieDwJ
K568iJ18tSRelXVQvWBgJgRtiBiNp+yTW5/zzvOFSX+MKBMCeKefrW73p3tswvco+NM2RWemFiSZ
UTwgIbdzVnt7D307cxerJAwT/yXEHYdPhZTNkKoF7fBPAeszNDNQsNCaGxhkT8p3TyLOrta2ktd8
znRtdgFi6xhMoRjaIT31o9RzbaaVzRrAIzZm72Gamwu50zp1o39LxBw8OQJMvXXi7JyX4rx6c306
r9s/eIojb6hHNri8scnl22Qdbeah4nXgZrbVra2Xd8UJ56EkYdUmMH9+GxnGfn9bpZkh9g+B78NH
eM9KmL5wLsgh1nClnhhXYvvc6OjecqVelIOrcUtR655nMiuZSwURReoCZEt6UoFDUrQQZ44Ri9qh
Qah2bepVIPkwC12zQLw1S/yP+fjLN85R9oueEr6yrvMPFHyAui4hCDbWRp0Zq8XDIcRLZFudEtdb
jjyahff8BVklvZ7te5RGjrTSJEhXu4bSHL0Ot3KoarVzc81uKQzmWJ5u0erwIASv+N7A6F7b6rR1
IWtJmBKrQKAQSqvHuU/DHIRFKWZ4PVAc/2k086539fqt3gNVjZe4p1BCyh9ucUHCi7BHmfP9c7Kf
Gsy1QgqeNEaLxpJ1HUxjx+5dMReK17+9ZwSitFOL03V6CbyYtjFG/SkMBK696JTuQtWciRJ1gkV+
jlKVVS6tX7m0CsY/ti3my3y6+6XPwVFrz9oy3hvsCJHS6PuIgAxbRkFXb8yg/9ooHgUEEdMUuFFy
noSYoTZ59F6BKii10OkD190kuNMgBjp5dECWYr3XwBpkkSjmJN5YGEMYF/1GHXQDaljV+OCtxhDw
/X8vMhshjn4pJJdgQLJMAU3WnJGq0bP7yJ98MxihGuhzsxb3Ki+vwiUOxxkWshv31XBbRABRAXTP
gCy3VpHNwF1myGtjvWyFdClEbDch6YuZPohOHGQ1tn//qgdbN+dWb/2UI33wZngebWwJKGYH+94v
OkIHrXG3teIFydeQEyR2Xk051bKkbNm7ewOFg8V0NSfyWPgQ5Gh/5XV44yKzmvOwfIZ8JOHmVe/2
TiDfNjzTazjk3Sv74hPsywR0cHf8fu/t8lxysD6TmU4mgKqt02im0mefArdTFcmolW2qdY6N5LMI
y7ulm3p3EjjajnskKg9wVOzZn9nmwtQ6CvlugcJ58GIe2DJn05jWVPv6B0Ktq/FD9TlBhxL3md7p
3ThNlKCtH4OMc6rMTjZYw5sr9SZ5qlllLg5LTo4Ug7aAfAX1BhVi/YThmjQEVwLlE6raYrkh4Vlf
Tg8nNLFaDZSaxAqhzxLJsrdczHbq6Xnm6x7K83mgQ2B3zLFuZh7bOX/q67yr9m3lqOODhq938Iau
K/dUUWCl+DO5Qk9nyPhu0TVE7vmzTulFhAtj0G1aZXCUoLlGkltR367KkDvx09m5q4jI1rgalwYg
3YWYmCvrnX6AS2KwiUTTpUC0d2IIf3FK9I+k/rFtvUOUGPUbxAiRkutVG7b4H5TkNMFbLml+WaR2
91XCg1kMCaEbBpEYiXgrxdv/iBiMWR/245dz4O3PsEnn2uQzLDjz8IpxPOKVnKUCf31CJLMIPLvx
R9QuaanaNrheVz6O23veZE9dJy51xB5+MmTqEjzi1MJO/zWWn0Hl6okSRscKwzuzwSE2MRaLk5s2
uWk+RiXeEHCEcE/wiCdzai51yotPNo3M3wZzY5eaTuBCrBYc2SbVl+3nrRL6nqi3954SDqJpxx+M
MNnX4dvgTiIjju0EySBrh3Z0co1x31EbwVrpCdNMYcZi3oBelUqkNqE6+pQ72uVHtM6MCp9/PKOB
n9ETZkfRJ27fB862LqQT9EXaDwEaCey4brnqCEV/VaJLpWAnGZEs4/l8QxKU8t7Bf/cdNTORgPhx
Gta8u5MavEdbpYB4rtb/S4oKvhEitl2ZT361afFKpAOkMYan7c+1a2Jsbpg3w4J/CykoNMAD2UVT
QrHSAOKeymvqo9RcW1yzH9G85VBA3MZwS7LcaT8tsN/UfdfYUIxlChxAZjwQoWHn7n4B5XZvD/Wn
1pDuURTU/GSeJwliH+UEt5OC8MJYoVqMkCfdnXZfHTzyCOr3kQbXbWVz75jQINC+wEMN/SH8oEmy
UrOf8MHIFvIlGl4QQpgrZQPGoT0JjhIP262tlsUQu/k0FyoAslmSB6TqyiQ1U4mya7Gh5p3atvp/
NtBHN/j2SLKaPZnAgMeWzVSbegPvuW2jv3sU4Q29cB8V0W2lqK8plNGgeKFwG2DX7nGL4WVUx/Oz
53VN2TA/J5GDFOBDuOHh0cyt0O5oDCn02ars4cFZiJBTFQFojoe3NNjT1oHmdhbt0j/LebY/yCZm
NVWZrxEY1cQZaS3y08DZ+Yy97SqbfvM2QzXJGotrCTOBClw9xzxTYZcAMQfuZqQQuGsTWgGO03i8
YSdB+K29EczOLdwSahU8tnlm76Pw5LdZeRTMOab3oDzR3P5BPcP9bMWhAh2HjgdawWMJqfTFd/Yu
LcQU4ZpWrmh26cNOCll78utm28TgBDXofiM2U69wtSCkEMnLZ9RoVsnnTJuSh89+rhi7sfB5rQ35
cfKxz9P7RrOvUX9IZvkszgr/sTvPUqEMMuVze7ZeZiCxXXHqlX+V2CGqIgoBmyZkKJNFn2WqqQN9
KgsY9g15LUql10NetnZZuzavnsyBqbb9tWwxaSaP0B5Hhn/kqb2m7JxaylM+XbQTFC5TBwx881ru
5f00UAbX+t/f9NHM3cvm6JSr+sABO0XjMk3HiLmihlnKQRLMnVP0jZYdfUzpB+pbgloAbmLBe518
EX9CX6rQI+i0XQ/lTUwQj4bsOmTb6yFs3B5FcWBhyJgYNBqQWJ9OfsPlCm9oUWEISS9DkwDMfzVc
pvL5IvqlyES8WLOUtYbQTakQ0hwgcmHm9mINagkhYdmAa9FeIi+wNzS0YBmvcfvsK7HpwCwqEYcs
IqErwFeX7/r7mAKXYo37vF8U3Qn3Q0gibWGBtJS+D3Sr42ZqEqWxwKcGHXCiVwmUO+iHX0MOfSHI
/oNjf1bgryY1+N8XgwYfg4W+bJe12eR6ISp7aibgWdSc/eion+cVTz/DAjHt+gvqwrZYYH18LYJB
KaTigqeXCi//kfxfHU69sUo04aPZ7462uuc2uplOYYr7q1VkXQoRf/H5GopgGoEYYK3r17b0WPrC
udUzpunx8uZWtAdte2d0qXCOnS2BNWIv0/OpNB9XEI+kI8XaYp513YwURa4I6OjSHpA3NUA0pryi
ad54G02N99IKEvmZSj0KsP8VhCXrO4dgwpOFH9doDZiawU7m8X3RDtuW6jG7s2+ikJ4HQ6r5d5vU
syQ/t/YXSkXEiFy/DrM7+FaQAwKU+Fjk5E0b4XTd6XW/0f+dLno+0KAIAL34MgAC2iXb4up+ahrG
+5qfcyvW2ttyNqzaXPfZi1qHG6hJn8yH0M4qtogbFxtbX1+9WvbaJfNx9r0b7lcTPTGcN0ikw7av
4vunuUHk6mi6g9vhC/2QrUL+JL7L4N0p2aOXgNXHl40aXvtTcIAWnbYcCvy93ezKvNgV2Ag9smLD
VtYYzmfRw1oApfSzzpJuVlrSwxMLEiC2f8/49TpLvVmVuyB31kTzSlz5jM1HbVlwVxgMg4T1pjVv
bJkE7Hax4+LDwU3AvmFxKcgeKmkpEXxhBnnVzG+dQl4L4htEEXSvBUMfrLdujLfq3O5rS/V9bbKv
p7irs34LUujBfSIzBlHeOMem40itG4qe4/k8EKjMUBLBW3SGXNuD0HZ+mYeUj5IIOmxcaM6rNPZO
p3/kRVdGQ2KisAfyyOKoCWtoqUH8Hou+2t9bUtRnQOf0H0U3lV05/UOqIW2c9KgrSYk4pYbRUMUB
EJVrbJaeaQiD0z8pCHVLdS2zOCFeo2WJlE+KJhuU/hkNuD6G0rla7mzzQSjA6LpUx7ajJqa/nM4c
+wcii+aHPP4VwrU9jQa/nu2mwT2zi9N0YM0LRQfp/833RnPknmHSSx3e6BMCclgMm4yhlc88auC6
R9qYRiPVFreDVwdKY2z6YWv1JyDI1hXN9xszZLKetrop9DGiwKnxhIFFoOOSWvCCtPwHFZdU5273
F/5pJOXct/CDtGv6PZOQEO00M0VZmf/bR+2M0jpAav+psaqjqeLc7270szmO6pmRB+a5Iqb9DTd8
dytRMnGETC9q3IcbCuZDdaka3r08lvT/+/jx1mzL+1TRAdyYwhJst8V95zV/kL6K55MVeI+Pe1iu
LKFYDU4XOVdrqTSjL9tyHqFkpZC/hzzt40Wyphz5tdt5QImVdeHBxFpRJs3BXs/ugWVadvh7fkox
QaWItuzrn7NQfGaMdiDEprBCVDbwEcPNz9JoCGWGuqhAK9K4YmANuSIfkZt9yxxD4Lrg9RXo5wsf
+ysOt1zoIz1e/0o0xSIc2O789hw96yvp593xeeiMHVRwq+huVp9zojLIPSmEuB1b4sjwuhailPsb
VTN2CzVYJLuC9PAW/tKUtu4zpqTvja87gp+1t172RFVDOto284AnM3sGQSzjQxK1DJqyuCMPVEq0
GH6l3/3VvDyICNnsI87K6JY+/9ckDrubwUiFYdYXixUDXEfa/FQmvc4yr6rMfwHgcizuoJ/opaiB
d6rIGCU+b6WiKQ0yJ8VWJ5Svy09UFn2vUQFqKVX2ONeIHmdm3zwlOXbs1BQyi8w3n83OWuSzGmOm
vG1m1pPoSFt2PTIvL/7fUygxU488RSp059Jev6y5vesCST0eaLI6Yo+RcI3Go1rhOOoyHcFo8pRW
nEk/WuJCHuppuYSghoh4zwV6L3Mi4ZU8he1kOziA64bNyopmdcc7R8y5Gjei00DzvYT/8YdPTU2b
JxtE7sBrVEDU/NQrWZzj+a9FowCF3WyH492ZVIUJpg1h5BvszdDiXoZRRWPNvc/wXgSWWzbIUQ1s
R1Mlxlrbk8/mrGSFdnXeKEqpXkwrog0VIqZre9kpTsA5JgtMEbnW9eqO8necLnAInSKthLNFagML
Rz41+0UbU1DSug1YI5xXnkcJg3VhA0mHZcWC3BPwAgabzg6v1mw+j1TQzugc9ZZreZrdGOdOh3tB
uTiUKxlPxNrcZysHSuPtI72lUmtl33/DqdRE5s2Zopl2Bs8OEehlcF0Irj2Ju+SiWTIh8P3djjKy
UsFrXTKSjkn09EJIJoAjIMz6zyk5A9Zd83AGmHsz42oKZIZNowvwBHLvZjwCSyaFfpEC/UFRWuLU
CynJtnZ2VHpPlMHzvKMJd360X3cRGG1krJyRUEfMFclINouX6xSU4IQsdsC9fcGIuxFYYI7anjFK
ooGzi9GnaSebn+pM3CEzM3LJg8xc1N7fKvnEwS+4aB6goSW0guCZK7KsXKXfF3MvFi17Ssr/xkw/
TI38OapK0FvPI5Jk1iP0E6lCULLem2GkPvScHthtRBY43pARUFPyS3EJrUitoxFrMDLZmlRq+4/9
Ekj/Gd97//Ux/2DdEngCau2hcNbgtZWGCkvArF6IckrxoR2FrZSLPomIlCofQBMPMSkCD69Ckth7
XI/jonLmzDBf0Y+fwOhRmgbl1I2CleFpefhOXqrQEZIhR8/wuvRz5KATxVCj
`protect end_protected

