

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hajT1eUvtcpbI2tr2ZpQ+yt3wRoxz10Ck0HI/Kzj20i705g6DeZcP+FvEeRZMeE3iSuhECQss2IC
TSZjW2KB+w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
i/I1IeDYXVmyWoncZmW1nYLxm0OqNFHolb3NRcBcmjKOMCITsjC1Wrr+uKyOyNEAzg8LAt8SApGl
0BkTt3hGlwT5vH5JpMyxisp39DIoQ/2rHyhelRgIJSLTMOjHU/hpeFRg/8m17ioym3ZBfIcVRSy/
8YqL+H+Sd5EIN7orPrU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZwMv3uHNJwRn2Ww5TFfON6zTPNrPAlVNsMdpIyHdq6Uz+3GTAES373CyUHUP+cjDCtRwMjqRzGuk
B23rvW/CpivFPlGt/mLvn2R/n+PRdHgtaqKJEYqkidXp8VZscndj5Jsns7Mg2gtWutKvoptc7/8f
8ZVlv3hAdKdz/jYv3JFkYYsQYs/9EMmUObpsbPxhccaLaqAcMcp2DPumqvxQeqn7235qfdKNrMcr
c6uFXng8fnfR9emT//lppNqdkpAUWD93PhLZYTwVVXcjV4e16eyGLhyZTZ2QS7WZbPAkj35kG18o
nJcfgFC/GO+Ysd8/MvmMgbWhQocjtlk9D4Q++g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F+8QLMkCmxgohq3I7y+DAO2INd7sZ10O4AWi5yw/qOjlH+MDCzvNaVws6hhgvB6On1+CWzlrQ+vz
8M+w5LD4ga5aEaF2/H5jzH7q3vP0dvfZN4yRMhZ4TVDJv5PjxyVU6bHIlNhOrXl3MF1oGoVIjZ6h
IEpVBqdC2ShJgsN6O40=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Nc2OtpFQZFg8m9MEwwFrTSX7PqIQjLT0ImG8RPKmLuLlbhKyDcq1HH6KjYM6DTZXkQahd7sF4tka
CU4JtMixX4Y8KRzlmswh0FCLw/Aoh3nJlGD/KZ3QsZu5KBZUxKy0A3ntWjfTg1NNZ+tsdv0ZU17t
6SODHMUk49BioUo7eB0yCXF8PR27Zd7koQvLbFKTXZjGgj0ayut3GjrNM8A+4/o3G/elRT5WscCO
qhmVtlygfHoMk7BWSkupTlNlfF4owb4C7/AqdxneLzHPlGWymyNm6olzMM4lJP0A39+MtJZjtTaU
VxxrhX4xVaQG4Msik48gN+qH3ORiExl++4Wttw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25536)
`protect data_block
WzNT6cERsmb/Wd+kFZFU3ZQegCskQlZRHwP4pirsxWd8Tfabq83ZGdYt3qp8eH0ls36e6VyMPy1+
jGBqmxMAK0z9l8zPTAKbGwdwGKC8MKhiKaE36ZePsKMzi2ifNcGNY6BrKwEyQXBnecd/QRpfh5tW
ydHiy+gEqyvgSDy75G+XOAO9i0O/38hk6XlUH7EHWrsa6BLHsJTHA58qoAx0/GC667Am7RPgN7GJ
xcf4WFjZy3/ahuT0Gf56boa2Hjc0BUHfAhypde+orhHF0+TrzwXp68zoSHrNm07od2aQrjB67vEu
MRBIOXlxhKUWAfr2LsxWFRzC4esKuDL86QUAYKqNRI9pIanzZ5PQP96zHV6wdXlMzpwqAWVk5Sow
pEpIE6Fp3+mCuR3I3Sn78WkXplyxO1OD3WrdUVSvoHYQdy69aUeeuZ33K2sPSR/Kn0cXn0Fw7ITI
AhsNJFN63Yru5Oy4KyGuES1ZMPueYop3Y+Bue0GMUhF96XHLDOyFaU+bWmTeuwqGhQrEKdz7Zp3w
i9QUhGAdWcCkFhMw7ey+wCVPZajfbr40IOaQWLnAW1/Q8cHNtdJxG+/s2zP0By+STY3vt23gIEcY
3moyaAiHHRsVC4dvI2f+y17XugZYVkLKyAEQ6NdLi7iBXzl+3nTiWGzbplqTA+Qv87LKGPfsU4VH
S7qD3ADnB3aNrKEuPysjd0TYZy+GcEWgZkREtLvy1BjXIYDJ3FMAaBrLbKFpTAh4mBfA5JQkjWLm
2UwqzdYapAGfEFF8JFqSg1JJyWuSC1rH6yAhaS9t5729Tkf9KDTIlJqm9p3KQSDc+ikm2zztnRKV
kRHzdkIni2vYsIVynpvu6Jh0MK6ICyrl8ohfJz0W5L/hW0w4S+cjIzBpaT9SR90QMLtT2QToQbW3
YZ2niEDztU31siIn/dqPL3WoZcnnjSLfipADxG8znVpUJSGaiCHhJjMEUco3Zl8gh4F8fUYC+uTY
pEFq/ReJoGZeThgcy3FFQvAM8+Xtn45Ci6vLU2offiCpFqNAxqiWNEKnX0jqlp5GNySoDo23u+fn
vPC7oiUAUQfUx8aRQ6ntfk4LizkhgEfe4aY9NfIY2+epEHlOo6fBmslQ2qPq4nnQ5ASf2h+iXBd/
8L/4NiCl0s/VeXYdG9jHRLJNSJ7jt43lSt+om4cRtz+2uiK+S3cEpfDl6FlxMFBIu/9LJh+tARVn
3FKgAIp6MaYDvmemKqiXVy/Qqj2EWxml9hzLzMVfIl6JV0GDLm9GlLNq4HD173u2hzYe9UrLOVch
3qfSHMtO0DBs5lXZdVH1UYOStAIFjlu2hZ02yZ1EPxLv4JqISSH5NaDBAVmG5TksdLYOpEm+QpxF
7/BCBNBwKW6AsS81m85pjfMfN2ulsya+bOTT97QjeA4UujZoXajcDh4Lc0L/a2RLgTJVwqcOxNp2
4lKj47VfJKaEk5CAzH2uZOLgQoYHbgrDuUpJt4bi1vfRk+2TR+cSz6J19yblzLEznDZ3R8JRHZdH
SOj6nSMtU2HwpIOzRM3YxwwSCdNNjZYNNoul9Jp13TzXPxkr/Cqql6x7wOlYOPfrPsAPNUfswMXc
emwJxR9K+sGEym4/aUfCU+A0gZ/rEBw3HwSTDPPhDlGRie5lDzTctKxKcM935myK6itPiEYwTqJA
5PfT7MJw12fEzfXl0D9Ts9QqHlR1Be/Ue3EM2Ypx6SqWR72FZ3sC8U7YAH+0owYTtHm7raUgLMHc
8wneHXxRxWVU6idBCwIgrE3mG7+gmKxl5btq28YUKmxwq/V+UHGyFWdQzfXs7DTC/lM3j6+f0u97
7aq6yyXMVs8unAn+oIQOne6houXTKds9ZOeeJfgaRubM+zngNDyV+Cp+zFHzepegspFUm3pGe80P
2prX822udaUY+Yl6KMAzhX3iUxAMc0vJbobgq/1DlWKZ1xpCAs/CQXAo3igkxOF+bHYx6aSIqwa4
bpFlDSeoigZzXZj80ftmj1XIcNFKyRkndn09CrSN/YHZyB+SPepGf4/Tu2oGDLpIqMYhCRkTmd+K
KH9qbcD9KynGA0lTK+f7Ewqc80PpqZB2B0OyfoSZHuKS3rWEpZ01fc5QnnP0Sq0+ORr8hmnwylOq
MlVYQnnni4Zb202w7looGhkEhV1azZ0x9xXAujdTYUqDg+iuQGdGXarYVuNSn2KyMM24Tz7ASy+f
czbegUn0UE7UHyLIHCizBlqmSX6Y/1vYW32Un3KMUt6PuW5SPAAtCk3qzcTO3wG5Y7xGiYi2rmWJ
nEXEvbXtI8njHxFYE2H1j06WNYVEDV6VZgaFqTL4NebKym9JNIzhKBJy4gvtAQIMPSxTcwoIEUw0
ps0gIA/n/HQaYOELvKYRCZzQMnO0ukQKe3oCkm5CurQfhWsEYKoBfnv3ILWu6NjQ6nmR1CQvmVWA
1zpp7P5D5WCTL9yo+0/n8F70Cwaht5Sg5+acTo5NMECsnS5S/O7RsRUmWzJuaBrUn7pkK0sJIHeS
u8gbwUtwkvgwFLRxbRpaUX1DsEQHDyWnnxtojEVf5aBvraQ0uHslt3YhOSe6Cju5Yn6+/uhOng0X
51p9Mi8994IwOJfm0HJHuZNYRM4Ies+BnfM8xZRVHuREhCqZarKmIb3vhwN/KXheGfBrLlAKEuXY
kY0aQsGdAkGZMh2TDp9JiEe5/EvLQIVurH5JQta3Jz4zNhugPefNdte/l8G8oQW4Zq42TWrJBAcL
qtbKES0EYOVy2eDQsvrb3JuBCQ145Ko3PFF9KGS+pJgkKsrE4izzzlqVIv/F89FU956PFY813CUL
mC8M4btiatZdrtbx3mwQNMlA4tyPoD0L+EY1b5nF2gZsSxi1HftHFw53OpVZk6AOw+/wWxMauOzA
OTOJ6OoVACxnJUJlRxxpBL6VGt+QLEMzSWkFQJMEMEi7EYrXZ0K9TAmNKpbRzl2KBJ2On67HSrLh
KYXdVGTNWX50x4WHlWIlrHLwLupl9SJdCaLfap53YdttHe/22C4IxktW554RmrkssevX6nJDSLbv
3KDzDfmf6bOeliPbGVL0BOOyS4CkbVn3D8h6cmf7KohiB71ZV29MwADqdPFV+yDTaqT1ra4p7sCD
VS7oSU3gP5DDl1mHtRkkXo4xZ+3Gtaj1XLOumQcqDuDXYMTFypEUM8eVCFs20cHNEtnp9k/HiLlw
gQR8qecvlh2HxdTZVaLQBmIt/+4UW99s+Dvm0A62pbfv+cAuB1YCt9LZzmQh/cpNrBa9EicRRMSd
yo1I2mdENddAQqWAl6M2tJwNzbHsJQq6d8faWc+PseuW2tf2dLETDwkxkXXpUuWyb5YWVK1/L9UT
SQIf+Jt1w3OwAo8f3unYE+2xBTG12j+AWLst8MXizfYimquBUA910tqTZFEMl5eVsT9lHrAfsEOp
+incL/tpuIucAP9sSLi5dOFSXVKnyjqfUrcAIHEP3eLWna9LehHfNyuLSqgNTTaVlkSt6A60SH/p
Y3ZUZL/T10SQpyNUBNz1P6+mm2meg7wKAhyC7gqX1JwwkmyHQCP6WaW28zf+Ds1ZNV6xLIhr3v6E
KiwDPrI/KOUw023+L8pdU9uao8CTaYjj+jZF3fOIVSmi1HXJx/AITCBVnAVjtP0QQeawcGeXf3t8
BZfH7mjvs/seK38zZt9QwhRr54ywvLEJoDXBfSLVMVejR90/ViZjfgKoo0jbTOgLgM5Ez3wMGZ+Y
n3lTtJOYR7VlwH9GX6FhqkrkE6pSFUHDx4536jgipxC89ZXSMQOsXbR+5yBlO94toGCPDLQ27cZq
jm+dJ/VRLrh53INmiFwaH55T072QttulQi3auph1EjnEM/+SC8mK7SeYPFG+w6S/X7dj7nl8USe4
wYOz8dvQYBDvgOQgdt135jrnseRzhpmjzr9Vq+DAosHiw7DiB1cKqyhC2pdtMeDhf7Uv8HMQKBk2
xFL1uzA3/Ss+YXTWb/wMyp27K+kNJ7jSaE17UpHbrTk0kwtUAkJqAdFHrAXwvkSSf1EQTqqZZTpf
bBb9R8PWOdVvmasIX1BNzPqGcRfAD12sLd+jM1eqiw5pImhX5nIvrtdANvO5w+74tc6gLqjtqmTp
cIyXTntbDG2DmlrXZqyf4fcb+I+xWjBMDISwjwdPcEusepFCrWaPQ/Ji/SMtqL5BKAv3ZLbKOFpY
4vg1YyGMEnnpwkk+TjWYMIbcQJzjEW60RpmoEAZiVPL2E/csA4L6x+pOuNI0Icgm8Vztm6sU8/h7
LVI/fcy96EQ/FXdPPbiICyzWU/YJIyMuFqts4kCpqDtgNxJsCkqdwODvG/YidB9Z229yLq7Aemiu
x4o62umbmEDiGTZcpqEwdU052tgV35Sia+gDmzj4oGnD1Me2Xg9sWE2qGqSPm5Gj8qQpeAhusHLA
+0LakScvnTDZn7QSdoQuGNc6+/p+jwD90peUGrk5MwiwWEmaP49yDirnzMC0mIGoaew2GlFJmrMV
y4lfFyYfPRrk+ZrQ+Mm6ESlk7PWa7lK4RGA8RpeRlFQO/G0LeNqwTd0uaiNSpeK2LyPDvM9lkWvf
OdmBsye6KNl+/4eH2KnxFeF30fBAabURjseo75qgkClgOdFtR9H7K4xB4k1bNYhiemftwU5L7y29
QFAwAvqEaZh3PZ4NxonzH9WHk79dcJISLCsYDWdNn6g9aljqh8Hdh1KedeFB8/rdV3b68PUgoqW1
QsvHXhg6SuE8S8huOY0LvG4cizm0pKQ8QT7T/FXKHNOFbyv9E/OaUyF2W2e3JTLvMC8x7WAjc+Ov
S6Q0ZFkQrS3eGslxF4KmwxRQhN/YFiXOtX1E52F6UBJfi2W6a+zRRz3uBHkiKrh0GAMqO3yIJ+la
sxRXxntT88mgiLDP32v9AyU5a+JWLma5mf1KYsK/RtFHviFayx79b9RmTpLepMtWDwGcZWYdnVnt
65I2qcemJoQFTQBr/LKiuoSJlfSRh3a7WzSnMoVAZMvDG2csmUgeNP/ayQ2Zxd4w/o/qWx4E8Wsp
NtWN6dQSnCyhBtWymmjiWDWPi7xir7uTH98U+vmvevTk1NvYDQi4r+KcGR0OR9p66jRVSdcXxwUH
0vIv02QUI06PRBrWBuvea0cqHPlEZcrUgmaVBigegKMcaZhGHMd4jaDLzXsp+2eSRGXH4f2C8m8K
LXmu9MWUuK2yVQg6IjaHX7soO/whgdJJ3NXdJN/g1ll4ysXqUiMZM0ICtziZcJMTjnsnVL+BBZf8
841i+WQINkt04YYfR3srloSCpDAJ4Zs4HgImu/C7xROuOaJSGbvjxQf/RFoP1QBGR1cu3LZNP9/7
knUBW+8xGdKLs/OQJzzCXRHW/obMADOLVGz3guyqDH95PqapldngsyKHMLLETOXZEqdM/W4/tV5r
dslADWzu1pz5Ct4RfR5ZFadMLq9Txrc1anQu7Tol77DQ03+aRmbBK9l1zO7CSQI44aIkhWF+MoKL
Beju3wnYKwfp63XrxNBgckN/Wv8l0N23KhOgMgesP7VkCGlmQ7PxNqVOeHovnBqglyhO8c3a0dMJ
ks3b8Xw7AOoTqmKpJGVMC3uZB5NtHWUZXHZ4fDZXtS8VZnPuNEknCsKTDjioIPNEQoBsltgrOICV
Ubacsn0KnuA9GfVOr/3SgglGatGu41RNm4cfiaRlQ0ZDCMZxBZbpP8NQb9kluZ5jkaSUxU7UhopD
OfKQJVcYD9/5XLYPl4MsxffG7U+LTKlyWmtUrpEK6D9xg4N5WwEGKHjh3e4uC4y3Nu4eY3bpFcWW
YlWWl71tONVYb08RImgu8JTY7CsvfKjLMGB3Ugf/paaVQOVUqEogTgqrW8iOgm86KJwWySnKMkaL
npZM/0Zn+IagkusdM3Js4EQoE73glp7VA+J2WVwYWjLkXQqed5L1ydl/zHTI4zBygzUHL9bJOmuZ
ogLgdR9lH1UwBmu0MFsPPPTBvqWUrrmWj82YOvEzImQ1UDl7rBZur7hop2lcLFu2EfsgbSCgwP9W
AqfOmf6TjWhRU5GTWLVNjNjIABfW5oAsKEMVtpN0gDN+sFKPSZjQ0PiE0Lsh6Nm37lHYfZl43+9Y
WJh3YNs/kbpOyK8z8mqR5V/a56Z2Vx+V9wx/tUzRyOrtQdHKwRbhJEM9MxyMEY6eqapBR6V0R247
7U/yHVJSkUBeK1GyAW1xU03YG+yrOl1Iqcs3acFiwwxDcuFGwoNsvATTYEIYQHqtE14AVSC5A6aG
bVml9cubXH+IU6x/n68smxKuao19BrZ27hQYOdTQ3oNfTCRFZR+mNB1k5SLOamtSN6Gqz8eNrpn9
ma2GlT1KioTXktNjV1LbM+25xd1qbimSVXRWW4y9bWiUjW+Wzipn0oY7S8iSllmcIGVLnksW4KBQ
ZlDPXU1Y7VZKIg3KvUhLyR/J8OHNMxRtnCNzrbq0t5sLsaaOntnE8J0m/g5NgNgkf3VvQwJPSCO5
fJsqVnC07AEUIU/LV8kmOmf1CAG3fXgXAXaz7iDWKX9yTYJgmOpFngv/w/5Pgb64hwMcaAgwuznD
XG25CzBB+wZk6qHS5o+5XxJkj34uibNnfYmzD7ta9PbjzKAcPe7WrFKw/8TKdAgofUNPJxclSKgG
dDRU9KCWozu2dMyphuQmpgWaxilydL8wSolzd4r14dGii/YKnDFxMZU6RV1fQxISblAkpzJAfxA4
NYDUOagttNLp4PKnR5EzciImDLxiFindhRVLCmPfLVRLCLtHMVtIRPpgaADcajjag511WWbNnzKp
sB7F0yo0RrXLaH3dcLNnx0qoEaUlFlgmC+UTuZhHwre+99gnR75F03GBMtqOKdbzaozXMrja05us
/PKY4Ph3GGxaB57DtlGo6u6SmNAYql6v17FREwBkq2TG5oTpYLd7D16oGfyDcA2QMgJqVDhOZRNd
J/flsofQBJ+4KzLjT8N0Pj6z0YGfQhRpBHpcpZ+3QrQoblrSVi05ObzTQB9BqkqchC+TbfmwfPsC
xwgnfFGREcEFrYvNZ0MdyouezjfYwAwT48CHX3I7RZg4fP2MmxPlEFt7xLoQLOiRd0/Kf+uVKkWz
LWQxg409HjLV5lM7Cii+pMiQ7M6TbQgMhRB/CNKMuWZ4D5UxnS0iTWGscbj25765MOs1bB1giYFY
wdmkbDhXgcwA6LB3w/sPBV4xxMobOqlSuupvITHNW6VLCXJoPo3n5L8IibFY4cTYr+R9ziA6CqZ4
jsS2JvOu/ilSiJqfXQh2XWB74T00JP11IbYX4lPvamX4WgBKrGPc5+TKALs2Q/YpLKpJ4SK1Vf1L
KwMYYhmqLcQs15P01y6PlYpSMuyYnzok5GpZEmaFIXZ8jnpPd5he9UUVx0CbWTFsgXuIrh3cdFiy
vhUCFVFCCBzgoi3ftSmWzzDt9+68tsSNJbg0/ohR7mX3bt+rY3UmkNLcruN6iJHUkSIhPMXCNCpB
l0cHReBO1fnrVs3W1GTySOQbifODprYqgWuV4LUjjEPPKGLW+PpUBQt98WKueMdbFIR5GFw+0CCc
4daAIHbd5LEkZCukYYRWVuyx1FBp47BcArujStnzd4FMWRP/IzkhyTHo84ketkqujRrKFXODHUBN
isv5ZCjjBLPdYgI839c8gf7cYAObs2XFFCn85CJM3NeGm09cfJmkos2u8tLewnMQSaToCJhGE078
9//M1z103xcwAzT4K/Iii2HJY+iFQ147Q+QLLBLc7LCVX84NKqCA2UBAsw7t2feBhlaRfKfKwKgd
u0XwRiGhVtCOzKnOs/JIgGNl8AZRScnH9/kmO0ReCi/9Re4+ks/ZzqN+Xjl5pAfys6t3gcAlvx7/
lyRXS7LRmyy7ChjzdHwzz+7qjiILcLvqvlIuNtzaqpW8dcOe1J+/S/nsU6fMSCxb246Ocu/jYfXL
vSWSoOhucYw30+VANzfl+I1ab71vaulh8ru+RMKE6qpf4Gpo7HYtsiYpWPHevVtxoksXGLxcFsqc
D2ZnG2YOng0PivHLRokSTVYCtQHvbDH02L9tnddRjTS53dGCxEP/o5Czq/x8wqbYE4jDZ0qPR49N
/qx+GFXOoe72DwbjID4fphhTgBz5QMmITnl+9oTzl5gqyFaNLkyv1a/YcmCoI+0lLfET5tEq5ATh
DHUyBnp2K1CLAp74Dnh5MPJhg88pH5bG3ukGPK1U4cbEJMnj1JDD7TGNoDxpswzVS460rrgWNDsQ
1BHoYoMixSZPMEARBnSTVNkOWN7g0xd1zl4O9wNy0OwqOD3CW0SD4T8C9IK7ErXqjZyfhsr6qxu/
rkVoMVt1L+DPYvFuBDw7NqcMGkzURnRs7AKujrQCWiy/9SndangeR5Me/yFC76OqLFi6aFsOjCvH
tXKuyjagKm9/O1Hib91CVTGa4VbfD4GhgimZ+OyxD7BINTIXcm97vK+MAj19ZLlzGwEPEDb7BCON
MZFZORLSEq2bMs4OtyDjVIDagZrRsVjFnp9+E6Y7AB6dqZkROKq+K0YAPicu32zOccoSf85uKyrl
ceffUFWkkUVC7YqFtI32MhA2RcnUVRCDJ6yEoxYjOEXz1+wNJk4bHHT3viEUEGT+wHMQLMc+JiBF
z0u3pTyRiMbK7NcXTDkHC7j7IQS4C6/Pm1x9fWLRyFAILsofm2oz0nrcLh/oEZOr06AsttvKsA4Z
aZFWVyBYuHHFYJ1OPGlx4pVJwLXOWDEwCgAnrXJxFWXKdZXbLicV0MyOd+fh3Q6K60ZWIGdhuft5
W7Ih9e7FqKwlRfrMgnmP6wfZnBPKqrDuM4ocO+Aw5MopbCH0pBe1ili/7uB4mePsItAa2eacujfr
fcsvffR2Jy0thx08hZSB7fIFsFSB9Ycd1+pFHCp2itUOQarLGSL0L5/VH2aHssy49lvqpSS68Jre
5WHdkbLUDRht+scy1fPoTaFJUBEz/lYjwwVD9EIRrlmMXly+eb9vUTaCOhdQ5NoWwY4exNwSssXk
9ehyTKUg2u0Qki6OFodAdyZhyrXnoQe1DLhJahavj8F7WUJ/wA1Yl/Qo7oVujqrRUQm+++kq6x5/
qCRNa/Cc07wT2BqOSP43yHmJwXVzENqrb2tTYz1Y3onPpkUwsFSwniwtZbFRlGC+au5b03iGt+0c
oB/1HwMxVHYkNrWoT4cmSH02WTscK+Bs4rPx2ojmbqFy+bFaYp5uEfqejx/6PVPmx09YEph9+iin
LQnlDJqY9DKbUU6o5E2mTO+GhFf96XNnDdAhbhvt1tJTCTYVmu0/5vOgH0ENA+rA6GdA8NuEmkll
Kd8iuI4mpBSe3HtENOUkqPbqjxw7tsuZ57lJwqeUMxl6wBLDiEMarX3X8IJMap2gBPs3S2MEdVjR
Y8pnXN5GBe9MnW//+fiu7wDe7MnZBI9hSKSyz9QnikjR3EsK33rGQexEgkpMK6EjqD1fKBgov096
AKEf4o49MfnWAzwHmPACjYYXefLVrYvW9aTu6Eh8FhF9Tej8+jcXZ42vb4NGAYaBKDqFFeszPPas
IIMnJJJSTYdaklf9jI41SNNUGFnBBEAkE3ICezrPp5f+/03vKF6MHxfqfzQ/nZ7tYUHmgT5cehyH
UKsIoAG9CrOlA6cpjUGHoW4jOuCuTB1nFgb5JQwVzrnxOn9Fo8yS/V0zVxw6wfelc/NSbxBuAmTD
K/sWF7WTX7alJX/qK1B5V3FTXDXASnT1FjGcMTN+Uv1saoeRzTvdgp4XGlKasfIwUAnBMnMwpi6T
BjYsnTrcPQNqCdni76EyPB+pKY3JKw7enAHf60xgollqQxC+pZx4n2CmiYipOvO+p4lIO5HXjLyO
jWdHbg+CMHfgOC5afaPmgKP5G/WHFBPHA61McBi9hAjUELrjRzcOMdPC5RjdmHSQJ9JXJEqeD0Jf
YVB27YZOa1S9lAUYN4sy1f4ld+hft3Hm0blZtKLeji6goYqQ/vuz7ZPVDInklSX9TTUDBtA7ZtqF
xLx76TlEpfZ7SMXZFNO7AA+wAw1v0UmVape+84Ks7vbqj18kbbGZhmdyFa2uIwG0de12LZrekmSc
/G4giQRamG86Q0nAcGU6DLkiJYdPNjUiWWLtmI7Fjx5T2/97fgK4wZU2hwvJQ4JSWdNNXuLzThrA
0Wiyv4psWTapv2MwYYxAlfZJEb6N8Qe145h9MGTvTJDe0KbWcR6SzRFET+d5Ibe4YcSl1KKz/Rlw
SvBXNsGQmOa0ErRKQ9jQYedLiyQskpNuz7dsr4iUuC0I2E/Ectcl8go2oqKKE7tFjI991Wt5ZkwW
QHKH/wqccjsas82mkAB+if7626UIJ0BOJ3K9VwDoz3p61hyOineWLLGhbCIvI4K8XdnKc+F46lGO
bqXpfJ4KLzsBNsbWBU5tOXURcCd3Dq6+v+o3B6WTfZRaBSY3p/fQEaAd95MCnACrftdBezJpzVxw
Ly7WYyB2fsTXimqNp7CjyfEGxi76BdYlAHk92/UlqMEHYUrPz/ZvDrRePyHXtGL8BoLBcHfJaWX6
CpH+wuwxGNGrinamS55oFV0E2iE3pM6bbx/M2ZRP+l+EdX9u2t+9o1AKN5ugFmWRpfzOTPDhUu/s
c9sEAK1zv8CQeE/WVX3Cs2TITrxGil/yQZSFPAAukckzSYUNx8C8gkvcITd3Njxx/Xs8cX0NpTn4
KpF+Mf8GEeD1uWRTNw6QZvDX7rZVuHSzB8hUvZtF321ld3aopHQPiIksS0r3NY+wJkKNWXD7NKr3
ZMWuG8V9X0I5+p8XiXbgj+bkvqxJ1V7fo4+ZHm2hbhwlhlIeQvv3YDkXU0JdOf4BTiGpblSQzc5W
aF1qBBdeBapxrpUZ4jk3VicvkMHYS6aH/EnAyXpAROcfTzrsFFyeWz8eciVSjWDkmP6ghN6iJmuP
XCxf/CiE4Iov6VbsPU6X1R3SZPDOCYM0le8TXzqJy1x0bo3KvJzZ/65GFj1SF6x3581O8eKeJeKW
nyuHa31aPveCBtxB7I26f+DEK1COUX7XRiQ7Aw/z+nx0IHbLRJatRoNux9+vgXCqZ/mL9la1Ynmj
oN5/X5pEfds5dQUvJvyCgFtA8KkYnkYhAauk69k6GsAf3EhK67CHIqQPwKJLt0w+1Sr2vR+DVGPD
UW4ndHievEpVoDhT40ZeYIrLPzxoGrEm76dcYrptadu7oXtnP4t/pSgyR8VQG1fM9sQFQBKp/nv6
tIXOvrhM4GpHcPYyx4Oz8a9z1o3qfgC2yaYTjsvXjfIzGdsq3MdN6NyUc6wM4+bSsIAFtfaiBdHh
mJYeHBNm7i+qw7gioWQ1ajKXOQVhX0QGBNrBzvgX+h3ka8Ha+h31P6uj8yl9cYPDjQAwZOXMJUBl
CH4hIeengNw6wGmZPCpJ91gGPWF2EvERJ8GmjSLdNPwq2yds2Bqb4ZhZ3yowOj+yYYvTQ8IM5cEl
CPWpVwRybUO6Zn9idnKlNtyZCHGssZVykx8pX57N3icwZxwh1lbgieEVfC0KxZ5hK3Z1eiLTwYA2
p7PwewsY6aBpYY5Y2URurNqItxmjdBSVQgL/WPtZrSsH9g3MXgiLpoiC5x4jZuqlZ0vt3WQnQFud
7wAvtpT+3Lew9wTYQUZ70sKAiRVQ4ngjAsY4hIy5m8Lq/Vap8ThunEGK4FnHdUXMPcxrBno33qFy
3fidYKB08LS0o2sekEfWEg+C7HJd0I2T6fOCIBE6ihy/gTMzaigWLpWeidg8jj5k7knygKl2/U9G
aQz3yDQDNdoaV5Z9mXhBKgnPnM+B6uzatYRwPeOsWVrShtFNY10eLV0jAAOHHpMii6W0mKDiIX47
/zGHl6ty5vT8O7EDF6amqgetWVUdYufVnUFaXu+aMyu5fbcZN8Ai+7UV3F5sogQppFV/j3LHlUA3
QHfdKfiG/BD6J+vJSGSIrFQrmRNXuGJBpqrSbKft9UQOZ8tTtcaQuIPYyprjPKCO2sQlioOHGg1u
htQiDf87Cb0SQxHNdENAO0Y6KRwK5qAXP7dL5vFXUQOmO8FwHVyVBqjLJ8rXG6zrgmCicx7Na+8C
8Uru/I4lzentNe6Ow4KddUs9H/HAQCZLXAOpt8PIKBZ+Q4G/RGr+xfneB2kXdCD9FG+eyXbF7inU
E15SeOL/1I79BVlVwgIzMFM1jLNj8mymZJbIZ6ieJWJshwIsmQhUsd+S7nxd+FZVHOyhMLvbSYWl
FkBIoPFfBrHILMmJ4tclDRkHDm9z5TCmgI3W/RWnSsZliHn1vvoDG86pVqXtvHnQs1va55Q2OBIY
NFbAYPxfOpz5k2FtK+VmLnk6UXjPspbiOMrgpi5PjACxmeoVtuyfN6hDq/j80Wg3pm2w4P56Njmy
e9/XkpBsUCM0+vFYjpOfGXaPc0o/2Qzdkz+BVLhMMhqq+jLdTUqA1t77TM1PunkKVV4TTN4cIXgQ
APuDs1nzbjGPMFhayw4wtRserrk3TZarpACNSoFc2SAkmLfaeknblxi7Ty7fcTrjh9XDjnIkQjMg
EDoj6RpGG0++Fx6TZED1B5UMutGqzb1sZ1ez7+n+NKF2GKPZGZl7ZNsR7eUnePDdss/R8Jbsqzeo
6bO92Vn8PwEWx78YWAIvtw2NIkXui6TfGEulzx5YZ7lqwP37UqGJC3Ex+Qv9n9bMY+bmmMziz1EW
taW93Jk9xLCot5MgM8ceKfXWZ4ouDJuU0RqUiGnCklkB3QuZoJYX4cmI4YfnOvUQJJNPRnoiw0DU
XC1mnW0XJm3dtMtHhhuyW7kCCFCIJq8QTqD79+e8UmZx27zGAzowne8uR5emfwJdFhuoSex2FXOX
dqcvaFSmEordDa23xKADxrF+SzzVshSSW8H7IC0V/ktYADIuwJB0TqGLYRuh1dC0ktsVSX3/KIKu
p/W5zFdLVuf3/2wJrNZviOIM/GPa1bxYvOQKzNuoNkF6Jc3/FmaOKOAA2oe7FBrhN+cP3Vtutjt8
qCkseObMgKndFZepV8XE3YWEMC55Yd4ASdDqdWaF/Ua4T+BIUcB0UWH9ss7ES9zO7PO6wv9UYzJJ
OGPF6PfJQCcnvMQYRpSoKRWfeIZfCaN5F63a5r267t2RvjsOWSwtvvguzyAvpYLq0eFDWigDwVxy
Pj94ye9TvkcrQ6A2QVlYNNJrGMKC+dkqnuEwi5qDRM05l1KpeekXJG4+MSWlfDZdIEhE0UcadJmJ
Lq2LwUDiVwQO1tKGly0W7i/ICWCiOpJ0oUy0W+4dv4IWJ3PNEkg9uhw+kKyv93lhbO/INOLk4cEZ
DnL4oBmfVsauf0D+CpgpSWJ/LP0G8dka3H8DlOw/yDfP9nBkj6HG7XmWiuoDbI4DHgodvtKBWMKF
yBRB/lowXeC7mL888aDxsZreNnuoHonUdoXK/5HIZMUlhFKoOVX1ue0iq4cuajyRFGxzHqj9/ExI
bdh+rE8yK8Ozv1ra/alKsFoxi6NyYbPHEWlfyKWlSRlfvH5qJVb0bAFMcn/TnkUADNvXBf22dWqK
ybatGlNmcnXgYrUXUHh7Tg8ueGdLM1L2qAZY0+vvnCr7OjRNsmuBDxsFZaeNfCiykMzDQhbAKfYk
3itcnBrqafSP5D0ggmLMgZFCH/4cfiFOC1hSD8alFYGD5EnUTIqCNU9ZaZYVSDzL3+3jA3i2EPnQ
THlrRzN8U+E62nUnTtiuN+EFjUOnoRKa7RE26DleUSWqS422dcMXx6vxK+DZRIb3rQVFxIfsmMx4
+tVqmosTmOgYV8no3jeOjnl24jiJ+jXxZQPYf/cZ6FsYFi05mCA657/dlV+vGxCSg8wYl/IG7Zi0
xdGVKDaDUSpJir0+ENuHwEWWIvk/xKDyyMdDUd9KE+1+HungVopNzNiRWgmY3/Xf7ZPYvyD84T/l
N1d+DiKmSYbngLesAtjI3UZIU/FbBo6wB4ohr7+l3eRfxBL4eayT0V/14HIkJL8ti5Xn7o3ZwUFV
LgetBdUkGMpuE4Jqc/BMqiYE6/eeL123p60wwxjhV5p6su7wo2QlA99X0yO/aTyXShWkSEm8p7hO
hL4k0FKwmWTIs09du2AW//hES6VQ07+hEVjX4Jr7yYAi8wCDmAJxYCvJoT2tkA2LaVUrjqJn0mbs
Wv4jBGJGsaZAHcxR+PAxAnZQuJglV99JG24ORiUO83UAdw+Sw9HLdBlhKq8stzR1sMzcmrQAp5ID
0Iu6aHlZBETf7tVBRK09ewNc7BEM/C+ggKdNTDAXvuA0YjW7g8lddevkVg/mMbOzrLhWgJ4LUdyc
tBB0+h4OgMR6Gw61at35IC/d6ii4LmyDHSfAfx2Q+X+rLsHDBJ+yJNa+kgq4bKcpz9blRSmNu94S
5RaX7adeqQokqQEw2j67s7koqhvUfwb1nvpVJfM9vwpkEUr651sGeTkH6FZJEQoZZiYPf1j+NAKi
azLbS+rLBwvnzINfV2ewPyztRCeI7udezb4ubHAreqafLpdCJIqJ1Z2lAw7QdrkmwCGgcOTA0rYq
pc6HeR3Cx/q36oJEbx136OGYMi25JGPKhGd19t8ekKDxr62xWHzyWXbJK1YVL3xfi/48E3OC25p0
x07y5eawyfBSJCgI/ox4bw49xxbNDJnKHWUcNeO/r57Mic56kwrR6o0yVCWOczodELhSXTjmlBH3
izUepmJueNVWxScC2KnEMx0cUfLXM4OoMxyGf4OyGAo8qjmC5N8l3v1iYtCVtrFrpEFkzqJx/yCN
kIH2SFFSkAxs3Pd+4OM3wmfHaxSF7uL10H/Rywyf9a12y+XmNSBu1IW+LYDln3S4XXaSZTldkvh3
GZoaaoA++wwJ6pfmSotPoIAcKLq340HYDn1gtTyMY4Ly/DgYtkeDKs0n+KjNj7GwfoVk5+Nn4FZ5
mZkF0hPu45FhP2YcJp+GjKKHbfyOPngovLVE0H+L5lLIMWJ2cKzJVmPEwZCsPixGZtVFRKp54TgT
htv8z1hnHzveByv/bcz+xWleoPLGYSjwNHL/FvsXoygphyWZaFIR7nz7lrXUUz0ZMOxybsCTnkK0
6C7akyCBRslGof+F2ekbJ67IhzlvptNIAVG6KWBgw5pxnZvrXFYSGVlP3ycfYDD91DMLrFC4oBUZ
dG41S6wnPhlAElzIbSktGmRJE1rCwyc8gIJ+Z+q9d1fgblqe92exkmmyzFSqfXYodC8Zn66CFzNL
d3BveHEZ547m7mFYNLnnFan/4jqkl5w6GBimI7bkeQLo2MUuwD8iLMzcJwg780fSqqGFOjdrPOEQ
6YCTIq3nIryRpOui5x/Pxt5M3yigCgJ+jILDZkxztK9kWwcRRvj/qSg6bUtI9aSy5ev+wq5r052J
mHhY+n+Wb3K6oFXi5X9OEF81B8am9hG3xL8DsAbHz+2hC3KnJ9HD1cK7vPvhPqU3VT/v8GKZR1DR
jhuOc3aY9SR0aemRUna8Hp4js0T5cudjHf+EDkEzB3nkj+EVbFrL45QfaBsI6cROuLcQS05xaggr
xaqe6O7g3NwcSr2y96e9kBHNXm2dSwQVd1RzeEf4Cq8P5FQOL8JL5QtchM1viJXti4RM8rAXg1wK
N6FBRl7iqW+suMS0cH9SkdpDwGfxbsGQQUfoVniTUh3QLHeJNGSC1Keg/m6hQGl5TyIdyNHPtwON
KZAGpPp5F2D+SofIKPOJtdBRAjoWNFS1nrkjU5QM5HWXXANOrefkC7E4+ECYTsmS+xt8Pd5zjrzm
RKo3TG+dfwjwx1/t0XYB5vleP9dwOZ6Mody/qCsk/WZy8jsjkbrSySSRL0h1Km1sjUlBjrDcY+pA
riAb6FFugdX0l/fN/fbvAct3vJF7uRAIZ9uqFtIV9J1R8lN3QjClLYrN1VcRZAIRJkW0OD4zN1T5
6PI2mqeFkUw8XsBZM9RbPysiFVZzTs4ah0hS2F/MIHLx2Mc0fPA50VzOvSu6Q1z0A/8/tYqT4QHB
VqPOVBzN7CvPmniX+J9kfQ8oeIn4izJfi+nMwjctVLS9PwXc/FhlLjcZmWmFRiAFUCtav18iEqEK
X3csjg2k4pbjElteR0YW5qo8CrwJ4gdXoxU56Qcn7qFyFdEMtkxeAQ/pQd9smC4h9VzPdgI0GoDQ
/ljcMyC99+FuZil3zmew61VXewh8riAx5f3Fs5d9AXKY8gIsoVw3MLzVz8QvfqTWrl/eDSFalZTw
JgXqYlUHEduQuQZtruAx4H8I8VXVQlsbLWluAZPjFRLTKzHqzWQdhxJownC7k0kLuHWQpW7Pb/Mb
/QbNTsue8j4VIgADt17kKpwS/9gsiFJAhL3VMFKDkZEJMSb8sMcDHqXv0v4uYK1CwAFL7iqoBHh8
zAolixVJhVjC432q6dNm7hFqjv5lGdUa5cCHV42dfIy302rySv8l2h1GpE9a86ECz+x716LFTXqi
6uYrL4Lw15sS3yv0dqkziN0IjLIrKdtKxnfK8yQt8994egIfMHxl05lwsjBgh/ABSI1HdY7scqes
UjBGO24j4f9wulJaydrggEREAgFv6HC+qpnN5+0T2B5d0qqjy1/Raua+Af8KdlURUyapA6ZadQYE
+MgbIk7e8QJMVfqkQdtpWghtdij+FtIUMZdZYml9ZRc8ivc69bV9cBpOjlznCqye+/EnATZSQa+G
MvTrj7dev8gn4oj7yC3xVAvpmq9OLXw6/a9RU8n19ZhVXlAFfrOUSZeyl/42SKGfdqAIDMFyHAS3
nKs1sYhNqtu7NNok7Ssx1fR9DJ+f65ZaoiHnY0/ajQ5n1V5Gszmn/g3fLJ+XOQtnR19o0rWxazvr
S8+zHa31Aiqd71wwCtIGJ/5K73ILRhV/MeOAnGa6xA2Z4Zhohdkvve4v5LybiXZKfvlxWoV7AA/N
q7Ob3ppGhMIq+VQZ4w2t3I9uYO6vYCTGWPp6QWPpZrMrwU2o8j/DE0lO1pSEZzFd3HkwX/FEh/Kq
Hm/BnLourkvPkYrQph8wDQbMH+gs7rkgBSoNeAD+JUq/urfr3wAw9OC5g0iXDUGFkdPfCWeXjHpT
ZdlNomX6TgyCs8Oz7FyB8WGp3e/UWz3opKjH622wKRIhzlJIHxrtYwzn0dP3UOXYPTmiR8aSUcQt
mLCfUpK9YeA0dcdHZmBJctu83X1IZKOnFHISrJdcnOJ4+7INrCXoadjPocNSm5+S4VCnhuSEbVAu
A81SmlIAMXuTn4jSv77NlUsdCsLV2doMsXDQL1SSh0VtQuTfGDy1pEynMJH89qnaXGybbUqkjVXl
xWNJSWroU3iVpE3EgSHKqopDcMma4T74lQdX4X+IU1mIVi+UeCs4Y963Pl4Z5/M4daZMAfRfMr7k
AV7pYjm2Ajzi6Pu1o85xGbQ9PVQb2/LpUhWZnfl/HO/6qyeLupvwvZhgETiHJSLYtczQK43JdjNV
78PTJOmqRi5CdweKLthwP2Q0eTeQhvjsic3woGqS3bJFRNiPJRXqEMiwXm28wjc/1iu3UiDeYcJd
L78XrHiWgvLpeIXPiHTPBxenRJPpUygfZFo0F3kYu+SCBzRVD74xPv+DHxrtEoy3eGiUOgyGeHRp
dmfOOFaCEo2IiPC6yBg4HwvobvIQEzZHhk7avWTZl/2EMRZSUxR0vfIBUOiRwkbUya2DY7tvxQS6
Cx7M3hWJ5E4Sjk4cBPGhYvW+uNWuVCxhLOkBCAnHkLcxfaLEuo12XXIhTEfXcSkj8rpyzKG+/qnZ
t2jT3tTsLL1ZOtUZY1t5ojP/MynzGv9/BGM0cKBaBe1ipf3c5G6g3vXsuV5G7W1oTNbYoccfzMh1
uzzkkkGPL5Eyv2Z+07RlKdK8L50c4H2NLeC3vyBYQdxgCMYUvkWZhqFepuovE4vzpcssV7Yi6Y5h
uu2/oYwW9Maa1aaahRZqercG9R0eLZOSsVGxoE8X9bjy2El6TxZ04eWOxFbmWC2IlvUgOVEURLS/
YlGZndm1XanuA+QWKw7Ps+tAe4+BgJWEnLPsnXUhTiuymB1sp9vQ/32bTTw9wAjAqSBSTgpfD85H
2nBMl2XRM2BP6XnTw0LU8DZOufZiIigEly6pUC6EUhD7DPmUbDHztG1sZOyMcv+BqCzaJfHCkjao
oNkxz7MtxFltSFPdiBw7VYT5RoTTtz9DAsYV4nq9f1wC56IgLhPtBht0qVs+/ULUwv/i3TTrW2BX
wk1NUnYWxur07KBMZwG9ITsXpJi+N4zbWBucxD6eDshMR7w2/GQP+wH/KRKVuNYiT1CM45jdi7Gt
NtkOvnjTsuCWmuYM/2wxm5paadFe5Yq2HPWMrXOxYKuWQefIP7x7njkr9QRV2Yu2wGpkngcaj4p6
VhyOOjljfdshAAX1L26TXve6/klFG894sUOMOT6rVVvZJhCl/HQAAC59UUQCqHPXHpIBb+kkeUTG
Y7IhVawBvRbl/IKz5+oOIX7FsrK03tyc9cRo2zOeYqMdf0tQfRpWAwEv+Yn3FICckj7sn78WS14r
Kuqtmp/70xW5hwQ4vxFYGqRTGEKtW/GkTv71UN2px0Go3TUj59TiWM27Es0Dc9UldztlkjygZz2Z
cxvKXtAzDzmsiB926gQ7aWi9HzwKCZWwrFG0lzcKWEzw8ZMSAI0KJM9LuMg3wBy27P/mPMkMebfc
Fdx8Zb+yBjk2yNx44TfJqn4EqBcbR91QMIPbxBnF4Dddl7c110xKbhr0nTPeAcpprq+jBQbJrUq0
R5IlsePGZkq+bhrlaBlF4SwQPAXbuTp/bY7Fduby5wjYKRcRHyCpFZXguIXfcuGh1+9AbDk1/Dvy
Isz/PuAnJGI4l9QV4NpZwCzlWynJySLwk/GtAhhPmr3Q9iRNzejKUzJw7BfKAbZMiCNBjZtmK7ez
Tn9AmH6QXok2vJTrWa9QHE51jI8uxywJ/N+6CEYU+TZxpTrsiW+uFSX+lkXg0PChWERSWHGJuMiZ
D0WS+9YAT3n/p1V8FYjhZTchvHi2amufXoCh5Uk1sFnm4a7v3J27bst6BTaAtCdUaKKwpyXLj9Am
favNhbEPBKKPh3ayMARvkl+UhviBEF3FIF+AvSoKZ5PEtK4lAul66pnLmGDTCfE7gF+wSvRfJoTB
yqsoyyi3Dt/Nf7uvabvRiy+055f/H3st+JrqjjPSkNoHGE9WhjVG/6YkpfOKz3UH9FhtocALt9rI
5fLNtocVYSlAL0PtCzR1PKf5SwqHaC9XnXjZw4+/Q2WECCjwOtDjYWXLg3J4BJtvUd2h4B7P6R43
NtiiP9SC3t1VBW16S8ISzxlBktMnGB+CLI1sZuMBbEtRi2DK6Q0RWyC/E92W5xqAmhZqC0/Z+cPC
5FHOo2fWfAORo//2av+k0Q2mZkpmqqT8JtYaok636R0tzFS7VWy55m+UhueTQmJMsAB/ZWtmRdND
fYryzyuHsI+NEiSzWXTXKDgL+r6iwTJtasbMsBsxuwdNTVyBgW9CNseFwx0AiceKfUUycqlwvS75
9+VRWqaAc+DUB11rFhtu1Fg2hx7Yk35P2bsSLtBVDQf8A5cXrgXmfcU1dCvHu5nOldVpVILa7Ubq
v6IH40Q1baAqcRxWZ0ISXXss9h+w10WUAMjULStuvMUvjs8O4LzKL3WdwLoBNxsEmn4WZJV7kvCd
Crmkd48ETlavoiIsfvjKIS5NJWuLgy14fUhhieE6vmn5wHFAZycFpSDEOm+eB+RtH86pzMsEEx+v
MnioKlOoLnOrcvk18xF6XJvdaYRiVMma3BT1uTorNuFkFOe2D1u+FsndWARnpNj3jg5B9LroJS+q
QTfkAYLLykgQt+kRn/SqlbmMGZf5wNxHYtFlxtbanbTIanxSZD7rQcYLZtH5NV2YrOugm0MkEfA6
X+wHQsSZnIvnSJVXviUow6RCkU/qnrnYJI5oyDJls+rkwiItGB+czVHYrAe0Rt+jRnaYts8/H1Jm
MlOKliiOgGx3d7GaiOzA+ZQRz+KsY1XEm4Ahi92SXm+x/W9PoOmSypxron5u5xAX5NN/bIo0PD1v
EWY+vPzUE2JGu52b4TY2xcBHeruIYm41xO61B8E0re/yBCKfqcNEWEL/wk6ypFsC9zQw0rMIFMpU
g1XHz3eUOW5KHkjO5JQLzQSGOZy4AEfAikw1yHoI1z2dw8xD/cJ8kmZ7yshv3UNDFsGrorftgyiC
JZOY8Ey81VFU3WFK8rXlgjEBB765PrqAztJQlVyn+LidEEvm9+uR16QWJyuT1KJiWW5dqx46CiFp
jyc5L+ymv3eypj1F11Ls54fcqQK5J8c/DQKfPXGHCP6QnbF3iXlbfWKB70UNfSRH2nuyOvEDI9ta
/3N0Qw2j9/Ote42uFxl8ixO83yV/L1st+JfbK05TyCWGrgYMfcGLXIp6mVQFGZUz2xEmCijoNqEB
bzOiJkAnUGxYAEglSopmTw9aJM6rJfzBNJxOdy38IRWYAQJAxmkhFGh1UXA42c3MxwrfFFQAtVQq
QO8RK1LLZg5f5MxazshRLc9O1N+c+PM4zfcv3ooPxlnGIvUhewlRbYVVdxU51BLijv/XVy8yzgwQ
KzLl9BpqIR05OdULKWIsdosCLMUxCuRNm9OYE4TT6qno9LpHltWf4mXSv225lbmAmBQGC1cJfFja
B7WUw3lnZA8g3Jah+tA0J7a6Qv5CmuiYTkNBQGHd1KKUFf1Z3UBj6u1ttlPahwBAxwOh/Ninuy1b
/TLX5cFJV6CXMORg+dt5FjqT4xDRDZHKxXflcmMbpGM8luuCNz+sc7RT/BgCx9l8Ha/mZN7WTnYc
tLTF0gHU1+N8Wk7/1J3Ox6MADhJkjTUNEDwwwYjzwaF3nJZw1M01g8iTDTqEVkQkuiib+Ax/RZsX
FxLQ9x0SNcXdaPssrW1H8tj4LKTqkAPqqUtRpOoYNiwT/VzwrxZw9IAGjLU4XFUrUVCH2hvN2tQt
J/7J95CUR+ZtxAZ97YZmbZJCXaIepECQwtpMheWjarqgDeL1zXMgy8oRLpnBgQtD6aWNkFU1wWop
ZxaMuHplMwUJ31sEFNAx0DQ7WLYY/PyJN0HZMgYBFDl1AN/w6hWsNbLBfUjYjsliYWl5WulwVHrh
pnuv0+PMsgsqHSl5RD1YyUcOrQWLLfU4MObEHSu7hjs9/d+mJKG+TPwxM89CmAo7gJjAQSjrW7ao
AT2RyMc2I0q2npdC7zCre7Lhs5nbiKCb0kddbOmBlavqfXtdfoJDH80Bwm4irGYukeJmCQDOZ3nC
7nNYp1EP9FX6JxTdE1GAnewhrP+pf45Uph5ME1So9k/hUOIIqAbzmnYv9na6Yzmy0btDzjcd6LgP
bifvFFBdYFD2QzHqriTwuY++3FS7AA+LIQnJH+qX+g63ZUqta5ALFIQCaJ7LFq4tPns6S0QetAy1
G4FPOld9sekyKTO+1o2Yizi9WX+kPnZWQJwceqoD6K23mUYK6mXFgtWvwJc5V9Sbcycqw4QJIMwU
tZkpcdT7z63q+pZL9DKRNrVZpwgOof5h+CV35XzYoNMlme64jX2+bApTsTnUif17b6AU1uJvnoYX
Rk1W6jUmyDJtI+lAT9h4Zi757gHk0cZKIhEEn5L//J29Ih6RA5VLaNi82GElAZADzwKDc5zYvvO1
xQXsSmDxmmKT6Z/vj/gYkgH8zy4X3bOrK+dw+S91WrdBHgjldHUDPwZM+OHpsew3xwYgNI3RgBoy
bpqkX5Aaj2jOcEUyO/q98QnY2/pt6nBRBMoMoP3Eo2ne/zw43YMot8mqOuTtkaqLuoMwlJcJkXnO
eEjpxw2/hQZWdHGGkqE6NSsD6lfI64Auh+G+rC/P+vJfsPB0/DNF+pen1ohnewrpnQa71h0cjino
3ERO4d6FKqpL3Bybj3dCWuCSVEw0HCfHEa6iT0L5oLJTq5EiNHKOv0otX3vr7aQPduKbSrvTNF+5
X4tEs49nA6ONjnXc1zRzAR2u2Xbvy0GpIfA/I9MsasoOXALq4t04HszkMA+1TJusvyOJ46sWDISX
aIOC4U3OhfUwFy+HIpDP0DYdOcfdxKhUTaQ9/yYR6ttM+rQczxKTPU/icONiAYbJH95QDn4r02wn
zgfoi8PfO/WTGx6T5UTN2EaLCtMbjTbq1czNsBCFW48IKxF4j0ZDzLfw7GSoMzqavrEZb6Tklkdf
uuQdX6gdWyDvhX7DySHjgnOHXEwoqgn3t6oohuD3w4Fm/9tisC1HuW2isqTlcrMSyaaxPU/clBXg
XwJectq1kqLbIcDNJAd5nMv3b4gQgInkSOSJRr4YDfpt3tlrO4BfxbwJBs2h/1+ooDcye627xbn/
os/fE5WQu5V1XEKtw3kVKXOdtW3/H4UuXbW2DgJaEyi39+6SReT/r0ht0s5qIVepwITpq4dDT9PO
cMqmK+MY2zfpW53sum/57r5Fjp63W5qYRN60BTTE1Dt3VuJ7HN/zUgawaHChQPneU6rMGBJMlzKk
1ERdXXS/XhrvPEi+tAgu9lMT0ZDMrQ+JAlBcqqPPRu/+/BpK6V4ZKtjQt7UE89GmNDLe2K0UzlfF
cCeX6X2GLfHZVg7XjVnTRXI6ezLrklcs74DWpAkvEGpSc5rwur8uw//pvIvxurwFOcbo/rN9yh+q
5GNpluHU6rP2oC4L3utno6srWWoT6qLnCqIngJzkEY9im2l15HrfEPuyZnec/J0k4d4pVIMDhhdW
MftxkUxC/hCqwUAnGYJDH2BvFt3SyMirwaFVSZiqxhA56dbPaNzXJDRdAC/ykvqwdr1Sm1d3SCYj
V6LNIl5DUx/25bKuZADQYkhKM4O7NZu4ZLa9oBHiWEufaoOat7JQBngudhMQQShvKIDDQF6IfxoC
7OniOCTtoqiDOND+ASS2gePU1ubdP7kQz260JCS+ZaEPYw05mFXLqPpYDMwCn3i5MSqp4fy9iBOa
288YDP7ySf8fpYcbprXHEZYEFAja1OlDuB76CyhsNJ08WwK3c+AJFvu6dy2pWU8mgoBVPeABTSZV
jTk4lpozcmJAkunOSuPXqru1wFCbTd2ONltIAIR1IGnkGzlgfXqp65wenxE1jTm1iCoWuvHE5LbX
ojoSS862M8yov3MQUBfmQSiwwIlOOAVBTAW55UMbiP3tITDjxnclikiPX9oY+borO/hxgA848TxK
zw2LuKn0uWz8yA+p7xriPQukLqsD0wUZ9m79CpWBMzUFhfdTePYSMRB68pTQRq+p+NAAGu+7kiYI
0jLtHy+ncUWAZ1ST+S2GY01XVOHPzLxcas7PGmbr4+i5e7AYvw+DFTguNLcNtazaOR345lZ9kcMf
HceBBoHcy5a6UTFDGfbVcX7y+1pP3+oLZcBWiX+IHAcHCI0RizUQsl0oDfl+Btxs7kW8zZoJoN2k
Vfh6ptPM0qRd7/cxJVktz75a9alEdFvONS5hIhtPICJ/xM5KSNR2jlrUzPK8eQxUgij/dF/97/F/
FJv24AlY1xbyFBNp9toG4GpOhcmA/gnzO9MrJPQpOQHoYKtdAbQ091IOvk+Zl1GYAN37Y4pEOYP8
aioQI7BKM7zyX2ddxUadMbbOuFKIZIwJH26JKZi7QF+ZmM2T/BW2hHGxgmY8wahI7GS9fhjKffKi
elQ31knjbx4sQT8+f57Hobl2u00H98xDlyGEY+Mjf8Dz/Zjsbmcb059SAFIK++v7yXI3uBnJVePG
DkU5EBR2CilkNeSOsWY4hVSTPHflf8QIkxDeAMNie6bL9BOETGooXxo5sIylDTf5s4mdBuqFTkEI
e/8utC0XugYkxYSk1p2c4LlOp14t9QXot0hnUCzgNwwlREaFBg74lU1xbGg3pgXYQ//Z6eUDDMop
Hn3IFeulbWyP3wUTCvKwrPlstULcvcZgkgMfWL0V8dx/iBCjx+L8Dgb0gE5Sxq8SYzfGBOnmt3WJ
u3GGeIP2BcorRUD+gA0EdeJnfzF20oRHrWmqPjvp05E1V8d/FjDYL+RRl3E5xHGTdCUGRn555UQl
sgJ7PM716v7Nw98e5TwZEZSvCj7o0X+FQT97G2VsA+0fo+c2dAiYORFPzSBgy7YBV7RbgzlvGPgL
uYa2+0td3mXKDZc8tlW0cm/Q5bBYMN9+FT/RzeAOivGmDMeM42D7pjHtxhBFqsqRUGi0fZsKe9DK
PSdGlOsLfZLGWA3HoZYTpXkBSJT5JzMWWCiJ0UqTIPRtO6qXm0ZVoEtPPtX8MhNzhxlWYy78Rhi0
UvYUL4Zly+e3az73X6YsmyH3pJbLE9C4fD+Vvydd1YyiThJdVWQBKCmxarAD2EWgaf2WCyeHPuDR
oCQxuTPcT5V3y8rBlXtd653p1yKnUi1+Gkb1tgYIdjuEis3rNytqeID2dK0vUCyX/pbtHZooj6W8
+H+TpIqRmHuczW6punAe50XUMxFQd9SRuOSZYMFGJFkg3WMctmNiJh8cO0qMYmWIHVj/n3PuSjLt
kZ23D/CwniZh2CGAi+taS/0s6RZbpqNzprUnOmWvNvgnfJX/pzsQ0aaPMkI+0c8Qt31gveqm4Y3y
t/pRt4gpnDlJE3pgwYRbQiA5YsYvMcGsl5S75TaA23B1pY2maNjhCTqw/c880/vi4Txo4fyGFdQC
7Tzvc86RPNqlW6Cwcq6myzzANFdl9uQZO1ysESXMvnNaN2XU7ph2Agjx1geg3ebMU3Wyy+Fsde2I
wAHBeXL/1yCgPXyVtlA0suwtdL/7vgMV9lOh/MONLr+x4+3lbbvXwtV0b758uDsiO4uRkzuFsJa7
IP/kvM6xlNjtOnSCHujcPDqyDRrY4SC/NbTuoNmb2L6sbIZP5jKkPXNwnsEc+YpQfc4MzUf4QzaA
Keyy0r86YIpqaeXq9NI8RR0urX1mlrAWg4/cWwmFjZVHXkOmOi+J0+NqDqcZSVsfx6TGmYhuNyXG
hPaskEOqPNKc4b83qj+/nvaql1L5Vu6p5A8zjeI+UygwUbywtsbXx62wEUywf91i6bJsl+S8Ydmv
aVu3GkaSQF8uUsCFEuvuwboYa7lCC2VZ6R0wjbKnt78TkDCN7CBMdw/hOUBurq7Yr6zMyGTlU3/d
XKGIHXSJGA1kDoXLLFiTO3mXvpEWqCX8AzDrqsp0VTVt7JAL3PwdgLNUqiGKBoa/VeoqqyXj8xkq
USUWQmMlE6cuIm/qqUfSnXUPLBOylHHJLtH2Ac9gENSvbxeu/wchnZkaUUMfKHpHFnJOY0meHhn9
QvK5R4Xg56ezFvOFpR2IarX20jCPBMhQUExYWmM8u/5utVQfoZ9qX3ktNrYccyfqzOTosVpL8sVU
9AVxkjiePS3+Irsdn1I0Y4miEhFw8AEaDTEp3r8mV1R0pOiME6kUCPMlwd6MJkGduzt4lj34Df3Y
k+W3UDHbP2vOR7qoe4uCAe6jblPqGrm7uZ6nQ4nMu7vCvy+QCiGrvLP4jDccbnFWvrbaUU2yAbpG
+cD+mEQ957BL4bszQpU2Wj1yrnTOeDHWZBeYJGxkpA87iabYDXPg21lNL5W1z8F4kiQY5UkO4p0D
fxBPasRZ77XQvfPJfJWvvyrSzrMP628G5ykowFHWzcSKEy2/pA6GLORuwbpqQaoYQsUuPVFyIas6
G/7tbHV8rphGsICAeJ1+qoS3tOAFTPtTRvQldJh5hYcZ5wZc763MU03D5e4o7KRQOcL6P7VhGIi4
3b5GySz1h4qtrRLcvWy6/uh47mm8ajjJP+xK3MNZucp26DmcbLcL5miRPY1VlrsvPIjdETwBax+l
4zAqWPuuErTr2qqyf5lUxtp78amgyyxBfY3rfoOpkmbPU7HUmw1/j+wia2S8+c8I1CESiLTniC+c
okjIXvw9ZwF3jMAO8okIKrAGmRrK+dbed8mIW5Tv0eqTXpYqh/nTM/48VufTYZ2s/RG2yr/nVcxn
xyPeH+YeT/VgtRFQFl8sTdPMgbOSMHVQ6BTR4ABiIUImVHzm6V8tLOcd0W3fkNmK6VFu1keqB5lQ
PMANUWFIUeT9F7/Pjw8C27hd6SL1eysSL9jegdmkJELsAiEkfH7b1jx2QFgLYQ1eOw2Va5RkB0na
MMnHlfn6Oto3Q2M8rJjv3TKyooK6tCLjcweVDcs7T8Oz85lVw0WHIaFHfsyrzyot+ML3wJSLbh5t
j5Lao3WcNKU0D8BdEorucvHjkOOaC6T/oAm1BLo/6SelWG1lnohHPdi97aXW0O/XAPBbq6/6Ym1n
bUMc8Cj5cBkHSpQRQDFfXWOsPJVVu8HvxJOq3ioODCQ57bX31H06C5BCzl5DOLWuo85YxSCebcPn
MNNc8HRCpTvUoF6tb6VJDeqRC6Fc11PID5dssyzZzLavlJd95YNf0S5FZCYv2U2b5w5As0OsY0QI
95BsMXCjNwisgC3omPRs/K3EvHQY7OqpZaX9nnuiSyY9MD1LUz8/s/wEuvl4QrdSXQwHihOv6PDU
fBs61gAx1fUypWfBmCggsXO3fhGeVPIfStUIhdWelcATr3Bby2XEi+xxzT4KWjwaKXrXYaRaWih1
1VfJZqUdgZYufI6LjfmVJQFfyXCytL+KyHJsYkt7JnEX3JMXI3SRTTPyQHKEryDB0x+rCSXJlNSo
OekdpkSQ1NKlRLdxe6VzQ7gjLQhA+DPi7KmJy+BqmP589dFAf4g1QiXCnWCmm7RPsyYY16fZ9yjX
DnInBEgsE9imG0n1o+8R47sstrMsmbRgaeK32eX21rYEwcheZEW1/W/Z8Gf/1ZdI99MMZnO84YO3
g+MCODJc8Q3wTbJfvZnlHzuxvGsuRt8Ih1jiS3mX4g1GJtpsU4jhMsNDjzb1tRa7vbJTCWHttdFW
mjCPnZqQnGzYlkoasy9bvmlo4c59ikwGBdZIBzdl2QO1ev6zaCnWZ4a/+CdFvXiuddsuQNUHbe52
CaufOGoh0zqomAxkzucRwNdrOwsnRqWtQGZ14sgqAy9elRxFT47eWu2PmD+bORdG1hN9pgc6majy
t3V5gRwNSxqAs64vOTtjrmcTbErmyUocs2eo5vIxfhRm02CvcheTw9LG6osvK8Yd9ka5/2hKEawg
7RrAymxuWTTo+XtY3od5T+zqRdvJwCR1af4f+cY1xEvI8LNiTPTPwMoBBNan4qKvPzJN7tAbWgD4
jZLGxc/EvhFmvkezyqPJXB+/qoXsUnIhMjQpVQ2tQ9fn4tc6eGYAxubNzoHUi17XnBIH89UFpdZT
C8x5BFE+xJVYj4kKpCVM74PttV00RkXihSl6+5o4Zi+7EbuXZBJOKRuamVYWZ6bH5hwWm1/rhfyC
gIVJe44Ye9YFCbVsLJieKpNGLil0Ovl3pOjUszRs/qyl43qqoMSG7vb5kyrGOUE7n4HN5kptsjar
LeUUhwkyRlE6+mqUTV78LmIg+Gb+PwBS5iJmU4TJPy+UnKzgdC/zyP1ILc6bUVFJmdnRhfloqk8L
X+7W7Qlnryr2MNH7aUjer3/8ODoRetLrLJa+1iJS5avoeJ10ELccLoSqcH8IxhjZimHZgxOkkZaz
2r8kYMtkXqE1Yx5yY7KvXCG8sUa/41ZpffuSU+K5y5PAKtssVZvryZdUPnRT85fHamwT1ZCegUW8
fQHYgo/dWObQeKNvpSn91O2vbfgJGzzc78Y+v+Gn/iDK1bNr2LGq4iXEgQwDMowYb2tXwKn0fXvA
rVY/aDrNqqC6bGKfir1LqVeo0JxKt1fdfeAw71wmPbuqeukz8CIG5AP59ZZ65UPrW5dHKv/kq85+
h+VHQ88dQnxioyvHHBWzPKDqojyCcYzIvX5+ZEdLvlNlelutqUpsnHgA+kEz1xy1xD6YO+5pujE3
8j2W0N2mVBWnHZdDNr6c1mshB6CbkNIuzFFVPkujHWIpRnIVoDOzL5Q+mZLMIu8E4mDeBsl776rN
OCQQpLK58e4guK2VGCJU/Q9xkeap8yupgG68Lu3npOVtEnD13AzNsHXz/JgA0Zj31JXCjRwO7B+B
XiAfFJkAMOtlVXSaBlGeyvpn5UDiJnWohuCHxpDr472cgGDPQ5aFarH/O9mzq9OyAnaW9ZomSnYz
003KJRfIcyblW3JbsjpGYobdWGfOj/idzdrR4JxEDwkD+hjrGPrOdn50GQD+LXnbKhIRC3CR1ZFH
ppIsMVHs+mRZBiV2deGZHRIRmCqMrCGk7GEDZZTX5ElppTFqPlSFLJJ+YY/nfmQoroG0UQen0UWR
NXb4stCzkGnJeBNij3snSaLlOR/q9Ii0ZtOD+fmnBH9aOHDZCFpt0bc6D5AyS9RW7f7Rg8HcHnwW
JA4r118MdkwNiXL8FSZtxZj5lnYGEZkTCgMDvjikfJLjAW60i8gtabtYQ1g+xJWU+DsE89ZhUs7X
5X93GRiIv9y3mKx+KbXCrv5p1lPt7VdQcEhKJ4p2hNlug92UD8fpQCYExhUuS963fx/y8buKIcrn
qqbNEnwVFl9BPklZWryI98Zs1Hvu80X8U+f9eFXkCMiWrsDMlzNgTceUG2xXJT1JutFtTrhgawwp
1NRfyQ8bGYzeo2PbAiNHcM7mOVH0+nnArlM0ux5JTS4BfbYGKf0DpvjwEGcUsr59NolEowA+ZJ+x
s+9uSqjONBKo3Rv34AwJoQlnfx6r7jtfZFko74R5G54zFxARI36tsMEvq7wbMLxBuLLY8sdtHW6v
raRmUKeOqoLTa2efAXZ347sak2C/LxreXc5AkFoiIyIvYdIOdjN+fJj1WzCBytLeA3oYddFxIPJc
RJzBsrWyGgeY9+mEexgLDDLcrbz6tpswVJcjcouQoYmHUKbb1Y41LEsgJWnc0x5NMWrg9hvpiAAP
l0r0XsMFpnT1qMIfTvaa37zo1viprpa+7w5Iq/6MTA4fa68mIrmw28haEFbyG4UTukTSMZKRWsDC
4haBoF/sYRjqkGC58/C0Bmg7TglJWUuiErfwSIuvnQVe8T/YQJq/hIk7iMYzW3iGB9dd+9E9oUKV
Jsp5dkOHIL7sA9ptdvJJjZ8Co/t9viNjfUbNJlRjFPGD3l6paEQE9nGJQV6ufXvbjuRVH3WkmPA4
WyayTiKtWp5M2PPOx7SsEind/GyYUipL9ZoVwnSBpzcjg8LmfXQHSuq+JXj97VBt6vnt/PIw3v+a
khOLCvC6mQRu+a8cWaFHyXy+VqzrY/PdOJLRYc7JzL7zS/hzQa0WyBDEvbUitTYlU25PBW0KDr+q
L0PbrXq7ZOd970D+j8RpfjXvlAb1I1QD2m3Y0Zx3kI7oVL+qvBY25kq/hnGJ98M9yRsmtI5FNEUe
d4GT6taKaFyykcYSTE+SSC+KPQ0d/zxmWkyQJ0bvpcfO3nz4Qtt0Ix9wMX3RLUJn66iqcmHqW3X7
O2YfrTJsnOcT9OoOY3DGGGoYH0WQ10HIdtezev5pOk7kmzBJj9jY5P4JHTinkWF/UNoFOnzN3BC+
eT6gE0d9CqFwzT7xxiLcMTCpE5NLgSakz1H8KJqs8vw5Lt4JpEjQaHgFpkvXJyTDO70XG37EGKgz
aCo2bzQbM2z5OCfpOZfx88O4OIOWcaKkh7RSFtXz6Q3mq/RT96bJFjOkSEAPqCdyAHp8aJKbyYA4
K+3H2VyGWWoGvNU/ZSzibM0BVp5AEPXSy9RWTGESzeQg0us2k/FrQ7KC8AKh/qdVNe9D+dHUVIRl
eBi7BRUEpA5HO6IfvKFUK9NGTO1pwCyZusf04GseGyecnlx4riamaYMh7e++Z/z77nY3oWv26bzz
vvW3dkdZU0blBHOTqJOm7OneX6Z3aYY/IiEP36WJXmGOI34wiYuDUTBKqi9vWpbk5WCLzOace8sE
nDKvQoQBg6djH1g9S5lwC/4ceggvtNmYljthTbELeKXnmNbCxVP6QpWD7LkqRu1c4CxVWuqm+HMz
eBg4OofmCGRCutLoCgXqjdV7KCyiPLM0Hz23qBmH1fG9aN9vjSpzJFgeB8G63O821x5Jkrz4F/xN
SSu8eLwWuKRAgUNIeSpmLZ1YQcGl9QTg8m8TVjAHfQIWcPHDbOPB9LeHy5D8rSqc+rwKnm605Nj6
p5KGhQJ3zXPM9iMw4uJgFW9vp5Enr9QSPbA9oYDoQ5B16Kb7EKhnxE42xxMjUVq2hOF+W4nYUs6R
ybEozhi6RzEn9z557tu2E6GumXdHaseofkJyURv4qzjPpFvqVtB2x/vyQmJ1JxZkz+1w5BrmtHBr
NwXPHo98RBRlTWz2sG8bXOy9gE5ZKT2W3hMZJkjriCWSNfGdUuneeaVOzgwqX+F8ntxcyvjyxzM7
4Ib1wSa4gi4P8fm0AkQOqcbta1Gapu8ktjaeWJnbl2Knc3nIG1b7DbsPGqLp8esbyuBgsYZ7kVC9
98nTo8eFxYWzS/nrZj9Ygkp37dS8PconiVj4I1QknR8cKgNkT66PBqbKcIZmyXa10/smVldNyc0k
1WL97vrMP12yv5/uG2m/2XfcuV04M24AYAXxUnczgrnqQW48nsjUMjVhp22yBTyDDVJ3Lby30Pl8
VwJ1JS1GwoBn5WTShIdgPOHo+67ia6p3pl3KcI8Ccygx9i/tY8csLGnMAqnFh6QqyOkQKGG+Uciw
aHvS1vEIUfM9VPbPc7lClMWOGXCmTvPfqoltGXXiUnAqpKv/TQA0p2F4IvD0wJ9Nv2NFxlfFVB6r
219Hu1KicoPblGN30jB1+yV2WlS7sPhTnx5cl/L8fO4hQqlUf5ofLd+yX4fNZNIvywN83a2Nnapz
nZBXPSrvD70Y04jAtYsEiGTfaNHUqYGZl0yew2FMnZUhuL+DAypjq52HQhEvpLuncxQynYM1q5bF
dR3MQYGVuKomgMkAvdqM4T+llgsd0Kj82xUvmc5BByseYHzCgzOevMo8Isg7p1M2uHPvSfbpSCRz
5Uw8tae44IkYPUJ0WgeBmgRRSOX0itwksbak02m4rqUYy7U+2gI7dR04v81dE8+BTVi6wy0L6Wm1
i2riVu7wcCRiLbwlrd3cCylHlVmFCvg+U95joB/NGoAmfo6AOF7oMQlToZP3xRKQkc4O9aUwYaOK
MLJifk5dmeMm9QhPWcjl2ugQKqmFtxoz7qoidOf2iZ2K6wjkbi0KRPJFjm0bTx8yAhanXbPUIWdr
POuoKbftREGjKHkfx6CQoJDHCRwqzAu0bz8OQInI/wzp0pKBrEjWY6BNqfNeZnJWWgt+77y3OwTs
rOaVMaB58yz5dVXahw2zVBChuXZ2ZpWV+d1ZGbPklj1O9j97rW/KnSlGYlWMRmJP2DEOJHqoCdwx
G0vp9xZI5Q37QVS9EIwpWYx2+gV5dPhqUBiks8tbQk1O9lkqncc1ez7pYtITYfFl8yiFMv/rwDYX
Ycx0BL1i6aGjZ6poSsL/fF4Inkame2/LiNuBp6Nr/16LkUCkGOBFYtIi5EVN/p4GfqofksfIPNVY
V6GYNSH8JP4tRKLL4twW0OSFVylsKRAY9aiOw1XQxdpCB8XXmEZ9bPmu/UbbMc72PMrJOE8Rt3CJ
UbnjOW89LA1FlQAEZ2u47EAfPFgeRNM5HKEQlDH1OevKESkSwzFqm2b+TyzIPQNa99XLO50U7SAk
JI+5gLispDG07GF48MtafV26I5nO6a5nOiLk8G+aMWfknkMg5kG5bpn33BYXuUFeHeTnVWcrVxjl
ZudKfFnoEvQGulwSQdLi1wVIwsoqTUswWqPFYZVgYrHepwR3lerXkqF/+M+igfKFM7drJ2OyybxE
VTWiq7EpNZ5rjSg9qi1YA4WxjpS6F9mEywxoSWKNdENfbg81ZFKZkyTQN/HC/X3JRDTImCnhHzX2
3altsErBPsLqKkh2SMaeKrdNyfCg8K2qlo8LQCXlpZq1i+4Dw2Ui/FqeXHvh+aMGq4lf0uTYQln+
fwfgNHD9zgUBNiqoTA1XOTWwXYU9gJLJYOw03OCWKAkz6PMvjcI+Yrpuudv1UsaIfDroCkcjM/es
hVNBpynHvB7lrKGdiaA8cS71NhN9zuBqHUuTx0U0IYNQWsw/ReUxrM+LtSkE9aSecMWDjo9Bm86Y
B+k07KJE7H+4AGis5RQ3vQs9xUK0JpN05xbMUOGXdwCAs6Y4oD/McUldDtBdGuAmQotO5zwqtkAc
jl34auwSJDvdkX1miaR1HS2WKWkhYNP56vllfWhU2swzdCFy1YzoPK1VK1C3YSMxkRU+mihtrl7p
Xa0FRm/v9zpSN1cESHcY6vaAcrOQ+ICXGQ7cqgV8zjqiqV1IwFsO17U4dWhX3Hcfch47ZCGJ4Ega
sieaUXZhRDn+DbkYnjnsT0OHuBxjkurmoqKNNRtVPP0X1ZCUsD5TmXxEtQumEyk+0AlOlIYU6ju8
9fCA166MPsQUOT9lasY/o0/KsD/E8DbHNsW84iZz9WIjn0COk2KaFDtpJsj7x8tme/Z6TPBQ9o6+
ENc5sIz5v/70Nw2lIZDUN+Vy3E8Vmfv7GXOA0KmeU9jgM6UCriaeXl6UP5qoFCz2NXafP7PO+AK3
LJcQKoXJUmlfCMsiVNLECzVJJYxHc7oCzPMGMblbXqVgTTNSfml4VXaINaZZAoNjUHl/23COj34A
NDTddUJYGwGN/Adxyw+djqZDFc4Rp6F8rz7RvdZ3bVBF64KAqWU4Z6cZVZgaDWopTFjOksYP16a3
kvm+ntpfMGwNBfb8ZYBJQbYBYcLtZx/7oUo/grcJ5F5KzrZwVzN2TgORSCbvtfTwcO2SwnnTfaQT
0AwG6666ojuZ2TEKFcLcUZD3JFIK1WW5xsarmYF3XMW6WOB6ji520sbDui9oNPqFMnZbzGSYeggl
CPGJzxcmdb4l/lvmAZN1SKgrFRVMJfbr7ExGplpK0mtpPmM0cTyaWLSqgno8CIPVyQzgUEPaOR1e
Cj5MYTxngIcnDgttLULJ2Fh0mvmEh/oT+WmjihNWw+h2p2Qm5ySoK919wi2U870M6pJGk8vIRJYX
FrxiSpzt/rvvlCSiADukIn0TlqIz7o4vkkz/HBhDs6J9421ty5wkuFA7ecKbegwngT3GB74ijnJ6
cdeRm395ACZfGF5ji5nea7qSftF6iuuedSIhGIFX67GUBccjUwmud602gBXF2UWxdKCIvRjJxJ5F
tNGPvBff+eAJ5z9DZyCbAivKvgTLeUCfZPvJmz6/nUkPPxv7Z6NpWPydQhqd4PoQUdqSedW1zC3J
XHtHc5rDWzBYgn9J0qldFHyN1eWSff4dgekKn58Z4uft9tm+ukcbdifBh+U21bOBlPWkv1pCGnvW
FQ6DM5wRG4h9g0N8WQqVTM4Oyugb2Ru1Vx1O9TT3neErds1/+iHTCzHDxn+t4Imx7l0n+f5GMYxI
u2QT3yy52Q8Nmh/+rISCtOkjDRQ8IDMWDIrvu9rGRcWtDeoz6bDqknTnrCgbZu4QEiI7vpOqfNa2
tsPbsngTnRBwMyRlfDfG76RcTfxCGYpklO/nY9OewWHr/kvpw+6EAI26ubeUnmbEqqca3a7+wj4b
IgvlWWAzj2wiUWGOz4i45v9x76U7Dth6ZGsvKDn0KfXhSLq/SOdDofBNspbrCgYGkMpOCc7abMIY
4R3M/IcnxmJ9w0hu8iLbBviqLJE2c0dnVCkUcrS4DgDXSFuYv70EGkIpiELyxGzKYAgulGJycBqK
fSxYd8jbu+dhisexckTh50V4f75X523HMII5GAhjLXcM+yshk/LepogkjNCXdM7rLsdzovMIWje2
5ZPkd381m3SiOB3fsoBO7fBKtDErWwlMYM5xXrTDouRcunozPMXGBGdpuPTqmbJxSr/hJwCmznRf
FzXcVprKilkh+dv6hIUJOC9yLPNMD8nmjBA9WjAyEvMohqFpI/R/DxBR+Mgs8f3zj7XOETxMAIvP
H4M/JedDYNFhI4BB/33MeOEHUBCk0556IwH53OEriLtMPPl6xG70Es8RaYAULXAUqFW5MqdsF5TY
qBYzkBFIDDiNnyHL92bqmvVcrxVSklsaFwYQvhe94/oJmRuIUGYtNnNhY8j6yCdinE4/u1qGYd5v
eQdem9bHCEd91BVdJc7ujPCkwHI1DG1NOE9nMEH4nlMavAN+1kjgxq8p1M/tOAdZrnmKgGblTP6g
lQe7o8ENy2OxyQ8B7BlUhkR/ROhuN5dfZsdgnadFsBKl/tzPkqi+Jlo8wKPRk3RNfZCL3qux7Xov
HhNcl9talk4Y15Tz/Bz/FR6hBPI4KTPwTSkX791+/Kp1WnsG76iMZmokWJRwD38t0J4GCB7m2FO8
`protect end_protected

