

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CJc8rmbxQK7PiD9FE9h/V8z28Q2yjtwOLUGOHj92X0D4bGhAiTKxH6Gs6WbTk3x8dF6WKWHXW0Xd
imaqryWs/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KUGgnJN/sGLwh1pfD6BBRkJkdz3qYXsMmFAG0D8TIT3kvn1DM/WYFdJfNjuI3TZJ+GjJhgQt/TQj
vszszvccproNtKL+iK2kDAI+dODbmK/3dk8pZpjNIY8iqG+SZd4LOHkCbGnDn8J5L1SCb1FbgOpc
lYLzGKyKMfpMp2H5zrU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QPilQnlZ7SkqHJ+uQKxasOWlKPf9SmSQp0r8PPqOPGeQK2aUl+9gzicjiy17/DdQAM7rwf++nyUV
Yi5HrcGStcw9bK+k96zmiNT/NPvXPX5xeKvpNagObga/il62MarkWpibvt8B7D5IQi80Rp8/xMyy
QM6+TtOf7NVahw7dZAUwr3krfROulZTDfEY3oalO/PlnwAGr4Z3udXzac9NTOUWxkjpW4cmTbWcJ
unHhHJbyMO341XtwkTUgKReezgKFOpi+gREeBT80YOKcPQyjGyGuc28HYVmxKisVh5P7BYL5neLX
P5GVK+HA7MCB8DsbsorDqal6rxwDeaIF/kJcyg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZE3LPHWjt8FXIcLXD6pONgldgtzqHVcVbUx4Qj9ztf/3D9DwoYFB/m8dT7Cv2OabvKVMu13QC5lB
rxR5Jhd+fouVouDNKYwIESeS4DEkgnwfSJpsmeVaPW2tqCd21tzGTVfcw3Igam9PcTjnI1q1568h
X1Tcmu9paLkGRwvQeII=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EV5YorhH0risCTPPpyQGO+wsA9egdTVjrRAwQuEDG89jVsb2NsTih5Y+XoLrashGMO3AtQzajDhF
KB2YGM3JfNSzKu3jU5R247s9Goe6ZA8J4KFFzdwq4blriCHlPX0eNqXwJaOF7SeF++njAnDs0TkW
tSOb3VJRRI43LgFv/CHX80X62oIhRm2LIRAjPrPj7KevSjFw7diU9sSURAffWyrhgq3XZsUY6ovy
nAWzeDeWY3xrRDkxjxQAN8xOlyfUxlNsf7am6Prp3DCG9ANkw/MCyfCVBJXBbghP4T6GS/pNjySW
+j4cMtiThQqIcJCHVcAXQA0FAf6PbH456gYJfg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4624)
`protect data_block
2zO6LgK/HPGKSlyu3HNnMrN2IKl9+5rVKhqtQ/eOJiwVWvre05ArrVpjo1rVa2f8mFLdIsGkmY6B
7MgyKMc16hHZO9zqi+7LGrQW6/w5yyY1OMUEJdWs2Jfpf915B/upUXoDhGBEtOGkMbacdMSnHyvz
qVGw7M9aq6Xjq4YAkw3swOQBJ51R/FrmHflfcKUCv7IEUTNPcA2k74z4/utACKRqy6fSjqxfs7FH
mBSQCgfISdRooGfuSTa0FSWIXv6KmG8DvJm+O7DxXFUiBPHGBme3vv9SdidFYOEXQqTe25bXhyaO
lwcQebS1aFdKTnSHDGIq9TWBjVm1q363H/Jom9M32uCCnqcwx664zPX0aP6MaKgg4JlQ0i8hG+Vb
pTGp0w23pZVcn2mXDxB7N5Na3WY9oYZxk6ypIL8ramoCOtMaS2a8SzAPZfvQnal8fWwlkucbZbmO
MpeHx0dobualV8nx2UuxLRihVayim0RcpEv5tL/caueBdlPpqNu3mpdfnS8Up3Vl7iHq1wmBpWDB
EIHNY+A+kqIu1K1QKG9BhS8tHqjuT8+f4DinXbSXnOzMEJNaxo2XxATrybWBYvAbTdtw3pHzHfnm
GQSttAP+nkgBxKZ9XVJJNrCytfPgaqgjNPASd14FAuiaM0DaKhSewT1++BbUgcbqTpMJ6kxlCAZL
nl1Mpk/A+keZ2rW74LTFqu/UQYl4TWYbxci3NYiw8Puah8gD7RL4wc2AhkqrbLnkKWwxgqkKKWey
2bFTKz9jOYu6HUEoTEuXAdKCzVDgFa1RNtnqo9ysp8fN0nGaKZ1U189kB1MvSl25idsJPxivn0du
nQWrB7YX86uH/4oQIfMBnpiJxGbPk/SSVQM4YbLtZBj/6MRns8BWk3+TyYZpurC64aT/NioyYYgE
+LAayc4ForV8sMEoUWAmE3xqgNWsvGlg7zn0LqHlHzxK1qEcr61mU+0xC7IKALcRgO7jasvv69UA
8y+libyRFXcNA56+ITDJT5C5qlt90DR9UQwiShlMOXVap6dzoyD/Xo74s+O7Sv974GzDvLqUZa7U
Th9B6b+av7OGucYdWeU2yXicv9xDHZS2c8Z6EKbY+NUCYaqPfx7d+RdDdEiJweFeXGIbKDSNTUkr
aMAg+OxuCRYhRzpI3PpAzCmeWLPStCV7iGzggG6ljEYrA3pglXhdsgp0dGDQX7X84t2Mli2i7ls7
JudUE7xQx/3c7abRaHBl3PufM1GbO8JkNgDv2G/MktFEXpTLwu2h0Du/6nnqRODyWNLs5yaoVF5y
ovps5fJiegojAKBLtnv/CfurW27FmEtbcqN0UDDWh/wLcI34c0olRE/0gPRBDTCyWJW2gz/s/isc
+++uYfZGQKZd/LDprHK0Uk42nU21y3Nn0Yj0CY8uoTjRUbpo8rJm9CzN7bhV5mXA2THtLoktqjH7
6c8IqSgAQSbWaQ/WSukhtv/JIlDuGnVv/U9mYDXg52RLD7wrz71VgB4UDIGVFDhDnwjZuswSFbS+
jJwL6/4o/+XStL3V8+jRdsgyPjSoDyH+LCKbri+e92tNwnDqtH1h02cH7Q7oY88fAXP1q1UWHN4n
QaP08QYCjPJuLBnt0viYLdqYYHzr4E91uhSZ2BTMLOqzInE/keUuGzyR6cVS8RxUkFlJyg5DVXTY
KYfT3EjIDhJSQqWau9XxL8ddOAG6Yrj2Oic7t0ORb7VNVvbSA+xdsEaesYdykCyU4eOQRbBrSOMi
uPHPNopUj7jorMVynDpWRPtAvi+YiFcSyWawtRDdUVvP439eAxVQZgSOyDgryX3LkTDgC5OyenbD
E9xDqVAGNgGVAqpS+G3lk+K1TuC30rHxGm38uTUNrAYrkXe5AGmZuvFS6Fy3MAueCOeNE2RDurX8
I5/lUIeu38CoZA7JlhorprLRBLN4jIiklSGHA75oiAxUWPVv+52IjeIkcEOhwX1i1CEEPmdBHsGe
5c3fTPqzEBkMgD7ZqAJ2kuIf9b5hEviIZO1Jd2LBhgLHoGmvZn9QSGCuyXwg+Tyo5Rtd6SXY1jvP
52qODNlxaanIhasWLC2pZnm5foFF3zg6bMw5/vfh9tzhGj8xhyAMjIMwFCWad3Y3DXFwc5Dkyxas
XRd3x4v04pkK7cwhEjR2ZUpTAJlBN750GlExHw9cfenEUkGuP1X2eweJqnOEQxKvHi8uTug5YXkR
FWoc0aOkbiKX24sUFfGollogtNXyLAI8uOvAA6VmfBAyUPbjN6+x6jUYvr+VJlU8K45gk9wx9k3/
K5DunP966J9+0Qc/SyQr2BOmNHU6W4hDgeYokGWUrNvgNDjgIJBIluemM9NOLS+O2HPswdnXSGji
pOc4+xDxjmmY8qwLEvzq70xnAE2Xbak7+LxBK7FesZPu0ariaUJXB7qvVchQvu2tofNHd+3fXeb0
k6e3boj2KP+ORU6flaM/2SpP9rUR6h3W/o6kEJlLvy5M/2lPQz+CvIuGsDu0fCQh7b8s3Xzroi3J
XQNmyy8fsE9siDpMArR8yiWCvgd4jt16mOi9fgE0a/PVTf5JiQzH8r/n2ztHxVDuZEyHk2/dLHiO
ZbrLIc3FJUGAMjRAXwyBlZ3fH93XVTgNBIedlCy8pwPiz+ITfYMG6ux0vyUAlD1Lqd/F/3EMMmOb
MWVRGjpH1qlk2c4z60GzcLZUtd749AnwxeTp99LhNBzZNNKuH4BScfFi5hYyUib2LaFytvp6EK8r
zQKh6nZ5XNb+RKNWKvKsUS6zRSk1vdJyiA9PlwWGeRmEezyYOoS4LiFv9/pyRuxs0u6XZygmNyWc
7S1GFUKbz6FfeyMEqr85pWwOZLvsz+uEaDRHGDHoLu+rf6t4NKwDSKBV92hI36nFxBAbHbqhNFhz
VRGopE9FiRQgrvm/1j1uUSj7SSM1Oor4vL1xvpgM+0XwXuPeLWBPrrJQvd0HcUP6JOTK0P8eOWm1
invrnWriSE1WuMBYpTjJh0putUo9PQRc/c6iGT/ccV7wFSPZSuXVjDI1Aq7X7t/4m2fuuZ2sFLKW
Dg+kVIM9Gzw4NSs4enctqgTybQ0effmpHf3bKseQVtZ8Ydh96ADnA4mh3prR4oZT1sto+wG6Ggjr
GQmU6Es/WCNHo7B35Z5kwZZwEAkxpp19/CU3xhpDokv7q4/W9P72ghL/rtW8Z9FYKnwltQWjtM9f
LuoGR7EfEiq469yHRGboOMo6rOO3fZn8JnCCKKcJ+wNHp0M1pmqOcHxcGxTZ0d62/vPWO/eHCaC6
BNnc45X8Ho5kZ37HLS43nDrHSqHng08/VADKweMd1ib/+5OOH78QkiU3gJcg/A4cJPR1FvfeSMCM
25x7VHI7YG4/GW12SS4nnuZFL9DH/lH7LgQOJG1Hk7uZ3EW/lwh+XuzYqUmnWAL+15Er7qsKTluw
RqciH2NW3wmHVYvT/o81rGy0xCAcHbBRrLWisf1iccWSZuw/A4NGWoxu5EU5akrxPc2iNF8KPBop
wY02IsSFt3psMMQ+RiX72uCFBb/GkeWIrh4vn7EXxv8Owvzo5IEprWCiMf0L/NZdkuHNwR6tY0Fu
aH8AR3UfNXVMkQaJ9A9jtZF7BwEWV/+PtD6ozzDf/B7hdvGbe74Oekj4qH4jagsDPL3yXikFatHC
PT2tAAWZQjSd19KjZaivvxl7otM/dpw0oBAjBGPBsAHyA1hkF6bCkGr57AZI1GhgnJ/w4r/PIBxm
H/5OSHOn4WDZrho6c2M35sFpj4K94I4DwkITApVjzfrhGOAifJe7DcKowVS1+PqIwd92fVrx0yT6
fvNM8FCjMokQVr/JoeLpbyC/Wp3YuQkAHtCDFwuRy2YDLBq7XIWvk1j2NFZdgnbHojQHxnhsDTZA
9e2HTl7UDZettIy1AV4fqJMVHffVqwynXw4yYZkURCemStZOTDHxJxkcswds8ISP0VSZ8xZhkO5H
812FmDo+VjPzKdpL00AZrFFQy1jCha8lwYPk+LDt1a92cE4H7VkUo0rCWNI1jyMO102SAGS0Wry4
SwJT6OLvqnJaOgS+YPxfEnJ1mklzc/g5+URFtVl7WbgORlbjkLNARv3yE62L2jfb5fOdLnFabVJ0
+gJUOpcdVeTGvnwseD8aDRcpKu1JbU+nG/vfOoAmeJZE94g8r/rKokbd+hzxHbN6DrEEbjSCKsTD
7YhaLJP7/QSDJR2d1FF7dvMEDMd3wTtiNXZ0lpZl4Ubwlo8M2gkz45CNUttuWmgACimnVhzU0aIY
XdbxIMg4WEs1NO1E2IJVfbS3EfOnoiVWyJ9ApikkA28ie0tA8mKLXBrK4oDXH7AAMrwq4+5Bt1Nl
NQr2euwGshGCpsFu3BcfqoSbLw/8XSUDh0W0ggKSqHlQIw3XDyy5OwFYxTc6NHIWADtUOFY3g2FU
UzzySQ/rD7TYdia02YPLCj/NhsxrqLlH6RmZhCYr8DKIwLGIyVPBBMsSitJFuulAzAvmaQ2nOX9D
vJUoBtwXIZP5zfocug4wcWR6Q86FYkkSgI2CXSPaawp6lyuP7Wsy3paENkIw3oRH+hAP3tF2yzA0
fxVFWO65fcy0dnRpFKep4waeWGyzRTPZo+tbbxeZ0vRZVqKPQ0/MLALIHeysixquqrGhLRZuJmWm
yk7X3ZQYqoMxUutEhxggHMzASHSbiLIAq4bcqcWcHFKWqWdWpMJy+4JyiBz3xrFqKdu+Oa1qavxW
yTRWI4GtLgV0WW3m6GtPFI4Gdx8KyTsFSG3NbpiafftuWMTnAZun4DkCEiuTJEpDr2FuWJpHbs6T
ZrI4PzeyC0QET0Saf3znglZsNLWSPU6AFeFab09myWj1LbK5zWXubbMKyDr3X09CkIuR6DXTzjdS
SBO2mprFXa9SomXIKPirbKt2IOD6/y2olmmNMYgw76eoMi0heZwbeny51r+SELH8uv/kpQ2b8gZt
6zFDDXSPOQaRTGhXA4tJc/PsrduTmilHsABOyVDw/X9u5G9q+jVVS7p7aYyCVMAv7lVDGtlANNBz
6/tKFoJUO1v3Bnqw6CiIUIjArHoniAt+pURLfKsZ//ReAFivs2kh1SUfyrLjLbXm7yCLXXxUI5T5
Yp2mtNH1boYIuLAs7qjALY+VWKlI6eZRMLoxM+86uaWQ8pzF5XGgGGqQkL2s1zPqnKtYTIk0yOE7
ujR9ByNF1forbASktXR/XLQ7dvOesuH6CD+BmKVGKPPFnjvFoeFZTKO38PhY1tdTDZsbIAY55kjV
hDAI0VbT2Ziklp2vfPyEF1TTrcKGd+52g603nFRJYq5u2v9FssAvRwr615Zoaheon68Tey7eh0N3
8A2s9KZv/RVTczutr7Lx9uOK+jk7Gk5PoLMcSoDrnW/i4/OVyUwd0OOUb1nqBMiat0MkH2qmRJbI
NqxV+Kj7UkRfaheyyTpwjhhqnQFy88xONBYn+9+WBzk9lgvoto2D/TcfNctEWLjyBkNfZLAFdm2A
Ixt8lCg3SSZ0Z9yDhB2/PDJwCeaaXMVcVRYUcFYmZdfMWiMPTTD0Xa9L3Xi8buDpAYuZUnGFQXL8
f3Ibk1eqrzrnxYMrzcak6Q3/PxeBcQiQlAxJ4xcXq1M+bvislTi3W0pKjwGnmDTXlYk+OoBvmIRd
RfHGnCIjsjsc65PIueldL1FP9FQ7fWuHIPKCKAraLl4FUAUjBj3dyQEY53zT3YJc54/vohwzRRIy
26VVVVeR/ACKHnWc8H0Yotk4Ej7RwZDuLwqcX3rk+///mwAMe6Rkpp7BA+privof3sUX/Y8ttlPt
rfGBkGfLmHjr0buh1fshU597NOz53afdbpa6Gwh11/hDcwGwZru2GUiz77DcjHIz18oboSLXK19d
udVksv++9X0RyG1yMj7/RUrD2+gLlw1NMKZbmOlxkSdmAdLEk2vDHz52bUZeJRmocJQrOs/ODaN5
7XGJfW31OvhG1piZv+3DgtsWVANh/w030YYOELV7cv7z9/fRv6ZCATKzMRATyzF5BzEugwOmVlE2
1ezBOuQ184lZ294Tbb8t0S6rZHKT7GuETczFUKsjB5yt5RYASW39rbTNo2aSgjAoH4UosoitCJux
pdcQuvEE29Hw0QfjB0XkVlwqJk5Pp6KAojLpr9vZ6BMOkUqoD83qVdw/nDKwc6/eQG9rJ9e9kWK7
NjLLhzgoKw==
`protect end_protected

