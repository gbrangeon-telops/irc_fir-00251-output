

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
J8nZtW1Q/IGk5bZ13EIEEDntauAKqOlRji4Tz7aOFZMrRrl3qAAP4lw8839dxHbOPehATkI5mWRu
O3oQzXKv+Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PO3vY49rlamMYJ9pWAsIelQmo4roKT2hFecsbIIwc9Ce9j1Gil9MEDKbHqn/9XWL2CZb1+nggmfu
MhGokjjD0xhuA7bkrZ61EFG47AtPbrzrGJmyawEAJ1PNLVKIspuVYNxaD9rI6pyGoENRti8P0hyl
/TLRO8J/SzWO1wVCE+o=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lek8GlHbeyFgFk70bzers4fkqEzZWIlCFJLfSucq9OzFI+lvPoCv9lLJF6jbu+G/Gu5TV4ZuNXdu
mi0r5LAo17AD7VicMD+MhRKb3DE2N3pAEqyDrMS1jasKAHiVpH3eXVPN2AI+lDAVZoDhvjSuQjfy
us+5QMijcCxvAveyXwnL06kT9i9dtQ6hie8/MMqHXkiG7OYqxKm0Iia9+F6bzSI9YxeA8Doz1sM1
HWlzlbYLDBCHp8//PX7kMS2bPsw5C6UPaQ+TKox3agXXgpP4ea6EVU3GCBe7nIo37nZIVwI8YFKU
1lK2hwoX/DoWAQ9zzkBtnp8rOkj66EFG574xNw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H24CFb/lxJKnebrcZ74EB0cwdvz2M6JUcau88JBt2iuFL0aDDA6OprhhTeP6OvCciaaGRsBEok+U
cbANkg9G0zLP53/WvEkpdYtezlQI3mkakzT3UxyQr7e+pL5MFVi19R/4mD0m4WBOiVFQ4vPfnILO
XObce3WQbGcK+NGRsMw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RFnK9ETQkPWYtdMW+yKQ1MaijPhYXOMfuPVBKnsFVaRScaR6M3W3RRHlGeNOaiw0ukl3q+66K1rC
RHUWrifpwoSOSO54nuXmCv6joF0+cR+UF1LUkBtOigSpmJUx9SscdsvDcBNzrLmtogpoKRScYdGy
LrKeBNVoMEblduWARlt0XQCFRD4X03OLybCK5/hlbwAJA/OXY8QP1rB1MFXLkjS4zFm16T1j7dVB
psuynNAT4Rwsqrw26xpeXem+8Ft+gBzXVIL10rNKj0y4I07ITYInhk/p/CsNH9FgAhYM9jsWml7/
R3A8DckKe32XlGviTUqdr3zXyrsrjZFSJ1kTGQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 107936)
`protect data_block
E1Uc3ua6x9u1ECvYnV8cltlkihwUH6jslsMqPHdWs6DicvYdrWAbtbq46r/jV9z/7xo7qbBAc6EM
rQAAMlaSzJOl5cJxSsNR61XwkjfIZQc6KBcTMCjkaTE486kWvS+6L3jk7jeUHjNiryWSGCYFk7pb
ixz3UX9TGPntLHp0FpKdB84DFiXM5YgY/2iAq2VcxT4EonGyqp6KK1wuiXq2x3ZCU1vVE2fCWGnt
mapn45UTw/SJI68RsihFAjopDQmeUGXmJeyg4MAlwGKlDF+PrHiGxOrygyJ0UTTLXz2kUtqG/zLO
OrPX101MsOP6jvRiRankvYH1HiMNRM5s9gFi/rhqJuDFBNMqGiWX7aMFRxbC7WNIBGDHOYbQ1J4k
7qfP05zktaAIqREPNqoIizXm8hIbDNP/GGp8El70iAsHwVrYS2ks/YRZvz3AthyFIKEjcLtGIAwn
lJWdtm4yaPtjVIZPV781TRC2DD3i9Xy46JHXGQ/mnwcuS78kukm8CS7GxCKYPLuc75Pz+9Hx9PlK
ggt48PRbzsauIPjfusor4r8Dz2c7h2DQnnCbNwfP4qy8GuDA2E6YbYUPwx17766UgAYCzqr+Hu8L
fwLnkIt1X3VMHUV9locP5yTzELc8AjwW6GtGHqJ9H9bDJojXtaB1jxs4jJzESL9rBDc8vLJIiPuY
zp6b+dywnaC8EQzuicCfPK9iTp9O6R+lcnEDHVDr3CxEeNQKGhYeKSvKvmsVKRxJI9bpFnOIccgj
jx2i9o9REwDS5cQ7hXy53hU1ZzK/KWVuztG1yHPdcoZIZcytw4CHNimQN03DaRwUsIrtAU2HmUKn
gxMCC/dqGMdpXMbEVUE2c8qlaTkuL4qP3eUXMmiIe/Xvc7V5NGB4z0Z6CNuXOyQfbvCV+GtvMOJj
+eKupPPa8a2hNYBl8r+MHhfiNcb1IKzw9vlSJdohYkVM/IMhGolsimA24Rju20sESAnAv4J+kzS3
7buPZlt2d1iIEGC+R2KYiYH8FDIMZNKmi/CFEkl4/i5Map7AklgezV/zVlArn2S1lXUD48kR69lq
m1/Agg83cS67Lw5LsnUUMgtsCgQdmtLzkRGFcLe3O9Z4bnKD535jrW8FbGCS1Tg+EVxykXmq8Bjw
8aYiB4OpZaafsfOHpkyzsqgy4JOgu/d+6q5fcK1hZg30pzHtFuxjoerhkKlsDisTrVO6gTZTrA9n
H/0j+quOELWCKVOja7syMHtH3lG6aen7H8CuStF4duR5F5Pryj+yupbhTFgOFvhY2JBRhkyLu/fJ
cHaa18bn09g2gHmaPAYSPA0LUEfBHcWXIcXoDj6JQqGBoMG704E3qO5nuwR1VWsL7wU6LP5stz0O
FeE4DuEe5LjPh+eP1aE5LnYPmL+nWGgiF3npedcsr2BNaaQkMoYW8O4Ay8m7I38KVPSa1gqYMUam
Prqg1MqSOuHCnx6vSvOpfPTAj7SN4cCV9Y+gxHP1/A/AH45moP9vk2rIBYuiArh46i5AG6CKjwm6
VFzBlfRKgVelHy62Rd3RM95no6h6vNwpI3zsZg3vxZmnlF39GTtSI2aFIsf+hFWCQik9+E2UfB91
WhhZD3Ul9+wvi99YgkJ81U0bxZm+jot1RjmASZLCcXiDSSpvQZMyHarJ33ZnSy0uIqP/KEe6of0v
WOmqtYxFNpCJsXs5RCsIcQIwuP++21/yjcsP6vvUVHNHMvtuzxB74NR2LJvi+w+TrUv/zz7bwDGD
FtPcTvwW72/zt+C8abvgZWsspebwvhzTOqPKtZbrNYoXsRNQZFy12wFdoGY3zy3svmRPkQ56nVvx
RbLSlseYw72V3a9EvQ33yLykjg4T4xMOjM2ph36IQ2LsuSD5Ley0ElP7Vp4WBUayD/mM+v4D/fxm
OkG14faUZvWGRRM7+XuPQ6lbKt+l8Q6jgMVY++w6sWCUOCuWl7HA+4vcp7PXYA9ROk+J3aIpYUQU
Y/daDIREAcRrFsazUOnZPCCUSbjUayk1nlE0c7a0fvdzi23Zv0U09UHszn6ZF+g//B81Auv8Y+S8
e/4uBQlS+GFMtUfabGtvYmj4a3yIKC0KeDZSeIHx+3Uix99UrtEEsE2Wh5cguGgg4D/kBqwMSmHZ
JJxq+gdAYM3yy9tOXz2yRdpwv6aW1Jg6J5kCymxo+R6JK9oRlTJhy4OpWkHpZQ+CbQy1IR/aqdjR
bvyBBqfO3LmkRz5tGlXkKnnV0McnMXJAED3YCewqH1BGcCPaHN/wbtywOq2kashWPpzIzTmoAXPF
6WyxoUOmiLH84oXxWy2u+mHkvyOZY2h5/AJgKY+c2kpN1KEaObiCsRXUMKWAF4jlXEbQXIS5hQ2S
e6ZOcn3hqSu/zu3g5Wd0JI8TW/Ckv9tMmOxl95Uv9bxJV0AQiXgHNmbgK5vX2W3DL8jjf598op9K
Hp9Qy+Cyvemus2goVHBqcBPsps/ACG4mHpEP5NFpf5fzFVbfvfmkRLAQ1A1iHF0tRg81ReoV/pCn
6aiFaA9OkQ+3CJwj65PEgyQAQgjtqNbFpTrt3qtTuXvkRuQvJYrHADCwPJm9erTn3eObDmt+vPWn
gNNXH0dMAeluxwzD6MeUB44CcshRyYn/nhX0lyyqi0O3t582U2N0hZi/j9lS2AIPNcsUByouHJai
3tUnkY4ILTGVw7IYiY48eNns2zYD3ORsd9qv5HflG3bU5W8rgu3gFJtovC6IiEFjB5ek/OPE05Y6
NLxb58sjZ4J9gOuO5iQfcmHbGKDJISG1t0iRsYRTRES5GhVCIWWVr+T1q/YwYTN4ND42j4x85L6J
ddUrTgJ3VumI6DTbX4TihY9IpKG4vLgKFPzB9qf8ZMbw/5M78GtpfjL/TzkIUzHqIz7Vo+KhTk+z
RyEJJCUhRCtofC5gKg8V8yXQQBsMINHMjTY/ntgSLR35nmIeAvACDxDmhTi1zKnctZIoQj4MP9V8
7FVOuYjC752nf7B61YNMqj9OVjZq3qeVKomAfUG7wcyAcsOiuSpDQzDILZG0/lF07/6WyoDAPaXn
Wpn3gTSUwFxk1At50Bz6cRrd1yS1N+Joj0am8OLIuoQARf/wzYkU5J+zkzTuAg08Qe07wARG/+GR
BvZ4re0I56KkuwgmGnOV4qe/hnirZTlTS1tcu9qPptECXZFhffZqCgJXx46fM+KNFFvCf+pAuUHb
xDxfi3dPeEPvJHCES9RWEaRo1qmXGmUrTSn2aZS5NttzY4nNsRsH0/D2d31+hfVw+T7TvKjLyKE+
CK+jEI60hAWru9sHBEKSB7qhtJRUu8wxx/3+wrqv3yiR4YXIS26gRpbzFSlpTAyVTl6diQ4JmyHV
ZFdx8qGkofA23W1XSIvfAM2CXK0FxlyalBc7IBTxKD8jfoH4AsDL6YD2+P2LHOMgf3fPznK4ylw9
3v06q9bPB+mc17ANMKUFn+vTp87cIlTtHZ3SD7SnZjTmfdgybETqLFbMYy4mRrFpiG9JtDQiQEp+
XKHN1H2+sGie3EeTxskXgNlT23sSz/cBHjd283XzsB2MktETKituG99P9/a7/MyCnvE/xwAViS+e
Mu+KfTkd5BjrtBifGcHX+ru70zGvMlnYlMJMl/TyUt7rDwR326J4i4cuLSxGaQK8nO1wRwPwfsZE
OTaweEvHO9qmSTRpqgx66QohiB7k8T80cJ2ZCPiw7o9ly86nlIunKJlb74+SOw3YqKP1r3HZ/44I
5KT201bPpQu9aBYKVkW20JcBIq8EHc6QJEM2mGEU+5VKTNSXMA4fei3j1gSxiSMolzVpqIGpYujs
zVWIE5nprnbbbgnrQ77Xr7219OAZLeOzeHT0hrDnVEpZSf07YJ/95H88Ad/iX34vQF9+gTsokcbB
aHAm1Gz/HLbUGGCvuTZ5ljHrdHvyVu6R/ABSd81Xlj+UjQ+Z+RKUja/H+F7R2QHqc6PxJBKal1Zh
IcXWSwrZvSAz0ZO2+dRALwlPUVBYw3OJtP3v3WpMf+5cUhzdMwEt9xdTKJbw/FACaSMGvsnP5XQS
iRwczEzU7Ulns3seJLfzekhx9+dGDwglW4BUsKofRNJc/GppP6VI4U8YRZ+CePAdzpaSHNh90spU
iWLtCU1hMsEFShJ/h82ZBPYpFd7BWrCTNuCA5Vrx0ZflEE1tgTIuSVonfDF75aSpTqyrBa5tZt5e
4lmVeJMd/a+MzrBIflOzjXr8bkGX1ff8urx6mIlPYWiUX/ZGT76c5RqpEdVvUXy2TA2jgjZCW6fZ
KtPBOLtYTu9pnDWBfR+JBcOfVoNhc4jyPEu/rmKiIi5iiihmUVdUO7fnPSgXOkIK2zLiSJZM1vJ1
cZCspocSf5XJF49teHcroZMxvTY0uMVP1vhjencHJfqR0znMyMGsLPShDZQzItpE1NSz45JCTbvD
XVV1J367LSOJGkIh8IxcyxO5SZGtsw1swt4k+Ub0p/aS8VPbdC/yBSDgJ7zmnq8dkLDL2zHl+z/n
hGpvXybb89vXMS7p+/QHYgfRdj9ZO+PRpeKhR6KUc3NHQSiI6j3TdrjH4Q3PCf6E60EK0XyBr6qx
zMTpkxNbjUoYyMYls/LmE9bCAdTGzqIrNcGzEU4bK3b9kecqiokx4D6mv6ABnb/UBUr0fCtch6sm
7F9XotWoKWakzsF/CYv8076Gbga6Pm2Ovik33+Nt7OCeVTAJkqscAcw6JVHhiP4H40+2jqy30lm4
NELQ5KnQMbrQJ4OHMzxubdDxlVxsLVU9c2R1TA7d7Q7u2rEJOcBI1VJUrZmj1sQetAWl0vf0GeiK
iqb5JaqUcvxLxXDAG91WyOmB5jdciTiibSlg7joKdVH0FVpCw2HlhVCrJYWjniw1yZA24TYgf9ug
tiRLxQI9SgOHJxwl/OwyBt5JN3QMHNIVsEHIwl8OQcJb/IfFqOCDoIrBUMJlQolCJqUb5IKr5cf8
74OVXzrViUab76Hj/1QE8kX0kLPfOptXHTvxi6yPdIhCZPiEqozNvzNpFJRQa1nWdCm3Mpu+zhgc
/uMgN+4wdI+gIgOhfSS5OhU9fETeyR1m5KmzjDf+nixR5i4pp7jJGq3QDeLIU2wwFS0vgUh6nkrg
8rAW/aYwZ6mu2e1pjP3jHyqVuSBJiH+pjjY4PHia3RKT9G8i2zkM4FLYsKctnQsp0kYr/x1e/FY+
/ZER1Z+oo++jSBs+DJ6Gsr5UygZtghT2jLCr0led7f9EcybyHDbI6NCA4PqWHHjmdveQXZYSveex
9lFnAzX1dmd1XJQhpguPd9/LAZ9JFr9xeC0qa6waXC3eSmtCTXvHZbqW15EeYY7Fsz3iUq1CPCGb
wEzWESEScYwPPs2wpcaXRWpof2cX1iN6JWU0jL4On2tnWR65AOM/upo+DXNxZooZQOjMEYcvVmUe
LTGveGphA+9ON91/JXyCaRjrw/hNzrGkik3dcX5pmE1xvbJ2mhOof2/x8T0sbxUIP0EGKdbxP8t+
lec4MAIvU5ABBUDCgtuQcnWI2S94asZE6PRCHhK6VoEXxei2AFldfFssFHtprjPb5IUWuH/cT9M+
OI73Tp33Qb2Q+M4qJXQJE3nHlOUX3usJUspn45oWw0pYmOxuEgEGITStbZ7JmgGmbnwqZ2OGWHTY
//2S/EgM138mDOUZ5ZMkYEBG8VIkCDlKD3jdQjAcwE8rUtrWN0N1U8FLjqYy1vv2ruioeXr3il6/
OgvXLs1XHkBHTo+BqSvyfPKuhg92ZQvSteyN0oPPofaPqMYPzQrB9alAwzA99Hj9andzF6v8a9hH
veMS7LhP/pGElzVra1gLGBezOj47rqUbeKML6gkcPfgBGeR1ziigmmGwSqOVd3+xe9HXQwgeI/kT
lRcMNgGar+iREjeJotsZJyBFkYS145zUjSrFtHMig8xLXUdrw55MxZRsyCqRwSGb9/eLsQptfF9m
yADnxDOkffcmANZYmk6pP2uqk6mNIXfWnVEoHMbbLNftJkJUz+yH4hBBs3r5FkbsGkfLnpUJ04Nb
kyMva420IcFhz5GGixQWSVFcls7h+nDYrGtqS9UDRUDuVOeejz79AA0N7SBhBavF+Cf9jD3J856q
r9rloLfgtE9znBpwHzuuFEJ1o/11eGWoRMey/gA7nF7/YhIXNUBgJDuK7G7LCkMik6cuU+pmZH8+
WuapPUNZJ3Nrxmd43/3rTcJwMSS26DKHCZ/RwGpNXqvIzt2da4h0hsFfpgsKx1lKwHfi40tHzU0V
WQ+KAtPkB8UNfwbmaN+Oze+SaguhAlcrz3kmWt4QHiqtVFVZP/eOBdX+EXlR2DH1ejPdCPFv4SIa
chpwOMwdztIboKUE0EFs0kbh1HURwdF0fzCovY3G6NQbBZL+ykQdCgpECrVZV3hKZrIFp0j5TMK2
fVUlKRIlhicy2XtmNeUhllIGyUCwRJ1iVH/fr8d0BN9BCJECsgA65x6ntG3DLf91+1av7I6eWNY6
LKiqZjYFpR5MtIFJS4rRUzImNQ/WfoxljxzuZYfhSNLC5zWbFCucYMbfq4QmGuoZRydRew8T5/2V
WWYz+yp0qkmjGHjyCkExoF6LvvU9JpKUrwQ0XK6HO68Zrfbdog/VAlP0RoR5VWPGukSfGOZzh/ox
09mHV4gfxJvAfhKigFjN+lX6dKVxbb8kJqZYuoQScBNkho8GkxYZANom3BXpBJ61Ng8VWv7X9xLc
zZfUxoVoLijd0LkOAKxu92yHhbQRVnrVZ5huY9IUbYpMoWHWr66tmKSiPf0S+iqr7PcOzFH277GF
Y2+9OhBozqGWDqkjsCvojzYhJFmRnZlUQUesn5QNqdt3AisgR49OqRT93SDTpRijbnRdA1KFyl9g
gfa9HaIwnL7jiz0W7u03NIrWoqs1MioA2xCcDp2IN7WC3yfXqZhKOxDtD07ezBVGz/NLiWucNk2I
whbf5c/C4/umEiTWFMWDLYFbW5UIAUAJI7izxR/seccpbVWpkv1cOXSIS99QwXFFdL9po63i+2On
mHq7jg0cq3f8M5P4q1UG1N0MnBR+F08U0QDzr98wwS1I/ufOf606WNy6uucMX4sM9oXuhW69yBiG
0n/RaFGEj/iw6oBUK2JLNXsSkQ3VAph22nlWQDLLTOa0mxoxuRALcsrVi3QgRTMCLW7GdSFi9QvK
h8j8ZKaJ+CrRAPdISbUeliEiNJtLaBsokQCAl7+nbri8HBjRaJMeh9Myry/7RfGRp84py02f/dN6
NCDY2QuX3REdI0KHTCF2fn5JkZiqY2fCF1szciN6NeZBR7uqTvEjaujds1owQRtyfxccMSgc3oYn
0T4RToG0CJa+uAn5YFSQBU+KwQQX5NotbIRMqSg70KQZnh3q38VmuGeizuCrT5RQpfqUwULnS2F5
BrrSwlo1N7YANv2LUT8M1vPliMcvITjO+Ryb2FEW193BVLbavF4AERyVAt0PNrAxn8L5/ZA+lzEI
9vx7YD5yvEZgwhE6C2HUay7ZhIvl91ChFVx+W1uOALBmj2veeuCLE4LrGaQPINpuH3KE8BBo+ASl
aEjjp/03MZfo88SxRXJIUpPh4wEbo7qAgZyePNpTkILIh/nQMzziburLfRAlOhDfRhlyIH01LS+C
x33NJG+q7FJTX5wxMD7cU8vGGEhmn66I0djelc1cxoGsi7LLH2dUuGNd6vIMluXDTv6hklNnPSHe
rlSTGnJb8UKPJp5vBhMoraB6XumpeVtta3gwyWcwiWIVRkUOCgXS/2OS0RuR1KeLXBK9Qi0AMHNz
4fa0uH8CzOahmBa7gTQrTynwLVU2PbZovpwMhnIL7Ml/iR7fWAofHim6ZQC/e8QyVbxF0swXfnGK
1/eNlkKJzTGjaUykUIwoBBt0Q15xFwIIKAqlRiM0Wa8gTyO2u9/Suij1g0rq3AS43JQ28yVec7eB
8EIELQdrow2a6/eKmcgsgyihxtARiojudiA4E8ymFvG4t93sYm6hjTp53mIPsF1OWxbyjyKVuD5F
QKeJKsy5E55tQZpa9kTWuGf9gCuuVYgNp7JAM/q8GlmzKj7DuwexU2l2bp5l42HaAY5NXBLw1bUV
Ixi0l3kCyXvYwVt3m1ZSIK49di2gpC/4bYLowBaiG3PXomq8Y6czHbtnqVFFueVUCXY+CyMS/vKV
FtDpxVrPFymP1srLSloh3NItMMLXBmZzD5Peo7mq0QpHzyKmRq3XeRv6MfEnFgy2qtz8rInlFgSX
PM0+XvTpQxliT7l3+IT5+VO3n2TpDrxTHKqJjcNaXbbbGez2qR53ArraRaYBmRzhuf7NP47ZFAJ/
hQUkpuwtn0pd9wT1Am82oQKHq+ISLe73YOK2xQxR0Iz4rm2MeSGhexY+H/+ZJ9vWbhVxNLvW2wPx
QH/w5jcCDOArhiMed87L2SGbYYQbm7PAdHNn/+BgaRKCTi4gST/54pOwkOIvAK+T3XJq9OaLP3uw
0/xbISfEqETkzjIckkqhNGw7OGsAClhEffoUGgRPVJtT07aNs4fduGynI9rbdeGSLxDaodaMzaYl
Hl2tYk8XoZ8sMe+XAp9Y6Rt8F8XO5aIDC9nFeqFpOZ+l6acDyC4I5AYaAcD4fw+L7hmIOD84jw2j
IUI6i6b4KOUT2xZ0/3WEENWqRTOzUB07piGXu2xe+eUu7pPMHRgpk740peFPfrtxEFBzBCsWL4RC
q2pdrPMcYIyGR5F7ogqFpcOMQlqaoS4YxNMWF3iHtx5gX1NiVP0iudNpyXHs9TqvH/2q+adJonmZ
4odSrqwBzZs0SuA/4HyIkO0joepP3nrtXTKkw8jAHZoxDdgD0wnjBZhSaZ45DGw8nZgGcr60Opgw
RvXiMjxQcxYhL45xoYTfOG5fvYgYtPDyLYO5CX5KRQFXFLimNKiVWPh9tiExtJvOMlL3lUHWXsj4
Fw2AKXescxDstmJqoiS2+bFWvqAGDepnShl+NC8K+L9r+cepiXNXactIpF4+C3Wyd4jCPbIE9Wc7
q5LRPjBof592iUxy72IYpAQrM6BR8Ow+TqmWuNYWq+q03OEaLKl6XNq/prq6JGfkaqLZ8kEhhVQt
f79S3NoIF3/2mzEmyo0ymi0VZMLmPtuGHdlpCVHj2TMwsXE+YOH6n4F40J+cI/pBLfdUX7ShQ9lR
2/2odem4quG7coag1+U2c7j7PhPW/KMV/SjB1WkQdVY4zIF6gu5KFFTM+xM6fxHocMAbm3QVnDOp
recQZ/hYNY1mAHcXV+gsCkmSOj9nxm2bMBPTy+4So1vMGb3F5doaR+CbYwFelHDl4ABRVhcG4XZb
PNFpcb6RUTh1WFEsCqkAhQkL9Ck3sWhpUEwPRLbMC7anlQp7v83Pn3FtlVGFXkTlpgvGJmwmH2+s
oXAverWssaBK5iMoJQVjNhKW/U+ZAlR9DwYDbCugtcfUOF5rhKU95CLnYoZugy16vYx2Yy7YN8Rm
Fye2SGmNgrac7bxaJ+VYOxO16MGhSQ3YihYFjo9FfLrKoaoMvQJvBmJ2hYgaok6xC2wUkGIzc6Hf
M4ZprAPF12MArlPHUejmgWs8uUu/+1RqSKAZopZtwcfaQLdMYBZq+kl+DNUhhp9QsQ0/v4u+xQ79
RQksMaLnxcpkUkYPavu52wpHx92YM2iOSGWWwZxjQpi5J5BbGkx+HbOXAky3FmhUudGThnj/dlju
ZDms54TtiFCxGbLx0qB8coIwpI6VZ2ZLJT10LIjv+vmwofzRFYpDsmISio8rI2MQntuoAXnFlXza
0YKYnL6JnYTGpZxRNKdcOGe3lMv8bcJiVMZoaZxOH96XHQ/IkHWOKRLhR7Z+iqQlQIxW4FYcZ+un
+l19qPa5uuaMPj1DaxOEkECwjLHzheCqW9L2l7LgIVeSMlbNOwI8qeUmP4Uz1dy6HKiOn+cf+Icf
O29d2wFrzjmK038sAKxO2b5TJHoeQ3pq9yqvIUB3OR5DJlYDjGS14zG9AOJormpQYhl9yX9mIE9J
qmJLJ6HeYNx9qJUzjYlPMBDcO1wQobKp3BEKJreQ3FcnLEzkpgLocQNZNe2tATxKFKiGj2P+lCfF
dJnqHfBiDatXNWFYVyOTvtaHwEu4FFVr7HoX3AcSzs2dQRILXdNjxDFO9an8MOdbhDKtTCvlrnSe
gOYoyQhmtGloV7VRAwhbcVKGu+Ic6F1vtO3REPJS2wx9UdqI4e4bidge9mzR/LZhnsOwh1U6wXvo
yhkU9seaDhcjWHoczZJ0+/ahK5Zymg77IJWnjlHNxsyVh5ITU007P3MSy3Sxnp8f0wTXOO7109ml
sRfXamYbOkOlwEUrl90RZ6HDqcTNet04CNlJA4OyPUQdUxC71XTOpt5bbQblYCP2GriiEGhDHDDf
MiJaev7ag6wiRPq1h+i3m10o7ChneeuSwzQ92+PQOUjMMy6UK4Ce5N18qjMf+gUhpbk2Mq6S6x1h
XDFgg/2vyQNeFsOoyOztR1TKzkw7UYNUGcQwAmmckXcAyLSWbOUj+Y5H6wzPHd68wPp/nUEzLYqc
PoPBMnO++9RNXqRl8ZEMHfEg1K3e9CcFlJaERy9b4xp7cj/q1iuYAS53JNprox3mFp9RAbeJ1OR4
sAO0yjJiJFaKia17DaAEziSyl8ct926i5vl2M0+xy6aM5sT2SqArPrkfoBmHUs6UtW2c5YeD6+NF
3I4gtvt/mMBU9oZIwtDLg6GGU8NU5/7cbLXw3fQYgtX/hgIGLHLR2sAMXy1E9v/0QUuBMXCvC0QN
+EUro6RZ6UGrbiYq4gTpAA1rDsRl16B7VDPbTKkY//GI7JW3QmfSm7xGaAPaT4pbWKqA747f+gky
zc4ANxUj+cmook3oolePerbbbXG14DT+wQ2DxXPf2w2/jHfHSLBKH3/nX4rvus7YKIPYFg3qzQVQ
s+TdhzQYvjcCICFF+Hq3yAuLr9aASpeMRoilVT+mc/7JKuiNz22IypmTVi/X24ELGhpwdk9+BPms
1s/dBYqFGztESlOv2QfkC3okV5KbAO/MHm4dEYAtzqq7f446ln+sBIhN73V7KLQVLJFjDL9nJH+i
9CkQ9b2HU+rAAJTFUg6wuyt/tF+tY3FiNVM99uuFwKI8AdlzTwDYVJ/D87G18aUqYbOTkZBgwGiJ
9ZPu5JxrgmnKo55Ui5YXaKLE2UHdhBOkR2y7JFWw4rRMauN4Uj+n141Igf2AsYGxGhFI5Kvt7a5c
TNOISllhVoebADYhlG0BGp2/C6yLIf03sWVkpLDTkLxITlS1EmtNLZc1Zgkdz7ko9YHVvUi66lha
MdqUE3vOSuOD6LiTeIME486x1dZC8rQD4ULkNgVynZgsGWTCZpJ/f2212r31jsafmUVGGsu0AdQ7
dv7tX4jSBKyUP+plm7XJkKJ6ZkkIEqTEHooxlHqCjjkaK7JUP5VIiWxNAfWg/jH5vSQlzXNxfFXE
SsYfb++DyLEkkcdjRrIy8wsmtmpdVS55y/qS5h4zbEkqzxGGOa3bx4g/maIJ7CTH9cKC/+le/e+j
zGlmqJDrkWJoDoaxqutlLQnZw/Mc36yIujAGSfk/lUyBUbpl0Bj6XaLa8UMfpjygRuur6LliUA1r
fmV5jvL1/ThQAFUQTQh8EoBC0cDs/UE6IUwBIhFIx1SpM381OMyDHgIWCud8M/tkS4Xjlyx2WZUP
2uuo07nDL03GT/B6UafoN0EofOz2qlYd4zYgKwEhVs0B8zoC4RhL+yv4Mg29IwcakXNno8b0fy8c
QV1xI8TWA61pt795l9Sq2uRD4tm8lxjZLmLsS/rnumPTq7VucaE3cbt99WeR+ktK0lc2UuddVkt0
S7dJjgmtP0eR0NlVZr7r75iESVJS52kOFGb/nQxKy9wOkSkZxI3bZU1bSU4OcGDKDTG/s+1Gx2RU
DPhYb1mtnLeuZ2pO730BZUSDteZc3UL+3+lnjxbtZLOkvRMpp6pUvSrIZdcdqhwnd2iZmY8/0/BA
/cBdyJGeq7/NnYOPLBgHKqJ9CuCWHG8EwOTzGmS70a08vLRCOu29J74Jk2IFkEzmQca8dkZ1qQmR
ceytFzyndfTezTvZcHWHAkIi2B2GjxQy9dvljIpZkienWEKJrRLPxPk2Sj0tEDfAesP0eIUtwZau
AQiXENJO5tN2QFPYBHUjhEb7VoqTOi89x6Q2tnPxkxXgAleoP449Gp1jN4ZqoCHiB/sevzZUdGVf
f6Pqiq12JVG7TjGHZ9OcaD5DsuFDCk2cJuVz3eeqHMJZnpNaULUl8ubm7hjAzphfrPRiEn5f9U1g
sRjNvBk3LBXBg+vwouGmxl0b2jpUh3pK77inIX2G8deSwPVS46o9FmiBQluna+LUHG2hmpO3UGLO
SKyxtTl1Pb8B5f3UC7iYIq8MftdIlF7xAmWTM6RNOVtJXYnbr3AzG6oNg9jB3ba9WxIYejp1P6DC
6+kSxVJS6bc0LnMklMjgza/8TTw0Un3d1JBddxDjY2tDZXhkgurqMxyMqUo/+W4g3aT9ukuWonUj
iyLIvp/pBPTvZaRv9Kx83X91r/JUiJ4+u4bkHjXx7xE7HJTmfjFILkM64dNj/+9rH2MIubT9x5Ko
m0TYQOfMVgjyexg5JZ6Zt0PgFOoV8wW7WGynGhK8OHHqqDRCquH4gNEAao0hatsnuaNLU6WdlFUv
XkdOSQvaNQ5AqcjL6shrXjM5PtNaDqjqe5f1DygjJcOH+yTje7YPm+jVcrW72MkXPeOhp+mRKc0u
Vk0a/tYGyYg3SmjHkq16uXy6uHBepRd5vNL/Y9sDzZ/JpVH9Oo46985WesRcDKeIMt/Mxl551Mfc
V+wIDltHGppZxSUmQqcePBu7Oumi8rUkr+YnKYJF8JcsJAzx8apok9vqjBVsyiBdqVHGvTirR7Qd
Dw5xy9Eb9W4+qJx1MqB+HE8hGf5agUGvqAyZx79RNGUR7XEECZYS1QwN8CqLoV/hAhqQw8szWFYb
rzbzFmbHIDIsSYl8zC1UoeXm9KRk5vE+zxf/r06o5KmENl0m+kpCj+S+fblYgq19C18s337/k75W
ET8ddK2Ci26sVoUcGvLtYBdTxnVL6Hmzy5gVNNo945iqDelAm2h+Ug6WQk9Qi2UDc6kAgUXQlwGq
MQIh5F8rwG6RpDvFGcfKJyO4kulWi9KAidqLzz34jx0AMNn96JAMpKZWo2StRxW1b1S6ERgtHiAD
dIHLySyiuqUEKa4XAiHrsbCgGodZQ5JUb/tIk4q6N+RZLZf+YESQowimAmBVeu2Cj5X5/6HDJ2nm
s4wocT3v5TWFD68NfqtjVStjdv+3zOWS74ImbNLl0TK3v6xbwDN/AaCTOcnmrK6qIXBOuTCZ85P3
hwj77q5pFJ2IyxdeVjUJzm15GQfrygW9jwKPbLvIOj9IYxQzHa4QZqndQ/BiKpcvqFCqkaRrGEZo
qvva+kg4JQiMSgSnvvYtVp5E8JnKn7ay2vA6O44N++IPAdK5lceYs6aMPj6CYKs52FT90/Rwsc1N
6SLCWIlazRxSd0WIwWVQ5RZqoAWdpKFAWgSfZJBjs6JOMrSNBf9Zd5269AXXkKnKzCPbRPc3/L3l
ptmI3qVmKzb7fHRgB4Tfk2sqkbx8xECq19dbV00eKvB6tYaf2V2n+CMEKlk+L1oBMfYeyBtw68Um
gv5fRXURWLYtUzQG+zEtb865YgtisWt2CaGEAkAbmtm5iaVOFubSK9P2NfxYMljSZxUBJuse7Pdf
Df/wUUTOVkLPFUoyMUagGyrECdribMOSh81udccJIlNQ2mykRLRSEL0wYVTGL7wbzRETznGsHNck
e8Qy2zCt8KIX+sPhG9dyF3FZi/ukxXPVqhsQvUYdylKFbhty1tA/NOzncfJ41RDlmCEuWvTeCD4D
gSB6aUQhbhtJayat75bp2wFwPOCyo29pa62/jMcW4c4bRoJ0CmKrLcIcaiweb/240yJM581bQovw
gxJx5EcagLwy0Pcv6xMynDEkD5jieouEHPS7N0fZqY2yOX2exTNYie19fOaqRuQKWQMDS3ueCgHj
ie6KmceRKCGdOsRvUInWUvQRNvmylQMDHUPL16eF0oZV96FZfUoDrQ6I9wjHBL0NpKzFQ0aJ1Kbq
GbidGqPncVJP40Gja2u9feeoM6V8mPhcetT5SddNI6zyOpCPouNxYdeJf8196Q+V56SZvF1xKWOx
3vhVRVduYezWEf/iQhoi3miAEj+ADerYo/PDo5Pf86CN+8oqnvKzvHzTRhsy3ja4wfzlp7rRaeTL
qBahPqBtVqFlvEQn7g4qiPMdcwTOrxShH4AyCeoLbew5Ar2X+zzY8fnDVfW1AlGJeWkYQcaiFSJ8
PePP8/P8c8SmDB6bxoDzbm8Jjc6OtnSjrZI3mXruBOf38KuCtPLSzAk4bqpt3qpjTrLF6J+gjEDC
3vgsyiEgrrfNBpue0Fhv8xnsjWWJJ8D14UFN4G3OTNi8a7kx+sy1TNrd2djwfNpkeFdozmCmyMhY
lcniFvXRRzgKiuSVY9tY6gnoT6/q777gr6x/+p9XJyuBZ5YW4jb/kpmYFuiZE/6hgky0cbEFzLs0
EYFJH3wnduSg8j0beSMX7tvwLWCx/0E48kFLhGeR7TNG+R/++e2YBfU6gAHyJBA4DTXm7HcIhddY
9IDZGUDUnrDUzZghlaSieDTvRIo4Xni0WQyczGelR9/GHzVjIjtdzMC5O7b0+jjJiO9DpXN3OXe7
ZUm4QimfFCCCIzujjaBz/y5f3UPtrwgquFHRbK/9oyTi2RCieJYw3agAz8y5mjTmK4x96vhRd8Cg
nqOMMtUO4IJgNlIkz3Txamt+ZI0HqrqW4BthX/PyI2sLCpLfROItrAvB/gJeR/XhqmfWXLGGzmPf
wLNkxdBwq1WRaS4DV4CApA4pj8XvAh6s60CCNh+NXxmJGQu/eBRirsYyHp6vsjnhIWpwPxGcL2mV
slHSNWGAHupqRpJ/XDP+qPSX3RoGxpEzdRWNg/e5pIc/xcMBT1CG9jcSMYcPK1cJfqyIXKcXyT9e
G7GUM1tZNF1mHL/dHl/KYeBDfImNzCdWXtNwN0YxV8pdBNcRm0zaYu7eM0OhtTW5nyPz7H9dH9K8
TggnDkVaMmzC/UxY4fsUW44Ty/z94WFHuXTkMcHJE1yFV5y4P4JBUKXI3MdyvwuruKEj6yOOf9II
QMgHXSpblXrXmQE/TM29K+VjxEMco/s/3BhAYEVSIUxNDebB6lFlXEMsNHPHEsEiufY85ke2+NXx
15e94OY9ToYzAqrkuvtlv0gpRCZvWUBNvmo38JliN6B4/ER0ubZvmpG4OGJukE9PWSoCCCYUpA5T
FER8UQawGFE4mZu1/ffnClm6a0yWovFE85r+pN/epu9aK4sAafAGbXahGfQzzsFmLwh8fD7fbVaW
Rpfjww12Hd8wzpntbG3LfYukW6pIrCsropQxX0I3E77LrmlEYZkNdkgFgLjFjwGWQba+Km96/1nZ
bHs6OiyIwGTY+EhbDk4/cE8R+N6Jz1p9Q1MO2n3hG8XkfZn0lKvYpUES1U0eEoTTOIh8v/5Wklgc
upHD1qNUkma1qKj97I2taiPJda8TL8mPQs8YRB/ZmmBTslm7onRi/+zv3Uq4lwI3GNlRjFSWOP6e
v4AmZv3FMG9ndZvS7v60XpNBSZ0TFl7WRYGvf7XFUwqnB+TYkwXDTRhUscgst0Nlv76txfjom3WH
4pFTp9uJwz7cRW7Iimr9P60JPJ+8D+Ka3MIVEPwqk/SN6SNw0dy59M8UAAvKqv3lEUh88YsHzUR7
c4LY+QGyapW9AoGxBKlum9CiQgZt6ansh4vIDC7YA8ieru5PUm7RRoeBs8W/WrC74zk8RnKM+k1b
fyW+NWzT2TEBx77SIJN+WrMdBUtp5+7QLK4wWFmMLir0Tc0I6MfK3lri/XaH5oYhf6siemWkESlg
qtSYXckqmaYjMaIzJp/6FH+pjgf0fwv+UDVGJ7NLA5lP3T0HifLHQT8XAlOtCfZUX04YKfbQtk9k
F+o8OBWhkgKZJO4NLAXVolu1H+ssMVEe9xO/UvqtkUQhlm/cQIL1whE9MxN3XJGrmiuT/FaiMCXp
PxZnnjNCR246EBkUdH7FjGK4sOdHyUXxs0/v7PbvI7z7fhU61K2QRJB+UaJkHlvUpkUftVbPPEab
dUco6lPhHgpZzrgZZVwsr5MfOi138tLJxkUG5udMUqZRBmPahB1vpOrkVQaLAKdGp1RTH0sKl6DZ
qCSnekwCH90lPEgKN/MOGDY/nK7yjNax7gxHC58H6fNa8jVIHjfEP/aDVpV9orNtTN1TXR4PTIKw
0h59dMA9Jc+bj1WRm04Pdz63GECi4HE9/B/gFC+Xrp2T3uaJ/2X+ABnriYF1HxEQYZV/vOCaP/q4
lznzTkf0HCTEebyQFCmpIMq5JEDDomgd2a04tt4IMVdEnqFluXNWCIEmXN1nCxeVQz9neJZJdXpK
LFIATZNSbMHDLsn/UVEiRaKm7F2fre9H8RS4LaUeGlD49aKiL7NzJu72f+H7U54tRdLHQcrdTccM
TOa4H3LLvgURpXO9cjDp05KXKUb3T60KXwzX8Svx2VECtD2NcqJJ0uyIdsCj3BjCA1q5inINQUDN
40RGfcX+U2ON7BiNNj3BUiBjyTxSIrvyQ5G1njIOmy6s88ujBgFumvUTzcz7ANN9e7EEPMqMMYBN
wUJ4k5pru8Z4DVc3fSHOIICkYv8AkwwkhUAecaRc5zbEveKxVahJ9RLjn3poOTM+VVmKE+6ioK0c
wh+tuMrPUTOBvlGemSfXkKbd8qbBZHD29EFhJLwsQB1P1tII5ogshTyO0D43zc90ubVybzNDftf2
dMSIj7OMVZ9OU33gn6275vEU0miNKWhuUyps6E6rh51VUHjHT0xoL1DUpbbcF9ljQ5o4fTQWUBIN
hSEYNs4qc90h3YUNUXrOGgSWLe1WTi2Kza56tQBoSyqRTqG415GWOdvflopLjiJb4wlAqnglhGyR
BuTn3qnJJv3Y81zKAUnBYGLD8Kr32qrMG9v4lqDuE+mZW240wAVOWBPimJLsbdHdP4VjyUjJoun6
3OQJ+LUsjAmrBMIC0HM5YdaJAmsgKPdGl2IH7NYJCZ6t23O5Bzr/1DhXSAPw71QmXSt4XGDlSmVA
ZwUABLNPhfqU17zLcm2xaid/voKFi3JaCzWobx1YWigTaVNn9A7/hXCTMTHZ9R2vPNKm5GOkW+Bh
vygkj1unDniCXFq5PXtEs6RP8iIOzeHc89FraUm9Lo/3r3M2Ym3Z7Glf7EupgLy2lryf457t5GnS
Dib4olfW2B4Ua1TRfW+2iKMEXOqMAEcV9Tb6IiUgIm5ue52V1l2R13KTY0iSR/aGaUNyeNvWutcI
pRym1jXFtHCep+b/0OcEMM/T1Z/ocG3mlazEt0k+KX2yknRakiQLpgFBKUe2VhcBMDVJPD7bBoKm
kzYA4sg85O4RzdQafoaJNpaFO6XqBw6gmtgq5+D5LXVmvogKJNAHfmlX6CO1t7FZdKKj8ssxlxvK
t5ibLFrbMRfu5k5FD8DbtbDyQE0NvegkaUL+x4V5u0p2Rh5Xv0aHB9h76CyYr8MY3AFRZeTL00ed
PTA4jRHSsnlgoFrM1nkJu2FQg+wKUzxTspvD5Fewdn+rrGFDjctFqsIf6UDjmy7sOeaMJyo4wByy
7WaiCd6/G3GvQkWdps3ZQqPM5dV0pApjP1J+BJRTTl09FqoPyNV3rPAH8wGR5zniv4rYwIyJecDQ
+uPPC6NqoLzmvIVps9Hp0oKOqyogWl3cFtOxhHheCByaMgh87mz1wBLPLEKbRhaudgpob1GWioFq
ICx3HXPUIc2aymKwJEimdXKLEMPz4bEhX4URPtrFnCCFrR62b40HvuU2XXmXqaSPOcoP/G4FHcgn
uSQm/WUkycMAI+WyH7mVA/yHxv+seXTZrVX3VuOTF7vaP1F4jA2qP5DKGXsQLEpbRn4UT40DZ2gT
QAIHiwRyNYU9Qdr6VXIbOvXltxcH4jG+sGoA+iuUXQ5sgRdbvCI35NV/5KFNat/ALpONR30zOvGL
5sQHTt0fXtxPnDkiqNsUmCYNcskBjcVV61qnLlQy/5tpVnivIygu8a09p56+luEY6gD8JkgrqylO
y95XZff/aks9/B3mDHEsw/MAuJ7YqeLlL+2txAG0gZVLPYylg4qb8Ywqyr9Kp8CYMexDbwPPaexG
5zElGZkY9zxPVlTcOK/x7l4f4uBHReTihybFM1f/dIRi9Jm1LB356KscvYVy1uQMwcApyFO3QzvN
LpOTsCOOFXr0lksY8l2bvBR2DBL945liyisdfWoLJ+5PrK3BupkiJW1f5uKKuRkumDOJsZMx8jip
B+6Ta88AaMyQrrZX7zgkA/ra5dGC35bSoVcEqT4nqTbBcf9UT8urtslP7q0JjR4thYpXPF6JMyE3
pw/J39PaxRf+wyYERPCORP0qOp7SQmJTU7RpmIhvYnuOmhGowMjhGWugHUaE6syQTuwsRkspdjNz
WX/yv1P5oNEsWUj5DPBaQdE9S/t0yLN1uUHlIppiTTki1iFFB6vFWpsPWFVCXGSdWjZjgpxXm8dD
B3nnefFYx+s4CKdCAY/DpZ2W0nsNfE0imLnEeEuroaRZSV/zPNnMuuELLJ2BskYfTVyZI7jXiJWX
2SqTuZOAuzq1B6uJsBYFd/Zo+WHueNmew9pXyss7ykxHteEhT+r840E9qxA392T5wrJAgpZEgXDG
C9BOIvA9QvgfphGEvkTJr8tCS3/IENfumFUu5r67Clfb0jlW8cYK5WGRzA//w2Qux7lIhIssoynx
oeOf1s9SC4e8Jqdcnp07icOEr05ToalybveFCRhEiHSC5wi566Za4lc7JDBfkxnEs6KkUNuxsXuB
u6a2INbOAu9p9mxMB9Mi+7HknEhoGmBPiHhg2eGYPVS1Zj+ga/ZHOWV5i8E2ZC3dD8ZM/8y7dwK0
nhp6hIbmMAPPTYK505PqZkGFwU/0SVEcfoNSM5TKH+vbX7x8Xg2VJgv1g6te44r9+oNE62sQHH11
6KNc1es7YDofT/9LALzSBdSb5wTHBC4lGJuz6nvYOv8TYlOYt31q1AwbX4rVE+MbX7yOJczYR6XE
6fyCs7ltEv9oFK9vi9CFcHMDmKuq3b5kpvXOtQWWbJL1WV8cbHIONnzstnCMFODXAfHs+UMPQr0o
LzKIETGjzI8YgGBqoD3IyC62dF0CtoMozZ15CYfX2YAcA46aJ6Ug67PxBcFQb5xd6ANghfOh5WSt
YXzAAkH1X6x6eV5mPtcT8n8M8wbP9NMn8hUAzIgb/09ncue+Ocl5SOBE49tqgfTg0gPh3Ne4rJcS
9oCWW3Cqo2gIhBKwGt+75sr4uNqqLdDekTaJO2m+zGdb7v2c+lD/WRIeu425sORISozMuVctWFqf
K4p4DQxA/UsriD20mLRc+pphQca+4mrYpPtNYwzDu2NXFT2IluRKP+61JCxf2nfX1swRj+x7i1W9
zMnzSA5F9yttpiy1qbTmJqJJakpr0HXUb/3akAmzSrnzWu9ZlUaKAAEzgMvFls/v3di6mFqmD+nh
ceTcLMod+J1+JfzOnHkq7HRrSlYPbzO+ajV5Luxxw16Def/m+RRtxkq2UZYVmQRRJpwj2nxRd+g7
Ae6mnY6Nwb1TmoSmHtMLu1jYvcq99B/YIQCc8k70YWExErCmfF9yRwo1WUN4GWLbh/SnMOcyW+gr
kUsLFV2hNFY1RGwB39U0NIesG7bok77AHehigsph7C/x1ydA43FuA6wqWdM3xdLmKVTsR5xGGHVP
uZbyEwX7OmlZX5ADaDZUv0lJWl9ziNk9hlsAzww6KUQtdzcGycWh/d+Q7UTnGOSZJHbYq8vfnCyz
vBpwG0I5jJhow0EJ30UKEwyeEuH59Da8m7yoLVOYzqJ+BW/JIxhasaCdEfgOtGUAoXblGOEa/+P/
jGXr1y4AvS9xZRG+C30idcMjoTXf0cXUHi8T9/A11oMXjcYmaTWuuvQ2UJp4Fkea4GhoS7/N5x1K
CBf22K9ENOGTeqf6fyz6xXTF/m/UWSuEbnoNU/LSR4mX9L3xyGxGfRLOTenZcU5CRdi2KECavFaO
gDDTwAA/zpJ4C8VjA+tPTZMZuij1NUViqjnx9qLeA2piruJaWsqVew5wTwX/BJtwpKbbxlImxmZw
LNS9x0Xl5fAMfpgTlkPmrgLltYt5cU5U+td6L1aKospqQg2fsP+zlLzlspAGJdmxDc6k+QIFqVUk
7IjMVxTkRhX8W/KtjZISirhD5dBL0xclIiIEkG9UKRDxi65IPwoUts1/BIRk8sbeaxJMV1QAWKc4
Q6SWNA3tB13wNhaXoBHZxYrDheLvfyjR2V0mFF6krNoBAqnYwSn3jqR/LVg9Qus9NTFBO8EixIlh
NvWrN3wrG4/VG8iogyQ8ToiYJomyghQYxqG9Jop+OgLpTE6lFi8iY5TAEr/ZTClS+PL49JG1+EHT
xMrUZLgyYy1Jnb0fuJ4Ci5ZnuguAN9TKImw7rNxWQjVXF8+fincr3NvMbRqfNVZNFhsQN39CxOv/
aKOkAuFDoRv/aomHCRRBCs03uwZHI4Ze7ki/GjuYxdy5AAyvqGjanmpjU22yAdSh0Oj+e01tMZPL
BdbD/AAYVHdirZDlRx6dt5H0edmO758rrim+gOYX1vtck4elz6QUPDbo1EtHil2IQHkWByQYe82r
7LPiIQAvcXMg0uNFRggbLOjuChynIY7hZwiDxoBCFsxJWYa/EPWhXcWzoMYtpLjEn6NXK7fZgo9j
7sedjULL08okxz0F1lLrMxSvVIJK7BTDszC8P7MjCu0qnY60XJnJkAO500X3yFs2t62pOcv7ekRu
q4n7U8ehcH7smGEys3E7Z9Ar62MUqWG5FcUTR18HGFw0m2RAbv8Y6u2pyDbVfUNS+OjJKFriZZjH
tVFfGReOVxQTMUxorvFeJbilo0ANWCKnlFofeO7r4hWQ+XiEjZaQ8BUo1KhqKOrYcj/XAtL5hHfh
Ldnk76t1eTC0znTv9/A3yy6Qlt14/2CDF6qkNmzzfetZ8+WxpwruionLDCjQwa41dJQnG8LVjcAb
tnl5r9FlPwSwgClz8s8mnyDLb2t3T29WRh+yK3keCDnqzsD1PZ8aokSDlzzjVYoiJfQQEBopG2e3
li2LMD/tkTwLdo0aPFcmhgTn5oKUqTjlomp7fNdhsqXwJfYjhp5I8nwcCOSJ9/m/EV7wBi8SNmIk
mUTi2zmLoF6MCdXMMIqtrgtDUE47FAkC3Ufy/G63EeCQ+xLg/RGDlHXwTkJt3B4bi3MzeefUfw0v
EZDfICpKrdjO42dRoJIlZatLyzgq6Oi0HqMjDoJ6ts2baYFj3mD2VDgH7L9VSKXlN+u60FPXWfcM
oKztXVWus/Mi9uzclZXpx3gQysysc3KeR2g86P7zlj9M4ul4LzWOKd59f7CrdHtss6sxx8SqC7s/
bxU7Bn4o1hqnsw+A9kA7KCW4wsu4CxWQvwgaDYAiN5ZpGFqDMjURSCIiRGM9FvPU7QdO5VaUZJyq
tKSHVLiGoh0BbOkApkaZkHfxaqLe46MGLFMdkezN36JuNxk8vNRgs5mvRngok4xqlV9suWInT4Q7
/tz3AaqofeGZYn2n+0QZvSwWAPhU3xLen6vKQyO/ux18GylW1EcOe5yeVLvb5KoH5kUuFelxT1VC
FoAHvMK9PPLelOm3rQswrdY1p8ShHURBzikVIrCf3Tb8W9JN5NfGhReodfhYUSW4/YAuuHtBv2NH
oQJOfzfh6uUbKpluce8haRYcQIozvbmD1XpGtd5F2+n/xcldEl5kbx+1UM5nhpdOTECY+LsDSfP2
ey9OU+nzHeg+ejpTWJvH5FDv/1HbbL6++k4TVqn8tKVY57+RPvVxabt9rmKK6FaSx8s0u1UWZ24L
8lbuDI/BZZI1UCGsZ9Gm5HAgxDQi82BKn6bzCaRbrMqDa/WKzjjTXaUSjBxf133hAQrszUz6UujB
h5HJ7ZWECOjJQsDWta51oeT7k9Zf6kyuHrvCG9Xsm6ZrGZzAnfX29JA/Uc4D2c95ru978DQ9NfLC
oajxjGKGmkrtUzbdFdhLTwUFJxlVqnLY/UipGxgUapsmVbGmL491U8xerex//5JzNRODtdr/m2R1
c5o3sJzZtiMgofFHfYeGtwbP5cHYTuYVfWhz1l6MVsM/u8iupD1JQny1Iu+LwrNsA+gPc+c7efeh
eHZ69VvcbKiCcr1guSF75F8yjlAyJdhIEEc/saxI8d8JKfXpGn4hNBlUEMVJsMXfabhZBqdxAG3+
8gJbkymvLJEsBvUKLhDVSTdaQxZI/BK6eG1/WhusqnSWIl/t7+aIRPnAKtEjYzkta49tGNugYI2Z
1zNsLkP7v1yIobDsPsOfgbeJ/kMBr00dvQcN0IvjMf24XhhvJHurs5GvLCTBdVZbp1BctttsGVDj
lx+Ot9xM8SZVrqh0SQzavNdOPpQnB66MvD5upV/11dWU+acEtqz6AjDbB/d/kv7y0+wi/EXaO/GX
UjsohJ2R72i1q4A/0+3NC4H561fGJffuif0GSmO89pSIytT8uCpUKRHZZIXy5yOzFKHTbMdc6KJX
CS1We1S0snm+RWUUBr4AYEq2Napbuqy11vuoY8OBzhv+a3jYW53ulnhCPcKNiZnuez8ChM7Bhhis
eA9PTa+G4tF7FCFkIuLzec7jBT7gk5ze8D01beei3+JNxfqaGxCkXWmpf3UkAdd5RZMMGXbX0Fpl
+lfn1WroXfmuOYvNqpAlJ+DuUbxTyPO2S41Aqpqyjw7Z7I/aTgtZZ1rDLVWrIcQZ3XHqaAkdqNaF
h+iPsFwWiX8ud41wBUD7w9KobM+BtitLYp6whaWSkP1hT0+3cObbqBBsGPZ9qiO0ibnK/OSDe/je
GiBUtYHGX0g+PfePgzaKbiWEHjVBEflwHQjqnscXg/KZZ15wgO+On98IiqF7SBtdkvfUbjxRtdYQ
fPQUYHED8ZnTLuh4/EJAzP3tYEMpsikgpRMZOd/q1YVOTx/Vq9K7+4aJ91T7SqaPDaCfeps521cb
zrQQx5tYKJYvwdc1yuO48Bq62WAIAzZb9ihoe9S7toWQjyVyHmS4og14UDOUlI7ORZdUGcBoevN7
ZOKILVgnyKcHTyjBNT3Icn1VenO9jiuePGwtvGxfXjs4SfkOQ4bI5HINRfn8ndkq6njlRw8mtrrh
Q07bWCWnowKqZEnVA3s/6gJrZ3BARhJTVuz91QHtdp5SVkG0SdBnmrTsPRdliUSqx9qXPnka808g
k1AbJ8tlp+vjqdbYB4/MExnhNDxB9w782QRrfpGR2sFKZlDg2laHyH+QAAlQYIxSkLYIxRGXv5zy
vFMLbDfpWFsFlGsNMxO1hXyqxyZGDRHawF6+ATF/2WVzzQJwJlO6vjdAYn/kTNX4mvznF0/XUFyh
nCJ3qj912QkHtjKG5IPG1K7T2dpNWYqpPObw5RdXGWv3pPct/luu48RDvEuW1LuUY8Uv6TvNbKpz
qfBfLbNTnRDzqIr0xuqLaNzOjwW3NXURTuI5lCpzieTsTp3FylAkAh7xmCWsx8u0JpwpPkh7bkDD
pfWeMU7GxqBkok8YoRrsaX1yYZeIJW6ZTB9WBKuIHqWhiMG2B5aLu/5C4/KVRXmk34C4UYv9lvly
btxPhYaw6tND6z8bqbVv+rEWYBzbfaseslFz5kkVyukTj/h7I63uPLyN0PM2gVZmEHks3NldACr+
3TQBLTcUgdyj4TdZu4xrm4V+HI8OlCJl/hik2TNM4fgKKYHNwhEs4jpeHCruypY393WmaZvAdmUU
1b+kfyEUIAbk3gEKGWZxrFEg5H6twSDTtow+BvidWbqNz/tWAIX8DUPxfUx2Ri7pjAPgq4lcUpS1
7I/IbQmjsXdjK7eJnYocdJ7QolD3uAZDruvb/Cg265pV8WqNJGHjulcP4ENi62o8ZSOQkScVSfU7
9EJ24eZbBuM/9LGN7DKrnLRqDqlHD6FCOvsdBrYqQ7G8Tl5jhbbfqOtAAkl+YGOL8CIvfn7z7QUG
AZaeGL7/zNtDdl+3XcXHgxPtBA5GWLkdq6gnPpLSseJO/3Dsl3xLmMV6JhdU2kcy9ucMyIdAgY+D
Xfqmtl5wviBr7zNf95fWJQxP3uNY0t/E2EppQjJ2e6fgtK8D8i2LnyUVllhRDaGp+f4LIq/bOGWZ
qLgQhnuwmG4AHEetx8/N/YdQFOlxTNgzUwl4kLwlwhaZEKtQq6JRq3KNNqJ+hCrvTLo1ifkWS3+2
0pn5y4D7nLCdHFL65JAMf/1spfwv0ZB3bjiWytEJAE8Q6iuqzzpoR084m6S7jAUSR6v4LW+oC4DV
ODG91dT/7vu/TLnTdSCZV1msUofSo2hQyOFlFqAq++Iw2F2zWEYFWxDDX7NUEIdJxdvP+evIusyh
dB9eMVWnpkqmttNEkKmkeS9czLs9nVCYbGss8cNXwtdvxAayRrpJ0IxoYOl4n8xAbqqEVtW9+hYa
HvVbzO/5BrPrCPU5j4gbsoCYCw5j6XJVaRrP4x7VmWru52L9D5Zx9MXJ5ba7PBpPtyoWsj3fSIzJ
qnEbU1Xv+DLCPJXTImRlPxM3hjkDxbQjiKnzLX1Ou9Q8pWwHva29jExAaXZJ85qqzbcGTtC1IO2U
uhDxV2U9XwfW89RgZIBgVJ31JOQ1lbjFeuUrSgXmE/05k4KUTg+ByZUCYYyNOgWkkon9QYP34Npe
RYrJd106NCNzQk8pO6n0TKdWLLchYmmj3ouwD9UZXJnmomzYXuWMvhsEsr+duDCzr3SOFTTA+fvP
n/Gufexf+8cDlgdfMQ1O+kuMV76eme/XfSDyuT1WipXGwJcW5l9hTaOIM5Gw84RJ7txRRqrXLkX2
RCIcxQbp7NXJIdzTEjeJns+e/+1xOOenPXmsSdabs+A+k68bSLa0usLed2W0/PJm85ltpER8zVk5
G6GHIN2EsLgkNrquDIyR7j3L5HaHvgXTmQKBFhPczTJjssMLWmCvQL0lsYZKh/z2QXvnQV3GDFEM
yeG5QlI9GPDZmet2ij0WezZio22ZlFRlSENx5nXUTcZ+muEfSulnrpaDsJHOtdx5laCHv3UTCO5t
wT7jRU1EJdzGKhhSYMnWMCPFHCcqU0ICpiFXiGaJjgTH2ZVckBqBVqzZ4aeBPit11Sdw0BWGOxmF
aes9xDoZA+7Dc2F98NTa/m0/2/bneIcU/w6brxaSwhPpygLLPtNK2B+ouH4I23Cdxr21FoHiIb5l
8bczxH1vXIw9WfwRKScOBI4Nf4vaJqo5spFlM8+7A2MR4PHaCF97GGU5TYdj1w1RZDbOI1r3CM69
2th3PZVVW70W2/LeXgETgAz4BzC5l+7ZDOxUwLQW4ZU5tVTcHgHBRNGeL7UGMKJmO8K9O/iahf7O
7eQdYFEogLdBu/2GZ1eBsMfbI6Ugnu9E7P+q+OBcjzUoBpF2QG3UzVQUb2aL08lagzgZncLHMqhq
qhcNoWHZu3JSa3N5Sbt5URH0HrVwPwU0iQRFEEOeF1EMNBTL4elmsxrAhkdKAMqKLwNOr/eZk5Pd
3k3TN1PHzn0P8ypVz3p8GaMPHxJCbnoOtsHcDA6vWXIzoqTulwXfNHNA4Bd2HGO8jTmyxJbRUowl
Vt7Dw4UAGYRdKujQPcSapkeuM340m/0JdrOVgx1y9rCfWMY2TpnTVP3216/rHS2rij4Ig35QRVek
AAWHjXukm5gRyvQHWQGMDgCuyjpqY9YAEoGWK95CSqhIWJoT0MVJ+V6LGKWaxCONXC7gJUKpO8ZW
MOAMDRZcRZp8U5tUkLTI//WbIHnmhlJ2oc/Pj6x0oqFBfePdp8I0ZHNbib0Iz3XMpEyectoxgvnU
XzgeeoM1P7YupyvoZvocDxaqOrWQNcz3pKh7vdcDza+1osXhwXoSkNpARK7H1ymn5CYnpWxjVPvR
pi9+mJw0xpRB/BYUSWzHa4vuRl4KXffGHh1NP2tMDv6KVVXyrmTd4e1zqPDUOXRt8rhpCygHsuyX
BteTvxGKRJR3/SI9i9YgaELmhdI+P0+DpDC6rKLfpr2S1Kq9FX3JZPsgs7uR+SEgHXgIMKp9sOwJ
nqKmhpd9YJs9kPICi4fSJYABmaNdlTW0I69hCpWOguJr9RMnCZh4WV2PyCkvP5FoV0234PxrTpxM
5o6iFqku5wYlnHtBjopNdKjd4pa7vooOee9twdypYJ9RxmMWjSRo+y3+Y7xVh6+9+DD+wNpHVLVD
4JibURx/ANKrR6YVmyRC9W3haUH5HfZBocfStiR9HJ1o0rr8tOaRkTfw58XRvLHpFYcsBkPqygVy
FSzUwdGXnEVxvpnIVYfjL4z7+JgaSkhhPgjYh75QCiH63++Lfg/OEsIaIFR8pOuXqWxaIhIad9aG
B7V/NMYobuEfW/WSsLeYANdG1qd3llGDjUFBK1N4zxxjFYymDYXxakxccvFQLQRAlCv+bnxyeSeW
BDob2lVpKfQln6iFJ6XgTSmDMtK5rzXNaIy/JGOjE6jDk1vjYa1v1On7F3G8v0NI2PBXG7jyWtYg
pwNGFvOPOZTKPGBhseptaqrHWTsOrZEBozsFuN2oGkXp/QB78g1kKbZ9cS6epS/ASBxz855WwMZ3
Oi37HdyXHk1dzkKfIB6W33XsN1hk4mXfOS+lvYm6oO9W3y4rWcZCOkHloJt9PVqFhNUwYSoCR5Fj
UwOcLU0bl414DELLHYzjgly0xMLb50LEmLHwZvhTQIUIOsaU8R04Mu65ni6AuTidImwZYML8NosN
qRO1pGhQPi+pMhrE/zf/4jhHTN5itXPlQGQQWWXR2l8ZqDphPoJdsNh6brplaFIIo4p73sR3rG9T
3hfD67XdP+33EyoLtKWxq44gWStGpbWRz/MHfXcm7/QNCPENsl6oXvhWA8y7yZ33iv7PQP35qbGM
VxXXT4FcLmZRytLMdB2fDWOn/+0ZBdppT/QG8F/4/XuobMNY2t+p+3LoE0JuhBIRANV0Q5c39ymr
Wi1JQJxzb2DuOpF+0PtW7D/73Z3Bya13BohPg2Zn1W1wKzE4rpcLWWXEyD6D4SCsMJhw7ON94DoC
TnaPKRdd3b3YeW3wcZ+mbQO9yh2HBLGqD0BqHiCfWDYNGek+r+svLx2Eedr3C5HvRf6+5CFVYetf
o9dkXYWa+RTXI5dwsPrRXoh+/1gTPz5iwtjZ62iCDEJLQIPK1ApBI9B5x/FpAYdvJJDW4TC3Z0iz
IiRBREeN77mpDBGov1SzyxxaxLkwygAQ2bh52n5KEeIwmBsfswbq/j86LJGipot13U5E8+r6VfTL
cC95CfCW+W5D03pARwyLoNj9VBDrqZ5rmqqrIK6sLTtitnn8yCL1STs6p6wyO8SXK35jGygHBjag
R9lwC41lZhPAIKgrybHNhYGs3Gz5RnDK/THB6kpj+7niDbj8QrhKImDLG0EPeS//PFmeQsfHRDf2
mrqZR2CEqmxON6rLlU20Smn3A5yQ919eRzY5NOmTDT1PzRr+11qUJQi4C3ogO0EWaByA3sA8fXMM
ILwOJhDsgRRMKtOrnOyBxB3EFy8Sm+cSgQ1UN1WaXPDSo716fs1gl+xPb/a7nwUzPEC7psKJf6Ft
IqUTbAKmy0BkcLHINz6iJkaMLP+q6xLAPlqLl1VEuVxBIComj0953OoSbBqj3b/SaWvspFUIgt6P
liwH3dtm3TCTpO71LDgBRtoKb/wc8OymSDYcf3Dxy9qR1pzjaApsxK93Jnb82dNgBhyAmRQfukqK
RUhzc6vifPgQwaKeCjXc60OJ4Pw/xdE1AcJk5Wt+O21MEqlt9ACKGG3cbxvXACkdIJIn5bgEulmD
y3ksQ5Tuh/cGbBeA1S2nx/TxupGAWPW4zlb1D9icCqympSWA18JYzqXbZd6yOG8o10ikS8pODoXY
3PUc6VgSX5gaOJPXg2NWNy55hhVJFr3QcQjtWL/MT0+B+84Mn/VeEhtVxoleoed6wJwhuc+7645l
zlgVJPqbwK5rPO6Hyo40JRORnD1ifJAaSWSvWezXjyAWVZsMjwYjxVhGwojStG1Tg6RFKtpncK4e
X+IIdMSpcDG+YYoQe1pP3HmTGKw5znTNvtzFS9Ew79rOUkCXvb+Pg58/oVs3Ch4TCzIrook+i9WO
UMCrgYgquzuqGh6OfUrzdyBQtI0geW4bGNK0jF9zRh910Xe5KX4q6Zia6CPmrpu3plt9pP+/dqyE
i1j0XBPqVjgaYUkWmsZox/jy95SYFt/lzihJfNSl5q9rFG9+Ub1UztgpDMlyGg4fh+LWwcNINQzL
pDQDM5gCLfGEJmLdkK2nOTEocoPCBKloupgJ6bYS8kC3Vl+u5fL3NXgY5zqPTRbWHwI+P0NqOIQB
P4Jw1w+Ji58SaEmapsJkiIKcJ/W8bci1hCIQMbICmyNf1ENGo5KNRVuCj/57DN0D/WJHK/ICO2oY
YqW99fQWxPqmuXPoV8YbiWtuxOr7CSLeEAzZ55Y2V9WImeBZkfV2du5jCk7TCGWb4IUiUtMp9lwR
vgPTReFITqI3PWd3PmmgPADtXDWMlfvuwLgBHQkVC5faE0Z3PPLNo43kUXfrNf0M29iDlaT2i1T6
1zvrtbmOu/57RXjJ3l9wUBBbp9huTCBOfJ6iHi548Egn1ww4fvuwq+N/dnOQJxKdMGaLL0SWc32C
B4A63+Oxjr5MfUWGTlZdLNj4F5eqBXBSb4e07rqt6Nz/r7ScfRgeAtdaQkNy44ViV3Z7OaOYcQT2
j33D5QNOSgttio+zSYO34eTfljSD4sD2AXMBkE5rYvGbLmmnBr4QURENb6tJjATvtgsNF01cozZv
GTFRw/DG0+nteUEglp1ycH9frEDqJhKi6YHxMqoJvkXvdjKV34TFLGbt6RyuFj00iHfSaT96lM+v
GZ6e3n0UEMsPjUWPIalcFgtfK+KHaYPsa8yWVmd+H67LRUsX2h3jLzpnwgUVuHCASbqEMwYZF7do
dnYNg9BV33UOMTuvjC87YdgY8tGkZZn3Osak9DbjAScms4olurkH0M0M7aoGbrBucVTn4LDXdf5Q
q9MQ9t+Al4EVPHcP3eQoMfk/LP8u9ZWqq5UfAxCgRyEvuAv+ZumRtcCQvhSqs7QX5FDSBgc2aIeJ
7fTOMniSJeThOGWtmpSrvqd8qEicHC8nuONyeWs/rsBn4auj2Ii8lO1tKtoS7VjvMvkeoExavYG/
NLRTqTcLIUp/YF+j2FyB8wCBlyLV69FVvnimFkx7g+cnE1KcXXQnslBCmJblQSC+BXZ1fAXuoK8s
fsIMLRgX9sY86XcVTm+dPlLw7c8YGLh6E3/jjn583llBEIUuDjEvDNVK0BuwbuWn6K+6gEjpzvgX
BINBXrDhQOlk1fCz0XLHszyl5fHU2p7+E8JqXaeSme3GoYw1+P/inVPfsVlrb8U5Rd4XkU9MWFpj
rv2U8kalPQxICdTanCYfQWJG3vjI/8yebXdqF8wWEsEk9ZIO+kSpt8GrNTaYEre5ycjOwgBS7piY
6H90tPZgJ528FreenGo+9dRde5GBOc5Anssb4VtuoukRFJjbAlpCW6m8G0OQEMPdqHJtnv29k7NU
6Wy6Co/E4ro9wriyIghQScZhShJc2ADZ805BOzhxiZmof/TPzTDMrljaL5VTUzzQIxLyqIRp5LBg
K8hTOGJAZgjrXkLamUkN6Msa4TJPckP83eEq9Qu19kc8SPzPaYzfIeimyd8+qC7z9wnboBOZE+pS
j0V74S+1PBu7uJnL0+78gwhN06Z7PMtRPGRteWhwogecuZm51s+DBSznOBr1UCMq8Ldz3aiCMirz
bqf448ezQ/2HhgFy8Vm+KWujNF3r+IpiacQxADLOHstvuF+ycPt1nUo9Uz8d90U4ureex0Mb1Z2F
1lgfpbKgLu5Wx7Ko3bC3R1f920/juQo54CUooEvmKiQU+UsnKWUn9AmpV2rAhp+Ih9hhDG3FdpWU
pcNPJY/t2QXpFdrOE9c2hmplTCS+7CIZrfsXDOmIGJ/aHpT+q9s9L+vBqYvr0+kGmHdJcKUC8CUt
Pv1ZOhp+jhaKDgPqClx+wLj3B+3N9b20MZ8F+vfs8kk+fEWa8wO96k3M62iZr09vuuSlMpKy6ZLh
AR2UwV1awNaJOQvyDgzvDYp38ZvaZsr56msszxfy3Bg2fvKMu/i+Fvd9Vhx3cRt59ssyXL4jSEP6
nS/1kEg/WG4hb5jF9oUYhxqNG1EQOz+guwjBgCosqZw/GN37DMALCjq7L04DTn74XOMgfWbBQ4gS
5xTEGtbzAw86LNQZ06DjVGeRizmTc2eIGf82vLNj760KftagzT6XYHmreeYd4l1BGKRzWsUI/6po
9xiP4FYVHbV6J19/FSl1HhuZ3Xlx9Ck/q8bgMxBYn8QEU0bdedluNV8fgeg28OPAadeshFP24RUj
DReWUCFBBxTfboCYVWiHlbBeIPPPDTnGuV5JgRN51mYnDXwWmSTJurAq9mSJoAoeY35IbUlzGXG0
QD2A3oIDMAqS9LpsoTXDunUDFwoWJ6wMYOo5Qq4Ueaikhu9EESqOw2CKqesq507QyMq211KmMFlv
zXslqBLZpkCSYXWfcwS2RWmHPqkw+4plk+lmCY2KUPCPuFWJXdAt0XSZmtqjik1pkyECjBh4Rmyp
iYJHmEHdZKAvbTf7DFdfvs5X6/Gg0l/JSMRYaFvM/7B9qPWb145FnvJ9ThrCUEQLZcFD6RVGDb3C
CDtZPDVFRmRGGOO5kOwEtmj09MLLv2ByL7W6ooYzqNP+7aZ2UclJkRp5jejb5MI7e+bGUBw+npOg
WzQdtqPOKmECTkwVtSObBJArJLEtrjxlqh74fs9iOvnV8wgl46CHEOVCgvlNEkL7RM+Ub1wGnEER
5AgI6FLTy2ekZN9USjgt1h95zDBNFiL127O661U+nYc5FmAU9pm9ABN0vPlu8Ygrqzyj+WJPWYzZ
m+WImeAakdG9WgtV0hPgSnF9oeZvgawMgxwjEb2wi3ZRTn2Mv2ftIfuwe3qEqeOi1Ke11sPMR8Wi
4AcPSyQ1bDzVv+LNdL2lSwLJM5Pe33pLN5BglK3FX65KcbEXlFRgs158FQb9NWn+LCYUtCNu1wKt
l6awYQ5f6MIQehJIMrmou2eCZcWkKnMBlXayfa/5W/H3J720/pdObQ6M58HNUGGwD7wFSSuy10r0
RyeBgfv2Q2LXPXcKiKTqI6gCC99/icQ0QjCWmqH2Cn/ar688boijUtHym5PXVDgC3ex2L+gH65NA
P3LEoh66X8EGNaETgoL2GCLRLVfYjYaj4wqc4glRu1aJ4Ez0xdjtXumVxKW0srl6lXEISitafDPy
H6ZL8WSYhTAwC9KQPrDPkH1I+xVHynO1zglIPevWxq1N0NImjyUm2pxENa4KoE9DLlisFJkbaMSN
prVJgq8x//PtYwJvV13hlrZnyiePppG9dU/ChZgkcqY4rZceVcijqljJOw+4CatW4jYMnlxvJV4N
d22pZFtoG9OD7TIJ9PNTFdEM5DztbMnpHQw3tH36uTi8zu5EGQfAEwsLL/zN3bIZMk+BPtIrV9WH
SeTHgDLMkH5HfR1cOOKpdVrvwBEZaoIoF58fr5+MaZzx8+LWGzojjjXbBcbNlmlHGin2WynsK0vj
ycz2g6GnLUkhH+P8G+buL0CVOL8+cEW4RkKnxlxP+mAS3SUMhJLLQwJfNWo36R2wXNlT5+8Gb4kS
H3qBhCPIg0G3GlJJghGjykGAXW4B/fKoCaWAhREITimFLOwTkD/A6/SyOa5jRbK0NTCrfTVIDprj
R7O+oOF85uw+Nt6YqlMaUfncocQ+7gIQ2pRYw3HtwHyBounXHdbsIOOy13LL/p3ftLR85NEN84By
hXACiej3UnSBZgNnMq9y4ui5Q2Kc22ul1Q9nC88K+Rbfk8iGGhAZ8gtZDthyiR9EwC/lOSRdqlTb
h1JUTqH9vXNHrpjI4ccA/q6yy7Pci6fZweOuEf/hegq3tXPfwV6RKixyz0zItC3CPrd8yjpuJNfm
lqErOxwd+HfJga0uccqeqdeHro4y9hO+1pzgcB6mrz3auXeat01EGJZ1Rgkju423PiJkEbadZP2m
XO2OE8Rt/xjL8XoEDL2J6pMvyycq6EuYV761M8ecxzGhWd16i5ww5U5yPbJ6QLyE1C0k1FBTppnl
iIGjKU608zpXNYXbj6WxHZPlp4T+rrLm2yjwVlOJBl/0r+NQDwSfVoBqV5XVyt1rAxuEIigNCmou
+RgxVEoTYNnnmTjpKsDsgJ7160L0RW/JsP9KU3B4wgwEiRlnB6YG+F/35mRwZQ8gthzYlgi08swB
jL92HUP091MIcgck8PSIlXoPhaVh+GPEZiGAUyZGMGJUsglBOJeWu/uV0bz9p6ErFm2nDlPrTDQq
mbrQw+/JAKurPpZWrURTSZvOBMTf+JgVFUKgCS2X15xpJ8JiWJA2sHB12+wwo6b34FoXrhbJ7VqR
8pW6Df/F5nRKBjXS8m2JIdPZM9RgghXvzIhG5Csi8Bt1SKQXV8UF/D0PM+s5594LXE4uUOOZjdY4
8H1HiMJgacztd4KtHZfHkF4s4/wTwxCla3c9tcpMIarwb+2H98/X0TNO/jyhZd5JxiZHUdFfM/Kf
6fGv4vKICJmV2lJ/+L5MX1QG/ah4u9OUmrXF5D3YLFDVSeQD7pYFX02ha91wTXoJREf7Uk8uEsde
EU4hh6/HjetloiHMXoZNlDJL0+nWZtJw77uIjaUKv927NVVHZasoB9gqOAFSYdR/WWk3VCK2k0Dd
mxni+USr9DI2N7Nrm5RSZMch4JZRUpBRg2eyRo/8vin61qZVJQcWiBD/wnwX5eC/+N9ylzt70GL2
2mAiNd6an+TnQf2Dcn7Pv/hsKUOrtmFwrTK/0E/Kua+Q3ByCRLpGnZKQi/vdXeHPPSmISkGBF9/B
InDoOjMESKWUu5XGzZaPYczso09Vq1SQd1qrPG6GTow12/hriUWyk0iYjyGqWwp3LsDUZ4GyG9Y2
ZTaNHh6nD76AujqSPSFAhmmRMTLMygcpbN9MbC9pFFXKb1gNJihKWloezZgafrp/eaBNXouil0bK
XhfOPreg/O3oiy4tKQte3fQ1sDXxe3JSKWNaLM4RWLvlNO2wEvZ+OKq5rzrIAp6phJT6hdShaPK6
OVmy4ogYcq6vTKor3TtwZ4HUJlrlM502RAHOYf+Xak9YdIqG6gqPowatpEa7vXx9u4eNWHyOooQx
yc69zGrEkQF5OfPV8CAEECGfAmdIH2nNWAu9uDsU58F0CgD7Px2GBqEoXHM+g+b91thHBe7HG0x3
Kzuz2n9bLr2oXhTD0LGiGv6WevjWBmyKtQ6B+elXNlqG7dUTabnt3DMoH/W1qRvpTghsLRFBUA01
5vI4dLhJ9/UihubNT/EOSuB+2y9fOsD9ngbRffuAKhEX0clU8tb6Q67z331yrBoei+LkxA9vQmSJ
+irae+3hg56AIL/AELNNFVi/3fInwZ59yW4tlOI4VKOdg4R1+L9mpMuvuFhi1lp2tM72zHzTlavA
eKo0TedoQ5z/w9QEkEk+dc8QxZhvq8w+2cq8CsGqQCmwTuq1fhuyFAjfTDlFWeJimR+9KoDskShP
DEPP1N27HUvDJE+5W3/Tkq6S2bQXuDQhKklMyr2lg7p5WV8qx6TbT/vYMoPGgj04aKFv2oWnKRb1
0HiQVV3WyDJD6FGnUhGmgOfa6G7zfk7ci40SELsBesD33BGwPV+2SAF5F3v5EWfWdoDrXw8UREZ7
fFHBCRVEQncCJwPriUAvFhog8dk62VJXJUZ1ME/FhcGYlKqSJfT+KDIvGF/6/9k9og3F6y0rGX6Z
JvpCQ032YNghqwbNAl2lujH2EZRhOPMco+k2CR6Qt12W0y/qbGLFcla9H3luUhYmBHVnFHjRCinZ
ttNTdXZ6F4vWkW2N6GUvz5GJyTjKYL1Vl7KRwfzDIYalYYQOupb9gDnQruuzaaj48fAQLDt7t4wp
HWhHySDBn3Y02t3pbFa4uBZae1Qw3yGznshGl5GskqOEb01cH7whEdHN5n3qtnyFqai8lH6QW1dt
gEOj/j6vEwvYtvJJDxJ7lJC33G4nzc7Z5VOYbhMDycvj9+IjTUAmK2D4dA1ltxBZE83yfJypgfio
hs7c3vsx4LSi/zQTek28oQ2GKG003aS+LVy+Q4Z2F4npp20QHlPvho4M+YznkcK85FKA749ctbza
zCCg4TzK/2SKMFyA2yLr3U9A+9QhD+kBSq6BKTAXSMO8/MC9nFc5yGmHT2fnGnRg8ERij+pdKuLX
cVBGCdNrPG1dzDRS7ZGIUPpXxTtIe4C735jeInvuuwLho3rUqdMTHPps15yCE2OUQhYfWc3oWlCf
AoLjbHMwhg1OrhcjQw24qyTKosgL3/eoJcuULVkbZrbJbQq1w5iHmp1gmxqcv9gHjWuFhmGU+pV1
NEZKA5LdbC7e/icUKi8QqfRi630REICz9b2Rx5wSqinc8mD6csqK8dH+eLGjoLQeLEw4Bx+9A5Ot
ZPZaUytRGAssbJDAzKpAORV67atd7MPFTcSc5xMXzV8Ipwmvf8LIHM6mL1cslpMWJ61eRPMJz/wE
3tItyzWoMsM9iedqe2tZ29JcEsceBwSlYb65oltTLLvbqANgpwsaVbg41L8khIzLFR2joBwk94PM
BjDl/TytuzDhDO7PYqYO4zrvny0jn03+Pp4nr2DtfI3qIZj8GcUK4yT9YJA9O8hC7RM1XweLZMG/
+5YabqesdtZTd9bajNjC0QRhw9MjNfue7yxqMw8zE4R4mH3F/ThCXfIuzx359pieh26tzyW3jMO9
JJVAoKyUr0FFN4lcPdxY4sq+CCWwEIoq45yBj8F4OXJM8AfyHnhbEPRZNjkr4hXKzn0h5IHDC7rF
poZnc3CwJiju2UcD5TeNls9AVIbVtJIt+SKiPm9MOu0ypf8XU6T+KqZlsflQW9iwPGAFm3SxEZnb
VL25RQ9VrwCPQmxxnTgrzwBDuH3NbbSNFqkbLc09poyivYfPj5uujWy30dPGOcdUxNAip3PnuQG9
0OrP1GhfNg3MNaDBDNdKyqwAwu1qiCP4M0wPXkuV7AbPjk5k0BTAV1l7AtKIbCJrCk7keClZo74w
K+NKU10h6CcIoVYc/UgERnyMtE6cfMWPb9QThHSqF5gAEuF9DuVwgUHHiGYhfLwF4tv9fWaWX/Ft
STY+M1YPzdvvV8ZuAViEdsj50a+3Fn35OD53eaUxGTp9B9axZsnC/5xXQew6Ap4XMtWkcYzLvaSI
KZjX1mEpWgLwThoFjwaq9sQKpRwZlTy0qRZojQTdDFxowzyKbApoD1kSiPsPEmVf74V1OcUwEqSB
3j7mSWgfSfxQ+gTi4N+IW0SKPg5Dcl4aV/tud16RC+lo+RWqV4ymZDEHi8/6BAFFivuNS1Wk8jBU
VQEqYcYsDBBWRummD1QKVd9WGMR34QaHKC4KBlpzt4okjWoG75G7gFLKiR0LorgY6NWBTM7VpExh
Zh86FCtJZIa8e8cTYkNmGjVJFnQRxQCO0J8XKpyn0KpvMqPew1NnIkHytIlb6dxLtA9BdnQidN4K
DUk3RVi6lp0npnI2Ou4c8KiTr/ia7IRcIdMYMYQ2oHgNXYgd5SJ9a75eaYwmBH1UlLGkXHqQUwl9
pHJtqm/0PSf6nzUwzE0GwE1TEh+lzJLue42QuoxrkE2EOZ/K0P3mo3oDcUQpePuENtyn1lf4BG2f
g37s5a/kYD4IG2+zbRbv583hNPy0GAygxqbXMOBEpUkwAVxcghuSPPBOXTPueXNGgwhLB5+qgwt2
o9gfFeAA1XL07wsK0Mw4jbxmhhu61PNNCEQYX52b08BQr5MdDocfAMj/zFPTf0jSnm8Zk0Wt4/Lw
a+20VI7C/vFekFwtoxkdQWN/5a+BqkHjkl1hjA45IJ2xe7HsiSGLkFSSrOyf4t1hBMgwe9zh3h9f
+ZXmubWv+in0eim0aEv1nswRrB1WK4KA1Fyp6bqfvhQ0P1N4VzeMj18E1Rvcd9E1MVOpawx9+ruz
58N5k/LMNsRJD/BrB8W9vteeiZRN/bBUFIGqqDlRFoGJWERC5+kMQaHMIg3YZhZxyjU+0N8ibarU
1gxrI2jFKRKkQbJKNU8aEMPd9Nnz3BnskDmXIHhZ9wPEz1b+DnwlS8PNMDvMC3Pf/w3d081vqg0c
AR90oN2a1O3wjdKVyHsDIFmcMI16BOaKdK6GW/rINdCvwQ3wB7Ru7qN9XIXIV4ivEgaWF8JGznC8
OlW97f7wNT2Rac86gb1/t42pKkopSh5SRnc64e/pxHD3Rk/wWCqePZ77b50kx/j6eQ53I40CAxce
uSV2+Y3/xhFFsiRCc+OmeWFVT60sfYp27oJIzrnbRrd5f89zYDe0EoEERrBDMH+m7ASW9AEqADoP
AayYdHEGinjMVyEnsD7nkTk7I/e81YadTMojPzm6uSDACrqk0pEveW7DeY6YH9fWFJSc1CTK2zAG
VoISSDkOXvqMOziW8ML6AB9JtMqvgKFFGfQeu16p0c7T5EBD+PH6B0wkOiOrUD31LH2dEr3PsYeJ
p35W0ZCTDgNPCPy/dMi/4fkWTA23jwKdQTDVrb3J5GzIf4wfdxuehOxW3Rv9FT8x4cGRKGhAwxEL
Dr0yL666nB/OXEu2oJrQFBcadGTn0llgaFVEgnlT4nSHihalQqacW0ACeSBdh1UL1ZdfzGhkuMS4
/cJmcgLmogIKfxns11NYsWpvOJ2rMDHIRMN3FOVG6PnY7bVG4YQwccwnItVu3tZ/0LlxyCkw8Z9I
X+7FAoyCVxunzILuvBptP9WfLldLhVItOijUm9lttRQdiJmloDwCjXERmsda9pMWs8+F9GVzz/dt
tP5JRzT3zGdfytWJ9HNQCVYsWCO0iaa0Bl8TNOR4GB9Az9MmypAFnYShHvbkdi/5tF7Ze0NkQ1pd
0rLZAENXMXnDYCtZ/jDxA1sRNVZDK/niZIpqCKrevSjVnATay9AUJKSFbVXzvysaL/8Sc5raEUN0
MIb3Kffe4F9aQWGTux9vVWtCB9VphPWaE3X+yFYIINVyum3YmTgQiLb29LmPewQojC5rCGtnb0Kg
sl6RoN0T1B9coOysxFrkkrTI+PVmOZeY/1Yrpw91ax6ST/i9DB45wvqXqJGmntFBuJSl48+e87/B
znARh3Tpcncm/vesobPbUMUgACPAkiF1AhAUyJA5DzvpAaSB1eUUTYNwFoYh0wJaIgbD1uDu5sqH
XZnf9HZJJG2jir3hd08WDAZsBbEQKcUDUI7nsaEJbZd8dyoNDxNZ2HD6cUi5wKv99Qt5YcroSxIA
lwrM+bjLSN08xG0M22PQtPNdO4u/nGm43bqsrffUGrJRA+UYkVI4ArBp7GVLVqVIMuyxUeX6QgZd
6EJcNXFjeTioPNAc5eJ1ZAUo5dFFYrcGC4RwGEHRhyc2Ql7/F854697wUYNIjuJP1MnujSD9GAVB
512QHLcmaI0u6ViVXh89zMJ/zhwVuGaYFXHIWxXTgT+LGI1kZnQLhA3+5D7sMAcyVmgsHliGN8/W
At7Eu3uYz+g/6P6ALvOMjVUmE+63h9CJPiRlme0fa3Yxf2ocKfQw7ZqlztA46OhQegeazmx5Irn0
DzND/qMWXzYN7VGkfUpx/WTHPgVz5oC4k2fkD+LIgAtPTcGfZgU+v9GHtKcqaVSlL7WQ3YoQykfo
ODPuSnJ0wVsX98niofgfwgoeP4zY9GUr4+aoAxvkRJ+L+/Q2CB74EUBuyeQMF49kY/SEa8EoaQ2R
IZgjrYsj0+K25JzGJwllYjyIizDeOtZD3OA8VARTK9rLrgcbIn6AAAFZVVdPnlxqNBJYf1eBZSMA
RZAm4NcSYA2A2NTwXScBYkGKybgti6G9W3Z2ag7Jx8iAqrffWgEyTAyyzrZGh899LKTPqkeRJq1g
YUTmc89NhgjXVT+T1qlhHyqtlw3hkHvzSlulaI1Y2+5JnWP4UBSyLzoiJ/tDGW/wzdJbIRjvGscu
jA0p4xLJ1VQlw8kLGbn28UNZMw37FFUYrObFCelKawp0aLRYCzmdxp5I+7fD9NMUbU2EdkTfDoaa
lI2GkBRe3+IUMvA1sJjcsZD7iRKFGTV9skP1v+E3h2RiBNPZplrgCI58LbuzakyswznR2F9ijfmA
xcMx6ZJiphdImPExNrGVvLGE7ruJGnevBg0gbYm9vBCKbQXxkcPzxQnEXdczgzUbs1YW9n4R8GKq
t9/S/ITX4R9QyCiu265IkG517LXNwvOVkeLYFLRtnWe8FCBJ+f1YbBgreivZQPPkqqxmoiGtYWmR
3pdcsIEGiXNdWBLAq72rGRvzf3v2cO3IGxh5uZ4TheWlMLFe/+40PwxYRF1TBxh3e/8H6wEJu21o
38XMhKSiOGQAldiJSL3gB3Ep+zZXRDcCE2IyWDNjspir7CB8Gm5e6xLZC9EVNLBKR+RXbyU/0QM4
1can1Iw71HF5uqNCqh5E9V51LfYg/Lj3ll8PjvhToU2B6Cs/1mnTkKcKmJA0gw1Ehw029Q9IcNr+
9kFOc2TVZWIclF7L6vU67XMpiSYzM/9R3w14cyIJCUIJg542rjaTuWnj9G6GTUVU2aVgm/AZ/1Rg
kDLIhzeR/qvd8l+/aEvM/BJhf3XvO1yjzJyyZKJ7Ve5WZy3LQ7l5qPy098Av6e9jJ9xN65V/YVZC
8+CyWgeyx+XD42AaYKIAsiHIVek6VnEmvsyRrDHai7u31biIsP82bfW+JDgnrqlpafOEkql7W8WB
fgiZeJ49F0eGhR1x8VF9S5TNRBnsFe9kZkRMRG0dvTTbOSsewQxLCeDowTSvNmdLUztluw21xy4H
w7RcBArf0foZtbsNevwrARztpYZzJmT2SDs1qn5dOQnZXqa/DN5hux1QqpNUzQbcuwjXnVfOL5xQ
9FVEdI1pjXvFhxOP3YoFzJERMyD6Uv0tnj9ZmrQQyzA8SxfMAYZCSFsQ5z+h63w1L9nn5/WCWMVb
iHpb/BKgUhK3I9gQlU4skavgt0DTIIG95uyp3+Ram4b3h2lI1N3Q5U7H3oB2ebrXd1SlvntU6vRn
WeL+jPXwytPRBsBLzuRKqlLDXxdhtAyzIGKyqsKdyA30l99AfC42+5vcuSyNk4Jmsi0GkmoP16dx
P6jMzYs0qM8uFXpzQsIMP+z4ZJCT58wDj8hpALkgT7owDgTYPufN1hHcoYDdQIbk/7oVA8+c6IuF
HybIsbSRYSia+1hMbjJzyVtxMQI7BCgAA7MRBvZV9zPnhsNWrVVuVSgV26hiw1NQBMrvar+Gdab1
ZeUi5wUboSjpa3RV8wDEgaMCsEUHQDZDb2ECuHkmulQGuQZ6YO+k+tMVPUD2lUrUmjltW/J5OyL5
wdnb+3n8eKmtTonRhr2fGeD7kd1ObamsCRf4m3LI+nzf9l2IEj/jBysZtR7nH84rtNDjlZcYG97O
kpuMERsDpxJ0YwkEqB2mZLJSv4nK5HtVh9LwhlDO8B5CARGcVJ6I4y7dro+mCWCx/9T7qCLLwrNJ
fPnEY+CvEyiQk0kA4q74MsxhCftQ0YYD/YJ7PSkciyohiXuBdJLhAmzcR5w5JI5bTbuYQwIwiX8E
OGV+20ObcMpw59w2/t3LYp+QjQSqUl3Xor8GN5jTIw3LvhGm0OnppiDyF9WSBIzx2TbbVyWA6jXp
Re+ljqrZC6+nKYyHYp51lGhjXNOr4J3lwOxdJPFkH/jPLbnympPRX4uJhA0OK8/98keqyOPrRAHi
0bOiFoJKvnr1Nz33mnmI7LDxmk0i5CyrEhVzbNSa8UQnqMsP25EXA0Sohgn3rSVdv8QG9PnbO398
LWxdl3oUf8EAj21li3OSrKYzpkKPiH140ixrMBaCznhkCD5sDj4iXBCUmG+3Hxlhb1micU2doh9k
MrUTmwRGiVxHCB/GxzblG7FyAG5t+ve+VdnnVOdscsJiWJ6SCIF5x0kM3/cwseH7gV70qShoWWYI
GD9xDcJVUOH8tAU3qxB4swJduNUevP13zPFKQ9zVKO8pB9WLi49mZ8UKNx8GWKdKQ+YT3cwa7+mx
nXV4FaZ+cWVKPz7DEuS9VDSmX/PuGmF/CbICCSDuEVrxRb0LtFYbkhLmkvNUGdse1Bpafp18t9Yl
xFt1q9jgNIWj+LSENVaL6YIpSSzXUTCQ+RTDClqP9PxNnuMiYH9f0LOPh6gLn9P+JcClmW7cP3gt
LJPRl+CwLRPAEeVvy8f8vvhXXlmWPvjcl/UdzSsvy/Jjrv0fDizVrIopo6wBGI9oD0tZQ2soHXek
/ORbr0OwbW+ZQsdG86Ph5cJgcHqT4huYFjVrBnST5WfRqbdxc+HnNaErbU6r2ueOub91na5ccI6/
yNrDUrULUOKAhruPFWSMWa0Gt2Ztd+U8W8wh6iDYU4DPF6qntjR8hXMcbRtfm7UqXMz0eeb0Xv9u
c3AQ5H+sLzaWMFEs+4ruXvxJpoP5sSfqYszGPw45nn7qDhcH2DYB7PVkfokgt6PRx7IDCVEyzvVI
/SxmMuRJefrX/R5PEsgjwW5RRkFbPT0gqutUCOdqnDIlvYXPLb6a6SkSCl1dMIFcAtm87jBgEsWR
UROvTArqPk6PlerxL/lhkuoZWfx9HWEh20VUPcTxhKT0rItHk+NZMNrWDg+BCE1u5wwrgRgJtPOT
pGF/l6kCWX531KZ3otUgg95Y8ttJU6ptjbqWHZFsQdzbxY/UToXxWsmxJZXHZVbtbp3gxkKtKT5O
Bgt0gNpdyVtnCW76xqL//yjwE1CJxc/mk9HMMz6k7XvW+A6Cvk49DwkUKJMSwEWX0uDSuaUuL9c2
U9ZDdjbm6dQ04m3bhWGn+O/AVntqesEp2hOoTTiweLy70YGtVfWSq7+wxFt0xtRsPPB19MpWWEGk
29jq6QaDfcsOP/mPTt9dOYuEolMBGIn7fnCPq8aJO9kzAyO1VET84gYN1gOR6+h0LPUsSSZv+7/3
YHso3rYWSKWqOEssX7fCnzgxsazFji754b766weGe+hqEoKg8t+lPoZHKy4CfSTHZAza+/Jd73Ib
GBIdIJNjRKes0ELpPuDLilqEQa8q1nJiq5PAh46s6MP4GBGQlB7Pkbw8G/YVbE38u7dpTgQKAB5Z
KyF8U4heea4LrellBbd2HFoiMVkzBQgQHEtMB3VcyqZJE+0+PFBecsoheoWJ/1cW2OTcf5WiO88D
Z/D0rxsSpfMihq7Bw/v1+sBNpND9upeTKjU9A/O8L4ALxB+fyceXRBQYg1ltnHe0wuPsmLzWl7kz
uam0ASLmfl7rkBj6JvcgvxMpNJG++P0nztfcGGxCGcwOO4mPqONqc65Q+ULvjb5GlubyEzezr/ta
LB3mcoRUxHuNORvnWb3FKZutyzGH+zEKMRFxlnec7TGLzxE7STdO7ooq5+srBKPP24c9+6xwEuu3
EEK18EdwTibMoSQAGowSkyxEbVYLNvzXlkIw/hoKsA+YcbQluHGXIzyiaD5kFs2flmvb+GjPQlDA
P2cV1tIr1S5CLQJ2gWpeEB82fGVbcNcTidS6hx9SE0BhVrceNoOV/hyjto84JQXfX+GdAC6k/Ubf
7xUA0j14UroxQ7Y1doy4q1OBHwMpAUzEF8NfKjFN1d0tTBpoY+HZZz1dze3DCtNG3rbvB0BTn2Gb
BrhIXkzgB6mAYl2H3fscaj+ZGm17MIyBEQT3ABW/bVNEg4+SD9vBP9q2FsS/BZI1xGJ0F7Qa9aL5
sDVXAV9DdMs/+3hbdibXS0+6ZHWJfv9D0GoBcXjKxY3vXkBt+xrN27+K/jSL6m8pH+uzp7CGb42o
O3OPCCqC5X1KwZJklVlJvuoSXTs0ZOKKBqOVgrnCMTPcjMPJcJrltICmpTlgeZ4nAb/HP95hN8qI
k9uzij4zitZHjwLC2UkduGBlQX1ewjUm2bIYJ8uTIrBpg4pwRoFIbYkIjs5SyGPKhMUUzwsr1hJc
KZZpHzk0SE0XnlcYJG64UfITlzU+Ep/rt2kcb+augh1aagoTM4I2GkIBcvs5l9LPHWizytTkErFm
dAHQaEhaUAwZqaTTPLlWmJSOlkJtfuZXRxMdBJ+B8IUTCyVeR3jtVn7yiT3jcVozPaKlvZXubs4Y
nYttLdEXD1EH8qMh+gBDhWEYHEM9srMK6RzwuqBA6kR8La5c02Q2NiCgqIDSEdQIYpxmCNENvSKK
YFVDM6xFlHBVUJYGLbz4DGCL9XMV3A8ShNqrj/gRWaobsOK1xGBa9Xc6AltzFapj0pEmk4oyezIA
Ws70j+FOdfMuAvNCA+KCqtidrWAqdug6X101uMvH9sb3V2CmlUfTxcaUxoyGwz62+GsEjacJXT7f
8GU1ISssN6IaB4Awp8MQJM9rfYEICy2FExC9KnJ+F24S6VvSsTLVrDxoGcUxqb/BJQ2iIAl+ZnaB
4UUL11Z3rW4VshdtxG0nTQKvFIyemKF4sSLiAugN3YD3eGE6M43vGKLQEjhB+9OYNskDQ2flB4s7
yf/U13h2jZmiWUcCa3xkBgfpq+iXiAlEccf85bgpa0/OxJ6GuqXZWUyqXJd1ZZjQHARk59EUK7xc
SubIkYzmIdFkg5+pE/m1kbhDniLgiHMJoj+9NvScNOy0eRdxNAI1637suWjS/s8eeR7NOAdyD2J0
sUWjAAW41toNwMfCx+bKwd/F0wvUbKRGYSsBkMmm/nQly3AhmLl9JE7qWfS29nzPOniTF8zU6zwk
ku/FBkxcvmI2zl9YG3Ve//ayTUAmoWHDawMxbkxgWiFQ73Zxb8I+K5QoDoc0Au4OIOGARCekrDuS
p8KXFIxZ6LbbjW+lxRH+YRpDx+UXGy4FKnLjja9efxtKESNrgu/pNth3rAIC5NKyx6Sl30LjDBk2
sJxtoe5vasTgPeZSGPiezkGsb0WS9G5waG4p6TTVQFPug683LtpBj6AlUpaNc/I2NpHnknZu5FNB
2aOGl7Ii5Q76iOjHe3BoFRbT2z6I6yJMtmXLZim3nL0v74gnKqxl06WCK4ZLdTxEmXwQrqwTk0fb
3ZsJ1GMaTcqFbBaJxpRJqB+qoXKUIND24xpcr1yxAR1YFHYB2JBxmNZBu9nxj2uCT0OGdOHWVRMm
BEvyNQy5nOE8un+EG62xhlNCzKytUifxq8D9ccQVxSWbV2PuQfXViAvjBEHOL4l4vbkZu7RrGBXi
34tdm5fO27Umvn5YJdPNe4GTHt8mmPuHb5gd2EQiD/w36zEPTeqW+a1FHNzHiOsCmtfPk4/9A5MV
x2hNBwrgdMPzYxrs/11Z6UffYkZqCjS7/MLsVdDUA9UFOWmNdjiVZgeJEub+i0tktmfZmGP0IZPd
4/0QG5TZVY5qLpKRWyJxgeY9/7mb/thOCBCO7IeK69xMQQhDs4KjHXovbnZx1dxzfJiigTVxM4mA
MApToow651opUb4+IaEO+6kwmtWVxEYocLKAVTZxtXq4esPo1rsaSwyl10mZUsjjXQjF8FFFc+qf
CfK2fj4IOcaBoUzQg6DUQMHxg6MYCmyqHm6YkSLnPu7IeUQHxGUxn31Uan/5eiGHAiM8s4udEivE
VrIQKmHSrSsslofD1i4YRx6/4bVDj8TBI7tmcL37pxS/6Cjo1eaOvAOraOQlcILNVLIDMX3CR6BC
PbgUF1YAeKiPNC/fnjgZz6f1w9KCITz15NLFykpPLH5LiyUDeOq/J+RjTpi1sk2SeqnQHliiBzpA
1UedLNZPBvqff4cYRS03/3SPMMT+KmdIssxIhw+Hw7dMeaRATzbp+ZV9ZJbJWd/oCXresYVg2+9A
36zteQjxjurlVkz+64PYWmzMcxO+DZAcN4HFxCTVUAL2kAA01id0JL+/h6ZDPBuZUPp4PAnjGbZp
Qpb8B3mqy9dhypr0gJe71HWZuqpEtAtLZtiu1WdbtpIHfvXTxvHDrOzSTnNGZNEbZv6uvAFrYkjp
C2ayDv1+oXUdWnLY2jWwH/iDY2auvKFQNFaKX9GGRh3s4rzP3k21cLoxWNeSw6/ExMs1elV9c/pV
QVDeB6811X7gWfYSAXmJs804Mug6939l4NANmfboIOgi0Yafhld5e1cFUF0ruuqfXycPr80UxsAK
dGceXTMynnh+8tToBWaRnUeobeQOfgCRa9Wj1E1FzSFmN+TzWPiohHEwGKwUmJpmnjZQcwprb6Zt
0bR+OyEEi+fsCB5lp+c5Qiioz1LBIhmzCuJxySoqacurvk5GoxmyoRWGHoVssIxb5MyorGoEz4jj
z7AwyKDlqqn582cFoU8Qu1Dl4cIK0q4PcSNgnufr5tZHKOK7g1lPWk/6hF0UhBj5riaqlXiyBrrR
/6Sm6Tq4Fu5P8F49rN5Cq/sDYmnEYO2HE2aXTY24wC30zvQ0qyl20pOmWAIgnMyHmPsCXqCRZ4LS
oSqjqVMff9YolhYRd0M0JhaIDv7XNLaf5Rafgu9PeRzsopK5p3UjStApU8HfwQzsDhw7K8GqTlXO
UVRKi13vttMb83IOQ3SIUYwl+se6cQ9KAQUSNgeYFKsqKgcebtFWxvtY1Xg0kjJEjvgS5vBQ6j6G
J+e1FSjklWkeCssWd2rEfHExFDVIsULWfGDotyffVhRhf3xHVwHD4pZ9goUtPPJg6zTwUXccQQFY
7zdTyNAt4sB2j145DR+KZ46fDsz2lCz2MYNm33ZLhf7XRH7SfeC3bbl6HIoK+w8XL8tbgQM6jSKG
6vSaQ2IciDHWW9DhgIEJ6ZnM9m/GPyyNk+2TcKte2ydEgM2YBXsODPgLqLs1BW1PGVVvImnQ7jk1
Kkcowm+9b9C5aHIPrhUu5F3Jn01F2Orfvk+5ya0cL2NuXAEZRJHUnp+Fjk20j7eE3Z8fwA5VHYwR
0IDJvKH1nkUGj986imKDXA77cQ5rk0EhF0ESx1D92iPeLbUyzy1GfR7hkGXULQ5WFQtju0T+sntk
aTE3VHfp0YsIAdU+TEMJlqjykNHpw7EislOW6EdErJJgoAp7tIw45quQzFtdEKigqRvl3VGR7TXt
lACjjNWOg4tZ+l6TWZYq8VwdUX7Jm3zROwrKzMon2Uwd6VVC3gZ6PzPaLrJF734jS9sCTPuRDn99
ks2vXhWjLoE7g8VSugjO1T2xWcawhfmFuVf4+U9TuA3bBWnUhASY3MPRA8YZ6LnoDZ0viaIneJ2V
FWZYg4TA4WMnsJj2BNbtbS8jwV1h1Gk3xoyIHrFqOjm87G9Nz/CkzDGJb3jBn9SWBs9m/Aobzjto
4OEqrGdxos9yh1h5WdjgPC0HnXvD6h3qp8RemE04arMKnw9uSWUTwWaepIuLWZvk4jWIJl77LhDp
QIxZNRaNB4gLzixQaGANlWjxD4xV7gTTfnJRROusrMvNmPDRiSqM1gKknU/HUdWTk3qGZQZ8/X8h
Fenm+qzZNn2Z04DTvljT8A226dbIQ/hpEc4Q9SD7CCnYogDseHVrImewYpVHTZPxbqPHuS5aDtgP
FD7kysq7ZrDeyC8eGCoTThRFRl9biT2w3VLoFzymyU4qgN+g1hypA4bCsHzmTCihA+SwTr+6IbrY
IFOIo1mTPqhju+CI2A7bSwvGCgQfgFZIjriSnuGdgyzsD6GLYKnxVLdO8bceurLZM+PGdoT0FHm7
TtJuzJrWujdvK3jBJmxzQJw+Jdu6NCzLfwLGuv5iRXUKEbf6dejaXRBgDiN7a03Z2VDt6HPJjzQq
A+kcu6vOEnUwaYnZ4oL04qmnS/orh5LdKYqZoe3mgWCGlpwYlgWZsL21fHPoFGtPA1AhyqYXxJmF
Hp3snJWI9i/FlStg2ghzRbKNmiyZWgP3gbJsLevxqGqlnVNDdXIy1kaoufcJyLMsvoy37l/D+rLL
LGxo648fyIjf2k5IOmsRqUv5qLvWEEIQzt1wPukixcPhZppFZihxkVAcf0HCJvsHWvz3gnu6mqln
3cboI1IfKuKKaKr5ZDWF4cSmsGw+d93DS6ILYPXlryJh+znue+9Y4p2x9bkAsda3RNi7vvna0rH1
4FwQYhD7F/tCyzTN/0UlRDGgVpM4vpAXdrWsaKGvmGc98j8zFfjulHc/SP6DS+Pm3lMQAYrf6dg1
GuQQNQjND7YgrA7Ysu7Ys9YagwcAvvDntCk2/6LnSExmOx/tYgCvpsVpnsi4iMbwj6L9rdNt8pBN
UJGlaFgq/jmT74JSecQYimE0hH1rNajhUop8hcMKxPMn4iQtMbOqsVmJhB/kCWb80M5jSlGbiKaN
Pb0TDxloTH+ndTSBqN8n/oseLgumkNIk1gA+nQH3GP4Gz1tJYFSNF9r0M2F04fpOhOuuWqxZTRNx
tte+UtN/0MMSIPFOiF0DFh5o6OPZXqUmwzWBDNYWenf+/vhwcFZ46DMi3zq2AwWPVXbelSWXcaWG
FeuqJTjmu/APF+fLL6aedqq7sbr/Bj8f76U9378Mp/igzXhSlBqLCeON0el2lRc/vwLK07q3KGY6
8XoBRq2Q5tnFxX0LIxkdkSTkfQbLoaDyj99cSnCsy/OJyEYc9WmBeSqyFHkxv5WOryu50cBk6ip2
n1UdJhsldBboZOc7p4CQZUcouseomnp2Lb6EefSz5AiQlkVoVnDv5FzknefZ4TyWNugCkwAQrs6s
f5PlUBi/a5WljAwbUcxRpyTMpolDt+Ier/vZWsZDeE9q7YgGiYMzrLFoQygs9D/GtjjO3s8IQ0UA
FxBKrXOBZaVRQxx/c13wCrbZR1oCuiJAWAmtrA7jdufAX777jwartRv57F1eqD56lnxTzeZRLQAG
Hd2QQkfp2mZ4L5SaTRaghTk17WZrSonOee/Q8v2mRehzPX3QzyjHpdjT8aZbUUhkL+AXY9hLpn+i
FQ4Nij24gCGGpn7CdAQ2gpY4pPNg5fEs5dWMW1Cumos5rHnhXkYc48ukRmZ6jvQu6gVTkKizbscX
/8amfxQcUut60NdnLVhhvbcAHvguK53PXHc+Lbrw9oB4oOKbL2H7jR0Y20k5Lvjuzo/a5YffXF2C
0g/WTuBa28K4kWxRZRFrE3NiVJTzLdbhYwJpgk3fBtNiKuqA+p+WhU/X9xDVXl95P7FrFY7FZQ30
L077S55PU2v9dLaFTmMxU86aJCS+t7413ZKx5i+6oGRmyyeZP27JvXtPC3vTTZ7fGMnTwwXX5AiI
aUNDcZLItF6kW2S32MA1lozQyBksgF9oLRZs37jDh6OwWpije0LiQ8D7qOpw1IzuLJQuxF1kWae4
l6Wnjk4qTaf/zX4gGW3u6Q3zN18Sx+oSy/Q0JeWN+pMoY6Ns21N48jjCzv+tW8+bjAMhONO6KWn9
wBpB/CW68OtaCXTGaSrkvbX5Fd85j6Ef20gmArKknWqUzXZonegIV2K7Sh2MyR7T/1Bf/rtuE7wt
L64nKTzsypCcYRdgP6eZOfGOpod+kHcjyNbs2V1wUfs/Exf9VBAwHAzTTz4JtD25aIM6QK+sH7G1
3DLePwB38dnzpKdOQPpJIB86HCDW2DLNthvA6ptyEbu7NLJf+2VW0ILQDDHYjkI7OWtk7qK02tyi
wGoMWZFnuqlL2uKYwxZv9IBXEOZjfAqMpaf3op0oVPxABD8f0Wqa0s1zcMgsXD4aTmfFiCXA+txT
W/2LHWv4MLpIlZ/EKTyYvJV9jTsvqM54ox24JRHXeZNzLuAqCLbMj5tfRfWvwdEk4co+s2HtSwQB
U6RmHzQbuJ/dyMVia/F0Bbtj6sy9v3+snw64oGIbhEt6JYSNgTchD2wbPKdNeDd0NXGOmf62R3Mj
nAVANn1HVo0t0YouufAF2cs2/S+H72UFYU9rLeEDtAFqu5yLXQNjw796LTlKIb5CWM7Gvt+eC9Gi
/qaY//iDa64AVWdWtBZHvWNKaWL0kTb7HNSdznYaQsAjq8vhYN6SkypHmiIH4iLVDAr7ouIhsfwy
GYL5dZ2ssz83zx4Gg0AnkikFoFB1+3LNNLVnuVj1ibD3BEgUbwixo1OoJHLKgaMILqoMFjUi5kdw
2dpu5gJRBqkoGh1q1M3/sV0WMhdCRTGsPIJRbmsPReb8E4+PLBW45/YjDaHZisF7mdFQWHLe5J0e
msR8b8HxLxXlTlg3jAfSVxw2UcC5JPJcqI1lgDuSgAp8/L+lvuaGNFHFrnx0IacpFEegLY31nZHB
VNujxX5lwTbwXi+KrYu5p+tpX2vqxPaKLJnBp96AGDKpjg08l2SOVfBjP9VpEREMbuen11pAivky
npewV9jBk7BcNb4U0uQoF8ua6+/+UROOC8kBD46AFxyVZLR66Wq87erKvLLOHjHXNHEu0viSGE9z
6nfuZkib6TF1MsHjNBmDatOEm7lgyAsElV5u5vYvZkiCVzqB20SyjU2ESviXzzJjfTeePCXR6U/1
i3RCEmJbOEJ/Roibhe6qesSiMWhyNYyha46aAwceJ8gbjENtR3jQbVUu9PVNHmasYSU9dheGlPn8
895QZkhOFtiUYHqJ8hrCAmzBaAwgQC34XiccBi70HSWCptYEpqzG7bT8ihfiXwvOAKUoddjhFWxy
EsKJjlmA8lqhitHUtWbGmI2X09VZqEQbVutfMxmyCejLlQuHo5AY0I3QSAEavLL1HA7ldZjfJYfJ
IVKOBiFAybmUI/UhlHEF9vh5z0a1EoKTsDHJsr/+WIrpPXm3yJr87DCM/PEAxFVVLWrKwQwNBZiE
s0whMuo2OnTcy7yJ0aoWGC19bDXMEBvb3AVwxVW9YiSob8cc1NUfUJ5LP11tKLp7dZLMdCaiLuEm
PVIUNMHJb83JZ0RBwxNl/a03L3mQl9uoD2GEzpbq7Vm/7iZWUo4CyFylkOymec2qQx4MWLfsYVO3
5SXEkQvdsC5l0eyQ3YOS1B9Va7yTudeIvClWrbKBp+V3hK2aU0zWjU0l/d0W8yc6YaU7fingevAd
/xoIrval7dk1/QmV8OcJONLhEp9bobIDODqIYRQmf88ArmyHNbDJ7DaQf8G6tWv8Rc3N64Z6vwKd
bkxJHqXZmW0n27g8ExKT8Gxxwjx0ukL+DMSfXmBjginS44k3ZlzJHbyoY8//UM9SNcO0ClCQRmTm
nAACoatjIIIOy+5YflK6waOoSMO0jTO4P8uz8tdtI8tWnIT+V9UlQUCVizHOeBiGmWMPJCJlXQhr
19SMaIZG282hVne86faN4dFnuCqy7PzikRH25Npy96h78FkhHIceGqLuqrdb7eNlXtmN60oGLfYR
dQJnhbZ5/i+CagcDqnWhv+i4AkHvU1zWO6JWSvUkapybXibqG0gSHOBPUWEClN7LrHkdT/fYhGBv
63WfxmRMr8T9AAQf0YEgDdZPr0w+pLlSU8+NdDv1/GfhQlDOLnieb0MRr7LnqSwqaD6Mjqx5PZp/
BZ1O01MVVc78R8jz2YQyZsZQTKzlfBDBfER3Ko8P/CbLXGQCc9tTRZBsT/9cEKiLKZzU+pW7eoKV
yiwix/h/Xt3bUNuhV/HQbEgha4l8v1DkSshS7EpQsRfAmCpraSsuRbvxkAimBz2Eh7nsCZ+a36T3
v19kxZIcUAgRsbRShcbDsvUBafe/0pnn3XMUU1bk0+VIYSkgeRGBp7KJhXJeqZAz9VgU5UJ+cchu
4xFSpgQHGwuR47F++KDvKLAVLgDiyCfv7c37MjZ0kTGuvfu4kg1uvpbHF6P/J5QNdjQ7yRsGFK9C
yEYuC9Cm0FYwpehr3VGy8ffYWERPcUee8RV3JnM6ai3AxNhJHi2bb1V9RGhDTfXnUQI2JZ5omDKG
dboi+WEjVtoYWFd0AQ9tT07q7RQjoNDauyzuIGET84R3idZkxoFXaS04KO32ww8oIgp7X7YIXkgO
Y8+bTB0V256YwkClkEcfgZ9deEjLdlwGJFEd1sOql0AOzTuC9ymc5JRvclussGvispaVHPTLXJdz
U6MkBdLaff77beOjYpyNs8j13SE7k7H5ElQbHL/K7gyKOhFWiiJQZLEqV8dT4n5IdAKZB35rZE9A
giSDw55fE610vw2uZzsSf5CfXSJgN7EzSEt/2nRYBNZ41GgejjZfPBBbJJLEJseIxRzTYhYAe1qA
wOmuznDHFtg/0+UUYmYrFj/MM+GdVlDNhl+tjMoNYqcCwmZlVfHZGTXKFox68Ac9gxoXgX59UPiv
iySzkriRCzHrEOEkEzs3gYvhWe0Gh+IVKFWzyZkhqCZjNbdVErDBQGA1dPCLpsY2BSLvcZ/gd2uu
+mZ6Pef8ktGgk5mpHY4+mHY/MVHJutntU9MBYseWXwbQ4l39R5nDk1It0X6Sz7ZnOVTU6l4JRudV
Omszo2RVwC2T5XJwQYDOnXKZmfewNwNl52MLrFRizpg9jEmECrf4yvH5n+qtvazDaHzB7lXcc7HL
kRaIvL80C8sATsVLaqxekpCHYPqNF5wa9pppNR7RuIDVAZTp/mtpR6XnbeaDWIyU2wIGLRMnYJEM
6EOjHRvM6pP0GhYO7Imesgb1NgvjT4Pn9qTV5SFFBUkMJpy+1A4y66e8bEKKv4ZJsJ0D2jah76WX
Q82djJJc1GSoUj8vB9BWDoWhfZzJunJVxZVAoxOoMmbq0quxeYHaSkX9jd+cw4eOQd2dmlEFCqjd
Y/x4VNsx9yZLUjPicuN6w+Ggj8S+ght2UTEcjcD4ogtuSqykuBNmKQmiRF5cOPyH/prCZkrzj3sw
pexHI9a8EwCW0K2dsGh7JyV+itFaCF/lZRkPyxeyKc3olM52V3HOpIOIUlllfp6tvkjOtvVPcSly
8K3wdEth7e+dDS3nEkxhxapKoygJ/SIPpt5Sh7YMnQf4kGXWs9bICQTVKUuqzlzQ8S3lIWj64xrD
DpVuJe//Oqmm23Ono/A0UCBoEyT8FPlJ4ubr2ZiUp2SGA5QZ6qTf8rgHyvYEuY7CMn1O1JhlY0vd
hhpzeuZJEHlwu/Ck7UHvwKp9upshyE0KyW4cyvdMfv9a2fctNaEwIpIbWXqSCskNyBPPDgEKa+Cx
BlBzHJLImLvBFefY+MLhS+d4aTk8AN5xScQUyYKAmlxiKotW9Kga5wCA0Rjrc5JmlpKvwHgvwZZa
I0LcxQ5vzEeuhFEvx90s/14ZBLnc9hO0eQTNibrLoUYPYSJiA85Guv5KA27d4HkI98ZjFyo//ahK
pegZAoHKkD613xPU1dNX4IN8j5I6v7xCL4msodjSCLp9yxlWj145+wlgQp+DAqhOeJlS3hf3Nw77
wu44yAITYeRg441ttiJgsjWbSdoqg+fo/XB5n/ixb9MIbr2i/HZcuft/wcCRQCC6ck3r5sqiy5G2
PlbBia0QM/2RFkmk8NEj9LoWqnecSR/Jii7dsIrHHHCaXBWTcOnbA+xMZG8lWqQ3pJgSwup6bA89
+jW6W3+ZcPIAr33C29srznwsRpXP46Ws8GHK550lyHU8prKAWEGMgpaIrKG9luqeAoToGcN/oiqB
5QY+KyrnYWLhV2w9TdGMMbEYORRGA6cjca4CgLgDKv+9AZ5UUipD/4EKxWLAlJanCKB0jvGMtmbt
HyNe7wFfaxRSvuzQMfPL0GUSIiVSiZLc/yzwwntjLMTMhq4qD+UrT7b1hq6SBziJ61d22sppSQSC
eB9wCUiDAu177V2rHBF4q0BH7GZRUCqZK6TuydW4eahgzDIYDj8LdTER7Qj3myzYk04TpyifJ1y6
CLkXWMcsgGa62yxxWNQ5WbdM50l6BzBQZ821zTO85vfmdaYUbIEDDzsIVnLO4At9r1KuH+dSNXTH
BPVXyaaPqRgz3muDlIG5Vvb4uE1utQRH5kbmiue77SZBiWI2TEG8WmAsQiuZeb8wASufwfIcBIjR
B2vZ/qnbWUxZvOJfPi1Tc3BJ5ogUBELadbxCs6Tiz4TEMuzQ8OIv6Hr0/wz/yL7vcSkxvsWJX6WP
uzBQr3ndymzsiTs2S8MqDZ4YvUAaxQh0FcvTejN8zIuYXJkdFNqEJhyK4OjN70SB0aJ5jJansJ4/
WKCM8TAVOw3JIZTeBPTiI6iP7ApyXSZvs1W0aKcLiJ5twlFQzLyAkARVLhDL8ooZrmfYgPQSNg7B
GYdkPUm+aCEcMaTTKm0RoELYaNybi3mocEJtRaNNkxhKkmcFzvrB1KqZvv6T4ynnXXinDYg/sGS6
nDi/eYBMKVKVJMexgQHba4UetLOOjVhcPo3LguOWWfSNoCK9HzrHnJlw0nem9ubPV6t2VIjiT5pA
MpciOwLLoEAVkY7Kl4ETvE+Rpbv6G5pOa9bRx5uFeUQ9f1c4k9U+oxjR24bP/Ynv5BHD1kORiV5/
Wmufy1EC42XXX7Byin7jOuCTNha+p+RMfbFoY5sEg/eJ7UUuHf3MgfXUu03xYnBRQey5wtSqoFwF
JkqMf2eZgngb/mkF6lMCAXPJLg2rEivvOyZUHy9Efkyk9gEuR9BA4m8qp12o4yYdxa9RujhKvvRz
WOrC2ltf0ngJJEvVa0N6rctCKaFtA4+z5MOO5mQ5nM4UGzcwzS+9p8dJDs+ljVfD7ExL8bBUwupL
5rer1skOom+lMsPBBQiltDBf7fUSYqS+tYxmC6UvwbyFDlv+5myD2v40wh7GSjJUwNNiTs3P4psG
lU6Nw+ibn/qnk1tk0rnGaTyKx4pf7cWPwmHFeIC21d/9jpKSk5iZVTSckbZuKWf+hAc2Urs9/eeR
ggNMED0rPMNjlzrlbQfrRGObB6bO92Wpg+oV+XsVSlE3kjvEM35WaJ+uToc2nYbIEYnpyoPW2Aj3
TfbWm57DO4Ci080t+Dtxg3to8QtN9cMV1Nrnr9Z8YV0XlbPr0ToHvAdSW+IPuA5TAHG0Gl6PtEeX
f4kMEJ+UViaJFW3VEzX9c72heajXQ5c6XyrtmLwyMiQBgLGob9maHmJmBCj/hVelM29fZkqFikhl
nNT38RGsYmf9MxHl5pkKtagU76IS8DLd36FtzgLFA34UGfDw7UXjvlt0EbFH86wP4RZUL78fW6hm
jmbaJznV8rNyZrwXwCVqr1yCwvQlQqLOfOv5q+aM+Oakb55Akd+6Y4XLW5ZeiMDIz3zWYFBShbmG
Ltl9ORqXg6TVT9luj8XBGadQBkKpzM00kgLSL2FE4xcOshvzwcFjXjWRRlFc/y487VTECByHPLOj
LCi3vvb8q2ksJbeQj4OIawDeVABdwOsNUgHNkj21ObVslOL+ASygpd4yopFUBdRKGEvbl12xsxnF
4dZ8WdQUN/XLtiQlC+3uomP+Gcvwsi7oxuei3FhmSk2+/vOy2LZ3yZ/MRJ7uKqjC3108/ZYUjil+
mvxNTh9SsHuMWxmwiZaJ9NAFqvl8TTwXFET+JBBrT/WmLz8GqqL6/t7cBaQOdzqD5df0U53E0p0I
klybfVPjubquFz11ImazStUvMHsy7P1RDzrgWXGMcXUyLFvrB5rmJPbvtA/CtLFmzA7mw0kgo+cE
7H5H03r9kt4Hwu+PjRkPpEvQWGEqiJhIN1Gg2w0SyVDprg8nmFSggMwy01ONwcHVQdtbDVqNz2ze
FIlou/LvjwCo+MxdyVzEw1CGGphXGCf958J31fhzdekUjnNhx7D7f1FYKr8UsCxetB1rIxIdvcIh
BmYwtzuhI8q5peTL0jKBKP6tDVyCSvvTYjrj8DuT5Z/Y3eC8snljs0HMB3fXBhf5jaHv+4R+eXz2
blT1JB3OjCqo5uN2JsLJ34NfSHxvY39+QUAaFoVRBJmZMisONhIw7LF/SXPRae1jp5Nw5KZuTdu9
U1nH4kO/IsYmmfF7HudoZfK0VIOXIr2R1K6go4r4NaSCm9+C5aduDkrv6shZOSJyu5olhipM+pDt
eLLSgtmIZy1VyfvebcQM+wpGbfK5o934MRspZMMSYaOcaxf+Q6v4+nZnmF3wylnRuSubPZ6QGt8Q
SQvA+t2p7yVFzgrRZsmN7/OLxErXctiXm3HUJmRwjCSLSDOdEQa7AsLInyKYv+GuNGDlyLkdVCxj
I2IrXF2MNWrnjSIRN2taIdvce+JDn+cJYDfi/DfZ2rUoL7u0ZXdUePToAJyZh+yYVigHnDqPI4Zx
TCiCuigvtLHYsh7lvxpfI8Ilph5Jtj6Bf2WvQB6IDIlRJHjWZd+zXvqrS5nuoHla/SyajrdcI1kH
wSaPwLcAh5JbAxN958JGKWJfuPVKTDEBQcGFtYBd5TVRGdregcYP/0d0VE8jWPx0zGaVrdIU+fCS
WotJZG55gVLQ5TrohCLWHExDn/s/s0WszrrFpjGZ9IsTFAi+os+J07/VV6U0JrBywXl87ZKF+mwb
NqZnnxEQVyrtAr+jjjIEtLPrm4s8MgUGfKqk7mjvUyB7vkbTNFNhwJvOV8YyQK4YqRX9tGnYULU1
ZiHF/sWpAiqgWt86hQWZbhnnHctOOuEyH0WGY53sZHhBsE+A/1FcJLaCpg0DvTm5cT9Q5lQHFMj0
vSvXwyrF7T0/rQgmtrGu9E7P4UoONZnlQ5/OCVrgXtOuV19OFra8tleNwyqeqZRuJuUJXuj+kADJ
Ovgs0buH5vcRSekC1TM635vZVgWOKLyKSEdYSkF2O+McCpGL0EvXzkluZ2MTo5M3V/PoSmjh221V
D+t7nB1D8tWsRcK7MrFnsf4KrKAoSenrkeAEGtFJkZMjUR7ZljGtMZIw4xoHVnY37jG0qouslLPg
LAEaMU+wEK/x7atphmm7m85MmLRRTPk0h9lclvoqTXA4akyvAecmvqZUAMFpoouVdWVJL0NPFdAD
V4120lkhy5k4m0MgY4qbaKua6wZfprzwl5aFZzyf+TsPOmnBv/l6gx1fPNEQWEGfal5coFJfMw9F
qW9StUC9OJAFFDqbG31+LJT9t3L4r4+CzRk0gXNakPOfCgNDlzrCZ+youXh9pig4nNvZvBBr8dLu
A+OQnOaPUeMb/jwVyBMnDoOayffi4p9u5loZxTxa8lUWoJNsewyZ5TkxbvXDQ4VjEGFsMBvCsJk5
l3hZhwZtClGHN0SKNr76Wzu1v10yaddzyEL/lylDUFgmAsQzySxxL3vd77TlRYioKk6L08YVCVl4
pPmWK8nhaXmrAIhqSZ9FriMPTQjtc6FaMmpzEO8DZNO2PyPYtIlfvne+rypAj0AN8d8SU/9BqU77
l2Kjh3w8VHgp4rSUlvCu+yuatuOiZ5PdoRVwpUKLWaEk5jmc3SjVgw2/jJwXM7Zh3T5qRr9T3+ez
/bx6ccQy/dC6CKWNdVvIuT4zGI9g+JpTVDCPrN+PMxjQLigL2KeiHOH8jXZsM9v/iLAY9jM229xK
9VHazqo6fNGnhIObHaqEO9eF6JEhnBO/i0l85Ulzvqs2ZEX1Pe1ko9O11r8xp8iaLpfNLY4hrZtK
9e0auPFttJb8QLxATlFoicH7X9G0t8BXnxBGGzj5jASW4VBviFBQrYO0uN5cXb4K0hnJqy8CwSPH
bSkBynGRKBbLvN3RkZe3b5zz/cTzi+54/dF5t5yiy+XNeDbQaGpgL2Q1qXYcp7ECA63/e2qzwdQX
sspRpQ0qghJ0v2Lky2Je90Piuh9kPSPUFDsdK3C1maMGeZHoCin02/Wchtewti9Rj/WdovsrfkWU
KtgPGOmsoH29pWzWm4sZX8JC79vJhpZhgKXkDITSvflZl2BnZaWJD9f5VeIkjNmD+ZOUj42fYAxc
ljcojJ3ZznLh9AlyKZvkDrh+GzAyfmc0++8C5hy/h+/GiM7xTBAiuynE1FVn+IwJuAVP/WGX0ikR
zzIwVAsCmxe8MQrCYqQVQEbqzxZyOsnOZ3MFLHPIWH3GyRumUKMbkqSOh8Py0u//BwYsmTQux6dF
JDyjATOjshHqGWVjuLw6TNuQdXDiy5TYgPV7ng6WjeJdpn42VQl0AGt0ZIvqIUeWBWuifij5E6JG
ebICNq+TwIhp5HPhTbXyOxfcPG226dztb8VORFSuDZATbZrS3cf/3aSpIE7Imm/OI7gToMxVVweQ
19fT815SpNfsny/MHFGIqX6EQpr8U3TPu872HgbEt7pQRcwJS+CDSkEo/mqI+S/X+XRfAGiG0j35
qBCGch6LfJm+ItirhuaiFIn5iVXa202CQEmCJUnujvd0DUBHJ+RPsrLnlB8TqvcPskjJDczfW69s
JPu9xY/m6NBR92ENWQ0QCxNDtw1qISxY/Kue937tZSdu587s+p6YoWV78nvDSJLEGuPLrL9dYTnA
z1dAkTi9hD+2kN/LrL0LhF4AYIUulEI0jKQGYbqS8R00smzAmS1xPlycbzdLNWUlK2v2sUn9sfEm
BDdZbFDA8YOXu9s7nG5d591rFHA8uFMWDR5Ghzt1OgTBtWB0NfuiSwKLyA/1jiEEJ+B9T6P5zfup
+lYC0CdYy2Mr803ngagIf4Tob5XIsMSfKUNdSnnYo0hRNcnTP6FQi/3a77f6nP4PUzxeOuXYQOAN
EdXjcQcK4RGCzxluQLQamKymzL5BMCSMoIslypy/1qC3NTHeR36jfFHL998GlirMrgneet3abmO4
eGdJ9eVe2aKs8zWtyPjuNgOZwmLgfDbr/TWbuJEaa+Scmf7u60b0YepQlSl20BheuPnEQZ442pwc
3ZUmG8gi2yIzEn5wcjhspT8S4sc68L1/DFxk87XOFoRdqeluo4niGGT7xiWct4wmxueasRyiTP7i
us8uPXoEQsTHfigYaxAbos0KJAkGV1yiiqU+72/gzF2/R5sBgdKGPRZVMKIJ4yBvVq+nbaCSeLvU
BHFWl5wy+E+wR8Kg4qQsTtUno8ck1sfZIOpFlgrXPA2HQieyONuAWtteJ/iHWmXFSpeGSCGqP3fA
C6t2enwI12+Okiy+QaL7+JoE0UTfLig0iKNYnCNXnM3hwaBLHFopq1zpESNSNtqXNWEJ4H7LjFZs
vRgksPXUKEgbmcafGkUyfyDTW9qWA9WBQKR5VkEZ6k1onOV5KtM92JZYH4U07oGquX3Fi4fhGn+t
l/O04lTyo9yBKMZm293yYGcCOX52xrRmtjP35QrFlw4VVoq5oqSctFCKbaM79isNVfwVj/fiBXvK
aRHVXssEAVZdnLFjLAgmRE3QrIDonQf/aTn0oqm3cmWREUizOCUO63/QAMtX+Yb8om+zwcKvAHrC
1T28GY404AEePuMdjToWVA/eYu8e4NQCnWsWC+BFpdY2qavHnaWOe12moDHQVDdhkWfrHBERJk+j
Tk/lGLzfaQaM7Mveh8XRjfk3Go+FlPG3Vy1tyYRwtVIEIq7vo5tRfta4Lsw1aBsABWwrwrcNaIey
gs+XE8nl2B87TZhawF2Plgrv7SMuwPlOiAqtivd+IjqdoOfOl1X7VYVbM4ugIyf+Vs5FcUXhEdPy
pIb1OoL92IBzByfOIYU1mKzqOQQSgFKzHlazh1WCtPa4/VRgVAz4+z4sYtVDqKARVCKCqlJMM/Wp
A5ymiRg0aqtWFqci4PLIeSMBEkTSm1LdGKFi9gbzNqku9NNEyKka2TG64qPzMXF+tIou5SJlrDLx
hA5XgUdD8bEaNnM8ZO1S1fo2a1Agq7cAPcXYorqxjfnoEWoTU9pTRRH+1KWBD06fRMZVIHDmQ05W
4GejsUjG08NzUOPnd9GTeKHj6YzXGALaexOhMOYVrJREK2Tov+0RVyH4IahLweBmkVuCFltfAWEo
0bOT5oT4oUkbFYeXdjb7YrFwIWBhpnfMEFEEzzrnNuo2K8GdP4ZyNTFnBpmEafEUNnzG3TV1wOxP
uwPxWws7aLAls2J9FmFT6LGBjETaMLWR0ZvjRV9wl8y7/J5/WNi8oouwzLAMc4rgi0mAprWl/iDf
bRYoapWC0DBduxS8y8MbdFgnGfx3twx64Zk3Il4cYiq8WDOA7msdykpMJOSOmU1SblPNggtNZ4Aj
87c2vPDvV4TSKlvFjAVQBQt6qtrR6wqzHkuf+8y09NKkyQbxsQ4oNn5geR67jyJaNfEnVVIHRz4k
IpR331ZO+Wo6w/BTM0fi2UJptL6DNNosZttVWTDxEF/ThGb2pwDmbOpC4TTQ9WwxGyOUQ2oU2PCC
/zg6vBE8yXXrVVD7CiRw+A/6GJjLFtuJ8fNwSO9ih/pozXBJ6HgVRIETU+8oaBRP0CYE9gznBJee
sYbphzx+fYOQja7oWoXXheTOae48A5ilYeygSpQpbPRH9MwS331d2lKY5A1VnG3DV+s71+DeQnUE
C5BGT4RUJKSHxL/vQXcWrfsbxbSFgSSF8Ex5wDUpVg8AZOWFV4GoYfXoSV3OiGD3W5cQvMU84ls1
LPPQTgrVIYXgcxKrTpQFMlnRebD6JAIzkGaQlW9zmoSVTTZyxoS4p/UMwS827YOXb4qW9C2ZSuMQ
77lDZTZl7Xdd0UV+ePMHXPqahwFKnyuGFk1/xjXUz6Qb0383lUTTxiV7RvAZRmH25LxiC/ixLr7J
1BtoVR187/myUrPVT/N6hWf+8hZ6Tr0sK8zzw3UBW+tuHCg078Q6dDwBi/ZkQQ5PKodpymAEYDtB
rcWFSiI4Nwt8d/YXqYpfP7ekxEdAf3MuZ/RG+wKIek7K2Hs4TQ5pj5J8ZZFXFas4vT2xjOwYsD7Q
C14TjqT5zBKJOrTpRFyOEnAIIE+2ao+8wJjpwRlDedsOPG9X0v0AEJa1iEzk7PZ2dAZ4/TyILbEr
3cB0bCA83EqCDW6uKCZw/roEjxEPazxzN8i2ogUE2Uxo46KPJFYjWgpgGSESvn4W9OvZIvVNuMDb
MwcijM9y4PyyHYCvQeGt+urzeNe1BjMhkoz3OSgickYkcZ/sr/XGkF9o5HLin0cNmLqfz6gC2eQF
mpKBZ3yEWpW/VsLtFM4tC1FJgQ094foWNEvJiwt6/Wa+11ZqhFRWvpFNScqoeFQ1ByfXkdnrGWfy
kUZlYJX/AYT0xKClDu5NP66quIhyeYGn7idcPSYNkJ2ugyzuGY6G4qbO2LpQTT4qMcTotClfKjIc
CygIHbC++w5L2+fYbzsFlJyZuwM4BJYsaKjyLsbmgVV5cEEg+WBdvpeGxfSiELA1QMolvbYi+IFw
TG/KxOxVvDdcs5IZ/Hhy1g+8DCHvVB5fugbkHj0jPq1QEKPlVng4uQr+UC2DeDTWWMaaJ1RNqWu8
buLGNM3vjioyGY/vxtblPiFAET5lFwasJHuEXUlnhIR6UKoHH4qmx0aJkjms948TXpEny/g07mZw
lXrF0e1pr+Tzd/5f3VT5DZ/q30zrKWr8PBz7yRs8AN2uffu7dsn8ICSnsqgtfvBgQYjr+/57Fw+j
vthhR59JAbHUTP067uCQyRRmKrJKQn6ZAdkytA+wpB7AzfeAD/5VNp/IPfTrf6HkBBXxOn6sJHLW
Hmk4edVndBROdEsWrsElbrVkB8Y0l1U+D5QU0Elhe/BjdwKnhO2gPNDTRcTw5yPywTjWjeY8ftJR
WpRYff70QgCaFG6iKzkCO0TKl6q4BytR6E4PwjCuLo6TJmmpiskVVQzaOg4WRcMl0eOBFQNBMeMt
jZVGLnCSoYj2nrBkVzNE3pjJ1KN/iskXcgFCNN+gZ1XKYIY20On/hcPsJHdhopPyutzUNJyauaHy
PTavvpkfExJCbJIfbnwFGbj0qkykjyugt1DaAbLMbZPL5KBiIKtyh2NMR1Hnlofndn1NnyXc2/ie
i6iGkFaH5lGf5i88rY9tJ0p54uvA5mq+7a2uL0KH7LYLjKomsZvW3E7UFuZ9RM5CJA9WPSe5qrJq
M7gsrXtBojo9GBicBO+t4Ymgozaaj32xMxgik457IGeWRQCAtmAuCEiHNiefpzFLmSAROJG+uDvi
PWqFptqKFGZ3XyCbNDYF/yzs37/zqikJoyQD4UT384+KZZl9M4H8ZIa+QkBVpKRR4EJWxjxs1jhC
xMpXL+9oNnaCsl0GgW3L58Nav61j4Ij1Ew0h19nEOAqmPS7ohy+WHeAHVRFnxxBLUDJMSaOtW82Z
yW2plOcINsLeMWJhjvmjVAkk7qMnghAF8ZHl3OY0smZlJWP/KU8wgRGvVOt3Ixj7nGfMuKdSp4wa
yHLamx2ngCZ37SPqBeGI3SFgFfzRd5Nzwnd3cBNi8NRRgrIKW67uyiyX4DNPhxJ/4IR8fGBjLjSx
R6I/HbkFjnbXoiW7BXRD6cqRquZ2SDcz6zhdd6eh24tIX0DMev8KX/fR38xzW7F8PJHNX9oW2kdV
NG1nduu44hHkVJV9JIGI+ogq+CRWeHa/GFup0tysVon/lT2RtX4zv10VODgNgVjF1RwZi7d9fNmD
VgQ0+bEpMlvqZTTDpe9TJR10YRdA8mTFSwlABG+Ner0hCgaT7wVUgb0+U41QzsY4r8wdQU/VxMQ0
E/M8GA3vkIHm7poY6OlGWld7JKcvOrylVzB3fQdeThMU1dl4poT4wQEZixC5HnSjaeipSyFAKjiO
znH6OemSW+qhIAsZpr+2dkyPOLVzjxXfzDliPQD4IgnmFJXQ/SjccR3+iz+pE8Stokr9hapSCxPS
HASNCqKOmHhlDeJEnl7BVmWnVJuMMznohMRQ5XH3ntRsaQ/fn8+NmsIQi6WCUysQrOa64u1QBj4g
r24AYjfrEx7LQnMl3f1Okm8eVQaqApUElNZkyexb1PKpk6Es0gPp3d873DFRreV1ib/2qR49zCVH
3v4VHk6Z5INYbTxqAaAe/p3GaIPaG+4HWO5acjgFqPI/M228q3FZYfHtXACB4j2KrZkMTwNfssfW
cdv0srXcTtmHwZt7gDHh9/+SaCshWruChCT4opaXUVZvTqgpbUe7Ew1e95peVWowCLfpzvstFA4g
0Hi3ZcX3SD75AQ24Qhf2cTv6efyH/lOXyONPXYJ8lSNCpa2aEbmT1OZIjt0RupycOTdgxDPC8eMY
x4HMluz+O/FlTARcIaoamc5Wd4XzrnlRNt91tR/g1VgkqRXh3y9Yyq+z7WuzEedvIY3PB812MLhd
9OIA21cw1ei6+rxGd8xTsiElSYF6AXQAs2rfiEicuvYZNbu7ZELFyDeIai+dcnF9hUVkc+T199L0
2ZyyX/2wG/EKkcBJDka3wu94q2vbuv3WilxfsXxxn+Nr2Ag9jVtG5QHQYzjg9Q4Ov5L7H1fe1P+2
ttrtxqX3IHYYNkFWe+rIj1qQJwAuPAR6BHnO5WKab1x1CPWPGxKQMz30jxvo+jHKX0Nl5PrqNsbM
io/1bNW9Tv497jl9L036hEkYAcmudW1qTLm/pj+YOAXXw0JDUi2fmVfW8Cp6A71+drbYTJq8FIOx
Xz4hJURRxABkJVYA2IJkW08Up+uv0C484mndw6esP12c5jyqgMor0vfGo9juWyNoRmH3m9hxTjwD
TmiGo8CxyEVxdlQuHmowBKquK0PnyUoLf6mt0Rl4wae39zPUMhGKjBd7w0V46k4tYrVZCdr6PFqk
agpD36a4mdxezmd+aInk1DWYoy7ZBwyAz1S32SFkejvXyFZWykibut2ijYVSFHeahRSq0hm/jLcg
s63e6YTzmGyepjX8cBycJ1Ds+L20x2L/GC9fe1C79RNOKsVp/AqDRWnemC+0VLKTz4DbAURTG5Yi
+EuiqtVlwJMXv1tMeRvR4qHkiMY0yvgacl1+FhI9LM6XQpBucCcZsxFMlkCctMln1gliMkQyp+FW
+O+lde87njzrGuPOmtw6LcHiBm/1cKyBAkNash3NML2sNsSlUxaT64n+dmKSqs5SSE6BuQTY4e+W
356St140JYqTN9Lh5YBtdHXKAF3mZpUXpLsjHDxdu5CMDBmCDZqSKH+Iuzb5D8U3CRAQ2t9Qcss2
L0WeI5Txnm6m8YBHcbH8Z5JKwAX8syBMoHRTEJWlEnR5e/em2QmG7pkOMvF6FQRisEDOGib6mc6E
UiLkDFyg42Uk2AlEJIJNwvt5+OOcO4j61vmLGnaGv+1kc7ccW+EkW0xKylAcnmACcO5KBbkoUKTS
oIKyagjCrrfZWRB/uDY0bZggKl6GrhkEel/14Tz7roa8UzXztwZBTVYWqGj0R5ogYUp9nJgefvuE
+XEHezVm53AjILucQHNANyACx3l38dGT1pgaY5JJ6XNkfmFgUiq/ysI1QtqjsbIIoU+ELnVtKcuV
S0spQcnOo9Ls/OcQPgKhQOp1SpUAthYoRXrl89qalab/jncx6K8Np65TkMxyicVrSsKpZVSssjvb
ZhRZU2rQGLq8T3Mf1ehwYPtOApkXct7hSO2wJlNhnNOEw9xG/TrkZIYwdpD6ZD2In0qOZjhAsAOT
BW6vxfJQeGKiQtV8m6RP9xCG2xhT7KR9ZW6+usIsDYDNkKGX8/Lz+0Um74KTUg3mUGnf757sKKeB
ZB6zt5cQ1YPYbkYNscoyJk29v2aeKfVCgfdSyqDY1g0IismTRkS61oUd16fB9mkp+A7oJR4KSQbj
Go+YwOFndFrUOHwAjm8kYwMthWBySyt6WVSrW3D0/QhOlYhOev6UgP2bLWSAGwsi+OwSJIdw8vHt
QGTcHot2kwISp/NdVK9VAOBNTdhZmAp5xur379AAB7GD7sHcFgLuiQSpI62nPU3j50dW08M8UJ3A
ihHRti5eQ//V5Faq9mCc+5UGtM1MwwoIn+c9xjfDGBAzyRzOIZT7U1zyWA+Pn8UiXvBsp8FTiSyd
fm7q5NZvlMJ+jalxC6mB6PILR8jDYE8aIkEHYea7j/SPEiveEaONDoe0NjmuaCn2l5DT5UHTJn6v
MSoVys/mMc5nS9lzsvC0OzGFpO6VCAVlYGvtBlepOVRdD1Ieck27cHA/OBjwqWLJARslJvRVyII2
95GjxLFEenEvSBvg4trx8vvNsuMGdacQ7cgjJa5f0WpTDToZTxhiuzBzn5WfAkpsiKYFdpZ51cFP
SAnLe6sEoTJ/b6DUYsCoQoh73ErYulAeVS13jV3osB0jRoCv0NP2UBSfr6r26s286uek9kkZ4zvZ
onBQ7PeqbKPT2zp9b+6wwmJ2CPLL28jp5UJuU1IQh7umbVv76JERhHvU1L12O29lbpkcjN41fB+i
GAtZrbfXr92FySWyjfVC3p9uEvrmkUR/eE45ix1jbM5esAcwbjG9z0Wq9jVTn97NfDFwGuI58B30
4MmrGGtqQEMnjXBR2oahyNL324QR+YxZm9YhRRyn7XI5PpCMps/s1xW5aYvacQCPLjcyBuet0CIj
IXozyUCcjE3SxQ1qiNZwR5r8hL+0O2Yb88Kss0G1jkjWrSov2MDtAa6CTeS9VzpjvSor7x2XhPDG
S2fuvuQrh1hEABxTYHECNKJpm6CjW2HOoC5s0qDXK65dckUbY9WaOuz6mPzQiRHzEJhXy/b/AblJ
p6ZgjNTSvWmQyDsl35JFUk832qCxqU1xQQJHH3AY4GeXBZ9s2Wf9rFRhE48NJUEoeAZM8sA/Zrw/
SMoMmI8bGbzbGKAtt+xzDmVwgWfxLZx6+w43Es66engcWlPPtaQXD4a+5AkKbDcTW2onkHmNZqQn
4bxWsCHHfKjS1Mmzl7YT0UDHVfmyl5sDxAlc1gRSCLX8IYP28RWVHB3K3jBSsOp/BExsTY20p5ZW
7M6lHPA8xtjmhE14VnBZKHV2Q+r5Q85RhBKZkcnQJrviZHt20Dk4R1RlOGc4ymALzw2u/f7Wg5uT
Gf2lW3T5/yZ5VkA6CJ+TL07VARYXSmjOg3XwNXA08JDq7Qj+WBnxRfpvdkSSK8mG9bn4URxUq1ku
RC9rIVe1gWdDI2YJWMn72rfUJsXooQmQvyBS+dMh7Lq48dNu2xbo6+1IyFRfOycQq+eczEkzEOPV
PfL0wSLQ2T35VSwgCZNVjbZs0c8rW3TtEcNcb275nKJS3b+UdXPrhkmC2KIlk9f1qeGr4NIyVgnQ
kXfnvCWyNpiRuee23phstDRtpCxSYP5cSgpNhwNomVIAqiJrlLnVxDS9kg0lfhES/BtFS+dBKdQX
alAvOhJvEMgl2bJZ/j/XHFO1EL6XkVxtlj9F7RHc0XsPq8eTYlNhHbJrgvZqqtsjU6PVXkSrV4fc
0OKlGT1bozH0GwgDQ3qoBr5sMnfYR5qzb0mFxlALROFrmkory/eBfpqHG3LPVRkpy4npHFTnz02r
arGuRdz4CUDKEZvlLJDzu+HunybDdeqaMO2wnTaB0J9fP8Wkesggypie9WDyNN6vX2YWDKhMFn1O
dmst0hRcNu7GV5qogwli4JbH84TX9D2zvfMUMNtSxqAiwd5lzYku/Gibsos2l8uXkp3lHPy8aTRj
YeqtE6HxqHuvh29HDYCWWOj1hh66JZBJBmAdWxF8u+2c0b8zhgFseq4ggbm7fCYz6VOvnYGbiaN0
uPSh0Z9/Wc42rOG9hft70y9bqFiHV6+CVCDTVCMr0FKze7qXvI7U2e0w201QWdEwGvJita3jqGF6
GzQZOtuUimo1oqNGYebOLdoV34EE47u3Wb/gCQapwakolHyOiFPixaVubMqIGh0rjRbVr2LcVhto
19M8Ba050cV4j6W9soLLrmxgEuj+s9e5oIPT2VRr84rVPQv+KhNVWO7w0+JtKrcg80fH7oomRbNk
ofEtjM5WNb6Mi1ri6bVw8TxXqR6jfJ52YIzj2+UCOwvLTxneX2oTOF9sQ54whtBf2yYht8G1gl1Y
t87uj1MkNmwbEoDLtC97WfOWKgYsLgRgF0F2V4AS/uXTigSqkjPNyL9IbTCBdlM25afi7AyECm9I
9h7vlXORAHSZ9fFtPtX03QyXHUDhsyYbp9R9BhocmjYJ9VNJyjF/b1iFfwEnhjLfX35YIgiPm4ur
snGMHfwxAcj3jRW3btIQWbnKJyRk1R2kQWktExtRhQQu8b2z2pcq7+0ZGE8KBDadrJlPytBa2p7p
/lOB+CobSFX19fVIsn/xU+KkyGdR81RPIguDXdO/kpKifNCTJ5sCb7BFhYLSlyw7u0/SfD91KsHG
2+wyxspeb9iCR0iUZHAKLBTeTW1dCVOitwXLyAYC35ktX7IExu38NvJTW9TOOXCEMBbOKVkKZlY0
GwPv7qygAKl49PmemQggNC4zu4U1lPf1Ma4+HMxSTG8T8d460YwW/Rd3XB9+PB7iZjWJ6OFstNMe
GApMahrLbmokSM1ki/aciKTVf2tOPHXBskd0x1OK56Kfs+hHq7WrXRu3+zZIsXKiVkiOBw5p279W
+oWz6/+sMm2IYPU4pEwPqWMzP/ewMHi9QANx09px/aMMOGzlUYZ8TPfDQciwS8AwjuAAFJGA6t2Q
o23zy3i5EN5LBGcTvw2iBmLUfmNHbNrmtW3b9m0Sjx/YxhtcJAQAGVZjtKYa/+MQgnMdWCm7mJeg
oFw5aHllgwHrt0jclLYFE7UGCI1kBrsPlWQNKP50fnQquEyacQcSCxI4garGtpMB3UwC48VIaatZ
YUjMPAFZfhLYLXPUDF3Y/lV3GIC92R2V8k2dVsz5TOeFykHLpN/CDTqJco/vyN/7xM0EQbGHLA4X
iatuY6ljAbjz7eypO1ux8zSuDq2ARvi9PJHmMu9QxAe2zkKWt235dxZ6FbJ34HgmnxnrPVMY3JT1
745XB+keHXSAD515fgeQDQymdXFtMw9t1Fh9JBPz41saKkPayV1T2cr8EY4DUyQW+Pa9gSJCVPGs
rKPic65IbPyOPTHz4H+caQ08h6pP1VEEVkqtwdPEuWGIPWOxJetenimaZIIPEf6pd4JaTZaIsmzR
CxE2hLt9ko1H2NqrQOIRrtCz3JRrPuFZcHdKi0oqpCeRPlBOOAj2rU3Uwv+DwKohIUMauZsTK+NE
Ip0676PUoqVeDbL//7FEqT7sW0dSguX+HklqGCvAsmx3juWOOLFziBT0aVXu1/2MpaGeYKjRx42l
jTCW5h0coOTQrw+Ix1uC/mApESbYwflmR3YnFZaKaKh7J0zt0P7qGZhgXG8j0ZoenNl3oQIYZnl6
SQj0tayiig1BTrYdW8Fr2kyZZlekSwNRpj4j/Jvfr4U7XlZ2uf1pCb+tyFwbECOCwAbJeR2kVtQv
2QmGL4p70oESEx5Q4altg5zOqcMOurcCnvjwGdVBgGTkP4wHqox5e2mNFrimo8iT2NRPkfcxTim3
GXWbhrPtN9ihrOce9naxS3nSR91KKJr7WpG2pzcwTE1BaAIyCkeSFGnSdPJlkRdI8ULPmMss9CPz
+OEI/Yemj9sbGZ8DlsIGqJcVbOugTb+Gpl2IJAVm5KmP7nG0FNzs0sUHqy+uxEVpoj7tOawzjA8h
ulIVBHjP10a0rExfAOhqqKEM3XzTL5TlSCW187Lfb6bM+ROMCTUCK7AvpUVTJB997EhFE7fG64Qe
CLMSrzYdB0DOC/ZM5ChMeR0KRtegMhdbd6sJRw6/TwZllWgJGFoks6538lGBpjCkNRdp12TRt1rq
0qSZCaDGvKmz/NYVPXM5hiO/cz1CMDkVlinVQgT4EVVz/vQ4egKazMY3saKws8PcX0QDlS/UddLv
DI0tzIbSyVn8QqXaC72roeeCuAB/p3FiSHdYThIo7CMe1axWEKljcmb3lUirJE9xMXM5eNNbFq0Z
TeQZw23iYOL3LRWPnugVthb6SD+MQe5+VqVafsHRKMdeq6clPmIQe8JUBbSl5YSMfrjuAKhF654k
UtpX5XYjjoa0nUzTnXerhcl2CPJci0bau7L9FUMaTIKtQlzZGc9eLLioVETLzgFSlD0RQofmc8E/
VvzPWovmmFcC9I/qISIJWmSJbKFTIUnOO4Nr/YEzjAxIqbIhS9tBjNEGf7uvySheysJL0E46y469
HP1zILdeFxGj/ATA8n1EUOKuV9G2JFWL2dSNLY/Gbpf5pCGWub0xAMLOeZO71EK8Zvuf6v03WE5N
yrzG3OyRmQsbzQq7yYkc5hX9YHQk0CqyacdnfVFl6gKV/QLgo8M4ghurnhr3KrzB+r3YXXexvQ17
uW8OHeKnR8VLuPrw1PFremN2o2NiCn2zGbPUj6Yau71M//IDwd4fghDqDhBFzlENDbeYEGejnWyU
mb41s7MaYHMSYeWvrRfdC/P0G3FY995BcBumIxmv9zUYZvAm9DkewyM4HG/gnDZORPiZn/Az6+HP
dfHa/f4CK5GY+C8bTSfjZYYGfCa/pDDjMKnqa5ZZ4hKp3lXlkhIAQm3Zmw2FqrOvdBRjLnCALGaK
DNSj6pzR/mH8mGYiOUa7aEiRIPXaKlC5kM0KvAzFVnrY38tLCHPoPFCMTS4+mywFAM9LqyHJ0d98
M25u06rm+ez+LqW3+fdk4MvWaoFB5W2v6oF3tC4gtyH7PUOicxYeDB9PHcRmWPYnbhyF8HTULYqp
QaB/ukUe2yv6DV6NyVJPT5JTfFAXxviRsXdMJ5BYXghrfAcnqPlGNsTIgH55Qz2IVDJeXlTVU6H4
4PDABIItwVecGfPffPONt09oqOPMuezPg4CyPIhGeGOYmH96U2xS9Fyhk4EgxnFoBBR5p6CptB+W
zufVyXltkPh9FOKq5x3P0SCXxTvARxl6NpwNBHmT6e7nW1bB4VqUHfCxb890sY9fNkPld/XBAmFR
mHAu63Otir6yl6ahC/PiK4Gwd4gB22Ebq9JT2mo37gywJM9ovh5X54fLXAaEQop5xaDWM3Rmd9yx
TPA1eCWBG50OI1eq7YCH8nsXeyUARNG+v1ecxFw8pr3IcBMDZsxZDw6i09z0Suodwscs9mOhFOmy
dJuvEVixof4YtFzQ5uCc0GVk7tbzVdzSm0FWv2Yv2KlOsV9vN+UYhTdcrfJC96N8EbmI89J8kAXx
LRjKgH/Dpy0zMgW6UKCvnq9D8oJsbLvoFr5rbP2CAhOmJ5uiShU1IuMilw53zFrOrMqp15P5bog5
mux1IGR04PWNhBCUE5D0J3l9QA7wen20D+xFxBYMHiaa7o71hC/fQj7XZ3XXifTOhyujQmkZkQKH
W9SLSpWz9Y8DDx/SD09w23eGE3IOanH3yf+jvrI7LBv4eytW7f/DtVky6ob2IVLrHkt7H9xY1JAv
n7aaiEOAgoiMaiG5H20uBck1ZzhhSE8cgpjZQYktEYoTAXT2XbZt/JH5SMhMGn9J+8rvfQG1bH5L
SNVA9ZfJZvq64Y6U48Mg1ZpSKpkwJfiihTwC9qy9HvVglXO30utzbAB+65Bkix9XeHJ6DVOlWWQo
hTQx07Rt6KlyUQaoAMbJMePdkMUyu43SPN2cA02KR+dsdkpyJT3DHMfZEzwv5f7yE1FBaIR+tfaG
fd7yilwHc+rG72/ydCHgz/+8IPul+DJLXfHaUjCqtuZ7FCpH+k1CNAjZf7pKVCl4HCJ+nJWpIuYL
lapzWx9oGdTGSzHOiTpFKe1SEdhI22yZ+nS2SRNb1OL59Nf4E0q43KHqZS72YQzzHW1j+VnpKQls
1VFnM+mNycridd4p/MrDLQ8b0OqelBZrUqdxIvIJn0h9ugAbPWRFcNZOJVRkB3MGZKhAkhuKCoWB
+U6Gxh++Zq5b/sffOSJhT2Rj2zLbSmrsdGXQwYw6o0apXhobI838KF+sljm1/etwddrZXURu4nVv
YZ5IttQbqBqNsmMyXAYLNX+CKH/CZX5T8S1ffKeX0Zp8fFFYs65UXRVpfZmx5VooY6KxgNreNHag
NXzZ6571Yz2OhopQ99LiOt426jSBJbuatPDy7pEvWtp6WC1W9186Z7CcawQx1L3ZLEQHa2AfpCtF
TeyAKA/DGQwzwgMHwf0BPxrsJ8YyBZvLfWcWpKu9I8QEP3dj7+K2hiqHsB70J058hIyjtLPEF/Pm
49Adpfa4bO2xtqBDD8kSrxOY2amhnQw6+ftxVQ/2huzENM/Yw+OY7aqZK7IH5T9BQzaIQaHtC6ve
Wav319hw+0UhB5KNhNCSFhmC2nvif/R8nLxMpjfCe3tXOGDttdfRzTSgZCUq15pYm/BYYr46Sg2a
3lWU0yhVI2CSlsCMPs6o/RLHw5PUgiFSJLK6Lof+/8/12yQ0PTWKpgKAVc1jqEMSw43Fsg8LW1uv
/NqtEnBNUOsw/4OFAx7U3hbbvf6/INy+moT4CnfG966wZEbmH0ETzYzGq4sd6M+0MQ4J6qIRB5Ax
f63SNp1gdiWNxTY07A8cnjVnOqjCsAHhtk2K+yxUNUUH2Nd7UcRLW2VTLE1nb7YXBLAwdZfxi0W2
VoMaFu2AAOUDZm+FdQ1WxoexKjGi8JNmPGIpR+HNahOW5IsvBBGlo8Ao0y5tZBPSotSjMcTy7bI+
FQekcrUx2TLzlpKi7MQ3HP3Etu8DneMhivZuY0GJAG/7tJB/Mta383WvyNSIsMkiadZWQRPqODG9
fLId4qLnS9pre+rjrKPYEuxtitrI3/iaW11iH9y96MxwAFywHq1kybff4bYukvU3amrPQt3s892n
XqiCR+4+G0ly5t6XUAHkWhc+L1gI55E9yKCclr8GToxKCCJULg42h2tLf7dmI6AQzz4R8CmrzbEM
1qrTs16GHchLYBYibn4gUEwM7+xgjZAgVdCQRhOCNUbSGIsdn4W2IJSRzrLPtEZKmMAyWkBNvChT
ZeAR/2nV5jKUGl9Cv8Ep8aRgmtoexBjuJook3l2PoBnN/qHEzSMc9XF+VZT8umrESOJTnxcipw07
AACZvmS7jJZR+ntWkOvi/XZc3SH+wz1cly3CEtLbW0goxQnISCindZ3OZ+jIHivNplIwaLWQTTrr
+SbmE5Sc8wkgX8soVWQMQDuqfU0ChzTa9t7zsVtwR+l4X+OYqTdQHJXWqClzCzFuJspIq132Eeya
VokSZHlwi+wD6fS3pWnanCoZ+q+JAARXmrCBN1uhJL28BzsM9qDhpyILLqW1NQSJwtRukGB8Dy0+
z4hTsXcXvHvAuUKrI/2ujQ4J1YJOY8jZuqQF5evI6Iq65/hFKK4Ei3Z0dNzRQU9dxnMwtWMGWkTw
6MqvRVfUJ9lewM4P/k5CUj5xGMlSNqErkUejlFgjswJwTZJHsWp8RnTxV5mtVYKkmdbh8lwhEi7d
tMFCX6cLHQPRByBlKEJLSiN05tSeYqLj0itI8UTIToVAGjmaQ+jpMr+BcwH03yJY4MTIP3ZeqjFn
9nGuqHbE17X0CR3mo4qFlpGO3OSXpcjfleIpnScm7sV0J0KXzhbN+SGBQzSqcn31d1VyvdG9hqpO
MbxmpcXBtlfjoCn09yoGoLJT+r+r3gKcIyEwkM9aT1SMygGEMDcipG5J5vlVsf1vLIMqG4WqIBrm
Hn+1O4RYfEy38nVxUq3FAMgtDHNReLKFGUt2Td7MwysuPaqbeSuXr9kmHu8Rt/PZJgEYSHPztwpZ
mkx4jozF+YoG3j1/ULQCp3hn/Hj5qwvzctWwV9K9lsdII3f4kR2vVaXxLvYutFwNt2neWjczudbF
t3or26vQ/PUu4N/xorxq2Qecib0Gi8bMiWeJK1ZhhZXuSWWDIXww8AJTbh97apNqMusTuTtv2nSQ
X31Ro3v9W9JgK7KnDAXNgJDb1A6zx6knwZlUqqPUNTepHQPNfubWuce8/JdhnXaGnl4mtkQn/v7r
mC6/ktDl7cH1xRct6q6R33becJaocGD9PcqYGBFVwVjOHFlm9VPrTFSbLvT1od0DXKP2/zJoanpU
TL7q5sEnyEHVw9eEEWEmW0JxXlChZzkz+q5n/AI2R7qgxX1nZbtM8+tGn7m75HR7xyyUlW57Wxwd
E2YE8G0/4Ztw6gKI6tp1FULkcUgtjcVcUufB+wU5QYfGcQahCEW6ruZFOi7Ek4myk0GPDeHICUmM
XwQ/FdTKbMo3StaDvuSthN9dYKm+tJ7GAjjnS8ZBHemDkOx/YxmVaXR0XMHi86Pu2EmPWHfzuIxK
XgXujySMJaSre7oYJR1MGcxYk/wwOE7zuH39p+ktcTh0DE/eUd719YNCY3fri3aa9EZjeflsFYrD
e9kRi0tSM/0SAtQTuO0fHPQr6LhyK+4aSMi3K7zlZfU21Cz7IuSUNPX9xhO+XgGaaxyBoI/7UZTf
CCXhi1G0zaj0jwLkRPPQCM1xdpJ4euX3/FX+XCOQLWzQHT94vJzPau3B63BLns1NkHRQBXyM5yU5
a4FlytJuszdt08Fs2JipLG8OTYFajb13Ti+WMXfSMP8+/vmC1H+sJkaxSDYc9jWEjpF2g1O9R0O6
4R40TlcTthNjxaCfgjYh7ySY17mbG7ObgmflYRliLfz6bDNeJ9Skycb2v5nMffb90AwcglO77fl0
/3NiR9oqPH9/bOaSuChtUjL+w/0VXYtGOtqPpx97NIY7We9oyZpP6AsKVWnKTX2oYyXU5E73otB8
Cz7AVDPwKUY2/c4yBHo3ZTCUMs6JSeC/B9X4i46BpjfzmnlY78YJw/dlUmOi0WNHKJiiFFpF61Hd
mS17paAfgvAh2ESGiWz95bBi0wqtnZmE3lOZSZedKQJpcxbiw3ui96x95sFi6/EsL7IaxRdKP0UA
Z75csw+vke7UlOGT7zoNUDdsCNrr/1j8ZHysd11WeePVufXhJ3X/aiI2+iG9/0uutxs0sJUN4GAL
o3XP5DQCkB4cVO6rRPDIj67FHsUfF1jGeoKun4KxYsg0xaHU8Z3hXwO0c9XR49glWKWsbGVv143N
UtEaZfdyb9/j5FbFgSOLP6hvpo1P4pr1gRx9VErsSbov1sU1rkkpLyKUza+KRTd+cgyrMVD3R8j2
l1GIWqKNFb1r61rbBiFxl2lsPg2F/25tMqU7oK1mW3z6K1p4QLyJ1OXqB7a/kDauQvrt4dScCcKI
F+Cfeb6DTUBRxiGrc8wgAOD/VX0zklgHoTn7vDTphAK7zVEAAZdCSaoRmqZP1r7WW/g84hgu8Wan
kAfpbq6LVTfTBlLsoi0EZtCJwJAc/QrYIuiXJECAlae4d8qWGy8YrjPwjzyoqV4lz+2nDwZcwSx2
o1FkcUgyzuHUCDkDj4I2oqXzjOFggjefbumpRu1oklMO0rxeqimMqFtMBX8tunwgkN9jAqBpml8s
cUwc2Mwi8hruP1xdYh4m6q6fw7qJNtkpto+5fxtV2HF+AIsPfZccyG+O6C45SJ5E0JHb8pz8WvsS
QIDazsEqtBXRL76NuMwsVwcsHLsDmMdmmILYTClVn2upEnGkF5f0Um1h9k86fze6OZD2ZmQiF5j1
0eHUyQ6rTjPhQfZNUF9IsnD2ZsXIJoW2pA/+2DIc6mSAl1Vgb06UIt7GCgI14g0tJozqWsXcUBHp
+7xjxKTJEQHH4G4u40MNRhQhFOmRbKDnKJk2sPEAzua+H3UtC9u5ebRgZ+f/qQYiqxHGDGJag3gX
b8VJkNy0I9ruK4yxoRwAElrwpZ3kfXHn/S+OJajqHXklTB9KwTRh/vJkY0mllSfXz8MApE5edzog
gz+pPX1vAAK2x6DYgy3QMyRAF1BOkdLjmH2hQNpb6DURWBxPUVkRTiNP3yXQIlaU1tWL9hoZEJ5m
xhNVZPh4CAiyVujlA1pmsRmPvfFxvYxREp00DhDemwpw36lZ142cuQRWjeyJRUPP5fexx3mivw5A
1WcHXuP2oDAoGiGifnAD63tGOtwoqxxXxhSbWa0xHPipFvVTU3kgK+xmZSdZy09H0psohS9Bs0s2
iTV9TuFx0hRlQrsafmdMKqArta8sjUCe2uk5I2h6RKNHAQQNGkgULT/QW4ZZM3Hvcx3F4XasTWrm
b+QzxCmNy0rAc9FbS66QZk0JLWq3Y5WB9Ew2XPtmom8QXV60SXpV7cr12yAgrAGsEkp/a6MZMRW5
gZUF20KKq6HbMV3DduE43Qrz7ewdwRrCLtr0W17LSwDjQ6GP+j5mKEC/XJ8VPSBYePBD/Wlikhcc
nOrv6DvqlWxGv+ev0W/lDNBMtLZlwqYNvshCtEhzVDQvFcf0oErZM/j/2K+pFzWZibHvonKxCbUw
p+tDHLSyJ0y1vCT+ccIs1PrgD/BhCnQzpcqRBqTmkYRp/Sc5rJnPqNYGT+1QIFf57rPH3m+EjkAF
rTXo+JG/PVeIThhIrEy7XPkxOWOycIuB43iDY/jbgiRNDcCFQ2X63TRl/b8y/rkufKe8fjs5FDoO
WHtUl2PHXMrBPfVy5eJr844H13wyUn7Nywvtl4DFALl0yJv1AJvCNWwIWE9JCNgsvDfTDFzDHdgj
gtO4EUWe6fADnwheDnV+TZkT9udZTVY7SCtvA1t3GqDkmIOngX/IcBeq9U2TutVPsEJow+ChO9gA
kw6hQ5ymlAqKcbNpe0oHepRb9CfMvluo252P3tcjG8CUv7c1YQkfK3GSeFQ7CJi/t+vapyXpogN6
lDr9K+iMvqp+ncqAsK7gBY7hHp1aplD6p+jmJjj4HKMnEkwIQhEoB+CRZXZaXaaMLRcgukYIakvg
aySqmwBwFPnmManEF4z18IkH1YkP7CtX/JrAxc9kWpZsS3kC9DwhAUrQa4OEArCEeTJpb+HFY7DO
ZBnjD44YBzWxMSdhi566TCesDPkyuguV6A5HfdeysrExpCOC7R0FhTJMqLmU5qvbuO8kwTGmpK5E
wtYFBXlCfQi3CR138YKVDslqh0xNq5y0lOzVmfUXMeFeGpofkz1giGNG+jeBompp6aYuHpoGIoHA
9LigjIuMqD6TL+M3IJoLE+aseK4AnfF3+kXhq9KeTX2lIJWecY/O4CtWvRHugwfzNC6zl2J+TIb6
PhFpfN+khpAw/pinNiakHEfyCf/qpee2Hl2hZPDQb+Iu+y8uoSzGm8bGMrIVM2HW93irr6MhxvTI
JEI1wtTEIwsyK6TdJL2/VMJYYxIfp1OvbcD1/FANtDxFK+lNMlNJc1qPy97GV50GoS/NWiXBX4c+
qahgUf+8yHCVeVtg/5Bs4P47BAOlUHiSnsxcj+pI8n8p77kvg3HM9hSw9wooSMkHfMnZV12Qurkl
Ets2f+FL5TF0D6WBR+06d6/q0VswSIL4vy+v+oXZ/jUDTyCA1orbwOOEeRxnavxRDeQ+sEGbs1a2
/cqJ4WTVEdxrAxQjXMQ15aOZEA8g2IOtWLgTXl2zJKUpBiem+EpDYwzMdzP/5Z7RohKe7Bily79v
jZ7Wmy0MbPz4DlWIYvTG2VezYCHQdz9+wd8+EEgoNq863w6+k7ZNod01zlT62AIAYvqIdszxK3B+
4rf8Z1KF980llJNZuZU2rsiKRh18wfOJ5HRiBS1PIshRJlVJegV2KNbnXT2WR5p1buwcGp6adz0e
XyJPuh4Xm9i25TUC4hyY6aS3i9PDwMm7vdBvAEQ/6zBiq/edkly+a5H0i2rMAmjdouYy4VVaoEfR
tvXPGihOZBbGBWcOU+Qzb9kXeTyQp7SC2d9LZFjVObUgKzYteISOL8+obmTIXhmOhqpKU9bJwKG5
SSwdyL77RiUDTpQQuz0QyNTc5C8cLw7jejPSVrfOE5NIXM1K6dqtvwkd+skYrWc0QY1aKLoEhpA8
ZgOt3eUr0jRdy3/LU7YTWnTA/Q+a2ldmK1tZ+2+EhpdYgmQBVc5ocJmO3H5LY0F4XACvI1SERw43
oe80ZFtOt6qje6J4z22mTgpznbmpTf47qvNQ4+406DNeK1vyoU5DmdjhnzklRb7YCvn0i0fkaGc5
iZRGwF58ZoQ97T1NFpKEjsnR1wikMiz1cu0zyz0bhEGpmKAjGb1xM0IIyRy+WC7azzKhyOjzd0jk
HIYVkH49Ajvrp2E7JjT2kJf19NwhR4I/gxa9ESFeumLm5xOUq8J3KlAAq1BOqebSBfTGrC2sGAoT
oBZ+vI7kOy7c9t19tLbiLcFR6Xl+NzH07eRi7ebh1y3SOq34ZGiFjB4/aQMrmmIsuH3wJkqTp8Ty
0XzTr7hSAzvpGdq5SV2mwBFGf5oJs1HXDeOlRpHLO5EWEYHcGySHc5sKf6c57+bmi8nslV2h1lXw
6pQcB3dK0hPy5teJY5d1CVZkOGjHhqLquli/7dE3pmp0bUyAwt58TYQsTiLAsJMGsCUuZfbGj9WZ
CoT6yAATgB3bSIC2k/lM3H76/hq0hM9VyRMzDHFDxHumtnnHrZuClrrq/v9P7l3v1E5mDTiBBb35
w2m907jgvQ3zoqs+rY+3FkkHhODKjCvviiXOM5J17Z2YcMQJ68+FKyGqu6xbJSJOJ1UZ0NNwoRqt
as7qijuH0Yyz/qNkIB8+VsWAQeqLo/azQ7KCWYOipWsbv7/HI05EDK9OC7zfXq2rUNkVyCzDeQt9
ab+7iwQCG+xW+Hm95F7Wo5eyecd4jSQuekpRxd7gHr8QAXR+0hi6wsdfCKW4Mckp4gxlokoaRh4f
xLo4rkRjhCA/nRSs3uUOGmTOab8IZpYNcCNBlJqTVzUbmk923vHHL3MxN1wYNdYMuzOgB3joCFy9
7m2qvUUANOh298HnZRcczN1BGFxI/l/BvP5dCDx2dkY7g9HIgnRjgm3jU6sTl4dH5IAuNsscIYNb
nDHkAZFLStMIGzNqMOzr91sHROB6Lz9cyl8MQtaBhPE8l9FXdsczTrqoHTDallZLse0xrVeVKpvF
NWH1oPha8pHPfR7bJC6aDWoWkYVHrQPUjliv3vDXdIAyPGTbJBeQX2oWBL5YpTyH90PDa0zfAD9s
LlmvuLsmajrBpr2jG7XylLUC2+n/lP3CUirycfyOw1sn+466IQzw4u6B94ZwaW1Z3wjgovWUs0hW
ldQM6I071PZ5DzhJEIxHvrn8ZBx6uOPMfxAclXvBd8DVPq0lz9Bgg5Nbkl5uruScgvsQ4ygZ0Nhi
t0/rmaI4N+F+2im2gP30QcicH8R1cuch7an1dz/XaITYGj5DnKGG/6QMk3yNrnH/hZtTHzUPjbF4
7QB59//okfJh/y6Wxl3QraSVPpv5OAScjBnEUAswz0N6V9M0PaEu5RqqI2EIz6C9oIMqr085r2D0
eI5v56M/jrEgrsz10KyFT/xQDxJQjCU9mugMS9PCKDEPsYf+jNAUfKxh2Nqe1G4Qc3H3mi0erGKi
OP7YADOSnlc+vf9e737RZa5wkSpwGzHsxrql+5v6hUmXx8n+xMdrllA+oYCOrVnXi7A5AXC+kQAT
B0eXub7PzI/+tkIBlIJndUc7vjoUFOa0PLU/5o/xgpOoSSvYCWAD/xierBVicPFgx8L8yD8lofzO
amLnAKe2J36sGZLL0bG3GJTaqkWiKt0jkbLqK9XZ7lxvF9NMAMmkZZdcaHRX64GoHnaPrP3uXhnV
x4ruhtuPEhajtz9HPCxGMb0LWEBAI8qYGuxR8tNgSP8SMnyKqw7lygxC5q8Izy3OxRzsh2M8XOcM
ZBBMj9Iqv3QbWVNQGl9OiZ5FuuhbdT1eYSnzOwmhr73vrQWSuP7GGaUh1KaC+x5FdN7byTqsVPSk
S05hoha0W8nMwGLLlLNdciuECd1yJfjuoio3umufkA0Oy4BPhpul/y8zm5T1rT0TrVNfSS1iuu1t
R0tiyVzwOOjrAQFC3H3n9c/KAEvlslKJHTVgO1oi61zmqqedeg9w0Zdl55sFuBzZhKeqVNMzO0//
uyv1b5hVucFqCLOKek8V6rs2RSpWQs4meHAKtc5osjWN7z7DY/2tWlPod7j4buTPYCvbFRKECusZ
DSJNWDWBWvuBiZSqba8vQ++UervEvHlsHfiDSFbCAqGV+c7OvTPbKeOfqHNdMA6eqrKgR3lx0qbe
DfZtf70Y/ITWqiWV3q6qOJehh7zMyq8ngcXr6AgorcXT9vZIa3B4UIwpDALqj3HjdLGNi2AtQEHB
FGvYQlAX2zKsVXcc4M8ZN6LuZkq7jIQQYdjJOhMIW0hiRSoDNERHwLOCJsz7mepqPRGO8tlrbPWx
aAXB8e3MMtjzMdHLmbEABLVTRtR3ItNJLT/WIE2LgmQ5NK0EfP9oIGrJbZ0MOQJtcVvsQWxFhz5E
QplFx9GZGEaWGYtUcrZiupN9PSLMF1zDQ7HWsed8XX+JMJNbXYTM6WRcqCuVZv5sMliu/CW2b7Sg
9XBVYutl00fEDwXKYhZxkU0fDLLfP4Z6IDRReYHA2f60HEAwOV7RM0XC1uE2BpPAk8MymBlAPEDo
xhLaM0WpiwFl+LcDAp02ZiOlWQwrIeFDbWwVQZg1u3j+p8cdP3KxcOkIHVIsWeXHVoUSrPRO6vwA
o8hD5oH7BgJSAFy8s67xH26YbEwiEvrE1siKY90qtgjYREWA5CBhFgFx4VV/YvIJuG3/G1W9X5Xz
xlHEduSvb2iAEotUREI1hyecWd9KITHb2IHgkPB/alOLLer4syHx0Fa9TCU93+NFztWpQmaUuW3k
BV0HdfsFN+GAWhguCoGsv7S5miaW/iP+IQ+yUG0SQZuks86vTZOYO5Qak0Nw1n1PzNdYNyZ/hvli
KbFmF1wHdTcBlRUQlKMIiiyzuV8C6NIr2B2Z5/H8HsIF8mXU8nQ7ScNngBoSwEWzpD7EFc29QNj+
zqfWt5AWNXjh6CTiPvWD4plJasJ5KjgpT6FMWnsMBfeEczPsbu5LSWWqC19Ib9iqOObCim5Ws3uM
1cWEFqXlZJTo1Xz1UIr2i1nNGECM8ZE0esi0B+8n7uxe2Yg0I3XnctQdcopn6wr22d5mu8UFVLMd
/PrDIAC96+XLp/2iQRlvQ236ZBFpnqjOTv8o6xZiW+iiGLa+g/pMZRKRqH873VxaNPu6Z/7Q3vH7
b61ZfyXbbj0D6JIPKfbcm7BN7qMsQBZOb3sTuNmlLNO0F7zqV649SYKTUtk6B934fPJMDG77NZND
juj5Dl+r222SxTUxdUyAvTrYDngU5OuttDiro4HR00yZl3NJ80lgVHTCctbm2SDd/Ibo6tLXPn30
6rEh7W9IxBKZO8fikQt+yGcPPeOXG2r1AHBZoWBwmDoqRRK0IbpPCMIaujTiVOGrjdFHQFX47Kp7
aDaR25PMLvFLe02T+WdX3or61GaC7YC5wJz7v6/sXo/ksHoA6/UXI9JeiTwzrt1N3InF5BYFixUk
a3hJp9YXYtk2xFqUvclghUHF7xkzYqEzwars5xe+RoMPfKnOZkmuO16UqTVrqo93Ih2P9KMg2/AE
iRkQM+udy3k4NKmGpDkUWsUlj7K6QrS+0NAN2YTdGYfAbM+8SXoFdaKxW4i4adaJJFA1z9VzMU8M
LpM1UoXeB4Gk2M806YVzlifOVr/fAaD2sIOgHYFIjF5DrwqZRqSAp9bO+EsDKebI+SY+Wbegp2/M
4whc7yEB/Y47wWn7uzp/G+OHk0sabrbYklJayd/WIGtxKt5Ma7O+d+qKxqzsLfvMpaol3OnVBwXS
8PtOszZ381P3jsUxt9h+oOeKXuzRYvLkBUuE/WGzDhWQx+y22dSkAFVzYFXS0xdHf71Uki1OWOmJ
8AaUyLHfrIPT/xsTqgvo3ogRO1AG/E8ETJY6uiHn9ReiBtSaQ6Hkn6BRleU4QVDjx5OQmxJgNev3
ga60n3Xo8xq+3m0W6TN/L4TgxI0g5zo4g7Z7hXT/E7jVUlGNlzvYgXVVBeBIwIPjyFe3hosQ7Bou
4FYoYZHH8/sU+80Wqj/BoRaN926f5MUE3Qd5k6lpqY0fiOuX9+LyjFusl8ZDp9Ohpq2pePm2Tc7v
H1Lhf/GWc+DJ835LGjqOY/Ybv5fpPl2Fap39yCMchNMUh+Q68RfHP9rGUWPVfM/3BM1buo4UiX9a
WkPgotaDAeCpx1QIcZGP58SmIPGuyCEwgPFwLNf8YUBeUOvKDPJZRa85xiNuFYCVm8HHOvdoNgid
tnFlaTJHh5mM2HvZadBIjyluQeo19szIgosr+JKfXIfd+uJOxkopD71bGjoA9lV8phfuKzW0+0Gl
LpkCkPDEDD3NHBxdu8QfRUF9WN6IavLgVOEwc5G5xcbdPU5blj1QMfTgiY/Aspu94EkXVtv02r4b
vluNGmP6EKXqBbvT/gGCqPCoyobh1bUArPw1gKPFYv9DuZZOYska+bayCf+VlItAMw07dQYm2h2x
NnKKntxEVSPBQe/grOVRZ2/KMD5Qjmf6sSwoslYQsFJzjDTaw3sN4lc/W91phTkuFgoM8uKjiWWg
GqytbCd+uJU5mKw0aoStvpwY8I0cYjCoHdyfayRLEI0IGwK69ud9pAy+DK9IyDKRvgJABs6GzjEx
aWJzQu7REf5klRUB7QtEUe1WwNZUYrrRlzNTYRxJMtrCkLyDHDkYJYfcABEfztAa8CbkrxqmBXuU
KdTbqZVHjkcZsrOYz7VGrq30Od534uqJy5bEHt4SpLgEBpPoi37cfBS0Waptbz+0Ki4RwyQHrlYV
VGO3K6UfdlCDfNdm8XHcxTj/QaKB7tu0YgU0sl6gAPV+HxTSZwAapwtewQNgWoMXi20pXhLh85JI
5RP9aYIlZhDhtZ+XdKabXD9W3ehKU+TMADwAUt/l+3ERhiwViVuH9WPQD7oEpVY7g/TQfUDlfHEU
wr99Wl/lx2tl4aBUUMWwIw4JAgtMC/u7Eq/h9Uts9y97v8Srygs1JWK/fOv1keBAFTqbff+Ja1Bz
5m8/HYiHm19W2BSxuiE7sdjX/VYREMCRF1ZG03ApFdMFo/cbr8fRvgw7RqNs418ygqbK39h9nD9L
Q9GHNhWVY7s6Nw+dOX6jqO6yOC6GaJxISUZ8WknmbBmnGbsb67T9ksKmIv1haCd6nK2bqsy++MRJ
CBMUZwpQJXf3F3MrWhEnUsfJoYFkJtWvNoKZk4jDg7y+sSM8V84h4BMLnl09sH7Foa1uKwvlrSrb
BPIoQKEOb/bdjJ3eH+ID0uTvac75VSWtNUlMjyZAwv70IYK4ptrMz3Wm0+gpBxuSW/zfvGpdEvE/
EEbgUYScMhYi4pMVdTx2IdthmWEK7kvMHlaH/DYPQlofj8qHlNBcmTmVd6qp3UYhNQNVobbzSMFT
0VP5u3zbUGLeS28QmgkD893sk6TCwjXE8/ttNJG6ord9PKqjVGTdr9Ye927IHa1oKspjXRjN78oR
FrrebMMJYSUPC6HYqji+x57PXtz5Cle4UQ5+o0p9zGA/x7bLxdxEL21eZ9aZEKOvceFIuh+zDZoa
n7HWSD9fi+ggWnqwSCNjmyPYdsOn56mUDKs3I7JKu73TxAYB1pv+BOQ7Ha3n7xWJ+nWzYerDGZzp
PKfHn0H7fI9nLrPIImZw49WNFWpsI/nI/LX7NnSWo53gFqf8Q/UeYXGFJsagwTReHzxcxic38CPz
zPy2wkNYa+zHWuUwq/O+UYO/zUFcSA+2x4H3SE4M2KMuHs9dVm3pUgFlPF0HzA4mcbJchDHxNljh
E+gvowu0wyVAfE00MvBrW2ToPCo8DWscRDabUay2h7UGJwevsRyo64TvO6alaoCkegjOhD1TkX2U
1TVvKD7+l44W7V4XtXXNKRl0IK0xCBdvwKct1IOhlbli+qaoxuMFwedcdD6XnCNmkJHakfVRj3CU
uJqAXN89VmHFNGOqh1e3zOVQhbDZQcDp6piLCreO6JgY0yVokbkPueEcTOmhze67qFlmmx/btkvm
7B4Dsdd7HUMHMmNrN7fEzb72j169Wr4lSLantvW57N9xzvJITYLxEt8NKZeGreVonqvktdyHeN1p
6rxPO4XHRFmIHjxfefLGrYR+dy2oe1aPn5sL9PYGP0p5Ka9JQPtL/kDoSikDPiGEkqoFr+d1qsWi
quImyQE48NVCXD3Vsl9L9kbudom3QoY941RaBbxNDRV0b7veu3mKDN+GMZtwLaSYotO1GgjwTFXO
RJ61PJzx8B+qcUXbpEgq3KlNp2NrF7XCXN1YPk2/UZ9wXgFIMRsSJflaudng2u+3rPfVVaq63+/A
NjIJc9TjGkyE5pSTXbeJBU/EijiumL8RWVj/qeaK82evczLsucR8NkV0l5AtzuD1yHYvjCMaU1Xd
3VDNhwbRSohPMy7Jx1ljiRQWxNGpciv6mV8nAivEGVSwi48jHDodthWb9uaglbTduWwd2R2M3YnD
d5lwzriVPZMJ+ZyIl74598XC7yOPUL3vgOmTxqQN3xn0U7V3Ln1cBtoc8pFIzKhLW5xwY7aMvVKA
FjpxYDRlbY51IcRYookK115XF4kmVuubOuO6PxSRIqcUxKWFjm6VFpKjMVjo6SOXeThTzwYDPnZ9
aYz39XvDkKI4eTEqz0WZHr3owcHKxKJTw0+mymnxpiFl5LwnSqoBQrye1Y+NUeLpM9O1qO5oyGl/
5x50oAxc3RE35uwm5rgv2s0frJWxZYJUgIsDJLRnKO3mdVSl7f56ghnJRu/DUNkgi2zeJT8NmoSX
b4/yKkgutMhko/HlPC3gRqusHVKYj/N0HppjZxV8ecqO0nrq2c4GznGMaR9isxMJ/+UGQsESbSR7
b9l3IhKBDDgInpkSDDWGU6Tqb43e6b7ui9BwamRi1cXNbceq2S//VEFjk620W8Kn9ubHsZrqsipY
bhyCTjrqa5HRb/4MaOSurLK6BLrNK3BkRtytV9ARX0Xz6IC0xAHFpNzvxf7APzRm7dZyUte2kipk
ltwuLFiRkR1TtQ0XgR6Bndj70/435OHcTTJxR96eDOCaJvMaxm/v1wex6tffqhsnA5akqoM+F3S5
IEBtwUQY8FK3uUG4oy2cCFaRX8nojT83EDjFOCWvjiAFR8DqYSo/oUchcmbKetiR6iunal7UO2pr
5U+0lFb2fjaRB28WDfCblvHmRBD5iP2uXVn3CFncYj4y/2qavbJ/RQBqsh6MsTe5tFMPEf00CAqU
BroTZzv3n1r/1ueJHoyIMV0BbzLSnVbYN/Z/I7TEJnNtcVldKrcmcWUkF5pf+fEL4fpG1shpDZzR
Eh4uBrjf6USbBnw8j4i01iRHTcgcdcCcNjcdaLReSwGjDh9PmTolnYer9QcCXxlrsyYjLKjU75ZO
q/3cH6LAROFUO0HjcQYe/8hqIwDFnFpBUqPoIIX5r+TZRifXGtKALw8D3Y+24aNRA5kmdVsAyaUy
vZsgbVRhdA9IZ3YgBGhf/YLmXM/+Y0DAdGCMNIZaEuf38735q7JsQIM+e9jEoGld0nHuZSDhzJxy
zO4TtDOASCk22B/U0J04j9Hjv5CdrC9ssOsfoN1RhM+kxVpEUD6lXWOplGGHesi8G4cFUI30Mkzj
GZZc2KL1etiZfta6+AwkmPLmPofqln869TQbn9Uvv21Og/i1Mrpu/KQvQp14UfD85GW1MajjrNr9
5tsxsmMeoRim/DK6if4+Od/b6XEGExmeIu9DZVaH08nTXuuY0hL4v8zlagfy6Dxy8QrHiXKk6pf3
GgR594N1zxp8FQif5vO1dq7qzQy9LAT8L9kQLERoxr7r6WdecYjmCKMpt2UMpq+iLVdNa4tqDQHR
Y6DHBbFZ+K+JasdyTpwztKPLQwTl0/X4hqrgFWNdDseNZDtvQiZlkCdm7vmlz9y4V52AqfRQVtcK
lGtIoipYj/CNguEjmDkB97v1ohIOvFWgN3Y0+TzlaSCmlTVbWCqup0BO9sjumLclzfAKhpDQE0zc
ZYxbCKAmBdnTu70d3a7XN2LO1ZBlnZYpxjcRgFIFtWci/izDVZrWVnIwqwC0qGxDHpVzwizzaHcX
+jd+1Uf5GdUdKk2IlMlt5QuaE3x/v7PWheIbdp+fSEy24SNj7A05+SZXeF52LfTpDwaa251FM5Ep
T7L9mWx4ez+pSthXLSINiIahY3E2YXsAGk4vRlWHK4G7rOoykCVoEwrvua1+YI2WSfivJGPHgeRw
4ynQ+oBPes3MNalVKB+kTXXGSZGfe/YIfNx00K/1QFfhcKJDMNIdcfcJ0Kjj+3bg14jdDLBConCV
ggt0msBLqCE8SFJCvzSC0qASIy1fRbHueIjoOFdXFjtwsJSAK7OSeKDlZqQMEsewanKYWoIgOOcJ
4njvJejwAFnJhSXo0Y4dSOD20Jln5WyHOthxlxv97V5/a+omf87OGFkPKDe5uvyQX9asuwcyGcox
Rlt6xD4FMHYsi4o4GgJk+tKCXI2LUQnHBSGOj29hZ34aEtRGrDi0UgJd3OgDstOkr9bNi9CSBXWN
khoPRcGDE9dgafo8Lr+S6imzgIyluee4BImBqjHM4jp75F2QkCHyZAln+eEzHzgPEJNH8hdeb2fw
u5i95dWLBk3NzgtQG4t8C80PhJ7/+E/baxdPNOTdPcX5PVZkBeMEoA6sAWJuwqTzRdbfw4Mh5KOT
c/EKs8pmBchTleFwAT3SOANVXc5Ti7toD+iMEPcjZjZH2qDFKJaM0/EBA/RbVxdqAklmGj/R5ajK
Nq4ZU9RXqsH5PUEFl4QKUsLuJgNKmboZzdK32fTeNRnW9yrsBndEpjx4TiEpJ+GOOZya6mVXkg2M
cY94C9pQI7chaWqsBPyRyhZM05d8JUpiu2wapNEi8qcHURTjvRXIIEqSNTEPqbvfyOVsxFPiP2c3
WRWDdbwwuzQX+fZVB+Y9u51KA6PR3aV5ovUiQi3BUyipVy/9QIKuhGfwJ42nvXBCc9rrGI+7yZZE
ZzCfp9wm2iVh1AYWSwURVqaKXGi6lx/UTS1VsTOcBau8/64mPqZbyEEEqX1dCR0PBR8tnJLJ3Kxm
uQQ7WZE4B+DXQ9DjPA+Fb66B1num6Ox/WVrHs4BL5BkgqsRLlNquf3r9F5LV/GfwQbHXrVXmpGfH
LDREJMe6iQ7ZtBteKqsrmvcx5LayhTTSGuKBbMOopyT+4EQNqbhMVmzIDPRRbprt7gl+s22EcpQZ
fzHNmrUuD7HjVs+IETdcmzE8Uy2SrBM3jYMma2uzpW9EPVyoB/w3K6I904Ua0IPe79e19w89aT96
ncraaN58FvcbxJ75yPpqTtgHvKiG8xJwZHZUYvhk9bbOtFd+G1ZdfcIsH+RrxWJD4rk/rQV+tlgP
q4bcDofWCTbzFnGZEyCL80gpPVncibt4LVTKRDjkjSEK6PCjLWzDgPx+BgUG3gvFq6Z3eqlWiDJp
1pA+RSM1Z7NMnTq98iIygXB4oWq8AvI422Sa8mJPiDl+5GctdOnmFpoIVaJrb0imsZLYAdHgGO7H
BlWBImyktvvRSIETZOz1SS9p/Xiz35LjDWP3A7qP/PoJ/KDVcsk7Ii46fmlPmCyEio8eBHAf2a7Y
N8/jlW45PuyT7lKoXkFfC1r4ha3gST5OM8sZMyPR9/Zz9gDENHFLYGt989Gul++QqIIt3hJEf2uG
L7TrAWUaCYA4Y1D1EuBaU+FZD1zNaUK3JomN2H/nUrutMIF/FzC4x+k+S4upcLjYmlxZzAqI2SK6
9anqjibe4fG2jt9lWIP5XhkvqYCb+6r6VUcz8lujYXsaJP7hTRYbJc/3t4g2939V3wv/bn+ikyCk
0QiQEGbP6Swce2R/CtF/Ak710pq9rEjdVwqMRRU72lnkPnCPVX3luQ/V/832OYBbHnP3uPYkNGH0
UvQuBp3Tfhn493Ft2OR2ruKQx35+fsSsdVGMu7RG0Zrzui0pVTocLBuL13jL7upzUJSsJlUBDR4J
bpXcVauFN05A/krgw70olSzCxR5QgVdZLVCRaHkW4ceUqxvWiM1k5TZ+WNqNC5oagb0ySZYpPKzH
HhbVXzgLUtBZDFQQNUbQZcf5R9LfVsym3KehrFvOQaZswHiZhBpaCzkAqckc37PSaWtR0ojWmwTm
iLV3QrJ3xt/XjANRHHrRS9ERVWMVbfJC75avp7g0+Lc4jWyno/y2FOUS0vm5uRD76BeZs6wPN5du
kAPO6eKQ2fjQjK6M/A3DPHdFeRMhACS6E2+oIyJeYo+6rAm0T984B/csxVGncAcKsGnfsB93nh9F
T5mbs88yPSLhKoxUL7ccO//r+/lJWGP6GAP4blH5yXfRXx4pLftxwWRNW4D+kDYfTu+njPVAxoku
ZwZkYU/zow5ALNtkscqpzdOX56A7NbcWpLGJXpj6fnIq/66tM/IudrBdzsUabt9gJaOJhK8H8GKN
FDOQ1V9HZUJ7lMV7u1ym90kK5jBRgT7dlA73Wh4NEhvCCyf89m0oHoJ93bz9WGTv74cByPH5QPE0
eP7ueImodJ23vkD/tiQaOddv4JYtgQPHAyEt+yNkjjfCNUGUuB/oPrff0Lxl66ZiWP0u6wxJ9Jzk
avhYCvzPQ3z1kMBbJP6jJ8x3VFC7VTaO2xZ01uk017IBkFkyHjMWZMnick1vyIdMn4pjje3fyoJp
tf5r1Swsy7gP6nY1UaqnQm2Q5s6mGQZs58QQx8/GQuLkYnJr9M/GSPzMuy9yPm5C6ozAXDA7czB1
1hh1exKQA9icydIsLS8RTKtSKtl12YAgDjdHReEmfiVsfRB9/CXZj6/5USRZ29Fa2eXkTIqmzNG8
VJrPdRKINnZFp1cMJs8K1q2BRTwjFi8rC1N4Y1IKw8SuJdikE6Yv5MUADr3k/vRYINea0GIYDVKq
2xoSFYAxPyJe5dGpudaFDtTC7sjuYcqKLVVnaRzg1kJs9DVln6Pc9axGKNrc8xi8UM2JomHz5rUC
kuz+0b7TN2JPMAQu25qjjiNQukJMsSxCUYMQGyvZ7Rln5L1g1RJG7GohCmsTUHaZKDAXVbMF7Eu8
cJoXbf54rZtyFoYOqefcVaJbpU5zHRTEkLfhqg9kK8a0eNBp0iOd1H1E/qC5cerfs9FdyZn1E0ou
OVKpD5XR73TSgtvKsbrHPnuLvfAZ2ZX2nDVqEYmYBt9yQ/AcQuHlCVVPP7lxcvnL6FJ0Y7d0wcYm
uQkseDHBR5VXjRArsybFemHWKYhbPZWdk08FqKUUg0VtPbCTyeHhf+aeYF3DYPN5fPJHspbT9NKR
pq5CnoJGU7Ie40RK1BkMfjon0aQW31ZGGbbVisUC3jxrpqi6bFurGNdXCOpBQYjjzljANfeOqToT
4aEVKj95sZabOfrob4torTvAyWhXG71VojhjP/FMAfov99cJIqWfLzyxpx+R8f2+R6pWAbGPSbPQ
GAlbgK+99fcY9SPPCra9/G6jIMNhlV9iYhY/L1ZUCiiJzGS8PEcV//uDuawnnUdFsUzBCG5MB6q9
F/7FRgsTTLUQpzGjRtjYugHY9e0pMQJVWoOyiy+RrHGb1cznBVPl64fgUy+qvd8tYQBGTz9wJFBo
kpVWqUQmGExXsuzjeQ9Re39VomgbTf4R/s2Cif1ndFzmgZC8qeJDN9/DB11eeVXF8Nf1vcbE2uQu
HPPuXnwPEhmFjLFP9QRHhGp59hZWh/+dZpMkW9HOxHc480seTk1lYKJgUHgU9Yr6mviFHOKtylwE
P+4Ccpf2B9uE7EnZ3yn//kb5WOWfmxEHawLhYuBVyorksWcrYhZuFXxK/j6mzn7nN4tY9vZ1bw2v
o7DxHzDciWKJI5bJkT495IOfhZAQOjYiZk5uvPBEmT5yDh26PAk6IcVXpgmGdVyUJALtq64YdyX5
PFlNQLoEWliU0A8wufEZH30Y30vo5JXWb0yInqh/sLWwGCmRURf5xKLmZkvoDQgGrfwIgz7+EV3k
SS1NiY7NpamgdXnPrNhRzfpPxmKdukIdAPzXOWg4hmtxb0JJYvE7WcxJyCYrEaSQ8kjjDUZhkrwm
TKxQZAG5Hzqk7LGTCp2h6vPDW7Hi1/OcfYQfmkPZPqVF6pbOSFcA+Wlv1/ajhjMVmDjF9bbqadBB
GadQLGvbAJXlOKdIUvpZtPrl+DL7W9vo7sINqE1FUaBokWsfS7whbzxFb9P5N0WrocVgwG9tntXm
cqXOEJlZBKWJ0bDpjYb3ukP8xR+eYC7X3zWd++KHN+OtT0OUAJkVzgrLGxaBmhsdEVM6h525XXT0
zcKcASwutv+Wv+gTgYEfBSHVi1AoAYRqhE9ibtklr2gjNUt6i8dByh9jw5AqVlFU5dgM9cT3mD0/
bfe1HFX7HAcy1uqVPC8qhGaZatApXiGYRsaVjDo0hWjdi/KN9fCfMMyZcklumKXFc7S3ifmPWdNA
EO7TfGpmGo7rXmM/h+8ZDAV3c4ns/cPvSqkuggYids/WF3OA4y6Rzcqd/OE9wt2iYiMYi6IN5SlB
fStcd7Rcq0e3Ud/bPy3tEUjxe93Vb/CMtM9TBcewPMUAy9w+kWUdxYPy/9SGPb2emwLVS5Nyk695
2tB40ahDcvg/QCMhdVERf9rrtcXtrXqlepbBJaHHfdbGruwR1S9uH5Q2XIa+itpTt6nDfUoj7TGK
qtJze8+v9qOnME2/nfQk0c1TT1HjkNVIOXwnUGUTirzT51oNJeodXLEZ7j4Ue/abVECc54ymmFZ/
X0yXGNtSzcO+7qPWD0Le1SdNd7Zr/lvksQuRhvSnKcXlw5gJ8Vwc6E9Rk9cSvl4CItWSKmuEWjBX
UYg4V2DFnMqRtUbyaL7+mRzmu0LAMew+FCKx6aG8UbF3XaXeUAALlVWGxquoI7QbY0pRxr+J+zhT
cuwgSQ82i4/D4uIadwNxr5IrppFmKYBusnrg4+pWDitUFVol3EhQGaolmQ8VzR1NADPGvMaQffYn
dFPsA4mRTTSTVRvXPdlYt9omd5Rc7xXgJSPe41ZspYDhvBU8slhzYVXpVlm9+CqwOt77fjFaUyVs
P0m8MMHyCNvFaeOTGRotpteopC3trBxczas16t8g0ilCEqAHE27/u+BroKuV6dlCYHFZWIbs4x4L
byhc0hwxfkIM7+bUhM0b0Vp+QQwuC2KWdAp8MT3ad7PDXtW5RChd5A8B+Zd0tAXII+1R0hLPvlqA
sc2evhL2Ex3zN/56YLXDSWK/4x0B6dF27x2G/KD1G6g6oe6LQ9DIssNjpL4KcCxOn0WvfeAe780W
8HI4sHrZJK2nPLJhtZWVeIl5APVuaBddiySOaaVI0JDLhgWTF1GXgF16JExR8EEyfUW1fRHeuq1R
N3X0O+5+RTw1iJwibdvfY0YhOZejvTaGCRSJFoSTRYMskwgDeBw6ZJ19MeBCus3zJ5gPPpQYdIhr
ORaMWxkfitbzPTh8Qy8+lQ5vMwv1WIrNBjHaEcKef5zTPBtxqM4nNLWllLQl08S0y9jeapIugY/A
r/lbMQuv15J/MQlN1sGaEeZsfCFIAZlJ9RSw/nyUK9ntb9k4/KWmdFZo4bpTyTF1MRmePvNvsfpk
1Fs1RSc97I+sG5zN/95nTQ36nXYcPO+R7/OkWSrZwVYFEUxqtb+tp5npjYBPZDnaM58QIoBFRhoM
18/suxpiTHqYWkueYYV+SEQQkPY+9apKAKbTjfKNJlu6hjZiipVW3ruhbFsMpR6Boh/FLX/r2toA
zEa7lNQAWHLKSs/ozkTZYbRvm2P2r+XNyXLBc5IO292IH4CFZEs2N0nDIVAJ0LnAogJlKOyoZFPW
VDKJCi68UZgLZm5ZhQGTLbZ/SI2nBNhInxJ/Dezk/39plKYRRS6x6qo6iRyUVACtunLtwk8w9A87
XDMq1NKS9XV6g4WlCdT+v64NWcUrfaYng9Rr2nLsdd6rlAzz1lHFCL7LB9u6xDmgFu9SyuUFmuJ5
KxMiFbpIU9DH2qU+FS2eknuAtnD4IVNxf4wFypjuv4CVa7KWU8HNRa95ETATTdPPcL2OpTp2lzvb
ZV3BNuRgu4Npf8VUxLvtRSLTqMTG22PmgNsx9wu3HEwhBOPjXAFZdfQO49ci74ac9UJXbjiJZwws
MTbK6iNmGK7oc9nmuvaXGfNEG6ykSpS03Y9i6G+Kg8PkOIHah8elxNnb4rKF/F8XvGxABfC3878i
3G4U35E8zkiNiHjahZhUIccO/WKm162Yl5WUQKLWq6FEaongtiIe5RV9o6BtYUVTXg6ioNZg5bes
+fYUpOMiK7HVrUDOzJOQY30gZZAAmB9U+7jKBTU/WOg13V7X8+468RgifeAL5RUjSUqTtrXKgtTY
UM3sV70iIqQJRJNSZHfl4IQLtgFJQl/0A0fQsOl3kEKAHeWPBALscEu4KGqvzo6WbVdHf4ToH9Fo
FQtcXZpCaopsm/q80bIu9qkvq0lug4mvfVp/W6W4zTVy0XbBrN2J/ZOmJ7Qqlz/8Rr5xTH1Gw0VH
Dme7gDZNXJU0E4im7+HICOPdmvh6X+aWRbTaVWqLYV7dUR1gF/lzuuseE3Ty22M595iZqBd5ZSV7
NDPyXjbdUg6IBUMVfPhpLXXM5CGP5oWcZNSZDiGvDtkTIpgApMX+PsbWv3jAEb3ZYZ58LgKEb1uN
sn4vO9Gz/Pe39ZSH+0HZuZjWLrCHNRxFE2LHx6ZwD3gKfCkIhlSPS5mhULzkRjzzQ22GSPoTCdu8
WhyfXeaccJGTYXjLFI3rJOKkGvPZaqb9qzq7Aj/iksWa0MKgMXYuZ9VtY/crh08DyjtvkEE8Xy1s
Jc8KWWc2wIxV7c0mt7ZoZw5T9mVXHzsWFcmJF2DM1wCHHGjTUcbpYNAoZT+3LZ3bbYVEUoCcT65H
xLPiM5WKEcQeg1VjNsY5bB8glbaea/n/CD1OelGt8jr/LogMWHFIsW/8m/yxM6/tXK5CZIkItbH3
WEI/zHtcdkCRcVhYpbJWYyQLJRVTJ7QVL8Sma00NCEQes30e6y0yhypfXQLR57L62HZ0Jl8rta3i
rLyvO86+ShE/wE5PQYVcizkpgDlPSYV3VzO0bxD4VRLM+JhsYjkprIue0GJlT0H1OzqRYIFpxpPo
ROQy0OGEmJLdLDZihpSwuMayYOHJrGMiUBjZmQ9Unwrh6+5Kf0RILUrwGhXYEsfRL82Uzdgo3QQr
KFiYi816LsGzAJww3cjjaeBwZly5PY+T6b7aRgagO2RMFtC/8euqzgJtMHyA2Q4F+kgBQUZEMO/U
kFDAtOL0FofuOHC4Zovf4WQO8aIplW/2CI+D/tAQKRnqIk10OBbwA2BLqaJrzQy3QDui/twoxaP7
olY/ypusj+m0hbDtuwVF8zm2rfYLW6dPm2MmytikErt0n8dQH5qInKZDH1uJFXlGXjFv7+znuKLn
9ZpROXDGVxX4SgOmJvc5bbYp0z2k56akaoscHs0oMvsSZPxXycGN4JlM7V2Ugm+csIUGQy/n4sSl
vKKOyC5l1Emkw6qpRX5QxBge5bvn6uoxWGgdVgm3I3L4RCDbrGP70t0d3z1Q0suC6XIEA9gpISbA
3Kho9XF3Up6AeqcpTF+S4l59isKpTRMn2nQQF5s6+9aWU+ipex4es/hSQZ+5W35uYLVwsh0a+c+b
bWlF4ck3WGCXj+6czi7YhJg4QwSfGJTk2eSutMVW4O8ggclNeztctKNNOvZ0jmNGqDKzG+JSKvhF
cW1Rtf60R3nlOVnZK/jiVw2VURJ/kuqBxbUNTLSfRY/uvdnkGM+lSluiiChOmYyISccQ8hdzvCkI
gpP24dZkfOC9rP6ixegeqiABQ1SpegGuGBoYglN1J43i736HG3ol0po0vf1oT+GCVL0HwEvPkb8L
Zy+5pGsWL4Hf2VSaRdrCX9DP0PJLhlOkt3emgiQ2joqSjckm4OETFxIkXjeud88TUcrd1gbGAOjc
YyBkLCtnBfgxUoyJSEs950F1u4Ex7QQT1ZRmidI7Vz6kdfwo5koJX/pFpJdk1sKSk6SmxrHPzOxD
FoB0XAtM5SkNmooThfzSulXQNUeAdivpJnr9HEpF13P4FJ8n78YoE7n+eCrW2coeOszJTjl+U798
G7PSm6XeQWi//Z5jdia97gQpVrYlh0I4VH2Y4MY0lQ32EJbVp4LoRoDBqmnXq9wyMJURpEuCI4Y9
8Z3es+ppYIY/9BwTi8CpNTi7xnsl9YenrK6DGWsHqR+ASUaA4vY0mR4/xcq8BCXQjpsgUgm10A63
hfd/o4kT1BxUfEwhd4tJykdxuVQIrvc3vG16yaCl7Zwp5wmR/jHqEmjnqA27ifU6yKkQF7Qo/wtj
vR943AOWFCSOiat1c4wrhiA2gtnWCDAI3Dr05QMdseFSx7v7RXG6XVRd4ind7p9uIofP1oaSxxYp
IjQZDxWcZtUqTlADHjkr7VbxxhMx/rOoV3Pkh8MI+szZQxjxbrdeiQezM65cbdyKkIxH0Zbl1Q4D
4pSALqnOW9aSTeLf+oLOaYWTiP3WGvU78Cze8AiIiy0FtMd1mzFNtfyLHiNW2/V9zqbQiuw6isPq
YjEWj80Hk+7gVjFDR1ery8tZcyVu3H8RY1l4jSys0vSjKGGEx+cbbdBJ5Aq5Pt4oVmKX+rWdAtXM
K9zauhrmeJG3bZrLsoJQGtbidjCdI8SLLsd6l2KHFc3uZ3FI/IdkA8GeeNbfwPi060889oXUA4JH
VpNceaonVuL+NbXk6iHCwxdWMnjh+mX/hn++g8TmoPWUMineoaPLMEamqyi8XhekwQ0/yAtYfQT2
fbBE9oITZORp+5+7Yih4u5lRdklNtVzSPNgIBfsVzAtpoVwnvaEx28RAwHFvg+EEzbyClUQfFL38
nh34KqSMpHSfF6K/qidB1LfXe7J68PfC4JKRcOL6QIfvpe82f4H7s11CW7Ib+BBl92AD2grjtXke
kzN9+obnFy+jbNLRYOa2QsVCTy2iZmG8+1G2F9i/xDq7NReHNfIg0P8vK574KlYZPan36Tv+RFIn
cZs2a0UtzUsVbsm12WsuQVzLS9lS43KDXfc/c03NuV1XgLSC3shOCk1A6SxrURI98JnwfwbViACh
MHa5l8JXqB0VnLNc01PwcYvMoqB+hkzQ3qb2Z4pynX8On4BhRJBDrcUUnsE6vDANBj/iZLGfU1y0
FhcJ0wIK3UZPbTPEK3/WER6slzzVilXSgXSW5qfnzaaDbqHxk+A27UaxY6Yv7b5oBokJAoHuq211
y4WzkqLpOvfZ8C0tJth4qNuU26c2tipbxBCDEn1hcx7dPu4T5G5h8ucLQx+jK/Dg7hSFtBxRsnx5
0AbGJqNT0FSYgRK0xo3x8N1A/hexypPC7Dx3RSCudeHG8HN4kmrzwRnI+0A43L2nrMaimFcoaON/
gTJeE6xLhwurGDQYFallwt9aUXmYqriimCRVp5uFWwX/qBezjmE0jKPFOIG/sTldJ1glFFdw23zk
a9ML/jgYRyXw1E4/vSOioIRB5pQVA+c8uGBKrjxMCNl4sEWgTV993alnj0HqZJ+FlT8pVL6T8BDH
ZpunDtxDn5Ejfkh2oAW9s2eTEwt/X0G5K+GnS5AbaOEkT5IOVMilhEmyHeeM+OVdBpdaewWqY8c0
4U9xQxzRtxrIgrOrrRuUrlbxoecdZczMzttpYICseIi3F0IfPF1/kOTtsbG03cmqMBbL1ik5I3va
eYHeH/h4VVNRFqKTDho3JoLvWwqm5qTKM4N1FZCvmLG58h6RpEuZ7NlVA0slYEZgkJ4GeB6ogqAm
yqnzhCFPu509hNj8v8InQOzGWeJTJYKCohG06jTRuYriCXOSA6+hcJMHQi+LA7AW7Nn2osFj0vfD
e87JzoeP0RtcX1Mq30ew2Bf/2cHLmqGUxVJ6hLLMg2S7Te+j5xiUR4SGQ2Yx8ScHPEES/GS+X0M7
dI3mG6tCD6WtwtTq4GsZZPhFVTyQTFiQUTUScjjyqcwN66JTg+cfI0ejna2q98CIwo9EDv+WP3QT
JWV5EBE6GWPPTcyNCxcovbROZflwRz7bVGoHSxeyAYQYk5mU7/ER7GLyi4cfJEJXGRG5xmZ2ggUJ
9xqEzC0/Y0MAZrKYojXrwHcokgtBrNCZDP1LzasFOb10H8nHywobEHxHRt1Y+Use1l0AMPhwjKS+
691QGp3DiyY/n5/H3sNPGNcJ5ZrUP2NJaUZ5f0X/bU6+h8Kp672hYXEW+b2r6VeTTywP18YiB/Kl
koPkWL+oGrICnl1KZCHjx9C5ab4NXTJ/Gs/XBnRYRD3Dy1LBrAEg2ySt/aqZdbSKgIJTpK8ZusNk
YYZI3j5dIArxBPZ63WPeo//zWut3KDxCToGmN8Zbc7Ukv51VyVGkLlw5oPgcMfRW0UwGDetZn5tq
BlFrWrIIBnw/ji0mMWjd2Q32CAqvGApEJjbFTvxhjejBWPkPG1sy+1fBDvEnANZ/ghE43TgydBCx
VCzAuxw3Bd+bC3LnIzx0fKKZxhZ6UgsyrcFoZr3Mngyi1zYmTTBY2wZyKHgA4VL5VztR1f53A+SF
9I+oVQgklgy35fywLOU4X2XnzzTeKyB71aLpEw3EtxEpb/amvxXY+AUZLwGmqBcKEKtwe57VfISM
KIuVTcdBTbK+mMCZZu+cne2Qz0jc79WCK9vgEqu3mrbW6RQ7JxhOHb2d0KNu550OYNxbPJY9DRa1
KMoNkyO9Hv4j8A9Pnzkg3Y9PPZYDuyY28xBEdn488cImtBIoV20lK2xpcunOwfSyNVJUTrMkFPbv
lRfLK/tDuCACxyJImiXD5UjcbdNgXOxOVIOn+F+AgLoqyoVfDIDkRmt/3XJQckEvGiw3ru3npirW
qTXuSx7Xu3sdF1vZpcS355/ib9PzTqQ8gx/iaxMeRGUP4cckYmQcmbhaZ8Nb4jmpEx20Y2KfVK0s
kqbIUmQx3bp2doWDuUUv/NBW+zOlqLDEkRZ+fkSzY2RMPXWlfVBaIi7oVwtA3Sk5tnbYfxps60L9
G0HOAOW4nbm4jJYAQfdSLOq7KNO3glh6TFFE1u3HIVYXY37wN/ZjKCM0oi1N0twJ5TWiV+C5RZVX
h4M/xUaA7BWrael0WOFUKxzjFR3FsM3NtVzPmSrVRtSOiBzmeqC6ZiVH3fPfm3P87aok+HTXXXnk
PZMlJHsS2A1RVWFohc8E/6mwRZFHYOGXnk/h7flEi4biFdSIUBX1ipna5DE9Ud8DhEL6w3XkSEDv
8KpVHnqZ5ZaDg5jF8EfpH/rA1Z7DTJzjx/bnZ3y38a0tCWuosjPej2MaMsY1EPg0Znr38DJ63+WS
rotndlU8QSZDXRSNCM5hoPW2jrDUw/x4mehTlaD7NBaD4OKu9OUWKcVIe5ZxiAs+/qfFHyzCvtj/
5WKecaXLXT5TMPN/NMoMU0uwZ44hyNufWEUFLaLtVEXz7bvN6dSYsnIbBLU1iLGejkBYhpKZOvck
lr/aSt9uAS0I4NnQmKZwCoLWEylBxbKaGFSYAiweAlwC5O4F2WBw0AcNuzlc/1EPhkLYygF7NfiM
/RdoNepCM1Af57wKvPr+okkSDaGBIBzqhV0hWzFP2cJep4pGEiIIcXK9b5iGMuEti7GhHjGvacXE
1RpOnhvjJ+2Lq1g2SYoEcAaUZAa9KMXGv2tcW0K4GgPD110bL31FoGz/k1beZlDLEhYCx1ZAgUzD
l4nRih9ykGxwlYgXx0EdLzPN79IjokVovYNxg6Ye9azlWqkpZQvi+/cWN+BsQ2jqgvofhOrEVGE3
b4tSgU/1Q54lCtVZQaX2CjxN5BF0GAehltA/kTJMF6Lf8rFwlmXxqEdHJF7kP6DmHaR5yhMaCFrs
EA2e8K215Gfzu453VgpK7zVJYBVRakc6NBSIWL1/r4cElNYcHewwM32k0tUkZZcuYyAQLQnK/liG
JTK6v80XCil3s0+XCfD2oSFJL0iKi3s2s4CM45Pptls069chYy5Pox/YcOPtbLQC6nxFIV4S4BOn
qqmeAVY+o1+SYlMaIDpOte9F1FCJWNSSqZMx7+Kp40KOLnYkDzWFehCeiZ7pUjCOGzR5WcVfev8E
JeW+j0HqvGu6nfMohGzYr5HD5xe+9DpOJS1ht4vNoqiEAuOyzpwJz9eKraKbTWWT0tNzMBFRoDv0
S3DoYv9rbR3Bg9vtKh31gyp77mFegNfS3GOoM2cr0kjxSTaHWIctlM7My1K4Ejor99Vy7M3oBucZ
K27NbVRSzGV5aZL2XmBHF1CECkkOU3LZBX4Efkj1+ChPlnh4tkUyXN5yW+KIPcqPruTEc2v0jsxo
AOECUiLgt4DvpEEdhClsbc0PD/EANvxPD2Ypy/Q/8Rq69+gnzpc7mibZ/PHRAnMHT3/lF0ARU2P2
lC/6WnxJNJJzUgmt14vns7j1JO4AHrOYK0dJR40MAJrTNhpgk+cYDchUJGZOgTP1wEceQAijDeaE
n5J3TMpZJDtHXYArvHFuuiFJF1dnN8J5cYfKQj0nKJ2Ts48dwMb+Xjdl7qpXlIdBUxtj2S2K8hMr
87x84d+m/RAdPBjFMjF9H0B/ElkUY1VNYlxjNFPS/PklGXt86bosKbwcNb2d4oj5JsrT1WiKvLfE
9ZXXP5mfwESjn3nwSxis4/5y3InHZqL+MQUkeKVxA/kyQ6LUI4lZS6i65z82/QboWhXowDk0fuCr
S9fozKMiJSmNICGY4RDuo57DyGXt1DOweEilLu7lk38XCFzvMzPgaFXZPfZFOiSJjEDusLZqHb+4
/IKn9eqVDK7bpvw4mU5Zj5rYfy/yRYNr5N6ggjokx9B/bxiixwzXOnyjsijyQSa9C6exoYPtmfj6
vOn1PDdWv4HMq0CstGNk3Q7VVnVkISyDmh6GFCGaFi7sBUtkApasgXnaiFvDysL553RHO6T2v6Cd
aMP+uuoS39S32uAa6ByiGRJSi51199ZmP7Qz7yQGxoJzjiHUbP9VTeRuKiBQVIo4oZBc1dmsnneo
lIZhRv4wtJtsAJxQhRJ5j2KnpxtZMgJPQxHjah/0sCjZsj0yTZ8z3DUdia+udn0FEBc2WjM6rFxG
b1HEl67p+HL4I/6FJdEOrinV3StUy4XxJS6u266mR/7l2irTugUeZAMeAFVtY8nz5GCOEFeXTMGg
KpLwxP5Wze/oL07V+712Ul5Fahr/MQxNqnDTP58NILM1q36vt+EhDaewvOHVaZr/bVsI2P2kInce
2dh10NmP6zupkYA0F6uHFftiSX5cgOnP+UCIebL7wTOsjnR7qpOy3xJyoTsk2Fhsg5lGH9zydFH+
m/H/KcdG1HgsY19NkGT6AuVtwdSqNpBMNQgf/VBu4FkChPcyP0nuO2wSx5uOaOyOw1DL+QbaFX81
H3r7/5vvVmhVdnWPDxaqTXxjnC2StVAfnXlyTf+2zQmeVtKz2gVgiIxqIbj6s3ZH6pgxdAYZ6yj8
KObQaGbQpsVFtJf/N3DDAlQbPd8nBm7CM0l4f6iiIowVT7OC/ePcUhNH8XJFZWZzmGeWINHYjnRg
PsqGpOrKdS/p2aTTBjYvAkALlQMY54bNgz2gNTHzf4ggNbQkpb+/PFsN9gBzhZon4XSjjhS3duKW
qtieI8V2bwrZbq/sN7QsGlpEEYN4zZiWOITvyQB5DuXaIZV9m+JxcCy46NEM7Vg9nlbXYz88tC9K
dIO24ukC/SSloFwciiV8eXZNp5q9zmgYltwYom88VwN+zT9MIes4fXrl3/QhOMvV63oqBuYmgGvD
Iwa/WnAfrAgajj8qnyR3SHb+8DYMKnlwkDo2ocFQX9RG/78pUge4ejjCHU5Pl3o6FY/6nvg1xUqV
B36k8+g+AMRhz+6gLCy4Q9sSS3VopfGhBV5mYgBo5LBUReO/+FuIQF8EgPQ5Ll9i6Fp1sytfDdr3
FB7InYP/azCYIfvgYiIKXr/CoDGsn1NFQeqTi+CLVS2rqnMCSZ8AyrGZeiDQQOKZ/SItwszbjyhB
USoe+u3aJhBUl8+JJhX9qllRniEeggRVLp1uxzeWL331UOlAw+Fhd/O/euqYAVOfT/RLwb+P9VtL
pjNDLlZNd2zcSl4l2o7fDr/uBlPzDHqk0iOEVXSXDsAVmwIwAkCGFeu27KQnOlWFk9r3fwm1VsIz
wj7NN7M3lR5caIav74kIzfENMyjMTi+/nVZh1HdflhV42Ik0NJF5yp7qUBeLy+bgCEF5999K46XQ
jTLWOX82VntzKyiRd0s8foc6+7uh+Fp7J1Ycf8BFbE604ZRALZ5jKMCZaXqta/Z1V0hGsUCs8zwD
9Rlt2RrsemISzNnL0z23dUYQwiUVWRKWxhCgCON6k70FPcMOYVJaOuRIHuruR67ma0NDxk38WCFA
g7qoGjXmdRuvftABRDDbR3fQOGw3zqv5Pz6K2f0VYZ+/qBl66X+AADVnIL4pPIsjb4sQdPzBPjkh
CLZ0oxD4Qxs+sUSN0EsHTWtY2/l/ztSPuC50jMWzzWy5zSMWKzLqTJjGcoaVazW8Lm7DqlThSLz/
5N5SRSivClSLYKKtreqgoNoolmO78g/SaFV4nYlh6yjDKiyXR7rWGSGLSjwB2IxvC+iTq299j7+p
IENWcITQYZcbjX6W8cyCP7YlB9kjNXEe0g71vVGyjQNOXkDkOVXrte1rLv41F3EbniVVi228KA4C
2RSaC8Eovn0lm9ZvjnUMP7lqSOIyx2ryv3r0obX2Hmsyqo+hRn2J162fd/jwPjT0Q9ionP5JRj6b
snSqqLobaOUhGafdhYAK4lisdYq0x2T77wz0RuASmOZ+QWegfnKIu7XasickvLqBU0ZoW7mTcZey
wGvPeRRBezXtlCJKhBkBU/H48UrPb5xMfdjvOx4uZl0vGCSc2YUJ2l89FMuB6xrw/fqzTYmi2krE
mM7EzRfQ1UAwx2wFY4cymq3imoR6gU52rzQ6tjaFbVazHmwPhMCx+OS6qQH3MP4drxwsC6bUM68X
eo2H7vZBASmEGiHmSszAClX4QJ9BP+dQxbzdl0tfSCaXoXavN9KNf6Gcn5zveZ+EPMilwPlYrMmB
Z771J0z4hYUEikkJhiYmfSxmpEDFunpJqDo0uFR/np2mooWvKn42b8maAa6Yb6y9RgleiJagvUIj
SAyyPGrbhmjex9NZWg4LpBvgqtVjQpxKIocp/EKqpIydh7sGPOCuVApdC7MfDVMk/OPETCCFFy33
tQY1NtLbv0fhcMyKxddiQn+clIff6/tzNOydvuWpvy4uT/m3pTDMMhFApehqIQIs8hF0lprUoWUT
W+zo0tL+gj3FKyjal1q9eeD/Iypkvdpta1jMie8NktAD1OGDiVmQt2cMq/Ar1divQLRaVWzSbJ0U
i7AsaaJGZeamYqvE8fsQAqFUTb7Tk1yFUGZ8tYDo/bNsYfwRoQNtXLK+wwwJSja32ZQDQQkpf/ds
84R65QmCtJKwiHPsWPH96DMHTG5uqPsRUHws1qSiuau+RaO9aeO8TP6CVhA5jWv/LD9SZx8dngxk
7xutjQtAYsvzafsy7q0CLM+ZFZwdhQPtfuffL+lHmx1mTLr1G7rPjRnn8iEzlZjheeQotVcePgBT
0SWv9PJ+TDruZHvYqzkCDkBzpwt3mbKPTldV6n9OYpoK7tyBHB3bTBJAbH/Sfs80NQSI+Bp8dW8V
IZn2H3/EKsMZjs+alWq8s+5TCHUW3VqrCqde6+bG31zXka/9n3JfYzg5+t5uCreDYNyzA511iXzj
kv4jdZsFukFNInw9Ux6SdbvRcLAUD55Z+RIiKJirPgHdPaff0QJiX6pc/lRgG8jxkQOSVCyi/XmA
AUJ7/Rn0B2wdbKoPR1y3sfw2k5qGgq8XafjhEW6UA1oNDJ+370kic9aNERjOVWRxniljFEWYu3dq
9sRxIeYqXbHQHaLPbCs2roWSPMdyR1QQv/SuiE15l9X5BKsGd2Xy2a5qsrG+KYfgmYZ6iJ8gnjhP
DxOgWgPxoidOXkHm2zpdg2T6YmUf/yeqOyeNYDzJ1CI0Kl39ATOR8vhqP/fXscW2auBPXZ74o49j
kWxVS5k7zl8ZztU8PIJgLCms+y1E9yuFEFme6Pf0HEOcxUYseOtLyZg00qn3o1s4fb6j41PvYkEe
WNtgnBia6WGHboEXG3SyyuvCveY8c8qJEkI6BHUWxf85NzRp41ItEeuI+RjHuipvuFMp83kJFQTv
NeyOYurHYDIbBcrSvAstr8WMTzbPiGiXItEcdf0IzO/tD4m1EHdeEUk3Jxqg6RPLFDHuNvyKe1lJ
UWB1siJpyCaDUyK2+Pd1PTtxB/ezLa2XpweipPeBNa/LD261bKwB2o6Ofgc9qWPgmL4xma5e8Jiw
E6Y39d7qQaasBV/no+/SQy693cQf1iFmzC9cXhOGR3BD5jRXT5FM06XsY1D2HPzaVCknCbuB0b+v
V/mXdkE5kfdifdesNhQ/1TrMocyjFqPr9tqKRjDPbOXbFM2LrgAImnlktnrIkky6ENqCsE5ifBlW
H7+Zbg0vbjMxIKmDU3VVbhqqfEwhrraOdjDJmJxPtxdvsfnyB6apD6AFsBGjWI79PQrPUyHo5zXI
ml5yHr3TPJNQEN7acpnwE7VqOWL0ls9dqYcT0P4WBhjVCbFqzQoGT/9qIXoGR6psbRuttxCHJpeU
YiGpZCUPG9msbmoC/FfYg2/WN+OCZJJysrxmWNHyWE647cfR54AbxDm92Ia++W15dnkaSpNQXIfK
i7x9IHWiMIXV3IEaighvIY1wQCez/ZSNUAMogVMAPhDcAc/vU0itml/5GQ24pLufNZ132pwDzas3
bxoDS2B1zte+jF9Nw/ACirOcv7g6+dQxxeZUJFjBgVybLxg0wIdTOx667q/O+dfAYcREjbRVFs74
G3pSo778pJ+Q//hECZkce+We3+NQsGBFkxVwXd7rsWyQrxIt/w2E9yQ8uVo9KQ4z0kJlvAcPGrQ6
FHsrDp5vUApfGrPvMrbK440WJr/8MLOiZMwxHGwAmDmDMMkMkBGlyKa0rnNmFrUqCuNG1gyxfFND
msom2823sr2IjyuDSNEyqRTFvdChwEpyYHsKXTAAGLOMvRkoW8CbDJxu91l7IC8QNh7YQgYVCvV7
ld3ZahrVbEYnOXqJlqbZ7wJKeX71Jobuj2sAeAEXrmqrYewVr8FKeHRRJcKCkVr6J4DESwpmCIVu
5J7nrbbUxmTHidqfNUb7hgickdkgG2eBaziUcgP1esuyVvsNBROgP7d5H/jN2himvOdPNeoqekcf
F4cElWkVltcY/rUbRSf16z4YNmR3TvDT4I0+heKGTqpCUx7iEByZZizoiD4/9sw3JrKnPo4SXMUu
6WzdEuNTGbg/xZ8L+0a3GH35Y8G9/v8y5cQqIKrTgMzCoGlTgRhR37/wI7RiEnpepPGCIGkSbk/Z
3Lm2enqTFzUvZxyFC2pGxp5IKMIsWcW5NAYawzG9Xrucoi41VrxHpKm+7uCGeBAq3mG+rMs6J4nR
xktJenJu51eU4Gimt+GdxeZVAYFD8GytTKbEW3Juktl0OkZ5mUhPskrytxGi1D0dBFNpk8tqiEaa
1H+ZUClbwggsBgmwJVtFQR0LU4Y4o645sPhUumKz9EJhPRKaT419hgSuKcqx0vCL8rHNnu2JCIrc
Lo1PDyW31HT1IGgrQMOLqZaBJVJMmQ7YfgPHeNmWXmZ/+zObD69Yt3HbCftpxGdL1vRD4CqwgfLg
BioUWyKEkV6gu0UD1/7/tmajAZOIz22rJJxzy5g78BPPe3douCZWIX+E9/Gy6OWEb6MX9IN31fko
y3C0gFpFs7hRJV5WKxxuJEx3Nurf2z55XGgUMz8zuJMjcEVBLhUz849K4DzObXlWPfExEs5h1qP8
a0rRp+HmSwEu5gBtbQwjGW1fakqEsPmS6I5kIhTx/infogLeFxzRE0c2z8LXi5GUMpv+X6m5qN+j
X8XtRljtAgWZdxZP/NJViE29c6yxM9/J+mRG5Fn4h4BUqIHkjIgLRLNLbt95FektsnUy9SF22GgK
/Y8z28G0DN9wqRMEyxQlpsFrqfWtbCSPVHu9Mdi1HWTbiSts4TaSrEOSt4rRxZFlqE4w2HtvX8PP
eRMlkwlEbrTL6u78vWlrMBRDeVR15Nlll46gsc921y1ccDPKFP7jQS2AbQJ6HT/AVQWc6wQbSyAc
zvEM/M6Mx7fn86NgqC1PcdR7th3a5UZWuMMnQUBB/nyEhZvIuMC2HXkxJyAJO1Qt83fKaZpMJJfG
n5xr4HlfxKhkT+fVb7VbBRyUlTh+jeUjXMxZacBW14BK3AlvwiXbyrfucWdthRaBqh0ArZPvIgWg
4eIiDkJ9+tZ1l4OFOXGlFO0hLwoihb9k/QgOgyfvKr6cRxe24phI9BWbYKLdtqwWVnTvhEkk++LP
TpKBkwPFf4PIF6SFOg/dHPrXWxQoD+EgTr76Ne2F55GxRAviXeYSILIlzBWV/Gg2Y29Nf2ikDZyV
wMhMol0/51Ns8qamhV8g5Na3d0LJ/dL8m5BYOPt6WeCaE1Em2al8RRrkkPhRNsX7MM00AENZK2X2
6TJbjlepZI0Kje2k/HQYzPmn01VPYYkBy7wxzbDzCN8qMP22IRC6QHtvzM2puw2efqY5GFovze3F
JUbNrndl8mC6hvhm1wPsX0rtkflAJd6xMROHz7FXq2rxjjut/oyAwr18Ptf9Tx32Nx09EHAoLJD2
8QaT+mARRMAbWaLxuOK67n8OPHp2amzc+5nIHOBQjeXDm/FB9dF8WA7YYdz8b4EozqxEsrI4Oz7R
OQLvkWnO0VBEjeqOnlhDN40mVeGRTRSfmjwURzwy7j2Hd4AD9BoaUJnEV2XbL39aDgkMvEkIKULi
1h4qVGxBgtz2ypi1PAedAZkCOidcuL3fP0+xO3SB6J6XoQtrHkxz2XtAl2MDPznoRT4HTgcclAyN
zkf8igWjMCxaz4Lt5+J8vLKk6480ZowIWYfHmsi6pBQI0nUtxS1idSay/dRv/L9Liz7nM7ZkUuP3
LJWtAXL6mthi3i7xSXM+sSnmtN+mZIBVixxrlnTVNuFOePJHfTFz2dzz2ur80b5ia4eBD8d1RV2j
DbD4z6A91KYVMJavu2Nai70VJmKP/tK96ys8hsbDl6achv8TrxOhlgy419DlW9Ask4vAmAodaXYr
qnveJRgKiW9xZE3GnuVLjm1ZjiXCMuA5WL7dn+sDvDLt3W+50CDxUdC4Nm7ibTAc6Q+lxxjelDkY
4xfS5d+ZqFrpOuyilu5YKrixsTZ41bj98pjJls1wUzSp/fzWgrglVZnDMm79U0bCgIqS5qIpeCmR
2+DkMjWHo06s/yiG8T3Z9SIcMEFYMjW4LsobfBXVcTIoYhk76XpI/ITkkQYmmdlWN5QStciAXwLV
a2ukz0i8kcP9Dtec2G912EYFBypRQYh3WEyiKsEYnBF47QDa5lsSOwtZqlOPTqqPa/PCjmOOg07M
V9952LC83B+j4fqy1yvlC7GiFjz3aP6nmd7hHMTuFZ+AVL9seeVwbIRVB3nLF70QRRy+TGTa5Qbv
Ui9onY1xeLBqM2MSzOnHxZxOyDIBNRCc04haXk/hccISXqnONQT89wCSqtuTsUC8AZdEyAzfTc+9
OUZ5XfYcaGhruGjL78oLP0EOpwkxMP0WRHoWrcwEPkQyg4yMaFLj/uziPNRzxFMvOrz2C3k20Vo+
2gdD9MTmCNm6UqNsdt08xnW8Z1sEhGR5PesUtz+uU+UPjAdPFP1sh0BZ4UI8jFItfRfL5zIfWPbu
6Xn6RbdedsiOy1fiemSNYm0KOL2xa9zV3Q2kHLxdhtjdP8H6c4et6VfOOwpvEWUZ2UlMBIojtkGz
ChaBOde+LFsnm5zQfzB/WfH5Iy9P60m9h+Hx379Cwsa0hfJMbrgTDCxJ0eMDN+mc0+7joFZC6Qe9
jbQbZf2uIB8JHS4+clN2kGR7z9D5Nac2mvZRmKo4OEQ3z2hzL8Qk8lD18ivnV5gm9tzyRwiWxaD2
Dd70MP+LO2x/SugBiNCklmDKkHxEvD21DyyGI2HwiphFraieARYAzpFvcRTnTzQQ/UjgUvFTeMH+
ZxS7HX0lTNH1kQG8RqNuZHDWihuMAEGqyXjCxK5BnGtml5OhbfECqoLXERfa2zhLRbm+HGfWS3eE
f3xv2lh6EYklJTmpR3ycWFC7DDRi/87+Fz8vaAXnLp4J2mBenecMuj1Uy784e1PG0e9lQqZ0VsrZ
2OY+SwVsU8LyFtECCBPPapWyFbM4ItKde/r1zHJawC85fgwlRUfgO34M5LauC+TmU/Q8oy3+625g
/zXZT80+/tWi1hA+8PeB1bIUibgtzFhXUko3QjrcmZa+isitEj1mNVziU88niCOTnuf5Yaa6Ggck
HDUUaYkac2gra599HGVzMW+cVfAJaG8BMxQiH7rHBA3X+UWsAIdAqyp4qgrTIwoCEa+zuTGeMwhF
0bn705HhoCJxLhCXoypK/lEFnD3Spd8pJkAAVX4rTXnKHdqbbFNW1RE1WM7lI2bplg36tGKAhZSg
qsdrlq1/9nEdmQwvE1tCqRixbPwMRyLpjfS0221tSpKMmmU+ezzmID9LoRwkRcWrWryzI2TKV0qF
j/FyVmVHQ9uQnYRXOSAlzCDwoc+iufd+bDBzSxyHiIi/TKZ/vZpAZqRpv4DIVhlVYHCJd42TdraC
DQFKcoLeFz2+zutRmnnXmk+su/M/5JSXAY9wfrVC03G3tK+VTf+Qgr/Wh4/eKqYoexrqpP2Ashhk
wDyahB95ev+Mq7H5DJI2n4yC82iRL1+w/lPFPKr1AN8Zt/lVpCc6v39iVmsI2GlLRuJGB7cZBQDc
njo4VbPHaE2qRSStei5I/eLqWpfCSLhgIHX3DKvhOv5LbWjTfucUbzG7rqapK1anuAWi5Kamd63H
nYIjA+fgzDUJa2/4sPTgmgld6N/P+vTYLqmM10Cm/ckt0mON3nyTzXkgHdV0ervDmqeuLLGX0StS
hV8vJbg8/Uj04Fv2TgkhsYDzzRieBT8MjAlEQT44t0aTm4Su9cp2fwDvJEViyjIrnHyEd+KHUYPL
Fx7mGRajd+Ud8zHPDqlLEJmCoikYMEq0ea3WCkNBC2IlJVyLIzs4nZqyxBPr5f4hMXT82mjrDAqu
10sL5VcHzZjrslAcimsrr230cbMY6O6AwuRkVY3CY7Iq93dY4GatOhDjpzyV9pr1SuRHXJ8sx0pW
jteQpPDk80m9l+gUOWIQm1XrtjdTDRdIE0kCUrRq1tNcnAaNRXUzQ6jj6nIMagzFe0iQkduIgTA2
6NEuQkjJd0QCTUM4FDjC45Zqip7C/C1MhqTsIdfB3ByWG5yeZswyWXxwe8JitT9oVTl6rfOr+3zg
SsPqIAMQE+olxQ4eZG6G8wzFNX3fbpxZlmGYdiB8/kQIUckzF+BTZdxsZ5tf3BHKaqG4SA5FQ7P/
2Zhjnc3A2bFqWMbzEowamnzrSHZ0P0GD+y0riYqx2RX5hFZGYy7jX+vOslhlQ5Jkev769ii7U46O
AIVedGUeS4HUyOrKJy35MKUGA/+gjztw8GKAQTxN6rMOayfgR4q5QaVEQ03XFOq9HotCqr6p4Sr+
6b3U40rdu3uhCpajzyrqy5gWkgHBvUpYKLQbhodPihtCX/jTjqPPwzDpXCwSzwSzMVI8bSDYDGo8
Jv6C29NutW7/pNDkbcXuoRWppFKFMc3wotGnQgjc4r1iV36jQfwOtHM5X2JzoilfYmugUmqkbyeB
/nE5xRDzGVj49mzH4/H2tNuQu0mFPHmDd2Y+nZITRXJprZA/ZClmbUPz68v8H1nNrJPsRNdXa9RU
DoYM4XsDFy7dxC2Y9nN98wU4xADkeq7GHUCYf9mneX4M6MBaXaiR8J0u7SNEs2dJEFZDTqBOXmys
xJQIBsvqdEeX26fPas2a20v9LKLG/JZnLu64sFZGEq7sWsC9Og0s3SMCESHnEbxk1W0lwYB0+76q
4wEBsRHxuJRCqtCYWFcG1PJHMA1TuDZiH2DiBoq19JObdsSrrr8KLJaZ7oXRJNALBD5UmI8nb19M
JIcvB4AW/Hq4NTPrqF1LTo2qTzZxPVvOScQctTlTLZwFOM04zptPyBslgNEQ1+JCLWq1KZILHZj6
+Kuo8M7Ri2ur6qf5+kYzelKS++ELCh0bjwGlSG3QYXvkCzRr1nC/LPFOAOCSF1lNzM9Te90J+SH3
cXxp0GCZAD/n2+77oHjyd/l8MFYmlcwkfLG6hmNASyu8YpRF8PoaLAIcUmB5x7Mtbt35Sa1wdyZP
0V4SESHGNSg/jmk95mwvMv2He/m7G3qO6g9Fi0YA71TVePN2SFA2xeVLSOn+DwfrQA4RdGZzDW/w
GZqN6WW+geKHZS/SbbU69T0deISTFf+rf70fd3Vrye5QyOs8I2sxaV1I8JpUlDD/uIWntyjCpMGC
Kmj90c+V9ngPtFRm0CzemBJg/aK9CyqUzuOfZPDZUtGf/KY9cp9C71jrRGV7w56gPwZFYJVeUcfa
kG4y2BTfbExRJzCUFbrcAP5AKUpUDMBk592ElyGn4T7V8SHUHLCFcsl+FVnUJvfaFDXDaPSMXQVo
ZYA3l4j1p5N2Bea50oysF3em3J3Xwnv6eJINEPbPG/TAPxg/h68l/QONuU4o2T5om49Sde7qYMdC
CpZw13gWWiULI78cqOiVZWFltIbRdB1HlcTM9CF5SRPF8IG0Y7ABPD9NNPW6HggWYs/FXlgZ4cvd
MpNe6f9Djz/EiSDGotx99X6jsNb113MdnF7BoPg5XF9BbK6DyU1o95oR/ucNcrCBB0am9a4Thwol
ZCFgNTXrj5C15+JNPepXxD2L7J7MJcMEsU9/mHffl+OtW8wV/v1Ai6rTc4VzEkL26dqc8wk33yBn
q1MIb88NxuH7MY/zcXCmqDE7+D6bIXtxuH9naZsBdLXoOSSlmRxWxhjd5PSaOx2QaobG/mgR1c6w
CaDRfpolmuaXRK6OIl8sVMiw0CFQHPG8fB3DsHGGgJb4VebCMW86xwWSgRnP0vxRhJyzEBIEu8/j
uc83GBPwthdNtEqN6J9B7iiGk7wLxdZgrPG6q3kwHLrZjTvyGBgGv69hWI19ywifgE4CK/4P4hy9
Cc8v0guFkofkBpSwwXb284nI1HIIrurU5U5Sum8dVLySj4aeBqqArMLrdWJESCTiHa72BjbrYPx+
bUbLT52k2M7ExKE1908LnoKv1Ohkxzn6FBuL7DrlowS8fch27TlDbtqFaXnygzHFEFbcKwwolQaJ
k41jsKhHtIMDc/CP1JZm126sQS17b23sHvreB9O1gyLrz2YAOsRKdDktsjL73CMoOxN8BFp4FbUC
IplUhTFck62rA+iRMeHzUFvoPKrw8thlePMy1SWg2mSfUcqcYtjkjsvGwTFjRuaMLipVgTQ7PHgO
evtS260faNdr0fIDWid8Buys6mkGpL/65QvduO+GB36kkGm9uxA6/KVcU9YxZmlEVXbq2cUZXw2+
EYDfTsZEMDoyKTlDmLTQN4G2wqfsBeFRo/By9QTd3D5y5XfRUssFC2nXJApfq2YNWAgwwysY5jUn
HvayFqU01BYOceW4IjptEhtjZ6li1XSx5CY+4cbrfMrG8maFy+dfMpLZer/25Ebj/7d1y0i5GdhN
dhN6IDOLJKSqRK9z+PVtSTFnMgTB5UhLKCEzkpIrQDMGJzsboyeLj8g+FeigVhH1LNIXWRvDT/uX
K8a004WELZi+wV1wgjdV6NoUwsSykpvYXZaYDyKqO2SfHX+Cfmh7LSI10QMqzjdOJawG35n8qxIy
YafB/R23p57gUr56QlC5TOT+Jf3VySR/eERLdx5yGMocZS1v2oUbMsiIm/t/7X6W94c1sjFCoyNw
r9OyPPs/EUAUBtp+31sRHow8Tbn7kyCmzJRf6jL2y9ymz8imjIboQxgThprb2Ke5ftavmoJxobih
+mIlJuHEBnLwV6MJ6ntnHTYXazhbAVkysl11WdVrd9Cv1wei97Gvznyr1nD/mrQHMGJZBN4o5b2S
QoLnKd7NeUYQnnx++j6GuYskRzbehujZ24U6Jb6nqlEf5ItSvUpRxbSW2M07zHImzOj8zmtSJXTr
1bUzBacauc158wgDF9bQOOnQ1e6YgJtSxl63iy7XYyZs77sqGvodj8ueP2cYIb/V+qdyn0ShkBSr
eNjHzYrrxaRjGQhUywP898ZmDNJkziFFaQygi5r0RTJug/wIi/DF8pG81I6FblU+niqUfW//i4M+
EyN4b5bi76AQd3Je6Am0m7X1oWe+6sGG5d+eFp2zmTv6/lQrd1Zf0CTAPEFVQREcXMMvJpd3qmHb
e5b38ux4AOD9WMDG0JqydVSO/qI3IGdwJI1nEZWFeMKft0hyHbaf7BrlpjFmbG/AwdOxbXuWa0Dr
CN7MpFf5QGG+Sb6A/SwkLLp6/hoUCtqtHL+UZbtL2T2YOb4VXxnAolT9PGE8dPcoMTmtAIcjFnt7
xzDS40OdOiR6A66TXpz4Rbf64QSu0ogDeISxMA2vMvE4JEQxIGFpSuSexUBqJ6rtB2ueKR6dvxfx
55DYDldgAaQYzhQ1b+eoCuDAiyBAggVI88sVyD+1IbvavdOcxVIrL3GSYWZl4nLpbGZQNCz7/MdM
tpceuHXaKZaLDpoLEsPAc+67XOLDT+FLeZw5HJKqauzT6vCAbOBu3awFfDWWY39fxLhmCzKPuYAd
1zLg0cKOSX9tiDtFCFSLo/SQ4qi4Ru99bui5uyBUkCorQwgoAZCesgsXXDt1ntV1K2G05Lu1vw35
uN28pAKqxZqYsIMWO1ZUcGl+XlIlXxSoQcGetACuoltuQLAgqON83r+TSDXgG+8qoUi8w8LI2FX0
/FVAy0rHm4pI9a4uyW3liqvbb9ebI8j7LEixmiwjgd1/ghRCRZ81d3OqccUHS0QJswS2tgS+NDIU
mwyQmmBBqeknUvLuFdno65G81Sf8CKBVU2Tt+zN+pHGJKkD+jbELvPzK/101tBBVaTdwSrErZ/SR
vGR/Cu6TjC2eNSi9MDz+fSbtDP+CEBpCO6VlXErXZ0VTDq9A7E78rt85Mtswcu/P1hrMDX7gzRQh
DzF7/PMqekaBHcDnkrDWZ0u+d227pDtPEAn9monJQMeDWeUaMjHJJIpwdcl0SGEQ7lnxz8BtiZ+O
tm9uTpdLXT6Q+DYSHMWpTOLbOCYo/TX+OvSuQeLhOlCi4czZ0rKST2Ux6gT17Sb4hAQz4WzU5qQD
Hgbc9Y/gqk66UB/XL+Sg/UxeVY7eObQXRFnCH8Co0ZxBXpQpn0CAzGJKlGsCSODiomOBwALqfSFX
m1qqd5L2oDJ3VXJEp9bZsSyA0LFM6jWPdfWg0FSHjcEprFumvMBxk4lHsF1KEEenPbWcmlyGaHof
Lx016HunmdP+7GzYIrSMU5hizPte+CgbjswrmKt6HKusoXLy5cJ/A/BY3DCIN9ItRiYTm9h0zvzV
l7aRBBDj0rOtapD4O12jFmwyytCvsKPZHu5AADvdM/kmKCyAsl5Kjxr6z0n8pZkOHktQbp2XpH/D
RV1cWvRJ7LPWTLmi6o0mBi39HyTuQK2ZwBp8FH2dap9H7iBETKu4x+n1D2KmUBCHyaJMXowXbPmz
kRNPD66IrgvWQxCffhv2E57rOiQm8F4hyjhZ+6d30mEJp7cJKCbjReuUenCSr5aRUE8FG9W8LK0t
mdtrHu25+QLbZxEbY9NpKoEwutTo3oCGnBWK25j0kjzvChPSgapbMMxKFhw+iSjLNOfJp/KkGsEG
EH7CkZoun1m9G1Q8JPuT4isc94sytP7ML1FN3JXg+2nyapmrB0QE6LIgXjQZwgQCwgh+YsoPSrIc
lCzpJcR/NpoT4YSbn6QGTYJK8hPXOrlqm8DvqwzAxrijhOVk62VELfK+mbfwmkMU6UJJ/4wryekt
gBqT2pKwkf8QtV7aC5m7VrDr/RMhGWB+nX3v7sZHXI2GezrnXYW30Qn8rLoTqZP24NQQibrQGYAm
sz3wteDLNwB0ymiqvqWEpq4PLMPYr9qK5B6AsP47JzxIcDsfY/QbLMTK3W/bDmElYx9mi/6U7GQq
ZmEMJDgz14yMeT5/DBLnv9ASxVPedzQlAKhxpmjgCC1wkwG3JIepWYa6e9J9HSpoR8FqRdTOLiMI
MxZ+y3UQOLGg8NUXQj9jicxpVVyIlfQMIiYo4AhpidJl9/aGRfoIQJ+/gO/gocnd4bZivVszYTCV
PAmZXkte6tczT0EIs+gf93SO3K3Howmd1PQIwRaFGJaWa4NDYX96XKqL15za+Tqb55eVjDW503GN
XhtpYkOiEMmqPgxR8wjM0bpiowmw1zLsOaUzmETx+hFnP6UmUdCVWeo4JNRSQAb14SmZGzy7fcxk
3n0ZsksTaNPzcwcZ/e+6S37RYLvduBr2/JrjSQsrvyJ/vDVoRlf7566fTg1pbtnRK6aAFOWs0B80
DsmjXqtH5SIl3FW9xQQoK9FkyXGut9lA1V6g8gL5N9UIqvBJmFjC37aXEC3qeLuYq24MkASAgna5
fzgAGBnF3j4g/EtpBrVbBRy1wEySD/HZBFTQgrx/itV8byUyVgTV00xLAa25dSLMXBaY5bgAJIEf
Gy3rcC2mgHpIEWZEXxRDxtnOParR5uJ/JKUGJgy2JoxEFKurnrmrtfxhzSe0gU+DKYGjWhTngZ+X
5VgJIlQf2ITHS4a8D+jg+KJUfQg7OSNTbDlB+dlX2dIaZFH96AoIGx95v6wMg6iNpbUmzvAkV7lA
8djZm551stdHIyIzfSvpRtDoUTeLDNVXRjIE2SNlIgiCoONnVPs0Sw7UMVB5+DKfZPIT7xrnGev4
WFMe3GIbWUKVO9SawwZClGYYCnzfoIk0tiRTIm76N68SxCqwZ+lNBRvdqI4P3BfjVSfdBQ9y5jRO
vDgC6sWH0V/WE9tG3rcNkg03Dxj/fzUK4/V3B+8QdmJVA99N2qByQTeBAcvAPHjxKzmZGVMXyvY7
AkLmDywCiI0o7SswQkwgTSbr5sfYm0Gn8bGi+pZzSci9utFV/E//KhRxzi8d6PeBqCmQ9R7wT2UC
wg7H51fFPqUwR2n13KwaBl8dC98gozrxclWRvDmcEltYTRYv6uArFesb2QzegGYU9Xwz3WNVME8j
1BRebPIPQYCgPY2CNWnGIEwo9nrJdveGlqcqq4Ev7C1uZ9rLlv3N+ukRRnou1YcOKztW7HQr+10m
3eSd2+N7aPr29xqytQ3NTawk989J/+IVThXZ7IUbRsOc0oH1q4+suHOQSzCLsRdrvdJCGGGzWzgF
Sv3lb/vEoLNgzt63K0wTksrYPhz5mMAb7OibwzyQ32qKEklc/L2LXQBTau9hv6nb4NDyEX2U+pNf
iPGHNMQ7y73nf1L2HnqfWFeossR3vRmDDcx1aBnMhyZxB2SmmErHWJ2tGFyu+VJEiAr7MoA4cdTg
FhugMLwjhm6hKMir6eJUCoDCmFWE+MYBUfC2z0KeAVgoHi6nlSNyWIhY3X1hEulTHKmSD4VKgK6r
5/uXFtUOa8OaNomjEXZPYltEPnCKgmgEQKl+UYSw3Ga2iMhD9N2f740Hj0gnNiIQKkNz+7U6j67Q
vxGukxFqgSgPN5u6dgvgy1nwXR+D1YwAkW3VPUTyEB1RdT4R9oAqErPOAsz/D2so9kl0Ii61xA27
qA1X/ZNCqRkYbyN3i9ag3xIFD0PKt6YMmFR1a8vX5lnZmXe1lmDRjCfgmfiDRM299b1dvde1qTlQ
luFTzZK0AMUQNvGHlwUN11oFKTBMPTvrSS+adoG+09KdHr85VBip28D74/fMOS4F+xCpG/O18LxU
WZDQE0sflOV3jrHXJulcPtYSYjpAHy6Ksv2cbCRa6Q7YkAxcGqIuJR1Kr0kEtbzcRmfPxdf5VjRd
4brYWtDYYOrsB27BSE0fVWPUqFS0V7gG83du6RpemYeRdJrJQP6p9ExZtF3BiVsumklYqNdud0Su
2Eeq0WO1mhCg8HiAIoeg+KWeTwxRzfFpTFqIiKgMHhEP2MdXSCcn5nV/b080q2/2+1POzVT5bxX/
Msk3KKsV41cmA8qSiNXlOr9h/qu293WPsC03IAa65F8xYMHcnsdr4dHy1P0szowYUybRVID5odkq
VSkhep6tyofU+ZtOlqE+7U8eRxNNqiVgzVXJsFmwsPd6PRfCe5OWYZhZy2EFJ9HPsb2v+LzPiDZ5
w+bi7RfTFN2mop53NcifDPhs6/X48Hd1wjHkrIGcmcK9j41Wy0qFKsiT04tmQ4tePfpqBBYWvTom
wGBDNuqQDUeUgkdoXLlF0ksf7+lv37Ub9NMj1tD7Jw9jxe0qS5IGHe2PYuS+kNOqVHZlmri65mhv
UMRYK5wXvtzgln+9r2o/sj5e2s7EEcViuds9AbwKhd3RKG2MFgx3mrZBTjhjq7EqaN1qv1WgTRVP
hdsdj5f6A5XdP8SNuVNpdN7RtqR3S91XDAFmCriYrFUysQ40+vLS6FV3CWaPeDpFILNjHdDoJ+yT
Ej+V6WhA0Z15fwiYEoMFLUaMbi+uHaE+LxRrTcROAx0cdmdLgg7E13tt1aDEbMMBnNwSdgEIEmaz
QXEQWjo4h4eNmvzCKELMXuQCCAE7Ch5+K6iuQkSx4yfoO6f1ZVgkWVEJ4RPaJULSksgZRrqyQhHb
mqGegtN4A5f6/CZxqLyUmnlLIWtiu1wsWeIcoBk7xrXn4iDtddgmch8gBF0O1qDSETV27Wgu/bWU
4jGgnsSSIjY1I+97Wzed3WGF8vE2WbHNGQzrHMXSM0Gy8T+mEA1OKHpiGVZhsBGCrRxLs274OAHT
inT3XIzrR0EgOPG6NzW/3Sje2o3V3NOxfC8wVlz0HCyA5+SYyMSPEnlIFsJIhxJsGPozscc76i3S
MXk43ZK4IrjK738X5rjzhgMCRgnpy0dzOTwaq/ZO55gX5bL66NjTBUkB88mvXHc1a5kcc62mQoLS
E/WxQcrKkaw9O8pEhuRnp2fNrEZFMBentItzEr4a0Rrt1b9DaREnSIRo9zPSQjNCu5XiyFhy831/
P0/2e1SNeV5JgoPfIJ4u1IYO1DqkgGF2sdiyhOFAKUABbnFF5Q7CUU44s2BHHkvjEKHLP8Rmru9h
ngbcaV/VwfL1v9MC3eE4AgbPSSLtyyQslrBlaBu0EXI8i3gDinqWsGNHZstNRmCLcWdyLQD6v/YW
irjIuLiFYTDzQwpXySg14yj8h/Mqbl1ZihQY9gxY8cGkaX9Yif14z0YCuYM+xVdC7mKkfe2Oxhjk
QTCVW0DnEEMAqzHmzkbciUNDDFMbWGb6PUhVOkbpsi0nx9CWA0ZeJyWiOniGY5CVH/n+97V33ivU
i7rQiBBQr6N1OC4kKh33dS7KpKKgos5rBR1dlyHHbO5tAaGfGPKNVOF1WuKJxTH7z9bXulQQd14V
KVcl7iteJQe7rxb9UfWcvl1XD0TTVkmcos5QOsU+EFGOHQtSjlZPZKaDw1mqLG8kijZ3sdq5PFCp
ZEeeVYfwWCoFkI8WGD7qHe2vDPAsEhCE0iSkTq8kroHg28zkUWzT1QKq6OR29RAh7ohlmwgRr926
AuSu6eVXQQLANgCkQnv1jkkWcVRzBHBHlM7JWEWBFsq0gPpEYH1P0DJHr9rGUF5Vlwo4Zyi9p9U3
Ta5IjJknC3lMFn31SeFLrIAbh2y2Baw/NLi0NzjwMHzlh3yWq1Vgac6O/dVbGvGkBTfYPrF1vLBs
JtQPgjJp7nWCpaQqoAyVmsAbFB4q7YApI0f4UU74SCzv87XCC8dDKd665dotoKowGM8ajUQzRg0t
4SW2xPHYTwN3M4xt61us9HpO4lj7zpOdTQbTHCem7laUjiZYVfuhBlreaq7oya2Qdq3PyEFTM7QG
lBWAnhOp+wa9Cx1DkakAttm+HV6+Il5XpnCCcqIf6ceSPaq4L+rY66dpfuXJn6XLhV9Ckg3mMnyc
TShxOvxFdPq36sI7Pk4j7WZoNFdmzzAiTFJpvIAp5TGfZBsH/nI9cSOeY/vn7eTbmOGUtWDF1qz6
da1JcLrVudZhB1gByGu2LXiMSVc6Zy2MF6QE+zL1wIwmQw8HXZz+9+iLDKwkCs45VUOd9nj6IfKW
MV552Ck1eH46SX8wjhyWwBL2NFLmaU0kQ5c/HsYcElUXQfhOSEoOPbfvOxfEVRnynLl231EWdk6o
A4XZzaYNWYr1f/Ri6B8CyY7bef0oq8lP4Yu6VerOQf04Ee2Xq8Ja+O+eP95IPcvCzErVKdk0B7+y
7gXtGP9IpkdRZ58pb1UdCccbG11emR/Jv9SkCS1g9EQYnL2GlT2+04Hm5EFPqeDO+b+4azpakpUs
jmwP2wlGVGBPl9X9p5wwyauYjtDv04/cSzoPhKeZ1W3qITYtrFssjVt/qPGcP0YozSU+TdIFbfyT
GrDIfVfPq7KBOzFTLnVUsMBJQoVNiqvZtBTtBsk39pYbkJ+5IPKp/lNSCYwF11bgZ2ztY1gVLXDX
WhXfeFM5RfiZTWzvBtEasekjcS2++N+f030MZR9JUsN/5xUOp9Ju/ueH3APlbw7qoNx8/loz964w
K2/XpCQQXzplMgTSXJEPR9WY6UKD01/IFOv9jeuZM5eHgSYvMEl9zMUlxXvdpM0gYwc7a4Rf2oV/
GMNGG56PNBsKjtB0yFlwx4kGmNOgjVWjSJ7/9OKkkxoqj3WujaBpLOfE5FOlMQfoFdGlwLAtjCaN
K13dIRw7GUS6tns6ec+EFzfC0JJu/2GQ5OajzNzOa8K125pUFIrP731RTT2afVA4wqCINt+e8PeC
jXVMOAHIW7l0knV+tQDB63mtT1qg9ETqPyRx29V0TDkJ+f14VHAdJgqB/YstRnquIfM4qG4RNdnT
qtcedRGD1aNkjxyGbeNJlvBT+xndFdZ+NsK0WiK7WWnmrzsUkvdIzGfU5efiAXUGIQKjLB9tcvjy
uF+V84VXVqc3nbiaS6cak59FnNpc5W/JDnz7sxWepAiasGLACrWKKeru52KsKvgu2wN7g4C4kSHy
ovY+hIi7AreFA4HtcY3JDoPpfw+kKpJtY06ssVMH5+qtKpoofrwm2dY1Ly9UeHu5fyN56DzcnVjC
W3QgEjvHHaWbDqXsq+9LVeOexrOjITINq9OWyimQ8vHJnxVb6hGfS+eejemKK86ZRxBPPSLt4Jzl
/bPcYgio10U97Ik8Ik6GfdctRQkeYQPOSckgo+9D/CYuQ836pjvVNnMt8JpDADj9DW2+Vwq4JWLC
p/8vuLQKcYBEQ3UpxYCc2YgYyHTARULMUiNXUMQcGll6WtMDrT3TxrPAS/slSkUjigfVaX46tBu+
US2gvviMTi4QK2Lex/HB9QKOEeHB0vMXY28+eTkMUOQkUrITR2lpbshO0UICl3ldyw7cxhtxjaP6
/6wSxDhKiL7tThH7Pv7+DlO7LApZ/8iO4wZK99jne2BQfF3kxL5f5ddC+xdEXXDDItf+A9utRAb7
3HAKeh3F7jsOv3Na6QoZzK6LcoKnCQ53X08wN3MUbT/8QVt0SS9CZ+6WEWLy1oBgPkrIdGgZ5ika
X6cnTvRhLtZDh70ggLgzZMZNdyWm6kdVEE9LDoohAhCjVI8bjOfmRVhyrgGk4P19L0qGjVFOBX17
HeOnbY8WXm4Bdr5/7y8zJdOMunsPfG2jWuBy/AIjQ+d5DQ2jqPxf5rcLnQQKufaMcRPr9ur6Og6J
R2fGzLAZ9HJU73IJX+gqUz53dQANviySODiq0gSpM1cEsgXrnPEODC5CFw7Tb1oATfjSmq5E2iqX
uP7GzL925tEZtxA7Tp1wd7noY8dJIyN3uVZ4v5FRIxp5XfTBTkcYfRlW/Sc+BOUWAhiTi1cAFLlk
+DNnp8yfHkWDeys/DpxWTjB+VRohKzBqAanzNA9Yd1d4sUP6S3H9B6muK6/vUMUeBFljmHcPru1b
W+8aHfgKKUo/AWgSVWF/Z+fUVVzZ7Qr5ocJNviRvctOx/xKgpYB09RYvrn58C0tcMMQsy8YWpYQ9
7tycgkIXFY7EZI0RFWaGtmtRmAU0NRXiNcuQKbaB+MRlQ8oVyppu01zuStq3M4qbvr61smCYFxnt
Bdo8Nw48eReIMJv4RnB29j3enGAdR/6CuWZlsoJG5j9tSqQqihWsT/23tJuwJF/GLgWz6588KKwJ
SiOzyuLdprgOgpS+Qnp9/Eaoz/hsyaOlmnQhjK0q3OY8zXxe+Qag2kH6uwIoVWabsDhApGVeK1D7
hsqH1PU+aphxg960TSUA4kfJorFfjHpiYewc6pMt5IH5iUDbicoNYTtgPzMQQ/HPUEsRv1eNKhBQ
/aHjCDRXIIAnnwIbFMbqnVyHqtcdDFucy+OfpBCdG83iC6IT6AZ/Hsp31z7cSAkETuPzhY+jsyr4
QeNjiogXfzLkddQV5CUCsz15tGblYF9A47UDaDk9+2o4tAe6SAJuc5a6rDyVMoSrulRwbL/FrGrD
ZFnuCSIGtBzS97ahVr+AVE8Ga6EtytxXwGl8iQ8XHqkdNyyr/u2ZtrBrbYS78ID2fRbA7a6vcAe0
bKWmNm0iGsvokglyzUb0GYyU46932xRbo49TPuPjaRFR/NBhzpODv/CtYZKrYS3uY+xr3waaI+n1
t1/Dl2pa4rdVQSgkjXCfFLG5fFj9Sq0iLBclzhG9Qu2NvsWdmuChiqDszW7xC9ucq2VtOvwkzO+g
2CCnsNLkZQ22KTlsyKU143rZ6Ko1mEGw7X475h6j8IvMopoqjtMStHM53H8UmaO7tuaQN8yNeS6H
jscD2Dt4T9ts6b4N5M1YOTSIuP37ZTdomTWzKpsno9oiUfLLS0tWbZGxrzTjzlCO9qKv5m0zugQr
uOI1bylne/aQPJ6yeJ/dXLR/llXQ4IMKFqDMGEv9wDa/WHL60zr0lVW9Ie3rj+TaXZiNDFH4Og34
jbqpf1pciilcqBDZ3QNSRqFsdvD/Rggdnv5y0mgKubXIF21R7HB4TnXyU/X4J08wvw0CQpktCIN2
T8O31gVSWP6PlU3/jxXumS7uAwVvEA2sJYpXlZZLWhVVcKT0sosF1soBozKZtVHF/OH3BPCKL36y
z8rg1XMrPc3cP60BDzzkFt4/qO4n3VRxKssvpnF0nYltGkErhXNSR/rCmMUn0X62rldjGS7QC3eM
PjBxOz9mGoi4qua4k7RqInCu73gbIRg6eiIIscOXox5KLmBJzgFXcdhvlZh7IoEkPswiqI6/E5kr
LFQ9bIu4wLnnmTUHvsUMV9dTgzf5hMFycIJeH4L/f6BDj0JKibHU3vFddJxlIOFcXHj/ThEv83O0
JUcuzO0xxLao7CYjnDL5BRYjZp+mCuDpoJPJaiweQuHjZLoHhqKOKrwpxfz4Frsh4LoVY8ZGiVr8
wkC6749EdftgDJfsncU+Ov7kqCFEJTOTh3sTWLwL6/zmB8WsWsSE2Ow/GCFJgfkmOPHrbD7CF+Ok
pXDz32PJR2gnXQ87lxET8Jl7/+0bskCM85Hr8/CxEHw+45tMg++CEelRJtUrytqKIoONzRUtrOsG
qCrattzJVBuaB/qo6+z9+8itn73zssB1kQGZV/OHXTZNxEzt9bxxD1MovXovvbWnyku9xwV9CJrO
q5FN1KqMx0RLu2652W+FHMBYdx+jOf7F1NenY6sFIBiUCDWcCwShid0IN+5vsm+HGSPa2tU3VERU
7dXPamJBq9I7/Sx9TxjlEYuLBoP6bgvEhZWy+8vcTF1ZOnien/2nO8wUrZ8rEWSVzu/9doefUPvl
9Xu9nwSiwX0g5c0CCxlKowL0Tcke4ToFdlP7qB7GtMiCXaAzEZ0+mB1WNDxahKE2Q6MWC1m5X4qn
UXoesh4Sl5a1kP9WIBt8QKa7eNk1UctPLvHYzxTt6DIFrNVmHt7AKRTKeoNIWklIpTDtjLyjKyn7
JNqEsx1TLdp6kiVz8kZTxCZJut0A7NUYpDd4YdIyPmvd2DVyk/jY30ZzDbdnNM4TsGJksEfBN2aF
7ZtMFE2Bg124pbF36MtExIPzhwqffy7xEqmyQlh1ftaUcP2BVG5jVeuQgQsQiU+lWzwp4leSsDpS
QMxI5AL3+9Dh/n6tvTQ9Gy2KXjJd9uXj1SSRiOobZIa8IsHQ1TKLTNFGrwf++TwmmQSTdQaIUe3C
6pr3suiEJ7IgNkRpMhUDaFQSSdJnzCTrvaYl/Sdc5fI9SSDHKrHzeDDylWn1vmyZ4Dr/MXKNwUMF
sN5+O8Q/rOJu9cgXA6gy344lujTD715CBaQlZUgj9hE1/oHwaSplfbDyw0j03Imik1cwxmqLR5jE
RiX7aKOj6OByPC4FsirmZFBaIMxu7k3nEnqLj8smah5bUoEL3xR+zh7sJNZ8jAjd8Zu3E6qg/Q+H
LoETDLwZB2Xa6UlzavhsQEZ+KaWLR4rAuIgbppqu+0HduaXyXYudxRgMibYLQnnoUkFPXVaJSgGK
4D+rXMou92CltHZPQ9C0O8AA8eQw2x3WBRZyplH0rnpZQCv8J++Wiifacv1pfZsw7/v+3nMSoOqp
XPE3iYvlZOlGsJqrRtmdUoSyPrPDxYYqb4zJrgOIe3wJ+Pq3DrlqX9QlPgTFq7bnCzP7pwvpBCrH
hHhOuICENBd4GWxqfX//w63WAuBN6AT8Z60tmv0RHI4h1dnp8vkt4NTNQru04s9cab3XDwftEfDE
/F0rg2C0Jb+YiM+35orh33HsGDmMHtvL8tXI2ak8GHYeUu2paiBpKpkgw/odI0hSCYvd2NAqAT2F
yTOhpKGB7BiomjJnIscyE9I0nXyn9xwhVXBpj4Q007ttja0iEY/Bw16q7Nu68582BpsrAOZ5ph34
uOgAjcLi6mwv92arBRDQ88gK0gkhutrBTn0eAIQXnBWrW20VvLAfsX1ExWFgVnBYcH3IBIGNDjXG
HROcoDdv1HGDdfkufUiVuiFaZDndTP8ZyNeZsj7xj6JmxxNX5hdZKXH1SQ4WJkPb4VBi0qvOh/Mb
MROS7uhTF+TMX8zMFYAjNC6TDAugoAL7RmkEk85ORI/U2PrKKWf+iqfuiHbiLk27RCx7WAn8pKr9
dpvZ5PeOpbjouLOhB0G4opGECGOJIe/eWhw/lbw9ex6+9RHB6xvbCDrdEYcNUDJ5arjaQn6PbIyy
WIZOcewNqgMbdL0ni81c6p3T4J2BJf/bgpbq24ADchakg9AY64IKRRuTGRgnVkSsjF526BjUhPkO
CSD7unVDTNw9no1nddktnJns/YCgDvzSCz25eywg/HtI77Z93NZgCJY//lXd7FdOxdgLhDncVo1P
26YYGoxNbQ6EAvTIkRseboM2oPZXtcNO+P7Zzvt0/q4o1oIl3jhRKh0OL42QNnyQYPznw2FJi+Lz
2fWTlgxQQnTgrxCcl0gDcbjgtosmZQiIWL3xBJ8W5Vb9B0Rfm+3KP5sz0r6LwZw7aPNJdlzYIgSp
C6lGD+WSjRhLlx+DZpAGOYJNDkYuILACAbIkeczwvDdlml1w0ZMDt4HR86KCdaPqByE/84EW2mQ0
MF+lTB8+8mr4t/rijHsVsGMRZdKhz5WApnY45U53YEQ/RET6Bh5lTALeI7ImJWkbM+57TMEQqE7S
++W0wpctt8wnWRxXlk8Vg5bSZEJCZv9u0qd89pth/vxBWicxyqa6Tp9kJMQ9EpFIqtYUj6SWOtnq
ZrJ6xoIXzaYie1HcJWZz5ecHaEORaRm1Hlpg4QQhTJDHo719r3nPsm+6V5m0uIhlMyQ3dxs8kh+M
o6mI6FUAsVfGScmUFUFd33m4aERu68JMCSUC8lkKAfCYrqjrgFyaaJ2db9AFygV20kOPDYg4gUBI
qBSfdUXUcxguFGRTRCqwH/mSXdRO87bFancIYNxUhjPUzX/mPSzjTVHIpczNNq3vTlXQUFYf2u1E
i+e04F91nnAwfq8DW6hNLi9/cEXgJtWs75J/qWKATtvzdgorW0+hBfmHfpNrQl4rZqJzkpRS3t2h
QFnaxCakmi46rTm6McnTXZ7J/Qw2QqFTKvZuUTvJaqfHToowbSFw4YQ/h8Erx3KyrvTbgAyNdYai
GzSr8EQtF9E6JnLXyC//6YMQQI2IE2dLfKr4zLGWrguorRiS7yKp+awdEp0P+Mf87G8SIrSX+wTU
CEO5zWLDjLFQESTb54c+Pv+opPBs1HlsIsNVOy0vobMM4oZ7kUFPoCKrki8yTJVbi3n/G9TymKps
tHXFjoEp8kj1Vue0n8eqG5Q4O881BPuKVAhOd86lgBaqwTY5fL3AwaohDMcSCd8aUguo6IGGMern
NSKFh0EzSmKxiJXlWV92sZ88QmcGvx8yZR4wEBsVGvseyiH0c1m0eX2FxRALMmTH2uBc2oxduqBg
+eUJoKMaUoALj8SrObN1GpGLkh2KfnHbWVLap8mqHw/0ZIdDECwPh8pBJx7HFc5WINtuayZdzl9J
GOIlduQH+tbJw9WNozjxTrmIX21l+5VQF3qWVcSvVGhp6C0cSEWsNE6P5N9Dcw7WFOhPQnddD4dM
aVWufxfNM6/K1VG+JMhZavsgBlRVlsyfZ9ab10+VXA4d3Je6WWRbT+OW2T/dpZU3S6nAmNT59RCb
TkstNZTchZxg36x1AURgsbJeS3X5b+QukkLkggCqL7HAXFYBAhFNqaV06sx5Nf48wJp/3vUCIpE7
l+e3kH/gXr3HU2+95D5fGAXziG8ZvYbPnCr92mOtFGiTlNfso8Xv207sfMig/NtigvdB06j7xGLm
KsP5hkFPv2F3HIqXgUUDvHBQ713Eg42sv267cN46Ei9J/rdlb/tydtC/jdj3chhW5/J8Z3polVjg
TNcSk0I3eFJ43nKK9099X67h722EnL38PMN+59nB7JyP8fwqm/iYb3UZ3cUzPeDvXD7PxhJbVUn5
oZUkJbwTKpjvU8FaGB106Gnn4HNs9FhLe02klJxPkTdoMdZqz3GhTuo48nFVR9piSY2rZZh2Lcy6
IR+t2/xRJaNVPeKMJbeah3zCaaMTsCZ/7WSVUESFIguXGJ1lEFcTHmST/wPa/sisewyJhfFByQTE
fGcW9UXAcxJjdq8/E6fTgvorrtQegpaTw/rqpxxYtWvm9Lt0zrFukw1KYmPjPqYbEE3LNGH625LE
5iUUJmFuqpx0hHG9+gb1yr7W3rd5jIeOuHvZ31LP7QGv4Dnd6PL4hngy7tPkOHu1Vft4YSNhi7qR
MCMQEPwgNZEhBeV58VhyZ9C3NK8+bvns6vTteSZkCNIZ/6MtCeDzaRbnR5RP/fsynpLegW1PiDD6
PocetNbxTgVZdkU/xqOOKR7biU0yNnCB94VHvoZDu2gw5WhSqwrujof8+XJxF9taKM8IDCMLrSUf
m80npCgcWc3uMtYwjI3UORiprC1b/I4cIlFM5BnhTCYOGfpgGEKXr62y0KFC7M5WImWd00UiMR3x
RMh6bIE7+DFBSCweV7Sb0ZrlCXANwph+8Sfk8x7G6A5Y5YsEedUfK0sYLa5pyZpDrPf3hZuHzJNG
5NUybsoGNKrTL0GCQ3iKcDrxMkWqKZKl44BamYNH+d5AoR+WUrCFNNsfheS5optYHzv2K7kef9Wt
byqiS9zB0YMXMdY0BBbGyu3d7BWq8zr3pgvloqGV8Q2l140dumbp+Irc8dIAFa2EhJZAtv9eUYQ6
ABkEmbZsx9v1lWrtxIqIj26md0WQ3uoVArTS0qJHA1Mg/BnOqq9QloI55FdwShkXG+3GLfesF3hE
DFjDSX/I5Zr/Tmz/LSFK3M7FrjAFWGMDsTwrADxs+ZSNV3VHbM8QrkFFUrFzoEPZ4UZMzPJAYVZW
LMcWi/tsB4ixprauKSPFrpITv7fpjC/v9ti/1ubR4inDfownhwzqgBG55fYAcaU49VnyGApDLeL/
2XLGX8/SsMvBdj+S3b8tH5x9HPn71v8CJW2I8gPnn0UmJ4aKovHQQ2fATYXQzEJlC3dfXSQLHWu8
HFO6QSTFaAC0+PReUkgt/oL0oj9hP3hxhVqtLluhik7gKOwFysj1fQzsGi0OCief70rkdgEzGZhL
a2C0XzxTBbNViG1gg7A1aF/jUMoYBclLrMqWvyyXdTKBxFhMc0UmJD5cSIdZ0uIOY1xjOZcpi/qW
olc49HrMB6FKiiGAieqrgrPdVFUmATq3274CEd+6+L+n3I2YhhxKjU2A47FsjSTVxiaHHdOi41CW
WCTV1rhiDZgsTQvrGv3s4GVsjblTgy6uZIB4+Gs9VqoO2QBM0kDUvZBr3127C0RJ8QZqDWTGoQS8
LTV7k3+gJD+p8uVTKZN4msA+CidEEPmpc/jmGj/sXwustJz71MGEYssqPeObinvbS6IKCDBa1/ur
C39OXWIenVhXQ2523E8wCrC9LACGAsTi5IxRboM8YuD1s6L3n3vAWc2Sw1Yn/mqAR/vdGVgGf0eF
vbI3qphYCVsbFfOywZ9+zgaqA60yzmmJscVGRJ1SHSD+Yo0SohiNDFQiRo4bEyl8N+YMc3qPPJ+0
HV9e2P3IWyVb11nWn9qJ2AN9Ef+IZB7UkN9Wb7tvgdF5GOUOExuTQK7D1ew+P3rPAZLAQh2XaMcm
acUVPNXW4CpwzadTDCjgaEvWbE+3crlNwvnQfwIDorZlvroGcC8dx1GeImB2E6xM+4UgZEoA9KFm
LGxHRLbVA7PH+SnSFbhe8pF0hB3UrmJ1hKyzDzYuGL1hNUBAcgc03d06feDlNwPc+3B1lI9S0pwU
VpaHJNYSvD3nFTONEMK9lbv0vXMsQG+r+KS/EBF+gaa5eY4cKwv/7vjYD3vfTmwrWtHSbHPJWISe
FF1vZDkKSk9nYjl+nf2oJsvxv4s6nlp6lqE5JuBrwll0KXb7V9dgvGevgL/A5OOPi7fdYQUUBQ5r
NwGil0jAZQUW0ZqgoZNygt7V8IDL3Nbt0ybUpQ6ZFmRelh7qwe0uIKXXBFptlrJ1OmdnQtuXOCZ+
YXQ9JdLd8yOf3pwFfCvFWaPhTiUAXXVUWK7L9CuR0TxpXWCknaYQgOqX1bSIOVFjK7cYWvMTIZUS
dNKPpRP3GeybZagL0KFd6LRqf71Q9ojkigTq/iVO7KgfmsmJGTapKQhKThZgafGNk96XtgX6MqkD
vMaF1OJHpGPY0tC1V3/7o/CQpwXfFo3nHEkghQ+Wji7e9Vo3vCM0/3DW4wLMxIZHvUAiKFTmbA6I
7AKzOrl+U9KlFLkOWab4vIy9rARH4He3yxZ0dhlXBtUwYrxzyoXotL6vsPPDRgkI1klWdzb5CK00
N4VKvTMhAF38O7AiKFePNG7M8Kpta5PaM+ulZVSxzbn339YWnSVCCpY9m5RyhCNz+QL9hRZHuIvp
WDfgKUvplLika/3e/Et3qbPgJdw1QucGA9ERYejIY4kL/Y2Si+1H5nZ3UX4OBEDMbefFrft9/IqN
OFTsv/EXIj/ELCQaRJEypcoiypTFfF2flmakGwlRxCkmCQWFniYgdwV8QHon2HHECdTDvDP95wXQ
L1pxihdVMSLFZiHtsBAeny2T7uXbE8choIDMWEKZrqk2n0LcQYJT6UQSPOz1vV+CLzwvNPOwpooZ
r6eOnBQWtzr23pRmsHcjwF0+ZuIM9a2nYfIwpDW/o1DDTaqqfsy3Qbldp2nfULftUQam8pZ10ET+
9R8iKb0BTPYrSPMuUbShLQq+wVH9iEp64KgbgFE3wUqBxtnWfyJnuDQ327pthcBjh2SwwGo89rcR
GQOWrKBBy40nKkSPMRc6Q+cDKvNTz5vElEnS2n0zTYhUStA4/+NGZ8bYiWGeDXF0oQ42Q/1MzQg+
59soo+PnCWq1w9/2fJ9R/nn/x9kjyCpooqk5K03yNOzy4xh5Z2qSM8YxU8EkEC1g8G7z9pXI0q+z
PxTeM4BjRU+jwjbqQ+MZaOTzVE9+GCySop9ccgZdA0HnwdVIaPpDXhf1foO6lPjVv3C4joxt8h+T
b2UdmmNvITDGYXEtp16nkzaxg7NlRjfAFObMWLMmKXXsNbnl2l2j12IAy/PnOyTZa1gXKLkLwqcc
oF7KqJAnqTiSVh8lH0ntURYVuNR0YgSRQg3klTueuaj4cZ09/EOjLg6QeNo8zBZThG4v/hhQcIJf
0oaupSaGhe4SNqUsZ298jkYfAklt3PqBxDDqEsJsBCmdm5lb+57atuS3mkBkunFCsNHnIxkrOB6z
/2kazYzL5Lm6Kj8QCBO/0O7A1CsA9SmFR2ARizpsZBbX9ksuo5aNkG+yajv0QVgq9SvUkmbDL/9d
+aYLr5ztej3yInMaVSuK64FVXh5vQGldBe0P7mDPxBwFbPji+GwFTy84Lkm9tEPi+1FDetUVzSFB
LLYKNtqxKtv7e5CqJaZYHtIOPwCOYI4fj7rydbpUdBqLs7++cewaZhDTnQB64fFx7fa5pAJtoxTi
5O2UH79TMvWpxp4IRaDeWsjRs8BnD/2E3xORNtvQYJuduNMb2jNlcC3J+XokpxFZUhGW8Cfsxc3J
gRoZnqhIFFP17g5yYVHwES/bQ7qYJKrvjrYATR6IwLvY5oxJug479QnMykEp6Vg+DfnHwLaIReoh
3roicHm1ZRE4x3MmMUAcfldL+FZedvO9lUFqllDviOKmmU9Lg02eMmVtF8csiZ+35eTUc/06B8JP
hdOGYmtqvOpn43WNiwAf+Y8fpQGwle6Bzkqjo39FA4P/IktLrrnvKDqZiTcUsWSmXn8mRkffmEC5
1y7T2sdl8m/lS+w746vbVcI49JqndrSpQkmmWacchV9Rx81/XwyaO9GzeQQjbIubnigu2aQpVHb2
wAxiHjQPsPwkArTT8fzz9oe10lTjaQLokhB3B7qV79Y/kFaZ6XvkQZDFCPoNXDRf3vVlDykzaSQT
ELegvHuRKX89OqtoIuU+ybMkhRmRwmdcPlBrEBpqfP0Nl8g8S3Fi98POFKZBbOpEXZwJ5bILm5UQ
CsF92ijbnyHFq8mHHJdu6Nw9V+UsFHc0zeMl9nUR+1en61JvX3eLtwwsLyXUivWq4S9sLehBcAwx
ChwV+OlTLaPlvi43h9s7gN2FnyPsKBXevGqPY0fRxw/FJDg3fCHdRDeEdMs1qU1F+UNRru/U4PRT
Ex5hIJ3aI+c2ObdFGTUGtffVmql0ZTiZns1sVcrci5V+qNDPccoMNAMOzG+JdjJUU00y8cHFPRt6
KzyOtsJz/Y9uCi128trO+AfpAKQP7OIjBchMpdb70iVPpydZLJi4CNv1VqCSJGlpS5WMPbVoECqX
kEEmxt6g8iPDCoZ3w5JsRn6ccOVOaY6b1o+tTDl+nSbcGacvjlIBHH41rjQIFX3k0TDdFnju/kQ5
ChDLDEHu5nc9bEvCNviKWBV68gKwA+d5J9a4JuV/7LC8uhAAW9JkVTi3uuVE1X0xXZF/SORDicfM
yOzjLO2t3yx9Ickh84S2zMEbskL+SXBwAsNqDcDnaEQ8xdiNpN1I4cT6EUIVBAKYkqogjmtSpmc3
7d96webZvnNhs2lwoIqDgKaD1H6X58lPS79ry8AZtQVzTJ9NgthaZ7vKUJN8wr5vnEbEQjagOyzn
5OYbLka0HOPYTQtVkTN8jUehoLExNHxk247kR7ykycbZyPJK+o/QJl3LMebIs6fJw3wTaN3AaL15
kYTDYj6ZOtkePlCVtaYvNZUwLoqzigOoCFZup7LEvP627DsvC2ciSfjI8/DSIcULSsUCRrowMfcR
M2GCuBHVKt6HmEBFOfYZoETZMt+SG8mOUYnlL5c4nishMw2uzKXlpjvCZOpTbth8o67RVKKuA5nz
PIleQr9mYBZxo8KZGhl/TxSW9Em1VRNKImiRWY3b3X2IxSldBTrJISF420LCyPuwQyjFDaMA76NK
3Q18bFiCK0lDJP6sJVbmEtlCl/tXoyFXKMEbW+75xzAtq0xw7dGqCIqWNCXWkkmcRo5wmYpwu72B
zjxehUYK3iU63f6ltd+EOE81J4TpspnXllgO3T3jLdIDTRaOnkhG+P8rmWyl9TLgqBHrJqPOdLXk
zxFviIUGI/ey3HyAETHKnxm+PsuDnyM20XaMY1xphib3rUdoe/NQPv1JBMUh9B+a3ZjxnrdzGxDo
FPtYyzp5fD7Op3znNf8cv/kGjd/fE8sbNxqoRMpSfU8JAAL+a4an0HWlkkmsITzOn7T3ujvb9+G0
5xpa9SpwK94wl8hUweGVBd/CWjcYTHmuwTziB6SCkh5UB5srjn19Srh1lao86MIzxgQwpXET8ZwF
OY9Oprw11hF/dg/YlIDp1jvHuciBO8d5KZHeq8YsKRAcLxlfRvWWfcO4VkUVPXzNw6yTMrf03z6t
skDO7bs+/34xHj6TENGoWspmTwTU9eBg15VmP7Z5Mu/NwWpbcK+RExrHy557t4kUT+teDcSuLMP+
YQYrbP9FH6VCZ+DF2jaCmP2eFVAi9i4yY+wBRDUJWlgQOgSBkH1eX8WqG77bPKnqlgsJhvlYAJZL
lBtnznQIXbFGJ3XRLnINPS6+Q+01yZ0RDz4B2XHYoZo5YTfecS3Iz2rC6pn78XAAbUC4/kxutddU
WFqrAAetIvetPj4regKtszwm0MjB3Mn+Fn5Dajir4xkt4WeJRgU4epMDLY2HAoqq6Uttfarw1g1/
jPygYeg6fV/ODTndsVo2KVzFn0Sq2m5wcK2VFI69TCISC4cKeBJQB8gnXi+SgwbOPCx169yDTTZ2
ZNk7IjyNn1zj5fiPPZF2Kb0vtb4iSapjplewmSiKnDPGrphfCqeWjAMPJMdjWu6y9O5AV7VGFv+F
ezsprDouXtdEY97EsBw6aFeCYkGvUqdYbF4iYWQ+6J83u4H3+7eTHpvcRZG956AP//DBNfNYCFXD
O6bwKLrbkhmUzp0pCWBg59oLfjLB/9ZBP5FJ8//RC0w6flvSE5/0tZHYjdXiHaruH0jAm04OCNBe
q51Htrf0NyitobhQmf93JErkxgcuVe9Z9vYsFecZnVR754+d40Pnomaza8mPZhH4jhd+28SQvA0K
U+2WFfLu/svJ0jR/37Qux73WLa25SyUClLH2imsddz+z6NxICp6F69dHN9UaekGfvLfNIVg4lS2B
nqSuXitpQbGdTK89XQ5j6EpMTc1peXNq4ilNfqsKlzW58+bjHmuZ2+GgRukw+M7+9AEAVbB+thWq
mSoiimjXpUXJltXV2vNdvE2Bz2cgecwba0AeWcQ1tiKZ+mePODRC7qBQouhif4rOSWfBQEVF+w02
Z08eTZu8Z0RcRUzvIqzVHgRwPNR/JOy5Gfq7Rhk6Kxj3+d1TZka+1WWflQP7fIL4yyjfnd1gK3Pz
qxWIM/NmFGBcGuxw0OKmnwMkB6CfOa+vEP/kxtMs27Cq9FLXdiSD6bxmC5SUscI/R7bSic/3fLC8
XDkOl+wAe0Fan0ULiG8s6RwnV/WkiwtdyvDs4sGV7KSyDqC+dchsBeuMJ8OS9JlPInjEvMs8gsll
ryZoNN9XUEwJhJJ7w4EHaQYt12wgf2KmzJxab6UsVOfSO95zNweUqSfeWvY8aArUrea8yO6dbsS0
mvqc9qdVWprCbknPp3CtVzFsQwiJQApcbrq39dFli2pINtOQMB3AMS0VHfkcxXLT9mCbxEOx8E2L
zeU37oZr/G5YNwD3EGWTzcIa3Out9JU8C9arItPfcgHeBGMfEg2UoRAYDOr8GDCXUAhS6dwKcwny
FaKrCyJmlyU0HL7JSRYnd6oKnXW8BnvTERA1UAxKXS5WHCY5CyAdQzMGHVQe6d2F1VLHcanxqpS/
/jyZC5kmPIkl26Ws7j7dm+zDVYH6IYfIPPkIppJukrj6kKoOO6OVjxzIxlSEKkuwWFMerZFJ/3IC
cN6GX7QHaJ9rOoa7f0Qk2RFIKKt75qdDat6+TsErHvsSBIk9V8p+Nu3TrAg8AeztDzqlH3wTPT5C
qCd3zdb0ZCageJ8+cgiDyNmbSgXq9HuGhZxZv4PFgWc86cFSTclSNpY03BqqhxkyWk3X0Dz6EOWd
th3m3hhNqBboTYRJVE7fYgHBAp3UEMbwscn2hGHFIjKytug1bmB0Cv5lhUfJVMGPWJaSJjlfLa67
RKmGCxnxSKerSVG3UNcjsK/UiZIyAq2UN1Vfv0zyazxWdnH6P+HQIO2a/sKIzCpRBk2biPmjs9Ia
UpBDGQCLz5seDPzkjz+gB+UKj8o05ON3LNHx/5JoqTiJr9+aN5z25BGgX4dePz3ISX7VQQkrHD89
HFlglLN8kDS96ddRoFEFMgx7VZglIoEen2WWpAP9bJcXf/a7Zft3C5NYQLIGPxI+Z2TYOqMu8rSG
4ZBziMU/y1iUEF+yX4qrggJetjTN4XJDvFWiHkbyh53iqMm3cORvOINmTkcaAuG57NHGHyfHfppn
7EsBqtreeTXN0gCiWDomE50I0KMX0Ti197jutjbWzljK788HnKTvvKbwTooyYZDPdfL6hRieSegY
R02NtArxy0IYeuwdsYd/im6r+7IzgSJVzoMJ5ckZS8xUu5wWOQWoJrbw8xJnJd9DA70fdhg3Wcax
TEq5p4ZUAOPzfThj1q4DWzbKpKsGXb0pUMJi25beNgnQzIRzkLETbgGf03ejVIFWWd7h92yYzDOO
Pmglaj+1EEOCYSztNxyhWV92LrMvD+cytWKAacgI+EQOGRWfEfxc3A8g+WMf+9HK1MxQYNLmhX2f
jV9rqAoXnPEnZlmd16G0kNR+ioB5HM58lZZrUxBXw0unY6lpgo5f9ruy2XQ1PO8GJPB2VX8h7wOz
uiLDxaWLQ7YrPR5cT2x7pv+3KFssSvNWIJMw8dHVPgtqiZp8wZMxpiXkOBg06U4MFYExHwG5tHK5
BIHtP71GaF3wtTN3WbZqu1kJYotqg0SJHr1GXwaVKsyzMkhGSSfjhfYXEVRkTLk2G+li4ztaiC5z
GRnBIBp7uYadE5McQ+bu0/gLEsA82ofMDgpGbhAdlUj/6s0kyo+ci4Y8cfy7tN0qNyMjlScz3KSf
nyHfjSpXfakhXGk50fbFxSG7hOieyE4HDDhfOpiW++3RDDFmF6gpZFsp+xyvDGnjBChrDsi8TSf2
iDCplYYsDzkXm4s7i2v1/444low8J3JKXxv0TRrCTThid1aaH5RaB/kYuTgCqdBP+BduW6Y54abN
GKHrppLVDpDGi+44twUaZHHsJZmER5uRXPLhQf+xhVUmvDZwk4FsoC6+yDWcroPzP2Se+pp7l03L
QMILzE9OFM69/Sz7W0gOgx236J9QZFdwzQO96kTT2FMJe7V/YcFBWdcnFHVgoSZSNlpimnpPw9gR
Q34gjj3lLMsCfL/IG01xar46RVerXI2w4sZF6TiUN5fZs3eQJDF6cww8Cjn+SmpZig823nvUjONg
JStcH8wfqg2kdY0qY4tZfhBxgnsbmNwWeyf7KBun5OB+pcvr/Qr3vgU1taQ8wTucxWUGPpg62J3P
NosCFzOentLPYoz/jmrGiwBokYHOkOX9UKeNw7qVddW+PRo7/SQhYfip0TgLKlRujk5YAh0fA8LB
1sGj+1zMXYmjINw/kNgBWxzEdlGqaOd1qfPPL5K7VuwF1ThJpAEkH2j/oTYF+ZvdOpfRRfl/JnVd
9eTUW2EJ4KDyB1bcbLrMfTN5AO8dyRAKrQjXGTtJEeSRTUpwgk99BsNdHIc4B40mzt68dnHwzMKo
jWFq/9YizzXK8X0eNveNuaQxW9SXax1Bg5oGUl6T1vulIn61CnL9b2Mk/fASl05ycsKPWADpm+hA
7T4Q2CqMa2ePB6XS0MbSWleM3k4zPmpp6sAu6JVkFCJhpsSpjtSSnyp59wO9aQ8GjJ6NbncQd5Ps
NwPSxHcPzU0c3fjJl8yEbVRMmZZVEij8/saJKyvHbGdhOjsRqzeeiWEiZNWbaqegYNmYwb9aF3Ft
9eCbdtXV4WSUhnUFrHmrodxk26X0gVOM/mT1NZvkR2JkYgBYDsAmdSPQPGsfu5h5GDhBXnENb0S/
Zjoe/rpWIeqfmTLiftble0eRn9QWIX4j1bCn4eBogI7Np1IMm8eymg8o+HUtRnx4kDIg3wmb7JBP
MtnodSIDFOLx8clTgzCJmpv5zT37oTOVKTUIIo89ZNOirBFUXjHkxIkoEcBIIhemHPQFLUdiqHSk
5ar3FhAie1M79AupZ6Zjt82gLFgG0CRhACKrk2JAO4uhp69YB8lu2/W2tm21B5juf6yMhIjtj9gd
BAhTv7p6fZtyJ9RWAU7dynbAGEdEz1rAfOOdxhh8CQOSqMSqerF8nzbYBmsroc4zBsUbauJzvcvV
KjBoVtYL8CcHhy73aqK+Kgw5h5VUfGksF7VR42rjql7wkRWvRKO7QQZ7zNDbhELkC/D7v/lCvcNa
dRLwUf/1SMe9wmaax3j1t7qVdvX3ld6/cohwxVB1KNfB1qL7kBbKDoHtivx78zKPv4rtOVm69FlX
9xK49RESwja3T/GOe4roK2IRlqjBWrBAvcJba+kr6+OqxOpDBdSppMRWfaQxKZZ6c8fcjIeRleC6
EoPmlMSjTdx0FdipGDP5y4K/6S26HtONqvpWm3iUMNRXKWJWMpB0hwXzT8pHJNKTIowFYPZArxIv
HU+Y5JbitKxvhJfuTuA/Vbz7aJwztdJeskFnDEVSezsPsG+LN2AsyacJ5WuCi6q8rrvgi9xVNuV/
eRqQ2YGNKs7XRGo9/PS4DHUTBj3E0B6+ic//E9fHnH/tOYMD9GSjSGIaXi8siHZvyqprH/aJh0Lv
F0hi7U8DGfhSnuTl8L1KQ6L662s91BRz/qA4RBnO9DJ56OXcMBxntK9aND65cSsxgnzp69GcBBQY
QVMpBKLB3+5+kq3G0r+EzATz8QMCuV4zuxnCG/LIjZva1d4P8H+YE9cYHvTPOGYBP+yAK2PjKTAR
9mYwE9ZiNkzP1Hry2UBRr6Qx5glGKN/X48KK8LzFOW2upZoAROU0PZCf+CEkfB0K2dlfJEXhooKw
jwAde205p0wdYxtyu3e8ckglePG8OSaXWhma2vqkBFWdTc5uaGQfOjWXky3me1/2t07zGpfB4BdW
gtT5EKDHDPa6z9E9gfo+YSSjxy+1dUsO1QWUvqrBo6NfqGPOaDABzYaGogJJTwU3bNT5QS7awJTr
k94J6D3p5Wy/VYmji+dcEzNyzFD2IBF+DaCHYA8fLMB0Mf9z0KIIfN16PDssE0J6Za4yD5xvz9Vh
0yj7nhi3pkodOtGVtIGiaD5st1z8qiFg8dNfyKZ3m9JkBpQeBb8jyjydHepMZqee8PRfCTkQiBSg
oQFiqjZJQnLgPah8dVrRVmObVLpyu3OtRiXdgQI/imnE2Mf++W1TTbVWl5ejbo2qufIE0pySx2/J
5UmvNjQDgwEgBl1X6kPNOXGfUzWEo6LwrEl4ahtkFwPKUD1tC8sqbQeSUVKmd7Hk+i966u0U3+Uc
VbCERkcvt5wAFgqhFvRcERvPEccRgL5kieKcs6T+f6bB4DvQARf4k4yyNmi2xPbAagLwSpOYnWqx
ixCR9J25HZwZaULXyRTvsqulFUWVgWlNoyjTMsjMcWG48oNNOxSLx/SnS/I5HaobHRBrCwV334yy
K7xrUFlwg5nnKVlYMxNSdPKylmompbSUbuV75SKXdc7VQ/iQCVpKfC+GqVNAMkbvoBBoSke4c9SO
aBK+PXcPv0m7V0hINYcmVsxDz49Q+5WLNNJ9mzB6DgmUJduYODQZaKWMowPXygs0S2AkjOyln4m/
mapudN6vWEC9kFyMD58zIcaBoYNUT1IqiJ3ccFUiw8+cG28dNnzeLr+kyJy0tGSym/d9fQoS+vsr
tyAHC9EJGxcDt5NCYqxCWa1d4Xj4K5tN9EseVzavlJ9n8wuwpGXA5ZVP8P0cp1PuZ7A9MPOz7lMM
iW5rsQZFgIY2hkASi+u57AY6GLp0sfVhr3n5bOG4R8rShTKdCA8XlW7DjugqvFkiICZ1O2IVBOcB
eGHJyCQxvnZRg6aPEBf1XCmnl0TRDK8oyzoQgNptryXh7Iz8RGeUWfJ6gQXuZjYvA5kscJq2B7e7
/H7Yh+6rJb1D49PzsQX9jI/ax80zkVRatLHJQvJas2d4IJx5+gBl9vybssLnT5HDXyc/COlMKNhx
+I95heIy7F004wBU5N3Sm3cn11l5IGpeYlHsAFkiD33oIvxjuzCY9I9aWvg2hdp8UNYrkZbZathQ
tHcEi42sQBx5JCjZs/VKhYgDQLVjagkHmaS/Ts94iyUk8MYPRNeB7RHH5u6iEkrC7J2SWoNSbfvd
6yz43k1fq9t/6Vuz704ZTz0dasjDbx049AEyv1+cfytzQN4JKo6/JZlj1VSTRjc/DATaQnSDGy9v
As4ZrhTToDlP50ZAia8gXkvZD+kINxEKhzTmzB1TP/FwHXR1s9lWw6DjP7Bfg+Oesbdb4+lv9qU+
vfJX1AWyL4OYdtFdRbwl0+rbneouP0vPWt6Aaqpy4v9sNIw/wcINNXhrV++Vbi/2UgKXMJ06NxNM
LGSBKNq4z10aqzQglNmlYXT/Dx11/a0PwTbR/YVSnIKXWAp+2ytAHCPoLJwDTrCUjupHJlK4DQqi
71rOWN/qlcxNnDB3DlY0uIeJzQ0qNTNj7x8PnLPMDC+J6//XCIIFJu59etylQn4/WQoRRk5HW/1R
V1W765rsqQtDnphmMBambmmyktpppPQjV6TaDLsVJs0opZa+7+c/HyIprgtUD62d2RrTugCF32Y7
3VUUoKWbFAdC+6wDrlffng07tUBvJgWtuTqvR8fHekH2T93XZgjh17jPUwbHuVZWgn9qo9rBNF8m
NahNO2jm2uCXKwU/oBPtuWgBRYyT05JixQjEP1PKanzDfrW+knYSJcc1cO+g+TGAYpC1aaoyAwH1
QoGk4NHvoKAfuE8wuqKRjue/pq0tn3NBuATParsQDjEKnq76B4o1cULeJFO5YWEzwBenGP9NONQk
KxDpPe7n1uTBeRbGtDshAi+EP/dlxnaA/te+No2Mvq1BAss5eYhgnuV/D5b/++wlnv68cTH2uVaS
qYNIwykXCx4IH/V/uJ4uFHZrABozDyG0Kue2Z5b91u1/axstySJwen6FxkHpQ3hvNkS68zGEFMZB
svMRCy7h22PbKdi3Aa3ve+EnqBXbkPOXLzKkMC77Kk9K6liW8yu7YB+VUjQkbdhpo55qIJ1SGPE9
sCMQfEVo7URkS9WF3V43QESBAPoZPbSWXn/09wfXCgHdv3KtMnGlQuKRJz4dANMVUSvmLg5F/UJm
xRFIxsLtaYjcj/1x6FmFTpdNDwNiw8i9whUTbk/6EfojBMQLxoJ18k+R71pKVPSOWZDMZlz2G8Vp
uNNRSHNBvHMAGfj5AxwPYB2nk7iOEfzaP5OWkfjSVT/eJtSPduhXEfp08QuIZZcsvTGsjQ8zuIiZ
jdN1JSLvyLesdue/cYc0OfZkXl5p30RE2m98pqymeIbBmYbFtuyKHJ27SEzHi2Ze7GDbEHJKOsW8
TdGjEU9pyJjVgc+jrhyTzEjLW1FOv9nEo8oYiD5kafi9fJQyhCL/rdrdryBBiTCCBV1o13pxJhGQ
69sakTqRdqQ4oojlKVYqZ3ihSVEEDGXwMp3nbhl4ahXzYgmQNNRx4m7UzMXQlK+DX+rU01qvJpGJ
vwCEXo6zYm6AwLydNe6ocS0pizkC8Fj36/HWBT1zzfbn4o11YhyM4SqOMzQOtuPwRJLHAruF/Xu5
hljwIO2VfM6PGdqxVZrR05M18jXcBZBbKUxSxYuL42fRz95aEMqEYScuOR8SFnpYY0IcstZ4sl5V
ZZwAA+oaqZ/2zq9Vd5ILziphPRbnNEVLSkBOusT7XtmcxrAbPYXZRvcEcE3TNe3TInHeovKfO+zI
92P2KThWBffuG5IUqfLdbe6RPMG2KTQFqQpEcF5Ya3Ms+alSeCrUC6wdJH4YUWtnuYaL7SOa6R0+
+Z/+v1rCV8465sz7mNHzUULZBiLRRvf5KneBDqurw9B3O2qXoQeP7ziNgqaycO3xGUuTFcVNWhr3
wqThyuxGKEtQs1vRkbhb5NoYWYZrHkUbO8QdPRkWGiL15K+XsSyAZb6gz0DbZGvtZ0p3GOlZNM7V
3bj+u1Ot2vSh/QHy24FiL1Jr8liqj3BlcCWZUATAD57f/B83kPQAzsvMORs7Fh7NqlvA38AvihCg
Tr8R/pqpV6+Jn7kWTz18luAwkC2sUQTXVFxAc16JNFwz1kLP0m50G9dE9O47lhRYtxaeAxAtjbnd
cKhcOQVSWlwOXwJ3oWsYzPUcsNzkoio5PJcpii5Ayd/vBzJG3m24ccOspxG1AN6LQ010NPal+3OD
/IfbFi61uYGmkfP1ZcIeDILh889CNVLFwCnt5CcoE28T7qGKr4sX/mrhTwfk0DQAvbBZJLg65o9M
306Adt80zezpNghB3z2hB2jYlRlGBqwuFyu/bOSmnzb0jGWTvKCUDfb0B7PI0znjNa04zBqZiCsm
n99KQqpAffTsn7+sCBcKaBVIMwM60BW7+2STHifKPdUl3+h50TSVDmftAhbXsdtXnaXA13xVf1Lx
kb3WsAZiNBq7S6D7Bw30/oWmT4Vv8HHR95DjWi02D4FQlgctib6uDt81bLxjjkK8J6pCV3SGeY2b
QohABsfFJh0V6ejOJIt8X+9qLLJB0wqTKCEkW936hoOoN/BX8GSQSu+yQNpp262xAwB6k5KVYu6W
EtBC4ya17pnm14qcDcqkV/m6P8syPVyt6cJ10vXjx5kjBu6KGYPaT+KhFrSX1bmsl6BGzrCssycM
6AsKWCWDR9UBU+tXQFmiN2GXQrkPHdd4fluVV2ee2MzA6CnOSbwJauIf8/QQK2jQWYcf67HPPGnb
YbvF0WCYEo2ECGd6nRLPwpoP3bwvyjQP3WX0Ab3gV3ZtqjxYcV1bQcyXX8M7U1tWRlCI/aMGnXcb
913laf+Am+kToEGkQzY0JCnmVb1n1iksLpxUsI+T/qaYWQ5eHOJkUDvZFaXQP4ytdHaoCscmygDq
M120tj81KAwOiqPF46FjuOqN+mn1z/uBT43j5ObXFCuQkYs1ZnL8UcHRepQ+hxsrvsgct6o/eqMR
Ezz1vLk3lcMn8vf1Wf4DtS/XYPHDtGPK80OhVNaUfM0fysAmlNX+9DgdCms39W9Itk9U8SLSnow2
ymcoG1ND/G4WtUAeOyJmbid+3JcLS3L1cFxuI6zAkaWeKINsuzjq0r7dqKp+MMyhaeC2RWmB+kPk
T1PyeJL1TXEq1PATjEFHPzI6HHvpGgB3fmLHYjBVhr6nf/L1y3O7jLWQyqUvbDLnE6EnLcf4opmW
EUsHb+xkqbBJBJjAfPaNkMW5fvAPE06XLp6Jw2WF9jsd5YJmSuol6jCQ54HZnmgs7bniReQGg/IC
1r5+i8pYAEKRb8VRFbj7y0jSogA28DiRegOXJlrjK5Uiwz5ZclLTrwPg+01QP22hkv+HXP12yIEX
hW9qxWeMuIvttWKrkfQDqLAJptQi7RKFo7q7im7NE767plwQ10z5Kf8KiNtHh/vTexC+gufWikg7
b45RT0pbZjEZEeDDd1ZGTIo8QXO90ed/XudddYi41sCs2S4BkuwgZbs4ByCAMOXZ5URH1udufGXH
Zu4dmP/xdl81X3QR/f+tUajugbuyPyaMMPF5XRk0ilsYaDTXf0GZLEmlJSL85Gli2x90jO0PeBdv
wBmUXYX3sTsGF2X7bnHm3MnM1WTrksjhOQDi9lHrRklc5EW+GitgmtXCyzGjQx0yinY4e2NAPsEG
I6HIHqXCsy52AgH9O0QgGZnjAm2YaaZOtdsCIsHa9G2idDFmRxE/r8dAmaJGvnNtT88JuFb+PaqP
LCT4GimcDCJiTIh6ZWJRug1viWintb0273mlua3Nmc3/WGCngf1rf24dEQxUsvZPl6/kWFEK3WXl
SlQwALih5BKvxgp1+W7vRbtlwzY+OV0iT++OnZ2E4xHWcj3P6jAK0AODjRAUStGXiZD+6EyluJjQ
AcvhoPH9QWn+KskRHELYsOdWhxb644C6ibU0vh6yj48K+s66GMa134AzdLHbGD9uEI/f3WsP1D8g
i20AzPfBbOJ31ef8159bfu530sOFz17gJE0qvk2Bjdpixpv2XiyP+/V1LY/peKApRPteiVuVAHYv
WUCccB2Z54luBTISpBi988qQco9PgCb4EgVTRmchRxdE1sgmhNmAVDY2yZpqckvREwAEne0X7IjI
ChIvmY5w8sUBl0pfLYH5DnQhXBFCdXYgxWtLPA9WACWg2nM2PUptiNXUt+xxRLk0GUsp3bHxrhTO
zrg7FoH6R+ctKf7p09Tl0Eu//CDzeRuM4rCxKdqC5fKpXjxcUIbMwEkcVjnYVsFwOxbDuIV0vjbZ
ItdtVYfmrelg/bJ6oJppH87bJq19qKUYQ8XmYauZYIlezoSCoE4LywsVPsAFVGLUoHsEMbvgVqBV
dbjJTXMczGGOMdPfGmDmWNMIVQlzYDOEUVsQ+jRoACtTAZ0fVRTgMvZkx4GZq00M+bT7B6TzhU8r
JBNVpQXXO3fFEQVCvbIz9UqSrIcdifXhdaW9jNS2Nug4QtaDXGURGIGf09oJzed3yUtu100mGKUa
uvztmnS55MoqYL/Su75uEIgXuNeL7F17ObxG9b/OCdDl/Aq0HBkLch9JiVTgAR/ZUTtknLYIKh9I
sdjkDNXEK2ptFQHVQS5FyjdHVBXf9F5LPNAb4f2SAIyWzvrSBqNtVMrNZH4rEbDBfiL5OdFjcr5E
uwUWeQ1vr5frFrtqi+COkLVMETTp/ZqRM1AUplnR6OOrToXa2iQ/NWmF9wQUtrQqvd3Xv8zuYHjq
xOz57v9oM5jpEglsmWJGUTAMJ/hGVqizD/7Q6v5anOhOjZ340kWUpjgVEA+PlHV7V2mU1yeRBEqh
x6Nsqx6aFSy0hGzv1ht8YlLjdvahK73YaMmMNZmm/Ci9o6SXAJd2yuFBhN05xXXwKnTZZyxANI1s
sj5L//3ZPpDh8BuO2Oek7/r2mUxGiL8p87NQ7pKYzdKtTwhGfiZFBJMkE1noU3Yg0D4P+IJGpwfH
bLLpemCluu/rl1uy8WU4KpLSMrCpLucNrQgXUtKM8DGC4XkTXbbqjLcThSabTtSobi111AS/5Tf5
y0CRWT7cNdYtQ26z4w17kHZ2gzbLYk9V15E4yu3mewEBxLnbQML7HCgCiePTPlAAEvxJ36fe9PbP
iIOezMUoF5rgjEHqOzjXohec67llhj7vX7lwFO/KvnWwXn3Vv2ggTzatLYE+4tH3JNF7DcDMkQ+O
eXSs5o5ZAnm3NHFF//djciO7sY7XNvsRMbBdDN3ioL8YKH3eaV0G/nihGABtdeJSOz6k8AcjHCcX
RKJKm0/cil1nZPgDC2I/KkYpzdXqFHA2oz3dzRY2VS2doKluKkRjI0FSmD4gDpLZPa7fKXa9TMhA
Ih96F2v+E9qjYgXwxEkr9sPv02RhIYOpuAJtYw4QYQaDbACG0l6Nr7y+DT5WWTHg+BXJ3slr4yOd
hsy8p7KiYNizRzRLNdEIGY80wKmYO+iwjbEgbkawis3YtWr+aJ8vaTrAU+TrdMXNoK09R2XR7PCW
rLGyLodaNezF44i75TNJloBJ0sNQD3e6BYAfZgeZ65o736H5BLLam1+qHbzPxBMU0Vpnd/6sBswK
M7YxqP/pj8QM4sS55OJfXI9OQEtjj2n6QjPRoQx/x1eckG4veFdpedI3rJT7L/c+P9mnEnxncuG3
e9kn/zZXupzVsKFn1Ka+VrxCf7sjvl85SnCjMq/2XUAFyAJt9amUwADXXoonianq52dUb3K5v3Jp
IDHpXfRob6Pq4Q4w1NpRv5KMgbOlH8HXjgUckZWyTDX0AXU9fezwlnqhbS8/JxX4EThvcdTeu0GK
NOQilZHmxcX1HA61EEsQ/imJPqYyDafhBrbZc1a29mdOrxteiLAAsKMiLrkp9VByAMGp2F4TuPIW
ikhZKIagFeUXnz6jIyuG77blk0WC7qp3mylfli2LMpK81RpkJLrsvcycFYOb+wm9YzQBREIyzHd3
zjy7drtucQ9fZ7gwfyjWdxBPbdBa2d6Kv18LbZ0PWxHOKmR2ScYfPbrV2pwS/cLwG4isYzH1B8lF
jGaB1NTnoVO+Bl0hFfyGq20FvPv9BP82COzcd3rRWZWtaOoqgF9/JF6hgNwpu9anSc2yrK3IZfz2
+DhFYcmlf5n8ULIrnjASos/qW+G6F5rU1RqwQQCvPt/ip7Ce6MqFhh2jCgmLNBr7G16uOIvEtav6
c4LXojNTmBOIrXQcD0v516W2TcuWKOYBdK0hriywIRRifBboM11DCBL3oUJJV2PRPb93gcFbOZMD
gaDMJj/yqQnaobeWm9uUrhiy1YcVKjnBo+9NfId/qmTNdrOKvkKQHJ3+BjA/Hw6xTBUbcFDcb9XA
TH4B7j+5Vm3F56QQ7qmfKidLJPE91GOeU0HG2AyjcON36UxPwOGFEZYSUgYdvC6U8gsWerGqZ65+
5EEfQ/iB7G/QLLxSm3lJQ5fInrZnr3yRv+QTKRyMsjA5J/ppjKXbQVKLe0NszeW7PeeRqYERvqg0
wzlpLAtbL3s3TFIJtRUgpoPf/stkJcmQAeHmLw7Hy05t0/bWlMEmBTqw/OIBI+E9HUHOSy4oToOC
zAyQrPkP6IAH//sw47BVWTtjBAf+arnrxBQ6yM3IdnR4T6fwLK9QWrHJ1qxuaH+kG8lR/JmJ7NtQ
2ErcFXq9iBWB05aDHXHHX920gm+7WmZusf4STAb5QLAXai7IqTohvv/PQB1ljaIfuUMoPHlO4Rty
kHVHOnr6QkBrFIxRqsWg1F+jMvRYxPVurwHDx3pMXFZihnXDU1Kfr6vIBPFhdarkkDce8kMu2SAe
E+W5LrkJTTbbwEpI2QVX1SuzvhDjSY+SuoK0zKtCddo3UR+as7jlFMMBYfTNIz3il83Lqrkz6Ke6
7MawuUTewwWCIVjyreAkPBmxfrNYcfbHG0DsmtwhgMfvxZtMwL5o1dkaJwVPyys0I9qZHiVRrPuk
OrSi5u08qZgTnBIpxLz906d0N5OK/7F5cdTkGoQZdmQQIlrZt6nQmfcubvD70oB8ipEo3VDC1M0F
GWiHzWgMk0sH0qPuotTugbGFhO1+UEq8mR7tXAzgGhsuCGteKLXdgTBexRPQfcNZZi/+vaPUn2Eo
Eo7znUzdGCgqJlSJ7hFA9ArNsJX8gd2tPiS7d3q0qb5W8WVkXXuAFqIg9z7jvIwNw0y6fpzBiUZD
MH7QhaoyLGdTXuIEOxmB6+6bxPl8ilKRotnJCzvxRqmUaPussN1knmUzYp3UnSzJdGna33iBmKBZ
mLFYWsnkEsezzStQaIbiLLVqjmU/08uFbMHw8920IHzmsjZRH9lLalVE3RuxQTkgYijQxO6cmROv
jFCKgtriK+QEgtKYQgjxdQ6TNsNnaV+VQ23Va/h/w05KBnoPn0cCFcDU0pHajzQpEGgam65LJEVD
nWE6V0u0feD2IAx5q0CkP3iVQPFapx0V5qs0rxfCV//Bt0r2nY+2Or0cAjY4cWpK5PfW2Xa65mbi
/ys/K4Zs6OWxzmcxAUcx6VBZiW1hSBasxp2tm4OiE04ZrIuEx089GEW4+psfOVGH8M0isRzrYwyy
cun86KuXoh24pLbizFkpYcQe0SeRd3cRu4mrqHKpeKH9Nfv9RWXyvtlR/Az+EusDBFaBSFlGl3l9
BhTOXC9ssXBFw+HJ5I1a9zN9Q8Wjx9h6LgVmQewk2lXMXx21fvkGaiSIV89q7dJN2sBYPXwRxhd+
LLCQ4gPKUTtRBIOydbQeAJrdELnthVY8pUfOGgGZYEddlHjLaj+J0N1GuLZloJV8PfbFWgaPf8nv
bt61ykoSiEpIi8rvRBBClgpeyGb1o3rKjh9lJPlbommZ3h0eTmcHZFLenuobfmej1j6o9ZgQyhaJ
I0KgPXxovvCMlu0jiAEw33OiktYPUHOIfIuwX1HOkLFiDkIoMtQGMTgkCBWukGOarrepnmArcjCq
Zgxq5oNWiDfmYO0DBf+EW98JYX3Q9K53PxAepwbQOQ8qanciKjWkPjNAQZyN+erGEnFA1EeYPpxI
O01wb4OezgGR/3vIresFgEJWwfUe19NhcehSHSS2UBrP5+0LzVjEgbxMeH4QBU289s8HB++r+tKg
bhZ2f1ObAf/OzceChB+J3plx/HFcujTHitx5ixjjJ7uMhyH2x+WGyhn/nwdG5Rrfmq+YKJb2CQFM
Wu9skRi5mXejeI3prKAqdpuCblQMGrHxutY6GWt6x0FrZI0bL1ZPIDVRD4ejnbNtu/5TBs0t12IG
MBtQTADDMuk2dboch78GcQqbHozIazbP2WatuIFgpgBMfWWDzcrVGiycqhrUAf34nvUrt1Z+R4WF
4hY7/kEaD2fu+wPj2VVCNLQzmws/Whl7vSB6xWB+3w+FN4HFgnZifJdlojsxVDn8fsAq48/2eMxv
mY70EjBmPZIpuLrcsiLIXIHgzmjlywqURLvc/36OLLU/gXlNWfsaws7Tvc7pjW51+OtZrbuZzdHb
6SprnX44rj+TobbSC6SBE0T6Ow424X5ABrgAyKwwZupGeYk2RGN6lt7Y6AZcQi87CsTK2fS1lfb9
32zE4mEh3pTVHa15TB+9EeDpsp52nW+jRQ8BIq9L2z9/8PfBtWIGwSHa0XvRq6tqQJ/1NGbS/v2U
YHxfYzJqzLi7ni8Bq2QOwnicj9wSjExcmEiG5FbGMrcpU/IT7oesWipSPJGIpko+6zka+9GZ24Ew
0HCvWRD9nnP+bGoNmVf0fRMRMzSifbb8OW8Wcm4GpskIO7kcmET6iwfuVFF/Jvb4pHnPJws49SSB
C6IxklNW1/GENEqcRUzpvxUmz8A8fBZOHbfsI+OeNL5A/UAeuG+jO9IOpahrE1DvwMtSMC7IremZ
OHehcHNb0zY0VApQD2sR2zRURl8pXN0PKTnN0iDmgQlMWBwUztmei7vUjHRs1SBVK0aUQKQniUES
qkS59WwS1C3Obz3LJLmhNgnyAG3AiJN6vDoQoX9XP9AvhVwjiIHrX0zGpwl7nW10mseN2e5NN4ks
uUnOxySM1LdJl9a2Gw9HHpdd9h9f6BUbZi3fOADnEJsZCsDt4W90wwZElWcSlEGjaY0clV/P9E1i
y1hpu1tkCRDvNI+BgM0QK2Z2bB7LAUNyffZvI358lKVPYrkIJq95n7CvnHDm1wjg4SMG0yOfeTUX
J4YcsKFpFoZ8MOtgS5/+QgAw3lX349MwwuC3+tEcHPwZBWG4zLL2Pi+f65MRrA7LOdHyAG59kJWK
3NglHw7tb+KJlxqUc3/8qdK+MFaIprFHc2agzQO9XVWZd2j0pGm+xZ5HGfKVRChWA7vIZN/gvdcB
LgL5fjmuXzgte5I73llLwSa+qecki0zTsR1VvPJ9tGUym7L+eyzt/F44sESFQkGcVCNVz0SSWZCO
Yw2LryAFMj4mmH4B7y9dFg8lg/bKlo9/wgZMS3KvxcJGq4L2yr54VBwOI5r2yTmHMW/O/agvQNd6
PT+FDCCpRVTqXq+aPvynttnEZg8FSS9ISd90Q6UJrInTLA5bT5wINGCGPUsuBLVny8zdA+z7v8Wk
/uydC5ZvvwDkq9tdoXYDeHBVRhRUiJbKpZkj+vcEKnRxGj05/je6c+eu/5u3FC1J7VQLj1m/qMax
2wRUfEDS9XQABokDbfR/HWZ+74OmtXcQaPNwCJtbedNOY5WHPQBJuZ9xSyGey4Q2U7sa60BhtcOh
etfQn+7Xpkcmn/+qwnA9JKwm6sQqgpDU3e4MqBBoBFFrYwgZGPutaqJo8hVWsvOpqbkGMkUrXyFa
85ZqgP8KwRquYQyZdNwJwZg7WC8w358ZBb7dH674hieCZrkOoyS/1lUxpqMGE1VUYQWqvsg9iLO1
R0NfI39k9R+FmHMT2yJG1bTNXdJh3mKR909a2WB/R9I/zLrosieHCIpaowjmxyaWDe7BcxbKsAkO
CQyE36oTslVglI36cU6H9/93bAu5+iIO8qZ92woDTISdxW0MJzko/esUkO0rsZNXDVGixfU7zgfv
MQm1beSTPK2380+lR7QpghWTuJvovTSJ+4NVPU8upxCvJX2QTX+YDfMqB5ciMV3DROFKqUF6u+SB
bcOt8crxNIDsz6luDza4ShTh4imA2yH2PWn8QybKbqU1OXZLE3lsLlfpdetzHO5T+irWJmoQBxDL
sMEAu6Lv/m5kuQDwrQM05LVMsOJd2kFGYdPsrelHfVN6cGnbtU7jKLv4qInXpM+4LNhqW7zDFiO+
GmR9k8sur0o2OJFVNh0cXozPBqJ3ThumHO38Z04CJGXszVmj9Ww8XYYvx+S1H460VPetrtEEUQFy
PprPnWYQMPqvKChKKmDDDrT933p5NVySZRU7LJBkKQGQpb1AMJT18JsA8kMra68HBANX6dp8NXRW
Vcc8DD2Cx3XXCRZjtjSUh88O1OzlEV5oTsidLADhgpNAkwvUxrOWaKXiRIr87R000YHKkR64GC/w
967L92YlnqD7ihGNKywccmH9Spslyg+jU2VOQAvUZ6eFmsV02QLUXb2nKV+oGtf37ukFylDT2mtf
+c61Z635lWbBlUnL2OQWJ52dBw/i1Z7g0GZQkObKsaHtZlfbKYCHqSRQp95RrS5BuG9wINe3fRTb
BrEFnj/ziFaCUAnxtOhpIJ88BOgjfLKCCe+8QnnUhH9qYvnkdhB4an8x8BbgxzXFYK/fuVN9qGZf
ubVsSC6ikMWxUnlfO2F3UGthZ9sj724oZYiQH+AsmZCf2vXu4bpIISFqbsHYIc72pihbE32+hu4B
RMrhj7hYy72tZ2sPmFT2jRI1FMBFfPqy5UkKooRgyr9te3biw2U4rxjwrV4b3YeLRDM3ow9dsbuK
KX4T69W+SFIfDerDD/QsjkGjF70sPv8fHKX9j5mSGUctnvt+ceHXhca7go87FW5TWQvdoYPiTb9+
ZmFQe+eFjRSWTPzqIk28xJvrs27+Ck8qm7y/ir61IBF2jw0Npaj1IG5lZpI9GXilclPVpBPGpl5i
cwdVMLd29OO5JgUl0oOxn4GfnkJFaA6ZYkShzXz3Pa8tfLR1YH8xVjqIfYsyhZgIE3fMEYJzu4pR
5IE+iQ23DpdM4Xvy1MJ0nB1zoonttsxRZGipu4fhSdS9Lavai0hmoOctQbgCHhqnljwbFIpx4mWq
2/IPUmihgmjCHbNXymz0Hs/f6U6VGMbW8wFrFyC8RMryXWtKW4M0PIUw1czw4x6kyv2uVJIHotJ9
GL3D/c4beUKnPye9g6B41QzLUFCVhNni8P0EVjRXQVYtdO2y+Xl8GguRFeTun9u1frZx9QlbblSR
BHMAzzLwqb/mYsfsxFvRuazZSJ7v1TpVdczYSHruJMqlnM5aeTwKj0CLvAe60qhQ8SuZw1xvFEzr
FEY8C7Ol62V+CMqlmxyp+Hh0DoljGS+H3XMJ5EkPPRw1i8hMqaP6uqIuUWlKgAvF//sx9WMRUbT7
wpFZIDhxKbIDdLlOR4StZE8vuCKXsHoT2cTu035iAGOLvFzKRIre5UxI8mcpkn5tz2YMyBDzJ1tP
h+UIJk7Cy0mRU1N8r9vwjHUDek5qN87m48RS65VPSqUhv/LyQfQsT5NhfDRKyoOkSTK1Q2ZmzsMz
C2qG+xxA32GvpKmRb6DU7UPEFwuySgwqp0ccaSBNX7beYE1hG2pY4XVRxFafzRhTCHMB08wb8aet
luf+iTNpS/bD1q9J1kH1yddFDtXxH8WOiRkGDSSlh3I4++pCiZts6No3dtosgQ4eaWB+w+FDAKkQ
HuS3coOjxMIlGnQmjJzsFvqZw/2rslm09ngskC/IT86F1gthrQEBowgTyBZFVAB5Dp1mthkUlFwX
SA/Qla1xLebTS/4yOOe/Bjheps8aEOgPNoVbXS8A9YIxC0GMhc3rHgzTcwcsfbFqrffK/KvYudJL
vPhZE18mqP7pkHaXUEjpLsQRIpp4cMVhs/IITQ5zYO0aMS6DoIXeFee6E7DZoMAIx09wZfpa03qq
Ruy5PVjYFD+K0AQCrFMc2782AsF9TG43PbqMVgbFERsEFX0FyDheNgcuKMC9tQelaGTp4TYAK2iK
Y895jiQRz0oPvbv2ZQ1T3wI164Lr6HisTqGHR6QwmHTzjBg7RM5BZaQjWBtsrod8m+FzbOh7GFgF
eMiaHzyJCHih/uK1vUVUvio1aYeb2BeHlqUEXtsIuZOGwY5rPh3n5ZPfYgu04RqjCdXyRrQPI04t
2ecfgoqlkokYlw93zFRX0Q66JwR75gDjRVCD+xJ+dkuE89vd7kcTipwBLOepRxz8NSj6OFXULdVL
j99GdkM0CXILxBlL7DuJAOBHBgYwmZEss0osodFVbu8G2QVLwiUvsRZs6FeuazF6Oa8QrPuc/EDU
iFj5uOF3WAT2oj+kkQpfJzm/yRzhbpPgDKbNQ9QEtPm7Evvh9zeuFgAEdrdT42H1RGgSKI0zGw5d
NM8yRyXas1xiyjWnT0yfOfpVu64NC4Csq2gelJtjiq9lDToMpzhl2Zqp7uUjJjWYPWbJ5liSn8v6
1UvvuQcYV39wrLXg+RGtvy6KcGpP3IALL35QTkkwVJ4f/eeYHy++hcOmBZRdtQOczPtMDFdoqy3a
ojrHGOfpiGETxnLYs02zVwqPqMNRvLMsUuxEZmbdbfTLLugxEGMgfiuK226AaU76f1uGWztXLyQi
tRLh6JR9v8ajXwF9qxZOhIXZRxGuzjFnmgWOjLcLODysut3/iCZQfyWOZLWajcYcnHMYOrEC/8Os
vm0LVmI+GAbP7QjkrLA0hRnGM9UedeOGQkT0PuztwaxBZsXIIOCj0GWxkqX1KOa/rs4qFxWSDJtd
pO06l+QMFhYIDJnZOPbLUqhvWTGfvkVP3dljbN/AX0UHAy5/ZMeDvCMcMHG+hAIN3xsHmVHQuRtK
BbHgEq57GfVxbz9qRCQ6OuLwj1Jl/s9DHSNkuNLdkcn0WaASQpbrO50KvvXWwz1zqXbmS6x4t9r+
pRgcByuZaSUJmdoJN0I1O8uw+4Wz0xaC0WehG1JXNWZiVEbkufq4QH3CwGP/VKfG8S4TImDmDr0t
OJKc1pcBOXN3XvgmfWWWDtpDcwp7sFH/HZ8eZwjOL/HBMJK9AIH119TVwi5nsD0F4zJ2u2+yPObt
QYJksP9BFSWHrX+2kjUNN7/G8r4Cades768/8JLGe4McEbMoGK8pN1nBLwuNYDInKqCmsTtrgwMG
B+2b1MkANRcsfAiCks9oxOiMhLfYZ1ZRDG8pRDbyhlmJOf+6QI2PLZXyJRGOLWf4TRwhBuDHxYM6
NyUInl8AoXxqtqeLc3yF5KjkYfTPDmeqZdkzBpItEzPaWQsyzwk/ycUZCprK+i42djI31wb78D8K
Jx1JF6XjjrZx80hf6Kt7qw+hFHLYmwjmhjKiVlKzxPyqAShAbZdA1FMHjjHtVdqRqEFNu9YEKsSv
ybRnN5cO3Nb3M0KCZFNMOPA7wxs3bwKiobuDRP1fhdhaPbrGwLrBuRSw0ueeZ72ximLfrStIQ5Ve
fy5jJhQU2Ad981sJoZw43UyUdrcak44LNr35xB9nb4/QHqcaJwRDBa5EgvqsPeh487qd8KNv476C
mMZ8CXpl1sXfm9liJh3tF9g1giO6+v0SE5CKEUCV+eT9bnvrB/0bzrY05fnq9CWTP9Setuhfi8i2
ukvnpWA0c/OhPoYpZWEcBDQPcTqhkebc2D88c2XiBl25ZoQv4lqZPPswgY2AYH3eVo2mv0SKZWql
AHAgHW8+E1DGuhveGl6YU2eKy9taesuc+MCdto+uPG8PygJduGJEsNLFdF+2TxG0Y3W4PFrYvNtT
75dsu3i9yVPCB/AlWrX7aaCoL6jMMq0VsSL2HGA4B9fSWxU=
`protect end_protected

