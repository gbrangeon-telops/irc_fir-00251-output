

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qCd+mYB+5ZYTiHGVPy4TJGVU+1xhFKOwciEzku8LKPbRfJOghBFppfv5cFbq1oB+i1BSYIHhjBHe
eBlHNZ1Z7Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U42W2uzowOkwk+UQGZB3li5Wu+ZZMdyVhWtZ56tkrk6iW89qDlhJBbms676mTh2iLt20rMAIN2QI
nrgBsluV4yEsobcfFOejzkUO7m425YrH0cSwookeI2lEA6QsTIAcBHaB/5shcOjOwrXurevqKKI1
D75XL20Mu1iceA3triU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Nn+1VEi9KmQsJsZi+aKtcGLlFmSquXhfukwVLZNoicIm0aMjF4ddZCMvsg6rFcVwB/qfiEbWhQta
pSDRK+xrjxFlcTBesAmRjUBiW3/wICtAFebLqkLpSTW2uzkYDkrpfNE5IjiANv3SGir2AFafH3k0
HfjDFe0WiziIlRflhOF0bV/y0LPPvcdBpjP9raAJY0w7hoeg+e9PIbHp/PMxlJRxsOwGTLR7XK0o
em6r0lXpVib2l0JQy4vnsZ8th3GiX0bt/UuR0caCktJupeOBsRztdB3gkPhiKQLg0696Wa/3XX9l
8h+H5UXqQy9EN5D0ZK0mIS8tAdwDRw6O0hbAiA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2LRSSTguNLx2WvUvcdH5BTmA+6dHxBZj3mWZxmBysCd90ElOkYpPTP1RgJPbqjpN9tofDDFDarkq
+qbG4SV9hnaX8iB79Zk1+LwdXefyq97462WHnxaG3I/Bff3hJd5X0rJVBnbVgHIqHzt/V8g0jC8o
7m7eoWRXpC5NpNek3W8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MM8YGg7IvNumb+k802doh47T9OSqo/qSgWEpWTgYva1SqSP4phIChk0ewsR6o7XTxZAD05syyzDH
Qfzl5t+Blxw1Jl5F2WrihR2G4uVbXDgvFSouhPopV4gzzwlFtcYs8jnovuVf94AiRDosYHN8WPZW
68LlNRF7Ti2drGO+AuUCHhYE6L1qXzzHwb4c9QJYmemT5/44a67UOyG5CnTiIpfQTpVHSTGdVMr6
z6vPgkB/8JeX7+R+UD1AQWqiV2w63od+aHRP7gt7KRL+kgJ6qCMGiaLr3Wj2C9mfPy61ebJocomY
5wy3s56g63xqQQnm665jsZbjTUelVxQyQI2r1g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9984)
`protect data_block
xNmPkMrRTPnm+b2Rt3jpGjtCg9bx6dTyGrR6BEaNBs9InaXo/UwgU8eQsL5xYZrcA6jy18oIxJuV
QHrssBzWXdWJDZMvovaGQRpxe2TbRz7TomA0pV8U0QJ7uKnS4kxbVS9kzK8xjJxH/pvJk1mDHoyG
9iDEPGeNWMdB0omAeB0bAl8LmRV82S923tqfhAnTbmdUCww2ic3NFF2rz8+Rs8qmpLwTI9xIJRZP
JXBiUsoJgHXlA+ez84mh6+E2vy7N9ix8lFleeZZcWSuf1oTbCMYkj5uP2ZHisq49tdR1mf2/1Yqq
Tbr9QGKx9+IxQF3d8I9DvZT3/YCkxDMoQezgu7hH6P7vtpMQGYn2UtCoHaFXe7F3gYAKrlgpYMhJ
XTo8yUQE9bwwgIij7JnxJWyAFj1VEGKXWMaoPnDRlHZmJw6Lqvyg/xg3pL4zu6commCn6ibyv+FQ
DLS8sdEUrKxNfTNMsL37sgIG5ARTTYuctARSwJRSg4M+Z0VtUkbEC36fvfXEUNGWM9eOiTGcxRdj
x+97ajlKKgpyU9K78XCLmAp6GvSOk1vX8eQspubVTO6HpdxzP6iGGHWf3WonF9tgUQKmJig6+UXW
vm4vOhLebAdeBlfJnoNnKtfl8dMOT6yNbNlT6JIGav+wcbm8PwPiFeY+yHAOvXb6aRkMWKJZVRN+
3h21Oimg1sDEAxN+CzS2eCHgzvmURm/Euxixza7AE6DqXo/7BAXPLAihUY9B7Jf5cpGSCixunXH5
YpUbu/ExHDy61im1EeGCFwvwK81pV8ERy9vK6ybKbqcKrm5aSQGnXT/EzISh5+QzpZp0TUyYTtCZ
LU+tLLMH2OUbMKvs71tymKoEvEplDC91cioISh5hox9PSWEHpF/xwkQf+DqdXwjERT80+fzQmqy3
F4OvfWHr9vVg+uhnPqUJ6d37Uh9tFeHiaeuP40HGkNFsbQPNOKgkSAyEuNIQyifIHb5V8Ga2hw22
h+G4cxTD4jonTeyXCI9uz3fCQyNwEwaHx6Zz3h5DMbVptZz9khaBtiItsdKj+vvIW7FmPXnyhDCB
6bihY2Wss9TrioGsB1MhTbotwotGd3H99ZPVbV+1yNaeiVy2Iypovu7I/D308eHu7L//W3vWhE3I
74RrhF2grSJTT9tmt/S1hj0EVYW2gwdYHwkrkqwwE+ygsir9o3CVZLjHDFSqhJV+KrQaBKXON+Cw
Dt47CYtkste7s4KL0gKAcoLbRJTWert4pZuZinZKDay9bU/rUh1tbEQPvoPoWKg4JacS05mKZ+1H
FhRSaIfh14YwPyme8eO6kpDQh3Cw3qnA1rK3dKBoDTHjCwipf070Z8Fr/jlM2pzxtFww7WYdSRtC
kL670Bkwl/Jvu6lVFRLMLwPb1ghD2j3hcCNwxHp2HFRFCOQGFXP6T6CuvKqhSF9X/+get9oiYycc
lqcsDGs919tbJsBSZ9lJysz7Z+lGnax5LfKu9119MuAmOrXLKrBUJB+Fy1IGcZHvEDgrKcoIABDL
gjfo8vLc4mNy+36AkxOtA28F3GLuDOUA3Xdsf32RCybhNAq2N+4JKaWpuXUy5AU9u4DQtyWgHECS
8LnGP76G8Rgo7x/fO9x0FIA3ytByMfbi4yBOx2fOwienBT7sg3VVcMjzs7Az1UKwUwsKUQSLOCx7
s3CONH+ozRcmWNOsigQJJsLOj/FcKnz24s6CyepesZi+48CLEqfasyW+xptfzKkY5ZUfLEtGcreF
Yh6CBz1hPVczwTmIaArAa5nk2mCsCXLmjJ7o3BCKtCDO01Wx6lEgC4NVhAiSXvumPYUJX9JRSbl7
HxodiEH9OyK/5qg+zBCZ5ZB7q3Fb7SG7MizIL1T6B1a9NFyV0WIV+kbpHWuWg7WpKPuxzv94iVAW
T4d4jqstcuXRGzzuGvBKbV85YmbgwwuJAy0TCznGjVr32HdRI1EqyGmFJqzMeEXnOX6K/j0bVTka
jt/2Vfi8/X8yY/qDVObMO5rZlUIGpi2oF4sGuWY6Mnms5/QSYB4tXJFFr/glHPgH0x+kA2TaE5zm
eGfVXW6gj9ZY0Dksgp+7LIQRhrd8pqpRujYZrnjruR7P0OqccO5Clr4KmKVSIcqzwO4C4a3L66J5
lhhyAx2HNDGCzc4Z8IMhf/cMsC1AvzYbZraESPvQTWCmvdaz1dq5PZwtj7yW3Nl+iFIr+ioEdNQ9
5DS4K4XV5Tt6xNJdbt3xBacmxy7rHUjTFNtvzJ+XPw4T794DHVfxpHs2y2pEPR5wGXTGx4kagCHU
JfZpmpCQ4DETErfJCqebTD25GoId2kRXZ1b5dYNEDAFHv6D3xe336oxV5pggqZZoe6zQ4aSuIFat
ZWdZQzMgEwxLKy9S9k40C3cgALQEy2wj9eUUzrr+cVNeoiD7Ry55RB1jD5dH/+eX7TViiVcBuMCa
oYJwTFnxxi0GINcr4y6/AVY8rlxgULiuoEFpgIIZU5NZpehy/fmqi/14CQy5RBMkmC94IrLPpaaw
y4aZJaIjEiNEfq4Qe6II+7mmw98WC+70o5zqwyojBywQC8IYUsYlkAcgrxmYSq94/EnusfR1y33T
bcHgHCUf57v/bKZuLbtU6xQxWmFgjSG2Evux0IQC4i2MnyJUty9fXTcEbVkesAWnua2wr+rP28Zw
QgBZjMYvWL44dBJEfCj4b9mNQLWkwu2C0ETHtvstpE1h0jOKgQY8pv65RcMpz9esl49Y+i0H+PC2
w6s0n0PmusIyDPxZYo9kVKzHrmcUhFMFPn4mSJwHlgF+5J1uhSCFffsnZwh/GH8t8ftYz2sBnLLx
6O3I42cqxmTXDL2pF7TDuQHTTzDZoWw2ZaB6Pa9q0U3EL5paGHvltNaA698IHT4YeMcSDF18ocOt
Y1HWKKR26AqMW8yq3gNgfeQZywBSLLKlz99eRY5zaIiPUZRf2n7maecMznDQBv3SgmmLtie1pRiI
btw90hTi10gokOE5ji+hNy+F0L+T583MwAOkB4NyOvBLmWzsDpNB2FFf20ZzT3tszoEVSYr+VPyZ
ve5H3yrqeLYU5yqbAL3cFi7kb89fY/nSYsoCg07bwaSkFl4UsktnOorAzlIWb+Z7j3qiSCpX9vS7
Wo0IM1v0tSL13Wtc9XiWqtL4zWkTBrJqU3OWACFFmYowtIFC9QdkRpAT0/X+ShKn5afOKow4TmJi
P9wM9o/G5eA9QBNf6lq6BZUtl+s2KVfkYyYHuZ+pAhTjjAzWX/WXfksiSULAH/qCJttbZBLKhzie
rSGErp6Y2kabzFICyIr60sbZzfZ9lgAWrK9L1hkN9JiSz1ya3FXRivx2ueWw6l6QZyA9TPBf7KyY
l/qWHrTMFxjNGUr9CpeyYdYtUXPRGkpojva3hRQc9ooMo8R5lq+UqZUhkoeutSumjoLac4txuRgw
Cz52XCgBKLZrO6Vdpe4HXGnC+5EJ4PvJRK6Joo4iJIbDjBm6Srhe9dwhfkaGsyILRvUdzYilu5nW
JjlFJE/lh2KxkGlwpVT5xzgFs7M537OOsS0yLi4CO55PJeWwDMSpJdY0xGtiWOkKl+YS6pCAe4y/
APFmY9ySmjSe9jI+Nh9K7eYjrn1pCmY2ua73n4+IZTdpp1JSUGQOzTgD7KJr1XiWWG2W14L8FUXF
9oCYkHwmwFd2/8Xw3JaUGZsG+iF6DFbq/6Ye983zwo8ooh9Nvuf+D4mWIlHxWG1NrhR1x1LAd8o4
aQVwfo5yLTsR3yjv07KfLNBPCuSU54zE419g4VoQ+VRSSde/zVRccSnZ4iqSvDhIgCJBM2kZi+XI
p8FMny8K8cHpg6IdfBI2RINGTynmS+dAA7BRm/UMnchnSUna2Pk3XWYPhH2FknCR3+/bYkLlrI11
/Umhg8XCN3PSkiJ8CFB0ID6kaQw5NAe/7Ei2EQ74ft2lNDQ230jVkbiZNiV4H+feVXJuJUtdbjJV
wtO1l3GrF2iw3Ajl2YaDg/JvpW+FO8ihcVPq2ViywnqC44n3QzIJbdXzbIqPRE/XORGGVtAmaRH5
lzEeYl8CESZ4HItSgZSweHqPn2jAQ5GkW4swt0f9uh35C7NV/L2YMdwgWiZayxgheJA1H9mQGbAI
l4XJiUIKtszuHW86euBrR+CSr8wYrrEJCHUdTEDtFdiMD5D9xn2ZI2Swl9wqs/+1XN8qGcmIIV6z
8yv2/3JjZt5RQdIiXojaPhFHiGdCRPMHIe6vBD2rYXeMO32UrvT10e2wv7/Arpdk0Rx7++bsg/h3
oIwEmk/59GFw3wkWYtcX05sP9veCCmYudZ9IU2uZf0sJI9sN+aqzCYbLZTR4PM3pOtUpOAqj4dYK
ibQvLbKb4293fNvBmYVwe6+i4Qrhv7fOFFqf5c8TxXlsJL0YHDRvqjrUl4axdFkRYY4Yd3aDH4iN
0NYbRB9QyeVRFWFOQmWhcN2IFh8WBsZyRhAQ8b8pHQkfhYNubN75ZJm6kx8fjpujnkJFbMexPJaj
NL6qYAM0kmwp56dh78KGqTrg0EYmseP5dbo1/rUueo6tn+hrbQ/5FB4cfBeUDJAO4Z33OZVbrhZy
0mp0pZ2hFFJPlfrsXstOvNCfYVRVR3Xhjwq1RNjdmf4fQrExNaQUKdnuh2jkbz6rxHBMnG9LBdep
zOlvfSDogyumOjbm/LnvMeJ3qqbZ5iv3zkFgyykINCV3J6ou9t/2KQUg8EnqFlk9OCH86GrS6S4L
1zMmfxhIM792P2dq+pVpfOHufrTmN6pafa3BzkJUVqO0dizDOqizMSt+4RK145CvGl9BykfR53xC
JflNixq7lbD484yLPf4RNY0iYOwg1yhexCSiha4H/Ho7bqBpyvN+wsbdRdpNpGjtX9cVa7la4HfT
9qGhkVuRYRlydDEsvwr/divCgb24WOG9EVftkO8aUBp8GoLwHp8boVJpQaiUPYMRM5sgYxAW0F/5
l0mUi0wEp3uYyu983FY+TgM/MgfJzqDzYs1P5Ao3DKvCA7dS1rFLKBSaxkqxDZYFXJKTuL3l95HZ
jmrQl7qmVd+R5IK3yo0czIJdCQJ4QzDyGm9HKVO/sjNfv0fdjm7vfWcpItnre6FdL8P6AeS10zr2
tdYGtOt8LzNgC5ZMd9iniPRp6mklsmq568FD9GuazHQqzoEaxNkSs3ZPhO9Wt4HkkwpqzyNW0Maz
g1iJXjUQeEVVmZmEMJVwUw9E6A1KO9rLD4RwKE+Wkzg7MveVJlBrhk4hVFy4fFZUn479uG+JKTY8
m8hnU/TC341Qr6MFH92VC4mTB5aHJT1JtWuTuOKsi8z9qPDyrcfmbHW/JFP8h4m4Z22XSLahGyFx
wNO1s96/eooP2F4N0+eKSwcmi0NVe2224IyFWyHXncDafAnD5yIk5fy13KMiqntdpPLSMtWN8Aai
xzQM8OH6k4A6FMwxAle4kM65WziA7PhOPSJ+RnZE49DEAY5ZF5NZ6WrJxNMGZbLkdjcIdSOQm71n
XnIAdnyUon4X0oHkhxWp2HmDz/s//NKXlstdDg2efrmDuLW0v9aVTVARwkdDxAcodg3b8Lq8ICrP
Wd1B3Vv/8eWqPXv0TFTYseLlMeJ6P4tU4MoYsXgtzmwH7SmXMMt56oaeJkiAkh408P1WqYxifY9o
luR1OFM4DCvzXarRgJtbfS7t6k0nUXjgGiOwey1KsZTXrlo8mtOvOUzg/1ajP4WplQFJssQKt5l0
YNHlBzT8oxbmwsou6M7o/RBNXVAzzRR6a19nOACIRbeguatj6psfnJCNZQajRiuU499i0deZP8NT
ZCHLY8D0ztot6yA3m8dWm2cxgVxbCeXuHhhKZ8O+5YxydEBVpa4npjG+s6TskaENWQP5yTjzrQbi
4ZNteZENUycjjLGvtq47UVcSGuVP1WusySZCor3qraiGRHy6tY2jWgTsMsMBLNhwDkY9MIl41EFo
Wr+9XOiU9uFIMOQ8hbESLgCWubKddDM0l2+2osWoUXI2gTBqCySJ1jl77f8nzmwuc19TTylenyex
ult8mW6g9QmPsFRMFg2sGm7HUtj74Oy6pM76/JRGrhj5W1zA761er0lZH8wk1e3FWAB9EyUjfhC1
L2TxAD34QME1tznJAdhs3PqwRlxLJlnzrWHOGEtcv31gmJ06/w2bKwETImeWfoORyo18DAOD33UJ
yxrsielx53rk/rj5f2rx6cZDTryO92LHJgtfwYXJDCn9/vCx1aU7X02finpUP3B0Vy05n0GEQSPs
zx5NiUee+GdE1BleN58KDquUA9so38Wk0HDABwNdQLx3p1sWZZBGB40pd/RSx5R5Sig2cpvPkOGc
legIx0IUjzRQFn3+2GTrENXI3Rjg0Xpcn4C7T8kWwcgMhiNez0VfRE+KQpQqwYukh1NaetLNR39m
KKpfmiTjUSXcPxDDTuZN8Y1+PyRT6s09pjn+I+UA8imbK3aMGB223HyWivszhgPEwEyaBM1Zocbr
2Ma0qPspXC7nptKKAZHTjibTazv/NgIT/iUDDggzBxt2hURl15abpyH0neDOYjnPrXiYBtYLri3c
NWmgy7K55+49/U2STi3Bf2niIXjC5VdvUwI6kTlK2NohZ9yeNVJ2iFZgRdkZQWTohy8Y+PPAtbCc
Z3AVfnl6a+X0XtXwQozkz/ftFsWY06r8vbr44kq+pQZcRpXuCuVVj9Mh7DJgubi686jog9UHljX/
xRPD+4vD+FBNa+li+R8WvWCI2wI2vHbdjJSgdslGmsugJbiyVTeHwgxBqnNtlkHSCJ5kOyxGC00k
toEsKpvlq9l4XR/uSjCDhld0/UmBJnEmbWKDSqnOakv10VtZh5IhIHDkgfqyydW3lcvu6QyftnBK
k6PqzI5OWyjonopnJOJkN2fmncGpQP0+5Bet3iQnNihQFg9JpdcWoOnUe0Na28IeEjaXE5WXS+xf
UBHsNngTwGnRozgMn7kNdXIrwt86SNmBdfkonHiduKnLwoWhzpA1kx/Gc+Bjsyv3gu/icc/Wh8nR
ubPbjlTuEmfqZPR//TT5NLkUr6nvqtZ0soOW3tEoPASCeZuE/rwyXwpm5WX2Q8c8hZVIuv9FwvvU
KVetxGDeyf5KIVyZbUnwPAX+qP5ps4X7Gt0TjfRqvFIEWmR+/RjU4Wnygzgfn4gR/uLmT/i9PRH8
qlObAVllHiMyLL+n537zgyGLv1TooyQGhus+JnFnyjwnIYvj4u2AztIfJhIWeiIE7UNhFRZlT6/W
h9GvtCVMKs/NgXB8hAg3isUVTzNKcn3wMJI75g5MTUqm10WErigmh8jjW1Tdnxlec6rMjnQg8aPD
+tsi5lS1VtRcYTHVMzOIH3xdkDLOrr/VE4mpKiU9FQWRJi2NE1r5LDK0LAoulvsiLaXvB/nwVudb
7d9qfzCIiZOwIkIhulXmVFbnIjUUbKCjFd44y0sSC/Qq/rAK4wJThi/L48prTpDOVBsZTuiGb8U9
hiRzLo2BGEQ/cOhu2STEfqehS7E0JhXTpfwmvgskeFeqB96aW7dOjyik15oNKI6YRDUhyupSaSXr
12xeSZ9pHMBAm+Nk2awNo9hsIcrZNK9/UoenBGrD+prxuKNVSwKDuoRjl6b8PNfdHBVt37q7atSJ
VYvj+J2e5x4TzuqMwlpmWcs10bXHCN+BUIjO73wU3JAtXEG/OrubQAqgNCkFPtUV3pGCpxxt8nYf
iEIAEkkVX3XOZN8URUrZ/XWspfp47MEcpmGQmUkKBS0XkfT0miaC4vIv6DXyujhoc+Os/C873SqL
hwHhJnb2LD4JwFA35kL/2TIpaZ2TQZrV6T3Rp+qM+SHNiUCSQZVbIqFO3ZR4tQbOovapskbNLupY
98KCMxyGgH8t3C6dhetsyWhwxzeqS7KtstNh9UAryxkzF4o+oapiUnHqq+ySA9EygS8jdtfNSZxu
JZd7v7QFnSO6Y7kS2HQTZB9V9gtEfIFZAnECpgqAZdy9Pr/LcWPvhZVIYJAocyK9B9VX5r70EVTM
35eAV22Y3dQ8dHTWOaWd77FYd9EPLpv8TImgA/tbZo4Xd1/vuKYsOHKRcen4UH7DHH2pxiqRcqOR
mcQGjQIfr0p48t8RI+NaJ5iduObv609A6j8h+lxI8EszenMORHPM0iOmX66HhNl7uejX+3mT1Eb/
jf1e28ZcTcYN3bppuIne9KPlwXjQtxCNWBwmBM2aDxtKb8cPRhWe6P2/OqS3g28BPEprTJ22AKwK
EbUs4434sVYPqXlkCItwKthzY7xHkpw8Z55T1W9EYm355Z/M+/97d86JkNWWGewqP942qnh4z5mX
IW3ublxmwV8V1S4gTrZHbXKd/4t94rAB/hE8AmBMpjiGHAsLadMpSVdm+wo2l5TycbOx/zpEhzrv
eVk7N/jDI36Ym4cmyjf5dOvBbJrrktOr6dOVcRvJZuCSMFMS9xFDlKLuFaH6ncs+Di6a64PMoooX
nncCt9+xlCfvW4TGzwAFWwbUTU3cLNp+EcIVU0vykH8XICDfQS/4abA8rRZouiG0ETER3zWLKvNW
Uya7vrwTUQVGq883wAw2c4PK4le2PojqHBPFuQx19fZwNa+3OTh6IOIvHNU3VfbmSAcAneEyzpuh
jVPSZTGQXaPICPiteEza82jfag2AojwlCvw06DOFKT/e6yYrhOZuOIryqigz3mTy4IiZ/72/04Y+
0Q6muhmJUMisUC6arDoktaW/uHqGmnCPYOeuJnShz5w8GEs0RiVx9L26a3+wQ5Zqfo3Q4P3k1WZw
5f/kLLM34FOkGFIbUZK8VM3a3Mz5j709CusSpQCqumFcNnm+R18KN5L5hXNQYfDeBaVNwnazcuf0
CVWIKL0AWZdlHjGDxjeDBpkcAn2yYsAwLlLyNdWemug02oMTfN839mTxdQrf2BHeSzTZyBIE1TWA
mkuB9YuOQaKsbbpbZbW5bD62JC/YOuLbcGx95KW4mnuGLVbooCaPpRTjOQvGVD6JwKq25icNgEDS
VF627mjnjMFi0PyBLa+49MHJnUdp//0NMh+bGgnaLqC8fqmETgJC22EeHl3V5EZojgXhY+jf/Vgt
pItyL4BgaQ0f8sOUihF/dW6vdkhTiO6o0AZ8xXT0wmVs2CR7RAdvGpxUp7CwCCBWqNK0NfjFFhJl
6igbw+jSXOQHOdT2iBdbq14NJpCY6VxmNyJ/MWgUfVwWH69KXGkowI52RDD1zErJZvy3e5O3rSha
U5eV7S4CpDqIFjITbVCGoIB00uCjnhdETwTfOHJYbPw+3Ml2Y0OfhJecgExWEUGQBbmZzJOht+Y4
h7hva76Flxb/9QosTe90wH02zeeZPkYFZe/UV5jmAzB469guBrH2vPqQIB7AcALnVC6Nkb8/MJSq
MXfEXrji9QjY/tIHlmHFMcUKfC2EXq7LVAAC/voNUuhbsN804IJWuzHQl1W8PIyxQuKlemRcqpbm
071JNWYRohrDdAaP6kvl3MX7doREzaE5q8NdSEEyql5h6cFR6Z/9riyut1Qe48ZsoyldqhjmYqik
IG861Yr/cI0u/Y8uRsZN0KwWbK3c6PX5qpxY0pcmLMGE332vV4sDmXsTJEdFXaaXugLI+RaiWvcZ
boeyl34XNRNOAzHUhXklvpfXjsWeFMMHZb0vjF40vbhQJFutk44MAM1/VbE/Ry8h9QdN6mRsTTe1
7JLTQ+adP6MJhU8JAwF/Lh57noorlVkj97McXl0jCgGjybSEkZf6LFk+ua96Yx0BWHuDdXesmZSL
AwRVyr8iPiabsQSCBJAfZbWatnUKsSg8M/5noXk9LE/CJHea6flvBS1d4AUlwsCo+zE8f8Xsp4CC
J1jGDWerhZuZYt0o1p1Sc7qsfXDlQrOv0ns/eytSNfXhklapwxlT75aB+Ikh3iA4DbYqqdEKvx0v
bYXjQCzHAr58LbonUN7Biev+IS8EquGE+PX4irlOAT8RCL7RJYqI+VPwYZOvU2Zq2prxup0Cd2vu
z7qw/WF6uHnEWCsIoYjfxI9qgwfLOQBvDvVpnBK5rLFdXhkNluU8s3IxS29oq9RnLlFeaNvEq6wh
BQVcGe3n7L3F+JAXY/FtEyaojzl0L0bsbzY07m9QFBdXSX3HTsr7vtW6HAuKfIVl259LwyT3WrIq
1TsMiHFEPWTsvywfS0M49FruAxmLx0vDqTQtB4Ae68eskVauea8C1aTD4kYjIIl+4bOvNEVTYVFz
i75RxDEBB7T/e4/9CBNrjk2yO/bfN6F0SHfaO9Ei0UYwd6ZSQuPBvySUelDHmKPmtCO8YfTW7SS+
nTWQMlEsqAqRAxBCnV0n/oPqfU8l6MvQlWC2HkU45CRx83oLS4LO09Q9MnH4XL9t02lDL87djtXM
HjvLjD2zDrHtGr5JO35CD59jXw4E7i95JPIYiEZF0Sqs0Avna57iOKiz+3HqjerdabaPRDHj6pRn
CjFzQM07i6jM/j9jdzHvvQrI3yAq9eHyiAIM9oJo07yik7RP3tju6cJTcEoj/otDSDvmIG6d9jAm
gFBorkYDdY/JAnMP2Rx6c8p9ILxSy+8a2V9bLAkKxTTJ2WYIy44zjqLdLDiKY9U5V0zmP3DrcQyV
KLoJq2/QfxgqyPu+AvRna9XkOuZGt0E6oGeQ29Oy9EJ2EzQqXBsR5kFhkku0WLY4AuMX5bTWwztS
Yuh/bfemxxKn05PV4jUEFWJi5HsX5bmlBR2R0ldxGJbnu4dp3DSHNEo0BgyOx4co4yhJaolUMJPg
Nk6A/J0L4PC4ec3espfcmAS8BAoO0VGiKNK6AI5RhprPxano4oUHF+lDSHk8xkJf1p1yiWBFjDgZ
FbCt68kwhhUyMMF1GoZO6VKtBAoMcJ0a4oaocrwE1ulPf+FNnv+K3w1I10AZgGGcOvImLptiwErb
tETN9t18Qbn3IHdFZfAZbhA/Vs1XGNZE78i9KOtOyEQkGRQYhd6cZDqAog6EnnFxG2bl6vMP52Qz
PQzd+S0xVb3t+g0c2fyeiAqYH8UvFeTLWybLBDqnqV1ES/0Rj9HuqWST/i0S/i7/S02AsHmICJGc
kfb1v3CZJARY6GcGWOKRbcjMy9byO9fMqGr3viYx5hUtmgPjVXK5sd35ydP1h4bQfz8cZ4QjC//M
2ji56f9IMnhQZJvNKeDqaPp1bwSB6NtXCOIIhd9a2GfcgYyRTaFAhfXXLlcDmS2a1qWWCtRsZ4Xp
19KmgBHfO9XTtNkjt53ZThunf2Jh6oiuW/ay7WcbEanIcKyJ+z5pPsi0c6T/Ryd/bG6qI19zL7T1
5h1+iaLiHFX+YQdvwOJJptCyEhNJGJ7nF59Xuu4qH+SZiUoQHHS74HjwO9BuZTLxBTlg2DjR6/gL
pzXZLViNHbk7Qmm7Nf5ybt0qbqgG5WH82oM1CScMIF5SUe7ASB/LCpjY1GKPAef/ZSVGIHZ1xlg+
UrKJ/6iIj5fRv1UK0A7OQUKk/n28PQqE3xdqVQ9NKcNoml/kkYoWc2u37beeqtvRpWI/F6gJhLXD
oZj8lITqO4Z6t0ye21NhwFYzNesR7DZboVWuD0GZWoN5hr4hbPTZtBna8lZYPH1nWOoMxj4AdKMM
STcyo3FMYlkmqxasqTdqSn+Aqa1i8k3+XDbqBpb99a7BsO97n+Ajg/b7nbexAkZCtlvrlNd4Ejt1
CqOtGIuu2z57JPf8zBSQuJiSrhtvB4mlr/4IZP+MkEN/nmPNesjKqVcfzVpbvE1cb/4FMyYWo73P
5f6aYMzHwtY4RzH6AefOIZQ9Om+Je6Zr7hDzWHbBVi5vJqH00ZMiUHLr3/dz+72J6U8yv+I53Bld
c7yvD0/rAdFM+iwHSsiXs1mlcpFEQ4TIk/UJqZgQwFU+WhfQx7MZjS70ewcG06+g1wQvWiz9nGvl
jwxH8j5+7hYvvq+J7ozf+hdN9y/vmGnYGzkP6YKqP1pUykdioD63rLglQtrQDmh+noPrej43lufe
nkRmaS9qEIrHMAM8I9R8rgSdesrCu/mN6gjTjinA1NPHWlfzI24d9wpBlAevq5lRKoPAozf4vCjc
ZQTflXiDO5NFs/3SBpi1gA2fXzCah+OuRKZ474wtf2slx0OoLaJSl5kBKzfoOPn3d0bnffYztxN4
u23uEFfbBzcU7MQXMeV7kLW4pUNOPdL41uoJwDNyNLvMrmF89Wl/B27eaoJwMO8wBiN1ZAJHsq/9
yDfHKNVxSdDwW8jqtmPzp70548wl8SxQ131SYEEI1u9i0SQsKjhAInznG093UEvAADNGAcDktkX3
i3CvhWelCYYsXyaOURsEK7twwwPbmtO93YtKXcH9G7Dbte7QjzESls9R0AWgwePA71g+JdIF6zL+
DNe4P8VuBlVh6+SpH9UhyYWGx7j0iwHXIElaIIDPR3dvt0K+Mb0sgkGlzjnN9tQxKDkM18zQAYCi
f2nlCXoNsPNWvsSezzmae6xFx7XTBGW4WIhxwry+S580+j776ViA92OOmtPjqD1Spu06JpPVE2m8
MEbBo9spzWlHQ7IjTF8B47R4A3/6rDEmcNRonOiVwRA9DZp98iWl4NDBEMbvBLLfL4K2nnlvmti2
3u8FkJ+lae1Z0J0hxuyvclbxm4zN2d4NckVTZCUWhRLCqhMRrqx9+hqxbYek6Aeu+ihSYe3LOpOF
fFQae0wrBsSD9/gLoEdX4Hq0XiZmJD+yxs60v3yj98fGOXsUtqDJxglkH/e3Dg/v4HfMu5p1V0jp
HvnlLulHVqsUK475YYw2FNtWzmmlOStTIB8PvglQJlaIPm7ZwUUBI6UxAS485r/3arvm2ih3zUl/
cjc2T2cN7ofXFcMu6Ab8xSLYFHOTQv87jpVnALH/PyM/z1sVtvjewJJ7osr1xpmFVsuOKpKbX72n
7PSMuIhapSK/kUEZgzPtItesk4tG3sEOM6N++1HboLVA8bFPUE7XU2fYUZ0GPSd7kcwhPoHg7zcf
MbwCUidak8Qd3j3Lb3oja8Rf99BEu9+TaetHeuOdXpYVPudFe4L63svDHLSqAhjGJgiTJT7bh5lU
gv7J+cOgtEMDghU3GaIv5ChNnRi3TXa4T8kWdOd3kGu4K4c22M/DLp8ZT7vKf8kj8MC/mO5J1HJT
Vcg9ho/yTrXqzaLlj937w9T6vGU2K0Eq0WKhnDs4om4SGxDns4bXM24M4pbJJO6uMXGqRID+qtNZ
qaEVWKQk2JbLUdq96XSwjtsJQGEweUjmBjqj1pDld9oJwl00dzqNmfv6EOd3HDHRf0GaksDKiZ/U
2z12Zamj4/5gOXM2o4zCT1lGa8jAVt3rUj4O9BuJODrHJ1sfgW9no0TyqBnadIQM4QL9IGubQ7lD
kpfxUX3YCFid
`protect end_protected

