

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Zt+Kvzwu2Ua/vrjhNueC6ZHFBDEZvqw7CYHtLwQCcRpSvR8qcFedNcWPERpPju3eJt3nf1a3JFkv
PrBPNZe2dg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BgYona2Iv/0k72I3J2JPeYuzuEtaXjhj+ZWCoU9nVssKXxrxRKdrDHt5tFvberHeN9tDv53k+E0+
zSJEc8s7HUTXqNlaEROAMDRbOb7ChasXXdVxfl3WOvXTlUGfsx+NSKJ4/HfkR4Zaiz3A3zH3MCLl
LSzFeWSNT1Mt1+XG8HU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FzDw40mQxR9kpm1uxLfUoItwH6249dxMvWlSzzE19zJKjsyLJvf8oLgoShFkGPrtSiP79qKNxcUe
hzH0hyrZBcM+hC6bI6Mi60dC4BhdqclOgz1qMMvUNpZqrzZ5JB+kSMGHVFW8GUXvnFCCxYuu5mP/
ywkJGUeSDVEZY2th7ObJJlKEA7icdJ5tzO8g4W6w2f+MHJPOeHFy+SupHzB+1djuSlirLlm4nhaI
hraNZ0zRKoeVe6z0EIEqhB9JNsFNiC91BziwCnpzBdkOsKtsrb3RxMWbRRWbmc0XLssKg5Ki5yKr
zZaZTZk48RIng0NJRYTCGlINVIuaWueM3WuBUQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gVm/uXv2qQX1H4bUmXuUswxUb0GUskWeA1MPfdTQVCi9Xt+VdX6mOhlgO6EFKXSas+dhLpimNzTK
aBHFEULIiJVFga1QEdJchUQ/rBMO2ShyfVm62wP8vvP25+deZ0Ac63uVlMRNhE68fori8KTc3x2X
Z6Nr7gpu2y0w16PhA7E=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UyIHMrvI7wZyM6hLJ4gE4jKiSWW2iEuHADz2BcA+kHWTu+vXmBlODWfGdNNdgy52INFMV1nxlqnJ
XDvv73yssq80S34n064XoTXJBVIQ+OApIu1S7Z1OlLjdyiOtUW3Rq9q1U3A+hwbuiZ1x4LA5dZoj
5xr1PfS7YeIFNi86pALVL/xngSOmrya7h0pb27Yqn1ZWp+ZFU4zxAnMBdh6smb7IVFLN7MVgfSOU
BFsRwVHyMW6sC4c5q5LyBHJsVE7Cty+4Vqow0WWDEITa8OtbnNcM2JZrP1+VHJVzH4AYNHP/h5/v
rWvTg/dH3ZrlceYDFRqzQnHfQLNZHJkGerETEw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 42448)
`protect data_block
EG11/hpgGfeERgfBxueBbFQdS4n7XdvAhxQwjCQiwlT7FG0C2SLYOGKPFT+Ol/ailrocfUmjgXPp
1kC4IVebyBmPf95Q96ynUgQe0pVbyUPUpTooGN/9pvm0vqH5ccvw36+lOSbeWrZILzPk9zNDbBMw
MZbaPo5WTYLS16eGoXVB3DfoUpOnMhEOJ0eK0TGuzZgYmizYWSMYmaWdUw9mKAGMmzy/P6yqh5U4
vVIePRVuFW/28xMWXqkwJyPDaQW/BSRp1xonSl6fdedggJdxmlIQTSi4UMWhT9lK5nVzuA7zJh5D
JKKZnyZgqZxWb5y+SXIt1PzBR0fH10ir5od4eiGlenc9njYm6v+0j9ZoJDn9euuY3uQje4o09sey
oOUcQFXo6mHn9l5c4kaOFXXkpxdYhdXg8Hz4+E9pNQIgL35ck1F5iGuDArv83CX/gc+S54HpiyDC
F3LBOhXAwV901Xjn64Crlw0yNYFbDoxjV2X4j//GBxHjpE0rKrFRp7JGD73cMj+2rh2W3rSCAQ56
6jqkCFhPNjfuJ+gGicX23srS8QqPlpce2lhthLjXqWPU7ki8Ud+DzIJryCJJKkK/eAE/atI04HlI
rsNcAr6fKKWMglERndG6l11/fQVjrlDmRpKHO5/cVmjoL++JoJ1zmNX0L0Q6JnMehW9lWSNOfaH6
HPVNLigoE0atW5GZmUwavmmyWnxXPiRGrxaIcY8Gb7/HFSMxO8o6VNKrs7lJQZQB/HjBBKzU2E3+
U/6XJNUibnKgjgQCbngy7Bo/Urt0+EGLgnqPhueUZo7Bf/rfeLZ7mbZem00uBGbZ+NiFF5VrLxPf
15uK1H9SY2yN0MbYT1TsRGLiG8FLds5QWxZzz9OBB1q+FG7Z4PAeR9snudNUJ/9OY6hDc6p62gIa
xETQqqxGqsvfzl1DqbgrqOL2d/vOSuz/OGIqjEbz0OjnMjd1Z6/0SZ1jPI5Ap06sdyjULEKpRxYt
Ga2X4Ht4Auk49QjZcPXAj4D2Ak6smgut3LtRbozqkOr5fcXxQDSx8ToSpbsZDz5BUY1wGlS6oeTH
OtVYlrRu2Gnf5lndcghdbmbNt3gGRudhs/826U/pJlYb3ZUjow2NXOWJ5ZoIEzZpMZQwzfI2j0i2
5SGo4ItILpVFibHQeKPJqbkCjuxBRn05vsTiVECTGwCSe6Bc+3wAUmeZ84cuq/H9A5N0CPd5JDD/
BIs5hHHQNgANmRNEJgmWFgAE5hoZhK1UyHigWSbHhiMsKrJrzbTDvbyZrSv4BGt7wG3OZKMhLcR9
gzwZrRHjMqktbKiI2qFq1/m3lbjnw+JTuIpdmVvA6CHyl7T/ZOVTI8rWhMrLTGVpNGC2T5sHbcZO
RrsLU6Qi+lwlbCsFpOYl/jwWJkOMxqetSMAIIIUYpcVniUdIst4zXtgIT8EhPunW4hWn4rEUJ1lQ
t+gNuNAI/oRTP2jq++OkKo7gwZk4Kvx368CpgSBE9DdvNKQReyL28q7/hIqi5qaiDJPPgG/x1oxj
wUUre57EWSpEGeIIW5nMkexyTg6ciZgqhgRw0B7IOvUdYSgCFCbPENxCqyGQA5F2gRNJNGu5pnJm
QbM+UCFiFuGor7HXOpUKbp8iq7onUq6BatHlvw2PhSm1syJ+ZNk6y2zCTiJK0vMgoqQEwNroe6g0
KXypO/0jln1U2cl94qZWMnu2z44Ty1EkAJTwBkheMNgd+p/JG6/I5mDf7WLWmcw6c7ZWmc/eESFe
uJzKMTytNGJvps1QZNBJFjdIXh2skQB0sT/rt9h2DpzG1TiODOF7kkX+UzBYofmP0n/9N9vvIlV3
m9E/STymxVuhzF+RWVf+EAQyusxzM8t1Lv71ZfCofMiCZqCudgrkqYScJz8ih8ubqnJ2fAcILSsN
kyeIPypTtYK2h1w3MZc/XWdesSASRXWVW/nGtWcARkU6sXPgpurPPtSyFuIdF/7+q8tLuZI8dWMY
J+nfEzBDQr2usZ4v3C59aMU8AFaFrWtsoQSgIY5eFP3Dc/reUbtsKpSbjjmfF4uODwE64DgEaimP
Rtzegs96X76RGkm7CsgSPJXXxR5HM9A/TBS46b+1IfxvdflMI1GCQrHrynsfYGfDYM86kteaL6Yj
HHxJiOPJ5+DM27LPT939O7ZRQQ1QPXg2WV9Dq/Lw9GMHbAFKZE1XZrepxzOAzDG6xJOJD2hNxMas
qJi5IzerXoTJ7PeCzmj4na77GF+heRMiEAOqQ+6df7/4KahmnfFnoqzgvkMX8v4EDW6E0nJM3Qiv
KhTupRZgDWl8tcIjB07e/0b9NHxTDXqFtqRM8iPmszGdqWSDVikYej6K2hyr4jPM7vAx6dFB8LWS
d4TO1BSQ38zu5kQMBQDnrOeSTjeBFnj8dEDwo0+P5cGDtDF6iRU3O+069GE50YYia6cER+rA+obu
tdXO9BBIWoQ7tIF0sLEq9EssMo7B13enizprJiin4cUBESfWkPYzjWucW+AHxQEholACQURlrF8S
5TM+/QFfzZZ+70qJcEwqyF9vQW6yX9ozpa8gFKH5qZ0kFqKeYBs+Be+DqRu9zxSrtRi6qW1wZ+Nv
6ejqSY+ko807aMsuU77pSzSNUOG4TRMUZ4ukClbtmj1xrktfpOZUhxV0vqGGIDOACsKTnDhBbMzh
LvOtR1yvtsvZSFC4rraN3qOJ/4vTLlGI/Rit71jbgdw9gbH0Ibe/Hr/ZbUerWA9BmC7ifCQHOvj9
D5zhxmCtPUPUdPy09mIuAMykAhxDR/xlNyZqaxRJ4ARPUf08u3DNHMDYa13eA4IqCGJq4I9csP44
YeeY3hUAhakc19uErVQyyD/rVQ94qaQIL+vTbWjROsvhRiBG2VpLq2xPjQ2E/tyqqebEaBKoTN1F
Mp6I1uQgKYEvuZ0i+douPS7HVfu7oPixPxyuIxeRw9DQLPWRp5SHJ2mxyKRaW8VviZC37UsQU+Ma
VSa3QWj1TIf2Y4yj01PFHrmKbkJaa3TVPp2DqVVtCB8PcZ4luXzdmuQVBUJ+8zp0K3ZfchqVPN7k
x9/gDvbD+oGkZ4hFjz1/x1IsdNT5tc3QycWgyC42YLzs9WuirEsxKIDbFISwTLPBBdLUGHmwEvGZ
er9WfNrUKpQ+NwygKenC7rd9ZMwE5jhujYhsStGTJv5G1TXnhDK/ITpDqqh906k0n8TysYdn105U
sWmN6SP4bUgktG0wIye8iHkHelVGfhFLOk5w0up5vqQluQDcTdDqG5mlQmislh+lmo9nSZpTBhBt
eTWSiA+QKpeqHAIEsVZ2YOOiV+NFm6q6YvuLtWNRa+ZD00pXjpWxp0lqCJWExraleDDr/N0j5wss
LEBh/ascE/P3wqqzLSnveQkqZXMkMt4Wd3j4zo6x4uhGNyNAc3jork3WVlfQvXxb6ZpVXTE9FZuC
2DcoOKVdZ2dwSLBUMVkGvAtsJVY9gljcy2uvIlQucOtH3lgFaj1QnvqqWsXLONOPCh0EeiFTPCVs
LpiKk9mLd3h6pQEfZIjz3CgfRxlUswCMvnmP5lokvI53A5unpGEH3GD0tuUZDJPihXxWBOSyQ2In
vCwciMZIs6B4W1lo0kGltaRHqqAClnYdavmCLE0w7CvNFG3CCy2OZKOM6UOO4vxyWB7W3vY1FTj1
aEiU6dEmTdmTiPT+YZ9RPC5RPnMX9zMmL8HbC9/GJiYCSjBFNOk6Zs/e3/LEiLwj390tjmWceF/m
Jnz7wNq6indtufXz2GNTKGV7jrPhkLy32gbgG+Jo2P0/hr0B5gamuUDFzJmx/Kk9LEm5x0/r6dax
3RhaxGBQmxZgyhabTP5PRseAn26H9ofS/sXATocznLO9Af5KIDnNedZ9whQm5P2qB95ICmBgDfDh
i/6ckU4Hozi4zRPoKt6eowqEKMczSVsVNIDxV7ctszoRi1KHI2hstmSZEHW4kQDe6dLfUROczAQc
ZFDmQzZbzkfE+2rVKPo1QPv+Jq6KY1gEJ6aGdLjCXLHhdMUEQ9ZGj3cLKiMxiaBc8TOUOTOKrIHm
VHn1dX08ELisPmzWfI7FfXPMeetxc+ULRvjAciWI16Jxe6Acmnjp5VDDKB2VMfAVyZfgeZm2n9Y0
XKJWonCRSo9azj5XyBT8aYrGRHMblD7YfqnHsDFNDfjEMgOmkirmTNA02Si3kqqqX1+N8TChmnzC
ob7Oi21sQC13rO5wJieF0X0bBmQ7sjpHtNU8ggnF++4jWIpSMdi3EC7tm2UctGCPkUcsij+jeSyf
LqFVVuryHFj5PqpyrXN641JKbRmheekZholnnb+2Lqb71bc6RGWG3T+Z/W7N8b9qVO2yOIWJTn78
peWEE1qztBI9cdUSEJW+juoxO/IiCqWNU35damKqxeJaGTG0Bir+p0bY7bdo8t9sDMRW/ik5gV04
2e9yyRCpdb4TgoNtgsLYL5+Ti8G8YBRGdUDItn2eb5150XGGBsuNNkVHi+gowGGRkgcT7kgtIQuP
qB/aZNXa9MvVTWOfrnp49grrXqesL/HAbVe+MjsUcEULthZx+kwTqCi7raOUxT79VBa47X9x0kAu
6wXSYSAAkRsJluGX3pTFyAsVAVlmckfb3oQdrnqOKeIoocTK5TlVFyoZsKxwU8yipkxopWb3GPlW
vvifNxQ412RV+5LwoUQx4xFD0A1YV+i6deYOSbBWfzDdfUKvlCOsT8RX8G2cZEa7Vpo99Pi908zS
W3GVrF+EFM9iMGV5NRYiQYaL2SwCdHpNP2rh2+xeAhTwId2IgiyoPQl5O3GnhB/2za3CGMG57B83
XwdTPk6YgHMtMaXtqCy2EoVQacyy854tGRT+4m6wMteS3Y3wrl/S5F3N0RQSR7FJOcxgrkgI3CXp
6eLvosaaWikKp5u86XBJvXKsgIX7Qo6du1UhAUAujryW8bEJtDhOB1o000nxh7zuckiKBfSGkkUd
0XP9wwgMMQIYdFJCRB5FRnGzFdlPqGc/51Jl2GPE1nOr+E+0Xsnap6uPORe+OBwq+OIuHCmY7hj6
JY3rTqlh7typA3PFCVVa9Bd4pWJEJvkyas5iO+r7HoG6tAoHk4GVii8gUUU/gQUgxBT1Zu6VavSZ
5Dk5hwoi8LpnHipgA4GIdmkHaZgXdm+C0pyhA6xqsWg/zOcFiLbDrX/frMztXOjt86MMJ9yR6I8/
DNzPwlJnOXAUb8MDuqUVF0VS9imNDfjZvWgHmErqQ2XGjBfNjtkzMYWK/Syr0iKOThmWufcT5ZCK
LoR6YOjS5J9u7vBC4VK/0AALQ0s6xvTcaWeD6uWWUkMLViHBkeNz7DJjqKkzKXQN092RZRlKXCgl
y41weLtZYAWJXRo4p2PeiXzewKQHb7BNADM9jvMpRsK2YQi6kdSp6c5lrJHIq2vQgndYgm1/EZ1g
Cwd6PNlrdkp1h+Fn6jntW2C31ma9zbcqHZBQVoUBP0+J34fXFxlCyfWBa0KZp/mTPO6t+CizjFU/
U7Kja16KieX7E2bf55YkyGqOEeH9DXYMS2lpAuG8IzXDFiLYbOfOYaK9GS/oxOXbo8GCjt5C04bg
v9J9WGNTpljQosJjYR2ZwA7ndQ42Xj6V2HDVaGGkEV0+B+YZuPVrq65hQWzpTV8IDaHiTwIK4xil
GCMblzC5uQVXqHS4y3CyBsAx9vBjvBLoPH0UBz0bWQmKdIAaIXOfiKPeNUtGrJnzt1akP/OJQ8Kv
BRiOnuYGxx7gZW2VGpn9kvdcU0zSyinXr23sWZdC+eC/wUSImDPixoGmZ94XuMpIDPNZfDBSWvgN
mEPhCd7WFMQ69U2A0uipoXfScCgOjQ3Q8w7b/oWzp6+M64LOp3seQEbHFbahKVekz1B1R9adH3PQ
uFWie19bPj/bCXq3Zz5pX5FGcqujqH+7CrOnBxgvIXxT2tQcYJbgyPy3feqRODBIbC3Dkv6D/Exb
/HkFBdr4cuYXo0eIhjnbU/qWnzv5+pyqHm+LII1gfcgnZ1KyBRZNV565G1OUD7MELh2M0eGtDqGz
gPmsG032GJlr8O7ykZ+d1/TcDNd/pGWHsQ42XF10yXuLZ5BJC1ZNxD7pcqnl6DBLmP8QtX5chdYe
gP7fkboDgG20AtNPyzjKJvqVZFqoE+HgYx86pm2zyKoVGcM3D44FAuj5nNkxAk+DDfija2+6T7PY
mIZtSXyuCs1Bq/6ENKaherO9rF9DrYrqvWpvZfYP+DKD2hzBbfBNUOOTrola3fdkirvfW7kS2ZLl
2jKAe8JUZA2RbvZd0r1gEZoyZXxxbK8vfj5Uqf7Txdckp/kqNSkDNL/z8A5IaghBsKvT9sb/F2Kq
RM/fRHBY7iwgVxK9rzm6thyfm4DDMrAMkTxRi/aX+vij14QH4clu8MoMYVWxPpxydXM4pQWlR33J
sAJGjMigyAxv1f/IuKBeFulrfXO/aUjAPfJkYtkHhj/EgxLFyTj3sN1I9Eok8c2yJDtD6ArLguGp
cjaEHySaZLxdR99NZ6YXkpD34oeaV12Xzv3FiTbcD9V1FQcKTNKZ0t9m2i6rbknXQfmF/e9IUOJm
bVUfhYmq4vUCx/ZCtbtxt+q1Znfxk7b7kLONoMTgeB5hSQSdnnd+gMJXDxrJbf+oCM5ySfsrxhXu
GZJHIS5cETHmr/Oz8E7q3LdWRGbcMFYDDoyluNDXS7RybCPdqPgEuj9R0C13yyk00mUQNIiJpt/1
vWzhhZ2eet9YYjIgeL3iPugTw27hNK5eE5wwCdQyzGjhkbLIXEXdHfeVTLkzZikamHLxvKF1WO1B
1kC+oMIz1y5tkCXSi3ahxYnAIiKYH3RtgwEJMA2onetjuFgxTFNix5wJOF48w4zX8Qq4+DaQQfKj
j9tSX2DeJDG5EZsbUbBS7IcwGQyGmokQ6ov9EtJ0cyTEw+HmaVJajU/6Fa/9+CPZzODVoxxUwJw8
DXsL3XhNXJFuynt7wEJh94k4dGB4zJmxJyX5raRBYjMvxMx0h77z6L3mscsmUrNsxylWYxJ8xgBd
e7IRnJW5m09YSYkkGcUY/a7r7tWY/mO+fwq0XGZmXVjGXOTLp7iWq4Lvh8yTuAJPCzy9eNDIGGAl
WxaDpKHu3hKtfhpoIeGDoMwFFAxQSXhi81daUOuNmLhivxrnXNeXf5XE1QQa+pHqdw9zWhXyVgM2
zYFr8QURpi8bwy7zjv8XZD1F/XxCuff/Ukx75Q11yaYL7gjtLBV+JNxCBOB0jgxWtz6XVHqxF/bg
/tnKECuSZXGBwZxe5zLUzla6V0FGw/wra7h/r7M9/JFXh5ZwJDnmULgxP2mHjrWs+G8Uf6hgYZME
t1NY+H+juyNdMAxI99JQNHR2rESbCp0ucXXRl29QqsWUH1t38v3yV2CnNHXBpz5/kMJm8FDowVDa
AdWvu3oI1lFkLlHDmtSwXB63tjCff1oB94/u9pJzEhNsnSltUu6SbPSc5Wg2UvebE1tTwmc8DCL8
0m+LkwPgoncFSQcNTFLnqTghrF3tPzRREKjjMex+XyQgsfBiOIEF0wjlO0hBQyxZxigmGivUxvR6
8kZrjkN+CJfXo+TPmUuY0JmS0MAT2TDmkloFDJibqA2B7JYOJPYJpiK2Bc2g9hOEBNwrgTiJjMPB
K6Kd1wShKwDKOn4RlFRMWHNMks4oqRAkEhiSn2QO1DoIP/1AJ4AAYcyOnR6T85b5axnv/W1qieNE
w02XFj/E3xEXu4te9E7w50R2XNGfhqd+wvcHG3W0ZoQR8yBiolWYA5kLUempQ9K5jut6uYcZHZ7i
gC/HQrz7Cm8NvAtoFqhGsPNBWNnD//JSq3pd+ewQJZ5fkJ1iiwH3ulWGmFycrV4A8bQRYoUNg5uK
7G7TdRHOTc2mycBBb2hcvDCvzUUQWzDksV1ilNE12jefi0SWV62AXxBUPtWebbx3RAc9/NEOgDfv
vPEOJHPemEGWwlgzuyWcNrbJhOB3uMGOeXiSoBciwZL/mTf3UcOxTbLjCFSA0Q5+12gNeQ7A8hRE
MQ2efv1M1jR1DreYViizc8o7OExrgVnGmdKSeMQaZMBbccn4yMszMV8nSfPgMJTUmahLofFhk56a
3KQFhccHoGO0KHgMgsg/DnOGdivdQnQUbfWv10srIeS9Sv++rbPpw+NQd3cVIYfaE2p8/jDciAB7
WyKDjbH06VDKeFiG3UzZhgT0pLtpVCPKVwlqkkO1CMjS1Hj0+141e3RqZTXwy+J9cprbWKGQVEOB
9G82Xj/hWw/arcHhsFHHY3+F6ao2IEmc5AMYKWFzV0/fPANep24aqvZBgr78Cp61qzFStQBSr6UJ
w2sjCl8+CvREHewSsuYG7wlpO3eQ663yQvdT4o92zJL9V7k3ZnZr/gfbYfEhb+mAgm+XXhuC7Xu+
ipOmpmJZ1sbm84TAlG8PViB1rWSrY/Cact2BoTSD8v0ZZzgbSN/KrHccvJwGVqc8fMvpdG1SJJin
YnFXZWXiBFBAcvdKbaCNI831ByPkwPX0zkfDcyOXu2iUr26bHIEWqL7LngidX8rHD2ZxjtYPfrC1
8FkF61637FPmIrWEeYBRNKFW+qYSdAZvCRTGbTUYliUywVHlFOwQo/URK+3Ow1PmVa2jFm1CqkMe
gFEDWe/BKIVy48OG4QHoFRjJ1Y7hmzZzoBRovxRoFbxWbipysjQOWjp0EY97cVu+TFzk6b+ox5GQ
0y5HdjflLFJVID4Lh6xwUouhS94JYaptWdxMyhhdt7KltMM72nuc2sFXwT5caLU4oF325MdnVMM+
7oHzhUlaNRuHmCPeY9qDlH92EjYl74H0K/CTFEj2gTmKDw0lgisrMrw6cf5rwJuBBo1tTbh9yHgB
xdDDPsrObQ1e1MEzdDok7o5f833ulHEL6gIDYpKNJctJvmoVNhmkmx5MJuCr1Q+47TKINAmmeMkJ
YmfAFLXNk/Ei8T0xpwW9Ui3QJEq8ThiDb/XM0cV0IueIOsaQWbHsxeHHJv4exMt1MQWNIuLsrgco
rHQ9oRa8T6SpRo3cOogWXiKActMXXKX0yhsEQ1ynEb5lRyqwiSbxYd7lHu2uvLmlG7Ro9LHctWHZ
j9sFEvpjda3iamqqJig2XGkfagqEIuUT5kX3yoqsIak9eoORla6Q9jFToxq7RrVrB50c5mraN6pc
tExGnkn6PDCchMB0WQIDFBuHAYMH7C6H9mtDJmKcChlHivCqmuO//QikI2u8v9G2/iJCycmtFDzk
Ln/s3nwQ9OSrwJY/UN+oZQFQ8Q94Voe+3y8gByjIGvlWkX8ZVlizk9EaE33/UMEXDmVJsYPjToW7
dBEx3y32I7BZKZipnnRIqrt3TTagxrkXIdPhNJxN5Hote6Jy252Hrah+k3R2hzmPhLspZM2InM2B
TfHy698KpqePJlzhP3BhxCwxiYKJvOyMZszzAPTXmeCBFlXy0//lCiaSgKXIDeBMOSyPs87zQEoM
4HIh0qtGLvJLG5Q+70qpmwQlzBa9B+FvIP7P2PVxNYFS+9lbv5s+fybBgzg8sKkCn2s1F+ynWb0h
FTwWVtzvSn56qYnKkXb2KP/ZUAUiOeyGLL+gQWFpqYQBFN19fXvdGZd+bApPXS0Prhu09Sf0Yusm
I9uzGbgsAgnTJvmrINpEPn0JdasVE4HOOti1QPFB9V8PtaQyjp/XHW3Be46Je+NJvt7vftW/9Yuh
wXHdvRbLipHeBsNVZrM9jrecSeuOVA64rrROm24n+3tVcvh+Kk3bF5aIAn4aWGWRZHjueosaF2y4
C8QUkdh/YSbxSDve+PzaA9vSj/xSRbuiZ04hHj0uY9/gzM0Dyw/A+qdW4dTOJe09QwacmcfJx4y4
Pxk40iOW5eBuHFWk4kXBQPsTwrc4Eh/oQV6TbU68VBwjsoRLiRl1KckkoSCnQ9RGTTPq9jmNI6vx
DfjIiU2aR+R8dgfcgBf7X3t8eWYbBUO7WVPpGkdICdWF6cJu8h/0GVwestLoFKzOC6tLMBCYnXtr
8OqgIUuSGz8LQpWe15GSmnXVIxOIyGXQyOwws5v0G0r3qDdQ/GnUmlOcXLRgJVrUpekVKL0+u+yW
dT+cPvZGMg0kVRBTFMw2kDOgNYVWb4KnJLBIqvxvmLIPIunABJOHFTwsswF43SED/FQyXnLSpxlE
V3IsJUURtWDmlRHToY3v/ckvssZtxuC5ZS5FGDLnuAeXYwHueLz07u6M29LJwPloE3/Tyj3q1p1G
Jji084HI0PMIYphoaGvxhiTJG+579tT9rsAgKHIb9MEWR0WkWzzog/V9J+wkI8FOh/dn4uFnG9pk
sJx1W3TpchUx+pS8DimjUGq1NtfKvqLQBsNRPT7hkqPOKupY0WtwVTxU2L0swLLUbDOXQvg9Km12
VBR5Z/LUS+9FRoqS4pTwtU3IgiOUtxtFLnOF1z0d8PcnUEm7nPzm9MwGWe1bkQ4lO+8Qz03BbwtG
/fFwa05mi4EPfOGalaK8pgJkh4ZCqRxc+QlNKOutYHJUjArxiQeh67ZJCZVqC+/YBlkIsBmy9jjx
zT5aM6T5kZyS7XokYGqK7Ef4uGN7DX3wUXLMZQITFQSI8vV7yBEBYYiM11pjee/rx8pgEDXdshgT
ZIVfiDXZQvx6Oler9MFY0HNZjI4LS81kARcT6E+dYOg/Dh8+ty7eviWP2+fSoVca94Hlu6oLphpp
KIs7AnrgZlSnpqYAbY/QpzqtlCRyFkU5592v5m32BYo77XkNL0S/1kqxp2DvD4yTyM5OjHBrqy39
wxgbQykYsQ8knCOUI/4bQpTMbPsQOkqDxzog85//9Ka2cEDWCWSqHR14tqg64+gbTJyCU37YxZEa
9+EX+uEgG37ae9e/h7dDMVkB7/UhMtLazHPjjIgAMoY6f0DYJom+mxroUOlxDYydnoYqpZII8u0J
7lcwgVtAiZct5spwGtcorD9Zxu0WlKPJRdThXprqefksoKx3wP0rWVHfpvXzPH7bz6d6//D9UcH0
GoHI0KD+5b4Tkc2IV6NAXlcsgFsXouoOoDzjAtxPeEQE+7blbjJWZc8y/z3EKF/q4PzxTp+u7Qau
9Xta3lvfPMDCoyii7FCdevuWB0eQMRcDikKRJRppgUMZ91wRyNXtiDCkmf95DO36DSVtHCW1qbPW
Ej8KB8xvkJyeYgesOtwq1JVrI6+lVutRMFQBiRjCIzSRNWDTmoJd4iQO66b14YShrZVS36Z8RMzk
1cJbbXJR5J7cuocPy7mXbpi1e/8grzBNbXOpVCEFhbwOOHvN2MkvOBLcuhzF0Ngerf6i5zF1TuIb
zt96ym5CtfsJVTwZwtxAGDtR3E6MeiwrKZYkly/sfEAXf5qXeMNLQWQtX7vfMr4GT3j3g+ASw4Mt
Lfq8ay0b2R0xFLM/MatfXPA6aBJkXyAYY/VKMPN+Uxk9F1oR6p/7Rm8zTd0VXZaNN3MTCf2WHEu4
fF0uulI7UCdq2BxurQm7nP+42zdnXsB5PQXyv+4Ph8EtNLSA5Z1MvuwicgW3S0INq5tPhw7olCbD
oqbBtgr6exHD5ej+Ai8B+e36vTl1kIvtO16FGGXhfJCA0q00nyv4mq0niFwPkaswZ/eTxIo7rkJA
zMr7xIfq/8qid0o9G70osFIFhTwQxtrpals4xzXbNMKLHG5pVs7BEO23bdzPx585qtJksIAUMkbS
n3oCYpwOwz3qvfF8LY/37coCDBXplTdj911htVbRsY+j9BAmKJvs0sOOKJZVavi0ms1aiYztup0d
dtHPbg5Yj+fPJILoYx4yBln24EFigdNZzSjlTDI/HyT5PkzphOloO3yq2oqu06VWXlkhvh44ZN0o
I2uljJYy21QftR67BAdg1YVXxs7Qo8y23zILddqvGm/GXTOZrYfQKGSLZu0vYCUuLWzBwVFxXLgL
wQP7p34XWfIBFGgbEVIwf2HT9FCxHYrooGMaDq1GWIhBpnrSGI+9/qXA/knOskCM89Pax5qmb3KP
FuCiX0axoI1Caas6EF/kiSIW1nSOlj59ESh7+eMlv3cftuzlem1BtYILK21MSbsIVeSkhCiewrhX
Ua9BVUGP9ZISzXdjOd8CvZmq0Y+LYQTY3OWOI8q8RHFN4jM+SHqcwX9+7Oc7pN2EUFRt86VRpqhV
M7yQLY2CHfW/uq+NQUeMEidErqZZaB/ZfDA1eydswDd2MyPk13NA9or3GnTargENV372R1Nc/D3E
8zs1PcmBobuTwbtk/sxB4VMT6cwSnjABxZ00zmVcoqs2ESmSmOSgWP7bngvhzyD/amLL2y1aCrYj
2uFz1X7/zSqVFUU1VHGoQ2STeZ2aUhlBNtFM5A9DzQUsyFBwvrZ/IGJMIpVGNr/tsrNfsVkQkq7M
akqJmvdSwCjR7+PVLeyuha2nBqiNhv891RIsprwp3PjtD2vZvX2wxBuuPkd3+BASJftNp3ELkM4f
Q/RnHEVE40edSyO7QObONYos6A2k9pF7FMA3yjvKpjzVemXYpyF9sN08VRBsnaWjRatw/yOaXQMD
LUOoIHJlXDs5b78S5ZT5VFZwLbTbhyWap4KBHr55ypFVjIFNy4m3JBSRMshBw3ufRsggC01SkPqG
g3M3ySBa4fcKZoYE6oNOmXefZZN/gMgQxlN5IEp7jAhVnbVjnLWpiPi1zToEE7/NJvRNP73ve/bZ
sdDGfz8D03qXusmJfsCDTjetdC+BffX4TxUN4cDEJ7dCbOoDqL4r8mx+pnDM8MJhIumXIxTvWyRo
Zje1dglwtjVjywtaSP6A/BFUt9YXmbCz4UGKevvE71DFT6HsRJgkVZtEzQNz/ijvaMEckTm8rg4C
61yJn3rQNpXH/m4EHlddGTaxf4FHKiGb7HF0GLwmZpYt9DmQe25UQX64CiPj3vzW0j037ESeCzRL
0BD/h9yI78S8RswHiZ3AliDhzHCUSL2KzyQWlVPkVczwVY1kV4qqH8K/0RlJxkzbOC/3OAzBdQzC
l328mthBMqy+MrKNTd2yWQRzWy3o+awhvlBlMf1sV6sD0ZEBZeoDz2kxgOrR0AD6fdQNepshlnnY
wAc49zFh5G7AcCY5ENwAkNgjShQRGHbgbUL0zXsq7KRCjdBWFpNqi+KL/66WjcR0SIqq+cfo9ddV
kjyGUs4HzycCSaSLG63XpS1heP495cuH6aY88/Tm+GgYGFT5WWf1Ugyhiz8bN9vMoHuR2k0wqma4
/boIpcB1anbYm9GvrKxcq6RiWmWjJqfq2tqt+ZVQWa/5unfeg+DCghERydPXgDeuLVG2h5/fxCiu
xWdfRu6EzJ61UuRmwoLPPmkIx3ticpF5xWyYJP1rh5g27KoyScjOyz4Ha+I38utiCGtT3G0CNfod
Nbge2ah6OMJuyjbvuF9OafxgknvfpoLmNWpHUUJIYDs6Tok5EF3UN9tSkCMfMztXhCTDLOHKEJpZ
0ZAZRABuZH5tt5yrofrq9Q+Ct1uh0R9gXEii7Ftdl1hGtDUjh4aPHutfgjj2g6xceYr0D2w1nOlN
21yoc1tWjkZwxtTy033UOVfQoRUmjbD+gPd259fG/eV8uZg2a+Fv4DhCqG3kW+A7sQiLxtpYuUcH
61sPs8XdKbmVbKbmylHPi9SgkymBt1MmxcofjHExd4lhtNc+//QPXs0LZ/LlNMQRjjrUWOYFp/0V
mJVim9JLGoIu+iLtxJnB8UWFAcc3SS3V03cdWjCw4XtuZTWI+qy+MJkCwYULQrsGxI9iS9k2DZDV
P9Wi1qpq2KcW/qMkmgH6rZYYRp3CkQIEvtzc/mOmMl7mkVZp29nM+VgLrsZrIu2nrLzxfRgn/9fz
JnwTfOCergR9bwdv0ed7GacleHCNhg1yOAIbPL+G8+EVlKfPgr1U8lncxAM/qPq7loVnL8Zbzae7
mA+Utbpphs8AM68fL8MKFBMl6pBVWMiowIl1vnLF05fzi6HfuPXZnRp8EOozBWxRwhp33n9WE4l1
DDq5z+a4hDBapgA9p+6d+j+jsqqLVIOSHUFEvslNmArRPlFuRy9n7SulEESkVNsKVK4nIElig4Uh
bJt98giH9kSlM6mlJ4mQ6iEyTA2B1y1M+tjgC98H9geiBgxRSyQRA4GldZdqvgFzBfzCBQaojhWJ
CR9+Vc6Juz2n3oF3C72hufP7tIhQlXW0dnFVHAytb7W1mLksan0FiiOxYopI45oU7pmtGLG2JJip
fqPE7vKjInU9sobhxhkbzMDZC9uj0EyTOL9tMoQran2hpUYdCVqTUwQUZDKwHulfTEAZRiIvSlei
fITsZ0Y+Hx6m4Op0Ocgg8KtY9D8ZfOq5KPKxPd6BiOILCS1dJMPlr9T5WwjvhXUueTSVxCKwXJa0
Rz4+Ca+yl9QTZjKE33D3IRwasAKkd+RBNzTRsVeru4o99AErDT9Vtn7PUM+6dal5zTQIuOYdVR+u
NUkB4ZgFkwNCIeKfHDv97lYwhTTIa60uPC6z8YPGMu1WnAgwYM5O0PQf1p8s4KMgwoNILWpw2oCY
wcfU+tXuQw52d2QQHkvuYo1nPj8EC9z38lwyaJxSbUHx4ntzy3PayJfltKD2p0pnH4udPr6r+WSn
/9TfnG9XhMfzd4KBFIyMpYX98tJNiO+BEW74dDpblP22X7HCXxPbZscynsObJLN+nuJ7sdG6lt4U
ygyTATF4xoRtlz5nf/nyRRAmI+59OkmWkwXddhY8grO80rE5PdnZMhCrfIc6tl5GQtJUwOQEmp7q
rUhsund8nz/bsy1X0SynnyXOpTz+PjoCXcFDb49cwQlkXCXAiPGA9RD/kZtqjBFwEiWmMc2jj/W8
0Rz+fAushHZHo9+IkLvEgYgFSc7NNO53Yq9ZzaqaRx1cWQcdGChKSQbK4Yj9Ipl47UHDirr4HttP
8/3UENQ0nJQwBgDn41LEvinvQztoKuAgfKOIiLpVaxXJ7vDI6NDzzmlWIkNH2ei6oJ3+ouNEqcov
tJM5nUlFC2syyxciNNT7+nsAVdf0vs3iERXW8CYz8Fy9qoYWbUzaTh/KCqPCWotAJagRmi83uzeN
jL2pWMVB8jHQJU5k5nsqShaU8t2xr/t2eUGqfWYqPv6ncy71/utu8QFP3bqBrz7rh+vIGqNS7PQ7
EE2R8k+Y7K3H1i9gX4iK2ajFKRqGFp7PG6XIF52WE7zACwPYrC8ocxC6Y/i5pD9zghS2elAvX6FJ
xD0CvhsIYHqYyry3BdVJyVb4hcYbTaXZSngDnKhlxxRSo+aoqUSx8nD8VwvgiBaFXTCoJEauQ+n7
a9BpCntThjikDu0C6W9JLjxwrRjlRrO99g+zeEk1POmG/R+UAStQWpLbYGBlkJ30N/8fQhS/Jdv8
ZL3VRywjcEdCsmAri4fac/a+zcwd5+z6GqMeD20UFuorEFpiEUnbCpd79X85NBrE/JPWHH6Z8Ly+
dV1ERR77kXYcXMGYjp1peJqK9SDM0r/A9IEY50t3bcSSuoGP0dc3fe6vrd4zHMtan3OGk+Tsa56d
epEAhiZ1XAU9bOwQE0OZxh0PXzFU4M2t34EYXbh1M9I3tiW2EidyS410VQfp+5pgf+HI3DqbiRvK
eT7d6GfFY1a7r39YS6tWQeWkB1ZZ+9q8hVsAVTnRofh5ya4jtJ6IYjHJG+a36546QM0Yb8r7gAOr
5U2nthK6HdNZhnhCcJUpKB/m1uzi5htloRoOGeQzai03vnA/vPCuxTwuoW4kIgdhpVgHCtQT2jQW
kfVTAInE+Y/kSr774CMENGOT8FxXEeDDUOv4xM0ybBw7gfLC4cZf7Is1t3tl4hvL0d4xG1Hg9+Wz
vVKM2TGais3V9nhjbcHif61gWkyyJmzYOhyjkPXG5p16BZSUJejsE9G9f6eoCxVStSvzDVUVAKVZ
10T5+5Lkohyi00eF4gaTDY3eFRF6yRZmjrwUBYNiDWwjWLdXLeJxeFqf1z9UFM32ftfiMKdOYHtw
bng02KBg53rE0zpKpayJS6FCKwEZFocoa+1HIPePlVHlA/n5ytSWfBHRUovSERj3sFNZDvIVvV0I
u/qIwMmrFzVrR3rp1fmjwkIAP/NvnnnuQYmnYqkf5LVk70+1b1wvoOTSUxMOj9Z2ZC51pz9EKjzS
yS2eEs4TRkLSwcuJk6nGWXDQCqWnR+8CnmEbPFaL4+ejPGGPGf7SIy67YtxHycOApSbbE0PPdnQB
Ta87yCP9vRVfF6DJu0DpPZtzc9i+SUwYZhDphI41ewvN09nSs5MvHNax1ETeOsiks2NZgezGOwCa
xBfYCF3EIwJ9PGA5LcgtNjm0l570jsW540Hxt2m+ZxtG63MwGuuDfe99mM3AdKrXqE+9vxOQc9Wa
DY4ISYzXXSWj4dafkMOQ7wDEdGITUKNPuQhpu3pwJPKYiYHg0nOZILWggmUvFKzSR4DC/FEyp3I9
L7++QFVAL/p0z8wCvirjd3QdE2m1Z84NezSeJLTWBvZffG9FrAesppGHjCbgE3wyHRgfzr7w9UWG
D0d+31ZeYOO+LQq3FEeKVBq8dB4MNQQd8OWpLZRlcaUdl+CS3T2Zhnlhn2KfuuuJasguefNwA+jk
0aDmbxkK3za8qc9mtQzETlSgZSmw22QLPxBBM8NFVLERYVjiaOq/s4N7sKhYDM70ckLI4VpepSce
3WkzCDeojs0Ifg6jWHXb4V3sqE6acCjeAsRw6XibEz/NUS/GBZoW1/+n0/G+tdFotdWjXSm0uo9E
kapN8ID0msiqFK8OoZa/oWDGY1Oz48W8kpI8yi0RLODr0IndP2lQA8zZXJBfSa349aS55J1JxGDe
hgr5V1cJQsfV+0g3O/u/dmfg/F92115iIKFmxNHe3SmN3PCl7Lvz/+VKOCYc0DiiwWgnUMDjkQ3C
UQ9+yFzFxIkpvxhwKwV2StHqF3qWMhzfi8MU3goaQPfGKhhwU+uz9ot0ORtT1dP6nU6j/ZRZJmKo
YsCIciW8sCtDtQSl6+WiRTJxd5Sx6wqCpzvT4dWBB7UxiiUk8QmawesRXGMvD15pEDMJ4X4MiCLS
NudRXBc1P9Zro1doTPdJokoyDHiwAUFadV7OlwHuYEtMDkVYvoOJ/j5wxDKS+P3rgbvgT9Ewfjwo
IVbatbjfkioTcuCTl4xY8KNxs1XWdY/qazc5QskNmcCXl9rR+ssj3wOfkAumcp3DVI1NAXnimG1k
uZuAzKOdz9AKekd8bsZH6+TRa4inecV4w/2O4XkbeDT7VDMv4HV4RoPZSr8MNSDbnr6pgtSnLxaH
EVAoAqgHMXE/saJhSwcCHITsQ8O43l+kw6ugr6cJEb0WA2zw33WmS4tr5qPQqr5hyr9qPrvlZccQ
t1V1qkdYtsSYfeUTCf3r8kpbcmfiWjaqkzKGHk8sSHhrP57E7ZcgkGZO/ZDJmY5ADXGBOvWLBSRa
cSXHieKQDHflAso0oYFQ1GiQYs/XeZWqy3peRURUMPmh0wQp8u//SkZsyLrDWUPM+2L6MQJ6h7sZ
IGH85H300lCnc4AEFMVgmciiRYqQ5Zff8L+w8oH+/1jfyF+qOZiXLcDPQ+Q0OfoM9uhQZVubFrRw
SAErMWQI50UdAoVUZ032XonR4ANLVGe6JzzZE0X0WARQEK8yMDnH1cfGFx/a4b0YnnGgVnPPl1q+
RNV2YG8Vz5tkpr27fsK41XzHMzlflCBaQ0es9SIpiq2sYg3rzOb5S8Ps6viivqkMgnhuth8xVdWS
cbguDD/ix1AgDNFztNL2M9/PzLzKHX2z62I+aRVFVKb8vN2ipGjlcG8PmPtmgN6GrIevS8HDG6xw
XYw6534sN5hG/RBRDn4KDtX1FGuulHcPnpVONZa1HMDk1+ZJdRMC26nWOJ+zOdp+vTYmEjju/ESc
Q5X3qDpMkG1aVBpf7pDJy3KXi3GpF5KtB2RetuQ6t1u1RCBDTVeyCvlvKTqAnfYZ2aMTBoX49S++
cVMwQzIFJLMBOo+tuu44jGJgUMYyyEgTF7x8lj+bml/3AXVKrEgiO3E60X53aZMvKn7IulrfaWz2
iaQ45xjaqVTKReQ0B8RLUyksPzWPJJ1xCchU8T1c8OldC31TzvCpuGILzx6+eozUHylqpHJo3WVX
/xMiapVxSkoML+R3S+0GU2G7Ky67PO20vpOZ4WUh9mexCbICBsfyEyzWChWYrHELH20EQtCZqxZf
bB6lvGUyXOpUt2GRKrpEkEIgXSfT6fOBTuYTZufxfn/ssJ1aDw2HfrJWQVL36S/5owmj1rsfPdHz
Rss40OuyNuZtx54PdoFnXqX98yYwmLmXK79iublTz5HybZDm6khL7BgVKAm8hP+Lr78EhdF4CmMb
PzVfNDID1FI1f4vSY36JlETJ+8XKXrnhjpgUQ0Q6HP7VuazvGP+Yd9tK5Wsn15+hlybQCLfMhMbB
KB8ndRMHNaYSQxSMisA8qccpKYBQkZqQ+TUGW+Oq6zPbSGHw18cpMiCM/KRmkHGiiAmZgB4OX6C7
WBiHpIQIhRES3D9fZ0M16ZKQeCPYo+sDIVN0Bz6tIThmjZ/MHT1kctqVUSqbswJSC9B3ca9lkNlm
2+Xu0BltMCKZRCJk/sqP5M6qC01T2YVCb8Z34VUEUSumjtsdfMtRpp0jdZ7EwFqxTeH+TPHScRcf
duMYbJI2VOPTUlVgiXgJR9KjglDP6x4lETWBKmYy7bv3mfuWptmqMi6NfSrreBpuSm9pvUBqI6II
J2V8dQXIqYCWJcWqKGWFKUtVaq6hmhIx63z7p17asb2NiIwUKS4IEE8yigmimngaVogS6uoDTLBj
ZFKQ/6ZgEu5n0XtXEAvidF9rSonRyvqel0NK7ne8nn9Wbos4apnuHtYEidQxdIlU0OKMI184d7e4
2u35CBIwNRfnbLJLr0I0hJdJjXf92OsBoqwByaI6Ny+mH5cmvgNByvOHvvkqdYtUsyqx+8NdgLIz
iN0lwlmQuEE01k4hexn9DUT3C0rkvuNHFk5G6Sbu467dP1KMKCP6jmz0a2zoLpIm4cq3YnCvvO+r
9UI1izY95PxndjOLh47kUQKOSgTd5PNx+RD0D2bFsAAhOFaAnI7HeD88t2tUw2C8Xk6cK/g6Q6ZY
fo9G6voitItLH8HlaLJfWZstTDAjgF+OkLR68hf/jh1KS5aV5/DSygx5BjpyX/Lv0EImNkcyI5ah
JqnRscLYiCnJndjyGhcJF3Z2ftRrQTvPPwCTHGVq4AWKtMMYjQ/2u+5840FPhHAaK9wSgLdvavN4
WW110l4nZnYYFs/q6sq5KNeb62wylcSQfCPXWa79Nt4WJjhqIvUXgK31KAj/7FLU+v169+89eNuN
U50hCFN513AJ9A3Vx6hmc4VuwHpiTIBmSYDQ20YdVAwvf7RaFyPJLLk66tJxWan1RqThztkF6sPk
SlmckbTDguJtqJOl1XZp7XHwmK8BFs5y6IPRpZcc910mBrs+b32LLpLpLwCZ9wQMRrgTw0NNMm5e
1aefgYRqqqOuf6BI2v5gJ7U/NfjNYwn0vQUODcGcVi8IiiTZnzb1IAPhrtAliZ/CxK9P/W1tDOcR
bSTTPr/cKHdgr3IGv1AixzvFIrbwX5HKEKARA9M5rDrqmJwZtPDCobIj05iKzi75O1Ni8aBftf8I
eUkJo5IvBGs2OKcV/Uti3MFE4YvCEBnkKXd6TMxqnI91i53H7ZGcONSIChyM8RUeJQCQmudLYeXF
eWpMBB+H7LG4Ykz4gNKcuNW5ZuBQwPvf/x7wc9wyhBgfT59RYUw7N9eXjrtn8xRgyftQz4C+9iAn
4IqdNmVeZMZ//I/oZ5zkSDwm+ngU0Vjlshuy8PbhzeKdPyLYffwtnXq1MCxFr24TJjd3spMoGQSO
pJ3OocgDG1NU420rw6iqL7hqzvtAgJlGzFlItcq4DNTz/1J/DktpXWF+K3BQF0412pEEH/Qt+U6X
ZZS74nyBv8mzod7tUZRDNwtXJTraNLqo5nG8/Ettu7HkeuiNxaiGQeeR+7L3hS5kYtxwBjO64Z39
mjAzoTV/FPfc/3qE8p3Ttf3E1tyjj6nl6igeJMLTuIe5PTmSefblcl5QNGuE3WrX6B588FHGxJBV
JpjqAtCMweEUlRaiIhvhhWhJ3bCslsne/5sa6BktMeDQQ81l+NO1mAOjp1fKsmDIf0zWumm32Y/4
k7LkHKzaOVeyIj5/Yg/IBeg27Iid/t+vPfNkILftlVQ53RYjdtuGN8oGVMjXc0dRxqBOls9I+g4b
l1DOj01bwTKPEMJEzZ66tDcF7tgi61mC035T0R5Coxd6KHWmCuAlvh8ogNxZ2+EGVrlsllnTtdw9
9ecUWOX/twQyk+IyTKLHTN+yJf0Hxd7qSjPRNZARDqIyFXrO0g89R74qzRpN1K25qh/Ddhx8snT6
35xpFEXt93MUol1oZP1dH4coDpQVuFOkHNdFGw/95WQLgKBYR28rOyuqwaqb/aMwNgZapV+Li4sl
WqTum/fmKpMrcX55Lton+gzGwMzyTgjluobMyHakaWkH4qor/2RQgByY0iZHxlofwOlP22E2r0q7
W9Xo8fgYXymKN1xR8Jr+S8KFe5zBUh3911Bk8JvgfTHC85sUcYIYKB3cQZws9FrJ/OggnJIi8gh8
U65KtrMJlAiWdW1F1JoDdFREPNPWdsQPujcSzSuC9psPue3N/iUQtDFf21n5gGVvJ5vQ0F121WdT
4tr1sM8Ic0jNxUWyzaFF4SaGLSIYUHwyvFAujydvlwIEDAuoNuysisSPgiQ+XuqDSlA64F8U8LoY
EQrxtljUmKTKqOo/PTVgMvhCpfkRo8MknKoteJikGtkxotC6/Q/c9Mll0/9IM0VHLC+5BOadkRzW
M7xb1e/kHm3HuEZ9H1YjT9lbsKaG+q7xxy8XeENnmkDIQWWHvCyYzBrjN/wY+bF971I/QdQ4S5k0
a0ujWRlG2JfwLSFV7rOPAOJPw4mIJ0a8ccPN9tPTlUGB26Fw+0jv3dzciZXHk/WRLvAAPeJhyU6N
ZSZORJOj3tp7QPZHcJ98F2BUV3E9n7qZFzJHTq2N+Xa9cmKdU0JkolZ95zXsgB/VuQZcfagfYHT9
Es26KCuxMuxDOk+Wh8kI1u5vOfgzouWevtP+AC5ZPMykfbxjeMma6n2z1fV0X9bI9cPDxRhE6O4+
R1C3mU2QwgCV8x2SC42YoEVLZNkUrQGNji/rq3EfQpWP34N4702fUFA4cOLjhU6a1qcgL3vCO0Zs
sZTRHgNMatXO5xOAMNWqlFCTtWcqDCtcUqGLof5AwD6nn7QfyQLJa4cVKNi/GStof4S4E9OsnxfY
5f5RlvFTV/Ze6Yo5+5nYPxfBKGeg8zm5M6G6z4pccIVuAjZsJTaEWWyFLjPRsArKRjzJGckoWxyW
2oU6mN5PC7C3s6jzt9IUHT1bN9RID+p97MJXUunHXTHOQxL7U16Dmrek3B8M0e5BQr6Mw6uKHzha
aim1IBUNkwGCQ9j2NiVpt85jijwU2KUBBv85aSM3OOicsERcZaWh1fRlho7nb5r1uf4B14MBxstc
IKRZioJFTc7q7f8sz4Dfpd7rEXENvG5xW3mwkUwWbzJNS2iz4OzGeBCMmatky+OYTu6N1fqp6sHy
Cf647FnvyCI+SaoD+FYfUijJmbuafAJb1cImKhuuwGo+USaVSY2O+cqIMESDfEmGRII3qgv91+I+
XbEPiwqvfQq7yI9swHc69ydFwjvk6dfRsSK61Odft2oaPQ/ks04R14Ildiv+5WAooxZl/Vy+LRt7
/NrKvGEttvSrSF1IomRUsUZ3FW7sjaZAlOoujx4J/+EFDgDX0UStLHIYfFKKdZUyGrPIcJ8fKN8V
eoaGefLRfFBFiiKB8yb1ZiRL8YCQXz3uZTEct9sS0kMMaqOn7wfHDbSmktJ0WaXJxvYCyu2gojX8
sYi254zEhedd6mRHRpZmLv33sapWpU0pX55NazyDoHo2xVFQ1vpOkCg54sqWjmOt8xddCoGi1cDZ
Ezut62WRYNthPB9HC6v4+/W3Ya27TnE9iJIfvUckIDy47pqWnD1TZFuORUrCDMOCXY1jf8tHRI1O
rU0uQEU1vHmHywtthjZi/HSAvOspC+glb9DmCHi/R/q07jOol6LEli44HQwa+dqci7boGWqO/2xz
GUbAGhti3J9ypU8vGHKmE5iOsaz2+jDy9Io4ltWVu8OTBCFtBbbF28xQ5+Pw6jzqY2/afPdI+ICP
ueSnehiD30uVwFL0AkNheQqlxxZ4cyEq6mIWaigZlWutHk5ud+JuH2R6FngCfxwJ37wfQYNN+kFM
wrEmDdY2mI5tD22FyH9Lo5oA1pSaydf66xCtmWv1dLjHHHNDJ8M7uOzbrf3Eq/3MTru5PHmg4wLK
9D5DyFexLT8qy1mBSWvRJoDruWmuHMr5X2aJu2g7O/q+Tw1Xm1pz4DyS/CTta1frAvpJo63ZoBSp
B8QoGx16Hpw/lkA25Ui3ZsaNmH5ahr29EIbSG1gcd5NcWbq+WUxlFWPvtP1SxSAp/zfYc4eKyzjM
tMZpDT5Y4GafLc8xIZjTQkXqjSrFnVcMcye9RHZakMP5gOR7FqgxNV5L3pP/TO8pFx4X7ayqgBX0
BaLX1OnYdJVdnzz2L7aSSA0r9bK4EjzF0KsfXalp2qaaqRysgRWBVp64dreSOhDcdQC6rzuTVt+b
dNNj/kqA42uAu5CzgrXhnlGUEs6+o7ZYuPJ2n1peTC2/n2x6mZ+qAOZVqTHmV11H212eh1TZhHh4
IsufmZBovW37RGemHF13mrmqyhIj/jLb8T6FSfv0c61u/3cOmhfnLKhVywsm6hSWP/QCnR4vOIIf
NKUKlktnwFDyJfwyTcLmfHzc+i+lscZ7dIf7Y+OL7zv6TC6V83iluHbResT1pVdtIReswaiO2E2I
1/I0+6h5zscMFrISTaG3unJ5MB78IDItdvotySUECyCcNHAx4VU7NOpR24Z2eYbOHszGYAUrvqvU
pJCWmjTuS3emrpiVFJSPt29Jso6aU8oRqo3Mpbgni+sYjv4QTDYitm1EIDhD4MEkWdKCdsv0lqTC
o0PucAmlUT1G+UJdvA/sZG6/jVmY+A6iQagENKoM8HXRbmqJE/eRtFiLn/8UiVEWuB8FyPeJLAsI
l53UW+jEEid56VxYdxutK2JTTq1TxTGzR37wnZVh0yREp88YwuPBYeb8gA72OpBqGxqxbz5rR5py
5v55saLe3UZHpCziu1AGJljCoMKOJBc12q+IEp8hx9WCJ0P70E0yVDQM5FeWYqjV9BxRf85FnS9Y
fgwM+TQyR7lfGc8k3nL5FQX1FolCbxoKuGFgEDNvylV7wqVLgyIvkxqow9S/5QesxuroJDlKlBKN
i8Aqq+eb4kKeLzMHqlyUjGcDk7TLu8vxDOKQsGeO8f3A0rhGEvl5EwE5aA0QOquCb7lLX+rFUz2U
mOwYL2SS7BCanVw5xT1KMOnJvOKO5WuzzJQqao885ISeNOafAfymqADHaXwbP/ZPeM+bzlPyNa8W
KPyln5GLSFB41rmdyrK9JaWgWgsNMbV76JfP2O4W7um3Ks/HDMzgawce8qniMnCj8gQYWUCCUifZ
5K6epyhfM6TILJtSXnapmkxilayrmWqvi8UtDvkM/XyILFnmeHdbT43kS+ADhw0c6RAmKTMolgYB
IqgUUOkaOvFSmQC3LP9EnNY24s0GxxzJgmj9jVogjqogUe73XzS+GdRGatOcwBOui6WJYw0nLCXn
i/r0BhJrHkX/astN8hvH7YY2N7/7AMklpPa7/3R3bmCfOCoyuAjzZEcsPSLzQRW3tzHTDwgmt+50
+EYzWJBZLCV9sxgQwHbOEcKmZj6U1aOxXd3ncavDKTfLJZHVSL/gRTxzIb2JguDaQ+p5o68lFPRo
IpzmlpYF5EiC4PPPBITeXIHuirR1QxufQzIUH8cz0MBycq/oX7J62x/E4yZ3S/1/q9517ETAMhG8
CSrnnAZ+Yajyw86FoRzeva0O1/S+AGJMLI7nUGM9KlJXFbfI7pFyLJanXNlbUx1GBqPNBgM6n1/U
DOrd/2xVE8B/hBsvqBxlSB7kp228NDIvxY+YJqieAoxFc6gBf1SX4beNHy9U9eX9WbJ6dGG1BgK5
w6tzsOFp5yg6eFFS2Ziy6xopJJuKpORT+ZIkyF+ftyUTtGtXnbbGtoaVd60cko9+gV7f3pR07OKF
xeI9CC4d1bY9647QyxfclPwRdqKPLK+FDqEEas3qmJC/Z9m66k9e7M1MI5b+XAkC4uejuvTAcLfo
hcAiBLYNrpw33mZnj3+xf42xxNqThdXYgAwkNbIeQuK/te/v2APuC2LFXs+24+z4XREXyLXRNKDi
OKP8VpQoP6IQqYBFnLmGpYwuDCB8OJkzE45j/zbgHVmD9a3ko/amzQ6tVsseuCP6qMwkP7MB3c4c
X8rnflBvdZ3DptdON77u6Y2MGt9qUnTvJEnG2vJSW0e/5RvgFiqpGXberYPP/Sb/rHKLKIqCGYCD
m1ap+Xel/yU///WSUxN0n/I+j5Xs9T+g54RuFTrKlo6o071MDEbGZt8gfyqgbtAwyHvGgaVWvzEp
LPfWsQ+n3eDkCyS3bzAIotsb6J2GSoha9cYTDqo8Ojtrvb2GcUjdR2a6eWAH9vnxVx9sT69mQVR6
sp6qMkEeia9XC5SyXiTbGs7y/H6fV8Bggq7iV0qsyJARi4iJ8JifgpvYbRP0wqdLajzzFpQyRYR6
DFlq57LORjfdK2ES9Br7jBnsyjmJhZin1+9Aph7+u4JSYet2UdAUFuSwYed/GIfiSZFKzK2NPcr6
GLWx/rAOfO0MRNSSO3VmqGUMK6QDa2qPUa8oLrf7c88iVFf08aE33op5nQXmgCoZTNlmUF0uIcoq
9WwzUmiE8bVvGiFNN9m8lUxjjB0g3VNDGsjeq16fTiNi55UfZtkpfSOEPH2c0618ClZD/QC29Bub
Gf9ucrWi7SpYNqr46mxC26sq4H37cmEtLKC4e7GyCtCAkMc23FxfxH6c9UNvwXr/74mOfdfdbTA+
yDL5x8CtiJEjmBT1N6VdBcNgXwL+zynb2/lvzIZhMmuy7NkY+7cWlLATvw0+seXPhB1bf3LmZ3uY
FO309jiwmlYlQ79Gg2uPBpcdez85zwP4fCP0gZ3S5f3WtMeQ2WjQ5GvN4R9fi0MsLRXTiFERdLlA
Lk7RSzjfCtjrJDADKCCO+ewdzGF/GXEPuKWW2kHDggiekHgwCzw9ojwRRGJHTQ6lsEAV2ny279Ct
UNPKcz0P9dPcg1JH6A0HD/SF62C70xovnubGJe62VTqmBE8Im+8qpdujMGEk/TC2pfdpanN5TaJs
jY/9tu1dZbq74tsEmPHi/H6FDZp28E+PjCKfEjaWfeDNEfN65Uv5nbIHwPbjEECOGuupCDj35XY8
gr9XBKtDe4mxp2tyzscGW8H+MeaaysUyorFS+/v543VlThzcDJ0kYbH+jFt7Fma7wSuW8wB+Lo9p
icpttVQ1nZepOxAqzJK/SoBf4NlbuY4c+K7ovu2YnQMUmyAVHulftODwpoxbMrf10WjRVbYRVtkS
VnilQA6dnyDBL6Dg6Fp+as/wj4K7LVF4Sf++lTXOK7qhqkr4PfSOxTIsBeqN+wBOOyCT6QvpjQvU
80IIqpO3bBmX5Ky2V/lP/Mt4My1aSz8oB+V3EZ5gBjV/Bfk3/H+2qrUha1F5HXifAIeFj10B1iuy
YkZIiHVGi/Uvg5wYVMhfQ2Ii+2SEQSu7n/f+jGpkemlmGnqMKRmZaCPHHWOfwa9RDWgjr/sy0kx6
YlfRrz/Bb0ymrVQ4jZbXanfa1ZrAxP1M+dP9URseEtz+3qrMsXf6jDzOTfs0T1DXWc2QxOPe0GGf
hNWoivNmaM/KaD3X9abNByMyEEjJePZpoNcIl1sJT5BnVBGcbM3mKSmPgbVxMgKNkfXRaP7rkfA5
nKUm8CvaqPQBIJ7Zzt2IHcDdm0W2rchJz9XOncM1mflqz+eMdodc5Nd3D8yztKK+jqSVuGSJAArO
1Neq2PhQUT3zguzkL92c0QlWZmou2Kpzk4rwjCSfQaoAump1NhTg0Xm/1sCRlpBTs5sBxQZ9TwmC
K+3CLVNJBCsTnnij/7sql+EiKRRcKxhcS34JnHU2yJp1W68nSBCnOcKK5+7RSJu6XqfQOxp94yCh
8/uSGZjJcSd4z4B3QG6Gl04trPv8X+nlILwKXiHFGGWG57wSg4KFCZ3FZ3VG1Tn18zZesDwjJim7
0WAQi3MdOLDmWsO+fA3cg5b4/IAn/Qr2C0N2mEHw/VBtq4YLdDCBaWcHPq569+wsbbwQ5TLDp4MY
KAMhv7O7c60jOelm4lwxZty1YXOPJSNu+7tZAApk7zHa6k0r0kXts9mBD20bSAehMjED6kPhW+9X
rzV0iNqgeFpa5q0iA7BOlGI0voAL+do5qyDtIgYN8p9EDhcGFLQrGv/+wYyRm0y1oaOwQ+qZgSrp
/M/bzYdUW1JAEqtcQrZDqptSad1Bcr3OBQCOeasbUCVaqU54XvL2Snt8Ik0S3PVUGaS4wglXJWNV
Yvi0PyJFWZFGyZ4GxW67ymubV58v8aSpvlcI5LqhhK/nzmvK3iPe6aAGUaGTE8IzL5F0dn1trPeq
LdP0TPYWFebgxGlQ21yoLfk3+CI06NPtSJmnLd2MY1nlwRUqI1l/z5qz4CyBZEg+4Gos0IB5oi4Z
oudMgNYscUjkcybz3gYA4bUwQdmy3ddZOuOXdb1u/Mf+2tZGbR56tSWqsb960gfi1hp9FiqqfrYN
JPNvHXwAQpHADi4gD/EvXvH1zmgUbI6bZ1nyce9PcUklNMeReJ1m79z+R1CBs1lDztlWHzsAVLRp
UPaxR0iyVn8wxtnqVtb/DHu40cfAkthXR38ZVOlsydd4TWJjq4KkJt3CGDl0KwUX3EuBy8A1sOye
E17DyITSH1s4mXUGi+J1L2mrxeeGmUglxjh/lM1eR1r9xbV9wvvCmYTpX4qpkT2jSvCE/XmC/szW
NXHlgx1E3l/YZiZcfRam7ZsT/2k40b/IJvvL5s9EVfj5au4hYVZ567Osj06mjTKXTEkcaLwJTafk
i0oNk/xi0AJcrOdY+VVvqbcXrwUrhvh58hANQMAXwgb2AzbGCQUOSxnFXD8AI0eJafZBNFQ8MX8b
cE/kdUFZ11drdZjuppO0YSy3xi2D9xX7D5UhQjqwyJIC43uXAqV5U4+4EmWF0Xtq+cE6o+sfI2Lr
KL2zGMEh4Qz3YzVEvYvZ6pag/nxSbOQHETHGulz5iY08MhClaR28483pxwGlIUEmay9Deba+OGF8
61bicvnKhQame3Q9AAbLqINpSKJKZcUUxDF0WWxx63uzbx0V7lKfsZjYVWZWUR9k5183ZQ/hDK9R
aqexRO/km9hltGlorfTIQ5yuSkcbn2MIKgdyRhHGft/DR7yg26YZ3kC0OoiDgr6E6koBEAYNvGXS
fNKZ9UrkPZNHQFNx2H5io8sQRXjhuhtJR9pNolVYt2iyhwlBZzdsJpJpjyyUbneCMTyR8E6j2KIJ
466FWcTs4+dwJO9uLZRP7cOu0X25JO3VMcINICLjN8+JWM4lKyottC8EN/Sr1yOol7k/MwbR3yfF
Tqzukr6b+XKCIhqxiKbgKBBdCY/6ArEIAnSHg2Fr5s0LsFavnTxVALydK0I2X/k9De3/+qzzSXqE
N+6Q1YxlQ3rqUcEg55RQkfPOXGB0mVrnKgEHjqHKE9AgdTiION6RfsxmdCyIIL4VlDGMj7BDAuIP
3hk8BoaHxJ67/dFIXFDMIxvvYA5cF7hI74U0AUzUirzJ+olTIR6yhyDLejPVEs6qaXTEQHRtlmsC
3cD6SXgAQJJgv0ISyazvYOo5nlfjijaAyQ8QqnZM+pBC1Sh26E5IcFhFo8vPrOFD0OxNEnNPpfFj
NHUWWhero3Tc7JH1CsdVRY1lLcLDMH46nuL1uA2AKzYwyMnYuwRqprtWddnCxSJm6wpVixVd7Ibp
H5YFaRiHlc1j/SnIa3cimstLHcMJX23gaey2kgEOdixuxHoJlHUYk3SKocUiGUtopMECKSkTYEew
pluWyVEdomEgZ8VBGRAuMDI4UzAg7IB+rQu4X5ucAxRy6U7y1Y4rw9UvKIZn0qdWeraDHtoZphAr
hDVdf79YJtCb43k1LIY4K3tnEV/eu3N/ssdfUXQr1UrWUC0z6u+zk667qoOJ3oWqr4Thc8jdshfu
APvfqNeC6MoMGvp0GNtUx9ZVmiyNoCHKTYcJmQF1egJQRzE+baqXS5hNzP+b4WuDPkQrpC4WpMqx
8XBbfslj1Z5LPEq7gkCPtJ8+O+TAKMP2ZOt2rLeFgRDZtlSgcWanOfqtOSCCZ1ylZDPF5ZtkOPTT
WZYqEjqL54dHyciwUf9YKiTtBzX5oMmPu41TFS1IkqHvttL2/g7tvBKp2jtUf61LrpwE+m8KnwRQ
ZcojXCUH52G2opblk0tEwZGR/FJsIlU3xmc6pBNafZxOzsOJLqPl6uePjM+5iIHRNwhkaxIy3z7r
xQ0tt+Aiti9o/Db7pM8aF0MyLWe9RqX+YZU78Wt1NR2jRZK2Ps021TzRApt0vxdZvkJAJJw6SMVB
jOOIIspyXG9zTPiok+idiyT22+OkMX22Gpy06f2Lcd+wJk9/BO4ll1lyXuIbMWzFXt6I40gqUiNu
+CRfT+jpGa8j+StApl76JWWSGjShCUZAFKOi35MEQUUKyUBq+mxl/Ja9KsIdbaqek6O6xEfcbUtq
SSgqRBrGKh/qvAqPj/Cc8qA5QHI76aFYMAMn42EQvQdAxL8O0cQMjeQ8qp8ziaUE56yN/aGtgdE9
LLp2aA6gzHsi9/EQlE9SRPGCszrkP77g/H2QPtFFSlvX/Agbxmu8FvdteIj6aWjU1hFHXG2EdnOr
vV3Vv8tUi2CCWePsi+8F4ylK3pFiDHRvGOhdUVcnSBqZ2WZBGg/mz4R2+HTP+Cw6nFXONS4GjSW7
k4pkxfZgryudf1lUopbZqT/RhRCHLyKEvDcEIxZzuvuEKsaanbLZ34f/QKDSvVMpADsLCD6i25Nt
+fMYOREODlAk7FMNv1FC/F1atrUxg9zp4tsq+/2Ln9gsxk1tU8ITQhXmMEP5jo8FwRCKEZNVUihr
NvjaJI9mr1k1IqGMk2pn9JJOutdvsq0yPxWglmzIxnELEDlNsFXhcU9h9oVUL+cxeQttr1hEv6pL
r++dbGMw6gil0hWOdedPVLvG4hsT5qrOBQB+ja5FRmt192Go7ihF36TDAHZqCfbnU3+FwoLCaQdJ
o9jvXQFi5epioILsagDYI6VCV7J70pfHuQrMHDNojA/JoKSNFPmKprVdENv05duiO+ZOZIaGpc9x
trhfcE5u4KIuQ9wwVZJFS4mlWVkGbmOQb7fpxkb/Lt1kX1RIWw6PVbXpjDR6KgdBqDSzZsb5ouTE
jr3cbAgOKNtDrNFQC1PN1p+5VmNURay2/NQeBxmHyjtyVTcJnQ40oiKp0Mrp+/RySUF7eR9csin2
6iuSGAn9ZVB/DV0ioebVaqMzDvE+E6G8X/gVdv55SiNwnMXnIokJEztcLo6/mmlFvhV/l6F7q0iY
3qNfe88LlWyLsWw1h/IG9yu6VlkU3Bljuo74k3Fc3o0DrSUmkACgWL8AX91Faxku8PUQ0wwDqEvm
civSlP80EodEQqE1IDajGs335LGWUFLZNDAZqJ772ZWTCOQA1SzbaEc5OKQBen++X6HPBhpd9iDo
Yo+cF3Jd2Khg4fjvZKqC9hLO+46FUHMkf5Dacg2/jkN22oB8A45eDrE12rCL7LWxj9xHf/Kv0C3b
UC2pBnxsxp5fLvog0ExoTfi395c1mu08ose0pyqElXdiu5yVqSb5ApJZ46pObz9uOv+rabQ1Adua
DPZVHaoxUv5e8joPGUrpwC0U9JZaxSGgZ+7TNcCwn7GRrIkrMfvvPWzSiJL+ygeJc3ihZY52NTdk
FwNY2yvrSM38UgUlc26aBb8Ze0GMgptEkp4KjaDbq2UEsulNxZ3lpSwlnBIBGcpWQsfShjIM7TZS
fieBgUrQzWe/0IAMJReTm/ZzHfeTntDKHRbGa5Mm4KuIIIfndcoVAE2aZPYoQcC0O4R3VZebrJs1
ZrzBEAgWe5Vjm22tx98hRA2gBNcM5b+ExgM2z4MowgerlyaTOr6xhV0FMYTWdJgSDLymjnHtTJtd
s4nMY3szfuSOT04ls3mXifCPQCCd6copeqDUvylkQ4GMwIV7++LIgGrzv188NJyqHI/gtXAYGlKD
mSThxbptazaJUGrWDcO7seiQF3IyhtVCMeJckbyesWI+mOCMk8uaxAZYatBydoJVq39W4wI/AMtH
l7xjAVSqCex8YBd5kFdUSRNJf1rF+HnP+J4cGkNfW3JNICjj/LYMWkO96i/S4trdvDL+O/U0owq9
8AaoPM0dARMvyTJakeBRLo+XolK2Qhx1bgoHgvNx1HL8fVkknijT49LgSA6rlNm0v9dBsYc/7WJl
i6cO4GKy1Iv8MERDTywJD3+KB5Y6Ulia37YhAepGITMYV0HImMvuzocEu3Jk0XCQyxe+MbutW3DA
9/YbWAtzSqmPNcCV5VFNgU3SVBfbinuDSmUfJInfggOp9OadREbkoZveNmHKuE7uYOeqlCyfoWnK
Du0JiRXXuHVLswI89/W2CZ8OXXxjpUk2+VgQNuIj3kvz8BKo6pwPUfCcIoUgLI/8CuhElNFKdQfN
+CqdaBdHx5Pg7pRpTXColBkqjkrAGx6cXyVhWDQy6N3xGp3khjUhP2AeAjjL7nptZuJ9J1H+m89E
XxHzo/5CjPfr+pTxSVy2w0vPpfrLMcxitUyGsmQvETDN8akxynwpSOZmgy4Mth04qA2yQBD8+hs0
HQQM0WnwYa9ayreA2UfdXy3eXQKCJdkCtaa0KRoCMNPcVxRH4d2hBRc7M/Hqnz0P4+nhUD6OeTWp
20otqVHc8WzaKihN3TeV2maJQt+xigusdsgyBV9695mInn+O8tkkovq18Az+CuK87bjbx4esJhZg
0lZ+XSvPk1mYBezZ/3njJsIHsMOCojPLfCsEGc4TwT2khazgJDAVNAPopG3YRaTS6sltbrnSdp8a
nBrq77WpvHk/59VR5gdJdbMg7bytJPpT05VCk+Yq1bqd/RxmYpptau+ynKhwiiCP7lZMrPKSL1NE
nRjUxmPakT3H9qXm2tBp1Kr4bhbd7GvjNlCSNKbrzm2P9qfoAZWHN2ea6hlCxk6CJY9AA4GEhvk5
9+dSHbOSWG7o7itPFyV+/uTrbbw+JC89Eh6NKBWJQczXsyIrTPoAmnFpT7BC6vka+Sl6pJavrv+c
yfLjzbVSXqfTLvVvG+Qh6cK4Male9rHBxbqrT+eZpREhOxsehMc078PfjOXkr/qirBrjZilr2Bgc
+lUdCNmyRFTVcy6P6iFxDMEp8UFs+CRTkZT3yXyNgNHIdW5emqqlly54bNMCGVCZLPocoxw2pYFr
SfkK+gS+pJQsXF+KpEoKGgevyeUWb4Su/Xm+s+5+iXkcxWncf0HrzMpDpVCdcii3nab5jMrT6ySG
mmFIrwOKCfkNn5kAp+wWMxwuhyXA28maZw5N44cDfIKMyU8nNrnsbAnRcxWRqUlK/VElaaBDRS97
4G+eewenM/f8z33FE4mmmzznNxDCy7EnQQ5z+vSL5rUWbNM2iT6xWorFDE6EXoigcVibKKxtDPri
Jq2ldz9iLTwp+6uyUkb57H+DWVKTtiF4NBuP4UjoLnn5nq5M3CQjblsSpy1L/SoKixfK3xgv1DF3
C+UiguhCHXqOL7FSjSrP59QBV2zBycREiGxfSz9kHUgyNVD969aSH3EieKHNgS17hVKpLWzKM3kL
Z0ooPggOus6eKHixoM7H1jIiafXj2f9q5e0EOnJLXZvcPm1WMDmcosqS2ccR20Ed/5oIUhFeujWr
SQvjXIrF6StM73HUkO4/lNlt2nzIgxpXSKOjYm/HQ9tQ6Q9y/EmfDNdfcM8XObWKt3PCpnQl8WWT
Kto2FhQchYwAzbwPh48YEXi+fb7M81Ug7FjYJzCci5G84vCkYUTIL2K51PEtT+dVdZF0ZBW0N1V5
H1+K+JkgH0eiZEIJ6AN36WNI7Zw3BjbnELoAvSyCT9XtJuKiHJVVZaHiha3k7T+YSxOhi4b7myoa
q5gD8oyvGoZFeRTRzF/DwgZ13oe9Obm0GlFPsY6wjx0zYNMjxgHt5zpzy+S1Zk0szpnhSGvgNZxl
XLiOog2tkse4hKSC0qBt+ml58U6AG9k5W4LC8BfrLxdcV2znf1eQ0W29qz02SapAtl1GnKKuJfT1
jBUJMLzS9vNl+xQ4FerB/C+hyKrM/Rpp2RvD84YEogebvg2z3+zKGmg9TPn0oMQJEC00JgSHt7ja
BXM5SSY9KqC6ti+e2dp5/cCah86DuVvU5Yiw+YjqOquzPUbKVnXuPJqYKTcfTZxqz+/DOql8DmK9
SY9ppEfstWgAigZakTl8n4C/glx4p1ZSJptzzyjW6Hk+qzSWgJg0KK6ZgmNslB1y3EunuAjohz8U
fztTFby0Ph0aLzJc9KVFZ8oFPErQhk29ljbVIM1jeKBTZk9TMvn9QrRumat/8ev3E8gQqZLahipW
jkzEh2Xu4h15MyRSHxi/EYl/Q9DFTMmnt1GZNfC2/+CwdBuQqui20w7is5oJc4+JX6yn411v7B8a
3iHzo7BTPRomKqwHjh0XdWZCvPY6FoeHhLF0Q/DQghSYITwErMFafyB/2fjuz/uMFZTGVixt1tXz
aDLBRoaq9hHoeAC1npUqgAtaOcu9wcy0chPEFq0EDFlR4W7XAO7HhiHCVCKfmvwZlZXIY+dOU9am
Ho/+nIVifEqLMv2xk7XS6bXXjIWcEsoObywE9WOG+bzcTMYtBan3iuf9B27e1ditSOsi4CYBRnXU
7rTm9H+SHuj0bLMXbUu7LOaFhbV5t39QgUqw2w3ZtFzhGiRGbtO1PK2pxET/PdbJgRbJreSIjMHQ
lJS9BE/LdfTxhYaQoT6TQSz5/HjH9UcGTo5b5XAyj0Mhks9WOh1TQikfdwpU5mCHl+h9Wm7yfMto
7NI+OJ4ZhuUcytniHq3i6zmWzn4v4M84jsUpc8hQCInng0sN7UJpCShqWGlT4BS0eZXKAqYfW9bl
McAH2jUUsuaO0bUt69NSmc8oKBg3199kPRCvXEsDPfPDjwTvyv5DfbxDfXED+z3vafzQvh/w0MO+
0TTHlUQTIBce8GK2HKDonkvCdLCldAmi9Sm/eXGCOh6xfGIHLS57yMQFoYBh3tXDX0bKEOeWQBJz
so4yuWL4IS0zBwrj73Ox7yJmZ0s/MorSgY1VrNEP9FaL6YTSus9E+pgeN6eRlEHfdhYEwXcF8Ycg
ppSM9cWWtrkt+nHBE4pvl/kIllMxv9KW4G/1yiaVNIKvGA5qeiJc4xpnOwplJo4g2DbmHGyW8ahc
R9qjdJq5fT1K/ZWo7RGvVZxTamRL1GFtEiLGlje9ChyqTc/Tgi2h7L94x//ix08J5No4teL/UXEX
ZAdvxTQ+KWqfsraAQiBtKBUApg4etkCkILESZJUSro0iJ8F4SZ6+PhYxItbc+0lO2S6xWQhSPK7o
W0A8k83chwfcKrbsG9I8M89QhhbDUFsk7dk76i3DHZTgSSJCknoO350bJjsU2n/n7O18Rxis/IL5
oQm90BkNwf9hR6h49GSSWugvewkIi4i2FTPYwOHlXnZ+fTXG42nBKdg1sAe8ZXcoG+teSE6IaV/t
ucEvIiVChBGMYK6RK6jOCiuP7JxpGnOf6Ds2y7YcQnxs0bKvQYWNSXGSUmbJ5LGwHf+bjOWqnq6i
VKEkw8Qm7zFq9JagR3/D8LV0io27QulxJSQdTJBFJgjtbHEPCaHKt8Jm+JU3g5Q3ADHXOz9IIN3P
KiVdcGK69s19wVByDB1ajRR8TKLL8sADuq1t5/whvWaOLamakIVDK7Ko1mf4jEqAws7d+RowAALt
r3jdIP9w3xDT7oEzEl3TA1+1B9uvoZZGwlac36/40kqun/NRZrPxB23QTgwwnLueaGlnFrYa7wKs
1Y3L51WSINZAZ04MysdpA0AOj7V1t8wqYfIbs4Rp+zsivIjy38yHzdrqQRRVSZCmvxoSZ0gCg582
b5g8oP3TVROlMVm3YOksvIICFyYXdIYEgDzh/b0QhoETSoZc1rt5IVN87XrHez8n5noU9FR6hpln
ViN+1X+GAwOgy8EfL/FHfJY8E3hWA7Aj0ZN1JQM366Oui7QMYlWSd1eP74oJaAift0auBY3X5s8L
wfMuyGqam0Kx86toVI3B8wPRzDhQCQyMB6UtFs5kt/A58figDWW+Xc5XkcRWpRmTm5jO5exx3Ety
9wy1Si8xbmxVs6b3zI8sSnNKHo9uOYvzkzd/HwAA94L38vMl+ZJ9oIN9HsBHBnuXJnjwU9oGpchT
w44m9vUleSPUvCxThuEtvyyHlSsdxp898GMmBCFqnOca5VpLkMZ8t4JlLzCSk2ydhX5iYh9WcPU4
KnPiRizmH8Hgdzn6STc9DfX/UZjUWWdAyRXJ25am2buhqVzUenRGumrLqwYsWV38Q2M/HvgU7tOD
MKsuttSynthwS+hKhbgB09ZX6HO5gISq5nmemX6kb8v3F6VN7xf8VRvE9MSsLhUz7oGhUtbz7Yv2
N6h/K6IjjIOwaGRRO2ue0Nakq4Qx76c2owj2CEgT4L4ulXBgIHUXoNcDtLGy2YwkcH4S8uxVPErB
pHqKuKxq1IqH63kcFTJ8HN/P5Z5pHNhp4JMgPB/wXRuF/4hg842Gi/50BiHQnC+2TcPEUDqcJZW9
ONf7+n3vqcffEos3tvVB6a/mh41n2qGSRLWzOiJrJ7w7iKeurBYiZC7odfVR0GDyK9Rj/kfUY26c
OeI9/Ik+JgUyVZU2jP5wrMNHjyQTE2dHMdLALK9RpdOwpxquAT4kf/SkDnBe15ZWMONIum/BP3dU
Yjm/ZOiDawS/7eHoUjNAMNAmJCKldQpFzIr3vNxmK4jvQWl3mUKLuq6kqcCrHeQDeY5TAYga6rbY
8LMNsmgGAm8J4zUg9+Hkjy7vbpBULJ4sKwcGBwwM9Rh0KsvyIEUduoIgEX4MSpDBdtIX4MiPVnBz
FKpWH3tB7ecXJA5vvB3gCOwN66NhE7H7jEPs1Av8RygbB3bQ78GCi3SmhJCMzUNiG5VT5+81h/NH
tRs0ICgqODC0nQ313G9Xd3FhhQyQI3eqprraDuySUkMKzrAPrb2OMCmygkpF0ZoHi6nus+uMSEd/
B4KErOI2by3DYhoXdpDt1lHjaotRSA/WOxnQ5fesUpW5bkhd/CpTYY35wcmHbChDlNobNl9usMik
wQAmhVNwYRu2wNLieNSgJBgW284Xqhp04xlsH1hzez/FkwUjYR6PpcB4wMdtIqtf1l0w43rLJm16
EB9YC2x1/sA+TrqpT+p5H7bd+5eyEbRc4kyzGbkfuHCnIRsAkG2uW7o6i+h58oqRzTOMv4BBnqgC
lD9X/gJg1/iA7dn1JwmsuBU3Wy5+yk8p7aoxXc3zbWd6IG4VTKAmkjFLHksXoHkWw4yqI8yOYtII
hBhbI24fz73cZ/f2SNT+ba2ju9G4DjPzMGz5eHb49Sryj4MzL20/zij9uxQU0OGGbQ97shDCBLef
jYyibGKbaQXQIYeTxvdrczHf5/IT6glXT9HNxPLgaht24W8zhXxZ63yzofNC7W2i8e9PDQZhAiIr
eKjSeh8CWuv6GJ8hrKiFjvV7XmRTt/uxPEg+tocw+szHfUZLYq32Lm9yemwR3Pqwo4z0QEaN/Mpl
1Actp6mpsGZyjVTAXMlNSUTP9YA5NmxGyxAp8cR/CimW9rVOcUmXktDSH5NSr68v6XJUEyEKUcsa
AQEHnHtLWQlXyZSAoWu0ou1xk3rsIlw1tU7dDGyB6XZChRvCDA7depd27AIxbiBuRaTqEToyfqIK
5YYZUbaDg4eH9ZIO8J7tKXeGQStCxqynl7aY+ts23VbCqbDMBzrD9NC3GhDT1sp8YjhRRj/uGD5M
wcGV9sgX+lXXsArnl+1xsT3DhV47nWKCfFhcMrS17BSsb6Z1culYZn5EbO3MlvQqSxPuO+bP4P/L
TMlXTrD3sVNfI/GNuBExbhsNAq2nqEzdPWA3F1nQLXu6mKIRzsi0ROgU5f7DJFoNVNh134Oe/LWO
PMta5exgwzayYbQ82mAfWBITMl6+wLAvU4OpAH2d0bxWdsz+A3oNy4gUMTGMJn4xkjEWbBtxv1vu
T/1ZSg6SxNdXRd25dmZajedwj4yNDCod38Tgnt9Fv81ipIdSMdcpVbRRWRqX5QAD84nTWPkQBWcf
pnaWpFzQNg3+j/nKR5mFnZrrfmQE1UjmbsyfgbRJ9Qo62eFCiaMDPY4TaxPDO8cq2rf3Lkb8I4ct
l85v6/irTkLeEZBlQ8ViW8fKGS+jDjWTE+nkP4WUEmH0F+pJmAIcOyNcyn3QydaTJcZ9Xp58rHfQ
P7tpjmD3iOoQbdJfrso6eH+vqGgtmAXRqsmv+zRqEwu1ojen5fztLHUimYM8EInF9gzU8/mb8Ymn
nXH5oD9qmgXagOeRo8XqWrhVNy2qtU1VjKH9ZUg6WhaY0ixiRx0Dtwcxw+C+rm2c+ojNK6Xv2NLj
ns9MZ5mc8CFVtmzdKkruLOKJsTPvwac8mJEjmBFGZyMZMfMIFKjBWZj1yuOABLzxOFV7Q3ETZNi4
GLzg6gZOqEv4yYERVGwQygAxnkHeDy81YOyrLUscrzq3EZ6i/SMBR2z2/XuoE5sKXSQnc6Ru/7gt
5o1yccZwLwu+lYCQ7vIabczkBopid3gC2KjHYHZxlc9RBS+pXyHmRuJZy+BSPsJ8Oa4uGkCW7mq0
mzlplYHM6gL6Tko8f2EGn9ow16MeUYNI+oxlSs9Kv1aQTLBrdR5/vGAScTh59RzaKOFYmwzYb/bh
BhuCvPEzK20UCpwaaIpsBSil+n26dayQuVw8KoFtcfMjp9wuitq7+Tf7lb4pO2gwFr+mX6wHdOJH
D2/A/oRd54NUbjvjkzOsG5+nGpHn3zy2iRujKJq1kXXwtX1ryy37m1eKim9vSsJm5ewW1p9AsQQd
Uosln7tyrtee8J7FkwbwqAyOF31Q2HDJy2p7p7M4JLvGAGWoDrPzQTlrog88MIAseRqaSMNU18yr
poUm27uOUXe4jCmQEJgYXY2UR7voBmjFBQrqwRhSzklfafThH7n5ifAgdapL0IecmCknxvzqEMt5
mbJ+WaCT6to7Mj53H6A468UzWNlAxLgVcbeh87QvrpG2DACR+QQHyMQgPDU8N7trNAveJXkTp+lE
o/9i1kBi4PRfvJXpW37EJxeVvLybo51WfVGiRA6VtWSEiogKr83w17nOtZdSaQDyWo7esrwLEQsM
1PvGfQYP6vl3IZLzEXB5jLg4ElZLPybyKf/pb2s2oNgSj9gdeAqc5buwGKAj2cgmZEkieey7ITaz
dFhKsv+yHbj0+eZDYJVc+ncmVqlB1tRYZSGQrDamX/1Ymcl7RuGXc8N/9VtIpD+IfNighxg/7aay
nvEC5/uQf3J+QSfy4uTyGYWXZgLKOAZoXRbCt5Ev+w2yFsoYeeLFh329vd2mtGiQby7zGjfYqgkF
WV8fJiLfjfaYqSpuzJwAIpaTF3yhtm7zOvEI0cwFo+VEH4dMBbGYiwayz80peOZ25ppchIJfrxRG
n02Hf1NuLNZGv6moAVlAMXSGy5hkUBv7HKbU6YySuJHpJtxBVe+FulFdIuVxN5Bb9rpoA66h4sQ2
SWl5ozr/hipOtUivogp/+pW1VpNFc9prz81tCHbbsI7fWozV60icm8yTnbOxYP5xMAqdmS4KKmzw
Or4bgkhWQo3QYkFOEalRP0zbUz6qshTaE2y+VctsVkiJ7l8/FqQMhkgmOUAebAw/UJ7Ust+eumNv
6ttbDI1vYQTcjc5pOEX+8CNPoUAlHtQRZkEcRE1UiOgNK6+uhOy/ORYcKwdSChFMSyB9UuiUTlbh
vM0BqYACuPHTW7+1U49HiYPzXjPxBJCF4Kd0xBqpnuG4cYNiAwEu3JihuGTWSy6WtvUh4V9r3W8A
UlBn0iTyaqDbBR7c1dYCcj0W8yqaHhRKTGAjOyAfd04HJt+dBqOum35hRQR2ieLaGbq0gj8hXWM3
zNg+oRiKinhsacVInaYDJBzovxXg3RuyD3Wzgs9b1WtlS0knuSu36kRhuHqmEmLumnmcVD+EjOKP
j5EkUgPgyuInyVvJ2/aKHNvlMOWpzxrPQteu/UlsTG60QrVsKD5/74c3VfGcFl5jmB3tedQPCqBs
zOIvkP+Z9Pe47sEvjQRHLQuo/ds5/oRTro54K9FdTksiVWXOXr/nELQS6rJ7FiidgI1ERDBF+gvA
SvQg2Wtg8arx8zW0BxkRMLUWxMP985VW2QiGi5qaUxEZioteZGvzfXNSQKAS3KKQ6091Rd5ivQjV
xMBo0j8tX12btULILTMiqesKL61kolfl8HAwjXYyth/3QpdRCXnCR/Hww9hxl8iMek7ruxLfRRnb
+5Im5jdvL8quAs0I2QkWZdtTPI2K9RDA6jOQYJ8Kaafw5/Dj1tXRgiiKK5ndPq9j7Iz0DixbhvyN
8d0AQoRWl5LgqyoOpztnjU5VU6eRltxVdcqYkWhpDgtLlZD1Bm0jfMH9mDCVDybTLGMninF9GhfK
jUtPcqNFvfqSSupntsbs7+qDkAdX7r+s2QO4ow4SI5OQSNHI+9cRBuxDQ+Pv4LT2WdUdeJFgBCQT
kIQ0JJZLokMeDCxkXyUKAaYbPF/xx902PThuxL8xvPvqPDKtgG5wkY+DcmIQMZBFdEwJxtaNP0Yp
uOEObkHVGGu8EfRMGcvD1BKeU3V7zegy1FZHQ4Tbu9H0fD6VdBnOkGuCQoMaGX5lHRSZRK6C1FNw
vcXJF/o3TGxr2hwxDqpx821A9nHlergz/++pQwwv67yF2rRHDprERnrwyHoqLlVTpJx48b8Nl7RO
FTzLE0pKhNiezxTo7G6Xv/NxkA7akAF0mFSEQYMOIlNM3fNMD4rDbXvcTVcYc9aJcmSXZHNKzJ9Q
X0LBwBTHSavc+h1rQ8CTg/bK7avYuWZgVh/mGaLHrC/9Y5oZeme/P/pz/ypdBnX4ZH/WpumQfSPc
oif7ugLXt7ja7zzVeJHKXC/yZcuh2rYXty2MWc73+9HC7y3WUSm7x3nv/tovkc6C62UYnbOkxveX
I796c6qgLBoYRzmfORBoqfCVCZ5svZlKOGjc1vfF1o1YdZLkm4JBVDvLjMpgzkfihPgEd1mcU+Ms
LiiVGIL75GejlZKSlFtXNmREthhUoUBNbmnJApNK+DmRCIzJQnQDmTZpqfmXT+7xBiKk0oI1Jaff
PXoq05cqRrpFfDT0aJ17yXpctiHQpy+CMfqjLgG/tEXIMCjpVEynPAcd+kFUV9mwxbyyMcWnPQ8A
VhduNqLiufl6k2utcs3VILjWB383XEHkkOMALMfKzJHdVIjCEO++fxZXHIRPzeIj2PcUwqMdkzSL
UHb14i7RvM9EMGP2Qs7Jn5qBu6Hmgt4WFfMc4YzYzTOSkn7308SeubRT4EcnZGdDzCkv0nFy7QPX
oTHIdp+vhJx+7c5QYxljoTq6FsaIQdvKVoYwuCjyDhsDII5dvKu9ReRjnUY4rVw1N6qWDrD92lf2
N5442NWbYE/bvZ5c86Z6T+Az4OFpXq9B6Q+74ySJvx1QlbIXgkLPqhnNhphZyWWZz4PUEaa0hsjb
4NYQLg0DE8H0gnFnxt3Ga/S+lui9IRj04Mx8qW9bi3BcOrECUWEQllnTb0fAjidxkjfQynINFPQm
1GU1X6wVIu5oOqmRPjCXtnm/AaPMzeLrItsd1XpMn7lS3F/IrK4SHxT6UnlnS67YvxpyU2QzldYJ
jBLohFmbyMtut8MgRMEcawhb+aVgzNM8a/aysUlfM8idLQnLNOw97gk7HoUUvWeGoFmL9PbichjG
uTLx4B1VnG5nsYBObE5LVgiyaBuveINvLvK7mQPuRVNkFCAXJ/vNjCSegYR+I2If7/WnFKfBrrpc
DmJIDMSWoNfG3JB/9YwsY6fOHyyRkEKPIfpmYI/qT1ID6NB1LbiORzFMe+Dcy4GvZG91FA6TEMiz
u9Z4pjZJHjPZYyrIxlCiXZPe/QhWsOUQ/6n5ZIcBPx1N4vbGx61BTVKELd0rKOL5Yg2m8fUnP2rX
ZWLJ52atnozNJVsAqtqSMjBV5HIy1vAyz0Vwry0ZJiy1mglIK198ZrdVKFTXisHAkFk0GpQqPJZK
GgcXW+WXLSTKn3Mu43eRCcjOosGIv/iVvLlqUtNFNUH1bLlA//MZ56r7tzmk6P+u4bKHwrT0y+gD
Y/Ia5yZrwfBIzdnsUu7PHS5bdZVsU+bSEAhnZvIITRX/nYhaGHfubx7py6RMbMhjXmZqkEzfhfq1
s3tRET2K+br362ZGE3ROkeUWyMkHBqtjry2Dq6cCtkXM1AAU4ZJjAgLk9PT3UsyPDp36zNn7nMaU
Ib8DQ8YsALtqIvfaQC//FtrdjxeRNkfdj2pzXpfyxTd8hdEhF9L6obM/+a8qkjkowaQQxurMYP74
5yQ2Ed6HsNTp5OsvDEj/3s5c/u/cKgLot3/WfJOT+duagXtZB7L94ay+OuqadglUZ71GOWuC8woN
8HVjRVV6y7n11exJpJBWsqWlTD7aIBjh2d9NNKp79xhZoxBZHP9iO8mxlV/Ph1/3ZNb8/aTYYYNG
z5bCfSr/q/WR+s2V58+GWiBgkVrsc6X4TIOprUAdR7iXhEGmSGnCcCJxU7BGlmAOOlVw2KxI0c4W
73f6oMa+LZHG44owRVV16LZ7i/4QPNCUMJUVLbzF/jJlVzLqxr2d9B4Lf2WHzqH/pIXgXRytX7n3
tVB7/TlFTtFVo8uYEhq+D1woiWCohrLYGPNorIcRycrHifwqszHByjlmWke+ImwifqVCMZqwkdyZ
KPojUT8Kw+d/8roCJAi4ssW6BOY+ZWF9aQEIO0VY2a39ElnSp/als93Ll0H+MF7b8TrZy+9scrsT
o+HTfeJL0XCphlAPEP3WQf+6HV1KvK1g4x/HMHChZGPg4uQ4HROAC+VtZTvMxmhiFfmS7hYTD8tQ
HiqhaNgMaTIjbsIwLn6nPgonVicjxlqUHeiwY5qheLsGC8qp5OTmf4pgbrwxmp2236Zjfus+kgfK
/KR0iBzimrRqoALiUkGEUWIU3+6hJ3jr5woNBvhkknJVT/Ln/1nCT7rlSolpVfOZrvQxVwWo473p
cvcmJZ/i+8uNq8MKf9VW7wm4vVR9NTZKjjzMQAVZEXEW9bcth4XWSg8riHTv5//i290ZWc87+c7E
ALXkbu8dV1u3EBSvsl0wdFzBKO8qpvLTG9oYCTaAYQ1xElryfqxZtXUr1vRhJrXb+TwK/lxM6SY6
1QJcjuaDztKGv9C88iol4Tr9GJAK7LTM/LRsg+AXAdUj7uVyy/OrWGJRzuTXB3c1oz1PXA9ORdW+
H70Dl6B6KIu0AmX8tqXgERp2cLOnk7YOB6pQb8r2Xm+v6ca+wNsfGA0TACuF2/eOYB9/2fVS0TlJ
G+IiQ+nPm7oWKGXBmpm8pb9daOSkKtzY2LuGg1sblJx/rjbHf+ERPQMdFL+SGAifYfJF5qn9tW1f
UyaSGxF/UfkQG/TropPMI4Luh2IC7bZp/fVmlYzg+983hW3jgWSirMnv4j3iLgXm6inQb/1toa9i
35IgxrfOjN3u61uTrLy6QghN+jcxE4j4+mHNwqyrl6S6FLcHoOCJL80pim6ATIxQR7zQ1ynRy6Zu
NUHmcWSXopYBgHmImdGEPpg2XVk/dUmS6AEq9jNuYUBh5lGj11FPI9WPpI5XmujPPfCeN2JaW4PM
qNp8iwh59MdLWwReXBGYPmfse1BwcAf9s3YK8LEDoygW1AlMEg9WHvjmxlEawn+TiH7edZkv7o+8
4qvWEC1H3YTMCrgQhKklSYBqNQQ8vTY0gtblGZhd5fWChw9IawHYT0qI3gpO4bHK5de+8O/s6+uY
LQLBjaNJ7g1GtmbNUfWfUqX0FDtK7iC8sHBXIp+xr+cHLYtLE5VnKS17s3gAbQwcy/opWyT9XbKy
FG99EbFiXGiGaPq/54daPoqTMrpWY3boMAJ6qWMT2aXsfhsc3bamzvoOPKWDSu9Qmnwema5/YB4j
xOcfT4MeFs98CDVd7V+u1cvI2Mw22dzEzRLYBQ91KLW+qkXTqB4BbK9iuksZdD9ogToOVbtfXZSA
8f1sBjUbHrxjuzs/+EacaQg9SFoszm9aiYjpafe8L25Tpgbm4ATdmDmo7Cnw0cpeinMhtpTpl8rU
eFlZ2G4CGYpcLSnpHHgPIhmonV88HKJ7tT94AtMygOwlwH5IEARJex7XSIhc0maE+jQegjuazs5v
83mnfR/Hzl9BBfY+rLIsxTLcO+YgwdRbGVjEOn3wM/FC9g+UNAW3XoiztyJBZmp6e6B9tFebyUob
KqvlhbIT/VwVPv5k47odJFQbBx3IjvzvrWWzTwESptT7hggDQoQcIT3JVwY6dYORELWDD9F7QEFL
9U4waPDI/m+YXqm6/oaG0oL5nYq8lTY665cRZlvvBnmrFrbCWOwVcnnDL8qA76Xo0ikOcqhuLLuI
ePPX++AXjnUuhzMkBnsjgyiR/REJrs0SUv+o4Q/rPQfbi5M4QJ3oRQI6O5aZm518MRwnIK0MnuUr
Y7WrFqiMg+ULGF0jl8fAb0TIsd26sGlzvirQOrpgjA1OFanlSk6264sdTZdLoGsKFLySwKjV3mzy
kynVfa6tJwF73OrjWDPTlU/1igQDgpHVmmN8Tlf5VZDvOzGzDwGGqE9re967mXbPOvsCG9DwMf/j
UfebqinX6A4+H42V4Vn6JM8LOchn6quTTSYZ7c8XKHshHRgnzsGor65wCiLjCz72uJWqEpQOjpae
wZsRmQiquww46Lz3M26lRdgjzxeT1nYKualut04MRM18h+jBd0CFI1zXTA7ArV4YI+DbGEmBuAaP
lT3Bow2ACjLPsJQrCRRVv10XWDgz9Dv6+4BfaipMxqBEw/EWMKPH7wZVxw4GOPdGNjm1DyHVaSPa
ZxakR39NWb67mYnmq/kPhm1vBW/91wEFJAa/HQoK1MFM0UejOfLxwXDjTJHP6RndBrt/nIgZM+3I
dh/97Th4TUGV3faJAIuPGRcTiGYEmpPgNhl8H6h8q+0JHK0b4uc6E8oFTS65ZKVWYPS0nCWtWJaL
BJ//s20DIo8PrwNc3Uqt1v/klbb2hvMW0+UkZcLNi0ldBEOjlHDyfzGMJIHDilmD6pboJj/ZZsAr
gywCJAe3rl2Ev3ri+2kQxOY1UmSgIWuMfxgVHK/dQvNkYyCiZDn5Y77CDku5GN7ZAZ068KV/XspP
4M4GzyNOPjRIYIg3Fn2AKBbpk9y1kBeKfuYuj/HZ+GaAqinQc3iKOzV5eq26YOUjbzuuaNo0foO1
0l5t3rtrXitHCu/6G3tS7UzoXu6dWBdUALNdOfeJOV94FfdSuDytJB/QfcZ0nXO+7zmEeHxmfL+o
YXuVcSBfTTAq40ELsGAwEa1iVA+tzIwq2VALGCkmO/kAex8W5TH1Ap8PYMXBCje94kM/vQm/pV0K
dizGu7iZ1F9F2K2FHd9AVhzuWjc+4fOTypTSf4azgN2V+c1eWDEJLwH5tH5OBfFo2QHMaqIU+N6g
sKxFRjnm/gOC1ouEP+1W4YxNQ586uCMFpW5JD4qjHgjeIEqvIyzFcVfoBKenzbiCORgCCMR8cEYf
+sGMtffsslzIdfcR/r3y6BuQHCzXgktslEPknWBBr1jO33fBuGONGeDCp8wNxK8eyb2xzRVGOcQZ
cNrObPrACKDTv3PyCT/+c2GOFvYpbMhUFSrlQXu7xFhikAlW5s8X3+1XVPmgw097zSxCgqmp9uMf
+OYuogpGTODRj0B6O6Sab0XL+/CywmSiVAfQVos9KnnrrMXYne4IpZlw7QiLjNT6NORIOjHqDgGx
0HD1D/cAUZ8gBRKTS/7IVJYelyUzDRT/8YCGjjniFhr6mqDWDHdilSk5+ctyw9UShiANEen+KqfI
t3qgtgtCE45a5Z68cGZZ2NJ8CYdDujX7pYMpNkEShoR1nzK14w+vcYOD2arZxLr71pzZYPNdggwl
91BeJqfKfxqQaQBSCcd1ljHrMt/xziCYSkfwqURBNaJrqgzNyG2Dp/3cXrY0SkjhDoqiArApHZtT
CrpQYSH50C4e5UcyoiSOxq7+F5awRBY1gKu4VzrLykC547hOzX6NglPF46uBB+jPnIs2+KKeZxyy
3+bSDwSGmJ/ufHhC6RPXsTEvS4ZY4Kj+Df/tT4hmcmzO7TzK8zx0/Jt5GOS4CQVk0niCVQaOO+1L
lT2aVOWoxb95rsHMvlzf9Orgcljuyn8aG2RPtVJjMs96hd8/3lk1bqk64vPe7n8ZjIoEvnaQ87FT
neLBGyFHQ2dUqLAVFQbq6LPFR/EvJpoVB26k5NpPxv8gKNnbadefJDUsJOnWuGREjfoqBu9zKDg4
tFePhdIGOeV61Z9Sc5FFUOv/21iCN8V1Snj6I9D3PTc4tDhMgKC3vyMF2dGLnyiVUd1wcMDzd/4J
okE85kw+AkoH2F5BilvpoJ5fBc6podRov1Jzogx6V3etTKFtzhK+QidlPN57E19uKhYc0OKx95LD
dcfoa3aYz+GaDMicPV1apYsLrMaZbgL32z8fFqvMkcXu6swoJ15LDgjd69wdL2llXzRBsxujCPfm
clXizWNlXDrCZHkxqt/inIfOVilpHC4EpKknzOK2TlotSdAuiaZFbdaqCgAxI9dmAzeFkAQboF5M
MIiA+bNDI3qNzfbIANeffFyWFsE6QfMLhm21Pq8XPPQfd1B78SmQukVFugcLxe7hz9vyJDQg9hdI
6Qgj73jpCgfsl4YzgUgPlC+LO9nuKUTHsnZPaYxSrmQT0gJVu1WfCfNG0gjMUjW7aSHvFjDsULhi
Yars1N8HqYTIhZ7brFSbwMVFD4rSKEzkFBga/vWQh4Km8Q5uNpz9aJDHgou/PSsBH0jRxT0GlVZk
FrJBu9G3zDodAFX1wgn1XyxffpaWVLR7/wi2oNSnDI7jo+aY+FNyMtZocbWiyy1KBp8/Ri7Z9Msj
ehH/vUlafY1US+0SNBPInCDdy0M5QSQLjIeD3y4ysIeN03InjgPr9GC8MSCQj8rHuvNtZHIF/ozZ
sGuAPpZtUjlAiap6M8LOxiwvWg2B9jaU3skQfg/6fAoerPKDRxETV44oFyJuox1LLSHCHD8QTXRs
9LUBJ5VG1NlvO+Uqd9bRY4L1s95+bHKaWo7u7H/OykW+PjfZ5p4SDrZzYev4mlrCgODU058Aehks
fPa2iQFdrQoApuaMcXDf/zdSCbOsEHPYxJCUzZJI8dwSqp/Krhz4uM+PFzAbCjtkQxanysfY9J3T
gjwbARXQodsZSDDFQ1ztMGyhJZWm61+w9DrcUwo4t3DlNxgisrYqwfPskdHh/7MY+R4V888xrvKT
V+ocqc8EyeI3q12aqdps9q7XiIxYTqvHVTC0noLE7St+XNTGV2eZhqKcCd4CxB6E2MGVf26x/z5w
elWHQvuJUc10knPfDXKxGwW/onsXh6oxRj7rG54Z0Jn9cpnlLflumWbamX3enwWihp5Zhk4Ts4I2
9wWcfNW9rW52qBIt+6sWnASOpL4bathi+HQ4q+zs2mgrcNza3HW2nvV8IJO6AdSpQnFWkpMQ//Gq
mh8xR8gqkrAJu03ImHYvB41McrXi2J8xbEvkLk5ttPv2jrugoWAszu8S2X9JLNzOTE8vHw3t1URV
GzIq0c3oM2tGG+pgT9fcpjdCwOVB1XeWJ1pwwYO5rHRWUFUHuZuS5g4r4MJeC4+w4Xc+RxK0xLIk
nq+uL64l1hq7odXD3tKgrU+kFJvAodRSqkDbYnjEbgUsQCDFlYKp7d2ZkexzeMC3CsSsrZBnWarq
2i+tcpJKGiAt8ivUW1HcNh62ijFYPZDxzBRdMYWrOZRjN22hWxq+ritWoWt/VByRynzmOiMW+fy2
2rxoE3czOAqutlti9jN7bCaPOcCJyeXGxxEjPRC/uh7tnO+/y2ZFInr1oe7t104dKmPdJPl3a907
nVZJoV2Tcnsma93yuG1FcXKWKfJnkAW5XT/R6bHpa8/n8RmRJxJq3AxzE64Km3V4duRgBkQ3d3xE
Fz3867EF+/Ic3hTwbCbKcaSD2DkL3+ZpOLcUMOFlqHixEjg8jxi6dRk4xMfJHhBkUk6hYZa7Dd6v
kr5UiDjlwuhF3Kjrk5y3sU1709EoScRWkAsScU8xZoBUUcsbrjajYZ6fA3WJR5fwLJORogINAw3X
76QdfoyekGrDzgWbXeTqs+D2ukyP6qcN9nentLLf6egZAQur2cmYUx3HS8fpxV/wN97oGvX0RF+m
HLoXm1UqW8wmzvE124oYOoI8s/MrlIlAAskizUNYg4P92gHMrUO6uBuz47JHAlscu53FOl/i4T3/
s/9Be2gqdLaRKk8ZsT4DBsNOx+EIQC38dsgOLSKEfhhwYEnVDlioNrB2iMqU5wEFm9fOAU7PDVMt
CSVm6gifYHDEnlLUe/H5tsln/kN1dy+IrfQ3sY50HvxKMYo05OXpTaqstCyy6PorQBOHE9rn8Tb8
HTK9Eut5OerNADSKiy1Lt+MZoYNMDKHYUcFi4/MUlT4RIAX8ZBlUj4bocxgpsOZw7RoRAzZqHzrZ
e+qxKkd91XM/RYMy+YKMt3oFh+5DT5WQZGDiBtpyo9AF/kG/SigLAWojioNls5WI+JDkl0x0/6IQ
zytz3Tr0rSxih2NntUXwOeHhrfE9UKfMmffXBoerWeTBw27WUrm/bKVNXBczdhNUbWLPPk3EWOHr
VUXA9I4wns+iTRU8FRqcqwN2PEUekv9oKt/SBrumyimgEHk7A62FBAR9HZ792Ms70Q0Rg9+uR4Fd
nJwrMdtjzx2QWBM5qR+ukdP6+ulBcthjDdsjJUOxIbnrICDNL/LKGMor7I1JpeBEEVHvMr8tqAD8
B9bK0JA/0CRPRmEdaYcscdx80ihrfUgr2LkF2vX0fzx9kX+p2V4Vs8LRhXB0l5ejwRI/6281Njcl
FNXuOWC6y4jMeA3MssksPIELRv/eJCpZ0mVQ4cCBozNrpknH52Bjqk3vT+eDm29cV9ssRUTb3tNO
0iOvcqAIykcf8/rQ/CMV7z09sWbxgwhHiMBh4xkTnaCAVUAVNe2tADFE8Sqpah+bIalTVsuatpXE
qrwnxfz2zwdJPeXK4BBSLHQENaSBd0TS0m+gwp3j1kTvXsoUUdcVgxzFmvGO7fwYpsfK6CE4eR8B
+UWgMHikXcv9kL2jg/2x21mA6jyMNBsRUSlCfTM+mnc883j4NlPZfTPzoo3GzEwjy2SWvIvNkO9r
uXSFynNFt5HjJavpfYVO+nD2AwbkWgNOP7FflBWLazwlFz1QviSrvloE2983lo7Cw6BGKebG689g
qmComZecS0L0PCZcIg3e13CTpq0wNtQlq4N8X+Jy8VE7rs9IJcGJ11R7VhqupgICLOnp/Yp9QCel
r7kKmFdUfXBjb8fHSmSNk3sUFqg0N58cvUOwUa7eJZH/6GUTjUArmxLqH7RmAqCT0Qud4KBRtsGq
MrnKA5i7PvnF6PTKfGPTBY3y1UQBunmcOaEv+NRJPxjFSWZeQrcWjwcRMddi1TZpH7z1yslfMSvs
wd/6tCwe8Gwmi8m/Kqh4eUyjf8gjfiiL0IP82c4ZYWeD4Hok4olRehgh7kdcxhFHKIzwlyH50FZ4
6Nj8sAAlz/x/EgagS5vsal/1rsp5bTH1sulx+xqaLOaaTXqo2j4aNB6MZiKA87P4fqHSF80x5NGt
Bqm4/9imBM+fePnA1+mCFX57IGJZiD8FINs242NdvTLIgWmkpUwfp0zfNl2Qw/VYuQe84092zo82
xKdmISAy0hh5V0PWg2E1gYf2HcnEBBClhbQelIKXgHSqMMRFQwwt9BFSdwfHah75y7beZhMB32yB
Bem8Lzl40P2JSoZQsCtcT31yf8kWS6cEL4LpAAYQ0NbiqI6579dZ44UP+qfpjlaXK78atl1b+lgn
E/4zFIn+MqRLX2Xox8/5c4p+aFA8uQaSox9cWZ/eYUwBurdna2nW9Q7NGX935madLc4yFKJEUmgF
aVZqc5VfpIXg8fjqxHdV9NqXmPjEx03vJNzdbA0S6mUvlZJsFmSO40aM4tZsQGz02rq9TH+UZJdG
qHDCV/8noboUPTSL3PGSdV5xl8WbNrINklOZrF831pPoRXkAP//fXAbk+Yy3b79dJMqVkgOpO8H1
2Wu0ko/XsDfUvv9mlFUKBG3Cms98eA9f8AnOLuyN8KpH0VCtTurpSU6hA05yyFm6lE5BlBczivPg
HmKvp4tfj82K7TT9P57ojSCWmoCVBsK+4a4VA8vvZyiGijQo4V0QPNfyoaWGBOjvr17hV+DwZScW
hZIPSoC0X8UMjHTTE8XI7IpsGHJU8YJ2zpEtspphhrrEkjXbImon/FZVjd1aJuGX1hczfwpYep4I
yMtymFfb/CRnc46BDe5Tbls1jMERzs9ojKkjRKPs46BOSaH5URnJYC+rrCu08vB4W5mxRarRUZr5
tTclVdiSD6s2Kr/1uKQaGDiO/JInzkM6dnKKdEQwXM5g0RBFIhd3xcv51d7FhlJXdbBdHvAQGOsj
feqRJnwzeNcX9EAGq33jLcpyjBz+prwO3CTEqE6ciwxyydp7cOukodLBCYFdJpBkqlzttc2JMheE
kRho3UmHp5Npof7iYRei70ATMexRdsMgVbgYbJugeABQbQBruSjBuFN4DR1YhUc0C6sQ8aP5TQG3
U5sGsObfonbqprqYLsZ1KvShGaQKZz/Sdbzt2I2nca/uomgnBVHTnkcj4zrmcRpzFycCDjhGIb41
l5XFAqMDd27tx0MDakyGE+IHViHz6erZQSEuRaLw3aV2hDyitGiSP6tmEzTmBvM30RpYZfxpS4y/
ReiNJeaaAv4p04KeftZOv0kdNRDKUPoKT86mmG0qKjWpiATVHn+wvh+e0ViUD9KXbx0Hy/zenewG
SxuNt8FPDOdmWW1tpNhyzAehaLfd2z6F/lP+iqebF90RW+NpVkZUfkZBY7cGDa/R5tU4+mVSQzY7
GdabABIwBu6473Wnc7HM4Ae0rYAkGhYBY/LpIuUkRC4wkp9LWGOeIBIZUNpEAcJKAxRCR/smm+ft
77kYxzEELTN5RqEU6bQfu2wa9MaoA5MmN6z1sQ7DVNgQnSL8viLEdI4RyTeMdTQ/398kZN1+Fmy6
iNWdoIKC3sCQc2RESJt/mA+jAfvd/ISGqoww2zN9HdmwzNOkLYBkwo5tKRFalcXZ+7FKwb9YtoHM
9DNIqUpcj1/LUfkHtPW8shhuu0azpUeem6JPNNXYkG5beO2mpz7Q2SuEIiveNHzTvaSPBZ+qYo22
gRXeZZTke1ysRGMxvTQ7gBPyFhSJ53GfjbM1okJ/mA1hSrbdk3FInHp25Y9/CdXs5ApAzcGg73RL
O6FFpykN6x8oLoSU+QLomI4/oOhw2oCN/kAbxhkCHV9aWjjomyRxoY5Rcv9sn59DD+ZwtzFmPkve
uEqiRXKg9fYJ2umEk8Z8Mqv85AONbbAJLMk7+j51bK6E0kOjXwgRtdsQhx8GyFFgLpXW1nG8MGnt
GC/IhDOzVVupbgEHTU1L6PHrTdsKieBM2yHJ3gVoyt9yFPcmSYmK0/7/ei/E0DdpuNqUxCVD34ek
oITFZ5SMRNlpMAQB+kQzWsC/ELFIUrvaCxHxgUtEKruSuYX3xeIJgDl3Qnv28NZ1UZO0Xz9LvaLW
rADz5T0OfYRN9sZ1ULvhojFUZ/YqypxH5UusQeESepaC0JI+wLH6v2jq1dsdASEQ2X4E+5U3tW6Y
qqbMu79v+EFJRZnZvSO0TPPvDTSJYu7kLD+pidhasTImqUGLhKJcJCXkFGuMX/8bbiCfRmYj06PR
NECeeJRptPCg0wT9rcpw7mm4D4yvdxUNwG+et2k0oRtbY4ed/eC4Xwy0L6JYVcugyKET4TSj/Aib
yjax4aTchj4axdytIsGo6SrR2PQ0HuVtJY7GPENfZ7Jl/MY6ZoQL0vTVQw11TUbGKHl46tGVo7cn
qp+VD58710IausiyDX0/7ai179cF+q2pZuTbrWAL7ty7LU2cWwwgUajmkEaGY80BrsHEJ93xXyyA
hO672RymP2hGgnMCr66MqYFRkD2jBrUB0r9GAmrGn3AMN6f8tVO4+Egih5vttUgP27CYDTJFmu98
jLr18wnQoEdBVxTYNAeWJGpA+NI7sb5Qh1FW/4b3MDLTClbCM5KzfbxofjDIRsKajUV5Yh8qcGHs
T2Q2SMN6KD7nU4b9P42XbjmFzPq+aXo3z9ague/REncqqH/SBmRiImYjH2CdWnUPWzYP2IhDTJLj
t9MClAzSO8Eff7eK9PhMBlI+tqd9HjIHoW7+2W66HLOCoYkwI+/CkVk80ToJPE2RqkBTqPaUwluK
T7OhqjI3d/sxWzEJjm7So6jaMrUWLKh1/tcl5DEYLdskSR7DO10rSMICcOCxtMfQ0XH1LiFK5MTs
Mda4LYmGK/9Q09JU1/51Wsz+Qmrg9UYMdBnIh/feXYE/4XySM3LsjOl0G+csFW0yY8+Bjq6c6ySQ
fGEFd4dqFW0sWx2lhN/I2bIy4Zpw+hsBTouQpBqfiR68UjKJ/aAxwvbPCAwyLlAolp+mECh5fsol
Nn1znZ01awT7DlCukotJIFPEHa8qNI2DilZnwKVPzq1Mbf2Y1i1GE+GgSWWfqyIdOjc6qHe362FQ
4YBAwQwCoNV/x5cka9s2Cx8hBD8qPysWngqfaQqyh04XZ7JFx8H/kzgKOdKZEITZstf8wziJvEJM
2G0vFl4lIII2wsBIhWW8KZ/gvmPRoHriagqttGl2xR+8tzplQNdh6pNAcr8AUNBJy9bS2rzARXgv
8r197E1bkCq7y0rLb6kVVJ/8myB7rJ07pdp9pVuwSbLPb7k2/WWxkpIWMxI8dFAy6rErhTej/vKZ
QUjeNdWTzyMic74j8nKQbE3XoJUYi1F0w8KKXpRllcs93khtAcrDQt1LHquX7GmadeAos7QOOGyn
/qPLD8cwTzBKCal/GBrtH69HaZsIee2YsxSPaqmihvkXXMJzEeFssoWiWNwf2KwuAdkV8moH38Lh
9yr0XKjJz26JdOs2RSu7jBM77nmPZv/6e/IlJYtLn46KvuK+JbhJe8LBEJmt9PxVsD5upeKgL9O6
4iUraL3uhv6eiYSpXI9RjSa/zZ9MhSMSq9qU8Ld9iE4t9nULGP8UH+JeZRnUuPvmk2MC3j1foSkd
W0YEueNkglP58+9f1U6gd+0lFFbKrI0Y4MxjxIf9HnlfDP9SN8Kw2Xq1GQSiq6LiJKXaN2uO6ocK
egOzpvh87rnPVzxv4vGcRzTqUBa/mesqijhgBTnOiqquJf+8UhppK2Ksek/v0gVNCDz5x0stJXOX
3hx/olBoXe1XdiejOdY9gbMpajE15fgcFMybs6YzAABvcdc3po/KgVxlNyR5YA365glEe4dXL4gE
/nrZTGt2zSjwZCPSfzth9Ek3/vFFbKNHX2e2GdQ+bf7FoF8jqII82IzZZVA0je3FFAUSAyxMx6GV
adqwmQRbSAkhfw4wYjcwQmLsidcufi0gLXS4xEMh7NSyyQTB9p05WKjvhs+qqoThF7VJ9Sjg/ow5
tuyw9KbyL6oPmJf16RmgoPchfa9CULH8/AHlgoG5lSe4/YgK/1Rn5XeZJUP7GRMDJAoa7ZvW0tmO
4RQLt3KskPe6oargukN8pqKSW53EaG77haKHCc78yGk6JRtQyhiLUnO3QKdZJJf1cuvsHPhOEzmM
E1kyoU+CsQK5hVY8MuySS8wYrafAhL15qwJvHR49Pj2mTrbABJm0VhV8KPKqZzA/3vTgds+ZtpfM
PEoEeO7Aao1gFbjfuKI9uMF6uWCGjvbydg/kbCCwu7JS/Yif0+5IVNZhQDTVAMMbhAKznHAeXIRV
EGPchVfbCBsRYgiEEA77o+jse+1dGh+6pkCjxjHCOIdUYQAupEFHLMU3yX86ceXD9rjvRYYqVqv7
EgmpNSF4LFrwXYuOWetpiCtkSXPPjyv+yjQ7btxqaWozgTF7mIrprqcCRpShldH8hRxAI/3RtHYl
oFO9CgORcKrMXD5n3rQ2kmHBdducqeggU/+EXYcOB7LkRWMCBzwqN3SkykSSYLoXP7mqev8PnVyx
GWKic+CFkaBKmV4BwOXDS9Hqifx7DqaamnIQYffZXwdl55vOP+ECxJwmHmL9s3BaKyGdwoy/ajV6
2PPcZfDOGhnUB2zPUnV2XvE9cQ1bHz7RqA0Eh3dorET57eH96skwhJZ8mchg5o6C5ILDlmlTDxPc
g4zu8/a0s3R/aax+ge19JFG3lLBgky92Ie2bDlpkkq/ZBr0vvo2h1fTGl4oLuIUUDHR3hIrxzHLe
7f6Z0hNsUq1+oB2BA23Mmkrf0EDvmLxOfJtxBIteTN3Vx0ey4z06hOaOPGbmmkc7N9QT7XR5d+vG
0J8q7+WnLqkp5BJ15lmGEZqtGLEk30L6kRXduXwOSgQgudmUQ3skZCfEfRzOzqP64Exv1kgfTiNT
ieVjiRlR+xfH/N1EZDn0buYtFPPfTe+KsNIRBhnsHaJMEZnnkyLAQ5lQ4LV3BJyLVQ4FDQVipFEr
IULjFR3DZcF1TfGJp90E4fGgQJ8PrLgC4uxeQjx2KxUB0c5jndbgn+HkBq9195+kiLrMYkULHwyV
9oBbT++sUDwnXMtwVp6AWYODu8AiBo/zrAkWDJeqUbMpnH/fS91L9RWIaDVDi473wp05FTzS/7HT
IoKOKwIU5sa78trLnFoY5PvK7MxX14QDdhv9v3uKRhJes3wbstjgyr9f9dYCerKdXurCiDTe0kD7
T8afvh6ZU40FSPXS8sPR+2xXTWtQ4oSTce6XmObsvrPv4pdfYpaSmv3EfYaQjlBV9gWlOeDG7vyp
OHhDS+qbvwQHN10m0fD9cDxVb/0UA/QybCKUFV9xdGSHp9OKlcc2td+uGOvTF1zI+zYW8zA0Hcds
Y5tuc/MJkL7MhfB/Glutej3UI0X/g6OxCG1oMBbOqFuN7oED+YHnH2VucggppLJUYvAlLlIWdomw
ULCo0R0ojCq00FXiUy2qCrj0qjsc2UcITGb54irLD2h+GPusPsJ3oI0UqHj+jOUnOhAqhrw44xzL
W+pK1+jJtXPkxPqLmHJxDxryfEBbCVq0muqr92IDCRGuQwlz514UeHEo/wyDSfrOWVEwUsjZIcNP
AzU2wCKP7Oobd9S29yI6sblqRI6IIjEc8UJDCgEVPnePP1l8YgOuWk5dh8SAGCXiIFp1MT0EMlrC
x/uRgAAW5XnOWrdSoGAXnwo0tBm246RJ/Jw14NGIXN17W9hWA9W9wjTxMf47e9bhX4kvnp732XVq
x0pNA0gqjelomqTsz8ecn69xkeRAv1bJCyP7qJvf3Q0Vom2dlxnKth4iFUbDZ/jCi91kzLtlIATZ
1OEBViDsRJ2JvlW5/DGmulDv8fUcgdtwYZshCtreDVyFmc/0MHBhk5lsgc9F6t30J0ymxWIsJrkU
IIZrb7R3qhxtGxBg5En5eUBtEVFpPWBtbKxTig19g7BwVUt4XogCJ0ZMGqXcqZV1ExXeq23Dr9c4
kVderm+RsYxbjMx4ZN1eUQb9RY57ns0GFqrhkBrhUKAbBepEbhI04GHifo0FC3jOMx8eINknr66x
vPajBsacq29RW/o/4B/Zn78mbnafL6ldFz4GiaumCnl+8L/H9bg3Jnmhd0qEJSiGbzDqxJnM9V2E
cDSpUrM+N4N2fKqaXm6G5eLKIGp0UZwGV+O1wKM57Gy9UYDIadTsAC0v3xVD3rmVQwV+Pw1ygwPM
ZCW6zUW0rfYnmwQsuftBwv+pQEDo0xjwjkAadh5cjbva9BwLoQ5yLQ1FqTUc6Y0cT2q6u6vZzktF
gNjWxEO+e9xYnzrH+NFYirF/VvTYVOIRq51zDdeMUwmW7+HbE1p01u7SxYFhvcCxIVTMCspGNBcY
7qN3c7qdaJNut/PmBLq5Iwb7bZpGWR8xYn48JU/u8C53rOTldtSUNpt1CVDzLoyU5gkgb6oZNrCl
vRcDO9XhzfPcaz6/vmilT/XpgZZHuBP3e2ZUlORDtcqi4btJWYAFZsBLnnoKv/j0lLGmhLPWlmSl
YiBIN+Epxz38bU8wuJ9YUX/MaYF6lhb2SGQv+a0LHWzFgRqRv7g4xwATTOZR+Qioyyjid6mVCfXk
ERd3Ktzd4y8AuOnu80oGx4P1Edih5KZOLTcw2r++pWjCHdemaehflvm6yUVV36SoM0L7RbOvWLnQ
kTPeNCC+4pMPN+fFZaVtyLbejdLPjV4NGAKOmIu2Ks8UMgE1lliWkQ5Hs9HsDbeMxfjhYP/SQE17
TskZFrHQCeQqdPXjnaFeWsXiY0u8Jnq82Q2LNxQavEbfkQ/tkq02NdtoBFOMlVrQnMl7ou3gYiAz
+bAMTsrjer5Mg6hL7s7rgGO5QIoIBkxa2kFNJQijmuo5Xg86fktgRsIWWFrTGzc2rXUG0VbtL25U
WqwpyKVkumuG1N5iePy3/9TTCs/XePxw3kp6mkpi11JrMBOsllepJjxaTHKLEYSVRgfSeWbk5rah
V6j4geuGkwi14j3BA3PdTyjbsKd3TdJSosCjDtX8Ce+gznPLwvz6rfQZ2i20Ms0cpatvrgMUHdDi
7DVhQHK1iPCMzaxDuJjDdyWzahDq2mYhD9OIb26UG5sksRoUUg/LoP30HOS2ttPylngUq5AO/+Cf
xKQiO7BiEh7N0gFuCeRs2D7PR5X5chfwF7XsLxu0X2ocyaQYFhb9jLGT2oeNbp345teuJWfX6hOj
CuQRnfIuUf/nUkJJtrVj94mcWdddKLkgYuwiJJB6DZI6maLZEg9Grdw5NDWndm/cYQkDGT56wQcX
mPxFN9ZQJXnXAZVeiErI6gtqbYyXh22+ZtPKk/fk3/BQ7LDiyiM4A/5405zGdubATili8+x+/H4W
jgPiXq41eWrtWSufOzhOX2+PqNfNblLoywIBoDV9IAFqis/4zBF9SuZZYIBUe2ltnqj6unrfQaKq
M0DCqWroklGsEZHtj8R4UQm8z/Y5+H0eN4TwEAsEis341nenzaGqlVp/L4WKCWHHzDiZe10TIK7H
9vFYmIiXq3y80MeLkQKafqoh4EGSS406D/N17pUc5cSzuEZUw/0J3pajTFSBAVOlUrb5upZrJkI+
iUV6NXPiMEThTEz2tW3q8642Qp4v/Dqyi2HYCBGj2TaM4IKvMzZ6bpgK+HIORPeRSDVSpxDwa69y
mf7s79AGMYogFLljEs4tB5I0q4FeOZJ2wKiAN11m2bP5yfLrX4Bsa8FevgQ6asdVYlEbT94+LUyy
Nl2YI2hpFE61YeZnDipZ33gwogDxbWpw0U2HrkD9VxNZFT9b/nWbEvAtdWxu0DIIwVA1zPzFrZ3i
arhd+QEJFDDh8yRkkLon0BvOavBTs2atXvxdgTL3YerNtDEuw9X6iAum41BljmycLY6CH+/+WhAi
hU51HzXxgtZ4XEAR+05qO0XQqujxehRJsL7GpJJpZKoqfb5XNd3fXT6bL4Att6/snEAXMduv5l3U
NaIZw7xG+YXToCSb/ZZuJDWSdA+jZXMazdoi/SpVxO97PGSuTe7OzhnLPNcrg88UiOMU+xRRIHn5
N95Bc4rScTPGErf+qxCqlxiKeDAaui3/KihVDOnqeLdyQNzhlqAcdDi+AuOhEJs1tZr0mUypljjE
rfFdc4W2FmZIT+LJbEvStfAFro6hkkP0Sk/BlZOmG6oVoo8/dvwyrGM0+bDcZ25RdWV6JRyoX/qG
zEFXtTRe7rl0CGsnJorvE1sfhKpphTx9CwpI5DWrwyorT1w5aKRc4uQcItJGaWjM9kc+vW92fFN8
NgEDrAHtCGBnKLjSl/0ZpTasxUfHGCFLQILGsgeY2HBNah1e/UpTZNRZxhxiBvtfybIVj99NKH8f
Y6MgNnfpaoSdhLTVADOdTKsGPRTe0x+yd4xL7Exlq6zsC5fEA0ruvNjcx3+K8ImxTWYdoa9OC5gY
O7a7sikKHDGx+wNqhgJ2FVFf5MATwdrIErSKyUl+aHMqSAB0HHEIZ9aTxOk1p4kVDBmnYOrqhWTx
ZZ431EIswm/VG3GGtDItBi9Abb/s9bp+Hhcq6Q073KS8LnYGL7Ec/0xDaHnrmBFx0YVBFcVXmtI5
nTtYHYkej0QhgEk5gTdgIEwHbp9RbYmBibCAwBj6aByW3v5OVM1/JbCN17GaeUwe6zDLTEsLOXhb
MWS82lT/RG+IxEj2J7wRNjAGd9zcJn9g3nnt30id1RNnN9UagK6QcnNDd16IXnghEEciTr8yDFEn
wDB6cafUFKTGoCJseV109hcixlAoIRyNBurIwXdQD3zLd74LIcJm9WjIs5zkRew2vF40RIvldNxK
7upYJNORocESBTQkKIqENVfxTW5HAOeYsytbKBtKFq9GNso0a2ZEopAfozFlEojQcf98QPgmKpKe
0B6rwgEBlGQTgD+HQmtOjusVFMNmmNJBvhWIPv0gBB5Os6dHY6CBrw==
`protect end_protected

