

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dwCKj5yWv0+IePBqJHT08eVU+DwkTeU5oOrKTCm5D5dLE5fjKonyT8s7ehOuYqmaU7hbrj8cK+dG
v6Hkf9vaEw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ofPimz6qWDPfdZmLTvO15AJD3qAYPdAcnxW7u3A5HKCVeJi1plo2JwW0CBkFgjSMPqG4mB4Hkwjh
aser6hfQcfNXvJ3JUWr5ZS6ezr5tSrAVnAOcpabYJ2vlFEce3rPTiHxnx3vwSLvA9frZJO+K8rqA
zTaVjBo7aLNhP54LcX8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xVx1mMvfUwlXTa88EF8IX42tnG0cXSGFt8ROQqT5GxjYzkciIVjF2lg5N/iujDWrU+m+Hq1jVN/S
7L9ZrnRgKz1GFQOxHGVlrNSRcf8Ej88lKuK02N1SzF4b1/VUH6ht92N2p/ROW4dBYnWVBpIxhF08
xg1QHd1cs9lodA6VBrB5Eo1G6aluz2m9EBGHigHdWN9RnmtH4Lso1/y7QElbZq3E4/diAxIYh9aF
1JcFvli+iX9S3ENdEluRyVweVryo5jTYqJabkRWFuo9iOs/Ic616lgSVONZ4NUl4ItIqkTq/gP0J
z13d7iJ5zyP7sku49PKKDfaHMGhWx7ug9eg68A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mm3ysnbGmWPGigjf3cW3nqCJ7td02DMWAwGM3y8Ir0JjWwms2hUSloczYrXXwus0KFJrOvbcp8EI
afa1rxF5AlIKiPd5moyH7qLa6s40f+FTseHQnAhUIfuaGWVSTafXnP1rMlydXotX0OgXaf8ss8Rn
aesy7+qw+4loCzosrzM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
quGvQtw6SKSqCyA6Sp/eeM9Ow8TS12WLAPu5jebLdqM/ryW0A17A8N0thkaJZco15r7Owh4nFU5l
KZcrcDhvn1UKmGv+3eWd84UW4QDpY80dJTTq1XGSt54iFPTL0Mo21C1hbrKXm36H71Xi6xWsaAlk
nLsOCKMEHsujeF1naPb1xFZWSlnfCp9K2SB7wEzz8xUdktOS4rqm8CvHN3HMePG4N3SsN68l6nRq
sed/9GKEvYzA04tbQb5NASiphn6udoZq4W1cZDMS1xzdJ8v00rtDdh9Iinn05spY0CrdzbMqalEN
NkRAqp28PSG9/FiSfEP/QtuVq+XzCkevSe/NZA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 83872)
`protect data_block
L2Y2HpATY4OMNtrGLbk3p/Mvdo6WmNPteJSb4L5PayVCssM0o5DPh0KCHKoOQEB/N8xF9MAuxta2
jQPUcGtk3oewhwDLbYaqTlkmSz9r2ladLtWynK27X9GFWX3iJg0XDfa4LHXAsHywXjzNqhuycja4
fDm5PnEM4u3393nEe8H8miFvyGsNjiGSU7Of3h3xzhaEOtv0f4d+OwSgpqBAicUlQw9oBlP6LE+j
2wKiFrh/q1fquKk6KM7tTmUjELu1Fkg/3CZiKaQLq3h2qhyt3HIgiLrkekCVDP7NCJols4Dg8oD4
cTJ5ohRrKNACpDtfW9x9BgJSHKUhFMfd7Kdl6sPiU0Vp1GqNpy9BbHYgt2v74fAd50veRhoIdNRH
xmxSSMODUEhFPrc//iFZgeASHe+e+MMRXCb833UxSO1i7jmTPqGkQdodZ+GDAx7SPRl68yhTAJoz
VJ9fWDvxqz+fciC1xRzorb/RZa/Ea8UQk2/KmvBXYvbUyl3OPToE4uWCYkp2BZEj7LbfBNeUCNHp
Mp3zA5YJuII6dR3sa2leE2Jk71XdTtRW8J280zWJ2CGtHk9EDzGVTDPeqbD1oKHDO1b9awocESf+
ksfgVGolGEYVTbwy5vy+mSJom/B9H87MKGUZVw6Ks6XQF4+WCETEpuqntkS1v2LjuD8MQgL8WDwN
SKgly6NYxDPs3mqL9sXm36j3+MdIx6GnOEmfuQo24jRAU5em5w7IRp0O9Ok4/9zTsMe9YP8YoEIl
KO5W0b6kh99dtpZJog6slpS1P7ZiabWQCrd49JhYGk7nYPJz2NY1gYVPUnLl8Ke31q7ClNqranc4
n8PkG2S6GqCWMGR7sqlM8zRc9Auw/ZvOUm1s4Tbo/glnFzHZAxlzoXy73oLUkSehu27StloRSkwQ
fCdrPWMHu/3acvF4qQcJ+cWvdnitzU8AdNen4xgIh213Ht71fCB8ibKau1m9lrvndHCv1snGprmE
jmp0rsNovde043Uyb2uppkmd5MHYsuN0znb27cTXjg+h3+Vji/JRdVJCblWrMaMM5H9L3FX6Jzig
8ZRGMhCrcggpLEWWXs4Kz+msbaxUIvvXhDaqQ3CyNJ/AsR8rRV2hi2HRz5y3xFplncjq3Wm9PzQN
sTtbFCFx9CPN450UO4AfWXxuc+O4QeC/mjULHJrmOhfM+t3xnExUBO+flX+zBE+M8tr3+YSn3L8l
i5BcXt5ksjSPoqAbBfNfoO+8DdqxchayL+Ofgkrfg5meTjCag/srrgmLn0ySPJp3BWNmy886ek8c
/iARaJ9FFctpgYipSBiB/tOKP+4pwFgnPWoBqQ8wIqCcXIZPxRQGzcASFj1pAzceTd6uPsNJ4ac8
d2V1q6mTle71Dv3eIL/31cRctZkZYX5KGGwkKpb6WKmUqnc+c9LRI23VsG/aUrmdf89gR4Xv/6TT
1m6/2nCaoG7z5IxcrlIOPxesrpBouppGuuCOAyjD82VSi0RxepzLhEe0LVtQe1Lac+ADsKhYaF29
Vn/077o6drsGE40bS5hWEFIeHCk8Ug2ROliaW9ndtKro0TQCQ2W8Let8qxhHecujMm9Yh1XP19ih
LAKXlOKg8/sW9bnYu73FhbWKxg03e/A5KpWjvwfGxKSqJTlgCzsxDIZ99wXgzue9mYVQZ1zvplV+
h21LL7HQ0aNp4lQmf84gkwO6o77gNzDfKX+78Y4UjoDt29xp3VztceiWIvg5nRAOzX1rcZRtPEeY
JkEK082IGyp4EsyYdrv86A47gQB0DIQqUWReA8ZnGF8oOnmHinQ3QBvJSpM+rZW5ZIHqw7n7zlyT
etCTjqpirJOfht0FkLRHi+f1lV7sUepebcamO3kk2krQ7svT9esQXUseynliQCNAr9JWxv4lxi1Y
z4VxSAOqj2ISBEKDO76+8cs/CvZHNKYsQxLnNfIujzgSdayZjWUYw6HP8h67CZmGj9HAIkMxhn7P
jC0IQ70hQB/OeaWfPqWbddmL9JGHYlc4DuUkd3HYUKFXADrGGaNP5bPcHYHzHPJDGpguzZ6t2T7d
0ql3VZ/hoVGKCzILkjynpz6T2SLFoSxB+YXrWZKjOsigK4giy0eCZLaNSE0B1T8L5vzeVZz0lvPJ
9QqXZA0CAew7BVNdyOUET5b8OpXF4To2JlRYmQdMwGHtTfEVL8QuzuLFBqK4sKMSf9ozqrFRZgA3
p7Vm1pzrO8YU3otZIuWJUQ8J/uZ94r1vYs3fXLvzqghLX6/wnQaJ8aUGxSZkR1P6eQXibJDqK6zb
H88Qtn2ehuZ4i+4NbXGJAwXCoMATqisPOS7UBz5t3LfgABO3E27qKMugj3NWlDN9Kp2Sn7h8Hsqm
HjKOYcN5p3Pd6ROikyamjDXoKH0Iyw4PoRAUBdlaSx4/T5GTZ2yY3CUS6eouOA5W7DqfNqQ9rwvh
kxPCKPDsrMFOeeEDHgzke8+PEmLtUpfZLQ+aoyUhuSWErae11mU+cZp03/cNSbTwliIfoPL1OTIg
frIF1XGHF7hgk633TO72Cmknf7BLlbThE5c0FZllma8yJ0kdrUKmzlqyc4DQBZ9A+1xigrZHcXG3
lu1CmwaX+7Tb3RYQ6IaPSNeRRXGpcNuOw51P3hNf/uP1duvaUtDRSgNleCSGaYS4zvF0CAcQFOLo
C/JxjLKbcSnJVreR4ujD3uxZmvr0l/IAlhCxJVrmPHn+MwKw1yNwTDnh1GIhhKxTivlnrj1jlzFy
XW1rO923SO+gwaJYgqWMSa4DLIcPJYxr1MHzdHkG2aWRHt9bbNk/k0EYOKHokbS1JPme3V9HIPGk
TvlB0RJnDzYzgxYLfMlMlCAg7zcU5aIsDpRiB0lHeRawIAQKkzanIMIdwGeWvrut00F9FBqQ4P63
kUq1TKDyQbWNvRS3hKCLG6MPZ1rPIzTypl0zjyjVJc8WSeceJF6Dz3RLf4pcnoLMLa8sW+EU+2vb
5VUjYO9c2C1tm/XUgx5byR9WDT0aky8PzCWswj7qGZxwpL96H2oJp017XAG46TNf34i7L4fA+zHN
01xGWg+I7QgDdYJC6qVpG+ZzhFF5V9eUBZSTLcSaIvpxQO4tSvRfPhrYfNXlt7IyS2/bMQxsysgV
NxlbszIZlqCC/hCBNSl+XpM45m3ZmkU5BqSLSgrNfW/gy7pugnM3Bqi985V/OmJw07roC4/078F8
WLH4qkl35OlwRiBJDSirMkIqU1RN4jSym1qqpfoGPWl/mwQ1wMZR9utGUz7+sSYl3Kc0LGP/6FGV
aUFvFR5sEH48pAvf50IPf0xm1eNA37yjF6K/h4U4xwauwN0faIMkcgeYzmifONcYnO7BxBKmsLH3
RqHHydZSsB51U6kDIiRzQBpk36gOnS/tqaJN8e+57woM3L7YXeWBSmDv/4ykdcMIKNcnYMTO5Wp3
BTuBiZ6/UyDQz6wKTO4f7oT0jIk1J8EQFiPiEPyLF5UYyyH+3PwKnCQjZwx9tihkBcWqI2DRF4H0
lt06tQeVH5Ti4a4lw6o/DfFDXWVE2ShtOmP01zPOcxNphfM+AsSksGq9cznHR/OEnig5KlrFNEPL
6QlNv+hsMv6dhyMeAqZT4B6wf5JVPKvVw+xqwMZz/MGLdkPisrZX2/sJ/lXVrplhLc7X435D9Tb1
gLQ3Sccz6IlBhiGQT6VHH06xQBp7cH3BaOiDG7WQIkXIAboDIbkdWWg05mOYrT9/++yVZJnr9lJp
CtLx6iIm9uF8JiL2fCve1NAlgLbQpXEheP+NiUDXZhPVIZvCIRUrFuh80ZYKkOdQWiPZrUPOsimF
OK1zR6M8C2V+Rb87LqGa61gGu6WX5cBH/723c0veTOfC3V4Cix9j6cx2u79CLWe6GBJcC2bV80wB
yB5gjyRi8+RZ5VVRJwpQOYF79VUYy5CeUssScs30DuN055ImYENz1SKJyh1iPjPItl+TzljN3bxL
rWxGWDG5GFvH7JjYRJuExhEUkmAaJozpw3YKgrO5fkeh7XWuOIdK9GipwUCrFk+BvqexdoyvJeS5
WDtDk+xTNaN1LmWJ6DpnxwDu5GtVGxPcFrOVVki2zDJ2n0OryM8ChKupFWkYdzvrBueyQLfYEx4C
X/I3Qw4uUa1fjuwlzaxPwaF3ssGGesWAwIxheqbE9Aj2urvtjmRc0TkyAA1FkAdoOtnr1TBrRk+X
usiEWxQykJ57P1PAUR6QHQl6/1S+LmA+n5tBLyyMnLQcHTEWVlqj+isR1+jOw7kOYu8bGZ+r0nE5
nH8ACaVrx1WUqzwbgcg+Ao9Zrr76OmtzNsVrANunBcZpwnnfMb1PndfEXU5a+zXLZpgIHEaEdVrA
RA/kClOMtimR8ZLNB3mlxZBQ7mY46H5o2MqStwrqss7qijDxeE69brfstAwYNIceIkJMgAIqhlEM
8gJ+tv2aVPbdFwHFZxOiz7mFFyd5YWx8t3Ofaz1LMxCHbXVuISn490cgj6SO+eE46hhhr+ALSgLi
P2axslUsw2dzMyvvhAmmUKxvHWreH6vLHJaywcFyJXBgHW94FA02nCe2RuRiteviSFsL1zzNOXdY
ZM5LbrAE2NzFI7k6uMG/AI2UW0M8RFuZ8kkwFVrEylT3/9YCJfEmG3aad+aStUKzq6OqIf10WY3Y
Jrikguj34KZj6+ZLh/rM1V/s4u90Se74E6fIipSbs14wPwnvWXDpch0cI7BXEP3FOigIOB8OmDo0
O/HikP6SLQgAsS8jmXG/M5q+pggAlyJidM0qZ8tybVbje5KtUUH2eM4N+/f2hkrg8uvk7FtjHYfo
JrfLksvwZyAoUOEtFeB5thQMVZBEA/DzMLiY8fnQR98OVc9/DsxYWJ6PRZM87XVObT7wEs+lW1rn
61pmjDzyzMrw2NV0j25pJR+pk8fFEM7YAdAZXcP7Mp16tZJfzaSdZAbxaO8h8QXrKJ0mrZiV7nYi
oi/57An++Sy2b098WagOOJSlHthO56TrhYo+j0SVyn19zG9PHS5ZKuSWKz/mbundyvTK2p09CHJX
lnf2Q4MGLuc2j6Yql5uA6xpSZk2mBAKHpYHcwuUqz35xZIgiXATe1fma0XCNCCPolkn3YMHRf9gW
bHLStyXl1ojAiXjv8Ilq/Ik0szaZm7XJUA9emsL7hjBWfE3N+Z0ZC8hZuoJLwMp1d9rH/zPEwqc1
lggSJcxJxP1vV0vV0vHKqb8paBF0PtYBW7CCBfo8R71IxwPcUD9pvXPPdwcoAVr1ugCYh6W6DqLd
ndQqXbJ4UC+IvMpkDKJWsNqEYmnKNT/0DzQKd1fYbDBsUrYtmUy9rBowRBGCxSKD92Ue3bIW6ZPv
lzTQYVfQHkRn+G36u2spLqlyHqzus0nTCsU3AaCkeeVOg069jblQK32B2/jyOmvzf5r27o94cN8y
Eq+zncwcpS/U96+nTYsrCpSPf1dn6gti68tGku1Bk4BzzpU1B7plwZRfIQpNoBJdiLY4hUDHzTFK
eBjOxZY566h645WuXpI6VRbQwamcH4ygwn8OI3G924iAU8bt+lVzXubeBK2uGSWmul1e82ilkQQZ
T9P483ycmRVKxHXsXx8tCUVWjZ/clOBqSHLlShSP2CWDrqGROx7bfeIdUF+dNj3SW1moKyaq10G8
+N4XweJTDTyLRqWgEgVKOMH0mFvl9ATaCz9nh3HFN8YmXQ6X5ytJTP6HJ31fLvRwT8oY1gdGw4OU
s66fJ+KfhpEbmuGvAfH0c6NxM+gW8sgM0jRDlsswK1Q2xhbpbxpTSvPeF26e9rCY1S0/G7/rgTRA
q0loD7x3I8Ppej8ItaH/FbDsZgmF/SyQnbm/teqR5x/OHBPvHkf0q/wdtnuHDY8bjDm+WDFiNaE/
W681l9Tg6D94dXXaPoT4/7MYHFiAhWCSjTaLWfnZQRJCVaAbrEfBHb0o9pG3ivnmDY1KyGxww4rF
j++jthws5OJpB+vjMp9ZeYKfX66L2K+Bxn6VT90D9h+AtxbpmslVRQDBEirpicz2ntYM6pDA7mTE
nopNLxnJ5DOPtqI/9w0I0XQXsq8nYJkrJVCHjla21PudAr94VeLYo27O7FS+T3J4Ky+VcgIcb2yR
H1tiWqkjNvtTjMLgMnLaLerNopXLdLhSIdo9XGWN7BJPCuu0IS1KRQNFbeU40KMKfhA8jzcGCv/p
Z8yqW45BYL9EzCrs7PIkxj0GHsHex7gbaZzhUt6It5+zodj89RlQVLQFvKpyxHt3czqPc/6aFrQB
KsghEAtFGGb2rjzAa2jEe/a/m3DXomxyFGd5fVUj6qOpX0mE1uMCjkGK9TlInsrLVHjOQ3j/eg+x
qZDFrQrKaYq9MtK+w+WkfkUcg2Oc0ryyt7ydUP37MuqufrdHQoITb0KkOE8ldIatoMoyAAKgm4Oj
gJ7ZZ+2MgVpnWH269J8ywfkbwVwy1S8asGE1cpQLy2d9xKNcSn2dbNZ1PccLhLNKsEz1tROxWTkO
XLWpz7r7CmNUEsX3qAlcyt+OgDfJDVpI2HFpGkA21oK1vYBHHig+1IWCKCd1lPBEqTrgibs+sVkb
2n5HtS9gje+BrIEmsZHsAgzypvzcdWtN0WOGqrknI39qUu1qgGlIVMGNHZ754oqWXdFdIY3+u6OP
Foycuq0bZhNp5V9FV9qkHJwVSTl83x/puMzmjx6N63SmKJBmB6d7yU3V8Wumf5TaY6fz4Hm1oOVv
lEBMDMkRqyocrRduWTEsMvE1NfEqKaXpdGP7htdg9dYiCl8P3E9JtxagOE5wnNfSTVDGwI/PC1OP
95+Ww6oorm0kDWuuABDH9Z9qdz7pq4gBg9ByXnrsZiEcUtNyi+1X6jVWzA+HaMTYaTX7erERCYHp
L9ezjpnTJuzbro9GZAR1iFkOExzH5mMD4Jpy3PEqEuS2KwjtxXKpHAGrhyEpjEX7MwitFpqO3Tpt
duj7ADH80eQT7jybLSaQgW4rzB6mLWuBdZfDzlA7zoCExpcqyWrX4jrsabF2AGht1IDVSUbqMaqB
LLLM4XEEj04BKWx5YNPQ5k3oJgsWW/6KuNQt8k7digtWQq+e5i5YVhZw9/2ePHrACt1vPhNFQ6Al
Sg993VsxPyg/wI/ZsbW6z/FcLxxYHvFRDUW/C6uiFogWGxhwLYvuUyO++uc/fvXWShNRAdwSp2Di
QVyFR96CELy+sBXeHhY/q7lAJWAYOWuF4/NgTM5bI8i9861OtIvIrzjxSkLK+wqZndb5iziExCtx
Z8cgPVCMVypIu4J40PaeGnq4tz5mXMJ6LlLMKfszWExzgynz6bHDiN0qhphwsfTzeC4n8A8dDtYq
6Uh8jpnyiPSoxrtgCvnNGS6CJQT7Z5QzD3vmxdbmglIgBm1k9uc03et+PEU3AgghzWVmGT4zEG7x
ilex65X8RtNvWE1sbredj5dWpv5tqDnq3YLshm1xbwEVCrr+mf9OfHAQUa4/8nanemiLAUD61nM2
rjpxXqGrlXOe4D3KtIkakVczwAH16EJCkyN4H79mU2GjCCVgl+0WLrfRSo7WFqZEAGkaBsbgs0yK
9EPbHpEmAUIXmQjdXD2sqAfCWZbcyub2XS8XYp5kKRC5svKWwUPCO2dQoVTn0er99CrFmebfzR6u
c0ef0nMOqow9VdoqnlJdwIiwg9GRGxmueM2K/OozSuFTG2FtQs6qW85YWFOX8aTjRBEq/e91vfTy
mDsinqbh7p5oXWUXEbP6MOI4oQ36FO/ZHTZ5DPHJOMiVKUA7Aj8D2P1a0jCzK4TXORtOAOqHfbAu
rdlGuz5nMnC6SsHEce8N8ePbO1ITyvGjN3WWYk3JSnXVgsRRsdcCppTQfplvmQCIGTysecZzt+oX
uwlGjmNKT6wRHCVjSvEp+AbW5g9w4Mo43i32dnyqLXSzBs84866sTil5WM2DL+JbzCXvYQytLEiK
AizOsCN+vliSjG5ygvyJQZvGt5M/WdUBFXhFAt9UNXLkVnUPFi6F7IopYo+9rbfETF6xf7QOsq2d
LlYADH/OsBdpelq8gHa7DKra/0S4ev9YjLFynlit8wcOPwYqP6+Z6DZtBrFWXo0rkbVOyWZQkU7N
C1/7yfQ8kxxtQjhpwh3zv+e1XffG4jhuWhu+wIaCA8xxWxTrBvqZg4U9RpE5c5CJAShaL+8e4gtz
nmoQSogAKafq1Rq55HITdQoJTnhZAgH2UP5N9FRchgOU1q++DofTr1G/MTbmC07JVHOwr/hPDHZx
OFd7ievbswnCOQ9J2MU3J/oMX6ZHZ5op6fj6v2R++omQlwPNp0uSySEG3WaV8AZTbYvStlWJRwUg
ECUFyi7/9kBI4ANvtNBcGm74djYkjWk3jxIn2EbuACckZVns5xmNLv0Ak6Mh8I18EVrGKHMlkZ92
hMy3e4UaeTAd/fIR2+oe7jAWQ8CTiotTeIyz2F45FZnO2NRsnEJ1mMFE+B6bVNMdHqP1y+RET93q
3n981HZRMCOFOmWP1NboOgY9BfJHTl1/vOvV5Ul1bgG1DJQaha4JEwPGhloDBFkm/Bc+620u3rC/
vC5738rhrk1ZvBu5tcVgSjH8D2+KstnwVGlDXgl81iqQ1QKAX7/69ui3f81GQyAaCQd6JvPLoyBW
iVZyvHYWWWTRKNIktcov4PYaXwsnV72gADs4qqEAHFc6Ky1QaohZ0gCQ/O/GO4buCFbZUV/Jp+WC
7B2CzvA94sTsHwvBtZ3ekUab3+PqwmWn7l+EwY2zFeOBd66/RKyghW//gHyhkxRPaeOW7EVGKVeE
7UnFteCJfy6ZWKK0BFl/1Sb92cDA9crw+uUCr+Nex2vef50vccftPz3VresTI6HsSpCRZyK9wNcp
/nSm4/kXN6oHCDq5Ikj+pMHY44T4gbbTN+9X4mveldpz1yKrowavgcxoPB0/LYM6hL1YGSMwnJO7
7dk8p+aO5JxQj+1Fe1RHD8pZSTBbi2jdbql7vIoPHdp/GMLpp6sE9nfLeSrS5XPvDR5OBNTAEaa2
PDRn8lQSAPlUv/nz8ro/tU3CIz+l2qTZXSdiSzcq+z7eYzJiTIgYef70IRhAa9RmvIGbkXGGFHk3
I8whgfN3SWOz1e8IKze9Mub5yIpEtnT54Vp5inTkYWFdtVndbWc6sHQOjoU7w9Anu94yF9a0aNJK
s68U/v8r7Hz4TupK4/VMD48XL8/jDbkSHWx+E9BmJ9LQxGeNFCJGUkpObDScwZjar3AZcMnQUZza
Yu9+ZXzBqYu3YF7O+CT2fA/d3wvk3Kn5BWDdrkNTe/AqxummWxZ6hxqWNmaqoLWSFhoprqpusURd
z++5Bo1RejZBROORQXSQ39i9uu57oTK/lnz0s+LtCevZxH3aN9nG8g/CG4UxrhCe+hXIjEiyPf4Y
BWR9JzR4MpXcmME8UmtHBQ8VlbLrWK+/pYtsdcpvLIlpxCQt8RlEIJX6IpY/+Auwctq/jXEmbY8h
65zQcxgP43Q+jHnr7d59cxtsqyxotGACZY/j9NRjI6m6zVPD7mlUZ36kLrprmbubt5f0HtnO26Sw
BWD+Z6pt1psOTwj0EltMP4/SCDobOI8uTVF2vfrkhD9Vfe/Nnp8/qFqNe0K224f3t5wb4UXJGzXQ
5zHWntmoHpiZ+3C0OyK/w1X4eCjEvODAjklj5TJgrttY2lJKZrWyF+SExbxbeQjl/RPTQDpXxHyI
MTb2TCquN2qoI/CI2zVPf4grBt4GbHzXJAiJm6dcixCjV4QPu1tGIb2ajwgFGi+UXNYlmZHvz7fB
TLQBopki0PZavaHJUPiaixT1kahFiC+beAxcNWvBT1ktZwugwjkJeIKbDrZRx0ku5iKlubDD7Hem
wVeOwaHwUkOznGe6qDLwNpUHCLsFB8lg+O+Uz6gno9IKiQlQ3yO0VlkOmQvB6T8mIuf9ceddCXij
YpJSebcR1TSpIyhb4pZhYJ7dZ4ZBIdmw6g3K/Mf13Y9q+A2wHt8L8BNIAzIHIboGiwJsGoQRXiSL
P9VFf74PEyDO/ZQelVQBr0KDSdUp/2SZRW48S+mj1PbtPda2e7vvU0UmEWPKq83g2rR4uyxbawzZ
EHxmZ8Uz9vA1AOujcCfbPqbqcTGeatRktKjb0MLSmVmtT7Dtn8Wo8T8anuJcoNyjr3r6XBTh3UTJ
tj1gvcmoyIbv/Gp40ON5KinOborYGo3mg8wBhpIofwnFQy0bC75RSyg1iLVXtiSv1FkFbJJqQpZv
J7iFBpaRU0RMC2i524MJrXmd37mQd19nRCnICLi/CSTaK4aKHJj+nU1ylLudbpaIKoUhQRFmzWss
73Mu4sH3Kivtivxx5C7xJesAp9g/85gQ8PeccOmBalPwzMuFNW5zZDqLKcGZ4PuaC/sXz5Kvuu28
nzQFEHA3x3uKQd9TRG1vYcHWBACEP0Z2wVSfx9iQLGz1O/6tMy5zJf8idjNjYv2g14DJyFzSf277
ao3IUT4f86KJURnaJaVwoDyQEEZWFmaQ1fhvW1Aadz86hOnJa6cgx0rWrm8cL+R4GuqAQCTshSVn
HTSKJPxzLwEKMrSKchxt045q0SP0gjgkx3WiLPqZRNF9wJ6y3GNc00c+cmlel7xztU+lTarvSB0Q
6/tgVb9laW6rWFRNJvZqD3TpnRbpoXI3iBBPNGRRbgZiupgfSX34J7wHRONCxw210djeCbyVQuIi
44QJm3qDWBn6ZcVS8njHDSfrR5hkRVJDs9F78WgrJfStQUn6wzvFFkvbN+Q8Zwa/dMZc3oEe3B9h
K6D7we5M8sHhieapd7a8TJxqkxGS5nK0IJnKxwhncSHGasHk5rwwH38SynL/9dX5depoEiBeDV2y
IpntFE6uuQGTLcJfhl2x20VK7fPTJgozPcaevgi8H779FmNM9ncjOf4g65RTzY3iv18eZU97cG2U
jfZ1D4zyUDopB54wB5frFhV1LL5Ul10Pb7AIELsB2MkSrqZtT4y/Q++FEo9oGEXoT4fD3LO5gtn7
Eh8NfDMFu0CVhYJIzEx21baEyFkbkvVP3CSPuJlbtxDU2c+uuq/ZuZ9210QcFZAOfACn+QfLBsSe
BAVT8wPeWE0Rjudk+5LyayBUKn51OhvSbQIcHOcFOgwxpG1QoVEoY2X6UAz5XOXYzAztzgMZUn0D
9P1Pnm2uGJsYk57ZpqW0+wLflWcK9aFqra5ghVf5WUKf/vt6Nvb62Uf5WlO0u1Kfifxb+/9fDRE/
pQ3N6RRUS+pNXUxesx4YY4lBpcdLL5+cjtVLOETCAtyV/ngK46YDRhdBOeMFQBQqWB0FP/UGtvif
wseysU6yVJg9IkAw/UX6e6BMdXKPDfjHpMOSCssc509J7BbRdtNrmcf5KluXrH+hJI6qxOz9tfPt
TW4kBAxtXxx0g0iLCFAOrpf4mWKDdLgWTg7B0KzLKwvxA1UsNRVqtWr+863lnCiZe45318zh8IUf
OoNXK+tQapItQEior5HWRxTGwzwDnJsLeLmFPgC2H/tgUeeixjo5zFjC52ZpT7YNmQKdc85x5DQM
EQweAMxsDkBHqdlnUKNIZgZl5ZncZ7fYV3rR1msz4axWt4p66X3+mY541hRJiG11dVJU54qeKh7i
GDAWI5vTey5OhNrIaud3Sr/875Syn175B4DPUwGZbN2KcSda25eZKOaTDrvhAR7XqyUZs69aqqZ7
Ukkk+2quFNp8Hw3l2TwivONztWkObBqABTQCxGgVV7TiGdodOT0DnuT4KSgTvinZOIWCGEfTWcsn
3n3Gw9sonVUT6zK6A2uhMGpYpigTYdHFh+V3FrRnRlSGUA6ZGT/09v52ZfiwBrgOxY8+UC3tD6oH
JV4hnXJleUVP4qbgUYtFkykVxNiqHj1iXB3GtD3kjQol4cmkJwBgneGUZyWZkNyl0ykNb2o0mW7r
5EM1Grqx0TIqNr4zPZFfa2Hj+wG7LxpC/vKdAp9rm3LLBxoxIVPEuKRvktqkY5uLEufPBkW0y3cL
0XvYfBQM4L6AKBuMFTzqTgdiK33enNbJHGikGdyZMKqHNJiqqZdNQeipxDNBU7p9HcnkSxHO15mm
Lvep3BLijSiWgxQp1CdTNwP4PVnqOxTgcSRiKCYCMssSZkQd0gG9XewBnoY+nzrHQXK5TeWvagnU
lx5sevPSf+LRZYWnUte5saMOf1NwbaIsl9L7118Dxu0vtKN5dfp2ikPTlY4YZj0SNfP87SsZ6ciX
FjWhfvffCVrtNaEFWn6IthAH7eASFwhd9/LgED4wOrLRxpAjoB8ssPqn+E0FNT+gdIKQEvK8O+aX
Jiakfnt/O6c1LxrkgVn3Y7KCsMKLOpTHxINYq3mpnVsF/02Zp4SjGYdUL8lWtXTq4HKUVvzml370
QoC9vQi1JK7mDBG1YfeF3LGn90ns0dPlgPaplShWomxUb+N4vxzsn17MXTtGPNLPwuckvh5Exqkh
5pWQlJGAhR7XkbufoY/WGniiqzb3Y1lNsBtmctJ2Ph2zepfq97t15Pq145/XPxMN9fudThKAiwHx
cQi7ACxnP0paa0jD/apenhZUiUHqL4VjeAM7nRpaRat1syFWGK1sCG1HEtP/tYu32XlqV7bqnokm
UOlLQne/XVbAS1srkiv9/+oGTL+ha7pQZKlCrmshTaY3HtLEvaeAG7DWYLy0jptIbGSfRzQMtWVx
1p+4fplsyTNQbHfjJDfj7tBxdTvX3SacJ0joUKUeI+nFrNY9xO6CTfkH7QCMR3iIOnGMNp0i7yU0
/bR4TePBDa30WRub0Kdb4zuyZ2HEeL/ldOR8pSUD4m3uF2jVQV3DkwnVTyh84zGur8Rm8lU9xBCD
aoGbu1/beK5iBuYKycNH7XMNyp9XNpZoGra8clfsuHTHoxF/x0BeZvGQNAgGNG9GwCVXYg2vbj++
T+nK5SZnEfZ8fGxw1oi9dF73YHeAgYbTPUwb9tcb9+PXibhiwdwj3qe95Zb7k1/iWRt5hSU5froZ
2WzT8xK0u74vrRPFap0DNGQWWyFUFK+w+z4vuJ7/KQRxwwoUvmwDABSWm/DH+xiYgOoIpkfbPubD
o3KDRCsYYTE3DR4BcOKpLY8MglqgHa15iQShqHxg3Zw8NAXGrbSyzwxxQlIAjH/4ctXkgdUqnlwE
HbYi6KoHTuURtRojnlSxIE0q2BXtZmxKRa9aNkAtoq/idWbsg48ZzdSb0LhGM4mSBU6x/mDFxWZ4
JE3tbW/pkZjP6RFU11YUFr5J+3AVjKr3QH6QsROhvu5vwZ6lbOPJ6JCb1FdFij3RIwvfBsXHTNbM
xR1ZJiJ16y7mzLllUMFbj9KyzL2l+GUFbduEDM9gqkgxikp36KiNJyYE18GR9CdASnqenlDgCusx
hPFHaDZ6WlDJF4uLGQGhfJ4P94Rx2wHby1rMNVML9nMNU16SJJtob32N00q2MxDUDtqiqfqvJ+ZF
fErTPt9erHoFoJBFzW2VyODmU4kwa0NhtZAH76xP74RT8IGdJGnv5MoHHdgbsajIcYkyxM/zw394
6UbDp9uWNwd+vV6VBk+0OMjtbtghPak6QW0huhMKIeChbXsjxM7q37C8cjEPJI02HrlOJRpgswz0
epzzJxuAssHGVmlt+sN9F4/cV/q530oWb07Fp2DqHCUQlhElPoOalbxFbaIDunhoKAw4qSYhwOeW
bV3zQPiQ1QTsbyGURwNvMQooYfqJt6CwzQIoVo4T90Gze7cfiw7jx1vvop9/9VE+iLpUOAdJI+Kj
RrY2EaPw1MOyPmg0FXygO8BhB9tVdrp2h4esA5YGo4CX5O3xpjC9Y3V6Kyn5n4dC7xh5w2NozCvB
7iRzAsEGMEtrk/fT1qR4HlU/97N5I6iC8zwElVHc4/8N+5kln2xP3v+g/ne/xTbQhMy/KoBUwP6A
H1rcIdB+Ty+4zuCBk4/nWEYWfy2W7edWKMNJOdMfQhxJqx6e4OvJQRnsgc11e9AvfK3rNUWjzF6r
TgnVpFuStOyGxR/pr9khOy9qOWbSJVVeLcWPSDSlaQm6djj8kImqe93nwnEM3tTzH+mHFn94EDdc
i7qyF8qfD7gCae2Xg1oUlR+fO2mFG6i7p+v9iME8AI508R5CTLXcGEYr/wtu0d9r4qqZ8qSeBMnt
nLi+Ka+gGsucWSar6O4l4KOyhXGf9juBHgBOtIxYqM0aOur17xcqGiwk6H0/W2hgUMOzbkWdmap6
UCHHMKKcX9KOhAWPpt04ZzvVG4nlzRdka1DniI32MYObsjsZyiApMD6WjlATKCxTlmtqXQKPmLta
gbnydsZyfwacSdP8rvUsK1OzTem4CyErF9QCByL9I5dO3huOt6NHC2oNvOqHwV5ptDyoNm4NkcjC
F6bE0TMr48IJPiClJtlBJVR8EAzofVK6GRBstl8nnTjoJW+R6sl/b05QA+LmflMtS/5kDgae5Dmu
Usd98/lFFYGlGd6OHD4sLNfr6Z8288rKP5y2pTl+sQOqaRVGT7kHTo4MRuk3AYDswTD6Tt5s6jns
dY0xTiHIuNk016WkaYxuY0AyKQEISWkuHUP0QP7F/cCQP0nYqaIcyWQqkNHXYaAyZqDrVjuQksf+
qGswNbxMLYyyTCzkllWrPziqkrGIY4OvowbcxXvztD74MucClAF3j8UMv66gsNlM+Wn5LW97M/ZN
eVtU24w1ifmRLKqMmbabmmgWa+g9VB785fmi8q9/fEffl6mmBtJcPv0RnTyo8Tl+JNnnXoYMHtpn
FToUX/UYZPLQ+qEoFfUP1+yuYMOQdXejKQTNDurlc+0L1ykFxF6DgH02NriEduMZTXNLf4eK5/N5
jW5D5iB0STIQfr0t3SZ93G5CPdekHHEbvzlSWLH/7McPewNWLYuqqdh0nNPNcWChJ8S31ba0vgQg
C5uq7VOZyu1fSFtkzwtoMBP+SfdnHKbZwSatX/dqsMAO9WppktPVqmuAjV1xYQr62FhScA6X1IMr
jTErgelWbsT3ETIX8hPxA1Q6MNwlRmwRK6kGffhu+2boy6cXhg9MNaxsWDeAgXTuBFxCZgpGg9Z5
OxVSCkHtjSS7iwLnJqRjBRlPVzSGm+B1EZlHUHqfWPN9MjvtKKVo4mKtORRVn0xi1lQnu81/6tbT
q3Vjk7EfZTDy5E1UvjuSs7UXW+ffYdwebkc2wl8SQKjptZMskgWhvKzw72y5Fg9Rym1+xrwebz5S
U4VWL8UrYi10dKaPUZQc+5E0rzFdPqBny57i+Ii1/LPH5rN4wc3k3Tw3fmXrtODVZCNfA6ksDmo2
zGrN4NdTn5lOOqUi8wxNVOZybE8FA9NwUzd2aZUfInbRI7IoRtlVTXnx4YoDrbVc/HFUmSmz/6DX
DWR/Vs8wy01MyiFrBz/8nD0e6KTxLl3V0T2jh0MEXrRJYdwmVXynkiZDZI8ZnIgoAZ1cJjwLe4HJ
qDLzgsRDFzYQqckvWzZZgLc48ncjF11rxN+P3d27492+Yx5241MC1jVc5J98yvWRWUZPj55u8Pi/
o8vJL7S7YZ3tqqXkbFrswbkzspPURgCWlZYPKCheBKzfvUdlgTho3J8Tipv0nNABIIncXxDJg0+b
WaX/JIKhS4ytoXgLtjTc51nxjuB7c9IiVVG8Exap7pxE1F/wrTDHPG8Iu/ENxidR/HvCcnoKwD/f
rDEjWxe+0AmGYHA/uLOrPsEKyC3xwKOvlkxB81qgrbGgy4ywBAGmjQn0SpBxhqeMo6dp+JjlHjCs
3nLk8EQvSoGH0eJF5BnbL5j0qp/7LsVhK1oc8bGCKKfxe0EL1YclkUrmcUGg4C7kfTNhWYils9vu
QTb/KSchReQjpPMGP8ZZdhCnfOh7qo+Q3j/RssGNoPPAH8ASszevNFunh6Xu2J3s4JOQFdITdYyE
mtKR2GevLrXPf253gcY4prqLks2jb0KoYZoDizKcuRLeu8DKrOms5tb1TS0m4bGHFu43jTLE6+RY
2wZPFPHOS7CIswZNzCzr0LTC7j8dIoXVGffMRwc4fhrG39A4PQGz7CNX3TMSUjOOaJjiHXBOMKr7
ti12qrcFsyILpBG92HPjurXrengF2t5cnm94JlGJVcx1IVkQb3+osxXb2TQ4A3mMHhZE0ZC5XkBm
VpQdilfMsaFHeruY9fgC6it83Scxk7AvWK6u5rzYSEM0QPriDC+DyqOf8zbThaIRLbw5SX2UOiyE
B4sdBEvyJAQHh+SJ22GmnHh+8vgLiY5VzeA0IJWmjRmmRHERa6FRi2AZcd/vfRwC7RbUFGbOHZm5
iTm+ZUpiK0yxhi3CsQQnbjdYLHRecxUzXOPiksJtyy0yeOnR5erh7PKQK06tPGA/lbkPE4MKYTaE
08P7ihlFp6gS245Era106YfN8aEOd6BmgfIp0Igdpdy/E32IbbxTKskz/JysEVFPam2IpSIivjMf
EClvwqqqXHefOv90+bwyDHc3kP+uNlTuSKQprRvvggcT1QD+XMDCTfNiOVDgSG4Kz/YrkBufkkRA
Vm0ZfFe6Y/2sWA18RIKLJZ5O5UyjOltdv9qz0PYOibVkbLLA9HN/T6a219ehY79YOcIHh4P3NYtL
smFJmsk94Q3ldvdV0s+N+Rk7zRf4qJBWAUFc1mGDIJYAmjIB5gv+57PSidwXDta7y8xwFKJInhnW
5hlOzOBRs9L6Vb33e4ELSbQmEiG0/WDYyBxFADN5TsVkiLdtZ3r20Gji70P5XI1Hk/QiDH2hGAvW
eOH46A2KreD77ntNATqF0HOxb17jBhghWKLFjoIZEh3EB9GIdTSt8kFXV+fFPmyg8aK1L4+w79pR
cxh4ghSlL0MlyzJyv8NArHIgvgu9QU+z0/AK9NUzuEUxmqkB5e0cj87T6Fj1tldAlMxdI38Ds6eT
iPGhewP2OdL0bZJ239oEmalbUKycjOo4lVu947zA+F012VuZRLOCfRwCc+mxA9u/PyYECxP/chzH
+1Pu+01ElVr1FUuHdPthTb3UB+IFV8qV8qOXIQ3PNCYxY9K7snYDZvgMt8YpGqsH9wfFdOSgfof6
pqvrOXPink9K2PMIKKU6Qn1zGdfei5X9mclvHUQ+8Nvb6nFyrXvUfDZ9e79QHo5pvAWB4v6Arh+s
iZk4AJZeZd3tJo8hQL/PzOb8SJ1JopK2kbN896lhM38/pLH3dcV2nqg5Tjlse/1FsEb/lURaiN2C
tc2OSlWYRlWmVkG4t9/lC/t6lHWICX3yseJRd083jvsmVOmUvODK4ZfTLaDSBnVX1tz0NfUHyKMW
3ZKnURdu2CVI6tn+6ne3iTALYULaCNBCxZ/Yr/BfmW08dssl0PPm9u4l8MGqaCsW0rQYtdK2IDM7
Yc5XeYJ6NsqW5lae9VhmMmZcAybE7SDSCAew0ZxQIqjqF266zaERFAK1zdAK6DTejHSJQJD39rHO
PyKGA5IgbNxDSAEgSqWFIPrfzjt7D0C6jwRr6DyUOgFlBTjTah6O4vYnTuSqhHOcdz+PodfTxBY1
D+JtJKGHRp9aHjH2dj0gD/o3Hio7alnHTdkT/Ruj9V1a6T2LJ3eCbO03Jp6Ys5ByHQwgMp2T40RO
3zsDype82tuBS9T12ceaj92I90URmPcTKWM/afHlZ82fm1TXQkRNDCAEukHfs0GSPxWYBREHEX+K
tCpa5DZx0OswkJFPMY+nOahK1+ekkoh3EtTlmIu6A56XauAv3UqYQjATE2n0h5p0JIv0LTadjvvZ
NAjShoCIYQ66E8IG4Lag8Q9192rypjEB/zUvX397Bp4bpdacR5Rj2V5rNbZ+aB3Tc4dDTEuKCfbY
9XUzo+NAIlzE02VySl2ZM87oG0KTodEUr4Fbj4lqwBzDvnRNLOD5tCUFcGC1BM0xkzdsV8UvLtU0
rpmhVVXY656a8U/4oPWLGMY1WF0NkGXeN9kq2jlv0mME+fC1WfBP+MKPKBjNTGapb6WsiFylMlW5
df8jyxdsO1wBzG/YRQFXjLqQBcAY+MKwoTMJDPFqrBxOIx4anr/Kzh+Kj9Hazn/ifGhIH6uAuZEe
TjD9whp4cuxtmAmOwrDebal1XrtczHg2dTzRqWy72EDGkP/z5Du3Qmj42Xr6AVjV+yjlH2BgdQym
55l9PuzLpA8FuPdezpZSjlM9P8u1oJf9qcLEEIxf/d0Q5xQnJnjJnTLmqzkktIRNEqijlw4/uOsd
6sg+CE1/DVO4rnsMzcJgJeHFbPGbgMTH/iGFIp7ODLvVOhK8ValD+AiVnVUg8AhjYU7PsbqGCxZx
OqK5eBqAGa47stbqVfS11oLzMboqTBOiApxuJcw+dWeNcAVeFLt4yYIUYgSyx44a26dyDMFoRHDP
IYrfsG50v/BXNOci7QwXYxeo4Sgo8WypPTQ9Rm9xfDvkXytQNDhVdvxct/iU7SIv6oDU9fJVb+Sc
mlPfmB8cNHZ5xKv/B311QRJ/HRfQunncdxkc4vyjrj7s0cHoeSi0TVJWgrvegqb9pwNIqs3qV5UX
9jwvpfs37Y90gkyYJ03HBv73+cYgCi26/2qykiW2FnsmaJrd1AuPx3C+8vaFBjXKdhENxrjNYYpe
9uRiBhqI47WWSdqdGgeO8Fl+pW6nDvi4FpZ3wyJCdqhAIEbV+zP5wfzCNcSTxQks3ExqUSfS2PoI
yfoaKJKDr/jg1+tCgHMGXUsEoJIwQuTKxffUvmzL7iH7tPvSRETpugQYzJJJAco3h0z3iIZJfqQk
0w1N2/Xg6O8WowdehVtpuw6QQl1u0vy/zgFBsRuc4/MFVN7UlNvQaeagAJjydR8oPI56xQqWyj/a
x6txdjF3zO8xMvGG2LSk/9n1+1SDOrq+8sjAFMl4rG2rW81LbrSHCwjG5oJlkFuOK26nfjSF8spL
qXrrTzs2Tq3tvem5sXfOp9cscFbfr3RZ2F6Lvql1HAbDeC5h4Ks1LqXKdGTcBpTBZGFDGT+L3UIH
h09boaXN7iO2m5imkdLqT1QI2iAyroorv379VeEpmEkINukvA8iaM1Sf6fhbt50nxYrf8Fjqx8x8
e+4l6S2cGQH61PfO6JkgcgxfAn0tLisPs3R/Q+oB4T9OCJz1VipVTLvlkgsjHiyVX5GjbGeRyVJ+
/OuvFC/2ZqOtYPlW0mSuPuqR7AQIQFBjcuaRUeIhxjxwZokRCOGWA3waNeTo2g535xXFFU8OYDVe
H4K1NGNvNAVmg9qjHeK7iJaws3CTlvZ3dmsXQG+93Nl58bvICNpU6Bd9TxdPWRFLv9uYIkOBntzj
ZV6vJoKWky0fzJR949wp2x+j2tOaSMPA2POGbFsWbbDKCRS8xzHw02aHpm1/RRv4WNMcrvQ1zOmT
EILTsiJw00viHrVuxgD5aujR3YEUyOvx2CvAM7VW8PzuEmH2DYxg5EueHLjj176ofnsZYiBKtuZi
CtpGTwBOsNdjRiqS4gJ4oYRuV3/NOxE/3s2Yuf/ULBu6FHNMqbF+602XUqEsDrb71ACfFoRM7D0d
exdau7iuvNmiLQrYuHREfGuVrmBMVemcdz/zgihVuqNSKQitkpPjrHw2gjSyf2Wa+rOkY86tpPlD
bd56ikqetg82GLiNrhReCH7d0m7KvYs4Od9giFA3YJHEHXGP1CTuzziXf3F3aYEPRIwpA6EJckk3
R2Co772PbjrUNJN5/UvFg76FkixpNbdtvZs1eueTXXW1FgzONoepSMazf84nunBtdCuzGCQGosk0
4crvPaynBxSb3cB+8LyEcWkGkMTu9iMYcip+8y6IWfj1gvfi8VNSWWzvUP1dnHlNASS41cpqrpoD
TtZ9RA3LXaAUM71M5yJ45djjC5hvVc1CMYdPEJ25Ruy+9Z3MnUyd05mvMMFq9zxyXPWXjQVxy1Xn
F6ULm+bhvlrAETc3MRJR8zLeNt67hq1yDhxyEgWLWAEGQhiepCGZpBhuqvy0whv6GsVng4sxGhAm
9LYlP3X9XyFKDuoEPQnmi6scbXh7WIO+zNtCyOIHOYFoDUM1LUsyxDCiOMfkTi/0JYUpNT5Gu8YW
faR1kfUXbjCkuIzP7hhLXAT5EFv+snifnv2uWc82Elt05ssujZd3B+rTL9alvhFqu7cb97gT25fn
1F68xE3avO97Dyn/79WcE0HwJ3VHzV6dekNzq9JDtYehFVhStQlIMnK2Rwz7TKD64pMoEaqy89sj
FLZwJhB3xWlcXKUH4ltitd+yXJshTLkBx+KzaINaXUqwIjQxy3IDN9/RptkjDiCTLFIMj2fav/J9
bi5UzJOfcKJk9VYTiPxq4g5O5Z1IW4Ave1Qn0iRJlQSURZ4MSCCZXgSDZBwq3F2el0V7Lj8B993S
6dXoa2iXN2R6BmKnNDOv8Eqy5KaYlJWPcg21T3iAZNcmM3K/vpTapeetvU2EHwwG523cuzURXoPr
6nOPr33xP6cNRWuNSBCrHH+EI1qkZbqqCckEsvXGHxbzWIG9PVvoARBS29ZAU6MafbGgolTCTe9C
FgwGrJ9lsAUuiNQbziEAi2fIlmmLiTQg7Y5RY45M8coEO7oH2C6n0+VcXqk/gXgjmKY8pE9/dpr6
KlRkzhwF1zssnkHwSPpM4PcjkVzKSUxi7/aRlZRq5dMahqAoYPiaxPGWTuIpMc8B11FbudPKGRTv
jw1UKczj91DDLOr/J5Lo5DZuTGWfZYOW4CN/6cYOi6uF1a9QgcaQZOA+0uE2uc5o0pkmIE95bRRI
mXzsMj3eATnD0ipxR4E96/+ghLDQe6FeycFB5q+z+jM8DiqfqPC7EHrZn3LUyy9tYhE9+Fo0ZO1h
CTyfTVoup/v24t0zW64fpqUpFB5vTWcfvwcGsekYlDN3PGJM1VQ7BLQ8BZrg5NT4VhmNcca6Okvg
hajS5EfdY6Y9EX3tujAmteXCj/MpIqgyVwoS02GqcYJTGTDvoP79iWJatSsB6aWwl6T7l6tYpI2c
FpplZKGvliQ+1g2pyEPCqSMA2VWz3PtXZiFwwGq8vj+GlTYtFkx61+SyDxDHKf/il2pjlktl6a5I
V9MpdZEZ4H4WMLGxYXspQSE0Dn4xZhogaUuTPFQRJ5ruIGuUgOKBhpNxLUpc5Gt3CSDQQTvYtcZA
N0KrYiXhpczrAL8NuyGdJe6QybNd8MWWy6n1qT7aodGD432g7IcOmwnb871w6Ird0JPwxSleCaz9
mIws96oOmi4BY+e6O4Cu1QpGVEOG5tzsnY3Hfxm9e+Gyo/RCV+FKQ0qwr0X+AePV7dv/rbTvh5Lf
q/ncSwPZ6zuNuBULRsyVgDnq922UhQ5+/NCeM3rSm4Ynyb6yhayVVWOq7mc2LrEkZFW6XPCruhYe
OUxpF46CcA5g8/FYRbVwEAziJupsTz6PeIwWNj1LRU2H9AQVb+ilUXwx8Odeyxpi5zEvjFR/M45k
P57RN+nR4AKca4fqMWq5PFIDrcvLu97562R+H7BGlUrKpLgmPSNAjoMFRZBLPiqGwpl9Vh0ZivSF
vx2hrniPu9ExC6/3OQx9W6rbU7igoA1wh02Ojounsooqe4D7dqq4lYQJ7HcmnKhTrh/14FKa/Fgi
rUKKX5TzYOnawkTvF6H3IACs1YriSrUDmKEWN2KdMphB2X5l4ghq/8TDhRBtUsgKCNAIXR47mYeY
qBRforoLa4PGOLnq0S5dX2lMvusSThsJ6sAi9SzHOzGckDPmuOw4Vl1unRVCci1vwrx+qs4aPTkF
majCiRajPeG4frbw9hFCy7YZs7YdqZ6qrkquoC/ZcAqzoJ3mdv63gnzVCrTYNseDxfTl36G9iQO1
Rwz996vzmW/hLmh5LnHVP+MgWZVyMlQXRZdSflkPTwvG7BL6KPU4ICh33N1xM4K9oRFP1nMUcwNC
NqvxvvrfQOP5h2FxkwQQQK6A5E/MOV65JNGDR38u698LjY8gY3X+fM0XPEOHUoRnEU4aaocLibYj
/P/tc91BU13HnLinMB8bxgbgLTqp7A5LHlgHCdwTBLNckTQmShyzOHzDyPIfZL/twy+FDlfFJpQs
qrQU7bL/HPyvaLeFJsd5xbzEX+cPUOoA6EhDQkWgeiHiYbUQ6Bik1Ge2s36oHEZSDb8r/icymBIX
hlWZYfHI24ALHTeyDhVt0NqGLXiPvGP/PB7KFYflcLrI76B2VgCIMckErQL0YOzvCwnFl0NEOKZq
XyJ++Whmojg0HY+AkoYbpqm2fGb9VGU2kUKkNR0MhNrZS2daVCzpKbWhHwOs2OmrbkFp1gJ+YZVw
/jVVQfZlKUL9gcLo0WrYFf9bDIM30OGMs1M0sZjrtlRYai9Z0SZvr2tFBSn9T3bWRhpayxVYbBHe
QjvEw70Mjy3DQGeXuI53k9UYrdFSh7XuNTtQ/hg/xezz8pqk304DWYpRjDfqCI0wEvSvO67wxKt6
JTAPj9N4nk26PFt7JtEt3OZ8jbdSoPdZnDBBkmducoizl8lpLWcvKx0ce6GxzJhpak/Dg7NDm6xd
IfiMJYjiNLNbYpHemqGgy3jq2LRuthzOKhja/9v9zkUjwncFC+ITOBCgIKaXcuhNrVpgiNBIeT/0
CNTGBJ5Dpq7da4B/ZzL9ozKcb2ccEW7lmIdXILL089Lj6IUrrRjsi3pXd54R7CuVL8qS6U0m+pHf
fUs8nvz+1oP37qgduT0dE2dJoyrx6Cz96/nyDc2cQNDFNpjO8GWCpe3tEReMBELEmyGyvv2PcgK7
BQGredSjbKvE7rbpP0EupxZgXh2CTmlHrbiJyZDpKxmrVJ0SCMr3WvJXX8kz8vIF/qmPvN3u9/im
nMG5VlPf8UhO5zFdqsn6FqHrs0ejheNYFq+Ul02HnYeoEchgn42WV7UBN3/aKKFX04aCZHVmn9VQ
FHNI2oeSFDD/VtXqB8SlH1PG1mr8mtFNA2wPj/WBGk+ANmoE2jIo6K6TGwYJpSPI42Ld+lH2vGIo
E+551r+1ZKpPh3EeMi9C2KK5JefM267Syu1U0aPqVdmnQy3qeZ5wyIKywtVjSg4q9Meg49pn1qcm
MkQD5IZkaRWdBxE+H6YGI2k2nlcGbBGpz8ll3MXPfjsuXulrmgxuAmzToniskHXJfacOR7PyrB7N
QFMFtNDDibwtdCgQeWjHnC38C0boHqt2rFT8l1eGl0xoym++Wy1/A0wlCFTSGwJAS7hlR7tJ4kuo
LKD85N7PqZ6JWjRenaFOYAC9UJBLt4aG6SFV08pMXNeDS/LcJLlaHFeMOQdbYL6FV62Z/JGk1ehS
JdZabn0RA98BfJyJJjXSnkzFIdLBnk7mBkqM8o5LsA6ZZ3Pkwf0bBN3GvF5lm3cdXhCOJMz/Yqto
sBeFO/lJbUBI3McisZDIvlf/SfYK43rvp+b7ngZUo5hKDZ8dz0EphRK5EfZ27WNF0Kzqahk5CE2b
+Q+2F8Y0RWt/eMVGsN6luYTm+Zla6Fwm4aDXiYl2TgFs2zwX+j+/7Odi3nrhOzQRTz4tYV0UEqXM
xnwPJ+KWFrFSSsgkzH+8TDHAiaBGTk9mOz8rsMhCLUezgYebv805gMjUXGpkK/I5N+iYSP2byJqK
lZptgB6zukEb+z90TQyWba/QBItNDYeJ8bigB18a9AAJVuQkxb515N6/SpxmtdeBWcYZOdtIckuc
qpCMrZHFnpeQ5ncw6CJlAzr+AIMDm2pxuWIkvcC/3HVxape3VeJawMt7CqRBxmB/0B23KPw5t1JE
EzZjeu81758ZbLfyW26MlfiXNli/tUUZ5TibSk8NfE8EPUocPqpc/BFnUraAUKteyM8WRU1MHmBM
2xkPH5lgHacGW2F+9AmrD0wMA5ZbF5rWxZFA0IdRxUfe6vqH7prjrStAmKkFHdk0Zy09D7L1dIOG
SZUaU7fo4FlF8y+uzog0dFEuWhzG7DLEA0wQeFLXlfloIB6nk6kZidXIRBieYkwen9r1yCrn0cy6
zNDFH6VfiETtWfk5KNtuawGeM2jT3Msaf4oKqmbiRsf+WmJiFVhVLNomrN4pQ0KfZMABDVIbdzwo
XKHi5IybBc4+vwHmE/qXaWZznGaDdPIEBgjyqMUxT597YixWKOe+/m+yL9ILm6V+zINFXXtzswE3
EKUXuUj8fySYMKch/BP7+B1bbkOY4HPGX1af5QweRwjiar27zHi+jKeeEqeUlqFJW8xj90yF3x2L
9L0JhJ5S1u1SeEMyT2zwp6G02tJms1+Yu/n9HYrrWnu7WjXVgMQoms88tDJR+UUgMtLPjm6qw8Oc
p9oZoH7yclR0XIA86nSxFhQhUEG8wz/4KJCieXb6EATA96J1PZAmrItDDQnCcH19zMPgNdE0QGju
fkzecGQX/RIrGzEGSabOQ/3Bkx3ugNZImx6tq9FiSYeo0n6B2wWQ5a1HJGF3JJfw+1VQ20Yu7ATE
tFsQ/oefo+hr4f4MdGhiDZrHRtPreExzJr7KXyqIylB2o0YZ7vw0avBggLAdrepOortmPeVuJEwp
x47Tk2doi5ufDhuA38EF9YtQk6EhyvNhme9bhBz3nleMqrc+GXIpYhfvupUGnG7pD30m7yJpPJ/O
IZwyXYrSiYOBK4Tox9y89OjjnrOWQt5S0yNJfZFR2Ve3La72FgI/bpzX7EJkF04bkT4UpjL2DXZF
3vD+4HmhBrhzNwtetO/fb0X9iR8ZeeNjci0yt3XVGjo1JBePfyd2rElmTAI/rkh6KEhNl5/ykWXf
ep0sYJJySQd8xOMYhAlJRnYULefgYwhjhzYm1hmdozR7vfmyvZ/xXZN9E+RKlYzpvOFpArBAlrTU
G2IjzeB1kKblclJi2owuWrDQrTRDuRxHoa07LgLPPTQ5tcdIrya523MuiJ/ove3yj3+g4THs2SLx
xM9w65zILw4bY1tsTb0sUR3xB+wzLQ7E1Wzrq2m8IaveBdr636VIMmlsLm5rSAZ2gSHxTgVNxh+b
5cTUywRtK8RZD1P0prnd3b6rAnO79Rqy/0XtdTfelaS4K+/KcjaMgSkp2k8dFYt9GdprBKfz/2Jt
cPxzcYohM/5aM4QTct+nxq+hAHTPmS2U04WMl+QZb251ivEY0ydPv5OO5pcmNktDwfowSOVbVN5E
b7f4tJHNT/uhxTM6FWgSw1PxFVeLgraoKeJWcxkCMTB+HBw6q0FcIzMeyzBtyLMoIxupGlNqJJfc
bgrdjhbZlE5o554b7Dtud4Dlrkr7BEhiXqJ0RrH+j6ELD4W5vEfoqanRVBtJ58ITriyB0MHyAnow
fflJwKP8FUO6fioNs4+h+EqjyIbCj39QIuY//LbrfXivdaZY6eSZH73xcWFCCfsE5ybz5k7C/fr8
vwp0YZU8P3tgNvOUuCJSv5D8OmmkRIgAIeuWlT7exZLEyNKirgdDT+bJJFIKGf/73sswQ+Wz/Jkq
Y0uW3ZCTB/yF6a3hWe5bYNKCZp7X1Xj2/U4onH3sPOL7NIUeYONi8Z3rEYvSRj4U7K1xVdhEsNR9
kAUdefya9uVBlWMOb4ZeqMYSZoAiGA321bCgJNu3Jnyjt3TjYk92zejtBG5p4WD8rl7X3jzh3Re9
J2zQ2Rxk/STUeM/FCm+sRAsJ9MKHgVHbajhrk1hlun1bm8cLqWXF/RC04yFTTYWNtRjOP18J1K9v
C7yligfduu8Oh3ZPSIvvdtfvZC8jMgtSI1PE701QhPTEIGls6tiNTwZWVfIBHmlkBs9TnFOsQThc
WRe21pg7pmW1JmDaiKaUgC5ZzzxyhXpFqAjSLCOT1im91oww/J2lyuFz4vDhaO7Auq8T0x16UM0p
A1UR8INDRejFVnljB9aDL+U/PxNsPCM0drTrXvQEXt8aUQA0SP1q/xWgCN2sDm58vQL32AR3QaFX
v9/l06qIZaqaRcN65vqSTMWUz69GHzI7QkC5zZ7qXHuJdPWcZ/01fMwUaY7v2gRJd4kK4WDHW+9g
SZZlbo966hCiHxUUhuf2GjzabOUwZFxs4/B/rcf49549n8ACWpeA1evgprXvYzMHUGZE0H3qfTd3
6B2YXkymn9DmVTBaWkds1zQLMD6L4rYXVndUM32LQ+XWLC2Fserxn1vrpobnjgdyPK4j5Ks7vGbF
/mYNh0trC21W71dv7VnBnl08urfQAYYoj6OLa1t4+5Qwl9xWInrISy3mp9NaXP7HwdvJYLF65rD5
Ah2kenaQW10HwqdDnX/+LtNj3cxrB2qwFwpBnw3/T3VCtepBfcSSV5iv9g+Hm60a1xJUGAvyKdE0
BaE+VxecTvBEnn2BPwB0fpUYDW0a6oQPyqMQkI2Q7OPnq5oS0yxUJvAMILLt5nUHpZNzdX4LNheC
MStlyHjKUtj+Wa73iX02ayvQCdTtG/Fc5mBb9pOkyD3U/qvu9UjN4g4nypnjtjUAKM9HRe6mLLVt
Xr6W5Yk1tCcvq8+ZGqC2EElNzpK8cVrnsvO+l9kVT2UZOkghUq2eSS8hTeuLr6AKBh103HUalYfF
l4CBtPDhVBKtGQfN6EOhcfcH6B+h6Ygi27E9m5IM363P3COblqbKLlPKaxVL1UEnAlwpmYhl+n2m
DL2TabSIRme7wNgzJoh0Eha3Qe8wsnvfhLgrYOcfe/hk0ItQ/z+DeBI+EQY9hflLNfz5kvoL137E
grsk5wU/jnJ5K/iPfsSvXjdFomAPKlTJVhHBUqEY47s5numCGtnB4QstUIPDqdw+zw7sI6+tmO52
5syLNSv3LSLuaNb3LzwxSE+FKTcoqG4Rmam8nX8hKjrKun4AN1T+OXoknXR8QgnKkNfX0Uc05/ic
+lKkXN3HDN1bfV4EPhpGzyPCGgXhu+uOje7V2mIg/8ofB7RCDe/yAWlEM1b6xcwWx3GpCA6q8lMB
1wHnajHmPtYzcynF285qAGN/WDHBJfAPLyywNR3AoorYFnNbHMTxoKJ4edUMLDgmbRKitVpZR5ze
SL1JA6XrjjMSJFD4MOO1beTBaA1H+4+5iv9aGYp1P5jO3F67Ir0nNQCfgQpltJVvsrIW+GLBVp0x
/1/ACsgdXSOsmWc2VZMMzpQZUM7F1cYbdGm2TA46F4XuA5NOp+LsmSUiROXE2bQ2dVVGld2DxEKo
XeEZN2VJ85siUcxfHzHtG30Vpx9czllEFaT3VXL4S+2783EsJzgYrkhdwtcyE1gyWvZMrmUF9w8V
ka09DV/r/82oAG6vC9wceZlFq75qs25+mdGKcXZShRydOj6Dr40tsnAsVhpNpzRGWNMN0X7/F3GA
UZZg5qwDYk2CHTSrdw7RUX5b6ZKnATBzIJskDIsZUdOiVnlW/WiLSIWpfSdrGNqVWm8xjGPYVhD3
/eUG1yhSfHRPolIfbr9nVj2mWbRoA3y/HBdHSfHj3QjLVpeGpXlMQIBAy3X76yhp9coFR32mDYcm
75cXR83VkvS4tXxFAXBnVcVUEQzvmV9Jj2xk5QzkugZZrgM9rC14XoEEjwnXoO0zEEynuNrq5RjO
pnxgnQjQossXA80LaEXetZuE/TmY+uVNF/53zTWfGfO7wCtyk2ep3Dr+y9btmJtFB7JYJbxUrZOK
+osmS3JkupxofdpKClH7yeNK6ObhWhv7pcC7vv6xcEHNdcSwxJFjLqHYFMbfP8p3Bqf0NjY4DACQ
sf5/qo0hHp8ugRYfea+TavDAhwz3f5D1kYqJORdkfawgY17EEYl0XqGIEpXSgWGDuj+cnA47B/83
tdMK+abPlylckZzKjsS12yE6q9EuBIKg7DAU89oA0UXtXQ3kxP1D+HI11GFjZzRwOG0WGK0fUFu/
M5TU8pz7Yfwfcfr6+Ist+XJOaUMBEoZzxXyo/HFsP0/zwOYbjkhEdzZnyrRYu5XIgctQUBCGKlxh
Pl5XVsw/Xo6bPE7+BQuDN2EiiEsAV3nViWUvPN11tvvYhmv26EC+ubp036IWCBhCvSBONo2IXXcL
DZZsEAvCERzWAN4f1yZB0Ap32XaVEvuzj0MOQI/JpUydCdellU2X+h/tVbIfJgFoaMuvC27EvEy+
ry5fP4IF34yBLvJmLlHQV2pEL4dwGwMxeasdQCyz8YQSY/nLOq2XZR41Diqh0IxyT2NkDKCsYyvh
KldlSjGhITJpEX4iN2wgOqAvnL7mYkpAhnf6CJW5oB4UpM1aZTSYQ0glMYF0DgzEPgEQiirf52z5
39WBi6YrZPje27cZLaN02oTtFqwidJc11RnRtMVaDm7EFtTvcFvDamBRct25kgBzvmNkBclYCnBy
CdOWGtNGDYn4m3/trvQd8OWYkw5NxiDTifJynxzW0g/G0KP78CT83GKW03N1te8YSEHFJicczqfI
CgGJnr8sC9fZH5c+S5flaqEUITE+cMgZk5K1i20TpEM+IvO3EyNbXZ6Bq7tE0e8V9NqCnBirjd1k
ugJZsmscDj+owvwupjRXmfQ4qGTntxilghFkUQ5gfV6vcphzsTpNt7s3wjZQGPouCj5zGTUSAbgx
HSy+n9yh3lAK0r1NyAwcZ5q90kMXju6/XbFae3HKXDTxgWQr/tLwwxZ4KyanuBmXWeD6VMSX4try
8dZRkvS3rye5eY2QcDE3mBQnFMXW6mxVmKz1EJFSOGs6gQOJZimLiZIqA6vZSGoapWWSpLDYpiE6
U2xfe+Tc5CJzC0Pxhpn9GAfewXjEs8Bfxizx6ZKQZ3ELv/5JZq4cFGKebijXJeu7JpJthvZWPV1d
3um8duAkqQIQY9VLZ+qanRCgPMKezTybR6qSKmqxspuljZnNGwLta6+JvwmYXNMwugAjIgdJFsVb
3moRm9ExHboOiwBMMNvlB7+h+cfjpvEEyUoMaKzsI9hK/LhCgxIxB6I3sfeeFFIa0KWsSmGLFyKo
XfFz0GhPr90zwnIOFqgQw7CVjFozsAEvRVujQh40+A5Huav1T4aG2gO53I0OMjv0r1mJV8E4W8Lq
q5RHhojhiQAKdfzRqNfrZ8aezDYOegp/fl77ry6gq6j/rcTWAl0cpo26zqq9LfhOBLtgSdkwzW9S
jrlc55Ld7eoXeQ3U68thTCybCm8D4n7Z9UULOL6nj5U7VbZ2YSw2pRWC5q5TdU1XLnPfePUKqqX9
V9qjAEWFnGUflCUuIIQE7kEcdIz4Ep5yiu2O0W6klZeo3vdl4oGI0CXvwjG/cF1OMb/eOPoNvNla
28r1irsx8eRm1Ym79FRGiuv6hF+0fKLfochcMsf7N1OvrSOMVkVVuJYN2NiwU4fEHOc/OM8MgkKi
/ATj4lSEJmSGoiKJCyXFasFjp4YQzwngJ1NNV3ecYxNSIzBTByHZUh+msPlTUSYrfr391E363/Qb
z/cSTNfyOAavH79BubfDLqstrKtYOq38PE98hFizbUfjbFkgmFndZyr39E4r8NU4ArzeSr5QnYjz
Zt3YmJ7zDZgGmM/INLfI4qHOXrmhPhEV5eIk8gzZ1vJqvpiHc1P32MxZA11z82s75aDt0RJLE6pW
gJhBlXuieFPtbtn1UxNLTjPOzA+kAbUk8lU8TvV7ghR6khA6dDfYe1cuD2WU9tPp/X+nIlOEYvRi
16gLiiXN+flMeSB6F3xrfenF92QXHMutX4As5TJKi5p9meOG9C/nYlUvkFHC/CyY9v/2J37utUlc
3LR6qgqALfLd3H66VXnh8XEPzj7HJnjigmmRVcaI0rZFh/XlGVVFQVDxqylPXrSmv1Rh5ThuyBuV
CtOZ/uJg8KW42NKzybQF8xfFRFuVjbFHDP5vde6vVuD1s1LtYSpLuz9e7Emn7GBwiJvqZuE+mSMz
78Seco8Ja6zhcuJWOUoEEgsB6NFJ/H++6qNOb9aZtFJFKaIijKYE3zOYhQiljqY2d0hUG9fhjdRD
0CFKP4rKdYSSFYx9zvyjfmSn9Ej4rEeopRYZDHmqXvG1kkDLEXrNxIm5lTOPbOndxL9sF4JWoCs8
VppzS+2QreMEVNxFRvM6eD9VRg4GWP3ehys6jvN6Od+ks46sySuo8T1HoHhRcmaMC6Rc18HcOvCp
u9nhluP6bHOqmvTMMgt5+cENEUAfhsEnyVKQjK+b/u/QOJq2uGgxr+VyS7Bce9h7ZBbUG+z3mWhv
FMas3+v+LPBP1ufpPkai47ZJ06ExOmfQCvm8OUtc7jTu3Po6mYIj4K87hS8jcO9M7YRbT+dTbw75
j7FyiwRE9VVCbJWzZRhVuov91J/uoFwj5IM1yUDiVERap1l+cHkUIN6MxngPduH2a2KzCeGJBSo1
GBz41Q+DfdKMQNMvy4JvrOUOs/1yk3l7XZyY6now2IB1r00rg1V8AjsxI1g1eGswIvZTrbTr7T/V
NO08hF5ZoKtTscss6ySBO+1m0obeWGodyH0+2rCfW0W5W/l0rAXb0cbbGsLQQJHgJL4nELmZLtH3
8cPPCtRc0U4utCWFmmiQAcjn31e7NOCJaSVD8yzbB7GD42q6UBN2lAAx8REXQiRP4bqo0ZzHzZi+
buKPw1erXCCNY6AI8gbbmWWsJprzwCtkoFV8G/Nfwp0/2Elh353Z88ywE66waCkXlqBmlkT3G1+D
HIRtNm4aE8Ho/7kNaT02mDz1DU6ekuOnLUI0jp4xrnFULSJ7f9Ym5Cu7KnMpdkiucjEBIT5Y8HI3
8Vc9BZTswq27CS6Zxjocwy6yw1YHzt04i2/XJ2IqIo2DD4utxJ60SMRA0siVt39wqYWpo6Id7DI9
z3Jf2ED30qfRPIx04g3ThA+3wzc8Oqj3r59FobmIXNF88bXVqXBntZCt695ekOCSomiq7w0X6isI
bwOdfYJnvBTSbUev4VLGxdM0uJYkshnBJkbAHwL8Z7Ta4bn8P9DzpXWFDjD2CEyac0zsAQvEVS6+
wVFdEauAQLAWS85SB41NOqEbjqXvfBGNrMHQ/vt7UkjEU208qVjfC8uKPbs3WQZqI2ktVDP0GuyE
fxTeLygyoI5QrqPpbdSavjeIADJ1UIvtfXSZd0sfHDMEg7iOjVY+qSyGhxvO//E7iyaMaudH6SjK
iiYN/Khzg/N4B8+sK+qs+2aF35n7Nw2pdbwyfs2n4uWku5AjrzCMfxKoZ6vXXf6gW28NaJgRY3Cq
T2NAQ8hVkHPW9r4hjauWOaTp2eYITM33ekxLzLYDCFiO7SjViGB5LxjRnCWJD1noj8SSxvmG94UM
n618B46BKXYRPGBuAwuDtagKKTdivzaqRUZnWIf4Hx9BlC8uZA5yUDW4QJWABxpPd1IEf/bbezrH
lVBFvhZ/yGOc5PJ8f9CGwB/1nfFSUMQLLhAfKoMDbM6PoRx+zfAxDEZWnL3mJGmj3QLzySWKUJH1
gOxf1cJr/8xd0m1rLVbkP4BhtDt+lThoIHBcUoJ7Q83zpyJ1PK8W5KytT1KWhi3RvKPDhLGu8O6E
/nDt1M5USEC5R0cyuzxu3ctNRmnUtt021QDGuAFXikQBOoeOZyCIGFHP7+fBswvmXwlnPBFDm4jt
pPMP0xT5J2PI/pbsmE5pOMuon3gFCDuxwFC647QNKZFR+UZrFfsBv82Tchz1rtMunAS7ga7RN42W
g0XoaGOkV5LmppvkuIb42ZA+4bdMcRbDs9yEdYnRgKhBg9P8T4G0KgFWL84VIqe8h1bscuCiKnzT
g8Y3SAuU763cScfcK6UJtBpWGdCxExEIFihYWGSXaAdW9nTZnLmH6gwvZtCFhkijyvFhYsTsZdzc
nG5Dw3dFFnFS3x8eQseLaHtcL8zAtmGi6BRj8AFsb2nBOHfap5nRav44Km7QE3zV5sSI8S1Zz9ga
PPHzWWUiPl3y4GyxffHciNZ3Gcb9XelKfxEHy97XtAbshm9e/+w3xz0Nf2/w1VPMjmHbKxapbx2p
DkpR5LjHt/VBNb411Ru7s8bylzntbhZd3AlA+P7N5D4w83/o36L6pBtTjLTQ1rWxr9pp9NcBkntx
9M6wl9BPknUA/i0oeAZtn60vcZOwcxV2QJBDpDGZbQ70wlf4Ljfd4TqGePIzZwjiH0ooVvIrorxK
jf7dM8v5IDRVWQTRNFoGyp/4JNhpwPN0oNJOk8vq1xWv5kynywLhP7WcHa/kFxJMrKEeTTcQdbTu
Kt8O6V1SuRjZuIRKtCRwmXqXW6cmaC6gaMOGZS8Fd/NqT8/r+BN+t1GFcwX5bMU58WrH9ZTAEzpa
gEoUw1gqPlW0KhsXMpfBLbv/LXo+almhstOLF/voH3I0xLu248OadZMLXrAy/BgQPJ6ilsR7Bmat
PeQ37dJc8vTYnq9ihH8TcQQAG7VQOGp+jFz+jnILLcSCo11+VXAf7QNzxka9qUQLHnJ9mDmk4oFG
yVGcv1lUXz8+2xTstIR6VVre0D5pplQdShb3FscKr6+0262ZRWt603d8ROlIq0WLV6SSYK9937ic
VcoYehbkVGBn8Bz7rEoHf3NyLIg2EEdYyELBoOIUdQ114bLhE4VlYMrl6pCdVa1lYQ94JDmX1ffi
+AXHPIVPEjlDbLfx8b73/Yg8BLE+SuPihTrCYLLwAI54YeXY1rwb42aO/n9zlIdPciUUCiJ4WpgB
ZiKrJWHJUYKiW4XSARRg2kS5o87ZCmN62jnWqB90567X3OlQpdn1BzEiSZ6Lqt1M1v/8apOU0i2I
80ch4pizlOA5syWynpcqUGXZd76a8NAzlZk0/RuCblg16uJrhXqDF1CaVxSvNOo4B3Jx7K27IYis
SGu7qGsVxgm2Cp+vHLQY5xu6hjtVz2rEop8r+KgEtBtoN3UNEzyCtflSQ8JGJhC6br6bez6Mz+vT
IjN2I5veWUmuq65W73mEbEdWUDHyZaocJ90Ht9VJljLaVs1WdEJ+yE2lI3M45hXyLXUKKct2SW3t
UP0i06XkmdDeZ78UhAcRB2oi90wB+LalHNd1BzN0cKaQ771dxUoqrIHGCw5YVSrfJPBcdqJ7FrzW
mL6eAME9dhDk0RwP6jSRHjw1+mABLHIQNUbabGqqf8w5mpbDzrA8ZXrNPFjZ3d7v4mB4dOK1qv8F
mmynNd/KcCf6/QxN5s9NlH8dTrQyxrxtAFNjgukqUAJqTfdxaPpPFMEVcMznXyTzhfWYxpDP2C0q
UM9OHdhbKj2Us8PeokNfa97t2ewBdU0pc87yoPpnFh+iYpQ4osCh6VbdNHCZnAOed+MTQq2q9+J8
MddJu1tIHpQIfG1tlFI5V7yJm70k8KTaNXQd4a7Ay3PQfjIgHOv/8EMWsnOVARo521NeGItWByvY
j8zo5kCsGa/YL2oQdDsVOn7qitq+fiajtRaeiBLE4j+DM0GM1kfOUnPPWejDkHevG2IOMuNtJScq
vBFaZWhwriKKS27ywCiwWYN1f9NUsFAUgsSX1SuTiVq1+LadxYOhQAPKWUrbQFBJsp7rg3MnNmjn
2XIvkbYO8Wh9boLNoFTphkhDU/0uBUHVMvDmBMjLtdcmTmzz5PH/PQqCRry4OOL/0pO50p4uRGCy
LHHmaLeS1YPofO+Qzd6ClH2HmwQDE8/jzrEMoHiHqSl+RvpsrklXVZl9UttA67wiC85ILdIFqCJ2
/Jj0REYsbwQQ513bBcd4B24GbT1okVWjEqzferFRBI5co9M/Hd9hN4yHtRFHHwwSeMTRagBmTqbE
vPKxAlWFi5aamaGrmRun6lR0332TFyz3jrdjNtiIvRg12v4USSMn6TxPUgjFEjw3Gr6knx56IB5E
9lveuUS+oAd0kmrj2XBkBmLn5g0DVnyVKSHOAmCvLtPbYkT7bNK4BPkz8Zufdoc4+GBoqkqTmqmk
0lk+Ud8oAyqPRoEJEhIQOS2I5H+F1GODJY1dHeg1uR81cPs/smTC6jyH4Ux9PMceJR8XRfBIo0xI
VAXdAHIScHs2BR92fSla/IpRsEoBwfrwsLvoUaD+woODB9D0E1GG9c9az9UVWJT5nsLVNSOLa31P
L30vyKChB/xX1IUg/GQLYlPxfK13evfS/T2w139khP/NQIPqlAETvDKODLq5xNDHLs5s4pB4uptK
9By2n9EPEz2VGzrCBiju8TA7lFkLE8eKmFmHp/rTB3PVBzQPQzVoGJJRWsFzHtWfILSwJZ3mOKUc
WzQYjBl1qTXr2r6m+rQPDO2wdV293lWpArLgOqoSRJaVVJxK2StBSYHqA7QXg0Ql2mPOdqWozscj
YxrsU5XxKsSic/wfbKklq3dyIFCX+iVKU3XD8HtIarzQC6s5GjUhMlqX6wHwO5U5GtG7M45qPfXJ
zKEXQ5rxIdXHJrLzmE1OyivmhHOnq5ZY+buett0k8XvYheGrUzRm4a1R90NGZFbfvtjIJRaYHm8J
K+7A1cJvdciQSmkuKx7b/GCtAVGOx6P9Ze8FSvmSMkaFb31hkA7sFkK/oV/VZHFUcPtfSGcYp7fK
KkynbYGMYWAmlj0x/joQebjs09uIiPeklLFTpEkjZQf7JZAq/DAbN4PqdgNUXzlRsZpaVImj7IOz
Suq1a9MG403E7jc5ZlwM3ssjMyFx6RnzKlDTE1ry35JwcyBDNbe2qapGqDuIJhPeFRtvPtg8RYYn
+VC8McM8Qwr5I5XV/szDfcyrgbOPpQDC7QOEekSL6CV/QJwpKLKqpaBz3dWaNRv572LLx9sQ4A8L
qlbTUDV7hLlH31QFiv1e5WwxTsqO379B1lFrOG1TGtBEW//A5NQyFeFYxyDsYvPZopVqhNssIM+p
H7bX54iTUYmoDLEC9YQfqRtmiw/nUFwrdObGDvoKdh6NvHHajOVhxO9GtQYdN1pi4FxgyW5T8BOJ
iPCpIK+4rzGhkiaJocPyqT4RP65faJZE33p5w7QZZCFhv0P0LExjFT+CvxABi0k381UC/c0R588w
xpoNKSbauWhtuLCNu21B/9LpAXntrCy/ySghZ1XFYMC/yeMBmwzVfAAeS6SzKWH6aLI20xdtetxx
PPQZLnwtqi4TVs+bjH0L2BIwxVZdgZETd0XyfOThnBxW2NP2PHf7mJe7r+gZOpjxs2D2K/DoU3NF
nIbG9O1+D/MltZXNZsXsT3Sq36relINTV+U3B6K+1h2OO/MVRkIKgfmNNtMQQdc+iu5n0hBCyrzN
NMNum7mVO8zKL+Euq/JDEPtMn8mOnAuKbzNZjLyaIM3wcbfWLDHaRUMWbNNMj6sjXDDCTD1sJB+k
64ZcqtDo1E+525OqMKAJNObsm9dcEI/5VhxbybCEyVqOJp75W6mkFcBrPbKgxnvI5arv47MVS3y3
Hv1wi/9G7aWoLo+Yb4AW5fG2VF8qIWF9jiMtR8iwBIqYCalfof7gtCkmzFJenstF06ZHW6/01H7D
6lbCDUgu8HS8PH9rqH+ve7VWuU+NJjQtPsG4c2QbkEqWV2ZxeM940RaWcC4WZN5BqwelbucR+pWc
fUL4cnWU5cvAMD7n25hYJx+gizMNM1e7ycrpvBzgY8ti6fTNajOq25gKFVufGGdZ9lxC/NpudvHM
tp5aFTiHx65ubG0+bgSUfUqRcYrk7UAA1MYXbB8dr1RItBlOMTfdflMZHDi5Hx/5+NkD3J1WMMBC
JNrklgdNZRL9LOACEdZp29pghl1/aWGoKhk5Vx084YhM2qZkSHkkwJNmiUgv06NfI9bPbp2WbUg7
dndXwdSuLNEOpw2DR5AumP18ok5/gFmRmyJ0VfO+1umPfbQRg1h9A+6eeVGJetXsjUPyUtY+Nhlh
RxOxwt047DwPrukdTHB7Or3J9YxWa2FgYEZO+O9Ia4hJsubr6O5hQucBYME0VQKKdfc6gmR3GTyX
UjA7ZvYYlBfYy4mA4mKTRfKZvOlIasN2O6UYwIgHHJ7UYEJmm7TLB90WegywW+rxQ2moYKACE+R3
aW/1seKx2aeGbD/pwJPba0B8eBiIgOSlYgNvwa8ibv3DsEqNBZxnjofeh96ZuYeZ6ZtAvCoq+Dfu
vZ2KSc4xzW3SOu6uEz7kydop1jybllKx9Qp5ftcN4wSzR+yTkDVZMqe4RugWGoBgEENQcpRLQHGE
TJUM6rtF/DwM7gaCSn/hJkUv+mQqxlaLILr/FWzrGXbJQdraXfYwVpi8yBnMeszAvzssG+yuCg+Z
ybZiKm7N4xV7q7NO09QB7ORlKaSrTnNKqDIn97mjK6c0uwy9BR210KArqT1hz8a6tnji0NTIxUXl
lMDB71al+bW4sfwGWb2JBJYueYGlx050bMiStj2Wmn9UJFw9sRNvywEVCLD3x/K5pYrFM0vdIM6Q
4/WMtZgut/XJTkT5IHkwNT7/IzmkydwTWaKFQhDoynGeW0SjEyZELVE/mqzfJZWtNyI6UiemhA9G
lWDrWC0YYO6CgEin+GouMEvxiuAj7tXEJnHFF9uoAptashefaHUyaV7Szs0tx3mus4jIbDKHvoLM
wB/edcCE8yjM1Yfzb2CbSCSDckXraSIwUCNvSmHsVN0axNqrzjQZqRGOhcw4W9A/nuyxyzzvdS2X
3AbRwduiM71X6koT8t1zlfFWHUMdWAJhKnGatqAutXgWCWUXhO4sGjOMDz569SeD6Oh9+lj2Oek5
zJDiGJ5uaphTBY9vOtwI9BDlxuNjqn5fJVedJAqdaeXcB8iVbo8lLaI/lUmZUIG4y3/eUZOU/P2q
MPcUgr3QNDIbYl3v+g2DhL/Ov+PPe+eZQzG4sqVzTQFiv7mJAYkR4ZYxqRwVr+y2B+96IPdMQMYS
dGDic/hlOj4OSKKsTaB1CbV0bjHXfTAMRLk80ZVzZH6ArVFIbwZT+/yd+w7ymBFu8hlY0N54agD+
FrlbYJhmkuqTShLB/joDpQZsXM7Kg4rMs0Lp0A+VSHAw1b4RUDiIWRbQrMPrafwD5YwF13vamvEr
6PvNSw4rWNFXR/uSV2PHbUhKzKY8qbeNzEzxpimWJZLRxO3rREClSNfhSwHjfAsip3s7JvZ96tOp
2ahEgiiNAGKJU6iF+Ljkbx+t8m3MXCffn1gEljja3l+mYq0E4JHp8bDALB3eSltEMGPErzcJUecF
hAXK4M3Zy7uGJWVmsF+iVhzmNVxzv33mkKmYZBO885fRasbTfOGfMi2WXa4VV82ulKCU7s8UXFR8
iOTRhV5C8H/r8dvv1NxoSdQiXyOkoWaTp/HsjIIoTkfwXb9WV1E6+P/FFYtoveoTlMXx2nA4G9NP
LdxT1BjmaEGhx2l3JwwvhwV6/ScaksCpag3KSI+0NCrVAZHKmuGiwoCthe3OcDUQBiXjXjo6crYC
V+aXBOoyBxG0+BLnxKE3DjfaDmvBtz/4wLVgiRRd6nNtefu3n+gAJbkYGQptmj/T758loLmbQiyq
YPdjT8sY9iPOH61JmDKjpw4laDJlVQGqblvz6dd8vibllBmdcg/EBgd3NFtyx6V6GjT84RWrpvSr
JEdY48f3c3fNqvKI1NSnSG2w5gfYkneIDWnqOp3GmoiS3QPsDRBnFnI66cPB1WmH6/Zpd3Zd/Akn
kd4mU+EMJjWJZ0eJI4PL8/SLtYIfLWvWaSnJkhduVbULuoFNcOz+msV5Ai5hpIi6ZoX8MZp9DG4E
00y9GsYwcFwEJlQE8CstWbGmmoJvwormsM2Y9a0DPVN8e8lmY3uXeWPpoi5EcmorJic3KmTHUwng
RGayTm0Nsm3EQ6JI7DqvGtDPL70DPSRqy62OJztmYG7PAGWfye9eSWMDLTK9SNUzNsagQmR1qLRF
Mx1FRoiKJ/m1SXat1zM4zypbonuNn/L2cA8V00ymGxBowM+BQ8jd6TL42B/7XRGWDFu41ySXpPya
shEcMcsucEDUZdY75EOF6cER6TzdwJbd912/RbAXaF23VLqS/ZaqPdvLaww3LrOEqycTmRo12akZ
mvHRjWo/79U98jtKcm4dJS7Lm6g8Zebk04i8WNMBN0BzvfCJfVZXSn67G/whKGwLfWyL8WvprVdA
eMnme3uuF8fyA8q6W9RC/3wDEFOuGEKkTzA9nV/FuiTqDClf9Q2TUajl1XyXg8QYEHnw8fMR5KYC
7KbUoCo4N3OWW5xMkAKbcWwF/pjl6XTXYW80y8s3bgiTpYlIF+hRjMVl+Q6gZDj8Yf/h5nLRFyHz
/0XIew6XERClC4UbvdfOIrcwFf+SaLe8UvYp7Hub2cwkOVDyIN3+g/SD4ilLaa3TsQCZJXUBd8q2
8f75Sv6nIq15vAr+NYQ5qWh73V51lfVMeYF/a1FNchp0RnOdu+ScZy9dZ3HoG1Yc2nT7bL6o8luL
TQXVgs7eBgyChbWGznUcJt49bH6pigYvnuYo+gxsPfiNE5fsj9dIZv+a2zwGKspQOGMqdGlPK5ob
fKc0sHAp6+24aqdUNf3ECbHl6TRXh7oOLqwowZqlqu3rzptnhtt7NTFdfXEo4PqEPWnG5Tu1wlh+
Yqc+EbP7GAmNCYkBdAhrYRXHRAKfoozBdTTfFHBAjaUp0GQC/VFsJZPR8ImmWqEol8gf5xDUY64d
goQt1V75QgdkS4Mh+GiGR/hoWw7nbU+Ayis85db1jBQN0yrrmbpZ30v9FJidLEtXvfrqgIC2nVYB
ft3Ac5S6Mq0ewL5m0AGyTStQy5zbclz4e3T7Ef9J1xworYBoy44+NJbCQnIhiGdemRGpqT3X8U+k
Xu/4hBPU3k6Ve+NTQbY2ZJjMJM8qZQylGMDo4xfZ+1XGGyuJKcAyjS43j9eqGaDUhlTo4zgcPLa4
iWN+xohDya0nW2iKtuhm2FaTMz8ZpNpE+XbHXF9F2rmK6hktaqPCIELW27OcZ/AsvT1wVpz+Lg9B
zQiOMAsA4HDqZUFGurX7Ddu/tRmZm+Jfd0eewIW2R/Q2ZcSQCU2yTtGmsuOeF1tsyv4fgfemZ50q
WmXbtS4xBOR6ITxbveX2sTdphZetRVy2EzX91mkm/WBtBm9WrOkCta2KuQoMJgAbxgW3WcvMqlId
l1J0W7oxftHFRPbl4bkprO6GxTFxxh/KcL0hsiN4yYN8mbuVJSSKOvpKADLTX+JmYSxJBR85dgp6
wtQPO+Flpgn9K4jWJehEa6HQtGsK5sxEixgq4oXYeg8u8Yo4U1K5yXbEymQkbDzZzauUm+waC/ba
Nlbo9aekoMGezZqOlgrcsNhR3KGHWeNAXo1DFgbah7j3UNkCzsLtJ9lXDCU7Zthu+tD358qSlNPQ
6AxGa3QzF6n0srviWsSwkLQwzk3xZgVdi6OwaQj+j3fyzFwHL+Uzcywfcl1FoxmG0Uarn3pb5xw7
KOEeeAOCseLxQoyWopT8PR4hzlt9W2PF8b5qBZmXT6lqpD5ILbvexIiUSxuVeP4nfue55unve95h
lr8RgQrl1NJl8YpAIsb8ZHKqrlekedZfmQqqouv5tjmtzClmdaySDLT8zfjlopqdU0CJaVXZ8tKg
qa/WYJvuIyu8jdykyt7CdBqLn7hyeQqyAdOCazTe6wRImaBRYzXmvcY8xERspZE/EY5gMS//LSpe
cIgvP/db4rCW1w4zBUjTjM3gXNssXqGAXm2f78onf/WBmLBjG2+G+kGWiwWPPeJGYUF1G1an+RHp
CxCqWzBIhzXiRUU3S4GIRIE26u6aih9OK1IoynbZYSVhqjIVy7jCINX/QiZhqNu1vokFLf7wPPvO
X1rMlGV4XeeQ2pzQHLAaNplPg6UfCd3zp7oumFC72Viw5nWSQhBoObjlxOr0c1NgY44+28r8qplc
2w0apDdn5X2I/uhRc25PGxxH+4DRmqXVUKufMHTj5oeutxy8w7yZatAIye7rhm2NLtC3uI3SD6Zb
QQiOaO+O1+H15pheLdPzvR95hgepkeJJhWrGxRCnt10DYaoFp1krnG6XzhRo7P5CEF6Xtm45Bk6x
132k2zzY4TGcAjt4XbCuhlATmqkg6UkKoIJbNRsLGEzmEqeg2ml05mC4bntGLyANHGZzO5HK85CM
/CvLHSIbIgJETEbfSe/c5sWenejggzSQSZtOnOGJzT+fTUtqGrcaBAXyzPzRvwK8ihxY/8fJYnF0
+NP/T+Q9Blz9YBq4fn0pdOWdKFu7SH/BJzSBc0WN/6NasQapoQ2Iv4HsMxJrmOvzBLHUqhmco8fq
Y7ZcIzpkThYosiXjBRKOQrjYGogZrVFwB9VHJ7iKP43DdJ98nPQp+hR99IpSmhvpHOBolJEUAJoo
Phr11L2kg/XE1zeIEQTHKkYUCQH/3V9ahwuWf0Ua4fBq669bvHbPGhxTLl4SFDXRnr6D2y5W+gBM
cG6DLPfNXySoloNQ8/uW5JGX/BcqRu4bDbYpnLQfI9SKN+spmuF6+cghgRmx3HtYkmGwF3HEpivK
qgCqelkiOa4Bud4gPke2SYk7DlJ5Lg0syTDW/EQKUd0ipHmr2EkKX3WHe3ZIAEH1MG0DLkt0ks6q
+7pEu+f/35+D6hi8DGGMs5Qhsp/1nNo3J/MkMllE2kyt/yIPDmnnbwBNQNBnPUIZSEDM83Li27lS
wbYRSMbZgfJmFTdXz+4yvL1ojSMQVIj85qu4gdDXQVbhdei1zn3FLkQPusLUe+kxnTY1gZdFDTZC
CZ9M8IORKJ8o8eiBMNLn36SdIOGl4KlHTxxDbFI54SowXhSgXGGVjTnAeVIDidp6zVDLKNk0zHDn
tcpFQKM0tvn0cXZn8oxDxW7EQ1Yhb/T9yJFlRv3vSbNO/7P6zQW/7QglC5Sv0c3rqFPChPWEXZEJ
Ih5MtcwNzoVg10ATh7MkqO6++dzqjJ6Ex/km43KnzuLTzMg5hVYsg6dwbTEaKkbo/gIsyfk5Ig4m
36ex9TWK+y5Jp39sLvMUVK1Y/7NnrpObwnM60hSAPRPLTmnmy+RYmOKRneIVPhCHs53IlDoLtPbg
6k9NxrxrOD/gfUoEjfldM2p5bwBsewTdUi/VIZWyrh+dQ7r2KFZJzzmyJ1PYZwTgJ05SBf6rqvEw
T1kjbsQv7bF6s8a4zX44sZBvKPJE5NM9TzGKdHQ4RNH6UwZx+lCYiTEDCd8nMdFmQAjJYKTa3xHp
5dunlV5luj3nce48FZpgAGv04Q2dCL9+RpWt9WRbuaq5U89HbGFASw/3b/Y3VGijDqaCK2mpWFr4
fsT9QnWOVcjDL8jQ4yg29evAcD5trlw8JchqUzCdsfoNCnqA1x4m7sKdS3D9qApvbjm28O2U99pG
cOP2jq7jekEXjT1eXI8dU0nT2orVaO30POLG+BKk4kl5NO1jg2tOMjtp/VNI1MdTTbJ+soT6vInJ
AZof1cl6CG1isdilnocyM1F3pfrDyS8tbJ1/Clu+S9ifQCKvGvE1Ru1rzvq95wU0+B8ttSUDQb1S
O43Wz1FgEn3xPsgubXI0Hgs1j8CQAvJuitXQspixWlpQ5H4/NvmRSYIhySKcgZwOT3D1hBkxUz3o
DoOJGZ1c0ZI99pUFV2OnMkRdcoO1PuaZffIn3y/rU8+odJy0/Wy14i9Hb7fO/HpFtH14KieM4XAe
JRSSZTOmFwcGmBHV+0Vik+9wI7XFZPvRhwPPjXiFEich2oLtvEFhloiFOx67tBNDT697A/dCBpom
VDH6QAFzOMkZfJw9jqY6yAZZAaSLGalzcLLlM+z07yahU9xGCEkEcKnjMthdSgOIPZVUOskFf3Bz
ZHufNsVZCatL/zV8GNRCyAyurg5Lt8A+2xHMLbMkxl+HB34hvhofBvCaCZQeCeK9UfFGDTa3GZhj
wrlTtJbo8LK/DskUGTCV+jFMxg+2aFWz8BpRwjNDUohMfVK8AC0hpE96UIS+j3Nhhm8j5DrSLDv/
ZjOt2QwUL2O1/1tkYvdU1DAiJwWo9iDW6WWZH8+MBMDFefrMMXgb4BJKZi3DCFLsJtgkLZlEeexw
ky09uqKfTDJaQTERwYokIuZkxxJHh222eKwWS4mfTuZo6tWOs1tJxlHsaaGPKIapRwR0YSQQw9M5
8xKJP4uoKbuyjB6Xsrqi8vGZn2fn3Ez1Add7jlgXex2M3AtnbAYxUreUQuQW7nbzeE64Y5ILHFJa
BcO7ot9aQsRV0YQ1la/WUqC9psQui9Kr4PshEq+4xNJwp58cq6zX05pa5/Lej9DxA+9CH78gCmsE
W0hKc4cmUdekeo8+/BpfoHYyrJxLk0exFAMiukNeDVMJ/N06nP5CQRXeo/enNCPDJu5PMDPab2XW
eBRLZUmvGsGBtWvd+N4gP4aAVrqgisEX73bAnjlvSDHaG/O0/nBSoOUh0LueYNRNS+Jjavs0MSPq
Uw1Mz2EN15gy61gOvCdXCiVv5U+zOkmT081Wbq/Yquv9PbXaRLNNPqvbrgnItDR6kwqCastKuWlc
B68Ua1ZWHkLKMZgxD8lD9/qr+wv5meRGS+HZLvdJKz/W8XzaZXODJwhNdakIdzrf4jKjdhc0WQgH
8Ly6jZFC3/+h6c5jfVHzk7BfVD/jztEtBgNV4TaFPBRrWBIi09Ovc36j+A2nuksgKZJU/DOfKEn0
Aue5+HVL7owpcfgnx2+cDv1NBmt3csDpm5UVZxcEiDfjV2+3QnBU3qybRCgr+a4Lh7RmmLy/OZ0n
7J/VqtATCFy1Igst5ySrGQvOxTGvRxuOxN8ypUAZyrVe9wiPQZIZN9RSyQtlmo+jxy8AsQaTWmJP
OqQB3wv1j8nhYYYXUHPVyuhH8wq7jgqvcpDF9Z31nq30NPINvE8JFrKXyVpMZW60L3X0mgmK0W+5
yHYRKxwPEeYvhGcs3EqraebQpzGzc4FOtv96D7FlnXPVipeD83dcxwispaVMvJ9UZM6lr5JKg+Nd
B+d/Fwp4xVFaiZL1CE2lVoxsM2aTTM8PL7xg2Wu7vMpfXkYGCixsHHbxJ4Jor0JLMS7tX8TsfXGy
slFMpby+bGm81kGzP2Woqr6N5rWl7TFsimB+E0BWZST3dknIbL31SWYI3/BtYVoxX4+vp1xeeD5t
25kCmYH/93xIkmEMLsFbqg5y2Vm521CNyVZRkCR6URQs9WNRDjAuIoswhx+FH7yxjGS0z/WL5PUb
Gom+nS9xkJzPiWRGDwzAONZ5SOAX9fYh8FdValIYQqjZ89JWwbLId/qsgsTFsquLeD5zEa7FUXfd
jg/d+ZV2eQt1BUKdWJpVs+aMb06JDv3zTYJPYPvMQpY+5BNzLKNgFaFeQTaNxns11YJ9OcM9ZEQr
DXky6HwWn1GJ/fnIRMTtq6BK1Y/LxGizCYXXVspRo0ipfQULmTboY9xV15EHdt/rN+TiX8viiwf0
5aWb3GM4HYJlwQ+DAQCMr2bGon/52tazhuGYsvYlHnSN9OBvWIFAUbkGI2v4K15h7KZH48K49LKg
Q4yc9SGK3nivOgxcNBXqYxSZHdIwtVyTxb+4cfdAZcuTqgYQpijqBVHAVTJf3F91ksx37WjJMLC8
kNE3yG8r5LfxMG11q2Gh9lFF6OgOEzxLlZZ/DgLhWxO7cxlDYZIfUd8Uy4OQdO5OxWkhIW7n0q5j
b4ba7dXvrQaa3zpn/va6iw0Mn4FAuSbcMMOc2BeNgITXamnMejPrbhWlbFWNOiiQSnqeG8YjY04t
nnE8sYmFOv5gHwwobW3mwIm4JRWT+NS55bRtcIMFMYR//nH9a8Ob605phitBXehkY0hxGDQW3mJp
O4B8lm8x/EnN4N+6aJw6wLWWapX/18BHM+i/3FAJEIxHkFu3IAUqQiWMy5H/u1OgddYD9f+1nDl4
62y/ZsQu6Hd7qIT4THLGaAMRFO+XfeLz4ldgfqW62yCl1NGq4drdbG3IqESHCFS7Zun7dtRbbZc8
b0bPdrcOdnZriP7qepuOg5VuoM085urr+EUlDlPkjiPZyhqW031rMMNbrQVvui+LBs+9E1acfSlk
h0r0MBSbEXV4cuTUilzKuUhfId3JuK9yXRoabQzjOUlEkyOoGaGlc8fDvRpkcd9+4HLOfobmScUl
U8p4+ozxQZ5ITupHjIwpjfeaCg99caxStVO69w5iYFs0rLN0Gt51ils3punBzFDjuc5DaxwU8JPJ
CLwxnD4hxJPSADGRAcqhL4VTCL05agHtTIROCsdOwgLAN9UnzWvQL3hlSacjfKRaEWzMAPfBJ1cR
JPjonKHp1bUMysDQlCZN2YkiXLZhfE+6QheTQYsfc7GSG1lXL6e44fDXivxfY510cPDDEcL8Erqq
CqwiR6Mh13NZ8knlbXm587n9QYM+bZHpvcENjEP3R40d/Jh6EhxIfIGuMAeZ5CfmK9bLwyTBT+r0
PsmTqRmj7VAvD1+WahZbeG4i6Nhx3UvrGHNyNN7cgGxFFznB+4lF65Bh9C3gFX2BdfeBhaGUzYXs
MvtCyNpX24mOaPhPVFWhis4OrWbKV+L1skuKb7k3RGV58LLbBJ0uu2LNS0GfUMnMP7sHQWoq5Cpt
qjKjjSwIML4K1PqVqC5lZtI8iGErhe4fgwokWvsZmdpJmt4KuTrRA4AvzOLLfVzOvf5lhIUlC2A2
FMEL/sZPIdmVq51sY9HE/y524soNHYkh8nEnOsBCAhlt7+UhUqE951OKDHiIZWpVBmX1yfKiXZSn
cnqKieX80kMaIj44RFWP/dETGJYBMes/31Lu2qU8OABThwvx3lT26YPnEE+RLTM5787TBgaozd5H
VmUOkKYwgtBQ2CGSAVxvkFOH7vi5Ln3U9AwPAbKbyj0oJ1SXnkpDlYwFuLFPz7hGShalAFb4FFMB
vJPmQXgNBX+Jkb8guqf2D20KGCKKT6tJs7eRWYNXsmwEVhyne2usd5H/189jX+q8Me1MuaUiWXUb
9v2FXmPTj1ovbn1W4xSaZLISNqQcuGEmDOtOUtu/64twB283jjKYgadB3oTRRP+wb2uBEhHVgLIi
PT7jD23s78ViWjoeeY12WDXhQA66Zvro32C6cT1iYGw28zUe8SNFlwsRyaBdG7jwoXTxkwhzVLFb
w5he9+itT+4vo+pGjnUZ9IB+p7YIexRLc9oUdRwqEpKZAmNlVkq41+Ed9s0PYDYO6JjAN7V9wXoK
AQjBZ3gdfPCeBcM1KEeEWMsVmis48dMheT0AT6y4DHvjrmtyXsuRLKh9fAfkfc4hJzM7j/vicQUm
4S/v14WdyGo+Ag6g0dmgUGdh1r2JV+DJPI5q4+xTVrW00Mhc88Pz9teT2WUWiLKtMx/xLx9fQqVM
1klKgVHz37RRImV75f/Rb5n0NFVE/zJOx6pns5eF35dDOpdQERoHmczIKaaFVvYREodCHGc/14/V
KzsQa0TcGyX2R3j71VqKxvFvCjScDat7qP0kyas5eWmeg8dN/pz83c3mXo5ozECwWdVdgmiSPOj9
GVjEqOXbfFUVGNTe0izbK4EDiCOSJapfsKbbYrtVKAOcylTFqso9WcGqR1dy3QY/KgYr/7+6TbY8
xZU3kn+9LjKpWYOJ/k2wxSYTOMLWrGtT4gDAuJf0FNupZYvpRHYtp7qgtQOrh21TMX3FKrg4DGQG
W3bjEl+hnf2qzkwPPzZzmMDUh+dEHhZ4cmOev2u5QZLEN1aWUyV8SPr0w1+3sKgkXGxXQkmCliSO
rAJ9EnavuSG8BEQmuTS6K6sgqx8/mx87pLrutAtKfqHQlRrSVLOYek5EeQD04Rz/3TKUaflJ6k9T
r2mUWsrxg5/ljxResIEW3T6HstAo/+zgjRvAzy15sQciqIW1SF5/SlG2X/bkL8DmVxDn4RbLRWv1
jWdCk3AviOlOrzgt+odFrrn+UO+/SMqUihiEpu3QfsozlKm2L+/kfo4WwIJr9CESgd3N2EnCwZ2E
wwmmEb36WwEanivdfT7ZxElcTPgfrP/T+lwD5/gr5DRTrUh6MaLqprAkGtL9ZFPRcfrOvs3tIt3o
eTDLP0tnDWV0Wkz/d9XBUBqZ7cZVH41+XWlYh4p5btmsiGS8GhDNF+LUzLXQ0YnjAUDv7MpCF4e7
iYaa3QQoZww4O57fcocJ8PlxNlNm2mgcI7w79/Klksqonu6EWZtcdtmB+s4uFCGDXRx91JTax7rc
ghqdTnTbC8LEXfI7SjAjGpLDx7zseOfS5riLbCgBD4kpoK9xKHCdQGhFZQ7PDbWwPelULc2HQkgl
0DjNm+2wrcbga6SBZeVwKRM+9zs443wFWWS6PTKUgefCvAIGoAazkW5tzsNqCahyz8ozogUzGo9L
DwIcV0+WG6eCXOIDXHBpRrR4G/GvViKbWh+xMJ3Dx+uvo4rs9cGMDNx2grEn4BiN2oVWb+M0F9iL
bKfz2gZQWw/aZStVRhJjDZqu44eN5pFNNXBueQVdjc5NV1dipHCtGKQECe5mqkR1Vu1qPvVi8AlC
PUo9b0ftUZsrfZxVAU0fqQh/QU9PVFsxFFK2NJdtYhp8V1pCI5bwVIeCX7eLm1WGPK2RsKggyytN
aX2MHPuKdR9577wWH+cKlQGORnPV57yjM94G0hRyrOpNzx+93TvRvn3/8x/RP1xsMFRQRliBCjb4
B2b017ievUKfjI4yVhfPmYebujlDgOuectqrqiH53C0v9/45vno2I16rmOjRWLdMDNB3KUJPEK0m
4WmSb6XsCbyH52xcjDVr8IC2f5420fhRr9dlPcvlUc2GQ7QRlkfF3mhHEd+gGhrHg/65yzRdRozM
6ZTMUgqznzk9wyoB0//OT+TbUR60Nmv1w4yAaFAayRXfSIc5+8BsykgrvodyfU1WQ5531vZ+9aV5
+TI4kjb7BAf9Eez/FYKF2J0nKrIZgYfIe1AWpQnQ2nYjyICv0sUjAjZkFWiExjguxFV7XmkOezio
L4oSI6SRH5HI5/BDqByJdCSPWpczG4B+MQTpRmNiL1GdVTpjdhBiG7kybjYtrKS90+B4tP17HM1F
IVZ0C7Z5ifuppOf0ZnwAfgAY7P1SKieS0JvpuVkPNsJhAk9BCiTh1liwx1iWylicJyUNexLyRJed
QzuOHSpbnCrML2mzjHZrDaqiRHUyvRPsFQerTFqhX4ULYSzmOvsaxUymqSpdxW2m4FtNR1iUHxnk
j/WVHyP1mOWQSfHCx5hHFhDgoo7RGD7jEsRPtQL42tl6jx0F5xcw4niqJnd0gPKNgkOno5lsCpmg
aWDKPCpXAQtf+3tWqmQcGEZ4febT73Z+11OlI5/df6iKQcBd9d53/J0ijLMfnDOBo6xYqTZSFHSW
CMYFQ1fgURF4lmPz3e2vn7+fR7dXL/IJmgDgW+QnbPMu/Gs/4PqNs2hNjK5HAcuoj1j2qZuWIWpZ
2QWgCl45QC9GOunU2IPWO3xNSFQvcxPjO+zgjMpZMPUlzO7pRZsYgJQAkhS+IeC1Sys58fWYCP9t
X/I+ycPNuQP1WhT+6/lnFLZLTxUGdM7nq/F+MgNLzdt3Dhm/0KTvEBdLL8Fmeqrj43gwrXUu1beB
1nM31hrAigkozu6ENdV83lIhmRcN9zjPpm/o3OMr+lWJUxcRx9APMlCMeJBvAtkQMQox/wVkNNJK
4l22ph5mzZvyclriFtdw9HuX4sBgHAQzUxu/MDUBPsk+XQhFLsYQWaH1uLRR+nzHBiR8rIDxeMb2
LwmWnOgriVLGc/YwKtxpaVhgKtOpm6T+QDw/aq88Uq8b6Kxj3OYyYlb5JNJArG+8paRDJX8JmPhd
gH5tvQLrY6UgdzuyXBsaPDMtt23pgTmxU75klx4LO5PrtUsaU5cUQ/b1tlK9KvrbzQ2pvEiyfpXB
Kg7EWuOSLu+DYjD+2T3MGRFl4z+RgQIq7+kBpJ++7L5yxGU49+hZIA79CwXKO3/jB2jqziqNlFD1
TWggM01vxVa1CUbW3adot3YCw+3m/sB1d3KxYSgIoITzMPjOoXCUq0MXZJTdErDKRzGl3CoEhXgr
YronUuSRpBGAOnLnIypFJdqGeSImXUsRIMsmHprwU7lcmNGCQRxRKM2hFzB6zbXwFRMrcoCrZTYO
KABVHELgj4khOuTxqiIEebDfYfFmeWA476grYPgeiEbefqZdcIWyOoRceTCLBIC+QewtjnLEYnkc
Bjny+Ktio/x0Y05vfQeBqIKofSxT8yHFEYuZqYgEnhzEG6Ui3JHsSMxVPRsQnmovDUOdFtOBuJWp
QvSuFITU92CR99rCbbwuM2r3Cw+1/WjDQ52M4QA82bRmijl/Gg2c7ZHLuDntRORR1/xekP8ms2MC
tkygWoa+22VFcD2uEVrNh0J2BBi6pD1a9KA3/xSC/kk3ZST34DkEPCAaj2o99eHArulVYb3KAsUe
LzgGfA3vxbQjOpTd60hwziNsnZu0H69sxD0WkV+WP546xMYT8jNy7B0PyKAqEV69xybHQ/oQFIyY
eWDn0W9265lDW6CG1SB3WSWdDGEomj2Fch/UhCKF3t8oLtK9Nl5hZB8FRq2R+DZMAMp7pAhKd1Xz
Q93+P4F01g9kKihgcOPfJBu+OMMKyqQ4yFMZK1b+RkIGs2YbyFBm5x2am24X6LsVgZaBB4AiyNHw
SX/4YnPg28sF/XC7evnz8mGVjqMYTpTSnxZUaVVWPw/hJ0LC6dIEepTfFa3NWJI07QTeDKloZoS7
bLQyz6p+uP871yVqpUoewohAE9KjyWlzZXyCN7pPqPeMA+2lVH/J+ObDun4Aoyi3Z5zquN1RYzmB
UJEanEPwXN/zN/2uh+91u/+8+DK4jS8BYy1oTBgrKiC0BD27ZSEs4yYtGJaLTVtw0eZ8XvQO2qNP
UWp7TRR8u5Z7BYltb/8WZ8VvhRDTy0WcKNGnbJw4sYCVpc371Mzzu09Oqc6tm/floZpGjwy7R7vl
xu/A3wggfwKjfILcjT6/z2zcvAEDOPK2oqANukTJItigM/uqyLdWHz7vZ0sVCPM34xaUSr8Jkg51
BfaQYi1Cm+5818ClmEqqrwB2qOf4/+mf4m1i/voBUdppa8JJ9QeLroZxFxySQCfIfY8ZW0P+4+ML
J0rbdXOrYmS/DTbG9lFjppikIeSJb9Noiwu08EniUik1STIlmXid+52zG8Y0QL7M0ckdbpS+mBF0
jMksMKC2zQ3CTAMlbVn4xESXi4QcCMjDEMl1Id0QEXDj2GpKi1bbrJOJ5mM8XwQtLIVyUJiK0Uz+
VLbZrv4FOeqhU+o+YGGhcZfOjSjvX35l1w85shWGojWc5MOIMd55YrZYj5AXRPfS+DuyM2dDeSZx
E95uAxGn8aY+Cq7c2Q9sBiUdpKHi8h5z/X/hesurF0sUew0yyCeywEstdTKS1RmmFyb+gDSG+hxx
JPk18JdEPbvulfrtjeENc3LhyyfrRmHIX3AR7N5m6IH+bsT4GICYCa2xoY8uVIAL/2wTHc7BUorM
kNTHgK2BKHZESap7tD2oIvcX4gB7KbGNKTVyopq5ZUITyGMwk6/a8wBlD1pHGddy08BcCnCPa+FI
VOrz32xfSOvMfLOuA8u7v/o9MsJQfEx9LL0RwxjbkN1jnAaaoVgO4ZfGVi5n8uCQyveEHEgUagFx
iIelmW2xmhSE67hpfNokm5GOlmWv01P3xMrhGO2pueO+gZPRXC+oINzq6yJqYc+OPQzmFKQ4fMhk
4cgL9EwcSS582b27BR/PwdZQbZUiofBAJs2Dj7Vztph09gnYVXL3D7GXjGkatlzlkIDD8i/5emi/
Kgu0pHeFHNeaYG/IuDYBUxPmYMWraiSOrrWQUQubrXeb/3jfUYqzTstm/AIQv9xZPe4G09H0RC9v
ioqrSfsOzL2r8vYE/WTBnU8tD6u16mHh9ntK2T7z+tkuWcrQmv9XJD2baftvHXeKPTBj36vpwMjg
fnvUcIQx3sydx4ZTZipUY3xv9PRyXIAaf4ZR4uHANoKl+84Bu4Avhk3CoM//hoKujcE2gm7+3U1A
/Nn1TuD0ty7/JZIk+8mYNFb8kngu3l3JQrAjmcGrWfW/XFnhOZdQi1gxiu6y2PyjRDsHVLLEUdLU
UcUaIPGTflt57I/w8k2EOpMMrEI1gaEctUXM527YVKAmr+fRJfsfIM2TIYcLFvivelOLrOC2vgJW
dr9aqgswc49saOq6UiNre6hFbZ3xM3TXne8w4XFUqsKoLfha8mC1y2JGJ6XV/xJDpMAIys3PjOTL
WKig6cTXOoTbKo0zkx+UeYTFpMe3IHa5R+S+8OXudRw82BCQ5HnmMjB2rClSDM6Gf0+IfQm2WX9H
ZXNisA45Qsrvh8J9BbgegHNqhy4DFUdVpSK6NP2mpTzUfms2IHUEsHrrmvnWBe/hiTiGynvbT24T
3OmiLuqiTgdp7u2R+U/dyGkjR9I53dTdZhjmLFvZALWGWsOoFgeInohMLbWMcKmChfcq7TH+H/Io
NYUjPjdYz/Xy9K6IzfStV6j6UeHXL+Qxikekr+hnzLt7MtTKVT95t/ZMt5dGj49oo/SqKVna0YXo
5HrxEvI7dpbV0h4dsG9qVAa4h/IVl84OCIf1M0xnIZV786rcSMCcxWXTLHLF/HOiRiR7jTyOP2fl
aJC5juou2qCZrk9XF7egTLs24kWiGq6CwcPdeakDaX793A8B4sYwIraElZsVMvB8rFah+rj0ot8c
uwrB95faAGHjxpDJ0tuIw5lb/a0sg3MffrHAzoDD2joxiD3XYlNsQXXXSueCtL6J1+gsRbuL+hv1
OErlqEyfXH68TlzRn36b2f8WbXiBmTIlcgqKJW4VSpqNc7K6G7pLeItyr5EberY2I70qUo8aN1cn
gfHovFJKJ9iLvDdRVaVJ4mwBIkOzbEQubv1c+xFjDEx3+ZMgT4KRhqypE5zlghWqbuAbS36jn1uE
B+8GVRX2xWUphYjfVrnnpmJodhGsMCh0y0CQw6btqoWGy+DAIbMlLfSnGBqg7Hrm1fTpI2JROaMw
5EWb22ub8SJv9lyGGcRKenh9+hEXflOpLMrSzvHpTcTpQrD8FA1jhnKNssxbCboRs5CspxYQUMep
qTR6SVZ8yaWV++oAcIpW9dItVuGQAedcYpumjol2HViTEYWDkKWTJ+ZgWaFenBKooErH85MFoPHK
XnZI/bUyCgvyjgd3uahaat7qP7Ry+zFncXe36QikRlgi3MjSf6VdMvM1BgYXTnsFdl15MpSipYOl
VtzB+RXlEqdNcyAxdznB6CFc/eJV7ga9Eec4p32mh3tPt6XwCcpbv2YPI9Q9bcEYETQ5rcfuPsZy
DYAAsMrkeoANiFNIRdSzfYh0GgY66aXWB+UeQbQ1nDWMA3zIdM+3SkJU3ZEfaIGML3Hd2qnGql8B
b+9Z0c6kRa078U/yeUPnTK+DZ+epP/FGQ8Pr2iBtSKmqbmWigpM/FIHzTNPygiaNokgrHgtEaCyS
VAFgwCW/FnnxGrUTeXzubt7khpduvrx9XoOYmVXoYHoqWcYgGzYS0N20Y0ReDK0+S9urHxhTJbB4
Til67GZhZItsB5WQjjdK+llF6QBDwuNlBItP4PFkvV2hvvQkDar7S2fnhPYMoRhGp+YZLSekr4gn
IIOii7gt76PtG7ieckKrE1KWYUBVTgh4ZFNNba/KVQ+63l12XweWkb//uZod5A4aQMxjYIcEjn+R
1aZkakfCWWkKeMM/W27boE3sPxHkzCV0FhvYd9DoLmAzeIJ0h+ITv1o62EtsiEl4cIA5PLkFhnwv
jOuQDsdbbbkkPpUs5baoZwnpVvWyusy3rhtP7MoTu8u8s1KVA4et4YS15d1SBRotkb9taJIcNj1G
zIYAqsEsLPblmvBr0SOPoOuFwI5lpS+jq7+s6IvBBlHYTuE6YCMk31TthnRsSMVp6viM8rD2fbUc
E+/fOsJDegoKdAOA0DbI/08OucMKhTwHKXqyd9mWVLPAiY03d7ficFDjlTSf3gSAVPRVySnLPjeo
zex/W5oP5j6+uigR4DLE+sM2vKxvJqVKCIPUMtaCWkefWQyV5in37zCdfM/dXhLGiY7lVABLiB+m
JrBfPY+jwEqZv0LStj6nr01Kz8GksZooWwYFvmOMh5hZQQbbIqJHrmlNXeNhDDtGEmCLcBz2/zNP
gUqZJuxHHUNMflQB6+aXTKxQrBeafEdnnxvkU9lHcPGiCr+9RxQba85edc6j2s/7yHG1qYf4CMFS
R1V2lSZ6TA4Zyg4TuUW6mK7HqHymkYOT0jtkS9x0T6kGHj/vVb2QkXPEwltX66DSUXjN/bJutkuS
/L+t30cWpuaq0lf67VuvvLexWTqyvo86CMqATynjOQzCvSIPK6Iw+mnGJ3E4QXUTO3gTf+AJ/6Zp
JMS+DrAKQun10kr4KfHk/VmeW8TNIcrHsSjUhflK7BVA1FbfGTBJ6JlOOgm+87gr7zq1Y3mtYsOq
df1h8vwggs24JJLIbMmft+Im3khqcaoTeJDgLx5jm3i5T7eOgAk4ey35FRZnhMUfRvUxSJGEanNO
WcJViLd3SNhJ6qej+RxdxS3xYWX1SrhTs++QVPpqJkftvTewkr3HytjIddt1tzPrXLcLIq44lmNH
mJ1J1Th2EkdmBjE2KLe+VZT9fP5EcmM01zVfTq59n8GNqjwzoKTcZ4E3RiKwzvByd36QR18e080Z
Ya7Y/jSxmOFwiFhVdyY65929OeDE5frYBurZM3myYA9ZHEArmyQK7tH0YgljNyQYS+QTjjKrzewF
CNsBOmf5zv2MaZun6XNkSl6mALIwJKxi8Jc0KAohXBdOPYNq4ncFD6JDjb4rWK5TBJS021Z1MR+S
QR/wzbn3GfWugOO8cO2RAcO3a9h2uz9e4ew2VUYwF86oDhIeYUJ8eAxtX8AHGkMmFsGhbBQYNMie
GIZWrwO5QNCxCo0XHjB5LdwAztLke4En3YbHwfb4vxlz985QyOugh8GiPi/ORpSP3ArA7W/rFVwj
Gk5cAb9RO3fHQzBPhjDfr8LqqmO+a27eRsV3yY7d4Q64u2CFDYc03JJOOechxGbRzR+j4miLYsDF
9RUpYJVqGJPqoAlHyn1NEco9QcP7oE7cOFk8Z+VlH9OA8aNDkWR8Fu/TYTrX28OlJIJMLpuGy2XU
iJwrnyIqtf22aGDWgBUUmuPbecmFdUfGxamoN7JZcs4kW5d0UtCZceG+QpVTuxSf6WnXNilp/xw+
26OrB+ioLLGnGOytfrtgKvY6TKGf6AgBlvR+9J3hxca7e+FcrcKBUbwyVXiyijOkEsImYYwWkr0r
cZuMeTh35R5WRg5k1m9ZXGlcC8pWf4MWaWEFjIwWDt5fliZJzeaZB3mKTi2Ul/AZ3Z0nRnAenNtn
+fWkodGWPddkEmF0rGE+lrmEsaYo4Dav6mVxuP69IlShgXLbmgjVMY8ijEF9s5zC6rlHUcPEbF8m
X1mj/ECBA+zAgr0QNm+Jt7WZZeRCbgnz58wEc8aAWHXRPugUL4wP17hPfFnf/Yh0dfiSkCz4f/xI
flr5ZQCbGPzoPppU/synqQrSstcKW2iAChmgtaPcCUTgNJ7Dg+c6xE6+Ql3P0g5eHQCI0ABQHobY
McK22DL4t3fAGyCvbpiJIl+itkoZdFm3AveL1Ud0F9si74L6uAg9epV24I5mnTT2PXpQ8e9UfGrD
3DY5sLgkgMuYxWsQ7TIcAdwuUp6b1tyhfdqORUnKAr2PEsEeTtZn9fBaenqUuQZSf3GzyDYHnhbU
wClxTJ/JIQBNROrJttHXx1G7akA2Yo9grv6AB9X3n/FFvnXQkmJKq1qyZxom2ooPu65dnFf2Vo+g
InWV9fQT9Bj+1QrN613XixasE5fs365Ci/yTNnXfNfUoFWIAFYPzQtzYv5V3m7rkNY9CcfjnFdyc
4Ifr4+VXTYQUw+4Zjo9dtiOQu2E9o+2VvbPRTkiwfQ0d28tOnfSNY6TZXZl4vTfQDYrIjVH/LKEa
50uPsOJglyunsTWPGH8aXuWo4N1V9yAIO3q0LvaglYNQ3eIiT05qHJIz6BDytFkP7ek2loxZb24N
07LrFxff0OovDOiDKGRQv5HWnFypmdJCf2GpOZcy8BqeopzJ8+Xyy4cKhbloYFq6brjHVtFLPydg
uQCEqEufCe2WPqZw82/bNY1/khPlhALkv/Q/P9gJYmMj9U88G8IO4wcoChscMOHqDywZJbFSJ1p8
9T6eBIMVn84kIM4kGr13YpkZPsyBxjB/4+JHYMCWX+/ROljGfTBKJc6zjOK7FSzi7iX6WRCYwKIB
uLrtBKuQjQcp4LfSmzWR+BnHwm0RdgOfTdTfGsSLH+hb3HlN0l0csXpAN/e8bIu/5ktnRoI/ef0q
w4ueYQ1osB+s92j54zD6dTJ/b3hFi3idvDqf5bLHBk5jS0FWSa1xJivvbDQpROlU6qJD/s+xOUDr
57VzGLiSTwlKUR/MrRac7eZguvThljGlOBGcvztdTjyxluCIB6jSsdMGA4bfjHBQAWFvAV0cMYmR
zI59P2YlDDgHEzT/hWvPWGiYoQxjEf6An+ZJN7cLelJHNJas93vENlFjJzA2K7gVGAffoFpF4oKh
8UMRKP19bJHB8N8M3btb/mb7LqxIaFbLBuH5SPqcc5dtxucu6/8omNdL1L7X4YuFpv2xqb4D33R+
YWT1RO2nMzK2Mzrufplx3JvbmsgPqq3uX+rWyiHwwNfO0uM3w8Naty7Ez67jQRFwbQ0AYP0Fyo/D
NdDDGidHAw12xuZad0aM8Ad5qhXBPCsLx+eJVMbX+AVCKbBI/rXPBKyPDvtRto6SBOYBhTCcXd4x
LlgF58AujzP4S8bvgufa7zD4OdAKe1xi60qsc94lAJou/ajuK2FSzl5IVWuKgWQRxXvXrYZX/Sw9
yPT6hMucsjaF5sv0D+7K1fPlikpi0VXb3lH6WFr3T364/VhpUrODAkgiuILY5rAgm/cd0OzEO8/2
Wga9niJaRSHPhhKhyr+iYUiwxmcxDZV7CHC258t7wh/euVJTW60eGc3UcF4dnaiGTVCH06NX+Fgu
t2gZ5MjiulTUWsHO7SL5ssZF6FmcmVon+HWevME9nTZMLrpThGX95CYpSlICyJEdkobAYBgalDiO
tyKqrgGr5dJm7LaOPuDQEtbr+gUcH+tSMcGmObGKKfWig69CU91G3+2yxxyKmxHNmhh4PcUD9Q08
kvahacSnQ5d7aBMJvjHex1sl26ooSWHp/3jVffXJqd7sj72waz0jt3mZQGFvSiEc3KedrpdBbjWA
OKCI06lj2bQQCvGT5AkoGees7wO+AayCfIaqQFyrTIL2wFhevo5KV17ThK8jNrdTCR69o8cR7oMU
n8JZ6YnKw4aLyK2rj97wXCHbk/4ZLIxCqVKHOEzCeFdxwMS1sKyqHu9F4y2hBxeXUP6qQIc4IZu6
sNkMWExnufES3ZZ2rerC2Y1YozcHP329iewn0k2LW+g5wKbLH9eiXLPADeEnqJNiUOZLKNcOv/HR
G1trNTFS+PjyNLKzB5k9qYRuibBCE4TU/jsHWk1q4KdsaavQvEuR87uY8wNnvyxfZklmh37iPWkf
HDUbWJhrq4bGHa2krnGQdx8SVu+gWAXjOucKWNbWMQ/CS76bDXesRpIRwb8chYeRQji4b/MWXWKs
QO2kLR1K3oklyYt2ZWCWswxS+rrkIT5MSjJgdb01u4KyY7mBd1pp1UBcT4/lUdgS0ziRX01n9Fph
ZoMm8iR6a3KKcFyIY0rdTdBe/GOB7e59Uf1MlizM22x+UIkkpangi0yAPV9lppD7P7SQCpBKDWVP
LEEkqgFCNgoTRVcLseoB6U87mjwBkmBqDAe9cRUhz6g6jTwvUGA5A6Kqc+raQK7LSNwFDDFA1Yq6
e40Y3qRjlCs2Oduv0t3dby+8MqGI+wU4OIzZZY11Yej4lggp+zaF2KJ8vsmzonuRXYc34rBKSjDN
JKpeakKLAU4MGDQJFTnqCf38Y5FJX5ajBOpj1GxyKB7PktA7yOIfStvJa987an5hGUkVbs0fFlA1
JKf4KxKs0hcM49EK0FSWmUCTauKVNz7/jjojQdSH1mnIWtopATRmvAjqCJf8sL37hd78ykyAHXer
CGd6XyaLQ45zNzzYMXdUlmys/QpE2YQfBT13xCDVRrJMsMB7toYxlMnusxBAXDxe+HPgVvgx1GTZ
Qt577BSOPn2aeG6SROJnv27wQrHDpQeEPyD1xE/iDE9kHpEydQ6xT5AZeGih9F37KdKQo8XHNcXr
0jFg3zV71L39DZkTO2Gf7/sI1WJk2arNmpZAtc95C3MK2QvMtCGP/xbtE5sUeETQdm9rcLGLecXF
lqDp58jMSm82n8UUxWk1VCfgYlvKq37rh1PlY8eQJWkbdYEdH90iLvjAkTvXSwifdKsnDol7xmEM
h4aoj3YNrvOCuQUxfa+VenvIPwzPYQFizaQ90B3GeZSW4XLnBEAqCoJlpbshv1SUJiouGZlmkzeA
dNaD9EkH4F3Nd7eF4QGnEljfhXtdBnUE1AtSpYWnCde1xjQOV1ehtAftfOmbmn3YM0uDxqHL17Fr
xGFaHatk1zd9vtfgv0fb9IrXX/Fljf0jwRfO42qhvtlqgBIvMDsySgoMBqKsyJZz3mShUSht8FY1
755VXzhnpytbz/tb9mknhJ/rbuahgg8fEjSjSwFLMbXmQKXjPKiF5BfEifvBrdJ18/25CDDpajD4
xRV2XwGHax3UQ4ifh89Uc/0dyuPGT5RMqt7oAo+BisbR1KCnVrdzkilHZJfeRQKrUugmOxfHuRSZ
fkz5+PVRVkkXJPo5DYOuumqASAWAdqjO/hOQJnylaVf/p3bC6ZXmgH9KXYvEx5HRE9oLZdRr6gL5
a4Wz6YPH63jWlbzPptlrhiD64fbr2qNsX4LOasbCi3FI4RO1FGLg7CRCcVVkDcggBcVdvVOTA2cz
OTjq5BJcy20Y/BPJ9PPNImZWQXQuX1YAJPmoZ+j2d3eUGb40un2IS76E3/WNOhquVb9AJwZlfOn/
mZeWnZV2rYgKhaI1JGkixtq4hapjIpaReKASmzlEFlMGNI9xqDDFlIfeWWg7N1O6nwMF/LlO0khE
u5NwTigqj5IsVGqTWOo4m3Hjmeuj/iEEvxyEqhJIYpgsgXosgFag0p2lXQS8YsX2KKwdwKgjthrB
87seEW9Pe4D2H4RkoqRPs6BKQSdzcUm6B4M0jUZVf0p/cmaihSRDMLGEoqrNeI/q/7agfF3ri5Pq
ZmoUEK7SHITzFRKfL4SPEsfxkv1GqNthRmde7aSPUFxE+Xn1xrufckXRHP4KXUmppQ0cayi0yNOm
cVmFLe0ms4atEgWiWMdufRH4bUfXZA/T6Zqnk/2ziJEQ8taXeVJ5ngX1hWPnFzoMJC+C6Hg/QqgI
LpZ7BWlclMQnPuyJrCAQOvUt+h7d7n9Rxi+MBSWNr0yQGwJJwXbsWtJHRgmcYks14cK99SFpc57W
Prt93sMWDztoqC6O1JkEEPvIf6YhuwaZlssYZFRr7vExQOSqK6GwpZJDYJMTOKDBDjS73FMzy+6P
KZVDq1DNNtbsK1hNvmo2Jshyv6G123iUgTaBh8bTQJwmk91/2/1sEHAF/5oKuc6iVTilejoucP0M
o2olNP7zHBaPVU3B/R+eqdIpzej8K6waOUrn0E1Lf9iNGbh6wT/KjNswj+VbqeyfYrD+Fq/Q/S5K
P+PpG4r7cWDD3Rj5AZnqdJ51sinylOauwAYhPCSB9igtTkk3ZNrSZaIWY7ZIA7LRfEf6rhjs7wyX
IOiqTlYyJx4miemwbBh2plE3mRuM3JA3HB4vb7PxUolVhcwpNg+c/YutqdoO0RYJSLy6ZwfQADHK
3qlI2DW74l3AReR2ctpRu/Bo4rfzkvTdq500/XvCd7eW4EMfFFHPz3JJoj2aG0rtcYEee6lLqBn/
1fI8fja4oCj9lLEooVP76UatyC1VSF3hlPwt5yaHki4bfoNslN35W5n5GYxIXL+l7KUVypGA3mdG
HeuIBmMqmNBjRp0MuAQUcBfgyUdfmnG6FS+VDlEfGZJrKVWcusaNN8d80w5TFg8EE+iQ97b3UCIK
wcI58ALBo5gytMNFquU15ovk8tpI8lgYiMTw5cjE5PNph2DwQhWlQYfm+4iXPojip/ugrDUho2AD
E2gqd2g9b8htnRcsW40/zgEPBhANnWutpOpWOEUX/Tbqefmh+7X/bJ9Tgrqi0coDa88K1kHDq6R5
4KkHRUBaT1q4zeNL0GvQhdlyPS0Q4c6r97k/J9tArNqamdOGp77H4CovASDDBpqybKG0zgCGRfNo
4g3sfzaM1J1IdHG+xEASeI7nwzPOr/f9BLd8q3rH/u+ffVtPI7f23r1IRasco/n0Bu4bhr+UmpB7
SQjcFRrRZuI20E/fkFKEx9tBha/KQ5WAu1lHwTP7vH0kOaz5CdciLWvymVqj1QCGDcJFfeGtgKlB
s/0DhbIkUopYCmdgXudZH8nIjZUj0VK2t/W8N5BEPIURtz5Z+IPVhB8PhO0hoYUZFaK+FtPV13Ub
QgxeuK4n5GpHWxJw7ldrmKmTeLtpCT/MjwmRaudjE1cOj05wHjdPkwbX/X/gwm8y86ifXzIrNJ8F
BlyK3yQjVhIg4WYJS5VmCkBJ8Tal+4WfaORUyexJTA5JU0vU8WW4e3EVBVTrOSeIbdAX7iL4BTkA
j5Yr1SbdgbdOR9DtUdKfZwZuwgFQMtqN+CKIod/4/GUzjTWaT2E4VvAfQ/d/qiWkOLK7GJpK+dfz
LN6N9RyHYfvX2j/W6lFpIWSHhnhNXf4Yujgz4+OBWqnt45sN6QG0VMeZUWTTPtFtAPOFE63kGKtS
8f5fPNsXS9Pi9dSPdSVDNVAWI8brG8kiabq7Fjwxb+YEQ6hvVKtWLm7RExEyUjEmVsLxKuHnGpHO
7ojAPr/5LifJg55YCQ3JxnMpebOUfAFwMZHV1WTkS9mgn8cS+Ytns6nfyXq/4Dry+528n0hQGFHN
KRGF6ldoNIIYs8nxd05zcruUw2+avqpibuYMsCSgYHPl3g6vXJccVx67EnXlzCA4acu8fmJaNOVt
hjVgvZopjJGrfyOsoHiGoJjLakpJydapAvOA24ETnFToxRzGAfmNy3p+C3+fr3TT29I55l9yBgEm
3zfmvsZwU9Y0knTeWXVkmtWZocGk5V9pjmZeicgfWq9pmjCCarhnkuftEQ101Y+ezW64LBdU8UNP
wDQy58G8jSk3vKMth4QczTYnUXEI/8PdEmc3A/+/KvN+DyzYMyniOZOv7xuolAFZtZ5dzMQQdtf6
Kwkcpm889uZzeMcsRzX+4RqqhJKlkon9vuGr5RcR0KJt8bAUTZ3/xXNspoVGT+dg6MntM8+zcxPH
rST6ksGJo/ejBW8OHbvjssNxIfnnOxnCqNP0nd3khNkxTgDHoCyOggnVZ+rT3D2HkQ+FSMshQc22
gYzWRQvWmMMqpoakAUK2DYe/ojQYzL2zoHKeBH0hrDCJwRCgbh4sviI+0MCIPU2MuTeD11PFWJLd
14+eixfR0GGxnVzWhlUcWLfQLhMjtbuJfe3By47nKwVvpyZ5t7wUsIuqjnWv7x+Lak93Ee9PpQTK
ELEKXXhb58cGqo9rfUsIoWjc9+2w7pcWyLVI1RJY9bF/Bp4P4W20IH9OiylMyiWGhB6aO1g3buYl
ZFk900+vZCSt2ZQAGBJrEtfXY3jWV/IxdfRSczg3eAJalITYVhsCmxuMQ/PYvU7UJTasUYNBKw+6
98sun3ZzzqNR4dSKGFkvl4Vd0fo7oS7kl8D7kDWiqZimfnqYRdhTbQcjfeAmc4Y1v7OcWs+FGCyQ
dlxiKmzls4zajhcV9iVDHXQ26dHmelk1kA32kcpHwsCHau43fIqGJgwkMLvBom4IPEgBVx9DfG9O
fin0uOY1Ik20TBZ6HuryCIwg//Y3hM6Yi5ahXVy3tTCgk/w/L5kcRzAMxnmYmUlaCHhfvIjDEf3Q
EmgxVtkbREfMfrVrRplgiuy971h53Xc6CLP1wM4LniV1NtUjy8H3R2xlEzZSj3tODSF6ojbyhz7f
Mwr79AY1MBn7N/l8D+XSukYr8UOEwKfy3KHpMn6sImgOD+LWn2lNWjQJTFKhSs+2oT9e5QkWLTyl
DDX//Jd0JJGtgugkfUdCTsznpHOsmlZM1Zwcc6ThdaDaalxE+g/pX73idcUvK+QGjRcKUFUoSGfT
AW8bNUiwvnTEHSAiASPeO6hDj07cud0i4v6glDEcln/o1IM1s3cIRTQ323+sYo2JwFqKR2uXGQjZ
s7nxWBd+ZJdYhkKYtRrSxMHzcjjEBjNkKg2VrUc4FJNUuhpvkKpJhkVdNdYY2LFwjTLxWN3DeKif
uZn9DDYHA46zZ1Qm6cBvDiefu5JYGD/YsZJBcH30bmyX22zyqx+N/Ar8C7ggfEmC9RvqzP+JHw7Z
8tcDu+loO4wd9FU7MmfzXu/HHUp3FG3vvqj0IpDpcvQ8IcFlZhIID3J4McZQL3zoxRYSWtxYtBWt
nYj9pIQGZ4SQE+pMo7yzUDfb2sZlLBBT60AdMvDRSCEPeaHGwx8uRz4i2pDldGdwOAYtGoqXARsG
8Jz4vb1J3SAjFY42KrTtPbrYnNiFSPjzGd3v9t/c8dqJXPJ7kQk3lrqXOs409NLITLuWl+HxyVhZ
8wtiXBrQP4yzguFmUgJ2HXbiAVKTtpoUa6jwziLhEBa7bHMEibte1pZfy33u4Xjgeu7f8BUlkUCi
BDTlAQRnrgzbZmbT3qhwCWYnMlQdGaj/71HTKKjD2Q4i8vey5Ubi760XOLyE5SPykCVsn5HvuY1b
49lxRLI736fNcb7ZmZNLl1R7KEXFVMc2oGaGgaSEsVPFucYlNPc7XUnBPXdS0Cm1bHMww/381zi0
fvBzPVAMizhz/nS6YKrHfaTXz3eGulJfBGAR615/u4WhYKxLFIaRKAL+p+IMiRnDh6ufkHb7foHs
msJ/d2JVjNvzzXyGXmmoweUpXBNL1pTJyiddtZQ2Zsp4WR37B7TPN8Tal+yxjqIuulI37cn2Edka
xZsVxuouUTUbkQ+DIpCRPtUpUJ+Qlncx/nlPVWNQYIUgl1ly0iZdrO/frq0IA4v4Bs7bNQfk1bZc
RZhZpYBwVWY+iaOsQXBu2ZmGFKdlzJQaNstRaHQhS4RtGQPtzFtwqLexDqoaCouc+nS6ezi0IbmL
lnewpenpy2b5FDTgDh5JHWgYGk+qzcuIq9QkLFxxWkrrBK7bHYa38a7XRPxaQ+DZuSOcToU7ucg1
ryabb9biusF7NLP945Mp5XztAAKc/mzlLxpnNRmk+NtCawTBsqFc2BtgyRUOfJuh6r6slFcg074P
raU4maJl5gPj/7tMi83Dn1lF8u28urH1vmIEhcF/SzINx721KLnb3pt0PhePJbx5hJ4jwKiYRqpk
2lQh0JrpnnlGD0Hj+lcAm6nLflY9aspYBxUqSpGzAK+j4Yi/K5lLcZtJ7+H7EvG5PerMQOhp6D60
SJQH+ymvZynnG6vRQmnKuzvM2L8BZsSRXuh8K2THCKUiYn89yXHz4ukqmaQceSjcKXuRHFz5+l6D
EVhrOlTmKui6g/QKFOqQ+z5XbDQyC22V7Hi8pmYFaDgcc6VmGOh5N6+ktrWqquXz4S+2aDibXCAS
Fk1ErVm/dR0x0FCVYpAEEANn3Q+cConlXYUE2Nj18c3JuYfE0mwpiPmYaHzBint71/BSTRiD2sSx
yBMRPKBZOMJgULzoVq7aHwmYHVjDsqRRhHM2JJOOLRYnk9qx2Zmx0qTBHhq0c+lwtz8u4m2t0EiZ
/ZswThuRaAdRwpymcTmPILEYmqgx2vhuGypxClAhhs6AWQ9TXdpHORNc/Oru66XtSUBe8jkWHsoE
XaV3lJfRq05II2kPr/R6FBU1HYkknbFpOGMUFtVjz1AVUBL+Kq/6lRaQA2gLsjgRKBE1iPWfNZ5F
j47C9tY8qzFtNQBLHCEoWeUYzdFCE9lCHN2MgbE/6Vb61ATw3xrxvLr8d3E2pMbIw/FtWorjm3u0
kSanq+gZo0CtpnC+Bar63ZW+ty5/4TBkqB5DUJhSEeg2yoad3agii+3wVQEIqO17uzqygyShcWRW
hTGfIpN2bd+VHc4gR03jeYZn7JbSqYasGl39tO9H3+jXekTyi+M3v4+TxEgHehUudtwfgrsXglRN
gVl15rgem7mpXhlQAeOd8J6DKtMkIdB/koKYQc0opEdPZOgvlp/xmXs1uArHckFssvp4ji4rB2MD
Ga38ma6oZJaXE7wrSqfG919Z0HtsHM3OzatITvk8vUA3m0oaeYRoe/RtJXsySgr8AOF5ruzGb2X5
ybeWtP5rhOkCxrBKatTWVN2YFetUg/HS5e74lHf0YkoaBkgJSGVphjJm1LUbM1+51etpXKxSphJ3
c8vsD7A3d/O8t0+b1vPvBzSjzVzPxqPV0H0/I/jW50E1KCsirfBVK9p1S8/IR1olqz1l06lk7Q1O
EsKqygPm2CGw4OmCStrB9eqtmg7+vk4aNjSusH+fDu+rPnuwGJjePlDsUUgiD0pT26gXmpFngnbq
VosVPuyeO/aEuuikdHIFVwpEDbsJKsjotNv4Jc5syEByb7hxhlFc2V+U/jKLdLZOgu8sfIR1W62w
XMcdKY5qeL1l5oYseAv5OhD3LlfuaYrDRGt3VnsQUNApENfgnB4P79Zmre/CsSz6sJQpQWa4FZcE
88Pk9VWOoVmUXqbwWMRzWWR1Cfr8t07FdbmHNnq7Y2/q91BnPozFP3SRd4X8CKRaeweUfdUtgJ+3
UEpdIfEmivGpnWsfF6OIoeT0tSatdq5/E6Jey8AowCN/KSeQ5KiBoyS7yTm0T5vwtJuxobbbdCOz
EI5mVdVxVAxEPGqJcB3nFnXezceO2SgOibUKZa6tsLg+aYytuDwd6DePGiM4T95vp6ONDIIKtEpo
RKVkbvc3q0JTS8PbDvVEkoqJ98WdQPY7ltWbJCnr9OGc2DiaAVJJ6knV+EdEOhLxIACCg8E2YYYr
TL5c8llL55Ksg/jgppgSAMeGuR7kSlvxIYRzn7/2NQwCmBJbl4wXLR0pvLOq2eTS9ioWS8Xjyb+9
/JmcYISM4si/7UBFjXnnXO4h1rZkzeq0piV9YSngaPUg6gag62Gx/w0jiinp9ywQzzQJqNVBL/jv
yhBCReanLfQWrRScMDn47U9JwdWV0jN8uYmeUEm3EgUZlbohcLTs1CKbQGv+e487/0kOkNGfaljj
7nzXZFmKlOdtLCldVDcNY2M0EIXKFz8n61jEcWSuw4Qvf/bcgrdsoLAvp2eutDnwaYW9E+abyLKc
v7l+RHGKbobM+GbuVphUWMyw0fBM28wTnvZF6iUXFCyPOVvvqYWmssPVXkwpvHFJnFqocMoQXwcH
+T/WGqAbmRmPCEP1ByirPYooK5CmkpL3OyfRYIyirmjW7srtRltg88/1utlNMuT1W/HW4nJ8/xp0
XKRzoxqlnxOxKsgPYpnjMOw/273vOEBmgvM4EhSjgxRFmJa1jrmZDahQPMHytSLGKw1jqshitJ2l
7XoQoxVWb1thiypTxuu8tWomZyMWfmW9lSrWVZgMgL+JmMucILunIMU0PdnSOrDIkyh9Yx+31Mx/
YuShIOvmEccO33R/XLnmVNAWmMf1weHVnR9pCUx3M9QECA0T5JSzx3M9USnX5ABcqhhcJRTd//Yv
RYEuZMzDUYT0Brjt+/t+9FDFBzsy18WmcwUOMOVC1TnJMn93PB2o3aa6VPMnPR6wsfRxyWOe4c9g
LzajOOve9xg+0uUG7UCmgUMJQAe5pEsczFcjXbCw3w7633e7TcQD2UKuZiI3H4Q7bXCwKe3Ln76h
c2hF1UnMMPYgbP8o+j+H4X+0WpVGdufSGM5amhtmRmIQ0rBFrxhLQDLZFSFtg/gDQy4UYA+vYIB5
f8huqqcEroA4bJsSlODQrQPdlCnnO/HGefD/IJfmnjBor0Tnjx92vTLwluruOqcYcxChrCyWIggo
LsHLT31FRz4UQ3ofznJBo0a4D+GymhQHJIV4/Ltyy9XpQ+dp28s5Rgvl42sqgbSuTmopI2KdY/bb
k4EAeZmFDNJu2zdbEJSTWqY3HzSsy8l2LD8LkDn+8lnoIuDZd/4XC/wn8aj2rAeQSLTXjfed7dZw
uRlvSi3Sx8/pF+ZLBLovu6P/6jtLp9nbw3Fn5BWUWcQJjvR+w/ZTBckY7YX6a0siL3VnDoVEmeMN
oeMJegpOs3VJvk8nWpV/qYGFF0dQQ6T2DB5GuQdLysjAup1BVyQ8q0x5y7nqHNzdmM89r7WIRreG
7op4vhqDIA06frpydukN45amQ5YokuX2uKmTDh8lRLEisGIONC7gzhHW3TLnsywRipAsOk74USn5
Y0Y77GuDaWDFs9KARP8tuIBgjAP9H0BWzR0hjSDk4rJlZtUl85fTHscjqSxXF1AjyKOGqhIqhMdx
gqBncy3fcSrSP7gdWAkshuYLa13iyVg/V5JenTtAo3c4Q2NSla+Mkv0EJXCVNi8j/3JSWOHdGP00
HDL4BHWyYvqkB7qVm1dVLAkj/0z+GY23MNhaGFFjrgk+SST0Lbdv1Ch8adLG5G1XvduIKnKC4aIB
5ghKiRM3O4WEhF7E3RkkN5ZMXPLRgOymPE/RLwtFQyxvFJVwRiptXAVLlCOJdZYn6yOfG7dnpz1o
5+r7Up7U1NZejQAWR0Z8mnEqaQPmzHjCuAvZwZhSZNHn1ck0KUt0uurS5SZIAhiq/VUZuLz9zv/L
qMR8wnpBtiMZEOrSlV7e2mORZrNy75SU7x/1nKOXKsKQcbqwcGyIso/j1+ez6eN4zPQ/mg/pyQjt
O7SEwSKBR0F0mCvDpJlJWLO0mFPQRH2gspk8vrOuT8OGDku8Tw6StCtPaSn8fNsWJALX1HUR+ukk
U+GnJx8o8FTA07JmAGfmtXVHtn5QTOnjhVc7lhYMeNIk9bKHej2QyrsG7d2SOE32n0paKnfSpmAs
0y4ppe095Dx4oEQcLrRN9AAozVSz9fqKwtkKxKBCOauslPXy/guRwgBE3ZhgMwePah3NBHGZxrwP
sO5UVyX5G9fe+t3FkPrNxvEVYu+2h1A821y8QDsctc2ouRbKPKssRj75ZuXuh/QImZ5Til+qf6I3
l2Qf3EOmJwZqFCzx2zU1UlxmydLJyvAGs0VuIcU7uzsuQPIEPjq6BTLwIG22aAT6z0MGTydaR3xL
A1yQSerOGaImOH8XKxX1mNOCNMYF+UxusinrP60X2Rif6IEt2GzKtJKZXnr8TjdZaeThLUjemcmq
EwQS7G6uvhbkcsAvpn5cBgGAkZUcsV1C3K14pO4LZMDKaW2ytOgVq2L4E4cBTxpr8lzdhFTFX08d
uTNAOQl7P7L+jGOsKiXjJfQHd0ogpRoLjWiEq3md5keWy4dFI2apvwuqoKH4dYghhxhXtckFuLPc
Smh1ZnFlYTALSBFKsrG/e4XWLwnkXocbbO6JmQvalqxorMM8Gmyh85wJEw8V2Jo1JAZK1rWl3Kc1
3kraYGaqlms807haugjRsg5dGJCtC8Ca5L1GBLIoTXIlQYaVPOUpoIQR5qCrzyCrcUY7bfVZ3Wcp
y9raURMFp5AdWV2yDYlBwxr0I96PoN4JmV3cplnAYPdOyWM4XTOiVlKdZny0UfbpYgSgO71BOqlz
Q9k6YRtMMMFqovdqnKEWpaJAD5Aa36WT9M0wo4KnEo9LrnlaegKXnoeT2WDxYr8CNZ4T4U9Qppaf
9FRPyxzIbtkPKUk2zYZsKMeL2J5QmBJ2CwUjp8+6rsQ2C3pw7Wgtg34bN9H0KwGZ2uViA+rKaFW9
bNQ+6LsEd/zLDU1syUaO6vhrgEyDRsRNNqPDKJpMixKxz+AJnjthnx9oSkhVn+gsP28uYgeYRS0A
smqpXYJFTP+YjLgwW5hYqFej+xCqMSZWEsWLbk8HXU1yLr4OZFr/ngRLXlbRdHEEnmRxr1+HA9yB
sjxgdA/anu0NhBTPKPd6W4Sk6tnE8u7ZI5abQME1+fLtjFc9rk7pK4/Q/+xSMf4JouVXHaYrqu/C
8chgMACRNDJylXNys+IXGBXYThmXCA+vBqMkY1atg4lMxHt2ejT2nuGGqY0bT8UvcMM5FBTdtvRQ
9G2Z3NgzOEusGuMvVntnDysITt9gtRyCSdWji8VzO96twSAUWtduhyaJKHAOiWO6EcVRt2JVeNaE
+38ymy2R21u/iKFt0xbyakaEip/CZ5UqWw6vFCdQxZzfq8tplVBxY8BkMHdpMFOL8NKUPo7BSy38
bBOampQItrjDdqUnKYQRcIX4NEZVDqCqm6GByZZyLS3mv5xypt5IDmzy8QcKRdRvy2De4wz54szV
lIxq3gbTY8lnAemS8U4KbKMNVmqj47A6flrcxq5HmG6zLR+bIFeFmstvIaJjoZsku4H+FMnyUCj8
SCDjxnY49cZDKd2wU6XzpQDBgwSaVFBuUYuWItxnS7+Vs5ULlMiy37FDqKJrw5mlQVDJRRXILA6y
vGSUSVFva2OgRKuTN6kmDLHy00X5gvP/LSCAOUp/uszRC6/0tbU0ueeTcls6F2gfSyDW1bMFzIk8
KnmfHuCeHjR9MZaWcyHbgAhZv2MNrGUkUrI32RsqjevVwE6icQfU0DF9qS0a92v5Uisgvb6F+Bsu
PFPszb1QJ+puBAplRiGhGPEehSBa26T4hOD3hlznFbcOTKzoutWhZN6S5Lor7OyoE5H3BZYtkgZ0
r2xS4DbL/gwaO+21vJrpUbFxGIPW3ikf9TW8dbg6hcqi/i39c5ePZdZztCFo4xZDVqoet5uYaDXW
FR0GBsZSFLGCDkxMBV78tbqn4Dq8DcEU9qFYliKPZfBrhoNxmlozfZ4Y27sBQhVX96GS3XKHs2pI
ivX/Q57c4ZN7bRiRqLYq0zkkVXf7k/8I3hMi+fnkhTlUrVJB+Aq8EfbkYg/G4A69eXFQFUWF+ntB
ncXsJwi405b6qB4O4RlJvAZx2maxlH7UAP5zjPO6l1dMlODLn65ZbDqG+1/JGOkBEoHU4Q8zEhqc
Yav5zEuDsExoB0Qt9+q0Q0iRT6Hi7c4/ZHTJak5ihg+byLuF/i76nL16T+Aam7sX9WWj3bBAMomV
aqhW1RGZj3v0oi0X91eDY2hsA3VyycJKnYSqVkdJlWmHexlKLOzkvkF5FMlTJWNnWXX97cDHGDvL
XSgU/5rt6afm9e/cORRxYFwjXgt+mJXhK2osLsYVVWHRtMe9effOi+7gJ98yplexL1UfxJJg7kl2
xgO9ZB+TERsIV6Sv4fRgm2Ly7trforgxH8e1M6jtj4Jes/ON1gVW0c16UhpGMlzuQgF2Rwv5o9T3
HTmcPdBtdX8U1koUGOsZyR0fw2w98IB0LhFjzQe6drEIDDcOM+OfKecyXpi4d4W6zX1I3daINgjh
qFxdar/I4bj1vRL4D+IPVrjuBRQFCACN+HpMz7+blI9nPwZp7P2+nwJeq0uxe7fYGCZHBfQzbz2c
D0XXkJTSsGoOzhPXdVkR+edUQSQPunTWgRtwe/kwYIvl1TkDGxcv7v2B5mVn7Y2zZCgN5MT5i6a3
WdPhLutplAGeQAU6RY+ve3vPW0C0ak0j9NbgkNOJB6e6u8pBDy5Fh9U2nH8lQeUlGz0axp4XPKUM
z3yh9Q0wZIC6IJUYxY2m1+qgaKm1Nsmu3VJh6IYTvtAdmAo3uNHDEc3MAdDNhwNkKYIyg3zrNFMi
06VQohd61HthYtk7s0PiEBGSVHwtZMK23VWp4Fb1CMleQbrYBxuyA7zBaLG1m1jFHhd3WswR76GG
lePcL+wwdLcM6ajAX7eGQqArKReFUgryCDGLkNOGqRxcEXQ3NtgKN1Iact1KU1lkLnXLpzoFavjH
d3W9s+M0yoMIIkIHmqfsCyY7vav0A62XD7y2ua1KCeQazwW0OHkvnzNikkwX5FXpUqtWgCWikGf4
RNS8U4dRGImKLl5cPrudsmdMf+jHI4rwSYHITjoOfK7xdt9+oxtR5BHvZ7cMRhCVUNpwORzKUckN
9pzB7TphmxnKdb318q3WX6p7Ey8L4R1CjSrUVmf/sjvtfekqjNXaNNQZmXMYT2caRaFRLqqNoehG
wZ9Qy0oe8ptuRiH81vWrQhdo6SOKT4DVX3u44xAMH4+SNktaP/8sqLX0T9Wci2mCjefvdIoMPBUS
Jd1cgJqP4ZnppDn4PcjgJ3ChS7GaN5Peq8pa57ONAcftY+j1NtsRkx4DoT5XsXr8YEBf9dQXmesM
g42WbMxASsCFqy70Qw+Fh84mI2HPuepfRAzfA0MILpjtR9ss15Pfv/869sRlzVA7i8JkT3nvfXDt
MEUYLVzZjSM6Wq2Yuf7/zLlz8xG3G8AJTdFzyAhihZb95yV1dUEOZ0zopTk1XieVJxqpo1VdFPLL
TqXaTw/eZf/8cxB2BWtzhQYhpMtbO16yKulxSipHNrFU0XyfNaadTgwBuv0YmR+mBWJgB1WQTJsl
9GpOeMg9RuE4LY/fSmqu9ZS5dEG9U9oremIsVnnZmoWwfBV7WpPV5GKgzqcw/Njzz1ZMKD3idg+s
I+rsoyj1N/VLkXpJXQZPIQhXcV3Jqpo9Z+9LfxY/7XHXjEQsOl0xFORwkUXDJunhwU5sr9mFjNIp
seVsW8OjlDBtJd9xvx0dg0FLFoqDJvPToKmGGP2qbDEQkHTl4qdbnSfBS2xuVsoKJ+ye3rppmabT
4ktNlh0818YCQkeBVbnpbCiapNlLA1yM5Kyri00fvzR1MoKcMkKtx3ci4gZhOnf94GclCj0hFIFm
uDn8Qop/lX2AzRxG/55bVVqEtYdv46Orju2Ad4x3HRPVZHt2yP/iHRJseAtzsYvQQjhkXYXeKVaq
ZjHzdwFZw7zG53EVNbCH1IAUE/OKOeIIeTjQhG5cfrdUUvZS6mEKLdCfh+UNA99c4LrKaiLuRe9X
0a4Db/oYtrqlm+nsz3qIEoDvnQhsy7OcZ6qn0GdkxKDkf7aTTZen8ZyN6/3iFeLBcnPARSoHqLND
8sr+6FzXGr1xLZ3accsTd2vvqAsxqkpwR0QHJz4IhHFTbBAoA34S2DJI+mtBLepqfMnNn1gfgO9+
1QCdtQGk/dT7RZHrlUsl4F5agTstSIU8WneXlRSuVVt2TFplnE8iHjTsyC5mPwUisn6qAch21Apm
mBYo+z3wvtxwPMIa028maXrbg8jBnNDC+o5opQxQfOhh3aiCEhLi9hkpl2J/BmvvOSCk/Ucnppb1
tRXzN97VRGIWT6yUmPDySmVqz5Qtsoz4pPpgHlqB79oalF3MyeJHbtJbG4iiv4dHlYVwnQIVkdvi
fc+gAXM7LuGKhyopz3W2uMdyAZHKpNR7h0WjJAJKg2DmiWUb/7dj4TPBOFCh7tzB8/FwAshnbGUJ
m1aaUyOJwjNhO9ncWJkrB/hffCaRGpFfEuYVKh308eZ51Z9YSABRDtPuFr6GxARiudyXnPeEVHOE
DPy6/8DLL7Gfs4inA24cUhdg1bsdLoObGThdu2iHTA2QDFM1MAuQCzsMLyp5eQJZ/vO6uDq0OfJ2
yHl2RBBhmiOFg1IPxg8mNYbilkYHxr7dKgWWsRH/DOf6R72uhHMp+Cm07g5C0KiZPLYIFIz9XYGy
YBYC45/aFS8t1FtenvqfgMyJJl1RolybWCYYMZB+OY7mrM+teR5zK12xcbMibIyELHPz0Vf0uQ7g
yKX+ffvdEq5iYde+NjUG5Wse4RWUJ6gskLkEnyWe0TetDzX45/JyCbSf0HNrP/QIlIV0APGZWnqZ
mK1p/E9h9Dh4NNawMsPxF9DVXy+MNxLB+oDxa5179vmztglAW3waEjkvZmIn2tFY+djDrmagalDk
p5OojY2THfbK1mZJFU8TONOVMsckzlLwmvstCdCq0RsU6LcSw/LslrSKI6PltM/3Vii5Px7WdPcJ
qMQUYUEq99qMfUh5hH7IDYiFbjjup0UPkYWFAc2+VXWH9IOkPMIGXrMr9Dizbc6fOs8ZefxCELGX
gI5uKgnpS9q8HE5atgEqlOmB49FoQO6z47N9xGzegrCD4UZGsqZcvnUmLIgLWj2dVJHxYSSA1CTF
I7f7ispvvzz/xi6vG5MbpD3GvbsDrq0o7HwmolLFMFNJOp9a5jOCKPPn2u+n9wqguvyfxLt9+PlH
vl8glt8TaCN0+3Wu0gzcKGVbGVKw9a5Vf9ClMcGrm2fyb8UC0xehPXmi7B59A4xRz10PkjLQfidd
UfRcyJhPYiL6Cr6qegRh3Yf4tsi1+NhZDUZ8Gh2Dof9ELVDLTKqi6W+cCLXgWzecKjLRuv/d2VoA
ScQoVnNMZ6gVGxe/z9W+XWNPCWg4sL4zk0X4BANtQGaz0uVqW0hgAfe+AlU0la2GoxPaVqS161sk
7a1z8EDq325Xi295qNacZ4P4ZWQocQGoY9gMTso8IAG+MxsEs/mI0jsCLE8DrZoK8j8U66Q+860A
1UnSPagQv/3ijmMsyX7rdZDCIe7ZlVVbKj0s/Gi53oAZOKEhbBUqN/UpQWpdLeMCixu1bofHqmEJ
oSt3trF4ciszhDdQgpJVVvseq7TxSYk9yApjIFzmF641MSmvYfxusOFiI6XTRz1nF3liZESBn97c
TtDD4Hp4uZJUpfQPqNRJWTByo7ZT/FRNhteuCegONGHz1naDVkJWmy0/ZYpHgRBxwn4lZb2/Xky4
MCGR1tQHs64zZc6VfYqT2qmgi6MAQuG+zwgGGy+doKZRivF2XLaW7Jnec9EyANQ86lMX5+qXm0+0
0dM6YLYP03pLVGufXJyOMa7TDGIfAZ1IF5dC+dDpBDq15dGVWKo6h7h8mwM/AKvDw75IVTVmp/bf
sRX60JMSA0NWvekjQ5m8d+jYIsfmAuf9OdmpA7dha2jVy+XSNR5IhlNadS0n9LNrSUTxY0xEh6rE
clB7r32EVzinW+Xjwodpa/UOwpb927++f8ssvKtnfzNPIkuiWvNBaL5Tfi8YNEV39mKs4H9O+S7n
c+g9GVyZvPljn+5SvNjBdcJoPrdi0B3ZPvsxJdjMMLwCSSMvaK6sw974eeHg6iACTT32RPvP010Y
nN21Q3t0ua6DcVeaQRL1A09sl4N+IM49P1miJ6ZJG6mK4sA5vUvxtYeVkNIb8XG78I1W0OGR7WOO
NvhKmbM3FYTdcVtptUqIyd94z36xEA3WZsMRoeQqhys3UrGtEZCoMB2x657L3vVok+c0vcBfY+V2
pkxC2UjNLpmmMRTMxSDWLlXUATNooQYAwBCIw79VjuZRcQ+xKNXjtkw2KVtW2IpkLOLrZtAz9DW5
Ab43XcBN4RhwBjPGmjQjxGk5WzLYlQDiRfafrRc/ZKuJ+Jh/vNFV/ZyOLqGG1aAJWmTiAv/9WeR7
AZWMrxDRIO6bYn9t8bcRpfBdh8RP/04jOc4aw1KbQO37PjVF66EX2+hRGLqdFI8JwtgokNDTXnGF
9RMnGvn6w47jnY+E3X1ncymwHZHg7x8i5zpiCqdgOurIMKppMzb/kKtgbhO+sJYErpZjl02KNDIM
JQ4FDQ9BeaK2zfX1vJW6c9pbbdJtOIJJ6D6RxntjRbSr/DLD/NqAM+y6KrqJhzPRnM/n7+BybTqL
Jmoakurwg427/8+Y/b7tIQyj0MH59BC5gzIJbTPAOhGVkBin4aN3gBZ1DeNYk0Cz23ZgCoXVzsdF
woROKQtvHwvWTW2AolNVELsWB/KBo6gm9+X3fE0cFRJdEwxT6ZJAv2dzYyqqNMHx6bL2o1Os3die
ALExfBl3yNfdvz2t09fLz+Cd24L5SUecTOwVn1IJT1bddol9zcCacItM93ZLyIrVCIW2buMyMVG6
QSOO7nePds6IH6WFGhK5w7L+TgGsaJc9T6abrIvvJO15IHGmIL+v5klyPxc+nVaOnAAvZT7nPC+L
Drq62iQwIZoHck7AvLVOIZP89zekzLuP1YUqIz/Ng1hEa4phBiL69ek/dwKYKokCZR7xwKGLu6L5
tNn1WPJR36WcEeFDH7Lp3X2BuQ+Lve+Ib5vytcxj2P9B8ec2GSJmqFoFgZ4uF1sYUq2EJKepw9/q
cCZoOUttIlDrxAHwUE6fntWvA5vCycikMbz66Ceh+udBvIS1koVTMIHDP9LxLcszbS1P5TixqQ6e
pyUMC6utwCHnlp84ydJTI+4O2YJ3xpEE1rYdyVPfjHAvqFpCv34PhZkyG7p/QtCqtNe1xu/PbSJK
dyK52kGZVPL3glU0ycnzESI+tsIVP9zDC/wKGxrNJAG7k2ZE8I4oWdhpIJDpV1+6AU3LfpWNCypi
S5aYR+eNseSRIhT1S7sIeyoKfWsoYjoQj/wHZBGExPsBuYKR5kiRA711xb70JRtOmoPG+3GrmV4t
vKMV1DAnCgaR8sn1Jfsip4Wq0jQlHwCGITLUo2zswztPMlM9Mld4td9rsYUqr3VmNyg7bXuj5xnB
I/3fKfR+Q0bigG8SSLjiLYn8/aar0JtlTIlSCOddEhVGcvQ6hSIyJic6lh8msiskN5HDChgzqpIF
XMEL6CMBIcDHyXNWHnjuvQYczAWYPWBX9AL35uJ8u3jRGxwbGiYf+3mE5muU0drWK0YEWY/sghCr
9MUqRJZzF0o5q81Md0QCt7O9reT/hJx0fnHn9ddLfyNFCi567BrfwhEJQnOayRJsH/mdDxh143+m
Sa3RTpjxPlM0e6xhEpmz1xAcqkvb/phHwAlmLp6seotgm6tcnLsNE9L5UV915Q/OMu37Z2KOlHGY
8bJAFQNDace8Ix+K8RW5koabO9qktbbHnwT/BNTcPNOvRT1Fn2lFqUWxGCSnF7K440/BE/tADRnx
kio/0JJouaVAGy/GF0MzUKorJTOn9rp5CRgotaJXNtURfOth/lOn/D7qFHPqTalrNitvL6kGDXI3
pp/lYrghaza/uFfHmv+pXLtpDToxy2c3Dl473UULU0g0myBk2XAa+CSN99eqm+H/kI7KHmY1h13p
u5mWaZABNQdZFmBMN64tvyVKJqJIKhYgnc4N29YCJZ2f6T/b/6F5kEqf/TZyuc69BItlO2cT2lt2
RRQ9+4wVqp9Gdt7peIIv1gnuqwkkpEQR6pXOPGzASog1wJk3TxIONvy9tqAd2T9poTe9CQ8Sq0so
N8mhz7aAaLePo1OvYKcrqzBMHpTMIKIf1Pfy5TLcm6kGRcpVCFewv6/ern+NFQncB+yvgMEEqnJd
cdEGPnN2fyKVQdnd3cjTTN81Q4uPzIHX3myI/MaDAe54Sc2NLgBioejPCUOawpUL6I/MuQ+s6Gs+
CskTRzhb4C5dr3sXhpLL26o+Hr9lfX3aPIq1d4klay9x1EyucDb29cdZkZ6ylocrxTPkZN+g68lU
fC1+ZWOwexcswz2Dv/2IuuHlpdeVkr/kZ4n45NcxlE6DBsHVlWOkyNmPbWM6b7bOQkyL1s8vzIDx
KzqmCqga+L9WhI7RDjJgG7hxGH4MhYwOccEEmgepofw6gWO6d+JeRmKCn39Lo8tgiP4gY0bAk6Vp
GcpkjdFErchA9seMkKCvJgcFzaiSM1hemHIpG8rKTG9YwgCfV1kCFVMFncr/eu+oABNtvp8zUDwq
O/xFYHZHnntram5qaK5LenxKJciAME0BvWAdP98RSF6XuZjxf9+b08StYcX6dO60hS2IFtIfYYrh
nNAgvCNJd/bMqUgZfy6o3RfDcWO9lkTzIEAdM0typubhh1U5V5gCNk6msJFZaOp/Ckf7QSBu/pTl
dOTiEWAKdz1sjeR/XQFDZF0JZaAtivKRKGZo3C2xS8Sc3wawWHbmLXcYbtf5JdN8SLAP6kLhZ7Fx
pSP7RNXcdYvly8mypRcOq99X+JkiGzHAueKxF1K6Vm2br8I88j7rNn1eHsnUSkP0triAlISCeALM
fDpVrKaBB1MaeDzYJRiQLnVb6cAanrDV1W3EDTJKNZKB7UpKz+URA7rvHAZoDHJdxeuZPqmCTLTN
lfDr79FNpOWyeeLtouWsl54fAixELhcAfa699xTdnHw1/dExCj/qhm6cQzN8yshQ2GlVNnChyg2Y
ztW5EoPf3fDmBtbHce/RoY3+d4UEYAU7ZmFewIbX/JTq5lyErflPOuYcV8E109Vc9GUzxaD0V7WP
JZeUHo2hrfJ5NFsQQ52Lyn7qkx224/RZJn+92RIpz8ignJfPD8zo4cWZDk6p9B69U4jKg1BNqgUY
iG/5uOqRnVKB92Unp/k0RtkPw85U53AVLJyrUV+Mk2VR2wYd3aVeYs8TDPxJ8PC7VPjt9em/DgPG
FSCQlIWkApFtUTM8UYTZoAKqmQjKBU8EO5bbnv12qikR+MFhlbkHqH/Ulfy3DWupt8ShGSCT+uV+
9UnmgCkRAEOJjQp79xNUrPT9n9/gtbvo7/pEEtGCrSvS31kNx3gUQzx2VfNkWavb4jva64tXIco2
2yYV2jbKJ0LQEfmSRlqXilrf0udLCkxiWa36lygDAfnuB+AqQgNleESQ8NghH7iwx3RPYr7XVTRR
G2E7rocKnoyIt+5urApHfEJ5ptMopgq5XU8d+Mp9RfvlJ9FTYIhDqklw0yXMSjiaHhttqqKKq1zT
UU9b73TY2uIPcFiTFkLmMcbmQzG0Bx4tzdzggcQFrcl0c/a2nQJ5bI9n6cPiikxVmUn6bfD5eU3O
ob8u+z6YI45UIoZU8L/Y4d5CZJqna4ruc4NuRxeZnUtI/qPIEFnLQQvYIHxKdm/yAgs3WRFCtHfy
pojVBw2qRb8UWa0YOtOTlek01TwuVQWFCuGjSrfqfIhewnNt4m9WQBmEv4Dj/YAtlUd/wMW4vmFJ
M2h26522lveJEE6FNU8990oENrsBJoboDZsg1gDZz/g56A9p9FGTG85UPB8/o9Q3vVwbIu8ge/fC
ph2LD/0CRd8DJPUnPi810PYUoCdunMS7LsHDfNm5y13HIzmpq3QhrQOac6UiPMB2djLdlk9uMF2D
R2bRvzI/3f4r29ohO0YZyFCsYV7zeQb6zRqwkN4LcSznTT5XYbi1BiInjZc5yN5HM/cdQaVyPUtv
6FSpqOlUPMOnXlmyXD7em1/07Lc+i6aq7mlD9wcXOvIVi/pSGyk7uf9OxY/MT1ULvIYx753K5ykB
R+kgxxfnrT10ix0PsUGIMLc6tnyeADovPTkSbgTmUR/hPeqok+A4a4QZe5luGj7ID3e3ftcaWBlx
yzGht2GVDz94D1TxHWa4+KwGy7UFIIvso45lfenbk2bU/qmY1bUvGJ69286p5F3OOHVO5t7Kae/l
m0Q9NRcY+IaljoHv9KQn+HHKlkmVx9ftVgRwpjisqqKf0yxjEoGz4TGQWM7AqVp8zgRAblVqJLyT
J/0uZUkF8uxCJDzq0uhFhfCNR6up5mbad/rbrP3n9cn09H+xcTnX+Wi1TBLUrPsCmTn8bjJKYJ/t
P4embTqQvIyWRmX14Ohghjus5CDoIx0ZrmCAD2bdlpLqt2/6IFbeTvmXvjT7Ciwhs+z+HQVPNi5y
74h5zYS6Sc1rfuiPzx8UVizHKfhh23eizQKyNhUa9LUNRzp6zj+F+Tb+xJLm4BYr42gurSPRt4x7
As1dXF3UsBlYKsQm+0S3bbbcVaVf/dNzy53X7/sxoQGF0ZC65ffhCDpTduvQemBnHafBCeAd1+pR
aywZ7UHC0UDqmb3yfeEWAalpCEu0yaCMI84Vh4yLWqkOnLv9w6l3YFwOBtJM5gqpS+6WVw3SJSLu
9Hq4+/ilRr+ImOIxG6ZZGV/8mq7iIk0SVY40ZZaXV1RJM3IND4f7F8MTn7s3LhZRVmASq3uiXYxy
gmAoZy9SfBPboiFijvs684l3PedrO8zB4fzVkIrtUNOQHQrHqM+cIxxIDzd0Dq4xhOlqa5sNlqiY
oX7lAq6cDdg7Y/HczhrS/VUpC8Z0zQZJnqn7uzIC7nk4cMja4WVSVZlmSrkI/iKegiDB3XnEuneS
P+QPhIV3FznFUKVMn3RlOS6xVbSafWKKtZIKdydXk68vME5vg/QTgmy1tW+LesQs7Hu27nnF61Zg
g1JkCqeR249HsrCKDXC9PI4bC88sMKrDsBQUdM5ixMJgukFjkRl0gCczt3VV1JNLsIbK3MCtJSbb
1DiJAsMfzLIPEgmRaNBBlf66Wj30Zvqr16JlykQXs5rM4FWNuHJodprT4+BqnRV7cvHOqxI3/cbV
EHW7eUwAXQHXBZduuuu3Va6aheXZ0AU29zEeqTk5eXjkq05AsIryDxNZdSZqwsts0EN9F0MYs9PB
s6yptWf4S+B98epgMw8B4hjd+zZ9+giwgelyXkb/QGf9apCZKk9saWdKqhJh/6EOlZJviCKBbSqk
sH0wpD3Uye/xnc4ASKzCKfaq/ECsZADdJZbE0OOeq9q1ApJd4Sevt6/ZQzYo9Hnj4kifR/rW8pf1
HhTNZxdDDaQyCWw3aZP5KYuKt5O163XsB+Zm6VlUQiCI/zFFuOnz3IidsJTrTL6a5gaLmZ4WYymx
Ig4XzY9YsAOZnm0PfVJPaE++3IlYF7ize+0CvIj1LlFyeYOcSTWXQowpKWRlFWvvhz8qtdTmy0T6
6rtblz1U9O6V7Dg8cjrvsLoW81knnaxYHipBtW0nzHRzzu64KgZ75r+H/uZh/ZS4YWB83qqT2s5j
WUY/llDaANr6jgK9Ao9p3veAwrP95xwn5rGC0wOxyfFC/0ERE6m38tYGuc5EXSdmZB2MejzvHY7H
i91Lvssj+XRKvtpoKU0Bbj2rY1Qjj0d6K4yGYXfmjg4GDbC8+MEzdCvil8gJfxRTSnUAQv4HoRSB
kkGDFpX5qK1NCAOYtRbRp5I8euZvWEEyyH6O+krSx6rAoGUqSkOXXpI658CAlwVOi4haDBQ3kHYX
XWP/EHcprKQWoRINbDFEpKTlhZpc9/mPBVmMgD2OYEizVYzbd+KmQdoP5OI8PgKZTuv4Dhfw5+Af
7qHHumo5VsdZIQ7qgEbaOlUbbhocWmUGuehpqoohQQX/qaOTi6SdiIqsZWgk9KTlWFrxXRnHt8Qr
cxPVNPGOQU+exSpBJ06WyRRH4fpkfCJEws7Il19J/yzb3b8LNFyMXjmt0LQi/Zt9knb0BD9onrXC
qZVTo6LoSPcyXAoiJgQwumnXfBM3iG9HupLopwWkQ0fO828UnxWv29dHlPgFEzrW2CBXARzTSo0t
3FdJxUphGp7kfJUkBvI3OI0GCJVYKWnYQ+BaQLKH1bsTvtHIyY1xh0GdPWgea+IaG2fdSuboTVBl
bsH2wLxP94si6vRuq+ZfAsqmry1oim5aawLj5pg+c6WG6ETeQlUw9FWqKlP6Oes7FeF0f+nxUwg1
sGEU7P/BKZZj/s3dssZTv5l/qL+hwiRg3tAwNoXqkQhFt6G0vLbHVhATzILZnmpQS2XFgclBnqg3
/NqjAi7XrlnsfyiuvjhhzVS0lggalsTwBTzFsKZUarrvKDj5hAjj1KFGqS9jppgMnV5MRYhRV2jv
wX9v0q0+8jGjCwUWJpUeswzNHgRKFP9v/54EQjNz4fxCzGBzJ6fHyj1zkayqYa4xhKiDIF7sxP92
Vk5j0H8UO8GRuFZCBup+v444C0iLw5mmgQYm/x6/eV8BOy1Uu9M1CUuwtgSTL5Z0YtZOahsuFVwm
ht2sxZKyVFqpzXfYxTDLYrCfmsT5UXdyNh4ve/o105BxZRhUZwIos/rqH6e+EzXe3/l/y9kYiqvv
DTrxLsiOfXR3yy5hVcnDe5G/ohBOH6rYPmpqx7I4GzPHZplLZRUJieU5dNlbPsfn4MU+AY9zcA2m
+sLyu+cLsbGGKz17y8xtWSXw7AmJxdHDPli99LMI9R0LPUl/dOy+U438j295si+68mIoWfuL8FFR
/zsZzU9nXrdr6PrpnCrLykDo8YsqP6+jWa+c3HbxKoUc9D4UXTi8LvAncIA8fWpb4NzKtcCNKzrs
pzoI00ePmr7Ygp9AByTab1H+OEMQOXygUbCLh6nlYf9StdxB/9jmq1tMzJSegXqsaX2hPHbGuOWm
9Xv5o5CqCqQBq/hLzXDUQzCt88PYCedGt3HXKme1g48Cpg/Zv5UtTbh6dsiQD4e6t3HkNSoPffzb
EDH4v3KpGAs5tbypKEsmAHUejO2/tg8PVWF8JblpmluBczvgSfvoprg3VTipvBNpBQ8ERzkuBxMp
YlVBMpTnbsNJlczxlYyxwY+BiDpy24YAA+b4PThVUGpPVKLKCnv+ik3To5i1yBrja2SM35iDVSKG
1EkGl1CdfA1Uahj64PmsRcME/Ziq5esxM0FrGmTU2uQRg9Qht9Xj/ZH3G58DlhabHGe2C4jlmKWQ
7Xa9DGa831riCmeUVBp9BUNTDa9er/Xte28MxfK6oP5eaJ13w/zulfr0+HffsWwd4YddWHL7WGJ0
82lIdhwI+xQ9mTCRV4/IP3SLYcqXQeljhjfAMwRcqpw2rx5yFKSRMvMcG94y+V8V8StfwVsaV2fw
Oj39nP1kOFkQ5TMfLOY3p/XVR2rljpEm9umximgpWWeKzGE4QltOtWSNIiOxtPenyIVrPN+dn/EG
2wsm+KLgkUhDVH8oYF/sTLI+rUvZoXyLhDSD7qedJbtmgiLnJiUv/tDmHt8uPz9YjxS3qWLo+X8N
SvKAtDtPBUVC5f/ne9E/KCLTQwGPb2Bib8LILJXDvyXj9+1THtHwRmZDtwIedeahRFoz/jvCsJ4t
3A2EE8EjDspN34VrydMxRcvnpmna8KzqrTMBvALDd7STUTt0MfIP+sgWviVqLMkpyoWQTT1TTtcb
olr+X+XdgR8BxthJoRV4VL8MMMmShy+2xA3rH8UJNDbR2y3/q6o+/eVTLFx3VfMrf7OzEHmkY1LR
n81vi4pLrJ7nHkWaYRaj/S10T7cVSbj5IxbZgIWi/DgEtfsIwYNcUyupcruxADtpCG5Yqe4lhIIc
L3deRbsm9s9G//NIVsBmcXaa9ho3+VjOpm2Z4G3jibJ3n+2OfZLXg+Tleujrf1ORXP9J4ZcgX8BD
WkMOP+er/rJjt1tutF7UXHeyPQ6zKwKuGhy05w4nAM6leTeRTqVPZEHyvErGW9JUBl4XxhPlIVwC
sY6PMKi+zT4lFDcYNITBPf/SY0zYoUir/acDJtV9WoCW8gZVT9m25nUH4P/E2AExic8TTTNgeCs+
Oc1CM5GaDPyIsBhsTgzrmSsykBLPHs9R63Q3A2YSj+KysV1sGNcMngt7UKCeKLpWPcADx1x17mQD
nc7luYKFW6c+sWVO+4EZfLEOPFRaG/0buASdhxT42yQz+Xy/Ph01pCleD3gd5SMhZtP93Ehx+SYK
IdPUpmi0rsdFWf31M4LuE/aPXeWcNHCUCFaTditxw4Gu4mIGUZDxaJD+NO/oLdcMR1lXIdPSPwrW
i6xtdlv0XnRIBL3VKiOGjEArilmANQ7bI7XC8QCNxhaaVybSW8H4Id0UhY69gxGyyNfj286mruuG
PTdp1lz1oQ++0pJ3/oqSYsXpFNyji5EVj5otyzmzL+nWI9x0meEHxrWBIOitbJjQyEy2lfSsK9ES
bcDpAA26GpCCcU9RHhvJ8OVmEpYus9ng7GhGXOLKcjsfgK8kxRDVWTzXRzWC79dOPvorf6VeE2D7
5AyKPg3WV3AlaXOS6t5UxjEg1HpOS+SQqhhtrO37pTWuTbTjEMd0+bcueXimJgv2UNujPnex3Jj3
q8GQyjzhNCchcvp0Eqd73EtczCB1y5CSxvm+gjS2NrSmJBvK+B4ah/82pOny2TG11aOoc865ggjg
rqdTd3GCtYbYkbhBHxlnjMKocG9NELWSd2dCeUE174MARn9jXHZzaVsOBLlO8OckoUWtGKwmOp/J
GKO7uILWHH0A9qXLhKoY8wSsFmgi1QJ7lL745rLTAwLjyueZhXgRLSeSVeWqdCBwDpPQo8VV9EnT
zb4jGOHPsNsE8+Tus/BKYkhSoQpPI+ulPVVMMrqr7VZOZ3EFlpWdHdo/9IVKANK1qvr3TS5sbtLK
4bsUAIg6wEsfWAUJAtdA39drxH/T7rLPxkLcyxtMYfe57dmlW4l7KVMplnuudOySiEfmr2gj50RF
qinUe9xVQwcNN99zLTSrhx9pAYlPfQhjOl7bjGoQPqo07UsfkPspVP5L1zID0ARLk0KoZ0XfTiUt
NA4eZmDOXaDyYo3fERTFCCKEYCKmVf4P1eatVFfZEM14QWa9AngV5UlY4A8tEywAO0QxuqnHQUe4
ghK9mrFVNjzxIqA/ZGOB38HCSX0GHtDDihqXma/daggol1yNeZw7IVZHdXbHlii+3JfJMPOoa7Np
k+/COuCVxX9xts7LG5ZumWPP9gpARSRbnTZNdwZBwltyZ1r73Aq03k2gfdlo4QPTVkYKsVjzvhYm
J+x6GG50U/jHhx3ID7jOf6jV8IWJL5ATQ1bl135YLsDEPtYw82nz08x/Qn9HQsh9J8YGl7Tv7/h2
xZuFy8/oAK7LEs5eVF8bBb0CTAnzgnfEzmyohYWK7Xxj65idDEClgjHnG9CFk9WlDVuvsmUAoBzb
5j9xuXmQh1JrcpCKOeD8+Icrjr8xg4kL7acrfFgRtdil3V26w75rqFymQbkxYMQ9VdRzMr+A5Y7u
LFyzEVfU5Jz6Tuv+xWm/S86nrCBaDLC8Et+gSS4tQKBBg5fjElTQPPfPjkB89r/lg49SDNKEVnf/
ghCuUuArevp2Z5gkfXfVA1n/YEhkGS/bnaOMD6U475NI48N8+9ySQ+0pbYPD43cSfMk9ADgkIcGg
A17jZOVonPnFKaQpkrHxdQLeaqfIU9nq0dPmRPRCscxS4BO2aSCc4uHEnoKQgAm7YEXh5U+G6kAB
Y0JMjg8EVFWWNvXn+qtb5OqfKnkOXpyNOsKaQRqi+nWJEj7FLx/gb3nh+z7inzSMLq44QZd6djEi
Z5Ei8Pd3gCKrWmWL5QOwc3DNGSpR+wmNP35Ku1UcxLLCZ+AiU2PPh8fP1VOB4EmBUSjTfD6fvkkd
bY5pIMniOjI7nWhlUBlLZWfoqcn1y1A7VM+1AuZ25ypMnWdS9EMFlIgBkpViQmdLU77kicxyj0L+
Yhyo8Ikj2iuTrGSqVN6WdQii73tzCGleKiqmXQAMpdkKDyg5tv6Tfb8SFgeOQFgNM+9oI5RtTPO0
ZFnTXZnuOEaD5gE3spm+AaT97qfTCsP2gSK7Md/+9j/FfWRSKud9zb/prKUAaW9b9EnhX2fAo+9+
WTSzuuLTAUdQafGfqSkdOwDfzu17v6yzg1WdkdvKFSIUN8OxAS5GsVfjjj2CjZ/NCZCNk4ybCafs
md7npF4d+eMOjCgI6LbhDRR07ccYMCdKUHJipOa+UtCZ+FsJ6ekAwedejnynoq/YKKxDtmr2oT7A
Rkhe7Fkrei0RnaFGMJ6FYn97ymzFh8XTrEpI+9McbvZgKAeavmNC4vWqv0K5OiFj0JhLBKCxJ/kQ
KlMQmG0Xk5NjsswClRLq6Ia3RLawVsHbM97NfZMNn65T7n3hl1HEE1U5enIwWuWAtw6NBtl+SAps
TDVUgRuLkJaXVMirD80ru+XjoUviPtJ3hDrEgnkLJHjlSV31M/80YWG9WtoQI6EbH4iGmgNuqXL0
zehpbj3YlLSC9j3upZ1axPpfQZ6P8DLOBUMxqTDruLCd99KZfOJTqh/MoXeaG03DXGgVsyE/B+U1
T74HMu7f6dIiTDEJrMSLXQbLvt6uJKYkB3Tovb6rpGOJXw1YcxuIngopWaJyJv/RMlo7UsT4OeF5
NRjX0bzrYdtbn4I5XxWQ6bBwuFxCzIW8mBg4CyVE+XXId5+gR2p6d3ygj2rkj3rTG92Z4+buzm3t
kRdT6+nX6qDGLaj+zRSSbsVXwUHFFtSt8ICC75AEOijUsxBuNf6lqXqLdRljFLX4dSIXEsPvQ2Vk
MS/HO2J/Du9ofTx67mlFiHfBlD3rjSoX3QAvTIhFd0WxLcM/rYTuM7K5kkHJuyVW0RretEOjVHV3
WIUNPXEcn97qbbQ4bSNyP3fAZ9Wfh2OFM2cIVVJeIdK9Lgyk1lRxS6q6yx9zep8/q6YaW3Ah1bU0
djJf1M4pf0h8jHnb0C5BdeDwhw0WFbn44ztxIgkPl2I1F6KpiVkljki7RsmrHA/ZZfZEO2CNT9ZC
Of9TKNIj0MvzmZQvzGMwdGpgBzIYz7/ND2Ie938/9s0hu+pvw6hz7wgO6seuNfKLexA67szKTdfU
3JjDIXqHcx4a6caoES2mpvlcD4mkoIomahHFKIoLz5OCP9+ODMixXDRBCNkZkGRh6DcbzO1JunXl
dFpZ8Evvv31FxXlX9gPYOf3Ea/n6M2SGbRNipu2p1NT3VPMjO4eGklsv6j74HwC9dQRhkR8B/t+f
TIPW4LB3ijVsB1ujax9VXd0bTiycn/zKNQhWKAHywb4yXb7JKgY2HjT0g3Oww/G7MWjTbfGYL1nK
LyFWgDv2c5hHKwXf/EtLgatob6a1iOH77HHpxaKBwbGaGZVBSxXKKp6ptOVAyjXJiHzmLmmSZZO9
3CedgjFbk3/dms89KB1Nh8PfAtEI99rUtZuzLz07AGhlFG7xesJhuwlEuawe/n7am7uPmcLF1LJd
vL21sqTB4sJGRWQsjdjtEq3g+1BQ+YOzGMEFy4uOHtD5TYANNRISWSutbo19QFzNcDvlxQm0aBBd
Bk2c5Hah/xQB8fSj0A4BiL2HPj16RUFM8NgCxsE5EvN9cdBrjV/LiCJQa+P3GK3Y2GwrdTxV6Yyh
atfUb4gteL90gXcflbx/fmqThn3wggc+Z1gFD5vlWa8RZXgoS6/w63IjPSySUeLMWrWEXhHJuFpr
MOb9rssIecEBUQ3NkZtWQ8w/nfM+74D9AQog/FBbLoiT5zbEdCOgrV2Fj+d5DHJYaGyP5HL3qc5G
w9oBhUA72qsGic5ityCrO3ZQszt/zzrc6bXM7G3fCy7rjpGqz9y7aXH0F5CSVEfEp/HrQqzjfLpL
qalxiTdoxZMpjS4Rbl9MguXwC6WL+FzahWV35x4lcyyRG+LgvJvzdUBU3DvkfZ+gUDIWgzuO1dMf
i7u5HfeZqQpT8fPW+ZykM+grLfwOKAsDhiAmik0z5LBwIOGhreM0H+IsY2l/OM3UnVcGWl8aIfJI
y3HOI8pyRJNG3+e72Hjzjw1peuio96s61teqh0tZ/mvIAn4xq5c2gEdcqI3+ehMidRkWWZ+MnyDS
JFv/tuOUWzD3v5/w1kHogbIdQHzOyPtqr1Kbr608hLgkudJ1oqNFzgkO/7xQnJ7EPahs4U8+WuEl
4EZCfdHFP232l1IitkHoMshS0ow34lgXbjW6Prz+qoiSgRyvTRs1X4m2V53qiPuExieDBEB+6djq
qV0DF0ZFhKEPyjnNDHZDfmdkK5/2Uu4FMF9K7vKRbgsi7DwiRDWeBCOkAbn0mJmtnN7qHkQuTrXL
ENd9TEfcMJB/5yNZ/r97HSsUyAZ+Bk7VBFRlKu6h/tHcdWluPcHwzkcicrefbK9VGNDL+ba/fkXA
KCy0kSefvPrkp6YrZQy0qJIMIW9/r1txye7gGwqlE4m3FqFHS7JEsK56zixzi/kgvaugIBup2JCa
KEq03Tf+TD4/oXVovqiSe2MR+FMbKs0jLgZkFSreDJkVi7HNv+Kfm4rGrwfmhiaNGra/RYPIireq
iqVKP7EXgYn63fNhFx2uwAxeijAbClkpY/AWOYQhggQmQtPJPOqTQGsPJwfXgj4zWwZ0XlhYuTZ0
3yzd0JdncHPFGYoyk4v736YwYS4Sok9SawS7DJrJeMMyYlnYn5GNVkrP3JA0NuKLFr1BzuxRE1RV
6f6Y0kSoyKiaOWcuMM+AB4MadCbQyIGHW2FJoJfsb5VYDBi5URZBKYyXtT/L4kUXmnzY6YQdPvHJ
BZTb88nBBblmb5WZ/0gJFbNs349R9XcH90r2BzmhPK55X+8W9VpV8QH6YpMtHGHa56qsF4XQx50V
xOadXpO39TeXYAfBLzy4TMRoXR+2MuZcehEnfccabGYYmKZXvn24QuNHMo/DQ6bzOwLIcrMERtjZ
lLH4T4+RU6MVgaVdvjktYm+oaCmJJQ0Ej+id5lVXlma1LL7O4+LYAH7H1VuWDe3SgnZPNStfIBy4
n+PAtdFTuzhAvBj6oZPiJwErbyYcmg59fTMQRu7oJkWAoL6fugmlAn0Vwo73pVqz7VTFF7s5kgS2
I6oHC5lnZ6JEbaxyBgyOTEIJRjuJu4NW3YEfn7kOFP1gi8qChN55AMqANE5xfp4V2nrLNHw+5vqX
P/ShKO0EA5oeuETRAcVBpvxzh+0qraDpW6LlBCdnGzOUSoE/zEKG9B0kwTz/vReSKwxPzbG7yXN0
aELbNDZ2x4Q95+BFSgHbWacbLMZGkqs4xuRrcnoa8Tsw1ae/yqqY6FRMmOagkYt58CXRKhz4Arru
9RRulHF1A9EflvnVJ/lWaPybZktWS2VFfzciUdhMcu6uwNlPigZ/IWA1f/JpKP7jrLwUXXBHOp/q
uQGLRNiFC3vmM2ptRMhNA7/F6KA/ec4yJlIC+Hytg0q0Vl5Sk9huQ1Akx3u6BTSYNp9Y9ZXInIQ2
NcFjSbSn7jAShf+WjpvoEp1uBna9o/u0h2QBaj5mOEvSCUBQYT37kjzqhsGlTDnKvVyYXEV6l/di
hQYZsZ/tBE/6+/3uaZR3UdOUCNvxE9axKSJXgY3O8dV3mrUNlYTPLR59KIJibbolz+eiHyv9xKP+
GIBw1nVm9jtCt23YQ+cQpdbNGW4loBayuoCFUsrFSWFXAfJECZUW3uvQ4E4/hyMAlV+fAsrcOzgN
auR6Lr4lpHR3sxW1rRuaCTp7Bhr7stc7nZXD7epyMPJ4ET+cGNyRr3/4cq58EqDhVC0S/2DmDg0Q
k83EdfnTSmtujCy35zawMlfTNS8ELbEfxojELPO0t60vuS0VVKlrxvefYlEDyEd3yYNn8O2BofB3
n70LLphvRlYAgNoEYbgK51F3jjQqPEEc6IgmNKhld+IsDcm+IxdkjmaRK5NeKpJ+5cUOpfm5nKNq
4D75WtewMfITJQEUEI4SND+llU+gcSyOxzpH/VUq+YOi59Ch2b/9g1H0B0CjRyx5PAtso13fV88O
7TtiXxGKPQyGRN0u3xOG03bDwunTgzdZiIaV46cWn3BlUGANiTQlHesc+FNIypluiieTg/hyJ1Yj
fPJsJ/s+jSSVn6Bd1g0zw6Qf/DPCiUjSihupU1f4nwDCTJ2tiIkWNBda/llNeH2nfjD+eqdi7ycu
O3IoU7DRy8YCWbbNpbKqoOXR5HxF+3asneHTEjuizsorb/oEMJfY12k+9KvxleUPGs8MT5/e31pT
02m23EGwG73TFhGskBjMPnD9qHe6JPWJ1DfPLtlhWwRrr14AK0ZKu37N9+MRRG2OSXQ2CxkRSZE/
/KKoxu9Rk1ZxgAK9sytZ0cXnQ7WjFyuYRWxPkAHL7w1ycfrdUPt+iGCr48QXZmWRAdcmclllbhkf
vvlYUFqVhg8jLdnsEsCulVFIV648OdONehIjjlIeUeLe84b/mvNwINZJdxnLnTuSLgoCiS90n+ly
XQfAMtAIG7M5OesUa/MoZKF+FouFCvX0U745ncWPyZNRpBFsaDRe8yzCjVtgPyJARShxL2IAlY4u
3yfD1r0aJ9cS1GRQxyMcq0SjOy8FiiF4p49hxJCIYo9Ed5IBwDxJLUUmNOCF0S/XqHDQzy3amr+F
Rh0wF/wA1lt0Nvm8cZXe3zMAuRKgzGdiRligu2/8/yT5CQHznXFuaocGU0A6QGURQ5+CzXYvIIfa
rZMsbQL+1+d6T95nZW6sukKAzgflOl7MbY3KBNgU5hRpXmdZ0Pe7O6P9KDxWCYqx7cX/LSzjXFoU
u6uvxeK3d/9GC0iUZBzkhe3PZOp2Re4EG4IJBYl21LJTBWYd7YHNbU9ckpq+Nd8m7vy2C0y3EBgl
fb2QOEABBDJkyXWthZ4/twKrstM1wTjJBCmIZeOHc5H3cY2H+3vblTyL1wYLCEnrvIApf6LM5Bba
8M8bWvnFlLuHZvPMaJCgcHHowR/yVVU0E9zHOfqw3ydVPROpFbR/rBryhvSDcgL4mUv/qWbU6urR
opSi5ZuGh0NjyZAGg4/9GEMgOVBQatVaeHHNiMFpYbZ9J7oUfb2XrnB7XgMYWShGCBTAZrop5LcJ
tkrnpZXwT/P937kmO48b0MEdIFnRlDdLUnEGz7x4DX24aUJzkfHkjSTGvvHibagmlDi+u5B/y67k
ZF1P4QpJGbTRHODnnh23dslm/bK05iFKDtRA06t626wezIXoRbrgTeO5xsh7hUrBRek1gfTDgD/z
lCjACLCLpq4XdbIW7LSoj1HPvEv1eM858nZMqUg0psZF8dCdvA9Chy3xQXQ4bd9L/JXQkKIzCe94
TwaZrEffn2Z/t04+3C6L0nHddySP6l2S/6PdFtzF86azwg6BB1RgvD8RGXmWKrRtiCZ+KAJIIrfH
nuIKYuox8pXb7YYHcSrQWs77v3Mf1fljmpdQAOU0bHXtXNNgNHuOGUsoqowr8dB9IaUigaNj/rNm
5DF5MZVFnUoAhnYe+cvzTR0L+K3rnm7DckjxbbTrGYvpZqpp08GdUntZKpyeYhWomtLmISTr5CRQ
aJlHU8LOoejfOCUEDzslnc5o4fTAsoWdAN1IXRym3tOChk2zLFN5KuPY8Zq25E3ZF7QNXoy+cbR1
VMYpwOdGpL+GQUL+A9ISZ9nkYswzdsQwSda6TpO8uoOQk+NxMfrcUD5SbE62RRtnNUf+KKsZXIAz
wC2xeMb41wkJooRZUogpIosyHD7IpgvqmSeUTaaOmHy7fooVEOje3zcH3jiZske7gPNxRzh9bCTV
PIJfbdzEDb4ySgVVJRrfG7V7bUuwNi23oBRrTWQxf6q04NPwl48s/IlzmxzVUcj88LQEoXcI/Z0K
1/sMioarjDvtgA7SlZOrfgaxYl7vHobjlRfj0HDb7r01aEd6ugqGnQSJb1/Pip3wTgCPyxgoyVQO
6lm/2T30AfFrgW/mySjmDC8zgj6vbJE5HdHBfmJIRc7zU4MmSKSUoN55fj10J6Vukat4T/bPMDk0
Dvsr8SAApu7haocUxyMAjSM4ATUPKHroVJs7+tAFOgI/9mRNV85ufvj3Vwnjd/Supe3Yrq4klkmf
PZBqcsaizpgcWkD/ZrVXvOc6cukOEUZMdmbLgfIVC0E/P/sVxinOMuWcvwJ0tSklas82RfdlCj4H
10CPmiSKsIXOGhYsNcavTL2mFmiTSiJ2HViaUri5uUGY/yyV+gYret3kL3Ln53lEd/4AZPJA21/A
ag+Gil5nVchWa18dxUDZFCa7benEIOrWRUsfDkfyX3XFtHqxSsSC5jH+USjAVVzaA0b08jV/TwBo
LI3Ce98ZJewYij7AgStNkLZXIRyBmNoWBoRFRWy6OfdJoRBiJcpHJzSNzz/xHlbfKOlq3uvbxVaO
oA++lHshiw/b4u58GVUsBcuGxAHD3uELkEAKEwJac/l+VolQPcUw/CDHZVcBuyUkImXh7vb9Suxw
s0IuOQy5j+5TOqK67XCEU2c3O51is21qfut2kT35dANCvmorPcydPMKBP4pGZMOXHoTMgsRIhuhy
Rf+ixpsnJiYhloa03gKiKZlr1cL+dnXQobLd0XFF9f3CeVJVXR4rnNhwj7E2X4YDI4w3Z1fvRazC
v7salW42Rj5bHs7+4Mo+zWhjOxwUy8S7Dk082HfyqxYW/TnzgjWdv0sWJdeC33nUceUm5DfK5p8n
An+KSJwM6JXiPOD6k4mw2dCQLfeWPQOE7Q+AvXpovwodQCLMvUjm1TTyxhcFOFYjrxKi2u0jEYb0
kzh2In+nOeaqMKdsFSTwA540R/0KfiPyHn3HPwQsBf/1sLn1WSrXVBXvPRcCbXqWOw0LhmtOUdjw
ShlPE68gFKDvbV66ip/8bN8RUWH7epnE2YvwwuRG28eERZ2gd/VcnXcsTJDdH3Az2PDvfEPkWaM2
Oe7pTCoyeGn5b+fhQjLu3s8UYhTo1q1RaYY900S+UwAbAN7cdJU/iivRQglV5/kTBfFKo9/Ax7TR
QnecQihkC4l6XnRf7EGWXI1BoSjtFz1XoNMLFs/i3g4Z1Jx5aeOppWru2wGScszTTYyqhZlnbtms
mSd5ZSHQ79YsFQjgTWIFDth55DU1uq1rVKU4F4rz8jdOam6HZvsBp9CSVJN93kw4wNz+FudJuk1X
mdS99VcU4oGDtoZE3H7T5KJ11x/+/VApvGa3fUKCpFoGnIUFgaLBlq2lTjKYXCghPutSEbrh8A1E
P6EB0AFkH3+ZwKPeQdkTt+1aOxEvmhJzPa/k9YOpmPDofH07khIgbOaIVEuo92ae4igNiwwavJlt
fhc/clOlV3Rfyh1nzvPKZldEwNMKFrNlpkiIulKDpyTWewSqdD6OEkfjBA8z6GAZLJZEI7NyoaPl
mOoSifGUY1s+bI4Dk4Eg88nrr0ZPiZTXEMTgu6S4KBFpJCDYbtOlX0gZqFeyRCWwnlUzR/ydmiwo
X5e9RB3SmMPq1P5Rakbwg8iSFBHGgvy7Q0Mo05GpWON6sAWylkjv+hjIzIWJ2AH5VYoJsdLN5xgI
5tND4z0mrkwsTY7qxPsGJpfQoDdN2pRuWlv7HD2Vneh3QQt0gNim8+xpps8br5zRlP8sbmvLGcyp
+OJGhJ+fM/o8WKojOGWfy2VYLJgJUopr9mKikvB6DlNHYq+YxqVrMd4KFemZwM4mD9yFXuBV5nTr
bAxUztwKYl/pewmJZBQpAg5rM2aIJZSArGucENeP7//pj/2frkapiy5NmclVhVEXG1nO2WJXEj50
sjNP/4hn1jBiZIsPAnYvTQD7OpXfCpoR0FWeZNFrd25vxm/35G+voCl38ry2B6diJI07Hr4q8Bry
SkLPPQS/mAe/4S6R8nqTvI+BlEdVdimfFzjSGWfMZswbxN2G2aWKKIChqOFAPjRJJzk5VP2i+N6e
WbUlieJKxnsosveTrS1ntoOGDuugjcIycLNNU9lGxeM+nhJ70QLVQLloobQ6njmyXF2AnVqt/Kpy
hYlEfj3RMLPkZlhJHwn/ft2oRHUqjPC6oHlBAidbN+Mnbhjo0l8evI9BOYNdg0KQyAbgxmZ+vLpZ
yd1eK68kp7zC3SbyZbC+lFDICU+gjvx5YB5ksTefjfrYVo3+GjQd1s29/RtkTsSWZwwLV7tc6UPi
Kyd4ywH30MQPnXg+DhvqQx9LocludRHQgh0geWgrQ+UPq4/GwR2IPoO+9YJBgrGfoXKfa/LfnIqw
OlbShChTUtLIDXwlEgAXZCJMMcKRpCwwywqGkoDQBrmqsw5J/O9oPDzTtykuBVoVUWJRb2YZHZce
2AW8vcIMaZIzXujLQ134RDlt7s1/Zvi23SGRZPJNcaT2I6GUBqgM6o63pS/fOPY4vim95HTuWd0G
sTD2XzRfJ5TpY/+SKSf6dWwdH6lPd05wF4bYead0pw8QXMXXaOQb4H1pvafomuJ1pRoFxvAaOwY2
1h8KHJZcQ/PKvbY4EZQTLsddQQwQTimrFexjY5SPlo4UIojNXGRFGjrHUBUudPh5X0/9B5dUVUn4
JCN6/4Kg+FpUpzpxEtlXAVaTNqQuPKviyaeVfOZO/NKBI8RYktNjvChQL4YpnPqEBk3N9jnWB7r2
CjS7klcsQONZantvnafdw3vH6xoBKOdIkKxGgIPBckiOnV9s3d95Z45hLnjNVVFEo1GifZpCvuGJ
jvy4rzQyKnGWTK23pJ3uEI3uegIl+6vdFDZFGVaw/Ei2KY7T521pwYUqKhp3sPEjeWMLr6Olquzh
C9UQ+nNEqUmZq5gcZNEyFIPGXz1hJIEB6Hx0LEQWP37f4yWhiEftwGSjQvp37JnRXwPrr3cMAyhr
BFO+3JQdHjW2UPJGUYZwZTSGmNruvmSO8GGjBuzEfnzVQN0lETXa6JDIfh9TATiqofwWAOBCuHf9
eCveBwq+5UyU9Z9RaFvQt05fzmdbB/P0/Uz7nBtjPZopiiwB0qZFTIY5gdoFpsXJGRc1sY0yP0fk
wv86pwBJWH1KEq5F04ghAxhiRFog7akVrZgZpp4PLxgjsL7eczZF6XG1qd/pvRL3PXny7fAJbHNc
1neIedwUeuto6KQX3f+yHPqjMjfOsRv9nOwmdFUP1tw4/d3pQTxCATjqaEOUfHq0EScJg83G597m
jHNzqH5iyScnP+DPmhcVwdvYYDg7nDB2Z/pi8oZ/WzLdJWbuoPeqS7G/adbYRfIvhq6mEgJeA9Hi
JmCh9exO8dASCncxZGK2Meh0H6xrdEreNBfTswO/soGvu2so/OGNumz7HaRcOMnOkHWo1rx3AxBQ
67dgmeuHDslqU0CKFcvzMF9mV+uRrq4vECxE0QiuBldOPV84PgJxrdc8siknlRYdDlFPZRLNGtF2
EOb51AQV6mxKlE/NAM7f+zhIJdc+/Tde28epNTXUUlPLHTvs91i+hA7uUoSfV3SWe45V+UC2Ruuu
I4EcOv5S4NV+uxBfqwxsw02LORA30mZFo3E3nhZQUGrshO6jYKWqSqqW6VSyWTYGxtl87NhBa5E7
vB8eJpI9HSgL3lhlXsW8tmJbpVsKUXo5MstlcvgqKdlcXjEF6HMMNn9kYfQbVhls/DBYBh7vK2rT
9kUzO01v3dx+5oeG3b+SweouWKJ56EnbjRZ3vo9cqVNkrjCtW4uizYwNcCRj6YZnVOyZdzyr0jyK
GeGsi53C7uZuNoYaCfdkqRNWBpGGJ2J3XzSz4o+ErRR5oZzMJ7HIzzt+fPUzfoelp16NrugVntmL
mQrWkm9rePciXnmyPBnLIej2VRECdtmkDW48LXZPuLfs2rlRl2Ub1SjFBwpGtMDQNtDZdwNydtHQ
eM99jzpTitK+djgpqFi9C7oosSllVc91NfB6hR8lqylJTu8TUKpeWZE8LZ2XiJg8CiXPL3NUJT8r
8Jikrri//JXvl4gIMQiz2dtgsmdD4wRQxa+XdWL14RO5JGI2VmpyUk9XlknjXXoVdzm1crX3bssN
EXMQKUk5XVS7cY2Myicr25UcciRe5UhQpWje4Xs0tz7DoiQwrkLkNxE7cwGWe+/aRJJTvwF+lJFT
dI8TlDFD0WyLMQUgfQv4m4wR6ahLb5w/zJDEaSlAa4lU8Xrf1y7K/pI+gAcHjhFF2EZzPeAkvqJ6
WJ8CqQu7/Gt7FPD94CSiOiIKtgBBhOGL3pqwXcB+I5bhnWAKw9KsN9ZpYINcF+QUgCLLMRG8yDFZ
l6OS64F1FvOTbc2QS6uZsJDXQSzziitauLRqnHtouy9dH//VQ3zzpSFM752IzLF8XmWFSINOP5nJ
Y4USQccrovZgo9vwydyptdabhM7G0oMuuZGgGX9VsDs64n1IPQFGg+ISy1JqALO69cOoHmtlnt4B
NbK3I5qWdmFr2/PUoLgm2Ff3C4+ZTlLvndvvRV+g6KS/QdOOwNAJQ7YeoJ7F72ncDP9UnppnUM1H
rzt1RJahU6exrxer/1IjRMhqclfMs8yrxHX4PfUKS0BSHwsGAs2X1hAUuoIpUmJH1Vi97/8LKXUM
P6yOPAjma3Ss6o11oZvPcGSR3dYjvLhyQowGH2MMMvGHq8PSw/7B0jMLMukvmSuOIftpfbnLW2e2
WWI7BW3r94g0xZnzCo7sI7dugVyE5n+XyFk5/1r8rH24VlhboGtqLBgGMVLS9y81NbsXNRWu9182
1/6WWEYIRJIswdLkpzwOjGC63rIKjAqG/aoN3NMf4giWx1XW0CkZtwMnovHHWXykVjsdk0vDUFg1
tYnJwJy0AzBMzdivb8GLSOhPN+JAWnVH0WSA7uzip9NlwDZ9tOX3VFNqCuuIW4B+WyDl0WuDHALl
7dxgAYD2+NiSrxCaUqXxvCa4AiSvX3qBttCwbbkdOlHhXOe9lXVeEwoqjGvWVWjrLxozrgUalKWH
kxjYzhkAWkG5T33TJtICeklSHQJqbBvvy/8zQfiMi/aMbIcI+PB1VQ271wEjZPUPqaxsrGEISmb1
ZNB90rRahaCcYaBlwSeP04b9kh+vc8t9fnyOcTfKcP9FdMxuSHwTiooeKB8lVIP2Kt4BZhREWidZ
fzkBBDj58Fi+giTSsuzZ1qiTPfK7fRaFGs65jK8x+uay6JcIcGTInRU+hoW+TLYzwUonlrPUTGUP
+rkufHqACD1N1ijvZSj/SH6a8c7OoCN4AuuKMalw0q1ZpX5PvcIQnZRN5JVNAIhOGcXCRrIpjxXW
Zpyo9iS/ZyMtDfaFFvSZkYM+pcTtyWrv+oUqBoTxBEso6I1m5mjk6pm894T2w5AnEQscSD9BT9aK
m1XE54O0Pd5RuIGT3P9hjpC6wFcfXTEQyo0/41o3AAsoJ/BTKnCdy3WMU0Fr9IBziz8RHJMVc9iD
dGuTakjNG7W74BXFDZtn8AmhVIAGTGcKc6hNoYG5iwQrCPBDs47+5IKZQsp9qm4kdJeEJkpIooTx
jFxEQZ4ikR1XarLOBtttVDIFHaeVf8i+vkccHy6LARyGL+B+mQUueGpNrimxEA0EvHUin0NzNFC6
FjI9X0m7xrTYXYid/mVrLc5+jHjTAbfd6R6kZ0hOqcrJSEvU8PalZPz9aD5JLIpWE34TxJOoTYg6
7sW8fbG07Xf/lbm/Ey4w5Opa7l99t3q5mYSWe6vuvaFk/7e5ZzXyTVgIvKUhPPhZ7f5hds+bN+/9
13ZnxXEQ1lEzBCMyBYZTfKf9+VM7jMKEymARBsg6tRo7LtjGJRh5OJnmq6vk7q8dhCHKKZ5a1JsX
lDN+lbERjo/4XY5k8g5qQo94A4/04lEtktKMDaghqF6cXmXsXiiLTxGEdyt6F++iEjjZrynHDsfi
6wKz2982QQWMjFS9UKwCDdO6dnY28yZTARVGvhaoTMndOYxPLLBb81kpKAWts5ilrVHC3r8g+gbO
BVLGtTWuDrh24y0jUSGFPOfY+TKSV0JpaJSKjKhBQDn98WXxuEG3L8R1cVr1ivTWzU9z+0DmhR/d
iN4W308xYkjyhqoW+yryFMbzzeseVWWPZrdsRMRW/0XNsK8vaQopjQWDUHqJv0oTtWhko/4zJmg1
A51BUQMoaxK3brD1wzEJL8QBVqRbg6UCe0LW8Hg4vjjfsFjjz0qTVoLqpNJaKAqrQwYqdejpBz45
Jx5yQZOvqA/WfMFzRtHru/CL4ZcO70PYUkkOLUo22q7lQpgrgB+MgLR0ubTIKDRyQpX3yve+4gdP
kJ++w7Sp9XbWR+HLe7syh27sXe4Fw4IcFCziAXzfLGCj8H3IsudmbY1pbXTcUA9wBW0U7vAFiOQp
U3nLD/u2pgcNM6psrSfCK9+bpRlwmlsmFLfxK9nXwH/Ne4krL+IaDmB1CaYvhQYiD/GLCp3eprq2
yOFY3eOA37Eo949UOio8YRrm90T6JVeQBt2t2x/MbQgRimbqhuL29qQqvMXqptKnlMv3PyVytG/p
8ZbKl9pKVrvIEsFRSZTdz5SYDwGgful04lAxgMgT00WND8UWVTIacZuanFQZt4sP0IPuc/3WJZ9b
jo/CTdL/pKWnW+DkKBt5Cv2eFXE0Rdcj4z1OGB+GDiraVg5kSpiYzUGg3arMyzVnAcTPxEnKtwmN
V6AsV9Gxbj5+LsUXTIwgCafD9+ypKOWXCVS+Ldjpot0sflFFN7SvkitUsPg2GSalAGA2CtlnB3OA
OEY5ZWJOmPffE2mKLfUpVAgq65Ex3AEwM9Cd8hBr816aPoUfabeBRSIH6KX5J0NUCjnq2HvMJ7cV
8xPeQryvYnPZa3maTMhvZR1yHONv8DSaGWU6UGzUnX8DaMyL/IJMw0WeWO5Fl88MqLdjQdT50HRu
5/cewy18YWkRBz06uw36N8n7qxZtl1krrGMWmH1KtB8vXe6GE/vE3Mq1fXiVxfHxPonxo2wm63lj
v/APTIc/BbJG8jiSQbPZ0o//tCC9XbbMU3a0tNfUd++KWVq1O/qefHVVkRI4DZVNE/MuBDdUNjYF
nSGQqI2T63HazVUZ+S6G1QOqI+YGjwrGB8ZGIM/gTPEyRJTgXtB81dlUIRpTMhxiotJJVXazWPby
3ADFDOLCirzvIuQiyzTNhEJaYId1r2wyyTwwP4/ASbtiRntwFciC4nVczBUMGh1AyAHk/itwvtM+
jp7LmLdb65XNjWcXcZW7uGKMv4JJYyjZu4h0eI5UXqJwiYX2fF/2OfarzEi4c99j+C2Dw3n2nFJs
ZGToewFoMOSHHfz8fQi1rbK5SJsU7tvVVp4iO+jCeAXukcTbAzIl1uzu2Hr/1NcvUqJmlZK+eqvL
HSMaYsM1iOlMlnY/c/Wy+voMdXNVk/wwsjTsC7yuaC9XqEKAN0WHfchbcTXICuTiq+q/mX6zqol3
m+xlZUtaqd6WmvxO3ASu7DJfqgAchInv/VoWdZocwppkLnb6hD287r9UXfy0SvY+8SSVK92Fzsg3
fkUQYZKsTB9z0chcoeHll54o8oizrxplKCp1twql4IQ5SZmkb8M6Bm7mSjDZHYu7OE2m0CFJcr8B
5ZXleb1nV3Ka0I2PIV8fHi6iWQkJAxlu8DzPMw03pPRL1zaeJThig69r/7QWawTeRzYCS5S85C+l
dkNxkjcZ4bMYIxSezsplcSOcMmdPgwgLNgeGNOjaxN+6C7SJL7fvYqYsBCPcnK45x5nm08xmXfKv
K+x8VMdtAHP7poTHvJ6GNrCGJ2clnenpx4l1phgW4xgIfO6NSEXL1YavFfSPulBQRDtCsb46L+xd
gQ84XH1XhV0DBe1jbp50+sHNBZXvLQmNtZLFp/ZoxPAiXvhpHiFmZePBqSbz1hESBXfsd4Gru5ls
HF53/jj6FMGVBGL6Vv5O9DxK3FHtv2Bwr7YKjAHsEwjltH0sG8QGvbt7Iy2TxDuISEG4dI2G406Z
bKuKeYKajoAuTivtD5H1/bGnDLcKILPlwOB9oUBXvM8CP+y5Cu13hMUsiiY5R/mlPXjokpb8q8XU
kc75EUWbRGYzefCBxMtJv8syMB0aPRYKgBGtJSc0IYXM3PR+UJKSTHbamd/Ua99Zz5VLFSrDVMAW
SMQqYrW8KWrXFSxO6PewNMxC1BqkFhY5KNOz8U5tm95q5Sk4MK7/DvUXmvhLd9Ov60FTCC1v1b4f
3sPSosLoTVHhy1mAJHBNTwGKvQI1AFfCJt6mRP7EB6cSjWnyP2mzJvlekoUUMll/uDsZj5wDxyWG
Nf19CXQ4EXyinELpKWL2fm2uOGAM/tSyiMH0ltcr8Jg+CpYVBjIrcEufNDAWSnnbyMzxw7JpaOII
RCQk40ndA1/dql6lLV0dQs5+n2LKWLtATrlAylqKohzmX9xEjDGGhIfsVGZPD2zms+/Gdemwxmhy
MhsaoDk+VDRZJJ0GvsuzyXiwfX/qQFzt2Ofte9fJnqxLXn0WliJHzjUpPUtB0/SRWbyxHF/fZqTO
hMT1LonCHu/zz3ioqk4/Y6Z8ltX6JibRvxsvr5Z6uZKvEysspTlSNtehDQ4OKSRigeKr0Yrugljn
a4FXaHd/WrVfqv1IDtwt+KnrsDpaIurVKesqKXh1tI21lsK0RTaXtFx0ZfH0l2qqPIHpBnR/FPXF
7SITYAgBDoHWxuru/pCHdqRrM5zho3lRt5msArqkbkvLFCsZtTuDFwIbeW/hKtwht7YNSvw6ziC7
sHZVBeJc1NVGTnSSEb+EscU0b97b2GOnBwmPtvsgkb/60YtGhCGqtpEjbRuFVRma9P1VEQpVGy6m
xJ4LfIpobmG4ufc+mX6v6VkOsllkJiQhTYlZI/unSeAzPjxhsrVKLgCeJCqlkjYQQzGBkoAlZtCY
NEzkoObW7Yp8UoVTyuYLE8YgFnoXe9i/9+G0FZxFl3yHqm1vAlqgFD5dXuihoAIknH/uWOVNka0p
5GzMKQIq/a60CY/i+rpVD2NwohGYoV0jqr8iYIm7XLKd2QFhVcVNHUiEsaaVFb8oPgdjagfk5z/M
Hk+8GPRiUuZejnD3smhvooR+37QMf50FHbDwgrcJC5mls2KoWK0trWuQBuZBRv0In/oWdNlDTvge
Td7/uwHOOLKZmP7S2nV8snLUm0F1j0gs3gp7eH1OjDbx/Dq0sCYQWzlY3rxL6stZvYdTPcNFzMF+
HpgNQfrc/DMkVjdeyB+4Y7u8k0xy8HFZOCRpkMN2PmvF2gz/G53MZ6NXF03z/6AMgPjjumfmtYqp
x/a9OJ1uS8EFHDfXLRmu9nR1lb21hhIvm5Uk9VeVEnlfIHEb5e09nGHkxGpjzY0QeIPX1L2YiR2w
Lv22Xjmm+W0yqc1ibL2WAdsidVJ8vqCQnGcK/5NC/fvTnEJWI5kO/EKEJW6r0ai7NCh3obuwpwIE
iAq2bPl6bJIXOicIOBRvf3zanN46CLAUl11P+rpWk7uvWy/bbWbnBrHzOIvIHTayWGRqLfr4Y7xn
1jH2B6Z86qwSL+Tbl3uRs0mGYCT45zRWUra8spPNQ1ZAWQFp8yJqVjM6ZoXLJ7k0E38o+cs7AU9T
7hRbWyVCSAygl4lWHrdRYzW0ZBD/jtsus9Acl9jjCEm5PPBiTm+gZbAnYAusVu6z9X9LyEaeoTyU
/v+N78h9a+klWK9bvSULWYWf8a+9uUmeHysSJoJJDEToRR1j71o33cEbIiqZriv5CbevcL3o2Wje
0yNma98RBgGOf5y7Uai5zVXT3CPMLtY9aZNEq49TVkAXEBtBIbMpUS/ro3hyMmnfx8pmqsqSohxR
SSLPZ/sDwFUUUyhlAriKkJuBSNSUKW6ZcY3rJttrgo1FtbGsFYwoaF8j6Ll2iNMsKQDVAL64XopZ
ix5LRms65ro+9+UAgpue6Kcv+xM/yJAGmr4F8covMfZhMmXSmAgDssK169j93uOpurarMUm+ziuO
bJYNxwFT56fQ+ws3twWTz/5sIgCL05q0CM5Xb53BvIjJFYmy48iNKLv+kIF4j2bhfsKst6sTPlKr
PHQ9kdGWmgm8vosfuLyVgC5OSi4QF1G5HTY9kqOeo44gX94hJ1y0vxagoo/BfXEZt3bG4aUWnvqJ
9V92MoJQFGjyyCrfz534nP8vknqQMxj2HX3HfM7lntrYLQpZFW/GXLZS6GzEjfkptnogBAZ3Zux+
L8DhAFO4pkBcLEVluBr90ZpvaxVobKN5p0eBZd1YYZJcWCDGAAEYWrpaXsx3RyCTtVJTTQdV8y7b
cz8rXt0y+IGmMQG8rWLn9MF6avRqKaCjYuUNpAaWUZrLjsJlnJ95GJyCGXYzyoclh0QY91WB6YiA
0bk926ACb1VPttjNTqyVNO3K9r9Bqv2BR0VMpG4jv9XM6lCmFRNXvtxttpeRbOG6XaLHZEIk2Ul+
ZfWytpEcQ2RSmsqR6+SAE/vDnAUVglJQ/rAIRLbQHad//RHw1WmS1ZIMZ0sqH4KF4fvlqDfdsOvh
Y61eRbcVGtVJGjEoKfASEzdA45jl0HUBKeaaI4G1i0BEu0XFv9WY6OuwKO5NSinT5PN2o96S2eBw
t4baqv3RnvKZGt90DFRIR1mVJHw9x+JxgyVVPCS+ltcni1Nir7Ys0HIIrkrXkp4xWaDNXdW6Co99
TY3RaSJMMEcT8zn6cGG3+crgPDZS1mHJJvA7b9KChVmmnJZn6xRNONuqqCkG+EqpO6w1hK5xR3dG
wdsUAEfhmZgYjo0jwfssqhzH3jaxy5rRql2ZO36iY9jOwv2o/ZQXkZd96P86cjUdnOmcbap6meaj
Sk3BIjFgKxyP2nbtIgfFMWQl8eSSy3ZmZQbWGI0rAJQpAmAiH55V9UGX5B95asw4/jmeHfeUB6Gs
+64JpGYRDonbB59uwdcRp5ho8mRWPafPNZX5sUpgtmgIxVMhS/WAm00ZRIgVwjwSSok9kWxejeIe
enEiYhIkX/yMGyDF6Vlj7ZLOyyA0f6Lc2USAJVORXB5Mb6es0dmC4qeS0AfEERwm8DHHJw7mbQSU
DXRnEBQLMjjmrK63ZDsxB68Lx4n9M2GEUuU4fFyK1/IYv3UEvANAtED6TcW2VD+J0QuOLvCcwwg9
Y2XAQMtLmpejA/pLS8GGYY0QfuKjSDr1bh+Of3JaI6IS7JgbJRkOkYlOGW1UStESZeYUHf2KzUCK
BlWtvA/zXdNPavc0W9KbMeniXrckHHrg0R1eCevtGojUdQuOCGDRdDD8NXkkJmWXdpI5084T09Gj
btS0MJAfWPvtJh6Sf7watKK/MYwIxwZezR+TkMrySaXlNzhE21XZB/AGq/aoeRJxvHjsx/UXXMtJ
RDvuY576i3SbRw/VigVhjMmYTsomy9X6Nv1aUTGQI0ElNwahtbFBvClzoRrThTV6xJoV8ivUpujT
FtmBKpf5Ur7eX5Qqi8uLbjtnsB5dgunLHKDdQ2ocooo1CvbFuL4HPLH8cT4wstx+JM6hzd3ZVn0O
3RCFtLGLY1DZ4ffwnQyxdKX7COn73Zc/QvQpC2T2ClUQwD8TtI5xMDmCFKG0xRcZriBgFwmqaDfS
Aw3J9qwSKg+7z0h1QZ0n123o6uR2U20g69CppVt6c6rtG5u3+z02nSTpy/wEzcYbucTJs1WS8F/4
f25S2Sc1YWTAv7m4Gxlj72PJxJHpc6ZXgHG+sKjUtXb2mIubt4cEAMJNLvE3UIJBDS4OF5HvpDM0
AsA1/2MLtRftYcwaQQBJavVtx0J+JBhJfr3/TkPnwMMDy6r340S7lxEmsygY+PtMvXTeyi142hqX
9UxUqHzP2nL652VY1yDiaCebr+Qd5BMi7Bo5B0bzo1DOHLKuWDOPMSoj1a7DghaFAcpqEFMCzk/4
P7LyScUEWK1l9Q82RqgvXHgDSgyZKAirBo16LmA4MqsXMERyaaXqtpnPbMWTYBHZJ/arKpQhYfZn
iiid+IILSKl8QbWbAFd9OoqIGe6D6OIN8vw0Q6QnyWyqGidnT6GZbafGTV+oaIuRIBHV3iq4WZTR
3L378tMxu8XC83r3og6zOTADphFuf/+u/vySPhi0LcEA5FxtAHa7DnntQvkuE+EcmLelWriw1ck0
dAZTUeodlLvnFM+/8+wMGvs035xAR47pmCH7FZysWIQ2wum9jrVdJxGnQZ6j8vsV87UbjXE2XRBy
nQVn5za40MYyW6tFzv88bBGHQE25MilCVBn5+L/vjQ+tNmrwweBhy/DK1zZW6yl8IT0G3hl1QUQ4
Bi5KC8Mi99HMnyOW5DJ7SPgHVnGlDCuFHEfQYWt8MFFYyY+MW0Df7Z7B7kWIOPA/1m4EdRCzSFN+
4OM2edu3QaHNP1HPvfkMBzhXTrvs5yJXWPuyE6xJUNAf4+cEPjnQ/PXZZT0u0SPKhKMmbSJnk59V
SvrHQN+ohR2yv1jlfSwmlonfqEbptpcNfjGvWm6XM8y44GsgH+VHds1Ul4WqzuTdjpSKPxjb52Nu
9XV3UZQ6O1JMk1Q6ulXpq5vhyVqRUNqTzNL+K7/5PNNZ8X9zXgxc1vgRfxJ3WDIXmwKY7gjX0JZe
HbwD1r3REZu1fzPhnYd7OszFhlhPw9bIlc0znkxUoghyneLN/0OOHXs3MrvSDcp0r/HL8IT9KkG9
tjfW+zE6CLrwmslUIQQgVQci87pDQNM6ZKcedKX1onz2eJg1sJtt4J7GtmrdUAShxkTPDZ7Ozd77
gtDKwpggsjD4Lam7NwWHcoNI7GztHZ3tooggZ683zEEjHA+JQXh8QrZWXfpPqiVA8+ieymwDXnTl
iru87vB5F9GWZfY+MVv2jEUE59JzTlb2R+UvHHzdZvso06H+Xlf+Sh+KgVBdDF+V+eKCbBqKqTG2
P4UTB2ZbuouiVbkk+Y9QZBLelZEAmziOcQqoiGjvfJnVwghfhCLc6y8BXZweb/kez2l5AxIX4zoN
2Ok71u621jdDXXDVpKh1eeFkyZ1W106Mh+KPRa2Z4SLxrDmQlAfoPoaZnUyN3hSKk3cH1J2/+XG8
UCMqxzQKydnoCisZUvQTOrSiJWLugGBoLE+/rS2BR7dmaqUmC05pNhg4561YacQSEXpWDTTUxmop
4aabqWq8iEJZXI36FabOqNmGBPRV2BCqcO9XWVHht/7C4J9oe5JL9o5jXw93Tg9Ph62513XznegV
RqSygq9DailCRM/D83JKX1QMPt5TMuoJ4SNtt/CjBlouHQj/3zbfcmZruTpActao67s5we7T8o36
Z8Ge5vyxG27rTCnKAeDKS5aDlg7MR8Etb5RYXon5EbS/PY8LKUFGWLxZd0V5ZOFM+v5EhnVQlja+
7a3zgiStdYcBmcrRS5G1BeZEELnfhLmaDV12ZeVodGQIJFRVgg6nBS+PqUDK4QrZsRZKpwC04dMa
GJQSPpYbpXm8Yq4hy3J2mO0p+IASyZUuHHlDd6lpTjftvTz2IshFe9K4a4MO4kjDoy/oModJDYsO
1YGX/6RlI+4g3fjUXMFLv3pq8RrD3ODFn9oHDeRubLe8OiQ4ctx/KUiPqHGOaxzltMe64CS+zlvs
ZrJU+gUQZn3wqqhKrDHf/j2SjfcO1W31TVmtiejL91buPYdGCDpkHK32pn4hO0d5TRkY60dusS9X
aIuZqOhP/IhpEFPIhj2vE7YpaxClh/EcdtiNPepq2P6UVcJjfd9NhF9qMqU22DEymSWNzW2K+OK6
lZJBgaF6S7b/DZGWGvpN6Fee/766J9riNSSEgJY1p0Fk0502wR7/56xIa9yUV8TW/OcCD/kVptY+
7YSgmo1E07AOBewBM+xWCyD2PIMNPr4VmStOUrX5Tx7UWrdc36AJ2RQOzE1NTvuiCZir6nPnZv9F
PtBFrxO3drwPDCFyy4EjFYIweowWufjF7xAE607FdCdSer8RhEWGpaVW7k2DLJ7o8jt9WN1Xjl2b
jdxXJ7QqTgjEpQNMhvHzpU+ckiFvTBuBrv61iMs8qh61il378d/PVj6pOnaUX52lDKcSalPUesK7
jm97fsOC95If4bm5b2jgx+8OrmpK0gOmejVuGKtJVSe3vMqVsPcLd22+1sIBzeosU3HOq21viX3J
ouUNmQ9s67Z4FM3oEdwlezUavnpUDkqkIdQKBf4MCO5QKqLkutQ3lFhc636Htz4xovTHQeIUNcbe
l1+giyiE+xbu/uXX/KWo3A4UPv+ZuetLTv9KirNDgMTSEloRlJQN6GzvDh9ODhZIOWTTQTF2i2aT
tylrdpKtf7lK0dR46neBzD0RsMFMjtbOWOaXTc5ekyQ5CtfR1WCmuSdrC2l6tArF4ABMM2Sy6DuM
zW0d+uMhLKZG/wgBLgkWJXNEnq7QlqgBEm35CU/Q94uZT+YtqBAcLVoi6AMD6kUa0cgnUxebgtOo
wlm+9Y1EvYoPhrCHqwELWgd8FN1zoNwVDHI2TG39JKeYFDeDtFZj2GVrfIje2803bkKoDkqpGY5u
uN8sgGMHJKGEWsR1LV705T1RMDhpq9Ee1eEPgZ42Nqg7fwCaL4mfRi8Im6HrCkDC1Nc6EO0vzMvq
vsCcACm4o1C9vDSVJt2YaPEHRJfSpHkPN6ABuNGLvsFLN6cZ4Np0JdhEYeCK+VIMLCYmhtgEmxUF
hqg3PZ2WP0oz6w2AyqAwqzB4j3jRCKH0m6ukMNcftKsIPIB/4scykHrHzYD27Yrba1HA+aHIPXKh
Pay9r87Izx2RdlL1FRnm/+4h5Cr5fZITqAYdVb8QmzQhjwM8KmhJXpaWmKTwkGP8sxrXfo/wtW3e
2BHy5hFd+/oosuc+EsQopfQzl6TKs0GWVEQie0KEYWX5sp1jp6WNi0FvezEGdl5bUvhBhFYd7etp
W095OwMRuhmybAU9BzD91uWTX5NDw2kHKlgO1AAKV2w8ztrC9dU4OpXrbQYm2wJEWtSn4aXOdLCZ
UarMiSg3hFHl5S2d5x09l2+I7DdfFdpBLj81BvFkPwTnrzD59pASoLs6E6fsgHp3ANvoNHlTzHtc
fNHzuTblQog5ZLN6rPtLMlxeilQRHkupG3olzPQBf5FBLX1hTgH5qznm1S+xfYNNk7PhQezNrUPt
oEgaDNe1V3F7IFYOsQ+ouaQWdMX8Pdp5ZBiIySXnGDK/oN/xfI5rk8DQj3xafbMJlF8O3y3OyLJ4
Bj64n0KdhYCGDMTVAmAMVYLhXbp9lH7iVe2NHkPrPkJ8gHQ7nOGeYZhZpPD7YTooh3Nm9XuAL0+N
8pv6V88JNHTnIeC+3808le97GmCusWLNc6pO89Vb9MRkDdjzfIidsm36ENIJg4i1F87WNyGHmFlM
MBWqoFFLsPlfhnRLgRi2QXdPfVyQnTcSSUzEXzTgBPy7QheUm3RpuYJnqa6UEZQe29+ZS/sIoAfL
yB2ZnEBNuknQ9sMvrFdREUKH3P8tX1dNg5U0anjbp79HXzXrLxr8l/vsP92TRxi81N6MMUvpfyBj
CJHHM9EjkNY96nw37x5j6swYINq8/pWjhSWp7JwITmwCVh8IWxD588ZqH8Ig10xDvvKtfhYqK/of
DJXmYPfUoCXQci04PJlZD3X63vDf7dwojMLHJbKoIXU9c2i6FY0RBpDs4pxorhZpR8SEqybioZtP
/MkPNEVL7nl1pXDSsJ1YQ0IDhmQLCdDU4w5U8B/GC4/G+j5lxgKR5Xjv3izvMCFzFFsRzU/k8ViA
S7SI3SaiORNBH9tlSY6P15LhqcX7o510QPkzPK1RiIMMacK1E8PdXtQa0lwkvvknbBe450X8ZcPd
h5Y6kFiDMGlO43JTkcy5BxcGEXgv7ISsGy4FlQxKZDkzBNCmxQBOnkYxigL5mnsw0jLPNgX5MjCl
lElQeWk2gh5wxIprDUX15Sfc6PXqb1ALqH3LED126YVtRxrU/nIymlwJ0Ms/RNxVwfj9LZLSo4VQ
Mcg2WCjr/TyTgGWe/jL7vsEfYMm6raMc+gG17LI6DMkc0SoQFzfeCgv6/juwWf86awpNxTR/A2Aj
gLhFh61BfbgSRAuvJFyG84AILDc8o/VL5Xgn/FTZYO6wf3EQqTRQ9GBxKt+O1ZwfYikpblvI0Ue6
tXQjkMvzL/juij+Gawih7E6atTvpPsXQmqcv81uyOxCOtKeV9Dnq6rS8cx9RtAttHAg/SdGdhm9A
t6O2OTMv/Od8XIrZ9idQF8rQpJsA9QgNcx7MSEiEKpe9Wj0hFhuoq/3tVBV4BDLPEGHpdVuDeiBj
CS4S9g2nQJWJws9Og2EiGG9v1vjpAouMmeYe5/C6PGRRTTCknsGMNcWKRrG9dyS7F6PnSVGmVKXK
+2CeG515TXd1wGM+6M+cPeXj2a+1FLo5HfBGRHEUOxbbGwqDYJKMhGEZPLHzLiyMCza8Ie005/jF
5BJEnSQflakKJJKV10OTn65i70JwGWHxxb3k4QUCV5Vvv1hJaxQoN5L6USqf6UDs8FDRDyD6ptQR
MO1Y2ma81HqXeKhkL82/KxrK3nhlxN68EszJV1rwSNr3fWcOwgF4WCUVi6I9ESP2tBvXgxPPYPpN
KzQY5CK9ZgHYEALlJ8BC21G7m2SQ78R8Lnnbt7FjUWPCUPhzUGjDe0GWbaMVGbuVi+SNu35MTav/
5xb6SsaJHxi34TRjJRx4Iy8vKbmi4FxZcpI41I8uXbgSUGUImFoF8ckJYhaQkzWQyHbBjeTXNfya
CqCNNT9PZSYZgq6tkKaFXaFtx4o2FYgjrFFghiCg9YyBK9WimDis0sB1TaQG3HEjXnAwJtkF0fAe
3YgtYZNQdrQ11uyvuX3/KBUJ3X6qEjyXZkglMwLAsrC7oB0CljVXT9nR81pui8EfGQq04mHLM9AJ
NSCFLXSTIJ8bkiCJA1LdepgxRLPAP3hcOv5qfnIvZqo37/OA4/dsOwO9j/BROVXc3xYQkOk4QXa/
8zM5hroMRaeQop0MSy0ycazfR3yAJIRKmw5sH4cYJYa/3aYg+7wn6czZiy/hAVY9FqP6ZR2w+Vte
VtLl80xilLg9jx4HOxoTBK51vUsQ/Qzlcp19xquxHffd74YywII5a5N3E9Mb7jhUrAlp2rC5OLwF
kOzFh8oAc2xLacDTJf9P2G30983520bWA1+oGXN5DXjJFXfVKLmoJZQk/KKrdE7QgV+2ctq00vpA
frc9FjvLnknx/v1Eywhv/VJeiyIqKkMC/JWl1xDezRBKXm4RNR/6hlPYaxY37zhob/Ei4vQob3BQ
SK29xCFQLRJPqBxtwuKIEYDXhMDrJckaEzDQuoDxYgBbugldDqG9DytoWmIf0or8M0Pi2kVAc75q
uHcWTcaucU6KyfvIS1nOYDpn/fxdkWazHd2YVkebLLI/2iOuWeYEXCu2hfSzfT3LJnxzZl4fp9KH
QIYi+O0CbcbA4ycICYVwZOVL1o/BhLoeoNTM2obpgymlvkdKXkY06AsHVdWMKa8nZO2ttxjMWbZZ
MccM3iYvW25beWXpKBpMR7zhHPS/l248ECYLwwEjDzDnfdNs7svqjvgmG9qzIgY4CDjBYif8xoOm
Xx7G0vGhBOXPUORbp0BOlr6YViB9vykiTq3UkARbubA+9045Q+f7viaiw8xH01UYeVbYO0JloZWv
IFFxcrRk3c2mJsef0VJn9IjJrRdjA9cWm1++008G1h/T9FSQYgAl6SpGVTd0/EjcKmeiy64Wa9P/
fJbs70eME51nA6RCqFtfSTeAXVf3s1muBuSfqLcchIm672vajGDFk9fDDk94m8xor9cl3/QpUCQr
nadt+tCEK3NnPWkTjtGXMmvP85DaUJxX/mR3D1OQ2TnLW/F88yjOWtaJlcFvdonIY2ki7/PekP3Y
EsaqIU7w47xbodZkAn0KQ1DqmjIBqzEy00aOz7lDpIu1WjeSxuntlSIsSqScQu4kuBkJ//oGGXaZ
1gMXZx8ijK1Lh5IBxbyHifpV42DKIF2UqCWtqs+RaQX2+4ydD15DP4zXTbeUb/Vmh4Njq5f7GKy1
a/oMUzbLAowwT3Y332zBZqKK1EnBGr+anvxf/Hv036fnBNq5Zqf7VtvXBHlQ0wFl4h4OQVEKlNQP
lMexdUAgBAkDx85YCachUlHTO67uBxnTwaKWMp1vHxZgNgRBoZTO4KqIS//yIRn1UVjnQnZ5DQiZ
D5F+3i+vIggcfmYIxUMcClYv1v+nyGy5+bsljzjzFJshhW0Rq8lN5Jnz1hKXISD3uyxZ+Re8TLOR
RlOJqze5jRrk4vedJZMW7o4FNEgZ3s+h99mpp+LCav/gPhuWYcUYqORssRyaux8DFhRAA6OZc7Bk
veiJciZBSAQNXwrzLbViEX37ysJ0CVuf5alvoIYX54Hr+QxXThFM9fiQuL+2n/EKmLdnTasEqn2y
ngd+mwzbBwjcomktAgTWK7Wcb6mGb/XiWxWgxsHjc4e4Puu+PGlEHpSbR2g8ruGjtEy4A5klPiyu
6BLrY6UsN3jNr5ZQOlSQIiK0QK/Q5kiW6wyclZDvtAaZTO0cOG+2GfijqTGODsYWTGpJz5xbuw6N
+kXUpwH8dOdcDCeXkZbwxEZUN4Bls+MB6GBZoFBYT8GESn76sL2tt3B8mXNpqJnn8nRl0zGYxH5S
26m1uaV4S1X0krXsgf4OVUDWnXpNsQiyS5JitOi/HKQmk9SrCUZZqrWVnpa/oZ8NGCXSxgkGUaQd
L6m67gBkSsPhLcV5yQKOt2kF0xgcBTcMsJKDlWX1aCgvi5s4Osd8zC4ssLAmbIGm3RdVKEtV3pfA
Zc/pHoqTMCJvbQ17a8vmOwbZRlkegnn/M/cBKnLn0Q970Zn2o+15fiW6OYb8NbjUR/uk+u8dIez7
YzRGyjuedbap+EgRVSNQrZL8WroLat40JoFO6eSJ1IT9GIDjGpPfCA/3UNTs7mykABLPtLQlNg8S
YrKx+oUZEFKN8YSZw6SMbJIfPw4AxRZhHflkaDA6dz+w8ZNqOvQVQu3++hR2snJ7Gir++1Mme2fF
kxeLm2X4X+yepnMIkjq8gFyZQy32eSOb34NSgyc59Pa/PcShCGhWRNbGNH7pxoj4poKGsLJl7uWO
I2ZElur0KGMS9/g0iLaTdGwdhM/df/ZunHftkf0PQHU3wC4emQ3GBprW6wVottPJPbQ4VSORZGdl
bJ9aMGyXvqz7onjgraF7La7hH7rM8pP4PpiWUzXwEaFfWJQb/KHXyFa50LiGmnLQYEKeApzjPvDK
wQvNLty376xGzBLGaAKa3lWxH/UnObZDG/axnyHBeR8R0rP9KsSt9CDD3P953qgM5HaTf0P06OkC
4U+cqBOpjUz8hSvqKYwx8bwe7pJ5UEBTmBev5I0GUs+J6weyYe8lKD1ha9Xk3g0XBuo7/aPn7OEw
feAJNdsFvNoRL0zMS2zlgulW407mnh+G92EWPrY0KTHCzo/zMXk/HNb2Mj6owzdZGSLVpO5BcLB0
2MTr/POzrGBT7ICxcu32HBXYeFjE24cj6bZxopRNMbBCA00z0Hh+ImHrtwWPnY9ATTKlQry7MxpX
/zZWkUVlB6bNsPNSVk2Sj6xcZTQm6FMgIksOtVtvV03JeI++O/fIFUmoSjPF2QQv/oLGPKW4sG08
KJ9nh1EPIwyuChz99irzNArAMl/FCOLoWfLsYdx55fGxARY2KwKfquFHEAsk8QqyUAytcWyWKbwG
t5ZVwmuCFArpIdFgEzF6WwW1M4y1so02+xAJEWETqkx/3fWQN3bx48C9o0InuUXYhsfn06ufeqSB
8ZrdiK4sljCBQ5RhLT+6t7AgNffFy2MGIpk9+xWLF+yilKhjxv3TEuPhoPuTrIekndE1bWGKuqEt
6G+THJnDKcK720ckgY/Dd5PsJR9wfFq+vugLE2E6RpKNS9w4c3+jE0YoTdHkpwG7X+cgBGVm8hLS
B5zER1G+cABTQQalnKSr4ggMXTWJzC4gOA7OKNjyrVDrpJE3XiSNF/5bsvMB7y34wwVtNQSLseEW
MlXBfp/KfVT4vXf8sqroRIcLOz0j+M9HywU+7pkELdZswNNJZ/O2Wrj+FQDVN5cHTqONvToQlZ1+
D1GBlPjOfJzzYcF12zqlbFqsrFWK2b8tC3r1+isiXguv36F/VrGRhvdCXtTGI6GhXS7s77F4MyQa
0zJ6HKocQTVK9wDQY5XHpO5XpImRQDDnRt1XkkTPvE4AhznzTAf4/mbkcyzmXkevoKbrEg4uwORb
DAUHCpQr3Zh53UfbfjfvaY/KxcD52VMWw0XY0bhUGgNUHA26EdBqWFFCa/91ZoWXD4TfuxEXT0dH
ilmuby+juBtFMQRDBGeTDnkZjzU+9kTbXRGXQjgMh0y35ekfs+/q5HlUzEP2iH+qPP9Zj/GmWTJi
LJlK4JDnpWPv2ZKXvkWWdrwDmH0apq3iXaKAzvyjsz5L4nDPFwG7eZtTh/cpNegXRwiEW6PcUDLX
Ld7C+Ep7IrHCCY8p4wR+GB2kfCEx0FZ7nnAec8la9tWZ67qNy8hR6m59U+axuOH3yCNqX6kE2Y0V
uv0aG50fZRToipguOhdoQFEIwCWbcY/TGviH9h4PDN+fY0av0dqlt+my96la7PSET/ermo2SwGqq
va6DJsWXTmCrmrwmG5SfNdhDEh79tKNA/bO2xGuOUi4QbiVjlGYJpxF4yvxBCQhP6SNZJOpVh1n3
fgYsAD9dBoZAweys43tLULHa8qMUreXXQy+mm47q2evEPwj48vYYJJaLKV1cMS1BhNgspb/wy6uO
RPNp4U+8OmNZk1dkwOwCoRvOCeLJqwCtfj00xISWd7OSOBMarRo7JavhirZ9hwTr0lCM7ln2WTZm
EJkTCgi7qaFYWcu+aU8sxmnzm8+cqzZBXFv37p0K64rRoNB2p9i8d0V7BLAcu8tv0oB10J5xoCVZ
fjIhdyPiT5+wAIu9wzKmzWiXE+rEyk0D7HqO+6vrxnguynoYakEMVdhuUYo9YoXQG0OJ180Nspra
iCXuBK5zU1UAcO+cR4txBHKbgyujt71SBEDoXHof46D+RKrwgvg2RGdCkPAXksXMSaAhkNZ5u9aK
Q8+fgb1MzzhYzNynNTiGp69oEd4d1f/rXOFjcSgtC4AUWHpd0ayHbJBqenCdwl61KulvamUjW+wr
uQk+xssktfzJmIeMZ/h09j+gTGYepJCGP2sroIBoXQcIgsnkufR8pG1ew+2HtS5Ni4qo+J8alHC8
yiNzPjJUqEgeTNztInsIvfIBd+OjvLitiKSGoAujv7CCRsEy6zOgYEz0hTtBOaCUvbwh4TM/b7SX
V269E3eIPDLsjZehbSzTL8PkxIG8IZAaIBIhL+dzEupyz30MsWZM5BgoKXcja/LH/Q9IBRcIm4GU
h+TYnzrd1WfZbzxvQZHE24MDgprdicq6vVV3bPnQFDUSwspEPN9gNUdC9lo0zwD66PogyIbb2i0I
rRDPcxOF3Gppn0XQx7A3ct953Cu+iJEUfKVIzRw3axy8BigMHJDowlzv3WBjhLbDKYMv9VU4oEmX
WnN+pxbSKmfNAgC1HpeXityWiOIWKpDt5Gx2WjNc/zVjUOaoAev1xTR5bdr7YUvx6qPypYs1yU4b
g6G57mIHJ2eO1OapDFYbihdugcfpRPXfrLFd8XNQlDCgkFgj/0AeDAg6YLe66EXMgFhgehV7KC1e
y0Fl8oruQ+lPaGweOWQXDNa6d3eSik/k7smnXBZkH/jXl0yfcoyrQQCloV07Qqda0N+dF5i/47ZC
94wvoeYsJzN8YcEg7T+qBR5JhWVNSNfwnkEvt8x1HZgeXgX6Va+VoRJ+gKxyNTAleJyPi0yZu1F3
3vpTtbIyy62v3P82v9IgG7v+l6i5hZrcYN6m2+6nn1bNPKtF6JRKEOfj73tHYSM3PC8xxHVeikz7
5Sg1sw9zugAx+SasXjjOFc/rq+PaZzVNikhSS/0cMSRW3GOFq8MIm2nqGlIDKbifMg9Cd2GYtyKM
aQl1YvnWYeE4upM0dkRv6kcYIsr3DSqvEaDSK/U4k0vw0sA1OGwU6DSqhAtlqPM5t/7WWmKpL1Fm
jFfDc+vKAKOKF3oHorIwJyOHYBcBvCKQySC+xDYCiyWNH3ydhHeE1UmgvpEAXLNBhheHOgmP+Ae5
Uj+47c17+M+mnY+Nw7nLvMrNNKv0DgNGPXZPNiVhhhJdzx5Hn8fjWCPa/sc5/0bMlRsasMNl/Npa
TRca0R3SCkZcgyMQ6mLguXi7DWrFQzMtFsYwiofXmgJVKQQ+3GeBiGJ4q67lM0Miq1UF9MkL6lPi
ijryyljZU/N7jfeWUgkUIOOCsRpjZTsVnMUB3kfN/plUHXmyChrQTWRakvCCAHNoWFQy2EWFKq7H
YzrLibMRYTQQw4UAk3XWFfBcUnQ6xWjWlUQ7nxBfRzq4jWzPBUVW0YmPuuD04P2ZpUMxHuyvhEt9
E76adJpPjAS2sFWYABmIibvH7Xz8insYYC8HIPQE7bhqJd+h4qLNMKWZcZuEfegjS5lxIwMVVIX5
qLlzKFja/sHiQJTjEL95NrlMz2piTSz2jy7yU/vrcPAZAwRit+kZqhvTljPoYZk3K+hdjhkWqyNp
Fj3ajKnEPmvleV82TYMfWoYpAOGJiaBJbGp2sVw4ZfRWyo+cUnFMjrWhugE172Mz3237lh/umjuF
r11KwCilG5B53XozzIgkdCIwfExWC4W98LZm+OufzLsd/PbiwrDr+CH1JvDWDnZ/6K2wF3azyKUG
KnqYOjer/d8GVbSjKBI8VWSdPiGW8O07NabfZS41fp7Vw+r5NpB8LLfZg7cdgdRYc/gJM2vM8JlI
LxzkCjY5EJfMEK6J5O5UwMqcaXVw7cu/qa9a1/IGkKFqEKdKI1Ft/LLkCmuii4I6fhyUrDYTmRSK
W2PYuX1pnbG9coxZTobFUWS9UCOujidfjj4Nbbs/FDx8k2BZdT9JpkM+8Ccm+KOmV5PT1F9AJ8ml
RDfCErjCE9A93cXRaEBaGtn6Zg/IbGtcugkH3YEdWuexQW9EF1EFNiIGoCRfzaLcok/9y+LWkM3i
Ap3R7il9lXCuqEOvrlEMzl4vMaL3qaqNExGjLG4Si9xsrDOo1X/NXp/i/xVAY+LefWElN47Zp/5o
TBIDcdhM7n6CnJaK9TCSeFv8CDKMQ9Z0leWxktTwdrLg3hBno2aEQ8IdJHLO2xemLmR5+0pSr9xG
k93OL2k4yyFnHVmqRC/PaiovDpDx+HwfsgByB5Yh3LMwTkKoH0cesz4mJyn6b4enbJil557bOeKc
axVhPci+26L3e9AGW+9GxYf9KcOllvuvaRsMikrjAt1SLETcfJ6pknYN62/w02t0ncQkPz/n7c6l
M4SJLoSOuhkfZZVit2wlwT/5CF7WVp2o8VjYEaN8bW3P+UFgnA8MM0L0+Vq6rt4adU9XYm4K8D6z
fDy+np3/T1uGKMKezEXSGolQqHSYLQT3TYLogL5ImcNdS5QvwRgXQA4S6tt8rBwHtj5/mbsN6eOQ
N4ahrXfRMbJT6lX7qrcV6gJ80I+/e+ed2uux7KynymyCVgtCRvxKLKF+EdR/gzTIJnkstLemhnUn
01BuwDTKSRcea8b3DlXGMh0TLC/M7aR4e4vFKSUKy37s5o3u5LI+Suptcw6ybewPT25EAr6cQZda
h6oRUsE1FG8IwllS8FybNK7pLa5aF2XPTusq4YgPIZerE58jRZYcp3K5rnbsCu2ohdsJHjv5T/10
0OeU2ApBKfFEsPr70T+NREWnYU23kuojhPgZkq1rtqq45pXnlyHJKPxZRAyErcbTulxl5EgysyxO
s7T3j0ShLDYi/nU+z1t28/AXOWJ8LCoru0xeTzz+M17NSvkNEJsmRHSodAHV1FFZxhvabFkwQcJV
wWRCBCZ9OKY5vAWwDoE0IvEoPTfbQkEfPcso/w88ErMHt+a6wr5mXrabDbH8Gn7Gzl6DVR4RxUmW
52o2TXWhEM3K5iFJcldBRkGa845bgpdSFF6Y8/jN7fN4mglf/iJPjO6rADsDLe2QgaWdC7g2JLoc
jkRtYVKGWIT6r4/IvGir6XbJChrTid/7dOpr2U+B0GmP4STvza3p7qTFXbsDRYvXZJYmgOw+/Dn3
ZStFp4RXas7Z027yBEpaPPdfUN/1RRqCwzszL85SFtLzK78esNU/d/WTtUmMynVxScaP5znalfQu
HVhRT6GwqvWIehGVOzrokCYuG8MZOIzWdoAXyRj9zrJNAfd0zC2k2sCRKU7BCFe04p1IitidGksy
iJ5jwDlyBqhwfB0QB/Bf1W3IcnHG0EZoyGXxS2slFRXZuM7xN+ZeE0tqwMuEjmK0u9/yiF891dQ2
rH4ci6sWz51N/czxDA8Cxsj6h4ZuYDhDE2uQ2jgGULPOvChqBwnZ8L6pxr0VN2Tn6UR+Mjo/zcbz
OrWVuR6gIsvRTolsA1gGcllCkpE0WlIfkMDcDCFBLDplGdb7jvNnLquJGBI3C9GextrdXJZYFteq
LBb++EjgOzAVcG5rHWBR4hZF5h+TelFs1JTGtuQPhBslyrMt0iymp1PjB2VNhg8Xm/fMf3dWS/FI
8KoB4TsMZ3nQuAUxG/1O45QijCysFRL6dxncTTD3UcuK3o4zuzkjLBY13+6O1t8cVjoqgVnHWcZ9
YONlAq1DMtA85rJ/UJUVEBYWLcyn2GXb5HMD7eVhFpthgV/Ka8lJSujM0ohc0r3aUjqouQE+SEg3
k1d4vFODeZ4e5VihbWAC5oM1UThaM4QVsr6RpLNnDCddKJ8s85w1CWfbR7UO98e4Q7hpBnH1gJE2
3RDK0BQSy7+Y3ujjvXDsFhjLLXoQ6UVK4DWCXaXOTLzMGUJQLGCl6+aRZ/hmImqiAxLeSGxdTnA4
XDxYc5M/PEWmIqSJWhCmX2QPCS+LYDdWToKDUIoNzj69LT+FhpYTknwWguXYXCaViKi0sEaUvIsn
cea9N0CHKmaNqSVWvLZ/xPh3Krq864VXYf1C7tp1oPZrWh8jk3bjMFM0bSUsZy/LQVuXHmZftJTA
5aR6juIXlo0AX6WZntRYxmOilTTBxXUqdKQob3Vc8D0p1vU3hTHf3FCTfolqN9lxcCkqeFYSdrVE
WYX4CQqVixKfH8L4AgTAc3GGA3ssJDtOowfHHt3mENtmzF7uF6YHgw7anZVvz3wyoYDVffW4nUw+
Qk0dSAedqB+4eKZHJDt2vt3wfA/SNqTlTar8ETB/nXxtyoe9PuCJFmpYqDfKc/HJshdthwRo3vYF
z/0o1zXyt0A79gn/fIVkaeaIXBBrb/puvh9oHtvKJQ9fqMg4soAn61fFqjT5nN4uC9RPbNhUyM3C
h0fli20XraMGQVfYQVghqgRcxsqPJgv6NT3fxPNA3wyJsdf5f8/cZTvr5lat3LXn5os6XX/4wKKz
A5MC8nuLocwe10zV9MaJq8FAMyZ8NkED+PLqCr+Yua2ZRCOtGdHsXOS+4FxFQ+z86PUvyVpdG919
un82gei5YmfcTBojjtLG0spNXVMUe/wdXnToVjfClHH/qTaKkTJmr+8ASONKozgR5J6STIouP/Cf
XsbQmp7he07JxedMnqN6oag0nY4UwNU3vdIAJchXwMaXnvpysH5n18Mf7PsoJtwqLWUC2pCmJlrj
ggw+mZTYr2jDrc7UuUEkc6XwNHonKTENmQ==
`protect end_protected

