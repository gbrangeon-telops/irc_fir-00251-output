

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IoOiz+BDpEiCAzehQDaKkNxXycZX6DxCheIbVmZVnOeE8xp7Q+9Cdt/GYV8eq/1L+MpdyADA71Q+
diEx2Z9pJg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lwiDFOkaG5HcqeigSQ6a9WNJOSnncyPnebjhd+6IKLZk0I0Ny6LWNpdm2fV6AG4pFcvx58T5yWEl
Q+/SeuKD0HNAWdTl0b2fE07zxr+edW2hoGXyef1M8toS5SeJjbmVYB+jYYVGpq6G4uNelAjC+U6H
qvBM4HmLQCceNGUHSWE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UFVaQj8UYHzOV/s9ci9b6/M58BwxIhqPdXQ4yEijf72oAEn9ivW6AsDsNzmhpHIiBklSohpBNUDU
0Mva3SAcsX3+9Czy1ShJ5GBV/GrTCNonRWGYRXu6d9ADAsYZRaJCV+2s1kEifAqI6MJhteonJeVq
EumiTmv57LCQxMW5bGdt9ducpN0oI1Oavkx+FYROiHKMHPR5ux/CzqaZUlRJQvJOcmbQcmUZt3v1
KBK5x+Z9B/aBdtf5Z1OOegRTMkPGAdkXGlAX/Ax9OEiQYDv905iua1b8cAJu7PD39JX00W/YP189
CxrWyFNefwoc+rk+siGiD7Jjf0ooGeZDZmjyjg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HK3O5vzCNER9g8js4SKz6W+Zie9dlDlDlxGQF2WrvDyya1unL5bBpCJy1w0Xm1cUo/y5lNUI/ADI
uYqE7JGFvbSauhLZj4HImoydapRAa/ZLL9nSRfszIVrPI8v6qGNzlAIC3uzmQS48iAygYUrq9YT1
qPItKzIRjW+YafjsvhM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
haBqrpdC8sHCosML+5AEE8iaTVrDueP49m0Xd+C16lJUg1YPcQ6EHNHA456bk66+nGBPSp3B+PjS
04UE5wn9q/J8cGL4YbVE/GY5wVAtR6WtFplMeOXISx0KcrI3qk/KzRrP9Ji6/ivM1RBF/A3FJtrF
qq4E0RTyXYa205RDSyJAQ9RjkwZRwEtkcJ6VY2sYCysbDHMzh/lD130AUg9VBNSdV8LSRVpcwCzZ
sRog7YjwhxC0jQK02UyUpzfW4/xJ7RqEZDh6icr8dQvRuVfwm4y9IzcnYLipDLpn1iVw+wPGS0v6
ZJj/N7hNXBnHUH6mTiT5qnqc1qaRllFBLOzRgA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8144)
`protect data_block
hqvbFOmMDnBV5FhQhq4Qu6WsWZtHVr53rfFBXkv2QXl+w09ydUWbbYE+MMHEvIttUv/79Bj1Ri3w
s1zZxp+OLZ4yHuRZLXW1nmhTUwdR+tKzvmLggcBvvJgBx7dBTdbjRO0REHMEAuzZxilaxe720eC5
kd1f5Fs7eWgNyfjFjmoYnRo974xrCrnigMrhKpC5rzuOjH3w/a2YnqOJdkqgm3+nSFhFheyh/7IJ
UpywldyDbk6mzODAycy0yraZk9XCUQugEEOqvOGoBztwAaQu8DnFbvNTyNxg52a1mmWsiXn1wWgC
GCbJWkfGQTjg86hynMuNJO1QiENKPw77pY16xpp6NyOjgf/1Z+L+vs7fBrzeW5tFSgUreU5JB2A3
PUwopUIQWcun9D4sF3ZtzIYyj1686gUCGFney+98aCvATayN7oYRtq8eWvCRvLXE+aCtb4oSMSGv
3MxAAf3q2MkrCBVeqZcnlEFb+VVXwnR1A8k58ELdc2erZByM+QhgTJxptoR3DUao0hut2Cj9phy7
We24RLJ9VozYoZU3R768gg5apJA63AZVld+lhbJgc0yF+4yFEszsYT6UGsdNpIkwKjiw+SzqJUXr
Iov9APmze+wddoV2iI2dw7LXWl/4uH8anbT7H7dZKwlAYpmgaBKlD/7RMB/Wd/cGShr0N0PVg2La
qhj8ZcM1YgJeOIdfzmJ0jTJAInoBAzNsOqZnI7kwj2pBhFNDm/+Dy5JUZIVxxwsrSTBr2UTJSt47
0QFhOK7Y6qa7mBD4bbzryOM0kZEJPAC335UAulJ+B2IfwPQBrnVvX/REvY0pE5n+EDq7oM7IZUo6
ez35FSL96FCQqowaleK68KPtE2+vG0Pc05l0RgeIW7WMQsnpFDlI/5TISlvTC8JOKAZc6FYIpfvg
0E13wLMB9n3ZeiWgW2ekDTq8QrtdGfNdGM10kmp5kRdw6Ot0ab8Yrcgqb/rR9/SHLKrI56ij5NMO
3Or9yLg1otTbHCOdQ8KVYjML79Qc5glsUDe1eu02C1TE+DX9zJWuhsNI+6WETabSreolujG1sDPE
/UNXH0jcMPkjxxeOG7qvzjkM0iG2lyUptYytrxZGcPmN6T5oy5CC1LO0K6q9eYcDoqDAADp1LWDJ
vpEUUMXP+vhZUvNn+WaK67Dugqy0PknJPaXY38TdXZSWSVSmXYzMNNTfUkrab1BYGCBOY9Qd8+CU
oX+xkdL288UgpQpNMfC/sYiHk+z6pEkUjAVx3i4mg2nryZDp6uevGkWp/TpqliF5Epq7kCm6BYTX
JLKezQ+wUhC7F3UMHsQXlfAnrw83ULpZkK5E6DDyJ8vuzoDMN609WDNc4C5jGqpo9o9qOq8pfAWF
rKvVloBWC2MJV/Z/Wmq9g4tJfCTreSMvOLe9ZAwnIDVK2ErHK02yn8386VBa/vjAg0qJJ2Qgyz9V
wsI92Xr6ruWowJz+Z/1ChE64rLz9Daiond8z2m3xBth/u8xfW6cY/G2fdSQbdgAMO1G88Ls/Xx6i
Boj5Pn1IAdVuSMZiEGSDBvVRPSGHXRSVdgWN6LRSVYRR4pBuejKR72BDjocSgtZsz9kgHA1NZULN
LtAiGZQSYfN6kowaGMT830w0C7dbjYWwm5FNmUEn2+ipdVabZYGLgQcyrN7HaLBw2XGAocFRJVMx
099fHQrRAtQXtPsOVPGavZiqcJ0uZgpIhxM1Yq0Xyt5ar7/ENSSCmBSZfXFIznOAmKS0LxS4S109
oxOrhEWDMj/vgEhLorEQUYqkvQdSaA0BMSGKkjdLd2aFYGDILW8+FDmt8bV7wTkXtnWlnx/U8hlZ
VYa4DX2X5SLPatIyNtYh75RBik3xQlZEZXHpVBTOm+uYLAu+m7xWf4KNAS7x/fFoiHs6Klo1D8Gx
TuNEhhBdnlN8wRtqJnthLxDXGv/Pg3r9JfU+Z9NlMZW4E10tWRRjlxN4hTFvnkQvbhWU4twm03bv
3Afe90D+wWNzglJZ5KEV4smzvQblTT8RfvhlW4rynZIK0WjL8qN6+eyY2vuydTKb8jdR8HLBQUQW
SExr1AarxAfunxTHFPf/idERN4Q3OmQRQ0IoteX47/FSbV5Py/hTgPZI6upx0ThXAUGgNLWszvta
7kVVvWL4bTjU7RVDQa2Jf8LUAn2qESSwAmwG1sbBHEOyaZ4dH4j6wUT9p+5E+0dr0zI08YNj9wY+
ucDGpZUnQUSXbOGT4jE+OVuabqNEclj9v8gdkAuBLeWiZ77m98STzA6zhrX4LVanmMfVI2EOgkEF
hbSx3Om4NN01AhHsmhInmuAtPs0Wi3mpHBYiyjP+cMEFlBPegd1tvYvukoocgfidM7E3ZZPXNU0a
qA0NP6qb7m4LksUb04c6StKR54Wq/STDK32gIDeZyfdOl5FkxV2/7drS6KNGwjgpTc8/8o3Wq8WE
mdHaY6U3E8K8nthBN8pyP7RTTJOJx9XM887SyIcYSZm8C+S2L1l1lXLrX2gFkUJ81A6xkDqx3Qx1
uDrU1TJ/iAECvVnMj3HvcvFjMU36nei100bTa7gtQzAwFbZIzNFU3H8zjph8lW902Kfvol6ZXBH1
rO06cVQ1VYMN0mp8XAiEceO2iB/ZWaeK0O0PDUgc5tUTHXbhTCPIy4PV/rGg/e7eauEECXAT/Gfa
WK5sNFg01fj+ExsjV1rj6NRHQB9nrQ3OBU19KjHoAfOZU63NcOUVcOrHe1WJCheRSyvlLRg+KSFO
H1myvA6N/beyDrQ70qZXcIrSWp5MugfN4+FkOe2161vrv47hKFe0cm/p7jRnYyyE2giJJlfuzDXW
VBb/VCo6jKb8kwq4Dn4q+H8jORSBfFnZ1RMgrwSE817lviaulo2ttA6570FchFsqw/r19XszTxAt
wdOwgA3nupG/rDpuxBR6jSbdl4i0eS5wUs9uj2zQCct/L9P8DNMDaGKDtvEOZeRPBz6d1KE8zsIg
WojgQsFfNkkDRtNXt4bPFLH/+Z+qCKS6xDBjofcQdGhyb8eJvMoghFj5UdJb59+Cj5kXC3cReDqG
eI7522182wSjg4jzN4WXv6aSZtgtQUwrHGBU6UH9DEJgcx7YMtkHhDamifgUUMQOeXjeJ2321Z/E
VLGPtCii6GOgbCqm4HF8Fa2A1VaJXtzvg95hJILKPzB7jJeU38wfsrAZwWU1mCz0gzXomeffjpm0
SWRYz3SHoQ4CCXce5OL4yH9Jd5wMUAhO9FPNvJvf4YrVFVD7P+WtX7W3OxhuZ2XMp/Tdx73oeSs3
kDfCeJ6BkRpbPgHADLywC51krxzPeFuXx6HIfXI+DvJSPxrw8DS9yU5PGyHVtHvQ1CY/NHAxJOoB
ZLi0YWlZ2WouaVUSY6IbiSDDTcDlHdKx8yCPqpzz386g/5CZl4wk1yDatRIAgS1TM6CtJld+X9jF
vO7hL1eQ2fCTzvoTqu48OGj5XIEBJ7GoGTJxRp6vcv+8VkEq4PQmTyo+3/gmZrgmwKrfRaMrD9eu
e54qTW7R5danCN1Qf0IWShyr18y/SgDr1yLuqV1ZgU8oeNKuqufT5jHBXQpG8amxH/cn68EZKfkd
hTuKEgwRVi012T6cOevry0lD4aX5307fxfL6TYAjvg3TMI8LzCa+FKMIFzjJDLtPydHoso85MdAR
L9ZPtd1YYCQOYaFENPlQi4Z5PmQ26GrJxYhKGtFYyDO4nXWZfdaDCxiZfgTTOmb5Xrf0X6q3D9nN
Tby7cm3I2q45bBl95jmj+rAV8vUpyiLpkFOXS1B1cIulrYu3SjA/QGD7ynR0eJDEt1ScSoj5eUZ9
B2Vx9PMjbO9NrEbQ/JTmcn5F/f7L3fuaronMSqLZJ8/7D9bCcJcMgt5K1uozsSrSJdT0WDQk+KzJ
IiXuSfjR+PD1oYDgkmLVpbPmXCgXpIYOD6dqzYoStYd2PL4+ql7v3XTShGbQaZ977sbCRChPq1Gb
oxavqZOaWAXHwR1aF4/clEJuf555pn+nFkP7atRgOJtgQGKCZ6WDclBJ5DHrEBLYh7GKU9YHy3fI
jplHfXru8YSh0akri0xYp9+KUwbkkfR97PRYZ5fhsCx1t353fBNQZPYssiId69C3rd10NP/xdTk8
wI9/4Sf8+ytxTpdHUmD9xPHVIc6Pg3imKQvP3aCmXPPkBzYnWe9pdL7pzbroq2MXhoQGAFCfLcD0
U2yMKoAmS3PyLjhzSjSSUIN4WtXZiYWmaQ9DoXuiL6UDBYSI4wyqWKrh/KFO+vmR/k/vhzwLBPl8
XrsgAvzBMY1XCGuGd21XTyZRb1rvFGxbf4HFUssMHRmvXgVL6exQlY69YcKWLs6CbZxUnsexroGf
kvLK8VZ3kI57TL1MZ9bFIVBFryxUZmD6tfXFBNUTp7X7KGwGy6M6DqxCi6Lhn3MlqRcZ0fvaOV6F
txYm9lz0tTWPxkaWOpKsRduyDHoTNcIAVE9NgRoy0HoSOwsNwpSLSmtdnCPbKX7DM/lv1mRTe5Z8
oboyFrH27M/xCR+MNFg1LR4VqN0rYyiRpWTpz0okxKlQ7GcmveyLLW2HFrjjPsNNcLC1kgr1a3Gl
tpnzT+eBBY0KKbIuF2Qm/WCV4y6My/VmHEYR99a9dIHY7cDW/K3ufNKNcc1MCtQ0YgexTRTpQHpp
aIKjj9LcMUqKM6UdNYCtzXp8ix49UgRRWqYIPeBpJhqKotgwvZruy66WnxIFfmAw1O7diHZm8l6q
Dmj8AEzfqM0WxVWZ6KBh1+iewzhChAbTSC2/GxGXBWbfJouF1ocIX37vRyfriFfhFFoFTVFMW34N
WtTkJdTwMpBv6NXjJ0OeyEF6I+JKNtG8umBXikH3nvjaeYmkCUSwA/hRA2LzSsBnRX+atOBRQm4A
8s8/mdD5Ve9qwlslt3KuvNODe5nJItDtl7bLVExCdc2GP+S/vBkqw+ZeCF/LMsIkZYv02E3zxwnq
o3/jPwJM5g+N+DtrY7G5cMZBK75cUnSMP3u3VIbR2JhuAY3JfOatxpgL4wX58FH5w1Cjttvv1rut
B9A4uA5XrxmIBkmQV1OtPpr2hsPsI6bYRve2Dy0BTZfSOasGVzqnMCu+vhzPUBg3tVIvJlx1DX/9
Kpv3F6YiTSgFmuAL5pZpt7EoFg/W/7pBElk/hEWnpKeqKHbS9PYUqhzNt5cANxSeDSk7IsJcb48N
2u+MvuXxAgj71128/UKM3grhsSZUTxedUdsrs7NxVk83zjZ7tH+9yugZ6I3n9dBBGRGb2yBBq37t
lNATqTFLlTa7xiZh9vQP4lYmJiKpwJ+s7vMcQe2AyM/byZ/r/Ssd/LyOqWCYFpc26kzkK38ocEeH
A5UPAxSmxPjt7Eb129/EnIaWbSH+rveDiNIyxQpKPElbBs9yIYFALPye/rmDXDA2Cs/JnRGTMzvo
SkcVEiDxBemjdwufZeDfXiwI0woPNM1SI3p5vpk8vIUhJLgw8E/IEY1Onc8T/GA8inojtQ7fsolN
dDXTWG/HUkoQNbzDr7STF2jW/p5B9ukDRiOUzVcbIXAaO+grXG6SbGgTVhXw6iTyiR3mn4cz67Uv
CYpAiQcw1VWgwVETVA+v0dOx2zawBOWtJo+3WCALWVBc/5UcbqK7vSmU2g2db05XkT2t4XmF9hbF
xPjfPaw116p/Ry1Kfx5TDXSekpq/FVnhD+g3n5spnHj/oi7ps8WalBl7KzxNOSwkAsNUcIB6Bf4D
jRDKu1kyrAIaXsn4xmLPl0C7NjbkHY4NwXNIsaGYJWKTHQ7ktnQcp0EvGRgphnD1Zk4sZyP4Pqtx
7RHOmzAubaFlwX6pX/LoHTZ8gHf84pNKxA9sebKJOHtHDtVHJh/fx+h1fdW77ZUXJOUN5hOXhimx
5WbqEo3n9l4AgPfMOMXLPQjTtTfCG5MqHnYH1Fa5GnnH7Kdy6i/usF8dMlnL0AT+h/tu+QVogm0F
yCBIiLGSU8Im1F+9ZLaAW41qhykQVEp/IF7IryJA/0Ih1c0Y02rU9+zPzawQ3z21n9hkcs23wQ2T
kiftdFn/3Y7epUdX+QeWCuM+7bcV//CPQZgI48Vq1bTiXR9d1lUhd84XVRpMC/O27CbOU8cNZfdh
6Sejorh7hkGr++iIqmo9NiS/F92ZxW5TAhvS8RtMecub0alpR4jfCmYCguRHCQmz/36iKJP65Nm0
YjVmy7s91gE62k+7YGgdp7eR/AUPHQUFTziIFMgo/5tGmDqausP+Ad7Pz76hWXUex0wq1z5gDW4G
suqKep9GheqfcrR5rQfG7P/0uscq7NHIKuGcVSxKszI9NY0AMjp7/UA4mXdelx/uSSJg0b5rhO02
kSWwJPiziNfRld9tocY11SeLIrSgHJDE9v6v8AUrV1B9mOvttL1DEsf6DliY25nUW9riFIxqmtPy
rPHpGvQAgrz5MELB1yt9G96AEHfGLexblUSLs02G4aCPvz0u0UV7K+W6yFVvBDzQGIw6ohqeHEqc
aveBkP2ZeQOdVue2kffv4WQ/1TZy5N5apdMQ8JeUseX48210g3cE/cQUhqEMzbKf7RoCe6XoLN2H
uWnQOICB5avDuBPfRHxBNeyuwLKT5jZYQSnLHi9celDCkq8v9HNWp5oZyR39wepMbXRNUYvcx2k9
52Rlv+AisSvqWRjQyfXXtEXHFbcwK61mTGJ1aggx5EhVCbt2FvKqoOYg0ZzA+G7V52R27sffTFyJ
YkKwFSmAC8Ef9PhrVJeKry751V/sIKEouyFq/WeAsh9VKtqlKyN1FfEiAFl2wsZx4We+8seqAt6E
VgzJU1Qp2rpu/WVFCDtCCkbiPtSNhFpFjgnSzgPbx2nca8rhep4dIxdaut0ChpXzk2kQxUp7uQnF
HtrBqLPrnZB880S4P5zopiHf9WlzgFKre/GeG/5WGbYyYMnLU9DEoouWoED1NZKfQJFFi3yN8dgX
TxSykhiMXY65iBU0Pbqwe+DudVZoG7580RllElKM+bB18SRrpG2rOfALQlAcAsx7b5JrKE2Mvulq
eYRQnH2l70mcrHIdPNeBqbwZuJcUgIJaiVxrnlHWdJSG8x89VgRgm7WQ70iMgONSIrfEh9Ubk3Mh
55nSr9Sl6/gXO6vVKPk8xI/vWoxmmZJAf0jY2JwANgGgDHfjQ0Wd/OH4F83RsMPwEp5qOmjxpDae
tNDBpjKRiIPrcVKbganx9UjvoDkPvIZxja8bwNtTbY/Ar63bGbKYJSabn7IOnRGXsZeiMdgHqqg4
yFFHXKPEKq9K6n1MpKItcGlTMV7YIu1iTi1fj+7oAH55/uOfXnK1eHcLKEaypSbk7Nnqd2updCML
muJnuXoGm0t3o05iRgBelYjdtrV7uVdWszWIFMMm/QMAcjBYN5Zt3I8Uotp3s93wjox0KyiEIRH7
PLw+iFA1ec/4QEBdEEPGCeVigu7cuvNBNfWhA1sbXD0KhjFTwuAVzKXVSTQaDlMziHpPl7vRVmBz
9tUd0+KjGQkmIKUBmCSf5XZE5nC6aDUzXQbLADUHpqAOHydgUtvVC2fllTLiLTdt4RliUKiRC0oE
NV518gQT7nahZvNLrwrBs8+O2kNqn1GI8iKT4jRrNnD4VMZi9hefT5XjDcHmLUJ0ONI/Wa9ifiKR
ETDXDOU9nebIXr7p6AOzDP58L10ElLGOKtRvyhWJEKc0pjPyZe1J9e7eFhDj5TG+BjxVJtYSpaJ6
YP8mN3SQIN8yMAB3Ik07nY2uUzI/MdLongF/1w7czVdB5AxpGSlYmEnE1Fik4YdbaDxpobrLmfHD
OozssVo1xYuBDfpA3s+C4Mpue1b2rAPp4E240/xQsdhbNzOBiobvWaXVyb94d0QmMbPlzQzVonnU
lUmzZ65Qy/3Sm/J4lw6UV7Oq/Bx+L23z48Fgd/JCTE/hTvLhL6JvyZOVy+DARNgFpjApFO2BbckF
VCHk5no06bvCkqN5eA5f8y9P/fQfHsUbplnlWyvr6UVfMrOEVoeGwiLkGMUxC9dMcHho++RzhGHM
9AlwPW/RMInYvjnlSilrvJ2QC7oY4y4r1tzFHCjl+m3gtnSPlTmP5EcjvY/YMzRWZe09vyBgfPs+
X/H1cEkMAfhKlrXx/3iiz3cJTIK/L/Bpo2HcjPq8RmffLImhZmquFHmoTG7e4QBOq20mo2mSSD1O
WMYKxMOvXJd/60QmfJGK1kwarQtkulCU29yLg+s/w8rnNsql2FXPltcIpMFYxJH75ELuRl9nu9QH
/698yRoqQBVuSH/qsJF/P2M6guhtQSsoeCaWvUg2Nf/bXS7C84TnNIZR/cie5zGjjZgYaXFUpyU1
rPxhN87Bw4k/za+zBy7xx1bm5NuKrsLd04RWnzf/zFAU58B5x0+B6hl5q4+Y7qYJaM4ivGhAnvJb
6C8PKMk2IsJRSOl/gcHw3Q41QkG5c4g6iDUDK1SiVvHvE83/zvIzFQeVq8oApk3evm51EVhYgoKc
kfc55AloWAjE2iBljD7EsApSl04QK0MRoXNhLBbuR4Bs7UblPrjETHbSmThyxNZ3toqiOaKBuB3N
XTjLiXL9S4wNl7UOhBnsBZ9MNJDnZLOGN5KFnbGgbhtoSCcEE/vhpN7VGkV8yRa3CF/euBIFR3S2
DwCDVYFkCW3dWuTDSUnSNW3048taeDIA0RWebGQP3BYh47cnaJjgbyqNkKApC+ke12e4QULiPS1A
dRxejsWtsxgLArAkpxdLBLnfpkHdOCWQhH26iBf/3MV3jPAOwvfG7GUUQmrNQ3AHR7dxjl96TSRF
EofM7q/Tc7KwUIBEai82HDOAU7fxvrx2N+5Y30Pa86/3sUz3YatcOVypxD8XFDbZN4hQty30KuR3
K/JXkFBPlaTq8LGeFk+zyUydCXPTnhU/rpccSJ25mW7YkgNDks0Hxdoy+aE8r33QUOVXrwDWsgJj
3zOwgpHVnSa73c5qKGSJorCrsLp6hQLf30lsx49/5bzVEL3z0iUnRud8ah3QfkpXBFrFQPJHW9cS
AUit11C5mqE1PKLuLucH5ir0DHMeQiMIoaMuPrhxrIz8DoJ70EOC6myniuPMJBnBsHDqj1MO3vLD
RcREn7wVnaGqHrgDOsMQzTgL0wvAO9huDZtukLqKQ7KgScu2lz/Ys/P80vUxDQjowIQJfY+9rVY4
/lGAGApSnOBdmABBp0dY9rNqGy3sdk1O1DD48hGoEvwY6+PYx//2yKKoXEz3yEPJ2vlSu0ETB1v0
DN3aU3BK9l9GiBUboY4RDGDMUyxPjSdscEuOOxihMyiLVEKHb/J0pnEZ5bMsTeDHsW/jHYxF/+DO
fkeieDYXhkxHpzb+G+4dFudYzFGGnBolF4M1OodJIFPD+wIy6ubKaymAMjESdAlVvRZH/+D2OMFD
sb0zmY5S1jZiPLpxF6rWmJ002A7O0Pklon5UGx+GbactybRggOqTpjQo0tFb8rerg/3DL5Q2HZoR
eAOKA1imoTUCjx4oYoTLzTDThdjG749EEfwt0yXdlvPhJIdom/HbUK2FPa+hKV6JmYLUEaSlCDmv
2ysJ07be/N6Jv8bWxrWAXdMlvmHzUYggBGUpB63iTFEIOc80S4AhGYu93a8PbnSNI0YMzGzh5YLQ
2s3n6z9mNJdzJwEqW6h11i4tulOfDPK8p3wL5kF76Z/i9GyhOMMo98FYWpcmt+YfMUzJGFOX0hhf
ZSTYZk8s3Lz1Cg/6lIoKyBZ/V0kWBbz4QP9Pm0BgD4CILTtpqPDBax4R9c0UvdOkT4L6BmxLpwrx
cYlIlNMvauoEkJk+8w75xSmnF+2AWHdKCQPTmnsnPkSQ6RxQqcwW089qHHCZI4w8aTIQGsEaW1Oc
knn7SEOCOgKUpATMkwoOYaNbDMa9nBMbvpRSuAkkaCcxjjW9ZKHjERRuq89rg6/moYiJXVtLtXc9
FXX2R0lAwyWA1HzAvJiyoYoOEzAgRxGMZc0zvTa0+3SnggmUg2/RdYjB0gL8SvXO+TzEMSaotXbG
2WyiNj3sobvW9O71H1AsmsSczsX8h87YGViFE8AiU3TDTbBhyAqHSIlDIwv/B+FbuUde44wiUNbm
m92L5g7AXvv253i91WUjCKJvchZLqhka8z/IhKkg69Pptm/JcnqdCyrsOx+kfmOSAhELNfWOALKO
YNvyKou/cY2SwS++EWP0/F1VCMxJ0eANxYKjXGi/iOgnSAt2PooM3mYw6EttXDzk+sOlL5W6C7Fw
tfR9HmujlJYV/dzcUyadPDY1j1U96CaA8SMeddO8Su6c+r7SsUPTUPy/NhC/oipdkVpg3MK94Oom
fzpRjrcxxHBxZqh1n4957pcKPONrf/Zu+DNMk0Hvp1/AUdkA2G3eifescE7Lff3zGpEnu+K2fGF+
DvsAJEyTPWOGSaqe/MkRjYS+DW37g/RTbV0EZE7YotZt+66u4r5DPhC0W/0BeQW9/0PQ+b61ZzJB
udkFKWMZ98xmOkI+3xOn3sfOSl7fwkDqSIF0RxiG93nr5unfQEk4wKt6ntFX8pzPHbhafGgYxUQl
yJM9MqOB8Dy6czbHWc3aTSZffxPjlze/bb7iLCHhdbe6QEzvrz2LUQb+MCzsvJO3DGaFVB5zHPEg
g8y1a9tatjxgxWXCY+LfKd52cdZGCfR9ZGHsWnhi3CW5GIshYo6xiPQ958yY4ndqq9cJAkzutipk
ZlEbGOAEkg+Jy7y1qZMWHvBctFAbIc3gK+XgMMGt1PbJiX4duZwFo0kDpS7X4QN8mb8uhCniBqrA
6qJrO49INiSi0WRRSQCtWGtnrLOnX6RHZW0b9ntGcr+ydol92rNs6u9BjXlNns5BdB+as96qvqCp
c8gGLXSR3uKnvl+a4ALXp08rKfy2m8lc/d9UifW480pordEEEPan03MfKn4IttdH+ac=
`protect end_protected

