

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EHhlU67zSXzve/de+KpY85nXXvMNuZL7tYgf9fn2xs2MMX6KZ+NkxxVYV7RC95SlNzgUt4DfQ4/9
3ul1mLnDjQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UlAZFSxNoqgvPPKliBxVt5c0coSpd2sh9B8mE9L64FOLOsIE10QbDZBGLO1c2gEWIwuQ23M7QvQA
5NLCK/AU93Cer6u3Y5Kw85Zu7Q3cTJ6gtsPScNo+F/wtG37D/TBvZy9QIxLBvCRLOZx77GL+Y61M
X3HQ3kaL5tpBN9LRA7Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BhywTGDm5IJZmP+63CSoL/TDCpGJVG3VkCIbV3f5gGTJ6iLDPwvtFhhY8681GBR+EoOyUSMbP3AZ
DMFHBgscpLa8vafzBYp5kDkIAp6zpVke5p8WT0T374mfT86d/rJV4lUvVArJtTXZ7Qb2BRu+oMwW
4NXsxCdhgqbldJw6uUCqk28aEPgcbivrgwKY8foWfBnTw+EKHyn/oWDvwghTokcxfEnmhIMsR0T3
yD/98FKNKviERlHfn1BhQ/aqkW51Vp/q5U9qrKs/+lZwoRMsy8lRZRggDQnNmQrFO+0t1Oq/DlpL
Pzgpskdyam5KjVkaaUDiD9LunE1mnunv1fkvkQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M0G+I4o5qs/wY3cBNkJHuC5SdvD7yJrXn6vr03zDaDrjCzuSM2xSWnhAroxnc+rs8YiB5XG+kxRS
nfrpZghhDmt8SYAMsT5eb/ToWHwFcmxPkOwf0TCRf7UHox/rcVr0f6gppZYuBp8i/HMdTy7/9hVi
Jazk/jJ0qiENaXH3lhU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
II8O6ksX/NQP2v4t19inJMyzBruYXofFp7EnZduWuRh3lmwU4/uZj2tsoMzEFI9GURJGr6OGMrIR
LHPoTtEBaHFBnPNcL2m+mOF2hh90g7CmgF4J8nr08oNvCPZORB5fd/Cj4ujbrC4saBHdapCX/nOt
W3mratI2AGAl+T3t7Q0k1PLokEpC1hOrn+eLqLqV9hKaNBlW7DfM0Swj9M60AbHp0kL8sQjj6PfO
zKNcq6Xvq1JnJLzZ115Py+hhtw8g3az1/vAI3s/sf20/ggZ0t1s4m7+wPif6Tf6IZJCySXPmKW47
LjAxEb+MGgXZe5eFDZ4nbVPt5Q03mtQWzOAzTQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6240)
`protect data_block
/ykFRCRstL5zbQZBqKdO116XWRzUyfTltZbG0SNesags5PTVSIoubrmzUYlFzceeX8QoxTjQH1Jh
f7JUp9toF30PqSOJ4ReGZAMShBgKvTifsGyolmeEQilZhW6A0F/340lt40esJ7ANV67u7IFjGdTg
h2rYNjuAbTsn3Rf4KV9v8bCWlVC71UJG9Y12K5PmLKl8+Gc5KlJ3/TqHYKgv5LOS+pcLJc2TwXYj
ZLEixWM3BBS6OSFKqRsWz/uPBtoUA2mGF/z65aFuNnY/riVJRFnvXQGNOudUk9+dHcRbuoBaCxJc
2jf2aEhuoWiDEi3/2NPcE2C3BXEVQjbCo6vjH1Gcnf2aiNROIVYMaiofRpCvvBBKR4ZDNXeiDsvc
xdPaWkBh6Rno5/SoDkmORuGUfsy322jZzQmSLwB+KOrt1SmBp+hplFugLJufc1ISmScVCUDHtjDi
3JjWHuIgrDgKwCJ/ljlTD8upTE5YF8fju2poVUba1jMa5bC2b10tfCJw4K5HHW0pIijC0Sp6HjXy
t8VEerW9V3DyWC2cLFq+xZCxHNrX2rIId6JA2x9BWMCo2nHwBX8wPhz9IjrlAJFdw+FlWqRDBXaD
Oak7HWX9HbZNGMWbQDkKYLKnSfSfxfm7TRptC7//Rg0EB9qGIqXe5xGawo1sT0nxpcsTOPa7ipUG
+No/zFoBPe0l4a+NElx8j2Bf3geRIk/OupGHK3As01YXozOTbvaX9ORwtvRXdmmO0vywmwDKtf6B
k/fLb6GKmhbmMNhamSp/Gltcg17WiibFY8kG0We7Sa/hBtk0cxCkLTpODqgnJ+/bZSm/2vuR0L3J
O+27kMkTNwOZgYa7gSCPSm7OWa9tSJz9zAl1y3y0SmZocPLGDHc8I0p/WF4o92ff0CXb/xKD06E1
ajJrLH1COywoTrj4cgTZuXAxjR8bTNtPonCKV2w/RIJUnl0aBjXzBKBUQbj3OeCTOeeeFLgU5mXn
kPlM4EqadLiHvrJGS4a+O3xffiDR2dLpLhENVl/K8wlCTMFvJqH7mvbVTt88d7Zyucpv2m9seQ1g
BfWkNSslOpmdGAujClffqIiXsYh2YcOTu/uPiOpluplwQOSYDbxK9l4RSZtAGx1YmkZCj7Rh1Ovp
YkTn+5ggsXk109PBzu0EMUyTqUNhbQyHU6CeHGQY1eum3qSPbw1gfUH4vkcXTJZ/m2WsGWKKv1oQ
srBm531DEY8naVvcfovBwyTuo4YLpEKpwqtuSkCGjDimecY2mQUewnsHFiQwnREQ3mTknIfVx1p8
CNufeXaH8Bculs5aKWaOTT0wXJ+8TTsOkp+pc2uKym4UIv37EaqZryI/V5Kg4RexMcCF/LCU+tNN
3++BsMgBxDUoN6Gw/oHwChdEaw6QUokFsmZ8Sd5fUeZ9nLIcji3rhnBJp6XMjK07Q85zusKG41Kf
0ueUVAgM0Y7NiR5lVnogjykO4nmmLn3OYiFL5ME2B+omWfTjuZeZCj/E9U+XmWA/5tpHVTP9s2Np
kX6Az1es5t4suvGN5k2F/+B/QyI+ez0RgcCBB1NqjSpgaVDFJJ8qKFjgl2iYSnpsqZhVKIzb89R9
hDh1BjQ616aJG9ORR9RkbqF7sdVR/qT/0G/GseQWNi40x+ZLURTW+/R0v/DqHTmQUg1UdSq3ruz8
RlANvpaltb7RtoXpK3Hc/TOeWFoHm8MNIN1QKiflZ7Wu1W+VDrMsqNAcs1es6Noi+18Gzk3rx39D
RcvyCWgnXcx+3JAm5pTiICDGBzLmx6zJp9V1fmgPClEB1ogqeVJcS8asq0halydeVxXkBAu02keQ
zd3mu8khmCQ6ev9UbMoHFSmld9pHnxSOzCwexuQFFMAwS24c81pnaIl9yf6tiZmTv3Iyw9xqxaTY
yHadFcj/pWuHRLpBcSZTE/Hp8t6jGQ3+5yC7m0Z/LmC0HJpo6LlFuTnHsPKv5bInXTo3kQREhLYl
JfhLjhXMeTo6p65tuJkUEGFvhzQK2FTnDN9TBDhnAzJK2hUJA66Ri7nJ3bbub8lO45WwkQJnujL2
NUP3EI87Pco7kpZBMD8P7s3vkxnyaNJqe+hkG110MVfeGn8DZW7/KEO7P11gjRvQxAHj14JTUaxW
X41yDfdizrnvEEOHAB9Xn5w4N/1oMTsY6tnx7egce3F5wQoyM+psR9Amb0rPCWlyc6b+39Z3SGXh
MlXXMCVY1VkrCIm3rSOk7Yb8J0vliSbVkEy1f4D++IXSpaDdXIcrZW8N94fD6KxHoMC3OpN+oyZ1
861iwNzEw7ahtGcPaUXnUNn86a907cOKlZmozyAYmU+7JoLLrAxVDi1PJ24NSp+jTlrECi65qh+A
NE7RUpe6hLIiJOvkLNhxKGD09zXVk0k3ASLxdpgwDFbnvx6Q7hdWc88SpNJ7lWjF+dR/ue2uThuk
ZJ1qd9ePgmXNHFBstsJmy9+reNBC8pkv+L647NVXkVxd1K3HjoYdWyf3y/qrc1/5G1BmCqfSXPNY
yMEZHxQ0TrQt9XwuxX1gNRsAiiheb7Ig5gh8RzYvAOaDWGd15xgszb0boBCJ6cPAHzfw4DLnsECT
BF2V4XeZadv9CWNyiQ9gIAUp0RfhRG8yzzi5d2rm5MLStcMzerDmHy6mGHUBRA5GexsopeiKgMNh
kWYs518hg1nS0xoWrqpZDzwk/oWaXTSd5FpkN4Pst13AND2BsvNjJ1xrAEGlb+6qx0/1eaIukpeD
TYNB4jW/zCsEQrFQKOh+N0koS8SkYsSazwA9KT1UKabs8h5WzK93AGpvQxNamKXrtStyeG1jxAjK
lOAEkb9KIKjSPVh29Z6yYYAvEtTO00JmJE+RhGymIIyJSKNfxVgzgSCmHWUD1an9XUGKVM45hi5N
gtLVWtBITO5kpMYBuRRpl1ee3uwJzvC+7k8pz4ltHqOpwCSM6AaHQ9n1T9XeQgCO5iHE3rltLawX
/Gqo5JZ1zg9b1UcCsiQmRjJGBvHduyd5NVJpmxQlvr1UwuNXKbqbyQyZhTeHUak0CzcHWJ3BJH+x
v1ENKD7szuDWdadGdZOJss2iz80f5hRYab9agBsAE7ZBMEoDGEH560ncUkMwgX2Jlbkx6yfHp1NA
S0qjf9Pl5HsERDaQhEnIpS1lKUieHsLURxTjlZaCnjz/SJXlzD98S/7Ou+mpsr3V4+xCMBX4Au6K
9+WjkG9/L8S1rRXgbWDtvwfCJ+18x4ZXKO35WGisQDF1Z11tUlTAcebKGmM4YFNmYxYTMk9U3fao
3XG9f7y3tpBvd4CcZCghSK3WFBqH8ecc+r/bZZpeR3ypJexjsiMLN931afrQl+py9lGUMv70NtKb
2rsFLOJFfMV/kBKIbS6m7gIafCT1yG+SN38h+SWPMan8K7FPbcQK+kMxRHeb/t1cn/SCV6xEcbIx
rGkQh/v4hlTqWuS9ou+0bTldh7LaSrVQG+0//u3ns3DaV6LBSoNM1a0Nq8fSsZWQiIKwzTuyF0tj
woXp/6H5pUDWVBRxXrlI1CY5S9iLvwl7bcYVip486THZA+Zp8xRnXFjH855T5k9j7z8vxrvY/0uQ
lF5NDqfaIcYY2429urhsSMB8RQvW3KMxjwJDjBNwXo27ghe5Q7hzNcbzcOpFfGrGe5ubKhfk47nj
dy5475srfkxHeTt3XlJz+omxY53Rs2ZeHHP4+08wI7eRVpyydoPePCOhjEOxYZM8YIasJ90DkTFi
5G4g8E9tr7V2Vv50PMg7M/Umo0aYChWLu+NFXD5A7vr4EHHj8MPs4yLaZoXIDJtkmzIXRT+vIuci
diHxyCE6MuwoSj+EaXpkqDL+DAvyT1FtCsQPY1a6otzAjkvhx9CNQ9e3Rf/EJllUmNqMLtGDj33O
qx9s2WqUwep57IeiU8z1+//XBms/aYUz1HrRSvZFnv0nh9QFuzKyIDBupHrVHeh1b5jgcf8h5JwQ
XAbB4NxVPMdsYdCnuopdkyKvq2zll1f9uWgzjAhEo98aKgiYloaRc9VJ/7FWe8S0RzDbywZE5c9M
mpqiP7D6TsBov76vf4UJYHe6iEORkvVXo0KW13dJy+Y8mzPGdBK1CVQWCvrGW7H+BEqwZrlz/2xc
UQBsqRbJdNSQzLcC0YXKDsk1McNd7WuJXpn0dFbmEW8gzE8dKvi3hw+t9zMKbVgjZhoYmQKq58Vv
dP0XD8THhp9B7yOn3uH9HhYt1W6xoQaKhGlMhTAEPJASG+EHmLOGp7WdXdNdJJuKriOi3KXxiaYV
n+l1FPJ3WcsKtGuxo6u8t269EIVqEJisTf1raMiaMGhjRTu8J6tpfc4HWIJqQ7R5iw4hT2cdzFlj
+vR1tBJzu2VsvYiAsK3Mnr0FCqtM/FwTBEvPIQkC43G/9gtOSkjDo8sUc0hPfM7KcIES7xZlAMjV
n34i4bp+6vbrfiHhb4eEKYuLyNIHx8yaWkKFUaguexCubkuKCyCARiqfxCOlsV3zV0yR8E54apSm
cGSs71AgWWrd5VpNYmP4b3+JYOXbRqXUTMNuXE4//4AmoHKGW+zqqPqF+XO6QwSofyJqZKqZlZch
1xcFHcBG9/YCnQGADQWsVQXUuwWtAv/Doxq0cqOag73yIA80d7jdRq8QYYn7pDDXe2DtBllU/PAd
eXADFt7i+iQWKoe5wQW3Dx5aRJUKIoOZGGUUwTPt8RRF6/9lXQk9ETQNMa3n2fL6GpzVnrn2Ftfh
f0EOR/IMDtFiT/yCrD7YmpwQXOKM5kt9rbJ1IZ7uQxXy+74vLhH2Y3dsCgLqMYCOwTBwgMPNwMB1
k/SeVXD5ZvCHubMVqiMNgcC2Kd2b/K+zv6wgdZUXqSgvH1jI5L//VMgVJ6jcukVH3V4j21eDeLSE
UmKLxDJqgA78GVjxObL9/AYhP3T7fvK6i91Y9C/oEGY9BEqfldMuF4dWotThS3Xt/43rttZ6HqUd
ZEyPbbhjOc2mZPKTCSXpV+hs5MqjTUcvYuSfA7SPHp2Cd6+lz2A4J8O5IEJkvTjaGlfEXAWWJkl3
02DR27c8cWWtW2eiA0KdxrzYA2T/eKBACaNgfqXefbvOY2zdpGbC9wRveT4ljhH2G4h/XKqgvTI0
sqiI1osl9ucWgXH8+Q7yypTG2x9G3Vc6v91ikj+dYj5kk8W6J5N8uQ21jg4Hvp0s56jEeKJ/PHOL
PopxrwVxLkLgOaik8r+rMJZNKxY1s2s+3jvU+aA9nab+wA/sPnLqA0hicrZx+XMHFVANB8aKTds1
QCEBTDIEdPjGL/JtErq5SBuFuurRXR355gdv1cUHp1HXKhF4DF3mqhJn/lA4xbvZ2+RgIkWQLP4S
xKTUS1mpf7rQelRFY0muAKPjQGXqJfUScukGFPh/2Tg+3GfK5TYvbGIG1dVnRWUfYzk/KPcvhMJP
/s3TCiMmC25s87WXTY7zLyakCcxqOVOUXz5ZxtVpyfsV56ROpCtQBeK2l1zIR2NxxLUzkqS6WNXf
2blxwLcX58/51oL2K1eJjJIsbIWAvsk+yPbCg2cqUrmqD5I88UevVa262TAuHFZXvsjVrpJTdVal
OIhls5tiUHTpWJRUR7GOQSZcGfdQziLygNsXjL5lT38LPWDSD0+xSVdQ3rTgmyapTiExRoGrK14H
Fft9GPOs5+edmTOmGWIlt1JeRutwDPhYHddkFM5izxrMo0o++LZ340vo3lx3jtqQP2O4O3oSykLb
1xgJ3lfVjgt3GbUUx4mzqf+VK3qtiRI3CzHUYUl7gI2UJc7PfbkiB1F5N/7Nz9NmTfLbJxwo9SF/
3peaG7vsZ/NRM3KhN32bRm+68OkVyR3pf3un5buGjq7YcdI7RL9CscfTd2EF30IuWb6eyJNFLbWn
q5nQoEkUBE3MO/mdjzt4jWxA6IxK81U8qOiw/e6FUwIsGtG1aQjRYl3lDSPfwod65eOZexth0Qt3
NqJgDnzPJ6zvket1mjdyrZpj+QDK/xyNM08reuhgJjUi6nTkj8BZd/2/MIuBZsFcIDPPIOkNlqls
ojwYQxA4iHRWcn/4r2QB1i3aZ3JtVARrPW4Ck+b6DadXT3B3sOCnWN6efzsq2OPxyLv2orBUvrqQ
/UzFnDWMVxH8QMWKHWV7eJeQ7tzVGeGevOQfbNMVfAMFLLRJZSy261ec6Ov6lvKorliWCSACczAF
HvXjA/NdKfo4TV26WUkx0iZRWUCka40eTxsKHu2iH7aiYfhKno49W7IVbyk1YQKws9d4PhRhVBI/
BU5K966Cumyq9sijdrqUqEOoSGD9H6G6Z/Uni955l7fdZ3E5HcyFN2SE3HxE3+K/a6wAh3GXsB+3
Kf0k8Xs0lHycjrQMnrZUg2PmgeObgcpwWICmsbId6ohmylqNDwpVs4dm3wMZDjMDX5zmXKl2ODAq
q3Vzzyx7OTx3grLCyd1l/cIfkygPYRYoo8IdnnZjYrGdfENCvK6yDiVQnXBj9i5INWNveFM0Fqi/
90DdXCDLhLzR1utM3fhtl/bwWhpJ7FjrEOr55F//Ab2pbJR94II6shQlLVF/gPiLyV92LIGMRtav
vl+IPgEfvMS8lZz6l3JUOdQBRPHymKRDL4PlUxBW1C0JdBA7BpPJYZiLMjZtr0DoiaYy4xWKpVqJ
X5gpI673JPNH1AZQaNAuOI+9caMxsuke8sr4ufUqeBwaflCOXMmIZbNNs4wB3yzigv66wWjwyyfz
ukmeH+FeWAIGI2lVVLjQCWKOO3faDvbyevI5fm4h36qu3Idk97SFYCkuF9DdHBNJM33MsbitEYl8
qTdv1+gCiW6HRY0SmuaOU49vRDnGVYpgKW9/HZSDF9pVJp086zkwMDzicbQXjpNb+71xTQ5Gj3zD
/wzyai3coyp1Mql2RrOwFeXkOq1qRvRhxrPqJRgoh7C8rh8ytMhLPjXNVi2EV5pAYdTXmazFsMXQ
A3LMlLnkcuvr0xyc0t5Sqkt69YhWBTeWmVY5ASweoYnALPf/RbLwVb4eHrvUqKrCtrU5i+AIvlat
mVdCqzd2A+iNH5jh4C8mPW6RfXF21h/NNApGVFsXOfuHuUDVTR0aGamxNclLzs/NIjlbJZrYxX5K
/RRUXikKnu89tPeodkWGHtwe2MxoozTXgrd/G371lYml6Bhh0+m/1T/kWVF5EH3kfx3K7Otxo3wG
FYLAY5DuyPSD+imGLuPhvXrso5fnaZtGFBWEV+XkCSAqe40L35x3szof7hdKfbJcKx6wwSNaDKsl
KXFzecL/ERempPBNlnUL4OZy7HbjoDPlNHu/tIbvgYJLiqiRoC2cbcPAu1lTC2DoDtCN0ptLBFVX
mpqhhL2+6NGfKpUayBOBl1pri2LPwyEk9o4B5/4nvM8NDx/u1totMlRoSBFBOd5H7cCP3HcFpEcu
QciiZLn4XZeIS5RXv56c237KhKE+XgTTQkRkWS3TgeN+jwRt7O/hZ4pEIzE5PX4bc9FVIFSVFsuC
GD00GxJL3Y1vj+q6gwleSWVF6PKXeYtoer3UCa1Jhntjq0Fvs9qni2f9cC64zqB+mtSJAWwCrF1x
Dt2KMxpvCXpaTTp2ODo/roCTOUGt1M0N+FkxMfuwQydZED/wyAlr39QL7+gyHnveQq0JbLONQbHr
l+9l130suMZywqmnqEOwc+k7fD36O12zT5fasHgY8UJgPBsVorZlo0QyDCbq4XCEM7Ozomsed8Ph
04z/RngKhHPKfOzj1sxxO03GPjaTNvGjNJ+M4sLU3k0wlCVvxVMM165c87hyS7CNB3wV53jOAlcy
syJQit1VuUxnNTmBCIkF5SIopzXuVlusST7GD6iWgr/px1niBJ7keVQlvre4SOH5D78qZsmWk/Of
PnV6XgWUZGZtZCNPouqAd/9tSFmaGe7aiv7YUu2V5iyIkhyNUwBtTc8IuliP4GCa6APEX1XRy7NT
kA6vi/+sStxkBCIW/pJP2Kw+v8V0ydXp4YQH1pgvAvuJdr4i5WzCF+iZ1hKQwJSrs3vwHjNx4lmj
nC/r8VLiFMxOT4vAN2WAyQxCBWdiUOxPkzAhu6PveoqRnIsFQfBq9NTJdLJ0uOQyipOERyixa3At
WqD9fWEdNf5YwhDk3a1gNTCDYklznGU5VYNyWXoARSARjUcrWmzNWAGG3VbG+PB/51jvN6438U/e
0BKp7ufdQPiniD03vldH9KrfOtWg1uFhnBdX5yZ+DtsswYCQWdjb8TEQEWutdl6qzVXO6cvZiT6H
1VnDVNHWmv8iialVBLFGCbtYXCQTYcTZ/5WRP1pD2KD47dJQl1EO3qNIj5IQxfQKE2zW7m9CZBX+
37wr1nlz0guvkXkmZdO38+uDUCdowqamoFtY
`protect end_protected

