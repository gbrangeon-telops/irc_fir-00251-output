

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mwxNacl66MFUVIMc1Encct2aHZOcb2pREujQa4vWHOpoY4Ryx1q0qOlrkehqJnJB6VdIGpRZ75ar
fafQO/Fcyg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WTY81lfpic8wiNg2xUTFY/9pIQI3CKsiY3j1Z19a6adif1iCy2STS25TLTe/dZhZiWj1W1FKdbVN
mTJAkstRD1IiixRw4XPUhHS0kg8DebELiBmCxBLwbMicqplV5b6X9QbZ+d65v5AnURtcySKvK9fO
g9n8up28DiiTZN5JTCs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wSJmxWNG9Vaz0hV3ma6xxbW6Q/tt4VebLF5ALUnEWrb0oMwD9MOvKTVg9bgiL2D83XqOs88TpeXX
Ifg7m/wa0qnVENMQDpzrbdsY0X541kchr6nHO22IjxAZU0y34IzPOD4wlt/LkBIeRhuE2oOUmiUB
mj42HGuDYM+OLJ75MJFObfMegkawW+dQ5MXJZAvaZb3Gdq+Nc//x1D0rUYdDzCYkIE6Z7scW8Wik
/MJTbyzmOPOK9ZoDJMjaYzyR5QyLAdSzLEdKbGH7TxDHRl54Q3XCa50pfJuN0PstSuaixGzvKQtH
Tl8qJKpy3o7KeFGSzvILj3NDt+zm7na/fYnOyg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TWs0qYIcIilONYk/cz99Kwd1RIRPFnNZwYyu+ici+iMJ2JCkq8jieFKJjspKJpdZ8Nc8B4CnG4qj
aN9KKPyGY83yGWxxRkXLLk1fDABMFcSV/QWTMe6VkTZV7rSzb+eWC79VK61VEPbjbvhhwl9UlHat
EKGcZET/5AsZpsdS5rY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J9Mi5TzDBer7RNgnQmNNaMr/oObsCpVjypskaWXDXbsUL9Tz8WTWA1k8rjWfCv9Dmq2LFoNWohyz
5PixLjvzdMk+0EAtGJRSdyjvZnuW2bmu6ekaURxk6HvWMfHmukxtVO9c/su/PcWlhTBaWmQfDEOk
MXt2eXdYnsY9DHX2xUQnYdQty3UwLIiL21L3I3SO1yyv2PefA4p4KfovFGDUvBPco1deVqNYRLx4
GphEA4vKS+OANoIaExoVeJSpvDGH50O+wbHahIOE11SE2zucQ8cWichU4yUJXYALRvrOZArC8ClG
ouWj0ts+fBWmUc+Q65XK9XqQ174/nPdN3w6Fsg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38784)
`protect data_block
upWqknRD1BE7eim1QxpZiPJBIeOGmyaaK4vDBswut1/waFkhLXP0vtsvR6PQYXDhVCpVqyBsQ1Pk
8V+va+kVFJO2WgeXf/MyFQq7x6nuH9P1igIT6Yqn/YX6OzI3Z35doFqshefsGT2XZ8qNMw2PZJMp
+hjUXbAgjNywxO6SnUWkfq+jYsrUyWbXyLR9g4cvU+yXJWcq6JaQrr3oaumzT7iKzp2MwXQlAhsU
RnQhd5o/f508I5nikysdi7hdYlOAxgriPg+Hvx8EjPNUhuRZeMMs8auf7gyth3Unf/R4dvpEBpyS
2baSfqHZW8PJqMhuRenScSVG2N3gKHhCSARzeo0tYIImRVoP1+7Vy8ExsJHPYy9oAXDOec4AO7x/
1bn42p66lrlNIz31dTalx5seQSc/Ne6PnAA+QsD0hnEvfuU0cCcpiJw6rIZrciZdAbr9AagMnc6j
TAbq17TDCjvyAY9vS8RRLU7HaOXN2kHoRWgKuulUGQrLPrZ0OtAOB66jhdpFkdIkFGAS3qSDMbI8
XcRYUDVxf8E8E/svfsrTemm8pXf5kZlaiq0M+59BFCr0z4lppsIVjcENxaiXcrfifuD+1uxBj390
URVBzCtNC06XiO6BmcgJXh6JyZmazKj97AcbEDCMEyJAJyCCQeLO1nlLHQQXazOmAcw2PCAlOMvR
m5O0fsbdMHlf3kGR7MZr6I/SzWYNlFipMivgGamdHF0DfuQKtRARNKTGT2mykTE0QrEuMHsNskZS
ajV4tkNR5unorJ37w0e1CwdzxGRaaVzSY1ae0FvyL1y8v16nPuwCQ4cfBF4eAy4PU2BgR5uEpI50
ChJzm3sb6iJ8NdJo3wz3tye5tbZ/kYzqIzVrHn0KEBOdpeO13Zhas5cb7iD9LYTHvdVKIDwd5Dqt
vayrP/KARPd8jzp8sGaTo2BooSHI4wxfraVUa2xn3ghaRrhdYqdRxV+9Q+KEuskE5ZOglTmxD341
GRnmt4t5eh57CvkQdN95wu4iPAzNx50h/nLlo2Ohk44DN/gvoUF6/oi3kKA1pVQQy928QnT8Y261
vXm2hvlJRAwnbHClQp5vwHS9uuLSrrV12TQFeUpat/MtLrEmEq5SONcuwjbVCqOhwpj4OvpSxWJI
wFdl461cjwqYlWY8rFmUyqUfXV2Yk41IPBvHZYzZTKYsgRKrpEDDjhDqnXnjDeegfRV70ml3Xs9d
sGeS1p0Oz4l2PJTEk9p5eq9Mp6xqOdDFlAXMvLt1AUE5ZDn1OmneJqpnJcW2oiZ/xPofDDrILMDt
x2wkjlMKR364X3qKbOe9vRGrKYrUs084uC6kfiX6BQWKCupYNauUc96PVCHA0dD86o7pXHGbLBwe
G7yywJwRXgviVsyviArEnSBp5KBRwg9ws64TsSHK7q9MopEFLQ6MurUmWXkFF1aoTx1O46/mb7zL
QW6Af5AFP6IuNxgKquER5W/1F/+m8Yx8phvbwKZDfl1UMpUXb3WSwtNvl0xej3FIfciFI62IyYWg
JnHkeSjfr7H8Eb7CJqV3OonUhQbBDBmd+DZN2ZiZNsdEbQEPW4Pm6iltgXNQEWsrrLrp+xXbH0G3
b6HVwnR8nUQ2jbKTyHUssSZxRJczrl+z+TIrihZXYR/uXgocF+lnXkTZQLXLnVx/NycctyOjnre1
0aVsfOoxBosekOzk0+Xnz+RB4iL+tbNiqUFinbq9aSdQ2dp/zIOFX403WSYOGeRVZH9KbAoFMoEU
20b7O0xb6VQjrMjnGEl/dBecK3p1VGqToai5kfya/4pxzhg1gbMgfp/ogsdhyKrYq69jdUynQux2
NDL5/+bk8sZQ7bvxHp3Ljc+sGipeFqRX8g3GLZTvGw5/ycj3ulPekbbggPd205GjlnnzCMUsYxrn
1+68qYqcz5/ikFBw1VXcm+17+fMbiT+oITHytPFdIrsgAZKsa9SN8CL3Aum/NmPp3n7hcNjIEQyn
tF6ACbs6zxSIEG2838WnPWvKP8swh/hz9SzL7Y3Gjy57QX5jp7yMF71U+R9m/6QcP77COpyIDcIV
pgL9wNEv3AxHZo2fqP3SZizsFT89H7GqcdhhuN8g0oDCFr0r4iV+wo1ZVBmOOcFF5+5lUScC56/j
m/ug9A/GKX9GX6fHmuSsIwCOhn46YivTVZsaOtCzZBnZik8R0iBg4yQHbr1284LWcbJH9ergdw47
HtE2QAtSeALuVxpXknQZW3322DO6qVRPGacseMXqF0uu0FW+mmWduK2jcnDVahPrD0286LdO5dwP
lcDtCkkXEN9K0jV1+2yUPZ1oNB/txoThCoSjtl+CBO5+RJL5faBfQn0MBPZaWVJ2nWk65nYdn6Qi
lBkpuRhIZuGAmL5F6p3GynnD1l28+YRzNIYXfYXLZ7egnVNFXPDi51VOK1mxzLlTmJTt71bjwBiz
2nMAOHIZCPNqtMuEozyBL0ffRHY1leWyDYF40JUjC3UIUuVEfw1S1V0MFPlZ7S5NylzcqEYovvzf
tu7B5H5qBH3flj684Ysl9d7/gx5xEHBKgPfNRgvX8y7Z65SMILWja68mgadC7nIDy74JCOhxan+t
r6VNNJVFgu8yKU2SG7Gwb5DyYzbeZbxsUto6lm3lF75Ln5At57FocsYf11W8dkl9pTr/8Vd23tKq
gPRPAhXrmPZAQmVVJEJQaBdGfcSmRpeQAFbxHUUWOXJcKa+PQLijUfyQK4e81sD9wS+O87H6AZsK
GoPeIB1PYOkmL7xlnv6DtSXoAJVTRZe2NubyPULOs1/99LFmUqsySAM5dSRjrMj+oi47VcxHe/8C
vwedFOuH1hIXpDJKddiLmnd8zNkOo9Q2Xs6fd89+CwPI/J6aMZl+lnUJByMy2porHyRA9mEM6Sph
YwIwi9rH+2pkD3s2s2K6AmWNYPuDkQ+Y/VJqPRVF4jGnCCZsBKw2C4OOYW28LxXKw5EA6h5rY358
0TE+bpHZbPu4Z+ZMje6JWek5FTR6VYlIQqWbX3UJPpbN7K01eXbBEqZFnM6GOLu14W6Qjg1RHO0E
VJhJrV2UsO2C5fPhnG0POAz6BRxWxLi5YzQjocSQJut+OdUhQPLH7S4aF6crHqtj2hFFuGJgMiqK
Ad25OmKw4DP/m/2Myz8VY87FpbS6eaaCiXh+v2w87jHj9YU8JXvPM9yYbO5+2wprYPqypsRxFbpx
QYoeC15Wp0P+4TYAPH77ZCDPLW9mJbLvS1qn1D0AvjuNV/i7mLGz20UDURmIi8cqbF2JGxAWd9uW
8LP3UfbwDlUgDMQJsNiM+mgrdwHd0Cp9gseNRWKpyZxI/sqEYHEdr8aFO3svQVmB8TSixjQd2tPb
A+1B9xKE/dAWvgpGvbmBmnyNZ742xbn2hbcEos5mEyrstu1Q9Bj2om+inMTCo63wUuFm4secvqHN
ApeptrOxHuF0Sm3OgPQf/8EjZD1VCV73IgNvOc3yY5h4oKbm5DK7cGy/vHLshbYqg+W5SXoHdLUc
UoVpPG7jrJoMl+PdVIx0806jWMybvl2l7IZkPDo8uk6YaZ97PTAIqQesygSSaQ76cmJpxhdZd79S
Pliv6/5xTOFNRIp8POiMYqZyUVYLe9ao18MMxKc1fWsDBqYCxqKrcJi/ircFv32zKbdT0PiDbkrI
88VboPpg6hO7VBGNtktM4kwU6UnfOoMz5hbEciYYoWm0sF3EitAsMwePM+W9xbNihL0sewUvJsAr
A3nu3ZjKgdBTWk2ltrvX/Lm+lX42CSNgnguLoLPOTMNGt/I1D+pH6AQAkimyUuMCP+j/bPPGMW6T
DtzXWM8KDDtYwavfdEHwY9ibcHgmoE3iIWGz+OH5GhrEHqqNhjhE0+N6QPemHnVHHI4iik9G7133
ok3I3FHnlsaqve+rePt8Q8f6fYpXa+FxcHtdDc1f+blqqLdRhv5DSy6+2A1DQRadIdWqvXUFkouO
b2nSj7A3ym0ufvKl5V8HiPefofgO7EXTLrfw6FQSQ08zEmB5fd3x1mxZn+djtUpmZ6GjsxvDamLS
7v7lq6ttT6vOVNloVTSw/8IfeCWWZJhWBT9zuc/vIvSHBNdXVYIhQXAtXhZ/uRfYmZU4kUKQi8VQ
FaHadh3hBdiJl0MezYWsqvw5AjXtTxpQMDVTfAFimZfxrlS99c2B9Hc6Ib+qq7TWHIlyqlvto9yZ
h3V+zPsUl47gDje0YvcnljROBamyiDXLpxS9ju5tqH1ti5QjEJvotSSWmZGvr0PWmwMNaejCu+kE
T3UJGhLOI6EZUph/qfnrsz68hVXCK0JPvocdL8WJJt40ajVZiTA7kV10FgyJKf/t37dRjnIVcPay
xOZFRo+tg4aiPnMYensINtPm8lCb26SALAZUrKQcTrUK9xNl1ltbaIcEEQc+IrebvX4OZpHx45Hw
RzTRRYYrpNfK/T8eJAZYwaKK3iUPcTvW4EmnugMBhCVs/wwrwLAMVNlbEzk3S8BCQFNqZQpd6uob
ZMMTYvrJBw9Vn7cS27VCWQqSFNdew9M9Zj+oGyHKFh0wFRB6iOW9+WYV8gLvx4jk7Mokiq8+p+Yf
2tjlGplPJi8JQ4g9CTpzfaMyjROh1XkjOG/b0cbYZaZjStaII/I3uu19uRjuJ+3H2UXjSG4dYdSM
uAfMGzZFymDNwRKn5XuS8DnXpEbOlKp/eSBNLG6luFZCqbx74YXAbLwe0S1MlnpLsbs5Yesf65bZ
N8U0knFigdtuExxAGvLSnMu9iYt5MHD7WroSDutVhcyOsj8siH7+0z0ooKQkmYrHvTF01p6W8h3g
cU0gqlRl6PJKZl0wHRAWGR6OEEKiIpZH1BQr4DlrxlUiMEsmtwAogMZQi8zq3fFZ4qjNEL9XTBt7
jcSfyrm7FCal7gbLi9cXIhjM31gAZV+ZVrTb+XIp6YeJF5K6fl1AZoam80rNwo0p7lFVxG562Xhm
wyUAkzQQYPJFjgQ9Abior/exTRLyaQG8jrHwWo85ii6ve6OyJ730gDkwzQ/KuLpXmFJl2hCxCjPS
KvDTgEZDtZw4NZcppMX4OmmqDq3QlwdCNOLc6jn/dCosSMBVVDGIyRtSrFRDGnwaOeb5j0Yj9ZdO
GW76ztVW5a4MOZnTAC/3K89vO5pcytT76kRmS800flLgMEt/aIll3s9bHswZnkXNJHNLNyVrFLH6
qXix0vzvBwraRaHcfz3q5n7MI5piIgkjgvhGf73sVuTSKnIkCRqSJkv1Weu7qosb8+42LULQe/+J
mdo2YieDiHMrtP6FdJlUQLMAwTsMygoJrIckZZCSPKOtvgoyDCL0OpIhVNDZo1jgti7/oz0v8OPB
0CKhmZofpKpk+TU0InG1APhsSfCg92Ces7QGJc6amm++OFJAdw+QsOqHw2b2OeFp6WuzNL+MfGrx
Jr/GduJ2TKTDt45LWMzbT/Sp+6BxAFc0FTzpEi/0r/0ZmtF31lUYpnIrWWQX46Xq+pr0BsWq1GJi
z8n+YBvejoHyO3fT5JHAFT/A2vYgRtvxdMcJmHmTQ2ZEh1lJNsPz9zWUP1tCwQvYaj6XuPTVWAlv
ALhVwa4otXauprU8BYJmno+GeUf4A1Ku1DTqU8vUY/wQGsbwxCoM/qsT1z6o/l66WedtclFtGD/B
c9dxGMP6tZLvnOMf6WV9u1dr5OJw6X0sDSHGJ+4Swa/xu9pHIpt6KYlx/sD9NxAKFBzL0kL0MWO0
TnMURXgKdx4/CWfzUvmdIcOYkPcTu89faSnz347tMSmXXSv8hiMLXPiisQVNwkFSyqT8vE4zXm8i
9yHilIkEtughL8QpVz8WhNYo/8pIA4o7dm1qM3/ZtuUgJsemQeBK16RffZH6Z8s8SxNSN1fC8ewc
gk2V5l7F0n9WayqV87LcT4Yi1J9D4jh212M+AXfOMC5GgSeW+A8tx1ndpwMsr7plTWEjFbR2BWWk
m7jVNjqKQcQTqFMXpKvT0WukN+I7LbmMkmCisbHJXv6cB8Ez5htXwuoIeiDv6wBdWDyg7w0IsbgP
ccm1HFbTK8jxqXLPzBlHe2XFSpj6ucAaK7Gl0HVc+XTLNsLbNKVNPH81IyEN+3kGnK4JYllWxS5J
ptap7rqNqqjgsAbA4TKdK1F2KToD9BH0AvLj0GQdxomBUIgonnCjl69Ze8BqmhsJTthZZOuSgtyg
1JViNULREgTO6bSi5r3nyySPnRrVNlyuAvEXGei+gVOsekDj1zkD2crBqAGIN6GfEzYY7chULCZT
z69sjyu2gK4wNxxsCCPYvuhqjTxYo7lnlHnr/1pV1qcJZd9zeAeTOVe1qhULygxRL2XXHaR5N3Qz
gGgLXY8aS3cW/z/QeZ+Tkjefl8R+Hn1hAB6aq7bSXopjjtT9blVrQplw4hR0Sda5k/PnrWwXyOYn
j07mo25vjVQBXeIEupe/QnrFYs/TFCq1P0CMkP5ZR+ia8Xxlf2cf9Une2CChS4d2HtXiF3Og6//E
fpEC8Q439ZC20F8BuU7y/ZcBNRuHM6wLMJwtFsU0fARyK3pHhIMGMBrYUTo4N+TtvUK0DQP9GKTR
7MEAu73v8F2K3o3eIkl37iWGDtqYpDRISr9yaiSq1PZNRjAwF/TyS/+ayMbmkpFWZvDMiFzvt/II
5XeZVBN5cc/GG62IZ4V4/oEhJLlaMp0b92ESzTomylhGBYurYd3VTnSNrW3UUQurrrTslWGoEGqf
dc9sBBu6CeTktQSTeFlxRL1ezKUC5g1C61kSQkNyXwbkUlSKIEGbDxnomeqh8kVEotlRxq7JgLIV
7aeLvGJKW9o66FmCp6jMcWAkBEvSqnG+EG6lNh7ahq+SKCxiKe1oo00BkIq1VF6onwYctZWFJ3z2
gcQ1UCRJ+9Wo9sqDN8jyFKNhwXCBv0dI8/0RDB4OrmmDSn7ap7eCU5a1cdJ07MsPU61F3SVRZaaH
+lF/eeoNjVwYdQQJHys2GMc8v7uwpMsUPq+elYFk3AYDB7liY+eSz/chvQhXidsQRHMZBtqS757n
cJOy2lrJ2l9lgFtInkUXX44XssjHeH22h5yP6F/nAp+odaSxrkdVw/SltTSgiCmhQtj+NwFqBQnt
0Rr/TYEtUXgFFlSJMKbg9Md4eVJAkoFaQEBNsWbbzfYHmYh+qoNbzmAm/d4HuJyyqqWJhWTh0ZzH
ZNapVm8pCMdu4E4uWky0zAOygi2WdlUY6mIh3l8OtwxhK+GV/0lr3SFJ72XrNJKGuuMFPUVYkomE
KrEubTNd33Z3iq2pyw3Jc9dvMeoLMK1Wy4woqQaJb9MfDIqaTOwb5iN7s5TDKqahfp4wVZg4XMkv
3feiFTaxe2fJGNjMyW9QCN64sfglnCR+y6cGxWGGP4cohGP+gev7FTIttBJiAi8V+9AGyx4j9PgN
MAuBpQGQXz4MQqRpzP/IRAdn0DUaMettXwLNO9noTkZF+fj79Gppn/GlR3DApPAKiGIEFMYSnD9K
9MXFdN1HRCD+pzkE6f2IgeE3YdLMWzxRPLFEpClxeYBkWfPtqMgoaNRyJur6K3BmXU4kNOzYvRum
ep/UxBgG0Up/BaD1nc/I+pnjx2brRgoyM6K9LZlm7RCi+s7k40wjOponGfnioHMLgX3CrtuqlPSO
at1wrhzzE/Mg6ju0aS7vFEa9OpImoEPpco+sctpX0i3zj9omjLXNUnM8k3BdPI8LpwDVRrito3HI
OwgPzW7Pm073g4i73sZ2RcZbLlXJ9q65bRGi4qLSpf4otquOQarLT8wmxL8tL66Q3PH4T8IkOx0E
1P3UacozQQxZyVCCNX7vAYhKFCiGsTXPfkQ0WbnDJftAHH0atRVBeXqNRA7yxnDB02RNlrPAl/sn
Ow3YrtsRAVvg1TgFLT68EB6hx8DtcLo7jMCDGEXpGkl3K9q3JCOfL728HmcqL8rRDqNVx3Gym++J
bDoGdcLAj9eklrKVpah3PCxkM+f32W9kVGm0ynjDPqyDVU2rC0cPzPAn+LswGic9oiclEexpeYQR
gIZSvDrb2p1RkjQBx5S1hDXNSScy4LUOna05eszNUUG0NEdDa+SzIbZjHq0yQ0bqkxmdNI0phRkl
S8HTDgi6HcIyNZchz6wnFzhi7voubm0ks1LY5e8QDRvC7ZCR5Vb3J/zyPV93ZzfO4TZBLaYNSn33
6ImVOtLAUgvvmPSYerz32gNCZbQq/1Zte+3eul3Wa80huPyIYSGdFkudnQwagCevp5nB/Y6jdmGM
xynWAcC3aGWCp7zmeBr0adAbiyScn+gSmluK8W8Cccu1AnztQsKwxnALyrWDfj2Cd+G7JpKXxYcl
TTvMNpGiOcXFEPn4rNHi/TIvgM8V3SOxiBp97yeLUqXoyW0waiLQCHqdjEgQbA8q1mXhZBYBLwGP
hgA1gftzg3JPeSvKyJSPKqayMTH0dLGkVwVoFPy2L8A2YdzqCWw6oTzpAQXCsUYdHLgelWlh0R9m
dGBgets5wAOGIUFbRKzXiZ7N/xX9u/d5IHlEsZfbjDSXc9mz0Lzm15GFnx6jl6vFaTCAwcNcmHyd
Mjn4EyoYNELG9ywt+0rpPLwI5M+B1GY1IEXksi6aTq7wRe5RdLguak0uspRvyMQtFdylphzELyA2
yHPvQ04eNYY2FPPL0ZxJevdtFfe1Q2ZHT9YyCyIu9dCnzgjvGqrEdd2PPtoDNGCi2aM8LlM5di2O
vPBZr3BQtdYnlVV+hn8TlXptGqUYEl7jjCHQUhe1Gtv14u3Pa7M+ppgi/RnGXrCj78o/XxL/2lo+
o6bTlwyeZlzXu9AjoK9lgPAOWM274qmT4A0SvwOu04csF1waJxNczEMNnQ3uMqz88qumMWiURFil
PfkS2f4CIwQvos/hK5NA+6B9Tt0mmNjU2DZWD6A0Qft5weY55IX/ItVAmih5RghLuzh7WjRScdRU
QTxIw5eH6CCYWdLQlrA98VVFdqqoztWi4LI9lOzlAd+NK+NkhOiBFvUrdUpeozHX3FaDN4psvcOz
lOgMmEkeTsb13UrtolxMJNmiAYjbT6KkZesWyyFOVr782nMSUtGkohGV28+H1eBwyVds1+BS5xd/
kWTUgqqbC93A5+y2Jm4Y53FbXc5JOIF8JbVzos6nGXUffSza6Tau2uWJYBAw5D9UdRvWRHOTQL6m
m1l1Mkx2YtClDwghXxwhsdfYlxtXpsjeejZ9sazzLMzAweoxx7yZke97Mq++M3FZ6v390/oZmMs+
E1btEZztW370Qjb8n7Ujp/Vgyfc/9qM4WbV/6SLEjX5ji+ZWIg2OKgiZ5q6YsJTbRNHjEZfKV6rT
sHfDqG3T8TI5RWyYZMgjjulWon2omZrlggrdsB0gb+ZyoFEzdwTVa7I7GxY416SDbyzADHUSrUgz
iMkkAJEVA1DrHkyfF3VxPAQNI2B+OWoc9hjLAGDQbXBNC0Q1SyZK+Yj9XfzZn2m8PVsgvnmOF4Yc
omYuJnz/R5dIVr+15NxBskf++9TWeTETLaTC6uychjW2Jd5b+b8ohbfpHLPZRBTMDZDd5zDkXG0w
S9SYb4l+6Q1yt7eVuVJAKOwpbh0DInlWD/2flRmt+GJywBxs7THpA2x7RmKhTne/ymreKexwpCQZ
/eczeMOGw88kLg+u+GFuqgwoxp3XrjzL5akZK3Vz2/z+KAQWyhJ+AzK78sAcyId0JBQ0N1AMyURE
RXVqdV0kycq1Y5cXmmGoPgGX2m6uBoj2J1Q/I1l02X3o2LqmnW9PP1ElIJ6W2tzIUfk0Ql0j2Obf
BHotaFxeBvHr8TqG/1NDfzDahS5PFL2VXaqbf2tJDE5SzLCzzkJ9mQm/ShJwTl6k4c0apD9BDIHO
Zo5C71VTkrsU9Nqn5AmXwPoElSQSaPuERpZj2emluWlj2pHRmRBoj6yTrI/J+AJxYCU4sNot6I5N
8uoV8p+6r/u/hXB787tP9ugPPa9N8O/dcpRoCel/u+lLphTbKpw9rfHP3Ec+7ZdyUfYvzlrJK7c0
1HrXPy4Q4frDSpYDXKsVrGEqFDSVLrU+5sN1QaVy/wcVyj1KHJoMpkbVxUAE7ALagBZ3DAyr/c6u
v88xab0T+uIRn5+k8PNZDKvJcduIbsnOWqU4NIsaGRl2qaWvPy9+nhGeR85NEKWDXraJTpME4G3S
BVifsDogr7POIQa0Tnt/mY5Gv9zgIwl1o9SkoIbDXwuAOf2gkuHGKT1p2kXuyfF0XAs5tpW9Nous
HcM2YlgpVdEaYgYrs3KpNNuIC1MUTDuJk8CY1N2DsXJKNJJZcrbECaCv4jg+YUjUJIgICPBIqoxD
jZstHPqfITgqRxTMOzZsdGWxBmR3rX7pSVy7Uzj/cDiT11imrXbL/CCLwQAwG23bW4nv/hunm/f/
XgpY8EZxHd4oauFp7yGnaGaYC54w0cjy6S+QQ+M0osymkmTY0kwyf3CdqZNWuRkkcvgTcXjpp2Fd
kDtXpJYUqcc2i8EffunWZ2Do/OS/77OtUD0j7yhQB4Sk5SFrBwSDNAjrPexBXywe2dEEp2nWjUgr
qxNWFVVw+oHY8aUbn/ztWUU7Nz799s/8yZFteGMeF5SjK/QFk7hrgaTCsDpffgk1rAskTNhgHc/G
V+VO28Rjz3TnNkn/CHaz5EVuwryN4mp40qeYQj2Q3rb8AbFmVxkGmjSvj3LnCXgm0mSbZWuAhZTH
VBZnbUJ2/ns/Enw7vxDh9LTngUy3evQbTZtOqsLXrj3cXPV5AetGT3kPpuVp4bF2AmVpGofs1x4X
vx+B3WXC4fb8lw81+AO8ASbPNm+VX4OEUSTkEmmkUBUoTDHMwouyKb6ifXrkrZSvxEu5cijb3Lyx
aw/ZfCclNmtOuswjpNXPe2LOLHkW11jMGctvXdHdOGoH+JPlAiWSV645cI+wZLgxjS0F/Mo8X9mE
hRTvTbJqUMWK2extKR3brF634qJYjAxpvMf3ttKj8QBoC3BkkKxUN6guv0A3M1+EBLZI3gb/BEhP
/D9B8XaMGorhTRRG4Nwjvz70bE4kPHL03Z5ea0gUrpsn8q/7UtNW+Roe1RoHRMzpOdDXQDdtB0KU
WfIoBLxd3KowR0KT9nlItGawwaI22FPC4nnqzj54vGg+P+hUvgjlWvxPXyVkNuLIaY0VBuKUdCJn
tZMQJ9/c71sDv2EiBJcjZqPKi2jti7vxXwYSeWpPAZMidppGrZNwQgo3XO7VBB3lU/womnN2wG76
awUeTomeuCKPe/6UgAfTOjjH4uoAfX+LlipfrqyabtxzTPxYxDqlg2rT1zBeQ0qX4yiKO+h4gXNC
kStSqJyX/x5yL7iGnFnjuT+iuEzBYqsx29RST8cpQ893oo1d1cpLZzooMg7MHLNr6C2PFEG0e2Tq
KV8spcLBVuLlsoHcSeVHPdsy4FQlupYkPYPiTa9IjDFZOcLRWDJuHUe6A/4lPcl6DzTPdOOcUzzK
paSEm7eO8t9Ip5vrBrM7gn9dt3WnjgfUZJGnWydyHiO8pWyJLVRLrLKBj0pbaKUHGYsdG7xdYkuB
CabS7zu1QZTdyE/61AqBckHmuOESJRUbdWsTE/BQ61CXreN3PvAelWp8mmRAb/d56QVz8Bw+eGBu
XI1TN2s8PNwmXQevUngXC1OvPy3to0D+ejbgBJYVljkDlktgRQjcHqAqfQtd785kMIat0a7R6zfX
uYinwfPMmsFvcqZaNN1AWrusCbE9i7IejhkAm9exA4d+WYyPbaySGUo80dEu6pH5yZYjwTz5k/Xi
olrsPpB0c212EM14jBVGAoXpb9+GK6FzwUU4e+fsjar12tDOSug/mSnPYYkfQGRga02lIQTmjZhp
2D7/X1okHrPwr7HoRZNpI/XtyVFaSGAKUHJwU9rqrXaxHX9P1f0/UTY7N6LkRH6EcethPpnXTPu3
b+ZV+W0Y5NQXdwxVydx6e0nd8ggWjgKar7aJPRJ6Upc1RdgjdllajZ8Cgd0kfAnvQYQdDYFlG6v6
9mFv2cZwqeUnPMDY7EZj1FC+Tg8sXJc6QGM5/nEySc9N8KFXSDURuDzrIPgV8+WOw8YpLYU3CMaX
I0Zm1k89J7ci+oauIiPL6+wxjLWB+iGo4Jx3jcJ+koLEG8i/XWTpZNaMkcZUbf7s9VKfeD28nzIX
bdUh9TZ60vM1N+XSx/xqUTM2m7u2GJr/9foRCAaN27cYeuUo9DcHDWn5AnbL4hea/nZO6gY4VgTt
mWW1/SRePYNjUbMOeY5R3kIOfAmmEO0cy20JgNCaiNUNEeCy3ZMZNiYaorZ6h+aJhRgR9vqtSQft
FRjrRqr8ML9LS04mmfFQjlsWLt8xOLBrGLHN25WDPzHRiYSaiw0jyvRTIB5mKZJCP/W3mUtRotq0
gkLhL08kcJpEiiT1SWUOKHQJjUsCht2FmTQIstR3R5FPyXF+r1IK+RPlfnBI91viPyfyJO8fEYtm
E5021v7KkfR7kqGFfZd2Vb41PSFf7WO/wTybmNUO3mrmOVtu47VBTcbyzTBDCBQDkkWFSNOFqWE+
swMHIDXe6FY2nj8bCSmKds3rODgJ8aUOzqkW5tgirCkpFq537VTi1KfSKb7qOC23w/0WtYpk8hQX
F74M2KVWhdsR1KVn14owgVm5LdilIuVmXheS1b0l2Xa9Soqxme9iEASudVoNmyH9Qubrr6KA56GA
M2+siA4agf5eF8JP2QPos6S2Jbs9eInAjshaiv2jXlxLDze0MoXjNyx+zPYlzj0tKKuX1MVlUfRp
iVWZE/4pZTiLTynEYYfSoFsdsd7NbSIUqWlcJBMJYT39zM3/U/5kV41blzWNRoUNzW+TbhZupY4I
InfxbqY//yeWCmusamnh82YbfrVzMrH8K8u2ZN9yHd2NVHzYGzlhSTNo0lY84W7WDvA1/mV0Bcue
lXuw2acLx7mHjrbsi+W1ahxXN2am+rK2rvYXYD0krx6ZSFHScQrqT0hJQnjVH3wMppLteVv5JUej
d8Qg/dtvFDbAfv05M6EHCiL30Nx+vr2bivU6tGje3cF5SkwW2hk+Vc6KlD7UeVDyPAfdi3DukLTt
GkP1bT0fftiF2m5LsOpgocjLx4jeSVf6O0/ckcXUL+J5Cx2YgitBJCPbiv0BXTejN897ElxT/nCS
At7yW99URm6zbd4OYQwG08T6Oan4GM/c0cnSx2C8Abp+Cnu3jJKSDrtRjltHY5VeQkcvUFBIeU8c
XLTGdOZH/F95xZWzDNfSGNO6BBS3PlugSR7LFSu0bXslJO+U7irAgbjQ3RMK3Zd67y9Ky/OmaqL/
b8U5Uu8m1rqAKLMAztQfGtCKVz1tEjoPZPkDTWqGL51CyLMyBWJHuINKKKioCcINhqweCCzC9VMF
v+ITlPqEBoYG51gvDrDxU9CQ+HhbprYqsrpoUykwtHYy6ptrLpQ8pmRgznFFdzXC9UBVH6YrmXmM
FYKObRtZHMrLV+KcQRpTkZumpODMM+TxKAt+eWT2Sc4+fnS22jgtTnzsRyAsxU3w3uItVOTBAsiG
SGxdoLaWIF9mPA7mHXcnomU2P/VxobqLCDmnQYMmC+um4LugsNvzIYNdqE/f56MsZwMELSdHjF5l
9EApcJamNerXNQdrmkvP6VIIGLUDBDmtvcKC9aHI7DouraGvoYdSqOpy8FbnQxseDdUOhu5Hhoeu
uOiYhBLkcvNj/093ldH3Bjltr1Z/dsK8Fd1/txOwBxbxcWNBg+6jdmFF1kQa6niJpEglssKcJluZ
HrgcaKcN4l5MrRkdPd+zxl/bjnxXeg0stHYHJHeHoLpzYf97cypCFox5x3bJczqVbULadgeVIp+5
uPLOjkibJ0ZH9CoAS8be6L6/12GeGIlpCrgXNq+fWMvgejO//L0xtmCVNPMKVhUX1Z6pNDsyEiVi
Ji+qc/FFkGVM/0gtLK1gLUF27Sjz8ualuUYbiXKrO3+Cr39kzTca9/QxtZNhDNI+5bebwrDS7LTV
bJzcnpq9ek+1M3jH9ZsJ2IQiqL91NymVF9Jl5WwT3u3mlQnusgu5uzfdPY8znCra8mMYzfD2iD8W
Zln0vDI1mD/+Z6ydMyWwJ0ethYiNIV+DjNwu1qTWVAPhL3zux5yMxqfSuAZyjgODnzy5xrpUofvZ
ZJFBeluvvKDzvukSMWAOaS0YXKDLqPnlYNf9Bm6pI9+BhmH2fZui1l1bgo//7XSaHOl8OKav+ucS
z1ZuiV6hzNHBxsq/86fxZQtdOMWsQD37ZyNP/s4O4+FlT70Tnxa8cRwrRQts+36X6+d3rtKsVsHG
rZJIDPHaA4z5xazFATDWERPOYvzo6wKj5WkLVuoRLf4jIm6OyMF99CPrqua2F9GEPeYUIdV56WSs
azBgYCIC5fTnFRaIrAy9AofVm77Og3hcesfuuwSjJX0NYJ8lwwkEBf8KddptPUaJuc/rURvBHhRw
YmSA75oOH9xvANLPaEgFDyW1lJIJDiXOQ5hoOrmVLkLUeqWGJJUV4NfEQgrbjQ1sSe+RrEFwDug9
Cn41Df45a11IfBQBLCQcEu5f3sDmaCrSrtww24mnZcabUrMCJSxb8HDMRs6xVcTVN0ztd84VTHlq
KeBNLeVTwy9fcSKvmsQ0HyTlpUIRJfKT9VkMpQrjq/MjHuX7zbF7lE+GZm9N1kijJ1967yjkJAZ6
nVt82M3ayVtxKZLVZ8PI3mxcOfB1lrmsAR/2XnAFyMD37vftKhDiNjrrq3QFWYwWsFN0l84IPvKi
zlbZI8lBjiYw5zHJ4NlRMTnB+LN0SS7pFp4xNrko7WJMftd02ZUybK6qP4jnrDltsz74rPiu3D13
9Sr7IqbVdA5fkDJVQz06KBYgjO8EOS/dPnZGkKUFV8LvdfaGjYi2Oge4/h0sQmWQSEeCPhwGcfIt
YxXSZNrdWbFoT9MSS/ycEcqpM0s9FMVqQlAM3SgMIflDF50DIUB0tlXRwB+xJYIWU/YN7yfPY+tc
oADmq615qf+X1OijDLNosPr01FvsTir4l2LAOlN/OSkCCFvmUQvcmwqPUmNpNFMcWHvnMIH2+TP5
kvhl4Ssce6WntBbP/FIGLkRORRhUzkaeXOSNrBvLQAk5Fzzq+J0r9FsE8xWjXIwr9VktL6kX7puh
Zmuc+Rdt5nM3XrJAY6rr7gecD6uqO114M3jXwnbzI1enDeyxzJAymwmv4lrg8bBI1AfJe89HuzqA
XVFs0wfZm2FThsxd9PT/0z/gLuboBA9P62eOXjQV0BWjMnUZqwj0ej9nHNqjJw6DsLU1sdERwh5S
lrH/dd5gQft02ekX6iRJFwPe+X8A8syARQl26zDjaCIKfczFYHnUpMy0koyNfWSnuBMCarwleGKA
/9qn3v0URfV56nQ72nVcTO/B2VtHpkvMgL5UHCafgjjEN4rxg5Sd72zgxyXQWkpcH36zIuLkoz+3
z7GC3HSx01GYqGgFM8KiLrzU7vCCrYOGB5G6xO6km/seQTasrB0T9eW+Z3rbxJnBIIyOcw98QjWG
h0TJLsYzFim0W1bXsoaH9wrLg6Yypxrm0C014b7AEgM4GrWGQ3R+0TXd8TnFQDggufVTJyj1bo6c
0OjXpLpeJwPjCNSOGBPhVozM9Cbm58ncft4bo4eTEoM1I+cNDFbM5OB07ynqXnuW2iSu12FRp6AY
f9UdWQArZCzyM1c5bU0zI1jUhxs8bF3S09KhdXJuDW4xyPds3zqLCduUf5EcHZ1iOOCTG28i8cod
GsBrI8w897XWl5/G+/1eeTQKMgH574yt0Kad8dyNE6Z3z6IqItY/i8J6qIplbrkUZ2x4vjGm54eZ
Df96w7RdNyCmnbquvcVcfKCBOdvf0Xqq+udPwW3ZDT9RIhNFinUUGkQXJ0KKI0CIJ8ZcioVdX6uD
c8buI+y7c75zMzr1N9anl6nWCOpTqbVA4vXuCRSh4LE55U2+o6nPyoonJ3ExAu1NosKfH6Lb3dZy
L/WLTbZkHas6EsnwyuvmTWH2zcb3qEwV4pcge0JGtziYsy0srUBLkzQ/bNdUWCIOxTxBAnYXTIZW
a7WnD4+CmU5/Zh/AVdUW+GuUwaU+eQi0vAujLE1H9kT4xXwlNykkVkwBzJosCkPjzzYaOfjZeRa/
ZjTFHXZit2TfodC+wCYDqEQ5lNjSf4TDPsZVUqW/Lcdv22pFvuuCbJLuBiGy+Fhw886m4f48OMiE
QjS3jhj34KhIE1D21JqK6swODZM1ddiumEEu9FU84y+EvpvHL9C62RvLnlJzo70V3ggFfm519ovY
mQacrkag0KplnxlX1dfLHcUkAqhRATuj+sYkCHpZKN/SFqrO4Cw/jOV0HE7xIMSX9M7ZKprRIABS
g+3U5Ge739Iw36YbOQpJ2BDWoZJP/fA+qlCW0i8P3M2gOOEAWhxH/sliM9KtKlh/JMI006nvDdJc
mUu+apem98wkG0x/EaM4gED6VvP92XLGYwzCNzIcAT+BsgXAakYUBn5KezFCeBaYgpT6vDfOALrq
qHAiRLukNxDeNVzgUb69OY9cg70iViLDSGwEWDNlSDexTQ/UC1SR1Sas3HDO0v8hwpXVeACq8E85
LHmM6Kq++59jgsOx3c4eBPvHy38O4UydR3y5IhwdT/QqWEZlhbCm3oIr689s0r3l9g4qW0ieykNu
jRX3g7+cFlrUpS/EOCkVcAs9ZMCWTWxBHahAi06MyKGAYSnkLqNoxeAhWUOF8sXCqfzwMaVPzNpz
FSGOILKsR+RfR0nSvHsa9ADa+eivHTppe0jhsRAkvb+u1Te4otjTcDfuoBaQuPMio7xHlacF8VvZ
RRBpDUAbnw6zCmOg8MT8hyF620OQ3jFyPqv3lZfAoC6B0mzMEpKK50b9vj9A/GjEVQFp5KfA5WIu
7xf7cObZKh04LqXPb+dhH3nMZs80zsV98vyyxc97XNUK929vThVkI3pIJ7T9+6eoZq9OGDh7lP0f
gWhC6qiI7jUaq1RgaiwYfy0yaZuUq0OJHWS7wXoR6WrYyv5/G/ruOeC4jSvoBZ+cwG7mt/SM6Fla
Dj6rwUJ0vS89FRqa6Kq30ZjSYnh4bW8PF/lrDQ9P9IDV+h6J6sqZzdOWOOPLzFH6emG4WqUkm6bz
LoGrHuLW1/zNtpJmi0cBhb855w5grcoIOgwGgnV+sJlNjOfxDotMsUfyLlHRzREKKwa9Ox51IMUe
FxpIV85WBWD9wrWDxmPEQj5gsucZ+xf8OUQZMSEgUfSKVLuk5fJfaPZVxXH5uc61t4ID1JZ7Zi/M
35WfreCWr+ywNZuOi20W4bBlwzIj/052hZQWj74YlyZ3a+UbcVH196T9ItjMAVwuRKg/DmKijVlC
GHxJvQjYkiPXP6nY8SOUZrS3NDEIPsbjSBB5RSM+P0turhfNZsiUx10uiWE/Frn+yGOlnxh20Ig5
mxR1xQ2QoYBGrWA/OkrKWcM3IuqrV+AhTFRUdyPq5vZhglZco52mf3l//E97ekh/BtFQXdKtN+Cq
+6hml3C/Yxxnu+DBjQRBEb4knBfROFVcpRqg8Yv+YjHzdJyVGCbVoPPw9jSC4IKOYHeWfIzxq6gw
BSCcPArOno5AB7wEiPbtHsRhlR5pTx9/hq1S0P/H8xuPvpyOwsgW8piNUBOS1r/uFKswoSgTHNQN
2WI6hTrr1JFf424Err1HQ1wJbXyMLMRrU/aF6+uAlOz+WWo6mEm9+vbDzgjB87/32jVjyTI8ONxd
6/ASEfbCyZu7KrbMpxSbp6EDM++NvLpUwVpgZ+NawPKcW3yyJu6bM3FobSO7asWdTr9apc29xcsW
p04HLg9XiIPd9wYq9qQ+cQ6PLxTFMPpGWYpytAT1jK/D7fYLDySrkUpN3YDm10T6tiU9nmMsyacc
K9ZN9YXylaFI4CKF3r5u8Mx2vXUQhxFixrQNGlH4Ho4vD1tcSO80OnJU1Bq+M4/2OURCgrekOw+I
aPCOr7Q3MSzMlXql3zJbGzXskeJu/vdRyP0Cn8fVQ/JZPznpGnxz1RFBrQV+1d9Ob4xHnVqmaB/m
HmxJ2Sk64P2gGgxLemSiFn2vD21eis2N+MHKQ/1c5OkrKgRVGWvDS4WjbTlzM09HsW4Ori5/+PTQ
vZkWHkspCavsPVGXRYChegPpb5XoSoygNO3c26c6uB/BgWJxqpZGgl4/s7H7ENhxTH59WlgffZR9
ebqO4/Nb474e7208tuiEKx/cMkAmEStny93bxTnREIJerogmtLu0C4dineMdREHNak+9LYPMf298
zkk2bCrMdaetCIZBN8v+4mSSZgDNjLYIF65bcBJOp8eYqNQosoDohUuaUU0yD3jOtG+hVNAW7tz8
ntdlcfmlUTvERMmUnqd06Sw8o91atl+6oIRfIfFAms68SacL5yejiBnwAy/F0fM558VUeVmxR6ch
7y8/YYBl0kWdLtdQ9Am2QTrpf2Lp82a4bcQbKz2LBusA7z8G9dMwKHIM4O38B3uUNLv8raqmGRlk
GD6O7oK3EMwCmsRuBonxpc8fyo9cxZfHrdBPxxTT7gGtyvE++W7Fw3Rqf2/XcGONlhu4R7Kj5Pdi
ruZL9POBf682o7sXgOcDgJtNPg8FDwiznm0jSopjiUTZfNaCtliN1rid8au8yliqRqFt3xy7D7JD
L+1QoMbfvbi/SLp1ejE8WYzqLoN6Bo7+sy6uWSTNBCHe5CvWccsjl9kWe7Dg3JYtQLDu20HaDQEz
7QwbYvYgddsaAtJYrk/e/Bn8yRPTlC9XRHlILAqCYi5SBDejCbP99i/ioJuyoveSZMPP7Dlo0JhJ
K4EC+/FNDXiM0hg6Q2cK5MLeGGb67ME406JL4TX33qqsl+eyHURFPWOvt3T3voERPM7/3seVtShV
IuymspUBFnAvo0lp5ZxDt69K8gDHXzRkC+gQU7R5knESthaDGtnurxFXdCHSmFQ9lcsUMivLu8Kx
hkm5HZtGBwCznkSLr7DyOOhMJO+KQFObbgGK9p5bYTblDrwSW0tBOgYP7dvL+DI7aDipFlDu+a6r
csx2tgrk2QaLqunQduKpal5tZlToE/n4wzZMFQT+Yd6R7mh261ZoNyUSDHhVUY/65o+ubNZUWXT8
Q8YFtQRQJqMmEk3TLdoZ/2Gj3fQwCe1vXWIKfKq6h04YeL51HJSllil78kgXAJWqxacZBsiEl9wE
5XvUkSGDp4sxfK+gbtBNoTPFk2yDIqrUWUppHEfmBQOjQHuY0OdLDJNgRGPvulYtPwtcRpPkXClb
sN9a+nDKlAq4nbaecvr85B503aHRR4qk6ckXY14i8Q+bmPyDJNP8su0UbqxBIVWDM3UJqmBuwHh2
/Ger44VdltsV6+IWmOr/pHytScPoA1nyuDbyYRV2/tfGBdQed86FX2is5Gol2RfEkxGVlmpfuDt8
bN9XJhjMGrxc594fBOF40Isa6tRZBrC2c3wLTJKnDwGXJxAqQA+9SZ8BQ7vvCWycqZvsBngBuHv6
AyUjm02+o5nB2/Z3kLVK163/UceShf7AysVGyf10Toh4Hj8EJVm2Q5RZl/BjfLxTXhMeItVvTnBK
d2guG+OwdeP+nJ91AMhxDKwFkT7uE+HvPfb8QoeJHJzajeQmzJ8LOWG/3R81UowCL8UsNtTBYV81
UeF+jTM+J0Yco9CCdBT4XMeIkG6pGkG4G8Kl3fy6bh2TI9+GKGKi5nFesrcWEJ8ka1CwgSc9pf1e
VN5S5I/CoVT+g8NoK/g8NWdRG7qo0X+/28qWlVnztjLEau4uN5+IiI3vrkAxQbDRu+QijCo9+za8
y8ZS1rlTyVFlTaQJYmEP8A/91XzEeu9C6+ftFS2stQym4Y3K/QpJpxAl8K6qN8lueGoJ+wQ6zAVG
fMizYFZEmZJt46e2Ql25nyPMzadlBXeI+UoZKV0CJ19iUnGGdKOSsCk8xrqN4sESAQVN04oYRMgY
YpAaNU0TshXrKCnixqKakXW7ZcopBaq74fsCx/4mnhV7d712+oJkPtz7kVw88D+atzAfQ4aees2u
sFFTHgakWbiQwZG+anLLJ3HElJioefjIRXEea4isbRfzMXRGE607b8dsJaNfjgaDfMi9u4PUl43T
Q0cMSYmJcpH8CIANoHwCCgarZe5EZHwEkYq2chhkHFDkzfl4dHkQYnBX7JbYbh6Ezhb861Wj4W1x
3lVKuVSlUrVs5KZ5cM398/lWtBSrhGhYGOQzh26zx+h84q1sMe5+Mcl5W5SNhHsC7yP3WdDroUE0
up5oHx1ff9T7MCEsvBoJhjNC7N/sspBfFUuD+6/y2+zy0v/uibX4mlgDDhT42jiwg7ia9OJTUbhN
YU1/bx7kYYDdx74OiJ1v902//iiTUGunBA+NRZdmj0YKYnhhwneOFuFrfVlEci86dg2twkT6XzIW
E3q2Y86MXlATZg8KgeNI3GuIKdZ7l9E9vXhGYgBVQ7NfymB9zxBAXzDoRtR7E28Xm560QYYJQYP4
bILKDm2ulvHmroeiLuuv65WB97KlbYzqNSrQVtu9mPBh2TN1u7P+X5IBSsfXhWfdVvrkyK7HmHaP
vrf74fPg2MgMLz1WHGRPyaTv2ZpB3AUr+9r1fS9CTDNvbDizp9aQ1CplM42eVbHmdedCzKVEcgaX
2FUIhPlXzhRAJ7/a4i82KBMO3KZrf1Iui3HLHLzt6cetBDx3ILJV5F9fV9twaOm2FY20ZJdBoIw+
tzDrf/QhhDGsbStob2XECHK2F2Lgz8CYvphtbbmG78Bok1NaybxedCBG5gSRWB96XVovPw7fp05p
hHO/dfhLOfyZcWXsZddfdKRXeLIM/+0r9SmMHXYEced2pER1l3OBa2OQ8Wu4Mya4H0FXDij0Hisz
JTntjcjIA9ftU+M/p7+cWRcpR+/1tfy7Pw1Iri0XkA2AA869x4HbWcj1Zh4ATbUmSQ1J3jj5hPKm
TBEm05QS4jeAEkGLD5oLYdgap+OViHK7FB9ABeKRKasyc3W7VULiaAvNe4964TzujCjoN/aBKSOj
KFuZ74m4dsPgHOIPk1XN0ZxsJp43ChjkwujxzNfpn65PCgMVWzQcIgeFv7vevN0UFh7iHRlO97wX
uwwmthrHqRkFs00rrVSnMaNk5dz9vC3CnfUexoVrCZHi50L6ONw5DzO3YuxSuqyrw/LDAbGzlIqx
OEHd0E06W85Q3P+A4OdQ4ZAmFNJemr5DMH+QugBcRv5AcNqhWZelhtdhKLFJjVK9Wiu1t7IvlVGs
nHEekxn0uPadzlhqSnb5pwHA8Fm67Z9ukIqUz94JsU6r564PY7y5d2/Etn41c65QJ9hLkdnokEqr
QGkSkKHpB7GFfq0Jv/wgC65KxlI8u7MxQRixhh+ziD0DIFBbYL5LlVpBMm8QnvWWH794m1tr1Ssr
LMBHNyIipf/ekWUbRk6b3Edp961h0ZPaRxnYl1RhgAbM3BizRfLAz/WmFGg+t/9pjC4bJHqjJHC2
p9q+RkxmVOjSkWXrRUvhZubqYyeRLr6r6W811Q6Y1KHiQTzyAlGUoGxLtUzvb7IXRzJM6uVR4Itw
mhjFMaVROXotONP/K1Dm6jS7Rsqqkcp15CEPQN6uijrJWjM2VgyP3xe+sc9dfvLH+zP1pmYb0Rl9
g9G1RjLoJnO/bkX1GA+hztyrKRtihsyCs0Z7V6eqWm9S/wZUdAGNIgR/FjfYRFY3rmfLf2hoAt2Z
iYTf0vxR/+bPuVXRnUUagRQ+ZmcPQssoYglYdOYlKG20BOIoOerBNRi4lbElDvd6UvA2kJ7/6OGe
0nf9b9z0/kEwgWqSdXX6s3gMccW1SLSAnlC48d/iOHZ0+zPWw2+R7j7pvJb9POd+LfVUH2uFXudc
hmyAsN61S5JGE5x+SyODG3aeA54ZwCkk/CzlG9ovWRlIe6QFLuiA69U8Ccjw7lF4O5iPAg1CltQX
CrT78DNSaWwQIBMDSbBRxZMkowKAA4xjD0hA6IQ7t5Pp+pRn4I5BaryzuRNFOEC1bA6djQ0kWNHJ
UAXjxfoKos4eDIi8Z2cQ4xjaU7F5l/mQVXff4FEiYIWA2wnxrTBTkZqMgkH0aE17SWDnu5uu3/vJ
rAq66NqzguYA/IUjiuvTkMoDgUeVQedbFfhqICdCEanT9NsqYvB0iYNygA7mdF6lcJ75u0GHjadU
NhUTvmaG5mCexrlvPnGAWIJAmxbYVl8XZ8RzVPFKcNencOG6/LUk64Zi0nq3rCCM/0UvzUF0x2PK
nnRWM1qn8xnjGoyfibrYkn2SOfAGYrIGfapUrmkM6wAPCcBaznKQEaxunDz8ODvN0EoHEFs6wi9x
gfCjj3v+waP7djPE00SUbSOIHmlqWxx4Ae4xqd4QIaTNyV3qDYty9vVrV/fXg2mB6qdhiiSuTQbV
1Mg+2gdAo4487Cz/ZKL20IwHsTaEqYsejEDyR1tTwZUbUXW45BtEG7wiKMVZRg0jncaxlZm6BOhZ
tKuoojncSMm7qqbZfBrA3qRPWRPQ+Hm8EOG1T60dTXuFxd49D/BqRjrzgqCNYkZsFRnELyfVLHu1
HCH1ICPhLKx/S5Q+covaEaE9EP2hr8x+FF3Lr+jOl3m9LAio6c0bCvs6RqGg/Ko207rbhhTwlBbd
htmiB8KRSvWKBtBPy8rk+ZUZuQsx9PbSQsy1rzw6nr0HBQxJVxJ+ByjWtegron6c4z9KLM38uLZg
p91JZXnFMcxWHAS0IiSIB/G1So9YGSCyc/bIs6CPpiAe+sxYiOYp9IKOS7WcrhUB45ZN+1glrGrj
ceidKq6+qh+djqKCt0ndwR4RyaV3R+mMlkQx/Vz/AX0yUQHXCMyM8jSCO4PwmbytcpXGyXLE6OoK
YFRmqsaBxttL2nf1arm/EK4YttamqkrqRT3xfm6s4LubAy517pcsI67JzQc8n0f0I0aYaOm9gLNI
DCc2NKemEr05PJrmS4LOEXdILC/obVz372JiI0AlFuOJWHpB2EvGHwDBFs/dxqU454eicyPWu4lI
7yj91RMOKQYMOLBMn1yF/vGm3PNBWybXqO2u4A+/Rv55hLli9lOYH2vst2HNXAGdoseW8pWnmTvQ
FHpYZYRxhfIe5sB+Saqh9NQekRs0eNhNTiq6Rf8rpjuDgkwkPNHHW7mWGX5S+WmhV+J9c0QblEyp
JY4o0BiclRPKs8pGAo0a/588l/MKtfRktrq0hW5geAU1C1p/uj+8juOddw0hyyHrcpQ48c+i4dZK
pLPXiRLRTRbXQvthz7w8+IO2YkkoDn4csWSwEurAUwm/DIoqjcuMBYUUQ2Zd56jmoIF+nOTPkE4v
stGtWcNgFZcXKYGs18wGAgx7fMi0+ezQcnKRRpHQTWbVaAm/L6CD72W3b9ua9/YfRy8AcxQWFdEy
kOKeZr4UtvtXI9YcPvxAheLWGPG8xTpRD4Bf1GxXJXoOb1hiNI+6TMIFITvUPQ6YfQjtEM1cRuaX
NVOzjPRoWG28t2iGa/E8c8p5orvTCyRbJS8OVJK/2b7utUdVdFbZ9Zl66Aqekmp6dzDOat+B5sOz
TAkjyabcvVtZBxn06vki5pQFoDJ8uAzgl0aaAfOyh9vpYumZKGJPrbfoNfvC+0CHVVqTULzdGncq
VGLvkojw1xhiFSqrR4KeJcvXRfMMp98/UCC9wqMatv2bHwpUymDU2fWBvwyVpKHsFVVOYx+hpZSH
gj1T9gjFm+qftwQaDZZoGJBpChwlvQyB5/P+3Jp3R3sTWR6AByKzQRWAJCTlntLrfY21EgBNUpbd
6aLjULvXAklO8ZWkrF+2meJ7EkkU6ODTii6TepDDyHsUmHHsuIxGmdrjAwHcV+fPg8Bbvu6szedZ
YJzkN3JepMaYf+ToC3zTttpQV1uYZGriH1AElhqmZtiRLtueigPcjkvD4mnd69dzhPW7Yc2itg8a
Fcl4veBRvz4o8V5D3SckEm1DdPWQme5QTbkfXJ58yGDPWp5/C4gCh0r8TGVXg3bhz71hVE8z/kSc
YgV0Gm8PRRyuThqYmkTx/qNOfDLGNxE+afz3Df/4pdyfk7M2C+91TK/r3JkCYll/xuvCZogyowuf
6nmKSRy4p0T18b4gsCbgsmRfU0LAhsj3PNnX52DTDJy7VWQ4aPUSx3xtIUSY4sh6s1G6p3azeHeA
vtaNhp7DZXqEdZLhSY1lVPQ6bI3k3yKabOjqKq0OjKUD62lA8TSq+ytk/ktqs4yDP3AKOkb/gxRf
PoVmhafJe3ndGcrifI5aJd0encPH/o09SgLrLfLo2O5jOCFXc4epUBJPb4gYb0Cy41Tz9e53owpu
C7kmkr013KNN/5MKVTAFYJz255208j3wNMNUijMTTq70lk7Bj+5aJwxiGWdQM4yeHccXOVW3K1zV
TrLkPB6JKrE3DdG3EdsSbjVsgk3ZgZotFZyQYcJsuAbwDEZBoSnCEJ95x5luFhqMZxZFgQ94Ffto
MiiOmEswIFwdrju4ChD4/4KByxoWNzgBGd+3IVeR42G2jvtT+67QhG9lxlvLdFyOTRaCHqVsS0BJ
kFtT+2lTuMBxDolIDxeFBRDigY2hd2erRv8AFTu1/ZG9Uq4Ty6Wj8tZuJzRr8L49QWlPX+qvcic9
LUYjOxLMYqP57/OOxusag5AdIdn6ejms+uwtH4AqjSs3F4OyzAuhyhDpDui8YMIDnMVF4tNnul7I
ImRc0WteJ0QkTxZpDGrXeAxZB54mf+3tqZKGrlFn8zmjBSHqnog1aoWfsKKd0hfzakQUHMrws63w
AxT6Xdj8wAthZuDpNnLVn2QOXQdYnkLT+0AMpuMpiNdigNndQs8YYp50JtJMJhiPkN3Ca3tV5fAW
ge8552gdA5utxXbXVrxQkrlT/UPpzvshVSJsDWZZEiBW4+OowC1pvIPQt9Nqqu0gurJtyse+oggW
vZZj+VTFXgg1etXrij5Z6cFJeHr4KR+OtUXeX2/Z2Re8aT79gD/E3w3dNCzqKBPv6L9VPMgEbwtN
3iNYhg7p5rO1ShYZ3JIaC5NrJiwoEWYVAaRL2AmhydToCGtafZYSKBVbkypzcT/L3LdsZJO0/IF9
PY7XJ+ZQlvIgYAM4xJPSGAb0QHQONyouRcVAY4vaSnaDBPyyM/vjkoZgDPyNeMk27C68QCwW0hVq
DAfHkRqaxwAUYLXY5YqwWf1NZz54Ew/1IIXWmC92PhFKxJMKR0yP8I5aaK/4Ri8VG4bBkPsGVr86
Vz7Mecil24ZGhTbKca1fQfvqS8aaAQOu/ZdNWrONK4oqzyhkNd1pLuVtOn0ABIaZgJGYREAjEoKh
XqTKbveJZDjDCUEmjo4eSaGw+Qced20gVkffPx1Z/NxWxsCWeRTCKSrFloFcxEsd85R6DtDvMZ5O
Vr9IAxSyfvzDhp3hh8Wap7vIl3Mp8ABKLJF0B8HLjvRMyoJKuRc9NSSAYfX/X+hXm/cYzHOEKNrt
9XvnempDrRB0ijETskG5w2Qg+Y3/pxod3FKuxKpCztfNpPrGLApFhWN8aoHsSXghcoSYogHwUQss
pU7NIjeSFK79YwlVKI3uLwxN43l4Ge+6T79t9jmDqyZL3cNLZj5zcVfjL49vQ+P/eUuIUsslUS11
ZE4fquvZgmpj0OCQhM04LiupBqvyzXfW53w3p1h/qcwlRRewPpHenn6KA3yz6gXcXQGPpNHStvyG
DAMceBvk7QIf8YbOhBRWiRb5ea0dGIyE/ADbKDG+dmYdd+lTMCbZLmYCAHYWgjUZ5Udo8y7S0b/R
66cILjsYzsjnev0as5kn/RzoO2Z11tR8Bl7HiBxu3G3P+rsb5fOmWEQWY7lxUfrIHG29HHrXW0fu
jgtn3pEp5vmgT6+eNuOlAY6y7IR4AaG2CNdVuLyl1NEu3Ud/Vprz7m1VZ1Ej3MozG86Sg45pNQ9R
lnrFMhp0k8K1AgJ+dzAKgnWCIpBbLtLYM3IGAqX6z6Lo4ZzKf/r+Zkt+F7OIAWijTOUdMJ5401So
7FT+cc46/MJMKQpdpCUQfkYAOXx047JJ0orTxR/r3Rvgu36UlhnlilAMIuDrpADdKLTA51zLxAQO
2L0hsLu0qn298cIRFZO+SAE3F7w2JcgsAwXcztZYghkFFRiryEdp5GLAum4u59cEfmURgPIl80B4
8bdAHcJBAGeWvNv0n8aYuXSoQvTs3r6f3y0WIuIXzpPBvmwh+TOt4hAGe1XkT7LzGzseb3A6AOxi
6Yme9vcv1xPFSedxWa2PtRuAWQHN59e3sHAsEYoc4lt1OqN8tlA0yzpARSD3wlLxU6xzLFvzG/Fl
2nc5tfBNq/ZZ4hjGznQQCNDu0RqMG5JQmWyZofGIWov6uMkEioajAxGx5Kb0IA5hR3UGEicfhwFy
WeJQ3ntEtbB74BCn8IktRUkIv0qnLZSwDh8PTRX3jUaFdQjgofQt8Tht7dZRM7Lw9uKHxvgOvRd/
tHHuwm86ZUZpFJYz9Jtj2VkUojOimxENw0TDhIySk7gRSJMfcEdw75V7PpZ5tiskyt7zhQGdqGJ9
UxEqvGQHiRBHFg0VWzkKI7nGBmAiOC9fkkFdUq3wrpWq5/43HNIbNHFCuwEcjWTjBZ667OGEANvU
toObKuVWQeSDwMSJVEzwyqbObwCg25sJE5h3EgUDfNvbcv09NDSjZB3+JLN0+2pe1AoF9zDznws3
SqDEq6fTqQQc24vUvgRkVaHZeFp5jTwlC6VW+Tyb3k79cyjBDFbI5gp1UBr6paWIT6jTMuLVRy6M
wHWDa2pH5IcKAuWaO4iBwm7Wr8wXu2ukwdnfuUXTiU0vWWyrLuyPgukqApiFEV5HF94boXak9nnE
BuahFbuL58uyZthEpteZcXYfDi4DJpvnFs4M6MmniId0oS2O98bN6bU7eGmtvFJsFAa2TomXwdc/
AkgPqFsABCMTRI86i6CHTUt3yRZznpWjRBJiu/p/wNExilyP1GWLqtLOXz+JuT8yk7bcNSJVwakw
WNThw4Ko6kO2BrPvahtAnZ4DjHebKxuMR8c5NyqFSosyQ5zaouDh7NGZ8YYn1f6N2lcm8np0HUYb
tOaov1UhiyOTPg8uPj/j72YKdbEynS3M0310Anw8+CZ2Wn4IddUIpyU0FLvHNa/1AguF7gr6JF4k
Y5sgHWsuwxvTGRaQDgbBkzf6bJCkO30M+sJSljxIs7xeewnh9kZ8io3eSrGk0M9MjCK6OAfja+9n
hAqFop1sh82qCAjb9d489n1c5j2akaYFEQfGLOJyA+DsacT16GVgu4TsM50g3o7rrLHTMvkREjQV
Y1QdxMx4mOhicTc9oPmzdwX2pZhu7x9qYLhudE54bwyMVT3FllyYiIaaUuvxXDoKnVcLi535wdy5
GDPS8We00WjfvII1yN+6dVZpLJbpexzJbPpsiGg4Fllk+ST36KLCCnKOVrAOuuihPC3Qb+iM3FsS
Buzw+KVEFJZzOW5nEBL7N7OT54JcGKKJuLtr7T1J4h3d9CGLq54iSe8Is/HC/Z3HJENaXBYqn6Lm
NfekhNBQCAMNR/PDP9CS7KS6infeZToshkFWrbERjwyM8G3maa5VSKLm4oVukhfrV8uX/79EdNCH
hXmMbXes5DDnI28dHCxzw9/8rWUqgTO6/QJu0NxqC03MGaib1Kn0XjsHyFZ76JlaTzbGW/YpYqZe
u+HduekwzpnW73Pm2OMjwW2aacKJERI9eYvNBXNwI7EDqCq8ooMIZeAvGC1ZcJaLHp6TLaB8cPXt
2f6ZiVKxjqO7KIEC4DaWmBPXj67eeJLRJAn3biBbIc0whbr2ZH4uOOV4+dqw9UYXYz9G99UAwz9K
130dJu3F0l/gvkMwilrwctC7+BS6I04HqQA2B001Cf/iCUO98Wv0QHybID+77y0HN4i8a1Sw28PG
ztsKXJ1aGHrF2EMg+81BvTdo5YwiErB5OPbHQUA2zwNJinu78YwvYutPGmWePvZlBp4TQQg9aL3W
BOFsc0K9UjYixYT5f3jvqpVwD1VkTNLcLB5tKcT5i0teJ5nlyGstHli65j4O3vVTEdPFmwQx6VTk
JMidRW24HOUlUQoKzQVelYywaSItdWu/CHFGn+M5Tz398hKOAUw7CHFgcK/3HKA09VmwewDn6JkW
S0F+I7UEDUrZp9gZxgbEe8Hj2ZHGzfL/mQMNTwrS1Y5ybFvN3yFya6jJ1QBvALAn84j3kTEZoXoZ
j+ceNIVLL6gEzmX1LxBpEBPiiL+xpmHsKCplGZgczKsnaxa14HJhiYxbf24qKgAv/wQ+iBDd3R1Z
SUO9KVfrWs1nh8HVBmIwqvDUlCnM21+CPl06JByt+9ueNFvAnNyhof1iHRWCt2hwm4L/sori8r77
srE7/tJ1vtzvJQre8wt3MPFbOI8VQxhhGD0rtXhZoSuKynA7X1rKxxdjKQzDX2Gwf0wjA8ORW0JK
M3uscvH912nLmCvHD+Ba/fjJoB1xV9nTo47zUPdR6SvI9UXYjRyFrmEvx2A/MgVgHcQ45GrJxlAY
8G8Di+irCCDbtfX7s8TQBXpaO1KiS6u4+stddr6rp5SKc0qHvaQ2f5UXtFsbFtHQa+mLUMcKY2ZD
WHeQhnF+GcaAj/rLoXO8YlL8j6Lv/+YOz1Y0B3l2kZeLGp00RsVE+DtaJSGskIH56LbLwnSOmrzU
Sw5PcPPefDrFGFUTGOfqYg5+GeSvsBvGSD27N8yuxQFMeXNbTyRy3EeSVbDD3IXJkfPq1lHpBX5m
romyXK/rbu873tvVp0++f6yw2rjeOL1CfeNWouwZoD7Umw1c8Yd2fZbEBf1jD9kwZr4bJ/TT42G1
FQNjhaZ+7fEpALt9s/zY9pbk2599xo/yM00fef1vXBRs8MwyAAVDRt+SQFviChCHbst4MZ/6Cp3m
K6lQ6TRUxq9Oy8WxXYdDXfEGjCqDxOatmavtpZveFwep8qKSErl5jQzoP1EkPUkmj1cVfssXl34x
y9MHsubHv7/+aohjeHYuK3AMO+DHDdaRMxTppQCqoMNC4Pvna1+btRxyhqWyrJRYlJQTVejh57II
/47U5C5jiYO/DdyjFfmDILXeD/gbwP3o2BJKw2f3j7S9GblK/NNwQt1l0pQ3g1XxxOJumBDeeoCo
CgiJJrLgMC3QCxXjXNfy+OqWSURMFNuHKt1+ea2GtbdoPbMnkShFX1ltAzYnueQ8/KLVCsfFse++
xrFDRm1lBXiwx1nAPQOwu4eXWmMI0GqI/JoqbmKs87TAYL7HCUHPgqlV1BBL3aXxgdMY+DOQOZjI
33rs2MVmXJ7kBMIB7LFTNGECliePzijzl+MaYDbfmMp6WbnWYjTsroFl9VaMN+zEe/all/9Tk51k
iSDwuyrpR1SkOTRemeXpMJN9gleHi6QrwWKaQqnVYubtyd1adQvbXRLINJU6N4ZStq5BgLYoNDv5
t3L1lpKqYcSzKa4uAG6IhS92+J+iZJEOXKh7ojSVQ9DVTrzRaMt28A9ks+Afel1uBaNVxIfel469
AQomXHNR4GwjMCZYIiZdZYegIu1vXTNfKJkdA0zy4jSviZTg0D1Hr42G5qQFpSwbJt6JU/NKD9uN
3nw4c89+IEex8tqvh6LaYsh+j0jizF3yw7BXVtXAYBep7nNB0kz680Ok9lDWmBdVs/cAE/RRI+mG
WPOn9rteAdtFVMnAwc1eCsaspBHRIkAUZYh8h+7EFvSu6tR5SMXnOn2rAdSy07uTDmaFAUyTlawW
pFpKrxRg5W0wP0dZi7j10HecGRCIOZlPF5ZpF2u4q4ioJsXJJvBh6Mx/JKrIzhJJaaSTftmNrthT
o8L5utIRmrDr5cZfd5aDJj5Oqz93cWGyZ6kBI8B2mnvQDGgBi4D+DwDpxsYN+MmbBz3CGoUONdJY
PnZsbBzq9Ktwc86WAtvkLISACjSxjiFz6iCkZBelI0GNSYxQFqrpPtgUIrdethuSm5Lzs+aeRLp4
WCS+nh+Cs2mJLwTQtDMW11qs+PV/DJ11lU/FGsJO0/3B0GpUNJ7W1nWzF1DO0fV9kedtusll9KVB
Ahw1r+lMaPa2ahTOUW34MGqY+GNTljJTVZBg818acSeqXGlGGDUezLeUlXIoBcHCVYpSISWBehlm
9hkm9g8TaeUzrJ/3YHRH6YgDXmtlShKfwtiAA9g2frXHWAIKUzM4hhm3SDnFz+rZ0lSISs4kQp6Q
2pDUexfcdVY6ntZ00VcWLLRp3hkcuGgXTjye8+jHiHLbvn7cywfRH1Z0Ai36vjaVUv7EgEZDrbS3
eS8KYBomBJPOvs4PICEX0FhRjt1SKOEFWevCQ98ea5aiSVWpazNv0/e7CezbLhL6mQcyK/CY3aRb
nOMl477UBVNQlLQNFFst2fWdKv7C883y3XHiFpiKRHN/zxHRUEiOmulR4OnygKpCZGPpqhM34kDs
yWt5vKKs2QB/dE9p3iAcTYPzHzkVStHATmLChu7dNJQux4cZ5TEZ8TrAbqqxXUvSEl3V0FbTmPZ/
MGkgRrLsEYGARNTokFktZYIAltwB52bP9wdeiJfM8iVjQFpqeutxS2gImsf1lVhhCxRT0cNqaJWj
pT+XA2imtNmi3V9LxuYsswf/5hVoRT6Rl0UniX0HMWdLkweogLZTxCv3oxQNQkWzZ+MvcVgNCsot
twZ25au3SxicAibIjslrDyv7/7dNTFCZcqeF04PPbeb2ACgI/ZKs9pIWXuv2yGMI42EkzGc/AuaI
AeasNbi90El03b0ygjvuNaj0mIECJkxyb+K/wNbrHqIsAZwZlDkKHxOUo5W+eauuBe6NpSAkHgYw
/lQFsr2EvyMRMf3wQiihVp6SGdajA5YzX0XgxZjajf5kXdm2DTK+OYa6ub5+vGaG38NJ1vvB4zK0
OASrahOGpK8ch3CrDINjbXaj9VPfU0ukwKf6C5sjVGUY4EIsi0leJBHcTjRRfRPmcbYZoC9VcMrr
ys4nn+orhZohYrwuYo/EE7XVznd3RPB+XSRiZZ7CyCEHu0Je+Xb6akiinGeFF8O7lgQZSqIdjnzk
BSOv87ZFkCMqpoX+jCZI6e8Xs5aEO9WivfIAUOyWZVe0WEkcL+m7oPVkq0nkBJZWHO9HSHFVWM2i
NNS1txLVhwwewa8tvNjCMmYalpzZvuJXi5vGNLrwgHu1EOwNgKsqIssr3EDAL2uGo6W3zRoh0Vy7
1IABUPgAj9S1BXceYfR+j5WEti1OXoh2xbW1oPtoUZZ8zO5usHKbhzG7oO4CoFhrAbMaPkrz3Zad
mLUA++EZXyyX5J2nPHt0qFTh7q4M1QrGYIWp2vBblvobzIkCIHnE3Q8C+yLI83NhiI65/Gy5oDmH
StNLRAm0oAptJXAndljfpvN2Z4nWEDj7UXJpKNoWeva2GoHhphmPuxsXiBQi3yL9ZbPAGw8kQheo
w88EXf2dRfs9w0L8bbwigWz1OpefoMxOK8gn+FQDvfAXBafLBBno/jj1DjyZEAn68v4649aCuMJN
2dkGC4cDN1PNbWURIiEkScyoKBb24JwuKkpYd6od9YyliOYgSTgDefUPQbMmb0PvA/jZQiVYgn9n
n+dLDy74iSHe8Cu+R0lxQYCch7ThLmbsySLLTsXYIrQnKmZQV2rfvHdMYlujMHUw51EoZNr4TiEd
iDfz6pQdit42ZP6QWw1Fshj+3YTUoohWHhVrZA0Ru54YPe4zI3wZZQ8zAqhJ3A6+WI09gwVE0CNM
uAsZ5WnGOQblIKo5KT0cOjpqmGe5MEcwZ4M/eJUnvh7ij7pZFbCu7vNZ9T2ovghY7qcv/rkUbtxK
eCx2VdxsylDPOgolMurADK5OgY+mnNJgCJxg6i9EnkGIEHrFfK0kIyLOWm3tpflCw8ajpeK4OaYO
s1sS0RcvuOjqjKp9IAtazWzIhJoKMv/6e6jevdqh25u9QMcI0Slqn3ycQXF/kmNebbqry3U6YyJt
rYJgZiOKi/1nKDnV18rt0gN3BdBK9/F0FU2YTxzRN/ZhbCYvX66SqAN5M4IlJfJj/j/fKnqp5HQP
qn56U/8kSwjnszlbmrOy/k/VS0OBeHc3pQV019N01sBNW7fi5/NFim9WaU8b+UmkxbfHXVbI/52m
n1bO3219jhN+oBBRE5IRykAZNscMSN3sl7sc5ZQZKwpzSGs8jXftowgG+p8jUFzberq/mVexelhX
QHf4GycMZag0k4qT+Usw/jLg4g/4WwllA9Ve9gQqYmzHCfC/EEdplYxNg0TkQxBrfjC2TnhRCZ9q
ZECZURe+igG8W7PEq86nRe+vtvWgWnPpgaDXdLz5hGUU6MFNFXINXrilt1ZurInYTCteE0es6GgX
CdM+Ag9B8Q+vK0nRKKEDV0GzMv2s1Y9gyPUZLTM4fkVCwND17Yn1/l7atdfD59D9bTrY5sskAVPV
1DVPhe60zngqqIaS+2g281r8L5yW3pciNh20Fr4QzZstCpfp4OyDaZuBGwnSAFKdvTsx3ORbSBV5
gq7r6HxNh//5pAR8b+GycUDWrbnNnOTzHsTtU75c4oa0AUlPcavUExKKj/ufkNqPFqNsGcIkQdMG
FNZYUSjCTWAcOJZ9wa7K45Z4cXvYxvero5MP1r8p0MI9LqHsWDeXexiFq1PyYnQKKYfFqmEDzO42
sCdBZ+Vz4knSMbonfiFsGQ6FyxzS/B2xioWxf7Pjy0CW/c6p3Z5WicglLBbnSkGMXUDtZ53mS+Or
HIOnqx6iRRComChv3zmbbT50E4eh9l+uJ6ELmq13erWsPbRtiKFEu5cT+Q9+FLVoybJImyrsxqh7
n3g+qs6EyfOkRYIRZmFKBn0wgSpRSgDXD9Y8mIytGdJQWbYeik0ZxgQ9aG2KTbel43HFTKVQKwAX
A6nwErWAm1/VYEinIwkmPeYaO0GubZFbudx0mYj+OqjhZks1inH6tYCXBExZabHG4Nj5D776SYkv
QkpEkSPxDzUN6PoDbMatUs05sw+S1eHqEkwDN3rJiatRFJuLeE5dMuQdovtLjLNefh7D1h3gza8v
Alb+YH2Ag5wH9SIJa0OcBAL5FIFLy/u935qQfy0xgUcBkcD29JRVAnIJY+80c51QYEjYQCA+mV4k
e3ex+UqpMVc7eTdFClyYa95cA1NI6FLeN719ujkrsO26Zi/cGC+rG6oHQGBMWs2VNs/Bi1KESSKn
h0hsQwkUDrcNdzg7dLnvyN2Dfd1KCUERZ+r4b9KjGV4QTva/BIWBTC3COetDxxCpKa/K6syhQCvK
dm7ImoQnKxw7oN9V04pKBiXnu3tYQ5+ISSMlx3JYFQasN/2x/uPCLID2z9QzxlvjE4dU190z0/9F
WmdTsL8sX2hAvS8y6Un1e+Ez5UEHCZzY2YV5yFU04qfQoNWdq/mtxwIKVsN5POYNyMXU/Lpb8ai7
0u/7WUgmFnEGQaovmwODlU2mLkBsCNEFLeScmEeyLh4mjjtwNHO1zMuKyb/LznLZxA089h4d/GTh
tf7bcyJcAwXbhPvSAIEi60hv7y7wRSkOUgCoBXmqSmyVqF+0DoXPEnvDiSU4XOnmfmRn0t3cbgSB
L0RUJQrD593G1efz1Toirnq/YJIVTrgJs4Bb+8pqXc9JC6iR7faA5Ycr8p3kXYbAxZe1chKtlIuT
ya8fBvE7oDQ+5F1qMnCnzVuZIJzhxuZcS2l0SlQY5KivlWjBHleUPerJT4J4tcTZgw6KZeZxCXri
NgDUkFpViYw7kdEf4lZYkQsWFK37ozqxF4ief3lu6DkdiJL6I6VYIJAgr66d9pvpRH/rn15iPfIc
MdHlO5p9SRxKFMHQaFUEa14lIGna7X0RkU7Dco8YUkgVUmXVKF83ixJtd7FXMrgIK6TBFHlILvUq
6s4qGT1CkOkKLZ1meYXU72vFB8ut5rmVo+8HgCznMQJeFjWeZRernSdhxWXN37PFhjHoQKba+sMk
HRxbHiB/Ypg15fSfOawI7cM3cFXuvlWPPC3Wh0xypDxCFV+aKf12dlJUH/gK0WwjlltqUZnuqyGj
01JudVBsrmqKVFpbxk+OR3e2ujZdi9aR1tXUqCJ+TkRmKth9WRNanrSffelelfiRN6c4vUH4EVJa
hzXNB94c4q4OBW4OXiU3QtigQEMxrvydlzRg1/1b9C6N/xLmYatyN0MSezCsgilhiH3yV34idnQd
ACw5J/WAGmilxutzfrFxaNP+Encat1mLcFB9nwrzyuJKvhrjJg0DtJ4vzLVc0Z3mlDSTzewurinN
PTAoRFSLEog64/uX8IUbRh10F3QV9TZ9hSsIYxzXnzFQflS++cADS3s7T8f+9IKRrh+a/eoCzVOq
7p3LkDYgur2mCy2TAohomAPM5esGhdfEZj2CFbuFFt9ftg+hPnqM01pEyxOSgkDCCaDulXwJSDeg
Q566jyI2CqtobG58nXY4yTmNrB86NPMDLKyAEpE2XSQIJokb2YzRT4P+xYT1nooK9Ftq2nFGk2kp
fVLNBnNVCLgBVZraolwI8K+DcqAHifdWpBormKBrSVcp85hw0JKilDyusoaTYgoMnjHB38Db/ksF
YA2ALqRhgY8cIaTYkCDtgKVUbmHdBC03HdDpUHJBE5n6D8LFU++ItBH4uFWqQMYrBHUbTruUV/36
kaVgm4Ers6zvo2ZoZ0pajYcWox9TPZE7fchOEBm6kJwXRzBae9VVzE71KdsO07X5GpAu4IWgpv5Q
MfMIUuzW72COO0RbfBI6UeRg9+07BIB08v270pT08itRAFggc6WGSOlZ3CGZFAq1VLljTho+wXP0
TuQzCtSmM2RBxmJBLnZBV0+DyfPWdCoB08b14ur6+i+OuyuMsAryc/xWVVO0lVA9utkj1Oz9PtMw
m1S/jW/9ihn+R55rCFrbfwxZlhTG306xdPFQ0wrRqznYs4HSELHN/A5O8pRK+Y0HQ7LXyDuLCE9B
VnbGIZm7TuP/7v6MGGTfxaY/OXKXdtKV9lgN43sdY33uVHnK02fS1ijbVQvi9jWDbEMXMFS9xur6
MWCUIIV0o+P4M62fjtbbVj3FuM+fs39M89TBZdNjUkCj+50AUPQV5Shb/UAT85VVWv2HcpdP1UTE
5wCH3pzKJIhm5CRCVGh9/kKnGG5286MhLCqMWOjJzFkeHxuAWwokbxYSAndJRZ/HFsznG5FZeyft
fiLyYDHQn90ggBeL/Rd0HnI48VU6WHT+TqxTMmk09IlurNEuSDDkKy5BjeVei6uRTCwGeqvrkqiO
JL5S/MEO9lU1StbgSpAxnNLjkcwBuFTbdZNmyW+5zKC132ROWvEu9gs4IGBrpzt/QMrIbUPBYGd9
NV7XnDr/cIXpPiRkteyrI7qEvddJp0gOHtY68oi9okODtHoXL1nvypfkmtjktu8F6rpX4gzZsOQ7
6JrFmaAXsOcQ4aXMjR+uORnwrXkw5ToZpZPO2Yv6lL/eZiRGjxMd2YxYpHW0/T5KLFIPO1frtqsB
WWZlZRHWApKxWKSIYH5klwMNKsjSm/+7JgFY1lGfvGLxaKtW3r1/DeRQvY9vwFvuBUEMHkoKWwiM
JdZ9YiFlkuHWWz3eXsK509saUuWOhUCS9QlI0P4SIBRd492ZdQ6cpcK3EBRZYge5rF3NeWYcKLf0
OcSOOaJXIB/8tqwqnWDKYEIk1NZ3EEm95+xzcCpITXFIkkH3MEfmmVtMiR/H1cBGFQ4218wLbVBO
oj5cMtNah0dCn2qZtn85lqi05uu5EIiSQLPOstowalUZpfTNQUhO0kr3URvPT3Tbc8/gfBa3n+Ks
T7oVeRzoGA8HZd8FSRL6K1aAIYL3AG7wY7mdbaQg20yj71pHTcNDpknRlCi5rYRGQStpD8GS5m3h
EEWOSoSZDsfBW4bZMpJ0jzo9FFZGv48oVOC1XKCmEGua/gDm6B5ivA6+mD7VjiITxqBeOaxnAtsd
r5xWf+QcLGku1HY6evvP/tpKjSM8UWbQQ/0xmMTQxt/92sJco6Y8jXm/qzs6B0+JS3UhBqTKMJUA
cILk6yCX/w848aIyVCztqE4wWStK8/lO3HLHvmgdihB65tEfauXm4IuBgmlo8mrexTd4fps6QGkH
xgR27To4PE1IlTL0R6mC/Vu85h5AhNwqi7a6kDmZnCKq8P7cNK/sEmpeRukub+zk3mboEU91//aI
0dUd/gM4zOFF7/rqRqj25F8KRk9Gxy2sM68IT3PTkJTHMAdq1PS4xYv4NBXp/CZ2X0PmDd+rW3pI
JUnTQLyeFKekDPlEM0f0SzvU+281W91WVjayuqXvV7Ac6gJ3whmBZfypH4EGz7f5MaJLF0oJu9G1
Cy58Ci70Ellp2tR+x9X7GKhl7GtUQ5g2mLh8FGKEcKXHP9JFFusz0ZpRHfw6YXsw/htUb+gsBPfd
G7E8MYzrpNMazDpOBJbZ0FUT+HlkM688T9Xt3lkOdAKgq1F6UBbT6Bt+oYMo/QKXq2JM/UoKzsSB
mlEOiQv99+r3K2L0ekHbua3N2coxeYrwwIRiJOkg775qJJQ9m0g9i4jwpXAFbBrvsNHPihVQcMaH
XEq6XVbfAFAS3fEhmxKsezrDfrXXuwCnfwvLElDIpKX0FP1Mh0Pi+EW212kP44ZjIf7HLdQPbAOf
28yIABs7Mx0SJ69+zvSLvzLpHSab9of/MZ7xylICQuAhPdczjmzXJxvzcG5DT7fFHtmwr5+nQNzV
qa1/ju1WlkHkvL0udnn/enJnjMKs1B1CXr6XpQdOL/x2y/wHaxQc8PrW70jOF6VwELON4TQfBLe4
1Aaz3Df0Ylw9uJb6p6m6PSLqQbEPTEyQTEBQ4QBRvg3VC74EfJkjxf6mNbXF8h7MUT7J6hCGCqak
Jfldr3s1xd7ey/Loq3BQXFt6bCQcut0a1Oqao0mLZUd/ScnSsXQ3fCjkpSMjY050yAtlwgTUN1Kq
LBFjI1+HYavry7q4StaP7UnKWlwoW6uRkfStV8w1PkJIOdl+BffGQ3E9waZwr3hZQke4rLfcrP6j
5ecfHcSdm2mS6Fc7qOgN2xdsZbz6V1hjShxXmyURXDLn11mi+bNxjS/pm047XbhuLOOacN6U9Qc2
KxX0FYrU6zlJXOGwDi25gcdVoWzx6RngIuDV92WWMgEw4uKnGKWD5PtLSATPDk74t+mGRjSgM3kb
cv7F7pYMhMbgx/NrcPyiEUU7hBgOE0VVnUOZu2Kfk3rhGs+LpPOVFRWXjnpvHwQaRUtAji8NsNW6
VV0Lrd6uHSSK4vJvGCZ884qgu080aFF70Tflxt3DmHlzNbNGEpRpBjTdOPryDWqeMG4F1BDTnIDN
wUW7XQkOu7swy1M6iHb7LDyaNrH7nUqvxMgatT3AJwmnOiC/tocNACl6u71x6yiROdwf9J3JMqgB
pHtXN64x/s2fmUpcvWpOgeulfpqctoBfGo6oiKQblTHDTwX7xSWQ1N1U1QVqz9EarYpT3SEKBJbX
POfHY7WYMYn6q0R7+k4XsbVQP7lpMPktnk6AddXO4Z+Ey4AMS6uyEjmHq9cveQf5/vVRlGJYEfWv
Fgd0JSJvXWhJYGWbU4EqxCHKqv3gbCrPb0ovkJH0LoRy5etMltK3rmT5X9GLb8cjaL5dwxq45Cbq
30TG7yb1lXonoIz7fcewHNLeOmGNDiSWR9trH/jifNUwkPO4WMdzqTrc0DjMo8YHx2hv6oPzqrvY
lsNBT4TQKNm4TTKXkATYYcvBP7cBKYwE/bypnelToFBPTT2t7mLl+GyrbpniBAyXTmuZ8lCUG5K8
UgeTUhSyaECNAMC422BjbCze8LUbbL04HShgtPJElSJpROo8Zu+0NGAycKaq2615S7c5L6Nhu50a
VrLEuLx51odUgmTC89ZOen5uw/zLZYUH5LSLZzQWQyqFk3rddKxuKeti3i+lEUKhJDtVhga0t+Uf
5uY2MIuzcDsQHuRw0d2knlz73lw4CQN/HWaWIxXxVtA2ip1EypDxgMOfo2atzaszjArhNlefMCQk
wOgb4HrbAD1Zy5W08e17dvFs6KFMxob2Nt3B1Q3diI4U8xKllzQmLanwqNPMveNc3JR2J9RJuY2I
IRFhX+zVwhUVWI2zr4aV4kPG2uzqch52v41xu74lA0cmJfryAbmU48sMCxjtYsg6lJQwTk40gA9w
+8kX3YpmsbEuPNb/jHdnJ76w4LCc8UFp2hCvNNMaWrwyNd6C563zwWEA5X667AG57zDdbkrDN01+
FzFx0ghQIoUQzObWONRWhuWzCZuP4GAJFh6sWlX5cEQLJdjohIsTMBpvc2Fidru5LU4qo2FLy1lT
ocBHp3zbG83nPCzt9bcQmQ3HIDgYoajwURJaBgDm9eKMNbQTIFFSRWQ0IF87FXs7daMxEb/Sbb2c
nHNP0+YW2s/HRkfLIKhcf0ixkCUwkqgP4q2+M4J/odWKnMy3WMGYlQvE6Em37OcPnBiKYcE7ej1x
kbty04+XJwAD6gQ8Zf7vfBcVW2uFCfGjJ44q5NgHhxrxP4abk2PzwOoQLvZcQeMu71VW4YWcNzcY
5UiA+gG7a2aWNxjX0cKJqXfz0ty0z3hbZMnIy9xB+M0pem6DIy66Wqnkse5IDyKOp92TXs/ngJuP
vD/X2nuVtxYDtbhDZ1W+yZ6iBl5COkkdSmsZvzgToRkbvlTeQHuuZrrIOxEecRD6lXJrOygdDv9R
p8+7pMM8xbn/3zWK9HTYfOt/HajhWG2hfoOp7Oa/f6PUVklOdQtPvc0ZwS3lVRP7wDMeeGLZR46H
idObQKhv4epB5rdnGs9eKLmlU2Yk5XMcL0b8Y/z35xZJn5NOUo6q6mbvPorwM0TxBRkgr3lXj1Vv
Cngg7nauLcMUWT03bS+U0BfqqSXMyQKcKtc/qTL4C4v4muCPZH7yHFfueHs5Lxuozwkf7BoZaNoj
F2liVNvwfCRou2aS4OgqmWuspUcwbhvtHZoZS2u5Lk3XgqhU0Df7Wj6Qc0zsgCQbs+rOQ7aq4woq
wh3AT8jf01fmFYaY+KEFyv8IneQj4uRE81h14QSknwcNRgtUa4aZDaQWFYfJBzHSGswtxuNUDNxG
3nX/LaTFDXSF0gPZV7+0qcqHqBkDW9aLiyWbinmcnM5p/NufsLx3HXKhVxWcVUNGlWtx5uRjSxjl
fox8I1sZMA0F9oVAyDiSiZ+Oz19f+G7UXdlrrNkKHz6cESthxHrLPD/awnD8R1urODjssxito8tp
4NDhW+FCupXhg2F1zQzRCaakLohU5rXSbknSpowtmJectz6CVUAXWejhNqBDZD/zGpT6f/UFZsQQ
6o40KdUGSN8h+d5w+pgTj9UebOSufmqX0X5ePHlxuVNaVQwkTrTPF0Gf11R0SQL0CqA/M2MRAntJ
y2on7xDUi9KNgiVA8UP1RGnfOm/nSzCmhTyFzdXMIni4fLISHas8UbDNMPe0aCFHXEKwL4G4SxQY
i851e/s/RGCS//lPsS73bapzolXtKVf65IAHOEjDK/yU2DpCmwAP0g8bvCXlxHjkH7so3nE1UcOF
ly7InYiEqrdgqYhKNyhAfT3d+kCRX0wCcD2A8JR6LoXrLQuGIa69PtuJd0S5xeT4d92HP0gkgetN
m69bRbQc5HD30TPG/bTvg0W6l7pp1sCPslTJaNPtDtJE3qDvxSKKwhR7vEkMN4PSXyrWZNQywHri
f2i8a2VuPrTCG6H7e2NSlxJl+VKlHB4naiaJDISGe4KdVlfrYwwUO57/LQxaHiLqQroma9kLuLqB
UzXIcgoV0J4a13NtIFME+UQGQyFwPJk/BN3AZDLt8q4XPkVZAxwxDeRp/r6OLfA5eSJrh6whjxFo
mZ7ddzFrYvp22cGKo66P+u9yauqlze6/Ls8zvXlMDx2cQcedbb5hq7g/fDbgzzHYCHgNP+ktmPiQ
yIWXhwYwr3vehq70u8e9qmKBsfrwtfbotG3TcSduv3QqtdJAaBRWrxfGRwOMB4Cq6GwWVoSzxvHN
97Ddsme8CynCHWAuLn+mTP93/gBYhauR5hlCg8SofFRySQxC+JbaQaYUoDbMnZ4u1q+BKYFJ21Bo
lyS75zIqJUi4J55lRRwm+SiVgSz9/nRf9zcyYLBUSp0ktQZhbwUkG769BSntATksfqwFITDjBqk0
J7B2ck29txrwOIA6FV10Pfa5HKnu4e+utrhk1DX0u4mtH52yPwuZdX54HCvcaYQ/ytSgzC7qAu8t
22MvRQAnkY7KhsijJTk/GMabjAWwD9z+ACD0lirpFpfnRQSxhn3jhjxnTrswEI/ly9dwTZ158No7
E7Xvk9HKimP6Mogmdom7VArtpE39vRkcfclBm+jDx/bxp38u/htQW9wj0ksbaugg7ExFjMSirFUc
s/Yy0gOEmqv1MQmbKoK50nIsk0tudmsatQCqhyKW5cYLdWkwmwuU2oCmeSBCHHH6gzv8Ww0gUq5n
SMmcjtpbkTZ7+y6SlvKbN///vM9ZIc7dUnooPoYi3cUaG3b05VOv8SazzCWJAibsG30kjmRZd+ot
ooG/+KtkK1z4nx3hqFKITorkXForZ6nBXZJpAVepw6Z0J/LbkC9dUZi2vmpm4TfYKfRI3HtrW4qc
7ZhjRC+pw+wkt+fZDatCX+rlw56ZYkliJ5tdO16XIEu/WrszdfS7gGuZvE9Qw98JS1AUWv4Wjpv7
i2H1PgdvlhUa2cJNnxiJ2fOurg3BpBeEB6gL54BQWe3B0DivVpT0geg8Tjtmq+3+mOvZt8iEhq2L
W8f8L/3QW2AZ8NiWmYUIYfb3OsGN1GQ61AcLQdMjB90ERb4CX6P3mteER8Vgop793xFwLuE+tg7p
VrbowujPwYTvEmZ0aqbN0+p3Zwj24ztlXB0HMS1VVYLRfAjbCaq1232d3fkBvM7AO1xY4WThyP8+
AnsEVFi/CO8eUgmDLj8WWPeHdiy0mtB/h3ZNKR34gBCQoVZI7yuTOJco5ZsT5xfRrKjpgj0B0gB8
Y1+1KFciGH9xXoFkjkDCj8REYPvLXdAjeQbauBT0/SLcaxZ1fnsVWhLEzoBt+MhikOtx6Ej48ypI
lJEynJ85KkR60dKvvZSRZNVqI1L9zR4XTnB9qvkJXxk/ZgEqJlR4oLYoja34tudwxIFGujQqDsNh
tZZ+TfqPjlprvqO8aTOcNGMkuPHsDfvdfbGcbMgoAazugmp8qfxXQWmcRTEtOPbNWGkuUOMXKkMh
VYCmuvDw3KhZudzUbzVeP6W8/JQFlCx1iEhnlAnHZMwiIQpbrkb1cVartGV0OuX/4fVSPcWPyBNc
DyUZIv36dSHbGtP0PoNHvr3aQyJyshKkVlxqFzxKsKFxPT3GFkSdgBwDZ5cmLst9ACn59Zd177nB
MB1+3PjNUvIfyRpDIF3x9J441nBWSiqUklFfMmvfeXdNIYyZrEEGrcMOzvYPi/GmFZdIX2+NudVK
duoHpZVmjL/oJ4mXFh99v6un4en17hz/sSnDh74/4IJCfHp6V7JFGAVaKgMBrrjmGWB7JwCEPRXR
jT8IaWWD7FCXjMYN5AZQhie2aDrFR5wOIMGQ3TCXCpp9K2+K0TVqcmPeLgrHVNFo4Jes4oqqw6lb
WAyAvSF3PVXGxuHbMjiXIAU71gtpb+M5COwl8bynYwB+nfJiLnAxXSowyzsZ/7TEWzF7MKKndqvo
K12xOQo0k3myv3j6cuzphL9I1yb8gZ/AERGRILqNzd9/dsPfoe3++tANidHl9s2umMgU2vhHYS5j
1/PnT2yccHJisDY/dSHiBJsr1EHvP0LTxZwXsz1HHnqPg//6syg9Abvm3PFr9uMJ6nW341FDtG57
kXjax8l72XQR0ka29ou006Hpg0/aVxVRJndXxJWhHACChyM6e8nEwFYaD4XjYLd0SZ7ovOX9rG/Z
wGTngvoOZjKC1taZVYdrTbpGKyrA5eDF5k157tntiAwe0umDXvgmndDjfuPMu+Zbx97DKNr4rg8s
a+BQp2pyezbeosp6nTU17AFWC3FKxP2Tly7WCCmF264ezGW3cW+5o3TMR4QCusME5d4FqG7vSoVk
9DqpCzyzYDwfylHmpL3f64mPr7+5S+hyTZjWk0mUVvKTAlCaarp8xXucyvtS7qaRGJ7Kb/89zkd1
kzyhn26BWyssYwecZ7NaIQOXUofFlKLMg4KL2StUk6iOoNaeqmfikZPKNZXm1dz7f+B2wfy6O+j1
gT8C5CDQQpF9ivcVMqdGB2tugrfP9eGSbV9UQc0Ucz0vfi+c2T++mvBfylomcsoG3+vfVKv98O0J
5Qhq2xw+x0sR8MgEdXJF4T9qJbdGuxIsjrEcUjYip3VUBH7fbKLsUw8Z6X2fiXI20zb305uDDN/A
Y1cnHnpL3L+X5HEOuUPbHYmg4usgs6ryOSRWPGBBxbutiFFbJOMDcpLHxjdJZESumo1nRzRcRkqY
qQUrujnlmOz44mF4k5flJgmLQ67sXgfb8rCB/S0AUPKUBi00qW6O/LyJ3MsM/LSf2JStSuZb6jcd
236m1bOi19LDG6K/y68WErrzUbIkCDektA0xscDiwIDtrO0L4BSkJdB8U3eNTZftEY9+PpZwH0WF
a/r5mZpZ2L2vEvOdXYI4cxP2oFXfmshdEsU70qKdlN2Ro6lZcaZ/OGeJfV/GeebpfYueaO1uqXid
xV/ihD8/TIdS5RZEIJG0bYR2fHXqYAADy9o4AaIVWwFaIZfMNWFGmHCdrSe/1ussDRnhSWTWNO+q
lBP7Fp3UztmYzj86c//2h1ncTtmD/MpjDy8dtSUrAtQB/DvkSHWnx5w4AWo6rkmMtaj/dAxESyB1
i6jJpUEtNudqaqUfcHDO4l/Da2BUJuome6hEjYedmS3WXrA2kup8CecrLJomNyKBXhoRa3GI8DqS
TBTR5FLocIG1doeWajdwmVYFkvFwIKPRmg+UIaKHER1AmjD0c75uCsm8QaiYQ3GMsVs//uhVvp67
4dWl/a3Hxq6Ds1j4tHT743T8IUo4DAgLb89HMNI7RbyI0rVTuBzQbGPFgdR9oXOt3O6flbQd6r1K
IMH6Dc1KdgejbbLmZETevS1u6hccH1leWPRiw/Eyr5Psx84dflzu/LNi8pFAuAw8FNyqdSc5C77a
j7v+vzpIfbGs1CysmqdSUcVUMBKDZdrQFPhJ3i+EUiIXusID0wEhrbV0S1z5nsFHKxoW8bJZ9uop
LsDbjkQmFDElbD3fUw/ZcFLgv/HzzFCdLSJ7PnM0Iu8PYAbwUO4SYLCBhbHdlbxHT9UT7STSWTPR
h7/usDq6jQSA8pwrZw64MNqVHg6SKXtUU04AHTgXORHKZ8zO3yESDS1UswJC4f9NFMvgLt9zUdMb
Usvxcx3sHXRhfBG8WleKzaETJBaCgeYd1FkAVQyl+oWhPHOeTWS2qkxdJzekVEXLz2MLyaPxMpKC
jyiN77sjTey7oFA2kgHVCHv7uU715i4BvvkDTw1pV/L+stk3zYalZ4zfQE9E81p9MeTBMua+nHKj
JsUD48Yd/83uk8oaGmmw/uoUnxfMUe4LGESeoXHGMd/KTXz7hRKcXR/jWZDQj4OlBblaqblnfVW0
LjRTQyImpVcxggI/hsRQS/97vrjcmw9CpZt+yoOq9f//Q8ndIyubeSX1lGAZfb79Hs8If8cecx3q
mz1caZDO312GUkHmPYOr1zPsRKh7U5Xg/0sm600H+ur+ameuxwMzr7nSw14GmqFvbPoMIpbmqr5s
h70qSMX1ANHgMnCrfAMsoT0SSWmbuqmWO43FTmMbayGoIfDw3YBhpjpu6WMLSgYzYf6PRzU8Mheq
T4Ykn6uu+Dos4EaOar4K6gfCm0nSlJxiOIWnpZpwErUIfumqiBZoNwp9rebxoX+bEod3naM8/qEJ
CAi+BPIUsHZT5VX860XV29GvUyHQm/Yu6FGHJCkdkYhfJar5SRzfi/7wyL8Fcxsccrb9H7Cg4zl2
A0IdosWoZlDAl7Q38Ei3HH3dpwnvqjzARbPkhfSfTfHmxEWjeyrPFu5hlQHecG554e2alVTyXG4i
5UJq3PLd9if2BO7C1Dhg2I5NUfbO9JRVfbz8v8Q7Acp2WMFwAVTdOlOUJPXLBQ4eWjarRjQXA5c2
A3ugnIK+Q6DZd+/A1JnJBOEUUZ86dHsXPe/YUVBHz4LlIf5weo1Y6gigtPx/ZS4d+Vc/O8ssBXfU
6qzRKxkO9OJbt8fRUWKnXXenv1Nj9Jlp5Q2gZOUcb1ptltvF5k1h54u04eMC0VFAgRTHNQr/iOCC
M+0I1oAZnVw9AKS3AG4XKwcDDBPPlM2gsc1Qeu0WATI0xDFXx8GVIjYIPzt25PBp19VBLX9fCKnb
hHGLXGJmZMon0tzhDjBpzcP0KwCxaHd+n//XIW95lKVAjwVYRguANKXWPWmXbhzSv9ipH+HThmcf
jhFC826d0upMCQoN1WGK7uX1+TJzCQAsxmtyOAjRJjCvRrNEnsL8s8XSuEJlmmwRLFD9gBC9sV4r
nN9+jR89Uk4SekKhHpG2ANEoQ3eZacqWqfXcykW1PTWnSMDXsrB3IDp1ZfEL9OSvUxu5CrazXI4A
VUZZrP0P/0ffsN8gZQZQ4htsM/WjKrw/Ca+F6IwGWR25mnKh+MP7O45MJoV0alKB83n5I5fStW5q
moWIrsGTOGVT7AjBhnQ4HeQA3xsm22tQei7rOF+UA9TwGof7davzDLBp2TRuwWipBwwpKz4a7uyN
A1fuNGoRrlXEjB4633KljYk26emha0w9cHR3UDyPgEyIEA5zdVk7XBNxxmBPMnnDCBm/BrLjTgUx
UkFbxYgRe9XLUTUHK4zssG/cyYbWdpot4+00qwbJztjAhs5x9X+Zq115b4dhdZDVpT6U5HKrZrmS
AI34hDfaIfMzhQJpZt52EAyf2fsFeSzvDZkgmwgZILXbOHglktWlxHPum31EwWoGyebcQKuzf6/R
IxDZ1SUK6j4pgIpbOTKlnWTCOXYMSTo70K43hH38ar3wLIQXQSmztq9i7dSxD1a0btrr/zjx9q7k
FT3qJHBA6hSfoTWyaxLBE5+wt/CLgwFI/QfU80WblklDBeAwx444hqPE3hNwM5/+BzGTnMS0cB59
9UMjP1OL19fxYS33IHqN00HSeo5lHhu90MlpoHAWSC0qDvOp87sHbd3JIH2gA9ZJqIK8l/KkUti3
14L9Q2vvUEZr7bk4RO4WGnRdqMsYaqd5m1KasWnsw/8wjzCuVHgwKel1Ti6Ol7xsaWyJIqFxeCyS
kya5x51rr4z7XiCAtoWLvVZsudUiqCpun8Y0YUSsFegzrdaA8KTLH0o0JDKCXUGbljuUkcuAs/se
MeLmIA89BSYNz34KR9R4gp6hq8JpCYCxY2V3nMGFz2Nwah8GAhe/jOA6T6YTCtq+fgfaw6FwMxq2
20SebTJfo6Row7euYIbSAgaug6bWeVCTYYdUt1RjlbuPs5sg8rbEtzlJQPLQpt3z9zIukhoFXmUi
yP1xO4qNowg4Op21BPEMxHG9YZIUeM5zvXQzsl+yvIwNd2W+Nn43Xnxk25aw3DuHTvJsyNwPJtdG
yT5Ei3HOLr/JynFC7qPjgnkR1HDzbis/Xp14EUP/QsE0ejZ2RPNVMRd5z/e8/XdQ6LwnTLPIwxdk
E01KUrdvU+2cY1EXwOhasjYCv1uwvczJJk9KlyqC6H306dBhFEGE6S1+UZWfPTw1IRytAGC7Mjki
7TE4T7rFxbaoruyBoUCIcbSvfPmQAXKWnOlbSY9il4aQneQDuEGvUERVBffBHKgDj2mcEKPQsekd
SsYfB58u7QIEdrHWCo7koGJRU3Z6rtppwdnYYfWttMUKpmNXkUptUxjyzZLNHv/PbwnKGtJm/eb7
FBoUlkOyLC/h8j4OhwL+8X6t3QOjBm9ElXhfp3Tmh52Y7PgWUy3OAJItcyh7GHRiu/bcVSydnUzF
/iWtlxcGQf8Nf1BK7pec8zIkNvSIOdQtAY8bbAYXZlyPktmc1FrREiQh90XHsSftiBygBl5wgvaj
n73pGB6lXVzin5ee1GgUkD4mJ7a1X5OArJBimjtCAJrviAnioxTbt24LFitn1HXLHnizv2G3ZQ5/
1D5DeB4Pm/2cnpKP+JfzSSJ2GU+mCtiGV6J5Xm31M0qmHv6BSRiqhrMTzGgcJYm5yuNkK09S2Mfo
dCl4tdWfjX2FxhhX+zkVeahFvPGPPLdIAG2MdTxIZukH/R2h623XIODYtW/GIk2TpXopupNCKI2O
aM5uUOdppGJOTR0zLhhMnYe6aQE/HGWLM0TlLw+5UH2n7oqIEj+a0CwdCLE/wJZniLwOzYdfXwKW
E6HVB1OTVo4mVyxuPSMp/PaWkpYUqVM5ADTR2Fpv9qopuB7fD7JnqjvI+h9Nk3uUjLYT37du3EeC
O+hdC0CdKQzQP5UJJZx6Bkt1BCU8c//JJlXb7YkoZp/11pQb9WwFu6KNhhd6Z43+exXG/CQuc4hw
YOCxuIdBO/fOXvsRydOCcqq1WBDim8Ub6Hc9Fl8sMmryt5WhjiUcoHLAkXnJORCZvluYWBBmJoCr
LuLFbmIfsMysfw/2GSq+wWdXkrVvZHP9dL5tnUUhG0XqqFquyK2+3ruH2l77hBdezgsOsj8DyCOa
7ZqdtkWglAjlWXmkm8gUXdfW17rHl6ChHL4AR+rWAxybPI5NxWXVUWP7mhrhYVnARznMBVq6yi/y
kmWNUO+qrPJIfFbXimRcyiaLo8L7nTL17meJjMKadlLTbyLrC17XpwBf6Vlgej6pZ1lBI1qGE2Gc
JCBhkVhIIfy78XTN4WHm9mYA18UdUNx4Px+jBo0FSxjCwB6MkqTq91C1IvG3kPLfVV9MNnc7v8Fr
hIOlUVqs3pIhc/N2Jap/yqFm7nQEd+WE/QPHy33qSz3snkC+BWEowfIGV/OXp1DoJ8okHMtd62Lb
/h0KO9pKsYyq8DQrT+RFHxcIPQGtbJJCgKMTJPIRI/Sgm2+D2iurcQ3ZS9IA5zoqa2LVPj6ubaji
k5X6geWlG6skxesJR2WDsE6ChQXtalcDaag1x6X9v8+QzfK+BJJCw2wxJ94NiqJsDT1+klX8h4lt
r5xj/j+2LmtlO2SQplETpKKMYrMsxptyi8m+LCH7IiVV0zwASa45l+iggMvn2szfselkl72Wgf+F
OloRqa5jLAc2OgR5QhkCwO6KKDS1Sm2PVIhskbZ1du4eMwY4LaLzU/7UDBD58oOB3oJ8TNSr+z1Y
4XfmXb3GblpX+NRYUqZX7bXiZTVuDPTPdeAHVHPBjU3stkKb5OyoTvhfGkjS/lUnNTXnxz8rJrsY
1lhfsWHuzV97b460qfWoC+W3CufMj8emF0q2olZ4ADXRmmmygNMLkGyMdo4ovWkp0v6+cMN/yK03
Xemt7hfgDj9DP1WeZIx6zRu/bq81ub7nFC5IV2rjz/nrqMHkNB/TxKuH+rexCxftFPFyhVwPhSId
kKNWbYcyPDgDDIFSoO4Gbe0Q8bxvRKmTU+5HC/ggouiYO+msuW+OPbOQjgwyT3mKNQLg7NWgNQTU
i8GJG6SovytgASTYQA5/gjqaJ+WdxdOm+OfkstdDy/d8FchhuhHW00J3Txgjw4SOAyT79hQThrFX
eUeUW4H8oQPXwVHJ5e1B/YAUx5HAjDvtw/Ibf0qA0QZgmmqlDAyXCuKiICc5z3+FX7ct/P6ezZZw
XverWFUqnglEha5Gjl6oyr7jCdZ9BLLwXY/mjNoLOEuErAEB6bz6mCSAMJbF7aXGGKPOqXdcWZX0
XUNCEovp02UshjubjrsJ3eFFyHPSNEzGMYfth50w7rkD+IgnZVAg9Z7/gmyvnrNfK/tymoOa9QKh
Ozt6GGNLae79bCpWjC5M8ICMgzIhDhCwUcNCoMaD8GvMUb/N7saosXNFMcM4QlpWPNi1uSEvYp9y
GAFdoHQr+nRdZidqGzVngbWNYXNmB53fH5ErRhDlXtAweFYrBFFbt+xqH6RcUknYw9HmHLyXoT+d
b9+6vOjqKT+GuGw0oAIO8wr7UMaAwW/YbGZ8ckeRbb8tc+l29uZIFALPxLPwOU0K2IlY7ktUlkiO
glscB0lhENc/8OcpGKCYaPoTuvorOjZdh6E3LTVt4CqciiK4TvmOtTXfBpUlpPpz+VN6JpplxNEf
HOL4j/tRuvQR8zzJ8hLgH3MByCh3GSK80UTt3fBdcoWTJip3Dx7Ue4+FGLK/JGJ+2BAwRwV/CZ3G
ImexGeEcjV4cUmB4Xe9KgAoTIxkOOPNmWryNB5uGRyhEiLmjrFVF7yrzo6DIP8uhLRblxW4Td0B8
dO6Sj7A6e5jEeN7umqh3byVL+gGrMMp1XMdUbSv+4YOVSg5s3Vvmdznjrk3tf08tzv7kPJ+dgG/b
WHpuLfIE0hlknH6IDF1mh4+kNRt5ieNj/VEvupyb5/Axjel50j/mKEIjKbX0XynUXc9qqXq1o2CZ
9buHOZeSK364NE7nSAJQM+NEzwpaYVOsLagg+xx9g+Bdo+0NUiFeCGlCjk6PN2UCoW1Co4TU00+m
BDZ+gSErzSBiZdXgcAhXudvQLNzaDlEy2VboJy1aqvhG9/LsPDk4OwR7peuxiTk0XvYl1HjXqlwK
rPdZc36COy0HDf640xGM6DHP2Zi4OlonmSUr41EVPOrTCfvt9BeEqYdetVodP8c5IC2a6gQDNTRC
QnmyJqAxpCMynN9XYv7fdOFOJf/9CQN2cupdkmWXzyNjAl2iuuIWZaPFycafiakvqu9aXVJpwV0D
KXgXXiKp03fujt0aWrEHpQlYtMLDsDsYyaN41JN2hm3tnUeTkVFnnLX5lDVMgLsaDhzUVTwrSiV5
7Dy1M79LO3n14aARHOkwVVCsukr4OXugxZvQaAoIuVqptOsigqhOtgEbRMGn/RhqzfH05J3LYjVx
oR6Kjmql10RbVgGQMRQrJQkdEmd9TwyVQDmIUzSUVKqacvMh8xyjN74fT/+g6Of7NW9uQv1nr+UG
jwWDI3BidVBhisiepypReDTle2iAH/P62+H3O0iTjVuKiodoehMwH3H1BLn/1i1JKsEX1CXebcrN
XenogZTOm8er2rz5N6pW0Bpq4fweCj1UPHpaWga+ZU1BaKZGzHAZQBp9UQ/IEmpYaRWTnP9ydF8N
BI/JEzVeiqrXWrFTCbkeA2M4GmSdHWs94x4DKY+tunPhzVCj1gKAddi16+csIFodes4GB4d7dbF7
EG1XDgYSmUiKQ+ENSf5tlLxicOgbPdLg+8fdwqaTo0tpQ5LbUcoiLfApgP9Oiz+JDeqxNXblKNFU
QYHlwMPWT+9vdCZ9JnTqg2OUb2oCgm0AZ5VAPPC/zEKVuqC6RJUa6LVNZnYf7TDfcqfd7tw/8fcN
a4Orw41LETR8P2wBLvuBhiq33ODlMSy1M2+4SeGZhKoM/5Goc/lW6/WntwtKwoq8pWyIsskDBcu6
DnXw/upmSI0LmvxWmMZH0qEzf5E9yALoyMFtRe8TI8DaBWvMCdrIkxLd2RBX0bX5e681ndQLrcFw
Qbu0/Hx/LRmARt65R6sXGX38ZN22gEFpGleFxUA55Mo5kNfdVZa6qrw4Mih7Px9V24UQg10KvBnv
rJXxbX2pnZ+dFpyFtqz6V2lu8DrN5mN29FSklajkcKFVtHMU+n9yj90H2XP7p/uPCRSCtQ2aaWIm
jmt3D6DeABULtDfvfYBi/efjmRJNYWb0toIPfaff3DIHbCAJzAxV9Hk9cLo0kd3yheuvGwCSkjza
65aghs5ztU6uoXZDkGjz7T9S1PwIH1glIZPr4T5DKdggyqI55VMYg2Ct7/7g+hVVWKn7W6yYbopE
+zprn2xjLgFqdL1R9zW9PRJt3eeHWfHnbH3MojJ9eMOiqY9LdgJDsDOEAutkc+0LWmWS+PmmPols
i5N9Qn+AVOcOpjTH8tHCSFW0FDZeT4VRL4O4Z4yvw05AWPyWhYMV1+C3JUv0bC8ZfYyYNm0E7tO0
9mVyAa7UrE8CBh19ZN0pwWg17GHx7qC9id8srb+mqlV9t/u3S2pDhC2HtjELDlAWwEFBEizOUgHb
MkZsbTll/1xNoV1jz40C4ZRT/aslxlFIZk05hgZXT/ZjguNOTud8bype+D6/rRLQL6dG7rhcdsch
xo+Udd9d/DM8GpADvYXyFOSMxNRDVch0hO5z66z/6uvfV9iiINJ1GPuTurYNkzOGcBKruuVPgwHm
ArqOi6zcJjcBqDxx6fN4fyYZt5e3zLLrM/bN4CmbFrap+OQkBW7LyeaxO4x7aDBL+FqetYaRBtIC
MllmQyQJTcKKhExfmXQDE9hfC8ZeioaZJ4Co/sgTFs2Gc0L13uIZHE8OjSlqaokXs/fZ9y3Scq3U
geE9TFOboxrURGbq3dDgUOrWihxPae9xB7aijGDZ2iFNcvF6cf6BXxX/XszZafIkAsc6jshJnQva
uE7W9zW72K5rSc1qbw4jxVm0Ibd8+R5zPDtBhIUrccPcF0U7fxJ74N9VUaOXPl1lcUBdGEO+XpHz
kAk3q+P49sxT0hB3rgu3dAaK0v8Rrk5+11UbJfaLVhE3uoQ1q2ZvwNy9Itiq7VWlBqfQxgeqM3uw
b5d0zrem9wzPMGMxMkJ9W8cz1e56OpyQOn3Pr6DbkXEwXeX3pH3Lh/k/YOch3B6fm8HuCB9qFAeR
v+cXaVy00ACxHeZ+NHplOjuRypz5CcX2W5zkLJBqfWxyXcS9b4WQnlBM4Bv21edYGL11PWAUAWK4
M0HJ0eCENVvgVtJVQh6SSsOn5/pE5Vt7UM2cSNC3u3inldMhiVoTg0ParBnZuTTcJb0o1NjAd1bt
/SuLTt7+kbMYY8+IgGayh/8PhbkqpAFXJ/C5BiVmaKZHKk6PgbR+JuViVLdNntyzMmVYZ1IDGv2D
8u/iP8COn8I80zE7hWYWkwms9N1y8viHXKjBtmCnDNZAE1JoTuReEoitZVfWWAvDBrk/i8mqrSei
qKfKP9IbTKOzDAckH56cRUnGaeY0EPv+3PdQSR2MIn22qajUtRy8P3kECzIPp/mjjVXiRVK8sRgK
1mfZOLqurMigc/wovj1ZBKuv72qCBbbNjGLtCw+MVgfzbpMa641cxpmcvilQea9+7pJ1iJjvA4fX
+W9znUbPYheBAGfKLisVfEfStmGXfCiq+4UaEiC9aUCV3CxuQI9gfMcCY2+OOpJvNCa568NMjHE3
3CtozaOVMY5DobeSU8VlTj9KB8hfW9sefT3u3+0+bepZc46DNDhOH6TXrMWaQnSVxrOl7qUB6kLT
1HfVoe5owhfIQ6u7V6DkpKY0XmKohxT2Zwp+aUlfOpYsiiYxh7P9px5P9VH+zYc8pI2mee0pBbJC
sosehT3TsSW+H7o60JGwa6u4DH1Tc2UGfHtIHUEX8S9zuU5FjPBw2vSCuk/33bjYoJ5tZOQH72TG
w4zONmNi0+4BBnYemk/Q2seocUfyLASe6ygD2oIPIqjpH9POVNiyQJN6xwFFL4Y+g2LUEAxuKBeg
p0pX0ZXACQGYoNlZpR1LSIzeGGLDxhr3M+fRwhD8ZXRjiftp1mIo1+jvNLqnx5JsMrb9Jo95uNdQ
pvTqKTBLPwu8EFmeSpeS3P+7N+mCscMVS7Q8vh1AisOlds1NraCmfJZWLPgz8+EHeMrv+55Z67y0
iyAlvGpwNSbmzNzbFnKfryBEJ0aHHAhW+Z9UjgoY/8H6WWDNwvzZpM8b1++YS8fSig9tWlcSNfTr
WZo1oaDbmkRRf0hOQ3hXwzQI+DZnAE3hoFKdSCTo7rgLX5Nl40vkrUlZ3xAuOo5tjGhGUDIzhlFB
BI3SabZwmNQWOoluYUfh5LeZpZFMLBRsO4raiGkDTW025CMdPq9QNNhWkVNpBZ6qxGRZxtAhtaWK
8o/Y+T2EJIbUJA7GN2YAvdj3N360G6g88E2uhkI6Wl38ukt10A3Y9OHHTDNGK7NTvcNCITOe3OJE
dgyOeABRn0PU1KUR93HH6TEQjZgv9SmC
`protect end_protected

