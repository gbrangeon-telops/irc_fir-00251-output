

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ahdDAHzz440n+Z6SrLNKLMBChQ5FzHxmtmolGyaGzRzZ6AsdM11MYnHQlmkXolfzuQvsH0tiYFpA
bdhL84ynJQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qd5Te5HYUFbAOVCK7Nrwmf+xhp7iHLV1qESGeKRRemMuPlhm9gxKzGI5glBpEm+Bt6GS7xBHPesU
Rh2RxY+9Nst/QoTZG24XGDjT8gulIAFW/37G7vhPLNVOq1gP33zQ0iNDRVgAsbEBqL2aP8fzO3c4
Dl1oSNusYXsdFmxhv/4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0n9Q8CLs0GcRArqoXB7pbLNq/7iI54QAnaQ3YfVTrcoLuaPhMipi/u1YxvxCeQhStE/q36RmAWKU
vuVvb8WRD5dX8Gc/5jIRt4ORXRhrtme6cizBVjYhymzdNTAgbAuH8k+0No3YXlnw3iXuB/bUUXlS
9ThgyMn0i7erFTJ6h/eogbI8EG6TwEBPQ11D5xXxMjzz9Q1WQ4L1w3R2CAYnCrSSlQxqvapc2X6+
HzE5EzvdMpbru1PQrGeGwaFtvlT4dq9BRwJcYQeIth/77QtTOb09uuY2bIUtRjnczrx+97he8zc4
F2HQqnZwdLvPbSwwqlsUdlME2ell5wSO2A8Cdw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fXi1UCgHICyjHcoUzs2uXfr4QL3Zd6fFq0YYnh7DHj/Uz2hpTBP/xGkihvbT84E9/Kgj7lZnbxyU
NW3Mn3WgobnvsYj6dHFEG2LfnPYpGw5nhTQMawWoftBXy0o+AjB6W5RQ99l/hgORyzZ3gEP6q1mQ
SG+9quGTTiRQQEHy3Sg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GxP7neU6pelOGsRYeMpWhq9H64emJJW3ch5ZqO94Ja0S7m2rL3jKbNa/UebfsafxW/Jq07+9ZHQH
nakVk5fs+waKW7fPdCvasFZq3bHVoH2M3uf0FMGIXnsyGlgHQ4qCnawBWxPqrfn3SKY260XmNThN
PHkcyDSRI2OjZKzXzE7AHiKXBnUYqYuy5pZkIRpG5KuuXSL3l68wM2qwWAk4Dy7OFak+VRDwWWle
Ve26y55BBWyX0cVH+A1y9sHRRFBM6x678gQjaKYO8u10cSkLQEatg4BKcHaSLpXozsPkT0ktveBN
etZKKhExPa6BnJyzgqh9xypSTFtCXtbhEF1Eag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22208)
`protect data_block
t3ILwRga+bpviomJgcD0KvFrPJSpjLBzSf+TneKsU8cftu0gjl6wShho1gXMLKykjfTUov0cSkKo
zVODmERiaRS3BXuB4beaxxY0LWmGMvz3xBAJGPXi8dOAEaVZQv4uKHALh5AyQgqBnu8UJ78Rn/XR
d/UgFUpS1MecaCbCod27laOI4ux5uA8Sz7tgsLue2HNSe/ieqiFEUgY+A7m5KxYvXZhX+iUfEPxP
n+mZInKZJzQnP/dzAWc+QN/7kMQREsr07MMVsts6jP+EqiUsNDJaynX02ZndqenuV0b1XW8IZ6TS
ExQjyOXdauEGtVwL2RfhpdzXrznVNMfvugQQKkJV59xkGzBl4M/WNAeZvUghwJTAGHCmv0fDgRGv
1bPrmize4sltYHeLlmX+cHfrUgAXnrhH4+GHH8sxgIBdaG2R8KVZGvC7A7gyHaRD1V+dewAyMlh/
Y93qHnR+ZcfhYoUIhkIa21wIwO5c26Dvf8VsvHd9a8tP3yKUTNG+u/M0Z/rKmmXDFqPdNPMeaypq
HGMmKFF3uVuUW3Tw5SSFODqn9vi7P00agEb8HcWQcW/B7h0giAz5j2o9YmpnHnwoAPXswpwv9haw
hDaOxoR2HVUuYi9WgBkP/6zCgW/yF/HRxlQe4H3jto76C35RfkW9EWmIKcDnB/E3mHVY0BhfKvc7
UB7P5sqAeQTA4hi/5EX87pBOwaYxK0vs+3K1a5PQVuPQ9vgTAXjKWdMSUYr5ir+r/2pcVnquFoud
1e9kDBIr9PSQRr1Fw9vXDKB9mwcTHh8PY/Lsh3cFAn2mvrKeB6LDgfwxtAyrO77PRsHtUSeLNRHC
0QACeHZCBxiIFYla/WII7Zxrrm5O/2ozB/pW4X6plzOkpysML22ApXeYDZxdVXunlWH0YfP03noF
FIc+7mYwsLu2Md9/flOeW5QJvUTjsSkGNHqln1b7hW3WchUTlGCxNzC01WacHH/1iO5dD15JOG8c
mNp+h4vW0UsgoaZK63lcMueGDLd5JO9ZrzijFfFq/OauLKS5wbAFGIoKkfAZQzShgxckfg7eyrmj
uHlRu5D/HZ9OOerjmsPcCzskLn4B8FinHN3wlwYCtcS8DXpLidHs0s61+gQ7bPhd0hsCu5mx0xy6
h8tUhe9TMsZ4S5VRVbSImk+q2Sx3AC9H8vz+jMO8kr1/B2/dNOILtAF4HR4+gnLD6784gd6Fv9UQ
Zid4YVq6PGDuKncUyg8YxAZ2gstJC+Pwo8sGztCLEG6HQ6KDZmI9D9IiZxD3gsdE7lH8Q4DwiEWl
Ih4wx8zU/BPIoQRebcnVLqvsn2kdxL2+YPVKd34RQmwdyfT5vp89O3uw/+43ew3L5+i8GYy5AW5z
kb3wY51LHPdONRbJogozHRy8hwQHqPQKdFNs7/4SoO9Dl35K6DqTlhYtwjLRxV7rA0YZ8i/rR1ws
aVrw2IFmaCWZvI1ymb1ly2ky/zI9Veion6YRCD4MoPpCKncWDbmJzsivZYMBfg2cYw+wbSAAHgdh
cBHduenDrYwHOTnP02seu12WQfFKt1Hii6S9fQ/Zt2YwdaPEAT9VUqdcdRVFU2sbmITrAWD9zjaY
yB+i00slbfhF/AyQoPc0NhDtwWuQLQQe7uTZK004XmorecqxGKczJwvRvN+dIX/lkiigTuIupUOa
2NIFNyt22xnQLfTig7idfC8ImMNTpFZ54vbV+uDx4glEq0bPFsk89a5RzYMb6RM8QY7aJE9r65h2
XlLGswCCNXIUAAU5kJbtD0OwJ+TIuPmBTd053NCi5eRvJ254U8iPaDEvRJXAK0tMJVjTVlfKfrQo
XRRYLUtEXsysFc7vOiK+i/xCtAJeo9X/QebDeexqj4YKq09pOruaKl/9HIGheGNcoklecmyqJAYx
x0j7hfun2zOC1x7qnkapbXhUMumd2NRQnkgWOtSgkoSQ+67RzZ63KKms8TLEf7pVCJDvyxEGje06
7SL0CqLqLVcYSDMF4cA9ceOT/n4mNdsG1p2lv1dlFnrRdoWCSFcI12xEeiB5cWkzIMKnQh4Cm4oZ
2KDawfPBFqmsduDBmZWlFkRqLVH37I0n3sBlxagMfHSzu0oH63ZSThhYKQyaPsrQ5RPvXnaseLZe
X8koFgj8N7b729xDfhas+X3WMjfRhbVH4BkoFs4t6U+FhzqhQt/0Us20D4WoI7nwf0wb0++K6TrG
pgxGqLxEsSXEFY43yhe54H1YvpcXbE5BsTP3DZAbIXTBnBoZHnN4tPKvwEB/U6RJzvmuGJgPswqB
SJ4V7xwWyEkazchckYTfnF9yKUU4dGxC8URbinrL8Ldxthuu5xxN4E02cdZbXaKdx7zlt15SGuet
8se3k04bgAWFFiJLYAG5uRgEfVYUTViZ4RO/q395qf/4ghBjsoWXfwdb976ifA4PGY20zYXi7CK5
mILE24QyFcsiIM787FmkAekJbOADokjDFf0KCFvzHG/318IWuY4hka0rAJVpTyuNiOboWqM0xudp
qnEkcs2XG91mopQkrSx9NGVNdfu3YLn4iUJREGWUzFQsVtg+sAv1rHkCxZyTl+AV2pduucYJSU96
MvnPuNJpfvkvvRmu39dtVxyMb4PGtQvOskdcZc6iOKs94S1boe0AHfscuE1PExchqEVKfu4y8COY
Cxq+nO9bWNKN1d6epZ2XKnf3mWF7TN9HSz0PsiDHaXPSpxQSmxQLKVky9K4QILyUY6Tn8EZX3+R+
BfjadRrxO5XAyO1T47zahEQY4MTVffMma3xJlfOosoJS0e8FyiOHCxpR6barbVkQzudzdSxMR0G4
XIWxe+474ZVv9I9ItS/F1DWHznrZckgmtUpHcfcxO7VNQQSakEhTpTbVnZwCd3QJLV+6BqPV9OeD
HX/sn5WTEHyR2dblRZRd2nYhrN5WuCj6yArpMMErzFrKi/edqHooHageypq1OWsNTgZcT6+MXClF
qRwLbtEYgJTR6HjBKn1QJC4ktJ16oPG/Wv7UFXL2Ven5pctgqLZ+Lbg/dgEUHL4I+S5YZt9A+19i
WE+L8rq/fafQ7jO/OOw2V3cPCUAjEkKEXyMcK0FmttAf/PvFw024DAZkZLDKmgfvPi0qjJW7qFX2
vWpIQKK5ZUZfLFrnn66ex47W17ZVY4owyFxJee+mLYOQoPoMz2zDfWn1bILdcJBNXkKounxqOmNk
ZCox6rUE3ejtxhQwzO0CCpyNaOw8b7mBZRIq8Aqq+ZeLx8+h7zC6y0jcPvxlAmRr/JHOQh25GYVg
W1Gnp6HZBtN5Yt7/t38TFhd9Fw4fNEj6+smyzOZpMj8cBoMNiVMxSFusoUDtVddxvekPsu+C8P/5
2PkrFupR8XA/wzbgs3NMO3W02VqwVpAjju8dum1Yk+DakXaWr/J4/x+AZ0JzTLBq2uayVwJ6iufr
VGTOske3vhIDVus2GxlgqLoUluN3vEd8fWsYYVge9Bcz2eST9lxK+ugdSsyCd13f8dAkteZ0Ldil
qr9kb6NCIfV2D0ZjrVK877q9oBkL7r/gDyrge5H6BOSkmyU3Q5bsKOaTZLQuvYhApEoO9MfJbkXl
fG6wV6bJxn48CQbvfrO4CsCfIocWB/l6ePQZD/TdAfzrG3UpZ9nt+yp39J1FnK1QsdVF7NpMGPsC
rvy7HsergFUcXN8ST6qZ6Q/Y4JBPFTIZ3z5oeuoNTpYSqqEwP450pqTdDLZ9AT2bGJ23b1ZGkr3E
Lwv3qyFiR/x2nAYvWrHp06LbPm3shQzl26Xxbi07xh9AYDSBvKT4nxRX2Jd5zGwwS9YvW9ZBkKBa
naJ60JzxuWWg6aj29Y2UNcbiuzmQumepjxs831bYcmxDm1lcdblAWyz1ZXo505rGgcxpKkCJm1u0
Nim8I3bihBViwJM/ieMdL98nC6JEOKWTbjzteOC2nn3uc8C8nbUmjyhBWxjWzLuu4wNGt4n92vb5
ByzmIbo5z/40nJzG0C+vJCOazYoQozVxCHnmrCU2NZdZt2LPM735n/0lJNjl3KAZ95upTpSYhnxw
9hsiUx9DK4IP0RUSMRPJrtF3hk54orSzLJSMjAC58IIkiKOexG5ms85BhyViqwtKIcnbRTK9ZuAH
/DFOJ4qnsKy1FbzzSdw/ZmlFC1MiEl761GBMqT8qoMnpG2c1ISsnixmr4emWU0D53C1ZbkcIziCp
MaMyhJV+IHWrCfEfxsKXkqJmLqHeuuykHnK4L6XsnqwAliAByQC3dN4j0L/H1qfHxYYDJ2JGBheE
FwZFR7jLV46Fe0itoGD4aYrLWlxGlRopcYFydUbp0vXFQh3MK9R5jJa11iOI5b358gYTS+pMz9Ms
wbwn40tnUFRikfazG3SkNl4zytBCMFvAgv4DjOtP8WyCtv1NnAGPL9pSoMd6Xqn2Y3SQwRTwfwfJ
xgxuxL/N8osAQWtFh34LcACVzfzBd6GLR4Jtu5mZVux/XAmbaCRegqetzsT1M488Fbq5xWcX9Iu/
VOsLKVmIY8aAl1P2HakYOyjCaq1P97g44WLgpeisXKlS9gziovQ98qOD5epG7+37c+VSq+1jnD6o
i5Zo12KqBQENQx+7Xfu6E2tRijEff299H5otFOynCTsTkHb2rTQ6jAdKuRhVsKLeQjF/SCD+cJlj
SOuzgEKBlomqTCx4H22F37gumE9K2yl062uBUhrvlxEcA/9v5E6rDeHeUG14A5njTOcZplW52BI2
l+jvVk4H4aq+RCz7Fa4dvAp3kyqmDbgJnFRLz6klF0MnwOB1K9MMjMQC2DIcAUhkOFOBjAvZFRfe
QW4t4bLrqPUDydzCRu22jqyFuslTxazJAI5gkKIqs+6CcOkKdBhzL1k4cHN2SO+4GaKo6f17sWb9
dUIlAau6V7uLtZhPkbX9P9pWTKXzkx1D5sKWeXuSvD8YMe76rv+Y1JCbGbuachgljVnhKqxgSjzM
CdsiTFpJTJgmTYbfaIhIthzXwRNb5gGODID9aOAT5NskH6PuH3vDlhkMpFS6RZW95sVNf3hrl7ZE
heAugEWDWM1/9bi7NxCjRyrQiOGrkkpgmkwMeW9/OYZed97Z3xuP4uDdZdSGlI05iFFZxzFvAwgm
8RGtmqBQ/M3XswwNvKkirO/YPHRhWjwDYd3Tp2BtQt6SHkRSFkNY7jY8DmMQq2iDheUy5VbAXJf+
h4ryWcAOlfIZfzOQL25qYICH5055sj4hHKIlg2ENWetLhTUWw3Q4ewklYw+iAnzwjPQ2o7WkpVrx
Q3nHe9ZYuLuBdSPmZHf1XzxnXyEl2nKbxJN2xp2dK/HeCdl3N1oNn9ZJ401PjJEAQh4rk33eoRti
vdUKBKlM3UA4qh4WBvdilfIKIg/iEN+uigYV7xzZ/kfmJYEl9jhxoDjh3hIYF/NXrsNmTGure0IH
UczSQLdED4QGkCw/xXwYDAIsApmvij7opjKcHb/gohvWm2N8q1HWu3ebHF7OcZlWPZ6XzPerxkej
ehy0GWhhl7GXgzIW9FUrpBeZXCF5Is5okCKOvGGXm8Ic62g3UZ3Zz8xq3MIuq2Ujws87bSxfN+hy
WxqsjGLBbbI5c3+mN5rCDFVfPj/kPLHD3ndk97Aav5s1bHMeQGdkxYGL3+bUVgEmhYSvTPs4x1PX
Iw0k9hmswwfCFl28s0tdsW6t00opy2blpJ9UuhhSyU9BRcZR5NKbDl2N0n/nFw7jFYFXwrlwkrY+
SO3eTo+ZdqH1+Nkg9f3UB+b9v+qgKoVxt3mViJ0UsYWWq/yHX77KL9oOWfyBZSy/aNyxLycd9QPp
zf7yGAZbJc8UxR8jfUwE4kcnxUsc8MgtjCq3+9TjCe8kFhzKGWhVkgehhgXE8f56qxI4T1t7lFT4
3EZ5+r5FSeXmJZc5VJJhrjW82yBmndPcBH6WLDKG+e7RMTJDP2xgN4YF6l+jzrp4J3zQsTAaNAA2
8/rs5vveWlMCq7x+y/2bWX1PlpR0l162fn8TV6FvtPcdbo80p944pEioz5qxKLMoGqyTyIlbdR6b
sRpHPoxG6LqF2Nffyeirgp8Tmmdl9dy1ZeQoCxx2OgEt7bPJBKQlWpFy7HkF7fDw8OsUa3pgSogj
KMOQZIrUO4U9sjHjpTXaikt+In3XpcqtW2qTV8YCYZZHFYgOqa1U/bComT52Pe9qfnHrQ1bwTsvI
QIPdu+Z4XBbUBdrX1n7cX5+5rulW1kEkZmwKawW4Ik7Bx/KBZeEvKHBlxkOfXXLXSQh/241tNO/z
MB5MsxOl3XWs3Mibe48lalCcktaXMclmDnFxt5Iqw/myXT1QJy5Rw214KrYnRgc1+OxDN8MYL+Gm
HRKI9baemLebB07lByCvI8eIln4X+4LeFz63Fdn2JRBjp2Zy9fxgnr0hphuI/sprRVo2Mgq4R6MF
s9q7PLqmgQke6E1eDjM+f+FbVez/eIgn9Au64M0oWS9oAPYwBGDZPA7CCZkYrNvJ/qy5mA6zxz/T
6Z/8kLJZkNFP/JvUTgvOYDpRDzBnqP2isH0M1a8kjKXB3+Y3r/Q1rhUrarCrpVfy8ZwgT/9+Jw11
6DW1HmeV0LctMhC32ui4ZkpX1WazeHHhHGyHhKHNiZj7c6+WjYdmB/QbFC8OwqPS3mVdLQ8fNOoR
a55AT/mMnD/sAoRWBUQdDRG58FZg7jOubTivS3z5wLP8Ah+keZX5eGQwiTZ4edYv9BSzN4e1Ag1V
FZxLVwezrK1IFlH6YfoggIeJuZArJ/Dds4+ZOO02q530BSvoXwpDjqxz8PVoWdV4zfFSg4HjQWYx
76cKtJyzjiLN5igxPkBeoxDaYvHUKG2vgUT6LB8PnrN/w0JXdQ2+iv5RX+fAdMF30p4HoONTtYRu
b1hBesIzvFHByF6CpBCpu9n+g8J3vZ8e9aB9PhXcwo2Mm1T0FQAAbzrCkqh+ApUuJ1x5nNQkD2C8
8Uwb2FvcqH17Nsl5X91NKV04dZF46GpiePaiS5c4y1fxCp2j/R6BCXOHkSijsmBRx4DraaYrk1Ym
jMwZKgN0JLwz58mNL9c0oVk1q5I5h3CKMtifpw93cyWO2QeHDjZITLe2c+nqknWU2m1R8yBljpQ4
AoxCADzYSGPwPXKsVhan8XauNp6TxvTaTJUZYNkCOzmWLTajy9RDqgw+2Y99zmDgJ5ZXOqOvTyAt
wnhzDTSB5cU4xBIsOB7iV6b1sutatmlMyKnDkM4CLEbGrjXHV2UNnJV4TyH/1SlOMfiXN0agHdQs
FESQceyH4cyETdYAeko9OuP4/yEK78j2QPNwgLKGRJqsAj1LUZDuSVPXFGIcoBMujvf0l2KKibQE
Sn+B1UZR536ayJQ2BBENGyRxEgfscSv+noXRoJ4EHUI2u9uyJiq2FpXaIqSlsXoqg5th9e08Nho2
59ftpjfbVTf1VSo3RQT17Avl0Wv/O+tfgBk+pQmkJdv+Oy7IEvsGudZDN6J6mloF70POyxeVBLnn
wAjk6SLTj3WZHeLjHLkNDVgsIIKIDuVPe+E2x5BkfwYkPMgDQHfBdDi8noVW45wuuAHQxpqNB/bW
PxzoBVjC4HKpS00f7aMJXc2WBAtd0B+pAH8MY0bH3oIH3aLQ/9a0+RtzSwnwmPFhCky1nyQY8qDA
dMCjUDLWuOhgjJBUxD87vENIcE9CArG0Gf8c3lziMwEqYNMm+TGC28UzKZZ7vp2jAwMgEimN8VNI
cmkxwKHE9i//q2oMe7yAG8uLfXKG/FM3nYQYew6V2x1gMbM1JqnSPoCPCmKx780cUhK47zEjbX10
CxpL6iq7tNOpXEuZQOhr8V4N0Hu7wjNig+CJvO5WrllU8E/S+KPMLkJPJG/ywCyJaK376hSY9VaL
YKd7Ntyr28OXdIiHYT9a9r/NEU0k/VrYWwMvgLt3AB713h8mCS08drOOAsW9DajwI16lWnNcPz29
1JD7N8GBx6C+5owIB7er6BuU2EXCYHrb1ZDH01dJOKF9J1lqW+juFEFRQGgVQTmOxXcWd6BHkMGS
//k1KfWeiLdY29oujnWT+0PylvTbPKPW43LdDldsLPsSW/UjMS8fzlzUHaW148BDeqy28L/Zx7pF
pHFjl9Fp1AbCISuR+J1HyHKTUGTWC+BuGC95vHSHbf7vpSERKNveK8PzOqsl+UZAVRFf3bUJOphm
mPNZjgD7Myhd1HzaZ5okF2fhe2+5SohFB+li5LlGo62Vd9WO/evA+qirBrTjsvb5NpqE6mUWQmz2
/VLO/M9nmdkWxi5CEO2vWNj//Q0tT5N8VX0EU356ow2+FxDGA6k+yQvGWTYTxn10Q1Hk4epBwfAd
x/os7SS1czcxGjk0O0aRXx8EVqYQgcn7S25o64LUk8L9VErXvAH4jXICpSUjkrey2aUMT70ZA4aX
F6Z/gTdJhzmUSQyM6hyRoTk5817oUEhPmH+QS3M5MKTF7WhF4LncwhAbUcgKLVxY5KLSySAcstTW
tdxEO1OCrvZtXlWOZvJJKlbKYa8zQXaT9JB4Ig+yEzg8PPjTYfMZJkrqcZ5TgJKQZAJ8ZYW7FMx0
nT5KihiHSFIKp/5tOwvnzjNPgEoRaPEs6qPWlMMVxCXiE3gZ74/CXVGrAmA8u0tEiylBnzL0a6De
kHBcXc84VyAQNrWBWEmuHDHVYYiI1oHmJo2df1JX/0UBpKnOWIo6C2D5k0Zyo+vnWcp5IzdnSlfI
ruPgPIf3Jb2a0fd28mwdhzVdcBOgWqj8R1X9OvuFS73w59JpujOawkiD/VKMoohuj3HfIp5ZMi36
zEj7y7hPKQelATVaI5BbACFSF6p5578dMJGOwul3UNR1D1zl1X79fZlNyyNbHHvknTainhrfWbDV
HjtAm/M9xzqaUGLY53bg4NGVNeFqknwwvSSMR0TwBshhG5x5fYoPZ9Jwt/mv9lMCfcUAILQcDZug
DGfzMr5kij1gzglmoSnks7ZWR9CNFg696rdL8qH7q8bvP1u9C0SsW6MLGRtiH7t51vHt/s8qJi1n
AQ3gHAhdglWO0MqkEsulCtkcnyqnjNuI/2iX3E/3+K3Fo4E2g2yjY39Elzq00yf2GfM7WuukWfM6
LoBnXMvDAZO+mec/KYiSm0INk2MO1C0VxwQR1U7fTUsGrej8WT+272SAtZ2MGhXhxt5kxhlTKWPe
WPOZQ/oYwdPgrkMQK/9RvyFbjxk0WcykD5lbUdKBAxddOEC659HuvPPJcXqS42y1HQc67OUZFM9+
6Vx5Fokas9MyB12Z1lPoP80BnJ/kAtKKnPPUaGAx1W1gh8JGcAEsjkBY8Mxj6vxU01BVdCgxlTEw
tQ4KusTIVmQGaBKqZ+1/h21S36M5djqL1hbA+1tRkIVM2bKzCOt5/YuYUOsNe7/bN0Nx6IdJZoy2
N2cn5baKmZUob/9G+mJJ1rx0B0gwkU1fsFdYiRI7pK40JZdeG9odDMONQ4HmMg2q0oTsxTKs7J5J
F7mWyRj/78dzwpEfGTRG/rRIvXx1SyIPps+99TnPiAGDWDJsFtEcx1qAujvT4cLaxLi5VBxM+I6V
CSgYz19YijcGH1kpy3i/SvnrSGIERacoyzMrthnC6GjTxTCkkUV49Gy0uZrMjb5mpJQOkJk5sHTg
beLzRhx6WwZAQ+uDH01Ip7WKExMDwpIGBkOsjmmmgr24YLUrLVVmbIZzJl+AU2Yf7ZXccpOYhyJS
DaLLCSbrmb6t/9eXqAkSP1x1l2pP6Cvk7TI2PILafuHynlA7tU1Qsc7XXsobqHOdB1hkcpcM5jDi
niadDlvQPxwxK+Wx678BsEhv38xfkZcQjUvpBtn8hgM7EyHoWqEbLIymhPRSfx53vicbEykf4YTG
nI8xQ7gNjixOmu1kmY3NS9qhly/yyDHsWLXlaK+WPKRTW9p7j79fdJh9b0Hg68dRRM758zR+8Hzg
cZ0oyOa2e4PFKXIcZp9yBiBlgZ0JV3d6vNp15aUXYm2Vku18OQ5yknVvXQi/P+WTzV9mlJfeIj8h
k6P4VDTquCY71BWv2wpOHdFHOplChUIiEgP9Al0pgv54yh1Nyphf4RHCYVuU3KTnX3TaCcZBDc97
+Nxmy9moX7tL/Yvy2E0cYw5w3adSeKawtOWWuRSLP/EKuNlFi4b3LhBuDA/JrL3xihcD8cKoRu83
Q3/DfhnalVJspEJvh/GNp+Rve0VYnNt1JchBejrHwq/WRJTV69GGNP3autlFIOmtYx2yCrQJ9knI
nNy6W0/boIfvADW8OfjY6cnjaEfIdBQgd1Ne5lw97Ut7R0OFQ8jJwG1otZMnq5vng4Jv7ly26m2V
TgctZXdM+X2BqDixIbH+qeA/tag6ET1NrJGvqy6rY/0ppHdq2M8b573iSTyn+0WD/2MBoGZuJIkH
a/ZLGHG2LMJ8QOQqxC9bfp55caB3qwWjdhKxNK9toccDY8Cmththi5+bhqCCb/wWEoNjjAx8S0Ty
MqthnvixA1kTtD0QdKPw37yQ2D8Yux04bUhR53JfNmhucztS0UdrNvGgOV2E1IcoBFa5zq0NmKSy
1M62dGeBH9RTq1x6g3TRQrayRFa8x5Ai4edMaeC2Cf1uoeZLtc6Ma5ajARJu5dKAPwNw2/NLAjLI
OTKuRfHRrOefUJLzIV+ZGIG6K/n7NHYXXjqat9BCJDM/RzN0mbsQ98SlEgQmhP3bEPz0CIWNz599
2klzcTT+kOPD/Iz8aCDnZLJChPeJcoxTL6KwY9LIQvXTLn1xNmITz+NsDm3d1qK1E1dqGtI+EV1p
8+X0pUIzulg/vdId1Wt8ZXsY167m0HtieP2tr+qOPV0iFa7ipzA7VIzVwf2gti/0X4I1iImMloBh
yXD5dFgVPJE/wZt+3vlXEKTuieOu7b5aDS5LVDdCJVEeYIHq0pchyMYy1/qdzNPHiG8fSCqFXMAi
G+HWasISO5HonfqzvhE64fRp9ssEeQZIfOs8CmpHZiYPph24wB8czmVFP7PmLxiSpbsLg16Y23y8
rEPziocwenuuDWLxybUdT4u2nrYkv+khEkUzXo+2Niuu555gbGX6mImVlSvn6h/9E26FfKGG0xZx
GsgHZRfxHgybOCRPOzb73ItNJntxlz23A6QdW3T5U8ISRb/8z+Dzo2QLffDozfuGhjyz9Judtyoz
WcI1Qahune36D+2CeycwwCDOlMn/bGuKBSeTZAH4K8CaLDzHieYehwJP+x+TgMWz3mqH8VfpaTjO
+SeFMz3ZkVgD2qyRlmjjD1I1Lj29o2viGWHQrAObTWtSydT1UmJiWnxjznKOc01evoYyY5f+T5cq
aM7Trtc104g6971qIA+tnul5GJKnPP/tF1d3JZrHYIq0obEfM2Dw9mUb61GhPJk+7lo7xT228Y1a
lnLnsnZpex5MGk7WG9H+b7CmcBGBLfn2XUOdGFX2Htm4qAJLgru/CAt2vw1MDULUyrW+TDIy+pTA
n0TEKMfMLX62v/SSvMO9RyU3l5Cpu5Z6Y7/6yD6cBVOQ6vJC5tz8dPjNSt4mh2EyJyCfMLhHMiWM
He9ZG7mlSPr6EoEHl1aWuuj7TdPkbw02gXdNjF+ff7dK2a9dU83wHGkrZ6+jbTrE8gcI6YSl1YYx
UaTHA+QrVxMt55GysKPL/P+XFgbpitcjRiBDhQ0FEvJobz+pynZAF6lTXYjXOi94EvMlhJi4bdn8
cS8mlJLemOMza/yw67eiMTLQCp9xtd06KqtMhuTr0Kjj/UQTKEdP0M9vJYFi9wB4OAgEHGTwbLMB
Z+22Ygx9MYUGJ17TR7gF8gtUfTmeGsrGEp6ujOgdjGzP3QADXV4KN8NxE+keVdL5Lxt43ZrqkPvw
sREtpgY4LWHOLBhZrrEd+OsLgaHG2eMARhWB7j0Py1jRjOZhSrfRcn/iKdtuJAEFLG7m26+oWUDP
Z2EHfqszdwSsRc3ARPpTXk1q4w8nTIfgkoGdQrgO3/EC53tCeLK/OtfousVznQ6+9YDD1fbwHV6x
K9fqUqoXQtu4vYaMhTNMpmCFi8Nv9V7R+A48w5eR9dUWcD7k55vPpuz/uS9qSZ5SXoOUokDsw+5T
Qn0Rvy5NtpET7eEmvJx2eOT/s9BRG9wmYSJCR3EfbP2IKYRp+HmGHPg5kjdGmn4dQB1OkkulTTFN
gvFYmbK6AdpLFh7kgw5RvIZ6YLk5ESlMNdUrOTwORf3tTwaTVM4qmPdQVdIeqwJQKmogL0EkDRGj
dD9rd/m4dBfFM01IdQjLNyY6lakFYI3Vk2txpLDncA8zUKh+8XXYNE92jaeB19GmeCfe3bWykYKc
HVxZlIGLSFqudMgk6RKGvfHOWlUMctmey3AlFtsNqr+VBOqDciLCFgBituMfJaHaE05/U6I6XPW+
DOHnB+WAhZY0WoSo7nW5pVXsreGXFvkTyHhVbK4Gmxcmdnc/OVbgyYeydioQih8hEg3VXquGZiLt
L+3AvspZiXOhLCSynsSaVflsRST1iTIKbcAc7AHrNGj4EeFJb/wNDtOhZpXNgCa8HJXkWx7jUtPU
kycQc0XMTq+tL8AXBc+lKQq3kqgO1ARGhf/pguMT7gqnsdMQqqBApP8Fp/9CffKYofMsQuPemLyN
fwTe2Db9222c0f1+IVU3iRSQ/93glQR8V191KDm1FCxOShVhF0+TjUjhG1N4kianRuzxLoBBSy9J
rMh6Pr7dsD5nsQBe/MtmBIFfn7oXjD95kWACuCPXhUcQ7M33H+7a5HLUirjtc9m6/ht64tTRL+i+
Wj17jA5LtiApi4lMKU1Vf9VOKWb96bl5q+KrGY17l9dOmrAXk2JRPOW5y839v+rR0gZGOe34VtAA
F6yMOV2ju5N2K9WIp0ZTn5iRlws7/vWBom55LiZIegJeJE5u3FhMM8Wb4hEx+Y5u5nFIwxSr6/wx
t2IQuqBg2TuH9B43bqGP5RVMvjvHctC/AuU7PmNLseyFbDQ/cFPFlfW6P3jdUNKOU7pGMc9+/h5C
UoeAtSjHwGj5jr1CF+djenWTMq+aTNw1W5lW6HdZS8m7HZVKluIwMkWZydGf2AowegHOTQGwM8Kw
IJUBIHZOa/VmEJX8Rhs+WASYyRnYFhmlexNBX4DgF9nHbuoJbhnE1zqcQqiGgPC9aU5EwPeQn6V4
lOFMI6iihY/zt198lJ1N1veoRrBrQWr8oOLobId8QXojXNN2xyHt8EdKBKDEA4aEfXv/sy+i5yjc
N2GVre7gKFnKgJ7q/oo303DQs/oJ+IisWucYdub4PXLbaFYx/tpNy+45Kq3TpT6rQvVyvyai3L+7
jbnD8NQDkO7fNLwHHY3IEGDxB8eIDXvtRgxWdyY2n/74JXHpEOwxrK8SlAG7t+ix3RdwucnNI/E5
mBIDyKrGR6A4UpHCMwwIjyL9j5+oTrdCQ/yhNPfZe/OeLjwFTIdwoh2aFdnh2aUknNmLVNbJoWC0
DMdelFF827jb0MS+MXWAG3GL3yQnTJuDMcAs8tBdChQBrCMVj7TFfzAvas8Ut+okmw6fLYxg0OPe
afm05Au4N+s4+Fjqmq4r2X8PyPk6wtjsGR1Fcfmc0pOhErBtV8cLG8W/b1ChJ6wK6owh+3qVB+fg
45PazY0pvnCaW0AHTwjvaLLQcKmLBHjrqxJqViaSxF+GgyEuBxCada+SNXsKwSAR+hkZVVEfZqNU
ugt4I0aKoNyyam33Yunlq/OpM+Uzkt7LiP+S/F9TaXj7LizjKxrDQacDK5aJQTUguEskB/z42hqu
ZuPFymZIB3y0vlN3tp2RN2JggRGfn19ls8vXjlbu+D8pOWKL/cU2CvJ6yu8nYmZzpKwh7u7k+tYi
AMj0fBXqmZmnj3bYmakFQlc0OizDmr540VrQ11hnQVu2/ut/pQ1AdEFrfhd3XvniuDJXh95ARriN
0XPd6wiJlnumQa4QJk/nazHeYOEilemDS9JuhCzGF2creEnviXqYsmBVHh3zjFGIKfr/Tv7+vyrb
r+hr7uqlOJgyfaieJdCE52WRJ0H230ZYYAnY19VhL2+SPk9VlCtleVcqjD0+XAhRJlhmHTKoNizN
8bDeI9bNyBtpzl10fMjqmxWS+Q12qaU17ixNLSPLS6a1SDkCRLm2bRJXu2tuqFVUC/E8cX3ZJ4ym
4J504cxdrenPZwiV8A4usEY72eCe/6ORb0F5LKa1q5S98nEVGDv+yidAgJPqbjiK3IrBIfSp/lcq
MLpxBsIJO79kKKnCqDi+UCcECea2pY/uoRK1EBhAiV7fqLB44AUhPnsfqn8q4NbmfVTzd673cf43
o/zrTLCSBYQfLXEP31CEGTer6Z3HWKztwLC/ae/O/EHmLP53rgEj5X7VitKFLjxqQ9y4KUYvJ+2A
ybQdvyMlLZk6aZ2CPHgTel+h2jmV2bi8D7DtNh0rzwCB70aCRM0uUO1/yovcu12ekPHvycsDsjID
y+0dKRzoYl5656HvAUMqSXbNtHHTaBi66Z0ToZDtRSIyaZ0dGF+0UTIl+iG9rXxPyr7lp+1TRcNd
UsLLkQxIwvJ29oyZkcV+MnRjH3BXmRwGkqGZ6o+nkFRZgDBfbaJx1EpokNYczYPkd0dSKtI3b7Db
7Rt7QEhsCLb7mXG0xJYHzTO+ObzbFv0uYtvRBGj2ajjhuE09K0G8r2QmZ6fdF41MS3F7lakv8aL4
S2nJymw7L9WMPt2QiusMWL381+aK3IrXgclGCJbZwJRMM0EyZ/NrBcpWZrry/JI6dR/2V0NEAsl/
L4F/RM5j+gkZxQpmdHVTiOls9A4a3+PBW3X9R3iduM4SBn14Qiwi2NeFfDEthBiLcxo0kkdYh5wJ
g5qkUAfLTndd9S/MYb+81mJ14Snm8iVAZOwUEDuP/nEC0ox+aZaO2HJa72OJ4gss4tsbTPWzNB6H
wbn3XCQq0GMOR8hwMBWFJqg/zG8ETLpB6GOSJMyiZg3eJiTsYlz4Co6v7iZXC19a7Qf76YHI6vj+
d49Wwwte87aRGEvWJV5zZOzt5M5bGTRbafeuZtAAosZrT4pPJ73e1Prny8uTqYpfTbA5KusqIwJP
6T7LzePqPCP0V/Dg+GpgNGaQeuB6bpxuVxSShdeqiho/eRRx3z2gBhweuMfwO9ygiJLqaF9qVvU0
RV8+td5DWxcdZRnCF0fH2vmStTcNcq660dBg5hvp47HK4gQtcWhcJ0taoF94J7W2hY/FaQBX9r7J
5eDUJEqUQZ5Qdkbvsz4P2wqZHTtKNbhi/bb42svvsVgO0PIz91KBfzH1XOSISRhnFKhwbh42Qwfs
8vJQKEPBRXyfiEX2Xi3aXCLux3k/rw5TANz9wmq6sHP+6vjUC1jMT4kINSfnAwESoUq9iEN/Lire
jr6dQPkv+cmlK8NxKIpe0Jligwvvqsdcey+bhNxFYn8E5LNn/H9RbF49ujT6rztceeDIzE7olDoU
6FpxEGcdCQgUBmeWCpnhPGIsbHA+GP5ViWB57g270nYkHkQuXCsmLFQY7+5RF9vYAewEklOnenvY
oGycV1JQfG+Ku3Pf9lEJbnpmtfgot1uV2BRJTmc3hZEpOuSse0+ZcHh6tjR8psYGWdi2xgfzO3iF
AmHdIT16VrA/mbgl7sR005IsquRLFfE2s89urYqt2gjBMf4X7xUJUHI1wj6jFJ2RyHtMm5q56oPm
NUVF1qdiUWanpJxkP4lM/wYz9E0NNSRlMXs4zmPYSlmueqjcWCXdv46+TBWkSd+uHAt5cQfkPum0
Na67JjWqK/DFmvRTw6pMptUKE6cws1ca4zMmX1xWbwYaZJnWIWCMBzMN+33FLH2JDX9i7HNB3/2U
jMdnaZXjfPDxeYUYVc55YofAlLRpua1+uOWLHwNdrDVZkHoaVMdNlcg8/4qx2MytUkJ+XSRKfVsM
kAmx7PsKWCOYMyfhD2jv5T5gHNoR1KkR6TRBidB6bKyj4xhcjv3sln49/byxPQbZStermtJppW+a
ECkRA/1oF9JLaXLFcm4ooDXuAuogt6xRwMbQUHGKuky9FkBWVWim0dP3ZAhgB0rHRkJVZUss1vXT
ES18m3lK8VF2eVyxZIzNskiLo6p9oQA1mfUlPJ9Evqf/nGTWSU9FlKMjAJsyMrWXMM+BW7swIlW0
mGd8NkEvTxuYnjuCGnclSWmUcFTT6LMCkwI3FZcpCcwVS+wt5UdiakDKLyWJ2W+bPnrtLlMP3/eS
tQRhgUUw7HmNxxwPZd8oP/knOEmZQADo/T6ztcIJzZUAjM4vgS1lswGNnfCoFRwRCiOG20rxpkI3
iYbeMeH9rj1aeXwtgC79zrBDV2gAarLTcfLTqZ63Vjne2WuQYqxF7Xj8HRYZE17rc20MRZaTOhXb
lSHj5jPRHiEqnolvjUw7zs1ngMnBaOFSGAkSOZz4RXt6fUPGmY2DRDJnY8g055e84A6uEF2Kng0q
I6hUDFRAHBscKupeNZvLmXXVb+BGW9xGAL9TzYOinecPC+C/Y3luMrxW92PGhBLvxjpEGV5aVRPI
MwumeVa3tddlRSV7EOiUh1+AA6l/xlwiu+Dn5ltEJnrcdX7sWGq4+eaEH2BA9xT3Vqg8v2dJBCQV
TXCb53exUNKm5aOkUqLjd92ebQ87l44LdXYyQ5COSTjJS+wX6XuoEhCTUvlz163LJkNtjhI+gkqC
yrY+sq1uS0g0i5Bzw+kf7A0YshyeRPIr9tZbL7RfpHXRMuP7lChVP+DGm2qMh3Xrkh7rfPyU9gGh
kXPLLj10EvbtEIho3yWLLDjRs+n6OcOGocbDE5Oigrs19NbnyRlgGIzoEMQjTnqgNBW3DTGJeTsd
kQcbugm8v06BfXuZar8K75qWh9zvPKTI74Z5smgqapvcAxG9wANpEWkAlM3q9IqhDdTBIa+b4POB
tV7BIYowgHBACn/Lf/gBeIEhyhC9smeXCciMFwiI+bx2V4J5UNpfEI1QaIkQMvgJ2fhjarkIapo1
eM3uqFdULIHUIDrQeyJp0Vbe8kurFyq4Nwc3d6YZF0erXi9z8NINN6wYJYghMjuBEAt63C5bZkap
gVyA6OnfhGZh3X3114EprIzaY0AbOeWYl2r6rmvn7mLkjqL+9jovewxWX4W/Y73L6QLzrSO3hBzO
7rh5ux17HCypCsrH8zlOv2ZBCPmZrHweDuF8HY8VnPJ2yx8WPMturVMp7H+YR7jr/6TEeZ9Q+Bhi
e1/maHEto6u3GM1xWN8XeSQ3wCjfTAI0eQmr9EqAWMycEk/tjV+9nDfnXYzggJw2ADBpmx08rvYj
24PRUnjTCoYMKyXqNdIB8ib0tRcHej9UuMmksHiNeDExkFgjSjPYE5GJDZjxrQT5ArXvjklLQBDy
xBX/DvXSoTkAxQ5LRKLE4Sya4wpGhBYmtsqaU1paMrQoRvCJuO7Qt1ootklSipd1OeVInKQmXG77
iAkX3HVcSetjYzAwbTaHWhz3RowJD1Z3HCsrtfh66IciPdwbyo2M8rW5UGobGKhGImjsK3lUzlKO
v2ybmxTZwe836ENrUYpjtTXcYpNgVGyCfhakur9SOBk07sg9vri3QDFFBrUo+SzKsvVeKgORV080
+Fq0SHaKsRuU0LIHPUhcfxuuDUxgYoKpmDb5bONSZNF6aeEl6+eduQ66qRdjlrTjqVs/vaH1dhrs
33zWBe1wH4UjUo+zcWvUHonIUfq1S8Fa0xMufV6T8JNSXErIbNxQYzLwX1N3i46JwdMZYl2uJpzt
eWXuEoboZv+KNOCqaSqhPcbF/JF8K9w67crRh7I9Xy2ACnz7WVU/lXnobD0Xoco1aMY9oDHfJ2St
aXODeSCOL/hB13KpEPKaDrXI32xlM5+aoyh1sLCYQCuJKE+IX15djcPu0X7ge58ZyadUALhYdIqE
xyD7v7341E3sJFAi8p5JoPsiQ6u+C9yZ6zmzNVzPEYmzStkMB0zUgh0BlGNhvAem4MC0V0x4T7lm
uzI84l9DyuKOiKHoEU5cdVKBcO/NtKZzfov5hR8LNkbfFBD+lO0Fcg036r6IaT2dniSlkEBgssuT
drNUmpnLYOMRM6Ci0KKF/wGPM6fmteDm9UfWLayz77NcoagaQZwR5f+RvolgLujx5xhGjiUn6EZv
JXgb/l4RNMEAlmQlWQo3fn5KVvNreA2X2s5gMSuTqK4kT/3ns6aJqQ5E4W5DNpE6uAOEYtxhKTeK
Dqj6mVHfcOeWBMQaVz5DDMpW565orLip4FyM15npsHf9A78RM2gfEnRL3pVFFFT/uHzwFo2pyC3Q
tWRy9NAmeiLHPMlPQi94JuUpd8DZnKiBuP5v5fN0EZGpRHfbT3WiLrVdL3V0+E6tb3s3Y8fOrAPA
9adXNdqKB2AsfoR6ht+nZYgy3cxN9W3RyG/4BJWGGyl3CshAAgSO4Lmhog9jQPRJj7vFoAg4I0cg
jNsicJAdTLYz0qBC56WOJuSVve13N+Q19LehPfrrR1dXNB1VmiG1zrrelzZp1i+5fLUqfXVNaGxb
72NIS4g7p4YMddcSbOAIbTFIm1sXnXcMDrOmxkDIdxY+AN10McDhGV0MzJf0MKkXcmJPdgd2yr5E
Av8vZTyKJMl94x2H9Rb7nVYOMYC1G51a72d5dNPUKHDGHHogIvitfpKL+iaZLNCB234B4iGHBls4
cSER4GmtH2hT4xLb2fnPlcc8YKhUnq8ZqlOWzSmP8wPnRMvhRy+JOWmoartE9rsSrzLk3Lv/94Rz
PgcT7+E+b6a+d7W5u6h6ofuES7BLQl0d2JAiXyI88Sun7nHC0k42ZY2jqLQdEvU2tr3e3jVSiPkB
GTW82ejE3eQWkYT39pfaKQVT/PS+492fzPFoNvtFmIDhdHy98vW2mZLjdXTjEuoJv9BIyFHTR4xy
aahCYeu7q61aAIfyhwXv/Wp6UNEdPmNV8Ec1KRDTvuZBG6VuX5r7l9hKdYMXO8qMb8om9ZTjVBsj
uY0hFv9b9DmRY1JsGgLwfcdS5hohZlesddEAke/iFtbeDqAfx9kX1DiWR6AAasWJcvE9RKEfFs0g
EO9fP17Ag7dwbJnSH6Jp7MmBCr8GET2vkQNEO/RNVBsl/H382X+1O7qt6Gd8GIWnDgmp355ocYbW
FK/jQj1Y132uk9GvhB8sfRuXQVq63yexOhVJWAGbNPQulKC02xK0ExgkgOMIiBgU32gC/oOiq1kv
8H84JhmboC7abg1WHCk/l3z22bKB4T3ZiqDWcs0Yo2lNliEm8RQpKRQRz4+64/MIrnulVCh24baz
1ElXCtGYCFUuIgMdQCygGk9JHTfXfxiNDRClUWEH52QQW1+iPnW/mOjtIH96b0F/dn7JoZLBoS3j
g10U66JqY6S1cRZ1dnnCZAS5aGcW/gaF9i/buHvpkda9FfmGPK1UgD3xPhKftuVqWtH8toNX+8sh
H/egoHbY5c3SgefPHOJvYaKzoXezTs/xMn8Oo0AGLQxFs8DpYqQj5VgiFwdXKITmDse9pU2WoDYm
x8FWm+G9TprAm6pAJLEzDlG52kjN5Uv/BwCGYbVcYm9CUPT6KkuPyxUOkDGrhy8sBx49m5eotPW3
szczwVpUTO63jHaTdfTdCYdydsym9CdYpHklYbT28O00sN4DoIsV/bIXpWvnfjsTyE1wKzEgoh/7
911XiyQhfI5c74ro0TVZiyQAQoC8jVHsXmDTqjYf2gyWEqTO2668UYOxLjk9uolH9A9/j1Eam8wM
fSW38eAPhECn4hMsb3ko8bUzP9xMPq0zerqJ7QX/jtHW1nSlZh5rQqKNMotOEIjQbep9AeGAXXcO
SZDsjb330WbdTI/ivFK/KXI8Umw32vm6OxL6dcfB8D+DERofV3nMeyqYpEXQ9rHOjrb88fAkTUfW
uSt4evBRacaoQrZpzrFNroF30Xn2KtLYCHOsMFT4AdzpYj4Xt18YJ6BftYnLsuo9rmN1ZdE7fS5z
bVT0Gpu0KygYGigB2x/a4ScFxR0wRl/2ZLbCudQ0kUtp5uBz6hm9YUYJv2DnVzYySIFj9MagaJBR
+e2APz42g9B8YZZRKt87A+VkDOo5BLVk099vRZJZVrJEsY7UL1yLw8BiEvOPY4cH9/RZ/KEVK0Dw
tSG+8agdp+EmuTBrfxSb0denTT9d5Eq3DtemLSS8jx2NPHhvU6zhGEgmw1lUSAYP+ScbluzRmtq2
vMnRqkKH9s6J7WqYON5CK2BXHRnqZF1oRNw8JwJSn/2ccjI/XgKkSX+Zi8M9ij2Dnk9ia5LUQBTZ
Nhxkav9oNYa1ZCVcOi9t3jYveE/Y6jdm9pofK0KqoQ6ufbiMM78QLXWw2sGQXylQc4DaIh00mQkO
axnRZD+ZwFHW11+AMgM0yWH2I+Gx4zcNRnU0uEFH7gkaHorprKtzq7HZuvJ1h0dWeDDAUAI+XIEG
jd4yTW2e5QXvE3h+OCdIo/YW0FAMr0+vcSpbONDETnC6fDzlaEuQcd1p7TueQ6170PklWu1VOBQv
nflAaj9vOkeSPL6XP5EqAV0m0CrznF8RBggRgShP0Y19owf/Y0PotSOfuQTC2WhJoCjUAl08Udr0
UcrphE3Wc8/oC5mAimpeQAx95kJqVxwaNFyCsdXm1CujKiEi2AEAN1zcFBCr1d/ZWDlEWFM8Sid2
Hy59CvUGaJ4DYU3zCiWCuT5UiNj8uKmUlAGp0mfYAKg05SZJNI4og6yqKrGINsYSBqFlHDWur0D/
RzPShU6bU9NZ6txiy11BhXl5sLMxgWhfhwB6sK4ekfpaQ+m5COZkkYksKVPUYsG2puvKf6v4Rrlh
ERaMT7lwJl9Pzd0KOkwJDB7mkiaUo1BVCelObqel8Nxvi+DkOoOG8omPy/5VKPXX8Qv8pemawWvO
LbqIKQ1zDhhA4z/Dmil1whQB1RCxUs1aoEvjbqr7i3eyNgD5pXLYjk9+YH3vauQMuMDhwDiSPqP8
YyGp3ba56hFQ5aPGDcftrBFUwie5MO0tCEIV9Fk8guGF4LPnM2RboU6rjYfH5h1fvHjSNPhyNuYP
2ZreWjMX20v2sWfd1lTWq72S5r48BMh6E9nUUToSCCvqTcpGk1rMn5R3eboRzn2myrBBV8v4NVPj
qsv0KJA1TbfX/LjiWUXPGtJ1HkIxKRw/lH6c1ClEpGzMLPCW12a8mYq2H8KmtQC2hiUTsXxXJU89
qe8C8ymt2/P3MyXdc4unxPyZdaRI+UjbJIankbMKq8biEQE2gNam/c8gdQtCCAqgpEOpElUMfzod
e1Dqaw7IEqvAoXSK/KMbh2scFmGxsLXQi49azZiiEcngdNUel/GuxkxRtV686e1eQmefO+CFsV1g
elUBD6YHYHaTpoV26BKyYQjBZcIFn3xb5e0xjL9VIL6JesREnTq7SEOR4bDHL1ciqXmU3slSlkDc
ZxrVJYT+RhK83gRJ0nmjLU0/qRzEcFAJj7mzqqHQyMv3JgCGQTfsGuTJUd7tK2kT0g8VPKtGswL5
DbQlsamKBKF9W56RztOljK0D1qFNsY3xN6z+/4gPi12XRcdFwswrkYwPESQUdPcfMRiPL5Eibu+3
061rUcqypSZCNf0WMWXF5b8fOvXtWc3gpc4bIKhmbn17vjyQsgjMKaAkmkkCHkk5p3+Z8cJTTPPb
My9kDo2YC44pD3k40aZ3qNBatPAOlYDYrlAP7463DiukEpcBA2K7qfud23xu6Xh8+Ba96io51Z+F
y+Td3dcJxMEGvJZ9/Ol8NtfpA4lyQdB4Xwqs/ajVkUPjUAzHp84sD5Yn3L/3TwE7XUSG0yWxAsNx
avvc2/cxwQB6MK6H6SqVXAmv0F8SCTkCfS6vWt9Zeds5gwLhAGQJopp6CBZtwdIU7AqXKDlOwllx
TLtDLZbr/2MFLAKWVvh+I+oab2qCo7wzwtSmkTGYWJPCswHJlOa+gaBjvmhXNE8gRYAaU9X5HDML
M6ZKCvJM5L+Md0OqiwqqJ9QJH8DO9/f3Qo36R0TZuO6q7qQ8LxtYO1+jLk366NrLaGXL5Iwur8hh
BiQdZikCuXeU4gvu0ecuqYj04R/bCfRaJz0yAEuOygRJ6Bl5U6+c9UDn3bPUJq3LEKTzgXCwGFr2
KYaCUik2euDZfJInzMlb/atOXt+GaDE+/+7EJbhqD0yAVVi3T8Nt7mJYFx4TxOY7RZme5BP6Jk6M
uTAj0vFsYdGZ3COrVMT0elbtj6VkJj507Df0jsE+VHOj+aanQ25A8nsQbN1hZpqPydXI653koNDt
acTvq4Raf80r3FFj4LMJgWdHtA6PTSUWx98rRZhHY5f/4ZVY79oUi4xRb+ho23qRKLPVpMQHxsaE
t3BIvRgkl4sOv7yGBRe7gFKQHARfRKjMU5WBQmjuLgM9F1ujsVWfthn/ZSuUYRAdC1mZ7JMPwHvA
HrgO2PQ2OAE5I8yZTiX8EgJ6u/c0M1Dw7jbnanWF5B1pMYCMQgQfVMR+qftOfNPiOiAJvV7tEKBN
sdXIm+xnugjFIH96IrZKPyen8ggbpCmhUhVVMKDAFLcGrzrt/ELl755qMH+wLSpSTrcHmySboNy2
Ttl1GkeGG2RtpDNJPFogDEOGCQcBDYknxyQlbidyto/S2N+vzWqRFqoywARRDvVfmgr9Mwp2/ksK
shGzMp0S957eO7vouNgKcdud6dCjzSqEI1dbwFAx6WgZAFpwtTEYLiyC7anjwMBN3f3Eu456kkBo
JEoKwyMxg8g/+fyKIlu0YYcdAzxf7nmikfv8GGNhcJ9mBWIOzqa5OB3kmpFGZlY9itHaRBas7W27
7s6/OafoY2umaGHQlJ+g6QP56xLdoDrikt6dRrLpUHvr+zTqAGyozoTpnEgW/y2f+mlJuKMg7Eel
AOpOLfknMfHW86yB2sV9Fo82wNC4XBU4x0oxkuWqqplk0uevLMGfuVkvDd3P86H+qtfYtUgo+tav
OZGYEm1g8QODb6yk6oxbM3/jC8Zkyp3sB2zSQzKN8kwvOil0G97kSGak1L78Sj4ADWZomSohnpPd
cKNmODpqX18eB0r7/Q9U1VKqSkF2vRm0dJLvI6amJuVgFL6E4stdEIUSD3qJGuFr3FW/Z0k+mqfb
eKsCHVfB+YDcPCSAFgCZ4hUnkfNAieKfHoOgBKEYbRQJBpC3OeONskFlaSC4JK8y2z8sbmDC6SPs
O6UMHqbK1+iCtPd8+hs7xko2d/VSWwimG8yaavEYkjVCckWO0f3U2jtgnuMN0N+NviHUYuRFKJxu
LCzS/Y+2bM4hJ/6zDEKWWXSiyuELieIy69UBW5QkCY8oIDa2UOM3z5CGXtVDdteRpLgEEksQeiJ1
0cat0w/KldlI9VKf8gdirn421JOkkir8VSlDu2RDJzKZFa8YOYsfCK1b1YlPLbLN0zzUVBcpCjs6
okiWREWPaYYQLX/RXLMjPa3ryUdyPmg9hv+PzV9D4J0Bl4jqtBY0E1Pq6HR6NLuZwot/EcldH2ID
I4m33UKT3Xi6NJeC6W161zIDZA3EatTaribjblJtNhtjH4GEiiU2Zs/tHrs88Q7HXaXl7YzmNHzg
iMtfB80F6cZx+bJwLjAXNu0wX7TFafepa/SWKJdtVvM/GR/2Ayr66bgYP0N0B3ygMge2a7e8cYCW
mbB9MRZaXQAQM9g1e7K4l15LOjNRgQm6hDd367bFUnjlzxMCBY2o0L48ciMIH7Drkw6y+mBBdsid
fe7LY4vxk4YRKQpTqMECfucCL/e2XgeRSqlVvx4vIpD2GHMKLpEU0lF06qmRJY6u+BdpzeyG1o8n
8WTS9u5CGr+QtdoAf5gkt4vh3CM2Andr4njHX0WtIyt6bGCTTadhYKKDI/3xQ5w3KzaQ2ZQq407v
+38XxmFDum37Ffqx3heDCSu+dIjuSEibEGS8J59tfzEDFRgbnDo1N3yBM5UhqYx/V61jb5Z2Hkin
XMonoIH6xF/QNhUYHQryVnJvh58eQYhZZceQnUdDEZN6h7/kIWyWqAEKGl3h77DdCzVIFvBELZKI
Wx3h4ZBYNG5JKG0TQUfHltLJ/fU5fQVqjRdDVLiup3gw7AmaZdALarCScABysScWYcQtLqNpowBi
iTzP22SgoHnDLm+1Vbq9qkvm8ivu0ORIkRRFiv4eEUAlUwdmtND1/VulG4ng3pcsof1ghN9wI6a/
RfqaYLWjoywX7OOecqwiEXx3O6gZ0QfZC95MK96otd+a6/PYsesmFyMsZys/M5IlZ89J9cO6zm2M
YLQdpdWkGsEg8BVTbi32mAzA1u7PJIU4dJeNfbOwM3I2mFYhMa3BRax77O+noHMvhkA814Ydh0WL
hKSe8UZ9Hqp36Emv1lUJVBBuyA0m7zVuyCMTQ8SGtx4cVlMz7vFpuBU6xq9sgsNWowZV00ICrNSX
5dzXGYGKZsQuFXkEuAz1sfxH/xaqrzm18CuDP4S3Ft609zs3Wc5dOvMwzFoXIty6mybWoO8jVWQu
DkVDg15gjhPUTjMna5qRfL/ii7615v/l7UnE2ZA2QqaeZmEYPxyRgYdYVNLcFoleghoRcjdT4VhM
jVvU6AJSqj+Z0yPi1vOLKAtEZy4ukbSWzm/1/aeLANiQP5gS+kRW+UrvPBLWLigvHVYLFNVUIYMr
+NJa2g+EPmm5Mevng4fJVEivWW3VqPSPryZltfK/aK0bJgQqrw0tHfwVjklxcCeejki0FCZHKf4H
smsW1huYqh33rU/AZU+nHVg/qYU5mq/rXeQ9kO8j/A0kz09XbPPT+sxwtKnGc1rBxJLUViWl9raL
nR4nVfYR1TAxro8amaoQQ94jzvzIodfcgMr/hpeWkVS+tZGxGqXHN0kygvbdr/Fzl8Xa7by0eeR+
3/y/yBeEfaQLQEQamjLrOXZc2rGc+gudf8Pn2qLAa9haLpZO+rZjeYnwLua4bdbbnFJkDseFZ1t/
fkQKwj9uK6mSnydlzomOIGwSoppcdHaRAdrkyBZ6y6AD/2r/fGHJjFd01c11O5YqQPlu49QvZbgj
WXXM78nJBnvYJ9DFAkrj7HPvoXzUYpIMs/uUw1Yeir6lZ8C9AzY66uyBB1Hbm3kROh0DVl/mDK9w
kfN+/3Csj6KtSqK0jNRhtrhcf5+WkKM/lwrkws5QsKu8dIWcX3Det3kt8O9lEDS3NJ+WPDWhjrJh
i3zOVu7C42+xzrNiTp4SxBbprCGIOmL2fokAgYeDMH7TqZnD2rr9ukIvvv7B3LsLdW8Zw1UnhA0N
sBcuIahrmumm9NYTJPdI7ym56nAgh3dKBZ6duf6yQZ0eKFQ/zJ3NbGsoawFqU3NtURXJ7+IvLnyP
CyC+Sbe6CVFcHFp+w6SqSFgP4e8SioZVa4TWiNP/0PXLufEMyVn5nPyncxxS7Lz0sG1Rk2jynqqP
3l/fj11VAfaaAz4jE/LnHpOn29GwJseEMftQcAvA0sVQkbitDeEvZPfqNd/Dzdizy/5JSLVBAyhj
Uxjp5nuEA2ipoeiAcq1Ijij5aqjEyy4H5sAHnpGMhRVDyTzsO4GDb66ZsDMoSSJZ+sEXuze/NHKN
Z/sZd+5YFllIDEyJ17k7SPwX+jYb5cJ5djmYOv6U3viYJ5CZPfyPK3hENwS4x3Gaz+3WzzT8Dejx
HEICWVMZraJO7OjX1oWyextEfFF72CszVwplvaPtrFuebZfYBt4Qf4CdKOmu+l7FnXAbQntZQDD3
ZV45LjIev3aJE8+C5BJdkWbI+XwUq3fuZiH0dR6CneIIQMSDvwvbZ5wPS4MRd1Xes/LR+zcqvDoN
VTfVW+i7IKhApkSjl5QG+IeujidhY2qIazG0zAS0GgI9Ikt0smVHYEVmbx2599INZ2s0YmwMP9j0
huHzQp33DmFYq7IBAvnLoYWFpQOQgdhsscebBQhyUj7kdXhRauVdIXtV5+f7SpLbjbNTIusjLr1W
+koXZqxN1oz/qqAkFKNd8GmratUwwTqrebjo5FJNkOe8I5n1DKNxXJNwYncX/KGetzToLJ77nugY
KvZmS2L515748/143dbyDWsF488v+RhTtbaO6CEx74C5iIw8llxQBppnBEaK3v79zhkHpxf7iORb
r30FNwgrwaHn9ZaxgduL2sobP4wSYiKECm4U6nARrOP+bCIK9HlgR3P6FMriwyokhyDGcraFtYJj
EaI/SkmdjoEt2+W15mFQt/fSPliycDilGlSaoNIM70K8J+A3/E3lTxjP0WRterbyhmWovpoXEmFD
RWxwtbPvYjOTFRMBIOFBU2rE1BevlySoIkTxf+DqKvk3X/ia7+KRf/5/+iL0ssEUBcNLt08ViiUL
cCdCCx1FB9LsTIL8RVJG7yhDp7/Xy1V+GepweJRD3fkI42QtYYktmbkThz+/eH17AkuwKNmWsezj
zBnyh77ORkIDDXH/xafZ3g2Rp94t+bdW/L67XLjTwFfLJfrxoG05+0fEbze91qgoueuOxJm9tSbE
FApduWLp7iDN38Nf60SAkvU+WTeQOn0OZXcZ0qkDFiZueUUcvNFV8frotNF8btKhEKU1g8DHOH4+
yIuixODkAs4h7pLSOoSKzS+aDWeOGJvpbTSLkynsJasxm4b/2yOrKLMzghiOd1fvv53BSgEhqX8K
ISUlALj+i5F3ugPlFaYr3GKx436jkQhdmpuP4KbCxRa/fO+hQ8ky6zJaqo31LEx/gk7A6SbrDyLC
Fqo9CLOcnStzLdzeZcfMx3cla0rQ3SwDjodSbaBeP/52myGwkdfEn4tViHbU7fgvIvx5ER0s9Nvd
gLRL1jNPs0tkG6fp13t5/y+z0z1y8B0t+RK+CwyFlbIvgwSbeZZu0VYVf2crevs9YLOhGyDCTjkE
aNLEFqpTfGHxgbjAdRaw927ZNiPZis9x2FM5rnS/C/L3COpTx012NFPW4IptLNd4WJaBDBSTmxmJ
HPsvzImftDbqTlwyKYLTmoMQBAAZNU4gJPhZdaFvvw9jk5SKR2S8NSShgWN7djtiOYn9MVUs+ZVi
oZ+1iaeB0DBoRi+ggwoGA58ZCH5pY2OsUxxOZifqF68T25Q4pC9X8ORKJoKAgaMJzJxXlw8Hq4/r
HXmfD9yZ+MCCMeTPlEegzGcnRnimOSfpg4ioSYwT3axhrgaIi1OWOCg7H0w6W8kZj8TVJ0yCkVFs
WUmEd3qPO7fsflF1WBegjy8obv4ea0bIHpU27eErmfxvDBPzfPABMENjWsW0M0QSjJCvXTJNZxAR
ClZX4wqk6Rez4dzyMaLuOLhcOC3BVXfftouyFewv0UzAfS0FPwhiXIdQh7ztyhnDyg16H4jsVPjn
zmN328oew5eRZd7Tp5I9CutkKd5IG5LBeJJDdp2b3FaJ7oJn9a4+MTCXkZMgU8x61ehJ49Ywamwk
fHqLekXLXyMZB0HEIckJ85zK/wBEUYx7ZoOnLSjTXgc6FRikLpt1k5HmTaUJWt7b2b68YcJosnZB
KvmJ5krwiBpFpTeQtIeiQ9IdZ2b2IrtlmhUw9fC2No9+CZTLzh5fHYDFP+kKfXj6r0NqED72tuP7
FEvlKv9R6BzDLWHQxq5hcGJGbMvz0NBQ4P709TLiDgsXIkMlzp6uu7qlMkSWnbV4HZGmjRO6OimW
L4sq/0EKSgmwY2nXFHlzwwcZ4mF/zhBj76QQk9cUc74eXZJkzV0cglRrGr3Kud+7EmnOLvJKl6Rl
ZHJllFQ+kY+MyWyfUrxk3Ts2c3bKYJPhSkViP4GididdQHSciFA1mF4qSZj3ZPtxRkrhBaxerQtU
WNX47SQ1GJpPU834Td0YRf9ml4xXvPL7OIm/RtLvIT6MO8dxN8d/7/s6aCJNDzvLm5e2fu1Xotvu
Zm9gaspju7+r6ItYiNBzR3uyZUEz6UqCpN1QmyYJb3rRT+pEGWI5uCeYtYRujN1x+ZQg9p6nUxId
LtuNMRRPPY8AeNrbpKNzFba8sm0nQKqBdQwjD3y3Uej3Pkh1VYU6dB39kNQ5cZOyT+A/JP+OJXSy
4w8jLHUH+9+3ao5QQPDGPjFPMOpkp2/kA1LYarGQxG4v+coDagddOwU1SQ8t3y1GqSYs+RPksEGF
RdEFG79RMZhqqRc6lg5xc24sNMx5jUQrNocdapP/eFZac+3idvOaMZRTxnz1h8Txo50WfbnKozZY
tWbwmVy6oxmj49mkh9BG8n6oz6RO3InBVtauXdpBRq6fnawPeMij47tNcU3bM6567Kmrp2r5ifSq
eSAn18RGdUdVAWJkvZNgeUFBKa7NTnJWFSEOxX3mmbL3F4zzCDNeYKZvFpHUN3L7XOpWvPDFOBvM
tPl8/h2lOm2y27LucDT9ta4y/uw9Pe6iYJl2b5YJgNqdQA0s1eW+C5lMwGsDfw+kMoiQRKh+M6Dt
oEK7fROVMhWcZs+ApWPoCOnHq5V8hGplTI2AkocKRbrhTukma44ELyGM1lNA9fRvCogqdJMX0xNV
gjRx3fajJq0sajX+oWt3ZjjXn5oM8FkZBbX298gO5ji+SIGHZj1vPNKbtWr53lxasZHyiIM/koiG
Vkc2tS6fljktzkEavpgbfloRb3GakbZHygUksw5ONyb1PUxYKQMnHB/i+EyMYz4RkObwjcaoS/Ms
O1tMh3N7lq6wYeJPu1AISMXDk5ARLTdL9SRPnrB0TMRlIu6L8HN2IqbJ645H7PYzIyrWd8zXBtC8
WhGYeKTtur2RqALvOeXKxIvNX1BkGDuCZyvOx3oCyWt60TF0mReHGGfi+8gi4cNoUcqIYME3j+jN
cMVu+4dD6gojUdnYsburCJbc5NegIgG3nuT7dJ/qs9BnyJx0B7bNjVreyNOJjCddyq4Y62S9A1n2
NP9JyHgxIFiymbXRTUXAbm/D3ozjzJocPG4d7swJ/QWjJeUSTX4WLzu/kGV1YLm4Jux0/nNZq297
7NADETS9bKhEGS7ykBLyp6mqnqKhmwp2PGmItfPF3Oi6bD1tCISQ6vEU15nenavt6mF4gxuhWYgA
0cp2MIcdAi551nqowvjkpopQAIgplMtN6WN45BzUFo+/lOMVeh7DEALijg5+JrxdZTl1N22GTd5V
gqTQkZJh8/BCQSTvV6djmYeuEZ2aKPilIP5ashThL47Wtc8EeqQNZD6ItFICZo1R1lMJDOlF/LCR
mhiQK7n07VVB1aV1QFqVg6R0j8T83UOD5Aq9f86KfuntTieQu//EnCz3DdRqA4JOyZSrl2x7CtQ2
nD24lLIEbsYUH8PdlAO2+wQG5DSSi/D2k2ZYJzR7j9gzCyOeN2b/ZnfyN6fJQBZCouHFKQ3Id/sc
GvNE+Wx+cPOKERr84R/Tb92kIpLcRH7PovH8cxlkyaONBI8R4wez2KrNGyAOzoJ+/qnWcfkrafDH
kSx3FOsc2zFP1t0e0B59fV9N1EDICwURTrXyu1zS60jtj/5sChD741DTRjA/sPcZkP/XhYFuslFz
BFMNb98tfENn2z1O2NBhQ9gw1rX7N49HM4CgjWaC7t5JxT9iNA5VnkBaFnMSYw9gwZSC27PJV0Uz
mi8YvyDcz1wV+5nvgPOEb4h7Bsn67ExkBwfD+qEBkywISMb9TfvLgKfpoaY3n101HCYDkOJlNAtU
15VKpSJsJVmubyT89bYUrJ218WcBLwm6BHQ2+QUaszsYknODwz8kMZWsew4Mbt5RObNEojZ8NKx3
do9Tn/kfj4mAsuMyDQBzbXF2vd7IUeX9Xa7lybswHN+TDhof1a8IfmPtpn1EoyXzh91B80vl7i28
2VexdRk9hKwRsOVRsIsUBMeDd/HDAnhs0642s0vJLJhKgcY=
`protect end_protected

