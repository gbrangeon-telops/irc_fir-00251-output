

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cPZ8vU4rKWICMycnP8ASghxteX0KiiSQpWJpCIK7voNSpkWhaLkY+/QNXKrCWexA6C73eW4MlVqP
U/aYYyUL6A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LGoeeEeMUHkj3xBumwl7JSHXwdKJWR3APWiWCdcCy3wVC6g0GScQrp7fjvXp784YBiHqjtsyG69d
mOZ3fy7Gj87kc/h2xvc4Kp6GM/IiHJc0mbPVp01AJelfAExlIEaVGoQkcAXR2aVikeaMxuRKkb9m
THdehu5n5eHx4/tJQjQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aia+xx8RLMhA3IF4tHoW0Vw6LtYVDVgU/c3FBWk9RJ/SaLw9lkXng6eXJGNs7uUJXmkzrbSEXjkp
9p7xWJMhovE7nwsp+7RydSgRQ0ttqPUbPZE1eqSc4iNU9Q/KQ7cPFMFwb6o48JfKidjAmSeXX5a7
n8A9TbJ98klc/V+a8Nj+tTPfVP1QI9dRmdzaW2w+actp2BkWAgSALKaGkzvCVGa/MpfN/fdLNjxo
VsiL86HW3arw5N+Ra4HD3GVUtLt9RoCCVRrMaYywuIwp2m+MgGVDwi2f2wZCZ3t03UamXKangjoy
PBei/XvAf3p1OvrOrKNUCVdwEg17DQWfBwZyYg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iSq3so3iXhp8LA8lrAo4ElVWkZ4sJhg+rWrioZWefLcgVs70gDbHsh3ghf5w2wiNXalSfMYzUoxO
skfS1+28WFbvBvygndpiSNMXeXmzWGrwBeHtNO1nR5azyndKvNsun44/B61XF3kTINCJNR54A+3f
0Ezm1jX/FmstQisPDpo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fHCdwSqtdLKfkpdCYo92uS5kFXmPpII38bIISEYuCqZyK6/BVCrCUL1HNVeJEgqGnb0uRqkye2CI
eX2LoUaDxy6iVejnRrRRAgNtgrlZcFVc3u1KxZQXk/12l8pxvVZj8jnWgIvX3TEsZsoZ6w/D41BC
6xhd1LtUfJeg6bsnb+yBYV5+H8NnHOqkZuFtJBsUzS1+4qFALyFqcNVJhhbdB0k2hn6z9cG6wZBI
hB8OJAFj6xON517ug+qP1OJf6uK1rHsG0pxYXoT6xch+UowAmLY8V/4+ShcI8rx6DLYpPvJVhEGV
fj/RQD4+HY8CEDIrJcGjF+Rpk986lOFjZ/hvRA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11888)
`protect data_block
/O8DvoigFjWoWxIz2jJPtVuFDgx9XSAt7DXKcf6WXFldV1VxrtSgxMx8DDhmXW78Qy+ts41sakU0
RlrXpsTCWscwfUQcUEvgfUiucKA8J2ztkMFvNOApKFWA6qKSGT0wf6NE9z35bJEniQHGBv9slzVw
liiHYxcMGWrSAhVeEWHPIaTrE3HCMo+nBGsbqP3RBIBn3RoGrp0Ly8gz+iTu/xN3mEBm9J3iOVoY
sZOMMZUXBTTvar1SbJ9dpUMCukuwEgf6X8SN9lNd+II+BcelIQKUR2d0uxQLXbvjUoXfn5aIqZVR
IDzzfTlw1BR1sLElH6IP8YjO4PBxb9JeEJWd60afnkqRJcvId9NbQwBRvEgZL4ULeBDs6PZBuUn1
x2rmZBkjd4WNFRaehlycA8Dn8TOcEZthLYKVz5XSF31qEtgSwDLh4CEgSWGyYzPtNCCO4apR7pfV
KayK/CTyuxl39fVLP730Zwh8gNy5zsYMROLJIqhE4bvoFUkPGPO/rT/HrWdtCcb8muotPHslvf/h
p/8rUz1CxlVHnZoER4Sx2MMAyPETdchR8rno8ofyl1plCl0M9ilHBoQa3ANu6n5Avmc+i6clw9uH
gJQ4d1fuRUOwmabNlQScggvk74d4EqwqcJv7YyW8zfrX5q3/I8VP26gJi3rh8SXresuj50AEHJSm
32e+W9TuhXygXV7nKvcNtKX3XEJhZ94vD46gjRURy67AZU/nT3EnSLRa57qhvouj9vyVNUA4QBaj
R1HU5SxvzByQouHgV5Oqvmi93aChMOstgq8JFXBJ7wU3xNv9qiMyyx2pmrK29jxNFI7VqfGQIddv
5pPLFFsciwK1+4o6BXhp8esLmb9ciFy5lAzD9pimM0VVWEJt9VJDxpWNoQGkQdWvKAdKz+IyqUfQ
sQ7cEHLlu2Jk9FSp1jFLaF/z2e9wYsiOGA50I3vMwNgK/GfpNawPT/PNlOCHGnimp+euY3ufRvjp
DavSapQ7xRJzVYinURZT8REgNXYj3xew0rtON51895HW/kCT1KzZXzKso+3Z5mOd3szoXlFewudE
ndMxw1KcGc/2fHXcNr0zs9fix0UwBf0IV7XjkcApIc2wSHzqHloqICFj5QUM157UfdXnzpoHyRve
Z4oL3ed9tLCELPujjJL1I5JSytXStDcB0I2JY5dbYbOqe2wLXbsDNmcb6sBkK4Dt8nJPhVg5JAg4
YqFtd7FWltcBzJ++/NySngV61FrUCAr/wmkFMKwOAbjqkAxakMzOB2g7N3ZQoIjXMUekBlSURtqP
E2mxVmsJmyI3HU1qHD6BzDi1RxZ1nDm9nmmrLz656W0JXy1ThEOY5t4wHB00cTLb1M0mb9t8CHyX
UNFRnP3kamM0d3oNMgtPHp6nfH3HputWPQXACtDMBp3Zv4mUKiWl4NnVy0V5MJmsLA3om06rAs1x
EMXHLtSAp4/Be9mT21PaC5zuQo3nOQ6BKBz+//0LbJvNCewUfTvFL30VymsArPmmqYZ46SD5pHj9
gDOq/PACAfkE185+tdPGZoiPD3hQWhQFcHshZF9T1Ao61mIH/qZb6fA0AK4IsAndhd9dxRyAc6CA
dwA/r/SW6wivVwd1TaeCGMlNQu0qJMMzE4NTnmZHoXgWQSvzI7XHGyX4EWZrmmZCFqOi1+7/+NUr
tGAS6efENHWPZR0JrL41Fc27BVfe0OUWQK+Ex6cl0EdDXg8CG3GxlPsJSF03FnhYzevgWv1nHdxS
yFpTlB4rb72Pqj3R7Es4w2iB0M+OzVdDsO2Q/Fgk/WuAGbZID4giS5j3dDSVWyToBCoAdxd7R+lc
49jBntjCL+FrQ4tFYJbwImHsgYt6GgceOlV9QVNYdK5q8QJKJnEHeiGQ59qre/vIqYdDZgX+XzZb
7CNofMecvGN69YQ7lm0P5cWINwohx4ZdIgOKisl7CUG8/WphZ7wsOEM6IGNDEkDkC723sGfd8UQW
gEjCsTh+f5Wqe5OckJSyq/3yTNqp4G/QeNu8E+BT5T21LMB8l9K9biq22szIs2ynT8tI56K2v5dZ
HQz6nTFqUHBZkh9dIkVMR8xDuaB/Cjb68X+ceqAB9dGvoTyCSMSIni1OniHLmwzgqtYAznPT5Nwd
osQtY8R/dResfsd25QiJ4Av509vYvjLMX0vyHs5hLw3SqD3ASvT/M+QxCYrQKEe/9tord74+c9og
fTdGKbwbMUq7zZ+fo25t/mdCVGqsc9vph9c/inejWrQi5IyQolXvGheDpX77dgsCzNffJChIPEwf
cg3rGJW+eZffZA1IvwxtvbBXBBQx3FmnhlnNrpmhXjvPjJvtuuPVCDqVW0xct0bvO2uZuHdd9b38
YeE3IxBuX0kMhbyXP0ZtmgZ2qEvTzS9Z3XILxRpfvQ9bDopn91+J83k6mdQg5WlivJWFVCGxbxxL
LavevnQqXn67odvmAnZPRzwgLM7w++/JJep5YSGjwurJarMz+pkfIZf/7A/JY2kq3NN/1lalexzM
YmLPHFOkEPFkrNdPrgwptc1PN+bf46Z1On0cfePAP+3MRxNfPkbj25s8nFxtDDCcI+ePypChfVf6
t95tIuUaejpL/DLRfEOPGwujAoxffgtGLU0m32E0n+ksS8Wdgbuk/93B7g9UtdOv4TklBaR+AJZb
1/1Dj/2UE+bJWH/DNtiYyKWH55nscuHo+DCLRpE44WQzJ7JpGNMmzS5Agcb2SrAMkWfJWrbA7+yy
mzynVN98M+o8BN3nPH2svwkorCHAYPRMIvCXG38OBU/o5PjpH+TD+l+3FVvok3sBWQoIoPmBKcNq
bzAIUU7uliG3fGmbx2aRz+0M8NIMZjWxiY+nSMCr8kE6p23Sk5cgatjqbpdsedeKniOcMhxQcM+0
kkly8TFNOCYCYmGZejqYnHAuzECoPRwfNf3jGUXF4hqvs7bbuf5l7xtiQ/N/p2haCUB1KtCrxtjv
upaQfZkTlg/TqPCkHeW8s8L9eXKQBHHrZ67ADHMx1vqsS9+LGTT9MvgMtU/hqw8PVKC7pYodQCCD
Y7DV9XJxeAl3yEThlg/17EdIPvRPgMaVzYwWaZmGk05JGi0TU+b28/JuriU+/yczTHCy3bvw32p4
CPtZRw3kyLPCvIwR0A1n3RJqa9o7Az1+3tE4s+ASvyfLt8/kpzct9s0ZFJ1SP12JeeLqvsbe2Nsv
TDqUePGYc2+DvdV/QAzcYZglN/p6eNPxurHu62PuVnI7Fv3q7q7K4i+y92Qt8/kDXe98/PIBcq2y
MbmfGBjubG9RGFv23kUF2ECxDScHpYI3jFzqiSQBOPWS+gxV28ks/io429zbBdBh17XfoGQfPa6h
hEkKF10xZ6XnpJTOqrwWl/c3pOPiFnouhWHfpZwPikAKGkz9/9rLU23XivKZPCTjBZQZAbjzDaTc
GnEPNo05/77i3sDDStzHMySQ9fOezRE7Epy+PnmjAEMIzvvYgvynDDpsPGNRyOWDpgcQXgoIusJN
kWXQufpzhYoUrRtbIf+YQlZpXIRoHEzv0+7DQGE/klq0c9unQ6d0dbe3PIuW2pT9iY7Q1qcwxnDa
x8RtQbciZyROZShEzi3nu2H2sI6529b8Zsc+tnIcM4AHQdTgk5UovrPZfmRIuBNk6p9fI3tD5f7x
EyoTcKaeu/02vXSR+yykThsYDo2cbOMME1ZqjfcwgQtE6XQcLN1MxyD6PLQt766FpjfzRB74zXyP
6X3rX1h18gE6WYRCjh7h2CEpYXSQ5k6MHVgAgH32W+JEJapI09QpBe2sDzCnRMuDtpmSiaBLyhdV
2D1EZznFVcAE1SEPgfZj8Ong5hbMhrOfRq/qQaPDuXt2YN/HQRFrAqiTF4PNcWlX11AIA3zIYY1d
zTWED/VCRm/3ewS6Eu2jzvJVDQGhLG6Ou/m53ESt8GY1ggTi9Fayg7BcpAdZaJLVQ4RRTT5s73mD
PDocQHGnElM1YfdTEUq40DFpVKE8RgLv4briVbOfgc1E3HQGCvnfDKkuwXXCB4S44gk1nwFdKeKd
eKzx2xemh2q5EmgwEeWX0GvHT5e4SlIMpNvjwU01ISEMZLyWiSOm4NLteOKneCseuEemmXjoSt+6
anWR5w5H6SZ4tVjygpclaGsEkRfRdRe5JLzSUetOJblLVWDUZbcRoNlmIJ9xEDhXpqbg4Lku4jok
11nBZZrnLmN9qtoLRwBj3H92ZaC2kti7MQFCBc+GBGYgQte3Q0wjTBenK6//ikaexBz15w5yQxmn
Ltr0T8ZbLIi0rcxmfqFuu/5xY9xTiT0QcQ0wAABf0UkRJTi/xSznqwST8NibTGKRzDZtSQ9IyYgJ
HW9CzpgV5Fqd3cNooeE6NjHSNuBXTX3BO1hc+lSws6L9IAkcdglxBaqXxfys+xlnFey1IrBArWZA
Bvq5Fti0qN8wcIp03t5IiYjIQnH/eKVyjddpYAAzRPtkhHv/UHVbjSq8A7Dc4Sq98UUKtok4a4nN
Q1Z5ivNWvL8hfMqY5bH4zRm8qcrmSzh7nOq8mCZ8s/6165NuncT89kYL2CQ63G3wyHzNo4Tqu2Cp
lV9eF5z82UzFYNOAKq6LNSzv0Zi7HPncUcQhguhi7YCxqwRLbVV8dE3UJtOwNymyGLPWRVZnej2H
gCgnxVfC1EzQXMBP5UN0TylkB/bCTp6A4hdObqWdhLg3O25vUkA+LtkjA5KbYPHK9jIBGEOlYOaK
5EAxKx4yyFfAjdn6TRPMW1IZCoQwka5CY9xAhrROgxdxJAYeQLdf7S3Zhhqg0l5MHUgvBRLcHS48
nrwmaQsba5yaNMCcrOuYe+8eUQE/xhbz73V5uAf4HZj6tO0wukEELnrMatJ7/iBbf5yP30e62n5t
fkw8wTrrC3uYqI41IbXVRdnmCML+RyMV35h9NeZFyt0UIkqqi7C4xmm/RV/Nks71Xdb8ZfRgR34h
U7fc0CQmT35pBBAfopVjdN56+yR5Xb6+BCqtz4n30yHviEdLvA+axNGcoUTb4bsJgubxE5H6IVdU
4gdEfF0IdlKltepETrn3/ypkJobB1mjN5r4qFvZhod2LPoUjnva+5/9yqYRP6hM8xnTYQoMiBn+0
kkyHsux0b3VRYiCHCmtEu/WMsqN8/fLW+Ec+cu38KBzrR2h8TCoZFD5csAYUt8XWL+Mun00Nl/w0
jVuJRtEbDTgFmH4hYetfqLq55G206blTZ8luI/hNFHHQZ3ObaPAbe+/bwkaS+gRHU4Ftib+BtxpH
qZS1OugjtHMyk6hx0qQqPWRzwWY4a2LSaaY9wQqvedzogSK0Ut2R9YBrax54fZPwE491Ar2GhjJh
s+gdoOnuneU/79v7E7USrCfueZpENHYIo/FEN96Ry0NDdLx79ucKSo2gM9Ce+8swQF2THYviXBfe
no1MhaASk+wvyRitku0QQA/98/DOr6fBQhNGF/UaaAuCAWoxYvFCdahHi5tbNOhvJkpEoDGASau7
m3PuUVrdJZEUzm0COlaOr3HOIKZp2cgNmz8trg2gkXV2W/F9k7/0r48AOgN8yEzmKLpxJk2SqPl0
333GQR7f3F6pUadAfMwJdXjWZh8iY6J4e3lB3LtNULOVmOJy1rYf5hJdlxXCicaXWqTXuS8d0pz8
x6zgdiBfRw8fNr6u/kmlwao80RJ0uiZz/v/oes28KdyZ24ouV3TzLwbZpI0M3U++nra5Xonnniz0
RG+Q6ifWjivAmjl2zG7ykk/9YdGYebRmigLKZBZ31IqQSrskKO5F0heCh0gmBQlqMttBgcEtSAtP
Yfl4k3a7dlkwldIU9tLu1+bLq2S8GC7OMCUjFe7XvO5o2BHI6e2CtwuTgnpRoOAcAyQZbfCE5LHN
H3vYAqTEfU+k55UkS9rviMtVWLUW4tYQQFMroCJruoMOQg35f41RkzTlA6IWBb2/ACbJeS996Zqt
Rthj+OuIaO6c4oS2dXLHBWDDmhP3PSQ1Y7PhtkMMWH+28f95Nws/DiCrsB8AqxPHz8dO5b1Eg6C4
uYltBYej2QN6G/YKggxoy9f1YEY3yhD6UZIlomjOaNBFybwPkwA/sYx4uQETtTk8vxIdooxHOKGw
A+50wMyEGvPZeBf5uYLt1PpuiQ5k3kcXOwf36Knle9nowENaP8AUXpMYiyIS7M99AOKXT4aZ7NtL
NMxWqSkdUsJsr/9PXgxtoybXTWhK7GfZAyLpnpeuEbYMCph6sby2/n8McvFBNHmO38YpDy0Ak57K
QhuG/xsxNcyoUuBnkj5cWU1WBUJMc465TBeTer3IuDBOzplPVO9rfCbq0IP7hMCj7BZdw0lHVDwE
gfCRFbUviiyXfZnmN9Id+nNsJ+lSG7VtdvX7wqVVEiSXf0goL72t7uQpGA7jtY7DB+PITiNdgc56
LGFdM1Qh0WJiK76ZvAJbdIOjgIhDCtquyC6ViYbJnBoKMP3g0SC2ZTt0gp++yogdZoO4iA8+0E89
/E4Q6BDsn6sNqtE2XFdqDDU6xAfox6fI+TYTqhHaEcZunPVzaX6GPrHyzDACPXfILnABsx0+TSDQ
mqTrj3GCCL1OVRCNxK537gbdkrM12y/O8LuzyqU4DRObIlCns2hITG2jfketwkzWTW1NCljrI+XJ
gE58VL/uzSZDKJJ//e7MtuaSei9GwXJ41EEls1iH6AXtEvuKY6OwgeYzNWAlbwESKPduvLTh00m3
0/uic9oOzxqYI4IJKnBAQyRtvUOOMKgLViEVJToUZsJYVdZZ8I2KNPUKDEd26AciZLMnZVkXxtHU
EAQ564bFxyF/vZv2boeUoWRXszznqvajE++iYVrE+mPYqBV07UG+AzhFo0SDeADzs4B8yrhD+RCI
nQZ6JT356PRFnsAkRU2TED7JOuhdRBX9iaCc1EZ+Wo9TwxBO+SAyLy0A3t4bl8Jg5e5MjoTuPxBI
++n9A3Iufc73B5NrDEh0vy0ie97LodwQJe2ZOPwnXNpzU2LjQ/BvrUbVOj2DVJH9Qk5AmEDP5FaB
wrpoNf61j2bkUHjdGV5Xl/JW6lt+WKoG6/ZvrwkbDwCPFEXQZX6xr6FuqtPl1ICMosX13ybNV0dP
n7eU2l4u/lvIukm08AgoWONDkfPHu0xpMSIpduMmTYh6lZZ65fdMY1xGxTJsfsCFquSpzI5B9QAD
RVAHQUZ7bi2PDImHRsNwfWJom4VNqrIkkva5Gy+rB/InzEpmLL9Z0HcH9JByjG72byvgSbWRrMKK
eXGjXtfQPZuN119SGKaQXTLSgsf54Mh8Qy8Xi7rD6xlpVxmyotJhQu6l7F/7Szfn0i3MA0fSDe9e
bPbcQFgFDjVNzBSd8UmSCF0UV4mzojSzeyXIme4NLEHoyOa5/iHQ+Snxe674EPEtSZ3Ib0C8K+3C
ZF+GSNF1OUOwYnYkc/hu56IB+jGveV/MiiNwG0WJdFAFCW5JuNjOLnjcoyLLQC1Bew2wheldrEuP
REI9i5Gs1HQ4Qo/8jpdsa8HeDZetalVdrnYcwrOK5CMKpno6NO5ZmWMnSnd9W1/kmvU77v2ioPbC
kHApx49wNU6qJ/3WNHssnzmrSt9yZ3aAo20+gwEkeGih2xzqHaSJVwmel9dogU12veB6s/ororqA
jw2hbqLFrldNe6i65irdmaZv0ruR3lsRIFcOn5ws+UaJAY+7fvF8oFe1yoykG4NswnhDDnbHDCvS
tA1shK04c9I3Di+76NfIGZbRsPe9hENLhQ9leAOW56V3cGTy5zHrP/Jnh4oQ4afxZR29bqvdebg+
qacm+ZQqWDeY2ztq2xYy5Td+Lh9BdtiwX6gxboqChopoTNu/RXVsZcQFS5AVbPsGmHSSESK1ksyl
kPipWBfFYt2xC59kGDQoOUCFeV5sBbVE2q7lqJcsGdSCZl6FUNKp2+g05JIt7oczXvUqu8JJbBq8
a6KqC+BzQm/bQm/XxkSBJ6wawgt36SRKyu5HpWwV2GZFUdE5HuWtVVoqd2RjKqimoOIVWujELfWy
bQ/0rmmU/w+ZU4XYF4wWYsjyTUdmVKwncktifiS7pqebN3EoXGwebmGh06F+Gp7XqB/sBUgqiKJy
BimMVCt+w0LgZHd7rIM+ujMMJRX8LyiHRs51K2gA60Qp//ZLQgv1ipFb6dlsZv6N+Yx6VG/cMt+7
7jELNwN/d60694RIWPjLfjKvHYOWaC9lhmcdo9gspIKX+o8aGJfXT8Xc2AM1RMxdqxr+J74g6Khw
zJJgOe3IvZ7xvHVoP65DAnDNySCUSqKVGhhmrh1oQ5uMsGNZc/AhUVl3EEcZ6Zg/3WvDXXlWzkBF
WNz9cw2ZdmbUrJnZc91NZ5Ewt82tBYC6ZEDt/aw9Iol5ke9LKTJJnih+uDbqaAMN06DkHlI576JO
nKn3aaMOXS1AIflZFDbEkglOMlQ6mYhNC1bH52Y6Wk/Vs25v/ZNHufZYgkyWMI0XXfxkHKZjZ/DV
65625109Hc1ni0eADy0iEE1eDlnAzQMWqK2yI5fMNtWaN/N8wMPQGn4oqnKWTUd9MRnSyzqCr+Ve
hY3L51926eGPmYgj0FizNCjXieoN1zielNfGMVocDEegX1Q12AbCqBNxS2He5FXhUiPBudU8tDr/
9mc3TOqr2qwBbce2CLDzHnIrFkHCPZNWGD+lXpx8iN5GDMLujwZI3KWsYif/1wPpc0tCOGG+T+PL
37W7AW2o4yJIQUah3okpcuB24EHHQ3CCKe2YOl11kBfRwz42VQHk+9YyB3VXNRtuQxfIP5QHsAaM
rXfi/XtQREZTN5EQy6EZ8SkeVHyXotXczrBo0DPiBrHJvS3nIM8buFXEFEWXYStB+Y9dPVPSmVLb
+S0HqaQ6La2nAXA1zwh4w1eSgn3lkRxHiIHIilm8YuxlKav0iilyNGRGGJyE29mIna1H/s0uNnJq
gMyQC82B+G+w2nFvhvWmwk9J/xvcgmsQjTaZxxZIWz57xD4+mLuDwMC7OV3oIiQ5g3oCMvaCxK/i
hgDpO8KrsAa1twyXOsd91MuXcsv0pBsgcAsTe8Ev32wYZUYRpHsh66VraZchPsm6TXz2LEyxqPy3
pbDj3qMgikHAogBC5HneVjvZqBUFI0+EHh04M8x34R4FoaIeGdNtsz08oz7gBEB6HlT3X57yjx9F
B9XXJgAnaKME0NoiOJfLF9z9+41Z6aBw70+9bveEV5MCx+N6vmTzoSEXDhrPrfGeh+A4xesFad0l
WiNnjsjD/TKBlOzboS3hr9Tzf180E5hIeu3617W5He7XU9fA+gkWQVKHqRa0JEKVb6FG5lsPUH7p
XukXztEpLLMDd7IreiaLoFRnBcWWIwCH9+lhXz48T6g89S6VQ+LaCPz5sY87CTowR62AiUNcJBRO
kkqlG4lIpvbIGqsQAC00nifHvWONfv4p+I8Fy/szDGvpd7k5oTuDu3AMgno91ev2z4LR8ho1ZfHh
8GD8K4Manf6JrkltwUr7JA21/a2dNTxzndNQHRo/BuLu4XvWC6rItb2cjTcCfYjiWabf139ROmUm
DT66/enD7dR6NndLxG99LEobMfPg05ozCMfo3YSO1DRwI0T9B6XwXPpI2Jm+SzMKCF3RGII4DYCe
wDesDNcBJ719y/p+WE1UgcL+yfnfplTmArOllLoAG/ACdHESggRgJK0mYw2lQLWS+0nNEHIscL+d
QaywrHNoosmfkAxXd0HML96ATbIqdcnC/HlhK0zYhOV4rVo40oEVhcUOusEa4zuGfsoTTFmh1jZ8
lDOG+8I3Rn7ed7NE1SmhfBd2T5PYQ4BWXIeJNRHoHZcyoU7GE/lC3qM1rtvcyDz//jJ6oge7rkRG
gPuwxgmWJLuBdfWr4+0oOn8AOwT1NCPN2QiVa0noi/dNFubVZeHf4rLdsTpvAoZ5EYGiPcPts0ws
L8HGuAXK6zFpxqfScnei0AP9GDU7Mud/6H9GuADOtZE80udKSC3y8bolZUOrirK1zwCrfwEEoqUV
r509SPyfLLdggztBq0BFhAI7bk9kNMMjWDI0dBuUzxkRnKMfEA7mwp3kxnj4lsadihNSpqjJKxKb
FB67NOQAgJ1/L6pgYKWGTiE4HdTJRde51mmHeZc0W22vFnK3pkDPQK5+RSCgd98XFTHOt8oQPHIL
FIZAwE3WAdP9I+vk+JNqVWwrlczbWEz8UunoS/5nyHbZ0fBsGwHZ9ucmj8Rpj4E9MyYl3zu7H6Vv
KWoy1cmBTLehdjosfWOZBKtZrlXbalHw5G67bL8FZMMv2qaqdXn/D33lA4OqRLDoKdzqoohTsX3x
oy2CBNYrbr1USAKAgGVXSxqahYqtet6z6/d3zd3zNF+8jk9ita3Qj5xxn4z8hAj4TG7h/4DlYOPW
6M/WibdeqWiZpK0r99o7qctrc9baynHrJwEK6G5QH2gp/zUGA0G6gEQUnbIEvQS7U3yaDHCWkR0v
m/KJRtnxyj0oEneIPlkDXzdoVYhS4bYYKtvZD49deiWifJyrteGKCb32WWVoU52illDW3fUavlrO
MadV0cRh/64v5i4vZKN0dVjflML10Ae9fxYiRWa0Jr6HR3jUPp67EHcmtPOdK4DvFo4s8/UxHdn3
kyXc/Nrvuq84hnlrhKIx0xY0jFhw1hBsYzpYXBGiVaXafiWRv9OoKvASJpCrvGNcNNFxaS9Ma7Wh
RX/4nbxPO6+iRhg8C7QNA1T9NoCn7CscIdMCbG5gNWjiYpvdB8g7m0N33Pwz0Nx1g2g3HQWtSbc+
wboDaAAXXZxvxmXmm4Vj0WWrsQUEXSGKMQfeAKV6BGpeQDzP5rRzgghzIFnifQLmRh3wTMCAdEE6
tX1V4o/dN8qer55+cke4GPiKwE815OVYJfPOySdr/4zIdtAtZDxbRXEkmCg7gF8rbDpGBBwhOKu6
qne6sFwCpdEahPk4LD2nl8jGTPN01pQS2pasWCV+KbOCU4wsBjB4wZ82S+QR31L831QrxZSGGSis
Vahfv15Svn4fgaPcqtG7plzfSCg9AZUFlsbe5R6xEGgpCWO8d/1FTcVL0ZIjtB8t6k4emZmbljL0
LOunp1s8tppbu1BdHXDOrSpol9rMFoR0qwHwP815zUF1DS5LJuSSHR22/A/zod8p8gIA5NL8PfLf
i54Syj4DA5R5MUswPL9emkeF0CzWwCepzJzLSFqkckYayE4VIZ4vyOkPGCl5LLcnfEqJiG2p/kRh
KxZvXJrKyLDgIfQ4vbeRf4a5/GtM92t5ZOkWWPTYoobkgkuufJeEm/JBAkHh+qvYMmEpez/zODu8
QFkggsacrsS8P2+e58l5IT84BUkDj4vR4R30S1tdtsSY440gXrghHG0wU/4F9XIhWCCBG2RsjMpS
T5kqBwnmbLEfkOcgGDN2nAi5vlfYtCrdPHkT8vo0olIm+4uyD2PLudb9D09/d0bbtSmSroJRZ9pM
35syP0VFIaty8boOM3ztXHis+LqTy0m48+Pv7Xgt+zVEspKhcO+wJGgXTuX5jS2hSixH9gfiGzyN
rK7mmuWSCONmiziDNagxRlcHN2r1Yg/pPPTBDyOtkRdRGeFNEIy4U60hTj1cQiI6EdIdazjc5qzb
DWNRWQaDlH1rMbSD9nYCLnUyeyUQBdpjGo+4H9sYlpW+4P82ClqDKlJQgTHCATryCErz2wFv0Jjv
UnPKjffYm613P5ETqaoxFFerWA61KS3q9SiG4GHRj6kn7oxrAcprjgqu0HnCZCMc7VNd5QRQ6HAz
QHtQP0kCHQXEwqUqLFbhHtTvePswsmw6DN6rLLNT4PFuspWb2Ug79Kg18+4tJXbGrVuxFtUXSyxb
fB4COG5DJon1OEWt7hmYseZqCiZ3STUBqf4THjVkOu50UeYc04IRYOGvnhcO7EzfuobDRiRe0XlO
IrRIwaY4w44jj+yRJ5tO2SrbmCcfhr4zJSiJ8lHDzEbARRgHTcBwQtnsOpRuAl9fGTN9vRcKMWWn
nFEUeIXAWbtEw0XbKNy4kk4Wu7nD6Ijgksqy8EPT03aLZfsiT1funLxeKRJPMN27pz09mF6EifVP
+tOYHUAxaZyCUsQGA1Ts0GADKcFZFOBxyYyEQp6E7rYq8FvOyBs+nAqPzO+drk5XJiWFqfUYrOqg
dvXTgc2EeLpTbQ0DWs1+t3IwC2Lic/HvRy9HaEocTFNcECiU3AHl7jS4o18RQVIzyMoEX/NuEQAT
oxTnG/0oKNkDf4MF6PHbdyG28RTxlUELNjI8vlpoHx8HJ57yom6ogoejguX8CNwXYCFfEt6cIxJw
506Gbi9Q1t/fcggO5nwks2J+MsZL1KnM1SqeyHLmYa2Wnd9X8jradRkT6ht3VMnapWBc4u51pjVA
tSDOvSxH6J1F+sVQnizJRL3m9KF6uk8MHJtLt1af/mh/cf2gH64DqyX5HCAuxgRv73Wgf97AODvA
gJudxOKLmjRswG5JSjO0bJjNgU4GT+mo5mqdQ3fqyjznyvX8UwNGfrGmIMu1on3DpSl4/s22YFQV
ohUQvEjAGOn4eyIZL3edJtKteJNXF3y+/g0NN4QSgEs+YOcEp6j9QC7UvmNUeRmH5DpAkMffe/fs
1UNG/cyxrcjuZqT9CxW4rhK80kp/Vsz/BfjJk4kIXg58F6pezpx2vzPw0mtS1q/DtbFKQWDx9bBw
5yAGajfW5yAUv6DW/fhJDefAMpx+Cj84bpHsDSpPycO0Lss8i8XlTp5e0daiCinz7Muwpc5x96Cq
Gn8Fb3m9eDkEi3iEAkItiHUGBPbV7WmwO0XhZ53S8FOk/D4Y3GvZNgdF+sXEWhP09se59TUZDO2n
4emxmtNlnzJMqnV2OKienHZl0mDAf5oU3Pq4GaXg1NhtzEqXVTQZin2vUWLFUI17pyMLivM9Q6SG
BkijrMWha+kpA+YE8vuxJLDuOz2nta6ZPYSpqeiWJE8RUGn62PQIBKLGeJuvu8kFI7RHD/kNZp45
KkO1odT5mbVP3EBzWOSXkv23+90sBlqnJNwq+vDTF8azpKg7WtRH3dDlfBB3+zGrZZfq3H5YrG2l
y+9+uYTv8pRNKSjsxVDUspTItp6cdx/iW64HC8fy0iAQnMgv7VFbzbzUXCAztBwsoa3VwzltOzCc
x11z6OtJPwZF8emluhIw9XU6jhd2dhCnr5pbBTkdCt0voxJtVxOxR7AdTPtpESJ33awWx8u6tjFe
9UAD3IZOrP7gkKpYTZdsilOUkdXVWxgesQCrmJKqGy06bJxFe35UHGWLRiTsJFXNhUZyU9nakYMZ
p/FBHIlFGeLdGo9sO5UB8sUKGCB3tbF6hinwcupEpmzVGn5QYmDEBv+9ao3cDWeEQLYst6mvTgxD
v5FDeCUbC0OOg5r9/4o904+QIylpEaxu/l7YR7280OWDgYMG60PRmvR68Rtc52A/f8EMPNLVN6zJ
Uca1iNfxbgna5ELd1qGVfHMLgKEN/p0YhxWv1Elx//BaZkDp6CsT/InUYTsI8b99k31Ig6dzvUHq
BJ+CnLpDTGdABK8lTFTApTFHAeHsJCi/cjS43XpIRr1iaEsa2Z5UJtmcjBewfklOlodOrpCBv1kg
4s7dYi6tEyvsanz7+fZ8IldsKpuulKcrV3rUOJDyXwpjpBKQleMhg6IauW/b5Zkuywv6lDny2p5f
eqpEuA5WisUsf8wez+8mp09uBFqU/PvOskHWJlCFso9CBfkqj6LvFkjIta9SAUiy7rzBzDacFS3u
ZcIisRJyxa7NrPLF1gLlYEY4Z0sHAEBH6u/xn06cukqIj//kvtBFoh4rx6UV/xz5fwlFPHuwYces
W5+9gLsgSLJiHBIiOwIIBnFw3ZsBkHXDfvEZW69SGeA0PLFnk5GgdsqRpC76v/u4WvbB7tBj7yoW
66Q4jSbsFIk5IJ81ZGBsvowWrNz2kuoqZ93ftERr4HyeuJ/xjsttNkX0i0HDtC+5u204oHjxr80i
tLeXyhe0oV/wnT/q9eoRjgVylw5a4dhLHXKx4tvSKItPpxe35NF/drt9h7PRNZUzgaeA/HPEsHcw
G/zxmuwoqRp2Eh200r6GbwB0K/V+ljYnwrm4dYbmlpdWT2MpjUmkox3TIUloIH31B8RG/U5OzTqa
NigEJxB+Y8Hb9ycyEEd0rwKzh4VNJ/wvlcP8+PLcFnXiCFrEpgRZqIVSgUby3x5eQxWYzH1jZZy0
430unej4YF7YxZPSK91xTZC0hNmYRjG2I/chOAH2+cD5WW792kXLUE0KaPMwYrVOTep/M1HgrWep
YrrHKnqq+OMwjW4d6uMPfU6gxXivjxnPrBPysoTSDnWhL6YL4pdcs0b1NfLy05GgWDjh1M2GuKFS
Pl/AVIxBQgQDbb3UPyvi+VAmMjtR9iVkRZNHN9WSHXDwqF8rbBTqCp7iiQwPHwvdsQhdr+yrB2Zb
q5RDZGcYinwMsOfBmxY+VIhyrk0d5x79F4BdD3P9Jnm5jpTKzPxBHZ0vy46Yrp9NqpOtUjx5cptk
g1U8Xd2Txbo+baFHtD2NcCJvw4JfSO/kpm5+L8axPVEZaor1tQ4w2qzG+kYN60GWAEpx9AM9MaN/
m8s4Fh6UISE+aCmpCW28zexuPWplwKDePSHdQy7wX51W50zP+Fdima3D3PnERqw0IvM1Vw/RIoXw
eBmktBYHsBkq/Gh1WZJu638ELY6Nr5amX7PoZ7tvdBAIT9JDwcWdmsqzq9+bJC3loVRuRtbDOWdT
iahiidjqH4A3ch/76DLE1HQf4H5W1lBxzrmiWzZXpWHJKUrIVikgmcAS0iebXD8MSBc06FwuYfJW
6Iv2as+sbwgv2qU+ua3D3+n689vNer9oEjy+3qk+Mlsy/GEMTl2t1NEF16ANmtbFZAbQJxvkpFtg
TBlRptcf5PHo5FGRS6ACO3HaUyg6OsSOINcyaMdDEvdK0BYc4PtfiiRlL0eziRACdZ4A4Wq+K7mq
KW8/Wo3kORwSYxlk6WZJQouUsQVY2FKbuZa9Qt/9SxP1yHnp+1j0n3XtHJ937APRAtM/HRs1iWYW
D0l7O1fJo0VCmt4lZaUhx1AhZ7cHVgN2LpUT5/LAPPcnh9bi6VysnDeSx6lY7Mp4P+tYza2DZ5wJ
nLovocKfTU+5Iul9Bw+blcPPHAN0lF6hxKBC5rewkXNLRMNdhcfLxCDgBYQFfKAOeZFIRo72YwEo
TaH85N2maKrBQYHY3yFsq/xkfYUbeH+gcOaU4wINlN5+0np2lqBEmKKaAUiiBeVubdSLSdbwCLEC
QGZNk0u3BFBYCpA1ornB9mSs9oydttMEYxXNz5pFByW4WD4kF7sQjfYCvF2sfYsba5Mkdvy9Bbl7
PhBlfeVz5AYgq2zcGyD3Jr4stH/ZF5BnXTrFDPCqMDzLuz8oXDyYRY4GCRDwi4FhyqEJbRFIN3kj
hoqUEUdBM78RRe5KBUpShH+IYJv+K8v/YMVdqYTGw9Yqevaihvv+XY5WZz7UbwI8Ji3Ir6cx4k6/
4xppnuTq1B0F1TOjLD9UYETEMpisltuUoQCfwrNhUOisVKuAglVLTqdvrWg5xfINkc9x8o6WW/v3
fwKujiVxh+04HUyXWau9imNOd0/CcOKnY8xD/zq8kGPZSLFepiFfIpgQGT+Cnn51u0ofmduoyCg7
A+kUQctPE1/UdxSQcSOO5irfoCD/2FRImkee4q1B2VYAXZSfEAHRMj5f8kM96kuhIoZR4Yq8sH8E
zAX23BeFl4yBERGqMYk9K7OECBY8ILvFjhRkbvcUa6tBE21YV3vvaBm5FEiICecoXBoOsk+X8NXT
UQwwaM68ZSvL03Wzz3u9IYIHdSw7sINCOTn1VbtGT+kLhN6+ZPHDTOz1gX1164SUot2nfNhtvZ34
fRGWhdZD2nWMsSYX6MnkV7hc4A5VnYul3Gz98w5hCi4=
`protect end_protected

