

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iEtOB5S3Q/0nxxj3yhZWc1e9CYVNx9kxE38Uvw9Q5GTpbeWA/PaP7MHi1hZ25jWcWTCQq2m6lqXe
j4/ejpW9UA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Xuau91ineWkILAnXNctj7ghjv8v9lVNvmGeO8/qKPRA098IIoEEWbPkQsDw9y8PN0Kc6j93b9RA3
24AkaGw7vS3twv084InDNHpEnlN63djkx5ZcyOiUohe4xecSmu6QA9TFBRDs0Woq2jQD5/qd0oJL
/BaRHEN9wihMkCnRmi4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DukDx60lt5tRoBa9fYOjxQXcMx39PTzSzi3mfBKPNtGRH42SBSoh47iSUDQLozXc9RVtQC3PW07a
TdEl+U9LI0QpSHNQLVojqhahZCfYOg99dtV1mWPojzxtpV99k2zYX2J3PXN/YbIzV8ZxTpLcq1Jp
CAIcrPJ/34KYVzvzXFRsvxEfk+CxS8lIGg/nVz9ZI/SFfi31TG5Gc9nsiydQV6NxDLfMTIZ9geQt
WjMt/ZdcVbixfIDM01Blr6PmvrTG06LX8uxL31TQuw5SZfsZBAh/PoXSzsMleljAYXIhMhdSUOnh
qfkHi0I/YHOxbZGvwoECi6yzPk1O8e4p+mbfJg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfFouWl9C67kV59ngW+xbX0i0eu6h0roaptqFtm5oV4WYkqMJEDqBwmHay9e7sJ9CO+K40RDFIJe
/eeImbz2XS0Q6PwgmMgPAHRoOg4fHkGIAEugmb7hj+mXvk7iQo09CaB7HocKsvGcx4nu5U5a1pLQ
6UjYczksNjCCieDaJQc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RNy6OyrkxjF2nMK7NTVKf+mkYRQZVhnkvdhxFI69h+pJImlNAm3GMG9cNkr/rYPBFr0KpngtSqYa
zub6qdQpsLCoZ7qDFdEc1+wws1xQHHeB7VAyyByyPc8Chu9XZcfd6cEAYC55a9lNvtmKoAjppEfF
hj3OtTTwZQDicoWmteMIzi2n5YcjhwpDSzFHpmKq+NQje013CABovpP0/TVMHv74ZpkyX30HW4tb
0iH2SzLvUD7U/AR0ul2kht6wcMaLE9E6bQipSYn1DEnfUpMfQgGpPJCWjykHayljMFWfI9ucuNXK
1XTo7EI77uCstdWwv1uP3ZSQ8pFNDP7NXG8mpg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9552)
`protect data_block
LOXUn6JsNXcyzOeWspbnGFiQ9mJvLX3ZkWDx4KrDTRdqlFo6sLRdL4u3oS1GnbunopFVSQu7VNjk
vUmKVclR2xuTceEnEjA9eExzHI49B8pPjDff7zM3LnhiJkH4xjedPYNt9Q03022bPtOcC2QN6iUv
wmYOsY/0fh0Ra7v1IeW3Tc0SBlU9s1tg84Pj7tSgG+WeHcRhZR+CsCvnc1lBS3fPBZYsRdrqciL1
KG9jOudd+2hxaOpgPQ0BwTRLU4pwTAeTG9pazFEyw/A2b6z6/1nuF1NT1dY6lmBKgTMhef2TXioR
9JKxzCMLV8uPmRvOMJ4Qg9+36mHt0JcVrznhWzZVHA9vVhgGHXAuNj/tvnXdePLOJbFexm+0+MPL
gEUqLQrOxVYqyOnjshDSzhT/0XxRev/ZIpvENt8hruucuXH999mk/hfoLZF2Wh83oq9zUv/EYc4S
+Jpl6d60xZeBX4+3OQKxfCsjT2+YZnQn4sj1nmSqSHiyMTkkwLQcA+P/ek6cok0GFuGgSJr/G8Ox
SxXkWF9rt5NE6N1LHUYSECsUt/nhWxoeSwdgPj44My32HMFFVBC3d5SGXzoSQHBHjknBM1IMZKGw
bjPC1m5tRgLiScK9OdPIB2SugWWzlFOcV2gSB+r6jWghNqEnn+f4PC56CO4ANWxe3kqJWdNtyAvR
bE66bM/kI5+rwBAEgP9cwhHTeNpfhYbZVHP2G4ryjj7PhciMvz8ZHxVkvAQ1AKG/i9zjihh9pQpw
t3d+vWQ5tE6gPy14pnIKjZLndDgR43ph4W/MrukLoOhCapedP0qvgpLks9Ns7HdhGwe+qCCVcpIi
u02kegcJgY1ostBV/W1l+x+XBYGVG2mqCty9otdC1fvFbnv1eaVFaPossYkaGIOUmZKjpMFIPuqX
TzUbzxvCPE6WmSYVqmhiwh+KlLSz8XXbdLCnMpWpDmMNdED0V3acDLu2bn7bZvttM0IP6/alfmLs
meILis4NmlJ83REOwVVwXbZNsSoElZCa/XqRWjs8B7VCrTRyi9uUyU3b5gQ8sJj63gkJ4xWzN13v
clEUwalwsH0Bn7sNrlmIXXqV1QTGtzEw4UT6Qjkl4X2L1/3ScyV/JJWWavzJOlUn9IAYkl3tNdrv
KQRvxtZkr82T5ddafrjB5dX29h9FVP+QJOi99F1rPcdQBMOF8Y2LT+gaylJugcphuw+uAL4yNNTR
G2GkoX9NAR/ka/aMk7SDZs5iYLuAJWQZqTvT/HsQ/zXZ0ghr3pZdZ1ffxxMAU0Aevs0EeNA8YOdx
6JyydwGRID71pVnP2ITlykah0WqDBLfHB7HgFTchOse9ow/hehVph58y2QCXi8UWTruSSL4KqOWv
Mf2gdkewkucWQ6tMJMKjKtLRMccITZn8W0f1svKbgDe87EQtPNgoi3x/y/tgn0YStFUZqYQQOB7J
/VYActQ87LzK2KczkK1MK81ossTzU0x0+BHitaEie4VwvL/Ur8PHM7Yg7VFAIiU/WylJSMcI1g3n
y7I9PA3dypelhNNPuONjzbkzGh0hv2DimYLsyiCO6RhUTtqcGFQip4x03ajuBhVyPBkWIhXBFpFk
DyGOP65Rw4Yi4wZTw+7/pgpqAul5B7gGyybBQpbdfPEOuGkYzLkG+GJaaqh8QSidXZvb1FmDvLUj
htnGKG/s6iVxSNG3UIarw9o6tkEqQ/ZFwSqFuE4RG3gx6pfwarvPzgoBIZcsXmeHVsAwtP17dUgL
VQBGS8u2n+/zDuFTu0jTubPCZOGpUvpuyw6ehS97RNinpCmGtkHNdRoJImQ1WWCghlt0F5F15Buk
Mh0LdhnuobxwIpuU2EU/EshkYzeT7ZymfwrUm82OpAQClthGgNMPfIZmEDiWBeyztyIb6wVbdanQ
kY40sxtZ7Q9JGwGAbQfd2aw+/P3YRtaXhc0iWr1+H4Lq4Qr+lmUEdOXjxHDN1F6X/4YjFXg7V372
S3L640KJwahskLkB7JYvr87XwPhGdJ2hiTFuFyNomuZRlRWWQQst8+e3BD6W49+wL+lLYZXrWfp8
QE7e5E1WaswsUpqOc6bM5gYrSTJs2Dd/KFfoptz8HGX8mn0suXdDXT1knYgr8kk4xflbqD4XW0vP
ao3MCcGbvOt59G1cynj7GEtFRjQSKHzcqFAGsGshoAmTv8z8GS7DZDxIRAGDPixa3EfKirA0jrne
BC3qYJQ5WFKQMNHfcwnV7mlU0+da2V3ZZLnMMzD+kkY6ZIFHHbXthAWkj69ePtxWOzWqcVU19J0X
UdbdNv/9eh9Ol+c+lqJku9oHAbFIkgmPV2UYcycw+MwWE4Z7fMmRRaMcciRg5sotAcF3uhLnyxXi
LpAHFveLaqdO60nv7+nrvXL8iopxejVv8G9Y5cK9fUus5kwfapvKVjcXrO4IeZQtFAD/MRUYNI7h
dBJazB4NBJcTTxwqwqTAB34O2NLEmeX47inYALfhX93+KW5Qq+Qaw5kyLoCbRIq4FXdBatKldbpc
PLjUAAX9//d8rU/2aPYQ1S0Ibo/UH6KWgkthJwVl5PbaKPDM7LL0G19thAIst1qyZrJpwd0PhTRe
1cTOWV1PzQ8TAWq/FF4QatI7qi4AK+pl1HPX1mf2AOsNDaakkorcD+LXMDlgDkuYzUNkuLAdIomz
8w5ZKUULs9YaHESW19OLcp8tITtL0U0CeiuPbNBO6ZfAqDJuq/rU23Av26BNfPu+FUW2rvmxxFHb
nsQDM2JhWQ+aRL4c08yfYzl6xWARUmfTGkNsVl88/5tBHeARDhW2yduDslNjljyLdN6N43bLXdif
TGyx+WjEgHtkOhfjAFps9mYTh3YZOI9pJVsaAU3RBi14nLRbEJggF1ny97eeASP+1FVlJO9QC3HO
76Yp1KCtA7eqyer7lSyjPGYbiS9QFyGpsgWSryeWiCGaz7gkd0uVLt2sIx+MqEktSPWuwLPtsaqB
Y2PwxwS34V/RPpT/avO+8zEZR6MdSo4PLkEI3EV+4b4EhmAu4bI3p2Rlz6tDdgjEkdAcJu3vtT67
MgSo9cQcv/RA75eZGb4A5xwYoE+1pYWBrV51sYseP94FgI220jHYqead94boHejNRPEiAWtKCVXw
hvkDAElyOYsREe4NIqOtFu3jFoIvxlVjfrjW6LhyVvYtGul1DOrwomn47yKO6GrdXF+42hSU/3/u
RxhK20y4JJCuVoLE6G87tSmvnlaAJMRahEAq7RUTacBZ6/swqmOfoaKJreKLwZwyl71/UKRUzpwQ
Ey5RfGoBsLwDFaA+1zXssQrf4x/+pYY/NlT2ALFayCLw0UJQy3JfzZkBF2z15ZvFB9IRBpiXS1M4
aYBg/0CL69JeAjoBm4QluQ2bAzlgeooTmxLTKSrQr7LNs4SdjkdAA70QOHdiXGgwQ459WlYXdalD
sJLWhZO2oXcfNeg89BptBMn8IMk4Ij+YM/zMa897JP5+PR8CPraSB6QJdRRAAZugQzL0CE1rrTfH
/firPW5OoTX3+kS6h1IuSPup8NGjSp2TGco5TpY4HFaCNuHkyEXOhFPkOV9LvZkVSiMdrIAlLa8L
SdiB63b85tdGA4Ic35+izCLOc7hviu7dNUi25XSCnbw7f3YEgTPybipq8lkiBlvXihoQSwo+/tST
g6yJ4x3BR/ORzsAHZziIWRaoLWrFegVkgKsL+ijk9kduI7JdG4Rgwvk91QWNJBKETKXmzFFeQiDl
BFvcLbEL3KaEssxa+I821mfztLMQWzwbe/k8d/W9G4ixaxQPAnD8Hmm7S64LEoSIgZrrq9efryZg
7Bhklz/PxXvONO1Hsk8T81QW4plNBW4iWgoCClCiiZRzia84GgMUBxDwvgGCq8z/POW0FDRkyvgw
Ymo4JZLYNU2CKrWHTY+Xf6izaoWNgp+Tm/n7EkTgjbODis4nO4/LFdaUZV6n08ZLhRm+ObnWfJmG
o+qUhsZ6/iqXTOA1Yp/GeVc0UeMiw93g34RcDN5bmoLCDZWxlBF+t1UHdIXEl1A+r+Hc2MHRenfx
5AZoy219v+95YD7G30xlp7oAqEGIihOXPpO4B0IVJ3m4pDKrCOY15wg1/OY18sfn2NPIaf4vgSEB
VndIj9D9zwDe8Fxq/A05VuexWpjfTj56NJqpfpBzGlkYqxpMmNzDHCjgtRmrEzHZi+nNT1URJCQQ
UDk1TUWOwwlxXBzrJTqYWWWOpOFwLbi/XFC02xWUnUilXHqkaZW0CVrX0CdE7AB0gPByIHUe/2Ul
04YlBzmk5KhtZ9lGlKUotEl9G5lLnss6bSRCzT3wfpZuk5Y/UEyuU+7Ih91uc6Zlsmb/gJwun7AR
rw78m0ZpGmSMg4N8I6wwqKq88zQuuFwp37XBjj8orC93j1AAYcSwz2TuamKZeJaTQ/Gde/A02rgI
Zji1yJ+hlhpGYJiZIZYij7St4/mTYAe9RJwd/RNWc4iuw8x/UQ+RLTmorjzEN7VjkgEts/kFkyzM
GKRjtn7QsWCTJy3BgOjDzHI/lRRv1lP9NJOQxyfASwDreSGjEjlGCQQvvYyHPd8YbL0yFgpF6hUL
gpzW3qwa8+vcA/RmTmJS+BsbGnrzAiuDge/J4XMKDMESzUSfPIm4aBUv6wlr/XiwZXQQ4RtrQLsz
t9bUJl5jpLHiWPNjV7ypJMryex7RtRJDXcN15Jt6SNJ3xz4miD02XfqaT3jDKRwP5HK3/siDhfYN
5n6Df1mDzoiOQGKwRNB4P/WnPZ8o6KVustm0RsFoIjFVTJS2HKPxCHX08MRGvFMasnwKbE+/OzEj
CYgpkBMawnpGP14Hradx7z83KEWSknbiiBBqNcSIT1LCSePxxoGTODKKBr4m80oJRuxbXOJi9ozS
9jrgENu48QRNANnthSd9zbzf94IJcSVYfgcQ2OSbvqV8v9/Bp8y/ztmCu4sod4hrIDF41DIyLAE8
C8W350G2eu7KwniqW+yGRmWDHeB0Ru2HKxC4/cBMvXra1nGpiCd4Fpljf393nFQsJvszcIwEt8TC
ftQCe1GA6QXeel/J4+WhhJHDL1vkaOaY4jXTuAazOHf6fjeQvMzq5p1EQ2qx0Hpw8Q0g/r9YSsd0
aIcFVP7LXB9XrL3eNNCmnArZnR0ZHy2o0l9y2LO/9xZ2xLyCwr2VOlvBhAwg/X9pBbcfmLEv5Ik/
gTcoyvbRqSFcEASTY+L+jw8DpmjCiwgBIIkbqtRMOEHPVkJrqpqu6Dq9rCwCRVbo5OL7RohyQ1uS
pA8UsQ3UvB9Pnh+Qrpk9uxP57mjvEnmW0E0eJ3Q/Snuwfhgp6KHjcXE/sYT6hX/6ncY63hTBMuHQ
W1QwojNXKOMmFQM73Dh1zq5etEJpcnO6hWP5WR1Wqhh+fxh4ZrPo4p/tdWfk9KjpkQRgYJ7u15Ag
RrD8W5rzjK13LhCyBywGw9v2B6Rl+ww1UP2ASvRhtY7M13YouqjwZ4G68ec+OHLYir8c66p3L8aO
Dfx2J6O66jOTqg2hLgVX9phiKSgG0Vhxf5SQapg6UxkDZXn0E0gmSnBGuFBvFVxJTRS3zf31A5xt
kPdJ2N5Y52hj1MRdQAIB7VVTAtEeXPxhk5/FQpmZbfFIaBjY32lSD7h6FNKqnBxihB+DV909tirQ
kLPGKWg1NfRQzVJoamhXDWWSUNcKm//+DLGHoj9xEVvt6YTX9PawC19BdtifaH0ZvXWWRvuIWNms
IjGUnNkcqABlmF64EYDCfdxStoJWfmmacmw1KMHVFnRa6qcwNKeCseL28PcSWC3HHwNBL5cNl+N1
syWquH7SjoCjIZX+VDR8nAYNBItKzCTwQJLfLI7RidtIjgDZaGFAgyG1OAwC2JeCzAAT8wZun2pg
Asf6FvsUfD9sRqTUClvarr9x4MVes6hFVeKokfIFf//pH5u446Ojqd6D0c9VNVZ68oTIoToMrE14
0CnIJjj/Gsdnpds0c0AWrzfuADH3/rLnCqV859G9Q+FUUDAuNVJGf6FlM147uFIIG9vF6s+Tk5Qc
x0dDWrc9ytRwrW7LhwqZcNY+Cdp62c7SHbfGjW7jOcey6ewJjTLt/2MpN8kGM0uaVv1DWyoHjKZ6
K2+1PSff549SmfKDXLbKZhTA4cysPTBk2J/PDAg8D9VIjxkvXSlWuq4Fr6oVgTOQf40TXEPklyJv
UL7RYG098CsvqlN7nY9CZYwe+K4u4BhZ5riy9EAly/Ii4ZXJo5t3fdLuEC17qh52Fu0nBBfRSmr4
TwNd6Cgtt5+18blWZ3hqDQ0LAC0zCf8mzHoNPvHnWh5FN1zRNDMwrgHEWCYigSC3epHMDdex3ryG
WIz6inftDpY5bZZCLqRSpo2916MPFQtadJ6ZsaSS80YJ49uK1wUr1g5CudDYZg0ZeAs4ijqfeRRZ
elhRaCfXbll//BT4TDy9orbaiBaug96X+qKNoGUzYeEQqKDkYzfCwsyIroAjFZAAjaPSVKaVM/6m
TjcEcyUdvktvUJao7SRgQnxPLXzIze2aQhzArQMqV1vweHw0yAq2LvlVbu8+1aHYdV4RdBVvl0R0
GvXQXdl3ucrgyavN6BmBe5lv5n2SfNwhdeIkfxrAA26wxok0tHOX9SkRj2YS7Dz3DtV56uOUp7a5
gWTI8/iaOb7jMiaRjhsRodu1Nm9aUwpt/4BQad9nMJ8AB1d4j4Aj+vh3YSwDxK7fLiie1U0zfXAo
FvM9hkbSVH/Ncnw5K7qrK1/E2mxDnjYA4u4kqIuEnVX3d3xVoPjZozgE2JpQqjipWL22/UJKUn9c
vVzGtm2sp4XqXIm6o7OLSK18mRRXOGlyoP7jTtIqz+jERKkpah/dFaaPgHTcslaGMjCmUdLTm/7v
xCjAUGFGd7mbMReRiVwlAuH1IgHSiY1TKFi6hrC1ZGL6llPnwFZ+vs19xWaxjF0zFPdt+uUhyFMY
nG5PmZzwwDqdeC3deGuWAPzbwZZqyMJzZWHzRhKZIIjSDLxXwPKHxH6UTLz9tteLGK4Do8XBc+7E
FHrc51DOOFJtW90NMJkXYxaDgJ364pmsgwx3fNJwhlo7Z2C+SC2zLJUQz2Iib7OQ9+nsOGcuK1uU
ZlJAffprm9l7ERN/yZg+n+f98KH7y+ciA+tydH6DOp4U+UAfS9aDgPBirtXEJsqWuVkJo6bBNONF
6aU97dFxvzS2Zra9fmeQaNN7oejQLaLjZmfLYodBck/z+CSDYzJ64mIicdEl/NsSzs4loD+YS0A8
1/aoMvruo6JLdrzf6uQgwS7UMTeG7GYMpNlqy9f1/+I5R7NpMipxRmdjmPK9LS9NG+gJsZr/ZBZu
/46H22vjfsqQWr0Hp/DBTti3sWHaa1DC62b8vyAyiRgK8e+v4U1//AUepFL5swKBdVVx2/BOhI8K
mvo2rp5x6Tr0E9lHTXnuQ+ECQyd3qnOeYuojsVw5rBhEJG/fokJ2umgC85FMrllxklkPRZgIDBRm
74ByB5i0GJmqw1RX9B4IuO9NveOWugiJ0TmQ4ZbH5qHB4wI+7MY/7bPAiZthyj31miXQcl7PUkO3
ZS7mNDi5Cl+V9IhBxg5HKVN956UM1/t6n3VmQwneIFA7omQUblqv+7QIGzFP1PD0pQpblJCLRBXt
57U9VxPDsNNiAGOx4LWSl1VbCvmon4He5Fbbpb3TckdIPGp+3ZqArJ/t/nBCtr07iuwiHELABqVL
xr5a9iWzaDXxURAgFDMeatOpw0qsAyYBA3LFvBF9TClZ8zlMfhJvtbpfjyNxxfC9kJsmiE+/dzJ5
9laEhI63IS0FECqvHa2Dc5iFvwaU0+mRSC5JyAqMEey9D38oe59oSYxh65RFrYDoo5sLDK/u0r/y
NcoAbyIAO8itoRE7pM16IAZx5eUe11EdkSTUeYXURTck310wZKG+QnXBC/AIK2iQ0Sag2x40hB3I
+ZvJi26Rhfx/rcN92DLAVz6qFQdTH1rISXxXR6X635BqNbNGLb9f7MuTSy2bvevD1Omvl06x98Il
EzUYEOkQS3dYA7/m1kmS7gkGAo7NnPIP9OroA+eFzy8uTRQ1lXGcnxsNBd7NIfEYdBwuToAQVUVZ
9IAfjbm+A2FezWwDhaZvQMOjfo0IP3uyhEFg2hbevsZJP0FqL+HCXheUda8dKgOONsbi0Qw2dwC2
FJpM9tapdLr1Ed5Juj+8YQol/2drmiStqwlmXvlG1v/exBumgiJ7ZtBXsD2GwHkzpeA0VZpYGUMO
PxHOnxYk+3nxx5BRqQGdSjP5P22UAdhIL+VMclFzAYS1nu//BpxKT3WskV6KFabJKYUKgbIgcH4b
FxKpbbJpWXmv7TgTbMOx65X0yinfaVfBv5BXD3CKNJ29GltfC3kH7cY/GBqcYCu3X2zhVfH3zG6M
81PPt8Wi9Qy1JhyBcA97jvVkL07fQTEm3Lca/0xEnJhKI2Dacv7/3upXMUTBP4QSR1gHGkYmAY07
O9LY0r7JhfBYr+rk9NOkw0Me9bOdYD8W6OxjFAsvg9/0rNPitrf3t118zT5V7eWFxJWQxIwpI1Is
lFv5zJxkycxildmA2ogfL4ROatfPCVy3h1svnT5+qM2vKHwcmYKoxqV98PQg4osMZ+W/nxJ7B3WU
HySf9ACtuTRgCnV3FyezDG88+zbFbUm7apPY4TLu5DC8bDBHrXTl81qRYBUhHSyJjQOIk2orhSYI
tk1ZYXkdcJcJo1Jg+GxSPd4EydyeNrF52c6m7YTIy1CI8G1L67/zIGVnCl3/e2CxUTs1aGxC8Gsd
igUsAFkTWrojIoLREqIh7aK7S+FJ8bWVjXRg5/7SL1MfRHclkrSAUp1H/jvy2YsWtv8Dl4Kt6DGJ
3dITBjqCr2Epb/1NxPAK1072MP+KKZ73aj3mpEj18igpoA9PW2eQWI5eiT+FL/1FEwiVuPUv1Zc/
Nzn+PXSQ7+4PdK58qqMqNNzuidjfHKkKi5Lsx7OofwPqv7qqVGNVb8F1zQqhR9duLWNCa47j8tt/
MgTzXWR3NWS95FpsEjJo2elZXxnZExCW9QEWHCqNDBB0hWttSlBUHFm70TBZ5qnIEIot96OpKozQ
BVk8W637/0lu5cOX3sGI5AlnNRjEavgXdaeAMaW8mosAEclKsYfjc902DWggbrQs+5h+VGRXtk4M
KLRI2qTThu6spg6VWycIiTnmrxPuU5Jw2oCftWrB1WNgRfKKVOvVj/UrWsrqlcaYlpE0IDT/IIsd
tXxNTOm5b15fsrmDKL0UFu5NyYF1kRl8AgKt8sdxkyI606yiB1TItKZ191VlwDy3Yb0+QLMTaiyS
L0MiPiBanSzIN+nP8cSWSiEJPdud1qW3PqTNWlo1CDfbJpB6vEjZ3RT3ihJ3QL3pK/ADGDdDKqUn
TV42jgbLFcbrLQ/Nx/5Pw8As+V40OwiVc3rgPP8/nnsVVmm2RWvyLYO+dANduml5tckqn5H0IGu/
+Oe/batDNY7rO3ALKICe/d5BNRxhYc+THEebkN1mfYPXTup6iTzsHCzYpKz+0Gflt5P2on8I8GlB
bhUebFxAGGZ1F8TH3JYSUID/1ZDfj8Q8oR2JYQFNyKUdvWXdCZGfEBcLQsIgtz8HB/ZT5j3RT8J8
XUWd6jdrACew011m1O6P/93fRYSo7/f3hUga6CGP+0hVG0kQwd0aR9NEheJ/sEWz7E3thyRyBCQ7
xepcqaVNXGvaWgWg+OEFcitD0fNoCCXsRZ5lo6kVLIMv4jWG1YZa2SfYvHjSDA4xfSBT+ur6mHZj
A8fWSTRLv5tcL4sV7D5qK2pWm+WWyO+bQI+t/r7B1h14hBWAxtszRo+kjTzwVh/nKPz+uig5gbUu
8cyxWkA27jXplMSV1NQd08h71F0/N5VZ4cXANKlxNOKypbwxKraY0GqZFFD8pnHUqVZ+vWl2dHuI
jUIe4ZCSjjECd6veRm9m8zOEqzh/z7xliGZu6nvMH7WfNACx6uw3YOgFs+umoOhl2RtfAFBBNGjg
LVCqjvLnrdPga4lWMamx9CCLMHYifey+6P/4EXYQ9Zj21VANs3DfLddXpPlkN3Agj3dLMljLHd1C
HFBDeS8s9usFwATHYhmZYdUcTYr55H22uFLxZiMPpLS2WZzxvVFTNCWO3QE7GckzneUPrOGvZ+JN
fE+fOJUAXkQ26ciznQsYeIAju4pq+bG4ununqjnkjqd/znYn0WTD7MHzbLVImvQyPgGR+R7WIefw
ZCFR0XAB/pUXrqJHMRh49oG1iIZdgO2pquBYFueY+WxQu6tnLluZCsY6KJUkO/OrFYKsAF3q/rE4
NHGVc7PkwJ+djtwB2ik6jImeof9XRpnJ0ORnlAdDo/g8WSSvP/pCMGe7e3jkgqP/49EDjr9iMrJD
JCn3YmJs4PfKqpiIi9JyDt9I4ATT/Pe1XL/smUynxeXhs6YUUf86WFl/zniHGV7qBcgXaJZEDhRO
6+8FnawpaAUJ6beDmA5aeSJRcEY0o0UHz/L1iUiM/8i4mggfibY7NiL2aL10i7Wfpj0dnbn29hTd
JDSojldaz1gQdvSUnINfJHZ1AiKtZEVKyx0BqsDmdJ7YqHt4RWb0Rh49dUeXfJI7M2DyMcMRO0D1
ZgsHGKlDwvIg3auX3R+PnRWFpsByarAT3oY64u74htiIX88W0Awdbte4jd68WlgVav85AaNWjxDN
EzMLeDIcGGIIuDshHPSDjHdEon5RvW//f/yg/HHT1EpTH3GuxRRvrzD8slW1NYziZRRwiOm0Ogj8
oCGCPww0Hh8OhVKSmgvBsA+PSEVzbj9Z4AtruwFAx5IyLe+186vQ4703vGOgwopXhWsAAtseTYR1
EjKCLwDKu7DppJENRyQkxU0C9t4nkTOPUh5jRY4Cpi4pyj8+AK8smnzTfGBjsMHf/BRtQDFPlkMv
/aq+KxuHgCUS4pt4JRN48dSE74NSHe/Vc5iOEUVG0ZUeDy/sQDAc7yVGFEeFvBgonBsdiLAkc0Ov
wES73Z9VcUfRGL+RlsGhPhCYwxw8ziuSSQ9DFFvrvMBUbVliM86bDRzoO4WekozQTahGmuGJzsTz
hvp2r1IPR9VwhFU61Xzg51XVP/WHdyctmnCCSmEfaByaMRpPgTs5+wl6Neymp+8nzt+U9pym00Bf
y2CMX7QdhgdzyR3bZ3Adh9BjqMG68OBn6tbMHYxI0cIRA9bEN3kMy7icyGMD+wu85QiQlk1Wa8nP
8weJV+Z7v3ij3kUYN+Ft72fmL09oObXwjJaTqFFWH/oO1qLrT4zWb51TLD72pH6hgenKNGXHNfZe
uWEx3k3G20FouVQEwdESgOWWtic0YkWLhnmxHqyNi0tdOjnKJ/IgolpGV+CJeyxTggqeSPTGVyNY
KVFXwtqUaupplECtqcEEmHN0oHc4BF2i+7uGMaroolPMshEUfMR6g+Kv1bOQ6Sz9tkF/fpkqqde6
QXA90PduaROXSWl/U2AkkI801yQ1CJtFhYr70KGF3gk50f4TWxFSBgYNZVqP0wM7PjQmk1CLA0WD
Pivv9n7TPrs4+QWuAwPH3JGpomwLomvfuAhWww4Kk+DrMNY7v1/TNqWlde5oBQqZbZbdWWMaIjXe
Cz9slTN5KY/L6C26/+Eu/a8A0XSDOs1zRzWwP9xaHuUPc9nBRTEmpu2nO4Mp1vihAc0CO/LTEVJY
DewiAS5c6U8GUJwxY65Xou99wdXc0hvgOTzNGZt3mVw0y/IaR00DWiAq4JaGnsC761cE25Bp9gWD
7JqkjEUxALJmfx/ZS8AXntEmDHbnjyCbjz8bljUb7kZfvdyWISN+RoGZSwSaaFRomIL30lgft7t1
I/YM/IFGSwQWYemEwoLSLWPvoHtdcuuPo1iQbw1RpkuYEH8EunLgQtrd1HqKbr/ceeileWv4aP1F
lqMueU5Ry7htrxsBrRnc8nCK+Xkww7DyO53nGmnKn16CuXFqToQ6qoxOVL0VumI3oiypElI/U5XK
klWyY9ji07qUGQafdIIv6pHxiGqxUEOsKjq0kqXDGSYoeb2dBq3zLslNNeV526ad6olsxGv3GsHg
qcEszVww0KO1CFdisPr6XyuNSovVTwFq53Rx3Y3Nr2XkRPibNgUBn1Gh90HsSWF1V3s3MZXHwBiW
T0EuKNOwhXRxbJwVTGbZzdebpZeZWtTgiDmLkBa70aEsKPPV7KXohzlFIZzhr3YklGQ2kSycyyUt
2n4vL3OYgHN+eMPg5UEi+zWv74mXCVDKuteSmXLssyiAcOL5QW6M+3kLK2Z4Hs4R1zrZXYnRSRvj
oJaoPB04qSj0y1mtRdMEsItwtnRYBcTdkCJE4/oS87mDp7Ig0uFpcjMkUddnD5yfD1vzBrl3+DOK
r/Fe2nccDU39Sr5eV2zyB7xul04rJ6tIJf8f0tTNWXYpPzCzVH3rKj2GffTs/XWBVAw8grcbeiSE
Esi45QcIlUFyA2qoQsNlBwIckYI23d7TYcsQByMSBypLTvc/TIHKPKdMK+46lm6/atDggvasTMsb
xd2cB/uF2eMDwl3fVGWeO3+ybWbpZEYvpHZ3Po7B29vSrYXAdVWVw4lX/LZR/E9DF6WLnqKS9jZa
ZoyryDI6O76gyyLekvLFgbSqgVpwjPacd916hi/My6cSCoC/lyCOcvNEr+NYddezAqwuMdqhqroH
0zp1jKXTP64q2zHfUcDghoXJN0bZ7hzAUFqSTBqbm1ZXTJ/fIGX454KjnfzDlFLYX9IYL+BkSpro
dN5l6G7OiBk4eu5GpXDFFkGkzNMGzZoXed/Ac1Cvcy5J
`protect end_protected

