

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
E82wkdGPZb/+6GZoDi5HpckkoDtuL8TGRb/JCIEDYKunG0ehlHY7rWSAl7AxBVkDytYXn4VY0NY3
tD816aZ/Tg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aN+8nTYiRF19Ga2xgugxmmkjykOIKDSAJe8CuGlE1RsIGMA/TeZJn/LIOmkC0L4RXBBy5zkZr6mC
39gWvg+KhH324/pLiKCLqvJkIObctxdk1QghQFlwGyR5AgwumO5V8XR0wkFrGx5lcmF5I1Ic7QCL
4FCmeVtU3m0TggWFC7E=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aDXP5DZMSmAZ37R6bG0c2an3UXXBQ9f2UcCbZO9jybJiEbg3jaEsz9OP8BILMEuM2Gg6zqGospJo
IL0GjwnUkhmqiXNrUyuU2ZA9j5Qfpqi0cT39WDwUPJ8gireHKMW3Lk2XSOOhzAT2gL6kjlBz97a9
e5WZk5XJ4JpzHsyykVOoT9yBzVvTvBYrbMxRFsaT4GZ3NCp2/bL7FcAdHRGbG5cNEc+P//C3rwO8
4GNkm0wKVMVQq/2HclGOKJAykNBN7fGuG7zIF27nKqnI3IBVFzw28uEsxwVFMpLMQ1Amv9lQcw/X
S+F0+1sbjSvaH4de4WOv3cOUzYKQ/wzN6fSahQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c+SPO+b2cpVqItr9nAdAKH8LRjqZZjyv88QHjXDKD8kCd5SL0IXE6XqQ/EIjme3B6XJax0d6vBvr
92G/L1QzXOo8P82zgbpcUFM1hqtYFVROwwLTcIHV5QmMcqgWTv/CxjwYFY9l1w/ADUzzHakm7vO5
G+sQHpPE4aud4403sjY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T8GeY0or01NdwqMo6UKJMUTsmtP7APuN0oCIY7KzFu+PsK+FyNTk9rSPzJS4j6dAZuNV0qTymCiX
Xbb3asOZtqkbmx9Ts0TBudlU37PFSlhj9aboLv0+uBJsltC8lWgypATvI3dldUNiHT8HwKeBDDaM
ge1f8g9YSSRm9Jao06pgbL/b6i2WQcOEh+n+/rJDy+mhlYh4b7sJni6U+KkkIH+Nz+FTmo2KpEia
kiQmZaPY0KLlWtwgAmS9D9WXDnBy7lDRle2NygR7a23rjPwxBp5MqpWylPuquQQaCFWvB6BJrqSH
TxLzvd+PYmz3XQMRs1MJrzzaNEb2P8EXhMkKPA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12384)
`protect data_block
hENdu096VcnC3s3n7QlzYy5IZJYn0HINq41Jn0xW2faASoDFaDaYvDe3zSSr3GjJzOmQFGXCbXGF
tlwE90t8Lg5wU1FmRhwxxcMCYNhH9SJ0m5kc9gw2aut+PXfcrYE6nSp+DJb7jpBWYQJK249ReUBo
QADdRFLojwpYvFAF6jL5Qbdnmik48qfzyuwZH2Ozxs4qda70RCdOdBsNfqddFqXuiN+r4gORTJ+k
h14ZKVSfhDMaO0DNcaObfLeaX/Pg9jiSr+Oh5WEVAHstXMEVkVEAqhsbHNlmV62PY5JIsNzkbX5j
hbvuIzAIM3Uvwqzo0OZcqYpx7a4E1neB3uDbU4Rq/CVqOkmWO6d9xSus0vxI/LsE6b0zF7E4svOi
LMmZ8HR9WP1cMezBTJGUuiM2RPu+Aej/1bHNlkAvw8uMtBDAKJRJ1fjuYoF4DjIYICAZc3CCmttA
2cXWruFcnIlEIWMCvBtpng/mQK//plGMFroAnVHyVc6Ru8RngMIIlw2fUo64rStE+Vow+IGZ5bGz
SMFBCJFKpcWhyqpd+6swGG7zvSzX3Gi139CN8mJ1ei5OFqrdUUxIItYvd9etT48M8OLqMrpoFi8X
PKkpxtg3d6bKIF7XWcR2+22hpq/u4P3It7emOYPyvvr6VACmuB3I8YTc3zWZu9juw0m6oE++ksQD
UUKwzlujyRDKULJVpuW4/FWHsAMGZPT1mJQGbZPuGGT94rhSILYVYovYgAodOKZ1S41M5ckEU5DX
XNe5baGc2JorOATd4NxSG8m+FmCXSGUSqHxpiIfc7OlfdCRtBcELaaYnE520IgW3++1tVvlUZi1u
+M6oBrHd/mlTyeAkYNeGd/DZBbk61flPmlAeit02Agfxn3cuRq87rmnZOUBfkunGDySYdi+CmwdU
cVlx0iGAc0lSIA4gH9Rsbj43VyCutR+3pvGKsM8f6qcJjNi/P0EwYgtmEjrrZjC7pLgci88WpAZr
3xq6bKVi1Rab/sCIhQmbX1BrQZUZYmSYvDNkXBIl4Khql+aprDa3eH4EqEYbcc6zeD8pPCPVK8+p
qvtc1rXErFjK5qzAhiFjVdosoBMH+D+w+fI/NauzDDAI6rirPUH5dh6pse+cx6LoUsJI4BeZG6Fw
uEqoo62sovcNyhesYyPlIs73GkVRmNcbcwLDP9ALEpcAipzbjBNYP1EFxGH9HKnviQkkuJJWfi7s
LdAVryFHUghOibt6M9T11aXJN9d0kyns2rIaMCC9x2a4twFUdqmsfkNufLTUiGeQzQcFFwEyiGIR
kgZwYsRw8kTjdxDTZ6EAEQzN1TeoTTFTm2N88oZCi2VGj4kC3D+kp3946qgZUI9tmR4HjKBJ0Pu1
+xYlZLBnvesFBGSJTck5N1tgdc+Wkz9OnBptHVl+RjRjZOL6qPLp03xXa6SQpImgIdywcIZmAWMk
pQJuBuZhXhZKXOvbC6coBg3l0b1Suuvi6d9J5wc3RRC17rT9qgaT001MMTjUlbM2ZIFS1XMqd7ii
WwQbjjmDuofpS2gGkgw/UUt6Paxa1Xa+mgAqNmyL/2whbMHWnmxEHccZylgAPlIaBoQD2ZgeBA7x
EmcCSmJHqpdwzDuHuARf+m2LgTAIe2bFUv8gCJVy3Kqw/ZTh0xJE034Ee7qnZ5qplVPyPFYC/xnu
7DjX/kznVPzPff99nUHR6J+EAFx/KJ3lfBev1fwUqm4XBRAz/RzaqwX6z58iPp8qO2+3uo7Q4JFJ
R4BfbTLJWvh+NLwMiiFjxTmlDE4dEEegcpp56P20UwoS3Ut4XrKQnVqaTk5mmKPJPKJYvBcCARWn
OrXMQaySLh16UTXt0yScq3Cd5U5q2wPSvaeBgj5F01L9GI+uR1UUM0S+/Tivt3+XUK4SOjosJoCN
5XXGYLJWlNTC0rHr+QBXRRx9b+4RlWJD9BqPEUuTvo2tRRbJS6RfN8VpOK8qWn2Bmmqh7f4jI1aD
G+pKhyQU1ESbXL5g6tjq3PSqaxl4FH7szToDmOFnjeLclOoIZbTTTqJA26oSz3gB2PjIotZl9wMa
6viZcwk3eVJa3IYqc7g0uW+yNrJh96ot4BBl6dlxLsZ/r0pkupaRbV9iX6mQNBzWSxJAsffxaYjd
pR7Y/7baDOdybKWC1e6JHNtNl9YQutgbQ9cZXu2ffP6HqVLL9WWqjfDDmlq8OlE1f7xUDJidzRtn
butNHig3xSB9JTeyBAPIafXzlylXES7WrZZSA14KurrrugBU5oTR7MY4ruFtLIt3p0UpF8tsnzPy
XdWlygnIezHNEf6tkSUTw66GHct6E83QkxXrb1xrIGmEnJeTlRdUN3wb93r7bUGCXfQzSo1nJsvZ
g+CMfYjbjG3aGf72OkFUloSkzyyMM03rLrXPG5yaIsTRYwOV8AX4fPa2fqdzauWezZ0avqtkrNM/
+dCOJxLERJymWb7QSHfHJ8di28eIqiYRH8EdxY/rbpafWdoCqIuvIiefsXfqK7K37MsR2hlflUV4
/4G2/Ay5BGm2Hk/g+qKTp93hL8qdjwKVZysze7bNpTXOaL4PRMha0XheihR+zXJs/7MrLCMqBCro
qyJbD3iaWz6QCBeFnjZj9M+l0pYnqUKdTCH9renXbvL4UmL1rqG88xu3mTax1EojeCvg6nuUjhvi
hE29PxkRnXhoBrQeYKGY8UmwJG43VKPT3JaxVH9lSfFL4ftQDl4CMTdADhWEAMjVln7xLvpDHhEU
7eboAXo4IWxHHrRvMkl4fCrGNTnC4CJZaYBQWoPxIzx47pqlgYemOWXmlKR6f+oij1WPRjv2RQkX
4yMASQZ+ubOSTkAzdQK2i7LQSrPnQyJhxjiUqNLX5NbzP1Ws0Wi8MKZsczaDJC+93/VwRcjOXGBQ
MBiHYbw2fMvlUePxX7RCyU0KWhWkvi3SZ+BGulYfxcGHWx34HlJUrMkjrWGYPBxMEH/bAKOlu0QT
fMYptTOw+li96+ZAQ9IbZSVLcJtoHfEBH6A9nDaCnfvMl+W/BxCaCXavgelButA93D9rzRREH96o
8eRlWDqN4oKvMv4nMFCcz0PYNMFBehCYS93/vJvRun+wjelECJSUCAGpS4LujHJHYj9ujJlgIMx3
zhJq8UeMWSj7QP0PfjUARW4FuYdpLZje+Bd0s+oiKqSe03b2YQlMZjhBd5uqgSx8rQ5Q8eo/HEif
ZpwfKOs6kA+0UFIIF5Ovulz2SAqDFLNl7DYanwJSufMettAFDoaPDLXKe1E1e1O2GWycgL1lWm9W
aVaiwvMtQbnt4Wl0tIFw222OSpfnN55sEu+kcdbuO2LJDGQ3CCrY5qQsyvC4LwnWIxqdOZORY91o
Z6xlO1v2i7AAW/GmYnAbAalwyq4O2yiT4KvfMIZEnPV/fjJrGIVaBMPcWmGDnCP3eK/LT+8acBCa
lue6EpgLxbOvZW4vSwQ16EVja39XqleFQsIt+aQpiJ3qiWBOe4iPi+ISJoBSH/+RXV37IICIU7YT
rpsu+CTvwHu/jNINWWqS8NsfCd2hM+kbDzgvrGBKd2Xwx++MRAItu2mqHdWeaZ/ZSrgZqAa+zdv4
5z3ztLJxSzB8nKMECkT+uifHhhdxUco/QZGgzxuXSq/rNPpIxUzMsVNJKt1EosFePxrQFywVLRvU
LGKFO+nm+3oJa2+WzkiCCSpFDyWpkWdkS7AIy2difYit5JDV2zBiDT+2Puo47lfo0CL8sxEF9RYd
efJfoDGldw0ctBAnK8qWD+WKKWDSRnTlnxOfL1EDDxiengeNaW1Ky9/NBIUnVugHprLoRw9ZOOl7
Bt67ckSpM6WNhqKdvPh4jFfZ/kkwcGESx3GaMBERKn5ZZg8olsyySh1bI9wNVF+H/PBsINi3kZrJ
+gTfn/UGuj9X2NwqmVqKGzA5aaLbkjR718mSsxRQRxdtwTAVUEBJICwDLXafYabn2/S+0H4mFniw
TdLxcvMo3G5WU7oZEjCiOvxKslGdH1925Gx/dDQevGf7xOuzA5cbuSstCj+vqaTJu/QGtqMhhMsm
WCKCOe0VoMCPm9VtFI5ESCXQALIHbsB0cxg4gqQujScNMzBJZHg6IynkLegd9m7Tlf4nAQ0ZfdS/
/aQilxSe9+TlzsIxWRI3sbAXAmiQfVZfFqM1LplY20XaGeaPHl4UFIMiChXsqu5E55+MbR6E3gj8
ZVgy40+VrWI1zjQVSpz+vplEymv6hp5kAIRhCmUIY0yK60YRqmISfnzWApaYyO1ZMTdAyz8HFJoI
UjP+eUrimkVqcCEd6YHLWCwunwREW5tf8u2eHs9UtAowEol49+F0n29o7oll/pg3ctyBZayb9Okk
Wyw1wGyWbURHLMed5wT+QghcUULOaIfR3YPO3h2mJG6abW+Zx1EHl/V414v0Axrg8bXggNe1B0QI
iksN/AoZ4J97g8jrxA7z+WLIiU0yw/rmFaZGrZqeVeNWxz6hc6HRkcWgk3zSy7nutenfQfZsvQOL
vscLsmJqE+v/E+zmUUzouMNXHJ7Z3e1C3IZzdT3140h2KcaIDDxRBTZe4p5oCs8LkEv55+/PvQy8
K+dfnzyR7l9U6f1DJueraZPrYMhjEgCN+EaJbL/yZAAUhPukqYa7ZBhkmJD6KbJp9DRx8+JSE39F
NGl7NxBF6IBDb0sQJJFXUQVbYOFoAGJdGybwfX5EIljDYaDTX4Ytjle0gyCms1XcEcooM200eekV
6X03OYJyd0uTJdoaPIeBx2oqDFOnqfmT7qQuRnBjWWFU0gi8faPdRAfDvHs5TRFIR7D5oVTUM1xw
RfkMKuJOumu6uPdzCJjsX9jZxhB1EHi11TOQsolsywBCkKmUOaGICchiDi2JY8fTKkLLAQskHS/5
2rSR1xHz7DIvCUkr2XIqzFHeRfJ8Lhsh1AMQI18fnO0SWQgIgMyXe5ASDcmyWGCmnp8AcdlRslGq
gQwjIjC6NkKft0Mnh217qHHCRoQ8jmzT9/oh0wq8JsIJXBuyUTNOZAzZKDs3jPXglmMeUXc+ctP/
YLdCOtdAwv6D9583bgM+d7jwwFYiGWby/76SqUbjPQF14Sa9gAOtKgIo8B5D2/ALvAV/BjpErtKG
blSRV4M9ioip3glmQYcqbF6ErIuWJqtf+BulgFNMQ+tFlzrvX/7WrG6w6hv0t+eiwgThBTGEBfTj
gD8s9MlWOcLsLP37IWJr7uv8HG79ZenrUMj5HaGRDbhWlpI5/pqn16LNpoUqgZnjrCwKvp0/FEjT
ioyLbLhfzHA2n7tKe25xATxfAo72Aw7EjwVMtsfe7GSJH+hpYKB7rDj0Kn4iCuoMXPqE/rPor6Jh
saRwvWK6rrO/CBZd2M4G/HUOMMvUJdJN3oSOS266RoJHH0sI+DbHXkPDDvQpXErDuVnne/yTb/au
shYWcKXpQ3cOIt3RN8/VySjRz0Phsz1GWhA0Kz3G3AKaJfxWbSs/WJ20EBNJnaOQFz/qRfB16ioq
4vf75jtmzcMEjfUIMcvmSnqbRv9TYkPgB+afs1IDud066pBhwfwBAb1zZW75C3oavdTVQtaOA8Mk
ttW5ToyIi6Kak3jL+CbmmxuO4mE89V5B9svXn5qaIwUdYU+F2B9m8bWlJbCJdI/fcikjjvPApdMF
7SJiew+7Fslpqx9PXX+VVPiBQ6RbNpwGQtK3tnmyBGabutv1Vb+xOYUReafVZ3pE5i0xPMOGQApn
N6CqRCdgS3Ugm6eo6UzcEmrNV667obZsPt6/u3EKV3yyzzXyge+TEr7XOjQLOGzyDzFX0f0o8hs0
wAcZtvdBwfdJ3sCcQBBdL1/eA7jSSu4DPRirQdjS5CwUMlfh30d3VQBcvnY7S22tehQrgilvjC6T
Z1KCajYmP5hmgmeHVzAeQ0GDRxWVCnh65W5eY+A4IsKSalNhXvSXCi9o1PEPxnuKakcY48TXzwAM
1bcnnXE+8OyWw2X3ZKYeV0Fn1KGsq0kYRYpV3SVJjf7/i5VPBMDAVw95j9AArMg0wHm83/nbtC2W
5NaLmApvbp6YgPRqvWFVLkwatb9CuaUNSq3DM+mPepFHoy/MQ4IdSiW/Ud/x3/XLrfmUSD361K+j
Cy0WfgEbABA6Ksb9bRB1G2mh3MiMBcRuYPdQqRrVr/qZA379GOERkrZ66cnC782QGCq2nmSKxyKE
yP1SNCvwyv0PAi65jDCYWi7YsHVLL4RWYDJRg90ejLauEdlT5Lz/9M04szWNKnq6LUvL7+n6URZc
G3txRAn2mgMyaHMMnEOy570peFI3D0AOoeJvjZ6yPYNtu8bkMZftpjZwIvBkatSkriiwSgRPVBlH
PkQ+Mb0eRuUSNaHDTb9OQPeBXxAn4y2mmXI2TBsGttWY3fHvlg3pnyuCaUmhzQTRcIRUje7FyQym
eNEquGNl5V5taHoauVntWYmm8K8ROEDXbpdPNBFHYGmWXVlkW3cH/ah/KYnnx/r2HKT1nsrrygAr
yb2u7ao0oEQnjVFN0U52K9WVirru1zuawaAplQnJjptKRU4EA9A5m7dvtuwoTQO9HT9wXpuixgeE
FTSJFaQGZm4Rcl7fcPKJxm51Ba3GG+FtdYLtuWHiCw0uvkAgGptCVEnfzZm7GaC7NlqGXwggaupr
rJAHaGRu3WWSugNivgP2MR0CQ6tMOUD0+dmrFdZEzL0HM511/sqmFnmobUcpFnSiECB2+E5sk5po
3xTYlDrhAXFQJRJm6oYToCaq3wjyd8JH9KZ/sl75JkNMT9Q6xRCoNNJIL6KX8o2FC3KG9HA11N1O
QCoemkVXaIHAB0VLzFgdVpbvgF4x3kvVbdZF/lybCInhBQKOOiQKV6l6tnLycd9HYAAxZVvmdrVR
qjvdRHNu5f2bYUDsTlEvVKYmHtJ1GDEnIlOsaQ+88ekzd9O8ixWv5t+K0uoZivFc+t1eCa25J/le
Jhu4Otz7YpxTjxSX0umgSvrsRF9WYxzwZv6PmvOG5q0c6daxS8WZ+uSJ9FGgBpuOr2tAxKOv2DpT
uddWQBShLO1mly2XpsmVrg0Hld9giI65yLSf0Lfx0x4FschUCvqRMolnj0b0M0wFZ0ICv3IplvTo
nUAZ3HcP/O7VIUdICcNjCkJsC6UwjC5WtWaDr+4FEpdd+3q9exmgHKDq/swvNa9nweqahuFTOwfF
13Rlw2ybzOEvOXbAF8v7qk94W/KIV5RtAscXPDdlK41qeAb69ihkmytdSQrJB4QLO/HjREVokyEX
wKtHl/wajr2LAQEr8tHCpGOlCTRxoDxSBdXI67FenlftScxgiuUF3XFcsSGD/AvKOjoGzYHxBfU6
DKGywGILwTwRNFWO7JfPPpCXyxtqd1r851ffQJdy45ta8n3Ofi9INpQgn6PGpOd4gTkfn2jPwYLi
/MZtBk9goDq7rDCJ7jFux/cgRdrxUUvQqFeYNvFzFWw8Q2CEHpK2VBKTi5jf6ZjEYe1tYW/XjxoC
BeRYOuBOROoFYU0o8lNtt1rja1FPjroWr8JYwZif4GTERtIVofHT41BqAfdcx5LnZzzw8XVGJbAv
qDLxvfmoygFxxfjvrf+XObEXarTO72gyJ/NORqyOnaBbyGpnrtke7Ay7Up2bpTB1x2j4mHstGemI
+QMC+1qryX1xHvkJlm0JRaCBJE2eHG8pNI8wI6lGoBg+ldj++2rbbLRCxAYdK4BcOCdVOZowUmG1
djPVCj3hsoFCvD8N/I51ELh0XFNz5dSCpIkRGXDSB+AMLEBxJa+KaQ1jZIYExcdGgZepOYhNIHO1
5HtnFYvN0+03JjiSf8oK75TPRaV5uGI4/DDhmlB2yNJPzKw+m56wcaISYQ1+JVXwkslVRAdRYvWQ
agVZyCw3k2ypDAUedGWsP1tTGfeaB3sWZDxvBg5VYspcWc/W/BaKwFInjzkDFYeUhQoxltmgUn2h
ponKnu2SIi3isXXrz0qzfnce3q2UJGPRSYm+LYqkaqgo8GKSoZYaBeA7uefn+wKYn4DFzY5Q5rJ3
6lk5z+g7PMfNP3J6YSkb8T4jE9244wcgEDg/tsqIvpcBkgvzZg6tGtRl71w2t6XQxcC0nTvyayJA
4W53YbLl7zsO3sd/ov7kUx8Kph1S2feOXOw/P2hH7F/6SlPFj3tqVKY2aq8cT5XqWpxeh9jcQzLH
AB2rjlrXKxbwjqzCuw3j+89cAzUpWIQPAalE2OSPZ1k/oclinfQhaHqsYD5U0CoDxah1jCd4+sok
/eBO0GHqNTOrPPop+cuxYP7TrHta2oudnpK9ijRigd2Yoebqcww+72BQiOP/m3ms6Ywej1WpHhoA
X2fmCgAAuMl+pAGNbU9hJsumuWg1vnzd05/y4VsFwQ2dnVCNOSSuXlaUQYV6i7RQJuePi1NmvoJ5
7khl2nr37jeSPukksu+xaQuDewBS0X+16RKMnsI5W0dhjsYZ325LqIgpgnU6WiiaCKVoZZIU9ISw
CSLSzILWXh9EQWddQ80gCy7RNAbSy0VGHR0/fZwT9hn0h0omMN/G2gshidwpMpXelEDAzxpyZEP5
Rh/tB0EboiCnQ+2ZczeLMVUBR8RjzJmb9ftyZB0+T8TKDujpBxzrvYCwU8UFFqfVPAsmkvtSF9KG
oU3FNCKwxTF28ygCLuTN4Nij4HoDjTtlovTMLyD350ann7VC6484YEV4vve4BOZFfAEEmJrwgZeF
37bv+/pucIv9xLmT0fEPqeTbTYPrqFWAKmbyHZrbzBDr0kvwmuMhxRvsOzC7mG8SHRNYKlJmq3N4
uTpZA/eczdXfmNKA6K1vnkjqrtakPMFNVJnsAYTirkpz3InU2GrG9IdiCDoDnMVzVSFBiopZmmkI
YeCVzpRfyx0ga3vfdAezyLf48EZ44BZd0QoZtHT+wCmd3rZw5Ya4hOMHgrePZbdUfqAd1BajX4dN
SYtWHAQEFF+4CbZ22ev96/AJNHUi6RB7h/4Jk97l2lk45nHyirog7l//eE9kfpMUfKPm3bKGU6T7
8dBYuVOP0kJq177OgbAbzpjwO+3tn5cDrtS/IbDXj2kQaO4AlzqlF89W2Vn/lDKt5zCltMiKpqLu
JGwZo3cEEivSXho+tUTDugr9LM+KaZBG6l+G/2E4/qAsau3XfEX2+IAJf/rkNL4xFfeGXVkGASoo
Ub5Z4FyWFFsLCyAErbFyNINpOphOO0gbk5HsgNwP96zvQiNqGcOJupWagPyEzOA0gLn5SbpvXMXb
ifNYPuczXJyNmxvWZI21R59jAYvofVXbA3MTJoXy67pzN19scgK6NKVhKjsiNKPaXGR10l3VfpJa
C75/H9SFmDu6cx/QBRioidU4hzyV7siV9pFIl4T3p2Tt2Lvc8/42clnPFDAlYpueu0lUWzPPqqLq
zERriYl4IImaoe6ITWJWR3JuKDfP9We97SqFipkqMnApbDRK5kJFg5wEo+NbR/cMzdrp/GKUReT4
DqdIL9SGdkTQy+NNtq41mEYeGWqkcvGWSlmID5Yf4XXootUIzOAvAabLcdTNJJzpxDJxTNJrh5W0
E+mBZS2fwDLfkyDEZUneOlTc3KqpDNH4o24++s+cDeZwST3cZD9e8epKWVAOohZnqrTZ+5obijLT
RfLw90hOLP8SayM6RzFvkFcOo5GjO542tAhLL/uyp+r1E46RN10jbe2tI9pL+EgKubeP4m1anuEL
ZEO41wzY3J3AMsfFbhNS7E/U+SXcagSKQgSltqVFm+aDyDiegaiqJoPpSoS+sJfQBcrtlEW6r8cH
QE1ulkRwVLOut19gzUq8APyS6NPGq8q495OYjT45dczsien/3q8ZilvDwwrsSMzqIg3zXrAoQKqT
aoio4Txk4wcZ1RAFV3YQTDxVM1kt7vVO6NAqlXNHqEJ7TCNC1DOVmvaiGOpvAKUTfNEJxMJ6lxTF
KpaDrf1G3Hw7Fk0UastKIVSUWJwMARqYobCrWFu7UlcA9d7SUnghBiAsbtu+KiMJIXe3Xn0GEn5f
MV5T9zzDRXO2F/OGkBJeaekKz343YXzCsr5UnJkMz903QTAfSlJciU+paqAcylIinhmRHK+7T/qI
V8+Ni9XEMb8sNlDFUcMMXinww2KcfvKxgbWoflkmzqHcvuZZr4nye43vzNuiX9rq0A/o/SjwnOUN
u0XBjfmhyyV7RSDKizXLRMeP5au7O7aolhi7Nso6eIr7/QV2mumd7//VTYuMPN5YzC+vx880oppq
kRZcwGmD+xl+AgnapUuFNbPmm2wo++y+Cz53WwpLVr+R9k7xjA7kNjL7z/4ktKbKzr66qEzHS0/r
QNxWzSg/T/ht0/ypi68dIZWnd3f6fzlh5YYo6qL68ohSgU2awraVJfz1n8PP22ALFKiCn4Kmk6ie
n3cGRuMwiMmMJyPzJ7yNfNVG4x4RGQ7/GXE24XGCj9cuE7w1s4FUOE+Vd3WGWT8ORrLup2i1Dp/G
QF2Kry12/+lEHMF3dRE25eHNMWh1cNrVK0YxjAgmdPZbx6nq1jNKYTABqDM/RddXamN6HRvAIhmy
PZjCWG+mvFV0a5JF6jr7s3rpQR2wutU5vNb6mkoTL/ipI6ep1SNdlhTST3HYFYR8nspFgvR0xeKW
tA8chIx8ZY0CUqlDB1mzhqmBM8aCZ0A0sDVLfX75Lc0Sqs9/LceadX18oTLPbaA+F8jwqxNdSb8v
cq56w2hBgJ5J7AK8kO50OMao5mF+eI1BsrAzrU5dKQZGJLIcsJ/DBrTjT/s7MRJRnVp1ql+AjGsY
3NCsc/fPUARnPDIu0SNa2a5o1HJznQBVdkYJBFZg3FC7WRpbXTqlu8SfpwTNxNlFZRIGQmpDaO/A
6FT1EoZ4h2BO4WVvJofGtDUpPGuo/D/H0gAeCpUEW/rs7f/OkWf0qQlNU5jAkmTOuC34u6wKEDl4
POpFfsWN/QVMM4YL6ygF9kM6uV6c+NKkDaoW8dJY9uvxq37tQn9VeDGuV1x0epjy0xqa4shi4KWY
4mBEHyTNIgp9AG/doFJsTS+JuiyOeXnpxCB8tsUy6Xpqjnd8p4HzF6a0h4Jel9gFpGnFtOwIbiAg
4bWbVY3s0aKtyx1k0ePbYXv4mJKostCjh5Hhc8aRt28UpuMwdS93xvtsgq18NTQgi/G1Ub43jEjX
vQtM5/ZkJfeEzpTMgolalE14xJsq3nMlReymuQcabtVA7S+orZ4AMU2Dn4RIrTr+t2F7J/zxPVEu
30CupxTQfVW6zCoESp08StWKZ2VwxqH2zWj6YXj+R8k33LSQo1CkjZHgrPSy+vF7jE6Coxvmx1SR
IeVDy0Zu8fJ917EbKxpGWEUaOocioGkRdf0k8p59du49FJODJvZE/XEaO/+n4im6lO8tyBlvnOWi
9btATIjzHXEyAvbZbDjeH1nrFmylhaEh2vLNpSbaQsERgLpmQY8Og1gJsDB8SQhSMbRPNMeGJKoC
kA2K9Pf+XG85RxacV6LE2wWQj34R6yuxs5l4q2uwdNe9qm+EMtRWaR6wQXPGTKSVaYfuMiWJp2Gi
hXFHQmnOiQ5nRgYEBrJ2zRmvcHvcb7vUnd8ZKkNdCBrtMCPFo7B0YqN8algVxFeaIfpyqDDiYVSv
Bb8SUZuaNRYO/SxS3jMxcZ7uCwunXGevhpG8kYss/9zS2q+tWHfyvmRC47rN0JuUlT/rNY9qS9FV
JwwaRSCP0AATXvfU4wyaHBzERGZNwk17aPbi3ADlNtD82Ezm/8HNiyOXdJVt30d959Zx7/mvG6Xu
WrlqvlswKEFRAHAsDKvupWD8Aqtf/11+3jdtJMwgTwI32uEK9b3HJxv7C2mgmhHCVl+08al/QQKy
metPBSmQwMu+YK/62maiIOhA7LaoUp/0hugP7K9UgwMUgqG9E3e2xcecBmhFlvsXEOU+BLwT4keU
buV/JsOTG4XW8e16GWjhf9dEx+XgnMIHsD/omCFyHUXRZCGLQ6WMdCW0hfud8Y3xxm6MDrFDTULF
VkK34k1r6DAvQmBrDT7kQ0jb8UM1H8n+7AsvzkeDSQT4ZWvLmcurXP3V7tthY6UyAM6X4sEJdrRq
cHo/0wD91NxxW4keZRxGah1WE9XMGT+BczjrjLlRe3ChWANU7455KEavlWOEuSA4qdHAP7x4i39c
XZb/6kfEQiWKhpi+oqLNBuhIwcClDDzwbdZJ0q9nxQKWOrBN6Ld+e7XuPJtWFklP1FQrgpLj6Hgj
Ax9dUoPleBBcNZqkOGU+u6dY9i9M1V5kX3ksJIKr/ml4+tCNg3QNGuIgJvwQVgDR3w7br7VPxs1Q
+MVGblyh+FU3Fn2Eq4oY5f5FYf8QhbLJ4Kei4rThtshZUDZ+TC2Dg+0yBHGkU/wVs7s3whuG3Sdf
Y3hNAo7sCbIqUienWrl2HuunOFcnCfwFKzExb4sEOe6TMBpIi99Zc28i+dZ7OBTNVLtdxvreSDEU
X2Xru7qBvbCoqKv4ICJe3wpBurC6vAEXV+ZtIoOW/sFyMeD8c3am0oAd4ub40OsLD+2rCVQkH4vs
fb8FdXgBGF/m4cu7975RwHa0GJLI5yuWQXxalSQvACa/+h4JWnEYxP7kTyebuISM7O6OfjUvc09l
WltODER3zJ+TGf3iJ9wdS0GdnFhCheqxj+CrsdiCJ2d+3sWgYZFcpaQV0whAtkMCdNby68ahAGcg
ENqngMrqZP46kTn8Mf3iZSKPeH4x2SCzUgTge/d0vZR8kkP6c+1GYjZgBMyaZRJooC1fOqR1G6Lj
vGqa4p1Gn8fKEb1C96FWoP6/AFdWanY2EyrLte+uKc6KuqhB/bRROj0hTI8gwu9P9mH3rOHP+aK4
ugGBPNqlkcs3A6fFbfANYU+sRhcvcgBEEzy/8f5qigMMgB/gMO1qG6C/2+LP/UE9NtjrPgvex6A5
7s/E84SuWL//6y5GW1DKTF3NHI00TcDIfMj92RB5tgUfUz4/ybaSZnZ4Dy465yPR9INRZWoK2/qb
vdBOcD9jgsM1xSve3/JvY8pZw/6a5BZGcAxH08kVwTmoWguIj2JW8g8GyU88IJvC24KFzhv1+yGT
/xyLHyZC+syPmuny3mbnV5ngwvDrA6RKxmXG6G7y6L4m9V7xhQH65EC5hpPtWjfgAGh0gnZSMG1W
dU5VM4ukxxDhpRsF74YtacGBVy7qBE1EC5R0QrSrCqqB8rLUg4+ggu0re8aDP+V+CQMw9aEJGAlW
DXP4NYI0SCNDYayh+IeZO5/d2RC4WtPJlQHWUjGUcZQ7Dlhj8QPMYD3UnzZem24UmKqbwPYXjo7M
ruyKfgojTM63sfHxYGw5mhFaQ+hu2a74B9tpEXot801EOFKW0rmfcpZcXB+1QtjLoO0YFToRst4W
mMMr/SIDzAfoL9UNaLRwpFuI9jm+NYv/SH0nY0fAUKJsbDVf64h5Hr1C8lGeX5cpl8VgbxWHxqY3
DTnhj44anMzu8DZQmS0iE/+y9im2vjlQdMvSCbDON+sraf6PVDGjRovTx96BBs7P9o5fzB/L1Hfn
0adjNiy0k1mRe1rlEJ5noVDp0f86T9KpI5lPoaI+EXo4xz3NHPTw1fL0VavE3Zeb5lDpYY+s5Or7
vZX4gH2DzP5NafR7qs+UPJeWn30Xwf8xdwRW7N/0zYTsMbJxTg+Ko74xsAmJL2u/taRi0zbsdRTG
tIRuTCywLbYS8xP2oRozA8FTKoUg4MqEONW7tImBNTD3N3rGXZFsx3OcJIDy/YWDPUHHyNVqJWQO
YXgVoH/uvgZ1AxKQD0zLlPFCN/nVAgwV/XsSrGEs37v3q4Y4iQ6W3HaVjEVz7Yvf0UfT5ruQ9MUs
yHzgReh04DewJ7hwexQETvpavNNbhiJ9D19i4kQLz2S/yP6KB4FZtQOFi9wldfD3Svvu8PJg+RQw
AOxxFpeVbc7l19bC7Tji3jJ9Q5ZFnrQKUcDzpEj64vP0By2Hd8BEzcSC6NzCMB5HZ2kDoZMPWWtq
hGs965rv1+mJBRr1w6gEAR5rhQ7MOYwwTnpvEg9Ow5hTgZkv9NK5h3Vgm3nYws5+kzenhseuPXL2
8Z0ANYzBgsyeQ4cEH/lrnIzlPQiKbtgVD+stPernOq5t4LHlgjCIgiznYwrtS3eO+Js+KvLhNaWh
myXYGzvRxbwhyqb3hFw4DjliaIGmzfEh967K1bGq42btdgBorxcaO8nzFCshQeiIUjHtw39imA7v
PxiRJDCMwJnqDZRAxyCrnGcLT0/A6+CmzaLG3SD+OPuK+KMrKzpleGF1gCZo6ZIp0ROPrKCSHp3T
VbPHg4oBYDp/MHdrZyB89o8UCRmBfqCtYPnrkM7k1TXj3TE/6OFmEEUdTsR6CQltZPnKAjuN/ggn
GIWUVj+jzV5qIWydMaR7pPmr2bSnf3i2QVg7YuP911ZA4rvRJO2Xh44Vh51g/uCzg6PZ3+Js757v
h0qvbJVfQz4T2RVXPWenOlyZyz7JTQRHBdtdhzGccrszWNBfcGqcz/THBgDagIhD8R6YZmvdzE6m
/0aH2LfJouh0LTDytbKLjob4gmrolvBjb65UQTkB4DzSEN54uWWSUcW3D1RNIS0/mEU1PVzOsieS
tYQmiS/I3hDn93RAzd/P0FrsGImDHlWsmmsAntnSCU2J9L6KEWOgLmctFkvedyq/UfW+aOVZaxFP
X8n1O+Zf0M81inRBebEpe1uu1/P/okQaCxaKJSHA6UOOyxu2uhAkZfVuiSL9ISba4SJuOLkssV6t
FoX4k3WGtq9X4yYTOU5s8LBv+eSk0nlV5aQkUO5zDR9qYRAmx3FqHdbrXH+COWV0VQL9f5JFjRmt
PGq4TioID7j5ghXljN8QW4IheuHiPcJdypAJRwRpbRLdyHht7Woie8o7RjDxk4GNLFd7wateMSPe
Y/JH+M8PL0xiYlrMUOrtLc5hsGcMhR19u3dVOcD6XJ+MF1AAYlu6xuOJ/CRGiZLrQK2agdkxIJtz
qX85cIK07uBZuscN2tIZXRQBiqGO+a+fFTLJ7YgUshkoUb/Wy54sm1P4NigHh9cOB4UtL/DCZPC8
8bXx0m3KAr1NEC0OIUFFd4gioRtIBbl5GZCRYpokDNzyge4HphkMTxCxvPx2Gid8exY3eR35V4Uf
AjZ4wym0OFYZ72V1YOVXXICP9l4t8JXF/vIo4CG5uMtJEZfHNX3KkxlQIkeLZAL9rVHDXbWWYkkR
v9V0BY0a6HJTMV1zN1FaJJZInwTCVMUeieKFBp6A9u2gR1mi4caTVkO58V/6xUQeZqhH5zEaO6L0
kZKIjehF8s4FRIWrwleHhsjNoqW8m5K8HgyiajNnZ71bDtfbU7qq8W/1ujt5ZF8XQf00mOoPfonq
oVSOuw3SDFcvjzNTteEnxPlKJGvJfGOITgo+U6w+SENPK8RueYW9d8JrlOoVNKtErjswGkM8O4Rv
b41r6Yj7GWelKrO0cZdnbc3JQZfdCRFKze12WGHiFcvJmOtJe0rBcddL/m1JMoD60/RJSAEuZXB2
1uCFhHoRmy8KY0R5syxZiy9TJEMf7r6frCl4zFklO3vZC2B7r2XSPhyrRGgpGhPQJJX1d65CT+d9
Kwpd6BH2QpVe+j0etZjfw68ZKhQ0d6D23+3BN9o12w7hyIcZdG+c89v0OFMHxTWtGsBL18vXDR7M
4iyeKKAhWWheglwQRLkqbFxQE6u09dtTXNVpEq1+eRUziGPXBDUKMNku+gPuaA998CL+8nxl8eAj
Ei5iwPHvNWPW6JH/mGwt9Kzqn7CvOlGZBktf64leemDs4hhCJa2RJuY9OrYtPJSboUjuE/KaT2q2
QL6pg50CZStGMrpx2gQDhKwOudeOq0k8QOW8EvewI27NfmazXpil8NKYKFNQ5ak9FnazY9GsXUsv
chuy4VXnU/kFntJrKt5Pr05WLgoCnI2XbZsyCufzQqmHpxk6tETrLQ42HF78Edto/luMD1BnoXbg
wkRb3hsImWOWvoTCsugWpAPX0KxwY4mhLTCZ5xUrEsbN5Ym5rESK+DYeeBWHrLYs14bocDwJ4vCp
RZXgiUX04Y2UOtJs2JdL5lcPRwLlE4hVmvkqTGLqHcGd1Zh273QLnuwJ95/jWxPreSbAqTTVyI8C
D3UE2kl7GRC3nEBwJ8BJX4nVe61MxDN/pcLcCDmcBCP7mHTR+gxkBnuu0sqht7AUk8Ejw9vq9qZw
QAZB1DIEHs34y3lNqQXLCtrIAdcVpD3+esAN3G6zMIpK1dYVfOP6AsiEF/x0/3yM5/aGtppAwMNl
bZV7hsiDNNFdqMGNiKZ57gu4Moc/UOuzAkNBOLgnGc7H+y3UEhf45GMXBxjNmw7StsAcCs0H3sNF
rRQNEGhPdDBqvugpSHBSitEjgK7S//U1gQIAw8YQjBh6b7qpt0rldEtDJz3jXfKFnpRTsG44lVqH
Eru7ha0BrHHi+seRl28XUY2PjVFRQuGY8usrcbsu5kQ0BWTIfh3CaNNO0nh7l4KB9fm4aZAgbiIR
Jw6wafZyB/bGTfyHFUUK1686Q6HECKKxLN409c9iSL5hG2ScYLQXixlO8VNwGjgVBfQn/FX3TlbR
zQ24iSGlcmbif1R3PRwi
`protect end_protected

