

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qm+ahCoXbtCT96FlU7osNjp8Kf3rDAFQ8vMBTpaKgTo3EvHN1CM/XiHNcIsmMQ17hbL+pWxo5SQe
TeNJ1GZN0w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KB+ek3mkpx3N+ihSLNljgKYzWfCbUQKXGho6dSjrHEWrzL9W93J5UQjcPdLkP/4r8XQ5AjiJVm8G
O0+WgdiO6dbDdWggVe0UZIQ5qp9jotaT15XQQVVkD2rcK5wquost1xsRm7MTsEsCbzkhqKPM6ASZ
mpW7GzuYQ2vDPmY/r9U=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5IFnCgXf/KjXBNbWCJPfF+u/Xe3PWCvLt3/lqQEWvv6nS2jJ8qz3O+bSiUUxyt/rlAZZm5DvQ41j
Vn2wE7il4mdux1L3DFueP8Ob6UEbh6yobetr8hrEOpbRcnmnH7rXtvR+yuK3psDEpqbW7d8GyDcy
T6jGK5xIsUceYrUwudt7lxYx4bLnzP6q2c6uLhkxaoLJTWJGh28se0dzlAMX/BnMMfjK0HDKD6kp
1VwH2Gj4iT7DvyBkDmISaH7LPSlLhe+ZmQMkilflhi03bS9w9ABaqs6v4fufe3/pEUeBrvl3gRH/
oCU4QtUwSf8qfFsWdX+C6Nn7mzOb0WSGIH22+A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BAf2bWZTeSaPIqnT3j5aNO9C6t5/rcfC+/QtvmxOirWtcQ57aHowXlt817D+9PTxe4qEx5CjzmUg
9oMYSESB8IK4XXnHzrwWEKN1a7YOhI72J3KxmNssnP6jdEMx0znih/oPMXJaAdPPRUXzSczvXVqf
S7AhrmorMi/7B7tc1xI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dVk9aS2pcwcb0BrWR4Sm4FSW8QQWqHH7xHbqUaQTDLyPydXvHmrmxiDqUJWu8AAmbDSnHtBnMo/b
vhz6TIedlqcgp9o49Jh0CEli94frA6kGx65vbdl7q0c/R9+UB+XDf9B8tq4xwdSd4Twx0zVa9WGD
lmNliqJyvFk+OMbS2OJJyBNqK6eZPVzKMFkUG0UJu6TERfYV2nuxVMsugR94X7JoKx+W2jEprOdB
UQVXsqhudTLpaKEQiNqzDCaBK0P3FekkJJMtZNaV6veO7wX6Us6tTDs6pxGysSo4e6tLocXysaO7
1blW1S7foypb+e5LTkDXsQjIPmjtBTMz3Y2yyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47328)
`protect data_block
mjRVcCDFkwANXA6ooRX0mc1EpoF5eU5S+seuNHQNFRwXLnf9UA0Jwb7C4ny4zZ79KIysixX3HMuw
cys95ZfaSnPfd19eP8rfX2npu0SxcXgq05y/fGKxf0fQU/vX1FW4OiaaR55bUqbhL2qyN2K7y02Z
tiCM4WjUWx1DbluE9uvFY99I41RyfJmaayOh6SrWTOljgSLojM0ix7QMgXi3b3xUeic/WXZgp3+t
ew6xsIO0d6TTZ1QQMVTCsvUMQOjL7n1jv5PqA62pGu3YZcHN4d297KGVWOomwnwojPMbs7uPZZBT
5oiCLyeHdZd+zmQs9MQdqnWOkegLQj8g2mPSJ9rGZF7ejynX3KS7qmdMSem5Ob2UW2l1+zseeooU
W5jK0OJ7QHjOEG1ZI7Xt9oNm1mZkG0OFXJlWiZDazR87mC++lwq5oNsGOk+f+NzHYHJvN0gx2YCP
8Gqpg+Z4q+VwKb/6DGaQD3JCVUGkeZB9anEORVe0Go7vYCEoNXW+mvDBbjtwn6QC7853kFeZj/8C
0e6qMWJbwpkhrXFPte57bmTPeSpwrMppgBzIEghO7x0taU7rv1lfXdlEyP5Bu3rvNCJVYYelgh9p
5BpmMzM/dz8/dM61wNmXsZ6DoEpHJRoJYZqPqHvGIQe9Nm9SQ/+LVxUz3drDWKWXYpo1994zr6ro
Dlv42cgCUTwXq9tSM7KrD6QkHJhLjvXG3w6DI62Mtvy0/0oh4c7my43b7Oc6sSuy6QY/+rAgM8/w
5eZILW0AzUrbt14SzaHiuaQ2Q7t69uy0jn2JLYCg5WdTQbCbd0uZq0fIYhPZ63ygazfW9kBvTMf8
nihOZan6nZ7JMBLmrG8vMN4yJpbnpYDNG5AwMAIdcilaDwaF9SKgS38d71vDR9bVeSo5AXgl/Wo4
GK4Txrb3wSKZYuGPG78hZHBMH99e01iwBzbIcMi3zByREgVR6nKFHtuLFBWW2jG9eyR8eWXPDnO8
g1/sifETBwG2wxlzcidWsckB48QcD/z4tNCAGd294f1QMavV5c47TanGHE0s+ftRsZqQQpf12OBb
nqaOan8M3wIJMtItTpi3CH2ArC9ZZDOizAQ1dSbGEyAhSaVwlPySddGMSxh/YzeHqkAfGYz22xIK
Dgt5re9zsA0AJhayKBPnB7upkBPvhLtfBxWEGqdyx46nBY7eftsOchNa9eggh7Cc/tbzPMQdCWI7
i9WW5nj/32MJN6oys40mWg9+6IvZ+Q3uYtkkQW/4P7ir1DU60T/OvWonPo9N3V+d6bSU7Ra/ezAS
g0UOOd85i5WSTam5QolG7JQywQScSeJD6iR17+bFtGMgGAqI72ptmvLSggyxbYCVSeeDbXlcakLs
kaWubFhd0Be7fWi+toNF5LXK+vjKEmg+s67tA0FHJOQRyHM1WjP1ol2807fJ0TrH56TW0vl59I+f
fPoqe/fgY+Szzga1ssbjJgUH/oI2eb3Kghk9C/C1hR1KfEAiVcDJLL4ZYS5N4qG4JijQCrz+G07S
3AsAXSnZD3FhLp4vKppaZM9YduMFUj3GOzkPoXkpCA7oMuiL5kWZ/v9Hw03Wbi2TozpXipXuWPMq
9UIrjV2KRArP72Jq4DZBUBBbeFDES+n1mz5FAow/zjKsrE8ca5OwB/AuqGzW8pOWy1Ea8jdlR6UW
So29aMN/r/w3ngIANV98rnhokoSD32IKr1v2ZKqg3Rx8D6SQkJBQmcdTEZ1TW/aq2m9Lxgsd8s2t
Bh1KaKetsYcLusJsUKblBK/m6KkW2fOBFiPsBmUPfB4hUgnZip9qdngMEzDMXvMAxORKEi6MDcQL
BeKyYcLHLMPtCfBeph3dIgva4wAS2NyPFIX++k8aP9Y9dRo8Jw4l+n7veBv+xu05hcGEa2/w+/LB
CKB8qk0rNInjl+IYM9vqNkZsafCzE65XTbbLO5EgvSJZ1lwAEwVimmKkWw7VlSJxxcYBy7eRNvVt
xy8NM8jzZzWcMbUs3OrAJeW56k9PevGUjiGuw/GQoBvtGaYvJgYNhvYQ8hjYIuV042gCSNqOdDM+
PIP0pCgt/ApWZSKaKhLMnQ5gCoRjiJkHncIrzAgHLwOhmfqDJe0ECaPDxu/9azxteDfaDSysoxD1
jg8cSxgBZQ+lKXHxmOlX9BbVZqPlMYoMuecR6tKqqA5v85q6KH7naIScqfU8uDYA9eJRwIQlIur0
IkRMTgB5wkV2I9p4JuYfOvS04FL/Reg2oL6YbstZqHLv3t1RUS3YjG4Mvn8BaU2bdSSgV2SrYJfp
UQ4jLb+JqmUVZK8tFEq5tg2Lio/C6D0edcczDA9iHXUlt3nU/5VeCnD6mAToX2jHyzJriMAFLMnZ
JpJQQLUiyfPtqaJgnoEMXbOoHAHqH0MPK0imZUnJWmhft9pq5zxjU23PZBP+a34m26QeGjY1EBc9
fzrB5z+h70lMDM/5/tiR6Bp498ieF0ttOUkbJcq7EL0gb5+aleFM6XP1OWODeKBQ3aa1RP7WqmOw
eaKo7As6UEJn0xRcjj+tAislu1WGNanykdRMuHLHQZ9FafPVtisTvZm0pA/xRLPpyDFv01tadEaM
k0ArhGWOs1ePw5V7Q4Z0K4qF1sW5OkeMzdD5f3mL+ft4A5ykNLib1Thm9bGReIyk8NrqombAKfkX
ydFAJN77ZK3mZExi68JQKcNXPthkpOYIEcxTKILKyTpaME8GPdewiZJZQuoGA6uZRnkkHCUjZGje
MAmAwByMPRokbudjitA2uu4X2DXxDZeO4gTJlYzHyf3sITOFoyZRgiakB507eJTQC6CLIJTSqn1T
MTu39O2QXqrTPQHwgvtbup6OcrjT/uS4vxdtY+JXJP5jxRJeLKcotxG8mAGIAQp49k7GkTIkVdvy
hKJLk+sJIOOkJi8tacAIBQvXl+OTYUD/OlH2g1SZRT2ZrA/mTklxvXFBZyz/4zsZZbhlnSfqwPCJ
++/XYAm/i2cuG2XKOop90639x2muM8WM9Pa6FOeywbl9UfdLR35pRqoUEB8NFQ0S6BMpJj35Bbb0
GZrdb5akZsAttXUqLannSpJfmcdqvbaj2ZkIwBb9avYRrjlkA62wXMi+YeOxmKE0VAn5U1tPlx7p
BVvW5uDXmI/uGdE/sbJ1Z+dZOJO+byCSHBwllYDjKMChjXQUPPbe/mwJ+IZBmqUyvTXBerR24XWV
QUmTJmsCKvkJp+jjkKaRGO4bT/jyqb6ya7rHIVw0XgWHgd6Ow9KsbT21VLnTAPu99vl8+Y9Jibbg
vWEmjR1FUaAAOUOOa/DeTdpJeqOPcp7naMZ6lGtnBuwgzEC92Up4lNOZ8xtAyTsWddlKCwcZjAiY
91rsI1Ij9iOqLiNAfM6Y0833KZb/lDUptLI7OspOmzkoAAaL4PYIM28aK/I31KKBptbct4xFyP6q
oQd79Rus4WnG0DMFAXs71h6sZqk/uD7gA4WwtAbjCEWkhAgObTWtGByP3036L/SFGGlxFdQsIj+J
K8/AxRSe0wySWCLBDiae/9RT3KOIB8rm4bWfiXPcZiC4eexxc31zdVDB4st6g07PrrRQHBTlTnUo
ngq3dmLjoPvIbBB2ELrK0a7Lvu27bvqLbRv0QOC2xMqq6Bq+rDci3E7T9ELVhu+srJ3S9Ij29MSj
8LbeNLBVRhQixqVcRYSEduHBJMGgjs3uKyrBy+J1RxACZHhdyenIqL2jDuMnQ9xLA6/g1m4f+L6E
uXMBNNsLubArpM6Ofw9x9q+7GZZf8dJZs4D2i0ABimeR2BbXKqRyQGRXpUDy0Z5o3VDNxRKt93xk
VFwRG8PL9V3t58ltpssgklygmY4FAyWM6stV2yfUapMUWMxGndK3A24n405LCtK9z9cTj/ZJOh68
+2+F8zd4eonAgmevu19AHoRQJfZMfoiRYx2h7Ad6A6lnPAufKXQwTBKlqPQU3fX/3ZBs8NK4IvEm
sO1VOGiOUpX/Vx17quTJeA4xkDPYU0/E9gb6oX4rtBS92yUMRF9v6JmwIpisnY6ZZ7U7sEBMmnv2
EO00EkBNzEzF8dpAq8BM+9bniFnQeSkfXJ63Hl3YAENfcg/+tjGbcsNIadrn91Q09DycFReGJ10z
FBXEurvtVdk8jtuy47MK0fLI12u0mj+tjCbI9te4r4hPxiA8B5TWQneWbV8DtOkGV0OMp63nGTJr
CA8f6fgohZrO17CzXAqvnkFK7VpCZZaz3kpUzQFac7Lj7repDf63tLbdv83/XH0WHbxYAJy8tM06
ooEVFB31teB387+UJ8u/Xy1czSTB1XQpHwJ3dN9hcz0iLthbXV6Z9MxYcI9RNhD9T/HXbZnxAuPM
NZZuIrUMEDqk9tCRwLcIZpdOoltKjkYEEP+NZdgAU+9JYbM2St6QLLrCUntNo9dY0nDsH4ZP8SHp
zQEjwlZq4QpdKdr607DNSq3xzKAz31mkHBPJoa1m2JCf7OMa4zTZQpgdSSwFHNDdETkKYwsi/JZJ
5CxlkxlTSEZO5AsqHiZoBIeZDC0w+wMtD4bIX0gqXaqDjp/delP+XP9SNTGf2a0fvtxpCBouGmoC
Or0CRxUMytX5BEr90oPyBwamOw2oHLRZQ5G/EAPKB635c3S5uWl3lTyuiToPU8MRh21uMMMrEihS
ltyB3ZX95XXhWgnPfF4xti2//RZMPM1Zt/pvZzjV1+xafvh2giF9bUZOA/IsWQYVJU6EhZRhkF/1
rb0A/eKqD6cSdhAfMW+1Mz7k8tyytUFlLYI9CvLeXoI6TL7xsqTd5az9287GnKk+WutpjTY+Ws7c
DZbL6amKkI9wU8qKWsnYiO23VZ6Zjg4C3e5lKX1+N04Sw7lWhXB8JJY7NKC6iIZDOdKoE4z1CL28
rPWdqFw+PgqARTzI8dLAHgGGk2ePgCbYt1XHMpx4LEHpUo75oBZKB5G0RBepKtzxpX5Z7RhWLbSy
ARp8yWtV/KoRXJs77WKEdKvFTCPFgbSQ6zKNm5181tfT7/GQLQtiVTx5iN3kjBkKJzttXPme6Obv
C8Nimqd2Lu+6oy3n7nBz9AjKaNNVakA+OpvUnZWSmmHrsUpTtL6QwXuWvvlQkjIoZaCI33mLgCbh
Pu8HHhwMBHfbS6MrUhRL9RdkQYB7bEiLFb8A3Tq55FT8/1BYjNphsifEJGp8ykRk2XKrYEzIwx8k
ut0qSjegeQrwc1DwuvbbT0mndk75iJqfaRLXlzYGB0KgoLMYEpVGpkerBYjbZfyuI8bLaD3Kvj9E
wM8FyNgIR0RM7dB0rbjrPTRoG3mU36EUd6+n4q/MGAUfHxCeFp31RjjmV/hXAgwbueHbMijzBOMI
6YJA1paznkjory38Olv9aS1rLoosHdoin4FNKCM1F5iX946+FrndtUlyLQ0ixDiWdAKqsi6UYCsK
LQbXD7bM57vKvVtFOEja8QRMf0zLLAueiL5D80I0fCEL5qdX9TxhNggRW/3nCLOL5NVmxXuFaoj6
D2NLd9TCKPDHiWnlbK+/5ocwi4NiD6fP1VYlcq0ywUAjVGb9XEF7n4iFlgmV/x0OI/zTkGNEpKhm
7VULQZ6GsVv+kNfyPm0qN3tS2EYmZXiTOWZ2wO+OoaFLe/WBxqsz/wdj8+Rk9jelpwxsuKpp/o9u
J1w17+vbJqbPCMdRDV6w1FdSBN5ZwHa63zxPRdRx8JW3+iETCreZSFcgg96PjdCretHMC5nPM8Us
+M6peG2jss8CrR+Cy9GwbOLVVgu4bg7ENcaVcA93BZOg3X9SMOzkaz5la4dyNnwVWm8xnmFkOi6d
OdOQTPs2vmlug25bqEMfHcf+jzCGxHoRJGcmVqY1gByIhVm3M0np9KPhbtyeqn4VBEW1L+rJ1non
VaqoRU+xbqjd1CXi/aUdKXxQhrdQXFWQ0NprOLbAirS3qlbyjakgWkNQeUGS51TG1lDz8qR77QCH
tPT3yLVtaEMKPe4X/b2w+HZZqPMuUWFv9h8egSq0kHq6lQBNaUHtQcp1yilCu3h355kaKuNEQhM/
+tFHtVbrNMrpCBr5knZ1YabKROXO3CXAPlB42PLcIC7TJCRc8g6ZezL4+efkNULM7Y/xIkQC+NzF
kDrFSSx+qxFReRL3yopzuK5vseFV2u+CKyUxG+TKhgXj2UymLrUvtbv1q4S+OtBg2Dbapa9/m0VQ
tgpqQngEb/aX/wkCbEhc3H4OszA+O/y1Zo7SVb54cCXmdnWnY2rpquA657rITAGVzTvJk0FljRUx
oyziRa29zud4P1tEiXYgpXpNh58BdB3K7SFHfEe9XUB8kvGoobc18pbsfs13c+VRjP5mKePXxyVh
ryNKP766v9bqnye1GsCko7Ncpqqk7kE5DrCCk1vIiLGcUEme52mOUN04NclmWX3l+2MoRGvQDIE2
MUIeXjER0FZblCrtrYP6qJQ0ZND4M8RezC4cg2PX+qM7HrHK3cnE9frfRxIuSc51ZJ2hpJhaeJfg
HSX3KFq0mMhIgIV2DfYCHj6DHjrmefJJK9pTqWKI0BYyKRKQU+Pf0lUkECTbdrIfud7mvlKZmHD9
kI6tZquw6viZ9DIRfYrL6Cnmai79iEeUsdRjK6zO6vsMD9hO8oM2d+RKe7qGEtBI/2aR8CYGw1LL
IyxqTpoIlUg0LrMEx1z1bSzTcUswPZvXPerkfBf5evnmIZ7nJchvB1xeQvhjgByh4KBDhTpuzyO9
fdGaDcJmdnQA/6nvdI6/bRaN5jZ/sU0fuGMky7NcW2sCwWo/SOhpcFDTaF3/81HX/roH/7DpEQ1P
2O4yPpM2VNz+XR3IgIYQOlnjt+dxsXJHSafMayL1HdMLsc7cwO2dXNaT84LloGLp8XLnic8CMVT5
KZayn2kLXiSCbZ+eulR8w4suvjlIQkHmQQRrnP+tZsli1Xkrecs1Yhorjsg1dBub2G5nkKFOyny2
hpJZrwioVN0eQ0op6s+DF6wI9bpOB69puQbQLheg90jb1S3Nt0DTdoEKaq8ZCj41SJ0lcFLLsYPM
rZuIs2u2dTh2nbLkzfR3E1lQKpP6rqbpDQR8qugTLY9Fy06lqpBsXVb3ucCKJKC9vzt8sXLfBj9p
qJ/sKM0O3qePERSQDaL+aFEmAd/QPhmgKRADLu2qpO2/gjjiZmvd0RmvIzmGUfZ37tZdXNIPjXMy
yJWbkaQRxQlGcoU24hC81//o7FvfQaPt6e7SXaFsLfx0I09G7nXRmyyAkY5z9eliOejSn7hvBLAJ
R6yEiZXWfduaBPIZIrzcejm4Wy1YiLmdQhACYaEsE1fSaw8zS57StEm3QbXRY+r8CAD55rG/+uXd
86qRImvJvDTbKZ2E35leuuGDaIP20l+qgkiU7RO8UlGZ9rBy1bmPkI86s6ohbMqX8JKp4qc3ApMI
9Y2au/juMqeNw9+xzZQlpFfzCgvl20CbgKimdl1BBgkA9TkRVXYNZyy1+8rQmS5Gf6lur0NeiQ7W
cJPxfLKBcrbrt9jqoqRJmBY4nB+4m0qjSCeKbQRQAmOZfZNNi2WnRDMwOEmNL0Yz+aSfo7iT/Dlz
4KM+EZt769Clkruf/X64GFZZ8/6g5fDJyeB83dKCBQRR6zpIElEssqhJ/hy0sR5LAGnqvGWna0zS
9D340yoSo+O+/2dAzb0ha7WUNayuUclTajhi2NMeUAhMSUVi0ThI/MFCWhhJoLkcbbrKoxFH9slO
DC4YPIZNSPvgbJ3kqW94NN3CtW1PStxZnCeRNNu+bz26zJDC2jF5M2F3J0b4wwCzPKk/Nxot3UpF
4Xt43a0PG+ws50oKTkibfsQX4EGy5NDG43Him/fTImDDk/c4+F7LoFKpVm4+FVY7McxTyAcevfk6
prnWyyYyiWsDuRZZFeKDrNVb0G0gfroFVjOmazCzjXc3g4tORu2WpJgrvC1jMm7H+KUPmdRKORKn
/Wf0+MRIedSq8glfHskdP65dyd053sKRXNcwAHLImUWgQzs4M31bTxW46sk43kLcUIvngj9mneGG
b3eNaoxv9ImNV0R4Y87bwPM6NiCtZFwscaChpi5vFhuX+u+hZojWQjGYL3TQ/NIATAPvAWS58qT5
WVEqJ4DLvr4eUB/UpKGex19NOF08xqkqzoje0qD4w4sxQ0RkA64fuShGhZa7UVTY4Kau4TRGSy3s
lSbNEmoomiP597gUaMOY01HAoiEF/1VHG7/3ALAJd4x4ufL3SJz1QpZ8RW6P3o8vNYy++kllEddD
xyPT0NtDmHf5sIHq9BH8KIL9AhvHCbMKATtW8HHAGdqJuo3cEckuBQnI7BalcBKQMQQMBy0NFl7A
MzJRyzaEkwH7f3IYGwUVBw02ZGp669JX2mPBZmP4Kdtr/GzM7FovkBo33EyRzcxs6mrBtrvvhOnF
JPJbVYgODxwEcDhqIcvoITOY681qSOHQLmy8N4qvnorCDstw0ccQIopk344HsAGqvvJ92oS4s23C
e/jliOwYPHTvc0vGhMsxJGoJw01R0aR1VLkcNjsL6WprZNvgyQzaRhZEKrfOdMJxInCp1SJcKlhT
WlQ4Kg8iT1HPwAk1K1CYiiW2kiTDYl2OYAi0nDZF5VxYlJzFDvfm9uyZUGAXH8GfdeR6JtkR6d0d
ScSAQN0KnCC9DS0tG6rg0CreZIeigLmn9RNKTRrCr5CQDDc3zARyeLZDth0GNGtVcrdiWA8bGrtU
8Y5QEnCjUteQUAuVHKnACpXrjwIZM1InVMgTtUXpiu1XXqXaZOMz3x99dK2zWoe1Ep1Yhm6nk0/4
OBe2o24TG+UvmxwDIVWXiSuTKEAzxorg7jqhJ+W1DJbm12XWb4ziuPuWIA+a+oUiFAD0OuP7YdG4
otaDCM09Y3Uf5craKVYcd5bpln6iZNO7GF+A3vo3+Zd+X6NGuojHxNIMbvzwj6CIaZqWZyQF6V1F
lxTxgQuFfu7NNyDiaD0N5te21J3i5fMyGzMfecyEi6jSFUyBO2mTM06a0zBmTo+NjGPuFJEHxFvN
s87drEFGeftH9iQ+kMBpv2g7SEwJfM0BSOPv953cyXOInRDbA+Ng5MLFVCZyHC2bKnzMYlbNQW5R
yXwIXpJLUUrJIFXo/qvm+BqkjPVJT4wUzHC2irus0hddbem7yrhu3tpXts8m3DAUmLu8jVXNPCl1
qUfWE2mf4Yxjq0z+vJ4UzqMSRRO8X6rOh+JEo4QJV8TKeb/ZzNVpvc1M1unAEg/2NeIp12rvSe3/
I3HoMLw06CcJEWdGMrT8cJRrua3q+vYSObt2+7QQNuw/O3QEnoEBeCEcQ6sAMMzWIK2YxIMrXsLq
mVuaALWjq4y+brJdSnOVHcxUuBE0dyFNMoPKftlq43glbWQsC2qJUNGrApsmmvhe1zOBba3/U/8R
Wyj0OC2c76moFENUFWTZSB0HHtb1u3HjuBdb1Q1xtE7TemH1C8H23VFcBfuIxOC19LKckl7OMkeT
D2a23pj8+WeVqoH1gRsTKYWiHnkeGzjIsnmOWn563B6N0uMAEToZgyrJc0TQITVgk4Jtj9KBsUWC
9hphkyrxRpye6NKnpO20Swq36DqOJzEnd3Ry3EKaVBY8Zzqbn2dQYaUkx0EBvDqefAZIqjYraLKH
EHMMzZQHFLB4a7WFLJ579y86f2C8aY4+AjJAUT3RynG0bPEQ6rPC/2hW22mxUcxuAOmHI3IEcaF1
u1Qdqn+yBcsv+eV1r5QX08438/egYk9kqu2zDilbmS/+SvoEnieoXtY4RPALXVI/TzsGgqTWEVUx
mhOOxUEVkz5dXdDPJ7GjbJe1BHvvECbSVZR4KJDIV8lJ9SkqNdkZ86CW48Yq6P8Rt6ZCJsI54Mcb
kJM2VK1d2VkstaiFJy8Eff7tTxUEHha3tNUkXGfT8vvcd5ud5X+O62Y0ZbvPJ2Gg/M9tDLnBeewT
RULolE+MVbYTYRnWElGeK1QPiAWkXI179O7ZNSc2vdxQNrKQ0akNXBtiiDbr7r3uA7RBJVTA6Goa
U1/w54g4vvLfBthzKkujGjoqQsvM0SBjLmyW6hYDuEqesO/cbATzwyImXZmGXhtgVijTqzCEBbWP
BuHeJCCn4w4qr1/I4drLT6D98vYU5Ba7yDEgmijJduFnx0Q/4VOSQrOCc7bOgvuqCTvNaUIRdCjL
3Rs1SL4+ytwKOUoUKpjs2cdDBga+mVG2WpD9zygoLAVJbxwsMbBTzCZyExvEEU6XwTC6PNjmo0cA
X4ugGpLupOvNoxWCJUDTHKw69rzfkZyfWC51xh9q7lDZZg1/Dfn0TQaRFtVXpt/eaEi81pTn8yke
OSWAa3fO2VXQs+NJzU5prQ42hBondcYQ/pv5lgS1grmsTy/+tUIzH1P51hm6h2J/kagi1DKmcuZy
Pkrfa7CxCLesOpNuTmjBEOrrEnGJG0GQZqCPpoQH6d72nJOjDMxoTtL9i8hNNQ6RkOnY1D1g+Ury
W3q12OKkMWB8+JzaMN8xDVcehP9/gPrKs55FlMOIPZ3YDl4C2/1wFt7urwQJeH9i2OyOPgaPoLaW
jsY7N92kMdXz2STWH1QElx3tB1ZbAYTWKVCM4AK05y0WIkmKYf5iYLo5G0EbhVGoOrcK6xe9unDp
Ca+aEUyHj/fb2z4Tq0Vixemb6T+l9ZoYSzuvxiHmtAVNAp+kupPkPfhX1PPfkVOyiJCOCH/+TF0V
Nz9PvFxncXZwwo3hXZFRn31hscx4jOSU4zNlvXAVqIKbJkaFj7MqF/TX5z95aMF/UAFHXz8Vr+3z
uti0Ax/GLjt4IqfoeOTNDRkc7z6HvupQh3ZfggafQXQdlOVAbZEPtXUuo7FgPIQR/YEVO+lwh+gH
9mxoqSIl8oKVpzBeHZDL+nXTp9qY5br2nhiLCcww+UZ3dABO6E4XbzbYBau4+oe+oyWZX7eE081U
i0OUS2CHon9NUQvjOv4QHHXaTjneeGBD0fZPvL66TgQSswmc8HUDrPOIKueubhcWOBD3NtmPujQ4
jQNF5u9MaRC+hZ3fccpFBBvgfRu9pUj8+m7xq0NTPiTTYYXPa7xeN2+Y9bUE5BPEcK5G9oSM44uv
U14vXSn1I6tokBVVqoAY1fMnnhTFCzlrmDQo0z6hMDGTRwE+vtN2nwBIvS/e7IjQRgY+fdAmxSVN
OkcryiZu/yCFDfqaFMNTVOy6vjSbbySU+2jQI6XUWSIoBZU0Y9Gf6PUL3GQoA6kt+Aj6yRzImp87
/0MxCYRBWCETBWKaI86lB3zye9nCeaWrie2h193tE9MxjisG6Bd97FwpdRZxtwTJfG1iyc4A+Ll2
IaveWhShhfzKNSp/oemEE+1Lne3N1s6fwhz7zd+u4YMzdDPRC84Wzv/vuFCH99bfhfzXm/eTlRxR
2uVjMbm28RJa8zTH+NMlCu2UaxVJSfHvDjtia6+NSpGvaE1zHEKnaJR2TVabrnGBuZhAZBjlogbO
dG0W68FZf+ayHU+43zrm8PDH1xxVQV7f7d9wJZl9asOs9+1GhgOBf7K1HuHFXMDGog656lEzRWTs
oy+qez42KXGhPJlOxdfHbC8tFCo3ER9SQ40OC6sS9LxAjcUO+qOqf9ZR0ZgO4O8trzJSsF1D6O4I
5zW5BOghe08niJ1V2dDLZMfb2R6s2Qb357WOXNAtpEtZEzC4YIIQNymnLWKXe2Uxo+MBRb0+tGZZ
30olzIPG6h1o8VMPl/uSA9dPFNxqN58/faP4tA0ri+0qIrRzI9mVO5pDE8fDzXGAeYCtl7dUNL2T
xFMEiJ2LOdjRH/l2QinMYpC415KRUDD3VsKIEVph0okvu7LFyTTXHYHOtOqcpfM8brNHWBK9VNa6
Jt7corGUa4eDbypoe89ORFgUIlsBbvEG9OfP8pcZ3hlg8A9KnU/K5eJtasNnKX3EUck0GTAIJeNV
z0eqYy8igjwRRD68SfzfZV0FtzMVSltRTjj8JTXj5RpW31G2Cjm6ovMAN9zZfvlzlYMwsSuCTpIZ
eGJCjCAxRmEhoWPD05KNvXg/ftHAJMt/mn74tAJ4MXt1gn/UMF17k+XZ4ULbpx50fysDjiro73aE
yzRz3OIxwMTTaEFL25raahwt3FEylTKot8tsaqP9NLGOuh0HYIxhttk0dsw7uPV7AolgfE5WO5Ct
O3gXBaSrjtOyEuPX//I0oCx8uNiv9lE+IfOupTRlETLXl2ZOR5By3Ntt/zEp1H018t4VAE+T8R4i
RJ9sqOJFtaRi9IRemUk5Q/l8zsrwXo7whuDMCCs7Ssf8GbW2Wdl38KnjnDfAOQX9evxXtmKgpcXK
GpFx+D0lJiOGW0mfK+QzsUiOZACj4gG6BgSMT3PBvVyUnG8W9mYxYTtIdoTHTt/pZFhZLPu/nfh/
HUYd9SfhO0xpkkaCnIajF5VeXe1kA/eOSYBcmhs3CTBIm4d2YJfMRapDA/r64D/8lZAQyGO0LiED
sb+t87hHB1iD+OKxDBXj/YIhQXjdClaUenHQcAq0MQ22Z8rpREoIWX4EFQ+xPNcGesOyAwKnGc8x
+hnJuy+DfmCUi19wsICJ/Bw/aBbJg2rouNMtMoTrTacJlsjjj13h82E1tHDFl+EPNf2POVkYcO4e
w7gRhz1qRlHtlUowbGIc9ljTx6d0cy/uficlnBt/cCIT7xOccJHVeeG7JHkjPCgVSqt6IfsYCDvQ
WU3M4IbzLBsV8i0iSM9yoCsK5wsW0VUVUIt/QCpUS7ybfmNVhhKrfkq1QZKIULCLjtY7nM4C7nVJ
NsFLJtz4Avv/24feQXjmB8VNGm+JuJw6xNMAi3ier2f0R7raavtfDU08W/QxBQ4beyyDXDnY5s/x
sokKrwRTNeNK0nR9SsoKFrstCKTbNICv6IA4Bvci5NxOB2jckx8rmakggHWwGGkAp9pYvzclX983
Cp2G/kRV5tKQfN2GIIbwnWU97F3kmL948sitbkFg5lMnQ+TygwN9byCjjIwxjzZLx25oaMHLTR3z
lDAn9QXmfIMsmYQlZOk6ZYARSvWB9VJRCZKMEPlghrPdspiKFSlBFdo9nA+GEUImgrGXWgdTfz3b
KqaJDcIf2+/AStqQ2+HznQ5OJlhaBn7ktr00e6dr/dVXXKtArtcBPEDWVXxGnrU5FclN2s3usAYi
LHrHK/R7c5EtnemOR71O5jNl50qHK2BbcTK6f0azfavjxWTRnXiHxKA3WpNN+P8F2sE3+8TfG89d
AzPhdrPC6zu0cYdyaVS297V1v3inqG8Jl/ynh8MJJRbFWfar+IZ1ifQQ/YqEO87xOScrBVa7+qFY
BYd8E+1lpOhqo1MDFNthSGITAHzlJyiZHyPYh50bliRCgTsz+c85hsx7MJRoVdiibMF7CjLkng5G
0zRmOnmVqngconACbYU86pmo9ZsXwfEKHfXIYyDIEDIUoPdcpOnHIh/K5435GTdu+nVsmGkPSSPR
C2x7g9LwC/ZKGxvlbM2EX9U/OnyfdWFwHxT6AZ512y5liKfT2kdBUzg5weFN/t34hm6jcwuMaFke
JwLKOVVhOxdnf4WN1uLLQji18WfQ3ZwXQL7txB7HNgGzgHklU0u3pVGk8At3gF8gWBfZ1QQfgZDK
KHmcOotBIYDB+F2Tdi0xtHzxl1goyduVq/wDHluakxH9BIxKYx+TqP/Z6uDn1yvNJf0FF4jh4Ze6
ICSQaSoLA2BymdKvZj9GlBuwNTYoAF4GyJJmtCOcWNEBg4bBTaLVtpv1JancTZgWN2bPF24GTVZk
IDm1AXzCN3WEhFe6I2gdsi4Uh5yVyYOD6l+OwNcY4V6xh1KlgWM7YxaiWv7y//eXVQ51M+0JXxvx
ewbGEZHmw9cjtiMzyNcIlUdivj7KGAm/KCKlTgj5YCu8HCEylh018WdmkzGwWsX8mMoyYWj9PKOD
MD02ksW6lgxW7h9K9bCpJ8mXH8baoMf63EZIHe3l9j4wKqzhm/7Vdh/LH5dzTm5kL0E2rB1RDPJ7
A53/+CfXYfV2BQ4oQa19GW29kgwCU7lGxVq8580oAxxJsmqjVOyZqDDeFXm+J1a4xYub5MRY18h2
Y6wIG9aehVmBMRy4S1+WH2kmzuoPoZ31rAkMlDLxoVn6IhaeK0w2y4hf1Q1gX8lg5xjaDahFulLJ
npjiPb5yjYM+EEzyic3SnoZZxvuuXZMovTbCr1wLEr3EDhd7G2TfjKIjbPPZJWb7J9Xr6DXBMdGI
jdFDSw48q8REfvvkusQ8suw8vSMffKtf0MP6VOFn4Vr3qAmu6HKrlf6jJ/kPHKZuaFMQ+5XunpFK
y2uu2VCZg9cY2/t/f7BEJ9qJmXscz4bYe83us75ICUmB081CRKqdCWLC8iaoMuAZ0jpDcfUsWGuG
SriHVU3QdBP/pFVztpWXUAv4qb+lSSQQ2CNbp7MegTb2BErIyaOoHTSPTSW++z/o+DjhEWlQ6q24
bJdpjEd33slaAd+xMo3icmY0bvki9RaDWhb6Tq/bl524STbsbJ3JnZK/vgsW6uj03vOHXTNFWWOn
enIVJfEIAnsmpQqT0vxugKgjoht95MNMh1uncsLlZLor9d3cC+02ixmGYrfgDCJ7d28MvrmRRZX6
Llz7szVy/5bHekmmIsBRtIp/0oE56MtCwDud3uNAx0Eaha0ZXJpRoQ9bagEuj2F1rxkRCd0FCW0A
21XWWWxoxnODv1+sBfwnj0ifIz7tcEbRl7OhVtFq8ph/W2ibTUcVwCWFVOeI5aOVvTTMMKamc8Oz
NGowVz4Ke+AGLuFkqIx55M/3keSZEJcl3xJTr9wlHk+MX1kInVmmVGkJOw/49jltQqKcEU9jeSFa
0DLVdLHKWahlcmKF1CYnIkNfdQpuMg4WU++L6dBjIFdA07FoNCbNN6zFMmjisNppZgWP4MG13ox4
DfCz1ZoklYGPwuslSR2j02a5sem69xy9FXSG56F2ATU0aSyWNOLZS0o29Zt+/dVx7LT/IXIugSQ8
KAXiU+L8/PcuLf/a/al/N8vfflq+/xO5xMG+mDq8tlr/q1McDQqQdOJYZcs9UGfTMTtSN8YKNX2P
WsnjiAq/aEuNryS4yBwZsYAv774Z5sWT1A+qQQuhkcx1oaQsUxPeIU+AAC1KaGdj10ZjNquD+9hO
aqECT/ZqNYjEA+yK9yrS7jWceXesfpj8iLSM9LG7hWFQNXnAlXtyE4I2ZjNIMZhx4ybbReRrAafY
geF+rY49SOGJYftd2fqYbZmpSmM0LoSeG4uHa6GMMgsMJ70+Pr2XyvOXT4oHcaoUp7aK3EkJOJg8
uQsMJK1wLwe6EA6NBCYh51+kkUfLaKTQ1+pNxQHfxz4qBUJlQq3o9u//VMq+N8qdatNX77VLtsKs
+kQ6yhc5d6xAIKPg+Jv3vrcG+COO/c0/dUhBcAKQnRsJVvnXgojZxwwrAcw3Jt3zPkyRC4QzYhGx
6/0/suHWaqaIoQNkCBmfmq7WUz7LyQ9MlnEKgrtcgbILf5vBuDORQ5enBO/Oc2X1mBD8HpJsWqi1
UbRrz/rK6iAUNKBak/cyg0oYHi5iTHbGPYuiXdfSL/IPeFfksx1l8D+TPxooiZytJj7VZDIY5a1R
rDHXtyPfsaQ3smm6sbAF3/RaLzreJPusurrCOFRsN0J6IdQGgJ5t96msXbWDLVFhwKmCDNgpuWgN
QpZtVzbkSNsQBLs4NVuDckCuQG8fAq7DT1Ca285VGFlZN3LWgt/9L2Rq6RG68rAWiTS+zisckEVe
ZocsFPkyorXPqWtjAPb0ftI6Ga9zMdwK1T84cBcukyGoEvOGNe64qRPyJFefvBOOBlP1ZU2h/A+Q
PRNSSipRWMVi3lX4eSSvveifeu84cfIpoNpxZfMhzUjkX9MnHokWhu5VF55jvFUfb5HN5qUZeism
G6VOTR1fwCIRo3OPHeb+dDE/AP5DkIG9kye1h4npy7X4nC8ZdaV9Ez3x9+vIDgJbwftwoojZmFwt
8KEopmoCAW5lZ69rEHwMlK6+A3BX/HiDvO0lWOkArW146EU9GMEUHLJTl05T4NCdYcf8LahNc1wJ
7sbmHRttelFiv6HDMiokDSPDGuKfoRlB6w92LAtKVg0MR1T+GTrvFJGuq05dDXE0RypM330KU3kc
qVeo2JQWS6sehn+DXq3M18yWdoZ1/CoMw0GroViXpkmDUgHRtRvdvaQJOuJ0DZIQaGWasg7y5vbz
iK1JNff5lXOYdTZj9FgNQdT/NOrllJ4FQiR/Ye0FgKJua9GOHvZenY7giO2EsXST+7ignes9PNYx
f+iImmNuuNGBwOPXWeOZImG8t0CYZF/V6mfHVjHBekqRasiHzrnNWRguwfgs+GSNVW4DgUKf9tu1
DadQu+d27QLzKd5IwOCdwAedUEsymS+tIvCpWC2zP+RASwkD5ykmQhsunIIsnmGlP1vLnssq9SBm
FiexPuxo7kGTohPcPpcupFKz0abv+phNXBRXGOU2Fq/uDT5nQUOvB7GKgVHD+Su1glOhxdAmRM2C
OQ4eHXiXLZAVzifopFRkyPblMGNsrmwtqNfKCzr4yF199dRc61/wfcayXqIWFEFAzxXRa/cn9JZr
9Z1BN+XeXWWglqII//IhAJ/9Wp0KD4wEvhBOvVvolRGevC9jOevjH61P9a2FxHHk8VylnKERtQDL
jf53NC+375qqh4aXWRS4Yh8ZISbO2hCkMFDUo08u4h/suQrEPCqIxzZhmFUduEdTAJppVLG6RMXZ
Tvv9+F9A1kuh8KaKZjd8rrYkwzY69gKrjAZlm0wLJ31KhHPlKQDNWRr/9cXReyvGNsv3XfSQbkFh
Fhc/MCWGVo25n2S+ELZqzQhyXXoFFu4OxvtMTyAcR/UCEfKncHEDHYZeyo5Cg8Xt23hdIbs28Wyl
zMRs4nl3R5pV+v94ydid8qhHT3meJqaHErDJUl93u3EnmVeTgYnHTv60nfVlVSAwX7KpPrwjJr+j
SYmTXr+yGklp3jvCHT7GQBAPcQHNXODHhSOXb596J5kbShS66c0ILuXSYbmm1K/CYA2WIYoXFc0W
7NF0zhcOWueuzEHgqbjU8pyxRD69XLZEo7b9Ile87Lj3z/gsekL6Ayglhe2d4BA3n/5kXWpny3fJ
Bk8c0Qs9elux6fA/uU4MCmxUlhIa+NgRJJQGBEgYb43d51LsUNm+fhS5XxAnHvf9OexGA6O8FoHC
NlB+uFDmlPbA490K+KASZUHRFR15c+st6C4dYyKtgqZy7ci5zq4Z+vjCV0o9OnOmRbGbN16OeRdH
8VT4OlOQeB9vs9wFenat31yJDrCJENGArDJKlAGQygHdbbNZy14zSpeGrWvHVwBU1SmWg0ysF/T/
LPOIoTuVilX2nL+7YHwZaHj6Fe+OV9U61LDDfJ6rdzoisSEXaDaSzz3nCdcqWCtJv/Rfxa7bs1me
/MTJfxxTQE1bVhHD1EtzsBDwpTkJPOY4zFjIQvCjIXR+6md9OOpI4FUS4QwiX32ENg1wH22SjsRA
6IldCHvhF8Uyvv337yq93a6g3/BiBt8TJ8g/F5RTnnCT5n8wgGU3LxewTIM4QSc/MWvEt8ew7tEq
hWV8q9El7ufeYYW5uB+PB4RiNiN2rW54++6yUeFiFi5RzYXPI5UHPKlVe5kRXvHxQ1mCvVNSZutV
fiJVF8KhxR/muStApa+ERC7SVZ4R0mgqKA7/0sibuZG3krhyMa5g+AnGQVcMEwavRegS6ZDy9ycv
un5W0AaEqfh0uSpAAcqaHtH+Y022/AyuzWbFOJ2TETPsoz5BmpYVJLocuvPrX4zId9f1/CZq2Q6N
9Aceo/sZW7pxhAJFt61OCiQ/ZuKBPO431xlRja+2/btKXb9GvM71mVuSQawLbPt5lsQg9QFgh6YT
LHhuB4714RtDobVhuyDm3YOpWTls1dA1v+iWQ3RO11aMml6M3ZEUFl2uAcAHAplzbLsltDX5qqLu
Agmg15ViG1tbYTMHyuVIt6bOY+dexsuifBzJaiUS8t5nQN6i+sUrZPw99fuXdXVpDCY/cH7eREWo
0P7sc0Ju4gBZm3DyKa/Jo+qPpbFi+j0cdYeP4abFPiyHMXE5Kk1PQkhdVDNVogESEcQeg755ZXS5
xTwxCEgtUy+QhmPj1xbRURgtnU2A01QmcZN+NzvbWou2RzaIoAMKUgLSNEoSjBD5PNgysjoeEDdY
v2FFRO/dHZcy+UY8ccd+XjDl1uiP6j5i8ZoaIaRb8/BGEnjpGAq280oOF5vYyfWrQJuaqmzLxr7C
lyKk209ORYc/0iyh5IubE2fZ3BTCSHRxRMDLSqfxBW2IqmfE9FyDXuyPbIT8pG8uIkSk8JrxadcQ
YVWx6wodLLEv8JVc69Xsx8dDaKboHYyCRfAIkAnQnATl9IeGc8iU7yLN2PUFMOHr3AYNGszvB6G6
N+LuxU+Dbm9XXQfMx+/DECgnE6cXWdaXISG1tOZftchR/b6ROv70Iz/H1GszSleHrKyqxrXgSxeX
aVzMjRSG4qAZlMqorVIZ0rgThavaM5BnLWMygL7bGqUGkle6ULoDzs6CIMMyRoYZ8/4Lqx2QMDX8
QBLNGip7pUW4MPZZzEJEQun+Tj5xC8WDuCfE/LwoAP8qaOUO7L+V6ezJZfspZ0HWwoELpNmMq2YC
+y93tgMG6JgOSKo1PLrrokVJb8Pr4GPtntRkmIluMWLrB9uL/iq/0HeM2rJFGSe1Hmq2+DFriXL8
QGwPxNuVbJP74Bq9hK4z2sx3ghx2oI8hA3zCeWCXhkDG+r6aADSPhVeQcccm5YGD1jaaxHD1Pxxe
pcxijinb18qqSrcOpEQFOzgqAZDtuqVDNG/ohQyOnjpANUU7QKRcFPL4f2YK4mKesf4pj25M13hM
q+ckqJzFkjQZNkEC2VUtgiMP8L1Wem1Y6heIENoN+jCgm1Rn0MxH0pYMABsdza4LAjW009s6Nwtr
vmjV1ZRv9wTg0f9UMPCKYKAD9srCfA/3HJRt9DgEcjGUR2QDEZFkGi4LjOEBtelGYAU9KLwukMyg
VLzzBU/5XPr1Si0ddh+fcM2bF++WRONBHhycU8Qt+ieO2YGSDrqVJn/oT0uHxjTJnYLNnqKq6rvf
xcYliuamB2n/0vfFg02RGUHjpzc2fP43DG79wiTaeZquyPPHGvElwOuoyO56L1kf/aTA4hs/oV9S
xmpGCa1+jJLGgb8GSVemfK8Jowa8tyjNv9MNXDFAGodcr+2+h/M251tIMT5+Dj86oc2V9TVOIARP
hKNvyRQlsZS3E6JfSjCq24di+TSZfJYxN3n9dAVul/7dBjA8hLbE8vYvZbECyM1feEjK+s6pmmfx
ZTozVe30FKiudv7YVRms3wSvbGleujFf/dLzxAqURu6XGBpRu5jg5sk+J2E+oPwZcHTfQNzXss8Z
ATIoBN2PNIKgAvQi4NUG/lagjE/GwWpTGEcHVpaZcmJ5O1RiPHIilRLLNKd9t+Raa9StQLxIYi6k
oBU5uWs2EZXUvrevA5qX7bzrRZ3xcmoUcJZymImaolM7FEh927mpu2NwM9Ctm5UZGXnv2BkI25yw
z+FlAneWIYSSEUHrLwL97O+FAWM4wkyMDXqw9Y9nb6CnGN9igVISUBXnbPxXDMXAWWg3yldko5hy
yQxjet6IcxmTY+dXVMQuxkX3dWHYzk6lDrjbqV75wTZ/bZF7SRZRqwzsPunQE3erKp3W3hk8pa4c
mX3/CMGb8tM5wpIqa5C/LYgpQ+Ibx0C+c9x+p7+4lUY/kT16dVpLUQJakWmtNthzg6XGBJ0Ydm1F
r57gXFe2dKCm56MLClFE38jT2wl7nbESS812ONr3QX+L8qg/E9DvEAlKsw5waBjfL7C9+bOyE+Jo
PJmrS66fkt8oAkcjQETlgLi6wN6BRAI3KzVfyVemdpujHg3brRkkZcfeMHHEgJRGPAxgLRu6b/L1
rmwW376yX1xSFrMTjx/aw3QZb1+KVGxh+qLSBSfcx9i4UTdfpiNQpkhxL43l+CoU8WPaknloBd4H
5PgO/da2II81YsJZjj5xbDZXY0cK5K0mRLATmq2sKuOtmUjKACKezbITkWHuPJjiwD18DI/IQLtZ
CcMjIamBI0EoUCWTGo/E9tWAI7042dhttCamBiMaZ3nk386OB5cflpfi4y5C9jtruV4KX1FPnhzU
17BzREBMS2JGLQAzgpTH+k692JowvfSFeoTgq3Sjnmk/1d1xUVqxFNWlK4wzwKfj/sCmZLIMkhzE
K3YRJTLIspbVgHY84OOx2mfFV/1IMNw5sm53IA/AcAiRs/PTvnD6NlsTw8O+yMsU1hi9m0G6DBTS
Slpisl+5vb80S8/BRTpqYlnDUdi5Ecvyrptadzp9pLzSQ+DdW++0tA39i39E0uHP90qhmB3RFUhs
SFnZS+HUKTJa5SuGCAOpOLFoaX8tcQWAGiXD0PmpeEHJCctnuEQh9QUkjdeRD0r09QS1z+uDROg/
OhhEb6L2u3DT4XiSy34uchsGpRscK9mo/2CpsCWWLW1q7Q9llDG/lJicLlgtVd63TwSAd21nGOyW
EkJ2dZooMD4q8TY7CU3qZ/aS10zrJOp/9cYZhprxjxAdfkXXXGP4lQUXngeXtMdIKf97pZuTA5/E
VsP8MTC7aBghs2XMRRDTOsIQYW6UfPzxDLqtO+oafXaya6D43xri7TLOKfbr/21c4QbB4gBg/V1a
RFDpTFP8w3y3YSutSC4RUwfMTspBFPoaFS+dzmDzUFNrl8EuRLDD49kaAyJWifxs08feAlRCCJ+z
hHziKMLcAgADKwo5RRPd9v+Fl2djRcIqOnZFZGT8MOl8bn9elm0K4cAJFDY2RIhHSqdRwiK3szsU
Vaek3GUmbzGtS3hzGw0gYFeswQ+c7Ly3gSBDiOnO5+2QjEpF+BH5SkW5XTIpyc9cAeYtkxC99f/H
1dZl9pff6n9r54M0/nkXnUXpDJznrEBZNdHUI//5ixCbtqowUFmvG1smHl56X6zce9p5tzhWhI73
XXqf9fHaiHqglx1PzN/pmA0i++mv9ycf5TCBEt4cLEEHa7iyXhZJnmnUPyq3KXP+x9OysA9v/7l9
uo7CUd1iYI7w6wV8mWL963548T0Yyfluaw9NUgDxTXRPmXkljK6eVPDZX58cBz1Nfs3CYqmYKB2A
cv6+qJhbkf4pmxkAG2SS/i5CDo5PuJf+7vUhiICmWtCoYEDJrYnOXT7F/B5BXbnxkf9DeXqNqhcq
LNF6yVT6SnJ9iYYshr0DWC9ugYKryg6ID96oht5JcoxSKQW22xU/h5vszt3z1aesjau5Pn2RMUGF
utyowGl3aaAY8DenV/YDz4vt21SwaI519WU2KCRz8W8pLvOHFt38mBJufgatLXabbcShT/tcdYFB
D0gpH5xLdL/7xuH/IHBn9sEXNs6hF1ASLaR2IeDROKgHb/A0KM6vAB4qz/8SBk2QXNBe2krbOMJH
mKxhMixWC2WBpBs1edKLckQ2ULFl7ZjshaHrkRoDylyiOJ9vR9wzThdz4rCnEpRB8HrSCF3V6GwT
sVRlEDzf992RCEEMBiRbU+IQ5JAfK4/7FQHx1iNdg6ptKNPFH2ag3Eh9xZwHdbsvlJEszeUlecUg
c4/w4QDWZ6SyaXjPGQYB/gbDDvmOCOx3F6s8ASC4ssty93oMz3Vulies7J64HC2yCgTiUVTku5B/
2picAr1QWkvTfx+9eLpEHapTSDq/xaVMp4G+7PJetWakF3GPm5dd6Tt24rX80mILJXnKP78AjWZe
5ynuiYXJgCvUOtwSjSB5eSlC92G6sm0Xtw3vz4jkGRb9TKHVh8HgWqKlTDXIHMEWlN1ojY4jqKBv
7BSPZ/4Kp++pGiacgtzz48O9USELSeQikL339OEOeXjdTYs9apP+r8BnZOq+Nnbgn8ZLvfSlknxE
SVne529vT636ZvGFm8lWJoqvXCIEr665J4dWMPA+JVgZlBSJZepzk+Gddi4zckJAN1imwEA7H6pz
o5h3fGleh4NckeLvXiAzl1Zu4RPeLo4E5k6+ty0Vl4i4eeF6rElG8vaQQUl9Cx9fuhtvnPGsyqmX
RN72hq5e35A4RzN6hk2dmDXJwJbrSz8d4NN9tJ8ltU0P0df7yxa0t0TZRuVqCD+GIYWfviaTkVpn
PfvZUHlUdr8KD3ESK0TSmv73cSxrXr4SQpkPJsAyp8Sa9jo6XcaaNPH8RFjVgit1CRDclFSIz4Cl
fcaont7df1ThN2K1kNk3h8cGEZ3FV0T2AfRlPeBdOR2nWB9KfkNoX9buT7VjgGcT8Ue/ddohgWUk
jqG5J1Vv361218xKyWnQ9MF4UJtkMrAGBM/wHnGTuZ4B3jYqZ5O/flkVCeOiRKEKCcGLSv6sreDO
aE59b9GjifYAIsyr87uVW+EaaxfqxJ4z+JZEPOXjQ9WUamixIyjlJeY7UmrRCZvvKIjayd26/ogq
C+b6FHs0GT/gd62EavxeHz1xylYsFi3HV0hjY5mDCbx2H767n1D+DEO1W/0HqjL5j9b+MRpaAdXI
t6v9eDl8bWbABYc1PjypKBB57fee5GIrXmfSy87O2xChVXLf0LAp1i5TX17Kt4ilrSs0WarIXekA
7LjZRKpJvEyv11AfOHlRC5Xu1aFrs4Bde+E1WusqHQlpl5nBtp+JKp3zUUTF8ghDyQIjf/PwyqLK
ACdf9BKn9grFQ1uctSZ6JmYddw4J5KCZvB/EQCiEvC/BZ7gOA0fE2K2q+ddklJliBCyBn7fyprRB
hrlUe7sgzmi0Y7D7MRS/LW/dNqS2rz7fYJYN1Jr9ovtNuAyAr6ryLNCDp3L2I6zBrgb6SfwBluES
/fY+X5KHMEWcefI5G/JOwzXk5TNE8Pd4fOj95LBBloYDjeWiRPw/Et2j9QsYaukQVVU5uEKtJNap
aHwJQBVzBIY4UaSVmbnoVrs5DA9QIcwQkUEDd06gNVor+dfATGBm5dp1jt/RmpDwS36dP6yEC9WJ
uKbCKCLKtxbV7c3V0/sFJcwaS7VvYCA1qAmCk3TjmplXGfHeeCJbTcj15QbUpyGLHAf7idZgGRod
/9rdDOfOpO0RlM9xQlp9sKz1zjekA03GIkPj+jG+XDf3v02da922CydkZ5Fh4LIT/QJdsg2T0QD+
KnrA4nahU4LsppwBXD9LT0wvlMIqUinTbuhtjS92GdDaBNJQ2f1sFalwUySEUIO/xFSJTzMXHzgS
kg5ogicu4sCy8+u/0lg7dtEht7IvSqRV7CXMF278U3GiM+JpGBO+O2D7/HyeUVmQG+foCP6Dcry/
g7wEc4srbaqHIzuHD7fUGkAClV4vyKBMZuIfsBH+oykGX1ryJhfFbBtiWD7nNUKe/VJ54YsPdis6
0uZrP1gyweh3ts4VkpqA1PzGIACpAfi1Zc0qD9I1LkKNBnQJluySla6rCcOJNmEGrfYig5YAx5pl
T1p8mdMQt+Ck3W+eciPshUhEYO+kbwDYApCWBMX4WO5njoBEiRK5HZTlNZ3SOY1TTHgGLloI0jGI
XWnEHi+Uz8S0H2EBL5th7Y902vColDoJ72bx0UTqlSdMvZ8bit+sQbmsnd1L5R9Il4hynklBKTuv
n3nftnNzv4L8rnm2buZgQVzPksvV/hOyR8t/aJ/w7f1oNoCnR4Ca2Sp2La66veB115XSTJDgqb6t
GMpmgFbPL9I+EGMfIWHakMfQ3C6rQ0NRHoEAAzkdZSF+uixmKSv2J4+dHgpKwah/6NU+Iest/Ovz
/MkgAomBNm3foGDQbaAASP3odBJHssTdIQDq/dGEdHXtbLAzPAtYA7F9QQjjA0fLtwdzHzRucbAQ
DAyeNv3quGaMSUHVP0B4wO3NNZRLj1Bg3hasEaZXshmDvHQEhaZFUGs+vDtOPRAp6GaiwYAHJiff
tRC4gkR7M6//LFWMyAXWfqsCfhaZtX3KjEoURxldWPSoZ1MP+H+hJtd5fqX3xPBuDFxzVCFijnwo
bJVPxWn9IH8baHpCPRwDdAqjS6sLwopgLcRD6uoE7HhgGLBOhWrepeXcyF5mszPwzZQQZp0evQDR
azUmrCm0yQjD3kCLo61Qyf9Fx/UuR+6WwU5YRIU4VUTCj/xzeyfjJ9qJWBKR+NnUnz2EbvSBMf9V
vUQRdlczdiDzw4LmWpG+NZ3EQegJn9tf9D7nfhEi5Bnb+uspQQ3aAQNx3eRzidMcoZA/52ZLDyjw
vdsRXCFIUE5/8a8/TQujor5cN/C8aQX/GdEKCgKRL6RvZKcl6Wdot6l1TwDqrUWMK7VJshAXe+0X
13Rxh19mQswaYC1zRFV6VOLHbJziSLPGFqDzhFLsZOducFjAWChNfjGTdT/P7AjCPsHKttM3krpj
/wuAsjaZMq6YlXNA5uy71HOgNm3mG0dAugW/pzuXDEgelI3ulhM78y59LSZnzbcHX+bgmyC7gABr
dieF74GgfyhVk3sxK0SzI0z0lNRkneye0yWWmRjVDZJ8x3sT1VbQPGj3K7AT15bUGBaV80qmkgBb
m5XDb29sdwwry0logN1CgpRB6tkw8ksBFG9yu0znV+mrhT0Jetwu1iqgKmoKGW5reo0GG/Jl0gh6
DzGV44Gm5r0Uyo2o2k3h81qbWen0w/ENOdnI+V+GeZt6+r2Tl4uFHd4EwLI608XJQ4kUnYzJ906q
+Sg/soMDc7KVrgJCTvDCMSTD3+O26Vq8yTeWxYJch+eGPhsmr9rOiLNm0qzcMbQAQnyZIj7Fd8/H
R85n6Uq+9aV9z3PcJMNh32J0g7jBfVipUlSubqPQ91/ksVViEZ/bTPK4T+LozCFL9qfQW0qHQ2X8
KqBg/+EhSgEbWcZA1wTBi23Fd+15XT7wkshr+79cMjbMfbnfkOpZKqwspQRw15Gt+ed/xuc/aUf3
QwbzIiNwHwvJBGiM47KJDVI9JkwedE72NO2+npqGY+RZpv/Hgl66EJro0lWHYduto2syTKjbT8Vc
aEcO56ZC3zONbJHPs4S5qOvJQ+4B6tbPVVtat1Bfz4/qnlcjjabeh0rnuLXWRmPmGX3UEVCzpRbK
UCNBOLfe7k4jWqFREJBvYDAYQkTLZPdXpPNI2XCXWd+T9owyY4YpEGGGAiDw7FNnpvopPH8QJwWr
OwDJVzOm5KqjsDfAX0b6W9C2R90JUvt1wpLl1H9be3MBDGboC7m2TL32A7dH37khObOHGNeWd3/b
JCxpTWlqGH8TGAlXGLzSQV2IyOqsN13gnTHqxStL66dhCmuWfMP5dxcyxhAQnJETxMrie3QK/oPE
esXKDe0kKNdsCkX01JxAlxdI7nJ5xgvHG23IKMdDwKZgZYWL8AriQxL5lO/lMKR74/JeI+533j64
sNzPzEhC2pdKFrCaZXoLOE6F5gC4HZ/CMah3yZPmefwOYCmomN+MxvjyPuMLFAUa+1hoEsCKSgYe
wP7nsx95gJ7DAGsQNy1iIVqVLQo1Tbsg2Hqm4et+uIsnv/bUE92AIvNVBQUyYZlYHRO1OWMh7uHs
yh/ucVobDn0W7Vt16LQMoOAuCz1PbtSZilvsbb/a05EoLSLhOGHVtKAsTIpnENODK4XjZZY/hULk
sLo0+MRZUoK7rt69pO2rSJRE47DU05NA+lbWnGJJnCQZ3dAsbOp/Ij01bYcycp1Dc08zg4+2Grvb
Le3p2RniqQjJqUfDwO9xD9cbQo4dEwlRXTzXn8ttL0oRm1kxO57LZ2aIEAJ9qe0m053OpfMenTAy
QpMqJ+FL6BdfMYR8wsEQf9XBWmfzjkVR4SyyEWBSAptCCGG/Js6z2halOE0aTXGX5LaRFlnghzuW
fpRq5GPZts8dUhioyM12oR57ipOOFS5aY+TX/f4hJkFPat/Vai04mI8ADBgH0KtgS6l5fqgwtY4E
KvsJduLhrItlJ1NZE9Il+ezeEG9sbrF89cZAySyMjFUN0LBUAZ+Vtq7VfWyhjRiRA+7BBe+azTFx
b1zUjR8HEirXjVP069BP0p88qkzFCOSpWJ7Cml2cQJEs43h0W/dhJJa0jcDcz1sG8TFtkd+xqFFL
hX/fJnS6ozesUzwuVBFUMi3wPoGTHEJ/vJ6bUcB40TAHugAIFAz7wSnf5WKQHDO0hVNM9iChbveh
3NwT2QEq37dyEVJiXYZL0Jg9lMcD4rJWD3XoC645b1U6z84qDCerfYnSY1os6gIqEtpL8db30Hnu
QY7ckfPn3KUwHm7THD8sLv60bqpZNrHijUlyP31tEA9GxTWLkXli5aWIk7W8aPv+8O7HGxKlmWmn
t/i7cApm2vGZCi8TGb2NJPmDH6OZjCRYqjrqp2Bxoj1ggXkNg6rU6jRtkwowMKsRu2Tw+qTMP6xu
E33tZeB17N5uFl4+kIEtAf1xL1vym1LJOSDA7N5khHJL5hdEqDt7o5HZjzDDmGnOg3VNokN/3Xp7
U7vbup/LXbUjWOIsZmFXYHbuaNCsH9TftksTvxWf+eaFTJJZJWoSxOPrpOU0qBoKksTWe9ale9vX
nT9JM7y7sweAktWN3rSGKie91MjsS4To52lIsmmqksubBVheXiV5oXupplp3dioBHI6NpUIQ3RpC
W7ZWZzT6CdLaxJO58yFpsqq1DljUlXtNCHcnwUSgtErQlozkpwMcEnxBdYgni0f5mgnhnmTuflMj
uCsqzt3tt3+YFtEiobJfnMlWoW6/Gmb/D8ZEY0Lb5xxcUp7THi/29eNbnslh/mN5b9N8yQID6IJQ
f6Boek1TZxgzYeF21OaDwQ9i/TToFc76JlSy0GjBEB7O3rzGHg/WY03dbHuNbQ/cmg1HAYzetzky
HiPuNLwV5Z72j+BDU2oO8buu1tJijUa2bYv2eGM5HsHXHngQdexwCs+IEymvjTtrOk4oTp+7aAuY
QkX4FgRFm/3vcTqyN6uxOAWEDJ4hlZTjagggEmxWySD9xh82pSYAuI7lqSOaUfJOc6+JgBJh2pgW
e6IWNLRAaANq4686CzaKCGmwR1l1pUmSFTpr6D8BHJmjtiug4Kao2VE25xJF1A5FlX/yPbLLSJUh
FwmAu8VHrtv9EgHP6PWFuZjBGxbuL4kE8Bvcfo28yRwh9fRuorn98CfSNccwG6pLDH0rRcNg/92K
yQxPUgOaqhkuboyaP6/GD7P2t8ZBySXec0ME4emE3lAv32M6WQKOGLXSjE1iwR0gt/rcPkzD4yWe
EfhwJFvZzYwF//X5SSzLhhh01qXItF7PDZld0vGFrjefsTVfKrmQ8IECC8t8R0pH1GUiCCorrDix
3Hzokuo76/FybHyXKBKY/dRkUBY5CWw8Qc4TP12leTUVDCqdMN/QKJiJBZXt6wuwbke4SdPY6Jqu
Wr6kovWg3JvSIGu6aFsNY146x8rHZEthIPii3jV1qA+KOmA8+N1mjaxX/X+pqQ6FVjer2dN/G+Rj
qqUawxqEv5gpqPOnsNvf/ggJGo4xj0PC0z8wfwpdIfvFFVvOoQjjmDUPBLbTGmFvarveQBhOnB8+
nzqQhlTKwcQbOHRndPrIMEI+9wudDgX3HSIX82PG/4/Jjq/vgepOkhnrSj4rnrLWWv2GcQkNz9vH
9GJrrDV/hlezLPJMblWdH8wLXYENEWYh6z1igLVwrGW9fCSMOL2MpJLyDJCGTzIponGTDaja/TNe
QV1vSkT6SaVuChlbjCoCL6FoJ9G+qDcE1zpNdJrvNMxAeiteMy3URrb3wbOwI6iXMjBaoqZDjEou
crBm0MEKHUUxPLiNWVdfXNE2GpEvQ8Niot9+MEs7zT/1nJd/E41jBEp6scNcY4heqhauT+HuA4tR
yuDAmXYd11ksLYflAMiKd9tRPknRBLGyOrUojk6YCdUSU2/pKtN0SYVVwIpGI4MI0PytsCA45opw
Ag1gtjHlXPYbVVzq7N9qV7vPNOwBzP93xxaHx2vwyQXWv+PVI0NU7H5++q8zuJ0KQ+ROqw799EOA
G1kDFK3JxZdIbYN7p2diJempcOEe9a8pdyANgQ70XKt3iZI6Ndl0tv5EcAVv9PTx6AhJrouYvNBg
4ZQCDJqizc5vpbIKHPxoy2sO3JJLUr+BncbwrwzWZaRe5c9sDkfcm+JzQyriOgNExSPJ2Zo74WSf
P34xg5g7V1DVq9bTutAwp8ko5YCZZhFG3Ncl00U1sRenlyODJf70qP0vP+MXCtJxrA8mUr6z+Foh
jdNDnyDi9iJYGP5irtT+JzAo4wbAaLCRMcX/nHa4Z4dG+MoWdYgUssOCzquOotLlDx8f/mLeg+oH
F9HFAsUiW00bUy1GP4UEZ5mEccXlLrtYSuZIXTQA52q19uos7R2qEj8UXm7KcHmJNmu7e75Z0Ut6
YCKD/KDs8/C/QtQBe8JmK/4aEa+SIy+EI7aJ4DDqHjPFTsTmO8PU+e3If2cgqKs5q3aacpxPsoTo
OA/1di5DQ70QnzKDRKM/vQUAVtEpdYUSdogleKh2Omp+DDxJbLvzl2TvRNMM8spx3opRGbqCHtZP
pA6wF3N7m4RpAyYXuluMhRX9e00Ra/Nhh9AhMgGzZTv09OjssDAKBgaDkFGxDACx7GZgKYme6Hwb
QEFopKPzVIEV+8RLuR3WgqdecbP/AzKe0WiLcMal3Kba5knm6L2GSQtoWuf3YKQ7eHehCo1P2z6J
KtNz7bYEr7SFBZGKOK0SuGpZDgPVilGuzz95sF/9orHwsnhV/mJlUnN/F9XZ9izGLC0EIideTQ0s
9lwOVDqsIx16UcdmnyKgsuMlCNj0YoN/X/tH/WqjZGKmvjr50fTwtN8fRnWqSmfK43MdoXhZww4z
3RuM5efLnJvcbGqODBvM0Ssq0MTXhCcOR6YuQxtTVLiBTzL+KRjzWdY5ZEf2kL31ET0rVTxRi4PW
/mhGot2ClXT3WDIv5dhWkAkNKCCwvKRbv8AnJuWTGDeKGrXGqxfHo1NhHkXeInl9/EhlqG19e2q4
dVezbXLVpbhZD3MfjqshcpWc4JP4LhF5VJzXiAKe2sD6kElMEYbT0usY4eRRoAbu3jkbSOCzrWPQ
1Lcj7h/dWPJRD3zIC6Pe5QQ2HGmX19BIhVPt9J/dSzDvbilIsmbMxGpkYI7ZkmDnDfOQCZmh0Wqk
DC8xggqNLeLtOp5tWGNjmI5PSHdLKYJmM9kv8Ky/ndHn2bhzUjYaQ1IqhomRQuqQ9I0FvvrL0dMI
8NUkh+AUKGWXo+fz1MyMdavDjIwh1MYXddNCtWfob8YQfT0nI1k4SZ2ZednC87k1HazVET07GxEf
sVjMjT0HpekKSRIRefwcQzTM9riY+DGjbvU2M3C+0i+bHId5ghvyZ63NDCifqQuvPKcUJwC2n/lq
1PbxMwgjDcJbXw+PPH0tuP/8WOnWdGAz/9thPRhXUY+LJdnt6bEByoglCEd8hxz4PE4CrWsa4Iey
btoGth6+1mB/qhuHLZJXWyEurCZFV26TLwsuQJF3mx6NK0enKuPMJOzQSY+GwLjIM/ioL3hhADNK
4Zc4p3/IKbmRJBP3kTLCnIpOibcTcgRH5yVrYOAyXofTwdO3AEzR1q7eUdRBSTUenUPktvn0w4kb
WMDiXB9EiI0ODPgEiRRRafbmddVjSfyEG62vhY96tNtoFo2D9QZRnri5FiUktc3dxJeIQxy39WEl
BBTswFhCrPSBy7BInJAg4OsrHesPFQ6j0NpVsVnorOR6buVDmSw1gz9P8oN/mkG0/Q/tOnOyiUGC
HBtkzbAiGpswtNVaQIMiH+R+mia8j/FoQnqL/ekV8QqzvjyInQfclGg0gvjf9kbfqks5ws1KlGUY
2UZ5J0gnuoZ3mJzxwgC1bkRusiLUljdBDgPO8rE8en1+c6Pgb3H4RFlf3PSvAqgvcZOI/BWFys1w
ohmMqOTZtqQBNw1mgtrPvxX6kTZ7cKBqbVMBkRJNUm+1a/i3eYzyEBctub0Ol2e3JZcUF7pyTi1d
mXhONHU2d8Jp2AaE89vI6OWkIj29t0jAAa3nM+i/C0w/z/9V/3r/HZ/DQNKjgwUvpptH098SHAYu
D9RoHIVPSoGu7M4ugxYlsrG0KKUXAy78hoH/x42f5BfptazZn/PXRWgETa2njUVKybid5WkqpMl2
EQHAUy0QQCZwkfbahApSBc01+UAeKpe3HTzrtNe7N8f8I/xW+ruPlGQVaDemwhyp6M3fGZR6t0Bv
wG3ZEqMTNmBfTszMh/gRzL+roAnTsOrvs+ysYR4Yve0l5OFakbYltTD9L9iXjW72G+pH9ECX+qCH
Isi4m13lbeubz4ozVDgnjtrRpT8QanPmg7vo5Hh0w3l1CweY7cvQEpQ3lFqHbqlxv/cX29jYvCTo
9HBiIFR6FrvHIwpD3oaoWagos9PLiGhbVmPhWFRAiaD8OMsFqwPiGBSMll4fLZkVabn6BYMEgXi9
NhOz8Ju+b4MTbyuDXmWZDXdqD7nh5Olr7XqUc0G1r6w15d3D65uF+v2hwXkqWw90ES5J4zgrcEZl
2IQtSiCfpM8CLSnE8eL//4s6PJGuWMcnD0wC5Zxj8CCmQtoTLLrq/c2m4pAfiab3jcMMJN+pzzVp
Ue2p33cDP+A+e6r1QWBkQyyN0GYpIQ0R3P48lTfaDWkhicoz4UU2dgb3d6WA8cW7ScsbMDvZwe58
zlfPwMC3HIOXOpkoK03rrLQjqb+ci/q2/q1exePhUdcIXXCWNsneEagLkPs1mgsB2chRXY+2/yaj
ov1bbos0Nm9FLNjN9MaJB0SuFHzFWJOuFz3odhI2udLIdYNynyZ9eFdWlrDhCkd2YMubXfjb0q5M
mZrwbWENXx9stAkYdWIEN1zuMlGSxqw4uPzNDrBfG6oEmAobGT9M8dlyTbSOab2Xgd9HFBHe8vXF
G6ga5AxQMkamzmvIpl3vJeOl4wo6hS4T/Qzoqp9itkIaIDfp0+kp5Ixc8z0j+UsVX2UT2JEa3BMo
CwAltltfN0YRtppF8deaKTyOGIhX2llh3G0Y+HOx8BEvwrSIbCWVs9f0rhdqKWt9pAeQPOS9HsYG
wLvpmwEZQPlzoaJrNvYM2LD92hmoJoJYaywBMfA1Ms6wuuTmJ6cK88fOd5MS9fDlZkEpa6ryrmSl
W3FQPzlpFiiaN3z+9xCBf8M9TG1MToVybl2LHJM7VoloygLg4SNj0g1zoZn/GLnuF9z+b9GGPGlW
JIc/QrtJiQh+l1LrXsZWJladDbBIhTVBQS1USNxcLGGnUs8Dh3OJ6hSPE/cdrFZ93xxrAwL+UECJ
uKvjBP/UdpNa2TRgLPioikGeAewCd3EZiwGCodmdNPJtulrDSfOgoiUHBH58YVzxJEpfHCG5Z8oy
DqiKjhMEuwcah0oKtiMEHveRaJ6CsskpRi0++IGY5mfipaabHoU6QuhKJIYM+MisNH+yi0OtItGd
6oZOHuHXu94SBG9dNox1BGnrM7TU06MPE5fqDP5+7h13lxMMfFD23ZvX2naTckfIW9ZxvFXRE9lc
cZfPNDMUAy6sfUoqJxfl1fM7+/RJw8KyKHWaTUPusyYYL47EmoqbUhrHpEHAGBkPb1vbzTDZl97F
pUF7RUC2bMXVYC3Z6tvR5kzgQaro8BFUjiY8+McMG46RetnanO4hN/Q+TEdMgascNZJhLPNzhkmc
9GO2+9iunTxAOMYE5c/Y1Yhqu+x3K6nyNiQELrjLqTZ1qM4rS8C14alZt4g4TV5iB2q1p57sol37
0BIBpbUL12p5tgbV6y534Vt+TNSV9kf9sjtqltS4dFbJx1Sv3cs0Nv8H3amkYjdqWD65aoqcJ8sZ
xWWJcksqAEK2E6is7FYrIm20q30QlG/PMoICNCuH4Oqyoq6HVHYgFPSd76tkUQ5+MSg3Llms2HKn
LtML8gWbe9mvogLS91v4M7+Ai9T77bOM7ZPEw6dnLF/Q8+dWWKibCScVmiYwDYWMz28VyKhouJeK
AnKhfwPe1UT5xpqunspexdnHO3BUX7qKXz5J5bUqc5jIyKWeiXnBT/c9lajStLyOwBXIsg/fZFX3
HPfbgs4pl1Faq6vjDxlWjTJrFHlzp9ROMGgItA3qPGaakSlSGMbGLnTfMamYOy2yKowMlDT36PmN
xj+uj58MXOU/auBxzQKGz2Tb7/urGWiStTOVPJ4+Fl965LeSLCd8vcf6mIYlBq2y/aKoeoITCnb+
CFEzRmY4Ayx8FLvDch9cA8Rx5OEqpEyTTUfZ1TZeUyMTxZuKC6nJ2bUnlVGV7kpY7On0hC28VSO4
DzWbDur1sucsGqCVWdUxte8t18xTUu85gV7fvmiFPj7pK+IJeLhy8TDbdLLkqItS1Mpj/Te+z6oz
pDLd1N8SocJsJj11CyOt8S49WWHZ3SULDZtHOWxIV9eWoLAOSBCKNJbBarGq9ag+SjOO+zpGmVvY
tzeSI1Q9dGhSr6tFsDyoxrr9VnndxAEKipBoxcPvjAvd/IL0pS5A6RAvwlL/lXm2DUbmMlSL9uRB
CtMhZr9Edt+rTZJNE4uCCRqiQ1A+XdnpTHdvSvUHYeSX6CbyzLKZahJAhE/07jZXWtzGJyq52zm4
PyOKDYRYsgTcY9CBtXh5+0Wv7u4vcEkjoiTrC+Di/B12bzGZcx+PZYVPJA/lMy8wPCYz6aaZno7W
6QzgSqhF+m+iQUaoEuIUHRMMFScQaX9fhVB4MsFsWfTVRuNgwJeYD/CUJK0ecxk+LlcCAnNpEClD
lohDWWDnrdrBYrcwrQSa44suJ7UOcqdVU6apfJTABJq0yH+ev8xCAGMQEyVi5fTJybAPj+oC0xAd
K7AuFhi6h8UI0SAMCjJwGLn9Al1i2xv/LYH7UWl33SuN4GaHVxXAtfNFUxP/EfCkiMeUCtv2Jds8
tGL2b9EQwW1P46Ex5rHPttilC8dHYLYtTamKeKVau1UyBXtv3xoZvgAGbhOZTocj4yJElZqJgtB4
0HUMKIdCuhF+iB52NOY4DAF8j2w/LEBVHzZTKQb7R3rb5IUknikx5OnIXPimYazSDbpcoLvLcpg2
2GMixdxV5xDp+zFv1LG0UY/oZmm1NQqacDFjAlZF+xnW87tqZI26HqSR7/uGm5aCzlRrz51rZlXu
Vzt9u24/jRtL8wYhT0qRnA3WQmotxDrajWWQLB4t1BGlR5Y9PprFSYMaifKMXmdppNUigOjSP6ib
ZqpU97t6xqoVva+D+At7/ASP9B4JyB+vGAxI/2ygjEMHXkEhNtqwDnwboCZL5P7g9i6D/lrDQD5o
XtMt4tU2UyJCGFLlgvDUc09z+V4Yt8ZKK876tR5qZMc+6Qpj5R8uTTXuL9en6DsL/RM5K8M5Od50
ju8RHy+lxOpTwJ1C9YL2Fq0mkHslbqV+opVueNkd4ordxcK0N3eQqOADHEMnUCLwdGSPnQjZcKJD
UuS678KW4m1muhzPUzCCdeDAlW/OhvLlBwa5yzLS9NhDtmAIXeIQ+klHEgB+QR0MzgtRzOgQp5vU
Sp2G4TgvV0bAASdCihO2bvmgHvZ9Ttvufr6jVUpLxoyH4GBflafywQ/DgDpPe57Vi3wfMPw+AIpl
qXrQxMdldIeQwfWa036+bwGzPywR1eORQbowKXsK4gLjaY4JGee5PvmYWnUL9y3nWsi2eV7joCAm
OiLuCAWrh0Qwf1AgY9gFiR7+XrBEWZ6bi9aPp1/4cpjeDYSyPYwXBeK3KYjnsSR38tTZ48EZDMXW
VWDPoX3XlTZArVl/dLq3zDN9Th9pLbaRryTMNanWy2JQIRrDY0kqld3e/d6PjPe7BPi+wQafOW89
7h0tq+eoDIvDtlmpHHffFM7gOzhQDIyxIfFRozQN+SGsSdAJhKGkldKsnE/FUpS96muXr1KAAIpj
1nROa0d5qe/PS2tI09HyBPmga8aRdvVOocP8BuQz6eDcm/58gpoBWaGK4l1E9vB+6S7R5nF4AvrH
P2fvxkb8nky+iqIjvcZbGj1DBhX7y3FU4YmOGU6yl+XSiCKMl+BZz8pVSSarq6E6jSlz+gXjVM27
tMpriKqV5/qPDqAk+soYq1JhaoOdZxZKQSKitFJge7lx6SnpiDRpQC8oQlsXUJls2alMghQIDflZ
GBTPzKOE+7zV2l7lqUVAPZzVgurVmGQerOC0gra3RNIj2R6FMUGieZFJ5RKgZTiw38MY34Ogx5He
da866nqoHaeitdYmfTpm4Icyhac8he8YyE20Wz8x/EAJwy0jm97xi+toPPmjIR8wObJMSfAYPYYR
ztByG7hNoNtWVqcjB0FDTuE0kJAalNlk5L5Ne3P95xszPBsYfOQyNosfwu4W1BGSyxwMPi0jQneO
zDf+IG238NKwSzR0+8DqejQtOhb7qN2Iy43vYY78elTRXAhGxf5qFLnoORE8dBiSJ1mIQ8g0D/R2
jioIAfmfbeanBduXNrDpcpm6gg9ASScOoFvcEA27bt3Ug4gm4OgLA1MLirL0IuMTBxDsFCrRLQcq
KffrHo76CqMb6UnQ1MIEFO3scVAERBHxzd5R1c4qXVwmQILWGrxdqPhoXH3pCl888y7Ej3ZMoP8j
E0v//zk4RKGhKZAztaUPMKXiJdVOI4gB/tdTS3ml4x2vtKug9VdoOrnwFY2XiPuFEJgm/9Jn3T4Z
HsHi0oZu0o1TmSkIkPDFkxyOtQGrodBc5ARoSV4qgv6UGTVh59FXrL6idTgOvy0pMzpVzlPh3kH6
l3+b0cZBkcRve8LXA19NRVO+B54aQFMhXUsERRLLTwf5d8Ht/HGMESW7vz7Ufugwi6z8GkcpfWc9
3B51Db6bjvH5BD9iVW8nVJ39QWlmMkLN/tiW2dO+NNxAmLfnBTlXp3/8UFnTNchZnlE+ifl3hfaq
f/aqYFLpHZDrU4ahtF/Vto+E0Rj3Y2uN1ALKq1GBZc94PWjhMIvgHsu/mKJAbyqhooWwTa+luM+U
1je/jix6EWpbyii/WiGBY0RTW1Jj2QI8piJ4PBk9J0HW6jpTu2KUQoIQPcd7CoP4dydySn4eCMf3
KLtB7jkKvnLbzZJbJbVIvbZ3JEJ7Z2mNFCNguY3TjWHgqD6KQTZyNO4Cy8QynjLbyC2fG7ccMd77
7ChG43VajtYyXITdEXVvMMUhuAm0lr4TJTDpH5js1qsdCE4sI82WLPZFjCLfqZ0cCpYK8dNP0Old
y75qnK5CQ6oj6DnLWVZBjk5jxupQzXJnI4yTzdrUFqq/lDcDB/SMVvypuk0giXcPsWx2LmcOVHu/
6ljkdqV78Qxdqi4+tmzEWsG2rT255EOIA2kxxN/FiTmVj5nhVhmRY07DUoCXtSQlcWoxZ9ZyjfLy
WhNvFs7M2CFzcpU1uNQqoXlIMpP03wtfGwdiHX1qXOzP/sAYagy1EEqSlLB8lDBJkiXbpa3QS1wy
PIhSVNaVcv0P6VU1ls1mnXP9kVDBzO3CeqZDwXJEGOFqp1ljJILQNR/WRId+G7UJFoZe1//XGPVP
pJju44Sv1MEJslMx5FuaHjJLA/0ofrPy5LF8EIWAkktJ6b7TDYLDoRyycPYCr7i9oz62DeACjxF9
89ZSiWgqAQsbP53Mqx3egEsiOW8E8WLS5m2TnsOumAEZ5lKbQg1+3dhxxZBC3AhYNlojgkSCK8V1
KKH+iomKaiJ5t/d20waTFShEk7a+FJ3fRWwjrn6I2kKcRZfC/brvr/nEje5zVWJGJV2JHVZGq8ci
ouRbaFLoyiiGKfMONKxWXgvTeJ3lGI3+MXik5exztipLXS2r4VtEC7l0fPXTsH9/NwCK+wn9V+nq
fLjpjlfElbF8UbEHsC+K2eWeDvViZTgPWxd8jOJBhkUnyD9NYVku32aVKSBsDxr2TxR3ScvFiBRY
4uT+DN4sz6PJwle/Xy9gD/eQXmK+sW2ywu1iV3lqm1c1XhohoaEOXSMerhQCa+r0biGEeBA9eNPC
7UaYsR//1sUQWa/wWYNtcFNh6iYOwvJJogvey4dlKdHJu67gHGXXCFOXTKZ+IDuqRSvHmXmHPIB4
w2FlIVr6ryP8MSLSIPOkHZamL6l8RQoilDz8dqodGGMg7J2Y2Xmyqzg9GHj0hYWOSEY+YvA2G41x
P+lTgKcu4DDMKYBhq/V7meQu0rBrosTqefPb9troxvsnKKFFhBpwFNFG74VBCr4pcbXKTPm32rHU
Y1mvMAvFfAzisynck6Tt3zPWc1i9wo0cvNGyrP6cFHYcajEO4Vu9Y4mxyO7O0rCTs8pitDDeJtSB
Vaz3bz1aiIzH3v6/I2B+o02zzDJe/5rNTmcRySApAUuOcR7P5tyR9oeVIZR5d/hWUVjOfDO9o6Yv
8d0HA7sdSc/o/nkWK1mVVdXQf1UbJriokTvUkQxh/ofDq5cwnuEyTQUDCHvvpUNrZkViz6BA3Jm4
zr/p1v9CdzSC5iIdlMBScuoQm+E3D0EnW3/DUsggGjBLZ8GgLbV7MPV5WkNrMFH6mtVN7KnoWxrW
Deg0lfVQdZSq/u2Uob3zww9qd9+auDKn96+PAHh5S4iiCu2dPEH2rWxJ1jNqBJKREP4pbvFhiEJc
Bt4GV8k76NM/1fmAzk6SzeLqZT63w9a+7IUw/OMQvop8YF3w1y5EuVOgI6msizDGQCM3V0AonW3g
SpzzTD5o3PjaZs7cPHngDT4PpMF4g15JXPz5tM4465ghicdWpYyNFgxeRxiNJtqn3rk3nkVog25u
84K/SFYTDife7ccbi73GEiaqZwB482z4xMFJRdmZIkebYd2qC+mNSrwLJbqKE4eaPmCp8YhT/Z6A
rZpHtJUuQb21Cp9thFDivx/gVwybESTjtYBYidAaHc8AAgu98caR9+9gKUEGlMDA2ebo4w1hxE9S
V1ETSs9wjkwj/F5nPAp+W/KxGCQ32kLqDwbJGS5pkouRKCvkIEJTw78Dky4RVl81o2w3o3TEeUXN
h49mfVNhigJstJY9+a2odLY6ToykNhXMwCGVmSAWMsy9phlLcbhR01SW/uHvHKg4+vnRmRWp3Kb1
YgRIAWdbevIpUArdmQzhUzLTLYFNXRUgp2YPYlQwP0SBdDY7zFXehYYq9xSC+JJxVYgP3Mh4ufbT
usJ0ezDP9WOnEQW6YLsRpqy7F/2GwseWLgqW2ntiOZuBppszk8out0fZcZJmY9DEsH6ZPF8HJK0R
2Z6lkdEmDuPGvzS5ekD8OGs3RNS7YpqKj+j5fP4XYv7xo+nd3boUFkFx+t3kUcjgpWdjicPN3afo
bO80GSPg/ACnImYl6I2rkrFbjQhrO/HBz1OiKrjOqeYaUa357xCbNHdVzXiC7QJfgGJiy4Pnculp
j7A6GxoX7qZDLgSPiVjPI5p6RCXdr+Ez1LS3kItRprMaLTSNT3dSl8H0Wy2VmcJo6ed2qW6gj2dy
qs4O9I1BZvmTtHyJiIMvD4paVRgZoIsDIqhkZi3ZD5G6AZptrCyjGYjYl/FRnWC45dKAnNL5n7AH
y4+ZpzlLLnnI3rW2l75l4t7lNVG7cazrrEhYh8CGpaJSj3xGdapcyyiqkRcleIDiKJo8YAVraO77
1vGBXf5QLJ4WZjzPCuVtNKjwoNuKheeqDbrvTbeddHUJK/Yl6wvY3w5wclrlNf2aFUbTLHJS1cw2
+eRkkvdWWXZTiGEbwyZPYMaTPn533PaCvpFUoEn45HXsFYX71J1etoWBElZB9Sgh2c5bqOPw1W6V
FJOFJfagPuvtYD/PH7lbQ4HnmKqCbu18dLRql9NuqQttmrn6lytDY3+LC57lOn34L8ruv90SL8t2
wf+JLi63u7cWrP/kLgj06xWlaaY4UGRPaNnBmg6O6V8tXh5v1bBIuMH0EP/WdPi6Mdy4NnUukp6v
BOl1CcVV7WYMKLpl2HMkC0Y6oxFBgmrxld2++om+NeGx/lbmB/iLbXMnLODIV0rGU2Wmh0LkjyEF
6B2z8dEo1ze3un3QhpXMud6hgwRwis+7qgeXTExjkGKBo7brVmDxKChiF1rLFTx/8tm77MLoldxv
vrB1HhiXHDr7VRIoIgatP53jdXVSNPZAkDYifhacwRxpC78Ho13a/bnw6RM+b+qdeApVhdCrum6y
mQ64vZ4tg6KhAHhpLUXnQ3wmCp5upcQfVw70mdVR5eCAbKhtBXnMjYbymGtnVHEU976FJMPSRj4H
zmmrGPnNIiC6YY4sRc5qqh5O5eg5yfmBI8q0dOWdqgRuHqyvohGTZmrK4xEi5HvHc/fehJthg5Jm
QbTW27WChOKbPYIJrWg5/OG9k0w7bjxGj9g0ygOU1lwiVJrL6Utt1NSV98A7HrDs9Y+2+DGPjOwF
Zemi7yOSJVQ7kSEgyF5d8F4op2k5671CUDAvRtKfqvrFtYDqbPYi7iPWGP4qBBFOggOgYJWRkePC
41G07IY5JCIw3L0W5mVrLL+Ce5eAJ9sEd+C5V9dVjyJ7x0eXzWpLQPFseOxat5bbVNFjQJU1VWsm
Dfd85aSWT4E/E/P3gCdWkoZyyNiLlWsGLaXKiTpSUTKbg5wWVfUnnsb63qdHlK7d1T+DxbPeb3M5
yInAlnX4+BIbDRLTUyFt3+Uedbq01A0f79wjIbiaN2sAxuRYOVZ75e5hF4z8ymaNeDk9n/k5TdTA
1R0QUuoPL65pc3M5yL/l+2PKd+zNgegl4FF9AjUstxk4phoI/s491LWj5BbzshvZdVZ4kr6qI1yq
vqTZLWShlSJGlAdzA59xVigp8W/1trJrbEiLNgphScwTEt3vD2P+prt7+lWIQEAvM8Ee5X1fVQ0N
UA+NYqCf7Gsf8HIbX7D/RYl6yZsmAkVa/nvMyI/PodQbXlHw2CNJrdUOS5/MJD/a6uvxzOmqc6L8
+yUUcsJTp0aPwkhfMpqWrY4/xNFKl2ucaWu3ra37LLzATgUUrV6f47Ab/qXxVaXsHE8yVUxSDTT+
Df01oLWNXmtJ5uDN1IGsfSk4Hd0OYfHOI+j4ocb9S1B430BTtnCPgamW8YTCvgCQEvV9zfh5lbYK
SEqiwW9nQQzu8cgj+mYlS5tLEFxjDpqqfBqu739bPN6QJCcKnrqKDQZDVUdO8JDiYLQIweKlHvEF
vCs7EiTj9JZnJEi7A23/WcBtWjb0L0IDBiteZxbZTyioff4LX20inP6a5OpzoQiI/us6u6OXv+Jc
jB2qHnk9Hep8NcqthPz48HyMMuWo58sRsUU6uPzFIFW/aMpuoqpNjVBldUo0zzkNGtroUORPjRqW
IyS6JHImSkJ94+OvERqLXaPu3ENE0zE9xTdJH7/8IEF/dD98OnyI+3qAovVCJ1h5fIRcQ5EIMvB3
tVn4fuMecIyLqrDb/fFuY+3eDhDz87SVjMEUJuSxBsa2pjxaxxCrQSkkzWoxsEFWjXl1FZ5GCvA1
6VkVyJbzr3HHCMxUJGoRFKBFBPOlw0EZWsBS62QgfDlZKxqo9gOPp+SUf0Nn9aynmODUaC1BoI+l
SihJl8E5KM1jUa0LufqDvnzgRB1RNcMwFU7IqQ5EtroymA3u2GbZaCeFHlHhpIsm9xxKKeYuFgAn
U0Vdg9uY4QkH5+YOuFeqhTVWw9LppKzgSOmJJpBWDy3Fz4ngYwx5+lf3fpA6VslXpkCCSeH3kJrY
GgLFcvW1lu845PcP+RA27kCxy4Hz1A1W+39rf0vfdPZsaGXVrgdffKkz6s4krTBmCEiWMfGvf1l3
v61AHtSpdoNA+B4A5iC0qba2R6LKFRQ9nlFyDn8gdksNBi0mJJegej/Z8GSumTSm2Lx0r3Ae3mtk
RV7/+YOFvRzEsA6ry/cLDZfuUgWQBiuPWP/dxMnNC9VZ/Ri52VAPpj3W++3b/QCmbCbC7GQveewW
drkwh5WrwSvFJzE6HAKytydeCwkqU38z51GlYfv5ExPaLfe8JnsV3GWSeaIioG6uny3Hc5RQORoV
3T3a8m/DG3N2PPYZ1tOq6hIG45USzirnNFFCupBkcUIDJx2zDTRyLx0IZRajerJXKW8vDAx+XXrR
a5EAgzdIKQ7sdQr3s8uCfYrywVAAo/K/CfQWPcMHHOZ4fO22uVCpgkaa1qnUAPllsD0/RvTYGgKL
7rNNd8t+ul5Eep8VaxkWj1blvhAgo6Q+dWShvlJbt/Y1+E+9woz4heirDk6LZ0S24ku4N0UvMSet
La0PYeMzJOx1lIcJfLavSH5eTpMejqTJbUTl2f7OfAhf0QJ6+0u1xt5eb7WFf44SVKP2OD2nl63u
fL6+XLTNj3iVdgS2HKBOzydsYefkjfp/Ud96H3LL1ERG3W7q1ytvBV8jfGU8K2uaP03bHZ46ztSB
WVKsGn/eoshtwdAPfDhl+c6Ej1ojqQZhO2opXPniqLW9Uc2ievTdpA7aS+IVsRxAdfYWZzM0ekDy
c9sygpM8lzmkvgSEOiNaOqjrNcMJqFuzS+Z4psBfuu3+WWIjcvU8XghzMyHKMqy5NJVSJrbfI5ID
Ftduua/LBr8gOz1e6uQDs6KNXGrz0I+cNEo6eBhwKocW1I9nVRrJ8HorETbJTtowiyDC7PUOYVK5
YRoQUD+krwpNxJQOfQRoyVGefQodcrD5QpEs40ARcufatb0g/M5ZnO8wjNewmboySz+kRa7PW/0/
nnANrAn90kN6E3ra/hF1YwXrR4Iz68s7g0fQecxb8rIrc+VfgylMOtITYP9+CcSTJaFkltRFynhM
6PcZp/u8D7u1Qi+kJW0jPiwHUaE0AKKZ7CIIS+O7+NG4iLD+FkRyk+s0k98HfH7eNsw7uuXkgiD3
+U5wH40GcyOLC/RGhnZXxugdz3+uO9EA0TQ0hGMGcXzykklcF6Z0xxg0ITkcmzCw/3se82yzmGZn
MAhYDbdAqQz5t4tTcUgQrw/lP/KfUtsfa5B5AnvMa8KGz4szOddUrmPpNswtgDuqyuUdFJ9V7dnb
K4iQNoj0lyhSquSjWbZFa51XUeG4nebynvWkU5p/AoQZq9CbwfTfHQ/dE9XXVti5UDqwwWa13028
C+HISjl3p7WjjlHOn6GASjgtPQSGGFJmRkM/v5iLrRz3qGQb4CsFcyf8guLUjk25DfIHNs8+cqLX
LV4lHy4Q59a51ftNTZup+K0CgF42GW6gOYjN6DLuNgQMUYLde/5K24aCeCRGUD+xwRo5sU6KTGeS
dLf8V+dkN0oYFP1rZlo/wiJzl51aovOQ0Y3Sjf1FBx5Cezc4RRhDKXxIF12hA/Da1khGhA9YwUco
ZE4U7vXotibSy9tMVvuvnO1g+TEEJzzUK0ywXLYTwDJG/9dsXFH+ckX/dxfRLHjshBlXbA2R+ahs
2ifQRmAbTUBeE9qXVD9GgPkACNMH/el2oXu6Pp5jI+iL3uMA/epVi98xd8N/rMJiNyXSho5rBBkL
E2nit72KSCkEdXW6mH43LggovmsOO3Cmh7c/VLoGJrz4JGTC0dtbCrvUZ5efiQXyv90Li/06xYsA
Atfef/L6TcY8OId+CWt3abx4HkX9Mh7U9VobkR4kdX0eTXVZFnPhj9cP8wSrDBbwuG5+IM412Uo7
sY6Q2Cu26JfCcLEZJXZK8FFPXIhGtnhXEEC30YcFVOxdDZE8eiTAoYbDP69aluZrQjrF3HinWmNw
2hbNcZD5scpXopXpCeTMI5dY6+mBKh3mqMZTbiFHqiXh1rYyLhpsxlzapw3B3Xl1GCx2En2r0N3t
Wo8UasBy/Ljh/Be6yOAuI4tQ1iVZLlHG2ObNT8w8/rFN2KPFgCFCh4NeT6yQYfb9Rs9tLhdFV3+o
rWiXggJq8RBEQwTueLh4D1v7+PMRJzJUmrGWdXnEOmvYG/DYEXWFDd33KhQE+g8wgiTi4gifD73z
5e8WAuRJ/c71kVesN/V7j8VBjkJHZKUZBFOHkcYWU0AlN2HZ5PDSYMtrgKbgLDz0FnR/v96eCQz5
ZYWENs7TjBuPPvhP0bslUZAvstau3dqDBxMq2BsSw66GG4z1qnEKN6o1pcPO6RhmDHX3vbpuhqqU
0f/VNgUFOrB7fDHOwJAZK1uMFYzHAmYUI4o9raWoeLwhY3xmDrLVvhpqEOD3Gs7RTKVzC/va5A83
cUtRSxqaLxhPoRKe31pKuAyHKTbE84PlF/NzFt6Vf+5gKoawCz+qPAnBYtJOx686I0X/k7EjIbtT
+pyTQJCJ0T8LZ1p9mcoHIuTJERJwTjy8eVJGYHcPLLcu/3SY2AUbsi7sq3XBPUWtqGdI/p4JHvZd
+M6EPS1tf/6MqwXiJDtKWtzcLFX6K9Ug1QHlWbpEZYz2rcehwwQ7yn9/ODuByArYi6983JMQQv4M
NkQL7rqcdiZ3OOcMZrhz6rT5gxS0l9J0IOxmD0qiL8eCynNnfkF9dNvuUJA/qvhg4IraJ/4Xkzlr
4AeIZZC0/0svwLWIPqpHJ0ZBV/1wbA1tdFHA8xxgRmJOCSLzlWLRI9dSZFHAL0PI2ef3sqhG9v9A
uIGK2hxl64/rB7rs0CAES8lLufcNAnnvC12U2P84M8/EsYlUyFsDbjUiStJNckB0NuG5c9Sl8t23
tUiEZpaJh207mvJSAlCT7Rquw3x6duzBU1B/x3ReqflmEPviMDlCZ0J82d0v+itdMUfnVtn+5PUs
s1xIEI4EYFUTXmPoVwyv/a7ZqvyaU1J8MkCGl0eysM2XNuRz4osRVQ7YRi56hJAKM8vPfPslHWLS
6grbRubavamlIPYlYtaUwtlyWGb0cWYFb5dn8PBaJUt+wdeOePaX7gQrQjCXCeFV+Qt9OLNm0gwe
gEA9d/bJW12YUf4JwjGArPJeBEYBnqFjxmJwUOw9OuHkcZzrKkFlFu/fBTI06BUfbxO0bfiBUO+D
P1XPaKfbwdsIQSO+Jx/FpwvNyE/YfbhVClNjA9Pg5I5oy4iU//i7KKpd7go0QKNF/cGXOPdYbg5I
IMWxY1Jsg8jHNOVHuXsv7AivMeZDb9cwY8kIfLwqmKGsdOO4BcbOAT1fQuw0IRxmxsXnKi1VnCOs
o3eQq7A6eckLs365I6ZkG6qKEwLrbQpHEf0sFz997jzh4tnGDXhZQqG6xJPBgd0qbsJXGs80k4PJ
x0ZZZV+A5ch/cXbvv0aF1t6TKBTKz1QU7MQt+GSqIF8E9/5lbYR798v8TIR6NIy9cm0Qc8nEdVBL
MWkmOm7JUkr2F9Qhw3hTyV7n9unOfs8TkeZZwEHQPYQO6yaTjwfbOfLHDKqSR1dj+Df6clp0x8T8
rcF3EX2ssBB09gqVgA2IKt5/Gyq1BhPlxK3bIGmp5+5+v7WrkhegvDhWvQHsZ8QyA9ldD9ZOToXN
ilDtDUrqXK+HHwoynRCRx1zsVK1MwMSguJaIM3zW3bK8jTQLlkR/0cDAYb15Qkr4hsv6Mfc6R2hM
IAGT2iLMHGFbmebm5Ujro/UEJPfHqgEAfvVAbdb9yuphAjV+Q87JthlHpwdQqC5QoqL5HvUdiLdb
DWi9tLxDHC4Wh82+6ywaDcyMuTLZI0hmC1nlTIMICufUD5/3U+hYwOAGzCcpP8q7Ne2TyfBGrcwt
8c+saoyUcRCCVbceArQ9JW52IeKiM/Y/xWHDgdLoAAxLAXtODPKckK+DRXbQwMH2yJaY6rJA2fql
VYJ8ABARQ5O/C8Nsjpb2Iu2rQLqi9Yrf5suKcENTMHlf95sqbMzN1MFwohpeoX84HEsJmxvPew7P
PU2nREmtvRxj8ITq1eQBtxMTcxftNR+4/llANxK7GYxahRqDmmxA8d/RWibpIKFzkshNgG+Qg4LB
ds0DIXjZUWl7c4+txuNPDDzLX7C+7gUyIG4YLNfpnL2YAnWEmsOsH4IxJfauI/v86OF+ajkrJmio
c/BKVeT1CITp4ZKqOOJxwIYStKRxHfw85YfWQFKU3ksvlx5KX3T1fLwgJ+q5WQub7HXTRPBQnfH+
UPdTrBlgBhPO4YBSBicg2rJq2vkF0oJJEm7dIn8zGwU+1cWU8X2q69Q5Im5OFq1TScrXBbuYWtAK
ot7nWpNwCWmOY3cdqHHrEeh07cunq7EEXS4/WEbbNyKsjAXj0MGqqVmu0CByHEKM8ID2VwWOHMsM
SBCPIMrKFMdh3pokBPS5pAhRvnBRZTxpvFCcsC4UUoHpBj43LgpFlEgmZl5WvsJpjyQuBl7D47UC
w4fT1Lpms90zeB9mDW+eRKIC6h9BuIAQBUzJYVA15cfc0PIuA7B6YUTZJsIYGO/y2QYcTAv5VzHK
tgqNq6ST5d/nIgkq+AZgs2kEJGL1jrPzKWLlrUuDfDZS/2icwOYwHIomieEn9Io582lfwrIQo2SN
iRH0DGxIOFHkKJkYV0cgHluCrSGlWtXTSILQ0sSiSJY015HWnl6tW5Aq7Cwken5rZny7VkKNgEiv
vhSeONRKbQ5dk53GHPs5puaBiNOvfl81PTLXtfnXcUlB1GsUOlw2HnIYUT/eMVA7Y4xwE1DihAKm
km9LNrTcQt+Q36XI09opSUevXJnqqQTCip2gWEGPOWKLGTA49NZMeD8HX7MBkt235BmnBxRrWpW2
70JiJF61vUnaVV1AUz4Mi2vKpISc74C6eMk+/1t94IctDkr33EKjnBxEUidXRtI8WGcBRIKVjtYF
wUTgC8sfii3LXvk8p8CrfiCScdaBa08TuniLuFp08KDKYzloVj0qToGqKy9gNPGsoJeF+vZaZvn1
oweIziDJI9JHhl2Z/moDJfHsHR8JqdSRQnlArYxPutm+GIui5oSb02wpJ60gh2sioQ7HsfXfFXmA
vp01VCXH0mxmmYvc3wCqp/qJTY3LYnyptmzT3ld4ow7ssa2oXJ1zlc0zzjQpR3ySx0U8tmrMIm5N
sbwbhj5B6/pC0WQo2K7qjZCc21yg20XrgtTOd9hDptpbZBj1r2Sf7UkVE0o9Ue5OdUW6h4jnnJiz
1CxlbyTsQrkXT+pLyCxDEYgg994IC+fTdXvKyPPCF6GKWtpgQlc9boxMXEBuIjsnb+HmfVzyBQHd
rXQJw4YKcWM4OATrh/aMCxsidemv/QHQ+gPpuuQ5zJ5Y25C1CE/pwFmznIFzybf/efjgU5fWE0r+
/fmHbfJ8CGSUo7gYQCSBM6yabHdMXY8fvPwgAKkKuIN8V/BI1PFmCX7BgbgXhyVhsMmEZxsFKSyw
2c9MW/X60mDOBqDvRPoMsN5n8K3n7qtDP8dACjwG1vXUho9EGx5ohm26rZnC06T8WVypOb0vW/PE
dlQJxLSHTvmMLeh2+tqrhCmewibEuZeJ98xhuaepVLFs8hbdudIUs1QyX0muncPD8RIeudbWDmum
0tHzFKfZs4sShcmhiomukVhAy/E0pKeoEjhOWO0ZRo129hrNWu6tyyu4vV8BFYiOc/VMKUI0zZw8
joegGErbe9pb7jwIGmcJL/xjqXiSGPOVm6pz4sIP+vS7EuRh94QTueWe9HAkH9aUuZOEEcofVKip
qfIElwoR7gmUdHntwXoSfc0MTNMASjhKGzCvzNjdueXFjRXNhNNxTkQiiAVjVjKDQ/l3zCHksKbm
DaAGAnQ4gkX30vO92YOVv7Koef/8wBYBk/CwY2hYezY2dsy6XXLaknaa6cz30pMuUCGoxmeDHvkt
C3Fjw9i+vmwoVZ4ob8UhxJ5PFc1dpIxQPbWw9Cu9ux2Hs0ht2kl/31QRPAUDuqSK2BhdxpPlZyEE
JGfrBIRhl6phBhNkAzFSFr+/p2bFi4AUE/W/SjW/83dBHy6GB/W+53zsdCmFvVJPZgxOR4ZKB8Pn
2S53BWAwBBpmUaQzxtFpiNJE19uj7zWz+orjrKqZniVf2JmZ+Ys1eFFJTuCoQIoHTlbX8reCrgxp
kFd9ZWRuLO+PQkSjmKv6XNHjwpyszt7muPXo9eP/uk47gN7rs9LCJcbJc/0ewyIbZuEMpkMgoWrk
TJM8zhEMpBQ+J4UpnMHp9WsZDjzUjA4LxXF5kUXkDxNMzrNclKuZCKQBWf00cdG7gCc1oIOGRWMp
SVxvc+ZZeLPJOLO0FkLqqje9566s9K5OnXw3sZv+zfGarqf25gq2kntUmhJRCtlK3kEYh2VwhPEe
Pvpj5jWI2c2oiZiWCpX+iVK5wg4p6brc6RpARUGSOPnAsfAidUbs13IE2mqAflmftnwmVyrDCtim
yBIG5UsYYNJ5ZB61h7DQ+blR1racuOZ7xypwX9EwBUXcveX/0gweZ2VsAVLhKFEyL/9nN+i22xMs
oamoTdlHggO8lWV+rsxKJvky28w0Vm5ss1jDkW+VHPpx6kAVkTjql37atqXYHS+0EUvNHMkvAHIj
ZRR3mY433dMqZUepCE87oeogcFCAn3UBAca4FbtYPaaB70je43dylnjqUTz8Z7ZLJMlMMtgXctJx
hflL+tH8Sc6A2Fd4Y4NE65TA8VY/bjugeGWxOuV+w4gSihWXM6l8qr86YNV+JWTU3RXh90BqBwhR
RMm89R47ke8eqtbXxwDredrbmXvuwkE1wSKla9/vggfIPOFrPjZGY/jvfhqWu8jKrKBzU0JNRT9H
p83K/GS3eDCavn5rwEG0eGG+WwZz6c0V1027r8ezROfJCJla/FosOsR0tZppAu50CJlzFIMqA0NW
J6tpQc7cvjk3Fb20NNa91lSrS8yN0ccnPAjW1aHIOudUizxi9ZS8FlLaqSce8s1hoMAipdkHdBne
mnvVOzPsojIsQBzEGHd3XhKfutKuJ4NntSV1q0oAd/iLIKa7SqzJ2Zv7s5Usbq59sZx5DjQTi3pq
wtAAOGU3qfuOSGz13ssKvuatP2bai6as/3wjIYHXscfN8/dHPscpjYUuKzqZYmvfveM5WY7Cau0o
Eqi2QYBm0hHnpsCSQqOoGeXjRxHsR8Kid1zMLcqCEpptCY+eP4g+fXqhjIvT4+t8L3uuXvxkkb0H
UXzTm9tWswm2IKeIJHgZfJk3jN/I/iWnsHZ7l1fD0IGpXmJ3Snuvm4OwsGa9X0TyvPgrkdXDjbVg
qErj15vXBh4lnGF81fYIdqhGSqYJxhTQrlkLFUvD7u4UoJ0D3/BSuRfqI/hW7VVdk7tCfa8WyAmo
1fxv6FKs4jLwKQ8n4LPgoQ8GXeIxdO3CKV0hPql72J+UPG5SYoEF2f65O/HqWP//TmyFLWu30U0P
y83Zq43MOw/gf4564YxV9HCSyVPl9/92rjHUTypuOQzk1VEPNiRO/2fFEtNhIDIrTvVhtZiceHXc
kmjWJL2QDtwpHEZiVRYcnDZwKPRHoVmsjICcXH5kAvAlOjJbOf16o09wDGMLHRcczohATG8VtWUh
/663aGUWJCvGuOA1saCAJud2cb09N+KTu01lXn/wIqjamXb6tfbYrfn4hfglUr7VbCoHrYC/+eR2
XcL7NNFr8gOc3B5Gn7VeBjOYy2W9zib1ugW0wSNPDUfb0eL4bkILZ9yGcCvv7CTpFOmHX8Fy5C3D
bNZr/oY++quiXLMPA49GBVlU8n15jHWR8nXs0O7TVr2SLxT67BvWVagr68cEfHxRme7063zRKbQ+
clD5epVAhAWRpJugkDsImU4g/D/O0/oN5XC7uvUvPHOhTJEqB+m+nEcX8Qf1xmV43oHJ+CZ5wgqm
1tkyKagg+1gHfFciYI4E97EYQ5M+Uyl6MEgXGgzzgyGGj6hGJBaXTa634Mr70wlpntBvgMoSg8uA
BZmzmx3NTdXiMcBk5Z/tIt4L2I3JK+tLi2vkw3/YwEy8QHUhXY6a/4Bl5pFHBHXLuOz48KHw2Yp2
SNWnZIRk4HQ36dkFHbeyckd+icCdXqE0F179+36HRksuhnImRBdA9L6eW2qKeujIZpF1igjnt045
fHvcf6feQ4BDkEm7BcXnIkdIVJ5UfcyNSAYKNvW6FpGYxeXwt4AdMjoQnR2c044cLAx5G6n1bwvY
V8CPpiBHVetTAsYYLCJ7MtpodDkbTyS5yLlVd8mwyuwKk0Wu4wG2DjTq3KZANFWpoa/qnAF+1rRK
F9qk6TfwKbvJQztrN33T+iRBX7W+F1P9oAhY6vOAEuT5FsjaSCDG8YgBfqrQOgfTqHGKbDYSQksd
IaphAYiWyTlYOilGyNYDAPJYHTIlC7O2LfEKXXRJocj4w8wRn7GxLevUhYLQc49rQcd7HdN02xHd
gMscflLi1FZjJISBOsln99MQPTyhuxSs8LR7DrG+yz4Ney/PnlCSkTMMNnS5JY0ZzUDrJsnDyky2
84YlT8olT4/5rA6q1/cAz+JZ+EWY7uYhUQA5wv8D3q10aWkr+XDquUQTVML3n65mgTOCks8dFv48
AjjglW1R+EwzLgr5o5SNLEth8LmUeMvL5R3FYFTFTPxwvid9iVMTMqXmyAw4rDEZJZ22U4sWeiOa
y05Oi2h1CFnEDVBWhBg4AOVAEMxTtmwRCe5GKWm2qHWsCiUFSWt8hS/DGmCF+sZCK1ymzi4KZ2hK
DEGm+8OW9bMSUpPkkGkjKY3tBpbKWYJ+V+xZ3Ko3im6feflN223POrgWoNi9ma4q0a4JWP0GIaRq
362d2xVdWDtn5lQ6iScOuVCXshP6/01czJ5kfJXGSnIr5o6HSEdaS8Z84iqBGozYBM6LMTCNwLsX
d2fY8kAmPPwi0I8oWzCXyAsfvygXHXxdNBM2d2BsZVrMhd5ixmTxYmoxjvC9Bb2snc03sittEho8
z/NKRcExlFewdIo4YAa/VeXiFeH4+RL4QKLHENN0CcbuZxyJMvMizb5YPij5SBfOqyleHWDf5fim
SjR4xFMcW9CT2gTY8hyohMzZH7D/nHmK9w8I7tZ8GGRWf5YAZQRvUAMLYmXEDffVigqudkSL/ydC
jUMToR2KHV6NNtQ+JbctAKQ+ro487AO0xtFnqToRDz/Kvu8zn8Gq2RCKAJQXIHJjbSe0JnF69yVb
+fmlupNy7wGFmfeTh3Imwbpk2yUR0QpvpQGbNcLbcGWlxycfJCvtNr0/Y35MPsfgN0lkkNt16RJQ
7CZM0m1xVqJmBwpKqvQVx3Xe39o6eD4BcbpTMcdmMQJXLIoHt7hYhJIGc0i8m4E9NryLczkTzBQs
3CyMj2OmLzG5DyhiMD3N5vX7oQ+G/n+H4c+6ZctACbSJevjEjXX8N03zlHkesz/JOwjMgKs9JZD8
iopQ4dNUW75HWj84/ZrK7MtwEPKhYEB8h5Ed+QFzFymX+gLCitiwtWCaNIG4hd6QM/pGaNO+DKKg
FGLUogVywDekpj3j9BxlMGik/Fa9bE8zOM371at2RWMrk1npwGywXXrUHW3gv8WmzS3SgvYOE3i3
1cfHxT7gxcqOrVVor+7Tcg6HmluM3kgpbeBCn0ltRX724+TLDaO5NsAgQfa96y6r8DznWlvRLk0v
TfQUrMgMvg5CcmF/Iy0s0dob8XMFdyS25mfPkgxy0aH4/3T5UmYurhLXsKek1CDAGYY3WeTt7GPx
D8wAsHhIMj0aTgaOsoGY+EA78yDNcqY+Y/RSy/60oZpOtVpJ+71YC5+fP+rynjLuUy5ncsP3rpEc
5FasM/WclIql8X8GC8a1Mqu0A2nBskTVYG9knCguYRZ1xrFEULlxW/LJHIQ+cdvI2/KjeqBC9AT9
8a+LqQOZ/yGHBv43/jzegcK5d27S1YEdCnADK74oK8D560ZoGZ+fC6qMU38SCo276CQp/F7MfHBo
DEJAO/HH8kdCGpkeS8f+Beos1gj/qIegrbJV3iW/mfKRkHIUlTdAXBQsRi4PrKMxnR3e0LB7NyKv
47E4gSKz13dYYMCu9QIsAhiRUpgocCyF0oaR0fJMkyUdHhudoL8VI7xsfcRZzCrXlwvo+gyNWnD6
rIwuPeoSRSYKiY+KqJCZQrXOOmJnK+YblHQoFOqI1ywBmwNuxitfYC1Ufzgz3OdirEJOHoYUvF4h
b61t8fNfAupx3lnm1C2oFs6XFREVk1JC2EmZiM4oynW01US4f3gH5Td0cym9O5VU1/yfxDMq5sMK
4w4vS/z2IwCb3CY7Vi4OarpJi8aY5vHvtoO3wJ8JgGpZycfHpzJ6ywqg205qxdNW4iMML3dJ14Tp
ZXPhdjxzICZcRQ4qWxdRA++9+ZhJz0TqptbOopNmXdjAWh/9dDyNvfKoBHQpQLfjsgQrlPfgY8pL
jo0g8v6nczL8yCeQon/YEo16ojlMtPT1vuHO0x9DVNarC3+d1FifmlV/BEQvbzMzxLQhIYE6zqPD
JdIRxzhChkmzv+B4iIHCbBfFl5U15MFpcgelK+1FyCTOFJ/et++hexsTWCP/lqn4OYAugXWQIk24
h0NfGM9ew1QbNWyO9WIjXuFyEDSt/BQe8a/RehJs7y7iPBJFffqydzdYZs7UOIOxbxZpzcFflNlp
TL3vzpUizs7JDPYCV8bB242WZ77TrG4EQugY+gzPZy7UCqJAjdaI4abpuE41Af6dkVcIja+B0EbY
BOGn2mBrIyAqhUL9r7+JKT+AGgMdT5OTxqysZlkPPE6KM+QXdeYQ0zrlHPNAW458UxOgBN3gPa7R
Y3qc01gwVX4ROCdFV6A5iOAA89wlgQCbXPYGLyq88JuC53ebEtT+nHfnwOos067yyvd48OR0Tmfs
oeV1INC4L2EWj4vVqy7WFKaGxLPX06FuaXofpjB0jLO3KkQAk0vFnoAHVLDxXJXetoO47hXZUFlf
G2IVtoDApKFkSiwEeLjlJMuWAyyJHMOMzop5qgKhOdcGUf7LqHvkevym0j08R3qW8VMgVypDFrAr
uC2OcXuqSCmFHFB7JNvWjn5Z+7Qy9Aa2kRe5hGXg7ZJE6C8paCUS9ikO6LekBJLLXbR9rzDp91vE
YW9N89bc+AT5TYbr9XKXNie1jiinED1YGLLs0yAi/lDwI7bgiVs/XVPfezbQRoI/niauNQiO5qTe
s1Mfl0hWxGggt29wtElElm0tDhsKkbfzHPBBwjP9YXnpipW+qvW1t2oH/NOazI0hHk5oo89zhn57
08cU4/wiCvtLkNj/FfS2YK7VNhZthdo3waxoVIdBE9OrdfKuhkEQAteu+L5KmkfaLqq4v7eWw9uC
waIeseChi8ZVh1jQctx/IbN3QUEy76lE5KW92DpHMEV3YqqzAru+zk48Vfdr2CEXpa8ZL6M8E03K
HEppMsTTx0guivfTPMgCFiAtYbcS4shG/XpWyP5hFkg3j+ysCBXVwU20lXstE0LWCr2emQPiIIO7
2OYHUyz9EdxbOzb6FyLuGQN9QvXUBjIN2NtlmN0O6Tp1xU7D9WGz/SxbVwcrVLiWfx8kvgo41ibQ
xOvGUS4hYUOp/4R2yPmuB07LBwbFgo2DFho/hDU4NLWl5T/aeBTShvQiSqeBJZngzZTNO+mk8I35
p/WVjQewTCBuUqzLeM8bZEr2Tzqle7XtV2fXoDazvVDizbtTkoUWVrJS9MnEspvjNKP967vUdMpj
6DS4P/0xKjvvix6wUXns0l8l3rzPkIYps/QsmBVQt/LKi71WoyUy3iEtMQYRaQXiQFKjIHRJQGQV
bW30yqtAWEDbcf/cCijX6Ell6NmRuioWcz7k2Ir5pEgI/3+HtHLW/d9wkkIAHxFqvpM9eJ/k7cu6
w/UL0pH1IKT6AGFYbLrD4R8OrB1jtL1JfT7l3oE6TBkNkI9wBlnB/BGYUYvhQD+ECZI0N0l9C5er
+0OKewqkRPy/6vHh/QVosG3ca3U/tweF756Qg4RyEEbyNR1cGBlEkchAlom6OXmCQ2HXTbCNOQS1
4IYn8+g5lwlTpuPqndBf/ZeGEe6mfp0BMFDNEqe+YegyJGb+FAuXC1DBMTk03D3IE9dDTwp5vgjF
DX2tBYsdS0hwirFS6YmI3BXHOFtQ0NLUWaXci67AwW/WK1hVfkB0k6vPD9JtsisSSSDtMPxt3VUw
XUhbJaC0skhOh2MMR3y4UpLQHtvkcdDcUoACVK1ZcuPpLYdI4EsAQAUJdX7xw/uWun7EjyVl1wf9
0boP5i3SUs5BRZb3oQTVf3XALa2w+3DHjljGQxh/ko75c+ROt/M3TmcJ4YDMQwI50hsRAcxjILxf
km9BtfXQWLNAafgwD8dTv0rn5cl+iOcGPoSo4iBLFju9wLbjUC3jgZYyG4D9G/6uYSvcnWDmpBF7
o5OWHxM6yKEWgBri/8y33H9n8yZxU7YwvTGgp+O19QuyflVGBJaBnTFtgD3hrcv2uVpm8ufEnXdm
SPhtzdgmAU5CoKKQxz+6Fnwt701P/ZJ6LD4AUmfmaOaeFMSSyYhqH0gXANzmTo5f/JnQ/RzBlgtC
0PnGzvnkLo3gv6uBnNOVV47pclpzdM09ra1jL+zlVAEfulr/RTQ5cxXJVJLzf7oI+lvnoqSjFpCJ
G5KX04LF+RHE4ZCXwsZ9+hmQYit/6ORDgkm4wWXOJLHRUmei/1GuTw1LjEan+mKPLDGSfybaKrWs
fH9OswZLhLNkvjXOwLNbssLJc8Ov/e3Y2pNslkwhZGjicNPjjxR/dx8eIf3MnHePF0NNW2dcHfS9
AfnMAZuxddkI6Nc7OvFdHBLn4egnANTl5hhBZEQAmM2/nZXxDnszGzgc3DCx16N1sGxRCEcI41rl
AEZB7cEYbj8ifEWRwuPnxUbSnAKRIbBR57shYCYbFN4mUOk9UG+ajg/UAgJhkPFgYZxFASH5seS6
OWvBNm8Cr+wD4q0UcwJUJY48kpq98OiCB/meCMAwrGwE6CJzfv5YI6PsqG/8fkJMpCjFuNtcA1Iu
LhHh3zWSe6KU96wL7LCpdbtIz5GMHRDk0iyxh1IygmYM/miAfsQZwnvA1St5UrweQ/vk6y7GNdaz
alnSJ0yTDjsctCFzXBaBJRzeNtqoIpJmcl2bYNpciP1kmdvF2i8Zn4fmPCOInwyt6OoOr+u+3ak2
E2WveDie5hXGi6CuOqJZ2oMoF8MtHAhbuDyWcb3y51E2OuBOgz8+WubKnhuPWBCCFbT2FHe7yEdw
ZMiaUxcE1uM4ULMyNUsRmAKZrne+vsbQtJjVSJ+/j9K0iMiwpshm64e7n2t/rV4khkOHxTV8OLTj
KKtjegWAZa1pdN90iq92FaF+7dwNiaIRi7xFbqh/oJE1F24uHjvDMFofAtG44Lcff+vd0tIoE+x9
D24r92q4W0NcHXmpWAtfbipDDHf7OB6eTCJWhXB7YjjOZ3Hl/ZJE3D+cgSZAt7ONb7mbTDzW9d22
QYQmWR9HmQ8aQJr7AdX8V/nI4jZsfpTkPSdqZIO8WimQaqAGns1lkFfAtv9udEFQOr77sABQLTCa
aTGuJjzovKEncVDdD6tymY56pnG/tgkLrjoAhr6xkcVb2qi+Uun43krG1orov5Ud1Pe2MBy+peO7
NDJeyiWNVZe9Px85Da/7ZOnXDTq7NDcuNGeSTcF4oMOjGSovoR71XV9ofCmv/cg5gADGnIckUHZI
1qO8ri/oIbPP8yHo7Rm5pO5pE8WfVyMQzhGmNxxYSOa2ItjjGWCHSiw6ZCkPY/tmJ6Ha6evo9Ve4
VGsEoHNeUwlLV0JVwVc1uX1XVkO6gXhntr3TDidQeagl8g8UYybEByU9YTirgT0+1VVcoZHt5w/I
5MW6zPtOftWcG6NR/omTOas6JCEJvcWhJ0J+CLHCT/NtW2GpyVlP/JTzZqKHNlTNWcx6e3sA+l6b
HDd1GYMQgLGayh/KxXS3PIaUWYTqvffabg4W0NJge+Ny+VQt8tvXXE5+u/AHS3dhlIfdcVgCKQ3y
Xaoqq06ihcOeqqKUKI+od1KVkI1g+kqY7iV4SnHYdnURFGNDBkxdqmUtevEGgq7DiAMOifnnYN10
YP97OunKZQ2QI68pEqnMgvciLO7devPgButbCia6PU/gV1sddc9b2KqqtWQ8x1jDgx4ywa3XD/P6
nYmp5eeEPuK3fgvuPNj+h/l0YZQ+hz+Hju6TmvxvYFShqkgay+8fSMU/fHI4F4v70ykUgBNoLXNq
Bg01V9+eOXHKwgNkZRpnM8xKZea7/zKpWf2z7SVhQLmuT2KoOzznKdjYg0/qMcWaFzKCT91qaxTl
OCLPDunhszHPCnGmO7SsIsTY4uuQOlg/+yzwJj2ypMw/ahXPCWwAUl6iqzC8ZBz28KchR9gD02dt
KiC7bi2oR6l1ho3D05E6t8R7OCcIUCShHzfHwXuyhEkqyDb9tCG8WJ2OQ36lTjjpnhrwWlU7FmWF
2n1NWrKzzvjJvpYS+uMsFhJ3vBhK8JusJz/n91B5KFOXqbyue0s9glbRck9Rgl2vASXxzm1fha9z
f3Bd8AjvARMheZqfvsxHz1ilqORoV3pR5Fb08ETazaPhl69YxPcasoiEf9Quz2B/KSnvmSZydr0O
uTeh0DZ34cbszPe0ZVOEBdWrO/sajoaCAvf5PcOfdfXt5t0qO+Z6eRRtajMmEPW3D0i8We8C/PxA
xgEtQ1iB1L/4U1gc9bd3GRwIAa0Oow/lmOD+JPGv0kv0sb2Nf85S9+U75F3SHzQp849+JQ2P7sJt
xxg0/v1dL3vxjzJGrzcF5K9F69xKkJGe9lC5NMtwXiSfF24x7hcEl3xRJpvpiLyHKe2eOFZfKaRR
zqjzqLHQLJayQ6W05Y2ay4iSeIw50IRW8P4lFGzUakKzCBxM+5cNxmNXJsAlJFXR2iV771OIT37z
CcBVUuYBIfotJJxOZSj85RTCysPLCnWKMaiUZvlcQ1VuS9/Ko6T713NB2XrIYT1frAyTZsdxBUOf
a7sGFetuS3BzgGfVsfwIM5mM/75k4IcQa10MKnyW5fSQp1ThTlcxpd8eXrHRpuv1DLO0mJKr9w/6
0TB6nDnKUBn0zFFn4B4j9SqOGp56Gip9Px990R9dik2LxKqzOehURwJIKEPbSesSiUsiPgydnap3
Ev4Tzia+g2x2c7vMDjHyIlaDf7xms+BNO9mCKnN8zH4lndQkI6hcp0WryB+YH5zZ6QPagk+8ylmY
+l+TNYf6esjmnUj8E36l8YfpDE9i1owqdGe1z42ntcJw5cNqij3czm26cC96yiU/LOf3U3I02x+3
AMmlGJVN8zUWNKvGp2CWAfVlxCLZRORzbSMxmO1KniBAqr9ty0SzHxO2s3ddTXt4Q3gxsV5KiZlf
JWBE5IaO9pntQv9T0f2H3u64obFZ/I0c54j65K9qYtHkgUEj8+TeJ89zWwV6KrLdrrb69AnIYwGo
cl6n7JOMHyIvNHqYsZ8fuhfEOWjSs6PvQslG0Be49v9vVMowCvi3imKgVQUVEjEuoNBvD5qhX0Q0
3yG8by2Bn40cWtJKJgypWW4MHYYgEaal1tVL7vb9QhOH1K3O1QCgVmBboXZLJAOk6ty7pyRbS5Rp
2pBVwsFUWY9L92l2cCBl3kuc/UTDrHM4HbGVBY3BI42RGVkNp2+05NQH6xTKkhuoWIXTiWiWGrlg
W+ltA+a25FZMf3PEYkFWOFJIvKhUT0o6wz2MLq6NE8C8I0FWIbJi9THs7BTpLmarpKzUOsV3DaX9
JWr0kG3/40p9+kynWGPOROhZvxsjJELJQrIxhEC595inI3Hje6HuGSSntS6+n7k+Uwxblfpb0tBL
qhwFB4Ff+HGOPLPOZ/HSSMq73Ir5i+v7+CD5pgU3uusXa6b/eu7LvoFbOB9ScY6ZPwcajl/bjE6U
G7B/Fi7eiKjiztcHKL1YcOuA8TAbJgTxEQl2J5jmJZ8IYtOTje7HsMbVoi63zP1VUm+TTnwZvww1
XXRtb0VT8Y7Db75MjpH7Q2mmm4fquoMV7zxzPp550RcoSqMZOJm+R1PC0/XsEPLne2ShytZKAqUz
r0YLJdxx6LFGnk8kIlbwW6O01Pt8thvAZXIBn3RREd6hsGA3txnKcpUhn5Jtyyo1gfZ3zvlS4LyN
/vC2hmBpCTlhGBzeWiS5OnTnH94/95U7c9ogdPHq9Tg4hJoWpAFLPiz++4L0FBAQ4uXkTmP0ZDdB
uWA4iKM2aBmnD/brgATyBe81Wbq0IBhh1c3VhHIlVwHoCOlzMD5+SEBCygSRZv3xscrF6QTrgS4B
w5AQos0lXnv7L++moDqISfhcoz9evU4kus0v1coe4qAkbacq8OnyN+YUkLdZmv0RudEV2D+BXIWz
UFIFOt9AWl+E7gAxBH1qPZ8VwFKctMZ3yvOpLOE4bCw03ROJatl7hakYkmlBkZFbfxeLBaHAWP/D
BR7mb6BAkVP427oVDvjbsW0ss8V2NXY6jA9ClF4sjgT8ATATEqiHPikxZF0YNZEr2PuaWvS3HT1O
Dw0BE3mxNVI6GrSrvcQWRzgrblqeoYNZl1Esfa6nF0DssjzKwLeSK8SQbnxkmSd6iyw997xzPGoN
vChfWfr0xttk6MxcnPr6N7lR9Jn5c2GoECfcwPRXMtpnGth9Py9ZQ7r6jU4EviM/BqvdANgtNNCB
m1wiHqKLA5hUy8EV3cn8+17pictQTvGn/ZO7J7ge05etzSB1qB9B6NltiIKhezHnNBtO19J5VwsX
p9iYjJRMr0HQe5+Hb0qfqf9NDLtf3u+HQ+ADRrBlnlsU5H0dm3PBdEM05eYuxUHEAxpQzYtocFSk
jhQOvL7LotGd67SxLw3bBe+Zkuk2p73Ov4VPyJeXfdQdcQjtnyi/0CygJ5q7+pbvkfvflTSoK92k
SogwtGr5xdfRhMMP+qNuups3FLDh+Sm01RAscXUF90YxDPFvIPGfVRGWe9XrlRYTc2Jfl/hfjMgn
LNAYzdfwCe9wjM/w+/qUsj90wksEYwpd1KyPPrTROGq3fQPkP3vAPkxLUOL4Hy0e5IUTiWkCYWx/
oCW9a489wZaHZqxwH8+5AzhB4TxOkf+OUT5r4W8p5gH1lBMVi77YkE817r6L4QN2SAdpjVPWbFvd
sG5ZGBNoJ2Qwot0Lmz0hARx1VLnL3tgPhtiiURS8ciaqXjEOUFc4pVHIPijgXVZFpdzUR1u420Of
D/BWzPMT6b0TIZfU/uGRr3TRBCcpnHjxI34n8tXrauLVGIr1YP4f/MWPIKIvGjwf9ST5SLtAT0YI
1Q1JNAU8Nt819uY97ov2Ctg8RPRu9JogpTDwXyt0QJ4/eUH3anspE83/0ibfXMYwWphVSDBn5Tbi
s9HuPLwc9k5j59HNsCwjiIVT2sBheRhm0a4PO47vsc31gnWlPsoT5WNWPA9Hb7la7zLfOO4Z8HKk
jZ4e3sbKZJkMLqB9oepJvpNic7F6BuIPo6N73CdiwZ4p0rXyrUxVYMujzeRy0C66iodZ/83IjLZy
QBrzfizOqFlJ1F9cfbSNpm603pPytYbASs05ByaaFxt86NdeSs0HXfUdD7X1SXEV5y4C2C4ocA4k
re1mDbQR9MCoysy+RD0H9/EKLBpTWIAoqztOmdk62Fuvg/Xva/E6DVso45ntS0XdSJx96bQRANzG
JMweMT33ov7SXOnCUXYmgoD6PBJSc8/2B2jyMFX6FPFbu6luRyXGmZnMBuM+Td+dJ/drCvSHnQWd
jqimsWVq0KEh5kSbYmtsQuKcn6vbMCOhnkVx8TZFNPrC+5HtVNtIfcxrVOho8fWsQfOe0LAhChaD
jn72E0neAMczC5y+sIUphQpcVw72mx49yaiGDjxhp4aVXmwNGVBuYChHXa4nA2ZUVh0gyzSMGo7N
4fyFZvfFguc6ghxvEVNdQCEAnNOmDlvBSbCqEbVLiqaOG7Rrg5j1J3Yk9lZCb1MGDGW6eeT1DWQF
kLn4b1grcfjOJl+dP68tQusvsQvVc6zKcstb7bbU9UHCWrCQq8UHcfuDOK6iO2uh9Vp1RW3bBOlx
rPjbyeBf+j6HL7AZSfy/fXeyFxJyQhlSKSgchM53aw2jw33rR3eKLFhRAoM/E+gc8/uU6wMEzAPX
LrxHfWSP7rOxZAq4FRMSQ0EqFgv4CEANclmkPgfpyxCpKhfK++gsUvpLZtAjhieC6+M28TXVvaVF
2DLpq4XsX5Jzz/RGrYX2jGC38u9AWqAmOimZ1gtH/T999AaDSmqgGqb/LWj4F9FKmDKaDZXc+TFy
1gvupASUteDRB5925rPsowkz4iWHgyS6CY6fZROLQzUnaYRmHzZN0tHJHEgXgXNN1KmqK31P1H6q
uhjmM1Q/hwSzX0yvfG5PXsRmeFvYSbUNtg8GLt2ES+jXjd5RZmbR0VG2MOeV9JAygt+xTGOUnqDG
OL3SBQDg4SXqZjkYXOg2vK4jwVRaQe5X7QcLEWmuYU0HtKj+2LrTXpQNcZRKMxQGvOr3vkORvBZv
4Rx/H0wl/5J+ve7hgsOphRmXBPaC/kh00cfY+oZJ4S2i6UVKXf/mtTvacGOhphHg7w0AwQsTBqpN
a7UAwg00M0c0lARGMJ1iTrEaejATNVKk9NL+HW+to4HoXnrV0/F8f9yo0ttyfCSZcRkuShq5GHx/
WjiTBJrbPnGP4m10join8TlYApHcvUt4T9olRu780v7w5tf7YAhIgNhD28qBML+vPlBx8wJg6kn5
vIFfEFbu/JCLevTemuMCHueptMfRXNHVSaXh3z2BGV8CBOSar2nTEi8uLYOguT/5l6eW1qwNRwnR
Oij4IlsUlBiThkWAZZmVD4DupDUwAhAEDVrKEjwvYCDPS27kwauu//n8ib5+z0P58jmBMnF3i/68
ejuoJqa6XSkezwiGdFFYuyFIDVHk06AaiP1Vyj1mduJiv78w+zgcnqspFauT7C386Xb5YNpC54Ny
NfPb1LAXhdLloWhr2kSXRAjEonFGoq8/fJrz9vjpu/TVOR0Erq1s64uIRgKkrl98uyWMAsNH3aU8
dwrrUF5LkNUUX2HTI9h2hD36MzI/tThnl5zB3IV3LCLluLGI1yjJfrSLLm/sK70+9ry3AoMHMNs8
7GAxVr1t/laeWcyfN9qimYVj9iXL11p9UFVk9d1F2LEgaxXE+lHolm1F+ZWry74cyaP96Onf5TGZ
X/16fmiWfU6mPspA1tDyGdsacRy1qrgt4qrT1RwnIUJXpHih0s8KISip7H6CCLTUSy11d4Sn0zPx
0KXkAzbwAHOzGYkwTf5zXIiAoOnRiZU1bf3MRAPw1rMldgZLXwJxDukjAl13SjtpxVdfAJBU5nqp
JPrg+lMJV8b86Pwk3W+xoGApiKMzvA1Rdmu3OKXc99eTU98tHgWP1d91fkBCJeW+dMczg9lOUMGx
irRVwU2q3ksgro2j8BGyWMfurpPx9X40jy0yYSpuMZmFMc+m4s1YnQ0708HBDDlsM0Kk1ej2W+J0
hVxquQjQCuFA8vanjPr83wB3tsN70OMDgqE0euJl5MewgqyH80/8yKOeCEWiUqaQLlxcXy+TvAQC
ZQa45fjPH9LLeFWdGCki0Na7Wmnw50gopj66QVtPrNg2eRjQO4i8/Sj01tCjNSBR9tUXSpk4tA9h
Pzc7e1wRwVhmbljbYLLfnyxHyM7zNNdl43BfJA1YA6f683QQp1qEI19tSU9dFc4Fx/aqfmncjRG2
P41hAPdOkfRsdPxaLBzZAmthj6xFDzAvVakOKn6N9lygqIQ26vZ0H48oGYHR4TXqf9SxhNTUzsRu
C3Wqq+EV1d+l1untI92fqYSmr4zw+k4H3RqCVmnaCv9LtUn4n1t+EM2I1XkJEeXdnZkNZaTCMr61
Rfqv5Bgbz+D89XOOQXCy0jKq1qiZdbZ+WHUlmSV00d0yPUEJQ0NJ+RSruu3ua8mOtW28HkZWKNUF
WU8oJ5Gu2EO3Q3SRw64NFeagsyCicfjxm+znCOljBrgXuSWVgUrxo0TMrjx9M7fx3J6sobHPylWT
FkpTDO8mnxM+5a6Q9ZkxuOeskQsm9Sgdf/Byq9WIQf1tM5luHvF7jyRvSi0mckJPOnl6nZYmZMIu
6EPUiIJ7PUl2dqnJ3bG1KS6tCNhcCcWFWF+sTu6Zhv53DIEqP9zU9thLbfPDbxuhHw9f+xRqDM19
9sO2GKEn/PiGmEjjUMtcf4p1h7tyq9RVh7+6NQ6TjJb+Hu3bJ4k1tR9twF6nUSMXhxXxxZwyt4dM
ofcFdLqV8p3KgEnpEVlZBMfZmgBrPphjsRk2YdW8pYwZmPdbMzZGLOa/HsMnQ/+zLlr94STbIvrs
aDnR0OqMmYsug3znA1a+Zd4Vjd170K6rfDqLprmIiP96+O5c1AeKuZfPq2qKo6o5qJ2f7arooJD9
8mek1w9idihmdGEfXkQfsojt22vIbW+mzmxRKOWcPD8Hv5M7macG9C4zIWBOggxdIVWItlw9Aveh
sFYqrpBaDNtHOEE5yRNglAD4sbJPVOilLU9xK5w+S7/QJm+RvUwBWVauZ9ZOIrCNKIOMIuur8Vpn
viYcLE+JHQMusXnfwrC1VmrMRnPXUT027ep0dg1yDgLluMY35iVFW+9Bpjh5kRuAhOUOQ2zvWc2g
enaArhGnCia86fAlevo0NvkkYwMEU7Y9eC78dRs6LiP2AJ4uu/vyA7WI0MCMMY2K3EXu0pGmSZEP
+EgX30lBgSjD1WOZs+Snx5kjoCiy3w3xCR42XCwRQkPuQ7QDD8XqdikjU0WsQ6dNYQc/P2X/twmI
Fds40VQVBBOr2pv6S5TuA7F5WB5+6BwXcxSy91I5ERFMSffGvu+rLpIuUeDjVoIuJJzflxWO6AwV
V5VA3rYCzs4gEdGx6tj14qXRDHQlJ1VI3gjHr+CA82oY4aeZLVoa934+zAIniPoj6RActulrtS9h
980n4cGubdOdjS7Us1RLwfIlk7L/fPb0Hv8YDFmxb/AUcXMGIJffJ3IuUu7ujAZ/ROVa0XJabGNp
xdHREhcK4VFDz1Xi1ghLWm6t64BHcSpTFRgpuMc7EcJHkUjVjAx63u1kDya19upcXR4W2HaJB5kI
4/mmCaxN5L8RdcylCtryXz+gk2XyuwHEG7URsPZKPw+8BTd3sSiCB0IgfuXO3j8rdvDoDyrk2W5o
abiGfr/uoM73ha5iN5QT+V1+H+7gY/eEU8N/G+Sisu5sTpKJElJAwZgArKpRfnfV51qddU1sI2dW
KTh1SVQxHJdflt9uP00I7eOaVVJWMQw3yXfGIxAvFKJeXW9L5vSbZDuZc7qLOUZNdTCg6NPChD5A
m/YEkuzcpob8QYAL1hg1LAEcjOtfNNTr2yP3sWMB8V5h03jzA3VtBnkSKKj6RHCjNarxig8Oat+K
Lrsij1/6IfJBAQpYR+I6EAHMNBndodJZy9BwGl4kTFA/9gKLWRtLZLV+PsQWOqTjRZuTla/iwTnT
zH2h8fYu1UwyXWExFITGuS9bETAVhYaSbeF1hOobPwrEt7wHHPH2TOPOo7Qx1mHoPnbZM8ku2pZ5
+jsg1pvgFxtu1GWGUKaotv0Oh2D7pQMhdOzDu92s3V+Ixzuz1AfvMZc+mE6pM2EaJPBUlBbBRP9W
A37bvq/SGz/z9QUHnZJLI226uk2u1ITVrAO/VdVsWI7OZTKpWuT4cDtM5RPKUHLYPXYX342YtC5N
cBpUZgZVcga0BMhBEskejca/PR28SMt186HhNPFVfNpU0lpGD3nE/TJWLkgPgpqKOK/Jv/n3B/rq
AvY1YgY6/tjJ8h4v2kOIADgnaq/2bAnPcZPXCA/G5KMJ16R9S81fyd0RGnfjqnu6C5UoieqknjH6
av1sz1MRxuGl7lK+TcLlJNwudJlbK5q7iEAisWn5lF8j6uBhXzimo9F1xw6JIAdHqZlWjbfx5MRH
aeTpsQTNZkgStx14EqfZJ0Z/RRF02BpQR20DRode1verRT+GHlMm2z9mUEQIpYOMT1is6qeu7MjW
gLGj58Go9znl/7wldlYr4Oy4jl3YFDSc6JqEUJEzPBG9JausMbxCwPONFJ6nyo0g0VTMWJJ49LAV
LkW5p+Ty0StvzIHMB9hqxjGUwSi/g0U+mOCcw/kcbfNOM8aDUxxlufynb48JjdXn373CFQrnQaXE
+HG5sweTV+pm++vxjPk9FgBW6FKefa97IQaAE5dE+kQwU1obLjXUATw1/AFTWolKSDwXV53rWnEE
mOqTTAE4pQxYwkm0kOqULP0KpA9DvGaDYCLK9f0E1vjvw8RcYgfEDeM+5Hw2siCcaQdEbyWmQ59r
OHzZ5rOGJd8D+PvfchIIQhETPKzG2PmG5dRGP3/D/xAR9/URm1fAR0ZbjNM2K+7/6FPv/tiNq4CX
7mgHPB+sVPc3skDw0Z98WR4cNF5ZHDc9aCl2xsB+Qs4SjfJW8TpQgWPpZV7WXgigIIDx9tDd+08j
s6iwe7oIe/H5zOhrtyWAdlynb8s9frrsE3nTDLhbXYo5wMbN+ycTORE9pjzyVmPLABazndij924r
mWmBfsPtRRN8ZmCpKKBjPFAvgpx4Ilc4MHS+Dy8sVQ5Imc99ZfXAulRq2FMNcbfEyfV5ilVIlMUK
yy3W3w1s562EuK6DXON6bZRW1vvoAsrs5k3Ym6z2m1HRtwCqCJ3ennRYhDWyf8C9IDqHgTB6X3f2
zVJ8BtESsgDajCp44c/+Q5LcqHDBgU0IRfE7eghK1GIr0/gCN0MGBblg7wDUOqANCDIuY0VdxZ6w
VF6hIGpDiRdHTygPnVhFuZsqM4UHx3P75rEuDLXortAV+RJENucME3qpTcEg0DwHw2oGWvYguM+0
RupIbh4xIaXegW8RPoJAkZRwvmLCl/9Q5HoUdnkGxbReilCTSa5u/MmHY7ODiA+jNL3xGDXsgrnZ
AgGqbIRAjrrg0xA3uV8CfdKaaXV3bUg2UGInTNuaidNnGG5yzD995o1CT0NYqGLqDLluzIRc+fud
1L+3N0t6KyOOOMN2y1vU9DivVq7wngmL27C3f7RXHj+N02uvmh2kEzvxpC3VcEZd+dYTArzn6brO
3rIM9HNaGmGEmt7Plz+IqlQdiVxwxD1lEHC0arrOsKnwQpdzW5TiYFUURWBUh1cQhCxcvzvkAFWQ
+ZA2tGM4mFGki48O1KWFZpQJ7P2GADXdfGgu43gnM+jT0fkG2yx7ewoaNgSyv2VdOecuFkFFWzfC
7TQyMHipGUfzB2iOIreNVNWBMb3uUlrclxaTD7ElS7Wu8O7M7OJhL5CQ6P83mcCEqXJFL6ZkXxfK
NqoeUJGXLnzjDO/OMljDWMIVVmi5bgnzKNBdXwsWYHL+yaOKvMqzF67gHVp/W85mn0yXVI8cHutL
1Ltr39wzYDes8CO7terfMNfigq0nrkFBEpih6l4rwFBeMs+TLtKK92IT8ha6io2toeJmNtTvHgUH
Up2l30p8l/p28MXG9a1uwYzuX2g0AYI+sRGLkyoXFU/tEwm81G+z8t7YKomRNG08SAESLjpgPw4I
aYb5+m7Cza9ZrUodsDTLdwMEhYaQDY8//gqInvamAitxbtC1Cd1jRKPUZpc6mLOoLFRFwZ+kWeuP
CvmuG/klj+AK004Ah4KKOL9w1BwN+Uy/BSSmV/93IaVQ0Gsm1tezrfVgpW2QzdckjiXeSfpEvMN7
eC9u7AnQb4JBbE1z1JMEZUqvGHXIIdhOcpSsNN9Iv4/enmpyUciFJjovJywK6yZYCWYUSQX3TKCc
yq77driXuuJcrGb/qOtNzEEY
`protect end_protected

