

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Cqo+FjfIOIw/0Kghh877RN5JtWmUPj/KfIaTRt94dXWp8zshF20HfBCWrK0/KjFcQ6xaC5bYfJZ4
kTgDE7VoLA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P76DAxdsqqBm7Dhm+Xv4UBWtxeM3n7VV0uwUkGrQnJyruFJEvMXWtTIk68wS1svCurmxJblglPTM
AUuHl8lZTHelg/xsbfqIjFFpkYurRbfQPaEBBncWEUkGXitk2MsCEJd1XKoy7X9zf5gkivM+Dtc/
HmQtcrnx7yMmBEFf0wU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TS87/wLvg3wp8BEZbJFwjKct5crsKQKmGgle2kFCdS51Fi9lA3booRtYf7PKimLYtiDNKzFnNmDB
yS/M5Wwp3OXdwvzTqi7m8nPDGJzv9CPlgJYl97xwwfb/xlITgLx+mE3FLNjQYh1k2fW/YeWIYcJ6
dHaLGRiPpSzATplaiEnfWr4z9y5Zgw529sAAgbJqopXb1oauD9xMSn+2U51TKQlk6QzJOyaBGs0Z
cYN8i3mMrSJtz9+1CorRnx9v0S2lY1WHtTTmGGV3GXP4WDMI7lTnhoLYTdqSlyv31x9qhFidZzgn
WXAPS6oNxDavoZXEycPxfYnQwSx2gi0tzG/NZw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NpAOviX6Xvaq+L0foSrleTOrW/NGnS56aJ5rqqn2Dmt6YUNEPYGn9LoXqfbnr2nu7OxEo+FueCzR
GTO3m2J9405e67h9qARcSi/hF0VUlC6bqx3PVbV+Lg35W+tGaz80NE2OUHws+A7UXDQk1Cp7m/EC
XxMS909JUlXKjJHNQPk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P7klUwNMTreRZK7TaA1WE7CMMEOTtEjomJfZ7pHl1XNp0UR69ZqgBrqFP7D39H55daou+YH1hnHn
RPI1HarNWCxtLMV4hOqf8NjoCFBgrnnB0U1fZ2Lr4Pjyi28WQhnjcgxXDHuFaQlXuyVOq9XUsvMJ
ssrZQdiUjtMyy3njm+Pnbmk63891Ob2bUkQGGCsGTzQYYho8qCUxVS8K3X2BjFQusmuscPspGR3O
NvboEcmhCLzlJh3n01BooLiI/MFAc4YbNKfLIovvQV4EihZ5noxjjP5wWP91DT3v8RKOECGo+vl0
XfgG1PKzgtiiXSw82pyP+WwelLF2xj1qh8+H/w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13728)
`protect data_block
lUL0Lg5EKP7INKjYkJbmihMPHodUPbX9hcxLo0tV1dWbaTNAjiWRs5scXTC0B70nHKDhjFRRRR2L
aJroIlw12H9G/dQKV0/uTlrqRnCX9X/ce8V6GRCSwIpDN0a1hMO5t6vFgfiD/TgV58tgQEgGx1yn
rQ24Bp9sVyCaq3iukh60kBVRv8agZ1s5GYpHdOvnAEes/VQ69w0gakIVDl4gxXfnkDOwHkzOiG2h
wT4lm9YcjFeemiNViUhyI1IFCJmWSrO1gFa5UAt/Tp7bDZOale1m8qcHj/yxzD2mioN2VxW8tUSV
tiznL1eqKspiOA/0P9QbQ3KHFZxvZQhlVoJ6ib0VVxC6Dbu6BetyLxzNBd1Sh26lc+Dr6suOD2gY
3ahn+rJGb5svrbWkzBttQekTjZBB87QsOH5d58jN9Hi69zlSQ+XnHg3kQdaeaY1D9zSdXF43si9u
nMycPwm+0p7jNh3344gGXzP8WvweXKjOePY3tm9joSB2fJGOq3EyRdF03QUWueuDbQyDveGeQETP
YVCJhMETexKta6pLkyjeX5opOGwTxQEr7ZZKEAweAhwokm27+Jw6Lv47L0i0Y1D3NxYheB56NKp8
KOxWAC6AIFII/w1fPoJ8ZJOBY6BuH6590O5O84LClmSpyM7JPEryQn5Rh06pQEq063BM224CBuJT
dpVHfE6lYR39FHGf92sCSgPKj3w5Cr+JM/Gq5uezYHRI9o5+XgcblSwhHpwBe8heQ/M0SIksRBCJ
tV88263f3BZAM0EvtVFfg9xq1ywcbToRYBVXobejz5RvilvlJyOVFLe94F9+CRi58FdqTvhP0iDs
JUDpM2zr8SD1c2Ju5AjZr8oiLLRVxuSHMcaWgziYDiF8RSsmMD4MGoiO0/80sUuRs+66shGxCdpS
O+1t/pp0gXqMM3UKmmlcrVyLVi+289axdBAZ8eL3vRtKgyQLuBUmBm4ZX953pJ9HAdP5npZlCx3I
thKmYpM/zPecxdkDOGwVzoDzLCrL/YOYIlgBYny4AALBlQngAqFFrPnGk4KCNnGbw/4OvOZuLBre
S2l7vpgZh0SobypS9Lwt/SJUdsLgMA+sY7WETqm06/KiJYuKqr3eSyXTD/3oVdTPsslndJ0Dsc2G
+SEhUYh/SwpCdAO2cxdU8gnmrK6vft0ARN7sOIaL8bx4OUw25RX6ha/EmwvA+bIYKuOmYZhwBt/7
HWjYVYPcQ/qdSFXQBkgph5cwbhmyjlghn3m+4io+NsElT2J0rcwdePiQVlNjZMSpWPzNcV2VDG4h
ivAWyuyPSx7LdN6Q0VBkNa4oG2sLt1YxedSdNZgHJDxhAPuSXv8HQOieU6g6olP7oHOishu+fX2k
Aka9O0RXlioK9T6IvVCdpwqOFEIHFDPLDdKTLHsCxw2/yWlKYlZrz4M1wRLa7KrZca4Hrqs5ZAP1
4PO4EMWpRoOY0KFGthEsjQL7MRqOIIgEsrqGAqXA1BXv4VpiAu08FgsMeAU1AMIlMLWpilSbETjn
6DfHsvHtkEltkvDDqGlTmWMd+899/hfVfSl4FQUcF9bEUskuY3UQDV0bd5f1kUOwSGXl2IEFFKK3
xEpp4s/cX6Beb+OIJ07FJPnWDhaUX5rlE2ynkQhOm6MDDhZMncadU9VD30Iam2ter3g4dbji3kE4
unBDSDcw8LaJjseVroa/8Z4DD+cUSTY5rYRw9lT1DmECtoTEOM2NlCZ9ESb5SwtZT02Q33aV8c31
ZrqkSXXTp0zxyL8QuneCXKgF4Lm/IWcNQGoA3YODRxSsJc8U542tCKIT05Xagkyco3v+P5b6lf0E
uGVb2fFYXAkxIaohpXsRn+qhChqLP2Wc4MUSTOnrrq/XKlnCT4B1Igaigi9MOydrww9SYM0yWeUK
1aN+ApYLsvdsJg3ecSrMypGOb1daSb0TDRVqcE7cDstOBJd/w1Wo8EdEyYPnoYWE/HaG6CfUfX3k
eVKgbhSQVssXYWLHpWVX2IvsLw0VD2rkk6W+UyRSR5+ZZOGJ+/CDgIR5Om1OgOQVqgh3yzdBO2CA
TC5z2nOxAknOz0tDaCg5Dgid4JY28e9kxxD8kPj53dSZ70dZnZaWD+JTRLKEHkRReyaOuHuhGdv8
OIyoSAo7p+UZT5jtY/Li2xUhAhtyqXekmm2Sq4gHAW35Y/nBgvRoSVxuEoh5dpotWc7z4bupPrnD
Ffgh/y4o1I9bY+ONKGQPc6pqW2wgC01zovbV3CxJZ0/d+gpQhNX2JGBiEFqfJ0pIuQcbl6rKyQ+i
25hDlWvmJA7lQtNXRm9v78cNtqmCgXoO9hGeDf8O9MjHfOcSPlEE4qp6Armun+X11k4BZdyhNUP6
BgZmRd+ApXn0TOgFZWtdN2/7uPgCGsKLJ9q2Wtcu6YlYw4AhYE9iylEXleBwSL5Lu6qm3goauH7f
Hsh59YXk1FFFt7wL/kSLWJ4x6Z19nk1DmG24YTwhgwzrHqt9KXVpc22h2fZMNXU6gxqu//b6IYaE
UIKgoNjGbK81wZYVX6p/df7GZyQy4oQViSrcxfHJ7IlEZXGVtm3hvukrG3fYgve1IH5bqduOGQht
dzlQj9LrEt8Yyh1nUQnSznLUEXjgJ33F18VlW7ombHvkHUHKe1rpsEvJYDFiudWYLwLhZRB8tPzH
1W1+oNl6bTYlxro4OO6SDipgOJUvnbErALMatgsNce2jwAfaRFrWiUTyw3j32xKYuLrDSwlk5bMQ
cEDgVqbXmZr6SWaTBiseQK3fYRCmaQMvQs8nK0v+Avjsu1L64dDXZNeWg7+zE/VvhldBCTIGKacT
8CB/2aqDWtwGLkCjU4+JwZbMHYPxu560FyQw0go1K9U9rWEswHdZ/b7IBsWMczSR9SgFN+4S95m0
qFCDIZeIwTnIPYn/bNnC4mbrwp+4+QtChg85QHJxfuVv5V2Ry/ZJGf97yc29PBQv967U1Gc0ZG3j
9HKyWsD8NfWyKJXTiEnNBC904zdxphVO2MVTa+ybC3cvygJhDw5Js9aAT0US7avpbvMrlVs8Nw/s
Xmauf4QuANqhN0zKbYdTzA3Vu5C6kAnaYamiSPjVpOuTBpFcPS/Eic9cYN4QiQ9vnnS5tYJ5VPWv
rU5hXiwSmHTV6DNi/XYJjjgBiRsV5gPFWS/q212vSaBKnGCU+HoaNSVJq+zt09Qq0zcJinPLHBXN
Ml71AolfQmw9X9xW2X1EYjge3uI6rcj0apBhbc/lH3wLIWJCOK6iDEnnZODiTCEEH334skQGP+SK
CMFgh1fUeAXfoFaPxPx0UAmu6trlgiHskVgCzxoP806hQzqUpQut3L1ZEegINVw0XABxHqurbLFc
caFasMUyiCyJoTA+wTZL0coebTGzSPjkKPJQzp3m+3EkPniJDgi9mVJTsT9kDyZINFaRpZHqF9eg
ivqZpnOQVIXilYyheRCtGI5XYdWOiedX4PAkkty53HtWZoAG0W6EuniRkY66+/73ZDxVyMIcQpHP
vag3izhRiAoODreLFCbvsPmilEGy3t394vMPmvEptNy0QuRM6mkK2Rpx30TjY8dn1+y3lTrXcIUY
yUE3JLtE46x7yBmZJzLqiOIzp59dFNUZ9wmxAUBHyWSk1OiT0qy6AFMG0SXqeXfQ1vhtR4uZB5d3
KmzapZ9ELa3JDuwaafC8eQhaTyetkQJdkYiIA1p32RFbFY0mpfFN+VqhnPT6aXCAfyZ9rEqFJGL8
Z/V8UWO8yaHJeSF2LSqAUbRf1QXLCtP4FdlT0T0LDOW1l8qaxpsjxZrIvDrHeQpRQUR3V21JCWMJ
xfxfE0Obp8WTP/gxcInPDaH/4BhyvG8bsiUIs2CR/ZnlxuqD1YqWNXEiwcPK3m1WXTl5QcjhSqpd
wG8INy+1EAN1kzGblSf5G3aoVrkP8R4flVuppbBMGwjwP06UYIACTmL9Ru3/v+t0iLwiwYmqDGyR
lPnIxQnDgCnTLiXmJNG9NLVvsTG39k4OO5rIXnUSiaS8T7EBixkUdsC6EFs0jNoZdsbQ0BuVb37X
7MBBqUIZjE/+COPXuDsUJBLn8dCLpqrr20n6uUwMCB0e/v5BylZKnuauCqxYpUSegO7q47dMJBfX
0urJE6uPEMgSLoxdX4uIN0xBtuJ3B/iYOSWizQ6iRDP37etv8JZdzw6SUIpY1o7WYN69ng4KH2AG
Kfwc7nL0gC25WFJ8tRctZpwk+zizDlR+E6mB012arEAjQu4valQc/Vzvgf5k/YtZz0NYtGgyhD0d
J6pc/J1+sPOXDjZfu9nUzHvGmLnpRO2lawgWRA7tbykBZDwOm8J4nO4zndXZSpe+U2fgKmjMvEY1
zVaI/HU2oeGj9btYiDHxWV3HkTOH9o9OJfee9P75R5d2MEfr3umPB+viP2zWISUwMIMc+MEgK1gZ
QnA92pLhSONpf0Es3GL4mNnd/UxXfA0Fn4mTescJpx4KXy1I2pLWlrjrx2Mzn43A013cZoph8QqF
5mOSYJBnVxe9wFX9dJj3fHJGC4l1Dbix2VdM+hCjq+tBNY74Ud9EjMM3lDhvM3GbukhFJv4K9Tt4
QvN60Jrt1Ez775VL2zYz7ZFslkOoPY8wF6LBJnMOCwvilV9JAIVQXzqu4PNPMrJri1JtOx/qg7/z
1sswa5Y6bDVbC7E/jui6A0rj6wI/jyy2EoG2g6wGJPQcdiOU5mlOCgF6zZfpEZG9nZG463JXxJEw
qisqZj6aUQpZooRQFeE5PN0C1S8rmDFEtT74UlAnEln9pP0VqJvXqpNehtwZPM+0fJwBKyuOA1o/
CuYXhPI3VEPXAwLDadxoLXa+MYSX9oRG+htsI3j8EXc0u0ELyecHMiFznqT/SjDudq8druoP+Mek
QX1QxRMCFEPNmIvsUJlPe1f1ri6JvlRNjdYkL1G3EZ2xSkRyB+jkUl7e08FVwPccVAXDRxgllCT8
r4NE8vsh0LTkVuXl8L/uRcFJGwuy65NpI63TAUAw/vHrmuvApxDkALaRUWd997UpJIiadbKKYf+u
A3KaT9NYSJkU0rGGqKCrdLjWdN/cTrh205GsSmq8NbOz7h+yUR1R/TlGfwpn0DiItQLal8vVOQj7
l8lbbGMMCl8QPfmtAqUvKD2thpneTdMYHQS98SCYTDsDbbINEpXBkCgj3kTuXW7zy2UEJXuUaUSE
2Fi/nIacA59P6kSzwLsf8u/Z6r0KNnO0qEFj0xaZjJCuIAU0XyKeOCI2vGtbXxqHHPQYC1BGO7JS
NY5v0wjfEHbszHQXhEHsN0R7DQnI4MxO1PvrwCydCW/E0gLAljYmipBVXzYlwIDQuTDGbOQe9GJt
kyd16z9I4xop91rsQGMQwHvbYGLbrLYIJZD9ZjY8GcBIHDDNFFNVyop9T7wxQxEZb5PtcJ3TUO0F
kscK64L+XbqIBurDExbz2Urgyk5r1w8PTMQIPGz48norjnZdaN8Sregusz+o0WhGM0GQwR3J5wV6
oe57R9hO3uolLfg2ZRA1bFryEqFPha7SzcqPc9SFpHlg0CSaYoUTfadMCyTaCZmWqTwhXdRq2lOS
dVLM+t9HeyAQRHoNnqJ6JEKnwKcfrcWLN5Ywe+eX3hv0iIMhcmFmtKTCksLhsfzxK29EsVYjFpZz
ExcXYEtwy3SU7oiAqISaCe7DvFv1Xf13XUATJTHxV/t4JK0pA3nBjuh/7pvK7NVAEJ2R78PqxbnU
hWc3dln/mgveY4m91uSPjn2XQSF5lLPl6bRlruZYeB1BSIEXJNRaUAgD8Q03bGVKfhr0KLfE//jv
M2phrr+png6pndFygGJ00D7A9T/0rNyC1ZHfuVLelp9VzzgQrU3knpfAExzMKCFTWDGPLo/xnz0W
/bO/x2KDaecr195ol/F28hdi9VbAVCmzs9lKa03eqF9EIj/zLX/vI/h2mEFvTUmGp29vNU5OklFR
1yDcSrGKd06Y58r9Qpj9hWiw8E81vuzmGcJCD4o4il27QZq3MEl0/sD2ezeizyxig8Ab45oUm7dg
qgkiMSF+mobMve1Ot04fi2kii1xOjG1BVvOtH3o+H+ve02R01UTRhakdkeiAUxPVsNNyaSJjHkD3
anIFfeJXCnlFNfrKtkbidI0mHchNU+CT18ZqRzjiaAn7gpUeOvkm89XD7HmDyBXEyO3BIVGF9W5h
kcJLkDqTeu8AiB4iZ/VQ1rJhDhzlOZq8SJ3SK58uO55pY681P2IBzEhqgkYu3vabc7gwmFC7lyKz
SKoe2WHeZPyxuGTYQmEBEwncXTIhY6vHpm/AKnI2/GTy7Bd/XRAYtX9LxQjKZotbF5AbQBp96Roo
5K5hJFMzOlQwxA5CLMy9wwpAzoZRhQvOC/tinvMzI0rcmt4ANd9QfKeXHN4+fJwl5KofPzlH+XMf
KziDwu8l7R9Kgbee1IGsxTI1VZWZG8HKGS4DFb1p9UHpI3DnuVG3aYT0szszXBgKpPMh+4TPk+MA
bed/i2O1KIUhlLunQ4OY5Fo9XUMK6wzdw/B4azuSrEGI8mdnt4g7HMVHbHgI4R0eqUYGiEnmDd1i
EvpFD7IVAYxmx2IU5neKBrThG+qqA1yNClp9bjj3ZnbmtLtrt3VZy2gKtK9q7Qug3lBwacfiO3Z+
Gbfe6IvmGDaO3ymKT6VpzM1blCE89xt+ptGOxXyZuha3K4bno3lMgNZyZCkvUgRgS0W/vI2SQonV
pVDCYVydhU0g81ExhUHEOU92iSTr8UEtckyOUrHvNmEJe6TBzTuE2R+QFipRp66VlrBnzYSwWvXk
yVR3WHkQF0K+XkF+7/3XP++PvXrIIDtepk3WJxzZ98ajPWQOt4eVoAZd2U6DGmK8NptERyD6oLt4
wkTb8lgf/0CpuXJdJqhhXhrfcfX57bLQv6UrVxLCLmES0gQiv0fTqmbxliPZ0ssBJDBRj1CKcqow
8v9nafGXr8KCXiRSlzJXoNQkDJpDgfWv8s4mDK6gT0xMRyePpHAuBBEiligDZZiFJO+DdIg6kwwL
ut5spoVesI0ySws18bv9VRFwlSjdv+O7OUfW+dlwRha1Dn6WWWTqQumhkQ2WKJg59uAsVX/0QcOB
RfNNdsxq7pRmX+UaOkNYdNeUmb55Z/jpLv1BxlmC6dnjeVxiZym5wnqA/sFtRS/xEQv89KL9yJXw
SvRTPO9KQznZJilVi8Zmcrb95Gw0Xn+yewA1lDVZGbRBN0EyTxHC61Z0cNvDEoCDVbIMxlqxEXtR
vprBvG7xMBs2fu/qI8ksy8z+00WNLma+p+TgAhJOOqJ29FJSNUmL3lOsNHOsvZ552XXMEGCQOCXR
q4EufMOiDWdc8HPB5yUD51VOU9eJMW9JvGtRBXf252puhtN1VwC5sctVLA8EISA+tm63s0Ug+Woo
i8w4rZ30Nrb90UYqhQ0nfIc5pkv6BmT7+cO8k+eApD7EAiNhZFllV0OUYqwji23qAPPTvzs2twvN
DZf4TdSl+hwptFNHUUsH4yoUkYW4o6N2sPVEeoov0nGoEy3aOTRKemt4w/xnRGCYyXCImJd6ugRB
uau1QYHiqZjvOYItp51A5Mgx82kYRRj2HtXTS+giEjmX3GQTHhtw2uX9l44u5qs8rFJpyxhpDkiE
H/dt51T/2SqHDAxj6+vII6jczKZ3h6Ne5xAQmjr6bnuF9eseRHM6GW0JuzPkT6PcM2JOGkgx/+Ie
k/1DGqEoJ72r/Zh/xEUcD4xI1PsOVY1vn9YNiXTLtRdjwi8ZPojrJmRSAZwz7yvOl+WvOm1bzWvk
1LmsxU3Yd6IdV5prvXRBhFjIxH1SBUuaAjgcOkmT6JJFVaCwUFRkaYwED9kjecqZKBKs9OGuILwr
FKhtKyiyy3R/hTNAbe35ozhU9ZKyXL8yDgJdk797afJUKBY9PTsfhkgwO8EYDBAYkXWvjmkPjChs
mA4R71zc8HORxeGxu0ffbo9VGpbnKGa21Y6aHTJq+nJUZGa9N7TB5+80Ah6laxtt1o04ZeHbsF9v
33Ev3b/Vk2kPOrUCX5beyke8UqtPRDRetcd8UodjnGeoZcIqYketC5FFAAG/WwRkAq2H1cYJbwZ2
rMgwfJlGwXKVw3ifql8bFqcyFJffqaA7sgW4bogdadPt3PIFgoaZuFfE8Z0F3jQYP1C2w20yFeom
EJ4/+Yly45OW/mRKWVGl5oF/X8cGxd3ocN/Rt20EeGNrUFsX/rZlt4nqgdHG7O1Zu1fiHsqw5iHp
R77hOja2CFdUGvQxTrbKSdgsyWSZaxCvIjeg35HfJPd0p6tk1vFuhCqZTph2TmQrOoUQ+6Pu35LN
AXD7Uih9uCkGr8mnrsWV9XJlfwIE2OCtoHymXwIvpkWaC7gypReH2o3VPY4UvSE5T2Hh9cbAVKKQ
cgM3+RkytOcMe58pt7N/CJWvYl5kSJ5KQ6bn2aMu9zgwoU59qWpQz6JkUQfJtH03M+Bpwd88wf30
1X0ZK3BlGRIdqbMY7zPwGJTCurtofl3ZsxMnydWyuZxGOtn0qwO87+dS0L4ILYG2nOijFspDlVZG
chh9wFLQ0JYuMHhqq9jZH4PeOcltxe13V+hdhRUej1pWb993FR0wD4kPSH2TTBUEtVjRKugC/WF+
Z98iVNmnAzufsGmnDReohlK+wD4kWc8Rk0eWFNTpFA4NVnZCbbcSOisCYvMSiHGHhaIEpLlBh83N
HvLIAYK3/cop5zj8DlUnHyOoHmEKXgRhYd2KvArgCVlqDTu9c3NeLC5+6oUg84xk4WWY2/xZzXeX
3sEyA1UHxE/UY5CsWWjgYpvnP4Jb8gMMEz7CB7rvoQ86AVR1MRTUoSHOwgXPlhhAx4VYR6ailjiv
ASRSTvP+PblI/U0h+xQC1zXma0IkeZP0f5VLc9LsB74NgCV3xifa2Q2RYVTm2UK3AXDFRoKq6GUD
ixaGSXf8dEdiT85n87fz2/OiEYnlVIKUt0/C22nRh4QBMxGaJ9zjl5uKZEAGcxAE05+rm996Bn83
fxfP5U3xdoVl9shS/stq2k4NNtr8OhMJiTO/DwGkYKUQuD1TeYhpGFDkt0PYXK0h30hv07Omf8Me
mIbpg9pLgvSW4jRZlYLHGsUwEk4++906VY2ArYKbKTPRsp2xSeHI7iJTVYANILO59LuQwePe0F9Z
ZxZg29SmDzD0czZvy41BovCuWI1W07ZRYER5t6JUr2k7qhJlYZIOD1LoR/RQZF3wvUO6s/2HlJQe
75WcAYsPPZzfZ7RZPIN6m2++o9V8kuxKV1FrXeqK53wNv1DBA2fUMa6ZrwZ5HDUweQhvv+Sn06rK
PruoUgSWKiuHbEBVwkyfD+YnWnT58izHKJp28zLgPF1fN1BmDAffLhjAK5Jz1MVBvXiHpmKJA+0E
jVS+CoaHY7crEMfRLg7V7nToiSk4xJrZyQU1rpZAw1U9ZA38Nn7vTmqae3JCRgU15PxbvrBNytER
EaTCprcvipAr/mWxaEkMsGchyPhg10gO2sbQXOned39xoqNUHjw5KOH8lPjwiZ9r028AwCn8pLQd
BaWIAkXH0k2R2de37ZcFDL7y8bAr3uB+SqtbSEehI14g0I2nBsgAkuHHxuxJvd9thiVSTiYd/xdD
4qVdDxXQZFe1wTlh8GLGc7penqfSXSPDXY62OEsBS0cjjPxahCO7N7MuWVN8iEnS+OOmatzi5RwG
QdCYbBz6+yibNUDjcI1xvyp1pSxL+R2GqMc811O0xzv22tF1TTGgEt50ghM024shWsCmTKcilRfi
i+e8Zh14NdLmzgPfMDUIQ5elEJuygekC7kopdRA3aYchSFTBW4HtcpStFxSerSQJBxatNWXRciCU
IoOj1gQfBze99enwVIeqBiO9IoKwCONTTa5948WuS0lLe4lRZza2b0CPCeLouGhJH2+60BoSTYLo
7xSU6p5Ijy1lkh2LocuLXnb3HccaOdcFKtH47KUFvUaAeeNcCtSf4k8N98bSJQwBl/mEJ0EwM8P/
ULGyT4bA9KmTGD9LmIoHd7LnqvyKl1jgNehmwj7AwLzpMrUS1YfxOlgaknpopXvSK4Vc4gvxXNqx
pHGxL/hQNywxWDiVcwy7/u7JLkEh51B4YDYwR1Y8q4IcdjNjbPQXZJabpYJuR67ue/kKMRCa2YCq
HhT5A6ATaNxvJvh742uoJk2AJN7cHVdRMgdREcj2DhjJeEgaWOTQo83e2RjqN0StrlSWK/qGdomn
4lIeVOhi4EadOCkBIpcVTx2UtJiuwxZfZr72BDv6nJZTVz1KvvcxuQB72Xsv9C+t8OGUCy/mlBCQ
Qyy7t6HJpgqBDF0o5oi1T7Vf9DthVLhB+sZzpfLk6zJ4RlWJ6cahzfFPhxqtTHloY84UGWdhlD4q
ri8u0srqum+2Q+nRIBayabT1G+3d3Kx0tZx7s6hn8UQAa0l+qD0sNziISusAEkCC/wykPCMsYmgS
nqMY6UksRO8JYwdTnjtjX9z93fXrcT+S+T2gNIFTtQFO3lEp5y5Ddbi5+FeNszitox1PtE/dLfaG
fRmdXPFTEYD52Z0FMoWivYirzVfNoPl901ECpQ2xTAqhGCg9tEf3mEaY04MgCbtXYM5S+DQHWu1S
bAmvEcwd0Td1I37sKAkfonk0y64C1PTzGqHOiC/EbSTXc4UUHbumDiw77QAFvKWCk6ImeYESdv8m
jDiIQU2eRf+e7o2ihbcnIaQ9ff/9Z0q1/SDssyUS+doFVVchMIcDnLcfQOfbmfXHRJiLWX2BMJib
wdz+30vqjVrLQsMsKUSKy4JoSurCo8OBJKu4QhAtjZrttYrlSERoLG1CBECdNnb7o4VXH2UKosiD
MsIyMzO9SFxcbTcNXa76NuFmqAKk41YGeMjjCSexFomMbdUJbT2J1LArVn5e+ihThXPnKVQ0d/I6
XNLU/abJyzfjvQhSVKkQhbKYLJqMn4Tmy1YE7nb+pmZT8b6//618TvijvMkblvl6egl5Wjq3ZTUw
xoM3N+EjjUnm0usaSEbGanihTC7eV4Zb99ydVEaA/dimSkYblqUyv4MWYE1RTsqNyhu/fxGx9Ctd
uI3xJy9m8iQZPD5c8Neg3n6J5SW9XR3k4PhHlpAN8gABZRmr6vImnOOyAwJTleuY9IvP6EXjY6Wr
dWWFIF0xJOV79AMDmUcbFbkiDfJVuokad5JHbHR7EIzdJvkWxY48wnMoKfxo660b0mOLhLqxUxlN
yeXH2pUYIBny3KHAEr6P2WBua/1QNTU7hY2aZsqOUKshurOlSMqpVlSu39rw4jnw2t8cpR0qNg4i
o/WzwkpwR8shQ6imXa4ljVqCqiLdtjgVKlq1VFAdPKY8N84r77yu9XwJHb66W0eZaNyzF865ocl7
rs69b3zXyCIy8SeCU5TVBK3dYop8oX95ktE8quOQ8YUSa5V3++rSGMTv0eh168xqEfXI6Z32hS92
E2NQX8J7K+3Dj62CDtjhgeeIt9dY0Py7pNSig/qKwRVHH7mpv7nveLwyp+b+QtzLFzwV5uBmHocd
NJGen2Tsh0amxONQXcf/tTgWrDTqoWoP6xdV5cmEoEW4vgzPYqvWg2XZ8Be1aVSU4AlGVsN6QlT0
M17aWiMGAE++/YPOiGiZyOo7P7ylRFIGE9bh7TA3nhh1mg2Ch9F7D5V/guUdmuftSZzyGybePTOY
hlUea+DKgaGFC7MPiVtumJaBYij597jlmM7CQGBuiYr1pQWqgPd6vLudOpR08OIDwHoVhhp2QnUV
3F1RGLmrPDm0YLtC5UxmFL7A7eBELzlVIe8N2sEc2xDinLglpqw4pZgo0pLkIsXUieRJvc300JHc
SiyaA93zty68ENQU4M1hw2qLpG385Z1p+OxE5oWfrcvTbBirx1riD/oAxRDC07RwcJ6DPbxxcLp5
9QOj7SQ1Wu/VxEwqG7s1N3ACqMEOKkRrLsx7Gp5zSFV4tShEK5KARFT8iplV1oK+yeuatzl9SNZf
QShMO2r63iNmKPbpee5mBC8RwXwEZDoR6X8LMfu5d9kkKhp0Dj8qRCJSbn3a8JdkDNXnqEXmzyW0
SmNjhp9jqUBjqfFZYxEUw2xVgkVVhIKgJFIcEnb7o2baPz6APBPva+oPQqxc7+P5Wj7614ZyRzso
5Ojufq41jcAHS8LAvg1oyI811AqMxhBG9wwYog1ApejSh/vI4fEHcuOlT5Zv9NKJWsMANXuh5uGd
pN5NHqdtu+EKbGuZZiv2Aue0uRr42Axpv+goNHzXpQkXwpMSl2tKwHrYZbPDhctDLAe0W2k8cjod
fFHA9pOA0pxs4k3OlA8RVx4AoUs5qMxLMwP3Fo9RQO22eVDLCxyXZTx30+yLhti74LZ9j8QWUNgC
SJtw4GpDF5P51QwGTQ4lqI2Q9RIjXZGqYiWID3EXO4dUFr/B0n4b9HPJVhKOqZuKTN0tMjQkdCOo
Lk+U/GUIthd1nxFymv0oYTwzuCOi8jy1mAsh7fwrkjCjA6qQMlfJqjkeBB+8qXDIt2v7D27bKLCV
aCFl20lOJ+FNJiJkIXW4crY02DFk9zf/3kRdRnhOsFxZvgEqF+zkaT/qchitOsqzZ4qDz1GEiCfY
o1H8I45MOoH8L73cuSC7Igy45RCfyNfPHhi1ra1pZlXGTj/cqSGrKp+fc0VINm8LMM2RpDn9jENv
JNOV9B6x+lxqEe9NJV71Yom88T87hYleAkQiUUGZI37sFdcnR85b446MIhifcYW+AxbGaIcOIfNS
NHHFCgoE4hcWVFxBbMp5tDw6I1Fd7LouR/cwVQAmpd3xWRmzzBwtS8rgfii4oshrq09WcnRzReH8
D9ZM2okmmBytWzoiOnu2mGuGxFOUs2eZdusQXZ1dCwzYE5+KY99vsw+NR6N37tImwU22eNhM+ZOr
gr+LzAdh6RyNQ/I/gnmgHzg3MdRyZtOWESeM1J0Ay+Ne6y0XqmhgeFRmUPA6ajY9qv8le99GOSiM
3jwuVf43vDncOkFv1hxZN9jywwmD9f6ghCGsOEhPtE+LYluFx5iBJdM8sxDSgd+Nv3GOb9iUK0zX
+XlQLiDPR9bb7uQMCr00oOypzHAPz5+sr7vKQUK8jHEeEpd1p3HbvsmKdHJ+Kn4rab+6fIQl2aDk
6sApyPzTOn/T54TPC0ZWkvTWJCoKrA/vJ+7AzZx+S7SujTigCA7RAUDI77s46LhpzoeT+SsKxaZn
zC9xau6U9t8hho9ZDZgapWpHhx/56XSQfXmeAtQMe40DhOTvIAiXGUplIOzDPEawLjyN8HLcexTV
gRaDcbH4HPteQtPEnua1DcAeiypPjYyrIcWXRByqzC1rhbr0gCtOTxWspPNEZSYXtSF+HUx2paIm
0zahZ1x5Ktex8TDwYvilG4FhqHpEsWpuc7ka2rUDS1x0J8UEN39sHolo4CGQhkh71LiBifIIzb7m
Tu+zbD3YHnRHTPONKdz27MZFemXR61hslWOde7Hn//5lQsXEpA4wOL+rTGCW3hT8V/izgaiThgUL
JSyCqRQpGeNDhyfEaUngkyzjPmHjz6UBd0s2LJOwF6qj6B3GrdNTGt7PUNHFnviIgkFT5JoNXgXm
TSXP2h7KXRFjqWei2qf7O5tWs79PQKMkcj3hK6Jx2gr8jVmbZcJ9wGw87sulPNwseMHCo+QcU/IK
2mTE7Hp2u9NRvEVkgtm0EVq8UEFBtrE1Lj6FsTXJxpjbhykEcA08o3Fx2cKvXDzFaqMC9xm7nCwJ
HD0HkKPgIx26np9xiHQFHPmbYJF9wYcdLeK5FsHGdkUcHdy43vJSCzFlp6uZO3bd+StPnwEc/WRl
1fNfutVtzLBjsd7niZ97kHoi601tsQbhPZWv3d4qTQN//dox6T0T4EptQ+fHkzZbqvZXKT/Hxhs9
W1+SUYwW5keoH4Masd+P1Ae0kx4ToQ39To5OEhPpitGBaF0XNtSd69m7CU04jXyizb3ZhG1m/ZhX
uxR9JGMWIgcS2C2d6EoS/7ONOfewUOBAWj5SLf/ntq3e6RiVJBwMS2XRloLrdE78i6uPqS8Mwtfg
Pcm9JrmdQNGxLyn4tay1c0dN+ZyGtL3Lcv8fXjlnqLhUKCazWExkYQHt9cZ8wkzAkCBOMj149EBN
jVbFPS5JklAYq1ksqwPJiWfgzztoXRIXkaCcB4Q7cy9ShOPqSr4KQv7VmxKAJQeuIM+HICBDc4BI
R5Es6P3IITxxex5cVmwyZXdZqF13loWe/8xZqhFGq8BIKrxc+LHcZCkBMQz3+LFDdDPHdel3SQ1y
A/Pvm3oUGFtpNhg5n/ifmg7i9cMbNdut/+s8ZMr5guGlq8mgatT8JSXEqNcx8QW1l3vTsrUP7t6r
edKRf5rMQrazlVvmDXQsYku59CXfgPJYA4cJ/177N/7nTo9Sntt6d4RK19SccEXpTbSAGs+rYLH5
8ftvjyIXT4uC6qUhxxQKeAhq7N8oNg5LuCRBdiFDFH8nBlL9HkBV0sAXacbDiL0AuUvjsmrDHOX6
tDgfjYAUMV5/sVJ+jptYtRn9CvfuEr52n/m3h4USFE8PPA6I1NZoHPAlV6cpCRYqafZjGAXDJgwG
oUt7y3ZcpTc0QqdMCeKCLSSfGXpPsvM2usi+g35X/8vyXNude0fXnRJ5P+qcyHaFmrPpa0unnWMh
tsB4IR97IXFwl1EGnshwYZLv8aadsL4PNSQCq1DKnik9jW7f0l0bDK8h7HHSH7dCOJ2PbXSfO+KN
7MeahNn4DVVhDVYmW7A88iCWl08InpBZXepSOHjIKrYmgiMvEd614VRcbkuKFIrDXP7tDr58dexr
JrBwR8mbAkkbHFKwaGYrH3cfUth7ytS50OAWqqOS9m0BUY88wAbfLnOvKR0X5njmQhx98HrDOvH2
K8iUqSPQ10b4ww6d6JbRf4vMNOELUxdiKOjjaU+og1pEZPUefFleea7pWL4C2ows+/kc2KpxK4O2
//4mWyYpnJqUBxnOvO9CiEeSDNYuImk53KMuRGRxOGJtbgroVQ9T4xWpxvUUuoRGsVYNYWnepxhx
rzua4Rd/gsQZE7ADMP1LT30YfenbdScMukgujWjlszoNe4qjHZBRq4L2wIAlIK4KoK6WHjWS5S12
+De1vdwfbL1r370m5vYHsy5CoDkXsC8KZhvtWsiUqzZS+mMCCcGvay4hE6RAJIcmXAOKMoz9SUbi
AqRB6IdDuFoUdLZCZp1DGE3+ljmrLYT7tih5Zbuaq+vi+J4XDeP6QZXN1rCp0RkwoCvn101O24e2
Uo1p2VUHRmrcRPl/ruyc1MKHG1AJ+5azsbtZfi0Wa4FY4aNY0qubPfhOPy2vAanCJPG5MCfcuzDC
ik1/wayH2f8XSR9NgRaSPxvcTr4h3CarAwzwdg7z377zcmtFwipAiFv+SJnkKg0rn816rzQgZfEH
3nzWxrlqcri2uqU4LEBi8O8G17sUF9dz4E+ag1W3HRYTLSA7RqDbqDyHKPm2u/kp3tMxreK/kwAU
WzsmonIkYj5GKY1dh/HNTlozwCDlWe4uRr3h7W3hCPtizhQ9/rv8MSy/sz3GMTbcdCkH0nZN/T18
I0eaAtsWoXgF5WHHNI6cDalUQjDbpVYNkIjZut5QSJa8TXkRhkdXI4nZjQLAkzL/Se2lU03GywPZ
99K3VZnRh/FtGC3RaGH08Z8pWuLMbAtuGpZNmD+xKn5YIvVxLRG9SvVN1OHa6pBo24aZQ87j71M3
ngpacRX6TskYPx6ElD92jM1fLV9hqpTzLlvLAblD3NaJoRq3mGIqy3zwXXq4tEpXH9coSINAWibi
tphjyJRueR89S3KyRTShWR/B+MELCxA13bmgOZ9Z8B4QZXhABO1xKXO+IEQMts93CFRXDeP9Kl2s
Z2cgy21AbZrxn9F6Y38Nw+REeSpdw/jjZ7xyRTJ6yu96JzF/EcESZdraN6J5IuxkAAOYLLCPISTp
N52iVxDeijHC8z8pw0xFoILctc6XJwf2x+oPHmtHunSzx8jCDT/Qnt4YwbwVn5vm4jON90gsEI8c
re9NEp8DEiDU6GHQ4Eilqnvqf3fL82SGQND+epNkmZD4AyqGuWpEa/hCBoOK3oto8B1LNb7frKyy
c6rAOujZCU+aezFrEBp/fVrvhuZ9eHv1HGEIazsXMApr1FoJ/OnfyvYQDSqf0mOs/KdQ5aDdSj3O
JtOJJ7UDOCPUfOWMdJQME4S/FybCjHmkjete7Cq6F6ltdeDwTZA9jpqH5HmJXGfZEw6ovmaCSaq3
lXsnWhSysiSJt3fJTenpNbXmAi3iQkm1NG9tnAo6MLm1oSQVRfKIXxonAokPj2PEzsHMVlxmoNPW
IxDikHXsITbYCcQPKacGBTk+qGl9WV3YZiDI1c5RtpHmgZYoOrC73dFZhGV+Afk82IK+2BzH9zHx
/D0JYOqtdSRFQJtFuAFuKTQjIt2Qy7h8YikmezHpdGJltt5vGaxaHNWb4+2H0Ens+8bOYTD+Eq/4
ADV6O5hD641D2qAjUINfOSshhia5639Y/5YSz0X5O0jszvSjSD+IixcXL4PKnbQ8GvBFlThlaRJy
E9V1zdBz1rm9z4ECpu7OIN/KysgSlmeD+jVQnRfv6tdw0nM7Yrb3oJFd94ML6mvtKTVk9JVyNH5S
n3CHz8DYvO987BDouZ+/s7ucqamctoLaZ4bmjBU4GLeFeHArTxbNQzB5RIMEsdO9I5B+mEg+M7fA
ASWxrcFG7i4dksEicjHeSZtsZSn0Uzc5EoYeLS/9jLI5ZIQMS6m9bavDPFZuoVeYMwhhp/d83pRc
UVyNsXuqm8wY1tYSEhyK6AW9Tz+cLKVqCOnprJUYFmT7k52LLXV5dd0xKICVyMbJYP2rcOnSOhWK
QiOUcvYm3cAFpt51ZiryKksT0cN1PARXLcgimCxJZHs5C+VPAy2HzMUxVqGaw5i5YY9zrv8yTsFQ
fOEamLrCk7jClix7fkB2mfmAegGJ8VJOF+N7M4y9hGoSL0SDXwinXgT8QUQeeenqFa7Ic4R6coTD
ofNYV4eJgnL/du6ZvU3jjrgE+e7V/uuTakCW5HocABPyOk2cFXcsV1EArzHO9hbByJnUK5xFvNfz
WF3VWG5LzlLurWSJpMr7HtYaIY1seakiGc7N7gx5xJLkfZET7DPZffuyth0fagHlE/KCXi5iOdn7
ZZYdQ/CgGGUYqf0tlKVDBLwdd2hjnHjuLTGZZqcUYeZ5TmDVQJiHxTDMAzEfIBaD803CRrshE4FC
Qx9IFY+UPNQSxSQczgB8BTxZ0OJ+VsWgyV+coONDhMeyurjEtTCiICYhiW8obYkuLplLixbYQ1TU
+jFsnAVyR2jKFznGu+npi3q0MCyR9zvSQDzIzuvqD4VblMzEzQcQxSh+mBOE+dzT2985VKeuZEqO
sYaOvxDM2w9vDbovKhe3KBaLACBTJc0ARG2DqspNVDh+cHQ8D3XeSbbTaCjj0wdfyC2syTtpCv4H
9SJTC0vRN1zZfuJNJ0/TFAC31pTLOT+8aGZXU9FW3z8g1iwVLsqz1V6ELinIpdw65IPtJ9Mbg727
l0OKo/R49vKYpzC56UPotKwsU4a4ZOx5A67NNV0cdnlRxwuy/gFB9oJezB0RWXM2NKrMIu6bIoaU
XmPzVv1pdKeJTBArUxQ8x+fL3c5f8DDYCSM7REvPvqKIUFU9uwIl0LrQiCphgDPcunhGKJ3kAtbg
cQOvI86OhUA1x6Ax9GP1vLvVr5ePrA/ox2XkmhqVDK/r1xMCxR3gbwM4rSypb+0Uqr197liWRiM2
eDHq0j2DkGAQZYZk3KTAvzHshen489mhcWf32NG0qk6QK31bkqGqgZ479eI+07xVpUxyPidLeFPO
fHxT3qa5z3Ck1ao6c3ZYohVM7KKCQLmdu+8In/Mid+1QSDmIq5etdJYTGt0SyyJQ8LTj2jA4HPpo
Z1b6x2/a/beq7sTqr/VImKNYA7HnbnBzdOdcmjUCa9GlUCJWfaWC/excbDcTmdxOuMBb72VSoeXd
5qbJ0kylGOT3U5nCI/O4CQL0VINDxe+ARsiEsaTGcZB0BqFc0omFaiEKVFy7HFo4mW0NCkiIhVL4
8PJr0iaiTjwRWRVdwHXgTAF1ycMGH4ytLxOl0M4dNzp2f62FmoJo5B+63kGL2r4grJ71ynBa0IOC
x3TbPpODXhCAelBIUbrsJC+BHhGtW6n/l3p9m3cFCo3ZvY6OpZ2EwZqhxm201rK/WBzoJL12YHUR
70my/e1NY3gNqVDjAKpcvIun/nR6ZMfpPRagBJ/SFpW6l2tIE9IlDq1Jq3Y1PiMAlL+E3eMe0lco
xaddv7zUgvf1ugqSf4+3VMMJiAQi36eugqSXPMol73LXoMXfzF8eYKO95dtP9pWh
`protect end_protected

