

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g2RN5TBir43ECxFrT/y2GRXX5NGDYpjq+n5gxNTYWsuzDCjF5YeYUisYseKLr1ryeyQynd8Epzt1
V06LipLPYg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eJKP4nowQhkS+sdlDJ3aF081jbTFWdzdlOBNNOlq8qkrol2Z2K32WIgnl06Lqx6yc1xJY0X0kmV8
eOkRE5vog2ePPioAy86OAcMONOPoHTqykW2qaaCPwvHqEP73jf7t4R18PaTf0PZeg4kzgW5BQXqF
THWJ0viu+pagUeVYQuI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MDIZ/fTOzwhXm05ObJ3zkVB2FpJAN9o34cB0jHfFprFQZmUeUQ3tZW60svZwBPLmTXGm6NjoSEnE
d1b16jr2OvP7e61sGc1GOIzSD5lAxq6KYGFDCFGlb2HKuXZP87xm86ePu57tT4ld2oGvDNavbknR
LLxhx9ZyBV7SuzGo3PKuxBA2tnF6vIEJkp4n2dqwXnKJw+xgySn5xCMvJuNm4ghYOfBAsNQGJ39j
9OlCVz84SN0I+ZhsnI7KhLpJBWOyFN5hfdsD0RVsTRLOBu1rLKX6200sXAdAwmaB9xg+3o0vilh4
pIPe6hkIVYlfHVKU7Znj0kURPqGkJtm2RI+CaA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RvD4A+WtjqxHYEUrji4gUWEBsLfMuiFWzgBi0pzOF5kWQsF7tHiiAC+dbiIZv5TBKh6/SeRqqj5f
up1ybf94wq9EXJ/d1afld/HRqNac4VRPTUzPBHt4z5dEncFPVDK4ucOaLAd/3B1aieNd9xn+mBS/
wR5gmSxp/s9f+zaVsS0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NS2iEv8S/DLjr8oIhLcaUy30De4W+2t5q2cf287k87h3kSCMEoBnjvcyRcG6CE1IFz2i6ewnJ0mb
4oesPU8Xde+4KmwGSKnw2OpNx1aFtJHy7C5xPLKHuYCmY+9zM9y9RMguGvxUNsPvXEO9G/4BQZtJ
xHf97YW4qiiYtbOsAO8R0m9UHVOYT94pj/6x0Itkq5yeU0YXuubMwNfZ5ZRnrVKNyxQ5Ilm1kGqH
N2bcD8eyFlVJydABBBV388JKwKrfOh5ZHUd8//7U9+6XMFYO4OGZzTYmAvyyO7iRRKEjPElnyW25
UoL5ziiALbB2biJ+eBPz4dgChqDQ9nB8HsYg8A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16672)
`protect data_block
eQ3crrlfoUNFWHXbGQx0N81DRFaCMj+4BAIeJW8SZ0ZBVmXCDdgX7Oky1hiqeq2xRiOVipFPiVqP
BZzYGoOZklTRUfEe+nTAw+LWZlDcL/v01UOKv1L3L65wZkavIniDJQUr/iZbDfu7kehW4w0VC94M
okY52gdYk2PEV+wAMy2pso4VYqoar4tCmUzw4vH4Xeg2nAhIqdKL0qpdMLjrOoFvNp63oVOOLFIj
EE7yaD71CUmtgZmBkyO7LMCMUl/F7f9/NUOBEkuMiV7kaBY/L8C9oIIdTRNh7rn5mikpq2zA1+bE
GE9DppzbbsbLD1MXvHkvFo5IE6WcOLv59FrAHLHB4otSqC077qJBR3iJqxGXiMLyrn4s4f32r/pY
81Z+8ZSA7yHEa0NfOVrN7LmISW39LVsVXSyilB4SJA0+TqC6auqGK1O1VkznaKbIO3esOp1AChvi
oVLJTmAJi2FPmtnTH2yVHy/fbiUvtjDVNtE4AOrd59jRG3hiB+cq0MPnaIUes2vRvgGG9Ryvyees
uHHlScmTukyFobdyniiFO/zYwKOog9x5m63x9x5yVZg+6PHb0JBd7feQWmcydQeDU4/bRDx9nn2t
NxAVfOJ/eufP/Aqi8ZuL3Oi8HCce5al9Gk887n19pgCC0U0rOOWXnZlQn1Q+tqK2NOto8ZIpEOkr
44bdhEAlB/V3xhkAAF03Dy62igFf3PtUVxb4jVt3a75rntED1pcSCuOHBeq7P350s9CVFs5la+2H
AdPyjvKZMZewBLDoqsFWy6/MTkUl1PNdTOG7sdw8Qw2LfPrgMNjw8aTNUy/F7a1p614rd884bzA+
hmOQxbx/fyM5axigqVdq7eCzG0kvSHv+NlUcSJkEDfHfqSS8BJUOIR1hBaxrGF7g0KLvZlRF0eUi
RRksvKd9biIhcXG1XqdyjW9369TLRN9GfFmLRnpZtPzLkdz5ZL5ddSmu71gtvcPPQriiSDumh8kf
4YYb8H7iUmVmV5hjdcpNdj5DxbvM6YpokVjwTGulwicWyTedTFABz8ef/3ATaUXhF3h9A2XSZFwe
WS2i2Y6HWaN+xOEHR7cGWr0EvgEZ+KLAr5yHsahzj+NZUPCxFoXLkxQDrqzaPGGCTlqysAXHG/Go
eZL2cu2Hi+KTVE1v7fnwDLRAVkjUdfuwe5Pl//ZNt5R3FAQKdaTKIIfQebjJXUOG9dwAmw2J1QZT
MsZ11cRLofaBQFma5ptnUa01SaeUMphYyiMMYjLIyMLxgeOf89oRXJ9OE6XarryOGTEqPPdlHTt/
QVfwszBtiKqWsrHFpwQg5RmJObuJE71DZ6lLKSk9p1zokoSvVtqgg+WezR4uTXuJ/WoTmpPmdx4F
lBfxvPskrS2LttN4kM1J+JsKVnd9Lev7HNxokVXurTUZXPqELszz+Zy4LzJ8ZvJk4+9aYs8l5MlG
jGARKQbT4juEUAS9KKTPuhuzdAw6T3yCWaaz9U1V7NXHTor2JR/v8AU8/fHCt2+O9pVM6PyRqv1M
PwajV/P8y7zI5TaUAfPKKsqzkv3qT1gkr35PIXmRMjaAEJyp9W+/5bafrP4hxDIKLVDJoLVcdYb3
GePTdS+XzW2bCflN5FC2GE4au7yqCpw3yycmueba4VTR4GA7eq1sKEH/bNrzCYRcowwt1jz4Ci6I
PnU4DdUgqJ+hh6VkYA4rYdLj83Qwy9F3dpQwAcX1M9/V/EiZgPHLkVvP/w4QA7fmN7uUkvIDFYjP
A7ILe91YrvY3itZzKINAg9OIqQfat474MpPcYwJeEUGHIoyJgW+T7fxmO2EuTU43OMw2wQKNMeER
MwzNG5OcXyLDkyw8QEDdONmswj4I8Q7dbn3SH++f8wke3updF06wHMLDDK72uJWsCVTFuHf4fEfO
I+ut3PNP7U2z8sZxKU4jXhIm/qHRxcHlVu+gApZ+KKYUMlI9XyeypEmO3dji0Ak4yHY6Y2o9q3Y0
9LAZC5NSvzvR+AppH75OlzBlvfVmfimW9h20oWfCVlzG1DR8f+4QEOeoUcTlhYXrD6J0K1AZnl7G
T+BouI8l1OCraLwpt9jLoDcCEyzVDTF/apv6D+prW1R11kiQprfWjaRFcfwjzvYBuUQltTtQlnlY
9bKKI4Um8KRKRw0cHcNyJ+uaVEQ4EMu3px5ompf6HXZ9qPOzcewtWLEFIExtkQOx0uyxWVr+dfTB
ZcqST4swqwcsMR69ss5SvvqGa5GelFp2JFnCfZWTBhz327Ng7icyfTV0hEDvtlxZbiLYpXXrBS7n
UC/OZuYZATvLZWGyScBy/5cYiZLVKL9lkdcZybAShWX+Oc8T7JpSxOSMaUlCILA7cC4tHpVzEqmr
C9PsV4+wIGkaSYKOghVIjT+5XnwLzrctjf7C1q/fVW9P0BLu2rLCLujYI8Ph9f8DLkvEmkh6Vqqm
DYZ5GHnkJad4Qq6XvW0ifygDZ2v59Xv2vVycTMJadgbwZmVZ65tto7AzOSECZNEntBs5z9q3S3+C
/ZH57fCLRZ9lS4oTE4BwEbm3+Q+O5pgrTudmH2snjhMuSqT8/Tobz53axLkb7kgzHvuM3Vw3gm5/
vi/3NbdbRwjiAr8nG4X4j+tyAmmmZj+tyQNHPdJaTtQqV/tcc0yyBGw9zkt9ZHld+Y7pnEsZmzht
LTi/3KQqSLE2/hjhU08A+FRnp5L3ieDYbhHezv0wYKsVWWZSWbmnqHiIXWaJxgcLUylnymrAUkFK
5YAcghJcHnNlJP6soL8CZwyMjdEWVLL8KAARWJDc4TFJMR+Zw01wa4AWFEzsz4z0BXtrophGMDLx
26miKKO62DMS11GnT35FaCBVlqP6Tx23xr39JA6fJgBj525z/4PFguBb+4hhMtDBmVqONFVKPWGZ
OzIT6chdsZVd7QfcroQE1hUUtHX2h/jX83ujwocj0IBaQiBvv5EAi3XmnMr/wAvhpWAuzY/5p8Yv
4fMbQRhrk+2q8PU/rRDPrP3jW2Zk9zeysV7caQ1Bmgi9is3UYsdWKXLC2DZpL7EkdQ0lSSO418us
CnAfdQ341ih5N/sVB18g9i5j7Zo/sVAk/9XIQFjGhC4ukwnO5Y8fsXOvTMg0VBqSMm6TAz8EDLdG
g3QtB53tPUp/WYTeUBnH4JaftwLN+iH+IO3rcMTmFuCWliVrRaPIni+KxJfF1tPhH//+toxkF8h1
l+BVFUfk7o9It9zsKrhQRPgBcd4MAS5/kck5RC4uDewC8pFdtNqF64513VuCoJVlu6Pw7oIzemV4
HFhlonLVJWwUKbWJGNiFWRC840muSo2h57SKeKQFIu6FJTVdRiMkvE7M+vPPjmrN5KhdQ7imRTRO
oMonArRXFhewPi36oU1msvh39qMnG/4rL5qxT4vbXeg/6c05ljG48VZoXT+3r4TG/OMqQvX82VZ6
pFTQrYtqR+Ob7TPdfffQcYaDBDrPQff0KkCfFm+8lW/b9GuraqKq3+D8f7kYzu242TfgjZsHr5we
s53CW6zI/bbkQ3Mt4Jpiyc9I0Jj3Nsfpua8bviX+BOwhQ/CtXi9AEWlvm1lF3BCmTZR7gLLqUJGB
a0ljqk5UO6A1XXu5u1/EPqG0ASfxu5d8r1HgY9ChjY0eEdpn9lkpZBYrilNe3eVX3lxAsUY2Ov80
/nXZo9qDQm+TnMGbjliaHqLklY7fz3Bgzi65SFHZDllu2szEFCy7St+L5HZdDcyK1Z6qa21CAn3P
amnmVenSWX8vl34TLoYHVW+iGlpq1T1Vfj9F+tev4EZRvjiTcKJEBlPAohj6NUGkQychvKQCeYid
kPivypR0zXdrHUN9DVDWU2yBpB/ZM/G+V/PXc0+Ash7cQIpc4rZfQN8DY7GKyyivRm1zWaBLhnOG
ZTtiSeMmbPps4tD7/TJ69vNXuaWGcXPZXoPLIMCED3CLFQJIgN5TtPWXYdioQzqNuBAa9N1BNBRf
P222MpRxJFd3BtKt6cDJsgwq6bnIG4ITQ9ujXmKkTqcwPLWayXhCD9LsMhJugYmY0dG6U8x+L659
9Ego2umftgpn749IU0T9r12VEIgXeEiKt1IKvpI9seVnHH8GOiaY62bQmFrww2r2Cco+Mpg9dSW0
XH/Ng5neVgZuWckYUUjvYgSDU9L07KhA2UcL/LTbJnk/UpADOQFmj3UW27COpXMEVvHM+cvxofS3
PZgGEiU6jOdPSGOvs+qOvr5CtL5S54jm2Pr/aUha25PITt5LJt7XxkQLP78wgAql32FvHFCSaRmT
8WIhTvC5jGUe5lUPQ6XNzSzGu3I8OWSiPmHuNAaSbV5pQU0n8tW3+zDc4Z4Jo+OFZDZgQ9T563fh
RSYcVhfiuk4uOmlajI54xdRd/rAXNjT9OZYIENHFgP8rf0cpzRDaHubY12f3Le1P5JgDGPYWqG71
Kg57NigfPonWYf2FCBy7JlaajHuZfT8jT2Str6lVtRhlXBmmyrHqTY2sK5CRV1TsBL2NwOYlRyfW
VQrzInLXaXj1gAGkD/Ohn/b+cFO2PrWsY0mfUq92OKU7YCA9Ta7KhJryArkCO57CmnacDL7hrxJa
JlkR45IYh+1NBPQWPofQFw6iLEa/Mgmx837iBs6qPb+Hrd7lJL+eT3Z5oQijsUo5OvMZ1qOExxRL
t70RmomdP/SPBohCOn8XN+qZPlF5V6EshqSgRAslpqAwCbJeNKMV62//hSFouON6dmlqDV80fN4Q
hWL7GSWVjL/LrVXfRii1JyrZjONBJcc5Rd9VVsUuWE5Ce5nQ1k4h1JlfTGSF65CHhxNgHCyZFIWX
y7+myitnyF4WmgbB4dXKmzC48wP9zlvLHRGNuQcu7eqk6D7d0INgUNFw9AIJh7AZfilfpr5cLJTB
/EKJ0NPbAl8S0AUYz3wA2g7XEGNzkTuZ4K2rJd8+Me3FpHy+UkgnGoYdg7/aSzTPMmt33UFguLvc
SydV/6QE+DL65+esd53SQzpk/XFh6rSZuTrSbecHgRkkr2kM0hSBoK004bWjRwQatGZG8Gd7I13+
amRJzbTDCGhzU+EDzG/zC4WrtEp23B6ruFKZfSr5R/kfumqD6PjEg2EUSgMe+mdMXosNAaza7nuZ
+RymcikI2MDxju4FaBbyUf16vywqHpDMzr5c0riWKQ2OeD4i1aLan2LZHP8BVQJSKJjdvowJVyd0
vQPn4kcQcG8/XlPVuFDfPsG2w3JlJnN6pQwSYHgg9t+YLsDH2PdcCXsYzs97PTvzTqkurY7FFQls
CNsbNOj/ryHufVRaTkf4JrIDwHAaQLYgRJEiXMmp1jdgI9nTMaYKOTmjStyIxjIrn6DngAUrno07
mYubWwV3V0bn1j9nzejbxuB4WY4f20CgXfCPzx7urNl6/F6jNqryb/AVLRowGUrb0CvAZBYB/XYc
Eak+d07l4tCI6mYB/CKqVtD0zVyWA5fY6xo47hq0svYtfdUzKZ1ojbVNi+BnuCxGv4eds0Lb7PvT
iUYcAaNfG0khuRzB7PYTKvw61QO6/b92Ei3Js9LdOKqLqnQoyvNhssjhdcNvnnLBs/qFQ05EInFj
JyDjnRv6ktC711exNxXted1ryRbATwRy0PV0k3p2meKqG3LdI/3Q/y8TPzda6bDzTN+BrU6kbMwW
gkvTUlzfugZZsxY1swIuJ6w9JQWewzazAQ1+vuE0yez3q2QrOgyDP0i1V+oTvn9BWyRs4e/x6aRe
HgXJDMLVTMPj7PpPVO796LfyCRZFv9YGEDXCqGTzHwxhvv8pyKSQzeQt0lHJumautCJiqdUHLCzG
X3I9rZInQMuIyd9/5PBSfqda1c59pWWwvIp2wsBNrAjx3zjoRVvoleK3LN3ps/+DN9Bhsy9olJs2
IiN8bVEinG0urpPZMWlp0zcgKVeiQyOIPyZKszNy14h0ntWSVA/MwXzUOfooTQaxZJ5jcv1/n/BG
qHoPm2krisrXydIDjk+C7o067hKRFLxDjo0cTHdxtvXm34+2cHKvpia3RxRGYXp0KQ+2RLC1tGts
ZDEDAblrAz+ElTsqJ1WtiKYlE/jnBb1coqLmTBmrCa9VjrZAD2HDnrcT2YF93XJ32k3Qdv1p+CbG
HgZEpYywo1FnGacKJ6evP5BJIkXb/0iFs5bEBCyNiSeh9XfWFBwJy2vygUxoFyp11PP3J3Cn8vUK
V3c20UnrXR7o3XQMKoQfXquOoVWNAKhpxQR/H3NqngfNQY0sZyrvuxbYW+LPmYxeCMxGHRtZlXWs
kzhgxsklyHLnUqWRnNdohfKqHrk3ozMOi9emtwBEIY+VcMYFbemL6pHfmLwcCZbeFQr/zz5fHP2T
757Uqq7f64pQF7p6u1l5JbaFE1OySpQ2dBI/qFgzzS0/B1mAG4rPrH75lkJiHp6wzjcsNYndag67
a6J9UkgoqOf9t98uYuzE2BdArCrvhnYC8pzzYPIZpAA3OAiIiiNpp2IjE8T+6N3HQaAULawk+nqS
1qgEvAUmfXZ22LRvTlOnxKHyXrKlKmQW31arar/cymAU22tl8RrU4bo5rY4vHLFCiATuBUmSlF36
voMRDkj2zYY3Ek6UbsQdjV9SrwhI6zcmb28SwCAXRk/AC9O2S1ronwhh5+OPpUz6Mx5a9zw+mNq/
ORfLm++TMAD9ZD7WhhEBHmGwp5MCZ8War9u30Aul/74xO1fTiGdOWRQ651e6vyZIhyA06VAh9zyG
G/y4c7GCwdIdoQB39oFXn4WT4Lk1yZH1hxgxiKnRlg4hijBmK+g7t7vWWUpPAs4rXYzlpjvTkioA
A576ZYZuRPQonaDRS89cP/I7yWWzeuc9Ap+gO7UlUn/IChTpfcR/OfOO89zMi3ycq4GZrEx/2aI8
2Oomq7GwVh2j1y/A1qTwmp6VR7mcIGKUUVq8EYTDW9y2DKusmHnPaI0ZlmYcEebRjMquq62KjB+r
RPV1wX6NyR7N9gfUdRthxUDG+CXbDFMjGky2Pwod0d2txG8aWgUiYxuWxKzd4vKwgXczJrCsXKQf
WwGTWOgDh23fwHreOK7M6Qiy2eZbyc6ZnxBkYthuZsp1+2k3E5JRUQPcZ7iDQtbeepPd4I+Zq7cI
du7Jge8TswuW3zV5bBFbyZbDOMCEUoivjRBdO9YiSRghr3pW9/c85qvcMSdrbNtb7J5fxD7sZtF7
Y3dhRrZBiWgY5IvvtA5ptN0LG+2eSzNzMW/vYpsXYwmFaoiDIbS3Hy2blOEyB5ogfTwq4WUYXyvp
/iS/2rn01a9Gj8mtTiR6rKssgMjt/kAQMlHLu4ybbOixVSp7tQoUSLRYOOiSd3v0IFW4uPI0Adek
CkqEBhVmSPW87qvuytYXnALD1NYP3uSHmKRqfbG6tkG3vedFKGsgzLpCZLcCxqVhrXzshHH3XB5C
BDYH5LtKLLxZhVpyeeWullwCQX/vOcdpoTjNlVEW9QQ0GZBvlVuB69T7NNfymMngBGZyXU0FpI+7
Zn5mt7VcXxlBBaj4g538/nHxR4hYDz8oeg7WKx1ukszu2aVw+akMg/vMlLJAC921rIJgW47AXkbE
zTNvaoan1mjjpY+RYeCKHf8S2KdiHPv/h8f+NP6vCCVqqBzq3AV/mlUSJQKwnQ4XgeZCHyAdrp3x
YHwxJ5x8169GPtbVshXUU+wdy3BC8UKhjBCywUIGztoRGA1GsYkpL0piFui5q1e+C+KSyV+1XffC
mfX7QVzV0/OBNEElGiPkk3gid3lmQh9F3Bh35842wh09uWLE9pobi3KX9/HQh5Ckg7/MYTjcxMd6
5WXQwpTqeKEzqwLvEDsuQ3giP4Bszs3A3osA20CYD102BH3v7hPrW3Mw51q4XHPx7crPX8fTIdOW
6MPtwHve35mOok0+1eAExArOwg4apNW+sd30kVGjfUtHhjVYswt+QBWkev6Bq7t8/jHBAOYfQM8p
WAALA+CZzyi+b7yrc7ScXbR/s/rzwXULv2EpoqQucelwGq21U9O7eRUfD4cV4ouW06inrEeFI1wg
SY83r3rd7064wX3H5QCHQmNeIsHs3HRL6ULgnhg2BJquYOdqLR7qaq4VSye0Pi/rrG8vGWVY0qxs
8c/BCLrT5SIcb2xVBafRpik3FkgEMZ7GYovnKHagr1AgE0h46WF35FnGFMEg7wYLgLOjPX2+1X3y
fywt/j+NhRHUZZyTw/uMf4Adx0hxRLQU8wT91S0Rf4iUQmCMe9Ac4kpmugiFkX9DN3h0VTUmKQDe
1RKhpJCJWUgT7v4A1GD9RB3USpwPoCh9I1hDA6/84cM224hY51NrjLFCsVARPZxWLMjAh4glL0hS
T5B7FJowdsKTjho9Lxu8oC6BvbF5WVSiP8dulq4ctUs1yPA4DFk3hmeg93cueXyhuY7yHfKPwS3l
FPYUivqJam1N/J84sIRsh/+QQe7sMww9wdAjrxL6nYj4EbfKo6qKcFLgj1pJkxH9HyUiY9V//89M
BV4Sk4dYXXIl26l770bW8RTd7CtXkMVQdDfjwGvd4K0OGZsiAq3q6iW2/r78T2ICcxO5HK8y+9vT
nhtA1/Lk7wWRyEmzXpMIZxPew86pxphHRrribha5/d9GNvs1oaVDKLCVLk7CsgCrbFInM6aIy3No
3y/us2Lndtg7Uza/IhjjSRuCqAwSArEov9PgADPRXUDnksIrp6bHvwVs5jnZqtpHTslylPj1uB5j
up7IUPhE9I7ohY/ji6uW/gLpx2l6gCVt87asKuu6FrJhK+GBJtIdWwILDXkZXUU2musWkg/R7Us4
8BDA510MyVMV4i2GhIHQBJygWTIj/Kr83tL1yH2s4qFJTGaSDDBG1/TuIGez83ORyZ1ffAll7DFO
9yOcb1mnjjPqe+XcoE/7VcpAxE6lej5TFHJnLT8YFpCNQkPNTTlcBUsSuLgBFM8Hz9cig54ad8Jp
V/dmFE3+rMrko5T32DmRgSifAKgNj1aGw825XbdqcLa/7RDi0qbSHdlol6xWZdlWBoCbITLCq5d4
Eizux3nv6jRrCMJKXOIGc8yngKH5mHvr3XA9TJDQbKLIMdtsuwB2vpr2+euyb+AwgUOY1yDmeKY+
Bh6GodHZPgJt/IPD5sY6996ZhqEA7X3cA+fMlHCRVGZLGa9UaF6Ayc2ttqJ2Pb7MNQQZBoJqVKxj
liikGBOkmL4+xerVl7pf5mVpmTZVa8zAiGIMDB+8Z39me8CQjNB1s21GvG1PsfVnieJCnEdb9FzZ
FAkeShrih/y1jbWCZrjUxmqr+2YZQ17Pqos3jD1hvt6c54YWDOwL2Dq4yrRjMxcJf7JhIeNqcpCF
seyvXEzOMW+mrH9eau2oZe9SnGC3cQ0ERBxMsmrjqdNKfLuwTfUH1AZyXItKvOzIrXWFTkS8nlQS
OsI5rxWXRQW3M0karRxchEXDpScU00Aa4CL/EWEARB9nxb8xgN8zcO/aAlUn2fYeDE83fw3sgrxe
jQIMDshaej8jIdhZaRc5PfPLY4DJyo7Pz8+gm/yhTbINlz2jdwDtvhP0SYj3UF8hhkqfB9TM3hI8
WbBmEQSz/h04AWCIR4DZlvV0C65TQySexXY49KAM1DKYJUecJj584vTFF2d05AK0UBDxcFU3fO0s
oTMM3vDDNisTVoGk7AipV7tQGeQhcIHkex7Bt+XkeStdGDgGQClAoIA+vEt7aACwPQGbP14P26YD
stMBXfCEUwmvrhyFaNiTJNley6uonRnIEMWjxaR5Qtj2v4IsOa3wIie5RaDa2WQLq2I0eQqUmvmc
bE0L6L9Y8mMprOtxJ+sSiw5E9e90vxpTG1WvB8EEjjD/lSHffI5lUFH+bkYBMlUV58ASeHR084Cj
EJJhjnccw6A4xH7ktlwLlodC3Z8SversfS6nvumoSwKKKzx/irHCeEXu9eSgICz0SykRit/gU8Ti
LCNuj2TGjoxgPJ1dDlDOFZmFL+xX4O9qmqxBZswmdAbkNx6/jpsKgkYE0arB/2qNstC3XOXvQ1w4
xP1tbbQFkqFI/rK7VNo/KhFd65yqUW5VqQ46eoKIMnUge+j5hKKk6Eevazpidn4FuDw8M71JArtf
UkVG1cu6udY63Tkj3uB8bNApEURPMqUELevGs0hYSMitFanMSh2/QpvyEgFhdtYJwtKKD5mq8xRS
RaUIZj82+SYTcZNU3g5pqfrYAWJMvuvhCuCNs/omEvFIP/kTzBOjZQf4jtyLrHJWBeri8wZFoiiD
YWKddcDj8IDRfJM3IX/HIEe2gI4RX6Nr+IGknGu1cbzlJ+4vR5xGYB+Vk7M3vfKCYFyNdKB2UneZ
+fWlc91t0s58GbXxW8OOQ5m1LVreDSB2DLbdMw0ucIrGf1tyR4XDCfu9HNBMP2hgWTzxtUBGR7Fp
Mqjwj1aWHfQ3rTWkbuu8SECYlw9ltU8lS4rDn9xeY1VYtYNOMQVwNUCwwSB67LkMINqXGQJVoOrH
2HV4lHH9cVvRi9NUIWZL0+9m0F99r+XC3f4fNWUMKNU2LPOAUCxXntSXgM2U6qehp0gT85+8cBd4
JygYjt/jXbuslWdFMxkKdkI82OCqDwDNDMrdZu1bWfRqkoKkHGQgdoQ1azZePV1ghqe+9FjGWTi9
1sStl3s9lwdslZpQKtGKxFkNRrQGHpgb77IIOrcgWaZBAyDbOs6cogSDs8U8esHtVE/OeVGVZ0Uo
YQOzuFN3WeaJdspzGJ70KZt7u7UCXTouSlQA5nuqXCtl5bowazpfU4UGoVp8VttNpozvu1FK70Ea
kdw3O3F9UiVopAuQWLdS8Z3BvYv46SNfA/ISH2TOhVRm+8Dw4aSqb4qzGgEh1U59YQt/fNyFVNl/
ADwVikItZAXAJBd+cR+jr/A7UQZmwegsTDKWla96vdLKawudzkSdRYf1dXt4mN5KtHdPGnAVU22R
/+ahLBfW8yElTfUoNnyemyFrmpmf8V8LE2tcYW0d/uhZRsivf6Q+UoF8ZOLwUfvzfh248qH0tAe4
FvBkhxCFsvOHRW9lXDqBoDcmolrqt1z6nchQZknRgLOi8x6iZVGvbgh3XJgqk/IR4o/cxTrhRYlj
/nw5TVmTEb7S4xCgeqGGfLZ2cooMaWGutsFtfgvw8wCXZ7W++GMhHu+tFxAUJ3Iznu2ukjXak+Eh
KkdIfjSY6LAuS+V4FOy2M3Ov8XPhbhLMbPJCMUYJDnv3C6YlNXUTmGqZalAtVpsgWrT5DP6cJlF+
nH3ZECpK+AYMT5lZua8DOoiSy1XZnUuUcvYO376BnxlGvTF7rMj3/HAntsmQPcyQXFwxRmy9TW4M
hXhTTopXUnxZ7EOawQCMPF0PdlldAJ2xecikERt2AbjM7BF7Xf6zowBpPIxiZuhZ92VlxYgGJFMC
opotXO7zfYbzFR/trKH2ZvdmFNkKi5OppCheAB1iyQfOp0TVl0ZRkoT49Hu2uBCy7zM9CFNyHNDy
uFVLrsdblZwKGAl8KrSVDcV1kdBrqzit3vWeVTYsHXMNi7BF4KpQeLHXDn/Nxz1N9VtjyZ0gJdMk
ZY7TdYcrzUJDZLMxY2qm/h5zZxwHraYwFpAO3iDx4UzTNsPpeSUWQ3mVmCsCo+Dt4Nxni0/ztTl4
ujlDqboYP5PGQjteQFLHCU3xe2A9E/rXMYC8JzRujye+XZH/l/MNgU6JaodqnYuEJPwYTUzD6tdx
bETZESzsuuJ0udHuBCSIVAgKiQz/CQlDxGudtB6jy3sna9t4bOIkdV22bP3mn1msiLTbs0C5ZjiQ
lcZqRo3Og8Kn//Mlh/K01EhMZEUOHCB6Na5LOzZifbrePbt0PUxuL9sDjxZapZ1aaQfoW3d6BL0u
39saI/gCvdWrtNwJ0GzHsaPXbQhjaRq42FPt9F31Yp1ZAcvmRkqsX3S0YOooB1IXjdop+MigWFob
P9ymjxDqXn/7SSTQCpQwHJCv6SUIbdC+o6J/k/0DEgWSyQC5ASKwknBlrSwLv5UWpCIWQ4k2E9iZ
yjb+nKzPxmerkonPnPSEDAjNx5oJm2klW197vGHV8DyyAbHLEtMlrubABJ/fAFtwOhHdCBJHZ5Sz
rMFQ40XhF2rHrqHSHJS9lLE5SYzodqA+r1yIUuoqsNTf6WQUfgQLagVN3RMe7FwGSQulD0D7PDZo
7hOm5mzb25U+dSYXcPL2lIe5zv7TN5CPxSOC4kCaHBXuuQ0ggWRP4FO4svSsnU65HIgBvU8iAVNu
DjyHILcMzlF201gut1m9M0jrKyHSfpJpG+oivvYZIv51lk3OQZea+Wvk5Hz2zVlh1CbFWIDdHwFy
HtlP8aoK6gxgUsuPUrGUbR7S6rtTg3Y94gRxgWr8PuWdwBB+BbrMELj3BgEk5XDXPtNc878Ti0/d
1IqSgjiEnj4SuSIgSt1BtOtsluO+AtQq+EBi6kqchCJq2TPY756AKrQHS4qIB8m47tL+Vogh86PT
vQA5Yt+qU9HDOcpEiCIw+MYTqBpzlOiInhRK0xiUEOAnlFOYcMrKGZdN5k2zziEJ9WXimJJgVq76
0r/Dw7BI8TYq59Sm+U1cDCVKSdn4SMnAsoUbmDryLRDA50LdXi/8V3/HNTuFjKnNkuW51f5ztmZV
yD72rH08yx88EjWubiPXM27AmW8i5o756wsivmDr4yJk5mQ+NgAFYse/nKbDE4yxetUhlEQCzwok
sAXk5+R/Le6vZss9X8vlj4k57rp68RhQdbnNSXCfM7WIr5OpiKxTLbrssYK3BQexFfzwIZex+rvD
Hpf6loT12VFGSTxrv7JHt7gcBS4dK5GCIG6xU+bs9rbHRAlELKZyoUVy5bR7e57v+qGsGWCERIzM
uXoj7ui0LIqZLL28Gvs5axq6fV3aVRxuGaBbm9SvNKtl4AXprqACvSlF5zx9PPcMGNRflX2PkGz7
pEH4qQxMApof/f1SUodg27K/CUhcRMukgKvVDrqwOfms1P95Ozf7yll9y3fgkQewpDUzGyWh02Q0
bO4BrjuSCwiO2b9NECIJ287gu6J8DDnpwwj4kEVazxVEEh8CmYg0MQKKKwE5dA1YyB0bBNM1YMPM
4DmbIgMiiT4ViiMLCGjoftmz52e5PyM2M8FMKazGZW93bNLsSVzFU1bEzA6Vl/zIsUboNKiUxuqG
5g0OJpsIvSffy0cSOUUZtmeoQRx05QX8AhnEuAfALeDZo8y1Hplqduym0zj79yh7g+Q/s/4uRb5M
t840PhJqWyw4Aq2VZ/bRhiJL0pSviITHV3Fd7+Wafl9WKcbO4VL/JqnUYSx8c2Xpz2ZfTpqLqe8X
5gOwAddFU2kkHmOzTnSgzOVKhCM4v5prXxgO+YXsOcbzkuwLD+b2Y9o4hQOPeVV2PAYnKRT3jrGu
HoKlgiTO08XoUcrhj+q2vV2FCP3idKKq2I+ZjXSoJ8ubDY35Huig5S7xSASB8gbXcFA6/O+3iIRV
LrbyAyqupSje6xwwPTiMXGnyO3yMwd3Wfj7hJ/yLAiEi1M69GvLXxlLsig/WHJgGJbdtNdKTWYfN
HnOllT6Bhv0WTOTvgPwnWnT8SCQwlP52RJcXyDfl2O4Hlw7F84QPcGP7XbNV/Tr9hx0x3JHlkGwK
uRKbFUZmE6eNCDAJFbI98ULNVGm+OC/xSXBvR5EE+MLOa0GX3gZQAze9lB+VO9adFdZFAMGjag1F
3vd0gErSIoCWVkm3uNeT2yq94Q8XY0whkEwkuQ6TUAWF5tmZ1W5bcN2gIkNAo1X9AgAOs7g/9IfI
8kP9IjGZlyCZd5Y17d33NXvKEybnNZqH1Y+t9N+Rs2BEq/isEgwZCFffNGxFf+k08lnZwWBKb5gz
PxZdiySd/P08l2MnP2e1gD+VPlzJl3yVjzbMdu5IxLR8VcIb3GHaZaz6SmmjnFPmB7hryxKYkwoN
Xecl5fHEdFL2stSOeN4Ae4CxNBzhDA5lyO6ys/VzcyLTuPuSt0rxOjvw6IYvANnZyIn5nBYSQeaK
uWxVHUVJuXxh9VWUmDfFiJZCqm45LcX2tWMe2l3qEL4TYmhYFBFvVCUG5LHseh8qtsBFO0maw9l2
fdbZGp+7djDigZt0JA974/sva8POmFN/pVSAsZb48grxr/oXL4beI0LbFtg+6ybkNdpIZlDl91Pj
qzgXzs2S8968hvZNSmLjArSMe+dt4pLqemyCp0NXoX5oCYMyOoVOxKmexTQW0hozAzMKJ0wQvUuZ
M3bgQuIvSi+4B5s912S2y7tVdMwuiWefdHvx/770P62VpUrQoSbu2hcP3uhW8/ACmR9M/nC1qFzZ
vK1PTl0s3G7/bDvcvFbvXWRqR81VeKAD7rQ2bRK1mxnF66uc5a00CfXIOZXGzPGhu7FPCbUgjNOg
tc4KRN0A6B0LSX0HF082F2u1JJqho88pFvMoUGLV41G6CMUKRuNZ5cP5kCcujvrxLsvpRZDTy/jT
e0jJ4yDMN/YKpX8LX69ceKWw7rmXEv6332rVspT/40ajOhhQv7+G0ZM+6wjqaT4FvfdUX0sDQ0Ui
ekAXOug9KsebXqom3h9p5+d//XctofKv7hBsOai7DEO/Wd4/UcKrJbJxRvnT/pmKVdCLkydNUdoa
TB2ynMR5T/Ow8G6sktc4cdlwLA97EoWD9YatJcE5H/KIzpHUVF/CVXteAscqALh75aejEHOOI+eS
BwOvrjvASEQfRFO0WCncAGvatdaFAZ+kpBzCq8VR4C5pBTm29WtnCrOysIrmdENZoytkQAnli4g9
dc5a/+9p6aQWEmF5srzaDfb0/7dba7IlpVCz5tdpkiDiT9cTxH5KTO+0sVjiXVOBdFCfNVzT5pO2
ieFckZl/1hjFmqG3dpn1WnEd6IArYhD+/ubWUHgDRyhvRgj9v4v6im2KaBKZLnkivS9kjWzyPHj4
WtHR5n64gNZmTx5AZTT4oxfedS4GpVM+3EgTZcHWQiEk1eoPwwijBNH5xv2ZltTHInHYJRJEj/MX
uhJCGWsb5/cB8+RAAoMw3bhswRu9NMw7DNR0BQFgczEEqD08/NLMRRELaRO+wfTfCETYMG0wb3PH
vJTh/B239yqaeE68dKj1sV5xnh4/cMovuovJ0zKm8gwYPe78tB6WXYLv2NYUiqTtMQApyL4htNlT
7+3Nt7MrUvjhcPDTTkBVI/xfLqnByr5StxixKvOFoTehB020AJKr6TI/wqyzeP4pQ5rvCg+mScEr
c98VJvwu+VCqfIQlEMZqtMCko61yuPsnZ9H0fllVjNpb2JCC+UoeE2zceejTJnAsktZDeYUQR5In
H/s+vrRKZ/N4swvRQZZvBD1qcS13lAK7JyTm2Q8MrD+JvIhF+/LIG1USIvcQHkQfiZcK0dd4nHUO
tKg+ZBrvYE5y7R0lJ6I26n4c3/WiPZ7g/WVJEHWHz5wd4r3Bi7VmZoPWMa7eGHI/EKHh/870ennW
l2Hq6dkwjKbQUrcAyeKvOMJaiO9yagV354sOOwEkwvVjLEOvS9sLVAKf0P/r11iEuHsPPZYC8ASN
ulJfAFum2Ns/2u3GuQ3awwabHIu9dDBMdoWJK/qX9k+A4KWOFwqyt9F4UOMi+/ql0BHma4DsPoo0
8/nLNFs4Pnd9LgeHDh6alVcqZPkksL69UZcZChoJK3EKLcl6XjXuOXb5wj1wjipYpazjr7V77MEI
86KzFkhsLXPcopPgQj0UnIuT0BOSHMjSkMbXY1ChE31cSbO0TB6m6ZObEgHev83TUKHiScNpjxpc
/WSbjIK0UlFAyr4fFszoDkuy7wtnbaE8WCStu79j4dBtVgc7+6JWJMFKTYCLp/HzhSAF+k9usGaP
rve9b/rsuM91sH/T/rizERy0dbbcVbBKV5GAcfPyi8xa6h34TIxNiqGWcv9qZhkVSz336Gg0wLqU
ylerWZ62zUhvN8W2NNpDU8111I4gVbT8NSYN6sfjYTC/uPINBMaHUqkka0yYpk3+RJdiuAvtGhNK
Rok9Dz9UMOdSne5meq/X8zOICWFiUyK2a1cT40jHX5szjDh6RlKq2ymTfGzP7rcVBkDwzlr1d66N
fgx9Se7L2lOjPZhGoWCEPtrAMwI2qnaxY3cpPRXbtMvEw57DWcAzD/1TetCbzfB2ussvUGo8mOE7
EikxIHh2GrTXDZ9NBfjWGLG8sg0BZWTmi11Ajga9dwOWgMwhOCbnOUSDzQegoME5qnZmj5mdIixh
Acj/AM8Uvs/pWRi0ESxo0yec1OVsKwHbM6ZMYSjgI1i1LfV9c4kR+mt8KZ8I1eLVMUih8CFtO7H+
ggGFf7lnKJP8zYuzgkFXBXiv+B7HXNorYj/KYmIiM4ZLcsiXxCpuCzaX/VV9D4H8UNptc8YTfEt5
s5YRXrUYNDTh7gg5SfV3qskPgafiJVMkGPgvgkDtjH9cD+8TCKRBt8z7o/VEdjtolc2TCptkCmGS
XDGcB/lFy0O9czPFAkdFXPN+nC0ZMic9Rdo/I7aNFeuCffA3o+bJmsBbN7ag1UoZfndXs1FP/en7
394AFzsGrqqwdc3Yf/mZAOc52I8SvMMNKAYjyWmNP2R2YhzvGWbCpxCrS8/WvxeO9fGAN5LFifuM
+VjSC2SWEP/MhP0h5v2RoRXN5ZG9hF9ilM/wk+QGpm6MyAohVGz/dtUWCUB/iU8RYCqVuubz1qWq
343rfJXDNQmf+B7eRT+oQ6odlKZ+DVMBdL76bn4gPRJ6mNZW6lP+GY72TepuaJ3w311VOmzl9QcS
gRbSpNhhjUNq83yb4hPIggC3CuZClQzkEZq96BcsGIQWcB0fFs1GxfcZG4ZETTNp7mnpGIOBINfE
qvNMYZuKmqUWeEdPNXQCOMD0gehUdbK0atLopX+t7L8KE5doPWhA3OjuJI1RSMjPQYlJPh5r7JTW
9606O+yk9Tor7M3sLJh2xFMttymyAAP/Ilv/a15jO0q4WYJdOZXe0o5ktye/J1J1X9UplTOFlz4g
tA5PivgC8o0AjKSAWfZqQ8TQC4dKF8ofyZq7HOaYkM8Ss7yz+4OP4nDnhXDyc1qPJMwGWAudIyhF
JGqshd6IR6bEYwDflCqVj0b0n1etWUXM/IT3eaT8yMrb/V75MiMDsv1DtdTkPoRZ+t3iY1qQ/YMY
mFfReCXqdgSJXKzD2azHSIZ+3ASxzkCJTMjfdYqMgJaRJ+yDtZyY3eP0AaewEB1XAaCKoXycdvCm
syFnoe+MMlnkMn3hqTFOTP+ssgNigvqeO40E7Y0sb2ec2dA9JGnqj5VcgnqytvApP6098t/eEzth
fBwZ0Z8HP1JoeubO34GGkdru5OCjEECL7Q+2J+WtEIfnwrjASzvjg8J23/QY9YUy+wryJA4oykfj
9J+9arOy3k3uiuRzPq9ufLN0Xcf67M8evHrt+D8hs7r0+z3lkQV2BK/k6/OAWJzG99cT3CuLU9fn
LEwmkX+++19Iru8PLhI8n5tRyK3dbR9gzXwk/Bf3EUPlJkcLyXoBNZ7GY2WdbK44UdpULin1uCc0
af22dnQcJsGS8XehIYyE2U4GPjjsF1kvy6wrCHpPCjjk2GHznTZ9RRK/iM1eXmskaXg9Q7arGLZi
efcobkH2Cn9L80hz+Z7kWrbWfU5+2u9LX2ltK1j2qdWeNAgyljitVTxx36PDr6e966Wk3n9IUR+9
d4eDHnw7s8PzFeRnLvUIapRg7CJWLMipohC+c/+teZ83OIXdFMgzuyzR8KjbR18TLm55SPdqSlFL
8aOky4YxItYFywRK4w7f5/GFOPS+TtVgmMZw4KOTeTE6NfiB0TNCAJ4U+ydnGUFTgJ4pqWWTiN0J
SDUkMaTgi8eQE9nHyICmdwXvLMuG8HPXyNuuqMYHSWTMbrSDBShft+MhWV/zKlDSDXRuGFyzU/WZ
kV0ORe+0iWGasNVCvwCfnNe2wFo6fJjPolr8U/covkme9mxLX9BawgB8QZJTOV3a5JRmbTB1gcq6
y5TY/IlW01av0g9cHTlhMgGmIK9I/4OQoBFEHvFwb7CMa+/yC/QaZWN4laMrYp4X6wm+pQVGWOnJ
iDxuQpiVboDxNiyQ5AhFGB4s8Dw1008kvnwzHZ7x4wp/AG54ysaHPpGXxVSsdXzTzp1De/0kozHy
/Ds2FEadnQ9O3jfcVARziaYBtQ/7Qjo+GBdSLi2dOtXRk2vhqCp40vb5HaN/xtp6YMdhRGj2Bf9h
GbVFOwoEE++z7R+ZkF/Ft55TMubVOdQxUZUHtnpns2b2LJQuE35nctAOPtOGR3HYvp/Ww2aXzjQA
KrQ+mpI62Rsajdl6yCPss+2TYEqIZu0sMS4bssbtflu1c5EoD5vtZfwxxrClbJ7BnINXrLWdbGdH
3on7nOwfL4+xMwWRbB2CvUuTy1TheJkLD2kxkl5PJ9DOMS5u8J8r0VKkNfItmtE7Rh4xlye27zpa
osY37QamruA45ciDoHTvRszy0RMqAsX8c85s/ejb34YWqv6y6DVhVLNHUV7o8Pm3zz8dld880Xfe
Spn96UpAErA8fFTknLdFqB7yIrL3bL0v/UK8gbP/AF7CsIvfDu63+UAKn5IfTWg8kLhaxdtkLhcN
HNcqSNPiAJ2VWfahmxPsyWmzeFRyM0Y0SjjlMA0mBaFpqnLQdJvCjqSqZN/41n2QcHpMYXEpwADy
7HtfV7hxwV94jN2z9GzHDHhQDphgQIi4wOwFEcQpNZAnryqhVUNw1nbUngCS/zsW39Bf3erGZRfX
CbruqgByzE7A+d9q0icFQ60UHS7ZYKh5FTm/uqVmkOCpxpXnnV+LkK2hSeHEPvSdtCpk57L8i98D
La3He+KpmzE25Wdd7xx6FKhzvcsl0zTGjpUHKFKm4v6Nh2uANMayfbl2P91rqTVEtrpFDfDJi1Ef
+oO6d0CXgm70kmH6TGJkqml7dAtupoGtF5egaWkUcvKRyXK5x7EXemb8ejT3NH1gY1Y/NX4QR6X9
sNormrcL3vc5b4GDcqtONdmT2g9S18KU8cRbjEpjahvKcMvX7sgAenu42cxmcSVNhKtJzs1igiMv
MhYEgxViEK/rF8nCvF4JgMRqiSbpsL7zfKCQ+QWkP5fAtA5NNkNF6h+n5XP6J7X7/2wq52R8ZFtm
YP5TUpd6gMmXLVpefFCigJOggHZmkWb78gUlNMvyaeKbZIz7wFUP4wasqVqBbn6kuupbkWFzWz/P
/ju1UrmtYSkN/JUjZWQEIG21G5n/MxGjjYw1Mx0jhgG7IClKXuULs0t+tD+hmDhpp59p9AXaE57p
iRTjbJBGDOI4PJ5Cy/nHyvn/H3e/n527YYe066Q03wvNxpcSCvI/vyq9D8MYHD59AlKJKUKMjT0p
+VUUyKoSVTP+06VmAzmzetAsbL+M6VorzqGPOXrizNEtZKxg6YnOiBXQkBkBYlKL6SuY1wtSi6d5
qxe2YrJL1elrUfmed1hdlgwWv2+R4Ma21btF+KfGmaYHyLy7LUehX2COA7BXtLhuVpL1yjIdLvRK
BkVtGmgi/+kzCUG4Djb+/A/Xgp/nm29VwtbnNSKdcJWypPYCu/pmhUK78Lctx0cOhMXlKbYI0owA
PvvJH5PnV/vGX+iCVsfNYPatZCZy7qnx+FkKKhqmJLzg8rw0xHU6bni0kmR5TG58gi4E1liMmPtQ
K0Hf98bQyZFGQ1ZmTXhSFniS+EwBJRWphu8QXEtzgsi6safjNm17KsISbEzLPmHldbMx2YE4Sk6c
BXSCCpA8cCLlJ3F/dqIgyyOC5juLYzKcJcsv7mMZ00pk7FGkoP4GDuxKZIZ8lJ7peOiuMQ4ND1uw
nYaN7535OysDfdA2w4HoS7rdpFUCZIolMwxamS2DJesQLgzmF3bmY/B/Ow+cquBp3/nHYOYkkOIw
N5tMnsciJqQHMZn6BJL1mJhlvX0cNBU09ButzoXsGzVggNmMCoe4ufI5irNxVa+khPLDeP2HEX2b
k+w2rGQmn7iEvIS52tPiqTelxy0MmCcNtAeA0IVkZrkxKb6G9NWaPROgObmonuV1T2E7wbjL/zvL
35fpiFR48/QgOOEBjWcqwvPGVtiKgKsYK/xKvsyL0DK93/FqXLVdszd2NOdbbr1nHzPH3IcNPplU
5XwRW1ycDDdWw7zJ5KK48wM6WCPxFzmOX8yhzil6xKrULMw0PFxogbGJca8YMsT2x6PBK0cunWg4
I7CJWwKv6cYKzZTQTxinqewuhI89eSHUbPyIVKGGJR8iLfa29kK8VW61l3xCGEf275yp6zrlAZ2E
3REOuon7wbQwMqFp9k1Gfnc/6CWpRqY0xaQ0lD0SlRvoKXgal/9zIGo5w8f6BHTtdHjjmilGlDgj
K8hNjOQM2KmDj70/VKN2erqR7unwnqytA9xaG2UMvo6VnlGnecwTtQvipi6pLm33qmLXCDOIl30W
W0mWadyktUJ267+PzQXlNPZ+vgE4aZMVtovXBleQV45sadpJPKigGcJOtUaqzCvlzJf2gz69E2ZU
MiTg2rVM5Wnc3FwWjawLorfA+4IuTQKFz91FpsVHOylGZH31gbDEJRvKrURXH1Bqxzzw9qYRLJOq
XVSfdZZ2aArvEhxl/fTMMzJvLNgU6OlZ+VPQ10KjjYgEm5ezT9PI6oqjthUDoCVzsXaONGhHdg0G
QsvWHbqGe8mcUe/qhGo6HAk4dEei2dGAQm94F8LweJr1pLgSaowtSbQ70WhZTGmJNhiNtCYOMXb6
5ETslYIf3SyhrXf3OCL7zwsjxWu/vwOq9seDbf6nxWqDhM3H00aC304IPvKrhc8Tb3QOdYMDCzoJ
ZUaLzmbN9oZBgoUQeWp6/3pSenYGEmfnS5OOwyP1XD1zdB9f5Q2ZQ9tr9RdnNDWDIPrGojJ0cZXo
CpQzyot+Gv1aekh3qDG0TJXEquEe0bOPiFIqg81tAvpmxvPQQDmF4yvwKszrDwCYk9sBvfzoUTT6
zwkdMaD6eGZqs8JEseNyqrKrbOHsW4uPY/xnkhOkeARemXgC8bywjmOOFkhpZK5k9ecoZ2AzzGIt
05cuqKJbnEl8G/MyTz+w0Pj5e6m3zXiIJnR4NcVATdjCLtTVSJBPDmSDMC6i0mGn5FRSAYM/ywQi
qB+Gx0DQKaRbZ8RJLmGhG1Xq5A9sqEea4AZmn+dNrm8znW6guFqmD1e7FCljOgrf0egEIjVTwuup
FKum3PpyQSJ5lLZk8ewobK6quCZSM/c+3hW/kWJC47TUquUJksv3mJFRjUPcLzX9VdThQL/FFkuy
oALZxk1o12wqnmku01ddqYvih12aQ7n7+yapuEggYNlE9+5XDpTV/K6qAtcX2+KF0dShZiBHFvDX
gKUTzNvdeLtsMV0exw74cHOIKKzuU/x3AVmQJ7kP4ljPbmtLgkc8vq1wBdXRrSblGHKtFb4Rjc3w
FEzHvwQiCt/7TFtROcYMx5KxnOxHY3x7WEDQ9YGgzRhQXa9hHQbT8L2kovyDR/pJxuA6EA1M5r/7
49UuvFR1Ii+k8PB/+XCm8ap3esoIkFSx7Ud/fuHFE96cCJ67j/IDHRSr3cBtDVtQ6/ExK4GFwmUX
Pk2oyqon6twmGeAyc3PXCAu7/FcURZ6XI05cvJ9mRXhnwrHncpOcFakbcq1JPuHzPT4L34b9sYzL
AySs3COSCzoHjWp0j33w8a7JH58AzJvgWTOkjEHqI9jUyIy67ill4JzCxmH8oeqr1RTQZGtfFk1c
Lxnna5R0KBGw0TjyriBoFHqmfXzTCZ0BQvnfGSNw89OujSNTjAvm6yb7g41IpNnnECPDmq0Bd/Tq
M6h9DaJfkBJCtDj6D7FBi/7NmOLQtolu8mXGVTZOCeY/srrgJpcK/5VZw91v6AEWWD3+KxQTsg5k
dBkieRx58vmrNMOd9VUnC+ku07YLAmWnD4lmOVoSJSB8dtqL6hDKMX2XYQ4FM+BPVaF8EKQXI2kc
T9kt4Un2ZMjEj0iftHweJcx/FaUyhj1crnXtCiDrIZBtubUuQ5VfH1iWsZxotWypybT6Rx/LXGAz
SQ6lesk86iWdi7HIvusFKynS8hHq3p0fG+ZriUwW+HXPB4LiCoA/vnzMJ92CRrJRaclLHqwZIdU/
i+Nl2IbX2lUfPmbdeYHneHuvKH7WLKEes/SQ/y1z7h/1tjFUcPlFDmic7t4gHjl90Jsh8IKReTT8
kNa6dxPXBIhc0/84MlKVg2MTuLtcWSUTld3zzlbevJqmaI3Pn4Yr9pQhbqIxgJJ5Evel3H5rh/GX
g2X6b8mmlC3EsaZnHehCxzSJ9o4j4pt6hOoYoQL2AMZwtuQTxi/6BNpgdg626bi4v75m5aKSgXqK
i+Q1YOod26WD8vJtRfjPv0dMRNQjgVbSc9K05Q==
`protect end_protected

