

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hajT1eUvtcpbI2tr2ZpQ+yt3wRoxz10Ck0HI/Kzj20i705g6DeZcP+FvEeRZMeE3iSuhECQss2IC
TSZjW2KB+w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
i/I1IeDYXVmyWoncZmW1nYLxm0OqNFHolb3NRcBcmjKOMCITsjC1Wrr+uKyOyNEAzg8LAt8SApGl
0BkTt3hGlwT5vH5JpMyxisp39DIoQ/2rHyhelRgIJSLTMOjHU/hpeFRg/8m17ioym3ZBfIcVRSy/
8YqL+H+Sd5EIN7orPrU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZwMv3uHNJwRn2Ww5TFfON6zTPNrPAlVNsMdpIyHdq6Uz+3GTAES373CyUHUP+cjDCtRwMjqRzGuk
B23rvW/CpivFPlGt/mLvn2R/n+PRdHgtaqKJEYqkidXp8VZscndj5Jsns7Mg2gtWutKvoptc7/8f
8ZVlv3hAdKdz/jYv3JFkYYsQYs/9EMmUObpsbPxhccaLaqAcMcp2DPumqvxQeqn7235qfdKNrMcr
c6uFXng8fnfR9emT//lppNqdkpAUWD93PhLZYTwVVXcjV4e16eyGLhyZTZ2QS7WZbPAkj35kG18o
nJcfgFC/GO+Ysd8/MvmMgbWhQocjtlk9D4Q++g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F+8QLMkCmxgohq3I7y+DAO2INd7sZ10O4AWi5yw/qOjlH+MDCzvNaVws6hhgvB6On1+CWzlrQ+vz
8M+w5LD4ga5aEaF2/H5jzH7q3vP0dvfZN4yRMhZ4TVDJv5PjxyVU6bHIlNhOrXl3MF1oGoVIjZ6h
IEpVBqdC2ShJgsN6O40=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Nc2OtpFQZFg8m9MEwwFrTSX7PqIQjLT0ImG8RPKmLuLlbhKyDcq1HH6KjYM6DTZXkQahd7sF4tka
CU4JtMixX4Y8KRzlmswh0FCLw/Aoh3nJlGD/KZ3QsZu5KBZUxKy0A3ntWjfTg1NNZ+tsdv0ZU17t
6SODHMUk49BioUo7eB0yCXF8PR27Zd7koQvLbFKTXZjGgj0ayut3GjrNM8A+4/o3G/elRT5WscCO
qhmVtlygfHoMk7BWSkupTlNlfF4owb4C7/AqdxneLzHPlGWymyNm6olzMM4lJP0A39+MtJZjtTaU
VxxrhX4xVaQG4Msik48gN+qH3ORiExl++4Wttw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25536)
`protect data_block
qUidMM5D7zRMgtp/ijxisWOPWgXsMWBoGMEknCu6Ck46Tudeq3TcTkS5iTj00UT8TMv1Zc5+NyI3
UbKVUO0JccxwqLR/swrIogSdLBk6BFtnoum6hNp5IRDf3Ta8VPUANVEswzfKe27aNwAdAr2nrP0A
7pm+pwv80Gn0iObBCGXimPdI7y5ElXmhlJUuGyP4K5kmfAeL0sWarBHhHHr5VyeRhJw0lYaW7jS5
LWxDVL+rvbDHjB+AFMUmtarLVKEWCDHO0EqePYneBAqKxXCdAL/6eF1ehQXTu1HoN69F/aYQe1GB
9q+EuoUvn/bX8QX+1aXeq4czxPQzoXR7VmtqfQwLwwrBF1eAggC4y1SIkGxfzKmfLYln1u6C3U86
lRi9FBsPDb/WMrm9n7jR85/2UFEX9IC+lwckIsDjlO9GMs0CfwDGgHjICCdaZ7FPXAW6VJ30QkB5
20AOYyiAMzQvjpTuDrRHLZRTqDvJwO7wtYIoM2tWKiVZIXGY3iSG+0X9zlh6nDSfVZEkJJGURws3
O4NiKGH9VG93eO+W6AZFj/9VIg6grBUf2O1C5DQbQxebVZoaIMiJnp/75jNoS+BoC5Odl1O0IDqE
jRDqJyCefYRXVa1dDN+iinqO0f7zkuYiiMeNdln2SRrCW3j7NlKhXLDJ/pQHc+RdN8fPqG2K2Kw4
mYkfaSwW0ZwI36dsjCK15zrezfiKTg8wjkW1MGzJ/EHnaSwTk3KW21FJARsMGyOvMZGhxXuyObPN
gYuXEzwpYEimNXzUROywiyaWdlCNAwPxgA8iVVQecEzmifVVsLnkj3FqmgGZtx40LpJUfhtfjfI5
or8QXpft0HEzSNLAKie2/TRPISn53tW2daMDoHvulyN1PEzJgJ6rA9q9hWMGb1JW1ViFsqQo/YS4
nifM1y8CS6ffo5fxyIxYSXGcoM2bpiE7a5kGkO6CmCOdOWdVgWfPGoZjfJ04KbgQeDCgrl5w1HSn
MCIlMkjxvlNP5aWd/SVOOVaa9KNWmpqas28SmYvZczDCasFdKa9UsXUh6gL0urEnwV5XWFY7Q6wa
mlFOh3QsYOVXq+pM72oHo0BFe/Q7nXF648c37ng2hBDYaJrWQm6lLfs+9G7vg8KF+aueY1Bt1Xnq
K62b+dnTrX3J4q5tl2sFz2fYYemZc1DqlbfEUEoWhhi2jll9HEPjKzX3G2l/SgE28UftpFwn5P3c
yiJCdwwb1N1LdPX2c4MypTT5fjhUMqnKG4sCzOFGJ/YcdhYVgBz17DPSO8mfUHkQot/b9jSTKsN/
n/T/EiCA6HH6Kui7Td82nWtnFYScOuDrqg5BwEX1yI6rspiGHvBB4wIlWc3pQJYzw6yH0snWCVN5
M/3FrcoRbwx3E2lABDavpU1WD+zz3DyZ5E3g1H06Gy/XHAJsL+UObSfaOnuYEvvY5Gol0iUkiwZ+
a5ELNDwO9XKpzWuXFTnJMJE0B69qwPJs8b726RiKKZO0RpEfiTa8EFpD3ps1h60Hp5osstQXga9u
ZXa3cmcQ0iYaCgFqPcAlNks7yKMW8LQxqeT3amzxdzcy+b1HqYn1uaL/jI7k4YabqfP2KXk7rQkc
jN/yiRZTOLArBQ7d01Orih8jWMwWD1k3+ZiCkWKac8D19kjmFnGkVkHsUga/srmvUl5KCJ/FTQdU
RYqq+bzhXoC2EeWTNsdq1jbLV0sBXHNKS+og2ulMbRl1YyY+wW3qhaiIINbiREiiea6cQI8JiezO
MHlHa0QbshVm0hQ5lLYpaEQp8B6GboUX2LTqSGxXLOC3Zvqg4Nbo9Tlv9lv3ZoeoHP8KHLPdO9aB
KrCvjKooaq70CW5PZEjvm1+cXbCfaiAfgfDF3KKnX+fswcGMnrBNCpR942wt/ZI7sm9c9UyPf7Nk
mDeWXQnZ+6LgFP0p7OZuBpCHkjGa00yCn6h3tcJZ815tT3T9dCQwwwNYe+0vrxSQE+I+08ncxFD8
Eg/dx/IP6NFHfnsHIclmuRVecx619XRblcDErvThOdO9oJnwDY0aogIAzq2J61hlBTPcSssETmor
yotbH8iSdkRC1a8CEzWu2xEIS+j8pyA++5/KaiXAy+swuwMcI3lyDK1xKhorV96lLZLyRF81W0nO
/emyuKNGYCcQtfrdZxlBrRkCmZJ3Qxhtd19YOshOLEMoC72Eqp9eaoNIDLJeqtmxKoV+mrI3sU7l
nsCRLG6epP21UG49hPi7RZHePUZH9UBCWjOi3twCDH+Zn0lrDBSz68otimC/3IDqhzIIPPkDA89u
dKqDvBGg1MoERxp+sGOFdPTIpweb/p9/il6LGNLhKjmJK4WqpNPLmrVZYoRe70mn+9nzHHrrS5TA
/v6fsbu9Qqwr3EHOvKkI+bS3t9Ox8n03F+JMNZFohqTUhbuC8B+vThPJpB6Kii0gon4AQZirxAaR
7W1QYNcc87oF9sFyWw0i2oA6btbdlvjqpWyfpeESRqk7twUUZ9sSlXynuYnVD+qSMSZN105duSfy
sN8mkEK+pEBHBR09EKSUvuJyw9sn2tLsOWsxOFOy+hB6CkoVbWqFK57oNslr86N5tDujEnYvRq7i
v9yoNbiuPZmmE4aW4ENqxkMHBY/ViOcXIwH8d6V08gIjgIEv8PUlfl2fr9ByWrlepRfkxL5/2uku
Jwa5vNQBHi7XdrclIySv1iU7Njlj7zuAF882s1R9w5pLgYGNVKfbjr9xemrJA+q0W6PVKXlfab4p
RIKC24SAt93o1e7UGsXExqGHWS2Pn33LM3kB3b87ifrM7eXv1oezawwgHV90TxivJGnxWEStLGh/
wDL+66bv9uhhVcBPxSW3QW3ewi8ugg3tOTkUvfl1lE8IXb0GR83Sg+nGGxFsNXwd0UKfC9wTnc9R
K8MnDVeggj4CZXtCMLKdFbUMAPyG6FJ8wybXS+KMQ5MzzQgpPchpU164ri3Vm+W9WB6pu06B8Fe7
XK6Re0yvaIEmUya9mVVQhFkHJDiT4MavjCm4Zf5Z4NLmwz9/tiqo8gXN/5ezJoHFwPKZO6jks+nm
Pbb+Z6rdRq8YvN+RAwpW/E82MritT7QxI9df6jiBU2ZyF1q8mpUU43Y+IKOMrwPhKNDv1mRPs5uq
+gERQ6boPgxcZN9GhF4RRm8Z0zQX0lhP9l1bn5G3jPpWN+3y3m446+0jT+jktYEAI/+NrOwQk49i
udOMuWNzdI5NEtTdpsG42abOyYs6aBFv8Glo6r5VRgw1k44NUmoatFSrdQN8R8xpcrPtpDskG20x
l44BbBHTHCvzt3H7wQMMYunXiY0epyS5JeCQMgOgbKTbDm0uikuAuT8X5GxryMnm0TYizVaW7gQg
/+MqpOf5xLeploE6YVu+s3y60bkytqKmVRjOh7cs8Fgoiz0EoY3R3c/yUrRqv3hLEgqRGaFkh1Cv
sAwLPlVU/q0ehVXvxSD8N1igb496psfDGoGKJJK3tRGq5RBX3J987kmp7PIYgFzwIB+Kb8g3GcDI
nU3IVQwrsoqSReFSa9aiJjZ2IzeQSLrsJ3y43KCnRMy6Vu7ybL4sCP7P6w6VMm70/RgUUcHT2pyy
nbQaO8ZkBbmFh63bKgOmf5NPpclrDRiEcyMJ5G2JoDThfnDWVWVFlnYM4Ef7NxDDum8VUGRhCeuu
dkqRBPsTmepmb/wSyWlXnJvvWksz3ot9GJP1nkEa4C2Ysl88jBdTX0KVrJs21d58bhhFc99pV37Q
/pvogyeBvIPvcwk9LfRhV1wvxGFhNWmyHF+PxT/X7B0p5mQ6Vk5KZ6DrkooIE/tod2kKPGgEfrXw
k8rkI75wAV4np7Tj8JaFBo7lFnv7xzYGQPvyfcXNJ9Ikd3j5eI1jzalpbXws6nQ3mHSNtS7euZ9D
PmB7375/YPZhYtaIBVc5jKuaIJccDqMZMbcRrnk02cZ8KZfSukk/fbajTLiYfObBhTuAGfz8Pa24
pExogjEL40dyLGoJpZc3iuZ/SJt4084XCZfLTAv4bGVXexnONOSyudveyUQtKlm0xlEO+knU0Y6A
usb/F5qAAZulNs9W5MhBUuwioaUQMZNuNbDOdQ68jRKF087Chnv1+SxBOWjyyMmHw8GVJ8si1VO3
QKjPK8PR/8B1s91qDhnOrlRdIP4/RHPaTOmnl20aNkxYWnB/LhGIEfrH0c/kZ5Qhr2TCFXYV77y6
9sA/r2SB7DZEoTwcYGdxAOd27J/a540h4NwTrLp4nndsfzYnsysdpouabgQ1GSkKaadQ5nwvAVW9
iWT2m8f/paX00D3im/ruyIYxPMM9sJNH0spq7jdZ+00LZpebvJcetVQqkL0zd5zJMZD3xNvwDA93
/1kFe1z2Bctaf3fCb+9N1z5ZumWx9lcQYPkJncQKYbEno4MxHaUUsTfTHNNRZOJFT/cebAAcPMSc
JdVslhIbUnEf60hC5Bh1NBhwTvHACM7wU/MpBqJ0EwR9MONyg38gg8ydQqL+FaPCv99HHXiSA3uq
DnUo6oPDXMbgZdc8JaRIVIyW/pBIL3snetDvF0U5hvbaYQr5e2kc2KNuyWfw2v43E/piTcYanc/U
SbFovGd/q7w7Fl59+b3QCwtguVXbuAsKe5VFaTLqaI1QdowPSiB7SX7P3HTDNWwpgfTWUB4xm6YD
e+3wDFyFtuo44IBOH/BX8yMDwcI3vJ/Im07YpBpE8PlrnNAjA8JU2vq703o+0zILX5tn/G3rahu6
ebTjqpfoCcgzcLsOgmWx5C1YUJx4/XtiNYD7yByY3tQcXOMwh70DdbpaKCT7nT9ohxTD+NtD5LUp
z03IORjgWyLBaLohh0MA137hsSLFZxErdv21lIp8NyvgPnPFDpfBuVM4BfyJzoHxiPCAo9gA/8Nw
mUjtUO9jUw0W4o8QKpRmTELb8zX4X76xg58PXxDfiiDlOZzf76yVa8zUnQ/NgKBtsmOTwnxEc61J
WLtMda1XXaPqzgQMFSyIJ2G57PF3D7ER5PxafuUFuKE6S8as0hEuSNgmIVNPD6Kosgf/P3UDol4Z
VjYT9KiVbVCGy/x+lv6DP84jg1qBIQn1pdqd+I23vmdeCXeQvLmtAK+KY28QkD0KW+Ke1RMeGYRg
HClBsfWdV34CyCHXsCTSJyMw/+a8pqh5g8rvdOzvdtIryTr9dH5M3s5TP/zsURJVT3+pfpQsdKKa
66hNIWJwuhw37k+leBlmD3kuIu+qVHDvQlqyVu8qmeoXWV9j2Bp60A+YVOw25axoAlUFBwarpe0o
3afN5eC1BjNgEtkmB0WSSWe35nN3lEkDOEIt02XKFSqKJ8r01f8fdKM+0KQPMZmRrO5EobWlJRhw
HHMb1NkXQnyFxqpqeL9ZPj4K7g6l6K0ZhRx8vuVyygWlsdEvsAo4Vw5xmHXphq/EwxK04TwFK+ZP
MM6R0975f2oyfZDdkCnLhfhBwyo/CLsoG/s3fRpn50HhLB/jyg827pPZ7897Gk5gVaOlHXHUmOXh
SMTzi4ls+oxg9x+ArHz43tFeDElhW8HMHNHP+1r8VgBxCStG8D3zH1qH0oEzDgC80WQN4mQ8kySJ
xu5MHwGRYg5j+Aslaxh6qvrTz+MYkF8zkPrlYSeQag1bnb4rw4OFGWg8bzwW4RvhZvP7pGwjrvM4
m/rHG4LzTbPr8EbBwCeIUDL4FZyB5Yr6c7j+lm0qpspP1EqT0CtAnsH4jW9cMyoowdfSTmYiBtI1
q+YTnvd5LumDW0Ta0vqlwoFXGmpivT+gKsagzxedChVT7WZEBySCYUYsF9R8T7kNvIaLI1iUIrt5
/QlFAh52+xL9QstdEtk9yZrf+uWwTJ6Iq9UyX4XOc5ZgJCMCTIqvGJnYQZN1zshWrqTweYKCPges
4pJk76kY0bA2GZos7AY3Ix8vwr//Ds1YQ9GWr/hN3ysB5w474npqTRGw/2XB5hJV9/qSk6OhXS1n
8zIVRotJtAJCyCSoNHLiUvyF+TFNLFrgqx6u77oH5hskWTmcEy96movkP2RtNVd9iZ4oPsuYZ3um
AmzkPdvZywWg414ZTBzHwO62ewmNJr2isHuofEAdH1UdyPTE09CWsdQFzlsEA3JGMriP0lcT5I6D
Sb7cwvxFJLssXIoRpDIq0RbHVASctjm6gzF3F9I+EHWrHaBKdqaYGi9nNHOM671NCKsfJRAvpG0i
ECU9PWJ3ECGeAlDS2+ahLb2YpS0Uv1pnnCVC72KavvSSoLaXnBvyj/tWohLfNT7doNT0qI+95VkF
GLscVUVG5tRkkrxgo0W33TAllAq1XupBVKFdIyhePj3pzOiJlkOEH29lobAl1x3j//OKiJJvZ1k8
fkwkNNeeFDhefs7n/hgpp5GdWbSvjzBNIv10hnoUcjxyGsyCTpf6gVQbE3IFqMSwL+QkNE9TOFL2
4PM/vZrTbMCpbc+FN9zFm3dyj15kWhuvuMUBfvpIBlcSu77gzlQpqRWTCJVK4Z6kkZD2jVixVWR9
UjtTtbQx80e3rcYLTFSKKZiJyYYZ3gB5Cwwes3+CB5r652YOqKjPxCLQzMpEpiRLSuae5NrvAwBC
iC/4RY+PmJssmh5XACm4m23je9Y5IEnViWzaTsNPJu/sTGIsHcT8fhjoUJ0VpD/HvEo/bs/Vciuy
iaNbsxU9baC58IvAEu2qY9u6XL/rZjx7/VC3KvCxoSxBSOWNFuqw+aHUUuxG0FP6Ct+5xN+F/FEC
5KE0D2PGYuV3Hqa9tB5962n1MwGVzi+GbipRJYUnQxZdshYWOkqsLaphZq6g176QigEJgTgisMMm
zBU3pra9UwJUwfkYtrgvd2wm3NnEuvSFfEjWAuCCmcHUXJRP4PKz+r3438eBx2aOnaQ+nQze//Oi
Udl8EQZyrZFQpCF0fZIWg+4giA+HkafM11vmtOtYXBY7s9UA6JBpPITEdffiPH8uFOlI7NnH1d4k
Vxp92NGX1JGCOzL7nEexlVwPMVOC5LfWN72ejzORWqkYeJEUa4h1PjfkMkt2BO/eAzxRCW4Ie0FW
BWTWVKOMx8yFYeLNAZir00K6I/fm/H8jaLyDDXY6AP7cqwZZPudAAzCwt+qR6npOsjADGGC35uyo
cSbo5XA1y8NhGj2QJ6HDliygPh9ugVIeWdVL2dCNRq0UJ1FWxtK/HgZKxZgRdlgg6CFo2p6dxX7I
NlC9y2XIQPHpFT1YZpCPBtMzDmBA6PBYboBs08RT0n3vpkC/jBNqWujzGYUW4Mcb2NPHpnsUbWXt
+p4zBELEAngpa2DuIiSP4F6jg9GGidgrcOPfsRfnYODgYvT8ZxH4o9/1QlB/75EgYxt1438H+h1s
jykY8P3rhQe8MosuAiHTBT2ebPcJn9+Sf4nGGdque/Hb3TEluz9uCu+Rp1KlQSLSDxCY5/H5mtOV
sVA6LKK74r1md3mVXuxvzJTxg+KICaSREM5h+Xir4bB6N7YRP1VEuGP8TuKDFe5082btakyayCYg
Dd7PSOWkz/rZOODilDMrCHUO0Vr3gqWbZz3OST+1ugHj4NEgc1qgzLLdtYTJ8YGArpapFAjXNjOq
klyW3yhpQoSqK4N/pDVBx09Gh98xUcTQlPp8U6vvXJ1qvwWe09u05H0zPhHmM3RJGEqXVMRsbFSM
Fp1M2ma6ObD3KHsdNqiQTFyCqFurylrwkepd6oobwqeeHn/sXV0Ec1xjdiZ8djIw/2OecD8f5RB6
ZCrAKwgLOaTugQScMYgsnXuVXpf14A3wv5nMofqOUyr4oH8n+l3yt02ZIaFfdqJhZldDhAdK9r+f
IBW159YB86CozBhvnhhUyP76BZLDdrM9ziLyjTimALsFUTkHAg/h/ya9WvDLUjiD5/JzWuqVX77F
85QDzMj1rNuIQGiVQTldhANTrNS9Wq5hSnaifodTNOciF1II48oe+tFaQ3X7ROT+DS60AILkP3Q/
WF5WjvrueYuDaHCfPV6v/T9puoR8Nu2NWAstB47IXMDIyH/h8rzl3HPH2iK4lfXpUsLZRjuaWD/t
RyKsjfRLZFGo9TaFMsh9+XwUdFHy8159VtHgy69iViDG7ZTWJM3N1SO4/tN6/a7trgC8+nC9dsJ6
/XL+djqFGmrajRwy+uW9e5oayHOrmpwycp5gRcOuRmuu4A4NfMGcjwLXjNRqoFXYzRQ5FKjQ+HJV
u8lDCG0Nk6X2VDgeF/zscYCjb4dB63Gba1Uw/6qnT9KYDoQWyldlKHiQ2COFGMlEkY4cTMvONjL+
NzAt98H1YcB0lydSFRxO1BYfwESQiPF16sY4Z6bf/zRj5PD12k+z3pXy4jJ3jaaI4+1Tl/gt8D3w
imM0IdsdB7wKX7m4/HmPLZZSRvh8TafNy1PhtJcR6F1vdg9uMcT7YgJlp2A0z2m9qpZAUrFJCeP3
u3w3JMqu5Mu62FwqCuqe3kvI7HG6+bkFGHB7qKhqDyKQUW1O8WZA06GlVER7kU74Iei7WdI1He9R
jGTsF7j7q+JDmGMklbaYmkl/O3iR7jiMyGHiogtMSH3lGuQeE9hR1wEAKg+Y0VlQOXSHHfSoZVaU
OGAkpYIUYAO20SftbOzGwC/m0fM8RLquMDKSzM4ksUTgUcP4k3k56B8UZhv2HLnAMG0AtcOOFOgD
CYZ7febpPEIz46lb6khv/KQGlIjpP/HlR4oJ5zDURwuzExhAagsRclIFpc6kap0bxMugI64f7AFv
af2pgML09Ng1nZEsO9TPCsonYylq786fIj9t9pTGjk/PV8R8RWHz9w8WFPwYi71q+2ZOv+a8k5IQ
D7nVtqWbccgzG+SXxfE4IhROCVdLROurIL5YiPjrmze2yJCDIyu+2xAqC4ZaOc9XVWvQNXfpbF90
bNzNh1MrVmH7OnMwK/D07vTmPg37CpLZAZ9HVzs7q8QTp5TaAByyYzfSztAU7ytktqZrpp5hAyAJ
YIICpDG+pcb+G7Wy1Xeh4nPiYPT5qzuy+wgjP94JI+aOPO+l2Uu6gFJCaNwxrCU3SzsgYMReC2Ty
HQ9YdXkl2OkXOrdGmG5wccETFtWa6aL1FO88V5nCMJy4mAiC4BPinoY2P94bSdKQJPz73yNXVZcq
MWQ84bkWHSMbpBjH6ToC/G16abmbqeO9V9TzvNGYnfRaLi1+dF1JIvzyYC1X3wI4lh6yNCIT+rEj
Mlx1tIIligs9MHw/QllAlS2X0qZQrUwBXsGyX5LwjjZZYXpd0z1gSbo82ZdSzyZH+f2Xtjd/OOUT
F2Ne4PqedAeGdUG4SshgJuVLKxte1M+tWjKF49lCvJvFlVCxLD6ChkgTwwRtsAiDMBVP6G5zhplD
XJKS8M52g+vyg8ZXxnn5JGqjhTom6ScmIMnKvMuJ8AEwvKYpqf8+aQGwkjMsijD9TPOj1rAi+o/J
j1g0qbpaK64kcJpLEPd9rNt1MB/VOkTUklHuq74KTv/tAwUU0CaB1b4P8U/dlmMQmA+HKAPDKDIR
uyGk3e5WihY9uXoTgInRIfCVlWVl9fU3dmjfIBOjeDAmxT0UT7IdICECRMgOPlRhiCwHy+lFI0Ox
eChhM1msD8mzsKZM6goyLHSzcNEeLmkMO/5r8kDxg+pJ2/yf+5iBXJDB6DzPIT8/S7AfB+2Zu3Gi
g4lpGJeRDRB1yNXaYA86uhRxUUVPpN8zbPv33aGLJaLJy3x3TAYzfM9EiIibbZO7SHg2Tc9YmEBj
PAd0i60lmZsx1kMo6WPkk25NEZQ2/cfRjWghItUSgKYJ6Qf6HMh3AWTcrrbi6s1betBV23jQzKAS
H2nnauVP82h7ylEELGYlKAtmCGSkw3rNdewCO4ytPK9bEy2Ya1979AlGStmcb7UaN6VADASIMg5r
d5Ek59lt4VcCXfpsq3etmBH30hDgnyaAOgW1uO4ZUGl30FEu9f/rrLtJVhC8DpKCSu915gt5YjPi
HDmGu0P5uF5C7xR42758dgVBrBE0/O3Hnb8jG+Sr6++0nSSL9uxOQbgaMcpToVRk1BJzsO9MxN2G
euXe+zucJpOwMVJIIYPkL6PaUtdZOynET0IkJctmYAVnJ6GF3tf0SeKFeriTI+RwvGuCA78C6rUc
wUqzaRGt+QB6MGOCpwx0kHYdjD/qzEYxTc3KOKFsytBTl2E8gwulU/R1WnFww+gVWVcaiy1Y6QhB
TVrwnuSrm8W4/7nKFtY08fd0kCyvfmxHcLftBTbvl+8TxOAsdmCL3G0dUsmkwYIrgTbLLNBgSran
GUchN4Uf6/gP8i0Q1RrgSUDKFngRHaUTIGRp40Ue93VY0s5bsUE3Viv609ZO5ax9vPsUMmave8YL
5bvCPeLHIvD41T1hHN4+k1ejkTSayW3KrfH7WfUn4bKspa3FdiVbdg8wkxKMU7HnT5q2yULlfAy3
O1ZJKeiD3jGcgXUDZHW4yNKa2hVNEstto98JYPQPgvKpJ154c0yUCasQJLpusvA/fG1I3IlKohH8
ZLJOZjwOEPTlI6QcHUzfuCVZnZD7iLUCL4egUCFFuzTf+4iSWVNo7XC4RNPCpHq6qp7PvP+ZINql
4Ehh2HMUib0MnKv34WkHxs9zTv7cyO2zwu+dBbgLq4UnOXclDPu0MUqtxKFbCV5u5FERtx+7UyU3
kvaBFizmpen0dn/T4Dgx+D9dYt8vXv40PSKlH0tde66vU67kQfmJlofGV4SrzAgheIDbeRDqmHV/
ox16xlVnpveuMf6B7ic+7Q6kxZPTwY1hJuKqnbmewFmUeq82aFOZ6C8nN4ohrz4zB+6yZkSrMPIz
wiTXBUZvT7bFqKzL6JJYbClc3ckdlgU0PwtPp1bh+ZcTjk3yPv/vcZZeNpypJTwB8V7khZBIYAOj
wFycwvTFD5N4c2BD/6tcHC1g6lKTETvCLnoji5iP9gN5V3aoh3d8Gxqmwc0C9T/qe8evlDPsBmtr
gx9DLpr2LHhlKDMQsKo8dD18bH4S+R9sn1g3VLmsPsnTp6kzoVJJYIS2YZ1lq+MNrbm+jJuNokGW
x4Uz3lOgYdigrD9ZV4Lc9gYWGC4Q6wzyiDpQPuf5kXHNO75Rc1BGkFWj1Zxq8TSX/lpn990x5yhx
Va8qostQRC3QYJG3mLYP0HiCwqMD36ntzg2RMp6pz/MNjdi3exEaOsaK4MK7T17quRZYxsOUmVuF
bVj/Al0ZKwOiVKPTxF8KrCRSZDZ0WB2SU+oxMhWdGzfLfjuQGLEnQm7YzgGfNS3fXmfZMnO5/GYE
kLtYlJem936LJle3zzfW5s7y0fwqef8pXSbTXP0LaKd/zhiNJQzJPi6xBPiuC+Iq4fmRdAVanCns
x1p+Ys6BedjadQOvmnVwhTT72TjWCmdvJFU5Uj1fFWtx9FvwiQh2AeOV3Rb3VJBUDmdP+FQTHpdg
4e8dxpx6T8cEl7onAAs5LOx4x0eU8XoTuC2uz0zepWXdefKynmvwNv55rAqa3aM7+EdwUcHwzNC/
I2DYvfC/93vScweD0s+V9pcFR0S/y87j75GZdY5uUlKQesekwZJsjRGgdzFuhdAiF+VJKgHnweyc
kTNl/1Trj78jIgcfqCoKf0MjXfrFoVmBe4lANOztgcJ0Bryk2F2LzlQtMdXdOMgEh+p5KTZ5/8OX
yeoDsuW2m9J2Zk9SBTIUVMXLIOHcD98A+76VrR3H3Tk8j0CLTBkPTGreYx1kqUzud9cQp2rr+lmX
g7bvvhuoezwZSRTwi5cAFrvCUpf4Q0bfkDQU/9QgMVJLwC4848AHjiL67gYTyDcIbj4SW1Y1cyfu
GOUb2BMcMpmPhnMyQ6fYXDkWac6VL+VjEFBdecpLWXpfGqN3TthOealE+pl1Zhe1WXt5462XI3bD
Js6WE7hw5jZelaxdYXytU+Yo2eXr1CbdlrHda1Ph0hZ4S1tTdd0AakjSaf1mUXuEOgodw3Pt5Poz
rW+sRxCXzwS5ND/j2LdxNef+DkznhBzF6uezgatN1kUWMAnzGweUMJShlvY/r4mpNNBx3duJqGOh
1wHo1VF5pLQ/HjACMu/R7O4wNCSOCxkN/2kMydrl5fHQU32xdPRHAsDFgla6klAJcDhPn0/33Gde
jtKgp/6V40xSC9VIoArIM87QuzSxohhO9qvzPja95i6NV8U1aCTPThLt05J4eowb7M6AHwrDgPvr
lkPLBh2PRy15IkPuLMkGTyAgqRcm8cKM6sDfbNdfOvYhcEHmoa2UBeMSTx5XAyKLBqoCyxTEBDzt
utslVKnM4O4vUtxx1dHE8U1F7NLhvMatdvQ5a0kSFppy7zZcttA/0Q8VzNAxOPrTlU9mmUUV3oNo
p8x0G1URTs6fXTX3sbR0iKN/oqm11xj59Bf/aqI2b7GWRZ9R4RGsMHRCOaWzJOKPVvZuNcdDdEbx
Mb06gMzQDrNFwVUfjeuJnVKJvkJvhgNha/6zDZUjXva2yDqCuJecb5GNIKmBShytEE9NgK/vJtS6
FfMPHdEt689rrwwDKFwTQPNqdg7C1wjfnWOiKZeSZ7MUftvb1GlG+QPBc4GleTSRrTA8rp+TzSlN
LTHi9SW3NX+YvOfVNC6249FPQKyvoMlp+KBeE+KAa34QB5VoV723CmerXY2PoeIY2RRZoNl5ixSw
Aoz4mBJExqVVOrKLjBbMODSOL8mykxikyTwScCjaRe1HAmB0qNYRRmQV1kjKesmv/i0+IFL2EM4b
rXtU6wbm8E/AMmYytnPWoe8+PmUFF91pKumj2PohAsSlsRjoTXo4hA7of9yWabPktEhX0p8RdYGC
lgq0n6cHG0gq7T1STFSkJ4KEsFTEo2v22HC2sIVs1js4lkK61pWG1CVtrryPbVpMDIe98rsqYg+c
7N1tn6ukccpGaZAJKPN2zhzAGeHG0HjD2fEvcFMwvVZlvCHcCXitrM3e1ZGuNgaGdSyjERU3s4rI
cs9/UMenOpAM/4odEEsLdB8VMH3sI/NJO6tb5gX0HujfuU92D/hSvy7NED+G7ExUyoPcBkF8Vyqg
p5wECPaxgohCSaHthu6Ndahzwv/ezlb4BaE5KgQ29wFPToUMJ5sh1osyOSjn6oanc8GXITIkzJ6+
5opC27pzRiMZyiFxIG6LK/+fvr8Z34QZYWKm0c2aRmOFZOsJTB/FLvFUOUmrgBR1308nEBnvtei8
kG/45LHtC9ZDxovBnBM54v6mwD8xqjikYZ9YdTrw5OfGKh1AyGCRb1uLtDC7YEJy1rmkmYavUWLE
JMdR5RPKAhseQicI5EERc+KPKf+48pEYqjw+QaZjRS9ChJbAp3/Kd1gaNjdGM44Yq046BHhX8UHn
itkyKydnL1TdLCsBw+Oxr4wkZTqSB5q4M3l8BG59q8xSsf7Ik5dapn3h0CehRL9yXOzBjcE/LsMD
He09PTR/BEnALNZOx6g/yyB2iQqJ+5ceD7eefD6iI5xuxSVsyttUsPBf4zWXtCSGJrVObyc99gMM
9ZbnmyZ/fEdKYXcmuKTnbq6keN3PSdkeRVmT4xXv/GVLUOURfwc0r7mayH/YddE0GGeiCDKO3Grg
5fKZcK3eXs54R4NC5jJnomxJhwr2OemHU5/Ll192lKAkDSVJNe8DpteonTgnSXm+yfhnsvIwhzfk
CniQhOzn7Xc8TxqocwSzLPjhJyIjEBUm6ZvGjkM2PC/Ca72k24MDkbs08HI8tOi6Yy27i2M/1Y0M
QUFfKrlYab/VsMi1WXA9dNCtALBFl49yeP0nc/6KB2KnlPY2mb79BaBamcKNRfwaA7VOLQBtnrNu
rzSWWSLhK4jrr/EOgI68jqbRqu6BBSAxb7VejrRJEwds/ioQa91GEEstAUIEEIaBgWzSfe+6o7KB
BIqlsbQrFhIJvc1LuviG4tS4T9O76p7AAE+DsuQqAOSObVJWI2KRxcQCY1eLFvH35GJNJ4H03LAX
ZAK9sKweixHteBWUHJyNHqQmR3xJBEp2SENXeI9vmx6KZj29mFObdnrPCJ1xiztaYP+Hv0oQlavs
EeioG5n+POiyqM6IZIsFiqrGrQChly/u/hdlnsUM2lDThJGdkFeBJNaFGeIoGb3QlobLJ9dG6bLT
fbMRRWoRxv6i/L5f3N3TW02tcPDHoSBwmrTMttKaoL0y8D38rEzkMfkvkWLcGMbxQnL4i6q8I1PB
luMVo/lGAjv3tm4bqVvnZILQplRfBFgj5tajLrFDux8+bzJ5k1ABKOb2fhZOSaF286f/CVXpqHIC
wLesYsaeEF/awbhCNnE+3Cf6hnQDCP5wXkid7N+fNWl+LgCvph+yTtsF/4crT3s5D9JBNjG5ICJi
gUTl2IEyR89tT7VBo6AEnEFwQnwW7HQg1pOJvTa4Ix5R/2gEUI5xRt9WAYCMETCdmoJA3aiMhu+v
yRNiPydJ+N5h/qpF+HXesdhY75sicx9d/6Ts7jgpceTDKLErUVV7eH5jrrRcKc6gF5RjjEsWaoC3
pV8Xa5/uVuN1x1e6eKI7UTdDcqOSuBESwk8m+N1DktkSV1BJ5ygBlS+CsyGhA9Vox0qfOBp0aO11
a8LCbXTbq+YEyCZ647C34tPeeG3gAeLKmiPOoPvjU4QTwbFcXCkNfFY8/s411abqN7T3hzMTorfP
9zNgejCwT4vcy001gUssgiIsXjMh26TwrZS17SNJzoY+CS8tP4tKDNLfFr0gT3dh2E4C9fmIt3TW
I6AiEpW/9f3MDD4AR/P6dYCjbmSiHgmDWAZwfKeoKkEo6nBHJ30s/wvKLkEcDdm1HapD0XAWrWig
ZCvV4ILhK+CgCHq7URE8WjT0OFx3xPtUhEg+TV0Jl3y3x0k47UNkkcWJg/3Zn9Vs+8JGNN96fMM8
0wUHAyJsttZzKEMG6KwYXcSkyHbAtEwSJ2QUM7UZidOjC5vb8q3mHLDqsG/eSkAOeUGS3at9dMBz
2pUCJ5AGqF0exKqCmfIU1WKWkFSMFt7LkaV5Y+smJfCUcSudbzf8hAyCblVbZQpuVTnDqfNxXsoX
w6cTVNaFoB6XdtXDK5IQ2p7s9a9GH/Cp3dVnFsML2qtgs+T4rPIxF2ZNIqmfbHFD/Qwkv8qfVExD
h97n0BnDPXKLH6aahdHC/J7pTw99w+/2p5KvW1FwzAV1FVrwwadoerSCZ5XosfwDKaXB25l3mrQd
W/L2KGZhrGgymYgwdT4ETAdixlI6jttjLnAxSnlsx2BdkJVBUfcJUpVQVLZHy1bESmkrK6N2rWBL
sFsG+xgDqD5MlEvaVS1e1Y+dsrzi8NDeipafpeEde6nwubxxyT2zeaBa4MFu+2L7pZN+Qbzauq2h
aIu6ZecNjdrxtrJUM99CBzU7czgvJw4TDG5dvqlBd4g8g/YA6gcHW/QoKPz5XWmYk1jlPqHH/ayt
pTew8FO+x68+8RFSUbhSCuSgb/8ues3OF9MYhL6+g9TwYz46tYmtgmPrPihQf4d2EZXE0aN4qWJt
xJPlqD3+MvpA8qizAUh6URdPqsSzxAFxqCR9biH1V+VTAHOQbyW87JjWwN4MEUVUbwsF6N2ydW8p
7ipONzT09Xg6dDCcAkSlu5H6TutupaOJ6PIZuV0kUTMazBxzlWfDCAlG3cMI4MK6Rc2YjqxRDZEs
S2ldlRJjV553AcS9IEKNC5IyUwOwqOJA2tjyGOSBKPvXwvjqeZ3LOOrO4X/Armn3ZHdxERvjJ7UD
sdW+eZbXP2KqMkw/upDaIMiW51bFESLAdgBNem43O90f0IsSs9wlgMKSUrtMe8AwojDfido3cXQZ
hkVkgFTegQ0f5ms7YZ1oGwcZJumCVdZItBAwfKFIngQR61PuyI+ae0KOpyhyO/NT+XgQX3uzPTBi
pP/pp3/IIP0h6XxqzqvfG2py++5BFUfyrbZuFuKTUH0GGFL1L1vaRP6zyUaLKaQK3rfIzPBeSHwf
jinVDm7fhDtjYmq/iGtXQgsRknQxxNf3IZWPsUfj3ZK2Izud2w4QHxO45GUGlZyknCFDxCiXgdGj
xsjWW/VtHeVq7a1DA/mEU8cxPP/k3LVUxDZ+6QDyt/DkjI6f3UfNvzHsxSLng0BrwZjWrwz3MztM
N8Z31mUAqzxArGOjCe/g5OX8FzPOPToJQhSxXaZy3+k9tJJKDPMr4Cz+DBHedG4aNRMk4NnNfWNA
lxh6tG7N1cp9Sp0gT895a6qePPfaGrkOWheBCWaLzw9Vs0UTCMgIdcenmIP+a9vrV2YLGNGZgWEV
dxrdX4TrTjbZEJuTqK7F73+KRIJ5PlKawewfK6wrN7yrEpLtknbtVkemQ2bODTcVJp/FPG8obX3j
m25Qa8nqVFisRJJnzHJ4QK9Z8yrXhXGdZPfVMDDS6o5RPIFVR1dwivLBakDsnRYMCzGexIwrGhqm
B1URIZ4r+d21SDIQPFgU39VW5xXMBF3qnpO9NTzyK9KHgGtA/Ch4prbC6V53CbZl6YJarHWlYz7c
HCgREvf43d5BkunEXWQXsmp67puRhyzb4m1J5O4oMy4rBJssoxqiU5ncdhqUBmbJMJ2GgYpd0lU/
bhTDd6U+Bk0A5oF9FfSh9+IDo7ycJ57XDZWpguBn5W+QURovgFJ3Bw4nHg9rQ71Bky2wrP4Dj0sk
BTQ9DVmivRS1RCTGtv2f7BFt9d9dVtjEFpxm1nJIS70DSC+9v/JdgoRRFF0I0XCx50IBl5oIhjaq
Lj8hBK0KUBDyIVwsR+1NrOx6HlDD3QDwdyiXKlCje6TzG57bepW65ZojVK70mALsDYm4gcm7Tg8x
i755vMgl0SaDkxYYetf6SNIYt+VmLTm1fydQOwe0z3u/q046/GSM+ulhg7/uliLnfJ5liyaw+7nG
WvhQnJWX8RJTDSmG02L30eRXvLxCDYX8rjOYqzeXZe88dC3N2jykWZR3KaKCwJKkfKfdPDNRxy2t
QRp4SzDjtxni3RESJ7C/LCOaXBcYpFXjRKjU4oxYbTtHK1BcCdPUqf8/xKrp5D1wNyr5VsVB1TUI
xaDnxKnTMD/qrVAgfJVM/BLRCORjJRCCOX5yLCzwMuSxvZzOUArbHFG2Nhd3K/CJDqrzm9Pit2ET
mTHQETAWZF+LAE45nYUVkWprT88M1AsZiL/JOea6/4hTthDM73IP4OSzz0rqaLrW2fONL5azUUAN
HCyMAGLpJ7JjofaNfOmYMH1WnA8RjECCDpvb29+tE9x4m8if3PvnPpQl2Tq8q1SRB6JkNUsYJosb
FiGCFPcsGSeIHaz4L1qbAArHVz4fIlx7OxfSrBGQsHAJYVtabDWAQ7UAud17iRlvNzQ63PUcIW07
9OEKOUiwAWhGnaEG1teE1me0xQGYrRnc5PmC3PK+2CHsUwffJkAFv7oo+1ak9WHmsG5qChIjfv7d
5zlxs9KoNArrXLhgQ5/p9u079tFG1zri350VjotUUsuHf5IzN6kIHVzvCks3zXa0wTi7/FbheazY
r7cyanJhLToKSz4H2wxuVNMdjO7EFqAufasnDRLiSTU6czg57CeTVbXaRSMC1XA3ItVc4LxtgKV2
/drF+mfXoIvVt5jObNMPrlD0qmPbx0EMNomsXTORCN2t+fS/L2Jzz9CKun99oM7q/jSV6kjYPboR
iDiKqyQJW+MwGah+81h1wLDXGJrlEyZcVBPeBzyi3isHiaXxJN1gK9wKaBi25N5ZjeMZBkzokKkD
/gm0gPf4O3ZK6x6dYIPEhmuGdpTZrFDuH/UbO7ejrrENwKxuzftH5wO86b3n8NKBsx0zgxjYbte6
/wppFjixuZqhPUZXKp+Z951Ki1BSdV+IKcIegwMAxqlHs6qpfeNVu/5icvPCpnkBW7QyqUdLbyi0
r4F61HubpUCNzD8i3m3Q5Sdc5J4nIbUzKAFXvM1R/x8jaKX/Kb6qHIdJyti3gdGrxZ9YK8fBmucW
6KqA/YZXg6PP/uLhO3n3ZWxve//blHptAFktgGXOKTQD368ejaysjiZsDDgVkViB0Bo7zndp6u1p
GzOROlE1C1fMg6hI8JmXsmo7y/Zj0I9OioWzJwQsfG5Huy8ayR21X0m1f71BIWNRwu3DmIrJ8t8c
mlmg8b91NqvixjYOoOnilm7d4w3ff8cOkiCzRTXX1nsWExMfE7T+ezZ8W96/XLm9agwqdhYiXvxG
NqSdPnG8HJc5eer9UCXAkWJUGHzSu+taOMH/UoApm3APWTFVs65p+goH2gKPA66/D1vNVc83AT73
IUemzxo05HunbYEojt+ktJi9cIs1K36gl10ylYAPkyO/etT4E0g6PTv50OmpvbYzNQg8sAuKL9+C
9pIM0Zqe0WbDOvHB+w95oTlyIrycoZa/YX+6gq1H6Bf64TwHYF9qZnPLgUj0F+u60KmH5sKnE46W
JDKpKyanxXxOhIKC1XmV+oJSjpA49yci2i+vOB6EbCEZxPaPzxfgyXQi/M54xP4x5LfHf6y7MEFx
anp5IGo+lGDJxxPLnYhQN1QrNlWB3MUBopp7Nw28GW+djqxcDm8Nu46/maHNT5zOXvmAy83ceW6h
l+izbEKkaKW1ErfcbGkqdah7+uBvoGSVpRFy9McasiNCeXHHgOQ0LYkH0AO3x+ZuE5T64jCZJ2a3
H3CHOEZ9nyE7aBt0+N8A6MVlCS/XLyJ2KNFw5mxhWGylUyyaF1RMw/bixfz1AgdN7xkO4okE0IhW
tJFgbpq+mc9rKU3//wGVcTaATIYaRNEkRRUDxWWsDnBWGnK9YSkoq2wzR5Wtl4C8QIJqDpd/ScRI
dW0+uXMB27uibXKJkBcBjm49aJam3eD9UKvEp+zjcsfs0RKOdaJSQ+cFh22oVCn9XrOg2X5nnEHk
IfofJOizWoNIuDYs0Ysidw960QSdDVIxi+cCv7VEjf359LpCdew91jkVzxRq9G48an4flEzU1NQO
Aw0qJls7+UyXrLuvqz6+opUdBN19PMYBck1Zy2F870T+X1A/OBRwkDzX1WAS+mm3lZWTUNn5vVYZ
6wL9J2+B8VWykCOOx3BcBXoqesP7+y3676sSm0BpwbV/QSpFjgmOWoGY9DR9Tt/0/yypwV7T9sPx
WGn7H+4TFNwrUDSIu2Oaw17vq9hXoFXcO6XK+ZXW0f/Jc/Xs4lkuwC2E9eUtBOe3RrRKuofmr87v
RNMM2rDH8ciw5XJvofA+JqONBkAm1sFeLcxbzljXEqdgSGe+3fcjEPEnl5tQ3r8rPGso6DPra3nB
JP8vGAy3XpW2EM5hfcZ2CvLab53caVAZ1aultPEWRlqps7apLK4Q2Ub/wC/tEcnfIPbb7kwQSd0K
0q3kcnF+1bVx1p0UTfpDjTo1NsiJ40v7Q9sUFZyyXjEwQrbvM03luPQeBeSjc0nNHy/i+iRTq/CS
CCR1bmSDcVwnPA4Xt3z6IvOJzZhiJK0pnRrddrugeB8gvmgOiqJDZqeme1rQAe6EfbaQZF8IzD8J
zE50yD1gGBRsrQe2ROXAS2RHSZlDhhFwiE+d0Eg4g0d5fQNMUcF36zlwhHNK6o6E6xwxq7g9xtHL
scYZcEmLi2gcPdWtcS7cvYREwF3DH9R8GfMAL2DSTEBnjv0TdRgYTJYr5J2+HueIZ4hDq1JV+Y7e
2WctaIQgUoPB5gx5Lt/e/WbRI9eFMc3FbG0hKRxMd8xG7b0z/xhAo2a8mHoMiJOl8LduPQOKAhnr
LwJ5Rq3rauCFT+g57BBROKuBB8jULlUeKfLBul3jwkzGKr4FmuTNPT4OuLClAHFG8KALbl2+vZ5P
VasEiuZtM3Hg2OWN6A9i1twgiia2q6yHuPR0SVPeLotaIv8tJnBvBItV+2Z1KD1T0DJalKN0BShb
qpf+oMqeWvxekFdUprttA6QT0EQi8rfoUtK+uzqSS7oJX9F/TYXDLBB4kWN84tN/7S1Ij5mMhV24
sdef3SXGZMZXekCJAXGWN8SdJZLIPAb9IoSNUoPZBGVzG8yBzqpqnTrr2hzfPtkFnURHTZa4rWpG
fw7xZg/b4/BIK0xkVFNUwX3UjVuponuHV4lZgrT2yKdyC1LxiN6adbhvVLqXHx4TIdtfuU3xy47n
LOAcVaEHV4EocaWzeLn913Hw3LTwWf/LVt5c/DMMnf8gLshWaHLwQ+Zp1kVkA0lqFxw6FZzfGCkp
7cYHK9wChCecn67KwcBkPAz6gNFog1yjCv59Nvb1JQAQPCxQ5VYYnNMY+BIhAOAhEHJinjq9d2Uh
X//C9IwNY5zRswGIT45Ut7iGMOS5NMaAK62jfKWEYOTHnPycedzHqYi4XIqG50W9eRtsi1CPu2kU
+jwSR3khMxQ7cP7RLn69bFV10MkWaH3RKo3BWiB7bW3yXGLm5oT4NE0JA5KezbZy+L3GKf2FwsxY
JSxvzSHTwDjTswtH2nwGmZHLmz3vahv+0AI98ogZYqXRXYjEd822gHmsZYyS+csBQd93MzT2foRd
Q7JEEYKUcIdPt/cszDrfoEsD1KN56ghguBpnDyddiwDxB+5hNWznihAudnth5vLwVSLhqu27Daqu
sgV/BlfbY17wzJE9w0sMlQ5ax05+iprW7/b23ZPp82QJsZuJM+oIa/u0lxvS/Ajf+VLS2RwFrOb8
3GO5mVHfNRFp495mAQX6/FDyR+66PYBve6h5OwtDnGzzKcOVVJNEA9gLk052mwSX+TOikSSPisSO
Pv8Mw74uOQH+6bg6xpVsjWqEzplmUHF1y5EQ9NzaIqo3e38IPhlv5AOBnXF9SYxj3FgEpl6Ajz78
4CEvx+4Eg+P2GKdMSo3sbJXvONg4c6Zxfd4e6qr9upBgKNsaxzzdhfmbjIb3zyUWiuCkHEzwuADA
XnEo0xBKAhMAGQpCIPdFXUziW+dnYRlc6rZcTA5GLPFr+2ULup2H19a4Ps2ltwIooI7/QUTv2eKe
UwVj4UyNxoh9E8H7uLL/Hm/7aWatvp5AjMN8ekjXef+Y1jSiT7vx9h4hhsv5NNtMex344fO9dcvI
KLROsnqyW5fNtkQp9TJIG6wEp7V45qID0+HalRn5kd3VIT/OiBw1aWOHU4bMXYm0w+fsefyO7aj4
cuMFfqmjAJLSTuAfxEgfZzFl0Pla6ixeGlGxDu/RTR6CWK/aGwws37x2yJLoE/4cR8fZ3KwkFagc
E5W7VBypkzeiuwxgnpbvZFmbIb+iJ7uhTzbapTF20xalCBJdXTivr531inqdFuZISNr/qr9W8JWD
g73C9v9JGzK+HQXmZhCWU6FPSMzk0+4fBsMz2XE1QfTG4g1w/P9wy4p86eu3QJL6az3ji7lAEEzZ
+eRH1Ge+JbMhXcjNEqoL7+q0MM3jOeTmY5ckzvTFXOL5+M9aXg7CVon9C5e+JRsFVg/mqzfCtzDZ
szeFpbh+7MbMPzuyjMENrmbtn7f1DpTYNsEjOD0oyABHkXc0Dz6+7QjvHuXXkCdP2/cug/7Y4Lj5
6NcGtu7+Yoa6di3/DmRC2g83gYTH5peJID4oDXcHt8B8eKIjWLVLSOUV1Rdxmcqb0KBC5UQCNGAG
fTeXtu5A5mYcYqVjZx8Z3Qaz0NRyh9brlVNU4MPHcjlgmiIWY4C50bsVnWfXXKgGrjV/wra81ThP
3Y+7/wB5uMwm84zmPzBdr/t3KPF5e1a73z3nwUtKzKkNrooXOUrDf6fxLdn53DnB++2DMdMrdgYS
6ncEowwk1b6aINEtfNzZsh0FWi1ye7kNaJPijD1902eVuR57tndq5HzjLi9Gvq2XCuGl3BA0+g9t
S1XtldKFAa9XHcCZtYIB0k/1d9j2Ma44zzKJcvim7l1kP+S+Lxc7XBX+0dLMhufkOrtDj45VOzxV
wfmEJKvFSHXEyHt+ebJgHnjyqih2J7mQwNORsreAFFThHHLQKQQbE/c+2YEI9yZk1eAdpgYJPIb9
wqmY4viGiebkzqm5Q2JTqhL+pCgi7c5kNHLtBkm3Mqkk3FlhNZpEKxYKowuFRXR/Ua3TDXohLJxs
MyjNdu/E06j2LvO0RCTwBE/HVXV3m+kJxPdANA9+GRymHcC6UgysfCXUOsrb59i57cvvTSKoLIDl
E5eKcLT1/TVf88bNr3EUPvWqPr8DLuVvroJAXQP/GOwIOdDj8HWdC9iwbDDLdfd4Z9uyueNtnk7M
3fSQxvddrlaU7zZT1gOpznTt9kMQ6eKwlQEcZnw0HhPwydc5oL1jdE9RqluF2GwIkNhGx3lygUlH
DsjZM96b3lMYifT/Bgs+22JfVBdnYHQjkeO+0vdX4Zsmc6lIFNvYGDB5Z4PuCcpnepYAMAOgTXBs
ggJheaz5oUnj9WHdGxKbrn6TP3SpBVL6Qc0qpWoxon2dBfWANC3bZIuBiQyPOsX2mKtYTMoyLe0G
GDuXecNnkTY1RVw6gBLUm7w3/NSMNoAR8VBbLkNseA1e4Tv3GEGSSEji6frG/pp/shHd8mH79P1D
LXPZnUgykqkRugt5TKojltKFhPh8R9lltm7D6FIvGRPzLXtTTro5dWbeffA++oRxTLM5FVuCz5+p
5sHHzQWqf35D0Xzj/BrcbhtByT+/yEWbxbfG/grXBWq/a6Zoe3eH3dH6UXMwHpSk/csZ3CwSgh4m
st/5KAnjqoalQeXyW34zFcbF2Wcsh+2Du1kxbOP9xuLvB18SawfZkUJI2Ece4uptLJ/cX0v5cewD
2vT5A5ZgovDoK7x5eIxPpmVWQChUp8mDhcTtHYt5YqGEEQPe2ooU/hjGrPE++cz66IlHD3vtVxg9
xMpojg2GnPk6uHhe0E4FNGtvwNCcfVwyJgsLskGLK5BLmG1R9yD8Y7gwzALj9DoWAUzjXOsYJhgh
XVTvMye9SeUlSiimh0/Z9du+a5Sg/usj5hgBW2+WS0c5j/TTUrCRA7HFTJslR37a6AkH+r14jWtg
pgJq1AyRHLujZZ8OTxkC/QCKEMwJvXWQyV+CkPLshRlt5f7WI71bEEPPrvu9eKY188e4dBf4Uo/X
eyoxjvSQTvJstGPXh3veEEJzluyzFaqJUY/2yU8aIP2lj2sn5c43RoHIGPKrvKJ2WL/jj0h+Ku89
COn45SBpNY5dTpvXHs0dZAhs9LMXw4ZpH0iKG8IA7jULAEgxH+Vl+azSaC6W9yWJhNZo1bIjPkPK
MQjh0jsfnU3S5PlftP/cTm693uxHuhKBIQUHbCBPc1qOYKFFj5FSWkcbtXWUmvlDk2Lm20sZXj+8
lFhBtH0aeNu6o4tDDkJqjp3HSu/wtmYVOgyVv6CqNIxr+czZ8QsW28AC7mXZU01i9QnH8ukntQpL
jLdzOoQ+oY6nKxjq0z+RcnQMHbxAURNPSCESLaXAcqKJvEtxB/O927cDe21LW3bdzX/9fvbsTDJ9
0iNQeRPxZRAmKI6f8HMISqMJT/MJF1lCcgLB0VXsrsj8Z15AjiKXu2VbkaYYjVHj6gMMzcQUTNCu
sr6vixf+rJU/Ztz7aNKzISX8QgtO492yo2GSnFC9RIgox8/cPfUO626jEIy6U9e88De/lyQIhNmY
ewwPH3kdNBZWdw4711giKnQslhSpXD8RY2Jfz7MLsba3XbEODq7L5OyWMzui68i+dHM3GN5OCvAm
lyqZ3LpZp/Gx/mgTVv+Qa3Vbg+siPkhQLVwdx0EVV3YOEMOQETwH4WAV2EhdBhyoQrXw2QopHEQu
g+2wGSx3FqYDPZtgiriQU/2VOopmXrGej+VflXM3t12kPCQh7kcn/+Pajxj9SS2c8jRbNL3lRv9h
5Sg6Wz1a/jyIwUNmzbv+3jGnlmd9hsFNVZ/WmVNHNTFMayVhYk/zabOexZkTlLoB+HknV3zhzS4+
cGsnizCKEsGWIdRy8/Gu/0sW/Nz6drtymeEZGBkf88XF8SzaPoOpEiMdlzC7aMHSge8YI/AdYy73
IBIvh3UMG+lsfZ20JHYU2vy/vqawkGdll2YTrEVoGtOpRyzwy3gr+Ox500c3FTr7EKb9XWJ7DWon
WTZMl/UFebSJoGFY7QYB1nqsybjUbzh4wPbpznxb9G9dq7CIfkDQKsMWe+30zmbajVKVR/R5Fhdt
GcBK3gH5g8NlFBmUR6LWQBgnfAx/wBdUbC8paxrYLFKXmnMBXRPncEUMtEygZjLQnGQmfVH3BWNB
Y6NvO+ZHQkgWZupxhX9f3W2rbEHvfLqOzWq9+cCQAl9vVPHG5IS0zZKVZikt4i1LOdzm1KFWsx98
M0Tk+aH6TYwrZfiDFQGNbgn4FszrGZoxH9cjAs4SI/4qsRU/lO89Tzho4ChttQiykTyPR+YBqJ00
EiHKU30gfHLhgWF+Cm/908/yv5iZS3f8Sa/UyjqkXMXdEHzoRBfhot9sl8Vlzcu2D+1cyrJ4TDMo
O1eflFN6iPJ8cRLyQjVQsLQDuevKMqvrq0DIzjcbPNm5s1jFghDQ1YY39xsaW8euhhQcr4e/hkQS
LiElIRh3py6j3Fz61/VAlGGSyPxdXWhhP6cpayYtS5GPjENSAX+CsrZWDuDluKDvEwK9XtPjE/yK
Xqk4D6jyOMhzEXCULfXvn4Uq01lsE5icz3ib0NFAwFMhOpjDCrqTL0P8dm4I/qEjG/RWOoDZ9esy
mbT0DWE+6aVPD6B9IIJCueU3FIloM3+WBPrl/TKViqWGqA0CmRi9emOiHKSApHkRgUU1PYS30Hhw
LoZBiwUTowTn/pF7dLBSPIQhYQ39jFr/iIfRcBWFrkMvL/751lvxDxuz1ATYIQQVAu40IRyfu9A/
jHUW28dgGLGbS8/vxGT8K4fiYJIxuxvtC8CuXFgYWVFIfgHgrA8ojGBA3JT4sEXS+wBg4gJT1srJ
DSnI44y7RZcr8ZgNUHsThhz6PHGsytZn/Q+1VkAfV+DVUmNyruP+bQU9DtVjZfAmJmWELA5ULlJD
ucEeP2wt3X1dWbkXdpS/qbEfetT3TSeME+Y3YJQltnPWi8OXbDGPEtgdn9NRTXZdqfaxwhtQY8qs
qpeoINnb7ikcogbrfcwoifMJ0v5cpkR7FT6iVul+reGVDd7w6qoEaE+EEg/zcY6lI+sNE1xI54sg
VorawswfrAnk45Pab5ZDuPgLSyVowW0F9nZAJxQjG/nqB2Sj0j6E6C1l7YZR2tOIh2HE7Huctyoh
zQNiGt+qPzO5Xn1i5D+epj85ebwHWqnhcdvyk6n1fGh6NGWf8vtwWTjGnrM0GTbH4u2FyHw76udc
eemZ5J67jzxZPRMqNsMwpDrxpLw7SHmeATREYCiNXlBKwmVI6GpOG2j7+km1OBY6xsw8rIqiEwmq
+Ppa2au5FgC3KDlq9XolHwbMFKwuAgwSX2Seok4fKH8jSZOPsVb7RZkRsPWXLxc5cYOgciS9mD/H
2c5EOsXK4J5qKmuU/YM8l5i5SrmjXl+TBSlFIABuWKsYdR4GrN0pqyGKp9AH/BdTXGLdgX6OJXEy
WndQGomj/W9Z/iqDYxWHrhVnoBqPa/zyFeBzKR8QKpTAX8lokLt7/w9NT7Zpos1NHRqoystTNHBu
y+U20F2qfP4YP7mIDx5MHVZRM/XyszbbhAtBF6j6hWLGyVt+WAtwEFNmMA2zNYEG1lkp48cH9t2v
Am9A1PMzPNmpLH1amT81FDIXO70YC8nLvdk64WEVZB9p3gxSZDTyisabubv2SbhNE9FORRzaowoq
G9IFNZiWqaKyRS0yX5Ke53EXNIhqBdGmLRAKiWVmn5pytQHH99eRCB0i7L1qVx0qHnjMYPmjhknw
VALBVzUVWpv9DYBWw0nAlRFx387t93qh26TTeHfF0/fym93WPm54CVINxNpnnmHtKcC7c1aXmgtS
yb6fGamdzobx+EVUfUvXBq/M0Yc/w2iC9j9kWdepqr2z6WlFvT570nLaJ1YEun4YrcmtGJpQPB5Y
yzvhTV2Irsk6VIrQMHgDRPwCDLNft+dprMiOjaDywtCZaRRjN7ztQTEo/HNPwCd9bVGjpYiduh/O
TY/ot031+gc1DOYm3eOkPtVPPtm35ifT3i2KbtgfYnv7uTKIOp5oI/MaTmENBdo7jl6RGsOBFIaw
srEH4BO7PtEhh75Jg/+MHBEQuwtLEoPJXuGVxtH7V8idi259l5UVZr76LEm87Wkj+Ifz8fHglrJe
OXH07spxg3IoWd9O5lyat3eY62EWOTuCFiXTjNo4VIojyvKr6XS/GnoteoiCnYLjSp7ccxDisCTN
jq2CkffqWgnLSNJiS6mCnK3q296+wD5zNw372q/cV57ZOJfd46cwQQ79H09a7uj6pJVZmtrOVysT
qncUAT79fOdwrNPhoP/Daf+dPjQKXT5T5+RArjiG0dsMzoGf35XiQrUXMOonDGUtnM36XLa3JGNW
K8wNyjSnRaptgMf4B33dWWYICjaVZBRlFNQeYlt3C2HRGuvO6l/uVAobv/ps7hqBUZKjk3hXfYVX
zV9jemQom8D2PyKvzfFEYbKFIjFJNnIFfYJ2HoJ1U+JZIHYrrcTAP93ZLd2OqY9x3QHI+9A/n2+s
5YxWBBja6Si9vqLCLFV58EpmjZfYOQdQUwVW052qrRJ9NHqJ09EvN8M7ehBbqFFbc9vNJhFcagKc
Fj3DFnTGCIXpoIxvhyGdUgHN1jYo2fhSjREJccCWKiUSsSdckhBzBD+I0M3FYjWagwqjdonxuRG0
fQcpqXtUnVjFr4sReeRyq4yAp3O5FmEDNIibniVTXMkqb+yeosKUZG3rGL6kPZ4uJRY+xzeMsaXt
OcpC5td8Q2o0SKsGPsrz292BdKhfIKplTTivTQgFFSfd4OCsN1Yx3QV3pJUfFu/P1CCIaV1POr2v
D6sR7o2FadJAXnv6FL9x/b/3vgntsSptPDzrZxlmLi3S3sjbO6ORMvfP4iu3CC2G1RYWecDdU9Vl
DGFpPYPiJHS+pqV+LKtB2amo0syigAjFfUxvXQP3aCuUtl2lsK04pXZ2GOWzZ8YJ1c1SSlTucuBl
qhRLHT2bXmvs9NaIKxa2aTE3KBRzewXzlvj9vD7i/cHD0SMFSFVWGRR3AL4lnlnyFNFxYE03KuIq
by6HcKyoBtYOmSdlxwFvN6dAF7XzihNuDwaGZwZf/NYlUGA0/C4LHdpGv40erVhraYN4txdO3bs/
TxYvqtZD2csEuAC3eY3BO2+kSpqOzt6wOq0WpQrZtmuuHpDZm5UUBkiAjx0vHuUFsk3JSkQNBjiG
73cYTWwEoUnXm15dDdMUgYctT2DFTUZm0G2ovhe1T9kBaYf2Js46NQOo7lk/j5zSACLhpReTYdN8
NVYUsVuVQIrjQhtwxz2wJyowNT6kNA/M29KpAuU/68QsBgXkjcEp3+jiuJj2oQMteRQXcIieznhk
mjXJ3QcKByM8anLhBEAQLhkToQBBEPKpUWzqm/rTT45UhgxjABohlfqKCoAi/V7+d++Ub5I7QdUD
uOo+zUAKLMp5sZNZUK4RtYxKVmU90nYV9uezQfKrqz9HaJ01uM0n22nzkIcUd2vN5Vm/BA5w7nSd
vl+AbX0L64BlGpqyqelXqYijkdJPcdVUg3rtGmWGIwW/Qpylet0KPzR+WVB57ekgSp9gUm6xupPz
dgjWC1aIrtxJoEg65YrC73MtisbYE+S5e5+zOS9BASxUad6cmDf0mMgN9pPpSmts53Qs8rU9vUZw
UoEJ60CvmIk9e3J5acLaky450JTI4xem0XoU4X9MNCfzIt+itNoNfDWiRgZuaWUwQT0ME4qIRz5g
pIniNBzl9bQfz6NoToY46NApFbDompB0zKJM6jkMrZiH5ce7vIP71E3uZkS8+z3kynxl4KdrafSd
kIbixMRttpT9+oeSZNjgRkfsQjErqUURWqEw/u6EB/GzRaujSz4sy6AGWW4OffedP8n+2juClsS1
KmC7mroJh9Xto7ZO3NjITnZddc60lV8GedNFPXtt5KWDGFKB4mO4xc0Lta8mSlx821eEQP1Gojc7
v5efMsZPdYLpkBC15VjREW3he/f/aWbWk9tzjdYWNpJxNKnS9pvGVYvF/0psuTj7GlV2w60euj8S
ysCKmUWd/KMJY+dzdI1WDKhigUQuKzbwCxEJ+iRxdAxIcjTixA9qkBKh8tD92sTIvs0AkACbTQMI
G4Hnt02ubE5M5qOgncaS4SmV3gzofAsyboz5afRQhmQTs5mmOMnH4CwJWjplS4wmyGhRE5JWVvAx
yXJApYKWg2JT2txVeAvl38ohUkcZn4LeqxKjstnXncqP5N5tpkJEu9FTW/pCyKj2JcJL5BLV3BRQ
wNhJRdZ+9kHmfdMK6y5kXc2uBr/1TBRzuA+Q2T4hUDm3IwJU2CxXYd4L3C+tt+aRR9KdtEu+D4gP
wfOu1BEOqMaZ1Uifnml4RRWFoIpohF1PaHKPY/wgqaFSZqcJtHLUUTcEO+IL09vDEKzWMFYtwHEj
p1ifX+LETxNOlk31BYecq+xJwl3q2yfZW/GDOPTY1WfOtWoUcbOz9FK8zZKjwt9dEF2q12ot9dZo
PhBKiTPMzldtrvGXvVgupFZAGX4GWLjllxxH4ua/hWAYVyb4inIqP9DpMp2F6uepeB+cYdGb1Ebf
1QE5gZB7kLNLJURZdU3pcNIq3wU93dpid1jpEgat1ReP3CSgMlkWGXLyqlIkG3W1pYHIsk7ysCgG
RhOmzxZ3X0duRj+Z+klmlysuPUh+KvB9WZ4q9l1RHXhSLKYuIjoPcj4IFgJZsimUb65F/wqmMlA0
gsB6Q6O9oFqXTqP71ImeatO7kVFAF0ikmysH3j2so9XMfqXZz+7SUnyoDc5hrJUuIC366e6Hpewc
ZFZnRkUOT9/3sZ35PLEy3ykNPjPQ0dLhyLYBlpB1gU/2KsIwMGTzFrMrrllufKvVxfudJt5g+pq/
iDCCrArNeFakcohESbCW24t5sShHx1i4s3losklc1qYKOtCNJJjuNvzLWQh4ecNM2ll1o0MeJvtD
K0LBJm/KaFjqcZqOcmnibNCm/tgWMPOexSzYDVZiYEpUbRZeq7QieQoQxqKT1jBQRw8YxwggahJB
i+PgNN4BVelUUakl3bzYLrunTFAhC8KKHVolsdhdIB5TFSfKNkGhauWJO/8oaPghI/Go1ht4+NEh
pKqZ7doJ0lEDTHfksQI2eYphO135pGB9Zv1KB6CV04t1AMrSYiRwW7VLVq/Cap15fWBpNFryJa/6
cQwTNLVfZhIv92EbWHPEEKnN/O/4X08AoKVBAx2kG90EQZuXRLb4JCUrKI2YQJWk2Wwh2TZn843L
rXTZ/ZhU+WS9lcejAOnytQgIaNOA69+qoOc04JB2TYucKf0m9WcCDvZc9/EVCQ9gLCIQOH3oYnPu
64VnC5baoePBX508VsfMSOiaz2Md1aJwpIrHIj6pJmJOziXpE7uBjHJIJr3GvdNzsj8YMycd73SX
IUqsFK85Bm/vYP5/XShsyAKS6VMH6LM0LLEB47iP+cv1sd5r/fPKw/e9it9TW7jBvKrjX/PYLCo+
cRroNbhHG43HbSkKWAMpmMZ3YRlOEo+R5RVYXpB3e874cgomPu8xIfMM7Gqm5bp8vPKtZrrzafQk
9k9rTtJsV44zR1Ww022ZKXnWPoNtxZQhdAtU8fgVSG+jyL57Ml7YY4U7Woxi0decVYNNII2re6+I
woNoeqqH9C50LSZH8g1MqSyhAGg6Fdf50/gdmKRLN8ZvOTx9a8kLBQ+sxfviK/9Mstn42kLXDkQe
KPKvGMPX8rVSFlybVHi6wswlpHQLUGpcoGRy0eELvp6l4NJOe9WY48EGSl+Dr39/x7DY+W+DugbH
awfQOP3bxymaj5YjU0eJYSkU4XVYyazPeQAFb+G7ToKhmj31iZAFSelPrWW+4R1myMUWiMFsdwQ4
cIzz1hr2do8/VzCiOW8d0DWIRRqWKDkhjs6ndLS6K/19q+Zc5pZot7oH/Yow/a/aWmaCbuN8KsXM
BVpYoYyywdmEmUgHxuqN4tREjTyWA+Ncy6MqZn5MWs/9AvXFGUFHmP1xPSxEZKqDcdrs+p/pTOfv
MtqU7PrbdAsGMrnyG4OtO2odpUetS4Pt+NPTWi3TBUGIRpXZjPui7G8FYcTRPGJl+QXHw/G6LwQb
3cJHf+LX5ulhZRojsY5lZxwusBSKxjVX1toA/GwnkBG/wBcFD5hA3bd/p1bUUk9+6cTVWzjjrbH0
BwxqQZKNK6JMPbk44C/57CDhx38ZH2PkraWzLubgmNWWy6zdbpK0Kc7a0sjWgY85sQ7HfyA2lYOT
1WVpQGzuZIx1G6orZ6MrTCMS05XSyZwhlsMVUlCSxEkeeaKblEPY1xKEuHlwxC46XOmnI7J58Yo2
gbMHxmu7T6U9hjAjQ9X1JV/VjN4OJ/5DLHWbsl64uanWEtYwp4VCGULtfZ+o4ueCmDmIObrVnN9t
h0QFEzFe2X8SO/R4VKZYwdyhauSSXpPP1P09spEVJUCJJ3wnUdFmMBA1CHg+wRG2gqCmwYfKQqQy
d03Lvl0To6111HmJLNi08HD7WCsa0iLVMxAhYfQ3L1Hf/kv9gGugtF+hESl1LoaJpDRgqMA2X+Kz
XVQaWFdt/vFsIYZHBnYXRSpwGSSD5pJnddh87X8eUiGo8E0z5TosGciNTslaG+pA5Qz3cZAvKdXw
3iEP/VeD3Z7onKxqLJ5HiKC1qnm6pFSrng66pQDU2tlvblEngHVsufBnQ3jYCwzkiwcHkcELQlcu
ZY2BKDMob4JiDcb4eLGav36xzxE9bfQGR6IX4QVatRVluHlqXLTGbBEDqBqCRviNuYNUwYUcpW0Q
BccNwyatUILa4RnwIKDnbi9b+vFFOpR1MDWSwn1eNSk99eKSSOHdNSQPFPdzCpkQVSCogFb7ZYLp
nwwn0RwfbiCLgK/jpnuSGWlqS1J75b0b6B6prO0wbseBPnRawbwKSoP0YBolw5e9qbTy/sx5mnjx
WJTk4Mal60UP6lLkg+Ccmv7/n/zWGD2tQ90YhKsA0DHQfzWWvmcIQGRm/2xAAPVVfYDZu+lcv7tN
9AqnedemyoFXTKKUnto623FIxixtMnvZS3d3GW5Qztm3CQoclbSLfslS0bG5GfRguWIlMrimZRCi
BqfYn4vpIvwsKeqv/cdzDFBDv0NTtvj/+GCIEUhuL1W1oJl+i423x+xXcUUMvLXv7hZzPTYUV5gV
oHM4w3M84x3Ymc1Q73SvlMOwvy6dp12pGaFuWBOMYXPsToNkljMx8B/11q/K/goDwV0TeHCMIBG+
MYea/S4ELhLkH2wTcxz6Vdm+NKpv66rIX1gKNWXEd+bMUE3VLboIGmXG8rgVcH1jE/cDobNMoYlo
593zVFA99tl0Pfns4Tub4leHHrIu5txFJnsD6swo4yfEroq1s4zriafpTNKhh5otzCH8zzVamgI/
VSDQ6co/zP4yjs4Fij8RK0WG8wLkFnNq0gPTHLJKAOmkjv3R9El5J2lZS50op1g4qPVzO19S/+11
I8ep9KLyfi4qFwnLFnf2g2bkZVltoFrYQtBI0AGGpq5h9xg4E9UVXfXHHvRazL7NvlUvtHTNPSwj
b6wjwu0UP0N0E5wpaiOI4pXTN73vpIqpFAOKt5mBHmIYh3gqE3z83N/yDCkA3xHM9DzsYHy+gL8P
iXcu6fzI0/jwwq+kPb//nc0q9YMF+nX+sw1srqTPNRGCLFYBDSPLy6aqbwrQY5AuOFc/eLg7bq/d
ASnlATZc+0w37wdM0oWH/vUiN+W/uhfMy2fQOFaCJxYneMzKR/aT8A8SDTw99hhrYtkvm4Hj58te
E0S8sCq6Np3H/44YLPHa3EHBwKc8aNCbMTj1TxwfJxG93v/uN7D1y6TtHByoGaSA6RJn7ZRdphy8
MSGlLV88RYE+ekqbrHlZPDa50am7UQ5lkofASm5E8y9uDgDNTII47PEwIRBsL7W6aTC9sDivccZ0
V/t942a8wEFCNoABmjmMOVWz6KS0lbRiujaZUWc+LAlQEHyRTqjTwgOOH6ABSB5KQ4uB8eezJmuQ
0tN4QoVCP6RzrUtc7Kv/tzlnOvRejUS7OSZQEVcyTz3dks4HFXbCR7Q9ddAfd2wzL9y4NsuwaOHE
Kxl55eqk+BCmYYlj9q4NYDX7rJYXUM89DB6NH2WPjZMiOM4+yBKvHQfqrMy/Ese/kb98/aX8/z+j
QhtFuhkIOtYhridxqw8QtYquFe0U2dHFOSBN77uPQjXv77fSSxf2lyphWjSx+aj9TB0hrgW68PdC
qEylxQp5mzP5viVqLNlQMwgxzBwNP+VlmGSOV02nhBqJRIDiWf73aAVIZqFOMbSmqWg2rsumvjo9
p3H6wNiF4T/tFk7MlLRV9YUWbwlVxhxG9aboate4/If8PcmPU1QH9OOmpqYLACAL44W/j+vNptKj
p//zWb4dptraqOWqSTXRHbjdL/GZPJaBWhhI5lMAAERrReDnVDtgYtmO8KKFcWdGBTktXVBlgTrA
jvnDzQL8Ma8E/estjQm4d+MSbuBJg+0qxPEEoCOQwAyF4F0ZHfuzIOt3KpQPkymx6Y7I5BrJLTBI
SYpBPHC4AwFuZOl+SeET4bbaADdlZVbcVTSjxDIfHgoCPhB4BRdjOLk9g4iVeDmZiCqDBti+AyXO
wuTFqSGiPdHYEtt77YxHwNtVDUcLzFrCm2YdLM8OKU5/REaTl1XCt+PLC1HVE1nw8kWo4wLwQhPC
Hnt+md3+tdybWfGGQ39lYjExWB0s02fj88AaJXrqpk1znmhUOTzm2gpOAvEO55BnkOIBiYK/worr
YItdWvqcveauFbPJdERDqSVCVS1X/9eKkpkUaSdyrmYujq5clCFMgA8We/f13uiUh9MEJd0HQEI3
A5/zb0MMu/SA8NT8hs4xyd+oa5fpM35avXo0seDR4p+naerKNT9krbAqI5uxRz0rQnF6YcTqa/CZ
8BdydhlK/NYWOZ2lQiinOS+cYLr3tot+j7aE9ny6Jh/b/U/kh7LS8A2WSpNPS+loZPU0KkFzsesN
BiGuv1Hx2TdFHVf812DBWq4jrU2T4Bvdn215tItitCUKTUvOzhntSEY+ZrApFHWTYDAJbJP0axem
JKRiSn2X/aOSXa7mU7rXzyN99nbSKVf1kUyJcv0V5KVubnlI+UDHkB18p6KSYUgukWal7NqvP1cp
R0c4f6ycwhpwCfMLaEwQhaivOhc9D0SDiXi+MDv6CqSuBQ1NFizqBc4icpem7j4QHQqAJqN+WEcK
chtuiLrxIkeBqBzGWqH53r17BGG+uENcyJFRL/b73eHskrNZQZ7e9OE1/vry0xEZLOHx54pw/hul
PgG8HC1VFL9K2ivf7d/bIBbzvVkHfspOHK3S9qlSHjqCooKyyErpL3c4PMayLxa28fBNouYa6XuM
rYzZsv5aPboHNaSatjESv4KFO1zszCgW9fI104OhvVWlyPybwSgrHbMWNoALcRGjY+vXWMV1chcQ
0Y/sIIX9/01ELVAVwOSxwy1LHjmgR15dQveQEgUOzGmbHYb8fxcniWlzbO+iuCGKRqqE+P2e9l5B
/kB4AFMoYDSDZR7h6PeIF+UdVyZ+Ij1+HEcW5bMRLNq+agX1LvUxW0n/IE/siRZ68ln3yM1e+rmw
tDqoaN2rf0WQLYgnQZ0NqMu9leUMIwu3V5OlsCQ9e4okZeZ1TidY73Uzi+nZJYc6n33jQrpkNs/N
oICmQI4Wif+ncYX3k5sYQX2jCWksvva5aGt9PJVABEtfoHdARh3ml/g+nCt/aFlxEfswbXRMN9OP
ArmSyE8rDd4wqZSv1jWgQSxJQex9FpCJfZ6+uuitQ+YwmznKx5ai7cfr1sRKoU8KvcxQrzWgBXcQ
g3pM4yZ9EFTW5s0Kpg8qhEAYB7fYoCBV/JivC8Im8kUzF0EYoRVJHkGQSWGdgqKG78Js7y7NVDf7
+2Jj8iYgXmUVshKOTGkf0MYNJL29dweEtMkIQkepj0swrnpE2dSoNGa5bRM95ue3GIicbshkiIMn
IVigQw0du6JIY8G8cE2U/oqHkDNkAOkBhhXb0BMvn+fVr88Aw7KtfMtPGPm2rFicJjOSqauOsfHV
xoM8bpfWJ/jLF+F1rsO92vw4fzxW7n68AVk9b8WH7r7mhfCZmtMKtUHLl0Hf9E+1ufnKCXPdZh99
7wADYMMyAlCKwiN58C02Nye9mTAOxMku9Xuq5NYycTxDq1dws4/ewofFdKMdvqns0vKCFfNogQn9
CHnDv+9A43hQN4gBTSS6PBKqyLeR8S3g7ZdsVSRSAYf/y0uE+1xxmnu2g056JNO2H2+pqwS0fkUg
`protect end_protected

