

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DoylSncttFMA3kx042gUfpgfS9f7wYF6CWxJheifm9U5oZE55E7a0/gn13EV1/Vn6tAoLpUpkm/0
hmdlNetDYA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nsjL1A4AfS+U1MlmYTovZuA+LXs5hJP3SunimigW7xSFqc+G1o1qnLbV4BnmOncmqUv9X6mR1dbm
lvuLbnkHJpdv3qype+E/DkwUU+uuHlSP7/5qiYqLK0/kXVQ9CK4RGY/33UuCkCUXhFP+4VquDr0Q
ctFJ3ADjSF9u4KfkLp8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e8PwETDI60MBXnrgCDSTetYRVktLV/+TTSXZzS5MByZtHEX2iao5JK/khM4FDpq/v0uNsNW0rhjn
1dIPd1mlQZEDfzGgZ7rgxmjzboNMUH8CMdtSuB8lFy7Tjd1hDXqhliwc0PhPBGYBs/YEff98J5pB
EaQ7x9e3Dm3lUX43BX76qZ9cgUsaVwP5tX42M7Z1CZ11+5f7kvoiSco/DGzJuhCbDcHoQ2NjrZeO
tRQwYWFDIi7vBls1ETe/q8cjQLCZThAhSFjjijV74aEYat0gpNy4Hxz/UN0rUMO/XCqC2k8lo74U
XZlHepR+ABhyrwVFzKEwcRDXuuh6ogUCrZ1mMA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YvHkp5oDmh1yxPKtyY+bCFF9nl00iIDnF4JnEfzCQKeCjt2Tok2cPb5/9L9T+H/cQ1x5qpJZSOJk
cf36KzabCPbu4/9VIe9vwmzzbE9Ndy2Ov8q4+HYXDGn/u3gDUJZcIYEnVlc3E6se6bxCrEZNyRYc
iuoolgurhXiPk/HMhX4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XZ/Rjfda7p8W+LhE3BcXwsLXrN7RfTJezMmvWQf9ZKb6JJ7gmlPk8WkUFEwjbu79kr2SMWbEP0wO
UouQmHkylGRubs4N/1VfavspwJxzO5pggGGBLKHkmxqVxAWJEQ3Kp5uoaJSKWxqKIRLzeGXsW4p5
F/e0YM5v9fK6K2B07V0FxCP6WuqrungKJmSTj1Ji3gWd+VJATYp+hkh4HPUA/aDTgCzwwIaJ6QWy
QvHMQKHrEHbRztbzfLMH3RPC4Jl5v7PMeYTnCv8UcX2dwujd4zD00VIt1jMD19vjN2WZ7U8Tl83Q
sPvYlUbNQVTnqIBf7mqYAoAlbAFXbg0t5zqPAg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
0DGIAPIwonnLwA2kz+MAiCkEdLxCnaRGK7sWXtvZtAb87Oar4X3RabROdq3h9fn4xHHIrkxDGMS5
qPeGw9HaM10lbSeRgfPEKHg8olWGxzh2u1aSYVjyYPcAqAKU1LGvcy/3AkohQCvD/+Gy+dKc1wtm
arm1h+V0Mbj7xvScwfYOEJji/kmoL3cVu3WNndlgcRVlA2nmb89nNPAZhDvEVzWntHoc9lARh3iT
W6YAt8PKFre4nIFWE5Dbp/RzlO2pqouFx2RAy1/nFjYeixEqIlqC8a1VUfLzhf4stX+XEMndgpqN
M+FH56Avelvj+jrF3eamwI6/Br1RiTauu71i0i2zOXl2ogZJlh1AKLAJLh2nFLqsx+Ykj+PWu26E
IALkbKMkkPhonf2+oFqQha/nqUACkejUZ0tB0ftLcbaGqaNDRuBWABSXYrhFuRYoUyBnyFoHAdA5
c+xHxYJly1DU4Pv7x4Smqy9tUvKAn1n1dZ2mVNi3pRFdssK16WigVclMYejElY8weLXlMZgVfEXo
c5Xb8NUmAiLmdeeg62ZFeKn60nMoxqrGvpnU2BUGFlsMMXJLs/V58A9/uox1NJ9+UwDZBtBakpNE
/SNqWCtwhjLt6XGgO6gH8pDo0RPKZ0t8GXPEDpG9GRwW94CEkvFlMVxT5jOR9UmleSxSjogweG2j
BVlMC0QY2F8oDAES9jqtrJtsv9FeqguuGMrK8wmVn3RlyeXQalQBc7mRoiTCBL8LkH4GpYA8bvVo
dNPuAPcnepohl04LjEtuI9x6R1tO/ZkT4iKcnMOXFaAHNhKnn4QU3kskA1W5NVVuCTQkF4OPbaHb
vMlrPddZIWKWfsmuGsfJB6yoLWv6AcOFZSU+Dv3ySYOn3+S2Vt0cJY5SOPmJPhTM2ROANa58UJwP
w5bFYzpLhKNMLd4psdPY6/0/1TOEwdTkLcDPGZC8crrjO+wJjcx5CxXPE/L0iJDa+l9lbXSQu5gy
H0Xvc0XuatFnAGgRBYVwOhPvrqjw4vasyRe4qiGm6uk+PfS16UMm3tzu+MlfWGTPYP3L3Mxml1Sl
+g2itIaQGAL0kamfNochQZi3F4fcGNJqOGrvWF4EIkFyh8GfTCBXazpkRW8vyx+spQGm+PY8DyI+
xpaDESw8PyzFeczHxHyQcXs+UD3IaiQSkOPz9tHLGA7Y8z79lnUrpAxGBULApUwuYC/PRfwuBcz/
6lbtEg0rp+Ld3TTQpaLB3HmmAg7ev+AZRRCYC6p29AgRORD0kI2Q6A4rSNFFkqfWA4Q7keVFkhjE
nAdmeq8CncuGApIq4Yu4oPjVACpTbYOOrocA9p7/dt3YvEK5lWKIr4AZUmkRpLXSbxa9VLzYpGUr
+V9uqlooVC/BngEHnJLg2keeedZ50Mqn8rVSyCoLnuOZJLwpsgIafkmwN5aJZZfxwxdav1A7kXzM
wXqTl/wctFVecU96xGnxS7msaG3C7H0InacTBiCSWCgvic1GebBc2e68RFrzRc3rjSUjrk/ecKl3
WEhJ2JOloYfanIji58nVHLOxJVqb8dzxaHhuZC7ssI87b8fpjyoij/KTpKrxgCQehC8vLKzgPl/f
JPpoeEvmL66ZLN/Tf4sQP5FAY4/5wnSGMBTQqQbYm8WZBbTWkiZw9rCW01FNRu5/yRBeoytdBs0T
1SeI/OnBrg/IUYg0lYOMX4MHTsbitOmk6cflw7fb7+jyhLcZks2NeA+/k0SRofkVfESDcFsXiZu4
sNyl4TV6ZMEUsdxHuBuNylud6z3GIjJVRQprZUnwE7o18hi2lIterOKPH5VNoZVXK3DF1+k18lY+
r7gkn9r3oFeb2ORXXUw5qwlD+M/7FXygJWslTRo2wtxKCSCo161SmyNyikPzmsIhxwkhhIcg7JrI
bY3ilmKAAAVrVtfX9EReMOXQ3fSwThLMWUcqJaBalbcyNiIxD+cDGoSbRir7G2aEBmwBwY/w2T+W
+5TIkZ2jefN9vrBV1SfYKhcK4jxdwcB4NeeDAX+dyU7W+jpUVP8qEdcRgK8vmBYRnF3INSuL7YzG
qWHepwN9ViZy+s85rxSmb+/OncUwHq3tZ3QCGKYQVuxyBgY9cs3FvN33bgb7plj4xbu5l6x7MMDO
lsu0gqK17AcQiy4rqeYg5/AB2u/DefE2OlwVRFUaL+srNRlGusbL4Ku5kquHcMfxOl/0w0ONYErC
MWw5SmVse02LmF5rDiglQ7RdGGQbXxCoUBUV7Q3kIDMoAppRGNBbFXijqZNQUYQYn0k8UeT+4cV4
Wi2Jh3uy0tWGiVmWqE91HHfkH66hj7hfTd3ZiGpuho0g5qFTNXbUulOSHn7DIF3UOCL0n3ZOLoYS
zAl94eEdMGsvhfAN9NHFpBHpvdp26EuIwq3vaQTcj6njazFpV+3fbqlwPXCOLNfmZ1jvpz1JnyDR
6PwxH5ZjxCZUmpOajHHmlARSTS2pQtTGQFYux32D2gPRiyY4h6hAPYuy8GSBzsDQYHGjrUIFyFr+
NI+OS4vwsrZKxPy6Wre8EcN6NkLMecjW3nZziN2JutdQ/Jj8gJjub2DK0t4flqs31hkM87VUSx2v
pbj05wYtq46sGAARLHzwV+qZzzIyhgP3Wbuh0c8iaMMyoim+4u5Ta++IPqXsniS/4SgqidN/urNM
nHMCShnlAwbOf5A0tIrmRT43C6Py+gMV0ERd8NpBUE+ALAJ6aUWaDQwk1eNR7xEO1A16rNiVzHp1
S2qtEwvmK1wrruQBZ2TLa4XQOFoGucy+FoFAWRa6aJVcufvS6RK55ZD/GEXSQbsxatz++mbAFrTX
DxjHZU6nqmzCNR1P6Z+M5O1JI1sLcd4rXPGokyCim9+aeJ5zcaFhvSP/eL2naHI5rshv0wj/ZuM2
cpxOFiKrR/ivIdt3KftKgzb2JVbjSoo5ZffRhxPDkq8T/GL+17sbZglgCF9/pGbOhzCbTteR2YiU
JAlJQL1wOTuQ8yl+kBo4KoHnIXCU+xr9xiwfgjEGIrTcqaodbany2bgyJU84MK68lqMMZ7zGTTqF
4lkIt23IUFnJd1bEJAfId1L7RksQQXb6R+QefJhEMuHJSR2cdIqHA0ekXBzTJrlbxTCe4MO3eu5/
h/xzLfqfkFzJCTXBR2OuTohfYscuS76SCsbbdZpC8LGEhHUAhacEIb+mEbBMTWvAEvqhoGsp10m6
4N/SGThWh8f+Sd5/IUDwCu/thYF6SxRzqYoWAacSzkQVlg+vRXC6GT/9wlzebfZ1HB+79qEta+pj
EDEz1ZnjjHPWtiNPlu5o1aHWQ4faFvGB0H3hwS51BLXVyo2WDf4dEuygXYWzib+yzStmlsiOkWSh
eO+D8MKbCoSC3XK6bYTGhoSiz5SIAuGLmCIH5P4jmE0Owy2TyvhB/cL09KHOgu2mvADieHN3XEXj
JXYotMqh0dSwH16A6liDJ81BKFaoBZe3zFpqpqxlXwH2JWdIBj7epAl2t7YtT+e8fnV3plb/+aZt
rizkNFDDmfSr17++mVTxZdVXQXRzqAg4MPKLwN0TdXJ0uVaLusCzvKMM/KnUbiPnCz7PgExwc6Fa
rz4rGXzRPR0YbXDYu+QVFcNvSb2euurtlS3IUKnR5QrJ7L7buQgKV1NVYBM4W3akEd22Lf1BwGnI
5fIGPeaxlEEWx/uj2bcUGptaBSW2N12VMm8hl6MRxbgc7Qg99CIxRUBqrEcpHNgj6qsQ7KOIf2Tr
d2BNlq9EAB9Fl3UGM3BwqDMZUjMhNvbqbKYGioRlyifsnsP7ewtEIkVkBPuec8qhQGHjKyzN7r2S
3iBGcuG2yBSDjmhKTgqTVWLTrOhKi/nLlxtJVa4DuPL6h6IFye8yRm4ShbzvXOPoDx64IR5MpIGA
Np/RWbPKQtcK43pjHpj1WtEvAjV2OSuKgL8RBwIr4XUeY2rKZBLid7j05cOefTEXbZWiw26Fy9vj
O/FbyB4ezgwGmvYT+gq/hGsfRXF7Ip3cIHb783QRaBXUoumZ19wP68stIOcwWbSkWn18NBwEN+mb
M58Kr6zmISXIDg45o9vhSYHwB/bsL8Vsg8xL2kqNu0TRpXq4C8Ci4mGObmeeRXjtdBclrM0Pehvz
BFO6XdXBfk6ySzsmqUpC0/j6cWmK1jkH+k7GMM3U4xK+94oCWAGZ6JKshIJ77+kJSTViD/Z0/Lgk
VhXirqIxbVIeBQE+d4mRHQ0XjGDvLxMVrLfqxFylrUIxq+acT3TKPhpTaCJE9dx/b6zNTrSGDQgG
7lSP1/AGL7hHqvhTYcnjgdVnGGpJ3YP1V+P4rsrJ3UNaF7i0Ma5cPWhqTdKn6qagUy37JSgOOTZh
JKch2/SS5WYsGSuhwudp2AkUqbZvrCkEX9wi49+KUaABMQxQ1jQ3ySNRfEKvbLMyhbdDkgc8tPPJ
r3hkQ2/iegXrjHVYiAPfcD67MMClZ2kEO7N94e1gLCy3xzMXDRE76JoF9wUcvpIQzH4BjIi95ELv
2ChpIZtKEcl2FBLCL808Wbzc3DXt+sM1qfMqnVrMsG0Oc2DyKxuppNfT98eZ6gBWU0Or+7qe5bdy
38s81DCcD2O0D3Bo9ybe5EeOXtX4qx3kEveFG9WItqu2G/slyeNbrefrXFjoCYiVOXsltHFuzcrw
pMPx6HRCiSJW4VaFb8sPS6GGkVQBjyiILcDGjHwxgaJGPs4JgQrv8jefKamCc0Hd+vLn/TrM1kBj
n55nlevoCaNJQFTLxk7kRxbnm/Tph5fcVbhKajbqGTbLN7xRbiYstY+v3DWmpBP+4Ta+0F9PoRgH
/oq2LBqhW/wV4i+e8GhW3kWeW537ZMO+Jd9NRrqDybIBaLdLPbqHAkBEvGHapYRTnunJDKM1sUgR
DSwoQj9PZS2uROr09SVxDX/8629eYTXXlhx1JfWW2EVDCxfg1QNGZy7L7WeJxAy7SKJRl5QrArrU
ZNSURxtzUmuqAUJaqQhotiazbaDJCdeghMefe6k6b6bNUkPnL2DDXvVRq0a17v2VWYaJ521dx071
UmkfSJxZlrAN+lJKD0XVhiZW/c3HGo2BZfupIs40RdW+m0pUBdH92ZqKcz/GiNp5qWEGHLPX5OD5
kQZq3E0/lwgMmowXFXAm4rkmPCW072aOyi4WgwN/f6AlF447VfjpOxD+v6BUTd06N4pf6NCjBUHF
HRcweONj8fdLghrjSvPUoj3ItYmLhTaO2qaDzQL7WvhtYstfUP0UGP+3reCFgntZeD5YCmSBn3e8
j+g+G9tc4uIoTDhILQCqrj8FUHzPKQ5JT4Vcnonkkm2Un1qyiyoGOabRFA3gFrE/hqrlfYzanZ1d
5ea/VaU/xtokrtee7aHLVW2t6YVqoOy3h0IDSqFzC8LnekTb1ltoX2WaWRJidrntksHGfhbdXA3t
Lool/TGWlD8SnA/9Rlm5TNR7oNU716muR6VS/wuofjOOo4nqzlJy2MUSV+SNKdy1eAY9vjXhgVUI
uCGX8cMoPligQjMC8J8RH2SQi3t5UYfopx96CpuLG51EF+x7DDVnHR13QuQqRg7BZJAiSWPOESyx
UG3DUxyx9EsQik2Pc/GXTerpQnDxZbDJ6t+5Byxocc/LfYlA1Y86Z6cjWmWnlfPIT4VGG1g5PuOg
ghvBAqZX3+LP1pUXDnbbCAmm4Go5V0Q2UWnw++3owJZn8g2D+lJEotaGPqm2SSTcAeR0gQFbTehq
h7DQjgldsGsZoIMAg+zmnNaHleUw67HFRiGmnyhqb/MDSvBE2fjuTRNEfFLXdk6CuiHlxB8qt4mk
8OqHz/0LUyr59N9HjH8CKkxv68eN2l2byZxe0c6h7G4OwecwSIrkykCQuh+tqfi8H7+xab1EOEw3
JHk3Uko9wfQ2RlV+4cwjPj2MnaZU71r+Jlo27p0NibBX6D2u1me4t3AQAb69lPHlRMes9ie11WQT
DxGiN7hi4HE7Xe6BODCOqW5np9a5UWDYKFXETgKblJOToOnn5Cxe5kUnNWItqB8Ag3nmO+lZtLog
/nn6LWWuOIWGB65BGrTBo71XJvRJzfaPttMsoe9JwKD1naebCyQBK9jJ/Xbohjgbsi/gzik2sPYK
jmV0b6nIpiaOCtYkd76uo3HsJzom8TTz99bJ53jC8qORjpaRWVWfyXDVz3aE8/59/JFEs2PXX5YW
sw23sNXAasrpkRAGiBM+sU/OkaSTYeAorn8EhcwEecz6XD11B3x2cZ6TlsAvCm6Midvf6CHEpfuv
PSwBpIQqHps6troMgreJs/xQv2Wlw8/Al6QOm1WUOeCl185B2wh/E6DB7qN+0mJliU8j5pzWjvL9
VDzehrUISFMMXNCsENWIu3ZcrM2ef7sQEsFo4LoUd2AHCfGdIMOIiFl1D2bvpcSMAoDCQ0NJaWRo
fE3TgYAantyWs+HhLJE/O8R8N2p+jgnLu1/C9/n4LHJSCIkQ4PwcHYoJxgjM32agVwuOYqrPbOcX
W/lUI3BHv6/m33zbVy1a5zliD3TwNi3f0Fd76MlU9VqTPxlpAuBZyrFaArTqnHSZ7p7exXvLrGww
PAJUNOfC1jEyEmxvsBeNQWUoiiAYp+vfFmbPszVrUul9D5xdvJ2kMXVWPp3zDZABBHanFquh/gLl
VTNAp6znkDkRmojgny/SzZ4UNRvbqIg+NjvGWatrCYiO8KTR53k+zlDBRfgYOotPPqz/a5u7jb8k
JjfiQtmRx/wKzplJN8KNu5tI/FHnft3f8vYmLLASS8ess3mPeId4BWrJVhR0SXyXQEqiVc892WIA
OR9V0iTPzt3ewfhRmA/yPklIghATgOzLuzAbTWXEiT6kcWGIrxeGObjKLw0H6+Losn536Kcnkbh6
tEVxCQIaSmdloGD/MC1eH2V2YQcLZ3/BIm2u9fJnIr58+cxhyYlRpYQvBVwtes9dTQoXcFgFqP2B
uCEwxS1RD/BZ63OSxYtyA7PxpWTZOLOWLxrnW0hFyHSVsjJF5sdbhbrXL0b0zYRIlLt1eEq6rDbI
yihnkeMTSg4nqADfa1DpDcWpuGL3/SdmDhTHt+QNtMrYtATslPNqQpfi19gL7Nnd5uDsO2O5IWKQ
4JKbiJmG4Ohs3/hXXDPEU+jBFqY3FNMg04fOHuRsIomhkZJlUtQ6crdBWLCzpXNT08w/D7bJ7ZAr
+8ZixSNPbYYhOf3pkFFyH7vtR5H7uuslLQZ4tUj4+IT1YmJyEdzysK8kT1ZqcE/yQiHO7/9txpJP
5INc+/rLXRp/VdbicdqA3UNN1fU+jaCF/ps6q80jr4FkUMtGTfrtIYMvQn3kf25d5mVGNh3cWOEJ
aV9+kdERFNFR9LratnABIo7akLw0J+pIZ3yYwqw+PlzYtFx/YncrVKicMo+QxhSQbzm6Dvs2ub4b
yHV/S1a5JIfi2gC7YXn2/VYRkwPpvM/S/byJlZA3HQWFa3Nl/hEHCukm2ceZ6aQC/jBEkdvlN+AY
Cuf2kJB7LW1dwpeOcVnxQbU/GMbO6oeQhM5R8UKr5ukgW2rEdfZoEQIfsiT94CZWLZjPJCHe/NHy
EA1vjctNFPssY6mKARI/48GI3HP1zamDt5rww5s297rwJAtzH3NwNBY5uFSqFrqYB1XhsvagHqlh
3HhQRL/haau9Px5aewKcITST/EnLd1+cPxGS6tU6vZ6jEpgnAkEr4JSAe0rMJbggV19yrrHEQdqg
GqEsGrtdpXoPyuaZNiBYHvKyNStrrVJEaBjV6KRJ15cq5jtNaYmPS7a1zSpRPofIoXStDeP9Cb8R
JMLnWes7YUAC17C2Y/0qHjr5zeW1ve2rqoNnAYaonK7VNiPUS69zl0lLDLTwS+yFpaaPHsq5Uk4i
V97reciI6haVc6yHS05H4ko5IUNWt0Y1FuyqbEswFxUFOL1cfSSqs6QJuIxAB1370jiHm+nfXkGs
5HpQ/NXTi39pXBG1+qFEHgwt45V8ezdXB79OO1obRYsCibT1gLsko9ps0hGunhrTWumPVxkLncxR
nHEbLg2xsgDGQHpuuIg0fet3MR61aZ6V7SpGZc/YKbxH9910ejS5oS5luDAzEmLSnMv+zNRYLhKB
3aSq1+FnUYEzZnf2quyYzrd55iDvNev2QHNd9iqf7V6MC2iM9nJBhA0AJA4/9U8wXBH0P8tNLHaq
96phOabjzDYNry2VFDtUG4FDwfRydvvEY8M2e3VTMuUfIui/S3O5WpKcb02HWIFQphBIBw1iiRzZ
8kkfz3SlxuZfoi6/CCba76qsuvLPIjXT/KtjU/RVJRIjiBx0lE+4Da3hD2b9lob1C+MWSDl8UcaI
mZiLie9W1sLy9QKQ/6mWuLUTaO9sgBLi14sP5O8yRDvklRkHB/nnXckpcvrflhD9MP2Z5OF+D8p2
Qyhul6NZAKmbAKO5oDzWGaY8Azjtglq2zXKQd2VZS0INHu3qfHuOzrp5jWLmTr7wtJKXVU5E6pyj
9cWdMKAFL/tilXto9TpO5tUI/cMSwNSpCzZk8gFDQudl+3LKhpC5H7gM5xdClCW5oOcsGXvyLplh
bcBHe4O94IFOWfnCKX9Ec1HSluDsLGW6OlE4TjuhoXN/PH+GZlxzSuMZs//Liz6R/O+rykNyAbLc
OIsiSqtFNJN5SPM5UvV64Ziz2/tcyLCGj6oXE8vJ6vjLlm8cr8/r8QyKo0l6zWbGyM/uWU++CDwy
beSQ8QoQDmO2xmtJaau2+olJ0l+yjnEUXDullK/ByIjx1gwqHTeCN3FyLgip+v/zGX+WkGenZz7s
reIOqRIlGtxfNdvCebclCY1m2WPIW8pbLxU2gkpZ4ENdjKMvw90UPXNpVEHb61HaLWb/+dT9nYNG
6d1BmpsGmMcXnwCcbwndLSLiafheETS2bb339jIYQd12beIjNPlunZbYCchXC2DcXD5W3XXxNqKr
L9HP5Y8qK39axl3RCwKrllqWcaOrWGSD+vv3pTmoi5ba69rR35igfkZT+qg4k6Huz7fox7TDQsEk
XIiunb0jKPkR/THCwHkeW5Iqff97MKdM+X9GTlw0pByYAV/YLVZZlg6EqG57eAhNJeLZXX4PE7NN
JXlpTxsPPVY+HlLldByZbfIROxu9vQIu3b+JzzVSu9/QtJgPmIlndg2KqPnbCmLRneWSH+BwHHCt
sFbZBRoAzHl9kncUG3AvtEIKKhdcLVJ62Smjrie7SYtxV+wPpfZkR8mPtYDXBt1evnoV/O8e8XX+
gQqM1PTFCJ5XwgDzTn5CZ0NJp7krBt2JtYcWT/xpX7+OOzpmzXAASaJXa5hU0UApvwo9SRYLoZGk
RUdPeJqoxfGMGaOCcHNnQ5F0+4IjoJoRRAQKxngZ/jD5D8Tu7QgeR+34deP+mTyA5Wktio2GLSlO
dJpL6R/SHbLwomjGGeQRl2005MxZzGXqFq7cJo4FJTNd2wBQ7ayciLWJaAqo97mTUwFTpiccrXID
5g0kfEhRdBJns1XUJjBIO2tpJ4gY/oXW4bKMS3kkIzrE+1w7RdmMpl1J4f8tQPoDFi0DToI/jf0m
y5pHHKEWM9zxatqWGS51b4uuf1Y/izPtAsebEP58frYgFNT9wShtzHAM78i3nWZNFq4HjZ44Susv
yX4JUwOErkGTkZ+0C1Fxeo4runXjanQEoMVudzTGpHec7QAEJfyDyvZYCVGEHGW0wZuwep72my2e
fWITNb1kapI+ogsVKbkhEFY2Tx9HIexQYg7ipbWhZhv1ZdEVXlc/4Zu3uN+9usVpxHQh1VsKSX1/
Y99UwF0Jp0ZJKE/lNn41eC3H/8Y/j/YD68+lDmh8/EGArllv+HCNBYpbDUzvAVuzR9Xqc0ArgAkJ
WOHcVeW5I/7E6ZyxCbGz4mhHNR0YdDe431zu1mlIDaW03UhgwVRWtFAdnrC7CYQHk84TJJ3CsFYp
Dvfk9/MIN32OtijgP2mIqKQb+bRWg1hJ+r2Wq24Iz249Kv+cD5/gFmHocUAfZUMk1KA6R4qLtEQS
yNjgJo5um3dDWr5D6z2gYdnYZ0CMgiUN6bLDodXw7YZ5B0o9Bm+WVjVgvTa6HIPIofWs75llAnJy
Qi+lSbrA0ywof2UXjEk+TyFn/rXxvZ/IfFlDk2KS42lS+vYo/v3DIp1///opT3MyCkP/PSvu4C2C
paIfJrwdLr7ltxJruRiaak7TlYTHLgukWFST+Q1Y4VUdpZARqRIc1YRbMoJw6h96txqcstrMbQW3
1ufTCkVuE1MdVjhPpTmv0/XelX8e4zFuvU36iQ2aYU7n8z+ynXrf08NrcJV11q6JKdO3GVY/+xwm
5xgDYT0tNGDPOhfJx9PpxCpadl333RcY79JHiydMjje3uKpDC+DzGZn9kJu9b5gCUsZIPTfcucXP
21q3y4RVapfs9KtbBi6virhVc4PlYe9qm4tAMHVnduSIOuxmyz4vdq72prv45t6lRZKWvSWLP80n
bS6cDPA24sqQ2CUfuhRO5oVULqtbKwD3ea2ZarFL3W7GFNcJLqC19C5+A09oy3xpZJRFAD+h34oa
HA+ynJqwi8uZpgc1O+WvBB0B9AhryMNhnx1bbSx5lp9ne4AOOPyIMy0fBy0JROx3NK4DRnFYmlQo
UBFs5MMeNLFUXDBu1a1u8RCY4bv+n/nToZYr0O2dffsO5Z+CYUBbvfqGKwFlikxCL3gQP9uvae+p
pX8raJNKFlIcaH/wR0+9UwSSXcMRxT5lN6goU5QQWyk9LGor3dF9QKU3Tr1YGiIwbVpO/07XGpgD
mMqRzZem8U2E1KS5VnH9TOo9aFQONiYroPwsa273VHGkJCsLvMRtsmxh5+nsswrCcKiwffRx9hN9
PGkxcorEf2PwdYXRtdmsuAMO/q/sjinRRXI1pHJ2aPYNi+WKiHMUMDvpIyLUrE70GadlfTeGP0ZX
ooK/4Oj9rm+OB6Rj5Ge4CxbXHvNOWG/13dNaewC15Wzm/nTzOoTPVHBc11ZMjLdp2LPrTiIxyy9m
ixInT1ZFIYRMgYnKur+iP+CwDPGhL8zVL5Eyx8y2/eb4n1mXXR0WwRMnZ0IzwyRNA/rJrJypsm2I
6M5fhS6F+BinyJyRfteJ5IYodSZU6zpQT1yi3Kb/PV50GrkIHYEYgbA1GLH7zXPjrc11DrlnvDqr
vad3CsrT36P2xBcWuzev/R6XiYoYFc7ReF7U5l9llGAGTo+2VfyQ+SDA+6qopahz6QSZ5gjvPr4i
PwJMWs8QJE1nykbJynqhzDEHPuts9N31LM+IGL7NrrIyrk7KRHhFyVY8902FrJKK4ZPXbM53LMkq
1eYi78B6qkQ36CCPPo4cT6v9WrF0iNdlSGNknljLtF2PHC/ydZbn10AK4ucGfV2lJ6OJc90cR7Qt
dgwIERPr7GDfzgCVQgZwPqDcIeuODV8bo1gVjVMdobGkj7r5HP1lJeI2OLyd1jXW6j1QXGQg3V3s
c+Aqkjx0UO7hqHaSrTrgAemF5hfQKE2qXPYJHUZitR/6OLlhs+iZ6NBN72Dny5z2fnj77i0Kb85N
33Ci2SUTJc1lG/wgU1EwEi3feRRa09Z0tAb1WDsAe5049+Nux775ZB9Zuc69EOJ7j4TsZRNybzL6
APLLeFFlyZf+/aCzwqdtX9HxzPnS9lSTTSqXIffP5HkB6uuW94UnGtLsDLRrK5/YlXfrmzHNIkbc
W6fubmWnVpMuykzM6PKkjtAJw1tfnJ8196sNUWfmK5G16F7V4KZdm8HbDqTHErhQTwzFw4y3EdxF
QcFbnWPpuZCSON9AxkkOJdtyXH39yDfiDOEhGZpBsVrcporKbgSBIPws5yKK8uW1dkx7EyyYm0X0
jZMmX3e7xaWFOWK2wYHLLdjGz4LI6I8koGSM1ig1hNTp1RME7Kert9DQIPRTQjSRQn4vGQ6IoGYg
QPmIyANg0fsCb7vRn15XNGR1XLwGUojM37UeT4tCYq/pWuVkYBL9B05eW8ptdFu9LCZghPNu9CTH
A3qinuQ1ZDx5s9CFXAq+ZfjwR17xC7BEDmSqghIqn9lMoqWZ2DmFY8gwuHAES/DL0Btag2sHYdEI
M9YzfPXJ4bYtClv4SIXWsQZu+YknXqyBjVPCSirae3FdDm5tWauXY/E8M/8w4kLSJLX1Mn4ftIh2
IbjeZHFgpnKELpZjfrTgDJeRPBkg/SOEuvJhkHpGBWWTaBD+iJD6DjAlJ3LyjpWBA6uq7MnZ/Y94
SPftJOKUrpFrdE98+3PTS3p4/keLGC5aXGnU1+fpLJrzeHUkChNYfBiz9TJKWgBvtizVTDWmcia8
WhGGLRyFB1aI4f6uLJhng8vdoiblAieZ4y3/q9Sat/oZxvi59WI596nHpS8/2Bi2hNchAa/9o2rN
DQ0A6jYE7D7gNr7QxV5nX8uZdCjbVesdngKSQjUVcmXpPeztfLTxSRoUvxMTWezswT9KQ1YnXTHD
rmL0ZrAztjGqGSFtRhFSp9pCAn8IYTskHNZBzZIokkQXqyo70hSpIXv4Jj6oMbtEpgio7jRdjo1P
3LpVtyLs/Mzy2ZgDDGJrx/5ouAX1wBMoJlHsAg5Gk+Cma9AGRfBvbe+51YDdz0VzCpovw69+PwYR
P2auwNmmcVgjJYj7Erw+RRM/O1OxyqJBkKua8JqsIeZw0xDC1s+V77EfMrvjvmdfF6oza2yOUncU
7MAH0h3AU7NZzRS4/hsILXgpEpRMIvBrcwPv/0elLt0yoDEG89xl+JXEtXDgtmJSRuCGcCE4+P91
Ktt3JyYD+Ath3TVUZQei7o02FFHOsSzaf8vBvmj7IM2DwSawg5fC1QA6oyjZkLJ9NH9EM7pgZ4+z
3gFLTzS/ujxHTCFateDqjNXJEp66M9tfJUpHNYYh7BDtFulGUfenuYPqq4CAd9+pKkpEMgGfbwHD
WiDPsjTG5aHU2T6d8osir+4dKkrjXy78Si8JKQzRny/85qF72+jOmh61dCr2Aiv7oetw7jN/7UMR
4zAC9rdiFDKqAcuvtMReZ0yPV/rpBRK7MpeCwbzmp7EUqLu6xPu9sGESJ8MM9juwQd2r0toPXaWB
TPOe2jM5ofrYZYn3lr0fEoqpwN+BhLm/iRVFQfEnNVPmunXbNu6c0LeuOGfqlANzwv0O4p6j35oR
RIzI5V2qg5nkiKrtS6QuC/wwxxAeZz8pstDnmmUOW3tdN8MkydAlYys0faP7SkcCj2Wt/dRG50Dt
QE5PJW79guHfE9g7Fe1TCa/IfuhrRXKewsTCUY2AGOo1fsxGuDHhXVD2IBzmlXIJoWqhMRhshbf+
YgbbGJlb5yuMl1yca0pZ63s9e+G72I/jseE1NKIvSt4ftwYabHmjgj18kkuc1hgNtJvHGuOuaXES
ZAbrTcQ1BdJC74++ZFoviFzAn2n6rz7dMPhRmlD5ys1o8v0UPd+iFCBJ3e65RnN5aFTD9Q9pLMww
TFRj0iwr1u4KimWyQ9/cSdV+kmdvi9kqZ4qJ3j2UVpiAKWY82j7VZ0Jq+eMae/HO9KWMFhUYo00J
QWSc4QT3LWfBoPWx/76PZRV/jbtAQAJwzyZM5iPUby9GTq0I8BqvcZhp2v7Yi2FJMsly0CSf0iXH
PyJUjdq3/PS2Nd4HfZ6ncHyyScAZGzrZll01rgllLrLObjrZ7GpVlUntSC+O8VXvuRkIIIgGmgec
d6lARXGlMR1Sr3oYK/6gRbQhWZf5qCbqyX9waidCjfwnBnZY/5jFImPfUaf1X+zRgngwZCVNL+Lp
i6dh45Bv3rk2utwNM+39eN/5UFkgDhMHLKu5UTNhb/5/nOjt9NXz5WPXICZZ8nCH1nrwyIj7qZi+
uk7/sWT1/keYvt6sUwmyspFbG5lyG3RFI0N8QJzzFldwWA5l5UP1ko7q8OWg9X/Njs96Ss06upIJ
os1qZryV+t1sRSL5S03ddEXNfvPJ3Y6YF5jT0gg6sIzwtWVNEtq2mfpbIOuY/zBLxRiX0h8sT6pc
+e/kDtvYZF7lJOJ+JSX9YrPt1jB+CF8+0rVkO9LZ+R4YiJ2cdN1zeqb0lF5ZR03vbl3cFuaNmzMJ
npxI7H0lgmoNr1z8ARPamNyORi+KZSeQ7QPBTC6+o9ESo7BLV8P5t09dLYlorWjLHWOeLieVzLQL
2d8Pw1HZ/wUPNiQi8oE2j78pkv74uPGU7c5mB8B0FWA6zzrU0FgC38XxyAIC55zM1DFd84yCCAFI
tJvXBJUgN4FrxU8VrH+laB6MDu2GRWM03neXDzpMZaqi9FXzAXEcPnqplYL59GXtuQuQVHT80XV1
iGX2PVucyVSZ954I8PjzA+OgikYZD4xoaPqtxxe/Y+KP9mZ7y6bGBc4msk3TzcKfI99+WLSAU3eX
JwkvFnER9aZz22Lv7FXoyfvmSU6EjGDEZehzsFMUDhzi+zzH8Jf9ViQh3amu+L9Dk6ubnJLSys2S
LvsDEo/Os0TzciV9CE+Z7nu+n8haQlK9GVCjOh6y1AUIhwD9mmpjJbOkWUKqn8YXjEAJ6ZyZ6T8A
je1veUCF3dysML0AVQaJXf70r/oKFK1KWyooGq/1txwM8SXKhbTUl3zPUwaiRMqyaJSdP8PlfENP
Ddqh2pMiXHvWEaSlBWTH5piu7F11slaeJ6aZMjoGVthRDYYCEnk6TlB5JzKrxJtY7QUlOf8vvypu
cr7WGaGlebM6z9logluJPZN36tJXwNtSoIxAu1iNHsyOU6rBt00JCKxP+6DuMitR4w8AZ+Xzuttu
dReoXpEmmZqVEob+6ivwol2tcnmimcrmzuZ/JJI0aYGDXGuiK8dI836mZXaKZeABEyxhJBSyvDqN
8Fb9mGrjhUfn7U/MoTT2ZKmgmt2PG5p31oNTU1O0x1bP59Q5Q9b5enq+51qFXbRNosWxp+l4Sfgs
mlXw2/DAGMSfLOqxWYHmvVYjtu939q5bucsm+U95PDAHDP/5gABYxBu+sWyz8L42Nb90+DGeW7hh
PQyPXtmiXU9UjWWK3GSsCLA7CkMzRy8BrO790V3roiieA7O2ZyY7W1YGtKXyZ7QXxHNKUjdYOztE
jZZ67/RVIHG9cT16bPt9wao5re8DtOE42Gava8G/06wWNnNWo4ebrbYQ5KdPb3sgYJb3MAVuexHL
PQ/WNSAuNxRNtzb01ANT0ZX4ivbzwc5Q48GgChOTAyQtgCIo2BkYoBy9/tnmQfGTAcNyYZXRMaoB
XKzDPRTLrMbe/KhW+3iAaaTRIPI+ZMxBk1pmZd4Q9JixRYTzqRtuR5KNiZQUL3Ww/c4eQutd2Vf0
6P2BWRcOmuLufWbF9ETTvYIG12yHBtaaMS1X6BDB5fYSok1f1EMvkkt0HBbULCieM0f0kdQwqcGW
c5Cy5VZgo78Xk07TfcpYtT/95QUVMYZCPtZe1Zsu2vZr0W2cgdVrh9G+0I5hq9JrOAC5pZYU+Gcg
fzicrRyKA39LlQVk3Utk1tbNZVTK1Xnfu70SBggcTLRbWG5ja7KdeXz7d5doPebAyIh9H8I9NYCF
g3H7eFXno2ThJEPB9imp1P82g1s7A2C8F9CEE9JAdzhlX5R/WtSxVxV6EpOT0hUDt1kGaqA3UdPf
8IZ2RMPxJr3/1TrhX5L0e1cMTuVDNbsh0cBLeKWBxt2/Fsda1sW2cvItda4eSBhXRUl+R/lFucwL
K3xOZWK7pGbS2nHCO16lc1OMsQk/ppr3BmmPiqTapQixk4tN2Y6GQWh+70mMhi2HXRDJIEnTOppf
CKK4T+fj0J5eyPgMZWHtjIq0nLbDa5dkzXYDH50NeD7OMb5/W9t+pbmCHGMoGlcUIR2hvAKyt+gS
Qj28vJqNIxGogS0cPJ1EvBsmWSt8m9p1sVMrl/jBENe9qIuwpaId1drZnzs3yqULt3WwLfM5QNej
Qv5Alox98ePsfZOM64vX04w8WpQM/b46/EJsXdUvn0si55tOwObHNoA6DfGvsE8kRA3pNHEdQt0G
MpSmat7jDQAaK7wlf0JlJdEe82w6xp9nCDJrffrsl74a9bN5YI2uevhTjYu0m/3msdhMCIi6mi2m
348V9cXmRHQw8GJx4+v84RktKbL+Njo70V4Si5xffe/ir2spOZfEkSCVfsxqiplun+sR87yhR7Kg
/p22pzG5VCOPyAx2L1/65yPE3AsQspwFqXbFYS1QaYxRsKQeyL4m8gXf1C4odwHn4SS1Bs6S/zVe
+1wdUHXbMnyiaPSCI2VDypDHzO4gIIt7Ewp0z7n3/7KcJn/VC29HpRzd1B24WQvnatc/MRbnsZ4e
Uqy1PrNhls8M/7zbi7l5UA+EpMbM1k+3qICS+825yRWdGdamMSqFWJcLJ8/F9SfzzaF5AEuBjTPt
MHgAC6zz1Hg9z1AKtc/Z4tL2yORFw0uuPqioMQb6GpeusH0fo0TEr8u4CvkBnG0L9I7gh+7pyqKe
l6XxMiIiGij/oV+L7ILrJLtWnPUisNKjLFi8A2ZLpNSA2NNdtQLKKfZZ/UHeVeSpeojjEb7JPShB
z0QjQet62oPFfCx8Lw0KCNsuBIzJMgZryEttK0xpnRof3UJrSgcvJgp5QwLxCj/L9l39PUKDpn+8
NwZ0NWjyN1gxHqFkBoWqmxXAqx4h17mVmMcRCy4BQAShQa+lrHdfpeXASrfZv8zl0bsjZlr+BPg2
Tghv5qZoeuoyxQuRj12hd1rDSs75fk8GfZmayw0llPpXK5yMP42k/x+IRZ5bhn7pGwMUA0QqDvyU
4r62OEB160hygLRhgILfXEARCBO8XICXhovfeFougVDRtUi8Rkr6ZSKWFw0GIMipWA2+YJ/kZ3vy
uynlBFt52DMuJpjsUVq1RKr4pnV9pd2VM1q5M4vTacQT4lTtBwpBLeMM8k2nlORT/hcsV+R8ezfE
cJL2HSL41PL/qU2Snat30eYYOvsDgNuPg5j/z3Mtn+L4EK2G70HHnRBWTsqIvPFgZeqrKcmDHSpx
BeRHabHM2A6nPK3iint9ScZ1Ni0wAPZEsajX8WNIVePEHTDevjqgS1GrtqHRBt/wGUzUHSwS1lBG
e+DRiS2sH1he9vrJtAUcTIQeC5EJvmRAbOnp2Ea8Bh/jvc8smDBFlnt8BZCYMC71AWYc6tTq3ICE
fJ9QAYaE33CpnrtDhyUqld1+2Y6jJgo/m/abqpgW9SRuqP254Lk16z3e9xudfUVYRkHFGA48h7cS
cCxhPYu4tU1vvQpL3UoIAwGHJCLob64Uy0y4AGIbobAJMelQChH6s/lAkd4nE7Xh+bMco0sghWzX
3rkKXebN3A1YmBzUwXELidqNbDCuhFSLmS55/C58RrcY/GP1r6eRWaeny+zKlgIzVX1B47fhI5+n
okr/ITSUzhocw9JYgig9iKtR9dTv4F3SjtCpbOVcm1v/kWtSJCEDanLvxBwQAglZjjSP+0XJJ9nO
dRhAjU0hapWDfqbGbEE4OFE4H1ejsy5E4Xy6r5/jMXSy1uXoVuFy/4/JciUmB+7YNWuH1f3GlC5c
AErlIG32CAGoiLZi3AmgsOqMxZEmuEbbgUzdiqgyq4Ig5SlsfkeF8g76eEWr04c0/9QbCD2rL+CS
hrzaxgaXeWBbpcxE9po7wic8OICE0vacgn3BlS4jVt7SCzBUYNABVsAPw2u+PUh3CSV9Kjk7/MWR
Mwq6RvWqgN5yTNVoVEm3Y3Nlg85NYzu/h6LLDjZR9C7wC+jcIYHtU3kKJ4zt11t2/pJ2uOEAEKGr
3gFckCDueqyNDvTA/JmFL9xlQBt1MnuGIzxwyal+qijEieemODPEWausOZQM5fhGd611USX5GQRI
eyjJnmtkDgdAGdW+of6cmgro1aH0+W90Cc2W1BSYSpPC6L+vSBBS1q9s4rVP1BWeHUJkEyKB0NDf
1nwr7HiCRUCDpC/n9PI6Gv1ECd7UGOJv81I/xPZkkrOZF6CyjxScakN8nNNxXtfpH5PAeJz9F4Jw
yZ8UNmhO2rxpO5HncPk9K/dr4ZEMJ7UnhBUPCb7ArFUk3c2l3FByIdecFd9oDKkgQRyso91nVhR4
8+KG+ycRLSxzekEgy6fJBR2+7U6fD5yKLbhwL9YrnKjjtyGln9RV0OeINEGjL6GSnZUFYr0gJLfy
xKgAE/CbSLQFZpSJxYRskokDOrpXe7HIVeW95XNkqpJ6WJIrmTBrVRlFrWoP8HSYFguJ9IL2uPdV
pTt9cefpD9kHbmq5zwX+XumCklu5s5kMLKMwK/8avrZXaSUuFAXK3SCzLInn9ZNCz0U2lv4C582K
zILVweYb2Ty0dDZ5ap1zkuYRWHF72O7I/2yFkmUOPU/Nh+4nAUKT9OjPP06MS+ALMwu/YSaRLaiD
AqLM1LpyxBECXaDc8D6uQwfC/28heKTrDJraj0Q906TcG7UamkXgNxAeFibwlAKdRBXEbgnTZLwM
EWQHIkFOae3shWYuFsIK2Mse72rxHvJDaVDbG61xrRZNWSKIdUzvgNYXsSVJlTIQ8zgrfTs1VRJv
QcHjLtVN5hblzeQ06+1gEKHvl2TiM3PoSes43ZuBlD+U9o+8z3b0XdJKwfa0AGK2XzKY3L9gUZX4
hlmRR6h+RSenxllVathgcqs4UF/vNeB1Q519FIbhlhqA4v3G1qkUX3xKYb3+ELPX5e44NW3ix1av
4JRqxJC2+AKTuXaKFio6ub4LCjnSr3EeyHxurlDlprHk5eLHVT7hcsjxhcLNYwMTCo46u58VyZnG
J6yxWfv4aOsgmO5Ajrs2FORGxWoPF9+zZh9r08APV0Hk6dcDwhc/9w1hcFZNumam8bu1RZuXRWOc
2N2O5IfSmf1Ce9+tpuri2vOMW54ovu9m1lkT0vP/xvZerDTooXprSjKIF6gPbBtItCPa1eXbZ7aA
4cknkLn3159GTvwgW7BK3lv71CQmW6Hyl0FdyqGlPH56SWo7uzMUEb9TuWxH1/XBRFDQiEbA5uga
XtrNawuNlW2TlXahglEBlvCMAQ6XbnpmZ1FwZXrAZbohg85BPg8NpBj4NVUhxUZKhmmNkaELiU9T
iisXhz+PyYEf3bmfQyiDr+oansoeUoL7qTQwl4pwpYKhPllcqEtM6PhrLM3lAPDog4a+UI8KpfJN
Aarv6kkNaoTQudAlU1dphfiReDmi5R+xLYCr4MtuJDl1WySs1A02cltG6MO3VIvQBqeq8YjbQ9Rt
UiJNRr+oQ7yatE2yFHwMqHgo8+Ivj8d+Efo8IXU1QvW7Q5m+9z3fXblkvmHYgiCIdAl53YY8tJEU
VM1odkhCiv/7cMNQvenVyE0Buw148gSSzeu7LbFspJt3TZ6NFpusf1Zk4Zx609F5oq2qQtvHApjd
AjRoF/tHm6uw/sgmisHgB6fckDcJ72A1qc32ZFAJu3+pVPGVNMvb2nhiOGBMOvmvwAn3ZmNnAWK9
MqDY+QHSYhKGxwuHu/J5a4IeKGKu5cDh1f1xr8n3QO/RR7QESLQXoUBkAKI516s3DeW5Fya0WDGP
FJgouMfzz5eKqPq9D8RjJzFXHfLsPeuja0L+4f1OEMrxmqPaojFfv2JibzpIXgXfQMlHbwsPboRf
NfEGyXwu5/9C8vm0UJPcZ0qDRbeoY+Psw0Tfg7jAslc6cjzGs9MuOb0iT17w0Hbb5u11Qoe0DgS6
mutY/BypB/IauVMKIr5OPwOe2QUwDpB8vyWRnf0Hu2i1siGpaVh9czq8qGQtNO8kYY7MVQlRdCkE
yFb4Zj4NImoyr4MGcLlABq0ASce5oQN1xpjfTsZ0D4CsSEQPxCr19DLRRKcZxGGOgy8mhGR0k2xj
J6melRhFpsVgc0XyCcMeMw1fhFi0E43dF6Y4CQbc2J3/M6qrwp6G6nPoWv/tw1xjkDCoOTGbwO1N
vgSuZBZJTwia61fRh8TU54kN7sjL9F1eE+4d5jas7ecpRaepr48sCx0O3OLwTfrpXIIAldY9SaGj
yriPcUeps8yJlMy9CUb7tM3hwyCGehbfyLeYYkniUmC2fcRvC9Z/On6HxDEHcXG3RulRXXFVnrXx
NhOLz5ZNp70cAuUuA/8+hPBThg86BGA/sppsXy8idQMTwuoKK1G8YNr/fTBhABAVHNbsJ6eNooCq
nHuOunNQrLG24LGbcuryq+y1UH94aAxZsg/AOpe7VhOWOEpDjn+2R8OQb4oltDZSDq/r+vlGv5GD
zZB9CUXNZnfWJkTR6OJHGUflbf6CGC2TW7eXTlYnDicaxaiJw2xcr5lz45i3Z83r2Xm7/l2+DScf
6R8/BjssZfDizNBGh0TEc8VBLN+Wy3+sL4S6mYiSdEx7c0dqmBP2ctdiBznz4U8qYbAyntQXmybs
PqJHR7tRjbswQ6LgNwjoXILeYRKIxEIUeiWC2+MJ7nM+udkLdbRCdupZroRsqVGP6jFFSXmn4L3+
gPMpBWWoFbj5PeuKsjgBP6Mm0ZE3NWZF4lHU3uwvfIyUg16CRCs4d79sTNDQ3n0iKJNoPgRkrwB0
FAD2V1/ng1tBNGNfyhM25nn7DYl0YeTBRQsRYzTd/ykKyazz1zdUw5iKqZU9WnhcBO2rD3BDGrEp
LDAayA+Bs6ZyqnPfJCnb3IIPPbUZiqy+Rme8vav1f+J+pPyeANCa3PlFQ/0y/dYr68H905mkQztw
lAlNnjmmrgXFe1HJr4fAZDaRL24HL0+KSmtouEcuBpGrM9/4Y2cY3yoTkj8FmecpBYW7ivOZTixt
pa26Asvf38ntjM/tdbkWtTK3EcA9gSLbIus2kG4pXq3LRK7T0XIaHmY1agWdTkXfl64X2M4EbfIx
0eQ6ZpFy+1hQjVPfJMncrsp6frqRq1xiz4axljNm1V4Sj9Nv/cEABN3c2+zcwwzro0X+GEfO8fom
l6ICewHXLT/NdayxTbN3b588v+YJI6T08xkzf1AW+O+7Y7EubUCiHTfA8EZUd/0Zsvv59PFU7jth
yyxWDU8Ss+FDmX7k9cDhmTw4vQ8rUK27l1cz/aOUHI2+bgaviEMECvuYYfu15MP+3c/70LofrSsb
5siT1vAM8Mkxb2AE3zjV/9umGmL0hAaVQ0YD0tgkMjSCW1tW0iyhPXEgew1EjTRSlzVcdGCARVNe
FGjA5Wb+yxu9TVUm9dSYN0BveKLUP4KqntGPSQbPcMROBjeQL4Rnlz36CP6laCKruZhs5lmkHYRS
sFwlJj/qBEas6cQN5B3HGRZkCMsF0tfpqK/0E65aqptK3JnmSCQN87Ubrrv7myI3zCVHbCNU6src
vFqBMcjiomSxO15bOVWhdJ/RaIkILuhog5wdqtvKe7P55A+MMDJqDPtLMuXt35DErGEgCWS6VoIU
dedA9G3fjuGvSH8cZ2Uel/nPu+zbqA4Uu+hYzRiULhRicy+c2VObZLX4Kk1vxvTVluplOQy73SGU
3LV3Y/9IgRLkfMKpBU0rb+CtWPuId9O6oTQPN3UbsQJo9co33ZWsoohCUC70doHnrM9PHdUa2Lf6
dCgTpw94TAa7lN5CBYm10MMnvJAv8vratWs8UtqFR0KJ6wB1dc5EiZ4WguuRsf32B/7z/oAYh8sf
DjtR2StWSw3eAlsjYBOSqhV8Gm7jAqxXYpBKm7LOr9g06XhmHC9igpb2mUEzuooKYxhVw+eOMYoi
8cRlY0TAbxRPuOJPfJ8bA+h8F+ACbiHrAHUVYMgpM6XtuIda0WhdjjxSt51GA3BVFFSrm0kvpRtX
Mi6I/jmjdUTtCqxepQpAzQWDvCrM1g2T4+fNVRpyZMyQ/CPxYxhe3CEcxpg4/PkQ6tILglxz6NkA
YV8RzfUycm0YiL+adUAsXjBMJ4SouYQqruEEV5GaTYaniu94zgCEcfkh3HxuPku7/AqIwfWDkjpu
fp8Oz7/VKlb1DkM7C9Xeq1Ywp6xW6lXF1vtqZ63F9e/xyZ2UJpJttTF5tmlPy6rb0oNjoqKewTJq
kz+FNt7jxJtcDDQKoY7SG4A8JA2GS3PfsmUUxmS8+viOhAgPRA6iUEnUAK+puzNE8cqH7XYaqEdY
ty6R//vkMuI51RNsqI92/F0EqaQtCR9ompSH2ip/5ddoZXZha2cH0IxgW4NJKXGUiqLeqA1OyVNI
R6/wNqv5884CSgt38D7dQCMiR7Nurwcec2PMMk5nLB5YA2QMAHWeSwuH33dOt7RUi0ec3AdUJ7AQ
836m6AkHu1Y0Jz9uKx4GIFi4JW1K0IqKxLph61dkdHup5rtIqxxSYahUO0od2H4oTQRbouYfaCC/
8qIyBUrybfazTs/hDCEn8TIfNgkygmR5pT7LRAhicnPmUVtA3GHvLt+MMhf3xxl8JGTkCTGkOpFn
AFPQkLz8iBfHjEmPm8gG5fds0HkvXRgocjbtMMt64iqmY8HO78tt+glQyneWRAw4Irc26a6Ikiwj
46seDGYxTdR0noAYflm+Lg2cSRh1F3Ite0gWeZTvHTMLnoEGWUfGmuT1gl2altUVdQFempYRe71Q
Cuxb02dD8KkM4h/ootcq9KE/VOVcxn2ctlf5ELCsJ+iTiwd6Y8FIMnHslmcgITkFtcxm5kpxeT1p
juu5358HzEnDTGoQha7LrMWpypJiTctCo/QDSSjZlUyPzgB9mpRv2iH77VRTVxXCuMJWKfxcmdn+
mP0CGhK0XDp5W8W1m7EewVbmlBrO4STTPTdOXrkCF+ixpzK4xOG6HiezL9OUpkyf6rQTveCUEXx2
e2w+r5Tior1Nw62wttTAdZDeCc4kdR6QKyP8TIEzWR2cerj7hRjNyS6BZQDZ++amXVLDGZ+CfKyl
SLKM++jnmzufeEaDUFCGBUahsIwFLXWVD2V3JUEIMvzPQvKIGbzAKTY/jcYpbDx/3Pm0NVaGV4Do
LLdEDziv3qtWkidCraqiDzzDVA7dSf+s0rOvGvZnAuIksIntzbawmPiP4QFr2P7zZ9X72lLHrtxn
leDvO/12Dn+WSIMv/mekVVpaPbXEQIiW8sG3Pb6Ku3uX6DS2UE9TlTH/A7NbsKFakiCPK4j+QxSU
2UdCvXLF4nfUJmzTFhqoKhk8rhi4T/G9P2YPir13AL9dqoRMs+/CxXYC+YAZZ4vdCrsZmKpUtEc8
nnGRdsiGBPlsF6H+IrvBp3MdiBqhtuPk0uQejPLOmpwZJoZILmGOwSnITRgFT/08i1VZqFnrrzk0
CFCZWRAdZxYaWovCppQGGhWJGqw2KGw5JzlTzGXaKpVq+aXDC/dnwBDrAxb4JtIbF68ACfT737X/
jhF6zIJgDcjAwvOs5p0kXaMnOoeb0YOMs+CKvubUqGA1bjjZe27ITRlK9IvStEFuY0VZ+Sl2BFdP
g0EHSJFgW9E5On4Zz+9nhbFyiyItZpIF4smMHrLOzsSd6e+CE19VBbehTZKcWjmGxKgscKDDLu9q
8hVaM23hFuznRj4xnGZvb2AJpPXQU2u7jEKLRbVzK7gKyIDsXHN0dPy9XQrutB49levYBrT5tyUY
tg7bGJGhDtrwZRNEvo131blq+koUHOqZcj76lhwAfNN66i4twNsgRX0/LQc2HwYVH12czJMlCmRH
bBF8nVLWuK2FN5KT5RqNpgHiZk6fyIwztXtfgLZOz695zGqyquLrYG2+mUmuxH+pUsAtBlpKHrmz
H05M7VT0QVLizGXvETQm5DMbw1mNO2rwBcwvFlsRtMzxZEqnPtDR6nkUo6FzYxW8kzF6g91synuL
RLTBuHjKpOB82M+BAFfo7POLeo8l9eE8Ic0M7kj33forBNTRdKLhor03JQrXaolQGwja3d7lqBHc
wTRG6V76iHurFFx2yb/n/49eNtwhRUCq5HzmkLqYOELlAG33yfd278QUN5rKX9EuvsCrlpGdsRxS
b1XQypEoN1vANAdZYmBbCO7uq3pwIKzHeYaAm5O9Iwwr07uEZNmkjIepQzgNMlFqSqvpiEiXQpYc
JL3Vh9V0icNBWhaBhr1Mhh8EQM/PfsZr7TKSHUoXT4P5DD3fdiplAOeTYUKG76xGzy10DVfldS5+
WFceYVGDt6R8o+Y29e39YdnBcuB40opZm7F8KnwTN9jA3PXZ89Os5i8l6aRWY+tjaFsIQGAO6vnf
eqeEmqMDZyYgvSsjHmgCzNE/9XGIuEYLQAYS2OI28fItEl/5pJcPPtTiVnXNGCk0/SdLVNnrEG5Z
IhcdcOhLjLe9Bwi2PsCofFG6C24ZCTF566PdxtI1LY4J6sg6sNd79QNaXHNv7g6clDnsyA/nH2Zc
xVIUJ+AfKfymFehIDDK1jZbVqfvUUg4FE4RVg2L7zZZemz4D/EddUoaaUBG8ejh7D9IjlrsxLdAU
Lhn4dwKLsprA+wJ29aPhDlfaNpzDS6vJ1AfbUiUDojEJG07oTw1kKQiGU3uylDCGNuZC8dCv6QHM
Ai2/lAZkSwvS0PkGACi6B99clNdCkbdlCU7rs8Q0NcS1R54bXOS6L/HDSfyhZkOMquRcX/IT4Q/H
XN5A9GUsBKs1kZfuJefo++scvMYRxman/DDuaQ8p1FqWNugQR7F8eRbIlrB9J7MnvSh2/6jJ6hMe
4w2B9WJdzfYRxnAEhGC3AtvUcPeqGbukJ87toOqH2yHrikZzdZZpsVkr9GJP8RfaSeBTWj+HOrcC
4FYLVuOAU8bu4dB7krCbYA2cpxlOsg3yUT1ZjFLGrb9LkZC7VuYihO9CL8k/nQKi2HuDGWvp/koq
Pdz3njDgOyRD4qIxo7rGDSs7EHBPPEXgaUiTfQAfJ5RVJJE6MfS+/ZMdgUrC0LsGlDVsXUb43usT
szZ7tAocC9tnvSuZNUeNLLxUkVKghbScnnZpaqG9wIMwdsWdWfAaMV9uFMZ3qD03J9WcddZQILcN
LPJ4T3srybW1MjpAsHITc3sBwlx4YZKjypUw5aMBXy+NdDMhkGAFytFBX7Zl9qQ4FCS2l6hh+HND
oXtnJ3N+FiRUPRRbOHTrGdre4zB2IdrRAY2SI90+gOibgWYzHVZ86pIh4PjArFBFGNZNXut5PGMY
BJGwRGyUC67m617Ysp7POkb+CxyuDTwhyCpzleDd7hE7CccctnBHAOYaJ75NzR0egoYB1QcnBxl/
E/YkbzW3iHY8LdcKnhLe1lsCADS6M8hAwGLHsVMibpjUUJ7VYoZj0MSUiHQKmA4kF0l0IG2xNFMR
JaM5xtgSJFiJ2RQeoACCIO9VjSAoa2OiNIcGXtJQFo5a2SSclChRk+Aas+QaSJuDbV5OV3pwpGEv
OpEkI6mqx08QutHDPs3ZzA8ziqL51wPxGwOxlKOWZtZRJgi0eO+IyhlKlDcM6fmbpVuyvsQCxXYj
ZqDUst6CUTL49S+sa8OuPRIruXHlCHD4FXibZI2OKWBZt6FEaKSctuwjjVftSuU8lQf9qfP+1QGb
gVDm1Ka4fGUoTh2Y9ejw1BkFD0uHbRAt+auVWsQIZME6c5pbfcbEWY4L6C/LNE93YSEbkHOvXBHn
8dLwbiCYnmQbYRKW7kMh95BeEz+284dXdtEID2Ebc60xSuoLG+i+xDW+28hzLo/g8s1FMYw2tMEt
LoPKX3wV9eK45pazgXvAvHGLw976gMkXzFHTX/xo9+bo8sTzW9Nq9wADNCULYUqlmCfBJewO1tGX
76q58cWX4A3i8lz58cJqdy91ftSODoT5Hpsx+J8w89LNwFqn738pU/QdZr6aRtXrN+dRS9j9L/WS
BpTJ805GHF4EUYZ/JhUnZN/lSmPqvDt9M1js7o5BasOvl7ImLmKiN8Mjusyat4lbXu+GiPo0SIc1
yZxDrXaz/TP/9fimyvlsunWJsVOV1y1YcKsdZhfIPmhhvFSV3wjDCgF7TzzLNat5ru9yrdMJSqxA
PU46JRZOVW0+QjkBPKaQlw4SzQ6+k+YuE44AH2+c2Jo3IxyMEG5gVkbERTuHrzKZy/BGbdxC4T8F
eCEFEv7Tt+ZZTdFy8IS7+gRxh2GoyzAIlUDM1XhK1GRVgz6HULOAjIM6hUSGC2nNv8lfpC7tzwLb
CL+LyxJGz9yEq+Je1gGTOSFehtORLvjerRNXEfU4RTJ4WabK6wmFyNyETYdw7wveLnZFQfgFcPQs
+Sqi56eoyY+rXwG3gHoGZWN/elHj3GrQ+0Q2X8RYIt0opBvWVErZu25U3CMAEWJRO7pEBeZTkD8B
5SqEi8SU99+Khr+j26AV4UuC9gdw96dBI7Hobyz7bWBVSzz8dUw9gEVQQ3rIiPSUY2voNDgMljqW
Zi/ObwoSW6WWklOkzt8pPvEsNijoNYeWLLRbb3q1CB7FxezbuUnuDswce/24fSeNrXvLoBaDXKVz
ya3HbF0c5QcKhKihJpWiygKEvLsifG6BGlQQtPaL4ekED1huPR7l2CiD8nfgw/y2d/Hk4LLKhvp8
yE8h543W2XnXpben99OoKXB1Lbt0sWYzcExwAcNaF9hbokBm1rtk6QlPdXDflpsKTlZfflHzz8hH
J5rInxzdqkzq71pwB8R11r8uOZZyK8w0p2OAbCNADGz20eDsHQYqEyMf9e3uq13KM1rkWzUApEJe
NUf1JW8CO1rGfAFGW+274TZ2ojX6BpqFu7B/aEMXrYTEV4EU6zda5hCe5n2iscHH097OpZlpj4Tb
4qI4m86NaLuFfq23eGoXCOBF4DD3tPtvk3bnLIw9C65YPMbbhhSBz0kwl7wezXqYAugOSAczb0BO
6/zO+RSmyqIioHn+pBkppPNHY2tveh3KbMgd96XgCilvK+2rOSgumIrMM08mjnS1FC/Pk7RZCJ2C
tXMSurHE8nkbbu9g2sxue59Rs8Pv1kp++5QdqJVDPxHj0fJKK+hcBwD2bc3/twsSFFlZ4ofciw74
FuLxR8Lp/CFGtJOdnxbitOzLq02pQ1Q/V0IO2heHlLocp5DhEGVl0VE2G/m5ALR2Y3/VXSU+4WKq
QHCsTkIuGtC1TgecS/pdmKDJIF8E/btI4L4qyfQHGXSatUSGtVZwvDi4LcC/MHofU42A1H6ZP5Od
tvV8BQzziCm61lanZoiyiYhl0zYsKJ7NgEc6Um2E/nQnuGvuhls/BzqEGic281FNoEsBsZ2Jh6RI
sUF8seNNThmLzIBcUJwJsiOSrj8SrMBFYakkIYqlc52eskN5E7lAs3FR/AL8yYvGQUV3sbFnOo8X
xOmUZzxXYCvTxCqGAzE72X2On/Iq8Ds9hiNHNq6Z7MK+/cJGMpRUqQLtVsGZUmcLq1qraZjt5Iw0
C8gvyFpmECrFHnhTIwOfGarzccHSNxbecwLDMQLaCLJZg87nV+WypKgAJW0Z7f7ba6Gp8jGvgPEy
IOia6AAFbpNRbOqDb1s51StjSjLA3Rr34122pQK7llojTrKhorhEgCMWdsvjNHp9i27SVmtcvtuL
mPjyEG1wSAW/HdmFvEGl1W6s/1hIghsL9fk/hKsKqHslHKftfkRmSxcKMXeOV9eC4Fm/x2+3rtxp
438EqjuqVUatxOfFhBzmE690mzT6OBKmMweqUjLk7tpcuUX9fQdQTARVK0chJVBvx37no9ztSjt0
WP4p7x2t6o6nXJoH7Lf6J2L+pOXfrt5NuehPmqTzLsbwlsR8dZi6UeDPXPP+G5eDCnxOW9Uz1Zwd
Z77scyZE4fiRza40ZwJwxeYmywMStjvRBo1MUUSCIpmNWupz2w0iDP8M6uNRKZ6lOxANgvrC15tH
ZN4rR3CqqHPy3WO7ilA766jocQ1QVH4hKY1QPD6WoprTWjo/n1j9qdbSOQKpjDP9zJ6W2J8WkOAX
RXfLzB1tfCQ68J8DGtrXNEYnhpJ13JTWIVoSTRz2z5kX2+QwnpF2BxYZykwwDT+AL2a1/SnUzKCB
UUZiN2fwj9elJntrBfPAfHT8zK3dSAaVRSU9a2IcL859XJ6+gRxGvSJo/YpQZZJrsP103IhIaMu0
pveq1+M0A1UTnU6y0HG3Ch2LzBmorT3XDI87oQgEcQqAPCRWRstz74wnTA9YlFPQ6QEWRMgxJyhv
PodxcqxvN2BvWdbsmH9vbV5hr1SSdKvUmZBX4D7Ak02tCTLe46vrUTgxEubfVhpzNhkOoweTtlB9
f2Y6cZk0aqy/2tEvANsusKXSWsrX1zJISbCysxK7/VWP0R8sMtKtiYc8oR8ZQfl+vwlcY5q9AGaK
7g3O6/AfJqqJUkRzFvnxdIbsMYwXy8Yx4gmQ+l5kK88plpJnpCN+hCCQcf8BnkSQrMbU99mfKiR2
IGeGSauED4j2XFgCUEZlbUHCo7N5RGl63VwIU78mCFZmqVMWW8yuEKKEbYIxyIPPJ6o/t1/fu3N3
UdeztaRyowf7z2zd/nplVgDt/RlMamBdwrawiyH9kiZkE/LyS3qMgHQrszc2+22qM/kk/PyeJcRY
ztGyL3HAo0pVW2U4tfgpTgHtT/pV7GqOA0QWk8tgJEt1rWQ1205XaWYBHWr7uOR+REiAlsvJSkSM
rsa1y77u8Rg4pndz5Fwqb0D5qxkbys6byidsw6q6VDUwLffSQf5bW/C43pRqxS8jGU+1oxb+XqjW
Hj2NNkFtQ0djDO4KDbIxo19K/qHleuUhy3+El/IdoarxfXiYy2mYy7hxegpyKCcU169LgGMyN8ZL
UD7fN9JcF382Pb6TrXOSu28zYr6lbVQ6RLyWueSitedOdmSKXg2GduVj1cJXAK1lDSMdGZEud4LK
HuIrbF33/WYa+A+FQZwCvnx1uCPm2+INFdT5f1PVEBc2pq4fRwYKEyowM0AC9hzsuGiGTHKQaXbt
oUBItiGQ2QjViZ3iibKG/fyvhweSm9G+7EPJCesUwei+NDLXTvA2W/ZL6brIgDcfuwNauf74TahC
nvuNZrCKImyp5adB+wTdujP2m/cNl2K1+SHsImcdz0G7/nmZnDUPSmyxrZ0uqNAFmxPW1wfbcfDP
7dpbHbvtHvbDRIugew/jMDgToa3CDIVigvb7ErI3j6QG+2vOI+LoSEaDFseo/JNzFipQec+2tvCa
kvi0fzKsytNmOwQQ9qRMtz83minrlFwm8G2RkBa/+ceY2jCAAACowwqsl2SFJttzZOBwKTiTuFEY
6ay7ATT0CO05Rn7PMm0CgTph+dkbRZ+cEc5Sj/I83cpj63Tz7NbHCdmKzaeK6jGCkYcKYpst2G0Z
2lQRgsjOEGtZQrj+55yZSyeIJW+C2Ww2d96AzLcJ79k/uzVLZ15m003E4UVoDaK9lv6xwaTrHbpS
YuxBzFlgYcxY/vDlyAr9l4Nn3dhe7LpPhMRHL3aU3bmGMAgWBTM9jlTAPu0T7b0XUgmjIYpOReTC
HfcTiyTTGDMghJ9yulY8MADg773Hoy0aTTFLkCh2o8mzRGTwaE5mdrTcxQLG/DiIP0lvuDfzI1n1
ha+k1k9LodtyiB+O+gAbyk63x9AyDVzu7vEXEHzz4NdlglsCI/Ce05Qj0zk3eCSOd1p3bxR03tGU
QjIUUVrV3yO6kS4udSWHTSe0VjHFXd5x8anJk5HpioidMCSknxhwrIX1KUFB4KWcRR5eYFrsTV6n
1Vfz8ScdneO+8fGwqDmAvmFUag4/UuWCgLAS2HozzjLP5W8EfYFGFE01bMrur9ZOMoaY+P8Razyf
wMBMAmzhH4GbZICFfI37H8UWJtcH4pGOvaX5dQKN7OR4xFphpMwL4dzUZYdYOWf52QXg7cNG7+Tr
IqA7czypsD4tFXcdmlkmCTYIY+YtN7Mjs3A4wCCzoNXx4TBugJViEKsv0imDA2DPAp8gJouQ2obI
ThiPZGNKWPh/9UZUZe48p8uHuOY+m5/JO7eEzO2YnznaS+qgMSGP9jpfi/z7lPMFhUT93gYaEwFV
BsMGbyM9qIdNQXpBkRQdzV35NbXx3WsXkc3Opgi+9AxPWJ6MhnN7otTlsabv1cZeCXBE+Sv5k7UI
ly66dsQ7TfcyOuU2eYn5r7ovzYqaFfLuGk9PudIfEilmjhjK798B581P4uX6uXURVV3K0H/YZyVX
fHSSbK6zqwAvEcFq9EK0k+E0JqVsziPz6EPRXF5JYlyqfZ1D0cCyrlHUKePJB54NDWz+oA+oesJn
Ombapcyjzf1UdpF1lieklE8dm3SROXWjkilJlElFxu5xQ803OC54a/4V4R+qtB4/zY11D1Q1cSsD
5MS9Wp7G/SX5me7iKCeciLis6BybFzHrvus+cDTIuJkNBEfxNAFJxIyAfRQ9M5rC/q2gZAnL+g2F
wwzl6lmMEmkn2fzdV/vGb5wF/Nuz3XZIdpbSR3GbJREjKHV2ntD9L2jmCXHFrs+sWByVJYNKBUGy
SZd4jKfMOxeqoRxsYTQUYQGXT3ZZ7DH7Q11RiRxrGm/jvc31TC9aK1ULWF42INT9gNdCwuSXA54v
X7s+3acImnZjyyxn6WLGs0aIZBQVu4bqJnwc+9p75V8KEnbVlIThCvfpEL4sHNzgWi6n7QW/ND0D
BqP+qKTtYgc9ULJEQfJQ2Jj+7R9gr5ZgcJxpeQeG9Iew0ul1/9bssvJ39tQ8XFfN6DSvawPywhtK
uE5cw1CXYsoGB5tufhP0uyaBLzStgt80MKfwfVDlzzgeCJvXAmqrc2fv1cF56aXbCbqLbwkOB6gy
PZsUPga1M3Avkaq8B5MjYkor7pQRYNtv2H5l1D1t3b1XJb3GzAKyHAVycGPWbJ0ZtmN9wW/rGU4W
vY59azDwl24D9IP86KiyDQP9JY3gWSmUsLe7x2hUncIrRHfxESbpCj1ph8jL4pErcWHuENedjOJ6
/y/c7XgjPZyOng852tBDuHGkwOdxiJcLcLREvF5X
`protect end_protected

