

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mCyyeqqjg5/0TkdJEsEEwiyDfrhah9gG0fpTMwUWGOKZ3he/dpUva8HsS4xtl5XP9zdNgeOXA7QE
z8wIFX99RA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X35C+3C9De7vC0qODnacg9gsvk+3IzrNpqQYzh787Czr0LrIg4SN4n42C6CPfkCBLDXSXwC/eOXr
yWqN/Hj/SYBmrS5kjeF37AKShalo68kYRaZgUNEiNvBgjtaJt6WRpWYojbh+ogFdK3xIXCNq+Qxl
K0+QDwwSCDU/YMofxGE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n73jcH3HYbuczKsWgG6ox7VZK1YnHzJQ1B4KxEg4B/kZylbLOe/lb0i8/kn+CjmMlUuMK0WQWfed
hITAZaScEDQ3B6jcHH/bNliHMpa5PCxNetq1i73KuqIUSMzdaxGWTSuFoXR94e0GNel9SANUqOYF
vTOS9qeLaefJfWuMi23yYpmliTIg3f3fAbSdeAfef4vuNm+0XcFw60RpJQs3nrsFq9KW/GfqXw4u
TZNQUQbt6cL25X91FZ9ygQq3zmgha+CzhVMH2888hx1Tg3YKoHcpCHNpnuDfIIlbv8c/WTDMb67v
IK74ph/GlcH+s638TtetKCgz1jniP6o8owuM0w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lgEz+Sb20/Syw0As3tLsdRmvucviIYGeDJylwgde+NWKzNiVP+by1Maor4kKAxxHjnI5lkH0wLYs
PhqSC4UmzjejXWlU17tjRxtRz6BbrpAi6gmDH8SRbE1L1vIa3LM6opScw2kIKRT06DZ3npJLvb1L
GQYpSvbMBpeOoeXBKyg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cuBsFlva1Z5u1UA+GZT5hw/3RJ+t4o7i70J4gtLUlv3Ik7QI7QGdbqQ4mg46AQCjs/XyJI5tDPDQ
SIWqonbFU6W95Sa+82Fm2FOLny1XsFw2bfUdFeJCVtBal0R28pkG/kXPwJRvcecEIrS2a1k5PBE5
sZrJ66qcp7DI4wbfzpv3ic5F22QlsAxZqXZEB6lBkhSRHmx8sxDYGL3gz3qyqFuTzoFlxGj0D2l1
7IJKcs+gQikUKNCj4QKZQHmP0x55BD7tR2tDFNHuJwLQeErQDiAmIcwGhliqTf1RxwWpWFh5JUyZ
nisNHaWXl8SFhFbWbHjUNb33VdqRqkyTz+gZkw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49408)
`protect data_block
sJ/uEcngy4mv0H9i6U371cc1Z7e2xNJPinmUZuE+aJJ2L2U1BH2CHbDZ645Vj3svDBsrA81Is53t
8ErKYtwvzaSbZfQsmKAroBgE5t20zap12jRBG3iQZlk7sOf9InC+LVym/QAFQHI8XKgr7Xu92mCB
QYUZDJwPaWH+lMKZNfHZe49dQ/D0wCKd5e01+Lg1nidshdzZCG+C64BNx29FmuPoWs/S+LqEVlyr
hmwElax2pVz8ypo9ynOnK0Hk3+qMjcMnQveAI4/8jXPV7EDUYl5H38PL1zWWDIOdX8qBb8wEHrxj
oOdM9rxesRzCMlPWoZ8eO0b1PlZRFevYxJHW85ZcNXE1LFPwMgAm3GEaa4c9YW3uq1qvBE+P9H1l
o2M+6uoDJ8De3vA0nCv5xdb6B49Evkmm9GZWm/jioSBBCo+SNQf0uoEEdjVQNvEFmPOCCHjUusSl
XxbhX+MhM8CXUvWH1zvwKf6h2Dn82K4TcqxhJkWeDRuI8jeik7Z3p7v+nRdlA+Qw8F8P3DGfctt8
dqQ0aAXbzuBu3vzduV1Laf+GeTwuf/gLRZPBbED9lOZeuKDbOOqQABjPLkVPd4PFW6IHwgRojppP
tJ2AcfKmvjJ8lmxyDHHd65SFn/JOMS4cHRYLHHcm3ijfmGnbrlL/pQDk6Aqgx6oURqV9HzY0dhq0
KIYuW8QoSEjKraut4cTZELgVLGTgfB4mEQvptaIg52cwa7MKxj92QwTlknNjvN38qt0dNQjSOYwL
t/gd1/F/Uip4HePeF/z4o4bpS4BGsfiqC5KVJXWehJFE88AKXjIaSWEuoATv2yn/Q4LVATSrQO6w
46G0aOMg2IwunAZ3ESVn6YBjSAh0MJkOYPsmwb8M1Orlvc/xEBAmrE49ZJfehw+ifKCSDn/DNBnI
ZgtA6vzUg7jDY75hCAQfJdW2CZYD9FQkNESqLG47pwiSiWqO2eLD0riYGwDB3q+fIQ6asEi8FGju
jvoKAPdQioppX3sJj8jYHsbnAN1w3nJA/TX/jX+RE/aAmsV+APcWxPiviUstd+sR1kFkpIuS4WDB
KEjBR8/fIUexokFDfTnixKHEylBPGxMIoxlUNLI8o0qS5rjrObbbDFcJRhabC/WjI0hDVCpMBDSY
njQwX+7XA/myL2d3HdvdPju5cK5d7x053oUcXn7XwA8uW/ZtxRsbSv+forFKJPrD/Uo9Oh4EppNa
JEgS+PhqBjPZOO9rHQ/3Yvo4SsNTam6jqSdiC/B8dBzUJfWSW6FJaM6M3k8NfZiWjLfuOVcq3YRo
F9m3navct76E/VaKtlLNVbygP9MGzi7R8cpe8wmnrpRGtwznKdCvD+mJsbRgkr8LC9l0ZirjkVqf
qq8O0ztGLmHzrOHFklTT6eG7GzxlBKnpOoCspRYyS72U9vPyEoLctw9EIwQOXjTfbkpAzdRqKv3B
kQUYcYjSSVg0ZMO78WCDRdTx1HqvbYAeMxzBSnP/WlApDBuHHrZy/gYo+dYAIRGPsWzueFS7mYC+
f9Lns3detyymF2HnWrdzZ6PK2JoLImi+0r4kpSva+lMkxYgMJpvBoVZo/tCk4xLBZxygp5M3fjFT
0US4SSFHfRnakyumohCMNvG9Q+msrclZtxnkF1TAy8Hjy/WF0VpsBrUIfwocslpROF+ehV3+/5zZ
tRfVKzyiZAt4SQjhl1OuRGbFo2jp/2nVoUObOPPLWpNPCrk6GF3xkQJnvrVLRPEdwuj/MBSc8iFO
9cmDXtlWMooWzb3rjSADoJLpiOgCOIRag/v2DbIXGjheseyjYZ/XeanJkx4BL/wnflzOaLwboZnI
1QbWr54k1472VQGxqR+QBfsWPDGz6E0OOoJWen41ArTCyjO1n+mcpUnJLR2QnwgJBcQP4yrsB8S6
CLovG9zOFvouktjHEfGkv7a4XaI5Pww71hagwahtxXZAHJu+iTFjmzyXssRuGf4TI+Jt//PXt2Mv
/ZBPSh3/CBWMf6Ae5eXYEHd4tjT5rTC/YXon1mt3Jj00/KzsRme90tHsRgrHbES1o4+ehzj9Z9NB
Z5KazllispRsD96DZifyomaFPWjZjqbVtSzYPeUJL5YRjXz6/YDI6PUdq7oaPtCy8rUmnvPh9P4u
G6dhmLXnlHLA8tdxZ8B0PkLJFWb/QzeUJQvt2zJ2NzV0J2q//t9CJ7i+4PWdfUIo9TNyhsoKRqoC
XwlD4PpOhmyG6bl5/Z9deQyOZ5/ZVETosH1AnEQaU++AQb1F//fpZfAZk84S7WNGTvJAsVsFGt2u
btrEnUxqds6Q1irQnDVTpdZNAipBYF0RdbHTPBFPOupbZ8Mf/5I4h8uk22otYczYhu+26apg+ALw
AO9uS5CkN9I0nELNSIX3Lc30PBx5IaZ49Wg4nhFlMTn8b8+Bp39SXIxOiXaQWpkl/2WWwwrfFR43
WgyxRTarvDBzW7EZnN58dMM89xZNApXstOC6W3FqKYqsYkEyxdJWEINXuE3eGRj1F+VBdcZIlsH5
haFHJTOdCfHCm1ioocBvPOFtO7d+Ckg7uwvpAHyk+EUMndwU6KyGDWoFYERJCT3ZfMYI7q+xJieo
5VWYle/dppfNWJoMQ35IEwOSRe0aUdcWCQ4LOFQDCryFvhPBPPQCXqFa5bBPiMHHMYFKtKm6jErE
rVlYyfX/+yphO7bii/Uy49KVjPSrvrxAb7m8oRC+FhVz8n7O5V2vvaUGpDRtiwjTiaasF77UQDsO
UszAB4z2MuEqW7x4uEcSchsAlsTp7X7wun0GI7ykuQ1Jer1xirGA6qHBq6R9LAgCBV2dKV6xvpLS
b6S/pZc22/mJCEhgW0m1NfMFVTCWit1xlnauwuTouLGuSJGXCqOEnFcoSg+QiIAlvhMzvQOVH72t
FH8Ha/I+D3ramnzg1tiO0VctL+s4zuM1G/rswRCaXFR6MYiB53540Gt375ccMBRjVmTj1+mUaXgy
X2S1hdVcyGXnK8oR+LGL8kCXG+1VnPhQaNywl9CiA5jqYR334gr0PLF7jqMFsEjA4mO74vLVwy3F
MC60u5y6ML1F2G/SW1bUGowAXZkrVMxNLO4ZIR3CAmEOxLMpfsh9M/o6u97LahpbagmltZzg/HET
/y5/6vyICfC3MlsjlNM8V/eL4/linhOA7anUsglo1pSNoayt78C4FQqTQqeLTgDyQDt/WPm4z/M5
7bzZl9Fe4m0ME862FmOHSqoXWovGAQaXw6y9mr7BdoBQchxYa7pH8zgLQ0MG4DIqdkLBWmzD0MMT
Mq3kvXLSztCiuGG7lWJKxixw0gmyh2HOD0hhmrPkNyM7PGMTQdFPvN+Lvx3j5dFX19cHOkUvHfx0
beYCHBpbxY2kgRfPwL3K885GwTnV97ESBcuG+Heg8axFseHtypVYSJsCT1/d/uc1X51fnCgyPld5
5z8n2LR1caTr5EQU4lpx47BCzp9td+R0svQKYu/rwHxKBM6Z3Mu4t+lSnF1UEoX57jQj7IaxGcbs
SYpfISkSCQD/t0K6IcYOPm/DfS8u15h9LIyF1WdlEPbNDAAhDQUfQJwsRxiopG7P0XPiKifp3jeD
5hjlWMy7T2LNYZYUwjhzL4TgAMGCex+LEMYk5j3twxpvRxf7jDIFjEeg6pbVb7z3NHu2LcA1yf+6
jaB5ARlDGfZbTbApMDC/fdqdO0fwWJsEcqbNMM5hUY0uN3Yz4cVaFDFh82W25L3cZSNH1JCcjdBM
v32/20uGhQ1SOp9y1S8ntVc7hFJvZ17G0+v4r3T74q0tAURg5arHZzXcPgkR0YuCXgCETOY90yVg
l5c1qaF6rm/InZEKWfOO+G9G9WOG1+/+P7fgtJaBb0Xfq7Fx/zHwPfg83Utf7R6xUCRqIttets8L
ULPWJBTyQhI3heVp5MnoSmrWLfDCwIkuR2ugmSl+roVB3LeICV5bouULkWlDh+WvPRwE9G9tYR5q
g6e/omavBmDPssJTuUyHmHRAwagMr+mlmpsbNlKlPpj8sVi46n8oKPIsTBsmKkXkUlOHfCXGbFNE
ZE2rdF2NQTmyymzY6+s+jD73DJIjgVSPtN2NTYeZfD9LDl9LPjphsj4vgX1LgJJI/N1bgIs2MYaz
oTQ6kY4s8CJ+XT+ezxGvpsEX7vsnk4dfCQCUOIb+/EYXBgt96oMM0I902Ko7DxUiv0a4qgrXAEpy
nSz4XImPzGv5DkkDnb5JMBvE3bgNHkwOlMFBUehaPp6qWCWme9Y64KeSNNjN0K8ED7s+aGSUgNlH
0ABm6PkcF09K9evLzk7/QYPwAm5slzOrwpiqx0wxZx+mVd1BRh67pJ1KBLwLVwUzoXa20DDavwjJ
r8bGeG7lGEynR2YP1PN7f0r+LaBbmjbLTEzQIMj4CzLOACDNY+k9kPGl4s8hg+yFEIMjJvtxpPRQ
esZkasYHPZ/xvKNrcxwpBUqGKbh+qVjcbe2iZcHrdW7IFA7KpS8yypqKXKY0RE3jz0QfdzHL/zhW
Coow+jhXxTLv6EmjlFKJtoqRna9BD5YO5MZxsfjErycxhrgOCav9rE0J4IqTToJqpe22w6UznnfX
WrqjipSBGVvdYuwsbnQIjYzGL0opxn8YnN6+x4F5+KS3cFXNLgrj6lyneNjr00G0iKJYjWI9hITE
K8Uivt1rwIhr9Z4Jc+m1jp2lByJGxZMquzJ68oq1y3FOCYKZDu+nhHDwOkrGysTjDrQyK8htXJ4Z
LIjw0jNlaOIVoi5IMpPgfXTvnXOMUPZS/p8xXhsjAobO9TTHLMJmQDFPspj1+VLFII/x5WQQnKek
66Z68PB8OSYbLZhq4+op8rTIcZizw7/sCdb2ZB+g/BRyb0B7yzVQ77472x/FsEeSR6B1Hz1ECB4A
Nm74wus4I+9rPi/YldV8T7fD/7op9+7NSP9aQg28QcdGw3wFoWIStBOGRZYyuRkFzshteb2OHeJy
Hh0UMU4lZNBtrGDSAplHJa7GiOiQBYBaCZYSm+1RxMMqz79pvdW5G60iHCwdEtPTDXWQAVLY0LU6
ZonmsiCvC7z+xEegSdBpXIvbX/XqmGUze0E8RagxI1TCXMcpUzf9RIyA5W/NznWLDf6GiOHZzeI2
g2ZjyH9k18IfZ2L0HN47lP0oQRspl1K2AfKINWsCwrpennD+au5U5/gsDuIRn905pOKgFbDHY0fP
TwnTjVaXdmEP2xYB/4MX39G0FUNf7mElChxO9IThzvz7x+PPpMU+hxHid+QBROFx1Cmhv73yoGgn
splYnG/iFnH85Q75UFUyx3gfhDkk/uh/PzOjS5keG45XTghYa/h9Z+/COK5Be029BzhvMDLf9L2x
s6/qgvjzDFBK7atZdkm1AY/YG5+QwnOsg7k7NCxBe3z8/ViEi7aswb5HuWkgkvc7KCQlujfTkuHw
gHKVlRBZBAsbZ0/z3ubqpwYKiaY980fgbuK3Bg85yODZeulLX81NsxygrmY4QMN2GmACx6mhAjxS
8Wbjgkj/w7XaMWHDPTkD8mqbD0DzBDdbrcvNoyYRsRj9VMJHspQNr/ynEqw8dwRdfSrNBhd3MrZ/
YNAIMdiRGUDjo+IxiAiPnZhW7jUaywEVAMk7sDJx0H3HLGpI+cVGvTSNJro/IT3osArhcN6I7Uw/
6fcQUySZwmn4shKxjprvpwBqfQMybmGSiDIOh+8mpxWvSVkVkKOqyD49jYNpussnLYD6POjHT5YM
ucBlhNn3qFSUyoHgqm3yiXc54zWErzIkMa3MUDj653rHTZhg71Xr8gsj4iZc0l0/BooIyKKkT3Bl
6yfRWIMa8rZ3ZonAKbA7xbXwUgal9Ob7qWF5MtL+lSTZ0wbiboGtjzjwyGOFtLHih7IIeqvtHHqq
xfH4TDIGaTjHjSNxerGnh3NtxqPmhMe5p6lf374+52e02QeOMfHVx2OHneSHZJGhK8oXS/In89V6
898VFKRKhnPTTxzgzPGDoVgRavL7/8B4NQbaF9Yt0r9nTLhGF/rjQcTdo+wgNvOn+zZviiWYujkp
NtJuuTzs1Mx/lXDimyXKQBHYHV6gIDlg3RZ4u0mL59VQkS4bVvB+3e9i88C6YXVxVNjpCjOTvZBs
bI7VYB03spHfwtDbEPfxGvIHuuuX5QT3wmBtgiRsTobvBLOa1ecvQ+YhvGj4k0ksLrBJ3Ei1NNM3
XTGQNGotdY+pcAXrfoK/98+5XGU6SWwI1zh2NqTT4f8bd/XIvK4uhcLhN41C4CfmR2BWATjca1pG
71GOaroyoiH21EeUh4qHS01BaNv++Ct3nDIEWf0+Un+Lloc8DBjA/0SrpElBrbhPZyuRvQZywjwe
n3pHc8VIf6AslYGXuaGJf2u2x6n6IFCKb05Xd/eEStrRuH/cBTh5lTWDB3Bfi6SYfO+nAHZO6HUc
TeBBY/+3v1lH+VIT5pDj/TYvG8hxhkeeA78WGH4BI9v/gvwIj42HVfHQqWkTXJatWX4DhMsnnIfg
PA00ejQDE167VTrbJXZHYBgq14hiOJ4wLxprH1fqUgbeWwycZdrccD/2+ia69KNrEn3yiYeQ3Kft
rLrxRuiX0adu1sTN3MrMGDozA7S64n5LerOyHFaj7XNlSvbkeG5CktrfDZ2NeJ0T2RU/w1mBgnLG
yn06RfVWMn64bbLpLCvZrVmeKT/DYFgqsHIM2alzq8aQAXI3+U5bXB9j1NQu5saqsaWav+MtfDC8
IWfMCbig9rHipWPmqtE8pft9E4WD9metc4nUvumaFsJqohSr7zpuBpswxMgXhxb9Z1Y0JWOhNSj7
8yR9DyhLu1vusNbWSg5ef9qV0CU9ncr2a1kqCk/ahjTYQIe0Bor//yaN8fd5c79zKsxf4UKo3g+J
hQ7aLpcHhubdft8MKgNHtFa8P/vVegfW+a5n4Agnp54IzM84vfswERwoSgW5FA7VWvbZO+PfCZ2b
Zi1g8f/MO7wlQ9o6RqQEkSjmpdBoJmS/BdaPVMc7EJdGMyIyhOZuTBYXkxIFmMgGoGtuZ3dS/O+q
rTKVImhfoazoXqWxCSHw3+TX6/ykMxfhvpj4Tf6qoV4/a6iP9odwolAnlSYUF5I35yjKLKClPs88
7ABS5hiIwIl/vCQmm10jQhjqLH+0IOqLWQ6JMB3dI/IpAbSfMGQ5J/Dd7LtxnIXs4sImKU/vG/6c
N6op5pG2BEMpj2DbWJwnvE4dEHiUIOITaCa/bPNFtqnUVayN/4LqgzLpDIubV+7kPOz4LsvY88Du
vDGJXqRL2PoBwnDN0cHKHNiRXa7WlyPgsXGRduLRr1n/eaV/X+aKt0w6o26gK65rouYZ1ZdoVqzu
klLiWttHdUuwkuTHpWKu932VXW+K00tsM1wFiaENGuzDfvd2Gd8Wr5aXQ4M3DacTVqMl2outp2eK
DyUUYC01BctOKE3Yz9jXMd7rsVfzi6FFgSYA90BCZSj/AYA0iAaoBqfBDhoOoI+CRwaUj9XxHfb1
6McL3JhH6VvUzlgWE14+Kqxpj+4zY5oClY/5UBCfjZMQc6DOQEwMmY+GOGYv6m9i9SUMHtJtNJe+
2JswRNkifE8zGsd2t5HiurdeydGgbgfW11B/sxQgQcDg7i29Mb4hYk5s1vscthOlUQB36N+1JPl3
AegbxHzK9xek0F99I4DfNk2jP+uAD62NidZqyHEUE8riPpmvCMSRaaCZpqmcF1gaIiVmANdMWfS6
QMltX9kO8FScM0kRI0MJo/FckCKvUJwsYE0qfnHsepYd8Irg2etjL0Hxh9vYgfw81p7v5KGkMXsJ
qgokMyQz4R2e1ru98r4jBijM49VNumacJ4cUfNv/QQ5u3bio3TiJX8Fodq6/bACMF5INXpX5Sly1
3DpG/uHlUDsO11ZnDDsD3KU2/LZhnZHiOQJQWM3YKWdo2uot9Z4JVUr4WYSI9yhQh7LYkBxbNHan
MnD1tFftqeBLr2zK9i5fzs/KFrv6sYYwmTb/56qqzGLv4bwbGMRXZTLMBBnfFeUVIp22UFu19MAE
TvUQ64A49ONYU4j+m9q+lzynJrOGzlJMRlpzNUIoGQW0vIjJecKl1l0vQfIRiiVCBjXmyuLnQfKk
HZCWbdMiJTjAnFRMnfSl/Ea1wAxdg8vj67V9UDylWL2Mm+tLHskyh8O+ZcopsawB31yl54bCYACI
YrdOGiUUKHXqdINvTTezY2lJEk5oRn97b4S6NZUIYJeIruizERAbavViY3bT+2ZwhLtffollKu3o
7IMj6kDareTk8HFfLVgaKLHvdVnbAmSTTu8W91WSIlwE/k/69clsuG0IHgaaZLYCtjfCPy++K3/e
JVEHGhMnPHSRYvpzaoMSUKHQ2LsFnpWxKKDI+eSyzO6wLRgKP3iDLDPVPukd/BXbI0NvwQuv6Z8k
iMl/V5KmxfMZxfdZrOpbZG4Bnu2fvrBCfgJejtKvj2+dBJauGE9I2pAvNGI8+3pemNx6yRPuIFm+
ueCrOcKr1+puFpxiNPdR2Sw1yWIe6gCQcIs5zFsdHI88t6MHoZ6RN02w7VidfMP0M4LJSc5yocl/
9VUeB82FZ7Ql8MW0zy9lEc+wahaTedJJnN6J3/efAwXJBXtRMO8ueIbjc7CzH2ABNHQjlx/cZvEZ
Q3Ht5kmQtexow8mqjB5SQ+29vV8jFf67EtUeE9uDYKbZplOURzo+YRdYXYUQdfUkWeZaG1d4CNOi
KZVZ216jnS4G63LHcLtNtXffJcgOodNeSFKXEWFKC4wUXhsZcAixIKy8Nx+h3ZhvIcNEaNf3/YUU
tMKxaLAf3QfYGzjkB+GbI5eIGJPxynhIilrdQ8exQPgT9UwVOpbC0gUNLhETH0uADJIE8Vrj4bl3
jA5NH8bG4bl/DVR2Bs/F9R9VjvN8moY681FxLd0Q8ToyVBG8TO7S8dtrzdgAEoq6jIcPoVpubIHR
xf2mWY1u6i9OrM/59AF1GqqWkyenh2blmxUBNU5Wm3DYo2WUGtBZbXGdOr0LRJ7KrPmMhiF6n20H
DmDbLTndmm9ZkOhJy6lHkg9+4vV0sx0g2hWHl1be79Po22F1OE69ZukFf+uu9EUhIxPQPFTgShrS
3rjqk6tjljPTjwtmcTmUv62IuIHVWdgynjYEeMqsQZ7ZIqAcT33nz/adWG3O8CREM6sH+3RGvcvV
k+DgcXeNJkn8x2cY0OcDoQQ4giUPtHZT0Gno7GsQscMFWv4fm2O5XRktn8IgsLu6u3lxpELJhGi0
kAcSScKQ3+UBUzqrGtWdMzSYXVQYlSQdzSvtxihFVi6rYGwC0q/bMddoetWZ5NYpnWgx9hKPgrdF
4PdgYxGsZkioLnMOcOcX/6U1NA+ecXv6547Cvw6Wb0axlasb6XdOgSzpDR6H32y2txu23wAYeSRa
oZ5FcjipwKK8LIIzfiXzm/FHfganBzhZXHWyw5G3q6Eajp2aBhtnMo5OPo5PDBtnQ7USOSEGN1gX
87NKzHmbLjnBMo0OeDNW1Y4AW2SnC/59wsXYApeEblaAqxCMyzpuJysOGVvnkRDA5RmYN1+mc/xZ
9UppwmegDzkvkpi19d6ECnmUcCpI+6YhGmNb62tAph+LBuxxqYoGEXd4xiloqlkLjAZEB8w2N0zl
g2XU9cqVeUwupbd8ZSRXYsRQlCc+v4mbVZZ+N+6k8fISH61KRSFqLlJUIh0Nnw+HQWRuqmFDc/1+
hsDt1mqpBXTaz9+03AT6oCq7JhIygFK1g++DWcEC0npQj6wmIB4gYpzD8iMN7A2A2P0iQYKOffmf
k7LbAQsu0yZOq22RWHOxvpodCWEOAi4TGxFcnH3Yz9mvNuloFRnlDHgpcAdcz/P2cOM4gpJQFTh2
AhExz7adzBGcMv/aDIl7g23iLmg6Jli1oaIZA/bm85ixt4NPZ97befhitltHlSB85P4PycrAsOgG
6aYqFKJUUnfNdLq8a9NrjYCSy+yELgK1vM8tG9I2Jvd2Bii+hXZKQTGEY9LRt/1lJygoyBx1d6A4
Xd5mGiXl3VeFE5mHCUpZIk30HsfvHWGtA+lsTltD+tN1h/uj9/M+5jvTihJNbMbVjmBlv4SY06pz
j+T7J3d6SWIZsUJKlkNq8bHQsjCX3VCv7R/o2ura1LiWt8h3lhlqGw8ifDXAB08eDpfC87b+MRS9
BsSgUoW3/FmofQM4P+evKRhmU/jdiS2SvigbHmtkuzvlPWhEkfgZXm72otXMh5OftYzGWxhTcGxo
URoc/89o1hSUwmSfSKbpcrhLsw49guQ7g2QxRWjfGc72+7h/QTvVO21UAQMQhsFqmbGl4taw1IVL
LO2ltMWCc7IJYXKzFvKK36ddxtL49PRMk7BpZh/locuUnn6DKcXlbq/eOtwLtsD5XMDvmCPaKKjU
fW7bjQ5fIx1oXCAQggxpixTb7ydpwh+anClA0vglQ8wmUoDpHwvcMIDE0gIch6bHO+km3Q2mFgKt
9WV96Q8G7e535EA3U7mF1dmgM1R/OP1zeZJ22lEC+m4Gz3d3NuCm5G+qngkhNZkElAT2NM5/zSjY
f+bBABS9F/8JxncebQh+q2+HL3/Yp220TH/e3fgb8iXrDVgvcg93mSQhHf51wvs4zwK4Vbl8BJ6z
YV2lY4I5vd7kfOvrPW/k4UWGcb1xD8n/1KleNynzhgnhPYNiZKOsIkVWle7f1Tqrq8piWjKngC2P
wquSFuRg67GxFEPwZg8XyBBMhoIsX9HmYQU5UJ1RFWIM+WKFXPuy6YXVJWVZfButlDHppFRb0U1p
iwg1kniRiS118IUStWC3oehYloehyzg0kDeMtdzicsMWD9v77c3j2uo/LSJPCIKaDhW7lNzL8q5r
lqV1lS9NgUNEBsERN/H4MnOc3BHBympMabiJp7tT2xkqDRwgzAL7MXDcgYdpctdiRmJqJSHn5x4b
DjztjTvnOMHCwpSi0kOpAuADm2fJQcZMEJZOiSYxDdyNpI1E3CvCohsDcKhtwSgkIob32cdP80HC
OrwCwD7ku+Sywp3REf4Mtpj+E3I/F1hC7eXqHcQLGavR1ZiuOZWmwdbJfu0hKv0Ym2Tm23BfIq9I
X9pkHXu8MNb6vpWjtAzZxzV2w4dXV0QIkQwVrOqAHGBedWjIbozEK6nLWV7FoGezBTDTdkRTSCZB
S3+jtSxWNHg/NEQ5TKYaQn7azTtcSJHqfPxl93k3RVITet15dtBlihYL4Nh2oGTsY8SWr5Y172Kb
npyK+JGrHHqG0J/wPLf7WuPaQUQm7XeSOk4VqNoLiNrnXdPqFvfwMVswEHVCNGV1oYK+PfVthgAZ
jLDAYmwlBnqSIeG4sIKkdwbccZKSpZlcEKL23p5xoc6vXTy6EMF9RlwdCvcGYSGeWUyJWQk1Wfsm
lj/8oh3kiWZgXrmIn14n0L3CeDIM2RtiKSg+zrZERUJcGu6zwJwNugzbMBf0XeXwA1UiKwZ0bw/u
SlHe2zQf2KUI7qdmDA3p11+0Y8CgCKji+V4HSZAeFwB3LSWnNMBsNqkfD/pof/IbCkIY5xYCbizz
zxJf652iX0KsLIqGqgf6Ew1x5KCodg0/v4SFnTf2gDDiyqIGexDLDJwpVQ2U1miBetFWXEwzOuGw
roT1zOnfgZFz7d3MHFOTMlI8mc4+nwf3UfqsAbsJc84NS3dB/A6o9/qoIs0wz2fetTKQqYHD0aD2
+VElPKlERQaKnt1etRptaYwN/BUF6HGvhqYvf+zg81yPq5nE1aDsDzLy4KfaM1DRlik9m2kwZKcD
iBfVRdY+uGYexKuhIKCybEyL7efeTuRxiHDXXSKzGnaAQ2wsBkKKCi0WDJUmMiwVkApgskLS414D
ogJCFPJWs6w7EztVkwBlbrXHTU2qc0kQFaVvOvia+bgASM6Fbkwy8XNsoFctyHsJPFHHC+Qwg6kl
l4J1Xa9P6KbReLyv8V64MpfnlYsQoStBT1ZgF8t6q7czXR3U/xe3wPD6sJ+wwkpE/c8TvnmG2I9X
Wvkcs1EX0EDyQ2UCyjo0wqrhSMwEZN5t2WWJIlkNw7+PJGTJyM+aHnoqLCTYDnU5wv3NvukT/9Os
M2DWgZQl13cUmNtRbJEsj0l/ABtTQM2W+rxKfjd5dzcaTqLaXUvzg3SgJfOHfzvNQ9fKvC8Bxn8E
gQACNd+ve8ZEYKayT9DlLKAxQMMuCzTNGS1wDn4J0oAFDgxX0KzW9VijcqQefaNISg3nUHlOv/KE
TlgUW7B3gvdTgTijKxIrMjb80mprNpwIEeIaOXZqcF8zUy2+YjAHu6iTCQgny1Wds+Y8HXVOFOUy
TdQjQgieDNV85XvMKM/00nrNEnnciGGL7gBkwclgNIaEoO3c3A3GMJZMqVSV77/qH5lTLywqeYmf
pKWEYvRbBGLeLBAh8epaP8RDM4UQD8slCu1SwNPz/cNpw/zXtteVL1dYVcMhFFAnDrdLt24ZYsFO
NAa4Qyvb7lHjkFGpf/t+IiiQ6tlogEtFFQoveWPg1ptyPA6dn/2HshOvVtvi2KkBcQNsNCSuWOcf
u8zH4tjB+DRcKe9IZVVRDYhAxnMbfnHAvQBTYB4wcBL0OLXjH8Fqdf5vTYcPZWOuK7jd9R7jsbCv
m6J6H7DS4OLqJw+HY6qv/ErBFZQibpOqsvWvONIug4nSqaEs72jEDNnR5PBZ27pMlPW+4SieUZvn
LOhJczmdhx+Z04BHi5zxpPNwxY1YvvqF8gG34qmCLdwQ179dMjH86JAFeMtVs5UHryvYxs/Uf4uN
B1vXp92a3wMSZ3QwV87YW3H9s7xur5ZnNteqBnyUl5lmSnipDO83EPRLlDnfChB3OpmwGhBlINe+
zX3gI/pXRvX8+IYFqxI9Gg0reUkbqig/JauKF0EF7QBgLS/IYESscFj2HQuKZuo52nzNzy/UidEw
mo2dQZQIBobT94HiOEYA/We11CjtZYmL1RLzOqx1I2Pjf0/wNUvOsxfcnjNBNjeB+njoB2pTR8HM
rvvDPPt8m0HwYA+AMYQCaiY58V4NgTItCZv/7lPSEWoMM5gsEJXSNM64RfgpYVhH7BfHGwd74cpC
KZ+oaq+LYINGHjsnrWefGlNoE8fIxxo/8zaAzXH1Rrit4AeTXF0LT4N0vX2GE2blHk0I7NtWvQnf
W1O+rITk+m+uyEtYcLlBy/scF8WaIb3RXJHVSyrVVVTaO9TusZ6QSjq8rlQ3axwTn/GIxyyEK+tq
AhSkuEkYW2/2RVY6LNUUX1O39xOdGzgQSRJcpXGGzoO43s1j+xgnVOKPZq6TB3H06v6sKbYVzZpe
AeOr21izhOd823yKIHO6YqmONwp2ZJ3lZ0VqSBSUV3EKGNjNLNXAvnuaDWHTbaHFv3eNq9soxchY
IGve7rTN9En6ngXThIfTMOZq5jdl755frP3aeibhsmSb4UMnZyol3+0+/rzOAyfPhFm8Vfhkfql2
kOnLC9pS/X9maDqGmJ2rcZTe32k0ocbbKUF1B8B7p9yN0f5XuVlyKji6Kn5op0nl8Dqddz8WoZHa
LCF5sSRhwaZ0zlVRbmOVngPu7yWpe5Yu9vRVPmisnvi6mnCuazFKpqLu4A+bazNBVZonaFVNdI3J
RspzEFBjTkHkzts7BwpBBZDwazVZ7saClrdHQQxwh06GIg9QQCcNe/w9y8Rgzf8LNJWgD4bp5VCF
hmCWtjSYgpaXP+kUluqE3O7u7kohsxhYQfiDRgmL5EsRKeguOEobXqdYsuJMiKn8PwsBBalsHSsR
L2ODZLSTiIxQn3bhzfZBzpBj7dgopOqTwpFZsIz8Yv+URt1/HqutISWhZAmFyp7qDek/bhOZGAkD
qMHLp1VUx8yGdrju+nsTk73wKAUw36HRHcsfkWGfeup0OEn8zltUFRHhzwDtmG6GEeLumELgHmPj
fJWxkx4A0q7HyDPfYBrkUEHkbOsk4TVhlG3kqEyzXsWPYHxZ9ZgDQ3AaOGNL/frqoJb4UhLwEaR5
SqUTNsvsItVU13Aibi2qbYhaO4d+EhI4HrwP4lFH9DTdnpDJGBTA9Yox6dBjfaOulzaWjBM/m/vO
xfch80lMSQSnwlI32mZzkapRBVCxtRkbHrWCgmxPaxcOM6FJbYICOtKZIMuDD6H4gnDeKQPoFSXQ
xDYUACRKX5nTDtLo5QtMCbUzuySus63y5vl3Jcz2wScuoM4dVtLQfizcfwv/W64DyLlVrvJWrE+O
jS41NtNlcqbhfsCMo8nw6y4PQFOvCUGZSbqvevlnmcU02YVi3+ILZL3E27pEKtjbeo4wTyqPeqGH
eZTc41KjWRpFs1FE1ZFqMg1ztoQzDbWiTqFFyPXFAIQgRndBYlzlJA2oy4gX82FrAiD4sEYQcAqr
GDthoDW7rpRW0po/xhq4E+otHvnWKQTHxCTSxwFfgjQLSapu/esCtIjGT/PvvUwM9NIe3VS2ypew
XeVedn+bdPhVFabUblBcsbJRBhoG/z3Em0K8sg6fqbQajoi4MiVsn8H9MGKhRcJzCJe0ig19uO1B
2/jriK3Zy5j1bhuTEVQ2B1nzDKiCbdVFZg+HMJsJq1aR7jkoYTzMMyqMWVA9Dfs3AOu0A36P1deg
fSZzf3qZQUxoYBML8fulTetdkZ8FSt/fH1SpeoJOnAgi1hfd6DLA/f2+upaxofpX7cEsQok1KbcD
exylu7tKQibB5YlVCi4QG44QcCrtx0UZ4hpttGjIgySV/ZhhjjkmUtdjhetTImm+LbQbaBx4gf/g
fNSQWMOjpoM5wx0YFas1CokId4npfmaNXnflF/6ihqVUPEqd541HCVmKLFZHykJ4v4klc4fgdBrz
kXDeW25g1FBsydeywAgWcTDhSq0SZilFEpvoc+R7j9FhNOb8e+CtgfibWm3rNc3xjja/Lqu6aM5f
bB+Eevcsa4diBp0uZgrV7seZTSXbG6ib4+yftLNGoxJ7DUFE5VdzL5XuHobcMQ9qvHbILSEiIHF1
7b2tYQKMiMkXSTYEsWqPRWze3ZvHKaLCRivZXNJeITmKhz4lhZ70HFYpwCxDdJcZGPIB5NWeK1jp
pteTj+U07kztJ0YYL8AbkZxO+PhXU5SFSzagGDqMeO9BK37dW/XSxb/usZ504ap1ZH8D08wPgRp7
nJ94Gv6Knl0sYBdbnUQvwlp9CV0b5igx8Zrl229W/CQliPD9NR2+SUzskBlOCkDaiqog6GQj3GqP
/0vyNImMGTAjeiyl9lpGQRDJgMJEjm77fHUuVjnLNaXMWRyl2jd4sF90f+AB50SXqF58E3SVPT8O
468y+yQPI5D2yS1qXRW6txWyutYU8KgHCTzj5akGTCCY1eXscmffi4sx5pVKpUBY6vw11hk8Q2GK
oc1cftqpfJTC6fWPz0NQkOm0HnAN/0d71jxjRAVmh+h/0NwBmLRS/+PvWO2RgjDnTvjfA1e8V0NF
+8AVfp/NXA4+0mFvR5hsh9boGS7yNYbv7DiGm8i2b/sAPyL6xlbbTcImydOkeSZevs1n9QoOkkQq
7PKxDrtaG/pK7GqdBu4bZ1PbxVF5HkOjYuqSyTKq7UR+RzX4nA+u2A+mGfEUyAAwECWO3AOxQLbi
YTeAwXCKPvWzDXAzZVTn8DP5LgUvMRiHxQr3NcV3c70DMxP0RJxrdufkC6IP6NeXL8w/vnD8TkbL
rGrrStLaqPo6A4evgl7Ayueu6icXNdhZ8BiyZT9pUiLAmdsNtsO50oDZa4QUmpih5Dr4MrNXWwrM
MuqxhwRZjQ0cDp2pLNvquGV1FPpBCJ7IBZnhxX5jIUKV+xqVQYiRn/DrfCmGCIyMSyqSJ5ABZycC
Xcerxcem6GiKvKIIjl9aOlKGawnQ5N1hm+Suo7D/TtyUBsBnWscxsjmkk+rByn5vXWK34FhlaD/J
Ii3u7YaAX6NJktxpa70OHYjd0douuIAWom+jpCMbg7UIMlQIwAtoje8Gqn3k25lcEn9KMwNWdSj6
pCTrqPMaGhD8mvdmoNbllAsBPR+dWJrByIky8CUSwUP2uojF3JfZPbZbJLC2wPoW49aL/C2h13T1
0kT/VNtaVhXtttqjebH7gdk3uB7UjaFExmLAyDh++12vd2FYGXUkYrqgV1diQZtF1olU8/UPYYgU
+0rc9JbPLhNpji4Wp3aYRbT10KSzAjWm3flmoL+B1Q1S7DOKsPEm7+p9MHmJys9AsL2w9KiLe9Es
2uszDgbIo7jxlojZKLP77+GlI0pHgcGDKDSKGd7Qve62izY0gUFP97bnerRDeyrTVtiVXMKnuL5n
HHTd5QJEIElPw8tww+aDbOLmz3Q9CgQqnkIMrFcMx6UhpD9smcXsb67w2VZxil7YsZjmN6uVb3N0
6ahSPSp/JI3lun1oRjRKpoL1/p0CyuRVcAZLpv/sTockkeYw9VRirt0iwhyJV+QfkMx0lFhiUFbQ
I2l+z0E+5w42jL8LjmZumJ9MGxhtFT610M3YWNNzkpwlsLq24CRtYPTiOBZP0CdHwwLh5vXAhHlf
vfA913olVqCaCMKnSaidM0R4p/JidMcNmLEdojgpMBbuUbMiCXLB9QgzOw9dVg2ajtjxjI7CrIGl
+vylhqPSD8MhcpdjfvJi11ZYBAlmNZMPXY54lfzc+RAQoiabORRh+0tCwF2BIDSR2AKRFqnfe+eg
4kvujNcrh269t5zgZKISR+FJ6jeG4DqkVq5ITem4UxMGIdgHvOxWhl5/AICn1BLhwwsQkOfRDWI4
6rmThCQp2S1b7ieBUlNw1UDilkk0u8hOgvNyHue7blvxycdf1h1e4MKTQgZ/yXdC/Z/WjzqgFLtX
JI1W10u+WIUc6F//BuEsI3mRYKw0kTExejdHsPkt06CrL675AA9xHbSrZrr1GgXArCq2Ir2hSkPo
rZLFwFPrHqa1XA/nSiOrWB5l4xvfC5xc4XvoRkilqUARBie/fbLQdsMLbKMAkd2k5PTVW6IyNzt5
fWKDjPKJ2Xj/o8tDaUOtgGBpGavxqgoZSglaL/r+lcVqIZF0iuIgoeOrReGzbShuaJJzZf8f3p3s
KFiih70OjC3XikyE+Eu0E/4xLkpySImbnBlFy6F3d0ocGNNqH2Is3voUaEt9O7e7AFk/HnAFh6nE
hkqQX43FcwBlxWdWurf+0lVOTvgvJ61iBmxEB5WvPCU66QSoBUVKMWwf3OE028g0JzY8QSdpYNWF
fO8mOt7Gz0NC+AYmAkPZGodwE0W4J81FYLPJa4i6qGGkG4UftnLdC0xYhrkAV35LLN2xQxWiQIBG
PVmcVoOEO37LXzbJKXp+O/oa/PlV1vw33wGKWKpAoc4CO02lRVE/IwAbHjJXjaOUlDbZ20cIlv4b
p2wGHIXrb1owtmi50Fy00DUH92ZCjyDprWKCWk6iTHCkz6OKJQs3w2nizoSFMA4G+MfErS9YTFw+
zh28FQ4S8laPvPQVoNcTUUSpdzntDqcakCcLX7u6fhH84Lz2XSgf9fa/7Do2OnffW2X/8gurSMlA
E0r/qBndLq77j/59t0889l+TP2NZeX0/nPejyQ3UlDFJejMvZtmj4s6nYYhEPklBoX3TDTW2wWAX
uiU6jJPXj1sV/bz8DuT3Bz6QZR4b11vgYQnN4Bh+oylYhx+T2Dx7XsWcxZaw102G1JLk2VtioBDE
umCTcVfay6fXDKRH2IX0vAT8+B++hC1lf/9wM1tPlKxt6kvuHubYYZ7y8arolrW+EtF7/FtX9S4+
zq3l7IFba/tVDYsuk6bu4xKJslXNz6u7MQGyOm0RGdB5PCEp1VFWkBUWu8GBjZjd5QlsUEhWGupz
aWz3UHgPZDuajmDhi/l1ZawYqd1RhQtrz5XJ9gBz2fveRu1FHKSlGn+qzLgwgoAoQT9uOf4oILzC
ZMDLF1b8nM9aByit4u7+1mBwABxbiHH+8/q2npO3tpMBDKCsn5QY5farAFF3nbbWfyfU9NT0PfoC
3vC56IbMGags/51MzLj7IL2I6Rcx1j48QKWdfX04OHYuB9ABDHVWGybW19BUf+ThoUnhoSV8+WqU
79AmaDbLuhqFPnBupoA5IGgqLUQKz2JzHARTdjxCDFk6/tglQGXrYHmmr5FWtPf+OgMa+J9TqppS
bGYr0G1PMAefn8kFJ1TUwpvJuf5xIjX2D6ZT6PjkF/FEHcaX4AqYlJZYAzBxWd/xunZS/yFNMO6Y
j4xMLDj5+zYkwLKImRQmZEHdsFjuMuQfaUmXdTduGN9ml62GkuCNJoiy4/Qvgf2S5x8RZV2ZscbZ
5CKMWbZqhFrcEpAnoJu4Ugh855/xplCQ+0fv0Rg2j7jJ3vmm5BMKRKVrv4GSpK8TRrfBDbF2BogS
+KFyGAHMNofDSZ++1yVqe3tDuCb1V+e7E0Ty/cSBV4+pE2DUt3JkHALqZbt/3h3ajGx8MpRddYdA
w3ztkaNeU4diFxxFgLCw89ol9PxLqj8d02DHQLN4ncHoYq/ivoEzN+tS5PibaaRLh7AZ1+JTE9RL
JpQ+/TH3OuhMDvemI4/6ISOUOQECEKWRdx0sskdJkZlTdh5SKCzzXK8wMNIGGCFam26wzWmvUGW6
WSPhiIB2Fp4mMBMW72NFmy1zDumCAxYWA9uQxrDfBeC6RU806L4zLrfuydstxDm3JqppjpVJB+jB
xjJCZqoYqbFj2mIWhnKS/tcUKiH+4cHhl4PmPoFqpdRCG3MmYbWXJ2XGublxYCUAX5BPWku9PBik
h9s8KnGlMwvOhZ7svTwAO6S/U+sZ69E4t3VphFqIvHzAVB4G0cXj8RVPGJvmnZ4nsjjhsvXv5X2B
tfVoi5jl9P8aWu53Aa9tALIFrBuSCWR7MC5Fy8rUTaxXETe4KgIY0QQYFAxXq2hS4blLy9ev2cog
9Syags9BfN9DM1KqY+PG5yLFiHDzw/foo1f/viGDxFQ4id4NrnAo6iWtGEjBozQRTlB5WWBy6bLx
H/05fEnn2FFJ3t27zgzhAGSgioQtNb+sZ4PqG0ncnBZ7hvm7oQC47pm9TpW9i8gJHuq0Pyk64UtY
0huBThKprtkkPMeOflPKsoe8qUNyz7MeVXKlNNAohwkSnIMoYpcJLlbDyw5Ci6DZtkccQJKTPycf
qsWTtyll+5mEfTIXnaRlk6GzI0kARW6SpH5MZK0WzI73CBPBQZ4lxp3kcIEkFHXYDTH0jwEvEI0D
7eM2Iwp+S0QOfz5Bh6A9Z001VgbPVIEitn4E78DpG+mDEmsu7r256q7/24WEdpldRAelxvP9rT6P
7mQoLjRrdaRp54OGf4cU/hnWgMhbhIpkw7ngi/xkuLTjiffX1vcHGH989OpOLmoBQe8KckhtO3Kh
IDr6Z2/k7DnhpZB/GLML3AjE/r09ZmjM83IPctmXKRnuabPYrfGuKtj5rCQLhkk4a9qGt9jS8ljR
T36ohaGhNCLdLpsJVaNbpNPBR5hW9fd1aDmHKS2vdomeEQNpqv+uGbP31d6+V0UohgZUqGiK2NIV
TDSIYF19YIDZzLh4SSPhFBlXpPSqPb2ejVZXMA6PeBeeFldPG0hsCW37zPW47VQNDcZIJIopMg8R
IGUGSheV+9hY/EG2WcMNSGwuAPEYkVEf+uhcyKaBhF/txF2nnvCdQyOEGGr3uYB2m9VUJCcf7++h
2K1/yCYo4ZF3KX/+QwP1ccOE1Ze4HxDVK8+usMZu6LjvEu/+cG7zrOnbQaLRtPQs1NCZjtA7PZN7
d9ILXbX9WnwKEgsrFy646JC0hyjVnT9AzMAh7IZBZmHsmAekx8KhbozlyvElSriLY1O25GrTiZFC
PFOsRnl8rqGUqgGFZBIpwmZABk2EO9X4Mipv3RO1MXQWKE7oI2n6ESuL0yPjEcM/EfjYaKJPR7d6
wX7zHykwfQifsiauZ5aRclzNArj7P35I/77yxjcI5mE39gdT8RgumwzdXa2lxwe/6w6Rna0i16Cu
rf5MWgkBc+UAaHBfNszGQ8H3eCrbNYYM0UUq0AbsXmwwlb//y3d0/kDe8S6fD7EEy91UZnlOm6PE
XV4A1StD8Wd2opjc9f+WfUQUtTWBLV+iUQDPNmgnZOTZHcSC0u7w94DiUjQccANKwijxZK/Q4B+9
JMWs3c1iYk6/cs+vtyEOrlpjvaUIp2M0yTcvTACqClnxLQYG592wMul9tCnKKEREiniKyYMNwqH5
XIYRnqCj1jFhghn2ErYrJxzf9eRe0DXdvthzKMaWi5SeDbAlWOc6sr5KeXPjgYj0o3QSRL9XIZ32
v1OuSc+5hDAGD3WbvHMIbwZ/0hZr52bbG0xQIgDVkmtIuuhgr3+iuSterhOVT8pxRsLVs0I5Amtj
guL4Hf7ccCxCnhZrJUTAHgGRZocb14FW5cl4WbbshyJcZLZYafTOe6zu/VVT0WlnWxUCoZ0WvHwv
IXnXZ4+bIBl3IaCTwAY/+rLemQpJOwDLnGJ+Ah9GW1lpNoElAt28/y8vfGZSm94eG0xHRWkC2RKg
KSgYeYrf9C7jfF4JLpMsnrMs7us3Vp/8mqSX3hTHxGEMyAzNt2+oSPAz9exCsBqCgzQHDwQpxGOR
YofFu7UgRS3xSbxXNMNZlmuZL2sqahBwFeGvIgdUkwLdyawzUPt8uH3YFX6QGWgI5zVr+mfPxb/I
tpr6xygWx8SQkTTDvWsL53aa/7dE6zd96PZtO258w1KN7KBNzDdukOCnegwQ/3z2x2HBVPIKvvxb
3cFbpasPvbSKsjLKPATIE6ygYBu3ciD+oRTIqKpkbC0fIOjeMmbT14NFV+OG6wRbmf/kkDoCURHy
hgmJl//wgG/DtiygpQyUPU1Rk0cyaiHPIHv7/TPaTVvhxHdi/dA/HpmW43afPq/TLvaBxBY22JmL
EHln16Tky/WzA2ZXm6igjpNGFXl3kvTgcC8hGSyGbva9bXangw2WgAL+vCPlzhkZlDjFMqh42R5F
UZaCN+G+ccwxzA6WdfJx/0R5Q/YNbAPSSh7xjc9HkvQK6UwE2z4r8N9x0GvEi4cCNxcCQmtsmDRI
6YmQ+moe4mv52xGvnjM6rFrCl3knOqj3mWmzP0zz2rlImUztA3CXc2FG3ar9qO76KH03wQGaJdXH
XWcB94HERLZiCdP8SLNkArty9HNohGXRaIPalNhTHXYRlhdA1904TCfYh41kFNLnrzgZb49n8zsp
vwdBFepr10zZYxuLJJ+fBqqlC5V2jzOmvDc2gzQnAvOkSYH/m/vyTOrCa8bSo2q+AmeQZo7901tj
4Eq6hH52uV2+fAzXJZdjjvaYxjPukvnZfN7GQT/1lwbcyRqWmIrDpAuAVKxryJAzpqN52PUDP6p7
3i9KcDj1rL/G6qOzAc44eS7XJedrVVELz83+7dUKki8hKYWx4fx1G8ENoXWxfjO/eTYG09qVnG5A
tdqcf2BvPC+7bn9nyHS2BlTB2YO1uioCFzL4prriImp0943LMjXGP5sVoKI2LSO9IUBeLqQCW+/D
gdrgv6MXvouCcHeoAk2OWNDsAcDl2JWvJjC7O31lxt7W2ojeU6b/es22XLPI21w5EuWaADgUv4Nj
t5Vf6vu9DgsE1fEBc5bQsCYb4H2VdCMFT0AKY4kv7DpsAXt7JjHlg/1vAO19d5+ufhRBkLcCJpH7
E4rCD0ShnzZHTHaWOhUnDq9/9Gmq+Ny+hi1fP5tuQIWWgN3KTYv1cDXjRCywon+QtCST6cazDBla
xhgyMumCPO/Hz5p7rvdPmdtKFonUWBPX6QD/lrsyM9zwgVsMCWvf5ZswCDxNwTNws+2F3bXzNtIv
xnNOGura4I0PrUqOosiq9SZRPQuAJzju66GY+hV4YbF+FvsEfRf+pRhvTslLdzeudo/hGZOcQrvW
JwJSNaYWjofPPTSSjyixFrAah00/SoLC+eSB1uYAKy2EfRFqipr2R/rHNqOmX+d9MNjCvxZwRsS7
r4Dd7uZ/5o0VO1vwsItl54zrQAcRfmCZztTJILMjvwY2dhcJd4umI/Q5KCvnLJGpE+SBJfQvUeDp
b0RmXRGS026NKb+9Dmf8aNshba/gV2SmWZoumuxz6riP/66fwG8JAnbWprfL2mpBQwSgps4pM7XX
3LLcYdEWsiukuw2qve+2pEKEX3QGoTDoz+vOtz0VWtrhkkTO5c11WgCHg5qI1JRDiIQdzwlg302W
E03XFzXd4tqDVD1+Bz8FIjKZBRCKbotKGQ5fg6fBGkz8ip2fV+LBp6yEt71up9hNb7QolKEWvCaV
BmjGJtJGB77BqMcKJFrgayWWxJlthdm7W3SHseZLZUcljTPduSR6v/0FBZW7RX/mc9RevPTpKvWu
OkE3Pgada56O2X2+I4oaK8o0GTG1S3Zdz7DgUFdwT+oQ3LcqiqTFWes8oRch3piYVhFMDKqiJeFz
E7XvmBQsx0jAQGBBsQP6ldRHLCVLc2BYOywFIV/hzosCvbd7wlVNxy56UT7MIYljB6zILF3t+xZr
XxYdObALR7Gt6Z/qVEtUkBhIapsT5JjC68Qc528iGWW76tl2tWvQHeGfpXpg+XDqrfFX8/OOBHLK
jB2G0fKZvf1g/pCgc1VppLBnQuxJidIyBvntWX7qpw/Q9r911r6jFbE7ls2j587p+FOyaoP3uLAW
dB5JpAQfb7QKqc5HlxCjlaqqQ6S4W3/3LKuNZ9c/4F673g0f5R18BqN0n6O7fD/ljGVcm/6wRkVN
uKu+IAnIEEXkZ5s5jkbVCROak2ZlzJ/x9RU0j8ogdIhcjt6iJSFIxrS3ce68HtrfmR43eIUAyvdx
sq9K97GzkVfJdz66BiPhoxVQ3TlmnoiucHb/N7K4B58HBa7N9bIFjR7AmNDwKwTTkfiiATq+FG8U
MaVezfVRb3CY6ZlN2t8TrOxhAqoPHdDZ8dDbwZJGxjOGvFF4Wl1EWydLxCiNTX9vKEHFQzgpw2sL
Ef48e8zHMkB3DcpsKRKDhWz3nzPd2O+15zZZGahZzGANj+s6QazA7hoc6IMqvd8eegSyzKj8pZ4U
HnNRuJQ2wlcy4iQgDd8D+2WPd/fUz+LKwKajDNcViY77c4dYgxgegkZ5d0jD3izw8y0nlFRk4kuT
9pWcOg4yVqpe6qSqzDWH4QAAMQdPA3C0GYzJvDeGN9SgLkRdR6Obg+JMhBplVYmRScX9K1ATItj6
8OYqqMbDYmqilqjGQTanqnfbJzIOFzjONvgVQ4kKVfRLC5crDkZlKZJsCrs8WSOmZZ1LkjBKqyED
HstYhbUpDx9W/JclS21Tly8+yzXrljgXwVH1A1V3yZXy/Y5bdz/3xSmlF/+jD/fM7SECI2o9v1bD
wuf+3ed7s54wxb/G2DSJYdzX9z2OURquEzOTqJBfX6x48jML1g2kbdd7vXRmp3ho7/XXBPuFlKOy
nHRsgtDBvYmzEkIVB7ajVUbPhFe9Dyc15FfRnHpWjWub8si36oSGKMMthjEQL7MGaK7zVcNwg/UU
suHyce0Sm12wqeD9wKKfen6/+ouEAv4L7Kd0Y0KTDRBBCXVBWZUr3AJ41Vh+XfWVDoyC6J6jsCy+
64lP2V57In/MXG5rdRI384seN5/1HDGMSzd7HMaztZVoPsIYP+YZziwtc2Sv9Ixp6Gmb6cmBhjXc
sNA5B4v+TFVXkshiGo6lBkznUWLML3mhjVhCN13mmIRV1rPjYzOmHXpN4ST9dBc7EqScOaSZ1MEe
FHF/kfoqGRm4KrFwRBFMVeML1wOqXGtKFTm02VRaV0OOHRU3tZyZ5oQbGoNrQqewEwRbbadmVgqD
Ke8Xc/zpLpqnjEoTEleV6fTsLeZVOfRGVZNSny7zGCtK4EZdxlCXG37JkL/JLZK73RGOB9K0vkeg
MrTiinpegiT6fBHw6VfvRnpKs4k277/ZJQOhC4lgxaWo2UyFqCKmq77izJMBuWjvM8DUhTMbrR7E
ApF2WVucL8NZxa5WdUS64ZrAhdVnM8pxEMO9zwieMD1kJ5cPyq+pRZq8FuQxwutLpLFwRNGFiRYQ
Le1PrDE+E5Q2DfjG8uwj//dPi08RqLT2m9KO1Wnu/rcq86qPW4BfRLUd/J6XZmsNiKxqvu5+RD/4
FdIswwF4UrH0aNgqk/u4xlhK65OedwEyPCtGBAGsBp+pl517dvmBfuQjcIHwegrknnSQ8kBOKLpm
pKyX6QRrJLgLa5eCJTyER6djZuqwT4mvyhRSc5FrUYptAdQj3nw7pVyEKuGs9+JPDEy37PHGnrwK
hFA3eFQ8XjYfquuzqndhlUYn7WAQFvN8sb9n+W6wDq4ZZGo6zyiqeB0SdKjcTWBBRAweZLkcm25P
KQNlrz8lFr+FL9IgsctEEHT65HO9UkdYh77Ivu0LD8W16KDK6g+fJiayHqZ8qRy/coKGfKsD1Zlb
hmECouogvk5lNB+0zHhguf8SsPtum2GEiDkZQt3/rrmDzChjXECX6RhmZvjCbDD+PNmPKfOdQ2PL
sLZGeR3j4CwUMp7M6bFqbjrmg2bReCdOIf5+cYEtE4QJJX1gOLG8dja943+gT/Cxx/DrGmRJqYKv
EZ/JsGocu/pScb/E94BDywEctzYzjJGU23TH0gTcbJrYgwac7VNKvioxfKfLppS7z/nj23DIOuIQ
GoV2WZ8oYCl5ylkIedF1g6R7RA/snx3u88lA96/7iwsYNWgv9xil1wQBXLLlZPlFdyNBUrPoIInL
xYy3jCntI4MTQyRD/NyNJADI5ctmYnSHUDC8rmzslnvqVJTVeeD6BEfnHMPT/HYAEuQzBPYOjGn5
o7VZAq+cbw9rOj0LWKkoMk2Q4mAGD2svMvqH++HRI+f7UjXaid6ZqfAly6QumhILVR5o2xMuMY2B
JF5eyJ+J2etnn0DWj/WKneFtStA1EjOiDaVX1jqG/zkUtNXfxH0lIGU67qYRGdRTc/pt6Ob5GfE2
7ylWvCPUiJWHcdlVM/0n5GZezO9FXSw83bO6qZN/jbau6Id97Jv25syRrFH2mhngd5EDBOkh7N9q
SYwzG8rTYmgtHwfcjQABlrzRFAeOhz9nKIC50XTvSTYMUObF7aYA831shOs42ovxvXY/F7GkPhjF
9SV07uauvSGT5f54JLm460GVcWhrSDEIO/2osww9J0iJMtMueWzdxyq3L4oJu4sX3S+7bETG8gp/
l3w6d1/AuQYZyuITH70BL78+F1CgP59Taqq6wXwFHPZcrqV13fqMWUrsTXURM0Jm1KSyT6LgNpbG
iis4vjY5V4WKsfwdXdCkcr9/2qMATrP5GH28DcnmocOHYDXL3Fjs8QvmOGkAJjDjKPaLluvLDPFC
818/QUla0NOjDaevJtGws7449R0rzK6TSTm4mJl5jDRDKrMXhvYHVZqU2t/pp7qlrvjo9rvzzKTU
eQn8qIeUk3rVjujDZ4DpGehY8+SRvR9yqYLbkXJVu+uE6adpRdMVMxw0krJyY/RLnQJxtTCLdlig
15U+8zntGl9tjjNAIyjo0TixdWSHxn98tkbqSmxnqUqCgvvCcOuEmHud74uQlQdCeYKSlGJL+Jkg
sfzWu8SdXntYMlPw0kFbCNJ/iBcdi5ot0Bb9oMkFiL0cRRYxcJshonKeqqpsebXM+v+TEW04rSN9
3dkOOpa4NuuouQmT5+PVLPG0ID9z4xkKhjLWSbaVyne0iKrua0MdatZGaCMQHelhrAKKiDMmZ8Ai
aWZTduP+cq7+EpUOoVZfpCjGwetREt0xa3ZNQUZbkwXSwvecZSqNTsLMZ0rD8s6YlQrViZSvWDAu
UpVOMqYUVT7eelcX7OSTgSIeRRabQKBC9OiQTNgVR9k7FGHfnO3dQnMYXLWyY6OctMI6uaWjLQIg
na6rYoY9UhXT1FUo6o9uZUuNsyW0zfL9Vo66cOWkFDNjGBYQKTmlgKVbJcclm3gTCMJKcGIYGW9L
kOTw234NCsFo7MTTwXhn+21aQuxzKAn96FHghmLUgYDvo3pNEHuatymIkGme5Swr81VkQ70piUu8
rKxBOsreorDLuJAT21v8jYNrL5G4HMvH0GpXbm553h8V9YSz5z1k63HdLnml0OaKFZvEKeEAeKX1
mWq7V8Kxp7Z+s8zkJ8LaUtr2+w+d0npn967cGGy//pq5gYfgELo5R2BQbgLNEZg7DlX5D2YQP1iO
ePsCi0AlJUBtYEG2aTeG8wg085LuTodrzutxL1whSTYNyzIQOizIIBC0dr6u6owVafmhrtSUC3xq
JyhVxf6zueZ7tdW+g9h2O4MFjLfFNZRl1fCdXMfoZhSFJkZM/bfrWQyf5E5ao/lMaexR/mI8L3i9
6A20itt2Nbh8NaVsnxZn1A6EFdvpjPU0d163ZbM58Os8EX+UFdw9BwdavXUBLUjfctylnvM4QOgn
0stbm1KoZypYXfEPm3BEZgVR+OrEwuvHThJ7QEtkh0L6Ox2dJJLfwerEDA1DpYPH+k6a7olBoAxB
jcZm0GNuZuNTy6mgirdd141hnkQSaONYxUb5eMn63WT5V/8qsG1GV20U2DY5VYICAtA3eEeCCt5b
Ai2Dy8fiDwzSsJWBRc776F19IDhFf4weUVdpv0UrXtr+wQvqaNJ+mQiGVJ+LMYJ0SlW+Ru1py4qs
dYjwSkOZcArljU3g9axw4inJ4fOlkQuSejYNDePGDqPjGgQBVnETMuaU2xCs30Ul2drU3f3Xbe6K
M4PRAM5mwl4pPEAT9DvSulkAh1Lfppxz1Fh2vuO4EC+HB56tVQQ8EL0sa138RjC+TbVaFmBUBTSe
NqucFxnYFWqQW5uPctXBcpj5+78tziUV+WA36zW3OnWtO0ADBmiuntqGGymLYSzcJvdZ16q5nxqQ
UvfcC3FDPqqOxv0yzjJSMPb791Sw547JvyfwGyK4RjQJfKHk7fkgPlkJKbOKtpnQ8id9XMD5ZGlh
6rLvLV9vzGmHofRQqhCF1YmHepuiYdGp9XGTzw8C/waprixiw9RDe8RadgXhTKADbBWq8KjSVxE3
LhIRoyphTHlX7ud7lU0YJKyDyY/C5zDHb5WTyO4D8j9Ak5m7PTQB9J7geS61tlGBVUuvkAtTXP32
r52Z79/trs1PqDSgmqXwRBPLkJ2DzLqZsaXjS9gWqkndqEUwvow/RcBF7tJtPercT7qwvhPgxbAt
bK/7vPQ1HyDX5eUiCJ+ykDwLPp6Sk/B2iw53IE497rbp0jKlD5F6ILc8VXK6QROEteAguU7DqXB8
JPSKLc7FG3t3qpt+l9ukgPMvNsh6quQFFi6Hk3x5wv8DNiI9mdcvoMfyCzs8OFYIu8oqkz40drNK
BqPXa4CnR7eP5Dih615uCYQDD049j6PTJ1hdGKUYfV7IhVIQJ3kvUScnYMrZItbbCdR8uV4Vpczy
DhEt+V+qVBqYdKo7w3sk8Vl+vAM6E+1tWqi7iEEhr0psHlSAnJ4fBQKOvQQpHtyCxR/J/Tzq6lJk
5rGgu8+YeKU4L5uEdC9/Kw/3P20n2/Zj+QD3WQMQTWVw99hU2iW8HVoqQAlWg6XtjIWS2NNl+shE
2fd7QL9JTmK3tXoCVmGTqq8mZUbxK3t/VlvVtAe1Dd5/d2/+IHDKoncDp9t98cICgp5Y92rbHWG1
Yx4v1q/8wWi5swDq+gZ4DHF4bBCAuKJbLjGH8ig4A0Dnw0AWBgcbeCTqKdHVIBVcd+q4w+gkjwnJ
RtAXRSO8mn0IPTlb+4insE+MuKTzmnqci8n/eZy9+888/i8KlhVtsL069J+D9Da2xZiaLIZCLnru
l3YjBY/wZhr/CEqeqM0Q8uxvBKQ0I3L2rb4FLiMWBcxG+dYybI2wmtphSDjVhgLOHpGcfecslgQr
+gw20Gro5zKw/A+oMvvcZA9hkvwyLx8k4J8c2eXOv3/0pnldkjUSV2ZSwmrWxkzcPT3bRDdx7tSX
PDMhnIkHoVndVGUwoyvb9L21HO/nxBIMDAsFW7I3iXGU411sfnvJnVUi70RMKWdvK4evFP9jLpF9
j74QNPaeIrDkxFiGFTA3ZalJo7vb19t3oRQp/FvNlBZF8pmWsf2OOyeRCN8EW5aXlzY9AC2JDtS6
ZuOAMoASBn8C9Jxpq6ZyrmLCopOuU2jPGON2p1FLdmwobID/qR7kPPtj7iuOqo4TpQ3AKPQr7sSv
wMloPBhy0MJwXD2ld2tKzNY8y8kPKFshhLFnt7FV4hqczcmMB61sM0Nqzet7qdAFfvBsRosKgpwc
5qdfYk5fHtjt51eZCQATRwDLzLizkoAmY+Us1Dv8Cl0WR+m5DcdKoeNjTuDzUxoMABWng9BIkfsO
hrzG63et4EcAyhR0kyJNR3sYW5vhVz2+MJo3scSR+8wlYV7yZdLU6DifJTReoWJIA5IqFZENxbv5
OTMUJze7Bej5hdmwPfbxMKYCGz2/OefVRxPXkOl6u5qC2/2quxVqkMYP//worBDJszcs+tJCmt2X
Ps5B22Md36a0w3WQJy/wTiAXa1YqdkwISyvGSGnOMpvfkAVf+UA41RJDspA0l2fkGyrYbyut72Uu
KNUhVVySahNb+mACsQYp5fGbiYILD2D/dsoC0OnBxw4VMFAVISnc4kYKzI3wTthT8KXJqt+3q+g/
eC02kkzo83QrzjeI9JytlJy9yWzsdA+BvUnL9eAomyZr7qafeKRkXiYeUNEuSucc0Skx8AY/HJxD
SCeqhizXFw8D9008SYkzRVvu4PsKOoNUXqYXkPrKr1IjxIZ79n76rVCuZfeV6uaoE/ZFG8XTTXfE
KdZEZ1B4R1+NsJZsRzCh6qTgHbC7XHUi6QeSs9zG8pDP+imB6l3krlLyVxUpgzPHdQqXKB5+RtDY
sC2uItddpc9Svsik31UPOAUB44NanfOO2eWIFD+xppKF7/35kzEmH9a0IJtJDtGF5GypNg7MYGcK
79qno0ciQWj3qQ8BgdeYUVj2WsprESm9JgfpY5QhBEmHlHnmT4aQKQ5OAWZb4Mtt7wYHWdYhXZU8
V5eOdS63IhwWZxeDhwlRqvITjYqDrxY0GiWVTKWk6/OOSvtQ53hnXNKYhEBeEAIdNqIcVjMBwMmH
sEaN25QFMzPWZkbbVTyYQZkw2ZHIiSclY1CgFGCtafQtpmChpw31ut+vqDEhHeVdWyHRMF/Sa9ib
j5TG0kAks4p4Y6jUm1ZowoQakXc3I211FJZUALIM8CguTmlgDDvfjUZRgfuljIT43JGKAEGpRAOm
qsDOihv9+wgWbZQ9XRo7rzh8lUi9KOh4PPaR5FC3fjg4PK238b+Bk9YK/b8EW+1Q683+wNYb161D
c6MAZJxDH2FusenTQs8wJN7D5YBpP7L8AE7NITv+5Sz4MEx7Wus45u4cPg9xL5dMiK1B6haKa+/d
W3su0oQR5gDd+MCRIxt/PFDnp7hghYCKz2MjT72Lh5lGnSpfa5fOiDR/vTwPGBP043H/QQcCptW5
RN4eVwavqQ6b+C5eeNW4LPLs2UeqlML7cY2aBz7fM2z4NbbvDx8r3Y3UTeG4M/XEJvFJlJVHOGTg
eOW6l8Oj67r/bl3lNkGi1ARiBKv8kEBx4KSVT4gBWfGrb6kllWYVZTEERyApcqD25VV8hpBKeP1W
jC49FwUs3Ymu8Qr7wjVcxc7JkiFLBnNbvKtxgNsNNip/ewWJe9gzWEjSrAgiT7iTSsEf+8ewJB7m
yWUaCw4IBoq6yOZK/G51cCYfiuPk2UPJbyfxIqqFJrqYoGIPKk2hOFOHHgmpz68rniEygKxZOj4O
uSh3jWgpXfp9VZIploJ91h+eFz/YUnk2S6pn4MwkXTETuqAqzuZq2KL3Y79vaHQ/vGjmd3yryxz9
3DdCQTJKW0ob9PGhynzegJNEwGwU+2fnLF0xfiCIeJKQH0S/phFzJVnRLfPWkczA3eFhzWJ0kcBA
JDb1rvFSxDBbVvNxOAXObBZFTiogs9V4ME3a6ioZIxs6+GzdtoD7X59Z6b0PWykJpe1w+ypJGH14
qoBDiFCzQfqKCMpz2gvh3t3zZVaxSmqNdFoFDD6tQQFRdppGLs/BQ+eFB5+DBAA3z3j3+K2YPCNj
ohGLlYd+VfW8nn/5pGFFCnIupf7QlcvQnRnSY5Pa4K9/+o1oc8b3Rm3sZabFFjJVqGjG1Mx7BE2/
A9nnkdVLTHQTXZb0s16LRxzdgLRKI8kerOh4DO6F+3v7jHbNtcLjVigLCzOv1Q/9gd7o1bKMdRno
9X2F08rbxs7PtC2ffI2VEhHqpQWvlZ+MRT9XGhyQgu5cHWj8O7rxCmWMoPL3RbBQGuy5oxq88vXd
KJ7EHj2BySPxt4tAbOXmrUoKfbdwfgJGp5yoDUAT1WkhTH4cRM3Zi7va2dsRldiPrGJUJqY8QCHe
sSgJDfKqQaJ6/5f9qfxUyyKuhLvDLRe4yVVGwwtxuNe+3xdISNiBa2UGAxMDo6/gNh5P60DHoYls
CxkPuqpIM9JkLbkRExRXXQzYoM3sHL8qSYYBqfuSVzLBMNe6Vk0UlJOMcgCp3OeILZwdlA1bBiGJ
yGRvzdIyaqoiDU4WRri/yqMESvZKNl8F3FllkPaGBi3gyKpnOPqNUd1CWtXEtIHl54OOkEQ0wGtl
rt3sP4sdFm4SjVOAFtkMc1F1LYxP5w8K+Nwmlsn2tnwxd/LjFjv7jvx2tO/7bRs3zps4uGgENGyC
p+puUC1RzlKk2xcQYvLYDziUT/5DYEeInVzK/6ayKZVI2F6rMsPsRnHGR5vC8So1ypViRJgmX4Ab
2QVZ1YJ3ieASwV017/fjP6fyvlcEG+nTPJvNBE9c262WrjkNuQM/JwsQjuU6zA+BN4KHsR7XBN7u
yjYugzLvMGgsSvlPFFoEHO5dN2RjZuTOHPEvvIaBoKg+numYhQ4PJL1Iyde/e8UivuId87ggvD3L
4NTwGfwVS2/huQz1n9OVPUKNCIj/CObxPrTcrlyTGq3u2aYE5F8/TtvghGPKgdLyniLsMrXrJdV+
IhtD776IcgmuDhm2EloxLnGVJXKIDvYtswjexAe7CNkrz7jNcDamE/gg83l5rdoefNWD0N3JlNYR
2XHJtl/SP6OuPOczvBRQZJbI41SjZB1MzttlKXS4lJxgXlMVPwlbgymZgGhhS0n9qbr65kzrGF9i
KOJfHnh4WhMrmQd2zL77IR8aYRpT8VUOBwyOMX5EGGvVb4IZzcM90Z6mXJWkdwuEg6XpCAkGA7Ck
etY/JCjC0/novlVCk7TXwoY5DmBCUu7KZl5LaQCsTStiqKwsP7t/bNvAePQdibF7oB/BOXlOebnC
KT6moQTvlx3vMu/IcsYow1uKiq6FW4Bkc8WaGNRYE8qZYYZ0RoGtRSGsROFmN438Dcl6ADqabNYl
ox+ADdxTqyj9ZgjvEU49yzqSt/lweekg0J1IrgmtLWNW4WVNFK+q737pWyWGEHyoPKPIoaoQ/lq9
qc/XSQtGOwWUJeWa1d+D7Mk8FaNnMXJryFMeYM+dWdgIecKY+u8/38HyA70tgXoR/ToMTDI//bmW
RIlE/+P8TW3C5ER8PkKTu5BYfsWrqNQg+DwkzBltJ72Ln4+hQmNaTyg2AUj8vDydgWnWa7kPhZQO
giYCLTwyBczqn5uT/XLdSAN84i8duqEMzqmN1VQA1+ZXc2UbEekZUOD7LQZPeVNxSxP6AenrfnWD
qXA0nb7i/ggzkuEgNOOeXrHSlMOHdRRZRpu5lPf4vR6I93aMdVW87kGJKIITYUH5LQSF49e50eIS
q1e+j7QkU7d9/JZ9qYCIXprODvQFUDUuBFn9vbpqgINKrSquTr63lfO91UZXh02WN9WWecB/8ixp
IRSgj6jxbRFee6SuQFUq1gif9im2kEucxsQupumooO2ZDrANcl7/pFDW2hXYd6CRFM7OLnp3TZA/
6UlruNjxEw2ykbXCE8mXoo/R1BzX0MX0WoHbgXCgEwtOgTHR0J7CEV5BP/ipJcU637ah0luUAjbM
e6casWy60fW7yG235A7tGX+8EsPvDLl+2rhoFklKPM00udZijkrpE82X9kP/+pEi4vE8w4yDNUhY
EdjD7O8ZoI9Ktx4R9UYze9Rc3vFe7+S7dKmdpuu4wCZf5yQCIWKzecKvktObKRJiCvGRpUWO0ouP
ScJX2ct6qrA+sGmg399sOknHQDFOeVKv6m4E7GY8JHI2SINDOGMRRAvkLi3G/JhntxSLdk9D4gOw
0bMHYkAlRMbACOle2ynl8pmcViBWpS6P1ijzQATvySb2UoHyTefs11NkGa+D46eijpg4I7jNtXEZ
+5cPyaXv5dd/RhoHT2Z4ryUyQkpHMV0p1/wI6g8Fae53z3LtI3UzxmC9DeGfSidNRdlVdh+dHxtq
TtP9tcMXzVnG9U2KBWh4b5JqA92khNwAUkWy32T7yk8pR05HPqBwB8h4rcq1lFCpxfkJCz0wdlVh
Y6BUOPDH4qjLAi7YbJJ0qa6QLyTa6S9/NWtHioDYBC47e4uqxGyzY+nngticQEDBMmnISv3xZEo/
5+uY2QQ0cJvOzDksJXX8IYLBSxicrMlU1yA/IAqvZVPJ9qNY664u5a2c9A4zW1GOiKT8ja5kgfTt
EpXvxUzAqB0ZjNZ3/a58LKPfmow2ODpXQ/NhhW5oo7bfKGBuMKOQf9p/VKVt/OJ72cWCdHHASSvA
pyGyeow4xJkeiCGXtpIRwnv3exi/SOxB3hDiAzpju8LaPaMfthbrbMwr8/qITMI23P4aeCUtk+BN
mZ88DXOn8zgOpGaubPxdnET+sHSNYINAwKll841T7jdODw7YUNajlJGb0d1AW6CumF/DyndsGcat
BkOi4rH6VcVQZcY5NNpNc9+JbHV1n0oK9pz/Dlo2qLwijLy4UbmMG279nPGMgbHiack8GWHhH+H/
I7Sh2yr0jB38m2UZtJNYiuFnWHOjc2ruoZ2E5Tq+1Y9V2hgIPTZzxEk+mCGgSnVHHOQkv9Zug/5g
WTqQp5i+/cnCZc61x9IGmSEwUjwizW91d+1sG582LeU2Xm3E1LIQwSw9Ui5n9Q/19yZuwMkxMpHi
TVo7GC/TpE1SNkeLtZLWyckz6i8z2mtXEuT7SWfkgc7s/wJMFlRyUx+9V8SncUfeZ60+nJzUZ6X8
ZY68B5gmRfHKTxpCussq85NvVHAGoswI9Gq7Dp88pZbbqkUXH2mYGVh+a3tLgqCd9HipBJYBdtbl
RWZRNq95TW8D/KVbMSjyQhoGskElrFYXpBWcz964LrX527Aqj5rK6cX4xnz0s9d0uI+rHzAhDnHx
V9xAuvV+6IAJ7z/e9g6V755PbOc5yzTThRhjLS6f8h/5Wndsjv8I+4+nroqMhjz/wObXGdpgKtou
PNl0m+vsoE/axTuRMKxlqt4JRseq9CjUt6r2wrvWgcoJO7Rp+cMhgMRT6qDkR/Ed1mHy8I/y+7MJ
IXbFGo4CdCcMF9kJkplRjaDznd3XnTgTd7f9HySmKR4BF7fOWb7GL7B6kjoXyFEBMiaiR6tCq7Ht
WAtpEsTkGB6tUmZc/FsFMPr6Tj/+4pgUmygE38gTVLlicodbjohRjKE5aqq3uPcoziTREqmkOD9W
RMRvEVnQqwzRenxMyZ+4ddAr6CjBqYdJUbo2gQ/xOBUXprr1PbYmtkrg3T85M3TAIHAdjwxWr7UO
Jn+J/0wOwabDVYYZDERStE1bOJbCNk7ZZLhKkZHgqh3TYgbym6vF4UCKD6L3MJIqICQDbEK5uw7r
7UxpjGDFybFWw9jTP8qhC72QlxSZI3CB+PjYA4JJn0a2I+TM62NkR8ntZ8pNb2QOR2WM2dwsQNCC
rKmRIj0K47g+jZ6AKDy1Z/IwD51PrC2Az0tdNeO+UCUFQfmXVLyfPXyowRHW7srRESfVJ2x0ezpP
Tr/28qKTwjCjLfN5YXGfzXLCvSdluSLsYhzWvYP3pe5D3vveoKM49QnlqIh9WbvZ/pP3N9L1Hulm
FOTImvAmXnpzSZ9ztnKW49xkXUjWMIrD1fDhtQITcGxZyJr1eS2zvj3AGDMPzx+hRl//U0QOoUDf
ZDEK4cltc3YzNLvvULkMaysZFrWctuecmiifTkXW4k5oQ2PNlETztlj+w6D/+sfEKwFlyk34b8Km
oZvlNn+li8eIL+va4vzQV/QKymKCGjxsgkGChoAJuDLHZ2+lrLTBe55nMNqU88oMRMQLdWs8Oi4J
OeXBnJvw0bkz/87TsCYjRvubSmzXmAoJrZo10LirUDPlk0gQ7dQXFnbxvoW4mWDTXik+cl6fmUjF
5PUM0hXWzOC+cBmx1QEiyZfr9Vy818Kc9KulBq381b/xD9iikqnLfL3rBdTfzzzUhaOS32Rwx5rV
Jw7E0OEQtWJwvRehsaCyGQ/ik6yDqHf0/cVzCLkKClmz4PUd3rPeFdDkTI0pUcKdmkYpA09ktkXX
TF9eSSHweRWZdO7vOhME8eF24jO54lL15vI+hFvs9er9VtXAzPW/NO+qFhxtt5Kgq/HS8VSOeH1h
U3A+OfUG4Rgof9fF6KfvVzhdRtHZfoP+xGwYp7xShWXTGU3Jt+kIgKKANw/FvJHNLUFQcrJOUQrE
H1GkvZGexTGbSYjqdv0P5r21F5GFf78nv9QMSPJG6mvRU3Ro2E1JDkBizGSvwlbDWqULDY72A0fZ
RJq6SzBACRuFYBw7Kfu25q+BHlWzINBZF524+9QflTU4Gd1xbjadYk9R8VQgoCmkQXhE1d2n9vBw
fxolVCwCtZPqG2/GPPN3Dp2Gdz2RYLTTub1kxevNYQ/+OfzrnYeswvQ6IVEgPTzQgvz7f0efFSTw
eEDcMhUZ5rPzgRufA26kA7dB53+k0lkLvlcVm5Ib+HDVfy0pEG7Izc0JYk3WkAvyEic4hUJzWoZJ
BaMUOEmskq9IxMeVE83MN7mxNt8VtlKe3J8b1yoII0wa+Bno3UTD2GrTNJhG1clqD40UfAOZrSaV
rKeDPByQ89n32Th8xB58xROD2Se7vzs5TmGdU813dm8SclJjWg2DpPRfN86JISX1wOc5A8TRug44
Reo6ag7WBOxT39BjjjrRF5jRG4zafKs2qzxczad27S6dDwxtTWQR8R4X3adWIGn0+O6BV3/bR6BL
0R9P6oFhSB+7yTXewM6izqUdzDht5PZdRpLYlUJM1tbPnKMUYGsPoapesQgkP7u3blHGCTXV9fCa
4X3Y7PlVpLDVLEk4WtVpVszZU9c/xDDmEqvvoOrImo4XB/g/V35gxSsOYJEp6t+NCVn8c1qAPEtS
u/d5T2vuyzWoTt2uI9rGdj9QS5ojLEWmaRYaqPloAwxP1gH82ob4IrTaEhOi5QUl/dXDWtSgMSF+
IQtd6O8TO9X2Phmj9scbX/CuK949vXbC2ekNtA+CpcFbcQWyXjhXVCLtsszRVIgkEhs3zMsTAWHc
KeebWTgpCiiQR2vZSIIsQhwib+mRT3C2UOF/JdT/3GggYOzEH91CwCPCJP7q4Z56gyLBfOwT2l9f
ZzGuWqN1K4jldjGfR+l/vPhW/xH0YvPrKlDjiZNjsh2UulkHPwS51OLFeBV81VE55/SOX+CTwYf3
uICvq9iQ02tntZXVPBrSMCRtZAeh5SnlZav3GvXtwbtfSkjYFL8cbmjanvh8wYNTDXX3pYBtGPel
A8sYvwcV4y2Etuf8VBaq66STo0KfjirmGu73ZxR4cKF6u4WaUm8aYxMPGzDSe+QcfClQRJ0t/IYz
sA/2iSi79i5xQNThXQFU3pJP8Y62qsiw21nw+h9fI+X55m2j/7fHVYs99WO4Qmfa8RiV3WEtDNI0
qnIs0bk4ot4tQpo6aeLtcB960ZAgYyErDnu+5K0ObfjezvSvgiOXvfv6f1oOgNFrh9SfIn/O4hgH
ww6hEs8RxkuwQ1oxZy9xAogukkUsQPfwB9UARc1aEXgdty0yiwqm9QYy3anWt9ZraDbCofNZ2BWB
Z88dGH7iTGhUP6ZeHW1DtAq5DSmg2h4r3g/ai//5s45t1CRBDgCbA7NPJm7EZkGRi6oMzcdl6HWW
HDW3BQNAdKLNEA9sO8VEddqG0Q4z7hgJzE3KsOI7epW11Lu/6h5UjDSgodxpCEh6kqH9MZALzqin
0FWsO+q7wfqjq84ZskYzRcjnwlWqJbx38qszwM+HSqYg+S1alFNvN7B1qET0c5tBMVKAGZIKnXOw
tV6ziCw1WQPW+/llp2KWYZQXBkma/J4MQY4XxfVH3kFlQt6ES2RV/bUrNRqVXDZSgvutulbOb5zS
w0rldgpZlu343ibosReajFvJn7dmXouf711OlEXMbQ48BjXBAOtkzuOpKr0wSlwZMEazsrUtSa8K
4rIP8jL9dyqCHq65hVaMtp+7BTS0ilw5uql1D4gzhBxd1uV/kEffGh/FQFnkC5uuuykDiKf4wTp6
y7F0gLHXGebVUFuKji692M0jJ2uWKVds0F+P2naBkJnOj8Sgwso+sO249WHIBZooZyhbaxb70ieF
JkBxTQUWTpoD5e0bCapc1uRPdWbz0X9D++PwL7YbiekXfWq55EkvmP3gVvokGuFoNH8Cdbp35DiK
AW8PiS/LAlXKqHNyrvyJcRGnvR0JJ2LDPC+8WoTniikDUO827Tg0UgCLMnGxzg8Y04ffv7F6KX0A
ch3lJSpMFyrNx6O5Z8UAEsEe9OyjRFLMb23FzaCSKdcqr+yIcLuezntrXfKX1fmmPewL9J6DMPOk
OEUrracVlfmkYU2aM/vraU5Y6/6dk9fdyigxn8utefDDOMMGJHsXKlhderBfhMN6ryna8xcMmChs
8DXF9wQiA57aQTRE3JYp/q5eIPtyqnbc08AEmMq3wuIktacICl26eU4s2uiZHnqHuB0lPe3F14Ey
RB7oopQTGQ9WnUeBxytmFOvtaQUOnbIuA+ti4o9YUi2OQxi9/VSqMSIM5oMf0PEYH5vCWxvUtE/o
zkALzhoYPxJ1Fkv0Bq6rYl1pfjk2+R3BXTmSAP1A4QvKK2J3C8Owc7x/ZxY3mtLUkJGu9NiqSJoz
YgaAczVHQ6LHaqbpaUHdq3iBF045l2rVdpp14qEeIAGxEkehRqmIAwsm9taKEOfgqBQ9wfyg83Pd
s0GVdQlRcJJGQW9ETXfpSYlTX2ENqMRChRa0EoRqPOJlmMw9PC3QP5Ac60TSXxutafSCr65nY5C9
3S/cQtPYycHrt5vyzAk9gh4DXolhRcawZRBLraInro13bXW+pjfVp4peC3oQIXGegpY8agN6yEay
NQr0L/F4+LCqNMAZ7/FpDcOFZ5EprlcXpXe7h9lfpmmmfzXb9sD/yxDfpnq95VXlBC83x0PBZ7nk
zeQ+5JOfKHUbCOeL3/GXdTuI4tuMfstlJgSGEkoXidEYMCtchONJdKhsHOC4PEXNbCqp/Nx12wJH
5HCSQxhtKudNfoQ8uge4Yt7qBxDC4zEvZGN0z5wZmj2PEKWfsswmZBbS/BlAEfyJHVt64BJzfCrB
N7BFMa+zstugf7Gl8HmYugJL3+eQaKLxTeGFDzMC7cflPh8wsfumy/oAuLqiZP07k/2bN9UApljG
+h/f9KiSiAvK9OxPmgK41ezFFEHwgBXxuXVSxZUZsbECXdgFClqaVqWBxE7jmSjtncGCiuqwCpgZ
fSbbWum+oipLbhqLWtOTd3RLmgbAPLAIklnFCs5KkReDuxTilfRskca8T983GGyA8ZJRllbNDAJU
jSRdtEtk8dw1TLiLDhOvvOeb6xo95vlbbKN+bB78RdlC3TOKuFlGQSHEa56g/3KpCrJZMrq8HE+y
eHzqfbnZLdHa7CnoowztguIfTuWL8d8jhmL5XviUDiF/rKcMiYjxrJOJ4LPzI+vCNea1FzRvjFGf
sn4rQLPGcrzloBgwaYt8q2qNbZjFH6XCIhdKQbOgS57EOYeU11L3/oCVNCcszieoSOXFLCukCiA0
XqYbMksD1neHhdj0OO9p+BXsjJJgaK1gMZUKI7+zNpCigr77FNjbBox6wD3TbgZXnX6IkXY3M15x
3c7x7jo1jG81EVsou/rf0eDz/9a9PzWepZ1Usl5A1aubxUU2Dps8JH5zf34TycJGjVu2Qp6Myh33
tV+i6lzyrUUubmG28UvH1ihLv2Bz9dobAwp7QOsZQFYCezbzVSYOGsiJAjI7z9zWTRMp+EOntu5e
gZOO+GUwQjbLZiFNuWkIyo/GEizZLOeTBqDZVW6IRYJT1NzQouRi0K6O9pu0N8WM/kzzQRClkJc1
Tx+0Om9uQuvHpGI0r3TpetvHT+VzL10dRf0iDe1NQbzSu1krykFriramenQwGN+u43J7Xq7O6FES
kwKej40xxpvdAdMW+Lc/HvgFfDC+LIEthH0f8cdCXrYdWwz8u8BWBTFKrCBi3I9hnt4PSWMcoTDl
C69isQqiaAIDowv7MFT29vSsOnsXDEwOzqKje8B+pLDOsEEodYK89J0uy+y70K3kJ34RDKyO+mRd
LWVA6tWd89X/GioMoZreYBUoOzByVEjLxxK2UXbgajTQG1X8HDZ5uON0uKXN9EJuvnIko7o7nNGo
RyF8ux3i+3/PmJI46V2rhQhQhnNxWI5PyHXR9tqtrp2Qduv7Tkx6YBPqId2ef3rkpBD0PFG7DX0Z
bwyE3utSRtHpe9y+FeKuae+hZeTBOWMzKw7GPJqDHmcfkPvFFc3RRu+o66E5cxiP2zk/g0xKFHES
YiDPZaK0YKHeQc+7eZkF8KD2NPhAYx4kQLq3Ga2SAvdqHNiAqrzsuwuLLw3iJ+yn8jkTSZeYscyj
P9EL0c8+WQuCU3hho3+6XyM2WjIYfFjSQ9jKJDrbVra4NWJD7gsOQxUN7DUIxdYznQhNlmqzoXjF
mKjXtPiC968Cdze3v+6En8Tvf47yLG14OYgGsA82/oEUuq9bh9IH2M4cvHzqq49y5LLF0VpfZmmy
SI529xu3OmlJxrsHvjaq4LNi1al5n/TaA5Ti/1l3SEf3ffYSlDdoOmr4Gq8pS+wVZSrpxVXE/H2x
0bjRDa6bxxBZQj48KLgNwpvxd3SMXzbxfXSQqdJdAEjJG05F/N3K+rF5LItON2cw6gtGYdRw2VoW
wA9plf2QVjTC6/QWlhfPREcsAU2TP0IhebRpgbktR5xr5nzY6TxzywbJRSGzMUfHJrxWdQZYNmyg
/ty0oAJ4gKgeuVDlwZDxEapDREQbOLaNA6O1sRZyj0r+kQFbantmg7Qx97mQAJnAOt78yc22a3+2
t9lV9bZEd4TgVNWYPttK+EloPJkMZvpGiDM4LPlYMn2+pnxrE3s6M/vnf9qcb91SDSKvb96zLxpk
688+GXW5yHWBWF6H27AaLoUC09wMUDj1ZjOufVUsk7dfx0onr4jQ3dmLYSSkWxZaHlz1tdNF1pk/
w2GchHvY1aOHv91vc+uD34yg7PKJq4j4exaiK6YvFMV6fy1PU7G6TFBS+VSwWmdTf519bNBS4E7o
bDTHFI6Hbb3MyDGxoDKkqcamDWgACs3tq/2CTH+sqp5jHeEi/7Ro7WiatKhq97IyEJ6RRgto0y9+
S0sUpjt4NmjrexJHpPDK1F058rxyvLOG80D4gJdepTGi1LmDA9I3ltxchjXdwMk2isTqKlgIuN0c
0Bkiofs0C5iyDtmyL9zIsApSx3l5wqAcfgW61PjkFWQkZaJctJWRUAohIXkJ0yqGJMY1HhGxA0TT
pHBeJ0A495kMV1/VYH4N/qEI2YdPDFPHtysaUh+k+03Tuc4pgq28NB2WnUa2RrP7ilOgJ110qCaF
h/aj9Ibwbq1buQIB1eJpYDGysa9eqBEQ7JhYfqBezaFwC8hpD0kDpNgP0mpve3PVc5yeqj6X8hTn
Hz5OF0QnofNKYDffbgrVRyfJQG9iXe4YcW5FDImsM+mzIZhwREt/HGKd/JOo06kTafoJTcGebl3C
Bzd+sALOdfMwtAkfLSVEvpG5ACN8y5uyFOrtYr618Pcxig0fqwZe0rbSRipMqy583/yMp+yNEvGc
xRuuiQBfp4SsSlMWqGL+PSWj9qeydBnnUejuUdi3CQ95R7fy4JIXOxW0S2OEyP7XfMoJZ17m1OuH
UND9HaoVAuZuSZVvn+MhcD1ZM6BbwUxCpjd2E081VAR0BnKamKKmABhcdtusiZ+3VfzkPRpUunko
Xtxf9712LDlFWVicxd8FNpsraJ3JF7yx2GuwQyITj10uAmZ3IIeo5iQnJyvK/4dHuX9wkye3ko9s
7W5tFsU3f+Y97BCFfVVT7LpXxexf/qI+X65F0gNeKyqSy9+VCYz+4C2f0otJ1QpUYYKCkf2MBorb
NyfzqMY6aG9rNahHN8iC8Ki3lMb1evvYyPucnL/4oFRi2TJztuxXf2+XYYEIRzVtFMXcVwLKpo80
7/WsyWXB6BEYMrXJhI5kwTlVhV2LMKbuH3lpCtGgnj5uVANIkKgBm6+VpbKVTYzUqz/F/FNRCN77
U3woAB+ieDdmosOYwYkzfjxrU1+781IOQwS0PoxRKxcLjrIgJNvWfhQj1Kzc2VzEMkPJEbXGsCRV
40TOakgBa9fCMVa0iEeMI1aYNmgNYZSfs/KVR6NRIIyEDmE17RqJeQsbjUjr0JFX4SfrAruJx1iO
5uGTBfi5INdL44MOV9gVwGrpUxW1ti1Hv3lhnEzSOJYAL/dXGJNF7e0tTb4zIHt2I8Luo6ooUmFA
wXFNbrUxd6sq3ZFiecVgW2hSi4pwFf5Nm6Ce+8SgEiOgpQOCUkins13OXizaWGbZNeqUnVSSkKAZ
AkaQaRzFv4+z604NfCw3Yq2rbNi7cNkRa1VSCrqH9MzcVglir6Chzi9HCYN+dmYqwJnTzsDNTmDd
cN0WysF/XCcsUVZ0SVxEtlTd7JctSdVRvH6aiQzYKksU4EyjlsqjMRDYBzZWOp/qkMTOoTugd3rX
TKA3Zw+1lgsrpHJZTSza+ftpj0DuhCWFKJ4+2n3CApO5XyE7oQIP5kKYsRrXXxg3rwLIutN+wbA8
I1tnlyDtE0AX4HATPXqydjsyIs3EycJQ0yrett/+++zjRjRoMm2xnVtH2M5pNDiM2S8rj7PVFqpJ
ztxOaRWGee2IvqiW0mwXoXoqa44jZyKldvqpXZjg6QqXUOmmrAK0HVUyQlE7kYAA/LUiP2NqKsp/
KM0WXMblsulVclDpIKaxuIHlAEjNJaEqPyFNsfH07+pQZ3RmAcNXbJ3UPbpwAhHlHC2qL3/ktCH8
PdAZEtoZb9t3uHmHt/cbsxwH7r9DXq/Xy/ahaf1syMP8CFGgtiAbqR95hW2L3AMKxgckk+NAVgnZ
HTMZYl36kHRarnZFeixFfTrx0SX/vqgD1HR7VNuXedeUXM8H+udJfGiAaXvOFIM4HGXJK4kMwnJM
o67chavyb9mUlV5kopmr2dSkjOwq7b3lYjscVkakT2WXUTiPzby54Nal7P4bDrebJjwRUX/GnURq
Zjc/vGAnVnZ6uZMFKoi/ivyPoN9OXX2zlDXHb+IwX0M8aIh4IbX6D/KWdGQZnnMIubQj3DhW7COk
xEqnYwW3r2Rx3q+2PC3OS/VfLzOlx1YxG6ipBcqF8eH6aouIIa5iONt3PwgY16ZjLVzjzcKB1pJI
Sc1cvXYq907VckJyh/v84yAtzzuB0fKKDVT3wBhb++WD/KEDgqljfgNjiGCkL03pEyYqjSspD3Wg
/vbbBSBJnBV6fBlGlZYGKtRzAIsSh/F2FCSZQORPyALVebOKxrOtnCtK299WCJvHcT5XFuhmjsBA
bQAT5qqxDVR7XlN2cc9ILwuq/m7vm2LvrWQ4WPyq74RHgK37OtwmwHPs9TT6cI5gP68iBCPR1HAo
Wr15iIA1zd/TH/pKLEN6Bg5gqDaFnqehL+1Ed8c5BFImZVi0AHcosjiwpN1T+UO7JUtpt/kYd9wZ
X3WDPJo4ufiKIBzXMlhW0fOsw4Uib3djbJOQ0tiYBYzJaT4X7ZEqLSdNqKdu2RdAzEKnrBNIzcD7
kJlfW+YkQoJ0Eeispl1zBqm/pRcTGj9CbRh0nRGVFFrS0tylqejkuPJRUGPesLDCwzO8h0iyup8N
4ji+egsAPd5ppTc54RCLE4GyKwUAFLIdTqJu3dxkACJLicGCCyaZfaZTUmNBtitpQIruwYNL96vx
QwtUZ38mehS6eLwSq3N8/lKIvxkY4Y2fLQMICn9JHYmnCapCN0izeFjuFKVRy3PJznTnLCBGToHS
0KfQVygvyOo75LCGHwlpHTm5RovMWbkypNdYPmxR6D9ZpVfuua+EjiWwPbtk+WJBjKn+mN6LuHFU
5g2SjgFvKLz3MMe0nn3wK9N9AUvIzppAGrUCqKpVtG/gk0eE+Zl5w4sqcFCl9uQE6A/wHc+7l/h9
b7fStRQM3P/8ICC1M9umzf3Equf+O9DDv3q9UvMvvdN8vqA+6HTd1/uZZWE9BboF7V3slUNb0oTt
Pwqu1bInpA63YUue0hGJ5IBihFOHoSvrwYOIkRiZTn0WUEz7YpWJLj/sHFuMXmD5/8omIbn4Cn3o
TI1IpNviuqvAiiDunEpGZP+matM5NlOSuQVzLYYgAT6zOKGOi2JAzKKFLGc0rzlKtkjFID6+0quH
F0+vajFbvwlpsU2SxbEooCmR2bEUyoNX8NSP9gpYxeBnkxVqMr+6ANS4DzUQNOaT/Nv2313juPBc
ySrjGqMClQxgQS2YsS0cQGwFbYZFh0sARwZo6v8g54NP7ssc1YoZaN/gdCgSIj9357jTg7aCUMdb
TEQkl7UFj4QKmHF1Ae4Qzs2wej2WHj7vvF422gOFKRMFrY+EO1hSqXMGAnf1/0SxSGOP+jYrCYcy
36Oq1xgXLjOk4nSQQiGfftzGLdrbQWFIx4DDaUiGw5lqKTw/6mXkFdGbWnrlYxnjA62QtJQkiblJ
T0FBMWQlMnGGa3tJU/FnNPWbKxpXryzdRIrWlPaD6CGvxO66DZe26rj3hJjpi735EKn7D+6TCa4A
drZpngL8FwgRjLdUfxoN6D7FSLBn2+DVPhskMxtijINyhhZEFySlbnuyQlFPesOljqKBP4DOKRTO
KNi99OMkq/FCIOpoycZ96DgKKZKiFIHYJj5r+jok8iG/CLYqsR6jhizH1yykcIwGLLWy02JGqE6x
m5/5DNQMvYY98NHlVdQdorUUrAMzEe+vyD0RW3PnHrJdcD3o9GjXwCJxFCccTgMBpz+nOBerbQGB
i6CZn7dtybEwDt6y5mObbOO8STG5MeBxmY/JDSad9RgpYjvzVWBCH2WyxVzRZmo9fG6SMnMUvcm7
ijLaKvzeGm1J3T8meGU8GFBDC1HPhfXEmnzYnt8vfYnnp4J2Rm2iFqHgOxNsnDOiBqOUIJpWyX3B
K+xBDto9CVi034gh2c6x+tHv73+a02ggOJaJFhXQEzYDIJ350DFUmXkknDBYeKyqTgq0oLeNw7hW
61NdPtG5Acvcf6NDw+mBMZJ6CAZZ2kdKkanS3LP4qU4OlPnxinPuCBoItN4pOVha15TCd5J0y/5t
1FNqBsd1ksWCt9PBbq4iS0pmBCtXo8w/KBp9UFFV+t1WaqGxvgXLxlxbNu6Dgv0J072TNhAH2Mao
g2vK7xnNqQzxHEKS2Bmui1gQSVBdtPcQqL/vA/qaA73aj0j67JJlIpfU4i5A41s9LBW6fLG7/Qtq
Zj0RnWVAVWC9F7Rd8jcYOnCntba9TebeUAj2DS+OA8BhMKgFTHwKYPRZK6VwRCASiMuWKR+5bsAV
x3Mv1OsLy0UuYyxYy+/JNVb3z2c5QTuYj9heeIkyqAwL7N4J0DWKz2lhbTE45KdRTWv8tgAutGsF
CQbbVCGpVTPIIydsB/Kam/uQZ/UN3jUPaSP0kM+8TBqFfWk9hn++66qYkK7zDVSn1WUjtNmttyYp
SLhKPaMZkT2pjmLB/AfBwt+42xbUEgIPds3PFYGEsXxssXIKoWasdKT4J32AauoVxicMtqIMCFxl
gU0l0ZnzYVf2tORRhsqOz5ckf6DwHKpEzuz0EKZTrZPBw9D3YCDGgFEO+8rEau/Uwdlkqmhg/W5O
DqZVHeRxLFnR++5G1hLM/dyc6pMzOZpH/FgbgCtmG/kWKepRXpglglLalvjaRdTCh6wRMEIrGLcw
Uw4GVonP26NQc9K3zaTkqaw23fDXMjSnpRIGSufzmoKwpzzueG8AwXlk3pAr6yoKcAA+nHJ/i1JJ
dIitn31hSeHdGAJQsiTFftAFkKv9FypPzVUsAAWe6BFHdyMGmusO1D8lkLUhRh0rk/DuehFU1Hp5
gl/uYlt9dkoZ3mmM7DQPzll6UmYCVhXRHSps8u75a8AgrD1gw5BAkKlMUZRgChcMy5G4J3TRRvK/
+gJPYT0P+1iWNRIDi1/X2CdsJo7UkBezUwooD0wyv/EKU5JKDjUf9hYK2DbelD+mvZ1k0vCeur+z
bQh+/uJq96baqXS2e1LCgKUDzZdzdXgn7DcCcgQBc8byEdHb+n3syRIl4YeuHWk804xuDvf2uyE+
oMIzNDdAb+iQuMHPGhF9QeXVInkLhGwhD/Qi9WvcmdmtyG+fJenfiKpQ+eKqumuJ53W8f4BnVffQ
4OSbmiqauzqhu1rZM2N/i3n7ORFFUe6mWvTFqEj+agHIQ2Srm62mYDumuEK7lvbTLKqsLdCMbOrK
K3pKMxsPCH2OvXDzPzdVV4mkyWxmyKkF0KBD1Z2YLNXBvARXFP4klMXwPbKcAGjeUnSuK/E3Yhf0
gWe/exOIn/lOyjJ6uh6odv7eBtf7sWGbf2ZloenNNfVlYcFtDjIeGiJCKxh8hW7GuTZwmmHRE1Rj
7EXz/eKMGcww9iWxQ3BazGZw0vnN4F3wmCDwZ/Bs1N5g2kCOGD4Z+qyzcHH82Q05ry25YRYRHNFj
y5R3yhSApJ3Jl+iILFHGIa02AVGDJ7uRXgJtXPX9uP8ViyRPuMDB6RYwS2aB5aK21EPnQb5w0ZwS
QoZAiFOsi03aPXoopXn9AhmkwOoWMaSyR47fSAHyJCdU6PhX46K+LT/OiqCySx+Hm46L/JvLrCHK
wJVfwKJAL+vBxeIT7K45DPcEs0Zo5txnATJLhadVItK8e3zUnRpRHOUUy7UsGr5J+k8EtqM73HHH
z8bxNa8AxB9al0dt59VxPnp1vy/7nIyDj1uku4EvJ12V1G/uZGhCfbie5MoQUjG5V3abfEHZFzkj
hgKAkxmGwi79a5Pca7QB9/0B7ZkxByrCmLhJpcfzoi03bn4rrNW87wjNniCRyfk32IGboJ/2IkiH
G5ztp6XFfPCJs4xr2H26GI5c4RH5XGXcz7itEK3CP6wgO29ERZBu3apvfEti4D1Go1xZ1KM929Qj
rTpYyr1vOa2fBL88vp7Sw73BSYo3dMQafQKc4CCZmxABSrwcKNZ743mnqDcYujjxeU7FHiaSwq2z
OpcI0vWq49yt5ZtPrBaz8aGlmdVuooUmmpp4cLmko/UgLbgcUcnqqNwRs2RAy5zg9IqC+a5C5Vzs
g+UNhIRdZ5EzlBdodoywUio3HePfQFZ4DEzfo31iwswt1iwT0JXwXUJ87RgA/tFEk9/nOONsQbpf
lTfCw+nzwRb2fUxzCuGc7SFMPgaS65CiViuA5DCdDwP4QUs/yqsg2CYwbq+mG5pNT10M0+hEyq76
tMvWmTBKFqiqZZ1Xp3Q1Un9blcOeV+Tfl4QBGS+IZ56fkcWIiV6FOdBIDtgfZ4fH2qe9BTjQQr2D
YL+VY09C4dr9zPwf879LguyQTKMo9vQcRA6q5Y2ofTpiK6ps3dLvVPN4nhHtPiFx3yYzVNCVNfPC
raUVl128j8y4NrHTVqWPWjyy5ynpwzC/024/tbHPApJVPCpNNK0qSd6JOZ4VPupCrgGq5/dQ+O+E
dACg3ndPkBw+iKEr1t2n9xcAckfUa7TzAfjPpXyprMANQt4zqkxaKetQswWNAJMT1q3++tB59xHj
hGRLYUK01z7hPTHbWJI3lWqg12BbtdaxjkyRthJWBd6teWWVjGWQi/a9q5hJa/NMeHSOVfzu8/ls
TYCGNJ9SMt2Xrb1GvGtcdb3VDUjyShQKrRC9xIWeeVA1lAhkVeFGWU6AbdwOknhmZpOWXfgvkZm/
0GrPoH5p0YDUh4HAi6gxrJZ0+edvNOiyedFkhCpyLCTbQghshO5RGE1jGsK1Ac1VT/YwyzLLDtvS
LNA/IxC1Z6MGvpOIa09QSGxzNCXiDChtufuwqUdUxulAhKUgfjkJeareNAGKFwxXsKaCEh5RRl4l
eeU27d/ebghhTWUFBoQygfGqkziq60dybH527GzpLu9aNtSg4MsoYHCrT/IytIxoPqhHp3Et1x2b
vq5Zl79dOmwW8CRCrAHf58z7yxVqes5w/a2Fh4n9ohLJZvcb0JxdnnEvkiCjaarF12AXEyXSc7w7
kUqopwmTI9nrCx7Bn2knZC18PnExMNhbp05I7ghn/RMD02vbEGHe0Vcgw0gJ3+UdCVSdtx3GWx6B
GdXes4721dS0MUignFTaBzCDEXetM7pAkS+LR1Q+R+dpdtcX3B8NIExSGK5/Z71AXOm1aJg0R6Vs
SRMD5NPCmEFodeMuBbyC05W/TkKnqKbr70siz1AzlslnPsxzIKyoviCcGmkMX1nicZZ2d82osWoS
90g1vE2UijSzXZ5Z/cyi9ZvMGbiB9aAgsqy/E7/runhvsj//bnal+v4OmT1JzQxr8vBpxNO06n2x
5jvnAqnUAfOSxCmOGyYgOiFPmSF6xsOoMyPIPWJtCqkSZb5F5jN2Tm/nH5lq3ezkvCxGpwhTsmn2
H8JvZeHjGxMuMNYyruNOMAw6LRbHhmj7B443J0NJ8C8HFV4+JI9ysh8R+rorrM/F+V34a2BE+npn
U+drpMp3w+uYqyZHkkbND3pZ/I7Vzlj15YQmpE/9X6VJ7l2/fpkh0nXZ1IDNZafTzzRL+eJeesW3
ziVaa6iWDFQx85UcG9yGtQlB6ne6W2VJ5i35MH9MmUTzpm86rKK0bS9zd2g+bcmV2oQNPYs5ed5F
mYYleVWN1SAmhy+Tp1JLfVHq5fQyykzcFzDbmxyVFwEi3tkJQaQv4nLA/xn222axbjR1nKSh56NC
LRSk8w/bYmwfijJImFhbyu3FQS6JAWQ+rFaLyFVAI9UNTdb7MMA0swy5m+1oZknl6d0JF8JGrWpM
F6UZKZBKFwG8lisYJdEhUWzAUsT0n9q36KY0HQxmTEFlJGmEE3YPI1cFyiwQcCy57LUEIW5xLhYr
NCPHbFDpbusHBbawBW94l8xckwlTsySQlIiK3mPXSZnVTYLRespgNAOr2qF/A2maJOgknF1EwGSN
zuRAQlrkiQf1gV8wEUCJP3yyWDNuZILmjMQv/ku3GjS9kGa8DcG05C+m6a54YGJ4O0X+mu1Fjn8N
g9b2EPnZfizdy4gDpHs3ZYSmvEhtZkae5x0q57+GWYjmJwB03Qw80Itk6Ch/7M7kcSeaAqHOeSqh
1VXPu0oAdZdCj6MnPsiEH1Vx8BCyHVv7T+FRBl/Me3TVe75rCHMTn+Mo6qy+hOQPUOih9dyBpmM6
PJdQDzx1aVmXPkAP07VHY44V+xRkH35ZRrLj9SK+4OCzBQlS0f4facjGNWvK6TGs6j2Z9veThUIV
b/YVvmvxQGGR1dsub78MLOVLDh9goRoLfhTa10ozvcJLDRns23j7PZ6m4sQy+r98tyZ3XIxv7P7b
nRZZFovnQEVrUw6wS1ptYKqtL1EyB+ee5zqGkhXSdcMhW7mNyCGz1BMWLlPk7c31Tdzct5IPK+iP
7K3ZEJ+1rSQvBr4Z8Omd9/SVbLXqG5RtiRoDTrhMObhmcxQBps8lZuSS+yBR7luigHW6/KKE715e
wP0UctKzGJnLfi7blT3/bSKiNI84EvFFuLGFErbRaIfPSSlyDmLKiBsF7ie+2rF+NPn7I9hvWVlV
UiEldCnzS+LSg+5GCRuna1tJMbij1mRGoo1pv7df5E9CactS/xqjLg9EfoVLqdZAgglVGhMNgez0
Mbyd5sWeU0Oo9r7fu70GBL/cS1WzKB/wVY9scQWKffDNbfYsXESjVdcUBZ2HaXdX6aHrjHTkNU3b
tRdoij6noRO89nkgM5NFjFlsb1Qh7k+IFKjKmMUQ1GjsyN8rc1YAg0FQ4jo4p76QfEEMFfK6qcbC
6VWDzf5QqzY06n10/BPDtuIZk6JYErFQ/uxgDYBkFz4np1ryV09i1M/9fmW6llmUCvKwykYTZmV4
1JY3pM9r0kcTtWl4J43G6kaCxeQEHayLAuOVM/uFhm+2zt8UL36liQVjdZHJrJtRJCS1MrTF+O0g
oYdDcz/+g1BOhszLmPEq3wLTlscJEf5tWBHczBqNZuq24CxUweWwrg6Bo12Ry3B4z/6gHodOOj7Y
sxEhYIi9grsac/9VBmN/jCdJqwdXdijqoZ+qc0nztopuvtMReZdInPJ9f01XrMRPCKYKWvuGfZbq
W53bssPxujTjsuLFPEJa+2k3hrcUNZt+uuN0fyVSqDZPx8eI8eTKB3yf8GnekHsMrBkgUjQEd2CU
qO2lCxhaTcD/vUoch4W5FOcGz322uLdVTsaFQJLDuY9i+FpzWoZEPtCUyrioFDnWOHLc3JyJnDPl
AJKTavKhFRdEfFS82RG1DbLp1fz18HwPMiO6c5mudsutSTEt9msmTaO7883caz2yQ4lhN4i7A1V3
UBIx313TRMt1/8OxUQJ9OSJkkqxZzWKP2QRuEKnKPoFW7+5c/vDMpLeKgRwwr7STjh8qdowY/LoJ
dWvlv7b7aTBoHypo5gTxDMZ1V3qAI11t314mEzC0yh52Tr8VrZa+YsQpUAlHXRE7RR6wsCMsPsbZ
VXUI/saljtopGq4RtjwAJCwJFREnAuU06arCgn9KPjp29Y/6FO5lhCoM+CKCUKFPx0qbLH8fm9yR
E/U2qrT+tiH31z0sVsClt60TIFeQaaCaMrOZbu5sG7k/RWsKS3UVAAhZAZf9o9tqlR0K2hjE+eGx
No125Xac5fPJh7G7Bx1IDhF2av2KDHITZzvlKqUZ/QEUeBgOx++I9EsNiA8uDWI6NB2Uxlpms5qg
InClLHhBh0BHfK5klUrjelZYEU1rHYUJaTeAsro0GLMxDe4cwGRWl0mHIf0dICT1GE5yS9z4tmSZ
5vvAli0XbV/UfTtMXWaZJ7+HSadihFHp0VZWhMcfPEl8E6+ktJDkCorDMWsiBhC2k6NeZycLqHfe
/9fdDHrL4EH2Ts1NQPnQzqHG0ULhzwAEVZQYOgh5q9vcLVzY4D3MSuqGqFf+0tCykHIzs8dahcNY
4dllrvFLk73Wcm1MzJIyJJh/D2t5EhUrSAiaNhzGmPZU/J/4F1UtjC4oQCSKFXTg2QML3uRwrSp6
r+TTd8ZRNOiSeOPl2bGcxvqSzMWknXkRAVLODs4WKE168Oc9SdxKklz8aWZ4hV2Zey1OD2sOzc5j
4eVL9ruaaN24aeUvwo5YLdApyGmGMvtIM50ho8klWsxMEXU2QSzh/Zl/y/RgsT0BirfOOHl8goeW
7VACTiLWt/qhQdzWsqAMIuIPuleX8RzkPzfVo0PioMxaKVcEqSo6ATi02J5RUK9+IsaGga1LOcET
2pmNvlU0c5FQwUDD7+cvUldL53kiFB+nN6wRx75PmdzqR/NYBsoWaikSi+np8BcPEP0GY7N1RrH4
FYMbvgoR/WrPflDyOUruFsVEcKzoBDeHNpUaF77mOpO/jZhjeSrfin5p5BP7q+TzAGVacdtjZYkJ
YNAq79yeMln7+7tRhG+06rbUNI9SnRTLs3gyO5GiSkk1ur8McLNq0liv/oecIDsyje354tXOXOIL
bLatDdNw5THu5ndzmJ1pTcOi7uts+eeZs87qA1LihboLdRhnI8XdKiZxXccMtyaKfQbNJKvCd5m+
OuIZiJqRpdsd99D+IDkccOIEg/lMxXLv2hqZjzKlXEAsLV4wtUnCMh4vCOvJ/dMo9+lXRnBXwbjD
SQkZw3gcz8FME4oIS7g2imaO19kFe3M2var0j8uPD06KCx1CnBYAlM2zGE15yHv2srBAdH36n1DF
JSkEEURnVhTOo9UitwrSRYOdGWe9Vtm/l6qGWFd58hbgBtVCKUz77sZKTrWVw6SDnEk5vQlsWGQs
6fHkr7K4/Ha8fXHja1+7yeim5UqUvK4LLZro5cLJoK1Rxk9h6ZGeCVExQMBM4Up9/jEyI2n2va/t
AcN29W2WlBgfJEsAoi8aO+3+Q3rb9dJl+IVWXOn3ano5j2+yvokiMksEP6HX527EufzhrP/9tCmC
Pe/4mIwyemFit9FI0AF6X7ZtLPzTUj4FM5X2TQOPw7PuJEW307MNhZ2VRcsK4FL+rcLDWjaQ4DVN
oszifEFBM4kx3DHS0oCoLMULESixFBCtsvzRulKZJxYloqdRxLRP3EYW7pnKshtZyyLGRTCNb8qe
04/CYsJPH/TGx2qCQ2Bdk3ZxEYdh01Rk8VBA4Bc0R/3PsydQfEVAz8VBvJMxS3E88dgyDXQqDFen
Bbr40htpiJj3nN4by7V4pRFvlUuYJ+iuxc5VKIRDCwaQTbJ9izI+GMCzGQpNVuCLx3J6A+Dp9G6h
SpdPwsZxJtU9SRst532qLO1DliE7CUEXG0FIYg5M6e8GXY+3Mp26RsM2uanV7RYKF1GnAohWh4QA
uKFypu+eBrCgveCawOO1+lxrGdX7nkzPlBzE8MLJzOHJAAilL01pGNBtzinjbtLNGvIqTB3jbNxI
xB/arDwmp6ZXvXHBLIGMGBoBbwBwbJ1pMkk1QyD2EYIDpBO6MCZoZFTFi+Qb9tCinyM3ORJWv11R
hNBw7xZUyK2BfIfuieEiYLA8IogAp+pa/26Aax7AAVNKIsNYRRs1T4f6FzCVjjDAon704jcGbPTe
jC6HA+SAQ4vfglnVfXHloyXl9phaxNskeTvXQ1z3DwwTWLvWKfrBU+8XSFl2mOXCh7N/Np6nAISj
zBKGBumKmrEO32CWxdupgdr7DrIcrf2xpJxAhG55uy9XBcQgnyUr/1y2y/wnHlRTb2EZ2RXWlE9S
iIxu9XzAlPcd1dSdI5EOZv6zI3ax1EuqJA98rqperCeS4kw99K7F7SGO+sbre3MpLuAZFI0efuzQ
aCCIdJU+EgiNo6seAT+VulrYjVCf/ejCfIjePmSJ0yD+7XZh2kCJzovYn4/tWyRFIje10ChrHSdC
To5FZnfp0sSBixyrByIhwYe5oTKuZ2VPE7kjb6tEHvmO0GryXrljW3HRVkjHT7465rkWCxcuZ22d
tHtbZd8H9WhLu3siPYdrjwLt9eksduNGzPX2wsJ6Nca2QIcJXmUTY36mTJ9Y4idUOW6zMTfIgDbM
5uQnL8VrNeYfuOylKuwqDzO4roL8vw3slXORPq41ICF1ZVdElz3zgU3HrrWFI6esl9bbA4yfbFT/
kwI+wgCSgPoqqM//ZeqwqxvXqO5QBIR/mIzGLsPLlJ8W4qTBXw3E8nDz0hig+DXzSuNGNXRhVIIf
UKwOKNlKATeSrv4sUUe7+M4g98WGTB1RjScn5mSO0G6aSPOXZmVPfxbHSRgdUpr+9PoRcFgfJsAn
ILQ6G6xMz+QT62Kvy6wQosIDU/nokyjrFm7tjJEbAMVd7HFE3wLV/zLIVuhVafo4LKv6Ge0dtzUy
Bo0TgIkCpdDgaf4bJdsDiwtSUmiLOGCfPDlJthRrvxJfagPTIeOXVE9v40yvDPHvIrT8yF/zF21z
viT4P7KFz1H6IHBEAWgO+DU78s2lzgFnppszQd78x3zPwQ0eYsFr0mw0ahhN2ybwL+f8fVwGm20v
ihpVfliC4QN1gQG89C0Maw2Rb97Uu4fltmBSbzE0d3Dv/dYPrmRsXS4QX7TTBMT3nkkPX6wB694V
pKxwD2lsbOZbrilwdFUB6wRUXjziW5sHrPLjvWWze5NeMx7/yVjcNVM8AmYjHgiRdrJkquMtlbGQ
4g/gqefX2bDosJ8vlV3lHvto7fYBNQGTdyim4OjwcSKL3gzwCJf08Ip7fTx9XYVrbL7RJy8Re6HI
LotMT31FFlSv0gwNWmPuvkYHjFjSpDqYVT/D+dUZGrlzvDcyNS7u9EAkxv0aasRtDN4EsDV7Z4I8
FzDpGeFPa4jC/HcXuenbCwj7Q8rRMpze8rREuGPbrp8xZec/nw6CnRC5lLfPoSiXECtiRKE2B1VE
+wdlx7ovwH1JL0DZmNmsO3EMN/FhAka8Nz+ZVVEVRP0QjnmWkzD1Ls56zSdZno9nZX57lKv3WtzZ
OGf2KRa1sthg4TJRmbFvJpUIogVLRtljnhQ3oe/XD+mVKe82lpsYbmYol1leeTItQOHDT9Jcsiyv
tchcmaxuvITNsdFuoUaqQI8q44UXBme3ZTYA3Vml+nM5OOMJCJbsfKrIVghEQmPZ9R58PpjBMSso
bNKGI+0qZmYEfDsqxTFYudYaO+gzYv8TNzBHE8WnBangip7t1QYO5y4cxstnAhDDDq5fZBZcu2CS
ovF05ThCcjo00FCYca6jM1egngk/RVXIJWLHB9+euUd5fJaW8wDeE7yQhsr92EAHeRYj/NsaHvqU
GCzSh6XrytryUZInEc4EjtgyqUVTZ9JvdBFTOz2Dy77Cp8VWkAgF7FuK1NRt7PFjstKrAZN+A3h+
CIeqqvhc/GpD9D423N0pEvHEytPEVop4ZYnjzRRbDYif9wRpP00PN0WgkF5jSLVg7fvtdh4CRsfX
JoS3N/hiiYbAYsWJVr/br0SP7NcM4n4sOiByB9IgEMIoKf+OhbMp0z39TodMdbNohlW1+Trtm6Ra
viJo8Bc4Yi6dLrTyDeMAb3c2xyz3VcgkoA+sfy0f02qfCbc91fOEZo3ffwlDcveLwJ5CHOoTMkqQ
WoqM5XGmlV71uwyEjc/zdRfHyGHnAMHoijsIGMN1pAaB3rIRXCPXs4gLstTb7zz3uXl3cwXx97t2
tH1QxlyoVv/7u6Do3kjuxQ/y40tvtInHa132Yg2ZtamPHmfaCvykvbe7KZUz7p0yDl9t6SZp/OnB
RIewaz5FFVjGzsvu/POmWEwzkYR4DUfWFRuGzyfLB00F4icQQ0a5hYC+mBhGDl4/d1ewcFG99E86
jg5B9bQ30S9/AomwbAGXfUvCovsMHjTSwbOZQwWYk7ILv/ftJO4/xn94EYBL8OXO6q+q9fRmiC9X
8ZmMujPJXNpQzTEOs3pGdSkZgtLbxCtqJ9ePZtuVl13Mw14/PlLWV8Wpu1YuN6Vv8lxj0frvKd+w
Fty9spsV1AuGuDJHal3D6+syjl4evud1FvDxcLAikZeh211f0sDmZkKJibigCQsguZ3T2iS3uQ5z
qgjK5l3TT9Gd+ZV1NEaGhg+q/1LC7HAOAvbDX7N+FGxFScPn8n9J4UODkp041c2OKuGh4q0csQkH
V3kj5ZOo6IeUYzjwcpus+Gv8khVssN0uTz2QU8Ism0qVSDS1sSnz4NKVb+u1qWhGZSV5LAq0V7A4
M6WNL5u7nZucCyT4pG5G1yWK4pN11w19omJYxs1KfTCo9TgN4n0fG097XE5A7+VgzqrK8Bdz5o8e
t4moh3Reb1gBOQPrRoaetGxD2gB2zNmlVRR21Qj9TPGodswMpduMZAU/R04oDz9Mo8IrMdBXIx/O
pLDgw5bZSHawitqBPVgLs07cTBxIKaBPNNOfAB/MF9JTJZOhpTpKklr4+XTde5UQfO50dePB82V9
aAVsKFt6Hk5+ssNe1/WtMhuDdWZgHOU+TW7/e/WE02CeBEeM7AybZ1bK8Fk6r/pjr1skxCgDNAXe
uEHbsApMh3rZEuT1b3OKElzJUYqzHWlibWYzRfrmtBiIu3zijJyrBo789FsAyTK2hP6tTNXSebyF
gp9n35AQScUGR5WFqsKgnXO6MwqIVeP64LBeYky3sSFuV2abl5eu5/1m0M6nP3Fs7aLC3yOP+ta1
LXChApoatXIRZOkbQsxJSazWsN5Qg6WwyJtxIiW0Ee8S3vvO5WuoGnePznpX+LUjL8IqeuUPcvSv
9qnv8923yRFBpdq4fafLAlMUf/v9RuxgdAMOH1kGZdFbgdZpoNxjn2Oemvpv607bXT4B7grSrUh7
h2dAWL/70FCw3yV17npbvBB502+xhawJBP3mpWWbgFO/okrVx7E8J9oxVUiPGqGlQJcRZYj1Xp3C
uksQdP6PrqsOKAL/uQrnxMawtYA2NKdrJUBY16LLN3jQx+oKZ/0eSnUiVb6bL5RVzH1ftYwDDmbW
pmTVzlcEaEtXg5xXE+GgBmt9A7tzct4DBR78byyLgYF3vVaUdQjWN98Ygsq+AITKjKBQcnXcSTMH
KTnUe7ObLz3xx6dFNA5zHL2Bkv96paRSSMoFYItqlg0Op7NvxVEaOwCkviQBp8ZYZ8r19vGEY8OC
QYXRCtWb2vUf5sWMIfaXLf8sj1BblGAV9+Za4k1p7arZ4IKR4h9RTcFb9zbnU1y1WynZMVEzKTBF
p4Ib1YnneJ0fkBUgqfwYjLOM/6eqW5Cr9eszTf53lYS+CZkGv/ZORCgR6XuOm2juXBqQXdDDAoUm
BF7CfZb5Y4hn7froEzW1bJHERvAnUg27g5cdlCb89KRUc39H5mhwv2fgD9uL3NBxqWf9dFutGjx1
hVuzDtxzEcUszyjJp/Ghe0mcurzgHHMbVZX58omC4HJ85mrodWhC9Ae/nXpfI19y2p/ggMGZdvV8
SukbYEa5iOL6+rYlbfQpjgoahmCxu4+2mryKcKhxlckInzcnsc7bdGuluAqniunwP77y/kmpODJE
Jbune58v+axitY1SliZOaepKnTsV8X4nYx2Iu1GdQL9h357h5yMYR9f815Yqs72vCpq6l3OGwZM2
fiebZQ+JECa51xbFke/WI/ssImS+ZK7Uug7R5prOCX6Hh6bgijNlS3UhQC8vKjxY0VlWfNs1taXg
S0/EaaLJv+oYSUNRWOdY7FZ24sq2RC83eKo0t/YZFcfHZBFfFH+T6FD3PVk05KXAQJVyC9b4v6iz
bfGca/GBNH9PrZtuwNMxYWXeJadkd6/pLx8UU1t2WhlAtYXcLLpmfTjZh5X8LCsTD8h4VKCf0az9
ZObaXMQBFVbCVCeAQhVpqrMkSYTgDjFVku5Zs8QOiGjt2/GyePXYIA1wvg8zR1gvGjr8cUJPKZ8p
2oReUbeWzPpQcrRC7OMehlgJ4RxqnX8devNgqKhnSZkwrrTyFPLgGqV5eylBNr93Y5QGy9WmzOAQ
ZwzwYnWt+edyLbfLttcrsnWH78tPbC89sshUjzIKvQnqbpyUlQ6NqTPwHCcLNmiSz7q8sp/XcMn3
oLxJxwSP8OGo1qt/tEo167BIIBc1kWPV+sTAIarqwC8atrI7jev0zpfXvD6O0waNWeUjWV49RN3B
0XE/8XQWUrGevF8E64jqYIQtXTyOVl059nHg52Yo/ryOL3kfhTK17+XYrOW8JEpv/hTqTRKhsi0c
prW7avEk9hTI8O40hYsWFPQvqSoWBbBzmBNdsDXl335aisU0ydXQ8hl0v/U5jQYvSgP2diCGCJQu
qD1v/HcRE5jJAVKeqowz28chCGe+rUqjI2KdHWpJyhvbfPm5SjaekJ4DthBt33+XJ3kPW0WpcD52
c/Mdv99SotZTe+vO/E74Qp92mecT61rtDx0JPlBxYoPC9i/UJbSG1XCV4QrwP65qzbsjoO+o6FUA
2GTANoyEWeY1kUW3re3Agiv2cxk49umijCuggQyASOvceUErwkGj2PanaqniNoindwwGdtRVrNP9
MJ47MfX9Z8K/phGC1mzAss5Haqi5XJZ9A8ZTG+3BTZGwSFHqVo5r6Um7ObPuE+K/AAn1GDfXxRvC
x2gyknTNRqmh9mgK7yh96v0ekD6dpnw1dSKoieaMa/LX5Zj0GhTSI7hTs8NItESRI79Qh5BeXF8V
6pzL+GwOK8YAz63EvIYkUqYFswS/K3t+6UIfJ7uX4qK2jGiDZTknnPVO3X8gYcMm8BIm5zs6xCbk
r356p+8gnUVOmckj2MGyRIwazMIccQqcidWdcYziuEOKPFfuEO6XjZjWPSNRYz7x8aVdg7J3iHlg
sLW0W828DCLPQOPfQHuIqc4krc2QkM195N5o16OXZdYzfjhXoWsecyvAwitktF9jTEjBvrtO2tv/
+7YJr56McRDHrYhyF5iSHSAZlL/zx96mFqMu1Vmvk+YgvisqcJ7R4y3V75bAFe15yT4s5DMBckRC
FueN3FjEJ15OlnRO9XmfI2oVg34T1DfL5VZ6mXqI7ErjFSPuiKqsS11hQafsqUwtMZVmOgfNZ9Ym
+nBrdHhatX/rw2DKjDM2Gatswc5qyhZDGSElFrD8Ri7E5dSs3CY/QVRR8YAuVOjVtyRWA9bmDnmq
QwzOnkxRpZVrPjGLTOIg5Dqieh+Baj4GsJMdg24/YEdOu+3b5Ptu5FYO1kZId2aWZoJtow8702sY
+WN0hz0C1aNpWaBxlMfYBIq42ugbdUJaN8m5P+N1FmZqWiSCY+fKDy7t+U/DsyOHswjQxASK9DUv
F3NtKBjgRY1q1iNIgRg+lHd4dH7qsnDiPkY+dp45EJr4J0Dg0fnn0q/4odyk6QtI4M4axHxSoloO
GGsl7DProyR6lt3ACRDqNDheNRpq7FbYpJTr38WOKwWQCREwXeDpRLKvxm65NoBkOFEQE0gzaZj/
xH3rRcLyp4wvoNPD0IzLMg2jDSGSTexUOB7vQQykrV5ISba3lu+zLdFwIqHVxkz1TQfsW48zdN+Y
fIBeW+p3hBUUG7AMdrzJiyHD42ylRwwoVbyy72hDGKVqNW4ZxAsM49IBQ7jvltzKiOXMAyvv9j43
MrK1aCgTLSEYdcwxT8bOodl82qnWx9xJAkDzhT85F7YSppZshImQP/h5hqGZw/TbnD3t4h09Hn3u
XKOmct59m3dRrD1dMJ4CarH0W9Uapb/pFnk9QtguxWRKXO3h/m+zV3WC0TtbAfJv3dAmKUKUvvzr
l20dN94TkNG/Lxau/CkSdx2Ho1VxNu0ObbbPdmp5eu4IClf8osfxAH7gVTPimUigr6cSSrwFI15B
D23tXYYYIvsniZQUlIAK5lFRBchbbSvfbSiezlOpqR/KWrzCiojdM5UadTbK8O4y9Pegs6jPgRXP
KPSm/xtSzszpXpW7HBYVJs6sIx6qo5zRKedgfXoEWwIXyxAhLsvjPsPBbeZoRguLNOhww1FTZ0Ku
PtVsY/r1aGmhwbLaZ3C2YmFaKSAm362GXZhT6rm2sla6ur0JnHftxwOH8IDrHF6MVaBkED151zzS
aEeAll8va70bNmIN8A41873l9GpV4JeOti6f+LIqph6WEIWnRlTkNr8e4BAyrjzVisQMyU9aDSZF
MyVkzImbmasObxOSO1ZYou8bcLMP38oSt9qlyCvdRYP/T7zxV8IHL36+FANmcfLwq09gR0S9vium
nSI+X2cJ3iy9BdLq5hZTiZjq+KwObewjQ0+w8ZAq2/31HVz/b2zll2igLmIaXpy1YCzss9ssmWdP
DnYGa9eLwkUfWFMdF7xblRmKQSbu46xUoxH0zui2HuSaZmvFmyQkdxE0IcAQi+GLIdyIxK7LOKSb
e+lkgFGcQRlKbq91nA+EbJR6oB9H39pZFJrVzQmVUiovFuIs8XUuRUpxuL4IcBbCRztq0+YhvyHy
xHTTcYinKRwj0thO85g2ITPuFJjSN4L5YMITaz33xpYK55hwRdjYLkHvCpziBvVwD66pW15+LirG
nkeIOD7+qLIO6qnfoJyjxzzURIZmstGsUewdNXPMhLhNYefzweyeakIxBchIu7k2Pn/VEGIgPk7P
Etm0Ki+SSiAihJVtFBqxuDyEjRxDyNGPtBHPnouuQLCR/Oco1KCwG1RhNAuJ915ZJfm18JpekGf/
DILpFt+FEkKQn0V9Q5BG6r85hgnz15gWoQKAarjetH1SbSCP/ZmVW0DrU97DE97k5KLOfIx/16vg
0r2+jLVl/6ybf3L04ugm73tTMFJ8Y5PM9dEWPG2QMMSmwCE8n4Uk2v1dYTE1xv5jVbCtgBbvETkZ
1NfeQP6OHbKoTWFzZeoMYMnJ0b7qajltFelcLPUsNIYu7wS/m54IOFxpO9I5J+PymcaH93ncdKYX
7qQtx9u8HLIaahjNjMuah78onztwCF35tA6harFg1yWQqpUJfFpmvN7Q3K9S//s4Ddod6SiiS9XE
tmB43uzrLJ4N2Q4XwKQBCsllifKcw2y2wS+s5sDWdwU49p+j40ViUnSR+x5693b5xDt1o/+BOaeJ
M+DBzkBFf6fT5nsRcC4+Gzl5g+OqCToCzx0xXg6uEDc9dBzA3+YnsEJjnDbOrXRk1eYEoc7hpKFg
BSnLPMYzRf6ILIHARPjWU6vOGVxo4SXI8UPViRTrBjhgdP0WB18Ven/x44SIjbSQOYnbJsf8ulFv
Xoe9bh65vVQ/jJKr9qgecWKyj9Ri5MnSysh/hUBZafXo+4yT8j1rNDAtIP94Z3ZjdRGeGqaRsp6T
Fa+SYSvFSdMhcWQl4t6m33oRod1/eaONF2hKnUbtEux/PzoUhzNHI22OcPF6OYOFeXMKdm1dacF9
NOXS2ZQxFtWdVlCOMAbNJ2eZQ87XUJaA2VxHmJxplHlYvrxHKLhaOTb0ndrTDlqwnRqsxc2flmWh
lGyBDadL2AWQxNfxYd9zOGUBnNlZQaMUGgicmDUN84vRCEyfFcnKOJlSHA2SlbczDiWNvvgKxmTM
EtQdrkfqsm+2G2MQNSef3Gcj7sEtfnJq+fEfz8QGYjDq146VL2hfQTtAIva8BirEoJu1Db8gCo6t
m+g9hurHMnLyhdRkyN22gG0tKAB6Ryy03RXmxwbX48vjG2joYJyX/ssjBLiHL8qE2uK4XxH9rpLe
aY/ie+t8wJSPXcz2z0bIqTFuVnzSe6CbWKKYimO7RALJTuaPyjx3dhMxejPcYwQsip/CK/czsMXH
BfmG4wFCXvP0A2L8jIG4QYg+C0RDRTBRUaR9KdsvFCWLI2SgC6NRV2lZc76s9Hnys/Q1+F2PvD21
ir6bt2NN35dS29DZ/sAJ0ShSunDuWeZRy4YWwAFQSwn+IC0Z5XYOQedgA1EdEiZ9y8cUIYhPwtzI
ir9vgRt0M/kw9SQt17Hjy0pTMn2F9lJXCrqN0U38wr643jMgRjDCC5yHN6K1oQr5EwVCUmR8ms+P
GwiCPAHW14LCsS/Gs3KkMBkgKlKo8vRHA2r2ZTCBT7xtvD2BPFjzOD1cX/3/Dqpt12NVOnCBFkBr
MgDLRaRZBY3mOeIKAuL3TYjnKG2CqZBD/7SXUa324JQznruzfyz1MNgvzVdnn6ekKGdUi9bmS227
3UwqyJYdk2c8KFwuvP7UPPXF1DETzvsOk+1DSZ1O93ESzlRlRnvjz8ZgJmyvkIU+sqtldhUHfBDM
H61s/HWPeWD0YvjXJK3rZB3PcHN+SGN6PdJK8Y92xViaIbiYzpzyifUXeyc2WAZ6CtXDxJ09fCYZ
Zdh2mfUMlT7pol/C7wylpcz5/Gv5Ph8HNie+5PugjB/YckreCAaxez8Uv9YgXYRaedh5gwJ2JlWq
OkCoLlh5HQeXdmlApAqw9ibbC0wXaNffoKBFH3aQGFpzAUBBdPnR+CuO8aMZ0hRwNA7EjZ69V94k
axaIiIAS6OFSjkxXrRnExESepQOa4miR+8Uchks6NdHWOzQQSH15bdUUa4mTc54Fqa6SSELiqGdE
cxGWjH7GfpzOHmXlXQ43jt7lTUjf6Ws6UFYqx4XbiaBL1HPv+4gTRn7sFWl+UX3IYygKYAj85JYw
2sa33ixM33dM2S2WnU5WETGjMBX02umT698CEyhiIY/em9JCS7w7gbPlCerQFThwn26UbJGWOQBQ
TiyYveoa5CFwY4O0XCZdtbxY9/izp/xTkeABWO+MCC/cIl9Nv1BmStxQsMt+SrC59LT8HS3M2M7S
Ao2VGwAIq1XonAN1VeIOsddPwViIbycfOuWcGoWUG7fAUrYXI51KzIvOV0/gLfDLeVRWDgibgaYa
7/eCz0Ivz5YL7hM+YS8C1ws5iRkq5K0WnnGopfDbVbQ11taOxpdAmS5E6EqVceludtm2k5rUfyZD
cOf6XC7CzWah55AWNk16GOwiJ++QMX8fEj5GfYuQ6mGzhR0S/HWONpQ7nwvhDdQ94qPt/jOjLRX3
VkfgIlJyj5n5KCWWrGtd8DPVchIU+3TsJdkwe9L6hfLrPZ5A0C23+z3QuV7PM4oCk5kEgbycgrBg
zkHphyHv7yuq/Jd0eeGYvE7UIEChEugLjKEA4n8F5B4vWSR3i93x/NPmYguD3pPOwTU8Dyud0Ogl
Rovx/ibBwkPgDNZXNr+dDg3OKBPSHPVbMQArjPBFCez1fwLVU0dkcNbhmYCVBCdH6YCeb5fiXjpr
dlyk7NY0zipUJa62ZPJ39sxgbLYZgaIN4MrMmorxJMSXVVahs/3fK0JIjmhdjHzP88M2VwWDoTbm
JrOX0VI8PK5ajpzApRv1YB2gokURun8DPgtF2zMT7o/D6Rnuzd7IUbFchg2z+Xdr6nPyRRJMgPU3
yUkKPly4KBPV2yBux1bsBXZssgjyxJMBdFi3SdhigsVDzjMg//n6H3hqJtuY7u9QZLlVKx3oW8w7
hVBfiuVRJ2vYzyvxD2+elvDrn6AFv4TUYY8ZDqjB8ih9D7cIkHw6Lg3o9hfllDMDuHx94stlqNLg
T9DuOQFunxMrO049w29wJPkm5TRqYmuAiX8EKgdJ+zcH2EAxcQZfMswaHK02srr48QYJYM8klF5A
V4zSmwkXlYIiEGzxKD+TDm9k6sO8MybE3S5UJMJOtjOy3wcW1dpRFeYYV+vhXHzBdJKPgiVmY8aH
uHDZjq5QpLOzJPr6J4BxWcGDAa3ATLki6iCXg6iSrKp+fX8y3m1B6kFdKL2aRFpyt9TCtobDEc/i
k2RgyZXbzkPYWU7KuDAjOz3eTEOhFVEjSCO2uUr5/+/1atdW5Fe1Cy1+gWTzP0LkmkSEkpIO2Co2
TFD8YbUYwJeaZ8THFiwN9dnT5Ap7yJ9GT2ZqO6tDIFY49sPO12/1IByG+HvlP3T1YKTLgb+snYTh
oHn9fk/CVv6rptdgaZ2r1WUjnx8QyETDp1VSayvti+Taq3yhiKseOuAumGq3XljDiOiaQsUahPiJ
Y1tvG7OkV22tceRbqWHgbZyw6LzvtOKe3LaGAYZma40DAGj+2+eO9PBSS5LJ4BSj1L5XWxTL4yhH
xQA7Mj8eQgoR7dGA2KK1ZLmrr4sGyQuiI+EW6GOKnTAQPPhWHeSHe602GdvhZUe8IwBusFPOlcFR
QdLBFx1iUUA5O9iGHnS43ve0T8OcVxw+INxJXcZLi9/upDQ86Rn69fzKYT9KI4soXuFG6ewFqshw
XNgHOHOOPFex10gE/o6UGw4a0pC/R5+Cjz2QHj88MFUU3LUWip3fDi25Rchg4tZ2IhRkceNrAOoE
9dTQQc/0ZNDyI1fM0dkFc+2xYneTcY0+UGQ0MvVuHkZyTiZdDP6pe9Y+nARSxLXbN4Q7sBN/qfxK
voP1nX66AYdyJq7XbeNM/HOhh2auidJcUKqRsNMa9T0wXSRHUpTdJej1m/8iJXS86Okhgxcdq9cG
6afRFEUltdCAftLlcS8My/0vnA/gW5BmUcbBWjC8xVXD6ZuMG+6aw3oG3lwqeJMR19BCyeECLBdB
6q7NxSiT38hHgCsvX2CO5SHGKbd7cVw9knvupOqzsQVccgDEbOE07uxrYUQIdgUak7C0ydWXVzpJ
qhLUUwY0t6Xa7h0GMh2+b16+fKOpUulOpk2OQFGg+vO2mjFgR6ePCiRuV/+ZggE3C9TaL6VtT6E5
Oclz9Oz6fHFIv3k06uXbwAYyZlvr1k6d/bVMgdovdGCXoNSarSijOzu3tU+svAwaCPU3QcSsB+3p
S91Kb4fYcK4EAOMhRqCwMMiSj9eMM69vS2sRFhx26+mgYo2fxgdfUEpmaVq8Nv1FOluMu4gEFpg1
Ro7myLihs9CC/rNdF1Ih1QW3sehZS2GNMCAkDuLvJWdLruwpQDmriBOtQqDz37ypFZJ/fOxss30p
tM3otKcpDVY7XE5Cc3qZVAOiFvTb55PtoCfiarnOBplV5V1pErvuLRKTlstGJ2rAhhZYoIM9DjmS
TRN94PudRVxB7HcdxuEauoa+qb7rymQ/Gc8YKUGUplmVWkB02sFn4ugTcx/8huzt94eVs9Y0cRqk
MlEpW6lntijpb0/sXNp7OQVYMj4+UjYIom3OGJckFw6PoscnfFTWQtE6JokpZbKEYbKvu/2MZhv+
aTz6y5VRvxRy40QQn6GP8zcDQ0OzZ1ZVTg8BDMxGxnIWv0MiitpAJvyxmsvC8KFq3d4Bc4Jdz03v
sFMFDrSzc2+Kesjd81xGIOYoZPdtzsOee9JC4UN5JV/8KjqfXCT+FLCmMkRIXUscB8ctAuN1FxYS
nHyAWhBduMAB91EB7e/obM80gDzXQnftnwdymJ/SIs3PxHUXwg87TmM+pRRoLZ21LFJpuJ9HAxmr
Q31mmgIVhd/WYRxGQRmamgl3kO4pPxFiVWymxximS0SlZU7cXEwHs7Nv60YulSQpvezQvKw7cWOO
l6ApTWNQfVnBjP93XS8mO95tGr1u2GHg4NaOQqZltbe3Sfc+l3AMm1D4cXeBgaDGuSWCRilwZ3sF
rszoUuzFyrQRT2wunaEd7kPgO4BXJzhhS8ygLYTu2vTPaSBQn3ughJz3cD2Z3cBr5DidNNuiKqkd
RQ8RiWUmORKnht5QiwLyj9Q+x9J6jGR2nkceHOQnw/T75L/4uV3ISG5A0ljzB6Kl+zpS0vf69bS/
F6dgyQbqfyRt/WEdTWU4mHiUR9xARA+ze1Bq3+3LWDqC0YgSUCLD43ZJ3kpLcUcgztQkj2VwTKyb
oMSdjALBxQcY1dgzQpuKRamHledFa27a9SuOGewl5ZDQGoPP79ax+7K3/EhCa3u6aJgO2YLGe81x
vpq2PnaUjZCMmx+UqBh2clezPJdkiO7gAGhoc9S9+EP4qhOsXvZIp622dcxUnORt2hVjx33+bkUY
A3M42nYMjmQtlM3S6hfB7nEReFZg8Sc0YTaXF3LdkmiujeyQwujLObGL4Fod3qamUhiOQ39pFvrY
jmQHIngHTejHpcmzZ6TGvidqHQwv8wgzZT5bZoylNX6QXvC7n0qXPlkcwyE0ZmTFEm/wJHhdZMKo
Y77DVdP5EHOmNT/xWJSaQ20qy/JcMv879cngdUyBFJGs/bsTZc0B0h0F2rXWR2Q3iTvy8CEeI4+R
63nsTdt0JIrnyBVM5dUGDQW8vvL39LsT4CooLZ2//oMIFyrzYCGa0U5i4d2H2T3eBPTOfYeF/ASY
Zkr3pDfjFt+iUUQSvgPXatMwJDnsXHgKiV618sWDb25Zlx7eqGtKOF4iBJvuXt5kNOfnOiz/004N
GtjSwwCXSVtasrzixYg3CIdHk4nCIm8AkDLhvJVLaQOZxvzHsBDPsSvK/0kZUETf9QjfhcwvRSRd
h+zcpP7YsRVrmvJyvUH24I1UykVOJqmJwAv8cWGozCxPDH2ggo90ksfOq9bBjJWI7lFsNa855gpa
Yr6FUTOli2/aiHR7r+fnGSL0ZjcdAHF7X8yGMYKc6MxB/0e/gWmS58exIUEv2U7g7/0UwRlexpnr
logKkiXtUscS8LggC1OkP/GMJ8Al+f7Y3Yvgj2BgEkK4S4me7Sh/CkiWyOTyHT+2ZXLL3bP3IsvR
QLTAbIg38JNF7FCCm2e8qsb3p3d+fm/LeGhQdv0zUYfr7YKNA+/3Upi8fv78gOJ96kO4mhok3JNC
E2uVIhsRGhAbONfYu9ZrFsvYylMXnEO3h3t6mRrakDZkKjaBqg1pXoi51k5pwztaXxmn1WpgeFiQ
2LKee1clnsNL1TS7z9I3dbu8DWq2wNj8wEFhaPQGKqJ1qVNGJM5ZHwWwC2Z5rLPWx44YbJoj/8nw
76ViLpFlTh5cmTCV7GmAg9yPC0TazLKqTC807bLF8m6wkdHaT4KyWiLRB7kgUg3LM6T8qZgEBSq/
knWvM7BXTH8gDjhORmNPJ8vSC2egxjQa75BDrjsYh4vI5bk6pLqqNvO6xv6/pvCnn3mjjoJkPC1C
cDc3lvzjL5cideDn88TV3DBtctB6QUQkqs5Lk/Ndq6OaJ5wgvhYOJ86L+hf2ncFzV+2HhidVrIP6
HIxYMD/nVU3oq3ZCpp+AdACEbVtIBqLURN+izubgybydhH5AYALe7T+619piR/wp+2nzh2QCc2hJ
zx7pUr+Rg5WWkiAddtcHq9h3wTHGRDz4npjTr0DBz7QoYVPJwcOmCxHsZtNPfIOz04b2S5JCzpt6
3OOsPbi6+tkhC/BFpubjd5BELdM7YR+o7+VVZI507aDV/qU4R+bI/tXecYCZht8EkEFb8MIlq3O1
THRf6V++L5SoFmJNppZfm5gAYZJVFLgZILDkNVUYh1Ul7pYon5AU22ptxBo5dOxDrrSsiniVHrv0
6PqTh9K7bY8spgfbiy8Uj7CiqOD1bRagYZGn+xSXRfC4z7UvHzy6kpPebY3DUx/C0CWYtOU+TsjH
s89PxVOnYQ6xDpxjGR6mGn+P6xT7HzvmJHx5J/LePic5a9WwA0msD/G/Niyi+DaLzLAV0B4Xw8kH
8+ZvNTAERuDI+ehRBaq7ezjs+yxxqoaBqnkLY2ViXniRCBlXzF1AqolQr58nm80oVJWdIBUgfqSr
QAwwmhZusRfVIBRfDWE1kdbzlzTmjSVvA7XGFfbY/j0uDiQeHrD1WFtFaTpeYAAqKQyL/SiWqu2g
ZvHcmIk7ieGZ1/TrExT8jiBf6cX6Bd0g69r549M9u6wTskCNkeDU4YA0fFZVqpYENXtYIcUWYkd9
AMFWn0OM5hN+BmiZqxVnlV+bbGb0zPDNFoQBcfT3UOcSz19UyMy+XJ51LHtz5uOsbjkoTc3EkQU3
zlkqH0gV1f9nwsPCbJWmDETL1HgsfjEbqSbkljHdHDco1yfLbOTsy9rRZeplbCNKLdWt8Oc9O9mX
oZSMtmE8dlO7Mco3xiVZICmie9cBXSJ+RiVJjNfSEXVcNvXmgVk4BKhi1MoGbRkIgfng/Mlkp1H9
mUOpGEmcdFCBH0Ax1WsKS+ii0SzV2B4FMrZy4CZBes6Bbnzto1neOMTm4n0EJ4CMp3FvBghlOUjW
nYSwj3sSeqBd121ppxshG4KXwXWoCXLwy2jqfYEnXDskWvVAS0uwbQ3+151I7pfUmrxZgyCT8FPS
vYv18hDJrKOHEesL/kI+3W9HDuYf+aYgQ+6pW0t12SB9MB75GAmIJyk7XjkcwtcWANk7eXGXWBkV
QRiJ9LReeKHVOixAGLuOqgCBNwphhsysHIvwTptOokWg1BCYQxyI5kc0hp1f4PPvRmJChMfm6RND
1B12y2hl1Zd9Pt2BeoETDho3hMd3BWffGD/Omk1RxZpi+WvUo081pNePXRxzODhT+HeNTNAPA/Ba
Fu4nGGsDHymv+0u+iLzEV9PlEgqB4sCckayJHjzAxS0NMq0xO7Nmi+BToVXjjW5mdXxyPtvowNlz
2qzDmfAwl6CRJxthHzVfiQFDpGYG/UQkNNSYRiorn4mxdeHcFpKIcvE6RVY5qRHNaoxa3EPdyI4O
GQlbCT2o/0W+USrxBQki7jtVtFkYFcFZWmHJ6JfPIo+5QRA/pz4zwzezX5bFgKvkRLRnKXVakR/R
SPdrF5zNq9s/taAAai+AIIX5AwuPvA9FVQGMLx3zv64x3ua5Fwu50wpUJmJGUDMvunf21mDTVvp/
uWESvu30Ws/FvtllEd2DoEDzBrs0akqSDPSadtFcYXO/qDpHFivt/lIv6YZ0Km7lXJkIC1SuW8N+
AgVxw2E+DIAvei4bI7ZELiyX+xh6TOWxnga92kpZQIRTWpJ3INvnoP61/LnjcoeBr6mBRGvNMU7k
GQxNPL4F+/sd/MrUn+7uPfCoru2Do+Du3oYIQfAaPotjqAnRk0ROQVh0J5IQt5ZuMclpT/EKpT4o
wyum2V5O05IaMcC7c3mtugVmAZNqVs1lX/iLe7pvWKZTvEnUNt6Csx4+b/XwUNBB1XGoiVSRx4mi
e80SY/3oE98iTjaF9wpzsMRkQhE+rhNvyIlHQzJRbb/2O89ilIVAIKmMbmwc3Q==
`protect end_protected

