

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CZom0vHERP+sM9B2H0IfoDUsJRy9riNTVWFr3BZpkrcd8N+2GrPBLGYjWv5bwWNFs2qiaRKQWIBH
5SL3Ros2Jw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RCliXKg9Iz0QVLqI8b9GfxxBU1GhNUODWipyNqGvNd7T9Syer0VoYCIXvffp6DiDgM+PWpXEJgNC
ZPrITDndrkqwjZ0UurJqd8Mlj+O4jokuol/hbGtnMKDg7LMTP/mcm9YRpJxuqv5WE2ZWUtD1WAlU
7OzpzsPnbliZhM0CcXY=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kq4rQuO4iRu44woH6WSrRyNcsAgSUJbnevjDngvc9cypuoYRq4je1NTd7KtIptAfdlUTFMhOQTcF
fyvMO0ctzr5YXTPO+6ZCPBMymjnbHRykXwGANIGORUKHiAy8zVrLHGA2Tn1n2komEaNoM+u8Q25L
d17PGNi2LYc1A9ZX79yuNo063Qy3QX5dSU2poXOWXHho+u/vL1PlOKA9tvs+dS7HzKYxYNEywyjD
k9FyesJcGgO1rBPy+iEmTMF3cKMWOg5VxnjbUI6qOTjL5ZYgIsb5KR7Wy+RP+kUhXE6TZP6qsxFC
3QU0aGkYLyynNyIHyyLl9cVQHtYz+x8w0KmAqA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3w3EGD6E+efCt4Fs6HRylWTDMnbDGksrBmK2LrIuuDQNpphsT/R3PC062rFGmzFuJg/bLf5Iafea
N+aHJBb97H7ueY9YF/kPUqJvkNizbPUPQpBP/2fJ5zOg61lddHncYUooATB8NAF2hcSBgU35x68X
0+ZIEJC/w3FOSQwJ1Hc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sL/FJO3bDIPRCCsg2DyY6eC+YEqAvN4pdWi2+bTJiJBIOsoCbIwvgrvycADXfLHet65F7sNM/rTn
YIBRQ62HHXK4AhEPCYJ16a+GWujel0mLrgVipEjZe/PIBzOTjqR8RXDwI8IW2xOJhTKtdJhHoHnZ
fRLpK84QgF3/ft41vG+L+M5INzunmmeduLlvL3yJO7PaDzNzZxm4Yb6qxrxT22OrC7GODv7eJYeF
/B+o0KrZLuu0VxgdWTSijA2jO6/yo3BIW6TSbvbn1C7fQYmUfGWF6ssH9kJPORZ7fLwb67UH+6Wy
MDlUpxP5xevODOWeiaWV5Hs+S3v9MGrU5a5myA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18352)
`protect data_block
eplzQoQTiSq8tbNtWc5chM1W6JXRuoOsLeHWKJXzVfjTOXvKUK0dRZin69JvRaxjPVZOnKlYZZFS
bg9Y6c79lQuPXjBLdtMkclzqd09+eyoCTiFzlIW0ci4MPBC0tv0M9nJ+p9Zk7cAngNY5IPJ1gl9x
OnYAJsgQjcFSIGOCgBpgzHRBBy9zUW6clWy/JY/H5jDRP0YlP0rSQ4F0u37MaKXbdFd+XnAx4Gza
8UmelEvP4lGYcm/ldQ91rl8T/bL95QIZDwEzWFw1RCF8QlHFkXNGsG8md3evsF39ygINYIGMvEeV
Ls2ENgUZug8kuuAPQcfzKwkJKQnnkTVqv5ijvUHrOLWMSsre7Yi28oq+82tLreEa3Qiv8F9WT9zY
CjQLm57gkzwO5cyC2sOunHFDuVr5eEocg45MtQQrCAqStI7e7FJw+Qt5QDF5333boKPJAQt2DEwK
Vqlh+JR/fQi4PecA8rYltzdNeBfHuRln+wszRUR47Nie72gNIQSHov+435LAKdy4pon3yhIYB0rp
5s1yRcSYH9h85KnTtRvltOy+Y5dhStYUn5LZ4jLlgKKANwuU+4bCnp3jiiKkAepwcBfVpEp9lI5c
zz9wxSNZvoL1vcVhva3KoYzwCt35tkcxMIyQ3VSdw+f9l8XKio7HP8lFxXJVHPqzP/hUj7Vev6F9
bJqfXb12fHqvrAxg+YByTsEImVgRLjA6Bbt8MWyX5BH1/eBha74figpLBv//vJdnDTnnizUg5WFu
nyF19gxwcImiQ/cp3GHZtXPs9atgvQ1/CkWjK9THfwB9SpxyvcKTTXGmLRkRwGoIXSFMukBOQGqA
U5CdF8M1ks+yYxQVVoRZpIs3rCRM7QbAeYhGP06GBrH41zrYebhK8Uv8FeHodxtzwnDjwpdtwF4o
LvORpn5pj5b9FUWVxlN0xRxmr3wNqgCueYKlu/O1LBTcYBpMW6nNkjoNtR1bqalziHnBkSYn00Q5
yLjmJYQIYXXCIux/A/ShLgF9F12iqXmtWRdLu66uD4+yvHAIDxE+aUXNjiD9bFHoEbPZVXlT2R7H
pJbfJWfOo6AOx+tvpH0KWaj4n82pBhhs2fjIStnXGjIxnFP/qckY1s1TpBrcPajiekNEkyECGe3j
aDqN31+RXRjvW0Wkyvneq1LqulPLSnwWd6eUN+wk9JlPp9928z1VXUzXXy2sfUZPw7BODofTtJh3
8GQPuLhdOqddr+mcE8xdcV41fgUT3m8yY7Vieb8pte/5fBvIvhYeZZD6qv1Goid5NbnfYitj2xiu
2Wp7Uho003N9u3WA10pMInxWkaJO2VnKYIhoTubSFj1m5kQl41GV7fFlldVcha50F+8ezMqmIRpp
QnNVSphFH3KkVdmWmH/0km3jK33Z+fobEC7aSkCg37VLpdmELS4MzUkiuiGRKaodsUYhzCoaQOws
sPzEUVbqCFr5Q1HBlMVbayLgbm1rsXDyPcD/5Bh9GXDZXI/gmeIs+hlelZpflGU8bpC4H2i3smL/
1CkhxNvWZLfg7lrZDpjwkmOtGs3NXVHcpuKY5Gnx2GypWUF06nuPQ+W6CYgx7BoNPwwekp6iblnq
tpgwG//K3iPQKzTBi9OAFbw3hozxamDuLuuDpL9D2UDU/NnxjlEjMyNPRpune3JgjW1v7+4yyFc5
G/eRoDYg0EZnCVf1IjIKCLGE5Eq8qKZuO4a31/LCESpQ5HrSJdgKjA0LSQ1K/fFEWQ0/RUkEthIP
kX6DzFdU0BiwFCN7SxR05J9xnuV5o/XgywWBWJQl0WxhUsYgzqBvATWclYI8yDqvnq69d+C3o8dt
25KRkaLZkWPjYK207BB/Szsh03kiS2f0MI65GpOmM+syi1sDgZTWYj3nQoUKw+JXksnvjUZVIwgU
X62dJ5I2dVu6FVo0yIwWO1zhfs5nik06AE5uMdgfU/umAPada7RPDHhAypncWDvn3OM/HU1YxgrC
6FVQLUKZFS/2VKIM9LN8UN7QNEdMUONhXgOnJZ/gqq8pjIUqG4TxrVF03VjzIk3lTzZAnlt6l5n8
2rC2dBOucWOamqGIIIW9/wW0+U/4vf5rhlZX9VTzIb3TMM2fI4b0dm+/bgUnjeSawJVXagdm+Zif
Y60NUdI8waeq2TN5L1kOl8hZtaDdtT9n+LMRsZo2vpy3IiBThH5NqM/clNZSdzR+CcA2e2oARusF
sRs/yCJsUN5qL2IRye71isqeUnmxLdpT7jNKVFToAY87TQnCvlujCdO6AiSs842HY58fKBcTyYSo
BPNKxKfUrN/mWibyAXp8d/ni2qtp4cxm2mEhCBcwNsiX4+UqhE8Tbx5tqiDq898q7BzUdo7etW3T
6iBa4P1vp0lj7A0lEoyj9XNxIa3X8VQiCO8mM/PMPH2aRW79vHpcI/zR96RYwOipaywnc3/FAdqb
24tQkDwPrgJE2O6AzsIWhj3Xf25zi7jfQu7RzA+dgwDBIj2jMpaQCidQXU9w5BcxsogQer8JUU4E
7nOR4kasOunFQN6pgNHVFNxoveBddp4F9fBylKjMOn1l4nsjgN1IpG0LMSOYs3kalDjD/Tnw7Oxy
9x7YCe8uonMk0Q7Nnb0SzL/Dgv11UxJ+B/TKyeM4C4rxC5idpEYEqWEKM9lbSRdXvTH+0lWRfMv7
T0xGd5rXpwZrL64XPfX1NCCZBBbSjSJWovJqozsFENU/NPFAAEMofqE/k8X6sE64IvCXyGrQFbue
tGagKJlfQ5fbhk45sG7ln/7FYT6tu1Av8kDZ/ycplKneENZYH9LLlrPoOb7i0At2H7koV/lW2SAS
HFkFbUIpeysTSTgPp6TzQZERvwKqHboqYggNqAxWCV4c914dAM1nwK0JSBSvPUvQ5NJ9tnvu+Py5
U4EITSDdYoVt7aPvaLUqie5i2L+8f6AWX5iKIe7pssTvNobJHPnB1ScWAb93EKgjvpvHewVbF3LQ
ikKKiOMiHDjF/40JxP0HAtvuNRf62TkIf1yFYY4PU1YKnucAIQ8jZILtWnJAFQa/J5jpV1jbBdz0
uQ5PtxTiPlOlcoqy7h79NSXH5VTlttKWQnySG7jSDN0uILRU92TWNusxHc+/ZPgHXz4sUHM5oekj
A37uVGJoHA+O+d6/M6XfP3GBxKL2ubwoUh2oc81Ly6IuhqsDpbJGrXgVaIhESEn2N3JNr4W6ggqK
0IsvZGA39ixV4Z67wkHpaV/XGV0seMqLy68erQG3ac9dZQoraljw+Hra2OgfylCDS00+13xCv5h/
OxJ0M8RyRSvyEPQXkVFSrBurpEkVhNYDqjqsO+N25YIq3N8rEVKSgO8EDpg/UGSgFI+LcNA++P2y
rQ0o+bK8ZzD0DEFjsAIkjNReh22C66vIKYyqW9lEemkxHcIlv5mCXJdLa+bZUIkQ+MzWykcpSQos
xvjfJtp/iYNFVf15R9476hXwkvzPWpBBpD79Hy1/H/bLudnr0xZ1ol3oPtc0gbjSUZYAG0sSGxv5
/33eXQGC3spe/As4Dsp73cFt6DMXzRq1jRTJ95/5A5Npf7D/ID1PAUJt6VYQHkvmak1YtImFuA7S
HbSlHzHoMHiiDlSIofHNT68o6X16Lndi/UZolRe1qmjb9RzOmKfYSo0L9wZA2qFedhtmmKtU5QoV
qhDJ4V98occPPVIts5O2EVnVcpAXS/H0g0wO7wzkyMdrdurNIUKzaajlCNVYGlRjc6g+Y6RsbL93
cFGHAlFik1FFQqi5fMbQXXOmic2GmzhPHXGyE9y4DQNenhAnDYiMTD3WV46EpeN1aRpssFBxuoCz
YA/l/uLewuM8bO5WWSB3XDBVviDUqm7IWPf2TM/xoXzNxcY715JzAbfbuEsBiWkMQ0S98nDeztm0
upaN/1v/LPW98DVkHS0yuxuTnqRVeU7sHrskeydDzGRrnduPlHJ7FRznNOEEKWsINIwd2a6X7AdY
DzMhIA8bY8gIktOiHWnFp/9BbNH80Ra4wql6RMAlOPsugoS8NK7Nqalj/P5X9RDsk3I6i8bI24X1
70vlBd6bkLEv/UAcmGecMHJTGjiNz/RuTtYAk9vBmEVtn7WSe0FrbW/aRR3+/BNghvM74UNPUShU
S1Br2VlXNvCMANUDvKhzY912r6YOTVChYnSM6WQJMih7lgXY9UwGf2rF3Jwe1V2i8i0d9GjpHUcY
lSS55jXh4JWi4qyxST/he9v7y3FL56SMXX77qpmELWYYHtjuy8p1OfrGLvFM7casd6uBcA11lzyt
wP5YNQa1UottW04L4EdGE/Ui1VGgMhsyYfkff4gEwf0HRixPfFuwQDgXZ2WSs6YVo5ZkzRd77kbT
oQh1fi4j3eliOzNZtIGwj5PPCxNUO6DQrB5Cvb0fQmczbnwHj3Q1IOZd+yCYG53Lz6Y1BqejGdZJ
6p3epUKHQ9h0ifr6+fCsrCEAoogRqEJuWf7i7m8bkQu/RVSZ7WQrwoEOYf485EB/8sauCkG41DHe
vgN6jF/2mYImgiIo86O53mwlUvuBzm3BDD/R4qvXTa79yhmABwl1QfaGC/nJXaoj3mxURPIbdrN/
1PSwWdLGz71fFzDFFu5dAE5GbmJ3vvssi4HimuQVs6jSXgEROkyFmoxAhEk0rCLGgfpoaJV/v+fP
rqAXlKDB/i1Nfo00FtPPA7tdeSD+JHR0/eOpkFeibaDqo6nFISVV8gsM884QjZsyNQNHQdDpZKBu
g6QoUgH45ua1PQzV1pbjrno5ZXDDPN5b1/8D3zXbRlg2a1KlT5awUP0MrzNHJGhIzLqOzlE8UUna
McIubQJ21Td7I3o1K3wYm/Z8O4yh6eWR2AlfPCnuQBhuDTMI7w8etVuf81poMa5oc9pYJPA2MHdU
paejCwwyJn6s3h2MuAfyZ1FzMpMffJ6YJqEGAmu1SOcUI6AK7ZV88Uo5vL91p8wYMSosU1mSpHds
Zg4loQyVDGLpGkssnPGvGW/4edwcoSA6YMGYXlwCFi4VX1abZRJNfWqWcIdbf3jjmxzfdBk8PLhM
07uqIH1PvRTCBab2LbEPfhFD1csDbQjDgHJvrNVS9niR+mY1m/wQm0BhPQerKqEtgHhK1lvoh09h
rN1prunIiln+xoyWy2ePjzI7aLjeLvy4h/c2/4T30PgsOCPha83rGfC8y0bYxeM2pe4J4z2gUahV
Kmjok3Ch7zyIZ4JxmYkI3wDiNr7lSnUNK9bOrK9AWiX02vdDMeGdNFEvNn4pdO+yATdbRqxX26zC
aBZSZc61Aw873ED+6j+nFJ8XDOpwnM++7HBqRzFYOOtB5Q+02PtNvtnd98MQsR15A8ojMxt7f5+O
Njvoed5epkCywnUWlYAsww19mliRtPqMinNgrpNOVa9qPF3hdRk7EbOMTz4VgeU+1S1I4LZBQzpX
Yv+DNvyqHqOldiRVNjw+HTQd7Frli0WWhFbTGTevqQd5qaDGKgpuCg+6rQuQk3Q+O/wN7USMnFvS
Noc9WJjlsAJWRLEPBd7YeWWclUX4z68EOGCHdjw2T8pvvKlTV+qvGad7Ollcq6320LPdvippytVI
u1uR81PpfiC33baja3DUc0/UiZYxJcOgRSoKi9LfDScbNErs3nmQOEab+bbZmgBDdOhYwUYxsZiJ
hWK7jSpaOnpp985IXOxnPk1t4GHsVKGU8AYOqNqJYmweVtk5hwRxEq8U0RGhpKNFO4o+TNJe2GUf
r3JOEn2untUf1LdVRlO+zCIU6dI7+YNWin+WLQnZUGrvTbdA60GFh9IK2iRxaNZjHXR4UcK5Dn3G
eQcHs6w/ZvYDw4/PXKSd/5SFyZi2VmY8cPBbdNbbS8oIq0WS/26ikWGBrRfdAmnjX3N+7PR/JUUl
SYolwG4iovgle8IKibO6q7cFyV968WtS/edYA2A9F2Q21oVb/mUL/AlnYAGu9HHra0EK1ih6e+Au
5+LLjaKmwfgpk7aVHmwyq1f9cY8zKPUA2cKwR6YYExJXFNxnqXWJ7qg90HdZ8bvLb8BVfeBnZN80
5bdIKDjTofDdClDtX2DRZZy713pJbeRHP40fSCPQaaVaF5WfCgNs0lsnHZfzfDRIOi8p1lH/+7Vx
tMLPIsUNDw2VeoY9gjY+Zss0ehXpK+l+F8ITfcla6qBfvnqsNqs5bMRLbS7vcQc6iY6MUk+2RigQ
CY3Lhx/AaP/9nDLT7QKLCI+YL5K2kZ32ErsfGeSNowYOydT6s2Rk7MKhSxEaOxiE5dsHw38SfL11
N2Bxv8H7287cmo+OA8aweE1cGngirMQpNGyRHGk3TQ/Evfek/tn/lGVre7ml8ENqLrbjN1TpDp6n
/fpptE1tqbYdFFZ6oPhNneDnXua+c6naY+dqQgioMxOMaAcLe0+wkBRXmRwtZTr0fPr9wdwKEhlG
nVSixOIGwEZLBA88Nm5DFR2ieS4tYz9vpGX0AN5ibbcD5reM70Mo4wu8ZFyB7tIoUFEnLdaXkwwb
+oNd7zWpNmOh9kuVw985FTa9F/JRnw3qYfGGFnq7MYlFbPtME//oJFTJmsmTiY/tiD21uyLfE5PY
kugyZhb157SXI6bbgo3AgPAbXicENPw6MqL5GLc1o2ah6gORRr6dnxwzWbcHvUlwuD/rTA6o0DNo
qKs710bMrW2XpfsdAiMzcxymVyp7k56SFvcj3rfCiy//DF8NM/27QR6NSOsj5tv2gKgKi+aj3bAq
KIv0t1UJyTRYKxmHg+3uO+MWn1h5meUAkl95IZM/9tyJB3RfnBzwhXghc6QgDoM3J+1c2/OxITcC
i6Uu3xQRH14yz2P5zTMitN5k5+HOfe4qUvAaJNS+btRPJUAV/sncKnNO9rFcqA9huKs0Du0ne7BN
8nzDGR8iBRse9EsWME3K0qUEduJ6EkwH0JxpHKYa65Rn7NYFlzIKvaJECXOQvpIjOIMOyAwCETnv
KjoLk2m0qZEtXqgwSrjePkN9wMQvVLEH1SgwkzMP0j7heyMVf2HPKt7hwJXUay4k9CT7m48+EdL4
XRd8tuBJbKTM6xB0GYDrjbI1z/Sav0NLFcQv+nnlO5wbcxoLIe1vOo084kLa8apmvQ0OntR81Brh
2IWOo8T3NNHcAghzF0iXgzFh7HCZg/lAyeYKnN0znDw/9oYDOo0mMVg+wl/LjDzTELoo6vCkt9jy
U4A7qEHlnzaHI3/0BGVzi8v3OVj7uj4SVjpHhZZ1fI7Iq+tcrtvhrD1romr7Hm7jE+YEX6p8gg6i
u69v6U8qHAF/uZOAOlAmZS8dteKOtOF2VjG3VTSH8Ba8YncL1gEZdWFJW/Frz21n1h7a6LunUju9
1wU2AXBhadjRh75z4uZaq1Qe0WjhwXhABGG9zsrhj0krLWG0UaSXk+utP7+PeQa6nkIUJgAH+rmn
hXxXcsIkUyJ19kXlRKPOD2dkeV9PeflhR5O9hHAxpF6wS9Oaa9QzpD5FByDEwuv/FHyy7VS+R8ME
z1SvmOm+8iPvJDpAvRz+c5DmHtyZ5RATEWD8WC/92yiFA/QxDdlScABT7vw1bcG/90tqeAH/1+6K
D1wNxS2XTH/bar6dCykUJC60wSD4fGgeqhVhK44Cl7nBJb1i+X5GEZZ8RESSkTY0pVrQ9upoZlyW
tVK5SC6BVz2/DajxTShcGBiBfZK95TtBipctYrRLVWCXZ2jYHM2Mid1JY0tcjBcjl2nCrsQ1EIO/
L3R5665xRwzF8OIZCShyF0Yake6Tmbz2zEXt7yCwkZ34DmdCG1C9mg6iD1x7sbosECS5WK8Ail9K
zAS8X3VM93+596KcKSBTXCgD4QZ2bXoimc5P4DR+XsASARSOH4J0RNmKppc8zPunWy+dKEImqQtW
W+RkAVDGRhECxrehkTZUpKOpRqvnMHQvn9pOtrUod8Lyvw35NuNZoQey9DVcZ7ulHm7HrzZ97WOa
JdfG80nMbcRLbN7TsYwo8AeMFSO5SjmLQKO55U+tra8HVwCUL1Kn8NHTFipKgCkbXZBkcNVYxUJh
4yk5fwBGjJ7fMdmXR0gI9jz+OcaIRqk8W4srFp65/JNQdx2u8u9E6vLtu0NY7GbjQSEDS6FP4r7q
8yBKjCmm6hAv+uFhQ8w5G2AbxEekwT1OKpqFcln91p2tezsYhRVS0Eas+sGzy+hyCDWzCS2H09Ep
KiEWDq7FJIkhJQrMgYtdUrhcppUD5NaMWNnuVUudcbR7CJM958hUeacHeN5qjm2tzh0hrkUyqj1P
OCU8VVCdt5KBUgZmi5BLxeXNb5JMlY2/jiiWwfHgi1j7hUumhT5tNZoHZPgN6616nl0nuekOpRpG
7/ckYU2WBqAUADlFPNJEn8D7xY2DQsBl2mLJXc/Sce2m8+ssVfJJOlwjq2z7mUoCwerlf8e9busH
XQatMW9HzH1z0AwSMd+J88GzaadIAz7rl5Kv2pQHJDDPcC9KThmuLJQ00EUiixotP4ujntmMhPVw
bKhSvj6DyvgTTZGtY8eKTsVLqeaoBS8S2OQBF7nHhGNL6Ukpjs5n0Ub/jpTc8vJqKmAK1EafPlLx
KHzF9XUqfC0FqSYk5uL5YXf4ur//OJhT6+QKEW4C5ag7kG9eTKQf2KV9NkonKQWvTzMp077hvlPG
on09KoeDp4YlN4hLPEfsl13pq4jL/bsOJhaXsDNX/HCHaIldFabBQZtR+/kCDJc8Xkytce+OKuje
YRUBr02Rqr5cV4fXpQLKvQOcKcgEARyhgMZIhClIhM0i3uPgyU3KcGzXST+pE5eiFAkIcnNBmefa
aGQMHMPMb8Awk5bJwJQ4pn71KcgLDNOl99Zd+3BWWul3TqSowwyMObMNZBBmAWE+7gvXFDRwi4G7
jd17xgjlbY2czlVfdIEaizv8SdVMFr0GzFV1AnZDpdpA/xxF30JR9CF4d1lJ5JPSrn7Y26OoIMmZ
jMHnBZygsg+jg6h5qmgJuYSal3rJlEJ5m2P3gpverb0Ug+bcfH748oqsvMYq8S026kNUf26gpVFE
UOsBSD1lMI1VohurSdS07ezZejG1/iHwp6AXwcLpFfwYHo9y8krP59CkZFJziM8iqOnC85u1iwpx
tAmNj/lECpaaRqlSqC63fgq/SbjMnQdm8upINSR9RPM+APzHWcJcXMLOECJSTdxSSzocYekklZ/n
CP4qh9akrBXhYUfBwp+kQfESRriNoUWGpt9VFqSfUa2LV6a4j6EKo0tlgeiEmkpDpcSJoSCZezhL
bLmcc/I0G5be7RySoKVbMhhglpyqYxeAe5plZOY5yJmjxgpmtcEhrzK3g3RmUzB0xTEESzoa970M
J0Lo+XNmNLLyGcsD3EayWoW5LoAfXPHOBpImTT0k1WlfECnTzF6NpeU4flTHre0o6mwDpKMyvvsQ
avxY+WkzwwCgH6Bm9BCYJExmMqc7JEYjWEz2vhvVLYKQ985On0L1+pWbtTqoj7AQkYB21MprXgqS
iTBFWoJ7PmzMIYI2GYGNDktkNs8pWV8XHR/RhV0HMFDcki95pQGa/vSewy2nwV2HFMz1dV6SH/Wm
WkK89nQl9VSfXy6PFUuTUOA1Bvku+ql8o1GrfyoZY0tOCh5ulm9ObBQPi2/2bn57m3/UYlNmq31Y
bLusChQBW+8VvZ//i88QxgR6WwRZd9C/PXdnLMbsq419JKT11dc9TjZhNSR+U4jKR+VWWnolC1j0
GXJPMGYIyXwDsN6/T3Et9K5UNfgv3TEBvf+CIlqdFIOQUGJNEuZa3B0yE4BsSBI6pVR2NxgxYMNF
37jRfKxVgMqhv9LdxUTxtNNmD6iSqQdikrY/tPfCbnAP6+YBTC4SkmmRrweRjQYVEtU0mS2JWx07
RSdz2U//Zsj7+/RE34QGDhq8UeM47Thx8j6IXwhRE7QKgHx1z+1LHMwgtAdhsrtOt37MWgSXN6rN
O4eJdOBxaXfFmiW0h0mL1Dt5lobVzo8j3MTetX29V5He8/44abT1T0gQgu73zjamihAf7GPlqYhJ
qp1yv7kEmoVbO2KGWldDOg2ankxF/5/TV9e3HMRO2qGS5h/UGX6oSmhRgeP8ILdOuxrZQHLYpFei
KpanvTIL2mAyB4LR8XnBku/so6ZFBqWTS0rOogqYKupDoMZ2GjPgf5lN+urdUpRdakOfydh2pIm5
xr8aEB+kp0NhWEOFheeBF1Zq6WvkeR0aviOUYKINtgIqgkQ56Vwd8s5WYYXpLmC8yiv3nOBaGjhK
oYzRBSrKrkeATNoxh5o8NfPU+dRqW2Mb7iX5iZoTVyyEx/BcQaFmU1J3E0h4oD0xrxT9lTpoSMvr
wvywkNkAydXjSust69YL5l3qejGti+flrrwZFIWUJMj9NjlhP7cEeAqnGVtC5NF3diRkfB53luYb
jpXcObmsBetNgUAKEEtl181iN1Ck92+EUed88khcbdT9Vq6HzcuA4PDDlx5kGqIpRx8offwdwpBz
ceGl52YuLJ94e7/kKzD2bdiZFYOPSIqBJSwmgHi506ttM7dCidXl2CQsxyGZ9Ic49m4W2eIultQR
/6xq6qLXOtmGwQ1YlUDztEXdt5na1OBGPz8gcQLbdKBTna64e1j8uXCPW+LNUvhHKmeDQ4rLk8C2
KGYq0EMX0m6vERsnwidPPytFxfeHdqoL5v3anxAZrXJJzY03BeEflA6coBDqs8KU7X/cHJkjUkt1
O9qJXn1m+0HlsP3cG939XoWJG/+9YLLa0HW9WlI/2Y4ZxgfW9iKfrQvZHbMfSTBwDe+s7xwuTfY+
TorUx3yutFX5BErPbRtbwE8PIvaS6C/Sh39NG+uXNJX7lr4LP3u2TnJ2H0S9Y6R6b87fBRtJHOuV
kjcpSL8Zs5ahfg655evxDSvLXDBvW1K3pixQFCsRtDUwxzjHrAzuu4V6DjeiBeLF9y8F1hcZyvkz
GorzlM8vFhjdDKKjmEyusVrtRsTBPgHhyOEsopqYyh1SUcbK3nd+8UJWaIrBdf9KOUBVsqlsBnqr
/ApBiPfd/xR3qG+BWCoziy90Mf6QMdQh+WBe8OIthxNBCksFmMMWVc3fSOYWe74g2SWCBc2OA58k
VWGdCsSRFKQ2NxMGmDlbfR9WJMvbiqVsXHONhC2t5fj3bkz7lox7ii6wE0X8+tbjIFEVvKqTpjvR
RqDHBEdnfYSFubKCWtxen5ApFJQ9WvHoD9AKRn4GI1OVcDNW/khc+UeqNI0Et4yetc/MfB8lYI6w
/69F9xeLijmkWjUcVeGZFmAA3qpp6TR+YFu3walwGd5GWLN9Qow7jL1uC39xOhk+14ihNMrFlI82
srTQ7y8lo/xkQXe+QRakJpMbMTlle1o8v/zRECS7otn75VdFBaqXzV5HpGQkKxYaBaQ6t9qb/713
gjcHudTJa6XW0uyEutnkx5X7sYzlQpZqoH2EmTR0UOMuM5qJIdEmQyctGFnfJRHZlVklxA3Gevz4
jzVVIrMNonI23MhI9JACj9iSCBOuDc+bhyFQcx14GBte8d1bP9g/I4cX1Z+IT3XB+9ZxKmVwoeBg
BzQQQ4On9A4zBW4VQQr65DgU6306cBLSCx+sOj6u/DW7oG16TJpdBJmNyecZK5Ynqb+d5+s5MGig
y2AM3u99bU0UOHpLsfK3Kr+ItMVMZmwAw0Ty6I//v0P5JJiONVZtF0DcT/+3Eihqm2Ix0J4KYSUS
HBYEOWpMDaN6HICNZ82md047LuHR9NURuwvlF1ioP1GJbeZ8yu5z5RHkXG4c5/189YpE5gvARzJd
WqXAjWzg0l0mkktpc+GOivwbqrCOgrWc18SshUORrU7VFrQV4AG5NM09XQgos+Jk+mY24ahYBFK8
mNDFbcgzuaUcHeMfq7ymICIQvTs4kXMyz8MSyxET69zEquEJi5WpPz6Twq+r8OK88bDu6ZGCrpFo
pvrMQXoa/1BYwoig45NOYdkVztfSyslUtjRBvSZ/OmQEEa+BmPIOc4fXSkbMMf//Z97lgy9RS8Lj
/bCbM/6NJVVZgNtydYVpxrLVeau1XVK0YpjBcdEcXLW+MoSXGf+bq3/JCLTxpcIm4mdiTJRMAj7u
hFzmOfDvXQHPxnNyluRAN5mdECSfcOjjhtAzRp1k20VkouBXaU2CgwTrusQG7skOxJwTbXcKRaHJ
pzZ/QMV3YtrWpQasZ59HcThG624aidoykjtTg3d6BOx60XrFosMAxOwCo4pBqgg/sK9yOwj7Eyqx
oyU2IwpTC9wx8QlqUZJPHOUFmpKr/3T7tZQECxfqHJrm7H+fx06UwtemCR/ymNI0OGEbUWwU2wWA
+0Ae4Wmj2Pbk1Hofc1G7ZJus5+7A7z8xI3/Tlzl6ku+SZLro4GruVCtJuUCnkKfRI3t5W28huIrG
zIQKyGi00+zvS1+BaTaudnxmyfZw1wSB72N5EjhDqrRVgG/i2Izc2Rx5r7nNMMsViVt0GJ6tezq9
a2mQ6Kh5GIZvLUTiE/tof0+0LSLFckhqBYwUpyVSs02ubdJAgsJPY43pOngAP0P87XRiW2A4yK3y
GnTQ98acAq5vYw1WEH/9n9thvH5sR4RaNpoITy2cyMam4Kb2exmnD1+6ialw38N11i16mLYEUiCb
7jYW7eDsmh+MvwIzGnvLMMUoJxLzHuNz01RKX0xwAN3Rme0Blodw2LUZU1+5cxrjchWH+gf1QcCR
+9PLjQc6bOCSxZuFHfyOzSkYdaNx60WHwRE5dIEgDbLdc4sKa9bLk86AH2HXIvzzqY92e3Bgi+lM
G0IsDxool8osPsruUP1MbSIdaGPfubnEKDiahqsTiNp6GbGlSBngqePrpFmldoA16+/KCQNJaDjh
cSh7aWMx4+3WAKQrPqPH19Rklci5ZBiCMHS9v75R+PcO3qfQHFsn0Vpva4YXg7u4mE3NJ9ihndo8
KYBAEbnVAmIzHr4Qc6iEw3eIyKKBMpR6hOiXTPQQpArqkh7ZUMKKU+0s72cfUTFCbkY3GfMKii/i
vWHA1ke2s53DLZ0TD+lX5Tx6uQHqgAQg/VL2NqzTB7aYXiPMtB/Hvg6pTVBdVjK1zr5kZbyKtiLx
lTz6LoYYz2fZgEg6cuyCCW5hAAvFDlkJu45B7GdF0Qfkyo8+Y5u7Nn2r6QIYzeI2NIGTnN7m/gKK
Ri1OdmOPG3VIGUwDmlRuTZyHzZYWvYbbAS40uPfzWBIJWZSfvJTf1ybRP85ZC4FTj4SVFfZafk7f
GjUDRLovUp81NPvUaG3Xq4457tzzfpz9x7p4axS35dgp3XWR7Xwu9U3z8k3Ely7ZTEAWnVynZM44
7iEjSn0myjwRakK7bVdski/lhBDXkl2ERMpkJFtaYx08+bFAlXNsT9AAzwB9f61pVSO3zQ8ERZXR
PeUqEL8nQMDddr4OxfuGN/8e1O3IWwxucw0V6NcLzSMIoO2XJZGFxWB3FraRE3Gp3mQxmmue893R
UGa4Ij8HicffXgIxKexgywQNEy6uugy6pjYG17n3K8N6iytDMLt5n6EUmlzDZYZozskOBWQdXwh5
5+wSNXVX3uC0w2DPZSag6QZCIdmBmK1cyf7jnHAKJOle1yp5ZHiJtOKlQr4W5G8g4/Q5EDyHzlTY
28zno6uC3/xsmNP1HAoNSbDvF79lYCtNtdK2XzgCdQcwMOFoa4ycOKVrzl6xDQ4NwwrHjtM1VBqn
yC+5QqIHb4VLwAiRHijMxKm64iJ/oiQyrosrY8hS2hI0OTFfTTJ8O8IkLvzJm7LNITQLNdOsOkXf
zNodO75AN2Nm/waNTPV9h6hYQrOC0vXHuoDkAQxy6z5UNCQUfkSud+A9lQEOy3ikvDlftveBUbGF
SsK1hQV236y8a7PHaGVAyUj4vq1nb1UVJJdgj2rePsKNlkAUHu5gETRJakPjeN8vHaRIu7iIhfvS
Cgk4Yo4+tw2PMBB7LxOQZEogudLhbDnu9NYg6MOlu/I8Ql2tfmn7prUgLOSODyEKdz2zeUkTe9ej
kOCzdf98OjPRN7cUAUur3zld8j5ZbPDRExFBrOB8kZg6vGEbL7v7x4RAoHYi2fZiFvq32U/o4vvL
DsfBMQt8YKqRfcIn/wUQ2dyrGV0jO34FLRa1ZWzOlTvt7i2rWtAw0Y26Qq87n1kwcijIcPXhnkUa
Q06wK2Vj5Ce+OMqXnaK93TLu+5XEZWHKB3GmqTdBl2TkRyc6OGs9/G1kDPAw0xGEH449U9u40x4a
fN14cpp0OaLNt4gyNN3muVBzRzdjlK0Nqs+5lvmLDJ89vSUxUnNIZLHHqvd3Gv0OtG48NjrmxIfy
fvYM98PzbiM59djN7hhdtsA5VDt5NeTHLvel5NGcM2beKzOiKzDFODj/+MKzjJr6u3GCIgZ64z0D
+FgARtLji0VqCLPB/Yx/CxNh1I6jnxgraRWAijkc99Cyr078WpriO6W32+cjIyv7xze6DdPoSEg/
r9IieDTWB5l9adrUJ8dfLBJdYI6gR9dK6UoMIOgPfS3PdjZWUC2BmneEE+7d7oQhcaWJ/maO5mJe
hgJtM4zv0z+3MkXP3v3kKD2FR/HFFwRhf+uzkSLnnyvN08K4D1qYcvmI8Q8skT3qb34DJkG5iekj
Uf5rgNXgvJZ+Ft8mYR0Pqt6p+W++InJ4BZj+gW8C9Dsb4q5cD90ohxuOenqeym6t1jkkd/cfz+yc
6nUa69W3qnlgv/zTmJW5l+sf2GL6n3lNCwibeICcAeOxlJDwBQuSDr+41+vs4M+xzn0PEem+2XIP
Eaj8gGcKDZugUKYgMCl6t5v0EG4Gsfzwl86te/0BNb6CRV39rtG49Z2xPnUcvfiUy9alW+ea/Oxd
aKjk3OphoxzECNvYL42BMeI2eTbM7DNa1FIqxMA2i7uTxjD6RGyxh9ctKQ8Wpzi9smXE8r0FupeD
A/M+ufDE4pSrbi5QvJQLQwbmOZqq9UkpUoE8fdmu0g3+U0Sutlggy+DVUozEJsH/2l3CY5i8aMv3
vIWwTt7HXbf10XES/2gP3k0uNrkbFwJ54VFdIpxYSHfOxwzVcQNdCMl9R5vpx1hI9KXQBDME8CVT
jwokMpDM4rhyObRlAle5LRAje8sH7XpQY3cSk1NxU4xDtVzHyx3mEhLYpdv0ovSy6Q4IDPGdrZJ+
8Dp6C7loKyzDF3PXVDn4hqK9CUkpPTrzbvSapUGaqkyX/xHvmNa+BnFy1DHanhA64/5kPTnhCMXc
6REV89z2ZGdot4mg2zgYFs5PqhrslTR70t1zdAogODajWy0E+mkhhANosHtpIDbTq2hhtZh2/0J3
iM61Rmylo+BflXnv7sRQtJKdy84FcAStdh1LWEinATS3o4umkP+wtrREIxGk81m2t/O/hWpDqi9p
mxzqpFv8dFrcHOmRY6AImA5Nf+U9oulNYVmQl3s2dW5PB7oNTtDsh9sy59bD+YpnFoK3MiHZfXe3
Rezw5GHyN3PV+VfEDCFVQwNze7KBGT8IGGBUluLbBa2X6B8qq8CRasr1RnYV85n35pfthhpdg5lC
9IARDFnQYTA6R/Pux0bBQNabV/GlmLcmTEqpeSWvazLuapSXT5UO7aUub6xIU8kcnSOWn0wJUbKu
pf3KwNb4386k5CtnmJlpJG5f9xix8UJVc3MvPQh6YaGXggq7duSbz0nCIY5s1U4GFCORkD0A4h/I
bn8vhyHlNzWRNHiwNsHm/5CRjOLoFuUIYD0hpNTTxKYNL51QUUMTyGURupedDwI3YGaMELDtR0BK
hXUe7nDa3KbGK4jtOW9rjAdXAGER1iQPcIU89G8Etu2v3jFjfOVK1wJ37RC82QF5SAw+fY+ApbIz
Eqi5oBsMQjaa7VyZ0QS2RglX333P+HGy5BihJuqButW229BBE210KEADnSwmn23T+NqA30NIAsEf
wA7mrn9t8cI4r6VvYESGZMtvaUzlq0v7aJNlEsikZbqbUSY5Q25TLNNBP0y6p6KuAHgTWPT5G125
eYSTB//bGS8Pv/A21QRuK9g9lqH7ApEY8bQwqKfa44xW6EKViVouh6VRYk5pvjbn0o7bYBIERHD5
1z4xNWi3vNMisRjAwmoTj1XAULqvT+dk24WT/qqJaGj/HQYhYnTtTpNnVDKJN9fv7YhvuI23+fv4
gusYlHuu9OcJ+IV91vFhA2CZ1W7utBbmG5Xc/EkVo0a99q9zvpWRf42ShnvZ+BTjKfpBVQJuXWlp
l3gLKN5qp3cqcp3jltSStJVBrhP4WK5s9olm6EdjGvSn3Wy6UZIgPZzCOV5VYJkHgvy7b1ZtnXhG
UJ+4gHiDO2MWKIuRkiQbYbcdnLlqwnqXhyosNpK9BlMqtHvwHd75YZR5u63rr7MlNZ08XBemIPKE
gzpHVLF0HP1yUMK7ovQgtH9b9ZisYYQ7Cf1pFfI51oGATVCISiDj/aXJv9FOvO/rAtTfyYAgOELv
9hgdf5bsVwdu1m5KjQev0b+hgva5/fkMg6CRVqo+zI4EHIBt+VcWP1LJMxB9+ZmKlozO0RJEfrre
tQ5CECRxMcsgErzMcXC5+JnL7xYK3TBMXz5+XY32VBGfxVuRKjL4LgBG2a4cqKlGTbQm4Klgr0n8
llejN6ys4cPhxlrnVw/v0QYEhq2z/a1Xum/EaKen2GHfy4suW+7vv7zlq3Z3bvJy5JwyIQXYavDh
ChTQ7ho0bONgZzR7RBQfzBC/qgb0pkEA7Zh6xdwhR4scU9MWHE7oFBQM6cCRGMXuTXx4zg7WmFCW
EWiNyug/e8613xuuxlI5FVr19S0eciI14bRVr893h2LZKHBW8pmeL9FvkeCN4UkJbTCUk10z0Sn4
zZvRkRQoQWd/aJAa2IYQjeo1qwunjQvIvAQZt3446rMFar0lMUIrdPgdfn+FnGOJjmvgtljKuM8k
JbpZ0Mj9ytzhqARIiSED26ui7XAcfOziqSeqCV+CX4D1wnnVy/gWjNCgeBxBpQSNf1nSzHmVq+6g
/xf/TR3TUWlpHxM0WrArtBJ34eJh1x7bkOhxBiHWwVeMvXe0LKI7Dp7QcjP/z5/Q34PHlt4RmvL6
7hCol9vKhpJ3q3h21UhjJpRZvpXZO0QBJn9s+q78TAL7aJ68QYtb+oCqH3awucyo/bZJqJFFHXhl
pk6y+LDD01++y07QH8f89esZvMi/AyP+7cpgAXNGRheXW3r91Xh+dPclwWM90JeH6MIXzZuD4zop
5F8yzNvCzeg46UaSmQUgpGHej7mK+3xIUYkClF8jSOUbiPWn+7oEzSo/noWZpg9cGICADiwjJoKc
Dgg8BXbFyZyDbeP2XJ+d8Fz7rUgIyDhGZqyjHMJMzaqgUJMA7I+qkXSU9kZT28nTyunkt/oQ/EfC
D6hvLGl6wNHN2yEPMCOqfmn9ck6BZZDfl3Ksn21+aCmH9Fpvh1gv17omWquSJ9Uv1WbbqKOke/er
6pqoa6V9c9SE2iZY+iIbw5pQlErbYmqFF3pPhRe7yWA0QTHneSji+D3ZgAmzJYkxnVyMFrx3Idct
bzkXCJJSPGisd+OGLY8DZmj33pLDMf1qE9g+BTnrxOuNpKtQmmZI6gWl/RMyb9BZSjD51wUDOBjm
yrPP0UHivM+BbZW/nNBIO5ippXYGhh9IV+2zylz4ECz4T8fUyBrz8pDE+rB3ZmAaqm74u0cU77s9
dMM/U6d3Bq9KWEOo+80j0Jh1bWjItQ+DO/ByR8l5le2tqTEfPCRXX8ptk2wrpp8g9YQvB6JIYLxg
Xgia+K0p5lcGX+TyclgfwygZrDQxKtNfS9b4surQ/XaWf1SDNUBRqM2gmn17rlxvHAtXdLVdbIwn
E2OkSHJaLbEO9cnv9MPc441/ZDPKefinRW35WozzkeATEumsQ0kj+Kh3hFZ4KhHgN4h+fqBw+swK
VPrWi2VFix74I/7PJltWUap+cB9VxdBUHms7TM9dx2OE0e4onZrd+j3vEf92DCPwUM9gSTfsz0R2
c2PGD8PGXyl63OjNBl9RPpUO4bei27vs3gLfCUXecc/uBd0Cj1zC9tEexPp8STwd+F3mYIy6eQDM
cXX2Rz64MGyps+ejUR38ZTBy6JWG3WIgaKeRuA5sTsj+lUJ6Y/l0lmtekJ8X9j4wTDD9iX6D/OC5
Jq2OhU5Fc2Zz2M1gksPphZW0Ml4tha5bqfZ9MSnIB4x+vknyziRJ1lAaNrkMJwfPlJx+Sovbgzds
+FP/idR55cHFA9bsIG82hteRLs1BTvbLTe+jXWK6oiVkqu3vDfwoDUmPv6YgdpY8FUPptM+oDJ9h
4bWRF3PcVDThAMDWOd4qplD7HaUX4mG51JP/tx3vPCGdBPhXAHlFEr/ylt8ms42KJhPYCdw9FMMT
f+7pu7DwZ/41AscsX7AUN3ZZbr6Js9Z7R24i1j2PlDXN7Bqh4MHA21fdCooNICfpUiY5wtG7uNKj
ioI8dWAEchCBCutKdV11IT2zbzxltcFVKToxQijRyNdkzLsOTiOI/14m0StRd0XX3suQ2enll2Mu
LPs9oRMgOszMQV7o1PMnul3zXTxS/8Z5+wj7VRdy/Vr+uOlMlVf6V0kHjMGolA0iP45VWI7mJauN
ZUdu0gyCL0zouDQDIQrPGLdv6mPrB07mWw15eQRQOKV2d5tBwIsbyJbsGvi6E40qqKWsEUHQLBIJ
uYc5XOmKudltB0zByUt4zN9PW0QvvSygcD5MBb3OUcZoWaYkpzc3HlVmhNGmTEcP0LT+STaQsbbg
/PNx6pshgPczfsG/DBtzs4mMKUNEROqK4uyIYaFvdfrmpKP5R9sSnl+CPKGbNOWKUpgklCPnEwCS
KkUdWWwkx3mVF9JfMR9QgnIWFfMapxLCgjM2co5jGj3mwjLbpwP2yPbR/5yGsOed+18roEE97Z93
WhTsaCwyW6yM9vLX2L92Fv2OiD6FbxQemCu9yqvpS2DyqGaFMARGaqBHGHbGQDUyAPXP2eb8iv3g
hnKFuY2aaCscEZtXCmreJqURelwfcYDYL5aHA1dmIM2p6zJvqEEv1l3FskZCVFWmHTuGJf2sedes
WyO1D+TSzbCr1ZEG9ymxKt4NWXgotPseWw/xXdgCh3Ml9YgkMqF6yokRdAo5eoOm570Mr0StoqFn
dVUic0hqOQsXx8IxQOF1R13lwN8WpIaoDG80VevH+Y63cFmNvlhgYX/W1WwAvL2i8DzZuLCzTsU+
f8UW1/6q8c8SX4rCVY2UrxgVuf+acCbhYOVS92agF4jMxkaAleyM/Wzh3IXTMdd2cXwUJe9VaRIG
wn/6cQkDT/nL+7oCiVlisf3rcVtFpchvVi2LEnd4qHfwnzSS07M2RFXFBNDM1kLtbbdm0UYEfooW
944q65wzf6Aj7Of7+b3M6gNVRa0/RjThfDf/XLEfB1UBUppoG8a5NXt5Rh8jIxCvMI2lymtltZGI
9aPdoc4oqYpqQSH/dIQolAEYeVDnrAVZnPBLHx0V/NZoQuvvbUrPy3fdyXZEw6XTMeoCbf7pQflR
7q0M9g9xrWY/l+j6KBtmcUtPo6NEVDJ+g6Dc0aKke8480WmYw6qknt5hZHYUSfUS5f7g4ALmSGhE
oyUoI22VI1mUft2iHMWvcBx70G+hjT98GFCDTTdZ5SIXrFXgoYwCQ/aIXsgXICwRQS/Pf6y7j8f5
A2x6WUnEC19IlhS6X7qBmUPmOuF6BqOCiokN+YaCEnMoy7EWacxh/FimVoay1sEwiV0S52VlpWJF
Cs/kF04n/EhOJ8T3HxkEEyaqLNie9aLriHRaBhTwuJStR1WY9m1JKNLp1QxLNQkchHzYPEHUL0QZ
AnyAao+fH/gmV60CgmluuEn8Tf8OPAV0z1ulUA1OH+vvIcmy3ohQg783/aWqofnnaELZZ/33y2UE
06bGCigD1z73rO1uqCYk6jcjFsemgOIAaKHniNAM2eISm151lW9P3j4kkXrszbpDvfja6cT5f/fi
oX9jqGiQJu+eOU3dYl91EcWmz0uEIkkMjBViurqb6m0D0h3hXKN10SUx0w9YnQgLAc7hp44Xzw/J
TiIDeYzlJdRzkrR0uO/xQkD0DXd3X0/oP1meoGComt0eVXqWCY1qYehT6IxJD1B3XDt8LSf/5/79
z5JFhcui/QFI4uhknIVhuVIx2RLEQwIU1XpgyHHwau2nDHFDjWfvxhYkZOQgfmKozMSEnpmkjyb/
EC+UrTDbAT5/bquh7JcK3YXQ7uTwgYoe1e+1rFhpNPmjUgpdlBWMqxUlRvjFtHMoM7K93CPOfUAt
90VyARBtZzNYSv8fQIbQ2LruxSd4hmwHFP6QX7jjW1JaeOuExATOk7gkwJo3y7DdgOhX/Soj4mPN
K6vni/9flRPR8qBZA4VAx48vgYsUVGMWnEhRd6y5n7PpyWNiSb54yWYnm4ROqvu77lkhW5WILon3
E3LBHU2eHdIWhGK9Vo3iO/JUqxgoVeqaTy7kwp8f1ALRBokNeuj30Z73++6zXlBOKPu9SoDo9WhK
hvyq+HtNfVyU0kYwiXrIhNkIPGoUkJ05DdZKePxXdgp5Oh+HJHq/aaVvzoq2GbYpvq4p+scpnOp/
4611xeXBJVQrufX5x3U49STQWCWmAT2JvwNoJBo3eeVWK2C3STz95qkc6J/wm0iOQrf78/Jo1l1z
KT6S+KH21V0qd9BDZ8JHsaQqwEZAxGQ6PgNkmxjF9sSv4ZokIgjsvjWyRV5SLHYJ01IF99b5zowo
2wu1vQmPjX14Sw49CM1Inre4Brvc1Yov3kdkcNZkfGQKmlRucoGu/0hU8gombBWFV1pSiJACXJMB
mftgdd8/aZIBrHI7FxfNFCH93mzKAq9J/4hUN+y00vbgVWp+jmx4ZOe90rCjVNxySed7ObPZ6J3r
4bwBgskcoZXCVT7DkPttGBe5rVsF9AskTyKoIYcowCNcDGYsbLWsHzqRHbMeXo7Z32gtbFrInm3/
U/8SomusCkeWirnrvNLXWuGD89U+s/BRAIIhou0Wdm8zfeGx3Zb5kab8t5rZHbvH335kddsthBYs
KKvNGYDV1yJRd+2G5L/WWoVFWhKtPxSlbeq1NUPmjCj/Ocju/VwiTGMsj6JrXKRsYkMU85QUMPau
zpWCjZELJOb8ZTOYACSkIvNHVjBPlMh/sik5adZ5xOfnSWs9+pZOBXEgSvejBZu3SIxt5CDYd/rs
S9VUzjPI4v5QArDim/QKhO+ygeUzAuEIUD1PvHgudI6j6U63SZvhGC11Wbr2Ap5a2RgoBJWGieVn
FF5MWD3PcPnTVXx1T57G8tXl1dfLvWYbV/LtdFQOW0o56EkWGeiO8f64CBC0b0M1qeYy3uya9XYI
affeGrCC7MfJMqAvFNdHmcbLfKc6t7rhJjhkl7xIj+2x+ivZv+vbkL/ehlLtIdUV2Me3XI76hOoi
CbsxuPErLimszFSIsxb9ZOIOlBAAtu8oLrHFQeZIyRH6a3jq1Wm7F/zsB9k2TBm5f032H3xBRypQ
HG5BDyq6OdZlpOlyc1sESmzuJerf0uAOGWZjHx0027XnQ/3LPhHn79M5WohhCmtPwEdEMeON0xtw
/jcNTG6DrstBoZVoTiXU+meVCsSJLsILNIDdK6juAQTWiA7dBW8edeYa8Kxxc9/x6G2hLFqy420w
WexJUma233R2w1VjVS0Y4H4P83tYzCh/YU21HgN2eyOOAotHw9xzIlx9HO9jPsto/5/CodCt7yOT
qeAjBplnSBhcfVXvWDuyDIUeo7a4to80OaDop5k8F8kEI8ClmRZ1cxg1xfHhYVteppoweM4hpC0u
wupcrRF0PZydQWlaI51Eyv24KPhBhW7qHoH4rTzpcwdRB2j6zYTSv8YGCac9LDlrrze+f7JjqHfT
YHqPFQc9YA1/o5WwT4+rd1nvMq1jce/Vs5RL7Ae9CVLT2ADgKLaUemMtCa1EtF1z27V7gKVcMLQE
iqeKILUfURc8astggiVJ0FBM7tTWnsFm6QDs59FEgBVYcpm6oUScL6pJGRqQiHsKp6LU9wegb7LF
X4fAepi3tvOl90lk4N22B2U3heLp4FdS8GT6YCqc9whVZSYKFm7ngnTbaNFcJW1K7YO6qYm2B/TS
w+V0k7eImAChGi0pp44uTNa+9jC8WziCL79qB2zUTmLvxtLI64f6AzRyJ9+oaXAZLca0SqxebbaO
/41WFwlsO8cr6jQ+qhVsxESSqyTObyxDbBqpzANzIrAnW1XLkwT8wr8FbNjFlRsAJCMuTZI8JVXx
JZ0LhLsbDKqMH2jcV0S+UiKpDBByD0w3uOTqqz+kvZQZIdcb/8X8ChbV98F40NYJRHHKAP+ysmO4
4OTHveIeeB+P/052ua4lCUbYUO+4dFChhXcxenWD8XWgE+hkZN66DjHud7KmikUpyYdw+rnwt/Fd
Y3OumQnrv6MglsP/FMX0xf8fOim2hVAOs3xJ1nqn1FA0Uxx4Md1r9aLFxKPkeuVN+oSZ3txukRjO
JwnYXPXnSwbJ8eYgx7afgUjXfC/Fxws3zpNUcNQ/rpol1AD8HQp+GYW1Z5BUBTCGEuuxogzpoL6N
2kw5AnvHtyxX+qNVNWMxC2AzqcHdb9KMxg0WgumxS5v8W9b74AP1FUX0Y4yxaL2WbNSY2CjECpMo
U67eAYqhnUy36m1EwhhhWoFIcQE61EaxR+UDTllubXTr0wtvvQSCKEH92fyFPsKjyeFToXrYeG5B
NLikjRKI5EzR5uNqxWxILqKAfbH/A8RHeWn8XHCBylnaUSDlanf2iiWo0MsdugGTciQFNFKGjM+x
PX3Ao71lmgFDwEFPrOcqCqQ19erHf3j1YNDVGfPf5zU9bm0z0wiS+Yl7AGBdEZQ07j5aHTfDpZBJ
IkAwmBRbhmGE3/nKAQC7mFnkUmtJJc/P3iT7XOer4n43HtQEjNQt9H03xVG5uo6Y245KfSc8jVlC
E2bPVBMiW0+qnDhKRf8dn/hdXaHRVTk4XIOUy5vxw45fXnGHwM9dGTG97kplPhiQF2ZmSAo3K+8X
IQEIxk6Ea/0wx80skaW0lIzpBkgXG7ru85PjIWuvV3txtG0NFneXFAFNpT5rbEmYLvZ6s717t9lm
07Q8JP42WlNeTZthpPE1hCdRwPTmGbEpoM9cZueHj21IvwAV5pUpkmfa36cpSfZLDf8LLmPEGgxE
cEJTLqfziBCmyHJT/tbHByf6/CSxFxRH0Wt1Jyhwsso38ttXNSVNGtTnIeXNlgMpGGZJ0gdKPzTH
zcGM+C77OMwWrdU08ARbdUluVxGvGOrsj78/CdAZ1RmEVUnfOYjY/J/sahrYneC2P2ttXNZqtTeN
cGpauAviVxNs+cXIqwrRxod1hbZ6cXEFXT64Nf8B+RSRc4eavD41Y10VX92d4Rl7kxXNgieAnzwb
gVGXHTIdWPLb/aHBuXM7fooBUHgvGjsNXX+YcGXGpaekcE59ahcF3TdfiQgqhmbfpvZ1tlIi2fVL
cHU1EZPrhx/0uHO/xyyJAnIDoByc7fwJJX21I63gliFZrRPcPUA8yLv8d9tnpvERRv0zwY08hPyM
bMsJ/knzTJ+EA5mnaktmO+tj8ErPBAyosU86xMd21E+PSxqAn0Ho360edcw8FcEfVaMbJic8Ug2D
qZvP/MEN8Pa3z5Vxt+AE4F9AP2WpDEalaonv7amRD9A3cnsONGhSHasF77+UGCbJwl9kLTAI6CfC
uG0Id6Uk4f4jyBq1JtcNYjn4vhdNqHGwnPBFLUVGc17kAAlceDtT5HaWgoX5z8ovg9oIj7NF7Oz6
ojhI+mWqVsCckb1Ap+Xj3HKPIdSusVibRHUb/Zpg8bj//+dPGdQXqf9j0OD5mk6a978rfTJMC9Z7
rSBKBPqPsepWu8orI5KTWFKjluc3o+xAvlklatIMKI1pfL92i6phzT2Vgq9MC4qFCXe7k7X21JKP
vP027XnZjymIttMGNxjZ3FI3ZhRwLCYlrFFbdYjhO144JbNgIR2QInP5VhJQI2y7LQmgCwzygn3P
uQ+eMDuY3EoKdn1i+9PJsTrDXXK96kThmakUPaqppYs3OmLskSogqmYZFuzCe3iRWQGD3+rVdedD
P52gWg9x+miWh5JJ/nmC6wrthtrPIbSF55HJP+2FacM1Ah63CggK7vdJcD/87fH4I75DaTUAL93f
q2tpiNXD+UNWuH7YqdTnI679Bt/SwyMAUKqQwIMyhrdYoMpg4Wz+iLtcy/JWYosGnx3gh6YicV2H
8H0Syfi/XSqP68+BmKstuT5nvWEcJIc3abGc9yn/QN9qai2viuE5EEKUezHoidPd/10sNWzoFBXK
LS7wKDJ9k5oRCYoTtQMIkzk7qDtWchVOiEga1qj7wxmM6ljlO/t1pRYs9tIbqu8EWCaFaM4+Z0Un
MoXeLolPnooBklrlpqZ0+hZCCE6yt7baR2JgRrdV6RqZoLbcQKD27hZl2euhkarlcqIh3ijKxRSi
mvDMLNY9cBJMa6UHrn+6zpbRBPtmDs+0T8zp3/7FbSk2ftjyQaFvgtHQxMnoxctGW7w5JOMwAfpO
A9O06MNt0pXTl273xQp271D+vsNuKy2UyyWRgXWzQNzq6nIf1DC94AtkCAHVS5jfHd5vTVTsQA==
`protect end_protected

