

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UXXDHK9d3YtwspCksVg3cn1OQkWFk3QQ1bnN8kcpv130B5dMgVD8+qx+9EwjTR0JFb8FYrcL/7dg
lIwdmlKGHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lGlirTrah5ntgtsTqcFN8kWYeCxRHbehSLZqyiEvescJE+ORKShYIOu42/ExCc8hSawNVl9qCirT
UlThiM+Fc1evKMQYzaFIzbKiio/Xw8rjRfhTJKjaxdK3T87LnrHcsuSrci+tl+anpBCM3X47tPxD
oNmgZzATBY/NVtZsbvA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UAOAU0ylQuQrszr15mLZsCg4shnqFlxQBAKcqwUoJfM+lTESkAcOosPqKsRH4IbbLlaKiP2HCFU1
aKEFZccPWIgd9WlvneNU3oFbpPCOyV9eZTCX4e5jNTf/7OwRRATKc0mjpd4lxBL9xFrSwNaUKgs1
3vjH77tdesEDAIn5GZ1C/7l3wjwnB4tAiaRNqLY90lB834tlc4mPcP6x8L3rhv5EXfqU4jyJC8B1
4zsO/vH5+VVa1595cRZ3xWXEGVMvmWhY+6TDUJCMhztjp+p4kbQ87UqJz9ddvZWB4hRfjo99Os6I
PqyD9P7zikHIa7jafFMtZu0Vj7u4HDelVYnPyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qRFhWXCy25iIpt8SG9Mt+xW3HRp/MFye1jJpn72azeuP+g/A4uHCFxvcKVhzcuE8lYDqFZ9IBM4P
ZjcyPOhURivBaWk0KosUyfzbkORd8yS5XcayTSj5/d+90PPk5PXVCLjTrcMbg0+NO3tiyKtPpLQJ
f+Ih38e2az80fHBgiqo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tjh0p4bhQQ++Enuq/zxHJnIk+bY5nNzFWlWKnTVXUtnLIlVGko6ShpeQRaCrGzeMC58aHThmj0Rv
eUmPmT2uqc307TRbbuUeFDYMANj1kcC6Ygs+bdXnSkWnOQFu5reSEq5SE7OMIvzdCIaR/FDvSj26
cuj56WGV7WVTg7EZvTcQQsjBPGe7MBQPj6gVbjkHGUTFOQ09cS9h1BaC9UWWfJNQjyJE48PH9w0J
tqmbE8H5AkyiSVZzE1dyYA/E3WjYX0ib/4FRIxCW96Qs02ypuSbfnvJpIyeRwyQL7ko2qezd2p0h
VgIw3omrmALcnzzjpdcOgkkF7sgouCeIApSqBQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51440)
`protect data_block
WnPLmnLA1JoIk1YF2/Eu3H+RnGtwuI8sJDdqNcAhhHJ+rSwQPPRx8+v1OEzeU9FnwQTUFqQNJRIz
/gMSlCzssC7kSJNuwgMZ178xDUFnqkk5anrtR96AiUCn/Nk35XhQXL1u+OBMwfhLR4yxLKgxFbdn
c8ooZYVNSEtteIB94ne42eApWodFZSqrpJFK/BFnUlsiDx+X2+QLBKooLvWt0EDfpP9TWsqvdcfP
KecUrpjs4ptOOud5YdcPlUDgCWG2uqgHGTQqaY8zcEy1/VW84+eHTyQ9qQu5B9HFS1FAMHzhLsC/
F76DVA/GhRCViqA4IgTqCs3e+9ZxTzkDfbDLplQdPtUv2ty8KznMZ6YlDPCiNO1lK16Rj8ktAdq3
UCn/9XGk0iI18XDqPHzCJxcGj/xqWBCSh71gZqJ0LCoz6vftcml2wXhjOAUQJwZgYrj4YtiPNgN+
vCRHZTT4c9/xUXjuzScgd//tkZPiQDjTi4HMmJS/rORLDCwCLEE8awEr4E42v7bgO8chtvlAXMgg
7dhJQfinkAD6CCoAHr4ZLsdtp4q/9hc4NtgPv0WNhUjIhvhJCQa7+ReGOaK5LruM7aHHTVkwXl+t
doKXE6CjviVYQM459+MKJuSPRS85rTjYTCed1BQZ4CAsfzh5Rsy/54p9cmkW0bZNfJo5QiJcIcwq
jFShrmGpCemrW+NUK3iyg2Pnd8RcNLrQeKMDzLFng5q1JLsjuFoZkJ3/mIqmYhhHdQQyXMmFADw4
oW4L8uAIxr3NFfRYqBFnhb/pqlfpdsqdDEVUhwtxixX0J/MLAlcsXmh1E9zb5E5Zunn7ie+aQiXf
lBEyBWBfihB7XSMTseZ6OGxkn4MOrTk5oA7IuUwg49SV7ad/AmZFFoZnWP0krTqzWkF//W9sqXPH
D3Cxt65U8Clk1XCGgtdEC1dBr28OdA8apRFs4mOHp88XD/mxh/nWDlLRjF7aG+wuWo5qVOEUOQjW
ejxXTMfdN2WJTqdA4fsVZoUGEELWwSLm8T9KacMdZPS4p+XYOkcTngYFqH7+u9inwR3TGUs3ceJb
zlT/dzLDajxbyQJSmeHC0dsAlwcrJVBKkwhfn1wtu4hWyLAjsP8ScOwJ1rNEggyN7yCSvUdnfCLb
vqZE/sqx10xH65ENr5LvXQXgytc+OQk5QxRVXf/ImtV9kemzm6QomBYasqblKxg+cH1ClPMatqUm
CABXnL0cLjCiReOa/CsA8o1bxifsYCIWbBthuNJNPURCY0KdA2MB6asjpenuGbk/bT+voxSt6TLO
JUe1j5YxAQFrgI2gyUeH9nhYIQ9gF/wYVwLVdUxAbt17GJPBXxQxs8ZH+AuB8q9ViL8P/R1KZC01
572Wf+VWs9+jXlbqG8Fn9TOpHxr0lwY+9+dV0fB7Ll2UCPzNZ0kkv36A46eKBmvz/hqNCwN1zIc0
C65iF5DK4ELERpk7a7lmGOZUVhevrPEPNrykQ8TrNaCII66K28Aci8AJnr557uXW/9908S4Dtzrk
eFwm8oTvouoJDAxeZ3TWfo13PtQn15Sw7Ir11/xrMFPpuZ/rU9+Anc/x85FeM16z6wz7X+G4fsue
IZun+g07LZAKRpygOrc14Jqk2cYwAKWfZ/JC7JaPaVe5gaTPSCdwJ6Dya4p0IyPWCdRZrO13uYn2
gQiaSquSCMoeZG+WL+t0UeAoc/FEGLyC/3J8zvDM9rSN+KCBeYoiD3B8mWVNFTcXe/R9xyq7KoS4
XxVoWTC5W1cQsZQUkjRFz3JsX1alGXbcb0enJ8e7vmMYeZSrnsybKiQYI5QGGLp4V8Lg99x0Hufi
b0m6R8P3JhofiheL0BrdQdMDqHsy6u9n2KSTJ7C0Lwoo9KoTO/lJ+tXUugiCsKEazM4Y5FP9VZC+
QffTMPdCfYrjUoVyyGLOaIqluPkjpQy7rVpWDK3SGXEhT0EGKdSxYGwZucMXNhVteWPzXBCG3AtA
2IxFIyoZklRPFYei0mg0ia530GNR8mQr+eDx8w2xOPaxtHiTUqnaucqKi24i6nbz5VTGgh//vWJ3
iLS84kuPa5izYRbs2a4KRCZ4CBsty0S8PXaAMuGMpHqFThv994QsC242p/JrLxAXaxUHGd5/EzH6
JEA0JA8QKYfxveV7KtbV57fqGiSfkPdzZ3BG7zKB5Dhf2wQ0nif2FdP1p6TS7jzrpfAXlYIE8V5U
oVFyCiRv5NAkQMzXUoqPLHuX1mcPsgnKf0XXAyePPyv52hN3Zv6oe6bRBHehLTjuHg4cwb6+TO5U
Gavc1jtA81/w49XEQcxat3FVMbDAYltrWsZFT9zFC4Bf8cpF3LZdj3aODMU+cmWgyQQJKSeaBywd
d7RIfIcvhPWj/kT0vwlgDbPpEO6itR7cMB0WVMb+3vtmTsrDZc4FUrScDHbSy0qgtj/dfJtFW7Rp
GxrPo4CGI21YkZaX1kymwNVlTOOuOwhSPC/9K7yg68vBUzY4hZi7ElHboNO6Gc/KIRxAnyP8QBqT
I1TI8jNyxPZDpHhyj3aL3nBn68xeBkusnWwrMuTzVDfQDJXKdOKdeByv/EjGnNXLGPKhy0nD0BgR
w0flco6Rb/8BnZmRCeGNoVx6DdSFjPobCdqD4ql+Ea1bLXroXJMbBvwM4S/JK+SoJK02otqL8lWf
EsvpMwCKFKRNYEuBIgwee0sQFJQVy7S+yO9r9V3wQNbruxirB5ZTvejY7htUy6IwrbalxbpYsXJn
6z1MyqYSBQIcYFOMQ7cY+ZOtBR+3jK8T/YSsqliWjYlX6JRLoJJz+hlTlAOUeZhxGm6J6gP106WD
pd7ZjZYzQzjNMPlztpj6KYsDysSv7LFwfk0pRrQgZ5HmAaQiW3dMnx6AS2k41YKfXyFRNmpN5mqv
HZ6b2hPMGbVzEtmwXp0yLgQjVTtbaxuGiHWRvErrLuG5P+3H4MwPKcUUsatZV7YrUM0iMYJoV1YQ
lh8V/nIoq6yzXz6NOZ6heiHapsbOMsp7cvkLf1kryqWh5eDTL1z3bjatWG/PfZiaRhZek6fBK19u
w5xd5G8/TdTOtGG6k2oebmBk2wQJRdao4JXDJW0nROzJ9Gsi0vnIlxe7TGxvDsTZCa+l2JG/p8b9
5+rrOiP/9k6szsF81VQEwgTVRfYljsv8EFCajvfuFXawllOPxInCiOMWJEgOIh/k6HjGKZwksBL/
6FiwBTDgJHDmW/TaqL9/j789elNYOGdONkZvyXbiQMRqfFL6oFkpviUreLeuGz6/u9U2/lt3Qe9m
iyUVIzneIQd1n62r0Jp53tQ/lLncRCRFX5hu/IqNipKy2LQRX2wMJmy8AqjFwRhrxUuJ6WgDMyIk
PRjb2Thl3KM5E6trX7XL5qHj/MDfIrgADf6EXf3c1+BCmi5BV8qxxFpWHxQAcUdT/tkoMRbkZGyL
8mR4AFbKCNfuipcOSQ4wdLXZzVnHFOQkqwS8RZ5KyTSXZOXIEuttKiJPOmZE9IeRpJ9A/7yxjoOe
37V9qm0MoHG4BR8T3NKjgpFAdF8zI0Pg9MNqQ3BJXzg+weVuNAgoVS5GNpHS1HGWxcHSrqBlug5t
SB1lbsS+3Z9m8L6uwpywtv1gDpi3ZRprfsyOXkxOw6YMPb6v4qF8Xt5leYGMY5EjxW0IL2+5X3rt
u4dgRnHdm3dCGisGKkJ1MZ4s+JID5PmkIBcb5CmBtfj92GTDQItS2ccEgSsv7Z14dr6Va/mRmkUp
aiUcwAdZ+lYGwlUaK+/yJf0Z2W67BUjMT+l6KmI669c3qCMLY5+1o5FlyzLLr16ZgiHUi4ev6D4y
vvuzvQSJqTb3LkzfqsELrKh65cvUf9pgME59tIWhBg8Shy7HmT7qbTbKMddRncUoXJjq6w+tNPrm
wLfLGOnlTLBPj61UCdgPUHdGLy8jnoRO8XRO/VLEXlIwc5cJo0G/TZACCnh/PHLWQZlluNN6OgQP
vkvX6+wjhCmF+4yB7ZHrBc3we69krhagNy77+bQuow9U42v/5ogTyxANKnAo6FFWRsmwN6gVMNAF
dyjf+fR8ZGytFA/UVrHDNHJpAqGft7bcOC1IYp4iLMrVT3NYbwAC0UwpAh9T5TCWplFtVp94sqVx
eSQ/Xv5ojN2dADh8CNqHpVkHlw2kIHmRjhaUbkC3zU3Ld/IGt7pb7GquqMoGd6K6X9KlAGYUWMEd
3K8K9tFEtH2/rWmpn2IAIYsSVF1b7RjqMyzLgwbYaSL9fiB6HwmGFvwXlwNBUdtAjC6gO+rocxi9
31aMptfQMeBXUY2qSR3MMSslT3LNxpLy6QpizIq8MBHIVc1Lvhpjwqw0VubFZpkvonCrk4ligi9y
BaUo7To0boOnxBFzTBi/hYUcAbIJ4rLLwv22MSF+MV4AYktM0iHSslkV+NzDc/O9pfZjkCCyRWWl
UehNmOGa/4eOdBTf3OFGa+DQ0gs5/IXch5VGO7Na/CojzqLm9kG5aZIJ2dkUKDiR+cHt3HUMsATW
RhVAW848zaqr8ZF/WzmqirnekWN+uWLxBnYkBilKKeJb9z3Ey/0SRgDHbVDVBlp5X7JTQdg4ZmTp
BFHHSqQU1he7vxKokL9rY4e2cr9BFaovSC1SIw0O/YxHfmMIRWnNyTiuwgBe1ZXJktROgJsfgE2w
cce+hs8vj9GE36mcVFNPxng3OsP+edk0BwHVgwqmprQ++jcoqjJLy+KLoU9nte5t+DS+9sMuQfIn
2smcCSqyEjR5YfuD2skh9xPBZDEPFXbCNLZ5OiC/L17D4ir0IK2mvYFoaCbgeZho8Cb3TNWrzl/L
3PYs8FLSSz1GZyXUo04uy4MUy+OIQ8+Lt+1yDhSeLyh6c8we9Rj1Gcus8gTzCP30v2j9ca2bpyUa
jiyaa30hud7dIRlIxxJPRklx7CCCqLJX0vbUDCyfosVLklq1Ik86tcWn0mqB1lc+ZU6u1NDnnudA
9KZV073l6v9d62WzaXNXhCdNbG1VGuvgPx+r8V8j6gQP7+XBrEOY3a1G78BK36fjtTfcRQ0fAeLo
/FZmjMPo0qYX9weF9P47UAPxQ0gZbMsOGxhCMCjBg9MjZk+Zo0xjYRKXByIpbJIrEX8G3Htpf7DU
g3V1JSGwX624LSbc+u1w4eBl/oGuORZ4MvIoiJsNmDVpzFVV8GlA5s+kUuB+6/HVTC1QGAGaQas1
y26Tjn+D1nrQeWxHdbry24nLc8v/kWNP1WWzXohnCHavpciQYhgM5TtHGdfYMzlabUS2CrwYMxbb
mMjvhWDXUg4+UEkNg/IWLVRJ1y+4CCIX5eFIESzFwkYJEwpRLlGcqrPByHdxVXSMFP5eNz+9ylp1
TcjcNsrxTKrQAOlW6TffzJerbOeLz1IwylDUK5SppWcSjF4qcpiwWETw3C9IBCdHEH2fZ5mZkerR
7UoBdvHgz6EURF/NW+peIV2/x3wOFqHxL1SSa3zr5ihgtRBIS4/rPHuJ10wyyFxdSHA2kLr8/WqB
U2IMHjgbSYDOP7v+T5b0HPtVwO7Zs7C1kNbUek2p3h/tW+cnrBjrc2On9dKBKQLeq+ySP8kIg7x+
P2oRG7llRL3G/wHSYEI2Co7OqFiik19iIpb4mcWTg6EMgEcXC7hcZcBzZwAK36WmO4xmg/KG5JjH
GqIdspYYyy3GgTyHXkT0QLxxfjcqu6HuWRSqMMW8WHwn7VBYXAhixP6MKryqAcI7F3ixUv6n84j1
fNA4mgZg+yiVi0rpm7AqtK3ru4YQSh/F8bH8N+98v2tLQ4h08lJM/K92UBQQq/ZQiHgWgTbc5JX4
iYTL8dqJCBWYFPaWI9pIlhg97I9fUMJkfJY7i6bnwBiVygEGH6pF/urlmF53DwX1W/AX3ert9w4C
xy31yb0mNV2nt+DpOVmWCR9v1hZSaVwmTuZawXhuqP+Hm4VXtSxCAFCGSuX+9OL6rn5s5DffANOD
J23Ax+0WqBp41720hT9Pz8Amg4hRnXd+MyOkfiVThbPQAf10fMaOopLz96tbLyZAB/Zs0WQYGdBN
AaPyRHd3JEgm4yzhgcsEsrcKD7drrJLFJtDNjnU3I2l8JWn09Im8EF0c+H7mP7fqRb2897l24LNp
xcNN3TLAv5q/bI7KeNrukNetpUJ4FPNWPYxlyICQc293bHC8wKJ34VQDO/pc65bWX/d4PO8rAA79
YtsrWkwCHF2X7YlfOfiqiAbKDeCN1cIeOWyOzo+Uvq6HbQ0Uf7noGuW2kkV4h/wNOGQIgDr3cHl8
lxqwvucOIWzuWqkdbBF7AnzJBvToSGk1ajWSixkvf0uJItsIFikIoMGhMqbOVee/S4TkL93W4vRu
FHsomEE+rsiBso+sLO0VcOjGP3Q2a3Z2BuW+E55UKGzAdDK5T00Jt3CQPnbNIxRPiNY9EJdgClZf
avSpjr04LV8iiPKNcqB5psfUeV5sum2BJjYuTNfrAmRNwU6a5QF3AFd/2b55IWm4BJ7RI85AkpJZ
n4sPkTuMYWGtHCcNJFx1YNVIxle2cxVbBnyWE0Ym6TJWPbcwn3Exy+x3OrIbMTeWXhUXNQaCkjWH
FjKK5X7BpF7Hkd435AcTgDEI5bHqQmfn/5jbvN4EgAIb21gpi772MDbvgFWgSyt8rqCFcgyIUKex
Hd0CHT+6G/3NiNkaP5HUbubUzwXIEV1XKlP63LtljFEiE0u2RtqKvwo8fQPNTtbKgiMf2AxBWuGZ
4JxBiD1T9dFZxjVxnkBCLgF/omYdz5kCe0LAGYpHo3ytTMpHnnVbzlX4caoE+w0unJsC7z/G1ZY0
PDpQBksi0bYG6gIwRn9snY3aKLnyxS2B5+b2DIFgCAVpUH7AKCpftpy0dxDesJqJrestXQk+adsS
jK3XThkbm/wyyhSMhM03ayaPsio1DQqusMsSwc9hsA6zDb6U2NJy3rvSxwpNM+BY5QvsjytUuLGi
PpAi0epGCa25KEDJ29fZiQNrmfYAH0Fbr4CsA6H49EAbDlz8z/2j6fr2fAOazfrwXyg8hXwDEVs7
rmtmlwkVDAl1zt8QlJKQa8dfGBeG7jA6vYXMj1fB8O6DQ+S/bvcTQva4SN3Fr4wf/WRx8VxyDxEf
v/DkGphHQiWw4OFi5X4a1FB5yeY2j+Jqhcy3hqlanriDnaGOh3LUCuLZ4ibwyoW7oTWwzo4O3rMU
LqNm+gBdNPlReVBdPPNqpZmnCHfcanIBDJXXewlAzvyUv68bPqaIQh9g6lzeAtolQoBhTg/Geprx
rKd7OPwADcU93MWnBparF406byI0RfrRKROPswRq3QXByRGK1q4+DBMmWhhrSU0O07izlyPDL6Yv
jOAHteyIkgN+tFaG86Os8DkhkPrr0Td0cnPrIse1A8Jf0AItZ9+MWfzwvQoN55vC+qwJgveKqtdA
jJ70EzbLxuZcCNnSMeBzbPX2J2YEvQhDVWjIXWow6q72n0EA9Eg8sSOxA7qz68tIQyBz0M83lToE
hUGgDGqcIcTXZJ5Ag3/zsJtX0YVjZHSO93THq2ImH9HuQwMfOOuwPGtisB/U6+U55LDxBRkZIziG
v9E1a6bIL1fIda/qupHrkDouaBf+9ttwWZ42RdIPprl/EhMuc3Kf4FczFsKnns0vNczAIm5kGYL8
nV/V2PjyJKIwOkgR5dnj1GJd3IfwfqEZFemV5fM/4/tkSGOxhQNtFfl4usHn6lWBYBnJluTbMHys
uhvyQkjQiI4jDSd9su5nJEJdsyZsi1+HqC4ybCn2L01HoEPz5f31ADoEQ0t89orvNSuoZ949QWD5
A2FkvV7Mal7ufCj2q/fwcBKnUN3twgygrerrTIwqi7xOIvZbAUkyRTiDI/pLu4/FS4Tl35/AfqTH
oj+uimbBPptEJ8ssD+2cqKNSETKgxlwEf2doc7ARJpRq1gtYR+bE1eRgNLnHS+PSm9YJrxRNWRDT
XLRWxySJFx3yMEs3H++6ssYFPgmotz/93Za1pgp+Uqw6azP9jiigz3/AvnSNaIe92e2c2T+2FLQt
3GSSaK892PF1Anat/dojGv2+s6ZNx67X/XoqYHWu4eQqRJKce1xe3o4DnK60vW92btdgFQle+bke
O/fx5IRFp8IWX2cagDgR7+DmrVz68MlrG+v3eeGtc75tMqySCZiR8JXzsEvfsqbGXFiaYALgiMwp
S/ioDlhU6NWu7CmP4+TE1B1bxcX348DFcf10ruh2xpjiDVLSzvZJRYDI3kwRnkzaiu/XfWrmxbOO
9N0PcibzMn0W1MTzGghcK1C/MHIhDb8x25Yy/NUE01M2dV1puK/1rroJTuOIKqPBGSrWbl16+iz7
bxNPSnC/0LpowuQs94oxbBio8+LssLPP56Ueqry6QwY7MT6hcKPAGd2/LGfdbYmZugr2crWcZLUi
yrHwXVmyaIGh3dbFY4vQUa7JAG8L7dNo2IG2kIRczk+2GUINl1ICm4VSp22awG9x3eTv1TiBi4bp
9i70mKjBrt0xCAwECe1i2t0+fEM+HaXIJk9a+KDJROC9QOHljs9+dNUTozi/U3x0u+gH1NAMKplj
F/FzSBY+JJTNLZACEWp9TuqV7lLwJhagW0diY11c/M4hiHTwSuUVkpAEOkBlbqwTAtDjjhjaS0jR
jPUEmHeyQiZp2+bZPFRkpzn+oWeUcrGzJRtX3GuTjzNo63qg8fsBob2AlyAtzwL2DR7UF1Yodmbb
PjfKeOD/KQrSQzzkEu9JsDFkGcF2fFPyO2Lv85Ox1rqj9QiTRuS6/woR7FIvVOc0u/tcyzeaZqYu
0s4LFzacQqjhJBaEO/beF6rTOjFiVjbGUvMHsQCKw/wI0GXXxw3Ecs7OczBSvkq7ECMmmGl43lqV
6Iylmx1nBfM/qHSN+Cg9eXr3vlBP5GgGx3czE5jgbIwn32zhOI5+hQymtZj/3p0a0z/IQCJ3ob1z
nXaVzOe9E8urzxDl0In41dvth+Wun0Wlpurq/51EeIOHwdS7VIUI92jObSsCjDleoTgflG2dCFsp
5avdLA7neSjuRxFATkgF6aUIXvaeg8ki3/6OZhpS6LEFxgpz92LMmHZMwX5u4sXtR+8PhU4sU3AD
/oiQlDvPp1qbRV4xginXfXRGJW+uQFudrWFRsOM4lUaZJgubbl2+Ejp24ZnohF/H6C2OHQvfPsxy
Idab1Z6MdMCVuKOv9+OoBjpSPS5wcMiWd6MZo5k9mfRMUrm0C+EYJUdDNM2sUDTYM/LlhRyUwfJL
dtFjLZoA1ouomMF01iOKB8orZPE+/OI/0BAnOSKQI/cHNX7MFZVJIjkRra194ogW6VW3j+Nu6jXN
6l9KPoMBRHQALanosHBcu4Z88TO42hujFMrNkyot0plOgF0RIWMKMB8nxGu2FXIzCHEhANal7mH6
rMNYcemDwpn1sZx/nFWqObagDun3dpqVlPl7Or/tP5Vl+qzzkCdbGi8Td+4x8NAYXgnspwD/99uf
z5I1Plh/NJ+F0iE5D9ZuKGk34wfW0Ygic0BT/aavH+HIaofBAMHy9gWgvoqFLoPivQSeAm/NZ2TW
6wX90yZGd0mXtmeVJ1HfVo37AGxClk6rY5c27AI5hkh8aTWu3tabczTjtWq/mRFBZ9yDgC8p3Poa
UiHJ7swZe74AWjdoxrbxF6XvxNfMf3BTiigtC0EtR64OOPEWB9iOPGtxB+4k0s3GyD+mPaQVcxGD
6Z4GpPtcI8I3BBlOnfEbH/Zh979n5ylCtiz7gUjv9qfl0Ufn8yn6mPLHnuQEsHZPcp00cUcFwkAd
Qo7uLJte9QjWD6pBRWgUKro/uxKBEBkDQFH7TnutiGwLLRf8lMD3rmMogB1bfacXFQxgeiiMyr1k
DLy1c6PSzDWxAM5da475pu+a6WOyAgCIXY8CUYnny+Y8LSPraCxg4EPRTf8jt6vOWQb6Cd23pd+p
A0gguM3WKsAefjfSGn8CO2vPp0RXEZPRRAm5OEuyA9+T5orfqCJNg+DWUyDjy7szszL+BS1Zle3n
Oj5QucL5w1Oio3FbCDgAwfEaJXm1PVODUI3d66ADaIGIa0O+QEG9RoHYGtd5iuIE0d9B0Q8+5IXw
INd4jttXT/L29RECFY4alUULhf+wTZDG8RhH5mWaTNfiC0/CE06dT9sQO5UsRUOUuvg/81FQEAmS
tymWaLt26IQf9Md89Vocv42QT7FRaGQQi4MA0YMvt+Lm/v9n3HtKHf1sk7RzfGd5U3pJnMx5OUNv
JTVYt68oNjtDYCSZrLauVW3/K5cUORJWc334aGjZfC4EgykQ1H4Kq2jcwUdNt1BHxSsHnd7066Uh
nWQ+fI0YWGS+COdVO02mnNhQ9cfgX28wpHjFq3wRRfr9YiJrfbIMyqjHbWqTEkviphJbnWvOeI1G
F26TMyYN4ExlyZK3ksASfG9scQQV+QBUNvXLQcJgwsNNfBkp+bNK6Q1RcN64n6fRIeUTPRuTLTTq
Eg0yc5e7Mx13R4OzJu6IMwzod2Q5RqhG9p2GHTbsKqvIhnQWMpxVKuGPkylWa6czDOpSNLRtBBKq
y49pSTE1R5OCepvCzxb2vA91EXQSfhBinHDVnT46z8eCNIHz8ptziiG+3rnP7Ych6eYTNpqLsPrG
/jC1CUfvEh3kbs9uJoL0wvIPa3Q1yruL6PbkuT5pr0E7qeUY1VA1K4fJiltHPnEjkFZBbUeBECsh
ao9ktIibI+jlavgKJt4Aypx6MS+kBYCxp5+MWdEUeROu+lUJIsoUAorsiQcEVw62rMkygQbHYxwM
Y7krM3D1bKUDqZwefLEN/4asEd7m+Ya2vW/gozKl4/KEColDRyJJAjZJoW5XGfynsgRKoc58bo/T
9lekAq7IKnjOPFNPyvxmXnL6jlH1pGOYyFsnAGIC3gh63VuoBqhVno34es3H6+AOWXwNuwyXr9Ld
3B6YgLzG6bBGoeQSsLE/4HJIA04hVXjThXHRx8HgD7gdGnxUWwaRT0SfJQ7HuhvkAROGH6ozQQNP
dW9CFf6bWX/lfqCRfHSzxv19Ws2VgP9MX8L3SSWrJ7jFJNTDOh6bp5o/xNE9QgCiqojDGV6MEqjl
j1MQq3MrIkfpYmYtZ2qsK2yLWkWTxLnztO6IsFGbJv08VgbIj4XDY9IFKKDScD8yBOuIvNO09UEM
e2RiLZ2qhnnJLRkqLsSUQi4CdUu5y3F4NiCLWlMdYZTQsZJOO/bS4r32aqHPtR1J8n7ji7mXrTsV
AVChvVGWRv3Ukxs8ULdcl8+vcDOFiW1tjHvLIgUY8V7vPo8EeAA650+tlV4cRXqgbGwUtW4PWu0z
2JWDj7O28wmyOXPSuisr8luM6VSV6WuZgx2i8RZ2XThzDoo4/2EQhisI0pFF1X6amQgy7Wtj+Fwn
HLapgtZJUB2FKlcmUo2A5aVKllALUT6yGo+5JOhzX0PYnOaxMckl4+VpeirbmA0KxWE0PnCXhXNF
VdSMeqvEF+0bag8fq/sKK/QcRM+6dGVAdm9PCxdWmHDukWO9Eq37vvHtgFxlc+TTD9Nk4bMinwkH
hKLHpVcXCKhZlTSGcLWhqHuJUAP/F7sXxtqn1m93N4MEQVs/QRaTsg525Wah1mWIR13TAB1K8RWd
PHF7EaY+3rCDkJMS2jE5FE+/s/d5yhkDSlTJICRwL0eaj4CFV6b2Ku4Qg4NoNJuySsOy4drk3KOz
X+fvxOFls9k3JL1ilanRVS1ibr7WY8Qg5Z1mz7Zylgrc25DCz/QzduvP4sbGbp0c5RMx6ntQ6OWU
+lN2S+CC3cSmbulRsKzUgGdAEZ0gAdhOHIYzvfvBEdVkzsOJiaKO1a/hLetfO0MtPdsOy4Ue8plR
WT0jASf9BjilbwDEmr5+vrAlSF1YtL7X6EeIHCenzGL+D/9UbMrWpV2h7JcpOv3dE5VMy689wG3a
cSm/sK9yQbRzlsg2qWr29g2iXbdM51YiJQuKpdN1MW0Wp6K0DnDxu0+uHD8MiMw6FDGIqlBNIGfQ
tk9yOSom7M9fMBUrsH7ehO0iLlvRuATY+WOfIv49h2+r1CGJZ69gLwyc/dsQtNLxETG3t3EjaU28
GgsNQPy6m3JcsJIUxwrXlGIxdtB7peFMRbIqapoTArsbtLBTvZ2QZ4JHzrUUgu0bsEGzVTXKfI88
kMp5eqLOoc+BnxawFanJ4NAyYFlcCVauzXvRTTN1hHG5pJ14yQyyY4ucJAdLaeXo0peVR497bUVP
KtgooVw5NcGfng/7S77PMnOiKf404CByQXskA+y1S2yBTUVmzNdb/ErjFhHeh5slFu3S48tHJwFK
CehOE/h/dwkQMKWGcugcSg28377XLivuUTsX3VWVhD1hi26jthw8Vn8MHc0fHB1RfLVJBDaFyuk/
FGhcZvFLvJoKmjId0yB+GrC4Ez0yWAi8aup/HJ+bJpGU0tVGNs7q+zy48vGMEfJIfM5I5MA2cYWm
FNpekeZOgaiAmOuETu1nhWwbIEgDym7ogyGuCRfZwyrMm/D+LC8fYUwedhKMBxaUhY0HEujdPBSn
uKSLU14jwu8mKC7hkzDpw+RaUOaV6/OGkxiVImwvKUfHQWLqL+jwkRwMWACZzt/hFELWnV+cWWFW
UsVnbb1d+xZSjsgeCmuK7WusZE97ISVJIH0FLIySjhUvtj9aLjFqKzKlKNkvFEyzZRkKpuRDtz/G
DhFk8njh8Z5mRuuagkbAXmNyVrgL/fKLXCl3TIfR/1ErvkrFvII7kBvoKJaEJkveu+e1NcslA0/H
1uM+G40MhPu85yDG0wMVEaeJ4yR2fDSt0zKMuKF7opcNG44zLJG1CSBSmOKIzgurZ7qiUC8h7yUI
JWsF1hFY34YiYlPxYxdSAUNi9zCzN5PshlcuDHVVDrbsP1sPp/6B+AcSI/qzU47DAGtp5kuTjVdW
DxvTEOlGDL3lPj1HwA8DbpM7rbFLR8QM+5LjdxmwDAPPf7GXXiWZt/kHAoPzYDq9bxtu9L8HgkdX
5paScJDh3y31Vv2Lbaam5KTRSdiLPR7kDlB4mey9R8Ov7l6LZSO8VtzPvW+Ykhqyf6+kzlLePQge
iV6jQeuVCeJ6hNg7AE95Jrl6cTCqj+VAs1os4mSId9a4Idsxlovj+/LyuRWZb5hBYaCa2RG+yC6F
CoHj7hLMTyWVYzQojEri2JkrDdAzVkJ6Ut4vhiFl7QC+QW3V05SWploAdKVEHVfxhGVN2DJasSUP
qDYK2m0tXJTEqaoI0hlQ7yuFGDJUgU80mOHphoUbUkL3BZuPpFwGAdGbaTgFZWsEPyYBubN0Y+MX
EfUwWgI7XiFi6w/eKoqpZ+gd3u2W5/tVq2FBFjPSxxZ2ggH1ZiLGsUU/atDvOpTwon4hAzjOvpk8
gScYb53z4LFbAPzKr55FCWmiGP8c85F9ACKDF6Z40SFo/9sli7j/JKuo/fToBMa/6Vu3sJ6HBaKn
r5kDzwIjzKAGRvAd5SN2bf5SfK/q4NusLwqdxJ82dkla8O821e2t7SlO1A7SeKcx/+RGMSpfnifA
F/ZInuoFDG+IKECBUaf7oJ94p2r2eJlHYFj2LOtcY5tcuWCmqaHY6C+4jVSZV1rqMMeIXSWMfS2v
p73mx5615Y/li6cVDdK3dBZSiAI3HOhv8iTz1PbkN9mOhRSddyEbC4SZMkuv9xqYRvloLpSr/pnE
PBp1Jf59o9AEOYyHU/DgVnOViQophy0I1GGXN/Cc8yRaV5iLaa2MZqmvcR3Ka9T3ttjSNbVKNF1e
4xx152pLNJVvxCu+4kRvcBbsQzWe0F6MBlQu/FFddNSyCOHY9JbaM+d4Of6AcdiHoWkXAhzAJ0Pm
pBlJIy8J0eMkVLX4rpeF0E0V4FEGypcBui0Epin7svuRW/WjeeQNY/wIgZh7H8fBe3nQFE7iqePH
yXfcMStl1jBjKWQJlJkKXYkQcXDZyrXq0Z3WQ7xTMfy0bHps5w+WFSPGVXOwd2pgwWGXeN2LXW/j
fLamJUebzljtAqjsjy3R9rfVAY1NUqBR9QEnUU5CetkuGu/XHOPjBuXCpDKq+sZYy+8/KMR/4YG9
1RKRsrMBa3l7vUZUCCzzPu2SckXDhjLgP+ex0jbj496q3hjEmYk3c/EP+ely6uZOfW5i1m9mcQHz
Q910U8v0LSqwbhtaO1fTaje19FSB5YOIIaP9HIjuPpDcoKIsIUpzqioY8fa0sEJW6bwsKWQzUcK1
8EZok2d6P4i3Ht+qvmyyHR5ztpqi4OzkMxxOuBUK1+cSkYCTRaXVsLPq7LlfKWjKIuKW45yYme7t
ID787I7UwvJ/UARAcDC/fti8UqiSHhwHrdV3n84Wx1/TPcDM46PlgnsiWol66mwWU2sFVmYvxTM8
N9ZQE4O9txlQfm/dSfpBxSkAFi9ZPZMI0b5LKYlspGgRqJV25jVgSFcCaVYqaTHv5CRqfXpLXIB5
Zi5YEkv6MhZCxQT7dHz2PhhQADuR0hHkajMB00QO7b1bKlwzkJj9UnfdqHx/VRQle775NJNoZOJo
vmAIznm9dROBwst3swWhP7cDn9IDm2LnO1uVihHWJR1nrifG97RkeT5fsyJOOPm0AKMQDL9cVoYH
fS0jjHpzQ9/ctKlc8Jr9P3jNzaeU8Lb/ae0V1II8rjUoYZJXJ7Q2DwtnbzU7A6G0/f50eGcGJkem
raEhqlNZHW3ladJ+adVfi2e8DCXaQa0ydRyCXyAMZMkD5g/dPVNbd/tgRVZmWJt3rDl8dL69234N
6d65Ais576OlpHbxRef0LOzPYUycDIrK963zF81pnMX88xHy8+dJVKiw7rDy/KoXgYXpb0GYjRMM
GLOLUoaXaYtgOjGbzrJSTunvSG0nxf/KRaW7J/OAI4h9oX/ZJ/ERzAVgjegOJa6YJf6u9xndq7xt
MIauGjxSrjEhMkXF4lbEng4JUL1NfhmzIF6FxrZhUxCWiMWZrYCPS16AIfaMZdO+7fXRCGLS8qhf
VM2t1EBdhHuzXa+u3wj6jjZRsJqtHwaFK/EdjPHsD+b5Xlc1VtXBO+cEJX3cv6JSlv+/h8BY9IyH
tuDvkjZOINIwqOoEdMLhYyX1MU1iZ5Nxs3LM2LFVb5Ep2y+hqxiEGN7Ak8RJVVOE40R5pbVj4dsV
lQ9CSHsuxDGAU3gX4v/WLVd7pmeK1aBER9+R2w+7SmqDymK8bv9S56Qw8HGpSHlpvt+AV6iaky15
iAxtAZNsAP/0sipcVR7zwgWZrMpTSsHOU8QgzTRY/tVvhNrqwGjUTXfzTZkUJP/5xbaedOZbaVjx
PUncIcAntvpN/HTd2++XuqYNh3g7ai16iiO8fQph11N4ifO8qS5D5wKlZy+cKEeYZP5VU0kUMrnk
T5X0O6vEQFopom9WwwCrh3wCYP/lXqyuz1TroptzTf1ASOednNAmwJPu4RwzPqyN/6NunYBauvYU
7nMxiP0KgcU3y1oJYDYKDTGI+JNLfszb5jVksyiNnTgP7Z9GDtx9P+jM3iasVASNZf/fB9jHbzVZ
5U7k7M2p3CUntoas3eBgZl2DABHFzpmpx/cIhthIrJhZjI0EyPBatOhDqcYfIUQPO7zha1DodvEj
95fAyBhXcK2NgJOEHXiRYyOzVIoUHZePg4GlFGkwIo9li/6DgXoot/1QiLPkO73W6KOy8EX9mdNe
mBd+oxIfg1Ok2oOKxyNBlJunBTwvxoqYsJb0b0R3MN/U+irWz/q1CU1uJGyLdgTXyKDWhR+/bb35
MY6ZUSgTQerRj2gbD6H6x+dhgOGvtagEhUb0CAYe0L6MeZcSQdgtAq9ywYDI/WhWPK6ALfbkFfgL
Bb7DlNV4074aoBEknaHLbICL/B4YjvC+OXtD6nyYJqnXtALz0to1BY99G/TfFwECn3J7zd8gnQvq
odzcIgViB6J/SrR3J7IgClo8I8TX72tiRsSlQeZrlM0qGL8YNLW2QSNTu8tYImayz1pcgFUyPvQF
ckf2TdkFPhr5/7AY8BrUWUCIJ9jQaBf5Uf3/cEz51sMClkdF+sLT52Sg1OsO5VtaQdSOtjT53FxH
9/2YtWmP3ZEi17bgjxNMD305qLMP62vL8yXdbAS1mD6eDHKw7XZb9J1y+kReO+gFbPDBMTxoApna
qgDdpQOEliQPk+bk9P0axFfDF1rSqitb/dZpDPbUyWYB37X57CZqbahBdl+Y/TvxaUvY4tmr5sfW
vLJNYtO+bTvmjO85kc/lVMFggVZJQBiRuQCSRgbYz5PrCEgdU/BqIQSh3X29T0WzPlOj6KSHF529
DC2aDJoBXswBkfo2My6UmbMYjMjCz+P5A90/Q0t1ZCwt5t7goKDXV6UUn/m8ITfRvYT46ixmvkp9
bmdcDJNy5MJ8cfPCCv1IXtTqVkXpasOwDLHzQ8peDXjhIjg+BiB9qa+79pPut87KGxgYc7xBEh0O
H88pnCMpcS7d8MVvYieX9qJNSh9As7Rwobq7R+UqCMC2E+Ltn/xH72xHorc4A+eo0fty9rEgCBs8
KCk1juYW4DUoefwyUt7STkSBIqk1tS38zCjl5wo0vyFRV6HCNMVoqsZJtlhzwr1XPsMugp0NbaKh
/4O0bnOSR+VC8VRjrYWF3QfsdXq12b2TfiuMidzCPyZGK11qamOz+5zQm4c3gRxAMksOtObUKB5h
1YLST1Oldit2sSYXXSKzGe/PaRQqYSNPkQAUr72jpo2HrK9Oq/p6X8JZ+GpQruLeJ2sUJLGFxsPr
6ovww72px4OZLuBkjARwc/8m9CTxmP63caavMTk/h4j8Gum/8yTZxfLi+TcsoCYsJ2L9MBn4RGcz
VvOMa9bgFNZuIL5ZM05USfTpuAUg3xVOdK8TNEmyJTdxGgMerJ9roHZRi7i3qJWG0nFJCFFGVK7f
xRXftfFysUbNWE8sEwuaACVuSVOPt+M9OvKuaKnQ49SS4aYKcGnfenwP2FwL+q3z2i/diLp2HYES
Ktlp14V+0NDyKicPNXGcBItERunXPNtfsvQrgwwk6SXu8hUdfV4dqPLD4Tt6gvp5rODq9D5hhqSJ
ADmfAxmLgqLv0DpnnpUBK+bE2L8S2QFCMnQXbvqwq1a/b/vdJ86fttwfIgew8UjNg6vKiayWllxm
ORuIISNNogQl3NuTZ9UBJjclkdKd9cRiTK0XGKN+AdrwWC9bXY/N5zed8staiJJYGmXKov0viNUn
UPVLBVtKs1L+6H5Hsq2u/dEqj54BTJfBny03T+f3wzhMsFdqHP+RhKjoXIrpWhsFSNf9K5LdohC8
7iLKkHG7PWtfHM4UcEbeDpFJKxeGYQ6BeJxvbC8o/r57l85A7vE/2mK7ce2pXJ4VdmkBAqAFlb9I
3xA32WfCLF02Fic7TYvaDhdNf+eJEvNaUobm4XnLGVgqDxqtFta4UVIIKlavRJB+tZ74hqIeOZCb
AWp+0pKCqdXPxxQWC6o/MRhfslam036jayHx32eCWwedT2m4zxAB53Y5wEoQC85bg8bcSSfXpamr
dffBti+/OVYoqbMRMb8rzNwsNVseJSqfpSgtjrrilaGA38mY17bpcSm0gfsnFsrqD+9Ia+JqbTan
w3xiogU194Rd2GrmCmgvzE24ZFCMR7IGOVoXoH1VRAEa9Cz/WOKkqol2HGq0ZAiVL2a5tpDuNzHN
pTGET8mymH2+LgNkc3+UA7Uq9Rd4SDuDDPBEIIz4pxtjsme4xfILdkZ9uVq/3g0un36iDwD8jrnf
zBZbdcgPEkB47NXdWMVmtyENlcNKqu9VCaXUR34m5Y3Jm/Z1VIpCcnCtH34kxR/xskoKCnjhivp8
wXlroRn/3UQunHE3DQfb+lj0nnUMUTMZmhS0oeY5WDgB/O/sTGqarCfl3+KzZ/5pDC2+7bGwAGP9
1JfjdBUk99TESO3tx8+iBdr236kvr+HbXQJ5e0jFriMpARY4oGnWedmFatHRn8DxpmlZ4Xgh0nJO
/tYHc7jB6xQQ2zjJR9uxKsDKQvAMa5Fl2U36K1rM6yxlWtdAZKLgxCExZfHxMutmMKtBbpGLb9NQ
53RmdG462BDE1KkJD9n8YUWrLr+9Dtc92oXPE9xNz4k65YFSS9vT4q8No+5Zv/GKDs7NOjOy7iOh
VQOafM0Ff+M4mV7d/9CgAE1g7WWzE5teVfqdOPzpfBd2Ns5BklBqY7e3nNY/g/yaNS4mNqBu4iX4
0pwHctbCwT7qh+xBQJr/SJrmEa/XKsVzzs1ejcYCQIA0XQE+ICMB4fPrg8bduFUPVGHOPDsNQMml
iFJoY4juxDWFJuRA1+A22xvR4Vho09hoBUDyG577w3mIChYEYG8JIDNd4MJoLf+FvE5b0rr+ZRN0
LktO3zV1YMWHzcBwBlMa+itg1I649o4C9psb3W035DrvNspNWmAzuEvY20C+d2PayDwrJPLpq180
o02FdGzm+i0s7WPWZvk0UDJLc5q4oBHtTNGfSZQ2eqMhaRNFNLVcvCwBH1lnIIMIOcdBJzuuvaJ2
kv3hHvAfpfg06B9nFQXdT3h3IUn8fkw/UJgCLthvSmSJjnYqXG0Bf9QvPFXLaWpMKbH79CE5Jr+G
h8aRHh4bhIWjIYQVOVmKYrisWhqNfDtA4/KirVCL2iIPyvMXmSUJhQL6P01rTtGo4bX7FkrkB7Jh
mqje1Mk96IuuatgVqGyCEdBi4pB5fm2mhsFPZXoZDawEoRLPLpnWvYOv9pCYeJ9L3E4LbqBmXlzW
DNW4QGTOTvOL82RhoMeVvX772QTVp9B/chGTM9FypQI0rkHtQsQ9ydr5kULINhbxtITRF1vtIQeV
adhy91w+okmu8ypowwbO+4nIX2axHdBnIWvjP7/Ph9SsECdPekr1raQI+U9aRPaO7sDdYDx1aMFd
HO8bqgU4nuAJ6LfX9nzcQUNmHBYQkw8PLx6jBpuVzQod3PdnH9yO4ODCrx7vZyuFcgdNyYjqXFND
QUlzG6kFGVmcQJx0MhbEE/fysJXFUq/SlgQbjn0Ma7MF7j/UZ0wAZB1LLnQjo/8ciZogGKznc9Ad
xb3ddCwNkhKGTMg4DKPZ76hCMj3cj7sfORgCO+qjegU+jdEwKOEN9+XUvHCYfOWBXdYEVodss85T
Vrj9DG4rTRLD8OrDAVm6dP9PO7uzdy99Sfv+wyn5L1cuRz6jBz4AAKsfP/AbPjgRyyMMzKVTQCHX
LxT/5+WZZNyzHdRKBHiiJJxqijres9vChKTWg//c3MegGTNzhaNw0KxDJTxjWNeEI3G+dbcfe4Vs
l3r5m8lAkXAZKmNZMRiIper04r4OGjdOVwips9s8T0izvI0D26mCkrBqk1YyjGHq8kRPvoYPizQ/
kj9A4WvsuvuMk1eN/dZITVxwMSTYv1XDAxz0IpEauZ8NdYtXx90mlBhwiOccQIWcJSk3Sd2wSlOK
ZpBNn1gYSorbVfsIo3yybppoLeK6zDq1aRHiWqoeVnCg2nOJJgbqn6NLHhGtrKzpX/srxypmgM+d
YV6isEsazFoeVvZvg8bBX6xDnR6ZoxLM3gIp5yYprMBfo22yypm7HmjMPJonO98rrgk6iYwvlBAX
GuivCbncpfMWXxzVWD1qMg/gzFZQjjsN3c9DTGnMeDz+rGpt4WUmpI6+GtXkPKMDelHg/9r7JmYg
R2J3hSe4nd9RVy2XN6+i2yySd8+6dsFoGkMVH5EjvL6YgiL7FQLF1dfMhH+xpDz2ydmISG1NJLiQ
Nh7WNFjN1bvjhm8k+IWZUACoJ1E5rfWnF/WUVRS/AXIeCNwtiY2/IzK+nC3rZNRGcXAOK+nG7rN5
hcg2VGYx1IGJjsRMGs+EE2/t25irMJD8ejkSeFwvgI5Ch24FC6qbwKKEMmErOzXuXcfeM/AMq5kP
dtMwcYoN+MHgcoj/yTqSKYg8pty+cE4vnN7RfdraMyB0sEFU/hZcJ/VWSXURuJedgFpop0cGs/xj
WKpadrFdcjwgvfz1RmNXdO6+aIq3tZlGLi7lhdglCWN3NQOEFi8V17VF8Hl3bWD9pRfFlqb9bbBR
2Tcljv09cdxQTTEQceNEFZcb/DFRSVref5C3t+LlAGzrTC5btd3rFCZ7yfh15Lp25AmME81PErUc
meFVzlHIM4rqizLhuDBPTbsm/nF9sm3Oxn1BlUV3+tqIwtChP7wpkFysu9HS5k65LsLN97b69UVC
gKlfpTMh2ufFRvu0b3ppcP9i3IRWGuMeI6zKc4EVZXEMdJRuwwZWcilXaMBzUa/TNaqrT0G8TpNH
j1ti2PQ+PZeRXY7DLrcVJB2tmSILUq1xvpPuZpmso4f5p1q219QSQ6Mtw7/gOwyy9378RLEjIhmA
i3+XwcHDBmrFjjptWnZcCCB8e45G6ScbR3KfkyTaxLxC1xr3tsKz6LvmlFzXlTvI618dUKhOS0du
TwEicATM2nnEDpnAD7liBn0x1apJbkfYDgve9/nCZFJ+09OKzK6BUviYyNVrTJOtMdhrXYAEWS1v
/PAgpmlZMoh+BoKJwEc7EvuRwRD/E9YXs2JYQbkke9KJblpbCOqOGPEl1zETBsYVA3dRdwSMpoy3
AjPjSr7HH60vlfBSIvEg9d6Hteh0XfINzDAVUBfKOCXmk5qMpM4NV9lkvCELruIRwAl/5v7B1WHP
BFc8bUoI47H1kZxzZolnqvuoZBO1zQxs07/1e1oWPlgQq5JFexEPo1PGZYkKweqOyl1nJpRAvV1I
9wlwkIJJgl4Oix0axYKIe4h6hbKdhTnp9FtBv4yYDxZ5x51o/6hzFZ+VL+BZM2OInEYG9SOzuBmB
azysaSWVIV/mqsv82me46giHKAJSBDvyQ4vSMrCRT6cv29/1ni0fisd5B4NvhZoHbQPUxcGObU+F
0ZJ75RM4TKyxdZznrDTQaLNFpVprUT2mU0p2GTj0j71F/gGyPfI5u9RfmE6dkWIAJhOVXUZbZNZ+
WBS6NkzLU6qAltHVCGdOI2qWxNuZRLFXk+4xynShfkcI0XC1rJsIZ0RRjbqFX+P6RdH3USO5Hhtu
x8R/tu0h/cw0WGmtmwJ/vtDY8y8w4HoRSivwPgGejj4fA6vvpf/CpXZo6naYbJ3gggBv+YhDMM9B
h1DKwlGq/8WO6EHhyQbJTyCNLVjAq8dZNEtdXAtPhRs/UEqkAPuG6bFnACL+Yl89hp203m47z62j
MD9v7VNZHny+69KlHTWHH1AOHDMcT6hGWdWf9aCUVmuj7Pc9k2HQkmwQ26jq/YSb0d6UcdOkZtPf
aLRd3UUQPaQeip6yOgHJE9eaN3e2qLoSzaAXzNHU3qGaYWeqFN+aCjPc6c5FFKnVs57sCTr5Ry85
6uOkY9evM1V5uRdvwNR4BdLHChZjzO5UxaB4RmMC3XqisxrUzqx+/s1afQc71IGkyRoXQa9ftxGh
gXr1LH7jmJuhUkvsBoRpNfgZ1mCCtm/7Kv+mMat6P3yMZRHLQXreGk+C8GTmyWJvP1hKLorOgIVG
qayrrn4hepkKbzKKRPaR7n7smo7F2ZGrgsEghtK0uhGe9/olc5CXMFpkzxUpYD3CxZCDgzFH2aii
oZ9mFJq+pCG2GIkOw7ZkVBRi4HFup9CONtydhirhWHIXopC/p6t265LX9LuAP85TcAybnGR31AJB
DHnBHFCllEKx68a9vUnJXtwlLDhXqX/peNugpTFpN9tnA00rH+295dfroc/7VsumWoB5sSygn8Tn
9SBLmChbIVBTy7OIq/cqHgBExc/W/n5nmH3Telf/QWob2RBbgZQHbmIHNxKEaIZso9s1IkDB/eN+
lZLG5mTJte1wqeCcj8p1G1sGeJ/a0MiMe2U1szqUKG1kZSes9PCwUG3U5M1/k50nCMA010GYvN+v
KrFgvtkZ2ngHXdq5YlIoj3/48NIIKlY5vvwaeb68B4JUacMOzpYEVZzgZwnp90Y3kaoAKbUWFXP+
N/AR/WypHCLxtOx0eikLJxUZSKzjuInux/448w7K3Y/4+dd6iOmVX2LUmZD/KDyrOHTq62EN+7Vd
uiJtEsctoRk35RltLdVnzq+jFjjB425zOJvvu3wUGoDXjCU6VZf6L8CpZ9igzrE+qCkIjgErH4zV
UYJ/f66n/KF77T6j3TMH+dWN9cRXYUHk4S44d3f0mi+R35zX8VA1he0HQjahri6RSoaLs3eIZVPD
WchQsXVA0t0MAhqS8iOKPaBa7E9InSGDTxw8mM75Qa754jTqlIcqqT3AHgnYzLtSNXuxA5REJY9m
1b5MnpUKJIHqiWGGyRoc7Y41qhq2ea1ENAi0mXmLW1ZhHUQuLxES6R8NeMUKW0GmhVYEdfXvzKOv
Nql8ysnQNCMpXkGDukmW93a9lYdCUrgGntwGaPE7rdnQAB+cS2Mvfhiy11iTcqRUev9oO5nLyoaz
zR6NEORaZgpmi81b/PV/t+phsB4hGMZKIx5CBO4yycHWWBn0xUhBnTW3s107VgYKDRc4tOJUyYy3
LbzqOaulJ1vKObGWiVHfLWQskZpD4CLIWUMBLPv0biMnnY5dz9mCTI2M9jMt8jmXpBSTToD5nNAu
9jIlJgXZjUU9eoWRiSGyTyjsLzn9izUSC61Qby+kci1kH3VhVI6AVjIlc1Ron530/U/StG6LwF8e
3Lma1Pr422kZl3mVcUIYTaxW4Sa2lW+VYAvkdw3yvAT8SbIlJfbh2ffhyFYqlpORQTkXpapn3SCh
KYFlG3lqBUYsVgpk0QgVkS/Cg4KSaGlB8F7uRTqmBBxPiMjmU1m21GoOfHwR1x60G8s2aIYSVE7c
Tyb5fAcmqSFGbBhO6FGcUlA9XfMHgiCl64DvqLoc75aIHeoZKSQwt1XwqvLu8s0JdMTH7u/ae0me
N8RyLx8PCno465m27kQ1RoRCfueqIWq9oT0/w7bEoGp1pRXTGMIGAdd5vkq6ht9/DTVxryQyZR6O
H8/OvA1t6NnpX4DdTQW1xJb1o1Pnv5zldtHOy6xdweP7Ulf2uNyfh5K6Yf//zR+9h6lxPJuT0lf1
zL5B+Htl6xwBFcV73rT6XHqIpe6MiKxHrnw/YhLiNiCHLcHIMaHsrakWnB4fNynSrBZnAXfAwJWB
XMYe85EKRuy0HzevW9aq59Pen29jBA+KlgIf6LOlex8yMLgglI9qMMnr7MGsCI1t0ugEJMeuFXwq
Qt9/amPbDoQFMuVncBxBjE1YjTu4s6dv041gH/IWVT85YMDAd1CSKnhCtioSvmhCeojWKaSOXSD3
D1od2WdEvaKl6VB2CfiFrj4ydjZgZOWpETVqrbHdcVVuTQRB0SwFHOdhj/coGTQYEUeIgXSOUFyo
mjBYPKFmClPEYGlGuikN5Po6Xhhrp/73hqi/BWQEfWbno6djJ5G0nDUvnsg008LFVfki7dmNhzsx
lNaFzWCbiQ1ASDkTel10w5Yre6iK0owHX5ha1cCZzFOLaoDyaKzlck69fHQCPB2EWYyL4wk3ekU+
2QsVB7DjIP3s4gpKYoQOjYeRIFT9hNjz3mcWMJRtHLwflpY2H2Fx2RZb/vdJyUPxkKIKOxMKx8Ar
//XDOUwTYYDjmLpPTVasWXlxK+OK8jEfQBol/f0wbU1wG67axAGIK4QskXyAO721uJUPQmRD1FKK
jcSa0nj5p4ffR4aFY8nbX8qznQqgYRs0el4C1pHJc0hGLhLZjpkAqB3ggEAE/svrminfV6XDFrhp
HX08ROaVd8T5C3HC3TSqZBS/DbKer1G5/CXDupEfOmfESTvouWGpkZDtjpUIhv1wHoLACj3LHy+e
JND7KHzIt7IkSvjKA4Y8iah1Indl0dukaS3djHltdXBSaBtxypK2WpmXQg3RH+ah1GJHAzX5oY/G
5sdXGVTohEWld99Zg7p0MIsp4K9iEt+S6V8nV6UTHBqaKN9oaDx+IxxXWDY1HmSLdvfGEFDPN7qo
93zYRT/lGxpWaCwz/BkLxPLAgFuO8gKpXqwFC0drt0A/05U1QdYjlnPWvkeeYd2ddoKMxYiv0cYo
ZOMpuqrVvp7m8iyG9K3DLvBRxXGtrNqWoMOltOrEB8DZwdeil96WKSThJHcgX5tdo0FK38YCRqjg
94QAu8HTBFdEdwUNA531flaeZmmFcs/WwvSmkp5w+FNJnQ6Thg7qK9ga+4au+TemcB87+k40uxCh
KQXtOMpVsU5eHm/KBsz56uf7CI9VXVot74QCmDNBYMEl1lnwMFnFg+5s8C6SLLI96OVpH8eqEBAx
m5aZRUd9IUzhhU3U8PgRoAKZMIOfjxHVDZfCqAgALJnObvV4+nH3hVQg5Sng1/ud7BjBzNiblwZ/
zrcq2LWa1B9M6zeffLp0oPYBfISI/VC1c+33Zvir6A5L7fBdajmVAGUnP/ZMP4U49q5y+sxxCDHE
eyHT2ASau6YbjJDHaRgQ6ABbaZaQf76Hxxn6B0RPYPlzt+MdRpALXUnqCiXzzZnXL/b3Uii0odVX
QSdcqhBgS6x5whmlG+q/w4Ch15neBbYdvuqFWTkip0Qb1xUhr3oZPtRrLFoOGWkTO5ThxgYvQCNy
5vG25S3E+R2kf53ewIbv+qcsLOPva5uDgOlUM+v2fYmIGOLVP11wnUCzNeOeFX3PXqeHmeiQ1azI
lrqragZFIvwxgOE0bXIwcUPi8cUrBTwOCshNNbQ8yNsFYjhRHaYnR03x6V2bUvVEprLOePZ/WC9F
NaP9RGyAtbIsnXz0LRIrFQ1i6T+W/qCMQDNZQIQzZ4DQx4Red6Jr7ShW7c46UgEds5qnMPqO1pB+
DldNS+vRhcG1lV5G0PMniTJobN4Ah2cE1vsr0Tp2b6fbFmjqqrxoxUe/w8cK8eSqhkNT1obrmwPU
8K3B14OldmNkFsBCEcFjUIxP5YGApFfAW8GHqoR/t/XN39va8sKuUfAoILqvkmijFXvxNwkWtWmG
Wr4BDTKWDmL4KzkmKTIMlkEeuTpjWizq5JhXcx4Ng/3W2fzkpnNdDmKtVzS6X4bXBup26dt3MRBz
GwtFBfC20jUIzDy2ZbwputCoISVejV+etrnbZRgljaL1mJXxuR8edzYfvbKMeiSEyTBXtJlausmK
ytXR7CxaKkOnyDFwn+ajCHw0MJWYYTiNi0jdEAEDdW06/ioFJdWK+CTCGBi9MID+Y3aVfcwdu6pt
jzSjK7CS7V8W5G4XiKAM0ICH53TyGp/l9A/zYm0HgRUF5lQLAaa/wsoDRaLC2aO5vGyWBVXRLOS8
FBBDKMWjVkYqZ3pn9QqU5h+nnJb9D8Lj/hE/sGIloLOCRNF5fqSk4b4drzinCnJw1R6Ev1m3bmE7
uULgWvd9/pdW6rYaQX1KS3F4bP6ODGsJwlmrsfHo23BzfKF4QSOFZp2JHgCypCl5BELEACGSFsMe
/7DJAlyH2M5AVHbIJ4T3iZLI251Y4+FwbAE8fLcowUa7GAxDWtEq9j1aoYSNDgBX4vPs7I8gJnYt
43XIU1/7QDEXfMlretJNZrrgchp21SvFO/ZlZHrdhTsvIpF2+t0h66m6iTY0s5KIUXdAtLecRr4/
uKqz3UbUY1i3YghwYXKM3jMfpEPp8nUicrwTXl1P5ye6hFq15mVbsW9iOMSPTTy/NfL3oQ8E8Xqe
kAqVdDAxyB180IEVX8MS64lC6pNyN1gOJGVhzuDggL380h4dIBpZIudVkAL4oF/zLzyJ45PtOcUb
OuDihHwpDeTvapf5bnLO85gAhQZy13EtzuqmZy9lkCwrCEmWZjsrLo6SGP33wz33+7nfvK5xDtjS
3NbkJ8D6gsG3IXGq4WajLcvVm35GfDkydtgY1Xheccygmhj7b1w9uQKRXN0a6UK/3zjbjO3RiE/k
NOus3MxxDlDi1t+Ho6wBEMBnHTCzXnZLDNkktZk4XAUPrv91fENcv+0CxkpU5pOdNe+98YX1ORec
GcJEy9chuZpHEwNzFsPToWmg5kniDzSuePg/0+laqgJ1gm7yvjST0kOFX98/IJ9Ie2nKwHdSXTa8
Up6+6xTPlRxq3f/C75xbx9Vkf7MmlCCD+x76/dYHSd32FeN/aQTQAKsjxaYtQIwXKoSb/dMeW5gk
bxMpZOXLXym/WqVGCCif3yicrsqtN03a/WMhAAbksjzn2i6hwRYMrwuf+46IIn9J5fqvpR2ZtxkR
g3a+N6YU2Gwc0BN3I7lNttqZeGb6Uppt2QtFG6jnQXWwJARo0hYnNxfV/bw4n76GrwTjqzPLgtMn
/BF5iiJle4kMGcyAliN76SnikXvSAlp1iGTFcyiOtFmB4aqhIri8lWKz5hY3uq/RkKpDLgWo1iTu
LnNaL/6F7d/slt4x8U84OXPR5Vy4DuTQtRHLFFGc755VkWtvcvUVJ+ENewKQpJWobCx/izGA5oho
IZ5ALeQVZ23Y2p2rHri2RIDTTlfqxoB3EcrGRS0dGbCRFbbt0Zs3IeERTE9wCazQsbEoHGdJ1DwI
y9L9THGwTpNQ5DtAX9w/n4FsNsNTcBhz4yKwfulJHa/Cskv0gaMksvaOD282Ieb2zbPrQQTwMMMM
nXEyQkTgePwC1SlBtniavyjasiTHfVapjW6JqQU/Vhysxl0haaODsYIK00tnbxC3V9TG9wp1BIni
1t/BLAu9LnkmVrsgkyvc6h5aYnfBuPnu0tgsDW3J3kYUpWxbr3eotQFLPOSpJkNTBNTtXBe0r7Rw
CFJje41MLVCymLMOeVyLBvY+Ki5lnmhyHUiYlv/Yxnm/QIpAl8/LQOVlH79XROydyvuKJQHRbWwF
J5tKVYriVZLTwDhPs+ZY7t5uD9kSqChA4UBuPKwTc9uSnPBheXqWeK+kGeUH6qVrkoCAbdHXgp+6
PD5BcH/ZCZ3CrE/OmAWEXNp/SoW0GMA9k52iFjZUHmYfXxSZhGgdFpv46VxVyjS25ejW68IG6hTx
xPDcJwjq8d6vSOQtLRlDJRy1hOQOSYjEJckmic3Mga68IhHP8oFVwLR23gggRO06wWT7vuEtCwc6
tuHbNMM4F7/iV1rSgdhWG1pfTOdpUgm1PxYfHzBVJfYNi+jHuy1FeR2IeZtRMMVKz6F2WbuNbBKF
gsiIeZ7IPNUMUm5YGmti7nvoqHP7/EtCjd2+AJIH/aILr+2F1RrxnexrQN42hoHgtwFsQGa/TrLR
XyElvTajYh5r5zJmxBFacSCEbcOeDUt+xzpUrAkjfPonDQBf8kTnBekFV4UrVbpAVphFdn8mjI4G
AVo/f85ATmT2mQaL5y6gXdeqftWXGe/Ud8lhW2pUpKKLsy1amrMjpBCbAPlyvvd9uMEKhmhTIUjU
ucgvtr0WNmBeTi5OK+RpVUCeCle3Ee+O3L/TUBc0M2EckkP2nK6pTKv0/XFwKoZ76jQlzan/Bq42
EZ0/1g2wJAvOPmpMnrCK+qsLSJn2woNdlYYeKPaGP+ypNPQq/36M5mHt0ZcJbkRkS473ERMgPgEm
FJGr/ZXYv33WHkC2P5gj3gC/EhpbBkKwsN8Fpu7oRrQgeHqC5A1xs5xSzbyKklWjcy95pRo+thAd
rfpDnz5mQVykY7cVOFBucAalDML1cm+DfSFw2hJcwSehJ1awGWNt4GlLCADx7e2leW+lRMoKEayB
c1ogZYvoBxdNzY2omLcwuJ6Cmnjr/A78XUi+jyYWPeHlizwSqeESR6vwbHHbBroZqKDOiT2r35pu
oLpnkxYaA/LrO+18OoCu7vqKZRGhsnNsoIWQfXCzY8Cs0XxMureffF+ZxjrlYScaL5GBRfGo6MwT
A2XUuJ4tJKxgERE8GTfilQdkBgAhGjXYbHlTPISUory9gVb+0Hca9x/hP88MvttcafprgwMJNtH+
nkI8y/PhkLEcxA7gyEkX8D8OvHhjeQIbhVh9sq5WvpVX0k+CiFVxIx/qChf/G08fsvB744fYAVm7
L4xO5gLXCaA9VoRWk5lm5GdIUoKN0BeWW0nirXGm8sG1pgvFnWf19nLb9PpSi48f0ataRdBxXe/U
jVM8SFCRcZkWq+Gyey7w3BBZoPR/DUYyeAS3SKCywXfUHFoWfRy8bQBw36vmDnHXvpo6WsMzS6oK
6Oo1GbGpFJwlIEasPgE6AHrYH9GgIxLT1hWxbFJc2HaWzgREd3e/pViiPim0DfvZn8cAUyV9SpsM
sjD5MOfDHxPXul5RApMXJrHf4xISsouMFjUGtArVasP5OJGzcOYmUMrm4rLvEXBB0UzrO0c7Lfqy
mGM1QIBki7MDG1elbEvp3EsjWvB11YOmMRRlzac9mY/JvnG9qCWg3QnGFVDzLbOdiWulOhm5vfGk
Y7Ls9Pt1Wg5YeuRKXEA4Axi0XqrvoJ9LGKVuWw0reqO4F3wzrU9D+Pr3kq1UOz/3fqPuLqRqnBRb
hVygL8L+DWsOhkgOoiUwDloR9HJMDL8rENUTfenE2LhprOs901zmEn7kyMAg+Uk9Sgezj0bpSKpr
HnjpTO20pWXdMxkhvVk1GcogwpNoGQuoVWfM68RPPosrveFuso3FVTYk1Jq27q/Kni1iCRb07e8j
OS0felsMM9RrAgK0ApLiFhzPpVtpgC84yzkub1gAJh5AyaRqUo2fw2IjWKZd317+RG3JTkbWbFyF
Lrl/CITPKUWAD/W0rC/4rn6y9hhtzrOJo/TQN6Qb2TbrezSzWD3OT7DggOw6L1hs9luIzS0jvj/x
cnj9ULAcnu2Mk1Js/flMWbl1nA7DTS57F47aZA0JwmTEQ+5n02aTkDPr3+pbxe3quruENQT+euIo
FENJK9ElfjSw1VSC0sZ6icGFxz1RQXp7YHWxAWfwOSom1KM6/hT1ZmCr8pCE0y3+j8QQQ0c9pbNV
kf+J94ee+QitAvTV5HFePKoJJw5tO6qLPHqmhNHu9Un2TAugHa1lPjmgGMvVu6oeymTbIjQH5Dvl
EVe2U2fhjmXuwcO71zfSuyrFkrVGjE3jeOxoGjmwCJkS+Tb31+o5HvHDVL7X+3Elgq1ctYeyIfiY
3M001jQiw7comYD1fLibmAh/SL/5Yod4xK4LIUrfJYgNHSyhfaCjvURL4CWcPFyrRMWLTbcMxKCc
NQbi7SQQ6IkwuWw+yfdeLG65Yr1hYnYdyIHKU610icZGfHJUXRDNzub1MVAuwq6tdkYfEpMrvw3z
92IPqwaXsTI1xcL2mqZqUpRhfBXBCBh2Oowgha46HO/NmXPc8r1T3p0MKaoF2lDIpQgnmaSC77ZY
0lhAYQT0OLlVmhOpxT0Nuqo7onJYnwHqDlXtNVK66svaq2D2/vF4fMMjN5Dz1mvZiTQMZ1dZh1PN
iZtvlROsnkzWGS1xGkUK4zQXLjtiB6oKR3TNjMSi2an2XwEG1f6Y5DzYOmvqnzvbK67PoSKGQzy+
gvnsZPW/cbanoJLhUc+2NHhsAPSoERFrEbOGhlBxwWmgBmskysPa6xwm1xKvmaDRm2HXry/yK6A2
rplRmP6HExMKUYYuNp266NSt3Z6S4UMXAVKV6n5zbHmB7EjKoSdGb4CJ5chNwvvaT2GfI6n5PMaX
pxNq63UxIagjGzFCL4vb8fd8G49qeIrPEwH32t9juzg9rPPFVTCyjv5tajZKuyRrCTPMXEKKEPPk
3W68aVQz0j39pA4MhwV0urYHqo8lzH6mRCpf3bVlel6ZzTvSy/qQ3thNDc/NbacVsOOLWVdigeV+
P7lvUmmo5yWC64CtqRUqdByV0Xjth1v49086fT1EM80qzxRlZruNN8hFDy6/A1QQePVeNRTmXlX+
4izQ7vK+VT0v3oBjJ6DZmzG50Oou+IGAZsqGo76xNPsns8cLBX/pbxCB+3JKHiOgntDMc99SX7Qu
XpJsnh/RLSCH7vmRXboeg816NZ7MR7OwsVW4fGBx9RAHL1k0d7Gpx2HP/zJg2KFjS4Z2g96iR+4A
LR6NGQ/OO7ypDXZfElrA4O7VoOKurLfO4dG09+KSr+6rpuHguWiCYUkseLQ1VhlN2QcNDGXa82ZJ
oto1WuaeH4fA//6/J4FGRarmyZOilU0iKgVEoUlI/pfmAWrcOBUWgz01wi4w69x56LTafl0Ip7oV
OG5S0dRVKc303Zo8NLMbfUVG8PvhFVuAzK1Z/jBXhqf20+qH3jOJWvKGBdk+kkPoee3UEOZDf7KS
yN5qEeiEQJW/GfqWCwfHzTtYQGca49FS2KFOzFlR+B9DmAGMJWv/PHyGNelR9pbViqfefAY/qUpC
WMrBCr76YOZJg+pjSVmAztO2M3WFsfp0+/mZ8KzNMEhZggTth1ecVdmAEUOqbxno7Ni3w3GNnyi6
iiulWSH2rL5sxF2eB2zxzIbSMWLTfEUmAviD3ll636/5QkkXtwzNPpcTAOVtBNgMiHV9jcIMEuyE
whAARCrRKrwdV12Y2yAjicohj7Y/vIp8TVNLx72wtAeOmZEyngCzIAXcqTcH6azUwYsKA5VwBetg
xf71AYgfDV94GlBjFUtneo8gt9/bcsfshAkvj67t1Z6SzukRrxA2IXflutJbemXXVErjHI8yO1cm
fyR3cxNu0GeNBMw42QMWuNBgm2dE1M5H6iAHpu67cRct/pmIT2XAIjK3nw7QyPjazbrRvRMBTDqs
rQMci0lsSCeizY9T9zJHxOeBNb5BQ+QUC5ECOMZNE1MP3isZFIn0GReuMhQAuTkjBkcfvDNkUKkf
CFrmw8Jzfe5LDn3uq0N0hdgXwTqUsFNNPFyxO/goxM87bc7SKrLB1ITCpaqrfZcD6dyfLah+z34m
FI539NkxSOyk2xnxjM58J4m7WuwCvy+/Bhrro62nY3qLaAle5lUFvL6SIwA+TZvwgRNL082YmwbL
3Es+MfsDyjANr7Y0ou9VPULgGcnDnLMoZ8xNTblVP5j6af5gu9X48yiDT/fSFewqjRkTxp3VOBhC
1z/92gzNleRtTf951mctcQyZ6yobdYi6t5EXJg000IPh5ob5OD/a2PMYcZ1EU0oBDcWtotAbsdJ9
9h1ix0J1yn01qMAxU4zm6dYEFRIhHOTI8ElA+1dC6W3JhlBCnkASJhAuhepBgOF3JchWs8ct+Whe
JkE2xI4foz0phX5xkbs6eqOudOhEsRV3h2czB0KUynAOtp8bya/INs+svIGse7uNHMSMNifCK1is
RfXW2fyjsVbiJ/Iw/kJ0wn5jF9h3lOmdyCAv7qgZScvKb8n1RNS/hgD3MbH4nyBRBj58bbO+HUR4
MpFBJ3Ig8aoEgP0i0fl3nuOZRVWoNCiNNcT/O32GIP0DNpAsX0pRr7/n2E17tiPhA4tZinJxl/Vc
JvEEgBNgfrZ1J1nEOwpKErkxo02fCaT14tJWZFdmKuJEps8NgWKZp7crh6TxRom8wLdZEZZY4saK
KU0YTmnmQhFl/6/N+7m3EzNERSLv33xIGFDxG6esnNhXvd5HjQhjWCUBFP930DYtTA57V3QEG2VZ
mUI9OEVnRGJ9NsmPQr+nPBUxHJ/1L5AYMxD8v3cpdnK/efgnF3siYaVCjveO6QvYt6A6gdJTBGsZ
AjziRgFhTzb4Q+HD8s5+WSt/ZX2+gjJ7yN8i5qLWzcUuFn95Pe1cDhJEiwyEEnj1x15UiGx3jEEb
E8dCMfSJ7RKVLbA58OEuzVb0QSrQr+pnzXqamAti+BVfG9r2rU/ojPR7XM5Eus3iVmVzyFTxW2Is
A+WkvyK8bc4L59GFciMd4POQ9WjOD3S4bVj05wnzGM/KT6x93y5cFlFFHb3tQWeNTm3XixPsL8jm
MOl8PuP0mBRfXD2NNx6rtpxRja9eWhTxPalwTJIk1kd7F1hCAtlatrAt4X5zE3NklnyGdaWaa5Yn
/YvFU0F4W2R6ciillbb1bImlZqw6IiFElSPfkTih9G/fEWg2FLkL2bEues6EVRRgkWJr5X5rqBQ6
lLarMKTYs4gYBPv0IAVJTp5C/MmNEYx/t+XVHsLbrVAirDzciUxTUPPny0t29TLdtoo4QdiU339P
sHpk2KrUYjzFf14VlnSbiMFjVyKyhIeo+Yd/FY3Lhldh6FmNKVALf6aEhNKjC55+N8TGavezP+oX
v+aWhrG5kzGYbhtEszIro+4t3zHUPsDsdomdUys6bJHqinmbShAtsysM6/YJxO0GtpefFKNNQTJK
pQHJwZSEEjl4E7Chsq6b773rlHl9lSH8gVBVu9OT/YygfTPuDcFKtohfUfzMXST6VUhFaxXjszEs
0sy8B5/xqFm7L6+WKu9ezqZ7VyfwAvPU+S128rvkBB/pr/paivwiaWGhIlcKwNIPsqEZA9gmWRfm
qPzMjqs5/Jt9cO5BYTOvCMS8MxKKQ5DM6uvONtRRbbSk2l4gD5yj4ixNptqGH98KPyU2YhfnybQb
Dbf07LWDyPSJy/YD6xcugETzC1hws4+Eq/pDTH9jl1FTZxKmlF8exoz1XGcPe8oUWpnqya/0wRyu
uNaGtic0o/xZUL7sV+a4tf+cPqSWUZNui3SDFa4qqmQIqvbX4lXISpOno6FI9v/zj3L5K9IvFiRL
LgK2BrxdmZPyqkzye/Y40BDGc9O+xv/P36tE9/cmiWChqPg1P7ioeUVBzs9NvJADhIK1F7l82AyZ
lygZpCXHA4Qd0D3y6X6NCu8oGJwvbWbjGTDSmUppMp8pRTJOwWGVZr2MUdhtjQRBLeaJcYd+/iWN
lSX8WmMWqIWUqHCY80Fwf2IfViodJRlBIMysZ5QH2LiYQVqTWQCQN3CCLZQfLV1SSvZrNXGMExbe
WkAENlMF4ZDnoMPRKxZYYxCJXTC5epq7H63hzy3qG0FKcHhzcpFFLLOQfJN41cqfxd07dr02divD
AOvAHOs19IJx/7Kjkj73iKpfb4G/AXP13nXJnDrsw4cXgrRTg9T80qG8q+cjc/tHSVi+biigOMIs
5Zo45uFPwfH5iqrtru8tdrdxhljQU3nKuuS+wZp3wy5yTufG4T6wK8cvNCkDCXXvS7u99qXXo083
IoA3wQTTPeMDM/A9arYGWaAreqh7Ka8Z+bCfjNc5cr/w40FZgRF1q06d4d2Hta0BhbYn+KwBNJiX
i0bB7V0ww7JPzfN7U4JnOf3MAGMosaw96Y+lgPWY/9KFVXNKrIf+826Xa00ryAIJpcTJkEg8zAg1
vUVO3fAXmMqTzUYBi2HD7rheWQz7TX02mvdB5DPi72wCzVAGb+qHHqIWdsn9baKVts+JMjsEWPJF
Ts4dY1iX5KtR4wNddelm+SnZtk0iKhprxWZ1sH1SC+HFlsYn/z648qaoUIXyKZMaTio66xTCFDoh
hDZD+jyfPfML78/qAPH9u95h6JTqcMEbfleMBsE8+ZnNbvV3NPl6TAGfKDUMNf4T7jCIft+JI8QQ
fc79p9cIM7HVfKI+4dwQtZrYqGZhkIzNJqIdpBuso0y3d6GaIzPtOYbjkRZubaDwymTA9aqGr1Xo
WSfmpdMCxZqxbypRPYPtM36WKWdIW3bMMWw15P3CWTKU9LeOQcNUtn0ynXSkXnqoxxmT8WyIuTIQ
cn7Wn6hvRynNVuJN0QjCnNDqDx4isB3B+zeYq8WLle1QrVflIHgRlmIJh6JzqanTuXCET1nWuEZO
r2Kod+wXa3Y+srElJE6QKElXaHRv0meg+e23mBR/QdZ882lyJBUkCXntzo3OHsZv09pV6UQS/H7V
WwIuaR4NZrzhp1YmbOBzVJuFKQpWUhaa1WRS4kDMjZm9ph4sJqpOJnxQEkFUTv/rFzY+Xhc3B3cV
WJHuTr/9c66Y3oFbMUDgk1UXC+rkLcoqijCdUSZuhTkL+ZCn7Cw9cxyW/1ncGDV/MwCJzIQJCBe7
e/05y6iI3AOotcc1J9KysaJ83iflE4H8/dhhNUiOLMCDwq9QdteD5wva4sEF6PvjpplxN6Xapyj2
r3cPxML9FJWWFl0f8k3ZADKrruxulCGxZBVcEovyKDzSyzq0sD0oo5KNC6Mkj9EbTAzpT1ao3BgP
7xOZCjA4n2RCDPeFSDWoGdjV/r1xHNfe9TBrgIqS8spXYT4wGdKNjb5eTxLnfiNtLqFbC7POnUeu
YI3IvJkXci7Hw+iox7gNPILK9AouxpA5PJKXHInimJpE0VOECv3wRiaJFPE9WoVXqFTR3F2q8clp
HLvSArjYwa8/gqMm/CB41QvrvilemGr5l4ohsMn2hmP27zItgu6ysSzjheq8tTZoFvQKQA3r9LTu
e7ZA6fjKWjePQ/LUWJR34JANRan7xGa4mJGAmSfzgkMVRY5Y3QC2iAweZh5AMvMVZy3USmWtxJKL
SWUHK4vDaOZbrDiBDJTPzlUDnjh8SxXIzet00EUY7xMNFcDG4q/ICpAXhPLYGBU60ufCWvER9ZwQ
oY0TkUBOOQRhEUdugo7WMmbB/ZUy4/SkS3k69CVoeulVp3eQyLRa49ApruPuAJuQ5/gpEl1r6QBu
cP3YGkW2YB7IBPKyvtvYipHH4kx/cN5S6x7TArRhMwkKxHnLddiCRcPKL5aO2UaHI6YAFIQEcwvT
d8kTYcGVYF433EH3+vH+YTiYXPHi9b4vMHpxbKFRhzsw/hwCFIFphaMEebaPZ6IjPOWd81bE5x1F
1IekqB+3U6WFQie/S5DwsJ8Z00tI+sHCxDkxofgmH7nCCP7szRKLcD3Ggwmudfpe+fhNdWgfgKJv
WaYqztjBXXdyvILV5qoTonhqR7fKFEK8TfgB1e41CW8iwiieV65rv9F7g6QmaRX6Qd7JytyOMaMp
H7uhwBGEuqpYqcE+0pksSUh1LJyZ/yIoMbEYpTYQw8iJC/+jvbw8pYcEC3IhWHlTtTwE8WGzijBV
Ra6M7EE7C6mwQyXCSS1JPw7W9MNOwqrhpukvE7nDE2Z5YxXwW9CVuxIm0pP2gZTteEE8rb78pkhH
sygHhKFXFjaPJkoGulxpkvh+ud1XnMSWsBCOPvO0wrqzcVXeairYMXvHbooNqlZgCj4NmieVioWb
XpOJ0uVczgEO4cnh3SiPvMMdtzTKQBvk1WmrVOBAN4uPVcIVhGe44ZBfs+7wr6mSZxYD5W0GqeQB
HiXhA9dJaqtPmP3WTTSv4FAGLvsQE4cVtPLm4BR2//H7qc8VS8LyPR10T0yCXcwERIEzF8QIOB3z
7SvRkg0sV9KMj8CA5vIp1gho1MNKaviqs9u2NRs4QwlDgsJGzMNYpER8X8wVvBIeAOlSTVXcTjv8
FzrZSZ4tPK6Fix0zINzn3If52XIKHtSNLwsEdqKiDCABfbCSNQueDbn0MmN3dhXOwGdfsfr9fcHV
Z9YVIF69iFTlHZA2mCp4eYBDXBj5tUAE0G5GpOenuqunNObLtkuSfmAwzrsAEjb16qLTRlNsgUeo
vTHrRGj5EnjZsHzJ48iXHln598OcmVaa3AAYhPfZhqZKF24VPaTaPhBai9UFbrapU9YF57R0DlDD
Yz/LYBuiN7C4JCHk0WESERIWRanY3BBJxOGUM44YTuQGq4fTfpHhH5je//Th6OzNbaYiC7VEVtzL
H/6qIxx/5YUmve8pwG7ruaWRTQy67VVgiE8v20tDXI13zB+gUbXc7fqtxCj+tkcAgj0l9I/bnNQ+
4L22Dfqt3C1dOfHBQgC9bChyxExs0dz+O3EpOKSIdB+1foXamhEzGO5NAjxKFRH4KOZ98kwA3uwO
wFcgYKLBzsQ4HQaRDJUPO/VPqsYVKglq1pEmyeOdHZVShP7OPvpjl3uh6tlp/n+1OoN0L4IKJ/qA
BHLDcIRV/SYuc4HM5xkfYaHuYrhTrNqQAAkKq6h/C/ul4q9d6A1fDHCmOMf5y9R2uCBi5ko9n/O4
Ce65jlAhd0zUnjXgUe1QmMISTS66f21e3nOsqE42mpmL+ErTLg6jkea6Ib/En29RNYbQLI3SRUIE
xU87XNnzS0u7nI4IJJfv6OOBGmj5uEwpTwqNrLQJVnSPnBMOpRo8PADhM6tESam0OoV/ioYSG9qo
UncpOBMQoldC5Y7/bO/VG/7q5GagTX3p3oIdDGUkBwcMUR7zl16E6aIX2jaUgVI7MwbLDqI2FFsD
/3CapLML8CBmJGdQpLteIPKONU3AZzvgujyAAkeSb35rHF1LJO2xkC9x2fHmZrRJyk8DsGD07Eak
xJCSJ1p7nPAlgL6NafJzecS2n2zPhMD0i25f5JmlwdNvsvEj5Hz4SA0AKsuhwSwUwZdHlraJwaPh
6aTUHcWhPRM2CHKAD+vx8sqmWoZROsbN+5reB/qU05P+OvZyBmWI3gksocishI7FQbybRWGmT2ll
VNQL/SgedEvAos7594qnDNPByv5ew5AF5On1PK+h8cz5eiFmWPn4U3PL+GcSpAozXgzMQSI4ELS4
kQpYXpMWMuoBfECg0/W1Xa4FwBtcAkXUaqlFfVsHtQgcxFLjYmkxtbsdGfLroxJQz683LonqYg4V
Y3lSFOhqncw95MHJqIrAVvQ1s/jXaqADXrlfXfSfVelk20Ium2fl/aUq3VY0SCD4J6O+lUxbYb2b
jS99sWM7Dr+K2vGo0ewmUGc1Ej2USAefz2rYo4nzo2kQjBpqilm5BsStR0hCA3+xtD+zYt68qPbY
uPf0Sb09T5cpcrqpejUc98JHLMd7XPxSPZzcErgjLb853CoPqzzDR+aOxEysJA8VJa3AKhvpGKUr
PtAHgj5OaeKFlF/pZk8bFaecZIQ+x42M7Pa9MKoLbtuIvt5ygR3fIPujMlFTtH4d53dIMdEbOzpW
9udV4nmPUCW6wjErP3Q4BGVDWivuBb0oubRCQbVP1I1Bg1Fqut6C/y1ygqCmLAz4r2irt79bGLmm
KogagTBiPv0oU1HfAGy5O26XEtiq0DHTmsMY+jsBDnK8ht0gDhY5Nnyo7PZnCYBTt5+yZNoD8dbM
VB/Rpdmfb8T0oTkLd+sdiHvT6bO+lOm1JzWLTEj7gqeWneB3foeFN7SVwjORTr1fWACqxq6HZ9w0
vxWusjQUNKuRc+ye5edPcNWKnR7pnJbW8Q8k19ktRkjBNDYSl0OWtz1BFYa6ZTXFaZhdJ98PDD7U
mupXBnTcP5QI+xewaynuzCmprIlx0s/tZZSJAFp7BScloaXDOdBzsGteBzU6xuxT6NTKMPP15/20
kWH1cC9Mcoq0hlSqnP4qcopJzSyRx4ABttF3x/Dzdo2mQbL6DiEncE7nUaVJAKsZ/jA/UBGhiX+7
UvEDZ8KbTYZUFlhApH/gZ+qOqU2IBvpj7h/aKuwsjf1J5elmbDfc5YUUNdn/PgeV4O+7J19bCLJk
skjmzkiqGpsuE1zB/PCNsDetLwOXYxKf0XTmJV+jdj5KevnIuzkerYmP4UXJMoi5V+WWlGAOEmX6
cc2BeR7RLAUOjmaJiy1RztOicayFQQFhO0YNe0cXZYEMDOfJq7BLhKednLBtoWu6Y1FKrx5ERTY3
8ZTQcRzVDrZaIolTyMO+i/7IqbvdApKotwxJjs1hGM2hmpaPzVdg8AM7zqonUMrz5R5hH1upemqH
U1SBbuhMz5mzAWI0az/3u9pf75izZ48AqzsjSYlFIemNY/Do9Dl/wuwe1lUNq7gzdd1SQcUK27mH
8Pc10KfRxbtxLUwtJaXWuKiaPGVXeuxCtRSFq7T+N2UItqwL/wOdpmJxMuCCvAldq19MRqVaxC3c
mDhsUEhyOGS/rt0qzhS6CVDJsThp2Br72zTST34uNS+Tcjwo/nPJWI7Y3dL2rpkhhCjPD1/d9XUS
bW52FVFcJFugLmwbwztk2oaaFVQ8KOxBoAeJJOObppjGnziV7nSBXEM6b5RuCvCX+LL8jd4bEUB3
XVOrcklAikuEf0wVdH6g3H25waK5jNWRb4O/Zw3r2Wrr7jtXytmvFHxI2LwJ+a45Buubel5C4Ygx
XiwQT+YCfdXK8aUNN+acKPqZHHoALAgGcEIUCbo7KGoIkTxNY/eKJHXe9Fm+EsGRA2/g95WVcv+8
0OCUd+bF1ngEhlph0UOn3b+uzDiVNbscPtOTblma8FYYLA9K9Z37r+wB4ZbHUHIypVdb7cu0Ma5z
VZC/ZQ7nPrSlx0JSrDkz0aPMGPiVivaKDXynMPT6zXiYl1XPaX/curC23Z8Gjeo1efgNSG2PEoiS
pac/vjS1vvJmC6vHVwY7ZGLsGBj0Jzgq/rQ7G9mBSCXpXzt7KqE1Q2CG+y2qupqM0qHHqHuY+wyR
RSBkwOZ0SkBBn3sJKVK6zHUiuxin55I+0RJaJRJdafMmNdmb2MHRPIL7cgLwreSWXzsWr146TlrL
7MdEfkL1Knxzipd8BXpmfd1vaJ3YtbaAp8823YkAjy/LlixVMO8Yg41+DgIYr54mflfXPTi8hNgb
9PUaLg/CtJ2xC6KGeZwnFnz81dRlp6paJJtnba3VY5TlZxZiVdBE4A/qWJLYlZziMHSWsN0dZgU5
De1gPn3/Q+crfp3Iy4VglvvcIlm8d0TSxA1bnEL+w/LOCWn8K+NducSZwya+TIhPioyMu7nchiKf
aw5kUc5UfImXNfmMRgtiSGyww8wN5THNB6pAZpQC4G8W6EcSsUZDv96Ml8ldQ7q8LtVr2gL+YAC5
ivxVJkLCCYBzbS2utiPwEKuqmxLmpy91+1eDr86xu5KAQ4/6EJDT2pjbobSAeT7IubmAfcKmn7sr
7foZaeNYxDArCoHjEJweUG/HG7dLkTFCE4e6wpWRZVe3mm23i0yURM3K/juTxIntjwTsyyMsDstE
O+otoHpNjkDg+w3hpaqkTkn77YYK/Cf5ROtygXWSQta46hlJVKgJpfMJgV66YkM7WsqDue2iZvIK
1nX8KP9oPZOY+gfT4a1kn6k48O+EH8+r+mWgnI5mR0L2y7MGLNyxg3aKhh0QeFEQJnPNci5M4vNs
RlzJNHfdp51TqCVA8jxY/wgYsRDQYLZTw1IOxoYuC/8427GXwUKymArN6fxLAN9+Ej9/zLTF7KZE
n9DGu5ehHuw4fu2VS2djHrkM4Csgz2pPGChTKtpbPY9YcbmFHN8YAtRctSR1R/5aHwVmRgn1llhi
h3vI9BM0m0kk5I4ePP1Y7uQjS/pySlGTvgeXgdwrnpw8C/F4kgjONqPi85COjVPpZhw+gYr0oi09
0tQE5AJXet18I72OWmiGjp5PZoXHtT6lPR7GbSCY6H3eiiBUiAm1eg3yXjt3I8hQ5m4/eeRIVqKc
CiPo+HFSRxpUGGURurZv2U2U/oyhJORS7+cPaHsN67Nk9acsPlDNppBuvwSTCJEnbAZsD1rJyPiP
GQ3uvQNSIA/YyzN4pqsfqGbrOPN/M5jszxrAtpTX39H4/2abdJOn9QYtE3P7fMnuz+5RJVJfxQWs
v/RvqPm9JWY7iRb8sqdQSDShu1IShQ2vIChVI7NJqFqElWiNn1F39kHeragDfGGwOdfZkmxuLTO7
PX5Uwdpof3gxJPSE2upLONTPAy0C1fOglHNJqXaX0R5f1T9V4Q53UeVL/i/LqyoRikmMISylSdEt
4u9vG+MTEdskvrcfQGnJY5BENgUw8YcIow0x47Mucxp+v1Qorco8ssy/slDkDUwry8Xq+Dt0fgv0
6KleuRHBeS9DRy2zBel/SygP48f6bfdKw9ffnIwH6K6Wpz4xoge09+Vw16fl18sSJYVq9/Rplo7J
AOv4FFxNo2wy5qNIGnP0FzZppqpabNeykvskuWne8qbzqPF8pAERF2HQQrvW5hvob4DGdCDCCV8w
ElkwucZe+VT+nJBFZsLmdq2xzJ9LD8AFigPsN2mM4AmLSSXbE75GhbWmzphDMG/AgsmNzJfenpqw
mWsQNX2rwspajodwR4hzPg8JONa2sH0cbORLGIrOhIUniYw769L9gFhAeMrX+57vYVucQuyReYQf
qrwmv9RZNaz1D+6/cZjqbYVXsauIQCuwTaMK5VOHW+gd5u3xf+pAK1lzM/l/Jl9DqF++RtGWCtnZ
ne6pK3DjlzICLZFsQx3HsAZoL6uFttXnMbBxBwqq9mYg7pSHKJtV8513fSf/Zuj/ZrdK1gQ9Mphg
oLzXqniWs1JY6roI+ZYN0vAAGgUgPEGJfxi3XhWeyHC0z7uBemn1+bCLH4g0uHW2fTrBkMTEMopr
l590AeCeuDgN6Spr+A9ZMQjZakkaktEPFGw6z9iXa9YrQtF6MAIVSwR6hzCubbV1cL9+5338ThUA
nlBWipzlpAEPppHmjkQ8Pb5Kdb4lYqBPiOpa5JMTOd8KpuD4sii+HHzACM2rcBBExzLIOdRqQoIB
SqOoYbACN0HKECMFXqClSKd5WrodeWVm8a8aDZ3tKiiBYQkC6Xv77siEePwm34WXDU3qjiS8JAkN
CmG2V9gBh69piNi52KHlHSa4W2/AfJXVwBUuZrn98fpkPdLqMcW5yQnBzg0iDbzZaHB3qpRV9gbI
bIGfV34SbyF6c5HynAbb13eJCy4GdywU/aNxwJ7hWPQx2+8ss2ouaTICpqcmeOlBOUPaIeWeKl05
T4LXZTmrTP+SW95MgPSce+AF9DWHqWRTtvgJT7kFK+wx5ME7s8lZop8uRE7CVZd6tmKdGEOV1pSp
2hBtD2KhcrQwJmOAfZuUuY6JGdDRtC7RcTQJXkPO1Zkt5D4qFjpRztxvww0DGskZ+tiLzUrR5KDz
aM/Rkaoc9ISRxhaGs23b4tOpdB4SNixwTO40DR6lew6a4f8rIbGBmpxdOBnv8eA8478ksCPvBdlt
v91Nul9QnROD4aifffovZKX+cHRgZlrRRmMEh5s8Icpe8tgpcVyDIv7ZVIRxaxg7/FvapbQqMcPl
2+ph0UILdEREyfEgokCa9xjwRucLPRiOq6XuAy4sMxVNb6EqkYIoX0BcjnDUSDJZpz4ImSjqbdz2
Vk6F9qf6rpnvSrP+J99JUuBecVrHF2Z1ycVrB58/z9I1zt5Q7vcUK9Xqmbu5mXMVnKdm41KywIZa
lF/JJ+469gpKV5aR/D9EpgBNdmRebefgJM4iYJVMe9fcb8DDZbS9zqkMtjQgVJfHPuS4l1azjvpE
wTr1Ui3hUdOYT9GGCtojJ4HZhjZ3H5yjfs9DT8wQSmfItFxPi+hl9HY1ei/0jS5kCU+D3cjATXiM
jg5hcZVQ6tIMVsa8iePszs8VBJ1Tln+zvUjO0L80qitWFsC7CkaX2AXW1lFUs+cWo+d+tbNgZZGG
PkDNC2RRm4oXuWKvA4G80QpMCWq4d53o5GdmoFrBFUw/TiPILRY0Iq5FulSbFIyGefHGXFP9aYxs
PE+ea9vUWy9/wN8HvqzYfMcFK++VmvxHVK4fKk9yLRIujAqMgnKisNNAUwPOBJ5VdKLaQDuFUZhq
Lc2Yjor0QUHb8JsE+jORiLQjadgCOc7yxSm5P5G2d2ia8gQj+B2FHop2oTtt73nz5Vkq5w9Z+O5R
bzvfA1jMAIreh3kuvljRh/pzG+fTgfRtPRfETTG/KEEdnoj9gDyiM0kfBAcn3HS92UavQ3hDEDBn
IfpHk3O+aXbpt8Omqw/L+ck/uiC/4oaa2ICwfw0os97MsO1TakDX7X7CJjhW4mReZ+S0bl3hgibA
hs8ism4FOsXJqmOuCbeZTrRj9O38MRXJZVLH0YSy0Ares/Aq4ffGc5YEpDJqLDf87R/eTot4/xNC
FISHwdiseSNWLe2ev+10Zj2YulKoCPtcG2z23oqtwNcQ239bZu9Juvs+WmeWfE9UuHNjI1RlqnY5
dD9vI+h5HvpxF5C1opEt1trBBT8Zopk2NmydRLPPeVNjWiC5mg/Kmk6bxdoHKMnriHWgbszo8u1S
luVi8kyDw5/15oBCaAJ6c2qBKj17ZV9IhCd5qG9B7vFMvn8EO4/psslan+36GApf9LlBZk+iQgSt
zTOHOX8b2J30jO8YId3F2UoOVLW7rnm1MGZlo9rrePqHzMFgG47ulMG07UTWfJpM3fHFBOmzUVNk
Rv4FVUSjUlMg62rnuU5uQDEWzx/fDB1xf5yPIayfwJwXUuaY9YSHtrQhnll86erxB+BLgwWL0F+U
5XdnPHQrf21pJFGtsa1sIJ4J8UWIAF/qJp9VFNTnVTe9pmyOigifkXc2YPH9cWC0D9Ue6sr5x0/8
X/u4W8xv0Sl+5WfzyhLQOInmp6RNzqOXeCfzdqYrz1NR+LzQ3w6DnlO9NOdK/TGeWtLdmpuU+fcO
ypLnyrIZqhElrHvY0yfqNyNqatKBGPSzgnl8RHxYv4vikDqipus2C835iy1drZJvunDJceWb2xg4
bX3bUc2r1TzJRermqJgj4og0BABRNwrnW0Ej0xB9vPVTrjVk8Z5Soys/0BUHF64F3mz70FTOjK0O
p2RiH4MzqUjKgxQG9wPFdwzn00fAL84C/KYcTKRnM7jnGfRNOcAVNzecLwJH/kFEyVCrjY20MdH8
QJlgjqYSvpx0STZphcLI340qMoIaUde+FbO0u4F5AZGHjTq8vFJbyjIsCSJEdoWhM7zVNcjuliRq
JqE3DtTYOeMkHw+uLMt3rvUEZD5SHArHRp2hp9+JiH+jSuXL8gT/swzt6VNtQzcAirawUcWizCid
e4CZknJZ2OB3MUuLxgH7y5+FroNVo439e16CH1si16SarW/5X0AmRwhRBgtlxDa0wt8m+kDUUbHF
idLkIwdN/V6MOcfmafbbNxAsCc8+a4GyYQi8DFq93YuhE0+0qT8Ku8eHHeVlp8IYJxaQJ66L98J0
/KU2st1k6qUp7LkB98Wcg/05gUNX/U8brsfYaNzvZQNDwY2QRU5FKeylqY6mAq5cGwbXQM8hYTfY
Txjw6y1hxyy9XqnNi1GR1cebWjGYt66ZbcNQCIHgZt9EZWFQR2f6hnr7ZTHs/Jp62L33LhPEpCsv
CSFDCo1etvX/YYkYwadNDkBr1vTshHUzgqJ7Z3QD3dxxL5jsoTdjijgzmN/bnLoN3OFzlQ0PqutR
MiKuyg2dSmm1YBezNlV57lRSXrpkl/oT6ctWR7kGcmq6hDHRoV9SEq06AP0+LA6LKleR1Tk2McIg
m2aosqS0tjlI8vF+5wNGigKTMH33x8aB4SobRULtklMWHQkenu0F1VptxfNRYsU/O5ACmykhTiG/
o9nxbg/1cp4zX7SnsoVrEGiF2szzmd0MgTThqgmOSIFPnFhV36PuQWQ2k8HxRJR27MrHnb1lNMXl
+k4HKGUyRuA4xtWe0siZfvXaYqLgaJrVqTAYKlCKR5MdPn8YlWWyWk2ovWPEOYkdGwuF169YLkxy
1XRjSqr3JkBQYhgqKj14EinO4gff7evno34JzNgf1eq2FXdwDAru5mjDLtillMX4RyXx1btUeu9K
eiAQKX/sZqEI3VkP+/9tvm234VUQ7Czvh19zdCFMxyPuyCLkxdGcNB/Q85LQBs+3OHFIhmAteU2o
Bsh+vXVREk/HP95Wy+UwHlvlCrc27fbgogi3iIQUIGlx/+xl0r69q1/bmWqTW3L678GeFS+xhuBL
7oE0AlkwQ9eI1lM/T/PPyqstPHunwgKcbrvDa04UZX9Mf+aA2QSS13lzPCkRpSWxeau4hVojsGEm
alE5rzWReOJ79ISCfYZCiYjj2qnDi3EQukhngklEae5Y1EsKNMQysvGdmYvfdPdRb7DcpFKEy03w
9efo5hYUrxcYaUZH+OnjiUyXDm6Kulskfz+ZX/VfxrFyUEEUcBqcZV/h33LaPv8ZFlZg5l09h4vz
ITiMAckHIo5I2b2Mol3wN4HJuL1Yi503lQEln9+nPtt+Qwd8lc+ndXEIoj1rwZa/1KLRHu6pIF2a
R23G+53ucf4V+y1aj0fLBj3kiSTAgu5UelrOYTh/tb83dQgTK9iBG6m/PaWcimQBfG3aXeAdY00Y
jI14Ght6g7vbUXWVCDhiC8jp0ytYt8mxX2WlQH/I+gjlCrdEPWLUjF+cznRZrR7ofknOKuOLICZ2
K5Fr6a74n9mdhGyNu3Z2/n8On9NdSRVoI1JW7OOkugRw4JMEVu6vPg3ehNy9X60CvxUDBxH6OtXx
EMYqdDUyNw3XNprfl7BC1/19yuGIJElAvndUvctS4DcKltI4Wr9viEKSWJ1h0enPAGrdMSeU/5sa
gfh31UHOcaElLrXij7FrsMkEYZl0c3JlvEJs543RYcky4qLq/T5+5vkA4KDVAtg1CUoM/9f6/Le+
KNCjHxg2Dv1OFQBtuwSYEowCOclgrX1GY7PArMo+P2eCCruYdDhvcPKaa51b4SCCrwl5neCIsEEO
2l1bzgcPaIVGemEi8KNRqtpj5UakPRvrtqnuBOraUfvMpEmnTAkmgvmIGJ9bQFBoMd0ezbdBrTvW
orNcG+gpFU1i9yrEKP501NvsUGDMWDBtqNW4+1ydqq/0U6fLNvMsl4GsKRwFJnnig2DcU36VUZtu
d6eJIszrPtawLV9/m9sNWUcMt2XZgbiNQ1IFfJeSQ4+AkIse7GYVEOs/tlBnbJahFfTyXf5AwzOD
7m/fAUsZm+WslXudyqR/ZVzoiOu0KHSc/0Fg+DQqT3RX18721p3c5LBcgY5MsnJk4sAzgC2EPp2a
MrX7Yitmnw4gWy3URdNmXZDzMYr9xqYCb0Qe9mqUgEZhTfA3IOiDbnxCeslEE9XMr5QY/hyFRIQH
VD55n3V2mf3sBYB2s6BhRUE+fIfgoEpSzs1ymI73kdyQEoESJ1tWhTnE06Jd9ANAwZbpXgb3FcJg
eqJwV7vJJVsNH1KgbfsDU4DEuZ9oYeYDh9U5vEjB3nV/69x5l2AZVn1Q37cpeloVVn2oyWj59nSQ
oftoZWLG+LD7IGf1l+STqUXBobGKI96JqqgcllmAqhqz9gU8gTIi2mOdebQvL21EHjh2gnNhCGnt
3TXMlfsFyAil3x2fuNgXyJjVNLNvZ4fCzG8ahhWkYzyiAnF87+BBAMC/73SrROgo909Nt5ZoBSGK
8gM+yVvb2/5AYcunb4PPE5XThlTeRuYu1J64ez/J2fp/HJKk1bbnRaK9TEGKDeYoJI4kWxtzA/AI
dKtsXwPUAvgXmwl2b0oceVjvRZ9bWk+nQshtS9bTei2n1fQxPXsNOZT8A9iIRc5DsG1RL+s13B4U
N8KpoRHxvxnmqc7xleYqCidYjkHsLLqhyAVoJ9ll6ZDyRmeQ0o2R1EBH2t0QPepEAP/imVODzCkM
iyf3d2VamVLEw/PU2zkm7y2w4S78imPDd0jCwPqELCNYPTSaM5W9/vI1sbL1SmPsBEIBVyaJOi/b
5fGGTXCQyLrblPUTgcxwgOxzrZHB44SiM9UMDl7QBgOpbS5zM1TfZlwr/mX21J/1rScdO72NBV8N
fKVm2oFTzmGzsAC92Zf2wBSK0Z42hTGz6cN5UwqEdI/sxy1ExN5tt+V1kr2RVEqm3NRWctnnSBYS
tjO4bKaKXcNU4V14KeiZMM7HHAdiqr+rEPa1cn8lG+8MVCatWen70OWjbcdcx/4WjnY+tX18gP10
/qwQvtRic4GXePJ245TeeGaSZbHoMcFa2bRKkYcp9ZV8US/O9UlvCT4Qw4TB3HrmVkvn0dan+QkM
A3FbEvE1fcoNiBbwDYQ02jr9UbPB61mHsLGnIyxQECCHfoR9U95ypRqQU0NRt59POlBzHcwwhWz6
PTPQ9GY+aO9ogT88tnivFd6Pw7VTZsie2qWzQguKh0j2lvKWZ0orqb81/WYNsoPUUbFYhjkhnz0q
A+uPN8hLLcrZ8aFr7yqbuzkRG0j/wrZgFwWsmSdAlmqJA8NvKFfy+ePoPU6/9HuVH+7KQZ2BTbnW
LfZDIqVxSpusChBt5YsIiRyXw9W1t+MJYIRfd5yhmRr/5XP8ETB2ihQVkYqKBjPpHbPVcXtcLY+d
U7HiQdTnTBajOZfn7c2deA4h1UCHaog98yhQO/qZaCxjFViEMhhLztarPBijVKi+MsicQ3zJw6ZG
W2OmLPlBdIrlmVDTM9l+ksaGFIzuHPuCNFvrt7LucWRIDrio5tzEIXk7S594EYjq/OTnkXjdlAT2
DB5NQioEo16GmESM/cquyuo42QlAK9nIF5RTN2hYTlyPGOnUn/lKQteDF5yckV5qqxqPspUQCzwB
olNK/xVDIROL13z1r4lbFrG2x1Of/jN66cWOX66lw+7HaEahb6Op3/BiTDpzRvr2xjCofzsf8pgO
TTniR+3YTaCqDvpjRO3O8hvWJLhQiKuSzVbUIhCQ2yb+KSeS0zUsNHKbKwDBwqhvafIX4sz6ETw1
79/2eTXlwJFX+QcCfpGLLLc5j930T5Oyb395OxdZGc4PP+Nu7/3u3BPtVPwYK6qE6hykks5hPl4Z
KTlHA3SnqzzSdSrmo50qh4weu2TSCWPFX3uA4KX0g19e1x9FD0lsKqufgSJI//RBx7s1BjMHvw7E
Bhb5RIDNq9epu5chD7MekQEkmUmf1yXJIFuNacdfmsqn0k0GBnN/DEq+Gx1zgMD8L8twG0AkbZ4T
9nSvEIHLRTHIz0zf8DVaZmb1tOKEXjZ19FjecxIktirmssT9VOcIIcsHWJ8VSbbmLUCZltEawTql
GVVnQRWqf75cRgY5KBfQri+Av2kFnEKNQ0Etpn96RkrV19Xg7hXjdTM4liv1sJDSPPOw/yXFg7OT
HpGuk60Fwwi4aO7lHbpiymBIceLmo36+H6jK6Z+kuneRa5HTg4fYNdju2odsv2B1bqXELtT3K1RH
2SRmi9+MvEQpEMf3w/J/smTk9FjcxIX4NrRRCdGZGS1UfKUrlZEaSeny8J772j837Vu2vn6jzwLK
kjeS0x/yegHSFRhGa9g8jexV64mklV3iyvTj/w5HKzWuSwKsG/4Lssd56P3D3xXYv+AifJ2qSvAQ
qMTjeQ3CcBRbvyFeRQiQrfGiDkNcIXovg6QGxX6/VBr7qKE7lW+AlcxgzwC59AiZbgZvcETfGOZc
vkLfxzg5oMSezN6ceSOC4kCapiuSjkWXG/UIkd19mc+1jJCQtQvJlM0PGz6TUk7FdQyAhzsAYw1c
/ANFB89JT2YcrH7xBMpKRA5abW0DvVzIR9+F+bjAB2hiLalSl9aqKwq4ruD6PxCgN+i1wDWQxxs5
hcMlAC6xFK40e5xIPNvM/A3Vahdd5cVynowfN6yTjFJQVkGN7GMVatHP8xObl4nLFvidnzt4HApw
7JKnkdkcr6lzFJknhlfwBTBUjM6/hmtkDCo7cyP3sfrUtWUUd8UucBkuDfZlVvzuQFSbKqmvh1PH
IjYyijT4sPSNiFr4FbCgOPXWpyVYbJNgQPlmgndK9wPysmOX59bNq6dZwSwGR7T4zx6pQz+uIyRU
e+6dCjkUsaj0Jo7xCwoJM2ZDLYcfNsd3WyZluIZ2AOrDaqaQB4qLajBLetveRlGL8y6QlWZj8Ye6
K3UbNBBRwZCqfiFKN9rSKpwVQ3hCLhNtCXTkeGPGtPAWBTJr4n/pkq437S+a7sb2vDfcqU3S9xI4
fTQ7pl8Rfxkjua2FPs5AtfF0yJR+jS8mSueNWRv/2ZfpMtQrsxoydhos/cXdc6TcwxQzaYkeFhb0
G4Z7q1sFTIQ2AHoLioFIVlbB68aje9X6vWLxOLC4zUJ3YsskGbCCPlPRWGTXvlM2j3QT5Fy4pTTL
DVlx84jt1kLaZouORZFh1jVUoIyxlWO5LRBSpQXAd+rylklqCo7j3L6SCRqOptGvz0aBL//ePzJU
XYPC805MJMv7StPU/0cL3Q4hXDyuhh2lCqVxCixqIK3zXJgOjpEr1xJCgqyYsxcDdIW2fl/zCdUr
GXdGzMOBaIVDTqYaa0dJ4VpslDkn+aruTPB4ZESyDX1TSaKpxW7c20GvDIufFRRCsmfx5Go271Tr
WI3DQWtMfBanHubDjX9uEoxArloKHsWnhGGlpVHiJlrd4Jdezt4Ph75mNJbCgT/Q5MI2fcVW4FOp
SzLI9b67QikzrE5Y6FYh2q2FzdJucMTOD/spMEs1F9wAq+dBraiJMV0UsCI8PgDnvZLRQK+1tIRA
Jlqd4rcQJj9MLofG6h8Bteoko+Ylf7xq6wOwSjTAHxR4htGZjaInIOoRaEHIr+h+3gQvwU1mY8yP
W1v2D/W4Db+ZCgF2erC/O6Zw3lCHyoPPJ71Mgv1ySx59GHbUEnFCtsjxSgry/0VF7jnA0YeDYQ+7
hXP1LgvYNMHT3IjI91vPt27Jbdqq9d4vBL7BPSA1BN2YDi21ehc0aDUlIleQoYHF9v1ALnXXYMqY
1Tdx68V7VvA+XuZV+009pKj448dN2aLI9/dwzP8YWJcKu85kdRn4XI7iQ9NjDcajfmcazChUZhi+
rUor+gaUFjdk8G3ZssR8U6oRARYOAnXQM5vBuo5aKM1Tyuw5PKDz5Fj3dXJLKnAhbwC710vxbBmk
XRhn8+n0EKOzpiHPPTs7bhg9EZ2ePznXaGRJh2RG0iAq49AFaxye8OXYLla3D7cblsSJCyXUE0r8
GP/e+MEVN94a64vD7Xlgo1s998nbtpkXm2OheUrYivQFD1/A+KoG3zbAkmhbsfAUkny5poW+FDI6
yJR+REebkejwzin8wPdBPWjSFZdbh1itWIyk83ugcYLDIW4R82buHe1XniO9syrSCIdUjkMh2Irm
ZBc8zNFUAHAftp07w/wudLwNOJGMzMl9u5FLxo4uKW6IIIQ8AVe2HfRQAeo6XWwJvP1QU6yxVgEI
Xx4llRwbqt4o3USzzFZYg/tz8i2jmx/MgQgo1tievz6EyPYD5W/HaOGmTtC1XiDtaTf/YWC0Qijd
A0NS+48K8/lp6HutUmedIqI85KULYsaJAjumA2w0Zgykice8Yqwmj2LuBfzLzOrHqbjBr/miKKDi
+7CYY/yLyEVCs4WYQ0Yw1MFTNR8vSxx375PKs9kkD60sn2dU3XItTIT0O6xxFqW4jS/rxRLIg9E9
e7XpLlnNsuOOliYAOwpwXc4joPCktng083Gl/VtXMVUCEN9/gTpepq4qJwAX/AaKDPnXFwaKKeyC
+yh/sDzh2UfBpJMxZ5FMuzj4RxNQHqRkeMzvcHDUO0JjjnAZsz0T3/+p5X1DdX+2SMa8bvmFjQ8q
B52kF2KDJ8YOythFfh4DNDisS2Q2XIiUsKsW/eCLvKseN8UZ4kuE73ha7Uvcqrf/hlOjxdbc5dhm
wKfcaC6VDRZAop1t3n2G52mmuPfvPut226V1a1vhoUqOJ9ItoYqdvFla36Y0eAwisA627cjpU6P7
18PPAoZNa58P4+4DWlL9q2pP4EUp/BnvSCsuTMwu9o4zpFX+naUmdsJYOTQMAB5XK+9MAykypfWM
guwIdCPirxog4sciBsLX1usBg3OXJpwFXIGiP2KDzyDUxOmwSLeL2DbFKPxxYMs3lfeJ5sFkVJC3
dp05yZp9JXlC2N8qt9KhEykLeUEJFYfDlITu4j5nc/aMoiv32ztwmPJrbU7Uh2EoNUDejs/v24WD
h4J/8Y2XqUNA0nhHretIyt7PtGomGFE6UFYbjETXjZ4rYnXki7UBNI8mO4j8LWHbUFTQ3q8WfTJF
5q+n9edpmXvCeEDL9WhgR1ZHYIN2fXpKROuY0FGJw/iZJCedE178kG6zIuktukIjP1BLDF6FOUxl
fCSH1KwoV7vV/+YOu/aZz/1JUnC1w/aNtEH4iNJx54yXH09fB1EJUnnflGLmF1dzJ7TJ2R5g4TsD
ZCFZ7h2yHDl1afwNYv7PYHLUi2ASILJnb3rC/p3xdWjjsFCr0ISsg4pw3li1b0BUw0l/Vm6HxQkx
PVWa7aBCyJ+zWc5vzYdntwYTRAITcgLnXPlv0kCD/qP2d28+GVhhwETplLP3esureGwovEADeJnx
6hceIBzIDKSBKwk9mub/OgNmCHJ+SQkJt9HIylguV+l2qDLaVgvpoJYlBkDnIdVxHoCmJ9iNj8JL
dLkvZ6/QwLbmeZhCeTjgXnRuMW+7ib4uzaGRpdRIQnnSounflm8W6C/8m7uB/zdUK2EOseh/eJzA
tNPCq3XUy8ETmGLAIV7Y9fEcOeuYfaYqSOBXbM7lW+H8w1VJgl3lqOV7CDMmeQUN2CtcGGFVspLU
wMLXyemjErenL5kpgfotvcZOGQ/rHiBeA9ySLdOhKLdDlTVmvTA0nFcYNMtzj0u7XzfMU/t9AobU
INlygvikDN6HDyB248WLB1tO43fZw6+vV92M+eBNWHyTbNhTdEx0kdsFD+we47Btt3tFH/LmOTr1
A2AxHO01lIHfFJyqQGe6bRy4OWhe1TZwdBBjhVXUJpJt+4f+Kzs3neWRCxVm/NfL2d9FQv2WoRmS
82owAHN13oUnnFN9PYSryvvvDnD5wKNoQAbt+U+7FiqKT87uxFI1KjESGQJQg5KgGQrqaonMcVTA
fdG/ujozDaNvQ2lCCkh1l5Njq6A2APeF1VnJVO5o7qh0jdTQwbrSIPToXCkfMe2WZlkY51/qwXZY
A4GIKBR+kqd+6HnpaOoOErohBZ63k6tgUmDI8pxdZatW6GaonnXb3Y8qXCuoPVrWOvtYwY0SKMtr
xEIVM+3U9Rybzr96DgaNtsBzybEDrtzNiSIpP/IGJiop6TaSCG8egDfYhEt9MJ33CXx6+pxoIMsP
AMIV6ZhisZdTXNzg6GO/z7u2fvSRnW7sWuKr9UJj+Qhjmrj3INNf0iMmD8fySYR3B/ytZxLV6dPR
j7awARS2H+OVwGpbfUjyhxnNBwNONLa+hrZrp6bOyn9ZiwgW2NvCtQWrR0Ftqjg2qi2oX78QCqCi
pVI/B4WRvtrY7R3c+hCCtxfP0PYAdIuJjTVxArFdFgdrFH4fvJ767NfVC3tCfV2wuTHgNg9vYThl
ieoyt6S8o3HkC8DLIemsTMcJcYoWjqBjfcb39YA2XKb3Sh8zUPTc5oEMaEUHEbGZZ+aPWr1FAhy8
dVuJlOR4/yESNZrZMu201QTIkNwnHMiZj0ScD320/TBjKM7uvv1HlIcbjx1xiYUSMyYfO+M2YyAy
Obax0bVFeTKaoEByI+eP5kWqDGDpfoMAGJ1zbQhoSv6g8b3xfiXl+o3jgdUT5m1+QN1RQCLNkCsO
EBC+DgjIPAW3d2/UCVwMxvT/XE3eF2tJvCRRy7RbBjgYewvulIrex5SmFvimJIwd46u0hObzSXmh
m9bX5Zu40nvX4tLwfu2UKN02H/NPnUVAkmxNQ9kwknIUo9KqxnWbUZa1vddAhz0xPN5aOa7CIra+
zBj+C7ZXUZ3YFDqgeB3aAEW8Fguko5zw4psaKxZJvAkA+SVEwig0BAGG9qKep/hCKdWvw0i9PGbC
zchaL71gR+7nuSPpmIQeKQON4HvhHqvOursiY6Q1ZQ6A+68F7wo/DPIYkrW0J9712vp2QscxtDE7
UE89Xa+NI8UXFxonMnehR7qRr1GhasYmK8WhBkaLwn5/yRSoXBDFu1rSmiBIPcQMHzgYzbdM7ES4
ZzDcUxBf7l47xq3MU5PdO3EFWngk/rWknEjlUDD58FMEeDlX3g0tC1LbFjavuZlJzlu2aDaoxems
le2AmV0vAeeBfTqe93ha52UZKiyhBsfVni6sdJJTxC2TpQR6d4e8qCCo9BEQ0rsuX/eHcjo/4EGL
p6Xe8mNwWyHAfblOMmoVLgvLgHa94liiMNP6LvSs6kph9xiC2f1Al/2dezVjejOOwN7T9KOf/1zW
APhWU2PFzqVmZSe3uJuLNxhmRMPAikNNKshAThGvRPyBMkSsjVAZJO2bFOvZrfMp8w7v0om9u/Ig
qbxhnpTwjVkB97IuiHBLE4wq36KO32uuI/iZ19a64r5ePDZkJ2rTbC9shXqWlivcM+H4AEUFJM5N
U9Zj8WDbG6X1hIirQsQQDsMpT/7K0+0andT5fZem0x12GIKPoT3j9d1UGoek7p38MoB76xAshcim
CxrSkisa2GAEzxSpb8q8JX9/DNpOATiNa4E7oNdr9YX0lZr7GP5eMjmXCgqjMNZ+OAsXBJeHHbti
WphsrqCda87GI1Y8KB+oCO41Ol2N1TSeOkVIuD/08qOYAYNQI4brauQp+gKng4WkeTsNHUgyAVDs
uFklJCD3sBiltyK8rnaE2qLF8Y3DnVHg5tvyhJUJmH0w68tIeJvR+iMkyOFpo9Lk/t70S7OUb2pW
q2mOzVyAd7TIIRWI90C76q3ja00wF2TIY/A02DtUWauGHS03V/iyGwaNb6Gz4OVYsYVaq/1q6SXd
J3HgUDJjt2rJZ0wyzsbm+lOrQts5oP8AI6OYlK7vxPoHuwklkPyQPKeScVFKUiKqqjxKPvigfPRq
4UQ4s1g6RBqo/X5/VNJatm7hp6FTjEC73F47RK6FATANQJm+C0ynPHYSraanQ4UCQBmbOB+YD1kI
jVfoxzO5/Ubhh4itEGpCLUaiJLy1Y+IDbncA58rxwhrbsDw7+2EPazHtNqyJDCtdjMZzmkTRZqGl
fajXbiU9BJzboiVvFP2NNQqw2N9QjZjXSNFUBTvA/X1GOz1iobW4YOERB3/yew6kZ9Z9oGLbConF
AciAzk2xYJDza+UsrnUzviaZ9CJXdInX2gTxj76HAq4OItMRtamkBRbKAd50kdyMYh0yFFAYM+Cs
TKQtk1Ja8MZvzYNjD4xAdgXEXF7tQckfhcHSMZOBhOT9WKqLx0c84GK6nBdES4JQ6xbuy2R7ReJx
Il3/qVqxFM7fGKuCcWCmrY9RhcGUVxeUV4FKEPDQhHIzXoqjs6Vv0ihIZYkDUYYJo4/SnfH+ghO2
HAZ4CBYFcf/K2CgK4/omQaKshN98ka/9T2TEQWTDPiF0kTT8rMW4J1eYhqmni3clqfpLx2DWfoHU
pgCPNzUWSErH9JqZxq6LOtghoQE9MViuGsTWsEfPt/umvLhAvzXsXpFSm05gMLmhFL+VsQb/Ddd4
K9NFt+hwdIjZEaTtIHylpGCdwevasw8O1q4bRK9xQ/TYZci7E1gZZ9DH1TBvlbkMVIYuG0BIGWo7
RvphrrOO+W2G2QYwIxt4FWxKaHABNA2fxMTr82FOW02ftkL2nh73P2F68OMytjl8xcITbIiBvp72
+ahMGCd1igGgIeIuApJ5/K5pexDhyIBxhSRaoeKHVxDICYS5RulEA+attTVq3kcADQeOM/v+aSQP
iRn4UNqCPThP4LKIVNURKud94JuFGDlh30uQAjpyxoipNStgbC9bmS0TxVCVyYtJTis9xQHjqcSZ
HMjeSFXK0N/Gpml4WZT+CNpwZxVSFxnTV6s/kQlXk4aMwVs8jL/P7J5Q3TGMwXY395QxDbG+57WB
nRn6mCbts0oXNHbgAGP3AcyOpjW5ZQI56mHn+nTxmVnVX3bctJNASOyJ9YYU5vV1QWORcE9s3WVs
wRKDZRecvcpu2w80wRDs8nr5YUnYOeEBEd9FKXuo16GWLgPDhz2jB9K1gHXXDOGjStrmW+l+mQRh
fTBnnJHoz+b2igA5Bkv3V9Cpm650xGZ2kaEEC5qdVBkNH65ClNXeFTIQjnAj7TVLkx843FqV01Bo
fFNZSnfg0qzYuxo5YEznzJtKwMppb2ANcVZMAcDRct3P/x70/hMga6v+Kp+JHLk6siWHt/M4Pvsa
8/JetryaJkb6QuF/czDgiDND0nd0rirrg+DLzQolL/+65sh9KEXh8438VJlwapkz1mVziKb26EHQ
7iYPrshj6fXkbmZGOkDqN6VFI80R2m431/k1f10IyC23/QzkLab1AFl8qxbtFW/36MB3P80ylfU4
mrNN9y0NLLAYEzp4PIHuFTb7WVRwehP7JOhkX4llCRlBeballJY61EugQp+gCXkYgTcQ2UNIgtYM
nP0Rdiw7CHYhk1zIJ96b8uB58ToHQNDS6QiYeOg/1Wt6HROx6adKWOTDRsQWw9NpEMEE94aVj9hd
P+5Eh6RcL9K8oOt+bFhATu1Ilq+IrEgRh3W2uxvB3J5TCM6npos2EEEDGth8wDV5VxfY4zB4TekP
HiLIzn6bxqH2JMi9IbqsAR8Rlgu1jb9/B3ap80seRXx4ANYh/7SEBAXBBG8BB5g1KB1T0fwRaRJm
Nc5LD8HXbxaXWC3Pz2xmWAoWO+HtnPbU2fCyg2dFR9vQP1o+gfGOxdOLgVP4I/f9DNhh/PrG9w6I
sPPUy2h9tUREqvkrU9NRgh8imJ6+pyEkOEZAzBwmIAhxH8oxSU5RGxkNjp740795Pou+uetW/1DC
+gYqUs4x9Ut/v0YH459/0Z4eIXolz7Q5mYg3zoj5ElL+sAplD7EWWGxB5+e1W+OmXKp3IzgUBz/e
vSK8YctI1QRGOeXFtkGg28sMciF8k2fpinv8Vp9ptR/IziU4zsh/3d6QWTe9YFW3hlxUGxjh7Pr/
mTSI8qsor3tqRYiivkiZADoWCOdUd1/EFC5L4kRoLTcrF00hjL8El3g4H2Yl7rb/GGeExSVXGC17
xObIfm0bL9LpUZNXAwdH8GSeDezoQgDtw2vIsFe5UVK2YEDqP7s5xlzVwi7ZykT5fU2sBoYd1HXL
I70Jy8A+Eg8p942GgEK6/bal3/KPvP7CP83zHJPUIRLeXkIgDWUq0GzDri4MXefouqOkF3KvkcJH
1pe/rr0CIgykyalSI0F/T5EAQ8fEgL+8k5qWTo5Ll8Hqu5OHHY9dff9s1NNWd8IyTML56ddEB8TK
e4afRziDIvaVp/v/nxuMHZg4aJXKcdoisckPNSzu/VWmHAa32eJRKoboDscvunXnZ59SwHu7ZdiP
C6qI2ibj+Hl23BO9l9SHA1dltwtA3mhc2oJ1B5O9/t58QHl0a0QEMIXkuD8KvBc7axpQDcH3seeL
diCA5SAfxpoE5HLQ7zwX0RIL599uFY/bG5WwtCz9MwQTxPCq+uJAeH6Gz5uu5rGeqk4vaseGjIfP
C1WZWL3bi4DBtI8XBZ2DLPY6Ns+n/ZAyBOIgrSK70YFA/6eNXRhTwUKhtPKsd2nHFabDdzA4NNva
kHISKY7mqFReF+r/1sFm8Arx17clh/1W/IRee68Iv0Eihe6orUwg46YnSGYEGl3VZIFq6saRa9cT
NTY799ZCjxorvRbVRApP+UxtxNzdtUl67jzvbtK0xOWcTtsUG5Okv47fCxPI7onKS54HIgu/JtCY
7ItMM66XlwKuxNYkD0ItRxFWDOLlrpbYaZtzbDYDC7RYyw+o/slnQpWdsd3h8eys11LLSOVoCMKe
FYJs7EFUaQKY9VWFE+FhquLKFiQ40hxwMRX/yd1CcfXeOAMb/HWLccam4bXEtxtNRc3R8hIUFkU8
cn8DoOj6hXX7B1I4RVohoXsMF5JxZPb0E/MdTvD7gsalCRhIFOpprjHSz3Fkz7yn1rQFjYPLRfIb
MtLLw5PVHn9k1HXB6BsobYla23J9JwNY6q2UeyNTI/hcC0sWm4YAEb0GzG5e/oZ5XT/uuudhUuzM
iqCq1vKNhKTk9NmDkSfTkq83kdj48JsUGhlhIeJecCC+gJWJmdbHWiQOK3353CLbjvpAaU/vtuy8
hqhZACmQyL2vM0ePFksftbThf4bXykSYqvadA06z12yPcxjxSCVan2P6W06iJ3zN4N5SFFrbx9wT
qxE0JomKS9UOCTHJM3nNIymd5rhswS0YKMgG2Xom+4uUAG274EzaBz+coyFhYRG0DNNIRb19Rw+f
KdbtDk4oZbSgeASGGHZM9WaCAvZ+G5UhoTpym8hVHqToXJho9cMam0/yxIDS5edje3zryoKPLT4O
v7juLDXGtvFmQa4T4yEgaaVJwfzB94P1i9rk2HuLWtHoTz7bCGHtwJ3TY+6yHJXGup3Yhn2zLtA3
WEV8iuaV9GsfBpMczZ+wXeZpv312TZ0/61qpVCM2Kx6tlcKS8qEKeQXarwoXy54yy5VU4UlE7GHG
XLkHAoGxo/RUJ79HUSUJU976MJYt0OdCXmMs+O50EgqKJu/76kfL3VOO6Nxj7TrbH2nHPwxLzDqY
ob1lThP0a/t7JoRo8MvZZy2DzqIwJgloQEXpGdKLP/bBFmd+AzpTy0kXl9DCVxccXMZ6HrmB6LPL
DPgh08KHiyZyTJ9tT2tTuds2bmm2cCB9fOv9Z/V0eD3gTH65Zi8RHBlY++jhdqA1iy7Z3harg7M3
rFPoosjIIk15eJVVqkJiLqrCt4Aq09FVH1sfibbD2sgr5u8mkXgOJfII1XUx+4kt1TKjm9wrrQ4d
cylgp5RuegmvhGbaBZkNVAuSXC6MCHNFYxSZoeRo7sKn6Qy6xvsVqCT/xGIDDcUDgndXSG+zpiRc
03al5XCfuUnFNBRQRx9KcpFdvFYplWUE8z1roVkmm/7/fDMruhlHOo7S6FO097lssDfyCEqoNEip
d5SuBtoElnsPW4obGZK6zf+VoarttIfjkyZe5Q5didwFDm6XldrI0Njv49VkXPOzXWttL+p72obC
PslH+C8oxiZt3YwBPWbDmoJKiyfZ4nLH12WToLW5NVv9XB9s0896Juc1p4kZwVUpGVYIdwV2MnCu
gjAB5ZhdFU5/TYXy4B+DkwfHabASHJ28AV+lxIjNAyiRsFd3OZwJd5pW2W4wiNUxhgsuvKvL/j7U
aqbpPcJyDP2nOEvS59zSvo6KQegD8Aj0t4MH2g0toW2UJ89nVIih68WClg1klmO2R5ZSYHWNjHMc
+iIB2yR46haNDl/ML70zkDO1VrQhrdUiOaNPVDy6B0DYzkxHGJgF+30UzKZapDA+eqkfTULfg5dG
FohxmGjo/tkYzRDwyNNuGa3U0iaM3urdPTop059a//Yx4UjgehiJ/hErvbiYyXTmgwU9K95pUwR+
JUPonFW1ZmCuxmhKBIWn8BYJ5yuHvDJGaHWWlYVriuXxNKQGlJMQ/iKn/h94841WJNHqrJXQsWky
hED5Zh1aI6fDFO7ZgFkxB5VubvDydPBL7oZn2Ocu00hhTU241JNbSkypHbl0ayNGQLVF8KDiMqFl
szBsV1CrtcZJPbnnSf+M85ZGje2EeNKqsrG8AYtCKk+QRHUUYfPQKnWXbAXO/92sObG5BAvnJ/pZ
MYgJOoeoRcJ5kUrL6KBoXUqoyfhPjv2+HMor6zhTZp384VvYXiZPYgSXHD6n1NuuGNLsS8r4knMn
shrn/o1xZMVfYlst2rDyNJs7ftAg6ZeY8TsYWQbHCRw9Cthf3TBc6sOquBGg1VCBOzJ2shc7l+27
uyDAkatc/XNY8wfi6zZtlr4sRdNfcnfGtYWRF6ZmyqvMd9YybNikFOvacvewtzhsK7QUuCqeGEwA
UWGxF95nX8vUeMc7CkEUpeeM+nlX5neZiNypsw4q++q6aylkJ0ltXTcvUo5yObsFoHkaX5zWYpT7
1bPgkSK8+iMOo2oI0YIk4nOjnjeZxWQ7kY9Mxd5d5leF8tovueSUrXICg06/bSwqjvqg010VWhNW
TEnWJdxnbcx/+dL+YDhIOTri7OilFeeP9e2kriWVhpzC1IwLNj12V8TEkSLaGlZPYNbxaK0y42c+
IC8smYaU45zoxedm1e9ts/Iv7mrAXoz2ld+0XXd1fig7MellTdw4y+UTS4bPJoiqtsN6hsQC1rE0
pDq3DK+nZpHiZnLYte0A4amunlDT2shkxFWXCwJuEe4MCfef+VnIrZT1xqrSDHejB8HXf6wRFwSU
gl0lkBW/urQlRkpjVPzWDu4gxZSjHCXZT6MOGLo1MfYS+D/aapTc78LKC7i4l1D8ZYnZILRWMa/s
YbL0DQRr53DsIMNgyllCUzWYngJV18VqO4MjYbIE28A7sudw9ZdiRsdxx6+iuzr+VfV3F205L440
S+Lht+1BfrIp37HHZrkFXUCeBYXHT4iljBdf4xvDqr8wOKb+HShbrxyuzRG1uT0X+bDm7rTi/FZk
+q4/dJY52Nw17DdS36Br1gxk3b1rLUnWDGlWhlpTHTXZPdZPlzyLFaQqLt4OteX+4MfFEwdEfNUO
0fOdsGqFV/OtnEatROcpBkkrFHRxqG9D8CW5GMCrLMv7Wgvqt31CF7n+H/u6C+/45m0MOw3h4/xg
40Uvo2yXeIW7aycIzONCEGRTJXRHMNCcFUwOtiPe77/fcxC774IyTixjdayLo4iT7j8QIhZYuegU
OigFUDFjgWE8UTi1wcn5+pEc0heOwTibB2uj91Wz/m0x/iNc4ULauiuM6aEOFmmhkv8hYxcFoJal
fdgpv96+5fewWy0N6XGUfZQhTUtyX9mKyzzJxV6pQ77sHFLWU9FZP4gJzfFHEzCVhwVKFG52aqTf
Yo0GIYL77HiMk6RIpwd2NNiCYFjrULOcTU3Uxm0Brq+BI2D4klkCHSiBPgUj4rBFo7x765ZHvVEP
jK5e02JYRlmma+aeckMBFLxmzSfYKZ+8IxYvyNYK5G0mXmPQq4hAz4bsWSZZ1AMQ6HrTRTJZQIDa
T5CRyI/2oSx8kDyjyto91FPDSqH2/LPC2FXC0MVU4QThYNEYs687PCQPBEHZ8pQY744G3c5SviUU
VdWBXFsWOlYZKzw+jusUu0+XF7mIVe4p/adI375yN6tTcE2Zz3/JAov4I4K2hEggYqMSKmaQpk0y
5AWk03KLxS7sEk1HeGjtzuaVxu3cKYfI3Pa3ivTm3YiQpUtLUUcvnhtUIxaOqPNJ0GE1JplI8nIl
ljgwdXGANGy6pPntooP5DvSeYAZK37T3fKzlkEOfRVJ1Cx7pCCvn9GTa21RO0pGSVGm3631AH6s6
PzIEX5tPujIEdIc1UfpCjf2kmcL99UIqQoqbgCBs1iHZqfZMuTM2epeRaBv6LeaEboHa8+mfMSBP
xH6l9U0JwuBpUZjsXkpKx8uF/OeuQw3ptJ1Qnn2p5J/2cnI+igPj9kV7cUEmDaHcqQnEFeHu8ayK
VfxFG274+lqluLOvAUMY0OQEpIz6XBgek3zx9og11Gqw+EYy4qL/U3YYK4UgB6yApLLEfpubg8Sz
GLmaGUprrSAyjlLkv9MOreIuYYmTJ3CvrzB03Clxd2H+D4qhkhA9YpKYlwM9UF6fjJFepuTjN0Sa
rK8DGCnV7tOiVBDggTq6KO3kcgJ8m5hZjRDe9w4dSZkbIJRbyleTTXS9yL1ZCGxUoNnx+m56a+DF
omgB0hN+poa1pDS/lMJnMoU8EomYXeNRGhuap+qBh25sbyu1OAwcsEs0WFscB8mJbCm1i2kf+YdK
6QfPfDp9Ynthx1e5tGb86vJ/SBxChvp0i5Cp2f5P5ZCHLOKf38AD0ggtS5FMkqgC5PqX49bcGU+V
M8lSYtRxU+SaS3B6iELzhOCYmlPOgX1Bx/3N8I98SG3nHlc3ywfPGf0u6C0nLXfuHl5ukH8+4nfQ
o3QSNfTRs0a2KWYrgJCpdipbrz6qzLETwi9rDnpAubfl4NaSzM6+bfQLGQ7wZHQGEIKpFI8D9l7R
WFLe4aVUYba6LX/u3LEPQ3nK2da0iNaPWlv8xZlOJ+JI2V35jiyGB6Ilrc0fTwnS26yVzadQuQPI
pOpf6MTkFQIKct/lnE1C/vnXDBZd8fFWgWgtrbcjMEeDfjov15AnKMcG3MQOActoWj/EOKqLlpAa
E2RoHitToEA7y7Y62MBJayevR1xqYKDK3wSSRfv7XAIkqjzZKaEXSTEV+RxTdR3k04Rdw+7eCEPP
zcaQnaJx+YFjF3mucdAvazZSsYq223JYCQGgNV5UXrRzA69uS2lLldb/zMaBS3gc3zz6R2wvFG11
cNIfon9dWV3FWFywBh/jhXassJ+MflgwnU3l2ONYQ7SGBxNv42HFm8GtnKzQOZjapKZBw6E/7SPL
kz5vBJ8mNseI5WK2+IoLf7JqExWjyh2p/LnAHc4PMYt7/7D8rK0GAhHpTVEG0do2LQ+uBt3gm5gK
oCVE6vzyupezR9JNgfNjxIsGZRlxG/Mqo0vND9ZQUES+euqo8YR8NMgdYI8QVtYKdYxXS0JeIqvV
Pq/H1Qnm5yn+mqUbESZskGYP/SdQkHNjFDqg1ggdHHuoCNeTaOxPxnM+e5CCPk/Ye8XYDk2QOYpT
t7lVBnjmatlBkvfLa3lqna+klsMzhHh4X5+hKdO4JhrYUZ/ryTg04WEKLCoV/zsPPKFVIG2MPas7
ZUNnFJE7DPEL+Iuu1M1a9uade9WSYxtJNKZcDx3rUOyjusZF2jKBlQY+PREdH6+5fFKJYvdV55ik
+CMb9g/7rnA4Ov3MMz1UL2uwXxbGs78hD4h1u7KddV+Mm9w4UHL8/32i2yACWBU2GFvuQTBFzE8C
OPUIXVyNOMaADvz5a7QCCS3uHwHU3ZXfDKJVr5W2/ZK3s3m6B8/cI9BQ98nerTZieaJyq8WA9nrh
3OEc7i0CXTNdAuhZTmHc0NsGbErcqeVn1BzMCecq4ak2NVCMy1qSwqmVp4Ks/K3px0F1E6wYYxsD
5FCTNojIhA4qeTnt1KXifK/c0gsIKqFKFCNSlSrjxuKVnuUbb+6fW+T+7KpviNbGvicbhvvBUa28
M42yWmD6cdt19CiE9YIMM7FiLSwzvSVs4tvdiFBB1sY8xnJ44sJLo4glESioSM5grBiIjpDqvC9B
v2URtN4Yw6vkjJRLZqqDaKHYAkI1jqowSTnjiLYtvsp1wuoLNcrIrYHwv+m4i/BHKy0t3KkmYhJm
GHWX4W7UHNuMuVfvITxwP8/X1aHwLyQ1SwIwzFXj7HnLJvn8Gtgzg5CWu5RDd3uenu9jk2OmurlQ
chtKrto0XKr4BPhVRyheyEy4aHdcZPBV+5MVzyQVjq2b4h4pETnGr7LcHtAZfywU2x++CKULOHwu
PRR8mogFKfsYS62kDmU4d+SQjKkR74QDVMKBcHQtLvQnT1kYI2VdG3j9BL9SeQ8m/y22o9HKUdwv
Z1HBcRalQRqVfaAmG0yE5O/PSYo8HfJ/5pbecjk+WjMj3BfuloXd9tnBl5N7WMouPzjZqxlwQkMF
n7JB/Qruw2lUnTcm3BCfvyQO9ofdmSwjwljCJkphdcIwSKS1UW/yvR8MkVBVHpizIEsYIKfDXS2P
zMlCu8oQNAawumGTCUC5GQv5CX53v/tHi5usFf9O9Zzo4HDViZ2PDJfynbcWn01d4tOofGIwRWpT
6zx46h/okvx6klsAV/uessK/++AK69g2K96xIKwen4N4nnBkO8KdLCsWzRlgJB3CNfTkTnZK6PxO
9GZeFCylmEE2+rVx4+N7cIjiagMwI72XUtkTbqCF9SmBLyHTxZ3OH/ayLmTS/9WYkeTe11mwFIir
/7SW7unMdqRCVh7T0VPfHcvv4VFlgJ8l/fTQY3P/HJEusxOBP4RqIKNUkp0zsa0DpSS0rotKQyIK
MPhi8gIIlVb4AXEm807Wozd5M9D3rM71IJXU/YKr+QFNqrHb9b7L/5w3+vXEA0KojDKwv5P3oCKn
l91LypbEH6WYgIWuyMQUnCe+Ct+3mU9DovbVS/VL4b6KQF8h+H6XHWBAAedcYZkN6tahS3zPyEDz
0BchGReBRzF2BHyM0S4Hzei7vzEVhcj1PbW379ZrIIW776FzopzKiXW/0NH3c3PDlO4vmqrDISM9
t8Rnsn81z3p8dS+0IcAliGDfk6CL4DtDUFNV+AdTK1/DhR9Kh8yFEJMxyIFgsgcMgLj8fdw+9w8p
u6fENJIBy+Xx/CdOQjvWEFZjNiNeVFy3HtjVi2/LOZUnbfBuDAl5iTT6hfwF3c6asrX2fCGG8p41
PEeofhfk72sriqmX55L4nb/pn/fbg2WnU9xdIF59GuXcK57OuwAH3NKxd6F6y9yfbdERKGbF/ocy
bohFPe1sgamI9sjc0FhbOGrn6cAgz2qPvxWA2IYUbKOAxMEeIip2dSAyqPH7bkXHM/aN3M2iyNI5
dyCj4yoqFaOO0BTITld1a/GnqIGj0VJ5zcRqv0cZORu2/aTVu1quqX+/5phyiRA5GJtKdYkAlG5Y
yUPGa9GRcv6rn5PgnBv7vbALVY5xWj1BP+89DLOIvmxe9FRvi5FY+UPrME6wNu/rRyjeBSASirwW
AWbzyqdFPagvpF5bdGaYt7hJLzTLPB/TjCXgwIPNVskOiHmEOZMOOcRS2/UR9BZElALjrKlbG5x0
ZKbpYnNo6rfYotMltwqu8cIYjldkWdZEQB2lspIGiQehgbUMhU7xem86rGAlmeFRzHspaktKpdHs
qINS/1KYdsm3q1o9NY0cAcuxOndJwfMb8XNl5kc8kRhUmoa0SfIFGAnWZOWRro3tyqUw2lOOd2zf
55wA9RYuxV+0pr3DCfG5kd8GO+tGBIYQROSg+k/XObEYU5J6q9jlCgc+019HUzWBcwI2YRDCMFS9
wm5djXexFIi+kQ0ecHyV1B5UHPjsn5YmX4x2YbY1ZDyaKnxrgPm9q5tb1Qw7yPJ6VcnrA7FMAvbs
ePa1K1WJt803j9Gmqw3Levwppk6q0WmaUpaHAQ9AeQhYGO4jLnZbrPDnx3up3IUOX5Qm23ereHVp
wKAL6pUkAzsThQcFgHXxT9WKyhy7SkU+b6sP6oBWrH+ezxcK+MsX0bRTIHFf2taVvFhGzf+y8gRE
9mQERkyqZ1O6JftRrbT4gRVtLFYggIFEc0D6z3/oazXNB9L6zSz0L+0+DqjB+dhSAxqyRf5RbZPN
j62UHYB+ZQ2wB0fneh5VJBSUjWnE0vnVHZ5F7ZV+/X6djs74l6n3a3g0jUikUxgqebD5hai9E67m
xBprZ70TGvNNignRaYg3VIAUYHdgnYRjr3SPjvIM5qIiF/StD71ti3VkCF5YIn3ityuyWavRYgo9
zhLUDf2FSppTzSd+lYViqUSxwtEd+OBHtRux5rJ2pqBOBd6WM0l7lIRl8cwfu/BYS++kSt2kPCSw
bAlzea061VEzRJgpz1r1cpR9/eQba04X3V8h482gtitC2FrMJk+qOO849GTu5Zil3kVFNJfCYmqy
gpWEcpzUuxE6v0uIxeZDcaS3AdLlyzo6aS2bNSzy9m4/lAX/Bk+Q60nKEVmPe1f9K0840a/3ajR+
9SpvZvPL+EpZo4K1aSF1ASzSxDXR+l70Qd+dJ9fPOE8iK64JntGcvPibf0RMYpF1EvugUJ+FP6Q5
ansB8cvbLLoHftQymMFe7qu7dCrcdQ7Du/7nmsAYjT/1ZeLcGbiyFG2Dy/20C5kveVTVKgXWzmYo
3FZNt50mI+Nyu8TN6CWzOIkugIaXqrKIwxBE6lDk/WekoOXXvhz3Ndsdmwh22vHmDX4FCHiaGO1b
Vl13wcT5Ln4aOHA/5YM/WseVkub4YfJUJACPdz1ryaifQj3pvGANtk5rYrwWXRD97SeOHl0ulOTC
yu+pVRVbuZY+gbJspP3EO1nk4g4njKiAcFB/K02LLbTOfowkBzHey0hBNR9NbKKLdhMBOvAtQ7yZ
N99+I1PHPGL/HtdctvPD2F3akZq0yYDk+dSeKc5dLvB1xZ+po2+dGJzmEoBzC/0WkXRL+0LEn9yv
nn9Zb7mRsGWyaK0DbN9xVz00isnp6S6btOKD0VooeJ5ehEOnSspHjRAlyLiE5X2xiyr+Hy3DldkV
+1B9WJDIR6FnLhR1H7jy3VM4+aX0CNMMFPP6ZcoYEN03OMFPWcx6hpG0UO9BiRg5VQZI6F1/JRzH
dlDIVpcEPOiAB4bQ0wXTYl4bJ8oEbaEMi1J5dmD47xdpCWTFDj0aZDGL+VzScVKmG65lCVr0Wamd
dftY3BCctco9Jr1I+PBO6CVZjOTzPFlGseKnv2PJq6D2cQgoCdjU9TEQhsyMi5X2D9nmwE8h+yF4
15cPnI06tBDDHiaERn8WilrOk6IQ9wXOkrtQNJzp18K4F4+rhUmO3sOye5EfVi3ZxaolqcfRpFBf
CdeGbSlYBZO8tyk8kXo6j/52zAHR6sJ7xSJuqIN7blWrwVdH88Ifw85lHA//sMQRLEs2NkwsblbL
3Nl235v5ECbfVacgp4MSS1MCV7jdMJePChyotV78eO5zZbOfGNXOf6Z7WfwTOd602hNJmCec+1/T
Mvw6Mwa5oGAHi56/Hzcff0VRyWbqN3EuEywisccnWRfSw3yXPpLrQppiV8yJ3si9ApECLWdD+m4H
kk8yqxop9fnLl9VlOrFVV/xsRoWkjMtPkwD9s15v1PIJ9RuN53CjLRKcxAAo/UTk+mdl0bwxTPEi
9Rf1opOkSSug7YKR6ABmEYamKbBryyKqbn27muvw10n57a66PeYiqXyfAHc06sxOEBq0bA/exgPx
qkdyoY3OqzDEtTXdQXhthXULm+erKU3o24eMHWKTXqTldfF7boVLrqxdL7OJqU8+ZRkHCMe4DNPt
LB/gCkwmedr6YitaVQN00w4XGdPzQKYZPP+52ZWIA+hR5yHUmNgjfHeZK1FmFAfy1jlrvB8ggLSf
X0Y29BVWZAdpSqf2kUoYxDQQw5h7yOrq0i5EHfYR+iGcfm2UqFstUBVm1rWVk/l7BNtbmpMp3vJv
SL+aY0zVqWoFyrPCH/VWdrrCI6wgdfnegqx2XSKJ3RpidDUrzkUJUDsgaAn0twjtwD8TyJ4lTYSM
1moL4YqBjKpdzf/5J6/UspHY2mSpSJyhJRsPFUZn9bHZWuT8qvNqYvoTUzWwxGOB8lwtt/nLLPOK
N9gUtucF7ia3yHEiOJToXKtHOmFnKh2rHbDBksRA1d/zCZDJ6YRIgKgw2nCpUrofffqDDEs4z/+2
exWJAj4jsbooQeIxMYJYTfdgn7vgXFvJMnJZwWDiZsy4f0SKf4uPzeno1DE0etU74FN3PClVeKca
zf1GBrTOLWyPsJ7Fha8LEbh2wekBWbfhV9EGCibZIW8zo1cg2gq/fqQwHlXPd71Xf73KjaCOIKxe
FNOcn40hDtDWu31JHiJ9GmfoGIDkqkvKr/sPuIQpTxZ1QATibQuA4THxftcGvWZ2ry3PPnm4bP5e
YsTNo6oTS8jYDl4uPA/infcfycWZwNJPHhGxeJlYA91LqiUU1dsd6phajKCbp2baqFZ6B076ifjg
UAjt0L1T9hUqIgccjgzQQBu0oFAi+KkkqqoEJvVFR25xx6eRTMVa7rOBkiB2QGGDXlGC7yixvSFN
oMccXEUJ8tTlPcy6sjRIo23OTBxZDNm3lXNYqnVqFxjfPUFj5gGN+YqEDJ8E3zpTk85r3k3wdRq2
frgWaPEWBYmghc+EXLFLG1V4i+shu6LZKnkmYPgGQJR2sUp6ioLNvvAVEoLR30E2jnOM9niQgpe/
Ih7C7QnIBrvLrsxBeGwm987KhCyyCfhpKgsPlTAmFEkPoXpz5nt2POOyXydjzffDkZZETkTstq27
hlvSdl2O43ON0rQO1egO8fUqBHa3U5QCEh9KnQwtxL7AWNk1qkMSNqyIIrBRQZ8cv5M69gSDA1y6
Xd0O3X7Lz7w9xe7ia7cMTbpU+wCFcQekSsBpYdjr9M+VgzPBVVinOD9BMTQPAPIOB5Wx9J6TfjlM
hUdcFFC8PiKKi8NWoefIweR8bR2DLoUTBSOmSr5uLmFyqraC6VhQDuCitnySqBniY2HEyIiHVDNo
Cv9qWQsOkSjFaim6hjZTtKX3Xhxh3qB+WIGtNxpIskFjgRKekcIENSW+b5z6XEW41SvZZfS1+mDB
9jBil+FQpI0HcGFsOFu1q4AZ7R9efE9gTviuWZmUEr/gxNNCSIGc/KKjUjgOnPEienF0r30bmStQ
haLkqSWUF2NmQAbJ91dREvzWV/LPfOru75upg65NusGWW84yoUd5mSokFjW74peozsohHRiJMNrP
g3DiUwMaHbzCeN6Xygqr1Zx8CnzA80uNdIda9tCH/j7yOshLITk5gH4rfRAgY5wiO4LNnJahg8Db
XlAOMV+7gKnw82n+uSosyOJTjeGRNu6m8UfBi55Gxycjnm16g/ACbKcRJQvJF4Cp5Wev3IPsYA16
KyqoVj8xnqMrslpGmfvhpxHUpbCBHJGOt8eTS5MBGNXkfwrIyBkm/aNQNOFcO5pCa86VStH3P00d
5YV/ikhl1dW7JTvsTKJOwGBv7+SFCi8wTEuibfE3vNS0wGY84+XSxMkUOvGnwtJ6G8DMro/1yPya
/1Ho1aC74cvt8xTTNqF2kWEh1VXxsvbOiLl/lZ2JA54828EGYl0sxad9vnBE8HNfWMhMcMTJ47n3
hT0B+evbuRo4I4Gga0q5Dm82PRiNJkXrimREzINCwaa6vZg8mwlxZ7aIX3yPNC2TWPkBm3TXPuhL
zuFfjC6hLhc/XH2WzAu+vkggMGRmPMYNUsMo6ky0B5HmemPebiW4D8g5e7bPOQTxDEcXfab8EQsm
zLoDwY9U8w+09PsHvJkkd27cddwtQVj6gZIcOJQH56QckIlorsllBpiJsUuB/17yNf3RYw4YZpwN
/DMGzAqe3Zy2TG2Px6BxtwBhfIeOKPdTERYYOfueC0q/ehQSGSGdHyNvcffR1obLNj4MYWkVlNad
xhRaFJxEf4xx8z/hQC1dUGNdxISDmKQ1ym72z0SkiBxcvVKHIKiF/iwBSohNUAjbtiUjKKlEUS60
wDZ1YSEsdlWeZQwXn7FHGNnwcGBr784Xb9I3mlGpA/GG8AyHMXZbiAAfY1O1bCSyrO3lwUURT1Tq
a+tAuWjPs7GHVHS/C0W4lXAyQoh4f7ekgY3AxveKyQMeWvKLHcc23siZ9B+HKR6QgZpQZJzJYPP0
J2EItKoILr2kd+0I4SqvBLXiaeO0tVYv7A8F76do8qutSm6lZPThhlvQBLMOqehFWdlyjPLdVnHb
GyexMgb9ySwhVXfwOo/Ij62aFlj1KFAyPNAKriQC3KXApAcSRQiC4XjGGFLJLaoVpeHvMbbFJkUx
Rgyf1sKVwGTGXVRnEStY5q53EsTs/ASfhMgwDLkGZONzlAnwOF4mNAgLlIaYCKSJid8lwiPjBWSe
avu1dx2NerU3c/4cm8/D/4kPVVSvgPL19oQJSag8GJmgV+ncBgJGfXHxD14gSJS4JdMBdHj75ZYI
IDV2WmV01UloHeN0r+lbq7wqExVxvhUcksGa6CVKoXqnngsas0VoQpAmnuUaD2iwwySj9Jfgn1L7
EowoE28tMTyU3viHK6nqtzOd8Ft5CQeJfwBQXUc+mAQu6evbijcvIY64JrzZXOD/7wNxAX0X4mXQ
bLKSpwj1MIRqLfKSkH/jbv11HBynZFLQ/Vp44bNFjCyvoUfaUOtCu2nQB8d4i2xoB036qBaut7y4
VpE24EvAwkUzE3aLeoija9JUhTYiEJb5o+H7YaUdpdFlvbqmIs/d7RamJH2R2W3Y6qhCj/FxSY3X
D0+KovOJGKV7IIJYIEAnAL2EAyzNnN6io3WRsVuRovFYVLrkiSg63dl17FUc3tWJp3BhsQlVOqY1
wJ1N5kNtvAAtwAvFT2TVz5/S7daZQw+grxQdHLAl/YSJFnvWax7VV1jXMisPIrsNK/C7xOnYhs3u
l0FSvOxSzTh5UhpVlyjghpCaYgEqRyG5nuaEerSi72Q7Nk2JR6qMTiFRhhRxO5caVfTxLSN7fsqO
cAQ5m+/yco6ALRj0xhLyIFIPPgYH6m3fhL+6iovcsCmKsnnMVGw9ryhAdZQz/LajFgIYld4Xq/K4
gs+o+j8AAd9Mdk4RmYwaIwUwtp3XBXAvt54t4Y9Rkzo1cV+QH3XOg2xn2anwTMtTrHoW9mO/t6/i
WVcNT1Y8TL9M7s4qKHHhY4zTifmCht+v8ilFFgpdVgZ2kIPkBQA18yqNsI7ZRMssql86Vgs7pfal
5hwjMgC3Ycvfe+yvNnGVWpOyXgZG+nbTgOnj4Wdhg2sraB8WI4xYDpd9HmmM43zSdJ5f4SpxVdJ5
1W73fjZjzsmjfsUqTcV7YBWlk3TvTyxkrDBFoVwvxyFrkcRrpZ2s9caUjagRU5PalrV2vz4aksEJ
sIU792FUY9ydHwVWGAi9a3BHDS+QauTkcgnUD73ei0Q1ESArlQWXn7D6hJdS+tlHVxzcKSI7D1a3
GlRoEnmZCVKSgfO1isqj2yviI3AsBdGZBKOOVNR3VKzwEDzkd5aCP3kjLCXArcQWJSmgS/tMMxQe
Hol68L/HdExwc+SFEcgenrb1kmlk6xaBU+FgYC7OzBFFzB7BGIUti/AJH9PxIlgh0SCqhkFhlBsL
yUDk7tGTaNHRieYG/5pUBrsRnuFFmypC/gUORdajXreC2pxWsLIW0erA1rwUth8NPpZ9rKRhNUhJ
zxXBIAGXXLrWo5ynu6QDEMoolXxyOurqZH7cZJdNref7r8nA0Z7BNo2A2TS2r81LUT0fOjC3D7sD
CQs434UHqgF/OnIVNHRP3RfqoHHWXpKMTIvK0JlgABFdG0Z29tCbhjvRm9l17CtyyafeRXQ/hKdN
/jLrrEnN5kOV7iAvbbTpbtNLtkvhFah7c6wszxwsIoNJCvouyAwHDwzSF53KEHHcub+0/IGqm/Ua
r4gNArDBj5qjVX/RbUbPwEd/EfVR7dM96/OYdOJ4Q14W+eTGuTS+JQNv+FD9V3o5HmUqxBxkPsTO
VnkP0tImI4b+gBf4zeqFeEGFPi6NrbBKgZhntgxSMCz8yf/L9VedWXDRxThp+uj/Tzf7+zGVFLEg
qMBIsGF/acFNiWt50B4BYNGPgShSzHXh73U0jCfa8aeVkSF2Vr46dQIdV8aWwjXlohCvqRWulqL3
RRJErQFcnxbzRvTdVbmk7KxzH3SnPhh7UDAG/XOEgkep9en4q1t7tGhApO46OLw2gDub4ybvnw42
ZljjcYKs+fFrtGLUIYcNwBCm5OBg0xmfHHKnRghJIlKjuqpyDLSUADv63wRHE7eNRpDld8UDKpD6
NINhTrAwTdawAwVOzWn5B90R6/Sr/qD2MuVXYKpKvboU0o4ZdVczzTvRaun37bJsQ6B/YVKyS2FZ
I3IuG7ignNPa+sqPU9F8cDdY3o/thbFnlY/PQJIz575F+he6OeIogk+KN2LClZlKt7/leEQFXlIc
y+a34no8ibkXYlDPHsooXsIf4IM4iuAcUb2LPZXkprDlrVAMiU1JyNiWzuvP0GQQY32iOSitxJ9b
w56IgSpf8AGxUy0xQYeJT9bE/wWVgfcOQjo=
`protect end_protected

