

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ya253+37kdInKtzN3pd3f0ykMvIJsSTHE2tRr5TaFzMStJPqyqbq8G0/aCj9umOixPoTbod1oPEi
NM8lNQufqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZnAl3olUb+r5fzAKtbT+P9BDg9y9NfOiCUm1R2Jcpt91ydHcXeu+pZ8D0lxHNM0CXXGhs5RFFeCB
fQNmyCQv4qniT4fHHC3wrH5hPwmAH8kqSEyGt3c0SvSsHCYTeXhpF8Chp2XvC1WNZGYymRNjehFn
t70d4j3zNeEsu5WAW84=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iKnL/TA899sfLGiFOsNtfsGv8lNgBNaSxC78jj2+skMz/TodvgTxrRQVQ/h/L38N/D5FIkKYR4II
+olODWgmPzea4VBkBMLQ7z2XenA/M8Uvin39meT5Qbx7/ksgG2EdpyOtsmAvmeXZQgf/A59DevU7
Mrm0rcVFwLpmjNvbnBOl5iGpGgx6v231GzIUzFEiOeCx1PkRai2IOZKE9lG2BMKHN7Bhsm6JH1NF
XhuV8OyupD6h/Fr6EDMMNZqriSBB1MM7btJKN6VC9jmTT/Bega2BSYjqAkfYdUTeyup0UqEM3znP
2BL1mUmUOgL1/UMAmExO5qz/A5ddH+Ai46kqhA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bwfblhQfYU7J4v01pOh0vYth2hZJ6Xlf2qmEYdxkErcnbM5+VpJUpwU8+A/bDOJB4gUPbJHCeAw+
tmj2AabGe4D0Pf/UukkjTsO8eFOUvoPbwDwH6UV1AKQFszUSN+Z4NTgaKs8pxWumW0juNgJujhCL
2ChBu6ddPnHdB5HG8uQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UTW+eKUNnZFWLDMo9paR505jK3kaKnyoN1JMPNm5SlY5iSmlguqsHIHMaqSHkHrYg25dIfFqsLa+
ygBhaN4bDhxyus3QZ9m0sw/aVS4ly/5bNlw+8ePaK1evrFFnRWDzqTt8U+H1O06G7NfpkTmeK+am
Q1esOyihSrmjwIiD3aw5SiSY1J84QcBDQl5D2DAd5uRtMADgrmEFzx9Y7yHel0j2iF6Z2vom7g5G
7K31eIbiTPvCntdYde5+aN/nl/kdiT8a+6o8fslm8ZFdkfMYbKE6CsL8CG+5F82TWbIzOMfxbILY
sXfUaKwgi3ZDGoeeudit9zXCRYxReIG0hfQ27Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64272)
`protect data_block
14LoRk28HTX3/mvcSUvv6IhZclTT4AaQ13DuCCJPs57gI5COvGHu2MQfC3Q2zaRX1zzzF/x/4/1x
tJ/vwk9WpIScJHJh7QlG59U9WY5kpl/75H9J7tTXJuaFnutGmZM0R3c+xcmiJ88E9Bs5QTrN0tD1
Pjl1zalEFZGtrBPo5hff/1Dc7HNOYPO5pw9IU7sjP8dmb3EXxdrhQWRUqZujWVwdiFtMMDONlJ0s
J20ikWLSgxNVkegNJEapXMf6Q68beW/DRw0Tlf3ETml+BfV6F1eZMJz71Fd5gWvFl/HlJKba7MM2
Vxb/BMLzT2obt8TYZ9DkcJsNiwdxy1PbDwvcGgKExD6gdo8HL9TVIHVr2tBLhfnmIKijNcrLjoFq
bzmuMyZD1anop4414s+QRZgXm2n80uyfqkja2zfDIBEk8hUdx65MNSRHc8wsbAI9RBl9Wg7aE66K
g/WqDUSk1ZE6EGpqaEkKg8jIOy6INKysKLU7dTEAqGA9ltwAKnSdkyAzswcCFX7PZBS0NIFk9ldc
HJicv98SIGQ+pj8nIa+5TjbddSIXkgReeB1LHPoalyWjx8AyGqOX6CnzYMItfJZMDNaShkH2wFDn
vpldovH02bAoGl4H9Jopjv+LTxQXSEnWC3XIH5gVn8h/bmAnOZqAalIOlbtzA5A6NNcI5MpKQD1Z
wjsrK1tzILszafb8UJ+WrmJ7t6/nTlv2mtTgWPNgUzA3ZeGbc2DNxRRV0jxGdJwZFEmtZ2ypVeF4
UEcIL3b5G5AnAhRqVORGEPDF53ZHWeMDKjIyocq+OW+TgAGvhB5nvq4xvE/Mn7KFKd47lnqQzLPK
96O4Gi1QJUgvVVSIXmKsKJwJ/D/ZBAcOi26qLn5+A7SFXBjwBeJTlbXQS46rsTn7rY8ilGa9oq3R
H7rW/UbP2lIy2zCDav0U4siZVijj5A7zDtjmt+hIl0/LPFrEk3GnWnrQhq2U4aNIsr3qz9VazeVv
GHZ/IH8KUVP7uiMxylE81tvK04MXLOl8sVutjp4sPN7m5B5WB2lVunqstPKkqzbjl10VEBkIrpog
Oeelb2LOKnw6kTliBKuoPAcW6RYN0HHcsFF3hkZHJBa3V7Uh2gZmyhOJQNwE+uW5ca4PooekfbbN
/0y6pTEr3sDx3Rx+v6YMUCwtS1pf9AVo0a+JXa/SrUO+c+SP+qIL4GJCaJl+V7lEdelkcDC3Sg1/
Pz7mOKvtZQ1X0+q9TEZaQogU6o2Tvxs25qVitVuF3CjYGb8ChI/sjVc70mfbLA+t63Xg7PGePQte
uq+YrgWHenqCs8DIOgOQlNRQGCybwBJlZ/86Z4u4jJN6kRLlfloY8W51xu9Cj4G9ljS+le9hOLQW
xgVVU5iAtm/oiX5gToOmNmgF8V1LVwftvpU9vH4vHNVgX/gCvyhRGvD656+xWqK9ucdJ08KO0gGN
/CQ3CmbO/1kGv2yIsmksycFP/kGc7e3BKgIBwHhk303oxcROJNcFEeWL0djcT5LxHOcWDnFvDdDB
b1Jw0rfo2oYFuzrb5uR736JNvgDeqlmv+0uMIIwePic4c/uqZCyI0Ja3MBYVnCZiB0FDNHSqNtIJ
Fmbd1Y+ror6VLkZBiaiLloKZLNTqmV3zsAYPceAXdBCH8WqWtT6qQjRXkgl6Tl42csvssmw4gNll
CEtY597FJdGi6I98exFKa0b4Imw5RpkZr4wy/luwl83B86yU56I14lqwd9U7p/CcP1QqmsPlkGcD
LGnogttm0ArV6zAMdj1HkXrISladXwgnWhdBU6eRpsSCJa6Rca1WzIbaHfpzhb1pa9tZtdop5ujQ
UznTuNARPZhHhrVAMSlSiHBWGVugtuiK3qj18imXHEWVg9svRppKrwvRbtmy8pOBwRN5mOovLutx
n8qptOZjp0EkFwZaqXEq+R3gajy0FM36hfsmsefhfrjDt40YM+fExh693VKxtoqxngb6yHUKZSpu
nGeWyumZvohBSZTr3GAhdzEnHAulED85JWXUfedWxYbi04G0G9IfDSUUhD7HuZz00DP+HgDm1J1S
9bbwX9qt9/ct3AKUjgCiproGpq9WpwpZCHeKkS05AFtldsONOTiaZofseowVXkWtq9dJ3KgTyrlH
lJNYnkMQCUQAv6SpcM5TVVTV251IV88w0lpX8i7Aqpot4quErqUcDxZG7BVdoYBdGA3absfib2R8
SLjqjwJjFrfDnKVcpsykK7atH1R1Ks6iVOviOo+8zZthciHr1SetMlLE9neKmX6lcl7HQ6O1MUzr
GsDofEBdkdI4wNWHsDseB6o3WWhIrOwJuvPrYx7kXlsVhjUz+mI5Vh8l1LmcOGakOBHxG8L8IVcq
T2isXjdYXPtZtPxb42XUM0sE3h0Kj0BY5L2VrCsLWfg5sSGyv1KPvda/xilScUpRd3+Ukoj5ZeMt
DS7R1+h3AS4kIQHD9ukCxjyXHHTtTeXoALuZ32l8rUzPMlZ9inoZUwSvfSLDzTP7hs4liI1qMdR2
PNJBaLlLyLVjz9wJgqLmJs0/g/1SROHFJryPF7L1XcTwvbijT9f0xMSQqJfU7V8xrbyGF/TKtLvu
PtZMVs+reI9/1HWxRD2IC0Zajag4l0L/iq5o9v2K8T9WN9WslIxka+/sW3rUeFtWwr6YwJY/oL2h
peNSUN78YsDBAdfTK4SJ0Ke2E2LUSfsHl1LPemv7hUhuNKEgpSlEZW08RsZF159eed94wp1AtG2b
DU1cN9ujGpeb5Kh0Jvg8Zoc8DHsIpEp+t0tr/a397MWDmVQY4joau1QGmqFnonDBooIUcX/0aD71
WZ+c/YrmUOHs/TDRDoIU8jILjBjzOcCLUTeAIt+T6R1m5Srj545QRB7fbnCoYMFluyk6Zeu3LKml
jT2BAgoAPjPYT/ZwoJry4cRsl/eaqeK8Mt5hh0ChWKAaQ7PfRLdDdUXJwemCO8QODnT3WUmjM8yO
YfQ6JVneqvRPimI27rlU6urisal74txUZ1+3hNk8AxMoI8pWeanob65nGNTytM0Gl/Wj9s9oSY9r
8CEtd4EF58ZSYt0XgdZMxEJ5m38v/hXsO+I/wtDwU/wp8/pD7b19h9WLHQPqPzhWzUH70JqS8K6p
2kv3VYrC3zwSyXPYDasL5RqkVlFkuTh+ifgmvz7QLLAJGbPjdNDZiVcRIdijV+7D7AK4oOT4o1ip
4QJnwn9ZyjzM2UokRRI3jqAaxiAr7aOYGLvQSmceUuE4Ez/sLLRSSuJcH4zSf4Y+jeMiHShyOv1K
e0obldkRvgSdTWRKfUxjdfPIqKm+aag7OBSsFAGGxpzz/1XVJN9xtkkcFQYH346VB/nabr54qovT
KbG/OruaXXAAaHyzuEu114MT4PuM94velWI3yFArm5DG0E5oc/rPqjHMT634+qZIZDfKJ53SpM9e
PWgUgDV5JuijvYO5cNVvFaCEcu2KBGrGoK/yj5+2N1WT62qVXX7U41WL7wnel+248MH2QxgITHau
BiW5v3UBS6foQl+gAJEGmanIUxo4gnttFqU71yAWqUut7wsIctkdEGSRpRhfV8xExOHDgS9u76MX
HSu500udpuiiWarZtXasAxvonks24HzH6hhC8Asv+7KCD/aCYty/qYtrPmDj1aYVQZLXGsA+1eg1
aCcSUJ7IO+SlnN5s9PcWZM3dj9szBzskLAB7mpOgCyRqVAfXExEEwvMHaChT8yBSy3ZLZWaYHCdg
CmBlr98ARGGl0vGIN+bWWw+lxpWucg4ipMoNKzhj+bhYlPNldfP40ZwV9fvleN1skw6VbUHYXTEk
2rfMrfkqHQPK3wkIALSryksU3Xg7B8XjJ2ZNuuFwvn6gQjpXNQxeKJbr0FeRls6UBY/IbnnELD6X
Ywj4GrbE8hHky2/Ze2iSo6reXfoU+3J5QSGDEDZOmb1u3ryQjDV2TYGruFo0D7mKdajLhaxC92Me
/Ph0arIf7YfRBwE0fjFziH3TF2ryq+I7A21pr3TRqGluYcTzYdXMx1NxSUoF+r4oSgTPCp4uFKvi
FQ6LVd+McmV0ZWeAv3oaprFjDBmQh0NkzhFqpYGxmuvug0KvO30GQUQlD7l3SalzeJFZ+5Z6jkQ8
FO5tYYBuTtUHqV1yPO+LYM7Pw4BO5a2I5w24hzZQB7tDs0MO2r3g1Avhro89PkM7cMbbFzGPtiAR
VqL34wTf0wmbs/3D+wI9Aag9L6UHOVmlOamPseoyXBkzjwnf9FW380u6coIaduXeB9+cWwRDMmiC
j4lj18mb1qJvWi+xTtNRo4IdrI9MIqZ99f2g8CeSRRgvYIqzsbS8Ds7I87ho1fpUwBseaa6XvPDZ
eYKJD2pNv6SVmDxYPiuNGOnRtq9u4u7wu3JbDo0emKjmyASgHTTRecJZ9OGLrflFB8ODivnG10fY
GECzgVEm0NZZHoBEIJCKlOT+TeRhoabjyJoE6Y7XilvHjQQoK7KgYrnQ07YjVnFfoP10jeNz8+cB
yAxI2XHk9Uog0XS3EToYMeQG5EJmrv1a1k+jCzCQ4m1+eTvQBh5IMwqAGUFQUwdCc03xM5G+4iOO
9ZdD0bV6dOXzdy7L3GyMhQJkmYHyFNB+vECeiWXUr28C+ha5OJMBapASfEJBcl4EdlfSnZqsmw6L
Yc3tO8s9lERi4ptlna8UNhX00OHBwn6Q2AiCrm9HeZ3QP0yAFyooGcORBv3hNtilcH+KlU2GzMcw
09Rv6KJCZCocXVjMyuGJ0pvmj93EKrRpZF1C3wn5Nq5dY8GeIxrUpD2BFg0MFzsxp8HLYSGoDpLh
280hPqA0gNMYJWNqwzPaLrGcenUv1GHt5m8DRyyjXhuvtIE04kkaK4o55JQSn1PBV+kutwCpLBRN
PHEx5HhPDWRmtmA6ZFcTXpL1sJmnbbOkUVLHX8mfcObTYO9ujxotX5XeaTvKlcxCyG6V7w6YH1UY
jObRP5Cf+dIPPm6+x5PvL9UxgujBFLfkdqsQRYrzGTH3cV9NN5GESwnyw9xn+N2Slahg9xlAvzUo
WqXeZHuhbUS4bu1YqcHcqV88XHcNAwTu4HkMv9p4uGSd8nN8r4+b5RC0KaID0FTbZs1IMRHRrvY1
7UsNVH/l8Za0shrsyX3tCW0azkoU+aHxswpQ3vJshr2TeoYnpOhIV1bso4CPruGPAcbcyTP5FySr
2DLeF5cxvuxLovMl1R6PK8pFm2c97QCzuy5T03TsmAwZhE8O21IbLr0SScP9ZLZRGmyUfzmcCKUF
il15oCkI2WxJHOaV9EQS5Bcb1MDSZGofbWIlbl9+NmFvIaGw/4ZMkEBw4/8GfSjlca+M+e3Sz0WA
WD5afEhZnj/9QNIhHDs9wZEiBSUERrDClDEtOJ0s4NCUNKmSu0vNYLpgWP0nEkCuzPJOB8adPvO6
C41/Ew0d1sL0rIiA+emKIFu9YoKc2W4xxKatsh6zxlebiz+OvaE33vJHVC2K3kRn/V65uqKFvR3h
AiD1tgOq0Gz5HruZpgzEm5HDYk3SKVYoVqjZFbydxNKlS+DLm4AQRhV4GeOTKUHFNT/k7P+r6XdP
hgmaYIKykNhaCNtLtRJwnKBUiGlRLmqYCQbnOaUmZYF6c0QRYTRlIOrGR/j4eEOFhhJRJu5SFeFF
vCKyS9OExU/fMeTZl0+/SmM4YEfRnj1FOnaNmlDlqSilZ4z+MwI78cnfO/Dh1BT96V4r7FJtw9/+
p7m0rftxmDtb85WNhpfZ5wI/ynKPlP0aFT6epvYApFWHRYrhhmd1n6wNRLL9/Ir5aizdnT6j/TOl
+XRqtbRUu8GYb2S8uLYBru+biS+bMo5h+YyZ3KgQfmPBf0YluwQF/jqJEfSV81IyeswpQbgEGRuv
31POumelI7f3RIQ7PGCdvqib8c22rTMgKdceEYTUTH+pDGpy7c+7mJ0SJc1NK0l/FSLyB2ujfx2H
UKrAlMlzEU/WCaQsSTRdcEGhTyn9JTs+O436uhG3vRdLqFf3Bfq9sfBFDwU9Fp1PUEE5jucYa+7I
5CjX07PABz3/zjGPg1dGO75SL9C/NptJdYXOg5TG3WGJCokm9xLIzmC6MDxJ+FZHG3dVS5zJdofJ
FlKeJkQYbLa+Bw3uKv14cQ/GP4xMyMNScB+OrvpLRZe3mmevwvTtb3KihhdC9lejl8ZVaUZQOG1n
+abUhSj5bTnQ8fu7xTwbyMBxxKjsDU+HXO0Z2suKgm6QZmrZQtOPXmjhoZsGtU9Xm83KFcnNDsii
hmYtArQJ2FoKOvNPN4egXjPhWhvmf5hL0AdMs+WIMkZvD1mY1rr+oPyBZtGXa7elxZWSwR9bAHce
qcUXmmehyvJQd91ToibqGd7i5qkeIZPrGmT9tr9wErVFgdzCeTEKGIaFIS+J9sLb6DLOVUIxAZco
zT54nHtagUlCDc/tgaiaBHIoDkmjLDReEyTFeNeuhgLsGALJGVyamHPgd0MZQRlp38i0VmrcRLv0
dHhB2DrvpbsMLUBuAf+2Lge3DytquzmjklWnifWkQ2ecSeTxm1JhGNeBgPpknIsK4+6VkPvwWYP2
HNDt0sVPniCbYoXNuPl91SgTBPjMIe0XRMkeNzlocbUfgCDfyILbwRj8KBIM77iXcUrsNv3CyycC
Rh3Qcn9CYuWCAN45wn6ETpetxcVD1qMOTCnezj8iJ7UfwTeeo3/u2a2Q6PBgALkJMOi3YYOKfMJP
BrH7mWTjPl2kn4nvGlf7eJ/omCeyNA8/qkcwaBh8GIjpj+t4u8zn5nB4lN78JWQ+mTAViSpmfBNx
B10kKHqxgKi7bFy/489lIJjJu4nWKPpY1dEroGF91UOyw16Mi7yo4yRaBnpbjf243Zmlai/TuOWX
xu10EWzC5UuwQKaaIZ5koR38UY0XG75Mx+a4TfaXk4Bnm9Bx+SoRDBep9XRphiLyZPpddD5pDeup
s8J50OZE1JrhrF8dlFbdtc2dCtsIUErqYyIC/KskEiRVNVcN65Kf4YRInQZ3uOSGG/lAij5A2p5/
aj5a9rzCirQ7SlgffwGuNsvzfhLutY/Gl5BqzWE72Q4vEBb3QPEvIy1flUzoLyopuFqbxPqwEhHB
wpbsp/BgIyysGZdxbdAPjFny1tg9Ac76bbOzu5Xp80xY3Y7Q2NeWmHnjehGWsRu//PMh+OmcVCXv
0c4qYnmx28wnOwoaKhiCV0FLq02W9dh+iB+90/ldkMSfid64entQiZLUBAEgbyrUTO4OBSSxSt61
UFFnwnKt9SEIOLrDDSGryh+tsUkFS48MyeRy+Rx35maOVWtBN460kUPY7bPKGBbN1Gvu7AswKpeb
QHDly1IYgniH6ZIbgn4ugO4a4/Wuu5bMCzUYP6ktrDR0O3gdqT1I/0dlaKvWSTClEvfPTaWvGVxM
Sgb1DMABNqoLKHvoI9g1siNneCZ0BoJfIWai0p+QH5PWIyjz65L880IIhs6D7pBc6KFbHwQFmWnC
RLP+wqOPGEHWgwvxSVFrF+YzvxrueNeYIg0AvSzzIo/jKr782lXSVkNtJ3Ka/4zhTO8YWEc56yiS
3BwFPMmyFhvHi6N95vT2xDDfpIlCQMpnRGfhZPbvQ9ISZGN4Ef8kPWV49GAugscrmfrL3KIQ/6z1
1rWpIDIWiiKmfEq1lru3VU3ANulMl56SgXi0/9hI4KTnzy2mWSgkD9UKqX5tUW4HYHU21CmwJomy
5vddA+4XI4rH8NI1jhquFGo0fjnWSN+bl4JB6SFghExdu7NwAFlXPZo4lsbHlrSoXOvv6YXh3o5J
4aQYeU4wi4XGrRu2WGdmyqTcgf9vUK/6Nb0qOO760d+FXtJcxkvUUzjVfE/nyi8/le+BEHPvHt6p
mlm4GV9+XiCDXJZPOWuEwQITUixvmPr0/bCsT094KCkYUYU+ts5Az9OaiBgdXC3qinoxHPTRLeD3
CQXQ0R9HpROGHwZIufd6Dr7aCAUjiHypyWrgoSTdOg+64n2r9e6gWVErsze3dTfT9SeERLzDjepi
58TIsLEXt5V2g8d7j+D62EEEnVWTQfa1enYZTr1Ke7BkDgkl1HkOY1zq0x/tXL99kO3Zhq5JI7aj
yzmJQTzgCmXW5qvaEqwmzQW1T8zq5EsEREw6poAGagBTgXN5zL3jWVG4Ii6jxJ9R4Lt+hfnPV8Ib
60LDl9iENTBfOKBUx8V1vzuNPUdJevVi5n5IwggN/z8+X4MoIrvQRun+qfCItZHqxTAEldl5mJtY
B0Wx/dqLpPytkHqbRfOfqO66wJEgLAWPdacwyqBHXpFcy6kvvaxEWbx9Fp04QuE1+Vrv0CTWrfOO
6hrq+lVOsRELBJP4ycXg7tiVh8cKmY5DQmtfLqAMNnkTQl0+iu4v4FuVQJfbb3JSc6Ur+6Y9nUmM
sJEkhwIY0FFvKbjDkkXjSLWRJ31a8A5IlnPIK7KULbyCwHWPdfnA7ab5eXIrDSTktUWQHrcfCofV
b1Y2TmOSFV6SYgvuFdh/2d8F7FgzuO9H8B2iBMs1msjm3KaKMZ5QykXVlPc8XbiY2X7CTzzu4riJ
wkWO+jLEA1TWxW9MD0j2lRRBaR6jUVIYPda0fBYKkCFez3TgnTYzSea8XVe66rgOSb2uQyrKekP3
pCJFSI6w+yQggnXtpnkpYoLgqB0uonjjoZ83GEnMx7Q5lsZWapfJ5lhWWdZrHOhInoxMQI4bblS6
mR8ymAGqsebP/YVrV8DgiO7ljEOBwm23gfjZtmcEHAdNYDi9z89fnTr8HbOXMF89vW36pv7vOA6D
mkAZuZK+K3n/iP4Z0Zy/P8afLUynd6+SgVLrD1yY8J4rj4jszlAWVmJtghXUp0erlqkojjDIb7iW
Mtk2hItoeFieA/06kGGZjEdiAUucY2ai9cHSANezlD9ycx2JYnuh+SjF/9XI063NK7RfpnUOYXq+
d71CsxWmi/r1TxcjU0h+P8Ukxd5WwVNxYC+ig0Lj2Dg80lBBJp4DXvz1FoK8d9pYS4keH76IQoiN
ESjTd0C1lPTCTFVs2Z7KDDeWwlvAizAk83wj3jyNP31iqduEgexw7pSQrjs2kCRgQeg0ljwpT3mn
z2Ffk9HlIQhB69KFW3jSMMHT9pSQLdzHnEaZQnN8Tm6TUTLsf846ogi/RV4I4PTlMC+599Rr7kik
hSBdFCTkBEd6QfDz/rJxKxtGwr85i07LGh/hpLrG3fcpzE+TXaF80StuxoIlzZ3y9qxgZwfAGEfc
NTj0d1EWjXIzpgDMPpNhdmYAkpb1xVN3G5+PFW2rtp1UXfV5gCDx6o/XL7S9qx7/V/kFSrX1U+zt
6GX0LGCmmGexsIOaElljyPVjFFVtqgbn1HR7jxHuTnch57LsvGFarrFzP3go+162B/G515nw3Zgc
KL5ZSOgi/9f8pyW3Ll0vuZWJgmsVprSXJrgkppjeKYjO7aXNFh1IK+e0NOw4UnSc2On9q+Z6j8Q1
Dt1+fscN+vSSh1GHmte5M0v4+pq43ki7nO4+6KjCWeIa2gX+mBhss0LAfNTUm6KnjEkAapwiF/wy
XAR5j6BSiVhMfXSWIVwCA7f+eJ6+Qhz+7GNkEW3y5WqxnoSdqbgBTClXtdB/cobI3knWxwRCoYVy
/40O79zyLvA/sZP1V2NJAnX2xHr3G7/AlRc3SJ3yXYijjEKWWfAvqw4iLfm1TjU2LAOyhom/zp1x
qCze/PPmeomq4Rrik6o+w+wuNVP1WmdGpr+1HqpOjize5Mc9aTdyTSWHv+Jfw3NG5GYzgDWnuONf
VwDZxxSmE/4uwlZqUa+LmOKH0QXf0BvfpM3xSqFnJLbeDENKZ7el3lv4Si+v7I0m8i7glilYIJXQ
h8gEqsv3s5Fb3c7RD1CzBCpcG8ajXAvP6GCjLz2DWZfwBMmsLf2iOONTK3quT9LQLeZsToyjdv8D
6DQwMaAQHAVMzLxLQQgW5mXitLNdKkNXfU5GrZDO4yzDk4mUxi0N3zsRfPh8/Sxj3f1+J43xpRc7
v2TJ+nybKBWZRl8zVKOGW5gjyoHDiP9iOccEyeiAln2kEFNbAkRj0dwSaicopAnpjbfMemFHK5YN
4jC3JtJLlgm+lEaisPW1k8104Oc0E6zrKNUnVRtSs37/k2lCpA4LwcNli9tWpqnpE6l1ZfaieDTE
XSzdUN1s917TgafLNuCeZGpghjIGcc6ABoeMSFudYI2oBBGV3sYse931K93Lo2yGUNjVG+BjL/4u
HDfTDQgxLd8ntp3bBVnIsIT1Ycc02MGyy+F6rFKnqEDqgTeu2hPtyGENhJ/jjgWatW2KK+YAsxCl
u7bFG5Q0azEZy1OXsR/Mktvy9Nw2mSatRcblGkq9psVbHcjr25ibphAI4lHeyI2UzBaBTiabg+TL
3bhkjIHbP4yGxML4A0GWJWisDPyt5dAN1wbI9tjFCM05pu5YOG8L3EDYU60AKcmkI99KDdIJoCQX
WPrtUyjL/jriY8lepOJHJH03Moko9K+YkSbJ21WBh9OroAziroQ4DhQcKzQUcx3VQjNR35hBAaJG
A6eCRzzDAQXCFXPEElPC/okhXt6WCVlmvQeqAN153iVGgsQbRGA8sK3VGOD47HvgQxTbcPLVMrTg
q9hpT/r1Ut1g/xTTxLabYtzYn2FsFc15dkFjilPlOpfGstiLVg1LlI5/3Zkub3CLh3mL93L7h85O
b27DFhz9vndNCBVXZNtelVJnHA7T9XD3TupYP7d2r/jNifjKiS98BUNEcw8Vp2utnRS9piHp6tbA
DzyVlvtz3OOYsqmIOvNiSBKTdk6Tq8Kifvy5IM12+2vh3oIcyocIZhn9AJdWM2MSY1YDf2mDfmLj
89dT8UpZA+biBSBq+6Ux8tJh97GsvrHplhkZOnTleG44m7JC3kIL0E16sLk+t5xXRq/RqkxwYeut
m07lWTCXV63L8TBZUTjTP0m4RbNgaEDnU9nC+8kVyr5NdRxe/Aq25XzjM0gQ1eJMw8zwwmYvCwz9
GsvA2B0y6VrjCSUC8ZuKixTbDtJjvCFTU1nWfGyryW4kcs6NKUczENFuIZKATLNp3Zxe/gfpNhf5
iKv6fkuNwFbN8xGr0+4M3Jhc/HEfYYtMR2kX2G3xWQBx+FT7uzb1a7DX/TVWUgY3Rd6PPmegjfRS
kUuDOfrJ7OlMFn0PPdzFAi375gItgxMvOH76Zyh3JyY2ihWHHWpsLghGUJw6iJUKvyIVFLhG5fG/
c4NMK5SSmJxjAA1sdGsiTaygznosPS+B/q9df/RbuUvf0NDmJSy+SthHrPEVhX2de+VxGeILIIkT
7ZhRb0sKeh79xq+jAXQvKG1igcst7aAK4Fwgzn1FOYv4pX+VvzL+bC7WAfFCRzkncAZkJM9L3R9Y
y/s5vjomwjrSLfp1ZC+JKovKSKXfakzDb27moY1E8FFzk3LZKCtFjiXIpnycwjdstv7ejSxTNqQO
kCp4v6v0UAK0rwNLLKL/5+qEoftna/LalHRT0ZUKpd2uKRLQjIuZi+ln5Laica9G0t6rKZzRy1T4
PoenNniyILIIMln7piHiK+MU2rA+WPDTPfgz9iL6xFtrXg9HHCLrb3bSM7X7N88Tj6EPUOdZFdDr
GNZNVciaY2OiI+w5loNXTmzF6cUI6ZUeUCUQRi0MnJBkHSYuvFFtbutnhJTToDJGzFqsgmAiw5NM
2mu9tKgxbjVPPw2qev2BqSvWPtFREAE1jEXD0HHyRyiYXfrloskT77LkRF1aaAOHoQ8d2SjKlkoN
gzngueLjTbmiTnHnlaSbVx4JiosG4x1m/gf3cZ4xZiS029MGBgpAV41W8+s2H0zhkJ6uLKgdt67H
CL09iYeY5orntlWjNcC/UNiIQNyUyI40HUkM7wUH+gK1eZL6nGcuxKZ5SDMskj3t5s5pSUnpZxw6
I05U6xO6YGvmG+N4jlbE/00uv3eYK08vUVsjPU7scY6Sx9EVjbMcKLcxTB4as9YPcYpNqlO1yokb
HBtLPDFP9BBqzMKBvc0gWomoHrMCQLhpBHbrxCPPkWSav6Bb4WOjF4IBDd7vlmcykEElr4llBoF9
B68UPEbWvUBrHVRJws0TMdKHqTSceXf/QFcHonsOu6Kk6bKWrBns9IX18dzhRmvLBNbcTgFuAiiy
BcvMeJ1K64t66UsFzXqpOjp8nHHZvVAtL3WiwWRTobTm850tFVWEFk5uKZXBwN4WLW6A/Qf88CIu
Q7hRvI42A+jzvs4R6oaJimmcf7dINSpVhuG82ZV9OzAuSlFG5isuSbJpGsIXAdpR9QkzvWGQi2yK
z9DyY9nlEc0+GBNxVW26838df7Kx73W6Ql8nepRtIaMcsb+pVld1n9P870SMD0L6qfzZXJITnjQE
IqagN2sjN8cvDyMAjqmw52HaqQm0bDQ4UyEap4Ve894cT2okS8OmZvcIqkHAlGQJdqgBUMjy8YZI
T+InYXc7RPQqWGoAJKUS7DFXu5YN/55+OiJxIPUXhe/uFsjNgUCTEmSgurcM0JxKns28/xVYPVq8
0/dKrjsQyYDSyW5rWXZMyHWi9kVK1P2K19np1F3ClB/78N+8eaBW3mhggmH7FUxAAq0ty/Lwx7MS
3NQkK9vZH5lw9b3xMyt/mm7GkRzP90bMbnnpC/NS8O0EccUQEUXpDeg7fflEJwD7EaBlUz5ozPow
TZnTDQf2+xvskIk0YQ/eIJGa2i7lt+Ox2AYvj4+cN2CubVoBEB6g8IFRHsxK2yP+iqCkN8OHNyLQ
66hIWCkltCRPSVZpAOtxg8Oty8EltG1Z9MyL2J6e1Iid1yilQZSwwWlZ2E8MICT6a+oSQAmgmffI
23SXJYCR/c+dhtZ7UetVFZEL83nerkqtSejgl3WxClxDY5HGNon3AqqgVIIrMyJrmkvZZbB/fS4O
HQbucyQ1AL8NlDijcyGJ88ygFFPrgY4XlPqZWqpONPMEmSqI2yJHFhhUlvjOhkCc3O9EEjOi9owb
4aNdy2Ci2Nk4ukTMj3dPI3a7mwxVHB50uHaIctF0v6BYRw5vp3ZTL0yST5tYsbZyp/xeiWKX5zzZ
abLrJWjf2JqSR0M8R9EmUd+DLu93tkpE2GxEEJZoE7p6QmFZeuiUCCeKOg14hj3myVXDe633sCr2
tOocImD0Y5O3pEJRqg3lUgsZJhbnDav7uIH27r0sajComvw4bzTB0exit8/kaFY37NT+U8hB+yzd
2fHm2QNkVrSoV0AfvJBBMpRXvzechoInmj9yRrCL/at1u6pw5E10E9NctyoR91o6ol1BYK+FE6z9
y2RD/pj6p4WmUxEe/uAEpmCG7hr47nG1McvLMPnI32i7OVX3WmHw8ikgTT+psyorDD8j1hjNlBA/
+wU+8gcOcaYqLz5BNGTLlgEUey3WSTLSskWq9F3TauQVIdWf5hlY2XpgOpKXvPhxDvQ6CUDJbDwc
PlmNOVw+//DHeH78FBQxdY+MDBn5m9sLZ5n64DtHrdgYOU27Mm35pq95AnI66VCo0dOR/9Plyax5
/EiZzLVEZZBd7qKMtO4ArWlUFqR4w/VEc76tUb//CnL4w7aZfCnx/2/wKJT/CFnLcAesRpeE+O4x
p6VurkfvDl33OW7o69ISeyJr2p9u3yaDWm0NZRdLPRwEd0jY/aqDJyw/RCbqm2XDm9ZS01CrTRNr
We6VqvZkIww2yfQKcV6+4I7+liJcFqOmku1719K/riG+VUp490DULOWnB3zXbGrEF8FRQeHkLSZH
8nwl6NG1Mixa2sqXn58AkNvvd3PXMIlDQlFHZhUzkJkTkaIegcyQCoi9WshPrwpioM8pH+b1HV8t
Bw3mGJVlbw0eS31eu/e+IiAD4lFlEzTB3Erw7Jh/WhViXmpcjGYuUa5AudW2nNJS9rix05DaA5H6
4jExMHiLX9JSyDYeVgy4wMZeCH8SxmKSKkoxh+9Tku6qKceUpK40y7BrPigijt11TY8HFkCVXeDO
PQ+uQLVBM96XkvQFBu/HPRZ0zj5Jr72IttiBSqCDhMxgeliNzNdQJE6AD7BzgcBk+VNgggd8baVb
agZBKcq5vcbQmqI7Iq4z87SsHYYWkQ57daIM3mRU9d1PYUsynf7NtPhHhfy1PgN4Zsqi4TvUOhsj
2gIyMJ5FgUFp6F5vVgGfscflRlSHgzB4/Fdxepfb1pTOtJywrO86BXa9Pnb5AqhFSf8D5GpjmNTI
LEklKrmWCTEMTfmxwTSr8SNK2CLiUC6xIJgOfEGZeZ+UScpcsZcyPb7elL6D4AisHXrH/1bQDmsH
ISQz8qM2eAj9ZZTz5M4/7mxa0Kj2W++kx53i8oYEpdMEh+cIkhcBdl2Sf3GEekK+FG5/7PAV+2Z8
yIX3xurV6jNh+KgE7+qsL7T4ZfF5O7teo9bve8DT90hU7jkGHHvC23qifZ1l2kQ8H44lu5Dbg3A/
H1DhXSbxh3VW9XCr/2puN/WFABteubjnrHDvC6XHgzFF1gzh230vsrlg5ElXjvoAOxXw8DQofk40
uH5rS+8dWveFtzdTYZMylp0gw2gdOqvPAGXd3+YVR7UNPAlj+VemI8K1+4QU6/38yGOUpHjx2A7D
qPUvT5yuXCev/CgtRqP8P4cSUs51RwcsUC6Mf5r8cXeJVORtmm4B5+7S9KDHt7sO7y+39hRdptgQ
SRaG9c+gDy3BhFfQHg2v5weTwX6YuZahiHwo+HHTT9kVNEPbsDhDXg/+ebArVdab+IBXO6pOGfwz
xV1YDqKM5IQx6yiUACj8XpOPjm6o5ePcRcvXxpNFkSRX2MkMwdi0qpRL1lQHktEuVmHXeRnHpkyS
CiNvL2w2iXIr4Qlp5kc81PWEAKbz23HNMvBsdAys0NOFjG7/Ky/n4k3aoLiGHDGFSydswQA9L9hS
6IhqBAqYWzmTZeniCuIUooFDyiRNPnsNthf6fz/I2bvu2jZXa9v/xvuVrR57lvnDYNrxkPYFgrw4
2HTDNJG5bGEruopC5Bc2qt7FC3wfW6EJ20paV0YbuvojWzp+LSQRPNVLa+SbxpQ4+Cdh/11XMx63
GOFGkz9CQCnHvdLCZDpWn7tp4CEVzfdZGfEu2BMVwFKHNTPkDG/G/ebIkLFxenM4WxDuWodfdI3N
jgN3jKr2DYG1oWPpw9QdbmdzOcz+r1rqd7OUWJsiKt6uNhHM1eFWrFwzju5bHr3RTYFZc1l3XtIa
xcKj6TAeV65hAd97DB9l2klUdF4X5RXau51ztVVBFWGwGMiu6PwWq3AaZ+thKOz9zU+5VSv1bPHP
vyYSZ0G/C6e3Vcwk6r36q6GTJTv+41pTKZEaIQYb9wRYrOrKa5K+zlczmB4hsffkXoU/l+AWtp2J
m451mQxX6nil8QhYrCZbArfhIcsqU+KY3m5ayqivEyrB+DYMQLrGDVaFXTUiSavOTAZfOxJiEMyN
2RsaOVarMIh0EvmAy0kjbSIY+j4IGIx7IywhlvVYRaZ+W5WD2xLDpi5mvbBH77Mfg6Ukp7O1NQkm
W7RwmDxRX7Ydy4pjWK131PKKzk4TY+p+QlV8jCFGxeEuy17CYAsw72meIMz7D37jfV+9V+fytrQR
0BHv823elQ+qhRz7oe8GnmPwYDwQfR2T5or637aBgGktk6BC0REC0OzmU/4a6OzVXxntr5qxRXAD
aw7yj58HSA2vjAvCJD8X39IaFW2ZHmkYjFiOPGzAP9qlmE09GZZDWBMk8jKbQV+gZCDoLJPXfPsJ
vZngWwAnJLQj2hbe7sHdSwYp6KgAKDFGrdBO5/cIqpgMHo7B2JXJnSVXO1HSt+b6H2Fl07Slbhj5
KGIm4dAKNcEF7MVUyDi5XdJHh7D7zB6/sgeDhCBPj/wU87mdHH1xq6rPBFNx+NiBNRBwWkshsddQ
Ia1NpeuIzYXGnYRr7eLPIot+BMry5ChHoTg54eJdUV4TibVsEM1Wmc3ajohSWOm2P2+o7kYibSuy
VZuL3xmFoM5z5TgnrTJ7PFcDM2Fj5BAiA7U59BO105R22Q8l+x+5Tu2z3PL9ShdZS7fbephvXUE4
FT4IpDKoMCxFeg/N6xxCdhPJLFCiV4ialYhrLeoe3kE2YSQ5/v8IYMb5QhGCHCUe9FYHu7uWwSc8
eiidcIjz0bg4DBPWelro1KE8ulJaOIhfDleIgUExETFocuwKbWd3bb+XeQstP46lQGhCAt+aFFlj
doeuMAi1uttieJmPOUuDSYcl+Dc6qUDzEzlFPcIE5KbfaKCimUg5LZ7eVhizGwM4/n+TKY9AVv+K
MQM+sFVK83VGugP8AXxtQ6gttGoSJ64jX3ujVUw4v6mo2w203bv3Ps/BvKUgj6IdvnXNwoDL+1ky
iKX2vMdVKtxF4q1+58Vd6WT16VVllZf3KuSy0KHScAPr579+gWeagFxVz6vttoVAKxIvh8SxfyTn
7PCeW/DG7uBupCfoG8CmtPKAwrcsXNNdNsnr+fVYhOhBueiDNYkAQPsYFavmGiG9K8VNjzbs3LmU
jg38+vSPeZxyjj+07jMkkQnbj5un15BhSpPtTY45Et5E9vWIG+w/KPTglHNyEbv52487zziyQcKx
06zhguw+JZQSG+jski3Oy6ZAtpiFQAv9jf1SsePXK0tn1PjuX35Z3sdY8SAAR1vUeuHOhZSRXV8O
/LzsZ+4ZhmK6NCaFeJgYplfOVpk+m56lAHZiJsLuOc32InsGHMyMTK+4W7NDrkmWYwOV20f2crzP
LRwji/T6D/RsC6xx5wBXexrHaCCa/VXhRAImntvskZlaTMWneB5Qikh6aCTOqk7ntBxFxgWw81FU
Do88QSd4WpuL6oMKouLI5h0x888LcILvgA3zowR89XO/ZeS84YsMzP89KzEO9Q/1sOQnFyp6LdC7
xakE20jhQ8amgj9rzGXf62I1QqbDprc3QnY23Tj9CDfcwr/vPLLxrsTaDxzt2S+pF4Q9qrDYuNnh
Nllrf+6YBuCg5kDySr8qojbND+Wk73gUEFBCpWB4BYrovKeKMlv/edSJ5Gia1YjPPuQKboTc8D+F
wNawHOoXW116BrRMoJtebu8vchxMG6uSSoLO8ZIVLIEff9zMnlByP/UdyTw57QxAGSaBe1QFzxbZ
ojIdoYGaCH1zffJjHD8HXvqTGKNju/nWUhfBY24epCJ0PZVZHS7841DZGGGl9tJ/1yQmML1TuTCc
7mv2w9tE51OZiJ+6uJ0lVI3xG2Z3cX+z/erWb4OUV8UbCchx5GZWMNqTitvflXN2AKey1oOrLHvf
MuW3wGUUGL6F62+qsokbs6hZBXiWd5UazG0C7dnXNWUb5PkH+t8s93wNnGQEwANh6QZ1wueVI9+x
tBr11vaoftwmUZ4or3XC8p4JrkXE9hJ0oV9yeEldGzARAc+BtB+aFTj8bw3hk62A3txj88e86mqM
zOsRcRCrwhm0A1Az73Ve5u5m4ppx08JyMliTHZ+QUoG0Wy60whmmrPG1ms41LYPMwWgFBXsXtbga
2oZ+PjoWZ8V0SSg4KCo4FAdDf0lWRzHrMzfXf6lylJ1sVJOUoMyZgrkIxEYgxj0YrZmkeue5+j1H
GPaY6nDPTZGDUiSTLTrNWTFlvRBNq0FWtZvyg3YPNUZ4oUdSnXdzMo5liXisJnbCC0NwVXM6+zXV
ihUWvI57jq8n8x+ogSVr8AyXIVc3iOf+0bobEQycGI6naxM0O5polR6NNuFEaoZiDGgfYV71SXvN
nt3MfXiYWABrLdXwax7QOUkABDUTM3NaIoB8qutC8qUXKpK4tpw2zUnYvaqcAZPdEaHXnMHzzr8w
BH32mz26VUAQgc7JmcZnDMrFYEii6ahvIjfhjWDAdSPyJBhBtLH+syTdPh3h9qbwpX43tGPIphvx
Gr9Ytb/+D40B1QWb9wKsAt+ux/blXSLXwRutTydGsPbF6tH1Lv9kLGe/IoBKjperhcPxVkilbeFm
PsWVPFzvpWuqFceLMMchEAJYYd5aHFx2vBudMedD3cLqVqcCKHWSwD/k2lRPxBeFWH3yDaJeuhRd
5IvdQAniCI6teGXVOKFHm8g5VuU6IY5TgB2eW/lG41yfpfqgeC3D4QCSFlRtbrFmNAFP2jaacCTv
LrkG6T7HxNzCMmUdEc8Itn7gtNX8KzFqlLt5maTVtqOE1MDtqss1QrlXWUMlQZq77pg1TSm7mMnP
vzLX7QLjU92lmR0OReTJqGzGs+RrzzULQU4fPDoECXDP/XhDClafTDvDDzRYtos4QX4JjtcKt67l
6WR/O8vdXoQLSczWgg2ySEw7zTh0QWQEVCoRdXpL/94Hn0tGCs9PjxUlieJ7wRuGZ8odOJI+98Bq
U7k6OgdPzGf9wOknjcf5CKvvA6xUNgTsmLtFNaGzTrZTJ+9acv0i6IBaAzgneePYHDLoYebRQbth
atGQlfSepJ+52lQOS2jyZyKFsyCLZZQs+QPZ+bvPODGqJLa56Mnj9DY9k3fKOstQtU4AQivgTPoc
Fq6237chYLYBwdeUzqFmSI5OIZgGz65iLgH3GwpgFLW/X0M08Si+e6W+Gtq9gdx94+f0TC7fLItv
rhm11TGtky6R0IFEbhyY20DaLUOofEY197ReTRgLtXppGmpt9qFqXT73x7LpQ6Lesh+LIkS9M5+T
Re1lMNnP1HXeeaqQwTzJ1rgZl8IQb++N8jyAtSgomh/gfytGW4kNAXzX9wUDNteuedrKE49lnruF
OxIohaM6yfI9kYcdog1Li/1AMSEK+p3Mkub5caP7pQdUx3Gk9Y85R9OzCwrq8NUfUX7MwcfTgu5b
2A26PUvkhe1YbKxrG78JBzeOsnX8mavW1UyylRFxVrBVHmHtuayFElr98m+KF54xDuC+jf43+gCJ
k8ND4/UQgVCqiy4ROvximTX2OrbnFay2WOA26iMj6OR0kW2E5bYhsRXj73PlQ4DxaHCZDgpOJ0Hk
CWbo2qBRx8Z87SNDvA9eZhl13JcGFuzecQUocZNzavZGM0ikst9icwYeQeCQRs/+kLy8JqQmhTsw
w0rm73ktV7nzPBHW3WGzdR+7dalYCkSY8nzTGRNuUCTXPoixTBVh95JnZkAttHodwCQdOMZQ6K0W
pf1UZO8kBujujL3meRS5NhP6AqhgNYvHJsITqS0Yrsw25LcxDYxoi/EV1z/iVEAiwxkYDAcLCS8l
wPGUv3qL6gWeeEzBtaYetJabxWvx3ttsZIL4vQzpIokU41twrt4rVhvXDuXfh71Kdmu93hCzFet8
e589HiYJcw1J2Djc/w6MRz6l/dR0xn4KjUH5Lzk6UFdI9fCCJs2TbyVi3Ajz3ueLIExnBQgenxH3
AgWDlt6hCWuT3vu4msLZBOfZO336eL1s0KQFUhcdCTdT6RL7aeLBJjoqW5MG9h41Tb0LotnBAZq2
TeHTK75TEs867NEyGGLw3HNUUUdQlGU+C0XPYvqomL+kZxE3iZLmThNgbFdaM7APLNHvK/f9oUEz
/Hb6a4CfZqVo7LKJE72mEfieSRGgLOs21PePZF/PfuaeAQQE9rrGZRcs2ETp4X+qLiz0ohY2TJzu
v9Rz7g2KSNiKjravNL5FFJcymQBFOjGlEMgnjWbA+0tZ2aUwezK5BCtyNoj+FwrnRiNHNUDtrl6r
DpXYiC+KCMr8r5WMep3NjIE6XS8weK/hbczl6am9YUjRQ42s43kmVCybCcxwJk0W0CPCiqae897h
vrE1dU/FmZ7wRi/14bdVSntp4BTyu1KiqV6OF6WhDWjikkyECf75RZlFG7LahYHKDc5siXrAtsej
I+aOQWfk1Bf3A8ZIwUKyFEwL2oIPdgpOwX8j/eSX44PR2qZmTYEuuWZd+hmYBttxR5bcF/QgCqRC
L2IV/mQjJMxhsEQu/4x48aNoQ9T9rJdZn7elClm7TRVg6vMS4fP/DGJqS64SC36LUK9VeMKiYeZY
2YPratCKeN+2lRj0FXjpGN25GGxmW+rNu8o95U6gwDnUjb9+ZThIzeeREumDib1zsp2jv+D0J2le
5G/CIr5hwnUFjslFTWsuIfe6v5amGgLP9BC7hq33gjSmZPpp/RlnruC5zGYQXO7RDXRmHNwAFDVy
IbxO3Ues/vvhggVUSC8tN6APtuPnXxFhGMyhlIaSSciYxTd7aOjcyDUS0H58ld6cCyvAoPJG1TC9
HiEVVD0Nb5a7BHZi/7jEwYT+0WQn4XUURw5zqW1+RTgoGCcfjhgxy4VN6Db7C6MJHD2jEyjKHLIC
zJN3yDyeGDUZCMCuNZi0ZoF4kdMEZYV9+KzM76r7E1kyCV0yyRamTEuYILhvmJdYF1olmBlmhIB+
n5Vwx8/JXERRQ3hQPE8sckdvBbFI4JjZfXFi/WqRAlEOhZusqtWvihVmpdFzmB/Jl5hFMyg+0faM
I9Z3RRWkewTI1gBszhafLqc2Fi7R4Eek70SLVDUyOQs3uhVL1S9PMG1yA7P3A7gWRBIwazJtpcJB
oxy/0GW1JM781N+AebXQUxrRS829kYOS5dvRmMcC9MCQyRbR7pQk6bZPHKC5Q4MxVv7TD0QxlizR
sCEy/TcNEo+jCb/JvhWXOweT8SkLs4tRTkFbC5nIAQwQVTYBEZT/JyPEro7F/ntp8ScGPWrHQGz2
Sd2YxXl3bjasBPencyr5hu4diGApEHmdII0XIKxJnHKEBcwERGx42D3UE81TeI2oE9ohib/4VCfZ
m5gGPrGAlVDnISWVcgwSWHYm7zAwMWsSUsgH2GX96S32KfMKHvZ+xZsTcXGYMbLzPEXmYaf6gqD7
ixlLlKePB1+E1ONnwRASWjRSV3L/JDx9QhCMqEaZBqLyDrshf08G4baPUHAH5tQj/GCy6S4gRCBT
sYSWhiy0q4eurklKPXk4mZ5mAeCtib9WeJxMdF/zVb7OmKoR2r5rJ6qRtdktN32CpZSV2HkudcNB
jw+xXIsdt7ld0W9p9UcqkhoakZhFLR97yaiOIqz7/pJ6UA+txL7Woo3OiM2/ginzDm/VN3nFF3Mw
dyIdA0Jgmro6KHJNbnJnX3eTv/vER4/Tnh/rPbZLw+w945toeducsFQLgkp5ywWunfQ79MPcKQQR
2TUrCZdL4iQ905fnNXA9zJiKttcNn0jSl+yEM6roX11re76wZCbMhpwnGSsKtSmST2J8aLjbQCJu
b6HXS3xDHnd66BnOrSAaqopM4tVBsnKonecEd1b3XRrj/qYbCsRzSkr2J93IjxIXUUYv1nkioySw
C2TVocLtglRtqSKL0QutphC11u86SiB7vMYjvrBTOj2jX5iWJIODeWzB2kJFBw1xP+gx91p2ELDj
zZgYKEmxLiSK+LaDQe+y4PJknmzPYk8ijP9RgNZkebX89pQp+4gqodrc/3LGqF6ebxWkgZY3xbwQ
QjLUHWkEeLRw7KuBlZSC/EljUYTzmTTNnb9k79kmaw2ZUYdhIgMAUTUrj/ckN3fxVGnF4Q0q0UTj
0c4W6Vz8+TRQvcEGObWVleCDWlBMSS3mhgZ1BBX47govPCOqOoqzQV3E4Sk2Qwggqd3TZF12bjzj
nwlJeu16vNGdQxdmAhIM0aj/XqYxV9PL1rkMlXOVPQgvmp8BU1Qi1L3z5fvKlM7jKXFUx/LFqb+W
R7xzvwSkSTLbbtq2lkpxPymn8IqRzaCCAr+0byZ+mVIVZ8z7iBtquiU5xJN87XyZgdIIuf3wWcpQ
DN9WVaXa5xi2rK8bBGIsp7JilB8plIZPIwHeKjyrzpd++YCKjVbISH9nzHiaEzaApyQ0Uh+/oSfa
2qOZ6GA+1hUA1cHl123q+lqliIWOyMySAdRC+oHqGcQXkrUM7DSPJUuN053TWQ1wJn5BeAqjW4XG
CMA9mGhjIj7vB0f9l3AQgo90OeU2PykjPfzZORxUeC6eBbCbIREzXdPvqIzbEIJM5n4dpc/gOrzd
yp5R7udvVdni3Ngw7ExmZwwzhuwcbGxN7Tk2tEP4JGkJKLkzkHPhuY37Pnnfnzc6P0FYtEKUCwPU
0Amc4CTX/hKQmmXKJPzd+ZcoTqOA0ZRxO9pGbNJ5nklWX7NoA9a8z3ilHryM/AtiRIv4IXx9gJny
dkUs+kLXXF4zXlbgl6grOkjCKbEa4tMVlnaJ4Jq4U8tAuwbP58mG5bCfi8/n59bPu16M5tIKj7PT
eZ0zXNvTfmDhC3KFe4o3rdpIpINC5nD5qSEvYNsGMOqHqN3CtfOHOcy3BHkSNzYTLSOwNy7YLdIX
YI+3mLvoLyCugGZTd7cZ9GDADQVnrKb21K+1YR0xTjq+vOCs9vfYwBkYOdPktMau6AGw5cHCQmsc
XOkCyez3a9Y1UwoG/xqAPz7xddMQkFOIWGhQAaCn1M8eQVbnZupIzAD1qNoqDZC0mi3ht9/gG10g
BUrwUZRe4j+HCcRU8leda9ByQFWerIEog9gWChDU7k43ZS7trM63XJDXuuEQaeYUry3/5aRsMR83
vWp/vTQV0IPmVze0JgM3QBmrySiPdBn4a91uRz7oqv60mypzl15ON4mA6WF73QNVr/1pKtUtRnzi
7wbUlaY9NerhtzZTMXctUTS2PBcI53mx79EtFsTq1lG75ug8ay9pKWbX2dck/1SmiEnr2/3/hi9v
DcxoSetSaMfko66vF2Dk0HuS2WURQYRgTUnaj9dNCo7h/TJxk76uQ0prV8/CHGztW+eZGXsemFwG
foSuVd427T7sQhi3/wtvG+u8LPQaOT5dhfsIr4+1wCTsFVCHqbke6g2OObeQQ2WseH7ITwZoBWZH
/B2LUjmFWDEcM5IOgPaygjjRNnAADvaSACO+9MIaH/1z50yfiGOFy8DP2TgNeIQegAEbcb5d/MjD
j9iBO6Y4mjDyo413wvZtFo+SVnzOGvXUGFEMg/yNXoEpDv8+0DzUe0HXehLpYje59QtWxl5HSnKT
2XXoNsEEEuM5R0c0gxaNLQBM61FU5/BDKum7TPbd2lU+7feNWXbDUpZyq1+nvzAs+pVFAoMhPiti
tLL64Vl5owQ1xTkoO2NrejKDDXgBFIX5kOOrMfuJkbUcg78Sx7/9x6tt3myUbFuR3n2o03Kmpke8
w3jnbVDLDYfk7DLhH3Seb6YrcRWTWW1xDPt6CNaDwz1u9RjhYKbeCjNjohuZW+MxfVZfoXMi5OLj
AOnwBudWG5xwmZ/vcjQYHgR9nprnFHgNEu6vONB/ZAKWsv5Jh6qGuYZpL5htehavkTLEVofr2LTQ
y7UwFU0CSGrdOAi9KGKYErxRsfmQgUSKDcVVMYlI6pt26Pn0bXY3zq82XlJzRtTGz7t5oXiQwNBf
y205kix52B8FHmkCFM3rYMchmImEdF+DcOmalj7W9OXSwg7//pNET1XaYvTVdRvdQVBk724oKRAG
l78NJyjsl/6uhJ3ceLpDhLb4E0gmvErqH4/eVZu/mvEJdnGLYdKJ2r289VeO7KaYgJuDTdZ2lDDI
HL9+ERmHGBXtCVR9P3X76BUDQNqSJ/3fcGQAewUXZJYytwxnO21ooljec5K9bLJoHzYNiH+pUxsM
fRNxLpm3/s7qNYrp5Yfit2805Gu3c5ROBJE///g66pGfnQZNw2AEWmSvBWkHRXOuehbBIURrSlmG
PKbVFRZ49UU3N3P5So9d1plK1dGjQCdDzKGUoogVx1idDwjOuEytcavVYBDsAPSkNK9s6QXLe2I/
43Nxfo4V52xE0lrOA0lIlQ8urbTUkS+MJXbQqIPoHsMHUWmGapOgL7xT7Wtwr4fLJ5bAzwe3aH9S
hfVAlmZGdz8/Gqiy/ZS69zd7+13FqgmeU3yHCEv6Y9H6zZ1kUJhwnPijl2AjchsYhbiSnd28cEU7
hZF3lhQceCB/v3fKuDgYJhvNjz3IEF9QLoOAvboPE68kVlRT/OjmtIO2xHbiFVm+TI0yFtgQqvZA
UKh0tlABoIFnU/BmwXt+cCLu5wqTx3rwgUQKDBkOM5IpUhEZEr3bTJ3TTN1F7tU3uL4vvjekVJoH
NhrDHDs/T7sFlFGQtF/EjE6w2rUzdk+amcGZKCdt1zNEndC89VI79SiQCtwca4fm+7Gz3f9aXu8I
WeTPVLzMZ5f9bwewsiChjqT0UnbkpqYDYzrZX3GVDirVGfKFycaSJyuVAOUxKLmDhVUHOp0Yt0Kh
4uJ4sIXCxqgXZEiTR8hk9JQhePJIuOdvz3kYLqBfM12f+NY+IDp3A68yh4kCRkN41HfK+LJ/dy2u
/fZeilhCebqeNzE7pNU5QmcyxSKBk0zyaoVc3QmUCAsM2A0jNmyjpKZoObunuh43+gM3A75bzwmm
wFobf/gbrJIfMAF8YmHqkMgDfhvvceT3+srT+caUWd9wy7um673D1MzRKwLd/QZdsYGotRlYgItz
CdH7cg+2PUkIAOps8XUa43dY6CyvgmwZ+Joz8oHydeMCIAQCf+ZYS/yiE9T1aYgmbxJi3lrfkrHz
gtzxkAkluLtHR6Thw/CzEiGXfPHpxhHCfJWgAJpos2HKm6ASf/T/UGlaOoVaw3dZUC6NS1RKMYDV
Q0xSuYid+h4ipeBk51jLEjpfkCWnZk86Ic6eQPOhGf5i4+6xnfVojVgR/ykrDSYaDw19R0sUbzFO
YJJ5NiUEdX+gI4sQO0qnTzGSZotIyNTSa+V/0ttBdh60lMyQLu+cgaEs8jxVrVPItKFEuZABJfHT
DGxuy028Th2gDO4LMnkIZKqPGm5uePaN1aeES8Hp0ji47wG4i6NFI8asqAQodTRe5yCN4e3kObt/
0IMgxJ7vDJKeM+VcBrV0he9am/jefeJqw3eFuNBJbR3x+iInjUTcpY1oRa/q6xQc0nEunp1b8bv3
YSFn2CpI1bwxJxncEI1qZuduTassN67/90sTboZGsHNPKzrhpz2OPtWx6ZBvnlRpAUFG+tckrJXn
ioGVBf4i1i3DU3k9AJqBoe7rGpROiz/B2M0msjKEF61bFLlyz6t8ftuaOsFgtIUbYdLrCvrGlHk9
BDUJ/5P97e2b9QEqnxIppCkIyiHkedSZAzUWGry0Vi3xsQ+KDl53//MwWuZXbIYnYD+iKm7kICPF
mrAhvyAw9CNBkrk8S9rbMQDmAckDlKkK9fmGrVSdZ7YCCc5C+oPKPesEhCiHFcpKfjYJEH2aydm5
oqQNrqYYovb3BHdEFiNakmNqwyx+TBqu+H5iYb6rAyj3wzoBdjIgUxVELx20I5NB+lnf+Czrx+Px
gimzJIuH2DCxWRZz2/LEalrBNwEVJNaSaA1ji0XW8Bzl9aqTYw/LAucYKxNMj6rhUSZvn8dKLkp4
ouioC0EJ/oyZLu4c0qaFJ+Mn/q2i9Sis0Acnwx5UJ2WGb7Ve+zVmwwjgTi2GVuV/UAHwKUQu6qGy
UrxESAJNpKgwItn0HL1knQ4Lgv6ZDu6/VwVcSEi0fpEWVWg/k7Mj48yjou5pN+pkfBJLazM+GRIY
LwfI4TxHSA6bHQKHCBZ3e7KqetMYtD53e91tQzuu00YMpfwHbpqDXcCDo3uK66Thfv8dUfuk6ora
RB+XA1ri6+MuH07Qr10Z13UXCc4QOmsGSm6uPPVeQPk7kybYF4Xv7RdhyivENQE6SpSlbVD1Iu64
k1zBaMWTwSkBZGa1m5IZzruybCxIJVk0ulSbD7msVC2qrKpEmAggcWVlJctiCWAN0OkucN9QS3fx
BOmgT1HtYGphzgTc5+Ic3qSFCcVv6FopMj9PkdKex+IFiTDNadjA5wDQfU/61uX2xT1fHjd3n7Da
tJN5scNmXjSOo1WhM6J3IG0wsRNY2U0hCzoZHxNcURc49xumghyyXPIIgGbMHWVZI+dXRdzj611e
zHzF8p1XujkjUVA/zCI0wRt+vfCMHXpU36aJiGVbuCkJxdI5M+13sWlpYBVv+mRdJeSQvsscBr2L
TAm45fuGHXdJMms9foqQy5MmPiapvB56dODruNA2IjQzVbFkf69mjmEl4FPc4mSgQ5/YTI0enIjO
NnjxAeY1CX8zjkAgX2CGEiPvX0/Qx7ujRMy6nsPYbJ+PmG8ZSIlacAdXm/s6nc8kmoLLn5HtRJIC
GO9D0LL4Mib4+yTLwl9wxZFBEPqOvz7DytZxhodUPRJCW2uWaYP3lCYMvpHwj8RECmjzldawRVRY
9TsefHfN8TKnskNJMcdPXozQPsylnywF4YWs/+gqae+OVsV19uUrTRyEKrXGJhATS+GGaaBbWx9w
YDv5bhBETfefLo4QAm2K3t2sq6OAXR2ksr2cy8gW26/lS9SzfokDjOiMbUNBgqip3qa2RKZKFu2a
ePddIZukkTmlzThlS7rq0qp8r0L6ZlDoxKZ06Ok2w6GPhMAAQEVSLC1u5W+4EKDjNGkjUTyhK0Ip
Pr43f/DaL3J+ZClLVWMZ6T09v1rnK7tzk3oqM6DQel8X1spZf8QACftRD+hshLePJOV9Rbrr+O7j
biDL/wumySwdZ1xDuwO6HogxxX4xYUPZHH7TQasvnZH5M/N8pCWGb2zghlX8E0woq0qkOHV8YfK4
btFZMaNA469c1M6dOqDdaNQTybmOO+EhKONJjQhIUBjYSV9G9sGT4viR7Fjp2WtwKIb47jssIInH
cadjxdUE7FpDQfJtP0C2/UF3CNS8mwk10KIzNbkpaWPyRqIaZ2+fgshxfoADpWBXo00+v2Dyem9m
7yL8Z5zIxGrWO/nmnyvUdgKQNXSEPz6nIFk1VbAofcQ5a8cMQD+Vf4oLvpXSKy1KuPivD7udh/kD
kQuSnpXsZGwtNLRBwH6DDre6hArCP89DnYT57fXREB/DM/Y6vQp6XSVpZgeTkrAzM/oG+Zpd+imY
QB1aU8XJ8D4J/S9uc80I4Wv+IBKmIBwgtQo0oT1WNT0Yw8DpfK5ObgyGzhZY8lSpqjw/atNUzXSO
9ivB4Cx/KQa6XP0/2wpiuAOvg4OzU6SQyWbNnCEQmhCs8ppxQefk3qoahCS+P2XBUIYpkyzhiZZK
zNQpzXub5si9+6j014s74tB031/JK8JIB4a3U8zNWSA3kx1ukbikqVfKcbRtae2sw4mw21amCkMG
RP0maBdr2am5zxYwlGN62n6sfO1kxanywbrMoFMeyygjZCneg8n3Av+Uf00rHD5pg7sV/wOG7Zg0
ORaUBG1BzwxnFNYpmeSTLXfnisBMExEXv97vu3fU0qV8Fsl6oyEzdT3blggSVixh9iI//9U1PSS9
Fo34wltofmMJ730umqag+EYr3km5m198B2tJf2ZjfbGUsWKd73fRoyo3j4HcG6xNYONcx150DHRk
lJl849WLtKz2aKKqU5Nm3kZg3tvXes6PVbW22maU6sj1cmevxceNKL640vL4MCU/mBgPs4EMlvVq
thlU0cyXv/UGEqrMp12o9Adgqyh/rPYy63WP8CDSZYb7JIV0431tJJ5G4eRQEs01V0unZPyOnXd0
P0Ddknf9zSiheTMs+lmbt8QGySVBlSgsYrZlj6s+j9PLZgBCrzwIbCZclMQdZw02RBh3UT/+dnZ5
qddddHG7cxoVPFLv4h98gmQMgdrshywXGksMjj2sDTICNeqjo+TQvo+SR4wr//m+rz4Ime79IqKN
sU/VVjBtVfUcyhAW4UJBeV152RXkHjxDHD2Y21m1c9t+4WrubpF+gZZ5oYueik7tgVMIlrtinXRY
zj0G2uHMR8gnQpL5nPOUoKgeOCnCe0cxm30KPOzInb+BKM4PEKxH5F57WDxeO/1n2bxS5C6eWnI2
SUDYkFCXkZin7h7jKEJuNGxyAr5zGSc2859w8Gj0fq5esGRiZ7yfkAdfLWuGc39TYs6T7JRsSOcQ
K8HG6yCWB7vSSxNUFbF0rKh9Jfju+RLqbltZYWYr5wTcUbUKPzxe1e9IOuvp6XX4FgzggZQYqdy8
2weWb+AhEgvcGEr3XHIlmAYzWX76yFovTnNM6hQ2ESriliuzHhLjvO+75LbMqPz8E9lCTgezE6OB
AkxXuZ07mTX8C6wibq4KMv5/1N0JAB897+7iscmVRetp3u5MlULOvdCC4T13LRH2pA9EeIcupsi0
3+xsaKETM1t+s+tVQIM/VPfYUpSrzfgqRYu91+Y3T1TYtG4AhRCLIZ36PrjlpEF+jQj+8br4ZTPy
+6HGX7w+WwthuDapbv0NqqG87UFJ5RAKLwIjJmSJ0NB3DSG0eL/peO3A2gwAzUnWJsVOyXlakjbL
hr15CiTz9nrbjPJL2fnWRoFgUaH+QVsenBRkGsMrI67dK5uS2vLZd38ncJhlO13euUIdTqk72puu
6w+hNSJA08xDFmE/1I86UwtUumm5kfG1vozt2nnGPNP9j+x13fg/DWvKrMWO0fdVO2NNB6LZdjdb
kZDkPH4Nhy5Pi4R5fCgTVBvKGznbgOUPMfqJcqMuOVS/o6khpeGW1L8fcrKt/Uhpg6DQOVQ/ga92
2RYiC0ov5wHLI+M/9b6xPLw+jIAG4bJMN2RAlSqKxokTQt1gs50jzTkQubRtaeIgbBwjCz6Gl5xw
05X562tNsrthBrW6XTSdVA1kBYiqubPamuD5j38RxpZZFUEAVTBKE7X194vPgsxmgrPXU5W3IsRR
P1lXFX8dlO/jyeMD/TsIxetfzWwgnPFS0ngv+zQ27O1UwiYl0b4oN96iYj+A0mzxbYJeuOCuEUvT
mIsUfIKd6VwM8sXvYqCbY4ibVY4InJmhsCe8AbliVo4S3nl971EamSv66JrsBZCs4s1oLLboq0N3
gqGbWSQLXEuQTGiGZENvvnRfBt9h7G0WuIEEtSRvX/EXwALKe97vY08m83FrBDqSmJ3xsVILDNSg
iN7yalbz4JKMLPaWYwdqAj7MONYw2DtDdc2RtzMYwEEGmj7Td1csycxwM5+S5jwWS05oAiaNCKIG
VeXtvtr74YBGpFnhB033gAWWqvSsuIsXecI2lqxhEokMMZn+9DOsI7plNn4Wd7L49zPLpD32Tu/H
3iU29FUylnx1hjrSwIMcJEBXCwa8pVTo+lDGTYaW22kc3/Jm3s0CGSCvQdD1uXFrLsOnY1f4NaED
AoDf75ERDKmQl5C0mfWP6ZwwAfO8es0KotAB2qe73R3VDl30l5k2wqJg5lGjpUXCbatxBNlDZQAW
ukENcqWIIk9s6hXi0uehM8vSFT2sSef64ej5AwVUvByYs5VppeYZIZ+RfNJdW8UQyULUQnC9JvDn
xcQguCXLPOqM2w4ZsJR48ptR2JjQYoeMm2udxc/UYJ+ik7YQsrcS/sx/HYCFfVTcbFfXBxGp+cBY
+mbqBqUeR0XOn2wYZcwQ+XO4mgXNveLZmWmkSqDKC0wzo9rHDxapmCWPbXqPYYzx1Uua/02UV8iO
9PmH7QePugC3QFHht75gKSPeSsVY6rT5J+14ZgTHbiAhE4ARKpwwXT0O3jEIANMsC/gS1x64Q69g
MJGPzFzseZDgDq0cq+wTcOjb6EcdchDEnmvpRkkyjweJB9G7ozQnmz92+ujfshUud/0/09QZkzmc
Id5Qw5zZn2A0ANC5ZLuOsjf3UvM2On8lKcVh3lbjXdjIc8vNsNunc41cE53Apc3hT6h+ZlmxTvBq
85zdhhkoWpXViJRi6FCavzbuwL1iIAFOCYjq21YkKPbjdJYqYnzX7a3pDogSZbOF+kKOfJfS6M8h
JjhLJtLPZhzR1CkwTQOB2SxuMtGmkmKp6d+fw+8bVzzWi9qTsX7Wc4OKpLHrOj4S97O+snBmPJXE
PJpITtGS35+GDbjpEdn0sd+4EE5wvwktjUjCIi252jZ5cBcduRJio9gOVnUL5knp7LfOUKVJbLD0
B84T41dDdBiJrT/XmvdwPtqvP7wQPzCp+P8GYsd87WmT39dqLdro7OFV2GL1q9Bgw70ZezCTYp5Z
Qtww16Wjjnvhl/fPDhDb0GFFlmjxc7jL7rNssLpFKk0XlkxpqUU3Kd54blxDpDyRpA8ZVPPq1+W6
6XsNEqxUVKcnLhI7tQouiu/pPQlf1BScA5dBWUeBSV3sGASb4O6l0KcvgZPwME5dFrmmUjME221g
3orvUSqAkTGXr6S8fU08C8OUNU98+jJjzX5fwAPMDwq7vzEMxZ5+F/+AWM38AjswJTxp7KpTAD7v
cKeVmlmEy6hZ7uxdQupUvzxO+k4Ch1VALZ0sXiFkyGjt7Ibe9YXgGohaa25j77oIbGtSj00Nrkts
LWrGTdnYGXCmNbMPjS2GERaYT4WGkjsRd1Pi0IOncG8fD/VeNzPVRwiyFsNQemAlOBpT+4LaxZhR
3DODWFj8iIgFihEzHmAQAJ/XhrUa/31rpEwXblvYXuVVvFNm8bJwW7uJ7ubp0AGudVRqghs5q5IJ
TCXSouR9NzwMnUIGF+DR7I9TgjMol57eneMoW8EtJY0zkhDMRTtYg2WAWZQlI5DKiqTxvz5krqlm
1P+Mdkqj8wugQqZna+5/z5nQuivmQQ7naEydt25wMecUCuBj+ZIMJixeVGAyGrrJ1UsBAJh3HqoB
Kqes8Ub93hicdnA/EYyF8g30cqEjOxwdn2rW0IMzAIeAkmM4UedYW4UELckkb6yoy2KFMwSc2kZD
c6W3qLavBfzQVc/LATY48CDFGCynQ14zqvQVqE6YVXVgYeSo7VmAp3XSwd2Tv19VxabMzDZguXE5
0jQKUgVrdJ6hllTP0VoLkKsUHpBUXE9gbwJqO5KyS5c+fdfnvngufn2bHUejTFDEErehGgA4sms8
Y8a6REj3pasTOXYBJ3FYhuvqBpAXcg9I3OCr3wCfVAwV3Z9TseD11UCHVTbiSA9ggspsPT+i3BjN
Laf+pLCZ496J8EM6lNB72IAG0PTrVYiQE4Q0DIzCNnM7esBY0RcmTz+nHevSEVywASrVoe5aYrC2
hD1UABiQ3/5czuszxnXTvOOhbnsMKfk3WcKrpLSCvBbiKfz98pRCqrt4xGgnwfa6hMd3mhfcGb4z
zfE5z9SmjMBPDU2nmOXtxWx+YavEILB6cLQhfpWr1SLdv7hq+d15xwUZFe0GaFUasdej/nPz2L6Y
Pko2alAnZJQXXesaNu7aX5GySPg9gfSPU86fb6AGm02q2HW8Nr0LwCwIJfcmb/oyL6EHdK8FsQKm
Zu0bsL+rDk2Wx/6nRk0dyTUc8mCKGJvIo8UeopSzzYwCiczyn32K3RKOBRjrpZyvezXm0jLgnaUf
ZgWEFJOVbaIF4osBfts0cgtx7a8W3PjcvfTVKtqa/rtdDp4E0wNku5Nomex1h/HsKbb3hnf7SEZw
oFWLob4jmdBBPwuR0EyWvQdBqOR7hrut2TI7XzYvQQrmiabrwqq4FKc3lkSHESWqp7XLzWHZt1h4
59ft2A19LBPkhvtTC3zriw/nAoTO2XIYnuSC8UkVtMgOJIiZ9QXcMA89lerf6Oq6nr3/h1/rsv0p
CozzdxXW7jPVXPwzXizX4tF5+VPdJxMTwya4sYtvpcDXud5jNapx4WjUqYFecD5ISTz/AsSyTUIV
yyK0m45q5pGf9GJQepxj7W8PsDsdBNmQ/A5HeCVr5Fx52UrMj0GJs8wcUBtvRpjsjUkv63JSnjLI
ZZO12HZkgohrzPMntxkwj1hpMLE+YBc5ZSSm0/wHwYEX6r/pSY8Gfhsyg6YGbnhAvhRxL7+amT1p
JI75a3grk1mOM2+YFDMXI9SjwwRqj5+Csl8/el/82fxoQyabruRGuWO4d9Il76ctwjS7xERaxJ13
mVyYjdcF1x5eK0QppAWFVW1rp8xSICb9EAfhvUxRwXSZ7sVaq0kcQuvNf475XuWyQIqHIbXPRQox
qBi57hI8dLMTyhWENi7XlNDLSQl8Vluc+wAcnpcN2ZRnNum4AASD7qSluNz3t/M1L/0Zm3eXy4aC
NU7KrixdkVoFoTjSB9xU+djqKQdxLWvW2MZPkQvpN1WiiwLpAj3XX0Iq/Cv6yJDDaemXQGKQacxy
wyedNZ7YdQzHLJvy/KHnwKFO/UiM9oyKoqcagOGc3qCtDI9NpYefuABD95Gz83c/4yguj063DbdH
xaj419c2TJd3S0O2b+M1/pW4Gt/30shwRgKAOLADy2beQ1l4k0MCWSTSFNqd/KpmzhDu3aJpAGOB
CB2kXgrcAvdqhPq3IY+Uv4+/PyFvVDi4OUHr6JK8b19rSBCjrnCAyfZOH+c4ukUSMnmB+mLPBdt5
W5RIwtBdnJKeMXw99NlTOHbfFiPA9enrHPjiL0m3hf/WbCZSZHS7oHJMhdITFN8M3xdYQWtESAy9
aJXGrTgyaZ5V06G8gu6ttCm3fT4UorvAUSFaSVWj9UwZ4WOWgsP38sR8WU3RwwwxqIGqKfNumSb9
JExEBBz7pvIAzoratqy8cIxTH35kO6VSUvELU+K6+xs5AXDUNkQ7PuypTogjIpl0TeMAX4FC+FN7
M9oBblOTNRDMSFrL580ecGMaH4oSFmLLjd4Cv1PX1skzWj55f6SK5dWu0XdvfjSshDL59lw6ddAD
so1fEL6bLqptifO+uQhQ3ntX8LemAemur79PUMQVBpQfUXcdlugU6TqOLPrnPi4ltqrW/sRAJVqy
W7av16XXLKYSc9K3qShuRHsHsazFskbjKXMHjI/VnwWYTTpfeHbW+Icc3EpipNzTpdtqs6lRTvkh
lBAA3e4wEWvEJlA3VkeLAJgdntS2WaLDeREz8rvVDuQ1bIc9Z0ZiHFhFRatj1dUhLZWtzRqPq6yK
rIwafmuHmQM9DXttYodGZBDeLgHKxWwrlHd3BH95A8R8BjC0FOMXAiCTEnTtQa9m20+jDdMZdrUP
LlysRnC2cwYhOmr+vK9vztb0N5i6k1j0dkS91M6nDKOv4xg7CYnhqNJv0Y6Jg75DjEChz89OUrws
QSqs4xL+T3yR5Q7NoSuu3XGt+MfZgh70+bO/pGbyg9JbWaxEjaPQPffq5VLOuDmvPA+l+ZIH0bsr
e3T43raH6vbTKolpSo2cdRbhpKoAu+zoKnHbdk1s5Iwkg3b7L0CGATOtJrJUxHn0lgOC+zNhWAwy
ujsTQJP1t8Uwzg5dtPMq7LXfgavfmjhceh6LYgNsw8o0zhQInn0YDnL8++DtYTc3c7EVaFRLhbCF
Xf44a19R/4rJmjf1mZ4ohrzq9yabUUQfYI8aQSpxsmaJDl4NZpH5bzwUyDrPsSzZRjPYgpbsGzuV
hXXDGqNmwom+jQyUvrIS0Woh6JhCPq/+jgkifDSdrZCooaKxvx5tdHkXB02NaOmu1cuAyxJ3EACi
UEQhWIbzuhulsmZaeUJMTydQjffkHda74M4xl5ovRxjFSIsGAdwJd0KD4hqbv2kkrGyRLXOgdH4x
UEeR4AsXxULgBoL1LarHgLc0O4Ip0vRBR9ibYeWOIvgVQiqnqIuGGFbTY51JrsF5VwV4PbVihyGi
nHUr+EjuLGI3jAcxjnRCGJGjVn/VD8KvVbL21Ots/cFoI3N+UTmS/mjVn5GOgekeN0Fb0CdqSSUW
Re8qIwULN59kiUfbnpN7tk8AVZ5Ekguy3IRnBtxylMXecVyBDB3/gBooKD0ILTIDdetY2UN16mPs
MPdsZj2c94XfYmnN5bAucrtQ8ccgS5ItZzsMds8v+EqertwiiJedPQcBvJUm2KduGomVLa/EX2zu
mF/5VovG7mG7lwWMOvm7BTMIco3xDchhmapSGyyU9zBAjF/6o9Ln4hy0BopFhoLeeFofuiIzjfja
4OwFeZ57NnVpWwQI+9TD251HC0X+BlCjXlIlr7MsFyfNLVZt4haTZDl58/k+9zAKpthbR8DqWNZJ
NALj6uDgIwzfRO5vQqrk7c1naJyKgVc4iTZhTg3GDyzFP28pBewzxYPoDLopnZcaLFbBRZqizJ3A
eMLgi6Ek3f9Uu16pJQgVF213Vt9PhPHeZa8wjYKekAgKORkLtHkzMKWC18JOpq/gVewAzrsr1pjJ
b0bME+4czjZSFOfhimVKuDU5FHIzTUq96VbwtklXt0L5Q1l5hZLR/SVglTmNnmdm5rw1wNDjqLjR
mFewbIr5WiHvCiwBweZo8mzik36CSJYLotdPayKXPY/qsDzF5lo1NSJNsMV8SiumYotuFGHrVYN4
02VBfUhdKwVVzBUgD2evvxSCSYS7Tj3RPuJHerzoYMlJ2+E6XGB5vv0cTCpGBmPwOFxOWWLSBnak
Ek8qhtc6RqlP+Z5MEoHnL8JG0FNIZV7ToAJ21cP7S5F7DIY9V8U9ZMNuSwJh5fL+bneRPKxszJB2
6ZLKvSY10ZKPHkVEkA95ENDm7gQpu3usGaSYpBarDEY6PQNkUM8e7HNAaHCW8Ic2kdZljteyp5Lj
qhnshJxsw+09ymcfvaoBHvL7+5rO6EciqxQKilbHN1w7LmzfHW44zVLLIMti5mMi7krb9ontubZZ
LhnX6h5EFwcdMxqnxAMYc7ypa1U6qrNGTeNng6hjHpO+bH0P3ioSIcuIQpuNC7ib8BSKG6wbEly5
XJl9geN0CruGgge8z6xXV0DrU3MfJp3PruktiOGqBfZrtwG9JSYIw79ACcpHzBLev4UVO+MgnmlZ
fECnDCUnawfqGwob0AlT/9IUY6Mr7x0PCCxBm4rAF2C9G3gaMQeM2U4WCvd+KdMFx6m/9eN8gOF1
TBlOrgt5E9t5gjCc5zWR9/6Bmw7+zF0KB5ilO5oB5XAKWfWhIFb6vzc/Ucn//fB2yJ77P2eCwHfU
En9zKIWiob1CbbF+eywtdpv0mgMT9YzYC31YyC3rRViBEV2zCvxC+G21IyrkLE7Chf6RBHxTlySM
JJ+oYOsynDvuzIO9I+JOXWNVEbbZ5/QzrBO3n+Css8HONT2dduKVgLthGBsKtPoopJQjgiew7BJf
9F9x+IvbVtexZ+AcpS266jb2m09xLq39lVYjsljDSGuLTmjI6m8qEkjJZIkouKLcL3SoTfVLD8t3
L8AgnAzDRLoes5Mr1I7H8sTP0SF+p2DDASPKPtwbcI21RxJ0MpJfMU2WBjImfWcsSxnntin+Uwum
SdtLLPZyU9iVnVtPuiEPNgTUnyscTrn9tjmwPbvLJy3LrC6HMn26H6QnYUOu6lwcK9seYDTzVS/6
H8RP4SZt5vr7Sf4e26PLaBfQoqeX4B6ZNTfqft1n2k/m4txz3s8XJDny5iR6Yr9yEpAl+a9Jugj4
h8VKlD2FUPSwOCX39lf9mH4zggl4oSHbc8Vt9zEaBUKXb8u2sCAwW1sbv1cipmbg2WF6Vfe56qVR
S2QddhiwgnQVw3UwTJZBlK8szoXHKafq7vJedtI+x84gKVCP424zC2J44PFqYlfzGdYCYUlsQQb9
Xau3Ig+utzDLJtHST+mnCRGGqhcLFq9/A2vwIwjEyeLkpR6dNScC4xWb2tNEZrUfRHaL6ZfruqQK
dxR+n3Ud2GuYrNertChA7O3u/W2Kvw0LSKuCvtEhZJOKS/lMP6yBFvqq49peg7zMBt9pLg0j078G
1LTrT561JFMPx3f/QVF41LA21r8ckMWsBklVTKe8r2RDXlb0y3NblCgXebAwKEsOEv61toT2n5Z7
b8dKFMOJSMpe2u/pye0Z4cPj8anZhjlh6uxc4MLDlut+8i4bWgzvdmg/2wMwrRpHMFz0rkvrBKij
F3IqicNwuTBSa6wUV2r1018Wuwj+wBzlhSU4QYHCsVMNreX8hkR2Z6VPC0Gfi+v0RS+T+HgpXLKF
jjDzRukQgW63ZuCfMnYdstBOAbn1KrKIEBpBuK3Gfzd7itAgrNqrDwraVx+l7b7oMHmx0l694UI2
mk58lkpnlxkz71hbJIs7L7LBKsX660LzqpEZQqvE8ORqjgz4Aw3aV2OwApKTIaMJubCRA1QVxFD+
/f6QtiksjJkuOCNr7JTiCvVCavhRvUegx+dQkJSfHiv3ZYjLAhyyl2ofdncJh4USddwELifQeWee
k+BRHK3BnXlJyMZp82upkpCadsw119xu7DjC7bgtnR5Ql1mAHHLt9gKuYTY4W3vvT0bLhGF/Tf7V
yUT8ncdJEvne63TssDXWgTqpIPibKZ8OWYWjGopyntLioH7D7jBP3OxutEFMrW+p7pCbpYSt6U2o
t2Lt8nhl2BvLvtp5KRn23ogfqE9kyGOKmFoWz2jA0vGDdjgHJwyQ4jQBDs3fWiMdfScvqfVmUVWj
Nz9vOLkmM8fLUf/y6yzG57DcpM7HLQhjAfyC9r7tgEyqYs5/gzoe5+2K8NHVs4WLtoPT1hlF0Do9
gPCRUDY1/pBn5EqNJoP/NFdy0McKVDIGgQweR3t2nYJ48YG4tJhea7wbRbUqw7LiNVaaKSo0sNB8
R4F+EguMWdidb/SnbEaFxCGoZW2qleVv+DwkHAT2WCFuWJoG6RCBzMWFHckzi9dyUz7TvTSb1VAh
6aK6Mmr9vQo5Cex+7QJP2dThLLxAelsTgTMRpfa/QD/hVcQa6gz7vVrHWbBiqqO9GUeDCninRsuY
iyIivtJd2FdqYt5/U622DqCgknKmTerV3jNsffbLxuuCJH89WHq4f1d6JorQPT3QnGjjUga2DeQz
rD61mKIzB+YKPbf6U9oKtBn8sRCePuySHTA44PRS4yQ3d/8Phx6j3UmsO1wP/MiYjOLq0/T38F0I
aM5X2cErHRZ2+GyP1hzVgK48CSc9m4Z0YTtr9y5nFwHxjcWau8dUi41YWHIIdwvzGM6KMxn6d8GU
YY7I/BX1YCNf+6G0PiDjzQ6ABWPWn4VEDmbw3KGXMTAY358TVtGP/iP3KNKk5xt3BQDllZCMt2qA
QFWMQBLjpZTSZVaO1cEwV9mYecGNaynpI42dEu7qkAePLe4UFraiuMiyixwnHjKKHdaLn/2bEyWo
XOqbDTpX/jTCFbWvMMmtq+es/r+M1pjbinyZtVxdxgUvt5P5TgfUKZZg/AHS7Zd6Hpn2g+/0LJnJ
QRQzi0cip4WUs+7o6797WIO9tcKVQSVz2xundsvhwTYnQF1GS4udzd/NTawPq4uZMkAbf/LCLcpM
flxQkTUCGa1KCgFj9bEhX/7+rzJNXXk83K3mKj5qSKMEbWGpRGyk17DA1U8GvVmT5jUIi78QgtbE
DGu0HmuI8qyN2HwF3J5rKmRamfEbezxkBO6m+Or/FUNVpe8P4vomFtyQcr/3FaHELQMNN8P7VKDD
p35hXdwvmekMwznhs4EqwrBbrH0VzBOATBB1lsxQCyroUWk0L9QQndS7M6nigKmOzpQ6EtE0zu4M
SPSGE8UpEbO254kiAhqT08QkO82mcB9qZ+CtBZ+X0s3bvDheltXSiN7pg2fDSyDq+tKZRfPXHQl7
b38cXPhpUqt5wDYxFxVni+TvBrKJcOJBmP8pFh8B94IwmOW6cPCdoWh+N+OUdsIT+6TpB1ROVO+H
9+xVAlAo6rIyOdaNiqnEQSTGb7R5qXCc3heltFkILK3e1UXVpSWGr0ifosdLHXBPDXh5KHw8JfNM
tACqL/V3Rpeng1atC4YDu6t5NtvSVaZ0UznBYl8Mu4whX4oTBbv1vqm3WlC5aZgtU3RxKdTUeN7u
5C6GwT+FvTJp+cynpSsxqMtwS7iEW2cEjRZAhMVvrqtLwZKnF6jS6ILtK3Vd2uftoPqreXLkeVuo
VqmCk5ucMiBidXM2ugUm38AFAbNoXyNWBuqGtFfdQNkn5mYD5Ph/5exx2pecbJfNKHtJxxwgNxeM
m0e0NYPvwqZbdVgkkuI21Ip+bJK7WByxNw+PnDfJU7YN+BPex+XfJqd+k32KbZGJRpWGTUcoGQiZ
p9td+W8yjID0LLk8mOhBXnfTkYFEfOZNm3MtnNYeIoS44ntDIh7A5pN9kTnrYqklT3WrjpzVrfmE
OvDNNjFXdyojpOdx+Yw75YUTRvb/A3iu8fOyhW0oqKFG2ML/xSDKwLNUPqEE512kkErrk5IZLzr/
WG4dhuxVmR5PntsC8rSduVtAzYIlXPV6lTkm3d1mmvYE/mLPmPq99GzCHEyDAZmjfzRvKU6vurNU
L10wrekmcrsRm/ck4y+6FCBnxbs4VIRn3iu5k5qAJO2iTvcub4mt9ffbvh5r1CChavIQJON6G7R9
0/fO5OuTH8yepkbtuLaSlM6dieTSaIXcABGYppZniVUDGU/b8qZQzr2FIClU9Ueb4CRM/x5w5oj9
CWejJWzJBvAITfMJEZAa+c3LEswHiyDC1tMpUcRazvbt5sz6DEiVnWeeU+UGN3bdMG1MWDk2pja0
3789MqTt0unzPmINDvjkrXs/TaP60bkbfKt4zDi7HT0levWc1kx27SPws9vUPkuLPj1I2OWpmq5m
g19KM67JM1qjSUZXfou50kHq4bHWfGuInAJwbBSAF6qJMI56y5b5a5IDWVlxnJED7ran06l2Cg1U
yUGIwxi1tvJZgxj3SeloOa5+SQ28XnJnJHcg73c+0rGXPG2y6LV/owV2OMDlOTkqE2i9ktZ5sW/p
6zI3g/D7QmmrU4uC3swqferdEHuYWf17HGNXWHVVbv9V6kICuv+nPl1LUmeM+RoSrMyvndQpVgcq
ocD35yif/k74Jp1IfF8ts4X7wC/1r0E7ePJN3g73dIjLxR/k68fw4ZWgxVKIiGX2nZXF6pjPEjs/
j4cZObJI5baIuqIlepEsNIehG6Pn0CAe/QfXkAh8mHs49In84nKn9uqZtaw/itMX8n1GNkMJQM6m
RBawRNBTAZJBgPe4HBsCWFrHmhHsCuz76ca6MqJ9b3RuUbvcnFA06MrMYrmm/3kepnGaNlyQbTPD
ALRywpdMV9nSN+sXXFniWM9Q5Q54ok+DpeAIkGkaiLXpvl1BZF6Apv9IHzFWQf2XMzdT2Bzq3Ak1
G93JBxYIjswxSrBqPyzMIfWk3J1Qa1rUD200X0sHi3it7SnyX5WIw0QfVb0ZiTSvFPsLlwm6uIuj
su4u0tlDSk41TzwOFcnBWi9pQjEYNwPhkVoaK2raOxm3jylKgEtVKYI+1yztq+TA9u2jjA9sgdv6
PhXfNnqXrpwOlSEClVvzvwT8wkm2H1DvHFmvyyu7bKaqBC5fWDpc+0c9bHmbQbTVVlPrZPOfcLp3
GrD///KEepWANZXVlOsQ/GqD/UmT1dmp31fvumQFyak+nYHrQ76p5tMrr8hWfuNinJ4tOKKtVue5
R3RnLmYPzBqTxfS5brFkkGfbEiZGlDEI9TKq/Ww97sJzwk2MbMfKqJTg9S/tV+PlH+czac5uROtB
DyeFxevRnXfciSTwKfQGiwTcwkSU/CaspCX3lEFM1YBOyJkMwd9EJqmJB98Zpagbxth0XCfIsBIZ
G+PpIijPLYkg7R2CC+WE2lqO3YxSZODXVLl4GzJ3buTvbgU8IE1jNUFiYVX4ewY3CyhKNqObcnlH
pd5ZSRbDAQz+LCTzwsW9xUlYQCC22ODH51PuewthnpGlnbPZDOTb3sj1XxBCKuVg4C3oaqEUERuc
aFKgqhtBGPsjEWCAY0BMBMKplbVBenWZkoimGnRMccWg6JRKuodc2rupIWBCzMeRcP0DtY9NTyHu
ygCZWpGiwc4AaOOpJkmZPIZLHv5zHs1dJcpmQN5uTE2nz+9ZkGmlTXk8/oBjDRv88Z7o9jvPNcS/
OeLHexaWtWpfiq1tYd+3rfED+bslU+qwXG54mUHci1iK/XWaI0nFZJBjkssHaG7+WBeSksxZIQfW
5WNnwGuo9ZzBZdqNh7Irw6XdehOEDWLsZdCe/UzOBDKwvxcR8OlLu95TGpjpJjLnQPGRX9tnUW9q
fX+w57k0E0eX2xQA77zU27CsybZ8kRF7/D+SEwbW+ALvkaNDNb8wtqmGmvSmPseXwXpwi10SPH8h
TGjIDkkiI6ttL+S1ljSZvNu/dPv19Shc4wgAuwIGd0epLKb70TP0V0Cn1PpO4NvFtxLOkSmjYjqE
RJ433IiDeVTOvluTxYU5Mr1KjU67Qwa4kWmoDtEbBILNH8SDQ7mBfQCaY695IFkJir/1e6rd8ubW
Uyvu1yMk12fhmf4vbHPMGTM2Zn4hVPuhFuKDwZr5p4bLkxHlSlk2pOOQg0rz7XHECDP2rfklYL0k
soZZaMCEz97/hRo/sTjjW5WUqdlaG7mBFUnuhryCMQkjFiq1hLC8W/ZIDiqu0bsj06bqFuu/H94a
FPjjgoeLCTPQSMAt2Ge0P2KIfhDExagR8adgLUF7UFIB3KRnVYAJ4Ja7XrIdqAwiY3Np5MY73/YL
Z8fbwZa5e8a4wnTyf0ChumJCj+ReMAOe9aZi0vH2tAJS2RrpqjqhCbOX1Q1N5B9JCIH5Q9jMatK1
9mRmyONJAqVIApMXk49nyP6Dsyt0pY+5mwlhWBvl/6AfNhIBlPLNO5l9YHM1LmJMrjDSOOcle3i7
8j5PPOA5M9dFTzIjrHsX5ioOIW+FTJiWJ0f6BU1qVIqwcbK4iiJlTWOC5JSLTRY1jMGbl7ickMUL
jQXzdl4qZ6M1weaf2om8xTCqBP48sqmYRTboKdBwe9Dmajw5JZpXWP4kfwwmi2af/68e0ZvnRtr0
EmkgHwzoiVm+2ahQuUQbnxquWvlzwq5oe5LD1KeqMGnb2CHgdHKktv3jhH1HqSjk55MBbFKdOVuH
qBanGSyLQVuyM8vWz/zM1a0P18McLAreDAFiFHWHHtU5GWjQoHxm7lgIlKDGZjPTf9p8hMKqqcEx
y4SFjvbOxL07/Xf+2EbsEXXuB/VbpshFf9XA7hVftjDSfdiLUf/Zjz6nAYv17Ncr7qb0SxItswNT
Oq9kqEXHxxJDMY143zhWBZ5nfJNXeFeiaLCi1N5NheUSv9xuagbDi9v0oOErBGgu7ohwZM2zvRhr
9jbyEkEPTffWQXsctL3ARxUx9zeqcBhUrKW/rBEtKcWoKPB5kQym0OJ0lco4fx+G6VopeHC4FvrW
PTXqUDs70vW9Tdfq3QBqY62QIBpv67iuKtpCO08+sNeeMPug0CUYlpQHNG2rqkCUr4ykdzlMNYos
244kmQ+4bKX4v+y4BOR5Of1JL7M+Kok0KARSN8rnITKA4kAvfm50fWoAjEC/LMCmFKhiUEwogoSx
l46mxX9f0Th9SAwGWQAfOwP+0v84SPbbyh63kYgaaaFIFHIupXs7wC43u11GVSNoBEL6qp9rh4Qs
VxFNd7k8D8ifQvZcLnHraEJbcwmPR2o1wHUzeo5+qq4f9+KrUVwopnBkVRQ2E3NdfcmEqtUiKykg
ElU8v/AuuAJpTzJrsWGP0kAuuy9Shko3chfTO0DJgFuw39J0M3VO/SEzDwaV9wN3LMyI4FSXN/1c
SjHIO+rA95sOKbEn9KNua5WKK3MSCzA6GlPVUcBodLOc7pYGVizydxGlJdhVdsFGkm8m03Q5/nmK
ndXLKlpa9jrLVqtNJdiygoLv5K3Oymc7T0+8Ch6fRji5ScimWUPfc2GT0g97klxbk+MfzsRkAd/u
oRmbeZvfdMz8yZeJoqo27XWDSoql44oqPiLfDebpWoLp+/kux6P6SnOvLLNdvFaywwk+6mjL3U2K
v1aNRDloZJJXOtvLMV4N70NU1wMaq1+T8LljZXHTWUtY/12+WmvwFpIdHoKuUfaoxyOIEkzcRFhS
P48bdZS/JafphV3YawDeoE20CU9fGKHkJv0DOjqBjgT3X+5lNKHqntRMf5sMuc8YnaHBlynoUMA9
RiAkdzjFjcgzfGwmJzWv0eZaeckH2XxLBJ9kyZIeXQKJeSisMVStWOh/+owKUgU54gwBgqYm1fjn
raTnVOwrmtgh2+vZZqOlnc7ayTuSakM2itZKUrjsLjHU6TmOBjevkHoKOM/NOni6WHJHIHmiEArv
1FNO7eS42JAPp1n4OqiIaKugPp1SmrEsqGG8GcpKmjqqRReqq2KvbBhrkIxlqpJ/fimTcwFIS7Bh
g42gZKGn1Fyv2NVPm16xnfKTbF69Bbv3/uFH4aC63wGHewt5KECkNKQo09S5ccTFfyeXFVhuTujq
2anlv2s2HL5AWFI5QTCxU2mYLjaBlb/MMX836U+CR0+Og/2p7dvDvUtAWqpTg5mnguVNhuMHgWxK
b3NV2yUQgHnNvJjiNK5JarXQ52b1u6KkoQCPbK1SynVKHU5Kbz8Z2Eeg2G4quzdmTTmEUcw7rv/J
vzuiAB1sL9bHcjhb77EoCx3B7BtO2AFPUDNi8vtdJANim0CTfk6UbRR1s4rxA2C2EcqaNlec4bgP
Ff5YRxpLx7HVH9B0fqWAj1ddGQO1cMQz90VhKYyjrnBZyplxDN99hg/FrQFfV3a0hSvyhQ9MObGD
uv17LNZvxAq9YZTGMM7JZ63UaQFEbucaBZ6S6+ZXpTqUlGLqgiAf5OYD0Umzrud0A9LRGs9u4pd/
WPj2Znip0XxhTR9QNgwtXYNP9v1/1vYZ+S1BsI2fBISfypfcahxYgXjXfNIswWpuj64adTFOGpc7
EWjzDdML4LmUQAE2rSghMJ4c5d5UISh3i875G0w1e+4imsSXchIRURbuTRM1GCggSstO9t09meKh
zph3puBU4fK+Rl/jL8F4MqDoQJsp+AnFy1qNd7uvRwZ838RwkYHcWFP/WLb3qhVC9bGAXkrxLugt
Y1LqUTUDf4GXhySR4MPGNgpxs0t1/C0xC1u/ZH8Ck6ZyEH6Md+ZB9i0oIV1vxWfrKo/dNkdCp53N
W9SqkmjCSITtBH6N2eAjWcWVGg1M5hWuEWg/EMkZPTZr/lJX3N1S/UCRLah+aJbBo2cJHFXaSuEz
cexgQN6f31mJCp9sXW++sGICOeB4d7hW7tvDUEBUqrOrDLps5rXynV7LnGhecqbUrM2OWxGqgCQo
4rlrOLpFM6mar/eyfzc/FHqGQDkQClDxllc6UNs4EI00iPitqibZZwqTxhDTNK59xk/g3u3c6HuR
nbz4tmcCvg+6tGGkw/2P76oYU8386OWcpAf7QLZo6kqCHpfBVo1DlnVRP5bhcl0jv7g4j4Y1oP9q
NXyIEukq6khNaeSgO14pET4F0kgNZK8NavCpRJakAWy7R4T+05VDVCCMn9AjKd98c+/VaA2YJ9wX
BlkdsofC/732DXi8egLbz1BzPGOLSsiLs0cCPdwSJyU4t1zczpCMtpQkZpVJ9Q+lF/CSaxtCvO78
b7qXx6CGTlxYgMfpju/fvbrMI00qFVeK372JQQsVkXShVK6wlgkFlxX5dMTMm0MAhKmQ0/Dooa63
bZjxy6XygQRfe80uaS5oBESQlkm2nWvq2CX7IiD5G8qTDaLni74Vw+bQ4qzi+h+/nLO/f8DDPelM
iWpiCt42dxvWDk95MfN4qtcoUOr1NmB/HmDmx6IP7Qc7WkioONrYMHgcaxv4vXUDmwDpTlMnKO+z
7OvanGne+PltRgHPFLIc/ZkuNd28AEX/KTFr/xui8AdJgyQ1qAC0sYZVsV/5EAEGVambpuYL0GFG
dy9EtAb2EgseUlGks07kJ+n/ztcA+IYRsPz7cyDF2VN60AB3TG9BQ7mWGDjvopxEvYW1ZZzcWG38
XsnagS1Zi1dkJyNlAGCXOCNv//Use3SBvLt3Q0KHnrDu9eSGSoeoOCrvITNF1+VEzqU1Suqy7H/b
cqmRu3OJA6M22n19lv95cd+NmVnOAdcYqTeA1ArOmiqWqv5lh6M+v62SsN8nUgcRwsXVFAqdRNm9
2TYYIIwRywo/WBMoAw70adDaFSBF8TD6hEnmtu4KlanMiyw2BozvWcWtEagVuT64tWbDBIsCUtLE
xrLTj94sPtJrgxtPMP4Hy/hIM7RvJBw+DSYj+4PQLFDloaFBJwvSyurgYNOtQRgD7/8Bw4Y6VZ2L
3rxN1INU9+TEx3g78w4c9bdFGcsJTFn0zMaHtoYtgbQNXvqRkbvlhnGAMz0GbpCZTO6ofYU7+iOn
OegptaXZHodunU/CXDsbOywM4NUyEuag4x/RVfOr5xYKyV2qyGI8/eAedD3lL1mnDsFIXobSFaRv
nVuqBPrd9T0jiztztUoJw5pZf7bVAUxDgE4LbsWOfLm74UmPHSW/kSrVLL+20j2zBSNCVHKY2VEh
+/Ped+o1L6CEm+rlvO5UTvFoh6ePG8IalXWW0kh8ZgC/byNKg7Ndk8m5Vx1izE7tCF5e8cJisYR5
4M2nAZy9F8h9q3eKGDToYQyEJAXvMkjTK0VUDzyglffmcPbz5TWEEoAfREVTKAO2Y9mI18azVyWd
u0iEXNLYGbJ8qjFH1N13plspZ90R+7kHNB8oNZNv9bhEUIDq7L2bivZBzh/hWKRBPtxwRq4/rom1
Oo1ADFQXsdd+P0TXY5LbQHtsvx/h9rxsVzjYYi+CTexDRl9aDJ3UKepZ0CWsk4JE7K5X+1tjM1My
tbf585WK+RpIBXwCoeAZIEeqaiawnr4Z/NPNne/OZ0DFa87Rn+ow0B22HAnpd0k56ur8+oeWFU/F
jx+1ULXAWqokjPWMl+xjtoLZNUfKLZ30OfRAZIb6HbpL/UOaVqJMOq102wViKkJiD9ap74Kn7gCy
txYE3OYSmlvVmK1fSFsBXHceF69MoVhAe4cwJd1xI2tfE0dUel5YHFYXIoWMLAbAZ7HFyCv6Gs9T
ykVjTer5es/s2FRTF0Y5lTzpx4OY0pcfs9LJIY1g4Bo0nVJCB4m9Z7sOZKzGhuP59QiYFUSfXhM3
nAwRr8y+xRs17cJOEDMn5CtxQ/VokloZCvyUVcxSV7LoQHKwMFXAUHK+AH6fkNhnK7D+LlVSEnhb
MVQ55nuoxSUcXRsQbfmDJjUCGtOi9Km+LXYNUyT0cRqxBOrq5U6RLXYin+H5MkbFwD5jRSMBjnw1
N0JBEmPtbnbc6z5fPQXazkXmWmlmleKqnVkLVFVnL4MguHskOaTNItzbV0JVOAh5zsdtyKdD7QqI
XNbwnAYB+emzQ6uWoF6RxpYAptolKEuC8L12Oej4MTTn9oB+n1JUjSwKpxmP8d6CKFLnpaI+wcOl
SNZp8x3WbYJE7HV44z65vfcVReMDifa2xP0zYW7jfxGD1aNPVFPqVAydjUddbHN9GYvkAWkE+sax
DxjnwBZ1hDo9cf/pnQgmqWvfMuuWwPjeoQDuHypJQgkuSpts/bPGIuJDyAHLv8lmFQhGdD4+9vDl
7cmDtL7yLUrFYBUH406PFds2gSuhX8r6B8048Yj6gU1Roj9gzlizwiRWOgXmQl11pQhY1LqcajQO
UL5Hr5NEH8tshLjR61nGd7wF4Ssf9wxKSVMRWFqIAEM8i9viG46EYNM6AXYeZ6hmDtP1qzArzJO1
g0JHccUIhSld3Qy7O9We+0IISRCKT6vZ92QOIj9oGqMY+2XeHV8LsdmZg+V74ywyS1w9Kvj955rs
euJjds37szT8hTZfvwNEMw/Fz/HTKyypEjZaQCXiYbzbFn0AlbQ6rSu8Qg0OuaDKN9rZZQ1RTMQ3
PJPELOLWzafh5cmKkzwxnrWXh0rK1Jihminstpc0F4tYAdX3TlhTDBFhv2EghwjIl8nsciyfRe9g
AeqKRxoUsguxUWAx6cTfBU2ZepD8NE93e0jfRCKXoeoisz2VAbAfWz4lUqJxnnOUzjdXBjXJuZ8i
zdpDCIFPsI+Q3m+XNYpXzxfcsyd5Ow9Xw2dftLRpNHo/KCpCMOKz6E8ofuWEWRft7h/KZ+AB1QNR
rFlwIfBRiAzjYJov10gjk8Mp1cuIhT9fpHwIWUD6MmOke5qEk2wTX2uyq7YuOnGJCvBcoxTwTZJQ
mPqrVeFlbAFyw45G36fgHxIs7v1g1oLXABS3A2n88/ufhbY4QYp3HT4gAuhM+Bp083M6yihXxS5O
igN3wdEcWG3ujOIAvQzp9OkfcUZF0bSYulRH7FZ1rrJoZEqZlvQ9XwOgFpzBQ3J0SQdWZYWJM3W9
qdU891HhsTJlXLP/pAqQ1rhz07XvE8UgfwkUkib5RZ5zHz3tAo55KiA3ydBcAkWk9vN5b46Rkanh
tAr6zRhvLiF+8ntBvPsIOJcuacye4DohdSXg/pqQHAdEHJ4fsvEcCsN0vZiFKvi4KGf2NyPjZNzA
lal++DnvB/5GA6BPcXdZb5Spy22WLSgEpFXomB+cXUF9JueN6UL+VPtlDBosVvq1qI5SiSC7hkHV
V0cRvqk3ald7+tvjgNdoGTzixYj2WsYP2RMTVNTvCiUczJQZw2WtwmxXYROentwDDc3PCMFrAjV8
EdLUse3gd8nq8T6/Ixlv8npabtGqFcmO/u0J5WRax3sinNmhabs4Y4TNMaxp8evH3re9pBl2FJ1v
cj2ymygXDwO2so8uRtAP6yDJodnuK18+wQI6sT7MRUl+CA56R0bf0HTOeNmZPLg/4XJ9Le2bbmfA
vwY9I8mt9tV25HtUZT/DdoM4i8xfahLgBWTkaayle4Hf9yEauKxhJyxXsvxyfwtmzPH1Q6odUzy8
nn0GtsBImQcVj5khAqP/KhhFp07x/KbYPDmKi6XmCOkCxvbrSFVCtTIhpcIhVAaV0JrpPODmaoaq
0IRjhfe3YGlv5VqdyqCw9nttwAxssG7dT3qhGijgjnFkZay6rf0mqkxTNCA11c3xT3XTrp7D7EL4
9LugEyLZs6o8gRgLpidPrKyA/RXrQx6RY0ndBLqf4tKDJ8oo6yL2/yaYhMc2Ieg/OJK9kNKYfpQx
Z6fTjPJBw1hPeXkEExWQnNm14DerNvc08hGMqRHwvigqFHovLIx7n4zZIMj5r5sV9BxEUtftrpOn
znwwMp1poxKGyImFykh1/+L7rqgB+M7hEmoEPIoH7JzdhmU2f3mcSPT7ezmA0HLcqIHE1JLOe7aR
QiB+ruq2F+Km5Q1k4+7vmFF+i3KA1gse6oKccd+OXm+8YS+ijRjibE52XKsCYb8/XtEoyrDVMM2A
VfNrilRS1WRioZ85NbZpG02VUmbtOAjks5No3+Jwx9yL+MX0rmLnK9V96LtXhoOxU7alyjWQpcr6
qeIaFbQnRXMTdMz5mD4yuyJFYFzJTNKOkhUdWzIcmjjIGFEYpvnjaHBw3DjwkYYl8WZVAmwvbHp1
Yqc5LNAB27k+GJfzse7hZHzb7wHiMzcUSdCbHmOh3eP/CQLbnl1eLZAm9zSkZ1rKAZPgTpo9VKhn
hT1knBQbVkjG4R5+RfKtKG7CnPb5kBcpsoMiydm1uw4kCying5qwhK7oobE8u6IgM2Bt8EWO9Sj6
2n5k7qdP2Ic5+azw8fjGDTbyhSTBWCwOIgeaXBbH55KJ460JHVXzmIjgQrL97HEuB0iCV0Y9hh9F
NyKZGz6c82giDMSf/8pzQMNzXOdgg+9p4zdikveeefjA5rK0I+6Io1+jO13bXBRSLsOuCgilg6F4
RJZay6l7oyO6qqmKiqnVId/yDmtnY926msCbaRHO7vo0p7ziQCY31JC4QsXSQoN/rd6QVzKcZGZe
Vd3EukYTYKfiPUg8g70T/AMhtJpPTGLglPoesxtUqKBMEjt9XQKMcHQbE0QGiPUN6vEtt+e5EOmY
qvcUDsAo/JKwuGTsmG0cUKcLvXosum5w8408XenPjHqHf8w5N13YHE92U+llGzEho0GSyNeGGA2T
atdkiiLYHNoKF0kcYm2xhWn3I5M1AjxCZI5Ve4viNet5PW1oAcJSPazPy3Mpb+VtiBmiqwCilNb6
bSsnZK46YsXu9QTSDY2heKu1ML6p+7guqG3WuiZVTDaYqAy6SWFbPFIFMGftErPY1zxN76TEsZFX
AiHbn/Xe6zn3mC/LruegIQW7aiqW/RlbC71TMZ5OGlNMD3R8ms7fRMYDIshaCNWyD+PEnXFOszVl
Dap5tfTmGRMpLLyKlImamkekbAIGQnz7k0nrBSsAz+tdf0tEKLY2cOk55CdUJ86+9nR1yifnRmtF
r/KjPerUTUDB+ZxqrV7JtSNpHT8h7wnS/pEvsdqRxNblk2EAvw7lA14xvlRUc/wACe9yTx64DL6B
8Hwpq76jO97E20rNihkyFyg40PnXUugoIvEdLs46f3wqKwHwiwa8v3q3iX8kfRcvYgvT31w00jNq
KQQO8XGALqHmqwjeG/QpHOgLDybPG9a3u9aWB4G0e7R1yTRuG2UT+IgPAJyWJ0AfOpt/QPxQXeVi
b2FbYWrgabJZOHZ+1/o2rzO84FAaIrPUMfl0cTd13X2rwHBN9ihzQrb0lt3Emz7Dnys7yHCYpS7U
dcbg0Hl1NLPLAB57JVOmNOyKAcKaa0d7x8fz2wOXVzIt005MDosx6nNSPg8Uo7GH/cEVO4mbebAZ
zPGO5VTEqk8eM3toNAeU10jlL3r0uD+WmKlDfmhXmx0dzErU1o/q7LcyKFhiVgBBJsPfT2je+xGi
yCsSeXvRlJU+8WKwDLRZsX8MRBaFUy6UE9cRTiEjC/+NU3oFY+w+zyrmczHtlGLWhiNCaiNZg+Wb
1o9Jw9+ohwOXiJC9EoSQdaaPiV2iTM+mvfFgCsEqiZo/gC2K+YPMDgjAwy8BfgiwNQZ8msmYezD8
AuU2OYX2g4Di46Gj/2/I2er96J95wb3eq30NLBxSKFkC3aqiIjra8rs8SPGZRb05mM/EYIVDeGIH
oEqa2zwD8gckRVq9mKwKLS9ZQXTkWpDPE4gTH1XcqgaV9bsHZNYsT0ojvGf/DX2amrlSMQJgqZLU
JfPTxWJayuMttXGqjzjxIWmS9FIlfGcFFas4vSx3re7aDPcJ7+abYGFR+vf12Gzx/HhO0epm/SgR
+rq+VxanQhJLbloHaSQO5I2A3FiApc8RXzX3Dx/p49+3N89zi54/rIRGnG2uVoUPx1LIC7Q2Fn3q
AvhxVH1YpJk+ymr+Q31YZhHZ2UTozSJ7gyl4HKoLnZlig2xMNw9Bhhhok1MfPv6G9xFY3+PGISE2
ILAOJNh059/im1b7jR1QFwI8YEsDy08Q/hnZ1nnlLxrzQillCsJErR4JBbJBQnLb+dqR8+Od+O6K
/MsE+edEdVtHt+3E3eJO8BKeufAApp1z9SPNzeErzyBpZMrmrG2k488mF00KQLYJSdZsy3G7tjbz
pl7OeDI/itcrci0VtBmMpTdjmgVwQJzZtW+F9493NWyWtoqDlkwwTJ2+VJPPi4jlM9KTsC6kb1tX
BheUoAlrZeNe5Qg9GEz+epz3Fl4QspzXDWmIQHZq8ZNS886X+I7huTaejKrTYR+++DEBvOpJLo1c
EV0itdp6ydZCqfZDNIIoWQus9zfdVH1ihANeK7LM8dru7JJ2ks+cvD9jD1AEo2yQ2utA8X8stO1O
shyar0Y+prNXn2gR9NCUF7udxDoXoX7DUd+XIfMfYFweiALliRHtLnUER/ikpWitri+RycsThf5n
ucf8ay8NNcL18zPu4TSF8M7x+eQ4fJLtMDm5jcqvznm4kRcfUYzkYhQaKQtvo04ndD3rkn6Bwmyy
NDq6UPlPpfm3GtDc/6nNX1E+jnrXk+U/pk8iHd5hXWiwWSi930U/H5yfVq9yNQcKUMhDoKTFS/iU
cGf89m4y/RsOZ4+Z6EaNt8vmqCzaJ08JPMormUKjXR8WL/HRYhOct5whEsQEbG8z2r8hJObayTwv
LZgFA2AydC85Dg0wsTuZlJI4wgTkuos5lD1WoKZxqUGDkJEY5QGYZgPTBQ8MnDqcIoPf5dsEEBIa
PXg8XwUp3Ckw3qiUD0p2ExeFaTrQT7s3RpYbwWqb2XiqMd8tyPm+hpi0Z3HN2ZgSOauvTFjgWB5J
X+GFHrVQdd8qYgPOKeR3/dnDZqH1FsgtCdIXda7QOgSaQZKHyNJqJu6PzbA16yUMvMD046mk3bP8
2ASbEljNmipHr8zr7mbi5qqUr+rxDtoyxQuk4LbArwlEyr+uxBmRWMYYcClYKuA8SPv4YeCfvu8L
xR1CoTHTk67PWsVqB9Pb4CuQJManJUHOaAxy97XGhf5LlDQxWkt9uY+0wAxheW2yZOMrotd4oj4/
/SqE47tY+ETbo5/Tn5egkvxg2QvjoyWzig6sT9Ht3QGdW7zmm1/GzB23X0JW2UfHR8gA5JVvrdt6
7gzzNkMFe5VChFVOfu75Muxz/Bag6u+S1SYXCZayWZ4FgqJTjBiNkzGDNsQ9SjwdjZ4kAVsYlYKF
c0pPjRKaZYm3nC8BdovIeAbrZfZMn+9A2JSQor09fyjxpGXwf3xc7VX78+F2I5CxsxT86iwES1c3
6+cXtBxuYSidMzIy58TVXBGo1P3ANOWj4Me5mw5+WG5pnXwY3X5Wnb5MqlEzy1MfFfp2aV9tpukS
kCR+OOm8wLHCWJ/AaOxHyGV9/LkL1Wmp95kqSRu6k7TUgb+53EEVIkzsnhrcr5Z5wEl5/dq4VEGj
e3IrA0/flOpQgecsi19toO2Nhnd1t9MH0XA5cgMmSpbbGwb0seVOki1We4QhSvC5VW3q2FWnucBP
GMHVoDzwPLuWjDugMuXoZcGsxLF31N7boaqApe2lwDv++2gWlYPJSrz3Dy4sy8VmX5z50o6+jNGA
JAlDGAoXEoY0vevzrz4MlrlvqzdtOX0fGCVUMwPFcY3dAjPMbyzfGzO/hLve3pI3hGt3AzjRlu5x
+EEzXgrA06YYQgRAMgm0/ynY2ob4olX5bUVqADhVSxv68zYVFoiC13gwjUvUpbtUK5qxjT4L98lf
KDxaKw9fKFc5dUtxjJKx3BpfITYJfxLHb1DB5U0A6d7TfeF+oVbDL5+gBtnwiMSx8oOhkAXjI3pU
FJe9+p4qraiGvEH2xERnfUTxiFr9OrI+fQ7cgH7oXAWr0ciKgOQxEEQCvAy5iFCuNsn6Q50ApBgk
QUMR9qHzADxcoVRe36yFcZPR59bSY7dxUOD3od0EftxIKkJ58eulZTLelVvKz4uMY0ez5hwhWA5B
2Yc+zsY1osRBdIG5t59xWbiS6OzpJtqqIHrhMCPyX5ksbICAyN1UOn4sqjTx4hArb8Hp6jxEH7+F
BjdeR2y4/W1iYS1ql8YnDiI9jST/8a1Tr4aREmoVNAlsF99n1Naa9Qs3y7fubvW3YxjPtgdnhfwf
UXIXRFNNYWwkDo+3JKv9Qog9tDLOZnsNLR8VHPepG9IA6BhK73HwnUE8tiFeKVVMZ9UGc4DQ7LfF
3Cjjk2V1lJwhAddpc9izwFDEkd9wvYHUfCBQiNK5dh5syktgbM0uGRxbXBo8mUAqS6JtKMn4fltb
LznLji+15G5Ae+KFsrTf2lgbgedDZDNQ/ajluJEMDdPKGncDjgshlazYm4TdYF2aIs3Rmx2/VjUK
6j1GGK+9NksVuormfwuygbr2Qi7Wo1XBk85/h7rzX+i4i4Ulwr5nlsYZz4KmrnA40x0GCHIz+tqI
AKLQgZu+SRP9AsuD3p2uSpfBEo/TEiprzAaXUgj6UomHDFJyc+SVXoGWNIU3emrjqctB6pg3vbjD
oyBAXRZvzee4VpBmTCcmZVoox6nTsQQntp2TdKltJjnPIiskUt9gIwLa23lu1DTBSbxIQj5z2p7y
mxP369/rK2DexDziTDP+liPFPCG3TyPgyfKD6x1P0Zjuwm7p/POMiB6j1Oag5LOr3wcf6M8H2O5E
w9fu3qroalbePs6UhKDsiM58N2sefiNJrnLlHAnEZzOQg6vBZfewfIABUuEs4o8jDiuqXR28VR3o
jbMvJx3r99dIrZKi+bUrsyzMBXNxKyq3gRazNNlIMqD5GtqQCjrhUg19HIVQ5hV0mDfk7W/9B/H3
y1zfWDcxje6b/zkboqjcJ1QpkSWqGAwIIeukhlfHHyCQipRl6TBxqyOVkiiUktkYx8OEKO1kDDXG
Aqo9OUcH23rJnpDmHzlOF+Pa1iUO58ujY+nR+livBFV/Wx64Adf59nt5G1FhbYsIiRL4Mp2rTeNJ
qgzsc0lUGTlwMdbfTj7xEgXlvOCdPJPPuCoYDYdJ4ZJdA9uXs2HpwvqPHgc6JwR7W1KGonA2m0pi
28kwoiic+77I9xg62cpftEpvbaEYHCN5Ka5RI4yVrCUm0JlnpMUjLxKCMOfKtGIA81HBngH7Bd6J
8DVQL/FR3aH58/aVmhNvicOjbBFAFzSBn5D0pWAY/jI71NxSpjdBU2yeOknKXyWLcZ+aOa2sAw2/
RQdRO2TkErhejaXLgAPwpEMNv3QNxqI8GaBH4cvodGDtpC07ltJ+YvzzcWv5gU5FMWbDI2/aDBl+
xE2lATEw0EkDZuPQPQVUuv0enlG6CqQ0DaIEmtJ73O1Pk/BXHz9lOOtDb5Xw4CP8yrMCXkB5082R
bdMywKYfrfq0UZWu7/W4ReoeF4JE4lpiEEc58kxnBrMAM/kFQBuZJUcJiQQV9mzEQUbDXC5xKxsl
yb10CycNcTmvXU53AcUhrm5wdpODEcr4gTJZ1V5Q0C9E/io4AGKYw44cZuUfQL1VpHudrqqA70gY
z/R+RBK3PsKX6ceYqqqrwSumd0bQH3WKKFVFnMlm7CLcYjRUtjKNI3xEqwkBF8ehRhACrnePscAW
jobYL45IhO65NMi5sqWUgof707/IRDE3hSpzqKYNjLIpxMRkG578KXApOfp4CDCyhRNxw5So2FZO
kijd4N+rYHvRL16WRuCpj4xamwTBZIstQyBMPAWNSNo4gZ5Z8phsmNrXA77eJXJRSg8F+/RRJ8HY
SYvyAeV3MQNQKPsx7Ue7cp8HmeRitQrcmoL46zIbb/vVugvLdPukvZl0jJuZLjSjzD4kdqBBsXya
bQudgLQ+fPj28Rv17zipnMGyw1Jfu8m3AOmh1d1CS+S2VXNy62J5pp7t+6m66P2VPCLCYNMLr0xi
C+oBHGCrbBC/XSqXu8RFt1n/28M8VmcgYon3bjMwXfmvQkpngJ2foYIgFBr9g+9x6dG9eY/qPbW2
k7sWwg0dZGyJmO0ol1NO7VkNKF6VvjvG8VbVM/B4s9z0IaoStD4qCWliGVEevNNEwFosUgFQn6oT
aTDsAibEs5XDW6fcCqlcHm7HLzNytt2mMFWvrREfg+Kr/nhBv+euUDbp9sSumHcvHay6WmCIaada
4Shtkco7qRr6UugLx8/xPMULxPSRQmqjqLQN5cc2N3oXku88h4mtQ5J3dAbCUPbYVadnn5A/zEJJ
RMAXCIkzOI1maVmNcJATIL8J+baZDu07Z2kbDcXH5YaYkR1xTqFm67HnmLkahbv5VmYqheOcUL5y
2rejAMy3Q0DQUQBIGAyS0CG+u8wKLSRkHgidZYPcONnoRYpxlIcGQdDJ+1gPt6OVvZv3Mehpsypy
DxhqG7DxfxKeMWob1ULQj7eI8s7nR16HuYbwfloMsmY08ZibRs+thkQiMYy051XmN5i4dJKiSuv9
NUqgBGN00rFMuRL0VZFK9qXYoyuavlsiZxj/wpOJNyl4cg/HOL5bi00H0NogduTtSswHu9JUDhSM
7/+MgQqWv9LOO35eMHi4Id3yiSU92jwZOKlcLoJW+Q1CEPCaZ8RzhQapm85CvKtFWkiUpKq4UHTB
m8Q8tEgXU0uhkXgj8ajpgWGh8dCJYBmbYSytyvm5q7/YPksUIF9IzZOXm6J4JbLY2bP8aMnQk+6m
vbnwH1vgvy+F3gpeKnl577QBhvSUXoHY6t1uMkd1FZWv+ZovrirSw1Aj555XG585UMHMdBwpu7rA
XUii/xCEL5u0mmiR/5NcSsDxNKjSIsKbLp93/wt8rg1rO4hU4+qfXjKuDQ32Khw0vhcjn994+Byt
cdZtU6/paiE4yRPYv/r8L7otmwSdOTXjiQShb4aTNTFMoFTWhDNtWUy1el/5tekxtzFlIOg5sRqE
RGUS3kMWElx0OEvBLbYqzU41R49gTlrn/z+4C6tarMf7pEK3guylyLOf40+VmvCJzpn+bIE88diz
5DMY+yVGDFupmAKgSDIw5d6m9DY6FN4AbOXWNVsbx8k5SLJJi1UUMIUb2q7WdvLHo8QK62RdqnfD
XfdYynK761Vv23pEPt4+oyPT83mDVsx0IZGqPGW7UiWcL3G5fgMajXil5tPEInbiBSRWfnt48dSi
HbboDhNMw0iofFhxQmLkO+LowISE/XTraI7nn0cuHV7n5Mz6EI++6lEwZyOxyJ5ZjGIqEhuj4pvc
uMRf1SvUgIJxekVebUekPL22iZFtRxW4Z6fBUnEeNHryles4ClnZtP/R+KdZu5+DwBnUDWhSMlLs
vRHXQ4adqWH36B6/lykVt7H5DFjUDZpNld13QEWUam9i8dJzQLBPY72BimeM42zzmoubwOhU+t+E
MS0rwER40D5a9Ku/+IfFoXS8+VYhTxrBBePyKEyyNJVy/Tv5tsLDcK2WWvtbFb4r3LGZMCH6ZrNW
7voNlqxTfgHnHNGXSywDFp4F2Euzpe91LAYJiKt4MMQaKhqz5uuhTiwa4EvaczZYjjEkUoqed1iE
09a1kAu/4BhSAPYrMEMj9HRNpRfXpVOxxA/NXpmi/jF2P9lQG2YEkq0ERSbc5cNovnKF6813gezi
WUh1/3t5ZedP2ptMeuz6sE4LKQp/1k3Jqd3qGGLHSri3xvKOmSQLoI1tBom5QuJLSuHEXFLMaePm
XOb/xygRQ+b624+muTZcIuSfDwPkGTniqaCucj7YllpJuIOpjh4TWaUcHya/HY9kro3gXBSgr8La
F820s/u2T/rvtRIsgwVcwnWjdWc98WsX4uL6I+kPDTphn063q9PYAlStr4v98Ws0TgZOubd2zgJv
d0irLpcZ5mOiOjCQ0hfEzWM7Y7aL3iKsMNK2Xh7fsibhAxGWi51mkRGbkWtTCbfGquTHdoNFwdXw
09nXNKiAUMLQUQwX1O3SaCHlhoS2j2n3P8Vri00ptuY229fUd66t1D96GT1+uk4Q3RQ6Qgt+aWn+
YAYdcoSlcb0w1CbzwBr8fuG8ti+ty5CE6KL/DPoo42uWyEmBTGO2x83uK47qCfSByaCI3pq3LlXd
lUTbVCcf+4lKo5AlHtVKHmg0g62StY6USu/pvjCNIwWBVxt+nI8cT5qpEmZFscC7h4RTXGdiQiXE
2g3vYD5eaeSoIXDtAp49K0HyAMduPSU5kS6ghuSrhxWul8T/Ch+hTQaLzJieNyRW4XQuqhEDbMlG
U2IFmV1cWKmh6zWL43CJ4sURwo2PZJuXibsa3oE5yCg2RhaRzclwocZkQgOXNvJkLp7ihvvmC4uh
/Y1aMhfxLt4GTViGrltmT4dt1KWTt++LuZnQtq4ApWSW1ZRDU2LOn8An3u7FVHQO/BENVC46KfL9
uzxJqc9HiGbXxzg51rXYesozmDFCo4YDlrOf+ayPvSn82Z0UuUIQ6vskIHavcpcOYgKPhDRdK3Ap
gCYIcmAHporxK3T4RKxF0rX4/nHmQ1scJCdvre2QjioZEChy7YjR8bOd1qRR3mUNnc/Mb+dokxml
z7XX8Dj+Lswf3Pr2PYjAqAnyYzyL1z66Zcs9aym7I6xSajQ2g6QE2mcJmM+arckugMjqCDCnwZ/r
ZIXG5ilxYuBNgU13copPH4x90waB55tORc6X6xi3Sp8IAo86R9paZ6eowDslHQvB0YMRktYnr3Ng
iqoZNnqNfXO9b3hcOn8Xvtevsn7L7enk7eAWYmw2STRybsTSneo0VZfhIQ9vHz7nCWOZkXG74s0i
Zu0NODspt0PZ6rgQHLwvIR1rS4szJBd6H9LaE7vn0EwAaHAq6kFMpO8zdsn7EVR5msh7Iics2iLw
zkdPG0NQ5Mu7kei0vur7mFuW/kUDsJxmylbZERCWWBUssle0zCF2vQygo7UTYLcYPxWy7NxYQLn2
oKd6SfEC40kOmf2+zEvmMzNRDECYSwrvvg5C0f9VAuZpi76R5yZ6e3d5K6IXCU6F9tM49ygPvjzW
3BlwSoVG36ER+RX34BMWXrFNnVujPU6Ed90fh15xu/rtbUYm8pZQH15L1VcpYGKKJGm7HsfoJh62
nLLvTEHdCp00OjBz8b06Wa+mLHKM972x9POHoganGaH4V5bZSUllAsRiwqK+a2Z0PGcYbZl+n2DW
AhNhvJapex/yUY4qCwWssciwC5E7zALxDZ+pTlG1s4Bygg4g81nCNbyfmUY8jq5t76vTkn18QEJ5
36IUPPVA/SS+Z0eCROVhj7xkp3vVFOQvU8hoGUYiEPBqaMYQAcmfKCZvlP1zXLSGkRY+SBp+j0IT
KDxP6iTgwXooZrR+FUOQR613iFqL1iKklIy4Jms+SqN4d4SUmfJRaSXxBMy7a5cjDAxBhPIFIVma
NS5tNuDACXVUcCd2LY9yRPcLJW+s2wvizEVDznSFf90BaDbuWxJT6egc9e7xgJV7iHCsm2BsQdFv
SeOC/UAhpQRf2gstF9phbXI912SmKubDzK5AMi5Mgsn4VUVWZiCY6OlRD4Hlg0IleGpqasRDEIbk
lA8qzvLdCBcSedqiv+5vzVsSD9cNq6avkPPpF2+qUmPPIjUQ9ufkam6kYgoo3Lu46b9CMQY/kVxt
tVDhylT3bO9/tA8ySOyn6TYCtoZSVFnMdShvzmUAhkg6Fi7xH5W/QDqVUI2ZZb0jb99AA9dGir24
DqbovrKx+0w7pU2RL+mDcHqB1J1f28DGhjLi8jqsUit/N+85xj49VmBGg+kACoDQxy2dxNM/CnJ3
zk4JvcaDpvNe9F+F6zXnSiOcnJgFgaJ/hLbOpkqQVGBirDwU/N54DXgwU2ZMehzi+baQLmlbhIba
0RtpVwE/RKkEq/XTy2niWXtUEXoJZdxnr7rTur+HQXFJkRYrYL9x/iDQgPEone1YKGbPr+JJv32Y
2hTOcwN2r6hYvI5Vyc9DzwTrO5JkPjJLFD4nrb1PJiAZWXN0l2JogkvyRDyfbEtcjf46zqeR6i4K
bAtcyyHOXIDCjznRfS5gXtREiegrN5IvptfZYT70OWBgxzFSeAJRViBX5/gcjBjNFxXG4i0A9UOS
RtpjZ4vwD/VFYTXnT210/hNEr6gCxaN6YWgWHc5xNhTUM6HAjKXK+DDsG3eJ5eVXnKaN+CtOBQJx
GRlBVR71OMNybIOu858Llb+P0zgc72/LLYDAYdfjqcSPSq4OvYmKlE93PGm5aiAdjtzsdya7pF2e
kTv5Mf8fSyS3C1Pnxd4QTRhtqTdywbiG0WIg+gOjr9oY32KDYMbhKlgjhnjplQGWxSjHhfimTvny
A2M1OIwHhEH0AuzgE+U0LWKi2ktJ/Cdt+MOgmHX+Ur50WC/xZWjUbPSjQwGBuBMYRKSOXYCa/mG1
0OdJGTWNBpnA/CL8jLrSL9Yi480pkYMa0Nr+O5BCneTM/pk6X+InZSnR8Gr5JFyc8WHiuNmqvx7M
jDjTxv+pjpZbtkRroqREsBX8ahqzLX52klpDMoXfCIZaQK886oXEfFJYYJBx5T2nlXuKtfyuezIZ
pEQcvLkfLIVYWysgDVWml0LuTqU8kg2EQ2lK+kybvkyi4xU3ZZCVCxBWZwM2dY/zM6vEBSZR97b5
9qYqChkKutOP5IL22sY/w+b+vfJI/yLRlJEv9R8nxSpIg8oI5nXZiBKWJnLo1X7bMvg2Rq487IwK
Nw6Ecf+GE5PxlsuL7BkQsXcNoMwX9+2q4so/By82SbhLgrv7EQJyAqfrYnbIO4Cs4dWqjl+sg7Is
TSbaEpheQrEFRj7Z9ol2k2TXIPMQplMR1IQ62HCHDG5vo41iV7nwEFx11kNwTR3qbS3XfJYrZOEF
7Ela/5ieeRNs7SuGfMafTdiYXBqwYOuFBlU5R2OSkJbN9u0KHy/eDnFUcRLGv0yuMyjTfmnQPAVq
eZq5K+fyaaECzwiYXFlDm3MnPqE2FKQjros989/wzi9TX5SlMfO6bX5GVUDvkGcNVYlJnaCzc6QI
J+DV9Mo20yA6A9ZCjUsuoV6s8ypMYjhJ+6Jo5rt0K2hV01YOAr/ZuuRujggTVlk56B2graVl+4yp
Atr5jeUEvrKMPQpUQpeT0kNosOJMdM0jXhjScH5lRAbe4R7yJB4/rM2jYSmMWBxtYzYB6PdKBC+E
yloFQMeXB+UNy59qciNVVnWkpkwV1gIBdOtvF16bt/ISte3bj6LOl0Yq6yojOBTTzHjaZfSMXZvo
pNM7oEB0L4wZAwyeko1C+ejwB4thKe1ITII+t9UxKGOXBekNPSXUurU2LvIcDsSZ7f463hSrPysN
iCb7CjVnQFnwBL3oaENUbsLTQ6o/ByheOu/WpTxa1nKUsYECuXvOZCfLIqGayJFhHgKb8DRBRhHu
f6mLBTBCBAhvRcZ8eQ1WDn+XYSge42jQqtIJkEHji2nyHsVKwF4ExupuzUMRx3CnIziG94/o579E
FoEMVT3QJjSwiAzQsvBZ2fDPwbtEjAg11yVbQ8K1xJKucJ7vInqsyLk4K3p+NAxOYVppTDdR5DwD
4wFnnRUNN242gGwEqO9EotilCIATw8k1Iqs6L9N6hWUCVBhhDQFRJ5B7Jfl6nCIO5E9OIe4bT2o4
wE/31aUl70oTD0BqwPEvJcEXNYMYQN0/2IqUrzGekulSeYSFVlMMlXHQ5iK4LJHH90bkm2Pom97x
eODMYpB198YgtgFkOBy8lGu7/UjhZwAfF7UHCKZpig3hTw+/rJ09nzIx2VjGmjb7POGagg6EtnTL
ploolLLFnSnQ6CF2erCbe+Dh1Z98xBOjhFYDr7zIGEGq//rQBSif97klSVRYIlI5n9Veq0yjM69K
dTZVLFEJqGnW4o8GmRPmqPj2pz5/ttL07zfjypoRk0e/N7+oWA4CRp+gZzjJ7+xs7Hx3N3VsAKhW
/BC4Nglp8o8Ns75UGn1PGIE5GPvVnMm7N0oCN8pwbofp7wUYovAlVXjM8iKtjXbB0OYb7l72GAZw
1DbmfNCJANRP9oUj6PCAvFEB3WRAqh58+FRTwByWBz3Gidia8Z24KZbaFSW7n3hlwuZZiYh2L0xH
mEnLPG7jEazFsSjpANrDYYDgJPEj1yRaxu1d5Mmq+DmtcxHQnv99qTdA4HorVjFHpXrCVhGvYszU
Zw+8qN4+VsI9mLvipryXHM6wuVcCwgouKE50rDCMhtgFJciu6Iz+LI5xZlSHZcwUXKSbx+sPPdCU
84mL1Mw45IWoM/VAqeZb4JXFBaZ1ZywNUtwf3NeGb64N8JCvJZKjxG1cTmYQMI3p0YpZEJfKKHnc
3kuLk6ylJKqm0DDVveCwMJ9DH8ZJwPhkFKqBD5TMKIyXuAgDL02Gce3qq/AGbN1lcn6QDMSgOOjB
CHy8l/H4av4+QyALzRNEd74q4DtTRlIJFnrNLMezpDpqGCWTB2HIyMHEGhP/bYd2fP6R/VTq00LE
SVoN1BQZXFTB4APVpkFu2iSWXE/3qrCP/ZxIodk9t7x+FKikwx5YTGj8gl9wYFgSt6hUuCj87PKb
/tXWZAFGb8aYwhkkzioYjidDAwrdWNAK9ddRrJ8i/1LnloVR78rCYlzTQdd/sPfxjo0FCySgWLM+
zIaqFnnZboPsvBbocuWi1Vu/9iFlZJ72yQXn4iOEIrDKJ+O44DKe9hyC3nnOOlHjuLIv/ccjGJ9g
HEm8UVPUxMbZXeLoPoKT7WPyrvx1rKThKf5y90HkwFVl6mG/XvpdjgX9OtBWnsx/acsSWXGmx5yE
xIDtOx6eqWUh79/kqvgicsCBaUzFm2jdO3KIsTYQo+dTBH6B/ai/ez2rCBSDQWN33hVTb118o+TA
cJyKh3mIZj+IuS359Ix94UnBVb3GQh3zDYdV2gqVEvzl+dKVbOZsCCBh3MDW443X3c1G0hHFKjiY
OE2FEFFezVlRaC7/m5k7qjyWjo39B3keZies+TYFAlRPwFgeDBILqurqSFlKbIebC84qoRD5rGp3
hnDr0ss0vhQVshK9I/xNvRFkwBsJdTUUG9OJq7j9IZ3GlbhwIM6LulXrf5E1Oc/0+zZtOKbTK4lw
fEJBSjxAcg8cQefj92SDw0kP1lzNKnQmb7xuEy7TwcOGLG7A2x768sZV14c1kAg8L9DosscbfYq1
DyvfkRSqbTY7y4WbHKFy6Tlzz6mA5mNTxzdqGrybibV1oXa/dOwPQJQHo0YY4Qk8bvYNZh07Uq9v
YMp6ahnfzmsg/zg6L//RKsq4rv2JnSdHJPi5j+YgdNkvVCCUpn58oa0PJQPmbNQLJDtDcWf8QVfc
iva4p5KS+KtkLE724+vcr9a0J7D+kh3OxIGGsdLa5ha1cSlZ8HO5zX4fBtgF0P4+tKjKR9qswsZA
deO+IzZP6xYLdrzonyuo3YKlwx4XDNJ33Z0WcKKqb22mnsFRd7FvOC144TiBATqE9enfTuCzNhZp
WZwMXyZShU/EtNoGTdLEsZOcF77FK44HqCWFgeQTcSRzeIMrxde6WxQYwqH65yNixMK6BYgLlXKe
XycKVsc7lT3M2ZkT6gc2EaqeZFTS/K6RG0CmHuKDIb7/WXMXYu1iU759I6cSBoJXnBJc9DkLEGdR
YED4qCq8Gbbej+L4V7JXrBUzLGjvT1KoizFEIfNC/o/wqBMXwkmWqST6OcV6uLW79C/hiidlkuek
wND7onTt/+/unrXDj7+nfR3kwvlo49mM2CQ4xMiQUpx4siZ0gYrqb3tir5/UZ1SjvNS3Ev1hgr2j
O5gq+9KdHY/IXxAL8x+VdBd98DyJx1MaqUeQ8Rnwk6ejiQoHqOL/oG1oQTEyxQwRgTf4jRTBUpRz
v5HZSm2vPoAhHSGx6UFisUSyMEltZusfeLfGUqHXtaOyaeANeCbP3JsufMWY0iJGSLS3Lan2SxVT
4AUYlkYQ9se6YImrbw9yiMpHlEm4WTICQgOHawcORA7C5LAgmp66Od/xLbgUk3mkoVbyLo0DhwJB
tZIcU6eDDyntVF26ekSlDDqPtwWlWck0ZMoeuSVZJgHB+bfTZrzduP12S5gjcm/1Bo8v/9+iBPLg
8MHU1uWasTlpFFOXpLsRkbRS9Kim0h6E6ebDWyfL6kVOy9tan0MrchlfkK4jk2izqnSitPGrMQbs
hRRq0k/XICM01sfoC7FjXvIV2dQyj2AXlCQnac6pHqR6BEke9tEYnpKBJvbyfqoYUGET3CkmB4NU
VjdmWIinpyhIMsEFxGkI/4Tpj6z+TxrSuvvokBKAq6M4LkDKG3LBxOez63G1Bs4Jgqd6qW0R0zZP
L0BcJfSkZXWFUj9CzUm6W228l2iPGBi5HVgk6pu/+iOJ9bJ2l4Rt++ZGzMtIYtHiRo43VEwSp8iI
VM2bbMbFl/KrxPZPlxem22e8Bc560ZTbqMNT2NDcT84rrXhBdcf8SAjvm0/8mtvLzLOFSeLkvm77
qBIVxpAHPO7D+5rno/cebjdp5A597Speu1gWUP/BQpljSwPFgkEpjSclgdnY459DvofkvnaGq52g
SOP16ljIO3KrwuBaV/MfQk4bzAj7ag9YqrGMPVTBTF1JjuDGvz+9dv/6zzUOVmwOluexC21X/d0V
8WJlsdEf/zqDCo+ggy9akxJcmowIVD60TgVvgcWtoW1mWpezpofRWzOtbxMHFBaUcvShO+fEsGDO
naVMXe7psf3CiDDKvQs44xbYE2BcdQ2EkuBlxyWQKfVcIQ4TySCrS7C2oh8FkCwDX7NajQd8YTJK
CzUJUsHgGRF7OOusewFyhGWYy5LM4vbcTWw6ArwxHYO5tGPkOKRy5W5lDvw6Me55XHB0uc7aGNjP
UGuSWJes5+4FIa7Gmo/IuDbTk+oH36CyJ9PMf+Zpc25RJ2tIGiB5876PiVCU4HtYUYOjtHh5/VpV
NPJOfPCO3bUMXV0W9Drxmrv9PMf0PkVUghyihpRTuthrCTByWMAfAmjN5+2V9j0trc5ETRyxDAzP
IWg7AqfBPdSCbzRsU8YxfsN7XFvGrj/2QbKRQiNe7XC5SWaSBunAh2+ZTohcVCw4DJ8nrZYXgVeR
K/R5x2amZbFv3rUO0cK2x33KyoponvpywXkxG0vu9VS8Vy6GnkueoPs50ZdF0FaWNsTy/F6RU7kL
FNxKjFrfobC3zVqKxrDSg1xuoLQcXnRSbIYA0Kor97v0Nw+DOC9Z0nt9ZF+sb5G3vLzVrFQ8rZmh
zUujSXgEjeRMheAkHMY9fEOgAk0tT3Alp0nCdTz9hPTvcKpEmQfMPGExi2qc9FKxvRGn4Wel92w9
q69uCKwKayj5KNHuMJtOTyZ/9Vjkm5ehkQ1eHl3JMpfCZsvv2CQdtplBunoAPiFFBrr8GlfnbgLg
UcAOS2Bbx3yKqrDIWADgAC/6AspAFqz6t2naZDLvgbH3JhW88zNvEftGbZkEtuMS3ndOSgiXc627
rlWs0fFx68AkB6fNYIHsRVMojo1Wp3os7hIm60BTjkdOfSAJnnunkzLWT6+4rWMidjiKOeStQ16Q
P7at/Qvx5493afRGFDqsI88ueoeZ3S++KNEVOSOasQbs4v6lld9LneY9sNVpxfIrjsmguhqSWN7I
Q2R3d7j3NGki8gwF2TinLNVnsJ9ibfNgUQeotbelJZ0Z0WajsXJUsjpThcR2TsFr+WFdRE6gJ6hD
mMC9fGAtYiwe+H360qXYc6ERXw4rl5hNueS+sqm90Zj07UjJxBwqrhzhnLgjzKyHlRLNziWUeQ3K
tqwq3mnksTIOUVIbKYxf+Okdgthc2TSoSnFSN59x6As09/NxvleNNxn5lyKTxeLrD6KNfZKPtvE5
d7POZ7QwAkrD+xpV+CaRMIPkL+cwgH3XjqdSqyJrw1A39YDvo2Tc59ztnNV9AFB7fuZWc6Ia/jqB
Y1B8mzwrOhReJc46oTPZPYmszzSTMLUkVTtDmAYLJrNGbknN5n68VAsqEyCs89C1StuXhawHqzZ8
qKfxSNnVC5EIQIMLVJiRE6B31oSpPUzaATiaMcywQTXtuHonWIq+HtOP7Cw9zPAHmI31AI99tCy5
QwFb0P+X8HLlMjZw9QVsswltGugh6Fciynxsan8kLqPJPqxjr7t00wBWDzxLXCzTEvFf8DOLTsNy
sx2gmUjT/dUCAqy0YMKb0FR160ikwYArPxxI/LxM8BKjywr32MeSOGzttOtyJKdEuIJmh4RBatxo
cBEQArJSiZifP1x9M8DZ22PXKr1/+Tb6+hMPopDrcgDjUXcm5dxSdQJxMzQ5b35KXRWee6cQ93o/
bzSsU8ttL3UndgxCx0UFRjr2KUr5DFDkzlW8b81lrcr9uhXgLTSumw6ST1KsynKJhH48VrIEH8r8
eiiwg2HILWCeqIs6QSBrHsmeyKmcaz9nl0HKesm31ZJti/nLC+hVTBx7eySAovMdI3iJSm5Uucq5
cZmkonY/VL3f8Tky2DSKlNqSp9YfZ7XxaVr7otM+cXCAgp1eqRAl0zFU6Ka9S1DMeyqUm8uVBODL
3cqW6tnM4ct8BNrm0U4dqMhmF3+5QMhQ1BfbV97T7j5AoNzOHydwJK1c4JotVr3E8u5RbguniDnK
5TJt1Rp9L4QE5CAkKVs+T3ewZVgfNuLubvKWBU1/b41uQaxala2svGsvB6L10xo3sVPnIhjWOH5q
9j8drEmZU0oVn8kZPYoBw4tWy56OTp1aPEOmvJBrRRKbU479zJA4wlaB32jh+jw4oeR5Smg+BMPY
wQXd2gaKXkAFnLIiD6PnhsvasQvj3l5+OwS+4oCuFga83er/NYynLYjvRhddMf1MFdpKo5H/sajE
oQBMaH1uB1f94J9i3p+6XdDFqpT1tYCPNvpmuTrdfFuwvs7mkaJKPkJm9zIIhR0KZoCrSGij+Qj0
MnsEwC5KKgmnnRzm0+S5mrr4ld7IjcFLGCTyxPtAcIfFsqRac4kXCt9B7aL95FLm7eYKli6HvYXT
H8kFVqqZ8bylOz3DhHxiLpPVNSCS16qG8D5/W5csQDvkyauacQhVFK2t8JzHHQFaQ8Opwo/TAEvC
IGctiKAna6Z2k2H8LlRM+T/4R9mhrpcYRdLtksbMBUE5LFaPVdk7TeQItXtRDyKLnGRet1net9Zz
4KvBWHEntclsse3kQAfpywB5spI39yWESD3He6rFh4uTnbqKew36qAse84xvA84DYFWA+t7rz69Y
3vRGfTQpd7zctbXaQMEfFGPkA4q50BzE5nlUOTvTHAksenekpXHZle8U75ZIpNNOlPb5GEZfRREg
TuZbZJCOE8xBuRlrqMRhbnh/kJSXJ//LWgIP+PR0jcMNHnU5h9itKD/wB2eUQtjnNi9mKBiUCnyO
ux5Zsc8rS3zoMXoc6xKytADvVMc5J/wqS4dG6q5Z9wdPXe9bdeZO5TGIGxfmTz3moVtI9g/GqeKt
1rijFL7UAHcV1JXq3VNypcBW6s3c93NMPRbnfI7BnBIY8PbJ+S08l04CBZKO4utMSM0V2F0hM0j9
/k4xDtyNSFqmJXyiUgD1Bb9CMTgRScbWYnxrO6Xl8Us1fx1UR7+EDWjIXQ2Y2tMXYRfp+Isxof6A
FF9Zu/a90a4YOQ3WcJXG+4Igk3/l7zYKWIdYke3Ey8dJ9zagUmlnv0qv+hqY9+zeW0Tq+WkieRmc
Uy7YrZUiCIvqSWwP9naVJVeDXtiBEcwoXPRW4yVAdADYvIvGDY+qhERpQKkbXla8I0nyUJwbMvVw
IfrMw/wH/neKQwsRq2G3jqyWfy89+ABMHA1mWO2wuS8+TgmAZR81bESXJzV4yhcHYEuHTmmy5v78
ny8iek6GaOX6bOCcenm0L+BYPVBdUuiFsd9HmZWAsEba7892s3tWwccqWTGNhldIF9ITU0GgkpFL
3WjeuglCU6wJ98VlhMHqIcAnpZz4Tzp37keBXUZUww0CwRVTEIPgEPV14+M7175aiRuGH6cY59Cc
8tYb3bRl+gQaFEC5tJCydwVk/+nLYeA6Z8eKEyQdCegg/N52Urqb0xo7ViTQXs2gu8GZp6BwMa+t
z+VSIZHEWtpLJafPFMw8ip7b6l/vMEcLnvl4C6CNKYKY2z6NMJz3zHuVWFYOtdWNfB9J/MKa0DzB
7lxq8liERS+ZPKs8n1RotFFvqy5MVegLXjGtRlHTMBl6HEnWCFxzlAYAPa7N3eQGmOontDzO8MGF
0SaAAP+FGsPnIZA5QwsgakkOpb86INdIiLpWPrpZ/pRzfKZYY5lP/TncyR8dhTV0R/SPF85htfk3
8QJVYF5nWo8JCslD+Uw6yoMDovaNGCLRn6crrGIKyfUAHdAgNBEnM5WuVIpmkk25j9eR0ABpH+0B
GMdMFPaEg8vE2ghQwUX8Uc5pAMFmpkzuhbtGFYUG3S5OYWKpUHh5lf5Tf/VHb57zlNZCvbWKYyPT
iIhBaqX4sfbnZGGLTxVEAMeZjXVdOlZawS/Q2vVtSjPvp4IBfPtR/kOo9zouanUyukD44aSepVeM
SqVDuBDNbSliqjqQz7cWWlpurZ1GmMwKS2HLyK8P3gGS8rPjvdung4eB1P89l3eROhlHOOMTt8BL
1uJxAESoKWoNYrKPUEC+T4akGE6tmraZFT1BsWA5VVqU2BIaznj9k6QM5w+Lg+101vr4egsDWkDe
S30nncjbme09iJhH/YOaDmlmdlvRMRjMnlKk4Pl3ob8dkdf64KZDqDIVChaVCQiyQLl4qT856Px+
M5GOYkDDPFOnDvlDiaj5vww6oujfEaxGLNuN02RP7G9NHXItPqwMq/NkZcxkuo16IDtHws+AP5cX
2+tCJKnkCkdlJxwRs52HAIhPYzxbQrdTx/fjQ/U8U3gkAxKXmc93aTLAdT3gl5IAVAgRqMKtHuvs
LftzjX9fNAFWIhTdeD0QNCz7uszoZCTlb3oQVl82/lTNAZ2ZZPD3qtpFZWeZuJz7E3Btfpav3jNI
EKdBRMVPiwDaVEjFQW8cMeipeFv6lVMg/aNOzzmpKQgDTMdPcbUC6sgj5u7ub049Y2uqBwFvrpDq
ScrkMvzSHXTD9N6FghrTwHN3YNqvkEOu0GXPCLnDwMVsI9RCCMXE4YZQ6V78qz7kc+l7TQQwG7Le
H24XRhmdAFID6i7BjPPFfe6XgbKYnwsD+SKSqS/krqA7pqzIDuyhLrPJMwZMT2+yM3FQ2qAI3gZy
vsxCekC6uG/JKn/84GMNlsz9FE9xJA/i3NjBzoMu/NnSmNI3wi7n2nu/dYJzlWliUW/NmIw0Vkg6
upudEdb216hE6qhmYjJKvMDcI/t+7cjJXs5GmODXV8sS/Q78pgMv8Yih3enKTQxkivVCq3aSkOR8
2ViGIBY9YwDm68W56CqWuV6+96dn6DoE4PWsDAWv17n2kkzz8LojzwujK0ca+4fyesRmbu8lzjIc
YWtTZX1pML9nqFapAlW0NoaqCnPfu8aJ8paCwEdwUcK22lrXLmwkgcOXsQT3Zgxyz9delVHE5iZo
QrQpgTfOkzSwqKwZKyOcdQMm8ONpun9Fcx0vyxRPqdGAQ+43zzwB1bgzUXguOBc0itYiTQly0ok2
6/ZuqVXABmW8gWMqQ1DFejIt27gQ4N6yMfWHuXV4G7AVKFHkFTi0VsvztFqVrqQw7ZAFiWXfqdQb
DnQsrLa6nBsmcV8uaxWIEQshdvmww0ufohDfnUaO2ebroByEVdBp5EQRjEUc27kgM5ZXRw/q/SnK
NRCZdkW9e+zaPAQr/5b8fSIo5R3Zg0kdy7LUgk3hyFUF0P1VzqBKRPmODaS4WO3rsNIdcaTtTn/a
gzdwsviW0SYaCWTVfTzNabnE+GI8YiVmPdWz/lV8GYAFQMAycS7jgVNObHU8qPMRaSZIlRgBvPCx
hvkKIpl+biYPaha9MDpQcE9cLWrK0drrecnw8WUbZLLq9V9PI+JuM/+OL7YtLaQG79GWnSpNjgrL
uI28tEcQqdQ7ahx6gaYIz461acB3XZORKZaWfbOkstbhtwxro6uOkMrzcJt7na6cxa8h8FzPONes
CWwrH0Sz12+eFQYji6BOWcoxGuKa/vGPMlkKLxGMD7MT4IvDCeKbWhN6UN88+G+sMTPVYeXFtQ+U
5e7sX4wXzNF1SbcxX1KUYJY1c+jtMzOIplQE9XQ+XvJwZHd879VaVWdWb+VCzCxpkhqGbRdE8NH/
bZtslBAZZ3nFX6tRlXgBSbykMLdODjN3360BZ7Gs5CH27kMyV9KDIqXFFgDLCrSHfwcJu4xAekIK
5QOzkfe4T6iX8DdG32D0NepyPxzxl+8thzawFomMUwY9Kf2cFxUAvd+SOiZYTI8WYTEIQaF+k60X
KofUQorF8W4IswiIk8yG1D9YaMr0Fdp2YrZpKgt8A+ebWWCKxcmLWVtoRyFj04+6oQxfEs27lEKJ
FC05xQd8PkW8S/IzSf/cS9zMvTuL0voNy78nzl00KUUZZ9StzAlA/7TiCNQObf1P6S4SuIaVpayo
HFMkeFu+0z5k3JjznJMTbEqXV0zV967r+slyQZFMeZwZdU3UrGXEA15ykGBGq6ioCa5IsehK+hCn
O/3wGm+b5gbrESmJ3nd1AOKawdCJV/enhb0NhmvAY207ztpJHm2K82SxfM/McuCiR73qippgvNH/
Z9y+AYI3B+X+ysMZmFrbjt2xntk/itoPskpBxECyYq3nDsVGj4mLmUHmKPMP/qEPt0/68EOCLlnk
p2LRLLfBiwrs6pvqgkgijimhcJAKYU88ASs1ojvMbSS8XllDcQEo7m0v11+cZfIDTZmuBIvtVNtH
z7rB7JHZeSt1pF/jO4F2evh9KVLv5P69YPDa05R++1vVfITz0mqOi+WAlvKyGRHHGA2XwHtPhhvU
O1OMILVI/xWYLAewx2GBJQ2zTnGr/tXkk6NBNAh6a1+kn+rf/MkHM2vGWpoWkb4HzscIX/9EmRk+
Z7yWRNI3+PPh+Zl3FNHlAdSW8xwB5f7Lsa/YdDcFKox7QvT1TBDzmLAi87YRqk5vIpIcS6FmdoZ5
i72MWTpkV2QrkWCJMRc4kXUyqdeN9u4V97H+HDxthZkHsqLE5QhOyvdrNglVuNFBPwSjaNdCis6d
CuvZREOzTKqwfET49CFUx2aiNocZX9b6F2No43pkR20U9YO88VtT8dtlyUtCsAsugTz84d/C3hPY
yG/BHhpnMM8eNBMgAZlfbSDIBPfxb0fxVBAg7bPMh/Iwcf57e8e6E14ImOvXq2fCDfZ6dueaJF9c
sxLB3UZo5+wv4U2K8PYajagvcOIEZfodpAzpUwaR0MqkSkiVYZsbYZ5paxft/CjnxMCCCXhcM4Ki
EafRBn6XOHNrQzq6hIU+mpn9JT7FsFn8NM3H8d+x/DTGZPb35xlxByWfE5DejwqDdfbE2DBcgeqx
97ctmCGbzybX8k3VRbx3HzHmZpuse6Pmx9fiGyzmOZ27isEzznvuPx5TSKYohRGBii/BpFbQ1cCH
Vjme9wLOaZfPwhUdX82srpDGdy0OedMg4go1lyXEHKonLc2w8atD+dsEULsvF0nF4ZOU1kU5Q+st
nSl8aBogj8Ywok0z1//m7NZ27yBXNfDApSuhai+/sEwHfWYbzTUrbjBKR0K+S/DaTax8BpnTbMox
+OYtDNqnfYA8wFS3PcJBqeRmMtgQWmcqBY8EA2s5djqjjPaNHMf8vETfJxALO1qh0yT2T6Bqflpy
k7JZUfwe35abA4JacRpQXiLHBbyP66jWg6AR/IwcNUIGYeN4kAP2+Idrvd3OCv4aX7adhJaEQfCZ
lvQHzlL0TiRF0gml/sQUSoqFVo7pKzHtc2X0TaFR0mejLRK265lhTp7n+62djDtdXiCoilWWkOpm
5NdlgCQ7EfSdMlXe6k2lCjAYmprAuDW5KL4a8AjonFL7zty4Xf72nxAyEloeXXWA/AKImHcbwunh
vNftKc1+s6eHvfiwlcIGTyMvtwVLWvyTLvaAEXUhbyny5p2YN737lP20NCmxxzOeZHJCvH8NTVJU
dcSz+UaabsitxS490uS6MTu9YPQYIsFRryH9DIi+kToqCVhTgzMpdJ7Lmopm0tCrCY/g0cQFdI3I
N+/ulEs1GeT9d7x+g0/0pgOobPTie9ZJMpYmJu5DYTYY3j9v4Ba2m+GxmhGpBE1hP/dTtdtrHOAP
orR620gIN2nuklGgPLqpx3kWKRCnAOFjzGY8sRdqFxdLo7/Yssrr/GMjSYiuqBR3UBNdIJ+uZyaV
0r86y7nqcB561HAv+r9auriiMt1TsmlbyhIIsttBIKfuxnDCJE/2NfTjUBwJto8RHpqo04tJ1+2J
/ygZ+sdDvBAtiAK79Xc16n0SHOw3evHcB5t2e3nu/p/jv9I72ea2lFcl4mSs9C1hPil+RgD3M26y
654pfiNx4jc1YjPRtBFDYCuy6ucVy+pcH81hU8BQhPD7rSP7F+3ehZoAVzPdMNj2oS+4huReVy3p
jImuMwfOWM2GhLBT1gZnz8HnrQLO9/7/i8qjdOIiu3D0vyhtnF0s12hdx9BKTB02iRoZwmA1ajPf
PIJYBPWm8S1Zp/hgylPj46gX5kh7l9tyrkKq8qjZwbF/5L/zdfta19OTaiHgbpLm+p+wOlY9eLTT
EvUx4cA6BFaa+06Zsjr5/66LtkCcW8GGbAxqnEc26kKXveKQTz11iJpMA0AB1k10OeTOHni8jvH+
r2g6aAaCKFTYEJRXXCya3PQJoROXzghSaqy4eHXH+6ygvCoSlmgrRzuuByR7dX49gE6Th5h2s8+t
9YQ+wWiASEjeEQpZZUUECJPOSBeUWn1Lm02nKyegUK+H0UpiEJnT/rQKY1HfnWFVFTqPdLmDYZ/B
RnyXCGMvJCU7pzPP9dGcv35HGFbDbdrk29DWJAQ4GCUd9L8UGV729qFtXPqTte+Co+0OZc44Bg9k
IeoXotgGA71Q+pr9li6I/HSvrWe/BIqqSoZdxJbjTX+TR9gzTRT6FpgmYznWJ8Wab5EoKZPDCFnS
UWhT5FrlmAS5wTor/tj7bid1L8ifd9YM0UuS57GvXEn+KDN+RovkP94iQNwJUYDlQ94m8OwPY0G1
z1cERgcwGmorgOYqxCebniPvSlc8uaey1AcJmFjl5bO+RloIyW4o8ZYt57wM6cZ9kZLQzHtDi8to
wkF+AsLU1LqU3J0ur7fo9YsLgqVvW/eEqagY7hegaJALnDoC2Bsytk4D+QT+NFJJxOK2KSMPoMzY
+VANGM50EoiXslJiFOsp00bCp3X+nPARtOCzef3y5/QBwAyuYqKaHs4p2O+EK9uRxfbwZzvcG2dS
GUqjTYhbYLMjmd3mOUrBjh8yhtsTkP+j7vE9m4L2TMZF7hI3heDPv1/dot6JzcBTtrYectxsC/f/
qxea26a+w9H4niygMRnVstxh30SvujHEW9jDyjkqVucWrrXwIbFCG3dT/7e6Bvcl/EVlox6I+LKB
jtaOJM7cJoXWk4xZSuze0tSIbj42jsGyRio93mIJeY85r80nuBhUP7Nbxp2XOmSJPTuRk2ZZ8ALb
/e+f3jehBwSkvvL/KoFsOha8E0q7aW3xT5lzM/YbQu+izdIpXjmRrOf1JWhre6oaHBXR2ez6wguV
T46jSj7p2EP5zoQ3bcDzhhlgS9CJIGgSeHH2NBBNNuAAJbW9Jy4Yp0soMJJlfV4DYMGSi+Z30zys
ouEXMSWOuJJya723FPaNuEuZtMHY8zMuJnKpYUCPAOSZy1VUFgEMicqycrw9a6ns6cYAHqA0s4Hn
1QYf91i8HJ3nucCc1MN3luuB2gaAUU1kEC1EPrTLIv2Rb/FeMZRmAXO7WrQdUTLNubzbx1uEtV0n
/w+aTRZZOxVaAg4U7oNUKdGmcdLK/5PE6wsGUXoLsg3VqRf420y81+8S/S5jj1tiSjwdks5ozNXQ
GCSFH5wN0oo6erhisJ3cgQowDuSD6Oe9jS8fBpswAwUyFCSyMKvrJpwhDER8rbUa/vbNqA6QuvaE
g1LVTzgtpg3zZt4M9FiWHFbod8zOEgU5ykcsn8Z4WWyCJ9XBMXps7+PwddUhfoAR/LPg4okOomAx
+HZigxAbgQUts6xz1Za85+Xxd8DnfrbWy6abBvqVsebMo5z5XGZ9kY36xB86QExNykYtnDEC3l5W
fEumA0FNrx9A36g+jDd4TDenzu2yvg40fwOS+na0NmpZJgHXG7OwrbVZEbRAWJwD2lJZcncmBfEN
VhqGyMvJqh9rU2z16QNEf7Hpjq5VS/M1V/gdynyaDkCD9nPt67vdBvYJLA4ACcYH/Gab3Baqn6I8
Ees+MoWFu/EHRkqMbXPLiko/x9ko1YkUjsJwO3SvdH4Tn6HdPkl6/ENequq8h2IwjvIvNPFA6fpx
80sDUXbDjRyoUT29nAkM1Ik3uH9bZNAB9oFvy4l64aajnuVvCnb7ah+5zRr2t1CsaGop7f1MK6Zw
MoI350316X5r+jp4/C2z7Zq19TcMwH4GgTed9cjMUpOHzfbLncjHs18e9xt7n9GZS1lcxbP7Ynfy
GnJC5aTXtcE/9JdiK7Lh6Yw9vwEF1FfEqhw2O5dCeEVgiUb6HiBYS36AdQkVYcJr5O0aiWcI/wuo
52H1784inDjk8vpgqOC7PnIIjbNiee1UeO/R9PxWsGzhG5RQU4bl8QlFwlpwjSvofM+PgRAF93qt
HXAig8z5KJ73mLkOlOmqiQ+yYx2CVnKLog8TwFpL+TGaX4zz7FmG3xtfC7lcRvt61on6DLYViYwZ
4z5Ll3Z/hHo58YiytaYG8ML7V0RtuedEQvjMKFzBQWbsLe2X2BVqUHJfUeDiLx+XwawSJwXm3Ogh
qd8d5weRh5MIO6NG7257JsK5rvOD8dLPmGmzXc0tDddudpeSV5Zn5BvhLTsDXZfRjSC/80WrbIJD
SzUPCA/bkkEV0gT/GBmWshRAf5HTfE9E0M2RRSt7SEpL6chq9StjQqBj4XLQ+5qrqLNnVDF0bb5v
ltrfwMqC/jobLLVKrJVABFlAECnnQBRmOvivgLlE/vLEbx5n7nKWzItuFm9hYXRqRKvPptZ3I9hl
T9qy3m8NtAp4rbKJSVoDo74Z0cPWCwPALLRD9WljXTmLFimn0Bc/2/3kY/vMUcIoe5sygsGZWn/C
fkDouDCxgSHApnuHnfK132lyV5YciA+1ENaUIiNCpQjKEyYAcYReV61XX1o68YDPQs38Twhjmwg8
BX6ef14kwAh9WfqJZm1lASpD8ZkAb/iPdYJw1r8m4p1GaejLGIGSrQYiU+Zcg8KaLsyTEqX4oT2C
MZYJCvIZm0oQ2bUtadaFBZSfPVhy3IYy0Nyu9CDXoBQbA61fbSNhy6hAGh4Vl98CYaZZRsC+IzVo
U0KxiopGcQ/WxjYXXXpib76T+/S7KywXVgEcdpopUcBNEedxdk4ETMJqmxlIbF60WVGVsinoeacM
Tx/8WclIVDK44snyjT31zYL8GejrRJcoVoSXEIYizlxfRJ2Qg99NM78SP58Dsl0Epd7zWkN/zqyf
pIr3/Vq25PQRktLaspRaQ+hZZi2D6NokndnNeQvLX7QQAhV19V0FsPHS5MVgp0+8OQS31PEkwFtZ
sTjA5+XOjK1g77Y1A172evtb6yYzYI3gvqYSg32dltQ2LIWGnn3T+VznKvuRal4kHN9XlNGOGoB7
L6fwhdhN0N1Xp0LTVJM+G8WLl7TznBrf2hriONCJQj6Jss65IrPLlybC/OEE1nO2rKP3j43L/w84
FViItnTLl75BFnMnlVHl+tivFnaqcPtzpobEEuZT/4Fc01dRAsFWIoADXD/7igAX8HZKp0wFef7h
dhE4GAVNhlufl9eYJ1zup99vGfHb+PxK2icTNWxneFGdhY9X6E2z0QA0iQo47LqvBNikbs5luEgT
qdot4OC2jVyu7ayNkM5Lx7ahNjBrbH85+rN0/O+UDUb8tDDLFnNYNlDqYxus0uFKF15s215qlJrD
xgw7DRg06aJBEn2DugsMmj2dQBXaIm/GgSP4eaTP501z19qTFRk8l+9j1kL5x/h3t5MVDcdmQ10v
sPQDk1Ztyb4t1INu5Ox37RhFyZUCcO4l5wSZtaI3ltKt0I9VPfos85cilSl78t7+oGikmusWkW+u
GaWiFO/dfcNMGGZjgOYWvWVaLBSmXHTmqYwP0UF7qbACdeuPxOsmp/KhG3PwKiylQPKoV4ePFdcl
eUfL1vzwJYwoEnlDfqzoicidgr6F/Lt+lkDKanqDs1ymbS9Y31srMyxzp5lezw31//LRwqM/OGW0
ppXXCOcfKvUYrxasdsoOu8Edfo7APLdrR51i2RTf1S5jHG+EZdhrE+P9QUltKRLQQxqPcMWQB32t
iO34V9G627tlkbSIPO9Amx027n3iSjl0Ox7prwVxrJoumFZeE9K1R/HS5/s5VkaZoknMaw/0CtJb
tQKc6htzLGvcKTPbmBEIq4mydG1oq5GXgsP8d6ZqwqPuUW68LtgnoWkuh2ZEBJTWi8ZdxPMkjDf8
Y+RpvaR6FFDlwAoLh1OdxjoTQMs4Q5VfZ6FlpONgblPJDBPVtGj5qBoAMHVvRAnN/Tr/WPeDE7Dn
MZW7FCUdalISfCODIGongRBI8Kfm9DI+6cBUBZ7Fh8PfRVnYJB/XcF8VbmdisvaDgsrH1dLsFAU4
7OVZku5M5/bSLNLR5PhEaVy5MiLo6typ9aC/8vBKI71UciR9/grFLkYYivAa5WjRy1d4LBKNOoRZ
PVMX3J/0lvjQr9Io03H50JpmFkJ0v75Gby5MBCpaB2SYTze7HmN2XNlZeCPw91UMAybXQFM75I+U
pOUiA817+cJzPhBotq3GYvpLWpg9ozSfcQRNciNYlHD9r145TVoT5uw2jiZjsspe8U+oPA6GoGhG
5W6OuNUDotAPskp4w8Zlvk9H7hK78j1lG6lqR64CDoYZ46i12brKFT2WmajcQA7D3nx2smOnsVEN
1xU7O1+vNFKvpOsLh75N4e3kSmWgR3eSmgYJEQCajalJv1rQNUvRxcBYnzK6ZbLTxr+4aXPIM0fy
ihGr7BZ4S2h/wRCXz8Xy2GYOHLqNk1mEqsaFjYNxCAs4locKfE3CUfJ3ggr/WzNlYO19YR8df6Rc
ZMRrC4cRboMu2MR5TPXEsLjc+fVEhuLqiZBNT50ajb1Z9xr3cd2/p0HDrqpZ5BVzPKHeqmICMNhk
4QwNLQKeFp5nYbc6HJOL5eJhsObA9iXxAoxxMm22NLVu33nGg9nPuhWJKICXNvj1NFrIUhgO8+4J
Q7IDhiDBOT9Dj9KLWOWuMCqHOEymM3+py19DwfQHdMBxmcULNfzQ8dWAsDadZMKrZreXE5cYqwdM
Kfz5geDNfXGgh3W8MEYn2Mx4lO+kgkW2reNewCs47pSHfz16+Ia7OfgO9+ffaDwZ+OJGYnAVb7Zr
1OyJo2tjh65vPm7aw7DDu+qTNG5dwEeLTMR63HVVAliun2VYrRgpPWBDxHtko5YEJ73Unl5CijGu
AuXzpzPZ4vLWFY3oy82HptEvarZoVGfW82gVeZGUhbjBLuwYWa7/vPkftNwJ0pe+X3qbfDn9OO13
sN8r3+sbdjeZijvSi4AtG7nWr+sBEw2f6SKPR6LY4ULyVz484HCHGyGIE3NGVsikv+urmDs6JhzU
/qqYxbgTsQr3vujfd7BHDGKzDY1rOPIsw8rFJB6QAHbTcEpffxhwFlpF6DqAuyj3kNuhhY8Cf/kA
cVH3HsMgsEJsugsyIl1c9Jc8NhvxkMrFKZlVmRygqyVmuMMbke2p3elYXTvqjKPeTdE+nTLm7Qiy
eEX/FQiySNBfsxfD60e5sctXGllWA/OC0IT70aZGxJ8BaJpTCM2/sUQmtFvOi9Lvx3XApVKhjDkX
tGQPA5xNAqqjRxEHo28pNV7x87kgDOAv7HCOa3Q3b6orefaAZAQ/rDsqZbiMoLYiNzI77K4WAIWX
i8eFnNS7NAD0MzJuAWun3Bq4xfGR6AEo21w+wtznba3ZiDejHrGUa40M7r9XUs+S5BWqOEi2EWj/
LyxwHCtn7932iUpIxwjxWic5tNF9a6RYRUfrhxeSBSJ3BpeWsze3iEsI6VnXqUX2cT+MZoDZHzoP
gkvjHQaRVFuNBwwwrq/SUmww8AECi+IFRg33dhCk4tgaMnOeBFCh3oFIHiKSH78dwUXc7JYnCknx
PJ9Fej+bWuSg8B/nk2I6Oc4zgjUTIjoo3IvhiyyUetZWsk5IE5nma1TQyRTQ9+TE7bIpMiqIB1Bn
Qdraap5HBpQN7zeAUi9GKBMwK7kdeD6iDgslkcXBduMcjZZw6FQxpW6OjIyvVzDJwvebXUSce2Vf
O+nCjQrrOVTpis183/+mDYz/2/ABOVwZKxlzVSgXNxrx7BBaGxihdxMhex3bpFNQ7L/VxICXw6FE
vgZeVgqUk8c38zU2LPyT6CGwRTIkkNGfbB2dHtixXvVVdc/l8ghaUMG3W9WTmcWAuQ8/Ac4eALDz
42mNuv2QaLB3g7OWZZ5HvDUWosrMhATd4yRZkGZn1LHeZQnEzNbRrZFSPzRxWs+cY7Br+auFqGKe
gE49EV1OTntLV6OAcgdf1BxmelsbFlqrFwR0HW7QryJm0DLSDJ1v4mUWmcGx9f4XRJD9BNJtmieK
/e3CgOoJdnOLyq8wreNF5CF+91bg/NkD+qQVIjakHqHf5IflrXWG0qI7HoymGUtOfeoix05rwexT
9fSinVQkWRRPabz6/5+BX+m7Mr0qN0+A6Ew9sEQLIyhlIQ9KNAAOqH6GrFROjueA+4UcDaJwX9rz
bR6M3zmRaMpo8Sj4on1kXbVXmlWsYNOgVbJv+wWEizzabtZ1NTCtpadiKEos7MkKmqAbzXpxEFnM
zSVsWecKllnr7yP6GTL0xpeQmTldciLfHqk2YLky0Ne8+BBX5qi0aZMVZk5APxxKAeviPDMmoi3h
U5H2/Ju6ulk2KxZd5HvVzN9d/RrwNovVniZra+9KGFuEboZbVkg06jVxD5n5CQp2vAFIGDITSNj1
3jpYi1Etx86eA1gEKSM5s1Bazpd9Z/3HNPzZq678JvtAbgGWrKWkMt82MHKkKSeVV2OZt6yCla7I
4OvFMcjq4ogFd97sPcghWkzz3mgVzyMGjpip/bb0eWhVWpBaZcSUZY50VVesRH3ui8DIIraUMqh1
qATQ1+ycPm/tLKotO3vq6feTIDI3fKmANE8bYL8aHDRpPsJ1VgU8i5u7ATmHyAYf0Sz3fIu2Rl/W
mmxoTGz9pnYYFdDOpN+J4Mr4KPlECLRDmtCtLyCWtQyhVtrUUInTnNGfu2cK2JR15XhuGxprN6pU
18+NqatnJh2LwEe5+MVJE7febQTPNtpDBYQiccIgYwRQy0Kry8XT/LcOIxB9Qe++YHPwEWfGBTFe
t3kM7n3eOZW1HqCirWu+KW8EYWQiMnh5A2STJuKwOo/Mo07qNvSFXplDQ2KTVgtfekzcZ12k6L1k
YkXZXaX0anc0vsgos6DR+ATTfUpYnwY7NZm+mwNTbbJ2nTy4MKpHwJ/WhcGHSsel4y7Mo6R0KOts
5Bk1kO+t6nMO97IYljEWY5slliCVjSTz4rF/mqWJ4bqo0S0ORJVgcbvT9bMJOsX6roAPnISCX/7X
2wESRPe9oa7XTgJZ2tpZTnk5RadfvkKXe/gZIa03/y/5lFwbBwnmtWD2r/TWHTw5+ncSseiGqfot
YHIdjKCKfyil3vkajteMRdIgo68P597Nn/KUvOowl05CPP8Gu3lZ78zTae1kxnizzxK1QgX6iLPL
rtGxfMUpib5yZS8YtU7RKHJ631FEk/mf0WljPalfSHNlx93VSamsPb+Nj2/Zr9V0FtcuJ61UQBd3
15frK/CEsOKX9b5toHoj/wWsxbZBwaCcoOvZsUazcRLXQPLtLGSufXAQmc5PDz5BlT0678mEHUdj
gAtrbG4oa841xXfh9YS7mS/kkoHdfcDEAcoAxctJVDNfXdUqdV5A1uSU2lzzstgQiLxKvglSYFhH
5AIwvwMU1pFWXbKv6yTQ4ShTpV3dIIogFqfHbK7oV9rtUToN5SxO9LT94JIL7jiTZiYVRW1UoCSr
59z3R+mBRGNp+MkBebfF3j5YNsHMyoJhgmu5g0Ew6Vx0KYb7nPctEKO2khuclruQeAPvPhFtjRcK
XRspCY6ei34cjVoAocVn4C/+1IgbkEzRgGfOXZY61UUZCxBdcIYH/GasXA+J/IucEkeHvttQmunA
PrPMwkoKKCubvHxPGg0KsIKlP6i9fgCr5CJLIieR/cneoXRofYv1q9PfjI4K2Zd+9iO9wRKarcJZ
+3d0BuzbEnuGQqVB4qUU+Bly52j0JvNgVPtr5cRpBNSkio0nuMOwvPldLPkrzXL1X/3iH4uWp3oV
PU6pqkPVtylYP8XmA87n9udpnGNi03PNPiAojyMTWM+vYhzdbZ08f6+r039TDRW89+pnrgrsq79z
v0GuaAI1K86b1XE7TRySn4GRT0HF9kmW/z4XwWqFZLVJk5D2ridwfbBnCznaxGHAmNczqFWtgKHi
cIV6bEpVHkvQ69untcThBIyiD0QLz6IHTAKggjYoR0WHNN2OYB/PfV4mXRRIbVMowTFCbu3NSknc
lL9suY6nqvUxXmKq9Uspfxacli321HObKakrvmyZn/1iZeJk9/KFoo9dSWLd6ohJrzugDkzk8ANI
GFMIEf7v9QVrU2E+TpsDCbgLJKskjszQF3EjIIvVYwh+axbNvo2HGXH86eX0YznIaAqSqLeya/6F
FcdXDGYHWiHCB9mfS0xEsfs1Tk59OtwaXQhuzbZoX2eAT4ikKUJZhSVXZjPBvjAyOgpruODpgJ2l
pMhiqc3GOHH/0CHyY5i1J/Dh25N2KXSDQMN0CGndW8bzqAH2unXwe9ScnRoAeByPpjdtAe2vBOzg
38JbZpL4/B02iIOmW+nsDUDw07dOlsYRYUoXBrSugPpl7zQxImwrdQzjT5imwf9KCXApDoWwiw50
QofpIOSAVhoP7xicdXD3EetWQvmCbgegDu2Qlz1Yk+r/MfT9VLaHpJfzLh3oU0M5prWmtWwqkLlA
RanUkH9EAWjrFhGU7M1ik0BlvEj78yfGDwzqME2JjazOd1FkI+svhShwRT3s3UOT/jlGVnVCmxpw
gQ8Zt2LHT2NDK9euRGo5fuyg/dwNniDXpm4Ex91htu2syjnBlr7YeQltxboPOIcO9YpECq1ccjdY
5icvkR8x9wkiz0jSGlFNOweKrq12TkQwGmdkPfcOsACu7fItr6OmkThS23AQnVtI5mo3q0SGGdAV
VNHFpVyAIHJlvmS7x42BkFVemLo6RLKHhFK6Cprkb50wmz78T1RD1oc8kXBr6joTr0wjKzR2rjBu
xtRcwJd/xczR/7xuSpZNcXyrGUA9uykwNU/lWpExoa2pKdWKGIPQR94eAcBv7lLXM+IdVOe/N454
F3lC85R4WkhWgbAmOY0sH2FfS0a+de4pIFYu4Cv+URgpU7M1/vECF4VHG3apBFNtxl7fLo2Lb6ca
BQjGkx+VnjBhhSVTBlBk3hogP1lP2ZeEQUz5uDHHetxXU0gfZ9PzTPTGHe+F7SWxA19jxUdBp97Y
XQkjpkyLIk8ttel8ubHIkv2RdehwtHmnaMPwwbB7hHjO5SZceimSLKrjnxl3zGw0rdv4qtJanltV
59zCGCU7FWXvAig/QQ5FuZwjnKNoNYwOPmssBCMrxHcBBcu5d/3gN2ydKc1HmRCr7MCJrKmPAbKh
5h+/cVkRA3+KzSRQj5/dhq9ZbrvJxXTaZeBVMLhgSdQngb7zIQKvGP+mqYBRzcqR708Hy5BupLWX
2Boz9IOAqY10K/DdCtf0PzV88Ufm+9GhAW9A1f+2Q8qSJWUuyW9YqVP6xwAhnEbH+12DP2s2yBkH
yD2gUu0zU7icOp78BkT28X4+R7IADqawNC+TjCeXyBaP95qBei0SAGlteMU0l+rzAhl/uuZgK29J
3huyPI8R72FXnSv4P8sVa/LRr4gRhd4/0rE4yLPVt/PTRK2B2Bx7R2i/Fa8/Qv1r4FgYX3S37oq5
vtuGhyQ0OAaBDZ5ubeKpij26H/32ZELCX9Ctl2ciJSd9GqBVe22zxZV/CM3iNv92ZgEiXEdahbS+
9IovfUUmwMgRa9m9DvH6faxdkN9l8cF31+5S4ybFymyf0XhLgkGV5g2i8f2ZEs9fWHXCG4PcGXFm
UrbOsWFc58yXNNQpBQ465il7hHK5Ev1FbnjHNaE9f7T8E19MT/49lIBbl4TSR01Mk8C3PNgS/0L6
gdrP2JWwaPVEONEeue3+mLrctbTJrJJjVhcsWDfuLyRO/h4/sDul6RpDo5xl3hHvCU1p3mRDVpG/
bnL6iFNGuDLuLpJYSJRjkzA4drOoyOPVrCWqxJ8/2rBA069HGhHDz3w95JHnW1h6xesZxI89ggYR
OVBtfZIjVVE1VlB9+J++Q1IeiW9xB8tgl1hpvDuVGBPkUuT/A9+ImqwVjsfYV5QQ6+Dcw6SYfBYk
2rpJbWrOxgiRzGdiOaH2i9vtDhN/aEg8//f4fs4tB07HluX6Xwm8/g69PMpnOlktkOrKeChmLCki
gtOsLbeQPGRnUbmj0D3zh0KT2XEyV9kKjnP8khUBSpIvAht8SytEGuiDyRX7F7H8w9OF8nZ3T12B
2qd7EtZjGa0Se3eqwelMofxNhyMUiEr2Pqwzk+VjFf8huuaByt0kUAwxYfPQGa1FTP5Vts7ojH4M
636iCC/FHKuTDVY0HXosrVtHcVE6gg57gvqCChFjE8iOn7W+GgTk42vMDMpNnDVk/vAXew5epif/
zZqUljYXtHqhsisYihh8pyum0ADseMRDSMlGYOCNoxQ7E98iZLz9HR0BswUikNiX2Po5fdxBEBKj
/C23Lt0AvPQEIt2P9maOFFKcBEsBaOJWjlZl9hNvzYS/JK4bmRibWEHnbJ4QPXRr0I2FiCeDQPwG
rWyXTkgmTGHASkdVkg4RQe4cQhps40wMVkoqFc4kZ4+DXui3vB3GSfU1mQyLZPcNzkmCc7e6gdp1
KmC9nwjsixENVCFJesZbPsna6ylMIlHgPEVPECo9+1VpHyTJ3YICAzSHuFUYp/pYgqi+naWUwhjc
KLWxXP99IUMY/XKQJPYoZWfiNy9gUJKVi5w+Wt2McJS4o1nM0kEkqiuBBe7RXp3HabplO/gqm7VG
EuftuXRrGmthoK/NHL0t1537XSh6F/nKe3l8bznkEamjx67+2wvUr3L5AMTU8LF+x1eQqR9p/esr
iYMUibVd4AMUW5Bl5RLZ6YYXhQEtYVu3lxKq2GjuA1sHm19jXs9aVPEJgBjk9snbKUlnctq2NmZY
iJQ5u2M6TD2TNpTLpzA2wRm07gKkMtxx0s+Zg+qRnQMNNDtHpsGULcWUVSvtDlIT4yZKhaH3lGMp
hePp8QB0xXJ9u2ibwSJZLCNe6GZAVHP2v2Nyt6N0Ob6aJtwQZq89CengzIyC8KO1qKQvLwCQsou1
AWw6P0xJRLTcvFIsUuOQAByxNfv48VGkdvWWd+0k11qzg8ElQ8V9jpwY5vVfe5DXC3UwC+17bSQt
a9xHT37Gb+8J6n4WqK1YuBcyPjieO1bI9rQs8TuA8QvyKISLhXjsR6vzx4K49eFKKOxCuJs0BtKR
vXAldcksOcmkBkjGxij33d38loalimzFFMo9kLgVUxhBI6YCGwWFEy/NT21xYtzAbtsueeh2kD9z
LtGd7xCKS7+RtxdFfBsssr3tFCU56ffsfdm2Q70mptbgM0ZvLHT5fpgfWc3qy1kq0ShJuqTdtN0Z
PtEXhi7eRfC1SD4IU5FW37JsOq4uSHhZy0O03UtQBelHawLu9Jn7vs01nviN1zGQrsLRRpSPZNXq
N0kXmM5ZbhCw3AqUJCnyKoaCNjEVBb3mBXH/HbxIcoKUeyyBhOEPiIYuQAY3ibxvB9Rz8285H6Tk
qGW3jpe3sVOxhAs9e6NXvl88Jkk3+n5qixiteskv4ah+Mn6Sd4fwL3p7Nw9h4RSFWVJSgIe1BJgH
RYXzSd+SKySkKv74JSRwdmsjUpK2/VbyKUuKh3HDJ6LuYKCw/LPPKoCppWI3Owi/Wa06V75Px3W+
ftnh+RMRSdGyx+PEEDZTfB1G+awReRx6bR+w4LOVM0FgTShFNQlquZ/dUEQGDHvwd+8hfIC3ciEa
MvaeRgDpM8PfuUuzEHrmPxvKvFg0ztDj+r2fYVgPsaCC09YTllb6lyvAszZ9zqKvMv9gmhSBMOOk
olK5AKmNwgmWJ2EE91VypVB6j8jd45k1UQ0hFXX1MXiZeH0Tz2S68hzjMfmdsvKLqIKEDn6gE1yI
/Tov8Ivs+B5OQ2jnX8xlVpT1lLf4r6DRbkFYbH8W+mIDSDKVYOknGm4hkX4VmHP9pLWU2022ODcm
5LnKhLdBbQmkOpej+dhvL8yn5zPkJlnuKW/hkh9Mz5i/3HD1y3NRceHhe7YGrkOF8J2SAz4aZK8j
XlXKqmE4DlKIp4hpUHBNCGlLLiLNrbO5/2X12NTQQHWg1Td0thJ23GVtqw5zshFvCM5wKQ22AX0m
FQJnkpPCC+HoFw8mVMI/CzX9BmQPsBVlZbdIHdSycKf/d3fZ9i0Sqc/Ca911uTeno2bC6WZ/nWKL
Agx74u3I6FtDBhW1SC9tyfLMh6Jm8t0GHUTWcavvRvm9cU1DS2hPkwyNGWjr36pdw9EivNbnFrP3
Q7Kx/YDNF7PWnnoG9Bs3pMGkNlsZQSJVunwmS4BCWUec0NLy++Qw8yHGUEMiAl/7Uu2gFyWuAS4v
oLHALcp4f3K5xZGsBAWo3JIZmKH3nJ+cerJBOx8FMr89USdoPSowRdJ/5s8/LRruLahMfXwQoPOZ
4YCFp6e0kgq/2DuBo3P+QYvqYrf4mfOvbHbj4FDuzVyCUswVa23Sg4vqKDy3Os5E6NSmytuakOPF
xjqTv8UA5XoyEei1x2+bV5lBDQ7nGm3HYN9U7br5qP4IUtvCch7Ma7haqIRq61x03duBPgeKZarg
MSObuw7tdB9TAlbg/yH4TUtBSJgMlS7w0XwRqaNxvja7AbdChmZanZFWorMwA5RXqV91782trpaL
x/geXWm04dk/26Y/XPCbpgaHnWtIkMpvKJYOt+MU6kSW/iklDoxK3fecmloPJcYOJJhJPrVhMeoo
YJHB5FIaQYKDcatSXDPSccYRkyq71hBjbwuwcXAlBjKJU5x60/iQDDthz73N3fYVkmkFnw/TgkAk
iJSBwJHQW48Ido4HSsj6FDlXfgmnmmT5tnJTr/bonZeHArK/er7TO2H44BDQGP9ttfyV2v02C4FI
vNLZRJlPc6ShlBrSRkZAWDu9WUyzIIZHJTCGchCRMsW73jocshNhAXqJXFDF3ANxLE4idZgmQXRC
hljvS0CZGCS5t/UpbFuT/E8/LyQGpfakDZFMdChf0+pqRu53QKFsdXTB43mUtWsNHFdmgxqp+50A
lhnlxh1V+8km7hS3hE4cRnH+jmgxN1lSUFq40t9nDsL9Jy21bBzmz6o6nBcLzId+6uELq67jZ5Mf
kopHvAXDcxpDuXbhttCcV8UjzDYvMVmY6feCf70P6JeFso6umfHwml0KO+1v2UJrUv1GPSxvDyDs
ehdyL4Y9IW1vA3vA5y4IT7MuJQmZ5Ohhh0/9ZZNbefU//2Fmb7TyPqQlQ/1CDzi8Pq5FLySDWPpF
4WS351CTC/RqCzcWVjaYenwxyL4jY9OJt5LnmLonhS3bYmAsQzGbxLXwBx8I7IoBz6X6qsOk8K+Z
Yhf/mx09InFJShmpVOH/Dk4VkNGxDqhiKrdZdSDXKli4CQ+YR9MN2E/DtKB6d35zTsQ6arBx9GS2
licnKKy2GqCe/B4gVNua+kHK/GO1LaiklFicy1fhhy3WKIy/lPtlb+ZzeYx5J9VghFVbkZcw/B0Y
aB1aqwX/k3BRooOoUn3sIoe7u4GdjOZ2ef1SmWT9yZRiT+2YMfsrE8cTA2E/H+1MwfiO9PylZpWd
GW6DB8pblQ8ZGLuRCNYnsCZprk7wlQ6rG2gQwHOzEMjo92OaQ8jzqirPY5aR+OfKdQRX8x62rRcO
9h0Wf/EY+TJ3MfOS/mAhx/VaRTpncJu8gA2JQK5U3kktsJ/+vuf4fYZoa8qwDrXBZgtgks+/uV+a
ZJEDmtbxd7y63Jrrs878rjh71kMhE0/r8gqYoVv/sR7bpNsBfSCc5TnlHd58TLqK3dJ3cqsD9nRo
mdJ1Hu92fyoyllSzPjn7WZ+YIFnuY0gAZGCNthEgocvigTSxJErUVTt6MQpYIy6P0OtLLIeYaZz2
fF4TYAte6Rgv7At2I2bshlC/6W6ulgpvWFrs7ynyU2aey6Af64U473uWBNdDRcAaDrRsUdK8gTnc
YqBx9yJsJZtRzYIK0RFb6Up/adynes6Sfkudvur9Dc7qlUh8VCgGvQdiPgpiYM3Zqj+FqF950aN9
6pkqiQPaTWnaRCPaNTRY6fN0lXV8faMiGSsKRQ7TfSDgO1tMg4bWFuIpkwCvz5/pVLDEtyjLFWMF
YNPJdGIhoRZKtknmIkgpl9byhv8wbzNMPmUtNqnqOjNAbhgtqRiRy06abDR8ll0Y9ERPpNfV5WfW
59vEZ7d1uH7+N3yaNduCn59I7ih1iuDIcBARvDWMtimn5qFAurswPjfJL85KcYfT+dXEJGAeTSm0
p/Qe+dmOwFSAcuRn+b+nNGOVtnLa49DrVhYqPseiJ82lJ4hAQd9lZuLbRJu6+aXiR5x5BGkv5YAC
HK0fEGlaEXqWWjdvmekrczskP174WfGPA8APu5j7HEwwhmaGTmxJOjY+EVws3M4fkrh4U0mD/29/
aZTyDuN6EhL61Ycd2qYsREgSPIX7ZyMiHcHXSmoRPhH2GGeAs0A3OhkzimWuvkoGb21YABGrPRtR
WDmvHjFrWZNZRjW0jOEic+2qm42xXhZFx5M5juEmeG030qNH+LWwv1tEYEAyZ7BJvizGLpzbn7q5
xIbtVLKY+8pp3h4pj05qMz5TQ99ThMjWWCInbUk17Sz+tY1RTrQ5XTkaOoXxxhIYxQGtyjPv7Gn+
fSepSpIoQiYUrX4pMRHGi5cIZmXs172KB8qwaetGHI6T0Aps3FhkOzFeBI9q7rc1VbHOBPIglFOP
QssP3hC3+lcD60NahCknmiyk1FkleLjzVErKkZHn9I5ev1tNL4CJAKJ2KUtkHjgYX7f59Qh0Wkz6
aO5FYjTOFsXgoY4Gcs6J/lIOlGxDa9FuCRKgYoYJ98XfHeomJvibsvV2dF3VPJGmGhuhtuFSAg2S
P5M8Cxu0fyojHj9z1Qe0f8DKf2PL2/2D95HeQ/LRxet7ILWbhB4qsnkwAzbU6YljWT4T2ORAr/md
gc3StMLmyHe5gc09YMldD9beqH4+8kHD6ztJFChPkXUA64mpYtt5RJ5RnugLWQsdh7iQn84QBja9
JbkwLfSBCfZSFxleKx3WPbhg6NMwEUzNvsDy4UqJibEG490D3Pm4ZiXYlL3XJxagYfEchkfVnQhs
ynPrRP8NVbSq4jzaG1Xj48g67LzFTHCHET+zOJV4EiabicS8QyOiZx1i4JY3rwdruxb57Me+I51p
Lj409sRuFm2x4P0O6anh+mOPKoZ4pz9diJGuWV5SllBAkXQlKws9KP46JRYaqs6XceySFheKQigX
QxKGbDmcj7TUHrxMGRXr52acB+mnk19UE6059Mh5nwR6BnisNpifiY/F2xKOrSGVjo7KHtioy1Ab
BM+llalP02E8AVgon1NSjfARJoJtr9IEBG1R4agiqmiuuQNCkfcb6rqQAgdAmQV6LvwBd8ETFT8Y
8IIeUH7Sggt1lHZO7VGw4/CO5wpaEo3RVSeNKdM56i95JQ9sgcapLUa4HPcFLKGE9kDaasHSr8KM
yG0Mj8lfA9HZkFzKaNiR9TVMOAkg3QweDl9+yz5hF7Lwb0j5m6F76qDaqVWRjBBay2NXwoOqIvqm
LjqmISKP/wXbbCiPleSzupL6skHAOJUUiyRyxopTXRt4vP17XPf1yIR4tlT6DXo87RGTk7nIK6gd
J60jNv8DIu0MdW9/PtCTabKj0PgVHzaovC8ER4ryCGfP6g5k6zmq+2l0z0TSsDYnpCdaetnf7RBM
TcrRzEIgidcKDChcZAGg5JB+Afkxsjdx3oxrtbwMIdGqPJlk49FXfBGmEZgvRkUUXcmgM49um/eN
kjtYr/nbkeHLAuxNhR4Yqy69txlbF3hiTXBi5Fhgk5QKwsrDbMDI4g68rlWalCUHu72mBFnNvUba
FM+M2VqqQGEYy/Wpehq0UjNik4ZY9o4/Ds2q9+9cbC3xt/gWabfNkuCj+/Jy5Eq4s3GnujFENknf
BoEufbH4zNUyu6wbbnASprLlpnss4ATQYrpfUsaurFrdOOC+zUBLqMKiEgrEwbQv8mhiVrNs7eHa
49MgLX0kFwgXgLCZhE4aDR+F92PlPDQQm2WXubW8fywoaSVgnaBnOIewbyqXlcxHtmDxM4BTiWOm
GhyysKQPOmK7PFfdulB9XoUivu6map9lUTsWaC/+iYQUjlFhjq0UM79YzvDi2s0lRdSB1ewtFdCF
2fBLTFOpGmI2APB6VPBAs7eNZZmuoXLI7/MbXnIIC7OpFci7A7K0RmhCxH8vDEMsiQOHGL3PkBBa
vxFaXwwg1P/MndAzKvjviMSZUnkpXWsFCxDikWDDt5uYspBBGNf8tboxR+N8l+FFpp6xDyvSFuB3
ttV55fQCQPeVruuiGXIfqFb/kFTKvF1USV4/ZELZDkVCvcqkA1EW5wHGtcMQqL/QZqednlxDmF/n
x7dvZ4gdDOwcLusYV4v2CH01vnlL6YeanHsPEikCxFbB5KQQsJiAongw9NUwuzoMar5VZRhRzDJu
Ki+xt7HP4KuLBtp0okKdFJv7vbD7KAUHw5uuiKrovc9n5KV+Nsh0A/EPdSLWnZpM0s8y6Pm55IRA
PempdRhsgakFP1aDVs28/r+jnai/jmztAU6bL1FFNqOfEjjQs5ZEZacuPEtlJ7MQd2HtE6TUzIZB
WY7CM3lI6xtsxrfqOAiVEGU967Iby7xmTVyYgaUlYgMzEw2+afX+TaFMk/9+waXl9dQvWGB5l/CF
0giOPIu1eWzBPla7Z7+olhbJbdv+K9G4p2/egWXRHUzYy90UfcejGy4cF2LRoP7m2/L9vSKKCkFq
wSGYdpEfr8b4dO8QUXJV9U7jMvocMmQavnILPZ/SNfj8ts5QvjAdIRCLgzh9d+L655CSR3zEcGCG
4PnbqSu8Q5WJhUWD4QNvXHrGSy8QdltWbS80viTX2ouf
`protect end_protected

