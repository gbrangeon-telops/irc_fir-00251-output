

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e5xVIDBGzQkhDoQ5sfeAF2q83P6A1Z/qsmlSYQJY5xTravGd4CV8IrniJyUa6zNomwm8ijfsSBDZ
3Cv5fk91Hw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JTncam9YaU88Ye5zsiMSZerKzQZ8ndV/jFOlVBJ2+1NMrth4ym5MZgOOJUn+hqDs7WawEc66qp7n
dAXASYJYn+qFnCtyUAhIyvGYbamoaDWo5Ex6WN67wq/uxVFQHJyQE9mBWmFUuyQbfWAxdn0X8Ddd
XBKhuVWHjadjfvTndGU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WysH5jibOCiuNoaEF/J6UEux/f9qwkqszrQvmOG1LAQguVnzJ7+cmZtEvDLaeM5SMkI/c6AvWtXW
QAEuUSUqI7fc7s94OSdoy/EO2eWxzu/2PZr3+Vm/RDQkA2VgY92Mk7iTSAe4nvupzjwLJJp7MPFn
W0Qp6hutV366SMmocbalqT6lFUEm3BdJRb/waOPaQXsiK/eXFOfDC+OkXBIeDSI4U6bTS5BbTI6J
pFf7UmKKQ3+TO+1O/Q+2hW5WOgJzIUFjgYlL/k7HV9GLoiTkFeWQv9D4PmITDLLqEoJBQEH042D6
w9tSjJ90YaeXyJsQBc944KHiROaj7JIGL9ptSg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HfnNrIheX+bmcZCjcmnXLaiCn2W6T6H6Dp6dScskVGNGAylFhqrXsMMXHrPiUKf5LFkT6rGH4xNt
DnPlwzwiCAkQpMo27mNuJmSmEL1NZn19+z1IhIkgUjJMK+DU6V8j1HJvLoBzdBKXeOfEsIha7CfH
SYvgpUYxukUrvYeSdDM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FcdqosqcEEFjwfToDdg81IlS3kR13BUL9UoyGE7K0tYyJxwBRWvuEZwjlqyLvEdW74UEcoL322wG
MsjKrbrYQdHQMnu0VAIvQRAp+YUu8ZY/Amts9d4uoKQ4ceZKPNKKjhA2gLCTZlClOnHdKjhfnFhg
C4vFlIgGFFvgy7hYPvMYgUjBeujuUeMJVrfDQoBe2vY01NCaYs8PD38+MZrB1yBWXtoIH1Kudp5s
6rfzNC3iiU875HSyCH3s6Fgf+5qupOBLk1FOGYXDOgVB80WiCFsXlSgDSubN5g0HTJQJ5d2+rdH3
3+ADIpk9sqzMVdE2qp7yCA7kfUMNWwWOq2rtCw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15872)
`protect data_block
LRh2UpuzbmsD+vOEOZyz8uJFOhABzlOW9gW35QEuzmow54ebORuffH2dmwEGp+7FjQ/qPczNfC/T
M+lIYWGus96G1MaLPHLhF7ux5JkRWXG7QGPOkB0xdqTb2ZZ5R+uW48dXEwksjN09fGdiOPvtof1+
0IyiXLoSzm7R0gRtrGE9/Zy+Ylw3qghy/XfGfmGyLgv4C+g5NNYLr7nSx1IDdnrWHqHkOdcnV3fz
SQkMhW/EZqgF7Cw2LoZsY0jOkmHcq/9WU7oCYMRxxEONd8GDDLuK1pLtWj/2+Iam6Gn87D4KL8X3
BhpWqFYRXrNpO2BSpsCl5oXPZmQa4aGbiTyHAvm9A8wd2eYe9vW0duSfouvP33E+FTs99defxDJl
IU/DEzsVduVqpdrtVCV+HLn2e+GuzOkYwFbHbM2u6v3ynZ1huroHVGEspYv2DLS9Tfm1TxrP1mUB
m7PM+LBuKszn2YeWhMNckpD2JR7PBz3Dms6fC5XvN9pQE1Y3goNwAK/QkWICeBuVNlYyhUvoRd49
34gebpDNrK53uzmfmUwDBCWPFaYc/qQDCwgAE1WK91YPAWCpC370+qFosWYyAjxjmNqh4bzkRuck
DQD8LWpufQjadcKoraGmdlRPRauT1SlV4bT1I0Oqj2Knf591Na09ND/HdN75UjL8AKcIakITIA2F
AIpNUbOqk5q2M1PENt18sRL+BiT7GBM21NvmPFyZwad8NMGHcm9EvwZpgO6U0hmjhi2LZ/Mu2y1L
vtidWsZ6dmqnHbiGApBWWVqBJNkAxSpMa8VK7YoUWxGOZ/3CVH7/Ld/6YplrKDBxExNLRy2xhtcw
ZMHNo/VGqoFLM99ZthzZUGDJTHXyWv0kO6jHiKueVuCRBchjExVfKy2WHj0VZoYXoD3Nq/LTwdhf
yPFpuSPkBynb+w7dhLcA3HADjoOmBbgHQDpdyN+6w48vY/f2sqBXqrcOV2McMay3MCbuiPrDqMgl
NbAvwQqrOaZ+TQPM+GJx/EyOhQwRGH3XM/PngBjiIAaZDFJseld9/I8LNOhp5pTZgCfA5+/CIa0M
ga6/R3kDiUwvZqZp/Ct1uhYTfcOzTRTtD7/WTla1eKofn3zvFgp3YFUBspq7ZdGJHGLn5G0pAP6M
zjLBg5hJ8t7t/b+uZtMrEU60vP5ZaDEgYFe4lsctWkmA9QVDUObRs4034QzLnEYDVFpxpJpF0viZ
hAZA6aqBmmlH+S7jMqlQ6ZcJePYKipYV9r/6RhIA8mv6/PgGg7PMIVa2oKSyrU64wkqysTi9Bzke
o2kzai02LmEwmwnIahS5I0hy+jbLL5OgPKpJM+U6kuG518nkmBLDgUpCuTBo1cysCtYZIjhlHfaK
CSoUkUcIjWrKrMdZASKXbuWiCnndC1DzAjRxSjszNVJVV25URd3Bn0vF1ndHO3D6v2Mev9rDMAiI
A8NQd7I4KzU4z8N6GvSvGPVvOo4UeEkRM7N39b1kF6ex8XlaC5y8up4+C3hntlZj3rfPvmzTnAH3
Wy5uaaCclLiYK9b52tUf5EnNmLgYeA6ZnZ2qjnKkInJR4SonVOCYBNMK6GBeuFBDXGYic2iGiNAN
wBR9Un/FMpqpa0lfXM1w0J2NL9FOzuH4GZfe4r0qOshCQRoi35KukyJ/GjXrq7gA3wXIeWcikzIa
68CynEaubQD5NqcEyQoh3nCan39r/WzUnD6++u7Lrs+0SCfCWV6pN4+Xk7/zjgLv7qAev9t/OTO1
/sNUz3yU7+NZxnDozOw/wfbSVvGqrOqS27cXLFSipwjg+fkLVXMWmTikrj6rHoC7sNd9YcXgAMtl
FLmomzYQ4iWGcCF2YW+CDE46C2x72oLTMzl+DcM9mRB/DywljNQjjyjcOB/NQmDhsQ9OYLekuNQQ
cKv/6GEj8KdWwLBfu2mUIvjtgHcmGTIC5ARC6F/CkfKo7xHoGT3X7eaCulj/IArHajD1fXGURrii
nDy6xBrtjDOOI6au7OpRzjdvLoxspaMR1d5tT36qu59rTTw/Sv6GjfE1d1uWT9JC718DLOvZknzk
xoPNgdR7t25xHIUlq1BmydV809JWmqB9TQVP/US5hcWjjwY5361FUsMhDsH2T31QFT+wLN6Es/mQ
IYFSBh3lzfoDRzpGKZkRaYbM0QuMLGjEVeDVcJxtdkioBKSugxuh/l5+P6NX5zSo4NpeEqx3ajyf
FoHGPOPW3cy546yRy0YYITAwx3RR/pXWGlt12Q2JDmzv+Lyq7h4CQfZie9vnk+C4P5ZpgK08Jjlv
8r5/aVIlMAbSFiI/kZvkWmOuKeVsBP4Es7lhSbt8jP82ZwLw8c+WUaI/sVvrMONNC/23in5sATgU
U87jgODrlP5xCwuZtPDkrCesIThReUpUH8iMzPtmTY19yDNb6EOqfQt1yiX41BcedOonRqKY8RHa
UuxkfWKL1gbgTAAyX9a2CuK3N7nl4WiK0/KEqM83BEyLwlWEE0z9meibXoLx3vg29RxovFn2Wnsd
dSSLJphKvjeuNtEbIEq1NJaMtEdGEMW3C9vLMkWcoQ+Rx0k4YBdsOHqIiytrTtXvTLHLvSZODQMr
kqFxiWiCRqeUSYQLQYfmM3z5Ho+O8Ek+3ePRF60YcW4PyUb1GM8It4SlaJWSALQHXGB5pt8Fj4tJ
IYGx6WyfRdEdEELEFfQL9svDRaLfjHPIUt+nU90ZTuKJCg8ix/9o5+C/q/hXn+T8Pw8h2jqPdJny
NIPrnZls5l/92gboP4U2epYK3jjrQ3zbEBc6OYOFvIeMRdqaUPdbZsCNWEYeCuBJaof0s53UG2Bt
KqYZ3B/rv1/n6yJkrxXXLT1fK4Hls1ukpHkESCrp433b90LX03F/9MmVuYb/PLkZFFuV10DQjutT
bdaWWWirphlZeohudd9I8XKwIxz3gtRuJdyUDe6c5Io8LVIeMcEwRJ237shcOrHUwctjRMT1goYI
nixKw3zWmqyk5/WcjmfWnbkSGJvV70GcD952zCmiVlxUQ1IfUrlE4s/+tjtB5zvKlhn4/g1x6N2b
sxdmRQpvxBzuLCpwhlrar3nyICWFATOG12Jg8tpGEAvblIPstmyAHjW9GmXne/cM1OrCr5QLnV/Z
+ra1H0aeSCODH5QkGpp5ppEtrDX2yGjPEVJ9TpU9olxlCeXTYpcIgXDpQqNjdqxVxFX5rYXXgEYs
3IOP9LS0Ob9VTmwA2ZReEIii1LGOdqS4y32N+OGaHYEAk+0FaHs1O3eoU/kll3HWN0QBxMlFRyFM
BpE2iCA9FL+Mx8rJxRa5Z25xT4punzIy05glI9N5A9NROABOyb9xcUQghoQtvkDjxP5f+zf6qoqz
0YpeQ9owai3qogybI2Rf5/+A7ESsXER/jUtnFW3CCztU9zO4c/Z/HNjTsEVOxWZKSj4V4GDWt5bU
wXyPVv5NVuuPnYtm39p0GA2zZTQihreF/D2zDH6iXag7Jm87EjIHQ2bpDNI8UuRJhVa5BDn5GF2b
YhotBVM9kYFmAzqM7nVUsjVNK89aQ/Pa+88QSOv5pcDu/M5TOt/8G+ojdaNtfZrMdnAVuyxyZyhJ
PrhrNd18XHaQCJv2OR4Ypn2DUzXeYYErSXFjamEvhFzP9qVsr4aM+QN90v/zI9TTI4kRnMTNmQlC
KXieUJQvF9ku8ZwrrmKriExHVZjqEkeyBHRkafCtEYb9yO7psFnEpt/L6eR+QpDkJnW9SdXrt1g5
QhPoHRzs8hNwhcY1yPTeddoXP5sdhhX3j8eAaSG+5lDkcU+aHTkox0xmOK/VqSvs7YH0Eqj5gopA
q1uNj6kXbou3uWGWvMDcnQ0I318LkZ7taOIjQ3qMKnVhNtR7/+tm8DKt5Wa87Q65SI4nfrpdWR6g
9dA9PWqbRWs96y5kaAJ4VhqpVPSxP9bG3rdsKHcNwLYvwifcwxw3xiqBIhQaJvSc333/uBlVMNnV
ZqZRItGOHx7kBJnfA0bhgDuhWGRe83k9FNV724Pfv/WDTc0u6EDHA1q0IvVEyq//nUOOcK+uoMSu
MIdwESX3g0lCqG4ynp1XQoxFV08rSvdvc885Q8qlIXpvpF9kbqgHSFEhZp+yKyetcYN2Yd+bOjuW
v+c6gM+fs+fWZ79omizdBNziEDRVPJng6Ipca9+oJSb8ocaCmJ00bSoZp6jYmseoDYVG2mVYUqir
MuQZTJ1Mpsz53E/5RjnUZpfbfB0KNkVRIxN3/lm/08upiOPC75y5l7+O5coc7o++PK1oU8KgRXuV
9zlIviAnD3dvn6Y75G2hHeO+BDD2CpA27O1ferN7Qh/8J5DOHXeb/5akIJNv8VLBNKtI/5a1VyO0
H2GqDpfoaZOy9pXpo4Tf6l3JJC4spUQE6dOx4EEabNPsPSmKUrQSacMhKi8Ju3CrDwbnGmGIZbsq
rh0ThCoIviiFbZdcQZB0Kqsa+R7K7t9I6a4EY4RM6WbH1uLjZsFbIN7wZf2tNWuUnsHuhxDkXIvB
/R8zQt/qWj+hAZV13nptE8V6RdLsVGjJ8oM0VBEkXSEo6x4PLc6SXAr4yze912vT5mO0oYZwACa9
ak4HuJBS+iP3LH+k9RFs0DX6Se9YalZAXXnwIOXl5sxsZ6+IvG7N7/CrkxbWCUMz0ICWk4/TNfru
TZMPHZN+maM/26AOrPuqOnkkXnL1JekzVrKkIJXtscZ7mv4Lh4og1x33QRlV7yHzKdDKepYJYxzO
wMNA8UBg+g2P5eQMOxsj9SMCBEScLjmookYFPzMQJFPnCo0dG/+BcXUC9rXmhDnx+u/qIhH87YmW
3A0X3DDUSV1q3zN9HzCHveOiHJ9rYALLaIu2PZLaggguVGkbaH0fkyg+FjhkKgurV2Pa8+wmmABU
quLam9LZV6hFgeakhFImQuRcDgJvw/xypgr9Vq6jk4D6Re1hITSa7EojYFAYBtVeptVyrw7UHwqc
CZku0cTotrX+8pw+QsRSUDDCdvYhE/w8hqCCShPaz7IztR5jNCOAKyyDE1hYDjguYyL+ZhiyJ+pe
ia2F9RxdG05rLFwauXxjsnMsu0LWQe1O740yI0aOHQQhU1BuqzMRZYlKjlhRVyfG06RiGMba0UvC
GgNz/z+fS+qRRro8eU+ZS6X/LhzmtwkjL1Pya0HGeHvBXoH5qNkcpPncO8NLRg7QsY/DTKDQeoqk
Wo5vUJcV25A9u8R2US5i+Es43s6E0TS86dYt6kOJQPPgqutxm+kESjkBFqq0CP6Oexj6fPhRUCOR
qweG9yadk6aouqy9KMrPnEE6XFx8+e53+8nb1bcNhZwQMbY1RVGMtb5vFXeSe49sASyj3uYdwB4f
qmA7MlQpMOjJTBJufvCJe4ImMJVlFOSKZPoXin9TDbo/7Iv7+85X2U69iMUaIdCCxMj1JendMrcF
29my9pN7kFAhcKtPfgNag7WFlrHA9NPaJ09SC08NATyumhjzeue4ysUrMSV++py64dBL+w78/kPg
hrNOtLH2lkeADzRgJofs2Wb5Hn8Tx0q9oGtXEr/DEodoPRp0iWapq1/bXHMmk4Y239p/vm2ZEvAn
P5i8MPSLIEbf77wZv9DzQDhj+r1Wp9DQrcQ7cwIj81muNcpCCj+gy3eOnp7//ytYRJJIwdeoKkjJ
NF8z2wOHC7809ayKHBpelN5o2bcmrunvArdAztFlh1ZmKcpsj9FHx+12T4NMkS3mzgQD4yi9FiPY
MxJyd0j1Kz5W6Qimx6N5ic1DzgeEVa4+vpHztXskQuz+AJtDFeZrLjhsJVH+fzk0m6uuy9nagg1i
J+w8Ch/EfbDy9EhCYYxj6CzYWtj7QesamLmFcxmW5BFs9g6AI5JoLAIQDjWgh5husfyowFf0MazB
wN1TVoiVoDYj5LDpW+JSAo31TMEMphoD+4deioUqlKdqMI4LrVgWlM3ZjGUoCmLK73Km+Xv918p7
zVqtcCk+toDBI56fi7Cg+5cHPd8es+7hRS8Vo1df+07uJbyKEy/TKqS9DpkHwaO3pTxs2mZm7oWE
OHXl/8jSttB8tVFJbmtpSoiwPGtiUx3HF7VnTpLInM1wcDJ8zQMTNiMZ9PA7smldV375YwrVgQp1
CnVWc2SVT1KvQvxlVab0eCfTRJrM6o1NWqanbnkjfh2BHe9/mrH1S4L2S2cGsgy4nIuN3lG6C5xJ
J0O4XitSL/mtm/4ZdY3GU7AtUgGkN0c2DIs7eIrY+ViBwKj0kbaXbjvRHmHfkcTziiQ7lLmTlD+2
hRJOQB0uTITysoTPxwMigidF7amH53IhUXItA56xf6lB9ON4+f/3nzh4FsARw+EUs6IOa2WQWkqv
ER6hw1c8SPKoLN+Ya4XFSAnoQd9IUcoEU/V1CPPdssKx8ePzf6OQX6833kLlV0BCXx11Bs5FFC7x
8flXXhnlBQ2c1H7++UIBU8cfOh5KzstUgWQdWs+AWNzOAJCFUymwE2WPjsp7q+mScIduSi3GQ2H6
DxI4dYHe0xUTwNy3ASOYzq3OeTAbdlcN9CPQPxeJVeNal6cJ9NpE+2AAWCivALKTeBqjmXKtkZSJ
+wPc+j26mj19lnuVbbqZkTV0ZBE9NDCr6AFQugju/nVb6LtlkQZMvwbrINUQJI19Zj7oMSe1CELa
6mjwilEei7tddZcFI9tcg8kYN+Eq9B/3jwBbdbrUAUiOl1LpfNpxZFfGwf8Kx2bdScxrvpm5/PF1
fW26C4xCwEsiRSj+La7iCxbA2YsqgHjS8Gywkg6sivKCQ10dLsBwBLRFHxpWPbt1dxu6iRBS7p5M
489zSrpamBntsrPRMVUIF7SQtvNIhomgIU3rjmlis69RSTC5pi1GC6PivbM5LCcCob21aAlPQzwe
I2T6B1chD4ecxJU2DG+eI4T8ltBJn63SXMMciqFORSSoAtAscobugZwahKtpN0u+7QkC7FXSW72q
VBzGaWhiAdx2QZfIJXtpQVpV8a1LuJuL/pFepd7ITzpbZXEJunCuBfBPnMUoVOZWaJydL1UxRUHF
KvgnqMU0RxL0oT2nJwI0Wz2sY290IAjKaWUiv0/hVzFpmcZEajdQ+27qUdCstSVJZxu46X4hDdu5
GumW5OZ21ZihoH3aoXy1C3bfmWoZ5+6kRJfwfClPCQpWz75FB5yTGCQjVZVy4qFtQtjwj5Spzads
fH8JlKChIM2+1FcGtybLA81vvsqos0+5mK1+zIibdrO/uym8B3M/vFEKRz+q6V2xF9HjIegOSn07
p620UYNPLmPLQgjiK0Y9Gv++8epw6xRqEvVBzEtncSNEUAGGQ6H0FMj7tr2eDtQyrTUdA1HgyCCx
9VNjd4h8lzYDgTxCbQqBYG6trfZj4zGxzXsiy6WGoxhAQt1EC1gjVSotFkxUc3qXycOl7nVSiD+t
iaECakbpz2sV8bIa8WLqBzYCk0ETbsMdd8YJGTp6Ql1GO5B6lCiy8ZnaGgIgzB5igTWwKI/cfNEh
g8IuuAx41Um5aYy29RiDBNJYLHACBHqNbRqooaxvNOPzGjSlgkniXeQ/NILlfsLiTN7ho0+/gzKa
zi+RRyYP9ZaCS3CL3kc8MCWJLQ57Ityq9u8diCC/Ko4wtWLy/8sfRV9+X33c6UpPn6LG8TWaSluV
MO3mWWqP6aCGyxZfMaVE3fxDoQixYBldXJ+BKzVVsa0Uyw7lC52Xg5vb2q//5hMxk+qqSDbmRJDS
uL6SZaVzkuB1GDa0l3NLs9w+vX17Z2q0eG8RqqfChMDkZhDtVOZsJPPIP8KJ2FEpHUyqaCWbuZ8O
JFk8RqbhLg+2T4OIfCRZwxAvNwcW/16aVVdjvVHhXqSMr0Sd9cbMDUPVQau87YC1b9T+dhMdKZVn
W8roC68+1cO7K6nZhqUKce7To61V+l/Y20icfTftVn60ZGRx9LCbxaH3qnDV29Odc5C2rqChfxEa
WCh8z4r8H1QrNiwbcmy/DwyZQnk+EYc7kUaDn18DJicxA+GCb3SzpFoZeKC1LcEml2icIlCI73lU
tOwlQDvbmcMcuDLXHVHjvf6rTU/ikYg3VFiDGRUPDMIXqhywH7DcWARzp6N2svI7djkthTL2Bu6H
htH73psry6d6bj42KrTc42aqyGENT7qSjauHHt7cmrAD4u2PtXZWb2wn63xQDe575anSmRvTyoNE
kEzB4mTUW6VFyKhx9vTapWcHK13gQaBeG0Owi6cRlFfr4NLcx1namAd6qIh4uwWVy6VPlZPhRy45
uSljPBij6s0pqHsnm8EoH7e9Zm3vNjnn5EyBDX8fVqonyHmSsdt5dIsw/ntZyw6u2TOsf0MLxVVE
RHiom3HEt4wdmYBoxrUB8jYGTnC2w+dEF/Eo6wWb5Yl0tdHZXAPYdbNWv7wxvO9e+SFqMU4Yhd2n
trT5VQa3rj1DVjxU650LYtpRilPqHxdkcyOCCGnonPm3nPNz3Y8K6TbOlaQYd1LtXNyxsO6YcLUH
83ZGtAWE2Rbe7E8QCcY0SidphgWUdxKLw8jMxEKXS9zaHVXM6vNSxKYzwROpn2DHVfc6RjG5I3F9
LMg8PHaxI3dLRsiAAgx3gOr0019mpwm6w4YHWlKDu6pi2JO1FPl/kEluizYgfmSZJ5xWKW6x62sS
kM478hcPSp1SzBumDCNghu21gEqJflgBt+0VlALriW9sQXB41hbJH4cvD0E+q2ajhBic9QDK991T
0R5v5tg1jU9A58aW4zrIzDdcbNnocWf5k49luhYGElFVn+nI1WnSL02fZp5LS8pN/x+b5sGJxQMb
RQJMhBZiR+lc2q+K+BswShOupsiyQ1Fg+mH9BfByntPP3647v7VNs1mWy30iRqbB4ZpYYfNi+VjE
u1qGq8LigLysxPDvT2lTMz7qyj/hzuuxK+Rr9QyYzxTUZVC4t7SAs3KwJc/aQpi1vMXto0eU1qqZ
NAecXHt6A4ypmw37zDvnbGwKYNhM9W1pt+ZyVZiH97VqsyfIdXU+Hy70rcEc+5zsdiFxPF2lEguU
Xyx9AMli4FWMshb3QYyL6Mvwq+aJ6Gk4hMVE0EbZww01a8dsbo6sI5P56pn4uP/QPSvYtIy4zwES
COAbS1UtCsAVAplsNdSzYiJRG2pYrqWPO8YiFWO4LA3At0jl+B2am15K61cxIsviYK0klksTpdhe
Sj52/TqJ31Q5etQM5n5wkJzO3UFqW+2GSTkddT7mYHLrHLReLlUFtN/6Dy/fXPCZ+sMuqUjj2neT
d6cTOWEkIGWlMVmT0VlmSY6vuLm/EXTokfXn9shg9H+WCttqNUrCZdgEw8LQzAAfzaBC07lnrFCJ
qrZBqyeEBJq2DaOdmayV2yf0KpnAHhq5vzS7cQ+f0tv3lhgGokd2/aRA1o5dgpSoP6yfQpxS99mO
Krb+dEikLdPXlEfXqpgLscgVUMABPf88EKjLX+b6xfCHB1uJJxXwLEuucr4Nk3gR6w9Vne6+AGv2
1TiL3xyHey3iAQfgFmmgmJhGZoGBh+utLKVfZTAFkGNDFrAYCKjS+p1u75tRKrYSvjpE08QbzYw9
5ZGrHzdTCrRdA2oZ0D/APT9RUgp7Kz478pGL/qMrZUyiWWJK4PFZ+LZDn0QSCYuEUt+LWcVmuSZz
Eefpk42/f/0qpBJoi6iObEN2/mTaTb8h5Ghg3uPbbIBAqFNuFBMZju+HkBj+yTvAGi/qYLBnkSaa
oDcPbWTpKft0LluoMUw7RT8lutNeOTuy0BDH6kKa9a4A0Ehv33cQSsDxVkCWbLD12gS3ebiFJyfo
Up0taJotOPs2V/f5Y6j7fTZPW7yxvF/rMk+mqp6SMnnE07itf7lLVdb1rSNVy4q3qm5mMC6NnCOf
AGZhTW839zFTIukGHLE33W8solKYanEdv99sd9QNLxktgJDDjfubJEhl8zOUZ4Od8EYt7zaYolaD
HaxVWLlpvdd7lM6uzW+kHlmMHIyrhz48DlSgB4Drw14F4mUcYu4FDRln5hAzts6gQuHCEeDZcnXK
0hEUv0kP5d+TXgKvJZId2+yBe4/dTvD08DSognjeOXYYRmTaRp2b5mRe5Yv2YEIWp7T+OVvdupEQ
33WsC+nZCUNPW0C3TTWNU0yNOli2XPw3ImNoDgXuaph5WmWtpBoan0j04bCVPJGsMu7QwEQ7l/hJ
xyfcUbzLIPm3aRhvkKNKOqoOiAejU9fzA48Uj4FkkIA0MSMhA5mogLxW9U+pTAwBm9/imSHnSHXE
7+lbcJrjALAamW1MGR7TOoDUwZoaM6yn5I2IFrn52vrlKfjz+pWJOYjkiVGOSHU9CG/dBWQSRP/I
UHnMR+QQB9ftcykjR1iUaO3Oyw+XkduhVarQek+dYXJNyS6b+3Wlk23SL8KHFekx7XXjgAJUSLN9
UVwzhXw/olsqqydJxLZqodspwb69nptYstREs6va+/2DXIDs7Vz2kpUufF4OidflwLlrnrQa8JrF
76AvsPKvIK5zq4+Egq/WgQ3a7F15gE4IRxneVk/a+QhO7RGVgwg7+lUgCSnrnnmG81o8Nv21uNkd
zIyI9fVONxb6mAmmbZVEIKjQIMMYWa0ImGP7TioGtkgKo7vfxY1u0lbnmHiRpmcxYoAUP+34CgUZ
xNyI50ES3Ldhs+8bvfkAiRnkkwzKq7Mb5BBZOW0wZFPtitdVYGPvbuNniJeaaVHyqaxMHMnj64BP
dON4EWUPFvh9Ll6LeurEoCuPOgGizZRdq3Arn+M7wqUu0pjdYGrV0UgWNio8E1pi14YQFzkISUcm
/tsUgaSkgPZNHOwqaLb0Flup/D0Cszlo+gjLi8O2MN9cxtE2l6YtneymInFqZGlcTIDNPGgJMs1C
ryMmX50CwBhKovesxH35aKMDcn27mHz8XJLFqNC6ME4N33BebV8iMo1hdRCK0DMZ+b7mHSYL+bLP
863u4Su+h1GswEVaVWx9X2YGoFklLzXiYAKYhIMRNX1+RX7pGtv4zduAUN6P/PW5243LcWKj31yv
M56SZaidUBkwgaNgmRI0aKe+zDdYPbh6J+OC0+N07zl3wpT7b0iKynB8lUv15H9N712qxiyH13ny
M304xSGRMFLYS2Dcurg2fV+VZqddu4C9cnnMp6JvmbHjyhiLN7rrwwsNIP6uFYN1xnyiYwlx2El3
+5z2sLte2pLwvrdUuLhMkj5gEMQW2yWuVEnIu6f5dxPM3gAIzV5Kql46OrgHz/5DM60WoApyM+LU
wp9I2F98n13ZhCKyq8xciQKhYy/gVNSHkXk10Tptu53O7Mpunl8DIAJF1efgea9ExM0W7jRX6iCL
WUgvvriRWiGoBcSZD1IcwGw3rjw9SUn3fWyvwTgHoX35PctB4gHEuxgw5xw5pLvPFAGDu0qf2+Fb
Dcjqn3RqRDbFBULWEkzeYi4zNg5bjtDKrvSTpQ9sCPSWdtF//xLtxnsMe5QwpMX42ur7wHHPYuwI
E5WDbIfd44FZftXwy4QA5rW+/NC6WxJ7eYwSCD6if0Um52v6LSzw1hHUqGlyfsP0wCc8fcaXatp2
qawi9sV/71QuOak2i4eCxwXtqiZh6tAzlftXaPREtY3eB+qJWqDZKXOxmb//gMcYup9Kw59Ebthe
DZF8JpgxYCrSthZmhDkFB4GSWngcpeDVg0aqDhffU+haOjdPYV695lTUdQCCryog5pQU12clTRgi
dMxWt6sFX3n4tjigp//2MaSxK4XzmwSMYwLPu0QljcHYQf+SaQHkxfX1bFmP+Ax/9XGlTACx35TP
NDS3qXHCo85yrNgV+VQja2JiuzxF2hzkEen1dIvzZSA6vPkvedjwC0u8yY7kNO6eEs+eGq6oDxrN
ZiJomzKGl4j0y8Kh3ZGI83R8aRrq65URtCLuxySSYynY/y1sgppy+K5Fjc2X8S0+DWkA2TpbY8h6
+duVt3U0r1nQ98w9uYm1wC4m4OI04+0RYp72G9NIXWKIL/golD3a8r3tglrANaZIstMJeObR9wj6
z+kx/WFJMy9DIq55Vh9M4la+aHF/4RbRlYvikympa/Hdz8++fhTPkeKdmK4tfRqAbXcy6R8x+jub
GAh2vcRdTBGzCh72sb8NQPjmGeAZaNdtCAYRse/HDhpMWJPTvK8Nv8RXESlZL7KoZYfdx2oHvvVl
ioaiaxXPTex0g0QHt4dAbYxj41PJZYb0JCoesheDIrL5zW7JzDdjv6Jr6Mp7HDgjoF14KPgdsJGi
yujakdLH10Dn4ekTmnsU/2k4xLWF+hMKdry7Gfs6pv2SRBeF/yc06GuB5N0cTtN/+tUHSiuLkyf8
/62rfvghTDWjrg03PZp3SABME4xvbAInuIa1ydLNABEAby9w8F37Q7pzuE8PJYLa6tL6mk+6drRT
3CF/qci8IviRc22+XmNqbvQh6Xv8vJKRxXUH/p25bAjAwTU1dQQbxq/VHlndZRJeome0A8kWwfvJ
48IofCSfwsVPGxa5z6+4NNgUEXpIZRmMV2MGl5boimm1R99IQL7wPhuyfKOI/76DAtkXgkLqk2UF
aKKyIo/NZ+XbNi7a+Ap9C9iehbWwZSiigrwz3IJUoNCmdGDbKh2pB+pG3clC+BeYTRS29Jiu+oWK
glOk52tjCD/A4KX6g6K9GeVy63Z18oJmxUYThHCykomYW8ZXd5udY3rQTAffKLlKEu8WUtTr8x1w
daJDbbTBmaqnvXR73lFxOJuoU8goLsWkWsUOpGvbfffDraa1rYrNnylTQ6eX+rIKt+doNZhYVk9O
rSQFMpUvo4qyhhQs+8ZdsR5rSCE6ZZl1bPGsSDyPDwlPx0tCTWrohPD2OH5/qBDuFtthTzBbqFxA
7nAF6tdUEy2CX9K5XAhqRGcvm0ANd6iFUNGTbU5bKwPA+iZb3cgf7DhaYK2ojESOOW4/0W0Ci56k
nuXCrUTficFaJzTsBcT3cySZRyj1hD8wSqiC7169zwL4IskbUx1yakO/w2khCexTUBVERJqdK8vp
FXTn26oiCr0IIzbTv1yPH0DhlOAtti3biRHK2Yi4jX3LMHl9tJ09Qyw8u/xP0deFm01vvC5F7a+6
/mYHNX8CII5qKJhihlGwPN7TYJTNoRKxpV4aWaBI+Vqxhzuynx6MQKxOqdK4IYuJ5RPbXfGA24d8
8b5Qs5zo9xDi0davwiNKlYmQznze6LPDd+yY3pQxdJV+XdNB+eIOGLMJiz8wJyD+4wlm34w8xQzK
M6PDy+X55ZTCrMjHX44BJdcOQjno3czWBW4GIFAJlk2GLsNhPKHUB2tfJwEBPt2X9ix7l8QTaSr2
dOGH/51GocfO3FamIcDHlRAk15bAr+9hNrv6Zv76vrL7LPfE7zQ8mDQrG4qi7OffuRYQPocLuPgz
nmc3Qi0RmpaficfvbLwxrE/thf58q+Fcdv7b1AQrqw/C5kkDk/GcTjNgo4ncupAbFbMAJZVplmd0
4Mmw6zncecClpeBLJEMB/vtunNg39GD5tiuBOpCP/TdstPGIsUINT51/e/W6rIgvV8gi+isAx8Ti
wsEBgznWzbfTqqAkmjaUVqDeGUCYqPtDgQFFgOpauwGWXnRjIBt+oJ0n3R1FDbi2+SYLuiV4DcIs
kNBXHvTXP0wN3RaCrceppfZG5vfAojwa6ghk7RH3sZSY6jV3bkUwXeaHAjOycp/eGGby26wQYtsy
KaLh8ZbKY4grKc9v37FIzuxCukLIyWeC5oO42kmRd/iymX+kDamGiiwIWccRJZms+Y+GNpxFE0Ir
jbABSil/vLVeYOWmPKTerL0uWEiX5eTTQWo7yJPmLaSsQwimotPqyDwocawL+JiQ68Q6HcBFtEzZ
yW+M5iEhIj3mGKpwT+sf74Iy93WW8D/VzkpZ9UHTwqW2sfcgT1XJDKX1ihK4cOz4SD+RBnYisA/F
uahO0BFQ+uActUKUfDUf66Fzft3m+K9UnmcJWjAfVmkmLfQf5X2n3OX5260RSwvjQx5rwkN6Kfp7
xkzoNVWTFPyikOmn3bbrjxwWcZOxSAwNsFg6ah6OBpwzBO/DaQ3SMCM+nRdcFQ+lg2a5Xh767/HW
binokVt6JNv8cHbW++xUUX8sz1D2RB6trxGA+5Q3AmoOdEpPEVTc8reVGJhiTPMLJtutvyiLq184
doKrto8l/5g048vZSYACW2N3+vCPkD7zZL2/8CUA71AjnwDXllPwuyWNCnfP2iaqm1ftzOoHuTq3
hh0CdRCHJtAJN9Owg27SYXZnGzMcIA8XZYapytHrdDq2oskN/elcXXXocv2VlF55i98HPQHIdmKV
+AmPWoP7EJ6YHFv14mQTg0JBlHt2kQvacYFjxIzO7jWW9jACn34jjD8GgY6wrd/Y8+yGVVp2qVnz
P3K0jg5or8vzQLaK6NSxr0T3g6NhMEoRIyrzMisjGfrLsC3ZgZ2uC1oF+iNuQq5aDqAlj1xWJlxG
H7Mx1339yJZxVXkzkEnorDXzAgzBARmiXZgL9oB9AZQ6m+xaqJMdRlPd7Jj40CdmOyquk1lptJEu
EfL/VDRblSuSVUBoWb/HT0ksC7Bz+RcPLNPoszvdcBul662438GNIQ/haWRkI+M12bWwRO3Ab5aG
T2OMGTDfHNTFoHx2IIJsjaNDM+PS3ZrcL1qNh+mHo+gGi/zP108XmZLARESL/do8RqJ81K3gnI9n
Y/761HiLQsiCWrK+HC57uv3tMsXBspccapiQz+j4RR3HTvelz2941/pdQr4b0z75UQy4625DKSA5
q3sgODg/EXGKnmOaY+s6M4jLAZE+CM5C3KFXypCkL93n8/Aef7fHczLnMyAJ4180wDmlF4if74Na
rcd5WWwFdEKrwl3ANNe9M/rbc6W/7rPLoCMbRdENJRz+nHZW0KVUEoypYwP8JP70wImvkpk6rR7C
697jrpmGJ9d+vN+8o0ONzBT4EIaxE9bOORjlaXtAwf8LaHVpQi8ikJDYO+5zafTI412fBDP1N8OX
86ynn/k8ock+8oKGG0DSQLZvWUj5SyFqSQ1S/iN5hFB+VIhOSVnpgv6bxhCikzznOsMMz3bVKWd7
tBLcuSqCN8t0b3H7Yhriqs/I0XlRAqrYPjKpndHZfb49yWpfn8xHpDRUFkhb38augOOKL+yiOl4N
v5oxLcKxcaBqNJP+y61w3HdHlJx72jZqjouI5+ENQB+B+yJQWzgB/xkzHfPgYnMBB58IbsCzfilX
YMhEEzIqAdZ024JomNsgkoOPeOmAYxKBxWpEyLBLOS1fiE+btXTGFXTopwIiYlIyk06x74trKGzf
u3zE6lX46NrFRduN23ieMk7QqBrYNd/aILchAufJ5Bq+FWht2BtTA0x1g26LUN5EFVED/Y4ZKznz
wZ/rKxaD24gXdB/bFl1l6xLsG/N8wyOSJGQzIioHfTKopDNdbWMM5N4J3APWHPyHvSiBOXeDd48F
lVGMCs78XHgWDcxZvuqXGUOXA9/5P+SFCYa5thDpi8YjNtPJDYUVV0BzCoYyV8PgGENJtJNrqjhR
hA8trweIvbTJe/4pFq++RipXPRe99ZPN9hZH1rrSKdY8H3KF0kflPkNyqBfQLKtYHmWf6mQepv0N
YDwHbq8w2TXxTWf9wDASOnYak1K9rHHwN8TcRNYYX/+jxRLarYw/gQSWf5dThBRSIYu6ZYqumPMM
7Jf+bONXb+/PTOrjPmk3u7Wjmmptkv31lU+iOfntnt0wXIZO+dwFHEtSehbQ8tR+BweP+ykFnf+W
3Tn7s4fWjjSVRyyhE/3siOkKoP4RuqsjmYi6kriXOSEWjOEJX+E7w8SmPK/PWYnMLB3EYptLgQOf
bSNfRf3dMgvM4M+I52KATtWVwQm8frw4WWQ8TdKTcrBnQRzfKkOBw9KSk2JQ1wIOIL5myL1Ta3Y+
geCSeqidcCGfNV7GfcMb92vL4V4dpt0Q8Ov/XWYh/Wq8cJ3x2+xKrdkZFvD3C/dua93o0XIphDwK
Km4erkUsJin5d8jYiHiJ3z7pla82c7upy0d+yxrqvp4q2JrGEgLIM7HCzqts5YEUfEhcTT2p80uW
gppl47jK1w4uQJ2MqURwvG03YPHSzwHlFQde2E2zLH27OiH7uZbptQJ2elMr3qjonOHENi4sVyIc
/fFUvtSYS9Kmd2hbsKFqnkmOemQzgx85LjWCmoxk7YsplG1R8hX1SGgxF4Isq/0Q4iri4MDRKLA/
sAT4os7cj6aJsZmiuVGZjx7gnLwadqNnBLgliW+JXDfzfYdr6u9uN0We5vkTf7Qvy710byt41+xz
4lF8j9jDpisBK321oQEXrxBdyuhhb6Sb3/KuwklLMX7jymX6PCGgTi5o9WeGTTQdqHtHY67lZEo+
sPYFS80qVTUjtN9KhgEEf+jnMXamW87o/wbyJVNkD48GDkAINhqvGEsdf0QVOqcg1rSizHQ7R+DV
f3bitjJtnCD5aPR74jIm/A8wx68DLVCJHslOI/TGcJ+gU1WAtlRIh3tTE+YIfXVY3rTdS686Arkn
qcvRy3Jl45qPm6F+epZFhjCwX//V6j7QnoZL+E+3cN68iIfmrVuYY/9aXVSpZPzZ2ApgomL3P7Mb
kr4jPRWfCgtNQJ/R881XxTKMbKsKRWekSWmlMbgFfiE/v235lzEiJm5yIHLJyoek4LiK89g/MrdJ
COTTx2kSV7cUPg0vDrHFr6qqQtE/Hvq0ZB59jyh+/EXtYLg24XEyXUSP5oohbSODeYH3RjW9/tWw
nHWbYJFPQLmNV2H8s+fssCfx9IOSkzF4OxCcW2R+Os0mA5n+cWUNa3Z52VbIHxQ1VeyFTechSv4D
veo2OnmBOq9VvdL0KQKCrAiKdjkftsJMvx9B/y5THPIPUUFkwA+dg5RHLz9851wHknsiFpAM5OcC
fuQH+yJMUaW+uJH8hk9Zty6vVpBxEtKT+eFavoe01pnuxA+WTXzVHivjFTVKVmEW8v0juwyzpNsB
5NRYlX3H2NGze5dZZPmV5QLxrwm3MWcpPyPhAo9beR3b6aZJv71TiREa03Rp54vOFNnI4Y795b+y
x3u4KRW5oznfSI1H4eOaSYRodqju61qV7mRi0Cwf+9qF9HIZq9XzrlVrLuuWq52uH2SL3XibRSEh
NYDOxo9q25IHXIPCM4j+Ukd5/6MA4/rjvV8gHIZVXuROoC570Z+evaJDXD0gibrp5AfArgdZF7Hd
RzbsSvSUl0qvpcDlE6Mr+zKXlPeo5zBJ3+S7HYqT4CwlUlyxlZqyYxPtRb4GzxiD2T7XmgQTnYBb
TqHhkJMoOu8xGQYPObO2RN7+PTlpFZgweInyCK1bzPPhRC/JE7RReb6c1bBUE/vPMD0sn59neaVw
C+CnUNlp4s/aPaphe6NOFD7j8IXPUdxH45nET2fcGy4yYjwzuDmS9j8apgfbLyKRJpLGBKL2cwPH
7vQmyf5e08gOJIg8JRJczDgSenGTudXqbu/j3x4SOykODcPgzhR8Z9g6yS8dtdUpBkgZ9KprNSmg
WYebzUKK5OoUqHwj0uidZn8sg7ZPtLtgAtYf46OJM+pm6kszF949EM9/UpQRp7fQrYbJsUk2fWSx
afW9WjCY71RVLBiuEg9zUTQEX7qhInawivsiS04wUrX5qXrtQd7Dem2pwRyuvM3WKEiL62UBZ+pu
mgg3R9Ushj1WEjKLGCYH9CVRH157JuDwRweSL5DPBevWcYH1RrqGIunPndhZp16nXtG+YobTIquf
q7TMIquD472jyAELyMrlj2BCixSA9KyA0chifjcflgx3stEgNP7d7oR/A78aDTgC/XTFTAUf4J1N
vl6VMDGv9rwW9CSxk2s/773b+CYWSLoymQhv7fj//Qbl8X4u7pRVdwdnuLHVSZmXJwG1jwGI69bd
nlVNXZWO+1hGPFomp/KG3803l7yxj3+0QQdDkULHDQWJk1UvttKvPeUXllQCwxfNvokGE1c14RWZ
5RZD3UttZvDvlIAznWtXi9Uj5wsDUxhmlZTl3HWrXXIJxuE6nkSz6GH1jretEH97SVazjAyiUY/Z
311SvWCM1eOXp1pDQIUQgVRZYaDqRopZ7vJ47F8LliHN+7JqIKgGwbPm4jUpIsDBp8lA2FHL7IIV
iq9HZv6IAhB3Ax8bb0vvIRcwnZXE98iGNYRnpmRBEp0JppRXQlZUjUqhHHZ+aGExBSKWhZkPdNAr
NMJ68lfOu/GPvLPdynGPw81q9ggnWDrLUHpqKvAAAEdlOjPoJ0vSdWHFwV+Ivxl5NkClAoqr6bUF
Ms2D2krG6iNK/3XyGorZdjLHqQPZaT4oLMabmGzDMFWNUHIrlt3yFKrTE1U5yQZmzDpaXN2lBHaP
/8fEAH+rxo1oEulWcqT8bV08Ecrg+SqYQv44t/JPgBxbZx3NBmye/draTDuhwbYAs5mcX1QYdIZn
0jMsjVmNuGjQo4BJAxHf+Li3Rn4Uc0Y5PKwmJn05FCFo1w2dOKStEzX0eY9TUcgZ7Owm0nXRXaQ+
tkI1H6GKmpKGBn+Hll+IadGtpCm4x7Wx2Utl8EjgPuacufw9KAO9HbjWMcBT4+m/sErbdVc9HZaW
UX+LO84nPjFix2vsDb/5Gi/uXeuXzxGbIZlkr96McRB+LwiNYkzpX5ByGN71MWOz3tzXECRxelBa
/24D0DnIoF9zp2+kDwsNs+19pO7cULYlVhVVdLV28pooRVRG8htkmKhs6DwWoljTQyzgEJaHRSrd
2hO2zeNlX4jCqpYI+/Km0bFPqMklqghKr1rekksDmafbl67Dpjd9GoiLw5cbh3B5DbjSyp9KTTuV
J/m3Efi/PKoFXsV75Tzqx0jrqJCu+xu4OCsWu94+YbXwdwtvTfVhlkR6od1lfioCqQ6d37EKN8SU
mDmw5QfTnBf/jFyK/HRRGTEfniV0TTjSIcOVSckPTryukNktfvPytj/n1AcoQmRkom7Zneas4za4
hhZOS8TKn7k2oQycEBEJE4MyLMF5vxDfJ3SmMkh206r+69DUlb3a+iO6ffPywHI5U81tEs75/UyI
oYP5+VeCZ3R4Pes08H8bzm1sJ+2nFK1oQiCeC7++dtEL4/Bwq/Kjz20r8vUGDc9HYXgdfAH1aFcK
hPj2/mFAF1Xs5ubqbnhpytDg4i29w4M4O0c/rDb0AKs+kG45LLqElPBpjR6zH0o1nxQou5rHLH8L
Te892LHpBpOgfgp6Eh5KH5WWiDdzk3yzLM/NZtk1zIOzp3Hfgk0QlhX3/AzQerXtsPWxRTL3R94/
yFZoAkyBfQbWMMX5tup+s999sS3NneLtfmocD7LkehR+rRogVWeWPYQr7KTR1MtniLwKzyxUV5zV
ojr9VawRi2OtsPh66cuHrONbmcaD9j+hE/F4tSlCtqeDuuwc8yOGIWpfgFugZ7Rh9lHtkP255slf
tTmrLC6FrDmKiw3gaoaokC8jalxRM+nIV8nIPPTd/ke/GsMRFfiv5jZBnrkMymHR5l6rBlXv/6F6
hGuBPoTNl7ZpE9o8cDqvCYRrSDrwsDuHuPk/1K2WtlHODmUgCzturT0rY4nyMRSPOA1tniNYTjmj
01+swiChsTmNH3nIwke08X6fjIa249RWIz0wGX9HRgnPxRC+O/ERlojVdHjlBpQKAPpT3HizXaSU
hWfIJM1HTBCpwb6fLA5iX37HbzDR+K+Uq3umdif8IN9UZP2rxyFF/C2Yl2jiY0AWyuMnnuRTEANd
AcHtaXtX13vAfNgeaSNwtj6fLEjo6TC5oT67sqgqzVjN0yRhVbl3/bw1o2s5wZJbWQfMYN0Y8yUD
tb5IVw7Du7uNoAWYYFcZGmHdTfv2dcTkqUk4lXPj5VNkXJmKQOgj/2aK51oD3Wg1GWt76qGuSTYA
XHvGCMOqn+YiRn5Hq6wRpZQQgU+zvkQEewOsHPhmyhl5sSyk7YAUwoUleXPkfQW9oeuyYihC45O3
2A/T6apjppuNT4b/qojxDYyhqQIjpgytxn3SAQFY9ErbScJYSXdf5c5BQEi/91cIkNIBPJUgDslY
o0mKT5YlnYoBk591opb9sgYcoWjsp+q2AWOLEgiJjlRiBSvuZVSOlqYkCoNJH+wcjoeRCU8t2Zez
/iaEFnWa7Rt0hysh0m8m1GWIg6I/dYYWlCY188D5bTs4kh45/XABv/yaz3LE2w0D2Brc2piKbv2e
E3M0UV0+3ei8jwPE9I/bc/Et9JXipBors+zEE/97dRor0I0CjWNVuOcA9WNfODHSjs5jL3FOByez
GMF4mTI6jqE6UZXEXB7s64N//X7opW+1J05gna2OSf1ydmS+CcNkqKNye+iu7UcHUEyXlPrVpA7y
huWIlP3n2nG6KrmY0nleZdSszWn7DklPJjwZzYpAu3drqs6nvjR9u+BdL/93KLet/l5K9F1+wqy/
VORyAh44bdowpF+h4PuJ3rzEIDKsPxW5oduyqSwlZoR7kuyWfb95GudXiCuePmycqlQad5IuaXid
w11kVTaeIT4DtbYvQ4qcOVMzwtXhUlHwcZpGPGn0e2h861VY1gsvwAtcnYbJhT3JLKPHx8ybxvIB
+FpsHEd8Fw+NwEo2yIymHlc0AkQesV4KvRJVd8cMMgrxV10pUzDsB57ZV6ZTJXf4iPaL2jRp43Fo
vWpijXHqdDIbhDK16iR6RDV9aIlTEVz2YVPCZyiMPgX2Rhgnc7E5q1+6geVbJGCop68laUgwHatP
QyPEEv9dqx34vVZNYlumnBMh2QzAAxUiyzc4UMlgvlJVKKY7ai0n/hfMCiGEzSLhRa8AvOJcs5Ej
LXPk0GgnVD7ix/bce6OPl7ewb0nsAub9mfH4TxhP/Al1Sb8TGV5gzmwtOgoRvGcB9dW9BjthzWDY
ZVgwfER5+ihUVN5lxihyjH+HXPY70yJk1vLwXj8wGW3Xg66s1z++Skb4oCPkzOQOiqxjylAfEx0I
so25bNA52EVKkXEaPior2VeuWG8Oajy+lpAGRhB9tghXYjy3m5UmAjnZkQReGOlKFeJle4X0DeyU
sj3Riuw/5ETTUoEcDAoTZOLSTTeEc8VRLdoUk7tvvHyFs7/msobatAcrmmjOSIEe5x+j5XMU/Pll
WjL9jo3hHnUlZ6lhq88Xi4daDYzMJ6HBc4+H7C7gMtXX2lt3jfcbcpFXzgH3FwwLACnYVdlrw9vO
bc0z4Lqff1qZt7RbuGPW6Vd9c/3nNF2b24EOPd7D/6u2NhP0uPWoPRlsvbgxvBBE5+Iyre8Em7VN
6ccpz3gotErFmN/v4PpkZDTWgb0IphVkvVk=
`protect end_protected

