

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
b5iEwcuh/jbBlgyw+948d3lvWBbFsOTNVYtA4pJb/+7lAHor6DKhd4akfRWg+MPGWaTgwtrV3Hjr
bBdLdBNTBw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VtyA/tLK0cCJJRwkcmojHVnJYFSH/hY10K0O1xHrVFcESK6dXqpZL9jghTqU0K8Rgfgyj2mbpSmS
d3OjaMJOT/0rjwEIwUBTQhpYCQbUdyb5e+tsu6Jle32rY2EO1nN6daySTSkOW0tup2zZBsIOCr3t
+ejm/NK+miEBBu1xCLg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sf+0xczGTqZZx6dcqp2GTylMp6ojNl/Es91rC3p2Qk7Z8FK5U8FSMHtByvmeihj5pitp5aOxAIcO
cjVP1mZpqkA9QTc6UkTBmHGnHSpwqkUrzOtsT2ws44zFj3ryr3hssigeWwtnVK13YgLrM+5chsUj
26gA0jBZIt1YnLsbFPdAg3CFuuIkHWQ39NEQDeG2BTbW5KtUVyDTnpctdLn+1GQ9lYJeC7lVtfwI
4B4xEL5dhZYik7uaLaobO+7jlipeHv29o8EQsg6BnOj1c1kxrXtTLsKozU5mRUSyPYYAw5cgAAvI
P9ELz58Fq2bFhjjPjC0ULrxEE7cl3R3lE+lEcg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qzj1t+dWRPGHMv8nVaAMZRu2BQPWmF3UL/i0LvBgsHGjHy3fNoKTLAs04wnbPCVtn8n3ytCSqZ9j
YDEGkJeQd/ctkBALil+9bfKGzVPGZiyWs36ilhf0nuaehXbM+Zt3Nfkh/wd1LKqVrJhOB/A/iGYL
jRkozXf4ccRU53dhQZE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eo3jj49OyneaHUaTvAS2/lR4/3L9GHwLzRAoxweYog0SBxlqFd2rrO0OlKoc3GfXgogda87o4tmz
l/UHxih0uJyK1snlhQ6A1EHKpMBpfD++gCN+S5IJFV1QgpWejKXt+0a0zp/A429l2cS7KMD2pUZc
B0C4VRE2SAMGJhfx1GIRczPJREH6ZIkDU1qmMs04rSp0PaGn6eV7+euaxeQcoqowg8QlRFnxfvHh
5JrqhxNCP2z579eEXYXH3AWOzWM/EnKEFUTbEaxMGP4W7RzgRCZvuM41apmXDWTVjEj3gQq6xKn9
0OWO8TXN0ID1dcJmFJe2x6yA91duGkuqWQQaEA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43760)
`protect data_block
VBogWMQHjc4eMkge6C+BCOg0YuNRDgRarwx+E9YArYppP7TN40NulVKmGkmynUvR/M0tkCYF9Kb8
oIwjDg9PudPJ3P6fI7gOXn9Q/2gOCGschbC6R/ZcVKk7fm2FCnHz6/XyAMGYQUx01acnLecMBIxX
OyErF5UEFjoSB65YeDWlcZYr3ynwdo+YMexvP7iPxNm9oIuslppazkULxGMm4mWyfbMP4n8GNdy0
8HrY0N3pn5ea0jjWuLU2uZ0ZZEbLrBguHiCudLN3oQNTJDGs232k3l1cCYEIMU7nFYlZVl8HCPhe
1VNZEg+1I/uZV2rTlIiKNEsnkLTk2XqF5pB1a+2kpJ0Q3y113rQihfvpub0JtmEotTlIM1M/rWhF
IrmGRgQ8R0lf9ou4lA5HuwLbgINluF4IVac6/UbZXose8T+gyqj/DAWgYC49qJqpryESf0OWZRvt
TbuYZVaxEDWu7WC+//Dk1suqlADCRuishKeYJp8c5PKdfFQtQ4y/V6tzO1R0Z8B0w+95db4RsPoN
8KaQNr67NFg3DHaEhqBBmwUoSc42Y4vDLkPeWouOnUmMiHnEUunXAxO2TsVpAX76T/V1zYoNHnaw
GCckq6v1QIKyh7s1xViBSzDq909RvZ8IQSsVkRoi3wr++9PmCmTP335bO+vYUfnytKmKkeX/wsPR
IcbMKI//GxOMah+RKJV9UtOBf59hsTJsO86cMkHE6b1vqEwas+9ig1iufjoij0y0qvqSmLLTDDnw
I8hh9fwK4s+6WlswPF6c9LWrHDn9dWpcwz2snK0kjdcYyLzLOcBl5U2rhbAZE4HTYHR+MJXnsdIx
gxcKxbavZZizLxpJrZtqpOYqVGtzMlSYXn4TXJSLK7w5Nv2Blq5nu+fi0k0hQdRNjTcq1TPRfZJ1
/b7QndfAwKO6ft0Np6/whX3YfynIY6tW3p5XG64xMqRxLfrwQLjarEyofvJynIBKti/VEWe9bPqu
MgdZtYMOUzAvtHjKJaYGgiWvyaEKTcMbbRMKutcd2YKODPrA0uzF21K+HvhWBNbo7BC9ukE2yBFP
xDVpTnKtbrEo+4T5D7eC28ajCc76prbTxXLFaiouI5CMbZgUussdvx7wapwsEwdQnsBamXTYE8rP
vXRWTTwTgRIecQt5liIZs00AoT15HMPqz1fVYyOB6UwQE51Sp9hdX67zRp8qSsUFb2aqdHwbC+/w
uJYTqc53blkdEWW9t/b/yZxI9dFNrlEmRet12xx4h0687qmAUDNih78j6fbzZOrxG5wFZu/viR7V
0M++7NV9l3enh/o2c9oodjgc7m9U37r073jf00/CZ9pHLBT38kylGxRVUoqukfsAH/ltGuxyTL/l
dTjWLq0oxdMTMgGONkoE7YCGcXkdZieaAWDklUuuvTrBFiJHuoAHBN3e0rnzPFz5NDSWtsGkohag
ORA6nMSLB6wEfNl/eoET087pLG04ysEtqW5xLl4dav9ERp37/OmS+j3gQsBp213JqNECntbw2WYo
8L8NnVYfwX3VsENqVvkreyIrnb60OmxnfhUJGcIFsh9vymBq8z0svRDH9Wd+Mj+ojKch67ldo0j8
BgphmNy+XsEfbxr1/hR6ZpPiM0/irEjIZcuqU5qETNGb4ES+P3Cj0EpLDdtNmUQRdzsOw6oI4UMO
ZC8ErxjgBC87Icru0lXt8VTkflrsV2dPGF7RuP8s8adrGDzamGc1wV1YEgqdRbxFEyJB930q34E1
GE0WxhCCqsv8ef5TegHp5+TmoryWT0k4aSApGaWZ4uxIlIz/AUmuSFrFxQdSCO7dqOHSRGT1FGqc
W/KB0zxSlVWQAGWzNV/6dOEZ8OqumMp3UhC9vwOzDqOZ0HIcAyBKVsabRXckyWAc+aPN4s0SKT4o
nhPE44c9oZxFZrmmMk0vR5Udc8PcbficlFm2wv1TpkO/aD3MkAlPmovYpFzvJYzEGbttwWqnqhlZ
EsU8IvM7R85xt0nyARNozLfNqjv8f3Pm77yuDxlTtw4qdmsYXIMlVkDUb9Gj9pY1aw/DLsNmMIGE
/tPAvw/wEHMQC5oT1o/17CquAQpDt3dtAsA0TAklEgWXMyof0iIQz9nkBgPcqok58LzQCAlX3fXJ
oEpcg0bUg6REOchQJD9NEcqr8w428mVgH0xOUOqOWg/oDPpIFi1fV9ZzVGQfhB2VydJArobzxtB6
vMPnAiXNUBm7D//W0WctNBZUGUQSzIBIfxk8uuUMGGRYZDRkNpKP1ZukLQ3iDjtvCuGa3Tci/ORh
ygdkIDXO7XcLaQb8TojFRXoUDRkGWfwQJKNSSiX5/YEc0C0cY9XABAx+CcAawrylT47lq+1DonW2
oMJzKYRWosev324FQpug6T7yjKoSQbRDOzH5szacEHtqPTJZGbqO402PDYYEn0bmBjuLtaSMW7mW
QQfzX5oTl4c65NxhIx54Lxc8gonkrRwintajbAUQ7ImBOkMGxPkK0mGtYAglwlVUpY8wDMorsgVP
3JvyfO+u4gGCu0qFX5ppZ+4NBo6uQW2Ld6Asg0uiVY6wqDrZV2x3NqYmPdhQiAvUjLakYvQ7pxCH
CnY07wfkTz21NsJep0HHPA1rUxTYLJkaoB5VdYiUIOJWmVQUe15JgoGdcqw6UDd7yMY/blNHioc/
LsUGH9Ww83e+uU7N8SI3bGRwthH/0ThCNLYtOkOJy12SsJWoTO+BAmuJmUrQCTIcLOWBiTnS24X2
eq9HiDOuXb7gUl4HS+fg7kx1lTcHYUItEh3oxuQ+MwBHH9SAT+t13+LSQ4hWs4G75SCM4PgbNaFp
Abm7ATpFS5DAGTG3bHznJVTY5CjqJjhLQ8iiSGMlXtMhNozgo3s2oEYUGdVqDhX7Yhmefg8qmoAN
EYYR1eFBlwcR+EGLqHW3CFlmB2BVnBlZBCWXlrhU9le8Iw8ISueMly5xH06poh00t3QnSlpVUYXI
Dng/1TUKWB2OWO6TrogTb9wE0dJJCrb/iKxRl1SFi44ngA/5wStV7kI1nz4XsafrGbq8oBN9L2cz
XHnTIh8MuX+cW8oSMqpwXArp2Xwl+Pk2MKWSc3qh/6oWrOP20aWXJwmt6fosFdkn90A5tsR1VdLW
1DT6IxttjtPooJ5V6AWw47kKRzfHAWrlGPq8kU6NOMpkK9J6mvU1kbJEIrBsaDe5/wIs6onXyECQ
gjq+WBYTUMduapFepetMtT6ng+GxogOya3vQQ5i8Nf0qxiDx41K2u6LartGUbhtGW7Gcz8UGZrWu
8VffEKPSsAbUzLZ6OzGOqjxo0V8dY7bLtI7hqj5QzuTYAzBNwD8809/M1GtCrXxv2XC6ZbSzq6bA
6kqg2jsycdUS8Dup9IZ1fZR0syQ6JgJS0HpTGj5IEhAE3ZPZXseiEd0v4HsAApCLiTWrGqlOLEtj
cZXBOjNclsPEPWg8Gl9LDWCOnhTUT/ds4gj9aty7V7iC2ZGo6yv91sT73rF1M9wBlCjsNDrukbDx
CF8LllBgmaG81T8pkW4GL+MjWYOLh/6JJtUbUjjExVFLb2f9s622xagGCCiCaFS2yD+fqI5AiQMc
tVi7HHrC2QUw79AH8sas7lFYlVY9kx3yYsxEwbim4L6TtAwAqONMDXKOIsx0h+5kzexSnyI2qEvg
LiTBiuodk6pfiMtAKILRJKoSl8vUYwmMPNFtvRh1Pl6Flfg5NciPKmNfcj913SGaaGg/wKa80/6M
y9Y9IVWqJT+/3NieU9jw1rIM/dREdC2fQghcfMihq+TAtCQQrTsaVgkucJBDIfcmHkJJNIVTsyd0
zrQQCRs4FaDP6rQd1XOY2q7mIo9QtrQ1MpwJwuXgkMtzSPKas13T9XogtVZ9NiX56LpO0yssUKdi
+pljXQry212UCpChVXOnol63HRXBsvYOKiYg6g8xoIdf52OHqZ1jD0cmJ0wWr6/kiqfbrmM+hE1+
h9pB56NIFdvXog3Q7c9qKlPVSMzSQV5jZT0RpzQukPZw6ARTDMHqg6KNjojle9YSer/Wt7on+e37
lnltNo0i4NZqvQpazXtJB3pxO9FDkOTp1OOHsCxjjFlTwHmIi/s3klWkBcIiMMXgSfdI/kGgVfMI
CJgWMqt0N6ZtTrmL/+DjqN7ALtNYXxjYHH9UhWYehnuRWyvhDiKgUoMMrMC/7fvHdzLzzMfi50qO
MG6HTm28TN1tRKLW7RmVkdaa5WDFqsATvFk9B20CZg+0d1od8QJ2VwoCQkqWvzgMTZZri89fqLuy
nPFJ9hWBaBQHdf1kOgYqcdthg4oB9ALa8NQjF+5jm8MLUrik5U5U0Nlv6/OPQpvE/ljxwWLruzR6
f6fDVotCetvmr7xner6StSaie35Zdc3bgdRb4Xc2Ux7q9i4SynWAhtGfzGTaYVyo+iE5H9VzmtV2
EZrNIenv7M76ebyaeqnv/lrj9WXP7D4hERW9jvu6kqVamYXf/6OvJgkeqkdqXngylrId/yg0qvN3
LxqLfO/yU7uPpMAdj+lG7eRJZvpZAqv9NKPFN+gtWx4a0/u1uUrLMBpgtzF12XcZdfz02hheI6Jb
Msw78aTPPKUjo25pQzHWdHYg3euQKA30bIVw1i3OmDg4EyqRBW/Ni6UvBI6T0majRyel0EzbDjU4
Pp/rbCDg9oLykmTzGPLXq4PTKTieHXUeFMc5xBMH4wv+avKQL/R+Aiz3SMhG1u+PHIWz2ivwBR+q
At8aWUSIaLsY3g5bhEA2BTAPwLA0+ecNjumx2RreiWL/SKjpF1mEcsng/MfA3QWGAugbcuPljrJz
P/oLQn/5Px3GzUSkXlnWWYOFE/MT7vzMOOTqTrmIVVZeV8+SA7P+UuAuq8oHtMo51xSa+Isikilq
u/8UKf+mLKV4jdRXNbxUaNhYhtMci0Oz0lKaAO0ijP9CxXGN6GYzYD66W+qkwflqgOsr5Q6TMNcO
Y4l2+6yQiFDlIX98ZQb6DJYxm9eJ0ZEBEWGuPDDB2cYOdDNvaelEvMLWTmOKc9IgiOIDd11x3nap
KKJo2ADurDSUZsxIX6zq13vmOoB+1XZ7lS1gew+EjNz/f/o6h/le7pLDXj5EGYyukCKsqS0H+UJB
iA+aOLC1+PgDxYNVv424h/g84w8cob+TvMqEfnnYO5+o4jjzHD5tTiomE2EDtzltPk3bH3bQf6R2
+T0JkydBGHnlqrjP47FIoeHZyW+RBUxJHXc6LR3koAzVTUXdBs0+L16URBB0A6HeRxA50DvR+4m0
mD/FTk7vJRRmP9JZI2Qe+uJlVIrRTTiyfMvDy11UXFz256z7Ss+gUm9mpb6UnDhTREXo+uUBXak9
dIoEc4g3IzZ1P6OxpT347OtF/Vin7U/QtvYJggKOTkAyABT0W3Y3ZAgjLubZB0R3DEOD0esrhPzH
VJ5k5zcLbKjX4zkD5A4g/R3YjOpGp4vSGAnEQ5D9RVg9MLK78kNJWrQ62e0BKpa8paNooOTMcCHW
yW5ubMi1gGHpgA1FE8T8dODtxPNbCV7PoVWIa5m/rCCRF6jLl8TcgXdE4gmHiF1tAYlO/WJ1NZZD
ZWHXdeTYNdDBbcpcZwyohTHZBzYedp1gU55QR6d7vh68pEUdkA60NdPZ/MD4tkqYYLbvMBz3CXQi
0/PLZrFnHnMSzDkHXr3wLU2T39S1Lq8xUXWGpgjSyOlkgWYEWG/+RwG2sZ7OD9dAOSoSPhafsmef
YM62Z5LtbFjp/wuV19z1Ro+vNwcn57roMRMnY8wrtq6aQbFKSD9IrJReYanf9kh2D4ktsgISeai7
KBXiXF/yYSREljOq90PqCuDyp4p8JFmnHL3LbUBgjquO/vLcDyFrhEU8HbhoHvS1BYxBzJRhbHPL
bs8D0FAo/dA+FwV8QxDea+EKXKS/eqSEOLQN2XsM7eUxK7Os9Mc/MQAQa5LZfb8Ynx6fEIS7UFYB
FgxgePXG2aniJypZWwTvGVcwDKJfqX5k/p++3tmFv5rKsHUBSyRv5eqZMGUnX7u4ydHnpsBRxUE9
gy5oQ0Sf4B/0vIPEv9b7GvJ+/PrKyIgSVAZ7a+L1JwiVStXy632dt7LJ5PiSDawTX6Ng1CFVqIHs
9p28iG195F7upFyBSiRY94oNDT3j3v4hnUWtYlbHNv2wEEJ3a4hz2QGQz88yYwE+sIutx/t89gSR
RpiqsWO7Mo8ViDR7M8GrpnTkGKIo4kTm181Qqn3wDRegvOLRnWtTizaDnwGNvyeRoK7n9rJMaDtM
fBtqlsFH3slivXVA7ah9IOX14N9+DM/Zh3sbC6Dc9Kn5Y2vmyEz1xJYsgITDzTp2W7hV8lx4Mkin
gLuBvgvJCLXWk5xaQRXIZQNIFpFPU2/6D/TEhqaxZ7nmbrmbt8IuYwBTCI7FxFKXuQ8iVRueQftK
GqF+sON0sqHzMEOY3Y4k5pU6Ik55chkQ/arYrK9UtRg6F+99tgDzFSVa/dzeK2oAo+V43kphY5/Z
JhcZOqqDkFv5hSba+7xVHJmgKSjwsrZY7n8yepyx4sQonecMQYssl/O2VtaF+SAJ8ryFLMAvA2aH
tdGiD6MPgt4n72xRHjE7CXPSUUkuCI0D4lPWHSdP0vElx4Rjs1tAGS5k1lUimLzJjp9V5v/7Gcm2
3blGw6yiyazCmtIVmn3EpXrcmMZE/wfQS3zMV0YKwxuiASqBGMZC9tzHttWQcJ+kxSbY3pbPDsfY
veTKSEMNPOzn6hj1eWblT1tW8YhE/44ABKQ+gphCzV/d55uhNCCoKH9YXD9iOPbNOlOB8xmF34i6
AJU+sjok2bqJztch1YYJ66h4VpY8nvsc7O+mY7gW74Htn5YJOnte0sAncVPkJ2xqFC9qa0OXWV65
DDssqkaN94t0AQ9MRww+8ZiXmtiVPlhFtw7RAGnfMPhwitR2dzNBLxNyjf+xZVpWJJanQb9BOdFw
Gk+eKKqrE6ZlLBDCbjGS5IYCRzD514ZT8EZ2ax7IX93z2S60ODLCANBpKaq0Gg2EtvkUoJon+GDI
UQNa59DlTBaCnaQER+srg+TDA3+HgtMCgRkjS8LKDlDpoDAsULWG4GiWlDIxS5OkRPJ1pUBnEKJg
UNfyx6RLlZTjVlarH7gM/R8IcsOBNHpGF2SYHVsiMR9fpDGweClOaKVTUI++NRMT0NW2FTVX7Ggq
305Fo1Vcnh/v7U+H5urtfws83B8bzVnCWFjn12d1mI8QfuC0dDfLiH3OJB92a5jnAiej4iVwr79w
+7aZUh0pt3RmsX8zKmwXBG56WfhLPiOeVNYqOAcvNzKGaaDtRgqf3V1XAe9Y5OEXCmzVBiUrei2w
udmqaDzt/v8Grdv8B0hpqYminWV9HVlC5pwMe7NGUr65tnx1RRr7MJs1eB/XuywjpfvMe1VI8GYQ
F9+QsZtO9xKXa7/aQ0eH2k3wgg4ZkRsJN54NtBwZTN/15aRhYBZhLoTgnHLvUx77SjsF9GWT+WOa
+afeAh4qMxbD8dUkztrkBUt8YOwBbD57/I1t+qqcWYoQXMEmZ4l6aqH37ZT4PS1ajBLqZ4vLmhig
mGWQ8H5sMZchDS7MvQ5Kq8qaBEIWfo0wg2n1xRkusKkl+c2C3gSr9cTxYKcbXUUMJyvX1yzLl12M
bJz1rQI2Y4H0QBuhy/TmytOW5VXVjEBVEZejUOfJUiqDKsEPxtlA8zMn07+LDjcW5GcZFeaNyKcg
PmWA/WKrKB4qzvFagmY/lOi2tww9ldkgNT4Xgn9uMGvor5TxncKBrEbnz5Z5mm/gqtgEUXueeJPR
qwQLpBP2srW8XVO/BiI2xDNhtFIBoQe2YKWqG11cfyji6x9sFleK45SUgSadnkU5SbnJRcObtN/L
VdZWuIzc5ExW4w8ScNIvPLHmzF8tRk6fgzzdUhHowiuI4gXm/TmXCKcOSph5/3kVxrcLnEI08uH7
YF2DQtKZeNMESbTvgVZb4vTwYQQkxBpa67p54vNeYqtToWxDY2MyYWD/GkdU9oljyA/m6n9X6wzQ
dotVeDEiab+6NSh1gpnx/4qWQSny4osyvQ/Y0hu2jGfgzJQUCEOJzQ65vugxaVks+p9qYFT2HyGc
+BsiRQ+VwEYIK+uIyayBxS3yl49cvghGfR5ES4CrODokptaw8oEufYLhTwOIhV7KnXLifKPpCdby
IMwuYct8BVjFB1IkPkFJ4Sx1TP5gkvgtJsrnm5SQ+p1FLilts3PRzzPKxrKSge9u1jRncoMPafKj
AoM/sPhL93tAAFhHPjo3r7pvmXghDp+TjqJ0O0mVnQ0jvXNEA1n0xwU+7HP6WKiNcqROd7UCNRRR
u1aaqp01FP4W0agFoIqc0p8Eq5BlG0iXAWrUhMqwX9wGIjLr7d5/sE6rD6tds0bkxQ7Cn7zSrJAO
p1eLCmKo8S2pe0GLposuGjWJEsdbocPaKDcDa/5m+vSZk2CIW1u60FTX86FJNHWsW5o1m+fYD5B2
zRm8rjJK2/2ICXlejViipPrZLWVu2Nva9xiK+bgNNZK1z8A4tUBlco4PpP50oj77vWf22nBEZE9R
YKS5vah+SS36/NqLB/kbbHD7j1J9IN1xZupgArVOkeuKN8f1qx4J0I2QJtmGytrhNZTSBc7pwgQf
zQXt2ePfk1LxaOk14RcDB1ifhjNJeCtL/PoCJsbA24uWBkVovcZpZhNzWWQCyTbAFv2ts1ArqE0G
brSUMWK7QVc7rTdafkB2tLu5tH0JL3guhtL3GyEMrLKO6oc0VoeKtY57td9Eint2uTSWXbu4V2o/
9pfibMMIo840GviGZveOEIBM5V31Tgcrm4IZdhRM7Ba0GuyMU5RkvuuvQ4Slmi1aGF17ncwtH059
Y83O2pf2MCuRV3rWxGSbCp4Bq6vFScpR6wuBqQpsoVNJ165MyYE4tFJEDMFTi+aLES0aGLti/50/
8e69G6gMmJZMBXtAmlpEyxXcOLCwCgqwbX129IkftWJdEtiiEceLRAhJ5+AO1Chl0HdqnAie22KP
D+yuVxJ4zE3mLwy0L48rJNLroY/qPgAdUfFz19U9A3zfCCo9FJGsVBAbkhNs+b9rxoxacdB1xEV8
SWVBzxD9WlWls8na65URZNxiPshM5fWG+b3u6AEtOVaLrMxJ7cxWoJTqb1zmL3XtvTyH5RTXPi20
AGX469nPa0TtPRHDlkgyUeiihVCyvEI3gpp7UH5p4cBM2TQMgFBN592YtF4TRNnOZIPIKbR8fKb8
dYdLtU+9hQhof3A6Du2OCCccLXD9rT0KCwFpqxmomexSySZck6yeaHMHDm8k+qn5RtJpoIH7SfDX
aGWTj3JXiOEJ+XjVnj8KPRBUmTlNQDxTq/lkpLSrU9HKtxFO/N2S0nyLWFg6RNCTlEPBlYXe7U+i
Qk0pEeLKgATkx6O12acxtNpehStl4XwZHZgAwMsxziK5V6gdyJGvbOqDT/rIqEgua7v1IH6HudA7
+VtUB9s1YF4RYJPnw4jUlxneaHsxUP2y3l0rpR6t1Sa9mNqgPcNkawRrN/IQZwBqAKzv/NZc0sQK
3Fll4SJte2D/VQVnf0uTzMSSWT69yPe3ptpBdRWD4btLlUaK0J1FMgJddLKY415YWEXxDgLHf+Pg
BYCacbHXc83fhXn1chHmalVue84GMA2TJcQu9NgUAjOUPFCAqDd/ZJl5Eb6N82AnwkSANWKZwjTd
u575MeGVaLImUD6m/UHypBoiOM6nTOTez4CWYui61k6z3KEDtGfrB27xttpXL74EDaTl8Qgujt37
dqgUl4KKmbxvCXhGkKkOqidKUD3dGuS5DJEQJGHta4jF5+H9Faasakwt9rDFjPqWBPLW0E6u83rR
Gx5h+CeoakRH6tVyHpR9WCrOLSkJebsaokgqiNVUIWuhs9fSwbKnbscLiZ1aKKWd9xyvyIjtp6Bt
isGVa53PMCuiNB6ucVfbxQywkRpuV9OTJD5ONZMFUcLuZBfJWVe77mRTkeJtPwde8RIWNC1hRoW6
ovITgFPvC7QofD0iN0+m5Ao1yuD7v/jWgECuwTNT7bQDZSBfCnZUQdwSEaJPaKS0klOb9e0Ugru9
Ne60OwEPiwJYt6BX2fjb03MxRvr3istyRxN4/Lyn29/oY8ooqUJ8qerve/92NfEqfJ88Vpsx+vM1
ZsVaJpOdH/mVlp2/iQ8pqJBxqpWG3v42TnOyIMqGfXMNwgoeMUTzxdwb/wnCHTRoYL3PnNjDlg4M
Uq20LnxUCpZ0n+W8nectja9CVFllihFgxbqAuw5PetJOAZGtLbhP1KC1FcquwTcoSmPvzeypxjpe
yZtI5wch/HOytTDeVTOMfRGNf8VYJDAHdgMfajO8lxYAN3A3V9Wjhz3ENfFzRR5Df8hO3mBtjPqq
j0e+chN6U7DQAmX/qnNu8A5/Kgao6EKX43E2qWI0mOpRfLwGmjvpXn5uQUx2v3z+ym57qVLD9f2l
Bl8fy52x+haaEFEcWMhaxuIWSK+0BzzXp/dPIqyv7RV4fcvmpmDxXGeMIa47YK5Tj+TQhJvCc5lK
EfN6TkL1v6GnuBuuCUSYncg2jzcXxld2sh5D7D7aZ5Z0Lil3008/TuiFXS1okgf8Ih7MQ3u4bFbv
dJLkF9CWKVhre+vWjiC2Vyd5YI77oEvNBYW+IFvSKZiCfda9Cyf+ON0245u4Hq0n4dt//KclSY61
bixKGIuk6Uh0U/xYXLASfTqhv1g7HDnMbcBwUjQtffaKwVvqRfwbVpvXOTPwlA4/tO79hNbfGOFM
CMGyA/kOiFjfC1XPl6Ee7eq2BFFjOZNFrhleXq0sm74corb2/p6VZZi9ZEjjjShaOXVD13pZnVXG
duh4vmZ/oTNwawpmOa688qf8DCDQKx+kk/6NN3SNgEncEnSEMHe6SmRopiiJO004CtfAj10rBDuL
4anwutmQW+6i1pHwiFLbTuvxYUQCPaEKxFBc9Py+SOeq03AMQH5UtvJesNdqPGM05+g7gHNuhNWY
WZk7c6xBxWhKYBhfP+VAzyxCtM+zgTuW8g4J3ZubKN+OmYa73k76155SVp+Oi1zKvNAqhp3+Msn/
9FmxIqHfUZMxEKujiLADa6R+RCo8jfWadQ8zL/TvJG+5lcllcPRT0JDcT+WXcoj518saCLy/YI2m
dwZVVAULVRHilfnU0wlP1BM3cQDCClb1UvciWZOzQZ5x7XB4nVKZUweZcvgTpBs3SJ1wf7eHpNxA
Iirj22hzrEhRpjyxcAijzxmABsp9sMKh7NSkukrZ1y3VThQO/Ce3ZosoK0Sbk9LLmHgN1l6m5GeY
0JA+Mq+ygKMuUjTm+4/RDXiFAPn4edkRxAx4F1J4RmhieiKySd5qrTn0LrCFcUChvBYTHnOnk/wr
92fbEIMOIjlKLWT8LsyJncurYkfUtCqZj4TcLon0hmgaUXEFrGMiAPulRknD9iN+tyGa9ka/HcyX
6d2cpPO2/vzI4Dvj5fIkT70N44CaKvGwrtQC0SZVPrjK8W8PtQxWfOxqyDFyYNcIjdL3IOgkqUCI
kpa67VusSZea7MIteRIsmwq2nVj4fl9ag4bpE2lEO0doz1f3f4+V4Kww4yrtJsOlQB8qUnuV40o/
NPXHXIihWjszpY/AnX0ZdBrh8JBxdScY2EyH3yGkWuoyYUJuHTkZshc+hRgqT7oU+wWPjVW0K9ml
SQQPnfcaLMgkhWF8uKl0yvTQTifEAIzUSwERVRo76W0zn3edKPF+syVxWd7pngMDCAOpM1I2lXhi
U7sfzfYabAIRn4FDXR7GudnHDW2HByHjDXmzKkp1snqCXZ4iQzv4ScccwOcqiJr/QR7LnNFrZ4QC
U+YnthXJzH2x92pq3HAind9APiaJxCDGBBLU0Pzmqj7CTV0Jb3knjndqZjKKh9/JdI4DEOF8YRwe
R8eNUHs8PinVVuPD4p4DW9OWHMdLbtalDOhvDJE2yRHGgDjOLs5Z56m+nZw2ghPvZGEbc8D0ILOn
uEmqI6DjbnZu2eMrY28GfNMFqm4v2fVYS/NBZr4yLhaloIJCTvrsYTbEm+1Yh0S6kdztVDoAb10s
vpDdqxMnjViT7DH7QGn5DgY+BAUloYQgbck3CmBHkB6wuQ8ultCJExxJj+clspSAIYjN19m8rOx3
Wyimh2xo3m+M6gq1XezHm0YFSVIcvFUO4IwlvXnGT9JxOsX+/LAvlZykWDmrbpgsA2ZJoO5jlPzF
ruiSEg7JasADu7t9OHHBGvaMxsw3sS2wTSwNgk3DOc13CdswbVns04pcwPU+cOrSszKwnpaG6nu3
zURoX0ejupGQshAGlvMaOt0StNNCCRyfM4UImjXgZi+gs5VsFujEXfgqjqXyX73yUYDt13Kh8Y5m
hk/XFJdK1kmBD52+DVWynYwrz4uDD0E4Ps0BysR9VBdKR/rYNJiOmEYWr+uSUAiZ6lrX3zUJK+AX
Qls953JhUX3fWDOpY8umknAel9f7Zf05e5vzpoMq9IyHlpDNqqgOarMNnfW/bh4xBJOsHLox4Vv+
Ox2Y0iZgdem2VlxjdECuZOsj6qKZ7Zc9qTr0UW4Z9UZnrxsCVDX6N4LJzWWHTqte9Z2EGCmV/onh
Ma6kmXefL5ux9+dJOTDRcG1HRbH1Gug4nZdm6eOqG3wLWB7s3MJhita5NAhRUeBWtdxSCpIMgUaU
GLElgQ//IFNhBiuQ7nNbaQ8x6mNeu2BScAhcobBVjl0ImyItTAaFlQ+rkJVP27//w5VSS7zGIR3Z
SxvKp5FPvN7kMNf3XmD3lKrmZ0ISivapf3S3s+ZXIgWQNYLAuUpKF9zvspThHTwvaAUUbUmNUC2l
s7cOt0ycdCVijopP1gjGwivU6HsZIwGd5JMt9qo6Wm7jtchenN6Qu3KwS/c0QbS9lJ+0kwWi/80e
HpGFRZXci+aMn1wmvlV4qRM3ecWH4jOOcVJNeh7irz/udtYDXsVqG3j63goAo5Hkr8uNIRk6uP1A
c+3UJzNJUTQZm8Fq3682XZl5EVqGVNZxCsmTk89uGmevpkZE5cxiorPH1EMIFuqIo36MkNWhzw8y
FLpNIObLKyfXDshYlhTBrD0WIu7HS7EYXvNcIXqeUsvKxJTRPHHdr1XOm9EmsdUZBV2Kd3JrOxdE
TnQsvXnUTy/1IQU2AF5YzDi6ZwxEqUhoi6JFYmLb5XuhAhtsNX0zAWgzsdSEpY2fSZVhKkDDUwI3
ZowOJP9SGikXhVnZsUAP4lGp+CZFpD/lQDfnZFlK9upqVr7BeX+QynSxbkUnda3Xas8V2iLIeWr6
o54vOvjNKdgFAUIoYZjbPwpiBLSG+ZZ89ktVwFdDvkiwHIFokERVM0oLhaCdH9dTH+PUlkSZIumQ
Pu7UTNmrUqui1i/97+UZYyKGauNXuGm31JH8aMAKPxPLP6cpA3AlUIFg5sVSIAkkNjDRyV7iuTri
JTocQ42/qnd981jyn9idKC/SX43inOvfYzduSO7uPP0v3ZI8hEJUPnIHmhJtSFJ6Zx34OAoRLQZQ
Wre/Ld2X5uGP5ZThLuEr74uG2eIKx2lI8vyyBBxUAWYAFr3DwMSdU0IiVO4B31gdNE1ARjOghsqu
KmK0RyctoekOJlTdusCwOy0c95qdmg4Eo6qbV6Vj3IDq2VwSUKCt2k6qYKgGfdTo13RULiDh0Dsi
91fiW5n9Bh6v7a+ZFrqAYxvI005jYeV/XdbC4WFazuF/ZQrBKN7BmtRRU8gNS+g0R1mevU8zsSCU
twJvTxDH2HMLxmi7z8K6+ivlwmc3unPqn2TcwMzmEQH75NT6IkYcsdMq7pUifFZEZlASrxHI8yYP
XpFZ64V7ZMbT5tbOhB7L56qbTgD7dp2CzQMlo38KvS2xTChltL9Q+82H0wto0OuSj+f32ERHHFfw
0ON9th8k6Mgb96Xb+LLA94WRW/inrsl1H+IywlODzAtwW+lzCowk1q7GaHDlkIdG3euwAyVdeRfU
u1RLOTiKdCbDDKaD7ebCSfTXymh3AHZjqgiQUXsd8DLgXWe0pccdHX22qEWKR/2jPlRYVCf3fFcT
0Gti4E7tfCPfE5nck1WkfxgN8/ajztIax3Wl04h5/mpmxDzGYWMfPhO5iVtDN8asdnk+StmSpvEG
UBA5bJNdbPY9jEV2ll/U5C9O5vVxjxRznnPTWAv93zTto+ByXET3iRVGuogN0xmu2bvm63tTVEFF
tHlkzhDi5viXQcMD0by93HtUracljGj0195eK4SjvPgZiskK/CdY0R08aR0krvtIiWbuiKV1w9/c
YmdvhTPfkXa5kK1DDrclJlVYv34wLdp81L2wOn1IMKZ/5T+SyJfMXQEp505unf6SD+uLq6UG2ekX
uptCajzCRJ30C18ovCu7Td5lOXZ+P3xhdnFMvelEiLdAaOUNxisL6laIvgQU+b2OB4ZOS1ljx3E7
F8OV2+4yAyOVYgTV6cB0C8gAGWKBkfXaq+EYC4WBt7vQrogpVjwjFol8WrSAXxCxfP3s8kWChj3A
U0SfDFoViR1xvu/gHcbX7xUkyjZ0nGTpXTCLmiZ54FtRXe4qnnGrSNPGfAgzNwkjTBPm/vXUTC+h
Dx+Ck0NQ/gIrdZ0JLqLGmo3DY0fRVvezYsK3evF3rn/0HZcMoZQqjUuBOdTCK9/iiXnGZQv2OhsH
v/H6twdcBMfGqxwSJ6I7VQzI6J+9TvGwFtqRWL5AT35tUAC3Q7SAAd31VvvZQ0U3J+4PHYe3VaPe
uL6VfqtvcN42rHKwTE+n8CmU/xod+Onx53NE+EdAP3iB1EA39mpm26BNK2pceYb03OezDqYDpF3k
5waUYHMCsZZzItv2izNxRf7DmCTZOEl9yd0rUBCtd1zx4MsqkU8yMsbC5U3fuFonuTcm2YRyxQ2p
eHSNaO8SKKH76a0zR7NrGh3FsgEOgTsZgQktM9Gk1myqgiE967wBaUQyjyunRnjXMZMZZbCQl30H
iVEFmoAQ/Gdrq4Bc3smNPOwzwh+/YwrZ+vURCDdFME6cA3uaLmF8gSQE+nbJVF10tue43idhoge5
SyaG6qmc0JKhXKd+b8hk4Hxm07aGFclLah1/p71cNGJuIjniZkma5zbaHzbhN7zLA/yQQZi1WP9m
joj3CR8BlWqQHwTTTR3vC4znxmjTZ/ze09VT7mrq1aH2WNS3Mlzqiv2wII9BcQKjc3XsVrHsn0bB
YYCHCkfwo+jlwturqSfrQDw7ha7I3wyTqDDQSJd1ILe2PD5rMKPhZkWU4nxRbu9v56Pwan9ng3I0
uvE30QWT5EMp4sBRbRxva2SjHTFJARVBITcyonT0a9F5uman+jfEEZ8BZwV7R1nGuCCCY6R1geH+
15hrzQ/nP4+Men6aUM+xG43y1xBdIcWXuL5R93alol/c2+u9HhUfoinOxwKA45nSwAea4ZcS9vbm
i5spXhve0/71md4qQG+MZMQ2bKFxzMAveRfAIY3hcdibGyq4bjpedfRLeVhP6rdiL9hyfmzOcig7
KkrBh5hH7yLfCBfDZcsH4mXDA6rvaDIuoO9CNSnyuw4t7qwYvlvrY65DuolJQ/EFeYs20QcX+F/t
CG6v3S/5UT8bbJhkc9kWH3Le2CulGVTgHDZ8Zrbt0HHXR72b1Gc54ntPG8oa7wj4aizVbZ5jRkf8
30CrIO2yVxOswP1fpaB5EDykJHnnMDevyUHSyJh8mh1EtD8ndNeJJCjej+UkQakQ2xD1f+B3jvBr
bj9DbL+WX2n7rnXqErCczYCq4Nj1gtEzXv6GkLlJn/MdUqX9rMbkHZm0vL9Owv+zqmVLemT29T1N
lNUGySszv/nGBkUESlV+JhC06+vEdSzEa+SKDWwxcjRaafr7WuVRxAvlPPvrANSktDSaINZ03fbq
9kzOMxHV7Hm6KEn2iODIRLB+a5RqKQe0NsUipJxThJQjCeVnoEsKVrglDOmASoTmg/yxvPEOYTl7
Jp3K89erfjoTQIa4FTXdiHK4RU8O+dvE/VrEiGFDldE0U5KZGsTcnQcieohbQdXTbXOOkJnH9UU/
/oZCrhisB0UjfY4U2kkwDVztQbC5k7oAdyXvCZroNT284NzshPYK1AHDwrrSupSSQuNuaVM56qkG
2t3MD37qHWj+qWtVN5FrAgPDsB4AUxa2qVLxR5rWTYgeN+zdBcXjjKlKQxr7O4OWR15VX4PaS8HV
9mc5Bzw4ZSiBQz2CwNXXa0EhS9zTOnIBgbVmfuyVckt74ZZBw6pmdEg5yplLnEFBudAW7YQMFtNM
qOENVcoNnIw071oqvMsYKUXrn6mQkAS28eT2ii9Ev8wyrdTNJj5SfKN7Vj7cm+qYFky11qlKsZnF
FNThwDp8KBpvRpUf/mq/+/e+hmLDUm1dfSeCDP4H0AUtVyMaQD10g3JVcQff1Nk4sgpYbjKKUfUl
h7OvWpP8VKh/xpxGxPrqjO7z1wVKJ94AXXU21YPalTphkVa5SDUXATpHVx0ijxyzxMS7wZW4NzI3
lEoxfllESoVlmlKMNgVk5TSQtCbtk4ch2jzdDByo1OAUsUXdANd/Cq+80331GsjgIC6HaRR8xybL
dBoPUPfc52XNkP7i8+nk6sssIggnepvqstTmipifu6zwehcdjFghJLcFEPxJR0+dEI1DP1ObLvAj
xShED4RO6iXIdYoa9yOQSblpfWyVqotDRMyRJ+JIuHe8g8ds6nWteCFcbvNVGyA/DgcrqJXd9kHN
MspkZKGSR7cHla3S8RNxrm+c79GLRdAXariGa6BTc81vDx0cU2+WDQLqVQNBQKkLX2yOQRJsMI6X
illa8WJLHEEmWxxM2WzB6Puj8WNfpJbsZe+b2eyd9E4Psw3y0CmVJO8/O496rGp7pD6rOPkNKu/8
YpJqLD5ADou1CGyvjpiX0s1M2WtJgUmqFZu1/t5TVtsBQDNXHwK6XzGXHsz5gW+lhsLJvK5Kdayv
8yU6vgdNMTAotBCJ/iHjI6I73Xd95l9zzAZ4cGu9OzY1D4He1LHZ5f72zQ8oWtmEEA+toAXk7l2y
F5i2PRKREE9czop/4oDTow3H4I6YHtYAmfsbj3PIGxzVoFwZ5RsMpJcM1szL/1Hyi6emmYSq4cQZ
BurAbLsuDaby2Jw41Ytft/oD6tLh4wHrbebhRa8D1kRQHsf+UMB9+ojLY7M2nUeS9VtjAjKbFZ7K
Hagerckx24QVGV8B06OBYSAhDt+VuHhPykl1OSAzsJaFfEXVMWonEgGPwV10EiwhZMBeFbl38b2d
ef56j1qSlySJuQUhFlkoXzuKyCrLJFH37adphmso1AhP/rzGW2irOGZqN30rxGMCWYqlJWEAOp3T
SWgKNawWcgGkXzTvTCbI09Ss/G2q6ZnZUG8YHfk2OsgP1ufCAqw/fV9Mt9yQ1RnJeAXbrPKR9S2z
OvKV9YgodRtR+70SEDt3NljnIc5I7DMzarHnHJuSRRMWaUDABM612d4J49jtR+r7G2HXo8Xv8kvJ
N70EegDjGRBWibc5/OGpzDyalNwE/Bo2lBJTtay6i7Y4xnik8InDMUWl9KjKnseOfymX8hyg/r7k
9xjSnIupn+KlrzL3fCHcfSFUvzxPsvUWCKrpJT5iisOnVLwjK0w4DhtAkx3E8ZD9EO5DHJeStbNW
YK9c0YhpRMIPdO9Gp96eLhcvRqK/o3KwpRnh3Xv2cdJ6MnelM7noRGESv5ljcBfdRYCtV1c+mFov
lXZA2aZouwYFF+V0VfqrqqfwLdjUSAzoqX/fBddQgp/3l0sm+kN0gu4nuXdXRS8OaLHbpb1Bqnlw
iH13C+lN/GMoTRkDXSUcktJLWdE1S6EEnnOa0U0TOIbkPKIorjy+P9IILtMu77oa9wjJbSZcyk5H
3GnwcHiaAxA2amVCEMXQYb2J/REXWsygpJSLSfQU51xMEowr2na+4pWr1f5ChFmUOU7/4ccqOaZt
3n6k8183JZv2gZ61SboZDGjQ6yVcFjC66I+Y1NNhD05lyjzI0nGqkDM6FHVPyGdDRxTmL/Yh9Nig
QIgnWB1WX3Lu63NZYTPDldsTleIN2UgY4TwXGPu+3lXdWwqIGDuzqFzB84LP8PUXDfmrNGsHCUQQ
x345BtKNdGMvuZy4ediCMV0vyGJzEwCXbagDDyZAQEn9gVflOKNn5wSjl/03yuQFvbXwtkiB/Jh8
PGp8+kZ+UIgc0M8WCgGwBlEiBHB2wEHxspKfa8uh6FkAoih4HAqyM1yVZNUi1hMu/Gf/PmO2eUu5
yf2vMOFXI613ePaQ72I7GlzQ8nUeSoLHMcNXWFCdmpXpQPRcSHOd263xwLTFl0XjeuaMVYUw3g7N
EnrQ6LG/EGdIB/mDmZKiElyCQgFnEQ670Y/Xq/qYHh1ymVO240p5Mc0Q+gg6d+HB1wsL4J6gXZ7Z
DedWDSGqIj5koznxS8CBiXjOT2DFjhXbXL/JkF+HJ8U01+4IrRFnK2dQygvb7iHYAcP01Bl1tTk5
d2o7O6FHbcVjYqenMw6cxCxV0WLUn23JW3kmXaybHb+ECZ22A57by51uS/myYoSvH96gtjSVqA+z
C/nGUmleGMQZEBtgG7uy02wh6LtjV+N2Ph6qyz6R5XLkuOGtA+KYi3HIPaHjXm2b0bS94+ntWpA+
jZxkziwBKyoJe5vfdY/owgpNfehC34FlXpGKE4PVKwBq+SgBqJxiYXBm7MH1z1EwpEscSdslQTjV
z3x08sWGUj2kWfMkcW/mZAWw8qoOnDQi8LUns74fzXC5YHnO4BZaUZgReZFRXQo/HBA2J0tdcQm2
y/cIX6cGVG/xv5h501HB+lxpqLqVVWP50dOamMfU57t1O2yqjWfiZNChwMgg0w0a7zOS8I5GsccG
ReAPEg7u52X0hilNUJCfK5b1GJ9qRW/ccjqrtn/1mMac8fgATqXd1K0PcDUNHWnpt026qwj6QlRY
gRCJUUz9UwORZXhjK3+w/yy5QJy7M0ENR4jFCqv2KVXbGMRkm2bVLpgMy3XkLdLY2gkRWVjx+RKd
tLm2XzgvSonWd6rAcdpbfxXlRTVdKcSBVMpirZ1ZLCvK9DVKBO7eYKJIGO8stHtWmHmqYq++qLRN
GALKT4j/xYZeHc92GjkS44jsgtCNC0yITiCQhvB1WkrgkKbdNHidU2U9QyaJiImV5GnVxhSu963c
n4bBb8eJLXI2hYxpIQRw3RENZuQNs6qS31g3ocBo5BqOYPf5YAqENb76+952fJCYoccbYICJ6S3t
yndqgkPn6HPSpN+nf8/1+CWTXhyHTh795/GI97Wg1C0+68bacd3LBORbg6thWi+fsVAWeOUlvZ5/
FJQOBXb9i7rcIvmt4lEHc06ZPEwFEj1aKqmOvN1FrsYD5j2CNVJpBGD0zuNvfEovfosa81UceoQz
JUVtZmwpERuIVQlg9aRNd3Zl2KHAGtR4AGO/0SPCCkea2TbgmBKdeEimdPQGEUVK9T5dzHrMwZT/
xPlg8H7quRI/oXXdZvSJVEWAmZ6v4v356Yj7U90AEbyvsgrItvEWjOXeA8BfdOJT6mkglwcrNE5o
YVXd0wjB1mM7WOCWXBCfx2BE4+snJmQiNxiUrQgcEhfibDWfk6EE3rrwva/Uv7/A9DBAd0D/3DHm
lMafm5T0kbRWJoG0ndBlvS2imdz61aII7fadHfOc47w+1zp7Kan1wEv9fNGcGOnqs35w07bX9Mk2
aq709vIEDdDtLH1zIuxm3pFHlqv4bye0bPDG7bS8Vpnf8yxOYqgDxFpmf6soGuAeDaFMVjzr8qDy
GoxuLxkdtyitH+ZIp5BlV/3lX601OKF+F5N9LajDH+4Dhi0LJx84k2lniXn8PYkVi/kTB5cQdwNS
c2r+oJRkNTIS6bXMQa6oV28V17e5XF9qNAjlwckuVpWVkHQ5brCqwuSPlEV5uYCEX7sUYDWZQgVu
KXoYW7ouMEN1vk/ZYLYVfJBGi22EnD9teFwDy5AsnPxMEg1jElD82V9Y0U+gZFQAk2p1HhSSalJD
gxAof6iZ+a3NkqQIImq7zOFSHw1veCIOnqMgOGoTkYAhFMWKEBdcuksFPnfTPv6EiHyOs1XBkowz
MhDObLn/tBjdPriTtOZ/pk9NMq/4cYUMKz8nv4m3D0vVPKXAKRnuF4FNlSpZHRmrBX4+ybvBaadG
gdidfbJYJ+o7drqjo/NYCKpn7l0wy9CfgSm7YDYCQmQQDWu/vlbUlbpdxAufFPVMpwm2nfDPLpZz
wDF+zqmA+ljmwZgjxMe8VcRyRdIeRabKVx2xuUqrVMuO19Pq4lyC6ZlzNixoTXVkBLQ4czpE0xPy
zWZYrnSdfBS/GMgZMiupLDEv5FpkQ/8TBn130AgvwKcHHa4VtI/6T3G9olhiY1FMS/nq6UmCRosd
MIlHv7nhaZEpaUNY/i0A4LIDaBhSMS5jjtjXPHmNYm7EbxVQDLKrjeqi8pXIZBeYGXZDCxiuUUh9
/8LROnUUcM9lZi9igtaxTd4tKd704cNSI9flY4uhhzFFIvhvOGEwm1ei460t4q042fntWPjIODhi
hxI+zKx3n91leNc/e1dv6hfWa2INlcnhKluT+GB1ZmYODnmuO5/IrgZXXuN3MBBXv82Rm4Kkq3mV
BJTyY+8MffR75itLqEkIxCIuGA07IZodtKXnsjGmPxjkEPi+0ov7xBnmyPmUMeuZJ3CzABuaxPjX
OCvdKRfimHvcPB0F7xUwaHvsQkTzDrdLay1YHBHjQ9kQUnLumU5C8v70274rW2NHtCeW+34oP/Fd
IzGgcoIX/sSOYwhYjdEP1f9Vx1kX5A3vxpDJK2GOYlEcL3093PtD8lm3gteC4i5KKH1ZYtKgoe/G
P/263X7adcUa1ZjGVNZFWXAYUHLs7kD2ZcFJOlppYgRfptiKsp6+b0gg9Eu65g4hvex5ZRsde2kn
umz+KpCHQnLelJarEAno+YFzx5YtrJxY4MZ3csg7VNi7rpG4YY5o3LFHHjQK2lfN/8hP/XRwNXSM
ld33Zy0l2wuCoQoJ+hW/qgTdKTeC9dOVuwJrEctw9jfCvf+OIjM93Gzr1yhJbgEWgciZTuXVMSV6
bG74Hx0jHkikOygFfGkCkFz6HmcCjWhQSiU/+sJGUVZI5VGqaEiHsKObFkHBYCpWvCDv/15oX+Pc
zXGde/JpdrrYVhZco95BYBtozDd7AjdelKMRDg9bA4wyXo0/j6GZIaWtNzC+VBLGFCpE6H/x6hm4
vbDRpTrcX0qYZTA3tXKq/ffweWMtqOueDWBVGn0nY1bMcH/6lNvlqYIdlZyKY+ofhCvtUYPooD02
DbrVQnGAfsDlEpwbkPK2Z3wtSdWx5M5s3Q6kTTXYoH5ge7xZKoajVBgHFlGwqU+mL+Z4BmCGPd1w
xBkg9+0yxxwTp1JW1TpfbAPOY+nHN/Su03plfs6Qv/4YpHB10TxBMc7uh65uSedUG+gQBM9P+FXE
yzHs3z3L50jRXknFsHwJ9kJFd5TlxqLhosY0y6ODwskGhP1Wt5W3hDAtfszyYXFSxAExrWy2rhXC
EmcAOXfFcSANPNHir1rWuHGHamv6LFljxtEqgH9KjL+77WvxYvxH5dTIrZiTp1fHlsHdbOFEWdTI
WRf+gjn4XQsc0wF+43jZlsS+8Cybe2mHpR72KBvMKr547xWqs7x/H491ir6uBWqvZHRGi6TxqTeg
GcPapljEkYMRcVQw+94VG+HgQa/zUirkCURrpMshXcsRYE3VwKfEyn9rv2KgjS/FA8IuiDhqUxDC
TXf/oMKRAmcp6N/XXlcALRqPnsPvWdm9d99QsMXJrXUuLYGa1A1XJpTUR4Dj5LQChO/9WRdwh9eN
gOCUGvqa2taIfEfWSFHMx9bsEDjgc/p9LKF2+kDGqth4+/yGie08vX22z0D0O8QMsH6MzA9S1E9x
nWbRAjXBJ2Ig6GakXohM/X0tzSmoLopUVYeumScZh/ng/d1MNXZG9g/x9Nn0vgtrIV5JoLxqdk6/
dzaTBljthJOkoWOlMcYSspZdYp45UOrS915fw3pK0GwgdGgWMyevkZXWlKt7quZpLR5oh14s8a/X
pywj9lHkLPrMUTrCm6Dn7Raz/2cx+XLJHFgK7yGNMwwk7Db1P74tayr0pKqlJHsLD+N1z1NyD+zE
dIdV84KbRQKmb6lWAI5od+oCOVGDMY5bseJAdRH9gur6EkDAOKfJh+hLqq/ylusatxBzZeZAW35P
uqQx8SINUxmSaFjuDTpoxV0MuvCdXTB4eiUGmTndekTeS0ZbZe9H7ioaigSXG6H4FYRPz5ORoV6F
vEYUjQ/VI46VTWgzoN9nM9doXH8yPGyCWmmGBnoahTNj2zHpUz1mhrId1x/iPnAs10ZQJtS0mEE5
mmNv/j6My9zzWh+j1mM+uAvdMCwZT7w+YDDrc3Vpb6cFouqO4PkxICMoCNnF6RNjUjvDYnGjjMcQ
THccFNen5aUrvB6UhJAPlAxHbRwy6K9BWJTXZrIe5/taEVMH5NoMC6lAtBc+i3GeVLCalYRIVlQu
AV+a918BpgpxysxUS4oAikN7P6gLR4spgHqcCvmiA/yxpr+sliB35qsQ/t39H6AiIwSXYSkoReP4
EGXqQZ6i3Q14lgVuSmoz4THcwUcEDQp2k7XcgyREL3PFbRElO3KId9vnmnm1fEjXqfhtPfWzgfZg
OSB/zg5GF56wp1Ac3iX/ugpotz4qmNgbUAiXYpHCqMO7CxlMeIL0LcHuflHYEPhgPCkTmuxVCEnw
Ahveo8fBm+U/Aw7ueIl9mNmSuUIwRPGYjGx2/jjHz08MAPMu7jxI09azSOa1CePPokU3AVMFJgT7
ArLyKRIpECGa98qKD6ObIeUq0pRJJhO4DL8i6ZNHHFDcHR0TjnJs2POBsvb9Bi28q8zHjpllRTyF
wq/vVnj/6xixHqG9eHXyBA7YLVye/c6quPm4cRV8rzmw+MjcptpEcQ1Nt/7q7fO2TxexNH1Djr9w
g04MNkTRkAz5b1JOZtXo96emJH+aI6saLj6xlGXBnjhE6m+e1POltxFcd0JN3jkEleGxBt7uN+yL
aVZlmJprv0bhBtbnmKD6o1kT7ouy8+oZJ+kUNQR1GVKkSj+Mo1eWZ4GunGislOQgD0ysS0uCzphA
4pO1x0aHwo0hn1TLDzfLvrX1G7V5UmeHCmWWUeJtiZGv0uqRpTJgOle5YjZFfAlEBQYEf1B8OWr4
zZC8shRFrh5qRm/59NPrf/4tvoFZVpZBrj5tyvK0rjk9qmq8lY1CWxBhvChZJckPzA8tcc5lw/8O
arBjrxUWc5lULpjQyipjQK/25IOaP6HHV1lFrluAiS3mqDxw7qQVawv7wQ71iyzQcx1Hb3yzev+Y
6MiRvxFGeufqA1W5/g1/4OfRzI5QJy7pHhqlDbvHW5JEvaV6sja5c2YWRFs3mvpdFr0hNiyVzPQZ
pVQVvj5IINbis7bgN88VeFzacjcwyFf/ekIguYjBqNLrTxK4ZHtN4dL9OsffQIxlimY83br3a+vq
FcwlQqfgt9kXYtBcTxtMCF2amzeOpnENyTb4Bf6SAmEcvCiF41mLd1/pmm1toLMfte+LcNgUy5Eq
6Qd1fY+Yn7DS9zp5HUhgl7GQ91+wpDznfVKrSlBM7HC38JDehGhiZhcZmXXN7hu34qkqCSYFSotl
ajGXSrkmtsmHpBSeBzp2TxslVpppRlvh7BvaI1BQMspZwmX2IbLLrzgiCsQ412gqqdbE4BLRDSZh
u+y4NIxUHKYazXYA9HXpwebfnnqzsYwOfDXEXsowH/coB7YwrS/9p7Dat1SCAcxYYG/zwRTvenvj
LDpKDZgUgLeu9PRLkqIaBs9a/NiUCrxAOD7r1Dqgb2EhhS4Uw+nOkdaQbdppKGenYQLc+ivqix6y
GQfhKZXlS7PaK2LJ0HX0DtuephBmLyNXLkjIZWWtd9lt9MiiBSw93604JfYve9FcTKj1tl18xh4o
bf2e1m5Yws+bJnnU7I8NgfDwfcbxBnSp+NJm2dlurYjVm09uX4RbbHqNphPwzakrnzyEcZmOmyq5
nXhPP+NBZZZ9yFIidwyvRpKPQ1pGtzNKIxz5z6IOZ4/jCnBdrfPBC2m9ZlpWPkzuxCpihEHv95H1
M8EwTysI3jaa5eUMlcug+ZLDy9uHbn/MhD+cfqZ2vy0fHQu9w+HPIJm2BPHtEnp1EfaUyiAitDFz
M8gmGtkqf+WcKObKEIXzRaYfE9F0q3pRlGYBA5S8gpDDYV8w5D8nAtTCilkLXLYQMjxLpPZxDRmN
+joJkuk8eMcui4J4e+mj72ukAdclN3fsNpP3nQSkmALD+a3cz3T3wehDCzNfwZmVZmgmTZlyEo7B
AWk9BPXhXXail2NJ05c+F5WZqLU+KWeCAAJpqTU4E8V2doqje9rkGpOxEuq8WelMXMUO4DI3DSTg
enOgxa8IQ1mMUY35Rhx4dpruK2nvnTRpzyMpKG9FcPsJ+aZ86LrdbM7rvg9Ij/nRcHN56qYfFDfU
pymnFsjgg6zbIS03ieE92jTQmzg39MRbm5Obn9le9CNgnB8KuOkY9O5UgiAMFEpj7O6dQJWPluIX
XO2l1tPgCXZigLbXWCeZi/s0WqKPLb5Pq7eg6YbIERwtfuii7+jJzDf5fPY3KaPMlkFzNaIusRDd
jTZ457PzJPcWC6eA2JA6HJMdhA6k0WVB8IBPEpAKaD3MV0jl03+XW2FiwPfZwnL4vFV2AROHZmat
KjLX6hLJwuv9gFJOqjWFfGPAoO3XdmcexyhqJgMxh087/yhenB4m3Iag/yoJwpJnlCj7GNEwcB0e
hPYD7Q7/dmcDcq8Gou3+QYlXufV3fZAES6bEiwTDIoISI806CQ0NKZL/Q2t7WYmtcOe/4X1u3uRe
TQDNMce/0oM0Oo9t5W4Pk2oQTYDxkCClvyEU+xjxbJv715lOuAkqlscaAnWL5jaiU66u3yKx/6fW
jgXIqnBX3P6XSWqkhDWa533HBUCFjSU4aWJDj9IzMrzpHZAw2Y64NTJmzWfdwpfVd1zI6AvpngCJ
aGkOxJl8HuNXSMydFkHamCNY1P8KcRZsRsDFMghiP4ltnZj+p7bhtuyE23ObHFoTD9YfCw+hMk60
Lx6U5Tc7o8fqUqmJ3kfC77yJQGDeueatLWZ8lbrqiCLR198kCYXx57rkOEFB/hjr34ti/FR/4015
kd6FPzSulAezra6aCNjz4f7Gu4mUjLmCVW08EwNhPnkmQtF0UYVEooHlqPmtwp3602HejU4BFb03
ur9Nw6HPVevv9bAk4bKAcl4gMLCAai6d6xz6xiajPAeE9/3JKOtYTPq1tV7jPNmpNONzrWZvr7Mk
suFl3nvWN9wJssBWhUHQzOti9DH9VXK1F6VMiqFvzY+cKYd/+NTwtVR8lbwCuPX3j6QPR7ho9yhm
lz9jWuvetflPlDga7plOhbl/dYFPxRoJKSXC0TB2pi2aAu/h60zmU6JV+85/e2/rTiaSg6h13IQ2
bMIVqq8fKAWlWF/Lm45C3zb0lYGDSUejjh51ciULo8hTt5+ufMJEHBtT3uGNA+if1XoTKvevDRZn
0jHwHL6HMHUnicJmsXTP3RwJpAX7DHNhCKV5lpIMB7w4rekFbiYJCmtq3sibdkAdYkQ+EQckm1Gy
mn3c+AgixKf3ZLnWALZZfPM1IP+gmmCc/jtKgGQyMlRzbQPP26hav6xj1lXw2Q4+XTFrSsWcHLpB
/Q2fwqMIDKcpAUdvW6iqXJql2eVdO57oc+x5BaSzIrwPV/nMyL2ffmT71GFsE/lE5ScNxIlzI7bQ
J04GvgV3vGS1/hEVqmQ6I1PC53PMCQvlwEJsLcZIWubCD7d7KCDcyefSF2AlOykGzOmyj3iWfREO
PmrS1FDRcL4o1KuqGn+X0UGsRefyEGTHlNurK7Sj3EJ2jWjI1ZwOyHP1kkOL9JhMnag6kM9l/2KY
mGo/glh4lGtZ0Oqw6J6zt1L1zKvXxnQ5m+zS+q20p281QrZoM/gZujSlof8Oc6YGsTN9uC449xks
l9RI8pUpvT46Bu2duc+hLYvZ11wEBBRPctN8fnjYYWQ2Q1cdpPyGdc3FEu4RBqAqUAbmoh2g/Q9w
lnE8f2LN3bctXer7nV5nz8lDHC0mhSd4bzvpTBpEBdZwWohnXJrF43GFmJdkZTEQDdssiu08oL8T
lSaDjfvNONDApYIbLHGC78XV8QpIVnU67sRlMfqAop4ySHbNZ1iYDKMBYocBWc04QPQDk+5ADJZi
Jg0c1otTzV7N9Vu6X65VJ6Uz9FJt4BalzUkx0Kz4GeR4cmr+6EMkcgPvGAwwm8chh6uol5L00yHi
LlyHNXDowUfvJEYPGvejJqnPiKVIEtRRVfZ+1oNs/Tm9WiS5y543Ye/y98v73Z4sJFvi2McCr5Rp
diTCALibUVMeY5Ro4fM3OnBXc4Y/13SUymOV5S2EoTb4QHbmoQEhUhZvy4/LOOk32a+A0yDk1Mlb
DgSbbRoV6cdP5jrd3cP5Li1I0c0MVJRRcdGQyDVHaRrh6V4oD/IEjODSHjo/qqjpcl86zuXDIC1Z
4xvRkhBgmPTZFuZvd+XKNo1ogC8FsM9gF2nmPgYsGaQCfu6wPOQXvHSIlwXNBlpyRl3IhjnmwAZ6
tghg7b5LDkA/FnkXCYxgFUjJYf258n4zalFeZxYhWrFM3tronvSIiqkPHBLlMEAxyvMdwSVNSwiZ
QuBLbiCcL7ZwpZqXqbtpmqwIIb2bXx0b+/moGJx4iDLwV7mg7t0A8FVCng1MRMyPu8yoGkY3cHZi
2W+bHykofIEUAlu1RJgQCL7QFiI4AhYJX6ThBKlg08Qtq9+vctaXmvJT8eGgTpv4itqmrItx/pTp
08fjTX9e7FaZDJ1/WrqYHkRDhy1TgEfTKAzRMgpwq20Rvn56HzIh6GedK1tqiT8v46Oz7h6nGJqX
eAXHuuhQt7s5ia3fvTw7urDMLmeAEtrO/hm4fvny8w7qCnwfZYpQ1r60hDjoYBOHeK/H1EqsmOJe
+6tKQz5K6A1sDoyN8/v49iEsbxUnrEpgLnq7B6k6n4hvXRp0Ge4gHPEf04uVTHmfWIzXG72FDvTg
GhVRPTkLpouNJpCigMZbWKogIyTkjLdkVDm4bh1vMRCSlcN5jXLRkAT7k/duvYwspAOqglTtHe8U
xbkqwe9vESM7H3tMkPBLAV9NUuGGYEyYNu6Y+KcJVXgTsj6PrnsWoZct3XlZczaWbHNLhj2kBiBO
cdgwBPxv2f7j6TA5Ivd1EwcqmYHL+Nl/n7YH3paF6t3E+KpXx33UO95WkW3RE5O4/LNnz94pzOI8
kDXFFo8TqyGFzm06JdUV7sf1L6h/kF1jLCVDF1W6TT8N/r5HFxODYrvkGJrAemVzSYsArXMLpcMn
8qgJv4lb18W3rSugkIEkWfGYNc4Ci/lnxFZG0iDx6tXu5eqr++W5jxrY0uanh2xpZZTkTjGYZyfC
9JH++YYqUSjdVRuTQ6PZePRAj174NURVF6kF3i5N1VUinJeZkjYRg5XXjMJ7RcgsN8Se0tirzHEW
Tc5DluZm7MyJj20CbY0MmqXFb/dJBFdc2tDPIuJRjhOaFDvbVSTO09AKJrjS/3j4+i7XXJCA+K5S
iribD2MPctrmHkda7eIqckppssiZyTlDnlSq950PBZNeAIB1nsrTsGqZs9wzdUhx6lRQ6rM8Oidx
EjXdwQzCaFYncRANvhSZf6Fjhm8+pMQJ+dnTieQO5HkrtLaKsLIqyXawwolbyMLVDqpvTv589cmB
BJPeY2qoXWXGMp8h26zPHyNUOCrfjCNUAYk7PNyx2RbuOGsc/SNUlJCOi6P+JYLBsiexR1W7ndcT
siqSabGGpVARehrpy7k6q7t8Ov36ebQG1zp+yFzu1gOA+Hrs8bLpAfENXX0viNCH7qmToM7wFv4+
GhsEofoWD2ppyQhc2bG81RbRVOF8tKQ6amcKRiYHPDD5/5vyNkIbOgwV7SeooJ4csx/yf2MX4JGX
3EH56T+2EUbc7r7vMh/csYO2oOduRX730TUQOJ7LUtROYMfdHlvhKAsh5x+gbSyHyh9DiIED8wg0
SGHiVoMs0m2mVXAHpG8xrEgx6vWH+xjfzJJCam75g5OWQkeqPyQV1g+l6QgTbi4gC8Aps/Vq6bkx
l8gCalEsstkBU+U8fkEBVLxodvrqbLi84NZMryyofjra1koqLbyzyDaThVIRjoYur3lgm7KJuE0i
rSbRJbR1fc0ttTFGG+TaN/A541egGqbbcmAbsnFPqKknGyT3l5yQuBY3QZZg8JrLP5tyk7LX8E57
abI8ctO8sE5HzQTUEILCYtUuVs87JY72JugO4kRz+gq4zhaLzROR+DwwMrPNzyWyobdJ2lLXaypV
ix9kTPHp/6kmJ7Z7B143uhADqqfs0Qizswd6NwTNpDv8aDOx2twdkNlxYS+CVehUtgEcGEKNW82C
tz9IvMQSugFDPJQaeHTKoQspx5ywupn6Up9GM7RPjalW2z+sqHgSAZN90jDcUDczHGkZgmKBgHk8
dmQDtBFY0tVanFtiXWWj+ovBZCPAgXKUs+CIm+hstLYlyAorMrGaVfr9YSJ0rX7QsMh9MfXwTFi3
E3OIXLSmgsvbmynfjn015CVr6KgmHiDXaz2ZiM7cYESflw3P2yvCxIEFvJgpH0UHr+RCZsJYCq56
Npo3Yqpj0r+p7P/jcwbMzFHbsvDEcYnHhPHuNMkJdJS1BB1cMJgCaKzQeUrMZOSIFXh4VfE6b73g
9p5Gi1H87Jivt5aavm/Uxz5a7pnpe1/baJA5/2mAhctqSdAG8eQslzl5o7cRKyWJNK5CZ18G84zX
QFCQRBGZmmrzgvJcphGc45/QnFeG656ISz1/mWW/1KSHuFKOmAMxyzglXHafWAtf4tsPYbLs6dQH
doqTWYYAkR+56DZbVl40VcnHsB0y6qppZ5XXmBiU5ebMLQyz9g5ZYFiL1yxMOTkijdZRv8nmH64/
FcwK4+R+B8Se/rDECiAr5/5z61HdJZWmelcj2OXRKRBeHHcp2N0+QRt02OSvQaINb21K+bPkUeGM
hKhIumSrPghtgGCCqPE60YHKAjczcEPkJYtdLnPEtI7tF83rspB63ZpYqnHegOj+TMDc8E5iw2mq
2jLSlDkac+lp1t4axF2yB7W3g5W8YQhCC9JFs1GT9dXX6M553ShdssNzG90VMzH22hcJdq+/Tenc
oLCFkOkG1oX98SCUDmn5SKxUMU2a5XqbdQD6OlHhl+50D9W7alfQQCLS8+W9NRH4G8l8FP1NuXCg
zVYJ8vaQjZ7hklLgCthjub3m88u8FDOVD2+sxJAG56ybj9keuD24IT9YT10j+uWdxS8JBp7Ylph5
4oeblFXExljJzj/uynWqMTTEkh3u45RFZ0WbkhLZXLb/MCrCExqRx65zjwpAPyHcfZ38+4hD1Ob1
b3neOmOh3d2VkTo3VxqSn1CGC9Z24eqviYa4vGddV7lp643SoSAYbd/7208DMoO4en82Owxd5+qH
DayA54lJTeSBjo/iRLUtR9aQkBT/x9hXvUYxLTOqGWUxxRitoT9ItIeBy/Yo4vheP0NcnNgNiyuz
pUVbhr6oUF/MshklBrVmUE6uBoeuUG//nnBj8KRv3dEHKLmaKJ84t2eYn6ub1Dm3fr2i9FZqxbz2
UhXrVGSTManx98Ev4T2HyKAtX3E0fqBb+Fpla1c//lfhB5V2rF3V0VkSKVemVAYirlyAhfwc1wrW
vjkewY+a9WzQIwtMIcckgkyObMSPUBoa+0H20TrenTpbScL4MGEgJQXZ0bsr4N8kbsRbjyCIN2qC
RrYNs3jVyVzTARuSr9tHLx/jJGMXToowt+Yif04sUWicv0cPU/cPUVzvv+D61zYfhPRr3AvyOPEY
FiwH/2Am8X6It6Rcadenz4+RfUv5uOtAkkTKlE52RYiyqSSjAkyaDBLxY6cET3y71yUesjp4iWjZ
B3lBy+qWZNIxIo1pHFC0g44M2MDEdAL3Y+OG2Cwcbz91dovF3SydFGCe0rgMibYB+M4Ak5YiGCqz
kPHJsod6u2g7XPvX4h0j+dd35V5O650Cp/M6FHjNYNJzRGkkZ3X3juBnxyi0ZfX0FARi8v4XKRRo
9TaqhXhMuniKGFsXKNROaO1Qr86Nb4jW7k6gv/wE4n59k+olVd1z3c+Ng/ndUAlElCw7IG1tjWVv
WBbM4GTbmVkAHTubfM2L3pEkujS3u1WR3XWrBzgoiQ4RikVrT00WJNt5kaa3byQFFabKlsgF51NV
Q7MbDOmqvf9ZYhLHS2FzT22N1Cwn+BTpiFLnR872ZDR+47J34JR9KPnaWpV140fMDMtMzKbr0ukD
VNtf6iBDmqaXSrKg0KufPWvL/8U0894cKNRwJeXTMUBV6z4hNPNJ+1quGaZTjgnXZ2MF7wjg/nhQ
EAnAHQd1d/v8kGmFDGYKeQYp6S5dSHSpa8hFIaPEKU7y0qhmX88iKiyQih1RB/J6HFu4mCoy5kid
/ThXH1RRgd4FRdqte0+6bh4hrL84DnCrEmZdHlxbnV6nCqqWw7K//ycuqrc3YLPQrOS/hOkcsjQZ
r3m3G8YKUhiTRCQ+Dh8FLIlxqdJ55ur5fqLaIEI6FbkznOoOlfoOUdi2sY9Get+x9FuFVOkanSo/
bhW4Gimt+zWPP/wV8j4YsebAf79uVDPygB1pYSsrD9EuJSsZ/TmLkDnAestDwUU2CytpxpI4HrMZ
+TaCr0Zj2iVyuWcitx8YSeoFX689R+snMlWhKZvzedqlrUmR6kk8U/n19UB59HGuWfxQcaR/N69a
S9a1I1s2hBo6OmybYy/QWxuqUQrd2BmDK9U85uu4Iz/1KjQCcZRMSf3RVPCs4vY2YPCy1nG5gt5Y
YKcu775GU0wL10AeIoOyIjH6w+h3SaLBZEKHMwtYr897EKPxWEk/9/nhJeQWPOBRV9cEUAPHxywp
wmXJ4YSllfD++46eS4C6HQln2agKQqs5witvbl8TMWOiYcLI34nyfjS9/vnz7Ctrd8Gw8vmB/oI2
DsCjDQm6kykydz86pb03P6FmqqSW0yd2hNwemS6e8pvqoceHizpWfpLpD+a+UCa3UqA+oIDa8qtT
fvFkeQW/UfT2YeLnLfyJxadqCeIyvCDqNFFa7R0YTEWgYyfD7JjJ/H3/tqWzusyIrnFsWHMgICMw
RzkSSxbqpn06VsvQofxMM6pBHLVQmZgycG2G+D3kNgg2nrNuxeHVJ1bmoUAWcrYnlN6knPSqvJdR
lvViVAtgWnGfAf6eUCT284beE7p30Ink0DJRRA5KlVIBFTbm4Ix2dSxZLxQXEibO595bF31eaZxz
6riokAD5FhMZVaxK2999pXZDO/rKbVO/NxCOH96NruSL8VDuaQwxFnLTlMciysYViXv/5fXKB1F9
1ayZb8OTVUvONFYw2jk+1MumdUK1fFQt48StiNCG0eI0VklbdZsB7Rd4nlZ3GMzx/GgAbFb83NDY
E+eYJVOyboiCrPaNHdI0WqYez+ry9WhpE0gEAx04atDEjFk6+IW0nHjJ9+VQvJOjaqnijAcY4Y0J
qPxTIakeZq/JczyyAxF5ij1OA9wKC/Q8Ur3dSNAeIj+kUVcnq5ATnVrbxbI6eRaPRam6cfJQbFNq
LUJ4BsUhy1Xeh9PKJUVxUOMy9dsiE5g4Xj31hBIzzyK6LrvcUrteVj9/rMD/CqZS+YKKNgGItUod
Xw1RaSvuPTJ6cCOSZKyXlAJEHVgUabY2m6/WcLATM/GpB/zvBduKIhjoJWv+gLAOYzQQfqO+1Dxz
ZLkco35aDnq6tmLyshAkav+rzW5h4Njzc5j3HnyDr9F/cGN2Eno4zAG3BMlJAAkdJkGNHU5cGHgq
WDoub4ERSMi8qVxTld54YXHX09DQTPX6I1PhPsiSEYEB7rmYc3Hn+3V8wDM1Ypg9YvehYljwWbkv
BpQtlpzbDaIbvNbqMT69RkfTAMD2PhMgHfXNuN359uy7pBZHfrPyyTttr19F4gweDgpzntm/CD/s
p3lwwAuIAsqMQPgvsJy+HxRIy/ZiahuKzhCHybIWH+DZhyxoPfXFYwTP8T8fJ2UNt3e7qlVMx2On
frf3UkmZxLFsUSBUZpmzzt9bLbnhxTkc0HTFY8vDYhMJJJh0nvkgpyL79xAbKniq21VN2wEeskhF
H4ilSbFqIA6rb82iyxGZXkLM2PMMjaLllDZohe07GjOPXc/daQ+MSP+uyZ9GOvUwp3MOKDZ72v6f
jfUsdOpVkQBR/WljxDn+10NODRDvBc5SXtlr9GZY1y7F1eiEQsVh+ZgkteNhOrknBVeMOD62odPh
NJQiKWPi7CWLAhgRNx6FtcdNaX6IpwzrGZzy1Q5YARkNqgq97yzM2HEu422ADUoxfoEPA+bXIWtO
wskS3rLqXgZgpo5gX9OG3unzo6eiXPONm0aK1bszm1igXj0+yvvMG9Qi0JLdpHgxxCij5QbqBQIc
XUuyIX+FgNGoc8KfADeZbxQY1+ctSLAtHErCy0DsKQQsYDqb8B7f3eTqQN9Gnxlf5PmTXzRUTUR+
INKpQX90I/NKC5PWF5scuOCsDe0wnV0T2a8brf7xLMdeJpObE5dUrkYoAH/l0edU3L/R7WbKucxQ
vtIvwugRrPHFs3CdQFvhMPXGAEqklbJHBRAhOa3LRPsrWKx+Yr3MT9Vs2wstdcz5GtfDR/SoA2OD
3QCbDGaGv3f6p0bEzoGIg6Xw8xhVI55t8QaFqAPOXu6baSP5Sxya/I5x0jL3pQeLsQuuR37zj7ZA
8G3GSGgUTpMi9X1ioVZ+pWUhm/y7pZBkf0dqiE1m94S3Kcz4hKXBSPh/f2nM4cuybbQt2ydNfh8M
z//puhYdjNL2JZyAcD9igeCglGYjSqNpx2ZBqjkALpk8ne1F2prk1clJdoHxDBwu/RU5Hupyqo8M
YeJdvZCOs4Kq1JHq8CmTDOW8zBMLyJ5SYpj+zKm1ll0RWmH81t+6uJRjjnDgFoE0v7NzPj5GAuUM
I89wjskxrnEvLocJ5EM0T9bvB5xmphQoDf8lwAmaApPboVjWDKdl0D9QDI7ZL9P13KEAaARDibM6
Gb5HADrV8UKV1f+Nyi6EfjXNabkpBLG8ey535IGcf2MZJ2Ikq/GCnFvmNsZXwyE8N/ezJe1YrUiP
YLNTOS9OCsjtOEvsup+9CPh2Ryj9DKRpjMzjVtLvu6SLKs9HHBqY9c1MWeOuK34lNlf4qN78RnKs
xuQ+t7Kl2LCygGA6AoHhnkGtRFAPJLa6fT10LlSurx1084Z+tsvRlLvlWayuGQROiHoHKDicBHVa
FALX0+c2RrKIezWoOyr3pZNYi0iysP+dKvi59vgfDQAYwoP8ofMWMmkBIh4FfOcS0cJN1HenFtig
VvgGB3Bk1VnyjRvp5nH0iGJSL8ZZNu/o6/MuuH2Dszuwb9Czf5uYVvRnNlQF4wERXrFwYYfyhfw7
96CMwqP10MgUwvN+2ABNvKBKSfqTlf1UhCbg9WCWxRuT2+Ag5BzhllaD8AdZGjMaRv8vTAvUHh/P
OvLHT8GIMDtCpcolJwgRUeuWijD4/NZW1kEOVQd6JK/az9g0R4vYbeB4RqUA05/2fBb5NswRgMeX
WmjnPR4gGmTZGZZ89JmOZ9SOiyyWydAaX1o2OPo0ELFYV7+rvZfpnZgXPdch5QKkZEWCu3SyG2ck
LoWKscHi8fYciespkjUNz4ACnvC1IITjlUWp5ynHItkvHtmiADsOOC+PFyuLuVbJG2fJevqXqWlZ
xRHBZzDfOu6iZqDZh0NK15zjrhlFg5vv86ZWzkD4kBQE8arfZi5iyeiYSVkVmFn1XEYi4IyFgNPE
qAwNEkUA28vzewkSnNKQOW8sG90g3HzbpXP73vOco3VSTym/Bx3g0qBCEpJfop3pOk6o0Oy4HWUV
UxR4JoaI+gpwQSeDgatyrB9bdkzzYa87/WztQPLLYACqQ0+hNJceQZG1QfRgG/S/rgKhcQI+w8UZ
64GecgneF+0UzTGaLFMMNBGDl+gmB/3p1lFX+FNIKja5/5SGmmBZJp3cIUmHJbYNEbn+nLW6K/zx
3jZTejH+I0vsZ/b/TmqN8FK/P1ttYclwJCl57KUyIv2bd6AZE/ByhShaWi+KIxEU3eBsuUldrK+b
pmVTG7bgcKmqLBAP59e0jQXgQpbQcpKJ2fome+72aA+l4TOAC0xR0jYF45eh8LJYaHTpLHloNA4n
NkNxxPm0hiqdx+nltgzcOdL+tY2byBbhJlaRUzrseTSBDAMheJSd1Dylhv3eKCHuEwx/1yVKyvtT
fsyDiHa8OJTdj1vk+fvJ89cJutz05SEhCjPYlzLN5wCHfmGHaktkHd0+Be+1kVAOpQXZoaN01dMJ
hr2+QCl8aRH/SvwRuuJJzTF+TMYz5RVmw3MONMHhFkfBNhpPFbUGf93WPB0j/3BHfeAAHCuEEWoA
l/KwBG3D6OngWteAzFXYljXAlDADTgg0Kuln1omVzsiy3ZEkZxsh7K5aQJqEDek/n9dPA1DoNu0w
NPKV7/jwtX/3VVVvTrb+ZJF/f50YnzEU5iSjmtXmlDl4Xls7ogx2MVxtlajVJJMr6as2/HwsVMrx
KklGhvftvR7KJ3j1evjT+Sfgq0D6HcY0WbL/u6cWjDtkvi7RznJvcr0MWINiDiDHSmhTBDtyySiZ
AOMLhpyX4lojQ73hQ7hnbhVZmM8k/UPyez5axoE3synAhwUNreKpGOtM90Adnt0GlkvGbulb+Pqs
A4GruVBGR/JIrgQzRL5pAEHRgGJHDWaTGWpsnriQ6Je7xjAOa+zK1JqSp15oJsxpHZ5f5BHlVTXj
iOSVZTkm3l7drPIzDsA3EY8zxAHmmGlbuWIYTXb0+GbTfIwAqftpq49/xQlMIHk1onjeTqnUJl2c
XuX6GOTVHhF9aQTTWesaLmnzufcP/qNN966SIkVYPcr2g+0cc0obsR7WsmH1vtO0EsGMmzlg/fl4
VS/iUl6hk8n97WV8/NIpO8WaTTs9qRYBXMYIrkm64qUMfvP3LvdHZ+QuXECrpq3H8erxbaCtfeqW
86NZP//acTPhTNE+sFYhO4mE7s6/JapLjRdEGRxcbsCfbAqsPWK7kap3kfcMbhh3To7Qjov+NI9x
XEQ631Duvr2MN7TJkm7SQcwSaK4YHa5624vieqDwhvcpiLXb9H6QslrPtdwQa6Nh/rzm1lgR+OM2
0dY+p9cMWYQNNyxvGYEaf81a98LjC9QtfHimZ+AcJQojK2R1XeEKa824dMpd8S0AM1zY/wTjlQeF
e+r9BeRN1WAVz7esOdddQ1TlS4YviwBwsO7aDmFgKY3ITlXxtyrEWKEgbaGN12RpSOHm7tN4BAhI
gCXgKAHr+RzjJoDsg18raLv9QDiGHPrsHACOUWkSIIyzmQcW6t4FDxRJQAd8GTxVCr5pkERxN5Tc
4t/+rvO2wSzvZMXi7bkXal8q/XzV4EDJ0tJd5aKJcbn3S8d3Q6+3TsMCAUFFkIfp6cMh0h9/3I+F
AeTyQjODYM2QBh9YnEWVIGTTXXrQ0K39/OfGQ7wQ3oo0g2y4wBIAFvJiORTEq9rip+77I+BnBTFb
lv5e+HyTV5NJS7hB1nBfdeT3A+BXc5NXU2bC80Nnt4OGZgjFEl5IHeVLG+qylw9Rw7M+bbHKKVFt
L5nhoZMtRkTGREbXnnNjMRorSTdtbc4vALgGC0iM+7ywSxe08JBCAIvcNjrxyc1uK4x4VK3eU2fG
2Wv7vs8w4HaOb5AdVoLsNOB+iKUJOLnKZhCOUNF1fPH78JK5sqdFBwz5mTUSnLIb20fsrva7FonR
omSnUZHVZTq8Mupo5NiaT/iavlxhOrHnH85qPbB4qcxLVoGTdFtHvR8iDPeN2UHU1+1eXwmv37TZ
KOoGh3IiRrUYVzY1ramvZQ3iUyx+mUCyzNwWoXyRYrqvqu+ZikP+zrYSjGnyaPcqYZKoi9yv2gC0
CuPvsMAW0c+lGI5DJD6NmIUj7YTyS+lZGLMiulZwa5Ndedv7bm7VyV/gXgwVldP+US65gkaCpfZR
dStRS7CfBMkBPGQtg67kuaM2YwO6E9j8I1VsCa4NATIQg7dUIZrheNfJ3rkPMs20WckBbXuXhorR
ma4aWyb10EMhdtp0fXLJYa3SWT7HH38pWGrTaKkizidpkexmkc3iWQKyvdq/LKOj1AHjb2+FaqcE
++EYigPo8xSkEs1dymQK1BMywV6mdTTI+AC/wovNqd0fnSWBhxQ4gaIRFARPKRFux50OwcZZyh6C
QCs6u5Lre03F25eK4SapTP4Y/7TI9LQ/wqQTw+WXSJiEzgcG8tNvPGRjuajnRBn4B71BUCkXd959
ym8MaWwDHp9bGuzSyINEQHXD7cjYaGO4Nb9Snzd8W2AhaKfC2/sfHrfzi+pSqh3sQzgIbocSqEi2
fuwqdEIhXkiDMalsmSA1wADAL4aWZgWlmcJLDYk4SytBsQVDZ5AuHndsgH8vUp5cvbLKGbwYwQyL
vHrtNT3NFIJtHRoUIjmZV4Hr+7583hHuyZanYjVjd7Iz9myw4KAS1MjCMr4h7J1+83itgsVC0tdI
VE/0gODsvU/A6o8WfkrbMfVfRZhyH9hYbX3cXJ2lV6/QF6S5jQIRl6/fFbxoTMpD4ng7bYdLJ3Gv
lVqY29APRb2zGzGz8HqLOL73a/pCUVXoy9xwG7m8FAcqos2WhH2RUdeerPgZBG6qakYN8cu6w79I
f12OgR7nnFFSi8WnxThYYrBFLRlMxZ4OQ5vX0qmE3GntnkNA0XrXdkMEciL9vWws0BgJZN38XCGB
zWd04qlnvms2EQl4b5nGxHeLeoZhQZxTZaAd07qaX31oGQ8uJzzOJDgPRQAfDn31AGwROYldJoS0
Ctwr+YotnK1cL3DA5VXMbynlmBWCDbrLhkMermyR1cYY4WdddZErRz6LaFEvQfPquevntXa6B6/H
MRUGIHboapgI3RjogH2pzxgZSmZzWfIbKlFVVVxL1LLN15yyC3VR0/poXzHcTUJFuenYeFkH+7dJ
TdRCYH9Vq9ddXgk8Py/RI9G0Y2VrH7zq6l3/n8JvTGtRHJGl4H61tGQbhVNGjSZc5ohnSWRwWs0s
wsNGKSLhO0H1I+fkaVNCEXYTCYoq5GF0Yg0zEDDSr8kdJVoTg2BQnp926G1it8ayVjqJhJd+ROGg
6mjxuSt3mGCPg3cr1Z5fchRMOqPeoheagTp2AqxuDlmqpnR5zDlO7aXy+Q2baKVZGxEVC5Wsi95a
kCXX9uN7fCWPc1jJcHXNUJQcRG2hurkLjZ2bHF15EE58uOx2ccXqXqY4nDcEHKkcEBZESP+1uRIo
VOj3nTGWvN5ubA19q2tWco+nSmOQBYPeRBKW/LBl82rhZFpLh5MU0fadvZjRC9v09+pqtPEd8a6X
8UmhrZDk25qXP5I1IUdEHkjVeo2MKyzwr1fXu7nUXyBl4NUwK8DJSfEfeMG4+RbFBpK4PIaRMpGQ
Dg9Igl9fwMkpX+N7OnwbpwS+8eeuxlM5O5OSZJDcCBDrmXs49kHpUQLr0kcnZdf52Zu15OysMx2Q
FxON07+GIm4ql4yW/rp75SPvKCqjHxbGl+zCqXjQrNQ0nvW120OzVkAndgvZWqivnnISAfIH/Jkm
zmGoIR+RkKYv6ziuqO11SPe7h/D3IarLTgoyDFurSeHFEgZzHP8TaGHJkndTY0WHcFPvS8FKrNDF
SP8TpQDAldmn4+kw5PGdwOM4zy/9FLiBCLMrTWocPQvOE810q5gGr45iX8us2IsE/ytgPvOfFRh5
/7biyA0tegCCCpBQRSWSHEJTs/HPcvj1xIVgHyYc0MmtIzPXk/MhN2Yj05lD+FkI5lHUjD5MHyAk
HDNVLXocRgYcXtbXwMKUsSmP7OsvSsv8U3US1dp7JWdf5+TNQgYsYH9IDiqA2fbjRBY3Ni4dVHMX
pfh7EXcqsxDKa7sNhLPDYSTYBcxgAA1zf9vFwv/tMwnx12dCQw2dpDon2YdZQr+24asPhP+PGQ3W
n7CilF0aU4RLanI+ML+wtkOP3s33L33vweS9BGXJMWPx3om5BIwTlUoId4Q1f/zoIFHCzr3AzeD0
Ik1BtPAOcHEKmX+/N3+I3AfZg3LFrtvJXYdF3cjJ1NJp7PWM0RqyKsLdlTY5Nl/m/57qAm+jbXoM
LC8+KTw+78S/4VOiG/NEF/ZqPvFWORkWk+PD8vRG8tWRiSo7MoRIi5k15DAKR9GlntUf9AcwE6e6
ETyqdY83dvI4kU9iUcMM+RfwwXuhXLROn3gMfJ5TUUsbGmFjPO5J0bYf1AmWDYER6bM1+VwLRwdr
lcg4/oZPcXxCfcFlFn19mNszgmlXqC10Tm5Hr+zapkmMGfSvRCgWscDA8LvEoKXcY9lLFS3f/w6S
yUQMYi7NjaSTRhlSOWBnEf6KxEGcBYKNUCzqjrw362CGZcZU+lt/kcvGwbOMPbB5kGQ+U2B2NwJv
v8eGvl1BHPq8hbZhCOQsuJm7NwhEWsoaUmwGF/7nJAWb4Uy0o0yKiQtmBjJeeo8iWyg6C54DbJgz
d0kLOTrb6M+ZwVQocCpcrfuIvQ7XfcQdO340Nzc02LxKQ6WUoFiwf68USF7z0KKHXn/SWcZ0/BVC
yQbjLWnT60O9cioVb30A+uZItRVi4Jt72FYn1IqoEKJDmO9Poy6Q/0XWo/nqtSTpBY3swDT4Fomi
wX8ZE24hHyq6ABAdtK8Hkd8gxtVFBTsDUOkelo+XnH2uGrepNwuKOIVu5Smc39ITCujR2LVGXmFS
MzPOolbKQnkBdRb93y8KYmE7mTl6cnMaRe1DQumVfZema4NO8cp2NXPfoz2uskT58X24MugNJMtR
/n2aUvQAGnqNn5JUxRQDcjQjBcVVIt2OPW45HC5G7T2dV6KW1IjU92KH5EkHjFMXOEIE5ubXSN/j
tFDjDo+xRzDyyaWRiwLb0WpQ+p50qVHxSdiaUvMiiia+h92I4hUgL7izdz1l3AVJbUdSr5dJ2Ig+
wZcykSOXF4W/xxD0vvesU3YV7x45U45s1qyaV9V7HfKqLozV4eWWKCP8z/Jwciabo+ABDc/waFND
Zq79CvtVTwwrf41vhnxIsA0H5GDP+LKml1AqAfu2KYbZDXwi7XAj5OUZCu4TL+R2OEdQZMpSa3NH
hRYzJJ/uqGx+KHHknGiiMx7chZLAg95on4h+a24eRlUI9I+FKlnTIPnR0KNYG0+C0r4rZPY7Ihqg
LFdwR42ZfORto/5yEFYucbWWLELNV/MO647HWR7tREZZiN6ClUqekdhs76fFu9DfEe5Irx+kihU5
2AldWm6h0YW/lX3eZGtZWeLwAIa6/fOG97WZQzTS+6NZmhQ1xCNKTrpSFVw1+nGbxgqgXGfAMwsN
pJ5+XEKC+Uxh02QvhJgkijHL2QOuCKoTTQV8MKGr5G/Cr3hfgwIDRbbRZXE+uDlhMHIqbQnqMS4w
PwcOp4EIrm38p8nmgCapIQHa9uIlhmsPBQTCpHaLKLjRHQC8ZgYq1TuynH3k5LnJ18/1kYqOtwLF
CbNyL4HZPHVGP3cUAFAxPXVg66ofhqEGk9BST7kwR82Arx95OJ+m4PvSoVi2obC/HFeHn8+APbLw
YTNHdaI8nXInpiaOmJm8vyuk0qZmjAOW3am7XsBnE58GXdtDsv1OYncOr8WQOO1lotN55+XdXfFz
vrpljzcsQr0ZlL7lj/X4VXRPGKGgQtantGlor8OVk3L1BAv5ODNIt/XME/wfbEpf9VaSiNvZsWj0
a33DT7jze5MgK9vCbzmnqWHzFlL+kgo+Ah4hRcd67QCTstN/Oo8BLB+wlJLIfco7i3z3M6pp6TH0
CC3POcv9fDBek3rTB51baEcwN7B8ypaksqQ27BbckXkmqWvOC8OHM+G7kQNMBtvGeT5v58bouXLp
FKjY0do9wL8fqS99749MqjVU2D+MmXwZtjlBby1c8ahWcmdzE+80YPeHfIzina0XmaETvunalrfJ
qXgRXhaJ/5JM87X+pAMBvyAJhynzzyeGklxbwrj0maXRzyO5j5KGFbZPCD3B1rLoHnMIPPfODf96
CqAbyGMD0YyyYhKEsBVygHYA44qPQaKFkpVMURAk+7UZ8pXsR6/2OB8knPlEqCdCZf0MwykOXZ9z
aStub3/+1YeEmGIRv4DWIQlDLL1zaJdhBvhe4JtX2BQggttJFVhJM76vljjtZBvQgAfHC0pMmg5x
TP1NsF3Z2RJcbCcO7uJSX1u99+sy5uz/0ShL5ujBsP70m7zb2uyDpBfHXf077RHjln/Trfr7E5J/
0fFQ/DDkjSzJjMxxL/E1tXl4iJJJEyjJGTFbjEY4QOGfzA2OHVigksh/bKNWipAr0OxGF0wz3W7w
2KV9QxbMvbnSfr9tdzvSuav3196SIsqRTapkZOP5ZbVhbI5BvY/WJwFq1eMwqxpHtFHtiznIMvOL
lgSPFoQGq1Smo4pEtFFBLX1I+4ehNqR2a1clfE/1I3u8xYKaEmp7Gf+bdsmLVZTZseBgrdjj9rB1
vjxm2DWZl8OFm4fVH/Z/nPyj/E+uE84WLPUw35pRhsxaP/N6qyfGVI1bKJvsp5ueAXYUxvGYe2+5
vVjnhxXYXbjLqpjZVIaMPsFZhtn//plnaXihxGE8W1hoPqX0qMdRi8biIDF5ZzxgNrA1OjJ+8BQf
2AikjjTFH/B5a4kcJSEsHoK4EMiNJ/1zzjARZVvZq4W2KgiRWZPlmgca3JHtcuDbGio3Tc5FLQcC
idruFOyGcvrFbtMW7YLB153WSg4RebqIq8B3jPNSEkb+urwjCLowXJPwHuYHuudZYNy9lKbcR2Nb
INclJgahb/7XcY2wcVOROLQV/f9ZgR/0rd/0mKcvpTG5rWGloAMo3pbiaNPFeDfKkRcCNlICqn6X
TXiJvusKh0p0bhuJLz0cmsfcxDnwviybxTucEmzCWGNZwjkEouHTtjCqXW5pWlB+plMLoH7tNiwf
CXx56Wp2Few6rGn6cm/scFkzv+X5FdGby4nrrK/tiDUuXQTP2F6VquEUnIqRW23xeKLlSyLJgeNl
lY3kQMmQX672J6riunJyLvrK9rIk46/mv8Wsgjs/X7JG4WTuKNlVFsO6AuIOqiu0/6utQaDK24CT
pLjompFsul3s4GeklM5KBnXcmECh/DrY/Dx/CNK/RYkf329LWALHvUmTGizP/864jP4/o1ypz8TM
OQ6jMm9qSnv/oCQRq8HBEYKZQeGJBusHM51FeP7Th2cRESSdJZmUvMisrHqq/hHI66kXbFaCpl1s
LK/dEO/XD1Cmw+Dw9Nbx4DMRMcHEV2nrGEdNaFjAOHnRCf03NRzNI+xj9qb0KzM8myBZx/S6OZQP
0rdWkzdmeQ5JWapprDg50v1w+zmsZHwc0XwfXgIqHIQLiu/E8Aa6B54zPvf5jtndNgBQEgkaXars
1DX/HJrZNQULRZpstyOH9vEWWd0MVhFSTfE2GqANbulYVLErMTE6Vprl010bKS3qx9R0KxQol8Oh
BsRHi3xKnNzpsOXD1hHG/BsE9ldsO6jXarC6TOwt9Cf4zb76AAP+jHrWzdNfgDZjUBdz8oLLvHtT
UXMW1LrbzPDKU0N4ANPPpaN4zcHij6sEMibSaV6xISGxljVMpkhIO/RX99weCNw04GB5E6NfAjYR
Q38OM9fjKktPSXIBdurkZkMA6KLgQBSybCkQZlVsS8/Wbvv/0AkAADkPpOjSXmKI/Ll3qtYq3IJC
437mcrtqt77NNXNXAhKSVdsR6TvLKYVAAVbZ4SHrBJ0hPd/AHFKtw+NH/e2tqcKfyIgN5iMcsJYT
UM2fbpwSnUChU8PoVHM+J0RXoRLXn9/m4QkrjPfdMye8ALJgHbzHb/RB2nImWNr5/TCeQ0kfGMh8
AY2VJTSkhAncrO2ieJod/A/Ca3wijY2c+A6hnwH+TwzZA4zJSUaeBcI6oi6qHSnIlfF4yNiM7M9J
wC/oQjPcV/nVJhun8iXoYpl5FzIl0SZm5pkbzEe0Rw42J1bfbmtcAXIAcCxe1j6ayFc9UOJ3EFGX
q7Im0rIJhci/6+F0BYGe3MGgLyhO0YizIHOPSjjqKVeFKpStaCE6uQSLTHklO8i0ASSLGamLDV5E
pLzinVNBLzya+PXpFsX+La7BtnMEaJ1sQaSXAZSmjFbX+gk9cnS2elyNISZIxnuQ+RMbspzfVD+t
n6JZraCsOYnVtcc4Hwan4Tl2KA27u2MGR7oi/KY4Oo3QftanVMgdYI/kZrtv92GOmWyzDybI6yG9
5zESFA6VnXkI/YBHMh+9at/QsLQOTg5FslpsIDaJTKKn4PyG7yhepRj+0ZsS8NVagY7XE7X/FcNo
dkU5uf3JkTPfV7VN6jv4K9dieNWo6xOMDHiEBmqMM26OT/krWVH5AX38J3bIq+2GOOzIpqrZns1K
DbJdV2fed+0sIZP0wCFWEumScEDLYvvWMOsRlqTV3PgT0umlNd4uORF1N0oRs+OyjTDGDXi6KN8n
cKL0skU1g2OyX/ETLV4FuIGZrf2eXGQYG4cSTod4pMWRw4lXfQAoAqtBovFNVv86ajL/F+ucRmKo
VyJn6VzQNch75I4iYtodO6Umd9wTy9ChLw+AAnevOTq5jm6sQFOsfOQlPn8z1Y0LPS8VopUG6Ysf
Qdp83jwGQ2DjnPuR08H3wLb3clTxL19bEJdIwwWWgtb+pGqazO4WJX/bgyNEWDN+Au/szBt1JNDt
c3BJrqa+tgt3TG5VjESMU7uNRXB8M8HO5uXvKqid9oDZHY8nz7W0k7+mI6b/fhmYGvo6wN1MJqY6
ged9JNOWGWyzh5y2AV8lUs8PVixTCdEPlUdk32Tk3XPwLCLdwc7+UUR4ZiGDzpXcs9JcpQbfJn4y
VoAkUAPg7CK+4a4rBH+uziKWdWYXpuvinXTY9ywoU4Zy9Pqb8wcY9/BQxzohsXfZndvAHSKS4dnH
fvv8B2g7OIyERR2G2Zpmc7FIrvej1iGp+1EndPtiXKRizYWyuwURnEbS9bl6mjqDIym8LB/tVoNF
QE3Mk9SqsS3nqLJTLP2w9BIrriSOEz0N9j9sLxipDVf/CWQ7vAq/yQA9pkaSQZPd+ImeiQGQERcj
HfIVVoRf37nQONDJHWfM/4tfiZfsBcKZ/Mx5g6cVmbmZ4vOViZB8EpLMvrInUqS9sFK78PGt3tEk
HmYETfXqE6W9CCClVFG9wXBCMkp0j8Qpb8N0XCeJRg5XtQ8+TedahflYFAD0fsgylFXZJDVI0KOE
oAXk7p7FUc2Lqsb18PEQgOrYSDeksPSLVsDP0C+B8zxVd2KG2feTTUG9hPKjvmf2RhX2NtV7tOgJ
ZDaDHPFi/53lCf0QxYzE5f5bpxU5CjKEVhOvGD2ikKd7uF1qkSC1reiRxkr8XSWaSh4bXBXB8Re1
55KyLeBIcilrQ5xIjdJcxOVymfLo2jYUO4kbdc8O4RiBadBqVp/FVGoNpaUW9yW3zmr6nEa4tt13
0D6Mz/p2gZXZ4ap+j9QKKZFTN3MeiFqoOUL7GFmrSwAN85kM6elYozH089dEv7rXdvIdDcSE3GwG
R74KTtsrComP8HVeVMX+N2vIHbwLAvMunMr0fx8JDIst79zfCEGPN11oNOYpDisn7tMR1bdPVqPl
Vf7z+fU7mciPmWO+WR2w6nmij/tBsIwG5/q/gVIBqYGjunk9wFFo8CwAIMeShS6rDgK+vzinaNsK
Lf7X+zweBRfaBw9e29wXxBj2LZk9NFXhs9G73J6peBHNGzyqMBKJa8Igf8rlsRFMx8LZLZXHkuW8
fnm2zkg+NUnZP6Hzre/QUAyMxZ3++NpgJ90gZUDW0d43ROnj3XFWLh0tnf9zsT23kWKUPYyq8OO8
oh/Fp/hLzyCERCZQ2cwiQ5O/b6Ug68PGQ/pep+Dt7DH5TGMkYlC1ttJfU8DUfGNUaJcwdNE/gcv7
I9qO683g4og4o5tuLiZCiMOYPS49rWnygkIQs/G9ckt05CPlXRbzQoQvU/Aa4sOHM3BZFY+mR3/R
fgwJG5iNBJc7VvbaLpKIYgeK986nheooFrlMS0/YWunslhI3LPq/Ua56fmDjcrVj3c4tLQKgGMHe
PJlQ4r0a7pzd3fjaWkXU8P1trbG6wYXzbVy+CfKEW3J4FJv5SMqQ3izkvqLlTd4QMqcuNLbGJylC
jw9cdu9R6ULgs/K+G7DjUAxRcTQ5fXFIHeow/Ts1agSQKYWF6Gl1nfK4jApFDNNRMXbIjCZahOMf
4bAfhxEm8ME2Xi4Z4LCa1GgdBAywETK3DP6cU67ddPcpAc2KisEXtyfuN4XFrkxdhjf8EnuYd2Qr
c9UeYDCtat0ZM8XI0r1q0H2pt8MakdUcDX5vF+iKY7OC1v0SR+VfMK+aR7DRkJy9z0Wh1akPBzNu
WlfE3rnLH9r0MvhDgMBQRtEnfGxea0Rtt7FUa/N2JH02x7RsD7EWFcRQMwczxaM5jxBqbFfax0hY
31ZGUPOwdAJwWw09XTjUrsOOK3/u0hd3vzReMHlxSc9MFI/WylsFsnm/BmU5ICwzThu9Clfh6RKa
m2ozC3d4So60euUTprxiKJaQp8zEpUVkXKvpT4NUBqkwKB3EIU0wa7XCn+ppsQITTwXWxiRuPh/9
Zm/ySeQwpXlnj6ABWvqbd8m/0RayL6iQO6dHXV4Sgjv/tY9x1mE+KItERl8j6NKl3Jw9Fw1zNFHH
hcUX4BIXzgbH/Is3G6G66D+TE4gQ0Vt1tYgQkcrOCBY6l0f2JFR9p8vSTM4iTeNyJzq6RQbWqNF7
dfwMPeiqCMZVzlH8cYovus1I8NHwxZEPVZR6cjjwV8IOIIDeceFvSYD1Z9FdY6JNOOXJD2UQyDIe
h6v/r2caXQ4IBQaT6nN431pxZx+NxB+9QoLzeYqyGfhQZzTXGwlB5dzlnoXLzdtce5Mh1yOi/eY2
jZ0ZYsQt6zp/c4eMn1XfBoHCab1qe9K9MRgz5tg6V2l5dSIYJjEBxm0S6B2v70htpFIF/xUJdvKb
t34nroLzKh6BYhamTTf1SZCMmsiKR1s6cpVlVptKafSiKjUGIE6ScyvQQs9YEYseI+qqwLkMfXn+
D6h3/VOpRmtle4tSH/Dv9P12RLUY49C/QS6mVcH+tc4mAYmGzKZV3AuPBGAcLkpLa7WW3HKgewTR
Dc03qPrXvDixPhFz6CdGY1TOAQgm3yEjFP8yReN1GyUvfJrA6yFvx5n+rj/qGK3bwKvo0MfY7QY8
VbLwsU9NKcvSXoYeZG8rcECq+KZaCVpJogIV6rbP92U6UFLZheLeAaws0yEMnwwrWoLhJB0EzIzu
aluNeqIHEaqVBv/9I5cCdeyY5nw4S9u2UE4VDokWQ9fBuc1HxkFzdYr7D9tKQd3cLvz3AQubtX7+
EpJF43rAVZeZym+jDgNCwdkV4O90zKIIu+D1Iu3+ENdjlQVrk8IH7eNfxELIcmZVukma6A4zGOjR
iiOqIXRgC8FUfyD8lVh9wmUaL0i4shJ4KkNOicLgEyBP6a1JXAgB0YzSmerhxYX55efnwKIzQugg
OH67D9JvKFJv+/1oJjAw3riCU0hKykWGA18dO3KgQK+DmZtmwtYxl2Pe49Rccfk6s0nMnuRzggUO
vJ/GqdBz1nTCDBfLEUgVmopQ9Gfq3mnAYkSsT7VSIZ1IVs6/7QNhkkgBLp9XCm88fFRSrBnn0yIX
5UYEFIsNE2bZNdkzeCvAotNJXnAe8KUw1ucTMNkXmFwTRG79p1wqydZ5uA0eAx8bb4piVQn2neBj
jfb4VxGa6WKTni4E1E45QoyqJNvMt662dAZi2eY/DMFRE5W0DuZLP/o49+5HmZfbH/Evj4j4dasy
CQE0B27lN7n7rGD+XPU3nujKN/aoY3oVuW9GOZiKf54x0oVqQqDtSAHGnE0zMzOqxH9mnJHfyatu
Cy8tdxiFDvBgf8+viQ1p2RDqK65PB/rmwHbgA0smKiy7WQ/2KYcSElHywu0T2fo07prjsjAESFFe
nLwbDpwAuPCNqRc7HehApN7RimWgH8TWh+XRALbjMOXiRRKkYntJsVDLATVTikfpgPuuAmtfmWNw
zAt2P4AcxSCvCAf6QEMhXNHGaluvbM3QzFKgdM8JxZ0YdL/7q0n9pJScc5sm7jTrED23UVzWnivz
FzRYeuShx8ivb2S792TdfF7/QPAsfdclDQzB6/d6LlurRkkPVGWRXGedn/RU/hnnLMHhYLdIJGdg
FGTxLwi03+S2B1s7JJqVyAGJIn1b8X2A2sH1+Av65wvLTveAoAM1LxRTCfN70AI5z8HBJVcfVWhr
h3noIYb3rO7skjc8AEwCx98wJAP893UQYfPsLDs21hfhZxdwL4JK0+vVjYZE9N3h/CLcxH2stOT6
wOf/WzI1btNBuDUXI/Bu0E3UvA0Lo93vVOeWn19k2bQXHnqdNArDMrjF9nX1qzORRZWIHf6WG72H
tGyiMBViaLM9YbpbJNLrk2tfRLpa3P2SzlhPEC8EBIQ4oSwxXIhPVDWSfi00QXVi8mEFrbi1riCc
pODdJLkV2voKe6P3SO5qXCQTbHbG/4qEA/CxyKKGiLHLMq0x1IS8gLvTDt1V9ng4st1kP9W7dcvE
NuaYq0Aw1fac4PDo3VNGijtswO905zYNmn0kK0yFyeN6IsaZZDSUPxBUTc5QBbm7IIlPwvgRblWz
q1l6WV+Szbk+wu4Suacok7jaKXTvT/6rP4CSqKcMC0jXLodjUcN5VMdQNqdt+FYqOT6e4/FRq3RX
7pssP8MFgazoWRhCzdFiEskF9wzFEM0TeEArm159KGhaqMUKHLwhYCX1zStWvIAmCKtnzSjNx+s4
1mRE96DOYxvuFIZnAZ3j0o65yEV296xkTHJ+t6PYvvbrMkXi3P2UyHuJdCLa4IruiwtSpnve9lI5
g4CaF5vRG/mG4g+Yhjmw7TNA0JWLh91MlnADwsy30Wm1sKd8a7M0qd25IJnidz+LRcRVUP/K2uoB
lxypLdOfNA4WhgRJfICvcOQLRldaiFIRkg9VprZjzNIClt93+CgYN8l6GAASriw2yc3CfSlv5zTU
Yv6aMEoInq9VpF9HrREsWRdyEAtojiLzVHPo52BvyYIh/8r0A5PV5VwUtGWTX99W/avCZnOl9FZ2
hAc1qqnsT6ygHpZaewROI9JkRmvPC7p7RYSu4vGY3JDWH+ohY4FYj0j6UU7lh3mSE9+GpyFgulsU
q0qS0peuBzzBcdWXILPMYNpf2baVAXHt8Zxw/A/CFGWPbTy9T7m6pSdXJMaYl4UldNfUCWm08LX3
3+ESrJijX619s54XMYxFuQdiqSx5aYcgq0KtRm1oUfYeTF8ROd/tArbqZIc+V8/c4NoQmpQQp7iF
C0Ej6JcTnx2m42bdHAFW9V8Z3V1j3xXLcJgSzVlVFtZHKuMUdRYLKXPk6yq+5J8jZZlVMY2R+8CN
0hu9bJ7ejByHJZOpvxQ01gtXsb0DjTWtXVMvT4VipZq7C2wiOlECTEyhwoaq/BDu48vgiOk+jofK
AVM+ND6HEiWxYAhA63q8WRX9YGFhw27xdZm0MYl5CakPI9RynDNammWEJtTJF45UUQEz75NKXyym
5YL7ih5ZJJWtzC3Kgy5xLiEllzlvHhXvKnI6d7yhqITrSJwSNmIvaRSB+SpVL8AnghYGmx/gwxWX
JYxpYf4cvt4FCYhyNVCjUNLG2T3f9NHTCow6slvJ6X7VHt976EpGy4YOrgXCql4jd6wseeAFjO39
ExTrM8WqKhImMptemUtEWoD5Qnax7ucUGf9wzGERuaX8mQQObliQchUfARLTakK41Nbuk88CSU42
PqWV4cpuLtGbMnU4snqbBQTjYiqIz5ZSPzZLsVooI2hlAuk8w5uge43h/RVqK3F+RusDCBkqA9xF
Sc31h/i1WL5kg2ANdC1dQOKnvHMKj9Vi/vkzHENpdiaEqvA84JeuhV0nXYkww3ujYhEA2slwLqlO
xVyjuZNEbQs6c1wsAR4KmJY+msTvBtmGnlCpfkqM5mob+6UOL+IchnObNOxTAxWGPPoPPqdJRLqM
Q368rUMrdYuiVMf23AiO/gyW9ZkRiRX59H7gIh5QRURjXbhF886tpeTHagrCnRIMF/r0dZcoYomO
ELiXDRGG7iPYHD/ucllOWXdLDiSzU8kt5QKa+GHhZdKDD8FlFl+18dDU3cEmHwT9qqreifZIAdRN
L1iTzvptvMRFfNqsbC//B9q1Jt589tCoT7PRtlgW05qHgL5BqA619d/PAIgOT9IFmQCTs8aZk5i+
ElnVGT3jId3yg+8UJvbGtPFZC/Dcf/RI3l9OMCXF0UQoYI+PffejWYdImlIXpH1Se1spJvdOcj8x
OwCepNPWKVJVOOtmIV629np6wUQpq7ew6fXNc/3W/ob29T/9f4cWMaPgXa+jw1qz6U92R5o/PJd/
JKewRaFYljXhJ8KclBRDrNd3yS/EEc/BpFanR00hx6zxRhbbmhERsDDpc/lIYirVxYA/u+1YYa+U
2+ADZOln6Z2iUJB8jLxPsAtk7qFqD9+VHI4q4vi1DXdyLakHiQvfTlquUvKRenSQsMWA7G3meq0W
WkDMNkGx6pyf5WvZdFij46xA5YwyHKt0vAb+xYE95pz5Qu5Yy/kDfhyYVKQDnDo5n3ZE86OXj27R
kgwEV7qbtLlzHAMDLPWvGuPapV+pqAOcK2vDOK0O8HQpLBblq6QsWV3GuSSQzxDHzznmxu8UYZk6
+HtwdNjnrlyCocpkWlkRkBJSggS/e/aO4ly6V+11jsDVBlpDmgeZP05PwJINRHiidvMTcYqIcn5c
wMFUkf167I9j8WPcQ976NRRW5zxp1srpyvGWwUaHqtohdAgRo0y54UeXTB53jzoQPGjhJ9cg/ZT9
lzoNgM24qSVw3aQmelQS6fP+50ZFKMHQ5HV8NZ4edb0oIzp8W0st+Vcyfp6SlYM9FhMENNmV6m5m
jG7eLrhzf2iKoN3vlmFVKrAaWgJmM/OAdcqE/h01khUyevZTCxSLzJoA4h/HnfkGzV9RZPf/PINZ
dQwGw69VHyUm416sW3bKKb/G6fDFZms5Qp2RmntkwfUFmOISLRTHQrdkuBkMqsq3rpPbTiodRDX5
PPHIG01coXFKWZ+wVr8tSqCCZE3lv8U0lga8Eg/oBbymj46qSLHyst3AEzyTxbs8Cf9R382P0DAR
zb8g0Y4oL7dH6Q7KAy9yCct9QJ3MWsdEYEANeVYO8fQnFD6WNJ+ZXLoF8ogCEKt71AjfPZ66L4V2
6g+TArHD9RbUuI7I2AsL8CSEqBDFJDFSD/ezoAtJjf2XDdcjwqYcjAAxjc/8fX39l76ySkwZEHcL
iROcQ0hepUWmAazWVq3Fny/5qecS7t5tdTvJkYJnqTVuA3qFPE/LgplDpS9vidXtA2bzq9An0xD3
qpbrrCw9OwAZFinOsgCGh+HBqLXUrLaRjFEZtap9FHEiuYUM28+iycPsCDSp7Ruil8Ox/R9zlHJ+
9NbFnPCEFgOSJ0LxKpdQnPy7zjkJFDiuFXgkjYJrB1nu5nQZTlFrwBqMR/vB77C6TrHisJtJK0qX
8goMgi0yO4QmdVcl2lxHgSHZLdIs3Gf0TEZFoBFkW+Tyvh6stwdk9gH2BAD8/pp1lR9bPhM7rQUa
o6ZUrDKSvufQTh2+/OsonTc42oOBDecgkDA7GEA4KoeGz4MfVeU/szTziOq4o7nLawjKeSUJyy6y
Ty5k01cd0ntRcuj+dE2CtRfn05MKzc+pqTpHMVPncFJFRrctPCeemabRo+evFQVV4n/oWCoInrH1
IWP5B3KmyjiRTW2Xd54JBHReoD24JV+ijtgX4EJnlw5MnNoVJifl2A38Jt++ECwwF5nYHiPFrjxn
a8qPhFkybE2uhPFjft0UXXbQlejjbk1LCDLFejb6MyYbu6hWRaRZ2zvw0I6/259Lxv+jWu4Clnoz
gRczhCmlZeeX3J1nsbQF60uva4Lu/f97b7eGDZb3nXzTs1Sd79CYAO0iGJUsXbe4n8P1ABKbEn/S
dDIb/OiQst2uvGIQIs/2fgIzXJPI2uOctUTXCZYOp2DSayTSJXwMHuwomvxNua4rmzNBnhONeEq8
ViISYuopEF4u8gIa1e297YiSQaYFpu/Yd85slbNIgbKrMVbiDKRA6rBiAceGthw2NJbssQYfmuOK
sAruRxiKgWA8b76j8fwFmIEWqY5d+imO5b+1h1V/HWwPQH2367YlrhBkHb4TRdiOCoMbetztXZ4r
NSnfUgJfuBmfPdI995J7+M+zU9ghlnjEMD4Uh4ipPS7yFAki12JWygd1QLmPMUbsribSO1WUdZc1
euuH8DGTc5+3l1JVQw3IWO6ndyr+T/Nn6xcufJO6vJHNPUZZQYY8vv/bl0GfIYviXDB5JwyF2nVO
a3nk7yA0JcDh+E/TU5HcyzyPNhL76lnOpW83r+8KB6p8VRimIG8Xwi1Zw4W4wz65km8ylCxT8RUz
kHBpl0/VVml/t0uqUgSUNnIdT+ENz+mR9fKy/P4PnB8kEsmwRNmqzXcMOie8t79CJoArn+HHNV8B
q+FAzbamU2Le95pfIV/TSjVIpjeSCHFJ+uYdhksvsh8GCNu3A5Bxt+ki6gPsVZjO+oIuMeTl4KEQ
Hbhstcvod3GUkRbANrmKUyPgAPXDL6eN+naDRJqPLqwiXgfNZUGuZOSKLvH+GB1Tdy9Wysdu04fd
HNPEHVVsbBT2eqFoqHtbNMGK7s6Uf/WBzhUDjcSWV1fjGFlVsnA/BlclkwI5mwoPMFzMbybHcEb5
WupDimC4jzla3MhXc9DMycozJL/OX9gN7sMgJl2vn9NRLysEJ6StcTbTHFWm5SEG7YINNV/cP90o
LjJ+3Z4396icuDD8uHrEYH4GE6gKJpRYslIuGa1nx2gSzMhL3Lk/iy6dL7tUs+z0bBD8QI3VTAS4
FdkV1Hk/CvJqmuoQYAArpYjSVo+8zBQBiaDcVsO1rnNu8nnSHgiS3ie0OHWQl9DxiGPVea9zvAF/
pHljx1iVks0160VuxeRlg4YIV04ybvFKmXzuNnJFNGelZUunnGv+2WrvuDi9+UStQcPl8TG2PE8D
xQBvSKBIjj9704LrxGxBpzqyEN+p3b556siSzX1zyIhycKjwkWjc7D3RDb5rimJuWdLgNGL26yrQ
yEEbz9urpuiR16ixW+QzQnQ0rQ+umnABYG0DSPx7vV7TBzLSYvc/g95bAijX+nSG7Za7Wu46SMO4
7OKtX0qLq18W6Ps7XAzWZtBeNiIahSE7wO2M2vGd4kkFMIYpy7U6lMsL/xkLYsyO7byBVX7TTzuv
2GFu4xiDoe3L0vdQYy64PYZY+j/1fiAOB4G4PAMiMoDFlv7PL4U1MsbWkCqXuD3qpz+/6BAAc2AT
ZWVfI6hBBaMj8MDmH35/a3krlhn+DpqyxN7xW3XhBPxtrZTXB4ZUtUtObkMLIk0xOQG2RXTjuMue
0EPiaas6AvhzifCpsgkFhSL/qq8+s1B8gaaFR73noNsI4ESaDMUR963IugPxRm/k6MGaYk9Dkq+x
9Qhb6fqziRscTiB/j3wQ1kbW+4s1O2/AbRChynJvy3VYXoCETmo/4z6P/766AXT6p7I6UomghkKC
oXBl2R6TMI3RGNNqTJ1OxHhUu6bNNlMCl+5KwHYhIPv5zuqf6nXm+kIQ8C6rRdz1GTDoK7OCDQsx
yB3HFfb6sKCh6YB3CI3gCC9/p/wuClhTW19LmlLDFcsKdBpk6UWJlA6dwdU4unYT5WQZqNxn1Z/R
uWYfgTdu4EMWMp1R79CkEK/hgQcC1FA93nbojX8S8cbHAuFsE2aXPMyVwT4bo5pCoP+7JAlmo4wi
Vk4rfG4+A1RWknwZIuFHih61ofxlosdnJ6XmiMfpcByYSwWR9fh05wvLKGricEwFrySihbtemfzX
8IIpMqdUXIEuHm193OrU4IdZiMj0/ULB1Z4+3R/4jGhBHg9+wMCc9jE8VLdsTJZ7okK26nU4DEm5
nBvb+IIMrsGJEvtp4IKBP0tGO1rJV8IDZ5Du2Dpntk8XvIcMXjPUDsLPOs9JHjcJb57/kv7bMtvX
S3YtZuvtQg5AoJtXEKrhSj2DZhUWYirLnKGi/gAMnuIXcvoSgnxpO6eDnOxzQbfNrkfX7nPZKIE9
MN452NGk9gTgRewJX+JHZ+W84Q5gfdSsE5GFYpS13pJQd+ofhOwznX0UWuLIhIAG4iKMbfNLYn/3
HJfaVYtyeUrH/YrRpKYaoSeLWHFPQ4ZMxyfFm2SeKMZ1x54lcmZPV5uAMIwRi34tOMBpylvvW0P3
R2BmXStDvvVWvzz0V9lecqZ65NcSFcabbJIXsyvIwCPyCTzgPJS0q29xDjQZwc4MJaxR+TypTHdg
96yesMqZo+vV3i/hD5i39jw2geT8pebjdlHExtwRRUrIN9wYQ72oiJutxi/3sV7DkFDn1qYb4xk/
/4ENk81VxthnrveSBB5AOeI0UnR/DyokNx1FLCGGaeseoa5UG06e8/4PC9JkzkL/0ofUrcYHztb+
O4oyEUxEpk2E084JxXJv12khluHYg00MCia8UP6+tnZ3SKmOKuo8EASy2fK66JktI4S+On4q6FIv
RioessjYlYbfWjYNN7HUpkft3c31/owW2u91+K4li5W/9lAOfgjQJyzckar3fZweNGrj/+B/a7B2
7UI46tLsefq1SVf6l0IJT3vp5HPzncn8XtpczquB7txpLX7VLWG/aGhLwgYdGha47w7fdfW/SmIJ
e2/qE0BcfD7n92TmxcgcXkIIW9q2A9ReLFCpSAzIzr0ShP7lc+uJbHVHnXbDL8U8do6Hy5nP/HL7
/z8oxObSFqwFYkswqJeYcP+UgQAJRI2CDRgBAqqbOGBxvFCKhPM2XoGr3706NpQmZTh2bYbcHYk9
Lx83gvc4wmssMKao32nHZFsh67LJxj/mYHVF/anPNBZfq4ivjdj/m7KW4PWx7nuI0pdywiRS6nvb
xG2wisuRKmp0Xt8W3lDahQlXiwZVFo7YFC3rn6TRkM2edVqf6wX+qkX0fzvbSJU+urOZ67/PkxeJ
zSnVy1ac3600/CkBFI9tipKWs94FcZX4niBST8bAXmiD9E0JfwKa1Ubzs/6vrKqJ85LZk4R6R1Or
R30g9XLFoMK2zOMUO8ogvFBmmf0T1JnQuon9ZXWHhLdAD4UVAIJHeJX06zFUx8Ez5FN5JT9po0jH
Ea877D0B58XSHJSR1KMoXIEPigZxlRS+ZepLGLFyQmrulazpwcaOilmJ+UsMmRb/KjgowRQOEocI
CxgEaALBYOCdw5W0nF6Lytbn1272RNupXApupG2Zg12OEc8ClWBtJt700k4OQVHTxJx96s2Etm7a
pAck4krHIoiYQoau/Ro1iSXSQkK/p/UXHw2t+h7swjNOcNJo2YHtKPjOEMESitotaFLcV40zdtMt
Ff5jegpHs+Ub1sE3zbWTxkz7k4WsFoDUZmnqEk9OirStmBUo7Vv1gGRLrkQEDRRXpd78G0bbCNlM
Yt7TpEFQ8ktjqL2jf+QF83JdiZ751m/eJjzBvG5jMa0jW6+rLxBsu++61cWNsrGq0H2XosqXmqU+
pLaMbuIAEQGhhAKrVAM9DGbwst5+DFlabij5DHWsIElMn3w5Ie+eKf11fJGYKpysJJ7OCLkdaIeA
O/PV+JVyYP1WHGynfpmIRlWCHer6jiaJ1WMK6Fvs0n7ljSIxRPFeRwXsZzruLy+qrjsw2Uo4ZsY0
2quo4v75Ee1SD0GML8opNBPkJSE+6Dx8CGbYzW4gAwkDypKk3VbiYOxwixsfYHf5GBWlkGIe1csf
+8na211B5VgG7/OlcavNIlafufcNlmlZMcfec1uzMlOinj3jSnyRKOIhqhRgw05gf5S7Xjg+wtOt
3FNfTFVv2Inb6+5gs9A+Vd5nj6B1bbBcCWka6AEWm4gs80dJxx7GsDfyRdgN19KuzJjKCnVzRgrf
BxZzSWm5lIoAUlJ8Bl6/cPxjMwyUt73iryeXP/VaGEchrd/267FI++WLH9nqsDlVWfLGruzyw7Kh
eSauU9ZhhcKrclOuJvGa/oSuDhImERz2f/Ytl4nPXg4Q14nhHet9nxiaUJwa4EltKjyqIsVEjtK0
K7Ki5vp0O4RXHDkxa67cqlX8D4GMq/cjdAFw+5V/WWJrpyL7Fdw7Tpg7VRH6GluuYLRAN0ObuklC
mVNhd0yA+uZVpARLQrojYpLNBslEsqY2XdfZLxyV6EUC0A48RPTUqZuXXkCHmogxFW9+uawfL5aW
HYdiTJ3eY+bB5KnyrtCMTlSlSDBEkaDvSxXU3OgHjoXj0L9LuwL2S39h0U40F3mnYZM+ZKsSovhN
n+78P8KSzkRMm7bdW8P5mkNKxbx+K2nvw8Hfq91GzoNipqwl6fVn+THt2HgJpVKfW67nzEjrUGS7
nATmwKRILDkx/BKDHZzRyO5na0BpU4+0VISe7RjsHE0NP4rlfXMH2nzn0PjlycVJYCn4OAtXRaBS
FXNJgbOO3iESmquzgsB2BIiniNkUtjf6jhTxKV8g1O6jkZPJJfhLXACFods1RX/V5Z0GUAnIyhvV
U7W/ixZOadbYY5IxmkUPnqkUzk3O6eYtTgiFAEBFd24arR1zlGeZ8mWi8QwBW0fy9HQHJ0I8wCut
J2thzqPYJjAGw1LsL3Ug+RbvvkfFHfvJPuN004Bif1Uj2OEW0V4aEZuQ8LW4hBda73+7WKXvENRB
2rLYEzkdkXz4BZoGqkvXBP91yeHWRspjxnmN3z1/OADlERJ/yllVs6sUtu/YqXPkyZE42gpTM6SK
XkWjqbZjtjcPBmqMO45cpGxX17wNutAJu5e9kJDWyZEixxbFfJfEI/Tg67LMLu63mMWfCLvc8Bdk
4/ib6BrxJJ72zcXm825VXr2qL/8SU7yB/UjjcGov3YGakykywSteRdswUREiWekPB1RLbKbR9uu5
UpLqUia1DDe/HLkZCrGq7IRMml4hpNSUPkfL62fxpxropYgZFT/oG6ap/gGd+ROAJs6djntAxWjz
MvjVj0Iji1obHFG+8oSKj1NQ40AwGmP2IeuUk4Y82OgF4P7c2vNP7UdTrluXZGEwX26rMtPrMaat
RNJE/QCf1ViaXm6OvhZnGDnHjHp2TenLz3i3cIlQZB7YvP8sw4VqtKwX/8e2+bb01T1z1R8M+1y2
8laDA50EzxQ+pnuPjdhylkNkgCwvNYI2XD00QhNMgPmWH15GPPgwI6wnZnQNwJLdj6CuVEdKJIxn
cO14p9EYCTvpnHzZNXQhV6MLuc6ivVBVQ5ycPKjzlGu1N0HaN0fJbGhdV5F8g1K+Xh1Z6J7Aqivq
5lnB/jmPCBHE6NZGSh5K5vH2emFLnDO1KsqCUlWyGDmTVmj8DR9H8HQxQB4Wdd3ICpB5XNHxfvvn
quunq4zhA68GTjl5NLSXVmYDZn4ixfXbZDhudhrYGnA2woegyaR1JjA/qVrMwLDdufuUK4LfznP3
jwLtgbq1pXQVWaGCsTVE3UmzMgoWrgrCR3XcVZ5PSw847J+AMeXjFIOOdDSCoSdbPC9qfPl5bmi7
eStdLCFPssT6rBGG5lIN2kDe0xQAZjToprIRnKScHIifAttpQHnPxaS29M8l+cH61qe+gVwYBLvb
I9EsBTMouNduMp2WIc9yjCX6hBB23FnRFDlVYyjqeuoENjQA65Vn/XkNbQbYDSiK0Ej3aMciQCc2
z/RDbQRUgrLqyg6U5iXD6WDdlMgbxmOaduPZHByELq7nljLfjD6zM4VVqPLTOomL9aaVLkwSsgEN
ymMR/+N/SWi+CxITIKXPxmIHtmG2R1EKus6bPn+/mK43ycLNCbKIntLuf7T8bQMQMGtQqqDj6IMH
5dEK9prwpQvC51h7kXkKr0q6EsZFzvdpkg97ZVdT6Fdi/v2HP4RZ8bmjgsG+pvWK6m8dB+GtPKtP
1t1OiZYN6r2l5VGhMtrukvIgjsVvFfmvrDcRcRonzNYnO601bdGeUcKHf6Um8Nu1YHBK05E8QV0F
ZIAC4BCV0yoAYApE7L4Vg8K/CXk5Okh1Ulkes5KfD8WoM+tUqNqnQ+bcXE7nk+mK+/Tl7GjO9cK2
Nt/ezt3R7Fxu7GVuu6C8yo834oeJchQsSBJRBtOibhm7anwJ4MvDqcahMnI0cZ3QmozfHiVhmMdb
XAZN5o6KkMjridYGAtnVz9KqfhT1k1sJ/Ao13MHOu1BLAh/2QbVxbbjdAz3rMJOp4dVx1FXxnVjP
RNvZn6IkAKfSLLnn6Q3G6W5uVJphS9Q7GP9vRkU3zRTqdCOqhy9+zQRMvybYRJVN7h+lqiAjtxAD
xPPd1GrBEZ3v+wlI6y6YHqImkTTKofuxTovEuI7dTNyjkAUvrIdM9TShwbOEhBcY9QFDhQqygcQ2
5N7Dl4TIgB0BNW35GaOVQn+y54aAYJYmJU9KuE9Ke2o17wDfzUPZsNPJI2qbAyrDmv2K+2AkIqyu
anRBuIWfeqc6XFhbTWiRYF9rq9e/oGy8VKjTq2of7y02ZXeUnEvY5bfxMZDd2ALaR7+XglM4T8Pm
hWno3e0t0NkGVaFVteQQHbuNSQR2pl7sJjtRWE+07iBRzMO9DKt9CV2d61JPVQ4rjZwBnSbrEouC
9sZKAoDWc6QVqYQ1m4OUVIbz4/P2jDnW+tt/zzwU8K/HcSNImfA3AjTOm3Yf2u6cDh2NpU9Z6qbH
4uav+YwL9cP8QFT3OtOahojw9u8pjxLoL+aWROULT/6ezs1ZaEH9Z+3sR8GmVMKfEJ20cA/LdPeb
fkfj4FrUaRxlObpK6OfdfC9YJPVw7DOexnulpfMDeeVRBs6Ars9qZ1o/1ezTKWNkDodc3ZaBHMqd
SAuSZiThGNdZg00A5cMDJI5jZ/uzEWjIvDlNGsLvYJodZaM66mUT40oKnvLSPybsPMGiJUDAAbrB
5Iht28SEYDwKs+qneT+bsTct5yVp4hqhjYi7B387Te9zUpsEXmGwDuikxZRDstpwEE3I/OJ8iu+2
62/HcIGJKH1jwYUmAusCOjqBWxOEMil98Flpx2mn6hJL2bwBALvHPvKPDxmlOqMnpaROo0aYmxHc
nljQp/shLsKi8hAelpKLF7JCj963/6ueFdEZPYANCxwV2W4Y0JXUnHQkwCSVfhngE3IkP8Ff0IXs
5jL0FBaGZ0u5Zgeu/fDD4XGClsGz0cwxgDTZhktM8FECu6bsVcBDiWPwdu32SR5A6krf+z8xrdpo
cKiyfdKGhQnVL24umlNP1+wflt6TYw4UjDVBKV0ARoB7aKGykJza7Hn2LR6MjMIE3QIsYGQ4uuya
ZznN5NIKgPyeMondbtwMOYhxbiHXWzcPf9bSsT+GH2KBhGl0vpni70AMTHSR1sE/h54XqyOMvMIN
TgB0QM9HIUIaODvK2jW5ej5J/Ir/AccSDwCsApUsVzM9liY6/bM/ZhoZkt7WD4SKw3b8fcclYZYS
c8oJdE693jCN4i0/KnAek05hKVYBkSJiPJhqkLWoKfh9ohlat7Qz9+CnsZlYoCdyUJkNCx0TEV0E
j9JK1V4EFzjn/B7++RjrBS3TPAboXljiVdWMMnXRWRvXtJhR+YlodY20w7RkJBDxRzfpr/lTLLg6
NDlGwyAGzy1gCGdACvUexUERJwHbEfXZtGoBxFQdReldgioZYeGpZwgioFG2Rgml3zh+pOu+WzEP
ESURT+Cdz5P/Xi8aNaZ9Lu4vnmrDFcQfGntuhHs9sFLY9PP4FnkryNTUMpi+TSzq7uzHV/OShLZK
nxyXm9Ohmo2N9/MVSMdsGkWYmWsBJg/1n1HBr0QKthpGfQZwrRjgiZndrjK9oA46RPlB4u0nEJqB
xk7Rna8B68o0S6eMOgiu4+d2hzXSOftFmNMqYmWu9wpl+edmUV/Tv6wnvBTgGzgFK2vyLYD9ug7g
ScZD5oCZrbfuBDQBmnNNFCvnWHZ3xs4EofXUfB4DoaXBqtfrHLZSPfGc9J9ClelzqffaJDqi2jOu
TR/UGy4MN2gu7kFwhSTLuIbTrAr7835JCL8mN0Zr2/h1rCUdd9Mu41UC8GEh33YdquTewrd5uqlR
wNQlsgOpLU65/nwQhKeN0t8YkDZJfD1sg2UitD0QI4IT/OyNHorP6dGyGq+VpZ4l82yrIFFBO556
ccn77Ox0tkvU6NBAwoAdkH/Zp3CTzxPStZHYxXRvTMKVr5FlVgKZjUnvIlU6wRGVmfpq2l6p2it/
jlqNC2T4wT48jZIDHx5aMKSxCDL6vc2BRgE+JnhN+dgdiHez/gas5red0V5MTcww4eTs1gP8KjG5
dplm12mDyHfM+awEBoFI4Ix+TYo19sauU1AInA8xL1kdsE0+SZ9wSYbDdj5iDjDDbLfG72BrO0SF
seSrMtbDa8QBl/UOwkEsnW3Da326aCCxl7BLQcfVDO/d7NOyGLteG6Q=
`protect end_protected

