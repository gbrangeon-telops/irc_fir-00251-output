

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Syf21YU5JnKptD7LOLtaHZM+q1VIhUFTxsmS2r0ofwQ3ushsF40KxXOCQsGAnXjGfc9kVb3Bn0ME
1qO92hlu9w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dY69aEX8OSz52Pib+7B1y1Wvr7162ZPVuHYqEcMQ/oCfJJrpwF+oy+zQI55NVyz5aWKsTxE6uM7J
HbTWuphJFeGo7mzwyRD7dy/8IFTp8OHV9aN/fKWepd3R1nKJ/+bdmSsliOOw+inM7pfx0a3YODTn
FRAbVAMQuwe+OVuT0dQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q+4W/1zvXVAi9QMds0GLwNMATdnR+yvz4Aqge4tYro137XvQ9NhFGdF/mXOn40o0ijOuTLANSGZq
Y1fe5IvAhv/BzIqGLvvBSGadUyLWCe23JTco14xHGh+EcGpkQzSMsD+MtFlsKB5Lh4Pk7Fki+zjY
CYS3IH1yrExDySGaxaJ/xIpVmbcDUIB29ts6Ape06rDNuWSEZkqi5ATlUPCMrVpXs0LgVRBipzor
Mr/lCisQJrroeVDmbpQGOxCT0USTTIePtqKzCRURmGOM39JzikVR3QvCxX3V9zs6LEiHJnsAr/WX
JYHo8e0tsbF+S86/2TJe/j8LJK3VvghHADCdOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jFetHSEk8pl36rsszcvK1lxgvI24/D3eeWIqqx4SgMWK5zMch2RGKDJVjZdo+SXrQZtG4vIfoNJ/
M9NL/crW7IJ+pa4Cb2wH+GD2pA66Yo3aRE1Ld7EknU3x42o8aAXlhcPIjcxq9tmSO5RxnhMKlfjh
dMPsoD+Mezyol/EwGPo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Jgq62sziWqkTYcR9/y/ZRFUy8fWL8zR/UZTwiK9JRpmOKe++dsuUuVffmjjAGJoOkGM1fnXZqKj9
LDnUvlqAYGJAQrwT7QRdCNBN9eBMyr6WJUCOkpNRo5aWbRqVpwZihLgqtvesSbzoaKe4eDRdiEe1
xKR9vPyfNmAnPN1pwf+2YDUftVl5x4CmlqRUCO2c3iETzT+xwYzxqYKolk4Qa8DTTYe9PvjYqn2/
dj/jpAwnTcOKUqpa/3FaAU1zgLKWphnnTU+MOfKNP/ow3ZLVrmyiraKTGZlBmdJF18AzYgHb4rrc
8Z8DuRLa762hnT0qbzjf0vtKn06WBHgWqansQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19248)
`protect data_block
ZMsUcL5Wjsd3Vd6VWmbpcfYy9X0zDWdHHDcsyrAVIfwZeCLASr07+1W4y2xzyvNiqxJLUTnUOZ1N
SHPREH8PFwlbr3SOWqgnzGmVjr+Yg3N2A+uX9W0tqt1ZgEuhmvNrJQulR3WMZu7bXtZxLj7SeuBo
0ur32mgE5l4oaZRnB0RKrbHm2UbYB2rgfEMZjxXQme2aePq2UlXtr0Iligkiyg/ST57z6O5M8Fm3
iLxRlKOY/ekbK4Oeg80sRqOV49JDI53dww8Vqdt9Ku/g5gs2zsvaKGJC5r2kn21GHt1FTZx7PMB3
M8YCdXfWqb+fEAiqLHsbKiD5xyEQ5YA0i78Ibw8F6pS7+ojsA6abCxprG61HXWaEuqiilTrOVnun
ryRNolYurJBir5JTq5A0sTXpv1X6a77deGQ2C7WPMwky+WPLIKL63nuG3O6vgj31BQEFpVOq0dyk
Xg4red82MU1a5QISFcrvffmBWJyfgyu/VxYyxglt9q6L0toy8HVHgWsOpypb4A8Du41QrG+4TC8T
tt54MA2iLSTdrO9yXzlvvoipsNd3O4QdhUq+uRskQZMClS63bqJw6qSZM/Rlogd+4IdgryxXXr8b
AoOBtsafFy1TzUV0tjw9xXtJ+bb4h2X1tL5NuetQjix3zY+Rf9GpI27j1HybwN34bVnNCDYyhwKY
CbQgM4VNIyiIPBLPuXvt+DiwbednQYSWfDQobjzTNCxlO8x3LcIjvy/Z3uysESjVRne2ERi+Nx2v
CAJWFYBV+/vwuXccrLj1cb18VofS4bK21UkLZs56D3Q4/QDjAJDf5jLCMCnV7/XZzSBq17jtf7Rh
WurLF0fD2xccpv3wuW14XqgWOGSCDkFeSWJE3AbnQu68EZesOALIDj29W2e5PX8lGmOWxRBx+yPp
QVqpim13TmLQgGW4Num8F41+K0gAfao2zF1kUanDQmYbFdD7a9sVFm/OLJ1LT9+D11CyyEo14aRT
8T66xq4XStldQLl324NnVfKTT9ri7veH2LYvk8/AOIfKbFQ2WeREabXWgX0FkzFA5K9kQV49kA8A
X4zDqqwhq5WDB151GkgdT15qCAjsndeVVk1iB3z870Bs46uH0RlpJCHbIZ4MjbiQnKCZjx4xwsmE
BXiXTO+9YHF5Cpqm1CsS2AGBj0SfOU4xD+GC6Y4z6z3Uv9HyBII5bcAWDE1QSpNun7uka0uChuYo
7N7U1D7H0+I3Iw1L8apxiHGEn7+wrfzAwPPd9ivJcooap7mNrXTSxj+REXnbggV3cMaqLvY6Y2LA
NrNddErJUS12dDJ55YYWMn/t0eL5mBB6YKvhKWxwTzC+OZx6QGPvLW+JYKNIFbnRF/tNovfdf3w+
fAeJs3wiZr4qsty9ofn969B1v2MN21gsa46ZohyF0jhAcAT9p1RlmUQyvS5WPWJC4OFbMqdGI/NR
mQNwCIbC1pEiE3wE5BL2NZEtwYy3IflZnCI7QfyoRlpy0WXT5AUAUUAjhhMlMz16dk9M0FRGt5rx
TN0UEYLZ1gl9rpfZkAO27EDIwVeZ+v2NQ+ock6WX70q43tfCOnTFBRSBylTavUaT6jNOyYvWrWId
gO2DTL7PCx8aZeWMXJY52gQq43A4ePT9LlAjuTqgcWaEBl1f06hnk+J//isIK3jZPJD9JB6X3MS+
uQpMGDDmTx64QDflB2d3RpFsZzSCnqJ72InFyzSD+n3Llw2ZOSKjNI744EkAvDgIf6xjIuT8pUWS
DehrYGqUrRBcLIZQ/hrlJbXY7rnlECRp4UCezy/+ON5rVx5EnfpX97jxESnVfA3Vbbcvfdj1Rp+b
PDQIPNdOitVyewcissoMRHH/iDc4H00YtNMeCY6NFR1/X/ub/W6blgqChAnKMyJhhe9Lwniv0Qxm
/HShR/tquCZONe7IwuqiE4KjNJSwXM9+16PHKNjcD6CCoNprOUg4ejfYphdiqwoNQEA4xH5z8I9g
MALOhHLicGCeDQOFpUnIfKNRrgKtfzxd8RdSeuqvzaVSlxWD8lVc3t0m9Wsppj+bbTwnj9CSxL4v
vV7ViAokvdjNgMoHNPbRtEaH6VT1dfhkPy03bm/YiLmlBlr6CBJzRa8zki/mXzJOcmi0tOM38gVB
y3HfX8ioF02Zrwmp0800ygrulrak9ZmFhaaB/ynbZOGgroYzz1/IWqaM3lPWWkzSdMJ6pvpD61Pk
ygKJk+0wkUNwWe6qjqMBhuUOGpqsngPwE//0TwXoMr3y8bGKksbR4NEHOe3d0jEWeqxPP41/C2cw
jiC2BvoBA4qTiFWQm3ARNbTTm9va3/gKgx7xg2lydtDXD4mV3lYHncfv3ii392Bp39DYMBCHhfjW
8Z+0Nh4PzEOmJUjt/Sgkk0E1fn1yODZomHMhpF/08T8EK08M7bGV43lUg4NiCQH/c1IakXxZDne1
vMyYJQmltw3QMQGNqvmru+YwHfOJUOXP/33ZRC6vW6u768UfQ4XVEmjELBeQOnuimxiJI6HkWbGf
1ybSLfiwKC65RJH86N52rqWy4tmPDlnsO9TnqymshxHL8a4eE0887oX2XQ4dxxphucnyd3L/Bcoc
oqVQrgPLGP+jpakoeZM65wXIjYxoLgBpkueNBLzlQQyu8H09o8921Goj3QljHvyjyCnpF/ZuxkRN
JolwTQXvw/2pXBvbkwFmu6B3kF5ezwGbrU03AewtgKx5kMOZ1QmjByaWtfa3O2IqF9pAkGlHOYR0
JjUcKdQEQ9XtsIcD6dVDpFjFjeJO0TaQ75JCtdg+fGhvgYerBHEO/9yAZZAxpV/JvIp7qWcnU8Bu
4H6HfQIBjr+fEeAR/MF41kb1x50jR5GKef37uDFfRpf1eKK940aqLfwLYcv9JsmbhFhRW0SzMyfU
OmJ6rSCMNA1TKE3zlMMiT1E2fAfVg0PHEkaHUeRo0YsE6+3TgeGenyORGRYSll7Z0VdZ8O5T711F
uGlo5nmvMGqfPUoszoswkgGwDXA1AGXN09ImSvi2LF6w+N0To255jY1OEJlHHQlox4NqmGNML1bD
Eu9fYX2KIMqtz9SZgBnIoYyY3V7H1GGPFsQAzwjLhByRAvA7kMMVnVUF1qI2/NqmjbQ0MqZ2auPO
J7DF/OYTBipPqOYHxYHOaodTicA156TvIKOkp0EnUHec2dco68vkT2qK7un8EHhJe8wBOye5JnkA
mzwIsY95MM/kezckyEP3iryN4vGt7KvKR1E4dXv44xNfbjrtXnwalFzVlzi4phV2PFLcud4DgOvD
L0t500s+rE9cBVk6vLHihBam4suCZlE5pN8tgYqPb/rxy/xJYLJ5AsrJVYrrMNatCcGQyaHAFe4p
ewgKPEhO1DFV+WT491J42Qe8OanSzBfJ6jrADBtiWuE9Zq4pq0PIoUcuwEQnD5QTK1vdla4HuLgh
eJqa9QS3Xlb9m18MyGC+RSGguB5ODo9VxlXv2AJ5UIT2vftGI9IUfHzJlr7kytfJhxEJgRmb3tix
bReNXVnK0IfHNUxgO2BYw9Jmkdg3I3q9OE2F32awsjX8qC9riWbfmqrvhct1XhTVxNKAoRujGVdu
Ngo3NHmw9Jxw9fuqjSnnjNMuhyZWQXru1TGOS6+8Ny3YGhVcUl6K/WDI/46+dqIEOj+diiYFPl8P
JLF1BiRLzjA2NvQzAi9rW430VwxAQGYBXXmxLGnedH4Y8uom1mlf55/30YaVks/TCQ7x+Mmoc2B6
zln5D6H8tIGPa2HkUBgp9fXAK+uePHQbYBilf356iV7Aid4cJLKsMQMOnJmPXZLgW/f7SchdQRle
FFFSQF90kmUfZhBOeNc5v7bjGFgM5XbI4RQtX2S31hZWnsQla+UeGF+7gvcczrpSlWWyaFOBw0i2
VChvNMTwMSM07idZSjnlD55Y++t8g/exxQqlEoatZNsqYo3D9cutGicd9j21n9RNZK9xTlMy2w4H
lK+m2luHnTy8eOGJTHKzOtolvIAxjJQPocSqyg/SagYdzsMVxgCIa8JP+IPurGGt6urdukJOSkQy
p/jnNjvAABSdSEI79SGyNK2GcOkEXT3BFegz0wQ00yCSVXMLwOnWNXvwymZzwj4RUKtOaOi+xKvw
kHrszevVPRvtYF257VFM9lOSbMJDP5p5/r6f9//UBdNV4yGWsvX/k2pVFb9AmezlGwZtJU5xs6OZ
NfJronXmCSrjqWqwUs6m5m7OMDU9GeZXMy0ak3PqFxQR16UdLUKFQPjxm2qa00xA1bahKLJn40Sd
0GgYr76tgxGZT0J4K8yr4IIE5AETAH+nGUQXMsVmlkwFtGruFhgShT7XrkVkDwbNj/7qvvUs+W1v
IOGIY4hjw0LhriC8Dg4pFnvLiHoUmYD6jGPQjAmiojdDPdZjbwZcNoMY63yhKPUAgAZsX9EQDwF5
5A2fP4WlSinGB5oET5rQjEnJjU1di7IFL4sWPg/6ylI/bOf5gciSPpsgAH7mrulaYI2feKIa5vAe
6ufVCT16MZJUstA0ki4J/StJBsBuuhJbx1IWmZHrHzY0BKabcE1k3Kjn5bpDUa+R5v945H+DxStq
b4YreNAu1MTmF4enpvmjMRk4W1wL/9ljZauS2U4SQLhvkF4ObgrO83KOZue/Ul5+iucnHbRlb8PF
m0TlNpmVK8M6BZMtE2F9ZIv16he6ix1r2h9cQHWK4A/Y6TsNnFgu3DnMFHed3fFWj6PZvpH/DDvZ
HEoDdn3aRphl4xMnoMH3503mpWqm2wokpS3VciXR3VaIn9DIqa1LRlcLoBajGo2C+sKLWIRyDyWX
/o2OxFuff5SUWKnvUU0RXIe7BISMA7+e0vwFonh+ppUhHQw2y6QsURRXlrSSTzdAlHUNTJaZYC98
S0dbyVDcwtj4PuzIdkQZULmGi+Fh0w9T0edruAhcFtNcz21UHf1e2LNxnR5NH5iPKwJCZRy9Ko9s
f7utKT4ikaJ8UGVwMxPUMzR9r0oKNw5fzPnhE7eRGcy34/Ifw3Hc8my3ekg4VPLiCtpNW96Yj5yU
kHXTfcW2oDTkeqxXW0qBsxv3rTLSdC5Hq0laGVFiEcYqibF/6elWqiZl4TQKetbLuvDI/Zf8KKOf
l8jeFFHb/SSYjf3AQlY0msb8SAIzH5qyMtI3QQUTpRPE85LhzxPjEOuIZlAdcdTVCpkzWwTGcvZq
MJnkN4PwPts14caiSjX6nGox8qm02oNYjvxj9T6EYBDfDcuFG56lVhHhtdPiq9R18cx/npuD+mOU
DQJ77975f8Fm8SyPwxSRe5q1bBI0K7nI3xbbeYGGtQONxjLFPC4i5tuiWt90ZxLZ9e8LH8hTSPRy
rdy6SgL0nlofzeSqZ2rcIRwbh/i2CkflIwOXbsMkOTOKwnaaz6IJQ+d3UEHgKexSWs7OOI+wxmg5
AtaeQVLGFR1YOMC1gNI9XDIaRgDjE8VQfj609/dp8rbMUl/mPRqFkMKF/5mu8UbMh/k9Dc1VJhdj
o2wExxw97JpAZN3rgVHSNUdKwOfZOU7rD/rf3zrh5N3x0hlF36xAYcMU0VRWnKycdDD9TIWOjWTG
ASeBzm1nyc/LH1yYDEFv3UtbWAsFxDTrlbkUWABxGiOrUBOFAvQjzR7F+29NcjsVS06JyZ8KM7SK
YJkBquaXn+5mtWvKPiL4oQ6SjLLb/RQrnZbALBJMHeMHwlP1bkvrp3uy5MQ57GuMX2sUX0ts0XBx
OwTUyimfXucnUFFGuh/80U6MQlRiZWzo7jfOQoNCl2oiteNJU6uwMAdcT07YG/1gBTk9XeEYgCy6
URG5i45o+8NzFL40kSkIsrBPBJGkfajMi/GqL9LPBdcLeX2y2Md18FP9LWsXZU8inN/fMEAReXql
dGVHog1/dmNTTH5GbgZ3qN6HJlyyYm8Xs5I9l0+8Z1HY5ePWjnl6wP88b5xfNK9yK0x1B+s4IySE
uHmEJR7iE1lN8E2oW//0JIJuUbdPl9OWi3tS5k4L3vjiwInbtFGTDaX5C9xfCdLgehB9L2OhTNLm
Qoa7U2HGx3JZ04cV0CSK1L4DQvgcQdXytwESFMDYKuzb06fusUge4pDh5x2mZvuNMohi3YAFgE1M
PYFplq0weLH6Fku5pMC9MT2tSCPQ5Hb5kpUCFoIbzSTsUr7JdW1b/AE6h0TiD19x/hK9R/nVd9sh
Na20YH8KMT+fTKA0GBusO7QbrR3JH+PQSau6Co6wv77VsXPQT1AG2Wvc/cNfkWpWTskNhVtjLUx5
PolJRXXUDzBe32lojweDdBWOZeeqQujWexiqAfS8mti0rqqUBDeS2rASpSDcIoIddh9VRdDkdmQY
k6teqgIPwBYorNhBbHNp2Nh3G++5Hjpm2X5abwUxlh7B9n3KAyTm7FVW4UUYklpikXSS5U2V4FWj
tMolO8TOZcprLZtJt5p9hbp6SVBrjti6OZJmLtNiw+ZVLz85TIdJ6WNLBcIBzTEmXrWFnQl40/qV
W0YTlDiltw75OvAp3YpZF99qOvhy4jpg+nefJ53WBIfD53M8851LD929yxyuU785QHH+oXuI/x34
mwIyAOH1DOFNABiIsOqwNST4W6wmtIhrpQsI2tT5XU2kjkDKfZ9zrVYUwieofhiQCNId5+rX3qfP
3gGmEDvP6crEwkAdAbo/AhhBomostNMrAXOztma26Xi20wOrtUHndldz9gsT/70UmQmFWyMHuMNR
esNpC25gDves2dK91/LLctqECEPGIsT1A8noxCx+6Bn80xwU4xwGx4HonfuE56RwlUx8sth0PDhd
gt2eWbFFNrVh6r4anN6TJlouPzrDiRpvQVMlt2bK0AxZi3sjQS0uKKmRtUBRoNL7siOFAJSCvN5S
Mq1BXQe81kIC2OZQO45VrEVvT7nJgD2kHMz5N/8QOS1rlA0MNGb2Eaqp0t7xoBpMw6I5a2ydtBMW
ejZiaye/Q3XFTWTCQRyRME9EephriT5OM3bg/dWjDR3oxds3zaXXV8AUAaG0jkTsCMVoAHsh2afF
vCZmhJiAj6bgAGhJGsvzb3JvrDhESHq1r5XybgqGfon7X8wlDzf6tJHkaeYpnrq8ezKncYDtANHm
KqZihN7bRBxE69xs2ZWGvT1Tj+iwnBOLx+ouPSTJefCwQ7Zl17wJK8xWPJakCcWW/LPp9XaDrjC8
myWLgjTD6bv7Ycuf7zsFhA1qsi/+OWQluAFHZ70CetqNXsbU8V09pfqost4umTUk/DM+bZ2VWjf3
45S6ATYGFcCm+Y2jVbMF5RSZf20BYMx0EHyUAtMqPPf+MhS2TaPYiRzZlkXiTEbTPCk5ScRJvtYX
Huj+9QZjoaReC0pG+TJlFFkiCgXf16UTY3oVlrk4gz9maPDBIRwwPgvEKDtQLNZipyS9NyZ7AfSv
UD/X36XUS2R2/ayJzzfBbWmoeJGYbxAzt/1VQAciFlVvR82ULmVpjv2LzO27XffEcsr7tWpH47EM
/sPAmHaPvtgWn1CvH5xVEMnWkXsz0UQRULmWUiBSJ/79+ANCv93jve62DdFaF/Mk+dL4Q1mNozuK
b0OpImX3ndVBRiY2qUPLA2mghDl7dYO+kN/FMCRAdR5/PwSReESEcKFDMG4Gtny2P6ry8K7C/io1
i1GzDTFRlUhiyy8YeCFj8gHzy+OJYofo8IxlY8pIUD1LH+yvXBojNC+kjCuS80i7bJyAkjKkiOfw
pq8yFblqY/6kVXjIrj0zaaqZ5qSukWfqrmi6iNmLh0UWk1Bue24UHvbdeNRXDeRdh6Zk8dOabIVH
V7iYAaZEBpvE7FTlqcV5SY+1KXMkVyA8wgl5KLfTIg5IyFiWWs4/YyMjYLESON05vfmxJ4X3BRCy
UVi6VWZ0MB4Pym8MkEIKUtaxDhQaUOPvXHAwS9kUWddvouS50xR0V623UnNih486vpxld9DRrBCZ
0e+wWyPgqqHUX0FcCKfB9QoPH90ghJej3Ap8I6tpJ/R3buUFTS2+OmIwABC8PAXMtllgffbZaGaa
Aa6p6VeOa0tbkIq6cxCklGy7hsD2w9Wal89MAukH8UgkyjEzYuoOwssQKWaw+Lgx8+4jQuDdbd2R
M0AGEuIvURv5cJOU3tigkJnOwOhI3nL9OhPiQrL1QaoeHO7Md0B1q8LLfbuyZXtd0miJP81Tiqo5
DPUkpoPg82kH0AZpRkmNSQ16IZBuqvhiTfU/q7muuNP+rzMBrMDaO45b9iwn7Jkr2w9BdBR5nDQT
2Vc7KWYi6HaBpZ6BsEUt/SOzxcPhAxrAX+DZaqFs2XfLhFRh7E+ogKB2+8nPdBAIjR8jBdn/fWz1
H2QW72X18MxbyenPas9WMoZR8emLeWb6RgneJe4M7Rk0Y1H0xJGxyw4+mbAKgkxM/X0NDm3fPVci
Nf9uV1mIuII7OuKQkSUmXqsTrNl7XecokMDl052yxNglK/PD0Y2gzcmmRaQ+Gnx/lXmP3b4OKlW9
hoSjfGYri7BwcpizAWr4RavE7IPHu3z2+ApCylplSVy4UeNmPkRsrK+zY7A07HkYlI80xFaiakX4
6Ne4Evb73vBeBIpV7PtfNdfqrv4SB1LAaVoKnNdAuEFYcc6Fc56Z27I7uS4BxNQiVjcDS1lFZFb9
fpVV1+s7Zhqmc93mEPflR6pDM2hByulvopHceq9VP4kw5zsEBGT0MqryyJkFdKGPwNEgbyXmVMbp
H7S9K9AmL07L7Bjp99wFIHU6wA1jkudyu/EwhVZDgbQlWwJMP+dOhCc/D6+qRPqZn+ijLMULmnXB
Te7pba1Gth3Ru/Jhk0dE8Ot4xb2nJmyDjwL1mmEw3vW418iFSjee0Q+9+peOKf6dGzvM2q31uTTQ
FQi9SRg9aWYrXXQcz4qj+TOMZmNlyvyLrrTGaC0BuIsfMc2o7qdi9HNH8xXHIB91fr1pxxNTqStS
dBQl31QS6kBBNT6Lj/E/f/HVVpWPYTWX13gEmLocZSFoXJ+4hnVC6IRPlI3RTsDiETdGuVzult5N
1tO5UQpNwtBfvaUPIDjLzQNNNL10BTtFbMXHViDI+L1dYKVeqJq49uEFY3t1vU4pE8HPvwa9+AkN
dF65sgoV8MjMIsECtl0DMxTXbta2DSvgjwRWf3qHysvsym5tpvAcs2mmyglim+Ws7AHfCORpoIya
6pU3sRFboQcVv3QJuVat1U5nsh6xTklhgckQrSu1Nvy/V96+2qVF6LeV2t6XX7T5RinRE1vsvXTZ
EkU8np/vr1e0eQJ5K6ePFWtyzzkMvpVFDuCL4jZt9L9zgavFzNd/CwZYoY8BrI6GSVidmKAGHWNb
TRdZCEQludgQmOMxDoZWCzNnr1gM+1PIFAgBWvSn3NgF2+hWKP+4TLqk2I/vMYOpacDnR9432de3
DrxZzYzI1ht7kf0BHmPItL8/eaVDmSVZ7uUn2V8qf5mZC9gTe+xyRPD9BpcGuv6c987/fZ0ojg8v
UwxYuNoYgWpDlhqLINFeZqr2Jgch352rSND91NqC7921YyoWOdW0iUbeLikOpUD3iYQsKq3dGZOU
NwI/Gnn/i3xLVCDJXtQPzxpKwWvBCLmP9CEoOuUCxEQNUXxPntmrjTfv8BIOjDvEzcpHpUb4EWXR
13IU9Vpa+W/g6ifGpiNbopP4ADbcxlgJ/jJ4Hyo6kpsF502SVWGK5j4HWkhNW/a264f0jaT35guF
Dlg5ZBKjDnhWQeeqUYMHnrPj1yZvX6mvTYmcK11WuVWHwL1p7ZeN5VbSj+64GucmcVY/Jfx4AtGl
R1XfLd8fwprqWO5MCrJMqh47X4asinelN3eiCmDV1R/hSVetn71pKxKDYJNmEhXwKgOool81TKvo
lacPZXkBaiF4TcY2N8EcXHB8sYSYzNrLw8qGlPBpIeehkA+AEq3EOYzxSPOLs796gFaVAcVsuvXZ
jnftTlSkT6j8RTMyLYVIFHuUgo+RUKt7IpCrXq75KkVGChdkQVMBu34mYBsE0tbucS1d+QBdGSL7
F82AIaneFlncrgzetLXMW6YL+vlzFb9B+NcHVgesxOXaufqt1CUSWhI1b6IocBRC2yYVJL1uRTlv
nilo6gLP4YRHbyB/l3KMHPtBqmM0V8GlT2l8ymW2HFMNqM2lQ9HEfHYvBdZDeEYiffAUt0adggsB
/hN4il5q7fIZ9ohJoCNcCXb5TQKafhrpW+7BCYAlC6SBtXnN6s0w7X7xNRPrAtCkCWcUkbNUSbgV
3Z95eT2uyHqcwiuNtXaCc2pL0WNtAw8kmTY1xm2Y3vnRnXGvGCE1oO8U4x8hAOa8Ab2NP7Tog1BJ
zbGKf/RNrYohQlysbgRJQXjioAjD+khvUcK+YpPI8qto7uYUDETwSe/+SZ3BK2xVIYUyabrnKbLq
Y7T5eCGaQN+J67ad5Cn1DCDxsiXXnKpbmDjnyVDOzY/eiFj6/UXV85DiG4KQbjtKz65CQM3CXSdN
1nNQOUr5pKj3uRgT12XBLHEHWJelWXRK9t6GDi456waLJ8lTN6H7Dk1QMJm487hbAMFaLdLwEj7M
ogHLpt2bJ6vjM+HuCYovvgRayWemjwA3v3oRwAyXPSz68tSMlb/dBB2zSA/NDLXhGUQLwLy6edyQ
it4lLaEExJBJ8FqBOzVDoHceGq1qXqyuc4HbMlwo9ZkoDrFgCeBgF4X+CFw5BRI23LgubomL1W+N
rHbFAGDgCYCFoaPiVPnTNrUNlvIyaz6tuWZTvw9a1vmVUBlssvJGjAqGX02VFq2nEnLNIdi6ytUw
8kFYdVCtp8MJ9xp6XDY6KFazZIHfUIcWelwaeqoaKsoi/JQrQoPk+dG/QMvqUuQqrt75QvPFs+i/
7QgRMPe/HiVgZx+YEUkyESNdaFEDHZUO/z5p6g8lEtVe4UcwU2PWfsBsd6HmpiE1hOczyrHSvnGC
QgiGPBHd9zovVWeqzUAoacQqm8MGQ1vY6ITLSXgPWqBpmMDvfWD4YMUEZav4zMOtTVJQ9MfdOEEV
EbD2Dl7776fphyXj8HOGu4lr2qOYj3lIRfurBhAU6aciOzhRRp5+L0BlVUulHnPGZqGhR04WVSFo
dsEYmctpBqcKh4T7vkarByMmsuOT5MzH+nQnigdA2u6tg62gITw2Ht5vUIWFkQMY6opMoexZUfsP
2bNwxV+z8C2THUUCBcesNAm3A6DMouyjSTf1Intb2RSdCZwo2eYQ9FrULog2AU/3GeSXwHxXq0Y7
kucMIjNaA8ApcjD/2ZJjqUJzzzEH/lRKJ29n6uWIVY7a5IghrxS1vg33VD5AhinZy/Pt+z8iEqcc
pTDvjXxKFLFT4ArW7m+yfPdTslUM9yhLsb6GrWF00alNCnl+e2puZRrvKwyd3h+y34X1oe6Ftrx/
stACHkBBL75SQeQ4io1pbc+pJHSQOdrQrjmNmnmg1Sm9gw6kjec4xHb0r1L1UAZATZ4k6lOXSw0S
W7K2UdfjcYio0Yihtv9W+7ilI+vpsBbrSMYjjCfuA4p2wN0BSLx0+eCWenhcIE0rfLKkvYqMfFNa
OvH1uNxYjYsg5WpHyHKv5JAWi1tIxpcD+uvlomM/n0DWI7/YS27Gu6g74opEVT7Q9d0PJqitB3gD
sVRZyaDKJkTzsWVv9zE4PdWEW7hOyEI4NJ0oX7SOAju6+DWeT7mT4+op0o/D3fg7+lkimJsltJ9K
oh5EiotmoeUk08LJO6yLNQSCF0K716hOSL9p6IwtCxd3ibMG+Lgb5mqQG5ezkHxaWAbGHEaahS8L
yLvk8J74s127fdmSl4X6Ek43K+lUwaMybbtzHPUuh1zO6AmHERx/cY03W9PEUg4zWK6jVvlI/nM1
28bRciIcR743oWoipoakRCKFQek+St+q16sYdlT5nO4kPBJPD2cO75E9NS4OgcCFoRmqoaAb/8E6
fnlqsr8XRVw1fyIMhm0gYiqdFgaZhXAQKwJBgJSIPJh+VpD/Aq4JySm6Xkw7j547ut1TTIg/iijv
UPzmvGPf+YIIwHRK/SAZbgCFj8paUQPbMWa+w6RqYjMiqGmTomaJAs1hY7N93M1pYonewkQ5efP8
+h4v91Vao3Uo1iwKRw6KTVDYMFADvXJno0IOiuZhJpCTAn5aZW9Mozt+e99z0WomWUv62JFfIiD0
Gy25n5cF+eoibB3dFoP6PwN7Kws5Z0xtacr81bzIzKL8wnVDC0ttuuKiWU+49lil6Vv5KQYv1ZGA
ehqfBqT2ZieYfy9SCTJwkYnTo2BKcxXJ8QzCgwXNi6Ez+n6sWBgWaaacnz+xqSwZYn6aRL8MT1Vb
L+7l9ey73cfGO6Amh4qHSm9RJYffGZ8/m+HgkS8PpElC7+sbwHtiKmx2oKlSdtmJpXIWVLx9LklY
aRta2PSocA4B3VrR2ZKrtribOxNVZtW7mmfSV2i6Xe48AqD3X8QzS3lQ5EpTLaDflH6uTBX/zlhR
YJjTpqz4zH6AkVgHNyfzYhSv+Os1rMttT3JbbHwbtlg3Zy6MrMzvo4nv8fK5pvITznhXSG4oeRAj
lJFILvn8Umic1tS/b48WFQBwL0myZUgqCe+j+k205OYEEXyRJ16AMpXpJEQAPIexYd4s1Pmr1Kan
f1DjOG3o2+6try2jwj8Wg3W+gpKNbU+PE2aa/2Z0VMd0KrkHNjPVlrZJ/hjr3HUU7Z04v4rru+Qx
gmJVFdDonJ3Qg19WxTs6R5cj7cH5fDuGWvpQmH5NWMEJwkDvtCI8Q4lhp9dm4I20lLDi23JhTlsS
w956PT6BkNoqeqw42/GWa+T/0cRvtAKm2cPwXttYxoe2dksp62y280WwC472eB4fhBilU3O4JX6q
b6JrIxK+6VmG2dMtFN9F9k2eDi3o7gPWpBZ7PuF8V9dVz60eNj0vLmOzBS8iNAZzpGQ9IvNmOweL
pL27u9Hh2DqawMZdVnB4CkujJZHpLA3bmE6gPtj3693SVuvucRuvlxXimYXVNIZFF3wvC+HhufY0
j7LlUCRX4X7Po3R41JPlE+b4NohYeZKWhJcqQpmWIsaCBcTpOAUsIxyxiWWl2sIZhu7KQKpB5Qx+
vcNuao0cFEW9RKWUOTkPJ+xf6fRa7NI+qPdJM8GsqF2ptdBb2dCr9/59n2W1EBaZiQdGvkJjpc67
5JZx2d5q4fZzCmTyBeZzR5XNy0x9lec0wOSul5xgg51Wqf3r+OFAz45BpKFCzs3hWQ4uUG+n1E6w
hq02tcysbDrPPW3BG3fnadhFMElbfJBHevtOjz2J1InebaDwxvt4Wj3+Q0e68He1UmMAyf4bIMoB
lhMgxPyBudR7fMfdC0DdCUUQDCDIdmwTMxbQ4Iw/d82nBL8MLAE4utIs8eEiS2DDgS/w4ZqMWSPo
qtFqVQvLncQn7hqrBtWFnqwD5Xh8z5e68e32GMK2OBSOXc/43B5lUyTAwpwjwSHoJ8cR9Y73mt51
oehPndRTPA2eAzbEfpziaXNnIlcCJ9L2CqtRqC46MtPqYoDg4VmKLUAKPmlSLjrvacpeya8gxcY6
AU65S33zBnxDsKNvbHKYweTf4WRpHmZisBbSRE2eMEBomhRLLykihecy0IOeRvvP1+2LOdOcVIAd
SnEmCAs3xJas4V68ZWssyDIEL3PUHFrJ8Kf4BXs1PQ2ojQ7exe01ACcLRxdG3D4BxSWPDRfjSYSP
v+ft1iq7dnWESrn3O3AbPHisKTF7KRXbvdNoka8Kvl1NKZSYfdYksjA20SAH1vWstf0AXK6mQKZr
T7SnnQJQpD0L6dWOuC/U2ErU+RQnPZ2xpfrYpPlI297AQTHRQzWYWPGTQMfoqInVyj8Y2p+gs2Rp
mRXq3AgzgU3LT41WTQVowL4XlyhoTKRK446I3/0qhptofDe1BTMK2fLRZL1DvoFzANuFsB1qJzyJ
lr3V5VIvzfjnbHUPvTM+116IljttVpuAwebWXOzbT+/8kP+MVR6GHuD3mPu4uKajf/rjuGvlCKqT
1NJs9nT/EXfOcnAN2mDdFENrlJYH6ENUTrqIN3NFsKu+NYQKmyoaU8eHnqZMXhbwgYhMV5kuK3FP
lb3RTmh9J2yXqUgVtDYynRfbrOeDxxQxCU3X4w5/OUrFbEZgxre5qMmnr2ZDLhZSg0WXKklMvUtX
/WtfUkOrMkD9lgG7EoU2Wvy64bo3he6A6JwqdGwxz5lRGvf5yw5v3tD5X91e1TJ2Inn3uivPcN+g
Xuxy3ey/Dj0Zwm/bBQjpsRbWnzA0VKrLooMrGx9LOrrVWVDX88ApiyFIdzWaajkB5h7+IZMYK9sp
aJYPJUj2fRbSRpKdW19yeOPAEFHgK8mW/XdfCHVnWv20DvHWyeaoeAyefkolXt21kl7ak3ThuqyE
gDl29a2r/r4YYilgJrF7is4vo3H3Mv1WngS47cY/mB1FlbBfe2Ay1zl9JEi+Y/4MgjCg41rUxD4O
0Y0VYLSmE/5w0pn8yKkUTjQjDOF0Pmj+7gAt9gPTF+LsYjua+2nxV2AciwqdYwWGI6mcBA4S5UnM
FX9ntivRhhYPxJXbIZdal1pCxuOMU0efMcEm0H65uHGFyEETYV9gh7CngqMse6EF3exoyQ1XBHoy
kN4p9oI2miFyy4BVb5aF59tQFa/iRNlUr5UYglb57N4xn4k/ewWt4kub/X53cfrINmJ4anJxv5v6
ms9KQnZGq70vaEMmW7HDBAMpRYQ1IlNOLH1rOUS5Lu549y3x+XE93fJmgXOQDQLLwDvDV3+G9dET
+fkmXBGRME72UyU5zU9JxT8lk6K8RVyN26bRvCfaiagxSPoyW7ojwXGG+9ejyMsrrhMhVYvREtny
v2KmyEfJmo5vUQuS2z5B7Dcjdi8PpyAUQUkEB0Wt3ZmPSzK133UHqets2kI6nkV7HHY/S0rYvaM5
2N6u0CKdmqwma7/7kj2WnrCyI//cxjb8VXjUdb0/E042Imy37/X8mIU2g4yu4QO0B6Ac6gUNYMIB
EcP6QXwKq7jtjHmKhe5clGLv4k1caL1bZSdDXJphtuyj7lhsCNZ5JRR7IgmfqRqbbTbEzGWpVSp9
LUjFkyF00klNf6S/D3lBsrbRqdfl+dquh1xqeKF/IArbUwSqOi3y9svOtZl9CCwx4tjn+QCkgk8t
BA5warkUzQNlfT8xJ0ovaohvBqwv2Qak6E8KYBvBjRkiCElv8uW43qThR6FEbKK2SuQk6F+s4X1j
7GPFXWTp0p1W2q9A/swdcudr8Z5d3OPMeHXXRFAWeqnXaLnD2DpXRswdlGPFr0G0bd4M7pD4gtO/
Ruv4gl/XGJLPD8yY9vgiCSDfvMa6M2z9o17Aysxfordy7Bs8w38JTMbcRZLPwTh41W8n1AJHGzm3
7MADu8Kq8J2O/JGJ7QdN2PEz4bwvLGhr21Nj/ENanyeAcES/HfsbNWIqXeLn0ChRjbkWVWV8Qeg1
ntDwYfpAnST8TwSOvlHJfcLKf4E+ep6SGP2t8ut9AbOozKCNkES1t4HR/2jic5goma64IeCJBDOv
dlUE503Nfn3oq6iF3I8nTWc4RKIEUg5XtJkiKF/nVQ5MmAU0lRxHn1ev6r6UPgv7O0M/yE9XQZxP
jPxIwDPGz+1xYnMuR1GgP2bQBCbVI8ktyXxot01DFOkdHBv3aTXBnGQ79PpoIlr3H1JCF/tlbU+y
XYy9B0lzrDltcni4sYggo/U3BphoPtKY9ptPcZhLUouHlp0lDgO+UD6oOnViOX1NxDwRiVMkotob
wu5Zv753hw7Zj4ie28K7tyrZQfV3CYX2oUijz6fQ9X4KCU8cOO6BZuYm7j7Sq4ISMYYe0ttgPUOG
6Bm76EClVG0AnWz55Zvn5djd7uAIqN16MyGgGFWe6BrwtSwA0D+q1EqehCsdoEareo/cnM6MLwyx
rb0a1+6cTy964YJ/NPw+DNH0KiwCHq3KvXAGMMYu33J/93+9XwLthWqTHm1//O+GmIMnOFOgazyN
5erCzH+tcVVJsdHjaWGOE6GOo/BVicrpPGywUvG8YyeJqHE/EDUZ4wvK6zsgA5DMBQUlZmiT9Xzb
Ia4kTcD/HNzDnsE/ReAhD5pWiwWtzfdggUpMzXmBzQRw22WuhHmwM3mwQbBPVSg+izJG0Z92YYBS
s/u/IypMYLL0bBUMJdzbku5MVlQCCoO+fPJsBfa6Cf7sFJzXa8a/Vy9KEK9AdYJEY2cHoV/ZbGU7
4pLQ5dh1I4tNqwxnlQRmJJUsBO9SI7qMgb/WGvkG5j1DQqZW60bIA9/+hwvl/I6isXGT6OHEqtnD
6+yvCeIi+uI2jVW1X/rtzOy2ltk3u7l9RG3zVBRoOSaND+hN5zI/jkyORghsZKwuQx1hq3bDBf0Q
3Xf1IXNbhmnXJ7FjOLjVNsMOX4dm9mciQ3/ZoIJJaBSYck/unrDnP+96LEht9BLA23rzUzLz+rW9
PWN8pum0f0lGyvgyEVlIMLBsNTDT9iBYYcqQomx5FXajSYIoCDce4MFKwvcLXV5abc/ZMC4QS2MZ
GDDrSK6RtFp8iJgpyHUj/3XoFRqI5BmkZ7ATHrRQWC80yLQHRLf6Ky8mbrAVn6SjtUAzk3oFUhqX
4qbd9TQ9ZZ3EpVxBO3oh3IC+a3KRu/eDGNG11uRM7WqGnvHTbU+sU/XWV19oKRCBlLlNwapGtTu5
bfLvFffF2ULn0ExhakjwrqtMIjkSWHCh/PRj+uH/FXRcMlEpRzZ7dqGEzMq6c0ZIxehvm9YtdNL2
U5lyDeaY3gD5YyfVIl+uwo9JmukZB6uzK7bpCQkZ2XGlX+z0l+OY9ouIKIAVPMAdmwQyjUjVvY22
ObcS+1TkBdOJWMFoklkrP8r4toBmUZKgCra4RQGAfMBg+BsaFjmGqOTGx7INkm8HrwtETE3pFwsI
6DvVon5WOoIemnyv5gheFaz+TtEfmscJKndwN0XT8Vnjv7sA/hFeSyxxZmfsjNl2/2R0kwle8AhH
zHz7KZTr2hHSlT6BF6KST5cX4lBA5VetP8vKSKpTG79j0mTftnHdiSGkX/JxIMu4JM4Xc7aoZwZX
yQtWHOV4oUJPTxVDPi+ZnF0PMG6r5QMrGcUKxp3HQkyys7tZQE2Nb1GDO25x0hr/UYQZ2QjJ5kTZ
2cxjgit36lKhpHZTC+zy8slCv/F/yuQ2ONUPbrPEONLbXYZju2YkIhQIjcEZo1Y0s94QVE3FOzZz
Jl98WjIq1DhUZF5UhiMrSTZW0hGI3HrXjehoWqnvmNb48HQ4FZkZ74RGAnosf87zAy9fT6+S9lnT
woMxvH9lJ2BmeYjrmRQYkGG7DXFT51GaGH9MIpQRCP1pMbv0tpz5z6Qj0/32uxCduk+AgR/ItZkW
PxbJcQqL32iJ7XiU/qkma0h2ydVUjHWPPvTd7Mqlhvej5VmSqBnyuSg7I4R2C/MI6aH8TETmqPGX
k53Wqxc3NL7gJFVZLoiq3dysNErw2bHyjx7QzyO1TSBOankbTdPl4tYnvvfO6T4qNURj9+wT20ZP
CxSjnc1PyoshpYan+iKuB1zfYe1xjycUvW+dSOEvmPxJj3NfXQ0zx3jUPt6QboFox4LjhQ+Oa6N+
rIIUvcrUn9vUpEk5k0GdtMI+Vir8BqnwzqKr9aPiCv8exZtz6ZfVUzu0Afc0/pURmizNZn94Z+uw
vpCDmo78Ozqvo9A9gtBk1FJ5Ep0YTDXwfd/oOxxbE8iCb4yOS8OwpccrDeW3+CPoXDPMuB1vVlHw
3I4qJjT+qIMTMhLuhZrG+ijHF5YreNo/S4o+ZniUrmqj1z/pnhVh67VJoSg9ZlGcA3ZrBfXSGy4r
asSXuEhYVC8agwEQnTHOUAZUq7m7KgAcRDh/Fu/hp9TAtOA6QqREY66cgIbTfyPT7TTU2ERr/2I2
NI3qQ3QT6iJUYIWTvcl+PuqB2EB3HMuodQg6O3AACwmb7ggJS6rP8rJ2LrLItyTGM8NM8+8LPTg+
7AttbXwx/yfz707CAulHWMOeMrN/XuOAjkTQL5rQwWvH11U+LjrHjSZ9VYr+myKYuXRy714p8jMR
MVVhn+AJ3E9WSR9KlrkPfQnAFh//roMRFpjq/uGrr8es9z0tcxJGRyjJsTcvceoIFoU90yfk3Db/
W4YMh2uF4TnYGcwZGpvOz0thooh2sHm6avEYmy/ROuhEVUrHecSJLx2dAKWEzls2jU+4C8Z7sByc
8IuLt/JZ76V0YdlaT0zCK0Xd7s2rnRUQLNcu8g1HZH+Tfajubg6JDGU9zbJDr0HJpHv4YaU4TXk9
X5WE3Mi6KRKH+zJUrZl8R191JJ/P0pjyEAn7CFmMcZMlyKlh/Nsjb80tFUqfZQXHwT9VwcAmlFRo
WLEV4yJ+Yb5SXtLnvSmYAYLt2WUDsSR/TTnMwpJKq1OeUV3pKf4MT+4YiX+SoxbA9mgquaNUGENI
/cVTnAY/MelkFJUR2GpqNumRID4R/QBig4Yd/XsWwIdpIDTcmOFhLVG8raNAirkRSnvrLB/kmHLf
RlGUgnOaFnIKV6qqG5bXNUnV2+zjNg4w0W8wJeuX5h7OYgazHBmA/i1jQpXCA0SuOqYl6bVUPuH7
5M6gaaGOeXf8rdMtcFjHISB7og5xIys4+wvqGyC2dEaTtynf9hIgw5L1mpKhr2019iWjaI1xrmzg
E13mUBfjvWBQQ7BQfmijim1ra2zXiC9cXSxiy28LibUdGPUF/9nxmB2LRNNXxzhVf15XsKYmtm6N
fir+fEN0z73Ep5agG3oyfRSGviFvfjABmwPC1IRynlVRsJlox6HR1jj0aWvDqGs5mE6NU8LsR4/y
QwCpgDzg9GumZiQtJZveYlYVLFpElKPjTftw8CvBNYiV1lJoYIJ9I0qbFgiKr+mYgKRzie4WWeoY
LebrtoLoFGT22I+pNkE6LSX32yWlACp1MPHDbVz/t97d5EXhahzRjwa4L3iazJ5WAhEzC9VfIfg/
so9HNrUMPWuSTO33B1kyYUIaZD8JImchiEVgddLyr7OxlaqkTjZl+5yTIKr1XYTJbaFResXw21my
n764mmRxdqD7+7yU3tcJ2x8ORUWy6Ri8TAvdtf3IT20JBNc7XojcWWHRzMtHYc+YbR1E4jSKANLH
NDv9bLoRIuPB4OR/u1mLpOHOrTxKawLJ5URLDVIjG2BcZYbnDrwnzS0STJImjmDdcA9DaYz2Wv2s
8F1KwurXAe198tPfhXN/NbOtotiXKKx5rK3qwe/9+/veNu5Y0Jf3qK6eXE86yMCGSv+DICAeoCDT
F1pIUbvoXGGetBNsCncrZcbvROUX1IdIB05avgLrf0FHijR4byv+pmqcTPiC0pBbNJOPas7PgFGN
CYy4rzrcY2xcaMjXLShWuUw9IkDTKSLrO9JtlmIjAMKaDm7ekDQf3/M3XB/Fsc1+nOMKLmdVNM0O
XMGbzOtrZO468fpehpsHOXIb/P6J39eAW5eLMwASxJhNbsp6ZHSphjyLMAsDmpdcIySjQskAVEBD
LlrVb+NtQZTqijbIw92Zh0sCenEprF5OAeZCoIx6zmWDPF8YO7Y3JmYixAEuJZFEaHbs5ceF+/JK
dQkAmjM+I1K07bMU0fDSxtzJf9DcR7RwKDQd1hppTmOnEIOEua06GC5ZJIMmgMKzkpluqumAm9nq
feJ02KWgbVJqwsld/Y9BkIEHu9V2ShtTwF077aqlFrL27zKlUnxC/qNrFiofI4+9zN7siKv3bBbe
a40dgxxf3inSL4hjgcIDrMCgbz6L323uxScCaMEB/WzbUpECATsO+QbpHiDetTyuhmeiV5ELhvSJ
WM1o4r6behd31diZ/89j0mExsEYQ5/fYubXwt9z4M1KoH3HlFUZU1TpFBg9wFNjPgx9CIm7F4qWT
R/LRSckFdV7WHeIYI4MomSntsv6inZV3s67XZii4knKUN5XFHnRNYmDpcnz0ArDgUepDL2Lgsuv1
IVtaL+0iltr9KOcsmRWoyhwbFGVrof/5Pu4VLECSNLf3mm/vzpXlaXngrCRmXgBWLMii9uKp5v6G
9pIbvBEA6ZRRoE8jCdxqhPHlNi/TEcwYGreAdokvO5B+fbvZGP1OyMN1udgiaIqRLcV0onu5+Erj
G67FE3EblNg12U8+A3WAKzg0HBcJRK+O1iSUX+11Erj0E/7ISes0D0oCDMHXe4KvULNNibZFI8XW
NQLfu7LRq3EfkBfjQKsWI4nXJ8W3QFh7L8ZSaxfBCfQXnZBfXFX4PSh88ogAQEhv8S5pfoM80zep
7XA5VvX6syoRbO9EYBBSssaK1PJzDiG8mKhoCrVhs5IR1p3Q8xdgEueuo1X637c1Kvgortj3kVv7
Iu8Pyzq7GuanHBT1bzX5PHGgb2a5z8JEWXRfx5f7EmCYlxrJ89YNMSRg874bnbwV3M2ALQ53EoCv
gaBDOvvfYpsiTgoAKjI08EMDq7pEIXb6tOqmIwOE+INmjuDLhB0c4q1NxUckGiV+7ngx7gP8pUfI
+P2GNPstBBUNE5L97T/9qehXPwmYqaqXtKnY4jHHTA9KxwtmEB/CIANggETr/Sv8fS/S12UC0kRR
8MKSzPOIttA/E5ajEhMRleEYkVlUzoboSwB4oMn6sXuMEk5Obi3HGcGpHzkliLhpIHG9WlyzBDYg
9MUruCdGZ8t2HGcMgqSqDSzA4/MTQwgrTQ+kiYg2JRo6FpM8UdaknZja87Cn85+ttbZn+gP9PiyG
Iv8FN+aIoy0zmQNLtGnOARDBKJ7G1nT/dk5V/Z7UyimdJm9JCWlupQruPPARsG0zjPLWwI44v7ne
9U8iqKnLxYw7AW509gQCBl/gCcGBgjaNwmNL+Ml6J+XVpFRr+SZ2ldFhpUC9XQjjRih39+ENFJWf
rh7VfYmWgYmLj20iL/LFVLWJM7y1xYgVnJmjOuE/My3tsseGxUjr2lMZ1qmoqEqmNTQ+vEd0cw6G
S2kZ+0AsDNXK6N1GTdqbaD47XaDdV/xDkzGuR1IDM0P+XLNCda9eBdRf6QIIekQFSn+OsJyIDNPE
GCo8HaXozsYHDHTsWC9HYsYCIv4eJ7r+UKCjzF3I5RaSbnp8dzdG04ichwlJKVd+8V+5Q6GWyAFS
mK2p2FeTcWZ8hFCEGOL0WP3j7FBTEBCIWBAAE71KcvL1cssEMTlLYCr77daI3/Y1wqL7Gwwyz0/N
EfozWqwHibyrydAxMsX+86u+y3mFbohSkIzY6PqQTtQIk17yEHtO0WSpM0+DKJqDKvuob8JouO0y
WYZdvA8IzCssk/INoQWnJlCuBS+3j9dQnmm7RG5tTyZSHn8b5mQjOt+oMkdcAUa/BgaOqHc2OVBr
ifMzajkLT1UgKVMBSofdC1FSIIXlP6g0dhRK11YLb1XQZ7sHhcI5oJr/6tIhYNbcaMZ/paRDwyL3
mYpK+pzaPh4Ufux1MkUqtj9m6Lqw+USUk6ixl/+tOE0saaV75u309gKHO4UmX2Yhi28yQFHJxAWd
NIetixMfSgiFJ7u9GHkVJsTEHyvE8BD+yE6m/MBkz57pkkvGUNfbYKfkk2aakb1wE26kb93WpJKL
vjFHtrqXVdbqicJMFVvA1hjyBo4RnFnXfuuFMhfchLcqESwhJo7S+bmdEf08tgyCQMmItyyOGkwU
fAsbWHmkPigv/g/v4fjcLQXol/Zx9N80UuUFu56Rd0oC29ITFIdcSnUTAN6yKeGbD/TcBeEkqILY
nuOqhU9GUcibEvtA94dE7tvZPM99Y6itPpqzRQkQNALcPahfJLhVNA71WppyIMI7YOeEyPNXSILA
UFN6eFxlUxh9dueQWl3Udze3h4eXuf3SAqJLtWMa32L7uTkOKvFPwRwJPLcTXl7plFcnT5E5+mvg
cg5n37/meMVA8WSaADQ8doatLqgrYGOD1i6Jgx0jU1gPDssLD3m/3l9Uvvi0s1UFvnQbCjnvg93g
iOJNuu1FAnIP//TrcYuod1FZRcVrPW+VsOrVdo9NRcIOHXWYl0vnrajf4cd2uvg0PZPvhyD1EzwN
Hx/0K0ohrbw5+6K0bHsYmQUBW9Y4Xk+L3YZHNziQdzTUfhPHY9B7CtO/wg/8VUC9ffYh1ENV89IC
a51pb+p7SGmCzL+XbLB8vjrdgyur3Lq9gef8UKAme1vgqQm6/4fRrhZaP//qEzIPwob2ctK9z9mM
c6zcgl4LowXR5PrWSK1flcc3P0X/7IcHXcN9+SF1Bnq24PXi110G4mxW+MZ7Mlidcn+KXtzGYq+U
1qUoBd7FcjeDiT24NafeS6XQ70luri+jbhA5JngIm+1dWmlik68K9UwfEVzIqKx5v4S/EfKmtqqe
TvKCcP7tedYGvyvhzutlw/ZZrx4z4VmQrb5+oU2nFtPSh6knDhl/xdNUd89NX1bD9ugvyMPd8Rou
X6JGwugq5E+WTbZwWYBqW4i54GkpaPUuUHfIrVNLDmN7HP96nnz8dPmpaPNpNSIYqm+BqOHNYJRF
m8bMBpn2ijuLDVv2V+RoijFA4xh8boyPHe+Qc9Xbj8G3OobMw0tqjRfGnOFFyeI+gCQoHIS9peMB
hyyvl/dFgf//NgSohY9CpIRjZkLok6ooACIlr1G6EhCCj2D7HhtUepHl61JATJ8I2/atTXsIz/VV
FYtpYRtipnIMzFPaTHSnZhdG/Grec8CvgI5Z6cHxV8qCMRpNup6TBXj3GvwjVK7JNUMhXbQzn44l
UEyaaKdK8GOSdfhb3KR1mFN1kKifR6J9+Ost418ML1654npmpFKFc9/AJaj4FnPG1AmNx+IlKnfw
uA3O605XWPOODxDap8Nd/uaHWdiJ7Qs+eGG9tnImSXpvqcJnaNpXqLBfrIgPbDHDsFjHlexYLTnf
RRinqy1AJzKPd92bxOFDyLQ9vlAQsh8T09tQLlrJuupNhoknxSWo/4X5AkAPsLG+k29IjI5o56k7
8qb2qmCQtSsTP4ef9hnyfNpEvj07N9amOYty9ndoKi5sh6NhIFtYC4vY8mThgN7B3dRVEM+XzPeZ
Ws/V6gjHywvIfwLkrOX72p/+pU33Bihnl54LZV22j1lwQkqowkZi7O2ZPVwXQI31OZxkvEsAWypC
Ypjzcmqu3qb+TUxkxujCR6y5d40Z64oMQ7osFhSAA9ZEAVXu4m3kys44jILweQgfwqpBkvV1XVzd
WpPrxeTW9ZiQZ+LCqGjIHVQF4AeeudBZLGjwIan1WZflcNCIlWxQxw7Y+XV82z7W4zJ5nBJHCuvK
8ww6L6M0dNu0jKLvh8tK8szYgbbJETdpJA0g4yefGN9hZ8sAzhZK2Aor5Yn+2/+JYS8Hv/fRQmjK
34607BAeLUQZB5olsptjYR6e69728CDtGQ8tSGpXOZE7LaZKQBRfxieyz41odHQYUGEe+PFsa+3U
+cOUgcM7bFW4Xw6vVagWbDE/pEkQlucsd0jz6YNq8vWJWFeFkHkbV06/yh3s0nFj/+buQTc3Ki0F
lppeqPaU4t4m0vSnau+96rBw8jwZXHYGE0yGSVj+33JlKP585IS2QPV5giQH4EDhe+fhkYpPD3qQ
TQaxlOmrUjH+5gYngJwbk6eDaymqEq3WZXdJyAEC/ELT6s5/JpHW/EBo9qDX+A68UTGi4WcwAZmz
UvUFp/odpmFkodpZxG2qx9AoMyWhCSIPXswWVsdpGBx2SYfiiAfsaCUkeSaG8K6sOrHVWXTUTf9N
+iZwhloqYJyRJa5hd02mGdljVNBlcvEbnfWEm8ZEFRcYQZujO+Ohg04oERkUy2UCIOhkCeuXcrFo
AWJCUTT1gM4+tnTKY/BltI5rH4axCRijPM+Az84/7t59ywY+rJ0TAcl10bTvZYQgPuXvXQ962qPo
i7LXAreEJSrtnaYLt+WPLMaUxeV3iCnNMRA0OTokQxZdRInnsZjj/PwRhUI4Do6sW+OUI0l/wC3r
pIrxLOgoRiZj1kE2vXny58TksA99qMfa/KCOaX853q/oXwe+5qtNBO05nc4iBCLaGiPZeW61cp6I
X93zgtl80itzcDPgFAnFXIWsqs4CyzqWDsNQwrQXHIy6lTL8OFQOKQNMcCsLWO/jF0Mn8reBsORr
fwcwCIiXk4X9p5V1dBosn1Yvp0xvfuHQusi8frYwJWUWmCxgKfG8JD7iAJbVWrQMLBaKs+c+Nr5n
LDzRWTuDkEd8ic3jvtPQqy1M6iE25ZPqajJ7E+G9X1OS+HZrUDVg1bt2U0pmfklEVlTy6i10VnnY
vekAzM5ddguZC6VbXqCqH5tqWSoGE6D98g58JHCKDEnxote7bkpu4u9PnQuuq/YHXOpN9juvMut9
+8JAd4prw7/EuTlfbtOX49AHrWI84o24Kh4WVqhyTPzc12FzZlk0OTIaHj8hnyGqB+m0qJBWEqFE
hg0WEYLo0uU4r8jquLT55+FvVKqDHLh1MWUGQq2JYmRQwRXBF3CYCJtPSNJLVlj/ojmunZB/wCoJ
vY62Q9XPNnl60pfDXS2qtV0Plnr0lld3yJHeQb0mYyavKkUNnKSLdWtcE0MzhqFDNC6i893BKTjO
GNpLg/Hm1b2k5buRlSw+K2DrzuGqfB1+beawkPJ9Ec5TdOx5lEpiMag/zA9nKc7DxIJQwlhWZ4A5
h0+V6lJhJSOHgWrqEVpAKyzNrEBJ1AYei/c5eR1tS281udkKoS8twHAw4HPIBUEnOlIurdJ9+wIn
YU2getEGGEEAhA8qoRvfr7xwdIBLp3znslkn+8GQ0+yOrU9BLwPVlkVgXoGVQKLfnvIEtrPS5aJ9
hNn4UOJvlg/pa1kt6nzVLHaadE8jH1fRORat3m6eT6Wt1mjOfbNTJXUHLW56uOkcitEVY9HVrPKE
m5qy/P9KSTovd9Bqc429M//KAwVo074Mpyt3/r+K64PCjOhoJ/I6AiQ3spAR+7a9yztWfzkksvuo
arxxOs3LcBIj3YSaOqYriODtsWGx+JwjS/pgWVZZebkfPQl30c7P5BO+LWGya+MuSJk+z1VhgpWI
TvZat0VGsKmdj6JnRoyQ+TQy12kyIDBqhrKWcJsjbrDic4vo13v4oC+YtTXYk70rmCkR5EbUxr7s
5qKx0v+Y/QwoN4fnJPcwnQExaluacerdGRpUuUyf/62XKg5tqoHndZuF0Dfpj2nD0y2S5n5I1Sra
uV/MRjnLlp/yj1Etr5sGheo1OXXLENwfWmj6u5RS8tPIx2RJ5iKMn/S5PD85kIfOI/R7jSyh6/V4
v83llnzydF8p8KEKBL8X5xSxXF6iIbO0JqgLShNdJr9h2kNhGB67g68H1cCcNezN3NXUOTkLxro3
cmYuPYKqFAi0JD8ZN5mrx4k6w1e4gghqZcQWzMO3WME+FqqboTc+9ROEZ8shgvm3bQ8k0BHLkrSk
g74uowFCsoc6kvKarjrWAgTBgXyUZz4rj4y0lgtjwIE8T0HGpEUUdam8+NBSF3G6fCGXwTb4Htj/
RWL/ZfLbbN/mLz550PiIvm/sVqRaI0wLZyAE1LcNpALsamPib+ndzVV5Ic4DYVl+uWIYn6jPRR8G
/gPi7mHO6vXtc8kHIjQ8SaAsYlnLsvK4w1TjN57V008+s0pW0u59EckqM1zNTRrK38R/HoOA5xr0
oEPCmsyMKrVg1FReR3nNDnQos5uEmIm8sSzEr3ajeFAvuMeUs7+3J0fzHEaycuURLQDkbZRRsb/+
60bCmb2tNCGJVSECFdgfzHf9IsQZaPCpUQceN6bFq9wmO2ZKjzP78fSAJwGSJ5enOELBPOs5DhAH
dOTA9OORM3UI53V9n5KPa4dpZOWYLjeNngbyrq9V2Ljr7Vj40hEm
`protect end_protected

