

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HUpwfbtoJu5ljZH1PD1nirfZUiqEH4rdOJmHG3byOsiHMKK3LegkCLnxPuPlk+MO+z4ctY9AQVS+
qDXnVNabAA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J5amwDwAOhmwY1AI7aPhS8ck8cUzk3ZbW/PSkoxcoFtS5AuFiIpCT9Eh2Lt0JzHUUKx72jQhC4xP
E8DYUPCIo40JuI++9z5fK4HwpQiCOB47OP9CCbDUXkdRdGgF4e6aIOfD40xCprloxnLZWVs0yawE
2eWpDksVPZ7exWV5yp8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kHeSBUaR4Gb9xyNR7/PmBoZ6gckk9p1h7+VOSSxhgJTOkeDKrcZOdIV1GDgFDrDQ7kzRgTiYYdNg
fXk4UhiKwBVyrTjV2sMzg3+WqoUQIK6Jy3j+rnKZ0FHbaJ/B0H/GfbBoAdHe7Ll2JvXvA2JrUnjB
cZCpVeHDgAOSHC+pzlRSIpPSacSQtQcR7XQ/3XaxnZYRC7uHkv276AbG3wIpLBG2zxIX3ZP+ackQ
pH7/JslwJLo+2yMp03WDL60KY4dKN4/3Cbuq0p9ZXqs2Y5D7OEUZNxyvOtt0dnCx89ZP9OSkU6+U
STforoN1MyOGgJ2YZ3QN/z5I0fk2RYpfEM9JsA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lu2s7AKqknRcUE5f3UmM0sxhb8YGklEChkrpjNpqeFmWrHZVTV653SjxOWSucZRxKRWERgvAD5Ge
f+lfXprxLknFOXVThhIZcoGHsP1dAaIYcRFINHuR+NXvmYc17FBsIljnkMKM4grLGNoBCK5BU3oj
+OpUaEAqYZcR3Ny7rME=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZNNygMQdh+aYmFNm+RRdz6IwBodkqsu7V9fE3BGXF5I2MBgRK6iGinaX8yLwnKR/gy2F4SnWUzqm
SM6Hy+mVD8IIS+xm7ukIVwLbM9+0zez0kJn+qWOW6DSjxPXqHRWy3fQI42FtwyVBs6pb7/W8Q9NM
y83XMjmhW9gbYNHIHq5e9D7ao/9WQ1Ytg4YhUY4H4cSzY2tHj3tbIsVO5Swzs3K1mz8KunAK9qzN
WNyQE7ctUOauX1bPhyKN8vZcKzkl7x8jPe9GO6BDBcCZS9DeY3P2LTqajNPbMa7b+rdlszJkVZWF
aXg8+G+Fp5cfd6qUK77FET8A+G+lv6qs6bNgOw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26160)
`protect data_block
0nUrh8ZQO/5K5hVupgdjxqjE+6lvdNte2oUC2ZVfkJ1QJg1L5GI/zDFn8g5pZt5JC+QeWzith62v
xK48tJwh3/P1gdrMwzErQA9yi4BbGK+q6HGuWE6Xee0ut55mfgRZQtaKYFRBwo3yJMlXCmTZa78V
JJ5R4C2IjxKBYIBQQC9cDY6hDyi7FtJYW1Mo4/LjpgVzncSSH7mJoQpLNxaGuRNFaZwKChJu4YCK
wZxyS0IgZnMBixhuFjTyd45s8VymphJJ7HaYsFKoDBREsZQE53oMq9OgG4EOZYRTppGGobmC1OGY
2VFQG7HJfycqXjasNKg0lgtYL9JFjfrqJdH9gWzG++bX6ilHWqSW3Qah2MrKh4NGKXzhGI/76f86
3XTZqKQs9ZAIIsiDytrgQczW2c29w3coSa5Jzt2qJRFYCpWoWcUV/w2KAzqxk/kbjQ3hIB2QD552
Pu7KJcSER7JLVjPvDT1shJVJmfYgeOopRhLUquzz3XmJqbpkWqFnRsAVyVLeGslVAx74n4wJaRD4
AkLmWhex4uHtv/vSxPYFs/YDAuC3O2oQIx8zXnnEBTzuiXNGSqeKW5gY2EwF8NnerwXhTCfLpMao
3uiiPx+BAwwK0yoqeYeBz64YiHKPguHu2oV9IRCLdbyYVO7n3umti8K7nOgVHrB8YNqRO41uOXDh
vTrP5GB7Qplx6D2otbWg/abqHreXJ2XmEvyaSc/FPDxdp/4zqSybsMNKHEKsGzE4GQ7Dv9VEjj3J
XWpAuh6ko1rb3wW7HTA7eTdFfGFUiVAW9fDgSooxpkjQetOm8rkrfpxxTqIoYGB0q9lPM0wf84wo
jxpnHo0+L6ZCW3rwN1RCQnCOqRRmilZKo5HyIJ1WtIIDLh9JRhK22IxE7iLeLaovjFSHlaHg9rgc
t3FxXIM4Vp1jlWtTzqfXR9hgnUDl1rKR4SPP3BuJQNI0m5vFOL5LaVg6Tx5WDkoCf4kWjnJ7i+xj
TziW6oY3ZYqkcahXpOTjSQV/GCnlfkn0uQutbNXVlnhzlSUs6B3P92YevqM/ukJ22LtUkeJbqF9G
TyLrIT0zXIIV2/NSsAsZYMp5bCVSbJ1JcTb6puK2MsSvX9gqcpeQl5cFMr3V5yHrN9X8oJXZFKag
m7tbde7xljIbYP1Uw2/q83G6o4JSFDmU6F1xRQBh+HXsAmEDK3blVd3e7sRDOE5LIHrrDq5Y49T+
hFajXmkRyM6EHFB978FjoMP5uTFm8I1nGiSmCsw1kQ2TEqaVBv9SosI5v2x0wG3pjVi9yOmVT+6w
1YwFOfPiFF6jRpPQ92aD9C5TanOGLdNC1ekOhfViZCa8aEa+rje0aWx8krWNv31sD5FGTqFpZERk
pHQIfTn9ltpw1IMOmT//PDRG2npfnPCztcwLqA8qCwCW6+7WtKv5AFaCqiPp69AqjSPhJhdvc3FH
iLIJJvbiHU8OzbS3wLTAjz1aAvSPGOcPI3G9GHU1WFHjF9cD9qEHDCV/BAGwE7x0ijcqIstCcPgM
VI4Py1g+AgFbzEP1vge55Jde88Kn4mXVObXd+eRbADw+5GqG4oxhcyUF2XDIedHk+gBvl7csqWQY
71ooarMBJGtEOQxoOtaYFjd32v8DicXmDoovxwzuDfBR78ELSjFL6UOfhetXJtDHLS/7aC67fVlk
YRKJjZ3JqjiwqVn6VKpRvXqWzxRkKLTZoGAPziOheXRV4y6Zh3YoCeFiVAVNzxw43Cxu9n/oLq/f
hmbNFlSVrXkazqgzJY7ZeB5t9eRm7t4vsL3RZJXeJZeHLAvEF4cDBTa1ASV6j5RA/t41Hzejbf70
Vvo2onX5VITypVbr1ufFjdlfDpV+cfOMU1SCqvl+04DOY9Qsg21t4ZOnKMMBZ6pl2aSLAGIPSewD
8+yMFINrn1fOgD+ls/zJ3nNLHmJ+BP2wJwOycMfwjgxOj63F5kQy+ZnGIFeHuR3pVDYMJVKOmWt6
Z33iGvvykc1zERCyccbS1+4E8lCB/DliN5pMSmXDEm1cTNG0mxD+VyA167inrcUQtteh+k1VvPv4
5OrDXPStjQSwYENow+OtBsxCHnmpVZxYNsiYqJpFUH9Q5trVT3qKcEGByT26gmZ3R0fOpD7GDkGZ
xMCyPb01yfiVuiI1rVgzUMwR6UJL0FAO9HlQA0wO5pBgoC7f0mZkVAKoF4jR/40BVxJpTsrExus+
0iwoQR3CB7E5gh1z4iqPbGc6OhESUkOEDJsIRP4qpfn/A8Sq9LeMg8NIT3b9az3FrxviIEYeuBlW
q0996Ue2SGtvn6Q8WSoAVY+dY1nphCWzPoSKO43NTigHTAeqhJD5w+UZkkiCPUCAQ4hxT0urY0vK
YBjuDyxfADvPujYtaoq8shBbgLDwWevE3spkNimXsCyr/aZ+2ndkxD4BxN6a+ov3XNe7b7uu3dIG
lVrN5MDCyTov33qctkIfVlrmMIytF+UFhovEgF8DjczgkngTpxOIvPwzAJ2DUJWCJxXY/xjml+uM
fF9t1cVkf8IV/UbipB0cunM+3HXu6AxAZpjmzIClYgcw+/jSzALmEszfkBW5RVsNz+5NJkU587N8
m/LxtmeAmw8FOPcyhKnnHEqLdFukkomKJbqZBJ7yji79JVZtkdtvGQHc9MBroHG4Vkt0LsBuGJjW
iNB37ndm4tcz5TNElJ9s+tnisZ3PwrWF+RXoWNFpbkN52nfgDy24jKtnJJg1pyjIxeSN18agKE8n
mZbstgfG3UHbRp0JeOCer2X4kj4ai9/B9h+dQZwHFVQ7vKvJGCCtLCs+QMQxhvJrAi91j3xACZiw
QPANNmx1ssUbLAw25HPflk6DwQrzzne3baR4sbbcHrdRFplJroakJXsmb/Ev03YToK6MraSQ5wkL
awIdsLQbPUC3PUCw1SF7uuGvHm6WKxfvqLXE8rABCbjFPaeGFspOV2HeB09BPfpln2aKzIoKPmJo
NiD7JouegYWsp+OI0Ng8SYaYu6HfTR1HtGGjvFRS2vnLOWJ9Y2D+S2+ND8nclsyUQTg4qa3wHBgp
Cw5iMISopNkumdDGAEEkfJpdSJeOh+T1F8KRkuR8wOWbQICby7ZibpkeLVc6x6KQ9J/Xz/2/OSAZ
A84T6LS5hhoPnvTs4m612/ZI170VKy5X08lXAJYOWMgdKfgUI8jE5NLLMB648E9wLT+lr529m1uh
GocHXSVDXhclGhdM+7A/W9Sy9+qAaiyXhroOB2IU+cRInNt4cSTelt92Vyua2qrMPaUzOZer6iNq
qR3QwGLejOE3DDhOUDnH0BUmnmiD5rKMZU0IJDA8BIemkFOgMWsjmWd/ULvlhIE9nDXD5QD1OKqW
EbUojdZy6Wc6tjlJXuUb7lHtewZSqJLWqkP/coGsWaY3+RvEJbZZFwGzT7m7Jm+OSFJWwKCvtmOO
o+KS8TJg4TcTi6ADs1GZ1a5Zr600bdqODzcosbPDxhJBakr9Sf9CEc+uIVAEtgMErb0qHK4EuHhH
tB+ia1ZZWs/kJAc2RuY3a01nFd9KagvSoiTyNKHk+swrp0AhFL35npT4W2OAFTgGgjEmay0odFeJ
vvnze/x2w1TZ8gr+2rEsYfCfKZSCQq7msZpmZAMTfQqxrSssB1Kj9Z16n/j+JOzLosyxeR/7lzPc
8NXFUugWRdWJDrbdrPMUFK1K+WXfvsgjGpMRIt0qRSLLYqDeQI7KSSk+gc+CphnFeWevuvjGIGTO
U7BQdHf7+CWUkps8Dg0DxO2d12jHeybYG968O2bBMbrHW52aldzdDISamqJvIefwanR5fwnJa/P+
Z5hiXVlI2uPquPVgJ/st06AiyO5PsyBdimJ13xCk4zf73ai7lGzTDstjVGYi7aDEUtpEVFZqyMXa
YozpDRArGpEobIK1XXGwCEY+nThPNH/QZQ1p/CumQOPVS++lbzJ7EZrodZoKFFyaorpyZbGkrnG+
g3KXev6mSCEMCaYdQwNf/9BHJ6uUc04ObY6xN8ODdDYtmbwghi0IOU6jLZ2a2s5CZLnYm2dqNFLt
KXuv9kiu/QqKavCzwFkFuF0R39LeClNOQnDd/Wjhj22anclch0dMHm7GdA1Xy2kt8wNyR/WPloRO
oR5KH+netM1VoBNAtx4wP/qgZiQP+t+TtxzhJRxh54UWKRbJRTCUSVgg7lU+N0pNQi6okZL1ax3X
ZHopjz7ZCWWBhw2hDGXIt+S3F4Veinbv2FUquNBKepprZ5lgfuE4qsf4RZJAJNwh0KXb9+En0+bt
S4v4uM/xfEezTsAjlqVL1LJ8tG3J/TyMnRcCylsC7LSQbzZzCUqKy4XX9PxpXM08DWtSwOsKU91N
WWLyT/WVuJBC1oZagNSmx0emNdmd5GfJLhY/ma7nfI6tCcdSPhUcuTHOBOzt7LUpRXMDz79RnifU
lj8oJhE6c2h2PHuzt+2Hz1CNgw/wh2bFzc7DotISqxAiqs0JvUGzKLAj+VA4DteVjK8nDgRJx2j0
pD13pl6sw5mpPQWdToltGdcXKq97cVJHPWkrgUhuXhez3jJlqwvPa3Nokl9J1ZcNFU1BnDmm6sZP
2yl39Vd1tcp9LOLmRk26oeeynctBJQOymvopHrVWau1k/Dhe63r09CBKFJoX0eSZIV9sMz9bH42F
WGIk+8uCBdCBcGxTfGE/yCc3wunhP0xj5HMK1/RSxWjZKSye6rOVKEwYlOqRSDntsMW5Dpv6blUc
udhISZZBOqFXrOq5/cZ0cn/C5D/yThsZSKmolNL8+GhFdkTnyRHpibE1M0bbZdJxMarv4fiUfYD1
fTN5exU+nIf6qICCTRLVinFbzH5kvhuGLoWDlI5XCBGXOcDPRE+FuFXOgGCmgwtaIi4WDL3pGGDg
oQd/xNGyUXwhrlPkxHbFIwBc2/AOpNCKUaEK7l9qzQH7uquceDuJxHmj9wh/HtQdTySNpZQKe7At
Neh8k9p9ipQlYePhgUpeoY4YrdRe5BzGGRpx+gqwdd4T7W652TZsJ498ItOFqdoClyb1NSz+m/8l
WmyPAzgmdxnMVjiu2kJXCCd2hkUxPanKIaeSwUoVW4MF91XFzhpLIVW3ZQcPdCblpfNgvs2Xx9Qe
HoKgaMDeFVIeXK+JTtFWbrB/7YfluTsFAmJRDO8vESZUZfEs/ylm3Xk+4I6276PQ8/L+ZGAoH+zt
wRFCQLpTHtn3DwJdglxhJZBP7XyWJpVIF0ptSM3dEpBLGh9DJ2sLyz6Npi35O741nxDNAHIqb2kS
fHW5vfzRPiGnWJ/ZciDKwXoPKOuw+17r0A67tuH1+w3LR6h7lGEVSqGDDJkENuXEqGjnQd/OmIrh
t3OpdPiRt7prrCrpTk3yJEK7TcQUfjv8azvrcRqZSJtHvdI4aydt2YH3QpazhXrv30noIrDwjuEa
SZ2hCl/r305bl7x94dFziaqRy1VrZj+sMTskXdspBvDPbPB2gRUVo+nOLQ9NLq4IEXkcpa4hfRBG
r2YbPmmxdTD1zheXC8fv2NeaqcFOPVdmWte3M+48CLtawnnk/auPVhl7aDrEA1+IKmSotTPNh8yI
OKgXybzlTqpvtp8ZFEQmfBhOXHnNvxiGizDKhk9HYyBKpH+Lr75Je6eUJ18G9Px1sTzRVeqnQkec
5Mo1O39M48dX4GBEIua9CA+VZ+CQ3o25FR0aog3V7VbWEynxGdnE3w2k4Z2LpAQpQK1Dt1GZMQOy
NsRGCRGk9M5cfvCrjL+H9JnP2qi1+50MaDFb3R75qcvO/3Mo7ZUM7pQOVc7GGF0Fdam9KV5rUk6h
MpfgGAS8ZOYNvLh060pf/tvSnXGfgwrY9CaH/i5FbHyKDt7qIB4/90oMWTjw6+5+dOHJgBlSZBi0
ZOrlkgIXusSybfZDOajyVH2F58//8/KtpEP+IqQehWxx5dv7QHDR21/stVety/VFUBK/P7x3v68c
M2FJ5fNtyJZY3PyVJ9VKR1t90Hf4fub983nsjAudyWrjFBd7vH1+Aoc3KFHvDzEwZnyBBcesiD6R
fECpNWMSZjxPSlFZkLR6rDctgFlh2CYkiW2lVbNYjCfG7EcQfJgCfC3dfyfLa736RH194kjGy6sF
XWCL+jeQB7U9AmUgQ+nPBnZB02sJQBgBX7FQdXWJHSA+LAsP7bFWbtfUEocH6knTPhrbDVRflNSc
Gfi0fZ8yJU5PCSNdXX0FGu/XHJYMmfJ2OE62x/OeY71Wjo8JpqZCt2cXPD+kwxh09pIUiTFEU4tL
ATG92eXIcN2Lqg1FS6okVE95mJ0pZNJBOqWIdv02Qmqe5FbK0rK65rA+/Nu8neDd2TGrgTLGMkJ0
BRMrPE3W5W2pmQGHkfD+VUldKLPa6yHi5sbzyu6R25miKIppFeK67Xu71qZJns0oAXMk9jRacE70
tbBPYFCcp572uiOUwdOxal+U7adekcgqRG9jhqLpmLMH3855CYw3BjDx42TnQEm6k1oA1bt9QG9Y
T5N97dmaiLXDmob22FXGOOF0XGRfi49XC80dI61xlSdFwUvfNE/PS86NamP55PYGLxolq6Yuf2+d
Hrhs8EUX3hPve6oMCobpqd3IZMNuvJQGEqrpSqGlzdl8rpDRb/F/EDmQNWeV3ohB8RQW5iBGLPQB
Cq/HW+dbNGhI/kvpiRCW13Hv0PY4al/ZSuEZMKS8up50KI9mcB8mK9yn17SO5zeAhTFQTmYe0uG8
StUKETk5F2JO3KbijpOkB6H0mEuvbCBoQOkxeApShgEi75wnyL5Izhbo18zF7zJ7iqFnH9OiFrHh
1NgWjwnnhvjXWBw/mHU5VHrzqnj4YcjOW03SRUARHWaEUmckQGVK6aRIfDS8HxY/IkosIP6mXPd1
eVnDV/2IFyj1P+J3GgpaMLzOkqktiWh4r2bLzVNWUUXS+paV7QpG4jJ2bgtdbXYZS+xBWPJFXpVk
W6pumjofut8iSzqD67kjvl4XX8zR78GlZluhCc15d5JuVVdCE9xcRnMfzpAXbuvTzTyKFcw2CYj3
JR2rI/d/lBPirfOdk5eWxunWzXpS2nFjN/c554/1sFgGDL84hEFykuSXxIBWPFRnoJLas4/5PIaQ
tQUN+lc4s2pjB2whchWuwVoeoCzJmtEvqq3KbuTWrB4qQfdMWaFVpSEeijZSCFgAMuG7bbNM6+Y5
BC2mFWeum3T/P49qtMgoGyEaa/+Pg1ie43uVNCrqfWEJHqJ30hwr+z3VwSR4isL9VAY5GYqDt69m
zC/w5bx/NUqo8yXqStJVv3zkzmgAPr72uxr0veUhUi4KEkD145aY3Wfsblx7W9kMmXejxbvrpceP
D0sEkPx2rUSOt+ceznbooT1++J4ELhnezYwsGMX1rvZK6ZS1GVgd1cRIW0ETzy5MKRc8/kX7BJu5
KFhOGJsxTvrZwlzSM6y8AxDg1628b+nh1cJ3Fo+Xo3wgl7GH8CXkAGphDEDgLKxHTHfcw7DpfRCH
Pn+EdBfDAuR0gYhjqjzhiSi3ocmVCLpd+prsK8DxSS672g2W/fA2Egu5XYTRHqt3R+mCbwAvRYD3
+nC0ZQBqt3/8qYBiaHWKLwoVP+tWKkryOLMoZjNSl0844jQo8JY6tCOZhFhG282Ep9HJf/HBFXO/
7cVQMCLBsMre1qHNp/2Z5HmMHhvvfckNkbDYiqezShSerOB/PLHO1OCm9nIjip6IeOKMF8VGi6zp
1xDP2+bw08n1bD7g4A0giJT2s4xW8WcDM/RALppsAqu49USNaVcL1/+ITSs7pjo0va1GWGvNDhkR
P4dIbA6OLf4lyf97HD86nlTo3osXGQHtF794S5Qzm/OQbKZuz7yXu1CRh6c6h2hgYiTwx63dj2/f
ZLbGB2Aan0ndFwDndA+ZppKmY3u3bhTlhinWNSmlz85s2NEwVW4C7MJJM6rYQhQ0xqQhd3K6HMuf
YU4jUByoATIGqDYAsqjTfeoFRvuVR1a/yZwBCKjH1HiCIFqKv1asYpBFvUHLzzqAykoLr7lGpfl3
jHmhdrJ4e8DK0AJNrTsWyOMaWUZPRC77N+WLmRdeIeO0ARMFmLxvzv5McWZBK3EjLpKXXO4N7IIm
/WD06jFx+WgQ/vug8M6Z4zGAJJsVO14tnth6WQAzBo8R3HlX0BtZkGjalnUqHQ5k0d5oGBAOniu8
4tRdSo9SwPhcXvJgbN6Rk0aqRr6Ps/4/9q/HF7E9jD9MxZfHB/x/jh8l/m+/3xitXuwxJLbBLaQE
hYjAqKytM5wn5ZTiEiaUeSsBSOK9l1twdHt5STVUE+oqIF7+pZ9XVad5bovBzg6vmnPJ5vP2eC0B
cUpSuv65Dy2jRgsA9+Tt8fJQuF14k4utBTRgrto/9xTt3zNe9d/mKraC2vvI7Ex4ZFPupecCrG5j
hrMa2qF6m4s/r10aUdnRYBA8bIwJffUdjJyB0NPaIyGXnPeChV6z4jJWVS+xoZu2c5vtAu+eVtTW
1qjdjokwXIBtY9iFfB865D9z1lHtoiyWFMX31dKnVq9Xsxzl9WxVV/Cmg3PnViCfkBQZVqs5fiH2
Fk7rYCyVia6kPp0nzTZV+tw1d54OWjpHNh7X2cXzHej++A1m4Ym1A5RGbglUdDGpnvmNFzo9pY1j
Vg7dBPS/gqnPFL3Vd8fMlEFV/zHl7GR5VZJi5KQyhwz4PSUgJmWVEPO2ee3C7QE7Mr7EHEKx2yoR
u+j4nlgAD5iTgC6BSog1Wyds2ugF0Hx1V5lk9Tq+iHNdbOtYiWVGKqmoFBxNNmjoHtkRlOu1St7S
RVOKRwBekNR13D7Ro4QmHKuT+R3jO/reVqJaGaH9hjNznD1r/SS/PkrLzxCKlQG799948OYfzgWF
Xix4PFl7aa5vJOY1OvmAr7/0pQKtNCI2a791oBjEBy+oP1cT93kPs2r4Bbo854mCGHB/+JF3yHGi
B7d5pQSS0nweuU+UZa1jTk/JqBAx21BR9GQgZBBPBsvHu/DLTQpyA6DV1ooqQXAazD7+HFXvO4xV
8JYXZaCcFZ1CMPm2daXJlWmehmhHk374A8JFeLTWyCUAFGcmEf1nrJQUUZefSuXF8moGgh4D4kI3
tjq5eNUoRRVmhK02bsqmw4JqpamsgHAD1od12BgHfwmXeehPNUci6aJa+PJrvXy4y5xjjRKKurWz
nMueNcYlYpXz8kLmj+v3u9mmCuFpwKt4IgyMWkKEn1XnL7HxiVCtuE1mTqZ3RbMaQStACDy8j/VE
LvILd/7nTgUy++uaWjWszRa2W1XRuZ9b+XkXXm7YUM0XhHpYIg+bZNkQf3WaWA94pK8QBIv97giz
2vgYeJU/gjHPAgoRpeig+zOcVgQxkF23cjS60cx6z7YXQpuzMOYdNrPFK+a42u1kMxEClAU72XmW
Iba6nSNM47XNlKzmEM/1Z6HSfXQhWplunuctG977pzlPGEtmhlajy+Llx6n+2qWcmOzz6DE2bpBN
DjIqiOpq5aT+2Yu9nvkRWlvRKU27/Q9g8SGlIMvnWpBQU+RWugRqFk7KgCEMgx1YsKrQ3KN0awKn
kO2xpKd9KZmd7lbtJESpc6OIs0kGnWaBwqUDoDUt26NuRKirmjyF7f4THgHVXduK3hfEu2h4viSD
IFId6De0xwYZwFt2vq9o1Gux18yzTP+8rQcHhSAnqTTQ0RljHjd+Duv6rGztyJ2/FuvbcLcEkxSY
f+dmkGPC7wj9NDj2dFpFWjNZ78t7BBV7rL8U4q1jesWJRN9riZQdeqVbJplzNXHdIwcgOXSXgVGe
wRBVKdIHHerW/wGY5vvSG9NDAH6zEwS7KMSTSQNbnYTkopzo/nYAA3l5jaUxJWvPKAxJMEfU0QFb
6vIbYAG4UIQd0u1zmSpILsW4kFE1qEqPgokFsTi6EcwFt7EvoFv6x03Ofz05LGWK53vBZe0mkdXi
rCy73ulZ/txEl/D8fIFs274lVtLwA5KVfY4G2UTgpbEvGn2T3BQbGJ84ofDASy6G3m62qFMIyda+
MKKtqnJ9v2bkk45LT9ieP3PQ84cp8F3MgXEOBiVz+hV1btcwbO2ryOAKMp3rbjXdx3xlm5nxltGA
0oGe57VGKjXJmB+/rtE+Fv2fOfmwQi4l1cNRRhhjvi8QV8ldxoGOACPtO/Lsw3SGYtF/bOBY3jJz
p4zfzOwxuv6qN3AyWlzDnK/YRlIH54HrZl9MoAPRQFGMJE6KYR3FJUJ1cEXo3ue1KjOmDqSoprIf
cvrFpkaY+kLQ5P9qgC05F1o5BaGUiEX8cvWQHMj+eztV8neq5e7tIehKC3uCoWo6BTjA08VeVjDT
mnykIbnaibLRY/FNU7met1spg2ah7WdRBYspSaRE06tOQOqJ3STGV/KsDzFtN5hATbj07oE7Q77k
zyszOJzKL2vhjJqclP0M1oXDJ7hE3upOj3gMbqxTpfZ+1d3Uyc37pI0u+utthbhQU8jWx18dNcCp
BDU0TiYwb0rRdBHi4T0V9rgOkwc23Xt0IVe3jIaLsviJqjvuSe3gX0t/VJaaYuJ27ZLh9wla7SB9
LOncZesSri4aZj/kt5olANzWRxbN95l4hgR3i/MNxa03LJX+jYMPl4qwzLiBXIFSbYpnyhuwjLQQ
scgEWJY4klOd8Vlay+kS7x2TrKTCOJATx8KIFziGZVyyibgXpRDQGz1eLAU1GCuwDNMS8boNJ2YZ
HBr0I8fukZzWFKFTbB5U96/9YMZ1ne1iTWG9LQjFYjDd0Igzz4K7i+n/jdBpWpWlRub9VqJhfY6x
2ZdgREl1KoGR2g3TILuNDh16EB/LddYv9WOz/vI6cybDcZbVuzCu8gfsT4FlYXvp70g6MK89bsDV
UxM75e4BM9D2rofMd1iZOMPBbZZPwpO1hDxtsqzzKz570dNPtz90Axr49OGjwgSlnHbgpYheSfwI
qyH5s6G9amTXNeYnrYTqubna0mKIG044AI0/RClJ8hxKdzo9uzfDiP9CVNtAHo8BzoLg5+LWr+Gp
pkCThjSxAL+ZCwOjhrq3ZDw12D5UcPvx9JE9YbxT/Sq+z5XRdybCVgv23dGAj9YfDnRzGGbYfT25
QXzks8XybY6qyPPzP6JQCGDDahZdZvmOkee4CQWiQiE4ef2OCpgVtwuw/Vc6ClNBKlv1qIOYEBcF
Juhn7D8M934S+QbZFU0Nk9qHbmiVs3lHayxlS1SYgRsGSJi7Cl56vXiHOY9C6npb0jSmoU2Hcv3V
5bbZ28HYAfJMHFN0qQFJou/OXaMcR2UB/D2B7vgBUajsYd6Tg1Ri9abqwlZr6GXtIYj0m6ALrrc/
PCusbXIoWm6xBkDM7YzkNKpEXOJuAZEThl1Ef2iQYxFppJMoNJZvJhTzqhZx2MkwyzBKLU6AVWD8
3memEkQ84ZEVOCC7/xQvuSvStc3UnZujFpjaOO9u/bPSmrUct4uAO9FociqJs6cDvWyCvoGuaU0A
7ZfE8DrfT5C8PZEx5qwGcyhMZeLOluEUGakeT7J/ouNenIpJIg9rcao4NGlU6F/kXn8Y+NJ9AKmX
WYlaHtZCpywBTtfVKh8pleI6TVfj1WtI3nHL80qhh6wvP0O06d2HIPaYTQm5J3ka5mHJMzyVay5b
Idw7WIP6538KhEwEyzingyZbkcU0B1lwjYIPZrJDuHY1/otK6+Py0zIjc2pGHZ771Xet4TpLT1IG
o5ft7Tz+r5z9t09QW6lJtDD3hphoUVY6z9/Gvk11gsytncNpWKawqUJQCZ+ZQPUnMkByZZRs3BKT
6YCrN9n06+cBq0rxIorIqX05ppCowJG59+crCAh/nkbFGd2Meq13PZ8D58zwAL6oOHuoaDzI0VE2
66GgKBt7e+L2aZPYyCiQGkbypYHn+S5sPw+oGgewafncS10DXG8kWz5DCX99Mr/2L4N8P9UkrmeL
gNZ8dUAhA0rzme6r9KgTebknVgmZ8sP9W8sPyChRw96Kqb2mrb7VMkHf/vAzKyDlXtmZ0kZeDyzy
5NaGt4kD+Ot3PilIdZ4BML8kPbvBmuAPuIOYkZWTp+f0KuVi7GvU6BFsw1kYhy/Y7SeJi/xJlZxh
P5FiSYGvhmHS06nVy2blCyJFkngT+Dyzali9IgGOPjkZVy8Z6IC8PpxtsoGd1nJRNm6aD4Ts7mUc
WvVXyO6GUzuEMcaKhOUSJuo7WKbgCdP68ITwCSE6tEmc2KV9hAwKxfCMxUTVRSrcc+7RwEfmYSeK
xnU9hlgP6aLBgAcNHnLSPQoFTcYxto7JlGgQChlAsZdhREsAwxl8e4pW7IKJXr7l+gM8ZwKxLYRM
Wrxahc062VgNJQy5DAibK2l164Ma0NY/eIrBDNigEJIlvhuBRb4T4aBJDDakGg6VqQJcWvsKrxqW
pR3JK4qabKAW8He2cFa0F34AN9dHTc33SlAKAd9IKO3BQ4lD0MDC376xXhvoUw2yI02BcplNGGRF
PPxuCIceiyYEaatuUkaUDs0Hf0qUZulrJFGqa82FmHMHxaknWoGsLro0H/smLwOOm7F/V7226hDP
13KV8Ac5jPkqUfTsXv6+nofMMGueIKeM8Wo2ap/3O9QTD2O+80TaCChBLEiBgEUX0bjJAq3RlzUK
pHn/Xd5/KAMhH6f4MWJPQ1ePuRcpLLcw5fb80Mls+lznTXTs1JAGAYBxR21rRNObKW8xFP1QYODa
nGyhStzEsfHVkRncBhQpUF1TKODWy4dTC1NQbJGRaVc6/invPFdeww98zZPZ2PBD2xOvFXIBNHk4
dTaoOwcwcHRhk+JnWm6pMS95GJcmjRsfnNhV2FPRDsG/3H+07lUxXiIsBZb4w0BuEKyw+qy0Z/zG
NJNQaHmbvwF9M0tcZPGrEhvepitYQuiIlcRWhdsdZXQ86xMCwWIJnpjyICz8Q4iOsQsZalWmDYhE
F1kEHZ+9wJXo++aESioNyknS4TQLIlCXgRz847PYl2tjRkNGgIBFG1w3/Is+ykIwtBIxVWp+F9mk
WmLjhKNlujPZIIJw+ZfgMM7kT3aPbsB8RusXMdu4P+qkguFEC7zS1pc68Lp52P8iPLPTlFTN3wjt
tbUbYreYomw3SpJUU/8rXhmnGq7NXIiMJAX4pha5lgsglVMGm6LBsbYcFnP+0B8/4qlxtuHUr8K8
hUWZ+LLLKYJQROBrvEyR/y5/lnQQ0k+KfbU3vV2OYrtdVBnwNPSuC683EYHOosX6FKRJDblHyyQN
a9wBh5Aw+WA2qA1VCrO7XOlnY6wQUCzf2eggj9T8efGPaM9XDjoZPOsgIVBtxctRTRDWq/TVKlIV
u9atNX0xi+Z/N5lUD4cLy7alk5zS+1P5A/jTOnwGnHCewAHN3manvzMhWGXVjz0VLe9OX8DSszD5
XJtmzqjXqloocQyM58iFBgHNyqW171Vz5beoYA/0kZMsIOJkN95NSb2SyjGggfZz+7Ncj6yzf+To
6McGwMV9t9vkaMjhMCorHIeDHRKYfJnoHPHGwfhrPwqhOi5oeXhfMzr99vJrbBV2q1IrIDBBhgsH
/oGsc4f1iASchj2oSJ3hYi/PVJoY4lPAXaaGNfaCNOmwApItKYVclJNctuscVzJQDN8iMfE04Trx
Wr3WmDrtOqM5YU3hSjH5V8+jUirW2QuwinspD8ERKiKw8JiEyK5xGxEw9Ba3oJC94IGGjA5i8X/J
kCM4ef4IUoH0qbJM4TOQUkxJe/yLb8WxvbjgnBjqi0KXm53YZflhgP+c1E7t+r8vGw3uBgZMh1pN
eM/9xr26AoHwVK5c4KFU3Jb1BFWQPTMz1DUXi+J3hnMQBIYkE7M/hEDjt9sQ/y1h2w2UA624lx2l
uqxaihB7p/toqFKbOJsj9lfANn2kz8Er2PGUbXwnhbmuLdkljhjknX2TAcThk8W+q0f4tz25koDN
nDEZB9lwyzfCENZ+vEFqrRaqp3GsDAOdtCGjfglyjx5NNE+7guW8M0/xRyuJ/2PWPlABRgFBUl52
jfnA5Ny5Lmi3MQZEA4/f8S5Hb6WzwoKEcbaMmOvD86YVZoyzgZurYFwfTJ1Hr69O7K5orQ9TgDF9
xCxlOu3ilc8W7I3dPcpKIU3ucV43JVe1JUXYiQQB0vDhTVwf7FZFaVgjy7RTGHOc9YNOYpiTUopW
4z7tK0qt9Oet3hHdAJilTVZZKkUghoJzZahUkvwG+feJx7sDk3xjot9jQ8ylSUFx23/ZdxBgV6lB
d5f9I760BhJ3c70xcuvudUFsKXH//TWhZy5hW2i+Gr64hDqCJvw9TETvCfR2wUxOzhDduGoeBE9a
oZpnyeOcNak0TdRQDSgCr3fJSD/k/TWoBVfPBCEWO1N8lmNHxmzMTtj9IA3G/yJS/aJgb5dk218P
612cU5wMWguaJtj60qNdJBQyuatEXcbkqbjSmzgvLsqfZDgODrIjEOys7EoXe4Tk/LtsDXLGr0oz
sDIuwY7AxMZGFKAqf76dCkxFp5GsJnktyC5i2SQ0lJGsPlQtGmkbGZADRL/YZu7nkDhqT6f1k5Qz
u0hkLRO1NHt+TfxXFf+4Xw/dNqmjSeq47jiLBNT04LhLE+ijx4PH87+j30/Dtl9dc8d6JCp5f3Gv
22Rxw1JHZnxmByZ9/lWOvQIoc3FYb5b45G7XRnQTV3OdhLJeIkm/SVo3RYKnK35FK6q00Tc4Ti2E
yJoMYwG1EuILnWJbvsIf8vLC4AJ1xjhcmma4Z8wJYRC2jejO05eeVfGH5zytch5979zY+WlQj6zl
zb/SWokWktUIhaixqhTJPxaLE4M/IhMh1jOeRceLJW6hzq+PCzH930UQQhBtNhfAXpEE2oSkBar1
XlKdEXM7Be2dOgwzUpm0OQjVkkWVaNTR5IoduBvVUspQxLaqP2xOjuOpsQu1g4QsDNNdmWgsN8R3
px83ot6Qn+SxQLUd+URa3dyaRDrV9bUceLfRdOOkNu0guMsSNP81+BJNQU4PaD0mH73bMZeKyJgB
b5eGXHwMNOBseyHIFG1Hh5pj143M6gRY7GSDWmYDMd7glEEJD1la7VS04I4yxuKUc08AOEWIKIOd
Fl7XvG63mzgUyK8rdk1nE49CiyXNcKreR50+reXiPyavyWS3CPPt0ZERzpTpI+wRZQylRlHfsUyu
qh+S2PcVWTj6iyFqMLnc4ovYF19mmx3TNiet41Nx4Svl9iVSDQLYPcQS8qHK33XT+jZZRb+HfGEn
0fK59ZeCxDfMQxa7E5ZzfuY0mZT7KkSrUsgWDMnJ3+C1hOX0bxP+0FPl3SiZhIa2Nu2tTKYCtF9q
ar88RNAhqPGdvyR+5iVAa+aFZzfWzsloYcmYWm5sFVBJdEwbetTCI1rv2Iu+xN6ZQ0QGA0CI1FoH
gr+8ZYOOifu6jDgK+OMWEaxyvCIdbivN+G1goP9UmH0XnsD3zkl6LH9Jgu5OurB4HZ2Qv7sMo9QI
oDRXJMndBpKHxrPWZ3nkdFXLUBXz8PDPjWbcv9sU6fxEJSd9eZwxpMwsjhEFVyXK8+KW6tAFCLpn
mOW9TMDIVSjwis5Oy/JuaF/YEfvVSjipN8GCT2zXZ6iRr5Dp8PSavApFXGelNFVX4/+S0tWb53E4
V+w5Ka7dLXklF+BE8p5XV9RtZf4nCx2mJJcy3K6Q520NnOyjvVPjajDGUeronHd1YPVCl52vt5ry
c4vifaOlAu1aGb18MZtUJ42TFT6LGSxZ06mqOyIowjMM6Ibak0d4AB8YxTqmmzRXElZkiB1GmrNO
eVaUSgbe3efoY0H7dcR4UL+xo9OR3LLCNb3SGgWPjeDHaOO5krgnOVlhSTyAw99lq0dDbtUiflfp
tqj2gi9XJLziRitmKA+RgKfB+cFg4A5uiYZvzJriv9N/LgMGDSe7+ZgUNa5XDSPrZPEAwbIlTvQX
SAkpn80TLqcajqXl2tIdvM4nE8X7+m1KCsVxdEArfVVfiH2xsuQk2xERVYsr7/09L4/Y9NuWWeSr
EPyO3DNxq0Md04Nj3K+3L8AS1rcdlYcBUJbUX1WNanqB4y1aC2o0iIuhij4NH6MxRrTB7QDPfQ9Q
IIYE2Skw8pH1hweyj14jVrBGxulWjGY2T+eZcK+ArhK8frdNG3SHpyrt+jEbtVjYnUdjdMS6L+50
UrOXQzW84B/2YsuT64e73+yHsL1VSKSnFHqIPfogv+8lMpw2q4RURLiV08ki4QIQ2R4Z6msfH93W
Bhn+j5BuK6hYoYKagelPZmig901X+gBSABABeRsXNoQzWagZHKEXKabo+lh44PsioysfFeu9ZVZ4
tUxVOXan/4wn1QFP7IZDO2B30Vy5YijvpS04XCg1F7iPz0ZeDLSv+nMAWlnoyiW239JgUIy0KQNO
AP93GYFyZxosJLcNl0J6eQ1ZFX2uAs8Q3iilvvKkrUV0Ek4FOdwBaakXmWqpqRtcvADeOPloNoDW
farUxfgSHN1V0ZvseRDUZWDjo2Pssyf9IBIC2NnOJQixjJs4P7IGJsVSvw9/f1ssiQ4qdmK5bOIk
YvXEWaAzMfEg2Dl37etCRdaY6kS2VI1ELBUtBY+ohl4MnTX4A1dvf84+JyRqUdZJSQo8q29X2i0g
TcsIahB+EAARruqu7sjUtjwvMqxwFifEZuekSD+yeJ8Oz6E8TPdq6xoT6nhPLuP454rqh5b685XI
1q5xjucMBFo7IiWHuAnTyaYxqFJjIELTlFAM0eMTyLftQNv4/h23k3XqNQ89RaDbE4/n4SyvP9Kl
X/NrfU3F3A86mOkBEo4jMDf4TuGJ5VM78Xv72rLTA/u6EfhpLp7dnBWZOqh1oGT7KNvi4QLwmScZ
y+EZfWT4UAg3FZtQPEyULDKBA0uKsJ46ZLNmI1P2qtv2QKIt1YKG4/fwjpMmcogcCulMdd3aS9aJ
15l8GXolDxMNY1D6FDEtYidYRMS5RHgorjfd0alcLSURf/npr8JFHamrGbtwSkQjoSO+OunJAh83
L4NCXh02JX9s8sKVltrm3CkGvvHOY8tDSGj+cEyMBO30hZnCRWgKObKrNfrzQOi/qY9++kF3pOik
Gy85qE4fWCMP+TIpNUN644pXyO/phukpigkjHvPDtKR/Cxhpi2LC189EKoLR9l0FZISWc/4SUzTe
GTA2lh5Zf2u47SiqCpk4REOnD1cg8o8FiVjck0eHwF2Njlob05OSXl7k1iJzbMOsn0oPP5RiYAdo
40nY8B+o7OgXPZlCPmKX31ltgjDlsR8vUiMN/hPLepmBL8X0lP8s1hwVe8eOOe6zpkKyhV36mNse
wxH1cBX23rzCvvMRDfrf47DGj5M/I7vqBymSu2rCXs782161E/c3WpCtUqQbpzYQzT6FtuW15flg
TTDaTccnLVUvBF5TSRX0uLUWaSLUWHhcglr78ZkJ9m+yG3NM4SE5Bf/lzcVDBWEfIYfzjc103mYH
QPTSy8t6rObvUua5Q8FxwhMN87QW4SjfSTj2qzot/FDrn9KSt8L+9Zzw3a1VKsaD/lBlqtirj75Y
u9R/pPMb9MxkoA1Mnlbj1kU/WXz3Oq64eWqOvqQdc0q3jahxP2sD9fOoOJWBGYHiOF7T1FjmXNsU
E2fb14tC+6S0CUaxZmUSFphfL263LqBV2qdbcf12D4XebGcCiTlOskeqNib3N8GOm70gdG6rLsfn
/zHwgKcwyFbmTYoagUUx0JQZn6NsJkVxXrzBVLB82H1r2Fkh3DGZLPGs31vR6jTTqSkP0Jgl6KQ0
uU2cSoBgajIFVBCTJ+5jTVPavIRLS5ota8yjkvb/p6CofhqyLSWKt+dxJZ8bLpoZ/CPM+lcKKZ8B
GX4KbbOl4r3W12AWTunz9mkLPBDsDQ7DrIRlyEMGweiO+9yspBDERefAWeQkUFPxz+NZRkD29Wmp
rUx+hmEJAlAj4rdcJJC1FugP7hoeWN9kqCeikivCtOj62pfS3JdHxtyJ5BdY8sIvsLey5fTC3EA9
udFLpcrieGJc9Jl2QpNp5a1BTmEsi/IVyfyqQe7PgySBmMs7LCbZu9quTK8IRLr/FYnzTKyy3991
VLbjLAIUxFZG1JxD8GLXOJHFYh+UHiABtFT/2H2Hv6UdJZ99FHO0UFWkaiLaFLy5HoWhE5joD2wS
axMwra/52WWlE0WdLDjr9DDGimLaag+D9sD/GIf+CfBoQn9JLuBstVyVGqKPBA+r1NLq6DDKi1vR
hAIsoN2bOUSZq/Aic6kurEcZUG+7574umbCmaoo3r8AMjO+mO0VkGEi4esd/BZoy7q87wl2tOivF
mxUUuHhUFI2/pJZ5Y+X0f/Aj+hulbUqA+VuF0+LVqgPRIp5Mbt0yCN4fZGik27TrvRjYtxLUWAZL
x/1HWPfXiOeZJWRTCyk2xeUQ9b3AyvMQYATWagjdQJ2MsnR8fBTLjttj0hRdhfi73/XweGbCeZPQ
VpcRVEk70ps3mlnphIlda6nSFDGOAFTAgUKFS5vUgxkYHDfzr9QPDh1hwf8p6SZt3GiZFImEuPXn
oe9VqRUMKefWoB+PexHFOGhSYH7REspjG+1CO9IYniEkL3i7m64svJvl0psTlq8/MwmLQf72bsQ+
VllmDhJINOQBM8y9+kKZv4amIXPhuwYYeVtnh65F0Wv+Am5lF/9RfN4UykKwGaFLEbI8ksPhN633
Dd7+fSl6ts8RdlFi2AGITA8EfOoihvDV+/GYcsSDD9dpyJ2rNaCh3X82wlpm8OmLof6t0ifHIZLW
UCU4fMkZh83tCwugoH8wfCsjQ+0skTt4Y3s1M8+F5dt1x6j33sJFCpjFfuqmIrIpZPGtxJIvEzEd
LbLPPbxKRQboxnhiqDJNHoF8n7fRQfx+9dv4iXgo+KFejJRgP9qWs+HxlNbc6thuXVPNcKbJhE66
c5oXKMIxEPxvJfbDs3S0wHQuew1a3+CeuzJlrgqERXoeSh60K9JPNzACgiJB7pN6DkGlV6vTlmXc
7eIKn4S3HmG/hMYMkQ2AtKCTFDoXO/l5zfnkUoAvB0n1M/8lhpaw/yfr+Y4S/IfLsj8kmE53x8Cv
DcEp5iy9BSo8GstK+UQrz3ksS69N0adtoU70Tg9w+Df2orRr5ntXLDxEJ+32kdViiS5ZnAOfHzXu
8cN7a8GfeABgONGUMyOHQBRsbCN/jKlr6oWIi0X+oatSnGfGOV3FLS6GSiYsjbfnDPKV9AohYPH0
ai7JJ6KkjVYjSQhezlbVeNV5ORVFvB/XHNfHcyWgLtpmx9LtJ9aH+iYgvq8MkGxO/baM0hPUrjel
EscvV+88dtjb82/yLXCiJeZZwrh9FRI1SIf4dLPX+0WJbqpsQ7CArydplCaFHh0FfCVGwYpBa4i4
iGYsXrHC1+PPIqrGiu4yVBh/GyiLQ6E29ZVURoThvkRmaVW4G3hXcfI+MZ960B1xZPR/Pb63LXDq
+j5ayxycpTEus3oZEdD0PvPla3UPrj3FsmypwhEipHEl+DcsST7qY6kIAbL3NBfU/7snC6cz3sgR
S8jXsPLMWkWIDb33FdMkrTm0R3g3mQsiyL1eJkuF0B3otKM8zCDUVxzvAR9uxaNb7NDIVU5I2qVv
VocShiHQ07c01QnyJU64/rJyVgR8uLhvFYEh2p7NPZfY2M1ES8Q0VaaLoPaa7XIa3lk2aAg1cWAG
eecqAQ1kGbqUY8REiBUmS4MmO3LNGzFjX2cM8yhBuwYrHhtEpOuDgQIBVFL41qIVll0eakSQpVtc
tLp1KeHQR3tVSynlby9Wr+p3VP2kYH57ZmXJxXvD88hJZky4Ux2Ny00DAvNjmtn9GEa8ysUQsdXo
XbqWzmkiQbEBO/PzkFuEEj/sonS8Z1ZkIw/H9eITIbRjsnhkqXNggbEWX9CfxHF+4q3LmOWROlWO
jyq7+LGItEkrxGDTzsUdP2bnidwcn8w3cmE73e9Q+7JJ4MXkmFLFSPgV0JQcpnr9FeDz7UP0CyVM
M/32pv8y0ZMAiE2A+cCuczsmvi6OO98shtIoyyP8NQiRXLMCmlT9umv8GWAFadwWvE3CtkwNIAzr
/p5pt9ueGWc+9EQS1vlztRs1VI14YbKb4s5aPPpaAW6UTtgH09pryhGAwX484EAC2TQNIsw5jRbt
DHuCqWyN3PdTS59H5MB/cHVdxISImHGNRsGLhTBW7tqcZtWvKKWBg4qRdsXH5ECP269XkxQpRInu
Rvj5Pkqn9jEAm/qYF4DZ5lmrY4PYR6feWN9bcD88vkmOZxXy3ubIFF7hMaf64ecsJUVkbaRFzyXI
VNxZdv8WQ8jHGUycUhH8Xjua6LTijNEbVoAeyUJkRVi9zbpZ+Ed+bCkG1mLwJjHxUA9ZSfJhF0ej
tSl+7Fifa3G6ew34Xw60f8T9QobCNoEBZ0docKmPJdqR9YogcxSH940LVyr5/kkMOlkNRTWcW2mh
4eJU5RkB+MLwtVqw3Hr2QIIpgZxNnAsHE0a73xcXArEOPHmd0sA4EL3XNm9MzM482Q0vvnbkxGh/
D2tLmlqZ6Aha+SyDKGh+kAkjiI0xlZF5tkOtFkMUpvAO1BquMbGax9hgwjG0JTfQq0Frs+kAuKRa
gTS+fyTItFqZZa/mY7kqhDvsHHE2Rv4qFleqUVeQXzj20H2dlgApS4K2XHXrYZUN9QvblFxPNDBO
c84qhpidn6SXcu2+Cpox/7ZaxVlpJR+C+R4c6nf7Giko1UgFNZtxcsyjqPp9jD6p8xkjJZ4sRB2r
NTLpmlyXL8ni+ZorcTJ3QXjrFB1vd+inpw8CnwS2VpSsEnNZaUZpZAptoAEgHgXIyu/ELeRQdBLA
fBA3y3w5tK4wKPAzlCPrCJ222fIvZ7esmBMrnKflPtRE7Es9yM5T3ofy4R4iq+DI+B/uPxgWQXcM
Wra+Mk3P7106ApTizJdc04NwYFRR6fF0kgwsum4asCerkYwZVO2Kr36qHV8AmdorSznbHnDsjxSH
jDKzI5XEWIlZpR/vmFLU7iSAN5EDpCbk4Alfu3p+GP1F4wueYZTRdSWPYF9pexg4f/itPCvf8X/c
ZqiCbMZLw6PSZQfmnugN3LcMAOhaYt+2VWRJCWoAyiI6B219knPlla9YrvsJmtG1YfQavqWceQwj
TCe9AM2w+oK34CJPBDk4rSiqGllHhDt6/W+AmSoOZUBdpwub3rIT5fnFXbu3hfMmtgqMzPDwO3N7
WNfziZubEw2MXn3ouFZSjQm0/JIquBb63ah4xXf3m9iTkloQsCw86WUkb7WBZ+SECxTyKqyLJcmb
L+fXToAGhUYNoW3X8XnVt7E0HxJu9Lgsm2b/HrOVldC/yjSlDg9GtZ86bUD21qYzvW1rqgR+7Qs4
kKvjtDmeePDZIta0QYRpH/Ae4ppCoSrmOfQTnvdYpeNI6IzQWamsHOdQ5yCq+1xAwQqTwY2VsEzF
jyQAM4eCNDdmWdfnT7ohTp0YQHvqDC6EO4iHfFHXMhXYhgOzSmsYh1lMuBBHkWp6XKb5B5qGieXr
JhZDxQT9EKJUdyriCY4zMY+UlAsLxbkgvf+iefulfOZYQ5DN5hKi6tUEVZE4NGds6TfjYqgCkId2
Ks3XYR4D+fnpxH2jjsZ8/mO2pFtPkg4UWq1tL7v0DWOQ7SbDxFeSbj5fzeFB+5cyhcx+wJCIQ6H8
9Cg1+zxBAsRDyU7X2ZcU225eilCfVm2doy5JfklcTYJdfwYZL/wvoSs5wOiSIFWlJGog7c3g69uH
a8msruCNyvwTn9FVH8nUECG7jZiw0rW7rBCi3oq5bMUgqV4TlJUxVhQQ1RGxkzJY3ngSbddLaDUT
bhnym7TjR16OQo1H1ElDeGJvNvYrjhi2mQwb0fpUjP0CF8I59rC8u8nhhDgN6F5MoS1CxzoS3aNW
FfvuRXCQ4gdLGLQmqJSnqf38dXORlFEy1flmgvZi3bMPCm6wD6Vr4KPhQJwq0HoJ6y1u/qrVDGfi
2e9mrzf2n+Fg4ZUanpq2pRjxdYDBZP3mjliRqB7u+piYT4t/2FM+Z7s3NTmCZEoH1RsponO0uGKm
PUhqCshmxfV7UEwYtL1O+jo4TowwabRJ2JGXqYMLxMAzSb/LgvQa9nYjlCUOuFNIMZ6ZvRRvgxXC
YxuJVSdJX725v9Y1cdCjLdDPo2lKikMZzba2BN8Mj4k8miYbjcwfOCgI+yFKg5buLp7k8vcNI/mz
ZRSHEKY0pea79Eij2beJYHPH0x0JDoclCxJEIBtIn5OzvUw56KbJIASsIlETNZapYKzPHtsEsIXK
37QR8bgf19LuSB+XbAjtLBc0wasWjGDB/wNdlS54I7Tjd6ZhikIQz2N8G+ZNJs892UN1XmrXB9no
DwLH78MTDBCF6z9+/FUfFHQpJnwgWNmOW0tr0w4hgofhDgHGwJAyViEu4jaHrujeb9jUAu1Lil6m
DoOZCpDsYViiRujtIGpPaIC9ABY3MZRxbc8/L1UZkKSIyUYIefvCEbbUdm+nFWC0dcULInyin3KT
9M/Xmr4sWSgGsTLPXNJLTD6XfLUI5ydE/Fu9oiKIP42r8d8pwsGYPX7lR7Kc0+PrDo+DD6V2flIy
IUCu4sg0CJ49b4y/lm6pBQibs+DIRBwfpakkeKNB686mAwLt+pHpOjKYouzSUToP9MlKfj2j1maI
cFH5N4BHugBUZ+5R+0YvFNogXiRoRpnqLYO7kFXDgunt74eB7bEd50B0Wf3WGa5lTUm9LX2kticW
9Sx9KDVrOPgjbqs51j/35K9edh+auttJq5bT4rTUh5pM8I/s3VbgRlCHZZVfVZj+lXbL5U/u1OBz
OaIIWOCxBu/9Ph2dfimxkEXE2Y1/8mH0dwb63siA14p6DcNBSBtV3K60rKe18dzgTZ2Vhf/9QR0C
Lv8o4+NNELC+U5ehfR5JVbgSGMDb4NOApwxdL6OBAsAl9QB0XueRTx0fMQN4R9GErWadwmTFS+qe
vGCIfzeSEjj2dY0DaTPxXaZfQPIviImUEpDtjxjYEWAcI/AAKtZcHvTNWZVD9L2FW7LloeKk1CsZ
//v5izk3QaIx6NFrF3NO3hO18y47gokBAM7fqAXDh9rFd8onhkwMI/K6s/ZFsaHrNmFMXhQSots+
lwzdVK7tvpjv6xLs3+0q73yFy8zdZou2mXVHp5LuBMKReUH0U57TejItNqN0Ii/RHM2uya4tt0dw
i5Jp3PlSHAqzQ4kKbl1GLhH6u4iccQAKl6+e8VXAhImEsyPjCVm2u15rQ0PSp5YBmLZ1ddByHAHy
tk7723yZlsNW0kzQSM2KskpsnS4v8JYS+cOOMxO9HqHtnGG78Bt4mNZDy4z3+5CuRKMQ66krJ92H
sfQsMORLDJomtYr7mR+wx2eimC1iuZWx2AYwbY1z02GOcWZ6Uxog7U5+OpC73JPhCJpirIE9gqfb
7WdAeklAbHX/7l1hPQCKXCEQZXOXCUqMIv2OLSV01tFu+b58PmaMzKvlqX6M7dXUfxwvUqxLfGpL
00xU4R0okUDLYNrtYXhjtGgjrtH3bS4ckVlFco4f5zPFdZxCj6RFA+Hx9wlbwSS9J+UacghH4vgY
RlJ+F1pe0pinbzlPxkMYOaundvbusli/3l2DpPSiPwU+QwGh11CzHA+Mx0jvBgQdgd3RiczR+Dzb
fmkyNV1MvIjBNApPr8GgNJLN6CU/5XfvYosWg3VgdDod1exSlgeWqfiG90myIYJn52bNh998EBTL
O/iJH0h8Q9qr2GW+GbkeGpYj1TYH6ySPuL7Uzfd1Ij2qKavArvCAsDbO8DH753pGP+1MODbEC2/A
Zl6GRlQ4zsOqMAWfLc8gm7e+GbctUB6c/Ia4CcK5P50+MvLzISUX9kl8QKpH+Lj2s66Sx946Xzhh
UeKxSBzqv7h3YLidBcWVrNgzlIJzxcUy6VeX4J9wjzOZWiApx2Spi6uHqhj2c0pL161Qp0R3jobw
IAOVC7IABYagxG1KVXg75Bb847zGPqfoYBxU0TtEaqGsPwsJOJJBahDAMID50MsBxSC3ZcwkHGnt
3OIh8w37eCiJFXQo5JTHurJ34Xu7hquoicWbfQHpBOeaUefT2nfhvjJm0X5NMOML1PywaI3xsCvH
6v3ogf4EwhMOsTRs1lHGoWnjD5f8PQRaZd5a2pVUMy1iGOm1/fZOJhRQyZEyDbMgBuOKJAgFqoit
LkcVyvQC6dMZyVzLFo/bIPO9CgeaJnZ9tK1Lrt7h+yz285HHWB1RNQltfb0djLnArlU1PBus/FVd
ZwP9ZXNgEirXsYkNEWEL93T82RL3hLUrsAach5chGAViqAOL2Tictt5XqGuO/b6bTCi8VT3qiTKu
jjFCqBpgLKpNCIXoRAe00BN6k6NDGohvLDwNR/v5VaeuzIB5q+LehLnEgodvkaWrehzdlxzyOLkr
LUAkjAo64aBGcXx8czulPsb87++d56Xc5fSsIjuQ53A4DrXtRV2OQAumTD1kvEPZNVS8tj/eRxJH
s+tzIuuuMq+oC7bWL2l0wJqoITpPMKp7aVlipmViXwh6hWe01K84EoX/pMqbRAJPhWj+PLaOPXMP
sKGmU3OYiMdDJwB5/mOIfnpwRwWWst3N4NJJwwDX2ra5E+Gd5njHg878e5hbI04mYrpLOW9XXoyJ
apLtsknE1oU++Ut3mNstyhSfGpQac1Kov9+cnPZ9KHtJclXQlpwP0HDNoy/TGYSIZxvj0ukjazxc
lCHCqO8w/IbLZ7UlWlgH1LfDquH/1/lq0gR1XcOOSxPnRjfZ9P4Gat8/ugPF+/svJFnoPt5qoJQL
ah9SOBPECRGe6Olz6RROHt9yVlU+LM1H5aQYUG4uQ3BQyw50d3J0DcO2HYXCkkmsiolU8uBu61Nt
ixTI7rKT2ytDkPnvT8TZEGp3JAwsSiNmLLiBcsY4wUg55rBZzqa+yj9WrVoQTz4Kp1fic3KqcPrE
L9qwdkI2ndUp3fyG6LCfYl6p01Ru5pngpB3/a0v/6pipccdRbWVQW6dMRGCFmoMTpW/UZMDcwGRA
2jr3Sq8UaafF+F56Yo+zFQqAkbQE0xQD1hKz0A3Cml+kXmr0AyjX8g6YpM+1waH1Dtv5kNGSCEHt
V8qbmqSnQCfgoCbcqWpGapOXzfrymJ65sY4/uaGG8XXTDztI1n3SZ3ksJ6/GbWOvOklaBA9quQr5
+wW1Xb9qks0FJMLKZF4U3U9TUsMV/Vt0ut9HcLe6SSOWTCjlJ8uvfYuMdzrQjetzJ67wiBxDp9FB
MjomYoUU22hunTyhjYB5+sXXchuBSMl1ZwjFlD8wJexQjpdnhxx63de8WR5jlbF1j42EHvkq3oyc
dcVWcSm5pEYmh6UmW3QGIdVHjQIiTlXPf0/Iu7sV7aIqaHnlvdJAfGx5e9xJ+zgdcAdmlchWj9Jk
+Dz6fGv42B7iwv/2eGvPx7M9D9wY5aECaH7CmSv5J9ViHH3eEfcgTePSok5LxBZIIpnNpfKa+nrv
o+ACeaUb+j8C05AZ3jhg+vn+By9aMvsvHbyzDBQv+vImqnHiZfoYTNBUcV7h89wjrly6RAnBhjsr
b946JeGPM7I03FSMQgnOWkXJJkBinMfjj3H5O2t4/Yq3NVeXKLQfQOYr4CpM+Y0qsW3SEecqKSn4
+24FV8QI/qJqvA/co8P45ZB6WaxufHpGTVCzpCW2YCUvquZ/QKnkgIEcnQB0CTyVIUmuW8W261Gn
l+5INkfW3CaGOj5e0C7/7PI+JlFHI7DKrMCNoySxQl5Jp2Fe5YCxmryNYHJVyxOpk2dy9ozb32Cy
w4T9EG+pnfzSTmDGvVH6l+xJHDtPG8KN56trclCpApT3elCJejdgd+xHf3VmyULuA6Qle7LUWPjW
oMxPBaAv5XMh3uykL7xG3shf0TKlmbme0lf5QKXd8aG1wm3anDX/gR5gvLPe7IncbN7EB5nfqtcl
L+faI0jvxDqjnNALUCPrT+HcqvQBGXU59tqsOOL9FuC8/JgFMSQJR3ntS7//Uhaos1D7sOYe3kG9
OPKd8RNZ7H+lVaSJerGuXxckVUfLbOF6wRMIV+NixW2jTC8FSXjv8BdEbJ699ZNxwEgBMsLVfLeO
6n18JQeDAyiLC79C5wS0S055P5OUQ5VQWZ7gG3FmmW4V7mgMX1muK4n9yL8nITnU1RA5mp/6hlV3
Ngd+HVEMKtxlHQldXkmQRZzaUOfHNx3/XuBvY/LKMWxu038VxatxOKbiUhzgnciIbdbgoR2coZTP
7DO7G0QTZRBfoNK1l/56KkVNmiIgCBnZKsGrAlDEzS+6dVyCjWsy3w9sPqpdEprYXj1zo7RCk/m5
F5GaGw5tFtVVFqrkCSbrLi6jbjQ5AClZocmkYYjo5Xrcxu1m7hrXfDq4UyIMQDhM6HTTUw0OSQJv
E2j0eaq1DmMvwo/b2oh4CRNuHtMr9JDD7RH/LMycnDotVJx+rH+RyseUqJ0bDpi+6CnP4IpE4+ij
oY2cGu3kHPPlyx2HiImd5uHz37h9H6O2QwSNhNf8dqJfpYfYdqZa322xSScVY0IDw4/2CS/Pk55o
EUM5HLDLkmWkmAC0nTk9KCCEcjOnjZqRhp4C9MFjKUULC4bCHTmCD0UKD9QnE9ta7WW0QagFgJds
esNAmyehEn45deSZNzzp38IfHsByI5bqQxrT4KQRr8LKRoDe/FzgkaJuKx27QNpMITwHQ8D0i6X5
aS9zy9ZOpONgYmK2YLuuMgmdmLUnPqZmCpVAtZcPE/FAw5ADdNOdBgg8nDbdMR6aak2JifliEcts
Ce9ebq9ZO3SM3oWNnwB8e4gEXyBUcNc2MtCosH8qkc18vtFvLq6ogDUtiTYmxCK/9TLpmwpKhlsN
1GggDUX5aFBrRtuvYYtnSyfS9pZJ18qxiw2JwT3dF2/Tjt48TGEcBVHI2mHqtQPxoDeQYC2augr/
ySHQHcTVaY9VpnkAE8TDwz/+zh/HeL7W/87kb5p7kvtar17G9gz5pUVWkTIbrBlQS68lCXgh/gVe
woUPiis/DGlvoeFm1Lfy16rD+Yuhs73uWBBnMk750rDyjgx9p3sg0Du0x0k7cT8PAQ6YAf3yIukq
sfM9oSeNQ3jijZzfhzueSRGb6AvcwqTU0yScgOIGccAT83dpTiB6WkNR0u8k+MxJOKSdhTH3cBmG
H7v1XnzlpnayMmjfoGEpsAbpI5t8YpujzUQApQ68B11XlvDL7kIlcwe1XMERlPhhe6LL/WhLP2b7
q0r0k9jNI9oWmsbHN28r2ZSzVhfcTlOwIXgCeaQdVy5J+HwJABzN3nNrPsq9n3p1zEnep29/a8Zj
gfak9rQ5PibrUZwSycCWw3dCJTYr2QF88Qg70sVPCd0j4JlCjouLEMpUYbSAjRuY7BTpuFi9qB5p
AnAMwDrgPDF8gfbBMgwVrEStdfiuhmGniFlr5onbgSNCQDfoI6cK0odW6Zq4nxAZepu+H8pB8Mm4
iNwKUphrKqDwwRkhLXy++p9m5xpG0CbxX2EvIY2mUfBr4bqCfdZK74qq/yXQzF7tYBUZAQm71oJw
iTDsIizyHZMou9x8Ib6EBwSRPU16/5sw5FQ+u3oBOHGwEy63ZWIm/+aYUnvJcD3Ki9S1XEj7LLfa
a1aBoEaIcpCOnxPvzaJJV7OMAEcL1w09C/l3rmBlXw6l5BmigwoNrRxn72WL/TDtu7aq/5/usXpE
+sOjYfkI3bDZNQgPSRrbkhwU7zNfL8gIdoMrEG2keqzuwXDp4V4W2vHt6bb77DGeocDM+rPF3BFG
pj3l0iy6TckkMurmuHaL0g+3PjvInV+4K0ErVnjl2JD4AKS75bEa3UmWKEEmi+6Nuie6fDIeuv8r
sijuZZf1aIr5Wy725dUhdMBANmQVPt+O/e23yKJCgAsYPGslBYH8ATajT1vzm0yYAbKbwLq6CiYv
/PZg7xuxUn1uuPgGw2uLpKedxtdBkdsAwA0YHC61FiiQjDZJUxqC4hqyQl4MJb4kp6O5T9/Gz70e
wfa/wURmaDf0K7Pm47eLQaQdooM0ygSU5VJps/MstXN3LKMAcEqev8EDUJa4YL1MPzV3/WbtAHlx
05BvnjGYjeJv2cwgj56SZ8nggw8EUSaygf0ZOw1bZwEwpyUCDhS3FCKtL646/2boNzevupVSlKKT
EnFic1mzqaGq871/khn9e+/8yBqzl4gY2cVTacvbwzR8E2ln/TBNrCEnvEoSl2hMZCqpdBbPafjX
F5pTdj3HgiXrAEctSWcJJ85cKQd9/CD0YnJpYdcH+r2Nc0CEQ0PakCKBxXbcktwtWKO5EjW44CW7
+P+3Z+rmEUVHmhzHObomESR/7ywfXiDuKZAc34b6Zm8FVVt5uh5RTKDhy8kUQFYdu3iqkw7vSn9P
HSFMgUCh/l9iJlqJnK5SByv3ERcio4JniNYpjZg6WjHuVIdeVf7UH8u7ViF7KIyvt2OpB9b8Eif/
SsCCUSM873IkcRlGnRibq37wjm7NBsyXG+u/qag62NQU54qyChEIe36XCBWBhYEalmXZO8fDspxs
8suqTxZSieRKilWskSlTeUvYxtyJaxzwUzjvJV9TzLw+ac5o2TbHPFOeQquxU39lyfIMGSVsil8E
hB1GjfEIVU8M6jEO/xrE8RZdnG4yH3fhSQq/URVRlsvwH91swaAQxUgF/LsROfi6Eo0Xq0+Nnhbk
i0jogvbCbW3W4OXvpMEhztLBiUb2d3mCEiTMI4Ip/A/o2xnnInjAcuthUg0bl2/DGyxmrBuacO9f
GvTRmBxl522bZ8eW4tCtDGT2//AAKd3MznqOu78puqPZeuCe5yl5ANoynU2mTqcGYP+5OXe4KH/U
wQ5gqGf1TkoQ/ZHcBcaSrH8VT4avNw+qGVhBXC0wVtH22ZwjnFQO79s1ueJ3IQ4nPMvyQ6nu1Vey
aI/zmPOjwILUF1B8AXsqsM9Bh8Ik0ACZSI5gL7X0Fq83szmGEMiMy7yRh4FDyQxKlCPV82gXTR14
W81ebhBT1AqPxIb20MBA2WObUIi3xzTuAMkdx1UEgnmTl88QQ0mk+2w+gdpHGNLJibl2v4zves/i
ahXSro+DWxo5VHRUnaAOIulpqGj6EdeOdl+PhiJp6m3DhU+AUSuADgI+kB0qHF5y049Rbh0wfI+o
bzdpU7mmIPxIFRTLOl6uZBWZrLTlKfm+pPT0UmVPV9vwYwQP1yOadm6uDyT18EqKdTtJmzIuoozH
8VX6jzVSl2RIU5VhkV8CRCz1lT4c2wNNKF+nB/Lg3a6oVxaJcyxEYSrIcJfCmx87YpZPksTTYhD3
z5MTHIhR8DBWbCw/7UOBWaL2Aj7ADHI2rIAq/IiFpFbIu20Lw1DSvDdK7ij3dSVgDXAWhn7GGWg+
Rj70hfgBQT+KmF5N2Z0O7dJDLOePoH9fGGZvyL3do6qhmkqC8j5uhSmI0bFjQIhCFdEzbpe5nnfI
3ZAxngLFHOSZbg8yZMlxb9ERFrikmvSbflrTaqsDOmGkrbFt4ninEfBsyNa6KzAUeVyT3a8hDaQj
9TvLoPUX989mDxpC3XT2EbnXATpEqGQ812uYIjrBde1zWJRUoyXNk37jJsvfKD9L9+lGuXTHics4
DbCnVIoSJ5y0DcL5wd8u8zwWc80YQXuNiFZoubpsA+ztJJHSDljsRjCiy6F/WnHrKV0v+N2B4Kja
KQ7grMAv2fIn/5Cxfl2NNTeUa55vgJjNOJjaA3GcEywAHb5C3p1QypoPbwu1XTvooSifnDmuVMfe
ExOhyprh1hsRiGynXcpN/PdJd/LzSkeRVSiTSmrPg/VUdQQjex7LL8RycM9ouMhhoqbw/gcdRnRG
IONkEVU/AeYw767mgMQ6YFMAu+kdqU7BW8admZ0nndAfyFAUmqay/IN5hER4oLfKYGtfPVDvus0t
M5eRmKveddO4rPrjViKEQDPi9v+E/29ALeXq0+Cygvr27KSF35FX7WTixJ8Sxu5bdXmiSkoaSO/Y
Jsi4w/jiAbeqWWPVxPpVi7TmcmvdJ7U/pxZVDtG0SyJe6cdVPR5EE1pNShz7vW6kv5v9uJubXQyV
vlicvy3WypkTJM0iNBTtyo3WeNkjM9rzqE/Y7PqbxChO0NAXx2o4Y7dlETEax0++y0b/y0AlA1mJ
xZ+S3wUdIlyTvLKKB7RTGXIX06Y2ZDd3GHGOF99ZGJlxHrXHXMrFEtCuhR96lHriWAYaRSJn3/KL
jnOswvtQr4lHdIgRoK9h8Fmk12Ux8s9g253SHgMSOVtKZflUP6S5G4mhjduL30r7nUT1zU89n8cv
5SDfCjAqcENy+nfoQ71kjjY2KuYGdHA2CqlxH2DM+c3+jdtVKDpWYCpFFEpWJaXln89VXgKphEYK
q5N+94Yh13+v72tvjNsNfsjkerhkjgjwULuPwbhVFA2hasxgqB/9iYwUllF+TFsSrzgRgZYlHEhd
80sKtFMMV6ZNENRy2+puvQ/vRIbbi8883xneOf4kyYARUcrvnOBmlAOg/F1aMAV19ylbnjvDC/7i
YgPup7CdmUz5+KoDb/13RzTuSwnHFWVK57FR6V1J4LvLkuiZSXtJ19rDKVo45E4N9VO15rnqjT0B
dpgBxfciMi5BibEQobkhMwp37VxuTM+Z+uhPn/v8kH65X1tUecgUIY73ILtjMVceWT1HnYXNBybA
DqQ1eLSByMHTxWHcyeUce/a0PJi0QnoFFocTjhrncxkAb6V72Hrk8dGoCN4ReKOLj8l2sBNxl73v
6jFQbbUrATKK+P1GLQpLBbUM6b8H136OCwcDwsP+IV7Rj1F+KAE8P5JGTtbuLerGEZ8T/2Y9EA5s
xyoHzzbnyTzdgKHde6ewMU0XkzDmL8R5A5KHBUOAIpSnQQ5ZXP4lKCCkVLsHp6dJbF/e74T8ZDL+
Ju0hKwJWxfG4GQpzvOqg2wNh9R5MpYISCoXSoGzDTWRUfUmSz72dGQlt3kjDSZhnf1P7hIrsBxIx
L31hgZgthaapRmUYbXo5Jmo61MZVY5Y3saAt6xxoE0YQdQds7hBheVDDFJhujrq1Ngfa+Pocs7Vn
vzTPYR4d3cAW/9QiJhJ2PvzJBEWsQFed1HKhN+R5A85eJYGyqJUt5F5FLWwu9V3bkjlQr5T8WVos
/5hfuC5GhHbjpeyrKJDKyrIOpyEyy8tfGhRZWZKNPs0J4Fsme6NRqenvabGiu647JCwYe5g2Gfm0
di6vfPKTku6kZCf6VU0RxAsUrryq+XFK4XPrUXu0AA/Vii7AeKr4kkDAv4MiNzLYKfH+4lIw3q3E
YCC/bgPuJwZYUCujLoWsbNQ5AfjivR9jr+O5/iUCFjiy71CSIqUeAcSTC3N4HsVCkKEf3OynEziQ
4VFXb2xsZUqrOmIPn5Hxa+CXWAJidhVoBWyAD7D9SonZOesX3xLeGFQ6FGQGILFmbrkt6zmeeDba
K4eftK3QCW/rnpHnllnhfGgpNTR/ghCBfaZeHb1d/Gyn8NuLq9mIOJ73BWCbJlKiV8YsRT4aOn+M
G31KexsKPO+rmd28xWsIZOw2OGkcjlYOVQewygt+QhrqvePSD/PYlEGMKnRQufiG3AIr9nGP335E
CDez9Pu3nRYc87T/ACv8A0cjxEKA66RT4TTN1Qsy9gh0YNIdC/qIvxGNu9nwYvWWQdbc0ht16Coy
d3XZX2aQAHRBD4bNbb/uPaexfH/sYNGa0Bb+qS9CnjMPFixIVM3YxWHm3ga+HeqyvXXbmA0P/cmn
1vfVyllB7QGZue8UIISa+Yt1Ac0fA7l/1lOk+bx4e3CuSmIxtuYTyAt7+la7PN9O55Czxx90BKSe
gTO16osCmlw1fNnWMcTeNelthvx69mPQtdCl2Zm6yfZXFI29ZMp5IHBxebSx023uYbNmx9iMXP+L
wbTcENM3y+ff3EwVHgp03ae4EiKBySqysil2W8RhPsT2/iAjWMPHuhrU7k1yx6esQIJnsGOgMyYY
ZjLtBMEfZQz2nZWVeSbYZLYCHI4K4iW3qJ3729WSLehdjMvs5tz3tihAJYPCI3xE2ME1cDgBED6L
lATJcSX40Wu/uhNpvIfYeYu8aIN+wGxzhfXtD9KWW/R8lGJQ4DxX0cudsSBZBg99qslc3Fr/TPdl
otnEs8UfLj291oClT/7zwHP6Tda9ONUIr0Uo0PLj/NtoKtfw1EFocxWoFnISwXSDxlrDsnEAmtfo
5WA8FLQed5YpkvsqyO4pqa1oEr0qR6aPIfhA3VY7LyO37q25d0QAFfJ03iav8tRUHaGNRYRtzg1y
E2ERzg68hue3rDIVKNOUuFK1RqiooaspacJXvdVTyh/xkU0QG4cDZUMDBAtHwELx83NIvlax5tjj
MDxrEpL3YbojRLA9eNeqfMNGYSMzFY/K5XB5H+3q1K4UQYVwuAOnnxZ9Y1amOR6Pp4XiRIOpkS2G
zFiyxRzOak0nZnwVH9fbYsjIXI+DLhDxwl4niXPnzdszHZkXHb8ylwfrHsaVrjr6lIWASKOidrGL
1zCJF2uWkdHeH0IGZSjEn5li06bIRBUR1YHOXLctb2TEJfqlJrssaaLVbdhHjOTfWBAdk4OqV4D6
6DqyDI0qGbSgNEpej5nBb+Xc06N7gpL1FPsjXcQ6b5iukvzunwsjjh3hOqh3VdKSnKRa0sPig2SP
l6dSPhK7HGAFKqLZZvTzEywexglVyZ30I3YmYViZbC3JFO37fmhzdDpWPaEDTzGcmfMuwZn6n9ii
f+/gTmtCw3yRQpLLoLsSdij4eluIpBsU74BQYkDyz+dxWmHlGcu3uVpXGMZS0pNG18jz47JdUkzz
jlsy4/xNc6gfbFsuoquDDAUJWZ9CnAXeC1053mQi8UWzi8D6qh66+yCAaniILGeg1SAVmQp3wH3X
WKcxYPC3i4kp8DIkHnk1PNfyH2c9skAv65Siqpi3OstPFzxnwgB4eFao8pJ+POpN5y1L8WY5NtDZ
69nkptGoVTeApnGFns3o9zP4gadXMVIBfiBjwWkW0TqQZS2dGeIrjRSuzurs3ePkWKwmX6/4LioX
MMfGNBjUz02ja/ETKEFYjTe1/8lLLXPF7pWS7x7t416HwbN10Q0BB9c9InX9NyGiwAMI35YQW7/J
tKMZE9Cfh8hLV3f+4/+mmP/iROgo2qq3TIw08zYsYr28pU0G6sQIu3ejUGyGgbe7zt/yqPO9RrKv
ZvojoF6E4FWXB75VSgMYq8e1V85DsU7w5+8djLk1ftqNdRlVHLhVwSxxbkXDbY4qoeXNcpdKN/Pc
4d/0If13fDNs+hXkocD5bEjP+PibAxPVdbxnAJbWHmI+RM/avpkvswPq4yHg4gEclAyq6OTjEq+E
1tt84b78HKnE7Dg3EoBQy8jatdGkEXFlYZ7kCvUvH8gE7h6SHmrxvGq/quuANfqi8mYbkea889d0
Bo7UJwIGLnAC/rpoesPgJOM+JfCx6dovT8OtXf7A/ef5Uqul0lO+G9Y7AGIuLzZ7hoXXkXzyRt8p
AkO/Iw4rLPlC2ltia69D+6BzuKf9ulHqyA+HpxlkdVWTN5WOdaf2dKqP4POz8d1vdjeAaY7hXnmg
F62ZLubvdVsodbkxQm/frhzdzfA2/YIaDjdz5k/VNu1uKI+6o2QHqmHKt3EEBr7mCc+hzAd6uYpt
iBv9nRfxxZtMnBJqCVL0LSYE9HUnHtPROyEvynkl/9UAcRsm68PneKiTrLIS4FM3PxMxJ5VJhrZr
MlemkwanrD4jikQrdKx8ftRWaQ0Bc2Q6bHccmutKwmO11Oxgh06o45o+C7twpN9lG99FhKW4vgb/
7Sb2JWj+btWXNyDhR3GzfLBkdO1ns05QerXuqshc7DBkeJt7J2MEEzZ5d/HIgXVYyL9+i1nYBC1U
VuFL5xtKIrEKrLyM5PWWqLS9Sa14gVSk4Cdd2NPE0jy76V/CgNPQqQU5yEPLkJP8Rbn0B3yJ6eS6
7xJyrB7xrmwZGAN11Y/jemVFvTz3Qrct+Jj/rZe5vgxqN1Chzr5t40j0c0WnWQLIz0t82P63nbmF
YJmzClzZ1G1YmVsssFpiOnvA54XVAkWP2SmcaLbNKwR/JpGIll4GxHU/w0Ui1AMhi/LEZEh7Py/l
8zMZvSJUZJRTNh52H+x9LFtmcxJlByswrNkV8oSZSDWq7i6MdAdCS5lAFBrlwRKa1dE9WtG8uPDf
soaaqQap1mVrMzwIAuw31rrYhOS0MtVDW/cFe+VOtX8ZuLa9PGrPxIqRwxjOL5plaLnZBvXwi84f
wIoD4espmI6KOYvkkd6Gq3b5/tPHqFY6JTTWjNZrLxaTqAOJAKW1n99WBRnXraucee2QQRXuphqu
rSvFkFp0T+OTgGLETqqXXBpmzxHk5s2cDkgtI4XhAyLZfYCNJ+cg0jekOc3JPE+hsNluHBMKfkAr
UO85hmuhFC6XuV54W1fHSDJBnpuB+tiNcjZsfoTnERvdRs8qbJWEhCpO9X8rB7yKxo4Ut0f/VF23
EraTNPs5qR9tUmxWHwHw1CRvqL2TeGGDByvcIXd32DCvL+yJjGKrf2N18af7ZfGxZeYmVD6+Obyq
5QdNrHw31pd5fjtUIVmxjrMZgER4qU0eiqpVE8Vs0M6LuZAkj2/VXCz3jsfkM+L3pgP1Zkl9jHuq
81qOu7ewrlh137aS+soFBCkin6Avomb49ttfFylbXCyR+xZ9ID38BWPXdXQSioFlxQKAPP9GIrDu
NgniDVCanOFwLdeUK40SdzBKqrqgSEZi8cIJOWV60zw4Kv0Fse9nTH+bpesBncR5ID4fC1RRlYHq
5ejpCZbbq8fsm76uXSLHuccHRrDtiXfcDAs89P28+k6EU73Rq2d6J66FeRHyXTwtGVL/bGE5C/tO
mcwZFHf1W26vwya67WvTh07HdKI6THN9PSyRhLtnB144OGvuvWlCPeLQ7w6M0pL8lw8UrTUnp41J
S1L3uP8egbavh2rXgrVuyiTJEDmm42qz0Fwsld51pZNhDxNVmkavNTexDOZbMC5KcfdxBxCR5RSu
asF3zo/v5DfI02Ndm8egcGZSIcyqaY8GmUs2ki5/j6JSes5OabEfPE9CACPg/vzdnSnEfn8g
`protect end_protected

