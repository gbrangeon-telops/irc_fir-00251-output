

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PpoeUczC12+YQ6zcBW/hk7KVg+x7UTioMUTG7QSkaE8DKLm5OzMFnRnSP2RdM8C+WL55mLvLDYfA
5lOC4Ruqpw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K3yZ7/h8XZC4VnxKqSX+X1dWQEKELq4EziAIjvSKKzex+MM5ch0NyAGabLWybM0VZcnyA2IuBQRw
LXtEZmU52Vw900CqGAC8j1ob1JJokunlfDgROKOp9VekmhrNu0zlywHl+eh6CQ/t5W76EWfCnLXS
TKcvUxKzMPqBkiVg3Y8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NSAGB2MTAPfuv2AfQtQrWIP89UNTneL4Bk6/B2TdOO+6mmG5j3iveazvIvg7qIHwAqHfCGACbbAp
fGS79Be+x6ilLMPgwgbPlwYl5oARsjb29GILZJJbq65kaBdWWJCFrRmIDIFHXq65c5qChGV/7EF5
BRY2p2sjUe67cd7MFOLVO0mKHurU5wiieT+wdpbGs9uEgt/pGFeQKlj4ch2XzN03R8Lg3KmqOC6w
j6pa6lYe8j+sQMdh+WMN3EmYurAN2aA01NOtdnD7EoaLrP3ByXrwCKFB06hQfAMKudCun+42nXbW
17uiY727vjm9PIB2xOmQazUdPEZbwz2Eeua7KQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NPiHNhu2YI6wz7attBCDx15tEqFL81ie9/7cRUJzlr+aO842fU7+GGF/JOlqWsuQg2RB92onmIR9
gKmj6xIVPN77wRnezyej9aQsYy3bBfOSvbf7a7d2lZQT1pTZcYMfp3xveVQ5gTGk/1BN6rnnT8J4
QRALHC2oqPHhQZ427wg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aHttOHUQP+m+tZmSEhqIMk3Jbc86fWQ1/2LKPbbHBoOHb+XyETCjDqnDo9IWfpo+m+LC80obW4Zd
cXgM5NoQ9F1AYdG2ggcdGNXeaparpheOz+XWEe8nirOAN+Ks5VYo+yRWYwO3R0Y+0V6Yw8r7cd48
CXttfKVhu2QOlKTiKegYDKMRGhVyrdNkx/KDldRFk70rkBceBbiSjdBniOrozyhG2imBoMkKkCmI
8TwlLhPf5Ra+r8wceN6j4BjOnyQ3EtzJgw91ujnHo20MZFiaPiqLQIavDgBT1y7leXT7TIK9Z2uu
L3Oj5XHzPc1v3FMsMkjnu8xWqC9pP05Ha8xR1w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26736)
`protect data_block
4nct62pOgmTVzWSAG8z7FnHJ7VpnqDI77E2wZ6v0xyJ20jIgNxYJWXiVQLdTAzgO/oBGfZVJj3ji
gv0XsXn0jX6a0lPdmyEA85HybC7b0TC5tF/msrc4XENY6Aupm6dcgIlsR9DynfSH7A+BQMslTT4A
8sWG1flyiGbBQ3LDhwKTg6n1MfUxW/WX9x7iY4cqc4Xmfs7kfc4C/YIli7oCSep2K3kH91ZQtkz+
Zxqs+1HKrbQuzTcyShuXX2QpNdNixDp4jTBdege2M9XVFXbOS2YqfQSG+s6tYh1IM/0h7gbGcfNs
G8WfeT1WOPSbs5ecZSjiRwJOigPk2fqm5nrYES0uOLrezRqMcE1Bx3ocZ+okP0tI3+5HgowgbLoh
q7dkT4crhpfUWfUg6KGAeIQCxgYCMVD3EEB1j5NlWYeRXJuc8cmgvYJetfCz4pq6zFmoEFitFYAL
vG4nqjthhHJAjc48nZHgssAJXUc80+rYn6R31a4Hw6hRY9wbynZMpv63VeEC+YXNVVEaejjel5vs
Im+kymB9J39t0vKUTFNqCM5+TJxZCwNKN1HbrnO042YGY6ixwklXp4rlbLshU2mTzGuGjvCTtWCn
amIFgublUnElGjzVewyW7dSLMaxJURMt2nZocC30D5BTkEQlbAG9DzvhhrmnPyor0cPFYH6dO2SC
y8ijeBDLpC/C0nvxpaPsJlRykzD4OdwiFP9/sAg1dIcAR5Hi4B6T6giCUPYs2So9a32IDv/88kXL
vmFfn/rjmoRHbIA6olVmDkVbFF3EfUNF7wIpf0Vtg2RqaQOA/z2om6kVhOJu6aJmDQ13WndfkTZd
fHVTqLH024NB3oHaOu83yLfTfJlQy4rGrT6eAbnJAS1QReJ8QegoVEwYUExb2v3jJiQmfQeffRdr
YU5poZquLMpLOHLVI77C3lMX1FB+WTi1649Ad9FDu65a1I2p2uXfkWGHcOvnvnmNCKMSWe/yP86L
Go9QcnOW6KKQE/CTX2ODGCCDzsVgepOtvbunTf81vx0SVmwp8uXWsQBx7jRbDGHmzfMRZpzFIv6O
dg0GuDwTAKEKvr1Wz4ecsVCTTxaHRF7q/XA3BGO1fbOW64SsFYe+uB+n99p4jkc4x3wvM3Ew3I9H
qJ0IrDC2To4vplpe9ykPnoRcsEX/sUuQ06YWjVRRRWpacROH2S2TfgzNQ2qi8tlOTga8ZGBfxsow
svuB28wE60Ab3PJTqNw6C+FHGul+JSK8pBtpe7X00eKJ6gd20SX/Q3S2Mi8n+TrRO7IG0G3umQcv
fTLtosqmxlMoaQx+foe2rSeTMSEUbnYHJloW9PpAHUafZYfrrXnNUZIrgXA84TMVw5YVnomlmIXa
exVZR/YnfKHRcD6YI9YhEVfYqS/gjXIttCMZhztlFDgJT5RqY9ZoIZwRnmtTu68hnhEIuZ+cEXd7
rv40lCknX6eI3I7WyxT/UNnbzlTyzOEm2knaEzekL0RUFhUUfGRjjny+9u4YEasS0JMiAMifCLeL
HvkcgqpgO6OWX/7tGQW1GefbvASRuvQO4BNgfwz5Yrd0UfgWSfvA1fxj6rzvavmwzGZmy6oGdvFw
3jIkYkkL9/pUWa3J/W7S6MIfQpu/WdBbgrU5XX5hPKGG2Ceo3n9JSa+wC0/c8yHGJBx+GfA6KaXw
099nLyUDKmw74/q/TetKAVjXRfR66aNghQza4U5xiICn3Rp5UEEC/nBhnr+R8rA/ak3XI6KDn1dM
HGelCEkC9xH3OqBCiRR9vQL9W47S6YyeZBWVpKgTjRKO/IbyOYfPKYaS8/zuLTs9FJ7IcX3S6CZV
oPMbUsCyGGkh2XlnYTvtWIf3UqB1txZmStMc59P4jORI8ZejVzaC5fmrpZ5QXnONv/pwvo0zENpt
JYBu3bt8pUx3RNZMxoQS7Gt0YbabyTwgNRIxjoVdXF77ZD/kdkVLy91c1+yuwAfz5himI+hkED4J
VyWsCxJQOLWJ90THxHdtpu+dCrgJZAZLRYyJ5svNE2CTzDsOlvUfBxfCVj22xWQaDjELD5mQqCar
p/CHwoXM7HZ8b02uI9CO/e2y7jlUEPMjINGiDk/UK1fp71H6ioxlKXvugi54UPqQyydbqSHOnBl7
3Dqs/ghei0GkBntC7wOWCwjHXbytzpNiJ5jvztYiqsPkFa5Lp4pdu9EbctWiRt55Lbo3K8Hdu7mu
SRf/2ti7mETErIv+6ywVYbPyJuotWxZZLkG1x9VZv81eyNN93J+71K6fbyQ//Kca0TIAU8LsHxac
/QtYoKKJviu7HeletzX+9CpmXlMUcar+UtwsMrQBujR/Om/5yHwysZr+RITocKCYjEgxwkBhJF7B
eBsSfSuxOgfq21oXECTRcs2lVp6tY7SRgL4757nR9J8iGwzVcguvcbRaqx1As5SioZRtcLdDB1mX
VmDycNqLkXNS3c6aYc6lF1sNNDfG4HfYNif/J81+NGkp6aro4MHSzxvC5JBXi2dEdXdJlEEybP/5
DtaWXtes00sLYi3HeXN+AZxg+o5VJGZMRVOZKfM076JoeB3NNopFGbDM7kTnWPozyKO3YK4MPgeK
+pUDiiazbE3w15UKiZCvBENwYnY2Gi8Bwz0uLKAE+G+Q59vi/EDtrZ08nDXu5eF16OfcsJZ6+LmO
NKXNWYyfur49j3rvKAqVV1snaxdtBcD5DDalW1Sj6BNsQBj0XAQnQHvSRInbXE742yzmr/KNzd2T
Cxd+duzqqfDlE7NaGsa9cbFbOd0A1H+fXqSCcmrMNKF3D9lWBeS3f4d9UmnJQOsP93WL+GASm0J8
uOWb9XrUyREE7bYomBhKRwACi7J8fnRBgsHV/PT9aTEirlbn5ki4n10mBnMft7qMGuU7yaf6j5n5
cnXaJaflA998S1vxyALCd/2e1as42lFScAUPNlEenRmOaePwJz+2q+V6PDEhffjS59oht/b8QUSu
wBWpAsUZ0gyi9I0AT6vsqFnn6ycLIDO76ln+WML9T0TyFOTGQ9QhrH58I1AhEq3QtT59rYR3vLWK
JLH3irfRpgKhM/aPcH/FUHXxjuIdUkoiOeboDBI8xDaiL9v2qnP9glGpMvsfEzSkXlmCZZOXLDbs
XK5pPphfJTCx6PDtER0yESaX1HFuPATp20KFV0MiCh0TlJsvhOXMlqe7N2tJY7elYDfYOx4F+NMn
T9zdI34rMc6CpjM26qWFyaTaSeIAas271VGjYdiU6za7UR4IG33E6Ybs1hW3EeMSXgGv91lsp1VI
Be7w863Itjczi5NUJJN4AjNmTI/6ivtL8273cBuzxy3ZTe2vhMc7srbFnpaT1wx0MAJ0MBW5q/L+
HXDeqpi9XWAA8jYOC0DbSHgU+NRYOYRDl9J+w8U981es9Bpi1fOLmAgXhUYOzSnrXOFYcGmUCjFg
jfdd29C/RgeITys2XEhcrZZCcSj5Dlw2hxRNfF034lZeb39KmB8t/s0YasnVFn6KgLk1P+UInaVu
06wFxyWzUEpGMJliuuyxZ+e2hChtLx7K2TNH5n9rlfGVAVRc8BuHIvIsh3mGps1mT0Obf9mbesv9
OuYU8KVuVS22ewsY1DhCDJdfSaMBwDQX9XMAYpfYmYe1dHIjt0972UfHjqoA4XvPd2i2itbBdWkV
Z9jxkAJ3e/xKI/YCyOvXA0iqZ4LUnDqw6JOcZADmlfsD4IQxOoDLVghKuZstWyeiY843OWffSRy/
P5Q6VJ+FAeYa92CUdKi8McUsWW55tb/I+2gPMXVQ95QZVjOcpAlK2it/Lqb4m21TTXwDhSkG25bd
t2ifXtXbbMcz2HgCZRViVRfis6fo05pwLDpx2f/Ymp9y7d8IJ3+qld+dHj7hOUvSAPoedemokCCO
5YieWm4+yi0rl4BcIgbZCdrfUFq5cYGWTIJaxOfl95D9otJ128stlVoUmB7tMwSrKiYtxqEvdQp4
5rvqz53k57y78ZVE/rnqaucLZ5GQsUXkXxqbdh58B0sk9nH+jU57WjGk1rTkc2ltZjA35H7nBX5h
dA0OV3oAsXYXH8WJn8Azgc89NedmDl4+YWCqSJiE+dEt03ZbaeEVegd78vcdnptWWWXEQnZZL9km
WDaKfnmA9nSFGM8JtXiYRl09qPBoNJawAR2K/8Z/5HbWC/gYoHQDMW5cEAlTLgbFIjqGYqTzs/l4
8uEZ9au0qVWLPTDyZZg6ivj8BNdlBi5Zxm1GWZCWBjzFeq15/jUIBM40VJ91uBW8pHKigij1LR4c
jDAkKTPwfd4KNK3XxVbUb21pcHlUQGl/o9lh75eR3pXMjWtaCh2vi1b4p6vJ5ZvbkmvE0bYQqThs
eORKZQYrrlRkOlsnVHr/YFP0aS4rG25XziFKfHD8wW/4lW6WJIMy4FkEbfWTY1kWdZsgL3VP3iwd
icblYs0freKJor+U5dwej0xM/nHdWruOHwpFrxi1EUQZ3oWXn0gSytXqP/CEsRUsasXev4KgJr2l
yi91oPX/CxvfFn+3gG9cf8WJQAxSgd5/19gfk/kOZet59zWHozZeKe4q5o4krW4H1/LJK3g0hpyi
rmX0QzKPlEdsY/FheJBkOrcSnSAb/CxLi2d5SpYX3UQLZDS8XhanGbU4HhAGMa7YUK74N6/2EGnf
del/fpcff0EBE0XNg98hOL+xN3YAg01FQZ13xg636XYZpVDRta9MHVO05nOzuvNGl5Gro+9FSXmP
6c0bhiQVg70mOalSPAEFdnU/RA+2qAed1ZRiAv4tgW++/znNJ1cL0J789qrg7ivDD4D64SdSIjJc
KsrcZFVJ5zPNDyPpAbDnUJr6tA+XE2bpIB1aAvkrKqiHtt5EiKz28beFF7qbFuAp0zk/RP6i8mWm
dAsoKQ4XQyGT+izgEAiJw63NF6pZVVWFz5C9RW9zlDvEemtXR2CcExgexFtYSeQZGJJmasz86myM
a+qrM1WW6RXdkDV50Bdy8OUNvYUwoZWA97u4MAfZTvg1u1dC4XAFnnLmRuyhGVc/GcYeWqxb91up
ZsSHcTWLtjK4AQHH8EdzWRmrBENz5ZxABAD+oUJd8KauJOl8hYzv/zty2bBmshCtvuHTOXa+Cs07
p4dI+tuNGY5uWaZHl/7Z6ueDjyMwHiEpe1fO3F38gvjD5HUsh9lbEJPgCxQvdNuW7XJpnxdMtxbN
P1F2aCEMvXjIo3Z+yL8I2hBrywBCm1n9eHRllCVSWVeYC0S3shYdlAj684hsSTxjElgAhNmSjhvv
Tui4L+UuOojmqX46nXWZEGvdEtls4EcYK2D1pbNB7WY5IUMJHadSeC4y88m8F/ga9x+fnKntB4sP
hhnzZf4j4Vyhi9hs0DITRLhqUwdjgWnaN1qmw12XypOvrW7Jd2FtLzE/5cQhsQTtp0o5PSwYQ5Tn
MoUQtV4mdPFoZr5DsqsqZvqek+U/AnFCu0rRFbJcOwAaaIcwqoH2MF2DGkjS9TGbi9Xkwb9gPdIR
WFp5q7skchKOV/9GiGgaPcYqSURAOct9IrR23MAvVbTPO58lA/yjO+dOIs+hsrL82rC5vxTjgwWO
s/Z00fqo9woH9HrzzVYAGumSR7wLvfmrWPx9V0AoAgXpvVQIWzj2ghWscEMBPJPOf68gKSLA1gpe
iFgKD4ouiaExucf/GnU5Fxu/rtVBPcuYniDdWeRJBngOwH31twKniYsVXb7mbazkAl6B+mEkuaD/
MLNCvwBXCgqefVCjZaWDYfnFBQ1rDvO01nmVoD40UlYjbqckxJldLZ4oyoBWnru9GBI9lDsR9kV4
X6iDRQeFLDASzqxNtrFjLKkIt4VaPf5TK5q82KSX4GSKc0jN5gXZbU5hjuNiakVwqG8diXx+ovhC
+otKnt+uJEI1NTdgftiYKLruxsY1HGaUtW170RY+aL3eVYUIEx/hUoNrMhrtpnkyysnfZTS17tbB
PtY9RQswwnzpRnHWIy5Y0O/HvLmNeSay2TBgfwZNfPEhaMKvwE5gw5LCrr3p+MCX8wKim1+ubpLH
PXxMqwawdku6Q3yH7MN4SPCIqhwbc4QrSYSqDb5r9sbnWn06kVzRfZL8M+La5m4vyW1ERxDj1DkR
bpuVKg2lqopEmnx5d2ypRtNvQCbCGzZdoKfFjBz4OeLkuAkNxSIanehwtSZe7xTcAy44HIWDxPM0
qBwXDZWd1v77DT/UJAFJHIuahQYY1TPHZp8i55KY3Lg1JbZcSZCi3lbDaN35zCcxGaGiTG3DUF/z
yy/XeORUcKZQFS7/V2fCXMrkb/e+slcAg1F5bGTMxKcmd329EnVaE0tY2sJd0bU+wddUgBUkYQSV
E1vDQND1lmF0bsJQz0rKYrKaxlI0t0wbvVj3xQ904ORTUHmvuIVtTYpp6DcLNLH6+MEGVPWRCTXr
ZxXIH9En6HRF7Va45H3hpjf+5SfvQY8QBa/q0f9UJvrNelsCgyfghNobqSvHtZfKvy7llo/Iml3t
P7euQpKFGMkqNJ6jOsEJXohFLsai0+BhjMM+b9Mlzc/KLPvtCJmIv1hr6nfEnu8HweWhmXhPafax
7wXFQgZR6rpictihiXJxMUPPfPaenFtmenedPuEXhkAJAYBCNKL3AihreBlx9VPElVRpf2a/vAY+
Liagei9wlJcP9kE90HdEYu/ZWOkGMwOteVboX7XeP9LqjC/FC2k0EF3d+67pLu9uiecHOR/DNIlN
XnILV90ehSbA/wsmQentt1Vk4wRmJZlodmr7H4OHUUNp9PSBxWyIOrGQxsjINx5uGUZyXLBFH0dx
NDfCHqLWWVMXlN0XqlhKcY5mHpO7kthUf4IP+uSQUUqru9AngzsQxbjegWZQTpCdkElOlOSX8BlJ
xUb/JxzbioiwetIO9IUhJmPQBMAp0pQc2EbZxCWnuqYtdDWtcbcNyP+KeH+5PsBL8xS5B+taV5NS
UnJmbtTB/mX612O5ZVu98w/tOF8uZjIl1aFuUa2gcvZd3HhkP2uiVOwXL8fvoASbi7nmc2v8o6Ut
u2sM/ofU4HyZplHIfNCYd/XOV09ctYwbvywPHocB8mga1vZZkqhBJEOexljQZDfzM1KrZzqV8atr
t4S6HqgHlyWra+LNlYU1tbJ2mIet+Yt3TW/pp6M+1G3Qulhe5DMlIbFDam9kmd2T4YLwjGPME4DW
bIgd4OTbVe5Xc7HoEVdQ+3tL+QI1ZL75dUqeHhegc8HK1YPhB76Ab0wldaQEPHmB5nSIYTaaF1/8
BOO/pC7A3yE/9KQhT/wGRpLRlWPsNQzEepdqSJNxuzvZENxkPpr7KREYmZeClTzRaJqzMbxBir3x
805grgj6fCGjbqcq90SEp/QwtwpuP74CFFOAdCGJCWoZmFz1oDKkHV5sUJ5qSuUy2jx+xyEUBKNA
HI76JythlUn4CJDIlNbiCVpl/3U9lWUfGTXRuxk8TTzOBTz3gdyjK2oAY511knYw/rQGqbdbnK9g
nHp6KECilmMdFFWvX1AfnqST7y7F1xeoQqrOcNm78nhWDacl6q3UHrcgiO2LdETr5WmjPra6D+lK
/j04un5pn3b0gLB3veykCL7NsYyq+g0kJokVpFcKizLGqkRENYhWEb+ZmVSCcKn1QThe49O1Fmth
rqXPMyi7UQLis3CSlXSP/TCGkINfZmyOlLCCUXfG87huoma8AjA08hMWtkKe5KFEBJ+4SFbBYJ42
/KsSPyDPANuWKul0DEFTgpn/mt3KhW74GKp2uR1smUQVYDzBhGfUqnit1gl4XUndTmylj2u29Vbz
MibuveuEq0yaBARQnoNTgjNqQr8gsHq7R8lU3Dbq1dE0yBxXTxd/qJSiFuxTI5/81YQzT3DZTrIn
4eclbn13LDw450A/UFda6aBR7XP3yYOYaJKeZVzaHs2TJxs0IlxlOYQGCIPho6TqOIMWHRivDONO
+k5+kyaEWtvNcjbVITgYDDBdtRatDa3Y/PoX9uvKKD0adRHrD2LAtrKb2DQA4HO3ZMIKatGZjbKN
jpcTmf+cyUEDge60IiTz9FMOxf+gxQUWUTsmHfRZBsMMH7kXswtY2pdJ3mZ7Us9cKhbLcA2Ma2kG
ctMPp7fXrHcipyADILhlgfmQpPDO6HEhdgYRtHDpKv5YMJguoUbkXsvtQV8gtA4xLRbLgppcZh+/
tJ56RCp0BmUfvvhd8O2ynTHkTteDI4Wb1xtBzsQ0sxSeTZM9uNPtj4Rmaqv/vLZfHlE9cc6SkT7f
hzN/3a8FFS6eKs0OhaK7Qm+7tC1uw7VUW+y/0NuQQDhfYCOqr3D8RibRQV2Ibb2wL8D4yWoE/FeZ
GZg8tEbjqKx0qFjZdEDAIu28W6fznfil5Gwa76I+OpKPZD8dcFaZ9v413gcJTjzxI8JPlhkokmOS
EyZJEhLcJmTCwQRjAdgk9ttJCK2r5uiWE9uYTLhO2dLTenQYvHneh/oyxqLCcD/380C+DrQitiFG
pqlgcdo4gNsXkMk+Hb6yTpY7Hmn2eNX9x2tDh2pOicQ08ZTp5gsCpuFGTL/HfgkyF4JcqrwGhfQ9
cjtmBFlmSqD1cj4uFlLq8PItHXgniCqOrK92u7ngHCfjdoLZXqwVvyzfuEB0iYRM7OQEnEIHgv6Q
2tqk2PGU3mrf8r7mW6NH9A50z0rq09NQonuNk7ef1muJiHFjiFJa6NUZKBnVtEivBwCXQDVjiQwe
0E4mi3IJqe6aKod0yfN/kFAnt9SMXzXR1LQ71XVE18x29sVbQl69x8tSz8HRff6gm/AdVhWgU2V8
DHN9SMQ+fjAgCXksXkyiK4I0RrhVThSxotY1Oj+99vy1bwu06+3/c0odGcUvvRWTXIQVdnQ20vuI
On7V6GR9dX822wbvO9zf9dAwUe73MpGRVp+MbYLh4jM/KOg7XlHCsvVQ0h5CbXdaR252+eg0usv1
0OBjIJzLFq92+LZmCxbPwB5M3zO8Qb6silJ91QZZTfHPWpRJLFNZhbuUNdYgmYUeKNoFQfGtRtut
0/BmrZPzHZ61fHVQVPW8jNkrC09sPsJGvsowL6EWCFYppLGBXtSD9gru5cZVP3aR6VPYzN/MPh7M
9wX6/BCaNS6gywkvoRro/TDDenr5B7YNPoUvt9v616R96psXEtJT+OA0pnO1Eapd8YVNu8p19e7e
LQXD10mEI+WdGc6B0vFqcPl3AzT57d25CliY0d1xGGwgQUqCQpSqdROA3BuDKnGzhfPFYDo+r4dq
B1UCOn6AQSZPzsDqdrlDIlVMAnuSlX/vjsHMEaqyunMVxT4B/4mK652E+RRfIhjcjozd9mTKno52
5KV/sOifF0nOdE4w0TaybdMvuJb7HtWvcrAeI+rM4NjS2ASFZqpqGK8mdfGBR6UDyUnUo8Occ7Az
bDGMqYgCM007JA3gDZMdz+IQFfPrHh2HEfYE5z4rACrE9ANozP6gApNEzhaj/3mF3nSv82Lk2xRx
OaEJ7aD8dlgRESiZRk8pX6oxFCPF6aHrCX0XOTUCKThFZIpnLeXBUHd6Z7tUMVFC4EjmbH7gUbeO
CPGnAYicI3oZPNImU0J0723K+Jd4KvjrWSVI0fJyHy/+1rsYoPXEITAYcuv59p3sGfJ6PC3ZKL8/
sZBP/Z58VTN1uMxhiZR9vyC4DMPDlCI+kwFMcsJa14Noeyi33i8Tu+dAvPmupqzvY0+BWo3XIbsF
OtL/myQszfXJmsHkeDZBN3obCfF8Iy2zyvnpNhk9bSwWmsbm1QF5dVPgexxsuEHgEDFcgv3ue0ke
1A21n0TNUWb+Gf4HesawaN6Gx25hiTGs7PSMtuflMsCk4rLpG6m080F+z0i2eOFrzTO9e7A3daPc
uf5yA+cf3mQgmRGgc7IgNdY+NBtF3hO6n+kv+MlPoP7Q5OkcuziSfd2a1hLm2Z3VPBj8yMVJl0bL
Ll6DnvP7QRVQnVLJ7yVbj6kQ8h4RoRLRSDNzseO0f1JZvWCPa62jPDP0iFgRc4pV7Xe97Sy0AM9U
3HWyF7TnNJOP7Ntw4dZHy22kjfGqvaDnAqNtpTw6/LwjP2tL1fM8pzcAu8WOPIGpv940+W1l5jcB
G97zLdmt+Nva0PBDOsmaVYJWNIyYodEVP8Gc6zizNmwlWGjQpp7XRBTkv4mMRRrCVD7NSOK9ht7y
NKBdvqNVG4uZBIXYlQ5QmFWd2opU6UxJgHvjIMjPMpHzwS1wM7cqSoGu8VsqGEh54sX+57g/759+
fmwzlq5mI2JPpCw/KCv6/xAYkF5lnJ0pCWloTabpPt4EmsXegyyAJWF6oewiPmQ8iD7B41cmrv8l
or5BOEMe1fv6SVMY0Y6k56jq5nqdUxtgMTdARJfSd7JR8ZqmWwru+SIRlr6dZtnSjIGPKn9hNFx7
2RUC6bn/X4Xw7g2BCHk8dZLU3c0dEtP0zOkbQYAn51VhVwMfRPovzSrHW9bSVQgcuJCSiPcGp5oX
j4onhsmdikqZVYQmvuwlJ8Gh8Bt8AvTMosde7CprkvA831+OFbkQLtxu2DRjIGW6GB2jE9WIuas5
qL+h/QMoU9/PTv3l5sLoQGPkIe96ZDSdlA5Bws4ryX5x4sUv2OM/2p4h6TPf2IeAu99FZooI2vGY
YYRy1cXZaTStod/uIwlfEYmFQc6U8IkZ2NVpaP4AgM1PoDDDkZPt3SbHEZTlOE4CqyD7o0jppqjE
WulZFQs9gr96At6+/2QCMMlsBXGk7UwUiJjxADfE0SMOTY27VujY1vnuC/Ij8EEvXp4aJdyDJgXm
yDXoAzKuZiAPgcHCYKjir8TelSviWc43PUEYNDRlgGjNLWVym26f2wib06db1W+SXO4K1IMf85g0
UHxebbVLA11MlNfUwxXlV3/wxPopPoY7AYFA7Ra4sx57Rp94IZgvu1DEqASN2VQqHFmWRqAVWtv5
/kLpVteBojaLeygn3Z/J/G3GtJkOurqe33+oB6w1qZUrVMNtcrJcQmK012iYZp7O6bh3fe/tL1Nn
3uUtzE/rJ0/ishP71//AQH7NbIPVSecR3Gn6cPcWWMM6ZlVNvJ9fYN3BJBhJZNg/YBnSh9VhNhvJ
Vg++2MufWEdCwFpgeesk8pZmmYK5jrY3COCxGd/hekCjKVwAyB3V0KZpglTkJhneb/v9OuDo3wI6
qKUkZlXSlJkWMTMXnMawCX3M9v4sTmowXsWhBiA0roVrzuYY6SsybgVAWZ0D/dy2C2Z75fwhgyMi
RSlGdt7is0jCn1rQ4FNoFqzNM/H/qlthOVdIdo68RwW/F3xFKCD+0slH8i8Jl47wFB+E77rfxzp7
GKjoZRaopmXS7+8bJZV07uUA51vxpcMcWGVYFKcDjuVSd8wS53MyISbR3KOxupgivZewhb7SafbU
3e3s1ya13qqru3dPDiWkg2XxzlHkYKtQCwLPu8avjv42/77hh6g0XoeftvkhNrgAVDXqn6EpE6Il
wzmmOmXl7mFpzULzsKkm7qA8wENYFQ5Uss4O7jt/YByUb2I/nsI7VCjWnthLW5apW6Km2otQF6Da
FbthBoFiBCEYtUwSZbvMwAAy5ol52XE0r4KLhzvvbcQbNHXQw0KcQNogoaeR9F2wGtFbtXrm2vy0
G2M57ulKgEfcSRedNeRRsYTbVjgFcDbZndeA0SnLYgqRastBVQ4oF6xfGVjPZ+HS30L9w4hkywcB
7rZGXMOOPZdvYJXQFHUVG3hzRwRYv7u9zNPSfzA1WFC4eQG5hMLUqsVJIeDGxnmpiC4ds08VvsM8
YZ7fTo9XMRKKiLSVt03Ws/p2oa5krSMCwEkjTh/sc0mkEvRRMQYZ0gXVAYUS9fhsFFTn4bOV/Dcz
5FeyCvPUdHR9bT+8c2Og1zttCW8otNKO8mDt9iFsr16zla7Py9uYFO+CCbMdKRg52txOe5Pvw1+0
1ifdRiZxqtTJZ8pxnl8NHMoJDEUo7QPNJ2vKIPTk2cX+vTN9BxrAZr/1cwNzN100afrEti7foo7g
r0AoK969XgwpZI2dwi5kEPXVpPrbNTMAyL2+1PCj1z5jm2P3J1wyuCfEseS94mV8NsCZQhhZeV8x
ZzRQzHx8aowYucANLAkx1ztyaIQgDvNbeb1ExC+sakujDqBtfWM4mRpDx/osCfTEpwuH2wb/kUnd
rBEo1/sU//sqwmPHsG2LijWEuWQCMGUMqmF/PVZRr6b+2nAxIgwnNFv4ru8m4M0w5XE5UAO2tp26
Lf6P11PN3nYFBgTGp1n4ybXtVnvXg7oF/IXPJ9wOGbs8rnRk1K3LZ3x/DlkbgEHsVGgqk6ygEQPs
oLRrp2JW+FxbRW9kEugmFi5zI1u1OHpqGtpTWlN22Jr0pY2RWjKT2ghr9K1UH/m1ezY7ODeD2vJl
UCEGSqE9pKNLELj0HMCYLBZ56aGT21iOihoYPis4A2ftwfVrOHhU3JSO8nex4po8UMidxbx103hq
eDyA8jjKjfrrUvx98N/drA0oBUdo3eCJzl/0aZ0UdzYus9Yo189XaVUNt0AuIzSaJpPSOtc7G1Zv
oDO6bvZCJQmYaeURe9zHSjpxNaxDKQdpLbnFoaWWg3/zElPRSeFm6wEISofZRw3I5LTTNS6djohF
1v5lfaY76yggJ0szpE8eHGP7RDb8QuQhbPh0ner9WU81uJ1abbhZ1Qfww1z8Q+VTolODg1lxHnpr
cjVMH2LXxaNV+H1FZbWTXvEVxlQBjhhE9PzFeHpTWxqhw5aUl/kT8SZD25SYouDoTLeUyJuCOG5x
ihIWprsnzPUIWo/Sg6+9/1LrDFyK5Zt68Rbb8zMa/0LZPVCGgsZHw9zlVbtX+n6T2T5fdnua3Nsm
WLmqc8tmps4EY67rk/dyiCHYLP0fVKXUrO/vwPH2jnCfjlQHRDQcAnJjTpU8t2y8ov2BjpudJFvz
VN9y6iQzsVWDypvNfIr6mh5mdaDc5Bi7KlYyaUlyC1SwMqtiaqXDzj6nY1J7B1MQGuKevHfgB/8q
nguchfoOrUZXUyi48Jd2QnMFSqY1+mMhJNl5JeRsMjwECtZilKhP+lPS5ijrfghL4jAqp4g+Djp6
7W1WLoZKhyqu0HObQcMouF4WkQS8R4Ka0CkJsOSN8nUOcL3z0vgo6YGCFEaIhNshis4wfxDvL+zM
/6BjnVpFXLvoKqAJPSLi24NjD52kOjI2lwF6wLE/y0yHNE43mILWUznL9VpP/Db0uhyNsImJqDm8
NdUIQi0C5H73wN8noqGKa8w1/T1EUz+8H6zRCtPHOngo7LwGvLRI4JDPVxEwqDgTwCbcmWLRNmQ8
pPmRXihSTKTRPs7VXdQketJM6AcXbznFH+5XNHYtIrEtUFCN0g+O/TCbExQHRr3ZxFyYd7+e+MNf
dkcZK16z1JOP2t/p0hvFhF5UiaPD2sOuzhO+RPBXIw+qdTzN5oebhsH95GQNh30R5VJMs8Y3z+Mt
9ZpwN2V7B41pQzVAaMF4TR7jun5YNd/6MbMjjY5ICnL7q6puqjZRInPRw6jnawNOAXPCL367aCGZ
7VVUjVqYOzTOJNMk2ukNtNWyFcjincAHOp+ZFVbGsPyDCtgPRYzH1DeiqMjiWnLnI1fq5K3YZ35r
9Bt1SaUMkE9kewEa20DFw83/m5+0gyUDh6Dtj6ejurlQuQw4tLOltyEkjLk8sOEvW6UxX6mlpwZO
GswmtNGoJGp90+4GHWYEa+induPHyRm4JWu4QHe/cxxMFG097GdN/6pbF2BiXdhGzdczSWRAz+eq
6FvE1t4S0e2RV2ilPKdVsO7LcFeivuiXmpYbbTEaL7/TE+9K15GXxEUrTkCBwfo2FvaXfYjALIX1
Y/EYx4WsvK7TfubAhkJNJa4rnvD+9RvGc2NEjdSiJUkB0CU3LahmxZ3Jofaj+dIUtN/OKHq/WNVE
R4O+CjXdenxaVkRnmWfNhRmSGOIL7dQml3xvLUfw/ama9HOmotO4YufJozmXwV3xPCeh2b8jAgqP
qffT7PmVwgPaO/G39RzHNcrPKaizkhEKT+TgPcJUTmRyB2xtviC+XpnmIpczZmU3NPEMScoGDoLM
cycG06NPOxVX+tBe6uiG9kmu7Ip/pRsx4XmYWA1XIgA1QZEU83Z0NdIpC85EMxE5yqBbTqC8Cdyv
UizLgHVh5B2VsE+fz5Tgmaip6xvk022LBrAeJziNufVC5iYs45fsjy2gslo0alsF0uqIs/JrdhDG
FLdaxS900mZ3HFF+9jen3WzmEXeRWQY5+95qnF1fHYmTlVcntmdfCYzKE4Dc7e5PbplVpVDw9Lk8
jvlXzlSB3OURhiyFpOHm2qBeYdrgecan9TU28pnUjqawzFOGTvcTqGN03L12TW1LRQn/oGZJnTQl
eVrSv6Q4CSEIj5v/ZgNas4aJq6Yi5xB/4mbrTRAgTH7aRqvW1jY6l21zsy3L9GcXWbuylgMNg0N/
AwS7haAJoO+pvVkiBZT5CsGwetiDpI3zme5nJ07reCzVQbN6xq6fkgaVY0io16lXGLrTiPAxYHew
uzr5zYy7xFCMCyjrK20UqjLsyRTZei5Mm3c/57s6o5tnWsUQ+9haLl6r2E/xf/6JTePxcST6BoZU
ovVeQLMZqptcUV7RShVp4XUjsSZ+2tTc06Qc7kfQdOynMbQpyXWIDn4nrzHkzRzpwTMJdaXYLchu
90bsrQ4nQZ30upwLE2IVg+vNvLYwXudPleMqils4aD0n6TZmU1qSPrUCawZg8t1Avh3dQ1iaHCKT
jHPp+Ebozo6QCKPawkE52AWM66mjxvVRuZ4rBHjwZ3jlJ8fQ2w5kdhmtSzRjBZOgj/uPkHmXVfxs
bOWRvtRH80I40Ge2bIbVfehLpo9NnBU/Jr2kWduceVmXhsq5Wa2Gc+/33WJxxJFqqLOl5z2NidRe
Y+wYPvOO2sF19Zgk85elGejaAUkFYEG707IEg3iENNmXAp7ORju+eQPXh6KtvLGi/NztBHyj0nUR
WNiifkWahJR4O5xNUf465j46Jfue8Ufz2f4GHpZikbNdbJMummRl5nSH0+KIrEZYdfnthabgsChn
UT3l/KYUP8pUzrGvhEted0w/5yN/0ud6tk/jK6QpN4axRQZlv+tMJubd38ko+LvtKgohnkqzX8oJ
e+R7q4p2YPKx+y5SPCDj19XQqIxh58tI/ka0N3IAt3fnSRJXaDL1/xC5u+8FakJBYYZdmFkvTqGs
EykdVh30IPIz9gvqgZ3e5fvHbEyioPET5PFGL75Qt8xzXeev0n2ZJdjeOCWpUopiwkH5UWDV+Dmp
LRz0LSvwuwwHda8t/kUcbYDjW4YoQqJCChDga620l6HWXiaJcE3nWbFnYw4ry22bKkLUCDaNKaYB
B2X/L0YdZEbDIxqdbDHoSmgZIVw5f90aHmz3QgwCO56fQV2zsHFvObSAeEyphZ+kO1MVF9fBdZ6o
YLb1EKDk+2IWHY+RqeAX6XjYb74AWoL8xb19zq086R/Bt3QVB+sy3pxJjbAhgmU6RNiqDHeW9VOx
1qI08u4VNFldt8E4aRRRxOKpT+RC9UIob0A9cRWRE43JxRTbYH1Y6T1iYUQ15Q6LcAi4uIncoi2t
aCud1/YSeV5a7t3QF1/LbGeuruWe32z521dq2VEXpFRHOX7+fKCoxFVOA6m8jL5PE1S7JQ4JnI2q
QLMn94iMDvQLNytwB/RyVu4GkKeb1ZwJ4BE4nlr86q6FmRLV/AAqK3y5i1gGdnc6ebQju+kwOdQd
HmsjG4yz+LCYIQr2Xi+i3+2bksNRxmv7YjVjlZ9Y2rQ7y9/vD16nbCr71xQ9UVVih84T5BoXA1rl
Amc7e71Ibfd7iaapB81M6yCn6amYu2G176Gq1oJVFhgFZwxPr7KDKbF7bXkaWxwNZmvA6YV7N85N
POlHurztuSrWaYiF7+Z6H8QRmGyrQuX26NgbVj1dgqRhUIvTyhWK+EiZ/RiXcKEjvZ5R6rTuq380
41+Ux4tyu9Hy0+8V5OP8gKm/9r/WwAlb0VaFH7D9NlM19KkQV5djpxDaaFFDK6pw+jtXcJRqz2dw
y+4r5RfkP1cQjyhS3gZqjOqIhhbNubnYYBckauD1HjvN4g7fVew7D8FJXC0USSLkjQDVtu+x4KhJ
2RxQ9j5nFHRjgA+caQK4GPYyCeotA9ZMQDojfBTEFHadl8um2S20dgy2Oqp29EuYmetHxzXHWudO
NifnvTXG3Jh2S1ulf8rNa3TfBOuzjfJBEquscgcECQ3GIY05RiAYxjoghr+eoGS3E8HcHvd8R1DZ
RUXAFtjqv/K7syXDhWAAxEy9gXqx6t8hPcSQSMnmCpAODvijQuL1S/vsK4uPV9yFPhNtt/AkUZvv
nNpAyP6teFKzHxIyARuOjlC6GzpSVdt4J/7LsE0lqnEQe8sxfk1VFKkppOvMuMx/qkTagr+Pn1CG
E/rRLJIy0qQ0m51NZZgYoTNt5RJgXQl+E6iBmH1ferQkUEBxsmQ44xwiEs9C4Qe7Gu1Ey6b7M8EF
nep+dBvcTM+YVYBbhKWv2eqdyN03EGsZmakq4utcSLczrwe49h1atPjK0tShFYe3Z/spb9cK2M4+
kJqtOswndm1KFy/RCVClb7uMWrCL6mz0x8DbwczTBc7RtC58wTbQKerAmWO0jo1wDAx2zztjn22D
5LeeKDNZCqea3gXUEKEvxovGW5See1+/0SCQD614F3d94ahVzSY/0yvkIpRSOnLPpwxB0maiptjD
ZsM6byI35mcNQMfgOLJKtTlrgutHL3h007flK/c2iLwknN94L+xrvU+Vv8o+Tdbaqfl/u6xbM7xa
hzbXug43s1uQNKB6RpgKBeG0o+7SI1ib+GFMLgW1Lf84TckeoMNtjSP3wxcGs4X9iDvzTKNMdKz+
X+pFwRem2mIWFzlIlbzj6sD/gKQW1AedVcW4HAXhpT1f9A64r/I1JtsDbRM3YuyhRPp9Ublng7iA
jSXzF99HwUw1I3wrcyU09KNZVXLoP4H+pAwljLSjxLsK4MZLnyE2YljasWPkHPGBfB/ulaGPNVZZ
8janfBzCSOEsrtiYk71vF/CUXE/qHSJUaacuRFZ4S8t+br0dysDvBE5iR+Ggc+qBIutVS1055Y/u
UKmDFBPEc0zUjrxp/eiISkBSeawZpa5LQT3v3GXde5rMEjaiOGDYZ8pO9Cqt5//bdKz9lcVlA6Y+
ToeJKmYSTXVtCD79t/Z1nR9dy8nm4BCeq1nDsGe6vLbkM1/DeuWR+YzM0KQihyvQWltVmnUp3Ep9
Tq9DZ2s2GdOLnGBkG9KWyM+rj1etnZ4VnjV+jwgZPMAphI/+cozlq1ajQ5LbarrMuHFKKCg4PAmU
1OUA2wyqSozQ4nv6ngoSc3mIxck+RSn04WGIyF4gB7wYWSrtWANxcdIDYM33Rj4Mxx8h6W/cTABl
0pUaPsI1I/Uuar4WEKC+6LnzL9jkS+i2P9zjlkJeF2S4BM7but72bbumvXfeCm46VrVivNFzO68v
XqLywaeS/T2NRzw969I4KsXin4ONsgVdY0bjGnY7LON1b2KKn1/je78l7Ry+Ov25nvXGZm1jTgLP
vpM6ddtg0WEoGxv2Kz+rO3GkuFO3bkTH6vHGSEf5vuWaSj/wa0PqM52I+DkuU7corz82zpAmt1wF
kFU8QzvBEmiBP2iYEtBsAwTGXdm9G1273CJZuy4tlvPMdBrBzMZejmT1Oy9HB4NYRIfxuPZmWyEx
0nUiJRqU0kh4+KDeSppxoKHoFT2/S8jHj2rvUJtPaPg95gXmQIkDBSluWoxbuRQmtaDiBgp1h09s
nkIT31YQsxQd6my60zhqVOz1NNbb/fZgcGR6B6AIY3izntuH0XwFmJMqnVSwOC680Pyw8nBkx/k0
/jgAOrKK3O7KttOnu5BhPIKI6awcGkhWLaNMJPdvOr+AIBz7yij+vwa0uMs51T5ZRJeyqmgk3yjd
cUCC2dPfB9ZxUjuvWQ15lv9H03FZhH2azbR7K1ryaoEs+k9TGZu2LX5PQzw2iR9k+TdbyLIc8Fzu
CeZlg+n6ZKx48ZUgdGmpBSeHBVlR64D3Su3XTTKZTHgwSVHdHNUqxLvn+nc1P7kT4Cxhj/d3y4ST
VfqceVfExiPK2K+omLAphYbefEva8HQ7nOTqHWMn8GTJE16KgscTGGxkf2dgwS+3jl3ZvqQNPzo/
mhKfVrzxUI0/6LIsVkMGAe8pPvlel8dEbJA6PTIcAscC1PUl+JWcAztGDIRidLkwW6Xw4NOGfPNr
Cm7d4KCQ0dspTWQS/T3xr3nMW1bUFzH2Ndfo5OLsvMkg75ICazdwv893MPV3wIz1OUNeu0WZ3CNZ
T3cRssobPteGHlLuaXKU2VP//a5nJaTdaLWfIwBHMjd7UqcWjevQhp3EtCn8AoSc/EDYJ6KBcMuS
0PbzXHru2lEtkPPmleWOZymbPFnXA3CHFPbxNuynCuwTsxi5n5660vU5KdaitjQlHFI7ORCM9wfU
myx+3rs6aBZENLsAXjIXILxjYgm+OksDk2sWvdCL7/ZirKO/TB6PAARUe90fTgxXj/WENocBtQ1v
7Azi2EZx/VfQrNiu1wp0PH2R5E9tLzohzVHeX5b4jmRKYoUMvDeIGYTbZLfcXdNnH98Ft0nwnSZB
ty5j4gAvCl6haPLDKyEZxjVas2ksO8nRtaUSgvfAxWNjXG0DIDp+q7i3AdUoHKacof5HWRXqF4OP
qSiCM+TrBzPF5qRsidwEhIiFjmKNM7VkGFSO8Yl14krBsoQRmvpSZUQ+lQYAtDF6mNvqfj+wKssN
X8DgeenqB8jDKzzNwOnt+yBrepgibrEXb34Lfjb2vYMrdBxzeapxI5exnMvX2igUD/46izd/I+pq
m+HezNY5vX9m1ve9AfW1ZuTZ5P1xYQHbRt3gB+2m9iQoQairtsopwGrS/0x1wtoRLDhj+tSa1LiI
zub9fijIntf8CRS5SS7ZMjJXZUNveKgMsRrl4pd+k4vdFdhOaHZ4wBEPtMJoa25iiUCF4GJyiJ33
LBR4SHW7Qx55NZCB/a+IXtp7WPkbjnPMIXQUJtgDimON7OTqJxar8twZCJgHAdm0tfadfG94menK
vueoYzmlRZYIJsspX1Llv7gunxiJc1vpRvnVB0z3TsLs5hBEs20EZ8AfVkLQWnRABjnN8AZI3FQq
uzJ5y/8TP9LhW6AsatOSPbQYD2TtJ9gCf92MbwMlOwRQPQIRNnX/B2vqaQtSs+AtWlEP+pINjL/8
0vsR9N3bQMZTa7RcwjRX0Ri0mEW6Uc+NPuar2u54xOx568GJmVO+RDcQ4DLDE5AfdbrBqRS3AxUX
IMVWUL2D5ZeZ8zXgasKXp7hGvmkhMo8nLXYL+D6pkSQtOIfxC/nCqTA2uHWh+h6Y2W/7DJWvax9X
ZOJHN9sf6LCTXCdcTJIlW52XK8KwaiRsP3FOvzN3c5NSmsht75xSnIFefsz070ZhsczeM6PbjTv8
3BfW2xD+8/hK2uez0pltIxpUXCZKFs6UhreG0N9VBxiaG0u1tDobgNZTeDwET7WpKRAZS7Okroh1
wE/d9KSHJBqvwJGvqz+iRjaY6CsndxzFviaxaTjZGoz1uR2ozxz7OH2EnkGVp4jS83zx1FpW/mIw
5rNfv2ukeMt4VWlOfbFJc3wODZ8VnIAckXQzOxfyQWdtbFnZuLCrCfMfRgqFfPL4noYmwLptuixu
mO+qK+ls+YNtCzJpUFlSFAK3IN/TByID0ghimAtwAFp/nRsQhlnkKWDNEjIMg0RtRGDOpjwx5Ot2
ZQhDTv7hbpTJBj5WgkE3lxYaNQvDtDJXbVpVsm2EOD1YRJYQ753pXwnStQK1vUj89RrBRPb5rjEB
TdWsfbOsr75Cvanhl/+QFeDO5pZBo4zuP0DVlLgAEZXNLf54NuvrmW0Jgs6kTb6xFGPFtGqHDKXX
Ma3IZsaDuMFZO9UWphTZ3QHmbHC2qZy9fK91YmWL5T6958wZ5OpTDMTRD/UGVWEqujMSTprGk+Q4
IS1XVyPq799x5CB88KdPeLLOI1MDzHTIbLA3PYz51/Drq/tWLiIRyVgWvkMHo76nlB1tthrsKLLu
UoaFl9rEIBsd7DgiKsoT9fX7EiHKRkzehhb+d7KJwtMa39uqcLi/poIiV1E2Z30WgT+3zYUlENty
W9WLbuPaQKrCiB+JOf8beROOeH7p6LLzkIqU61rS48OXYI1MlCamNxh11LZc9G2SBhNT+mSxuxhP
iWypkJ0mK1scVSiK93ca9prwx2HVLD3YzKtHCw8e2Rzt+9v+iDhY0jjmg5Va2jfOxzDy+bDRSmEY
zjJ5Xn2aQmjL/DYhW5iIS/vp+EufRc8MmYZeHrZsJYLT7/0NsaQwvsprTTxGxC81jdbPGkMj5URv
00D7GMXoXSY8R9tw5CuIpkpzIEMKyLpYydZzX9tM4RZc4XyLTgvjuCINMn8Vso7wCUv+qBmCUM6M
6SXo6hOGgSIU1E7iLztQp53sVVuoSPPGhS2+r3DXGkMR3ZOlSRAmesnkTy0yUu+VhRSfXFW6PMa8
06pN0oXQCsIKWt+C7+NHf0aSS7i8/3FengM88TxGoAAPiF+EkG2ZKsWOG4LCJvk1JpMP2kW/DHdB
1Q9JoVNQISynOBAiFn9uzB3j6G30p94WoiVsRSjPUFcSMmbHVjsDslj3yVzPI+xHqkTudfgYg/qU
9Esslr9QY2IApz6o4wztZnTK9oXGF01GiQAZX1YLRXYJAFUFMX8sxhOCvXAvBYp63AZcN0+5LjeE
TsmxMIc1TsJbKLmhKMMkBonfMnFLloDzMQlMjQpnDtYah5KTLpeN+J2SdqozGgg9ZQvUepIrJJSZ
DffcmZBytLttK13Ey7mdCOHuQib3QidpIpETtACaB2+TMpQzo1PKMA5YUdn7OPBGGrsGjp36CuPp
IIVpM7ta4HS5mQGG1zMw06EnKQ09KFK/vM1OcNXP6It2eW0t5lbp7VE/VBIh97oBmqKLIYzUjeBm
u7OVVqKw/g7TxRPSsIf2dy9tOJhqv3EmUKgrZvpn/Xgpbud2n1/CSqzAr59pxJfh/WTW4tyAXgz/
q9x9oLyDceaJproN+8ccsqPUFlR2xBxEU2vpAafVJsZ4d5f66j0DN7X/FWP0uQLIkYV6n/pYjPtZ
Vv5sX9BqCUM6AFdc0JLTIDrER7KDK8LFJ55I1QavvVZBnyVM7cFn8h1Yi6JTFRyySqA1dq+sSoFG
qwLFjpwum2Q57ysW6HD7wd6Dho5aVlLyXJj08o0Nu6hkVFPGRHdTM3XGj/QYU2bEFqWse+lsqqjH
l9aqkf4DrYEMqb34aMT6sfASzb1qCl3z+CMk0Fyzj7yCCf98RGZ1HAbyjK2OX4Tec1MICHzoLCAi
1NAOYVO3tgkrUo9OYYGePli31vcNjt0eR4nWqxJnrUyKMmjOElbRhhYxL0cJxlhh9R2caU4TL6Dq
VVFueDx6fUIv6uEm95rIL63wn8BvVewtsE3bI4t9NPuB/0/mh3XESeAjm10MIxz8lGdV6tqSqBG8
K5zOSU1YItxH9pKUdfo7BdeV2zj4aV8tHRK9SbxAn75FQ4ziyXOvNwBzTy8gvYng8hHax8uZ7auC
8/jLJ3Ri9F8rz6StURusNRmT4nRLwvKBVkw37Dtf+0SddAV3UYfGvlPPppndDflP+fIoVUqpb6Lu
MSPcXr6nL+YRZsiXjSnSKjjy3yK142kz+kJygsG64x9xNMvSMGbywbhoWGC0YpLPY5clMzCuHKQV
TNfOIV9nSeQEbqEPdHab1kvdZg1hSz+NDCx+JN6I0DCGl7X2lIbJhaOVwe6vSNFmmRNp9xR3Lq1T
11IBqgfV7cAdAq4JXkGoyCE9oA6V15xnpPqkdH8RLy0x+aDZdy/aQeJpVig3XwvnPr3D3rix7tGD
9zGBSFPQEaqmwDRnBRZB8N4o+4/HVsE2dv7X7eoLga2uHPINVzwzxSvE5j8nU+3XxKyowpqUyfT1
PSWfSYasz84797aMmUA1dG9laZUO6heMMn3a59nS1mswpgU/2lR71i+m8/hxmeyRzdenSdx2K2yo
Uz8n4aFt4xePfDt8xw1BmTYKzEm5T91qp80/UVYy5osXWRzAt/rrzmXuTDSyoY/OHS7K2mP0H3o7
MdGqSlwGmTt6EWEBnZnmhkihMsvABTtB/5yxVqdrDfJsSLyrguaNSvLZ2RkRSw/LCB0PtcQpUGiM
oUW4yBeguir68Rru0UftT4EYW6KHcxBmnLBVrPO+7WeMG05nGb9ckcVcrBm37MV4PQ4T9/aVZBAJ
ghVuS3tWRi8qt7W47ZkkBf9QDVB4g0XBWOpiYs+RG+7CLGfpDvBmM90G3GrlhQZzb80o3mScvWod
5FHPB6p21nSdfsGYkOUuQTOfn3LylFIGBMj4zvVBKdMA5jEM46hbEbCMcxsbTvJhhl4EZktw4/5Z
PnnfpYGPnXdcs12cnx8cRUXjD+G62xVuuFht/PMc5dEsuEpU0v+KIsMvgtqVqPVjP1PAZR0W/eJu
MG8/hRaxtcv9DLR1yi6G1g4e5VJCmuTBoVbQFwLMz+4jHl4KKp4T1Xs1ARtF7mf36Oc3rAzVWg80
O1KjmUQJMXW8gStkb+G97+14kYN0bD1HNUKyBDzGmgUAN6r+BN6PhGxY5k9+cGEHtebml+ycfCCW
z34hUx4oUGCJotmVi7qaswBPYpRQSornvr5fXTOoglg7VyYU5pRK62Hi5tDDNyIcBpHOYUTmvbz2
5cqkVb3ggw48ZM8qCu1VDlJXQNosh/NmH+sDdGL5fiYBqrnOHUksfIK1ZtCXcNX16W4QDjS3fe/Q
AX7b7Gn8SO1ma7cm/X5GcdcqO7vMWPvL1d+rjUgfb+5oKwqLVzcwj5jmXeFZ7/xLFl3Ra782GGp+
ncYCP8Zp7GzlH001nh4ed9C+h1DAmg9igtZjIfmj3RJfemM0Mg6qu+CCyYu3nQyBDhhSbz19BrLO
PdxLQpgdY1IDsGQ1EmvtvDchLUk7LdGFXxrYW8p8/seUZAD0ubuysoGUWzS6jNNCwiv5AaYKD01G
rvRlBdM8EPRKvtcfdOiTPgwuI4PsG73aMDyaNVHXoxpB3gDlW5frX78U8sq5l3K9ps8cYw0yAP7P
8WMfUiqyvPvESs2mKjXpK3LGY04oF3X80XWnMrXDIulgoBxKhB62ULu/cf2pClzOpwsgHwZWUlvM
VDnqfET6DZBt0NUwiFa0btl0/f+McZRTJSzXRxpogV/vmlw0e53pPWPeB+vV94g/FCeOnaNERxdS
p95YQV2H9PGac32ECRKg7yxqrdzDVmetP4doW6nRdeTFuvVaIEKHf0WQQIIRlIYxgBqwU5jF6BSE
pEID+UHzYDSwQRvmQ+1kFFToBQ2/UlxKE88kJXbJ2f60QtqQVZFhcC1+Z9WcOf32jivnbzLl2E4l
kkHBJgXz8IUduwz2qAmJPBrHbIOEuXgXurBFZ0N0yP58iKXc5FDZ+ro6L9KfRYDF96sGzp915+Ao
x3W0BzO/DneatmeH52w+W+yDNjbCT0MoGaTl/Xe92Sy6wZP8KfmFvd1qe8BkXCSVhevTsCIGSa+j
vShW1p3iAcdHnwdNq01Utf9Y+IkUPO8Pabw0ssDuokW7hU3pO4InH5DT7EGfJM7JC+B+sBIyD6/+
G+qIr8ETLB1kETkLLzA5iBp56D+T0saPXEoKpWiLBFoe53a9SYvQqIqnBJ2Vy9VPlZ1N4sfKIsvQ
JTkYeQFzp8ZXWfJcriGiFEqj+GRnlnv0OaO45GaFEbJ2t/VAfqWI+3P+XCHNqc8b7myvksgSJqi6
Y94TwUFzmV0t+/v+0IdQhKvl0VQcwUeUInAbcZeAKFIE20CoklCq6JNwiehpQhgCP30d4QjX3AVv
DpSrYn5ynr77itKRkXLPz3lGbfpDbk6Fgx/jQzWznjrctgWjw/CQJIuyll6nMmw7ZVqg1RrY+ESf
CUETKCcYUD39gzb0oo0q69C3LMkKJHssOpqM7gV7mKz6XbMzCQFEPT3GO17insCbvg3yHLNmr/lo
0pQvU//k3fCvh45b8VSalkLpHdhO+v4eousjCsepE/cNJSCOMikezfVyeVUSqdmraqHL1LxFtFwJ
1ZN+WDfNm91viYK6uyLwEKSYzov8NSJb3XrdttXBKFZt4x31knWu4J9hxE6HgGgrH5Lqp2q8oZTH
gPaHsBmKFUrO1CwdeNZ1I5h5C/z1NJiIOyAyCB/CVp/Lb4Wrr6XwuqwmlhBdLYyrKe3aWeJLe1Gm
FBog9UDLabSHUsZb3R6bEil8LjBaAzGuzjrbA88sKcBkAyVuObEpoaJZxPX8sqTECYDmSgHSTsGk
EHfvuamebs5uPSs/0n56TsMSVU9UhBoLch8Z+c4lDyqloHVtaXhTNjKzInZmGS8qcNvV21WaHAbH
ixvVYhON2eK8iBIP40a5A/Xnkwt8ZvMIdyDOehQX7+sFUxZiERtlZbesF3GW2+pedTJrQOfCwepT
Qv4G1mYSPxixfxjo7pEKzEwhHhGFVpaCXjbLcVYgRalEpdDaYXujS4F/HZMCJiAJ4HE+AiD6ql25
VbihYBb+8eY6SzOnMJAkGL2GrXX9g1ImSjyTisgWYowOWHMLxnFfv33ayvqmJFOsENord5hMExUd
471WToyT0EEc8cAsXYqQq1yvV8ylzgjr2g/Oj+zJFuKMhJ51eIhUM0Zqns1mo7xIEFLRe+gvwTDK
ZAqRo2rYL5we58DEIxC/TuuG7CBgq55YS3L85Zz0pau1+yXOGR1a9lcSJQjS3BrysCXGAY/Zx5Rf
yYPUcDkolVNKy39sOOmmz4Y2cMLMtzern+4WIBwJiCdgFaN0C20L2Wm6A6IWDc1/WoTPKS0wBqx2
0xH3ImrsiPyHiFuv0LUDHqZvVmQ8C9kAvxQPDhpapVIqqIQFtauBKm4bPdRptv+9drBPcKRA6iDI
GEiVuPrpbjBStcXVQKkYaZ6Rr9NS35ZaaVqloH7GTpLVHrkEOaeLq9PvvFMzTfW3Orj9Na1aV/+t
w6SZ9NrT/aIk7Q/HeUGLpVE410keG2N4MeM7yPykjUIckGGClb2Q6HpqbiC8qfekXXaZkRzgDi72
L/ea/3qV+nm+6BFFzd8NA0tyE01bP46AX91pWivB3ARKLvn+nmFcG9vBiUgQfGv4fF7m7CSk8Rqt
5rEV8/Y6aUmAwpEdB44dRCFK/HMkD5QCKnQoVzThEqyLRc3YbOGlzTYs9K1jvK/b452hQhiYEcbX
r+jv7OKrZpg0Uf0o8eb2Yxm+h46U56N59ihoQyHxFQdurt7m+Krct64JEHG4kZUYbNgULSRfmrZQ
OgeIcyImLDBx+PnkJfomLdKc14qjF4Os4Y2QU+kVae8LAYtmY8J9fHUY4cxp1WcHjC7fdZ3yn/rN
yxscerl5rv5iFQ5zU6PZ6Rv4KeOHcXNYWsS5SKCQx/if//lVJsAntCnTmmUTw11xnkNFRbd8Nuri
P6XZJRmWnFTZuQIourTm7OqThOOaBBKkyuqxhx6fmu5m3rpiBnKkjCibpCEMScM5T7l1UFeduqf7
NR1efdZzRRRkg0ba/F/PiHWmK7cOHCkxECBvYfKOkhTIC3p44edTVZP8axkVjWYf7di8gaV3u5vs
hEcNeA3ZrjTcgnhRmVmAkBQ3kcj2w1+CYO/VLEfuJeIneKdcjvaV0wrSHueSlye6wQbjcvkK/DX+
XiZ7yYDQo5MJp13M7lVaM9813T6jf7CHcqdqNzEfSiR/yfxMq8mBREE6968w4Z+zVokvautysP0t
T8xkawnjhubb257PPGM7zPpqcCPrgZHY57RtG8ezLdpXl70YSWo90jKyf/jLsT3bG8jkWfi/ejnw
jw0SUvYkKEDKZd/kdz5RgQwLAnPBx1GxyQXLBSSa5brvrWuNmCDcP/9dLFrj/tTZ/clOgGIRMBR/
wBRzQzXM0kaq57A0gGh2WECvNrFEWmC7WvIjo7re9u3kN/5u7woDpw1SQ/NEv3MAraktLP329pj6
UWlsmcrXmzeTHOYSwPevWV14qTXZ26NJELULQbZmZqnu/8F9OMY/kWymSf8UGsnGhl6gCh+2LIG/
OvfEqeOYJMMgpSMI5ez0nIdqyElMlEj6u7cQa76d1KwE2jfjo0nZ9KSDd2AcDTJQnmvNVppJhRd+
cb3A+MJR5Gi3Jg7wadoQJrWtm52JrtRQSIk5UVS8pV0rq8122bo95ulCpA5rAjEP6G9THm8xW2pI
+FVkQElkd6kFx/slhnxnnzXqRQkVsGPHvFSPX9CFdqIz9TWxBJX+nqJRUNcib5vrf2XRJe77ytWW
nW09E9kPAqEwoSrztIUZ/kY4B7x9W5lh2EvIAX2fEGv3LC+71pD13OSVRieXHgGGXZNSRmd3kOLH
vnn0VHRPQlznPfaLmuAW0ASGZIF3dzzaktuPDu1KqNwGzz7O6YV3psExAIDrGbpz49Eb8vYMAhXw
KGI0XAtKuaFh0Om7A2a2BLuZ255pROsNUOlhGsCVErAsn643PNZ/2eEnL0Gk1jgvpEgjkwvI0Uuz
Gq6rducBhHhsx54ouiGz5O3RW6ZcpxHiVEl4mo41aR0py1rUkmuXTi5R/rC973/yznDlINYXHIsg
nG4mgaEcExzlwXooIo+weGvh/s7/fOwG/x3q/QYSPKMNUkGgIuud7D2HkXd2j46+9h+CIobwDXjq
D+xoHC97dLDQk4YDurk1MB6zmOKeKhglray0Rk8R6CkwQlthp4C4nLHUXociN2NIcROKvGPjKZdN
iBxn8j8Q9nnXwc1kzUuhKgQqEwu3pVP21ESoS0YdEa2/T3PcPZcoqDlBNS78Vv9Pq/si+WDr+c4N
eSLUHnGaXp0CttQngm+c0QMJpPhU1suV39PRTRWF/IcIK3sDK5t7JMKNvFW5YNdIf9K6scK3iX5j
EYqCleTRCLXfIoVg9SvRLTvpnjJjuCsH4pa+pXSJx9fFAPD4K8Ctv+n2qu37z/SEgpr1V00HO5a8
nd4KWcFOiv/ad8ksg1cdsX17h9B0I14uHaZWRGAvCELVskgcCOylnnHDninvu+hVEU29nZo7AY3N
HkbMJJxMAE+j/1X6bxI77KOgDR7XA6AlLwZPFiLRaCEH+JduT2x8sTu/7iibeoPYm32P8o5SM61a
BltSPoejgkkPOREyFm1d+65jl9KtoOq78wMdfIzVTrgiZ8scJkduVvo7Ndyx98FbQM3775/W4SFA
FySVQWnCusFO9jAuy9/XO7vKhPDPwDXjBWsNlPtNZhiDPE8txcIN3mXvR6pa/g6GQQilUoZOzeFF
4toUGy8MTQlENW/5bcO/obgEqTl1N7qwOazGpbRf4aEVQ7Q+ZkFYidN9a2GqjZz41UkB/VnXMj+M
iQ4YQv01bZNBm8MiZP8U+CdIfBpnlQV0R8GKvZhGzm6fZE8mb8v8o8yuca1Jk716lve2SUyUhZsc
QTNGAhLQ6ewJ4Ju0tGyCqYBb9vhgT3zEQP18mUeLSDMZywJwY9efjniVwrg6KznYtpnLQhe4zLxB
qIK+wxf/vyF/NlSuqNDu82x0paR/ZOLKNjuZcCn1yRkhC9i0y8MlKxDm/okKtMZlDBNmaPvrCaW2
TXOFH7Wbsfi4ekWxlLgzWLt5gJM+Y/mtuwS8j9cKOVTLu34pV72CGleuoO8Lf1E6w2gkvIf4C7Hy
6NqIHcciVYj4mosTdtGj24NSXoiLijhX5010AxtMAkZDPOXKkItPEUPgz35XIr9OhuvcFochYVKF
gXCesa7YyvD+kIUw/N5r8yyZzdtalA91pbMgLPUWO11YTs2lCyKksgXGUUgrSAv4Y4O5/8BgHTxy
Ihy7bQ5L9Y/e7CIcDFa62FSM2NIsBOS9Qi9ktmQ4G0u5igj4oF3361bRoFt4u9eEMtYAuBaYwYXw
rVdEQXF7ayJNf6RvR+MsGKkKlX4pjLg7aQCixFP2wK/zODBX6zeurFgt4O1l/wHNKuv/xx5dSSL3
24IQ0EaptfDg3jV2njnVWaPCi7dZcZLgNNWlGnwuAghO/qiHyG29b0F3IOPnYl5AFOeA2oDrSaD3
YV3asiY+B9jrDPZbTn/OY6g1FgEwv+Aj6/SJJXoRXF6USeM2k2POSloZ6J+/kZB26WvVHYU0SZzm
0WO4LzYCQELvJZTp+UutwO3WIZfnptyIe/Tp/KpOE9iJHEKDlszRB8YC09u/pbfZFXOjTNJUjXwl
9VVtWtBdUD+fS5aHWJTOyu5nKWXyhUEvLr6aXEaFG3o07SevfAMD6ovhHS9jp6N6jjAFK6Lw1UOu
JGieRa72ua+4sIwaToaYuGbT0DWL93GmZgkPCLE26mo0Ss7GlVJLWEFNZmGuPt6OYaJgh7gCVVyq
IVvxQK4mP5nWRsA1W5Y3BeFxoSlxuwwcnk0UaeODXAfmBezueQ8FJfy7kgaBPhvTzjfw86ccap76
5VfMmxWResGNUpb6Sqz4S6CL+1m2cj3D6CfQmiU/aFMRuXp/ASEVgjLDhkNtI1fqTVHMtUjE5WSt
QZZZOchzk/880rUISHA4r22McIFUkkz/Ha26mu+anXKxSK+ikEVMLYuf1R43ZtDpbB0HDWrb+Prs
rYjYVDpT4ITMYHwS5fksc4nZb09slPVHwqqqny3ZCvLDI9OB5xyXIqANvJt73Qkk48pTg6GtRgje
m34hcG8hDmMGJ89WF1iK4TAkCxqqVm2fFaI3ed8OxTALLBuhKW7n/6dTkxOgQaDzWiR9N0sbnkNh
IslYGio7jNgVOqC3yfms1JUInQ8msEcla8+CyH8+ht3VOBKWvltN3GmzOVAx/T9VdTwFgq7Pd1WI
B07GQo1WmK3gbAOb7rVzlcaWg9Aj3b2fM085hFcKnpwJD81etOdW3H2QxZ3OC2Ku3ieeiVs8Kfg/
WquNL9ai7FRBfwAc9pTq25VmmK9YgvPQpwhawAxkWRx/+DykbvraF2HeucLkjVUa+yZ+cUPZxc2I
FD92SvUj6qu5gYAITHOAnjLd/5Qs7kJg8BC8IffScSoJL1n/VGD2ZqQUFYamHnN5xALqBsAP2+23
4xAdadHLdYVRzhXOabVoTHonkCzYiOjV+iJbKQZx6VL9alux2CS6cCrIoXxPs16F6zM3d6QPeouE
g8mlWU03QPA2vNq5zXjs0c1h2UfdxeMYhDI0d6LDKZorFzb9CBzAZeGsiD/d7mQoJEgVS5LOmYFf
+4yFuUgmkd3AI3y72/ax/bGiXSi3gKl7WRXm1/6q0NmYoklGL4sBDLDReGu0COHgPXOu27iRjlXO
GDgBEbDlVcI9T2AjbvP8+o6RN3ypprCm4YbwRWuVmIhzox1oOxEIAYKtoDZsCCQH8AOt5WZdk0yc
81zD0nnVU9zyE56ZjDIegyOHk/ERWRR888uKkWPIOAUkLtne7BrbaPh21+uLGkh7ycDeyh1QBbid
K6R7rrndoyI7M5sGZnLmPyKnDBeFjOgoTsH2jweOgPJdF+HYRBwaR5hk1h3F7aOpubYacdLH4GCm
e6jWJFPugfNciT9itphJ1c4VdHVRSmP7wFrqszvN/gGUIKLzIOayOSXg4N77utL7BtFvgpHA8S84
4TtqhYXhz/dJfY5uTYLG+SYKGMZN9WNrBS7mqeD6+7vwoSnC1qpgm4TIAkZygYerAeQjS0Dv8RZJ
LsJiO9Za4VEsgMNBik/ANscPr8FtUYg8vyHak7TksswJck7tjrZcjiVr75K2nNdx6ykqQKXHx4f1
6/5ycoh3BYa9XsyLaMWbkRQepnjJCnWQt9ZIdPjVd89OV9PSJHVivaCkBJ/4hQvyvCkfFaF6r4QW
OGbJGTjelGxaJDtKYbG41sd5r2zj5xYLidjneX3rqU8LH+Mpz2jk09CoXrf6cRs8m/VyfnBaYOdS
R+UOko/x9uJVikKrKbUlWV1/Q77Bf6QwoVJf5nzHSUVMvQyysUm8KE/T4KFnCdYn+mitA7mt6t6R
cIKcapoegEVAOmL/qB68Hqqd8QvDt2OF1T9LCPX2nmqGtIG1gInCEteogMTQaasKBwixrfZYidwZ
STxDTpnVjJf0O2MXA70yFZYYygZqkCpd7EDhu16B/Gai0ODh7/YUcZ9h6zSO2KB4OnTiG/usp+5F
grNtOe7j5QLGDNalRROZ76EjNb14o73iCx+sFFkBiNsjaexSccXN+cgvUf2sHgZYAJbbUwmzr8Lm
E/h4AYSqOLHPsKQXcTU0WzXkyPpIDY8ndfI+GncXo8XFH0+YKYK7GA/S9S9wil7OMGu3U74hAF1L
i8ZOtpe7y9lUo2CiQM2Ieu6Jugho+NCWsrkR/oBBQcLNZYEB8wMKe1BIAKoO7F1UeiUT5tCosDfE
q4CR2HJmUGDnz6vMdFmSSptJYyFwA4BywKIh5NJvSQSuVbbtRgQ8p7Q2m+FKOp+YpK2JgngV2oYT
sj2LMr1BtIWK/g89lZRhO/ZSB0481k6onhblpRyyBQAYhS0iso33zW6DNYnH5I13jRrRnFwFjGVJ
PFXg+21jWn2yOqfK6My8xSEZ4IuemKd8sH1H4kdM4Rj0o/cUwhSSh/t8tQQHfh3OlVF7wFsJJoPx
uqztrF10Hb44BrIIun4/iGQFSYPf7ZB9hfZOOH0zwNHQ7TTcQbubUtsauvpg1F0LW+U24Nm8lGW8
6XNl6t4gE5kldHWWKt7XihXGt9G/kFcyJDg0EzOmzzC+qUfm9fFB7fajzoWkV441NpARIZCimEqW
U1wQ4+WMA9X8houyRdKF6Yhli3Me9Vp8ywmBadfhIVFGOciaGWMnzmGMWu2iMMgQAVKxHCewAl6N
K/BbXi4ewxk8UfiQJBryyTBtO7wmrYpl8fD/mMqB4bYI3IbVp9+ZaTArGJ/hE/Ivhkpk8GCMIAc/
QMxYTh1yzQkuBqQFa435W0gV/AgR8QKerrl5khkMevRqS5Tb4a6MK1uT9Xt6iKb22VNiW6aMoOco
3WCWSDbCQrGbL24qhgsKcZ8ZnEDCd+qf3l0gf7yAVaryu5CsFkRe9esGGdOgf/O+88ioHyIs9PvG
LMW2eCtgJZUgMryioZDM5yRnjRKNjkvjt+897qK8IhhOYth0k/5PHZDy+MjOsqHcAH0+LiwxRHmS
oYgByBINX6o1VxgBhGPa1WYGLQLWSsacbcjuloZZixmD9E7PkTjxpo869GTiX2XXKkURABssWdkU
6OOw9wS3jf/oa+86i2xo3D9Z+m/pIpaonhdKBYOYRqtkWUwf+amJLeub+H76b7M6yifpgYXIYARk
D5WrDC/IeCgpf2ucCqRHr9tD9ujSvF0CU0VmFMkTZuNwYmBeoUkwAiQUR4Bzww8B0bMDUhjRvxnf
jHdKsUTjSNV8XJU5W6y0o6k/R1DRVTIfOuwpWNhM9c9UeRal/7tsNRUwBKLamTf6QL5H3o1sEsFF
e3BKS7ZtSm4zfMp9KAqon/1m1FiaFx2ptdD5BGZ1IV7wJRk1DeIVZwug9lnrrHFJMw5eoyjRcrex
qtenq5ihl1S0FqcUFYqWI7+5ssOXc41EOmf+Dzu7ZwUNTqRf9Q0htDxBy8Pj0/7zmQbkXjtHK8Gq
xZqJgvjWlQBpbykHIJnldhS79hwaNwIdN6NrFoLFwuRPVt0F1aSBXHmFtMDIQIz7+yZO1/Fn1HtL
u7DwXDmEphNzRKWzAl/KXAekQlRT6Y/pX5LfblFgAqi0dwmEgaOcas2PwTgaieC1URwJ1ai82e4b
tRuNHEQ94rDGSf3SBTDE2WctYJJ6O3C1d4r71kXwJ4nMFmiVpBW9Txrpmueeixw/nTd4tLijJJDC
8rEozW/EzAPDl2tf+0tYn34SBq4/c6t5fL9UtxN+idVPNA97AZDFVk8JjfaQWDjrlbGWLX9AoLL3
+ZAv/r4xDh8kosJapV9JqwTQZh7BFx5CUBi1jC1jJ63zjB/TOl5KA9EFaJgCfcExGFo4h3wK3Fwx
7q036zECElL0JLbYJiNHOFdzbu+qJlFis+xvI096BQ28pvXS0u+g4XnxfHEtTlIcEDU4dkaRH/Xj
1quZantAmIhK46B25jp2QkTCfM1UhvGSCJI8fQpEomVKpXU3U5LtOVHcKVLEpvkfzJlCPF6VKTms
Mdg7QVdXr0l4CkWx3//ZbtNKaEvjZ1vpYfJzOMsyY4gsTj5Gd7ABOLUUCIF07/oyIYCSi41VQarT
cFFPa5bHFDUO7DBG5M4/+8uhE+uiCkvMGsK4zNMHeiFLm6QpFlQi5MI/I6S/FUvgi+F2F7IfhhpG
OE7yUvudzGWRlXyFSZxR0FSiDV1bf4ijZkPe/i0T8n8mJas5xJZk8DystIRvy0S7U370Zqvjc2Jp
T8FpXfZHzEet+Pmupf6gO0jFJrBkhp4shqGHXPpBMJXIYxsxUEzUH47gWW5OEGFTumlM/TO0osJP
t5pbuoAYcBzzz17Y2jC9TUcGw6tQ7Rkxziea6cMCNsgiTrdrsPQyoDX21nPCcz4SymVauqfcRjaG
xyr5g2Dml+pfb7gDcknPStre0JuzdwbLU9GMUQ/VNICqcK/Mu8C4vt8udo0eHDhrwnfS4yoB/zNd
0oOGW4VygSwJkOJ2l/5uKTRhrHqJJ8eXgqvkTIOlvP82CeyEjOrKtU68H3Nu2CPhhslvHJNu6MMT
Q6YpRRZjML7nWSfvmSakM51vKLJuoZHdp6kKTQ3qyJMlB2a8KTCacaBCJ7N6TlB8ip/eH87PsNO4
sP2/F1JW6iR2dFJcLkf8Qpz6obh2DMVusB1Pcvc5imGggP44Od9IarwK12+4HPf6WcPgDTcCUYRk
PDcYH8ikXjXQbMX4YXoRtU5zgovB8fO3XPK/eqhg3SsJ/3yRMwaKsog1rAiVdoaKfBHLWFD7bvdC
2LFbIS9NuwOUTWw8hW35aF33+gGU7Y8tJkD91UDqJPWL4uJVSn/AC7dF3/i5VwcO4/gGMs9GTpMY
9JMc1YGoCwB7zUp2eHNpAC0bDCip5x/pvdCPv3xNuiEiE3E+AWJHSlGE+qLtaYCt2a25JUFx2If6
QsbJFZw695BiJh5PyQkUxTyZznP8aBP4IqcwVX8tZQoXuy/nnYH77+FyeL0FiLVTsjrWbDJ+MNdv
8tCaq+GCfbRscKXcEjadSnOBZZwxtiYgcwHmxbliF9svkVyK8xb7PfYAV2kbMToA3sHejKR7ERld
bHMkvqp2pToj3YT+j15wvGN+LmC2cjs5lWpiS0kkOcV2OwaKHewxCqMMpVRGf7h+CGYOJGXLcix7
uE5oXfcxREvb+fLLCQwBFvGbN/QPKnyJ+LUCiYzsCL0kI8rmtzeHjrfC+wNewDvcn2dq+a+GgSCR
ou5imu9qsn2RbnzEf+jR0T9VgaQl+AI6SyfUrdQo3gGt8jVUTV5v+NJ6WjO2QyjhT5zkR3nZsR2p
A9YkcCou43SgYG49a1o9IjIU9nKjRMaaa0qhyvg36Njkjxpz5p/a6Ylfl5cprDRiS+ZnzHSF6DNg
zhfj2JDMYHTRdGXPxYysLednixcqTsmrKk+Nki7EhSBvtneNzS6O0Go+iWilh0l8+IrCuwhdIAES
zvVO4fE8s+MFD/q4GtyaGYXuBLK/MlgY0DT+768vy7TbG2RiCM9oE+oYl5hC/k99ngrLSD0f9fmI
swykl2iFoS+idYbXH7fOUw0AgzULiD8mJZ/fNEle+Qq4wB5WG7E7WNHl39biYGvmNHkuGGPAvdrl
KKHJkYymfKpmWYjvOdU/htqZvtEGymtgII3E3JWKWrmSpjbrxcLWLmZ3omNf0ydcBymWSf8OsTfH
G/2J4nVdUWfPqKz0xDQVZOSeUXYUMxJl07oKE1gWwl2zVw+g5Y+KIx+JZQKJCmsb1LgPTa4Xhrde
Yki0V9wUAIBsBRlv8Hve+dfk2b6WRo26Z5sr2NQxZ8NLXvjyMvQffZr7K38El1eWURAbnY4tiJye
ApHyYfoahMDG6Xs6kZdxFAMbPrnlztx6EkBVG4FslDqPf56Co5e2BvSWh+abyBxUTY5DuxvzCR6d
lZf2db6nMMYlp8Io+217tbWFi9kapdTX0KSdtmng8LqyQ9kDlUg7ja/wo3IxENfsoiLvqwz8+bxE
IyuE6DkVs8rR2/VJOg4nMTWGqRJwuRWjYVz/XtSzzfQIS72/gjpd04KnHxSmmRVP6hmR2mV9ISsm
GIZr9oaLrog+bzn4iYZS89LO/aPu+Pe4Eqz/ZKo8bYIP9sh/dOeMmzeWfhwF0NaW5M1I3UIdcMRe
6cuxPE3xug+sIhdMO0uIjZdGOi02z9JFH46kR59LIeSQ+pK5/W6V2S+NzyAsk9o3+wwWlLm5bBY7
lFEups59aUoOMTobFZQ7lC0HMvfbFnCGKpZBlpCQxxnFQpRml1FzMpUJHNrcNQbmNYWVe1RqVL4N
NZm9X5cajH/rMDUxy6JhviAT8jYd1mg3ho6z5uZJaOy8oKwXtOfA1mf3Uny5YZAQ3gUuvJBIQxIu
QfpjfQPXfswmo4fI2IdVtGU8A8EtJQlLdlSCfOoPnybyu9Z1ue+mWIwTQ5x5BvGv9xCZQt2o75IU
SMb4z9kuk4wcj7AF+vIrBWZ1O2JSkRbfXnNH/IIRY1AGQIlN0wEU5x/o9js2YA7f4MUXqJdFwqcD
lESi0zADFrC3tdL2dhfwLA+jVNoVPiOZfGM1mRJr2gnh8VEeFn4Q0mVmNKXSGnLQ4GAUczmOL4aN
H1qAYcIf/YD8Glgq/eSGwmP7XycaLWhxgE2mCVTBAD/Ol3ccYoJCA8/otm53huk5e0lWP4G+Bt0v
p9gvjeFMyYKgDjwTWcb7nVzumuhTP8aFf2WNt8q6LXOFyJCkP6D1EIsF3XssKKJS2b6Nts4UHZVg
XDmILv21tp+iTu5NeRlSJRgGyRYuLuTu4iYw8o02M633IowGSwJ4kccDW5TT3MgUb8UE9nro/ngj
Uea/jHmbXArot6ywbjmvw0uHhkmXZDTjfJvRsaeK6P5Ek8eRRA1TdffpSsQfBXYnkLNcpNKrJkgU
oQJBrEjESdJJOVZ94gbQu3I5k6qTr1wVcAcaohCtrzrXvgxqHefQk+jZjNb2y+jXLMbcjDnrp852
jdNnZa54uBzfSBWVgysenbFSEAwdUL1Ye4VQSRs7lyrIb0AdEpdG7fv+ZNRvY8OVbO42pf1MKl/G
8GObuVpIFaw9F72Yr7BBLtUldhoRrK2aFthuN9FO2f96njhXJ9vIdeiz+ULgGDdLqhtJW5f2Nt4E
bMh8a2o+Hz1PmgCEhr9SWNzVN8WBDy7oANSpLGTymZxqe8Yk4/JZHXAZnRiSiUtJjWYtGpMVGgYi
eK+MZrw70Sf3xhD6HvcwSJQnEEBxH5y9ZWCWxDu0GEIqKb0/Ereut5hhhwjlyaMFBilTatM4K4vZ
WkuyMC0AYMnEa0rbT/g41CpkkllzgpuqE72UvdgRgzEJp/Znt6Jmn28HsdDZcbBhG/IxMiJcOOcA
sLfUHebtzr9YE7el8qT89hpbOlYXxS4Cu/H77LyrUynzAAFEeanoNUkBVboOes3HkcMIHBXVFOmL
DLj2oKzug+CCnX/tbMjcsVDeqLwTGkj1vUxW89tL/bo+zxMJWSUaj3moeBNxAK2p8y4QwFwVmrOQ
LCQ+t4Uyfsv/jAg9+bySXFyzo2w2uyORicSHc6gGr8sQLHZnNVCV0q2uxZa+33vRgsHs4es2TC87
5IQ1/Tdi8qwgvGldNfzVA4saRoL5+3EBDvnWzCXQzRLS3213ui4q2rQFxC9DCTkN4Xzrp0CrLcyH
2YqC
`protect end_protected

