

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MxpeY9fwU4EddFSpExWohS5o9i8UPinR6kQv/f7rVpVjW9v1XPHFNv5NQBBqnxbGk/3GroOhKYHi
zeZXd9sb8Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
genV68U/jEyVif/FXdfTRcDdNLXMaB4JkzDnEPHISJLebDAxHBqab4xQb3vzSMzS4EZxJxM3czS7
l6/Pa+/lUNH4iHFgH3/d34ImoXy9UrVsNWI4O1k56f8CO5JZkX0ENM2JUr2+jZNnrmepHCpz3pyr
N2xknPLUPWomWT5p45Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
4dyOi6X0ND7jxJKLfQYpMzBQUnXRUvqhIlWd2qdz2OgGY9VUivCAp2239OkMu2rIWSpkdV3gd8Tn
4E+XnpveIi4nHAn1AdqR2yW6qJRqYI/CpvcG8E7ZhuUiWSAPiQ/jcxRmeyzLFdVhgEV4hed5vk+9
Qi0C1DUHqDNPvc06f+xZUSTzBSqXkxyUqGIa+j3ZmCrjq04hmRDILUEkjqmR0K0TOLNdsLd81gAl
LqIfeuzK3hLcVWnnJG54RzS/q6bahPN8UaYhtJREcAC9BD1S+QEdDXRxFczj2T1LQBL5rSryR8bI
LV6YqNl+85SCCMZmZV8Io9S7fDVIrhzNm4Kcmw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PIdLn+S6alHzFt/ir7zZvMPdMeYQTL6BrWSuIGxsOazGugSdn7m2jtyII74LXXAGUQ0h11spxnUf
W/HpoHHxg6pfmAZclwmfvLsFiVi0w0hNMmIWoR8TGPdAC93Y5+aRfoAJNuDfUDfLzdBM4O7G2ZFx
YGYpvBcNhzcFFuSCCK4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KkGw0OOEdMUjhZKEmICwPPGTbEeQxk+K4HH0ah7Z5cm5dbbyDDJyn1CdBy6WY7ZD/SXDbXp0Ibi6
BH7Y9BzUsE3rhTUVWQo0OMHXc+hE0CnmrdIq6Yy3Wkf73IKl+pu+66Qo9W7SdJGNPpreGME4X4AM
zBwAv9xByRwGoY45EIIGTaE7VL15piKgLihjK8Y2Ee8q921qHsI62b9osdj+stH9M0nIgGIwpsIA
DiUOa8Naw0kRMS8QCXDqKr1fJ0jPj3cnclvP9Taz8J5tp8Sf8I6bs8irg+MGD1MgQIfeKkimA5VH
MerNz8gbn3+/Vz2X2+nKanM3LebAMLyCO8EBfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35024)
`protect data_block
gZ0sXTxogON2oz/RGbnBfekOUZ3fEmnCjtc0zWeJNSv7oBBwpy73Xuy39LPzEKLRNeYj5BDQaFtu
cjAVKzrwXqr1HqA8zfhpb6fLghTQ31CR0IvQao4D2kNgk8G+v1hGxM5S0zGdIKpu1O7UC6R72RL+
Db2tynOP3gqK6tiavsXeM93DsqrnZcCV1LOmKKh2d2MyqBjvQl2iURX7WqiHwEuu38t4y04yDV7j
ogum7cw2yqROSCyg+YVvRAMBVN+eeR3LWDPUXp5THD7X2stohf+uO7NNg6Xz2ZV+mb4+j4AvZd4F
aql/lpDHko9aRYg7bkNCAJ+pkqpS5M3s6KYzv+NobYvMtSSSEZMXYDLOKJ0DCNKcLJnRVPGIBDO2
hwx6t3JfGe8s7fRLjjOnIq0Rr04h4oqRJu9i/Ct226i/OeqowZDe/gQaV18Fgm5VZriWRXqDXHse
u59GnjBHaWDVaxJV1lEUZrgEQZjefdH9EPf1vncDTUjFoNEjlO/VBXOFcCm93fK89yaY1dWd/7Oy
zZY4MJajMGP8XtoBNy+AlKHH+CheNr1isUw2WbCRukH4jr2jmsxD7wKcaU7qvLtD47RYQE3I8zqL
7xzb3Jsq+BaiCeaf+93uKLc4ipake/OBzFvIlK8G/T2kwlziAJydJPZ75shWQL5+OShymbF/30gJ
aA9MWgs1CTpJKl+w5oaaKNTkQAIM32pEEerbjEum7CClDFcA1BjwZ3vXiSs0WGVbn59jT3EjqxjW
z62IOCF5DEMkvny27KFfC2uqW3dJevrgsdHF8t9RWrHU4w5Y20kW6FyiVZoaZDKNm+hWwsCrRPP1
dd9EgxY26ZOnFhqPnbdUmaIGk7PLl4/tYvYCzJ2HrhFpEjZ9GfD3A/BlxecSEsVwqbyj6Fo8bV4T
uxS7JJtE3TL46/LqCvgRXMVU6YEMYNRIQ7vSQBuAgQo7lnszpgpmcAIo3n12PJaqqrd5s16IHgRN
j9wvy4+FBXwuMqNtn+AhGlLsqm5z9i9spMdOhHVLgUXRo+n3DqSq67ysVAXIHoiVM7jOhxyJw9Hy
CjOCCRag4ktMc+Ywu6fIr8uVZQI4Ug8tbcFPe2tbL/42yZPvh7APzmV6Yo0dEbpOfKczOxGAidX0
C5ECkXpAczJEI0LN0aOb8rURmOEQXUPjS2VmnToZQQT9uHYd2aqMdGAFPOq8pH/iewlDpSsYErpP
cdmXe63OlJ4xIMYL9SHScEn8koUz3l52O40682Pr4h824YEFW/yRHCaJCmgx5W0Fp+GLSWPtErY4
HWFBz3xgAAMpimUkdN1BIIl2i1xfGDVwe+VEY9K+nddkFHEHjLVBhbotf+TRRCIYYHoQgn0/8LTS
6/cdIcWVtsM5DF3JGqmWY3pHjZxM8kxUw0vR5hE8+D28TkRM3EstfW9/8KkvgHgCwEDQj68BVf4z
sC155mOnFzzdfXwYJhDGQX9UxUrUphAz7GrPvLSjkndj4GUeBe3+o+gT1mgL5G8UguJyTCZlCmnt
fJobaFZqqr3enEIvpTy2N1b/0l79FVLupR2/Qn0UB+V3FPBYZFnrzogSFa6hq8h4HzzdimU2Edht
gnXzXVxhs87alBX1LvEiTGphiZfizG1YC4wNO6zVORAj+BaIwNZBfG0YJ+W5tySJe5P20M8K8/iu
JFvL8EnNZhsZN7KJ1bzXF7aaZLxZ8WvdFFuXm2ex415DjKerzfOrDRH+ix0T1yudeXojjOk1p3mw
NvjeAEHF1zdXhyfA03MdHlXJDTnWNW24sLlK1OM8h1Cn3RgWqy1DNXVgdWYQ3mjnayIDClTH/Ytu
RdBKwJY4/nMF63VcOmwvfVE0xIw5k4yDFQnJFfi07UDxG08adX6SWt5csPQ8YSFkRb3JjyW48YWq
KBFI1ANcMy9uvaEyIISOFfEEYxC744hVc9no6d1tZIhx9WR9hLhLFUfcdEG8nmpX0GPGpr/QzbJw
8kIfEda9S61z5xnMjFxFqcCmMKaqrrGx9XiQcW8ZAa8w90Ki+W1Z4caagleSarHW8RimRldlpBsh
J+qi5tiI/SK5m4/oAidssUK8vi2Ot24JNsJa8NvKQCjbpAtjMLRs70JAxH+wuSU0jqr1MNkQrbvd
gLxPlk5hiyX81aaoyuCN0tD8lD7F4DNn2uxJXDq2fKSI+m5nvARtITZOX+9F7VXRu94qm8tOj88s
kQB3oL0cH7V7JC8rhs2nO/uZe7Tdre4RY+WnW2syOK0cSwlBDawW2jVeWNA0x1+RXQHEO75BAOvo
AcGzXJzb78oCBi0EhoYbEKAdOlRNxWn54sx3PpvcYjVJoemLYw2EP9t4MqP0EGn0XnT8YawNIYpZ
bVjhJiEY0BaLhm/T6bB8ayfOCX4etuOq+VN7O13wYzsEimzsi6/mn3JfnzTTtB81je8jfoiZbZDJ
b9+/f8bMcWUOKJtjg2lnOem6pkh8zeFTnq6i2/g8oV9xg5fo/j6cxyc9lJSthc+gBQPEoSoil028
W4DzPk4HMOgBb1nWOFHHD8emJyA4LLhcfHGzSqAOvp7Iv8O/DbG6yqEP7t5p4lSyNlHhmD5k/Mzm
jtI17ooYoDvHWxEfgOiDX4P2lLZG7ZxQAtdCY1ZjFVHqI87WW8FklT4d1ZWfTqKQ2hgGZ29C8fCv
zM3E/u6JnZYM4GdSotMOcO5kVi0T9lTSpcpoUHa70GQ3bB8lU3m4c+EOnwikc5nY4C7S+ktiC/aF
wsNduAAWOpi481NtIi69DZZtd8kVWsuh8FGXOtJafTWSCRdjgeVdKu1JWqkstZ0DMfV2jxb9QA1c
pi11xpGL45dpGSS4z7vAnnK7Zb+oVmezqGdzYCtQ83UmCRkEmAMWVI8uW8tlBWjgycoit+6laZbT
Gb7j6MxnVcugTC6Ew+iTUhkt8ZgO+Cs/wiNel1jJ120HlCgvSJz/74gEHHEBxOtC6jesjrE9m1Y0
FQCcha1BDk8SwTrefl48/HYSCjQOjkgbP5fsDx+ft5wm4CC+OOkJSHAJ80uo2XVuRkzvoaX7kmgU
IhHTloXnSojVDap5GGPoK3QkuPln28ntaiZIyGsBfJ+LFjvhF0UzecZfj5OAcieJTSM4G5+LusmV
dI2v0qwCiZKFlb+YIpSyNcumWoBwLLRSSUrk2M9J/fhUIRdLOiqR9axLpw6cGNxrvl91evyGjT0j
DDCEh/AVtKhzqWZehUKZc/v7SQxvqBEAt9mfLCcJe1Pomd5KaAQhRgGGY/xE2YZ6rJ2/5kMUXUUI
x05GtxK7fiB64NYjX6LiMxm/K5XvViQ3HV2FsBkKzztdZFpJB1gACCRaR0P4zqHZ60Hfawst25Xv
VZkmjxXsZ26w0B3HbM1j+wWG2YbmIJaMRNOF0krY7EPNwur+BaR3w60rwln5xtWIKq5k6hRAGJEt
74S+cK7T4mzLXHqDSDgxI9BsZfoC6bWiBgfow4KoLN3QBnR9R+r/A6UphTXuDxXVeNRoAcUYysnc
zbOhxfXNZfTTTSJa7v07Q6VMEDakRlCxSCFh+cC0JFMJY1pJBWlT/oCmx65I2gfQu2dgC8RTGwUN
5mzxsLAs3hFv2oTE9TL0w2EuF80dPvA29VlYxkEYHpihv9UldvdQhWu9ySx+wrYEgHVA4Inbndg8
XGqUcQpQB5NkPA+/Xqt4IuyZXZnM0tzH5c/m7TupTTbFQOkZdrRjLEnRtSjq8KlnBrJnwlpbkU98
kxLCufw1NFJQa2Sj+cAjwiAc58dkcqkbFstn8K7KrxQYXVG0v6coJK75HrQDIX8kQ6m7SmwQ4yxT
j0MYNmEjh6T/HN7I5LVMof+MXZDgOnZoHUL7vhSA3lhtMBwJqctZenYLlhSLf+CaoGkizGdFVBXM
eF68CmT9ZrsYkLSiEl1WgLpMj5rPveQHvrnycWELFguKSAuaY+HNkAamxKoAQy/YruTABx9lpPj8
bVqqgmWlXo2JRG3fjwby39aEyRxV4jzZJQ6vArMb0udBQ5yNIUuZApwWoFsVt7daHYqCMQDF3ppK
dVbzvfGYeeBMYOc2sndjbq0QaUlyHsAF3ku2U80AVxC4J5TeDhukWRht7ZdOJiXvdxV55hynQTJT
ysW0yd8VIVdOdiyf3/pYa0Um76Zk27jqyc6s/KOdCoQmI9ePzORlt8tTcK45+HhuyN76BGsspFkY
+HEoDKVb9P81GtUpU5q2dShw7r1RPyuAjasFNxbrb80uAZOzqVmKgBanu24Z+r+AistkfbRI97+5
CjNPaEB6/+3IyPV3EbjCCftlDDX0aFzi4YyWj3USQbASGEfpgN9m7Mz3Xuenk6/K/ZMfSl2BwHOH
s2f9UpnYV3knWhGJoyBezwz4SuX1jymTzeB98ZWC6mieCSt5u/16UYsGF2xfrrqTttiAfJ6uA9CR
KbWVKerUlNubl207knfEhTO4+QV3Y3mUtwRbRfZgSVg5DRiymGn0wICl9UAtNsEM/WWYaLdD/mdM
Hlg8Kbx+x2XilsoKULXULxcx2Q5Aud7nZaPif7lhSNS9mUrlzsbR5I5Pl/hjx+igq+QJS5f79ngf
gCCMCGBpEgh+5A+GDaA1Xh9cJsqmOuURw0fJCjc/n7Z8h6h7jKzM9uGSONpjFBVB5/gCG2jLGKwf
MqW+PA7gljKgmWooGYjbnlMsc5IQE1mjW3vvRC+bDxg6lzUe+CfkhtmhUF1BdrQqEMAkHiOU0Bmt
o4A/RvS8sNwLAX+ijP0vWf/ZuKcebZaSWWpeKCZxJ2mUfCwaxC3FutR2XffbecBNQxgWpfBKn5WC
wjUixo2/dTQWWUYw36Pmlw2Oy6dNwZNYx6MEHZJW5TQ3AM45jdhUxJxI85neImI+R1ul7LYK8P85
24sfsfGo7l6NS+UniyaZxRHLNncrhOq/bPUFDbMOb8PjQYuUTpcr3p2MacW7lFEuy84aL1gOe5e9
kvlzgyQLOtCO81Pw8L3bQgq7hTce11sz6CrOpFnVU1NTlrE2g0buqcVNrxshk3n+69MrrUrdhOYd
rWi6DA0RRVN006MbOTJaTH3RPoRxTFs8nmS8hrsS+uYxksrBofHj+Z0Q+/o0GJoEnsRwMGXwAjqD
9jc06d/tgTeMC6pGq3TZhKBj2J6RCIRqMlsoD6eyJgBUju1XT2eJKBB4pBPnXhDya+F6Y/AbLUgR
c3ZYldWY835E6FcQwU1Sc4+ajyfCXjTQJS004WQtHS8NsYB6cqZzE3teAE1LLTpeN0H+6Yn2bqlA
R9H2AhT7gxMpAJeY/3B84J9dzKyP+RCj1KwiB7yYZcnPX3kDesLeB+S2Pb9X0BNNgpbPsE3wVI/t
pqUq5ZTTyd37sR1QVxwyQCf0vU23VeQuByK7BFFV0gA0apQLH9+n3aMQTOyIKh1low78qLJrWLVI
IajLxHmxKxevEwjfoYyLOnZkTRTqxH4O8txJAw13M41R0AsnndwA5axnb0Qd+SD/QU5kRczaT1lw
a7Wf1diZk1/WjOioQRkv1XUp3dCd2u4ht8+hq6r9/yaw56hRf0gfL/mQwHms8xNk5e/dmyW7wMj2
XOqqPDsz7FP8w9BSkjnuVk3LNzI2Kf7DmGUYSd9tpZ7V81DNp8msZKQuc8TXNyMnOs+BZWXhQ0SS
lGPG6ExEvMD+O4QZvgU0EJ79nnqvB9xqS34L9/0kVAiviQawiPNCM+935iu5Qx61BE6VwgNsj+nq
rGOcXZnEiZL2WcQbJC4Zt7vVfkSP85676g3SrgkE2UPEfym6sN8mVwfy5rzaF6NPsGAF2ak/hX+S
VGGGJQLQ7g5Lbc8WgkHO/YHDaIcizjxmmhfoLDqT8xMtueObIYcfQAbtvGAdZazPPF4QDwbgyOL0
wAvXipRnaABsYK32H3/5HMlFTj7CwEAmPaRpFgF0o1N+oq16FfUtnwRlYkpCcFCj3I1gZrdXNMcE
tb8jBE+7dFyw5Y+/8aZcF2hRWksirx6sYOd6vK8wXTJsBsCEEZJ2nQILaz1EIZ1YctyA9YDGuYUi
PATtISAbcq/yJG/1goK8FifaY8zC4yaNK9HNdmKaIhJdtUgxXo5MRK0u2Pl7IOxaaw8VEiaEiRaJ
dTW/LKeiwRlUP38zAf4K0xnO9MKW9h91v3gPys938z54jua0bo33EVzkwrBOEESB+c9a3mdFZIAl
BecrlyNEIpWe8NOFUQxxhIBRqp1jJRvH33M/YxIs/qBawwouE+3myA7rvsm87unjBQprBVy7tdre
Si8RY9dVKqkGaB/8ock2mLQAKonKxmy3+oYPUCnlqQcHzV3tbYfM8Z84fSctdmiHwQxxBF/dUJ44
wZviCJnNYZPwTiwz8Lpto5MsaXQE0415uxjrUQmlMRNrdmfLwzcStyie21a/eymldvYa7mnyQIeq
59Aszv3WdyKNBOsWqJiTV3rEVkcMVMTQkC0FE05yIyNdK9VLRF0ZgWqlMZFRbfJLDucqYdsngze/
mL458ycsMh+2jYOZ9I7TMWVK/VICrJ+n7/BGpR2jJ/2YJBSEyqxOSrRTRZQK6w4PuyYHDEL87ce7
nIVwCwo+q3l4g/yi++bfqwohbgSF3g7Qe964sMo1a4FzHvA6ZaNTrvzobGvrUhj2IuFjbla8nwD6
xBOBuE1cUdLbvhuFOvp8YETfp87T2Eh0qiGe0LZsvmMl1KVZXUCvFSr5DbNvefc54af9irskMe7e
+rk2Ep3yiFo9VUWwiRqI1+Kj346+cTDrFdVnHCoeJqjVEN5/LbZQKFZC9c3kLVSWxh5I8788LLZW
zK76p1gIogJfTqq5PBlu75Y1/rXJYHYZxOPk2fEKLghCrqkLmxmDXKgacr8Ov41rDwOd3+sNA0B/
0vUgVarf1aiZU6kNjDmDW8beRISNaRbfja8QCOmg4v5hV22ZwB7jaJJdwR4HU52da2JayOF83/ig
nEFpinG8xCqXsnRxWoknVYaaTT6udD/FdFCPblZZOseDCV9kQvRmnEOavbsxRFhdD+BJcCKmDosc
LLMjOxgZLk64riKegHHw2/jTsDYPd8zpKvSoV9busqs8GzzNMjtlByNOZpI1ZNdLrkyNatAJBOd3
tapTbRrT0ZqmZKzdEm1SJSU0+MqfxN+8bRDxwOQHleTCCz6AsLkuXz//P96AkEJ1VQY3bTsq16BJ
JsRYZ5tG+cgibb2wnQO8MMIcHZzuV8R2HBf1d+zZlbdNoRBedphwewOAzg3q24TrhV070LWj9f+k
6V7lH9anrLUfB+MMN9coCoQaNfFKXeG5CMW3dfwhJrw3MpoA0MK952dBDfAB8jQzpEy9oUAnK0mJ
Oc+jLf9HTIFXhGHv/xA5S/tknMBiP1FySaFM3JEH84SFS/mcD0DpkbtEJgipzxOXhv0fD/KQJap9
Nf2QYv2egD5Za3ItKbCZwC+FnyDpbm6pTG8v1oNXli+7W/Yjno3buhkj2JkGTB9fdq/XI0n7uq4M
4ommTOm/s9S/e6zYntRUfHaT3PFBF3JN6oA8F+h7hNmOP8u73xzKeWhsnrYOMkw4Pv0HXS+rImdN
ZJf6TpYahgxdmarakHqzvj1cymmV1JQblKe9rZ2LvhRr/8jFWE2eZYinYV/8pEFXizKQXrNK/JvM
15TOLQaN7bNj5mLXbIFrsDEF6TcFKEhZyZI/mydjp/tYlPtq2HYfNymGvfg+uUgqivf7+ctEinjs
IVKxrWxxEKbrfhbPvA0H2Q/OOmf/nWlRSDS53zqTugt5C618ZM9O9eBBt9NyHBX2KQj9ptf1ImRf
UEn+qOxUTqGnaU06gGnWJr9FhSN99h6LUiH2wMwCONARCg6VgE4SLwrszhNBkUCJO4dvXe01kVzT
N41LLzO0Avr+1WPd07aUXA/TLGueetrDZLwrgeoKLGADBoZu8UVadf5jhkLX5Q207U+a9Z2AYcPM
lNqSCKH6OIvnWuBHtsh9YavR45xI0Vsu7wxOCvFKuusw3HQEiHVN6XH36PvXys47VjSqElFYceeg
BPizU+7JwBpLxiqzt5lM0gm/HdEFU857TH6KGCZ1Cdu31lumLbFEEOLPCGJI3oHL1q7YXyqa2TwX
YRQO8YtEdFouZ1E4vTyxuDGym5Sbno6oxfF9FQmhKLqQhC+SyAipG6z9H+4mxfKQcUSfSzFgWdmc
TgitgcGJmRIUCodi+1+JmFnKrERNe68boPNL68sPczHWEQMKx7qHHHQJKwshQUX2tCgITcy4kwUe
UaYM35ta5atIpNLY/4eQAQHSlgDSOmqcCQFkPBHwxps8CJis2ZPdANFDIFldZ85o+iqF8K8uQQ7C
UJnyjM+vHn8XmVMBQWTrpJUCfYahJNiN3h16eE7HOArZuTRh2P768MEclAd2lCTJzYb7Pn+y19JF
O9PWzyFNIsda3I9NUkIUtVnLan+jA08eP1wozZ7FVy797fwvQa9aOxTzcjX9E6eQulXTQkPk0Z8z
fU3O8Vk23qvSaBLhYWfWHGnFgbKrT8bgrdMxu2LQZ4s0CA+B6vG/rMGLundO7iXFbO0kNkMGk80Y
xxl3Ox9T4tws/w53RC07dt6U8KKkxuBSYg4EfeNFyrrAt7tnpnwxwX9D2f4aiYPMrBNV6khmx8Rl
sM+82oulDMruKq/u9uRn30Ma9VmxrtUi1H6pvuDKxFYhK7B+Of920alq7yjBfGccCSjwbWNNE4iG
qfngijpzG4Ev7bfnf0zzaeWJhuZV5PzX5qHwI1rFBpE8U4ftY+JY/7OE+OCoFTO7UDdUpGUFGhfY
gw8XvbBAHYh0j6uVOPgu/5+fRCugqgpcgq9sO0pxPIp887ugiajGbNVApUp8MHf1AtMPUst8eZlA
Wq49vcNJjtPDvw8sTP619Sbvww/KE1+5FhRO/B6f++ggTTf0ec95VhqXcYrg5gW7oLza+VdXtpa4
TqZomAzQOJhZ/Dq6sM5TsJ8q+QzImHGrWgzoKhxKPVMyCjec3csEWCTr/bP1bPN4mAK9V9uQc/Rf
89ILZDE+DyszU40F0Fs/wxc5UE1x01dgNaN7AfKoRtl60nqu0AKGnk3/zEuOUnZEdxHhTpQp3A1p
bKtiPeCVd4y4mhsu37PKZ6E/oUQCLbv1ntNIVOL2S0gwEEUtp/+JUnCWdo3s/Qtz/5Er9i/GT0cS
05vCYSEJdXgricxvRps3iaEAGfH0ODO3qxvAa2YO6vNAu9AbT/qTqjWyb3jNUfRVbQazh2TW5uv2
JbIK2k+3XRJTe28xBebNJdlY+YXL07UChnqq10v+lEj+N9b2E7SgG0mgBQcGWbDapmz2/ApjPTrM
iMPBKAnUrD+e2yRs1kUwCMYfoClyzgWSDlJruxLM3OWauvQ57DEDleJd1ngCLXVj65Sitx8IhS8X
3tTYrx36N96MTkQSBO05FFA7OmRshonv8p/LQX/ZdHmLdvrm4Hrpm98gbFnjjpgmCeeSDS4CitJ+
1gH5cHVSgd0heMq57IcmecW/sccGEuVoFRPd+HRD6qvFFiJ1enp5vfORy0tshfTPQwmqC6zG7/bX
2HDkizM6XGkJB/qGUee5jRCoZ22gVNXAOA3UX0x8Y3t+p57Wv1WaXbSDGGXtDRIr5VU8NRyovKMM
vPdZq+fv5fPWXLAaoPH3sfG7ToSDc0QMJDzaEhMfj9EtwmW2FkCxpNyrfAkTjG1mnl5CcEatvOiw
Gc154dCB1eVp7rtnrK2drALVStZWAdxbMDLrBGt4Edcwln2YzVhERoNoHCC6H+LIPT3LsCN+aO47
QTi2BDhw4mGJOpnw2OBC3PU6/F31Xmgi7fPrG2RJMs69uj7ThocR7E0iomS573LRU07NU3g/tBSZ
2kg9xuQ0D/ZLXUMu/UCdmFZB3hpRjlRtIhM+Tp7d/pe/4VlMKkv+v0vTYPEwNPIN80Xf4zuuVTRw
bU/nA9W81y/u+IKg4UB0oFImQXCn229dJEEZbQK5HC6RW6Ci1K1QIv55L94K1HNCydc+XHj5qV/z
+cGTDexn9OPys6IlIV2SZT1wWZp2M0Q5UDv5+DHOkmEVcpX+dqmIAY4eISHHjlGsFyHuKJyu0SAQ
N8UYlYXOJ0KkNCRON4ooxR7K5oG80OsoWoilJv0/NHmncMjO1ezClGndzi/DOT5A1Pc+3v//DO8n
pKGpue3+k0TPPtBzKRHiR9zQgYmi5TQtK9S7sIOib8sv9sYtNOcTygpw5rbbFPk2TW/JuC6bSN8N
mvA4ZGR01dhU4ddGNHoAueA55DRXYxR01SlngNInwaEsCWPb78Pl70DQW3UsH0yzrPtHJaCQKPjU
y3feGkNVWbIjhYP9YP0VD+Ysb2ws6puU8hst/8EDXbFnlBJRsvnX62rmhqvAm2es6VxgmD4FxkbD
yu3TtPh4bAuceFTmOITXqaB9sxopVAGcfx5LMjl/vQM03aWRwQxcOnCPFtcZGyKEzsJblwCOoTRv
OhGsRs0dcjyo/p2Ok40kFZKZG9vqbdlAHECgh83YNcTbnVDXX6syD8zwGBUF0PMhS705HECmK/KT
3P42drurWlmnbSfyX9nPGjTqaAokTBeob6C1oLObTzaX9PtVccxJ3NBbRovjbw4DwWfe4Qzwb0cp
EtN1Z9J+ug7Wc4OPyzcCZRAl/IYPkGxsgGPFtA88veDIYAUfc1F0ykCzqsoSVA4VlNJYBoJ3h8ou
TtQ1F7CiPmg2yGWxqXTBqt+anrunDg7H+pzNN+Em4FzIN+9S3Wcv9Bj0125VppABRF10eGEek/1m
AaTe3zFXl5vMXkO/o10jWWjhQFW3FxrM3h6ZU+N+s4+zyrHt1y4wFmVN7jxVjA7ERVKEUZi90GSi
wZ9W23HfBROcSWgsfTDmwf6d0fEnsYr7c9awmOAAyIt0025lFlXK6rzwVepkiAWGaNo7zNgPEcGa
tGCG6ipL2fIWJ5MVRlFH/yN7I91u1kVQ3eRAGOnt0Q5VcTJLTcnfOoXhEk+a/bk0Ef78D0qdiVOo
NCMKy975lw2nUimO2c9eMkALUlWe/lhnaFUkx9n8+JnYPZUdYvL2DYZBbKOWJjSfXEn5leDJfdat
pZnhJsXUFQfoDbTuxeOza9GyEeoLz7Jy5hwglh8aPMIe63E0Gb6xNbCdN2qZi+ohipopUrxgSmEM
XHN8t3hlZU4AyyVdfips1HEQcsWxEgdorceCcI8rxk9zSndA/OeEVdsu6mjTIQ2Brhc+xeDynGWg
2os3oy/j5a5GkjnO3AyVkA3qkUt3IL8JtDhC6KpuhHjKI94mCCkSzYGJudz0FRMnSXwFII7cSEqF
mwZfoHCgtNUlhWh9FqOwRxTEGvRR2gd5pbq55iFJO2JJAUWjfAOESgCQFLmzDd5TtlG4yS0AWxRz
eHjH9ZrHTSmZdywkluBYvgTAfk63FaEo6qCxHsri+vjezUjTPodOz9eUozNHG6lNyBWP6eKA2ObF
Vc0Uz1/e2+Gt0UMkZZ0QkIoucDbaHvlIoFUMA234N0RwXg40RY5gp/rxYKPpuqtTjO89WiY1q919
Ii1gvf7/emQ9HkJekFJkUIhkO3QOvTLHZ8XwkGPSngFgDx8sgKZxqVD0G1rdWLhJQRJ/0SWE3CQk
dJkf2urd69kt0vPu7b9MgDl2Ema495DTc802ewv4y5Kz3L/aj8qZKshoeHph3s7GWSAKnES/zOUz
4PUHtDCIyOnfwNp6rT9/8TfCQ9nliY9AAA7tIDIMn+ghcmdczwOjI+0NqVr8ZMf2H46+nzFdYJYg
00dSUYkh9UQuOyQFh86PCh9x2WLxJyGx2lUpb+ec1PSr+F4T9uJpqAz1lixU8i5iGLftgXglZ0ts
epUX+TtqaoJ/MmUqI8bDhK6gESCI5hIyQk1b6Ci11SxEkQQnDdTnGFEthFe2Zm7vHo0P74euqIvY
0r2ifqHnXHyBXjL1OEAadPlzLycDFYbu6T6P6C5zNF/Tod6Ee71Vrg52cBuufRfvm5JGEhZjuXHs
nio9aH87DKBmd1AAvTHbvlcigJfMvvIsuT2L6WvzV3R5YLjSXQsinDWSLV8H7TVQWVb1wQN4LZXC
nbjQmSUm/48hUD8dyiD4m2TRz6zWpO3EvQfo+lnB6VTXx1zWQwiEPL36n9kHsvG2XnpthdD4VWgS
J//gCa+TO1eHY2G7+yPoHdi3Qpp4vNMMf8t3ZzoQl9MbarVxJdZFOKq+kJEvSwYif9R2DQUz6ovt
duF9LV3YxCBWyXgtBUwbv82FnGjpj8+sh0tIs4vVIhbMtHz7xc3UKH3raaYhn3xWyo6yIX0Mscfb
qF+v+FNgKrwm+4f7jqGPYPpkQ14O+v5xWXsw4rNTrRcG7UtDlKZluIkWym3iUIYH7KvYWTvGUZsb
nqpqJlZ391C0vUpHgzxAmMP5k7irfMKO9gJs3pruWWuPqV91iyuazT8Dw4VkGM45Zd3NLDQWUdmK
Q3W3xRfvZYR9IzL7UyFAXotWo3Ie4Q59rZ2xkK59l8KhsUG7DsS0pgS1vxj6SGX7i3GMD4zY9FgE
FrIH5GZw/9g6Uv5p3egqXXVRGbBIKowJ8v7YREnyf9AO+XcKDV5jT7aG/f90QsCQktJQ4OClHOvL
fEJBg9TmIYCd4en4CW7pKL5YcD0sMtNKd6CxKH4y80jGg7g0L2oak9QUxBswXtcdeJSoyEEvMs3t
8r/qmkcyYd7JMV+nQoDpf7sAPuymLeOfbAXcY8H7ZnPOT2hqv5rGyhW+c/5B//j1DhSxI/54KDA9
9bQXi3LwJSIaFpe7rhAKnaSSEsxs28F3ZUJq2sBqwE5YiaLLttv+TQk9qxHWuNgeNztHRzZ0qcNw
TceTsdanUufuxzLJY0M3U9yLZ6c3t1sNblXgzF0DzfKCNIt8WG2K0sa/9v+/J8BwotxYzGumOyE/
eEtskl8sESj5tVU74Lr15O2+UAT4Ym6zadaHPXdt/M4rVQwpYPqSiMJrd5N1+dPKszPP0kzbNTGu
kENMKXE7jn0ebJ2Y+sUY89QfjkPIFMr1luUka92CuhyDzehJApqymgmvVt85wLPne0xSFKL/GGtm
pIX0q8FypJi/7P8hgb2POQwh9oRR0iNnOCyAlu2PFLJBNTq9ZMHNfJJKeqUofppUz4UxAzdbClmi
22QltmGioAHaDV8cno9aRa/ygctS7R68IxMGXxNOm865/1opZ8RzVtgh+a0qel3e8dX8ufxIjHe1
UhEkhujpJ3T9y9v8IVsf+6QGhTDsNik0QzHb3/yKIDyfNpp2sUBRMi06dp302KTRNXMfMr2ss1wn
5PzIgl5+gHDeneXog91kWPI2WcuaFCzpUSZjWg/hZTUZNT/JmPwZbC/iFDcCSN3Perw4v//54nc9
YtjS74usTJWKFC4EnsRtHykqDnF9k6kfgLcHivBw99rShtvCR6YIFFDq3zk2H9A7N840on7a2LVM
3wKCF24RvYvzj1RiBJzioSsKHK05AJNPt8pvaVb8qUGK4/bB3KVz/6XdDvaFKkVSgmtSqtTQ2aWW
4/On66gglNw0484cv9qNWJnmCs9Cg9nWkJ+gP+RGSmXrEoKXAe0yVt4l1n6KSVztuvr8WJCIVPu8
hHxbK7NOmOrmQ/asVU0IQekCWQ9P8M/ViuLkLUOfBIvFEoR8zLfx+InrOfzvEgKiNHMNjgRkJ+oa
dOUO2tqof0EwfBjPf4/GW/7suj0MwvS11H9z1CGOQM/O/Yivy89xbwPyw/NPLZu/CcMT2P3yIx+F
nsV0WFF3U17A4DOkAvGPvbPDH+MjFn7gZnxgL+OLxBI8JJajgiI6LuJ3JhF5XyKrsDMEkl2MudKy
s11L08/2sQK/Ld1h3urnHzjLPRkYltAAiGy9THGKqwjmJ5RWWSyD90wmlSP0Fp/qm3C2SppMTmjY
ufk0J8edaK09IyeWfs4bu0Y//JoPwYdrQiVg16ksaeOZQOoWbSNZcuQM4S+yKN3Id08zI7wqywMG
18WZbi7iaHs1Hgyt21meohg2p8BH41fZ5iNM30/DEizPuItL1zQosS15J30WUbSw5bsctlEfHQAn
/9/BTbE+RuudGGPHIZ/k1q+k/X/cirHGP1htlJD9Xf96OyXcjFixPDtCP5SV/lOyeyuJ8yjuNA8E
2YvNUjPd43egw4CYohW9rVeOALOD7UERYDr963Q1RjPTc259MzwFlt3F/5ZnWhJJGvv3bLYCuuGV
TO6ZubcDeBINmYCX8seeRAcTojp+5pjS3HX/XZKpYWPz/Y6ywkqePHVCoq+xSiZf4EquZuiSrcU7
m6O3qtSKE415iGanyuqUYnGe5pRVJI0PKgPif4XVTnA6YaT3Rv6m3zhwwSw4rrQNygHfT4ocpzV6
IUf8YMhGHwJsjgSV+GkN3d/Tsf3ikXIBPJYLSd23OeqqlaZ8Q/X+hl4Vzp4xZ4bTHwojmN44tlKR
2wIadrJr2pzsfGyFO4zuJ3fiBCSeQ1mKc0SKXBU/1yekSQ3LLR45gBWR9mKcPH7N2flaO4JFdGJP
n4ix2pAlGEa+WVfff1AP+zg8LRwUPfBukAZvkqqYtDrKinyHWBJgLcbOb823PVnw1cZvoXnqKGoq
6tlO7RKdIsdwBTYLBYXOBIHDy8WTvts5KA99/L1GLEYDE896sZqz6VxD2VKI2yj/1rw2Gg+uBXAm
emMgHdjt/ki1fJNx/TxgQ1FjiZvfow8J1KnMIlUzmnlQau6WDi+fSKZ9Lm+1ud4nF9Ij2VstUK5r
aQ7XLI2Hcy8aru3GOyS7u4vWd2ZpGfJf4osBUvs/g7HWi1koszifinqQCFrk0N6kTGmwCJrj0aLD
lTQK9BTA7XCgHfs9Uy0H6u/UpogdEAKxjCxByAsEgvkVzZGFpegBLMxPvDg7zfRKv0WxsB0CBW+T
gje2Fc9jjjLAUX4IZye1mkv6tYecq9FHMZG0ruIDTZGoGh0+Q+vkDMY6GEBNXkL0bhFejrQQB3O3
lgzUzzEQSCVBABqW1a5y833VHa6iklEC1SGksRKiMxvt317JfmSZAsPwjTFcY3LDVzepkHZKHiy7
c+BVu1g6yOvxoOz4IDsUp762IxJCfF2fG2YQ/IbTd95Jebi2c4di67sGimw2AxFZN55JhLm3MSsf
kg872VWRhn81W0HecAPXaldb75GWsWFn9I3Jophm0rKv0PjZ5c0S1iDsPgIVduaqffgzGFAhiJOX
pspIOW+82leVx4lk7PJs/uE9ffYP2OJtnQ+InHJVxR//fV78SwV8zTQkDDEVBFeSR3wU8cngH5Op
ZOgN7XcwNNXIdlR7eXDKleMx4e5NOxCI4Klnqo9a07578DkIPcaBqwLojZSSEdL3ubpHCub83FnT
7x6JeUmq8yEHeCN1/RsixGyaQFBQGd/Q7FmCGofDuiIRH1r9ms3bAQCcFYxT5tGs7D4kfT+zPUQl
I4POJ5aY1F/MBs75/d5vPyO8iGlqEUlvWKGEWgA3WkJPRAcRoj2tqyAX/uUbgikqxhh3jhMsv/jJ
Io7Mvgnwua2hwqqTGd4dsrg8D0JqzAKh+WB4I8P3Ur2SatUBa2X18veIyvyHOtIGXsMfyIhb2X5n
hLfXHJm1ctRB2QPcDL+I5E0U56k3y5ktXpjmdsxD1RkV69PK44EU7E+BdYttOfulxyN+n8NmwXh9
xEB+7641ATYLvT1uGTwidaqwNhnm7J9ZvngNfURuRQvxjH66F0EqfgkQVsGECff+EjOiIp7r5Ky3
Ysg/YIL3g8mwJDBzpr8snSmDpvM4JCynWn5JQCVj04YrbNhpPFtxBBg2KiBkVkpH5EEhRZ+gNOCS
HutqScHggO3muTVmvuwC16KSVfNdj3tYRtqcYaMMzOeiMoEwZXh8KAWCTNviGSfdb6o+Os6/lRjM
naTwxf8ltbTlRUNTt4nyaIZSRqgq5S5wLnZ6Gz74npwMwkSLFkREZHUOZCE2cWZeSFZA+Pjf8lj6
7R8bRUbojFyq5+pT8ddD1ZGtcER4+DNb6iqwd9EgbRkCk4sC0G0bgTpCtinu7ZnxUrkQaLYpxiQb
ebXs7UYpZkRjnTgVvsaucdkRsvfsBc9JTxpd0WXDFdnrL29x/CDjfNyk/jD1QEolDQyMB5g3nDJZ
gTCgVqDCPYLIxwLqopmEUClniJsWiyHwFle/9npSmMEV9kizCAPcTzovCq++1YkDXApDabfVR+fx
vFAhQktNbcjPpHgJZ29llGm6cGHWBrT9QkTpkd06kIYQk51LavExsWyo//m3CVY/8gupDYzRozFL
4JFeSstRt4qMMlCtJGyycCIUFzGFC7evZ1RHqpHKNbxWlAPT2NaQlHIHcMpS94uiUw+vbKQVU2WS
UlztqgrDzMMi/nuY3o8nLRGwKhcxj22cuBm2Lf2ZWcVZwijUFwNN6mQ6amgemqPsya6WFJC90PaN
f8LKaCCsF53e/HwLEUnEEWjgxm5r2yN88XPm1u95UfCdZhBnQgxjkRvzWLPw+v5CAMX+zs0FYEJU
JrTWKHHDaNxd7SQKQdp2dsZENwMM6q03l4hZqCsRjVohcJNKNGXuJoO/rAL5Eu5LMztokXG+yzcF
aDr0QY+iJVWm2cG8DCTyoExink4suSyZReJSGw996JDNiC+fUGLix2xgSm8+IvTKCHH40P5phXBx
k53zJ3OGKEcmA1q5gajQ64SeAppHWKRHbra5Rqz5DaUEbCN6ane7KgBB1o9SgSD1GWGQasRAQPGO
64WniMvRYZjSqqiFVfNEwypV+RksoOPlx6D44uXY2qQxF5E6e7G2zRf/bvqu1dMenovZL0vHi/oo
/HFtdzRDQ0o4PlVOCp4q2tkZZPKmzJ39qdumOd+GBbTTE5NgwIhEL2QQbMbjxKwJEktWZIDr7X4q
akq4uPtgZ/f96aZTkV5qN8jc8qnQFehyMegQQO4PqqGW7gqeLbICgqXv+H2YoF9teCuzxLYs6NkB
vYJx6qQ1aZ12DafNs49pHtVaLVuKhNcTwmmwcZTLdLkmmI2KU1G5SwX6nOTj+j9LeDjaXVu8QrNY
zChOsvPI6mPodPGDFggVihWzip+H+UaAFBCm/AjZpwM0zAk5T8wqAyKS8sN8/8cPPscIHOMQ9Qb3
bVdJ4n3Mc+8s374flDcowE6IL1WKANlPucwimEQ3wFYJ2QjZvbCQf8K2dJnujBNVR7qmq37w41uo
x4lwaOt8TcrV+maJ0LppFFDMtV/cAw3Zhcznn0UjGKKPEs052tdPgy32hcgjXCivLG2sELEa0I/5
zLmrIIbqC0sml01/C/ZcOT6CIYzJOy5jCeNiLPe7HUmKcla0z2KieflcZXjPVcxK+xY+mhBQoeAS
64FP6BwSRT5MFLj9HzFht1Xbsd/s09JFOSC6tms9/HpQevBR9aIDqtKDBIXQS0MFHvIA+v6w283B
m24YBszEuxoQphmdzOyV/Z0GW0MgGlUMWx8B6TucA95LJHg4iK1nCfCtT3w+0Pn9mJzRaRiMhp7e
WpPsT2NtDuwRMrR6j94QzwUKhbkIi5C+eIIMEsbRWm5c+RQUx81KRn2HlJhgnB7DF1/OycajfM1W
1MbwLdgeIuHBiOMHvv2fHEcrz6C6oVK961EajzWfJHgkvGKIkKOPG0vQ8Q7sBtNI8zCufIydUbrd
S5qRqKniTxAVFPuvRG+w5azNXUa+cWcT0qYjqzxMhTlZ19NHlvhIef7hzyaEESc/NkxYZ+6oVkLn
hz94qQmObdssW7g/RYRLyzyQq+7ZRAw0ia6nxifU+VQ/wOuG2pWI3mJp0GuQgoRcd9UdlQXHeCDh
oiNEgipit6XkdY+eADmBX6cnVAIweWWNtlHNwaL7AFhYpFB5ayeLlBVSbkzV8K49Soz/iZoozsXd
nADRCunWGL9uhPLlCwO0aWRcku3SDgurONzsv2CrDmraF3ObtCaJyeU+KItgsqirJb5qaJs7ILFZ
RPoL/5C/oSuTWa4A7EjgYdbeI0/O5O4E6aYnG/S2HmXe9o+yuWIfQ6Vt4EVwzl2gahcQDQBxfZeQ
joTpWnISPEYS66LAXK28JRKb7g26AnDlQppcrntJk5PGhAkGVHFYsf6kFvBiAOiXpLv43uSFdNH1
xliTzeqdSIIXigUh/iMqH8KDbx70d9DC9wvs+6CfF1eY+0CP1xSUs108Mblzpw9BnZJT5kHWMPcZ
Dk2nqOllRnUy+3ClTMkIDqjRiU2NAke83R41sNfBKbwkf9f7TxoZcPhjHyd8fAziv7jUjAm+FH8I
F2cmbrRbjcSA/9H8ngmuprRtPpgzvLFgzNlkOKKgLk+BoyLmq2e+3Z+iBFVIU82LPsIvHf7/3kxs
UybeQPfuCFnMwrJs5Inap+N0uW4C8m06ZssyVNtBC+jYQLd9/Oyw5m7We+WvzSFXJ+qhvynfcqOn
ZO85WUoKicyGoWVXvgDXVSX40kuvQ4dBqK4nYMC7e5lnhZHAF9rmKE1t3G2TONgSKU8jZSwrA0PE
MXpdZQsB0x9CAgj/3SKhxp/AbPw0Yz3QHlG7F5LLHkCnUJ2PPz+YcuaDBBnpgV9g09JQy11Yc/GO
NNM5PUZvYpyZ4uhNxVmvfn38eTrQsVB5LmO7O5dRs4ONib13XBBA6/KinMWTzwIApZ34wbHeWaHL
lmpXNrAEUyjhO4PmrHiRKl6TW6dttXshYMQNWtHcp1psTvt12LCZpPHHEnIvFo5H/GNIRU+SKlXR
YkoB9xSWiKa2FpUAweS7WZ2HMDpLyyRpHUIYnjXbvtdNndcU3OicrWV0I/yO0t5gwHSwl4VcIVkK
aGbJy6H2ZEfM576KdYltSjiztafRV4RG0GQNSOaqYNn7shRw/53o8t7PkHttchWI1xdm0ysVryNy
G/n8ScHrJVszJPNRY1a8y0IrpKpE2OrmpC1mgzWpczWk/K9mA7t3gDUHpVVYmtm4gzK3aNovjL9J
K0cWZ7ctJ1132HdaOsykAaC5hGzYcLqP4hSK04sdIUCzU8n3zR3JR3GIzbanwG1Qvp7UqTEer7W+
PZNUTrAmW1pCyYeBbGf7Brzb890eLNBitS2qA7+PxwN2bM5lMy8ARRjKBhSnG/s6kei32cOvXtuK
E4k8hOeE/MjSMhOwGHD+tDcHQSevpLD23PDRsqCOgyLIeKTskRQSp0hWmXQF0bDqiRdkBzpRo2EI
tHuFV+BcMvjEABDLR1rwE26yB/x5Oa8W0Xqzy+urQt0ulI8fDQ53K1DgdahHAMdFpUXif5m75GkO
CbmLXt0GbLWnuVAO/IhQuUx6rhLg6TdZTGoTGS/5OQaH+mwLHH0xZozVTADqlk6lDs/Jtxlt2beK
xnk2sjaFDxL0+m4jxKKYziLFYrAgVON4s4Yo52v1RvgCyWEUYy22E2gIJwgZ+ilM+OKhWfsIfos/
EkFLQSnMA4rMF3wxJLhgp4Zfy+RkimtsBHowK10XYWorTUbtMstv37D4z/82HZwLYXDxPNUkWqDZ
XJxJe4y0QPF1wbOHUm5JRFiXvSjwHWUXYWAnz9PaANsGCG/yvF7WJkxV8/5iOU2uBJUo20SwAA3V
yJkh9xIw8CZfnNV1uEMaMwrnUTU+gXX+yk3lvLF+T5BOrzd2wfZiMrfSC5peT07Z6Yrvuvasyc7V
IKlsEEt8k8uVdvxW5LTPYpkG5BJ/rp7Cdkz90qTok7Q3lDWd1z59rAJVMCG9xBdZses8rdEboXl2
KF2rP7SjihU0WlT+3WjfQIh+6JoKNNngcZQ4PBFLtgBCJOYB7rcbV2b8saTUtiuYb3cCPZ/msVqB
FZisFIb7iWEWCSqt1B2gB1LCQcr4Cy1OKckC08HOnQD4Xfl7K3BqWpShbsLRJ3BCNsVlnhOZv78H
FbKRbK+6Dhe594lyfEQVGJ0kS4cdqBx3BEguoAkPYrLrbJ37n7MT0upYrclZU9jhn4inNK20S63Q
sgAjdLl4aVBVLtO/i9XJKJDDSdh9QREsKwWwyji+Q+fl9SOTqoD0bnNvSE2BQ4tf2lw9jhuXAYvL
bTWhiT+vlDJctjHslyIcwrDmv1ba4NoNw0J1MlUBhr42B7vToUlNWDUTOGaRLNfhCiaFlk1YgDkL
AHZlXhSCsUdJ/1xWeK9RD/Bcs9tXo1Ev7Uqepxk9t2u65eFE98TLhr4snkiUnhU7wuVkcsdvtl+s
eGF6Mnh0sOYnH3xeYvN2mIM1rl1wqE/Csyk6SpHUzIhrFxvdRgXND0pV9h/LHluw33eCuqlGfleg
0SIgbcohxHd8RCt2XOIwQ5A4pJ4b/e7Tp9OrJ2mf4PA2Ar1abaHaSymC76tZjP2N7qBV93+RbCqF
YUJRT0Kq6mOHJRWQgPGr+TSMt+7CILtAJ1iikDbuJ3Z23K873Bhs+UrzERgKsP6kBmk7XbFQzXQh
56Cbguez0DL5VxdyY9p7FfhTJHwNccAx2Jqf5EXcptrHWvP31991mfA5Cnr/MvF/EjUAobb7Y+72
1djVCqFT4yHZin6IEtRnfx+88/+IKZivgrlYKf1FBgGwXbkKMEayteD/JvTNWI14LRSgK7nw7Ezd
HQT/hfMcq8AvRZwApbSxyZJwAuddK9OdSNT295Zhg6KlwtpEp37u/y1uPwVzTeJRWwW8JFgMpks1
tBmYN+RHDCklZ65hahfjMhPIcrYoJ2DxAxzVbwBqPN+gXqNUVLIT9lCaaWztLu7DTlQbflqGUqcS
nEUHymb1Nd3P+6JM6e1DHLazwjx+p/eiYvQz6mz96x/lTl32JAJyJqEFgHenJqrhLybnvmPlsCuV
6Yf8L662OGVwzhAFVzM0T0xSDuzHe1TlhazUTwbHjHmOT6O/GpXujuXAnSY6VTt5yw5Wp1jDkLbe
m2B0UDGeVNDFX+NHWG6v0+pcjPeisn/50m8+TMuvdRxO2lKmYqx5Te7sGbBHq22g7hVDopp41Cmr
V8m/5WFchZsYwc4iOFOY2ci2SVfAmdh985/7U09AZmiRxZ72ybaChwYHOP49mwmm3UwGKQtfgSIL
sLdsD0OOYdsSA7l8tP0E5Ia/Z8UKJ6VhSLjpEK8QIZB601PixlMEVmRQmgtVvFVg2PFWQ6u3SXwf
5dgUmCoA4WvXrzkjkTyhBXFJovUOPmDNp88thuY2PLVM3kbcbuCJLlZBAkRio7bf/VDSl1QV1S16
qpIxuNYiX7XYjC/FuVldigcGEDf+QnbKabW1JsQ4J/rV9/2kpYjAZW4iGvUifw6idmbquwxRpCAZ
2mnXwtk7f5o+a8jiVM+sOfOSkTROuWrnUPx0vcOVVzKjuf+jIJLpVD/9KJ+rzdQwIKZriqr0LaTz
reScBOh55+xkX9wYqY4tqnhZJnV+Y5f9BUSAwYxOMAWw414g1sM1OXr3SKOgh7VEydGc3IUQFFrb
UclQYhPSCVvUsuAAsxiEF8YvA1FCIL9VN22Oc6tTjVYjKn/6qpo6JXE3AEBZ01k+40/9Pjkmn8/4
2lWOmKfsytj5hVQXv9MXo5ZOzn5m9SOQy19DElVUwsoV2hRKK8por2cPDwXzjLIz3yvDCH+QQ9DG
yR6a1h1+/PwYxb9XG6PJfplzRq1w3vxYRwWh21rjvq73ZGOOGxCRM//9V0Fb1l58c+B21IFV9U5V
OW7y7E8ZK2uqEcuEJi+Eoj1PDIcsktYGtwDIyF6l2+va3ddBXO16C7Qt+rnquVpGwFgRSwjjPBY/
cP07+OtVP1+RF9bmagW9jIjsHm90UaDoP2g5io31FzzoCbGldfqpsgdj8loBmoLIGXPdFITWaiew
mGLdNq49gcaE+fHtsZC4//E7e9uNj6UfayPGzercB2hBOUCAxQGWBXd9VQ0v6Cq/9NSuLPYcNqFv
lZPKJIByrE4dKltFUY0Br4u6/uG9Q1B5kyI0AAw0ZvOpK18n9jc9lCB3crOaWYR2glzYEZZFhfht
c3LVnW2cQL4Mt5KOjIY6x8nfKV915aSeUikc+O5lcbgEcemWtcJ3R9SFMGrG77SktWgUBrkAkaFZ
3I2iSi7fpwwVwS8rCR667zfS//JtKxgBkxu0PNXY9Nex5X+zvVFz+QL0TzgV1mkfniC1ynURVndd
QOdPzE4v45ojg+vrVxobZ1/KSJFIDoxrE8kMN/AbD4R6+4G8QZep5YQQGiv1XLwMbb1CXWNrvMti
zY81NNFJyNL2mZFwzuzxnUXAZiQkcbCOTglsni269ZtHpZaW/ief7s4WLDP88QZFFHJEyhw72H+s
uSqy4zyAPAQMzixbCDIAqjW/BvdTpjCl3pBodsZ9ucfiPU1Q8MQl8eyhEGVBzwabGFmZajvJV3da
eO+LgmyF/JTuoUPFryA0KJtsP+NihquxRF2INRlCQ3OegodYRBZocbJgg+fDHrkHyClkBEWO9uRX
N/cRA+HtseaFnf+kuI+BwY6EQPR71fhjq6qdew393Yy9mMeTkQVV2v1yGeWXsDwQYQ8EGSMfTSD7
4SYsxzOmlLBIBjc9ExiXZI2mjZ9s+dbq1UdKgy6d8oVMrcqD8BP7UC4EVcpzlBVyKSImKUBUpwBK
wuE2rC9LuMKB0v1t6f+7JihT5fYMHiUXrLoMoNDAZdO8bJ56al4L+UKWcY+0anI4G/85h5UIXV9O
G74ljH3UD16LoN2GU3shIj35qWToGvyl+UI4Vs8e5GatUq3rgZMoYYxoepzTaelyQnChWoGYxr3L
58JLa7XtkxqbiuO1zTlAmupu1BUp92GuY4K1MQRP+jJ0vhE+6esOsGuHBXSh4Zwc9+jINyTXQvkg
ilaA4rLntgQolaTWEXffPwJTTN6T7mXFdXlzeoqjrQc5u4urwjBjhcmT3hnu2cWaFkkiQmkHkqqb
rVxqNUkFLu9fdwUZBOpNwMpiwb7MO5hbagBTl8ZEJS/k8pn63OamMUfZG2Cy2le6sDvpFLuoNOop
93JkBNU+UXvU3zuwyQefdRIE9LbkiQBAfDkP5Q7oNY3G1F3NwYohBfZgVa3iJa1u7ld8CFk/mOFD
xk43bk8HonZzHS+AY/nHTKmCA4aJZnNTteP0Ut7NhA0dDLoVKKwhpIGhFx7ufrbLj6TCqKHGWzUd
ug/3Rs0RdU0luW89r4AYAb0I/E+QWFZU6szlkmYAcBbUsX6LXC2CYz8VB7QWsYEnNqUzcxWTWeTB
pzKUqpcXkWjy1wHi6laGC2OsjqxqviokdSNJC2xDhyxBkrRaBdPOB3SfscgrhfE+vzat+yy5xGyQ
NJblVKIpk+ZC8SF9vJZqDaEPPACLUuCEX6FPGV9PfL1PyBQ0aDMNmusUn7gFALPHiOpeDWMlNNci
6+TWuF9kyl7xXiZy3KvTQc0CXRlWEZRs/Rv++ualdQNl1mLS+Sd76VI1VXqPpB+s3BMC8NqnDtZl
ndbC2TU18dFWhPUHNtziBHb2rV1NtQp6t4AVe+c5LsHX0vZibZGf3hz0Dlk/gQd5UQ+/7mqtJhwg
yfRYEsn17Yff43BBjLdMTugrzp+ONpCEN4OGHTUSoeb3Bs4d0JVOALd1H5jkKqO6nXO7S2cL2V2Z
0OCDchQuj2mlmIeoO/8rkCsho7UhurqVka++oct3ln85D8EUMXi6zjqjCVCS3tbKxKkYsE7gOVOw
Fj3p3qspWOCEF089vO+DPhEtxr5bQi7KfRkpSh0r5WuWmjkeUnqlR00D0CmX4KQ57a8Xjf4AOcpi
+QZsTkKS31+ydoOdeYYIQF4LhkoQHCVk6bFvmddegGwkn2kmvcESyL+5/wVJNXepjDQ4yttDNwwv
M8AC1IDK5F7oIoOsWUwkgROECx2XgMYBCzq96F/z6RdTNoI0Fs6r8E6XF4S46bfI32riOrU2wEV0
0EkjEpY+oJSFNXhiIruZxlUCKwjLn+gURnaW9MHbhWhPfBH93LSCnsgytSRcxHRMSvvOQCYzS6Ji
Zg/ZN6xa8RfLTOwr8tNK6scNrrSAD7YuLMsDVTMkpL1MK5yoQX6lJFhEotzc/HQzbM61TMKGJrGc
n2P6X+HDRHYvzHRy6BzczC5+ZVk80dTa2lixN1oKFkFjITJ4w8JQs0YA3J1hqJ5BtrvM0II0bNPx
PMqUZVhiCLY+0OxPFBMC9baCsTidcGvI1N1pOHWKuZACWSJMbpcxj3tB+J6RCTBAyC1GurOkxfOP
p5pPope0Ald5CmUoBb0/+WfSt648hdZkGqU1jK47RIQwfbY28C9inIFLNWqJ6AEWPX/8aTZHphuU
2AEh/k/vYok1GYx7gegmnRoT7GVKM7bmc0ex8WQ0/zGMGz6KFiEDqnc6tzJrvevZh/Ck3xRUhQaE
cD3YBV2EHKnAVfO8kxCck+OVioTHXtvYURqLLhRuXC3NffMWX6BGit/silCyf0ImNspKLevNwV46
ZUQu06a7Gf6OBRC2WNTXNbCC0nE0SuXym1W8Tgtj3mYpsnAYbQ+r7JvH7WHNBQN91AiI2rJ0PbEh
izFayJRdbqFSt0zE1+MPe4m0EhYjt1dQ3+TOnf00s1jVc9nqtrtOL0JwrGm7L+9x8CaswOTQ05L1
XFhi4wHlxRstXqzTxl7kXfHbkkJAbYnYZk9EG8nCvHoiIk18vhSehckvV6V78YJERCDbh77/G7Pf
YgnIA7aQwWQJcQn9o0eDlKetvmqp/IBODiwT1KnJVH7yTaoxlRqkWCRDkIhFZ+ZrLnWNAsxU+Wtm
8k70pdSRPcxnr7zzjMiQasHycHXswdT7RqfinSRYc5nfGaJrTtIOQhTF9nxAk5rKVE9H7gGxApn/
WdmJoD63qjMZrVndBpnt4VqgRfaTiIMXVoc5ryW/5Nwt7FK85tCJgiGEVjoizBIYfPctvq8AHnRj
KdN1DT4kwtQQo9BZaMOeknu5oL1x9/KgulCR40W4Gw3shV4Miai1D6A1XziXPofTR24cSg9a+RQH
Z2zSbDnif5cB56v4tWzudRsOilGi3VMZB0t4j03jXYpLMWD+92w3Hz61TufEyW+FUKlukw6MEO1o
lREq1ktl0BkoTCV/zaAalVz6mcksYn1OqihW0GDZvn+g3KRV1uMoqdDnbo/xd2rDjOT3AzOyaJJe
CReed4+34xIC6wznHxDJTFoS/DUmogO+sap+xeJQ37SFGRSGxoaJefj544pSI8Kc98c8lzcOH5hX
6I0WQhwEkoZvFh41Kn1dqBXt0q5gPeD41ShkcEOz0nlYYVeoTl7KwvpfP6HOF+qBeOwdDIpN84li
aFwyONcO5EHbD1Mqw7ewxiqwDJ38NX4UhYEvBC050tIbBcX7F4qoMu9VNMPjbPOoB5ua8v0l+/Md
7gNhv4nRMx3EGYq1lioaZmeooqgJO1LHrwu5gZG8Szcq+1Y7jOuVPzQYnpVDdLbdhxrUd2yUP8LC
i+iaMOqzQDG+fFNWlxDKHkvdCzy9oX8MwQx82JTy+/kbdmqJ5JbnHlDeqgJW6EkvwQ97ZN1HrL/h
qoaqZ+B9Jg33fQVImSeODBa9w7JXUKMmsUFu0SnJadjuvgYXOWg+KV2tAU0C/9+/1Bxu0xygbgad
8sx1/tEZT/3nO8r6/0MoD2yzXRhWra5dyWS1GcWpwB+CxDYg2xeAAg4EN5ORNq3btVlnHHlIo8Gs
oz9INhtx7AquYG9VWIduH+qJWt5IS+yeMwYdK9EPXB9GqKLGZ0ZGmnSYPdpP1z0mcw5offMXDC58
ewAz6EJJrynOesEax2t43rg7bNO4usef9ekKt8suRIvHSLx9iQqAMrJ9ovJk+8mDER/A1Q3AL0td
tara613qh4ViMnZKP/+nwfv/NmUgp5tOmFiuz+HKYk1/8l/9fzHX2b4Ufqh3XMZSHw77w7Kt0kZd
MqiIwOlCc8AFM0NpZfNDgxW5c2btOsYXjC19A2LNZVr8mcMjYJDtZlp+VY92iDzZj3OQt2uA4R0Y
PExo8wdf9+FSP4Lly2gHDZCaQ6Xwj9fNbFtuI18cX/G4F8tSuxLeGPcLP71YRGnxchmbf98ZcV3a
T9EO8SGzKC7Bq78pjCnwQ5GulissynDnh+k0QcuG436e8sXCKpIP1HHxKMoHvHV7UHtoT2KgGr6x
I/NF+DWGChwzz0jXR+0bI0jdtexa1tds9JFackDyX4OlgZdYY3Cs71M5QLaVOKH0yV1+2U3RNpKL
V2GITEwxjfYln7uTiGwpli8QY/+HpnnBhQKk78M3v5p7q4eHMCoJ9AohOCYHGOjvK7SB4Aow9F3C
4+CJK+yeDxp66IE2G519zg6iM5tjSzaKco9vJ6HJ9SbkjbSi1axwttBorixhVL4Xq6IsRgd8KFTT
FmvJ2p03uqcxPP4bwo7/Fbph9bFKrPb8sGbZEFB4M+4nfgSwzGmkylG9mcfxovsJpGVP4+uyavwz
UOmhCZqvZRH/j0Gp9yM8PWG7CCNhLUibOyLgKgE61o14bcTfczy5sn1yLwEDN9kvK1rEG6M/wCzX
lFHWlRciiPvYg012B8Bacexmgqm18q8KhwsUe8Ug8ZDNyRfb7+9yT/mFuntKQ0fjnzmBEkvVQx/m
mOHaoiMum9lRJvxE7V4CukCDHS8Hcmm/kX/yGWoGvnXi2kCnx9svchFmboIpP7jxM0/u4B/4E8m/
2mKJjtSh/9t5//QtvK16xwSQwJFCkeq4+l91I3PLIlYsweQPQvR/CWwP5MxoGKmfGMZJ/ywU9D6v
AW0CNyVdlOBsyaWvbwZ/1kQxfza6u2eVwfnq0dfZoCfvcpQXaLO57RxVWvHc1Eet8FegmeUnKhpt
QUXNseFD24Z4N6oQ2Ll4qQ+eyGKv9Fq/45ZNC4700k9RWAWizuGD/S3q8341AJAek1XosKv52xLo
m3OJCdknhkIV+hkaKCh/3cDCzpbduKM4hWnYKTgH/BOhiQMnq9yRfkLhFqNvSnbUEDY6OauhUXFU
ZoJLBabut7HXi1p8FBmm8K9U7fEZqfh1GCrsxo/DCIiJVwEKA8iCJJVrD4UofJ8cFr3lL+TJ7PvJ
x1E1bsXIa1AvBfB4f/exCfTZ+KWWAQIb+V8DTktcP1+1q4tieaUzaXi27sSXj5iADMKd/uAv3qTy
xJHskbCVsTc9duz9LOWkW7RUeFLQQ5mM3wNczsyllZyv+86PyCZpcHIdFf7L06DGby7Fpa+E4laA
qPrGClReqgx8gclpWoNvwvUxYZGTzVeN8oopyCFW8T1irB5tTP9bBCIYPLZ8zPJ1Nsg5LZ4DW20l
/eoglQJICGP2PibnNrWKkixEhAfsfDTXht53Fe0qD8C8/8AmIERpQ2YXs/kpJFfyrrG50np2LNQ2
8lJF6RPe3uHmsEkxsPa0iBQYv8R5OItrbUSRu5A6V40qns+ZtzNxLrkEsvFn+vBftpz9zvtLtBpV
OMBsbqA8mwNk0RbtY8dBTc27PDMq68/lbhP3jq54J0qGCuJYlSxuOc1t9QvpgG3cwTUGHumLgs0U
jlImnkB21U5/2uMOtOpfsC++jtTJSXY5TVvj+lxc2sSyWTFT7EnmJfymCqbK1rU3V2OkNdRcSpl7
Gyq2MWX35I2Cd8kFp/aGY+G6J+oSFiLJmB87AJlAX7gwbrgPzS3E8lj/WsjIWTX9CjzZ4rt1WrDj
opbRgJkaLRekuPRXbBf7nGOCOtkcgn2KuTQH7n4SB4GBo/yDWM5b8BVCq2mmfVPlSer6pygUEEFZ
1s+/Y7jYtGbs5z2KYGApUV+3fa3YaIpvL97rkwjLi1K0oEL/o9jcYKMlZ+YnDRQ/aWoozjp5rGi+
R0hdEDem00DsPwuhhwCM15cMcMOWKNwcZczKvQIJLLlyW56nw2gdrsF//Ec8x1TSDQYZPmxrH+Eb
bNoUyGT6AUxUOlhLLW3+hROmQisz3Jcu29USDnVgRUSPiY7ZAWZW/Zh0NeK8OU87n8HgL61cBjxN
gmyb18yKTIBlem0bKC7l+FPcMhkoHFOI/m4h6Dtpw2AUq2Do1WrcTh4WKQi9g7kS0MQ20WdRoHbr
csVxhfd696n9SzOBJdmpTJ2O3VfdxSMcpidPq9w8jZbQDDhRjFXcVlV2uQV3cdfYbb8V2NKU4a3W
FwWNZ+WhNIkEaxPuvBK9i7dOKKq9M2h/oIlLe6seI2bDO1HISHWenTXtOQQNkhFkN80nN6BjQaO7
2dfteyDQZYTDdbuMSyA2Us7QdxU4pTAf4suwIQ8wtL3V3fc+AiiE+JVUkTdfaUPLZvh7n6eT9VgO
0c1ru4HudkD6e7qkoHPnODsMIyLZQQ+sCgBht2v8/34k4+BBqeHrXnAN6jKh+/w/2d/WjjvUin1A
6c77Tc5B7ibThrGX2k/Cmy34XtvZW+V015eXn5b/6nuVSf6kvpURcBmu2NGSjk3WR2wuq3w94sky
/LiD4KnNmVuaXqYfXCnge8IGw3gaAvYKtrl55OehVudAXE/GT58TT7C6LXpGXMvUEK77cA7KOHZo
QfDiHCBUtBRnuW9gPxi0Mucpryw/0V/WQYMde1pqCSxptyxPMttQj/UXapCBZCQdZHrGsZsq1uxy
vY34I8ly4wPF4d+fNGfdFlIWSMoPj46IpPYCX9aGoN+IztOqj5jGEVONpb6XFD86HBmms9B1f9T5
EvGDhXOsTEZO7+JieZ+Whgr0eC+I98odGpwYHModSaBl8A2QfzT18a/yT2NajftQ/ziYXHbFKkYW
E2nbQlOV9EIq//8gSsLJfxCC1aODBWL3RYmd0bci7BEw0+nBIODn1TrTOUSau6llKvJbBouQpTQG
BqmoScggOJ58gIgTyagex7nfc1a2hH9EBtkLxxN/VjmhXgEdzXG4sz2fRgeYuR1PpUVVoE1UeV74
qY5H7TdFAsKqwVfq6iTL4mC/stxgOKbONtEn8fggSNpMObtxB3eBoMBO5nxaRrTVLa/85RssY6tN
Bfom5SP3hcvYgSHu1fO2o22Py5COc5QtwrAlW4VoSiYt6i9YdxhK1eJZYeNqrj/66UF+5XIB86VG
TS7ckOA8JctrTHhBCawlvTz+ctg87L9ikfZPHBin3D4r02+si0Trrt0LM2dgdOEbu/wJdOHcfF+K
4V+jB7M396ZNktMmykRJByQ7t3bFuRcFbWFbRN443XnJQ4p+GodhuHKb4CbGy2xAU0s35wMMNzg1
jcN3M+FULO+5fuzaHaWJhonHbmYs8rwP+B2+iTI+SIzK0ji17bhmAvEH0mXy5cUsA9a0Wr7OJ6Ts
GmRmJUVjgyk4A9MP6j4J85SGY41wSjZKUwpLcz2EhBb+wq8PFHMgcV35ARKEYsw0sjzElgaT6PVU
NKP8DuYRlpiUe5ansGDUji74eujtNPQNNa/LPrQscUZCV+pmhTYU6vmb4y23zrGsf48DP8jTE5AX
DzhJ2Sp7f7+JA93haKS+LeWUOuAZq4mbGsOf/b/wG+KXyaRAvsymMi67XBqOC4Tk16wI5pN28PSa
i0yYj5wKEXmBQejmEFp46M4HbewZUY5VirmNd1zEF8c91/Eh7EczBsXEGANjfTkGPgIO4N4A7f4h
MHhKkzE2vir84mJkSl6sQFmUHud7U8CpHwSzmmqGKYxQft6w1LvtRYpJoS4UXlfg7achayTC3+tQ
7HKqJPUAzft564zl98tHUT5KTKj/dUVQV4ch563HPVaxA3GYCOZAl1drwMUD1xIgPiV08sCAuK9c
5t3H7O6fX4NmlhcDIHWFIgwEJnmqvkSoMAcpNn/ueXl80QBZILJ/okXFUXRqV4rMg9mrKeRtsCBm
ExdmytvE0k6QksrITjJnQo+s2DrGAmVS8g0r2o1s0+z6IInhJOReJOgp5+VQ534V1bp9rvbrhXrq
YDZs4UIERMfvAGex0+NhKOLLDZRnvfQRKYc2UrtfcenuklEzsTtKK9kdRF0xwY07k3bZUdJbS0Rk
hPdNrD1bZh5Intdi7oEAYI8eG9D2vVA5RmCqowZ9Xg+4b79Ys6B1LnerzNOfjapAZVPLs7qQGjsq
ydDemu19SpsVr1+RJOIsnspUSe4pP9HC2zbGdrAUd0M1NllcL3gmsSsM2/tiGDq/J1oT/GOx5m03
26JiU68Q5nINfGeTDHmlSsbjjPTYMaKcVTOL5KVDKQy75R9WU3JPgbQB+k2q50n1JQtWmG4vDygI
dFwQi5qDLU81W+heNJ9kCZQuN6U3N3XAM8HDTf7E+3xaUJ6xg7B05JHA9FOfI+Lln8qV0K9Bk1bt
lAV2oCoTTsm0ERBVbBcYA72GYePZJYGgFNa3iDZG8OU+vEBnZtacGl+g+MpAaPuoK0qpN/QdHSW7
FSpRmLxgy63yAfroWwU1EbDds2oZITijz57LqmtfmTDM8fOVbmOdurOufvYzxlS2JDpon2802lhw
3/OrklZ0vKLe+vWT6TM0wIQOB9xd8QHB3CpV0FEgiwt+7fBVW2eGZ2IQFCX5X3PRzxIIbltuTkTw
KhuMuT9AxIHFaM5gwGps/o3lFzdn2JYrev6ztPCYFeEkQScNL89L4hBWI/vr7qmNGZlrUC9fac1v
GA9zee4vTnxsv1hdi4WCQbyOpLh4gNjbuwOUReAXCWWtIfzb67xYLBBY4PmU+8G0tuyvbc5qd/x3
qet7ogt3WxGmaPOb7uTWV+Kzn4f7J6XUAHQC1t09B6mwo8K28r+pR1GVv4Z/RUlfTxbCLEHTUMZU
2VBf59qXgzgS/UPKhLOrw8Aofph7ljcvYIrCZQDYRmat6PDIavFuOT/jlNN05WcvavoD1FPeyyXx
5u0t8vFsNFx7kyacLvePZpaHxpKjldWj/FozZ405oTfSaH1W38l4SjXMGRXxHhdukavn8C5a7IZQ
Vki7Gnhw7z6RcsoRhHm0EG6xQBMFTR2SKYeV5ylUvKHy5UQpV/UdobG9qdptNzGNwZRNLSu3gN7d
bsbzosaFGwv+87H+pm2+L8jJI3+oZgCY1gLJpjcoHEScYC7VsL/BZtYF4S4OAo2fc1x7qyYi7goD
tte4v/Rj6CIBPNvmlPOgcNHX8opxvDhUAVIa6Ys7CSJtbYBSbb00P1cp9XLcJX/+7rYkukAgXspn
VF0ce+PRpC4ihd+Rl974597FK21DUpzgpUymFNP2qoGU3Qr9t7i4TSZt7H1GvI6eq5NO0UVLjNL1
fPjhVAKd9Ix66ER8HHyxS3m8vNwWLuwp8H024st3KOqT6Jg7LswpVeQFv0ZD3RkAQdC/uXqncp5M
0yIISKVZltEMEKSM+cgrccMQIjIrm+X/UwvVqySSwRvz95P0+piJDXqYV/QjAjGA1zwL0P2o1FkP
vv24K+a+7H2fJzruEB1JwhsVGbKroLYaFdl/A31RkbL3an4TyiFbevGFIUl2rWcZ/xw4d1GYiYbn
YWOGYB3MZhAwXkXveME9sRRsoErQZ/BAhPys4wsKtUV0XDgs6DdS3TTHkuYDtkGoy0dfsaWTtb1i
9X/e+OSwePyK6c5J5hSwneiM6qmUoE0Q12P1YS8A139dNBXqpTp7T2AZYgXSgWj+y+e5Je6WRw4P
vUgglZC/FjNmjInELhg0r8bzSBF0Iq0Nz49QSsICzwmnn3stk6z853UfkXDoiTyeOlKo5XrbfYc/
MNfuczEfdy0Ir9HrOLqjmv7pVm4jrEw1IrHMz8NrKggebTl68jq3Q/H1gNdscKUYvKH1aQE3fLnH
5MgAWolN2RjkpgS1ai+4CkDdGsy4uZNhRwpiuYq46YAAoK3vYz118kkfufBhAgDE3U8FTOboDd57
3GeTOGs8C4b2Q1tiWWTdyorgq+DnFxZFK0MqzOim1xtEmQlHjMboTlhpmKgcANYnNcAYdYENlbAM
vua7COEj5QQRpBfJ4Aq/nm2bVvLEkHPcRZcmHY6qpESl8Z45JRE3/rZfLJdv0v0OHHY/5awI07PD
4Q0jDqKrEx8oMuYHeP+ChWRl11Qqj/Cf58h4qharnqJoWzfRjQr0s3UQXyJqf7+uslsW0VfcShWu
wt0QkAXizqoVh1/hay80o7gbYebREQ7jpf6/UI2CvNbuN/WkXDwlx6VEuNONGOu7xrPL6HSvrEeF
3hOwJJSJ2lvbQc41QMfq1KHfNdltDWyAjFmwAE04YQJQXtCCRizWAym6j0f9IJLKpTclpAgX/rEz
tCVIgHui9P5rhro6POiIEsnp6W4+f9T+AtD1VfQpFIktxINotulYohupK/95/SQrsiahQpadaboJ
e6fvHTwFCdwiP+3VS3KvbXxyvn5i2BOM4CteP4mlRwpanLphktw6ZL85K1pVSbJUdB9UDTUVTtAN
K2nvqP9q/QBeQs3nuRpf48OUTzf5F6kjYfkrAqIcfEt+vg10PchLuy0O+vn5VsgKxAIaK1S2jlTM
yUsJfUMgkcF3xI6X0sFHiJwt5kXFEUFNHWhSW92Tb+Z0JqwDuCGvSNEE23To/BVjUrYG0iRQgurB
wWWj/0Vc2JLdFFIB8tpkWSn/SNvjD+JpR9P5qWxLXQHXq4NGdrlbMuprc1OYpQeyCymjT/f0M1IA
y1HMSoyxnA099ZsgpR3k2DEbglzDoNXLTu7uV9LygWv0sWSyNAwqw/EgTLORlY5oduyqxnZKQKHw
ZM7oaduCA9VXxCBeFL7pwZ9BexJA1StSFw1RGaAB6MOgviSVZbGf9CoR8qQyKeExATCq26EWuTF4
LzKQy7cQA37oKkTlxvWdun6/Fm0COJ1j2AnVLuanLURTzKz7d6WwKWpcRmZfP16s2m/p1mXeSJ+X
XLkssRcxNlZPx2NnRvgu//Lcy9SeLzrOqepYjtrQCl9pGFc0C+Dj9CL5i8ZBwmjwNtQo0mzPEHI6
ygeJ/pNsRzG805zZ13YryZvUyIg9tT2TodG2XLXCujljEz6irykBSDpnHyV1ki3fqcNkn6YoLged
D5VMgWq+epGuM+AyIBzFxjv0X2cB/1kJY4WEIaEaO+t3d0mL5ViwijFqchsGoYFjy97LbxrWMkyk
3+aqD34jHaMbvwwzsWfbkI3OKn0Vybs9JqulPsmIFLRdGrjXhvu7WEDanphO4NUAtPiBUAOD966f
0Yk3wHMbdB4RAt/Y4ex44IHmZpC6QEbTZZB/gxpfc6s76DUXNhyHDb0fsTZJ/DcIU2RdwPpfm6f4
uMd2M/Y7gnzLbmZCp6MHN0Lovhpzialepsh7T5bzHepnhPAnZs4d63gdioSJ/6yMALsJvy7mnt/B
sRs7u3skFLh7rb0NdyjEAGj+jYokzdosPyrH6vG8jqBg1+7a4rMDK6G9oRkNI8SUnsOkSHYVfsaE
LV4pxeegZH4B638lUHLX812aF9oZiJCVgNbwQucC1ssH52ZEG34JsB0lir38JOK5Vz17NXaeZ9m2
5as9YQTUotLgLyiea5CJxDGVRp1u6e5Wo0+zvUE40g7yrpt3s+jHspjiuCgDZCBo2aoH8ai1mx9+
26mWdZz3rBgYKX2Ad/tEe3A9JczVyG+xlIdWqW/eFQHsYi5/S6bnfaF4leT4GKkfxVqK1vTBKjCJ
dqDi3Z8KHyoOq3A08Xsx+JammFO/hnMpYme8aU6GD04bdP+BTSRmL3bsftTz6vyV2TGuv+sEKPLZ
pZvCqmbb6b66yLf048BrvDyVH/9xYVFktKrk8eWCH7fIxTA2/0ECor2E/WhpHAarWZLdAG96Dwh5
Y99c1UfmDzMO8WrI36Ce1S2mqNmrKqDRPRDDDjLu0b9yoYBJGES+fqyoR+mZVBMbwbykYNcuWvbk
CjYLHoGM8f1NyJC5Pbe56QEqdDCyxa5Fn2XmEB9yG6DbuLztqaI57P5EIf1eBz0cSUsHwmuAN1rh
8sGcurWezNa/OYV1QyCXwcHNLbMwhsjr+j0PN/736La33aszpZVV7eHI/LH8NzJ661pbVe5aoZKu
5n47DJmYyqD/WT/K3J3CBUvAmsItnSJzXjaNyvbLquBNwN+6LJgsV11eDhmG+7UZlvIBDq9ZgR8Q
agTT1vuv5ZZJK9a7KXJ7RbTTQqhIdDXZ4IgjEj2oEthWE1mTlXYKNpKi6vjMFLXi0pCUL4mBHu/0
oKpPjVsyLkcXTAFhDuZKhASKtLDtOotOnJJ0JxrH7MhMTbw6jSuDrST+WnuC8Wc+1I9SiC0To7ks
qvwtrP/dHm7lPfDjTpld2kJU3o+VUjeGKQyK2By39/ctjLRfl4YMZksh70HeaY86TuJGAXelYxjT
Z9vun0jHNkD16m31zLaSZlYtjfIbab8SQ0f4iGo6S9D8Hj96NoxyeMOQKKf1wNo0rE5o0aVWFS5s
EIdVw7Axb4XHKvRENtuWa16SiBsvdpsTYpDhULvdfsXyuRXW4hiH3Qa283JiD7ekXi5ZKfm28VaK
F2ID9qPSjwTpoWvnKyxbFqzaPQU3oTGYNuZansGzAY6MN3fqvLg3Pp4R1AigzLYCYgtbEiXeOc6m
kixTzqj8kL4RnlVxrvKrkR4mBay0lYONiHwWgf0fWWrKUDkabCTTbXnoqREsUOwHqCvuRYXYQuuI
twOYvetH6FLR0LWCODYHLRP9J9W6xtTzekMTRwl/l3VKb0uqhgO6ugQ8HChpAoiWI3/v5lxeBLH+
t48Mtw3ZPR0kMMGE8kSZFO5M20ib77VlX/idhO5XN1XDBnFZ9hKz0XcF6iA2+6UvCvO9a6hHEEHA
ZnzXic0NE+H5p7VAMq8EWDlfNWbJqWzOky+dIyL+y3Bf5a6dMGHVmDdkFnZ/lbnTV0JoZluDz+S6
FQpo+l2qwNnOl9mfgop+cB2WqI1SWW6eXxQrnz1flIDLnmzfKpP/nhTrqk0R2V9L75lD6vfuQ3mb
9RpDK9rI+QcgHZxzaCNMkPjRDuoRuLz8sgIjZmfqqEb/Bzc1vkmxzDglv0PiKXGsj8yTJKAzl982
dzgdkf/flCfHPxSDQphoRL6feEDXOIT9rBRYjZiXLbOAgXfAXwCgz+DWngKOZNphGm4Hh1xZ/6ie
9hxNU4VZDJ59xr+oej0xWW7w4cyTQ8m1yTSoJf8O5PbF3PpEhNLydT40A/ynb+HTV6HYMokQM7Gu
MHYN8R7+IMeU8wlFIVyFXqbBlQOSrEfYEnl9iDCwzMX4yeOclZfpWDsM2z8wLDWvFCyTiGviQyOA
FWsdfapdOnrfYtavJa5F1tk+FEvPkh5Nu3Uu9zZLmsZs1lvPcZbTcw2aLaBPbXLWs8X49yyADG1K
yFxpa5PNSFIChPCIg/yX+IwfStGekRpEzXRxwcfHuq53bRNfl14h01PtVOFITg3yplEc87row3ki
1GwtTWTpWZ6Vy8lpf+K691wcLbCVX2wxjLBHkE4TkvfIpf07q5GPRCKfT1BgFu6NjRKl7BjZCyYu
PD91D+aL91u/ls3xspQ03saX+eVGP+YGH+NrxYNjYJEW4PrKzxSDREugfQVxFnC/36oNu1oUVgUa
8H1lE3IumMsBY/tyzS8/pesaIz3yzPILYhNs9p2sazSb+efso30OwLX+bhluZkr7/v5HM0vBVdfT
jr4DxvU5NGSdzaM7d9XoOFwPFIOgoI64C9ZNJp75J4xlpUMnLvpCL7btnfAfnFv6sxbqq4Zezngu
I0Br2e/xumrLpub96BsP/3rQcbyngjPlhq904gEy6zpkmciO5caodam8obZKbHlHeievCBEVyPXh
2wCJRX7+trufC5NmdzdfaiV0mgpr2jDJPzB2wrCg17DnOz3MYD6bZn6MRH+0Ixs/ZQkB0kJurkqG
f/rf7vbD6j97wgiNkAXqMZidhFcIFciAW8PdxAXE1/7URqxLoyoCRJTUvFep7Nl0P44bIrF8uuTr
7AYxRYmcMvMGAQ7nJY5o/94aFi1kSyxfN525BTtyrd/ZkbEFfg1QE/ug6BMxhWwT4ugpzsho8OnK
B3q3uC40uGvaWZPf9OG4XuIyLqLfMfWNjIROTFE48l8LatP7e01B8v61eR7Do4iAL6Uq7Wdg0fvg
+VLMxFoR6W20INov+l7/q7PV5JlPubI2Wfdv10706/wa9k0/JslhzBjG7j2l+NEzNXgmGj4wLTO3
LTuLXKJ2YslHRS3zWKlTN2ZX6Dd+q33kCpJ3VrTklskgrHX3ody8/a7nMWYx1WArbdZEr1hJMj6n
+AdoGf115urfab4WZr9IUp5r91pvlgPHPm16aLKXXSEPeuDguIQ71wfzGY3hnl1JTtcjS/m9s+6z
luB9mO+a3kI/NkInTPxcnt7yZy+Muq/RPlOPEdvAZ63Wc3x33C83nABial/d+dnAVUZPeokS/7dV
QQXqtnGG6vt+0gughUhd+iGFSU1RmZ0MpqtPxOWUQ+Gd3qSsM/HyT38+zL9pe2QoC3Sb83h3KSea
HzWUr7EObayh3LA2wOXWwD12d/NHmC2H7K/uRYbzl6dFkP9WIENwVUa8/j84V2HrkMoEOwKHuqRM
ORPihas9+Bgf7fIgF+DDcJmsc37b6BCL6tv43RSOfQSLbTUY4j4gJPa95RpgesC7HE4L4aRjJ34o
1mVZ265DgnODAiXJVsB3rZzLsMUECEFpRxWnBs3usfE7sxRB2R+/XcfZ2aXgFsRbNhiSjmRtJOBb
M/wpNCFXQxwqwl7/HrKZgW/WpzBkRfyNYTRvumBxhLtk2OQLJhkHKqRMPEdEtqxuTibjg0pGFRUZ
5ExewMchJlkfHr342erYxGp+JaSP8vUBRZ7IuTIruXlS0OatJOPdpUJHYn3bNz1oJfjq0AWlPpKg
H01/vE/kocf8NaOHhLNkXAp64j/MeT46l72pUF6hg6OGlGVVk5cOOPyqT0R0NOH0G1BL4IFqXQSI
L1Ws2BGwREMiSGiJIMYC7YKbw+EICtFSuuS4Z10WDTYOAkHqpJhp7JzzGlBahCUWFTUz5tUVsX7B
RJWkoWfErNSD2bSk0SFJ+It6iqFB8grzG9hxpfwHbRw1QzXB4l7l58TeapzSZTKPW3NKBIJ1pYy8
2f4mubzHd790YiuOuvxHT5ZbYfrVZTOnSym3JCCvwRrn0eM8DuflgONWBgUZW0SOt2Vidv5pqhKK
GXuR9f00VxPDKaLtylOPiZNWENHho4Jvx1yLQDbG3+5zfCuUuD8UySZNZNjjX1j5TjwLis9+3sH1
//45vMJ4/FU3s67PRXuDIg+Kkdz4icFY7tbhDGsNW0/cpedIrGD8rCKAr5nymLjGLehjtrqtyfWB
Q35l8/ffraduotpqUxIXXcqytwdYA7T1+SWa2D15uIsegdc4izMp6nNFs3C9GRmhOnvD2sXCNZJl
o9BfZVmOEuPopuBW6tYgxgqMTFWhiqaZ29l8g7wFCheu3BRVfgvoAAwHC39BMn0BhFp4JhXibIIu
Vohl18pbyE3cMWcDzstMtisCv9hFltO2k+iyQ3tPxMmZ7U7E4JlQbG4l6ZuG1rYPgwiVP/OR+K5r
cVtOeTiYkhNlsdKDbBf7w/gSEuhvkd5Cfgg+16T4vS0Rnq490bLI6LRqPZ+i7vHM/lTXVDTW4GhB
tKEoK/Kh2cg0LXMTbrRw5ZfQ+dwIDO3s8MWP3eRJKlgf54yacNdAw5XFLkqaj7nzYX/rvvtpjwbY
AGxo6dcfVfJ95fFpt2uPaNe66+c+Vg0pFipoPqqXgoQVn/Fx0Ms6VOdc9LtcI7+pgZr9TAUT2i76
W/w4vmBojmrW1UxqHfatZC/FVyuKNRpWWswVrE3QtyEFaE+ij8MseYTap7R3MOoP4fF26r84eQ+J
pibkjPnWdEBtOdgkYxijGRZJ0gDwBRu+lVAPe8Mq4C8UHZUO9D9Lznu9LwzDLA523sfir/0EURu/
ACPBQPGvRb6ufKbZdQHM71TK4i5exbkJD0/L/mdcEahikV/MEvdBJx+5gESFZyHjeppZNgfJEFwf
WRaDg1g/re4fM4xdexEjyol2N5sxM4sz6NTxtIcC48fUPltex9Cx5p5dek5IqilqNOmhYpW5imvs
0AR8RIfsw66NbS5oMKFUSzkSUqz3U/3f/ZpciOcRIV8/q1Y/D58UwoFXQtXIbRGdVgRZ0PN1Lmhl
648NYzgMJtAkZkHMaZlS2oqEftRtBUNXWaJNqEwbMOtFJPCkG0/5sDhiPRcv5ztGkAB+gQhd+iUO
F73J5zknmyNKzgzcAKsIRb+Jge+KQpxYnnsNkffUDKnha/krMTouYVQvYhd3ZcKEt4TNtYc4mhan
jGI2ioQLcVHBQ6A4NDfKiUF9ItIEWw/xLGnhn+ddikXv2Xkn5V400OYau7aHB03avi4XL4SQQApo
agFPzk9dE85XJ65TzH2IgVP+TVGYOVECiMmAdm14RmsCkb4Zk8MN6zf8lPrrfXwlEeNQ12ku1K3Y
6UQG2HA0kHvzx1kj/aqEaJzur6gDvWG82Pi/KYbqvZZV1F6BjUXZQpq92LVkKiDh0O3w2rLhPVc3
KQfu5UcHxiNFR1jF8hcdcALFjKEjcMuMGUZDn7s6/roK/yPqbRJ6iBfJU4y25jDdvEwlAzHggxB3
pmxtnuiS1t/+iHHSmf0tLsdDoAMBUcBlt58kzjB2ysu3uFvfJw1FSR8tFoUEkxJaOmyBQcxJ93uP
ZFDLqMhSY/fATkgSviVN8WvYb9Ype+Jxxs6IiZ2xC2velsWtx9RIydEJhnGcKWAkyVvImPqRINiD
QiPyEsqttZ0iJ/PgHimGhVldw4rEh30mxFQd4JjhMOthgRPTCKdet5b4toV0AIc4/wJ3Z4MNoxtn
LITtDXEiRfvaYDnC+4/VKu1FDigx+o4oAJ9l3eBlDL9IsqSzPXqcFeXVg5eYpMuwWVGMTOUlyO6W
tVyv+AXi102ArPTsAcae2ZuyNvXg/REGM1MEqkBMP+qrXUCUhcPmHWEZK4K5uN+pu66GjgcA1R2w
oVl2ZrqjZoENO4/0MAMKH7n1cB81OlCSLIyPP4bK8TS/+P5vHj1lVRBwD1dOHKQ0Jfha06TznyBU
gGbC+FDsU4jlVPLNYwJXFbFUGnN48uPn9sP3krzsjmHsu0hshqSamEu8PnssK7ZnqauZAu5sZWrg
jxYLgZGnD+uBeYWqDq2JujfgHrKP9uQH2Ff548yWzZyAawMXACHvKgfzvaKl3TVtiaoWgacnUVGM
TaZMV8v1mvMu4YUK3AvtZp5Lj1Kbr7BjXb5zTzdRDpISVZ/1inX9IkAMWLQfT3B3N36I0VM619VK
TplqsUv2XktUJkw58p325wv0C1jW9filjzVbD16VkKLuY9xmGiFFO/zqaMscbJDwpExFh4cwbpa/
9hpR+eb3ify0e5Qnd+q/9uZktzHFOjGCRLRyzj7F1dpWB5V9AweA9i7lCehau8x7vz42lG3yKrZp
p//ZVBtICNsa90VWjE8kMYnV4kOJe5Ce6Szjzm+8uQldyascd/UZcnJ7duJ5JdG6hKaXEhK3FK/R
dAOImSJqvknh3I7nC5GYBQFyihMeFmp8IadhNl60AJErzNARKqgisSqVWcFXz/yVsIJmzm6LD+Br
EO99lAHYgxBa6eSMeOnZyVrsxH7d0PWO/uoUlUcrMcPKMt984R3SytLV9w4R0mssGtpyd3FXS9io
ZzC5vTenCnXx/8Tj7uS/okEVQ6xKQMZqj/V/i8UqcCj0BVVZePN1Y3Eb+4EOmF/nH6dMshpy0Jak
qOP5eGeOc/+h4O48LMX5UGBzdl/KeviAoCz3qbaoGOhNV7mosko97KuVmRcxoSbsNByH3IHbFLEb
9FqPX5NOkYIskBhN6IZ0Ce8MFUo6OZzj8stmkNX6ASJJvJdMhbO471NFpBNH7YcfrrOBwyQmXvSm
J8qzZrMVMNmyECMV+7YU7r9KTVkDaPQjnbU4b4BbkyeGkQqLqaXxdxMFhOJF93cuhgaXALg09Jvf
5TS0Hm/jFG13V0MfOuqo95iA7bih/WoL0BgKS8iCEND1UQZC7nSsrlhKOmcZpK340OXH+G9Kly4/
UG4I6+h65ga188xNmGHtr4VaWSIWSvn3Np1nE7huo66nncn+bYuolrS9gvyVrMmQ9f8KWCK4SSki
mrD837X0FAScYaD2B8U+M9e91Qiur/D6KIRpvFAoJ0ZkugVAcxVgU0gr8Ilws2VKeKsfjqABK4kZ
0YI5Dy0Ihp1JkSu2/FyxDZSsY/6qOevd2R7jqOc6XAUm3J2fCffdu/3GA5FDGKjQ0yK4o/NIiJSe
SJ/jAQKZh51sAxJsu5YVWQ2n6WuVM35WmY7BdkX23hyE8fn18sCSyxYzDNTVTxzx4+9TDomgqpvr
gbf6ogGBqcM39jD0Bs3IC/KiCEPD61tbVhKm3ER1IEjaVLD8Mebqn9L4C8qCXx95us22UcZ8xQ2V
a6Np7HDCVafaOtHx3sGwCVrDwGp8XNLArSBCfIuy60M6tp64hTRGYD9j3oPK0BmyYyoIbxiYExQy
Qol4xrVzGSh2C1OeM3aWIvBOI00De7aBTaSqEv1v40l3U482svvRQ5SuggzLeK5YJoYcdGsR39Aa
WEKA9ojFZcQFqM/yrqPShvXRwjgus9TmbGXJbmHOpid41p00DEIMEmltCpBEoBXGyea99E1ZWpqG
96zdnzWBO8TIZBu9FkdFNlFF8RsXA4PrrCT/Th40rda4tvQY+1qAlXsS2MF1RN0JRFi0TitZUdVh
tNPax4cMjCOber5iRf1Nwjvp2H0fpWGCyi0S5/QUjDjxxZEeIhw4P9LDSBU4C7oBIG3AnkBjvbkb
RZkAjp2hinSCJ2lnlIoOXfNsSOTSb739VOXiuTYMNJf3g9tbRJCXPi2cDCrJrfkI/j17RM2bLz0J
vwkGqFbgcHYfjj/aemUK91hMFljm57lwnryGOiey9X3T1pvuYMZxqOY6ZkD+VaR2ZCX8Nz0L6rrn
yRIcWKJ+3ZnnpVSrt3oAt3SqLGZDdcflykGVG5Xtyff1cTKKO4EcJs6yj00B2SIo/kF+0o2OKxwS
zE2DdSUGQLszfEMy1I9y6h/ANq5H1LP3FAOrHcIwgKeIHw4tNWiUlq6kBolOt1wr8XtPSybfzd1U
Q7R0B51P4/2UMRPioK3EmpQ4zC+ywJBjM8pCHM3t4PkhlWprm3bPaJoueM6pEcSnlR2R3F3Sv3BW
0f0ucxzboXJ8KRj7dno2LYOqV9lM+zpvPVUaro8sW+EG/175hHEY0AEaY4LiNlxeikHY3X0jKGAG
VOYgof4/kG9IEA1OymsV2LdUh9i+0WL2mzN0czXO+W3P/cY6+h0XstgzbcL+L43d2zCd8C9YegAU
Y/168EbDk6eH4jzF25HSgPaC4FkH9JszaivqtkNNrRmnCXluFgfv5MBKJ5LQOf/ZJJrMvxq0CxVJ
cEUq12Ds5tfCSX4xJdgU8WNyMo5/aAseeKlkaD61WUp9a+wDt1/iw3iJvbWEA/70ARZRuYBYicmu
Ne8RK9Ha20cg3zozpi+0fjh2w1THbGILq49qWV7rF5AMFPSipxZas2ev0CbKWQPeGqTrRP51NbDS
U+ccO5Vq/ZrMBhloX6WW5EG73LY+xB/mMl18iJ5MHrIi+aQA4glmfa8GLQOvEMbyLeRVGN5+BD1z
VjeuBAqDs5C1Z3p4/92jrA15hucOVm761dZgoQWVH25Fhikaj5RqWP5q5NS8OjEqbX2xN5lZSI7q
wCQ5tYhKZIPxqDd7H0FzML21Z5TDRocd9k+j9xJIeT8VynVxJ19Lh6uTR+0FLY9Pv4q8ZmROvXX4
SM+L9pyshYhJjDgjA+XGH3WgWqJxlI5qd4KR0GgRsGJlSFZJlC8KXf0Nkbu4nrdYrJkJBXfynIb6
db8fo9VBVmj/ncFmsiYVMOaOdtH77rY4Premlh0+FOye99QXPhxM9QJ+vfuP5ny7sxSANF5obx51
mOdNdL+FomQmLkHb4Lwa3m9kY6pxtNESAsfSCo4TAluSPq+Yf+K6FsIPqEPDWASTlGQ3vd2e+aTA
0/3X1r+sGCOe/fpiuCGsvUy/htLx2F8y71BF+pZoRuOVATdXdS+mKej9LZ7Vm4BeWxUjovPxk4Fc
u5upEtN2/HeOpdM4paL6u5m+3ov3IEebXfZEqrYN6TJVZho4T0ZmwX31jWngmLQ9SVbfEjnPrn+2
Rj6pStu3kcLUjQ9XYtBVKtZhEuVEXyxlIyHCO2C7qQcejV8bN/l4k7EQgH5yUv1nHrmkblPtSh4k
WsmkGbrxwOQRTCmTw7V0Ezx/j/uS0Pp2kl8gNTZEyPkM71lQEfzP1Fi3QADGnfop57WJAoumaRCV
WskvGASpiJa00HBPg0KMZ7lquB8GjfnVC7jQhlFR3pAmBSyxAD6upkpWZVx0Wt7QPqtf/CRJ9OSL
qTNAM21j0kDmpcOYTuk3+qrIe2DRUZj9Dm2E3sO7aPbRbzp2RqIxN8CDoGUPxf+HA9Dkz0A1gBIW
73cP942Eqgf9nlThiSURS3obfEZJVyP/y6b9CFacRF1i1WihGgExe2oAAg2DisO1XIgMR1MyshXz
oWeRbv1xFTb0qHeJ4mHTKs1W0nBBu4V0+wZBBeL8TgsB1PyZSpfmPtHxOTx8HEs/mtINpkgEPtsY
XXGrEzOYO3XYzYg+lCgpJ6lRaUP2IZlklEtOp4mKOJgJV0sp83ae2rPwMoyPFWU9do8vJ7mf+mcW
0Qfdnp5S4X8V7b6WfemsmUEBRK2vJg3Q9sUqgiOeJ9bbz7JfsST2ATobNNTnejjnCKX/25PV3ldy
9RtmF3aqj6VMBcUrC2KilEItTNiVxeqQ4vXiyddgYNFH2lM4p9i3f1e63e+P07KUtIe4Wfosmuk1
FSSSCreSF4FuksE6gqqfNaE9hzJk3bzy4GP/XlVKxBdkPC0AWme6miM6pHE1IabTHSPY9z/0VdBQ
P5gRuwkm6UDRpJdNDvEch82svEV0cp7vxXoYz/zpHhBf+79BisApdQeJSIfNC43JTdsYLU3j4C4t
7ewzyOpcD4E3NDLwKuUfjIVZWvCcW492Ed4fsUn+X86fnrzZfx/4hvvWcDzLl6JOU3r+HsXn25Ta
yOtOJvc7/om9cB+vOC3pjRlkymEBkUYMY+8pbvsutaUdvJbu0yAOtd777RlHMs4RGeSxq0C3QYRW
c9J+apQ755xmL7hsehNlHf92Bu3Q9qELcwudP/vOyyG5ef6BBBqJ12vmRyLy1gC36oLdZnHyoCjS
2igjMfLjcmexy2DQf5R3lPcMc6YjvVD+VzI+5hGDPrVHV/ut9HtXutGUVUVC32JsB3vV5GhvsrH8
OL5+/QuPUG5L5sl5AVMn/3D+5GvABr64rSxFc+mb/hxJzQkct6KiKzIvgwhuj5XXWU6Nv59SjTpx
IIen9IMSKVYYr3+yCcacl9pH3pxMDS+CFom42a3Qxz28fIxc1xfc953bT8za7mTd0Tl4LdCo6EaE
mhJqNGmHYQ67TlGhIYJWBabmwy/9/2cWQxjxe5wPeQGgOwpeNcuyWhHQRXfCOwFk0LBQd7JPfVtQ
lne4LwrEVmjoNnBxCDXJb9YmOsstuSznj4qjPzy2EAhzne7d2a5gt4D6Dz4EQKKboRopsFX1FIfO
F6TU/S4jY+E9VLwATOkR0ZEgIssXHnvkCUgdadCl3WACfo8Be4+pX+ZQolqIHU+yWU8ixzbwzuBx
+xb+GmbXqY3kJ4wwIbdW2fhl/pj+4NZA6JtLHLf/j0yFGMapocGa+ex7cHPDvcMa/U9DjUJiNMTi
uFV+hMdNSAAz39CipfNKn5TdKMJMg7HTjW2rtHQnIm4nR3GqykNvUtBOFKuIDBFsINAXcGzjYtsr
4rdDMS+bENRZ90CK/g6gSnbv6XAne+cWxRpWEmu7kQmJtrdbs+jysLxoyIfF0cwhoGqRwpdc+QZm
gQs0nvXfV6b0az55IGqYIsMHs3KcQT/SXQ1Olu83apZWdV7GBIHp+qxZnP/hjqqfvdwnch26gn5K
S6B38hXX9vfs6uJWIoXK0PlD+mXmclthNFtTDvS076Z8a6/6zynQTtdZNkf8Fm8phVWqHm0cPI5+
5byYUrZGscRXRshK+aQjLF672slEsnuEGufznDt3WAdXhHyPLCwgtF03a0p/F7LYbAAzOPZYwX3a
NwVsDd5R/X50AV6THLp5hJcbtDYDaE/Ezygkso+zCElCoy9OPNDSRrLx3mia1gcHoZyF4GzlOTe9
bUMpSPFTvGMRl1pIcSGi0xcKFjHlItQeuSt3/5vIzguIRgx+JQWMOENho238pUE16v3P6y1/MDco
aD1dYBA2Jl7HgUdd+y5IKq95z7Q9tNeSoapsN2mD38wqz484Uh+Fu/QxRxpWP0gfSE4qiEvC4dn6
ryqvMW0QZNCX/B7hofmVhS3nB0+p4ZKejgFkTir/QRgkVuvOq3jsuw13fr82SbpNb2ioFf9ljST6
gCAWsF1D5Cs0mYJEDPSkW6GzNRPsK7iLzM37zLCETwkOe227evB4qGEOskd9Qm4FHe48HGwbFHmq
RSt6VYHXfcLUM9zS1DP0Hv9lrrOeWPvAo6DusIgNVPO55Qmp08yhIsuEDe4szGHG5acXrJqfVrQy
77FRPxtdg57qJKTY61wF/L/6ZaSgsZc7VvrjNDorqeOxN2RdrLzxeCNVbevDpeviqc/EukxSnWdv
df4OqPgkT+bGXsU61Cv0uAJyAdw5b8pink4alhpZQIjvXL8isXHLGJesPQkaJmUq+bIR2Hjlt1gk
qBL3hwoe6TN6l7F9K7jyUwnxk5VQKlnzgzP+MOBM6/SrDI78pj97jWVrlAPRJR/za79NgEz+vppt
5639lBQo5SzNh7vXt0jfZlFqYQr7gV5FdM5ffsz7mWI/Lk+/7wXP7vX0vyiJ7iNs1j6ezygWmpaN
TT9yThArWJGo7Q+Herq+U3Ilqi0qL/hbXFf0LoKG6JbKMf6qsqClhU3N/bIuJ1DdY8VjxvSfsN1R
hQl8Z5Cwu8VlMNHqyFQVzqQiHbHfppeqyZzhStZAHH+zaP6gY5lVILzVKVFhmW5H2zuWq4tyARNo
ywgJCOJl2EE7AQCaUu4OI2MCwGfpEAqzW92PisyIYw7VsgFtx0EJzVoMEhmVOG7563loBpohX3FX
RIdAoS9lRrsXqAAbfhVLBtzY9/wyqJDAU9pSFLLihKw2YcqAhkRIzgUY90P1uhJmg6G0/c8nlJb0
u96MAibL8iXw+8sSBdNL2EoavH3JKeTsFqgKeKgBjg3mgMUc8n70eHqA8qDjT4J3Mdoi+8cCqbeb
Btn/tiwGKndcvAJD376HM6qpTI9+gTMHciCC+2PzgLcn2DJLUfiiHxpMu9OQN5Yoz9WxUvbUWrDO
LE9+YPP6mmaJ5BmfEA/y8McUDqNEn+ffNrIiJgE9CctiLfiC1/7d/oIqi46XGiVd5l6A8T6yKr04
BMo5SsvOJfzYgaPKDX0Psdg1Z/Qk0lGSr8qToVHQ5z0zKwAw8Pv03icyOUQjS87MCxGBSjQQh6H8
qEpgY7rrjPgNno1BMjmTf+O0Fp+tJq43c+wYTbH3pas2qHHEsCeCce2+VJA9uXHiDRtaGjzbmHsb
ZmdZq+YfhwtbYvjrlcKKOISivlCGNIfFgpygDteZQlFurPLc4XvivGGNtQynS5tDM7BR4BuQej31
RLy6EO+1fJjEhklRemjwYPIArSMw5L9XrLmsRq3WOA3xFi8gCv84ethmYTDkwILGx9fkAxc5WWaE
TAevnwZ/ezZtDeBmQ94U9GQ0zl/hpgD78+MbnU7fctq1ndMjsuH01HJ8Ef6Fuk0/XG8xymHqU4dV
+Jw6LASUuS+655vAXBL/Mi6vH+FkdK6abN9yakzvZolrlckU72ZKvKRQljk4w0c4cw0PNJnsliAz
obwMHBhSbDJwxonktlWcCRoK1hlD6VD0XKJEkm+6cFDrOgLITNK7JcAwTc7cKyhATZ3szvl/Z8wj
K8ogaG90ZvATkP4Hyq1RhkVDR7lheMLM3Hi31DPXngNev08q7ilzCqo+R0rBdKc/fKjnPLgppaCO
DNFhFliBgxO4wBZYjqLwwdqWiSdIml37FJRgTk/u6R2qbI2JYTO2YFTGXfuooVeHmxz6xaxBeAPy
oedzz8enBuChrE2xvDy+tnWv8xsiqEDrAxPqJPnfgEdSfVI+p+Nutx7IWpW0UgLxHUg0bBMOXDRD
YM1KyPKiXgmoRw8B5w2ByrFRbqb8hYwOjyXqJmFnvYIvS7omew6YlI5zxm4Dx9WtSB5VxxCALuPq
jBXzJGcm5qSLJyeZkQHor8nuJZ9UWxXpSaEamsMfXrM1NWWqi8/Pa4LHa8uqiv4l4/QXL1O6HS5N
3sU9fTkMhfpruBGG+RCVI4gdttuHRjx1Mi7nECTyy8OUVB6S6ujWnE70NgIksKl0H4ZH6K1L+HRL
NGLOOEItNqtUhqf1elEPFAn7z24jY5ZxS9aqnMrEkiTlwwaE00m4M/KqT2dTERiVKOH+3p+vKqAe
7lu42eVSp0++bh4HltaHhNmp1yuXB6XSr8ycCJa0398DtEZdCHmGNT1z+wf+Wl7jtKXg7Grp/A+c
xLhFooanGJvwg+XadcMy2iTk6o7ochSqZVwKguaBtk9EtpiWNMb7vlo7bFYv2dTktVe0TP6Y+Nre
CAkcvV6AHeDnAg23CMNX9MMHSSi1um3k7SfQGVUf1VuVsSPztzDXltcwkDlv6cT+tre+3whw3Hu3
KoW2ZgbwGyGT+aQmh/1hRxs3dbX/EcxlKUMsqUv6QeyuDMs3nOeEpxOlTSeqQXO04YUDHlhA5/Be
D0/yo0ugI6whfLBUSwIKvYNfLh3UT2o0/Dv/zWMPq1glRKCN8NqN1Bzo3a12SR7iZinr3Cyn6Dua
i4a9TkUUSHZWgnXsBhNriFbzeuV0Mex6VQB/2VJymatHhTVgzqqFGD5kwnLxgv0ZPcXEVSU/JDV1
n6DG+Hb+1/Sh5a8JfnsFYwHtVM8LXSwK2jKqC6qelO/PjFJLCCRXliDFUzlNMrfmgrKS1V9sLGfO
+ec/shhD7YFVmdiyAlkXxdTAVUKinC2stW8=
`protect end_protected

