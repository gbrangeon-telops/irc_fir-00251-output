

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gjKSpUobpdaEiN+EJKINegy9RfobWzPNNvSuynmxBaCaiXpZzE42DUdhJsa9nuNl5zrnRUR14CdT
xujtPqnMVQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VxmOSrOiNTkpjQCdEraeE2yE2mnMFQ7pRVDUX9VslB9rFCGD7dNvbneDVpuQoePUk+nSB0IAqnFe
/NakjC9Wt9azzGAltfbGlSpsCZYTQJMARswgnWL4Fmc2+3tN+okF6OFM1YLClj1yRXdxl+CDsxQ1
FBT8tPlhn++ZNTP2k9k=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aXqd6ynCn5cZfxJpxEun0CmjLX7cGy8EmIQDak6IkAJ5uWqWXRabnrZlR7iXAJjslJ8VJzSbOvYm
rNknXsQKfebDaT1iefkZ0I0Z762iOiWvIR0eap12f4JcJvz9RAzeBAaW4ZyAkczx3IYLwFNzh/0g
2pHrl6Pls+OFuVt68hp3jwzH7c003L035HPpddZ6HFBcZ3MJeQ/LoNxx+FWSqyEG8xTwd196QL6n
uNyNqC2ytbe6mU9D/s5w5KpomKyiSs16Q1gq8Rj3swuI/cDlyu2A84YTnDD1OVt7+ooOZIymcF7C
BaBzVPlYihS6ibZatAmcUNJ2pZYltRbTtDOOXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S9smd62+t/cc6T+Az0vn0kXxFJK9ox1swzdVaJK3ag284vMfjrlnVswyLQNkD6M2BaUNuZuzevou
xaHfzJcTFt8YvMUaEn6TameCIs5/mTCxVsde0MlJlF2crCf3fZHzWj5ooeKnlSFJXuUK/R6CGS8a
2vO0yBw4ZENNd3h5OqE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cOFUj+LOfMo1PTF/10pikQPB0v1eZ+hPEU+cjnPIX80Jf3IXfuV5X+QqrEh3UZH/0+YwNN5uc8yz
3GcUBcrBnY3TVkMqnhGUk3sy243Fxp5BXFf4yGZm4BbuFXxSAKu5Q+k+UOvWrFZfWdNI4lYLdSEu
b+Pg0ebBc04YBsQL8j7TFN2y60Hw4npf4Ha1Oh0Q36x952OAGQt/kpvEYJz+iBAv7Wj4b3IJAFhe
Hz1SVdnrXpsS0DFFqDApZsueRszhz8yuOSjC5Se+b7SzsP1onkP7OL41tcS1dxgV6XpqQDe6m87o
cIvrt9MVp/aWXYppakvqJEuPRZUIN54B2pTOpA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
yFcu3d8R8qI2bGKGFEP4X3dpsfj9YpgroFBH0sRUGmYLcMI6RS/tpYFFg5+2bWSz6rjbdiWCpm9f
ISim6hxeI5YvpWZutiWYsYxGMMtWtmW1dhCE1158wHQYvGlUyo5TFP5te7KfMs3b35qTe3MrBGLz
Dcegy5oIG7p5nGDTo7685fXoqlZKzE+niORj5ffukBh2Y0Dw2H/kfMFhzl6xhZFOrQzkFB4lkn7J
hDO0+YDZwHDnKfV6SMx/AU0FHROZhNtKFNSgs1OOmXC5My8fLIHIMvpJKz74OEERmhnVCl4nr9jw
jbChUJgcuAj3CUVRjYIbB54d0IUUfmPR9lsJ89x9Okh4hFLDnlOYLwE3ayWtCdDh2cBL09tD1bSO
1LXqLULMVX0k83TRK/n01O7fszTg08QqyOgPX5jy0Zj4JU6CcglPG37VI7RGFwczPz16h2CkfGZc
s67G43TF6HkZTMKuZO7IFU9goxC/c1DUoPS2nCzISMFOW1VwG8H3c3ftKzb7t7RQYmMTx5Vt9ntx
W3ouSQPKQ3e/N5gB9UH47BfuRHvQzusPTbpau+MQySdRKEpVtPvNpYoHwl6tC15ei60h8e4wkx2o
Wv+/j3oivHBN3UcZlcFqCgsFgg+VEzr4I8ddQ1UriIXN0LhJgHCjEetpU6GSvoB8ho0/RyWcQRev
GW3+mkiGSDwEJhki0rFjwzhrglESGScHaFgczrX+2uY0sXQBnEczrCqylCCBavlAcZSz3nXbtJrW
YjGnz6M/KkaW0YRIZkGuY3eLlDU8BVOhaE22Mcwv/7vvrt7MWpC39fUrN7g8WXTIwPpYo+EBA76q
0Ei+Jf0UalPCZWljwB4MTk7KjKoPQL585IHoH4LagYXShdtxsnzI+Ze9ZtFkcq3APIyVfp6c8H5X
5t2n4MvVHbzd0Wb38Ane5kNZ7DavvaAjLw79itP9//m79pNm5xAm0lDG23YX1Vr03c6ttKNXfCGr
GDkjieBGVtsDczTPmxjVxjBrRAJ8ju8gQxbxPc/H3tCwQRQfttjPTuRmqRAHsdJw4Ub08W5iSzeC
RXoGuOmoveXmTsTVLgxSkyv11fLPAISYtURE63xJ5MXx8WhOlfbfQ+9o3EhqxQb25ciIgHMHYy/7
2C6fBC27dLa4tU806X9xBCJUOxrAgJyJ6TXt19n/OXMVvNcRNpzjlJo+ugm+HE87J0mKNMLMzf8k
E0s7g90ZCePO89Rh7WbV3BY68jRoAGvs6mB7e9tMyGRhj4Iadef+ilrXHjumPqw18HXNCigul82e
MoyyJEwdXyZEVm8E5mt+a8HedN5fof+v2repfC8RGi90qZcsLuSpXuHq2DP3VQhxB7MnZWRsqggA
TkVN9POkuF8wPBobobSTb4J0N322YlbufSwpQlu4I6zFVo6sAqCO8+oIn68HajKXjRaJ49jMZhe3
Ojnk977XmxW6Z9S8ggDHMlAnCMP2WsVWJyqJ5OQA03jVdc+rjXsPC7PCSww9B8SyVhDtX8BIUjC6
iEaG5QdOK5syaSTCA7HGCO16abX2K4a26PXkefCj0WjB2bnlUUESp7zS61AL3IuBanbzISFLVjCm
W3YMF36DtRvDaPKoD9q/TEgjVZws1uGM3uDFjijCQuUj6Q7Dypb2C4Oa2xBJRfKXbGfCV+BbXz3b
ps7Mvdc2bJ1xjqQv6l+7wUZ7f/4YT2PZeTrpQ0plN5JOM4+DipsELxnY6sccfWFLMlHQfxLavTY0
956uvRtbDqg5kmPC0A3eX/Cilbivz8ynJlYXvxP2ax56PDUkNJgXJv0RDrQpAjrJ5ICuxT6COm76
yu/us6IwvSIFIaqGad/pYUVIihDBOjOkscgi5UZnl19/dV38YCvJy9t+cvw5n2fHP/hpgkRCdQVp
JkqJF/1lobaWfydemuW7cTBy+6ckZr1dJPBGeGbDfbWXf3YDFegbMvR8+/kIM+IPTpnTX5Nwt55W
WbDuYnI8t68xDi2VLGEYgX6c2FpdotqR3/XR3VwN4Wf4PuRRpeEK4MV1PqFkXkf2BGnPIuTYNZZW
aw60SEJfY4M5MORi66i7CZygprX9JuQVVuOkm3g7MVhgugqO4DbucD2Kc5/XHKfMh49DOS1Ihp5k
HvROUMG8nO6zRx2LmfHf9bLP8qPHAPtVAvi/03PD29bGIwRmiVtbbgyGVhlzSIp00hBJ1ipjNl1n
fOwomqKVwt68ksAITtxGSdBcEm5i9kT+uesQSf/Fdgd3v4x4jXTZ16J/p1/i1NzNPU7cWcinpbTS
i0XJySXOpNBB0dMyd28yy1g/IEiybQE2vdK8SbLPzna7NAl2/TdBDJgAsSpxyjOplURu2w1jXYGj
1+V0ksRAVVd0sxuzHmGLK0otw/c5VOgg2pwwZ61C7K37TNHl0GW5xyt+7zhL5xIKjlbYzmj7isew
CURJIEvmr0oa8L5qStmVLeQbO5RAIeayic/r2iB2FOhbcLYyvAUSKymEorx7XNLxbxRBHV16KH1Z
sH5Nkd/sUl58Ceug/AiUbPu9ifd2Vru509mG/Z64HZgH9JvgBkBIngeeU2Ak9IwwqH6iGgp83rmL
hI3Yz+9p9VSBD4Q+dCFGPR1fMZciwwEA9V+D0p5M2wEnLDdwMWhkUBfqM9SvLrOi62cOjtsYa2Y8
7HEbnIEoOyebYMB+gkL9zPhuSyAAA4W1xK2Fy5mJcW1krtjqXjm1IL49In/GEqh2LWt5a0PVZu1y
cPXgzekeFZAHb/B2/9A7+aqIihXT+ELOx+mAiK/Htwp/RmK4u45xGajWzAHSX0zehUTunwdfYiHS
tcptw7XKwajj9Qhw2mepi3b/1d4RlLSxteGSI5HbZixaYpB0wRwJi3Ihh1GW6YswYc2+DM9PacPO
ALm2Aw8Xy/nWTdLXG9V/0byOf9iPZxckkzmzF0Kes3TzgMy+Ad3WiMwcMJTRVmIvABqLjd5DsAe6
uB/ixW3+zbOrJdSfZCQODyfmmpddOo2B3KEPDKK6ecboPignPppZ1zWUAwp8LZ7SOLRf2xP3iuzp
N/9dNvKpebaNFL6J2Oy+XxnN1AeRQPl0JDZG4Z7v8PMVMy9SM6JCo6hFqRDsJARGWAb9h5HwzWWz
S+oPQoD+Drw1G5L6U+xDhem1Y9m6Oig5zke7B/A2448uPEQUicnwi7X8aZQDYdOn6o8rIhCDzoc6
oYt6zn/QEUNYiNmdn/u34Z8Fzmwal2ZuRpq/aBoOAFTlrHo3RotapfSJ0kzhviYp55m+xB/yGO7G
quH0pB3rZWTGBuSjyXioyNZT9W4n/CQcopsy8StCOuBZObj2ZOeD0HgAy7Fayof19oYz6IGcu3X7
p0+4PmITEmKutyGqUBpLovmSpZEp0B9GJ/g/ivLH9cRPa/uCdVCmvYYKhJsZwZGzXpuheC7L3BEF
iHFv6hJJcjimVDW/i9qOrhMCi2viHIvDzKH6plpxfQ8fFdSLMZG4gywP0L3oehhUyXeLYwVqSBj2
r60HFItSlPbTxuJj+2GD6bb81iXtKYEOF7rFV3YU+xv52V5es9RyhLeYr1aVKsbxFNbDjCJMvpDG
HTCJouI2rHNNLdASvkx4JRfaM3FdqfNc0D1m/b33KGa9DZrj2jsOZsyLiYOVNSuoSZxG/p4XEXxh
n/Lk+MU0xDCMLAn2jGBVGTLIlSrTGSvG1/IAEYdS8O8BccsPuaiEYaNl4BMh0BJouhWkkJAtgzsG
5VthWyZGOYyFVCGAuLy8n3HzSAurKTVi6Y5XhPty+4drDYE5gOUzrtXhlPXCixYXk+Ysfwlo7fHe
NcrV/PY1/yZIyCIvSm0fk3pQmPUCsEMgDNmAjgC+pqAax3pU8WmDp13F8kV/oC6uOx27hVtOU6XB
s4mP0t/lC2VAKFHIM6jHyn4KyzeVQZAnVVF8kvDzZIgjkMadKbAJj4ki7Ab/4tTlK1ue0LdIZaUi
Q2I8pec1dL3sEgKXnD3CensqG426sAHpopebvKb7x29rVQbaLIdioX81RZ4NW4YIrYuCgW/AUoeq
/XxOs+ReVyDOK7WQbBHrg2xmXgrr4q7I2h8vv6SbGwjvv6EJYVL94KO4ICQDzi296+sMvuAziW5y
+ULQ0Ln6y5nqFUkrBlwrjM+AmxdqcrZd4JFNzLaa5J3lPwbqG9NQfvZw22zoZTFGq9jRhJqa+sPC
dRN7NgCNrjuT0J45KLiaSc5HtZlopJ4lLFMJ34x5a+exrB/E4IRLpi4bbGMl3wrNIC4vKKQuB92I
KejxOYmVRMH330vyG0V3bOUqpyMGHEQiICxgFGfHIqR90hIygA2cLTH8fiFc8wVMG0EHlBIC+75l
r1UYn93ejpgnm6/5MEcswWioHs9qCrijfj2OtLISfT98Aq/ax4jHdl7REeLDfKOVZyEqkwOZvdZf
IH5k+Nm8RFxpb2wMkETva/9dKXiwD+IWC7gb6Bl4oksSrKP58P+ujETggBYXEx2h/URZ5KS0zaiz
DeBf0mfaMRlTcWIjMs5/94IavxCw2GrVhlhICoNywDVHiPEqSQ8ufwUO8KWjhECHn3NGALZup4j9
mIhS0sc2Hluc51r50BlROQlenCjLNpi/RrpkMKKKmG2L/3u9JZ5b1l5rlU7RWxtUqrQFZAkjDicK
Ng3YXLhM3v/RPBTec06RVGd7kQWSSnXcvUPQRloLxouJVYv/hA3+7NCKmsbaJ+fl9pxradA6WvNF
+A/1j9OyJ/Tuw5XHNH6BDzlktbbr3rtdvmKVXEqPKgYdlanhI3WMuuF3eK13FhZrRyuDaYrmc9jR
/UXKu2Qk5znnLnDBCfo6fJNgoWZ6oajnA3yJO7hf7RBc5TJQH9gvnOu3XqOUiT/B93SL2lKZap0L
sTMbRqDiVPvpS72iKleq71KQLwiZNOXCYf/nVSFjNnFkM+SlUx0EcJ8cXnZeC6LWf2/UlKUnM1Q3
tfa32/35qqDq1UXyejldcnraYvCPA42bso6geKqGboE75nzqMz46YZxx2iBlaE6Mhx6nGGSBPSSu
pe+JKmcVfOkr9gybJZG8smsxmNvS9v/TeA0QZ5UOVvGauxkFnyJsGye1+f8tnc85gXeKon3Wjaoi
OWsti1H1etwcggY9jXJ2bMzFv6AMnUvjJhvFTELCbyqGMlTedCDGLc39w/psVeCYs0ETNVsDFKv0
8oFLOw+CT9U6d17StbNhrGUyHJgYvjV6tOCSRoLKyI5Ahz2GDAXVg6sO9UGR9dUPwciVuoKaDOpG
5rps2kTPRqrOr1RptiPG+wQMclgZOLGOwK3l6nvpsA1caGqjbyHWlWBPAY+vXrY0TqFrkUFr/8r3
qbnrVnujJVSxJGomLUKUPOQGrbGYe0wDcO3vg7DhEHR4ILg6LurJycpCXDaiHcQDAnJXAqfUml3w
RAIpuMCtSqfGR7zLfm65o3k+tL+uVKwNvtieTJ7CKRgBRlUUX+gmrmfvnxju/89sfiEii5GtixVk
iYQC1hYJs2nmxxgwwPN3kFj4xYuhalGZHtSnzGMRvztxJGcKbjk15/p3GGxVYOdYTfYTmbYKInn3
toPnFj7fURc3PjhEWt55k2RBZE4hItLYVIecd5AtJT7wtCAW/6NMG+Z77awgCeIbdb+oDcrKO8/D
3MczR4kNT5DbKdo78Ak/HFC3WFRBdKCkjifrG+CIdb2A+fGyLiyu3tR+5DRuWuLAHxPI+EeoRx62
jYJjlNw2SAy05Zo2ivOhilWdyVoNuh6FFAp2nNQdOIpA9r2HcDG2vFpRvTXt4NOb3Dsciy2WDssk
f/fNqtNcTaNZuAQCTIDnFS1/4f8Bl3W5qvl2x0QxDNrdwowJe7tD9txR0zfHB/140nS+JWMeZH6t
jnM7BoEx7m2cpjyz9ejCC5FI7JcP1IDWEsw2GjN+6S1z0FbVK/qbs8x+pvqhrKPx8P40mNS7Zlhe
09eQ0Cko6/gg2L4lKYHBvDUv1rMFaUutLSgvVC4JaY5IEiOhKGlhTM0eTHXxfBTZfq6n4Q8933+m
Y4/i4x6DnVa4CBG6JVNK8fyT/EzeJVnidttYNmxZkQLzQoTlVcmnEVcAA0ISeeYmi0BetHfAfLCp
oZtbjMk3kFn08GYgSurGXBbf7n4V2DmAtsbpnbNnDi+89hi4UgImGg5EipelM/oPrr/CjiwSotlV
SD0MmqyvS6+QpdkFBUendyDZ9e0eQU8veo4LjCKCWM0bMRd4WGDYRCCjF6V4rsIYx8Q50WzQpum4
SplepDWl9RjB9XkEoHP7OGiGidxMDUGL+Ccdu9NhS8M0PltI97JaNXRpbcEOJaL/m0lHroehCtdm
PF8QWDNw2TUoyzA1+DAXj0qnmVwB4NNtZEsG4wPwLCJlK/PIY+hVbJFPOCAu0uWaUtCiOOL54JkE
PXlFJw8nHzJD1pnwelSm1NdQFx0KA69oKAGS6xqhwB8ew4crcIbZe8aVsDLFDm7wtm64B2TNupkY
q2mxBJueMOIzTJfK+6pFhLH4xDj5EnYoNvJ5ghUoN3jVUaE1a38zq1lP8JMdQLzrhAhPBkdqEnUp
jPqIcUpChHxlXuwngaQCuuy+HCsd4BnAlGcCLmRKHHuPvUF/E8FPisfiNu7zBZ5dV2fu2J/qcvC3
EOx8na1QkYcdzkKJdXcS99dZ/JGUTZm5hFb7dmkC9giH3wU/lWQhfeXkxGcF7nqqVb38hcvYUY4p
se6tMzeoKuV3I/Sm/Y4/EaPvQA5V1Gr9VkdvxhnC3u7vK3oMeVJIhvvudfOppCQXmKyF8XNTCHqY
/MRgvgbswmrvHjhI3ALhujvRQDocl6ZxLG/a8HBKcSoGu2PGc6JPsqALXABylC+REoyK1uLEKX2k
XzvjQJNqg2q6RcqLdiKCJmU3/wKf0wmB7E9+h3Zdou0krk1WBfMDluUCKLHb//vyDPIr5dxf0onE
qMaM4vdm+HId42Y4cNY89T/Oufsi8kvMaTpLHbHgkclpH5yY9oAIImBeyYOxPqZexMlpzG/02P9l
EW6c8Z0WFRER9uXwcvlvlhG9qMVwgTW8zoGY1xJMp3Y1CxHt1YU4+igc9mJO2MjRRzI8q8OWfrwe
49BXNYNJfPHsCpcoEIixRgSxmbN+2EJsmm9tnVJmxttOl3FbEWVEO78X6HlE+BzuJ1OQilcna360
OV0b2JJPRDZlGBWSfAWXMyGcjolT3sC/Xa1v0ikUmCv0plXRKfrj9iLnsg+dpeEyHcUFNfAsvMiR
28ThlUbOxCBf8dhbqvKCzHyfFJcqUwgDk7f4LStOaoL81RlPatavsFYZASyCMPafqJnJBE0LQsYn
ecsDDPsk5sIrjf5Swu7G1TEO0RPMH40bZ0249gRedG0YlK9on0/xakYVHg57KkLbFsb3dHXGkIv8
Tfa5HoxB6zIWZaFmzzoWTrS5ZMCjpMUJOr6p9Iik+gHLJN9LaKmgRbwY1SIy4OEggFSIo1HOLpZC
tNjq5ib4g8ojEICeOXQblBcacdk2bxbYovvuNgMHIWytccFTDy/Tjh68lRn9r9C7G/AanxrypAhD
L+Xf5odr56vmiSqsdRw8ngPL1AeWu1+rohFBewI5KINRp/wUQ3hepyDRmW0VcsALOfgK9to03pb/
KlKzUpXsHJrpa9A/cZDL2gu/QgnnLpIZWAx4EnqjKQmsu7cukyFbWsa23H5J1lY/IsrHv1LClwmZ
JERzlvvkPmjp4Iswwi9a7g8kC9Ndaz1dc4toa7Rsncv7WaOKsRMAPIAOqWrtLFjr7jOpA5B/nUyj
eO4DJ5UDJExBEQfCW5ZiY5e1Q3m/rdCJ6tjob/rudLUU4wG1Xog08VZR14q1n5YsLO0LTiWDHjNL
8tWYs6SeGt5JbXhown6U0wozloYdi8Hu49MT96fFgt/lwiwpj8A20oe4CnTy/TAIUHY59d5CIlc0
FR8Ts2kiJa+26vJ5F0xTPnCwc70++DgMjnbXz4/6XSmYEp1DjUp5+yhg8VBO/zL1Lk+6a5IeiRHV
pn+bjo/MGrwlD14KskKHINGIA+Hy4u5oHdPbxk3L+jQ+g58eGnXL2El1ZO6r+1lpgH4Akd01cWNq
RoSiHEM0ar350E2l0s1WeEgrETw3fcypv25quP2BKNxsY17GZctDD+C84bmrHStK/wb7+aweTZOI
XqG+6pPn4MGw/BX1/Cg694FxBZVWG5zOyVgEjzg5O57Ysw8OakBLBUtXXarfRDrXd0jRhfeeAmrN
HkjV5CJijy65OySN5DBxqg2LwynFDDRgFepEmMyvalIaXFu0nfmiHD6yD5F37YxtuethQzYD94Bp
redA3mr0Kx6rmVd7C5Wx/zZetLKK69eCuPajl7joY+aiJYRJcC3LOTP5rQ==
`protect end_protected

