

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Pb7E+qNVEP4sE5d3TkwQJMYKTR/FjAPrexB6qdDJcLdscPV5w27UvNCqw/kg86JgS2hNrfoEvTNF
uJ9eNTpy4Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Egq1eCtVuCp02bpffloqFi7UMw6fphk3UOZCcejhe9NQNeC0Z0b1+S1NY8yEfAVY74l4oz8pZ1vA
hbrAzplanZae/BDY57rCQ6UjD8G9keaOwYv6mG13f+m77D7Y1nVpXOE4Uujw3cZ1QgwXR1H4YfYp
ysjb+lxmo0pqYRikRIQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KJqrZ5TKkbTlecBRrKRCsxKhAd1omWJvIin7DNafgTE5a5N2or7GsTSawdWWjYWHESLBvStvRGQE
jVUeK8m63dYVJN98fa8T9iAHTDt9yiBRki/VqfvAejvDOEI+l8row+LhhHMvCd29xmkCeQKiq4Qt
hsdsz+jNufnCYY4Y1CVO/4preMZeG5Ow85vRd/341CoWEOBji8o4pk0XyIttBBgjBzWO8JyhLpza
R+Z8LgFoZ5OTfgpyTJ4SjYRWp9IHP2HL9TShNo3PmM36nFNBvQSLoEjLgk4+rUr657++ugJH31/C
Y/QScvwJcbqMK15awb6twj42y2gxJSFzAPzSGg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KxmYEF19quU2lnDIx1hLVbiBV1iU7MlwBSbpQKNAVv6HLtZNpIjv2UPtz6sPs9Xac0T26s1Kjo2c
fAw+uaSeKdgWE1BMMV8ya3nIO40+wJlyaPYGp3qW9dt6kM+FZZl/3MCpgIMx24FXg4CPHrHNKu54
/3DZJ7o9x/QjyM8WSeM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n4InNydlMoO1IH7Kq1VdB5tuRxM6d++erhleefbfKU7rQGdfSjRtqcQ+h67LKfA/jQJYdDdZMjd3
Jp84+E2i9v4ovZP9CPOifgPGXKRtOz0XzimXarAjLF+OJp3As1WqoTrPJI1DspdbqtDWx5caLezn
hcZVfRSFpZUoLc9H0HW6DXtxAWvJT8e4ntjJYO6koEzzHlZPpMhXvbbH/rbArm4iRGWLOVN205Pq
oJcFHv1n/e24XGuCRksBqssUXd+D0UgsxKn8Hy5kQi4Q8xdFEXxEOVBI7ivvG+HKnJFOOr+UNhLY
+rNFOKSwlDtT8tPfpzjKS5GdaTuv7j2GVoF5Tw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21824)
`protect data_block
VU8sa0HJv5QiqDbFjOukrxTGkD1oKBx8PWc0hvnPQxcL8GWt+EqYRCUjgSS+gpeFkhkT9RzQfRzh
w74LksNHPfkMOKQrRMr/QHwxsILtM4a1o6xDEnJM0XjgDRH6HI2uJsJEqyU/VimHgqZJmSKOmJQE
AhI4NhQ0E5/j9TN8Ms8N2+U9ri51Gtk2IYB3BIKs8Cy5fkqKfJnXl4huC8tQekKcYtV6IceReRKR
Sb7PbKQDGXp9YMk8jmibQ0ryMiccWr82gUO6z32IR0hcc2kt9iu1hFGD/Z4vSu4a1M2Bh/ITUBGu
uy+EeDwO2ZcbtDUifeAriTZQN+fHqBL4jLJSZA1RkSIrOj5hqEXZ8AuXob6SvIDlyiMwjhlXKAlT
POHJ7qjvdaCcX4yUu3X8OWu5iddN4OmSZPlOAy3Dtktf+Y78GyCj57Ij8+aBHxW8ywiUItEWxHTn
esiwL4HKaBqcbUXFGShLNrzmnA4rVYanRlxJnKtozNy5cirYe6SIvNTCwWry1oGIXZnlYWlM2FMb
6DFpnDkTSQqMz8gxxuZefzSXjmGQ3LMBX2/IBpbTdyj4xyuLrMM6sCZnsZd0htnnYbBHrqdDwkCZ
sptrwfBm5DK9QNQ6wKJtKMlN4tAGdrtWtPRXd1CUmfxFmnsmuRkRB113dKO9lXuEI4zFv2dmjPIS
V0robbF4uTfW0dRN/G16LSU+RvMVFRVezlTUiFFL2bQAr8zLdz3y2AVoy/tZnZu6fv4E8aB/Kj/o
h68JaRUIpXr0U8AQ/x5YqQzsziPseyl8KoZx6Nek6rU1F3KpoS4k2UbZO8gEcN9fmK22ksoD4IXd
D99h4fv40dp6jxx+E5+cIe//Ngb8wH3z4JyLormfgzX4nRHTZhvdyBxCxQFeO39AdbW7RO1VKEyK
dyr6k1zO05uShlz7xWVcyhFE7nISovpl3Z7mO0nEITmsmELn9npN2XIfsgkLxC5U1glt0FjTWa8e
+rvX/OpYjrC78MDDEYFPts9aIASEn2V81abcy6nwFbDOMF8mpRwocRl+Qv4mi+7/MBypi5+sN7Ai
pSuN9g2wB1FwJjINCQOV3FG0uI0gPg7gRZfbOcMbdnUUm8PzA45Ib90z0Inp8TDFaPS8gim30RrI
kEQNf5Q0PWuVgLo4TgXRwEUowgC9+/8kT/IneTPprQMLNPmanw+zX/s5sckxn/8Kjyxvm5gMnNFg
SpPC9jC9gUK7bwuv6vNSsiEVsuWn1e6tt466rv8I3L7lZAFSpSM35Mm6KljZWdeyABNDNSRe4JB0
WYAOajn7c8VGf/Kw9xO5EwF8dw3q2FNP7N+0r3YeJnC0YK9237m6EugKuhhU0wZ1unVFCsOws5qZ
dx+l9Xpc6Eoqs15pfHJ9gsuDBNhJ6tNBvIrg0PJ4u0orCqTf3dRuRAiciqdD1hkuAuSOjNprFtS9
MB80JoWb8kgiggKEUsKJ84byKP5DnXyaaWGNgBuAhIgcmOVa+zAafy8CndQVqwDi45RXvi4/spR5
rzyn7O2E/wmSlNZmZ/w79YgzNpxQKeNewq9WEkqb01C4fTCgs36dZuffKBrYjkVBz6vDHGDyKFQm
IQhEzcEvmNewr/SyrJiiP2UBV1cC1jEDB2BPxEgfMkJ+jsamTkRsy02uIRXSAFsfGmWeXKK7nQ53
PR2Usl9pi13yy83UOSaHNxXYAi4Ka8iBKEn+fNM4hQVBem32JG2EqwDElXaFun1XgWR/kjUl86RD
tdEGDbQpghmAp2d22CpUQKXIsA63mlRwGknhlbSkqHwraGOdvFyp7nhfHiHj4UA9cSZjoSyJ+gz+
RDQul5kQpXvptO/kPL4ppq5P1Slja9R4bt2j5IFlGGsf+k62RYjneSslVK1mii0iqz1kWYeXz/BX
lezwLoxXzeW3ye/t/+z4Ic2cjNsfclEcpLCHgrRASij/aHjUsgS5Rjsz7GAv7SFQENHg9NcnyZKV
3iZP+DESyGFRD5U/wNISRVGOQA0Y+0khavxjA+fuZanMp5JkZ+J+HPNyB9R81bhOva5m8EN1wlpl
+dzahOF208dJaWmEb85YXbJHENyYEbTyY8o/rYR7iGvxs44nrcCs0vyD1BSvvgQuLqsQsgezdeEp
mSJvCOVX4wuGnjL7BwTCMd/6etOxkGKA1wjVarnu9uDsBV9puLlBeeSXc7MQF1NnUGqoOYgNvDDj
8RkTsAMfV4YiKu+7kKXAJL4ynebWRqry3xPtqG4v2YREsAQmhV+KpYItKmhSpw++VXqN6DljIwmp
yFfSEgnMNmFEb2js4IMqiFYzLa3jrEClFH2k9CxS/nQaq97da2LbBXdU6fBTtnZE6vfvui0KGgz6
dgczVi5fy7gMPBelVbot29/X66F+KfUsNDq88izTIZGlh6aWRt39CiKSsIh27pRV+MY6tlLOHWIA
QFj3Srh+UdmB5aA0/e0YekGMmPl0NMCU4ck5bkaOS2UNeTCyhs9OPYwLHwXP5lNsziR3X0YKPoW0
+K5TG0g2kPQpZy0ge8NgViJ20tje/K8tamkWQat0j7+G+cJRrnq9XhN95qx1Tp/rkbHr0v45dOzz
PBAcPoNZ//VyWff3NXxteyG7NowOHguS9Vbp616P0gxOqdtRG46bz7Bxv5Psdz5mjI9PaaCCg5+u
gGLcnGeH32TNIdZFEyDQoqQ1YQDk0EMtPxOB/T0f1ZtLloMEv+LEpjpa6kmPstdjSaKazhpLD0n8
noBAYfexqMV+lOF/NU97sUAE5+edvJKYbjswtYpkj3jaLxLAj4vXEvaqVkPfCnGK3Dkuz6TTUEPs
+M45c8jLaE8wUkwzI82A/8/N7SArPoaFP2uiEooB42KS9d14YiCk+s0qdLJB0VOveON4BKp7hBAr
N+GkyEhe18XKkdLAG4s+MH+Nqzku9dmdD9iVSMc3it4px57TP5AsBqn18DQYG9V276jd45RontPx
b9G6IohiceNgG4X9rJhTKVoeDDqX0ujCJ+U/kac5GRCprbI1OcBWJ/ZiQ7JO0SpGqm2hc6Yu2lK9
Lil4d0QeMDipoQXQ3BQBIag0HJ/O0Aee7vLOu41H28iwqLkQ3i3n3RbAJ72jLar0k3ZCdbuJk+Rr
4/gkHXyvnRbYY1UkZZFMpeKRHoZInYaDA2II7c1JijaVPB+BMtS7E04bg+qsdfj9V5Q/OaN3V5GK
OkgLuOWHfhAu8wp9eOnZUkumO7nY6s23gHKhEV/zek+8Usapt+w9KAAEkmfF6u4wdvxI83sXebbF
gRgjJjzhZ6Y51Oyp8r0PwjPB3PUhmvYHLSsVOflKURAEHnMScBx47NJXISC4dF9Q+xU/cALqQ5Ig
NTP+pZLLIGkdCfNq+n/R/1FAKSfrnHPr7m9qrfrsea2nYsKp76Vc0XP/QX16NzdpoZP+yqJo7E0Y
Si6UqpjmN3hKcY6Q7ArAGeL8PX6vSENBU5EsLQRtCD/MKFJ0G/Y+tAc4Wz0PaVpchIBWfRrim0Z9
L8Vml2cqr2LhQvLal2P9ErxcliZq6YlnVjrw4G18gq+TuxxLcUcaIjgizcI6f4nhw6FFo7vDzZS4
QLBK1i5w2Cnt6n6h9vusxJ+rB0mIVRvFUXnf5XFFciSLdTlzQQPubOUZEUa4E8dlkUhsArZ8CYov
nGOU7n/oegi+sOTd2gAYdiTZi06Of+2SYgG5lTkWYtFtm3A5wVK7PhWFUu4+jaGHwBwCfAEJy7cn
HejG4DfoxhiW/KGVdFe64jpQ0sgpWSlYfs3SdadJQsjB/mlhYg9Rt6fEnO3YgrtjV0P0hfBwyr4d
wBqgAKWQ5XZ8k5g1F7LZO8wOhVSbnfKvCvr521DydlFUcSWAYm+Pp+qk4je+IQw6HQ0Eq5X8RaBm
5asCvNMeJ2rc942qoQV3rEmcB3ScXGml31OQhcdm21aH7+XS2OZnhvo9D8PKNPamT/HBNiYNdidD
uodp3022IAwQeRUbu44kJEQTqh0pQkxArzdgh20LY1lIzJ0iXsviXbmjUMAMHDuXlzTvSPgadvmn
iLtmoYEX8B4preI1age2knIRWluW33EXIbk/6WCFJDb8Td0FhhR9P5zSaunDVfDm/8e526bZP0yW
b3qhI9lzRGJsOxZWdygIx2AHh/kpptHAe0nnPG6YICwaMH/rkV6sV3RO3IbXJtXWXZ0mhP1+NXzg
+PodLwibGb+ImfPJHHbBB0ZWctYQDjN5tA+s5MTGiSW/ABTdMgd6x/DNl2Ngy+avHc3CihyNko1f
QNVq25F85wU48nTjDmLJqT/WUgAFEj8F4UpId8bPYJ1NqXMm75cbnK74aniXVl0HxQqi8cJsk8tn
ml3jRV26tgpMX4mL42ggI+sCSwQmF5y4K4lSC/wsLS5MvEjb68dW6ifdmyt+JTWDiVQLwmpBx29F
R/Dbu88z8CMyO12r9N8kxkxE5kg84ePqGs/fakoLKvFSotX9AhUPSgYZfGbut+FW9LReOq9Y+Drq
oHR2sSHqdppsttq95slK5AA7/1Av1JhQFqvz8zqTZYWxby/8pHNsHndZbNUUxV1sjiCCX2hEfUnu
qNsYOE44y1c7TIYDdJr05LV+h9GvxXnLEuUQyrhYhmOEJjwqerG4DEM2uIb+bvH+9HgyXpPNTKRv
GNIQ8Kr3kE0zpabk30g5DPu5eCh9NPw56SvG2GsTt7wVz/3pkS5CjDS6eoEUP9BRNUokOtlaOtp/
Om4dyUekvCHkvAeGjCw0GEmqNT/H6ekWzifXLLT0Cul8g4fZKMC0iIbt+ZQO6jk4Y0DRLqS9Gc4o
3Lg8G9x7wO1MNipyUSzLNx02b0cOCs2dkXTBJ8NdrxBW3XV3BGPct9GH8stHDT1yGYnh4LVsgAtC
qbEQdYvAmDBLiPOL/SEzygTvcGdaD5L7LCREdGbc8M32hznFVaqTCUOvnmbklj6tTloOMYU8thUs
HAIDT8a99R9VXh245/EF6fZLhgUKM+Y8T0moXqwishfwm9DQ0YDWbghGfrefPAcovemiFMh+IlX/
wdff2ysklviqdx30tLk2Mi2y59cIyCkkpJ4h54noh3KywYkHAkaWW6Q6lC1Msl0blun27wsGgxxF
gKqE4XitfRV7y7pF5fqmjxEX9AVRSr7/h4F1fk526fxjHQTXPMxi8M74AoRzIfYNWTG6BwRieYHR
r13pOyh1SVYOggYi6uzsY2FMkiwBpdQTJk+hykVZREf0AtPt87M0SdxpA+TYgoqRdHEKEZpJ6suS
fLS1BtUVhv6bQFUpBtSuTdwDvjq+0eE2xBvheEYq2BXrwF9cHyqcxPocuiLGJ++0WXO7PzlcHil5
G6P4/ZKaXIr0hJX6O8jaWFJZxiWPOhBzTrcjQn7dfzao2BFYdx75qfw+2aIq5Djonpqz83EAZJPQ
YGfEY+rJPPVmL0kOpjHiqI2RCX4hohrCbQaYlfx4i6dzkzi1gIukiBkhsZ+FzEdE+zBwALrUVsmj
phRUehy9bkiQOcdx27WfA/FfJS2CbX/vFpJnCTmxOYRF0xYw3VU59NXkkKGOEabPJz6t/6gPEWhm
/ON10gkyZ7btVVF/CneipFtvQdRjSmtf/5FDnQn0ADF/Cng12PTufluigAZbfM1q+g8U1i6FC+oD
dU4upJpayWX/DDhbL/2fvX4ZvVSIPNuzXMB/dwLCUDL0Q2rHyMtB7VbR2H0x3vs8kmyGb62OtBXK
xBkbgyn4Zhq4MNFvrST7EsivBJKY/Gru60j37egvruDaLNHejY8l4WsvEASjCv2ncz59K9IXnIuS
rOFq/S8LWLH+iX0dDY79QA+BgFl3vqO5b0b7dMRfcbeBZMDqHx1tVPceRyQSwq5R27qQErv0VMuh
Ls727gEouNk0b9oJjEppgQlk3hoa06GV/JVqz+Gump4/o3pDoFRYQS6hARHDX23b5imxdNTpxSJd
vSnqG5W0JjOM1mcRPkt1bTP2Z9y2cwDmoithPPzOR4FO+4rn35OCkmhI363tpjAL//kTPc6qgNW8
hE2lYYNLsw8C9bwyPzpvo8AKHNN48KvfVy3wBSdkqoV9EEPjuxRy14gv8XW4mxKandgwLfLR9DlG
BBdtsKSUqiHsWp28pEtcRautRWYvunzmmlyOHP9DQgqKf5lQ6zbCBTP9KrUWoe/gdxV+G93oSuNW
FzBCIMsyI93lWm53hJWq40qUI5yfMRCjJ7ksmf8r8bTuAdzdyNwodwg+VTkg4X/DwqXIuZvSz+np
HkfWjkmY/iC+2MGab7fxBMZV4QxOTxKL+p600dNS6w9oqzPMbDohO8zy3LdPN/Mjw2yLjZpSlQUa
Nk8g0ImvTCHQn7c/cA45+4j7fPwEt+whl7r0I+xgW4iPq2FsOwdtPsKnk0PMuT3hxB/906HjeShE
OQBNOLrZW4L4nZIDufTwi3svTolOGMtYTNitvS63hySDiCvK6Z24ZCrS3wMso0MoX1Ey3pPtWM27
1OvfdzV2bNil0hRTFUMFh0tsR9WgAVXQqQxJ0xRf4NN/ppPKa3hcRRljmq/WKzY9cxEDvAguMBAr
aI3T/gOI9zrdUBIb5FQwp5AOCB8iJ9qLRx4NyRYynlmoY2XCMSkXjBtAeArbfnIGavZIZN5qTOQt
du64nJYoh+YOxfohgTuB+yjAgiwpwOaJmxKdk+RkpDCHVAzebri0jk7JpdPOTXGwAtda/lb8wNGE
QSjAb/HeU77IpNJl4d6enJw8kgpSXNondl/Ro3kZAyH+VIYKbDJa93w+PylW6HD+iE0MX9VDSLpi
aohcwv5XyRISH8NO6uBLYIIJGGqBFTvLBS+i4n+BVyF6TjJ6ccFcm8J4LUhXW/jSkH/uo1yN5o+I
oavP8Ik6XGoQ7cicsYA3wMtX6ZST0sHZRgaF20nEoE/53JhL9g86IyVJIrQA0IdosWjVtqTcpzpx
HOsUQVci8i5+ZmYYJAQweK6WLuNAcJ97lGF/lTEXzTPgx4cU99/IqEfAHefakK79kBYGTXsGwKqo
5VfwiZMfCOXEmArWbzvozeIjn1/7KKzSJ/CCdqV8YEXAKj+KZ7XGrrQ7qURd9GrHP3gWdmgq5k/6
v/wEhsOCVfBeJ6BwwuYEiK5LFggoxqlcsWfCBRIOgSPqc7LsLZtrmQlOptc1PZLdFXCE5k2flz2r
RWo99OtMCwE2KzroZ+Sku42zB7o5kZxoYGlzxIumQAs8hi/XdR0bYj3wdh1trJJ7868XhF2HYaLA
kxddmiaJaKXbEbWDaYQ0q5UcGpflFMSzxm+708yZB7pvVwr54Wjg37b5gwFRyhh81aXdO+bIpZpF
yKOSYBW5dYCrahWy1Psgix6mar1DgVqgV22cszXGMtVVeCdByevxszNz1x9woDgNzC8AyeFrUn/M
emu1lYruqfSgLjrI0yVu1dBPouGCzOFeD4ATZGI/0Duw0UjUK+56n7V0h5vClk8pTY2Ji5HoaA0i
XjwG63t57nnmhM0wn3a5nEFKip3knV62Tt9fA0MnyrmPfYxyatNdsUnIf1Il1J+TEdptR5JI5DwI
tox51gKc30QOiB4CVWfaa3JB4wQKMis38t0hOsl3jXlWk5Brrxwna2KTxTqshLjuGJ5J90709C7w
GXQoJ9GtCoEeNRr3W4Y+GwTgQ6g+6J87x8wd4WCXOA8G7x7Bw0Z73KP+nuxRzt785Fn4cbxP9vdO
gLQQtS/xSq24NfDz+dlVBW5SByqx8VWPqjgojuSDaGY8OllND4Hnm40pbKljh7QYn12qVJ6ISevS
0aK/rVdKQjBlE/+k49/9wZAWpXnMGJawGWRmvbWFTDQaS5XRwfZHUzc3XJnLWrW539aPrPMndeBa
nbZEnmyr9nKoKK/lmxHikQXN9jl1gmo50dtb2DKmTns6gepxIYz8dQqjJzJbQPuCZ4LPKTtjQANT
utBUva3ijNfhlHdgZgmfrlMpfOLYh79LLjvs36KwsaK4Zq9a6VxR27zrH7kd2ZtIm07O6k6Q6skM
5zr+NX09zTzXnQNnEI0yzgUDvQgeaJhJreBJZvZ3JHPZJZSUcOAucrq8TT92+MCkUsLqnw5WRD6T
rC+Y5k1jmmQcFTbQFJvDCXfp0Cfult/VYViclDmMRqSAv//VDF90nT2fx3l1Sx6VOkLRP0Zv+zQd
URDTLYOIQJl1TdENkX/EIMPHX/5yUmvlYsQyUqMoEelywfnIgcgbZ6dpCDTNL05aI/GDQWFQAFir
9grD8k/vmu2cdZ1MApORmhO4VQUj8jp5minaurNN1rCQQlJkHOmx2neKptqpH9AHP2ALPE5leWbV
pyloIs4Zqin22Pqh3auLYf/JucnVBPNrXiiVYK7UXr9HViALFkAJqfwfDmhuzAStpi+RIlQG8jb5
Gpw/rkVuJ8sJ2gr5MkcyT3iyEN3ppXCpexL6TJi9j/Y6FUFIhWG2FttGjZHJFyIbuUMsjGbMQy2M
LQEEVtMvZqYaIhl2bLQZTm62fGVM/ci+2DdTPzlPT8uqyZkXK3n6B1grcld7XSe65BOXNepk5m03
4U+JUxiVkbNJEoQMMSVh3OgnFWcodSNHQdgz91qh7b0ySwmYBfd6YO/n7txIujbSZMvqoar4dadT
oiO/d5Fm+AQLsrX9cLjNHXb358wBwEzzO3wsv3ByZpyoIZjFcDSUvmvkgvPPbZ3p4nR3XnsGpAnn
978h3/Nf6vmASGOCI1OFNnnD2dSdV0MSTIE/iEINO2qtUH383LGEGoc6Uh/wsQ69gID4CPqzEefz
BBoZQev46PYD6C3L8fO1R3KRms0CPC2nPjfyLGjoHDdMA3unOT05vVH+EhpgGNNXik44wkE/erCe
+zLWbR/IfWeDvjy6mKorQq495rS7LHw5TLd6UOismVHAbNbimt++yTuhv6WqNg3IAUoX0p25vmYJ
s3LePiSHvpIWVf0TRNtBFrDEi4UTdrAfp+H0AQFF9udZ+RiWoNx/BPqhEHxgZdyqYNk2pm/Gm6tG
oRSe4xrcYUKvj7JOcP1QLvr9XeufXy+Uq4x1gNZTtOXMW6yw0Xs7LvJf4+bUc+YW371ZIg+Dk81Z
4QLVFAQqKvGWbAlGQTR5xcNrSoFGYMYkCSwQyU2LecgciiR6HqoEOQW4mNWQruQjBb/x2Bwgt5jw
zXEbY+C7ATQEebsHweutwalLwogC4mrt9cu3BWRebvzlfq/2zUeuTWJAvNOJRFxxsZg61ze4YxX3
rNL/V5Ru/0NBlp8EXO18SAYBwjEyk2R23P5gacymetvBr1zzpG6bm1CKj+F0F3VeM26KjtpTR9Cq
KEhum1UdPYxjiv+7JJWy9yw2/yBNUmulCj3wFSTvgdOJyQTUwBVar7kmatVq8OkHM753B7eijUnr
Y9lVUcKQbELxxQlIOm77EMk33zFpbAp1PlQ+GHF9fiijwe4LASIYhj5qmxvlNI9QGA2Rj3d641I1
4FRlNVTvzrNNfaA5na+OMAHswukkbrTr0xsgYUW12VVUlPxXhPO/9cgLL5jcG1DdYjr4FO1czvQa
Ydagd04cymgWbUCkuTCi3mG59/qfYho/NlVjObeAyNH+6alVtOFqHEAPUiMcOxyw84dJLEwJvwWK
pj2l/YiExCZwb0G+s1f+tYuf2udxX4i9XtqGLFJ/XyRb4U4Ikrdh4j/vNqnWUtx6iUJiEJ/Anvi8
6J43TCP6VhVdu3L8DqpzlOE41ijXfhcLMLyS1/2SqJRsj6fYuZqjrc4wiwNoaOL0O3eWDa9sY1Rn
QxwYtgdlW5lFbgB4rVnJKDHDeHEE25N9DeXz6xo0LwGGbAdpInqkTOO+5ztJb8DM9mZtWwCmj06X
W7jC5AsdNb2PyCnrAd+jTG57hfX3H6PZj+VyuFpg/VGZ5M3CBIjFiZ3p3WnRtbpJcyQgFHnssQZV
S9dB2KusvNYaBdPinKcbsKwWO+HHnH7obfyiVa+X0rTqyrDh2O+Ziw6hYGOInLE+Dz9g2EEUoc2E
eK9nOQu6b3/VnRmwuW4bc/8Y6xUf6tnhZmpjlprqat2Iz+LP3tFhPnnz/flnTbJ2LzljW19YSSM4
aDDIEI+Xam86fFyWvv3XnUfCHkjNqa/R7+M/WsmCQX0DGlr6JWcpmHO1ZacYergd44jui3txZvII
dYQLofD0VwJ8BnyVDxB7xBBAyDibkES9q3uWxWO9c4ujTGuygnJ77rEqhAazPI0cK51OFPrjPiuP
pYSu7AxiOs3CuuFy+YjupYXKGAFy2+3X/9AZRMbicDNmthiHjWFlki8AM5GeI4UmOYHNs5cKtXWb
M9zeyxuTiDRekgZMc3fIXXtlRvxEdmzlMRX4K3xLlOB+gyCZJ72H/iyewqIeKNTGcC20DRfjNcsL
i5d60ZvJ6QsrMdJv61l+76SYf9hGJfBSovWvd3v4xPPwLBtNbdhkUtY+SEYreziCDLohP3Zu+Ds1
neWT3i549TdUrcnvEf9SCbNsNIfY9Yd4BTyS5iOI/YxZmGemvZaFTjX/bS0eVM3Fd416m+znl0AN
knig/GxFwfCU5SHeip6CdLmJlgJ+WTHGcRoogT0Gol4y8Kfnv3awGaqwXjFE0fau3DfijDUSOBWi
m6yCRHfGb9/Fq5/5V5wFyLuaF4iJgwE7xoqzjGeGQYrUz5APrJicWtZmadOtLp1uG146TYHs4KwE
MaTp/hMPwhi79s4BCEmt5tjyETWcKpCHKfShWoilWSu8CMTsHINm0kEj9q/uoSKJsx0BxoSluSiq
SnWsrmQH0kuWPzkvz5xptvb+C8A5PX6sjvenBLn5frwPtbmGnhNDHuGXlMewtn0XpYvYLAIa1uhG
gL8eOkJDF+6ZvHXo45KrDGMrBg5OInbjTWkVtG8OKq13JBtzbhOFv5gEQAA5S8SdkrRy8T0EQwE/
do3idH7pYftE/k0IHlGW0g5/Oe74lN6RlNnfETac4f2anB46U4eIpiR2XH+XQzO93yxvuhN3rXSX
zbxBUWg7aWOlfHslvyPXDunlCy4VtvxNVBvnNC8Au2D0CECxjIq6eZJOXhBmvmYLMZP2UyC8RO8e
a7FFxJsImMcVEXoJaITBXj4j/pJh5k5g9zF55VzWfEZRcx4+f+z2OpHa7sRccm+9Wgi95RJ37THB
15MJb3Gyad8AzrQsslrST7j2jhmI+Nt4naq1IjigDo853gmZzzj8Kl/MHR7X+XTJ0Gz2fdyR0A4O
PNpcDnHm7ar1JxGcECTHuPHL2rsUvPGuRFdEsUndYUPr4x8biEEoWsrQAa0rWZHg+tPrvxwstAF8
DXk167JEWwL3TJiiDQMXUhjP5ByDXR7HOkV1s4ga/57dXLiYksOT9KIlu5SjzYQPXvkCTXflGjQ4
3lvfGAKrE14OpEUkA3aC7gfjn/XseD12wek4R0VkauSV0n5+LsJ+drZuZp018/51jVBBi6/YQxPM
yzfLwpUamDnuHQkzEA1b9Ahi9vPe9a0u74OWHjvD2avu/NgAORhd4oxvU3zroHnNgqeCTCS0wff9
g5JzRfdZdaePUVkt6XXsz58N74uyKphSiz8CTREBNbx7387AynNd8zSZZIBaUyAUwMCV+GIlXD9Y
afDVSmWQdDtiIglpl8gCw9FZwXF9Tx6nUo/fRiTLxTh6jrCCCXI0db0WzZR/jHiFfi27COci099Y
vq+FNOxtjSXuU0DGYL1CCDdjS2eTU2yIIwJD5nQqYq9gCft9ZFyyr5UucEmnZifzoYExXx3p/YTH
XMpwGAK8AcCRTRGBtcyPrzmv3cvUDQ1amaRwfc5vBY+iC8LBeZrBhMLWjZEec/v6KQR673k3g5R7
5uUwdO4uKSQoh/yMSyCTUuPQFs21aUkWG6C72AeE1M9jf6IyiDqNbKEbH/GyLch6R1nAro+50CDj
XMe7WiWkOGdcmJIND+c7tnhue2oUFrUqdo+IcShVkjB8QKbnCuapCm1ey4+CGzk4+03LcOUyn77J
W4J8/umKdCgz/4UuanKOuqsLB/H71fJlC2V+zC9avtRpLD6N1OdJKzZZjbBdYm5jVZ2aI9BmfJyZ
VO5/3zVhDZNUlTEW5ZtYEUwbINUKEVBC/Ox0DqU8hDyydPaBf+KhhLsAeMCXFRAAy5yhc0N58BqT
pcFdylU7hLVMswQmWklmiSQjfi/tgD+Z3BLknu8963O3LgjDX2vo3Psreu9o9jApbGqYJkWa9Mk5
eFv7Gt/U+NtZadkGv4U/5fxXV0XorbkuAyDlfiATez2oj/e56bS/rkz8y7i/wOUntXxpx+AT5pS9
OMODa+oR8EOPmlQQiehh4zj23XMnKRAqrmsAc0k0tfoQtiOdr2P3hcR4/Fr9lnkb9rmWKt8Qavwj
g/UiSdzZa2GYaLFqWr3h1aM5X4XQvEh3VQGMV/atMz0ECe+akZc5Ux7ad7IE5ZtEUCpu456D9Cg2
07wEdOfbCwvbvPK2pvtDNvaBvtrrV9iLt2jZN9NyrqG9I0VP2nKiTK19ZAEvJUYm7pKkT6wvuyXC
JAsWENIC9PdQmi1olQvzoGjdrzIRwtqpnJWERkzN2XUUYDSqiiT9N7SXNQ5nQeaaC2+J1kapwlE+
11QB2s29RPocx56NMJPViBUNjbx2oncDw56qKU8lM0cvtPlj9QmLMqHq+f7316MCqIUvnTmXE5Ie
Ai0Q5WQkOZAPfixTkicCEwOjOCdBzptuKgcnTT4A9z6P1dPvywAhkS9Ns0eGC5a0H+Yz8TPYiFmQ
B1wpOVRmM/XYfqtet3aZmkc/XoJEUAgiNIjuZZjY/VrMz4yFc394RvQ8JprBL6ytOVRCzqkWiQ4/
2qB6MDVir/74Dnz4cBNkD2uZppthD3iQI52+wV3/t03KOX1hgFVdigpwRqKD4cYwQK32oo+XBp5Q
n+trVMI2dCXgtbKpkmp8Y3isib2GLpNbuzw3tFiX6diqWWrnyi2b7joy7Kd26W3f78cmsymMpojB
ovJqbXZRZXqjFnKi4QoMcpRtr6EFzNQEsdcc2QjGepaIfSRI3+yFZ7E6UunPibOJ5ctpCHOy5L4f
1KArODkLBVnYDgOiqC3badOK8qf2Tghc+1hR7JAHjgpieANefOYUJaOGjEIlERisQfNbJ0gOGBOx
DAwTXHFoKcaHB7bwulWGfo/FRWQfCu+aJm3+pgpNgB2KDs9bKQljXiRjz2Xthum758xtwzqj8u1b
Z53Ey/7JatMdvoCWDrgSkqEB+vRk7Koa+sorQjPSNOs4VyCZhGQ8FL6/ffIXiidVGkVeozk51yZy
aSjHaYMY1loXG8w0bFHcUfPjCbRCmQLANVOsxeqbnXFCw5BAYNDj/FfZbf/hckcoFjFuQ9pqee1f
rjGxDx9QBEzrI0aMtEHThQx4zNssKaDZDDAO3N92yuB4UQZEOUWFvji67SxUrgSYCaJHsqt3cmve
99j7xgZp8ynH4dQjhcHtg8No+lZvLWGi9SW/CQoeqrNDjv+GOH6YKI2I5irZnE0Y0n1/I/nXHvyk
oEGbZQFFFG+r0tPxvqcCG7GfFeaX6TYKWt0fcnBg/kxfjVGKGneQQVQtx7D4B2kbbfY0yv4SUEBN
EKDsmpeLBK6phWyy5zC0jBHt5uBSSQK4z9zgLBWDZvBlYPo7CVvBpGWyYCo2b05pnp+LZOHmHIhP
TkuzO/fTHojbKsl0mqxVzDApGfuBAKZIb07UAmjz9DScH/NKmH7eCEAd+KIuJu9xXI7725XPIjIw
x0EclRcjfkEMqbQStOwZzAc9mOhFt5lkeJg20A7yJ7Ca6H7mtUlKF9WdkzokS/kGwjro/iZTZFwR
eKIJX/wHpUnahPG2BgbW42NA7RS+f88mPQWHBbEEyTe7uxZxTjqYpCTFrayecDQjsZxZB3AvQNRp
3/gYLVJdquO6bblhJ//Nq9aUIQllh6mGwyHeXgVrQ6r0nKNbrqHAL/tadETddlslTJ2VHo/vJn4n
qYPYZLprp3mzqehzz3ijvP4zQtH0ZxsMltKF2Va5M9GNv22UvglYkfstNEGR9hFagnUXU5v4EhXk
sdR2ErDWhyiYmIbpWSnRcyFbU5yeKKZOrFEQnCHxpLL16+4rciZA9O0RxM4ujQ1CB4ijfygE33At
IZl23SWJECWkK5NA/Br46Ay7pSuBZwsj3denL/bKXEVEjKZauobhK47vnAK851qbdFbUmltDxIni
gVwK1voir1Q+y6er8m3L+eFix5IZyUqRE8iDBJns1jVG9qJKpp3QrOplMjapCD4yBOxcLgmu6O+7
bskhz1GUtCYwkrIbVwF1HQhXROkas0QYDhd93ULGbGKJ7/nIX4s88lN5jA6kEPA479FsrfC7nYyD
XsVT0m422xzBoHG1Cl9yVYTLdsCa23o3C9aWM+562+cXS1OsDnOroHCHS5DkpLb+AsMKOHYaEkXx
ecIskxoZkH8vHgHbmgTkpyiFK44acsG+/pw4cXrQvPPLYI79jf9p8HQMNgkqhsAJzbTOp2347mGc
nJNXDCsJX0z4e/HAqaMVC6tzjb/WKMd5p5RIRZZE1mCrRRJ/UW+aVdSxp/QMTXOLZp/LLqLDtwoK
Vx4nOFp16LGRUFMKGVh/UiRoV5lNA0OMItFVT3W1V+zb6x+vgzA1JlrOaMKvngfeB3QV/BINedzN
uvtYPSj9McXCNRKE/sn5DVDOg39y+PwXcdVtU3kEP22CEY1RhF/5lIhZewKBGkNFF1nd1YHYIULz
CTuefWq4NSQnSubMqOsuUHNrr1Kyy9cPQ9seiv0G2qD7BcC7mrEYmISogSNuh6KHU6S1xUKtrZGB
vgEn//Xy3XYKeUXQhDAUfU+T6sEeOjKpIZG20pN8X0PvUPgDMmn80ykSdp6bt+pvkv0C7qZnkcYr
R1ENSEBlVJMyN3I2IzWCr6YdiEkAsQsF/NTNWTd/ADgDCVJ+G0foAoL+Rs1PUdgUdB5M5vDqAa0H
eIrpQpETndaXJla+m2aXIesZuRlEwMyanKW6TZQ3u4QTKFAVff8vJrMAj48IU7mMQiV6nN0itwRt
+cLRyLQb/WByllhwGcRrAU/JK99o0VfC6YSHS3uob7qIDvc087nrCHIwgdSMiBxPK2VnznlEt7Yq
Hub8LG1Qv0QmPMVOeDmvHCvhf7MBB71BE2vpWVtUCNkmUyOxna4ECbaI8XwrcHaU3pktFi8vdZNl
uK1VSE5jLzClp3ddqATsHgc1Ypx3FOZ5AkrjldLeTXIhT+sDV4aorCqS7IfB6t4n6xEdZhBxF2IH
7C2gjR0YDIR4LsRbE4esFcHNTp14G4zalDtziynFJS1qJsvCTo0JoA6DyVQ3lp9MK3Y6spZgTpFb
5y9epGNQUBAo01r7ODs0/tcFfUC326Laq98bh96yVm1ZD0pwv/UfjbDo1ctQuOSbj4FwtPkIjqfm
UClnsb6c51y36Li5DIZukOm/dXsQ7Vgmn5XlsRgHkHPnRUr7EwagtW815x8b5zOFc7cUEOZPUIia
HTQB+pow7uatnLo5+ysFcnMbQ14FjlU5tT9F3ChsWZqjDYp/Bh81WxOOYQt/i+yLSU23A6VrHZpx
VVZ49taX/mWzAqEJ6vcXflcQMyEaxVFVOQb2TM2QQKB1tsAtuH8Ym+rlawrizJRJYOST6FRg6e4J
MQnRBsMufxFmK8Tkb6fqKUGzC+nIQRW6hqkcdHl72AUnKpo1qV+CB/vNZOkVAtKL2ctRjOCW9g79
3SgzVnagvR9VKAQHnOYZhauDHy9E5CT6tQ3uL2wlu4lExvY4XTLz0+II7EvLRPdfEllE/x5KwvFP
Wc4jMwlsCt1uFSAI8SuIReeYkhYESOBtWal4KrJRsw1L+NNgAD4HDMnCwJfxO7hU+KDbvkVdeCAl
bmt6wzXMsfXkZ9jRdARN9rYprmAoyJ/0/bRf9YxaK5Aw7OqCHMuip1rqQVhXwyE+5O+lM95YFNPw
ZZB5wIES5+iduXkzsFDgEFT+eVo71Ul5QoUtzRRzCjaudVNL1M6R542hcQ0X0qWrkzIoXR8KWuJa
eP/thWKz2dhKJwXJnAO3MSFAJQHnuTAtd2yT1jk0mXlfOkU/2jJwVmSkfnGaMTqK4Q48JMgQdeFb
x0jbSPYMMHVN4c2kMgYqsLtjjl8hPIgFR91X8IvYfBZ0u9yLHH29p7+hLa0TQrbPP8SsF+qSnMuP
4raQw5S5yPmAReMZetEtwWbCEq0cqF3Fg58KvTNaOjvh1il6FBUaESp1Y5CYmXUQhJl8FZk+K6AH
2rJNyMiCgVDvrURKrMrXW+rn+hygKRrkPQ+p+DG1G/bwvHcBouzDtdatPYDXft8Zg8bw1AgaRd7m
AEw0w9t0RcKE3d0IwPl3SNXQQ+TM/4s4B6Uligd7ZFtdcNvZWwp1AIQAQ3dj7SXMRoTyMPTs4Hr4
spQEW+PQaKU1OyNTgUnzjyBo0y9hp8PnQSirOAa79M4hySDNY4RTjZSlH1kfiKRa/t0SpwI2+sTQ
k/mewesyBAtQWUZrymy17EvYc5XimrMh6uojqZZkxPO+HGONHo95/WmbZK9ZWz3IMZQls7aVVzER
OWZtuQgG/FX9qu3MOIDtbgxCca3KvVKDSDDARWAgYt6cYY897jjqYBU17eXf8/TjUzV2AQzEDaQp
cHQIyTh2Bt8butOJuGUrfWYCB6Oc7qq42xSPPPVOidP/jNTHWvlOHj+c2IJc4LxV1i9znjHgNfbI
T2MbwJ0cmZeYptSA5gd4GIzxAdFtLD24a8vBQti/6QDTSW0LkPI8M/DbiqhOdfCeTCDXmN8vmHdP
QJbYEh2s46pbgzKnxQCSC6JIAKL7lJOhCV1mW1doyt1KuhpaEuks+04GeFjYryP8DzbzsiGyw/D1
xoa8xlY11aAl4yno7RyCwidSNvlCeYxrONxP9GhTv/ysavFjKg17BaERNSVCPHRjXoLkdV/Es6yj
96uttS1S3GDPEgs50erCDLY7hoWbaKmNDCJk+lWozay7Ybg955EEyl5XYdmcEq6fx4NrRwfyUfGv
xj4icECW0bejDSOU6jNTM6HKz1DY1KZMCQg6K6V0sUgYgOMKCTWmWeA/vBRtEpS5siDCtcmBQgg0
8ey4YR7nm2/HYv8J6duJp6xs0IcyO0sgihdvu25CJDYWzidEDHRTH5NP7IkkkMx3lIqz0KUFIYDT
Q5P9TOrSTkxlUk/SwWlK88pJcPNG31OEZ+62oZiqEfHxpS9k56U4PeuIOdGUPK9yiucQG4qiHk2S
azujMHdyTvADFCKS9J/O7uWW3YA7hWTN2vXHm94EYqEZzLNyE1bn61qZpxKHZaXvyTPkB0yNuxqB
UOeaqcKXdKwnxDKRzOaLQWAOZYzH6sePD1//AuHETqgVbd4V+4gYLFo1qm7erUFbLU4nE04FYZfc
rKV4m5HRbqz+PgRKJqqt75q45hrqmi0NZ+0pEELp6XFsFund+9b6WZvkkFh78Ulwe8W8GwDpX4u5
iKzbdoosQPjJDb67NfHz+AZpE2CEDd/PhONJ3dOOUj+0/GdT/1wccofVraazPoqTGW+0INolj+wK
jUdcdEltrTZOSS8IXo8ODh1S0X3pPS7F+huHQxY4K2IDHzPCUw6ll0Wsdx9FG+hZVaXTR+QIGAFc
QOlMVXwWtvirCzPZ/D972oJsxYdfN93/sfKeBNTMHkcWvyGUbZPPcefBNJR+CK+YZ/oDOfSAQJ+E
5dzNb98DLXijfbBRGXIgFEUgMU+bZB1lth2SxEF/4tLkKyzy7+iQOnlVYQIgIDl8E7LH8jUJRwuD
EgLJpmqSjmb05YV84f5fdge5ZkO6ZG/jEMMlZLedq0rFDVkJyQuLwc3ucyZXsMze6j/f0nTLv1nf
aaMX7ibJFemQfQi+OmZ08xmcq1X9eKgIcB3m7Q5/X3iyQg/qSgtyTG7irdYEn+Rz4qa2OLp/hDY0
qGkgAT9W26UvZU9Ou4/RPSRzcmxpbDjn3HTE7I9Jm1MdfqmnxMXaif0br76jyFWFJuKrwnVDyTTI
U6RaEu40ljfKwfr+LpPaT12Q3riOccM6H68O+zlHYQZoDjdnyjRmuCPGKewR17UqcAjQhoisl51s
SMpQPs64CQHK4jtv6M6M3hzozUXFRN5oYvUPjwMgLmkUrhy3EBvOKft8jbuWXY2jRrkFYjdaqOeZ
rK2x7u7nI/q0qwlBmpB+Y0RmY12eqIUQqZunOlErzYrzGJucPdDkB5Nbqt+G38X1Y5KrCeeTCSRB
K+b6EAK64xwzCydFoaLlt/G7c8QB52P+Z7zsQnm58fCqGI+oZm7w0dknyDa3jYbxy+Q0c+y0RlWY
XN6XNXxqnwo7bRo1UERqkYUzoThYek85umitMfNV/oSxLdeVW6K8ehR4SQMTtcyPP1AVxvfwQqDE
Z85Dmcly2OjEm17voVSQalyt7jVQcwn8V0Ja5OVeXXT15zCMfNJ/VaAHoOFvFztsHrjDCg8n/Xa0
zqnpYpVAqQu//Spz58V07cbICB6Wr5kRYZHRMG0BqvuJg1+2HrSRNUXAF9QZd8m7oZZ1jrljslFl
MQO/zOBTMgoLDgzvelXWYH0RiOAnMx7PFAlPvnK7SsR2TURhh9kQLYEC+OEPrUcZL9Q1GCKIf/0C
pHB5iknRdJSCtmv32i5Dbc5t4ndTh9PNIVWGgWlejEYfeFtCQqhP1+QywSFR39Dfe4exk2CTjEvf
kXBNUeSzHgjbJqX+/1S6R0eznxYwMEcUdfDrzvV3u9PBcsFfSW0zaH7ZLhRpOr38Ey7uJcAmktIq
moNvAck1PgFYzrEkTRpIjLdsLgW1mlbtvnTRuFhS9zAIllwvcNRZABMItUrdPjgw9DL2Ag9XkG3J
LJgQPBYWRD0KguMAV9vW+EXq6fS2iJ5KxKEU5OvYZ4PZR7iwCKeZxNcz4znxTE+NU/ozUP0bBFhu
6FE399bsVvqxCgwdLSkWguWB1TFyn8IDkrngmm8zX0vR0zCj6uA0wM5aLeXIzq5+V5MAE6c5I6zT
NhH0mmKihmqrnCZRjgmZqHAx9S+aghmXak6JCXxxxmxk+FWNQrBelIRtMVD8g/TrPPnScbpZkcoV
nNXVy84cV9Q7d1PZHgpy9perwEwyLpe+z6+XH/TIE0V2vRmpsA2/kBreHMd6ObkyKX89z0Fif1SX
ldZoL1sppitH/osDoUmuM6Z5PtpdhTi8EF+56mDh+lNP8At8YOMs+iYEPRWEad8pqLz9Rnr3K5rh
o6OkhBWN/lUWTO3AWo6KBozs8zA0+N0dGA9e6dPu4RYBfn3AhF7Q4nTNub8WXXY2kOhyEESSP5/J
6h3+VJFNxb0uoB5hEhKNK36mtc//Mv8vdeKu+iVnzWvbBZyCpGKDl0FLoxfYBCtmQqcmerdeJCZM
PpX37J1JHxvsDn2i65rJTVBxOkhqnV585lofp/yMQDcUVQNPoHC6cgIs3ckLD4xbK9MGpLxs0d6l
J/IHbTpDXhypla7hEAYjoTbC8OT4qn2wWY+ErcPYCzq3pzHGZSp1h3W2pRXqX5KNJ8+S5KBV3TuF
lZPD9mnG1zv5ruVh/MJUcNb88kOcVI4HA9iyh+OzNrzMlRMwgGvU23D2EP7BtZVKC/j8Safmbm6H
VFi3wyjQTcqI4s8nlidaKeAkrzaRqHxY8xfVIO90Oh4VjcZ2Ox2LKK3/sMWgXtIGJB03AKutTHcW
bgB+oJYJNjveRVG2FTKl8wLzeIj95B0wA5PJndXOyO0FiJN4sMCQYNg5WzXKhWQGhmOKA/GOOWRD
8ld0Geo73YLGXz9i7LZyQMr/rW4cHlyP4Ur4V+P2rV9XioxeQ8kdDQES4XOWobMiOVl4Qo5hjX2/
hqY4dWiZUo3ouR+TtBldvFVsHNbbcekndXVxElicee4jm2pgrZ8n+PAIHReUFgnYLV1tYyDdANwZ
r7l1EB7lMWuhuWhe913PvnR7pBJCokVkaT+zJGVQ2rS/EvMjuMHrSo7eXsKSPsVZom5ShNh8uS4T
3izLYDHzJw3SUwjU1KxaEC7vOR6iSHeOIFrjtkz6bxvnn5bH1fEB0ZN2PPcqQFdaeV1ElJGMG/Vh
9FRtF6QlEV1HMBaRJIvWEN24qr0Wl1cLMm9M5EKJl7AcNndHreLzMY8vyOFtw33E3I895Ee6w8Pd
QGShIZcYlGUGS4sVJNq/k5CI5xkSakozkzKdVZg0X/v48XI3e3z2U/sg0kzsZUiIDyUlbSkWoX0+
+xDAi9iNRYE4fZYjoWgBmp1FRNfUw2+iriJbRm8Nf5u7P7Fd8RbJOnIQnZMixuce+kL+PWZFAyn8
O7g4KA8kDFde8kQ8RXWw56lXplh0A5e30UKM+hkCw6rXGkuRiQMo6h7vb0J2l1AnOe5hhhkJMJNo
V3S6ItxqamNnkgVAsq54Nph2kg6Z5NIMFLrA9MG5uEKuEhEXNe8w/8lgFUCC+GqwMUyU4gUAYuTK
o5rZUxz/jKU2uq9zHFAAX+toAS861gtSdlozpGLj62v/trXD8lWlH+tk/CHht6YpWwlGNgnSc1aR
hB7WP9jQpzKdCzDACwgwzFxfQsaYLJeuSOrJ0Akj9KuecOZdxV8AjwbvrYO1f+LJxJqw6GGJOPTN
5+zyroiAKz0Aw7i/CyzsDE4mo1CIZe7Xr5wxZLtT9pG0QdTg0RT40KAZhSz94nNR/M/CvyqqSheU
FPIr3xIU8/KBn+d8zOjg8R5n0RHaZu9z4P2rLm/leF2zEMLv7xIXx6Vd078e7bYlOeNTSICcf/82
4wo/QrIQWyrcqrmD0kSQMTd2RMesw775y+6oXUuqCarOyGC4IhVJDuNqro6EgaB4dWAEp8AucXVD
/HF9UETGhzABdZ0oSjPeQHIEqS1wlk0IeyVdyYDLLgMl9aYdd/MAmjXhrfc19oiIDaOTumSzPKvS
GQtsAssAlC+fWfNC/ObW2Y3eganC7tGs/sfjRb/0h/sXo0VbePPz2LOxe0UI5ll+KX7uMb9QDqZe
Ty6jOucrd+ju9p6Cm7vP01E/o5PfCkVf1ajdvHN0+3z9N6dX2ZCX56Y1Vcsenm9CsyoW/0j2Yw19
OUnJ10YfWU5S91P11P+iaJCKN+gZkdottRUpr4yPU9y3hKGdsk3catPURVkVuBVwAifxscd7Cb5e
XG6MVUUKXTi91whyWg8nSp/AA+mDlQb2wjK7W82eCOiXyfmx+JbhOnVt6rKMD9B5IOy+X8dAGJpc
eZ3sQwS4VY4ZW0Jr9KcfFsEsXBNlMA/3vInHUEQD0+WOk7vT1WhvMfjFtkUIQ56a6SEw0DkaANa5
Luy3RE6RyaAlsIlAG2pJqryqHSsgazt02//JKhJxqkZqQHZCh9NYA14fZ8YTzAVOzZUBrgKJ2Avc
rPvuGwHWovPsQ/yy+KLIBGq7va6UBaF7itwyjfe5yRzhzUCIGomS4tL/Hmh/0ZcUgh3D66r82pBr
BlBg5n1DAabvdAAHxkyQ/bS3qTKsXkX2AjeKOJQfF54HJXpm+LWctAz+kGWEHjcGfnjAj/1/Uwii
N+k6NS4tGAP8WNGeUzgU+L/W11XBAwGdMbdiYNiouRusmUT7S0bUpgXLxKGKUJk33fBZ4N8otyYO
MD6IgU78Se6tcBFX02KkHRVTqAloVgqWpj9InpOJpy82WEqp4U5Pbo121qobs/9+c9sUmVArabbz
41Z6ACMIVBtFuBI3jMzD/UTpPiLXKu6+5gB4UnLHuolrPvg184fTF8WI3vNiMB+78N4mE2C1SZTc
rPOgij0ieOG+YucbLz/VL4+W3CcmU5roDkTCqvt++bZKwJitsHqs9cC7RcJ8UQKFa4Rv917sW8hT
/IY1HRtOLJo1Cf58nkCbJN+4rLVH7NbhdwDFbKrEv7sZCzz4JE0WHYkC1JUJTsSn7H/lwjKQiPJX
MxKmZ5+tnKIPGWaPMorPbYHad36NZNPL2nnJ4OZ+XM6XRAk8m3qA7WvXGtKI1XgQki3zdLo4kpz3
XVy1OuXuFcVJuJq4Ds1w78w3/KwlLhcqnouRpopRDq71yiW0CHkZAfPpV8NQ/K3xWg0cXpZxiGsi
zLLNWNn9sH4CAQDKylV2uukppi6XrUXgx6z7+ko2cFX0m5hcA3fy3eUp+U2qAFT3n5fxT+AbjUsk
kHVRtHqv39lWBKNSZqLHDdmCSK9xAqrPXYVz4wS63o9z93hHUCDv4j+F4hlmbLfzF8Gz6N/jQDIz
X1t6biuXtwnlh8qdUrTwzOqx5hlO2v6f/9ucLlgeTMvkGVL2PS+tUUkOkMiO3IvWHLiLNMKDrfPy
7lYBGU23ZvGsHiEW4zeyiciYoa+bcEtrUiSC2Yzw6ABtb8GXudferOz7O2giny6+lsg44YGRX+qc
saiGnRqfj3vV6WY0+FJLzpuFQ8sGVh9ueG/E00mcO/vIlNJD+f7BVWfrbx30yWkGbBWa1AODvP4U
1VEoNT87DjGqRMpI2HspYQdIRartURP95XrGkCemqPBy4lmxv0LI7U8P5NENVf/jMT2SNzSWpnNC
0bZfhHEd6yF5TFDW4rhcwHHHT5feV76Okk0bSKmBSQ1UhHik2yFMGVu4i2mvGNvN+O63MLXsghDj
9HjyCN3vsyIGSOpTI7rkfUcqUQnfh6KZQvPBP2ai+wDyvwcuWc62oUvPoQRs+1t+W3prUbnJEfIn
VnlbloYxMKNJntZ5izw25b0lxMm/mx5CHaXuYOuCGfiM0FuYnB0gFvwVSY+ymM1TsDG1lCvQLRMV
a8bX0Cs73B5IBPdHAyTXcpVN0Bw/8A9yvtztkdhWPS36Zb1ARTqnvDpMKjAbi5sslGCttFIHrLFP
p3hBc0BI4ItMds/3zW53TV6eXt6157Om4ieSNK9Ep3lPD6+dKRlCCiCClYGnohzjh56816IQWrlq
FeR8dTBaMukb/OtWD3QKd/MMs3yZG8DRA2NxPO1tM//2T97zeqMyWcGqDASAWkWaJsZGxwGKcUzE
QT/Kps1fSn4I3pBCtpSOFeY5pseAI3USNymLS8pIuMixHK3VFK0Pv04Eaar1/0gw7vZciVhOPAUn
O8mCzpEW65JMh0o/mVr9C+QcT/mmDy5IJasFeWxykRdsALQtuu7qTD9cYZIh4yeh28Tu8A7/zJTm
Rqr+JzPoFfBra7rAa3C72Espza9AyusMI8v+51QDhZLGRNZgpu7fUZcFcGswmNojUp5K1TE0Ff3w
4jDdAQLL1/EmIt3Yvt6XRbW6QCvcyOmSmDlc32sP838w8r2+lWhySfGPWAuEGC2qfPk47Kp/E7Gg
dI7G+NkOlLtaSjLymVy9sdRlfQhQGObB1458R1Uf2JY7cwBMBNXVv5IHVTGkHO01sImTDCOx0//n
BFATHHWjGMC2hJrAJkaAFhappoE1659K3RvoP5xogXPf8YWngRMzkCn3amyPYskNOss+YdoQtJFc
2lKoMF/CUKjZRx4jmOxcwYshOWhfviBOfi5j3ne2gwBWBx2jNTYWT/hgRRmjNax/Nu2/G/V7kPIG
8ioex1uQYo2EzRUQAKONFpdjv9a8C1hJq2VPSSQZX9myH/Hv95Iq19lrHI6zHL5Q1aY37DHVy8le
izpVPc0qOAS5FbLuzJsFaH4a4m3wcu85F5HUirnwri5LX48iNkqGN2F1mmGTywFQvkwsf9KyRlGo
2l6II5iyLxRe5T2qA+hNXkYmdzS7nHBPD54WA+hYyERcnLZO2KJ5PsMvmh/EUFIjmCD8us7ARsIW
WLmVSPan7fqVW4dnmstMalg4Jlnfw7UNf0jJQIHYq5q2ImzMvwSLOzZj4M1YwTYJqgYRXdxDbZSL
SDRL5zhzmq+qseww6vMJzhVHmXgh4V02VGaMteAox2sZivRfCRr+KizHMEtxjnf39M0bnp8lh6c9
pH0B12XZ3yn48iYBpGZeLwnm7Ux/VgiYK/KiOFOP71w4WofnMmGFLz75dbKPIgxQ7hN3YqqyxoS5
SaJK8sqH00iRlarpBHa4AgP22gMxQdpKK8nLQsPdtWO2N5nwUZBhVj68FgpI2vqmjL3htJ7l9vbz
OToQO9ADWKkgFyLZyCPVMQt2wTpPY7szuYO3Kth3ijujyVPljCQvNg6OrE6J3ehcsUwYgOrpa+HG
sKMr1J7rI8uvAQ7A9V+pSTvRcXfeqqerfSrQJ1h0giNcSiEHCcRmtE8Cgz2ribzOnYjwW8sCZqr4
m7N34xxD2+7PuD+8Ze1Bxo6SKAZ6G7U0h4jg1cF0CDxqfkzbZspmun4z2DnuiJ45cnVLZSGp0uYZ
W1JvkZT7ZMx3toBG3kU1bcA6oQJqGOMEM83ra3zAJGugtpbpv3iLammFH/17/3t7Dx6GC+VpEWCQ
+IC2oThF9wBDhKnFg0hjhnuhF5F5QPQQEiQyO5JeXXaBH8NZS6ODtHQnAkXhOCLzEQKlsYSEANWN
QSt0mElvem20VJx3IfeVrtEQfS07RAg3TlaYwOSOqsYgiE8TDRi45dOewwmXcpRRtyHSW0bar40P
/qtyn2sYx3p9ZPHBQU+Nm64LfscC5gW8X2hvXFTVEn9sKYYMX6403gya9LQI+pB+/1dOiJhojfj0
S5MZZtpcv1vbAcT1QwwPNPMsrBGZd0A8h2CVz+TZKb6+a/ZKZMGE0NEWtrvjc/8bV5efI6DU9YIP
g8Cg5x1v5qiikoc5/2Gd68oJWG2XYiaCmhJlRnf7Rj9AdbqPZ51imVdAE9lzRVsUQvj0gqE4QE2o
bI0R/yAXbEkFjGYFmEn4qWehv6aMAzjvh/6h7AgAqdBX1iEiU7spS50+PmTkx647fGtOq3v1aNs4
UAjhrz02Vd61VvpZ+Lki437gWubMSjbnhY44unec3MCpqdExa8FWVsaHUub1Sb0M08LN5gzxZc2V
z+3dToOj/ygC2gbwv5jdtGUOtv7gd3rdOQ46owlLqWDtrUnwDPc/s08akJn6fONBCXxRrY4Pqr4L
czHBaMDUq6IxUutW4ZmUyPk4bHa0lpX10tlBBXU5uNcRLHFK3ip8XT3MPaIUYZUqriIAWxmtBot4
dnTBL1A2o03HNKYXos8mcyfeJ/a2TluP/t3rJj83cJJCN7bQ2f8MWu9+r0QikIzAD8CJI9EMdHWF
dEL7kaBApqZvx/3d9WGZnMvGu1b04N/bRJ4ZqcIUKhyXtkjYkgVAWYKbO9605kK7OK5iA8hdeQjY
Bqj9CLp8FkLtQk9iZU0Rr9XRyNUZHyp0u6RZ0btSnQ87tfEHu5rBQZ4ELLJxs59BYTB4uE8WXt29
7cHOTF9RF/KE109HNOrw+czU4QBbGoTlFWIQE9rzRp0Z2Uu4qRyZQtbWJVe8JV2zfiy4iWOVmHKb
mi0tsVsaIChKmsIATaUbFo7KcX3T+Ls84mvx52x97/WGRtBy4tLB2w4Qvj+Jc5KhSSjSY3yGl06Z
rHLmkJDkb8/ij48koRd4mNCj235vCo94RKsJVJfCta+xDLAgyK3N6GHbY21SrXYj3PsOBqzFKoxP
yIYjXk+FCXIoiBfi3+gm088Zqe3QG9mCy6pi0pecyCB/RIHJ2VWalcu1JybY9B9SDYrQ1bT7MHdT
5fVLRsN8ZTTy3zXrXfrAGUGIWHKJnNXvBYd7VYPf7o7845Hmw5cLsXKU+Gxjbut4YNfns//W1L6X
SG+tG0H5YdEUjawxEKA54YXRLeHF9FmTrh75MSkTa+Gg4jd/VyQCFKo+GwcUi+NVDgqs8UXTy2co
PM2vl7lLZKsMF/KF0Rqqob6WyYbZTJeQLwRh78duNA+ispt6/v/gzRy29J4+T4/yoW1GwlvzvEKO
lDmhNNNBqmwTtZPPLThulg9jU8sQ63gUgkivDcfAkoykGJAL+tINYx7Js+DYrl7iRBrij8wHZHk5
0TV++ymIwSoYW5Si5pgUWPUShjpUza60he4or0VYmex8ksFsKlWpy6yXm3N4NTXmOE/miZRLjJV2
pdrkfLLzAXvk6HtMBNDbosu5bah315HrIUa9d4nE1rKX/5QVCIXRHRt78LpGyIF9j3qrJAXqa5eb
lmHPjMrKMRjCEhBdp9cNCkp9CXUUNNQiBop4m1JD2jdtNPwzHtaR+aG2YxW+0OSZJnZ4Hacuon86
c44zFmqWyxIQ4XAxMA3Y91abw4R7OtyQ6awRXL3vgMEksPCRcy5fg5Sq4gsXWKEfDV5Ih+acVv5/
bvLyxfGSEU1FrgaNLLlpgWjrrp96oyQ7v8T27dl22FkA5yGFP/5M+1FedYoXm5VKciQrS/4d29Ig
RjdX80V5f21Isbt5TYe6cd4OZk81Wm7Smg3iYm026IOX80EI5g+RTzkodPN0hFjpUmHwKBeFkZfy
gi60dteBNZmfSnYs7js4tSToSlcSJAI9POggxSjL8xGIka7JvFr+J+LqCPfrN7wwW6AUkYPl7U54
VZVM8b7vrRsZkUMIWv2ken30nc3XYVSNMjBZDYnEWF0O2bKIn7i9TgrA/TEJviVD8e6P9MYAyAxl
LEMZN/ork1kxQHpZ7i5mVXBFL8yKDlhGrZ+SPQ/6uSkl8rTlwXtcSCaF2JpZlEoL2IjRQap2WViy
m8MLYWh0RVXDMytBG7/cWRWfp/jRd1GdFPTPkpxMOyH/b8oBlt/EbAVkwmXW+aBD2L4sA1e9Hk61
f9fL7kIBkKijtxzwGGrN2WZQlZMOoY8yIymYUt7Ai3/lbiIbJBVISj6wL+aXKZ8R3/pCLFNOPokB
hin4SwwJ9Ml+OqSE0Bvon4NQAX5nSA0zt0Q8oOrTrFgyyqX1TNdetHoFcKNv8gbOt9Eey2E2EW6g
XC6wasi/xw1lmfRq92nPERUtlKpKVanLDmyvQoWR+z6onoumVuABIkkXhhpbCdyxMn7ZB+4lzoX/
VDR7wXflnIxH8odm4GUX4p9QlxlnTkq1zqkbWX7otz2u5Eb1Cj1FF7DX0IkCB4buj39VWhNDgLm2
cLjjpE22wKXyH63YBZzEBPyVyBnw1MK+2namChN/c3ZEJqO9qrGdQcoA8Kj+Ab5BiPvQ/T22trGa
UZTt7pK3el69y9myqIngNTRuA5e1eV84bq30mSln9BQvDdY5gbjwyna2vKzdROBjOcoliD5vwuBN
ey6YKHLy4ySa+Muy2BtwEP3QvellvuDs5fw43pcTn053ycpr0cOCZEvBHbwRIaYmi63pUuHLGEDn
17If/5p+caI2QO2GFJ1v+dRns44pPMH8zVVniflYOnAacTO8SQpkIHxxg46ozt+KaX1bDOc04iyS
FSfQzsT3wWYaazvYa/C+jWAM5XJWf8Icx8gore1pk2nwIyQEue2NEoJuNiNkxW2qlRaveZDDAgfb
un3KwClC+Q+CYwmndoejHbZQcPPDPVvXYiphTyPXzOgcZnE9EmtkhdRrKOGQ6DtM4oloViiybNu9
IaUsORA/F3lvnrRuyFEW8eRUpOpseA59x+/ZWIIg578NPPHSaz+a+WhKOVqfH+W87B77Pf+VXUYM
pmUEYUdARU90Lp45gnQ49StHfjn5sAuNZXjIZ95cz0MKmGqMRsbaqqvlNepQMSSFxlqPAfqVdHMQ
JJJ0bi0JDmlRm2YoL2hJzQ2aWXjlFucGsSxf2U7zzAIMRsiBqpHjgz0BHbXi5tnS4Qui+yF6UFMK
9hiC94B/H9c9IW0dIkIYRdqCeHfjOFDDWnASPJVyegT5AHKil0Fp1oang62WVA7CNXrwvWwkmxIS
9lqQVbitSPnQXqI/jx0vWsnCC8xs1u4KL7zEnZaGGAqoMjo8IDJbEybzC22/1KxoaYzsOfNjDwOV
7XF9s7Tx5YuopmO9Q21ZKplzUso5E5Gs/0ikNaVHaMY0BIZTzuf0fwqRde+k6PNBzLuVpMKBvvIs
vt45UQPoi7sjP6UoiCihI8iE5L8lTc+WxpqsZFqWrZ/HZRjkNXZ4ep50w7vh9bvGyRNyV2DVBJpz
f2J02ImSBkLfD+mWjjt12Sqp41adWldWaqbssb5v/GWYf29DUvZpCtcOefhXZBTOoxEylh6uP7XW
rnwClXJ7n2flEazjXo1tMPjexrrJu0TvVVBmwhtAvDPc8FNGtyeZ7uO4OPMnpkCNi1cbm2Lqzg3S
XJ18eNM5UQ4ZX3pNaKWvAe9bPqCNQw9WikOFVxxbOQlC5ybFiSDB/fslxv16t9bYJmZyx7H2S8N2
LgJbZpkvhgPsGLebbbg56ssKnFWw5Yj+c5o2yPmUOMbk38mtcpcTPlPFUkMxg7ztLgnTpePLY6hl
L55hSRbGWtIbg1nk/hFaFKS1yoCpmUlpEhJq6swYstOMlrILMpIxdJEmFHtUJOGfmoFhpoNDKPCo
PIo6mWDeljnNQ6mEkKqZL16g1tacAMeA0mCBN70AxtQzOpZ9LM0nY1PLDmL5dl8qD3xOQdvPLgjO
ditgaXZYOTAndRjxDqf6wC4LdkYVpgZotOEDD1LlOLHKr9uXYCkjsTOyMsLX7NPiGb2pfWhgmbJt
YI8Wxe3jkbX+JYO1wD6ktg/dliumhIHHos9WgJRMqiSpTr6rY6EGJIGng9atHO/LYfUCpBXiUCkj
f5Uf7lbtyuC6togAHMhDh/4rTrk2irPP4k5J6e5feddLoxZqgJGTYrwwHunKq2JKtJ7JdUOQGN0c
M/Fj0kMd9ru8xUMSYi9cmIgVbiLbNMI/CW2GmYcm2OoDqm6VXRKYM6t3g/v1CCcVeJIxZlRm3R4W
WEGmsvky2QYXDcEl17Yt+Ydz2tr4EJs5zMeR9H33wGv6ocHWAXwGgOj6zQWzliT0t6Q7AO1E0eNQ
0HMeFNixD19/6BaWxI9YrFb3lbTEjFp8DAh/C5Zb4THKpZk4rUHvgmS7IuQ0ifbEp+Eu9y9/3AIs
rpXRAx1Je9SgppE5q3Wlt5E94azXfB0/b/FMeE7RchkFgG4tuKluGnw3bw0JhE/8scRqACLw4oMn
YxarcBBR4O4DfWI81NPCrvRFUO2WoD9YLBK3n7E/qsB5FV+x6wDmr8T2d1JngNck1rGB5zINpBP2
9me+scqyJezN5HSMoIqbmvJqlrYtWvDN1Xn6fYWe9hnYY2o/U1GWuNggxvJo95X//NaYZEtNZBgv
7tuBiwKZejinyTQ35aiCNgQkJBaLtTUJzEQXkWlIOld2tLv+V1NfD6olcALCyR8LalpgTOxKjLIn
7ET/PEZYOQERxa4IblzBV1cKT16Oo4h/r0FRyNy0RHzzM7E1DKMQm6f0+ykiA/Y5+bM=
`protect end_protected

