

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Pb7E+qNVEP4sE5d3TkwQJMYKTR/FjAPrexB6qdDJcLdscPV5w27UvNCqw/kg86JgS2hNrfoEvTNF
uJ9eNTpy4Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Egq1eCtVuCp02bpffloqFi7UMw6fphk3UOZCcejhe9NQNeC0Z0b1+S1NY8yEfAVY74l4oz8pZ1vA
hbrAzplanZae/BDY57rCQ6UjD8G9keaOwYv6mG13f+m77D7Y1nVpXOE4Uujw3cZ1QgwXR1H4YfYp
ysjb+lxmo0pqYRikRIQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KJqrZ5TKkbTlecBRrKRCsxKhAd1omWJvIin7DNafgTE5a5N2or7GsTSawdWWjYWHESLBvStvRGQE
jVUeK8m63dYVJN98fa8T9iAHTDt9yiBRki/VqfvAejvDOEI+l8row+LhhHMvCd29xmkCeQKiq4Qt
hsdsz+jNufnCYY4Y1CVO/4preMZeG5Ow85vRd/341CoWEOBji8o4pk0XyIttBBgjBzWO8JyhLpza
R+Z8LgFoZ5OTfgpyTJ4SjYRWp9IHP2HL9TShNo3PmM36nFNBvQSLoEjLgk4+rUr657++ugJH31/C
Y/QScvwJcbqMK15awb6twj42y2gxJSFzAPzSGg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KxmYEF19quU2lnDIx1hLVbiBV1iU7MlwBSbpQKNAVv6HLtZNpIjv2UPtz6sPs9Xac0T26s1Kjo2c
fAw+uaSeKdgWE1BMMV8ya3nIO40+wJlyaPYGp3qW9dt6kM+FZZl/3MCpgIMx24FXg4CPHrHNKu54
/3DZJ7o9x/QjyM8WSeM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n4InNydlMoO1IH7Kq1VdB5tuRxM6d++erhleefbfKU7rQGdfSjRtqcQ+h67LKfA/jQJYdDdZMjd3
Jp84+E2i9v4ovZP9CPOifgPGXKRtOz0XzimXarAjLF+OJp3As1WqoTrPJI1DspdbqtDWx5caLezn
hcZVfRSFpZUoLc9H0HW6DXtxAWvJT8e4ntjJYO6koEzzHlZPpMhXvbbH/rbArm4iRGWLOVN205Pq
oJcFHv1n/e24XGuCRksBqssUXd+D0UgsxKn8Hy5kQi4Q8xdFEXxEOVBI7ivvG+HKnJFOOr+UNhLY
+rNFOKSwlDtT8tPfpzjKS5GdaTuv7j2GVoF5Tw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21824)
`protect data_block
N6VjYkwYKj2mWI8n0VIOOYn8MzKpN86HzrtqO1fATrvSWtm4BNNk6rBTck9uGkORXzq4I3wZVqV4
hfmuwYiihb+QbqmCbh8pzihS1v1bEycZ5W1T1xmvBgLjG040oP/F7w2tUywhSm4dUT/L8h5kfVvk
3NyqOiC20s7Yn8Ei6RDSZVJuuyycACB43AEqyJf/ZNDFDI01OPsM+bzDNSvn+KKEHt7Ccdlu9/pU
8aCBgeKEZ68/aP3gUkAk8zp8oncOLJK1yOgpmF8Mm4KjxoUWcvY4QyC4zfUr0nzN1eFFVO6ERdWY
qKaEngamJM+DbGfChTtrm3Mm4Fbgi67zW2dCeFCWppqTovakWyuH0NoooyEIZB1oTOf4SjHLWl8S
wabcteV9PUn7eMJ1KDhET/DycxigiCGcufR5StO9MaB1ybWCK10TdeCbqMB9EsfSdzmOrxgpWbmt
Lz+aLp0izDs/rTxHyFyPnRHl51fgOb9pxhTynjya5ex9Bru7amdbLDwlf/nTdtWpLzg0sxiafJGo
gONrXh8DmEseqK4Barp4RRLfXIwI5HWjtA38j+b7w+E3lYZ683REwHaZwZThx1QIc8nJSjHu7uSz
wumww9lJMyZU5fjXuuCmY10E9mYKbZ2R1kBV23ph/dYBTAGrUzKi//DjD5ZnYELqgLsUFq5WzxRN
UEyk/5hkmtCi03iwWyQlkwHlSHT/RxrYa7fUp2/yJAh+7bRIS9AtFBZn3u3xU/Z+QofNurCP9R4Q
fzfdG/C131NV2VKJMYrnxBCghWW+/3tAnl3kUw9WC8fo+meh2qbgZuX34BGfzEcelBJm7kvSy9pi
CjblEIxY5Xy27hgiEhFXDXoXNSNZ1X9Sd/WZg3ALgiafwwMVXpd8cVTL0GjBVlnfrc3uWTZHSPTg
qLM/18rOf315bud+/14LXN7TbtBXkijiWeZj7K9F5WAdlA0kts1SGWrGF+GoCgCR8sPbSl77bxfd
fWOkQBi1eN180Smtt8sw0X6CARGPAIdAKSHUNgf4I3JrmkqPLljpueral86qQs8trbOVFfFKtrsi
K4AnU4Qe1uXcKSaiOgypTsNWkiahgI7X279WBfgXC8TWlH+A/q8KlthtNieJcLRUYtbbSVj8KZ5H
gwFEB0FBE3xOVssfQvOQUQsdLyGnJHxRPVZkL4g5yVP3sphKaWWXfqV2LuIoUs2V6WRrMHGlHXo3
+NpqkeOSxduGAVZ/7/WkxUmclpQqFtcA0ana4Vw3MO4HYwPmGZN3y50L+eg432TPLLDq28BNMSU/
7cI3ddEhibTOPqc5OMOqLzCXXQyGnNfGICe3FiDxXEHSGAcpYKO2xPJ2DsAcaLhyKjkpZJsfXGOW
PVYIIjRnpjAVfBX2cylCcajH/Bm+QpLOD9OzWD+Y6ikw9n9/WvGTXHTPRsDEitf4XwGykn16Wrum
gLzM2JhjAYKhgTG3ROqZwcokXFDZd776rTtwv7tmAeOEGSEPRWHZvlINA3SnCUYG1hbyju0zR422
bS3hbNQfAD0JyEhh5q8GIRaZLpQRVudzCzybIUpm8YGdJSHitIM2YPGu5x6lea/OVD4gMK4WlQo7
Gpl8w2aGK9wiDuUoFoyLjsvn72HUVzuNRE1lVg8r4qKSRRZi7lDOP/ALpsgABTpBvktGDprjdsec
rKQ0aqOPEv61lWjWp53blE0wD+aD+6wKNFIEo6S9wulnTR2uVwa2w8Rc1R18N6sxlhfpk1Mqa992
6R39FvIe3BY8HQO59pdyEyEu72J6Ondh9+3lXa7gPVITDPS8gzAxXWcil15dq6X8GXQ6WEl+8PJT
tV0Yj6Ms5fcZW9khnAkBu8sKq4UQUzH2J+Hvh/z3WklUEMHPSZRTLcpiJnm5HvCGmHx6tMAyLymY
dYqw5DYV+PvID9y2mqvwn3rpki2FpjnuCmFNR5aNCUO9deMrWARbhpMQRhpmAHcJVO0myhhkBOPc
EReDmB5erB5O/UJO/UE0u+bMszzpNw2tbZNLvnsS2tahniPgAZvzZCdaj98JVxGysrERkzwamfJ6
AiJpTU1H3D6ivNJALQvfyvunsZEUffVhZ7+4WkosWM3oe6OG5EEOH0M8p64YLym43DiR71mZBPpM
8sUNiPNvP3VGUq8dgfjWod1G9XAKLVKgYplviksmM2K27fJvYdfNcNAk2xjvvasOb3myKHGusa3R
tgoEtcgx7gnp1tF4ANITjNOUp6+CPLmvmXM2wr5IMXk+1YmWvxZJ+4Z0pBYCN0NkEpJC2M6RJqnR
OwSTjoKaHcoj22Tpsc6yNZCdKqCx3zzDfWaHZwvE3r+IPifhnlqNRrtC53bwmhbfST+v/2mak6k2
/mzuEr9SMAVheV2Muv8U/o5q0FsniyURLoJ3I6CQxhYYbRkr+Piv5qwD4W4rHv/gZi8GlVqTo++8
v5mk+325CXpe7MM96ql2+9DA9hgshn3pucx6AzrmmXiexc9xUnwE8HI3oB3b403oYXjlGHDbzYe5
dXzzll7AXsNgcLFADC9ivHzAeN+UEfx52846bRX1tfPdTk7DHOehKya/cTrZalb+7TiQ9WY4IJlx
KoqbO2vtddcJDvK+l4wqUR6YJ1n4azRbhVj8+tba4QF+gOI/XGF2tXZE1rCT2BfTfD6scPdAZ5yP
2F4NQhZM40IqrmMLjXnpARmY/gF0w4p6rlmTJVUxT3fOfcIDD6M37tFsNCJCa+fcXAYlwzy/LmoL
c6TregnV4L66lqNGBYfSMr6kJlUb2MEvFmrYHcztkSKyece0c4yBtoxshz+9BfnZz+vMnngnp+vT
qDda/3i3w671cnnv5Vj4CeeWngdg+Xsu+8LXbtcQFDJJRHs7ioupHFN528bdcNPcRBKghs7WT46f
5qnIu+zYodS11q1XsljEDh4ezVNf2bBbEX0xZbfLvkWVFtH3VkW8EVv2g76xdnCOGwPM7wh7M2el
iO1rMlxNqv/A9xmsc3gwb1aP8yg9itnmPQ9M4AtrwSbi7BrMG6ZHbTZ/kQjwzDKRKJCnrqYShyfi
rCZsRk6DboEb9SOYl6dz3DrKN0c/xvsQnoN2/UrMCdlFD2G3+u3NYP1wzizp+xWP18XwZmbKrruZ
D9OR1wlzXNJyPnqUm8BVvm+EIu7SUGtQtZdOUjEOiWSRTkK3kjHBqeNI7HcGcJNcx8uRRQLrig+t
Z0vhNLBjVRn2HoCITzc+Go8VGEYE7acystVm/yIkc5QeoWXgd8idZoDWRRdYKZOpsWRPLlDbi4AB
Ld2bYrKZAUrQlQCCPVhBwNKidjZ2+m92cJ5P6q0FeM0+Ivd2RbYYLOcjNucJCfOgpgz5g1d4pqZF
fX5FbuJkQeiNIKjIe8pUym8M9jss5DftDzLYa9YcmadEfZf/yqGH7qwry0lPeFif9EDG+m5D/GG3
f72MDrl5J2z9oZFjZDvuiEU1d6GND8K2drLZVOSoaXPJYd/kyG6vNssTKxXMcNg5eQ1JdljEcosm
gGGaLWSMbPhAYuH2QBEVEn0kAB1hlYE6/nGpLXqtrFRRdQkzQ+nednDpWq5RqfuZibRv721kO0uj
7mYLc01bF9gfcOiLN5GyoNRP10htsMJEL5OxWW1NxbW+Qu4mw5QM800SlqauggfuVXWWiLOqKP9G
6nx8HiNyO7qLSqwWIo1RDF47pNMgyLnku/oAAXdLuBYuBoLPr1DkzohodmGGmbZtYujlEvb4BPUB
Db+LfympwLGThIZo77SN+bEKvwu1a3+zlxP38u028ajEEXstbFb+oT8ozBokvMY8NgAlad/K3n/N
siYDqZvhbmqB1dNAHbjzeUKgsHTycwNVaPFRQFXbUy0eaKH2lpcn6XuCBudHaCWU+/fQLmHXiZM1
EEbufIVu6YDumCkwqfqxuMGLAN5VcMPCzx3E5J7iqxkYIgJPfN4YRh5zb/pZiXS3V0/3+iPssI/W
Bsis2RiyNThb17U+hvuZEd4s69hzyZ+OZEZbp6+p3/wDnGfqRQEIzpp0MTnpG/dwcjiz18OM5TDB
BM7h/eWRbbwHtgpLctUGhJOCalRHbOgCbs1JzRoCZZXxaPETl2ZviQIvx6WMXvm5FrDDMXs/O3YZ
GerfpmBCxcg/2VDqmzkOB39qdHJa+d6a2PyQ/BpZGHpt0X4NoGaP4Jsu1XMnQND3JTccJ7E70Mvm
3Qp1mgpizNkFS3F8fljU67ZDOkITbeNpbKPZaZuWWLv9NSdGPCHpdRVFNw7OU2hxUr2xkJiBBjrX
t/w2LGRS81my7bqX2Oph6oCDI3ultWM2bwIGpApWdtuh0cPzneZuZYGi68+7zxokwWh6sfdJvWxP
gR9WiN0ONulNUzKAqzGhbqAJ72YriHJLfz2330Gz+CrvTJJHwtRUS8g0XaYwX/UvnW9yGU4CE023
bqS2oxJEoBMNSp6nVAImjZhy4DPEYUIfAHJ6OEN+mdO6XpbJ5H0WWaX2cNbpRccUulgIi8NBQ7aB
s4NG4+CjO+Ovp1DSsTEuAR9zoCp96Ji2nutObFwd3XzzpyFt2VgA6IAyZ2EwIgoUgn2qTT/laqqJ
DoUWVELeqQWxLYa44UA7DUEyKRLErbHfj0mDxF/dWOd2TkuiOMirNIG/NnafR+oH0XpfFrDbHbVk
C6iOh2LWeUlPmxJUrZAdsK5q9tFwQpLvWU1IzWCbJUueJrYLgRWdZPJmHVK91B0QY38o3hcoTbzv
6SegFqDhh9qo6bbZ3R8CpnoRT6Rr54dVWn7NcTSYMz7e12k6eRH+jchTt585Sxo+dSl0kTV+wSty
7T4HFAM26fp0sSeBhRmbZU3P8MnHmpVU0sKu2KhbYukNQHdEyezR+5H7VUTcTdzoWxczwxtfCMtH
0kghs/amqrdkCisnCUU6bB4KfyfnP6rWhU24v9MNsgpHtYmSb1ljhbEti7q7cSn+NRwLYXQzYyn8
WLl6ge9ccC4pX+RdTCQ8qfLXBtWLs+lXMhGQicpJYDCUm5le0osu/IGRgXbFpcuISHykA7Cy35/g
KtrMU1SAILGYn+KLBFjwYwhfSiMpnJCYZkyUzqQcetXK4/AnalXeUa/KUbfYjuP9ma9xT9gygSyo
iyUsV2TTPHMlAxp7iqlL0ZoigVQYP+p74QVWhJB3EhBmKgMqrSvbVV99d+7PfI26LRCzYwv2q2Kh
iw6FBcfUy9jHX9/5oS8TE6daLbUOPaPzpjUlty7MNf/8a2PZNOYlozJczW8ZxcSWrVMaXSN3a0BE
F+r18by9eYT+sc3MhqZ2ucdaPwwCOn3F1l4nE73KB2d5IbZRD5s80JbeDmZaFnHMVW8qrQzymL45
GKmcfLk+TDWP9ed0h6EG2b5sKj1ba3//G/E+K3aUjx8Nq08d698t8QQFD1434vedu1vIrY2Nhf4o
rIkotIKYKjPlSiwS8hvM/liu2JIcsHSY+tITXFG3hI1SuNBHVmNJwgiKVfplYY0P3uCoIGEUvP6D
hJEy14srl2aSfW9LrkXl2UT3UTLFNdhGm23Hj8zV1i4KKrv6v8hXbdNAniJ4ndBmOOlrs2hldQtP
UPNkcPDtGbskkFsP1vRG29/LF2Q8mne21w3KrycRMH8ogdHZJbmRx+L0INHbM1Hf2qyJZoxNXuKE
9pcNQlfb5MVFQmDWIeM1SYnMiNWB9Deo1O7JB3GNKl4P4sN5cZI+vvGbKNMTLoFkxoAGPcMiKIh/
7DxRldJKYhEb0YWlOrA4hcC2BkRa2L9NxgHNMp4joQQFjRAGKerB7X4qkg+W5JVokb5Rk4VxomY0
bPyQqYFVAAk4Hl/f6YAeUexT8OgwU+lqjr17aa+3DjTl/V+52Ls0WkJFC0RpjTg3yGFiRSC2ax54
qde3eDEljQHdtuiWFmLOsKbbeTAq+0THRru10D9xztntEw0yTTHrbRJVNI+0fGxusHGa5azI7lyj
ZrgbG6fV73D1n9NT8b030/jt9RWQDjTMYPjlQB9HHL0BHDKyx7/1BSP3SqATW8gKHIR6lOHrs+cb
TQ2r4Xlyr3I4liuQ0Vh1duuzcE8FyRIltCd06Wu5dJ68mgOlAj+koSMjk04PCgLEFGDpC57zG7Nr
azyDJtgiVngMqQoGWoOuuVNzIXyzuEtVG1/PNtIZ/5RwxBJ7arWWy5Rgt5zS8402WFzkrQ5kSNeg
lfzK9dKToGRzrExzVnpexUH25P4zmFw5ZXmmVVioZdxB9Nz67HCfSFuWwrp+JRYW4ST0q0NM177H
vtWYdso/ARWAw7e8vzsR2QKnKC5XneHctdsH5RiHXkRnoB7CIpqVAz5VgiogOBHCHw71OIDlxu0+
vT9NasXHfDCN9h2xLKtRJJ6ATkuQ6YUP9XVgYHsvtk/toa3slFQLWghhzRgq2yg/1aCRXT5oGdBT
GmSPBGRP/yCy2veFxntRXyAQZAD3WrrV6L44gLDXu1sjrW3quY9PhuPmb95ZKrJYMyLDVamhRerF
pIBFjPJh1xDXaGeKBZoaidmnuS90xS78btpz1fsSKAOf9UAmjL+CrfaBPbjnrBX85/BXmnSjoH3g
k2tyN7UjIM9qiDUyyOpu3lX49LI+P8uPFvy3PbEsK9kLt0xGW7lTu83XYtS5q7wzjnZVEbEi/Mee
G3XDq3tCoxTdXShmBrgGNMzh7K9etQjTvpF1S7rVKH6EDP4vAGMuoHkcSREpfYT4CyBU8RkjNSh+
1pz367EPgLqdG8bK7btMDWust8YSa9dVdcNoYZIAhT9He85L5Bw4OG5rnsdEc5XYMMSS+H/q8lBb
6bQaCm779Hu7H7Zyi3NsbS0xPgWgKiT7NXjj6UKjtH3miwU5n0PP5KjMcCGVp8YidAhn2lJTt+dy
/1nMCuv6ed3juwvskDifB1hNDPjKcKSqXbWTSCQjAGo1YY4bOVBxftl9lQusOulSHDSn1AcD+mRK
mTlA3ghqnDtOC0CButKEZI62koiVHW3KnNK264FCe0kjZ8ViR5R0m1aO5qEGUq+VKUUq79pOqaTY
VUuRTwqE4rCSK3LWwxu5ou5OatrVMklJnZg3YRPvun2C3Vb0wJwy4I7YXErQCU5izZx8Km1laLWS
1YwWAl0Fl9xQsSLEfTwPsJdU6izgWU2V+AWcbNa1j0xhBktMUlTmw6GpHKuUwFivihA5UL+DfGZT
a80auvI6TqCiBkmSQ7yKV1j6KzKxj1nt4VvOPG/zE/CHTQhk/sIs5iHxT8OvaHCugJASY6Msxbb4
oFkO1CXHH6hKRbKUOn+C9uw60XN7QYOGM8o8FBshwklBsdIder1kSt6d0X2J07YJVTjovoPozSNY
ItCGIFZhtvdpPtzLTPVO6k6L44cTKfsEkIpRCkOp911YYMfyzcGQZ+Jc25MLUqP5j8phx78U+JpI
ZfEXl8ULvv94x1NzZwyHZ/RTrbrG9snMCBLg+f4xRg8lb4KOrzlWcHYQ6x4T7+gWJI/dJJhCCHl0
rfmcEHAFi85ubZEgQCezpIhY1p+n5ehyzhYIPLh22d8GQatC5d6hA46HDspnGiygIOcQFDxyKnWY
zrdlcxApsCevZrXQ8RxtkIq1BMq7+yQeqObxj1EdPrFALg4B8moOagBWkiwQSyDo2xkS44DKYd7O
h+loxHtn3/w/TBiuxrraTSYpJ9A10maR5MP5z5FAwGdHA714EBK2Bpav1xRJDm6gieMwbry9JSSs
UMJ9cd2RYA9pOFFqYig1GND5XZFWOO4xcRUjB3amAigYpsJDWIGSTrVBUtroIz5k7bYYpqb8cjtH
a/bXaMsXuKRvo+RTMzOEyUrl/3j0RAgKwL5HAq4ipDoNBzWlzBxXkOaazpqUsmmFZHyP/iAUAXMc
SqD1s8Ds5Vgh5X1AtynpdPX2bwQk2IDJ49T5qusOiMOolIigR7XeLK/dH5OKGd0NAZKxv3mgBaDY
BrPvLC9ZDOkt5rmUO8f3Ov2iI4IhFYOqpIHVJdMBQFjlSHWmK2Tl9ueOrTq91jrfnst+yUmWE5/9
5c9TOrOGQj/1kOr+OzhHYLA3CVSmf/VLnGNo7VqE7R0LoNSfE8npk9oK7Q1ZPKkJHnYARDgZEcKp
oM+g+GIBTiSIYDOXTI2YH3tNVRj9DnmMMGprVMFzfX3PeZboSm7iEaReCZ30ZGCxXDDBDqWhQGHk
cbYNd71pptOqwh4UbJkc07r1dBawhMJMgzLlSdnAhNdCjmgzwfl6WLvTduseLYtomSud6A6tPFMc
c4Kq+Y8n62D8xeFhgxUjxTpRWBKmio8ce5Rxmz2FtrA4qoWMSOWFuNhBIv6QfZygvVSXohS4KSqh
DLjQW3nQArcvYX4Aynh1LbSvWfX99yqyOc7JmufURY7MT5zcHj/GrsUl4gVGiTCuFGTUWlyul4Kv
B23Jvc0qVZ9v9yDvhySMA6NbXjEOfo7DsIko8rC2XNdEnLnQOcUnl0foRAVvtQLL8rnQMkGwvAMw
KzklUZtKujSIMtcOw2BQ+dbG5hMkUBZwgy8im2kfprmqo/c0mXePwn3hI2AB9+smJ9BFhoWnqD9B
OGOg4fTbnXEplRZjEBA0ONOUuYSGiSSY0iX67diumTCVz8DDMKp5hmK4tiH8iEzTtZ+6R2tS7WZn
7dZhv6nmmlzzj9R8KpOsmrBaWYn30ilQY4wUnGzDL+Il56to0aLrtw4N9Y41yPIMmsJ1QKO4vKmA
SMxbX/8KJ9YHd629HIYpRnRu7nLuQbP+uMtDeOhsZs8L1FRgb0E3Edrv9gwPOWAvI/mKsm/SxIog
ride09LMTRaMWz8Oq5+rfnWmTDK8ZQuU6HnHb7brMI7zIyozzZfm+5wRxDqenrMq6u9EFrwLEuOm
0gdicxj69RuzqNPMZzPGpv1RChr9hbdZXAef4mX0fNBB7wJ7c+SSatZCon3awkZ2OReut1coM0MS
nAcZWsygDvlizwVi4eqhr8HFz6v+SaqrebjmNWPI7nGB0vsaGZw1ILYfJ9YW/4khsYip6+XTV9fa
TQZkomrGHZqkxr6viA0vt0T5LOx57bBspTOt6q9tjnRPiWJpJu4ZjlIQ+yMR05YsN8kNJQRynCrr
5QVyDLC+EcxFOQp1Dy+fv4MqlYTjJy9gIvXVSPjxsMIwbx/EeyBz2x+Mygb95iAlMD0dA4ux06Li
MTFxYpufj0IxIP/p0I3yNr3N7emH+3y4vzDeDOtOl48Ubp9+0retr6XgRY41A+G8Ah2G66NufsyP
GNCx+let9QHrcfQv66LnzJirQOsz1sIe9AkZxPJiSGB0MgET68tBQlUq3uuEt3gEWMvXMomGcfTN
tKpJulYZ1xS7Tk8fjPtmj7WpekJmQkZd5aCGR3J/CBbzyEtIwOf7+BvMd6zxK6TxfLAHdBXJiIeC
u0o91G++VY9hivyTDWmshmLlkEH3CFRyzeU/f2t9BEG6U+9Bo3XPGykYpJA1Uvk1t7zcrFgn4XS/
rx5MfJa3KFB52JjHYq/MvrT8WvZoeDV8CuLsB1lrltWMP4bB5slXEpGV6r+bccWW62/AGM4ZwngD
/3uZwB3QY7ggFiVxUnX4MGJu279a0rEj7oAiNZ8LlWgCC7gosw15mpv0+msKmIWR8stzTtrQnd97
OJ3rBGBGjImkQju1NF/f/UnRrHevWZv2R847lsKCHvyMqvzEJtrHMeL8T5a0iufknBt5y/zgjlhF
VdV4jDUSAMS2B+hkjfiCA7R9lhLE9vZ21lie2PBCjcxCXXs47ZAbN9jgKgVsVnJvDu1DsxdJTrH4
rgaejFwuWguaA9OiL53Vrl5xCeDTCZqIHshvY4d52CoyUYOWVYHprzKBhgGoUU0zTT6OcgyJGI1x
Ifq8AvJ0pTATQlXqXOynsGUAFQvkkme428oWb+AdI7RJJoX/O2f4SkjwGaxrCtwjLEI+Bt6c/K85
avsaevVOFOnWNvlzhIKS3XlEnj9Iiudp251gQMwyZ6ON5QgDI5hZRPQidISd5rU+2CkK5ilIhMHS
QWEyC5u/2Emro7l/cgq1YJ7l5jrRiHWc/3PAC+9Sv8dSQ6jMxGURwDgADf6/VjJtsACpunu+CuSc
JVw6WyOcX3H8OT6WsaHGCRe9wgT9nJAYwRBq2kbMaP9QEFuKyaGcgcC9x78LXVvTMI9U944ICYBH
2vgcgPhPzK6OpCyyMn+Md7YfdBIBwz3zHOgDl3WJmsqLZfvREyNty/yI1ipDiPo9mokGSiazf30i
qwvBrfV3DqN4gN7IB+KuI92l3udGFuDrX959SmWF9v/35H2hcUffLcV572XH+HbmI/m167srTH6m
sV0dqaIWFgJNYGCsA1yx4d82zULPOkDm7myNnlhMKQ43xxRXnFDXT33MeP9Eni4AN5+a6/i7+Lk3
2dS+8ek5fN5qYh7Ro6HTeGLbgLTqX2DAS2bj5LaTSHdAy7+tODmpv55euwzcau7ApuRXEORN+z2A
gm+m5q1xs2v+CAhcnk9Gm9MF03QvO7OvTtYOdo/JiKRuVn+OJ+jMPoCKD/tWJiPv36m7CoJe01uc
VsQOsrZ83LYLTIuxMh9RN7SBl2pjFRvGmc/zk6XorJKZvInVnWtcOP5kXX4uAQ4nI52ZBtzYlKyJ
xwYEcWvsZCxzfNzAISUHLBVtJF3YeizxpNH8dBJhF2jDFiAmWPuBNaZ4hD+EZ9Bj+li3pGM84Bbh
zz3q+HunFhitSSrQlDkRtyhbFeNwIi0ifS8GUf5xvTXaE+bdnU1F2MEz6AlVRLSKAbbbutCCfvkZ
rQnJ6ou3UtruIhQxngOqLqQLjXnAZxYEYLZYFb1w4vemQLgGtwOeNNoS0Tb/dWrSTd7fcVcKlPd/
db/J1Fn581Oq8zHjdO6PIKhNZ9sQLlxos+DZr4gJhdD8RCDOcbYcf/5DbUyqNd09BinL8yyUUw0G
WH7DjJmU7TxJoz6N5r7ePyeITIgpH71jyiIe87cO/9myTtqn3uAdyWK8NEfatDQgg6vQVDeTMfMf
MmhAf1Lu9+EmZlJMwWZ6uS2VolkFjz7AujOSTG5x6VY8Edc1ZIPZ0CSH6RkaXJl3tPXRQmWrCIpY
xChQzSUcCqWqMNx+p5540/IYtRjw5l9H4zeavOF/HPfRhiOVU5eton/Q+XFigNWk/lPDSP1ip3GN
QkV2uoIS+CETc5j2olmRuw+UrWirk9rXxf7FqoTpdQIMla7aYV8onXP2yx9EAANRGO+HgADNFzGS
Uo7e/CJsOYOZ6VjZCof/qjbWePEtgWINWjDCW5xMN8XNt2NM/MfKrtVvQGaIfX7z7EUoZZ+E4MOP
p2y8lqWZo6NgKMJRmBiNCgbTgPxKkYliOv67C/Nhk6dNNrSgo3S93KLJqO9qWm2DEl1Sz9QEbJL+
obUm3Ec5iVR5m3zKTucHdFAeJQsFnjgp0kjRghyWULt+S5YCMR46OdOubSpX5AEOSBWLCWnPtDvr
+rvUoMcvwkm1JYYJptVvAA3j3SgadN9vtcvixLT9M+0T6JzaGkGvHjqmz2QpgEjEgdVZ2dLyoNE9
kvJ7QkyOy2uUWjlEDuBwXCrVDyaybN+7wVrKo/uRC6JDdq0qd5uOo+SP4h222I8KUQn+SxLZbVro
az9pcbloFTRS3886iusVIaSyBRqUjIMsWwwuOF3Trt7N94z/J0sJB8C364mxmhkDi4Nc0dW8kyHC
gowExgGgJ9ifh4JzaUKqLbN8xsLwldIxpmOfCPJzTPcKh9G6unANhY5smz1EAHVHmCuJOb12ryLM
AFt5BKUA3uoDbKUBypIWQe1CWm/h3mfyHoLfS73VFlNr6T+DPEvVVOrGBLdBZnt6g+Di6GEpujA/
RQafafRxiYHE4TtVuogANBZ4r9o+tvpokYMLCMc34kE1rHZ59G4jqTmwwC6mTLv6Uchl0g8jrIDz
o0QRRQsrQPG14Euute5wI7WBDztJ3KsqrgvgSUboIgJ80Avctt2MlNRRJ7UMYFzNKpfqo0i1/OT+
xhbWPMyzOG0Qt63qpPJGwNOtJWmKey3NAvAhvgvWD/2iSPpVudgnyMCX5YfGRO47WfC+2mlzg0sN
NVcRcED92KiEeDL+N+XWEqpRibwQGYMASXFtKQ12P9tNEzWsItRoSjJhz6hubf1KLM5blDEK90yS
zlYwfbE1onAlaqD3nohmpaAg9fqq/sKRTFVCsohe9olstm7pCSB2Leq1ApYFHNv6SGMdVbcM4TtU
K/94s7i/LP3LaxbzDhzJQSU7QuX0n1+nvnpJG9mUrPtJtdY3og4rb780Xq1Pi6UmKlqHX+yhT4WN
H7v1RIk4+KbmReedjIjy8c+dGsfFRZpl8dufKrB5NXDU1sgqtXdKmyovQJy0AwoEQt9EKj3NhLRQ
ZvXoawxSByW+k9peLmRiJM2/lF22TJx+MrNniNlnRAinzHTbIJfvf2YUKyYo5VcDmK+mmhbfM/mb
mv41/Pfm/8RlhfKL/myfH6fr9YaazDQHm71WHEHESRK0+hX8KFVqF7VtvqnHbfhamT+VLKnBrXpG
vBkMyRhArz9ZjAf1n40Agx2gp7NrGDMAdBOjwQrVuSUD/KEXX7Eew9hyE8E5LzfcUKO7wokGnZ3G
hGBPtMCal5RbllOHWT/nd8Xel9T5WnOrwsqC82HVn1Q59GokkYq18WQ/sGm1Tenu+LkhFygHyF2O
w2quApt9yNZIl0vGvEV+JU90uDO+zb06Tr3BxvQobImUIL0rKo3zNmoJfQoF8x21FxAlZwmhx16U
ga2OZ7wEFtE39q0o5ScMCucAihd0Hh5wg8qKrpDpPfh+R6O/VBXoS3/+vkzl/D/Byne4XMpyb0Yl
h8uK8J5BpleeMqyVcSDKHFkYCy+M60KzI49KZzj1ibrTtIDYP54pjBXUDiX1ekz00gTAPbpihBX2
sRxlV6aWnfa14ihMIoStKd7U/I9/B+66A89A2xV720dzIdlLCAM8NNtffXo6Gc50FMKxo4hln7HY
NgGoJv0AfhYWr22kb5eFhV7NsG60ixGGNj8njenyW9j6mvQKBoHJlGXX8K3Kwt5Midvkrvx50+YL
wtehkUbwSd4zgCC5agiTCTo4nZ8ACJMXb6g5QmtlfhjH8rDUH/jts9HRYuMKLa8XcgiEgXxlkk4m
Pyavr/XAx5r+gaBP4GDX8VjA6fDrkMxxM9sLC9W7DyHR/2p4//OR36Jl5N11521Kr1Y5pwg++dDK
WPcI+3flzsqB09Rf0G5vWFw5fm6GC0S4avra1nEzLBfpv7VgI5mJ/jRUEa532aWaeH9imfrh7vCe
Hm3P6cLoGwIxZr7Z4hU0urqQjCwQ0aJWoRybbPtE0Bq89QO2a275KApvCkAH1QYY+heyNxnFOKK1
3Z81LPZm4Gv/co0MuWdZC1xMLe9rsMUUPuGKwUBEaYBAkJlPZ1FnZSIyVAb9IdCyAo5cRquLgklE
afno8PL8b9LiexGdMDb0edpAVinv+tsdFB3sEenFXhaR57xM0FadijwKMMMYOwOD+qwwqVV4Y1a6
YWjXz+eo83EOTPhMGw/UbX/oPUC9tzoz4ABfty0BzPDRGVLGZojvIuprI1EMaYzTRwmz+feUIGkr
T8U6qNB3muUGt9R6nbeBxyLXxImyMPgUEhCulwLd9TNhV+LyJEcau7QaoW0HyweSD+sPKouSo/k5
7AfaBsI3C7Cw0pi62qSUc4UGrz7FdC8bXJg0mQujIAATUumA7PZXB3UAv7xoocqcIuOwsVdtIs2x
w5Nk5qwFirqEmz0DIalS4tKW3juRNfm95OILuA1yaDjRx6ZnDllRrBLlxvtuWvokZzXISqPExWZk
Hxwr8owsPFLvvC3iYG2bpYmLKlHcSpLQjtLJRt8ybjqhcEaSPKtkeNk/eJjTRcespj/KmxB7ksx3
CmysveLH2wuIGA1aUSSYn10P2iZCbW0705bq1RgmI1jk4/373bP0u/K4RAodGQw2+/j77MOzGAph
P8iaijhuMUWS3GozFa85/4gglR56+/8SjbpGKTsrLucnRlX19tkFuOHRlUPuC8ykklVjDTUxoip1
Deu+vt+8mhN1MsKw40qLE6osDjdS7wbB5YhS6aK26SAKNus1QyV5CFUj5/FDSAKw3gIcuwyn7Cpr
jWY+OUjWDwx3OME6PgYG9YxlTRHO5nKzYiX6guFkMMwcFR3C1jo5wtwzviHlhKhdUdm/thZtNx3x
ut4kSpaovzoaHp/s2JHBJ2iLXrZDxc5n7EeA86kKILJDVKhdwMnx89oq8O0NyO6QFAw8TlLIVjf1
25+Z2HPVjDu5nCqX+2eKNsn4wgLsAM6JHdKSCNtn3TXkw2eH+vanUMXGIkrODNqY7OBRcV8V8LhF
Z5piXzb9pV2AevC5KP1avgW2kopX7hPyRle0Amv4mZVcliHPWZwfjtbs+B36bfAYQqbD21NsjGhg
upDgXet7GsuXV4K+EirchSfgi8E3VzfV7TqxiAmlSIQxijVq4ZUV3zal8E6LifqhmaIJ+aWyzMAn
32wv+YGDwt3elnQ8RbnH4ZLGPbgZQIv3JBIkI2VGgcJgtln/k6aCcRnR9vsxvJ8LN5G0SwvydZz3
IqYvFZAQzkj9jAzgq6Z/LPAA24T92obWxvvygZ+kxTVwdbNcgeed0Myj9zEoVliHUwZDsAtMtvpk
crToQ8dUvTKbhXKsRsAt1x1dM2zyxarpTgLIvKIENgjKb8VQ+wYDZkfRw3j0fsRBv0hC/5XG2Tx/
fZkBmnF4xZKFcpHFxXXStPoPqCrSkq5xYKBmDm+BhXtEFKgVCFQIk0tmz7GCe+N/bKOK9TXG9wqx
yCTLQN9OFTALwfEuAvV/+xB/NlpxHfcrBOoQ69BjBAarynV33XIMJ/FzWzNFrumAS4JhZJlwiSXE
gWT5Ys+OQ/6wUkUFE5HmScAFYAUOLXAXiXjZFKJadJaixbuPurgqIIQ8klLfqf6GdxicEIzPiedl
fTMFh9Jio+uW0KE41cCyShy+FuIP5MNkUjqUdaz75x1Ru+XQ8WFqmWyXveR4DP1C/jFzwmZkYbcX
Xqk35VR+qNqLWUOUH8fz3Jz4I7nKXby9+2IQfg2u76QQwke9wahAXXCNNRk5Q5x9SniXjcvz7UVe
Za94LCvCQQiSNPkcP5XwSQ9tpP79NSuRnwJHE8fxmOG13LP5N3yRdV5x9tHdkiycJbXV4Nm7FVUg
l2nxc/AxLtEzY3YEI3vhjaup2dHvJN+XPDLpjhj/+v/taUsEnphh8Z5Tnw+79iTVCySI+JFVavNs
fd+oUUaOQKkQ9dFbOWH1+0uGX2cALf/6srxsvNXpC/33+8h9+bbS39i1i7Mvsxp+lID7ND6HYB8g
S0dRUOxWZ/aQuOLMChu8lInlKbn6vCXil22b7qmTRM/IA2z1r/cmhpgtw3vxBkoHSpQmlwUh0O4H
dC5jXC/Ot31otQv4+R+qM8E6sd1vOzHjCwPArum1Nd5rwLUYLe1l90UdCW3Tra5AfeEI227TuVHJ
Jo6DX82wIPbIxALz+9ygN1IaCs5TYK7cldJkx+WpUdHIH8gFWUJXyH+tfHuA+e8+d1LMaaWKQzSS
IYnlqS7aNCWaWyPdqJXyP4F4wSTaknM7RMIUvour7Mehe9JT9oBhO4OA2ae1QaViwv2/SxhCCgLZ
NEuNJyCQ3UG4V8la8m7UkOJ+KUay7nxftOEmbU4XtwomcIVOg++u+QhFkOhEuRvtD5vykB8EAAhn
PiebICMhPTNViJWnyUI9K1g+LtHtxlSlk3gMOLLIBv47kKXXJq8aMSU8pdT3aMqdnaMZQ1ayvFW2
fMa5GGKPgdeMRELhum55les9uZEa8+KFFTJwfU9M7MKHQnmPA8ae3md2ohpe9T1Ycs6FGdd2PrFB
fbSR2tnk+4/dqL1SjTWgZSgbur3JD1cpDw3Ba08eyd7LrR5KMl4XQWS0zgj0fJbUo8Why33nqCjZ
/knWmeESJFQVyT0qZN4UP3jDcRnAz7yt6FubmZ4gL1sHnEyJwS3Zhl4VggPC6utvEh7Z2Pq28f4X
eugdqr2dfEv/uG8Gl18gNVXlTccrP8jY3yRsGYMf5YtPS1kLDvkP8SiFVabTR7rvNi8AWb9pqXMK
0pB8enH05lm9m9sCOPGETgI38M00aegTeW8nS8AmGZpgZepv/kvBzosotmCIF6i09ukMsfpDqfbX
HtJVwpfOZx+aZ+QbXhZJ1pBI/cVYA6EURWHrxzVP1wMGQ9+2GOxv3R1KaK08IQ3FbsPUtyyRW9RL
PtBfjrTGsOukmlje2iv0FyjDGWhangn6X9jTEMHG/k1wL6I+ijEc7uaoEo0j5+5aUIKKWslsM3DT
2MVoir5IHzk79ycm2NhfMnM9nMln6VjtIfYZQ3Jlw6w881LAQZwIsSrsx64f+h4mI2ZGWPBPpHBS
gnZbm01b3Ny7PPelAFE+CVPEI7oO2m/AN/kA8cWlenknzldHXm4nMdKJEyaYFY3pEGyCDEQX93S7
qWuabfeIBFTQBMYBbd1V5Bu7gwyhRZrRNHdt45hwdATi1J3PJm8a09Gl1xEvfQ+HNSRefhqb9EPv
1eZRTtlwHB8Tu7RhTHSRQkBfjaEu/RKJSgMEAaqvbfCimbGzDZvqhFXyNh6WR8/syoLkLVHk6c+t
Lukcd/ueoz/iu8rKeSqSupSWYFMXTmJgYD7B9MT/DoGM1hnHMR1AS5Rw2KAuOohxqv4ISgnsHkft
3gmQW2sPTKntRZrxsD2xy2dfzSYrefOtyMSfNH725+qQnjjyY5zuG/B7vrpPSuhEaiIceL7EZzxE
coi5e5Iok2E2XgZwicxIFSTs/W1b5fsQ47yEj2HgYN18rvFEiKlxq/lbRp+BxiRlcvbCbr7N+i/p
w6l/zT3B680ubSvePL+lXJdrauV2hvAHJrHOc639acNpKq9tBip0XD2X/oBtrxWUaP2/cyi/bnAm
pThMf7o96kf06JmEdbHKILu1fQDoj22S14U167P75SGkxYQc5JRNm7nZ2Ez+PsOcxwxEGtv3pRl0
/rGojedvOzdgVlnrc/MoejoHt7o1OmfvJPw2PsVFe76auIIX9PjWtosPB7vzaMMKhPHrakF0D/AW
RJJLhbY4cjW/oqf7TvBxOM14djMf59qxJDtXuDEz5By60n6J1fZqwjBoU135YXODZuZjO/IaHgYG
tVRpgU99v1Zkm+sJEKEw3hRfV38dajVOOlXM6AUymFLSHuTefancfisDvcxhwNg9GNIhsu38kctd
yi+82b17hBiPcbLR8V/cxDieSP5guXqtfuOCLpieHrPkLqionYu8pYKkUVu+gHz6AVhNtzyOH9Do
aOLiIRIbUtyNfqDZl0PZZkptvFS7Xa4Z+JAuW+mSPsX6RAFmjYP/OBIRKVGLE4PFUWsMFPMDHZ/4
30Wq3Ljx1NGZeqnkgfjALI4pLEHCinxY3962Oh2aBkQZlf6n3Yr0ow5YmgUZenKeCtKZklxRhDj2
jAyKxtMaKE7m/YfWNB57K64D1yOOtd26KhsoYyQ4nM+dVL+LUEDtQD/Q9RElb/x8sQ+3lf9ZakYI
7TgHPF8fzBMm1YuXs/70traLJ9JN10SEpW8dou5KSf0zPe5up0zWNL2SI1QiGvqRg/6yBP+6sanE
bxkqruztISW1i4YP45y0JOM9AUB3ywJqtZ3a04bW1Ls/PhMKJNJU5mtJXQhj7uKy2cAtAx74twkr
JAhp6RTEY2J4pFVzAd4Vp75Qz0ek/3wSQvQuAyU53wsEMTcncwp0QY1MHyRf2XMPrKoT/1ANR+g4
lqj0YgcKfyZxZiFqvtzKKjsoNmtHtwrXmVf6+xVk13317rt8hSf6+emHpXLSRdY7H2CBrDYVM4BX
JyVviRWMXS0zVMjShWOqZVFyHpeVs3Mqt9V4DVtKc2vpBFEYRg48kmqWZ70ayCwKYayzI9ZKmh0C
3+jtNVs/JuwRxKWiG9lHmlICWExOA3fqlFVDqWfpSu2DS9zkx9EznNyTU3lV7T+FUOCekeDMGObv
MNRf4kp2JcgNS17mU3SYZrH4f7Ol/hAHhjfcZWiuwAsu/330YnYBuKnQaPcl2E7XMozacOTL48ze
WW0N22pPmmiheDoqfl8hJ2FI2PW84vNCJ4VSsbKvEF+Voqf9+IRcPBFiOprQBFV2m/Sqp3YV3841
v01LA2kc0PdrfE0rWMLJ/qDuGwOw1tafQ9Ku9lhOughHTJ7bg7cWXH4uJ2SxdvsW7UGqCuYdDIo2
RRauB3OOM+v0sumxuISxBQcTbam+qkupEX6mdqmn6G1iE0TmepPBdVp6cqMJzDI2+OXm7Q1l7E21
s48ARJRqxJnngSUOnEMZCJIngevGh0341Gpz18j3AL7behSUg4tjkvbNXRV62Td8p5ZQG7wEYsYe
hJhE7pwJbk1IR9evmMImZbHtoxGcn3mGFu5EfJZgOeTE6lJkRnjBKHF8glWt4c64uOtqen0SxeE5
OGOrcHiiTcwWJq6epOHDvaBOx2ZtR0/tZOuYDbUUsYqoy/R3TCzYbos44W99VECDhP33wT/Dgp0j
yiMgmET21/TqtIzO53BSm8ir1LDACedFu5WDuIkRWZf33BZSx/3v9oVilnFy7oVOPw3cAlZ+l0WH
avH0VeeOGUsjZkZYsakLWKUl+pbKCcmQMYRcN/K1QWnDH4KfzoPlgVza6WAhQNfN60s6Hlt7V+Yp
eSjnu5EsgrqvdQsGnJE0pmvMxy8uziSCFxp3JSlLtkauWjmHN0F+QwBwpVt3lQxIgnxV/TUiW6x8
N7KiRGuuhrLz3+BG47uY6Ffo6FaeWevMXC6whhTy2JXv4L6sUMIu/F8w38sPRn7IL8t9n+1guoVC
4Q7IWaJNTUeqnAaJx+p9IM/KzTG5qfmsNCUhuKalBpaqTOayB5OBQSw8etwSj7a04OG1drtAJ3eV
dbW6iygia0Cmnkvbmk/Gc2iTRmQgd37/zGV22F+Efz98oRlR7hhtDv1eVO9C77RzFVOZV5i8lFma
fppYOzchIqs8091n0UD+C8xznsnB6NMCYeAVq+NuBabod4+D1M6Z6VBopRmW5Zd9J+Pp0jCvZUZs
sjdaFK7vdE/8z2kJyfze1EaZoA6gsKjVI7WKqOICn4rrX6NrQrZ6gG4zG7+LkknQbFmJA7sQckhs
S8q0yWkvMlE6FJ9+DJXEyW4vcetHUp+s6vDEGtypYDe7Rp592Z1FLKB1xDB2km6nPDT7R6NZ5A/p
MEbX7xaYuqv7HQqJKM795KTJ4QgYAi75v0EZ0iJUTUjvhFd/LpKo5g7GT3HNkq2bWVT9OYuQq5tv
1WDItIc6Anorf7klox9quVNqN9rHzYXizA/q975KQYCc6WruKggK7eLu+utfzyFzujjHtgaUsMN5
HErl7b/ui7S045SGUWpnQ4FUiX7UGwxs1PZwGOLF17GI2NFDfQJ6JfISmUa2T6ESOagO5T6tCob0
vfYKr4D8gPSYop5elaQg1a4c2KwyxrQYU7muiNgauSZXPzDu7LlyR0TOS5FmIEU1kv/DV5adGMbV
Fu54MLQ0JCPxT0EPcBhE1JAOfPSwyQS9NL7Q5vFj92RdMMFuQe9yljqvcDtx4KZZiJ257lJJHA7N
a18JXxbw2NVwNVvMSHFau9fD48i8i86a/n0hIVlAyuCZaMToH6I9ynh0Nbhz0JUm6MMa1YYG1B+W
ApSeJkHaceMWbqJ0C1CTCgpcpJ3ICEMg7as63IUP21H4cxOmbuz1N9CtB4X99INE2rEEWUSsuFJQ
U8NGSQmCsroIt8K/enJt0/atgx6tnmGJkLMDIuRAleENga2rYcIFmhqzy/uDZ/YODn08q/opba+U
TBR1E75nN3zcI65kMsZ9enTnewFxQpdraDxp9Mw+cA3MhCaTkwJmES2URDpVUE48Sli2FZksSmhE
J9isgEK85gSRM/y9om0hAxgJhK0nstLB+mAgQ/0NysQjcRpiMgzLoYTHwUNzDbpZ0AGSXJoYfM3E
AIQdA9EmrDqjE2uv9n7T6O5EEKvR3rTKgdBxcCsjingsCBdqiHWrzmqZQfqqABUdnz+uHw6lOOWJ
8/iqwbgJOoat92nFBcA9tbC5jqLtkj7sgm+oG1LD0jeEl/9p41Ru9FafVmTz5VO35KeDF5yXzHkh
1qj7YbCg2hMKXNWsWPQpHYrdCiCz9r592mBdGEaYX6nzFXjpFUF+x4Ey4f5O0e1UibCcyYwfkUaT
Fgjrpv/HEhMKj2QVqWDvF649DK74s7nbyXST9xmFOGmd2ahtwHUwkLhJFFrXhZ0SRQRWCuErPVZ6
rv8+DzwX7ZYizS+/D746meKiCXJ8lYipuHQoEg54uO4Z13HybR2oYcCUs3pKOS9XXGyokVHj1jXV
ETnDX6sBzv/KmeNvfN5JgtI7EDKE0vYg3Ffv/FADnEYD+1xxy8anBXAKvYab49jtTuee806FWfNB
TqnIlX+HBEUFJygnKFRLfxCtVtewEobB+6lPpnDIBKQwbZzYWS5ve84752q8SUDO9h3QWdA8te/B
14pyYAKE+aWTscnzeyz1v32PhytmTTWbhh+SBqyXjxTCrj29Mmie0efHJ5k2ffuQVwawf+Ebah5K
kXydMEbNGZFUhNptCs2HApTugXsyrSSYqrvGt+gx4ggaqLPDeb+WadJ7BSGxgxF10nUtEYtSTXSI
k6NG60G8HHMPboElMKwS3AvVSExfsP7aFFlUM20wJLdy7dI5CW9c12pZ7O1ITYDG3r79USuis4te
47oeYzkeGuza7DL/LXehwhp0nveH815ng/v18+nqDjoh88uxkMFoJLeaTE2JF0qQtCRlDyBr8SAt
5dimQLklUUh4z3LeeUEqeQUUbTymvt7IDkznCmc1zX8qR0y6fXA6svMOFSppQdoc+7aGTSaiVOsQ
3XgIP9r67X8GjMe9mwdZTCEvmIFS+EFhBKYfg0OpbqmzPT2/+PU0LVG3JXDNRHNQz0SJNainDgo4
+NZqXwoFtxfXriwkmMZN5c/ZWvnGZ94mR/Z5SGcKaWGJCFJnBdsIXnZNk8SaSyT6MZr/koFAh9IP
vs79VBOlUHtAobGBr/5uEXVALPU7E0e4iWC9yLefq5GzRhjXEI21z1uUwIdw8b36roChYgG/pwmj
m9CxEw46MoDs4AZMyp4GvMf1NrE5e/uAeeUyiQT2RjWEX1bM6MWOeYUe9YFh4ql/j1bL8SWNVVla
lPK/vrNsS5Avw+AO8L9MV1gt0fwRO9hJAFaVc5yTsCil9yoHAxRzBPQ31DELkpmx+aSrpdkyuh6l
vlhTt4uS698uW0Kk3uTzE0PLaaOy86SGTm1F8BS8T4VSzHZCEdSWz900MT4NuJjo+UvQxbjaW8fF
3V/WxTuM3T2S6hrXxZlvRaNSwPYMFD4x+9zF+tQow1rAOXHftqWCteWyoK1+JVvm6uOpCoNxw2KO
mVruMMWLgMG0QAJ+u2bYSbNkcpOPLbBjtiZdlQkglT7k21/ORQeC9NtuW0uKPEuPbc48F8N5v6Cr
6xDEY3i4W2k+qtf38/P5XDx/iZxclML6cnqRnUXDYJhN7Ys0ZTIUuppsgTHyZqSZzBvYRchL8Wb9
r5PsNbr7Om10jo3VbEZ1iB47/tRroua04525ePKjHX9g9jO4MBCRoYhz0dzOZdiiHME3GCrNYU8Y
lKUiTpQ+387RM/BM/m3T29MM+Lu5xVZMNzTbqBwjWLVPYxvDm73OeyIG1d6RfbN0Qd31GR3f/avm
pbFgdXia5CFwfBoWFbzlwBIW+vBua8j1QWbfe1Z/iWuhLRrW2moAxE4HN8Jyd7FNxn+hQWsHIEdt
xWKcfPR16s1aPRCCfCKcRRILDij1pGgUBqB9jLNkEL/q8+zZttXgpBBncZZMiYJ+siGbF+XmS2h8
X2GVix3TLmCZ17rY2cZav6ODqSkgtZE1RozwZearuRiHDRjxeOuLvMuEPLaRyC3OenGHKaSl2w1i
opB6dGeNjpULXBfwF/fNCEvCvlaKaoOsR+mh6NvhXhggyvszh4Y4KUgSHgoNNb+/6azNnUWQSiCi
6da13sYJQsoFnNue6Kakfb6o9snj4zXRsmY6HRJcqwK5Qobhgp7o4MMUXNnSFTIaKb2s9ZdoCekq
vrmzus2Iv97uR+ugjqVXMfw15ap1/shI2zkrOAHDfF4bKxCfjAynbWvzHBq2fZyYyElMfsUs/Fbx
fX0EmSpVJkK3W7sn50CSu5r0gXAkMsQ0Sz6qAxsX3K+edDn+7XZUsihyxpdRWfkjUR5z/nb2QIq4
uZfh2Lh2iltX2l0E+Iija1nA6OL0TDjU1CkS942GA+z6+Q0L9dpmt9nVKUrEYOBJ7SyCDu1qbeHO
PQDiXRvH4t6Wc7awLnuFoO3J8dQgbum70HCubNbmyXS8EbR5iHwpNQbsaFD1k5WUuwICFJnPzxj+
spy2ZSmbA6e6/b1o04qG+DYcIje/k0V52WKzhNxmmWa75Wkk6B1qhbIbqOFD8IIOI7+NJjLc5nSq
+RCqijG8VFfpTIfBnguPP9nQxyobZm+CJZNzqGJ6pHw9e5fD+K0coN1UK+Heg4F3NKxGG0QcesaQ
EJTg5tjXVf8bGTnUbrxDNFKLB1jzeJed3TjUWLC7oDuuFlLAoItGThjAd6Wy10gf/b8moU5uoaXq
VPbq4PCqtp2zdMpcNZijrQ2/LbKKi4Gg4wdLDoo89rizJOZWUbv+hMzbDfXMoMFRuhzojJeynHl1
KQ4P/lsvS1ksXKBzEmIX2ilWhm+oBTp9ac223d8wok1QTm/8z3o7bBpl4KT7DN59Fa2b2efco79n
IHHW7GEohQst+7TYoWnOpdnBqkgTGy8y9ZrahEt8k9YYqEV8vDmNn29lSCgpabEU1xgoAeJRZGnA
PtgLK81i7+mJcN25PeEU3wDmAmOeGcWJx+TG5FxwI/xaR3BBFoaTna69ctC19YdSQVepH3z+37ox
tVd2IwqzwQEssjb585ho9nbsI5s3gjbJ4/uOk7Q6rtTaJ2q1piaQ1IN49FYxoM2Mua43FO9pTqxi
I1n3f4MOk0xS8XrKKzxs616oHFhiJsCMwi52koLUoWhsb2AOJ2dDFt5/APytytCefVN/AjehrGR4
QAWS9+P0srS7RT2g4EEh5z0SJVkMxbJekEXkS0Rix3xTxwMh9R5USwuwGBCmqmv4pNTu8KaiJpdb
dm8x8C0YLpEn3JhMftfSON8c5w/Q/h91G+KhEfbIP9UjGZ3fuH02fKhZdosy2vmt+7dCPAVBlApN
I1TZwREkrEtFuaGAthlkghrmoajOnS2TTqxZ0CGWrfcpNXfW6k2fY7D7ngwrGmI3582jyncbWXZJ
NlqDa3D896TOsO5qYFXUlhchJ4fImvSgIDhUkftTeW7O7GowjsDpy+s4MpwX5aMOD0pOrtu+gl89
lVE066sig1LFoIB/q2sUDi4oQSAtGh7Ny63AsVP8fwnJOmmUT74/7bmf5cGIdC7RbbYKjA+QcLpX
/hwGbICxlQqGE/erjYdmRQO6l60f2VVcDFxu1HD7ADla0qVyTpIwkBSOgEG25bVUA+UGg7zcmgVv
aO98tvH4xRM3RuhomH/GMSEtvQAAT3Lk0i28U2YlSj1fR9s4Vsy/bQPIE7QqZWYWNht0anuyjSQI
OTQp20g7JspuhyTkQMrHStCtk+jmNbP27jjEVrYrEy9YZfxGYPJx7/Juld6CiRFTPNjTfbt+eSYl
rMzM5HUh/NXBCSQNXow37WrorGce1x7yNX3b3Qvf1zPWNA1vXGt6/FwIsn+t/mEAWztjiUd6AR3T
EU22Nr5tUp8/sVQ/BkxhwDiQHoIyCFkT6UHLxGy+dW0vcw2OXQPBL+xWqrzIvNNuf5VzYK5YVsmH
cguf3e40AlWkblIzapcKVMYQkrM6KrHSMxR+VWRz9ZRYolcoQBk0SgvaXkByuUNOnA4iuVzkU/RF
FUZs8XX+wdd7EDCBnlq5JJhqWzNRJXVe1cc9WCZMSIHgTMs4Z4WJpbWxpIFediK1oAR7ohD129RX
JsFxkwgu/HltMH8DtlDAqY25jUzMPrHw7JAzKVwn9qGPo25B7Rbg9klfc5VMiPWgp/VcLeCm1CMS
ocVIwB1nOtFEHaXgfybEn1luQeyZ+2IdE1n7SiIIs9c3tvaiZRwXceMCpg5yiDUSdkLoXMH5+b+R
0Ul7lTyVm+o0Vj27sg7IAIVMeKwNTfvj2czzyim9tDa0VbkvzueO04LcvqwOxnXhznkLKRjTKmUi
x006LBj4NeKt9Iy3bjbKgtiyOTisACUnOwV4XjNXlqDz+tY6RZ0zka8FfvDe/P3/c9qGDX4brNn1
vtUIBVrHrNzokmWwEmzKDLeCTr5EnHqrMRL+iQegty/OI41cJvV0+9TKXZZDh2fMpC1nS0hYJqY+
XGGXJi/XA4NuTxAj5D3hh4nbdJ3xzRiGGxiN22e0bWOEXTq8NVVnU/x0/V17prIljLCRgjHsL0EG
JDM9TtaBDUuikwEscwYZryuvdJWOecpkIy6I5HAxPpW0LMfxuST8+01Uv0N/gxp8GKmSAkz/RR3J
akXpjAq38AQYwgYj7DmdpR4+jjHe9XYFUda8QG9T/8MIyC3oFZJziqr+1C+UbShi3I7iFdi9e3sy
MOugd1MmYH6hHHrVUi5Q9q774GhbJMzwBTA17SVUymgTH+FU48MI0e6KegtWBlNAdai7ysn9wQa/
tdnJ1RKNcQmPMYdSvQJfQdUco0ovkGDkFxCxocQW6qhERO4Rg8RoeOFkoL1/K8LsecON3J9mp3Cg
KQimaPehHr5iibGlQzC4sz1lO1M8XUZrQaIiEaNOcU+WvAL2Hw1Yl14Z/KNunK0ZBxadg+ixa3ZU
tc7mq2a6aP7gGGRrXBbsiZj4aQUJceARdPTbHIQqbAOUpJVb/JnPbUZ+xALtR2bmpDxq5MkGo62i
u6yTyokFs+4G4FQ34N800k64tJnb2EeCMNhd5MZU14z48meEQW3tBYYFj8IG/RuFZmI22fxY7lon
teaPd8yrvl59Ldx5LkG3XYwBqvBSb71MkF584xRNp+U1dAljL309tGUR4IKJtmYKNBLy3aLuWZ3g
T4uO3tQzyz2yr7dTdRTLHRcd+HVh98Mgjl0Fm6q+Fh2nlqHlibf/CEcaI71PaiRjZMWsaJlGWlVH
VocABLbANnNp2sevUKMpZdP/91NozQ6DjexX91MKjcE9iyDtvKXVGTfO/6/YGZYkp5114KaQ7J1L
XVoJA0qAeLRRz0rXvShPtMtLiqMF3LCu2oKvNWFiDfu5jtcHKORzSwGYxGZXZIXevBUQ8p6wBtn6
XJVNNhWUHQOWi/weHwm2ye4eCN1SeIP7byJkoZ3eViQA5O3Q00ZL+EkPoFaEEwtUOihYirAWwh2r
NlIs2YZmxDol7lNx7hQAjUJzmT53CreA2ax5cMfUiSrC8xf69ZpK4gaKD8e/RHxt0mQHZcHUAwGg
37uvFkqlZtqy5KfBdkekcbQcwV8QsEY4BF5J+EgT6a6gx42wedhj5IgE8ullUzbybC+vgECjbwe7
ttKFEHZ7f7VfP3Ps5hEFWQ5Z6THtZ1vAUW32dytEb31BZOisDLhmJ12Wk+4Nai0cZ6ScmPEfFddF
jSAw+aCoU6sT9z0Zz9toqrsIvI86g8e/ZockGIU6vhbO9O/MKERfs99znx8xRUZbuCGqkS+ZuioC
3gs2cUG7iS3KDswahnPyRd48F/6/XQ+RfcHL7VZ/nIVM310QpjKsA5FY9AMu7XeOHOHgdLMZb5Y7
BCVDIiDc/cSD8z+tem3jF/Sk3thz2Y7MV5HbKVIxB6TEIaPvpREoZIj30aa5MuadVMeC7XgvHkEM
SOI0BM2Ud1ZyqCpS/0O29rbEb/m3mB1HB5ovew8CKe8IXFmdzEtxE7j3D+F2sRf7/FPlJy/XNEkv
JQpNIDC9QiGsm+LyPLQoP817WYUw6rrhXfxhATb+3FEj+n3xtuLtB93oa0mTm2cnts/mlf9Y20Ou
3RKL1KAVSS2e6EL1JuHh+LwuVfDZGPN6h4NolDxYYTuyDr0Va1BrZ5oATbDOXDw1vdWkDcQaRQwl
V6yQiBwgLUVwbk2CkIsWovx1fQz+SKNC6xWWCthl6FWFouD7NTAmCMMkGmoAFeeFrbKvRBuTB1/U
QCQqDMtB/9fT1+PTxZu/v7jxc/5yr2a09m+Spmz7J2idY2Ty3upGrCtCwwQK0kOiYHhGzEcLX62B
U3JlUygqA8Uoi024EWxf2HPow/L5FF3yRP0V4WU1EhWBfyvcti3Kae/uWfhTPVYMfezASC82x5lh
TfQXO9pqaKdJ9rAGFO0XzjqsWjal4lyguiZiaRwB8IaKhWgKPsO+UFvEnVvpAkQWu9XatsTvzWmY
sGzGwrmu96zn+8N5x/xl3AbnIp8rH+78CY9RqxcKDecS3iSDHslX19VIfI3xf9+dBqraoe2aC/f4
+xNQmYdlx1XNLGdBgBr9/UOMs77iVaKcutu6HDqq/yYExkIAK7vuZ2F5Xez8hMEda8eBX2XR/g69
0CzNKIUktMi5Nm/IpD75VIQ+CUL9iFddA9YCUkdWrXvj1R9o9L0DvdYHRriCCBQOwJCa647GCCWu
0GVFM+nzV5eHnVQoofkLcqR3hpByKh1xS+45nHxfmf5QIE/yCB9oMjP0TvoxZJPXemuSaOU344QJ
RWQdpUHBjR2gpy/1WMYN+jAbwWgmZjCWzu8MpX2aJfkQilVSs/ki1nqXLVVtdHwSa/XJkfE/1++m
PUgfAX/UyqZ7O+gRgVTRq8ItSGemWi5PcmBi21uhgxxDMGEz+h1qP3z/shjU4GVQV/+M1RsBLCXU
s9x29b+uHszR7uvQBDl3HCkeAQUo2YzjiTOv+EyiWhsqBVDAbJzQjBYMho0QUvG2ORqP0PReCO0q
Wt1+GILGFIn4o3P4JHxueBfPrAXPafpY25zwGts2CFw6BYemBHvN/gI+Ezh0TNblTwgRU7hPpyI4
8Xuq/f2+33m7gKGH2MX1tSZ5s3OXfwT3I8yITaV6cKLTkuSsLL0leUUEclw8TrEXgbCU2gYm4Zr6
dlVbrTJUpmIihuVgpuWxD3VNSdYT1nkukKEhuWDznh/bFe/yee4/D6Gz1+rbDp1Xg+/ZwiH37tXn
Wu1OIqWqYZlFS5m+GQh77faHQxVt4M7EziGurnOZrcGUqf5NuE5fHr1/hEXMkUs89n2WuKuSGZwv
fF/9kTr5X9KtM/iAGf7/xxjNvdtnpDcY9aAm45to6psZdSOuJ6TcAbWO2IsqA5D1FBqMeFivIPrt
vXlVz9dJb5F6+BWncbEf9LqycxEJNBWzQ0mwH15LaGYCs8GIhGTOi3tJ0QBr14CGsq/c3IgHjzpn
hOx7aVquWoYyIGoLfwulYjRn0czFJMli5/WChMZek0E9ma6gajpwkI80XDpVAUo4mBKDzbh/wg0p
SrjiOVrT4lA+2g+sY9LU7SNnFqSEa0an+YAwPk7UEe3LnI2xRpUoIyAxVMZQVUwmdqkUpxQO55VT
XbfwHsH35mR7pYc+10QNpriVmGU4JUcI+rEifzdL/hQFNBumMG+zkc9e7UAPVcOJ1n7nN3hSsk6X
vdeq/g55t3dCV0CmoURcSctuKqhhArDibiQ2TuRidzQHGrbLIst/Kv2FDGtsSxxgmc6VIrUf7vBL
kdq2vwWXduwsSZW6npsaMv8rhbtAcPVhyxwv3VdpVJBdivJq19hlvwNEMEVf5qn8kxJpLBc97mm/
A8E5g3pwErcLRz1pqEyiGQn+B2oKP7zpALWO1/hF6Roije+8pkurXZ4xnnODMYR2xRUQtQLI3zy/
CbfyMHR/Lc4KgGerwqQvS9VYwiPz+4nyeqHFNCvIwrFPjmT3cGqtiacm039qzmhrzrMEjHwEj9/T
SfuhQtuucQcTtuGdM7hsrlo9N/L9AZt+lX6QOjPyb2AFHiQMV8q8qgYRKIpvtpSbTNYG6KnoVUOq
n4lnMsnXelOfYcOoQ86LXWWYCMADw0xx45xfc6L9+ntGMflbIA1yLsw6m5FYYtA8DFVDAJxrvM/P
FaAnCWnjBi3tQuk9D9kudouOPPGyZMmkRjQSVjBApqEwHLYBCSnx/j/W90lbNzK+SGnLx8Z8NWUD
2HXwL4eAB7R2wXZHuiAiZFZAbDnsGfT2Z6xcgNzT7nr/x88Bp63ISedGhRchtRxycHDAyhNRjGJ0
oTGKgk9DtrThqDGyDM8ThxwCAcjhGP5tyV/QDxgTJpW86eniMICGJYrJrtY4pZihEoFYHEOb/0Dr
gSyadvaGxIQIArat1udWxIs/uC6hk+oWVfaNI+NypzFePM2fBo05GcLfDma1FQnVwtUsJXHEIADh
jviQTnCAs+V1bvEUqnVE17kQcmCW4014kK43oTXVCckojh1DV/YanfALAr4L03lUOY21shhdq4Md
Yo7ixYbQ5ET+osHX8WXSDT3BC+Ow67H+OsYl8Rl9Ur5XyFxNZde2SyfXYY1Im+dcl4nSdZSg1T9z
LaOdl3jNHez29KDfocchXe+LlZCAqneeQkG3ZX6nelH3Y4rYRCW/QP5cNocFkERKcgkE6bnY1FQc
W2SukeMUXmvu3CRkOc26mvj/5FjAuzJnpI6Fh8HjP02r94ZIwf/mIrMHEZ/Oz62zJs/6kpvASpYO
CSd+TAgGrQ5shVvQgZ+5A1LTx3UvfZtJ4PO4cUetHM1r1HCgBwTTBe65mA+tRb4mB7zHjsN2RTNo
W5WBOdqSrmZsWBs4x8wEoYIasDnY7R+16Yonvn+fi9pDmD0dtEmS4l9Tj8iPhRhBZSh3Ic60ADIE
hA6pvYffDyTg1369JztPuQA4NavciZ8r9lt2/V2VKV2TL0tbKaT7EPP8dyRKg1N+hSdPp9uBCisa
KwEXxujbxAX4G8uYNxQYIzDtY7x6kpFPM6CKUV4qWTIvg+Qe17aPYUjBEFAu9lT6IkHdDY48XU+/
Ylexwjk8tPM8z1I45LQQzrjnzy9SXsdSBVdfzXVORGt2WThDarkOoa5Ru4Y9ZrVLDQZDoFLe1LWK
BZHqqMoeV9icPHOktIDKuVvtT+kRXk+rR8AGURo9PV3WgoYudZXKLLS1yQ+PEhCmR+TIDuSdwgel
aN0ECzmPtJLBr1PirAsUnQEwNJGoTwXOsbdObmRXijR5/Jh6B2rvIHuw07DhNatjK/4=
`protect end_protected

