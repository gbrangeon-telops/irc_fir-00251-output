

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
To/0Y2C4coh8VFh6WzI2wbA/wXer17nunFaUIFXEvO3kBprRAlXyefibFdeqGdMCN/jPnm1lnQge
X/HG5CdHuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nnkNk6e3rHUR8DaNj0C7aWkCs5LBgvWhHhtsF0DtIcgM1egO9JMHLS9VXFoTsIgw40ekMylMZAif
7Mz04TLeS83J8LIkLQIVFCxUoXkTdVbP2vwAOIuzbV0fNimpIIdRDB4Qyrb5oJF0cClV9EVhM+PP
xrslkcRoMPftZWbNXzc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fa9acIf/jWyoTf/ZQQ2RdBUZgeC1x0Ej+f6KiTiJLxfGAO1lB8jxkDwdqife8FqrZb9GuA0CC+35
3eXgFQAQNKjhv24q1nYDvGkg1xQe+JaS1IiyitufBE9Oqujx03ehRV4B4wJ5uK9qxFjJm3WBZQeA
cWZiPDwrU8E27DqZYUHGXiufRSfFhYToep6g7NhnZGCmAfAD7Cg9pLa/AvxaXAS9nnGeBo/RPlyk
G/XXEB6YF86+MUOkeRMAxi86Vcag14njI42hNh7J8Lfa4beMq2Avi5tz5eGJq8y6uRjal6wz33O+
m0Nk9SOLFKAmJ/ib8Fpq77uCjrQp1T7Cl70Ebg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h4sQ6/cKFAjr6toNt8WCtcnxvbT2RbQqvunqru/ZMP069wFljAWXbbabme1u0tsoVT7hQ/OZYU4t
+qXe0sbPKDx8M0x1MxaKDasoQ543qKQAHxR7Bn28bTi4sQCu/+YxH72mTMVFjRAGH6M6e+MhTnGO
FYX19oeiewDQZSakDrY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
C8DUdaX7Hd0diH5RVXOZCPD1GItaWr9F/mVcGAwJsPm7j/BsnnF1JwcYxytFDkPy0E+fcaWYKz9u
7/hZwJ449yH3vkp0VWbVjDe3BqRjhnTwAc32kEGR+a+f8HB/6hGM+mJkcuw5DhoveoZqvYIICYqz
iQAjheEs1g2k4DBWxSdaCPNW8fXVd3J/pZQSuvaNRnCtPGOVMt3rO5k/WAzjiaWwDL0KdanM3fU6
uD93ZtkLZCLilGdf0EAax4p+pGVd1C8GYV4+XW66vJmZoT9LNfQ7rG/mL7dKp2aZ5DJPqw3W/O9c
HVwQSloSjbmiN1Fhr9Mdj7iCZycwuy9BYtMK3g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24720)
`protect data_block
krn+ELRivkcesI62cmRBj6XrcTJRWhXtxot7hGlZVI+rf4QHfprG23cNnFxEeEfbp7Q504uByxDb
qOLLsTg/mL9GICLCjtcDNPw6E1RVRvPV2u9/mEpXjuoOn8/UL/E52y2Tw7UhGkDNF9JM+uT+kAl0
3nzbPct9jAWMdkC8k0uzWQzV17q4Tw3/u7mD7LtBcKQH7a9y5PBZnwnmvtOqaTwcaPeiO42UsrkH
wQ85z9CU3evsVgIwh0EC2evaSq6EX/QcetgYP5j5DHESH9FTzt1dvdZNjHcTo9zSc0KqOy1xwgZq
Y+8wUlmDeY0hlKHM2Eaqxh8WsNRQ6MuUgjkQLRyeXwS9MheXMzwBpeYYhGXNSw1yC+boZ5nmvOWc
/zEkefV+L2uVKqD9em3BRzI1uTHwyXtSbCSViISp/zyfmBJOiTMUWpOmS9DezDTAs0+fdjbswZXx
6iHoAO4Q5Oz97yYPJlBzh5IrQP4tTyZPNvIcPPOPO3Ym866CIhHcbcOEv5p8y7gbvpL5ahItdEWW
PThaIsTbYe1M7B95qF3dxi8ezOLsCTjiUu+jrLrfGXJcxgBDecRBw41pcNtqBlipAYNZNbgtNg8y
j4gCduaJvfudd/L4xMBVXhw/8RIRXhfyMIvJVx/J0/6oX9Rr0XnRgbnLZSHL3zp8ODtY4Hlw/qr5
quezZu1ZGcVB+r8J+kMcATr8emurtbEBDf73r7FM6BhbPTuS24v7s4Efb/ddAq6ho0EimOkACvTa
YYaDiGcHRWVwOCGhQuDww5tGLax+FxRvVEtIq6NbIjfa6OLVeuA+OcZFpn2nRpfPHRw7omrn+78B
ssSn+9fkDuLxoNuf826l+H8L5dIg+gay5LsWvwTlJhQaOtXEi6ywVDPOk4BAT4y1EukJxDORTk5C
smYH+XZ+ncV3BBPwRyiaY7oEAW8zlW1GqLzqt+Oovn3lLxRNTdGyBsXKg1BhetOZEjy00cIwCMWz
M9H/BP+mw8fOdZ88+Uqd/myOezDIg0L6IedlgxL2k3R5HGprYrCSO26g61ZAV3vxIidP+dG31JVl
LmGFpKSmP3AyaEghbWGBKE1MOxfntiiEhcgY3k/LS6xBDbz0gWeJpvbwar3M6eiFaP6/cIqKioPM
rnDYtdAvXb0Rf7pSnt8Yo9OqcLTwJS69ct6NN3dK63EOAN3IZ8w7INsRmnoCPiIBjMWd1omnEKDl
cyDwi2TLBiehGlOBd2rFlk20MMERIRfdtM8X2iaXdDut3eh02vDY5zjms/AeZiuKij0kZy4Ed+eO
P1mSlWO9dO6PJyWsNVmdRq5J5txg10/qSNI7QkSnyJWdMqYV0ppB6n1XdBAMOK/33qnxlaIqls3k
lXhmpn7GLuuCw+5u5391V8QA2vOUxVcOEcJGIZ/7btyvRlfbe+HgSmYZgK+EAZaX5Am/Zd5LoP9/
TtSnZMNScih38LFh3XTS3xhWz6dGrZcyDdhnsjJT1tpnhOZaovgshH+2qEjz/H0RwSWHWZxPignr
Kr6Sg+/rwkMfS89c4tMtOFgzUvLodWi67FHTlJ+mC0gu0VgACdMiuo2L+3qXkteUKBICVnE97w/7
gQKk+JJOi0c7DV6zc1vp7bz6ysW41eGk4uRPJEAahz3eQRls+ppuvEAnQcWunZceCtGocNps4wsF
yQCz82i4p/w6Zk+2GuwKKAJeT9p3ezXX1thn3e6JrlZszsbqgirzmhheCJGZcAUiFZUxCSY0hQX+
iFAwBfaWvo02s1SbjwKSHtJgb/pissZB555FemYrDPqlolOvmeRWdqhQinClRnxjRmh3HYjEBjj7
EWmJZGgFRI8fDbzuioJDG5hr/+fL7QUDmmens4a5G/gy+GlkNDTAgxRpLUrfHHBthSh0VCBUKAHF
x2neT2we3fFvc0ZKMb3uo7gY07hRgffuLiP0VyJFFlcMlTMbJQE2pkt4wjXjtUVjo+iJE8zC2RlY
JRbyYWX04qjLgXcT/r0c8Lx2RxrTpf2WjTnNm6sPMi2WM3ZuJNj8j3O0HrupZsjhsy/mDT5RQu4y
j9tFtHmNSwkDC2fIJdjBE2c+Qey1HYEvOK+xUZSnCsakgNPKRI5w0ZCi0Rsw+2KKpP++lXEFL1QD
VygzRqgXEQ/TAZW4cBu9VdhLy5QPu5QdRPs+E9ALNMCR0p9sy63JCLRiCfL3AxS2oNbIFUAYOuOQ
sgYUcbFs5FfG8ITKW5zN2eKmk7xoYO27wI8zwqF0V3yTPysrec3FEFRvdnAVVB/GQgyXvrqQL4yY
yXyyMJYALVK8iFLSsBEw9hkOzm1OQ2O2i5h2pyWVxfqY6uAzZF379mmhzk2fMHYFE+DW/W5uXAvM
gGc+np9wswCGrge8wlqOr1XDCI0MeJGDG8kKLXtxHh8wnzWOljPJVZGsdD8ZU2dJq9tGLpdl5qGk
HiIzpuEKiWs1AKtfa/M10ucr5ed1k5ik6BTFAf4DgOQf78v7B61kW+ZXjpHt6MMmSm6L0Qdtwmyu
R3XDApMJUPkKRm+2YUdsq3CzURh080eUR3pfRdY9M+uYRCGccCP3Bk/8s6hzihMtrlJ19mkc4soq
DNkGLz3jnkpYEdXjLRDwNhOGOyBHhfhj3elkWa9EUTCQFSO9oj7ii5spsj1mu25JHo54ympm0+eG
du1krobCkA28jfm0eEZK+BVldVrLLN65C4IkOrMjGeIjCS+i8nt84bvDFKYEomupHYDMP9GPf6Fc
nLPA10r3J1nhm0Ir9G4gFmBdCI5HTOkysOxm71svEBxNG1h8bHU9AuN6LjCOCfEXhz/8LPWpHOLN
eKua1sVyhl+MGdw6DSua3ug76xRFFf5Ofja/lQEihESJmPvWvzgm2qtUN94YvVZSI59yl9E3Pp0h
IgLySj0ZbiChsrDhsA3o5BBWqQr4dLdxG8PV5MNUS/EF6bw7R1Pr6TXs3P5l019KKq1artHio7Su
x4+4FArUFR/zmITGLHQ7fPLTgkIeegeakbHhPUSRdS0Lu5w4oaB1jufdh5dXxuILgOCNW6h+gNZk
rzZaEdmo1nEMZGw7Jw9pX2hE/Ff/9Nzzjzlf3sMSldQBGnd8D72Ole2toFbAu40MwaZzko2oHpIq
MXcBs7CiAz3cEslXMMjbnOzNBTxBanyPIL6J2+AOL+f5aYF/MIwLtV1wRjtKdTPYN7I/gjZ/vIB2
Lq2UacKs+Z2/kVnna9NhU9g79QKbROYRkxmoGZKeIB4034usPsDpx3+Vp6sj565GzJaOtzKk7Dok
A0Krq7+f7CdRWAKlT83LUDu/GYQyNzC0CImTHYq0bWFwZRmXLg6upDWJEZz8G6Ry5Amszqv/Nc9e
itbhNctkLzFNN7hkrMD+53c1Dkv1nxKJeNgCzx9739RNQ1Btok/DToF1G1k1hyMPsWgcNIG4s/v2
NilppikqyQBw/5Du/YgW5mZrMt0sdRotkKbY1kboyvlCz2OKR0J4GDoBrgo6QJPXs2oYsafnpanw
EeJc963WB9+ggTqYbIEXnIw0ApuCoCKy/Z6u2boBgVvt093uvgHNs4P8eGkIL282so6Lv1olH9uZ
P8eI6qhK+voYxeF3Zyk6ItSOXlQCzzJqGTRmPW3O8S/Uu+rLL1cZ/CztF04Yc9loY9SeRqySwP9t
9r/xb92EWlFhbIEGJ8yQCdzMKSOB57EMptum3/Cpe9Qp9eHlI0TUdxuMr/pALeeH+aCh1zVqe0aR
TRt9JP1BIqCig7Iv4TTovsuAGhkOy4SUq2B2SwwhrYktwUT1a4cYxqdnoGcQnkmlb9G/shT9+Qgr
/im/K2CIZlN0qTFrMZbbneWLEnmz1Tq7i1ktWSVTdHDUqDX++9canRc8F9pbGa7uIoIAnUwHw4N0
BU17X6mw2m6CRaGREhkI6H2Qbi8G4mZDoeSH6jwG5CW0kaIN2525tgPTTJct96qdr1oY1M+gLClG
ptSX8GCL1BNDlTsMCYn38qM655t33cd3UV0I3Z97IT5cewoqXRORcMM1AKW++Kku1jSXnCv/Yrxt
uCqD+CNAw+OuWLz8d8IYykNK5Ijjnz1jxIu39zxoOqT8FrDYVWxkZdnIHklVGrFF7b/CoXXcmA7N
WJo92kdye+peah55nQ+LHXaodHSaKauTmOGZPTY1PqA5aE403uYMU39U9qVQWjChnPW+YJAAfbEY
xnG81iNLFW/IdrgmOgnbZjlQ5/w8g1emUqORNm7lu36Iqqdarv4zwCTXdEKO/QPh5amr6MjaQ8Ur
7k1mCJ5hDplif6wRMqnTUHCe0XquSz6SEyEHxiz5OlCkDCCfqxWn6xqRTbUM8dWHByLLsXfUh7LI
/rdlHdXCbwhPSGKdsg//RMcPUXb821wXq44gIm/10KD0IVqumaCstP9XEXnC+Z27SDjGkSpBjTGr
l/KIfV7KG7bWVP8SA/A1iGK+cxcQ9pEvwhdSYDQat3emNoijC64r+uXb7+GGMJJys6m/da4NaFI1
z/apG0rkye6eZFBd8Q646daDrZSYdQERpdzQKHStkDOns7pnXwXZdZNFEk7oM6q0Hv2r9QPHafc+
nCFR77OAvAq63uDK+/7I/v4w3wTUfrgg+25pRQPlzQCeNEkHJyVhGCwM+/5KOAe+C9VDTvdsICJX
yeuH13ehUAZNd3cimKN6ItjSGygyOw6/aYf8EHzHtwtmehrFokaB4amm2GjZe/zkxLm4jNPM1OFm
wael+XRmM863IwWSEeP/hxqMOmdT3W6Vsw6Jf/BfWq1I3Jvw7+W6P8C83N6+52lhmSX97/K67Ipm
3KqXndb37tEn1Tp6oYNHmCf/T/3M7qPQQxk63ke3UDQYAm/adVVDwoJaAIfE83FU4mI+UHAdnGdM
Y/ziEplrSd7VlsQ+TT9A0doP8SMBdC5m/97413sWZWMNDSfq/oq+S9AlR7mOvwjR+NZBE1l7EOAi
nMiOPyElUVEdZo63D4SdF4eCV/bsl6vIwzqJ6UN8WpyMLGmZEm5JfRG5+lJCsRAmwNkNPE+IKD5A
in5YNvPz1aZ4q+AgGzuvpxUoFfo960RyosyytBYKxaAwOgGMx7SbghuyfOrjX9VcSIvSe5a+kpb5
p1KWU2ctvC1GDJNgsXcw3yxhOAFhXv7hqJ03wJrp0hjdbYUtHsPiIkiIxtvx8t4cof9pvrbY12xF
nm7PSKPgFnpmOPodfnJb7ePI+aQraQllUrfPxWRtCypDcc9X4cfV1UYrwPvKJJzu/GWhTxKjTGn0
9NQqFowQFF+q+xcuugprv20Qu8iFR+z3lC0z/wMjxTDh4Va2pNjub9TrXTtuEqh03fAAQXn8VscZ
pdaUCm9jSmZ2cGHbYm2inVkW2NCOoXu+iatgUxBvMRMuoH1M0i95SD9hQOwk2goC22uVUdXPBhYk
36obfNJuhxbn5ss9B3cfOzssgKUSMyBZPSDrPwqzyq09rJOC2GA2pKP6BKyDtHeM1CwqdT/FGgOB
ngpL7n2c7s1rOHq5tDw0Hct3h41K8N0hsqo+s3yfvh5GBNJmNQq19G74L1soS7gQNr55OYxTTE2a
JSiPUYk2D+joQ5aog/Dh9ZsJoN3+pnpKZNNLa6sQuVsh0ZcQ9tpMD95yTWdKruw4NowFZ3gIRQpm
u7rVdrxxFbM5z3bXy8oK4bqtdOmLRq4xrXkvZcBTdOrcz4R0JagX9y7gu4KMPUNWC8NKliGzO61b
URdCpPMSvIED+i75+MnHM06Z/PH0lUTkkG9hfQSfFJuJw8c0xlaPc035jOyENHPXOOo6swx8quej
P5vAmWN9Ygp7nxWDmmyYBuR/pTMnxCuahRABseafw5fsfRZBiNqlLE5ulObqHMpwR4TpEAUB+Nka
huLdfTBxIe2Ds3FNRy3VGZteJspjcJHT9bzrlsvE5xZ1xpZgPWivdCNxAQwxvcbtb22wV+cjybg+
FI53jo8fpmtI1BXLI+8TOohmoQQKUh98G0InzDRbY3V6ONTdJzQiTlQrJzLGm5c0FT6U6z8D7+mC
WqJ6ofzLUAC5VFplM4AtlRYGzAVYRp848JU41T9EXbhjAuQGHTOcF/fYNPM3xyARTKz6rrdONHrX
5tiHtaNVS23wsKxDJwUMo+rU9rP8//quHFvUVCr3VuMGDjPKsVWoVnecBfBRJKZexuFtcp6dCGzU
kV20S0ADDVKYK71b7Qfn0+y/bJQVtqjIYL1+1xuoV4CwH0TE35GaJE+lfR0n1O1JcnTmNPx2SjjC
Lccn3rZZTalRYmtBfrTPExVIvxw8F9kmQfkHMGBswfg/XgBn/smdRd3nSptkhHYNELdbEl2kg4JO
yNkCnKSQOImeMpvoBeh8MAAc/I5fgI3bieCTbtVvtlP6CR3WCSlz40uLtRLQu7LhckXp9tBRxjjL
tVuEMRRr9iBcq6ZI0jmWIa/XqusQ5TrQ0v7AVev3hrN7ORSjrPV+MapIuB2ul1Rt3XJA8vrNEjD9
9A3RyQALGBLyUp0cJoWCgBFuS4RYjBsgXqkFWvvhvfPnP3lJ3jCA6ilNTdqvDqW4K7qLtUJ0tKK9
rfT3Ri2DQzUSEwQTCQR0TWRIN+Qx6248XC9P9ock1mBY3k1hjwx7YxsI4gkkpsghGFvHa7HJibfp
FQ/dVwSnrPlTqzQb1y+hT/UQgdmyrjTTHj/s3wlthwhiznVd/WSj35zE/1JuJ7VgG8sen3iGki6u
eIH+7U6fEOtpuMD5fEAizqsgkrYiYbF6Hv2gQ9wUWIdx8jEnQ5NBisUNrI4bMranxZIbTvoAlFN2
OUzn4lEI2PxjVPpKX9Tep+YLuAX1A7RmKNtY5VwGOoAFbS8DQIwSRfEWtapLtq3GnOW6i7NXTr0D
f8HDxEXsi7ZokJnA2lJ0Wg7/n4e9pImELHSYq0wscJhStydgKnIAxO5DAjmu7nHlenZ9CK/mjuFE
fxuu5pXiTdQ2t/CjA5naW1/9cEdcVArgDW/fXmRzxJlXoLtMPYcDxePhNWuyA1cKGcBP6jjQawAJ
NAk+FVAcBR6fDqAS1mgyABrzV1hiiDXv+PLouNV6F8e41BRW3nPIl1lxloSPv4wokxLSFpsPlXTx
WG6k7eTMm8LThCBVea14tAWM2AhgWXZXiohO22jxcJy6TCXEiY5AS0s/bvrUkEdOpVCTcbqlykwS
rwrw0C9Y4fru6dC6ZuxCNWqk02dI98e/RdoHS4O3tCnb9zqPYjO9bTeP9UMbl1v/aDHwgB5c44Qz
HwMWNovqfPRwEpRoBn45Usx5ipW9zl+C7nv6pw6amaG04tz6tcmnwfV7IDa/09NMnzXfX098jsLA
NCiMPDNk/wi0UL6E0rmEvZM9+qH0PTNNVQmkLWC3oggJ6QotKUc+QZLS4gdWvd4wtm5PMD7jB4JI
ap193yxoaFI+OABacAbfQfWCijKkKoRiY3Xrn924hDcVR5QAl7a8uaWVYhPe6QnL9d91dnruIxa5
ZLrR/qHILYBWSGMOj4/4dBa+GjB93vFeoarMTm7rmCYNoFGPXz26XTlu/cbCO2zaOr92H2f9FDEo
aO6a5TtFofVLdkQTteS3M993sB21+lrDknis5BTziA3RXdujVK4BuMUqpmWQ9L0xI06lNHIfqY2k
HExa+0AJvALgNSiEb2wmkY8aujNJxE260wLzUlMwJCCpNsvWGefSfd1+zJWnyoBZYKjuAf5cJdpb
VLmHwg5ZMzCuehvBc+6x1jnIVbzkMI1Jse7Oos4/w9bksPyFRR7+K/Y67+VF31O4FR49zmWuClL8
rN0SRje+1sbPMC6uUlfGxPQeoRJrYIbjapqLRO9dsmI2XVr81xPceHVTl919f7dVx+lT6v9lZg82
ciMjvVJCQwfPH6UUvmcXiQ5u8acTZud2hAEf+oNLKvOxlLi0WMGuJvuBXIWXJsMhzasToMp8rZHW
3ktOxV8PmGrgjVR0KHUC8mOcJLpwb0r1RKpBlaVEULS9dFVbNjVqO+MPPSVGThIGdlau85cfdZbZ
zEnwlvU6gs3CP9wZhRnJuJOynO485MuwDjh1x7AdF+TL6AYqWlH3kxIiHd6jDAFtGGFG7IW5tIlL
OG7f2vBgHLoMMtLRWcinZ8oSOv6L2O0v3eW2T+IkPeYBDekxvl5EXB4k8pFBVN+IFlyASi185MNF
7JElIebXUPQP62/gOtwqi1mgb3x916U1nZSvOsRgHot2sIMx43RhWV6XMr4L4UqRWvomHR4LKUKP
9118mUdU6BJcmYzHla8fcoQlRGzQOW61+CKNXNPo+Vg9fmpN7iKbyeBvjIIZoKXL8+ubp04RCp78
Mt0iVd7ykgtSFlXIwRzBC2mD8XPTZW+6Vyz3Hj/qF1yhD/jib/uHHKoF9NnlX8CjNeRo++yu/E6K
n5WkgIv2ccaoLUE+ZPWrSIx+7k10+YTS5d+S/uFUEuYc07MuwzxQZRNfLBZCtK/pEXbDYsce8mdv
X27OvfZowCZfcFHC7sBwRAM97QAwAxwz1k9fJT0tvfy7OS8aUWGjEOA5hLMSf1RmLfYfvELwjYz9
eC3CrQOWszTzU0hHuE71ARp+JioL0a+GP8fuAp8eWupi61OyptASra8MdNNdCRbQOmGEayjfaIRG
6W+R2CGIfN45oTzAuNflE7TB0sylxEdEEPpDHz+S0IFFjkU8ZzhGEMF6dSZ21vaOW1vP8IZkjuq3
OxoF4tfTFXDZxs5KjAvIGn5NMCvzz+cvf4QsjJP1+NIl8NtHJP6frAK4oU0jC4kjm5OppNhdEv7/
FY0r9hw98JL1V9Hl/EV/9rB3wFUYJWWihPtaqzYCcrdIHHdInvIswxu9d0R3RSj2didR2t79Unid
eXe1iK8U1WosT7vQukIWv9CX5VkNAT479AiUYJtbLIgCiXsRt3RWB4QN7Nu8RFJNU8CE8dHl3KeM
8zkWD2KgI3BmHkWLqz+4YapxveQV8RNUMVYgt9Uu3OR8c5Tm6JuyL1Fjw50YlJenJsxcK+X5vUtl
HqSE+bgwctphAvvxRPC268EZiSczmw7pMnW0Sn5R0gXFInW9xRN6Otb0Yiyh6gJ/rjpzvqGXHwLJ
RXgekmx4lJHqKdNQyxqAqAUPVJhSbO+kCryVHL2t8jCz5nocUxLxksRvU2N22/SWHapOkyyCbNgQ
bCR+/qCwc7ydUYyB0/DMzWAMR0D17n2CszDCOE4t/yc3PVY5C/iXVlU8ykpVGCmIlsTFKsWdfoAk
yYXBu+/VS7TTOrst3Y3sCcDRz9Dwn4c8xk08Arndc0aTNNisNVE98bGROIZXvqK9X136ZxhA3KpX
koZvbldT7Y+lyfVpEKsiq6VmbFJtb1O0vKgJmxb0KKopxU796UNbeh5tszm46XbQ0wgps5wxgjMi
Kgla/VM/dgW6GpwBcy3uHdyxHOOBhF1PIxVLrygWmnum7nRqjoKUcx7yrCKHOq7Rjvlx7B5+p4Hy
hSpxG5dsibNzoLAxbvX97vIdqzoPKJyUK0iiN14AOFCN4wDhlZ0ybOHIOKPTtx2bsaGO6pTD94m7
aAOKdgHmzGHt3UfyytYIDmmkjj2gpjrYanydMxHBDHKXBhqRjvW/ZpI0E3Nmn/H5WRnPkXRyShcw
PWJeGaOaHXCUA0AmPBhFPGcyrokz6qAYH29nLzMs2avZ1YenjY6g5rEWoKVWrDmKY3gPHrhIKRhG
r0YT5cj+8+F19hwknGOHzA55+tpekEYWT6O7RUPBOUWMicD6E9za3Bau5NX3pnCk32a3nbrt1dPx
loHxeUEqnTXSkasDCM57nw6GTipiZOihnSBehhGvpo9qTlIZUtn7d8v5B7+POAIB4syMOpr4ASzZ
MRNyEtfgrYT7vkpQr7adebLK3U5ZGwolr0ZrQQGB2FWzcBzR857bib4nu97Hj5OKQT+hExLw2SCm
e6rgALEQmNy6TcReiUX7c2SoskWU/O6e9+LCOwl79+veo+Uum1NmCku3ZhZNkcWvD+MRId+C1DoE
peTTUsXNhaAiLrB4i33Gk+lYS+J3W76jp+8iAoqtJJMrZVpX6E8wPr5/TiBlwQvNEoH35fZw5EF1
0MUItIkzP50jUckyYBeP//gjBXrEXzgo4hUZAZLmq27dxXcGOs4+RPGVnE95fTN0flKSANzFT4pD
F4rPr94zJvpBAiNpYqNM3guWIsoRkiAC1ztRdqhSFKi5y9YQMfxZN0NgL1TZr1f+n9uQVWc9niGZ
obUd4IFCR9ciWnmoVkmkGBLnm4lXOsBf6OjVzCd9sWXmELFR9DTVQ/0qn7UjeEFT6r6TNHiBlgxU
swjDClCCLwShYML6Cwxgdzw6uKarrjhCD7lUG2IIJd7Rxl6vbilX+NThBVJq9TVbXi/Qs34C+2e7
zKVwj3GatibozkoKvRdsylYReVbc6qyi8tDJXTsV9yoKnAtXl9ZI3/7VmapYEYc1cf5NKksrZZrp
L2zA9KyT0/MHxn0Lm72AtEdgKWoKHezWjgVBXrbmsPi9KRWJo0ym8dkQMPEY/XR2R+uFKGPfwyrD
xu3UT8dPWLufRoBWp1OL0ozt6hS8w/Cwj5VKiBvCpE6I7sbOviyv8Sl6ojwzpoct+4KwW4zqEmCs
yekUmzpgIP+EcxDl+mKPjYIIvAv2elHYIaLidrOP/7XTEyZzK+rGjBtjtyWXje0Kw4K6rHoC7wo1
jO27PDphb/xZdb7D18cmuxBW7BSbVnfaaVLElAwhmzSepYZWQBUF/0cCgbZlVfquBsKODeyR4nVA
WcY4Bhd/5CvJxq0dNcD5Q118THbcfcNa9NrR5e+l9vf4xF/J98ybvrrAFd8xzsH0OWezdlpSjRJY
jIULE9EEYfOMKbXkYeBRfKnFctxdRkfXx/UMGSuTkxUP7FElpnwmrPLWomoUct1NdN+H/BCakyYo
gvBPgMM1e7DShZ8cw47tBn+HV4+MBwttURatswefFAUb19qCBSKhwvuEGloGi+T/5V26MAXWdrSt
jnQe9eCdRXlIv64hweBWIOWW10gkf4SPg99nnfJgomYiChZe0e5DI8a7H3nKRzG4xV91xyzK5aOG
f4q392NEpgINdfwyspp6Y1JiHLZr9rNONOBAzS3Ac4XGvSU8wqJ7nSy3QS5M34wxxoqonN7t5q1e
zb5nBhIzvEStp/CrTs6wmGMUHy2uJUPLcNwAUT7Ld40HwmC6gwkBUc8z9Wv+AywAN0jjmGw1NeeU
LTsJ+d+9SFcS5ez/4cWD6Ub7QtanlSidsMtOCrWjozpT2AOskTkoadnoubwcrI2Q5IfPKCbqQp+E
tlSN6zk2gaZRmHfLCG0uG1sqQC8b16dErO7kfXolUs9hEGLA2W3gHomW720UTl1H0SHs1GYMD5aq
WyNIKHa8KIF+po7etP5BOhzA9SeBry0fToVzG8BxpUmP96QTpkR/5dUZih2H+J5tYCHsDHL/KXUp
wwacSTBbfcLAfmsXLFgu+IAPzDWOgs/3qM1BKFnnFTolAYCW2xcBxOWFYcAo05TPM/GFMiR8kHCv
BuCa+G5NId/ggMXpDmnUTNvOlGOxnt6FJYBNBtPv8pJIh2VX4HJdTUjkEaQ57DstwC+UDwVHDgkl
wBr7aD4JyT9TqixTCRLPyyP4EDsal0b+xvSnt1U+1BPVdk+vII1QGREuP720PZrl41AKRvyI0eNx
sVWESajrR+wLBeEgCMimmh7yaS+0MkY7ht/Z0p0LVniZHWNAqTJV9FbRqLdQeKQ6QzDbQf8dJRNN
PYPy2N91Ziggv+JfjagZt7a4bWnRl9Q4gCzcW3C2yWgqP/OoK20bfR6hlJ7CMV59Epe8FR1dhKwy
qMUj/KfA1Y0EwQLO60VXoqg/bIzxTD4XuxuZ/Xzzkt3Pk4JD+Cyx618FqLBtpTqKrZkk7G08QVnR
NZR+vVQbGVUT/q9vEIWonRncPmJnQTedzn3ZccHT2MihvxOm9Ex8hC1eZ6mZ2NQAVRUcoN/TpEa8
0vNqhRVCCLeul23hGE88aw0+JZlfcEliFhAvGCp/VQUuY5OOcKRngTuAQynJ9SQREIx0V67miovV
k9BnEXajK9z+atJOjSW7n1Eu3jz/4+HO0fg6m4+Bl9ecRn4ku2gmejjP3GZL2T4mM6lgpx4i2SeD
QgQ11708rEM3PdJGY0e+RjmBeAFIgcntVIjaBBKbDe/SaV7oq2/JT1gv4kjY8HGTbhapRkydFOJd
G2AhCkm3CKmH5KolqgehTjqj3I6wJnUrRWJ8lySckBcfllkmO9bBrCd0IL5FD2+yqLHsc7qbkQdx
PcAZhabtU+0+VZd4Fc56YLeVPx6zMOaT+gCPXJMiRQx2frshs5RnU5gt5WBl7+7io+vpzSKs7hMw
XPN5s7D087qkBEDKS6ICP4xus6HE3Ru5r1YL3DT9y/X3thD5+/kplYiljvSN3kz4zUmKVgeHlDPU
1P9w+MuVT0XHrvTk6ClEf5iRTgqPY/nlZVVCJnnVGNRFtIoAeZhTGjHh8b54OEHBKDWmZQfB36eg
HZqHmO1KdWDH0tQ0dfvBTIi1R/X/WvQCACr2X5KgJrK5r+GREj2JmiUpHMDvAFdHBVKvWoKU+6kK
qeHecQ53fC+eWeyNsFPhLIoE+FCEMjaVcwehIFqM9n8ywfS/iG99oJtN/AVTo+9lL+48W4Nz2tII
hT/K/J7PA08Puz7TMJNVWXcWuneZJUQDoUeA7M9wVRtm3m7CkL8wdjhEb4Opie7y+E/MvfJwogOY
wlgi0KY0Hbp0H9H45cr32CVgLqJvNr1hVi7MmV5Q6FsFFt6y1EpEWY8rSXxJWGc0PVN4DDkXjTp2
O/5MbNU4aWJdFVvfYNa80L7q0zKpRxCwSv1cPx3tvqD3HRdGWqEfgZbCyQKRwt34DHNyYr7+YnDK
eHS7W7WEdNouRARsADYaxprxRAJR/7ncEtZiEOAT2boodowL2+kle6vGR5MWDeN6HcooP3gvKGdo
Ap0c31shxZgbvxDyaFLf8IG1v4UkYGDGXMfhuVxXq37g/f6jGixBB/qU/VRVRo2MiGPOSTaxO83e
bHWUcRVxdqHY3MKsFSF5B4nnjtUNIhI80fW8BnFKK7k0BwJI5w1xgmA4lCDyFUZXym31Nk40jDFF
WQjwKYn383PlX+qBZBAcIjFlpZ+Jr62gwF6bByBuSVQy5z5N4HQlMrsURk5iXU/xlgykBJdkWrz4
DvIMRjB2hbRjpzToi6P7alR9KF8ingqLofq1uD1b5i0IeF1YIszhSX+zGMxZ83YpeZJVGerjLDGZ
sNOMjCoqJdYCNvkteALF+EF4v+34s0gz7F3xOA5iygSLDp5nKGKEJ7xRk37pkS6oduU9faHOZ7ne
2crFNHpOUcgcDPWcD2ao7AJxZCiXOdtHFNtSTodT4bfqX4V9seo0j8Imzhvi2FWQPdcX7Mw+EmbC
M4JDTrzXlsd3mxw4wVkf5S8vCzkVH66AcII5Y1FK8YyzPYIOMJGveGT3KVqk1OSXL24lv6eBsS5e
Rx1ry9XP5t7ahLJPyhLIUBOXk78j/f3nAxcQs54G8CwZn+gyq8C7JBNtGq5gZQMCWezQz1Tpbo+c
jB2wtOx6Izp3vRpN4KYxWs0p0MncXZSVVFiZ2A7hTzscuSkxNzUBNLiu7ton6c3Y09DcGQjJiBU6
DJ4dmuoEWfrAtUBW6550KKophmKBM/PtZkPnN4CQn42prCKgpg70CeL4lkviP4wb8mwuLjAreN6n
lnCOQHg/OHewuEPC0S7+Sqk6RpfShc+HBFbzK/Td6Pl+gg9AnnRj0iG8783F90U3n1vN4QXVmQYb
uoZ6jH6yTaqlu2EpNSX3+NffeXMfS+0yB83rXneltDsVnhfDeWNOWF1iD9QBSyRQxQU4N2OnGR37
4PPJBEHU7YMFUU59p5WTTyiJfBxDxLJAbKcNvk++CcK17X2csH/x/Hs3E01+LuVKyiYcGHNitNy6
k2lhS7FejiFearEG2yPoYAWyvoORpv2jv7rPSszZGppAXHQzMORZLtKJQZjZKn+ffhbLYYI8bnRc
ZapZtbd08yygmmGjDcl5QsaBTNJ+E8FphjJlessGHtrA8oYQ0vsNQ6bPnMZ5IZdugFggnbm2giYe
ZhiIqGfHIO/+xDgtqqh9Q5Z50Fcv2QYt6BkFTDZ7mnJi13U+m0B4TaKqwaCYI8M3nB5kk+ro45nv
Ba0ue0SctRO3HconAufU+hrA5HfGozjgiONZpDqpkyK39Ycx+l1p6aYIzfj6A6aPctxt5As0czlw
345uzU9cfot/NczMzzJKtGOoKE3QaonsUtmCUcK1eLVhblt51E8pz55UmbtTL9nplv5DAhQj5A9o
aNc40zxl2f9Rf5y7473GGYwp+uIiCBGWOb2rS0cyDi6AF4YGf13187+N+JM+XsrFJ1kgYZ2K0Kzn
LfSIBsIREdQTrbt7GcEc+Npjin/NHo8HF5P5CUh1npa0eZ7vibYUmyoms5bLLSyumkddS0dLiRcE
u+u7WLMo+IJPOvxCxJPk60JWwP00UsluwzZ74BDcVPXmmoRJYmpbAXdYQFRVCRFwvcz0CsYXeuNd
JU+e4XtBcTvIldOh7IVirOi2Xf1Fb4teEtGr/EbKvhrf9D68KsAJ1z72QMq0BlrYrZyfBM1HL6ot
gIaWjIdyrygMo4du6rsmo93yyKqTQ0JnEVFbUtaGiKZX7WSR6cmP6KlAzU0b7jzgzkATwnSsZWVl
d2j9pTgsiXhF+NXMxXaqFk7Oh2pK/rHJUSPxeYfZmQh1bMwhppGlQCpO/uiaYFHdBFeu1i1U92tU
hmk5IuCbBUlvs6Tn2TQJ/iOWZfsSxWTeCXsK0Q1Vwi+h45V+6Wn8q6fQjMkzufT4qM78WOrJ6xbn
G6+TdLLDU6nWAnbIDzEZmkFbuTUJtwoNDHVGaOrXlr6KNzmleOTM2YGXQZ5DmRlsd0h6LEvjJlpz
BqVlTlGz1ZiC4r1Tuafgdo3z0AKpbTWsno7tXC/ZxfzyjpDcGYaCyd8zlU/6Lp+sQsMfD/pJQOH2
hgQ9BnrAhMpX5oH07r+z0wJ6XXb4MPmaJSoAiYlDqjfPW/Itjd7+w3QBY2N/vrt2UME6Xem0VbyL
4HvceLjckv3GgkMmNfJgdXFN73K1/+94PmtmMvG+IOgzSpAKE15Ee9L5DGCqq1J5JEJ1nM4YMnDG
Td4O7r/2Lrzq3tCrfolWm4JKB4hlM5hbiD1u3MZB9breI5PmX4XRNdW5ds8GTHF7XSR+IyEOVYjI
cSFDfeYuh2oz12RSVwYJJFj95rR3DpcZSOlJczo5mLjukvmvc9FFtkvDpR+BKb8bVDZ17+DL6Nio
+34YB27hDeIdIfSDvJRG7N8R+ksFtqbZ/sxSKZ+kbO7tSVq6L5CZ7pf3z/VJVvhz9I9NXXQKyhUb
y2BfgUcJAOI6QyMQg9CIWOedeShV1adMdRGfxKUyosGAYSLZx6Z5dJaVnVW53d+iPj0dCmveUTRP
TgHArlqemR+VqorivFJ43lCYV7oBGr6jNIY87PQ6Up4aIrWr0c+N9xvvrMiD2pf2SEHX+WrGOHdX
clkvU1MzhueihgsASpxWCd8teHLxk0QFUds3z8J26mSyz2ZSewc/qISgXpZ6TzQdYPIVKiZdP2qL
+KhtEOuGP3UFya5vsKGZnh5b/boKhWVgU+Nxa1Ur8vaUEtwdpVCMBnoXOIWArexmBAUtqqXYO/RP
kCPFRrOAVDYensO3Tq4L+1NTrqCV3oveqzAk6VBOD4chWIFPkmbNUL3ZpgxMdopz5FE2EponwCGH
pXYzVs7RDver0U+Et3RQTabXLb8Q+48sq4GDnUuYeoOonKJOfd+m7MRevwUGp/u6Tx7TmapHoy3L
8lw6eLG92yVuUqzsAosTyy4GMSFBGw0NFkh2WKsOKbW0bydIEiUngX0s41p347IYf9ZE47Tg4b3E
m70hAqjFJAct8CXD223q/m41klotS3AZZZNNedqXJmG8bJpVew5YjDs/bU8hJqtX5oGtEtSWHZ8Q
vLLK2iRquASZXAaeHUAy86kYtFVu/okrcYEWZp0V+bwe3VU/LbeeeN7ag1dC6RfndR7Ihb6SL6hn
Vk6OaBatyuaRh5v7jFzIwh5rJzlBn7Oz40bpMH4e40JqptqvPdexOdUywXP5Yai8YSGdQxveEYay
AES4wYJNOJkTC2s2bJXwJpB71nRTzRUA3TRqNAqQwJDbTrEwsohuMOJZpUtlzpGTxNDyu/PigzZI
cnEoYOA/Tyw9H5dz5rvSY/QrDfL2n1vc+hzh4ln6LHeSZtvWW0GyBsdMnbRqySJKO/rZjHuZtJ5C
yiWP2gl/Mh+03G6dPrp4vp0bHguBnDQnIeLg7sOZodqnnPCI6WVP/TDBE23F1L/42oPKGkhGr7wI
tbGwn9CPN9STngcC6+AIiwjZgezvjcs3JzV/Q7fBYDFDs/utsFxcq3gztk+t2VuCPu1ObDXu0cbN
Tf/ea+XxNYEIrvf7QaFa5f1mfLOQ7l+5Je9rHoqiwDioyzKP0p4F5kDAfhh2ydwn+//jYMnbhAIm
zSCGLrgZWJBHkAk26R6C2WpJSM7CaMTa8uvTzwQLct5G31cFmiVlji1xE83gdyoJ90+0o4GP3dwq
2Zob98GSkH9ywfnEA2C5PhlLPxmAlhBsI0cVSUsVt6+oqtukfmj7MGo312IluGrvXDhHvaBbQs8B
i0QtDC497/PspPrvwLL7fFOeDheO80DiQsenLclOpLJkYilE3Z4q+MTBM9hkYvJByGXFJ/PZiFIs
MTx5H4VD4MT9oGPgyaTb1n5HTfgqZFDp/m64+T4SQI/rqbfIDv87FxMyXi2aPe5dmqJIT4ddLSZA
23YFMrzaQ8I3u6+aCMJ5DaqAfKDIh5yItAumFyYD2Y+lO9eL8i9tMaw1PXlV2qefAAC2a21Xjxbf
OvtcnWA/TBFbOrJuUTpU6N7sUPwoavWi/LsoA6stxYbOG4Y8f2w82rGtrRFazS1G19S0c0tTCXjX
CYMES1v/bq3cCksrOiQ6IX1SM+ZaRsz7+zYEOJxdWO3aQ6Mbj6CmgLXcR8zaT5L4pYQSMMToSyIg
nJKcL3ixhuGRZJ3/2IxuEWiGhOBIXuzmBB+jJg1rsHJowNPyXYYsZGpAxDk2BsewOIaJwlklhXyT
kDIPHmeVV4VG2HwqRMBu1geAViuHu91T7uQmNzbt3sPPCFGvNS1VKoSX7X1y6/t4eBVWdD0zs4KE
zfTms/nSZNOHaku1EnOfNf905vpi9+aDBleRwuZKhc1e433S9eBfyf9Cr3UfKpUQt1s3+ICGEle1
hwsOHrvMUIWo/2We2up2i57RiJXtY64zECnR7pLHlYyNPRv9zmeKioLG9wyQGTepBGINFWXO9znd
8ZDRNj7VqoccZ8s/ozLYYgxZzk1MxVID84KOepOdT6Z81Z5BXMEnwopN39DL5bFI2My08wmgXfX2
rZ3S9k1PpAPeEfaNziDAoKa3TD7aQYHAlNkGEEAHNgOoT/tVyQV9MgpLMFw8NfYS6Lu4sxppBM7w
chF4//3aseW30NOX6lOboDT3HJEm4dYYyCW7At+peqhFmCkzwnbFVijNzdCpwGTz7D/nCorVWx/r
jXCLHQckG52oDuoEgWxlGp2LEjUgNE0H3QC4Ubp6ZGg1dR4mLI8FkRr26SnTal5/Qzx1DSB3bIEN
0xTbkuAmeZ2B+Ecz8HfB1IhpkqjXrOJKlXU14xcIuaPa2QgdV19vcziztDMtnWJCZbcC/ixzIb31
wjire+9GwqA22HItM5mFaKe0s8/tlvuP+rH0id45Eobw64zaF5W7nrOicHvOBZ7A7VlD8i7g75Ms
WnFNCSWD/nJ7N/2E/q1I9n9AiyaixuYDQnXE3keys29L8dxFShJRM0EnIO1oplvae531lWA4UrLn
cMkWoOXsal0v5vyS57ayivFPfjmuerasOuvcrKkAq587f1nncKJuPpl3nNWTffLtGkWVn5jKPSGb
7EiOxae6395dhXxnIoRX1U1gcCQnxbJcmgbk2b/L2q9Xnj8AwS4LBdC+MbtzTG4cDVHq3dL6PgX9
qk1+1UvbDmsw2KYTmrlIXzYLp4cEAaiqpE70LeVpB9CCXo1XK6gtYNUTz8aDL52JAUhMboGMcFp8
94aW2TSvKOPUWiUclhcMp5Jcgo0NnrdptmBCqCjCfUR1pIZbqxSVCLFb8AkfMix3U7wEBsSbQtvY
AVME93LiehQWcoC2goHMTMjFNRn+Ch1nG7dbaMRFX20qWyItBoL4BFcaijJACA1W7cL/N0FKlU/L
zUo5b4GFWyqCUhKyhYiB8cZuBIpwP7OKcm5MdRrsna3y3u2iOiKVngy/0qI3NaOM28GTzOUFPGfL
zSjdcua//M+86He7tX0g2K1BdrjdccUceLsjHd31kbAtOmZxAc0ZOSTdpKUAjDxMbLoXgb22uiHq
09qfcsDSX7T3qQ6d5QtTgci8kp0aaRpsjWd0GXLT5pBLx10ZeyWY1csCyFeh6nkTx3d2oc/wL1aT
1kgWw0u1v69TQj9CV1p/5lrziSiAaoVJQcseJl8kb/uSjg9KFipp/zhCbkn6yjBm1bCtpeLrhV2K
k3GQIbWyTMVtxHUkmofcE1xXBC1u7l3uilTguPpryU51eWfWubqh0uhN8EK+saU6GM60uGYN1gg9
m2IwD87mUADRO1im6XU5oxJ/wZfvYtgcUyynTytImlGM1/GOcnsbacWg4L1WZLUB5Zf/zI5jgNSX
HZqpuqtQ/xE59D5m4R5kWEf19c6Ua62vnonm9u5dWT3iIwszSh3Yj90tfmFI46Rko4N6dxHR02SQ
sb2WwHL5h7ubyKDANySycX+O+dWI/el0mjZdR+7gWwxSl+6xkd7RDMrYB07tmANIK1efTi97GjRX
r2pVI+9uRh5Pb37jZonJvVVkqB7TOuECMgCX72HXIiHEkgwO64b2zmlOLChm9KakLwewAUAbfu33
KVfs4RTXpm6Kko0h9a0hT439J6Ns8mBtAkpPwaA/HrAIgxfy8y5ioZoSNSYWC/wDIXNiZaADZ+el
m/1f/nyeM036TLkdFfvc9hFqPtGQxXYU0Aooe128YBsNVvfMMfBpv6Ff5SBWaieSDOmB355EeLCW
P8jQpkr2+D0ACYSxr1dLJjp+5CPA6prYeyXTD3xLRJ7EIjqxJ4E7UNOiH8ccu3mHnaz7Ig4wH3ox
LOtqJAf+rvbQl4XBtjedwQaw6YU2lA4JD3TLwb5pQbeVDH7BluNqEfuiAICprsTyAfEJTe5I3ehg
KbpT/e6kOr+NgbPDWfXKUyMlBUc1Ok5xYoqh/wMFEe4LZQr9p7XeFP46LGkanhUyFFlsScBEeJmK
uQAliJ/c0eDElHGt8nxPWoX+ZnX+oWpaD5M+fcFB4NPEsYnv0uAhh4mf1dZjeju8/l8OXx87feuT
0oEnVAFftY1dtejc2e/qlFkoK2+eJ3oxKxk+mzU2B3NIYdxPJUWk1jesJEJouI5Em7q3z1uy96bU
TKV+eofIk6FS1/deY3F9WUhICzaAVCTxIInjMfliQZza2Yg3JhJZ8BeTX45LVHEe8RbdVdhdJ8eG
8mwm1C3nBNGF3UY08nI1FrQXTxRY+3EA3mwPJBmp/ppu+6M3TW66z8TysXQDrU87lWncELFYp2Dr
ILAvbfpf5DQAF5lhZ3IfDits/Uo/ndpxN2VZ0GM8gLxFJsmQeChvSYfW33Qf2ZlLUsTwwbQ4BGOr
ywR+IGyy15rgG6CZ8mM8N8b99cNV8tCfmNvTBK5mB2/3l9CN4EP5VhH4CQDClK5wX7sezGwpejjI
OA7Y62j1WNyS5b8kYH4WbMOuoGOYLVyTFjZ+QWUjuxyy3MfDk83iZoTScoxZ9NFPQVS4lqZnwaHX
uPByIwWFrKJJhEvWXjz8VvOYn0eiUjHWv1OJcvkYTlyMuO2s/jR40o1xz/FFFvIYtpz8tCghSx8n
1evsa9sq3JYgGGS/DLVuG5rYRcozdsD1LOZNTB4YZy6YhPWZbMTbFbiwg6noeXZP7ZXH5ggGSQh9
lZzMxlgXqpMQVH5+Pb4CRYFxN8eM8DOMkEUthXR71oD/TocQYUDIapFp7MMuqkFawfSyG+qHQpPX
ED86s37/6w+V/AWczkqCHilFMlQ19x5IX3ItPoo1CwBbv4cFS84z4N3bZxnjYF+DuiKOfi5jm416
dzXZtRVEp4uw9+ml0xB5Y5/2jZMXh8TO+NOPuBmffN/bmHJFh4jGkvVPfme+DKket3pMq3rN1YDc
nBmo/fZYAAUvU+51X7uy7R/m82+tZij2Avin/LcW2zTb7k8ZHrJZW1YdWmwfLfceQgTfxTnUNnZK
nytzE3aPNIZiwqmQwLXXDjdhDSJz536XthCxJcvPRMkPvFy+XuxjjpJkn3YYWQjgcNMs+NM7btPy
laztgduad7RIBFtNfjIGVRC6P3JnwKCiXtBgfTUMDDam156DLRmvQLJj2EjWr9zfUbEawtbk7C1q
9pzIGgThWshxAjJS5ALidUsMK4pI/EQptCJLkhDfg1FxsKitEYM+SVWP3DBKeoULlkcCSjiKdELL
5cxaVUXACprh07jBBGiMBXJBQ5Ub9xPil8aSxtAaCHAWvU8d6aJ+9l3hSDdu/IPLgtdYqe+Z6tPp
2Q2990BR+D0PGF2uhwh2/yYnZVNl3+4r0FBGzBghop6pTR5XJWmMY+aF7nCWT6SpMfEC4NyI3cG5
YV25kujrCBG/skPok1Bm3wTsTUPviBNBdLVURVdKAqAPs9h2XvIXR3UkPLVs8NpKscr23Jk3JTu2
R8F8bVmV9BwL+mCNFNewkjtVsN/DO3r5j0vLasVxzWa4IlhhLPahCJcs/oQE6g725aUCeRAlZZzf
U7JHiYDfsMEsGsdaUrjJVcOtheTKwvC+LI/4cJt3YA6hYH/seydZsytyhPUnGRsyyEra/796H10L
IjxZr3B7Q4dbUNAXy31oDuYagSLBC1Xl54H0uJgzOD9DLZZNQHzdu+5QgJJFpfmoy8zkC0Bq390W
WgcMwdFP3Vh2I5N3a5ywGREqhhJQFUzyPjD2g3B9HvHDwHvCI2OXOAAXcs6mPWEw3dO+t+YvKGpr
v1pQXynf2XpKPRO38GqWcffoZ2YYrCiQ6xJ3qZy/xdAMSBvzuRufbSgMXd3GvIFLK8KNTuEb7RoZ
XU53bdSFYT1V4RrXef58EG4pTea+ZpA2scz/HkGUFnazTWmL+SIvZosUZBAbPLggLyWpabtSh0Ci
WJSRttvn11QD8kCXwDl2zzL3ClKx7hqSgqdzWM91VSa5KcKVsDMOi66W4lCr0xstaSx//0dI0L3Z
uK1b+xKroTUP3kMEE59x5cJ9076Bi6Ws6o+pzQvxBa+qOpMKe/pIbMmpRVwr4XBjTxhuyzI5wlVB
N80yuXQKuO2m2GMB0WHd6dD8C4/tJiBeNO0uMuvr/VlzBRZi/PwtXNMSlVbjq4nQEShlYHZG2o8z
5vppyFhGLShQwUeVBxMulKVcWHaFlsVW/jP//KYEZdXu3LRymit9uL4DY+wR8uIrEoEDGNnyUeoi
/lcOqOf7AivVn+vFMM7UwafDaBdhWUP6C+9w6qulR0kJxBpsUMJM8z24DqKvbji78ohozNpMFsZo
eHwB7mtpz6TIV2teLjim3iFYVpC/LDLkokNbDafykplGaCFQt+XTFbVOl2lHal19ZNs6inCL43li
+HrtHSg87iUh1L/wcdMFB0OkGzJBSbnGoGM0de0JcjR/7RaSA5wQByBfdbl409G/6XF/IvWGSZUy
ZYrvmMMW93RmIITPOTEiwAFfhccuiR0DSjvvU5P+mXudjsgwsL1IXk8B5e+t6Vw1KVGSAcTjMms8
z2oCqr1oERMfJyYFPvoMX4Xe1LBisKAJNAt6XGvcR9BLYtYpSKfIiqwmqLwTU/utUSGWfkYepAWK
EM+rwK1b/NDJiXr2jFNsvU92hFo6IqNoiObtevarjmNcXmWI2n9JUre/Et/+okjALegfzjLU4/s5
YjR9sUAsjz01ZXuyoCbgH6ooK7ck8s2DwHHk+5VvheGu5H82tERFkLkUMWnp6Bw3Y0k/B+z0yinF
sm4OlBNvc0c+cs27C7f6KY6tSJNVFziRanPdnoSRcgRAYK8g8A18WrxNHvI6Y/JHFdDtCcTiXdz8
Rcta6+NhghfBqwiyKbw0RjquUr+9RMaSZylqZv3NXmewUh85e7YQ+8mIEFLmMiRHOljHsNh1pTL+
md3Exoqx/wc7YlGTI1lFq7EWoCorBBwF/A6ocxm34TeJr4ncyHx+7VQ/3bxPx9uQrwXXKgUR65Mv
rLEC4j2WWRhMUpbh2JrzM4aDY57WkGfEHduavWrhFKiBKBqyn2MqIpN63U8CCEe479oJ1S6mYm7M
3eiCmkTq5ifxk7uh6HnJ1IVAHoM/ozVW8141PXqx3EO82E9LU/tbtQ0qdOmMSfzi+/Bg4KrzVuF2
3g520K2dClZykBmDnXxIBbULkzPY2e1n4+X2mWz1gjcV5Ocu0Gj6VKgm4b1xZGPNO5YtA+xK4uwa
VsCx09rLRITmkajTZvI5TcNJUhRrxeOpXpu+z1JVX/Mdl9RHRkyGDXpR76VIAXA3EtCdpdn292CF
glK3VNFo8j/WefmwD2O313v8DxJ/xsJuSUfJrScTyy+KJC0VQ9T2BkN50bjQh2idxWqFeaVeJz3q
UjfjHl6wFbpiGQjzshl6nmSTSLi3cDyaiOnnP5JEvk/Iq5CTZXmJmlj5n8w8xShesivlPGb9S9p0
7/GIqLwtWJJkMiLdg6Ypb3/NxcfvsmpUTQn9vthmwtTKFhkNL01R2hYYe/g7oQhy73+OR0/0HUoX
A0T7Is1rrzP+UaRc7+VgqcKRYmUqcJ4HouU1RdD73uF7vmsc/ZGGqP6CITt/JjQchRYYPV7jODyD
mxPH6HnoiROngkBsxe/8O42RsNorW83bJ6eMDfmWbuZtGIgdc9kIKwpiCAS7o5030l3H0P+YZcJO
XWjiVXFLwiQAR3QFTyp/yBsALYRzzpz8w3/7+wIEvyciA/TF+cpPA5s+sf1bbZ3nT5QUqZo9PcFO
CKGcXXzHeBlwxbVfzwM+iahlSUiLuM+fS+dUndoeuJnpCqpRQAlUlDoo9XXWw4OMWXMKxfbUz8n8
YVNUjBZB21TWDl0HwXBwxchNPQaBGMaSCzu+usDFR6cKNOkBWjRVVFTxdhw7MoXVcQvYlvdGYoyS
GW09vRgCZij7rDJOt9pqlQNR9sfsgFA8cogg6n/qI4XEkJ2HESn4ZFnNJEzrRzBOqLEHOvAjfjj/
fr2g4Kn1HIsehxKVJBlINTVHuOQEUxRBn+bYRNSehjIoaDuI0GSdBw4rRHDSkBIaLP4H0sveW7/8
x9fLg+g4svkAuEkXqEsoo9wU3pEksELWKBKuaBu9xCcQDcaW7BedOSs8s0MfSwkVam05FoK6UGy1
Pp1Llmt85zCDoXPxYNkXl74xqGC7B71K3U9adumrYMHkt6QSJFsCPzuzCjJvnaAkUwopx+AKFg6W
nD2d09CD0JIFIh3m1CTqK9AlYiXZIcQj8uHrHEZjmxw6e6q4Monla5MPz3wVC0QRLxIvWK4b+ufK
t8h06wsyuvnVrhpVGU1a2EElJR1c/UYKFbv/84voOrW3DyXmvxR6DO7QQnZAskoxtqncel/ZSZHA
Tpt28dDuxhhXONGth8uefSNlULjUdPQzf2yHllG9N7HkzMcXaaMMpIxuM6of32aklGJmtBuLhdgP
kcvN+UrEdtYnVzewtPRnolpLmezYbDYdJnDZdkr8fcUVbk3mEPfOj86vtNmIb4qjNeioz56EZ0Fo
W2nRuDgqsGQAefgFkJoBZGelI60IVkcL7ErbQd1aTPGEMNRdHFHgIn9J5hs/d3HLwn/Lq3XlvVtu
CINKud6cT9icNW5aLemuFQDnNyJfdVz5aPcRMUyHXzlfENfOIW8vmRKzptOsgz5Zb1GYM6XABOYl
6Bw/hLLyDjzwr1mYmrP2ImqIN879jiocRSTI8g37MAfOCb6NUG+ZTfba5YTdZ4LMH6uN+r1uLRBA
IDjDY1KFEt7UV5ij3dxcbkji2psaZDjokuZ9BB6Wjd8VgVweaSmoTvafGtSxhziEfadDAUElfsq9
MOeuA07jCwu0wkZkeoJxpy0mCxLw9HqhyOlkYA6/P8XT09lEZ6ASPMchN607YbeibGkQkpWkDwLb
Ugd4Xl745UWC/S9YwXwtdqw4yUnSrvaR+VWzNvp6g4nIIp2e24kvLIIvJNRCGxopSp/lThuh40/2
PojUvikfCS8p/lvHgLtmZVLBcAd11mbYmQHu4ovsXlOjVPGozF4Rbqm4u99iV3xMEpnxGBc6PVj+
XZo7JqGKMfDdDNF3BGIJVM1dGLDciVTOy0P/5+vDMrldd3ekQhZMK+UUOy5JzyljOSG1CcNb5RXw
it2oia56S3n4zWHsVNZ0pgCoSX56cVqtCUX4GPtILlB+2p3gN+/aTlxmPq3pmajMVzz91ThSJs8R
Qq7yrg46JkN1e+wCmmH1Q4Y4tZejWiZqznACBnLV9xMhl+T/vlfUdw/VUFvA/nJNn3xd2pbRIXsO
zDB6BsWm9kXgLYqJL8KGOhVkFQujAyIVKFKcnmYcQQqn6M5ytKHHGAE/gmA/aDztGZCazXaqi02T
+v/647nFN9Apu91q0MBEVe1y9Jeqiyu7x4JohwuMlni7gFH0qulXII4E2DzKugEO2gtldWFGkZp3
UQvpUmeF0NYTc/sg5JIaMstMGLdpDujrzxP+odzi+2KnrNsRAGILkStsbFSV0J/5bd5tl8+0mEeX
MzazNC4fjCV87LvEZB870f8vaQKqYdzf/5uLgh7gKmL1LmxSWrMsj5OnkOwc5XITJmE3Pw8miqbx
dVnhWpOLD+QX+NZBbGnYstK6FuQf1EchAG8wbTQb26JoMe9oQ2weu1LB2fr/CrEBA68qiRor9hLi
qbRdOVNcV6zrO2BvYiPjiu6xeL7vDsWIpzGsoj4AIxHtXBNHzye276zC6Zy53W3Y+Nfki/HjStDu
lTUkq+Iv/PFFGrWIRMXSuZuLtmo/7bvkwmemXqrGY11OyhKWWJiOFgOOIXj77XndZeFXnHDI0KCN
fgiwVEx2Q0Cccdo4teRd8HQPxrypL5WjlmyLo4abZOBiuPqJieX18a5iXYqNEKk6YGlVXcGL+tIe
UAmk12NNMG5eH2SBUOKiFGS+992FOhFUMc2355AxnzliA/WYHKCRxPG8uIsoYRpkuPedqXL5OH3j
KOUEyE3qR//vJ70JqU0ZfR2V3x9gYKLWKzXBF6BJzSOc+/4QrMLIds3QOgYNRn2Z1uCM6AaVsKrV
K5/wq+kLofi9zeNmeKNOdXeBlY0YE+vDVeescrlGWP89zTQfYqLZdWGWyas+HRRfN6i29kP6Yhbg
D2mlLOWfGzceUJeXOLfhf93Nlph86oB9fB+3ZLu+euCTuTpB0BgzlYlXugKd0yfar35HYDj34B9V
2EeVHKLj3vckGkoBVU5hyANMXyB3NlkvfrdkaKIccSuiqcFprteS3aShwV/til5GaUntEYfBDfEg
p/UKupUsXTcw0FRArasqeHd+bbVKMuMAdauOgnxynmSRKkNJj5eictt1M5L6iZ10eI8RKK4ik7z8
2rLqTaqxsY+8RTMwinA4pdyp1972BuoYrYohf0NKwvX+mu7UrMGG3yla4H6zC34CXNnsQbMwXLxP
NU4zRXlEbXGKQp1MqzxlRPUfq+GHvc4GxwDxxjfgwTT0kgfKsV/K0xBdv6iqJ4LpheF5CJC/AGMu
zWsMIZeyOMMSwjbrm+tmmkibR6h9BuAuYUKgK4mAPADJ5ZNW48pr2nVJ8sGx60kFJumB/k7GK8Xk
LbkEjl3GuUf+gKkKGOfl3MmUR9k45Kfyi+XssFlZnpAB8RCMI3sd+zZi4SZuhRdnx147QzOMpiTE
KGvS/eyFkyubu4sOke3IQu9qRjAMnAZ71fn9j3SJq8wtP7ltjOlVL3WgYET7n7QZDZh39nK895Tb
NtltfCvk6brKvNjFH2RmgRILrtY6k2m92STCeMlu7SL8xW73JAgd/ASlEtOR/OEHWtJuVV+7gltN
Gvv91uzQyPoNhg6nDxQ1VsAThxU8/W75tB8n1iOc2RkJjtOV1EP/8XIpSI4IgesOAfkkB6U0OJ6z
6hbqGUk4fwL5bYVO3nHn1uq9EU2czwvGC9aL9XkKno5kI69VLqqfpTAtOayWTBM7uOD0zf/uU7XR
TDWRPgmlH0cddk/pSk0TrY3gQkJBpfOYIUNwr+ZJKleApWwh3GiCzG9Vuh+3PPf1oPpMatFDKH+E
PnqiMyRheOFCNOtCY2t8Pj5J6TRwttvO5N6h5jn/1yBIK9LvWT6T4hq38F+TPYcX9QiwooQgKIRf
pQEo0qrY3srXhDaQh5oE3E6G1IVUyhlTt2uFiZfe5GZ0of6HBh0rIjVFgCoou3GPAGDij4WMWe3Q
c7TMA2lY0V2mfY6a6ediywLe9IRnn2Z556OfCKlNpjGbEU4RB3yxKeQ71Ox9zhNJGJtWSSerS5JT
uJmUlJyg4/AKkr+r8pG3qHLMbRXWegi7DJc1d5wbwtsyxJTxQUrkmOmO1gyNt7Oqx6+dBV4RTMko
TqP4Bqoo30dkj6nJVQj1mXc4aO8TQCPt+Y9iPPfUDhcMg5I0Ydl2xT8p2LXZ/lL8M5HerbAmwWNN
OFLRozLlmNBEZB1HOW2RuaTHWo+wgeob4dhcRVHhp/NzVTmph6bG3PZEAB0l8jLdQiTLcQnrCSpm
QUssufv1CX0LsxGlqT6d11zGSwdgecLku2wnyY8+7gmMQSeHsWsTgcw7pjm4wi4U8P2U5g1tQSFc
LyXobwl8ij+kmbmuFseDugPPhGDOTiCX4jRVNFWC9WU3luRcUFU7kakrRJEqtl1+i0nytdmNNuBp
va9w8QrJlX6pxDak1Ac80cyP8X1Dzs/93lTHuXn/rXGdUTkVdWreUc6vbb68MEUecC1U7otdkjAb
2auxprxuO1io3fiViDutTsisp16UvncT/H1PfiAuXhWS/iHbOJ3GSSACYMeOtvq2YXRDyX40OEWi
648ra9P9WQkkLYbmAKkuxtrggeABOwsSOyG1jJxLYW7czBSEMT+C/3HtzMRGfevCGYjAdAXt8D+B
3tvJhQfLy8X4O/b4z7I80QjeehaliLX2GrNIdUoYgdkb3S6t6sJblzFqo/LbfRCawCpU1B/+eLzb
HvFxY3lbtFRtdzBFFF8hiORjTalbNWUJ3epUTDYlPqHQy16NqyabTCvIY1SIP33YbM6Qu3wlGjnA
XIjiGQou6FaSKiHDc8fxBagKCF/BDeIsb7o5IxFe3dlS8VnJIn71P+I5IjwbZc82uEQlhm8En8V6
FrC4T/a5seJvUuYjJA/wZxqBZaSwgcy2gqFOnS9jsUAH0+gqgD00OLwDAvmImi61GMk7xfEH8ak5
d5QYpvELMf9R4EpdERYzW1KsKCPBMBjJhm7Nzkg++DliRvNzOU5MYD9u5Pw5qyj6pD8jzyouDP0M
RnX0vT9yrYlhLwtN6a6J/SSOoU0vOoFpTEyxZNg5uWAmUPsca1qqYD2HGmoVet2/6eqp/At7Nh+q
k9f3blkZztEbO9pkMq8gC16ZCakGnTDeOusSjV5h45m8ZUcnhGPkg0J9X7zfFK/pXcsBFUGqkSMa
VaAPQedPRZbdmzE1nfg10hixs7N6S8KLAJLr2gB6Glnsl1GibNwQEb5XYzzSJEzi1Fh8d3g4BBRQ
qCIx24OICE1dA4Uyh7FaU6Vb71Ds5pmak0J11aYDJr2ZsEoJtKzjmjPvO1sq/reeyMlAuhB+TgAF
nDGWsqbFcY/rfJ22LY/UCLI6PsJx0Agz+MBVn4ayXBnBAL44roentahgZNXXGCKQkHVPezMz6mHm
snA+4SjzdMpvJNf89ZsiAzXul8aF2aVI/135lXjjlF0V032AgoT6oeo3p2+7/nzHlUQ8tW7mVMmI
MmITh2MMbf67c6ti/FZgIkw4TwzzMUa3waNdCAa2lQ5MFZ8e6ZTBkMPWdGH1DvcQ5PTCQCkca0JL
loNLIu0+tiYB2KCY/1eEamelhj8BmOhNTpTuB+19QN/dRtZ03hD/lIi+GYWfnG2dbyGNZjl2EaFE
b2Mkl5X4moa+xQlQhDzTD5YuYGWEHXZvrpOSz9+OE4vQ1xb9jOR20NHmr4PBcQ8duIMl+TnpH3oB
pQeSAam/hVcnsycg+D7fP4iIt5TIPkXsTX5W4nbwfOzgwJVmCsvjfOSOT/NbIK6YQmcg/y1L4u7S
mPXUjTZdxDa98wLJyqgGjSzLdU4DW84aqndnRZyxC7ZvDVyQHGY0VQuIx+lFDJMOxPtCjTfmYpH+
DlvXgY158UJdipSyu5m6A7DvcN6UGwgOw0vwTUS4+6AQCO58N4+U6vcPB0V0RuzRK0BYeOq5mKJS
Lbiv3ht2kieIEDWe2Lfmeyr+2sB8Uehh1wP7MHEYhHghwp/PJUw2I+DgjJsIDlVxCoA+bngvWJTy
JzxXPxVWlt7YfVuSnM9Szg+lICu3mkgrpDvgaaXFDloBUNDTz5F8kWpZqXXW5I7AbWYEwuM0HJju
jw3hm3EwYdCAfeENt5iw5nDf64uH0Fjm2Y1YUsWfHt9VB9WgexDPXu0ygyfEU39TbfYdcGigSyG9
86Q5plJgSgGhTtHpkwyMzMnM5AHOyAtEfy7OEeeh1JFvL5aB/qA9QxNGY64NN3x8kMbnvaut0hIC
eMsDT5ZHVKAcLJtBy/coIaqinFGd52SlTkrxHRcDc/Sg1jqWqao6wDKivrvcPppaXSD3ZzKKIWfY
e7SXzO4DaInI3w9wi7CwT7Vfct3uCC1+NgRZlMCPSB9TYGy5e6HegMqPKeqi71mcIN5SBO6hQt9V
iAgSj2zubFc9GEFU17zeK0tXEmv516VWSQ+DCnjbRcsZxmf2KNtBp1uwn80K1VJkg+/d3hooVZ6l
2NehT2QBdv+NkF2FFq2NVX/VRhAlPhAhD6EKISv5/XCjyQlBS2quU1/VqvPFIMrj11vpHUs/TAPe
ACLgphpx9K2iru9oKXp6AT8M8tNqNvsTLFXupKMAUa5d2gZ+MfLxRWH3bTA9nho3xf9bU1m/5I9G
k1NypubOh2aNoy10cWRqSvKjH30A+kwBOJLkH7Px+WSN7iIUOTjHuXTYeVrNXpdkbCktdRD7U5f4
2VTvUdtoLOEDLj83dpgkEbT8gprfKk9DCVUlpjWEbsG6t8fz+KTgixLIlVi6XjfBskv25qKUqrCO
vibH48ZeLvPN0Qsva0BJgJW2w69b8NZrT5tvSJsfLpP/nQtOed4VG4GkeYF5QQ7H1/Zx7NRqlRBe
5jNPkQEQmrxKzOKl7nFrDxTiWQe5GOfJ/brwbNw8qRtlH/V4sDBpBGpxr/3kFfSZ1V4yf3p+IZgX
4J8XkSn/cwRi9LtQlSYawIcbE+xYrI9XzUZhXPo1bHEQTBskHpEkhH8PAR/N6Xzifay8mwWYNivA
XTCYW2kzu+ajqACNR5JB/gfmr+wodS88ms/aoszPuRZivn3/CIomqvISEPQbarf8wBluZNnfF1q8
uNAIQ9BcowGIOtKUwHP+UIXtF0/a+JZO/5GTB3K1akzYRiydGXieRBr2uycnHPAogKHuXrqILO9U
+tM+QaPt5uimgqkKaP0WyBpPdQ/6/AZiUqEUqhdb8rsAms1PLzK5GAujGOw1pnPuL8AWUsg2tfgO
LHkERCgp+pgrftkDKBWWv3BLcAwmqT2eQXFmPNpMWuZ1cisfACOz56Ls/KqeLFRyX7/F/0KXmoFp
Uj6/O7aiW4+WzUgtN8b9F2TtMX1cVpvoZsVILImXnrzMw2s7RmyMqa2ryEvq10iGVDf8inU5Rsjz
ywX5VJLEiNB8QwAyhBzmh6W2O0TZE10QvCfjopLuSbhIPfXa3kuc3abmPFoTNPhAUkio0kmKpF7+
nVcYLxmBZnZy98RoUXA4hNdoyx0/qeg1k9vOSnssp3pW8cvqubKfnEOJNeTA0SJpAJdksn93aXy7
bqFCoOFQ1OsIV0IiDFP8eeo9/01QVwoFFICCxht+qGEypPDRWViXWI+RFIMIPWsipDUxfxTzwwlA
VkRobqE7yDTB0tNyF3FOwF6igYmlWWlnhBn3DXV12xd+FSLPCwkUH/W1Q1tpa0wTEt3vELcGLL0y
cWd7JjnIiJOcbXT4rtaYpxAY2ripejwOEzuKtSA1vPzxPR2jMmlSR2fkmyakEBlucQXZQZR5EeHB
65TaR0B+Jl/WhCIvhJkoNfI21AUPycyAi1kB5Yo7dBzHcv7GUoPKnbjIhH7Xo9ls16i1mXkmixDt
i+P34txv8Qi3PLnz2FvvkPe1qU7naxcvKYfSVN/Vi83SLaqKFisub312IBuYWLsM9s7KMORuVyfK
w4hWIvW4zEVU14XMjp9SQ2jSj0cLOdwIJOMriLcvE3WO5oeMtJW2JuHu55w1jwctKUlR2fLjAk8r
OjNHa/xHJSKwhbx5XYAmG47a7lcEWmvn6ay4+OdiRzMd3jc+sxYkx6EzPVJUn7BWT/KfrF+5qxHt
63sPz3r99a9VWnlA2H81f/tXknDYBkzWBcQPuQw9IGHFlFzIRyCtiWJcQMS2HQQXi7zV1f+WKgto
nELCOx/ZjTYGqhsXjkAqJBbSd6iixXCbeMklkOejopBCzUJfAS/PHh/DIwaqwyS6qqfrj6+b01aS
zBxHpS9CFXkcZLVQGHL52/RAnkSjOgNoZADEiS9/m8TyAE0PWNJlVwnSxV/NzyMB2tL4A5dMaFYH
4ZcU0l2fEPHwwD5tdLqqa0HSaHsKnLIxOBu0bLhMQdXlvbj6Xe/bMjb5SexST5DQlBOygsMn5A5q
ohN/sko8/X/WXqLbqSdwM9BMd6lu6ONyNDMQ/FFiClGgA6AwfPGpraNz2dFvjoT8II27GgtWbRLE
dkKIt90K96DbEYFmyYXNABbSm5OWMXZGZyySeDUkmvu7kAX26MUKbHhgnQL6EQm2lzYVWIuxbK2M
6+z1HJrN5I6oYY+Sgw07QngfcWR+3xCEOjoHTEUKihhgOI+IxWu8TOAV5A9WlSx7RugVi9zzMI4D
9dtKd60nGTqWN/JytMJZ0nQQhafwSR7l6ajPWLseBiPH+rZGJYPnkkPC2Lnwn68AbJLLdaDLItmL
F6tyQ2rMxkavAfZVv/kCb+ocCKFormWWE11+Fl0vowaMnBMlvTiGg0GL1lS3PIO56fxVaYjIdgtH
GMGgUUBYG4aXHbFVMA5x/LYitIggkQuocZmYDnFp/bjCKsE4Un4JRWdkSKpmUa3YKC9JgsEvZEGH
rLP4L4ZKNjo0plK3gQ0HOTqzOmrgFzznEgJhXvqE5b8dujRibGOQSwtAZuHFpuOERG/vIYs30XyN
xcjBzh5xF5RgFazW8HIBEnY/V0jN55Ofiy1xbjVk113c7tnKcIe0P+NS6lqcIjpwapFY8B3saPqQ
IKEZRsN0Uu4Wa0fBz5wmd8Q0K12aZTVxaOdY5OMSxjkO3/kAj2GVi7NQDN3hqs3GjtCYeYOy9eaR
D4W/f14TWw2tXBcdhHUhVzL7dQCvq0LIv7d6hD8/IGa/d7D5G0hu60p+XlXkblX7W/rdgY5dyXFn
rFX04b77CxeKc9XgPZ5PMWvGLX4u+AejDO2lqBR68dpuVRRHBRoZzHxVFZredtiPOUcwg8bBilcC
P+UXW2Hs7M3VBTfLI5+umJGxjrXwS3WDwsfRQRGhvHa6DVhVg2Dbv3gaD3GZeQO0Ypv+kur/7m2z
cAaJIeop73gnDPsRJMQZpaWrkVtaJNC9RA0rP5TxT0MyPZ4o00aY0Y/I844T4uDEtXdcp+4dNRPa
CoxgRZ+QECUSy7X4fIikDrfETFotylJbW7L+3qChj/AzgYG6af3Mwt2moAvh7nmbC7Zoah270D8X
XxiWGes79pGOtaz6B67F8YAOS8DK8UG1nnj+uJbKq+je0/ITqJRt+UCS0r392fJFQMuNo1K+LG3k
PpVdoH01xBIWpFT/OTfvft0yDa3qu+jTMnXSM9LEvOsebJNrJ+dRpvBHtCCcE9i7DDHgRXPZlMIR
BKUfyRaff0fEgjQBzNTyq2xnx0nTmR1EX6v5yL10Al6F7fHWQdB+pVnkA9g6UgH9q/0/arA6SgID
n8DvOySNGT6BC7TFfMXR0NvmXzybWmxBL6L94NyIP/IN82P+PatQEK/86+RS42J1y+/PdGSAhpwi
m/0l4dMOxw4WEbTDXWYoET0UxJqNxKIOs/YP3t76bLOzlIJbeQPrsqnYVahKOyFm9UHqz0Z8+6Ry
rOZiNMRTCptdzmpXktMjZE9tUxoVEInCkmzPYsHSxgtL1G44tsl342/fGKwqM41MRPFeR8lp5EKn
fUHsoF3E1Iat83toTSq8l049mTjEtg91ajFsw3LFnp9UrrBbcetEx37e9V8asyVrbHYmDKsU7A/m
UOnGSQOIvehRK1ccJAc02oBOWXoDXXCqT9Wptdcs78bVU4wG0QVWfx3uCD21TgPjgeGTqImhvNiu
59UUSdurK074+kDULDP9dOr0wlzMy+3LLC/C2wGk3Z9GfAiiPFnjT1xNKewpzG5Bx+YxwaVhoH1U
+DzFCD/ChpwUh0RYiud0qgXYgafZbgwcan4fi7X+lukwgkT/dSN9Fzt9mPFoVK8JrplblzGjS4IQ
A18iWJQpRHSlvYiTOiWx2aEWXhEreGbFmeLCtoEz2WdtL/miWgLtS5k243svKiljhJ+Cdn6kAHrq
l/2EUuW/eNmkvYSiivWUt0b96W23kw9kLjlCxGcMuq9WFdCao/1sO7W7wm9EzmIaWLR6sEaExtnF
V6ZE9PsmsaGwAyQPfO/qf6gum4XF6PYJmVzrtkRjVQd2O03rj236O8RakHt+3EUfLtVa6hfN7imr
22+4kI3AQ+Ozs/8o5L3nrndT3gaXlFfFjSFHx4WIWHZM6jnwrD5C
`protect end_protected

