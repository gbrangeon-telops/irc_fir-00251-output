

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SYUpj6do5sFTflpbsRmqzQKFPQDYrJyRQArefGItBrRpeTStPf4iOexrlL2KuY5Tjxr42gzfz2no
s00d/SuK7w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NR3ykkYMNFMRKu0xHAyt5DYiOktc2YTf1JOlIURJ/ThqHJccRXVvH+Sc3vg9x993epLj5za38fd9
R5dBjv9keX+G5g1u3CtBsdqXK+hNOz/uDIy23yxr7rHw0ImE57TmiDkVMvMwv3eYKhw+6jZKYes/
orVUKkqCIC9qrUn5RTg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HlVxjhtCNCKKX+WIZOv4bglrDneJvrVwpTadJxqH8bLj9DfFux8A76EOB2zOay/g3B51jEHFXs1k
cSPeVifBOPOW+4hnoJ3TimbzQC2WXDZLrgI3HV0zvi2+v+260AsNylQU2ks3dLwbxExBHvawkhdm
qLdLQIFdyzjRMD/G+fo3ZOpvx7tOdM4iBWXd2qur6t8wJth9ryhPu98XGfaQXlmJP7Tzn+0ub08s
DCWHug4G341eF+dWmcugGtWe2Ca08XjibeU1gRioez7LDJacBlMb+me+eJNl34Hg9trbjeo+4u2p
UhjBKGy0TbAWhSuuGKcCtfIFOUbYcwT6t2Yt0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DoI+R7m0zbJxCq9A8c+QbVnIsy2kNMG29/strbjpu4rQhHX3C2LKQKMwC4UXbs35yFBTN82oCtQE
LCzB557xK8srP2DUb2FdCBqlo4nmLOUDlZKHLRnMjMktj2MJoV0ExtbMFAErwe3zZqIBchZgf5Be
0C+OuuK2xw443onEGyA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jkJi3dDxF04M0w5noeJKvbYmN6cGn5suzWOH55jYT8k6r3UxrWZdHPmAWJgyGzXTFa2rcCzw1zFN
8CUT3mqhUaMicnmv3k1IZXtmQp8LLIMHIhFQWUBUexg49lQQHlMizPzJBAEcyMQJQl2JrQBPC4y3
FtPjOGWfsQSXXVoSz8O8MOKUSTmbuzqKeAR7KYOBiW1PqJBZo+vP/teWIw2p1h9/ADBVH7fQiL3s
cyUleDPcPx934u+grxqX5IGh+uK/gO42i4Ms1tDDhMblp6piYQ998xcC3XiMWw8hwmR+KGnfqU8Q
VD22eRbZMxNB+D8sxEO3PnV48eApa0h9wT+rpw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30848)
`protect data_block
uWLXK37lxjwj6aE+437MNxFPrhdc+0z9g5RsmhhjDTBm0bPl/ORQmkAau34LZPqMjGglVXARjNfL
HAwmHm5BJdW79hEEuLwzO+yuWwtwcDpsqh9aci6l+hvw7+Aat0nBzksYa1/2KnnPSw/9ZaMK7+dj
zroG6G3Sp/u3Ojdrf3sBYqVFLtx3J5pHLk/fXCzc00LI7pl1kcCYGirx/VeOuMIr9PPj36JEzbLA
rZpgVtUJJxOHfMTwqHuIm+ur2zwLReNGVjJT6XLweKvVELNniFlw/mMOxFOU6QbARzSvQW6YzWnx
l4EZjhyxRzDk9LuWVXTjZmZ9OkgH3KKZDbxyN/VsQ3UviT7xe2o/AIsBzy+M4fvPIYITxWC4++UX
/d3RXD2F9kL7sd58ss1wDU5VZbcWZT0Fouxy0/JKISV/opTICiqAFv3mOw5s+kiMZFktqKwefwc4
wCSnP0LKHL3/BardXyfJmeVjKgFa+WCKPwnpwkErSPADpUIFR3J3BizqYbBXkDmED0/PALrpIhHf
ixzyeluIaJ7pb34Pw2Z5ECv3eq3uPw73egBeJpwtH2yrug5vvqOQVa6gZs9OSYhykG4+p38b22hz
B+Eni02wD3JbWVrqAdIQmvflKBszm+AhD6BAPCiJUjhL+qrU7Z9OihwE6UFleU0kk/9j7hUCHSxS
vo2PYTOvbwHlkqkKGVusRS5JFLD5K4oSK3eJdL16rRb+R3GxFxzYte7ISa1PqAyucYpTDXulcXez
88Cpf/iSER9jeu0k9RZn8mrO4glpHVXTPSfRP4NToQ5l82ynPJJ0Lq33UZWHcgKIsl4YVHhdTEl3
DzsR4cCrzOYGYsB/bu1/aG8ENdcmPSdSdesNuZcSN0GZAGMP5sV8/llsIODwG6r/tRWvIX2N3LH3
WlNtbZ6Af6sDD39ELijqwWkxjrNfSbU0w7FAMHl8dtJgrM1vV+ojEY8Gag8RxEY3AfRUh2N5m0O9
12kwyeWzH32sArnEJ0jjaI9ddM7piqhJH/gbCI7Thod079xZUxug6IUOVQx2iGBY0gaqtFbMIHwf
WJ2ruav9Hr2Vn8HRMHdyFwZg+RQG0XJvKW9NlpFdEraAPAOOu73wcMw4ZZtP+1Bqf2ZF2xoO8V0S
UluDyTzvA06Wt9kF25octusOUBbiatZnARC7I7DUK8Paq3XZwRsqMjg2u2/wKZ0wrz8+iMWGGoId
xqZF0ETOVqPZ9noSCu2Yq85AHCGpGI83e6+vhasT4b+69CJUhZSrHo6vHI3hNxHFDokUPJ3Bk9DE
pq5sybnBiw4gtOklmtjYxBt925Tc/tSNM6f2yJKS1j4WTu6KVRZW/jjWtQsEO8jgsnWA9ktbEEHe
CQJ6YxrlrOuBNg/ABP90+Q7e2yZ4DRSxRLiEWVTFLN/Up8kyqYW4Xlps5aVGqJ+XPk/Cqotjot4f
5xAt0nbhDF5Fq4PzCtwSXKaCuTCGQuIRsiLa+PYSkIqd45knyNfdFmeygg6KXysegdtrbBD4ZbTC
4EizA1V/kRNSf0yKAZTyI3hVjDF5HTQ3twtzCsEzVdQiHZEOs7+5tfnV48whV04vylvkPu0osM0P
EBKcft+fM4Xh8IXmDKkmsc9bowosIazKbgDUc6R5gmkzcnFt9x6qzuUWhqNcbODLF9RZOgdRz8l1
YHvcZcJc7wzYx5ykcRk58XD75DKurbba8hawRQwsvnvX9msh+JNWmMK/6XPmfPrlCbMDjAX2t+Fb
RO2SkJwTmdKZoBL6V23rOml7WOoPuliTvX6ktPvohSM1HbwEHWWfheW200AHywu8A1Mt6+W06heR
/HsCqLxy8eRZ9LBAV17c/4O4E9Ouj79+mlG4OtYUqQJTx3K4xm0ffYnXoLu1Z2oprgsfijUummA8
fOOQHVu6DikbmLYyO6vKv+25CnKUnAqLiUpv047nVY9vfJV9bQUq1sPd4vasuBV+5F/sFGDi/iwC
Gln9sjqSjlz3R2OSqMCv56KAJTNcnk0omjfTm/aOil+i2PnjiSnrN6foMMR6pF5estS9mAELuQgC
rFb7slGA10B/fguzL+//6yhBOHhn+1mn/hLC0hPFGAiOEIHErndeefYhLKYfpilFLKvYBU0MI5H7
7VS8PZSIXI1x4ZYqtYK4QmAZHIQU+q+KKv5xYdIw2qVjYC5NMEdb0olNo6gzJ3bmTaZQyZCXLVm8
VuwcGRsmCWa1l3IkAOjbsdmLrJfPhxeFb3OvwUK4fvfgX+RBBJtbibhtKEuQwSb5ZRUtwd7L5Sr4
w4orDihScsw4MGEw9alZC2L6eNwTPOiC4iYTHU8P/ZzkXnNDWgax9xxITXtL3D+xMq6TDwybGggD
Rvr4IGjbFfe6dW5FXv0Q0ePmmrD+Qs8InCimV0Tq8lBx54O5PPQfo3BgS/4jRBBnK+rDDRMUrHrG
6Lg/E+UJq9dLRGq40fXRXy7t4WBNjB7qdIRzkqtqCZpNTxwsiY5ROQmn+c04GCOgMZbaCQprXlnN
c4Vx3hTjFG8gb1DNbxMoMEgyAHW70p3KoMX7qaS27SZwB6/a6k5B2so0MWN5xV56TLP8PTk6fFs5
4slT3adDKeAgSgMGlUC0gy9cX82pUnHjbCjxlqtVWpbqFGLkZV5RephaU8wsaSCLZhvfGfCmPDtS
MOtcFg3AL1ADuV2PVTVkNUavC2YuMth/gDxCAkP9M7yhu2u/JMFhYge4Nz/Qu4oWFu3NhGcI/lLU
DtSKmpQlszgSSqGqjlN5SMsbiXjouXE/OgVFUZ5cIM1UorV4owXy/3i0nQxOlU/WTBjIEwy67ToZ
xpn5zyGbE92O9y0tg4HR/Y6jAnRpWSH4zfVsXUw7Kc7MpVX3ri2WAjrsNk0P4E7VsHmURMZVW+NA
p45d3pTwmEZJ+JuJSf3JAKcNBpHab+QZf/aWQ2OFwhyqcZ8n5rzdtNHrdGNnbOTaTkajZ47Cz7SF
BI/OtyK6uJd9VsWpXLYiA77SG8sxRkFaYUVbC5C++ztf/7FC+SXV9FSmmZWkVwUzAzejYsa0Yqbu
VAXeuP5rKKJ+mgDWpYqlrUtr4e7Q2V15uuCMZ7R0ML1nD2lFXAKAvX8PnvCouw+UZUF1n/91v9Q4
FFQ1splVA1aubo5RfoJu4Z0h3QgJxwiTD6F61dluCNadEPm5JOEVA7j/+oG5eK6ckZ66fbekr6t1
Yw5zuS0qzaP+Dx6WhDSrkTJ3K1uOgD38JnKtf+KVwEXjDiqNO4v5En6ujo1z4/qliEN2GVCYApn8
oPnNlXljNihG21AA1ZTXJA+ZKqAk+nF16G56twDnXIwhtIgNNRg8Be8FYoWXNhgjkdKZ5r5dDir9
GcRgfbm2pAhuGqNBgvCxvaqqZHiV4rZr3rxDI3zQFbKPk1l7d+L8pkSlF09Y6JXBshPcQ1iNuRMS
4U+vfS04R7mwpsfUPC/3yHIUjmGw5lYA04IvERC8NK6za+MGGDzY/4BfuRTxberkQfUwlNE/KD7o
zbUArJh5eaIKxhBM4/o3FJt7soMjcmyCiOtNAeybwy9na5CqCof6xh6Ax9VSbRV1lVakZFHRUuC0
aQo93nP/Q4jfPr+6AbiZUE9f0l+FK8iPfRZy8v4Mx1kii8luYq7eu4aC16DL4ZWszdBlz1QuDeTX
NHIfUA7cbImzWOypJovmo50Yl97JmzIH2iobEXESb4YTvxNMb/yz2PtpWsuWysQN9SioM1qngzmu
Ja6dEsoHCzhMFKa3oHXnjUOMbnqGWZo2URY7A+4k+uRD2u9RmxH/mJByPSK9uxRGMtnjYoDZ84d3
ncPIOhrDbSqg9zV48O+M8DHunxYvCmfRv0jZJiWbso9/oMf7VTzU2NvPh2YHd9m0P8R9KcNw7LSz
KEuWkWi0PPKp0o5hFvrcLjS4LRMdqgm8YxjMfP/fuKU8LoAhGLex15cve/DE/CFplNs0C/krvkQG
G4PbTgivNDBwCs/c6ggnKXlRn4Q131WAYkQKAA6S/Nxzo7AZ+3gCBRsd/c7hHJesObPeO6VQFEwt
94BZ9oRS89J8fMt3GuoPgqklyt4YQ2jztYtSQSFfv5kelttBTsb+odNdKw1TaykN7u1V3ufll+d2
KWSVTYdMIIuvO+Ob9asA/pUzxlrphxZku7uKkaP49YrervvrYT5EvO/w9BFJyLo5ahSdYEpMDJdm
L0HkyCfbOdo9MX3U+Dvw2UHABFbrUs98UpkvO6i76qioxxFrH+rPxVDLbeEpLWAkw2vnSflwiCRe
fjLXoNwNpsNa1JOsTauM78f1+TiK7c9jK6xaCnhKENYDTsQfsOgsxA+x/n3zubMrVRBUBW252kfk
RUcmBeTyvty7iZ/d4qaL9jpvqDHHxZU8xIQJwFPmm6Jo5jlNGXfis6p9ql8zo55T8aHyYWPpW+nm
Wg0Zn6PFzw7OnRRoTXWRXs0srhhGEOTYEWIn4xbPiCgswj4NNxjic4CD3TBtdDyu7rG7/TGSt47u
8p2PmAQv3gOUPQhJ6JW4yQUWXmX2//S5xLWGoknn/z28Bp+j7NgNk7isFfwGbramwodxjTv3yZs2
KLBFO/Yu1wemo9Q9j2gme9FoaNqe2wkBTXfWlGRZg04CLDeaP6T57oXpgPYn2sA2pKGUGgc185Hf
ma+u7EB7kODrkU0c1FCzldkEA1DxEMlDkWtEdUS6r1EhMmWdlK+SYK+5+8Kcs+uleWU/BIJugjyj
7fSKU8kXzn0o7rh8r2Pr9/p0ODVTiOAQj6vmtASzqahnIlCBVpwvzuQl3uiYUpniAugnReTJ14JR
kWEnZ4y8365x4oIxakeyeqSWDNEyFRi42/bxptDnN5a9NDuHTdn69OcfjdG5Tam9W0ytzgM/40m0
9a2bf2kNFYsrHzcAuN8ooctu/10D9w3WyzcvhgfpvR2nTzf8OAZ5GdB/nZhK4u79nRLkbQ7IavHF
PTG6OyPXYYFsbYRPJ2zjUS4q1SQOwO8A36Z91XQWjBDPwCoW2RUSfds6k9Y/22WRmtVoKZpY4Ado
N7oKUkm3Ga42bWk6MABQGLVApCL1Gff1/86zECnIg9PBjsWn89t0EdLOZ1F/aQDHXQ486cnoxmTR
3f6JsKHUnq30eg0C+x4CG4H1bXaAULliM6A9mVtSOhO/LtEvHbOEdiGu2e8AuZizQik4R9vXrUvY
6bBHWZOdtIo5Wz/fPMh9+vi3Yd5GbkVsMDGU9yIMz+MCQoVrR0/IX+la0uN7W5bPuwdCpVnotcH2
E+Z40ujY5fq6I1l8nTHo7W/Q+MJJtJl0URga0KdJ6nTy1Ux0RPpvyEKxkxmI/5OHgqyZ6juhBHfe
KraYyMqZ0Dvcn9SLS3iFlnbmnR3GxoKz4JAo+k8FiD9UWj0+hcpg0TdGEgvXNc2qELxf7wj3D75m
/2V3foV2deKrRVuX56JhBnoLTnlzXR5qSKX8BiXCAPmmecdmsANhCi5EApjNWwJT2NRKlZNt40q4
+8dNmr3P9xz4cnoyq6awwkawnFSMb6D4vPreWR2zfWiaccB8RsB9MFaKTgRJNDHJLK5pNyAatePF
5jDZGGatRJWkTfFHF33OPhHvKRNCeywM7oegiPomeplvj9QtkeTWjn4LdRgHoOcyhoLYPP49s7ve
SJtWaa5DzjlX1h+PvfC8nbZWWIKLEB+3lkSI1aJVF+FTPJySfv6dAECnAyax5hO9gEbLEXkHJr2s
2s5iLP3sap89PMpt8B7Vt8aeTip4mRzHMVfIvsdkZT+lN7X3LQtLVbTlHL5nmRkvzKYtBfHDW3hA
+oACk7rz+VNqDkY3wCP6XIE0CPwNS7c8CxGg2kFsqQNc/+Ihs+VM5Cnh1IVJ66sECE/CR+5ccxMH
jUtWzOvQLR3rvb6m3HZg55uEYdb1bv4KznrVaOCWwpPYSIITcVfLsEMilkmZ0zm/jmCzIkSCsQgY
iIEe3aPiN1JbJHmrwTceQuT1iYPKs1mnNE5DI1LRzlyd6j3AtdmsLNqdTUMF4XmmQiT7EVIioCXu
QAIbG8voCDhNgknnQaBlINsUWVm60Tk5hb70QQ0MQoSk/0hnu/sfseg1ozASRpHzrDjnECsv90Eh
T3cWzerb2szTFDK3txukWILOjE9qbYQpfBJafhBN2M10DhaqW8e03bapYM76VP5Epnbvr3oGB1u7
PXHud3bcvKqzCqzMDs9TQs4VQ9wn8T2yMFaKMi4isAQ5yKMSyE6inj2owQ2mx+PgyO/x8WbLLPCf
GiBmJ5hirIMV2SEosS6BD6cm0E4g39frCnbNsuJfQEfSctDvk2dl5WzNMAswOC225/93kbBOS1El
J3/CQ8bZFtMYx6EwCttxMEg3s+51+qmMdvclTerR44Wlh+bvLfun79fSj7ufj+0DYshzE19vNLS6
oYKO9B8oCsznXIyIFf0raCop6/p+xPbRH9UQxVJ0rjWEtYqVDqS7rrDbC559JQ44YkfSJ2IsRves
jtpJFJmaS7AlUYUNIwI8C9keaU0sVeUUN55qUBV5TsbnJ84ywKdUGeniWp2P/gezYUccbUrz/aie
1X3ydjasxOjSE8nEqUOHMnxeMAG+f3KYD3/2Qq1bLYtA2+u9VOT7uYH/lkcbdY/FUnIZtXyE+cSt
C8ntASJIwMYOo/LL0Hmn97jKo+HEc7hkVs1owS30coLfCvADRH8iP9s8a89dsidWWvw7GP4jRIln
qqA7sQ12x+8KauqwOn9qPmtnSC/MsXBfj7vCEL2/cRV81pQ5Ive/K76dfjAZbBZO6rLLmTNPJLPS
f5QWZaqSe77ndv/HzRpyw+rfxPu/jpMiIJI+OJDtAoUxDgA4bxBoKY+EeC75efaS97Yx3X0ewjyl
HQyzUWrpYYmBQc60dbpkhz69Wz3QS/2W5HhyeSsdG4+V+kn0JEMZd6eUXqwiCZDEWkPv8p9WfmR5
QM9j/lMcAslYIIG6kH7gwo9n+Ba8MfoCFUkhYfJw/W/nemJsTBc/GCIc9mEaPCLOGHQXNWvhBZ9O
eOSDIljYNpACldO0luPkBuzZxhRlHhFnOPsnsg2dTBBhhZ+DEC7l3aIMWzepE/maPmF47volE1ln
ZsdQU7kFlsmHui4CgfBW3rLPUnTpyoFKDMP7RWRYC8F2q6hjn/O6dV8Rw2cbNJGdxPJ20KPlPR/s
Pul8Z2HSKLdPamF1ka7nRbZTLHP8u0tTpBWThtg7UEywjQP+tHuWE+lCtQWGAD/cJ/yEVqL/401X
KxLrWlFBlEUe3fc9kqG9f9pjIVGiwxyDAqKK9aSXZDML/vBy6OdLgjY+movXKL71JQyAXqiv0tL5
iZsAvj2F/SqLRE6dA058uwBTqclvx7y37UZotqDRiT717resFOMTK0ki+OQ0MOgS+q9t9MbbUKQL
HHjOa7FOSeX3kYhVTpG6bSILOHwjGCNR/K5VtGV31sQphdDTQDFkx8uDOgoN6AESuSa4fsJnLIFK
u1wBjsdDfs6J9nyFVf5OwYbN1SIQ9k4WL2YS2NDqMIW0pnXrjfhsTvBq9q1lxWO3Ai6TEe+dzjkp
ebyPq4hyMwZAoWd+/eztwKfEuV+P5WFSNw0v2d7gHbaVLdG3/1z19DivS/45VEGoyHepLO+j9H3U
9oarSqajsdTCdEkVGIDx2yitBVv0m2DFkLHJPc8pU8BThCLmH6h8PwPKCNXvhP3amhO9byWDOQBl
31G1Wp+0HW8bqONfdB6vK3zOJ2zDBZVjhNCJZ9RAV/bmGWW7Np1BaWmjVUooePLrHyJaX9NbUFBj
51PBFWErgkhrpU2e3drEh8S38D1Aoewf0YyFL0oxL9vesNVt2m0f2m1yKyirWDm8QUoxUH/rmWvv
TWw52fan2uWSBh5f3UdIgk0pWzNITU25LoXhmjuUAbM21O3Z6o7m05b8EXziPBF8NS3U6L1WoalB
fHz/kJUu1qoe2MOcwn0zW/XjIS2C9mQkgEKOS9dMu/3feVrmUDqKialJJqszoGVLckh+71zcGaVr
CZ5wW3vZzNQXC06HHc4NiB1k0bO8rxmWovatni6wU9oC3qR4mRqlSflTI/gyaU/svV0VCYKRfucL
/qLdeC5h/3dRsBq7EDLtj5luFrtQZNrn+ZCkryqsIcqZsK9syuupNDe02rcyQysKCDOe/4ERHUS5
14JHvUK5rPOyBGeNY45B96d3GvPT4HP1tQ1QO3qdmmqouCMmlLC5oPEPV9uPwvlgpPcsk6cPQB8p
OnrfD5Ci6oxYxz0D12TiiDVzIjiVOaFIYYV7e/cENfsFXrxy+Z0uDR1ZwL+kIimtp29J1rlwNFj4
Q6RpB1k78/L1aqQYfBhsdVyG7/ak09faFlZNAaxqIoCo5MlLnxtzvpUgOzn6qzkI4jdbTcfEA54g
VrPjtoDXxSWpQYbSXGwgh76HdQOzkD35890m4BbcCIk+QiSn4ecERJTIu7Lvlo6FhNDDPdjfMUp6
NNr/j/IMXzb412FQhLj6Q7UoG2ZsTjErh8sZRor62dcLM+hkVaOdTKqfpJa/s5tnuvpj79uzhIUL
2aO2+DBWp7nh1lpI9Ojq139mTgtk5a9L8shBRJK4Y6nq6dHJkVJHBrK8UL3DPaSwGYH+hef5Adw3
WJ2FiheFz/hjRY+rAZKTk2si3ZTeXrrKOnSDnNW8qGkTab+8W8WJDnnWdbJ7VEhoZBmObtDfc3p6
eQfjdZWXrLY3LdnCtc4loG5U8Jz9DAOpwg7zKlkgU/jyWpbi/UtT+PTM2ofVnH7z8fx3rGGBORu7
q8f0vf2whQ7KEJOFNyCJTRszP0omPl2HdGxO1oFZjta8DgVUQX0HdPLG6PA5Tftbk0ZCMCHTrE1U
oxmxcr9FonSvfHVeJR5RdOQ5p8mU6iCqv+MVsDL8jr3PfsRGUJOveUJe9J5r3YKomkH0fUVAweJh
Id/HNaOgQtCpRcZyR+hQClLfrFGZ5qU7GhLKFH4uBN9Myr/z8HnGaTBpsSjCCXSnBMYpt1hBfpaG
BAYuU8iPR4l1flaBSiS7B0kqHACaCc5TVVZhtFSMq+P/b2WC4CS/SNVcJGkELq0G/Q2K+XK+xQsi
PUiESdHeJFgg5MG4QTEH1TE/vycLl47cjgQpmxdU+7VF8oMlOplS6OtweCd0ldj9LXfoRATRlIwo
iz905nBf437iOGVjuSevNsIJ/kJTwtDVw4UYDZdWaai7Dfi2KNHdhCLXSu7fGBk6Cj1BmfE1SrEn
BnMBsfe3FecWzI0p6g3b7PsYAyKnmYTKarycbkMcOoiMGJYrDH/dtPpgCHiAUXipX7+C7IqkRP1+
ObPBf2uqn0g8Nl9lzBEgdayI83jd3wHDaxfvMtBpLpCerK5WvY/RXRQJHamvZwgBneMcQsvKXV7u
dsHqgWbkHq9X/Urq768LM8eSttRLkcpaSeYPns3MfeJQchX0u5gn3PbFA4897xrtJkgWNvPC4Z21
pUbISimJ/poT9kTZTckpJ4dXx7pJ36UMv+mSvq0311TuYwiptl2nCIscfqJSRIkJmPfpCbEG+0hr
lLXhKDkLjtaTQzrWkuloMbjdP/+10kxG51tWk8bo4Wu1mKfDXNKOrYYH9AcsyxYEnqxReU9ZCn5y
8GMz3rK/4jonZ28DOlo8RxLHwJp9ha/3xXC2idsHVnvPpuk3rmhjFVMgp7FdJ38ohcHeYVArXhgw
glrKEovSb9z/oBDz0GdU5lYOKoAixQEQnxo7cEkQdg7X142jZX3xH0aOakpThNCrd6OtEic+yeIy
ciEhu9qmmWOP4VcbathZUxZk1Ibz3Sy5LRjVSZg5+1XMmYxtBTDX4w1DaFigJwIJ9V8yHUwjjDhk
bcBvPfNY7QeMShecr9xijUkvhjEvanK+K7AprHX2JylPubWT1Z1MlJvLV/m407w2MPZqZoXJerTp
H9uGHsYAy5t9DzxPEZIRp+hf+38CMhCDQbKmxWWKrKaEoibOpIoJlW6g2cMTs+aM5fhEBe8xG0IC
X20wp0mK3+ElOqodLYlD+Qq9z3QmBdP3Edh4w4gP2QFTL+CQ1SGExW3gnKxjw9AaR3R/MVmRdun8
NLPwVCKacPJYvZ2x/8VuXMeNuBRggsWD1Ax4M+uCYgcaK9HjkW+bEceklKrvaZpWsqhfiA1kApmh
tk4/xx5Il1SgwzO5evWQbJ1O6Ifx3rf5aN17ty+bvB+qC/CC+4WDgzAllY3z36cyc69bGVnAVwzx
6wVFYa4GC9Zt1WrxUdMOyrNhxs+EuVPOsi7zmsHTwVCPye7AidUgqE9yzHtQbVA+0PPhoSjwGZC4
i1Nksh6CR9UtlCgUj9Fo3RSMg8iaW8FG6QSEfb639BgLZ9XikeFsNhHyA7Cw6+Zogr2qboO16XY8
InzATn7FDswL1EdpyrmzOC90KL245ImsfO4H88B4xaNrxmwUSqNQwr9DK4awHKdcOElIWaP+usOp
cuPgQiIxyGJXA/PX67uOpbm1924wGTHv5z0i1CR79Zs8a/E1r35PHRIBuYIeSGt7ZO7dCTEryvDr
RopnavI6eg4D/3X+lWBFbzPu8sYcbP9lr9GEkXo3AmcHS7y6C6NAn43dptKj+fJFqDDIm8qQQPgo
2hvkY92ftDQ0Z2ijx9kONFp36lC91WGqBRMqQ35O9HA3ffqlXePn3Its9uBdZjQfwQkUQqFwNYtI
LCcKO2ebHBXnOSw0sbB+grWNhAuqY+R1HshJyGn20bd3l8AosP0bFA9CRQt+2g28chG1KN9EHSLR
qN61+k8VA3+GJEJkYJMJXCMfU0SjiIbSMtlx4Jxu6h42Mhbmg8wgS9VqG4JFsYSdRtNCV0wdtMaL
Afit834XGuxgXpYGpIYI+69tgs0qcJjzVWD5i3Vs2euPeSNGZGl/Ryl4VgzDsKbR1/lnYIDUzT5l
YpQf6E/nUVF7LUVYHtQfvNScVhhwYn/RTzUSH1SFafVCuHeV9xQsq5fFVmQ7ZW/mmDwmXgux/dVb
Z4J14AXRShJei/GheRhUsS/RUXLO+avAxgvX4T4CeSwpOGhb5t3yv2m8YDAlj1c+Ant9R671RXYk
4i81TphAmtJTgn7DivrLLrG/Ov4zblRXl4Fi9fL1dTPIGFus3yQ1ypRBb5zebkSiEfa8uwoGXER2
lP8LQjQ2uEakvAl2vmIMPxVCaYim1kn4QsQQogYppXm0IZoBiF6vo6+9nysKgaSEUwqohLjTM/lX
qmrdkbejZIJtURoww273fsNzQ42nD7b1CGaJE6UK3Y/2xpcujk5R/Hnujhnqb1ZXaaxrYO3l2R5D
rDTno8qBETV9CKTXY1GawuqdRI9S6TRBxTTPzeqlPd1EXx24T8Cq2IfPxLdZCdcVU2uU9++L7lcJ
nE2nAlaFcZA6Y6NTrGQZM1lvnLcLHwYKRW4gGY1Sw7PB/Il5uQ0m6h30odXih8V61IMXWvS5t3/t
zUiMuwJaF4F+SajVotyQD/zsKXV/JJQjyxAz3HF0d7EVotDSWH1RfIUGjLS45vvuKfVLzVLkbgyp
Ssig2bZs8swhi14hO492CJAKz+hAfX01xPwC05L46LC3Tq/B2FCp1kZ/KlkA6MNL2FcLkIFvVyrd
f2JqYCJTrOnMmOUzPvWRe98cEg+pRswwnYsaj/CV6tbCPAD9uO6zLWMk5qIfzMwhhqcdnKVZDxaD
xDsTHc/QVJ7foynNLf3Bm7/lZOKr/0PqyVUVd9QtHsbLwtaTJeCsJq9xRD2gPzKFCoYIpfQIBxh+
BL722uZnhn9xGVhV3Lvj/R8wfjs14YFXtuA84EN8wNzhzAzf/mzuK2n5iexAwF9eVfwQ24H1hsTq
d3OGc1pvAuhixyx0agMTwDCNDetklG28x+kfGAh79Z8cerWmVbbcEDdy8rGC3r6yZTitzbMiK9/M
ihpnWYF0tPTY2qrYABS4+/6u0uteCBppPTtzSwzqIahNnUSv2TFTR9jBY5sC5MJyu6jBmRKeMqaW
GPZlUEUb3FVuvqODhw+UTfezIam4+dUkloJVNWapwrrsBMSJlslAY2UNurSigVopACTiz+guDOu6
2ddrx2pev/7flrRmZucno3qk6r+wuCdxiT/66zV3fckYk5KFiF43zxns/3Ou9F2aJHJorNNmi/G5
o44G9/iH0MakudxQYJma3WX9WcA2R8zkY40kWmWN1lWrcRtVsH2+h6t9Lvg9By0Yy3nOKFQU1OmW
1fISgvEDgjnBEBEAsYfiVFWCvQ81K7zJoI0gpD0YLOhyFTEGVBEN9PNn9xnKXNH8Zn3XHrh6mclr
obNrdDQ2g4RNd6MJCqsmhR2I0c96kJrH7BQp42sdapITOh3UXJvbi8nO/SopZkksVKnr5CUxHT7O
Bv0DssLM0Fg/BBNWEbmtmY2SOv/pxzQ7RGbOYTL1FO5EGcNdaQDB1Ns6Q+lgvSbWaVBFtRHVaYk4
xAeiL0lAbHxbq8fS8dkmCbiW3SeAP30SFaFjenGzjteh296RXtt5/WTO0t/dAQbrt2fY9ORu/qNK
Kllv1clWg6I4R118E3z9/iBHV/5gZFD12TAtdpbzdaAoAvPTfgnEwk2f21TGCDu1BJXVz+yS0+XN
6rGiK25v3jRn4QqubAwva8Cz/tKlAvBq9Wg1jqxHqYqoEEldnbfeneI/s6JCencKbya0gWkC1rbh
yLWzBpYpFTvDaREKcv9JdcokxyRYyjO5Ugrra+anR3bp/LqpPMrH6pExFWKlDBDYwQUKn9s5S9ZY
T16uwKvHeIHfHJZVHnnXmCFusnoz41FiP/ReOX09Gu9Z5DXB1NXLd5uwwFRDxWlPdG1PHC5tbl5x
9doaZiLfzW7LA/Gn7esS74XBxhtrjGdhI7CQrcU+Orf2n7tHim2Q+7Bhc3wQnydB3PU2iPHzW/Fi
CN91qKnon5LWN6EiR2bqgBz3aAGXnHEA3PaplK5PCKeEsufmzr5vj+aEJ3C25QmcZvGsPurED/7J
PVrq5iT0TyxPCY8pJYXyM0XlCe8roHkZYfPfUU1wMVYkmpinXwTFJkikUJl/f8KEXJggmfCkYR9D
LsWbcYoj0Dj8ZbxQX7JRm2g7cjHnSLf8pidiUR8Pc2pjA6jT0ZfII8qhrGAXcGaOM1QoCn+I+/5T
bvPeArgJDkO071ITY0MhR90h3cwrJlmlSw6D2Jkc85dlKc8GtgAURrolfvNpGatyCJiCFtKeP+Ps
koo8+zd6eREnl+T57PpB5WyPrK6d/DsCNWYpfIrykg2qqNIzMsRRqa5FHKdetFuxahblU1W0ZNMr
YH31YIiCU45WF6rPUVSH+ixJcIg5IlkXUT0TXbHyBhI7nCH37pTH+NtFa5eOSv2EX8F0OFfC7Dif
rAMjGBssiuvatEjO1NKEKS6u7pEqnyp8sPEW8BezhwDyFKXg6FnKrwvh7sWZ88Jnfrq2xklAp8NF
IAp+jYhU1jLc4ARuapuAKHSsy2H/OjwgM+MPXd4XUUjtbWOwqas7QT7ubkH8jSPOoOR4PLafizGo
7fqugInIn1G6IWZgHIlN4A8qtGu507ifynF8BZpv3CXX/t/pa2ZQil1nNciJQvttt7S0F2ngfAV5
6GxZYATC/Y2GH9Lc4vD23M0Nm/YpnIQvhTi59EBu8u8wS1RTw2nWWvDYsYZnaEQuh5BYd05XqqCD
eVgNTB8jc8JbmKR3QLtkVNIem7Or9b0wNvAXb5fU24vk84ugJSrlVsFDHZ4+HFcCqADucFfn3Oem
zekCKjutVxkg8/b5dS6fdyEqm88SsSFO+WQxRsBDr5khYc+hFEd1bstUNljgdjU05vg0lW1T+l3S
MtWbwi8gKQYaZfUrkHSF+4FYZ3h28z3hMzDvO4yptFIGmLsDkNqwYroRKHWR8d/JghUkHNPs3Wi7
pYxEPnR5sLQ4UZDezCdgYbfcLHxoiZyaM3ODsiGNUbl4sDUSwvJWE9TJPPvFJkDkk7JOMSGgLRt2
c+0N8JLMe1qkp4Fb5p9HGfRnOyZOzuRw9DYeJve2xJijkXFfsJBeCmEhXuGubJCVrHFjzTTQpIUJ
SC/xbZ66tAqnNjERxPyLx/+nUjYIYuXpPxiT2xqRYgasiU2DTTFecJFJ/bJ+OXu40Hs8YozRzsUw
r7NR9GvUnUuTJxcZk3eAd7tmOuD2XdG9caCD20YVkxh8KYn4xKL8YlYiRKIKw+ZAZdvgCxvDfmTO
/yO9eU5lOLazx1ISbeUEgpcXxDofq/drcDuJKyX3BT+ZyeVr8pT2J59NveDszP2sCN/W3gKC//Qm
kEYqXmGTDyWfup8x/U4hG5VR6aMSlt+x/uouwqwYG9l+zOKs3dvbT3sflNex+GnFDqiAF3HkKo7N
+AlkLEDFhJRNxkoJzJ3/kD7A/DagMivjbogRT3pekGPoDvgT33U+Gk2liQtyFMw6XT+54FjA/jW/
eYamSnHVeSuzLcE4cnlnyz/Gt7hK8tQuQ1YHFZGj8Hha10/vFSI76354ud0NuozFaRARjmxsLsQ3
NhoObMoXNjBtOU/Gi0BHTfXrkLM8okaARozhPCmEg1eG+Oh8XSsuM7tFUARCc+Iy/VUidsSSYwoT
ByisRXxkig36PrrMZgmL6ypTIKAFZUOEbn/S1d/8rpe3Reml6jiRz3puYYqlVZzcv3iQIOLJFgzm
hmrboegPu97TCv7E66xMJd5/Z1tG/x7FYfeInyhDJEaKIX5MZRIr9GHi1z4c+aAhguhu+wPvl8of
qrxQQ2PyqZypVg17uyLmXYTUvJ58JqSrrZqv7QPhH+1XNFdernCipKg/6YuJmT//+FS6XKPrEjuj
K3iybcXyXlBgJjjJao63EQ666uswmzb6MIY+Molt6Z4J3buiPhuXLfEYkQcgoPYAtbU/o32LcVIM
lGNCAGGInMkI7H4qp7ZSo5Oyk0Ay0Hcw51jwblnrYuPQoDV9nXCFsN+4MoZbqaFBuGpqhZD66nsW
IalZBmBqNHDNchTmRWSOGPcG7paLXAtmWnGiPW4BUbluKdt4YH4KPXCHbM259GxND8rQA1+2VkFu
GTXv1oOvM4NcUzAnczhQfERXQvQpebeHG2I1znIHjg3mUnU3qTEF3sDssnfITy9cVciZtEs8DgT9
kGoD7xzDnoGzjzJg6e2tiVT0pN7R7r1wgS2/3Mfhj5IQ+qJmviYLkd6jDtBFGDpKc5WfM3uXThOE
I0Sq9eAn3r+8TtDuw+7vzgoHKBpSQAJf4kyiYXTaz7EcUtl9oDabXXoOBI4N1MU/vczE2MQV2Com
6o5R6TmLdtplWHTSRiyX23o2NUFZUG9JZvmTTI8bcFObvZfPKX2Ssba8/cc11lBMxiNWWVtzqc8I
wv3xgYqmAqhiziKrNSCr219VeGsDJ4FP341QgsLDL0Q7CMRT5O+ADleMaZaDHbHa5OrCx9KfTtjP
92y9FXF9x0dGYCpJ0NRYSuAvSnquwML7WoFSJ+mn4SeuLCqP10zQzviUj8h6b7+gjQamabC7n71m
o7HX+DV859XpHPvoJlv/oViLtP1mwcDGqbhvqNSoLqc+ka4DIR4EmmnzuUBJXAE7J2U+uMKJTByn
a1EnywIAQssBhARRU3s3AHHEDOGh2E9JH/7PumxZAFjvC867LDRSe7OY5uq9hRq1x5zMkz37/o/V
LfPa93X6VOkNOlJWRM9dc36H2QTlcXoqyi7nLdWIO3HG9Y3UJvCSGZsGFeepw3WOCEKYqGAW0x7w
Oh63LkCVO1RFka8y8K1MyyMakpWO9pUNO/5L5L51yuXh6Hq0eyF2q6sEofE7TnpiooTJRBdcbFRF
t68ek33dmLY+d9kBjEUs8vLbieN69kSzS6mDhP90HH0mmLguykpG0Pdm7LEL1mgG+V0gh5e0/nG/
KQCrUrg1ZsS4wj3Qw0Qok9tTgyjwphjCOwFJWcVQYe5J2V0sXP3RDXvFp/g3oOBblKVZhqPZnmfs
HI1x+azoTCAMrIYesf04s+H6z3DaufVk5erkgAlDASxeVPGfxLiC9v0ZLL9p9uVdc3gwNfeZKh2u
f/r4B3hzmNWqDFLm/fX2vVR2hTFeLm6OdVPMzED0m2nzVTRhipnj3+E/fcMhwKv4q2Bl2ARvTjkm
zTUhJVtAN5MKHDYUkrqy4YP2nYYDqy6WeJ/V8XivNsnkwOgOFNo9Nvi+YAN9djNepg+n2vq+y7rT
yyzbDizc/XjEOin7lwhqjswMjzrPM8r+wRTR/4/swOIyA0Z8iYCqxWBDUiKRbzbk3z75rVOK1jAw
2BrY6oRtKmRTt7cfQrMCRuHPo3QWyUTYhIIL35Ozjz5mxW9KmdQwgHvCMa3BtUhFI+dmmVsg+OI+
+2TjdIiMCLFKZSgKnPgG8ovY34lfZlmTrBicgsxSCBq/F662LRIenW87FQIvNuWDVg1/VeS0Zuwo
1jS/M5e6aDL20MmeQ+dOmVq+uARryp4+uRPCtGG7Rcv3v3OcKZ9NsMHK/EoWc5rsgaqlb1Tpiz3z
3D3WF6yqqcelgWXNehMc66hID13WI87uktekEeyOahxRb31UBJVC+Z7t+ndocCQoyHy0gX7ATaU1
tZgCyn1Eg83gZcGc5GINX/m53UfpHnPTgdAh58o14lAR39vuse5Sq6i9fokPVivdObokfVARTOy1
lNNpkVDJckujbP+frxlMchuoRx4GgGrhBjGmV3aG0YbAWg03gWh/w+dr6AMTxS7hjJZbAX7nztvI
YOHc8waipmT55GLKOsBs0QTF59vvMRZLh2w68p0BF6SKMoe9nc7b3Ni1zPuznACTAZWlMKP89uAm
nPw7DOAWFeilEU4yL8rhHU/d9ysLBHQs3enBeqN1KyPIMzVktIb5dNVsBA+CPOfqHO6GIm89cAo2
Yx4MrPb8z6naF/Cew1vDTTha/YE7y4T3KNmavEjiRubhZ/tGzy61jHtJ2YWd/92YAz3ibcqOeVGF
dbUYHR6fOstt4JR41ZTq/RfqFW3uIE2OxpRJcJvaTYYHJIgzTCt3ABQbezV+UYcn8pet2aB43jtE
y9dhp7RiUKhKPNy8L0Q87llW1iLtmNj7DhqxljXk5n95Jt/4l6hJWjhFmo61zuYlOLuYhzKQvcrl
YQrFW46WIDlgOCqaR+h/VIo5bgzNm9UmvbCVz0k1AKWzxM/vz3fSgqtbIFTV5hsrTyIC8RClctUE
TF77oIljn6QH4sz6zEzb4RRgdvIQzguBJE0pbd73r8y/At9O8z7orsC9tWJ9xS9L71TdImNxWJr0
cSEr1hgom97AJPxamsUZK1wrSyyBzNckhor2lFVTqtfO+bzUrza4a5odG4x8tJDRGUuu7UsaFCR9
cygEsmOTtW1KMf1v7jRZN0ryriKfAvg3XHlvtdZB2pKb6ZbaMGD5U1YPJgusknjhABuhufXAdorm
Ka6LzZkNBHsUiGdkeGFwRIGjnZ9JDd1puZzXQ0UDwEPNa874F5etNDfnJReLATWimUM16FEZl3+d
ytzjGhlj7LThImyfJFFf32SWD29Igam3VrwGZGPFOfDOgTsOaZ3B1RlQYseMQ4eL9nW/FsXYkb0r
qBjAznonc5VtrC+fcrM+m/A25dreuSzTXPGKhxvai9l9TyJlF7OQXKzmoHHV4Tpbqy3u14Ah4i5J
vtaedfaZp9FDGRqyXi05PVgC6dj2iUkbrACJxKmFSvNfhjLJdNri4zXfliu8qnpG9Dgv7vqFr+YW
q913Hvdet6Gr/4sPDlJyv6jwjkn4bSfYXdemt263L3y5qQ5jaYdsBS75YlNAQJd9xifhf9hsX0eF
Yk+9PAvdcha0ywrTmOlSU3sVZEtHxDVKLV9AfcZZqOXcE0clzLZgbj8jYtZ6Kq91wQEVPtWc8htI
9Bq31Y12npbCw4JsczB2TK4HcowQoNi8K0C2alPbIEZtNY7K+ZL1GlnQq46v4rBN+jW0zcjqSsIj
JeIOvLVxs/nBN7nsSM/XiH58VV1hb+oxXkxhCr84cb6y+WyOE7kCm301gexhTV4jkOEnx/47N9xM
A3BplQprGTSVhzd42JeHQA1AnXxX0JKvQgDoT6TdY6iRtz5Lf18nRsEJS87/zkjeZlcAtMDp7U+2
Bsjl9jG+MsUpeAwKvihApjYIfAfz8JEchDEYum1Cs5FidJbJf6FasP+AfXlPchiqJrI4DXhytDzP
jmrwml9vIZYFB5uMTdSq0zzLUjwTi68B7gGrc9grlCryCr1WgXOtzPv9QrmEFAS2k6u7EWbeBvld
m5a6+WalECwerh+bVJiPb2/PqiwURKAWu115qSUW8JOphfhsslp5DvR+ZozmnK/g+uic/yYQ2CcU
G8ELjIZRwwZUG3WWDZeUFUJXD4XeYJMf5rSQWmlZVIcMkXwAyVJy0I7RpnfSzxa/Ee5UmUoG2lnk
DJF24TeetGY3yTuRFT9ERgmgP/PTfc/Df6uHicAyM4vOdSTag7ZpzPcOf1+YfXxrLB4iBtGsfB0H
6IDpJTTRKKphfwyGujTTSdPwvdg75lQOq1pq1dUMqib7whDkjB8bYIf5aEdLlOWNvXHBPvFqB+jt
BrDk/UfH1QBPdym1wBL7T1ybNRZBnhQkq9bD4BBruOo1JdQPV2eVWgYAZaGfF4niukCU90qf2Xsv
Ggku3LVmGk1DMn5igwAbdGfuPGg9Vh9469d9/xicHdNh2McPv/FCpOv3iUAXfd+51AfJLvgY3Rb8
QSec6xdn70jV2W9oclstx8mLwDSLDRU33jB1r0lKY7ecs/WE6TQZxhxqEvMnLE6JdhUvoUMoiJwK
uKu7iX1OTyK13F6StFeIBS6YfBJUuYQKeHs2YiK9tTJlkE4a585FOVrImojYNYngmibtw1tpRrFu
d0oPil1xcHu0aBuToGFBm0GcSsOGwmL5CqCHuj7+zxqtBln1b35ysrjQnL6atpM6fJbgu3Cfd6qM
dpznEE1xBpo633zs2k1XL2tm1s7ZhMcZsMy8FzHlU82QZkC5XhKQQecVU00+8L7eL7oXyT4zZOZK
qvJD2eqMMJYH/8DBU+HS4atEDyuutvtz6v103cNZw08N3lUYW6w8ditP45jZVtmNAOAlI1GT/8YY
4ozMhTDZCQNXO0RLkPyU33+96B/vokeqXh8l6/bOBTGlWmJ/BP9G4uA7/cksISd75exMMA37yCPy
Pk59UHmEu0nxRsfStjKNXa517onoEz7cOu+uCfjjN4KLMTv4YuUS26OibpLir/+XHzACoRD72Pgk
m+Qj04sNYvjncutroLIftj0DFNGoWGOAGekY7LHF9MwXbs6WHtRt1w/QtiWDBS9ri+Je4NceRBZ/
kXeM3MDAVWY49GuVCcLbsyUs9rdohslj4LDHxts4Srk/dQ7NPC4RUbSLlZuE8gIMMqsyjfSWX6w5
DEMArzGTJQMdzTFL3PXfqMth/o+tYC+6MRIzPFGOHB/ds7PQW/7Jb/Il8tfUHAdr6kTZR89wPQBD
Mr+CG1Y+qbbKsWcGmmZUBOBoBh8C3Y0mcqnfa/879fQ0Pah+Pm6cDEZ+ifM84CyUsr8eFz6vkf7/
ctF3hv4Kif1XplkGrX8+21W1gJvSIDM4vlZrtYGQZi1qGnOHfFK2X/Twv5QnXyg03acBZtn9YcL6
jexqPcOS/4lJrbu9BjgaAfUcHl8Yqqodp/dl/f7IIg4GkgHxn6i0kJ09KRLKS9v6aO1rWdyX+cdK
TvjuV0qZJpZVRsvrrI/H01gzuG4WB8Un1EghcfIb/EEL0rI0hp9cEv/R7Jnn5awsFr1G4aqaWw4G
QPE8eK/stL+nLDlHm39k2qJFykRSJn2DcF3E0OyKH8JgZZBWCd3lYBpmc2Osjfq2hNNfrzxxgKwf
FZiVpDY57GJE7ABbhAC+pmbQg4Rbkb06lzQDD4EtNPoPexo9iguLD4o4e11h5VkcXKWWMun357Lm
jy5HSEakRutuONwoPAM+urHUIb3VS7g80UyeKFl7Nq1WQAwWmteJ3HYvAHIhulxGfRjs2nh9z/41
4iNBkNU5xFDmz2+c8LQSPTas/DI2x3TMVwSaRdJgLiWsn+fj4qTXzq49iD5EzG2t4d9/K+/NN/pj
xqYlPdsudXydtGDwdRz8GconYN13v8jE3lCVoCeqJyF7xmVaay+BCpcZYaP8zDaW7pPrpgogvE5J
vzSxoFCaG8L5U7qJ1voBL1lCKUoSa3VSJPSwYvUlmEHk8Wz0pDKS+NViWRAQY383jdjKHAo8VqGl
HvWi9/buNQ+zBXFl9tQOERRqLPry3fncpOo2SiuTWA7HRG/bOgCGZAGsQXBwnqcQcrZICiW/O0n/
u/mGmSeepv2Zvr20T+C6QDTbJs1pPrS2Cva78BZEFSQ5Rz2KwVd2oYhdZj9KgWKlc/TruaK3iLkY
BtdiwQad78/LWRxYxs/PPDsMUY9TkGWhsxo7Iw5T5BfRVKpZKSC83GUEhZEywpoIklFJZydaF9Oj
9pyKm6+ri+57y3/wV7WlJx+uvWVnapVXkMpxdh4lIgE+k59juB98ii+1751I6a+jwgzlfN+xDIn7
pd/6N7KqATYEUYMQkkwk4ZLDfzBjAcrCKjCdzqhd3f/8kBYH5QHDwGUPUI3AEWVY33e4u/c2J+dX
edG/MRxN3QCodiAoQsc0v8Sy/KoJu44TqOOeWzwhV2MLwA7/uj1lGBBkOUK4zIO+/LqY8THlar04
BxUFMtvkw1o21MLK+wz5P8syKbrWqPVPyzKPJNWkEpXY4yvl7tA/g3jewS/hf9v+7l1N3Z0+UnkS
qcS/LPh1U7y9tbyYRSl4ul49tBlGTCJ0uv/IL/WgmcLuc5ottX1KBRADxB8EOLYJOToQd9bbULUO
PUBEvleNm2qbzwx4OQK9Eek6GQpFz+Ld+Q3diB8MW5UCDSxjEwqydiOpoUGeNH73wrga2DInV4jQ
qltFvNfl3G7EMqSYrJ0IQDdoqJiyBc+okL+LdXkMkJ3/zuU8Trev2SMyFlAKuxRe6+kbGa+x8/S8
oImkqJ12/zOPP1ULIJvuk9CY6zwze32cEAWmdzGRrb28U5SnfCG4wZGtDjPuoTrLI0HVMUokgl/r
fLnHpYmYXev949+88Fhakn1gj7/S6iitz105sgv7Zi0wDCeh3rpjIxaGkLtLQSpuP20CR8NkDej0
6L4i/J8nJ6mGqTpsSpHcdZhxo5M37o1+qz1pnPADTnSSYbyS3DJ1AXsTaia1irwwf05Y6VzwR9lZ
7CQ1ZdPVW1p7PBv5c3KJPpt2LUo0tRVWuOoWvil2SwXOgYHASh2KtPa3h0HeRx7DongZOTvWHr/x
ANiKThHlc+dxcSJ8XIZTSvoVIUKGraFW/Mv3lle9F3+UQk1dttu9e3Z1h+N6hNHGe0++1VjMgyPE
SP1gRbJa5Qj/9drj7V0sD0iuzrSsTKe3Sdw4fM+9TKyRKFrJEOHR9sttLk7MEHSdX/6McjIbkHFM
zBSOgh49aLesJbt2OgNq6nr4Hv8/WhubPlSe2IFchD6v2H+EcCTO5hynC5fUDqf4IlPZ9ZtGKrGS
Hi+5RAzgjSwebWKnNOm5LUL6uE8cDa7Ar3S3+4+7GXmf04Vbts4FQCGKJW19pPTaIEg8TpUNgg6v
Adv35YTK7xI+B+gnJuRCRFSG719Abq7m2gZt6uhk9jjZq/+S9H39rN4/Ty0ni/NeTgBVzY6Q847R
YVS2IlVweRQES8kPXxMD2ZGfXzTmyrbeRPBANjBwzkI+oopJyP5gP08W+qMS3XFKFNQVWU2wEUo5
tp1LJ5FvYB8f35Q6HdAaliXFwck1g6+rd2hWKtEmnkjteL2jP5J19l4JQxZlBeq3OGEToDgexy4/
tFjWbeR3NPm5242lvOeOcwKVmKhQRLYC0yVvmBwgXoxVZMvyzAz42d2rr6qq6CnCUXK8Wa4rJfd/
ZyMgnuvxDiw7clzPVmVZflrjyobJuXC9L6foSm33/c/DSpGFGMSxE/ZNqpgIN7a3gwj81ar3sIzw
hoKjDOMfE/cRHLvuCk/ioNzff9vkzeTi+LjUDxAUdnsci/lrFqxS5uU0AitpUYe+bWgSaV7+Ciez
4uzbS70ymJmMBHXArwuareAgsels7S7jUQIUnafDiBGaFof1QkGNWt4n2Cxzi6Qu8KCTnHndKzH/
93uTOmhqCGEwaFMU1Qetsr+WuuoH2nQe/R+RudHGVKwSQpqPFsy6cCO4bhxpt3SE/McUq8h84o0M
61v8BX89baRnC82biG5OtjZUF2F1v0dr22dNrypa8IWpnp6RYre4B4J9uhRUCtzpJyqKnvGrDQu9
APNulsYPQ2d4ZWuhcr8a9/vUXKHPY5AyPzFOrxR6zYv4gB5w1bop6Ut9R6LE3ZpK49sHNQsAzjGM
FquUECARx50ZATCGtJ0TppPcoPFHbhrXMQ9F8l+n1pMWdHpmeTd5fnRhHsDGaEO9Gvvw7FOMwK51
pVcyxW5Ql522z5dXwd280y+TCWlSR/fBo7et1l3xDwTwINayj6QQT4c/pqDr4e27w8XoAfPcbQq8
Yj6+KkemZ1oXWvgh5IvO/0x7b/9B29kVxNHsECfVByjlyCJw0/0TxjbKInlyTBuPsymx9RAG3SD1
fzEEfVolsP+cXIZJg4YVF6zCaZnTV+q/pDE1gyBXXo4pdWZWjZuHwfw1Awm1MqB3NFty922RP8S2
RinRTCKgXwsxVx1oLtQ0ggLEIAKL8knpwrrqG8LxTGRxQsbEhyPuTDMI/kjcE62sR7RkD2A39HVS
6TU4KYeh5rzW4ksRlPjnk+hdxHDIfdDw4NdxxGsZy+Xn80D6daUUosgfoEalNo+chz8HPNIzqjY7
EIxs3sptVv264Ct2qGGx7dhGAAupnVYl4HcKbewy5XhR5xW3cGUE6lYfDPL/gE3V9d9U5szJfyK0
wFrwWgri8gUBy4Ydfdil/Lp7ffca17nKhaF9fJS0TbNkMQSF7lpmL+e9bfQOH8CUDdIBtovXYzIE
5zL7JJNRqkihlJJRZGoLy8ifnPiiLOPnfmEu8vtbayRYE1qPJTD7UgKZvbUNnJo7O4nnqrAqVvz9
8PWPXej6doPnolTkvx5TBuabacNndmC/uRTcIPkwoabEF2IqbCrH+MV30P/Z9Px2Wp1Db5xmck6j
nwd7pLNxqEDD75n31en+pkPUMRLuQIWjKLuBX2m1TMaBnBxRPMdZopbHbhyCOwbeD8g1+I8p3UAc
iv6JIQuqkAf6Of4P7uMkcJBFqAK3rwWICdAPVueqitf1nPP5KG7viRN6PQ4ZBGoHcrXaQZwB67c/
noc9JMTS1zmDYjV62h79sWQAUrZvMvhIijq+IrRa+8CEuhVjhEnRiLa0bFm/lPN9AreEQifibW5Y
W+XlkvwSrYK2xX6tTtqzaRPXBOG5a+ra9OQ3bEvv6rZa8uA6jQ+MNIL2HhpXkupNRqEpoxe93dv4
VIB+nwDCdVxKHaiA5hBBN3DmydMC+axs+DP8WJ1ztLx1CsTIQcJ1u4yAPqSL9ROggSN1UxrgtWvA
5czjQtc0ZURSQt23i0uR8iewKk7NJRlh4qyys3Cpw5bw3Q9aoPq0gbEVcHkDtYQct91caLj7fb59
oduJe1otpUfiq1xscEXEBfuWwfHlGkznypVajMWvUiAy94y9iCCfQG5nNsq0O/bSwCmRUvEhH1tx
FoZntKR0toEBRH6zcYDkK8jp0mZeot/zH8AbGTXB1AjR0k/5Ggjdmpi0XS2SckJCBnAyW3TCCwah
q1d2gZ+/393idSRNSjOQGczsEC79XXbYqbxU2RGBhH/9UaIw2c1TyfBSoidw1P0eDzUll6ooOszl
vBKwnKpMJZ7BfMZPwtoSQgmp6qPp7EpY9Ds14p0rcNWtFwegKTy6pLaHIoGZZunyLs/CgvrU9fyo
WdcGDKe9ne6gP58QMxX8z7waKR12pQLQG1tD740mw5NlG5ekzxQyx7MtQ0DOQSnurtZnV8d8Dq2n
64YXa6E9VNy6RJueqIPxmN1HAMmpvT5Fdky4UWAkjmmLkpcHMXnVYPGwWbQBBq82RcEemnY71jch
7Qbh++JyQF7B677xXZuHxZcraoBYkUq4+n61CAGo74JTvBwJqfDzHjZL9dE+cFtitAGVcanlHiI0
9M1vs6wkCAB8SyrSYS7Y80c31YeG0FN/DHJYycAr4boNiI0o1jUEdw78xKeg8mb55xNBDcnVQCKo
+CIu0qQHrqZMzqCSB6P0XU6BcroeuOpETTW4BSF7c68JifYCZ3nb7k0428hIVBPTGlvbcdzGvxUn
gLV+EaJFCQKLHUfv1BbgiZP9K9hx/lliVl0Wx6AvBtSssbwG9ASU1QbO67FUx0Wrmhbboy44q2/m
AxDitLMNu/aC0UiZf0kanSa4wsfTOrlMbvH3PM32xr2Dkc6gSaJ9XTk0WNBeIlFCFaEci/I8RLTA
BbhHMfKGmoFssbtpCIZSbtmr44bYmIxnSAn7s12cmADiKysisHBKPLKKEqNBm8IHPwf0Cn86Dc14
mmz0ff8fb4JMW3e8s+pt2BpFk2UXRVoLDf0fT2yBUW2ezfUe6YtcKSIhzEzWdWUBEulde8XljahL
9aRTXc3nMI91RCPqER1RbqyH9J09uFHXLQtzfIC1osP59BkW9WoyvuAprobhoIQHZNE5e430hyxS
ebNRF3lcJkkmC1VOeAg3FwuK9bNnCmt/3HXza3zef3Q/AhIyzavKDrvsBGRVX6MN2SYwLpdg3EKD
DMx3wl0orXtY2h4Qr4JWT1a3hJHfy9bWy+6qyyRbvdRRMwR1lvamxg1J2e0incumoXO/bQq5gOv2
+q//uw8fcRphlSyfhVBPAnlS8Kio3P9ZRAAQ2Y1VLiQN8IYOfgJke0s7yGUj+36eKxpq0+HJ/JPR
QNPu0XpufoaF1StCoS28S5K+zScGMxJgk8lnJISlRiBbwgSaXN/nidxZtynYCIxHT8bcJMquyfJ6
vut3yxgJmOJUg3EzsOU+KS3qz8XIa1E0vNc/7oi/IDxg+h6nxwFw9yzaN3kUZP/Gy1gCX5Ui+Awa
W+ZwYxOTn8Pq957wAH3ixcGQ5dxAWJwnkc8gNbQ/W0N5appqnn1guP9iGqFJ9MZ2RqpbkDquhYoI
9jrsKa7PId019ykPCDxiJPLYw75y2PWOQW+pOFkRkrEqHStraUCCnkh4VG+YE3S4q6DhAQcjmPA2
7SS984ArCT1iZHq3Ih1aY3Bs8yjdZHB9DBCifYuCpEuIvW25s8xrcKwYmSKzpoyItinN9PX+lDaf
D2qpvS+cty4FuiTFKdZtazu7vibrEG1cw8HBQwgf1JUI4F5j5Uvm2ytvddOPS+ppYkVqCoo20LyM
Hj2HQd4qFhmjlUEpoElpp5rz5yp4BQkw5ncfie100gUFcC6relw8htmlVQGfBearYNCWGq5IbHAq
0tRkKDp3Z8by0tFbf1YuGHLB0TpnepqUq/zEdnbJaw3OBHKg+bWvNT93xfZJA0yi/WNjtyJLpjth
lmN5SOC05X1jAtpSrbTbX4UAhNgzVPLdT59HKAkPuWyVPtQsjyaRUPXMKu+42RBI7mCQ7qaNig2j
54ZifCUejFY2Rvx3r7FlnMLe4vfntgT6VSAts3LCa5W4dR0VcWB4dm5s6naV6pumcVWzYXJ1fc2u
u816bYE1TJexR4EXy3XTlq4YDqzqedA5/QEbh/fhoA1Hnu8GlS4kpsrfSUbtEP3C0Cg0Y9oI9Y+b
zJ7hdx1iPhw+T892I9nquK1yqKBuwX0SDzvg6tQI8KiT0wBHMpGLrF9cSfNDY3iKPWjDjI9CxszM
daDiq4u7PA+sIe+cAhZVwTtEEeNLAoMALcg6yO30UEvbD/WkCROh7wRb0K8aqptqVZIhhsHafIQe
9IKeBjDBrRKHDGNpNUPgwaxgOBT8VufjglT7AY2SZ62v4xyZm8yKy8eGIBVnZnlC/Gg6am0z/Rry
KK8OoAk4/jnXG2RVv/59JxTV3ItjrcSBD6RkoaSXufJuiqQD7+OeLrq6wCs0A27kxCPVFhutcQmQ
hWOtU/ZZ9Xrw1xsAm8OhMBYegpj3JOLgF+lv6e3trpl+GReJaEwyQ7tsRQ+tJBZY7h1dGRYX6opn
UeK0C64wZ2/S3/7XITeg14sowNFvVtfdWUODWeeg6e2Vvzd+wkvH+4TzDi966gOqWqOTKDv7Cr6a
/EolE+/1e5cm5krbcps5RO1mAo3yMXFVyUnGViQLqqUlZn9JQU7HFqKaxMDS/nqv75p1utiHGfRt
D7ZsmKoUGPiBZg44fhOFE7+XBBAa5Pp/vmIgrM+WVhQ1nCCf9n6mSJB6skKK/LcO+Q3n4lCEXbAB
Lf4iB36ZN4BkR5m3p2RlABscNqdy7y0L5VPslq08KL3D1rShn0O+PHoNiRtrnKzVh3BnLT1kWYYJ
4yoXmn3BnV7hWr9lmhIiIjRikRg/XVjqX2Juan5OVIfal2xhkSal26IhgLp4o+yGekiASyTLri0L
etOVsB/aX6ivRzODU5kcp6rEa3gqnxDJK7Qffwe5Glh8uXWXYt+LwTHxr35N6Pis7D0leF9k9c7W
trFKE7HIdC8eefh1lLtqeAaM7OCBbqtvlO2OwOiaptKCwF336NRgaKxfV08nyfZKOqHWpgfzYc35
ev/QjSX06XDvqtZ9SNSZ9R63lKtfAzZRFWOkDZSn1A2Jaw1dx7topQDuPqkPRc7Wz3vJTHPAERK9
XYj99xHharmeRXSkx0/tmOOSHrsc8AbHFIKBr0xA4wikNbmzgRQ83f+DWW5W3MY4tbTNHjYAyQ8b
vxFsiawmt81K3z8DulSY56V2LOPgye5PbcWGhKnR7jq5uFMF6K+FngO9Bl4rpo6KOphNG8wDcKww
N9SahR2lqWWxJhF9Vr9bsUtzbF9XF1To9+zNq2tTzDDJdSEwM4ct9c7zg1Z2yF6GhuxQQtS5M/CG
/3Q18F26xMIZNsdA55X7IdWCyPlQ5ElirYtP8rBdM8ZJHcG0wInXPHNLdsmhtXgxp51aSa0h0Ybx
Q5RLqGQPEb8NIZm2bhH/X+jP87fqWd5TZhFQ7ADlt8UdWRuIBAJcZfClLxh8cXpxDdW9FrYgHl08
/4e+/TpuUStsQV5tJvsdqvvIUpA5FELLvAwt7gvInSS7JZGe1ySI8bT2Lpou9oX/CmWeuGVIcdcY
OfjStpwnOYbIuyrYIBUZuyWRYNjYWh7icSdC5aODg34RvypLH1gXzQKCSA1K5FrSqCQgsuWKc0iM
3NK/dHb17a6d5hYIFfXHUVHeSFUv3eyJjsKj+nzZanlIc8OIqs4lTsPz9DWEG3j0ND6hHYaHAlv8
acswDx7FI7m9s7eba8ofUB2YlOtwdTVAovnakNEZWsQwDw9GTfIeMY8Qf7ONp9APxgdrflEc2yUY
qLs+ytaxCH8q8K+pgNQciv7Ff/AoE+vgkEsPkd6BxEgB/RLCYHxmpTAmB+KwffHJvCdfyqpN2i+6
ggkvm4TRAlh+r+TUv4XX84bgR4UokPoZLr52EiLaSsvk5GyWe+HziL0r6+QuCbnQUoZ96MCOeTJ5
yQGCPcxNt3mhu6jWrIFg59vzCjEQEBkvCw015Jdkdip9VS2eqrTUmNcEhnQQLjDvgjjyuqI8Eyu+
1dlkOnISfyr13coBySouVPm3AxAIHsoQ8WpY2O/nVNFXKFP9C3sbrFAXgntyPCEg3OJvmzScKL/f
bMgdE4BVWwifD3d4Oc7QutyWfW16Ua/3/QS3E16a4D2jeU998t594vQjflVRO1pqkbdElIxTMoOO
VMdn4ZoZ8VGlUfjNpWNnrJ0v554TlvIn4dPJ5oJrFn/HvsIB1IrtucAiDON3bWbDWiGJJInDpMt5
Et1gnWFpbjl2UpA2RSuFxSRKfyUytC+/0kW8oukz3Tc/DOS6Z6cexQehWkzNpgHdK8nCbZVfxar9
sqWvS5/2U5Qgs0Cc3r5ngTiR3AM2WFPHZjSIynSmnVKrDBcanRr1EqpJeb/8IOQR0OjF3wIu9Yjj
GqSgcjGNkSlDxMO1SHO6ZZqox6ytgJ7EbCbr4UPicLqnzCYeFpae+i5LJQ8I5kgP8IHE4cqAFkIp
veJZDzfoIIUnpBLDji8koX7yBPVtPk5GdVQ+q3AW2X/fSqe9eaBE3OX3ftG3XFCUYwxN3bfm+m5A
uQx4wi3gIdDINlX/Syb6ZDW5uXDGNEayChsy7u+c5bJr47X2AdMBpdFju1gGy4phMNMiPGuvthQW
1bCZhwC5Kq667bDqkc5l+OT4U3vuwam/939pNQUcNdmE7VG1j1iZJ9mk7ivqfFcilt+xn9K+pfIX
7ZQXajG7mXW29rwUV1xdBcYnDfKTar6MVHuNl/16nucO/k0bGusPXopmBhGOdOFuEX91dBK2bWP3
HUbUCL7vrihtE1OMXMp+SKAEIPbCDqI8ldMVqoBMh8wYWK3WQ7rnX2jzzUM8Nxl8rFvF7PLVltQd
Swmu0lfDXAQ+La3Ju4HnuK5K7R0/hnZIsyOUP3sOgmS+AdO2f6fQEKcD6gteN5jCbUeLUmDJAgTz
n5U4bME8cQMOuUa8vPSY0DIYqTny46K7tDDRvXJMUt62HrcewO7BarIInhEUHAo1YRFEo/3cX9Wo
0w6891dvnrG+pYHvWnZo0W5Nl6dL5TX/zItaXfybTje/S+H/Y/6KPiLkSPDW58LFCC03+qDY4QAD
02BBcf7ClIhJt1Gs7Rcbm3JGMODtY7q14i7uSHzH/S+KcWxkK0P1c75QqLx3rT1JNevnBxqRIWT1
BiJbdnJa5GI9BMuchFCPCsHKAHeUQus4IjO2RACeIJD8cMc/HZ5y+lb4Fs/4ZDWBlq+pxpBl7Wbh
3V26luoYswaVDL0pFtqz5YCHEC9FPViD10flpBYwKM+PQ0U2sTYDBe15yv0yVQuARnBT2IA0AQS7
J6YP8wNui2k5jjhZuxlClJaxwbc0TOrCESeIO8TzomvSldP0fXuiy2/9rnpHe21uJ5bvF3MZhRJr
UI0Q5I511GpUu1nAebYy4x0Vrp8GQMvlL/SfNBIjKd5uCyqrhfrWqwXshGCqhqcrHX3HdrurxjJA
RNmG851Zv0BNWxb2jFnCShA9AVLjKr2lbvywaFIIm4wOibP2lxnK51ShqE3ukkkI/hOLxYcKeQLf
6QbL1I1GufeBf36WEKeRjWGpsOq/4YyFTrYXCgJ3u8SbRugd5HGLkYLnU9JfGGAquDUNDioQvY/F
xjOrYw461Ssyj46sHbhsVDwtwqjrUg9Bl58lm95Ahq+gLA06mnBTOApzuSd2FYAmmn3xmZ6yjlkf
eFWFrrHp44/y/qXAUGg+wPozrvA2kyFyVSazhjNzRj8FJchYUyMwVor02K0fv7XCLp7niP0w0KL5
lgbAR23uiiKiDrVlVoqPQRBF2MvdAQwC/EkjxYsCqKGge3TsJ7QtRZ9kVuBQM6j4MUuhV4YVLUey
DaGhaW4ybX4s9tCk6dQhaS0xvbpmMUzFMs3lkBBTNfsePVr5flreLsXVEiiWVjBkIAezvUtAjCJ1
GVpRjo0VYQTlupj+XZM5IP9l4Ia5ANOS9HBDdV54QvaSk2Kly0F75eAcDfWVQhwdeIEQEIqKt6dl
JGoGpohXr7qpfqP35o9Uq5waB+JS/N13IcprkJIq0V7KBylcmjHlm7Cnr0x/+a/CcMacwmndcQjq
A1nYSrw4s8IYMmmmLgHuaXpAqmXF5xINZeKLWp9UHodkGkxRCAooyfHZvwS7Sh639oukZDm7RZDs
xwv3XLyGr+BtH/eYd/TBiLTCHa9zY7aNr0yRLv33HKQJsxVIxVBImrr1RnWMahuvUrymFQDxZKzF
1gO6HT6UWHPwgcnF98PLE+YKLy8kE0uI5EbM1lq10lwnAJEsIa6b5ltSUx29aO2cyWTjG+rov3ap
98MXhL0svciwH696JL2fZLH6m4SPoXBqRETbqCN0ul7MftRECHR7GR0DbuQDSnAEvfrDaTwF1bZE
QqoiA9R/w+LH6ILgzS8T5Aiswg7gASweg97+CCk/DaIvO680mlFwFpEVbq7Ic++kHKGy6QKjm8gX
+K6CiBIo95GZh9/WXIBeRqSEfZ5y7BLMYhBl4Bx87J1CLGMfwHzB4x2TofDqmDLnuTBNZe2acF5z
A8biiYgJx7y2FXJajw4u8+oanMekweXkTyaoM0Jik6mcNgMBlwh4/OJJUdeNy71hqpTrdV2haN83
eG7anGtrFRqHlPsudie4TxHoiweSPmN/FPLsVQiQob6kGNbbK/5CELBypW9MgydZegMPI+vI+D/l
p2phk3VpSRmeIKJKiJTxHEANmM/no5bLCCP5Bbku8pFe44CkWxUdTHz/XuJaX5c7NP9+f8uR4Vhx
LIp3O6ieVAUf183epiCloagHe0WF9MtUhQ5PjgGPpsPdqaUGlonu/grSuCkGKqBs78X4GzdpEIPW
pC4JlMU34p348c3iiMYel0PLOWIkNcojcqqH9lLbbgbrdmVkdxIFPlH+NqBrBy0Uq2QbIn3mbzPI
2FyiXClKHPFparROj0i7r/b2Pk1z8Yrk4SuaY6Glo6lTmrWftJjdK7KIUgPi+uyV8qcDD3yGgczJ
wMzayjC4HBmE9wMw5XCLVjJGtKmouz9BjSjNiyvVICH2l82QijmH9dV4n15vQXAZmKORASKUKjQN
unqVIbaP88XkBF2eN+IMBhm7KXJiZ3H7u1lVJIH1SPHgC+7ylAYspXF+GmNO7Cpq20hd0gKPLUxE
k4VcmX8H7Mk/W8SXlQ2NhIWcoKJW5i2RSfR8VACnjnVYNKHFb3cEFHTcF/p3dFOgEo+4QWgojX7C
aGzh9Gc9bVEXaVKq/Xv8hkKUKFnO08K4XLItrZidQHeSZNDIA4wkuzo0OtXjsupJaK7rX3HK30IV
v2qm17taoLxYPPwqtT+R1GW4+x/z4vPFyjS7itlczFn4qGYt9QVpO/Jq3qwV7NQvqU4ItvsqTIF6
WPoX2UcLUuIRN9gTnkE0MRM6RIgZGCBv827d05qBgitfXe37qQqrCa23SBnjlmN9yaVXP7jv1C7i
toCdX2gfV8RqxvlF0FchgyW1T5S0bGw4SFWGnpDDuACzOFOkG4Zmr4Z7roBREPu09kx6vNvxevBT
cTYguuSiinAxe0XG5FQfv6a3XRZ40IZe1zgzHYIC6DToVtdTAxz2InFKJoqR7roW854ICH/sWQ3b
5MOAcKtflEuEJFbc1jA1rj+c9s5JzypgO2ICFy1ZKlo9WeCLjVtYO1U2P9o8O11iA3MDeKplsSi/
utNwuDTb48L/q/4qSQuQCcHihVU7tSzq3I29EZnvT96fEEK/vqVsakxwyZBkVf0TuO772/6rDlW8
YSMmk4vxAuyGtk3V0xXIHtYzSoxg0fc3x7ZjTnTW6sbKq4XvMhjSSAjkkx2uNRUqRCCVFWRtNPDE
O+ljldYbDaWa87KKaLPmO0Xp5UbGoSzga67EqChEeevLRecjMIUEivOratcHNY9GLzKJ7Z1VxZlg
w/zi+W052UKt6gf1Iugbr0hzAky8Fs44GYHeklcuuMsQ+F9BIPsv6zggZjNcsHAaKUu7JYHhQ21b
wjpkP0aXloubHLuVoQgCXBUqin5RK1yEF4R6XcXTSHWK8F2bOrwGM2JGHGVzNDu6Ij+ff0Mw28+w
6/FfW8SaxMlhg33nffSXwbMyv+J9D2eSlyDrQwJWW9nnjwBi9VeVBy621EqylfbMUrTp+lSeKdte
YAO/qDpm+m0aCi+cmbnBoVQrdJYz5LxqeInUsLRobDpFJs+PZhU5AyggtT2ao8fsMzKbU+3pM89F
GwyCm6DYXgJjrCLu0OtDdPo8S9uI/IChG3BOmfju88m+RgzlgoZIdUYwkIxjKRa+4K3WT/fkTVxB
1R7q3CzyqP2dF18l6UhFTxyQL3W4JZqlx2Q053HMIZ5pXOXaKZmG+a20psdBBVKAmfZ3HNYYfEWg
i6iVKxshp9Ozy3mptTlKApC3P0h+RDsnqjEPlCW6X9ClkufZ6zj/EPHrUWnOARHgKMCHxVwWCaHm
rLvjqIyMbTWr052y3+L6cKIUK/54xF9GRmuZRnFhT6l0Td51W3N4+u6ir//rj0x28eHrCYDFkCrS
gepBFnGTFufME8WnnQcUEjqspxebfc1w35Cx4uOasfNs/Le6NwTZmfItHmBaHzmzNzPqxmchweMX
YS9I7QARoTfz6rlEwSwXpPZDNb89C0hZkTz2+5TpD0Gwj3VjG/avVzmfkBtgKc2rXzfTux+b34/z
w+XKdjDzrDSKm53N+ME5HGlxFSd9xYIvIDxgAVmvyPVfY+JYmuDm51NfuJuAyYszKSzZo26w7B9w
GJByg5BGBj+z7NXVAyMjYYc3bqgEnQ4xtKABWw2lLkBvt8aGz2+AUz+UHWRVOTR8/ZIOk+XZ6+CT
Hykv+/9k93XSVg/EliIgm9wuvj3QWsjWR1yahc5QA8dznH45z9U6IqykpRqGa0RYfSFG9T6Vjmvh
w48wSl4hRKTu1v6an1O7NaH8UPW8kwtxdpd8sxMrzkWNGz4tzavuFACpCWpNDQO767LwjsoMaO1Q
hlGRYioWJF/80Kwyfj+k4baY8ZfFMu9waXfd+LCo+TyVHgZ8OrlAtoDXFAml+E0Cgb+YgFLsbDhd
uWqzrOXz5z6K8oI3aLGbtipTOpUZEWR+wMNmpQr2+w3Xqk3f/TKzsKzZtVagxDlCEm2F282FSIPP
lcOXmMoyvMGtJIuoNNy7UvZVh5LCHRHL4R/ngOuSe3sSY2G/ho/kTUmNtaTh3jjc1EKVMPgu9HuU
2py9xizEMDcd/JlN04G2A2fo/+5Ws+W7azGyEIValf1TDslVLhLb6Dtpi0r7YmzLx6vll2/LJVB1
xBDBO0kPXBxpGfS+DrzDKhYnGU7LoDmyx3UJEN2jxn+a4lYHXiSnmnboa5JkBMpbwN65YXaTcYMV
n0OL+ARaOHEKxlRSDJYLNP7m3y1hGUpU0EyVwOxCQ4xPMGKMocWYEHXfgn7IlvnyxYfIPyvKDhcQ
HBJ4eWMLUYCka0z5FKAIiSr/8RaxZk2Ix+AZ2hJXGwbkYqmSwx9y1W7fSdwI16qZQ1DFjIsQbIZC
00IU8UVXMMQq9R+ghUWV9V+etJCVsvzxvVBtwZ5WiXr4GUdslxXiQ5xgVvvqbxUUYn+K4fG+3C5S
jI5MeDtG0coNQ4tmhkzBLGLN8WaBQcthM8ViXkNurtc9O50hXVtl/61asm53AmAbIeIaAGdFiEM5
Ach0axamcY3ifqvvoAgFd4ATGExAY8abtP0A2pvg9fglGWg2KCdk1+forfTxKWg+6aMkEblQ4sNS
qreMZKqPORQUqIbmJMJGtP53Iij1f/QJ88XzLxgLmLdBKS/KSjxfwDXS/bmv4uG39ySBzzuNRDdC
fZ2E+4jqJHe86VahhhsHOalBn/z2VSauFM8QycyWKI5+NHEbxlVGa9YuRFj3pDDeGFGTFCmx11y2
Fs88zd+IRc7DpAUMynEH4RjW8cW8GXW2rTa4B9pcfU7ey5GQzCKU5AUOvPkwHYCAqu3CWD+/NC+Y
qiveu69EPfzd/ftxzzZYFxd23+GdpIW2P7SsIEEgshjcQXHkqwhOFLVr1ybIEDjPAgqIMPJJyVTz
NGaEHNfFVeF7ei9FwswfMcmHyxMQKEbasIKn5MtAHzZZnpb9N3XIlG/kknEPFF7/7n2eM/Put/XU
2XXyAHWmnnjRUMwL+XY3/eybQ/TwUwu37djxPuaco8SdbXn0cxcGEAAP/+AiMYfXmTCM1r6E5Wck
VI3iMbMwCNuqU2o95z1meFZ928lIvY0fOfVAolfYyx6aptXXc3fHHoDA+oFjLcaYhlPGeF2eyNPP
G1zs0EYZnkYuTrR+IeDd7eqFxR0W9rFQNQRspZiEue63dSPuogZiOYhTcEBNkjgtoiIcS1zWA4Uf
ZmAAFTYotX43yw1DwTyNZ4aq9L1B7ynvkilLtftxEYInG6MaRuv13ddEE1rVDpegeDDJarP1DHQ4
viHBWb2jUiWUj5/LpgpJ+L+8MHVrc2lFoCTgIhV43wEqkqVouaSgSNr+g2mPTXB9gyr2xcjBVx8L
mJEo20P3ZNT9RqrvMEp4Ig/8cwIGRtEd6Sb3NiynzL5z7W/GhqX6x0F527XlaXzLwwD5IiLzlJG4
lbs9QzoPU8Sp+5FxEg86woALIfI24EnebRJEJ6Ee1NG3UxgX5nv6axrz5EJv8VLYtSRG3gbvqov1
UBc575ptOQ+nkV9N9ZcKoYByFXTjCjzkUKaUiRNiNcA5BqDmA8RwUibvAY9wHD4RPlPzTpuvTuHv
ZqGs+09EKBwTrUwQf2LnOqViCUP29eNkSVURP6HHkAHuP1kh98KoksFdtbRv85h9zOL0kBkeMMmQ
iA0NipcfdivrFvgiyjlTdc5gW8dutxTMnp8QXmBiXrjOJioh4AdQR+bncdIo8ODIinRi8LyCdK6J
QkSW7dlbg9UX9ysdScifdrI7KDnQqMtjLXbYMlt04Ltq5OUmxTMcRZ/Llhi2aL7vmu6lPVT4bijg
5ZohbIfe+fjqBpTVFq+VugOBupN3TD0sP9pvIAF4U7pgh3qMlj3W6PApCHVM53aAD5shZOwve/U8
a5sI6QqT2aNjWsBK74qgrvOsvG9IqDxhUMf/OrXiJ1mBxDDr+eUGyT82PzEsKnrYTK3AlNxGtYNU
fUlgFBUY/uw0tk/qYU2AjzZ1Qdql1kpvYoOWFdjUfwIpxDPS0YLrbipjLQ6LfgPCTZbVFa4eJ841
7NuknfVptqTCUnC9cXbXccCLGaeudlH/LH+AedzqUtCs4RrvTsAueDpI6Cjn/5k/DitqvgqjArwP
JbvRVm+EVmvEbLSkhF6+B8oP3IuHgVfe1WSlWXpsyl2JzPM8DjXGNJ1veQGHXlUFztQwZ0Ed+Q9f
Pcva3z4xJcpCLFXnNQqI0tZ9k041ypu71NlYXFCfbL2Ec4/OMK2vvY4HggMWBO46bFNhnK/dUxa5
hv4ULDmiK/Q74eHEEnlvL0OwzrtOv4EQL1mJOhGYrntP0JzMvgowtATbGH+B4MJ2K7A1ENTD/xfG
lNBj9Za1+k3k2wvuExXubvRBRhesbrWBVuIHADLjACIqb5Ub+tZfZ33j4ZrmpHv8wjJmJqjpu2ow
qnbQA6eeX4eEUjxmuYZoz7XUzxBlq92KAdu33neWpKXXkCG8lzhEc5wjjEImWDXuSbB4J51fLSyT
tApNn31Ggs5oMLRRnY1TwRdqyagWBR171eJ9IMQdAeAjHVv1VuX9F1PyvOBKtokoHaZb4gCGjKUq
7vGELNpFS+aRviZTaBh9/o5kGg5dg2T4j+xq622oLRJxCKwPV0jMOhd1cWQOSK95bDVoBTrk9bak
KX+9ynmDxoPy5457pVba3APAUDcMkaR1vesgTWwm0NFQg//kmu11IvCUUbv6XrBXB9H9Wc7qVS4l
DgfY4DzndzuO2Ohvzx5aasgUEKm9/unh3QfT6JI+a+7JUaWn64iy5WCj/+UgMgaqL/eBz6RkD8a9
O/v1Lw0/26axYn857njDQF0yKcgOw6F59VKmn0ue28dtKwA9mkwpEx3ZLMAObAuT0VLFr+JA8liv
FcVY5tlHYFSFKu/OgZ9l1pjK9WrVrijG0PKqhNr7mTHAWRH21jOy44sqUP2FpXGwoRw0qNAV9v1j
pudTv7Ca4ei0xm7WDgijdNXD5+FYIu1nA7EhWr6mYyAfiAfn+l9s/StxCQ2iB97Rste4/roySGDT
fon5e8aHX1QD5nwIBz2GL4BsQH5i3l073Yz5fdLdyzvBRKR/fMq8G8c+TJkK/2I76jNdmriJciM1
POTfaHTWSWfhY6BIP6lnUV7DMpjj1blN331iN3gvzKUchaI2KcrxdlssF+8df7CtMhlXkm4tuKkG
6kNVY9JnYaSEhudzmP0q2EkF5De5DH0V75FauImPY7yJTjKmVNcP54h4GcGZY8DhMaWQJx5GJgnL
jnHAQOuqEccV+tLKT13v2YuqzNDRJVTmdYawtaT6GsjiVgT++tFWIPF/+ovKQPuKwW6Wugo/jCkk
lTCaohovf5U/2ek/CzOFptYMXvC3rcoT+ouo3pFLQY/c1JgK0y/vN6P1asprqlObCzBjVuan1QG+
I3o/K3SOJKidfhgcQd/hvrlQtqDEoxJPbTofkE2260u8cbB/LOvVRkSSERyj21lo1zadCznz34gA
l9/BDCYg2GtyEcNUJv0ebeVxy3BQS5N2PXbqrZO398MiGTrZ1vuLIztCTgZ9Qq9N7XVw8wz0nanK
VhqB8uqka5eimsqSZB8tXJPRl9BOiVfnwQr1s7eYX+4OZnFm27bvLOJ/+TuQRw6peefl4CmZLL6P
iADC2EjQM0zVd0Ybb6xLVLliBF/RJdbaZ/HNUa1WMroJSfmC/wmr8dhK26wYv45qx+za1HKFZDAZ
M2J4z5HPXP1csxs9JsG3oSdTMqI85sGJJ1vsypRYca/k/L0Tiu9GOMVJd7igDQAcrNgF3MURHLDq
gQLtqPHQQOX0qmMknPIy6MeRkYi4nYd5MlHj9XpEbWDtE73AYl9qIhPIutm+Ac5TLwOBeeR4us0F
T1r752pBUs91opynBiwhDaoqpS++03TRn/i5plzX+h/Es+Z0MiSbwVHEEplpGSvVFMdNE15jzBoo
7f1OEsjP1kJVgh4+VOtUjW992aDUSLG3k3rsyvi3cb3YtbRtO9/hpcH9Pw+pkGF4wO5XlUdr8Zo2
ZpQXzB2BhdvK2bcPjD0Trf4Iyra1FvdBsMD4OeVhdcixlovHlNWml0c3NHWArXTc+b4CdTJU0FkM
AW6GVNmcOfSTWo/ClMfwX8eDpBsjFOt4Ja0Wg0+9p6lvh2Wm2s3JqKny1ZiPurgSM4MGvp5lgqSb
1iGq9bJZWtplM+fTgjOMvGvfHm00BIc+21zkb5t8MN9nkdbPRyGm620QdehL1lfHDrgrViVIZLyg
/0rrurcpDB8KNWwwBjwnJK3WGkY8I7N2Ze+yxTX42hsImOHYiOMEMRZtWXj+lwXYd7dmQ/WO51F0
pUlzxisCga+Ngns1jpYbv0RpuzmsjTPsoSButjETI3Vw8oPr2Aw21XFpq2Rq8EhmMxD72BQgdGY6
7Yu2E9bl6nrAHXdQxw1NStvlWTVTAVMISdqn0b5wCypdWQ1ionrrz+Hl2Wqjo95oQ6dnbsEwC7CA
giQ37EHTuyldjpqFGnmkvHR0joOX8Jx3rF8jv9YFkAmYOLtyTlc84fdjpM5yto9RLn2z0FFw56oj
D0micKPZsjqLl1P3rxGn6RvEbVaGASpPku+6DJwzoL1PB0djwUJocagrQB/kmZGMcooUwJC5Nwzf
uaJmJJ6xYwCeGYHW3S7mW+Dz1g+WnoZO1brgQyIEpFQ7ZyK+SePcsQGuTiKiuzGmYG1FgewCkZLh
Fe6c4FrfIrqzu2fitgcehozP840HV9huka9OlvP6xgXhmYH9CtANMbC+YcK7rqrzv0hE+7DwuGhT
W9lN15Pen1C/iAYJAba1akBes9Ht1HQhp0RW9kosASwjiL4rqBgVrSf6Mn3J2O/C6TFuhiE8CcNa
+j8vlq0mPHu1oXAY34ySRHDjOM2SzxFdTPjeUJrYT1RWEr00UOFzbjsrJeMAOeF6Z91VRmAepeLy
MiqMlPJtfk/P7LN1j56NPk+pyrSnC3XxcpXbhsnB0oxxXIRGyea7yx/L1Teg7qNw5EOxiuTRdyze
91b9qutAXxGO554CBYB5Wp3wfh+SCzhBjb6ImLEvMJtEosqVHNroZrdmDd6uM/zfk3gyc+sEVDTF
DE8rWHO+W1znsIUMuQUOrAEI1C1Apv0fr3EMuaReSwjXx+bpr95z+yWiGJnGmmvuX5z7bvwdhlFM
0P7VE4uwZ9dLdMG1YtUxAX53rsDoj3qQRIlrBEqgCaDtzmnXxQjzcQNkeoC6IIW43qXVECqhJsnd
OSVxamlBPoya2Qz5f0LAovEEkHzGcT0xv2AYhdfeFgj/DaQzuYSYmvlDob15rVmvSwQcGbO2oZ+s
mSsffWIJDnGmASf8ZBh7+q1jpWSm1f4o+8THL+a6F1KlL2s/q3BspUcYOSJOctDK0gb6fi7Mhz6x
wfudZK2efgKjR6w8saZDhb7/MyOOFauIprmMMSx3r6t5Tw5F14WekfQCebBRt0KjuhNrMiNtbEFi
dCuFIplpy0uzJbyk0D404QIPM8Lo+oWXWrrsvO5R/M+oqfZAmZWIou43T8RpmIf7ZLPvw0VodJwi
32DEnvtMQoVIUSF2xsRRh/SWzTupnY4gtm5QmTF9TTrG44Xe2kLzYpuamw9C0l1je7cQ4aj0CSls
kP+XFSBECX6FBaSIBzPBK+Uvf/rYISSQh9yTy4tPv9cJZc+6dUROhY74RyRHbRXnfPIFXfFLKVxx
IOWAZZANWiJdEAx1fIFccavL5wgDngIHpGEiqXDK/4+jrxXUGFUM4RNpoovYny8cU0jucNKZO565
z8SCSUgtbrEGZvmqRcYp5ePbHiydZO0l+gz2GZdUkebqO1gaoWOCl6LDGjeRWbz/zuxCMLdDmoEl
fziKGUOb2VbSe3XRW+38fH2sjtF80hoLTcJuVvBcSEqUzrBwk7KCdUmH0yJ6H8N1e/8shFjNudyx
Oa9bfg2yL5eFGSNPD9BPPUJLoeaZo4VJGVG0C1L3+uR28lWEPDQiSWfea96BwEqYQ2ipKMGj1BL5
9jnFA5+zdR6LemMSCoOwOAn2zHvjsQbG4c6+k2YAQ8nEOMS1JzIKND5R5HzXp1QfuSukzq4X31Il
7wPiPjv3ho01YvppZWsZurbx0kNKl5Dqq6nPQgjjU8Z8x+XAgzjDu5WrV3y4xwzUIXgUSZgHhsuz
hku1nk1YJHY479U9OR8uuybIcrmDDFWfuZDChqj4dDA9g6CuhzaYx0NAsPgXq4vq5px0xbfaNCHz
cP/Rcl5QkvpbBn7VVlvLOwSoGRpqJpgSl6V7Klm+S6AeMDPtevILyQc8TT0166sslp86IJhDh6oW
MOBkAvPb+WMETresclp7Yj250ISBmr21XTi9z0dQi/1sqmWGJIMAhObPBz2+RQF6qzG4uFqd1kjQ
Vvt3HpoWX+QkMYx86+1d9c9aEtETiVmrzQIqlX3gSX+FWkhweuu4TCIIPF27J0RyUAP3QENVoClh
kCP2GDVMBFGxq96usDoygwj04DrXd5bOi82udOCLQOcpHJq8VRPblyRxy/hvmeoP1lEyn3hvLG8n
sxShdX0VzxKc/FdKGqA/8KvpRD6P/Dmj4rQI0HAAvnEl5YNxrfZ1/COK2gDjsOYfRz774D62fjoJ
HEdaDhYpqP9Uv4n/MO8Py+xcJt1smhsH9nkZx8QsYhYCPLjduF0rGpw++QpJqRVwt92EmNkoq6EK
9wKkXQAsmx8p8WzdhZ8T9sMR132LOw0Vimt0LCcb/OqyORc5N/aywCG6/6R3pbB3hRO1xvJmuAYs
eKO35F+ytlX7KFJVw/+0LH4PQlBxxCkc3QGIS5XWaVDfU3wg6o2SE91Fh2vQssdCYUZrggI3UX5u
2brVG/XUXYzjBnDcAnJSh4Rdhu38P7fjs1vUG/s++tI21cmSJbxEVpafG4TN4jQgBOI9N9U62WfL
Mslkg4P+nZA/0WRES5yML7nZwaPyG86BAIZ6XVE8HS0fKc/2uelVAMsMnItdcCWxJZKRaUOhXj2Z
GzXY2LHaksIMjQdOaBiqLNyPqIsSoMTCRKemKb0vW10K7LoB+12EsZn/dfNaAvsorPPZmia+mkyY
ZUDoGEd8NUOQxvJJB/RFNJTuseUBfnqTwpDReQPjtqZaXwQY+ELnb04dndLDKM0uE4S60owpQR1R
CgIQNXcEC+V3OJsXKrj8PQku8ZnAYF4MK556Jpq5wIYFgSAF4jXP2z1I57WH4SXs9owcDEo8/0Ik
ZriWSsP08igQoSSxJ1i2k0BQRoPBuQKbZFkqUtLfHGHmJXKLTBFcNp6Dh3xGu5LPcASm4R51KqpP
kUXu7L/k0dljPSb6WZ4D4kuNwoMV6UvlizblbFpHsn5LkD6K7qAzz3X/JxNjEwPcSunnv3B1ySju
wxH+x9DLyeNn0yj/FtI8L9dKq+ui69YAWfI/QQiFKW2G1/SIs3VDKuJCg+MJ5gjej9s5CuAAEB1C
N0OBKqJrTeuOcBOggiVwxOFsV+1H+Ew1cFPtIsr0UDmdF8TQZIrIoeLJRFSE7jNYBTKuQgJJlht6
htRdmMB/q+eNDbsHqGUq5848G8IvfqQWTQ5TZ3Ea+rgiKBnPAg48G/l80XFhjkUgCOTBw+5KJMqk
BJ2jtjlhKs92Gf/dvOdxNioVGOM30Nlch9X4kjI5/lJ50YcmN5LndDlgfsWzHDqzVrb2ggRxhstb
8K+Vj4mGqiUuNymLEgUZRQTNreYJTGH8LbdyryWSYSNh27ljX/JL8wMTCYkHQhP0PZo6U7znZwNF
rJ3BaXa9hn05GK2W9YxicbW848T/uUHbTgi/lqhURPRFPfAc8rsTw+efLucKMy8lVZTTr4iaW6ED
wUXp+jrnh9MNDTMD6rly26AatSf/jr7jPXRnP55m0b4GWSe0jUeMqIBDD9QI4jPCCMQC0D/kwT4A
sTyQSY60ht4stilyG0C+FRDRitDd6QBK0wEEnEnSQN19wJIpj+VY8d57kg91ug1DkfOR1DAT2GsI
tsMO5PIS9i6lgqSM7p2Sc3ea/fiykJoT4ppUHeX4IFtmixMDp2jHCmz6H3pbW2uXUlAH1UspcJmk
60T72ZynrYkcGitYwd7XfjR8q88XeNRYmyYs+7zsuC0Ygizp3r66CUdjBdfs9Fl6uiB2q/PmxVnN
vFJIEGoZ4oDGxmCG/869NjU6O3LTc0+mxu9w/zxNogTMah7Ie0SBkkK9T+FPkZiY4NaB5B+aT5BP
tG252yJixcNCj6/7fpo+49MnJDXGNYZrupMOao8yt/XCnMtJ93TX4LNZ+qd6c9zjQ5B7Ff0fduo1
2GZlK02KWxpS3A9D/pUAREtbKvem2oSrBLQh8XHlJra2mysW+cBMkXDcQvj4va3hvw59YEGHVrEB
XI2DpPEc7A7ptLqDSTgDFAN6kBmwRLk8zHc6ZzbsuSWhP25+OabWdbWDzOLvaS8L/ZdS8m+Kzr/0
OChTDwsc6SWGFkCRs4MmGaPs1p32WvVher/MbUK50wbiHExuCfIpjQa19w43j6xOUJ3NQbNblzFi
WJOkON//SXoh2yI=
`protect end_protected

