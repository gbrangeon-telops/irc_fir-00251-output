

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bdlZLEAewQqpv1o7OoBr4R377V8Hk5Fd8+q/Az6G9nxroFaOnD3V9+lWQZaiTQ+UR8tYlBixiDT3
2rrbvlUYqg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PNj5XhRRPylbuLUnq16m36512+Iu+tuxUNOB5vui/U9Vyxliy5LDYUjGyTrkosJ5RLmSfgYfmdaq
x3GXyG6MVOiZo15XiDmGz5Xa3WMM3TuUhfpzNItvR+cjVJcfSX1Vpo9/m4Gf2HbgWDY8/uge9Yz+
pdDWTg9IqOS1f9m0bhc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tfy6e9ewB1av8IAVBQg5F0wJVpezM47U5T38niEmKqoHE2EAQIsVtLXdGuC0EVCv8iR27vcg17Oa
mBfBXWB60tzPu8Q6DSJi1RmV8OgW+NgUvCiTMpLKqqsw6FnhMEK3lQVXfOtnfyh9msybPw9byzXC
dambJMmCpKtH2TBazWP4yb5ww1Nsz/1jL5i1zPiiJqwiUek+yJBHinlLsKOdmxiEOjEIxiuXMNyg
LMJzb839xkVhlMYTWXZYlSQVwwm/sLGnZ2Znntlf9sYBoE6D2vYri/PUGcfI5TqvvhrwG3MMHoTN
rPYZvU5TTqkZ0UHzprP9ZbAAvBMMlhHGjyKLgw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
enscaK3Um9KpWwQm1hA2XwO16XJLOAeYZ3URNnasJSAORmdXiuv1QgNvxstTqRmJdf6aiVcX+SBW
QAS4XOQmaHblVVCTrTFxq+i8/M/uWIiPlKdwfgcbq6W9GDVZEH2g71B4sNE7sbY88daOW+dsFMn8
evKdCCrOhrfApxD2w7E=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qn8TdDpu0TmAhfXr6OjdWoz6rfyBW7fFZKyqPOjjqWteCvm3OM0JlharuS1oWtO6vCpto2FAzG/S
BlRFnD+qM3W558gotDG5xKLXH54U8vJ9P7HSKDrDRZfcvgzYnDlLOZYqIhF3QcOp7QlIfdgIFJFF
P1RDJ8d43uSYKR66QV0gPXuT19+tneyhi0YpcaupqD9/Z/vQdGHiorXfqzI+zmAX5/7dF89mvr3v
Pvp32AibqOZJekU7QCnp4VkIAFQi2sNR2R1SirejbeSwa+gfCdYZC/MT0OFTfQjM0uxBSK/I4IyT
gWZgfuPijqASxDrsrURmKezc4hgCDujIExBWaQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21952)
`protect data_block
KEvMdTL86QdNUIvBxorxVf59oySAAbkCdoX0zkyQyun6YnIy7EQeNb2NZucEylJUGvQZKe1FHuAL
UKa8pszjk6BWjDquA60T9W+UDu0VtDmC3HO9Aui8+vOH5daZj9IS9zBPArQpUCxLTnfQbJOWAZCg
Smt1cJ26DfnFkPK7v3Zo9dEg12smGESwgH3LvC2LZpFl/CtuzFpvh3OsFOXy9hhiw0RKjwM3QmFP
O2qfm4bqXn0fMVjV9n8eJz/YssZpkeHq7teFULavBpMdipYRx0T1odsrMSJLqDF8wXFOLBq3Jdwe
Y9sGfm3SiNMHIuPedRhMnSvt/M0Vb7ujOIl8FdpgofgiiKh65JkyA+egz4qAuqlF3sA1PmJpJvOc
sb+p/t3f6IwYglJ00dv1v6TXNFwwGRm1FZwrEjciclp5hCm9qU650vEgtoEn1mo0dxOSsqPmsw+r
OVqbAxXTvQs1istU0uReeRt6+prbhPq91GNClDsffg+a8Ll2FMGgLF0NUs9E4Mzr9/MrcuoUPICA
6D72aqhVajDZE2SPTyQxPbfRWZt6gnYk4JhGsZos3bY74qc17yb5ARyQLq4fmHOZUokXxGoqo4w1
AZwzmvmxCLBWNs+UIWB8wyiDnPTU7Ax7SNf3XAPg0x9ZrSDsiwZOFqZyZasWmitnQiAh+f1rMrex
288Arj1uiIhBA5bC00r3Lckqp4Lj8TsXbikj7dG4qk9wap0s6VODhcr47hW/i2XE54/0WdqeTz7a
6LrWhzQjteQDEC0TLZqJwUoKKKfY5iN+pak3yLOVt8urQEFPNKwewZXpBmgJo0aOMokiFIUda9pn
RIQQvkYuKK5Pad3yaNnh2eEuoDqs9AYN+Zb3xCsejfFCP/d7LinnRS5/AnlBdSzuM4M+Dy0DEXae
gj4BPjF/TQDmy6J/91s4esFQlf5XJf95UnXvSVlhF0B1i+RppDcnMDNQ8zlpvMPlwgWA9bF1/36V
lMAStSIw2XsIDjOTgV2AU6VHpvMdkFr4/G+c/z5w5nIuiQB7ZJXpc7kXKIspL054tchkp//QPCda
/zmimP70vDgMv7oVqPI4hzV8zDngLGtulgL8QPM2kxYG3ngIhzjXy4lCgRk+rkKXQfO8kf6MqSvO
krbQmKMlWIpXX7k4gO8tIEYDcH5a1Cfj6gNj7zea8Jtjf2Cr2oui8kPkEH3lDXkx8hnt0gFCQtfW
k9dYltCYZ9+/CyyXlVeD968tKaYs8+PplxEwfzwxlEk2RVytWWIdkwBIG0tRgPs2BbbRKyb65ptW
qL+e2nK1xB8PCh0yduK8sFa7qPvAZNe7KOgoKuqVCOrqizGM9nFm6GKZc3u1/hLMiEv33uyMzv3i
7suq1GlpzmlGl/GBQ82uoDh3iBLB1yAolfO6yW9vNRW18MQkKF7snJxG5lhfD1qtqAXPq2/3dTPk
1t/K/1tMcdKymotjf0kCCSBQhwCygmQ9Jb7tPpYet6/1mwqwVrLUal0iNabjZxGKfRm5jsTh/AQX
93Gn19PBy6XDroT9ZGyeVm6u8H/kcI1qbPLoqBa+BPUhxIkfANy3cuV7SY8t7/vqePPajnHj1I/l
tGo29hILUQnCv3fLj/IF4z29eke0mHiDogd44FWqWKcABA4A3P6kM1FqOdRa1xRx0BASVP2ONigq
z8skWo/f5xR9AfLG+zdTtJjzQxQOqQE7uy4i54fru6LLmBsqrDgbBQHtUkRvgt2P/xczPSAslbe4
VWJCVMaMbGRkpvF7+/O8u/m8GipjWC6kbqYYIOigI6VwIRsvb32UbR5KPXp2z50CnQ2Wc7AaEzDy
PgZ8nU3mtOpTZ4Xpc/vwSbKNqEVPrcYDnfoB/0SxFmik+Y8TSpNzMXulP4St9RQsULi91w4sd66L
kYcrUKmbp3RSGFPCfu36xgnwhQ/3pICsg4w5jXBlqXOItD++8sjx3Uf7h8BmubusfBbTBTXR8/lI
iBpqqpafKDyEKzoo5YNpyP6Uq2wWQasRnPchmiyF6Qty+giDSoyhfzIiawFM0Tu3u/8p+yLAuWS6
2qeATlNri9uRA1HlWPvXcOqrJmgh59s9E/x1bN3+JcSoSxDYK23iOwqR0uQ9TDo8QNWYt42OhJTp
wYhRd7S3SoAMYKRDDzHo8KVQRV2Qia1mBZhO9GwYWa5TiZBFXr8s2cU7TzMGQToRRCGW5AdVaf6h
Q301LvzTL0fbo17WM9/WE7pRpDi/2drHV5ZDqblEyRSyIf2cTyGb1giELQNWkX3miFFhhmL7e8cd
rIui6Gi9IMu+Bwzkp7Ksk5e4wfqRYjWq9+7iiP1HcEEofrXM8PDEZ4tRaTAqmRgmlOD/ww10MWvm
8RHOzpwTPiP+qr9rKw7+txLAqWKcDBN0CnWHU0TitdIYytdmybLEfhzsRRJ6xNTP75OGDvqKPp2u
hWaQfae7WQCHG3spRWygBAqkqd1133okCGc7ljTAy333zSAzud+/xOjWXoqZx/xGpvpSMcRd2WUU
3h/5aLeAlkjuK/1KjPEBKQo7HF8IpRCNvou4Us3VGijmUGHq94EuWJ2oNg033svajKKZPfKKtc6L
7TMi5xeTCBrmoPu5FjBBSOnh52TUx1f3vZ5WULwX/4MAJGqNxu7+DSM/iORWnOZoVZc3n/jx7+iw
hdsLU75Yx8QU28QOVytKeBxl5nGMUFHUgGexucURL850zIlfKoIY30nSRjZezAq237LHdZui/jxq
GCdtsx1zdfM6y6yHSlEZmSvyY1JE1rur/e5I80iLf4BVExuzEOtB94dPBSmXyJwPNaqRLJx0yusQ
7sq6GZ1K71r8eYUOSnUISyVpah4v9OaPrLGYH9Ix0f7puyT/UquZBi++cw5JiHsoDhTDyPHv9hcs
NrS+o4DWuEBj2tjz7bl/fH4O5tK9AognVprmNvJYlxzPOXFwZWiT79NEQoy+ff6Ej4TKyTUnYu8n
cdRmoN428BMCPVFZmQ4Byt1C6ijXik4eYXCD5aqvojTRcucLeQJeH8ImApGBCNHR/AFXUq5uoFIh
yf0I79ozEC+B/3vTwkjTIvenHZ4eSlSvQVQDD5NkV29DOW9PiLNhWRMCqoorAFqZw3QebQJuGEG9
CnjP6Y1b+6MUpjV/PBvmGxr2AjrA3mfYY6UC3FKN6vz3h9z4BsL6AEsDgZFBVrZnsPbLZaMGSlEf
CIZbme2k9D11lQHtLz0TqHobgYidXDO1PO2sTgevRP6OmkrUOZi8ECZq6MxE2fPvT7wALGV35CNM
vSarapYVIgl2XSERiKMdzfmxbWEwAxs98qWlcBmOcstZTbUP9J7zywijQr+/GxpYX1GPq4X7jW7i
gngkbjV8tqkp9FTMd28xdecxXfzThWvCsrBiYK6pmj3OB0IrXl8DM6ymzvLoh2tsh9G+8JSgkP2V
xG8X6fe7jevmTFsFNuadYuOQK8DaeSMyBqj08ee9bg+hhw2I29VHTTANJbudjda5hKECsBNKefWS
N0Tw17UWg7QweUkmP8aEEDEjmUxR2kpLunNbqrYvkQdJxqAO6syORVZvS7z/8yzFU0H2EASCVftc
X8naMPN9iw25JJVkPTh/S1c/2xi9WqbZ9nUdQK5MRvhZ6XKWnNlqKrBOpxSluBt+TxMVARgcZnzI
0JWyRC0MYhtdvcr4zhItMl2pBXRqJe1w2Cv/4jeHsMIiAWipWZZzbB4KQ6pcU2LsCqD/V8CL154X
t9wXvMqyXnNAlVOtNfWQL7dyaZDW0mB3reI6pav/N4OfkG7Lp2FxQVr0XE2yg1GhU4yCZxTTcjan
cZbZQH+dEhGsYSaJblcVh1pIJcciJrPLue2LEtD3E2Tcqyv7NhNkUD73CHzq9f9qatcelcRoYu8q
UztlJ0GZvob5JSX8q0sCUTJ/Te2Nwj/Oc1TzhJ5OOYxfjgwnONb+bxMLPhZvYGJuf83wIH9WPyAV
sJp+AXktzRbIBUE6EiLp0D6Pn2hH5mxF1uIotUfmBXXGRrS0I1Gq/F5MbcRodX5WMQfx/RLru3TD
/oykLH+pzfRsPBGb+s54s9TdcZsUP5pEWm5EhvcTb7XoNAMxyP46Bks4WfwSvy3aYwFh5heF2FiQ
V64Jm+j/rHTBfjlXGyezX9pSxucg7k5b1R5RdzTHd3z8ngAnu1Zk3+jeSChh7BeOLpxYG29TNW5a
J0HAeUWW0rWN+9tWk8YWsz9RHUgzg9rhOQfXT+rvlr7goVpYaKSsy3KV4XFMYLBbUwk+Gyh3uUP1
x7a7MGWsG9w05BVN+IfXgidg5ncMkMOoFhqLv6ck68R4oxTplJAoRP3eKeevn2cuZX0sEZbIbjNB
LlwmsgwJUdn/YSVFQBqU9fRZ9Hfrh4meyIXOGopc3XIaBNpsHS6vmZOvjvOVxxcxmMw8QXdGRP2K
Hsr4Icu9wEPTPEBATwA5cPhQ+xCwxHHV0rtrpO//4JEZ7ria6YrdpA8ET/6FVTc8LTy/aVuCH2gO
ONx90QOJUFmTFmNaNGx2F2laFuWBNqTZEgZm75mz02z85EcDb1hLkJpcm862q2W25KdSuaw/WZ/F
wkZv86JjHX30tJMJtDb0AEUkuXmNUjDEASOpVjQ8G/NX8VHlDIqozIBLnjIhcoYXpBRTdywpXW9I
yaot8LCL84R8FSTbdlFjDngQ8aGy2oHmt3/58PhwR+6uOQxa7ky+PFAuwsKOTgkhAHd0TK93I2kR
GLJJsovK+fFtOiRHLb93oRPW65o5ZHnmGsxkNU4z4bJfrHRJ7LEB12hiqGAppayrmyrXhdepiYYO
JtRO0AvPf5VQ65BgQUdZUb2A1jYkESS+QbGAz/9g/gF1LcYKRlejX7mxdXYGNGcmiBiKcTxXWtkb
keZ7j/XyJfeiNPR3P9PSdp9kQo4ueHyW16FYWZM6niiQz7SdXanKA58C/wokl+BqeHbFxEgBp6w8
ol50dJ7xOrqwZ4Sa5R6p2ODrnStH7RbTu1bD+Rq7YwbCMEynL0m5YwsR4Uyq7PoQ62kYueRHbklH
wU3DYDLARplLel3nSftYq8nquO61+ASyDP1xRKBqOa7uCydSwYbKh54DXMrzJvDf8epBesVVbyEP
60Rh4U59bMDtIV9gZD6HJpKqUNDyEkQJRYUukDS2xEZoF5ztju4p7aGTl6H7VwGosk78eCDpfMgj
8F7aivFc/yf5HALS8ANS3d3A6vYoNQiplv9MsO4iXdaUTlBY6VN9LikjlZpJdPuSa187KjUR3o0C
rQpDMF6DcQ51HF7tAsE3ihHfu+6muz3Qn3IBIKSA3vVAXFg8WSZbg+nPiLaRzPjadt2+EpRWXTJc
kf+XVghtp+UmV8VdnL5+l3RseOg8o9WOWGGYvGn/ESSWMXXBgSoTzYlHhvYeiIZl0GswOiGnUCJj
wssdQ4KSXnq9uTZNucqLI9dqxd1tln9mB2+TKHnIrCyJsK0G5XBkLtT99yacw/643SS2VuirNlns
dFQcTk9zagRVBM0sfMfEZXS9EprGXFYCfK+s0mgbqTNpGV7HXwt/nbLg6sGs6w0tc1BuXlGCMPqU
Hrfw8fp+wV07xx1il0UNiqOCO+DGu2EyosQf9JL18uPpXTdwB1KUTRhlMtwXuS0+BrK110dYmvBK
AwyUY3b3FEvgZVbujaXGIaz1VI0aKH1Ho2mCGAxQ5LG3aCuLizd32uCAuqu07j2kD2FJisoibLt1
0KMsoTOWib1/ZVM+daB3GqAUrrwijWgP35n0H42cyiU0MXmKeC+er7+BkZ3e5yxf9PFNMcoYVl2x
v0fyrZe62P81EVf9gfry8/8Cep0vKxzvi1RD8IiPklz13XDATpDD23ra9fTFuepi5NUr7s5+5nJm
KqUwGHAAbf0AA7jlSbQW2kvK9sijirBdY7E+CDqMOcOvHos0jXWSNzjtQ06rzPIqzVjj5sjaSXyI
cvYtv9RC3tS8JYCiuuabKpcvyKl5xVJCg1LaHhuOsz6PaNCXSXQ64I/B87VVxXmUodqap3tBMhW5
QRJ+RYl+yHQ5krOj5PMFNjV5rFFSLfWT1NLEEYbJe8INmzVsO9pUhq/yp8ajQCh8+eY7DQY2Jn+2
ILXdiVfrvoADV5QlG1zdJQnWUJlpIhOigZTma7LmVElC+RcyOKBhEQ77gmFsSmcogz0at+pnYffI
I8kAVc4UzF2RpOwst3BtPvnsShkaxxkJoCMPz330gz3JAfiFPp++9Vee/GJa7NvHuIfLE6gI6Lhx
apbszw7v/ncQZDWf8M5k67tNUByXuICQzsmjbMMQhJgdJkmjy32NZeNqx5iGC3jmxisfUJf68np/
IbvntCmgY5O/z6wHmax6eWwseLzoC5L+wbHjh/llDhrZXKhMoDsrYH0Nln+ZEDEh4zCvC78ZPvk8
Qu2qcegzqX6+9MgnZ6sRcS74+MeXqHX/nbyB+dK3wojGdH2dIdh+3wo9dGMBf2YOqqD4QQT5tQ5t
9WEU8b4gd3iLstzM2ZXX/2kw2JYoPAezBONVVuYJXzOT0CHq0FrVp6VyN7UQEYCI6UgiuUaYeTgM
iWwdLVcfonMqx8Nts7Lg1v7s8+41Vohjbef8m7Ap0d+4LaB8xKTBv4pQgD5f8kV6GFZ1wFpQTzt0
ilvRj9O209IhUHKu8ULd/v8DQkreyOBVqhwr9BiUJukRc5e1LjItABS3aJ4kAkIMVuchOtFjgIhl
uvVeGSnHWchxCsgI74w0dxHABKUaALJ+PeWpFjTTbDjPB8LM19djpcoCC0iZcgaqRoTbd4H5x7zd
xej5IJD7DwlxJsLE/j9hsdoFeI7BVUE6XlmdPnV16SFzrAevyEmAbVDfXnKy/ddlQl3GLqvtFucS
CI7ZdLlyyME3WnA7HJgMYsbQooODYysf/wKLk+Rke3HTdHhD47xrdTxMStpOa0XWtAd39ePFBWbh
1vpY9peZOZMcJugU18pWJxmv0ou5gTxMyh1SiR3ZGzoHTrpAEJPJt717RkqCtTKgxG2+Enj8jjxY
CAQeqIaabWk+SeGu1+0xKq2f3otAX0nFiJtqh4sAGtF8OSkRlXRack+AAvVACM2NtFMtqDyleyft
Om8+LP73g0zBJXToCXB4KkaparPVnmbbqb+m15q46l5DoEqRHGrOdroKeOdqQFdQUSeZR+8iPq3h
Y6S9aLkEGMFkMbhVf3bbDJhkmD6W8Z5dfRelEYhWyr/T0RRy+Bq2GKJfBtWvOI7LjhZ7+mnLnDF1
SSmb0OLHpCCZTCflVvaoo/o7/K+GCPAm0pvLJWr0z/SJQY2LBzfnjXEZdTwlFiHwKSG62lM08S4Y
zzDk9YfQKg1cOc8yYNq2PgFPBf/TbpTVHa3X9Y/P5SC83e6FUHbYLEbtlmvmc8CGALrxl/0Vhw3v
xy1USqMLUgMziAacECNwx+KxMQj2yj/LLhrnoYoiLF80G61zs7U/RDU/Eijd6w8jGZ/Vr+vTQt3y
GkA3PrGy8C38h+PBCmjtbDPPPmQBvnwM4oYdfUd9x/p2AYedOszjouoK1dTOd98/xE4mblobkgrT
oU77SJJ9QJmeA4fqe7eKB534RPSacwfg6Z16Y8+ZsW3nuGyDkR8Nq7hyt4cnx3kj3ZE7x09i4t9Y
Ni7MIPndvYAgfsAVZF3Im9Ml71oGMGPSPJKQhgzZwLTcWw9DbrpFhiLYUPEHwimiCYRzcMAREt6H
o3BIrmtNxBHrPBx2A07otvIMCttxH9HqaG41RjtnlhnCP9O6oEpMJTU5mX/vU6jLz3tF8XSvejtV
fQg8+RsgOZ5pReEJ5YwVzuted0jaClUhhgXQ1eVItuzMXJm/+Cvs6WNDtCsOC/H84snn/uT9MOiK
LFoSX43mxefHusdeZo5Ku2GhEEsHZhUJsRklK7HkuBvp+IAWCZ2gjZMIVGt32Phx/EGo+Uik0TkY
hB82xuLCkGoRbjs3LhJR/34+43t6W8ykCgU0h2LPQY/73OemkB8+3WTuABttkjWnNfuS1fhnBq8/
vD9J51BlOeGSpNBNZYibPDMobTba4gWnl701DQwl3mfu1oXO71SFHaeMTXng1JrXh1wi9ta/ocda
L5sFmit54wYqwoPg5CVrYCBZ1p5+HPVpnad+jgVILOQierMvPYXw75OOsweo4nddvNRd9E8KX1Qy
cHn0g2QSvbaukOYMJzsWnVlAMcrvEikm8V7lks8vxufOjpgfGUeE1JfQJhlgC/ze0+knTPwE+9N6
ZOIecu+E82wbrq2pYQE1IO0Fdi4EWzAI1TpFtX9YG6YFwK8frXRpH61TdQ6uuMAGmhnYfHti5+Wn
y+hPC6t2iOesKIfc6L30yoWAwctj1cZ0ymhNDH8k4X+4aFfiQw3sNKebyIvoXiEalLY3NIB59iYq
iC20ED1vG+suVyU0nRDFoCUduvoYLCBkdF7GEopfWYxKJIYPAecQgET/KUadBgQhv9wd+njDBdbZ
7m8L5BInHXXgS93LsShSTkVb6CwhAMG/UXmlywsdMymcIHLHwB8QG4NaImq/DR/QIUAIZC7g5h1S
Q3PtTUTNjesdsqH2HInufD9JjTjfPETCzUXv4CPux3KZPQFVVVwsDLeNO48kypHzaNzGDenEYNXR
9/QyO7qGtmkqAip5q3RxHBKC4Nn5sV4TZhlrZ829t9aYhAejgkD/IxlePxxNQjLfLRNE7WWMBdYz
dQ95v2yx539rEqK/pBWCo/F4wHFWSWKzihkrH01MOKS2u15tUTwdcpD0osa5tNT9NRDqhvOHJKnq
UeFz65aRRzqXMi0aSDKXNadklQCLQI2IGwgpRp274pVsxj+FkSM9IScVhANppF5buE/ni/gX7SXm
v6HZwqtYQdiFPSL+xGjCG4VkHsk1qIdmMO11KbY5qK9I6FA+Rt6WzLdmeTAg41CxjouWNziElbxD
WksIA2NzpJsqUhaDPfQIxLTP4pt4h/N2F1AbqKmgHo8O9WqI7frZV2PhFUdngwSR1Bt0R3R51OLX
ZxJ5BKDMBh4F7sKVwINNts9oOT7dQQPy29dCbCxLBmuzuwNQdSow8sz+q5P8oeUiWnMWfq32gBQg
M65nceK9Q90dQAzciBLn7O5a36tbG4wjk+YRaV84E6xxSqRldBD+AMp1KS/uWlHA+2Ja2+1s35mq
xH9HRIuuvKZ+VZ3+wDe9czmXgxJIv7vd4IISj9UIAj9giLIXDtcAGufQK86t0NAq9vpOTp69xBzu
TnkCFhDmIbt2u/L9wyiLYRtNJOsDrb6cHbrUzO7NBZEIKjl9/9IyHYwh9IxO3NpB6lqtDxvUEN+C
n4eF8BQur0CFiGLXpSWst51tOrPsC3HqEQDKSd1uFPk76Fmop7Hy3zd8oCzPLl79W1eHGWwXsSeb
hSUZoDa8jpggetQTcllxmwC3avvlWH6Sf7bhwXed//+EKju3bn10jb3rzyLogl80jAbP6ICZpL8y
1ICk4cuIhdTdVhYSgwfT91uhgxndml3T1+4EHhSBZZSg2sKy6EMu8rdx9MLzfgG9POz1qjdoNw7t
2mElmuZAQEsc7F6LmC9x7cr0p42RADZBnRlvVCIHGrnfrgaQehpdFYeZtGz6/rqADOhphCRJk5ww
nBvTQfeinIl7blzFrjcoyf7zareb6WP9lWdZQWRqbGhvdPXotZfepgFgStzZw7iG17kDDyXiVKif
Fe9lgpOHpx97cbLR6yrMLXe+ljMn42KjhmqQsLyYrUbBgCZtH7J/XqQoMlBB6bS/++Ggsyf8t4//
83IV52BGZJM+eJkfzXHGxcCy1u7HjE03ZKC6yXG2TGj7v2abi3mN/xga0+RtEF+aUTwnDnsfSo6Y
xiygcgc4N+Os2Y/8lAfO3ZgNCwCZlQUPy7hV0RQ7qc0Q24Q5GzWmRIZV77G3qsDeHXxaz+UJgibu
Bl50mNcEUUxWXZrVy7F5TELRBczS4vUFZUHHA56aogDBudz93Ro3e+QkMiTvddjtRZwttdPY9szx
gt6ssc7f3aeWPCEZMCXYf4UyuCSR5Q7nqx5K31qctnYPz+mh0aVKfQa0ug1jF1FpGQNnIYPbPh2e
AJH7BmYDqkfGX1OwBHxsqg1YrQ4TLrUZ49vmwdJUlxJS2UXPZ1voaxZvdGs4SRYPc3Vhhv+pJJsH
4Kz/aBC/H8l3a1BfuEc4IU0tQO0L6kEafRaIR02UT6giQz9WXHsNlnZijdWBgG9du8hIJ/CQ9Yv8
CX1wKmiBR5AIN0+shlWcg2lNfG4rYteOVEMj0of2syMI8LKadftg8x9sLmjFgI39XZGxdgxNtYtg
nDXriHH+QjGWhv08C9u/dIz5GC03atWtceCK/cgW48ZsX2rTi1qvzjHNeG3nkv66+u5JTAXLlkWa
x2IfJPv2iBRSDlCp0oExJxc5dGjxyAt4B+0QDAzo4DrWVOydG/yFQatJQK5ZFTfyDKdzHh2v81uZ
KOMsorp4gyPfdaXVQaaTcamWGHReAEuGadb67FIcqlv2HZneqp0PW4YzjVLgg6G7Nn5a7NGiIM5t
bdb7NgwdjfUOb5RtwAP14ROC4XPThGXyqA6sDJS1B7AJ6wqcgp8PVFeekWLeaRCl6YOO4REIbdy6
sJ1NENDoRgUg61leR7EiuPzQ/62nREFzYz8NIImRkfXcYS2bp5ZkJRlnR7blp/FfZj0rupKFD1hH
/2b1O4n3tgQjnoT9SgdbnRtuRi3K0IaHixgjDFbGw9ZESQ8PKiqh9gsxqXHezY2Uqtc9IY1WkGdZ
F2x8uvxni/VwLMTRIOfNAjh05SII+VZaKdz+rh3XYT3GHa1bz8IH9IYrZ52Gn6L63D5EVQm59IvG
XH00qV6l1YIuWB11mpkpuBJRHmmhUlI3ZqQnVPAEvmMM2IaP4A2vaysPZakPcphwrORo+b8LczBQ
5pD7ifmqcrALkHtjYpC+TM73taqUcpfffPmrGNxJn/KG9uJ+4cl5uRjLuqkBE84hod8X3t3s920p
9RpspdpjXDInlcn6likKNOmq7g0Fvidepn3es7mNfkBB/kB7BjNhpHwHSzgJ2MCIfnHlsPoay8ic
ZpKkyY6OkGnB7u1qyriMkcKhDE4Givin4tq99OHBtT2BiixgeuyXngjtjrkZC2nHDfeRlFtiZ19h
loRgD56I0XgAJCaFGoTkAKbimtNHHM+/zsKJeO2G5zQT+c1uKW0kcMZ6u7FMTB9AsExp/ZZgKfAf
0kdDCqW1kRvqcOLnKO4pzDHIIqxMaHDJEh641aXhPc6xsmUUUbNeuzBu1dmQd9p0Z+oMZRTErvTj
kcUzmi5udLuKBwWwHjYKpK4GKaOEBMEG1aFNWezr7xPrQxKUHePyGYnCHp6HyY4i+3d4QkpGUwjH
yAAIXpE65kLV7mw3FcjJUxEHUZb+dGjsOoIy+5HiPwAaRJH4e8S7gVIi3MFiWiMxVOpkjIdopUfi
eKDkt1oxAll2lG7vPpl7OrJ0+dUNcBELUTMwcONp4JQrMK2VjgRdthTCQSXkSxV5zu1vC0l2CYFI
Op18ehPBF9BlE1Zx4e+O3pCCDbMagUn6dRD3102t+wVq25yfPyreTc9nC9taIBIQZxkERcxIYrji
G37bkiuXjb2/NLEPige8Ch3F4axu8nDe8sT0H7cd9L4GzvjVmFmGwrhIuSKeO78ngvxt7krBIaKs
jW3Y0iac7VWkt99TLhkKeaz3laEhTlgZYSA51e059JMQPegLcZsgYnSuTdUwnt5CaI//8HpFg5Yd
X93qxhKIIf6KfgioL5YXxe4uD5tn9NWDcRf0vcurreWZ+K9QNlpGK1HfBzX2Xx1Z6Kb55H9mFrdP
gpfC2MzT9HYN820SjjInlp0OTFMb9/Voq/KeXyhDPDLl+HFOsm+gGselT6PzDhbeC1XosIs5EfHS
VypQZ2iURw/BAsKNnDugTMx8/jS/HAks1eMtizlyoEWo7NU+VUB0s/kSnMEYhdCWzuKvXaW+g5Ym
KSbZ3TCIyd9JC5AuUxvTV4ZysLhSADEJZrPqg5iWH+e1AenNpcneYiM/FQq2xDou4K17l04MuVBh
4KgwvvrmqqX2GSNapgtar4yMZwYpDzqo0iYRczyl4n+rMm1m9CuXIp1aYvz9fugFwDz9o/5PDt1f
4AHtoPtCwEYBKR4hclNgzf7G18wGq8MttAzBlXWSTT0zssNIHPNixpGCeMfOmJoODT/0DVXCxBwH
A3FLQhpJLLFAb/n4SahmsqhNKTvynJU2SQquATdOMuyWipkdxpIYWtJ/vZga+ycKcltPX4928ygI
2KjHBEVK9rn+lu12ol/ZMNuTKz9VYTUcowq+M4Cvxxz4PMFQ8tynCmxamVwJUM8LrVrS4PMABpuQ
w8ZpsDlpadTsp3F35Nj/VW4HpbAwkA17xVq+zQ76Ls+LPAuSQmhhVvcg79go5N4WaiFXjMkTeeKK
o62St5dyLzDFXX5Ihx+onH+q8suRhk3L07G7bUv9KB06izo0PqXe9pLrup75fihPp8mgbCOym2nj
B0i+tmcUccU0SkGvS+oSIvmGugojy6CdzMY4aeqEwety/N9CReoxx5oyzNWEVC2g/VoQec3dn0u0
rQ90liZC7bHDfFaPUcLi//M6pK5Ef+dN/6EPQdHRRHHVS5LUnPEtFbkzsFx/1iZ3d2kTlk50pCs5
m6M6WKe7X8WUvtFExhxt3KAXyqTp7NRl/AL3ULGkcO6Zp9w01fWs0gzX5UutbrjMVJig670n0teZ
TMZiwWjUtoGgkFswXn8YQBiCyJXDpSx6AMKo5P8clqBnYhqSrsWfprJicUSJzCNLZ9Lm4ATT0UZA
x60HgzGINAEx2UrIKZUShAvYPIe/Wr52yfjI57NIQpcoLkCGWKXpg0zBFEJTBiue5DxsJgV3hmcQ
vLdP2kBn4z6aDFb36ATo0P9Pju3+WZtdYCZF5K5CLORwLwbNoMMBkRwE+Lb3FebgeA5mP4ssuBYP
NY2UtBEtzdxLhg+akSpNSVSCLmoFllFXjUj3tIjmTq3bID+z6ARRKsiup1A7NCzUCplPRLdqTdYk
fCp2aLusUEPaBGhTuWy6/LRFmc/a0rXEjoSWks4vIRrbI57EKwM2ldYLByv7MxETDfLwuTwdoOjB
Ut97vuJ9Gb8u4Tj8Qa+u3xW6dLtdUEZwY2Grm0O2RKuLc2WCS/0RcwfZpclbf+zN6OpVjEOLwkJI
XTt+g2orvbCU306OwLq1oajAUfcpKCB0PQMVVEfrKK+qQifEgzIkdR0BvoRN/7wDeW4l/xgqMP6i
yYZn8B8/qorWhwnEp/YauD9g+vmwP0kcZANWUzOABZhvwVJrOVOMhKcnKaCiQH356YbRkvY3F0uY
7ZKsP39l/QcTrHqjXH/etHbMeh8eVt2S3LVyKN5t7Pfy7Xrm3VwHibz+ZZvFYYKiXuyZmwENxTjW
5KzIAknD0zI+jSKZ20zRK6KlufKoKREJuhAkZXFcZOuHhHp3Gh+Z12uNaPpRkFRmbuAFTSZ8RIRI
v4vN7qWnnOADj+Rn+hODCcC7e0p3ClP5EJuRGQKu9vs+GfKAeAl/gjO+5fTPVysZxLwzMuhs0HsL
j9LvgVTFtjTeWh+O3KKI47HNo2juy/FEMxet3wL4H6UMwKjRaI1xcAi79KWtg6v1swIp1YSUM8gA
pagBF5rgca6SyzLWVkLQkGkzU+/Plf9Q4SD3PuwTsnyOhIXuFxIeEzISZojudge7DwN2XjfI/7SW
DS/I2ed1C/0Us7/ZdWAm8BDRBCg6RRXcy1oarTezEENOf30WX3eurVYhv/OVfHIvYyjlkcz0KgkZ
Z5zcNwiF31RGuQMAg08rBqaDg/b6mAz2MPLUZTIxTGBI0gYZFZSfJQHk5Y+k7d6KMQk3LoOkHQ71
72y5fGP7hyZKjM/fA76X2LvI/elvFI823TBgAVw3fA5mPNXuaxI2YT3ZeHmJNlqiWluLM4+w6kVe
7Lq0Xq+zu9MHkW3AtefGT2YK9d6WHQNvqAed0ovMn6pjK1B7hW3vIBKahXzP0Gz1aHvoknNVEO0x
CBv/9dY+2PK2IGCtFBAV92UOiGs6ZL1kN5Ycsla2r/fkeOYwRTs3gUEPM+cEtvbdDimn8GOV0nER
nlmY2B1jdtVQaT8RlPjjBbYlzX+9zc55lfhN9/GCIOlF+iJ3yE6htnRy8IJCv3rLUMWl/4vcd68h
w8WGI1MuaYTqdBRujdugmzZEBCBB3AYabWZfoDev6ubYBW2vBqTsjI0781xwrRoxhpOqgtR6zxru
9Rp+xxP8mZAJqGe4dXEwnAIURqlFC25uyyvYsy7m9F6d1wcXS2d90NJlRt259vAApx4vpyXzS/xb
rGr9zrYHL/T0ziTzXKXiC2nIaAR2mK9jDvh1jVc+gIGVIyHP4NRFYAH0L5+PlYbOLphYgXt3Qdtl
yhs7qbQfbuWzIQwrzLFVRgVC38+KKCshPI1YRWAUVjkzX5mpHazje3/J0UDW7+trCiuvT2bZxMAy
5KBN3t/O/2Gv/e1fwtLPDVY7Z/uhwIexhyU98SezsH6YrOwJib2YUKNKd7or3Q05XYhc2IGP2Uh2
vSlQCwRy4nhSBfKmWbO/S8w34b6apnhOuPvyW720gbA7ucw6IQDLmCbyB8ciIjQXfiGcFuo1RDQ+
VFCBDVrn2CEgctoP+kAsI53YeCpqkp35Rr2qfT3qu5vUuZBpiRGH2eSk/o5IyxseZt43pHgrQdZO
BEgtHYAbTtihl9YfsgbsN3BMFr2SusE5CavQVSmZgSTVt6BHp/snctEX/xmNkKgNyCf4aO4fzfaG
ju4gSsHo4k3BukvNGLCZDFhUC2AE8bb41lTtFD8bTOH9eCo28/yK2D6OCG+2QinZgr6S2A1BaWXU
kuHLr47XXFPwRgHWMV/EzoxfmZib9yDSBbpS/xpbL+EZFgWdZajgZLwyDarFFdW3tKwRzTXxs0F3
4TFHQ6IUnRCSpy9+3BL6njKLu0ElOh0WsGm1SZVBQUos/7JA6iK3CxQbT82iDA1isxBhzwfbE5Yf
Sef7RTGRdPaBNqCiWpRxYka2xTD/nxHaRKxmf9pl+nDv/CsLpiKRet+EIcikp5uSGLPgMduGCLTo
eMENTU/t6OGS9/uD5hLm0jx8fky6I621Vu4LVBtc3Wndxtn3bdxK4c41jdtoqUEy3Be9dtgKHzZG
ddiNiydBvNgXbb7/y+lF50PJvbEZEJ09fntozDeK4dLuMbYTvbtuF4XGkFMCkh9KA2afDdaEe9HF
6Vx2ZEWTtQ5sGtyCcDsuY4M0T4n/3cVGaeWN+fM7LWzsMfGF+2OoOMR+JpxNj2cHTCVOgb+keUFQ
c7N3frvzdlhhVo7Sbi8W/geN5jpVhYLnce4Wd6AY8xqk6LnSAD4+3nPzY+M7Nq3777bcOXUnobrW
DJXfpBU9h8+OHIp6MTohk4WzkTg6a/0HtgbQvDUOw61qmynVSE9+A8g2CNmtNRxLW+tihG/J29BJ
SThfCJhxT95rJ2WiQYGD/e/ZTgPupngt+LZU9YEhRHlWl8CsTFGN7pSpgPFQnoqOgTl6g56PMKil
sEj336fk/dzpg4R8Kg6zxI9Q5qcbEYWXjx07qYFbWSbod6xcQt27vtPyr5Jkce8bbTkL98/LrWTg
lBwq/JxQMJdIkgGToWfj6TVqfwfvi26VVP+XhhCVzpvlVi51iSUm32Tj0tfjzHB9e/IGyPH9EpF8
Edxn8vyzAyoEy6oc7ggHd/8WU+KZJ/lThyi21Jr3lXRROazDybK4YfvettqVvaO2iRY8ppfFLymE
VtNNaXmRFPel1VHWGtu8EAZ1rmb0hCBTCWTwWqdw5Nic5OYR70OP4z2FofzLisWlsFMgy+BlBJEj
8xHXRQEFryR5TcDiTIlyYlYQBTR0ncyog1rqiPLuF0QyNFhkTyGv27KbwQ/XPjVWbOU2VRwmeBPz
JaP6/R8jM9TnVniY4v6oJMr6qK5RHRGvM15+AhDBakJwUqaggpeXmleFR8B3PFxU6J4iGLayEGWf
/mHIgq2H+JgninCbwO71pYI63UJdSwnY5v41S+Vcn+AMD1cVrgtQVWnSzs717NJV7HD0wSnGjWWN
bC+YkxlqIe9P+WkwZe+MF1Kh1RoO1l/hZ2olvVqZscHXVRIyfgCewrahXN6IDtx543lWRXEalwoI
DIKBq7dX3Gm09opGGJs3qMQt7iDx6yf9UsOYhasPmRbjxjvt7KT+qnk3sUSyKAKs+QK81CXcmgC0
6ZQs1sC7nJdqO4QbC02FqzSWhY6tgQKGO4DS/PmHv+Cn7xsWtjdDC23Dd50tIUiV6MwdE7bLSuAh
k4tZz0PVMpEnNhYc3Dznaacp9Nw4S7j12ObDd9t7RIT8qYPonGpkOPTKuOKvanGlcqYtQWbqQZUn
dZrcs5GHQl+4i1MEE2eVrhMJI8wcxSL8ofEBU8CzKZ1x488Liuum/T87K94Ptc/1TGtqAy1mgw/o
htHB8y8hTcHfnfNbZdppatIKeIzkV14fdGrw9TPMfw358hFpEkShxsIkieNq9t6Z9ox1zU9MxOzu
OOpA/0Z5MOg1Tj+8qOsOzSZ1VJG1YizNIhQvft+bRowBSAd5v9vz3uvyueOo0ncGASlKwd6WQlZj
wRbhzkWeOJrWYQKUwCwGu92ApK1VcGdg6iagXMNi+h9sCd77syIu/uYf4r8IsjfDiKfFnZjm3NIu
GRns3LpjxZxIXt5ZiFm8pPjKu3tjcdqTQzwIj4LlLireCvz5sxYzdgpqFRzqLWNpS0JCkHf9t08e
hXvTfBOAuhZwom2ut/IRo5d1Lqb/9I4eXezLFMtEhe4TOkKtJERmvpKFGaEn3ICt9ji8WYwhcZfA
VSIM7cdw3fzcPFWJVHKuEeLfTjU573CzJ3QV4V1TjVNA3dfrqKGC4a8z9J0qi9p6hjK4r7gPknFz
r3ROM7ZjhHsG73RqNac+o5mTOu2rCFLj+3ro1d7eOoga7pZd0yLuHXzXZco/nhM+p4Vt4/ZZBygv
LBVIyBrm3KoloeN0vzEw7yyEkNaLl5Kl8DsnGlwT7hONEPiivPTeeCvM1NTjmIQzJmAohNXamel6
n73XyGwpPIkkm/YNyNzcweWk+/Lhe2TKzckR9M+xh99NV4xzn2/Z1uW/Q8CBIjKTQfPzNI+/FVfW
ojotTJCkvO0NsGcP1NufqmBVZn0VACGoWfrDeT0BieMPOWi6wLDxgo33zxzECQoEePkDM1CfZU8B
mqR9p/L4BtJjJdJYFF+SSLEUZJyxDJkAoee69uNB8pKiv15vQfj9Y5DGdqxXF5JiBapjRib6gmsS
sDV00ilTELGiFOX9W5x9DmsNUG1sDB+Ip7V1RWHdQINfMxR5DfnMgxsrCBDP0ywr2se3W6rzUKOX
SX1gqsUoA0CWwoIgPqXVSD/9rq1hMHkDeBc1O1hPvuC5fTQ03vRFjPbLRy/lD/CWhTTIMak4oj0n
0SPSblx9gEPQvVGmONFsbtlbGZ37PuuU3HfAI2VLvQ1YaPqlMH9I4XnSCqhxcTGHAtablx50YH0e
0lo5Qb4Xawvx5PQXBzU0l0NkiyNu2PliTKs/G6FNFm+7W6KNX2/evIX6nnFnL+50ZnXpNv2XWtpw
5utmOrAkeyF7sH1y6WB2YswB6wlrNbtwyeCCX0PhPCFzjupKQ6bmE7USkq9jCJo9m+7eAWi40F2x
JyohJ8xDHohVWYr9EmGwKBReQ6UvMuf+ylHBa6L4NykoKdVQSj7u5sSdHZKWcRHibhFs9giBmVPQ
Xdp8yEPW/D0UZin3SND7N/NIxNx0A30XaliZmnB/XjlO8ZYqUC4QMq0RSWBKNl3bEuiTVJIMQpfC
S0sq/ZcIryi1VAWDimbymSc5YcN8iNefT6VnLD7Gg+O6KCnDXC58h0LCHYLvKi1eEKCRH841K+QE
QGtU8DArLTwFWY+UzVpnY77HV/KyI1nGFjDo8r92fVhD275melOuvQXZZLpfLI8q/+PmHyItcqEN
QtdQy5fX6MIEc+JPUjdotIoYTQ1hQ7/v9nODNPdrqSEqaYg9qmZ9DRDrtY9vMxd3axbQAhHVDFDt
/2Qo3CvLLdaP3AI0ee6TbTNN/F7C7/SN5CuqDGQ+mAdZ8kcLeXNG54FVPRBET6X1/80UTGaQCeqj
d+63GkZU2I7w/fF5S/JzKRkP1U8I89X4q03UQfONZbysNVcB0VvmfwEdvnejXra2A7l3eOduCj2E
L9stGJv9sWu+jdanHEINHTxRC7tdCvf0G7wngjIxZl0b6Pps/ECz7+1510p0fELIkbzs5JQAvOmo
A8ZjcexsD6h/T3bGFFcIukl+mXnusjFBxdfSB9oEL4v059Mgm1tNWJt6H1J1qSbmSJYp12oITAeE
kuj4wTxObooBhCi4L09U+Tl4EOPkW9eXi4cWNWtI/o526J4gG6Eim7bugo7vC6wokwsySek/uXne
tGOn9mDH1+3wvKgdiiAQpIssMVLabgBqavxZephIhc0V1LrWW9Cx72WxXdzx6NDQTus1QGXRw51P
0nUHPGi7dImiYKT3JqPuFBWE5Xy9ixCuookHL25Hu3uoPYDxYxgbQuCgFL5C7UAYuuhKiaTkHf9L
a7/CiwXEzlnA1pkuW+7jTKZ5xMlYumVDbp0oKpt2royCW58BaepNsl9Aje1V15Uucgdyb3+7vyPh
DbeMj73KfJsybCjaYffp3afDovJXVi9xhzFzVWJ9ZizuC8F4HhlqMaYPUiwui8WPblRgkL2njiZG
7f+PM013NeHrSizbQiwlCCs3gxNC7XiNHyLMwHDHyktw93aXH62lQcXkrWTQUXGZRT8TBGpWjuyV
8voDpx+mEaG+DWvm1QV1iquUDXyDvcuK9teEHdR8OFYWAmC+SK9UaYYXfXaxfvkETpLmSRcOiidC
iyIBrut0GlKcsJeN4KdQ0oK1fKQ4YubClauXfJuZd2x+UBkRd8u/o1RMXObU7DIwzslhpFEM2obC
psD8pXckD7Ii/Ykse5NopWz3c6PDJlIlz5sqs778cSZBHLa0rPY2CsSm4bJKKhn6hzWgwK1x7rOC
Cv4TxguHtZphemxQr9UqODQue+GrX/oMc8ERvBax932GLZFx6IFQOLTMJhv1TOiGZLf7UkhmQpIy
UASYgFEa5B5AM3XnkPsTejaBSbCxC7x2uaaR+hzHSptHXSj8qxc5wzNzhliMa6irVeu7H7hXWCse
ZplpgqZ2S1fyERYtIcGk59Jbob6Jozq9Nsyza96xBTQYO8FY2FXmJXu7LIOijctE2ARinerfp3V0
ACglOKk34czVA1F39NMOpCDFCjrk6MZJ2NDewLh58yiQ2Dv+gjvx6oxj0UEBvFgQZg8X9g0uvg+/
XYoqLCzyrsycQFEmh/JYN9jNrew5GZN/I8Zg9jqQUbdr2KDsaDXRORWbnjRPhVdh4NOGgO0WAqL0
MiQZbBNYE7pdjBm6cc+2sG7uyz0eHxvKvKL7y33kJAyceSerrS25QScLe0Oy0faF0PhO6hXUQ50l
rcpN9OooBZLWBPeVhSaRzAL6vWZTAESYIJMhKxvkFQPrdiZmo0dha6qu/bVL4LJkPmDzQHqCFdTG
BoqVbOqXNOzA0obAsJPnBKkzZQfC1wFj8fxlf0b0AbihjMiPD7pINQs79AHhCxl2sZNzgfvk+Z3F
d3nLLtia0u2Eickk4sY+JpQdUxyP4yC/aBnKCI2qtVG4lJP3tgvK7vyIFypyU6X9QpdEv99uXOtr
7xNziKGbCH9VtU87FkpVEIWz4wTVZHFNfOb4Zr6ntvhTpJ/TpBSztwg117pHxeOBhsIBC2yucTLK
OI+Hywfg8h2ivNWJ7i/fY/otwzGLA03koOXt5jwsW3ivAWctTgyKp/gUHtWN8KDYCquHoYPKFHTl
l/l3Y7oz8cCAhE17iNv4ZCJmuyJ8zG8cVlpW+dufgW6NQFbiQDo7D7ijoUyYrYHM+cm/bEV+0VvQ
3eElqupLmxfXJaOGCG7njwg/EG+uK6QX+V6LxvZ7+SLRULtnqz5V/AFbFCnO5VRtxODAz52LTHXY
IF4Hu1qg97cYxWKEVWLCjOn18g3QyTXxgmTwk0YQEJ8Wq7IdlbMojb2h0b7Ajn2HwYYXdINJ1w7Q
cz27jX3J+QqkN6ywAeQ9EKgbo29rcGpPv9wvZ199IFPbeqHw2vd5utmbwbHa0fAQb9EOTbNjxOPt
CFAw4V/g/i8CZmDWka5rDELmWnxH/1RE6tfBoOy8jAbY6IJv8Tyi07J21vGhmKsHP2HyffkToHXx
4TOxlVkU+rgsX4SOi8b8fwHb05Xakukk4bz9qGHj3t5MJalQKQLNAMZKpLrKEqmVILEoRfzYPaC3
VxRgVrSQPCKNlxdQKVbbHp40V4rTbY7lp0MxjZ9+QwVT7Kvh7Ra5aTgSTNehRMOq2Cd9gqflEH9p
dF/1k/EMjcLQP/EuCm27WgmBdDe+RO6cKKkI22bBbGDc2iCQxzPWolVOlW5zJ2Mys8ALu33WNgfg
SqDot3p+2OXZBH1Fywz9ic7UMuxxvtkZ+Lk+TyMLfpBFhoSWLAxa+HdiR5DtuF7NuZyi6/fO28t0
g+xJ/kZ4SYQep3YmX/hYu8IEeUtUrE4n0XBWbgsoGZ/GZHRteA3rDC6YNf3II/noUAaUy4o4UaX8
5oWx5DN76Tu7kRwSbqpVZJ2WCQ20uaaoh8kZ7T2YTxsE7HHc3vJsvHF3zz4ePHe7woWrh0Sbg3Vx
lym2M2LnpTqhNySuucYh30pE+CSWG8nLbJqaoUJ07h+TuHjwWag7lc02rItdN1/MiOjKMWOhteNP
0nI4GRXOUq3MLmXYXYUg0zFsmcPwjpzX3OdvU2OPOQVjz5OjXaVdqmocBRm+9vLf/qA1EtWS2LEG
Q8TsHYI3y+xJuuYLh95hiyeOeEf+9zMG5pTT/NaPgOqqrZPfVbG40hxWGacgE1rg0nc/nZyRUEss
pavNlMohQqsntq8fTH9PbjrHpMgpxtG5r6mWlI4KpFwhox91i5gFXesYeuq7BNKfTU6BbkdeNtll
53E+Y/h+dbD7XJ3gvDYfSS6oC4Nu75xTf3RtvUAzuQJ/ZAemhwbGzzf6hvAh8Te8xpSUmukihAIO
X3+vNNtkQWH7pI25BRN3Mv3nyQ6ksr1t87gzYK6FeMjsOWBKcQV2KIEo7PEqcbpHI/vsVF0qkLwS
yyrdHruTmbsxTiay8mo1lJFcQ0i8UjkjRA5VX30IJdlhxx9P3ScqhKk3/v+joygWFduYWWI7OkFZ
ONQDQT+DguSUetnB7F9IwKjRSVHSqOMYbvBfPakqtWEzTfZUFKuW3LHdD9/WeCAudBR9GKQDHglD
j8EJPLVV3fEW4JOFxF6hgd6wDN+qiIrCBxtC04W9AcYek11gWbFd1QICHHVNJYTKYQKTc6duFm9y
EAFp07dlG9lJyPfHhA2MoLuvzDuqUD7Jx2f7guL07e48lVmK0UlKjdgpAnvN1o4VJ7VlVDI9Z+96
Jlu+HVH6u0/60oWjBnhJE8F0HMI0u/gknocTjR0Th8Y4Ws4hpbgKuOPkZDzBI8AMo46o9VLzUJlM
pnVrHkLouv348spLe3lyJE449VsR5yNbNukEzcQjt/o1fwvE/AMsKmQhXTDZaCEyqv8g3tU24Yb6
yTfJutI7guFn8D2oz6L5xG+f8ah63vE9g4cZtDdYvXMFqOAdZFu+c4jpO0F7p/ksX3mljpTpfmap
kMac0wlakU2jv2Ix5kCRs60DX+5sDXZub2MGkkAzwDRldBpAxficGfqqm1p3+FBgUpl5kw1NfAhF
OuHS0FytfILMskCmhIBeXTXzf/f+/mxLlh9N9uTy3vP3sICyPBTeCFAg/1G6lZ58Xp2gakGBbSTP
qU5nvSa7KhPXU2uAi61ua1MsmvGTJ1N9gdEQGyH+uXzgxPYj5eGddXM6uV1ZLs9038Ij58tXu+Mw
dLu3cyNOj2Ft6rno8JSUshaCCPBf4YpK1JZZn9lxtCIEufY2/q8416x6oWrAsBNaGJl4G2///t7v
pjmL849KDN034Qy0vnyd6WGCj9oQPioh6sJSm2mfy8Q9H5vToEx+CGzUZV6n/lfyneuQwdfrbvRn
PSmL0S++WoFVeq0udGo0UFmI0XkhZzLpF5TY36Zpj/z7VK/Jz8MaDQkLEsmPQzOrUoltj769TWb5
zMG8O/zfuxxgY7zu+7uhknA9zkDTVxnrUEg+cC66lUQAZxxcoHEcdsVUBICSryijpDKXullooxfE
z3O85osXjTj3IdObsptj+K90G/NJeGWsgk6ahh+t7/EluqwLLd8QRz1ZxsR4wKtphyjjs/4109eE
JSrocsA2K7JZiEEQfr/S8oM4u6uW9Nq6o3qNXv0BtVlNDJMhbtN9/nFs3rrbIFdlP1nTuW8opnfk
tyfxwZ4xfb9zQ/ll9BtULNeWqrvYq9ca5mWObSdRA09JpAO/FjJctmdWN6ukteh+gIJorEX1X9ki
eIbrJpk8zaPEOonYU17SucxX41qfe2MJt82z+hM5/m/uWufvTUAqAnWIRMtIa1L38zVee0bkJTXX
PTOZR/Vh3fJPn4gzZE1dgva4S7uOOJJsVc5XySQJ+OOHgNJGm9Yq47Afn4M4AVXarQZ99dzgramu
7MVRgut/vddGvFtCua9z5fyZU9uhb5xAso6LpxMoZW+54Xk/g03WGt7fPJwsDLGe2VRS6AOhB9G/
6Qw8chrmZItnQHFKoeQUSteLMK0he38GEUzPGWYsAwIHyxcJ4OgvsHvIVCOOuHw/JnsYpFKupDan
DlzxlLLG3N0LRFmLNwRTzCaMrULjG5+BZHPH8A3Llpt2EcaKHPjMNODGWczOd5q17MZaIHmLjMM5
qNEcByi3EDyo8OBqtqY2Bxi15LUswXkH8v9RhpbKHP+u1UQaBU6HyI9+4AYBNhvDMwtT7XmpHi+A
XoetvNHgxREasxnA0YqjGZUG+3bnje08Ze7GWRuyoZzMb3rojxWXPSPLYaSB51YwSXpoiIUF1ICb
NNF78InVzvfz+SQWto0cOir7IZJkfHOZuwcwhiLFeRWf/5bsuNNfDzN8aQz+1bOvlhu0SGUl5ewy
VG+Mg526d7hltgMq52mbkw+scJi6SG9gn7FYe+RvCQp51Q6lAax04p1xD0h1OfmU33anaezp6/BJ
ZarUJEGctzJ/CzDb+I11F1ybQh7RYqwS3veQqTUuuyPuHUsGPkytihSTjOzPHN2Jk6w9Ne4G9+ZH
cezQcYqcOHI73+Kgi8Uvt6U9g7PRiOKfK/pTqvr+H/rW24BvN77EdWRP+tduVOWxk8u8yHEnIcuO
aZU2T7+EXbyCV5OCdwskJwWf8fdnsqR374CUY1ujKc4/n3G5G66WaTE6i5Cplu0WuQKSWBi60XCQ
jOCfmWm1I3eD41JuHfmRElGnEOhs5EgcuKQ4rkQu79vtK9dFhPYpr4xV4iZqRBUNIlFk3bdLOrFB
IsC0IzmjwaGbbMke1ZimUZWxlIou9a37E4ivaJFsCrmO6NtFYlvPUXftMqws/3S0gAW58J6HJdee
sczrpQo4riz+xSJ6AdKKRZdImTFFXaTNigG2N61TOtYPOKd6NufZRGoVEMW/zMl+gmfycmf6ih2h
7/YWKBBUie6uCsS7ZtjD99xh6gQJ95pn8fm2Yf/JAj98HLCmwUsylp85sEyNJ6A6iOlJHtqLigUZ
iYXD+KeRAHrRZ7f/lwHEPDL9on89NLdUC4NgfOu3MTflwFtD8felhMnssz98L7eI9vCgXbB5z3c9
pk9gTVbENz2+3f61ai+9P7bk/zD5cJwL5YICTVGhDa13hMs4f6vOU5uQ7qHh4bWx2Kzs/2DMxsXi
4FAZ2SXikdapdU9+wbs3/subtCRja/zS+a35as/LGkf7lw4twKZfVDqmSBdAlEvw2dax/dW66cFw
To0hxTLCb+3ybIvKurM8cr3NzUFKLi+fWhyAZ2gKAi/lojr7rxgjXG202V8XXeT41HdfAnqYw5J+
RGYsDyA3gtQCwgCA8wihS/y59ZdigTRnEiB15APCafbuc5k7dXdbsaw5yiN+4WQ3HkRZ+QEivCbl
xrjaL7FzacqwRSrdcVN3Q+BsReRtsPn109gyL7ogbtZi9gHEUbdw9K1KLoLb7JR+RGryJoOHI+Fs
5MYe8zDxUIO2lnfWQz1udBiQEM1xtQxp0lJRw3wIPnBEPcbP2Nkoh5bizagmWXvYXyJNlNybJVEV
tCmdhjk/lnfXL+MVJRJY9cBtsuJ3J/w735m5uFP9lK+bPpPVK5WcfEmTrHnoKEZEOf/GpNbb7B9d
MqTrkyOb3xeh91aJkQci+l1Q1H1iRR8ANJDiE0b9U0kVWWiBS4/WoroJoobdoqnJO83vP4Vic8n4
dQpGDlUooJ151t0yxCtAZsZzau1mhF+9hL5qjJkPTWFrc9RrL1d7+nWYP9hBqtMIDaBbpCt1acg+
SsCM+9RrKDupTQAGmlOG1AHPBEEboyCsb0jVp7xN1Ejt/7NzzPpFLhyP2Z+kpqwiIWivArfWPcKy
X4/JP59FEHWha7ImvTWg7CfOAtuj4Sp+7x3jsqzRmpuNwyfNc6XWuz47vEixyXn8c/A1HAV1RtMl
1gNQlVov4cxekR36u8xSkXblytJiSyLIUjW9J72/VLP2alx80xIw2fEw2RBeGciHVdzb0GDrH+c4
LxCH1OVE8gcZwM0ZhVvtyYRFjbE3bxSQlsSmORvW/IRXcpih4gE0WMuceOrXOgkXsMthBrS6/Jh7
78MtEub6GL7bjvheEz4WNuPhJUNAPAUo0LHK6PtjYB9ErSY44QGgJcCoInhV1uiwHkw5tOmNs3Cu
u4aMhAZPfLv0DgYI8Y/8eDZxh7fAa+ZZJ9n1sY+Wze7QsJyb4L0BmZEJ3KjDhljoNImt/xXGScFh
g4jAtfC6U/VbT1EnCe2DiJi2uxysxRsR6FmrtHIZKMi6wMKA/MU8NYdUQtyeKoMKjIm1L2VjYso1
FdXyNA/0UOn3VG3487lS3W4naj3X2YDC+c9j9xZOZgOEiKYnGuFxCYEVQaQZRtynUT5pDSgjE/sd
nX5V25BJsOhVitHqqYB5ZwQL4Slprw3JnS7Hb2fJfmAn1CslzhP3xxmOdwGTG+17D2namMKjMA5O
PP5BQg8eMedPrM3dhdRaihfMcdm4kJiy9RxtwJAV7zgJX0dn14AQ+Fw8j4m4fUufxMZFB5xxpeXx
0bcjFZo80/MEKgu6EqpgU/3JxVCdVdZcBenR2FnSW+OKNY5tFQZiyWYAoP8bhx305sTUREXSsuPl
jgSMlQ6XTD8+p7vdeTN/VrhC88/WC7eSQKVSYyD2EXuFAZ/F+tNeDJeTR4iLNZT88mAAzu1LMN11
YdGynX7Wx2zE5i8bvBo7YBOY5A35npx2U5pqjW5xn89fyojr+2Lop3AaDwqRGl8Keqiqs1oudRaM
SElDaAqJe41AYROZiW0l+2U6js/oEZnuH6GZWUzho7K5mDdik7oC+zT/KKz40z+SzfVLTB7s0FQJ
gLoc7FwNhwyHp42pK7vlHU4pzZERZvcAmYWWv47vSx3kvqKt5frgG4xPOgZb4j4hvHOZbb5IDThu
USI3czy88R4pfXzFG8V0hW28FJ7SKDXUQIAWEd6O84m94+ClF5w2DBlgwJyPml8td3Whmf8rVSU5
TO+XZEo5MejJzdJk1ZmpYVtaHuplRHtJ21h36wviheThtL+25EHnejxxZNUAVI3/zquj3iEAht+5
Rl7T0MFxdEC+fSb7qAtbHWhuFcLlpRkrBr56xML51xUrgb+1SsoI/lLqH3mK7LuIeiPvxQSQwL1I
27igKuu3KC/7shHb2901BinnAwSj6M+cbLUY6A5jNvZpCTbJhRGvfMa1fPpsLkhqx278HPxf/Udi
LFvMWdpEnk4KZr0tzDecRUYwv6rarKwwB95YrRFjzPNDaEAepj+uvyX3nNZ0LXyd53gYCHsQO9vu
GWfd8zrDf4cj5kwwxMiCTVoMD4TItH+iVP/A7e/gV49I2n5Q82Ij0DQ6LoXGxjboPX3mw+VcjGxV
Bj4K3wzx0hxo/02v0l/R/YxEwxzxgetnz1ofJ/8hH+4w2Mouep2ET/gO0OA+udo/9jNJmrUQe4uz
dAZeyYXAura5p51wc3/69Ssfuqqb0uHTgvWGbxq+HqeZkCJoDbvF9VE+SFz5tBkxbdI1zzNDBkrQ
ylFayUGanxF+SGHJfT+UNKLCkRchwmOKeOU10WO+vA60WE+WwTSFDZCXXjvDX1bnoUv858huaEV/
RBn9A3zMsCN6qQlR2Z1rTu4qqlY3KIVX4TtoKMzWcYFRg/t8AvB3NRj0HZnGcm/J5Wg1sX6VDZYs
4UOe12u4xR3pgD6BY9aY8jqEASIV36kqOa41fvkNE4YxBSfBG9QUG4Lxsm9lkUnTcdZwH7/KNror
yqcLumNL16YLIU30rSRpSpE6AKW5eCm2ydPiv5S6Af+263pwQZQaLHKGHgc5RkpSJ6oIhiKfnM6S
1PXUIoQ1oAAHsX3Njd94GAP39UsqjA2fz3T/xOSWpNiQ8CIjgp24dvD1uMrb1iS3VxSHDguDCZND
C1zuW5TX++5M3M8wrRmu4vnmFy1aUFgh1hkSIUNAKJruA3SvaHp7zxk1a96cUvoTWhYSImsoZ5bP
+OA0R48yBX5K2ejeZRuSAAyP4vlawJrXw9Db4DpVwO2tb6+l5+nH3WKoKvghu7LA8YZM/J369cUG
s1yvHYLBGZHeFd93Kv/XiNRoH3cGO+eG12q5ltXdsfdm1bu6LZvNpXz1ZJpSWZG/0KnCGC7V0HkJ
ccitaszM4PYasQSeA9EIuG+k1sgRS2k5sTeKPVg/dQTfquHz/jZrJgtmcGTcqbmFPaDIiUEvro8+
Z4n45nA+lZ1GIw8Ib8xsn7olXlhsXoQeOjOO5QPnADE+mIiZl04V0hSN8i+3py4WhaBqE+cY/5uG
ysqSDAHlRz/GBRWYGaI5XYmLvuTY9myezzeYl+W+VdFlBtao5YRtJ/hF1DB2J09qkubFJrZsmgFb
TVxVKk4xs9nUJYYV5rEQnAunsptuFc1E7gpkOy6gGjMVAjHFtzqBel0rlvOKU/5lkatG3s0nUAvO
W+5jmplzauPuuFrp/fyE5WhXmFFf51YUNnOC0aA3TJyLyrlBZTMQmuNWl0R66ujJhhUvXgyXJyLv
Dn7hv8E0K9RHXqut5bj2NRCXZbHdj3RaJa9uov9r0rrLazmK1BA19P684qbsqx77+unWTkDuLbon
fWm6zm5UIQkqoMZCg5+jRSfLU+bszQpzMhvJuE7wqg/AJan6KmSN6yXtRUUmDkqMP3j5BLuxf3OP
k7BVDdSW9hQDvyk9ODv8hamaZUNUq5mq1wTKYt2GIJBSy/GdRRj6ikf1sRuUxXFgeHeSIeNnyM9H
ZAF9zNn9dN7Ho94HTOLLxARugIuCZfrUPihbxcy9gLrcH91RNbPlnvg0D0ZgOpHKPmhYJIcThJ3y
IbnorqFebRKhE/lqkQu9po+g/hdsS1PSZbPSQ6J+ZtAZv7eikzuYZeAtSSD7WYVyLIJW6pS+5Sti
Dw0/Gd1oLDnJ2dQEMNqkCNpZ+spycEwCuQDTPaLSYLbtKOicb0AAEtVTmv4zgaVakGUFRKOdfEEx
kyuZ83Uic5d8UIRfJ+LyqPSQ/SOonRnI5GtYVb/CMFPgJovjbM101PGdf3Q/Zkd+xgud7Lhe6Cuw
TI3j6aTWAZwzgn4VuKkGoWKb3v8XxAwotnCcmbY2akRmzMcsHPifHTh5aDuLGDK/Co2GCAfcMm1q
5X1Gu+nKfNyAjN6IniKIlpC/ePWLfSi0ETyV3RFSkJdTwFyb4fEfHLCX0sPt8Ez1cI5+JeTK6c00
RihAMOF+Zt52mZz9eEgLlOQIk1zQ8hdh1X9E8vOhNZs+xE3Glqld6zAxUsJLDwfXM7nEVzf8J7wB
A3wYWGYC+w6Huc8fO0A6B+svT7PHad5LXRQiOnQJ8o/Xm+kGZ4HDC6FSN+xLJPz4AbrhF0SpAYXX
myOsmp6QHnOwxSXJUkQBiI4W1Vd7fj/27HOPCp5EG7OON4wivV1M52Neoe4natbPTeqfxZ92jmhd
Y/oZRuMkEIhsBLGJ0r/myININUGnlZ/ea0Jimqf2SDIiv/DEHHOzBb3kpR5yGpNJnqjdpfvWiz4Z
iv5Shrgc/4lNs3WQAFi4VEmhmFkwGT0k5MruvTM+gp3qTsldR8RDJfQFQ0O3D3OyDRSygSUk22dG
NAVTQccYF8sIrf5cov0rjngN/dH50osHKL4S/iPth0oXlGDPlM9XCOliZGwox6ekL42GE25QG61V
W2atLK+KTJyzg704U1HKfT0EtPEiio2i4clV9DWs1QPTxFGlmb9jVkQO1SsS6RZdiouay/5CDGto
i5nbFLeT6XdikbVXquwB49NzxVuU0DoKg4EuGzi5XDVb4LKoAubM6pLKvu7v15x4toUHDBdEIxBl
5Us8oc8EAmGvhRUYBYSIS7t1sHMA93guZIcEJw42oRtJFylMg5yYvOIFKKTsdbEghq4gR18o/STP
fXMut4uV/nPwAaER/mhXXcynzdFyMGNjaXGCyk992JQzBSznn7MAHfejqAfy0FBTg1rAkI/Zfv1X
Xwf3qzXAScJGlgOWkDn0PEOw/qyPiIxRzxhcx3Mwpb4hHxZz11e7MuaXKvBFRGswuwJdX5X8TGMA
uPv8O7VsGluXUuH3BsOtfj9r4l02CuOZLYRLo0XGtbKFLnGKL2cLJ/tnpLv19CwU/+d/7i59rjKB
NC28Tdy8phEp7FpdkYhDK2oQa1er7Za3SGp8eiNLBG3kM4ZtjeKP8/KNqir1f9re9ZlAU3utop2W
IMlzLsUhsY/iJ4mZOmOopXQDMkxgSgoDOWDiezYOcDQQCUI1GQx/58GKr7hpuikX43lwzyadnzOs
OLjGx/ktFfl1SheaEPPHJcqPOeqwqr9daSy+d98QO+FCbAHgVr3UoB84L9m+zXxvfKzhH3xQTAbG
urEZnMAepjhAPyegKqo6Np2O860x03hKFUNP4bZLv8ebvSVmnaopK7A33E94agzjO5n4ff3UaP96
D6xIJne+qZT2BLhj8xFJ4UkE4L1wO5VSekTSMq7YeKiGMLZBxQaLrT6PyxMGryv6B1kO0o13NoOG
JiOwuj5UqJSuJpa7fmcWAwf/fWQzS3JV4EYhUlXHmbP2FOzK41/UAHq1yQWIQe6WP2My5epggiXK
NjbO/QDrAi/VvhhDNPlEFs1SPUHq3LdwWctkluu+RDefFWV9Z3W5aPdzGbYgZRzVglCFrfw0lu0L
UtFIyg8c5w==
`protect end_protected

