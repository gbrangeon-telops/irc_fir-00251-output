

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nqqBtmqfflVo0LfdOWD2OeylbTCJPLX6XaSqFQpCXkHX4TF1QAXZspyiDVaQlwRkat06cPZ5E411
bTzbr9/qZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q/X3qbnpTyRXgHhmurX8chlDRL2XjwnbHjo5m2aoqrTNSVAUPYEYGIGJVoJhRP1Bd27KZbGI0BFX
fZKfju5H4nz84jXPUC/rcsp76WTu945qoXwdo30XI0Qhi1w21P6EhLXccz1l4c9zfTwlHtVuYV2c
xkxHRh0F8KrrR61HDHc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jBFh6UBl2pQmyl/KNdwY4r9ld/Frb+RgwTVitzK9Y6Fp+6xDwrsib4d9Z9Trd2PuW5z5/ot40n86
vR7VZpJnONM8UmDjWgdiB8rXNXaI1rBfme4TQ3jj6RaF803c2cAi4cdZ4qM3X7V29W2B5HXbYsfA
+fn+v+caVjEUXZHZm4HMyIR7TNVnvmCWeeLj52d+u3MrD7UjjkqtqnRWdy0ckM9p4TE27eiu/nsz
awiAJoiVLZNTMmdaTdZ6vB/sS67SAe0JjX1nTwssfK86UYU1+n0NLZ+SLB4lkqxmhepGPNojfE8p
9hJaPKOTV3d/umJbTV97L90iPloNPMXpGK/m+A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cwUUX8orCEMoCaO4wbzIkA5h1G/QOLlup3/J46IxMYEEhFnVuE82RZ46tcCa958uxg+L9/l1SnQ1
1Qa6GFDzaEz3zEcSDS+t0jFMPNI7VUppaIgcalGdkOXBIX9fihrhASeWjqmTDrUSlTt7Vzyo+3TY
n3HFHRbTrCchXcVswqs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z1XHzIMnint6AvJuhSJyN/+kraiZwIT5ZFNyZxcRS4ee586ZcCrsBlqjvo3awgeNWb2yZNQKbtJY
UBJT2Ww9PtMdwpg4MPuZFMCTECdiBOLjqX7gX0K3iBdA+35RXRVkpnaon7ABi2dY8SU6a03iv3ph
ed9P79UVGmdGucbzSQNo8vkiW9pS6ZJElXKmEibSc0C9Vw6VmCNdLosnrss+vUEVkPDu65r8MqDO
9/2zcjIio0kfnpSLOaIDXqGefGNR89nRv/NxKymzLnDjvK13FSfKq6qNfA+cXOtnv8oRuf0tdkh7
e8F12j/LQajA5bXDfmPQ3bNX4Qv06vuQ9+MAAw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 89616)
`protect data_block
3QvD12vhncjedeDDU1Q7W+gAaP3vJme/lhEM17U1EMjDIfOSMm06H/yevbvPXkZJAZFNLRZSlXmt
mk4Uxf2NL5U8pBoG3tMI5T+SRhMeAFfQORXZktmJUiuPB5XlX05R0jmhrMc5+CzTnDkyOW7VkKeK
xmkE46bQc7OTQK1VS5tdFGzWnGxv3nxr0sa2lkDp+njaqfbGdiWlDmSoTGYhQ/P3bDTnyCfPw1Pu
n0vaalUZjiiuQDMz5r5ngxy7lHAhQt18z0BNH39ZObW9SwoOPy7m9OAk6GCoxbBtE9Nbu0Ytm/iI
qN9rpUeQvY4gNgkhmXl65zJlGy08bTOEphrwQUVfd4WzanE2kOrZcpJkB6rZnLX8XmZIECAAbruH
VyhFsgJOirnD8i86BtZFZN0ZcQCeN1v+uWa0iSvLH9zSkfMWxfqwRIawNY8EDv1itC7M8EBbAbBF
veDA/21BZkb7HF+CGYBunN5reRXgGyUWwjZSyJ4emP80oPNZ3cismGNFm63Pe7GtpDppH7awbQMz
R5ceDTgQq5j9CLAS0VAhC4zYmcHie0fGsNaUCJyjB9cRawxWpGNDzdyKoOhgG1/xIofVmltIll3x
mfYx52jvDE9QQxTgiqJ2PyozlWdI8aaZgw269b39sWnH1bbyHn2ahHmiPcsX51fdnqL1MHMdVXg6
NwPqNyLQ40fdoaxvZKEjzJUcoW8Jr4O6OcVzFrP9otKa4PN0TxF+qdShP+bgX5bVPCnURBkzeSuh
XKbW/gTgaNQD/pk+au3d6h1SRcfPM0sQSpAfkPHEjaDgW213vZtYerPLJzS8UOqB56XhWV/gLlnI
GYf0K5B2dtOdjZjfy8gSndIFJq8yjgjwq9ru/jZGWgMfUzg9suUsaT0njfTp2xjTcmBsBB6l1gxZ
35rqcCC752HV/zoT/MANLlcEjpPiI9ZzaJvUkxQY/SVM0CVKPSeJ50kMbui5DUvkcR2pyfJJ0MXq
Qs28g+NsLkbQD8o9+GrRbzFmByX0NA/BfWME2lWxPtt7ILFWWcvwboVGrMlbKQepctPnbsSz3Zif
fcJtjC6+e3XIc4FF7pXijp4VBzhj4xX1cUJuMwKvtvePk1Mx5zDuqX7wH17sxmL/qKwuU0Rmhw5Q
uhTglZFMfaOJgyZ7S4NIJAUna+5yMfueDtPhHvUem6z96TzAE8izrjC7VkHIMISA+OPwKxmI1ILX
vsnZ0Ni9FuAMAZ38ffqEmYGiXXgbrXgPSdL8yD6lQTmxunaXOLu/EMSTckYjKoAluGyYpLqkY6xD
8Ln+JuA4QAfqxnfEIP8bCyHOB3F42UuCTADI3Hsvz5SXyjPas3uC/IbmOIDN46hSvFduVZ+x7rR6
U/1xj+Y/z/fbjPUyteOPiCjAWgo2h08vw5lIDaX2cGaEB2yJJMnNXQXHU7vvysXSWh6Lob0hTGg1
FvCKQppzXdweAStUCgoJnH3Wl3uNZ/1E83y3uQVE42JdltX9HpLEoO9wiBvvQNN75g3yF1SbLfPP
zjyIFZfUSmFkTGniikODv4Ixi2L/fGe3coIKrvwvBdH54N+3+sUdi0vXd5Z0BOAphF5mogMRGX+o
lJWOz9rDGUdTJCKFHlA9tgT4ryUYrDVPVj/a3MxvrHR0ydyTGYB7IaxOSzWcdOEPxIEveXUA5QEm
Kv0ALjSpGbwf302KlaBkf/1tIbZZepKgddTU1wgX3wm8irg84IrKRgNvB3jdS8cb1ZPp1CCjcvPd
7HqiNPTTkKk4EAoggedH+590mFbNBi8sNzXUraklseJAL+nQ00l8SWnftiXbVR5SLDhfUQ+mpZSX
+8u/dS6woveUpC2PpITWFR7oF4yXgz8XUY4hQlwaQKd/Y2/U7z9nXM73q1AF9cCjTsauw1ypi0I6
14L5eIMtFD0y6xXfdVRRB+7tlB190pfW/ziR2pYpuLNMl0u3tB0NpQWYygbsmjFU2/AAwn74Zm3Y
pDk/94wPRQjv65uyK0j9NgmJwE7zaUjdgpLBh6+JaAe+TNrz7zWd0lZ0VHDj4wsqFgbduHbi/oPf
vb+5JjUT3fmdAg1UV/iQtCYNAFkgnc6maN+MoaUo1jPkh/qRd3/idU/3x+Jai98fQ4gteDqWzn6r
5PwoOOCKcPgLuzimgrD6BuuSOB6gjhyjwUj9GQMokNozsV1siKIKc1MX/Z99vLWirgEX7pbkiI0x
AEWweqgs6XoAl363nepkObRFrghRLJlpsyK+gM+7kPzXnKByCFMB3l4GztuSNtD2w6+a/Ckj061T
nZVI7VxPvoHdrIUM16LAW3b6OPZp3Hbw2FJYSXHLX69zwaV3ej5fngdO1DDk09dGR46DxDwwxDNO
r8sPKc4Ha6RwXWwIKTcWhaiDGsYgedT5i3+P4rH9/NzM7COgCx4Ha1Jdj4Ft0ZAVwGPs1+aXCeEk
6DYKam20g7w+GOYSZaHXM/Pmb1aMFoRMIxmIU1ze8Tz6k6/YQzKyeXlwwRBIeYPsqhGkmAYkem3q
1xJ2wTzdrca9YKs5UJVpKG/4GSQzVTsF0BWP3l2CVysgiWhQLHAYeW3C7gczIZDxzO3wrgHYGAo3
fGvcyZFJwuj2nhGKeFGNJzViqLhk8extQYx30w5eCmQjkW1rn6V86c2iWIbIqPyayj72TuC/bgZU
gbvdT2t+iK75FJ293+nk3tx5EJuD5QviGQd3+nVh3MGmPsrM5slUj4G9We+NgPU7nq4oduWV2QQ1
03SlSwauSHpZ4DLiHopCi1TPhL5sfjjpma9lX6aB4mWuRL2v+qLIe/a0SNBBK6cpvEHfqoBzZIB+
w42oTW8Ju7aBdyNU/TNNyFrkjzjLfeR7A4iLac4MsTDaftUDkm58bz71S+SOsYzyBYeK9jdFPPIo
S/GzvnrK5m54wW/U6fhK+HgAMjUXc5RTAFeOoR3SHLYCjMNBdT2s4ahdQg6JGKCCpNlWliRDLI9v
Vz6uUtpWJt2QhqU92+6aSN2R1fVKYBFMDeZVQimzdfeG+TtuJI0X34oHRLeoQNT7QaZq3EIeyvqH
Tn+VBcvd0HKvj97U3SofKXcGgMdBMcZF10GjPguWeMuap9zNhUEVE9HxA87Vpj/0AQ1MvJCsr5Dw
Xuv6Z0Zy0pGyMzTjMEdi7SayNKoUgtt0CfsRE5oT2PhpXnABJRShmNhR7o5VrLORW95a5ie1bDxz
fnanMYZGUxrYJPXGyw6ZcBDkweVeop6Huff2vZ9E8k+DmvqXOBIS9/odQaOOjmQFXcUYEqztVW6/
8jZIvwsQz3fmRotZyZv+E/9MdUha9l19JqiVU3XUfI8UrrYFhJ3Gab04+8/eHv80VQzc34SHWDjp
O2riqxPxMwDlIu7LqrKaTE5oyPjQ0T+AW9WvoG9DAcZ6ZwPWZV1VOjZ7nSI45IVS6JInceDMEXmz
I390IrQxIqTz8a1SBtJs2Ec8hiEVmLUHyp7fFCznUrlU1k/NE8bhs6bA4jyf17+Bo+LOaIacguBe
g9K3LMxg3Tr6au8DP3g6Uww5tsT5O4mg4XtfWDioovKcP+sjA61l34D6JvOYHpjGI7arMxSBK091
TQTnEpMGDq7DSBwdrG/mnXPS3Gh+XH/iqtMa5rKyOz5h2ogx6uvIM8qPXRuG8ChGFPmtEQpmcFll
CJUTwVo1sJhncIowY/bMKhngO0H/7CLVv+UBnOsFGU/ISO3TEEFDgHj9GsDRwKnOtt29HG/4OFqF
pZFibV7/+sTwHhpxKQ6JpPDvjKxI8TL0uOwhwtvF7TLn+iOf0tACROA46MuTT3Cf/EbzJDp+h0Yd
MTHZ6sbG+/hmESX9RHchCQWR8ERf+Tl5ao33lZJTjHM2AbjUsNEvf4KOpOoYcEXDi1/ZAQ8ESWDK
ujpWKwvGxNy9qII+56xJmE+ym40FDqztNuhJfk9F1SmC4yeKkscp+HMXDhjaFnRmKTbyzMB2p/lA
y7MDWskY84HB/CB/a507N0DTm1wGLi+z+gnNrsimE4SjFOJPUmQtXYTSPxuxL3TbFgXCpTgcb7rb
YLVjAjD6s+jTYkgioqkGn++ZixYSDoXyz82kId2sxGpZSrDvgXHlpSJ7xe78QAZD8Ll/UTX8n/dD
iV84X6gz7cvuv02DE12pExt3APee1Isofbp54CZ54I/h0xUQj9MMGG0l7v3dFnTUfTKVgIO5ZRmD
xV7z94mw+tqEp/d0w7K4K3Lf6qSIB5JJULqKU6ugqCZ7PKE5/hVR6ZQij747OaBOY3ivJhAj2IJi
0W4Qt3sSWcgUPZfhFAMn3eO/xpeqdaGyEFO3XJvAHpXXXtAC3H4EjqL4Cv248FCWUcsyTCoXgKpu
uBnp9z7Ym/Tf5F+Cf7E08Th6uMnR0PiBuZwm8+rTBjVkFcgIT+lKEtB0NspymBb3mOcpRtTk0w2I
bs9rYrVwz7HasqAJVnq0mmJGKAodh6xbkmZiJiXMrWHfZTkRa+LT6BFHAvHirL5fivKtmcp3xEoB
bTYU/62nxX3tZsSupVcIxAOJSDeF4py2feJZWvfkZDkMtInkRmTA/5wjRyjt95JT0xFCjgd++FEQ
JMYyKVILEvWv8zswhO3wL2/ex7ylQKWIlUaIocYzdOfmihsi1hO/37uesZKsc3anrPOj9Klhkoxh
uHVZcL1LVATT+TWgWfmNwV7E0wiBekPdzEv6UOZk4A0uxYqTL9pH1zFt+8sJoFVp5VKtVWr1lTdJ
fEnWZ2XcbRJx5QeCtUp5jGF3oMR4ZOkW3leja7SB4Nc62cIbVoRyq7L3ZNsLyHddZJC4TvnE+xja
tZmV2eKzgV4zNq9cQhQOu10A6kFOypeg2HA6Kc/A14hx8KuUo05zMWFk/6Zd6E77luhklVgcNBYh
8LRvGuh0ZzvuRkF/lo3iKk028y4VwxA4JAh/j6FLStpreCYPDPWez57JUaikqE37g6aWldMeBQc6
Odc3z+pigQ9O5S0BAhEabjoQKKqEGRhNiMlOXPgd4onIxPIKQvHsSbSczSkc36X/llydEji19iwE
BpztsC80mahWF9xEjHqCURZytvVjVSgrgQNbd1ebJdBNrNDTp+A5JMgSJI9AQbVA20HLhVYM60ak
0fjPdi00BOxGC6Tjklwwz3R/V717qt/a5+SSvODbo0n0CXaUKonTQVKW5jDog6lyNfYzzb/UHIq+
g8+OnuJJVnSa77D0LikuPJUZIJOQ3z76RWZsb+ybolCBv2THhRnGiBvrffdMbh+Rlfdz9I8L/OLZ
guWhvK14cDCuHnHjnx+Cm7HdJD2OzuydvaVTlPhj6GqpiR7EGxzdlhCZYvwFgBlqz5i20sBFQU3j
DiKvkfjZ1Vwf1/0aFIta8o9OAFgwCQuwkcwOakNLbS8gGl8FN2Ybl3I7uZKcMDmQVrZ/MhQLgwdA
ydUio0g5TIZlwSb701ty+vjs9NtKu2YBcV7ElYTt+7rfXjH9H+EoPwNSKq80YCYluu92iO8HP4xm
3gcLJwx8vIRiywhnuxcK9h0kcKH7iKFHz6NFL0CmjymfpXvZYbpB0sl6G++4xD9Uda6m76q4KRv4
l3G6sOZb4qCO5oPAQ+eBD6fmtAreF1C81RC/i1JFmILT/BgHO3jIh+llcLmPVklxlB51qKPXwijS
WRQv86icjYBJ+ngnzg62xXkXYMzl5ueXv7NJabDc2UHgHKwmH8iygsPzXMguwHxoliby0EiF/rZ8
I+dfalWb16Rg0+cfaC/tjnQEdbW3BdWO6J66VawvhQ/nwo2/EuA0Z6yWBvXxmVBpVQwWhjiXTJZA
dyZfXosqLtl7ea8jbPgHAO6rkAOIlxXLwqGC1pxVQZrD/v3KreyIUHKOeITX0ebxAiRxEIJooqJZ
MbmkZ9Uk2MW2FAsFVQ6ru2f+az3irJkHLdth1suDCMRbU9HFFvFI5jEV27wvoOidyMttljVN3t2J
efFPtPao6kAxFgyByYHNFydFjPhSob+zdrmvxguWihMVdrgwQ4Zwz2JU4uNXIls1qFzb/ikYPt0q
ChHVe6G1diUaLESsiyaEkjYMyyym5M+1+Ix6f6e9tb3+1FvvnCTH9hkDDJwkPpLQ+zYzJVHtDqJ1
dv+o9dxOj58SYkc4t09LLh842VYjd3URYcKtdo7Qo7CFNzduYxlLqVzfSPuCq0Ldc+OsEE6eS8lf
w2KBEve/RWfQ5iTTtnPAh/gq+Cox5ZaX8MyS0CbnpWutllkncT1w1mvyVPt/ZryiYvmNRtpYsovw
+A3Gk3TiMrMGHMgAODT1qwkTAj/k9NTU1lVHeH9D7OK/rRtDxCqQBUtzZ/yghZazoKNotheRuEBy
m3Z9fsc87I9D7tTvC/mcAPrNmlcLnMIwhykxQeaMAIBfmeT5MZobTj9P9eKqFPtxSBgjbyM4htE0
8h9HlAvrfiBkOzl4XmIDxDpmpkIDsXCcImhhrUtYoT9yO1fNNkt37i4RB9LmlC7DA7ONBxUX5IBO
s6Ko8LMvY2OG7pt5p8OnbyxSVdlAhIPFWAG669qZZApJWJroU95R7JlGOsoh2pJxrgGuQ9pUWafS
wnEV7Xse4fNKvZiyRWivKkwzyQjJwvQ0esr5uLePJO1MlQeEennWRIqWKUwSDky7tzwSKy2TnlX4
nk6eM+nmRA30WZa6t6QIE0F6gTp/l/AeuHkyytpg1aZL/E+Gq/5u86Jv8MOT8GDw91a9AHcm2e13
RRRqgsL+AFnpP+lxQrWXRz6uVTKfPfbxeyXneeaJAB0JPfvo8hPHfviIKCQUtqS9STXfFsFkwMwg
i86ND+U9BbeYfsDEMW/ITwlvx2USCdMCReUBeq6pF/Lqo6kUijG3RPQ0JJ+57QWeH4KoUdpnXrwS
+VCoK2y+zGeL883bkNs4hkrug9Y/P+h8VOHVP59wKrzLy5rDCHrCnzJkflKxbohFD8C8/T+WCh0C
xfCGEsUCE1SqFK2zucT7Bdg1P4WJ48A6USptiZOtTTe8qNRcyJqJZ5oSeLN9wrL8jSJSi8gz6Iuj
JFqb8CL9TAiTofw8m1kTCAZs0n9MMJPfCYjQyWl86lHvBDc00YijknJuDav7/1+0PYAuM+YrGHEa
fwAtDUyk0FDP5hO4p1hUYCSx/MJRQPJBjOhYiDtHaQ2Yb9bqFIqf9Fz32lqbdSinnGh9WZCZol9e
WD1XR6wu1wVvCdGhITBAB/SK9TE90N7FTUUz6rk3yYbcBHamVdscbU5za8i5utm/pXIbv0XlDYdw
UwZrL+r2HC0YDf8q7rfTcq6TE6iKKuEQhyElH5wbAyc7tlmfLx65DLCJ/5sWsswnK+bbEU/kgJ0M
7goNOq2hzcOqjd7R8uybNp7mbdUkK3CERCGrWp3n6dEtWQKqZ/cawETfzEAbGJqTYj+LFq9r7DXk
dNK0SE5vVDB7abWwsiElV965IdyBI0ykXL4++CtYw8EI/aZPLc7UEuo8KK1efSV+3eiIOpva2aUR
kEOItWneDn3bxt8KLZXSRMlEdpeNYovC9DBf+KTv+Wr8y1ZifrcP5hYaUbuQjByb57GQUttNzcC+
nMprouKhpxR/eRChscdybR4MXcJJvciQknM36NbvGFYFcADRz01OpExClR19BXGhdy3YJivcGxyb
Ob7v1BtcRkh1clJUZVFIK8wlBpEuY4xvyRtUQIBXCoixST8reD6IRwjhgtZOD45bDXTzG5voEmei
360Rpjon6zU+H1/3D151cQrANjwl8Ut+YWI5ZR0j9+gOEpVK/rmPSh9je3AvSi3xMMWmMir1I9Ul
qP+scfMTiL90jW7LXdzedG0dJF17axwzGr+ljTnHzsx4vU55cbQmoSDF3CuuXEyT8WdPA+smMyod
4soFbm155k0FxEYQXjvPAOrBfqHR81fvPWXAeKCsLJCWDaWWiQK8e7kmynAQB5EDyNFJk3vw255e
nhm053GZM5FGTatu/lDZZEcFSepl2A4xSLnRyBa4W+5uBzd5e33oTHuqmzS3qRXH6nsR4k5auHS7
Dtz8Z0QfwdnDyDd3AiYdsL+O3V06ph+v4A3Ka4AqPhFKjIxtUnzOvjpco6V09tcBYpAt89cfWcOE
LZw8UXaTrzCwPaZt5KbSapRr4iqGZy1IAXzZ7jWdvEN1nDkDUAlW8znmu6r9/vLA7fU/jJZtQnNp
IDJkIuDRaR7OimooC7H0lxWKZathwH8fUEQmqkRcxi+9I7SbmUrUA6FUgqMHOYkLiMaNcnatptoK
bsNVQgJyGYrINsryWi98URogpIJC8i39th2BtPdAUigqJOcEnmbbVoG96MBPimYC+er46+lXkKaW
rkKJ0HIkb4jm0a0MUmcFDdWSsnZUvPrRnP8Vqr4qj21bjPyFtxrBTPdEMF0rx8gr9/HbNMssqQcX
scfsmBAlryB6djFMg12D5G1ppuezFIm2zi8c1Rf8R9QQQEJbkFrH3taaM/xxrJ9WoV99Vf1qHFSm
mq7Gez74HvsCRiY908zZM7oiQ1F25pzvxpecgoEKLAcawCl4KI3RYydlec42tJii7JgZjNeBLrvV
Yh7PpsC+yOVeTeLOor371aLvGPJuxC0vhtb/Of1lvop1YHcHqjk0PTFempSKso7r9l/nNMn7XBOe
p6RHCIJVlo82mljcOYctDPl8UOOKVvtMqFgULzujeqA3xdOaf8Bl1jJoL55Kk1wIosqQ9DGV3HZY
bn+aJVOw8SayE1EuIF+ovVFOp5g1KqRAn8OGyY1vpSfn8Wi8QQDV1SF/DaxJuqcM159K8Z3g5OJL
EkDw342/4N3bwfhWxAUE7Rto/nfUipBtAKntPSP9dqHPh/MYYa33rpSoQjh0SP0dzJ1wbKfhPmyp
BzZ4QNtyFI838yOkFTIQffgS0tIEj/+mdE6of0cFsDmPcGNO0L4XOhtTSiohXeHcBI+KGLtSUQKX
jV/tauPTYLAXRLff6dbSvIblSSjTMrx2p/Vtd4j5/99+4c9ndFiv+2cQ0WkcBiJU3E6KgYTV9t0t
FD7bzKHQ6YKZh/g6QSJiHYJ3so73t5ykjMqjqTa+gn7PUwSues3XJ/7aquJMV/h31yAMFrHhswuS
QkGXjrOTEuanxMEvLfIEpm528iuhcJs5VVhg1ISbsJ8KkP6rrdKy2wh9a+suKWVmRjgjAvPFyHCM
hYTIaHV4d6tjb66Ahjz8VIBD0W4YQUArBXnoDO2ur7ItYGWdnrblZj5tTCdK6q/3mRLvn7hlhvQA
bjSfidYw7LlWxr6zTIgxF2jaHk0CNj6t6D7Ft28CS0CgueV2Zng5/sR1za65RyOJ42tvM1MZJSTz
OenwxQX4YCutukEMzuS7SRx9/4+nIRsMkeGXgGgQQFFrHcy+oPizk+RXxsFXJ5UoFttHwtgFbm+/
karaZePkSDDdAyiQOuuJgdVBlKij/IdTKwDdl1EMkFy9qCzPG4OaS4gOztX0PzDRPX6WoHmpnMd6
fvYYquD9qDuEFTiSxLWEbc/g6ZJXyME/fUL4p0yHcn8YLNXCeMW6clpJshseFF2BMYUbdTdDkDwp
/1CV/RW5CEHSPmZDpneJI8Ec8EL7yuCjfr1uhZ4TUb4phS8EfqW/kZ9AOr04Fj5KF2Ih+yiexo8q
U1zQYcUFQySEtDkpva2ZEAeeHM5S2l83ScmKKdRfxju7jDx3qTPMSg9wcOIGdCf3JTl/w6bq/43T
urllZCnwieHBOpLxzNb+irz5lK/9o6sg/RiparNGjTVm3RencCN35daMp8qcvuq1xlheyybB9sD6
jiRt0qEu1UVvUMjQsCZ4hfHZGJNVy9MJJGHQ38tCSSFw6Je022MUMqI/JPoDibcPmKc6OdD/zcVZ
6RG6st5Sui2QVoePzXOo75as41bIx2xm5GHsTTbVOU2vRRanYAyKyRKUpG3/5THLrm0wMoZj/i0G
wZY7+jmVsb8Yu4KGr9qqBFEMn8n1+2kWhivsvsg1cEe94JnFczeqNEI6Ea74QLkaYRR8yE91+WaO
guLpy0rmM62Po0Vp4s5ZUoKyYrFGtwUSePKnWnLGepz7Z46kPSql9EburEwcsCp9RR4NEiNoRLuo
I2BQg77Pc80Cw5XWzEX6D76SELc9efF04b5UeYssChQdXzHCq8+W+cYv0d0ufdCQASrxJnX4wL3P
9a8LBHIG1niotWG0rHOh5YOON68I29F7Ax18ngszYrrttI9oZ9FGgYlmTkypwcrTB7VzKUxZpvRO
iBY8F7iV7f4iw1r9fMneMUaefihERMajFAAtwVqHuzl88qWj+AERFkngks9mOiy5jAb23238eSlt
e8QyxJ3BXmPLFgNGXhrHDwsxD566g7ztnDY6NNu/wmAIAfxRU+u8nWmVlQewxWG/MyC7Nc9HMDtY
/n6IiSo5Fx5t4OxkUdm+O5uvqbS4eJlhwRqtmze9ZUkUAROgHFDnpyuK4w99LKCMiEWg0lKtnosz
GSs/fSsD4TwWMb3dwDNsz/MdN+8pHdR3n9wo/rA90qW62QEB5UaCpVKcEW7QuueCnt0f/4QIRa0Q
oCrjcwcdk0EE4Uidiq+G+qFZiujR+j5x6nXIEFi+qiga8b5Rl77+9VyNV8kiUZN8ijE3Vsw04KP4
T7VLz8mfeb8l0RSbcyYqd0osLoaoJiIRpNBaE8JRDwaikzyjkIyIYLMp2JeKAjqyhmNLveyTKO1y
LGc6P++HITV+dCHEM72BIVtf57EiU/XtSPg9qNpYlkZpGwwjT/JnXHqpf8rZ563woatpIzEOCRbw
KglRlIifTekGoTE9PVTCLVmLy8CH+PxflZ9t6n5g5UqauKha0gfxzN9B/wqzVQE1LGEY80E2Qu6g
qjO1JiXyOVKdFwNCaj5MwAckANwYTImtBNzxlmoFlQSDcl00YoYX5eUlNHMirf5H00I8OjuR2pK6
NGBM6247SbMXEodyKwiiK9WKaw7ihybtNz1Uo71YSzLX9c54Hncx0lmnroLyr+lNYfVTr610Alvm
L91u6b6eDouE6/D0xoQmujwqfiKQO00Qfb6fcO5OLPp7s/I7J3G/TzOUGF+SLFDtxAHL8nj35EfM
RLuetnbNkBYmnGeVNcMx3OYnEYCv9ZaIoTKThnD1mStJKusPvTPnjFZB5rXqTfRrAoeXVJEnqdwE
ncwIpJBVHDLGiJ8klpW+eNa3dbSnh3eIrBzwfauBTaNgFdIVEuY4Mu7lGYDn+IkYZv3UAKhauS9U
fWbVcCyVNNv5fL1OoPCF4YHliIc9XMpYmphGwB/z7UQIqvF9KPZ4XWVy5zQc6LVCu0+FuwaifdMP
8gLaVy5KpjsoMuQLd7LjOdohURZQMtbfi1F++zcUQzSezjKuaQX5zuiupckwbYQh6/65YW+S3sY/
pLQ8uivSl6fz9JgB4Mpn4BaUvJDHMu2beRy1c0KymyjUcEATPp2phl3MS/dF9xXEdVt9yDngqNY6
6ObKwJSzIBuLDRqYcD6VIKAo23ezFhTywv6dftHuhP21tpVtBnU4u9NveDL4L6Ag8bL5rn9m3K3c
mtOXjcGHEO1ySRBg/Hff+AUvGSzDA0hINonrFw2q1IUCHkV+8liB5m25vCdhkkxBcq+GdYM+FobT
4EUmnV40QfzX8yeC+UJOFyNjkdgCFCtiJWd0q0Oa4tvzP7YMcoWuTUd1U9TOKMaGT5WWSSfznBZr
LyVyvdvWn7/gZ2Ra6SA9T+jYtUIH+I/+Wk/Hj9wckk78M40aRabs88lJ1UKtiM2I0gHQwHpWGBUK
u2TLFyPjRsa7/LouBqBywcU6W1PnxL7WyULuUOLWak14Hw8+K6O3/FNwhhYDv7ZN6Y6Z/wGV9RUe
xc8atzc/Lp9u8d5Dt9BMU4hxquON2QZ1c0pHnwjUNCNgv1b7rE4+HPzc0tlL4eIf9p6Bdih/QzY7
EiDeRpo024A75qBmwwKIYshXDXzDxLZBSz/LJ33RGBXy7pKAbSc7W7gJauHxCBxF25/Co0/tM+kd
IjNBU0qbFYhxg3xydYSzDasLY/6iuW1bcAk8PQeHELxqqtFVX0HPAliqFQ5pozmKwRr9AK0BsanG
HOGlu4sIVMbx35zvi4MVd5qHwFpgSSMefMCbvWLJ/swHaCcZ/hHwCfU4Z8qG2FZ5kK++V47XMnya
dpRxFZLlfsPTCzyhZdzb5rTvsG+Pdf6VbqcpYZFmSeAB5VJM0+/JA2QIduhwnZyo/96haqKmlLva
/6Ro8e6jHjO1Xx6jmiK0A3+qspqqrEa6xF1ODJ7S8XLvfsqPVxKI1xbTVboL1bdP8nc/3/6mozo0
+fxT142wF2ZeUKd0UiOy9qca2CNlWXyu0kONKWfQxJBFOiulA2jeMfKnliXnnMs3FAXnIFONRJp+
vdAzhrPoe4NF8b1sG//cvt3w7lW+sHoIW/GZCyFpV17VLnImoPR46zG15SPg4hFaHTSdrRf+3hHN
B6y1N+/gKCy4URKcok0Et5zxasO0cvIQ0qrkvIy9OqgvtcNiszeZSY9hNFmghSrVPb0z2/1r1rAu
vsy0Z6mRsgI2O01ZNAoUWdV09k1UgkwuysJF0uUpCNuMKNWPFvpfW0JfBLLGlUz+jsJc0ue1u22L
TaSlyOY1tYfWuI/ItV1SqfwfIGRCX4reYe6Q/Vt0gw43pwO8VUmdLkyinxTZjMPtEhnzrQih0BM6
oBU0H88rSWdmfgC+UV8ZCNlxEBLhzW0KMskzRrrsJT+hyQJQXp0jAVMrGCptUUde1fMzMKF3tpSv
vAXONcQ6Cw/+p3jMJVD+xO+gH9f5UnWJ7h+dGsrXYiLpa9SR6zVfiv6kJqhN0yfPulJMjQcDnqDk
PNLPFaKOdwTGYlotDPoR0hu/4PeHwCFUnKhhu+gZ3tp9RwrMxiM1dxumUKsqbUfFCtWBcD7YgRg3
XNwYreVLT91dEcCMVhtUKwSEZkHfd6DU6Pc4GWRqUl7/pzpK85SP9g+1PAHZrMlQ5qdfXFCrRsDk
gzF4jqa+lAN4gxS9bXIg3T9bZS/Qr3ROYHU5RvNNnt2G9HC9r4ANo5AD3vJlJqWSdOuBvZ4iwtSK
Oys/CnqRMUrhNJp0xxPGNE7L9xPjLSD0AMiG0sO4gAWq2qmxrGAnyqqIavN5Ss84rMx6jA3nLYLZ
qqCnc1kcr+P/DXR3JG/tf8n54ADCtqKeII3nekDAAUxgUuoJBZNDWWfkeVBil1eNTZZxPjI4cwEm
0LeNsF0IM1BokMotnK84YfRi8bLcZvxmJ7ens1F6W8d4B2rJXo4at1xZ9nrHu6x6QEq3BNhTJXIq
1YX05fOnCakTeW8wnMDvMxE5VAck169SNepK+m0JnCLSgAPzSvOcJ3he/yLJuUGj/ivDgCIOlcFG
YUdby1WgqFGDiL+xO+LEkfE5jgatZAdYifB+lubZzVVDfACf2NtC6J98g9FOhc7HbBhY6c9rUegu
0F8ChwDhkhlSXdfWzJ3C2eU9nE0Mgo/AQ5yuR61MpRcNkd/fE9VtciJvEivE+PQDmqYPEwQ+0eGl
OrGhXQzmUXXi0AitZbGy67XHkLSB3QFWK30yPWfRNuqqqejT//HPR40Wiq/gPmXIQiY6tsnj4abF
TT2F9sLzCjOyZ+ffxYOgPgmIf8ZMGtfEoeJCn6A9fXaSaxKMW9m5GpqCka3OXzEWGt99m3RWMFK7
pJ4aWPKqECUMzq1MvwtzxrVey8ZYHxqiAcdSkxK48g4EwuuizCtm0CdxN37kO8O9YJefLRpXCYuj
JKra2BoMYtopw+e4mWHSsuwDIPLPzfhXZSqBm+Z05QBn3da0IrFLQxkd8rV2a8+UoU4R9tzacDVe
lPWYO7+ooseShLA7zwWu3S67HPOaPfzUe6qv78LPKOKapLCWKKv+tjHKiqw7SgFJPhhge9VQE1sI
u5RWfH40jKE3nXjIq44LaqpqG1MoPbQTT1I9CkUNjpFUXmwt1zcuOv9SEFiON2Z9Qb4/jBspbwNz
h9YNtbCV0QOh+1DQpeQBGTgwL79w/a8/nxbicZ/+iliMzfZgDUiSKs7cdV+HJpdjZq75Jjeum9hk
+mxFxYABfq9YfS7RA1HEkoN5glbsUjmdRggvuegYW6N81cUveLd6i11gGoRYKYrdqwMX/XsMF4bP
vXQuUSIM6ykJwgWLSr1Blzi2efsr3VI+28zTE34HyG5qW7vGqRM9qtimVleKMbglKcZkvxTC5FBb
vn9KyK+6nzPJksFry/KYym1iPYfrP+dDPgIpDMNf1DWrttZ+wFDimf7o7nzi3fOQMgcbUYk70XLD
HHKiQbxGhTqJjxoX2IjOsoHvAwsTVg1SbOzHFHOaIrh5WVlCQ+jmu4joH7KnWeoq9509B1McjoF3
GCHdeYNFVPXOUhDaZD2t/ONkQBlRyTMBYl0C1Q0k47yRv8wcRS4Psbi3ZlVDshQBaH01/bLYJ6NT
nQW9xiyTQDPSaiC9YbQT9e14832TsbfYCTrjpWapRyu5PrLh8QbejMzhaqqKPBp4xGLMc5/mty5J
m6Z5O5Zo4hRM9bsmXyO5sPO8UmRFNAmuamwuQx9tHjJJw1he1C8SO6HzyF8/xgKWj8R8C9HTkUWQ
+XDX9lWmj8VL0db6XFCRusQKLk6DcWsEgAzAjopPfdcAAsLOr4EWXjM1/Vw6yXsUKyDdU4hs88K+
4W6ZfAOgqY+oldG29aatMdePhvsDJzhS5vfd5jjxCyc2QyeJnLZBMG9gvvcUc1ZwQT/whH4kEiet
VwDbICP7nSfM0oIylScV3YDkkXjPIohWtDsJiNPEvZY3mYRUjEM5XXI9J7qssKJqeN46XjoTTJRW
yKvgEG38rAiKHE7IAtaJozlI+C0B2+TQF+VgJ3NZtBmxhgAj7cVfibKupUsC7MAsnS2A3f9lu0pl
z+DI9cn+z21SC1b0cJBBXpuEeNbVT8pviXg4me2+mDHuNLkjUBfrALjHWtjVqQ/cGmQGA0V/5+Mu
eHEqNnvrcgwLCJK9Cp/hjYxv+5zox66tW8/wTdmEmaVN13gjRncldqytTOYulAtqqaEw/aT6/NF2
P/JtuO/Yt/c82deM+aWNCDP1w9O+LXtnOxgHeKd72IbBkGkDN1sFBMu71KanwbsTUe16paTOZgxr
xpd2NMD+Y6PvGqNAyzHoDERFiSf9jIA/w7FUreigILmkzzbySWrP9Kj1rr35fJtHzN8rtzCwuGzC
o0EaTS3TQ/unzhH9R2kg20aJPfxaEjJ2xIoNI5/aXO3Fm5jVxgG0rwDK1ZtCVd1S3iwEcMgaalW1
ndCIlTUO0/qrDDVV+lv/1BNflsouqEeHRyUo+9FWGJh/XoeNJPutmSHCDUfn0mWTNcDqgc77EqMm
4eiSqZ/ULQkXyAzuRPUl13rYlGhvJIEcEAGGrjHcpXVTwf8PlJQmk5jA5I38mIc1EXzHk7DQHYKo
qRA1W3f+hF3GUcU964eNoB+oJLCpmdFtfTwXTIr5+eBi2VV06qcZMbCgWIwpf8q1dn1djwIBOq5X
zC78iQ8Pd78fP+nZOsxqCsAzhi3ez8GqntBjWZ3sykESEjW+oxHTFxFVRrmNY+6l139YpyqPAUH2
DVT6ybwpo5PC1h0aEf1WBBditJe8IKK2JaHT3xISbKlT4yQyvP4NPHNbicuSetsQH4eZyOAXg6T0
yEZ++jtt9P9uooV9iHb7vFaCVSDAG0SaJpglcPK78Jcd4EQRHnNQe5a5QysWsBPP7DCT1gWSN49S
GvXiX/0fWEvJk4Bw3o70wn4EJhAm6IAUeQz/9XelDzSFJunTlhE5rFl/KZou4vJMdWVPqhckxOoL
Nh+1oF+o4hoePeJeqzTw0XDTcHyYi8BZMIitv8GG/X71fXDfixLDEllgc9/rMgGeD0s3Yobo9tWY
eMlMhjC++FKZsQ2FHr7A8MxjNJnDObpXcgWRxDl7tTRH4Mn/bQDLHYMTYJIwyTeeLDgaJFAkOkoy
Ep0MH/1jo6JTdWJNWweEL+0KhmzjKjY9tWzJ86xxs+K4SzRjRquUCDGKJZjlP/ikqZL5jO88IYfj
YP3OpprcMtIAGvZxJ/DvP4gU0QUCuU9NAYhDq/URJ2ONJe+Qv31P6P+PTmhCx7UN0RxSo7mj026Z
FKgs70oFqKZxS1twUsVDo0c/l/80zd8bcL/t9z4G7j3pMFOJzBmt7uRmbox0fmZcOurMalcc7nl0
kKr4fO6eHSG3caT90IVD6gCMW8gYM9c5MUhDvZfCMJaPtN64kJvkhAzqQQIV6gq2jSuYGagJzkR/
cKPGTQI8IZhMHGYkgtx6Bd9lIxUsLDiyUAqhmmzVVoaDH47650s/snZBWPV92FFZlW6suJNjZhYW
dJgvvb1zC6X5IvG5LaAIukJRBWDudsIZ8nBTnLoZbuoTb0jDHc+R/DGb6aMhuqU733T4hrWyX9zr
wGpIFK2fEM6mpuuE0pQjr9FytPlgXQpJyfpmNoJBrfg5nVs+ME4ACcsNDxPJS6bvuQj4ESfRuSCV
2yOgrrMhhTd0PUVTPcKajPB7qHrOgwECJEOxvj+H3rpriAnN6XyLZ0blD2EO/hMr9m82Ay/QQUmr
ERJxzF5kSODnezk/TwJNI/Rf3sIx8wQPRDSi6h4dupykSu9io1nLdF83TwRyQ5ftY/eM+IAPhl/V
rsWiJHZLABrFuHLEJiRBbmbdKeUv4OsuosM5D3OAUq+NxXwkaTccXN2XprzQa9dL/6FOBWcSbSk+
nhOn9zw8Z511m3kffRqqNc2Nrlw1tAQKoWlqserXCRflCbpkFiI3hgC9MTw3sIcZLBVsL78hLwzh
cff0szd22W0FMhJVqElZlGEkt2hjY8yKMsj1roKpdidI9s+p1NgHaXN2hERf19OSiQQqwXIAmmfC
I7Oyik+6jt2E2WmEApfkCv12AJKqFIlI1GXvJuNKJPf8jlfzgYiYOpMXwsRc5YDf8BePRpAicpPY
Zyilq7bqV5BS5Ia0VoAzKGdpM0a2FAhT+Qn7q6AWyixs7uH7hjxBJaN9FRjYHIZJ1yvPNYhMTzH7
y71/Zpd4XeLTdj3o4rLeNj56JtYdQHPx/p93rkWGSyXKsnuL+VQadAv85aS9aNp8IOwcRcVSL2tP
a8n0mUrhtemB23Nhf5jA9EGgdbUt+ygzNOXjL3eX/C0h4sPvaTpRmEgBXev5LsKJVu318KtF4mLY
PQLneyNzDqfgUfRVZdyh3BB5CPj3UDHwBOMv1yTs7XoHnW6kxjp5yBBiHlmr4WWrI6IyDtckiy+6
eXkJeqH8ni1Jjw9rgfRUUMmKvMr0l4A9co6Ioa7rqNMq8gh4zfNC0Rz5DMEqB/hw78ALO9k05dr9
h0V5zH4E9W2u6HjycJQA9At8EaciShDdE60RlYsU8GMAM5TVAHRs15A/LROWlVpB6WsJsbsODN5n
UL6JvZ4Cv4Qo+GW1vywyHfHmKpA7rEqQKEQSR5JSnNxSDyQTwNJcGyX52KXbXnmxBplzEqpyfQFu
YvvC20GF8cR6Zd2FNTqMl+rcOyq8ZtmUMB4AtYgdQ+JFl/0poWNXucC4YoQs50CwKhj7M/d3JQYx
QuIzjsu+Vd2bHsJFZdMcXw/NrOiBoTHbcP9QDuEtdss2VQRR2F+NTAT5BpqaMR5L/IuuxACfp8nB
u628qTbFKnneOnE5hdhXDhI9tsZpwvxo7VoK5S45+eJlnw2Ny3eDodpu7fhu254VluD9bFNJStIG
zfvHu61xCmQlz9taR8h2W1sDquQuhalxu8/jZ9cY0ec50H5p+c5PCUxdWOW/2cFXRUK6/mN0CgeX
BNjmUEqJB2ma6VXLuOUdhPOgtFUBryiY6idADDV6Vu69OvBIB9++xUo8+BjSZIgm/3in78h9HSny
O9PUgjz9nSc9YSF/6cpZP7+Zq7qdiL1hhCoxW704S0pi3nbnxW9/QonHhzRDLm2qMKYEXjb6gGmE
2V13B61EKqetALkCVdPtquTh5xyC1DGn7bG97E74nFb6VyWKKoE4mys65PHC8wFvTFby+YnIA8px
6+ImjTgHdPUHYT/KkqbZ+usBP1mORDgn1F0ZLf4DtY6Gv5rICC6gu1MV9b16Trdy8TS+/1dstJPU
ki94mDRfx8kdBtkwPSldQAPRiGWbtcqiEXqxqm4iOMbz356KBI14mSTWQcTH757paiZzBGMobBn8
xVbMh0ARsnXRU8mQT78v819xKujF7ufZuuXYsVJ2Y45/OjGj7+lYttbJ4eRaCccPHMbYg+wSZOH0
7FVqgjNnM3C5T/0p8fkNy0LH4zw9JsJJG/uYJcXiqZrSibgX58Ub72PUL0ysquI38pq+xBcJ9UVX
AVHgMtkeJ1Sx9GxoLGHm8aQMto+Ra5jtP/2VkzE5eIUuNgK+e1mdmKWLiT7KpbObS/a/NtVzcnMX
TJa4DZv3LTDdFCj6BlhZXkMofq+MSZpRA/akT6s1XDu0VYd/R2BDU7ZuCltISx158/xAqVWls9I1
myDldrTZRIIhvT7tS1wv3ym8wSjtdU7+yUjoObqQw+VpjMs5zwNZamFYCkj0tHn4kjF1gHcBolgQ
J+RC0bv/adgx85Xc7/5l0xLLxhhN+QzKCQzIdGC0rJ91eADF88NmmfnJj7SWAzxP2sBm279m7E5x
3vknj3YCSPJAoMK54myi5N9UDu+/Ex4CC561ityxUvgJUZLjbqpZ1ZCohQHlPc5KRjRAU3PsE5H5
FtT9kpl2AmFBBGtR5Ug68wQmgVPlghXXvibvKEwU9ALerrfI9VHOhTHPDAob+74MePPJj9Xjxe2p
XUlzMSMYQNzSGVbrcr/z6RZOFrLPHzlvehyDMl2h+X8qJ7MuM4gSNCWqqqaI+8P2H52kFLSnfB3f
qYicr5Kn6GNh4FroPY9N9rAM8QM291gMICtK21woQ2nqxBoUmUgPXqhIIincUfc98y7I661M3vx3
PgjoB+rnd3fawK3MJQRmlPEVwu4wcyEY/XYg49jwO+RA7aotQil7FjTXefZ0St9x86pLQQVeh132
0SV6CLXCq7wa+obZr+PQHoQ1WKlO9waRLQ0OETw3g2ZrDm6EdTUBzht7BTlUzZt+uUGnrqjX0d4B
7zzvSjRDIW3KKlDwAKPEP1z8lUdhGKaBdjU4jOai+qX7AQirO0oI+pGUuMPwkowQ/SZbGipCdtrd
v3kGDXNDUcWCg/YoOGdWgCyye4sOrM7zDT7Mvw5BX/25d5gKie01Uzo5gR2PFbfNFFEB9QvGttnb
dWHpSnjsFmOG449QETlo9RgAn3cTQmynmCRI2XP9/QfqqglH29iUnIDLyNMM6dSq1CM4PN0fkyEG
GGQ8vJn0mKY7Q60H6d3RVt8lvml7jTjvFbMOPQvl9DDRHH3bzy1Ji/b/ka5qciy2P0q+U/1OieRz
R4tPjxyUSkA5JuIKCrm1hDmaxDuTwz4D30LL6TloCVjWNPkEgn44bbGUKEvJ0I5HuK7vPlsJQoMC
a0fg0oGJnHcLwnqtZL6fo9zmThrYE6hfRhCl80JvKHjM2XGSG/lJDlIDCxuLzpaGmYSRSadFmUr4
JxARPTiEZKAInGiCNKnUX3j9r6rJ8TJis8zRkClGdLlJSr6EQV0aGgqZpQZAcII4rPR0VApnqiam
JgiIs/ZAaGUNBQW8CsnDQkSZuseOa3Hx94T4c0d8GvEfIjYRr60Bt5t8LnsF5Aj3jA6E+4AOtR8k
9DZAzPu7/84EcqBZMfJRz8Rn54/5IrDVJ5mwtyZhCSuiDgNezCVYeLrCrAyPJ1zGp2bYCauyXfij
blORVORy4Q7Qc0BebymUi6zOM4UJnj4NOnG/B2tbCm9s00UrSN1mT81dtjwT+S3/vDNaextkx5Le
9PQnLlmCQiVEaeX1GbdNYR5EZHHeFBb+MXVWYwbjV/kVJgfWccD4TNQbHUmP3ue3cmbx+fyoh6Ts
/U2GuTpMDAeE7zRfdhDn0fud3OHfmxTiomORpCYyYnIk29H5q63uo5KJyXIAeO3z+q6qSk1MMX3v
kLtWsFNzMjsFMfZXzpT3f0xjT2CE9aRyMfizC0i0pE8IufnVY87jHMQiZyYdOeADtKHwAkEGLUIq
BilPzYGPjLCeDQf9/VSDnNIHINxtOeUrxZan93F9/YMGRV36lkSeBrf4Xd1cScWgFrC5JqOuTOOm
n64YnY0UwesyjHAO6sqZYoTv0LP5tRgT5mElT/LIXqsx5A4BNJb8D9Iigi5nF2JuqSDb2KRpooAc
tZV2S6LOAqoJyqDr5CZ4vLib0L2FdpWu729X36Vs+z3WhvRjtlBubGEZWOk4gzOPIcMLMFqS0NWh
eEk/G3I0VgqM7PE636IOsUYEHXP8xHXpkYUYvWP4+7Nu8y4RzyLP9pbnqRTgtaUs6I2v4Ev/TU6c
y8HYtdxl+xOX+g/3bX3mmtE9H5wt7VfGfTbd33SAJLElsSENM28gSLkacyGYfWmM2Hh3FknU6S4D
uYg/QhW9roKDiep72TEweCT+EH3shE5pPuDVsHY/R3eAuZr5ZKPgX6fEspGv+dN7/q7+ZZeY+3OC
Ly9HRyZmnc8/FlK6GzbYsy2U2erQtl6st1Xqm0qKfGrSIsszrhFIFVmez4EcAVklzeMtYXfckqy7
VZWUAeQKRQlI0gyJYTHTyIvUQwUpPhmPopEXdU/3yHATZqOSuVscx+pWtBG8EmTnYut+pa8Xs8us
3IHZQpIl0nQX4hcKGQOGieoeruLxjJoVKH+IKE/PqLe/Yk6NxS0kg0lrtPA6hEmsvfRnhLe3Vq/F
LGq7D8dd6TUmxwFy6Kc0/fvq0TI38RhmauU90m17iftX/xXqMHpvi2m6Oo6YXllwdyzkmOoeeX6f
tc0W/sCS9F4QBmkWu0FX9GyLfXLjC4/fINXROcHSrEanVsTGCD/lJW21VBzOBcUnQE5F3NEF2cQ3
RvFMx2IHCAd9ShMwp+otCPZHttnsErJLJ6ezu6lNBNTwW1C6iGRu62wyDqPinLPUfU4jD3hgCN7Z
mpbaOKSlTWle1Mr6MAcz0q9jKpd+8L7Xm23OAuskMcfmQ3OTXU60IE/jmv5QBpDLz939Kx3KdcGj
e7hkxzrEvGrZVmKsjteaRNJy5CrTgC3TMGPsCdEtpDefNMOXlhA2hfuLrcYMXvegNoBzGlawVnB+
9OsibPIk+6yQ0sajgHaHwYjhM6AhJ2z7MvWyXqM2f20dkMgVEjL1wnM0okkiSWVXZaiyeSk2sxeB
OKwF94FSpFb0VA/WEY2NML/TdFbE4Gqzdniw0NMS7NrgQvxvJvfNMhhTpxZsi8mDAkbMMWwQEyOW
D73BH1NgY9XrP5KtlO5qLJH6YdHLPYdwzxALlZ+3CYl5XSFWciUB6k4iROdhzDGLIkNLSN2QnibD
b1G0B6hxZsj0ZKO8M4zrGKfN6Kx/Md+cZpBylNwCgJNy4a2UJ/UaeVtgZp7ZTAzgwZ9kYCyWLNV3
T+QeRepSlDu/w8fmUFwvPYZTpqFxBYU2BDHtAvgSTfFqgcENoCaGg17Zk7KV2+ttvzBNMjXNar1k
GPw+GUgnB80bms3LWqbzimV845cWju91UHPHgXeqQFVVEj7dv+tVKUiMVoQtXa9P5rpi6D3LQ8or
JefdoL4l7pS5fVP1WHZ0NVnFySkab75vwSN3cVcd2LiCEpMkJaj+vp9odndN7SaaxjYV++osnXE4
WN/TJOSLhx66mVVgQ5BYt0ka3Ms5BVSURDEcGjLKazngKjOr9lDFNlIGhodKZsbkkoHnF4R1ZTEr
COtJeCvzKzQLHGOqExcd+CZzSUbZU6ZUokPOPN1yqPQhiqFRHtEVvZjFzOBsD44DvMO51zA3SUHl
ru4y7fafZuMbfc87hi8KqGFrxLv0yFcgmY36uVb8lXnNa1Lbo91JU+5A/eAd7cV0iPZnb4lN3MUr
OQ4hs8k7BpaF/vEJRxleOc0OnCY89SvZ26VuJ9SNU8tOhoXt32DGHUzWASDOyeB/O/bp91qa4riL
ip+iDsgPkiPvrUad8vGxn2bJtt31fiVXPjEIer8ronpKeWS64nLxqJnZ7/ReqmtPIJx+ppAunhus
YZFUJeDkD8dY3e0Qn9ZVyMOpfM3LV1Ek/gg0ZviJCPPv/1peooM/I3JfygSYbbMjaHN604G62oS9
b2a6Nx+aMVRGiwA/ZzXe0qZXdhWXNC5WCUitRQJcPBkpEq1Rzs9+v/DBuyWm7sdADpJpWTTN5vAR
Rla8LvZwkzPS4/pWNfiG1llwTY+Pgro5wONmwP4tapprOcR5a0xyy5YftVuYjGxBC+lBZ2O5vqfF
Qsck7TzwsqoywCVVgzpppZkgPJFLtW0zgmiGAm4BEZGk1aq10JRckyqD/0cpuq1VaZPbYM+3WKre
06sVUfllMkcibJihWPmLB65CHxz/QurtdxVM4HalhYY404P2SGrEOew9AUNMtl9+ywD/Qf1otYMq
YQf6xSbAv1L3nDq8+/cajatVnDhHpUY+v2ym2dZ5Xe6yOmecapJCSdl22gBp9Q4KWudblOogXi+k
CtRhUJ8mb2kpdJ058WBNMRaGsYssIY26ZCVkMHt++9Ohub+WtqvScXtEqXBoW3Bi5VpxsgSjtxwf
cElzhjGWzE9x40uU7iCFW3sTmsBraYSNPPeM/JOL37y0Evj7fqZ1sUDx2cvj0MQmgBko8anxW0PZ
bwPMpJTRuOLf7WyGiTBlhSFOO40So1CGP0I46HUPs/qto400665V/+3H4aJybG3b0vC4RZz9w8+o
JkwvWTepLrmEKYc3nwEl5aXXLiA7/LCaPBay9EK+E0CT9nNiIJN2UMl1XSpwOUp5tiwevCQ0Xqyr
791qwfCrjqVFe1UHPSSx7bU5OWbbLZNxDl8uLLh3UEcfh1Jg/1fFtIc/rNcWiC4ffGSkEIdI8Fal
GZtzB5mjVQ28vB+gkCIbPonutLWNmh3UVXrdfKSOSZIT25zIBn8BYoBOk/DmbXTqj5I66wUfq7d3
N6HAhWWBWJ5Kf4oy8usPu7acqqB92dXrBWwkfnxj4mCLt6qOQZVI5et+o8M24JKhoXD053NptCwi
8NrCjEfI7DW7COHhW4o9x4/V5RcPhSp1GEaiACF1G7WDhh8jPNFCzWaCqqqozLFoyr+65YyPsTtU
2CNZSh6O0/8GfUUbZoSs4SQzWyWg2UlXO+Wopextl8P09TaHhgIS9D+4aovIC4wIPXqEzV6hDvoZ
XgE1echm69sBq2BUbjaL7Jxxg+caWShQckoSHYZQiBap4zygaBnJlgWTCTdTljVIkNaqnGM+G1F7
0bNL65Pap+cL+BPKKbMRg0+GiBZVpCTjnSqBVXTYtACIwmFfb9gvoXzt4YqpD1vTFfsme6n/uBCQ
t2vI7uKouLdOXW7Q7vTfXA5ZSQrmdfrATO2G3wm4YnnAnw6qeug7AT7TYsRDfGFtFBPBvSNxsE9D
PKGMl76j7wTO9j1mYgKIcpnk8v5h1rkEsWVm8mTCQ5Y5zNne1PwfFE0vTk8ASlHyusECbCvyIe03
ApqDZSnFOXp1GPX3UnXg4o70fc8TX9uO7ZoazU7Nxu41dZa1KXRU2S+OsKSS23lU+sd2Y95lbR30
2F9PNWH/7bkKo+sqtZhqA2Ub7TQRoyTkba75N/NmE0vjxn/1tJXrDAxkpQZuv+HEmLrSMBNFKyox
8IxBQb+RsJK4O1YN/rkxAXgV1ae2Iw+sbM/zmxwNVCIzXxtPPIsMxYf//z7AaTRMWF/sCIB037XM
IteN1iN+YK1vlEtva2xjIHrwzBZxu2cSsc+BetJEhvg6Nm2v8MXTIkMFqEkJCHAuaw1Uq6SYjcvL
Kw8qUiHdYKSRELQdNpwZEWIGQij+b/kigI4WIF6/oSfa+D9CdZsglIja4VaIW3qp027lr6e9PFyC
UhoTWtzXymTObeZGmyoHXqBteS3PQuc526+Nj7XTNcdr3lnmJzduNyisuLDli9rEeOIBokM17Q5w
KxxOWAsX2zE6ZNG/iGCLFe0QySZcvwMluq6O/GYwfGGljwsU7pimX2LnqTVUhNFmc83X+qjn3+Pa
5RL/T/QeI+vdoQ3vKdt5NI1RqZnie6PvxTUSXeZyLmAaTStzuvzTSaMEqzNqlDsOgBnD4wPfC70y
wKNThQ/H3+/1HVPbgvii6MxaJhaxEE9LfJ1a+4NYxzoArs7Yi+vFJcT8FbQRxeel+yQIoo+c50Ik
jmCUfyfmuYmJqSFTqF56ioKRpGGplo2/iKOjlZsWmYBcZQRxhHbuzwABQhvTtHhfyBLJUsqivjwK
fP4zj1nPEMAb1tEbCnOqg41UAys6ZnkZXw+DUC7Tg7jLZQaRI46t8FKVuZfNTOwUGp8+1ooWXmgA
JLCy6RBx0CiGrkcstq0HiOOHSP/1k+x10kFb0icYUqkQxM2qgaIHqGe82nia+SzH7DqM3f5vL8uT
hzPDjRzPmv+q3fFe9oRAPkgRTNbc2PN+S9cuaVdcqCI+62jy4iAjIW+BcmDT9uMerb3rWgWORCjX
4Sp4KX6LGcwiEhwgsoy4XHgN0mwrvbz+3+EJocA71OEe0TdvIUNLVtf0NG6UxU1vHACwyKWIgoC6
lLZ8sP+sHHdSvFAaenkGLAvARx1XfYWNxiZcAuMdHLsMUpy+w9QU4fe26+NPi0hZTvVgBmQa6rPk
glHDBrxO4wW3jTsGopiu/8cxkXs9CJPrJxqYhoBqZpYO7gSWFYcQOaNR4yXD/G8hAs+PaZn8Euo6
oQ/CvjvnDjsotyv+SMf1lw3zk7Jj6XnaQvx3yxoafkEAdmWXvateTF6OvVy0m+S2Izg0W07To3Fm
ARv4lNqjmRZX36/WGp+nas72U4XEEK4X6vxeDZtXZ6dnWjCsu4SuSjgG7svquykM30SofJFAIWy9
yQr4woqdiQ3+niRi9nYo8lz/M3hdWGdaNY1WPR5KDnFAZpwg8OUj+390PaSNIvM06D9qs7lhUuE7
qWd7ymV7x35gqRqQV8TUZnFzdZOrTwO45P0rBN7Mb+Lmo5dPAyjjLl4vWMPG6K9cO01JP93loGu4
6rCotVvlU4+B8rY+IPVcJTe5QqkGcofuDazjaup5z23W3+o83lW63wD4IelQ+2HLY/8QRLn9sZOd
nXM+9bHJr1hzK0HA2LPb/73UsT9iaI0QSd0emCbLIZXHLzWxSmnmqtGTD2qgiu34yh4L7MwjI59q
B0oaLATC57NJfJzDlmYVofa+kxB00DWRnkPJX7fsT3jMLarUFtTyPQgCYIj6SyqsKJxWF81+JJei
1vshatlR+AaLlVh55g/Me6TzgfgIxjuaOaDtp/RxhMfccdt7aN28VMg5vu8eqka51Ylo3XZ9nOnv
HnhHAHZYw3OWLzH27UECQAHXhF6lnAN4XQZZfP/g24lqDw7GVb3xvKNnTI8e2QVk1aPlGE7vtAan
jeuaPYLKq2bunSST0eIUfU+DMaOG3gDM2r+vz80Jmd/MZsruZIopbDdctFMt5HqkFQUPC3TpCv9e
biWhI8jD1h+7SnkYorLia/Wkm+Db8rLPHHT1tAfM0wGp0h2SV9el9Z017TBE9NxbLtbg0+fYWKb0
d8yeevbkcxEPUNto7LGv97x5/2fYNr1Mk/yeltCItOwZPGkr9NAVFKvzrwGnKp2emBnBn4IUCmTC
dtqgy3iYe8UeglK5tuUIfqIGij4dsZAaFTICDsp+sftfmBywtIZszvltCsQ0PUcizfG63+oFYGHa
zbaZ2sF8GbdJWR4fsKJ6Jef7vh2eBJtVj6gKr9hX4zU5uNZiACdUO/d+3G0Y7ajFxc2a6ggEPWa2
4PTjENUOLHltpzJLx98Q2c3hllhvISKfEczTU2iNE/+cQtr9oITmv5ZI9nZixvo6wr+DGJMgfgP/
yHwf7SjXSP2kaSpBHkSelbsSLkoqPf//L+pzJqWkqnh00VCYuWUsTdr6bB5LQPkxcFSFBrTntnMx
nkkPkYo/Qu+svEAiSLyYVBwEftySIMwU2QI9RoMk58P4xCkXwQ7NWL8q3eJmMBkd4Cfc/3pbBR8z
TkYXv/lBXDv4vuYn7tIOE//loOlYsKfYq7/VxaTD2wAZCXqyo+4BDC2icWsn3DAos1NedvS+j3Vq
CszdhVOxT9P4+1ETJGrnxgcq80cbVIibnaf6RbJCnCMUMG+dv+JeqSPdmhXjCrMUWMPYVEGnytjj
BisqZH3MmFIuyGqwzMfaEwoChNtwjDu7lNc3Iy85C0xiHrKWELYxesROI2RfOsvderLOLhi0t/fm
dg+KcLW+9FgYqm3HdRaXjWK0eFeaWrVDHLKh9jlrNLfHtaRtcLqszhcmhMTWum2ZRUsxbKcFvojH
E9XDb9bvce+YgzpEnXnAbwLfF+tx6gZt+wJoBh0eIu+BADPNvHvqKfI6/n0l6PSvBQLRa48uXqM4
3zm41WNeMgO6g1x46klVF/keNJVN3PkrXGyBiGRanifxHZvyf6ARUAwcNMhgpYGIzNGqgdTQX/ZX
zHoQVQ/xfriniwAzdueVV2s4xTKylT8gky8ER2gnbuZ0PMiFzNO7l6OWztZ2R1pocCK0Gkc+/W42
oP6aU6deE0zg/Ka1xuBBoVIDMS8aPmqqJWRBO6RQ33rHUzl8iWGEruEiR3hvR9++u8QxSc+kuv/2
BXwb+QwNwmmS0dk9Kp+v5AV2HJmYZZogof06YBXg02fc+ZnMJIQEg6CXiy7wuDhrlnQNlJRS9YgD
Kq8oPsee6oODateOgRLpAApUW/EKpG40tIMFQTgA4z77Sb2kThF9U2XrRI2+nnxbuKaAzdaZX2jT
9P1jZKdRjk8eOzOtHvi+W4I2EEmK56+HJMPE7tkRn4j0JXq04u2swXz6OLOKBEizFudzybPaGRTJ
41FEXb5Ln/ZtHAlQWrOJqxRtf8gahyTLChyQTcsch4WGsbNGuCqLiCGkac9PDxzEfNzS4baEvAqt
UOIEF+4K44X7+0f59KEUpSI+2loZBpiFqktxB/bOguEDWVR44UNVl/qbXPmgN20FQzwP5w39e4oA
IHe/3s2l2fSxQ64XCW8yfpIv9FD9VlUc6Aj3zw2pzCErfxCtrgQcRpYd+j8IDxNUZEQnOfrjqF0d
p28rPjK90Rg5iqL0WhWVXFuX3uEAZ65k9Wef2vi1+Hh/r+kQTQ9WQl+oZzL7Xl6+yl2epTajPNUj
MjwGwG1uNPvxI/kQ6JDcDpU2XR5LkpKhDcG8A7N7iy69XulffDEJkhvFewvtZHUm+2+8EOXZ3rnx
lo6TA/5n/3w/PxsZtmr4WvepI+ZU8IUKRxTjwN5sdR0KVUx73CUYpQw2EpICKBvQu2U4GceC8NKt
UVMjfiOCfE8vmM/gTMrJz+1OJZVLjnnqlZpm2iPDfDYOLjJJ3Hfh4zWnzerEKvVLlT7DetcaQuyy
9hMKMNJvSkuBvPGQaxR5u8YLB9+vxOFQ1qyb4QyjzY1tyDHaLYRBbnopdnYcxMDjq5lJLzdN8SkO
/dOCqTTivMquo60WntQ69CkSVnHD4Xlyw/TcB7PTX1J5+QGjon6GfkYMSMuUeSpqd+NMEQssXB5W
yx3HdVRJojYij7wuEQqK4z0xBC6khgNTfIdjEKSkkqW+kCe3ZIh8iEPzvunA2BldGJM1SdoUTcNt
BDwOtrWp6GZW1mjHDseHZzqbEwh+0DBP/pz5uHumwXxuCbOw3ekgMl5kt4WfpDNDrSRU9T4W0mgb
LxUa9fmfF5kpKnfd2mdBisNu75o3wzIx9bqq1rOmA97li8ROeDWUrdSkfMOXVyimqFZuu+Fe/ZbR
Y2KGIgPwmHIpIQYgXtyn0lwVcd8BsI4JI32p3KVyf+w8pSqDJ1uBjuGioff0oFkdQwUOqr3hGbvX
a6ZFC0GnsGMP6vwOeIBBXGWEksMF5U6VbjKHkubp/WKNEoYTMsn9IHQ+TbBqtgDOlVKm+uoYK+cd
TMmNlm8AM0pB5dKlQF8K4pf0I0WAxjJ4K8HDtKSh3bp8/PpHa+yjlxS2uqRENwK9hbybPtCsDg59
NpijZIh0/UwoMON72tMZ0/IHrDnvEDy3F5wICmV4Ei78xZBVJp3+I//We52Irjw8XeujbWifjKOK
hGlBWTbJ9lQi0LvFJ1wBUAdPalEEgg8hAbQQ6Z9jicYQv9GNIcpD6KTXhfv2f0kyC4a8JwoVWuQM
dqMPVG0nfFl1CVQOsUmwUujwVMal5UyMe49QhXGWDwbnmJb84eICeALMqQ6Z9hEfqS2NyXpC4RzP
Upu1enpfEs3higAHL1ZOXvgCr+Fab0J020gzx0Cq6JqhXy+sqYi36h5uIhFtBhggZ2AGryB5DYcr
xB4KZRLzo7aUyZb5SxMLGwhAO75OuLvBxMG5xNNuOdmu6EXnrbJur462YtF9Ch58S3jIw0Esr36y
nlNBe2KDPmI2MKa0X9XDkAyIv4IN1OWGgtJIfQDziFvqxJ+JJFLgaou48D89HoWg+R/5JPSakf4z
XYCSGz29N/xmiZqta6OGqmk1XjkcPdDok3sNp6RQhW1iWTq9mpC+J9+o1wjswCrQqFdOxh7ysRRB
+aCEBstCQ5XMJj22Npwtm3dIXRUt+0YprWp3ft6/B0Gt5KEOiL3h3srLTkhXEsBjZsSF72ZuYxM0
PpnyDAUrqkyNOYjtT0prL3rL5LxUgm7n0FtvnZ9p/z0s52mcW9HCOm9YY2vyl+OS/ORNxO9YHZFe
wvH00jjK5FmHxTMf/azDYPAjjk5nZWStK+VWuOtGtfcj80WkQnhjIvb/Mh2Lu1J4uEQ8eFzKrPru
+O5qHCowPYf4Zah99S/0RGnY0999Pla6yg7J9LZATZ9r1M3vD4kxG/QnDJMmSP09wkPdbYe4Y2WS
0sUGAbLjwC2kCsORqeOb4UsU8ti8rg7PWivgO/AQrscwocCH/BU9f0K9S5u2nqlPEZ6uuQQKLUV5
/6BdnEaXIQ4DMYLAByBcg5Oh9UciCYxkfUorNMlFrZota2UbSmnxgGsnjgdlWw0LI4B44JwFrQbE
w6fXWgBLFAjG1AKTDi70fNFgpV7T8BeCNLGDJtfPCWNCUnPlpTJ4VXmQLiM25biWX9JQyhQzm3ie
TjbuJ4BuupeG8N9JXMIqsGlAzoPnSqZrTby609PYGJVT4vsdZ6NfhdWdT6X5zDBhGY0yTWpN5C6R
0XrwZx4huGhS57MmqIq5/5ZZXvRICTTeh2L9praAUc0BKEHPw2ZyfXkhldWZG7cQitoYsjKn0rKO
kVTzaIQ3+KNeskacIMAOU+tp1z7NyLlkazg8dgkH1ySs/kYZQBy5tcU+YycNjKuhlY0mroym0Coz
Nb+tul1yP2G/RdyLj29V9qT74tnys8VJp0efo0LxqrMT8INzlKefPyDUxOg81SoQ4SsA1HBty8HP
KBurSqbhDADoRU0Xs5d8nYLerfN4XijoDsqhX5tBMPZNE0fmTycHj3ZYxpc/XdQPEWod5PF7jKa2
/SeqybK4C1huy8/ob6JpvG3X0R1zWmad+593bMp+ZwD5DRrS/IZufACHR/HS1fdunM2heNZb/AaO
9iggsZpLqW1UJaIt3vl1qqcTDcflst7nDNiKxw1Xt02A1zVLlRYwlasXKvl5euTLFB/zl2fYErzs
80RUrWa7mfEme6HZqd2IqcC7MOmLTnEnhwAODVJChZWYgH7K4Gvfzi1JkJUAzcxwExFNKjRm5Es1
m5RjVG19ECoocbyPnFccmv/w0w5V16PpUo08pbTKppjKcoI9j6W+r1XJiCSEUUYLT8A4UeC2PhMe
4FIh2szNHyK+LM3mnmJdrGafDOjyyaMQVqPRW0HRA/Ibjzi2uVMgKzcWSHg/RL452vkCJVZyE/B7
wxohTHpoHLBDiiRfZf/Beje64odv1UdjNK0WDo/s9wJzjmsSklDhtx93pWqJwBWEihOG7FcfXkk3
xLuNgtn6UNla+tAQ4iCakzBSQ2VZO+ylXqFHJWzBREtnWiIsw4aP1j9/Za6k0poogkGQik8nG+BG
ja6J+kf52l7VhyT03YD4O8JWetLAkoiOo7HyeGeuGm22A38pUWz9OirjhzstTQCapqHUi5p0xU9j
8ZuH3ISyR/jIx/M1d1CfBBhgTEq1jASQ9MwZGOltPjtf75YOtW4ze0JxxSFKeC+saXi/UtEVM5md
BWsj+pckO5csh3NFdSX3m5taDXdTugOCuzt4qqEor3eh4RbQxF5GrNxWIIIH2jDJ9OHe8OrFjzcl
HqIF6lKNRvFzUVmqfgB3Snp42EjEd3K4VTHs/6fnEAah8RCOrPkSmo71rMX+cuKjVzAmArlaOSdZ
6QlXgvbVhpw6Da04PDD5IGlY/Iu7gcZr+xrjxbTGoXsx4TBgv5bW/IxRel9mCcD1PYLrnzQIvMYd
gimmho7kmCiOqURHiZg8os9H8P45VAw2JdMeegBLDxBtZXytbNivPTHwq4LOLAEQrVp81myYPeuX
uehZ90dgcl/PGvYxkfUaQ1UTwe3OdtmZbJiWYrcpWTr1yZSBoKMt1c9pa9ktIXppBckV21wC+bb7
PZQmVUwGx3OxS8xmhiCivN6uuc4F1uDvCYYuxp3LcEN6ICdwT5F/Ua6NrI8YwAamJTJdtEPGNN7m
NXXUZ0/Yf2xPcj5QoqnMH56Er01hWFUCFhu76gSgKQFyD4JQtsKnAQWDCYX1ULphyz9Nlu+3t4WW
6zBQG37ViTz1q8jWpG8m7R05xDSa86Dt68HEVlgCuHEEbPW4J6O1l1mBGsLwbrgz5MBazgffgYDS
8UNzpXNiMfLDf279SEkdxagWHlR1zxAq81rnkHjhLnleEzAi3ifjflry7qJzLlgkKzjeOdIYYm2c
o4/nmgiQIvQPN2eeHMbHrofBegUpeDLbKAflpHGeo+37/e5MM9jP6YEBx4X/wk7709d88OuF7YOz
Q84t/QfuIkR97MK9HgR0lAP5cetns6KGE5fqZ1ZBbC0onpIs6XR+PlIwTkS/R4jnHRQwK9w86rsD
XXzBE1MRGCOMJape7eiIJDRyxKKmYMSeLTLRkSoFm4mAg+RlM7PNvqj3uPfWtbNk7pAmRZe/hsDX
8Y3EW80U9HzdpXCR/hi1CYCCxsOGoUIvC6qyFrwWUlNSmjrK0TRrJwn0nEop7LGdgh9pmgbiChHZ
AoIk3NLsbgnOFLy8EvZlLFo/RLoeA9xCf4iX2bddzboWkvVC20ayjv9neQJjRDA04UUbK9Tf5Ykp
K7duOsSjZdsekypy9lm3rYcAooONq/sMPbui+h/35OnmTmaXYsSCIQQgNZZHtNY5Gz0UvaPP3R2p
ckduN4e8vA1wpM0Z3wLxrsf4rA8dQYzP7B889+7Iez+VvMP5drTLcVTGaYgaioVQlfsNde000Ws0
BkKP8DHL9YRKpPMopqYMomFLxw7iUWSNj16OmiK+5xB2LFz13uZssZ+IRfQmwccgd3xF5Py3UDuL
BKFbXRMBSyB3MfOvHvZBWe7UVjMqTvd+/7xpD2qgIwxcHq/OPwS7z9pW+wT1uNoIQ9OWmoqAnQxs
Xl+lUlGyEpwJREARo+9tAM8LhznU44EIvU3f9HLU08oy8Q8v11Bs5qHF8IjrrARJylhW6VoYnRNR
VzZVWKhmykm6wFUE+Gb66ZFc2XDdbYolvfuvDz/sY9/fNXgrpz01bmLkG37Ysl18RIbFJM+RJauQ
ulteIRGMQZtnHaB20RxUQCA/pKu3lPSBjTwFp86kV3LT4d/K3js51oNRxKOwEvrmpjUf5v1JNmI3
8AXJwfyLDfo1jglySEcARVL6ZSzmGP6P9/sVCDtj+h5OiWf5f/Hy9qgFS4j4bA+F/QlObdqOREK7
PTqM3FQB+WX3F4PjdT02aOpr4dRJX+C7RGnG0d9AGPznqTN4x3fLoDJ3/npVbq22UNTfpfpH9gbv
nN5udan3rCbJyS8xETofZOsYIgW8s1MDrtxo5PcI7cAenjxlK+Zi0B4nvyElwe2x/7eXa5T3nBjF
S1W9I5zs5XTq+K7s8SySdI/eD3EocO7sBBHp+RvFbGyhECeel0ELIaTtud96JfmdBPuMkbKoVPKG
QNq+s2e0LPAUPvyXJ/P48H6PYxnCCJ32FASTXSiGFdBeVFawhsjs0NJORP/BoLStjW8nhPOKqd4n
DpMQj0oND+bPZRr7hwSRSbSeFiQqT+BvfPC4F9eobtr+F3OWtA0R+/nkSMNRSA1FiNSVwUSX6A6F
nT25/lE14oDxHGoooeqgvvs45w7hpweWAhHjMk12ulXrI1kOGjNt+bYBgpilm03lLdvjSvnWDY7B
FP8ChmBjat3IOkjmGGzifKx+Hg0NWJNpIU4fizNmf8rPxwfp2vzQmILH7tdBC6Im+29BMOTS6MzB
vZn1CdiE2zaVQx+54w4/QdVoIB/VqqsKSLc15ic1ifF1ixanjrgqxaed3d0UrGAaSRvzaLX+PZ+t
jQLae7rBrjyJbvmSk+jegZb26d60d97NP5lYq0lAWQF3IIsiier8/buAbf3n2Ll5TB5t8sGFj2xM
Awj3JON2Q+Z9yRyKSt5bTxj17cLgtilk8OP/J3RAzyTR1JcOFmrKm09dnnSVIh3mcHYTvKZmbNLf
l46vpGwT8LxMs8rwoU+2gA4R1toImwZvgEQYO4S0o1an8dg09G839oEkvhTJs6LbPSQ3UhZzuAxH
GDwGok8h8JLqGjV+SpsMhvo/ONoxdE4NQrJnI+GPHm0ms+Xxox5VWDXZbtMmIozHWHDUa71KVlqb
nObHy7qRfBQhXdYHS3qwoLqo69dKZHEu+/ZOCdY052JW2sAhJqcZTiPy0gJg3uYtxqsCDw33t6z4
lxSJm7HYMriIrTgaw6f+SPBrSUvCms7XEr/EPuf4qxJs9A0sn8/PFzb8czchY3Cne4zhHoPVClzT
jxIci2UbmE/xJNd8tMpVa0nHC/31VLSWxqKE7Yrz7PLbdjxRh+mz+N63pq3NCUcciUgqcVbls4CB
6yWYkQcfKtEw8aT5674aQs4GVV601ep82SnZzid36pEsjuPyvzj6trkqof874aULJNUl7bGR8Fr7
94y1WBXaQ0Dl9mlKAb9ypBC7AKf421gRsdbznNLxmmZqxe3Y93iuyDcDSRQkwnKIarr7u9sjkzYv
2MVQGxiCjw3Y2UnyJLciJzQmAU/H4v0dkdkixSGuomJ4xkJnewipandTQafORaGsB6Gerxzgd1AD
Kb/WhqbsIg8E7xmjPNxQgodXlOm9QQU5J9+BgQr8wF8NQPEvpuOPnszSuJuPRM1cLeCiB84nnCm0
5GWn0O6dm3DI82iAqZuTsbPd1zjGun25etjBHqiNyRa5ZgWeltKA0g2pxkwZ/uBMf5DufMkXi0jt
JOXuBOaPLYpV8k7hhew6XkdHF3Q/62luH8hOUrssaprl4uvDEyHnJE7+8u2CPnefQ7cVxDL8KNQo
q86r5QqFDb7eQnUvxan3/3uIEaj2p3fWkfMeyr/XmtLaixI9zuNplyar6/f1lUSXHpomBKghCAjs
TrcvgmpH/A7IFrvZMIxLl9t8vfQus8vQ/BQunwl1WyHZkyC8ss760HtHt4/sqzg77NMuCFsGaNFC
1A/SMPHPAq+3lk7X/fP81aZETRJTmfdIqFlE7MyKN7lcZihDrcx6AQiIiI/M4AtgmjknLXlMtVMf
HUX4avw9+tB7Zd+1BE5vtFS4w1sXM+ytgFivH+1xaCs/4fjEbLewGPV5O+7F5i624oQ/ndh8r4FJ
fzPFgklQ9e4vSNtu9qFUvRxBDJWa0LnC3JjdXGWkEljNipsVNzGSIDo8alCk7q1jwjB9R1fqzCJg
B+7po0sjASY/57jeqBd+JBWB3Y1zTAnpcTrLpjWIwgsw5blD2rNW8sA+sRKAWfu+TyO1BJdfJvZQ
CSjI7stZgAxuOVyEWNy7LMJqDMtU6wsevPo8Dh3FYubTecJQoDW15b2YL13fhnYL4qapiZWLCWjb
G2KjhwGzSfthPCWi7K8fPzTGt2Lqd2hB92WMUmDk2FRIGfazZwV62KjSIMXPO0AsVdSXNwLlZGEq
4Z0Y2RTfIOVYX2n313JbRZ6ppeog9pLshP+XL2XH2A1TcpGNXcnnvWI5pn60/hTMDkC2dAEhU981
nxJ9aGoKjKiHfY4DGGJ+Jjl2WrppBbLiyu/oE8TM6OvzEozmSFX1pbqkMJ1bSWyj88PIpG6Z3Axt
w0uIOu2WdssYzpvI9Xwm/UhJ7RXNjwfA6Ig0zlMsqK07qe8V7yEuMPos9IMN40lAvlxK/l29hsA+
gTbr53ZEnVx3195Rdm0V7pidfZCQ2d2SlMQI48i9TDnKWo+oRiom4v1K2Ls5F0W9qmB8GL2ETZ3/
YVrsjazcubvWLqa3kXtljmMxvPShY2uDmJB4OR7Mb3ZHGZYVyEfugop5wWobpPXiqAd88prbCRTE
+CLIkZ8aLi0wKLSGt/1MWiVA2XCFXUyzV5+9AYtd2lOevWTQR+0dibuQ+9AB3cXpn6kJQGf8nW5k
tciosJFW1tu10BBHAAE1WO6pfcn02e+8gAvd0iPTofI1ApldSnPuDcZ8J30Fsq0gvR1yMZiBI9l3
kLRJj+m62awAdvs9XQYz3MIc/J9ajg0RQ5rgm/bYr6SHb5wJrXwwLLZeLO5xP8k76zXYWcfQAR12
QbUpWvEcX+WBaR/M+OLOW+ti7R3YrPEnMsQclCWV+XGmHuRjIzZkZzxGeCHEX2Y27/HubT1Ce+Dg
TSZA4R3mSAr9AithFWObp5HohIByGH8czl7ZIng9hR+as28vZQBs8XQFzPlAbGvfZ9JOADT2YrLl
P3mg60UhrHo4rTo+Q52FEM0OWjlIlYcfXEW9I3kwuSTF0kcnZlzM+3/NihFMM08zYxw727joSDcE
HFAP1TO0SRgsz6E9HIFTRuY//BOGaJbk8r/Sbmr4ugOHj9BN/86sgSIWv8KfBqODRRQNbiemSzVL
QB4mjmoze1ruACqkTCI0Howg7FCk8/RXyxRJkFxWpAgJz5faa4w/S9ZDo7TjZLtThTjZXKqisL1w
P7i2VMPBhveCF5DXFN1jcDHU9ivnR1k1tZ/rFM+DigJyr5d/3WUoSYpqflQL3aJehr0FNZmycqg6
y/31vsmqT7r1t5z6e8aO7001zsFE0cAT2BO+VGQzVWgwUKVWQu3JZscWZU+sS3j67rMOijVD3yi8
1VhtG0PYtdBaDejCTlFXA7BY08kCiws+5Nqi/Csukr1pddfUROhG0YaM4/70FvhCZpCsnNVNIiIw
KQbxbmFGaToxJnvjThwF/BjQ7Ps/WL5h46C6DTn5ighA6DZ9UZXg2bUwPW0SocxF4PGWV5iz9wYF
jSzj2OBRxkZY0mAzIzWLd+65pQ/dcmMCSG6kSVpW1CxWm8OkOT9YUcBRci0Lp7eP6r0/3oA7F6UA
E66NEBNTgT5Vazzg0Evan47hACW1DQzsjjjzO9yWAdOSORFLqogLkzITbFAI7eT4ZFEVPfqm8ANp
47PoJO4HjQU8Xg2DRF7v2QjOjHLBFMsmMNiOoStU18/mC2KKfUydwE4e9OditlLq1e/Y2vLZOyP9
XxqOZ9KJRpxJM9aJrLz0VkszDQzuVz2/JjQFvitwoIRIXsJxk+LDIee6niGOBPxyKg0Rdwxw6yxv
EKQgVdhxkILbpL2xRvKh1+yJvKDz4gNdlC1i7e+0RF2A9yNKfcni46b4CzfFqb2uK9HvAjbfft+1
KfJk4757EMrzWj7hqDnAWLfVNRdETVS0Ii/LmeQXnEmNYKZSyJDqik/+XUtIeryVpZ2fqj99JGhi
4dRmpWRopJBKfOpmcNv09BWLC7HbMernFkfXsxluLqX9HeuFu0YTSDnaGp0+2xyVvi76i4ibacld
ocvGOsSuHCMxvWXc5fkJBs/wX3PSmVH7NBmshvxE2O4KpuRYPABxNqMBDWrfJBHTH25bc0HkW4Uj
pMMmkuxEyVELl7Z+hjyA/TVfkIwd6qgm+0DCYAqGRSCGZLzQ5ty58q/GgUns9vvRttud3wHGQ6ik
49L8Kx/ayTCkmHhqMNpl//jHX/8dQkw2UrFhfqbehbdzBVlx8rlxAjfV3U1yLlJo1UO9d0UUWSOg
I8gZ1F4cqpU7V2KgxI3beIzDf3LjjZIJpgGZtbocv4MmYL0m1x3n7XYqdXU2/vJxcWro9iyH1G6k
0O2NozQdJTiUbxnlCJvSEWhD+Iz2EYQ0nFIEHIVxL+lAD/fK+I/cDYGUzDD6uwNqrVMSBN65YuCY
nDG9yRKL7kJHRtejar0DsGWIHS8lsPUKZ+nLyt3wEcj5PCuN7l//Lkkf4wC9GsXC776BjbXYCjWM
9tt6J+jecH3I9T1ZMRy73/hI5ONUdDZwgVwjkgo0E8+1jNSQCekw3oa17iv2/fyngBEPdrUkcoz8
7Ry6GUnQkVtb9Y0kZ7nmiyPmK8BjG9aRvRIPddIfyt3k8xvE7Of4UV/cZ/DVL4i7eR1fXPveZGEk
N5xeuMdkHTmARu8PWXhuYdEFlGJ9uidykeG4Wr9aTV3bjmxFy9qhgWJCUC/nnmVtNVNc0YfEfclk
oibyd1fdjq30MKHG9BpBqEhSQr6V9HGSr/hKHyngNhlQrebzn4dRkRs2lemHueMERDwkz+r9yt0T
H+ss7/B+QJQpRxdVzfR9/rWtsdrfF2oJ3zimDaxPdsdPTxeJlCy5Dz8ECNtTbJ6ISlnObOVE42/i
n5Ou1kY3mlfaE/K9Rv7GYmaVuuMCyAYJnczsyriQ4q9StFvU/xOe5kfjwjhY7H8ReCDSwq4w8/s3
FOLQLqKBwmiX6mCNulVXOw0eEwQmdyR2YQbabOVgJjeip2GbolKIZDEi6v8vry5tEGBXiPUzZ3+v
X0UP0OZYhqRIkntDrB51Lquw9F73WogVOzxV9Lxz3enHSFODLfM6cwRJ3pAY4QVoKnCBsyGHA161
iOQQ341XUjuWykGJKlaCr9NepW+TyypFpIawmlM+pw1vcRVShROpBLCIH4Y4dyI3Irc0yIcbax1x
SUa1X3AnwRa5HFReOZVrZI25JCc+pNZaz0p5spT9jFussIj5ilLMyjuvhaadjj1Xtn/uxbFoowIi
08OPZFVAkNi9/t3CrsQqD1Rt7+QUK9WBPOVYbInR2P64eN1x0j5NDWRy1P5+7SoUkha6L0aKimM4
VDhTaTMk2fVF0lgx1Y8u5gFvdLhC159tSmkaVn9dymGsZTn1NrjWVfnk8GpW2D7PV+fVQnO8uusZ
TF+iH5x3CyHi3yRBG1Wr5w5gJJ0etBmpFtSKGyUjvJttvx/4sGSafZ0MUlrhklQ9fp6x85XnHwEE
ZgJJ7AX5681L7AAY1OV+RRxGElJ8KRR4SKzSk9N8M5vgxZWaKM64nrLnQ40ZTKgH4D51IfabXFWc
yzMeDwYA+u3m93zM9YpNJ1BsqLEOzjo+B+zycBlR6Cnyect+YEM3ojQhJivsj9F8El+xEkwUyhQN
Kx4i3mU49NAhwJAhIK3QW4GpS0iEy/mSM0xt6MW+vOBlkbps8s6TaLhhUnuE/6uTqoALFahq9uPx
Wpxn7BjwwznXsZmdukW3x3dPBFepD/nW5QeMByIVPoaB1Mv+5HiNURemVa35dz0Fp5OnW9OaVCRz
ZxCkzUVMba+5zm1Mvs3yjggLv9h/Z84qLeigQ+6scy4/WzqGpslwtpZidm8yecqsX5QKCX2Mnifo
VYh4TuufChbFXg75QS6Uu/uvh78MyXdgELYmqAW1vUjsBWBYDcYOtjAMtjnlPc9EiIZeu4avJGYP
wsCrsMKwFp58/YbPfN9GFy1XEbYPAWd9gVZQwCbdg7tKpPTgvpjPXhGtRx6Jewc8oapbCM5rBTml
ZRa+hKMiF5OPWOBV5/F/1BsSLfyfbUhbC4L8TKQ81zbj82tLt3Ne1WlZpFY8pkWDNLeylt6Kn6vu
HPPgOgTld6VvSKCUGNgtzYtG0oxssjEr59IMW6VtL7L29Lxdqd6R+KlPJZUxe/PXz81CMrEYF5Lj
k0EIpXwdogfphGwYx7SqC1l2d6Sk6AwkCoI2aj+m2CNW1bnPM0Su7NUsWYretEKn/palVcxdAjTC
BBHsStjxfptGFTGrhyZJOyxzq+u6sRZ/pLvxfdaX3HvXIEbutX2hty8VpfCfctBV/QMneJ8Qe1Cg
FWy+jR75o463XbiCJgpmOLqn97qAUkPsMuclFDkU5cYgeRyl161ec9DyEOu9T9++ICw5TG558/sn
eqPh/dWrQM9yaX5EdcLCJpJlspxMUoheeYG3qzID0+tOSZQBIzFgHXkEqGJc2cr5ouiqeaFc1ERV
EAFq6hiI9RKsZRHufvQ8eqN6LvJVpUabqc3qtfoiwAMniwKtM/AURcdLiFkOpXboeIuiHXigCjTs
OQBXjOd3aO8LjscDxJvXVtpkiIt0OOaUeUcKTlKVZJ/YDAJhboc3nJnTgCosD7YBwd3X33AEVrUl
SKxturCEx9VRnWrtKs0jYf1oyoJW6oJR1r1YQdsJF+vxli8xB24OU20qgvY6RNXhkeqVHLtnBBhb
qRsHikAf4RGJjbodg7HTMSRwnvbeC1h6v9+JRZE7nQ5r9N0ScRqpLSSgrNIp1erOR+8qTzzGkr7+
ia/ykSPy3TQ6S1AdlyY4j9JdUTP/ASC5L5xV/FgKxuz2BIhNWW3o6l325Vavr9CJOlLCfCpbDHMd
1pDQsY2Ua7zFK7NQ1HB+mDH8V2AirMsb0PXkvfA72R7F/S9OTvQuaR8lEOSZr+ZMaNhWVFPjUEHc
eieiV3JeCp5t/beHD0vDn6uD/yGpKVZCb2+274ylGZAXVYfSN55CpSHVi9dHqioQGkBIplAkDb9M
A/+rbVpbZDuoRhE5CNZQol2fNUi+fZNmDtlClcMJ1slG3BH2STQAYtSTPDfxas/ZHOF18wizYVbX
OIdDZp+7nvR52TJQYC6IiFKMS9C2evNu8I2bgG8sbmQS+lFk6aNKYwdPapyvluE2WcWAx8N/5ioY
/37isqdHodw9ZA1tUzroxJqiXibljEVsxtAtQXDxRcdnDGDMgIUz/W+1R7AVQ7q6CKrYnDQrA2Ph
iTStVFGHLJNTxcsMDypfFhuBDPc+8YfG2RXiDuT4EG3R46fvAHvYxvzKDxDfSY84DCXj9sf0Xg/p
eulqjdNb5QQ88v+e9cKHdAtA07k5LXdtMvN7Hwndm4pRvshPmK6DILUMH3WuRMhcKzdMV8qGpwBu
+Wj7J54um1I2e3PzM5AHRHKlt+9AWARZ1VUxdERm+WIAGuk5tmbypFY/5RTO21KpmNeLN4w0dbou
knBiu3tI6xoPzC4nr7q8EQcYx0jflNWjYsiwuACQBCPdpzzz60lDtItd6+MrMp2JeMqeeMQPS15H
6HoruWFufVNR1LOLt1ZR+NQEzAdThD8svoIP7PV5PXrJ1T4VYgE3RzskLY7Lqif48+IkwCBpZD+n
SlF1R1x8Up29Vyp6FE2gT+gwlWAqR2AJCch85IysacawuXsZy/i+bxtaWg6fRWZ5gAQzOMmWxqGG
1rZZgQPaMTHG6VyHs9jATyCO9o9jfUINyGdBj6Pft1vvEyOg2dA+A1VbcN46ZiL+gnMmopSkROBT
Z256nDAqhmNcJTMQbQcflH3CYMcaB043aP/Ow97cM5eRlvEE73wmQobTNf3Cpqwdx6FPx1a0oJ4b
6bcfKAcExF21QXbqJ8UM5s4GniNqanzKDlxt6J3Vs+Ve23P7cksqnaX7FHBIOMqhUUzKUBDmrlAy
8ht+kdoghJK2laV4u4SrHMeVHMMGwcPmQQF267LqpO9udTFpwwATJIK+Yjs/W9JGpZFUAo0RrHsS
eIqJ/WBtk4CNW/htbUzaJ2R0h/m6rUXDAFacP6YEhxJYzvmbiRrQOhwHVcXz99bqr/gTbChUfbr7
I7GyV4109pHRHq3pzSHcQ9MwokLL75tWCnN8yTsQLOtzhGkvUdoxgyri3xLp7oSwIu2qZZxczboy
/YPRzbXsmJEVG/IKGcgvRvs5d+OcneyBeVmQgUWUz+iNPRsYZ2DZGquv+eCDiFXmGrnaur7H+n7e
GhZlk1IFiQ6MWPZDTpop1PEXHeP17YdXdFpEGd2QKgILtGegG2isNsLyb9ZZlCVOLdKQVbfGM+qJ
OcEv4eu9exX+2Ei06ytJHj165iIlo0FVDv4DtraEX3g0A6gOmvmK5yS3CvF9JOVqSgoUIcF5UBwI
KqW+58URWpZ+8VNce0zfZby0Pv7BEv/qyo++xTJj2Y+CwpbFhNpURcf9aU6zwddRJUw88lOvbnGw
aZKVxT05oSiJIwpfp4Zj0O4X5qexsvJdYmSbCBhMHZI1EJQlwpkHjv6ELacKhnb7+hFXbK8Wha1y
1KCr+C4gG/aTCqha6Jhknr1gArUP+RKo+m2uDbqHeggQZ3l5PwZWnDfg5Gg/FjZMHXu+PsdboWcv
us9aBKiSLfviF+NPejU9Y7ZWcScW9SUHFyqULeGMwQ4LfNvCJT8/TJvyFz83Zk0GegVJ13QYQFNq
mt1XelMs8bD21v8LV4r1v8B0mjBhfKrJoKI+NJCd0WJNorayBSlSHOT7yzjZfu7NWI7tHR7luJPT
FqCp7ONmCjlwRq8s0WcjZWU+G483sAzASnMRAL88foWh1EW/UFyBrTOGVX+BZUhgkaovavJtvAtK
fDKpS6/1d98SKVP6OzTeZf12N8TXUGMy5G0ItMk1jHuHdIe1a+63uZfwr6GhAdfppUryeRpXPZv+
9cK+wJyk4wdQ369Fo6D/+2ewtsu27RSFVW2TNO2RzwzTCmYseRgMGuFDytem5ERonrVcB8iXCMy0
ZAbpvrT3fjPTiM0crgEbQvbFxMI+v9aV6XLwPhwhrHJc+9es+awIPWhBaDG+niUZ7BN/K0uH6Xqw
Ty75oFflAzR0Dn8x4Jbn6Kfl8FPFFApguJ9CoWxLPLdY5t/qL1ohezrlB0WvlLxNVMgQaq6p6kfQ
8KXPsFwseePWfDVE/BgMwvmW9VT4ayAKKwH4e+T/n+EGqR1v4f200vqPiKeHifBR81EsM6SmnIRD
JpXEgG+fxxWpFR+dk/y+7sqbw3ZstHjpVC4r/6fbI/KI36cOa28+6b03p4+614qoUBYDLE61oJlB
aa6OA1V7XmD7DLt0Fi4T9ZdH/oFq6bj6sct0/zMLYR6uHxhIHlzt5siz1vryYAwNFa3XgIFMgjA3
VrrEYXy6U+9LoyUcuAwUU5iLZa+7NsdGG3b4d0XLmO+CjeFofbLIkpVTgVjNCba0e0NZapDrhDqV
/Y3FFupCKRdOYBcuS9AxhC7JVkmmn/LsQnHNgg1IZC5CZDSUS9JJAJTZh15pId6Rc+UlpBWKdf3a
NmpANFqYYyrsRPcXdfH7v4DsO6SuDyuHpI7It6mMXXwl8EUL23/ULFN7LPpvpzBMxcwqX/sP2tII
0+VU7SQ717aaLXbhVQaQrqRVz7jMTMD2pBG1cg9+1SxgIKJj3sUlINX4MtSwRORQ4QwuAdahhKd4
szwpStQ+mkAkIf8thRqBPIOm2i+kJvpThrDGETV+5NUmwi7fZGlcyc4mtyXxV1JUGc7egvbBzffe
Y3NMYwFUBDnnRQx164Fm6P0zPPvMxGdvZF2mwXEvtP8tuQCl0rmdju7YMfj8hsomymff3NWOoO5/
3Kj/MDiKBVigIg8bkQ7pE5JqP57W07pygNbl4rS88tWwuDumTqsmbnfnumHN1KYPw9yLc01U4ljV
XgcEKd0ZpIB5g5N3bEO0TIobeQzZgTy42RaIbF9XHG/QOCbaho3zMs+fhb40N/LKjmmUW25MrJ95
pRuode2WWxDyLhF8EZiITY1NDaixYIK1t94GOQh6ND3Cq2/JX947NKs6tfq69yoNldNgqpi4A/9P
hkExuB1ufvndoYqoWPQVVGwugGkof8W76jw5jL1lM2pQS1NQm0j4TT9F2j1IycytOIBnBws2DGG3
R+F9R4Co3SNwFkaP0jdSeu7guMP0jyOxB3+1PrU51omNOb0So63KzUPEzQkXcqaVYLSZ/PKO8B49
luAJVn9xMeaShAR9xlx7bKydiwLyjbr4VQaZuUGeoPt0pGvWmCBJsqzX3KWyq7S3nhX0WxawieiG
CBiMYu91qT5qSGtFZWvHWvKCdxBUnBuu25PUhBU8yK5OrJYbNoRdoxfrSEjpXD+SjsYwFsJDeIaM
2YZOJcAtGcFhKvlM31VzBQFdpcZXo35WfbLs3NyJD0FZplZMLutrfIjaqXgDOCNKYTL6SnDacfkz
0sxSw6czSZqnmSs0zfUxIxdDPmglNPsPPuksxhFLRuSUf7vrmfLDHUNVVpY879lkgnXK0q5ZPFPg
AvbYHaEj5MCNi4XeZ6q+Mtk7NWDAe1+O9unwHS9aI845rStCLG1ss5kMEE/iNgp20WrM0MEzw0ez
nrxste1f1jJB/yPAOE5AWadzoF3KIG0SGyTrsz4vIQzI3oYM2N3bL1SAwd1QXY72/076+UcpY3/t
zfkN1MkPjrQPFzynGhvWGxFr//lBeJKU0rbHs6EJvezlHpzPeFt8H8+Sl+x90qxlcURSHQwJ8DEw
etvb3tcovlBxvnnM42liYnFjfWnZvWlR13161K851vnTx813jrje2pNc6xtdmYxN8epl+YD1oowt
jxMrFKSkLKAdvVhx4meQeW6m4Zzen5nY0hrR0qjiBb8D46NRGyxvor+eEalbdkzmMMvBRN/DPgrQ
PRDnYi8f6bVh1zLohSvm8jW8VqRYQfLRMJ2Uw55uD9hmlXakXQ078B21+A3QToY48E16RmwAhsm/
ahya+QmpR1jxSOk2hP27XviePrD2A/7me0Kj325hH0TaQX+2isqxol7JoKr8qKZbcTdjOGfiDzid
1ZKMNQfdWhbhpKHqlux4HNzDcUJvjvJK5o0pAk3J+KDaw58jvVwmPWwpK7Jdgd0NxAcTr47JwhGE
SGvnNdsWUIIClu6gGljFDPuPIFQfxG727vAPd9HZgIsnt6PdZqOBuwuWoTUNN8PX704OEhbY5Qj2
QoXphFbZNTE1x4hA6PAqbmldrJd8xeA+Z6tOCDXCBZcv0DbIQtfG3rPVvJLphqh4ErrwpbcWiCFG
uJOyB4/YQWxC+DeWwLoWVN31tsypFExPv8agt5R779V25vO5ZwZutehhCtzEWDQPxpz1WxUZLdHC
owZ0nodM/MFk423HbBnbV2ofZ6Cf4/BWeo8eILQ54PrnBRxMDWvw4WVFSyNjESs6W01hOzg3Cy9c
V1lHYog0/0EgacCCBqmynUZHq2F5w0XPLxO47M/67zJF6gm57enRJWiQK5Ul0HteHqsiyFelNa8u
ja2JWGg8IMf/UTWNIw0o4LuRKtWGfC8nc0s7uVGiJtM71BWhSDhcbO9ZSSicGD8i0h7pYqyaJpre
ezNwVQC5BcCGtS4F4Eh3rgRp/ZKk7BEBO+HTfUC43ZLlg0n1YtLPB3ytwSV3E7jvqhHvmyXOEBoh
BlGcbPNuaUX97MY0oFzpdaEdh/lze2Zjxdj6QvshDPfk8sY29oJVI0iNvWIYVJy8lMffkOYr5HOo
iWROHe0/2U7HkmRq2NZDf92506d4MdAbYB6+L8+7cYPSEkslWZ6IJbU2ehlya+xlvqVGtlaGhhFE
HbLw/xNSDEifBuMusTMqaWCMFC2G7CB1OMRSluJ0D113YCbxxHDyUseBVfKKiydSAG5WBq7JdNO7
MQtim7LtFC3bJSPv2O85Y/L3QvxcRP2FD+dZmVnWDDs9upLewwBpRXqxECo+u2Mr9eqKq/O6SmRH
Y3mVVB3Y4B+TN9S4zqnH7lX9nxZ3+jB5fi4ZdELcSkvb8T6mO9XSp+le1IkO2tPPN/Impqn1c3kT
J+RO9QSVEufyi7YRfQn9wjbkkWBKYqe34lj7DU7gBWj5U+3Rdc3IuyFlGPrJF8khbJIets5xq3ms
T9KXM8A7NZi8nQcQUL+8v7gJ1ItGDCP4kRaDAT7qcNIdf8p7GI2vufnTX2yB1yVGCli0qxVyHzIv
zelhp5UvtgUdeXfYzduRcLn2QqYDdpRhLKFMxT2OsLxTeOuA0bzjztB+FTrhRoY82XLGQDZsPnAA
oXQ4U8UgqUIhZJRleBCSZBoVnyvyZnOX2dMD+CdqaRq6xM+rD3ejQkAvz6EjVrZFylayFfB4V4SK
ZlsRNSpdp5hNa41k/ocCDtxjyw+g7mRbnOdiBo9hosKFJHmPgdC8J/5ko15GH3JSiNVX3m1wdIdf
/sCrKhIaDPFvNgjzBrLLBB7vetV4qYWllk6QvJ25qqq8CfehnyP5EG6Nkw1MDBqiQ4VkFbHYSv7k
l9VwHb7qcck3g/PfO9BroJ/FK/rl0HCVFEyvGBSZM2P/smXo9vTcqbvOvY1yU7zOPiOAcKNIKU7T
FaXMKSNEfAtl2FI9RGCGDQl7TQy9YoX2fLsNnA1LH6U2zHa3+dYTbJnMQjEVtFTNZGyJADaJxwEo
UeF5SWUXAN0ntdVH1uQu4af0zxzbgyzWLxRV+e/I+g1GK12pjFoQM4aazvRNOaBoLqfJuSTtj8Gy
gmiUBeloBELOzsmKEttLm/wLU0UIPpEayJ1QPWRx8e6JepGNVP/kXKcqMQ2AMTO3k3rrR965zPYC
oF3+f0pIJVtMxbzSIQ4IuRaO6FD5mDd2PqaCneQXGxh/XZaJFlOQ07goIk/Du0dt11nxyMlYYeXO
v6Ti17XoXVrMTehmBjrmuaWamdTpiKmY3G/nKa4FTIXXzzugKJUQXhkYdTvvNbYWs/dOELE0OUUE
D8r8h7ZvLBvDIh0yT6L95fJ/0uu+yUftSLDZ7lwBSFoD6MvAY6qG3AHukxr8aVwBTy0NGQe6ZUiS
I9tEfk4Uwx/Rl5S1K9THz2YnPO68Q3ddTGv4O5noTrWXoWLNSstoitSCOAN5SX12uzlL2TARyQWp
gp95XnoZM3JK5z25QUVQudM723HowPDGRkBKHh2F+bboXtLXTe2H0Wpvs889XpKAKiS5XwocnB9s
FFt4EBEeE49H6o4AJHHU1CLTfX148zDIhlA5Q7kuQV41xzvp47eC4EFkScuAU3wyPFAfPRx6C6+4
OMRZaTS88YGApJzyvBgkQEzYUZLUs9tbTuRnhSnmuDZxfX8p9rz3jV++nlqwAj8Op2s1o5iYlfOt
rnHeT1xsSVL3f3QivzzvQR+ChnRe2HXbIBTkR92wzoc2trRQxtEsytjc/zxUaJlu6dmTlr1zmC1w
SXFCQcpPKzmpystS0n8+fB45sW0AB7KjMPMDK6/BuIjGJ8vJjrCLSUIFD7MHgtaPnnRw/haoQaWh
ttsxz+3pa1bk3iPueKMPgE5crnmC8bXookide1gqxHGwqnLuV80frktPBV7jeCIM54VkMUKcjjHx
m7os/EEmpb7ECCVyVP7n97n1ViS8TAWmj3ZbnSg9PSskSNuHddQwmdpJ0ro6RzFo9PfgdMN/gC+B
xuYXThZDzB8jBmIJodTS+mdow3STwQFZc7L6Ix3W1HU5xLg7DQJlLB2mU3s+Qfq1xE8Uyfgt6u6y
P/H9ZZOxLNAGd5V3vENgw32NHMHCtUqYdNe/FW6EvAYJXRF+c1okc9J3n5v8MgV+JN2PqKLFpnV5
KO7afAsDk6UwanP8Zd8tBbnsXEL2mDPNc7iKC12ckMavkfVfQ1hZfUNy1jM5jxylpVS+Ih4tFnG0
MSTsqOApY3kFkbisUF8i1y4E2SdD4ble6h+l3fH9HOaBXWQwCeHd5Te4AvTEM2+bKjaVmLFQ5zkW
FzWZwujyWP5vik9g6gMO7h4kS8iz6mmolpYpfjHrQHwl1atLuedlpY+ZAQhJ1VQnLVtp53cXcmlg
KCCKj1JG1ZDTXCKV4WRGHlCbtq7ctqg3cS3Lynsfdo0X+140ezBvm9s8aA/iKxbhVeNLwAH9LdE9
fo9fh4ObrR8o57DNVgK+pdcoEHTPb0dYDjh/WNLySxMceVAd+tm9Kr4auomE62+Y6QQ+0X7K4W0i
gvyvVHZqPQddtWTp3r2SebOdS/cwuT8cedxIQw9VN8VgKbKc2mr/KYyBTz2ae/RtV7n3WXnAx4xq
Fe3bxfmGvXy9x36oPo28JrOg5OziFgo4sJ7bIEEWZ4gC8vvfyYSuFhj542WoUTCl1rMYhzLvxd1e
NOoc/kUKLzk2V0Xa0Vi+1WncTBm44/89zzl27ayFy+5J3paSceDquWnUQr1vUxUk0paX65dbTdQP
RbAwiMJuvq3p2g3LE8F2gOr4n/b3hWK9c0BQl16jGoQQUX5OAnrKA1F34RgQHx4okkE3bIiuctOC
7Cw2xPtE/IB2kVjyyBSdyoxknIt2sPPEbhPEblz2jY5nmj4M8BZoO4DZ/Au262GeiaghtqFydcd/
0dDTXc0Os/Mubi/fe5nxgvGCp0zWgn/aJmlq/c7VClw3yrGXo9rosE7EHGE1GF2bpSWcHR/dSkoO
TIK1T1g4g/chgo7UKk6NAMrwnEL3KO4q40eILGFnYkCGWHmB4nGjGi7xfZhUQzYuBY46GmNo27kh
GDlhErvsiUO5pgFAW73VDKSrl4LFCKGCtft9ZJKMX70MPzBIXl7txeo2VZeLaEhh8+Oue6AwHQaD
oQ2fJdcSeT/H+riyGhJ7MCeXyCH97GBTYdUrQkXu1nKej2ubFJQ6eV2/97ged+d0LoJRQ0d7uVcN
bDE8kvcZj/3VWmSUvD2uu9aCwtpciUCMbgQiw+45hpfv9X3SBmny+gj5rhhDN1QiaXqRufCmNcJW
iwfCi7eR5/Rr9fZSSG8xuATHa/Jju+xpf+t404fvBcUJcF7/l+9gQ2KJ08/KqDLHP4meViL8CCzr
UkNlPmsyXgJCrHDF3/vBc3giwCJpuuQ9Djz9VaAWJfBeaRqvCL+P+8t59xiesCUJJd7MhMc/p5y5
fLWgcbgBVUoqd7I3RtKZUYBQTJU9j9aXPQJZ7/1+RDlM9y6H9avTlQbP0qplRaN1xFTn7izFNVnA
VKnurB/e4+E4LQ4rneuVN33kSl9zzirfH6aLAnkgdrcCrNeFTOoIuQvTxa6Hw7f5yWTocLKuuCv1
nj8QZJ1rEDPEAgYU/ozmd7/nxI5YGjOlV4Yonc9CLnlF3vVQ/b4oFlamZ38lveMFQMbh5sDo4VHq
pwc1PztawPyMASwtHMolKx8tj2Elf1dbNQy1vOW3D4v3xHHxftj0sTYNScJQeZzFCAiqJbl3YeDd
SJEP2yHnr6jr6TmCOx7Nt01+OAtWwSYUdL89eDIw+LDv2L7rRyDNb7+FfUAUBOj6aVrFdL1oo+dY
hG1lUPaz4mvCKTYjs0Cba7AF9C0/lQkRRnZE3EnWcH2vpvzFBFJ8tm1AiYLeY/rFLlAGfHebttNz
etV/3TQPxaaBqYmqcASRE2U4ramwby7pquQlKgHFx6ZgfwBLQfvsKr3mbnM/GPsBHHJb+x24f4uI
QMDfZpRDdAisHzpVBp3irQTbMHJ3ur4QzDi8Tabojy973qAFSQVeq7W6FyB/rA3wM7YG9zrja4e3
Ai+2ZgV2REL2jCaFp2PYaS1xYDe3FbPnL2nkjUBYSs+n2BVU/nbwIBqGA9jduS+2ZG1srQckWB2W
S8ayvsmlF5AiUxWx997YX4K/qYaBzB7haBcOx7I1tOhXBNhLAXlu95V6371iahp1PuIGONN1O4/e
/AT2a9sqm7dBMiBm8JRujgiBDSjYtwm2RMy5ktqeyzq9jsq6EnehfEqJX4IWc4jhvIUIvM6BOg07
chgTmrkwxjVN5eXVpPcbvBPtM8g5eIO9SE3qUEYN1xvXgwqXKD3j5+9G2L3Ao4rg88VaJGHvJe4B
LQA2iS7sh1wsite6FffIl4oP+6LYb6/77bGwlVcPHWdMKkE7J39PB6X4z5R77yC1s+x+M0jSk5xh
ONqJsrcDhWyRRjqplBR/TO/XbdpeRM9pduvdeADhj09eU783CP7QiP+YhTF7MLWm+XrdgC2F2yyK
oxXM8nKuVrQiZG+GKiu28fGv35aR0xvD2mXUglHt3VKXwrMvHCPki/UeWqHQTDBgehlfGAug5Ux+
QJBxGmZLRuRTiKhMQjEFDgcMx1VODnjEFbDzuzXVMqTnTU5pgvshiiQEDcJk+H7aSf/gLVnBzxp7
/tnlgZ4J/B1C/5xyrKVf1Q4IWum6uuwskE16vN+3Nqe6UXm5eYa/nJJbmPzgz67vveXR25u9jZSC
c3gockGKIKKRyZ2UtcHgETmCZpsSPAsSBtYu6+gHM9bCZc6GulA9qzIAFXvdpja1+XQDbV9ehF5/
9YFWjBRGbnsrEQxOq2L9CseKpUVrnbMFHy4/n3PUtlIOr3u3W7/XK3+OWX7EjoPlP1D4Wd9P7rUI
9PHliYwtlp54Me5+6+JOPyKbBxuR1PmQ4Ve7eaOFLiPw3uo9OSrGl79u23MNkPvRhm6il6E1dB21
s74Q+wCePMh18v9r34dZ0YTE1nhFigEv3R7Ta1suwo+beUmV7yNy2jlCRBbqZrTgs30GqLm9OPM3
3h2vhBXREtrbFcYv5zjSe8IJeBf9z0YsuoU8+4p/q2ZqudplnA65ntx6NmSj2eje9i0bJ4p0z7+5
L6mghac7H+36Tn47l5opRIk547YhD2Ors1yxw1q5dCd+kb0Rui8xWzE4RD++KRyAmxtqtpK6sJ/U
aLnpbWXLIv8AD3H3HnlXDFxwB6oX7pi4vVt3zh09SmwfaKaAuMhZ/tTEg0SmXQGfMxZAkSo1yQCS
LRyKe9Y2Ro4vyzHQTEdkWCXKLc7xEPiy91aRrCguEXGW1eZJLiFATKsetDGvrdj1OXQ2YySZ4tnS
Opvg3oo3JPVnIEVO48wVT8tZ0q0cJ5ThiaS2ZKzYXr9XtzjjoC69zt16DGCKBoccpnRem4ORM+72
S0lEZzyPHz+TsERbhk5f8phmQeByOUSs/sn66qV3Or/V/Olkt4dj80faJTkgBqc42hOIyqFzD44g
p2+YgX4n0sZnCLg1G4hnuqG50zymvPBd4+ZRdQxbM9fnz1nPi1YAJ1+fT0CHfARYC91ZPCLHZ2j7
sZSWZYdl6+NrDF0to0lLS9xuBOvAAPIL9lj9/LdYPeRAXH9iCSr5kfzIJ5HYEOqsii93dthtn2Rh
NzBaTAGllic0qKuNyCgNdsHcqcgvNoqUNL/drHuXq6sHUE3+OtYZSgVCbVlgGvwCrk/HFotDu9xE
edi6QnFb9X6ZixRo5Jp1N5i6xlr7Das7BmQ/ZeiSjtG2PS/92fgwar3vTaQ/wn8GLWfDr5QKL7c3
I3YnEmIFp1Q7DDS+eqEPJzHFAp2WQwyKQpKian5IbGuLuNIsNO5EqEnxHunHulOidEBTtklDAfmx
FhjdorDZi5Ab+K39ChOBuhiPrJhUcjRYq7Txc8i1AMaCPqNRfKWP3kyaB5YmRanamSot16uEbsKP
gWt5IMkYvz4Zm0nr56JkdMDQvsykr45f3qdWtB35wnRnGecLlXEZIvkJIrXDgQrrsLQwlfVWNMGL
7J+2bELSew/6aIeJwk3qf6PaNQt0M7+tnJF4mEaG00/vb5UII0etzHFPPVzNKXumeBfF876cN6Zo
rsKMUBUHtnNj/pLVv76x3u2w8djCD4aaReEBu7ypM7WN/eB5L/tJYZLUmykJlNvkfVuNBB5f+UWy
SyVwp9CbwIIbsuc/GLq60lkD5NEsfRMffX47A0PrIk4F7aRHtb9UfIaAPs8U/htRQoKL+UbpUu56
rpIhzYjLRzHxkGWgxbw3B/508VNQwPifgBifk3nAuhsk9Tr9pA7crdCN0DASZCy0qF5WNzG+iu77
JnF/KYO+x9fLoI61OooQD/3ijCYGGyaK6vA+jO+UJC8OdxRkHtJIIsD0Ek5EHJJg/pH7WoYgWoE1
LlqXjgy4JFAoQPIemXoG2qGLUhXC2M7at0DjL+KJPv4TvACSrKBrHRw2v4q3ih2V67p+3ONNwr1M
vVy+eVUi0NPBK6rEeHIdddUYxxua5wnkg2b2VwLxYdirGFrZk76BlyBpEYOvP/FhDzAWYphEl87z
5lV5Q/D763BLtAi4i3bBDWLUSSFbMyix04RnAAOGC4/cmJ1X2QyMEdD159gou3LMd0Pzyp80TKmC
LpjAwHuChbMEoWN2CzUalN/8W2rxppMUanqlW3108sqUd9cr2JZrL5EsMhPO9fwdHLwOqGbTTCov
4Raqixtx7lJvBaRwmmPHY7lN5/qHnM0csiEvOwx+sA7qr5OJUUkfzhKGlrid2FS8ukCITXlSDlHO
CLtdFDgxTRcx3pYG8zQHH+0p2ywrR0EfQmBH7ppNyit0iSAbgD9d4VmzT1VcfWUxrr3hT4SKQvMU
9gMCpgE8qwTzwpwXhsVssK7EltT4QCBfGIa1dVEWBFK7n91obA4cQRTIrQTHRaMJ3YXS0DcaBp60
ANQX7N4Qg0FkLRtcrspFq+6X5Uf90g7wIMLjRHokFXkYy+IVnScYAiEtW24lBQbPbrYh72YfUyOo
CJ0b/UrmmrznfRS7yddSN3IBPTSeMfJTcLtuoTOvEo+PXdZw9494SshzyRmJnrgglwocQh02b2aq
g1CZieKM+gxkPyvygKZP02cV87jL+XIeVUWKc7YAE7W+T0IlSYZszeA1Kfqqhtow/5P9yKCyOoJ+
Crxsq9ANVlG6rcA4AoqzvSZLdbMmkTJQPkwM/5LoLOHqwxRQ+W9T4ACWyf00s0aON6CBsIloDOEq
oi9YMhBqUdevwqT5Tlqcb3vygOTRdPTkCIICYQvPUgpmb9QEwo0snBWDcJ9TlXFomkFszupKd9FT
YcsICAulv4gceTt+UbNCbwrJ1o/xcax9vDWFrxXwC1iOt+N8CI79jMhp0VPlXkUZsg8cnD8tNot5
m9QAqAynjAemiQzswwHJViIsUNwSJbTZeoeNeE7EBNtC+ZdhJT8pa0PnyAo704qIleH8e2+wzo2C
bMwjQerdJg6BrkmAjFGijSS5aanZEY9A3m59TGLO1/FB9BmIWiCWyDXkePdWA1VhrQCsuUo2aSVT
+qHau5JXkqsaJMwE19l0fwqd+ybpmQeF5WpW8Hfpq61KUHCPjdPfSJVZnyG6gjWceYJmVvE5dQvr
xoUXzsj2O6BuGNUqq91m5UmjnXNbKYUF3lknJu6NNNund49UHoo8oK9x9GzLU1GhYFX1vtoN1ODO
hpkOpCRB/2SINQmBsCLmbs65Nhfxce0ALeC40LHMoRUVKF+nZ4bi8nIs+z20fqRXVU3n/dvT5qMV
Z1wbMRmaAYgKpHwzos2n2UcHhorBDStbga2fyACvQqJ584W7m+8vuhaMLobJ2GMxBl1bxcWtubt8
RjM6DzjEDtDby798Id0PfEMrS4XFRC4RGkUwCZ0z4/6l9zHKa1dDRww8ihYcwYLJ9fmVC2Ln6a4P
3PSiFERImHfmi6eghfezjXoKrsSNYQ3epxHAp1CnYVrvZdkhYfzm3ZGkRm5Bfq2EyFZJo/qeLRTn
EVICnJL7IDf6LWK8VgaM9pH7TgA+DW+OuwbFhLZAYGumsmJJ/Cj3HkxbprAEG0wl7Sr3OScfyk8X
k1YjkNGBqAJWr7NZpeh+oceSFdAKf4LoKXn5Gbz83CgT8hVq9SwegGWQB0k7nCX4yVj82MaGwrFJ
gouqsWrGMoN1eY5OiT3HDZBUEcJeKhvd6N64G6swYFjrlfWpy1KovjDy9Nvzi0YQFWWfdRozJtME
tAleNQH5hW6M5Vuf3AwBB3k904tupvYNTYT65muBvXUpXZsuRJADJhI/EQQiOJ3S2JBjrkmLDhE3
slLNn9wVsoaKoKD2rNRPkaXv5kp4FU4fDDYyGMNM7pWeRdBvGTZ/eaJB9AM+yKN0Y/vlT+BmquCg
0nnl5tP426R7+HSiQJS17FBul9xx/U/RBfx5U1yxqZfYDJKqGpa+DrpsqiF0VaQlhS5J/63E6SpA
trNtQUFzjy72oz9uixLGL6S12W303Gt8KR6i8wi28nNgWCfCAgj6OHXiEeUw3SopZlT1VHYfbnyZ
GJgA9gfQx6dn9sLQr+L3EK9jcyhskicxyUlwQwFdE7M+a1cgRBGfIFczErvk0bSPRxGvC4KW1j6M
phOrrgsg1vbNNxOtul6KW7XflEDqvP4pjb0c/X3bC1jPIgM8Tn07jq6Ey0OEg7xRyEZz5omrRVSN
7oLiZ8MStFj5vySyHalqwYvHS/OICBEWewLMnquyVX0T6mgzDC3QtnPYtaR8QvJ0MRwVhb3ZF956
AB8UuYEmX44QvCTGDlnpdf4q8jeH5fbU5UXMQ7xfjCWjfM+GqiIRKNBS/6rCpJNmebjeE2rmu8bH
sEy853vi5mC3RH+bnw1TSonZkjES8KolA3VSO1Aq3O8Rd0DI03o8GfHj/QfPUA5S5kCAdeJ5dZZv
ByIZf0hYnq8GTbZdwxgiyyrP7+ZbirWtqBzgUP5FqDoSKh7klSauFOs9CTvMygwd80F/Ts38QBl3
I0C30y1bzKItnAfnGOwNq8STij5vPkS6t72x7AdqnEgIOntq4SDviO56sg8xTSfmN3qZ6HO3zLSB
OIgjdYLm2VhAG7vC87p9wcSyljmyMfYtZv4g4uHgYb/aZ2v0kWwhAEm578TV471QZM7NpbFZsVXM
7Sh1SN6IZ8Jv8Zv6oNrvc+xxpY4clZ0QS3aKTDTArhv6rWidufTeASjn74zKCB++I2BuUiBskp3J
LXREjt37mbj3DHwhsy69mTpApibKrGiF79tYkuR/lFsqeJeqfQZRWur+2TC2jP3ooPQTHf1VAWrN
LHpiFAeHmcIHpp2lr/I3udfkTGJlCmG4qqRlv/Af/YbynA81B/P0Pj8b3eW+phyvewFAVeItwNUM
mORv1OG/mRwWeUGbxUgZgnx5cTzbD0XzUeXE8cP1Ymdkk3HkuYZdwkf+BOheagfyQSXvaROSkv06
CjSfXMUzNfJwCLstGWlnkMgmBO9EdRIheRSvHyHO6tCq8lRoM2B2S+OAOlNnyLll0rEwElddewKN
y60FYPEytPiXupphcjbq0QFQNpsc/ejTSHuYgWFfJ/ndtAW6YMT/iuxyQFwcxFDYuB98xrs8gPds
NhJehPCmJxv5Az4x8DaOeuiZaFOcrRDaIe1BJB4H0FZkA7uflx8KtN1rLlbOT1w6wxUZguB20zQf
sDKNzb93JAMckPxRqHV8RXiHe402nOCh3Vb4KHNBYkyGQGKaNWsPfSos93xi/TwtAUGcST/aI10Z
Ei2skjcsZZ3DwItQ8svWWiIaWm8aeQr/WC/ygKAzyyAocATdgO8ScAEfqOH10ZNatOxoAAT6JElL
qLFYIseqqcdO7GiG0Jk5nGpGDXopAecZXqUJjZFsUdiJw9FBc0SIGmOotjnJ1Yb1Vp69VH7DjPeM
TgHCxRfNe5H6L3FvJt7Nvkiuwkq96weJXGXcumdLE6teSnDgr1Rrpc4Dy9BbvS3n+9vgJqqBw9UZ
Y9Nk0WY1L6wPylwAsDkMi5/6U+SMgHqbsiL+YXtSN1ea01M4mlw7vd6HzpEkoQXAp4Lm7fNP3a+t
SRWND7A4lp1mnKoqfkbjomnZwcz82FULBAo3I8KiZqQTpt+0qY6SHZDcEsCdAphzuoeVZwA82/cX
/nkDEQJxavAHotZjXqM5E3uzvIydZEmRPhUyiUgtB7+r64PpxaIrAhKvm5noohtH+u8dde8i28+b
FLxtj6pjSX1CRFPNDQpEqS2qzUSTSrJrdMrDvZZL7XkULsjJrjxB4xwzzjjr0KG/k7+t+qOCGYuC
Ij86msBQHnURV8AywngRxx42aj547aGWRAD9RwkpsnB53VC1zK8gu0p2xgdz/Ubm1SMvHcC9H3Yi
dnI9Z1Y0IUV/L6kNh0ni6p0R7EUiWSWb0vTOqJnhE2X8X65agC+zrkoBtWr0s6wD/0pF0/evSFYJ
lPcOcLDc/LbWblntgeKS4N/HZnxVGsmBvEAyUD+TDGDEbdlb7azkuxzKH3XXYg7+QNom3mbeD3DK
w0kHo+7KHYGjVAuZk16YgJK9ZzVTUPlhJzfW9+S6W/N41gwC45aoMVnzutnzCgpLLOYu9cY5/m8s
L0kMrCwYLkZXCuq4vP0mT7YoZUkpLgKP2+trBXAml8MqOOsxBkzdxeGr1+mJVyYpnOYvJleqV45f
9DbKIHlKPWG63V99oX0vVBCz/XAfw8AboHVuxsr6zhhMgPSiKvxtQCdDs+cg6hj7KGFe4eWqvOJc
QdUQAMKzpU6AOnBRQMz4Ml4y09gpqDvTGerqWZvEAZkfkHNEgO/dTz+1GyvFVqOuBsi3bDvUWhEY
0nMsPTCZHGUjxYh/+8RjzW4ciHMeiBhdEVsJfHJR4gdmx+YpLOGeMtW8X99pke2pf9yllLbcszOM
12qfufK+sNNVD9SZMVOVE3Ikju5qAPa0vYbMmop4xhoc4lwenff3HRv7dMDNbvskwSb44CAWLsSb
2s58ok0Iu6V/TttaMqNeqrSb6mYhifM7qFKdI7QSz9eO4USsEs8KGSLNEICSon5QYfUZMhVe2Te1
MRrtPorfnDYUuW3UGcc81zpFo5bhusEhWpiANdE88yQyrv1CfHdxyv7sl5FFYFIRNwtfil9OQiex
+QsLlA7+CI297MxLU8qu2sfUrlaewiqVze9TLRMd+ICuzwjVajx8W4SkX7TIu4lRbRbA8QhICBxJ
ZXdYOLWxnzTVEh1V7wFLm9D2fUw2my99kogos0S7a2K0WYCBaFvRE7H4EqJYsZziUafnIAEuXhBp
y1d7ggnYoMphA1xVJFtg4738ruHvWCZLV29ZZsnvEWaH22TizbUANDUoohcwMwvY/QRT+Ify84f+
Yk6O798bZp4cqM1kqlT1v2aWctCVPheuf2GHoYwvAyp8dhRU3blyxtzoz7NQcvMd/8DobWfo5INK
V/bEf+ieD3n3UGlURxZQmUVQBBKzGN7UJ5abUAAR/wENe7WxlWT+Yi7MjhfRBMsixdDHU1kU34zN
pRIadzOqM43HGyinhBPh+OkkEA0mwsvwahqfoad1H/VIF3YCbwDGifrg3n0K6Ya2OW9fSwGQ1SsK
8s1I/lpCOREaQdSYMUEPg5SM2nxqkJKNMHJSC8i3gCzqwYW2wQCPe8nofo1QjBBlB8GkkoMqxZOE
6T8LHPhNgJEhMkFREJsnmiBJG33IkL1pKmRgR1WdyDKAg0KCVV8pw+tJkYnFXQ0VT7d+4gZVdVOb
daRcLS7OcX7OEzR6iAExD/VQ5zukDJQuUVg807JBPI5Nu4TMGeZzKJeLpJogcS/PrJeVptIoQvZR
WPykE/BHerF1Cr8O+ZKJTYTiaK0yiGRxvUDN5WVFuCPh0MwIunrhqx5NWCgbFllrxAaHYgU0njPb
4oAAgiBqEGJY0ZtlMofKNFviq/b4oIZH7WBIA5KDLUmSenA2Wgl4jdSqUoivgYV/lnxMcgNHJQ77
ZtBQuyZIlXMM49aa1+9toezxqF93zOK9joeH8sGZdiASPQ7y54N9fik3wmTCp+u4baPU2XusdOKW
DSqqGIgbucqJYsa3mkOnUbIYeMyb6rwoneLaKEZfL+x+2JuWgHCiNGP3OYv7tgF2S8SQsUOAUMge
1NYLJm56pQkC98lCEafZsWsUa3108uFQ3jq49VhwY6WG8cfRm1HKY12fczz3YK2L0VYvRqqiVhex
dvgtjuxWi5IBECyaB2wn4yxNTGUTvjpr6hsOGIxIj6sOsaes7fiqE1PRxELnnIdKC7z2Jxiog+Fz
b0A5J32O42k3LuvsKjkUzPJ/A4QGR7P7xm6ueVAXOPoAh/gJfr9TAzUY3rIbbJBdHc/7gOe3v1JS
8Kq20dH5eIEqbJBHQc1BUsLrIudg8ZyM+21mOF20rIIx6VrIhV4hNjAqWLsavYBb/sHBAQFh8mNL
oM1bgNc3BQ48qksCzECXayezAhj4FTCl0qO7mx5n7CG5FAvnnphE9o8Fs9Qz7yvt70WbbbHifwt1
3PEYnmlsjZaif5VtOW7z6KShyIju3DKLgNTp4SbrkkVdp36uIlKtqWBKtmGX/holvXqXeqrpUvtE
CEyDB0zpIOGpZSHWSl75twgXf779AFbNPP1LSWuEOpVqnGLBKUht6PwCR2P4VsyiW2qD6wqpWuF0
IhJEPbm3qTYFYzhmH8hV+i3g4wizLYDc7glMbkz3410scpEOMeEM77MoFeiDCAbqMGvt9f3TrI9j
jACJjFrDICj2xvpHtpySl9XTaZV7/n+iAWNV5XNsDqFQW/N9mcGoclgu+84f402M77zC3AIZJc8G
xgYVK/py+DIO/Jr8egFuCjbGFEPZjHtd9237ZkWEpHcNzuubCmSU5v6BYdJ7sGGn9FSObMITGDuw
Br8BMebICG7JChvHFAUdNCuisdSrPn0A6hGSzy/vVUk01Wt+PIl1y2cEUJaSd4xrTAbbAbUNpmf3
J7FNOJzelf2aaHO1ujkSp5YC3BR0Q5R3KR5hGI6ybM6eBgz83q70M0bBqjEoPG5TYMgSc+u5hJ5q
LUaTaVWzhmdPPWSbpul/tZeY4BqfK9PstX27RHIox+E3DFf7qSKGOIIGUiwAtgvt5ZwrMQt6a3Dq
c6yQlb7HLbW0W5dREIJfZDoaj16zzp9z0BO0eP8EqUcFQyseBt1fhIUiKlozFrL8w+NPC0fcmjn+
+IhWzjhUji8fqhjgY9sGti9ErRVJLDY7VEggnqjuEwW3IWMFaTwKdMbGbjdpAbMlJUA+tTSsyOIH
waHpapdcS1q2cluKWpZvGEvHxSqmajOw6CmGzbjG83H92bYNSHKM1Gk0WeAo817EcoTnQe15Ghk2
vq5xJq3fxnJ5CluIB91RX5SHj27XwpH7oAp8lWDVeCSPhZwlbtO5Zr2yrPx8W5V+QXPmzxSA9jwy
wmBmkggERDZMdOqrK68NOr3Vq86oIql9UYzdjxo3GJWBleQJWgNNdloVA3z2F9pUpLf3ioPW9osc
iBLdvdN0G3HXcrzPiR0oaeWfU9Tfheek6a4BLQg5fKHgAHW/Tig2SlFkbpFroMARgP41HOPzR4im
cBGA5C0xT7mxVksX3TyKhqV7Zxh4a5gsTVy9hDNgpq8Zi53bnnIH3w7XSpHxdl/pILbi3iOiogVm
ZbLRF78zIwdwdJEXGCPFHvBSWvNIZBA0GYiHwwecTHf6j7dFQr4mA36bIqfvRVD/QwK8SDwTTvjy
LOVYbBnzvInJ/bS1fCpcgpUprhAiWT31t8ZV5qlr4VgYPGxw3X989wkR/4ZiJxavHlVphYapS9cz
3L7SzEcgAib2JGNRcqdSq74ScSWvGrC0f5MCMWEFHU65NFK3Dp8mL3m4F2S9Wsd2N3mWHvp4/gXs
mURLHcISTruTSgkCrzB+00EAZBlIz8lOzRoRIgWv/3fIEBnYOTiS1ISMpDzyzpmVv7cEaHZoDx+8
U+3iW31JDd+EFOJt7gv8TZCcV7VlfmfeyCQ3wAGjyIoWpwG1XMzZtWobr/g47A7wkxe+Kr/9C5m3
445KI0TsVzJFsjiDodhQXAZ+9fH76l4tu0Cc0kUv9c9CXOE9wv+7FnF7jNLOV1m7O88vQiax5CZt
LKuFoicYXjgNKY4q5KYvf+PUezlJYlPOKR7AX17ZKAAuTKaSnSTUstbHXKIixL3ZJl8GmzxpJqx+
3CEha+2sgWsqc3lK99pQqXYTPGhkDtylB84j6aLclOTkU0zIoLzTn6rVsItEyJQOXg9/svb7LE0q
L45Wp2XgT7ivj21E99bOjI8QGZAEN36yL/v3lDRmtZO+JLkcHBXtUynX7xzsK5WcnRB0s1rD6xkv
wkIgblTDKinAOL61CnQuJsC6lYNYNOL2yfBmcZRgaqguufx2x638H4iZ7WLITwxOB1vNXrKQFZZQ
QMQQHGEpGfTbzeZf0nRpl0c0nm8MrIUOxV3oUOz+RGQJ0Q0HDnfN/TfX7wPhbefFlLMkJ1lHxokX
6cZmiF0zWpYX2UXkr7YfODQjIva9WTyLlW5DinyEWZuO4eJiRsjpueMUjhc7NcNIhI/WVEot0PWo
azr+0Scklz7kPYkTQS4q0LTlFiz9f9ZiDA7JlyWToOsXQzKx12kCBe9590BsaudX2M400ANh4/n+
6/BwxkwvsANpqJV54FPafq9K+DWzg7NsngMsKHlQTlAif8JCx+k1sLQRWywDYKWB6FNWMHCIJqE7
vsZuJr4qtlAJswGwolde9gFTdhz6xU6jUtdmGmKN+VS7kG+vEbOVM4t0COl0ATV1fvYPOwYJy8vk
XLY021R8MJ/7ntZvhDDuvzKRNjidlBBPZRhds/LLUKJW/dA5m3+LvGeSXRNluFsv1G2/6gvyr0XR
fjAjcrpn0WGDecMrdOlWPQIcAACjTnm58XaD/tA8caWLdCqDMRpNLCvFYr3ANqlMm0035Z6kyuLQ
tec2oih+fq0O7BBrlq8PBqD+D2eHmdkEDdyMu5ZFqIoTOWAHo0sNCCfTA1RAzb+OOVjxo+B/v0ZH
IC/auyooUQdSy62EB35y5ywApzYDYCuMVXFuwZ1PHbD3vZluk4hbDOTNUTbhIc4wNDIAn8MqWPzr
0KgMdvc5MJwOGqm5St83zcV/WL3O/FulHmDnoZo2t7I8WwVlHzHQsmf/1XRZBb0rVduCeMAAT8IH
+z+fh9AQv4dT4cY2cdBWWXVmnjwbQ4Kl3k1e89fEVbZJV0faFf1Bt5xzDzUFhQB/NiYElRQz2n7H
OiKV4Su0J1tP6JDJmfOrb6OU32urpG5XOtAMzb7z8j8quEaKdGnpDRQBsIpDqCXrJ+ACd4PYtnM6
9Dw0wLkn2mraRVM6xJWHpEDRl+8MwVSj5USOfMhD7QpS9dxyNtO2+YI0NdDN2sFxuv5d0rNnIMOX
THZxl2eg0bWQ7vkz4MviF4j1BmCfwt9635hJaT00Vl4kxPxDyIS73vd0rG5mrKXiP1rjqo/LjOhT
q8CM4fYbCjV4ahWVrwJHOAVuZzZvnH3dAMIwAKAV+KRcmcRDefVz74CT40JbAVQ/RtKZtI6r6KYF
OxNswmP3ynodktzXPYIv+ReJGJNJ2vH6W5q2mOD6PYVy8lq3HWQknE91pIv3hpbCZ0zFbOJCcEDi
NP/syXRjvWbNKaO/hunt8JY/HOCJVla8SW45SXygW9ZLRsAnCDMvfjzscv6I6SIWK5Z7kMNKTmMw
Er1/qf7Pol1eytM/Q7k4upug85S5tCWa6GigPsa/tTf3D2d6pwW8l2mVgrGFAF7L59krNIKg097L
kklWEzL0biXYsBH4o9IY2SaYterUt9StGXJkNCl701ZMPiseqbjjo9RfGipDZeJwMUu3G9KpnD5e
LUQ4jEyzWIgWgDnmvF57R+tfl+RWPNO7fE2aA4BQAUTYmfMzyLBzTHQbGzfEusaEsUg4op5EFHU2
T/NxVbf96YCfcBwLDq/oqDbr9d5/p2Vat/PpiB3RBQgR/orzPWSUnJ7ZlO8f8KgmRqP4p+sZRP+L
ZQujJeRE9RsjJBYqgkwmQK1dj/5kw0ZurlSYWe4jJ8A/nEUELz6WTozdypttDmq0gwrO4xc5nlBJ
jcCR87MTbhTlLbPsg+qeoPyiPN6sLwsXULyTb/wx5cWMyAVJlIg7yTZkIb+nrgwSr+jTpuAhhgSB
MIftgR8P7IOp+fXVUpY5F1zNEivufI5MznrNYm+LwYA5wbQ4z3aVOftS2Iw7KFIEd07igQUhX3hZ
O+xezNP9XtZg8kOkAMZP5lvrNZKTkG+pVT/Gi+U7+grEQ7CmYOWjm0VYHM/reUE9N5Lfm0fdrW+3
sH5niiqPgUiyI/UsHHTEig/NczP2D63jcFVW2yiHk88VNCzxw03Z47D+Lei5uxsm7KbMlRCGaNig
pF1pvvABI0ggI7xcUbqpJPPzsLjCcFQK8GN2onQMxQAsws+sShUGPENrHnXwe6z69GFnV44jgH+w
iVpRa88ST938DHXT9Mcfqozi+seuGQUwz6zOYNyo8E7GGJmIrmcATvZB1jt3o92HuXeolEoZ/oKa
ZPWy7COSm7PCcPVsazEisXJLOl2/RKGXE01PTgqQ8nsHGk63Jduv2g3uJaMlWX5neQHdjtrMvmms
BRBI3ZhR2sLrIHhVAQB/e4yVuVdhY4txJrQEx/+ta351GBL97qPrYVTa3Rr/WUDh5v5Vc3U0c06R
Y1E7Fgeip6uGoGSVrI3VLEBFcrYqp+0yxFKjMqmzFoRrLDJwuGAokFSPPyw3oKKTPfojgq/D4M75
rQ5qG9+4YUI6bpF5IHfWVyjy8I0N1lsk6g37UczCOcC+lm4E8H2X40MBTBjPshEtF/zFJ7/W/b1o
elVkPIUJhpbXm1htWp5bdhn7gSjas7vVA75J8WeH6W/1va6apdBlXiGYgtqZiGMPTMeBYqv21Bey
vHqpBUgUfCUHh/TuaPRDcXSe2NppujAKDgduwfw0wougk7lAY3UaHNomdMsTED8Cx3uAx+4ikW03
YwWIRwx4OpVCdU8kL6nGN3TYL2430SWihxLqvcFdsq60VIjztlk4CmYrpsTVxbEwNk652nUWbDm1
ughXgOkw6I1uoXQDgj88qHpfd+a+/E6pLkk6sxEuWvcuWYK8uA4CtVr/lPlaRWPDdE/UIqkWSX7P
7VYvyBNhIQ4WleigT0XOTX8MAgWw4t2QbOrnjFCYZlnyNTqjB9wsrkFwNpac8mbbCgV4XAN8ZRPQ
NDVZsXeIpiBGH+f7eE3I6/Ad3VCs8LyWl7yUJUoIg/1xjp+PLEONAFrav9NFETydH+0a3RW+78es
UalYcghnr1nwdO6p9w8qGsb9VVLxvnxO/W9HGyW9kH5/cXVI0EXzYL2JTpwKxJgauywIVi0DHDC1
T6oEUWKjBH0Pm34Awk9hOSdV9cNwC06k5IVf/ghOrKNgjMZ6IXz0GWvrsrGoYPnPJtueQtqzXVrh
rK/z69hBbYhAL3RbglLug96Llh4LVsxpXd9pZ7RrBlbpOk+JXqZY9S8GyOG7UM5ClBJatYz0VI9W
mnWzbAE3db2y6C93ro2lqOTcHo0tU0yxr7loIt4Wf4S0jhRWSTt5nAX8sMBBPo8B3jkoeScEIz5P
5VTto/5YonMeBPfg0DCUp0jKKdMupV7yg32DTfKaNO4z4Fe/KFlscTqvxRNeMrcPDPEYiCRBjdWK
zv4MK3xbnMAm5Qeil2DTmz0oUaBTPTP8RPnIrBsJBMLbOr1hwbtPAQsODpmPMYkmVC6EhL+fzjKe
BM7akzbPzmKIGrGmRipEV/djYGN+Zxbdhz51WmLkKWC1CjYcoSZeAl8AexlviWjdwA2G/ZQdFpTb
iCTQTW3nPM4s8YvIuz3+vj8oVd0sdk4XKrNiTaxmK4A+dNKAHqbKcrxJCHWRmoAUb4XXFrv8L6o/
eUm5gT2FbMNGAYEvhcI8aX4fZPLFY/Lk/KtCHibqM02VGsb7WNQHAUsb7qhnEt5Rj59n4xDQAW+i
Nfy6TdySuz8UC02zgoZnYKP5z6ona8AiPpEzV2fGrYaIz0lqjvI+uIZcgxReIjPNzWgvHeBUTwnV
HazCEe6Yg1sJ/Qs344lO5HhRlse3sPwomieelfB90SsrGsofRZC7C2z4nguGqhYW8+X9Kbff2oev
ep7vedOhurOoU8cpHfu97G/mpjZGKh7ufl/M6EDhJK8OgM99hSPAnEzF7pZw/MF6fgdtmO6QLRU2
s2LQvSP/IDaddgoYIQuZWJvgTXehz++rGe0rEFI+DZjMQaCk8Xc2cgwG/AvwZVLCqBTyxkAeXWdl
Nl2w8BVlOL305zvXd/CH8OO2qzb3KDTYV8TpEtSBNM/6+cCY7iGC/FdUZwyFNCoclTcr2pb/cNfJ
NMzbqPAZv19IdfCnmWClcZ7SHdDQnCGuUbkNpIJ2v5MXyOTu6v2JQcfER/wPDcvWVdkhnAj/UcNc
ZAmqH5RcJzdmEpVcYifZ+F3VgL/spJUfW0ZyXukIVHMOehHSbs4Vjvsic5WaaV6NYyboAttezWbu
BuARM8umQxQQV1N7BChMJuNfE/PxkUDoZ5SAXmevtI4sALnoPFKkbt9FfJvVs/zXck4sqNDY/8j5
A3OeWtCm9851drvQaMQIXkoaSikanwSE9UcLBO9aqBWDesfVCZZvfj76+GIeEs5+H95x0l511Ezy
eeK+H61i04NiynudSQkELjOiKthHBBe3oetmDG7u+UsLMLcsDQ2qUtirXql8L+Z2kKGsigbm8QlN
4FMzf6UAHMnZHDPolQTl+i+15fNkX5EKpmiCbi7hS22d0YGOSAHpIsqd2vI0oix+s6RFeUEXN9F8
KFP3d6YcXR/SB8g3xjslnU2ohIEu/gsn0De3BOmPjCcBLy6PmnuZmGBKUvndJcmoQesgxrxAN3RL
f+yJTFTWvtdWzz02w9i0o7PiOAQSbwr+eaf7hK7w35ikIyOjZLVsijVi86sLm67nxWKfhbkuAfh1
UKw+KV8esZ7CgT8ceMGgXyt9cGTxo5r40e8Sg/59jl+Zd1y09890G+2sC33Ok32QjkymAL5rXcIA
6TbYyk0Ri3/2r7VBIRJzSaFhH2U2IQRbvBjyTDNRRsfQ5SSOmYIEZ4BwKeM0HRpMk0PV8nBxiGiR
nam4+hoNhNsk8g70AzuoYNV6PaSNDtLz7gr9+cD7F7bxg8wkQi6M9fj6VleR0W3BzthLTiNH/fw/
WexOOgOcY2OhhnJofUqN0ED/k43Ix2F/Q1QFvYR9nl2rRvkpQ8xjYP1Km6cSBmljfLcTdIWLIo1m
xLsTn21cGFSB87YSHeSOtdlblwhLdZ4IALSSGO4qzRFOt+T7gxfibbtQf5e0W0kzoS2bD1xUoq98
m+5NGI4ICPk6ZsGWfUdZ10W/Kn1xr3eC8fp9F+Qm9y1M7x5L+Dz4NMJtrdXxKk2WSLR1iKbCj6Mm
Md8Iy03L7XmTGQ46lPEHho0+wYvFw9qsRiCzTDXwrgVixAKvC2runuEbKMkfblidy8qxycAh+gFG
6hVIYrS3YOc/jggS132rUzTfUiQ2qstOVeV4taYv1t8+W9nitCX1Qru4YJ46roB1uTq7S4RwMIz5
PKPFKnzOQXn4HfcqUbvQJPslrgyyZQVNUjlrDKqpq7+JR8Er2r7B5j5f7J9ACQV6EAc1PTmaRBDG
EbWLpJKVMjrwv1V3KhhbF68J/S/Y9sJvh04rGdiBGa7r+R9jWf+K3nrdP8XVC8Q73VIA6D/YLclU
up4rQrJxdEyjqbO9KPErpAVncuePyMoDQTr64j3L8ohXUXHwG+qSFfFPuHiV97I4tOC+3u4buqBX
7J90MdEzYQO/GEovufzM5QUEo5oacfjpeEKrb9SzljlOjGd0bQ1SKwzbpJ4/aQz8ZrI6s3+zHUf8
78s+VnXw/NPyiizFG5znDO+ZgDaVfuGLuA9stREVlXd4okUmdoijfBI/sp9uAqajb4mz0XnvXs94
++4DpuUABefqHWLdmwh/a+GISoh1UKeaYVZwPbi70ch6Q/DAIIuP+2EMEQRc/6FFCpqHtVc3aui0
MJ6aJNjzi3jnrBteYg9DTHWrO0vDHFkVFnmdh9xDI0Ip6Y0wi8X2SjdhyOIkHYblz6/9diIASwcx
+3HE0ZFdMzp5teeqoolLSxzeQrDa8TDfMOngfyFD8sfcRz9cVau7vU40BLtsoR0TPofuFpz6/P2G
4GpTb6qOejxNy4HHrOJGsAsr86Ecp0pZxGISwlgpV9KvoflHin5awsYQjyctNOjen2YO6Xuyl+Pn
gKKrXZHX6a9hbHYmTNpBpuDH8UgIDOit8oJSLFcV2LhzYa1Sy1F6MMjrYzTGWGdU8+2aS4fFjZts
Pdhup56lL00jBFJxPrKTKKXZJeFIKCB2iY0hz9UgYw5XMzv9oio6CJmN8wEVweYZdwgY706Oz3/Y
Uqw62XZiyh7m2xzKwumthG4Hv6lJpwCNLjpOK+hlNN7sVHEUZ+/Ew8N030o+7WeHiW8gdl7Wz7Zf
d1uaR2SF5XHZ4bQ9hWj78TiEUNGPxHBBLOJLX7q6ZUiooyYZUBT+pJUFM1T9PPZ81dq6+JrJlEA2
Kxm9UtTLOrEfpnESajVF1wzVOTyIcIjfjVoTqe3Uibid7I3tmDcKMPKfaIIbxS3Icrj5x/ife64+
MScpgK7s3Q8qC1wkEyaTrbXcKhKv2uSodJ5xCClPAhKOpRMmJexozcv0MMcrRCpNEo/0U6IvV95d
+z9MPYthBdLBfJuHRTG5uFmAbleByHLJMOiRn0U0RPEWdRCtIvfFER5OiOaxSl7caCdr3qLcgyqs
49sJC5oUJEduXBy+NiCMnta7WTebgajYDrZKK3218eMB82k+6E4PuQN0YiZngOAyitf2TWLL7BhP
O0qlXoA6jpef8sCv0fCQEXPTTngyQ/bzeJvZUVpmMzQhUKoXoso6Imf5KEiSnnmSh1xrZFnHEPu0
E64Uc6i6m6EymurAOsAIka46U5Pf5n7o1uuXh6h9Gr4vML4LeTHij0fvXl/j4zuLKbIG8fQjuNYj
VHPqD84+eC2/NQtgmPJoygRqzcJ9UECtU9L6TCQc3tw+9Bvk9W0DgoyykNlw2cVIkl7hHyfCylwb
QZn7M8gKYvvkBT27EneZ60OKnliCEdVUzFPM4kv9LR613OJGABHgIwKaFppVGbO7/16bxX/cODOz
Y5vuKpw2epoRi+vsNU3UVzoQF5Lxcg/ziihZWoUHX0QGXU7sPXZXwuqlKvO8eQFDiHntEBUYYAdk
UhdVQD11N4bNnRN1/EcR2VZY1NDa1rMSLH+m5wQaSMThjgApQf0f+wjCISACdbRryZtkFXx3D7TZ
z3h6Rodt9cdBP4ej6kxRzIkeBbdJV8HnA5xDm+5mQZXw/uj041whTdLUxG1re0SMo8QvFrtWbYj8
A/1pXKkUeRrGfSTKMIKPqu97sYyIQmMGhdbu20EWjP3Z4oxbX5KL7Cs//2ao/FgDMPFg1A2qZOE3
v0NH5l0StmLFg/MINOXOxWpeQXgACV4oFFZg4BAqFMQTFmfOtuN1N6FxUNuznpuqaUmQdRYRbSTs
w0YrCE2RAzLgGkHOZ2im1HLk3nBIUegoQSIDoVTyGkR+XNTRCd2Z9q+RfhgKBkvK4mbpgEUiEiQG
or6faEOLN1/nqUOEdC7kRfogKazBKoLoO5/mklKL8EwoRVNkGlI59VKmq0fAzc/Wo3l3e+Uy410Q
fdPRmzK9g5yDsVZl1SaklQdPbaSwOcr/K/fRmZe5uqht2om3OYhgLLsiaEXt4geStvMMjfako+Mu
dc/T+ujEWY8cL4x+l1wniAtc0jvtxM12Mt2IzdiV0enjTxTCYQpzh99VSYAzHg5aPSz2S/Q0p8zI
v5T/5Gp+Zs7YrrHtjFedKN3empKe7Dn2lhOt/PPWdTiACRMzvYlls7UTteJvRUsq1fU2skJdcmS3
wXH68lUHvQvqb58rdbZVdmnxh6UEFgWHFvl5btCeHauOB1xkbCkkeiMQDA4G1nLn3V8Sv89kzgM2
+cT9gOzthh5L5FbQpJY0uvZIlw3n+D5ZF4Qr2yOU0nvgvCIgPscW2qLo4SOe6B62wyxnIEz6cCr1
z5Dc20X6sdx8kYEaU+L3BfCiXu4ve7KoJFXYV69DpXQQk+nA+VemcSvU4l1p1nJSnNlIO6kVH8VT
QzjNflCm70HOCv6vc6FYliKpqF7pe80vfZLkFgmDubFOsnthWd60rC4cVbS4Bp2P0K17YL7+3zra
coWSPL6FFS5IFWcPi8wdqgHQExs2gYD7N38pWDzaxOS4cK+fETMewG0BzP8KrNlBca0byt+JETjT
AThCkxIa8+UZse2+Fzt1A/EOn89DVckc6/QmE+BY7SlwI59TKc0zoGrNdlJFD3o6utqSXgOXXFGJ
faJ+pcj5utaCGMk7VIyK8nCNiimQGwUB2tptaAQInnK/kFNem3jA3d5ANiTk/u0GCTdORJpzvvtY
bTCgCGVaLPp26ts+c39OPBBQYujBSG5UFCkmjqQW5V/KPsdSd5rabqBev/cCTmspErxBRALGPtRW
+o9f3Hnx7t9juYy9OZNXd1ieKzs7wva26OlXZqEGenQMxdL4/rs3RSt25WerF4bwhnAZPqjajzgC
hrSZoarsy7LnLkAQtz1F6cuZeLgwmHu/UqKYlgJ8Xkml2qaRd8i3l8/ZjuLByHAQcJsgvrfZTY3S
7Y73gAPYEZT+qTFRZYRBMC5Kslo+umc1IDnCymcNQhnFQ7EyFzaXTxOoKGoaCjWzk3xfvBswawSm
omPAm+M6b6vMHgqSLh90pXMF5q/Cx/X/llg8CIHXnVFOA0els6fNtPA9Y3ghQNWLs2egXULLHWjV
iWkM101YzUj+FWcD+IsHfCXU4MOP5+6ioqvnE/lTwRoqYpCK5bqU+PzP5B8E+TWoNfzwj0YKWdK7
u765FYq8Ikhr4SkZwU1fxBv9wOR9fG4VcfUOD3tg2ftqsD7Ele9qWcj29RF+xy31Qgdpaw+G6C42
C6CyrutmjXBSQRzbKwI/fNUk05NZ6d9tKEbeOnb35DVjFsyltzJ0Q9LZdYYxSDbhlrxXY8mUSmme
PdKEi9ld2a5LkyglcVKiIFWcTsRN7f5cr4OdLbswAeIs46gfAEw0ThWTT3HTE6QWD1LQBXQ++Tou
iiHOwg4NxM/qlGvJ2Er5e2CqyNLtRwuwH7EzN2rI0l7KRJjxt2tWqUJyv7kDokErCX/VLE+dFXYd
UTxPjQOFSLuxh5j+JcTVruIWJPaOMD2TwuifHuV+Eekbj7tC88JUCsYJFtBrNBv8PZ701Aro2pgd
y9xpXX+OGrUX8Lk3IkCAozw6AHnbKMRVtkC+j85+Efsmu0Eum3Asbe+92sRBXX3yRlaQYWRi1Ub9
T4yilWCdR76IwEk7QcPh0Z0k9to8fQjHfF5lF0J/JyLSHbbGeHiSk8I4GldumcoY2y0/4bA18Qtz
HocOwNcuotycGmMmZDTnfsRnROfu36Sg6WKIG9xMlAr4apK8fAVpgAgBcsV2Qarh+oDwhc92/dpi
Uy0slGPdxoXRuxMHe+lZbRD2XJQgFyaxUvaYCOazTMCTQZw2A6EqQFedEAAMgiy0hp95HSpsorFg
FqDR8w0hK60MXDlPa7G3L5HrnxRImn6c8NIbE4XJjkNpAu+YY1glRo0b219uonZiZCm3tG1svsn+
ZDWLTu5w5jpQ8gQyYxK/2U7pZsGIZVgas1era4nxAYgpiv8gLxwUd5MX2gak/J9lrZDzknr3NclH
vBYCebYF2D9UlZUzBJQzvTLsELnWOvbRPOCjY7kRYcT4SNszKzRroVf1MKxS3uzvKGwYV1EuB4OY
K48HBe1Fm8HDSWOf/aO8DgpjsqoEsBmMI1NqMU2h7ueXVZWWlhfU2foOcnaPAsN1vph33on5tGZG
5T4LMvBgs4xPfIRUD1ApOAwVho/7b0D5bNEPlFInSp5HVja3itpar4Cl+XyaAissL3HK/V2uvNrT
c1jAB8a5hBjQ68JqJ7Vup+y+DdhBS1QHxUUZh83qt5dVzP1a8FiS9UNRTsugu2AytbUY2RY9y6rY
sbyTOVnsuwtFKW1BVXhIIYNq6xCnNJ/mue2U1xx4x0V6KDQv/ePKtv4OgeAdX7cQqT/r6gRDEKx+
oYfcCJIoPWfwCOULushOGkZ0fHqqK/wDaf9z5pud17NOQa9Kx7pHMeivT2NvqiSFmqxCj0leKz6y
H6Mq6m+t69aMOdnlKyVXF43kjrI9fkrRTJaR4u3+GUyKmlkRK42oXNduS3jKA/PyUin1MxHH0WMC
TIyvLLY8MX3U95FHHvMk5LCp2j6564LNGqDszBlKoWjUvGWkv/8IuvU6qRQuP2yz8u7/mirUtezG
LycAz/fsmmgjcWc2JO6FFf2bzxRVfbEefgBer3nyy/McTDAOIFG0ve9H0Ngc7cew7OSwEINdTjpH
o44Hcc3cu1A6ZJ0zRnOyj3XnUOSVVrJvlZ5AFSbha9Y2joj3hoSYeR/KOkx56mSTchvlmJjuiFvm
e2mBnPVuF9eynNB3RN9DL5rR4KT8lKFMT3HBplC1d0BZ4esl2jehfFIwgSMfn44ehBjuzngTAz8S
LPnsXelRAwJ0ZJkEPlczeMB8612HzUplJi6pG5iseVXKilUlCzrfFl93wb0UnAY+XbF13Opq/yZ4
bMY+7KixWeniAKplEvxw7xZH4MhL/SfGNtzwt8HTsPHMoD9mJk8x1Lmfc/7viPxgtkdPB0onK2ij
JK9w/+Nmlc7NlFvDvUCC9uUHqHlB902s8WHmGTMr98z6zqhCeG+Haa+JMF5TjY4BQQYqotlUPx+l
KDOrk4SUHNEA399W50WZDHEK/HIPXsPMvRMRw6C2ZvTTPGdjpv6h5tWVmpqQrfQ6ts/xVnRf2Jrs
DouS5PmEFFYmrsYLp7i0Re/QY+h+QfE6Gq1sGvy5zFYk3c5DDfcOBES5EXYcQc4hCzUqDRRcFxFk
DYZc5oMXDd6u82ls3Vi+1zsynmBVlA5hCaZj8p7Q8jIMnTEIUEkafCYeEmLLAQ3zmVo2vll9aVtc
MaMTAJXIeo4gzos3uDpbbBFE1fa9waDwE37nZHGBz0bDwQJf3rcFQKYBGiiNCb0AwRzE4bQsSvGK
bPRZObZMTqFSxaSAN2mu+3Lomptdyt8uFgOoq4CNp3mUHX7rqDY6QT0r4zoONq1IJBLiYIHUFMEo
4pbjeMmFAA4msboncaTqBnQ18ZIcmvJuItRqhKfn5Kisq8SroMf4/RFVWFO5C+d/O6PYPcWbjuFG
nZHmwuiUd9yJGmjcGpO3HsACtDJR2fbXdYYE+Xlv1/WFlVxuWhKf52onIZloy8WwzKsABfgQT7ki
CjM31DyUQles5nHqiPhoHi9JAt5ZvHgkSMArhcbK6LFDzjikUg2QGJo0o7/q6BI5sLgw5LsudlqQ
jMt0YgcNOOtYrOkSEnPy+Ss0Z6qzgcXfsD0UVvQVh1LbxHaJB2nFYDdEzWBR0neTaNvWUbDC1QlL
Nz6LslvMU2KnNqsPXaY88Akq7sHaiNqxSk6VidgguOt4OwY/LcgVJ70S4CO5e/cwfB0Y7jSxCq5y
5mMjea7LfKg1Pz3a3MyWv1+9olCrypISHKLnVZXDgok3nGztTUBO4bWZcTvRyh+2h1/fjdES/FQu
ZOt//YQ/BEJPIsrbELOJnePsRxEcT3PQAIV2Eyqqut9ujCek/KVebAWEQ0waYV4E/qle6skuHf9f
7V7eq7qKMsfHij3sIVU0aMYFk2LOOjRWGsMvhlsQXj5VaV5f+m2c/e2cT2HCYpGLvtLDVyUB03UP
Dur6zMq1Np9aQNm5tpTv2GioIC7GyXifKgW+3mu1P26J/NfetIw68SaENTx+ZvI2uDANMVZwtXuW
gin79pMVMPZM7emdhBW1e3vg81pB64Mh4jJqe4/cgErRBfWQmMAEWH1T8iNSU3traII17pQfSqqP
Ee7T1FO1WcHoGtilMsErxPqMEUqdWDnVxTjGQXFbkAvH8/3iKnQ2eFXJma/P4WD5VEhR4JlhBbPe
cX0Dloxe/U9Yl4JntHLCgdUyN851TqMYGbasWDD3+UC3MmCcwdqzLLu+qzH2sbsggyLjaYMcvRdI
f7IVdCpJJDSOU9yoRVuAzxUN1BIHXEOL8IdETfpN3OfhONr9OWUkp5mBC1+vuMyHi5QCjIKFZYgg
nnZWgeesh2DCFS234avOJ/pAADnZPvVDXZuXiEE/UojQ1OZzLtaNOH8dLzeI35uVlv69ygSqUYy8
bQFPNJWO21NQs6snz5k8Zjsnssq4v0pQSl24ZT7NEvhOiaQdx8+Jj0KW99A+72Y2jJQkw6Hh4cRQ
hjJLqdT7+smaUCuqlAZYCjmqCKE7ZT4cZZRPwioIKpcltLZKq7xNanwKW8+mkksJsWxkuVDQzc6g
4yI0fyKhlcp5jkQqIYpLgRwQ5isdZ6AqQhLsg/km0atTXtbfGgC0ALFqE/NfpLeAGPos9NBVrJV5
PvWwY1yufXgRlBbI0GOLi06CvP24+5Y3X8QXXGvOSGxZaSnDbPIswg1MC/wuNGXffJm5CbAxLVhZ
+Kpobh77SKixaHwABp2DQ1igIFuUQi2TRcwa/9WdK9hbHnTlEjYZE2eu6cZPbEWy/RBfZDlTO6FE
41h+PHZc06emyIsduVE9dtnxUsswvRNuhW+NEaYQMUX23OzT77WkAWNLnpVJw1nTCkzAX8ImYU1B
0sYNMXDH6B8iMeEK+e/j1FiPtCFtMdFIsVYIK7TAvhsg8+nqfvCBERWcxtafFXLCjNOzg6gtliFI
6z/Jxm7bXiyCvsTRhCwIp6dwCw3ndtbHK4sjXd3TUUO0ZpRbXsc+t7CIGJNBEoBwYHa7w1NgasXU
518aSwZ+0PpQVfBKSTnK3JGI+xThco1IXWhmNyB5guojisSdsH1GK1B6iky20swHHnVV0KbXAm5z
esTI8s9F36X7m1hz/5enWr5/cqBkk0DsG0hvDSf2jo6TTWzlhHZ1F2wSpxOAIc1gKVdvhLGPdhgM
jo0CHIxBGXIXasK1XiKSW+Hc+noEsFyaIlUCEmJxV/81OsmteFJJEvQdMjLoMEEeZ+YeI3QxoIgb
PdB9et/V5S5oXXzmHxFUF6nQN9iXu0rfrAbBgvTZgkdEdky7I2F6yQAOr1cRXhLMOIpS4mhi/x/r
FGMbtAr+QnB52Lp/dgLd97LfDmhEY1Vu0jp5z4IU0/7++jpEkTnP5vPaprGyEqzy+o7h27UnSl2x
7Xa00te1GbSAT6dqTdx3H41HeYwUdO0ikq654o3EY0TqsPyZK3NlvmZ75bKc8bxgV90cZL+maL1+
TuTLhkdgjWl2zVONHa3CPhDYTXsouIwg/ylvg0IWQkhMUVQe7YscYs8qyObwygl7CjqgDfAy72og
tX8A6HY3vn925cEJcU7bmwVOu4uqzIeEfid+mISKDyXKrEa6NqftSzpPPe4TVuFTPdRq1fSDXHPR
nK7btZvOjEoGitbO5syETZCu6Y6Ae8OzTU98Z1iHYzCkAT7cRuGB85NSozraiJlsFrTaEuANoJ4e
GWC+47vGRytE+mRIvohOkAP+LqiO7ovfqwJTQEuMblWUlg76V6bWHUKUSd/miFwvHh8JJ5nIiXAP
GWWX/VQneANksKwMbYvbk4HRFXgAZthn15jyFqT3DQxhLyfMLJRBSegRIl8xMzQS2hun4gGtSW2R
Y/tUYHEs/hB4ChEZejLdyfORcag7zaVOsM/MQWc5jAW0pmJueW+lJCtszTLv8+FARS5sDbIo/3WX
vke/hEGpF3xw3ed6eqoRyzuAVvhotOsvLfD2Ff8OMv02NkDd5zEyUL9wFErtOJTbHgAtaUoTpLKt
wd4RXBrfWloadXwntC1aVleFL5n15GpsWtmNmnXZ5ko4lhL5Aa/ohkbNxX/Kl6S0YVa+/ZI8RXH+
d8tiJ4Ksa0yADpXtKfUsZAbDkDswi0JCFWCqbnD6/cS5KuDDIJphzIcdKsiNbAJyCEi0aFAL6C8B
hvKvLdLZJtjZHrdw01j/fMO+EN5dfxA7cU2K2kVpeBtVvOcjfgfP0KF2xWN9MaIguEIB8D6F/6o6
355qmA7VpRKbIORyHW6GleMAyOHh7rLiO/agw9WLvwAqQGH/gelo4I82WdEx/D/y+iVEIrL61RJz
9VL9LdQg9fhL5fNeSFVvXpuOcJAcWxcwyJ3q1uiafMjlJi4gD4klw4QYuiPIWuYqrAyAYp0aF2M1
JodrGxt5904ShajNAETWNJ0yeoEhCuV/Y7rQrfzScXUJzGlXmLrgcY1AebsQjW+P6/jibUYanXKP
Px1T9y1KXgPiNWC4hOLtiTbG+1nzofZqRs/5TK8rBb8duNunm7bS/BFlmrPbodkFHF/nXuBLZR5v
L8ZU5DwUG/UmgiXD4eTvw3HgKnKXVxfYCtxT7XZGeneQ84yhyHQ86/EJmVMTdogi5z7Wyj9DJqLX
xNv5DzWCZO5d8tZ72he5RaiRHCu8HmSPX7dmwiY9+dg9ZBnww+CJN6fpoH+QWsukXZWOKaW07CQm
Ntva7xCQXWQEFkeTS2qg+SWnplUCX+FaMo5ukh6yea0mAsKrB9jUgEt+zrBXahZvXs9jEj5Hw7La
8TapjbQwz6bXA54hkL7Byc07dlCkSDkMjjNthGcXIHR9rRFgrc0y62ZVrovZ2pG7rVe4Kb9jd9Aq
ryvfnmQCBB5zTS2aLYfCw07x3EQKe+N6fngu/sb6Wguf8nMVcYQo+IYSS/GdfKqocksdaGv6SuUS
MMQw028Hzfb2B6sy8isbl290ajHBUYWrbpaa19/MAR6G9DKo3msoi9qotibC/kFIPEk61rl3RRxl
EIFpYV4C8nHSrAjxdsiNqmhkMUSyQqOniYi6g3CbZHGfXMGLi4zhbexuym0d5bpSvXRMYBVsTy64
jW9Rk6VlVzMOlrL/e1E6gMwv0TG9snI9/+Ni4RKCHEBARQjRusEQbKxAv9vscWSLzWSIwtriRUAq
dFhceA10KaiZrcfZyqeYYySS1pb/UWGBb6rgQO/QaQLZP6TdUeLSZcaKJJTSzfNX9jqWNN/KNajN
NTChM4QjNQn+iifFXVMLoH+f9Itsg96b3E9cjhRW+G0OVs5j9pKCwc3xq6XzR+PRFbIFIefGeLqS
+ba+w1QWcplQAgkwN09K9LrMZJZwCWjoEB+YZwL/PDCzfDtZX31b+1WiU0e2hIUMVic+WwFgHtal
vu1xXMaK30rcVqC3ZAA6z3zXpRjpi0LR99P3jS9kRmB48oURzE6Of7lSW0SrfzdoV65eaYbdNCjQ
QjdOc5w6bfDOVqA5n6sHNDUcA2+1+xkRpDtMRlw0jwlrOUkpwQ8CEUHT8z4RPHgImBEfUvhXq4NS
pcQT6Xfc7D3zztAkYF+5Lm+Ckk2WHBF/NbWRK0+y5KaPAEwgw4ec5N5dbJaGuLx22aCLK3kqeQSN
r28JC+XYunTwh8xhluybI5K3BWVvw0tL9NANVKbgIDVIINmCz+yOZeSxvakeminLDUqf7V2MtGpf
aQXh8dJzGiLpmk5mwTnpJAJqx/I5+dU34DArfmx5Fjd+ML21gFwIChzaNKy8XqX82uaY0eMwCTSM
fIYaMycCxspXjbQ+ni4lyJTLac8kkcKQZ+dk+VOb+fzqK2iUQ2mKUD+uEn8gwdgYTGTPr/PyyLjE
sqLP1JBwXpl6KeX6kb4iO/KpF38TMYpk5T7Sd4KJCmjpoQ5vY5Xwsd3aHbZy2yLcz5ADKom/p8wr
7XGenGBQUCUU9nlwrcr9VUUE3BzPZw91A5begtJzOsWhLBBn3jhAm7UapUPS3mvDgSJtaQBfHm4K
TjkftdJyaP/odm4L4Wtt3gHD5kCcyrXF4UixMZsjyAckiohM5PXZ5jNgso3yGG6sx5IzEmTi2F6S
wnklOAf7N4eJdrUf9LZKauN6IUyGK/zcA8QYVixxzPo5CSeWTCVNgcT8l7lxDNWIyljqt/OQlXWM
pHDVrYSWpQjuaaSvabd5a5KIWlDQosu6iDzsPGDYbEYaj/0tTLNgwlS+mZVP+AFURsj8zLPjMVf/
SiyZxH5HSfzpzVlVEewvTxyx33n/cC1kseODErPdH60weK/6OttI7Sck16DduviQLNtFr8cMZUk/
7sLQyYXXmM4dLOsxf187twREX3EI2xMEW+tfycdoJDYU6r2pbsS24C1Jd6OPKj+U14t8ywhyWj+8
JlbV4wZSKAA2+4tQjqnQpah5LrdZSaOcnY/oY1d4nmV1CUMF7X90t+9lCM0nxMzqOLB4dJ19llfx
3/EOxhMu2oVUIwPKXyj8gYKimTfk55YJqjc0RRFoizrt37AZtWXy328HKLBd0EReJCoQW9p58rZS
wzkJF+MOpqJRx7/IE9rtzw6/brXmTloPuurX3nRgJoFlM5y7dvtXCI2FBzxG5vw2sSPE+leHWYBd
3FLYcSb28pnOrxtZVfym8l4NUcgYzck3TO6iSXVJobn1cBS2kCKYJMoZ45TMiQhLYPGGUglcivcf
pOOMB1f9oRZzKNHxwyd0KEw3c87PYIQFgS04+pnGwPMo60qX0capRCOJe5bd2XGQLg3777RHa/JC
Hiwbc1ESEJXPY3Fw1wDEOKqokqOQ2eghbou618dX4ZTl0c2cq8KatuYFfTcZ5sRO5WZrtnBqZF7q
EZZMj3upLXpGkJsE27Wfc0dsg+l3kL1FzuD44ESk0A5PSIaqF2SGJ4OnyY5WvaMWEujwS6/IE/pO
yZpMVFMTHeVEMxxNfJYtbRYy9a/NuLosfLKBlJkk0cO8+mvQCZwbxNXaTp2L3us8IL3p4uyBxcnF
/odBJ4S0OBg+B/VNSmJFJ9n6mvWyyvFVfIWc8fQj7Z4mz5ixlZqzFTKYLkcFTyNLxCNp9dO75BFk
9WRUvaQt4uYVwXY2UtHP5Z5wfC5BxMaTHs4VfiRYzc68xO8djemLtbOSe0lEc6rzMWCXXKmwYavf
fVeb+ShKAWQGtqWqSvv9QcfkbdJBEK2bNSA/66hywTGkDAdtT1dJi5wizR6XJ4G0Q5pCmbGc7Ays
JEDmu0Sl2d2bhE+H08fT6Mba0gx9zpI7ulnYFjqWOoAcygu9SvyS8y3+R7r86XRQAN1PWeupiOQc
oSKNFSYT2jtzOG4YOOLt/4g5zTQjleDrAIZtrYSm+bhD0Cm6ktOeS9QA385rPy49KvWxKfayyFjP
5Xg1XocZH5pGCIOUM5MyawhjYAuzQ13xY/U2MW2nE0Y/VLVED3Npzrzjf7meaRrnRLIzf8Z70+JZ
V7wwqN3bdGTY1XhnFjL2+k7NOiGszqWWN1W3ntkQKjsCxFXmywk+PPE01mGOvva5lj5gaU/QDekM
R/ULc+KL6cGr5zpA4GxxqgioH32xHNISnGm5aMr9Cz9fVsnYI2xCA2hwjRkeh8A4Sap+V1TC0dF6
2lHjeI5HBMBq/phkb3xE0sX4gLPMRYEk4Zz+SYSkskHGLUsdamZgOay798PBC3OqxMKUBoRaZsIH
6Ph2mFzgl5BX0b+yJsFDGAEIr6jaOE0Zr8T7nEcWvGcOalQM6+4AtNtZp0CdZWuIrcJwxgnExuaB
ONgViErAIdE+E+3VsN8UfAf97FF/aGa2vX0fH4mdUocy+9f+XHWNudcoHJfyLwTYAqSev8Jd3YXc
RxD7tOHzaDTMwjHmtwak/w+uRfp74k8m01sDeWI/l/mEGmQkjIWVcHd30+1J6l95Sa3p8luAzfi+
aLgYQGpS2Nk7MA5YfbxS1DJLLadVoMAuxQ/3LKq4Qk1pTItNpAm81XLI9CBx3R+noAuYH17oDuuq
DXmXLPrTSTLmm1CLuTHeEUtNPrMs6Vgzlu6c9hVnx3aksGilTl70bXVjzZpxyvmx2NqPvv9Zo0Qc
KFRDwVObx1EQ5iQa1lncZCAFthNHZbBSvGZgJQriNOTsYVNsZNF6IMdTivczXuR9gD/oTjvzSr34
ftUeI+01sYuSWQWyjpkne8Us7AVA48yidpo4kZPT5+EjUkouylEPrWKv7KRL0SA+6p0mElrOsUrT
CQk7tcr6XnZe0qISQyEl+WPQVdYxUyW6WsH9Q23INASrEwkvqo/AJFVBsYYjhOJFYqpT3L/rVngn
GjksUtfcgh51GNuGb6TuBYhXMezAgrADFH+z8Tdhe+SWOpNrq2xDf9VDN4gq8Endly9GnweTageC
UhXaP4plEenKCVduxf6lHJRoWQqeYLOoEF3UEUlOA/DTbQ8fsvt9Azk7vU2zvgGTHJpxOXX2QAJ5
w+5QiKxt4FCmZYrKUAJwf1kyvvjcVUpNIlNmBstRU5bTpLjYIDw8IYyc1H52c7TEhQeUxLEhdDeO
MZ36HrVECV43SsPjCuScDO2HkkdA6ZGa1v8+qSRtBG2glL2hdwMMnHJYDyfMn6zakpZXWEuOezQM
a+twpOQ4/ZZjBJEgm9JqfMWwRaAQ7plJzd2OQJ2kw/yRt0vC2bQ+pDYSeVnK00PUkoMVvFaVaDgo
S1hXlNogICNUowNU4zZYvgLV2vmJQscJvaT+IkqibKxschfjl20gcfwiJhfcDxW6BUOuAGDwiOvI
00C+yNb/Qi3h2zU3N//MleLNyAaMbr3TLoAZJECQ7lbpMFHO+3qaiSmsYq/kMCJxbS0xP5cahac5
6cGzFSTzd7XfwlIBNTpefModCwSbP+UVJgRqmuXPiSMrkb3BVYs7emQWz7iUvS3DSghctszQk2hK
tpHb/XcsH7jEI8Kkiwxf16F8PpXSKQZP8HJifCdCS1VtsUQVjAZEbcVc4O3XUXyjA/cJHlavUpYc
XYv5r0O34xJjvo64tS8n4sEh/hemPFL+iFNC6ZlGYirEKBAWXH3/Cy1TQ0yuehSVppqEZIclh4ez
x/CbPHdkNtHL3G0luxIin1nIkzpjKDIqrKZE0TvG7z5XMv03DfhfcsEJJqGuO1ZY7tjZQUulUIXC
hZvjqYS81gte+/1imAmaGcC5SHz/uNs6U+Vuisyc2MjOZsoezt1pcR+0phRBOckLeksBpvwlM10p
h24qXAXJvr7xBTQ0537y8e5Fq5BFFM2fT6UH6XguLgIn7Jec4eB0LntnajgQy6qepLxBA8q2Mq54
tfIbk4Djrn4YWFHLG9XIIHymK1qPTDdH/JIoltn/uiuiYgHiDhoXCSS9oLFhbhiUq8t6RaaQtGxG
A5r9b/8RQEqQ+yKszQanF/4Tw0rD/FVSCLFifG7zMN5w/9dXqFsnFOIrciVXieon63cyRAPF/hJj
JgrXYKrB/r3sTyEBcDVWW04KaXGtReKeULelMNKg6XVseGJhkcwthJCFyjGrvlFoSv4rRrTA7sou
IQjtmgA7gv0Nx7SsFbEsvFG9w7rTHGLQLymaRkj9xjHMtQiE8dsWM5SzhpEhSNNNeIP7OVGHh5Ad
+Eisc/hdWsfQ9TU6kNxJV2qI0e7ANHWBE4F2XEMJR1l4AIHSwvuo7pGvI0hqMBnI/nb16AVhL+xq
COp3vti2yGZlu/c/Q5Z+n4sXXDgPR2LRXx2bH/Lm6ntVgyYkhliVIuu/pDJaYDYv57iqHfB0Laj5
G0MmLMrEowp2SuiYOCbmYDzpiqQFvp/CydJ5x2ZN2EluLif7Mv8w3rSVfU80ijpD2WxJ/Xd1tKNl
wqofMSsq0qdr8zqZ+LdEiDOveRN45SNPZZVkt9Pb7i6TaZ9dbHseS+cflxYxfN68DC5KzFuiBshG
LFiuF0kzbfJSZ/Zs4grU9DxxFlvYBuuIbwV1o0WzlZ6T6UYZe7Lgcs2YEqCcEirN58GPAVu9CTSL
rqjty2AEyQU0AvdsckZBFNOoSLb9CN0Sd9k4IEdL+5+zi8D2PYgSkxile1T1t3+j8doYVStbU+S9
6nXr8cRsEmOgVJpI5vmXSMMdJ7l9bqOiLS4oHPEy4Rxq9+JDx5PL1ij0SotuFOZFWPByVDszK0qq
v//4ggPqicidifdm3yXmoqYQpYF2LCoDtVU+bItUujUEK4BzkFo8LSZDXbp3jT5JYzsvqbA/iq2y
V0Bjwl4xFYF5lgJstmYYNFwENA5EUYgnDFsrXzjoMzHAwJA5NB0p/MEzBQCjXVXFnpUGEwZJGCo4
zoy0mi+mWbA8LXcY1mmGknkGvKvc5oFHsjk15wY8Y/jN149uhVYKqgG2KL0P5rdZiZzpjoVKquIe
gya+nxpa3dwCEqANzu9vllcGmeVyS3HYUnCgLiW87D7yZkCZA/T+5/O5rEl9T3NMpBSelNZyaVPu
dSGQzgh87AtkvYz2rbORE/djq4IfmJMJHbbWkB3xCNf81xcnKwUvqqqP91kFnaaH5sy3+jqi/cOE
EeAub+PXn3Qm5Rt1A5yO1M+Jj+tLa9vO5HqTgYxuNmS1k0ctwQEJ875QIMpbilhSHBU40Ok6myv+
w223nBjdRYi8SKsp7tlMbcyoYvQN9EPhykcwEB/+k7BuwIwONdVNi5iGYL5FS7rcwsvJMpHTnUR9
VlUIAHrqnEmi4+IIm7Gh11aiOjIdco+K1Hi0jxkI1GIysAZQhg2eD8IAxvBdZ9nz5J4J2wPmVgjB
ii/4nBH9f4P87kCYWfS277dN0Rw2ZN9Zhk2PnBulo6C2PmqA8jUly53zZP5DhHzTtaLDSy7PxTEm
jTKrPP3SsSv+sJLUsjLEzckCb8y5XTY0WLJtjZXiIswNVrpL4yidj6lLfAg1DKl/r3x9Lkss1GR+
3tZBNGtfRwIv8rGlZWvHYMieziOfPJ/ZoZpXQzbJuybNknFitH4XX6PJgN7Unc9KoV646XipzQgF
h/BSuKzn/ZheZrX0nxMjZfDLigpZBvX+FFFwSlXNkCzAFHaMzr64pudDA5yg8wwwaHzRwokYT0H9
nWC5NgB7skHsaNSA3bYQjUX7mL2e2MfONu2EzzO4g16VbDjBJ4fM63eKNQwsJQy/J3wZp5xTLNL1
aZ07hV20MwDkMojueJp+uTsMM9x4JPLFTmtrH/9k8IlLkVMZr2P9hbrajkdA/YGLut8+pCz9wgy7
baJ4lBG5XAI+bTZUFs7lLrCId2XzNJYool5Cg+sO0H8Hdzyzw8CkhpNUfyiz+NAWn3HZPt+Uzz8O
nu2QrX+vwqG4I9dy3yUL6te/eIYaZw4SU7PkHsIE64MLnFCrgqeDwVrIVr9vfBEp2ea1QQm3I8VM
65KW5wvXYw7V0OLqTkuEDRR0LfEW88JjzCgcaGa88BBejC3ZCgTXR9OiJu6hNKymZU+4NuBqWlwi
bqhh3E2nqs+ibcErYmKDc/W2JrPv6tZJBi1g7+k5GmdYcAc44bTbd/JU8hDxnhdBnYRDlesCrxxb
txE8Xr2EhMKG2JmslOppkLdbapU5OCr3X8kRHMPTOH+LJqpT/Kn7H95JnJzQ3PpBZr6QldaA0LH3
O1RwWVP+m6nR8hvFuJTqEpMa0MI0SL9D3orpDtZwoMMtC3v2lMioN0MxN2rUE+Q1wuEamt5E2Zb9
z6qVJ3Ba3Iza+/Du04a0GDKA3i0y1/luNj8e+Pk/fk9pjKzvFMz0RyHxhiQIHQ5bXk7KgrHIFaRh
SUJaEND0TCwr1bqqttTIKeFB0+tvfvWAszv4wSclYw1A0ak4ps313TizT8PbjUdxgrFYxmEUIiLE
ddl7ztt/Te7BBplxr1j3WOPNAe5O/a+zS8YxqIVFYp2Vdmdz1mXE5rv8qxdnzhpwpyue6E9L3U1S
FeXMXi4kWSqD/UGdC60p/buYvePxhEJzGlEhsHC5+vWvtyou/iRHu+gfS+MMrKfp/sD2V2JgcqbK
zTWvJrz3Iaxkfp39i52HnM1wPXnkKi+y0iJFhy5P11mwmuYp+WO4qDsoSwInb3J1Q6BryiOUu3Nf
9SXrKdwxz4VE2c8QZA/3EtPjO/Q9f+CUaCwvb4vReEMypHU97dE/457fwxJX97+0C89ijXVqMkLq
aoqVKG+wRpgnH4eUF2oaGmUh5DBIjKc4r+pqzokvUTq0cijIM6CiitputUDjr3PY/qPepKCccOyG
+y3WRZSWlTylLkEfhG4MC6shMDSRHdcGWocYwHKrml1GwWtc7ClaCWjczmfDzOzm6k+DHMaTGtwE
ynpYRq5ya+OhkAAXKeW6uneWbygksIr45C7Ip9K3m6O060bbd2dRrI+Mu6SQuJTCYB44xDzqw4yl
4+6XW9kCkOJTr6x8hg1GhIqo+SQ5jSo4RONubvexvIHTpf87U9cnLmuGZ1DviA20o7La+Sjx5h2E
8G56bEVEXyXKQWPz5stn5yKqzcvI6I+BRunE38OCbBK7IrfN5gJ66Qqarhua/1nBbn0sRlBMFOh2
DDc/pUuQRmf22S/kMbTC8iqUKPPJ800iErbMhiq9vDilvkqnGjkSLlSEzNpGQ2pT58BJv8S9Wfem
QB2N5lK55iSGhnpJL58+c8o9MXZWYFVeo8aoM0QMAaoWyQZIsg+wPlaxqh01HQTW6PO3e2ECuDia
2ecOj/R66wHLbb7qFwApt+9/GPGeCVDe/6WiQU1eU/htbmc6AwfJiTXhfKhTtXyDXhiCEcEoDvbe
Wr4N8lvO2JiBafSQ67jpYmKBP11RI7MZ9Xp1aXfMht5RedFZebOaWD5sp30AmkEm2mUQOAtrbpO0
OtqcLpnAljN60EOkr+DTvA6ZGCBTGca1V0WSAr0ethHe9fvYuPxz2nXp50ZLj2OmkFi/cBX6S33/
NfV6/nVTqmXFAzuZxGuOaHIFmYSDLqZjCz4QTOE2KUwkz++UMiNZFxicg2tTA2ngZdrLhWM3EYdA
HJKVKqcnFypfXI6smUiGeMIyYlCC3dHs9Ud4Kwil4t9KiLOvMO+ebzb/+LJjUD1+BgJjG7bVvcc8
AxAWew5uvsqkeGKBR9j4+jFzvYDUhJl91JP+ftCeaXnyknMzDk02r3CgYzRUVNlkN34zIGKx4RWD
Yh+g3MluMfHrztvpUePi7KHvHC7bic8gOMMXp27mcDcpD7VrHSp3Rr8ycX6nQ7gRtlkKXyn94x9f
ln/7Gg0xPWKFfSdWan9G2qOWxu7ZbHek/3b+1YbA95hgKJjKCPub9YoHejCwT/uMxB3+pLGNp5xn
LN1R8tjMRf4/Nli0419p3hTiIlZhWECbShVZKRAgrIFOHUby9MGeW+XRz75lEuQizT3wX+9vLvsV
jbLsfy3kcOfYPwy3Q+XSmmHLmpWIrrl5vAInrrhlEqTBmzW15yTH3QfgQ1SjHlr/WiKxvrkuUuWz
f95avAfQK7ud8BjhVeGkjEnjSpKeE3jO7dIbwfv+bETz101JOktJEx/dt0CUUiXdGnFIO+cuNfyl
8g8TIhM2sQTZScy5x5gOnCUTL4XZJWbEVfwDtFz0kfYYfzyhyaGIFNwAnmXxw8lj1EHpPGJSJpu4
O/UxdVJ5RKU8Yd93p/B1GwLmY+PFgwbmZk9xESahDnFy6Cz+If/Qw3WJv0A+JM+fbWzv9PBHEoKb
F41UODdCHNCw48hwgwKl0HE/oZg3JV7FJ6xDudcbtkcHkxkgqSQMwj6EiFYKoDr8NyIHU/HNDzlE
lnuw3vnqYlh4GsTIhhWtZrBYEbFVf49uuCjhTb91wT+V0sEuZq5Izhk+gMgOSa/VbxCtR942BPTD
/Ux/xvD1QLBVylQxz3BeeCCqNxZ0Ut3EqBd7/ALsaY5UNtW42wJLf9KtJfx6iujkEUv+8Iju+Zd4
x000XYYAdbzMt+9KJwLSErKqWJ6VyEse6cc9X+di4zE8Ld5FfddCFAPNL1RePJ72QtpZLVtrrq6K
TaCM5mEEEAgtwf3LhGzKeiBs/RTWGEPF4jg9nczZ+vQdwedP+C+7/GrzDqBdv1cPRiBKbi5sLvzR
tEtTnsnKXkoMr2zD2m+Nbmy2s4LFPKSJZxPB4vPxrJ5b8uRRjOSNlPDshjIAXi28vVVt9xfeu3XP
5LtIt2ITQJjHKnRZtDjBAVEkGBz36aXqIt0C0hkV+qAh1A0LDGEffJiKOShnG/iro506ZWBCvtqI
wZK70IAEXQrDWGplcHbTCKdK1xPz/JAi2qMgDxXAnB/Q0VIZ58rUE2TYOmTKb5YleHGx3qOIZfU2
dg1GbORVVxllGKGUr4hY3pDj52dztnH5wu8GukXTPNpmfBcxtVyHjYHGZxpXrcI3KVuslJu4866D
g4vzWLaLXJdqbsT344BIyoUlxSprYek2F9qo6alIsSRwhIS2+v2sFCcqGAYT3aykrjOi7NECBs3o
v9J95paJVcG/0sGmArD9XuOWJ1+F9uSwMCuP3zyVklQxsFibF1J04snuqeJvh9UgjaK0ngeyXoxx
1BbeIqZFyY+Svch9SqucvsMt+BGu19OEfjqgKJUTaBHVBhbTGrJRH/B4TcJpNccm51QgI0cLoU2t
D+7puj9yFywygv5NLAu8Kml9diYqEyST022G2irYEewzdh6Iu1HG0XdVhB5rs9/7r/lXP3YlXIpF
P5HC3Pcid+XeKpiUfhBNl6sBllaPBnTz92tqc1HWlWA4fGJfKSNIoVIFKTynfXNrJxrV6EtSDbYE
FhSMJewKmnSUBnb0XPlHtp6+P/kYn8WVc6dg6XZH0v2SzC1Ae3E0uDAta6eMKsA9P9mtRDRHqvgJ
sc3Sm00awbUuL6M6cRdN2fz5N5JFHFZHtc2/dCU2bLJbQ2OvHn86uNgEw7JCyxD54psCqT+Eqq2D
i46ps5nMVhExjdux980n1CD7kEkAw0mM+dEgSuR9CJxfZc0gyIM5yoT7aWrXOMR/nrPTX/QSMidD
JYXWJDiCw83IDA9UxAmqwUCVKFWKHSiqdzswIJW1Kw5+1gylOKjgyvvR3rpK5yM23COE5snBUdXa
EsZyz8fRgHSYpTRJ3/AaRwtTzW9fK/Q5YYfIt51IGN2kTjs4BklmHY+JCulES+z0F870g2E7bS79
lyNIsK0jURn17+QbHNE1oS3gzeSff4ZEjrSbiDcIbhgIbTLgxTXWD+G+o6mmTy/kezOBQPyhMnwQ
PpIJVSggWqWhzE96qHKKeXXO18B8/ZjbyBJ42faZuYXv4zoXGM/BYQEUsMTAb4UE7EWUY74ykqP4
JLuVBeZn4t5+iVNOjIlJoZ36/NXaffn1fej33jWqaoUVet625QJ+h+IotX3avb7RR3ExxKCHmLTv
7Ah9r9ie8G6V06VKYwhm9Lj3uVaAP5DnkGA0u+9Y7rOkEW+EGI0KYp7d5Ir6j0wqlnkGABuaQzgJ
oTR5QXwei4PItbDgiv8qIjob27Y9Ouoy4O+IsvIhW4ysmnp/eAfUwKUGr52pBsIOrIXiN3IR57xY
WshVZOZFsPOj0gc42OXvsRj2eo/td7yNtcO1qk3fYt0U4aPJD+51kBmuEl17201BFrWiEVCoNqQS
k70sQ6uGzBQ0EBNGcUglCUp6yquhS+8XIMEy9yU8LRvN5nJR0WShz3GJyx53wu3o+N68LBKBMSAy
AxfyCG961JTq8m+XKJF0t/s/e2d3jzyVBLLiYO6zcsHp9J7gROssth9PI9RaUIVmO0VuPvQZHGNK
1GWuMiiGGCYEb48+jfI1DSvhYz45NT2dRrz+TXL9kPWPuESCUHLnzdpwSVQV6zZzAt2oy3GGaefy
0hB+szQ1q+wO5NinzeOPxJiQaBLB3f9XbaiQLVcw5GF0Vw7/SoY4i386hdjyvcsj57kiC26/VqvV
l0ykNm8r/swyS8SeSYztLv/8OuHyUzy9r1dPnORhMCKZW9+xhdu4D0ZHiJl64PI9rDehxrrfNrJi
qRnsypTkry1kaA8Wq4t8B0uNZRAA+rMy3DZZfdWOqnVQE3kh12tgmeaBTANEjkGIpyrX/UFGl+sH
RYixbD1oLx/9OFo8C01nZsHj7jp7aKpr9aA9CEOYDPU1TZ6aSVuEIxD7qfBDjfq06CpzBW5HAkyM
+EiQgAtJwpsgpLML25bkXJEHzOpf0faXBFtDlBbLw+yKGX5i1XDO3c1ClxTtAYcxyqYLaqF8gsPv
I17Ap43enOhUrTnnU4+VYOMfWkuVz4qPeOo1VRHSIGoqfpXBF8JVsmJTUPoPVDXORDcpA5xgJcJm
D4sN2ktuyICUHqIc9VRuvF4uTDTmMjicxAIDT7KnytUdBIkqBUhr9zW6D/1eOuu+7qk0APcmu750
/L7niY02Ga3Qm6PDNtWaNXkSu5lv8YcJy/VRQY7PqKZqShMr2JMTuotHgRwq/8EoHAPhd0LP0GdD
vhSYaLQPy8AG47Hwmo7FAgWcRnvah+ocAfBOaPTTDcs7wvx+9ajCoWYrlkew1a5pMdQJ0M2J+tYi
A5+DTHWV6aSJFhTCV/R+m6zdfuykDr3tm6Rs5UG/FvHY1E7fDmAAsRFlWORERBrM1VCSAZPEocnC
zrI8/Db0WNY4fk1IDJhW75wbGY+YKXkKQDHeiqJlpBKzwqvPjOUxrEiZ+dkdxzNiJXPNzw39Xh5m
maDjS17lbkmLXMAHcoj0WEO6QAajA1exFza9fAXesRkYbhEd8MJ50mA+jE7QZSKi3aofPFo+MiPr
TD/VvotTYiTfExLM/3YDLvc0v4kBYVWTC7Xg8UXWZjHbqZDQRoDqRlUjNxiSU/jzcvU/g0VWordN
25zR1DTShmNFNep4dHRdEDPi2xr12PzAVfxjywwkim7sTpwEfYTMDrgEcX9Ch8R9bx9xZg7WwHgv
ZAhQC6C9T/meCmX5wnNekxoyy8PM014wKuCsVIiAJHOdArDWWx9r4zPlLmT345/N7FXutKKN2ZxK
uf1iSvwRzSU7qscOcZWEMKZHyVtcG+QVomf4+5VF4ClDWGCtxHlnXFsfgOrTVIKRs2Fz0ExS6I3E
LqxQOlPIfR1QrxCrCTFVHQ/sw22VYbXwv4XQUR0cFcsiw+HRrsu223ZwT8HV0+9Mp98W9lsdBm05
i/13b5+cGw/kDwr0+EYAbpL67BA03zOCsfQCNDIyvLh4kpFnfh0PTTdEz36f7033zLgl3qyN+xBP
EaXzFJgmM2W4MKqmOyc+MOTmGRCA5lPxpbe0SRBy3LKBxAW2fMJvt+GNBPLbTPVztp7dXKBwPAuJ
0M0SO4pAJGk+rupVAm1swXqBYuSjCk6DL6Xk9wfRi3Di7bm2i7vkJeqDwCZu0sWhKkhoY73LDXqS
gEN8UB/Zpq/69yJfOtfh9jvON5kw9xf4ts2PXYHek8wHJ4efHRVtkKIB0Bmut3EOlaBFDa37yJjj
LxSdveoImj00SXyW1y5jsjSqV0/NSMdlkUOsV04Gs3kORcNEDjfJR77A+Ak/+hW7r5sr+lx+7KQD
a0vDQsIFH/PWUA2WufxvWiKX3Kz0r6llruZeZF2V0+O84RTcZTVW/sIQrPEnSRX2X2tznaHBgUbw
hbV5ocEtTjTfr9LXdWxzFFeTfKPmCMAUiTJjIafQSpzT6Y9HT1hhfUAYPqAXSy+FcpGXHwzQblEV
jPQi9efiMR1fycNvSCEvNDFnETt5A9cW9MbYfknv/7EkwubpAkHqX5f5mWqkkUt7Cx8ztp3TwLo0
Ah0x21PBHtfmbsE5WrgUf+Ea5Imx9AG0OSR/HzIxnl+qYKe5At83ZAm9Hp2c0nBgRQT4tn0Tt1n0
wRSemINkhaD8Ph5xqi3uF2aJ5pUrP7JdqbxgV0OAKcAkLfcvIJV8YHXVr3T0Yf7yL96zVoKpYHI+
jDJk30UP4VIV7aIHt50CIyvUH/YSHhmyY5QexV3Dtffm0+phxJT1LcIk28zMN+a+HUjyCwh16hpi
nUtxwkOBf9GAoR7LEI8VmhxRICimrJLGOy5RwCNFmpmIkaxq9nAGlyE6zHXBRLNsMXDLmfRXbQsg
R+x5OMnrKOVfVqWYBVEEZF89TCFoeMBzsUFqcmCT7U6wYPzumzxNWlpCby4GyNEfOaSgEEcwjS10
lR7UiXm4GM4EN2PA7904F/QEBjg5wjxVVImZnfokdSqgn0ul1IVr7/3TlERMwDUg/DtLJ9hItzzv
YkjJhr+aTru3BvupsIRTEB564PkY3FEcu9d1t3n/kk4r3VoN/3Y98LZA2hZkgW4VYmkV6K0vqcec
ZCybLrbxWxVqDv1Kr0Nv0Cmw5iVpZinUeGFufWOvD6R/AWAZ0ZVDBUp4na7cgkx5iFa4cJPt3QOC
G1mRAnBpmjJGLNWswRQWnsi4qjw1wpSNbs6241bu2+gY/ek6x8Drad6sPAKbNQjULcjtopPFyykm
4i7JfJ68HiidFKOFTn8cP0hBYLWNKNfj4bmreWjHg3Ft4lbQdQQucFxUUzarOOoBXIQax8b8s2xn
YAHaByH+BO88ALAzwCDxQU6xIzaXZibSa4eW0TtwdhjUEOtyCbaVVz+RrUHM7w0MFU1Fb8Qpdwif
GjZYlctpIeo+PT+sjxPNrd6S1wD8i/+YagnadHcAGT7GP7u8XZfR5z92zKaNeaJP51LjpW4D7R5E
8pgR3lFX2uQg4qghunbk0GZv1WBAivcAdQYGo3kiR8GRnowmhumuCKeu7i2+ocH41dmDh3N4EYdW
sjYLqXpwWqOuAEum7o/PSPaefq6TOIw8S8rTvgcp3WWAo2yCQ/4aPjcZaPLIFVUzFTizXthA2kJi
ymxAsIj5qos/lseGMx3V4bynjusV1jnyE8WUU2VqECDPJhNoSbHEMcyj1gs10dCgMfyYN8axflgL
tSjxxG3x9kI0MPaiQbNBJ1b7eg4wMpmdRFtrEyoew5j+xxk6GIrwVR8DUTXSJCV2rly6E6rSpzrL
4hDXes0NsODU3I7E2q1JQNKI4z2LuqRnuxXqt02KtZxH6Lf4vqCfiyMJyfqS8dlkv7s9zQjnBG1F
XRk5bDAzCFN4S6PM9LN48OlIG/uaU7lDntULFkJwO6+g+nykwUNM2kPb4f/b7oOkxDOsE2TtwsqD
mW7fJBWHXrlFvoAe9FGV+IIBltyxMBA0zutOxtx3r909rmhPTvfWUqTBBwS9h7HLwj5Fp1k3JTzD
zDg3X7e3FdAckU5VHDQWUUiCYucH9Bv5trdgYxxr3fwELC07xT9/6k32oEGFP5xTQrMVjJW+4HxL
Mcbt//kOZpwoT5E5vLfciwxDKyDr1paFoBgE/PRYrPyzlnR8X+KFYOfLqhHfTTwe6R9C+4VbCI0a
xuYETLj7ZFKJ9h4hx7GYHCQi79sclrovFbh7f/SOB3DvnyLKztSTF1mhyjHhFoH9djhZwVHLcpsM
TG2ufsjj9p4Pw6t1hMKxd1C+cmNbziEuqTbTUBa3IfF0JTgudid32qvueqHSc0TRzTsXlHovbGlv
KlJVa7efWMPS8Aiczgpti3OKYnEENQcfABx4A+/xIZG5AYyoqnqgDAiZRGm9qghclfnsV36JPi21
VAIr8w9FKIGlKsQubUjZTKkSQtlPpqVbjMXBEwXwerWbnNukw/yhZ7lzycojBSJDTMIQZy4JdG4S
AqhOfu9crK3eqhijZ9Ehj7a0K8hrsZ5mfluukVOfptYcKAQZrbozO02lue1CNabz6VXPZSjXmUOB
fSe5aMcNTLqhTnThplPLrnAOc/DlihVotu6XtyVhr6OqoC22ELsJyo9z2gpkgcGi5At1GK4wMDie
B10/C1LSlmnaeT0TWZNBjvJ3n7CQVkIwbUQvfh8X2q/+VWycDbGi7UFVqVMJhON5v4kFB9eiz4pC
AsfuzfpZPHU/LkOJT/mimnO62MLhvb6tbp8pefzVL8mQxUPs9LhqhHHvFCHox6s41L8GPfDR//ko
RMZQhwA/EIDm4Pzt0Rp+8lv0KSUKNIuAEQ98YvtP9TkIKfwL6qUPVTmqnzzQpYiTlItk/RSgOCLY
SIdq9rWfUl3GhIl6wuwxiOXfKAVXfeQJerw77GyUFKSzw0K+CuwRBx20nt4+O8rc9Iuvtw18gz5e
DYCde9nnNS8tcmOV2c0iO5OLpngFZapJUxOvPeHIHe+FGZKMCs/I8AesEiQuUgc1l3uztINtPZn+
8q93n/rl6ARMQbyRxhtbq0huaXVcZC2/IBoq7pcWlK83wmE26w/RMIzxhGkreXmZl3xgnGai5vPR
f1H9aAPRfk7DsZCXWS/wn1jBE9qJAnAT0C5a4UhsVZmB5pJGUt2Ws3AQhoPzxqNZJLZteq9giJPf
VFstAncksGtj/Tz9CuLpI2hKZaOSQQeYbuHC/yGyjTLcOtuf55qk17CbRa9oClSzgFJeo2geiB7i
jDzhCAuXzvHFzyR2Dg7PM+DkVzkIbn0YmgreARHI3yZYXaj5NLU2y0rPlqALV9c/o1pcf34RYMH8
wh+J4G3KHwlEKQwRriDnkL/YYDu3RFuGUm2CG2S/7gtaAxX4DArrMPVVGNcZmrF1AiEGtDg2eptT
op/801DH7vGzh+ozlEw1NUMTgnTFiiHxqh1/R6sLL2u7P1B16KhoRe7ZBOWqgr32oj8LcM/6cJSK
kdV9zemu9MEVrEINWzOYVd/WNY3YfL4/jrfdxY+yirp1zSKNsbqwNCjkeWc4ly/Vm0dUl6SVI6rF
K7+Q9ODY/mJQAr2iWS0++7kbpqjIQL6q2Jx10B5/PKRfPwIe5CrmJjfXmZeFShDmkpWU/qTXGg0E
+W7kjXV4HwgD3ltS5eAMi6BLuBskKWnfD2MCdfcg+TnkR/NRhKDQOHFmx1KZHqLdM5Pv7i2tmFgb
EuzLadMui1wtPXaxl/OKmGyRpADzfwLPHFiBPFSuU3ZppTO2VaPLfvPezPSNqV+cd7vZFuHshfhy
T9YupmOTWNGo8rQE3wYz1AvC4MbjjJ9ZOedvA4hp9wUhR+FWuPhuALjOnw5UH44PD2fqciH0Pih4
xEOeZYyuWH3Jbr/QjmfvUj5l/rZrWR8xeHa0Uzl7FcWQEBIXfHJMFVedYp6SKdlLsUlhA4aaSOGk
A0LEWQUlUQRvSE4Tvsx6gzOWo3gS9ktjL8iJzP4aLGcYbWEfacPFGg24vaT42I9gZqj6yWoKCOVA
DpaxNZTzMbNTket3nVUHEE3Pef/hb/D642AmwZtvhYCCnZi1gGQqzHnqqXvmqTgnoFTLrrREBx4e
bvdSGBGWVERrV/wPeNcWJFkPT6K7sohJtGbsLkbrh5loEjIo6HeOI8MuFXbV42Ium2XYARaZqg4R
8vzIx+TpHAH8T8ctBJq+xSKuTmmaUAO3tsotIPC08jUXcIpmvCIawzTdsL4+ByIFqPpissWmvve7
QD7S+emnof3vQFL0jXHyoNL0Krq34+u+s+i2ef+Dwo7rWLyRxPZ9bsv9VsfCdqZIin3A5a/iit5b
OoFMvL6yGeSSnYDqc23SdXj1eWRY7/y4vrv0OtyxHuimr9lrNn3Gnd2iCvvHLD9skSmA10KL6REx
Ry+5Nq/RSkbuhLijhkw2fnmriB3ZoFIwH+VnNQMXgZWG55S7MgI9L2wBwvi98MoFPVjFY2X1n1Ux
V0e38P5domZ1KfvEvWzE7bmOe2rgp07wP+AuViBF8oGftpnGefGKAU0ByFsTAzvUFUVUpgwSkEKa
sBKpm8b/CjbIRpHmL0IKccKo+n6WHxfDgmnEsZ4xV5c58T+4uqMgIUPEogUq7ukNAQvb0Kiw1wd+
w//wHG/Wo6KJXvAb+cw8qz+uxrN7RGB7CfqaA269kWczKSGITgf3o2bsdNXWG4tRjPDV77YASbN+
uAD+2soWWXHc8g9ioKG5yIAHbmpAovTa9dh4Gy9KN8+9stO2fb2cunq5F2YyTuCKTh3x58/4Afyv
HHseH9f+Oeuo6SljRT29XFW1vTHoNCCsckoYJGzSQYyCbvNHl1i5MdlcWnjbBSO+yrSui8Pk6yiD
OCvuTaZZJaWslfbiYBQh43hWT+3Vk1uBGmGedvjabx5y7XQ0En4yLa55FWAx1wkhfLETFCMsQqoL
cAkzwPw2MiMDxnj8XEZBuxH25g4wGi9Gjdk0x4rMPdEYn0dX7TIcU5xKARd9MLKFNZfYjVr8D+91
gMWOzWIoW4xw8PoLLeBm0NP8YV/IFww6RM+RYyH/376ACk0DIaiYGHAf2tjIsASl3ROURwC8MwHL
2KjKQyLoraMcTELpL+7dfZtJ0kdx/ylfUyxHUytY41oIWBbrm7lrVPbBcEc6M7uSqNdO4cbuhk6I
66nwlMV4Q+5yeAtr0vZlw6NKk40rZ6YXms7dxhlnxNQqRwwfIdqDHwtveS7xg2BOkWEYvrZMt3XU
GivqlVvGgs5WLY4UInofmmy1vHUUWa9FCK1SPHjO2Gjh5oQOG5X+6ZLwNqD/rLXWf4TMkN461fDr
hJuYKxA0ZpU6lY8LjqwS9terGJCjz9kzRbzuLPzBCdabeLQbdupYEqG+OHmBV350sG0TVYGgK8Il
mgTxumETHhTBH5m9ZHUNlGdbhYtVmOYwlP3SL/soUQsFQfk4mqzocQmTgtcPF9W7Az1yWqxLpXp/
pbaQ86EE8Tdl9DCO/4FcAVrxzB+tZ9kPOSI6IPsf18Zv6Fvh0FS2xoWThVot1TAf05fARDfDw9eF
bGUsx1tmW4wmCqIF8/LfFjE4g7t/TyFHAownflf9To9RiOF/PIEhqnDs0ynKPiWUWNYnHo5YHxUO
zof/OOZjF56gm32xjVzslm1jAILW9cOI2Hq6rHrvEuuzJYCaCywj7D3yk7wmuBKhloHuYHcmzA5T
jslSu85F0ohufz6IPXa4+i9J4xuu6/AVOhVQCkyTW5Mn7/CiGc7PnjhYDabiDm/xurpiUyOG7onV
qN8B/5pt+rbhHz7h88jf0Orwdj2DboVAymTWI2XtXWj3wCrh9koEuhB+RpXy3185RnFvFQcxl/7v
GFnBu1GUzt4Yfn0fbpESmB7oOg5pQRe6Z3JWEPjv2CBI/tqkRxuy9bEABxJ52YSW3gQ0dgT3rPbk
OrmUCZLjgU/AseleWMIR59ShfnNelEqeCbd1JTtv6oSpX1psWvzNzq91C5TUXlZhXLcEJHmUDghZ
lvhFVlVDHKPdMdaOkr4JRu0G3Q9p+XWbRRBbeC2hXMJm6CCtM2HsrODsaA/EFxggmw7/P4r3jZ/l
2M45Vo+tYYO/iyJWBHijGN78qpOV6C1IAF/ppgh2yABE+jrg3us2J2xsPOjxlALP/MjWUTCSTA5Y
lh0k1z5fbSr3RC9sPgrtJaQQUeopecGDsteypMPSvb2qS13Swar51WZHZMFEt1lj6FJaUL1Pr1xe
UDxyA5Q0WUAMZvz26UGQe7mnH/tS9WjUtZjRM7lb6GT8pjSI/PH/jt71kNj3IQTaEnr3wQGMNZza
Sfoxlgt+leUsGP+B1S19Ggq1eGoI7dJIbHp8FNzLrX6ATxbYkWzn/pFH8RLz1g4oQEIkTnPKDb4L
PvN7nW/9hWK9gjQY+4PgACXnrQCZn4RO8ss8bZL6QL2FqP6ExOgmqjtDZ7FJZK5JpRQy/bG3mMZ1
Nyg/wocixsCOZWELnh1JztV+O1QFSJp9Jb4+1TS9AgurGPOzug7PwzxkNFSUIs8yS8cowh35O56D
YSpJ3iLjkSCnWbXYQj6qyLmYxKuV2xdaSzvmB7n4PHo66H2HoiM5/pO1WN6uW8e9w1t2jTb7xvcB
KAo4D0fNro4hZvR9bid17l6mhta0ZZZMyAmnOXeGsDdpOmwACt0r0YQk6vPlXlILYj73seDDFrpG
ETtUsO90Awu7Dg2azH3tEWA28uHdPA/Ix3irQvTqiH/CN80++aqs+JNifopjJTQZrvW2IRmmkJ0s
PVkEIAjAM2rhpTklbOyS3FIFBGRXuK2y1ATOJcviM7r9saHGz6LXY7wA0SMApJnDIhbx6Du1k3gl
Zl4P5ZrcpPFF2G9iLRRmU/KFddGZX1BvPA9FchMx+rnaa2rkyWdTNn9mOdRe9uSWx98w6BeBtdMa
nFVWQ9/HmW16/zY0QHFH1VIbnh45LT+0OD3DK4gnVe2r5J642aAX7gOiRmFwU3nWE3Po8Jnp5P/X
9jcXLN81Dn+KB5ERvOKTnznaCDmytuAaX2iXpEgkAzA9istvRQMs3bx1JM4FT91RbraJ2KnTfBuW
YTB2WEUjhHIxxMaYhtP+TeqE8/PooR+yy/G7emXiDlRURIxn8zZ203I57rsTgP0TvRYwOVUfhAGw
SQ7tqMhDOHL6CL5DGlmRbkAE5v46phzAzXeBwXsZPFMuLjndbfqu3HS6U+aAJ5FjI68h/ib5x2Di
rgD2/Zzilu00oSfqQ1cn/13tiNMWhTmB8EVjjxZYSgg2v8okT7i+HEneYwGbVsP/Z0YrGCjXR3nJ
QDxwFnRCsPiXuLkeqHvf7ASZ59f0uTQXpa+x9QQSX3Kczqg8v/J4TT2d/38x9ab79lChGU84a4WI
VzbwlZP8b22MOq6B9TW/PkqycyPP37T7ZwGy2BYIfbPED5EuqEweoQuyMh/+uS5tH2Di66qgJCQU
QS9/D88S/6EHcNCej/X9rj6qLuH/BJS9qKZ6nZ6HY5q6NJpJDGotP0D20IfSHYZ8eEuexTdlkIoZ
Id03UeO6hn1LukEx3XKpNSdIow89RoGh93IoY+kAAd0W0teXOw0xbFCSeAlZ7TuiTHYu3eDnzwEu
LR9SPCd670p46vLoxc878hGGG0CZUltli5yZGCLUC4o57hKEs44kjEUIxXSxffY4M5hfJqZsOfXF
CbOGfUtBjsXVzy4H2v7XAp1Evb3nahRc1W3Wd7U+aPXmiiL2yXcybBCR5B7ofaqNT1+ZXYwwvAek
LrK9soVRA4VFx0XDRhwtBafyvGL8hNCxy5XUbkr5raOKRfviun4ticLKA5flLSx0IQz2ZHjf/h14
O71EUOQb2OPMBbujyyNNCWyg7Y0kSmb4bqpS7pWsOpt7tfgA+XYGi376m+tHOp88qOIRpYSMsUhh
c3mufRfvU1CrcntO7VXXm5mXVvQT72/vCHG3UMIIw1LdKZS7jiLaEteO90qrkrDNCriFWE0kxciK
eQCb/GuOhir7Ecf+dGA9S2ESZ19ivsFBp5iaRHyvJKyfGOJMGFvKUv5MrAUi1eh0vtXoFFFbiyDi
z1/3W4UczcXDBPKpCrJpHUa8ct+qJQD1m0P3+xYs9DnuUxZB8OiDOnJyRbmB483J3L9D/VuvHdjW
VGHzgA4ihE0hPwrq1io+a6QhSypGFaRC+3lIqbch7/fU1+uVxCK1IWWqDPDD5sy+OhYml0ZFuryh
JMrVHUle3Rkf3cRBPk2qPvxvWWu2XIjD1gM+HYhvZVkpgID7X7TTpbBhBZzzBM6H65TVIy1MFoSs
YPggKkHdjry6ZhnMATHYIrrcX6qD/OfQ3ZcGiEMCiTBQmZcHe/8mfp6jMM10MIFyW5JnqtJaRS82
jJGIwu3ML3yuXZNtybD5gFiWklxDgc3LZEFd6H0aZHGKQ0GMyhFbhOIp+PDqfcz0HnpzEiJzA8km
f9F26imK7s3VsQDDWBvNckJqlM9Wvtzn5K71O6mU87HZm9pskgxekEOHOcGUmVSoJc8nVJrfwR65
QQGy2MZao94FnDqawNn4L3pI6PfOemq4E25AUwQn9u8IjiDP3dDcRKnTOp4rmgHm3TDGhuK6ot63
OBdqws5bIpe89dwIQRvBpQCsKMQNzOTAEIPSt2TjvafyIunIovyjLGqLZwZz5dlN4PUYskZDQN76
5/4CULEIMf/+/JqnHgz/nql/klGiYA55TE/2QhX+NsDPe01ttHmqgBe6CSxfI1C8ZcCPUYa6TBgY
3UdaO//7A5JnbFne3KJFGCcWwzJeoD15aievmMzVObXOdiJ6u9hPHXaLRTfIJsJYkYFjuTJV7g2L
0vrk9azlJNmgHVjPH64Yc7ROezkhGu2o5WyCAs7LELGxOHA1w+ZEzV1ow8NnSmsZ8nMCIHXz38dU
UuirLciAy5n/uoSww7ovRt2+qkEC0fARHXZ3y1BjzbYzOeeyo+DHNHyJ/2JMv1QBJ0/M7emZzryl
sXR9A2xR6H/xN60BrYjFwi4Do+SKYC1I0jPb2VkxFjeYtfnp0g3HvDVMxetDAL+MmkdHEKSaR0BE
wnpERgB+ZWylNEES1NCLVmTFPjKiE04z1q6UFezWi0UVNs4RfXxExK9vvss86umi+0xfvj+WJUu9
1v2wS6vFnbiy+dO1Z1eObfno9Q1zPzclpK9z5Kx0ewQ4cftbMauRJ0XPTNuodL2mNwkSG2nuNGC1
bHMy85MEjf+nKCjOtCDIqxuHE62QNs8evHDXOlOCmW8ePTtTfmeMkQkI8JAIrhWqsf/ly7D6D82I
ooYMeiw/pf15fY9T61cyeWMMVRXbUCqK0jerjKNkDm4AgIn8Z4qb2u/3I3nrgo2aDSR2CHAGhXkZ
cjNvtow3rZTezjuG/ORE3X8iQomZvGlbwiKTpZyrr+Vgc+pO6Z1H53+82I8jPOqkMeZe8TOXM57/
mgkPBdZlCVSpEanUxdjheDPD5LPi9NkBW9rSS7EJYr3dvOmOCLu6Gcky7y+Ng+jC36MUgQsuDkMI
Fp9BZMlZZmUxnVXi+Xo7ATYoRLe4yMKtP6IZlvgK+LNjlTLaGA5aP/9MwNMVksI0SpY9WPo8rtgw
Y0d41YZ5qYw5m8NnkZzqI8ZLSexmI2xyouegKiwMkvpwC3PLN0IA6DvmjPHx5tr37Q73QE+bveSw
7FtVvgRzH5R6QSC4H6iWtEaoNuzVgkSVKO4L7+iCIAUWljRjnU4QERrkz8bNyV8NnHmkc6zPsyY8
AKbPDVhbBKcppIWAPDm2Jui6baNKKxpTLmGpuNepXBVKydb5xHXvxGHWJQbrrozC6Vqd6l9kZtXp
TNkIG8Je+Z1VIVkpc4Wj4voorKqmkpJZBGqY+5fKunONV6tCXIfWWkikMYqnvQxKIBteadvIlQFT
3btdZpUOCr3bWBUVYpKOrk/rrirxVPpN3nVqI3d0eibnHpTcNrRtZNgzBRegOMOEZ+xxLtEknCEa
c6NLBvix/oeakDmcP9Fxn8BqasDSWp0KmKDRAX0RaKJhDu4PoN5dzXEgJj/dQ73/EBAJjr1G2/6C
3pEe//IILly4/oQOHt3WZw2l2HNE/UwLAoRqa1HhLupOPopoHc4ko+sTfClyTlBtd8EdmlonwELg
ChXJEbqxkYbLV/fprXPxZc9tpi596s9yTUt+FreYBSemTt92fzuL6AHwQ4jNGyQq5ekeIGdjD4Fj
fNqgkv1YW0Co2Ygf7s3LP9IsS4oIFShc1xaVdruUimbPzDUUAGt/qZJXwNa5wsVb0wOMovh+8xhZ
XCBW0X+Sreqp9nDH+LRR8wVRXTlEHoovIjw+FJUQAWRsRHMVcbLnRFSo4mZoOLgok4tVn4dNWWhY
ATBF5NSaD7zCDDy8eNs6bg+FaOjWhZMHdt2y2LM0VF7HAePM0nRQz2HVjRgALikKFJRUpoIQU7UQ
xkCW5I7MKnyX9CvD1GORGsqkgxoZ/aDuLEKNQSeki0oxMBiqWXvRkZZbo99RU606DqWkZh3c7vwX
EjxPQP58QL5NMM5bs22p1l93u8JcdEBhvWQiYZqPcYomlragRfnKfRDS6Ph5iFx1n3ztQFkazKt1
1sb8tSMVla4Dkr1HgVITQ+9IradWUZhvPfA1p0sA2NrWwbf3YDNbD4PoebolyaazTiY78TjPWT31
1/cgMKQ3QjQuEDubL9RGdsvfV+SACh1AB0Ud3FSlGfTwk9Ue/3jMKwDWrl0yfUT5QxPfX2PSkjhb
iVWOfUIOvG+Cm/UUtP+xT58u87jk8ywEYKSD4bio4+C0epczIK8VZ1uTp8QI0k1ppdZ2NEQMwy+W
7CetNeruII/C8Rji4C5Y7f10DCdKj1NRmOYDz67+l9UVOYG0uPP6g7p9Eb71eKiP/mxOWFEVLFvQ
LZ7AfG3h0c1zm8Zw7XMEkHNX5ns+7jiOFXfr8+nPWqYn/z8igh8frMrmY+i3RtCjPS8Ocdiel/Vm
uNct9ppKmJkQiQKIr+9SepTryDmAgWXVyLKjyTLvA6kmkb778nGyurzueoAykzszuqC4qo8lf0/Q
ts0U1BBbURfqwxr09AHamDkDUKuiIanRYKKg/7xCY+m8CTsy+dq6Ri/J8We9UfDn0/2/4cbWbL69
3e1KsoeDkJE4X4y+Cxxr4pcQ2UqeOJtcAYPMm14yuuYhqRe9l/3/qpzH/OjRZixwclgnQ+z4A5K+
MmcnU6YEewSMsrdGEfayU3rVSbWmC46UBFhVSZOc0IDsG/OTCsESnzE6rQHoAI/4CqiK4U4PA8UI
hJQv1HDv3l2P5/MPhgajZdmD6OoAHBpccUL0z0tnhe7hI2okrEA6iZYV3+99FR3x6hUmQFEW8Xr8
W+Bg3E0A0TLgKaCXALHWpmQH2RZRnAqVaqSAZGzbqDe1f13dXD966F0agqEIG237P7yRRUjdbIYu
DTmMI8dqbuZa+kvCKkgoHU9zch0kZLyBnmAzKCd+WvxYQ3Rw6dIm30OYfjY627w1+H//gEXqAnPX
WO00+Cn698MazV/ZiAxgFTWU7lpspENSkwxhSlC5KjhGBTzw8EYxqtgA4QOikkCGULx68H46BD/j
qm05ktDzSaNv+ajNedOhfk9DLfd8HfcxHZzmFVMOQoATG4IAz+9XP8KI5cvmOPNYzRYtqhyBsYZz
g226HMRk7h2yopCnHmY5lpVpeG7VRG8/77pKxtnDHX2ysjxds2PK+Z4Gwr2HDXDsE+17gTj4PVZ9
DTOuUB8lcavn5zAZQATBlkZWkaYOoP36lBMSOYiACJf4Sc+ajcXLqS6uAJLD+EdNrnhdRbzon1Wq
JkjvaDCXoSuSl3ZecQfKdLRYHcYE604JbMoo9STqpdM3hEanSeL/kL9KNTpXdqJrffRpzlzia5AM
tDL0B30NuI7ocEuVRg4bO/qLENqsIRzPo3SImK+CN7MSncKVoMzm+itnNi7BymzM4OE30ArMY5KL
+T131qoIwDeflW7fEGgRR4tR+aRSTObgRPcNn2/72KdFj6hKeThJKvA8jRf9ek2v0tfjp5mHhA7C
ekvyPVWlU6eTiNlmnZL0vD5oDAu5ocGHG0LoPK/6zERV/pWFtKW/AtpPwOXzg73jzNdVl795dWkM
TVTZjugivyJfifto02v/fJKDAL0LCoDBhUw+Hqhdbvc/TLZHyRe/axColAFS9U+B5/Vapu+u6dL7
T96He1o++NdNZQBTBI4PbkR82/amgYCihPatU9bImu/ld2BKfaH1nUOaEDJw1bdQzRxiYceEZtwl
1TKwir+FG3rHIMAUTglWzua788FBz5ch9rf+pBc/jjNzj/Vf1Gs11pUBN66naUn2buBzHQb2/i8y
PLwsToX1UftRsFfR1EShP1mbz/GTnVrPpH+CKvPVeODjciOLOF/DUf/qjHscPtFspFHmiDwss2qu
WGWH/pYve6KQc2fQFZC2iLU/SS1j+aMWiNfQGtG+KSsBbcUKHhodTl+YAP+6xLTmA7hKAXY46GFR
uuWU1rtbzD7xbmToP2LeGXff9tV9e0WBWXW2XRk4cTpFPfPQFtx2/LfcWUOX8iVlD9UvOKxyo8qo
Drb+Tj2SxTNmUOmQ/WqubPWMin9wot1fp3E3Qs8G3f67sEx68kZoL+2pmjN/NBzM9LYyMditHz5x
s3Je/nLYcmZkGH43V276+D+TxxizwmC272jCDPj8X5MH7GA3cVLkuBnR4vOCtqNP/QOUhTsxo4um
psaMFRj52lJONYdCNv3WMQWS8ICE0s42GUEbHmjHgfXbBoeu+ITec86dCE5iYR0CFj9hGb3dlU/o
XfPxyEp036+Fn17btVQiyOBfWTCaARVbRPK2NOCL7F1mMfD2g/ur4Hgb5nwT/ISfyMsXPp8FhkJ5
UMByt+Blwqwu8Dxrmog9jWFZ58W7hGkH1WHtsjbUlsY5rvTNFq6iLDVO/izl6rS043jE3vx6Fny2
xY/DIy35m51ysqJkX6RqdZWyvEyYoY+6vPh4L6Mzgsj2OHeeLuaBgTQsTX7YG7xyqLHcJW4Ib11p
wb++Ixigr65bwMlGjBUCW8jttcOBNaPk8vqmZ8J7Ov7UhqpIx6UBD3ncerrIM2/KhgPb800uOBZx
bHNxj+i2k96tCwxyEWMjQuJtSBdBGBdBsB3ueFvPakU7eUloHEn83d54Mj/u7NfPLth1JOvb/czm
sru5SLg1n/kcAz5SrBQFOoVTAxkd2PiBLi0im2H4faGZmbUgpfXe/89zilJq8R8wX/F/+QxHsXxn
vyq+gpEffw70NAf3LlH0pWrsj2t5g7cmBNGGey2PIZutyvavJpZfzMvAUEGMe70zO+3rGy3g+Yaw
s7CJxhyAwLJ+iHzGR6vsKcm6AUJTQ0joo7NnETHnaFA4Z4ZYHMIiXo54Qw4h+f/GFEeeA2PVpQCE
3cpm8jyv4gHzBIzmvcWG5UBNpuam5qyyWme0bDd93emtUYYPvieXnz+0HN88mOthVyCYy6glC46q
PEkjzo0gM77CYf1jawhPwuAvKr2o8rSIsSSGCW8y0wduK4rctTqu3KEm3uUp+ep4I+gHnNAmClw1
iCp0k2FRXF+nJFck+BEuId383rqfdcHJRU/FdENDE34rbyLNWUD6Sxh0hzdx0asFe6NNSipUhNdI
BvNdK+WEFcYOXmzOpGSqsLZrudI3LuPOnjGfD9UotOXfBkzxzrR52/eP4vSjM13mhKjEUXg+hA+K
V6uYYJk7UAHSOYmxSw1CaniM6qU1hXek5LlDinY7iVuzv0kv//NrnMq23j+LnCy+uNovMQZgWZAa
gVCuG7B8/HZATfHQ9IEU1AOgROMfHjbDBoW4RvJ/X23bgTZOLAykDcnl4R8uqhJUyfC/wRiwbYb+
XyW0LAw/rXGbTB71+HBskwbobujV39AOD+c2qTCy5biVyUjgxOfRUkM8gDYOTWXzSJe+efeesP5A
j8zzu7mgFkcuwAylW370Rfa+1gtBUTyJaaSGj79lQNdRejqKz4ns4bPvnOqKbIzoQ32IfI3Bg2F1
ufR56uIpn+JrvqE1BSH6lm/2DWkFh6/xIW7nfLxjQfaKMjXiJWLC8HtVgL13hd3ZM0MHXpOy2vbL
Gx0On/DNRcXOrqzNISUly3jJvdN4uo9Qpl0XBfimaNm2kpmpi+8EYiN5WwxJ+5inP0yypdgsvoEZ
0Odzwsuhu2Pu1U0WrGtusvRQCTEDHnRzw9F6T/pPMyKt0/UOvyoicLyAHKIiYXuu8LCnfCCfo23c
LX73KKm6ywA+MI9ZGYRebLxxvVcbG8s74M1U9XJFGnaUEpmMuw8lZkZ/RN48Y4pLnQtN2rRY/41M
n7jnnJzW2tbWcYufpL7JKDHnQhxtTtOtrvZsn6Z9NQ4h3W5iIetWajNg445fTeQrzD0+QHIqNF82
E421/XfLUZUgZhaOe2hwrB1yijkVZm6v7QYAAihqihnyJx2r9fRKEPTOvMlrFNh7VyGRSBWORKxM
M5c6RFC4s5441lWTxNDqIpggfTAeadXsps116tzJpKwf/PhKdemZAOdgcF/l9hceqsiIHdxHZf/U
Tl8HrqaXZbFJcwJp1Abz/U2oEMNRiVveWAad+umeyvNmvNSluqn6ulYf7TKn8MR0MeGUr2jfpZib
4oLD0/W6FKunZ1qBaD4sXqun/Ady6KOquAEZ4uZ2i3/wiPbUfd4PfSeAqnjQW32uH75LXb092HgY
Nm/Ws9dB6JLaP28zkbnua4UK621iyLpOMUOqCGYDqxmW+f8WCXBhg2IvfZUd0vVPtyXOox5uuAUt
cYCaUsKwHKWY+bKPWBjaf9kieuVocQq4e4SiLvus8lRggEuP6mr2LCfJJbeMw307l4wCsc/SiXqG
HsfDAniFaHvMuUEvwqeNP68wklsgnausZx1V1b8VrOI5Y/G+SJQ6bADmcmfmRY/DKtkrR5ly/EDL
K+Df+dl6np4syUBhU4pNmKVKzi3BISW5JGyfIzxQ5uo+X/1MB0GlqXfRZyTBedp1FTV+RAS6+jtt
SmwIwmUUWPQGk8DjTBAyNzFH3zDWkwziYfdn0SRxi4N5DgsR2SssknmGT1ye5GmBuZxGfKYlkZqn
h7Rl+aU297HJEArNADjPlRJ8+op+64l6YZ8FktvQuly3juZ6MdE2YM4JkB/eYDM0Yp/iZZ3mUW9+
4Ytq+owfuZY1VQs2RiA+dHSVhr+gdwBNINr7RdVIvc7js+cK3nmpwaAqU/HpqKSDg38owK0bdYIe
mRU+SHeWFOXWImTfHcK8GqvRrnqaPZK19aMoOTIXHLNC/jBSdced+WVo1+QoFqJrbSIah2FMTquH
GMe4eT70FjnjXu90pOZVoxISXGP98/+DWNBIrtycWup/Q8jU306qqhyovhBMcDpirqGlhHlK52lM
fdyhFb3o6iIbYzAa/nKgxEUShHp26XP8186elnaFGOamnzAPOxhtbzqCgM7temuLQx2uxbtzCdcQ
vlGCnqD+CYR6sHaybr7BOk0Ci7wHq3eWmiaYtkuyhhDwnmiM0s6bfJ0Q0TuzGFTdeJXq16WACxH4
LJmflLxP9yOOm9nmnFFr5DtnyQ2HVLTuDTFV8JYzygnXaNyhUu3lXEYbfRuBbPQKwoqrCPDoJSD0
i3Nghq2UP02DJTrOPaG6V20d8PpS7Fl7Mc3LqdepbfMgDMPF5iiVSYCQizk2mqPW/+fsEpnTyBsG
lfwi/0Gc04Owlk9jLTQge1QlEB3A0Tkk4ZmQqf0k0A3RUA9tXog6lcaiqEh3gu2h5HbNpALNGdA7
S20gkLxSLbB6CVEjrU0jI7bOI7XXcx/GaXWYMkaYfhWqMaj8yKMyPhkngZGgwG967F7En3J+7ajS
aWxuc+BOtRHq6ORTSV2e2DE4AD1j0A0EvKJkyjOc6o+6u7xuXQuKnmlz7oOW0zp1Sl48KQI43P2z
y+StWvz/TxFZiBfibxF4ggRaAL+OD8FKz3ffQ5Ayonl9I9pcJvtedJzmnau+luihyzpu05MV71xe
uAOHdzFe935uBozY5hRyuk/DRGdYGNQQ96tA0J9V5BJw5RYRYNQQUKqPiTRvK36AKf6593NuRwHB
SNiDy/nUczOJA/7gf2e5/dp9kPBMFHQExTWOw9tpqNit4ef6afPmEzTw6Asw6ggE8He2GNU2yl0R
XjfDOnKXnKxlznBed4NBCx0lxyAFTucThnO1h1pW8wFN9WL3hgN6QRImlGT4bLj2FtrptBUT68MA
I+Pmf0VmFHDSKlIZUDc111UNpTq729dyp16/H0pmYdFIXw7/vVADNuAdKcyqKMQuhcra6PgPoNwp
nG7H3QGPs0M/J2L60PNXMho5xavmdoEKhpnySdvsGgOfdUdKxqGqAwlg/5uBabzAMQzYHC+aMmeT
e/yNJCUR4NswcuMN60fHXvYFxdPjQ9T8fq/dqs5Sk9H7LzyCp5RvcFTZgIzrQTatGrwnb6DHFpZG
YTcCqXAm3QIBvt86ENMdJHM0IzRPidtAfv15gWF8xVY6nki6Tazqi8mfz3m8uWvt+VgYAegiKMOK
e7WYDeJuwpTgiYxFr/cX5hBKV/vsKetxUfPGez41isnonDGupHrDpEUd/6xlv2IKiVdVNFzE2Mof
CAOD2U0u3w4FkWXcCt5zmZ6G7EpRAnHR9KTRSY4tnqiUzNYBa+C9qPh3+I8foWTSjIRh0kc5djK/
8W2JC2Z24/3Kw2o/m1uvf3McSU1zm3H0pGCKC8kHYr2vNKgXe2SGeMe3tHvr89akYxC1CjYKkT+j
KQ93O8r7czctR7EngLO1uJCCSfvuEgb+qMA6C3cZX4OUUu5AVL7W6ucrtREXI2J8kvF6ZlTADCSW
52hPfLu0O696A3oSdNlH7u4TOCulwKg9NAsq3RSoieqGW04buSx+jlgz5Guep59NrKfIYslPFqUz
YfbV64AtZzBG8gljAoPQFiejwgTFI1+AUrT4yULGGcWxdUbcpn8wPz07l/NBYKXPJVwM8Ldn8V9c
ElPi5NM2buM2zuNlJw1Lrk8yqyalnIF6gTJJ3Fcbw4aQgDTHyOGqdc+lckxKzsUTSLR027mMrq4D
BlxTVmW2IeDkl0iwXOPXtYv+u+kF24xxU9zJ4WXoN+aMWoVTwjv4nFhljyeG/Jaj881WvVmcwYDK
Ol/7bKrCQOAxMaNKHMnHrHJf6xPY+oz8cHwssICcd2F6DsTQ4DgqtySH8Aikq++d+meTHeyywhLk
3CZFCrQdCkVmjg9EMhe8K/QJU8G9/5/J+VZ5JYvzxDNn4dxs9Ce3C2+wLrk9wtpcB+RbdIzdpFc5
bCZeJeng8UFOFLUllqK/VzoDSWB5SRacHT+N4pn7dRcwvkRd9ThckW7qediX3ygS8LKRRvjdoidP
FUW/lubzU1ggux2vccAiwf+xKGqkmlQLLnN3fuC6Lcl7GEcFUTUb2Ru2vmlHnrK1o4nn+sx1RzbR
BnXLIwUMIYq2lSICYXtIHlvRgTOVrhiC4dk/6fOFLnqcF/fVGzpksnRS+uMNKx6jJwH2x9sLMIH7
qF0N1bI2/d/tBpLA4httNv2Ymexm76/h96IHHpC+FOQREg+ZUFPN30Wx/cnQef5SXnhaMDGvjemi
QFNJnnVlfDofy7E6QPVIjxeBb6pioG4Z8a7WdQ+mHjmeemSR9cgLkIQCqf3FBiN3KxaUWj3RWTJY
Yt1wilrYAMbmLir9OnucqWBDSHOH5E/UKbowE6e/iGGjz2EfWZ9WVCo03WbtBJMTfYEroAUyFXF6
XnemBAuHQL2UBJ4Ll+42sHMb2QSVS52sg5pXr/saw2y5lIw9Rwtqgea964py/JnzHU5c+Kuh8ejy
zEH8yR2S0iuRFcJ9PSXhPtkuRx+wrRIemAruQ328HY1r6nXXG0R7prVbv8Ye72bMtC8d78PIKIJA
qJMUKcEyC33w3JntCmfqW2RG7Y6o1ZKAAgIluzrREO36z468xYxeSK5F60tR5H2LgBsylvvvWbSZ
5DOPl9YJ9kVOil3DX4iNZc5m4qgErVaNfeYei8gghGX8Lv1fhTMHXEcRilb+L1vmzmz0/IzQ2nWQ
wEZBXC7jVyZww5URa1dLz0rtzzQJHJGSZl1A0ksLPaF8+07oDv/RTT1R0A4JI8nIYbxBdLjNYoTp
Web7dXYCzVFzhdegRZjy3+raK99n2Jyll7POrwL04Zjm0EA8GXlHoKoUU1p42LxyCYQw+ISXw6Gl
YALb8sv90cViEZ9amNZKMD7GAAc0/eeBzX9AjZa2Gs/jkTQVMRBq4ZZR4p3WioWytrv7K8DwVEAX
j6rAsdRcqptxrIa3yIxpbmaik6gSIp1tBKur5BdR2x9swTmSGdesSiyiJdnn5pJUkA9BMJaU3Zb2
c7fYZJnAhoLX7TDxMY81d+BSbSM3UQQWrBbuZrfG20QOH6LTsmegUHsD8RJzO/QVpgXiB44RZ4oI
DAPRgHm0t4uu4lmbwAt7Sf1M8Sn6R1iR1mjWTDjkkTLx7zTfOy/Mu3kQpYVfUCakbFW8KYaUGtrm
OOo8krfU7GoWweWi31AqLXWHynjmBGuu0OZ1rOrpnwzNDPFDU9WBJtqoeLZ3tiTkGNHFMARS23TS
vKnTQ8Ye915iKsnh8NgB0VtSuVK34QIqIaMhCrD1Oe93cAi54pH1H0QhjPv6neqqhy18O5SXU1B8
xsHhpcMeXM4t21LWwGdIjonp2G/oJaNp9fq0A2SmNS+L+HHmfDHszYRQdTHl89c9fGzqCpoFKM7N
Uov0A+v5pDe+mo0mKNmtr/jPObHW5gkXosYJQCdszsjtKOonXZlaQgbo5H4pV0wcNQxQZ0DRqfLg
uCHWeNFI16Jvq99O+b6noxoZqYNbZippTExajJ989gj9WGtFBc5yFfFZk05Ok0gJLZ2mXI+rfVyC
e0GUXjHUqBUEX/NLcNAtK0xyZNgIFYakdUa6Mlo5FRTkbXE09f4ITR+MEcjA9m2ZaWTsViZKX2in
6TIG53FMdf4wMrt2YIbqWc8CPqxQIFpsq1anIDTpVvthPANl59YQVsjo0/cEVT9BGohQoRuGYWGq
VRK3/d1V3sUkhXyO/jYn4Acw4Iw6VXXuZo/FoiBQHTsaIZhJ0S/W4F00jy2DvTRVhDFG6G8swNp5
PWM6k3UxatAyTe9LNht9VM5C7naQuSYR+11rmeyXqzm71HSzVUwCwuC2itunD0UTzPtNA/3Squ1e
mqA25Ul8ubtpINOItGygoPPVCcHWArUhcqnq88AaJtXoZf6PHiFtaL/64TXqr+VPPyQM/YjnAbP3
dYERohEwx0CE37PAs3SeAORZG/32bj4P9iL8AMN3Yi+92JVPd8XPHLIXiw1BKLvCFcDRVX8Vbkpz
Bt3OmHUyEJbdhld7gh5jH0R+/f8z5i+dUBXkUKexrBKu2s2QDfin6EC3BM4HBRY/w4+CE1peiEl4
vGGBv1wXVp3ptkTxYdiP54BMjYybxXws1FdnVdwH8p4N2O0JWr7MOAAdBJ2wqqxHJwHYkvVltc/o
m71CIU0djVbUZb+V/w1pmX6lwrTnJ+5lUsqEa89XBJFiBCKlh7cJ9UIYoPgW1J9rN25bwoYk6Sfu
rW1zX3FgzFO78YEzxa5qdHq9SBHtLkVqxtFjjXweV5+IyvXAYYLUX3cHQJXllv9nDwyQpOww6YLu
aoqfHeTnbhbSX3veplPZHViMEOSSpIXldsrhljrNCNIVWkG4tbdK9ogI6iDkAYx9Fp2PvIdiVDy2
OYpLapPJKrXv5emm99mXCktMUck6823tvQLTxL1LHNAOQalIaVd0kfhDfY2nfXDPnL4E+XtQWh3F
lp1pXsx6qFL9oBGEs2V99bqfUmb92JhZCs4bjGqGcRm5Ih/c8zS79CteVAEk4Ssa/htICvZ3sOex
APRLttJYXQcVmfRGeAXDcVYFqfkWabM8M4JpHYPkjUmEO5IjXMmpJbfAU8W6nNfuiKnB6lRTpOSH
BNCf7gqE5sjUa+aPPv5d7HPV+PNnhxf/V9AD8jndcsqhh8Hkxzf27ofqJ8U+k20TDT8eyCY9K818
pvjLqx4aq91130mcdMDh3/xnRfDTqi1z0t8Po75DwjFxyKdvaUYm3JbbPIUmksHhuJ4vPHOtmC4S
cUKnktwb10G6GfM/sGEO40EVAoDlMrTsMej/YOrdil6vaEXvdA1gGeWR31PKBJ+Xek+ITHbH2fjH
xhyRsYrcW4UB0Qb70CjtZ1kwY7sR/GB2ad6Bq1lQ1GJxM+YWvYxSMFoJlReKFXM/oTkQtM5EsoBF
OleYuuQASCLEiDvW+6MhVq3keeYuh534hM5YNmczhc7FkCKE0SmA9OPyxn8PWLKDqJkqIHr8ziQV
g6wNWaJ6s2GkAsQkgRAPjxUqMZ9CC4Hm4QMwBoXDkF2yjyKBGbexidynoYyssxG6gFSx+Gv05z1u
hc6WW68v0rtEYHbFuhCHuvR9ke8En2lP1TJ+yMCXAtTUN++9q1uJD9O4s2wQRnFw7ydXlGy0K2Fa
wmGXkq92oa23+ks3M2eCkx/LAc611fY/ddqk52r5QeWafTWNQY9tAJkGVNfeG+8C+Eb2phNlRhTC
kTYmwMVkWjfmPQJEEfs8/gX0SqvPWt6OE2vm0uaNX7rfGpsivAj1GFZXKJlm8YlgakDLcbW8twtC
VJlOGy9Mm+KnVxlGb7oakBkKRLdn1ZS+G9TVyOYelPmd2G49iP0vY8HWcBuo36L0uzdoBW1pAs+j
k8fiJQQG1FUX8PLqY0oJLVcQDt5MggfVbsL8oNQaVE3TiI0VnXER4gdUlhhMIhRXp6W1k1FlcXn2
rPsp9PQSw5aHUeY0N2S2Tl3XWUD0vRf8LVQVCj3npvVcuiIfm9S4zip9WX8K0bxdZxKYRWgzoOnJ
Y757u0l527J276CQkuD4oGCKSHc3akVO97GcOmyQzeDYD/l/D3rqNhlvCgWCQ0mk3QcTgTP5+5RO
qL7rHw+PvL/D8hBxNtJJcXCTFRxmTsnuuVHCyfZdJkf1zsjr3MrylxcEEWfgeE+WQEnxzyfjN5D9
i3wNHqFxGUGxMq3YteuR/ypRReEIA/Vt3vHWxJmxZu4nvqr5TS4V2MYCiTGLjDZFrrUSBAOB+8HP
L1I+9r2H2HQEs3ZCrgurL+Nqe8Z2nyAb+Y/YuGhlSKrzpbi0uGOLuuvi9ZdVuPBd+eUHoYdPb+YB
r8j+bR9AzmQuVRPJFa22jVHHZXfd6CWH9HzjCSQv2rOg2hWQjNqb3FUSZUGhfII/cG7jUXXioFrh
Uvyzfxxe+93e6HN57IJ2wh4+oz8eJ0VXhvG8Nwejqv2H9sHcWTSixOPfrU/VR/PkZ6/Fr9YwLXSv
D6iolgp10TgrnyQCr8InN9Rj8VK5qglNSRpUEZj5uY/h9qDjvXyBqIyu4hpXm/NXt2GrsfXqJcS/
t781ityLPWq93Yaj+2H9R8+XbOuZ5W+qhyRlRew93/jswRr1sHXCUpRSrcSp4+5mpep+r2+ktACz
ayXldK8Kdi+9htLVLhSaepR6BeLKUrpg2A1dFZV2GwW4z+9rpTc75rS4QxXGJxqlPaXvJUMQ7Ioy
vZgfBxPHeu/6bRNmzEnkjtWUtnwVdo+fwSBeoADACp+Y63qigdExk3QOTbJH/GA+31EdbL3H4Glu
qh1BfzsF5jAARiQhKuiJdXq0md1oFGlUT/hh4WLEFXgn0X7MTDP8eYZTis3MMEFueDAB2FzkVQCs
6NE1sBj0dSwDOkDqxhC4JpgVgDBmQiltDi9SVDVttJTD6E4iqv6i/XVKEWAe4P0yJv2RrgAXgsNY
8s8gTk5hc/XskqKsDmeKeWPUIX7sH+7Cpch3EthWEzuEwTqtkv98PoRRhFmRWDbimFYahoStyGVp
cTEsN1YZozEzLoXN/sVvbay5uow0T/3IgWxQAqFgKpLThN23fhVpCGy0lWEVzAy+SCtbfbLg1NAy
+Ih2JUU9HMo0coBAagmAhD/HzFl3Hd07dBBmPmha4XFz4vg7qaJzoLytwF2vyzXqTBAhI8WKvx6r
Xg7xaXfUrXPY6gWFRqJ2+ZBGWS1kflgLr6bODWB+uMitiXGkqcV2tQaUhR1pBnNucSSpAw0cjNVw
LZj7qYHiP3yADNhXsw7Lbv+O3DtdwiPAUarvQdtvFHB/0h0Mr82JMm1z+WOujKf2bXMq96FVrziX
ToKoE+/r3STlxjhTmy8vK+b2f/aRC4QCzEVAdL+T8s3fPfihATmHkYv/Fdo69hImK0V+zCgZL0y2
9KO+TDeSbVGlPBlBWkpUKHkNknA9GZzTZr6MCpKhCKWZigUBkVcimLtwuC1iRbVQt+Gu13epPQYO
o4RPtN+VZf7fZaa+M0iVlbnhFCNVJ90DjJnQ2WGpE4oFkvWqM4ocCmG3FuaFnQSJGZD+6iCX3RM4
fFVq/I6Ak/DUa43wq9MiUwmdgfjgpJ6ZHq0uPq0mAxTE7AFaKG4HhLX1KnEx6K9Y3xPf3xe7kKvd
IAC8KiEwPmlqko6B/4bOY6PpmidwgriSQAX5RYZzdDo8F8IxBn27X3CQdcu3ZgCp46RWNhbr7UKl
6BWGlZUI3XcroLaVibLggNnEbPYiEnKw1gyg3eJiBHkS5aV4EvWYFXRawmpOaNLnGzqBPcC1Ca4X
sZei6rhd2oSnA21FQL4GXAkpdmHcEtxkKjBk1CvIYX/DvAftPLICr/gmlZgxsM6L2I8wEcvmBhhV
LPRf151MiffkGDgrrSapUUK8ME5ZQoZo3UTh2nKbVu2rEoODHwlpSz/jwhKW0QbSnKfn2D/+GQGG
98AvGQuOGHjy4I0L7n9bs5oaDhs9+GDRTDzGMa1fpl4I/36dGN48HWyMc3GmoVXpSPPNP+pLeozj
MMjejf/r8TwUHk1ST53sfSjNJ3HKp++7BQou52f+Ou1DKqtxBEk6ybroYpav3Ly1UH27HPiP3U0B
3PWZSfSgb0M2u/Vh8tpJk/H3Dn8Uzj88mRtLBLVwJNYTrK2PpSMoq+FwgSdAfLLmfOdW4LS/zj8m
RQdmU5yLs/10qSpxviVYAju4pe7N5mdtrrgXxzR4csfuoFIKHo/WenjbFS6YB6Wb/hae6G3fLPOP
Ao2oKzjJVp+bWMZPChJSnh8Q65Zwri6k9nhdEEKwWxeKe2BBQN7iJwZdFyxALscw5ndnLewcjubi
Nh9HPBmopTQACP60DA/V0g82Te8RRO2gxgjbddsydL/Oz0BUpAur/TRSQsoSzaMApsElx/5ql7xu
h18Df2JOO2A2fFOa2oX3laAigsD3cJ231UaRgEmdzIEzxAXFGGexEuEBVqVBlhVwRN00og4OElwa
0UxCIP3nhyEGFRGXoQ8nspMGR8p2NSy4w/IpYjdIzGMSjoBl8XLHy7DGihrDTjUEW8LzjKVXkSOX
mWvTTFzXhwjMJ6KBr7pi1KbclKRFIzC36sLRFTztqMDeevKX4TgDXeOlKLmgkUkbp5xcm9CGcLnF
bmM9PWT6cOWQeAd5vm23cwIXj+PeHMXLuG/G6YzXKPvNyshlvLexlyOWRIDcjvlb5Cw5xxNX5wmc
0uN6qQRrcJu/VQRgBregXHGQhiaJRfbneNRu7X0FU5THXXmQxMH9WaDBV0Ussn+mFjgW6YRaws6F
Pq07lYQJm2UgJlGqBfmOeOiyYvQ4+sKFZ2DhZTeUMKb00HxcKUZwjN3zVb/tDslYevvHzgaTLCva
q++2eSiLPEvOaCSJwn9RMs1WkB5brgfbZyd6rW+kU77L35Cye9NVRM9xremAQRin6cN+ca9/4HPi
ocSFm+dLHzBx/ChW00vPOkalE9DPnYVeI5pzBCkTyUhjf/K7v8Qd+QEzyZrxA08EZLnX1fH8EDsJ
I4lWZiRjDHg1eXgtAkVr5TzhyVDMoo+WrvXIlodOD5379tie2BkJBSmOuJU2Y1XX3EIbcmFRoHUu
ay3eahOEYNhwA3yaNCta7qye6gbouNcepDI7tlR2+q4B2dK0NEHDYBIDRgYYPEGBHmuKpG64HxYv
qM9L//e5OMgDA1fITeqT3u3Je+iSlbwbX7Fg1UZg09Yfkx5HFkY1qUsKTSsAcyZRP5uPtBbBIA9+
cus2qO4jfpYyW0LQIrzUgJIZnVCrJEtGWd4TUbDialkJipVYav3BCNC/0Zy5bKZPaRotPL6J5ltB
ZRqkibObNQPO0AGNquEHPuwtsPktPJWYbwZtAcnkFf62ltq1oIUEHAfYKCcQ2G5l8Fy3NHEWs7ZU
2wY/o6YDGJYWE3vFrwOcFEvXsrz3KZq8oxeQFlKjeVJCmY4c075uarJkRjoe1kvT+rUykEm4uXF5
PeA4vdWToa34gGq7EvT+inKN+MNfBODYLwG6yQ/LoMlRd/XTpvVG++j8MmIw+Do37KLg4di8ga2u
m8nti+EkmoQCtIcPyo7G3l0BMgrqwNgcbu97yXkPefwvYke9zcZqPvPpEla5UIEvmSahhKGFVpTP
WVhY1Hm8jmwIDm7rWhyfWK+ckIecTF95xoDEE5eHSe2feQFqNyYnKmKtWtKntKHSzdjKfxE5y62e
8R+xlNxbYeVR0g1OejM637m0lGbyGpyFhqYSZdcicHkEZjfQNK4nbgrxLS/i3rC5zC6DvqGfL2Mq
XEBpZ6loJ+abGR/LMxmCicP1mXnTKAH9hDzImVYYLHCo96kbxKrlWzt43ywz1SJbW1ZCnsmLRdhQ
5GMs4SHmLGoNnbUJVqZvbau2/yMGPGfWtSTg3rg3wOvIB4yALgO/retNbQFOm1PF1IzdNVp3WVUB
fE1UrEqzR+hnhxLEk/wgBeIHXuvuyfPTLk5cRihb6buMz8CfFjjEbX4O1wrodkFM0UF1TRvsSCVG
YJX7dUBDkcAg64lpAuVZGz0TxzXUjWAt1OC2kGy7y76RFazHGX6FtQmOFLPtRE/DSPrTiRZfNwsV
+FJs6yIiIYCyFAKJKnI62VyU6ZY+W0P3QJDjOWi/2X+Mcsgam8llEK0yW/d0F1eBWLBntba4qsNt
OEl3cq6kvV9yD92snLkrhmrnuX4OUoFQJTE4OHO06DVUaG67sSD0bJUMGuWYe/KIHnkwGekMe/6f
4ueHyEavqHJnv6cEhawwJciU1i3xXZIlYayQE0kMirCAbUj256EGTDC6vjcNHAAjVCmmu/S8ChcC
scQKhFlZcqtXJDPNJfuaJxoVbWGnLy0Lr+5s9UiDp1l5uEIwlYMRnyG33uPntETrR91xDFeNQikh
Jrv5KZpN/ZERXRFzWQDEGGQl17cuH06V8KkB3RDtlx7lZzL8H/HBtuKfMf53j92RIh+naQs4PcCj
FoujjoQ/TxdSPqJIDr9LQcJcs/R6h5Fq4f9NRAXKS4nBgT8CVbXUC6vu7xmUb1uwJ6cBZMsyOsM7
egCqpA+cIxF78bE5YHHu/jRiYnLDN3cWgQSG701ySmWYUu9u1TSBkl5Tqllb3J+wTJlV9tJKXKHm
vaZ5Hg8oCRQoW86D8oY6ie7QrbuTZFebc2sVf32nPy9j9EtfbwqYW77SgX89bjulogbjd/a+Rhz1
WMf5SOw2dE8NH4iSt7W1nKTNioXz5cUKQtyYAR16pCZIWV2iM6VYPOUhas5MgiINxLXdV21yLirn
Mrk9o3jZpIteGbHQZma+rj20foAEP8MdKcqXtaB+36CbVr/SmkZGoEHS3UR+0RKqglqMhMEoHhG/
BhB9pqkdKjxLyJyUygWfLcVUs36dtpoMFtJquhjl0PK7VR2sQfAG0Tbr8ghkU7ltM+LbPvBoIRug
JL7cNTj0NKaqBbieWFTPpxUAXP95eM2p0cgB+NWVMupcCXMnL1XgjwoBq+iDoeEHedu4fxjs2UKQ
ONbrPgyTjb1NOgunXaSjUSC6MiPt3+d85Hl25rN70TvbqSzWKL7afzLFW3kbN4BW95dqvDCM3Upm
bzlIHbzoPdIJyzavezNOrIfz0QOUB3S8emdQ4i4z21MyoQmMiZ62xrloOIG7yGaw8k2dcGRDUQjW
4G5K2rz4xHJvwAbehuyY7sWoOBwgJ5j7qH7X9x3ACDXN88327m1J56KVdlG+IUHGxiLiOtBRNt5T
AefXMZUN6s4esevWv+hIXRSCg+rwwwbmONm9iGTwOTtf2si+660z8G6NVJrpCd1NyLlzoKFs1GRg
k5EioiGUIxiqzC0/lMOcFJQ/mGtIHhQrYXFqzpk2SIqTTEZi1Zskn5uvm6Je4DXCeYG2iSJqEyNv
OXdQXDMaqqODx1sQXSXb7R0wG73ifsOL4ab3KiDz3/d/zn9zFhD2G+naDUkqzKNVfEXF1ZRURdnK
lfDaHH9+4MYGOWdJL9eVCqdxYEVu1JiIcnmTjXLVWMGDjpmwYV6c+XYRQJoEOXodQjHTM1i1Nf+5
A+z/RFpIhNJEvzYVuAzg3dhrxdZZUWrTEdXLNLMZzjObA2H1YbRw49HAIwMnoA3GLy04r/JHW2nt
BaXyrFpgMFvtQScf8oYvg1xZ9IWRoQaz8WZYaxMDgPYQ9JLTUc4DwNm1DcucR8r6zCRVgsaJgDEJ
ZyoPIomsFezaGgMGW8JzjyIFHaAofw4mapRDbxXk1lpl7M7Ip6+fWpGfw0NwcU1C98K1gZLn/jwS
xLqkknLVCKpb9FwCqPynwk5TxmjUxLUPPd5//rgCcTIE+GiU+K5YYSvMbYWwwEIb/VRg3T/Ca0dY
YlIhFC9aepDM0iOSrwk+OOlv+tyHGZevkw9mwylfw9/dszgr6HmdzTVvtqxZ6t4PZ+25l9yB6bAS
2Xygx6JjG/0hgQZl6T0FmNc4UgPaMWqOesXlj1I9iREzHReoFMGnGp9XKClipOi91WJvRMsP+fZR
Kv3r+NPZeZ699PW0+LtUZlePwXoDI+hq1czFV6AzxwLGeUsP35mhW8bHI1Dw2/vvp7iTHcKwqnEi
dr4VONAyGJFgIyk7edZwgwRMVAS/Hs4FTAJeMZEd13ufHREfCTzFAzLuaP99ltJdbSax0mq7jLZn
vessodn87rJDtMgWu2r9JNUt8YYmx2v/rqHWu5HT+zsVrFCdV1BwJM35fZskQWeW+NK6rcEOARxX
HlHSCkC5q9oADspi/6ugduaMDgImHpKDrUWw7GB7ePAyaOoXK11ckRn8nu/f++5rVRa0kfpnWw4/
pu8koeaTnr9dSphoS75/KnGd2kK8Ycdm0mDw7fYukfXU0zflTv014sOH2nGnxKl8GIAjwWYB/xvn
jIZzzblb0MM1Qs/cTTrwwHUeOBtry6WchX8wl5bUoLLC4EiDhusunGkNizG7UUp8Bm60Aru0o34I
LobMSmqzyT4ovaSrlVfHhL/KhFFen53o0v6MpMZSLX19ReSk7SsJhAXd/NPgZbXlB+r4+xA4bQpG
Jl8NikNff8ucuFuCU7AWGDmL42N01nYPUOZ0bK2egvF0M5nv3eGcOM7meEDsEgA68Nfy6Dr9PZZs
S4x4dIAiIPWg241wccRlhlsFS7ZTzSZeNc+h+9CUo7ueZcbZRuRcAW5bSENdGv4t7qczWGROeaXg
Q8qMBLhLCVQ58t2Hv5no3j125Uvv3cxMNPtUXp8af21aUaqOsW6mgH8NkwLsF8TxLGmWRPlrmrSa
LeGbGU7xXiPz/XufU8pcywLKikiv7GjTgZ4Zo5O/bdliBSJy08CO6RlLt10/UvY5vjCuRTUA0LEw
F78LLMyiXyOWM1p+8h/FYEqtkTrjNPmqT0EjAkN34401qWa+9N0gBeyx5/DUadTy1rHfDQAR/YF6
Z95XwK1+1v0O7i0ThQ39fOUbHlN8SAcgOC/XYx6LuonN5ty4q7rrcL4yzBIwYMm+DVfxJ1k+aRHW
52mmBilnC1c8inKq/yKGiriDeTRHwo0lmDkpdFHqN0DYLo4C0eLDToLFzzbyyHpBZHjQZfox2wAG
Vw5tgNcZdlOzuK1DSWP4ww3jTgCTxxKrg1ACtVaVtEgi5kW8TbdNVeaVkH2miGbCEu/fDlo2KF/2
GQmlaqS9hlMCd2WSHT4x/vCl7Thzn39flD1u2etTGu3Q8vmxvgDSTHhNbBHVfKX1QYFKPU4apt2i
vTXpwXMP4rXf0Qn5IrL49qWoUNWwjkhnLlpVYsDNRxR8mRs/i99FQutarAhSTUO7JVVqMsvVFG7w
Bicu2vCOVCmLHOxPd/ORJKkwSjhsuynSiLNOHi0ncfg1j3NWviLvcAE5R46X60wpun5ifMQSH/rE
9drrqKum4cYtTzhlu9Dxfyd+KsgV5aKDhT26a/azDHEbd1MsZ5xasuUpr4tSdDTJ+qKtPxJCuMig
C0vf3XCyxHhBBd2g2a4x/XcNI6fsQwuBNLH8O1WTc5jBoSgFrMqtXV2yTeDA0aJ2r/BRh179iK1O
OxbNqIu7dBylg6V2enZ4L35cL8zp/IBVaVXgcjtVRjALXVweQZ1Apj5zjoNBGcBTwEkcfhdHWROm
JTYp461wh3XT7RxmHPrcpRaMo33qv0fOzrZ1FievrH6ttTC2PsxftDYWVmffQS6HofRVHy6c/LJz
kVCpkZtEWRDdTeeTOrVD0QjSJuMz7LojZVXEq7ZU4XVn3D8mfIvxdOwKJM3sJwZK7NnQPMOL4A1J
yX4hGYupDwt4+iyMLMazgIQTvldEf2LO1ZZ+o4ur9JovJcIh1+DjxpDSJoqdXCoL909awkfXUW+P
ZuYMhuECEGGemeQkALyGoXqkMJ8y7h5+td8VyABNp3YU9dqTzJgoJ2ksH3HgmkFmIcAHEXu9OFEF
oTR+gFZKIgvWle6yHbGiL+nag+BzWtoePViRFwetb1JMfCF3OFQeWL3iHmgkYPMxaXE32ZhBomRj
hqFQdicIowxiG+SY3DBW3RFGaL01yS/im0wcyr0NIUgk4sG987E1jmmqwDzNJEd/y7OXrLnHfz7C
Z/KMQRi0LIcZlxdym1ROli/kT2T8gjyBvZzJQZUErDoFYc6YiiPbN10piwE/Znpu7uZI0lUacisc
Lkxle2mE9CpFUwJV1scNe1CUZhKOE3g5TRaUh8QYctonUi6XnZfKR2R6LEuxy4qOeP6hjYjzD5ua
+FfKVQqZa3pzUAMJrBRYxqkscGQUwcQRKZeOrI4RhpBp7VZOz4LaV1PA/wBdx8YLQvUXLaAVnYX2
OgoU0QMyXZxDwNxmZq0jA+21LydmI5uDKst0OUKdjmIiA9LdbIp7Ul/Z+alF95LtaO/ksQ8nNSST
TbzS1PfjmVkBTCzApxkpNH3fWkne55oMw2DKtgwa0vo1mU6KryVSf9BC28rHkCm7nKVEhIZ2DPnB
hsFUIs+n7RJRGaCeWYaNjUhf84YceDp0VMnG/8u6/Y20pFEQpZ0OROPJPUBbhHVlaYxmP6GryftL
zcsp/QTq4rZIMHe/nlc6N7YFo71UdoYFrFBA4K25AD+cTbK/wvfOaUuuUDKEiLoiKjszEg2SDABo
OhEdxtyNgCf8c1R9OUrWmAjLKEKwJrgGl6xGf3NLoJcfYm4gHdYvEVN2+bA3wTIbixwdXcylYEgZ
A4P1ANbwJiSt1uM6mMm4d8zMaNZW/TEPUregmjqMPK7SlL3lBc8oRbCzrfAU/osIv7HOe+S7dZSc
OEykAUhVhQ3gTB53fAJjuWia7Gdzw4sJy4vCCc837sgmqlW+eaLAGwKOUIt3fIaHCATCVtzIHu73
w/5UdocmShp40C9Su/H4NePUgF97EJFrFN0/MUvTLXpEk9z9gYsM8H5TXMfF5hcng2j5Nkqt1Coy
5V954jYsCYWPZ7SdAYqk2Ot98oWrWpwzEEnO/BlQVVLPOXHV87FKiPqyq6Q6QsxiFLPQIrvVyHpI
NkXtkNLBlvUx+CJGyKjW0foQo4wKpIBiKgzSNIKn3aKPE18d3Jre+MMbqzIwZKV9tjzuJWKdetHm
igWTB4PeF6h2aJiUnJuuT1A5UqM7qHdMwonRFNSZ2RBLYBQAPSO2wM6zV1XzIxJWVkYUNZHV5GrO
bGnVUUzCB4BW6JSvYWqbrkZUdcBABmK5TauGZskWuOKDye+TT93kl84jwnOQldai9BOTryo7V9dy
hic0hIW7TsPxu9Yu9cePqPtaLxHQsQnpb5wNr5WbQzDUPH0+4SBc4piYq6OsDMmniBEZuah5kHKM
/IDEB259evWSZ26STCiOI3IIHyKUDDwggaJiIrtZNRfeBPyFwoXvOnQQfQWUPZUpOS5KyNEn5AFc
HtDTsx7t9/M8MTA5a6+fbFCCFf4jWHmvifd/V1qDTeBDnX3z5EcaffyDPRYnDX+fTP1kGvJoWKmS
H86Q/GZjpssTztS76BgWiKksvRCJBJBberqK4aiuYx6uPyxLk/KsbDEYAjqcUOIMn266q1G6qT/j
vK2numlJY4GgBIccw5AEJ9gCpcu9uFO1RT7L1NwnVvv29anATKa22ZzUJPeQQZq/YP/ivCeVk6p1
hxuLvD/Sy6O/52XKzqtUwDPb4vLAkN8b7ABokgKOZPnpBqWIKMZOE4fZDb5jUcLJbn+5Dt1iuzmf
RDHIziN9mJJnHTWa49idLMoY8Kaoqm5RmQZeCqL5IpxS7sqHkm7Pv+PvU2En5HEe6b/ZrYJzrrBP
Yw9yDzw8NP7umtrmoP8/T2tFPUXX7Avr7ICInSxlrNNuSysaVCnaP9OO7wsQDfZITbHNaZuaW7Su
77URZ0PrV9+65RT8nnX9/Puyxil8u5q8eZE+hPvjgB9tpcN5u76gh5WmG6HBO2lBbVmHBdSV+Bi9
2TdeCwcrMiTkqFSph0AYJQ2CbC+31LsHcX83Tj/EfXgYI6LjfqGS+uqgri7Vt2vt4J0Z8tTm1TeE
I7HTxMPlpKITiI3FUrNk3F+G6hF8ZYa11WKRwqMV9eTTgvowTz3gZo/gHk4fKwGcs6GLLtm4r8IQ
M/HYRNGAyEAv/h2Wk0t3DudVqUQY21jMipPhsYNtSqdnVgeV3CO4nFx1HKUX7vzaLACDq8b32J6Z
Aac+IuicnuQVJy7k9cEkiWrlokq8H9yCbqW1f6BbklE5MxgW13+ffdb/qP6xsgqRoCIYI0+so5qz
qZESaituKDWY1WoqnYO/x+WIaQhjUh17T+MUFBSWuNBDjoDsPVlGBJtWjiPEdekMpYTJTtthZdlK
8/BqJlo23QmJVN3lTlD61A2rHN4SYXFoUnY54C+ZxlElY7CdJM6LV2V2WLq7xmSrkPIJ6IdUZ6NB
xWuMQg6glfS3FsMz/Jy9LLxHasZIVtLZXT9SS1fL2CyF8UPC7fuh2k2v7ayiT+yvt0P3byruTlcb
1pOXGbWZGhFuCgVnVxmZYEYytD6zQJJFSAL92HQ3PbSx6zt/a4sdROHjb6yA9G/KIavM7MqeYmwx
U4bQnKOCiKXLcr6FK3gCowsA43sVN58pl8UjbfeGJAccAcCe97Oyzf7TcuVUXh9r7cazWnCW5Hff
MIDFuqlwqIZJl17VgF2gjlqlqKv9D1eVtUrusQqKSfNrqqSH8im7PMQBVou6pc93LFG1JSbkgReX
qnlGA1IiziB/fNvs41eVwbI9wTRZmvwPPtEEMLhObnIamJoQcbYIPilaSpY8wKWdjs0n09hq5a8H
6VuIyHVUfYz4IhSodlNLpce9Tl3XpfqixFAmxwQs+Elqt8Ot2V25fBZPlCE6HJpcQReh04zjsq6Y
nCt1pU27Bdz7Y7AgbMvdM3jcFCIpBnS7vCPMfDWK/JzVNHmumEElbJ+ekNQm1dJ2SZi1q+fOJUzX
FWv+2Z/X7v592FG/UeOi/4aLWLlmip+Oo3MYCWe5suE7kpsbL1yqYCkxGDJ9JqhmsG0YaqFYWwD1
GULOzUpOHxL0KOvDRFLlLqHrHZnBeXl9ENkPs6yApZ1Xp4CM1tcqMFcHTdz1egtMyUkeqNdSonWG
CVywd12ov5kJCOZ14EGhtLZvUxdN6aUV86dXhNkIUstboqmy6J7GIi/Q1/p68sYj50MkRWRWDXeu
MapdozIN5f1UydybZRjTxEcg9RBdoUZnK0hfbRy0k74kkzDV0mlnpPwPfSq03CFDR76MyG8jU1Bm
xDuUlCSLMsmXqM/4aTaZdmtsbpQyKw2FWDTtt9tQgOQZ/UAPLvHAB/bnZS/2SWzsDWKs+jGYZGvW
VQ6yIIYlV8wQikmvrJi7WKss/Zag6IghCEZcSuGU/5pI3zii3mvqsvksGgvxWDrVc/zbp+07Z4Th
4xoA4Mb+sOkC4CFvcUOX8j7IBPVTsgM0J86xn5cSl6hwJYCfbQyGqWIpP1n+cO0jXjUpR8Wy0uY9
oJwE4P5lSIpjoZ0kV9TRoNGdW7/n6UrDfQ3y0bRPWosr1axuY42YSssidT+wSf7OGXDAHXBZy0RJ
lkgzqy/sIEKRu5ftwB7OYRIHr7JKLASpVt758W/OjLQ+KH79yLsRFBN2EOihFAEfAocgZhXxgyrI
rUlfxOR2tVtZbG4+UGuRfJMvbtFglPFAy0c2WGMiIaZf7/vv339ToLQ8SwYGYM/V4uarzS5SoMiK
UfkCp8bDNasYB74eUavJaMDmy16dqfaSMOrdpTigDXsUbARyelcwbmTrw9r05tV4io09LxTCKoHh
KBLI2dqz07vh1UItDtvSUcR9Nug/8HD8kL28Yw+MU7jlvvuVwVN1MTQbe+R+iL4kbCeH3uQJYimy
DOd3S29pU6nxbTOKd5E3NtvvIWi5ltvyxoVnnCOUXxhec6CSO2rnXFX27r9LVhOysxkhc2W4efD5
1TXfGfrKfb8HMPugQu+aD+hQjg1OqMxOoxJWan4iEDpS63WlO8ovQA11lRwc42hbG/FbkC1rmJeN
hjHB8WyZ70cOsEbTEIdOpSe/Y67QVCbUQjVdFkgfyYQZuza8H3NGOyIl6WPUR29ZUFpiI9HMlwTa
jXixc91OB3+FsL4xNN6meKCDtW/uuK2gWNAE4rrXr5e0/lqVD1kPIDgjLlYvY1vshpl/1nNAiX1y
tP+A32ZDPRO8pjKfb8vJtDNdSQxbMbt0uDGlR3RG/nGikDUQ1/8eTyM4Fzd7rS6gpTx//vaHQU+1
IHsAMphAvdB99HQWJW0FywMkMVTS+3i5Qi1+y42cQ4zhOMdDh9G58TdUvKuz6O1Dl6Luau2KlUpH
UoO3UX8prBdFARy0uiXxOvsTLpP/aBMjdJc25fi/7y1Kdo+RH3BUFE0ax3/ZMD/Gn+Bh26FxVKIv
fnDRh5uchfvO1ZrteoGQyKJNlat8zW56KXVWEI0qF1nPSpWPazbFg3gUeJeZErwXAXjFNJKsADfm
qJTjZEbO3rgwoNK1NlmD+jnFiqGJvlqn801Nm3gV/NzPEt8G2moFyzd6N+kFW04qIlFfC1I04imZ
Hw4Ws0AvIax6ebmHWcjxZvTGQ7ZGOOj1xat9XzfAgQMZ9LkofcAYjoZ+z4+OYGySXp2MrhLHLZ/C
17A+WjNT/WNdsPggTOI0bLQYJYg3Qo9pTEsp+meTHT8fF4cqPHwNgPWvbx6z3579BKVvThEyJ8RJ
AUXVPywAwlvg7mObfg+ZDpS8FJYOl6u+uGnC8uqrDijSgk3pvOOALsutUXfSkI5tPFFGH6dxULez
RfFtOSnIzSYf2L8k6pJYC/B1R1k04n0WXRMTrPvm6vWaejS8v9cPMmrb7SQax6Qe25yc94GnwtlR
+ew9ayrT8Pk35yX/pAkcpupzGYfpFI3JXyTkKbbRALbneZjShqMpG8HEANr83iU9PUEdRtGl0nt4
H1d8GRIJLG/AIR9wZ+NTLRcYVeBNHIdlmNtqjmTfgwYrJn3ThJ7Z9D0pzQqyaWjlD9J2ywi2AnHu
SZ4efHF/RLjchfqiz0shzJXrcnc3Wdoobpn7bWBieBJ23fG0tGECjFSFJunVt/+SC6KAB0w+hAOY
EpzMkQSFOaMk0nnHY3ck+ZhmFLsIthpbhtpJhLCGXK2F+JNd+614Uh+9sogl108Daw5Ib1serhwS
HNyvSDEY4K/tTZSYa/1iC5J16X4wu2yqNN93PwK3srv5CweAE6vwlzQ3YTVXHABmYzq/WvS9zf/l
0TxpdcODbxTpkSGwwY5amzFdXZ0wtAoJU7nOj7d/qEb/cgLkH+s8wX3MQz0gJFWVeWCbJkYN+uSF
MaAF0v3cfnqe5r+vzqrzzyjDJKGdVAyJg25/GX9y2guo56gGsWqufluL5fjLqz//JGwEuKDvXjFf
starKb77UGSC6ML6TNdvboPI/umOmalUCf+Ej+TNgLneVG4K++8gkjfx6J/L9ID4J0mwvYG7wWNg
0sAuCKgSKYSJbj6zMLcFEQ8eqlYBu6RCUry36nq29HNB9CQ+a8TWrnmci1Y9iwjXvw37eubXY00P
IIF2yJPWtLqW3fTOeVZlhcR5ZKFr2oDtnG7Hmfb473+saINq7R6F1CoDo12CNTyX8Ixr22yX67wq
OfqjngdZDaL2FxpbDWTQaJ77HRj6GZEhXAKVvjdIcSZaYW0Nlcx9OfxcxNhtLItWzZveD6awaKoo
KOqoqTVldY+eP/9sTCLi0xNwGc2QBzW0PS33oMRLq8hg+Esh70+ew8X22keFRUKl8XGtTVPNmxUa
Qmi/QlsUcT32h5UjgdDy0ndmm+VhZ71FExmgTJmLmubeSbMFgUoT72XSD3EWY5UlSrSKMroikNCp
ChO6D4waLiOGXVrwWL0D5Lf2nwXNkadHz8CjSmRNkwZkYSFD/fpFzzLNDND+/+yVyhDqAPol8gyC
rZTA8F85gWip6saKZjAwwt8eyLn4DeZVzXBg2/tobNIwrgDsAswF7ZbcrTGsyXnujqKi5X3uNbeL
rCwgtYseyIK7UT0kzi5Hyl3MxyXwMuUmx4VCnOpl0u+8inemQzSpRgmTwqP/8zytacvCHngvT8lk
LvuGESdz204UntMcWKQFz34qYXeWKtqeLWQYng+9DP/q+G0F5W4uo45hnVRlZ3shv/lDL2PaMJtE
ExirhdZ9kPnm/kuTb5HFGc8+TdyZx9+GXQeGAqich11/iWdUe61wKT0Nk7E/KwCJSieX7N++i+/5
U5/sc09oxmRxwNhYzJhxZ8Vrx5gEBAd8QWbqhDiSiX67JyWSUfH6ltK6NUNOHQ6GTRdOTYtmiR54
iFe/t9eIP4GAoxaiC4v9TJVPS1FP2ebbEW7+Xs+d8fhf6u8FJmynyoCr/NWhLQziLxpzzjE/X9SN
Bob/Y+90CsJTyNh8r+5Zq0S4akGXhr8SF++kIJMym5Re5P6qd6inLN4K2XZ+LHQSJBrPjErHAATG
EpHJrB4Ji8EDdSRC4nm9YPG0O0KTspmEBTm+DZ1plE31ptNzHId/LlvV3M9+qnI2k4hbjz6V2Gok
5L08ypEUjw93Qw5QtGDjvDg1c40uf4EglqtEJJCpVxupf0BKIddM+PxAvqChaTLoStB0g37E82uM
CRoPPEvrLaCLUcW55f3GkL7ya/eFTXeRXiYhlVGeYBP8dQEa/fl58lN4VHH1mxeP5dJKJL1t03I1
lUZUYP9ktigaOUEP
`protect end_protected

