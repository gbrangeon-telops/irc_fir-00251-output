

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PT1CWY3UnkDDUklMeaNBhV6BliNbBJfbhqNG4kOV7Gat9/z6WihgIxC6lRE+3ldfsLvMpYhy8uJ+
25GNPlskPg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UvJJPlyuv70VHT4mYaiqDRKTOeGm/bTLqTJOIy8dhI7h8MQzd+YE6IQThFVGwKNg1149OMGabrJO
oYkVzjNGF4B9Aleco2wvOpKfvWGZDwt0GGcY0bPwCYhgwzblbjwmCgPjWkv54osNVTW8DzqpXiHT
yqTtBlllC+UP6StZLKk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IvSnqjuvUH0Q1DG87naNrsoN4LstR88Fpjj6aMMwh+f6Fho6xAvTtV8qJudD702FeycqdNzlt1ai
QXhCNPnT2uuSCS75+mdCpNaXrbRjxmX/iWoxCnzawaHjNORHnFYbE5ycb12Je0b7xDgqmfK+x/mm
Rr1i9nWC3k0y2ultNBrqag9B7JWz2UiAxNLz9gIhkdjfo9uuq7n44on8tD92VMcRgnjXzhfwsV/R
WQcm7g2SVj3bLFjNpwKO0qkV9egUmW/eEov7KDZj0D4B6HRqmpo2DevGwrEmNSVhbBsv+hYHPySs
vJezY6TBoybQdPcPOmulaKi4zQJv0qMBHUSRhA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
N4Lf2o4qQIsZJ5JVKzqV74g/C10RJITmHA7UkLNDA0jMmd38lQ4sUVhO++1w0lqqkNK7gbVbdw+5
aHqNf15gjyNPjYW1ZhVXHrYiWWCWKhn1CmdTyUXz9OVBdu2lqmPJnjbOZQNbhaspal62bK34xeW5
H7uey4lH4qjMdyRPWyo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WmWXhlbOXU4TrFQt6FbjizC0tiQugH2eLLLRZI3zQRGusS+51Hgzx4mz/p2wkOrjF/inwb9EGctX
9EIb301sFgIc2+iI7RGNXRFy/HDMZa7bViPHFvPX6IIbSblSMhaUsZnDGZ9ShEIypX3t04pywLmp
oC8cxeW8KJ9jku9s++a0XQ670LJrlDd/u67e8zo+xwxrAToVkNJSGwQcgXMc9YDwrXqUemdrJGhD
qf93Ms52+vFz6ikE9Bpwux97WA69cn9Tx5Hhj95T7V3DeqQDYaa0G162sFOeOncPAYjRFsxSNp5b
cwcMCxbjJE/oLyWzhKmrRPek289fPpANZ4f0zQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45744)
`protect data_block
4T9g5R6VHyoM/D5OHqruSANKRPAYzkCFbQMRgusSmBNKHwX1eXbQHZ7lkEALj3MvckqdIczWvAJg
raudSzFaOmE0RH+YIoXIXFw3QnBD4vqGOjRTFSClGfkg3h3FNIr8g4H1db9ro1kRlx2IXR/bG70K
IP9jA1mERBJ2FxCYcLoDiQKyTkPDlLF/Il+8oir56ZYswzVG4cUnTUGQX8TCN/Ny5m0qfmCs9TOB
1co4VypSZQx+Nh9zmWUdpo+sOKmRJUz8ed0mTqLE3pMIL3mjnaD2lhNi1RG6OPTvZxi9i+e3lAkJ
ydLWEjBkdyaXeXVP3DVMev+dRj9WHxdtQRRoiaCpEP5bwVlAgnmzbHVvzLV0j0RuZhlxRsOuW/YW
OdrCWUYgLA3SJ0IQI+wbElNJbi6sCWUFfDhijasYTF9TUV74asfojWZEka6pwPxZpTN7129qQYep
tI867t0wvVm/Y+f772rZxD0IVM27olQpw8kxFP3IMu9bqFwddhmCEAjR0SZu0KEuLzvksC27tqPy
FpkOtWKAcBP9WJgBQA3RTyCiRNG06GH/XXR5oOzji3PRHULNXfesl8UhrocaAIij73nh6ir4fzNQ
eXLSubyNqgTNXVuTyOXajYjr0mHKx6C2HFvBp9DHTvlztLx9mCNzkh0IE9UmhUVpim5FoBx6O4Oc
AXGpT4LPK49LXodk53jhjdR9e5orKeO14FIjKGa1acZr8YXEoHT4nvXf5dJVHTQGs/4kFvd7lFny
bNWlAVyNTbsUtEWBkQfisfZPhkvNeozwwgAL4u8qljr+gMtQ5u9+bddDKe7nDZaZaoJ8gQ811WUW
lUvI8O2J9Nef03JzjwnOrt7ZXd9ElSsLZnbJe8UDZpMGDdZLfi5tzzd3/G7RD1Jx+LMx8e4l9dvl
pxc0OqmaxUqWPCHLXqmL2KmWNcpnYtj+GQ7z56cKxChau8bPc6fuD8QITSHE8nco1SW2wiESs7FN
y2ZSX94IK2NYYLQunQQEtE29l0OYxu3/9146bgNpi8vGtemaZC6EsocYPl6oOFG21MTRx+/58Zet
XWa5p20M946Wfoqj6KnnL3kYdKs9n506Idpa/YXvf76nrTTXEc367Mr0c7bpQTQFrBqkMz4rs/cZ
wAID5xDA5SjrVEtQzMb6paFTs370DkKHACucM5Ryfg9s/ddhFiYG+oJpp+oypTUOHyWH3YRD2Ne5
+chyKMduzLlHCrQcjYEEqMvfcI9EvLg94X06IuWOxxz/i/aA/ma+wWJuePctTNi+wtmV6Sg6ule9
LaYuhHHueBlJlo3tnV/5HLsoNQz4Clrikq73vC0Xw3nuDlEEUNWe7ZTkTbnFHWvSIwCiEY480cla
L47Whzif+iQxBlRgVhrHAekbVKtfxfHyrvwoAlC4PdCOBbMv/kzf3kzBh3ZT9V5Gw5RJlDBAodMT
NuDaBnVQZcUPDFnl7bE+k+A1zR0sfsenYNO5dgdBh+ztE0Cj2SEtmj2OudoCSXS3PZK58IAciSOQ
pTgnvHB/zQt/yIj/QEmguuZr/dyyB2io7M4esW2WkPdJwM/X88/f9Kjn3LIHG3tyS2axLBIkUYeh
64Ux0k9mjqFc+4zBo6iy/g/rrwBGoMrDZzpds631e1wLl1DwscGE/QHJRC3gpwSC4Vf3EtKTM58t
Srs+YR9Ll1HOLMu7iwTJpQE2bDCnkpHqwNPpoBHOA8Mq/z/ZRUuIiCfzrYM3KlMHG2k82Xx2NKLd
6x/XWnK5Miv+D4b7cOGttQtnIzkG3WZ0xNFjzt192ys7uPUbjjI0Sfd6BaVA3m2WvuETO3Vx01sv
ADwIkqC5ZXbxBMeWROFfjJwZW6yEEYiH9Pg0rcp346xCQM///hVnYSbNwVF9IrUy/9XoIRa2C3IO
VSeM++0kzVjJQ1AwJuBmKMHptlworwO0uc2WsufbrFXUleMeY+xph1P02uDyPRlBV99b5N+hKN3B
ztNntl15tK9C/lAFdysJlOdB/6sLBwSKVw92OLlSf71kD9C8pPW6nWba2X69ONxpd32TcRRQHYyH
hqxPpp7UCCryNFSizRGO1ey6j3giKYyRhoyRm7GpKhEJg9rkEh/vaOoESBSPJpLLwucuEoyEwqTJ
zzO1+O9oDaG8jLgxRhOf0GiSGP8U0unfpb+JjKrel0W3siELdQ2UPozfk42To3caITUs7dYgPtos
CIvth0SvTNaaBNvG4YUZ/8jL6HHMA8AGCk39JLeN1+Kz0bGUW1U8dVZSN3aD89X629LXhncy1o5g
RpXhaZov07EzdOZXC9cejwJV7PA2vtpDzFsqaiN+PD86ePcSZs0E6lCl5CTf2YVjPCQEcktoDl6I
96zNX0VD7fZBkNltmZNup9rdaQVlRXuY7Cjaidb5mpYhF1FqL50kieKBv7v1SHcqX1V9fRrvK09j
3En0kzPf+ej//BvxazH6zgRj6IYrI03tHXI+xZ9H14s9OReY7bj5/+HjFoZquCX6BvGsYg0qHs2l
EwrY3rJso2bSMYdnMAiA7OObzgvlQMQk0dOxtZSYP8riAwF4PXaAIg+BomUES6ncXYMOYFGsHkCK
LVC1/8xgHpx32egOKBBCpRfSwA2gTd6DbP5yj/YIAOeKD9CeqQzCFoAnpOxPvpJ9NMfdSgt5R76H
c/K3pQkgOn+UsRIE0p2OCXyDcndgGrSJRXk+iYEdy59LzCbjlX7LzwnOZyRPgkPnp0x9GWYwLdAQ
XojozZRw5+feUR1dSJlIVxUrfw7zFaX6vAb0v4LWqrqcp5qWVCFdkRhFp1xO3LHA/vxcqR/+SziR
p3VmIqKnQktmEIOKpPf4f3d6sQ1YlKEiVTbXiTLbjS4ZLbndFo5X4jY5M0XqNUEtfzsxeqP2U8Lg
pIZSxupPABwDh8ncRGElpN4kgSlayP+vVBIBr5y+x+WY5r1mJOmHsKVSA8WpZ+mdTnIs1B10LbPw
3d1ZHMge0Imnk8GnmwiISSkrM1qU6wXlzMNsVaHdLdNQyoy33sfZO3Tgd9MspQDVyUTXcdhMBI1o
Vvq0H543ilIQmF8A6gNGKP8OSykTNCigH0F1Gc/2V00ZK+imTfyf34nlCyHvFS5DcPGyIEjwxx4N
1ZAvpFLJiXZvoF8q77rOWU1Hl80SuDt61xiWP5INERRwZ71w932cmuNJWIcu/Y1i6blm+XJYjcvz
O+BpLPZdcReN+WzKHloAIC0dwlygAmTKgsHMleX5kYBA1J/dyCogAMc4FLJP0+e27XP4YJ1cqAKs
IDQ8Q+BXNKpGPPBh9UKB75TPQYmt019LslHfRPYH4C3iAkSZ5f83m+zlquMfiwwpqhQhKRKlL+xp
re6QBh4Wpo0oYc1WyR3wEwUhuxvK9KQip8RZp3nvnwJOwEBL/xsAbPIeuVSd74UC36HSn1dgSXlp
GwloNRDN+OaZ3BTAC6iqFXKnro7djQM6TytsqKXcrnPFJWdbyJ9OZh1D7c9EIcUpBedc+GrSNpk1
wM+Jvp1bUEydhb6mCtyT9D4wb6VUm3L1sASWCcgZSqeWMzFutCmiAuqzIsf88sI8+oQnlwdxaO3I
msmFEFlyTLdDAqyusci5/nU8wpGfkldB1Op8BfSETuCuT/hoCNp8hEHHSKNDNrcFr84A5q5GL/9I
XZpNdF9R9TF7FQDc6BBhDCb7vPbJXGTUgHiViIsJteewsK1IZvEL0X1p6jJkmx0wWOiz3Y6o/6lw
6CCZxeun1diFDfkhTmiz4iWjuQuWGC4rGQZFM5bYMhD2O3AxHoi13nD1lEXaozBLjwNKh399M7gE
pawv0YAGc5Aea9hiYyaefKEorW5lhz5K8beS070mbMN2YEEbjpSSG3A8Om3LzSr22vbUS0jS48EG
yL8XK4QzeXlFfjiS6XKeHE/mmf1GR3j/UHFX+iUX/MztWCHggfrnZT9jkCtn1yqckhslKbFSAnNe
nkd1VhYH6bqfPQy7faEdsdjVEsdB+DgsymG2quMn9+LOjYTcUtBXDBVfCUbOR0/S3iOU2tcvO2T9
DuxOFe4/jA9HJO2y5Xhu1BPSeWJPfZ5wQP8zT6gYEN/SweUM5ObFZTunIBM38ur8oB4EUI9HYX1B
AK1Yqx5WoRUe7GARFp4UMqvcGXtkXRJTjVjDUhOe3yJSJj1n0M8kclE9Q8DBLXlJBfy7ZfCsU5DH
jZN10s9cUcrDNxi87+s9NAWvrTGBX7HjE+6s7ljK0eSA/UbJ7qOLxIt4j9nAtXhkdU2XQmSh+HoD
X6Ezbei9r4qRVaK+KXJwKPDP+TAF1BXcO+cuOb+RvTNQe5Ukv6WiFlbZ68KR8fgrnfMvJT5fAiBm
F52noC//kYbAboBOYXyJVdLxxT0y5gtBJAvxDdnzkdW6Y/cRCFed7kGlDK4n2LBJ9zO0OuZmF3B4
IG/g2e6FpokCjj2IXHVXw8WwZ80cqjo5KI4bcm7z0K1R5Qf3T/4nIHuTncPmPRq8YQbzYbKF5PvY
PqFHxCDezR4JmFWgNVEM3hqxKh+iBDCi53XJYSYEvVNiGAo7uN1CBs3PEjqXb0mGDYD60a9+pTyN
mP0j/hAeg6KpYxYZxi6DwNfLuhkFm2biwkKZwg2UKjx1D0vidoDj6irRiQ5ajoNDBVlzhLXRdKqq
BU0Bmm1JjkpBPcs8lfhNqCQLhqQgCtXhXohsGagx1/ES+SG/2n3v660mbcX2+itPj//0NVRJlQwt
eO1EeUmbwgpEEHwbAVgcANNXziXCBkGOBvOO9nxp5gZSEaQcDX0oZarlZjigoc7o91Bph/T4uj7r
q6RlgJAnvKFVtyhULVLvMia415znL2wb6pE0xH04RfiEQaVq8/BEurmRufLZ8xzrztmMp+rAKoxY
cNbghfQWSqT3gGG9Wo6jbPO0rjSeZecty4vmQ+ULnZtdFn6GEEZjuxs0hFkDQqarxJtzZm1yn90V
r6U10LytrKkHv5QsL0H0hZ99c+lLlTx5LqX5+uA4yGaI7p5V4vd/nzSS5zwThw9KOM8MrBLdTgWh
61aUIsk99RPt80rpk9AbeRWF6WH6RjcTHZTZ0tdThnQaPrkdJ07Q1xo1pMV8rYkhw/q68PvL3a2l
f7Vvx/f7gzi6p6UT1SigXAZhCaUjFzC0ZMSmbkPAOiQoTyE2HoscjG45lBkti891NabbQAyI2Qan
diWZxBHmex5PzdEJuRtI9VwfPBXcDGxapkP6YPq69KrXqJ+8DE46xNypLZqouOYdXJHgIBCaf6Bv
OmJIoZLx65EbmC5QkXw+8nC7Sd4U769rCwdOfuUZ5fBwxua039GxW+ff+PYaSRzJzU2vxMbDJJ2+
ArVc4OgogqumXVnzbE8GKD1gFqnruUOfF46jO4xO7D86GLPmgl9GHxeS/hSPblpuIK3mfY6QciLT
YpR5sMZ0zaHNYfJBIKuJ1BLLqqE2k8pa1IKeAJ26aaqUwh2Ozjv0MiuboQVaavPVDz1YwGNEe2sO
Kq2ueIT8XvnpbofuwkOyHh+JTtSRT5GpzS3/Wn47E5wdy5kHg6OFKzqHeoasE1yWCXc/un6F7EcM
y1ZsLQ/8ahaK41KMoHQPgdmakjsoay1+NE3PNzR31ViHiior4yni1ueL9jiYEKcfcraxJFSHinA/
Ad5hM9M/N8MfEZ0RGyJdI24K2zsX6JpKRRjaKJ9/psIExUhPktmuKExsJ5ab3p/vyA6yEMrzBIL9
oEdjeM351/2LUToAlXE20GWcPrfcLJmo3vXfeJYMkhFxVDV1cy+B3v/LL8sjRNPrbK7qg9uVWv1R
/nEFozSNiJkUnW0vo0WhFmILoWdMP5OWE3/MYfBBzjkoR/a3RFJySzWbAyeYhbrg7q1eN3oZ4Gjq
2L1BWJ2qouLePy1x++M4iD62ydkW4psyJs05XFx3/1nzo8DKFfkGjinkcLerk39Ur+VSdgVRKR+3
uTXv/u/NNNVy1JtMQjEBz6TfS8nfQqg4GM2W/e7eLNwzGSVaop6/UHKwGDurxV9HwGLDvRJ4Rd8G
Qbi/uAsgIj8n1PerrVNy5o6wROWMYkM3lTpp/EKgJwehMFYJJSuIIFlc5e6YlVHxfnq9mSxMTJAU
CoN4snL9y2UJTlrq11WEUfVFNUi02B0wMiGz/KiTQFfTqwr6H710vX+IEwcdjyxI5VrJYpvHLA8u
+D3VOvOub+slgtymj6XkT0g68IRwrn6cbNVA3vjq7Sb1CnCO4imYpaqTcmWmhJufWdrGWyMtqpzv
o4Ne1EVkwG+kXE9+0aSs+SpzUfk5luSVN1QBv0sorC/AJsjATidOdS6gzyl46M/MTkF4uVajAML/
FPYLdxxDA1jvms3IYXM+derHC7AB5UIbCq5qx2Qk8nNkDdNF0PRmdBUF1jUw4249xv+dFJ50rCzQ
0UczZtxl+o67ZQ6g1nqZ+XHKnje1Zq7eP6tA2kcf4lSw0PS2HkygPkbK+4xr5psda5fcyrFMibBR
j4qNSUlT6ppWnOgwzAUi8qwQP5WXYB3FNj5tn0N+z4kiSw5iseqWd5MoNCLLe0Rij2GYFBdZXBCY
3qnzUzEh6PItHQrfWlAYybJiXUrhqSyK09AFLg53lht43phHQ8TpoYZVBEdncTMflGO1/FpEwOdU
vnZqIUs9EFheXPZmRcNfn6oyDUnmug5IkAWfg8AZLn1SbVNJc5FglWxb7s99mdjIr9oF2ooyy/pY
OBLc1lJBYW6dv4BzrHmjZtEJmoboCGhcTGO1i7ZhokvsUcF9130obnqCGfrp2qq2ut25jSHTcGzw
r4BCJtnDbNpFICOIzKG8guh3TGxyDlM25m4cYIKGelX0W/gjKlZILfhBdRdMRod5m3jWPDQBz0Pm
MkS6QGOjKFXSSyNuZCRMgPabrJJYtRWwCk0PNtl22VZosBxWp91FGKCQD3DY2u/bDj9GEA6+5fOE
gnwWeqy+9jhY1JuIw19iyvFgxasFoPweah6lZQXTvz1CcEx6hv82fnzkuILUqVgVQRevS6/XL0bR
Qm9cCGnSmvMX19U9NqgZpykNwJy0CjY9Ai/y6tRph70HQ4kkQ0mgC6zNZN9adVc0TXmHVqbU1wig
cqMrvDn7ZHLpF/UwDBfdsoYo1Gc6RwGtT2xhFhqNthJwsXzgiBUywJCEjal9LX+9wyUnvNoBW0RH
nF3fUGEEer8Wp5mnvHVqPPwKJuPIQdyUeaTKI8NIhS2fcVsDOWSPtaXQMWZEmjA6zosKtJ3NZjzf
U8dfU1bJrarzaRWUewwaEcJHQ7imLnmNA+m59WV6LccjZyQn9cBFevCTPE0bI80hAMcAjuTHZNmm
pxAt1R6O7Jz0fqobAZNIiHo8Z5Qvqk/Vn0713lVjpr4X6nK9oyuhCqdMugXQRkPCqi9MLRndtz0d
RX78AZHZ8R8eY7RMMJ9omZXHRAXIkgN3m7Rsk1j8+EZUcXYGX9JSMFn/CFeLvkEzUFsxOBaciC1Z
ir4wP+KMQDJzCjbFnt6joYZ+IDkdxi3ozutULe+BZ8nLUmohNB32CGWhq/3SABT5AwIW9o2qSE5a
XApRA+D3g3G/vZbYbyhzhm7VrlWNj5VcQ+IE/5qwZ3HqU306u0+YQ6MpUYLpqlC1AOl+BD4t48jW
K1xlu4/L+c/YmNfQUq/CegG0JGEdqCr9t+LDijeB+G695Nxc3ZsTjQpsMTsNc2J/gfq3NsiLznck
ffjsJXGBbo6xetjaXlB5POjp3Xn0MH4kHW08/4pYUhV9m9gB9N2k/m+3VrJXm/Mvtpygfolhd+S9
Of+LkJvHTLg9eUYCVwH2eKdsseJjcp4yEPcucR8jPXlZ1diY6F478PX9IZvd5GN4mKC/DfTEBASW
L+k8nQNJihou7aNP0f2LEI+DElSYFFePDiQZ4ig2+oc1MvI1kjcHJ5hKp3f5Iy3+XOBx5/o3YTb8
kmJGOhtGMDvreyvFfJMYREcM/zKzaRUCPd9fASssCGEgbZ9broGkrbc4/LyVgJTIkYdCmowIf7SR
zOFTyGSVQC5k1V1X9ATNae/Tf5xBkOKRNUJgVF8rw9NbPmettvPfqpvle9VI71uZs1MZn+NYaw11
POzmZftunS4OCFJ26+Nrjk1cbsyzZcd6RuPThKY3WJYfEX8M/9uekpxuK6LHaVwzdXZEtDfdoi4F
WlPot2hiqY4rE3jtDwfVOwdTFy6d3UkfjicCoB0WUDd4n98BzG3gwG8UzlB9XkJtO74EyKcgy2AG
vrEOZhz7wzWUs0CtHsdR9o0Um/yJgx3vQxFjE031UiDGF3dbI5Sir83IvHPMXyvOVTICBULhGbmh
9GkJQJzlHPwBrPOkzQUysCmOQiH44qrJg6qHEeUiD9ghGy0io2jhT8uYfYxvLhhw1/orn490zp04
pBgIlZBgmttSOWHMAJ9NOcr45fKP5uflTlx9YeJssIVi3KJ9aiDDXXzv3tUsdz9b6JNdTbzGxnpd
9Osu8oUr1W0pqzmoDHkuvVaiqXEPuAvOYYLBQZnG1ynQ5v7YkEzrWJXDGra5pnCgi9UXlBl+cHvD
eqHLVcCFZA/3obyaEN0K550aitnVOMMe7hSVP42LmcJ/rAjYrnSpsjAw2Bk4DdumGBsCMM1idFEZ
R2lGnA4ErDR/247CabgZ8N9i4y7zCHiVoVIlcnMXxrwIynKEnX7C4vdQw2q/EhrxFeqKP054TB2G
mZW3HngQ+iXKar3Z8LHlUwwZLAOLz2VverHrd+ByTlfgxGvo27LwNsbm/sr0ucbWY7yEC55Lyr6f
1M5E4sJVMiBb6zqCiBKPE6i7bT/I3ZmmVkIgawcR2SQEW3J6RYx4EuMQgKpJRSur/1NPylpHI6Ia
iRaak9zDP5wx6JJFxWiEwWdDE3G8PAQ17F/6PmbOrVArh5ORfpQhPJ3pC05I6mhUy6HM1652dtge
kFdYcLdqemixIVNXrJv+ZcnFUlFPdsfgqfSPIWGZz0LYkvIzdvhxoOJEz0s41pnFaMSdgdfYDgS/
jcORC7J/brPzqQ12Ma6aioY6tNgqi+Cupd/Adfcksjkb/IhnZ77jBFW6+VhjFoCnfAiYtQB8l2Mh
nySJDFRK0MC6BM31ILdZ3tAfLMtf5YBMTlXoyG4mHJEx7LH4yRg2+hF3JDSKa1UBAmVMA1tUyQG1
uKvPNWg4yOqAD8PGZJJMTgQNUkrE9l/1xYPml/5Z8EL4sRjroKwum8kS/dW03+G/p/uhhXo/LByP
n/LKglfl4fxcmEN/sRB2nVPZkAeIqSd4/vxlO/+OflDP5ewk9HtiKpGmWt66zrbYo/DtxOeNN3TR
t/iIX6Wu1yNn/0ykSyE+34AtaAk2Uan81S7PkHgvVHhzwsg+emiVhJYs4AnI2JGnh0H7gC5HchHs
x5BJVTjuiQsqj9unhiNiFvENvGyJf6wFqyKY69P/fCvzVKARCSW5tNp3e4w3O+0f2YZZ1NJ128Tr
lvwHNr40X1J9wqYLP4z/Ru9ZB/2J3ilhV7a2GTnvWkhNyj7p33j3PRC5/JHzpU7gMZ+FehgwrglC
YsvAfhCvmCD8qyikKWKbRgq1d+p3rWmC14tV2Vz+rll5OCovACA8WZrJLcxoDpSOrRK/dSqpOLid
jdhG6KdTiz3Lvoff3qfc4az/FhLtMuq2opNq9k54RSrwY+9mlRzvsC42QNEbSHyeolcVBmjVL8Yq
o6Hgxx+qgSuvzXkQGTWEcL+nHYztXYq9pgfOrtLswGAkAFqKjUdV2UjjLPpURwRr1urilG7AvlD3
90oFX3UImF4DjsoFcSglt8+CDlHsOMIlCl2EOiCRDJNjYz8ceQrUmg3SWR3ngiXHhW4ParIkaMUn
CB4LbUr/rpSClvd+VEaH1tsQdlcpehcWkOARPjjK3G8ipbHZCcNxO7VMFVtuHOrFMOXZDwEGYY90
6Hg+u8uZxQUCmGLZe2egpSgmtrEJVFVQtX2fwo1MDbRIXmogHMMGQl8VNdi1lsPDBaDbFGGUvzqp
e7AGHSJrx8ruPw1Jal74vjae9mnY48upE0/6SxWjzt1SeXTljfVXrkB1etI+eXdOzXqwOcE5SIVE
4lega+yS8SdKzLXi2iGjoIDy7WCe1Xl0A3SoQ/q5GM9/7ZU7pxivOmCIij1XQJj4bOMSidjOrT+K
NOO/pNEX/+33hdqUorew9jY18KrFm6BYnsj2RYiYjUg4JA4I4ygwn9T1b+x08lwRTlfieZrGBNMd
o5jh6KcTrT+OrchiT2fgdiOhD8p4iXvQXDbbLurV9RQtZ6KtnofIfHyDNvcx8icuxTYXNFC0k3IO
VOd6448QPv9W6ziQGeM8zHCGZu1BQf/iWAbBq/wEVAfDxoQEmQGg5o2w8ZavYomEhXr6MKWgwt1I
uzA5lOX/xw7o7tkk5X/gKoIAND3ScN7XldTdipkzsTFKMWiaohl47AZ+hxoGWj0vs+iQKddFNZjM
qb8lMu85cm5yt/1R/bfs0oP+EAVrUdb2LOms6fXaMO5MmdoqBMUgkvV5J7mfJ1L7hDQeCDTPlP6c
qP6rZ8yTEev3qmDiCu6lpUvbAVeGwV7fiS+9TuuvdhcI9qrVSy/V56l6ZaIfDfTozgCwsIbekw7T
VY8Gb9J4+/1+Rm4b2t94rzKrnlwSvasIXLbjBBvPkD5K2MdSaE/yc2MBkuuqZmvcrAPr0rf1Kg5w
9Id6guTfoQyDXRmLBoX8kItZEK2iLBOO6iWOyt1fMVxnPeOPVD8JkR+bJefYIchyZXp2KUSMtdl6
hY+o/3ynN4etYUKmU3Wg/1/OKa10TCczLDkZ26RbXruFQ+pAjdp5++FN0uE+HKXULZFAXLh1iC8J
rA5fWn4gF3g00R55heZgfQNLHbyFVZP9UkRRPWhuqeDhMzS1wkAtureq4/Qlggdj+AQvfBzqGgen
337x2IXEpz3lHMmEt20ZKh2ozLA3T5RREARr3ByKkHZOBmsQN1KDwneWgvCbwuXEjkz4KCp4WV5x
ceJpf6POazj+w5Pkczgfh1r1DdDpKrM8NRpGZ2dZIMxnvyZRI7mIis8IwuSoCkqY2CIOMR/sijIJ
UNY5kDdLIiJBkD4rjHIp50DUcOzQyfAS5j2B4MvaT0X3xrY0STZZA3UqOR3meaPw1ul5RsqazxdV
MsuD7kbPv2cdvI3VeepSXeRmbAbhaXLrJJbqqWvNmaXSzVRs0PVSgp/YUw4dRblRD7xEisRQ//Cp
bjjE2T2cyYuUDtZBh7zvuDdodAkINyUXwkjI3UfdDUvlOYxwc4muSKX0R9SGNtGCp/IYW9DELp29
Ed7xnGEgkLmVOBPrBZ5EHyU/0SabfkJxGpG84UER2GJdgorihqEAdy5Kg0T7lNO6bakegTfF1MHM
geyK5FL8spC3ev2y2v2QpOlZDbP9xVrOv8PvAC9pOSD3REU/MN6L8Lx5UDLPri+3Rg9meqkjIHTD
PCop2T5RsJ4u5mSBS3wdC7apxuMZXJAveMBKs9CRE/fGNhhS84avBU4z7t0rcuqcLz/LLMeIJTBD
Qoy9hAHfXVvI8gVjOWhV8sPTMfurLXwA3rXX4AhfBoN/eKn4fFak/TzCt/cOpCaxk+wo+agVtTj1
A21Uf6iJu2Xnccz2d87aPLyaoYHZdJOUVIxI3bP26qpPFJyczrTT7WBi0gbAvIqvT+h2dSbxMFj7
P5AaqjNC3tOUE33EoCf8BKfBVqw9Lk3BbppD80ahKB6r6SlbkguUra2QUPDMlAywfQt5ebz2+i9c
yL92+5dpPbt2PE+Dk7SxAcssOUP6PlBRSssVeSrDEAjeicDg8Teywt8xMwPoOES5TptuXVLy9SHh
8Rt4HZYjKoeBqADpgELfuH2ytdjFhmZk4TaeWYKv1bF1RagYXlJ/CFX3RDqIWIto6iNDtpBfr4Kk
ttVankyJeOsOfp+7AX3JgYbD0nMkEB+cyX42Skhxtz06L5PrkZ+WxUbfz0/eOlBYKAGDT0wAWqWO
e/D2WSe/HsMStqv8z9PnVyk+TWcaOMb/musYReZoT3D5WHPhjakcwBcsVN/fK+VMl7kiAixx5o8b
nJd7i/eTodsTeNlUL7opOXwTiJ1iY9xgtDDHoF9KOmYLGubYJ15tyU+emv3vEXtvFmx/0HoAIGqC
oK5IMa82BBGYfgNamRwBOKyOq1t+OpPW1cwQvPNIfKlNQAUu2NIldebEBkc/+qcaxFiPcd53km4h
6SJqk6iLJ9Q224ZFBOwILKM5b5odl2BLbrjhNBf/vJGEeBc1WSqM6lQ6ibVvrpuDcplGL60OAiFD
DNzK9NMcFbSgL8ewDwEsQCIveA01kylIlxOKAr/NqNc1VJYefC2qxhsR9DPXuADM6azmNfVhBggn
RWC6ym843S2ZbnYeOlUt0nJtrJlLkig6L+2O/ODIjFudMq6JVc+nlOw9iHXzJuyLUjVz2PT6MGzT
GXwESYmsz5ugSpL90XRxof/6QOaIju1Ero0ttkCYN5qJ6N0CxMfv8rLsFfcz+WvXzNn2HKLCtyTi
0ERWeXyZ1QwQF7OKvq1uk1BV5iH5QJkZdcr8u4+8XEeOk3QtHEnc9sQ/sWMwEBj3HIFFtuXVeKCl
9lsfr1/J0woXbgaWjHYy52ymlRvSFzkkU1haXUpcjnvhwzleE3jR6WcFb8D8tThED2W9ZjSTI2HJ
2ZJiP1KtEpikJxHXhoenKNkgNPBxI7D4hIcA6pmDRgeULSwq5JWozeWI7gDga9E2qGhXfDMemDZt
cqq2zo1Tlsoxj08RiTUQ0NsKDs8hgKE6wIy0SOPotiuVUVDzRcWSjlspKICKXcC0+KKIA9eBo6sr
4h+tWK3GEs7TgU/E2m5OJPiVQ0t6fveWDtCjwDgjoQxi9LLmNZOlWbB2HHBse1QPhaFphjMl73B/
OP1JfkicvThFSg1tPFF1qZRAxeQLsg/bLsEWhO6/yYNqFn6JNoQx/mYFkQdeIzMEJe0QQL8yfyPZ
D+y70WIu+uvkf4AYj6evdrs1/ET2tHuSc/rqDTHACS9SO8zmyc/5DwcUhGR2VylKtk9ttnHMr9o6
udxlva8B5LMNBzm9ZCUwEwgb/PRdpvQ62ECi2CBYK9FtH3ttdFSseuX4jaOxG4dHxi7MJPWT2O16
GYfXhF8lMZSJ6vaSIJTM2enkhC2qNXa+8NPIrWNCd9+AJzO5QxkBSKFbdzuUxC+hupi4hNHuJ4U+
Zq5y8itvVpLfE6TJlsbEDe7r3KVpSIopsMtardmf+Mj6W6xY6tIJ04n1njsV1XyaBfi/6qon+/QJ
dDM5zZn6nyHMx/7gqN+IKFyy6C23yeErvCjpIjGihKiJ+nKJ5Z5ba2r83iRsPxRymTpjgowLmwG+
JEqN77kZ2G77LneP8Y3n/zDm+5US6qY4UN/TCw/rf937vlMEcwFD/9eOTXRXl0LV7Ug+IIabFCYP
J5Om4dv03FbBZR36KkAh/Zo+R8/OCBeeL9rAdOQyQXgycorza4wWYR8bHHpW/L1qVwYd6oxGbGcZ
wjiN/SE7Yu8sXzxmtH8dew1aKKVrGSSCizQ6N54q/sW1rY3Ur/GxjE7z6Dke6RpYx1JE3YSHBngZ
bxTE8bD0MA2Uz0Z5A8YS9kvsUxY3G7+YN5xlc9JxvgL01iLDyTNifCV3UIQIuK7vUelXReS8ryp+
Aajoo9r2nIFZLbwAt0LuPanjV7deGSkm8ERq9MHM8R+g4UzWwFr/0V7hg/0zQm8MQO23tSgcc06w
ljyuTK/woQcvTFlC40fcJVhhxmJSNBfssekyTVSHObz8LIaRFECYdmoLloYRVpqEu+WB6hYkNBag
fHkHaPWNOO2/kRnUFcn4UADW/SKeVOWmugzDRrOlXEH8JBYYo2hy8agulOx9MDR+oN5+AARwkyIU
sLmKCpRqo6O6QYbTB2gUb0i4aFxt3h/5hFSUmKLKlBCBJoHwZPGROuThMgjheT4KwmkEb2NpkOcv
NfkZGN89Ya3BMvrKGwYIlWLaNK/Yo+sMo4MlcBjhGzcub49kVnXAAwFm7ZxUzYGnPG7+oXhhX5dX
3tuqQ99TA2nJmon09mISWG+mCQ+Q/ZqI5wIA4PZuhltyj2UZM6bpfQIO4G/h8ZtgNJJt8NJb2DW4
Cjnlo2crrzvZqyhIbgPAJOHz+9o5OZDPbf7rPFkgpIoI0VtzzuwFmFENNxSvBZwkIqMoMvcRB99t
mP1SwA57XOUYwifXfefB+SbVeaVyIm5H87UFX5SdLFTYo2GBiAMfzjTDMWhqnANNIOejJvqaDYO3
g44osZsc8O0TKrRfbZa5e3yznqufmkMfdw3N6zpPgmBXEXmkTUW6a6F5bDzxaNI2XrAkwPd58Gs3
NM/J4e7tV8uHzwEFfPKuglnmHXobrA77UY3VdOKG6xq0m4v1Ep8btzt4OehcxOhJg98ao51EQHwO
CP89aanhpFGIHLHSkkpEnydVYo2YbvroCSFD1e2c8iLGCw/JGw/F4R/yihCebRIabFmw54i0b7Yq
x8OYpHZfgKtRENBldB00qiKqSVQNLFzpOBNYhj/yuzGjuZqkD/lrziR5iQITtrWLD/30VpP92mNc
bh0+umhoB5wt0jvVLVSGpSyvvae7RlkuWJSwcz4Wywf+MDmeD8X0Y0mM/LqT3Vhcwo+oEJ9cmSy6
+OVeCy5+PBlRjIvhCDHS3Yw+l0J409knaSOXtpDVMrzl4yUZ3UvyJcWUFolQ05aqIg14i/TLWEoC
vhG4SULiYREWlpMNkVhXzCnxBp2gxEx/QwIm7ADSzTjc3BvYeAYgllYmD3v3AKAXnsLUM0K80Fa1
EKYQtUsQKrxUfLGIdrfScRO/Hy3BBCZT/oIE3jyUeDGkXKf3uhZoth+xCdsoumWW1AZSjLAMryWY
HpCK9zUGPPZOyZgJ7gtFBm+1Wx+ZxLWTy+JgTy9LmKANS4wgDWeSSggT9Lj2jfHR3bioJXcbjBD0
K6/GZFJa+2Z1lRsiV7uo0UHicHofV5RioJQa4A0simpaXH/AzgVPB+Q/uKEWirXLRPim+hMHWK0V
ogw4HeMLBRErFIdYqj6+OQ2/RwytRAc12W2JvfXIkV9rJCwk5wPP7PNIVFPwM2y+UrGDsMcQGtGB
0qjHEuFO+UqXT4Mz2uVZIk7PMWr+83O9t1SIO85RPMIS3fxlntAHYaIvTSBX69gZIPxIH5jWXULs
qq59trt/StPs1jcg3Qz+qCKPGZw79TkmLvDZbg5Ay1fRe9CpxzzhbAtZNt3uT2niBesnBqz+omwH
3AwBoR5ZMmOOgR7Lu2IDNvg0TNm46j6OCZWaEQhaZacoHkunU3IZVGGIScvph2nu5d+Iti/vmzDS
fBe23k3lJtJetL1PVQ+EnsZScCvpwt4JbpR5GtjTPEWNRuvdlh98NiqxM6T5EIXz2yOU04van/Za
AyRUT3GDDPbHo9o6Y61foCoG5osy/pp2voq1UpIxxl7h57uvYnbr1xV5/lzdSmfkb9OLfRrRDlps
Mu7uO4yrQyWU9fGXSIqq7j6N6KJ2fJRuzPm/enpw4l4e0Ou3d36ixhTBQtIz1sN8l+rPIdJZRXQB
uX+9PxxghIYGn+ciePH2vcBPTvAplWFpYj0WkH4ssapt011R+tFY4emGkHDKQ0VjKt6uWyohqvV0
VabUzVh9AS2lknSRri2qj0D8+DCkMxQZqxnkukUf0IynOgQ6C7fZ5HbRhkmEqPNQnGtA/WGHWNRy
xDJWkadVcXpgwV10eAtTK/yEWAsNYR26dckDrSD+6+BkSjcxUy2rYBHnfDF022JDRBq1z7H+asDO
5fWV9E/tX4JT1fgdsSLtdgFYkIJ0RV+Kp1tjv1tGNePXG8vrGNiox0VGHLSvgAlp+/pUPzAfYgWv
qlT08GgOmAVpHcP/ZzwxDCer6ufnX0OFjG7frkCbTc9KKBMSQlSjkG7bqqxAa865i2B33Mx//hUs
nlvYUCI8UbRTHODxtgNbb3aOdO/QqOZMDJnXDOCarlr52wLu2tNNUSPKf3bdLIBdtELLXCY0/9aF
c3KQZkomvTWYcMUrfVEGeFmdGaA+MGXwTHhCE2Uudm5mqiSRFKTbgkd2gqQYIRMZrBKFhJhNhrsw
gIRuD7YC+9loc+7hEh4HOQ73UcLIfoudr4n9y82n9GnwrghZjeo7AFQrnmz7PR100Ue5sZaijqva
E6b/O44gt4Xx79a58vVxSvWVlez2wz4/eCoiytlYWna6fOgtqkA2WvYFLVQtV/Q5QnYArcR/j/5U
wUuTj1LR71RNMuDaRjmSQX6vVS+YrtQMArFsCwlgaHxsmcYPR0ghgANBtngzSwcgJkxI6ksrAnEg
me7f1bb3gIiJw100cg5uZHcQWJ8qbk3HqveblGm3Ut0dUEjjxg1+cbMfP74hkR7uKeg89mFhlZdy
HbMUHnR+LnT0dScuuT9rBxB7eMi1Ari9/ZTzBgLrNPUYrtqFQPEoLVfqZTAQnhMu3WFGT2jNDGke
LI3J1hN6BbyH64uwaTiMpgSZW+JZYOV6DqFJelY82ZcuvIU+GfIhr8yileRI//phTOaJO8T8CimM
2y136Jek2PRde8BhNJhWXcRrDUA8uFWme5EQLK3IkeF2VulFkmxyX2ZkWPVZrrcSjDStOk3JSvJn
j//xA+79FmG8nH942PGGoUayfQOEWJ5ecsTQ319+aqLOub47sXXBlXWjMYy6nJCPBmPOLgsx15Vj
0b99i0XnWt6IGxVaWivsB3HDRrHE1DNKZQVlinzXnk/CqPDuDIH9Cnxgyb3m163ZjkkG5L3qYez5
Tq6hldny3qXAulFjODtW55eQssIRfPiKkD/cAieHwirUaxRnzM0KGuDp4Kv6FQYmjBaOG4KpyYmB
WKreph9u4eaz9yg8VsMPgjHl7eVjLz9JqmA9xja0YCT0JqUfpW+gLRFaICPhrQiIqtEGQYofAbOJ
YuJfo5BrVC0hIrNFhX/fBSEOKPKX7n9xwxJ40hGweAOisMmOotiQvMrhRD7tJWa3Qi7NkpmJMGuy
VBB8+ughVM4omDyjDlSKLaPlX6w7yxz2sIoECOW+0P9yri7l8uLn1ffdxtGg0DX1MfdhEm7LqbJm
rvE2sJQHmUMbuHMT2w0oh1cl1vjOeI1e1x9l9FCHVXzCRbyOUO/fHwR7QnEvdoizV9aAWgVUk2ZK
9gGBYJhudqfCa0ymTpnblXn2CIs5CdpgwoSAhSgFuP162KIADc2m69bAn3pUF0t10e0RkYmm1Kx4
WX3HcSlNreBMgyQfVCT/G0kDHTvCc5RoFn6uDuIzK6xBD5UHzgdSZUlrm/bjPuEZRD5rR4noWDTV
5Xgd0QFmFQvCYj65C7U6S1m81r8L/Ym+0UyF0WYWl2I1nvmkxBCmk7Gv8cFG3CsWuXvH4FZU7k70
oogfsv/xcBtocSDcUXh5g5s9ICqARQbUDFrwrZtZ5OvjF6/0qiXMwSK07FDlfcJig/On0KgtUtDu
JMxL0K1+h39ic+MQP+TyuOTMPuDOi166NGe3TWBF7Imn9PKfbIpxU4UFupaRXFaA4IP+EFfU1sSD
TWEx+kzZ9bav7el7CVRpS7MClx1KeTV62En2ufcIIKvNnspfBSlscff9NlfgXdD9CZMEBIaWZ0+k
Wkb1RmkHwSm8pBvivjqJ5LLedi98v9mR3JumMeLUNz3mvSX15LejgL9JWyu81/deUDIoCrBDFKUN
Nj1UHi0lwLqktabQjEZ9L9FHpjtEwwVAOuv0l3GrnrVAX9rErYfwlcYw/UQYFV+XAkV3jVscxeMH
F6BfnuN3IpIHD/T7jwP24RX1uTEZmYt8VfeIeFsIjhMrCedJphmofYnGklNTaj+RyGd78BANCTkI
mNfaP1vQSYXhvNW3bhBZfqxG8k2qQdvTgiJiEIH+PVNaTq30kPVp4CUxon9ouHWDhwj55i/bclor
Ct1d/E6aTF6zqRo4/A7GWCx9ZzB7j3Jj0RnLb0jn2huHI2va8Rz/VhwOGiz+tPCkhd/MDUGQxfwz
pHblKhqNxot5EnxZe8HAqodGFXytRkFJPZfUMDucvU0nSEeQ9yoK7X9q4BMSJRHT61YGcg3bpjkG
ZbL2zUEPLJ0wTzd0SGXlzTGfy5JLo10Ai6gZcHu62z6ylI+/bB44NRSLYg7B0YbcH6EcUY5tN5jv
99fc+R/i9WsWdORRnoT3c8TfdA57mliasxV7jVRO3wLzmhv9MFb02XynMT3HzHa1loqxxJTlbREM
JBOCI/cRhIOxvKotDtn8ol6YSjRLpygsN1fIzA6c1WR/P/iYhruUj4UWerSnnabdytWVidd9VetT
lsE43Az4PMo+QnEEFyiVnvgTHI2Jf9iNtA8uzkKWZN+PUOSn6HvNHMpge2Ebru1bV4cweVi+KV9S
x4jUWDi9y+2ojUigx5PFHkPum22cYkNcbIrZ3cEOUZUC6JAoLuvyESaPDV+NpwG+2wNiKrXvzkXL
0PVmfBXJB90vaawhJGXA9zBlDvepGXM0W32s5fLCh8KdcaGle5pxofUKlo7Tqsbf5NOAxgwGe1Xy
fQo9rIISrbiuKlVd5daEVAIscc7ifrQldwY32Aw92cmWMy//FcuOrikTOVL84IMf417n87IraFvv
4Yv4kGnixPHt8ySMQiC81BmcQm1gs5CNNgbrsgbjMBbnxXe+rsE7f8X5wSOHBifdyDTrbDYQ4POF
Xq+miVoOMjdO0rexzxaxNpoURnuVivI4vppbK3xIznM+lfToWvm6ICjL4KNMsFlH+WhP7B95lGdn
J1kJEnzGJAYp6kLTzbJh+5b9VuzC69hGEwVXTWInG2w+JFkj4aoNEpmxASmmHoDAmejFg0eKy057
JEZD3+Su6nMDz0rLFeYqOcrqTSvRQcamWBtigbF/4Ohm8WdLNc2qo8rT3iETq0SwT6iMN9IFhcCa
2XvoqvAXki506mp0fB66GtXgZ9QUmIvbA1r+XW2Iyhnu61LNYY59JcxXBUcdqFwXfQA692QhSunT
15JcLjHXNnqHyk1TM2cUSiBzN4whIl0bBncQZrtS4ll3ufQx1MwmEi+8mUPtpAd1QiuSn+Eehh/1
LBw5vMbXGXFr5cayfm9JtcXd5vyOGexOAD9llXFmlPAn+cK8tgMELJvIi9KDJg8Z9bjmIsYm/9HQ
pXoiRihrgvQIAsKsNthVbDiHU+6DIk/+0F50dBS+HyFraEW+nqXFW8zhzfhVFgw7Kds53ET+H8xH
diH3UkrtRqzPABd4IK02VlcdOhV/6pG0tAhsrbxJvPotdPT1K/pwtDF1N34fwmNLU2/enXv+7xI2
XMNd7GLpzooOLrPascIOApjAq/AYadMtts36ejcg8sJt669i3F1UYzfgp6Z9UzVmGlCaxdh8QTop
T5qOoefLymGy+/8d1kQCz7AlxcX+UPRWK7GRqrecvwbij25JlgCHbldrMJEGe1wrQZc9wjWPb4oO
3NvKi67EPA/9XNWLUncQ6/ypuv82jwn0aVmjuCDHAoyug3/Ce5hj5z1hTh/M/O3YmRFEwDNj/gjc
Wds9MIGWrlDl/xSKa7Bn36Y2yHzwppHZ9S0Pig3ivsU5VrAYvKGxRhUEnvMNuN2Gq4OA/zZkhwzi
5+gKtmskRrWCD9LLALL3Vg6bRHmQ55mg4OhGg+yIftrGwC0peHksEmp+qUU9hE/QaLD5N8A4eKci
iFeen+QrEbJjomE4Cq58G3MoSqFMXvpm5MKUK9qPoys+fzoGfwXIlVvh0aHJfqRHBu58LVfD+9CN
r416aSiNxY+KFb3j8QAC/yjErBjYIO2WEOMjkyDeN4GlU/6PpTAnsSMvqJa2iqi4qpxk0MH+3ZEX
Bfk/G9ExumNT4O5rxEj7ThqTZqkI4SbiwxD2aPTSBofSlyfQGZ4Ads6ecmBwGDnNdox/noQyhBUM
/nZZAv8SkiMlApS0wlADeu0Jt8CGbJQ0aUSaf/o/9a8wAehkwWNJxaCiGE/5j+4d2F9DCrJ26SJ6
pTRVQJcy6B4hf0udCYPjXrwumr2PCJIZeMJMsML9EseBJ5uvk9K0sTxXxouSh8risfpmRPfPSJqX
RW3gdg8voTCI3UROeaMOnbD0vK8QT/Oqi+CElVrFkuCZuDLcrnQ6g/ZGhH0PpKqIgOEJBAIbHgBL
dPABCV4m0dVDf2yIurl9B0FPT4QRZ6unx3QDQs169rZJq0J9HFslKzHPB4lOo58c5OFctMl24ePo
tcV9fXNmeK1yFh7MzOSb2GcVExZx8Zifb4fYtk/Gu4FevA8t77YSVnhUKZyqX7k7Z8gvP/9Q1HGY
S7gxm177iCYM96XxLVbriviViiN5Vv2FbOJNG96jI1KDy4xMSe03pvRcqdtfD2zdidXlgknPG5JS
0DmHq6BnwPOkWYV3K3beZyKPdsu2G/p1vF5kmUM2VvH/Fq70mVOLaojnDxkzB94u48oHZZqze1U5
cXp8BDNLbMSs7/cCm0EzNz2zaZ+HlUpyZIoFj6OGiBPLXPGP0G7+FK++9pJ1tew13dUacefS7g7E
QblHrSB4Rz1ZpW/SEw/R49bs4QhxxsV1pz+CVn3WWzot6tu/ff6FkoJK+d7/lmcmCbHELpIPbvRO
CTStbia/BsC2WUPTX5jPUCsGlarKs99d6mIhqZr/mjUY+wT7xeHpIKGpNpu1l7twb0WXt0JQq4iJ
sEOW5OosxUKOOHtbS8otWyF2EO7477vpiUK2rJitLcnQc9EcL55Cp1DJbT5bE5CtPl6jYiRJkTL/
pmKjSc3F1XqCnZ/P/4/NWsf70mgsIOt+3/gPdmheqXVv6XBSD3ws3yNpVhb+DTgouDW3oHYA0A7d
PfHqoxW1NLWhFaZOJP8IDgyjdbnW7JfI3KPeBEr9HyzCAhmvO3zBVMlPMLMMOx+JtXKsHnHOw1Bd
SJfLky+Q3g8Y1v0ElSzoxGtgp8LV4NKonlRJ2IU42dc0Xj1+lRAlSJoomRc+g97EIq9Bqg0Cbem3
9w5HgvTcjWVUmSV/KTG6Bdr5wVl/64LE73m/3i58J31t2HdPXatQnEgwmHqn39SFhXaCuUm2X9u1
L8VW+mcjQWP7yixUUPezI9iy3PQoLj+6OInC7Ds5+x7WEfKMi/4/ZlzQTWLqTLF2Mqr2ynrQEMl5
LSG2blbHgc8zo2I6B0SGBhdFRJrkyMym1VZs8AcatHGzbk3I/sJ6hHw0S1EDXaZtzu/4RjPOwBnh
aa+TMXFdtu18goMH1C/lLBsYd787K89+Dkfe7iZFxgXc3360xVfJEcOwOWN9bKhvNaOiQH19TGGw
N6UvB2GBo/HB4h/tfs7ErpVEmnhFOgwBQyNQ5btLPLKKfyZXm01nl2KqF7dchNeTF6qGZjfAs1ut
NFgaWSYKqqND3eC7nzY4DrxWLkHYIDZmCz52TZVOSzsR7xwoe9jZkubIzVYu1lsokAg7ywpBQ/5g
hHz3N5VCGsMMC11TLG6V0ZoegFamggEJ8d5hBfLeGstIx8xkmBHF7ZAliDP3KV0t8uUJ0ytKgR34
AjI+LAQ8BXSBygLLSAM9wd/bAGMhFPRaJtZSIUHzYBmQxGPF5RNmtJumFYZ/sxJFYQGSgeWf6A/k
NlUyBJNO1TAY05A2w/RteM1R1/cSQucXmyH/sNP1k4qBqhQ8ETPxwShSHnRGtbq9QNeq7HYt2ZfC
vZ7GZgOEa71P+T2Mcj4Be5lLZP8XMxhNJZ69qx7lkgO9bRRWBJF+398qTqif7BoQ4sUOATgl39VJ
GAxS4HGD2xeAldLVqYsLLhT+aF5LTz+QjixYkEWr6AOEhsJkaHGSx5r9CNknj1yY0zu+bVVqS53A
QBpogYXmvfKak0KM0NmgjbgBK+57onIhYgZ+Q/nJVWUNZMCOgH3uTwvCV39r95vWloSpC6QTWjBg
vPKLkL5dhs0GNwEgMbMdLz6o1JZuk7tPoUcLwyGTOz+CctJSXsFKbLpf8QGU13+7eY4+b/Kdj356
oKhzqwXVlKj8kPqx7JL/l5rbsQDO71NCC6q/1MotiEiMpamhVi8Do0aemXbZ7JpCPkopvrJQ2+qa
37EXJBbEzDzbkcVz0OjiqwnnZITaR8h/5TtraycisnUp5QEJjFxRhlTswy8hBoMyyw4+nl11/iZU
APDUM1k8RiVavMCq6nRd2QT7bwuDZi7bCoN6ZlxWDyby9hrc+hKFBhTBqu7OO7ZZG6xA0PhrxmCr
f5KfKOiEZfZepBWdgeFGyORWi25Y6aHG+X0k8x+EPs9B73Lpv2TTn7zpsgwA9AWJt+DxXZRdv9cJ
DxGqXkx7nZPDYkynmPje/YJmKp/HY16wOyXaP5TdSDlDwmDeUQ6PKrVTKul7wxAqlKnmiRHW/Fi1
v9KeiGmFTBxG/N4oaWVHO6mrN7V6X2jNpo45yfiEzTGydSbXR6yEBr439OdkHbea9gWwm7EiY/aS
nhA747EzEL1rlauPs5Q/3rTG6qt6VojSXhPaqjVBtf3WfiBt6unyQ8VAW8DVdrr4zp7r/f9aYF8p
8DtU9cGSLxaFwleGPZs7ZBz5P4L/HtdYV/qoUPyMPifvlSaIBRXeNnN8O2EcTX3N5a6TFOt9Sv9Z
t7RrpvTBXmxlpDdWSh5eTqHryuf/+bC/58ud9Pf/dhyoOWbHO/2+KN3lCNSh4yKzXY5rAyd6Qwsy
iw7smGFcXb8smVG/Sc5/OhAaeHnhkGI0CkKCCSK7NP9zgiPxYiKevWuJLfg7lkl7+9f8HnxLbVS1
oVLz/N4if4XCNYRdciamwBalIIZD0CyrBbkGun2dp7KfuObCa/fzCyZUVN15f5im+zcd4d5n62Z3
fCGIekrS6sm85cQgN71YTdHRAEcTl6yBgpmP2TkRT3bRF5DyYYgC1Qkhx0r4icR3thp+Zlk8oJuh
ZfblT1phqyBxyceg+fpEVpRQDTI+8iI2IjIWuPX4+Yfw9kYtXMR8Jlmyo2wDLTWXGJ1sh0cOJMEQ
HkaqavZ5GJAlg8VK5NTLkQEGMVCjnbiN97lWficuPnzxmiHX/9FfF+HGuX1Kk/6yYt6e2NL/0Bde
2inkWBaySAarvuVv1o2scNFA2Y5Vveas3vd+KoCbQPB3M6zQxsEplmLe/EWpQlEmLHd5bsWNpMAp
EeELzqN52k8x37BnmQ4SJQ8soL/glhoKc/AzEnwwUQHGGtp8I0lMkMiJcFhq9oqANyUC22Y3gtZA
d8AmrXt+ymymauDVz3ir0sjkVopCKkkH997hZvjAeQeXHWasmPP7VZulJPFlw/cPWl2N8OB1YzEz
yvRiBpAmgSYGKMLYZxCw92QiPIJcRCCHZA0juBwCFWbT0ShxSDqM7ArFSwLr+OmUYB+vgH8yUhlD
JHr3qG242CsDtbhCHGtv79b/Wc+6d/e6T4DRo9a/9a1jCss0Q4anrFdkNAV3T4So0Ngg78SxkKLi
Qur6P4qqoWcHrA1yzEs+BsYKdxgeGsy2214I8gud3tlE3dYXm4xChTYOJpPCp6lD4SscwJYarVpp
mDJkS0Ls+OxkphSc0+mvC/90RH1OhSkrh48PzNXwJO6PS5mlr6upEwA5n5Act9MK0Vb8Z3+hwOss
cYF7UbSHb17XPQl6Tsh62ppUBV+r5Ji2M4DOHI8lkLxDDWv/oMn0Ur8RgltqglVdZ6Y5mVl5OC3+
lW+rs3jWNPQbFfgcl4m074ERPu2ShjVnGmub+BncBt5ODSEkuV6Sk5zDvElwYS+dv8ZR+e3kMXsq
oVmJnKnvEPTNf7/Kl7uaM33NdTYRdCIFTpbW3Uy+ujEhkf6umv/z4ryyXqJtwoo86xhqH4mdnNYW
EsrdLyGhO+uPVn69t5OlKYTRUwXmkHYJCxQsho8JbbmBA4AL90MUVgFC6MEAZicUfoLOahWcNAW2
Zi0VrDMyF/6qqDJ+VGsByBhJISGaHT0esXFugonfZOChFcBrbsJ8FBtN5UdJpyEBjcAl1QC150Ax
0XuuWcOBug9ZVrwqY6TYhVmNRln9SK+GhIe1n4K5/34QaLsXX1IpIuL6BwLfqR5m0MFQFeSmehGn
f8k5XpFz6cHmrDDTMl40ZHPr+NjdOdH+YZ18dMSdpf2u21zAHlFzUU8fbruokf/fQROHjpC3d1f2
r+IQ6tNZs4qYVj7wqFsOgRZatquKdW+xnhGZOcynh2NRVKinf9Krhq5BKGwdbRAfDp4LqtIFhxIj
OmcqQSxOYJN+K+ACeCXjip+dMbGAkwnp2xSml65ngKNJZzx9MZEHHFRVejTGrf5YUoebdDiGc6Z8
5Gs2tsOcMj9fb8EkLX7JSfOLbm1Ez/Kz1T6snQ6V41Z48JGVzOBseGBKIgqruuPhxOou9BdHQz51
c/XjA8jwokqeLdE7ZG7p0yeDitnVZk2KhDH50zm4r0Ij+gGRFNJ1/BZwTJGbp5L77QmyOUCoq2qo
Dc2ZZWWBmeXfrpfDNo/yhi+GpHxqpakeEg9m2OQStD2wSDOQ3uBrmxy9MIXMf0TTsNQRugPBhKTv
1RmBYo/zIlgcpDQmdiYwLCzWDbvK+shdQYR0p7Fiqefg1ongpTyRKIAGFtlfm+fvRbjfDegu7oGj
kUWfJUXzffhQmyJyuRZaTlGjBM+2lzb9EFnESmIIOGIEJapJe+/dA6GvyFogaO3fKyAP/SFFXlZe
vAdZvQdNYaejbdlOOUEooei9WiyJGwtOTiiBkddrq0ZLHVuCnVHE/CHyNyA2E5iHCO5iKoCzg4jR
5eUIeWNuplgiJVkWfZD7koWQV6G1fBrZH93P5oYh2TbKNhVWHCWjJuGdS1KjIwQOYtMJ3TmT1/9q
GzRO0tg1wuMTIgQ6+7O2pVS3As58JHvHRXcp10b6Pz5udFQrZYUd7OAywQqJDrJ7Vo9fZ9EVNoZ6
9Q0DAFnowQG8ljiAS+kBl71eIKyVP145VaJR1FXxDpjjreQVfz+CkW+XrnxkRR+CDMavdPpsHcBk
FLVbJH5mCkGGRb4Ho8giXC/E53A+VAzyUmKavGsGsQOHRF5hUhubXwDkgNJlHFmIlh8lIW2hdRQ/
EhqEy8eh1nIxDHmCx3H2rU+5rYAmzpF2YzF97cG6FOvi8LlTiNfyTGwk2e/OnO2VYTBFx1h/rlRU
GSGEpXQ2Ov/ht+sRhHxXIt1y7TuT1/bYblUn1lylb3IvqMzQ2Qb3ryh/SKlMR0ylEPCIeiVElR7M
+d0Oyg1/4c/J1UNNQbIOV0vuAssWjqhTpAOSg/KJfxmfoItPisoNZqnHC1/wFEb9+eF4za15jcHu
3zXezbqv1FEZvyEK2KfXxsysJMYKYLAh2G/YayI3KJfDjpzeg8kBX+7sYE3EPDrhw0/Y0jxZig0I
e3UOiPexKtEWJHz+kmjoGcWcszyXYcwJaSfWJfqpCyPFmzl4ALZ/4JtcLOUobnq1Mm4bXCa3KVlJ
lh9RISfQMFOm1Xl0Mnb05/V6PXxGZtllYtucYe7G31ORYdH+ClHldSnwXz4rFXhYGXk152bymMqS
6hBnmD3iM91BLJBV+AMRMATELrzlOqpekY2JvLgWKuCw9JhmdOQyQ8KkZGgNtCbKafZXP51k//E1
Ge8PoDI6atUvtzUCisMNZRE7GuLlRAmHBAkxuhjD1xkdX/Q7vgg/t77ilDmQCWyWzBHUG3Rkf3d1
k1guAtdBMgspiQ+XrgtbBMCsVBoJcJxlGhChS9xbT2zyM2rPvkehdgRCpU3Wj2M4eAJtlMUZzjTQ
NhMqLv7gcVtTafha23mpp2yeOsccnQyjXIgjRmkL6abVqi1cDskNBxqv9mjxy7Q0SVqKHENQGTsC
Uu8uc1aIGxqAUtx729FV2TVCx4QuQGyGiZrfosSjGQCMQV7jAJtPh29J4JVeoRMYG755ePCutzPD
l0IXD3kQ17LZz2v7ctaW8I+TWKkyj/PsXtrnWJL+YkQjJpuFCLWqxO/GJBBWC+eGS3j29J3dLDwa
H+yFxGW3DJBTa5VBFhfwsXUtwadaIycxlXgjrVACMM5y4MNuL9avSsd9FeYIbYkXXm9sjvtoi+UN
owy/ZPidPqIk03Qn0x2IOt3rRBcn16Yda8oq9V7t4bZ9UckPtdzZAVKmEgVjd99AtQQw8PeDsa2v
8aRjAgpukCnzQ+cTnMRsGF6X0ggGBksk5rf7kXv/3mV6KdnpZmul3B2lyOrTREIgyrM44HqwA910
iY7hyeEiJgKvPVRmm+dXc/bMywju5uhabDBVDYkPFaBhOX9S1SJKAvv52Kh9evvPI/Tv6UjGedZU
5CvlWlu+bdTdrcq+ZIEGMMe3L/+NqFx3t3Cvhc0vBG5gm4HdRiKKq+Jr2OM+CqRqlxL8tD9Mge2/
5aTxKXlRLKBdGGIBXtG0NcXZBQGgIFeSQURpqrCTPzm+3T3/Yh3bBvem2b25QDK/EZA1+FsIQXwD
D9AVNdcZbMJySKcDyiJRJosP12DWHBs1UolK5CmfmvfG3Hg/1tDoVYKshVMDV+7Wzpb0JPXq8O6G
rNEEwnMBeABkWopD7QJ0THrG56QxD2t5wflbaFY49gK4gzTEHjgj2It7VaionOoa6VY+89Bo7puU
OIdCTcn2BgKmBTLCPYzqAvxu3OeOzGDUt+ntffX2YH9O1+99S1lqdQVTtqzHPIlhKbuxPwv3vNGu
VcizwRmBLph3X+WPIvPjtqhpmZ+AJR5yBDehhAidFf/xwkDQXWXwn1dUQeJ2TQVHxDvrHhv+kAsq
TFEArUNHa91QxLlkyxkZzTnR5HPnrqEs3CQQbC2u4oWvetLbh4tEht70NTLtW5Dqx4/Q6UAplaRf
JNw9Celxk10CXg2nHZrhoXbnu5MDoG5v9a5PcW8ebq5DnWWO+Me0UewbizTZJxBqVxQhId4Er/tv
Qo0JumEdydkqO1fcb/9bxASSLbcxwmjtP7KgeZUcLr25nGzYQNiLnhYpjSc2D/hR0WeWlfPZtaeU
qxanfwEyvPT85Etmfk95ctnEOCvOOk13FMabTocnpVML1fRocavUN3CMME2RBQ4qS6yf1SFdo2NC
LZVJbtAk5gCs6s/rK57jhZSvvphPh+zUAtQGlkyTJ2wIfaLJApp2203T++gKaJmnG/xXexXFoQzP
zgv8E6fWPiebv3uEtRvXZKpWplFxF++ziMLRPL5DpQd6ii2xL7xLA0y6P2VBz1RhFZgAd783yhVo
WR+FPt4bj6cTpUzVsOhbcr9PWJGCxxNTYx/vgczT6Ew8V1ZETmUnFbbhTL25DJIPLuqHNsGzAxsz
115e1QYXGkAi9yXKcWlb0OqSyvpyT761EgpUgk77ZtOIJ7qchSS7u1TR+g6H1oKdYEXzD7i5OYGK
XAQ7Ycr1GEBzLyaJQ9CAYLdSsIk4RvVIAqRich3y+jQiBq81Oeji1beIVTc3wqKBVQRJp+qgX9mY
rk8cvDGf4NJc3QpI3P2LXZxEOAn8/Ld5ycOT6/N8k+13snWzaRdwBsJsf4dWauKsirqkI2SI6rBr
ySMdJIw5dGinaAjSHFyHat88hJrQIDbuVRRYiOMK49OZErDfLsZaNHWeqnjI2TCTTliwOilxai2j
2u4bGCbE2pmnCAu3Sfi6ivOzIEsTWZhj32txSthA8aVzxLqu3b0I42oWCKwGe+qBBqEwqr7iIIP2
b9mCrGwTGDNi7RiuxFsIx6jwqfQ2CDVvjse0qEK1RdmaljJ3tIGZNzs0E4a1L63HgNswIetqmDEg
TYIZuJrufhASQI0g9hNmmkzQhh+Tcn2SB5Ml2WlmWdjb8jRm+4azHIBTh6QTeswq5xtB+rDasa0Z
n0nr/hqbtre6Q5zkiIyznYvHDaA5DJAw9oTZkCxQ2gN8X5HpEYCPR9zTCTtG8k4tiyVzdqVJXxol
Q1snBmldZXcJJGIlerTE8bKcuJmIdXC7wNRpNkmW8kVA3+D6dCZmoSxg3pQYyXHDCHzW22wMlhQL
s1b0ePmxuD5/jDDPI0esDhbbDTrceFIS4VFj8qU0qkx8b/W/n3kDpojXpUz/rQaWzD1hQ7Wtouqf
Tg3ZJNCjU61Hf2q/AoTGIe7/CUgHLg1ba9B1XskG3OXlW/610+q+zOyAIyO8WULy6Jm9H0jKYvan
q5fMrE3Rv1kzsg0wCMrygRKSnOE/Imdc7Qb0w+1uxQrNS0PUcKgVucEGbgJMJH+u88c6FEAEoKlz
dv1SdjgBf54VIvD5kH6LLiZXdt0RQzT7cK6tCkS5ZFAhLOS9mP+aAkO09jKGHfHnd6q0CFUaYIvn
Q5uN5Q3lJ4hh4Dd2iiT55P9WDBFxirXtMQriYxwn03dIPvyTuoXdYl6kCFsCRJoi+wi2kizUsUMu
+lyKeruECeK2z/E5crmHIy76o3YJE1hBPV1+1HjllXvnpUGrKd4ReKj95SUT7fmvYEy1B+CAvykH
zKnD3kBITSQZiXVTdFW899FAU39p+xS5/5tL0LtMIiA5daJHUiK04OufSwuTOrFE4i78vouPcSPM
s3cTPMgYHZA7BIN3m1jpRGv2vQMcJTMlejH8o1Lo+GEIgSCIwWqY2HSh0vYNNQK9wlRT7UzLq5zA
zi3wOknRRIxMcC7qe7TymAG9jioURKQS7mEXSpoGlVrVTAzPmUoVXa5e7ZM3osq59zZxBRzuig9X
aEXrqr79MCMXtnyyQqFtmUmRBWrqEmbF8edm23boqAUZ15d0fQHtppWSjuHW+sifHKKB1hw8Ws+w
lkIBRNtv5n4GPABYSWGt31rlu267PLmZthikX6p0ZWdmhqaXQP6BOWfXlFjd117L+OoL6LWL0JB7
dcEq/QIqA4oo0F26ANYpOvyqBP1GOWiWJv9CUoFRYoibavuzNwYN6XXB1O+jZ5eMnaKyugH3G0OA
Q0T69dUbJb+iwewIqi29OBh2xHGFnSH+R/CzqwvlfZNLIJtoJ3IdXX+JcZJN56PtxyJms/srHGET
lDbOFrySzJATH3KtjA5RE0sGq0q9xZwx+wdxDRWdBLngxM+eBvUiejY0hISQpGxnb8tgVB45dM/M
DmBjyIHx3reXLGqoPhyOh0QdhLM3/z5z9njm83nlpUDVtDP22qO2Ez0wGU2yU5SI7zzqWEJ54cMt
cJoIqTKf00YdMtjKkJ2BXqFfE8Lc9RbOQPBqj4MSPpQkHVCtuvAMzHKgQHMxFZ/QXgAjM/UdGfgJ
cB2usE+VsigLlzhCz0g5Vo1/B4T8UuaK99H03dGQGwc1uDyILJxy39L9/Nplc4ohoogSYfLcCPiQ
/51f8fXRyUMxsdfGmXQq43fq7jkFx6YKZt800zVINrIRYDC+q64Ns3bmB3SX36Cnd2ERQ2l/VV8S
5DShcM1pMY5aiYS4pNk3l8dM85vgo37MiPP486VTIIvA7AUKOsgRAkJiuTo7obkFYp1H6/XbJyZw
sZv33CI2HHKEpfmwQ8hzD047Z//8SuJDIiMka43BIDjn3kMwe/3w4Bs5ZZ/tFpacFQ1/U/QxBT/r
Mccx8N6fZzxBI8xIex1EiHJaOAJKme3apV66orSqBFYTmUlP+lhQ/TyWr7Oq7aRy+/Y/yPlXXwLG
6dTDqhHc7NelzM8lJ9Fh2EPd7SQ/cClYpX539C/ItMkT3ib/JfF/Mb2nRmnIlceGCd2Kd/7ykXJ9
ed48jGTJjbsma3Kx19H7zyVUKlcIq4EVf+fN5mv4ShmBJss5C1uCIHyZFlHmCiKQib/Iyrewac6U
/XxlXSSN0I8PPLCJah1Sor9RXBOAMXQvGedrCgSKDRWVBekmB0K+jkovGt3w1zIAFREhPzU/uDpe
vH8lt+KZ2vz19W20oRh54F5J/vHz/xtlKLGCiZl5VL/eRi0XtfFkelBILnN2UbeTpwhA8iuqvkdx
hHHSkURUQMycKUD1egX2GuktP+ni2BAPKFRZDhK7aWCVdCyS1trKYIQEYonr0VYhdZnf/BAio+88
VYfWopgbN9rkyps9SUusn0Jeg3GF7oLAoyVmDGDwKmWE3Lb7/MFvKDfKSgCMJ/I9tseb5897Ch4y
vi/Ox0ctYkg16q3/p2HD3ELdZ44N74MWkhGBKnfftKMrmhLYutyHQeb9HQPu4kXy9cACaKLgSfhm
KS248e8Zv6fZZ4DwscnaAxK5VyzUVobClLcGKvkoGSm8XGFwgMnJBdKnvp0hyvxgkKyupcj5UpUe
RWCi1tx9P4V/pomaKG1+DM9Eit5ruHWhTXpgyYeFapmg7o2dNiK95OHEgoU2WFWUh3NSFSLPMZPS
z1RtDaJ6uYvOvTqVFiAIf0VdkEtf2eOMUMhj/u9JFIxCaKj3wJq0djBNWJJs3PM7Yq2dFVR14f1i
fKNdnIGSHPXOMQj25tgbiL/Cb/cOWFuGD42qvxuRwwSPEQmIJ7j9eEtNv5IDgfnB7v8wedXhxIXY
aAe3YnIty/wjLTKRwreG7Y+TudcgzHZLDNvAfu7o0ovHUUm0A6BXirRzN914F3WExhGJ9i30wOzh
Y4WUQtJxO+EXjzSa1LVo/HjeD84Cn7VZW17opaq+rJxFCSjsdvpWMhbX5xBBWG3/pxwxJM7LX1tP
GPJm56HXnJ0SwmHhqQNqMlNNNUeS6e/mk3dxqpzjlTl5j3W0MynpCjHbjYnLALDEEAkcK4qTGEPN
8+udFBd02JPetMgvSWdUBRtglWFIEFUQp7ySWlKVioH8XSklWDltO649kBcWuiH21neZRtEEh1Tu
9HQdggLex4s/mbIsUkvLETW9NqF8bb7AK9z2KqVYHmkmCPO74xFQtTrGYgL0h9RXBj+3Sc81Jrdd
GUnxJzQwWSqpWEDslttVo/6kuHjgzIXxhI8AqUz5/T/hNonNz+laGtHcNhWs+ottDb4jy1SP5cZ5
01ojixMgPlfqTiWLHqJgeowzgxte49qCjhE98UoXwDklix8mT1MuXuWd38xcRuZ0iyV7NqYEcWN2
g8zuV0SFnvfty7cmO8c27+cByxSD99A54yUyJpXiyWFt3+QdvGDsvcAO7f6mNPajkNaQWgw0yb1x
GFp4QxTV3nn8OCK+3/t9lXO1WHd+u1sN1fyxMcLUSt8nAdhMMNlBQ93q+nrLX2T/lqr1QXKIXJ76
ygYzO+lPhRN5SGMIhFQaiDeEHOY8VPr3NGX9YYr8cF2mvZb+ei7YIWlU2AFIEh3x677SKo+lDktV
OV1vgHyZ8LoPrkT4C9DRdsB+WKmQeeGx5NHlkqxkkZxTfg22tF/FZ+4Q6xs5t4egbI0dDKbr4lI/
G7PXwboYZ1+29OaTD+T3u3GJUtfGt3Nm6ZKpKQT84WksjX64rzbeU5gsAhtzXDqRHZQCMgXxZoC6
r5XnYC6x/qg3aBj7Sy9sPXkOQXTlROm+KvZUYPZHjhC/+JXc7e9wYMuIYOnHZOO02HP5mLOcJhvI
lbp+zGHKz9imiCTRuQeYFPGetJDG+wdIsNtq5IO+lKw5vKKOUE1AYzU2CZMwjyjDYzUxhnV08Sm/
B93NOYcVxPnVkhiSKigPVKJdDUmYIh/X1twy7AJJPDhwuepQ1a0wWP8rSj7z9zC6NB4gvW/g+vaN
QzWz4Fem3iPLJPsqxCgwzcNxnGu8ooFgLGUJytQJ+PxlDSuPgZgP+ynCV2w/TI5uuC32KY0IktUV
xhW25PcZuccRv1PVfjT+MDiS+oUEpYEgvM0BLtPY+yEbRWq5Fo9kVafi8E5cMoekIs3vMRSa4D65
jjtGgluIsapDUULG75YHeGeMGHqfkiFOq8bbaSU+WWrsSZTlFk3pDX0+jTtaLmxk4fCrwqpzXuE7
QylCab1DgAd7MM4nHhzq7vH8qs59uPZo5JWEATOQ/HaJz7YOo+I324azrnWNYwJRqMuJAQRzx4D6
k5lPXwHVjffJhtpG3fuASwbdRGFY1/7FZs/bHoz2btJTj88+kj3bP6mZysNpdrbNf0+mWKkQraoa
wpEQrQdR5az8ULTrZyxQIvbLcWMv1afgBUjozXFUUq1ThnhIDAQQQcn1xDTAOJCi8cInXEVVJmid
4FKBsri20c9pTCDXVsS2HXH+qGrWQaFi5/mmy5I5YcOwdLNQs2qYaF8tUnSBzmC/5ZJuj6UNdPju
BhdwXc+ICK6cBUNcuGne0yV71LV8u/nGoPaBzaWg3204mhD7I5bQ3zwMWYFZcsLPYQUl6Yu8Q61W
aCXcexMBpbjitZGjSY0efkjqYAi+b/wQi8Qaakv7syI5KuZ6AyYMv6uZj4QYasFLQfXSfzAah2sE
xsyP7ry91aGEY7KHThllDvw9ebIDNHb51/DmoVdRhfzUvalH+SDa4SVqsl2mFT1D+yFM0byuMjiw
Djri0P6CKtPf7DwqxOVwWf6EA9go/bWx9FpqscVOTtGUBdHjI2u90Zny9Ov+Gc+yP8xiE20dHInb
G6/a26KTma0HpcLdkm9LjIF/bwGchsd6pNP/aRkY0TCNGNplOp0Jn+gc6aSzSzwcGctYuaH9TDIZ
C4GwtdMfUfS8l503K+8m5ljOdxszeTao+cXsc9Kopq7VG8vGT94qsYRrHAPGnL7Gm8V2GAZ8+Frw
WWrx8YnEyloBGyWonIEYul9yQj6pZrI2RsMVCshAkFbO3N59M+VT3vEjo4dfk00meaZ9c+NlHyqz
J123zu0hEL67v3gogDGX3e7YiB2mq4InTjYIkuwGBhcy7NMuPfficgO7rOqnt8COzRGlUuov74E0
sPBGQnEi1W3p9ir1VU44Js1DZaELGrgPF8ZzMUoCbrWY7MvUqnE5fn3nPY7OfUzWVyJGZd1EOydD
zJogmUKisIFC/YkJA6rAC0p6j3S5a6dhAPqvRIxgjE95j1hzkWi7mHKVKSGKydsonS9IKt4IqSew
R272Pb+7m7OLo1GhCGnejoxncFzVfCdKEmGBK8O/yF/qF9y29+5hubDvOP+hAl5s72tGgk2qRk4W
IcS68FkO2wEd0SQjklg1no3swpSC7cP4MOy4sru8u7OeJ7XIJLCH/6zMnRKq5MKZNZ6Ldr53UnLc
nR9W2jVVfEQVoIMVm4o1DX9f483/82Sh7jx/x++sFTecfVvwnwiq4rmLKK+H/R+7u7gixQG+fzoH
tZzW6Esp2z019lFgBMtZPwumugYKhL+T8WOyJ5Pvq2e+06DPENBq6x1hxtUi90jaN2rmBQ9d5wiY
7yWFNqT9Mk3/DycRR6bK4RJNF4YKMM1yZL10xYnu8lzewiXQjbfXNgqqjUuSXI05njF7TeS0AfDH
XWNR4r1xUC/O06fjSCe77MrxDfMAPFlFnUdOt8bSfGGkdRHNV8pLna4pjlipTVFv/j2ngIaZXO9z
qnj+BnR50qujLFEDJZXFruGJuNyQW555EuKfJaFNSBFJkRb596T6Vfx8AXWMpFjFaZk0y0H9ivko
wW08h2q4WnCe7F9EuI56tkUmCNJBeMh+KD6LKz75zG4ZFoyJSD4XQ1VA3sWRf3DH2iVjML0B1SfZ
Y8/0ThIa9PsCO08B3LtO1jZntqB310+KFm5ibCyNbnxDuFFcmlchpoILpwZ6b5IA+Qa0HMw9Qd3A
LoGU+pU3ywr3dGMXuldK1CCw9TpLhs2sa8EehxcGyAKQ0hVdj1cdIrKzTvq0YT1k/axTLgSIfzOS
EDo2uND39dAKvGgE/pwPZCXwRrQv6QPM4RHeJjNylLed2ROZWrIdcRqvmB3JX8L9pGiw6PqRGcf4
ozu4EGC6TyaR4FJFaiK0ZYHSUcz9iJx+E2CNNLA952H/BKO5zpWcDgNAU6J1LiEzWwsuzJe4MYzx
ZdGf92QDCQAYxQ/eZN2MngTMFFAgwe4vSOYVCQuzPk1JX3qgwrZMn71mxnvdSN4G8H6i4r3evyNv
G2wPbdhTw4gkmWfxjYp/TQWVL5t3bX8mTkz0z7k8nwOpnOXDAlKw6T3SiF62g4GO8Qovu+QfwvoA
uUsmBV+lxmG3x3r3nGMkEF2bJ+9wndJj8nxA2qFCo4bu5aNYWjOdTlICkXjPbieK0dgy6VToSxyT
HKTlFamad9eTQgTgTzz5z0XuuuiIl9cwGwJJTjKAF7Di4vZ2hjAZUl9WpZwJLArBOk3mYTqMuvGa
pceET5cHuPvnWy98jTWpvO9jp/gwU68ES+E8hZFiUFp12pDuaUK+WW0ykYkiFrcNxgoPC1Hyv2Qx
X4bZ2ho++0CtYSa+/PcQmK+pNQbDtOuWwq0GeyJIMcb1/mopLplF1xqtPnyUoapcpRpc9hgOMuTJ
eVDABNi6L8vVDcLC8OEOnXaFMOx8uD17trnhsCQ0D+hP5DPf+tay66ECGIFzsb5Mp0hLoTp+PKpX
bapljP0d32rn7UUiYFBYISbQe9KX89ad4gzJMGiNMXne+jy/snXR5F5eieingBG2uAhcq1UOrWWJ
5zIiJMQVcSNlMSRooe7o4UGh0+El7joeMGUL0z4xE3JcCDyeJl+vvrcqJ4Of5b8HLb7QJ/7II/nH
W7MQYIrpWTfcwKvS7JdJ2Hvu/BpkEOkOKyn8NdBpb/LJj5Xnh6rKzVdjAb9igdADc2nNB95XoV3j
0Bkh6IjbUY1HLZkJiVJABgK+HEELPTdL39r54sGyYkChCScpcTB2XqZpU4la0KCwjnczNucmSeG3
rsSqHbuer/s1kYxyCDHRdD5Wi2RumZsmjTHREa9QKMgywfhFPoGDcVL+Lw2beGmYdBhJbVN9N+AB
eQ4ipAEPuGyGe7//hefNjS4vpiH3yTUwm+xMWB2dS+kRQOvDHA+LOEe7DykJBxt60FwfNyTo4/Mv
mMxgSu3s7KnWIC9mwXurUAICO5FI22RfwwvWlb2c1gLcAhsyAY3Lxfqo8FzYZAvt9sqlBQjxFtHN
XHY1Q74NdxeiMQtKkNzhEscKpBI8Pmf2X8POSMk9U5f6F/XhqoHjwUv1QNDOZX4LIE0xC2pUBzla
t9jkehzLSKSgaEWnRcMOVIeufyF6bjzkZ256ttPzRlUflIMHSVexXJBJvkDohlf9hdpbWe9lSuER
ats8+QPG0/hpD2HxawHsM9z9RFloAn9gcPwbf+tW4m4+cb9lZ0VzIsb0YH5WkmOosF+G9nbjeJyO
w4A46UnksicneBBO18g0awGg7ZyS/6qTWLAlTLycqldHx1eDzp74n/hTTCrDM3ELfTqYDtHM0EiF
/J7LR/6Pvj28EuVqpLvVU9qUr3M03i93C7BEPSj27P/Olph6zY2lQpOkm4TNABl4o/bj2CHqYJh3
GbPXEDNusKPH79CgCHrEQR0cnb5siBoXYm5G/BYN6Z/krLSh/i4o8sBsGPLSqzGurhjic0NiLUS/
z0XJhnpDvvdk+MVoI6vG6Jb7gtGARQvylxrD/NGgjqsrU25C6ElElAZHengLKR/6NsN9qTTLnll/
pkUaLfso44DdXWcFMd/Tz6rg3kPgE2ZbwDYTmxaej3zBZdSZwDiCnmvs+hmguUKqjS1Mm1FXLAtb
KIk9ij6dU0IWZgzYTM2O5GXF7JmuUSrJ2s3CHYkEUnyBFR3A4Xs8z926jJmJx18+FEXhe/5GVC04
ke0tmrh3MPUwCdpV6lU623/vpBo6eWRNr7BET8/rBxGfymEi88LDSV2ActufTkuGs4zritEd9vWS
wE+SA7/ysaaHZliRggHH2t6Cc3IAsreb2wiVC8/PIY3X2MPE7OTFQ8MLpH7m4ab3cJlpIoTkJJes
ni0O8LKOlQe5Z2UyhTORWesxd8CXVI3AanjxdHuNZk39rdtcLxE55s3SyCnWqkeY9DGPGLa4Zxsg
NvrLCvUGMxd3ccm5PJLKwaf7aGplyppOGd6FpnFVMsPVwB3YsutlQ6dzWMDJuW4/m3LRSQBbNDKc
ggZQqFPYUh+PcA/UqT/Vjj9ZoBkzoZN5CFufnuF7p2cA8EUYKeANVmSCajfoNbdR1QTVc4k6t37z
tf3hvZW1ueo70WnLPRQQdHUSPVCRXfXUoOrn2GUD3YujyiGkVwg0jg6OZ42BCdGygzH3UQtU/WCH
r2atHDArwHrTCk6bWkvg2LI1xsbeuvgGhqY9FdIQt0zFdNpMgDmWxHUTY2J4GtxMW4CqiMZSaLZm
eBQg1iM3alCBcunqqfyuadRXV7uxFT0i62kNSrId2fGb4b05j/ij9EZhJs7XeR/wZshhG4KittlH
h8bkKJ5jRYQ2HGcg/q0PAmDGlmpUwOocijKOZfcp44Y8ppvySVLPL+XkywS7NWggaGLTr3p1ZSLp
xDJIXd7ga3RJeiKgjn6AMZUx8Gz1mkWM1PyGCW9cLErGzMFuLasrbR0JFwg5N4yPhuglzzG6PcVb
TO9BXjRXpnwaIYkMRV9dH3me8+4VKDFHQl21OGx1EhF8xMdpnZzW6VK1PjDO4EuNV0kOqfbEn7I5
5woZ5N/lxgHukiCDQ2P7ew1fqSRf2nqErUlYfH/+iebdR3YiUnvMl0gbCWAKaKU5W/1eWRWHNbdq
4mDSeoW3+kMIUfbdQCi51cpr3bNLT5wWZ7d5wnzkOrKjPNVj+Ig/4TZlILDQFpQTriEEkvGSRSGg
eGj+Hr7RDWn4/dWU3pN4U2tCtHo3PK8SSnypQuxthoMvhaSIe4F41gzIL7qCvUBw5jM4t7C2oEfw
vsioDXFRkkGyUFyA6qlpudZpbvzROirAOJyDFYj7q0OZCR2pnHkwD/fDtUdkJ9z63V81zVUbASyd
TEeXDZlkx1UQrj2eB3e3hleOv3fft10FSVBYwS/uF98OsaJbgmqGLZSqsx/l4XSZyKhXr13UlyfV
WIN+IWHOLkXkK8n+WDS8jrOT1Dnioqo9yDingoH1ArA4WbCWXf0OE8Fw1/Uuu7fcmAFLFuaMgqk+
ZVPRz6N0oDGc0v770+JW7C9iho0Jl9mRgKwNW0lwR16mKxf12SaKXy8Ehpfp5ctvW0dVRRIdZQA0
t9XvfrhSBdTVg4sPUQDs1WoVLHzn5eKL52soH5LxY6MismxiQrCHcnZDmp8fFksxyovVPp5n8WFe
+ClJL45FvcoBDynJcgoPfqMoSmPRyR6ldXpATFp4case2Z7+0vL53pKLaY04yC3nl/BUkXETrSCU
Ga8Cf7hRpAcJNtnzgVbgH/x+jFeTeGd8VoVxILcAFV1WsBvG42qyxSzp366ncWUq1aghTc+ouhSm
SbTS/cftKEWqcMTkA8g7diDGDYn8xBiCI8mkwDwtGVPdF+D6X6N6k0/F3aGhjz5m2Sie3HhRvuTQ
Qui5uGSWsJyAIPyZSOesDoC4QjY3rUmFFNoSoueYSYfsNMCv1V1EQI0+o4wBrl4myjR168ekdD+T
Lx/ZIkQS/+1Nc71BvYijIPYhDPw9D5nccZ1Vz2etMyhXTOkN7FiMsD9zMR31TDtf4IIkWkDD6uIp
QVvWRXzMqdqjk6uKtghCDpcImxxQG81FlIiKQuby8KXf9UaPMeuXZnVRHHnPeuNGDKW9SLDYxSG7
dNHaFNgD7ZZVVyjh62TLZswtBDKQ4wBmSrQEWosOZa9EEC3U6KT6AkMXY8Ixdw3cN6QArHIw7TLz
YBEnuq4eMRlGI5x3R1kFDW0wXV6HL0fKKNKkk6pTj986MLh8LDUNTSIc0zCJRvZgY/QGw1OInnGM
R7mDUQCFRDr61BAiaOZrplCBQv9XegpEEG/TfFdzs26f786LKpSf0HX3Fzcn+5TC+Et+MKu73B7z
N4Y2/ngBCVR99b3AtuK+K9YLPdTcp3OopbVLpikf1MOZjdAoSKzpowL6DbtQYKLttBre8+Yzjc6b
2vhlNnAgpli08IWDp1Rst8G45x56+2syOsDuQG5+p4xPWa+SmzQkxszoDjlw811/tJesdpiYvv3u
hcEIfeQhlkksoGf8KLXToyiKTt3eRsLcOOrZQiue97o+ijcY6ISi/OJ2HJoLhypzvebLz1Mf1chk
2AGZQ2TA39s1FaFzFgPgCDY8uvyXuKT/EIiIdrsnyvqDSARxf9Ppl+8tPjRPkBNiw4Zzg/xym1ih
WY5yx68XxgQBzAB3nN8b6CRTpzSgWNyQoHmuS5ZI5VW8wrHjw92+ZxUynLkapvzgG01+XlxAcaPh
UQ3Vclpe3Ao8JKRUeu7Pu/kcXYIv3E8L7xY/9BekRfRwSfWvIbZ4+DHmIE8w7vRlz39XJd50aWxg
lVkMR35fwsBiD6oSth2OZCoKIKhT1E+SxotER5yqRAFWL1W+DZMXK5BZydW4rAsUVoUIZp/jBYvA
0pIB9xTWOTksB6YVBZEbWSffTygkCx5e5tbTN4IECPWtOV1i2q8/2nC9IYS212mn7aV9GZ1mHZHp
VexsRMd5dXiMaPN/eaOe+vjZyCoJ9T3SSbntrhBNPH0O6/ifpY1QPAU6KPE/d8ZGC9m6EE2k+ChJ
FSGnk9uKoAqIj+MVIC3+ORpG+1aGwjCqf4PKHtZo6a+UQe62O5wRKKFaIZpaBeQ9VWiFnBPsm239
DdJOlKwFmLKe4xIsFWaYrBoGFnH3xhdwao6ziBrb7TfiLVRmzpw+6fTNQbwuReN6DuMsppZnqyHV
N7d0Gg02j/ebDIt84qOOdenzdVGj+MH6GWDzgB67j/e+kOFO34zd9wLWCeFh2Qx0sh4QbWNjTQ/j
3L5QEaq6Z69nRznHpbtX1NSaXXeIKQmnaQDWRwC8oz+KV0FY4VwkRlK9z6sG0pf2aaGotQh8Z+Kj
czezegWwc1gVF/pRV05kNQppxZi4+OGYXdHHj7qyOLcOUzZB5v0fQwuLYDBn28zI/YuOmoydW6LZ
NEfKuWI/MNIlCQJNvjresxvVb4HJn7r/Bl+HnRmJmrfOWFPqnGZhe6YcrVqOQyNnpsbii6pEcXYR
IYadqqEVNHHLKQmDRWwa0aRf+V6dpd7+TtvJzlf4c4jOXkMz+hTI05Y97Uvz0o2u+d0oZ4fiCZsR
ynsrX2F4zMuOs4wicwFWkHbsyFxHQHRn7/ejNOQ+KJmzbDZAaNM1bRYuphEnqver9Ff7DlvqX8Sj
JbEjbX5jM1DwZDKNA+0Map1ZEfdwiGNcza/VsI3PT5JP1xZ5GFX9TpD6343eNy2XpSNgDTY+qV/t
jXGm9FdMkeHiSEfDL8Ho5Qcs5CFTguPblIPnqAj5HvvZ1/XeOhBt3fb5uFA0ix+UPdU3oAA/+kvR
GdFoeKjgrpcgfGGfDdc+6K1WMtNFSR57taxhpisBphiTj8Qzpmp99Twk1FKsalvaml8kkPGVNJA1
k0LEZABra5YgdRJBXjqvtyUJG+0UMVGuHh0LSvkHHTn2UihpbopxBzudVmA6hWtlq6VctRgnaY8W
bTOqG47bgS4anQ4a03g4XYIT8uUQMLijMhjYOZ8Uv20+vefj1Jvgn0t/U1eQfyWVJ4g4GTdbNt+e
22C8HfBxIUeQljnDk28ShrWEC3sfbbhpks57r+qEZs2BtSVwQZPlqDitMvwsgmqWIKUkUN5VBIML
Hv/RLRoG/LxD5f63BTaYeetDkB5iu3QpNvYY7gN3i5sNLMBvGLdhj5W6NEabf9Tajvl/upImI+Ve
+bAEQNOnbecALIjGR+BqTbrmXjUXYHBRsfgI04HpD2U/A0A/u9RzcO7bHMh8/yioGwZAxkUA4ght
z4hkwAkGwL4oQmyTMW2pkMb11AYwnZUk3vCEGrO3BpPpyFgPyDutTjXsQOkQ5Pqe0WZLmuxgbKEo
QYe8zMdgrBbkRTFyTt9oELoclpi6jcGMUuDXtzo+pQNKgpABy5kU/z50IHd7MoZfxBRVkgdl/CBk
qrj//dQeDF6wOk88G9hWD/rih6X8zUH2c+IdYapGRLJR1F2CV23vpsTRDGtIfl43HtNn7irbAblq
Moe+H3BD1VRuSbe+45Tc0G+HjHoB7iFEACaZJ8HqN6ei8De6mmMymYHsFSlnEh2CrmMtPDxhbWrQ
OPM5fieI3TTLUQQuzOAoYNTQpkmp+LCuFnvunRMpXoFgdgm0/XhJUE/i1VTfmvjs6dlvclaxVv4S
ZW8w9DfBDYC2ImViR5TC1aowztkWG2VywOX99Q0FIiyETAa8Tb5+N+xklyh5veYQj5hjUq7YnL6V
/TzQIiJ7jqnjVrxdKq+xv2UMLrgiIL3LUzaf6MUIPlPEwL+w20MlDzUHOFN3Pb11IcCmOqtP9bLz
fnx6DhLszDconVqozHUBBNzSBkIw3uQkeRL71IR3Ew9jtSlAfmeWUGJfxT/y8nhDUEs+2ILf71Rb
51ujHoktd+xa4G31jZT704JeHwplCuCHm6PlYUt7u6lmEw98aDwJ6RyrQmu6OlZC0q/DskiC3e1U
InWl3Bw05tguolGbtDQ/zUHMT1vDmMqxRC+RHyZveOJLvRw29cHILRmn5GuazI8QQDoyPNUlW5C9
uptJjSf6esOF67PIfj5Gwf31+kwsM774d+FTgwH0hUQPNdrpWeQwhZXA4kyJ1jUF0D2dyF+ko0Wz
rq01kUy6L3s15rCOREsijs2aONWB7cPh0gQbo3YdHa11ggs/mxwAc68gd9S7SWKppMqoKawVszhV
4fDH+w8UHb8J8ai+eWhCOKMwoSj++aMdqc6M9IfNE1FQGmfEpDTs9H6RtIka7didQRlMRNjKZ/Tl
vbxp2gzN686N259+j0sE4W6YcKv0LXNwTi9KlRvPtY5aGGy58kbKP8ueQ1/RXtPMhfdchX2C4xsH
ms/MxL/nfsORjNbCX0rvwrukDC37DA7s1fIqFFD20piNl1jWeJ+aFfIIhtKPxrRjbvG0u0xrKNbU
l3/p2cEYFx/BVFLqkG47IfT55ez1ZduKlN/4fbPV5LJnRmbK5gGD0tYI2nNkGlgW4yWDTHPS167g
Hnhs7eOw3FhQL8zp0IALJTp+JvgYau5wMuQBuuZGMxte5AUAzcavKoOGd8GkAuOel3dUS1knhayG
WhXUPK2UvRogDLcl21BSYhDTOFzsDEXSJu+8bede7cHT6kWMNbLnwjxipY0jTVP0P+L60Zam+0Fe
C+h4fX3UOWp+8q2/SaQtgkZg5aOxcHOz7v3wk/usyasuDLeoZ9mZfjVHmN14R0luLg86brpNVR5n
uwZpwc/MXqRPLKL6vwGHL++sUkk4qMmfkBZOGAGACC2yDm3UuJaZGm2H/4m1KtGsi29/pU4+Y9Xq
ZO6k3M13nbVlKJEkiGrzdwDj8EllU72k8IttF2qm987fX2/S7w+qKcl8S0mWOW4lfJTc9mAGOy9v
f8e2y4ZDpUgs2EU3NUhkV6Euflb31SiTlPvzIgMlndp9J6o5NR8hBFrt8WRr2c9WGBLtP9MAQ6Xa
L1ZjiDUSBv3XroHrvhGJeibI/+cRdq3EHGZxADWiQKBm6shLqIaW9fGgHfHRwJ41CXb65wH6jOei
uaJqgdHakWta6VhGJfoopu3na1bYVkxi1aL0II0s2Iuvb0KIpf+WvGRwLhZ7o70YhgUihq+zkMF1
aKR2DPlOzHL7m7alNk5ebFCsQJQpzLtsOMYQfWXewYMouGmeCAeFT1vwTHbEep/01MldelxRgKBl
eXna69JirX4fUyUGruG3dp2HkP4p9pd5CFTPVhzca5M0N7aoEIurKkRR7vj3n3NxNj+WZtPvpwV4
rdiiFRYpvSQ4OBo2wxxfeRZ2Y1n22OSEIRAeqWXBJFL6f61cry0HXq7LeV3m23IH7nUQwr/eGu03
FLcWKH5CqkiAKxLi6C541v50zjJGg/KcToHhNQPpYdYv/IkjietzTHbCdnw1u0hfwuNptL3f/nuN
urin9nD1Rn61ngEeZctS1GtajbTrphl8eVIj7exCWMXCNqKJ3d2IfKNMGfSle1R3z1b7IYJRdJ3Q
c8CbvYe1SwEU0oG2Uv8psMb4HZwEqc0pyt1cpguZyssN7H4nlLt6hZZcJT3/NbF5mYsjglZqlGC4
udBtPZ5Vs9VLaMLdNioGhV4Xnnj10bYepB0lHZVVqmuY29dk40sC3FSr+tTtDZQFn2OG6P8SupXq
obmbtWg5us11Q1M1fG0W1aWR22dnh2+obHb/0PrIfhnPAtGhxOJ/Crk60I4OljHRPYrZOUk07EwY
fUJ2eXxOXiJuYx7/MWdADJvwfepNf3+TBDnznHTztFtjDkRQuK1MuHeMfgr9s3A0jE0JGM4kO1vF
a1IdA9ftRpu40Ye+RixMIHDQMR/EgukWs6LeN0Bnun+miWp7IsPWs++yDwgfWcHM5FHSI2oUXMZt
cpiklxgSfetpr9VQXIV2j9bDzOpXVNxPwydCS3ieJa5LwEwjFLTxvFH7zx2ZqXVIwPLdwfmxMgmh
cSiOzE3W6512b871SO9Z4msm8nw8JhVpsn5qza5/saREdmDITl1h/E1giZK0V6N7iOSEW/ViFoq9
x0lofvoQyPh3H5wPUzkIhOXG88DyKyXAsY9YBB75bDTcRqjCnVZdPcpo8iytcs3/bProISU44654
xabf1+O4xqc734UQ89xHt3ip05k4NEQkNTSTFXlbP9020F4DG3sICI2t2ZpsX8aTuiNhxtQor8ub
9KTyXtw2laMC0gBzyCzH0krU9x9fymCQam2nO7PyLQ/7g87NMV3QNxp9uSJouSG9nnV4cromvLQe
mVPpv29pXT8/WV0lrxtzjrIPPKQLKzccDQzMgc0Y398TGGoUdw8g/HFfJz25CY+gHDUXDEcoXhpx
WKjVfF+DbLCQYYsrH/8FKEEvncV8n+/tkXewk0mT7bJkknXtWSmbwOe4ZAVwboqL0d9qfJtyBfed
No+Sx6/uvkyvC9fWfWZ9pSyU3Hc+VAZLc+5L04SSc5p/nfEdapyw0wqJ906NfTAZPqhIcYFeXYnn
hOvH2PQ3VjEuW3tbPUr4fS3Apk98dFk/kQwrwOPWefryh3TMAFvISRjU6bS59CbobNxWebMtgGSY
8DFFqtt4v+GktPc+lfniK4g5PYKrNh1r2OqGuFYBailAADy9Rxtg4BQA5uHxobOVl/gA56fk61XT
Z6vy98cKOFYzUlZWJ2xpGvU0IdBeVaewstCVLYM/yYdtML87nFrf2pn23jkSBbC2Fnd58V4WZu/f
S9rYu0tpen2p+KoNGEUKagJuuGoP6gX3Nt5P826N0+gHI33/9bgTwlJkWELQZ3Su/7GyXY2zOh7q
3ac4ZzLdq8iOTREVGIUN03QTrxMW9971fx2/qC5xm+Hdc1iQvShzO0chkcJDgP1iJ1+jWkWxfvgM
mIBxgmocEKFeKkzE0+KnmrFvIEyysMc+gKMmF09wUFUdYUTjWl6yh42vIjqZu3RESYw06UEV51W/
avq1F0rK9yQrWzLMD4yuWopsoqwCCHQUzP8eG557GiuluTik18HyRwk8FRjjyZ97jKE2dQ9QgxPH
TLbsWBZ0hx0o3q4MWn949LofRjRIRd8sY5GyMarIKk6OW0GnEpyvUvHtl2zifLth6/Wrc+QvucmO
lMxhkzIIHvR9rAEs6i3NM5aQpV+/Q8cFGSpY1TFHEub8aNEZUutuI4s3PLIdV8jxu2USPeHI6wjl
DYL/ufIlqq7C3fs3nk3+Dw7NANXX6ASucv4bMMmgyua4+SNNhN4wlAeCiE00N0InUvg5vA17kfxY
08fX6OYN6TH7vqQCw9sDciHp80M7dbTEtw6inK/QvF1IKlMuiL87IsbdHrcpnyp5YKSLCFWA+MSd
bLIWrYCk+s2j28N+a3nDT8GvxiXsAhDQ72Q1Nl0YFrPuDhkkTFRtJG17+U9Lw+6/MT/B4Et6LddW
1riymVGfbh7J9mIscyHbSPLQAEMKteVLHBPwQL9KMlHOgsoIjZPT3bLL+vcdenhd5TWkC6skDiU1
drQM5oNNTiHXITHB1OlcWHWqriK388cLvz01m4qzRcB701aP9AyMu2wwFDlRZ/hEx5r/DdlwznMM
AnpOLH3FVv4LWGwkcovls9IfK2RZ+1oKZz8t9c0+NjWvxaPnP0WdgQjjKk6p8v7x2Mf1JgF4Jz57
ldYoGvSzML/yXjtRIh5ZA9smxjzrdP3fJLVI8HeRk0ZvhmuVTE24UNQWzFwnKa7tVN1V3WweEun6
Hl5tcHGRY6qsriEBhzRwEFLMIIKPE3VhX38Y85G5rvZ81iHMmEIPdk39GsnSLrpxWXoiCd7J9bkk
33wn9seXtqL/4XZp3LlrUVDGUAk/qkX15/GNITdEof6YmaT/3LDE/ppzVSy9JT+EZ5qRnm1504y9
8/olKutOTMyKIX5Q9NMQtFlzMMRRja/uRkVrZLAcKxlPPDZ/0i8N7aQ+B3Xro1tQsmLQQ/x8aS6G
cxOxSEhR9kyJ1SvrE408CKQ9bIahJYvz1I+QhFRmhxLe01Cwodw//YgLuaYVS5QwzYEecVLApoGo
gDX8jG3vwaC6/u7uNtAHH1uNWPbkQDHBZP6Tgeth39IYdvvOENtzHLzmXBc1ypOBhGBs4Trocnso
scFVVjjSDs2UtSipMlRMa5xBuUmzsdAZxtF4EHHP58eg0jjyuI9soPncatMfQQujkvxulE/oZ3MZ
/UCVM99Z0FEXUJ7F2pSVI9qB0FnexJhfm/PjjsCP61CEaSM9TK3ZyZq4wkfuUDEN+srRtijYiWi1
8+QPSdz4NTQOAnv+TLj+m89Q1H7DeqwjYk9rhO2wWW7Dafk/lL9A/QDsstRLjVGhYTG8Aw/n6EhY
fM2i6cxn3yXz8PEcXaO/LuEpc0iHWrt1s6aofQ3Xk7blD+fOOAMkwX5JZ2LGpwnalujBXW6qvdEX
pPOrMrjHLrvpFwCkaRpwmrjHStWKR94kpoFppm9MohprBftOS/RUgGlQFCwQbRMmJJiGIBP9Boob
wJrb65n97OOgOd/rGHu5/a0/bp3k31wcG7L3dbFCv0zp4AXqpheR9oXtNx1V/89hsmUqsyY9hyVV
DBh9Y7opdsp2kFVPPzYZhw1t1jT2Nj0+woRlBzGk/b7j9LZ9C3rIIyVfi41Zena8BmJKt56R2eD1
ymO2mDgZ1CIxkXwjhc1DTF2OjDOMc9eYh/bdJQdsRmvk30j5oWm1fhdpVMU/fkRBHyy0bDlyTYLO
Kw3W9IRVPgF8nsIG6ixtyCXeTrfOhPQ0HQxqO5zTbNrWrFfNuA53ACfRzUyN2pwxXMH6FOZrqexf
u4DNQVNv6V0PfjYFddyDN/LXAekmEJeWOY6h0U1CNOhwzsU0IUGKAqa9v2ARXy1UngYvug0dhrby
BCJx1Ms7UgdKvbuiJz8VomzwNE7GItn1A65KDYvSf3dgUpEZxFycWkofjRky3A8RwKINuakj7+Md
bUjVVymF8BV45DBi9Pbb5oMrmhrVs9fb+u32+8trHfnSbry7EUOGBwcKcR+RllqLlFisxlt6sYbS
POL5bSm3aWvp+QQYxFV/7YR+Ezo4lQPKPvf9upQRocJhP62Q5OQf6+sCmg+T6g+hsyMVDPGfbhux
eUHlt6yAsCY5L69kZt5FWlpG/CV6Mnss0pWh+6wFOGsk+N/gF9+kaG+n+S6CTN/XPX27NFodwraG
iZJUGti2kgTDTC8geA/IpjzWZ0Ocf6E0lXsgeZXEDI6Y63AmiwdGwLa3HVWfCkCBKtOLs1C32bKV
2LVqaptLCsK2pus0elBx5UdQmyzjtQLSNZCXHLL5IrMU425wWN32EmjZoaEQRdXWfLDK2FgYIGKT
CXgQD+HkKug3uHG8ehmxgPpguFov6bYOaZsO3aqgznKPe5nCUractIyGW8y/kt/PIVMx8+uwMJvI
R83VXuWoHwJfMvdtxw0Z++UzINiJwCT5mCuYzpEqSthrCxoTevkEyl+DxECQ/xUMPm+cDB9RYGXm
zbw2/gnue80EHpek2bJeYnMs5JT7AilFGGeh6zpROi//vKD6fQjaDN84zhYHbNrx3caYqkDQBg5b
3G9iQ6EcUKD+r+eVykYOi9Ay/o5D20UDpvGSeR7Vs+gdmCykQ0Q9ddruUQHZeet6lq9ccR5RcHQd
V8RsMFKxrzuIpOZsJvIFwjcZxrGC40hKBdM8WBgYjq9uOgCyiVASxnzXaLL9aIFKQ1YV8RHGEOSf
/PFAM+ePoVhRncbv2wAf8yqA6fsU1/0GJDpYr55VY9qXPn0Wkri+1IPSvfVtx/YlQY9xZj5H/wX4
lkUddd8ClTpyhKWzHaSzsAFlDFVVxHEh1EQ9n4mecLTX+ny8xK5HtALj4hREiI8/R0Sbxxo2irkH
ISXMxiyvsWuO3sM7+l5W0eWzJkfWOJ4pbCBCDulM7ylFuu7LwV9srznUEeOv37u1RZKVpG3AE5IR
5oxusyVdcH0dC7p4E6Vv5VbHD85iZmKKx0EvI90R9ovhpa42TeVwHSnC0e56jL6WCWdfF06OU59s
NMcUEY8SIAsoi5HJSxEy2Rsg1JYrLxkI5vz0k5hU6m/m8MWSghwX0ePlvrOsuduASAmA6mYfTzt9
uyDbQEE/zZryVqst50v4RdDakpis372JFLP2tffjk/i1GrMJ+aLEBdV3BrSHtAmTjiPbFDEPn1UN
d3aOXlV8Yq+h6CkJ5oP8C/mh2152rdCj/QldkGmFWO2/weqTy7gFMy29h2wxy+sFokb/BX+zcIAf
YrQVkMPikpHSIp+E2HrstSuIagnZQZAX/6mmvTwkeX8Wq0sADG5qJGuAjVvZoEkODA2TTuYIvKKC
IunTwHxI4HQoRidSETtzU7Ijk/FWdYPnVn8KxeFUNntg7hZFrZzGPnTasGGt+urqeZFyEc/NfrZK
4yP+wezf6jIdLbDYgDQ+N3NrEMbKsaRPmW6q53xFAZnnQccwALDHDwkBrePIKiYfBoI0Hoduh+Dh
qk5+CLnXJMET3WlZbWqYP56BV9+OrUeHmMDLLjNWd8I/NDrPnaYBnuZAV7cFk5EMr7C/OeFVZ56u
HbN47p/fPF01fW/vWcTifsDPPxoYCbzfLQzWfzLUV2Nkb6jjjVe2oru7nSu8rGyaV5kf2YT2F81o
SM1MG3KYw2ptP2sBFzuBQvtENwqpTrcPAxRml0F0pRVfzrjVsBdWINLby/tJhfSVjcxrYYFuAHeS
WQXVgOY7zxnM4pMxMmG/f9lquY7YSf4zjpwEvzprTaNXJTUDQG5T4IwZRgQCmTfXS3xDFK8sFjpx
Pxw3vzohav2txzHJk8RqN/DeJOMJ7qpP/n4JYMBd/v3QKb7TCwx8MJzPvt/9LAclsgKNYAl6QqBw
wNKoFffthipfs186HGQF0NEczmmdNmRQK+wcJQci/RXh04hs6ScRzMx8xEDbYsSbpmbaRCSv/wYn
kkyn4nUJ4RPRWJ8Zg60h6/TBry0s/FRftsqU6sIiZp1VkFAGaKGksuE2ptF+iCvSCTR9bV9I0zmI
KdZtwponjTIM2hXGGcheE12qek3ermlVW2giW+IvODjgzJ1/Dn+bCl9tJJQ4WmHYe0nm+JHP+jlz
Fac4BSoF0w9n9OBSEj57Q1sa85WWXJPGMTuc7/JDz+BYwwznN6/u+E+UbFbykFrggIxRiTFQ0e0E
xEBZKh2uGWgpCR0fL24HyrtIS5VcSBx3CjLNpBg4MJUODydL58wsC9SS3GbQBFHCXAabZhfXuOrK
64KOZ8XINZiwlrZWA7HN/M0HTCiiPao0/BvQBILCf3ZsvwDadnTy3rC7Fu8LSQHST4kTwB6kO2Lk
y6H//XyD2pSEb4TG1JxRaXzBkKB7mJT5hm+u0Jsp3Ex7W+dK5fH4E9Vg49IDdM/EspZyO1e0wMLf
zDj85Q8sN7yxAQxE/y/xRFlh8KypFIQDCHot3ZtXcY8LjlwewHW0HvvC494t/NaFuuAbkO5sNxBw
X02w55N9n0rBTSEcTd3EJYPU1HCtkT4qqjDuFEBcsp5X115kkpxGibr7xSJUcuMGcn8NEMjKA4nM
FroTgDrts9B0G4qSV8nnX6DmvZnezhW0Sy0uglOpw2ZSakqNlsOyREsCN4msUNe/BY0uRp38X9IV
KjsDD40YQ2LVHd0ST2hxNBPJ/Y2rxEIEwetHjWJ/w0pgSAcuCFWhXWTiKvuOvEeRNZcXMXeuzZ9a
v8j0d/8HRQHB6oU7RgeQ7+y3+DK4vaHmpW3BVQiY10Td28is26aTWS8kSDWMUWbqSmFdz4DJpYVr
IPKn4beNZx+9sA7vF52gOwQ2w385E80WCxoPnZgqt8Tcm6gka2kDP+No6DIQ2XC0uXYLbrAPf0Wh
qpxCNt09uC7vaz6Gxgdv5khUi20COWgRlweCYWFlDjDmT6iZ0nNTtJjOOqTEeBIpCN4cyk0ZwLIk
gpzKo6K3q3sMiMt+4cuiV07mMSHTbXA5yXH1pfZK5mDMdmOsr3JpX8zSJXVXVmCaAmzkomkLEgUP
IElspuGVwB5TEcf8fTOoGkHEE1pWR4omU+lZzLjhwOJKFUdvpMDZXoTnDpKyxLv9MP48cUMj3mit
t62rSOYMvmuCY5lxzxQ413qA0QC8Z/b/K54FdfMT3NmcNmwuStGaZzTAYJF/vTuakqUz423d4e3u
8K5++oRNc3eYqfklSu0+r3e8SJ223kUBDcHGsMM2/T2N44cHxHrxkaemComgknIzRCn0vttOmJCH
6uxPYnM20xQgYBf8b3PRTo1zK+3L3/lTIgBL9hgINnbZzPuhqyIhgxCk2R7pzdNrWiNtqJNkCdo4
W0SYHW6eeU3/qLGA8wTrSSzzbDjQkCzqqFp+VN78rq3y8NyarPkm6sSOfU6WUvY5rF7cFSyjKB1w
bY1T4NU1U78H0zyiGcF1lV3Fd91FuE0/TPmrskAbD7CpBkkxLYitQYllJBXIlV2b7i7ZnSwYOCV+
dvcXgCYQmUqHJ4QPXLl4YBxDUvzFCjW5oya+bPYyDItjrMq5kRDQkWpR2C3xVAYBGe7gchSbHE+6
VjIAKVu0n89CI1vnFAMOlqCu9e1bxMcD0T+oepJPD2ZGMvEnwUiYJYnMbzziQDQvmf246goa1rvn
1rRjRqxCxIrN6asmMRw7i3vDZipZ/R1qH5zkTH6CrOqakjt1u+UXRuEy6OLPzXtpsaDTJE2BZ8kN
1a7cbz4bvcGy4fZ9v108ZduJ6HVWPnnJBgGm5Vr1uGEiwDVn+dTIaP5txC+7/QK3OXzWsPi+7b8A
9Iu0Acu7TfZIgj34QgyfzpbQgiLbkYTf6MBbH9WW0OLBRsPGhrEKm81QJWqHXut71xSG6BssZIZr
I9cyK/yHgHVxypHN3VIPC8SZQN4ydSOB6HoWz3++130sW8pXVtdVX7GOIPAUwjIiCZ0wTWHnirAX
n/AwCG3XghxRa6DoHeJZMlOfqYMbamXdhWRvDTWPQXiCbvmH9Tjsp+LUbcZ1oMC+y7A77p23/ecw
s/88piuvZ7MltEr3IUWIzgPAsEYBtHEPIc27LG0TCJYLGhTGAp6apZAicTs1EtLF4BwvM/L2kxOn
GpaULrZwXxMWID45WRkQtr2MhgMcRVHAVJkwWB/V/2Lh8Zc4T4YdVRgAoNeB1SVn6MJz3gcuRAHQ
oFdKo1/xbSRVKlDrEpFtJAhb8dnl82M7DN8lbj3kUY2RX3HIcy/5PQwvUfCRzbhZifBFIadDd9hs
6f66R+eZe4azFVxs2imJYn2SygEqCxf8Lc4GJonhw/yQI/3IjYqnRYUlc5wDebIE87W2JNrAob72
c42MEdF4wuXxsKSUJcus73YWhHOmN85GzgL0bxg8rzO4TwbGMH//wkbrmv03g38Q+dxjZU0+i9Rj
sjo9FrpRSRp/c5wkZnEKkdxK1azXGgpQGH38oRBEOBStbCwlo6N9Zwi7xryNfFzZ60mWFW+4y/Oj
EDuHIBGlRkKA9dexcAycwC4OJ3o7GfkhMV8CxxHkwgTXeXLLYf8l1xiVWXGbH4eFc0JPwfyQHZXw
Do29NvRXpVXA3Gi4P5FMaIYhklJI/KMQQTt9HpF2P34letWrTFTuNVXj/YR0gXseR4dMjk9mz8gs
CDhONV4BHJ1qdWk02Dh/w/p4hpAxRHGSfZ2QcaIZvTRkpV+jfSDytIHqzjy2wEMy5aIxUgu3Vso4
wCzb8HdA2kEs8J7kaGY/O84mXy55CuG64G8ecihNKhE33zEEEM6ST0WhEKY4nqBBaQXlmQBDAQ1N
ZBrDmBpXu5Hh5Padl+Vuqcuda+AKVyc7FY4C+fu6wgAH13DMYHE2rHw/PfF/r0XuwFLH1wsS7Naj
TI/pEFOMARqQJvYsmqPd+pSyrh+/fWjgJc9uddqHfWRXYSNN2KiYGBvXd4eozltkH/Xdf7TAlkZf
5jML/9ROY/Q1Csp9Iac7tCmvPsGQnmvdumwS3WkJ3P0FKv2EqjjOTMKm7NcZ8eYA+sI42XUHBxO2
UbDd052J8reNv04nEDlunOwm7/ZCMETdawioRZy56Grez+Kvx7QkWofFs1leFEUebxTyPPI/t0GB
sWrLcuJWEVzv+3J60tzWBE2nZ8ZGAYD+Hi+g0uvquPjPE3Z75ffRLqyf49ScQwpRLpRbSGE/acZB
CoSXqBnswababj9STlziqykPA8aWiUZ8w3NReut3OElii2K24bJSDz5img6qRZR9a0W+Dd2YF4e2
BovPozW0YaGDvRrrhsFVjKljjShNH+5D5xiKHl6kURASGrimheik2d2DRHQCDiyjQOFCBzz/MVNX
aeCPzNhDuyailZTh0pdQr85UW/DSd5BzVjKf1/xc6PQg7ytL8SeJxTp+l8IzuwzsDZg4Kc40pSFJ
FV5MGgjbBNL+Ja8FPBCa6BGuHy7rA0OT22iJ1Zpt45y1FkPLVL6CkVRrE8wUv4kcvqDob3F37Wc5
+UNt07jn879uJizGbZRjRc8/vDBtpgaSk8Wx/uh7u290RqBpoVj8N8n82dJZ71NOEjyUc0t10enC
zc+igBk7RK1W6WY8wlJHvEsHaVVRYGO4RNkqPRb/ygZx5Rw6TcwKJMk8rC2UUyJkvNb0KMTsRYa6
8Bfhq0pyHGGi/QTEVHDdni58ChASxleCOM7UI2Uf/v/LCzVoYD0W7QfCnUApBTi/lrYoQWhbz5ai
JSvdvIVRt2gGDMByKPp6szLuEVMCohJmTI3RpmFlI2tuI4utp9ZEUO2Kw/cvLMcZUYTDV+B7ZHDe
YT4v/JyWM11/Y/aF/3mcLRuI1YXOn4Tum/DmMLw9AE8s5DktD/9FaQHVL6yZf3lYjbzUU1vasMit
hHVI5sS6DZ02lr9rohjNtrUFkHN3SnpzIB4kRi7W9y8cD10pXgOPTSav5BjX41/RoLGhdsNoYNnz
rdfqOmhPhJ+EQI6145Kc6Kt42M463E4aGaGTbYcxzOzrLkrbTdQXuoRIWgyZVkB9OMzcMg8gcqDC
j6TiGbSMdaqidrBPqzsOUU8VCosamNBTP3SfOuLQa97889c17r2KP2124D9zBOOl7qLdTnRi7Lb4
fq471sjtpxwv0BUgPuB5xajshp5pqYEbWxNIZi+yOMd68ZRtm3DxsgjahY1jEplNqZBifBFI+cyY
HI/HnMCkRXQWt2kmffTHM1s3J0mYOjzuhU8a/5YwoLLJPGsvPqf/TY48SQQz3CNTwdESk71dvB1V
IeeCzHElmhgS74U4POzFkgTF+6pXlkwkHJMasDZznA979kPykkE9BAOB5z/S92ODbM5bmeqqclLs
Sbq8tqESxQOmSU5Mo32apCN0nGuchujVBkF7tCk7VB+Vt6na1vkb3K2GghYQnyB8hSYnw5OxhLfM
i+9Tmm6f2w0PkEaDJVk5/mioKgPW8Z7WFxr98LkXzIA1RjlAiDZJ1G3JEUdlhJOVBqhSfu3TmFip
7U2hHEGmJfQkrsdR/2EljX1V3WJVAD6Uf/3i36aXwm8hTn36fDcQMYh/3J+t0xNFkllNxNEezu9N
Shh5RkdGtuJXDGhv/wXjRezJCE7HqAEthsVC+DKIMbKJHdxB67qVn0yIRIPqOvAym4gY+4ocapcG
7nRW0JmxLYbf8N9kqFIXRvKMt2BWsaUSxwZdkg2rQpSRQ+KtfVO97ghoC5kXdQOtPbTziNOawdPC
DRPryCy0uDPdHO8L88TxYQCMnCXGOzZ4NOQsHdBuwIas7g/VE6W4u+cqOlca1ydx/ZHhmBLdZTBZ
fKRgp3cWBW1BCS4BUaOcKrpeUzl4IyXWmSr9wzZeZMpvbua3ROz7ALjeKUHIqofpNefKSgLJlMZz
qjJTkfVJy7q7iPY2MKTedZj7KV98GkpNrfOTi2omlyxKErsrq2GvbbkuEUNW3iFyH8iH+f7K9bN1
7l7CtykfwpgT3/19ZUygQY2HFdqKnSQuioa3oehciOlXhstPO3YiTlIs3K1Z56HL2I54tKD/yJiD
kK1OIc2ltiEdcwY0t2+ldGPLpUWg95s3ilwD0o2TDe8aGh/CBNplD/G9t1anVmXRGlOe1U4WjJMu
hl1wz/Nb0vbLJOydaLJAQLEgj2t2fyEzCzJNKQrNTIZ4dhlQsu22rAtyLNpCN+gE/iD1+m++VwyG
f0Ex89PoiY4bLF3h11OpZspSSpVKXJQnGi4YGC4dXHtFzpBBBN0rnqp8d+PfHZ6vw9hQmHO9a1Xa
DJEuodDdS4Jc5KbLbAk61q8o8C44rtNkkYQ8TqBBdYKuDY5XetQRJMR5Q9keyMCN32NS1ChbSO4Z
EiHD3CaCyynFDtbCkVQg3nJN7oXsbHkJCQhEvNLY3wrn5H1fui3Yn6bl0l8Y+ISUDQA538/0FwJA
/Nrr2Ba+8KgkUGhmrBvu8HAjQPgR9J8XT++2h9YQ1/YnLTWwxtMYNQVJnRSNH7dmX0q+KfCvJ3Hm
+is959F6wprhv3O3602dXPeg3+eCT5ow/R7AIY2OlIEf7OAGtl0it5XMcm5gvhzEc+yo34Bim3JV
AotOo2iX0Bf0zHh14fbUoEBJgVd5l+gx3EsCHZhBTTDfCYRLyT4K4t9wmFvXow+033Ezd/shQ6T0
ISUu/oaZizYHHVHXpqP/hrtFCUGp3fym9wff2EXWdODhvt1hCSR8fer0KQWLGajZuQvhTlrADETR
Y6PDrGz6KTezJ+sKmYPwzEp5K1dJ55nT5wzkJbc1LHCV1RJDsEBJgkokeNCGSknqgKa/vFbgx4am
s9oIThRhOsct3WFbE9AQchkfuG66tnsnWMUc4+dI8z1NmzpN83Pdqd4VFny2N3CLUebadrbAVauw
myRmNQ+ZJvyccNd7F878m6H/Z8zVXMXRZIfwFV9aE3MBJHAzOK5CPQNzYruXqNMMgK5EsxIgJIyN
kKT27Gas3qof6upypNxjBTaGgyBCWpZsC8Qy/aatruNhL2uAtJVUHccLSvqkkJYFBc4TGiTypGzx
AJRosN7+Clnp6ZN3p4XIq0nNi7n9lCOfm2AondENTpxDlPWUvIAUMbELmmlOe7/4NWmN8vyRQ/cb
2D+qtY/Yi38oA5o/e5iUkjW3EnrUUj7tPuQ8r4ZU3eYeLIvkR3wNwfUPCL84BWJ+6a0voqYnU5MT
MfxwkTscN1ZVTreNnL/pXln3yQOaw8KMttxoJ1rDKujDSNS2bBTpDyDsimX8/odsVQBtbTvfoofT
qhYLGwfulBtPJiFRwhEWX+tdmCsr//Iyvi+PbgWvMDhCqdkBW3aTrwTGQSQBpJhcxL665lL3aWvo
qNFUI0RBz4JZk48jvuWa9HKIPw+3I7ZyltrNK6xMRub/3wdthPGUQxG/F561RpvoW1L1Dh+Q320U
tGyltv9zPKB6/PfcFoBGM+R6n7RX5cjVOLY1uWrunT3xvxnT0ocYD2UYAjbaPX7QWWW3Py26RoUE
681EqQ4LpkljE7PYoTHUzPJjA/81MzmcDBjgalNoV6l8OEW+XFM2QPvuCXqt/R2Y4hOalULqhMOW
tD5i5w3R/BQnzRO0nsVbqrzCQBtVAKOd3prEVUmpHQRw+2OXqcHWPDjSfADV2TqfXXW2Anv+GJIi
uu8hJCC2K7UNAQWO98oajp1ljJLNxYDgJ0JbOfJPgQfrUBMh6qBTDW9PphoJFpLqe5xRCe8bhCM/
VyJSyx4DS2qVuUzTt7RKeWvsHDt+FMyAxeLVDRaE2rxA6U1yuRoBbrqTD41Y9ZbZls+0j89Abfyd
4S6anWPRrTD2Jtxt6qMWVipTQwes1S/wf2RDTPb3vqqHLZFRC2Hs2OweuwfOqZeFfgkcvyXw2Wnn
Bmp+S+rnIdYvSVwnaOIKR9lppIDLoOzEbGgPD2dDK8XbkWvHkP6To7ERysIiey+wR0CjhhcFDu85
lBLtFBzlxpzu71X1GJH1DYZ7ikr9VpHT3tLVNUQyNKUQCxLrqPux25LYs5zql5IFwNTFD2J0VZee
iGuBJv0hyEDn9I6yHb/hQgPTeQWf2sA/E7yCMcaao9IycYQ0Nb6h5Om4EDgfBjM3/JJvl9mlt43z
yeHNGZhXE+19h8cBvdTBXeGWPph+98v8RtJc2oFBAUWAwa2EROPG7D3jniLARVKZwR4wSTHSxBS2
v/TPOgy5Q/B8Z1Ii7maAV72UYYPG7wc1nOvSsPecw2AB1OVzZMnJ51GorzPvHLQMJ9XihgJ183X1
UZm9QegQWShSUUVC+Nh12m0Ds2oDpeYYHW0a9zqYqoBp/l3+sGi1XWhwt68saedN2RGDgIt2P6Ec
8HTcpsQlFG0uYEuRvJtt+w+zjGvegS7TmFmYewICUsLzm76vLtDNox4A5/uiuCEasnZ5M2d2tOou
1NfY/NnEaBLm4vmsjTnaYISsId+mGEZnxfvsGgONfyw85erso8s4INjX2XqrDuaM75wmZYmNeHip
rvxkFoVX5bhUXycicCPffoepEuxd9jqQLM5Xo0iqMPwvWnCw6ZOCLKVH5yrRY/GImL+HixU2HQH3
621R5ZSPm7IBcBovMyzL1sa6fB5eRgKZT02gQpkb6kXydJf9MOodCT/v1asOyUlRcZJKG5yrxJFz
nxt7no8CNdNUDWCWCf1va+gNtWgpsPaehovXKHNdHH7RkicEOx6lyITWldmCug/ly7ICN83MFmVx
cOXnBnckexgBQvsj0MtjunIaP1gsp9sSdCgvFsB77Va0Z1sBeDjI083xnjlTaKjdJKTxnFLGBLpK
8ejZp6OyhQZrCeH019ArZfe5IProQmOcOQtZUv5VXeuOEmQJ7IybXBGOKs9i9U2rAaHp5OgB65Wq
xJ1Rx30K3vq5Jd12/g0jbjKaJq4pTvcV6t9wjwQdbIgUyXuK0TW7E2hvedHn1dqxTKzrCgag9De6
asJifldEI1AaDBjhPcwDnkEQtOxpGH9AhBh0aezhzFGMQgAWAsOxjxsw1Ym408V6XX1lW1AvbBkO
oQd+/Qwkg1qEAojlvT7e5u1yEwv6NJrTsrY5L9xmc+jd6pzBmcNmT152cHwkECRl//5e4VTrv9lv
dpKYy1wna4E6QyiIi/vbXXzCAaepsxSax7ZKvEQ5AoHimkuOxIk4jnyW26/pakmK25tQyLYbNwnh
Ypokr3chlW1aCwRWI9kIk5FcyADrkSFIKOvatVUJX6y2l1Bcd2MDIcQZbwHdo7VnlxIjf9JUWDWP
h5UAO/oSNz6gyn1bGt7GR5UjApqPmMXlUVIpiq17PHqaEbdHO2Y9um4eyGDF/O0rFOaLH+tqU6rH
sq03MC5BPjNtjzqHf56xtGHbzq5wSi45TWL0XvST7jQpI9hl2/Zx9Z9FP+DSRAGIq4zrZ9MuVzBS
l2Hs0L0dSXvwRhbA9Nw3+YLkmzSlEXnPLRsC20dk1w+tqBAx1PzOTwd8ZCEvCCVXs67S4HQoTteq
lpPP2Vr9kJkfhXbO9pzNHyP0jLUQccnkhahAlHwbvL0k3NI70LQV9bzCED1q1Zo3XEfkIfbrJ/pO
ZKpubN6dxuD7IwehFIVz5Ia06WKsS74gJmqo5ikFulWH5b9UZDyJEoOlaJvc86frI30RF58Fbuj/
mmdXpO8OEgpUgfvCWk0jOJBG1wO5qKqUa9INNu+0yyvm17N3ctUqaPKlTHjUWLuFf3xDoUiHsH2U
LNhe4yNNtKoI8VHsIdI9H7dHpDil/QGKQWEQfxw9kdOgUQkgaT30abLpqgObxPgWW7zH2iwFP7ti
1Uyj0WM4ZqKELhzzmyV7i705RyRBs8U9TF8xIuni2PBNmlk5TrMPnLkHDW3Jzd6GhrRCeARSOv70
zLEZhZ18J6I7UwDi/TlkoYJXjwGG9nzy6zrWIiQlYAYj0vmNdO4Px/YlGxh4cC0S2409MqwHKwkw
uCY0LletKaykH5rnDenR3wsnC3+m5UGSWyljWePhn+xL37fxl1OorbtNC4swWsg2b0PoHeir73V7
wW/hGMITsljG1ne2EKcZGpEvyQSlPTO9UoqbegcgcV8yUaHWOWOmTuJt1J5JVjtfyPlhCtzalFtO
Rn8rCrPNCXITUaMODV2HEalqOg8OEZmhkuWQFaxyilLp81TLzY3Ku2cMcx/AECWIfsyGozwLpdpj
dHN5rsrQRHZq9flCumUJ3xwoVf9TgnuY67IppnTsOfDr6H/J5qscZ8s/2HYb0PIzPdpVCCdAc0Eb
iK4EHPh6ITJZAet/v0PCjhzEzvLel2VaaMRBGG35XMFRD2+W2qBSE6quPby7xOqVil2xd5WsCQpR
Pmncne4xACJSLYZ2EUMnz0RIJmoRXH6CV6e4W7coxoGsvNECXBOAMrWtlBUhZkf7aQNUR2MxFknC
u19CIeDiFx+oGltM7DzQ/qO5cC9oaAptHGUGuJd+Eq5wyEHHVl3ppxjzH+j67vZcpdRK8TcZoYdF
y5DzJp7LOKEJx3KidRciryo3qWBb51eVoBqAYFy+/zCLQZtzbdkUz3hy0s945rdgYb7KhTSE1a9b
6EtiTTbdmvYUeeANS1rm1Pe33KHMiS7oYqzM0X1GegD95uhZg8WV2o+/bjpAAspOwZcsetppgtpN
I9uu1KrLsITHKGLLDo79S1wTty3QM5L5Np5WCjR24BhSb5Y+x/Q9QhS9cjiMo570/O+lQpPRdnDi
wgMty2Rblp7QC1vPN1LN+pL4uYWZ+8q/w8yvH7+uUYr2LXe6MiHtPCWwOG5TbbADB6is+TlH4IEB
Cgk+YrkO42Ojte5sgQ0V1XDEp0LVScAIPNrJdcqH6aZf2Vv3g6piz0NjcK/SEZ/BQsPY1IJOszCv
d9JQ2vLVrg9ALmcnVRq6LVkEwiengFIVUrYYvfzHi5MdV0eqw9wEkLjk/LbEarryHBeubw13BNpv
7CvwjqBso4oZydMnGK6pqHoTO3J4/xeo286iGYPSSO0eIcwe2Af2TCpADdZWcMSL15IM3W0++M6/
A/Y+0IJ6YbeAfF8C60zuhJadMd34mSyhPPreUqKLmetncIE5A51F7HYiRbb16UkqSVLXM2NhAo03
ujhRLqEIDiEuuKwtPXQsJZSjhRZYYdoSwWaoyeBQUxf7sUweYSnGGSB62YNThH/EmK1yCffAbZE5
Zr1DV1ewyu7PHDWPOKsyLGMdoA3cbmdwiBss6s1qXlY9Iqdgmk9OcXC92eh9GUthy/jACfw3nkJt
1HazNFVzB7l9Ae24r006Aq7ykzoQZJfc3cNBErwkNJDKh9S86es3csLBRKmU2RnsOtx5AeZ9kVvF
t3tPz78BWnR52eyZg3Kr2MHoA93244Qygn4M5wnWFYsOfkY9qUPkNMqFVhpUS4pw1x8Lpbt3bKSe
iujafSOGeq90oxGSIgslV7uQi/uZwTpUCrFgKt8yJBNrxtGwvc09/XlQE3bc9QO1EADCcpQsI28s
5a5doQOJa2fm7fUmGrBnNqwGLivjOM33cvev93bL7ujmaIaGrchadoBtj28SRFfbrzKq73qpbnPb
PoDN/qhKokm7kWEfv8k0x9lsKk5ct1jczRyehLfFDN472QzGFuiugVP3nrpwZeMXrRlUFmwEHKyo
jaYxeyG1zRdnHPjuIofOn0QE98bA5KSSTsqfGwOHBR4gT9+pfCO9XPPtKKcSBx03ON8v1m1G0Jcr
LIOFFIDT0S5NKi0b60iglNdoSTVs6C/uK32WYrPNyUSuAwcn804VcZx0EIFV+kDro3MOrLrG2His
D9wen6qim/1q5YoJaCLxxMZ9VTYk7rOi9IPpJFZ3B5TfqaUsIvOcyvmpUvZ6GQVVEllMTYCGymiS
4lQsrOHgBFEpMXhqkTn0k8uLM/2yq7jdrRBUdOD5wRfcuU5sWXFrJIoMClqrFywtgyCH5AHW/Mhq
dQDa5ltsuIdKfTsHfXRu2rjIS9E5AntZZStjc2ihpfSKogdHs6NHGVc4IsqGEXedH659CsgnwTy6
g+IB/7H2HV0c8sa0Gof1j5cyLc+Ojc2Ph7HqS1NEL5VG+8k2DwRZBYoTIsjmm2I4oSfnf6PvyVVn
CRjRZyfwsrIc135JigGUV/mfWOzKIgSXC3a38fENytChZBNtr9oH13jbWpB2xBXPU91jZRwhEWew
Lbi8zq2rttPBhSQwdUvTl/15kPe+0VxkcavTDIb/DtAYfElOtd5NpuRuNvYrRkgHIA3/c/kVP4w8
C1LtDzCBjK5LUySkeEioAvBFqmuixwjOYHVZz6SC5M0dXqZIf1KhmEGdffJiLH01Tr+3ggEEpfwN
y5CKKW0Qe37m93T8/PGKk/CMKWptxLRwReFsKH4jgSKU6s1UTb0m2qOIBP2/ba031g5LprRwxdau
5DLNdkz6Thtiwgif5MQ1ckZ+EuK9R4BFZ2vm5PsDKWKAkQ0vPw4YU35blxJY4QUfuMGomjHS0Swy
rRv/dsdUeLmI3mh2T+peNV/Rbkfnfg/wh8OPjLO9KljpRN/1HrkUqca88VLO/ZUaWCCfXVtOJx7X
UutFiwnzWuRb/I9nXoyTeiW56lUaA0RxeCzVkpuP/ggGjHp2kYGhCKYxAjsMaRABfFmQOoGN3Ni6
p3CeqP5thCpwVhvTICOd546hlMOKHEHqS+bmmYHscpPAxAq6XjjzMh5nlfPzKXbWeMSvadeO4w/l
aHZDkKJBpgRfdFZXwHO8WHa5rMdR+mKcLeudfpVccJqekb+Hx4t9sQlNJCfCr2gPTIgMX5oRgM8d
Bje6FlUvrzP87aOgChkP/FsPy2CDKibPe3NUfoVXCgOeFZgzsJuOlkHyPHmwf+HzX6Kd9HEeXIig
hEiuVncBXXCD3raePMNcGGsF7yVsmSu5sziZg7cJy256wjeh10I/SDabzPP7C+Xb4MIHyxuFWTaN
wBVyrxTJeREHkgHL2OuA5IC2KEqNyViaqT4qQsEwhHQmhaTNThXK0NOmM/XJTSxI9+H6HOUtAN5G
za6r+taBtsnPdTkWfTLdzEAp6Xq2VmeDabSFRdlGAl7VULZAKl+w9v2oVDas+r8gUz48JG3eKJFD
KzF0Ytrssi/TNmkhPEzif//sQPOLuEE434s0IFWF9N9T/QE6YzXSBb4m7pP75By5lA0hyIjRGDDY
X8SlbiRFfPyM2lSIwv8bm0Cv7YEey2Ek0QvtyZ7liZn8esL6rN1vmjOwr1rKVFem1xcjoOFZtOIb
7VCik6PwiQqZMnXIAE4V80FC3OkElZMwAgqoYrEl+4KXVY8qaJ/frhgvFPC0t56EsplN3gOuCcGZ
KkfiekuiP14UVXTkrEksnVKhAKkDyYxIdN1Xv8M3YHof1cZwEp6r73Dk/+70EzYDZZkFp4zGtTZs
JJWQUOlNn0HTHZjEq9oG+DRmqsiEjGBavO7M79ea/6KWBALIeg/WNbC5y9xCveDojtP94+VVFSxc
r7VM/7Wb1as26P8XcM9E7nqatlh4v9w3y/Gylutbx/g+XARPfxVZd6zC8E+wxQYbBnhB1f44Q+EP
H+yojTNQ6PTOsbgx6wN4pdhlS8vZ1YWBqSMebCva+zD5MayTAA46L2d8e88eXDULSIjCYul2vHFE
7/67TdAzKTVDIMeCBykNmUzLluELbAjVSbH3abXXZPSA8NKT2Scrb3O59wxlfEeC4Ukp4Ka1GgaN
365xc41rqeSwyKKkA906dI32gSWbkcvVLOnzgEiZQVnCPbSA1U4ljoYsmILPDA8G/qbG1e3bDECe
yAanySKHJ8X9ZEQVH/dvy5FcxrskGA+WI5QjGCCWfN8PgjhRqWYWIa95HKi4mTtUqlZjEMdWaSsH
1pnn/HAVc2exqRzXp5G8fMEyt8fREQXQaPnVFmL+rdxypOJWbyATFVNsxf4seCImpduXMWINihQn
+SEUtxo0+bkbrAJE07gQ1ACBambW5m2miDuGE240jZ/RBdrlD4vxiTQKqLlWlGOzhtXcCEp5TpVh
KzQj2QTUP+J6Y3FWjPyZCNM3pgg4IlGrN0imw8VvWTtY84fqPbTmy6WYTp7H+ZAUzS+zLldSI/zu
wSu2xKd4+Lsa0EGF2xTm80sLCcWmdtLX5t4Aj7H0M1PlfP2ZJXtsyQR6pge8WQl/8s0104uGgWLc
iLGQ4dZdlajxoDjl2grNfzcpLjWRT/bBSOtweSC/tBNx/euzl8gFtpIMdFScy3QQOxwa+w55hSc4
42vcBkNCdCNXTw4Pme6OFjhqg12G12P+LEJmTvj4x3KNhU5ydCV3t0eFgooPSgb5sC7mNdztj0HE
qjJC5QWkifGW8EJt9Jkw1mNKniwWWM1LA2VsrhfCcHNHbteXCM1f8huRYFbc/4+iUE4ez9w4ePzm
BVUE5JOOl+SdtNGOWmVcUj7B6F7jvuLOfaPU5C6HbcD87/7eiLLNENXo+CXUiTGeKt56Y/aySkLe
XQ0nOVq+/bUlGl76GbjTJgz1CW+4Uvyt1F76fD35FuOG8aePI19ts1+9e88W11C3htAabCgprY6M
tXH8N1SPgFqH2u7j8gcGM+qzRymQIofp3b0CiCnUp71vTo8t1nk4cSS+/7hchTk/p5PRASyHkvAa
UndNUTkl1jlQ391MfN2IJGKCUNxznWlnWJXu0qsXXVIHO/+SFLP3VyPA0y2KEn7/yUrQCFBBli7V
lEhrS0Snh/2IjdlMQwp+udMvGzpjbJYXYJ7EMj1NFS7rZX4NVljFa7x2JZh5ykPLPdMef6wAc3xF
Hiq2+g/NP0oOYduAEErlYJ5cu26nNfpR/bilNvD6ZzGtpDT377cagoCkjY+GzxCKCyYaH8x5xy6q
zpL2gd+YWj+XB4cHeLzQ2EU4FI7lMIDxznK/iwEsXxNG6h+sc0WPVKjKl6So77IftNX0UVEUEFJ8
Onkud1O+IqqycOCJdCGXCtOQblwYdB7pnsbt/HlpMvDE3unYzdtOzlKqp0mk0kKBSIsXdchs26bs
u4Cfl89VNHAnfONrIEuij9igKFgb6lxA+dg4K8UTmzmc4MiSYFfa/FCbhq1AFS7TgQy3RqDLKRJc
N4KIequ/lP4bVGUqdgl144SlWOywrd1i//rjDn6A
`protect end_protected

