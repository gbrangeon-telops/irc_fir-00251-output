

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WOJX5Fv2S0CzprysR8KMEndET58Nnshq5G41sUF8nyr23cEOOYS3xFWHzDNrh0BglAkKcA2/EcsL
0Mi0zP+UFQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Gc0ueCwDN9OX/N8ZykP2NxXOhHr0aqi823TAFhXP2T3sZajOBosaRN5Om/T8R3LfwK7+baNKGGz+
UJk1ogy8JwdYWmJV85/JpyrrDFtvClJsQxdfCiEg0IVlJhvJlhs6FCZi5Rj8qwlvbn+/sc8hT0BX
IEC/9Hv+yH9f2HZIeiw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gOAtaUsYvJmoKivS2pd7kBeODY1Q4VX+agLZ2/SaxV/BkQgGuuCLHYg9eGdXBmjxTqXO35IrXGnw
8lzEMm8YS53SBgfLbyNKtLJ5Qej5jTli3Hhz2BXRqoQonahfpMOh6WT/32Mi5HxamPl3+Ad8Dyj3
AbqGosJ8LBJRb65Babsp/E0dGGngj0nJjmmY8NHpqNTG489434uBxC5ykK4ltOheXkVJtXSHoR2s
c+RXEPDO94CZYlHnY9b3pUqLafSVqXTeYuw//0PIJQNmrXYuvkdozgm129vQnlKXVGzYsK5DUlRz
Q+VO09C3aal1Ga70326sWIG6XdhCFEnAfQoucQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3INKfUgfMTydNk3PjPUP24H0r2p1C85cOfDxce4LgEKtine/HDrFDahWRWORtm3mNUVaknW/GXSC
5KErdi7NyQ5+CFdf2MMmaC9h7nGYKW8O4nbf09hLlm3blRBSd2i3h46PihYy7iaS3Q+Z7JKvWuiD
J79EKDKw4Kqn3mmg3iQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YHV/PdEXZA1kC+N7hsk5uDSJPgfJRc2Sgeu6l1dsNtZhWFmXeBe9vCszID1P11I6wOICxCc/uQgT
A2JL79m9I3kuY9Ji47hSGH6+xG4kfTKsYaTVdl+16SjuG/YaIhBwQfN13p/8IGQ6FysnYNYR5siA
+0Lm6CwAYBXVRwsuIA3R9dSPKgq+Sbk3MQCuaqKXbxHiA5oAAI2R3Gz78f9hrvy4Cj5P6dJ+TbkJ
j9bOdpZE4W6tXHasCVI4EqJlfqQQ48uWK076fFPDGpd19w+K6NBgkvxxlXDC1t90ZvbdFgDD30L/
SOFjS0BafCCf2aKaRk8VIdeBs9pr4wj9gMwZYw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12496)
`protect data_block
DUksb0OhCQnFdtJo44D4mbymtbIClEDKVbnpwN8Y3wPzdEgfHqzz80BWyzC+HgwyR8ZKWwPHCZOk
IGgBQnfarmeGuZgmP4sRujifLitPNDsgirDhZ6QWY+YwUICEbREa4H3MXgI/YtE+k9NAxS9wNwHj
AcYA3mbodAQMnPBotGAVNdZI8uPn0cLMfzIsE23CLyvWd1MWGk91KjJHgCXw4nPMyBMtZcVIJX51
vrdeAXPtmiSu6JIc7Hnqr3HJs1Y9s0b39fdIgLRIZJrHzwYAhKFq/x91uLT8ORyDnaQIf3x4gsOY
+IvmHgDndtm4fNNYm7+p/kOUNHGHR61C690Bn9BZU6wiQgSokNkypjwCNQkII8g6G3+wn9p6kZo8
l6EROIhRUlcCna+7HpITe1DEpFXrmvLyU1j+rLz2GjjtnaSab80vd981Xrb3/UTd2c5NZ/HTDTg1
OwHDbW2N4pYjioI71QN1+z4lidDpJnAn9pPgx5S6ia1L5iduq8qcmqHOL4zFnBiMy1f/B4dteSQH
AYFSiTo96SKPhO/5nOEv2jkMKwQq0SsLfEFCscRBspS9lliss7OHTGI/a1COsvfIu8ixpKKTn6DV
pVa7FDVWs88S9cLEgm4fSn6p4zL1OO59+Dk9t2OrGrejEkRGFyDbmcZszEL8LtUPaQfqkytm+Sm4
q08bMEb7bMiMdezyWm5EdyvLqt79eM4fkackYKj6/MLH5xPzS2MOtOsohpPbYILPYeT0mRllJ5oR
J7U5PNSWkzjEz0Zt9ldEHtU/Ye16veIQYzPohGH8FqZYluJCL69PJ9RyC8Vw1DgiKol4kIpY95nR
3E8UUC+ZEcPFGC1fk0m3mvX7VFj9heif3yIi3rpubdKtjsuzHbavOZI/J2+Bv0t9szpbysXvcp8s
IYnKrxhBRL8pxJf2q9gv7qa4lws4esS767KTWLaKZ7XrY2ue9lFQdfXLCX35xbtBG06g4mtxjvCi
1bVBPRHbdoPwL9fKP6wwJzJXJbYRMTPH+vUBaeYsWMefXCyOtcWBbw3FPhlSns/1mEidD1MlRXtX
D7QOnkqtiZ/TPyFQfFdtMRgGq4ALFxkGb4tDFODBHS5DMxdmJwS3MqnS6wfDv2qFCTjdT/5rUuKL
ak23YDyXfqo7NvbFY20NCfyJttE52P/2VbMuvG4DiIYp2JVohNzqJNksJf/zsK7J4Xqe+m3ijMP2
A1XJ81mz01lgvsp8nPQcMQXIDmz1xE3R8g0zTwqEg9IhxZgVJeAx0bqVUzdQmos/kPzPdAwQMJDx
y9f3578sdcukR0wNSusjqcU7Xe7U1eFznGoB9dDf9HVHPVyOj2MJ9DNf+de/9px4A6D7TSkmsM29
kYTv/JH2a6gdle9aHwGGfFVjLRm9VBynyBZbM2SaXXek5y0Map0geK26j7p0/REL92wfz3aWdBmS
h6tFtOhMH2Ef3YIUhUmjzcSGmJyQtlI1jMHCOkABC14SRVvIDUi/tmy0dG5UyisRLuEcISUXo8oD
9WaaDVD+m8jUpa3Kz71qbEO2bXJJ50VbZzl76yL4Jo2N1GG887mhncWl8Ci6M+JPEAgKqwvpRnUq
TMiyUUM2DodQtRNGSz/+J6fIfxpU08halSkxzksZCRfQa9azGrtPQqdDtDcUvL33i/8UtPT+WCBb
rDKTiRxtPJf0vRai5fx4zpbILxcfg3GfBI9nQkJgLmBiXGUaKtJS7R6BkNrJ0WqKqO+o+PUTqtQz
+vHG5bV/Y1B5KtyjxSVoL1kuj6vLffWYmKjRRyTuuMN6nnzw6eHOSywoiIdSaQdK97kmGzY0/rli
a+mNIrH86GyAYJHYYLXL+w+TW4dL7L/fsQZeEBktapRTw70T52E5HDQ/MECddVecZFJspeEXlbVn
aBk4psn5vY/6oqUbMEGv5WXK3rx1nho+xUsjMhU12lFRQcgFHW9ymNU5/rhHTs3mwQyIDS1jIFq5
n93iLDGs7TyNLi7tp318P58Z2/e/1BvaD/ocZcuhqcBUMzItZ7KsKud7ZXg44WL5utORnjyk2EzH
liX24+AWLuUb3p0GH8fiPqPYs6JeQ4SOhPnj6vnW1VK7umnA1cGe2Kkf5YWmGT+328cYd9pXHe2k
DVEPGdM4Egzrb8zxSmmWmrijTM72i36jEyDDt9QyhBxEiMWHA51UYo4+2/UugMF0EaP4L0m3hdbR
KbDA/8Z3843gdXo3oquR48wom0yX9oclE4aQuVQb6QlpvUFoRVW+tViARtIPR9PQNZDshEMFZcGx
66IvVhRU3n93erKa6B9NUDF5Ud+Hj0PlIrN08jIE7wA/wlHmAsCB0kLRotSYxG8SFhyoZcAN2g71
QZ+hg+4d3upOz2V1vvBVZpYvME0K01MNHFwz3udViMMbh3Qkr2BtenEloZbyAyjXBUbleAUqFzac
e02TmagE/0+vDyyWFt5g4UuXa94AJBM4c7inpgtBqVEKpAn7Impn70g7zdR6uldlbjbnLIfuSSDA
5wKVvs56tJI/bPA3XWl/sXx8U9G6N/22bipr7STpP5nuqXEoUSjP74uNm8fxmWZ/b6n4R6t7pLH/
bmH2XIxIy4SBY1yWXLtlD7h7MnsIbr0D/Gjl0a9707ft53UjaUewji5TPhT2u2BG2G6AwVCQdvBj
CaKR2BYXsJoe4O1z6ODEhYU0W7oS6N4KnATE2UQjqLwh6QjC36WnN1eKYiQBSFBhlpWogVksJLUs
Xvz8+s1/8Ui9HCnGI72lWwtelWt8M8Andj3jBAQtJy7xrXDS1L7RUUiu+vE2MeRcgjeShQQH+s+/
EpM7i/f08Zaa5eRxCIMC6jDkpR/CksAqWtas/z5IpuwAvtkFJPO3aJvljrDRBhNSJta5jpgSk3/h
Z5tTD4QZfUV7zN3+wFTra5mFh5G6AYMx5g58eH+o4bXw0ILNjMvLd/OBpvpLuGBBfgqdjOJyZBeD
YGsQv8ogm2hey6v1q1mmW9+xTQV5/KXEcjgHdOpN0uilcO0NexIn0dZdMX1bops5aRHeBqMyK0lY
Fk3tmrfxnYNg75bMXtEUKi/8KBTOVgOawxIG1Z8khuFS5uCu95Dzy45LYV/sOPgUx0h6l8KKIJWm
1xPBAXcgoNDJQKXD0fhM/oCIr27QvMM2qc2aZ+08eAKmRGPtGYoja1oRJKpq0DHlvReFz0kFcnhH
UH8qNmUOw2ZK79kNs71Lv4h+ulWR0JlClyGia3K8/VKjXXhvUwVzy6yCS/Rdn2sIg8J8l/L/y090
8rfUPEEnad9tUF7gQELGjZp1lgBeLUHzmc4cr7Zey7pUCMm5KM+IiscT2nuGixXIjBReNyyBHgMT
nP4Lr5+3P0p7nbAlBQOItVUM9ha1MUBfIjWcc7AOsXQIZ21Th9gSszHvqBpTujNJEj83nhBUGW4D
xFNuoU3mE09cAhNeHjAXfGIvOr30oV67kYYjwh+CUnNUYXKzodbxZBAqeQfMICwNABGYJKOF2ERK
pnpVRzJUR+JxX0Zi0Vyj2G7C0/RePLkxrqZIYt/1aQhJ2wQurP1bTnTV5KE3ykL6xLNsJcDGtP1x
zQ4KMcEc8zCICe141BDyBMBQR9FW8oAcyoJUOKEojwITzLj45O9rLRX12a7VaH4Ue2fces2TKZe5
pP5eXMFmxMuH7Zioq3PWv6069CxSQEHmLdXogORyJ2O/WdP4uh6PoQ63Tv3/uFeZWfeL/4YLgzWO
y8MUYPzqWbrlgG0ZmRr5ndgeZLj5GQig0uxTsRZlg1s3A/cz/a47y/uP/KMyJewoozYJlg7mh/jk
n4W55h90ApvduadVrSbpvBa+MlAJ/panu3LSLMPR2d8zLVa7AX52vcjYnu+YNCUwsGrsqQbCBXwA
KkDrTbUdSZInGZu3/cKaOY7Ilk6Lh9ijLtTTN48cbSHKs/unx4lpGaZAN90gGvtycQ5V4OHLT51Q
2MGe+vbpSrPk/0rzOxEKLVk2y4FRLSA/FaGtiTAY7DAXfyv3vewt8YfOGDXJ2oazJOiy7R2HXeTD
CfSdGdkmeNfBj//DRSrqaQL6WJ+Rh41nQqHTBI/TCLYOmV8v9yXXaf1nclrUp/z6uI5fknj6etyl
pRGhIEsv5zZhwGuiseIpyqp4SOCJl7IGmQP5EmGZIDaZIKXHtQ5ReIBA/rQF1Gq6bse54H0xCUm6
tUcRpTt5n9ACOjK8nr8ZAtnCgtrZerSKHl81fRbwIxFdS9WpJ4Pn9UxycIwimcx4WcSK3OcIwloc
9fY+r+Oc+DiNJb3VXgiW0FXYBHHXyP0iU3lDHj/yVMHGrjDm4Soi16zdHjDP2k2MBdHEefBvd56+
NpCsCiA1yjrMD9zGNWOYElJOE57j2dq/pB81JNKiB0gow0uE+6hg/u6rkMv7/UavBVnyarX6pbcQ
NcyCsLPgpeuGPWXf1i/lOfgRK2rBAhzqyPI0pu67qymFzCZbJzqgs5SJ7eXtDaU725MSZnAY771R
M+DPxh9yCzEcEJ4qroyTjKj3PlrsOHM06HoV6ObhWNXmmWdMX7C+gLr6S4sWPQNzK0FaEBtvqoj4
lF0kfP+f688YkuqZ0lFvxUOMnN3UaSVhz8tN5zxPRNsvKFQB9dn9A/30APbB+cQGbaDP5FifEJ4K
zNURLUEx/ZY2ATXqQnQ4POxwqgdkE503qpAyL7hZh6XNaC+zZxmrSgYZtnwrQqel8lAqjls7LLaA
aij6kGTXFs+Ejux6aO13L4D54wPFYG7t4915Qbs9W0lxqPS2YoqltVAm3fQdw5ADQbpnEvjJZ94p
3Y+g4SE0+wcaJgCuN2TRH3/uRR+4gFfrIqiwJ96jjSJAl2Oy4FdBjJVmHWxPiP1ApmVxZEKaLmXj
lvdkYX8pquCHeLubSi4q+jWHfBOHvu2tph0jB0ISseLV0jBvLkFg27bLEmEXMjBsYrQ+7BaMIGNy
rarvLYE0QSf5Sn3NmhRmmjniKq3NiIQDhzNlct5glCW8pq9OK60Fq9DyosiKRdAZi41lV9BzBs5Z
PaYLAxGnvKuPpYNByaeMJSMNYf4TblMGUjBy9WJ2h9MwCGDAgfC/eSOy3uaeQUYrndeyahRwIjjK
gXNPX7a7uyJe9PAq2lXCnA5ol4A2POTlX4Zf1ZECHsXbQ8Rpm7TF8hNbxh9bkCkgvxCg03lRzSjK
ZmE9sLuXn9hupg/K9p3Mq0zZ0M6EIergUI+YVKlRmmpoymuoEz5xp8y/sD+3zKxWR2BGj0R0JwUk
lSRVEtWNMfRumNSpQTgtwQ+go8M1P2Twbj3uX4RkXLZznWV3uWI9/l+/q4T+RCwnhmFRLCTf57Wu
2GQFExn2UzCH0vz+E75mesitCdsz5LW+UbvLtmE+MzrSb6RrChf+q6rPgijxLb0NSco88UtSxRaR
4ze7u4cRIXHIoIbtAZBuYW0nY2+j+U2GUtWsvXyDrzep7f7xE7NfSCKyMDuI6+paN5AsetpcGato
NEo1HJNfAiljJQY7YkX2g1wfK/0jUwRYij7YwVUUGexcw0RBt8R88Bf6TVC2CmbExORipfgFc5Sh
+ndAvPxPjH9ZcmlDBLDpBtrZsNarZI2yss+GxQ9dEEKP96YqqoX7OYjcYiZxqOiNUNWIVtXuKBzP
flZviayPljvt7oeVyUed9NQtR7tYZ23OrKXh4rhxk2Rb8Ha6YdO8tqG60sOsGyTy+X9BCl5+es1j
YjQIRQ6tX//1iDwu3VrWhQkEoUhP9vvAZ7Xq+nfcabma9wH1rB87yl8MJEiXL0WzrO7/Mmo8S+8n
VXBAUXKktRtOOheH7FvY2R1uGuG3UntUVn7EntL6qwuoIGznb62JAOhPJ3kVaY4uSMThQL6WXKco
UgLXaXUjs68OZUtlS43i20xGPZTeCTe/WS0fK89XqBMNMmoGG/yneoTksMx3TbjJgbh7YS06lPr9
ifdHnok6Sh8sKKyK6ZuYOjydbFNw0BXvLQ2duuuMzgRTDXL7hqEjIYk95P1fTb1IY3oiJUL5rib8
WU2PASIdOqr/VB34nZmGpVpvQO5pF4QSLU6zENsF8A0PX1V+6TpUjhtZVmDUwCNrAwxLlsrqfiWd
UKcFFKQ3ytpMsvpU9L+E41KsQE5P7XvPhWW2IPf7RzRTsgjEIFoQt9pRigAuWGr00AA7DApwIkRD
cMpD3fMp7eyTIdJBjfLWnZzeW1C00utuJtfOaRiKtaneiESBTiTA87B7GAVy2KnW9DzeSPxG8lZj
I6aA+7NFUxJEkS8zxgbdA5NAGAmQ+fm2yRdh29XaT6YUuH9o8gd1mEKzcgF3i1a/82vJA/JcZnrc
nnheLTcQHTBhekXwwu4s+W6tDzd0QepragjTHgEwiJe/YG2VRs/KiYdbMjoTK04yRpKvD0VCkc8C
tryPzDdoUq0dAlOBER+6EIbFepScESqaVfZ79sjwEULERP45MNpQCI1nzBL0sh6W8wU6Ci5xMxbV
PnMIPiEpUbGICrp31HReM6do4VsFtpJpdIlL+Yuc+8mLFpx0mgmazqIqqVKszL/L0/6Qhp6jMao0
k9UVe+7iN/I2XwwS8elpedmmXfou83O3o/8OZWmAy++oPWNtSLJdB0fqQKNFySEuJkb6WUZM5R6v
6bPE8xpqiNPB3UmbbVOFI6okApkJ4uQpxiOqk0DMMFZyH0uerfj8cVCkzaENY24kY6Y3NfT9DMxM
K1tDH9wZ4uliXhCJstUJeo3AWGYLT9vbkRRsLVJI3fKFR0fYUKMi8Ta1CgmrCFq+ABLDHz89m9Pa
rnwj6Qf6bt2C80PGjcIwTxVy9pUQ9znNwRmjLTsSY4+zv3ebAoygGtAH5TD7ZXX0Kj4/ezT7lXJA
0uYDrs/IcjdQ5tx7v83aae3QJQTpgD2WqP59b1iNQwIYKXOU0xVfUmSkWiMjPCPGBfbelFPMC1XH
jyF03mG6CH4h4hhXAHl8QNXyt9d52R6bqhAwt/i77zK9M5+dYqpCrF8msCuKY1kUGuz4cPrD3KDS
4eFEM8kXnRmC3erPpGw3IHK7FYdfHdsTQHKJgl169vTca68XmlR61p0mN4R3/FQesvd+OLwA6r3V
73WyTAeSN70LPocNaGaczWI+vT9yBrjk0XET/DXy4HHVfmRWkLlw3inIWWl+nGGIbDnMEIhE7ajc
ydVMJX0wkE3TELDO9JhEvifAg+D2h+Y4PUuNg+JFeRi7n+3IdI8fUYYLK+KmyfB9KkQdudmd2npi
d/j/tqXRn7q8GLv94y8dihmoJUM55Snv84k5Gf4ui+d6A29r4eES/74d7BOzHr26PsbM75Ghmy0D
UtQgfeGC3gHPdex/5IWXOlxUuDpUbx1vYWjJWz01kFyZcs5e0jPnqJlD/O/KfPvwIYCxg946nTbF
dDayTAryT+qumATfa0bAHfY0H5YxxJut3wPedcxS1iuwQSIw/jUEQhyGHMG2SFpPRiaRj8CCp9PM
z9HBYi+DY8LsvO2+o7zgYaf+kwcG6VYeR4RC8cL9xdnXuRDb/DeWkYNx+as3Kr5HQzhdhL5fR/ik
cux5/Gl/Ep5d1rQjOgXAb66dqyj8j+eTQ0HRUS4/+PsSEgz1MzRw9vVGbrjBXksclqSd6i9XJAi8
2tpc4aJuYOvyFUrOZ1yizP9XZHdJZ3jVuPrFNKXH1BjRC3ymNx3TxlSmPmJaM0Hn74PE5ILwVbit
eEtIp9fyEoTKWQQJVGY7LryXWmvyvNJs1FX2O87H17vUKIj4p+NpPTLWkRcdn7mijTyXS3ZjEtwo
ZG66Uw/tI9Iz0aTNDCriQ5xJHS2jYIwTfhxipKoaJdpaejCb5MIaQfoyvolu+i7AuzEpj+lrL08A
Hz1MtFVxlLtA1pUX43TLQelK2H2uNxxd4EerkOMAW8Z5sEi8FKdhR5TzFHT6NkC4RVA4KJs49r+1
YyWgu59DX8AZ9lnmKgkN69t9GvjjHdVVumofrz9DKkJRh82zMaX/g4TWwgs6am4W6MpeC1Fi9lVq
gHvIJBujcMHdSJRtGJzmoYD132yPb0Yo04y51N0rAWs/J0IPILDOhKuBTmXJ7tNK0zOtwEkQdvgM
jjks4H+iwiPCD0TFQsJoRgc4wYuktW2QzG4H/d3mENJ+vgIpZvbP7txjdFNu+7YJzyNwK1RMl3J6
dOjXGmGmVBDqy5mVDjuYwSlbgw/mGfayd92KT5mU1p0yr3o5Zj4PSTa0oKTaauqG3FTIsQkCLdSu
YTQdB4VNyIszZIDoe+9ATnce2UKAOcc7hZwGdpl6II6i6yeOxccqaACEb+HEoWTNpVN2YEDyMRSI
8fKjVjvq8nixyxwHiDM42AMJ2gPhZmVHk84D13tm+lYjcEBeSVmE+9ur2Zkbwt/thawSW4oTNONU
/Ri7dHOqiJNiV2K8fw6n46cR7jOWZjgYYzwe0Maip8vIbJaAZ75Nam/rpTZgSafQT1MHYDpOwpnM
6Wa3iC+d4N1TBfnucP3G/qAUh1pUT1J7T2j2j5Mhj5CnfbeiCEtn6GXoIEvbCgReP4nqMREMc0p+
uT5B/7+6JTemnnqdiM0rl1ZLpMZbD5a/Mq1OPv4hFTOZIPhbEM01NngzpI/qRjdxjBUzpRIINhey
msuoWdn2Mzfov4oPnCb9nU7CuEoXiTMvZnNtCAQx2C5mPnJF1RYPazCQF2nPukbToYmoyF8kHcia
BvEz5BraWX8lenUvkpKVrk9hZPpAZ+pH9/rCJu9/VbGjC3LlFQeILVj0IGWaeKQ/lUZ7fFKw7dv4
NuUQymPIfiFFgJlzyRrTGczsP5wLjdvdKjSbnuUEqZ3jRcJwrL5smDKLpJwExszmajB/s/ywYiy0
enbiNZbjtFxWcXMpv1VTCTKimxcJazTVwuJVcgkFTtLPN8KlLw0jZRUzCBTmRMUakMkQod89ahyU
Np+AKnFzgYRt3bUovTJgXaMAHT5w6K+wQcLxT3Efr2N30I3zjeOdFth2p+OgKj4ulBz5hSiod1X6
6dKnE6NiaMDX07prkwpNTLT8P4kPAQZ1A/xKQJ5zXpA08n6feW6UDQuQWQF5RcVvU0MxRmyK8M/F
YJxhGidMzTgn7QSRDp3XmJGtk6M08hvBg6/owms7GWPEdAlqpMdo+7WnzxNFzgzCHWJnbtJffq0a
II+C31LKDsROH+ay+0CWaQxoL+/anWA0KUOjKBMLj3qkjEYcwseknP0/G/C+RLCS/XNrQ/dQfeG2
ZHue8U9BuB8KgYhq9dKjrmnPdtBBXAAKoGoNUA6gRJ22fTRtV+crXN80JQUahpKqxAG7TIJ9exqL
WfixzQD4cL1SEKvPWAZFJWAoit/TNs6Ubu80bP6LvUvqJzU/yFslrA1KKhcG4iq8unYp1cgvZ+FH
GWzEomrkPIoGuzYWakprnJt0zMaby3fsT5qxdFVft+F5vPC/UXcisDj93j7SXnlLyC1fpdcMR6/+
8sAqfp83yaYBe6ysTDJRQHjFvv8QM7bBw9vqmKLXsguGqzgzhlegeXdt+GDuQOOIwm9Ri17ttwr1
88PfQHPiqZSV5QmTnXw3LTRY+m9N1cX2myPMSWUB1rJjFXIlzFFTIifnHlRUAhlOG+NGTs3ppe0g
QvFUefPejXRkTtgE9bDiXShMy8WAoq4ymo5s7voNxtNxhOGJLyL61GN0PCrbE0iBtNKhZr9dat7t
xj6BU/ft9wNJ0naR6c3ntY3wTGJosmRTni0QESDqyTv1Pkeov8ynlWRCN5BYfQ+xndjNznzZDCuO
QMDJr7xPwMSkEw8zogVgiA3xC6gCos7f7yJgLT6OPX8+d3gx1hPbdc4WsQshpONz6AuNGdgOa2N6
Z5dgAie+pEz1m5stusNPoZtBTvIwLPEz5m5CwsbF7tTFrdNjfPHzIN8/yv6XBsIkhEQYi0IaFqn1
hM9l2RFJjdomZh9nTMQ42B57PF6yLWhRjVhq6wSx1gdtbEQ7idPqg0b9TNe7KBVPDaX5IxTQbrTs
aCysgW3XlhUhAbrj6A2Ph5413mO1PP1rDB7lMX4H6lFd9VjRxfHohvANKYvhKuqkgJXjSSRVJx5l
RpmfZ0jBGbSSDHm+WCfbXZ8aunEnylgmPCCB6qmw+QoTJf99g3wiVg1TE/AMn1+ku4RBDfXV9Vx9
BIA5rihl7Je/YAieKglR3feqJ8PTaxsYvPg8HE9KUp49uObRrXvKDY5nibEc8DBSbDAsJqIGdydq
CJnpv415tMFUqeTR8Pye6hPRRb5dklwB8/CiPwo+OJaZSxJ6CQHuey87bNk9YlQMKgUwSOshvHD5
QDvN9+tTAkSpIMKYaN8lj8Y927RV4TY0h4P4RFWm9a/kDfxq/BQnmgwfOQymW2DMUKEycMCQWcNX
STN7+q9XpC7PzDQm2Yp5nIfE9MEhg1fur4nWXTy8cy3J4mt2W3+phxvTf7mp9KObpb+YOJAcAkdD
BPAP7OO61rbwZd6UB1n+DgSfHkQceCEp8S+M49/N+ifrwwFS/ACKkYDTTAYx2s9eJZdE2kQdN8XG
mh3AiuRqszilu9mYnl2wU6XqT83KCCVRyYNvxJ5LtYIb2upR6T3N6zWdj4T8do6YsXewPKn3ur5h
AY5S+YEPop6zyFp7SQ6r+2Co7xsaIIJGEqm4TbdtdzKFNLhMrUwl+X6iapnOz5PpYtPbcXmb6kzs
GJYayxZ06itm5ujzQcvvBjN07MvcRIuBDebiKj5pKmfZkNa+4nuWGEeCF/uJLrs474nq2Nu63Ws0
eLC4NLtwac4uvZTTIfcnD/b4DG8o3ry8p+6HXVWtmE1G5pFUUWMZpUu2HtVE4F7M/MoAdsXXyeQv
pKEd8hFm+fhXKlSdcnHDBJhvBK97Km5UHhXc9ifFl0JmDC3RIv8GdlxgHBasWJAa26KzYxhEgqIa
C3j/Yet4YkaOxHCtuFgo4dcMs/2N1rVNxIUVEeNpsCdFhb33dEeOOc0sCkLFJ5AAURIUyY9i3OhT
iuDLYoHsP5P9cdjBB+9PwTHyF+uPKrB/0mXHvXclqu4hsvyJgpuQ9Arb8uNAhknx+UIeehpa+00V
dVQxh3HZUPN1e4DABY3wn2wLi4bInztGXQCrlT5VyJgXRxnXBkfU7jW+8g44xQvrQUseKpyfUXBB
rDrmCJ9FJL/BKeWQ5C/+c8UNmiYCnEoJD9tG5r4tveInPEPxMrZYcl+E0flK2v3VoJ2V/OxT/IiK
JJy0+rrGMMvJ4Zb/rQB0w8a4ONhCGFvdy627pgMaJyvn9S1FZZyJuiNI8XANM6U5/f/53CiR4T69
ceyNJyoJbY8p7d3tkwG0qRwfwO2tyHP95+D5HQ5o0WRJqCfP8TlA9Pa4XaMKE6zNyNcaXWFAwQsp
PAQwbGxtWpsOZwxd6KRKefnWN8Q2mZr5trUOFjSMIePHOzyAZC8PbQDj3jrm87dMYvy6khu+56A1
kCEMIMiOYlYmUdjlKqWPOg88jY6Ec/XiTJae9XsY6YslPUqfAPcYm7/oARu+uZDrDl9+CDqN8U1A
WmUz0mwFo6RHr15GX+yPavN8FosIm7Qm8/gNuX450uLbmzSCA3aD+74Ia7en/XVyPuatXUxeaTXk
+1sG0Psf9XkaABTl43Yd7QeT+aBKlLqGLOpD4b0IVLDFU90R5QYO6C2HlLIi6+BmMq4tuOa1C1jv
xIK4kiUjPfaH+saGmsY1jsUotojv72wlI0GI52xCCZRlE8S4C+7nwOY7m/xbjpIxPDArP3pgnIPi
9vXWZAk8P+Fawp5x8eeOzDDy5fedw0ePf+2pcJZRAad+gYf/0WgsmzhQndpQB/fXMO7x6i8fn30k
WWnT1y+lDRhRyT9aXeJ7XTSZrCY0239EGyEECe95Q4bhCyaNHUpW44cgbf8m8mkbtRG78mTDChT9
PDSBWxtrl3FZ4IIviGbola14kyfr1Ust9+7kHxlIA5ynBaAY4EDaGjynxa/mMtjK+e5Qrq4/mcwM
rewuf0oMxRqwyz5SdhcldKYE18VY4zIRrbgWIQlYVIp3tmB21eLtn5fXDa5EI+QdqjRQ45jxLOSX
ZO0UztkxVB3xdvHAPMGiLUWuKABuAL6TiLhhj8sLbej+ZRdkaUg9/jupJTfq4/gvR7GPhtLhKC6b
h1T1BJEsguiFeClBRUDykVgfiPO3OfNMchZG4QFBBHh8+KXqIFqKnWqQfG5lDRv6TCbkOMc5v3Tn
6q34UTwBD5+6NH90ex60ZhfQMszaK6rjJXLQQ7wMjkM/JdEMm9JZEFpZq+r17NXIpsV3qzYdM5nq
ejhgeMi79tfAM2Y/6hn8WVNvIrGL9C0T6m5r44te2Z6QqFUKKAoDvaXYKEdLr+DIdiRYQ0p7WJrJ
2T1a+7wua4lw/jGh9otuReJEQphNRFhFtN71IE/VznoJ39fhMiGw89iDQvNC5zlyGX42D8oLfRaG
33oa0t5ESPI2PzGD4b/J/BZN5jH2lTvLIxbmHSlE75XLDDygGKM1VPXfJrnxAXFR+TzjVgCWansN
gV0I2ikIly1aohJa90/YX18bKvFvNpn7qoyGnuNxTs/5gLQiStEyLVAWRY2Mzed6jXu+iIXhHhzw
V5T+gYouN1sBR31hCDt7zRaRDmwoqRR23ukx9qCidAEW/2GW8g2CEAj/nILym9MZTGhvXhPYvRSP
apcRfR/kK7kVzE3d2iVLNxQl0Iv7CvELG+TM6VXC2fgxJYyvCoQs7MNAEHO3PE4kFgIERd1A8sBX
uoBvKAaOqGaVfWeKIW6C1kZh3Z3rel//WdG7WwJrPjEJnJRD0k9Un4M1PCpvqbXCgGS2EXSbEohj
tOJA7HaJyaA6q0wzG9FF2jOrTHYAZj3c9O8XUCk+iBfFs/zMH41oaDCmiujzoSO92bgqpB1JZZc0
C3qFOB7yOuVMdkwLKe76KCDbpJ8FxJomlp/fE9Vw2ROi/yzSyUzl4mYYs+iiGhoxx04+BIpSYZFk
E9RnVsmUNExxRGrO9qW/6uTuhiswTm/L/OAGiuq9fdVux3+LYnVbVLoSUxeifzVLJFc9bFvlhVKb
6nV3YZ/OumQrC9PBq3orT2LSrwPphFx0dmjps2qUkXcBAZn95A046ZA9kJyTObOR37d/2Fr+KGJw
GWGwtVei0I/VLD7pf/Qa0+l20z3OFrchfUdTOl01nNbN25EjPp3Q9FHha3lz2AIrUoTeKi2pgNdZ
atUyPGc7WXIA60rFhas0z2CoIDA7ZveOE2AGUaauI0gin0AHvCqihObFxuJJHW+XcTHw3gWSpHAo
w6QRWKkxxmyzyG/W1JWLuZgqyVW52lU7Ny94EblDvpVrak3s055HymYJw6sONxQs4YXhWFSr2Fsg
UyEvz/L6NHEXfbHm8SFJZJf2rvhrXIxoV5chkAN03dEN281glZW9o258cN20Ps+/hPDjfFiiRFhi
boa3y0vQ2dsxC5+COjBNED/LzYza7En0/apcYhKp4/s87O3QCCwpbEQdl++ZBd2EQnwqXKkWmXEJ
/c4MtkN6FZgzYrfXrqYFE7fqmcY/iFDjjO5N65TRP+8e/zC/6FW4kldVHzh/NZnj1agBrI/Jxeut
8Eio0uWRk94V2rGb+tSa97jb39rCERzRC22Jo/NDjALTaY+x6+lpmaseUfVdzOxWxJE9128lNgZS
u87mbEJcnr768NcqyIWR7pLLGmEaqvNi7540MBfHEfckyYw8RdnM7kYc7pHBMa7quEuAzPHdXlHs
VYpB+9Wd+NzZ4L4CMeyk34vycTC/qapMg0brbOo28eElHcVusVdrBwfuY7jheEJ7u5hbk2ZCyHSr
wJRtyV8eWdukiOnonclEEGcEsWpz43UfYhM0g8Jjs/M+5C3968NtsUUD9wMnuDjMXZjxRmF+lJC/
8PknVRamzAdtEI4t6KEvqa/ofMXn6llGmpQqYJ/0uOfxC+6t+hiJgFBkPltP3TcAgQEo/folvfS1
azb3fxJiV6GJMeR8YhF4YfPwExsu0bQtoYjmIYa+tKBe2oTMMoLbm5uyF/MHMSjXSo+rzR1SrDhl
Urot84KTjEWxpwOmKIJ0KcCyN3MVTbplDxTSx2KzPn+U44S/b8rZBmcx18Foj1EqZbDrjxxIuxj0
T8Gh0s/H16IUOnv389Ioc0TWvCycEN6uXAux4WI23dzMyxDb9jHmPxTF9Am808a3pDpI7xCNwkDK
zD5pqJj/iE8l+wy2gb9+JOgxh2YUPnPe6ShvCPyXqNmal+PGDQ130YdW0R5hSFW/CTsHq0wwS7k+
8T6rI0oz9OeXDA6fSLlBkO9oibFtFCmjcwY+zZfj9nBl1vb6SAKfzx+r1CpiOtc6aYwUXHAkWZnX
1DUvWImWyQS30Av8/BaiP/ZDcYPpwvAL3hEogfZrCi9VJdkiU9331ZIuG9y/Bq9DlYGAFWjZycpT
6Ft/9ES7QVFnGG00Xfa0kKjQm/Yy02+eXQUAJMM+PsuXZpvqKb/eJ8sNTgdJUTzD4hQy8JuBmN1T
cVDjSySaELLarKfW+N8esIYZjIsVElMBHENcTvGSu3H1pXyYv2jmYcj/aftzNN+BVpQsCpPHBQi3
qo5JEwLsg3DQS5piwN69UHpZZ4ZAGOqILaWMZtwJQjXVECr4jV21C3bxrw5Of/Wbd5J/orfDA9dA
oFOtpogL+zvzd8aX8mjVpPWN5qzAi1+SzQBx17wqI0OiJ/FeawsrPRWQRe1Nn6KPmcjjfeC5IgSk
oV2x5/GumzaMn25zWE1Ym0MIcQJlnlN1lkDbFxmswOkGDoxE6ubV8Llkey6yTwx7hZpRTEt2LCTE
Vl0haRUwL5ceEDBLXAcBoaHp5GpBj2BrGW4PeodHTaA5cnNCOaEWsxCYI30WgMGanJuF8ur/G8R9
D/EF/Lf1pDRUJsnE6H+agW3Pz0jqb0z+s4QSvPdIvuM8HJiVK6/7QcIxwI5LpYHnuaGhEIGRTh0c
rATIPIEmEN3DGqk9aFdeLTD6AgtE4+IRQ0zjeDTJUVcVKaJFjnrJ8yLJ+0o1jYrbQt4NRv7NesVQ
eTR1SUVZorKpM7kFDyEWexn43O2iZgX3S1spc8xndmgUmAUO1LnGzKA4A84q99cGtvH1iVBGTZej
wX7wOpPUnQzlehkJkVi+BfIFx6ViNP7LpYenAnA+e35l1LquHf+fyzLwq6cUpJD4Rpv4MBaDe+bI
CGnBjXAmeZAOHN/tqbTKvm3g1B84GQYt9MZu8D2xw5f5UCzTGIALXjy/QKJ5tr6PUx6bLIzpK+mB
olJ4pWtT/HVqmYdbV3GCi2bmE/rF/14iqMy6/pm757Ivtc2mk5uN1n/Dr4+FCcA5/ghbyiYbMsct
WxCflWEU5NdcYxh76nH8hIWK9o6Xg118hB0zcEq/kIq6YmrJUmnIPbIYlR9CoH92OMmnbzws+HYz
GGZ475IUpm9Bs5i8cGpZ12edsw18t4ckN4cDJjyJeHAaIwA66f7AQlqDnHpoGu886H+B6SUN9IrG
SJD8ErDrpmkmo9wqx0trCX7KJY4UxWJ6rkLWqgAuBm3J8CRtsNjZsSztvmg9PM8LjVJUhH41AR5U
PZdF2J18MU3mfTsS1vwZ+wTReXzikhJ4O2+kqfgln+wHfGQiqFln0bDuQAyaaSumQtZmHiQHe0eE
Ybc/jn7HJTJe3mqYG5DRWtwxrS6Txb6sy7g21UhMUm4m7WPH2aO/J7XmPWMZt0aE392WFh4sCvUD
g2QPBnSOzUr9WEQXyB+Y0ZYOMZJ2KnIODoXMe9N3r04LciKcQAqrYdecgzk+OlVzV8UF64la3OLF
etow3NPAb//tVsjKJBeITwG6zF5stQvzlbDltydm28DWabLQGssfPFma5xuEObU9BJehSlNkzlwb
9aVvUaJr8rG5M+Oa+rm1PWTwI3E+zQ95cYsQA8ewOpe52KQYxfR3utKyoUIXgxc6a1Ju7KVQNOJr
n+ePpcgYEUHH50etaiaowQ2plRqdU95HJ9y+YGZkSl3gkca73PKriVqax29fXDD8CzWPQVTxqZCe
w6RS/186BBNVh6WYOn3BtEqfFRxKXVqBr/U/ny7Q5I71It2GI84clIUtZUugWDO3KqOrIp3aBw8M
JOlV5pSqQcU17IfnXXW/Iszr69i9HkdqmT8x1tf/979eq4P4HFEhMbz0l7qdNk4sgklOMuN6dLKi
/wruE/ivmhk3eZqo4qpOUjPSEZJLw5Pc7jMk508vJfzuz0HOUFJeSj0bMXQgisJrXm91M/9rCk2O
PGFLSW+1x7U8F5y/wLfFKNC/5xcD8SwILOYL9/2FYWNJisePae3zCwv0uo/FDAHzogSbkJVox/Jb
oT81N7yAVrivkUpOgHkaJIiJgHbs+GwPp0Ie7o7JXZGnx847Z/7ixH9BwBTiQ5KYxSajqzn8bYE5
qydtu1lT2ZpELoJbV4AXFQtTJuBCxZCqsZFK/b9mP0rsWgP8plQT6VEZ7FqPfbidGvr20z/s3J1h
qzhidZtYGmn8su3q7hEct80gujSKZClQoO9AKvbkhAKsRCpyyu48hQpxkiftsQN0iEDhyYamUwcn
QLW/eC2ZszI+5sFA6WXlwFgJoBxUhd85rNUCeP+L53GNaiZ4lXL4CFzJckCLE0I2nDePbiCc/kBI
ZltizMmMNVMd5/PsaIUqhfr5A1n8CIa/62p5hiRCrr0+EzmNC8fczkHEHrYZqXTvOlS4zV9bnLLx
wRvaU7kTQRkP51qsSQ==
`protect end_protected

