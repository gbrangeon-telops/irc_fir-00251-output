

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XZtM4bLmkglBewlWavfkobXOIMkrnElgJo+k4jE78ykb7oIZp/SGV6Fmfr/ogrusY/kHxxmgAde8
wVKEHfi+cw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qj5OXRmuDbyb7tXOe/IIP9hVzpHdYEdnGFMGPum5TPAz9WJzfNr2HnR7yYGe719tx6wYAvdRlfH7
1KYaZqML4WollrpclochLq72pgPwbtC9iEEWlamVuKdvYSw0+IzNRBHdKqTykxKbBvXaQ7+UOUjw
UnhOWIyi6vA2XCWBMhs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wc/9BtL9LkvfKqZJg7KOk8nPkSL5jxvAGfC0RV814LDUHBZcOVMBTQdouKf45+uYbzuqQuzhrFia
FyTrOU0b+Dpp/D8a4O6aOPezhZlqDF7SuDaIsbNJNkVeEPTzKN3+pib+HJ+07zD5sgOQyBLQtobI
4fQy7ggQ0o0bOrWPzlXO7kD45yraaLu2CaLqYlQzcDjqnvaWtdvg8Q6aRiloz0plB7OdNZ9a1tRM
Nl6v3ocdKRatScwi+YnBgJn5ewXMvGYuuBOXAkUmcc+AFWML9u7RnCLEmrft5oAR19N3inWP9hTR
9sdW8LGJ406SdzZiv/gZpUV5t/AFjTB8Nihgew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RuHNUBMTP+a4VfkYIP3nKug+Q6Ygohn4DcPwrCybnrM/u1NLZNct3nJM51Ftp2uYn4LtBCAEFd4j
J1ykZQnUjNHc8Om8TkpAk8Xoe4lNd9c07VFQ/PdNEPsRZobFbRhtaTn5kYtwFZszGT2+NVjW60i2
zzHWmeNAYn4vMcnLRnc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M1UhZ+OMYDjkT/STr81dVx9PmVVG5A+2IqAmn0405vupx6bbRZIy5mB6w+gLHolhJXN5SjXXAhWo
hTPhhYqRE6WXBSt+aNme9SGwhhYQCQHfdP7l6de6Oriyjp0GyOVTMXW7th225i4gd1/MFzrJY7uC
eTxBA69zF+OCz0UpsBa0iiqA6SmkbUtST66y3rCQ2iRlo3MqgxqTXadwVQPjyKh+YrZv8hSoGQfZ
859BObwRsVOuARh2h2mJuicqAywYo8mWCsE9MJAhCYkJvjGEbdjUCSpq6KjZZuBtdg5UMkBgdSnW
7odTSYiZWcCz00u/B4xtOP+tFTZhOrGrUTKipA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 81744)
`protect data_block
hiYSiBUfGfvyKwao0C0VgHXjfJWziUXIi7gBoyPaJaJsM+3UxxeMfeJ0gv8WguIB4erH6EgEWAJD
/1Vsw1GxA5vkKsee5407dDmagnww1UzHih2qt6gxdnRLze8pRHdon/hmrImUMkg8P1qTq8CH+KgA
jENFOWHwSvwIXJiYGxNhMfoufHF6xSVgW8gzvzxc5oLy6uQNTefyGn2f9h8jGdzYLjVOegRhh2mb
lPMWhREBGyTZ6GKkQHup1OOaVcZHlqZqDPa5CbKGluxMETQECgywygs0dHMtZJoISBBAnOEORxZ+
EyeUQe6xiavJ6ViG1jhEi3E2HXvawg7o6adGGg2vKtGX+vVXmdqe70ttD9y945EIfIluQ6tIW6N8
de6UcDWuHD6M5qqy6mP2Zefj6qylgvsa4fC5keXwyZQZ5a/tlJ2j8a1BQlAad8ZjtD3gak3vb61C
B4AVoISAeDjYGIyccHny6KiP94GC028qn04GMZ5DGH5ZA5T5376AAgmARN6VM2wW06MGPqka3rCf
cH2wKhGgomtzclU1w1VbYnxpPLKdHr+1Mpj3jwXhgRYU13YDj+nWuHv9kDV0e+5h+ZyNn7ls5e1t
aT1OMVz8WFWPCbCinIjkiIfk9ZHI8XbU7JyR4UwFlKIRJIYoDBf5KQWwVJhaCxjvQUQqi4eTJXNg
EFeQ3+7OFBQ+T6KqTjUFIG/tmO50EpiePcQSKXkAkA+ElS1VVsp1P+dyKIwFHCbc5IY2sjBfg967
0ag3/LSDK2IrQkhWFivUUuJ6XaldO/ZbHXq0LEkJ9DTk7tbjRBM+3MeQVJ8G5O5NlIFXgG4uTNBz
PycJUu0RPrY6OJxud4p9wH0NdpGaPclr5Up1f1hrb3IDiaQNrkDUYJQXKl1N66uJfJ9qzSHQ3Spk
brshWKUJNO99opLXurYPEw1/j3iTqIW+H7N70uczeQTzxFcZfk1jtG+8IDvgWhNjzzGOGx/2r14G
K3OdvxRgfzmYqOvvtVXiz1BnKn3aFYEpJYRdxOag4V0/gfKHqMkG4v1a4OU0aeGdGinY1/41f+9V
baNB0rla2uWv/zUUp4xFTE9YS7NJmVu2WylNbtdhehSiPU/QVeenwyFKyDZP43vqrLNKRD+naYUp
1HKZ5KX048pmDE9XykbumFOpzp1jNAelMIrlQTtzqjB8M7pweKhE19CX9yvTtnbBDVygLodJLbT9
2187zn0OnI8YQ2DNLRMH2sstf7UDt8LECxnoRDb8iV7edRS1vjjJLt96OHwxWRdRF8rC6Oo12/2O
zeiZY5qbu2SpwDQMSCYOJYtjcGYg25hyqejLflIzp6CmJ3Ula/S5skJrOqechLSix2fswHJXR7eR
lEKGzp5WdLYcA6jQ91cBqfNZeWNR7QhVonT1BZ3DGlalVlfqQEZL6DpbbgUE70CvNqiVF1fNXLs0
Kd0mbjldPUHN+aG0n1+rcoMYfCf7EQQLFyTqgZPUTNWCLxH5erjM9VFCWJiglIz+5OpMTu9dXL8E
XT+u7D2U2PC7eCO3TWfBReqJ+wZwHApw5OaoyUiok+eNiBE536/x5oXYTg3HXCgXmYv9iqwy+EXb
BUJxxwLQ5F4g6TmdeEciPvFOZ+OPx41Mf32Xmx3MG8bADhjuCOoeGFznAngu0Vxh4UcEuzwO8KET
o/+Dm2i40aZLJuv5MX38m30i7w82W3DnVr+9ZdnvE4ZyxPOyqLeu5XwheHsDKPSCA0hnKtpo9ASj
dnfHCpLry4gwCVudKyTO5M9/HUfSaoaFcHauCGr4Iuy/j0UVwuAgoioTIaEmkB+QgDTc3nX717p5
40NnIBq01bBXwgfAbBkxNV4fK23GjpbquNCZ26zTctOTzOtOUqkFqCa+TRUcUi6wehAopTAP2e2A
PlZr9hoxQXN4wjB7DpQeBN0QjqIdeb2hvLNoXQVnlq4epIcNxbHosbi1T1IrIK3oXGcJW9I+uzGw
4jetCM8ldeWTZ0pSCAOvC6MoshAaXduMvaYG2xOJoJdi/A6ufcCF1MnUiqRptXH9RWUTp/ObiKpk
MOvy1afsjmCC6nbBIs0XfeNZGt1TtsnpLHtPYEPET/tVevG2q8cT7XPsBiAeArQ3dtMdOxmx1D0b
CNaHQ9x6etK2ohO/H33zs2jF6d+kafEmnx+0sNC1pyfA60SFcSF1a/PkxuucxZWRXtDvNMGUrqEX
l5MvznuK0YZ5y9DT89tA9GMTWoj76e3NVxD4zmHd6f3dQCHGaHjJ4jxFvPyltKV/++Xy1+a8xf1x
d/cuEh3z81lw3WysRii1wwfAeZDUB+iC/mAFgkgC4d0uq6e7njfEjH1O5Zu333CujLvYQI4DwN8G
l+2YE2CB2YZKsmbW9ISiyU1cpMxhWrE9NTQazd7dpBtS/xcDCCsfhSlMSn/s2+fFcbkmm12atQ25
naB7s/S79MkZkkbivbwrzOKSsfFORw4IvYsLqt1o4lu6+KCW5O+5CflaSKCU5ycXD2aClniuPlOD
CTUfeju2k8ca7yVVyddsdQDz9xZ9CoLKIv6nkC32NyzUEgSDWpASeWAmqGp5eHk+SHe7INfxtCSg
LA/crKbmukwpC04ncxCn9mIz5OR9toE0ClTbPQ1YI5fTTWtfXc6/ouNG2vO1bNQ30/LuA09HILrs
q0vTLJ9p4cgBpzjdQOIz0l4ZJZm+OTnmQuidnpuJ0VrPa3pmrHKqj0S8zr4tyLlIMWTOhZiwXfMI
dysTdrRkW/iJfzAqUsFpnHMoMuoTHlCwtcG37ORYcbq1J2KBJhsc8mzfeAMeMRPMxca1roY8K2gg
AHyyvhDRLMoSYIIpWg1JQFTMuNek/N6Tb10RYTnPabD2EjFg4ZoQmDlF1JgS2N1xC7bUVfIE+Uok
P2BzBO4bWyTrLa4+Jt5cjzprw2Of/qWwFscxIOOuQp4RH/89xDB84j3hgdv24eitpa3d2amJ/Peo
M85BNVvZd3i+VUHAy7hSKOfd+MYnvg6tDZLviBL/WUJNbc77RalTiOYh5ZrC1FAvPXTUXeoQQtnY
CaX0VuBSyJ4oazbjO2uyrmc2Rbwmv2Q+k+agZkbP8QZZYtyRK+5nNC4w1weNyL5nan+U1cxgaffI
6DPCJLm2sTdSe0kuzeKFxXTC08taP4tHVZGejtmJE/uMR0IdDvkhe25iTsd7nzHLh5qknmA4CI4f
VMxTgVBCUKqNQdFGR1eKAnaS5L1oHdZP2785gXQZmbMUYjR25Mfp55NcZcbSZE+iQChbdYIi69t7
w8Lg4bBNpzShrVhSysoLauB2fFQqszPH9YGE6RpeQ2irpCsX1Swp/P13m1s6cHhQ1P/D9KJ6aajL
6n/RUas/fUaitOdOEfzlkIaZBlq9ZapBBQAX0cXpG16qQBcbdcGkxOz1eXpNu6LzUpEnDfGdomSv
jFK/fpy7FNUzxNPHIGpV4IHfP/oU+c5E2jJkahvBrP+zhcviPCBkECH/CYwt9IK8LCFykhrtdajJ
yND7kppErAD+3J7EtBz7AmERdTQsDR3u0hMu8oXEF8xYIwyQszk+Sr2YjIhTK0eK5agyUsnFHFnw
rotnqcJ+HptNCBjSyZadU41YOB7J6Fjm7fH5G7yLXoP/8Ju+k4YQ60LVMk1PVW73urWZ5q79LEG/
vIEUV4E4JMk8gTmjl6+n737yYcwb1dkzaedmHYcK5nvg6ecqRYkskTmaDfP9vYx+vOLvfvX8gfkJ
njPKfgC+BuFlqxj/zqDezjY/VTw3sXdZ5h92l+T+rZFAtqPlLlJ2D8IXIlCowkNOLwQB8DDFR0kD
eQ2DL0y+/6mop0F8MsA9GsQAKk88lKZh1rE6ZvvKPitXio56iH/x8IuoU0LDWZ3G8F9oHnNRS0lm
I2+eN7rJEshMTqzdyxXlNA9BG0UNEY8ICxAS2FE7ZCgzYYqojcqpMg1dGAwfkGK1caXjQHrHfDRj
phw8sYcoeR+AzEueWIMTzpKfmxhmpuQgMjB+/I07bZ2H2v+EaJYt94FFmL20S3ovBp3R64qccKIx
EnqV40r5KuY//4OEoOndiRvXMsEp+hlyeJCcc4gLwyiL8Ie6KnubutkHZSAuVS8v3oDYsY1VRFQf
O8LqNHB25RMVPhdksvY4C3IYQ/pRYHAPB5vIowzd5sAeVxrDokhvvl7e08URkWwRDltAXSmhGija
1rugyGDyi0bwv5FzCfv8yymNdLyUL0bVztbQqA8PGeTuuxHGgY9C+QUr9Lr8TULNHtf2CR/ro6v/
fJxd9Nz5rrC3Pnc+7Xp4uY44XrF5ba+cknIOhDU1+n7GgZMY/CNzssMxb1vi78RN6Ly6bmtUxzFq
oLblhIvk9rb39zGbDKNbzsFEzD6R+A54dDrN2Z+OMX6y0Fbk38G4RfLPcPYjrPmHZIZ2SUCaKvMr
AjN6pboe26hEbSnE/EER6cfvxCrDWAdUm2vJlnq2t2+GQ3uTC+DpNqLxD4bkUDqiZXikIbpxGyt7
FUWoB5v7i2CaKbOxGRBBGXBLcU2a2LmcVMLckKfHqjT1QUa7FJ4yA3/x04VbM2Ct7uduRUgSm1rI
xlJ/DvU8RAOrJFc+UIpF9/41KUkMzGiPxY1RiEokAuX2J5UYVsw4EhtQHRbd/Urzc2r2rDQ5q0iS
NNTjKIq+Jx85TBA1ilJGhnkfGmmuU+W6sJrDaROpuFnyyqNyU1gq9nsj7JnlRVG8NdbmcZAniNOO
SpaeLuUCAVUc8mOBUZS8yd1tMoUbCoWThY5dnSPtig9N9aj2XKsqbCTw+AWWxuUnZ2RVRecduXHR
RCBGLjY0k7zFMi8FsB5fTiyrFpslGc+DPZenQWNY+Ygb/Jvai2HP/2JiNCEokyC4i+xzSFjbsNyx
CO9gYv53uo0F0e6KjgLoUgkHD5vkDBbT1xP3po9OWxkH4DwZLfjjomGD5zw6GmSOEH+8mz5ku/La
B3TP2wfYcIrve3/p8IO9WbaDvau4tXksV2YQHrsOmXK7JRSA0ayrGusul9tsqeusAhQ7I1l8qpAT
/adLCnpe4tGSbxGWPk4KWU0H8TeUZe/7RzPL/dd0o7y1OhJy/i23wvlDVm6vpSkCfc8JU6ZAFhqp
ff+v8U1whhFSuXeCHlCBsBH2KiUGG0+Qax9d38729jkIdRYOiWkbYjSyLWTpPohMGGyLad5IlZDk
WNRs/giuICH2TcF8hVIsqSMiPbCjjKHD1ChfOHNxJXQnua+b6hv9MNL2nKbaIcvjCILmJF8CvEmm
1HDjAb2FSaYFtSXrv/3z9DdFc76FEDwk2S4mu+QUePHESGeBux8TC0bkLx7Btlo+U1Mj0wNGLNIE
ZIH3mCpEgazkcI5pu7sg/5D+s9xqN5d1wLu0aCaIFgZc8il0FQ9w9M7cu2O9WXqs4Hzgl3X9WSXi
ZBLJKSh0Ty5FYwP9wTC1RJw8L5tMvFUTvhM2KDd9HGBoFeFtvvn5cyrutRN6DbDmUcnNUZCbF/ZX
z7cvCLTtxU4uECNJ26Z28vh1a50zNu+PDhXEtuYP+xoIedWQ7QaXy9vZym6PDBgJoFYMfslErnHK
ClGmZy1rmHlY3lW7TPPM9Bd5URmVGtLMJhVeBbBZjW+5w4iYgXiGAALfi9r2iMFWL0BWBJBD2c4v
WPXm42GuGba+JzbRkuO/gTgT6l/ZhlHtDAMJe8BuqI7fwI9f44N2xKCbLodvrkjc8NjDqytwywSV
w7YGcA7afFsqjZNXk9G6QT6LRa8EoxFO2U/bmllkjtznwWo5dgJ34FJmt1IwOGkYKCYznPqRUMIH
OUyBIc+73rWSrhAl3SQj15Jh1nQ72dOm8OkhU36Fev1ctpDHQS+MmS06eABT5F2K0vVolEPQZEH6
OGfad6u3s0W7n4jQh0aaompXWQKw6i4eKXI3BdXfJvPEG0dYZT7BDANHGCNCCrZckFtgSwR7B+Zj
5Uno1XQfyZfFGFaI4TEsHvhRPXrUeOg86vn2lmSpJxLjaFv1xTWzGDda3pzt9/7l3btbQ9WQZF6K
90NcL/idfljFMCfo1BNVAoCPUen5AUAlMWC6ybaSRh1tyIuLgR7qBKZhk12OzgkFzBm8a5VKWem2
geX+AHRNN+hsB+JYqP1WlTir7h9cdbClTPXDylWI5VOuAkhh1DJdYs0kabG5/ZEkk0LiXiiP9II/
jTjV0HjU+cdZUGVFkr72cVspZpSysWv5c2bsKENteOIZ2r2ESjGsw1zgvWvqFI1vMK1R2qh98TGJ
wV6FnNvfAPc/oeZs9BehqtClx/aEmUDTYTLqXQbFopUWalkmxUeJuwqcGfSaLLiFVBLicXWWTo7E
LacF7svAHeaZs4BPM3Qc+iy5djrwCwXCwAXeYy9wwJVW1q5IKhk7Sx0TDzCxfx+vJi40WSPEQwel
Xsp+9QHpVUIq4x+FLv3R+UgCbMd/2aigkqNG4KepN9Adltz0ioHLA0VJKD0LgXcDniJBLznOnTU9
z+UIekXEszT9/n/V1FxjDuXHcYGd0JbUSp8WscVmfhg5HuEF7FUhVrDNpcg45Ob6wvMHRJrITOHQ
i5l5EfuD28MYOTwacJdZ5C0MFypfTxXIxdkF/gtp+vSCDo8Q3aL/K9NN9wUNxV4FVMcbYroAepXF
oRzYSldz8sxMuBAXnXdRE5elUuzJ7pxaom7piEmZb9MhVTRqN6rAcC0HGgiMR9aNvZWbCMEbo5cT
fPA7juoYLhMVCOqLmvteo/u4sdzpfVOoCxBT6YuJzra7kiPJ5HAnWLKvnfA22ctj5NDexPDXamRX
VjeKv6B8112HvTthSk5+VKJKyZNdwemMnzQ09zKXXBZ4kHYs/rEB4DlalsyKq3/+j8uC+JDUM9Ub
YzvSSn721Lap1Kx1VhLdHrPiqWsvHEhra/ikW1NF7JLVhICN9Mt+IXiwt6uKr1GQ0D9CAYy+D6rC
lSU7yJSRJlyKxAlk6GZfnih1AvqqGTXihbPu/oEoyy+YAh1ikx/+2EIOYKUO0zMcsbz9j8PKI9Er
NyLXO6YF5ar3FIQO4ZWiH7zOVwl832PtgkPaWoK5gaHPrrf2+FIrDinC1uYq+xIf+e4zNV/NoRdd
KpcvVYR6lKcxryZRqZW9odcVOquLgXxmX6lc8sv6Z4oQ6+dg5Dg+Iamzo3al+9oJYe7K8qrKKbr3
WEqz+bfVyv26fJC8U3R+3Qd6CmHIY104ymk0gv7jtYOuZPs/ZItYrxcarf+PwO7C7pTaaD3dwu1D
3USeNJDwjTuV1NnWjELBQlAu43CeVxt2TA2DWqVoZUBRW6FqMs++wWXD0mLDiCIYT1nZPcmx+O0Z
fEA/hxDS2LCZa9fg+1JI51xJwg1rsztKnNNA865Emhgl5fv6SKMKR+sgeLlSHP75VY1NXwb4Uuu1
4sHMuIod8HX7qvOxLnW6Okmu/1vmFmKgs0G2Z8pac8FJhC3x6NBrkSgMjpr7y1J7D6Okj3rdW2Cv
Iwj31eWlWKUVW1s/BPdVE/r9sjg5I7YLSArM1ULX2G+6BljHHikNAQfIC66/E9tBTWfVnChKmNoj
f3WjnU19cfLOfwyY8wz6E8y0IElYC+0L7w/0RzJYu9/82FNCtSAw4KESRB3RQ7Xhogef9xS408LM
1MgkRkISLTU8Pjfja72qHq9WQYp9fPY6Gpmmr3eSTTPG+iUCQ+k7mQ2XQ49+FKceUM+g6VPrqtqm
2qV9SV07gfg8t3VNva+drfDg/82YNweWY+Z131wcwtOi16X7MecnHVvSXykIgQPgC2slC8S1HJtb
yXK1AViVxvgPkkHhnN714dxFuEz/O6Ey5KlRXMDDDOsse59m9OGm1u/J2jwINJg5GdpB0cYl01Xn
vQ6xuUzh0hXyq3duTBBZn8Byx8p94P6tcf1fFDhwsHEjAtXLd5otuFEFcNAT7B0FqBSH2xlv+zm/
I0PChfaWyE1DN3aTEkRXqKbgXBFqpIrLzhnI30Hc/ogNyp/h+UYpPCM2dsFgpA2bArSSmPllk8Nq
ysA1fp4k4Q1x5MQDqwwg4y5DVyTYwT7TtqFpb9OOPI3npsNGXeUc6+89lWjRvxVNKGI8G2MFcv09
yJ5fDjD7kN+o4xhnlJJhnUAFCoUj+fNXgUttWZvGM517tE9cMXkItyV6r8y6jsHR2NRDRu1Fyoqg
kIoux1jdsQRIBl52ZK4PFy3swODVNp3VrD9+AhiAXFPXuBlM/lIO2cFjo2KXkdhVOI1adw3vGFRr
8CtNrXHyhxV+sUvMHYdUQnjhdyfqRBrr1iuD8sl6AVJ2c7rbsDt0gGGWI0vJI2DQQRRlh7BEfSfA
leVSPkGmfZon/OhcypAjGJhw7JWh/X2cPYYvmyFohRCYW0v52OfQxmWYbainnCjNmv//ifEjnLXi
UL7kQogxJTpL9fVk7SCQtfLYKT5MO3t3nRfP81AkaOxyC6G5pPIpbHI846JjwnB3TV7MZK939506
XIk5KJROFKzXCSo6DzOHNabWi+97y2vWPw5pka3Y8kz1sO3p31keU8Q6aTPmF6xNcFL9haj5TnWS
7j+0R3roBCbyQGEB5kStkkr32OH9z1Bix9RoxStZ/eRuH1bOoMFSHaVW0IXIRw78lxYvYji9wMnX
DcnwQZlFCOgxdkj7O8H3QeF5PukiieYqxy21Sn153OtcOw66vSfWZ4hO/xxi8jeCQC9YtAmuTRfX
7/5AAZPXrgttVmO/0jsafrQtOQOH8MYDqNacli7IirksPfqNmpgTB0xi+2ka5blzb4Sd8sHcS8IN
qcrjrP21rcdMGXUACIVYB9hWCgCA6hDLQjna2NKMDqCYS8/dE5lfuKTKCI9TPChVVJ5A1LtHbrhd
NvBi+yElXnpvZToTefBCjl1VV7RWGiZffCt5M5O84FtYujhefy29nJqi9u9LHAyfYBcTLgg4+VOR
BZ9QSJUFMxVSSl1mSTZz6He26PP8EffFeC21uq9giCZUVd3UN7gD29ZFxYNhzDNhRf/Ds89C9mI7
+Z6hHAhBMD02Ze5wIt4vzUpmmo1Mfv3M3+RWQkS+tul7m50ZMR+vc4z2iAdcq4477JqjhWNJdCyC
ulMuk4s34QxsUurtQgGw4HDRf4ioDosOMW3F0JPDoajMbbsW+EaatZtYpldH65J0jyRb9vTQNypD
/UEaivrxPvVewIHnMW3mvWWuL1bf8/79MNUtTP5fd5e2Rw4FY8XBHSi3gc1J38ZsHQj0BrNz53z/
XzkmZ4UVm3u/Oa1Ba4poEiq681u3tsLyzqRO8hm9WZnZXm0yCYQiuf1IzmN7i8K+6vKVXf648IaE
4u/WF0Y1ulsNAKrkhx2jZSh69+3VCz2jTVtFtwOvZmKazf8jU6JuHjthk6qx7Oq6vIYcQG7Osjjy
SghrJxcS0o9QPYgXTONDv9JOFZg+PuHVrjfGL1GSL2ptQ4izntTnRYOXMwPPd6tw+EsaiWoyU5M1
2dDMpPpDLdGRjFWc4Xr/nNOWSm0xIuoMrqNdwlMDXh7RegBjMI11HV+4o126NXEA1i4S3S1piGOY
XZEtKJQSEEWACZs885a3OLma0x1RaSVclrwx0QpG080ni9qtDBedsXcqv5aFGtOFvODX47E51Iwn
k7hkQNfbeAzE9fBJCZBJgCwc4jHo50aXr6qGoTz+iD4xe3nC3zTqSl4rSG7jS3IIqk2Kg5mhEO8h
KSCpXMfK1gqisNEn5eEOzA4o8MnFMjQmWyctHk3P2rTpzbN/bRvSBOeTk9k1LSXvPMxVajXgiiLH
+j3a+8edVSX9/VlaBYrX2/D8Ho3MnkAYBS2Y5tibmypIvBIPTnBZ6hwZ1pMdCM42H2zbqJL0XUmf
EswWKTtjp9UeZMhpqIsNa3V1l1gQk6QePvATB2ESwpdz9wqERUPwMJR1XJxcR6XMmpbYkSbIh63i
UjB04dzFebz35HM3vNPD5045Is0L7AQsFtP9qxn4Z+vUpz2qGeajXHrGJQHI9nqQ6gAN40uUrTGc
bhKEtS5IT5QxTMaLi/Su9LQ96uzUr/SoIDP17ENmRoGC6etF2MqvhEpuZ6SZnDJrOfhGSoz136+V
Qsp3zPxQ9OJBqcy0XVzcv4INiKKcvp3M21m5CMhWxdFuZTye+vPg1tK+1upZPLTOPLmq52LE8Far
OSWK6E+NcPD/JSWwwxGtZ1gB9jpLaKoKUpby9kyKcPy+ENRvcXzAL1BpUG6qlveXUgve5G8NdFfc
iCWweGjd+isIevKljzAdbZ4wRO97iESCo/ZsZKwMmSVCMKe9oJtwmK8rBIjuf49LVf765yjyg/oL
hxq/VtHIWum6CCO+5ncZOp8HK5ZbJUawqIZniXpcGsSwkj2jyAfAvRni8OQyykK8x8dpayR4he1k
vkKEXxRiOIV67fV4sTedEXnSh9G+PE9ohY66M/hyFdh/GzqoR3vvdUSN2J4QQohn5JgVpQPaCcZc
Sm9WG99j0gQkayduVMmnOAo1hQrxmI3zTvQOLYMyni1RvOEew5FKR0NS7FYSxOPLGX0F3mEB0J56
5KarPHkDMei2rxlRKc+P98aKnZaE4QG6EJal/bVchaszloVHqY05ZmbxEAgRCrSMh9jddTnK98zt
9dAAwgbeFSWG+D5n7c05F3IWIQXA4R+JzsHwSyxmivQwXS5lGccsaEmRo28he588ZODR4bZiWCsd
RZnQJNEp0WPgvVjH6MD75ovOGOAUT4xLPFlsGBx5bR/lpnqN4Sm6PW1P99k9BumefmCRyEuHQ18C
3aQllWnHAPa9GkXEi8N1qyYqslWdYECSkat167MiGE6Z3MWor1JngpWSlu9p1tsRToIBMTu2RJLx
p+MOgVs3U6mhTFs3RCBdn7l20Wq059ArxUfoYVYTUrKPoN2JHsG7ImogqAbr9aS0Yn4CvbNDZZY2
7MMFPl0/1XCZZmJsyGYpNFJAumhZBILeZrgAWoA7X/IPHML3dpwXC3Cc+7Y7ah2mjP3aNIn9HwCp
vFKPbc6oYdyE4Ofz68c8m/o9aI3gySG6Fp1Ru98vmwnRbnb2oA512SmPg3Dns6PnAEAQaMLNNRRS
23zBEQAsr9s+RJMRgs2ndtqm6bSFxV0rMkF6mwwrGrF1jt8dgG6LfwS8l7NZ9eQeo8tBJqsIstvg
YcZZR5JfLX6SWysX7dqYDWeC9yV/D2eqJyX69JbwpCMBBU98K/ugy0rrTJ0WeIHlTtIOFXAVbcgo
VsRj2LmfQKwgq1eR9iqZVU36krXSzLnYl8KclxqmtXKhP/tDVtEvqBNqY7wkEUpNa451hJWXWBXK
sBfbeHNVkivDWSU1+tj3D+LwnykD7z4qs90h63LxUHZOQ3TkL+Xxcl5m6S9LO/vor36LDSZyN0c/
HVxn0AmI1PAQnLzZ8tZDRQ0GMLvX+itoMlfNnZ33SxvOOvURPs/uSI9ZEyFKUil7pYUHxwUusqr2
XT/x4Pi6sfXhpM0xXTsrnQr/ZZPomYt2eEwDvnIfein6lCiPbMC5t7HQNTONcx33vKc0smZO95QC
7fCRDPB31zYbZclvMievRNXqZ9AzmaaVOV8ORjridOizAfqPOjJ8CwRkH2pZuX3hnCjFA0fXZ/8p
E46/jaGi1uBv57xzjUx/Q2vZrj4CvJUk7dgyWt0hQBqx3EsO3008F/aHtpRWIx4reIyLMctQ/VLY
jIprV8GMvROnLCOJOP1JmZ2SNLklU/OWcrhu0GOZHH/7vI/cZBiT6BLAdOXyQaROSnbhDjUMRFBH
zpNSFrnKLDIO6OVxiD9D1CkKB7DB3HIHLQiXOPtz0OVzim8+hQJokZuEKpOYwuJuKLU72gEyiX5V
aaEVSz0EyS3i+0AyVhkRu3ICj9OcyqOt/yAxom9S8z8mkTSs7IY+sZfMnsoOmEJWJ2/Et2KUGJyY
8pOgu8KtydVffuZ6JI0dILAKImkCDexgS4MUK2i7lXqxJJsBAlxa3kKyglf7fy56HkdY+00ytzeH
xQOkDQfUAbgOzYqZCp19j0fJS9uSEeKciJxv8OD+QdWDB/DP4vCjQmbpEB6y5VGjvU1IFUqbV00D
fDPytAdhCOCXRWi2zq9+LACrtTeCwdFUWqXkC/YO0GY0VNXNNIyCXs3WIMHMaO/C5Nt2BZCDAvms
i45XgnqeskLkFzu3RtXQjxFOpe4yEzivXXAr0+joPcfUyeOEPL6aPfpbMiCKt6SdIlIA9vB3LVET
0/8F4Wwytz+feDZB7Ntrw3QU/BnmChHOGYOmgvURlQnzC7sWqXAwmGpvZQ49rLoKCz4gS5H6QhiT
ONszXQmQKV2GytHzM1y5atJRk4yNzPUpwu8nN0SVnII0gOh2jzoPnxu7JL6ruRmySojFqhLyxIyo
Cn2LYG2fAVvZ6jUiVUvfIQ6Xrj8StU/d9R4DSKNhAtvd3m8UBy8LHm3nsiGiuiVNXHfWPfT2LwdJ
ujAGpAejy4fq8Op7qitH0kpTuslCTwm9Ewka26OIZEwXiW72KbT81cLcSgapNKUbrorFshSF9yzM
MFKBYwW5SulnAmxw9c40wVoaxXVc0m2pW42tlsb3Z2s/0uFhxyccslbklsXAsefPLO+lUEfWmW8d
jAet8PmsENMP5PWYl6lPtids6RefPtcf9kpWDD9xNlrm3q0PRESEZCRLgr59yoHnhQlp1JZXNsf8
3bIzvR8kyL+wMamB/6PjA/ImfDXZtSCFR3e5eTwEPtiVUL9ZflMo9IjMbfWLOVDsqvljFw0b2kJs
K6TJKV6Rx1r/e528d/JwzP9wzN9yzmUdJdRBO7RS3264na2mVV4WCDI329dEZY7s7DrPRj9JMD6d
XsknoghW8vo130XpmM4s+fsLSJ0Az0h+BDmn7MiqALSJEHf60xa2d+hJFiZTphKilGnAgQ+2rJUk
euYMEIYlm2SyDqtXa0g7Lem4X+nhgBKjlZrXjaGU/7XlhEme6SzMGeo/4Zp4LhmHZxL3rQx30x6T
FTjOqiMvRixN0lt6h8h7A7+t8L/VlBrtAJXGQLty62+ZuBoTIC6EepRkg9xcOghTN8jyh5YprUgo
ROCSZ4KciEi5V11JglNpmQlT3U9UpC/g8ZwY+V8ppurBJKIV/6EWY3W4QGpe796IfEzmcUIpM6ew
VYSN2SvkRRGmwf7RuStLgPNkdzChXvYUGMt49Ei8Sb/SnT70Rl3NiYPxC+HHuWa8bqLN3B+MxwQa
Y3UGaUsFMZ9tzHixxsZD5H+JROkcDmGmUw63DdQ5WWNFfl8D/vi+4ygPeb7IEnGaBATtbghHyioM
e1jN2tqTX53kOeKaZBZdq7Yn3hxPlAF/UNYVUIOjoRGQyb9RcEUol90mypMEqENXRS2w0/f8wWb2
nGlEFE85vRC/rONUeQdHHhCzrvTfL8nWe+vj0DH32JyDv+xpmdyHbMsb7zLY4iaNZH7wFtTYoVSD
oGFlExL+NCdyilYOf0iNv8MbjM17pfSZHaUz5/g6adehwdZmi4JxZjOx+dc0H1M6TE5puGFnpQ3Y
dLoXelg8vkPFoed2DEW2dQBVJS2eXrflQS5Sg0/hRpbCxqw3vXe/VFbRN9vXZ1RkqwNcHlISSIoq
XPR+0KPUCENwV4miSxKW19Reio+W0pf5ip1aOJT5mSKVs5pZkyrayILZJC0Qb01EHQJHuo1r28+R
0HWcDperSEECb+1ZuXbnRpBbKyorI6h0II/AgOZkpf4aK0UKvZ37oEQFG45ISGI5TJW2JKKIIg4U
HWIy4bmOYjbeBkOSlB+fxmIm87jAvcjqDh4O1QS4bjFO2IeKej+pik+8/aeE3hxWsuLItdiFpPry
FLbGnoy5GhQV6VJs2/9hh/NhUFwd8sKqADtHREJoiFY2RMAncNPKQyODe+Ag8UhyG8fieWaLFtLy
6/jDYv6uiGkk2LmJyaUNgs93qDAMgcM3zub544cFyD2zW9lJtgtJEyZJwZl4hUdFFl4WIMk1II7H
F2upioR4a4BC5RuuYiTW/724cF0+u4GX5NV2XDzO8cBrPGNe2ikjuVoEjy2hnjz9CMe1ioAUMh+y
IOL1DcxIdifGAYTNfDByWPZKjO0E8JiUZbx/BMq6BYxd7CzHJZRF8AorpsOruSslr4DLHkSyaCnn
hG0FxSNsS1KWpGySM5J+3/G7kSieg99Lag3olLhPp9vNbQmCTozkLvG/s85XTlxUhqDq/4XXqqmS
xyeHpMyfghuTFmvRYDpzo0Vt3cAqdS39ij8NaNtTr+5p4BltYIL4V4lHgxHjOIulRVhpj4Nu7N9u
UGHU5i62DhnjjCUeOtgO79bQEkM98mZrG8yxyO81h2AaF1w+lkpYm0jnxGBjoHflZW1gLlGeTqZ4
X1xzMV3+Oic98fp1rfcfhU387mJ5vhSthaR/fRlR3NmLNSopdYucnlQVpOLPVa7XzljbkBs7VtJh
is/nYDDCakTDByO7VofbZenmexiJYb+hGgJQwdYB12crzf36FMeG0G1VL+rpOxHE62/ad74OZnwB
nhxC3gJKQXv8m+d4S901TkjG1tOxI9/owuyyLEV0fWyZt98zLJiA633x5IEowz46uxw587vIXXf0
9xD6uH9+9MVH2ui0o7vDQbtgeH1VKmWW9ILtsquUc0HmBpskpa2O0hPvuQiNWL5Djh3VoslZsNXL
5F+98QIb5AVCOKeHVk9PSxhNrnEpw4rvCFQvCQ/eFh20JKYB4cGK3MnlWEK8bISzzqBVG650fCMJ
5nsZrY33FSwqcphvkZN3juftI2It8TpAGcQEpVK8nnNMx6gnBiWKT2qlBaZ199K3/W8e2pVbluTd
2lEGvsXmD2H8Az98C5MtGkr2mia8UDji6Nl9OnHq7F/iE+3oXhj+qZ3AWLrcWKthesAllh/P4uTw
xiC7d5fCYbhGqJPO22jCT+1ihvWf67x0yeQJdeXs0R43ePUjtWLPvlbLgLPKsbiDwqeK5DbErBX6
PpVLDTckFK6ZNTRQ8ehdhCXhPhP/2pCmMv/J5PmeVBlRXwWOlTeuXEIVBev7VOgPc5BMsV655ew1
7L4XkRo1leRjNpxgLrpOxocJ/JYMTGCQqOANSZI6AFEf5JPD4UZ1Hr0qlPSpNpQ40/4nus/YNH5+
itxz2UVVnxoj1yw/cwv0LRoAjGV9haPcZXizG4tLza/32aS6F0WiiCBWzbBv8rmfR+yAmOUZW7XJ
inuOpSGQOJm2/PqNntvyIqvqy71emliSdwnWiXsggETALC8VRESsAoeUMbI82OEEi+5cEHsC9pFv
T1W4c/mPnwGZtEoZ8TJsST0CsEjEYMf4QmywcAf5N+74FA0w6VyG3FEvxYlHAKk/LzJxNWIy55ov
qc3KT0KegODALNEFTFIjFtPONWcYnUQNx/McXYoC9sXHXYp+s58DC4HJwavItwHN27P8AQrX6LbA
QcAZubOe99+FV+XN4IN8lTbIkgxCcuPph5qec9kPyObmx5zwb12prUssLe5iOA9TMS4myr8t1fdw
F8GgpvdOkwkRrDPuztn7JRMpJkLUYs9hBxUMCYzyWp/GeDWomEuV3GsSYHTx40wgtT/yEKsesTmt
yq4w7CQb/EizvqdUbsiIjWGjSn7xq8GtqinIAtHSF1XY9RWKFzLXX0TeYiTGJjRECmgHIjvW6G0y
SseFJFNU+S2BFVLDv+i8pzyVFsOrOhvTKrJ+OQrMTkROmJIsBa3ucUVo5TlHRvHnh+pZt3IdxWRo
W2BH/A32Oho/4ockn/ZsC4IOM8N9c36F/Xht57ELCc6bgi5T1myMBOKqy5YihYGkpDzKLdTbyv+8
cLjtN4J48ax7i9kRhdIH6PtzPaXpHZX1yyD0BPhYRGhvbYV2VhuRztgwJIb1aPDeuuGxGg8ase2n
El91kvcUhFg6x82LJg5eszlmNZtCSTI9i5MyqWa8GBwfqNED08EnnSAQ4K2so6LZwlB6u3n+FfaB
6/6qPgGr8Bm8OX0ie7tYGqi8uLTfRH+HH5Jph8sZsj5s1MJzEwfvI8kXb5Nu6rTnBYSw984GYcSB
lKEsOwLTGUT0tZbLi5INtjdm2SCgfSaRtQbA49R2X7+/i7C3dOW4SWDI1efxXdszXhO3OdHwBpeX
V6RQroK5Y4Ck7wT/ra/VaID3rBNkyVwj+0QTuGJd9c1p9xCRS95xD55O++Z7yZsbbv1ochoKwbH6
e2RmYFwVjkj+MsX1s1vs41mjvYYpuhDjLzf0NAfEO8GPBbcg2994X0XMqJYFUKsqNzrcnZpI8rlX
aeKzVPwMC6NTr9Ol7IQgOdRZZqS416C0wObEWDS+5p6OzWOeGKnVUFExUE5JvCasZAw0DSIQ8Kgd
EUUhRWU610V7aNgBHLk7HdHI+uwbnu7EKr6zxhz0GvsRZubtwxW12MJPTq5Gzap3i88goh3r3npD
8rwTPnrjekN2Bh3Nw4UFfFNKgZU7C2dEzjsj7LbG1JzxBFNjy8Zg0jMxqrI8UgFexuqKfwwxzd7u
0sBe7kQatJt6xJpfANgB9/a9grHl43gxPZisKmMKFWm8tbR/DZkiYFb+XHufOXLdJSyqyrogCcQ8
hGBL+CkVdTUlhMVI2yLjYTUS5V77Bsaln+pzY/AXTjSq83LoI26TwDbWhXaMM2xOgFr0xHpVVfjO
7VZWh546T1cmJUWq3tWbzoagN8O7aR1nEhCJZ6TqYQAv9OoesjWN2FSr99lPCTxL3l7O6fMvLVeN
dcpLi1fUfExDlQlYdYv412Y7mmHZApNJoGyjZMQi1htzjqg+Tve1RE6XuWjN1H7K8CiKnaJpzGWk
JXNtG8d5Qly9rzN9KIYbD8q+QidU2QyGI8ghfmFLuoNELKW9UH9FG1Ux5FfSMtJjuj7ryYotvvjz
Wz8IsNtlWdFiQpJbFvwBO7B1qTn3pLK8K9AZWYvlEfleaalWgdTfitbIGzcMiSUehYmorghYqpry
6OZufbKNPjwfo28tzcWhQQxXqayfHe0FE7P9WrjCnu6DXN3faXGgtRFhGzGurQV9coUdNRQPM58n
RSzUNhpjLXjKFEj2IAZ5LtszCVUdMtSdZdPyTteyHN5pNWM3CSqEcHZd20UlixVAbCNDlfrMyaAQ
1rdpM1ROkMIvxVG8dxwO6MMVMDHG2nt9K1bAU6H5siIBK+Tvgs3+RBjP+oAWDhdnOHiMSTSbo3zc
Zpk89+GdfMXY897F04Y81P35JD4XcEKsAFtl+ZFBCN0An4msUh+LwvHlE3M3vjQWRHnzi11dL6bt
ep9zfqUce3NJr15FWDlXBr86pmP2jR5JXlJ3esyIm5gWGsosltTXv5n6hzGtE/Mrj2w2nDpNVZP9
Sthak1ZXG9eIQZEkYDqJm8aTpfaNUZ0fmrUeFVb8gFgqXzFLVv161uVZRvmmtTCMxV3WeNOjzj+a
exBMifYTi9uwfHUUBImp9gVHcsxRnj1YrL30Ijx6za2H1M1fsfVbESb4aHPnO6wBJgyO9WeQ8XLl
s0wqDhhQdspy48hc+IE7BVYFIAkc/axCbZ4+br6Atb9pPAPCEfxI1aKxuihxrhlqf186Wz75SB10
OaIZ/gwfXc38LosAmZn+KfSju91GiImI02+m0LiSdqNXtl8S3q0T+jKGftnZAGp5OtUmaXqtIdQQ
hUIp4mmgSbvPEkugAzTndtPcI5VMY88bG9LJ5mjPfknwvcVkxc9rduGlpIdlNWEIXY3iJYd52ux6
+k074h3YWQcKdbncNYD9D1Q8NwLy3owd9s936+GQlHVvf/YP9ELfTWThOooD0j0MI/G4TVd/vrVl
fmUWGCRoAt2xCkVyt1BdSErRvcgFu7Nzg3Mz0Ak3GBvozn+Nr3F9auFnDHJvV0gXS+HHv4DTE7gH
1a4w44LS2j6F8PPtmJg/acCgpjnmyFYX/AnaO33GSnl+eO8kyolWYtEr9wLSI2mDRLzc68EVcBRD
D3V0CJZXYkeAXgeDAGlFoxNG8mAaWNTaGrliuyC70vkphdIo2z4pCkGxQQlJlYIWYeGsZsO1MRk3
x8+j8cf3WyDk0WU86VG0AsFjIYCWScfuJ+g3gKSzmwD8nGQQPWiZNHxRXmEBpWLDzGAHTzDB/JOz
oJd2siSYazWRYcj7Zahb/HiEWqGo+sPnL1UwHjtyymH88kY//ibBlK6sHN7cudz+/1FwrP/caJ1j
dr32dV6zkFIvdB7EDZWVmS7Byam7Rrkpc36jqdPyn5nikgODXnC+WdR4msyQqwg5gGoeuJxTGsvU
YXiYByELLR86lZtbOxT+aTL5PgqVFTr/8I+egQScX531VBiQoIiuy+w/LA/aYmCTZ/Ds5MJM0N/e
a8DDWSpFlNvIXNAvipev8uuaFgjrwcncX9kbNSAabEkSgXKmAIgDIH5RRLYphiXNc5m6Fqtz9MMC
ZN1xVN2kD/EcklOERkydgA8NecTsU06xOI4Ie6LoIW2ZLXczL8NWhxI0KudE6Db0gbBRskG0BO/P
fPYcUznK7p+p08M6sXsqnz8bPpbv0yGqsbxMkD75LF+4P52y4sWLQUDRu0QubS761vrk+xrtyY5t
ikNDt5e+VsaP2XbrP0loVJYMlXVUUksuYsAHYgr6N6AMLRYgBzkbsT472Q8+xRRpU3gznwNBoPhV
mm+Qo7vSGFj8IupGblipnLkpbvz7P8a7rOH8oaKgwM014/+1ehb2PGVoER8oCKOXDdPozQIiWWpc
/nhW/8Ly6ODGEceQoErYE5GDwgGrbgGy7UFfWUbQOQb8nHonZwmIbzuxxie3dy5RHbmZs5qB86Wc
bVWX81toH02ug233ecbqrDE7UTley/AyadN9tpAGha6bMgxFqClt99di2W4C/CwyNBiRuKx3SQOF
Ext41ScpZZWbjNhqBTGa0PyzMrOuX40ml5Nc0kyL29h0MH1ENTFPttjSV49ia7PDwWjMejuC7rjf
Iocl8X8zFvzzJj4f0WH/ZgR28Os66vgvKSCYODxg2n2WXq0ZkY70kBSyqKiakjXB8Fd+SmFgheCy
1YQD23sb5QBFh2c7mXg4e5YkAfMFURzUsPtvEhHjTzWcfRsVJ7iGe2tR5ZCoLnKBJeaEWGdkcOlj
gkP0sg69KHTUW+6Gp6wxwzAjr1gReaT3ZzSFdRnRX90U+L+DTXO6yabyMrJCcdM68n7ndTSOpPyy
BHzN434LQS3BG43o/C2ZsR1UqkVSSn1ekVkDI3p77uqnhjOAS+MM8VhgSfKPbQcusBAXyiGSa0vk
dr3VK4niJSQb6xJz7TXgW9KYlxh4kxbVOjTybFamrgzRCNygRQ+ghFue4T4sEes2G6Y2Q/s5pi9a
rhCmHl2PzUbhvrCJ5rAGBGWEINQ4ipjIR7xQQAd0iHDuDOuY9A8kkO72bxvoOfvjaJ+si0e5I9h3
fQ5P0peXbLXTjzvLIqdfJwDaFalWH7d7bkm8btsNDTMjBJlFddJKUYLpBKWq6SCL5VbyFDmvGgqQ
4cXMM0o9XzpqwMMQcvI/schqczpkSa/7/ADk/MRT0VWjCnRJV7krSrmDAmNX1fuL4mKF30/IXSpM
xntEm5GCzaVrhQzK81PF5ikzXUbMd8AZXh9OEtnIzCkRNLqz/jrrs40rm7AB4Gtrfhx5VngBBZjm
TTu/3QDx6SN0b9tgca1lpCTAldoOZYy+sQ2cIUZhMFMMQbD4EWupgGN2MseoScA8nzJ+gdg8TalQ
VTUFmwpdck53Z/LuBp8pIz2XTkdDyNmuFW4Pm7/NNEeRegiktG30ozzTdyAbPVfnfZsmfgKdGhbg
kDmhxWsiJy/WDwIlo+jdr+gkOTAUeKjo1dQ7BdrPfdsqGWN5Opjys9NMVevIM0+jL3BCefi86UM4
8JD77JkBYUxmcg8lR7E41moN0ldEUnPHzINMeKQCQngmZL/O+1b8ceod4zFb/dVinQtSnUSKMoh5
ACNVTYGz2KoN6fNwBJwRDdnun8dwjn+bRTOmTsarcZTd4GwsKdI9SuMUeJM3OT2cImD0nOlYW2bA
jhmLkDZDURkjSSyHGaV3JVJGk9HMXdtmgZ+fZTxY03iCeNyQ6umgfLCrJHGU1+TWU6aA6J56pLFR
t/I2i/8K6EJcvRnTJgC2N4IsyyYPaJZA1/Hx65pEsDvbkF0YunEHoBb1ddn7kP03tM67uSnAiooF
+cQBt4mDCkaoXWdHY8Xwrf7ljiLt/Lp73xjgdGkRaA0RIu5D9GD9aVCwBH6LW+LznCntBJgdqlf3
heEOyjm8Typ2u3u9Zrux1tuv6pTtXRoCHqG+s6exhPn/Xad0TdEOJ5DqGTa5l+cbaRko+7fW7BeK
6sSQKdxgEZx/Kdm3qL3T6YzlPjkzXJ9nVjn5bYorWTOH34Jgq7mgL21DlX+YNCqMTLk1mXVxw7J0
9YK+54VmXOSLtoi5EiPYtWONRA20wYDCWbF4YA+VJIqT5j4YVae7wFrS8lXzqsANJFtNKreoSH0Q
vVgIawkBOBBZOvWRePHRbCbq7fIyz80y000v2lYHZv/z7OkcyNQH1OBT0VdmUacEAv2QxHT58JpL
68nja7XKFBpPxTQXchyeSggTeWGs2/pxrZ9IJET1yb8ehyvLvJTCaqsBoffW4iTM9h6Kb9qPDNds
V+QdDbbzfoGn0nEcoGKqfmM9PSLtUaAO7VCsoFMutUPo0VT1gYkHNH3FvVhoeFPHw64ZlEPEdQi4
HSvAf+1Opp11XtheZhc++Ho0Jdwk1KK55HGV7xRvubS0LcT+7w93gC/6cVD77PaSernoT5L9qeIp
OD30+vECqqgVnD89yTdswpo16E1RDOMayhOFWTXSXHjVHRKc3L0QeSxPIg0pkgJIYGF4n+7WJYry
WuMe79+7KmQXRT3HoCbXnX79rjXfhYybjLbs817Tvb+Dd9dOOZZoLMJjqK0BNND0WPKfoh9StB82
LZkhcSWDENSZphYQqlsKYMZ1MdBTYx5oDzcupBgvmgMggHLa6sYyfgnXI1VsaU6QsrXoFNiHco5c
BUo0B2eW+l2vu2pdwtBgHRg1r1ZLdUSjF7/sym5dvJzBoMScjvSE8AuuuYJEu85lYF4fR6VZRSDh
wYQ3e9kVpkshq20O6WVg1Bv2nccaGPgZae4hnsDnUzVzNlOuQZw+iWyz1arzqPB8jlvFkOBlz+5y
5tyGF6BgxNTiy+BoZh3H+RxiiGDyADeFqlw+VkpEtMCsNOt3qwsbNjq6pkIwD/8Lom2+FMgYcMpy
zHUffqJGdsgHxgvV9PA8dFcCZwxYK/eUCAsoZ0ZiNvsOPbus05Vqr42mM5LJXXb9uKvT/UvwjzjA
s2bfaA0okxmK4IFTy/xSzhuZ4TFEXuK3g39FoBnZWKlMvOLA2xluxIi7A/j7NRc3yDu358q2cJ91
qEPKWogsQuEme+f+FW9KfR7EZIHHLKz5OtiAy1q+B0Qxl2dT3cREY3mfp2+deNfFOweEyS/W7xWP
UrzDcnpRvySAZNEVD4CZ63dbE2HLQEmggGp73sxPtER7WErHR3q+yZmCwhYaro6seeqCE0N3wWx5
F6MD3TNP17ict9foutOl1+pQdnpkqCAhGLUY3XaOzmEdWPyEYMuzJyBm6WfCwsHzSuo/B4WBlzPU
1EIpi8dwubhWlMNvWOAZo1M4Il28i+L/ikQ4XxaQfleHnxzzNJJzZhQA7VIkI+tbJKGPHUWIPhbZ
H5iH5sWvDxmuBt6aSMHnUVUzgAJFIuaJ0e+jJUYxP5Psraw8zZ8NbE0jk5suvWT85VVX00A/N2hN
CLEzhwpBsh7Ujxvm6J6gJ/1rvmp0qp1f1Iq2vy2/RZH/q8posb3qXJi8lCCYPWwpaJrJBAvCVVxc
SFpuRaMIYZ7KwFrhS/bpH1em8gQPD2tUdJt1pMBf5o/7JqiFCzNxwG2qKt5eAjE/UOg3Dr+dhp7y
6CDOtTqoiXXHJjSWbioQfidNy0loruaUrAoTGFnOSW2mBSxrtX5Fd/PXbLsK/TqrOHuuujv3l9TI
NZ47oJPykJIYN0CI6yWfJCibsOzA1Oxe2SOfPlOxGlH3ofVxOqv2OuheU76aGoD8hft+OC4gO4FH
DB0NZK+4BroNB/g9DbieNZS1f3tpLEQMgHJ+IPV9wq4qDL5AKFnkdmA3WxA4YAjOGx9nIYRdq79t
QEpVplxQj4FiSbDXMjxgUxxS3R2l2H7tm4L9PMXc21VNLZB1/YCUCBC7R5mYn8oOFDEuDkJOyGm7
WHoJsMpF6rDh4Ew77dM3edfBqKWwTR3hGaK+rAsen/8VAw8Pj2t4E8IwvbdofEFZwJ2ZWH7d7fzs
tpOmiWTaUVUWyOkQLXMBsdyqje+LNtYL+vk4CD6N2ywuALxU69mTE27hQEvd6O7lW+Mkx3znIqzr
YcKr2Vp1hB0thRdjvTr8T2920LUf9cHe7wLjxXFq1WW950hmStrMWMUXUUure4mHvPp1f1qC6Vha
xjhBsD3EffkjZrcKPMHC9yv6RHCzaNpEnxprLu2I001jYnnZ69uMh+tfntMgY8mrHOnlmejjLu72
fs/u84ZIW9DBthjUoyj9wLcm0WIoHIyxqyAm5na9Fhl3p+x3OXTxbA+hAN0DZaddWfIIgEzwAlaX
AhJJoblMQYcfdlx/vXFLh5wYNACX5A9lfqMbcZhUReia6tXySugPYqdQkfNwovoWLFnEy0Ejw0Eo
TcgvrUfdZnEMxaZdovVLfEmnBB0jaAlPNaFWqSxRk/wwSI8vw964+NoFx121ybJ9nO/G7hXy/XFQ
rDJPfp1CwrgDtbF+8DZwIK38jJ0jGkNlLqghrujHnNYd9NrVF8JYeiEgTuLBczKrxiyqtS0iY2Qa
+QACv1FHriYpNUD/sIUkraLUe0WuUjJVVi3Y2ev5eu23BhWSTxlUJ9NxVLE8g6sqfGxaim6hYSE9
HgHDYWyf+JD5OKzeCpEJQRv5DKBKIOOJE0AW0QBwoRsVKYfRat3Y3p9PlDlNYrwI5Dk4rB+QHCmI
t1py6wJc246GgIc5xOHOK6aEqQVyKhaco4AwaQgHUjCI6dB3XMKN01nlkmukqSXMmw/ixtmN8Cal
ssxb7YfQESVTLiWjX7hu49qdlSGrz88T+FoHI6J96tc7Fm9vW6QBqSvP7tUzzIvyNOFWDj/aZzvM
uFPE6t6hsa0Sdb9a3nD2fPr2Pu/BegoHR93GvH7urUi9DScJnql9KCBHfP2ODN+AFAGrvBXIoeRh
5vGBf66526w/OOV3I7SFwbBdXr0zcXdusodBZ++DpyfqQ3aKpyZ3/AwNqLPdSP2Fa7NuDNrD7QRO
TJa6rSFIeSZVzgrfWdQ3syfTKpj+l6kZ2gElc2xyh4yPiJSiLNZ59U69ThtnsT8cKYbLQVRw/CP0
LAV0y1s878mPAg7lksQQi4nMTLycjTisDeoYe49p/U8LHkKgMcoSSRczNAeTErFYvTjCKiv6FFxz
EqQFEhdH50DFQcjeL9DbO4tEZp/77C+TPM/B60DfESJPoZkO/U0rjo1EMcL+f6C13gBepDvCkdgq
0CXhDXGhzoqvCO7EuUzr8YxGm/Y5omP1HG0tqkd/0u8EkuniGW6ahMk8/l/9TXYS381OVYGCvXQR
OLL0xG+qTj9C8BwoXAbgru94pmCvqKzKMQfRKAzU//jmUo8x8tJ+i+snfViul8kK99Xh6rloaFkB
uCntFf6CzK4wHhZ+2hDrFOsGWpphVI+Qdh6rzy8AEUHqA/pbAJI37W7cwouFodbSNU44UOxtwIcu
DoXgvWRJnKtYXJY6PmJnEM4ZzUFiqv++88Sf8WFPtAHQpwBlNAv204uonNjcLDzk51bATg7ZbAQ5
zRvGB0dp9BiDL3XTwI0f87MmB3OF8jGVYCGRn2shHmIvTv524pN+4A4l67uT0JKXhWMtuWuONeds
jrI4rRDhBrmDhCq7j3AhX1Wr8LqD67CiAohiSxSZRXbBw76mIwqvm7sR8mHPSdHglbl1qMlTz1+x
CXhgHAkNLrWhyKrq7k82LV1sfWIDJU3AjwfCjN3a/pW397uY9lErNQwlYc8zvoXFSyzbTtwIBaRX
74gltKAMB4QHA6iHPfwrqVD2fcw1ydwOMAGwA0TUIfGnGVZtZQA7k6zwuwmj3GqSx2y3FhJRvK5s
N92+zwXslonVlFuoGzX40mAxuva1rzuUetMF3rrYgi/FDzsJDmcInGm/5x2hzeUeH6XDUDE23NtW
wcJyhkEtkyjZ4bMFpHegFh2sycfn5X4Wv3SUlYb04K3tnHEh3dtJrt/16y8X8mB67GiLbKHg0kzA
0MAvSOsimpUYo0clVCX7+MFrKxybyFkdz4jeHvFTaOxCqsSg2czUYE4EUzgyt7CBM7bsXvD2ZF8r
Z21czZSUI1aXcDDstd7p/aS77WkSwdLpGlj9xLPZt6Z7D9NGQnJfyXuoRKcKE2MS4ONQaeRjhnim
GwfbVvQK3yZJ36NpXzMBg9DrVIsLrnLJpBDzPwyIMOrMto1/4JtEPRteMgo7I6dMMllJzf/F8MAO
+2iMBnuCrpYfrNNWhMo5vkOQuYJj+au+O/FlcDAEjTgOO4CTgghySycVahZmoCEqzVnz1sEsKEyy
DiOdy4n6k404Cr6DkiINn4DL3hismKVsY0GFtaKs61dWjpTSMTan3qXVVBhsS6L8NA2WFVEObcGo
gFSumhPOdqJX3eiB6P+5BUYxcqVbxOcJNPadPRY6Eas3MkG0Bq6H/uWIHK5Fx2ATQoeyYzg5w2kZ
wKHWSBN3CRTXDaYyoMcnfEPZfTkKGvyCCgxwTlDVRHffj6ngf8AAZHxar4jU2twytwslyprq6zpN
zXMi0BOR14TizCNX8wTiqEeIu7hKwZWAIsDaRYXnQyJMpr6r7pLK0PrxoSYhc1MIj67wE2z+TeBt
HRd87wXxz1jEFKXgcPX+b3wvH9YKEu8LuShuFgl+ZP3tqnhCRb4+x7GguL4N1CsMBIvhucF8cemA
uqDEnB38iJZIKEb6awOGMV2bT3bYlZ1KecQSl2M8e688cGQlTM/JqaUvv50anDHUpjoXyKeyDPhO
b5HoLl23I1EHxhxJYndglCVcbFaexX4r9sKRebVLjJxK7m++WA0lXSWR7G4w2Oo5HkGAdN/R0lq7
kG2ya/kuXAQyQsKOiGIzDsjj5Rlnbm7nSI/N0mWrtlxHX1VW2MacC9CvTkMb+NZJKUy1D9nwuicZ
7SLjdMAKLhjxWtNfj4mZXvUcU+U3irJhFCAGapHJQJSbOs7ezDQ4+wYfu5A6rk5rwoVie8+XCPjE
DTHh519dBzDvWXOKaaK12mYUmrXaz4amHvn15Wih6PiyXSl1i069rRtoSLkNa3mJg7cE49Lhcl4v
xKMOH6MymDmykp3AD6P4zX/H5QjZIR0dAmkgakuagK7tLuI2a4DU2CMtqKkQ8PNUBkB4DHgPwweY
/EDNSlK8M/aCkPUtl4IwwZqkGP2ucJjvXnM/o+F1At+amsEj/JVRLCx+uUEH7lrKN460lWq5yweW
VqDdo0UxNMaqQsCf2CzeT/By1bbb0SCS6zkaI9fLyMQOBnEEpb3392venbfwVpTzrYAAxWbfyEHZ
SSlXzggXfpMMEqA9ZHQ5qyZDg7Cfnf343aN2exwdhW2duPJ29tQ2kcEVZOqhOaOe9qkxkmFHU4Y9
0184/yOkZK4nOOi6lYV5/JVtN6ia7x+PL0flso3c32ufyS6NbjaqS9oFv5o0aY48oeGDqq0J1e2I
pCEHZ6LRbOMRWFO29zGhkwYAMFn5JrSE9eTPxZq8L9CRjk5duZJE8MCXKYpKXTnUNAmfsteESyg9
qR80b2/N54/ObU25JbHbcSE+5hvolbD0avvg32ftAL0yr/z+JWh8Js1KdEw8yr7nC3SPz6od98lm
5w64t4HcBeBZ2iCsOXVLrm53Klblh7N0RmE2FB/+yZIzDwAy1XlmjWg3qzU1twGoCIFZlfgf9ztw
mftVEvRNaMGOfBgkD5iJhTXjlTZaeZ2igLHmN9IQ5DRAMCOwxUO3DS/+b0jTq3eYhwCMvdEPVs3K
HX1AV94ama3oowYfi5KXhkIogfIbb8Ip8a5ocrMlNPsFGNAKgRkM8THSOCkkEeeTPaCiT1GfgB4V
rt9IA9BuEQqb3PGbgZcsXQdQ0GBEWeHFM89ns8mLCq6XnclFKD5UXGBt3zn67iY4PQfFeFthKRoU
XEWtMkYNJB+FI/7d2Bx/hafq6Tyun1ly0c4LD3ctJyYv+B//OCDkoQRY7ez35qYxk6+Jpu25S0fp
LgBjyto2UesOyUWBWcGTamua9UP+DELEqoWZv3kyhz9qqCCF79Fo6kAHVx8zLJzbjsnQDNpFnO68
OKrjU0x3xPT8SpxJTiiKI8WlkKIWpksDIHQepAUe7KXwhEmudz+lMAsl2Th4L9go5Pcr1b56IyRu
H5Xh7EzgS3rxAgu3AJRI4d6AjQcKIlkvBG/9FiGUmfPaso0RE0dAX2bRfXRfBb3cVIje8OZQoUzK
TDgs4U+rULZIL+Ai8Xrrm6Yq5RjaSZVa1SYDA7WJ+2mtlYeUvIemMQ5Nw7nFByJHU8It1MEo/TUA
pWpgZJxy+4RTGHA7ulr4iwtvI51spHPyLPFFLUIuspUTOqLgX3cj9/v34JdTAn4fgX78ObIfNVsm
cmtEjPBahqMe2JSqxqA6xikMlFPkRi8ZDC1VXT0AJs4JH1BdMxp/9p1NXqntltV5bVefCfAbtKM4
JicIVA1o3S9lzXIB55wrT77GyGyV6isSOtpQi/7O2dFSsQsM9aBEsQmhRegSGHUCJzpIjXdIIjJr
ZfxGTZuGjAK0Km42W3wZZc1M64EELB+Xafj97Azq/O13aaEN2NIYA2FG2Xy2h5imszUC2cUHpQwb
P0GUnhodLy4wjNefOaXBRvx56oPDra8rP8hTpvXwmQiKXSPpPPyb5JdAZN+O4G1uPGCHqYzmF+2t
NpVFNC9zHwnqPsLwvdUitciKQYaEQioiCKaaIl+xYyoBw5AzL2YAAYeW06l8cXxMVTMnRaVlfCdI
cJ5EnJ+8GufB9VKQVLB5re3FPzRGqIWTfQBFHEJs19lRLGdVeuh08vLtLRqnCSrkCITAdysYzrOV
Z2sFOw/OA9Kqzb0Fpoo0qYbEYvguRjJkNkvq8m+5xf92RB1+LEIOPwljCDw3VeSWt177qR5ViErc
DKr/w3v3h1CB7LNlXxA/rHnnRhPvdFHb/zq/UwVMpT/xlIUVcEsL2zzUXsEApIq3Z2um/x2aNy4a
fXw0UIl40BNF2lATuRVOzQJatX1EUvQHi/uJzXCzwHI3W0eM9Y685iD4iE4bcF/Vnt12gktXtt0c
t3k68ozu75bbymfN6H4ZTwysCFEyt/n9eH83BfYsann6OUvZlLpvPKskle1tyh8Uh52o7uBC7ma4
+dIIGiwJjUTAGrismwI1k1z91XoYMXXUoGsi2bgsbsQKuDBfNlCbKhteYwTFsdBQeqxaAwg22dBH
ve6MzEnn9kqK2C9ADgGiao2MneXcVrmn9VrTykZBNDcNuHFG0+tkN2O7VQ2s4rgeTrWAi35CrOSj
LQEWtsGKQNQEHdQNrV5uLf7eGlhEL4V7K2rosJGJl6AghSky0jPqn64clabbwbVEEimDXh+lA8sz
AXOsNZFbUGw8fJaNV+b1eVesNx2qKJqB78m2rCCFZx7te7I39QybKJcShRYtoIVE0TMtk8CKI9xC
HnHTtoodncB/Q3SD1U0Y5wUcl+iz/BhRagDRDTB/59wQ3FLIReD8jodwaNYrVTCEM0hBx/c2BNK0
eu2bynPOzDYcBDFi0XJcdJzReVAFRdPaYYfTRBmLIfiukPMSjoeE/OeplHKa6NJhLlouheEYY7SF
Fay/TVnh/3nvqxT/6WfiZymR7RFdRhtRcd9H+vBQLPdOI+ScALEWd9Y5LHGy5IrBT+buFzz2/v9i
aX0g6s3b3Bj+myr1KSNvHci5X0Ds6VDJiIAwSESJmMExbVRXvXxFmfNo32mSmG8isBXvBbbvallc
GLbznuzsZaeYFD3V9qKH93St2+Z+XGcYZSUwqZV0sw4exj45ifUlsHStyp0JoVNJRqZxLKocwUAi
Pc/XZ5XpYwrsDcgOiEDFI2q0kh+W7gY01bYLxFc7KkFBxmZCuWJNBBOI4U5Xljk6RotGypdxy20O
mQIunT9mtxdF6Eo55QJWaHprWooNOq8CHaI0MZkEUT4Om1f7zKZFLjhrYG2nhF8avQbWwfwlBPzh
5IUGQPzQaOwka/8KO5x8C7zPg5Ai0x1dc0STSkIciH/xxyc5qJmYkv8Yf2SqQjvv++rdNpKZmRl5
e2+CEOc9RVv0oIguEVlQW9q0T1Y3N9tOyrYsKBhZLgDrIHklX8IQe6LthbFq4oNrZYJh1GLMr+H2
Jkgj/EKMeLYM60p/6e6egHzJScMOmaFTXgw3GP6uVGoECp7zxAbao6YyYJeP/OI6fiwx7bd46VUG
FP6cMgR48wXAEIgVWpvXpd6nlrv/ZoGP5YUEg6jC/DtoUg7EAbvv8rDKnxgDObR3Jcv0HrJsRm1o
S40VpeRCfTBbtt59Q9OIyRCzJXS+EkFwkx9MFpTksga7avuQ3NkblmE0n5Uj6Zp4+iJ7k+ZW/XVN
Wh9A5MFMoUTVIHtqsef/lr1F6Bsjtd2RlApsCGaoWnRUZCus2AOULFMs8v5mFvI7u/rzcrI24+qj
ozs9HuMqoHzd0TwM29fdsTrMhYkpNCR1MHyuo7/QlCSeCE3yVPUlxPQtWmS5DXAbOPAHrEykft3u
5feNoOKJ3HjQZOJSXJ4bm5o8qX6aQqNJ9nk0dhYpXyrMCHXBrYpjtvPW/IBhCHVxO2ZUyfItiI12
dfnMzqNfZyXvX0CLyqqNYNWHSXwN6yarE1+AUznD9GQa0dO2LYrq8VISFseWLKV1VbDDYgpj7yH+
H4WjvmMhBEAgjkoZ5v9wMjfGITfJXawi3KBxCxVF+Rp24dbIrwh/rOw//u2R8TJic3cPMvE/ss5B
5u0G/StLQu/mzvHAE/tRCcyoOlpgOLZbnDLGnI9+zhdVyUM0HUOlyo1KuHxwy/uDOZY4El8kGH/w
hJwePU0ir7IJVuhh9Ttz7qO2H1Nw7qAHR9NmJFeuKzMbFmegGY5PJbXPCY3Z/3nNg+TaF02UEgDF
hFghH/Uog2ClMjkLQf0QOFt8af39bpfjvphJhqZYwSlanfYdqvYfWl0zX0XtjHUfCo9/erqxeO0o
MM6CcB/MiICpPn0fLAOcxQEK0/0q1IzTYVw6UCmyzusvEk8YgPJ3p21qf2ZfGRC22zlZbFxj6ttq
ahMTDQvGBbXdUBX9uWLnAdAOYp270UgS9blUam0GWyrme8YKCuFLDIblJEwjuZjscXtHFBF3kIgX
dyzA6mjSL/cE5edXZ8ri9TSU7OhZRa/af1TsCrMbuWQbuHT8WXGv61pRVrqj8gtTNAQ0eOC6CMwq
REM6ofaYtfes4nn6+f3v3bkJKJl+VCHK4a0+ChDZvEAbi8ghsJV8VEglYe7pZ/3EATXa9S/hUPf1
Rx+KY9kbCCMPnpt5sS1sibHxm1K9u3Jmfz9f/qUralG3Uv+cXnw36oGVNNFHJGTgYlKMDf7zZKBe
NsH4idC3tfYpfDHSEev2lX9LqdJvyLuKNtG9Vsq8Un3C36UFtix5XzjMg0/SjX5QHPFZ4xCKglCc
Jb8eAnl/Bh2vwckSCx0vQYu13l5yr3javasaYD/RpbeDjCM1I2CsuLXlTHG0VKME2Oje6Kp1vs2L
xtre7TDgqhnqObDBgIzAkY/OPpEgWWZRYtnvPdwnYsLWB/nZlL3cNfR7TGXQ24yT05J13N5puFGw
+5NKeNUex3mYrFNlm7Cp8MrXk0SGYOtK69HlTZwB4Tlk0n6HXTB3n7N1CyX0kfSrrVNpY+khfJWF
KAo67dYjmuju8ax/ulFs7mZscjgFD9PWWgulQJjXgJACjU47iHYUZ56vVVJZkSN0Rp8ZUVMrXGtS
AHVbXOjvPh0nZ4PXZopqEY4Y8U/5jeIoKTxWHHDZO4BicDKnUQ/tmbedQ4fa5ATBpj5FaYm5oXmp
Fci5I0nV6Gu9uOdMnhNpOM5l1QBt3/WS2V3y/COaL5PJ6VJw3ztaj7HXTPUjYTCZBp1SaL0cQxZa
QjnXGdTStCOz7hYKqtX9aKemMaNHTr4WebG0ND1H6BjIysH+R+z7l9mPd6IZiNjHS2OeptPU2Dha
sYyVN+p837sN4o3ratof0M36dLMSaveOB/m1h0Y7g+vd8GHgzO0A23xCWDQH1qxqxUqQH+cNfAfW
61y2EvqlOkybbF0+x1nXaz59AV5nNCcljDqD+3Llx1ghZUeMjHtZL+dXS/zrxL7xxiQ+r/DYxA0C
JeeNMyprWXm5QZe9Z/shSFFFfH0pgB+aG39+jvt+9qhMkp5JtWl2bWsSruZw+7YmtluwMk9kVKBs
b0Y0Avk5iGY9Y1Dh3tr/gmtxuJZN2LTPZfgcA08MZ7gigrWLlTwdegvic3c2Lc5OuU8L2mLLCAkF
BQ2KCAGRIJIntipAvVaafDS58Rf3XrhRVVgVaNlFiNAmjOVFYcYJ+7Wz19X/NBQtHVwL/5k53xi1
6YNl1L1J2oqWij67ygZVa6RilmhGL9/Tw205oRGmm7enBjESfYyEljv+uFOvSXEIYT7m6t2Bd9RY
JAcjH+CtSyBhddKN5D007hkaHcN2BdOHTLWxUn93F6kEg2Uu3dYuWuE4gcJ0lNwUii1rE0bsF1cA
Xcic0t88RjWuypzHe8hZsnZFbU22DlqznwYNpT4MIIfQ/6PUpJ4vLkqv6+Zw6qa/FIvwSQQWwt+l
boOcO088H/E1eHQR9AC1hpvFu0UUkRCq8Qbg6S9w27ph6Qjc0n/tffAJJ882c2lWigFAfsqvyRbd
sKcmOsCmpu/QaL3+5jILdlC+3DcTAmdUnA42n2VgbN1Ffy5xxwXK5CrkgZchVXI6Fi8hIkPSsJP+
RCoMuC96Av+RllRmrJvPrt7kNFeywE2wcvUOs+dpJCPki/hq7YWUpD1hK3NCz4RfdPBH8ZwpnTSj
lCrhaaMdv39E2zEblPkLr5k92frj4VWZo7SudL0t1WMIoD6hmCOLdHzHrQZqtWwbuH7PFt6GnegH
XLc14oJxPdu0v23elo1g1XDcLf5js0pug+9OzkaG7NmeRtJWX7Swl+qv6KODEyqh5H0LdbwNc3X1
oGkrbTvMfVtmofgEr6VJOA4MTry+nWYT6jeGioY0KitxH0OfxNGEVbH/hK6XHu4vmfWSJZq9u5Kw
cNaBsgpj20AqpxJlOvkW3Ux4moSG5zzWetEa6kASEl4AukcAmT3vkWu6W16SwSW5P/lHTp8yL0uN
vnEwXSUOg3/x3g8PcFvnpc04rwYNeh6wtnXJdEPGOuZfe0KNh59ZNauOdxN/k6WLi9uVshsoLr6j
2J1a52Ip1msZ1HsxcQxYqElvVEepJyQPDZ5gnTTkBjnAbDeD7UIrabu/71AdxmZIQ875vC29B5yJ
gFLU0y6gQ8sx0lAks5LCG1458R1iud0AvNPXko8+UFrqkNQ8dVwOK6a0TAN+Nht2ihRY80NsSsV/
zIe81PXhORmRlHVH4mYdJ2NGzYdTWQMvoCHjv7T7wQegJuMa8Qe93suk1JOSJCDaAPdiHcGuaapK
b+B8npyDZQWq84QrfboxbzI5f8hNaCyrC9Xbc2aAouIdNm6Dst67u/lRMOpc+W16TiDDvs+EEAXm
J4/YC8e6sjU2gbvX5RM9qkV7aLneq10k4IOc8bsth0ji3m5u/S5Ymrtvkxc+wQc3w9wX3/0BL510
Ww/VJg5WckRTxmPilhGyZVAVfsg1ZZQBj1nBY6wbTd3ny/tyXR9KLfLQuLoYUcCoBTpaXL7uIhq+
FaWbEeBfK323P15xzvTxEo/P48kODoGyj8eZGfQtK2ewBp4pYTh8D7VQ2A4NyZZv6TrBytICibfd
HNeOMk4dJPfuoPvaVFstOKoICy1rowjRymNj8ldJFCGS2Q83afnXkppuWwrO8+p08UaR9UkGGSuC
pt2MVMfVTJDb8CSr/SULfuib0fEkV4KtkGdQvIoWMS9JtGCdsWoF48xNGfHyg2+jgweDJUtVRBvG
4CFpYv98KgIyZmnZiLN/pUtwwyHvPVDDBdAdDXTHWa8YdIb2x0ocUIcyZebHnjFKazl6SyxW5avv
wauDELsxs2OZX6Um3T8mLcdtILvnyaeagTea92hxG4fOjuz2PGpUqVp177aJALhOSUF3pv77bKZQ
2jHe92jFjURxssOJ3yCSjFemD4Oisb1t83Z2cZWf1NJ0vNCcu/yUq3TcRs0WpU+FlLyuqfQCThm9
JqaWCC1+pPPWLrjuKu0MpYGsnxEtxva1uiTo6cPP6m4AU+qRZ3luqFoHJHxaKZj+Z5n/dlOIxwOC
oqYzuM9gpjnvHthGjmjbXP1/XXWmbDou79kggVpsTERFpKM/Mba3fZzAh7gH4DaOS3+D//QluZAv
M7DjQXLA6njkS/4Cjg7/vSo9PconDkRcBTI7et1aPk5oNnIwVqQYs12Ty8WAQainZOCMtSeO0TGD
lmYn4hDtLiCSwY7SUcrbGopqX3fwEQ+e0w+A3+rBKRnJ9J86YLdLfNFk7pplTuSIjDmGDJ0z7gN3
TcJ5znNdePAv/DvDJNZpMrib1NkvE5wE6Z575qe1Dnbei+uGw+FWbGM7h2/x711r34LcYcR0hNCD
wMZziLYxsjbHsPxwULYiD1f/3HhYQrDEdnFXjXFxGl3xB0uD3S+3fAHNweY3os+v7XMH8xqt0pBE
pxJRXcsub6sl6a6yE7geBFKxCGWrF52lDMLwtyBbxx2/s3qg8CT6JO10yS0dU22bMjEeIcNLvUKT
9MjbHv/lO5/4l0FGfZKOOno1cb2ZUk3LpQmBGlBXt35zyPNnggydYDgwIqI22wcx0P0DQPlxWz1R
olma/NAohh1Wfl4rdgnuA4mAytXixETU/f0y2LEbM7OMfdov7dqMt82KzRCd4on5fYlAGs6bqndz
z/d2eGE/wIhIPN/eevwLce+NnSUEB6HWuEiIHQd4kdqK3yx+Q1LJPhAaIm2v4ygIUFYonlzi2GZm
a9xp+nmCkq44Huu8PyQROQwG0piEKH89NqGPozGzGnCDcJ9c8qsUrvnGa69vnAipc0MaVlSONiUs
xyC9lZjbPMFdAF+ZpFLMaVE+h1whiXwF4mGGqaGuvYhaBqoDMj14XGJEF4Qwku4nJJbVCmHYB7dV
XV3nUP/xQhqxi2d4nqXgiCL21oVEC++jsxZL73Tfcqoxh6P8QRnhqvMR61CWVOS0ZkUvUUHYHnQh
N/7eIF0bz0cpVOy2CoxAHBf987RmfBLHp89V11e7oJcgnJWwuBngPzN3vXTDMUw3+3TR2Bskf7lJ
OvhMJh/T48zWzAbzYtvXk/am3a6luEsb5Qyj7SUMylM0wEP3c26dIjYPb3b0SjwNuxQ0UzNZWabq
jyDuzRx76yTf33bQ6zrXLMipnZLEbw2heN4HUVswEWdcz0w+6hFDth/HLZI2pMEV9yyBe7PeXbUN
GF8uaNCh4M0KsXMYWAjXdQy+Qee2RoOSCMntyvRqjXqk6vafamdg0lbv4qi+827h06VdHu3vRgZd
1ZKxH/3KWTkW5OI24d3Xic9tPJUb37XFnxre15Gn+GqrPzCXCxA+rTTmWJZDBll83mKZy3FBmAfx
gixHQuNRnGPf/78YxfJ1p7MRqByU17oYMe0as+mUrk2QNfPT9OzsjwQ4syX7FkUw/vmpaSxw6VBS
LZdzvIEE0meXF+bPM/dxEb/Qqsk9G0N0icCeh1i4Aw82/h/KvH+OQJa1hTJgiHGg9zAUo7TgiDP0
PFWT9tjE50yYJvWSvA2jZDtzpRkW9ussprzLooI1nWi9fWjPVqCWNI49cZJvUyiU9dCumwgl1HnJ
+AVa1SZIwP/cGZivGleIYGF5Dc8pBS2d7Vof6HHRwcMMmtqn5SkVkTu0+st1KyuailMI9q70VKDU
VkB/fIoCItueyKBGOqlLhFrS3zRqE6idbl1kXzX7vt55n62qZqFPXR8Dq4FbTeWZJEQ2JFsw1H1c
murPZ2lnSoGFl2sMpJ73wOmV39DG9a0dCOshsNH633mFs7eSL9vABJ5X/1PrvnDYqf2uIvFDJsJH
8dHNG6jmV/w50NMeZyKltkOEazJuP8A1eGSyEHoE/NhjJQOA6Z8sBQl9dHpS7TI+d7LiwfQJnKwq
4qgCRGO/9Nt4MJGahazjKDLQLi36UBdOjd4TncWkZMYJS0z8vDizfnnRbN4b8UD7YWviA/J2+fT/
wPx2opGHY2VRRX6FJcNYFJ/HPwkLnr9z/Te9tvR5p86QRWI5Qu9SAamZMcuivYfvp92In5KO3r28
6PnVcKOhnzyTkhZAPrjbVAE8FZCnh2UkFZ2RP3TqiFP/9jcIH6lVOe6WcIEb+2+pdk8PS/KuYaW6
Z2rJECX+iE64bJGTVxEriwuCHOjW+sqkFwPlMN82plM19a7Acyg/BFdtcVxf639J/cCn9MHPV49j
bw4UoyRU4Rk93ZZVbI+T5CAd+mkvQWZLHanPZNKeuNTj9ZAvioK4nk2xEgq/4HjHrDNhXiHhcuIC
SP1eDN8Wzsknhcqe442+CH4ovMjYWqFZtpz3Z+iuMrDZCcl61zEXRJTx413NbrsCJG9CjHpqy1WE
Oe6KAJU4u/f7SaH/+y7ayJS9rTZCtkCfphsdfO0t8P5VTQXIb+VB6rXY0vo4AO5OFQKbSXa19cqm
9c5tDxuSXpFjNt9yyZK/wxfrqvcUQwoko+4g2W+zx4k3HVfRkeukwNmfRTkK05eUToPHZ1OLUv15
Ac7Xtw1Vojz2R8IIP4SJGs15k1i3zUJJix2RwFEBEvuyJeSbKW5fQCLE9yfTg7HCkPCXhD0O2bs5
vLZ2OVcLG4HFsREinge77Mn+dWqAT5sDkIog/Dte2whBtY1Ai3kqAAH/aWlwpX+EueGQB+X8Ofki
XIaTsZJkqBo1uSuhrRxXQKOFtPRY0T39+vprVe4OWTy8TnplgTnBdOlPjwL/ajTLgDN1XZtsZhRt
+y4JEOFreTbmXq49v1DksXZ3vDOV4E1jVZXs6HZZIS+Aj4i8mpR+6S6VglU7kJXUmHIu4itgL0W7
5+hA8JO+Sb5B3NpxKjQrGjW+1YGWW1N/iwSt3h6KX2Q5mObnFZ+n6tp7RIr6VqeJYBwfb7SCSKRK
qKgekNh/+YbjmJA6n69izFS38cU/ZIVVrcE0YD9ylMhAz8B07C7kpCBWXED2hjXdpxkulh5t8feY
sfTEjutv3xLCmBYCXORcktD1JsXxCnmdrdAUz90Vhj0A8RetPSTkbR/gXnj3pSO+byFEjbJ/kz91
UCZra6M8fj35FBgBOkG3GichcJxxFZDUZZFatSpx/fZTf67Fl2vi0uphtGxJYSnPYSZXcDzbI5iC
dA/HVyBtTN8QJPVnJRtWNtptZaiLZUnKYOm8CyaoJqVLxyOZj8j2fmUkv+Jg1q/MYVTP9zqB853e
RJ/32Nx9L4rm1ejCbjB7StEAwX+SPkIQR9SOTLcD3OiwVMk4sUmu+WvZM+3UQShB6OcLJ34fM33G
KSRdu9FtAXgOib6c2JBOvdp6cHiXSVX8tKDkiaZZAodydlTZniziESR3RMbTxOd+96MM0veRImKV
EnSfBzvw7adijDNLYEveYzYzJ+21O19Z2YtXve1/hndTwPNcMbFpbgvW/7HNyNNuWrjNoUUtI8z9
ix0+tpYbd3s1ZJ0tnMjwjn/uEfdIe4C3P9EmvaGz4xSFep5ditpOo3e9lbDbUtp1jpPrPKNEYWv8
M76TAusGGof5VY794PBNSzkXqVWQUxD8v3MNA6p0o6k2iQRFcjUVBPN4zLxAFPhVTeiZFFJnpWbB
IJmRJKRkrtDWHLVOhSCiCgdIzsA06Qd7t4Eb9oekW72xqI5OD0LIv8S/ovCRLwzRkUdEAbvO3s7A
9yBAgBDItCX10aLPSFa3/8tm8G4BUvCPjr089DKSUW0wXzsLrNiNiW/8TTJtvRMxSpQUrTh6cwUQ
OBG3stkpHMVDK8wrP3Z0W0uscJjZfnEUb487vroNZRvzVrUI39RqxRqEYOcb+BUzGNtQQgn7KdU3
slXySJbOvI/CmAOYfdnhLFY8Y4FFwU3f5WBhkwHnhiL9M+Q0ckbBnR+i9ZZJhLy2CiEJ+LSfmF2S
Qu7W6ka1U+b7qzUv99LOt62icKhDcuu75i7PDQoTMMa10hnQjjGl9xuBtsedJ1KboU5QRu1ulCLG
KCVATWNbM0w6wK3+AQh2mhSmolBx78MO26Hxy30Amsz2aTNpnuCcOuvQEwWECMlZyfY08mP86jhf
MwtWtrSFBrmiEZeRLDAEWvp4U6Utgwtlc57lptnMN4dovlFIyMjaeSkAqWWngITGRTB0hDCgOwxg
grPziomMxtOkiDOkEKzcS+ZyVt1ql9FbGQSsVC9pf61Zv/rEQgk2hu1fpijPXeHFik/3V5CyztX+
+S/Z2Y0cQIaHsDix6Fltkd9aLPk3ktFOHR08DpOe+C7UAvT6sYAIv2F0PVBCqjPYxcQPAwH9gU3z
Zo11yrwDh9cWWzCpWYAto3abHJd+6Q1H5vTRNzF6jn7abRi0meSrZi9VT40mxuzU1vX+JB1UDAu/
wDTvelF4NDh+wSYCxk20XiOMxlZFBKJ7MiiewbyxbG/62xuRJcRKmzkmjG5DWWQA2PWsu6S8sa5D
2tgNB7sFHaFFBZSnDgHqQWL4t1BR+HCSgLYJ6iZ/c+RrJTMJ7cxVzCVts2WpquqQtplyQK9uCZvS
DzMYqTvLLcZcL2t2Tr58WTEaoJYrhW7e+IxmvEhViqBpOIMEktyt0X1AKBHdGYLtRoJBM51EtYgx
wNKjljC2Mdn4w/WLUzzeR2iI9JO1ITFXeXQt2helzEASIPgBrnC3Nxt21itN8Y473zqWBWzJZhxs
4/u3bv2jrHlHiXIrh5MkJcv/YbZWi2Jc3j/DnPfldVdguf3YodpkVs0NTeDjwZ4VOwgh5NpuVa6N
L9Yz4kVdOWtEXUw9xW9BT66EC3aJlGbHFf5uLzAomC1JgM9vbxIN7e/DFjswvmAtmJQSy06woKX4
VSJmTFobPOjWjDT5tSI8R5ssIc4G6aP1kl0ZiYbDtPCKm1Qa1x5k3J0nuvyFHrJ4liq6TbvZLCjm
iIeD7lEUtBXkO8ufljHQWUdyH4SdqNMrgAHtS/P/qXW4L+6ysgeqMsGeLf2VdSsWv+0ExYwGXQ6b
YZq6IrqVGihuk2sNlw8QyvBMb7VRgXGIC/1qqswFPI017RatrHHjiLGc+livRB0c591GXvgEi9pV
wqsMtQjDJqPysJBmQcj6N2I/N/kqQJbmNDdL2AFjqYKk+eu1k5NKSW3/ETMntQqpp8Cdl3QhUyNv
7Zj0fvac5GxgiunAsWqCHBcxLSQjhehCUTk1wdyFcPgg5ySVkmWplj9axz4dYvDwJUlbSHtMtmCZ
tyO83y8vtIeGHqkcmcrcE1vKvaPiM2yUMdggn8ys+OJjeYYUOVBrIWvKRI47CMtNQRL+nPb7Ot3E
y7XfLJ6pz9z+4wSGBGjogRPSVWs4AVe4Be4Pgx6mLa2kOPrt9XfSrbMHd+Gv6XxngRC1/IyR2IFY
9Jnv5Q6yEAy35dnXCHOH7EV9wmxyXhx9qCMkRqXXyu28H89mYwaP/IWNTQ2eQBoLJ+qwhretFe3u
7zsSSn3Q+Vm/PPKndOyk2/j2S+IlZDPGdj+cQvUj6fdLGQGAe/I0MUkLNGoCJ3coPDAqai0XbFHC
z4/7CKkxFYm3du8/FPBOFeKinLLV2fziWffnyZEDd+g1KQHI5GqUFwg9NjKgqDaWnC0b3eoqR56L
LoPKCVtkWT+bhdhK9wTJsIdu3QaRcsseqCsCNDdIkZOXhAZ4sbk8LTQVgQST24Ehnle8/obZyrou
Z8xWzdux98L8jGRyTpTLDmBNKV6UMrRI2BJ1fsc19uDCJh5BRc4An+AHAYDITfWUozhBHOKZQTUy
9Mo/CyZ4KmkQ2uipgrnjGSke6caaOFqfaLqYll0v9EQ6p1JzrNC9qemxwTaY5cV35UAck8wIyEmg
n/n2MQULIMB1efiXGIFFUJTLyiTUJrIsFgn0LMBVXPX34upm531WjYzBg7vzGB0YMQjE3AaGKHb/
47mrsSeH9vyVkqJQG6KEiBoeuLdxWnZCXG7m3gH4nbsxCsgh63JCV8lBklAX5U9EY7Rkg2KOauae
+4krA0uZwsT385KrTCz15ygdcXoxyA+lVj0nq0xUQgHS4F4993dEx2X8fEUD17mjz1JSGhijGBtC
q/NzOawFGuPxVDBx88RKv3u3r5zwCxDaX3HLqD5bCO6se/evvtwfR8Zz2NDZpR+Lh8++Q8CikDhX
05HMlJ98kXnjHW/2sEwiqIIsvyZMRvqt/IWp5XgAgAv1Wi5btaZKpO87eHLCZsIjFKEcAre/QWHw
H1gfwZcgXChFPOkyumIoS2f4+fa6bZHpu/yn1zcedvLtYdO+Mu4MF44RXjIePnncPng86PHJCu4P
LDe58FVDlTpTMxF3n0zmsmlE5z+nvBApdY+3O3brsVIqJbzbzgUx2iEXM7DZ8JZrEOZ/SO3zu487
Ezt79a/3u4y3ygty/+oshDcHhPbGX3bWaYUPC/VGEL3vw1Iw0Hqec4XxmtsHyoxjVZuuI5DJa/eG
DmSeK8VQYWvIKagBGXtvJ5sxv4fy0aWNsvwZnA/YcGOhrMSDW7p7ijw80cxk6KfdOMdSI9IsaLvP
lWuuYjfDqcMj7sursas8FT663uoDkQgZYUM9HZz4RYf1pQZLv0ZxuVSD/Cv/j10dFO1/ZJsAoKnf
GtYB3PxXCsNNpAtLnjtgVY5zI050LMuCHpRrNG9b9aMCp4KxmrdSmn77iR9qyulq/2d0DUQoloDp
ZS/LB+ACRUKr57k0D5iUZdnKd1BZ88aw2s4pr3SnU2EkdGtlUk4cuoOoLjzWxREsW7O0ft9yX0Nx
Qsthx8hMd6z65Zyk/w86InDtMpaBW3Z4DgnnOSPTSLIW3Cf6ujEOA6nWDUO/uD2uUJ0zBroXVUFO
nkUBQFiDY36LWA0ze1NEN0mGEZxgqB/n+yh/t5DRNiRVsHVSY8wt6lDrjWPkT5ItSI0L7C83ZHJh
rcLnzCt88HdXfG5qTSIDBUm0+stcuQcPaxwWwR1cGPletyNhCk2IahNalhpPyKRzKegMewGF4Iqr
iLfG4f3lk9Kx9agR4k0t7LxEIiQGSj21Zy2wLuS+femUM5Ec0bheZzZhpnSSWFTRrZ0Morzntcqq
bIWet3SI9LZlxoFfaZPXhGW3CC4okXSVeB1lzQ3BdaIE6y3vGdEAodqD/KLZQiIHJLYrEf6ISNpb
JX4zVxL7YmvDSMeRQhzzDumIeermWl0iS/7iUpKK+jzSR1ZbfBKkjBstzx92le63YA4NeK9Omo+d
BK21bQJ8s28IA76iQ838eGBRhazOedrquZvAQcBXcltfk09kVCy6iwxlY9xsVXPVn/nqv6XG77av
FW7ZFNNrJtJpAWIbX9FoGNDSYKsGL4T1PS6I69QSzpyEvbLa/HO2mjNgmU2Z+DUy5k+j+IaiwdrV
Pj/ZmxjlhwJLdGtVx8f3t7PaBuco6vS62e9H7Jj4DtMAnKPyiFI+22joEe3whZ7F3OezLVs+aXfq
QHtmmOKVcdTUefADZWjURizKe4MLCRrWTBdt7ESXRPna9mrk9oxiH/+ERIpgLdSaMHnzSGXMLUSE
bBbTQOJ8oVCsf0YquUT8JhPvpQLFk6vQ8wHZHX5srYKmhLHdsMOHfnCa9knVi7QrdDOpF5nRK61L
QBZ5ayGySX3RZ8TpUr5ylxdP6NyrzU4kq+QdNdmwO32krL80GZEgWybWesy4m9qReeK+z2txZ3+w
QKihHVZcOkstJgMD/10tV2FHQph2IT+6UlnsjrwffMK1Lw4BfN5jSwGhjmEd7d3frANLvBwSTUXe
nmROQ1g/cs5fn50zFJrxgXoQkXI/VOIK7A5vS2mj4/8cktl9Z8P52xDKukE20/tc2AOZdYSMn9oD
tQ7QQKfxLQLFfofuhTPLI1bIjUc6Gb1AzHW0NpEXzwEWgJvyZ09YvGa5myGUf9Si6evc62yEuw7f
YES3OkENj+wMva8Zk8cpRCRf3DboZgQj7pwLIP7tOYdpsd/DNcs8hMYVr9a15Ovf4u6crNZoV8hR
24B+FD3pnkNzuRdAZ8eL6rdmQKUB2FWJAnbS/IogD2GsKJHbWAjNs+JvpPkHHX4tiH5s2Rcig/r0
tM64lWICTW30Skcf5QOrK2NyrDLMcT8Vk4pKblXv+b+vAxbw8BseaABh4lqtvGAJihRChyHPbIas
lzcvgQuLmdrgMcTTux8mw9DwkAdY1tBSp1IhGs/dI3p9YqEcl3c0BImEFc9N7fUoxlXRbTlI594E
XOtyDvacJcKtSvN9NOIhh4wAlRjPKRqG/q3OHoPwBEV4mJh7NVVsfuv1GI5yuS4MzkaaYCvOnMzZ
0A+mHla68/42NLoCS1NImrxgmEIrclj/LHs/CrI0HloqX/tbJ7OMpvijTHtJP/Mmq72wSqZzfYsh
x0blc+2jzDoOkdR4OBi4jcEmaYpzd8LQKGXWXXzZYj/Urrku3DwBAldMwrxXhBA8Gknouont2B70
XDMF4t7ZmuaPSMyeToET76Yk/P0Mg6zDkqjhkiNnbPNzodO7LMMaJ8eXb8PH1jsolYXQgeSqXXCa
E+5lyWzGjwk399Sm7QGXmFCcsPRWY2fZ1RuuJnLD4ZIypgBJbFi0NXbInvm+pi2N9MgtU2VAFzjt
vjAAri1BKOxifjgXgvRVJK+EbJpRjidrPPlJccJSt54PwYb7wNI4H/GoNN54BxJMBg2kXeVspZzN
JBl2rvKO178n+gXSnOL+5z4o2vrnagiN05q8FsoWPKQJwDVa2FFK2P4kA7qeuU48kjzYVGZFnd1h
GU0FI4TjHuhxPeHbPNUAZU+zhpcPwEvc6rSIHXhXBIEPSdrAkq+2e3mftjp+qqFWSx7knmallB4b
B53I3Lgsn5qo4R4Ld3Cb4IHE9cq98gyoAwAMuGgtVZrL0FC6x0vn7mTrirvKhA0jMcx+IAo0tzUy
6kBpp+XcBEKWGtf7F25Z41TW9/Rmt/2Hp+Z3C4SHrn0apIZTUiFPJKxWFrn6n5t+PypG8a/n7hhN
867csCQIVz5y8AtaGxczS4rVXV4Ittc0hJFYoKpVDGuz1uI0FAeA/iX5KNIleZnKhhtmeXM69SsU
CAtodRj1//fQarpO7lIrAFIGtTCO4Xpnh93b981zn9ZhMe95auoAq8UW/sPrBG3ZHuUbUGePR/hO
ZjQYYsmFztXsRi0dgizQa8ZsDgAvwN5b3dgNggq5Gq55lM3+jApgfO/PFMt6jPoFX7VQTz6n4tOn
FSg3i/CXkOcrLaS9hwa/kKsI07MBeedht6ZFchJlu/kt51zLI1cCngHcG9h0X5X3ffWrFbSijpzm
psdjPJuxBN8pLAjtk5wLuM5Vp+SjkgcK0mtioHD5TarTDTE43Yvk/qzSK3ZQ+6QzXulDXffxwtln
BCFTOVuWSm3L8A+N6BYuSwLP9vHk7m6RsNXNrhUlsiVYT50obyKXIXk8gcJ6C7cc0upBaEC5hKUN
kdhmuJZge+73LLKtGYvo1FbWh9cK7uO5+4xze63Z74PFilwZqa/IwnBG8j1WER4MfhnY7S92q+by
8WbkRB+hR2W2bpDIZax1IBeRkwiKzl2y1Z7hOgyfulQVUR01eEzraHIlpTpD/llK7cKuuRWw+Vcn
4mQkaGUXarGuW1mbtK+laTxATR1yrjRctAVxTexsDJIA3kp+YloY48s3arrGP5zBNry7DV5ITvHs
60zqklJcKiSQOGyBa9HjbBtMvOTrkGx1GkaIKVj7KFpnKKs6CdhSzMd6Q7hjdXWDGp2wEokY4bIJ
zl4furWbv/e2txV8414Wr9A5/uClJUDTf4+RRT9q7VePnlLxardiVzvNkok3VPOz7O3Vi8OpeqAb
fI8LX6K3aMiadl3wWRVN4em64/klQWsvzUFZvdq9MU898KGhBHinRdQeP4xgKQ1rnt/SDpLLmp4o
1HRDkWocyZf5e8YNwvhok319nIP9hnbe7Auf3IcGiIwcGUVZgNAmttg2mjYJC1eR8bGksolqkMF9
sKMCIIT1xnWQZuldJok+mvy7+QT7frQKecpu7SmPK0mueoeS59IGXSyAz0y6e9AW+tkeZ6jdUwDN
N7+/m2lMC16s07ZViP0leA4AXRkBiNs+tWTGgXeVQc8Y+3AH1X5qx4hFbMvh21BZMi10sFPTgZkh
lHZU8PC1uqJq+apC4bBLEw8+hoEzPXyS76ms0MLwx9kmmntrQX5TiLGtJhbM1KbAbHSWBDu28xc0
Bpf5nA+ejz+HBSstcyB+6JCh787IknAnz+J59j2TOfQJfLTp9EKElxagc76xOUlgpiDjMtJZc1s4
gLEXJIeGOpiVs/7KoCkN5rKWGu7+zitukOXy5nEFmR5Kpq2EbiOetbCvziCQGcSkphTfJyvninft
lBcayz9bHhAuo0YRXHBAub6YzHIOf0VsuHvSzTjDqS1T0HGstUtF54U2LkQ2NqzXCRH9WWbgMa84
3dxAqpElr1optTC9nAeBFdMEDxNSdA71jIGUk+c+m8RT/BzC7SKmPNNssv1JLrHe8ToTGrGSxaGv
k6Y432dZ8AcS/ktk+QG/HZTBwygV1Fxge+ZP5hQL18YfDpodSerQebgXeigpfra0r5cgNsYoDQsD
++uYQhM8POV0gQ9fyTDh4RQac3l2QEyCeRd0b+rMnxJTy2i+o0GDAm/tHtBcmeh2UFc3R8cnASfy
Vf5BED+IDJ6nfBHMz0hwZLuIFeerkOtMlZaN/kRKOifOxFA8m510pbJIUNA2Lmj0E9fHtk6Dc/DD
mtfS3r/vdKUPMFN5Sfbpm9AZVFe0imG0/4un03seSJwifh3avUXMRsYE2N/Yf647XHuTmlnZyl2x
f7huomBOg2phzu31gbspG/b3sM3UGy7BRYN/oGUwxZg6/M3s4QrQ+nqyfSttaKhjBSzGEt8fWn1h
F68zO73bSRHxBUxPuB46z3Yd7BcIym3GS0J9oROIfWwo2K3tiJkg4y3Uecs6kJD3rsw1DSQJxElS
mBJD7R7DohT0CGdcmyEzcvhrIHRQ1eZFhf6YMg7XhmB4xpF15CUZosMfJyTDd9RAAG8ksfA41xsY
i1T/8D3G66PM41rZoFTGgO/ObgJedHHlxHDF3/wxobFtGnEPe8FZ9YRHup6UzhCd0rNeXhAb+AS0
aSedrvLbnRg943gjoP8aWaOGEgGj8bM76HVjUY3r1myXSS0h+LJsiAJSl20xS5DXNS5CjTkEldqY
3uybN+AnMBIr27xXMH/H7nRSjygn0/bD6FemAH3YhI3iAFA1NrFWRsISkxdx5g2QMm4KdXGesV5T
7Z2gzN1SLpJRyyMOWgbnPtcolENf/byWavGYNSVURC6fBsJh3OzbrIdfGPXh96UYShU8yJYVg5mB
Y1CplpJrgzaEhE4nW4mdiJm9rMdITsXrlCVygnpm5khgFYMBVRPqK/sQgnx+S7qO4FZcGnIPnHhu
CQt0M1YOlGJHUWRmjuUUCgv4huLmuPNw9uPHO/SFAgEQbTaNlNXC8djMnTlFITRJ+SzT+k3ocXPX
eKDVU/YnaVrZGU/r4cCKsUZkYl2+oVAo7zHXSgkYPwEiQVfJaAM4u6G+LziwfkRrzUWMUIFACkvv
qo1GjnZVIs+ODR9KmVpWNPaIp6/9FhkRJCkeMI4wocMUGc785uh01tWS+rcnJiUIJdphPXWZkcOs
FvQyANAAMoToNLASc63g9Dw8Ms+8I0prm08NBrwaZAlhQzLkodm3ROeOp7pPPqnuZawKpoRSLPO8
XFCdVuTUN4Ym4G4elaha0vrLIUJWo8ecmiK1LHipkb0ZwOMt4kXsXqefEIVAHs2n8opZRgJjOT1J
6p2RU6J0OoY8QhG+Ob6E/fHwmWagGKgvNb/QUSV4r/H7pj2pU6Td1PYULpNax+0LIai9ML7LJcxm
zaRPXcRDYxaNQqHa45zcB/G5mXuNXQPvOMU7mLLlB0qZTLwZfVV34YZNLNfEwsGWeUfllFqE3R9E
HdiOhMGHu/WIRoLsE4qzX53UJ7I/ok4/qj4RwJR4dboxlBvddQkhFqZQcVE5nZYvYZMrsGNtFWZ9
K40m+FrGn3/LcECc5DpBxB0T9v0X5KXaqOjbQ30+gUWFS8BEVOXD6Ct5AR7r4MMg3sFWgNB82Rcu
uFm+zlZ4bLl7TXYhII52xyubylnWCiqzg3Gmy0IXC/D0M1IfbZovboCzvuC5jZdD1FztF27yCQnR
FEkzzJrMYY48H6pN0cDoAxz48CYhGmRsNNIeIdFP7rqszsCXcaKugWx6UGZAqErEf9wkmpIGfBVw
jE5LhZg6Y+r9hYvQq/Xd0n7cf0FsDms4GXJxuP4aDPzzb57IIAL6/mVzmoBgeLb8yZkLSkbO272B
yf1H5jngN32L6C/xp5n5d4irBV39QWZdR/B1LN5ZVEn/VmvfHKK/2WBCourCsYTu8c/9NwzCjkf6
eWoWBRUBGAE5m8ocnQzslpbmdY8eEamqYQglqpcZTB2RSxgdzTi3YMfVEqRnJit6FEmAqK4bWPeL
sCBCbJinnNxeblYX6rr6HXNtxvkxOx9/k3RE6QCEuXMkcU1KSLB6h9aFAh5THnigEuf1PCktfOCD
O0gQDQJ8KbpxFZkPX37Hkh62XzX+G6X4cYRKuk3x7LIt6Lh50O0QR8H5s71vNktXk6sSAwK/3GXl
2x1sqsXvB1VRZimd43v8mGcvhdLLIgjmBAuAzZq8eiyF/i9AOL3trwL4FdJKrFK3gEgt4ZekBOdG
2Ep30JTHPa6vRovRCv1HulQ7XDtKNfKr25ntCngZ624GNX3VwsVlbaPNAVhABbDT0P9095pvO8Qw
ryDWKbMkO3tGxpNWQ+vIeQtt57WmvYKJ6Dnr5nzL8JhpHBjUoQ/cQpuVo26ZJCtg7Cp3GF5uU1gG
u+nere5BZQN95G6j/eQE5qJKg8SeT5AeYlo1ThPuzod/dSg1uT44Tul4ef2Kdf3QD0N65gz4DMSN
IaXOkUFFr6/8oiVbV+DT1q8wMDMKBjmR2KnTqkTJ0UN3+C86csTlshdyTLw6ZxUniFsARkA+BfYL
77rD4v+F9N1/KHPIq7dqLL/JBe+co1Fw6VNYflc4QlxajTQXzp0/d2nieQos4GQ7hfbNEU/3RnD1
ta9wwYBYf4XmtJMVKgdJAz404YFIezF8xRJJKF6HoTTHVKEqv+NR4PlOjTJ1vgZdekFcUQ4RlItC
O3RCPypr4qyJ4vOCd6Lpz22zp9M3KK/+tvYDvJgjPybirQPdHpIM/m7bLI+VA8TjHQVBDVSrEB1Z
rUXfU1ZxA6ZAGDukpuacvNsDX7VVfJND62drsu36BOftlnkBiYPfuB+UDWXGuZPc3R/D8k1c8+9h
gmgbMuPJQTt3jgmWibDBUed98EkB0J2eIV1FoOCnwdKmRFfKObyEwW7mrPnil3rWIgfw4PKHyLoQ
4bAbddVH/IkosHqBdd2KG+1GvfXXQPsA1zj4dlDXj7/tSGPnLYl55i5AieW9EKZtZ61fHMgPUCba
BkSSdBFggJCdLpC02u+YhOAT7Wi+Few2y7UgiZddu+6/tbzOaHi1ZSmDFPvGlLyjgSz+P7aKjU//
hmPJTOACh5DGtZume8ptTrSEPYedXnCozgKGZfZdB4pDt/z0mgsM7XVywH5soSURPVraF5SupVDc
uW3m8BzpJcKWpGIIy/rGf+xBFJdc0G0mYmxFJenI8qRGfUG9H6jiR0uCKqmRaK8QBD+Vp6/am/VL
e8yZ6DDvxfo+ojryTeI+gmCxQJ/j6rVTPVPsc3iHcF3/R+KvWUqM0HxoSAnX+mSdWg0CzQpfqgr7
i/YiTybRop57WxIkmyh6HP8KDQJ0VwBBnN/sGv8jU8dH4HhjwlkKOYHTN/ib1Va1DdH2GRsgMWTP
QTXCzHNMV5j5mQ8Ta/C/q9YE969TQ5KP4egzTmCIP2cX07bnkjoixp/Pzo2aY806L9Xp/6VNPpda
97zdSYeHNKsNaflqBuSL5XQRah7Mh/gky/SqFHZKMES1NeS16GZm4v/K91vQibL3N4yKxQk5zrhq
WPvmcuLrERfQcDl/ibctFR6NBSTWKOD2AmhJ6a5Mc2wS3qrjV6L+xgXF3rA/PhHIxleYFOAZKF1L
BvB4Euc1l7UMLqbstKpU68nNYXyzQDIx2XQYcRzeO+O0EAYrd2Be73VxeJgiY6S+FucEcc5N9woQ
66bzjwUIFsCAcncxyBKaZjJ4dTxcInXRTP0mzpLyEW1Zdjjhaqs1zbxYinZOuzIqmyn/C/hFywlm
1Z6+zzRHqNZXVXRJvFOiU0y2VH2C121qIQRSg6+Qqp40b0iTPpOsHsWCbagjR3IR7WqDKryZp6hC
/+8lKIOb0BiuRKc7bg1HDEizmLJ5gTmO880gwoLvzdr4XVxfdKMthV7X9ukvQNccpojA35WWLRvh
ZidVzD9ybSmtyi0gVMMM75PuUeFLp0/+f4XF67oqVHC4deBFxmFwgvf9KRNDegMa4P218ceoigsV
wnozDp+NcXA1DbfzRhmQfjvrw0r49H4/yJNZdZpxH/0DzbwtCqtC510+QGELMTN933FhWXtVxZCw
eUiNMq6I12C0+BniMaUijDP8ul8FLD17uHfFGUhGU72BZxLrcxOKRN3G/q77TbCsJ9Uy8tG1PkOl
HddJ/ypM+7iPusqINfKS0MrfJ5MwPob49uEbO0Bs8d5nYgwsW8V+LqGNYEnzq9KuAJQbT9P12U2d
Axfo5p5IyC+OlX7KwkBQcMgrlNjyJN8wH8NmvLdLnPLax4AfgEN2aWcbP/mJ1J8VhVI2LPwjnENF
+xtFRWa6BaGGhOKQUNLDvB8rtG4zdvgZxVXlqfXOE/BADkGRfPaLZSDLg40VdqVyRabcNUe4wdUR
0bddGtge4DUElEeeBxYIPYVAbfWLwo54/OAYM2+rS0c0gpZxx0q+gA1RBT8IXG4RmELGb6dNWwnf
WofXN/FS1y4hvQDsKIQPppSaReYXlETWVBT2zVG6l8IenZZwdrJJvQ+JN6u9gKnH5vUsQpuWYtqH
jYrwYkuMKC/fC6sOZl56XsYE5fj6gWHurfK0zPBWcl8D2vOaWANmbbq/qOpGmfd77pcxYEhrgki8
2wWI0O8w+mjXGZVV4vHryxAQX9+32GbBBYs/EeyRF6P1O2oMc4noFdM+EXe91ivTY62jAARZbjE1
+fwQ7eqX2IQQAw9K/QQeRx0N+ZGHsPuL2d7biTFIVKEPPiYUbMtwhOUUqkVj6PTGik/iYMPNdm61
3qHGFWShAbnHS9stHIA6E+aUG/sPzH5eFYpkTUhUu72xz+nCIBfNiHluFYzfPuv7BYsivoJ3TTN0
rK64mUlkuiA5LjHuF7h23nCyvGhY10iJZ0AyiN0Q4HGHrtP1VkUk9QTHx0HnTbWS3NhrAMZ+h9/J
dP3rVkjGJNl8zZPAMxMrWEK+FdBnLAcmxesNZ8XN8YXHwZJp5h3LRchDCuhVmTnaKf6SIF6Q6/+w
p0AubcrhP+9GBGvO0cv5sZLgNk9lNKCCAebllP1QJLmU5EpvfZm0E5D3Q6MfIOCVEhhNfD52RoxI
gvcjhfQnxVpiMQVYQhlO8vAbmPyyMik6krVxwycZezRnm69r/CP7N3ZwMw59/QCmTxXumAw9rFWS
1V3FAHYIQQJg33d17/nUsvGzCyL9nOGk2ye/6u6SBuhl81/HdAtl018Oagp8Us0SjKIM3Ji1xT5K
kkWhrsSar6WVw5mS/oSivXEiVcoJrgqjwFALSPn7SbFixzLUXju2JlDd99FFKIdKHIknh9qWoyeb
TOdQIgYvUpKrfQwiqyjPu5ELZwHnWQHSCkfbNW7qVU28vmgHu64OULsi+CYb3QcXPPlwD4pJq86s
XYxr1AomXxQw7gh67G8h62zAirbRYAPDTubAD1t3aqpT7fL4H2W2mzuduzud/GXBS4NPkqrVn7wb
Z72REvmyIEBWrVcs/r60kJnGoBW2a96Y2P3aVg2OX7yNg4Krjd5cptyUb65cN5KrrRc0OrUwWbiG
6y8AjNWnPa4EnnCd1ZtojhJ5Gx2TeD/vxOB1YmbLVu/rgR7imAOi+6oAjV9xNT3UlVG8OUXaqCN7
2Ez9kRDFdh8WzADoWNF43HfPUn7esw6rTprhCY0oL1hk7UXCU3G5uXuGW3pvwCsBN62khQZJumyk
khi3xTc42VFpQNWcHu38iK5IZfI0kj9JseWbD9InPFd+iIWPtr7qHtqiQrpaZZyeYbmhuh1feIWS
6vw7paa06lr5t9UXgtVdkfFGLn3vI/8Ew4MzziddVzQ5lc7zB1FrMOeNStOztZbL+H4oioGvyQvU
geA2PWZIpT1iTw+wMzk5po9KZUL2ZZPUrjXb1QCzmkqnlgpAHMeYXdy4Uk4Pcd7hly6+N70pYcjW
3nJvno4IjOzyShjf4/AF5kKXM9rRZN/BkQ4828RTRXSZ3cjDVr5Mlt9wces1PWiqZaWwHIv2LX2y
/OfszBLc0Z401J7KcfyE4EaxLlhsluo841yYmyRWAKcm4kgf0rwH59tp+KcQ0bnUnlVqzXGhcfcT
caT+kpCaN9P6EIgDUdUyQajjoIy/6Liedzu+eNqoRNNKBNz8b7lMCoILXX8ffEzDzLqSnqWDskhg
lgJYDECrW/4tt45wcSbGVQpEtIfHXVDt9nwubs9WZm8w260hEVtoiFuO/6BRK7Sw5qXvHH5A00/W
78ZP0y/X1JU1GE2rocCcQAvJj8CrQuUF1M5BXzCf+ea5JhHUjH9Y/3mE1tKIEETFiIud6/oaB44D
YcSA4wIHp23kbvvmUX0w5WLza9ppMN5KE/ofVRhCo1W4wzegVe6ze0mA9Yh5rhg9k0MAN25vYUs0
o0yTFn9BzZ7dKqKirPLIDg0illGeRuYHd5w2mFzP3YWmVogG0kKq9RQV4Z1/6IJ/0mrAaz9W0zH+
lVGZpn2Qk7WhxygyndKGtSOdREhnBLlcT4HRCx0rfrHAg4bAMzmp6YiTKfVsz/9CxGrshYX4NK6K
RsIHNayF8ZNCV3QglMK37CoKWoVFm+yxIKQQqrFDDlHng0cdas+EEEl80d+mVoNN9tDJM0XP/dXf
HX3IUgYm0eMHPZf5jgTtLYApjIkewTr9/ET4A/UMl2jKvhnAsdIsPt60t8OR1rGNpw/JSxYaRdst
IWvtVIP35kMDJ2EktLuPSwmoMueZYlzFUW7Uyu6QukHF+mJuiRBBF82TimrlCq7tyLgSRdHb1HBh
lUWfcj39R1JqyuGzF1B3vwDkPJG31M1R2U6wAk16EzwqwEsR8cF8c63glLZJNjxn2myfUhRgysCf
Ye0VAoB1sx5obHFD/O6TN8JAm/GrkCijHqShHjYlf26Fvem3kSKIj165Pge4CuPEzQ6aNcqkEK2N
W7rUjm56iZBU+syXnvSZLk7gX06JZbtPSsD/6Rav8mvh6X3v17YgqvWyiMrpyVvwW+YBAqcBizTt
y0mR5JoO+mtLAiEP4IjFck8df7n4OUoxHdrcIxsREgqnnLNz13Ukw/DqfTLpTWEHYtYRwVasXLVt
0+H+9/ZrPHv3mAW4OGm5qhHCyoK6gfT3+hw9EJkHj57LKXIpZJ+TxlVBJuS0PKwWqyzLmrV84AVg
AP1IlDZ3FY9JgLFrGI4IcyamwgloAhhEiGQRlWDHUZF8WPTpjRNzt8SHFdUFIDr+tYln2TaInMmx
q9jMxSPEEkJUDtn6ty1/4PlWkj/XPqDlRe1GKA6k6x2c2eBCeYBDxD0OEEwhZfDZQazUGkxqQqon
bn1lGY9TLt7C3g3Dy3JEXlczuv+fLLq6CawG2ZucGUAUhbd0lQmhtBK/D7VSuFgaOZQPxev9RHOx
WEjWCcuqq0ISjoSI9zj5ABIYXVP1dd6F92ZO5eNzUU8eHh36g2GKhNnkR0hq4azE5BapnEnLxRcZ
X9uZsV2pQEyHQBwUHZZcRo7k54E3+aiYM1kULsSSLNoetEBZ7+m55ZdqxaKoYHQcZr5Lz2Ejejoc
6E3tFEIZvACPqalKQjixmLXCtj3Bbf68PdjYK+sCVfjMpewXOE05Zb5j00MS8t6JzA/j2cqlYcZR
86jQhVv353DTudP35cIFZ8GdECWuDmvlPr8joPZ8v7JVvKmq+j3/LYIBMk6jsqUJAkEaZoR9tHn3
fOC9ehlvngUju6VMY5DFgxlvNwSyM+/Rnxfk+7htCpsZtHBjvo8evfHm7eErXIgI6NxfZQJ3edHf
Cc1DPLjcWJtwf122pDZp3fQMihXd6WjjcEo4hlpt43/sd3CEadbnfPwp6KVR/BMTATHPBQX0T1R3
FlZADD7JUbi4t7TV9M+nFZNNZTF/S4V5iOzW48P4cw4cgTrfq625+xTwJoJ9PrkoS0Wd0jGRcVed
hFxjVpAx3Qz2N/yRIrLMArDi5KnNX8BTCuta3gWQ4wEduSh8PQGy3MoajZ1ulyZAGdIUdd9hws/s
BG3UfiEBz2tw7KFEMtmxgUeu67NfSj5QPAXoUzzVVwcVySvnQurnegM4L8LaRPtsYdag0fjAgE1c
MCC0onBBxJnaov97yRSdBs3kJAHN2bvOXi2BXBfjIkte/WpxP8Y9KZc3Np1JQIdNZohuhiWgQft5
X8a097kl2eysLv+95XaEc7MBiFlym2iBtIFv9jAhmadFOaC0JtKebT/OqXkj6uAE4zhfy+JnGzp9
9ozLGmhmv/5ipjY6XH1INQO8KCVwPautO32oM32QQ74TRMov1Cy57H4NMYln94LifBZWsPNT4rfr
OdZqjB0zVS/p0ocdB7+UVz3QG/okk38jqRsXvIWCRGtGlyyyu9y3C79GZIWc3GEXLMk+kR9q18/0
f6wvLxmPBg6GziwFMn3r0RnDM8AdkowismdXHT2TwRbAAzpPWCLSa+/eHR5M8R0Uq2888GSAPG+C
OxIVym+cje1ejCSX8GXegiEJCTOym3BD78VYLa8aNDXNqOq/19YNfzB2577plwQ8Fk9XvI4kA5+A
mckGhpe/84YBaX5JsA89ygClG49Qj20NzbKK0b9MoVyOvPGccHghPnUtwIltT3672nu4g2UycS0F
AeWHPUYIDvVAgwo+MIHoRhd/vRLCBJEpJX2YF6SPWR48Yf5+pmX8W+lj0mK7dPn+ZTwTNiQg9xu9
LHAF3+2clriYU+m1XZx37+nsa2JilRm47Gi2Hc0CJ/QQyGue0I4qab19fGMyGD10hMyCdoPplnwi
PmZizEUv4a2Q/+60XiPtVvnH10yfDUttYyDAR2cvkyKK6Pe68VtRFMQ8+uxwV2oTW8DMWeUtchRm
B7A1V5nB6iHjWgzUq0iuOLJ48Mie+dsp84/JL9aTgkochbokTE3oxdB6eTt6+NsaSYQM3Al28J8E
WQXHR72+JljJZI4mpBPcblR7f9JwaHPsViDJgAIdVzoLC3Ecy3tco0DInzji0MR/+HpK3nIbDQ+5
jReGshMJxgqCtis0lC8Le0TDXksWB7O0iB+xLLKy1Qn5pOi4ki82fTamGvXRxDfxtgddFTDnVCmP
b3aU8o2ylal4XeFm/yleBU1YupWRXLr6dZfilVddpp5DIyo3lNAZCzGoPyKlc4eUNZtMea2FC38Y
rCj/kKpDGkfRksaX0gyraoRP+02BDpmGGDr94bdBR3DlDK70Gw+yh7/6wpNVcgxwcInIZ2McHkAQ
ITsPj3xoNqh/0X3RGp4QxTfSermtTIw6a+RQHH0LrkjbqNwLTs9ie5n7lW9gBu7bPta4Htb011+Q
IXz5vGlRSpHPox7aMi/et9QrJ7TaYsQyd6lfZrXYtScF7BGVcrTmL7impXSdYKPVv8CZ9oGqQAJO
eHZTJgWkphghNLN3gpuDBR3UJdmECcFh62miv8gpsJwpUGEbt2C+VeorNHkZU9hY8PDaKv+RI3Fs
JGsevoQAkQCTmmrix9WnExT1UT2c8grI5k5MnVdcA+MNWip+4UfdCmRzLe2DqCNnP0qHuBS8rlPz
kr2Ervt1uAsd3msi4TWXEnU/Cpl4x2ZYJpybRaJHObC3Rv1Xw9OK5/pxQJjwVr9yXIR5pb1wOk5T
lZJ3wuUIkyV9V2bZClxB/6Z5llK/CAH5bdisp859UEyzxsCVc0HGjeo8ZwfWL34oJKcBIMZVae70
EhZia6d0jTzf5MtB7QKLorSMnIxHwmWRIMoVQWWS1w/CcP0qDrLaoNvY6HdWGqH1FcFsgs/0pvN/
FDmkyGxUUgKayZow1uwhZ0VSn1CFYbm4l4iboj94lT5/LvkIYw15wLkkIOJM1mM/RpD0hiLls11U
yK1af/YSFHTzZTCK038Cf4pVhsKkfUA1lCNJFTUlyBTYm20SWOQx1NqShOPeoNLR96X3TX/xn5Ww
ViAK0bGXUqHNj1WpX96XcmXrKLA2eYoJCNyt3vhmiKpacaKXnQflqCyc3ZQpn/P9FYkxRRCNifSl
T3g9LVR39jOOJL5UCPOgHwdyY4N0MH+JXi33ez72zIYL5uQ7yz650/jGI70o8FkoDrofs2VEDKxd
X99dq2PP/M1BNWPMAhvY+gY0UKD8dGnfV42MsSzixm69iZxJfQ08Bov0fnMA6c1g+COUiyQzId1z
UzO1isYnGRojaVtZ2BhlX8ZBb5ZNN1kReSGWFqvanFzkMc/6pgGVWUIMyOK4TpUBfjtNkvt1StNR
SsF8moRzUHUyeHxVkEWfWuZp/bfsGhDpkchBB2Td6Ux+6ObIc5ib93Kh5vnygFBJ58hJ+/Ozq7de
MovnqDTZoal7vB+k1wp8Go3hTwFWkgHxGHhWa4K4AGxpR5rZPCzMTXiaB4+0f8NdnHUUXLMtf4Gb
4bybykePyxnkDrnG3r94g9sHtwUB4aGDE2XuFFIPG3+glY9kmhOoVxopGhKjgnNdR97uj4M76TOo
pxIw6V4/zOORKokzWFZof9VHlxYMJPMBlIjz3vF3V1fVQLJxAG5oEMJ7Rvrw7M0AQg88nvsJl+Oj
FmGgmyIQhIAnrsuAsR7vIhTDp8rkmSekgmlniApr4j70wkeERn/bm+t4pGzMmsHSCnewvPPG6ds+
ELds/GEOF8/hFBtJ3J4uvPsq1Sbnh4A0sjbcGQu261hVoEHVMWw/QZ7Etx4ocQ2lCbHrV+ObmaAE
zaTj26dFB8Ck7JC9p+XIrzJLr0o2H0anDJqB54q9t+77X/ogPgS8nAnBIVeJEz5OtL9cB76rhAKQ
orqEK90Z1IItz197sPuBDshePNYrPOw49E9H0sqlnbOrC28jepb3cFrQX/27TgYMtqtBwDRb1/Hj
l2Wm8KMQDZvwmNiwOfTnxALW8BAGBcweDpaeBNSua62/mspzEbaLtifpt1dMfoEMae5bx0+J0hJ8
/bqZjsaRGTkiKAjW8b/4UDb/lc1vpegNxpyTglBC1jkT/Xhg3+2qhQAReH+yZKr2LT26xXEkyPci
zQVRUZfl0oubHHs7XSqn8GYHexiAYhX/gqGeXuXp67tTX7VwYyceos1nkVc6yS89UG22w+vO2d2H
bOL1i0r6qdZ/5aIOUtRp3lEvyOwpmkZKrzhgp3TsZhf9MfV/uVXG9Q4eZIh/Tnr9hm4W7db0tHSk
jRczDlxO7GNIxzmG+CScoiUqRGCzmV5lAxudkA2DZ/ih4vRtzM+R56DuOuh8nsXfDTiJGCgkwLvm
RDVaBf+nGfaFplvYdonWKha4ROdGQZv5BelWVAwfbRUasKSqTC/hxGKu8KmFGBbvODRpgS4AaPSg
rooDsPpVaWEI0OjJ9bd+f9/D6KyEOHwo2aZZfp/779VeEtq8L2qzROauWvsca0HefNeIPHKFeDB/
UG5Kfle7sY3h/H474Kgt1VwYgsBsJy9SZFRkUrw/u9IEJLmz3Na/ARtTATP7FTNXtCVHMWS90blP
QeHzcch81oi47gmO4ZGu1vVp2Ioq/2Ww6jw51Cr3ZI7fhxZl8FKEUt42Og5MDimNFwJQAsHoFNEJ
1O9Zz9x915RxgjBsoJe4pxYp9W9wjJVOtDyP1udNWlABeTJ8prUk7FEpabbT/IbbnSxMs9G1NnTu
kDzk1GtNGGR5plOPgUliQ7GBSFxX+qoAjybbGfqnwpMk9YCGEJcM3lZ0jZSKglntvt7b0dS30yCd
6GyFm+MzA8XUknN7jMqP0i/DCap4FSrgaTjmJo4CmSUQ3w5e+FhnnN8nTBRZOQty7AABdF/jAyu0
5gqbDsdDZOF6kAzxwXX3ou6SVSgDG5oKJ0PSL75TW9nOr4fZABKw5Su2wCWl05PMWCGhd2zIEaS2
n1uVObHYTpZ4avi9PH3DFFIa43Ssb2EgTttzLSOJgAx+x5IsHY80CqUb94782DhVRy37egALzgZw
asW/vttENNh1NO1bHJh3AHCukvV8fhuoxyobiYQsiWIKD273EZtjddXDQj4IEz36H2o1YNIisKmV
gkUZur8Nl1zBcRUlLxdMwlZQoKTg6qOOPza7JTHwC+wQJjS9wA7kWKRrrWfu8MdoKI8h6cknZxJs
DQxwkwE/e9WMQed5I6iI9C7o59it4KoVIpWxZyKIyh6XRT7CzBe/GIX/lCeofIiF8wz0/F0gvAQh
avysOIRiopwork3Z8QvWqjhIo2cdN3BFYxFuiu84jDMD/CpsN2+E3wzlT/bQXdI4wLh/YvZtBHlA
+ff4Y4FAkra9oaf7R4beYh4f4a1l8qHz280mRjmVNcUrDlByOuLWAB4WuvCGs4Tslpv2+61Clssx
HSksbEinpkGh/1jttMo3fyY/iHmuosHOd4eHG1zo+FxS0UOJhYvPnHeOArhNYgsgQE8oCGNkB+wT
H14IG8f3sicBeK8mVfbHPNznIAMVcHWYdZgiLp7GHlJKGrEfdLo84I9vS0CoAGJbau9RIGm2Qo05
OTAbe1HP/0KmnLx9pReiuVnKqrOjsT4/G9DtnG77qRe+i9dzA0yGPxodXTytew6KsRdjvMa3An9s
Us3gWlpUcqxsoy/y/XYMUptFN7NvF0LOGPSILw2PrceS1LR7Ts9Caa3gwzfxoBC9rR9ZCGpQKLBU
GN4b9VU0Wumky8nIfjM/OeKzq8dT6rFfAJRUkpLd7gkmUIEUYIAWepqyEWFHrqUXVAYgD9gmdTKz
xHMEW5CJ9LwSLiCS/usbZnWLZfSlzw3Ie1EMIdlCJd5ingTXet5xtNY8ZpbiSnXQJcyA0GuQpJHo
KY+TAjMpZ2l/fHiZp53yK3i3bdDZmPV3zqsRKjbdVXLJDX4ZjLwClwsirzZzIt2IB07k2Q/ad/4o
txKq9350FNl9vWIzxiIn/pNQ41x3YhloK3U36s8F3VJknJrwsWweEEsICDu+vcULcRChSXqV2YUi
3+v2FSKuqxPZfnqQRCBqUTWncAWPidnuu6heejh30MaTFNxy1wz31h8SRt8fDRyN82ACzMNC8pRz
7Yo4upb4U7txaZIw427gRPK7Gtr5sLUVEHDNmCu3YMeOVgK/I9rl+3PjxtyCml54E0C6uUURl5Qt
91GNmhOCzCf3vOtipLg6iqJRetVPjuBReSoTQl/ghz6PKQUkVq+V1gI9vXejR3UzLLdtnvxpRDbw
2KUSZTwt6t1rRFdkXmGMZEWrrSfbangOrlEFbu5gzDikqaL/QtEmUmQ7V06Pz6ERlG+otHPUj4ww
7JeEKxwgr8Gte1FE8r3IT/TpJP5dKywFG0iIU/4R8O0uLapulGG+22v7aTOd65H0wJCUgmKoQrsN
nV+U/zAvClPgs7ocberFc0KyAjHBg33Zxlyto25KpS1cCSP5ugj8fL2/T5JY2+HeL62LLIXczkVL
fPxEHozyjvMzpON72XPwcw5j6J+1pr0ADr0TMb9uT+lGlnrV+0tamllJp7MWQrkcpFHSjvTlKcpq
gHoXtk02rkJSXrvJQvgKOfbSy39Qipng9IEMDbSLhtob6LktMyj2DFVbBDX39E6NA1y/K0t9/Umh
FFt9uYgF2OtjiFhyNHuXn/3PBJl5m2D7lqHlE+bGoZbUVos9bETxY+ug0bzwPkCUITqn/B7QKH99
pw2U3u4MyBwOhCZEJwJeS6+onvvFpk1r/DTKD3mVSGNPA2odgv15+QVWoGCxddffCdq9OdCwXXcf
Q3bxAXxs4fpNTj45hwPHhY6WpDgN+vXwue/OtaJ5svVE9o3gZGIzwzhwJA/OPoSN041NZP08+f68
eN6ozf+7MImzWIXRa/eZW/bKp53Onpq5DsdC4Ssgm3tQ9Oajw99TPMlFRlqesh/S6pEKB1yE6wdc
aRUVZuL7zD+laq/5Z9HAzkD7r9DYa1ezbWWtsOU5gAW6WApUs9ooKl0fdL1mTuLVYcHR9i7AwVr+
8uNhFErhviJiavxMM58tKE/DPQhk2pQ2wTnIbFOizRVL/DPdaCcUaLPYUcbzfEjFi00AXgJvJfy5
QLTAnpEK/053abpWCOBsBJ3e8ANPip9DPUwrk5AjuNvb/+p0r12FvFpcFNA0XzHZOvDXEYbd6yE8
Zu+YrCDywwfFjo6ndYADd4slSEM6h3joYCqNxMdUTjxGu3DVTbo9dBCJ128M8YGcj0MrJTAfknF5
hWNXLTSeAKARz/sof8ps2ZJIGiEx5LRSbcoT0zk7XATn3eW8U8DPyIRFFFnonMIv/CS8Cuw1MaEX
6RafGi+FNektSwbLYs7Jmp6FbPIWy/tZHvf/GVvNtoDiap9sTe6TTCSpSUNsFvQyKA3FSP9miNuq
vS9wjPn1MbifMDJhhugcVZ2EdunemGHF8SZ6lLvxgxlJ0eOVT6/jca6MC2bKMPHn9qKK0Zndf8RS
pt67OWdn52IDLXlfCVWI3x0N2YnuvNbTh1wPuW2VZBx1bevvsrikE/sJ6EFLEUjrHriwGFDs3FbZ
nUsXjLyeR+BtBtN4w6/ubLQDaUnYys3+cB/IoLc8xgu1cxE4dUfjLqKjPlZTu4+Q9hqKFtj7z8o2
+RlmzrITrvA+z76TPQCpyEiAkTLDxpczKIzunI0MG4F7q0Runu6HY18fTa7rQef6ik3gn9toTaUv
piIXD0xyDaz6aijnwRhboTBaUIBJaDkzlICfTKxJyk2248JNJjmxQ8gXNPSu2GCiDWOztdkX9i7h
w2sfuA0yF9cYJu+y4TEfjITVTylHslaXwHmUEk6z0XM0YnGX8jvHBicENer/c3urPc5g8wHhNy08
AHwNK4Wi7UewAh3w/G08nSAGiapQXTrLFvttTAvgj1HtXxu66ihz79JEYtcyQY0niu0SeIbNeQI3
Ikl9wd8ePRNnu/QMzpSll/hzNQz3rJtdDEWVt9oCOd+Uh3hgddRaHhtYOjLMd73RXuBfflpJdZN6
lrdZXGqmnfLfiH58GMQIMZGv13+ZPrgNdi+UbrpKQeLxAXmNFoIdznNMNf1dnIb84J7ezl6CFBMf
7q2UvFx1XNsSRvWDt6kTXgsADU3TAJmJbikgRJym7uxsfB+Q3VHWxXEGQUvqn/WiXaAj6ZxeqqJX
8MMJbIgyYg/Wy3XqHWkRFV8OapXzVLwFcBSvFHfAFCvd+5vCENa4PQiA0gTyNeWeZoTPCsS3xWWL
aM/SSxCWqfqHxk42tyPczmIDc8MtxqCEZm6CujTQmM0VV1HcQyAnMfidj/FA88XFVMsMeKPav0BZ
TwDbODy9k/Q+awEC3vfnAr6OehCGYblPXBqoWaQ/Dw0+Dm/WpnIpB1YlWzuEV7ulb23ZpfS9z6V0
+yLbLEvcr6/JZ+WlMgjdUj4H8EtQ5n2gY6oCQw+XEViEMOblfttIcWFlKdVfpqQs3ZugdJpeW2aJ
c6bgG8w9XrANJLiLdBKFLm9iGOhPTxCJZB2fPXEIzZ73VGbjS1E++9C3Ny+TuqhlsfdAfQTn0bnk
Xd9r3/wnUBLUsT7h04TGGKHp69NFwgKfT4TTxTItgu0ooN8y164pxqj9+qHQglI+RAbeTPJFCzuF
cVG1Y1crj/MdluStUQvGrKWCh2Z8r0Y4WLhFkuLP9uU2ZbID5CrtNlFbgfPCFJilkgnDHc5IVs2n
RcPx+3b3AaPAzTeR2Dmq752RNc/8ke1ohWHCa1eLzyuh+05bRiiPmrpQUK05sGOh6eCT2vwnPpRL
D4HYhKcjPrc/fUka6Rx9EPld7B28g/6uSImWnSKHn2jZbp1FZhzPYgOTMvMCEWrowTDOlgMjAbcP
AdyMjFXuKwHnHA4NGEa58MWo9GtHnc1SisxSbEa78o9k9sgWSRmKnvjrkFEvviqRFgA56MCYDzmo
7+fx1M8Nt+Zci6T0wHMz3Y35t6axzXWkjUST4xPWuMEyy9yfpiprYcJ1hW8LCCQXg+QywcFuq+9x
Vt9Xo//HlGe8vByBRT+V166tm8XJQ0w6S2GmQt+mfU13zWGLHyQVVyN/MbryvYQBRmEJQr1WvSJo
ZpNxF0m0WXl6To0JswZkKBsL4crJv/INon2Go6F8sgfXE58yqkRVZsTMCyNOgwO8jjx8S388fJOt
B2UM/oruyp1KjS+V0W5PFj4eKsNl98tgh52INmCpd/JbS3Vk8QbSc5/hfJfCNli0IBQWq8BleFRn
Vsni9ibMaraaK/3d24sOo8Puixe0hgkmN+2J+rmfOfv2ipgqFHD/vuZMipNW/oi5zWCa7myp9YUc
1TVSQDOJRnNWl9jxa8gC1COFg4e2h6DYzXQIu2UHMdDR4X8dFgBC1ELuo5R4S6kFLe1+/vrRl6pK
z2h3T5+s8oPB/NA/nl1cuy9xaksQ9pIY1/yFz6uLgHAa5VoTp4zI3POrl1Qo8r8z2Im5/7Kxz7YP
JzoXj/pgpcg3+eWavuU1eS/twRSoRNMlZILHp3UPAkjdA0qA5bD5/DecPnBEDmzJvkW9lb71/cvm
JYwR6aIKdhk7U1ZVq8+DCgzq1WAQp8GtpRkD29eRaZVphExzz4w7o6sOps0X8ysmCmFPZ8bkPyK1
+uKXuT+oQKhlDlVRHE/Kp5/S29NFLes1cMjvKRVN2XvMVk5q3f2yUyjen8Ym5KVj917bJSWyeWxz
2EMPGAOm4Ecg49snmXN0xw3jXnKKbsgZd2rLjxlEInw5y9gL0S/xLk4gw7HhZ7Pa1nMqKENAGQK/
tYjRkzhWnvntVkcqPndqjoWROtuUY5UOKdR4m5tb4NSA/kuyUJmLNd+WoEYPADLe1b5VHrgGUGaS
sHeUdjKrz3MnbxMmd/898KmYJTu/JlKQORgNWXPdpEmV7UERwgnz4ndDKz7xXnCu3cQBufFbeJkD
WMq6bliHMSSXALo1UtecVJtyMQma3QvuRXQW3JB+1+7EBFrpOb75Cs3ehjR2ZD3volHvYkJ4MChC
Rqr77SMnGR732YhuNt1j0voQ3bIEZlXd9faG+HoExZMu/YJD0p/Q7FHOBSKx4ubNV7HUWtgeRpWs
Xts32bRpWr/WtwcCAA8S7fcUpyg+yLPcxuRu/8uhU3IUzecfCDhIs7uZouy7e7FpV7fhBRXxntCl
0HMTlxQoeMTr8YcOV1JsoMX1jESiUpfVrrMJl17sO0uvzzLchvtvFG1YoQnNUKcZEgDlRXsNr4Vu
bMKn1laYqbrG3yjkEhWhXixfljgjx/XYRQiOJvhTqZssvCnt8tWRvDWzFxJzuo3IakjNUDc99A01
QO3fE+Ty3puQ+bVYrMruwWrQLpnVV+BgWhGNoOBbJWCOko1ENFPePmdJ49SDpOqEGx/3S5Ul34F2
51KlV6IQO6PPmGlCoU70/os7397krfnTGtnaLn6gb9sywyrJxZohCbcing50z9h47QVdicr75RhJ
2emdXyHCZCPHrepNudFhav4TQq9A18vm4YABzyayu99fyu/94GOyI2iZwGGZFBvvbCBFFPy1CPLn
drhrbqVY7/0CVohWFlBc6598EdjFiuhggTKOWTijAIEEsjuR/EbFqMcpjA20HIx56sZERB/sc3V2
h/777fSLFkaGPqrw3QBVDXhCFnSfZeUZbz1ADojb9StMQOdt9O8YL5COOcaQB2mDrcOhAJ+AFAS/
jBd3m/yZajAxeCos7lfv+GoCy1umNOieE4IaaxWBLkjp6F1bhEomOlYlxC8xEBhDZ5lDZyN2rm/1
0vYv+YS64XUndRqeNImcHBipBssCz1PkB83YgD63rJ+YCe6hXg2k8WzA1cjF+FUBBhGB2vcTezPE
fHZkedvpVbxvqvY9aJiw7OhT0acNlGLkq7KiN/syGXON7EFvZygGLdKP6AEf9+lK7qgF0MSh5TGz
dZFWSy3oOLOFiW3lfGE4IszbKd6N++mTPnedjKsssLLB6/WbQyPj3b12cwxYRlVQ53DPSKAryX8u
LEqwYqVgiTu+yoCKxVXwVY/Vm5XN/psucznseKvgdQA7EQkTp8gBFOFSQ1j8reZS5sEZNGdwbcPc
veyGRQOU6sOrQjRadan/gwHznXIz547DGamvYJHpyZILK/rR7BxmQrTba51CMa+TEK/zkrARfyX+
GysWQ1fhZ6Ix2viXYXfHfsEJ6cMr4u8l07vNR7aU8QfPfQz8wfs1WSIg0Enug4znqJ0l3zHnDt7r
SCRmX3rFOTrkhbRDqm7Gl04uNXmcgZTfcHv4ga5QrM+RJO4YePaW/TnLwqhAiT/osy0bvQWgSMY4
gfNchR40yhikhH5LEUO+imiN6Blj2HhfBM0Im5+E/EetofMLavKGMncUUVORPQv6VAS/R++/LwKE
dGuzDzIwl36jrLUpsH+BmGy9QF5URmOTg5tMjC7jtAly46NToCV9D/tAWHmQngKz4rca+04ICq1j
ZMDnyECI67x/WPrYVPejkw4osXtuYxVpYeZjL7MHXsMPVID/Wodxs8NmMHKo7CekYuooWK0/CrsM
N6NKalZDlvdJ2Ys//jExQ7Ej5hZYN52b7d7t7djyTDNT1IX1OQe6bvnEcx1doNxe052tta9EtGl9
eTz0/rMC27vGOLMhXOvkYOyr2UDj+cBNo/ntH49XySkYi8YbgkegWOUig7QFTVUurM3Rh4nCdNfV
8ff0MMEn5ofVHjA/bkTojsmAPPvWGAYJflIii1S59VnFIOwPAK7Put+ryToEeYJnVL6/yGBWB2WA
7f54xVn+aWmJqZprSsfdSVyshbx7nDGaG5KrQw+kRn1T/wD3D8AZzGUZEQlW3rJwV/VEvhD5xaCJ
TebdkIyPkI8CNMt8IxD3/LmqGSA+cvW5e9Jnb9m/3clpHtGqWobeoaErGXp6V/QCRRu/CHu8gnYm
WjEPXUUsfxv+X5oAqn+VPvTvJ1BoOJLfAGPJNchZPrEaPMGujs6oQZR7IeNvno6B6RZqPfxlFKwL
CQSU0Dq9OW6TTY8pbZDbpsUiIYfctnT5U6AD3ho0HFP9PnXBAm44iGhoqSLvIhSKFjZWl+665O8q
pgDGu1YxoCiobhh7tv61wAjpUumkdHLCWLNnJdzGOSNlMIbapgxo3ZIVOZ954IoA1c1fDmtiq63A
rL1b8ni5CTO0RKL0aO7x2iqHtXeCxTGSzvM5QKRMo9gmKYpawHeNAcO5AU3G9GGTFKzBtr/hYCzs
8pGEVfBo8K1OYe5NaTV5bchG67xrZS/KxsJDkfCfrhPKmKbCw2Smy5T+VJwuSRY1DCF2jHGslRGe
OFfbqxmmhqVAnt6VPD5fG/h8MsbY9SQ2pTcKy2Ve/T56sN0Vstl2wj7b7yYoxJ3vBP0TcRIMPJm+
HDpVxV909zRSWhhhrwlpuNnh+KyRFVChrFEq9jXeSeI7SUGkH9PwgPPeiaBPZKZYTLp1VY69MbQA
M6GH7rcPCZIkxtirVFPiWtUwLmC1uorFblaPKPnEvtioT2DHNmKqWCDcRkyWFK2bnpemJb79jQXN
3IRjRDiAL+0V/5eOfATEOSqSPLff6QI/4+UExn+4RaJWpF8YWf9fIEAOh1Ge8xQ0kNGOH6xH4Rek
dWEtJe2W8b2BFuynbE67loeu6LewqiQaXVjair/PeLYuwIkcvJjsuYIBxjT0anYM1p8FDGeZEUx8
e7BTBgubF+zzFlblP5kZYwDF3BjZYqe76/k7KGKh717p5GL0o5hdmip4+Qato8i9WdShfcEm5baJ
UDYwvZXZN7j/OiemORkI8dqdG9iD5Y/yWBagWYvCGfSo5xic6KhOg6i8nByr/AM3ps8VLJBNRRsw
kBWUUT3rrXCUUUjtuWYLtojRaUxR0urGGNeOgu4qctohyeUZs75EaAiI2ckJC7e6L31TkV3DAj81
TKllN41SjflQn4Azi8nsBf0Us3ylx4TXN8fdGtpfABLO6kV6CfxP2bhJaXWtJRK036qxHgGaWaSM
P/buMcgcXSKkXBjlcCkyFs2U/arhlo/Z+vCc/PhRXgZMT0TLFY93a5EdG8yn4gHzW8M2iddlMnwT
W9eDx05Bv1mbXlyiTOjbRdNubvgenD6clW9wSOLTcETCSHi8UT9M9tx+dZJAYtofN/6EDQa4Id8x
TE1F1XvJd5m50oECB0DQdvE7JYZqnPlwS1oygmA+IVzznCw9ueQxN6jrOuGdERtjdDVePbvD8ktX
fGN8Fm8dwVoWU8iEgfvyTOAzm/U8FdfNHeyhoezBNjVZoXbnkCoyhsCQuIwjY3J0zlHFNV1iw13o
qCzx2F1JGgpaclfWNmbEimmjT1ZyASJX3y9wHhVEK96vfOtL0AuRGxjIwSfnKzJ4fUlF4pq+4FO8
j3ZlgaUNV+emVtR7Z0tV6a4prtoapKtiGClEMNfSUhf8Al8cWjGmpwWe5w3JUQ5sDtviz2LVyk+H
jd83vH8QxGxVMKCakzpQlbaSIdweM3jfhTSkTvKyyZLZ4KZz3aaAYhh3+pDtAAPavZl8oAkF0LdF
Zoe36f7iBbxL8UaxBkStbl14Ab9+/TQj7yPtyscfWPbz30/HpZIo+KozVzyhfIdKGzGR7HDXYVHG
N+6B1c1G7GMwYO7ScslFrplz7NqNl0/U4alEhztTyiJ1kcrQXOL7JfBNdG/AVNu6HTcdwy+zXS7x
xWpDzfoWWKq0NSKbcfSvkZ3YCjkIuQQNZ1gQjxupknxK1kAdffcH037ai1j2fTZ0n0dkBnMQfiuJ
BrzeH5FfLXHDjU1hJeRnIxNhVERpH6LPXml4cMxa+mrTOXj4s1y5i/NhlzMRmAa7XKmigQpnL+cJ
H8LQVF2/obnEfzYUdDm9QRrVqaIWtGE2w0h1xdLGZKsTZIFaylTfILhwqlLxsev7Tm8k/szbM20t
Ld7Y7WRv3D3RSIq9rZzMrIMqAd/rWXPzzL5SznNxylondFfRMGnfa7ULeHCj5bQ3EKyguW44TSoy
YX0pat38aAbsMzY/cThn4Nacs/BuG/xq/rL0fnMAdP9DDf9QDFiiigtuPjB7aJh8EVVcI5cR7WdF
haxJAm+v++yHGjXpr58x4viIf5i0/Dp4xvzKrtO/0FtyjCTTquXXOW61suCXUd21ETtedPC4lQYm
vVxqX0b4Gm6CPbcn/P+fknQjmqJv7Uz4B7qvtbaSltdc897pumbrYQsAApU1o0anMociE+5i9q/w
oCuJTo98CL2beWqZ/i4dZ3aWp0uYlO/GKlSzThCNewVG5hzXpYcl93S0AYe+3tdImMH8z09Up9YJ
iIaCxOaBRXpRcOnv1PZkGqYygFqwouckZTitgJBP6BE79sRQyw6DjSAoQX7DpEj1RWmalFDPz+/6
hneQ83RfLk9t3lr1Z7D6Gw5AxFNT+M3yuWzGAtKsaUBuE8LE5B+0HRitQ7RHBCJv8SxCnYTwiMJz
ScL0GxMv1tet21p6s8zk7bQ+x57xpj39TdykBKP/KTtqUSkPjFqUmYs9080VZOZqREh4wjJTuIJ9
6EUv/yS5lDpvkLoDSLKomE+r/byL0Q2Z/v5GeYPqciXRYgqjN/oGOROvP9C41764nBTu4C8gt+Y8
I0Rn7Lj9L0ADnIdSR9eJ2JM5mf/TXrlAmE76t1bMJEs7JxmkQJ/Y3I4UXiJyV3Qx1J9CqhNvcm0I
53bF1OyFEhWKPHF8wxfmKQ3enigHtYceJqg/mL9X31Lwd/jlCRiggAuYWTZcPfNPBGUES03vnEJS
3VraEPVWRbqaNgnEZApp6nxzb5IcgWWWzsAkNxPerSskV+woTnT8ueFMqeiLk3VV51Aq30Wk68QA
HXAXlSn9evMj17ODjdJqwdijQYbCExnMmdnJJKTzaPKMHLE2GhV5TDddbuuAGmhd85cQRMIDQXGt
C85d5q9Nutao6Il17IGQ1jJZLj0k9DpVe6nfw2N//FAoA623ZwTw/U8mYEd5QP4tlDmcH/5lhj0a
DMrjjUOFcs7Rkzw0DqiRRuEtFVFuK/P+adXFvkIh45gSuGN+M0z+3QXNd4rBULK4BlEF0cUWq3FP
ZOn8tK/NkEmOqleWUB6PiRHsIoUOzkdUEducHOCcS56BjVzLlUi0dCEoz/j+68V3XKfFUWU6WEgQ
gPH2zA88gUBHhSOxhc2BVc7nGOMSVPHcImUIswyGxNuKj6vMYlGZdX7BMWTBk8XzO0MVqYnrvG9M
SZ8wZ3FrpG9U2oswb+AWr++RIJaYkxtkKzNBZpo0RLy4ElAUz14u8iEuUL5H0jsk2aX6gUYekaJQ
AEydbpuvsx7TkoFnYDa0k95J/GG/nbtWKKJ73p/8gF+uOhQs5clpQ9jQPOxy5tj+nflNGdeTCVcr
hZJkIbfB8n1hUiFYS2lafGTNWDYaCrS6CXQPvvXTQbQYNI166V6eRPhlUANh28h7TokK8gS0AfkQ
YDCub7bDy7+sA3aWa8hYuggbLA7Vg2qkh9T3gEYuiWbXu22ycdCbBZ4izsWIRMTZENbCbybxEEl1
tntPY8GwPZGPjC6+R+xHI3brnQytoarXxfaaPr35E7SN9ETqGvS3vgTOO2c+bj30aJuBapT+0YuP
l/jC/2ADRa18+8+ytp7Ob/nvziBX0mHSDF9fosKTwTuM/f7xHFpr4x1BLiyD/PqFI/IBBbkTtBuX
CCXw+zYSnMwMJIxIOfKtzLFM6hz0210GkTstVSE/US+Dojk+vxSLpv/sFtxtCcjY/DdbXxAzqJ2L
1nYAzSV9rRKZQ6FVjJYrXE6QgqWIIIlOzCDJDiaOcCU9h2w1ZcUaJuH/cNK2+fBKR790B3YfkH2X
o/InbaJdInLz3teuA2WxTPtU5vvvy5ve+0d5rBNwBe5XLb9u0dX0W8zNxx00VMg71D2X5MwzheJm
Ap0BS702vZd5fh5MKC0v6GQQXRypu0nV69B8pz0gVl2sek7ZAZMAAQBgKwDVqwBAw0RE7pRJnag0
zJTHiy+10RYGrVYShe6RsCGRT1ULDQFkIS2N9YNtH8NW9ii0krF66W3XhghhsMIY/tav8HtDufvc
3S+WJnenYDrVPnqe8gIVQ8m8TpKDU4idPE7IqmCvs60cQq9CfWqcFZgErQnonF2jVXaTrmW3uEux
5o0HeGubpHE114wVm0g1GnO1UuNxTYHj3WvKv3tlPPUZd8ub2Z8J4Cmhkyz3B1E5jzVZbjkAgQgW
u7ILj4HLWGBfMbfn07Bla2vhjBtrLA3mHAGHxqMc580utgG7PtUaaeU+3gLQBGOu28l6LRaPilAU
1MW7dvkSUqeF87F5JjrYwQlWvtWf4asK8g+Xf+VKPy6LgFVNbzNOx1TbN6F/LQBnKSDaea+CbP+e
ORepZATJ/kDmy+aqlvdqK7n4tZrOIohERXxOaoJ4dNQnwCKlSRAb3y0HbFIGVYFLtb/F4DW61ehU
HpcgboxJfKwq+s6B90sRGpFye6kYMwhFxfmmcRfVjkYTGqRgS2uSt/0vM4j93NKwMDzzYmFCBc+o
HJ664aHgBJmLZLs7dNyuxSmVzxtU2Wmha9DK/5oHY3SwjHhvgi/G0TlO0IWJFRGN3stX/lXraFT4
bR5magN5h70m68C+NqPt53481DzPeKfOV2Ym4VExULGeAhfz3CVuSo2+r+7tFHJ8ZFZSz4JMP90u
JQ+Wa/qK+za3F9jVwNm0TJ5e0dNwUQPlpXhr52gh4US1dorV7UhYpA2qrfiRQTlHGm18JXd7UGyV
JgrfCumhT3OzXsiMU5GD8goCvg0Fo11sg5zgTna3yKfatbimrr79zW0ryyYhd6KCcHaPrgwMaVZt
M0oa0/tMXKq7O/B9N0pQJ1iLO2w+av/GKdvyPnRkk6SF4xijxHYX9yCCLMj9dGJkKFD2LAn5iyMc
xf8gwcPKZmy7MH1/fUIVA58A3EzQtEZwp8MLTSrDxtfMiswpr/kHUeeeVEAAPPkcEwquww1DWBN8
21UylcfpjftKNbxVr96jFLNH/vIKTaMnk49cdADU8BbpRR4i0Y+UVq0YXhuIn4vh2ROjKSub4pgQ
9RNc9qE1SBDdr97by7Fe3CLj5syO09YlT//wVFnVdRcdGvLwZ2a6ZMuepMDCJwXjSCqDlLh+X4nU
abko1mu10MmbWDYLndBlL4oETk+l6FsnPCRCl3iNeOpIbfcqEZZtaUlSpRGF6yNSWN0bGQNBAI7/
xv+vI1+3ByX5jZLSfsH3GLd/7FjrdAkXt8bFv205DuQbazuB9/lWdjcGxaxG/LR5cCoJiGg2k6yI
1MxdhwjJdnMtDEkGhj+TAlQLnWLDuvNbEXb007A3ypkN005zbM/xtouZWa7CZhwF8vxRrJZ+RP9M
vH8U6hwdwTZNwNOp8QOpsCOgHGP9osocMXg1BC07fxMCkZFz1uwy9mvPfMzg2n91xx+X+IbV60bl
FjzH41otXwMn3NZL6q/gqThZoxaEw86aiNIoVH3TMZ5LsvHmvEjDMQxALzFpdhJ/xDxIBp2QGXx0
po3xP5HrnX/msf8p+5B2zKL6bZGv6eSTMFeyxs/21Dp19bShv5vyU0k/qJ1f2iVUTWSWwb4hODzP
pPh514yBvdW83hDlhjcZ1w3acrixImVct8P++ImcKHfxzjCwl5eKN6soxhF64gG1aqlbbw/pEUbn
vADmnHFM6Spl7EDVbodR0yxsg3EjEaOflfxggkpJU13FDLs4RdIicE1gGlE81kFVTMKIT/+XGOlY
sSEnmDrJXgsfz/0tUVdvhl3wdbzSdTJBRfoZJzxtblyRj7dGVauyD3ZkOWtEMoqxjlsERQT334jj
JKi2ACVLGoAfucRKbC559rKRdKT885qNSEumRAu3WA5t07M2URr3rPdwPk0suf0LJpeu0Op51jOF
My4GDoszhZ/nXMDeUjCRjKlIdZKy1qSe158cyxJTVJwExe5syyo+0x6TtcqNWBlYovqiGGKQsM9d
F4TcEFgLhJ34JBw9d7eCsFIx2GqA2UVg8m/0usoRpIwEZ0hhKiyTBtGg+vugKUou2J9/8fOyyWir
vqNZ+AN2Aq52/tQWL3Zy8LwQSicepVvtct7PWTB0zL26kRQY5hc3P6NvOef33bu2YZEX/bpon+rj
W+kDUQxZvn0O39DMO191nyVvosCYqiY9dIeU8Mqu9Rc1Vp5y2l06afnnt3aSnyC5rE174d2ntDYp
zZNxiFPQl05V8qJs3Cy5QUKYev3YsV/V5mtUQSXNOvN9LhX9/nyYz6nlG0HP9elduJYd3wjL9OTO
gI7oGfAmHXu5Xip5Boz4Wt+v1TTg2fZd5T8/UjuVwmg0RMhRHxK1JGvmdLji/NGzoXxtvdy/Dtmg
e5dU+pYY8DNJm5ReLz3HGp8CpJhnOVyabCj8f6+u4ahzrR6UxlEBamsb7PZOPYSKtsACJ0Afb7Mm
UHuB0s2N3nx90mIDid9qISr7739kaDNCRxSxllKPJqPJHaYClsKjKtrP701m4Q6z/1PB2c63kIU6
cTcLUgDpFmr9R1u9UMRmnda31HaOi8SBVmkURLr/Dk/LGi82PfJTsGeKzUn6MVw+fVWSILQXjnEs
dkRAm/9BqKGh7MHKqybs8pIRwNUtTqhjgHQqBt+ghjLdw1OACSmrhOZ56g9tjofngH+QnRkSGy6f
H3duyJo08at/F1v2BK5anPjPhbIwt797MZknX45sZ4T3ASNFGXWc+SIcWfqqIIqqrM2phQgYoj/9
k3/wRR2lH2XE0cJkXLrd5gq9p5VCND0wQBDuCTjoqTgHSmEPhcbH8lOEZ3IPr8BOAagbvx4q325u
7/sEDJFZALrk+aST024YiBOh2AgiHr4sbzgzGyWviau2ST/9wnuBX+BXZw/7h6lVtGB7EgbXcuIP
q0jp3dyqgiVeJjVHXB41YMYLksJ16a27wMJb0LU5lGtrPSWc3Io0nOSk6qPKctXeF/2vk32s3Vl6
vzLaKQKI5xUwet6Zi1I9M6qJ39fE349u5Kl4hz3acDHAbzhLeJCWWR4a/VywQRFAmEiEgq2UYzWa
v9YSCNjaMC3PLBt09qGz8OKbOAdXlUitjNcMUkenv+AX6AXbqIxdixxWBTFcJXinO831PmAdYgFT
C/d/ZBK3+hIfHOc6q+EzCFg94UZg2nofz5SfqG/iEoSVQ7stSC6fP7K5S7GkNFVIG+CiY98n6e7/
VvbRwiX8uK6ztQjLfBHzqp7LOSy4+pZBPvDjH54YRHBtJdRdLUz0eS0jhA8aPoOrnRUJ9aGSOuRA
k+okMC1md0Ckyw+LGE9Gt672w73AF6vkVJJOlbMiTb/4oQYtACQfaCWXbhGhDpav+gkyrKnaXpK/
d2FhSpPGfxlD3A4G0sqb6kMqgcL80gE+kA64scyh/wO80GYaYBQXgsZbAFBMEMkNEH5LLYPe0+0u
TOp7RS1/W3YdFZdopTd9BSY/c4sLHi0JXNTa0/AloN8phKTyNc6IDLtxZwsFxw3rkEjuSC7/LfLe
WfQWpY5flXefxayiVDwnaJBb1CLg1WQzbooVrXP0efolmwL9FhaTJDtWlqcU8LPciHp7WjL2FVGH
zB6HmkY6FuZBpYojpSTX72MSUCh097GqpuNC6VXWX98v5sjJR70oZ3XFyiGDZ0byqJ83Ed3OW802
6v6WG3nxepIGIFm1nUN9D/1QQnJkEqIcZZKpoc9BPfJepXgybeHrAy+VvESw64ADld0KyapfVagv
ycyMQgwrmU7UTXuj9/gXC+EugvyJj+0p5/PsXEw/jk+OuOP63DiSiqSpx6dnCFpc7qPopqp49Aff
Q7NhbKEdUzXYnkeo5ioe9SW8m2PSlaDvs+W0ypxjr3evnlgNHyxeIEq8WSG1UFuKoCwjHOLn3NTQ
TC2Y9pciUVqYKnAnV+QMQAYI8WbdT+DusDqtWi20Aw3hFNCAtSzdqNOkFLLW0jOSPMyNn1acthYO
YV8iw5W34PrHbm/7VHC1kFm/oZoEtpa60ZInHhjjBqykAWMw+RgKWzo24r80rOwQf9ZRe3ehJA84
YDdzLA5CpAFI03NSBKsJ1BNRioTgkaZAk+mVmc9XaoWACkv5ZrEBkf0EitoU6TBp1+Ugrzve53TZ
M22Gg29OOhY9bf6VAaLGAXI4zRZZYqMEz0dUuJwQea6OxTE0H2i1Uy6HXFLz2Ox6PQcgnyBe24Cz
tDqGptWqNYoJN5pioL9Runpb6QGJraExx6PFu+CI07XY67dCnp3O9zfJRWZovgAlGBYgIPsLPlzf
++dB//BtjDU9weZLeqaZsCWVZb4JFsiFmsDP0sd9OpG7fAkxNQgM69ilAGBgt5Q0Ma5bbMgpuOrD
V1G2lwzRyTu1EtNkv+O508JLgIOtxRQvK/F3WBx5yn+ltsxtEvyrbZLsJhjlxPY4n3qDe2JraDX2
sffiVomR1N3pVz6V70jOj+eZPcBRs4f2H1gmvuFRM6yx+1sqTVKDnEi5m4J77gP1uXri107f/T1T
HQ1NdJaMjslz7OqmZ5vEMVVkdUvzwATRTUL/Y9VjC9ucALBWd12FmeVCQjdK/zsOdg19xtNh/+A4
ce+GnyHvRugNFWPZelWL3ySmX/PGxAAd6lfKlQj8YaxUxkUQ5WqXQqUd6QHjzGcEaZBkNiGYsfbi
zcri7XvsV4qpUbivQ+YUXpIV5SKT9aSGOmt4HICD9NAw8rZ8m2W+QOdhGacv2f/DteVfa0btGywg
XMKfafh1hDC3hRZEqEGEI0k9aj+Ebdu410cuQjbZgl/+v71JbJ4Q01M+GY7boNtOLnyyR6GnDCsO
eZk8hK9Bgl4J3gS1gAJmwEq0oxQLiyRCZI/6je5nZcy/trEPx3XEkNRmjMXy5dog3/95jGODG8hd
C+SgGKWmUOSo13Yryqc35VeKS+oKVrzWGqnksJntOiRzuEJNBZrx/xm5gF7twP3G5Nx5R3wia0Z7
WF9gs1VmNQonVspYraq76s2KezD/6DH6Uh+U3oTuCghRjEbYKwnFHrH/pGPDBVZgtDu8u2Ccwxw4
/fGJAOSemSAgvBJo5TxTrj4t0VeEY3P1Yfj3Sn7pOL6EB23Lvdc5SKcF2kaAz7/AMmqSIvGM+lSI
ZS1d/rqk2OaVxA6ErNUTEL7Be6+W756okjaRostdpcl4c75gJQSWIfUmBmQwdE+iPOB2rpT3qg9T
3aCFa0TOD8w9pm8nizIiskphKJTJAVAnnR1F8Kco97sEXhVUBil0326E2tscWJVRU154giLIdtVz
9T7f3exyc3AfkrQ3WhYWlmaOKfoSXQE7dUjAeLbvO8jS2gaOQPXPOMzwRTDJ7XRVqHcpFTKPG+h+
ZtlcP6sbmDU8ejxy/3BII6GXaZwOdu9Ens4TTCoWBJSnel4w8rAMRKjfLs5HNmL6Ap5p4y2hcovd
HeAXcP0FOmknyrMrRDLmLaJtf2ZXBwpJqjMZ83RC2xt0+i1iD7nUdV/gz67Tn/d+58kjAlNjwwq8
BrNfuFbmDJvFT8XxdeJlDZtpQ+pMZfARvwnZZpr2V+ey/E6c+7JnTTw1vbNUu4YhxijF4851SL6U
x1Yy8mOUAkFfLjkVnqs2hG/7d7DZ+mbM0E/qMcF6/UVZVANN4WrzwHDhg0NYbqdMarP4+sReQnTc
KTgcZxPVw5uw310naP1JTJUE1nxJbW0DP25AX/OTCYX50RdpgnYxJUqsBkeijwViChRla1Z0WyZq
l2vecAqRkJWCITpe0iZpjly5UYcrsgVrSq0juWT5L7jh6TUwfCgQbnGaj/tkshrKzkAg8wiPkkdE
WSWPza4Eg72ebH4l0bk9SMQjfSXiL2qxV+71KXH6E8fFvJYhITRoHjiqmniwlqhFTtsqDFnyCOZj
IcfKAu5dOGppgdQ8oDVJ509yoheaXipSed/QXplgFnKIveD/mpSEN1uJDmEq8yke8z9MMXlt1U/g
9gvA045IBMrNBzAbCZzZyzvSrMyBA89oVf200WmQXmEPIDmxnEHeBaSv84/pi+F5YG2uRcE1Iu9J
wItcIb5uj5k+gH54oE3SZ2bYbsq0Et6gyWbuqNIIEjuEn/6LUIpA0j1ronbSMl44vxE1MD6+r8AY
DBk7MzNMZVoP/fK51YdXWBS6NtB6yQyxxC27nbBXUCbMrdhWjcjVAscIeLXr8h9pMzMXsAI52Q5b
+YTN/6mutESWj1NyNYjfpY2V/7U4T3NU0UGIuiUGYkxKL72yFlcPV7us2zbRN/BEv8JxkMycY9hx
KBQ5X7LlAxiEccHcSBAYNOYm8LHX/MEt6vUc6UWycHPi9aEIPAL5Sf/lR5Vh+9rEJksHY3fxXmJw
EWVF5X2rEacGf/dSujLWe/nQJKhT/0XBi6cBE4FNB3E2HtOr8hnCGRlUc8L0Oot7Mdyyt/VFwVwl
g/oRMeilYEqOCWfl8RRnw7kWwstSCTD02Ad0GBvuo3kF2GED2din6YeiOg1qkBABFbVgRetX10iU
+26Cd37TA4vYKnP0ArDfC/+5FcOSNWGW2tIaYVVQltdNnApQRY/msV2V57lVtaRJpejRnScAFGti
MG+5rdLSYXhKY1+V1TpKXKAxqMeyeK8D3xxPWWDrhtFdh6VBEQhVP7bndnxYFajp9FU9S7hcMyGM
CRgKmflRX/rPEqYtJ2D4d2Y5CEPslsXzB+Bx0b3r7sfUWoqIR73F2wJ9y82nGvKXsAo5jKdT2aR2
kPCAiZbhXenlRyq1GUwGu+9o+LEEgxCa1tY/I42SrwzAvVooD/HzfWFAeaiUO1YKc+j3sALlFj2t
AMvGAUDkuDeZ1tko9TpGE0IIe4/lZE0b8yvwJFTErTTTUFeFL0g6E3acTNVQhsFHV5o7v9EwMDVE
Hed63/0SbOKbJ80lnvgI8Re4g4ZBgOHFrejivb8/+9PI2wgQ0T/tapeyCqVvK2MRG2qswObqSAzt
MI9ggN7XETrbD0EJWpcxLDjfeK9rryUZVjSb0B4RCtxaMAdmupfuAgrZpuHoBp6gBjZfPiGt3Xlp
nTWap6BfdyrNNi8KYgGaboW//rBoXzG2d8fZ3An/O9WSAwFEp2Z4Yds6FXriit7eQZ1CfmKdBIE5
5aOCplM75jhc8i8dsYHQl6UW1v3xfnVDWg5J6HegLz+3/wWXeDBGzXvDAZpR1LL2sFUlRjKdQ8We
WZPOm9iEJBocNUKtllpMPTj8kfBRigQqaQhPo1NDCYUbLHJ0FyiXn/Rvx3AJIr+6Kl2vS/cSznIp
xvGpL3D2BHTTADftiKJwRAIwCwBRl1hFcA7IbYqlbqBKqJOhbqK0Hl/QFQXCKoUJheTG06PTdlN5
m5+bzgbH0JhihxGeiz+TL9ZHs8/h4GEA11mkIRpFS7vXy7oF+VaYfLKu2ZcM3rlg4uwvqbrwFBoN
XvS+MoNvTEAL3zBJi61U0XFprjS3PZIxCQTPm7xSTep+LriS5sTO3XDAkDZYBY9fbeJcyF11P9EH
e29jVlMNJ1lW0xyFjxauAPMrq4tbFhGM3TP9XdNvMZ9QET+MrH9NlnYLVOFAXEzLT9QWwVNKEc2B
pCD+K3I+IN82iGKSbgmyxQ89wi5DPqorXoNJUh4W+aDZusvSYXOAIy3AEv51NhdrgyKGixC315u8
jS1e8eLO9X/yRVS/AEc4GiZWzBNoH+fWh9FTa36/2LhnSUflGS2GMm5cuPjUOj9p3gPflJK49KFs
4A0JSOF1A97ANDbZrIXo7QenffG16ULusa95l4cuBsoVs/kK6V5FtT1CMLDgk3RgMFShKPRAYYn9
en6IxgdlizjZTUFF8KnKCJOCgiogKC5jLgdjl2pT+nq4hzwaMvsNGL4hyyqGm/CTHXDUcegRogtv
U/smSWLquLbvAs3vk2wCFPcokqtAlhdz2fdFyXznTB9fji59PULgH6id8YXyqa6D+7PcQG8Kt7Q1
hb1YxnCKj5NRq/vMbLIG0xzJvrC1hx4hsDnAHWGyvo01jUHnzMy9N7p6WYVBesdhc2q8XNHELMWc
3wjVTTxbAj2nRCKvqLFVksPbB6G8u3GSdB5tnhn4whNWbA6k4kNVi9IzrJwTQnOEEwq8xOzLd8dw
55p0QtyyIruL01iOMTIr7VTKowawD/w33UPGF2NGrTv3LN0uRZf4qGsTO2gEfsjh7PnpNG4rE/pZ
G/QNmqck3Tb4uCLtLCV5tq69UI06xbIGPbzmJJVvPbv2H8frp/Am45xWiHCQ7xeWLLmsUa4iDVFj
CdpsHa+BnAF/bqLOO2zPj65YXun+qKUEnG5PF+v/TFVVfC8/cs2Zab0l1JU0db0EKjIeCPDvlj4B
6YWp0xY/LN4ox2O5N5peZQ3cOUunOs4R5xmJzbQ6pgEzzEgtyHfop9xftP6MSmeA+r5Kjsq09gr4
5QHWS//bdEv/xBNbLLhvHJ3AypQKAVYBSoE20xfpMYvbKUdgknnCvX2v2Qu4eiZ+zpvHBU1nP2LF
4IJnTFluNbUqqRFXf7MxW4CLQFHBgNfznBGT7v7iZLiBX0EB2qDnA9uOVywUWp5Rkmnil4SNusTS
1h2oph2b4odIRrakJPh+7t6h3Hsac1AjbI5WUtJRFTiqszTKJjpOv7xS1DfKIV8Lkrttg7u/C5cm
J6WI5m/urysEEMlvLCXUByZKNNxhegSeEFzeDvSiVva5+xYIjOrxL3IkICXaRMITsVwdfhLRm7H5
DhD67aNwbE/bnY+y8QQve/us9cIwhMgTGlNwOVeM9O3vbq0/E8YzFv/LwhsQuMegYNH5BnWSGWu4
bKVDeAwJhLnnxf2n/MTAcBhCHH2LpdTVnGF4nhtDx6dFCXbs1Bk2o144NmkF7ATR2JPPkmR3x8Qg
U5epz+xa3OJ5IVtpXvS1ImmforqnEpRjNxwKxoYb9lxtXlIXtOW2U+9B8vUwz3AoxEX0deXFYFls
MDd0u08uCsE55QugPPBnEQPKBMHsczdDT5MrKXE59I5BP1IinexCYKmb+I+zuArIQGJMVFzynqSl
DiQgjeAaSyEtA7qzsRnlqaClNkU6evGOkwJFC5pouG5DDq1nHJvYHquF+ZNvzZ0Km1qdiTrlgiQt
pKeM+xUho92eblfGRGDCs/JntcmL6o7WeLf23E+7fOLmctcdvz4CVI5X8q7P3XrxxMMQ05qSqtyR
e0lj5NavCpUhWhGZu6kbCDwnQZ+Y5QWeL1bjf8/DcFI92br1tl0kYMOV8TQmodVjRpfRUsfWv+nf
NSJnNqVtuAwMdkdkbYV9w4fPey7lvxHc+pBQr2n8RNqtxOrd6Xx0XAF1UKFYLO6mq8i0jFT4VES2
fiSPnAuAjlwhbpWXrS2Ad+R8jyz2Hi/DfI0adYUcbNtPVQlZAoW3oTe7YGCWMeWnjlaByKedGxdL
zodmhz/7tJ7+KXXzZFbea0fesuHf+2HVLxhfW+KD9DeugEo9i6bDRMjgz/mufBO0Ulvijzuo7DRT
L5zfbgTLLkBJndsrDrZnEQTaMB/fAogvAvqnBJQI1u/OklBbuXS29PDL/bxfcXCZgwftjG8o6kFL
VA8QQyA9EPHvMbb2WCFJJHEuo/jzEqtkv86fEtNZr2Sc36oNXcFoVrTr9Qtg+L141v85Te64IAJl
FkVW+xt4p5C+RwikcRx+dKawNZ6yX6jw0wvtGz3QlJvUqYg38PrDJEHLAP4o5yt8MwWm3LnhYta7
rOI2fiMCxZqUtyOnMa0LU/IfNpov6kUMfeS3LWBjWx6U5txyWxJ3WLXY6Qe8FqLK9l22YR9eJi/F
V2HiHu2huv3+ACJlWkn/SOnrcsMdQtgQQ0BfXuHpE7Pzkx93ONozEQEOy3FwtIHa5pIKpenS74KB
pXHNySMvSzojnjHz+T4nxYd1aSoKwP1NLVMDl7OnAbBxi2U+DxQ8GUZmWZcw2JFLQYrOUQ7yx2/n
7l2b1RRmPS+DSWnxNo2vXXYOCD3YLWFF5yCZJwjC9MGXcC702N7eGwdWm/tNdH9LCg7x7iOzKDb6
aVAg6AgxJld9/IGy1/96Y5ZbjgvhjUhOfnCN72PipwACBsWOg8ZDs+0Nltayix6Jr78mVNdECYhr
lShRRV7E+a8F+bGQbk20QV46IooeNGbezzhxLj3eGua3GyetS+TjwkJ6D9zN2UtEmmtdLoW5ihaI
jTSgoW5mWbQ4VYBjV7W4fB8auMJ45yAejNVZzkZEfqfMgkjonT6i9mfbZWxaAtpOGHabAmYNHby+
9t00QK/D5LZM8vrTXg1QWqub2VSGFMIbp6iepUOgMk39pNrlO8LqPaU4toTRkKu8LI1Cy86sEgNP
gUTBFJwdXoUBz5wY60QkEjPYhNi41cA/7hi4ukrIHeEqC13FO2T8ISe/AwYFieyLUks1MlZBYmly
fX2lTnI1TLKns+oZjdoEtznETg+cjLKvO+OnPFYHs82/vQUIDLBS3agOvyUM/QG9bIEa9AZEZHI9
8CIPeSrbdJ+I38eC5yeoIxgZmyh9Qsqa+ZqWXSImU9tmd0Zsjgr0F3gO1GQjDuV6LDHVohv5OAEb
7sZLejSdGA2AoPfGSSIoni1StqGYABkf9WIXjAHQ+onxD78ijDaQBfBpnRFskgoxAUa9vYTDllnk
LkYLWNhyrQQ4grzkYzLQIVqrJybXbs4H4lAIQTzsrAqyexVs/+aqAlBkQjEEWGXpTDP5IWayHHv2
ZMeop6BWL7CVSNqtbKXCfaZrpufzfR4fJvkHdOk+QFI+Nt7uVnENDTIsG3sT907k3VkHfImHOV4K
GxJ8PkCTVMNl+CkGEieNS5VyodzVgyUlxUKKm+z81vyqsE9pmGprDf2epkffAtbFYdPjjFCopD/T
e23n9vFVE0DUY03LG8sIxbDhz2ifQVhFFnLsl0Wd7EhZ2yEODRFpLswKHt49A/1FyWYwCOPVE41h
gOYWsDlv6AexvuSU8+8PjpLsdO9XaX0W31Us4tWKZ52ZlVisWOBgixBKrWFvVNx0/m37iUABZW+r
gcvRFf4Rv8M8T2bsqHjpUCM2enSr0ichgUp53Oh54gyFq0CCRfFAhKkgHtl/f/sSq9zU1B74r48i
TrKvDeIP2UpVNZu3Xe3gPQ0STSbN4gN488+oELu7yqJDxk9bgkeBwdJGyFC1X0FqCjvONK6VqZxW
i1SQ7pgKvuZno5hK8ScsodWyQBal+G+vkuYWa2NnZ+AmmRhxzKj9iQL+bNby/4WlCeWzLRshDBOk
4wbadQ2fYsVeWjIc+wwjetoGJix4KcEb9lrlJYDf1ptBlY7w4SOw4+RFaf9gC1F8giLokqka05xF
X64WVuRyxle7rUdyrW/7/i43ivEnBAFbUEGrUFaqR2EWuJlzHjuvSQmJyeVLhATqQZ9ajEdPLDLi
hg3bcrWkslb2k7vXaqB1vMEyEZCU40syGnAgIfElKf3An/MzGVr6LZqLi9fI1Q0iymMCHPG7/Vrh
Ci8zu1J+O/s8kMbUkN1bcSJCBAH5/qyxjBklqgD3FmuiaKf3gG7nmIIGnYeBQfhE4wilhBDHpw/D
Ko8vJa8O3LUPpX/QikMBbiLlesi4017Mu36Jd8HZ8Ohvc989Dl/hR7R6d7+y+rHQDS1D2S1Otj+w
u3c0ftCoef3BV1EZW3/eZ9UqgZTXxUn8H4xXkBkSeiG5xMjmYKFCRYJiU67vUE/XeTpSpYydXYdC
xCpHsu4ZSAE9YYCpfA7fx9iUe2JKoeRcwIw3itRg7kRxkZfCPxzxcs3cRfoNY0yknqGxrrTYbEfR
3Yr/EfrWJ/lwCKxYBlS3IxyeOW3gKQrHuiRipqgKKl0/WLRzLoJJty9F7oiHRc4gOobH5SXJHAvM
R/5n7oJLGj86oC9/7GYTx3hbq0bZ4RAuwQ0+zIREVnlkqUXaVRrA209wCtQKXibe5mNkT+MgQ56r
fomWZiqAxyeNaQUmW0gee/+Ae+ZaUtNPsryFR7ctl4ShJH5ClK9cIpw3ARMiV7ET8JPuKLNtYpqR
U48SQ+2pOZ4crEK/9g5vS9laLE+bplRyOvY0jx8gv9DlrkLWJ7IqyBiigf2hKDBk3B5j6trMI4c2
6by4Cm722Y+oqTWYmcEGomUXJtOa/5NtL7aLew6JTHb8OOTYJNSyVQVPWNbTl8xSJzzZO7+f7HFe
tDALSxGt5pXnDsF5WauRbZbc9zj+yKY+pJfuFTTN9NqXgyTNF7JO9EoViq9ZAmL9aQPJA7CoS+hM
be4n6QBd2qD5oVRl2o1693tje01mGZfgazCshkl3E6Bn62HFj1MiCIwfvI7FFgH2F6gFWx81MAIW
8qJVgDnnjRi46l420DRAF0a88S0rZO1Pq1s96jRgaW7Nkeayq1HW1uo3kWy1YxGEuMRXVnWAy8G3
QwXDjHOySm4UmVHVT7hzvtdurCNLeI1Vpgq0U1S/IzqCPt2KX12vE7N3XWJC8Jz5uHJ9AEy2jbJh
UWmpy4d148g5X2H49RdkSjewa6iTWuIf4wdn59j58EsDsD53wTLFdUaO+Zn381qWJgfS003vsbYz
w/4t1qFnRdjnxNqdL1QWwnxGoj/3LvOaksZCKQ42PlCVROymUVBOlRleoqMsWXXheM9Tn2peUsJz
6P4Dj7UyFfiFVF7zXXgVQkLHwzm4sr1xzjmoEwT1R85dkqfQSGWUdD1IQPEt3IJZqQl28V9gJNMT
IMVPT85MB8w/jbwUCPw1LDZKgTBHsFD5H+73Yy7Bbbc/+4QY5P3Nlw6HZ8ER3s66Zjlwz1ZDui63
eFgbg720O5Hqge05hdZ0/YMFsy4fOS6w2COCddkWFe2fCC9mV7dGc7m4SSV1MoH6dL6JsmuNu0bm
1Nntwa8RRTclHysdgqF9oGC0RJYqdDD3kzS5WpjvIAso0/MbU8A2FSLsTSkZ/X7sd6vjHrAZvT1q
yIpDvSHMhnyfSIbmc4gw+GkVbLe5QEYYiTLiObeD5tNOHzKE0ZLTXA1Slke482+pjdVqJli4eutp
BgIprq+hBghLLS8a5+J3BNuVS/C+jTeg106gNIvpvj3eTEo2OUAMCx/VPn+9TtwJPTyenPWapVtI
lAQlTY8jvxo4e84NVwPIh6pIyWszSEMUmk+p93KsxnJsSeKvqdrvL9MVyeN0/gw6M3AsLJPnP4Wl
eAJtqkaOyvRv1N6CrvUNiXjZMyCkv/u4al6/I/iYohCzC2XxtkVWr/0y8h3GvVEycaHwiTXNeQJt
9ar2M5MdbnwlUAMgG4QbC37SoXyn0u53oPb7FkC0v/NRPs+QP6ccf8bxhgejrnIY5rk6neDy8gsT
hptDw/z5FybW7VJ/jsLFqetBfcpKaKqdpi1S7ojdZStCYDQIJe5L4sUZSXmzS0aAVwmMTnLXAUqk
YD65YTLNjZIZH8zf8qfM++lgSbF4/j7sy+lziiYtnYn2Ii4QvMfCQzYnhhwCP7sawxotnShOg9Dk
RrzDx7F3fiH97jqGean8Nr11//BYNrmXLGPEooakKEsoYeeytRU5+faoOKevUT4whuqMEpCA8baO
n1+eMQH6J2A8knws8wvZi0uTDOL95E2THbuZhfmuQ09kCbv0K6zgz4AN61hxBphshSOmKQfHvjWN
RNbfyc6aBDM25MksMQn+OmjWtPTNTX3yTOleBz7bn2Lz6NHtxIIFcBBjjqJlLbvPw0+pTEovVSWX
B9xqC80DRqS63mIN3RSEf4TfvWXb3iP362oAYU+miWm5FXWMA8gAjw7RX9kHjmc3sKfYg9GV5VRg
PU9xPjjWqMhcCgP/JTX4zQho54yfcXDfi5Db7dIspj9buuiwLCyFyrZqV7/LrjBrFbVkZsoVUaif
AbqlhAliUadTfsyk1xfAD2tnGOjjYcMVl5stcHt+Q+Wj93rv5XGoCzaDcVQ3xvkxhQ7TajUyhtvt
yBQVFT9SAPdw0hO6H3YmuJt6Jz46ael24VSQUTO0IOPhnVeNZe+it4GmtellU6iFDrkL8FElJQpv
5MzVnGYAjCkT/ylmEBWtKwB/mXA5QtKUB2Ki3Jr67bsu2OwfJyAHKEarH4y1ALXtgrp6eFiptLzw
qYNL+GMIHRA5rDPwaL1dzs6rlEKc4Lrb3pVvWG9ub/BSmYkUTmwT1KIZYD/0uSIpD1+ky/0/hHVR
ySz/yVNcdbXJfKQQtO62tNO0hE8fcB3XdPBHAezXkaB8edAT40KBpc6a3wokJtKVaT9NXDywlMOm
Lj9JlT6Fhs2ZrUbkMSMK3wSPAP57pGM2iRX2YEoWxvu/om0nfqULWoMwr8ejdBRRPfM7m2sdbsxK
eSus6UaSHy3JQk8nkjp68bMNYj0+KEsJjhlaqo0zcQqVfeDiHT0oIKaDQEKTfnaI191Zcwz5mqtR
CgH2Ij48r8rJORgs6BaFiHaWn5pRvGK03phhEjoIjBkMCCKTyOBZu00mixeKYXS4+wDVjtcDw66s
Gn/mRwEOMH3e5olAty9EiTgNcpasQutn5AXrXOs2fzzqwniBbxm8Zpr3tPM5YvnB9xGavON7Wu1q
ZhxpvdPt2dh4+Ry+LOgG0CywhK/pe+MFxAoHNTnNBEzHkUz4iHiEtI9B/oFFRC4+rkpzPm9Jiee5
kvE7nP8lbzITzdLZK4LRLrVAofJlwNCvvMjh4ELKWJV7uY8VmgQiUV2GSjs9bxgL/KtG4cMF08y3
fUm+B/IuvJCHTBW3ttD6V2uXbYvxkmD2CKUZqJr0j9mSuCuKkdG3r9gkfVfA+72Lu583il2nQ/W2
zds2sDS7BjfJgnSA5pnhu9JRd4lAWCKqkG5RnryHbdnKXEVEmGE+9zfjbDsOZtymIxPFCasKodhm
UWC0qK3XeOvx7Jsz6lp8ppakqqPs7F1WgZ/Of+Qnae3XVYeQ8otuwMNiWYHHirnrU/IQNHMTVUXh
Ao0sE8l3IQgwekdNAeJjfmZbmUtIErrth+oC5fvTKzjSmZ+BN4y0RF/KDO3BfoMarXuhJpfHRkz8
9XT+az3f1MPYkjY4bd7zd+s7lVRcC5B9BHsKG4HYyoULSJhQzmmiw302rgnDeg+mz/lzcY3wFUZ3
z1iVaBVeRe5txmc/F7mhb8fs7APISv7Sagyw9d9LGkVAlHqxW/CRorGemvaRd/oQlxswl7S96hHv
64lELPj0ysvPOgOR9NIDcdetlnOaOirMn08WeRXmabkTwGSxLnKaCcmm6ukC5mURauB+XagT8Dzx
gdSoN+9LWet3ZoSpPE/7Pa9GJyjjiM/ddEYGl0NXlHwQ874CoYwIpYVaUitZL+PQW9L9EaMJEJ8Z
yXljA5BD6rurWGV6e4vuOQZIWUrOWHM5SFgKcR7u+pYlJ7JPq77EF5XIONUfIHJE+IyH4SkwRqJ9
gjok78p5aLBl1rEdD740TGnT8Arw4KAQQWLQ7qrhtqhEL5Wk+I3hZUeOmTC+mOPowrJ8aMt0qu7y
DqVKqGLsZM2oqLgZSt0IhU/JAhJ3pcqlrMzlJkSmwCN7NEpVGV6jD9Pl8z9epGsg1epf6oRPyV20
AIfUHRUOPsGX92JtgxId5W3LRP6seHQgkdU+knNqhpNyk30URlXdtaS3PM4NotZ4jdGcwruw2GOb
raDMa0SyVun/KTZ+kiwzLs0+3B3YcFgFpxpkoNGYLC022PtVVsMkoDttQlis7PktMc1a0tELWh1T
516AYDWelYMBze8xOPack2LV4WUH9BD4oTSvHRP/g0sCQg3wj3Ocy/3y/mL8eSepacKclew/+b9m
lUvpJaxEH6Xzh1I9bnEquS24ZPatm/gdIo6c5RMTrjRxnlfpkTQebb57v83Lr699rDuGQLMbSR8c
opH2pk0Og1c8nJW12SdZ2p4QFnfPBvWgSiwok1D/NBYZ6G5HuXU7r6Z6c2dVK0zNAp8fYpi4maAQ
0iTOlSDmJxbF/WauuB0G258qm2nJwECaGB3kK/E83lwTRlFmsYolsl1PhI7qK9jIua9VAB4hHs3w
QE6LKPrITnR6zw7pT4N6KMgLt4wzMNQOemQ5aazemwMNc0bUjFJelGN9aZfYoT5DJcDLFWFLPy4A
lvSh9TYhJdYoCHE/+GH+3MuPg7IuK71wJ3USzQeNNjxzDGGz6Qa71PeONWwc2zwtAviSKBIqSML9
6fAQrdvwli/EyVbm3KXLg3X+Uy9uCwTpdyjHSNIwU4KVzfpUVf0uwb8rA4tmoBEs2GAwwty37gvq
CL8zYzWRPkqB4q7gj+/dfRx/cuJpiErLx4pjET2y9H8BHI7cEsEfOydWoiwTSdW6Hg7HUj+HXc8A
PWfhhV2Tv9ihkCrUZFxsFQjWla3PXq4B9jfOY6yNvo6UOE2WoKq1YtWMeKQToYTk4Dq7BMgHTH3e
ZQY72Q2Oor1/3gaFZxtS+6o+c0CmbTvr0JIoBm64HD5TXnXlvvLDk4hNnGLjMZuvOYuoskQJv49n
yKw8rzGE0NDgRHrikVj0x3/jUDPXhsp49puVxzzAKfPWGT3FV3dz5Ck0eawNiRvOvKpe3+YYgvjI
b3YTxXPIfMyhuaBkE7RXROQ64EsyiRILSZ3Ys2fxmg0fLfkOAlz8sFW88hsb2d8xUyC0WUu4lge9
2iT7HddW5oNCmq+/DmxZmLIrIHnVB9N51CcVm/5Kjw5eDFOpxSSJBdufnGycetFrDVDhs6CO0ozz
7Ag9wn8sd/ZvfwbJNFWLvfwg3fVKxfZLQ5CUnyCbjKzbN/58yV/05Tdk6HHXdwcPctAxcdswAcsS
GH8jNdeAfuLwHEoKNSPuiRfwQ2sSG7Z6ExpnQJmtv2MZylTUMZhOftqc/bMlu5G0SXvRd7iEU2fU
pvlYaOedTmRKCi37Y3SO8kukz1ECcIDg36+DbA0CcDBYolrsS5ziqH1/hvpBGBYSLjzd7UHSEzKr
c/AFQOsEV6FjEwf1OHl/7XL8zoFm9YvQ/OdpBQHwpGpmt+WMXu/SjSdXczFnNwPLjJcbn+f+nY0j
nXAyLCZvCx5DY2yVZrD0dRV1gC21TC3/SfueRs8UHgS/F6xRY8f79i6pH5fDRt/6riNtvA4aBq+i
voP1AVocDYa88eoWHMFJ7YrLRP+ofEhOvzEwt11i08ANPBTZPj+avW8KO91/6EzJywM3nbJYk0UF
69Dve+EL+rR3vh3nvVp6bEQ8vlOlQvgXOu25f8cYk0cVVs2iop4LpSIV/bobZZ0XZLr+iGSuHavm
Mr/U/1sTYP1Pc0lmuubQna9TBkloXvD5IKIdi1YT/HHfs7NaIyEhXLFfUmzQCejvAHSjdc69jnvW
ldrQHBbMnU9B9d6DVTkhSFDRM2MO4msoX2zXG4zNxBaIx1YCqCdLZqVa/08VixEQ8GHo9dj7aLfv
dkL4FoPP8s4YuCjBTEZohpP/Xm9QMuLoJf7GWcjYuYhaLgUTD/x8plXQB+nGici0XdaxJcHj6swX
iXEL+r3i1otWx1MYLPh0i4kQWw+n0quGSgqTL2iQBkqXaTrKE/V8wiDs8NKJaM8B73ycm4X0kCGp
QLIvBpErgD163E4Yeb9M6uSRWWk1iw0N5Bu7uVfu6ILUmH1++SSTOGnyZp9PI11CL/v0O5waxp8h
RrEzDXbHkXMY4/1dTRcizU078oG5nonf4I2fe229/HYO9fsezyoHK6nbCn8KQ+o0+7xYWUeoe//+
qUuB8JV9dVyeIxhlZUdzx7vGL3OuoH7iYfLkRoRbr6frOaVs9ZsqVBWEbFDvScxY/ANMojTPWrC5
FcuTtMtw+63/7tOwbShWwf7EvGk4ea0CIP7iV+lDzwqURGGp8Wx5Tpp6RzYBBYNEjxD1Wu+wOnyW
NFl3wTQXnqjwoNLUowFVXzqRTOQjor1k+l5y7emrXAf5PbgnqDyFEkhNHHyU9dWNzIz1gFv++jnB
8pGcaOTY8kJUE4Gg+f+pb1P70glPBhGBpaygKD4q2bt01JBz1CGdLaMsS2GnizmbywJApnTzLVYV
XzhURQyHC01IncEomYnfm+g19/F7ndHO7o8g884QLq7yVK1Ez2Egb6eZ8E0ArV8jMpvlniFJXc6A
SdqVHyoVd6SelnBWItm0c7hfz57juK+0IRl9AB+sh/nMvemCz7aYGEcwJYcqsf7ZJsEKZQfqDxA9
cF+uQhpX8BHhFy7/YKFwTEM+GaQ0/5q1Ujuk+Jppj5/8wtSfVZlEPv5xQhvI2MwLpSgJNXW1sR09
w58rNSTvfIHQnD5Nk5/yBdqimgczzXpMXxPsrX0G+iZ89N9p9/t7iEbhBJPCwOxlsrFweSQXeIUh
YH8LN3M0mGidCEve7EeGrN7EyJhDtUXXerW/7XA0MtLSkJXB4mT7C+It9FS9jfSbPlBtOcqdPkkV
X6z9i8VrOjGdPTOH3cX7o2oiSMhCc7jbCRh76YdpLLBSRNd7R4tLUdDx82Jiwqldf9NUnvOG2pYF
pu9Pv2pr5sTHDcuh5iHdNVJrn29epIKEviMAtkXAII4yK/i1MwmoSev869QVzFgDAV43SVn+qBXT
oICJ/ET9i/MA7C4nQgN/ow2e8PuGcVO9U+i9ENDmMTQg9qDn1+EDEnYBbHi3B5v1ENtBHatSSUf9
FqJ5pQ9sbzgAOk9jQY6+8MTpa0NVmmahFpUF1nA2UF2ACO3pqRMVxrxWGC7WD7bfUlf5H//w1Ahr
7DQxNvAkVV6yVv1jIatD05bZoWfF5dCl9eAAIxDzbuSe4NCLzCKTy2XPtqsK8Gcb6wZbPdpvKDiN
QRWRRX2mt7UIDhjpVpofhH0Q4fbHL+bpvM7ZeftQllftE47o6p3We8vdFA+yXmEk38eIG+ZseGs/
QH1wHTAtam0fhsIvHZui4nVK7lBAKW5bswwe10DWY7bDOtEvJPouCFg0LBh2dSHvGTuT69xzh6R8
k6hKup6m6KE0zPjnJhuOhH/sSjLKTg6bdh65UF5/Uc8xdKlcQiISa08tksQYC+cxaVH3OOTT9mXj
03eK9yPaIVk2FFYpuN9fe7rDG40AYhCb0xtcLqEqXkUO7Dnhb4h0exERodJL6AQcSIDk3NTG3YLZ
BzvpJsymCzcM+YoRtdmIy8K31GlMMHphm8gMwlQmEV4OS/V+b3Rud580Zdqf5M773Zc8brvK3JcC
xyf3BUGc6QEQNiqstdt4QAxJCNAEKvhEPwVmIuIt+BiLYIwapbe42/UKaSHKIHk4jDBkDhk2M45p
eKLZ/DZqImIJDJrmDne8VojtY8Q9XKyGHDQeuq+6f0nLou9sez4+n8zHkN47mc7UVc5Wb7F6B7mr
qrc7h19CqpEXJCz01tsYrxAohET+zUSKcnZUiKQWzjYdAcPbp83mr890T/MpyVDkyREv1guBfFaT
XdOhUQOAdtlcuevdd+Qoj7HyPdL0vNhwnopzWKmJ5np9IGZHTu00FUFx/TW39ebE1J1AZmYCpa2c
89OzEulh3PUkLb6KXMl70N/FfsF8It+HWAW5BvM4RNH0Xse1fij3jipY34X23HSwVIROnZiJZXNa
9IXYpjyCuQH+s0gl7Y0c65qECWbirwrQJJQYC5NLM61pTD8yzxUyc2wKGRlGrcVf94XxSk6PsUKo
4FmsXZCsqYXAXzS+fji1n/S2OmJh6+YWfqH8bUGKGjOgsgsnZxzBgrPTTTdfv6Bg+gwW8IwMEUyC
uzVYblhe5yEMmzzKerL0HWUfU/+HU9h8aqIM2tlMIirFRGqLVWxADNq2g5ddIFCXaElyd5Ypce4S
4Ma83M52hwmkYCnahZku1zuOZgdWE7swrvXBTBQTavmuukGJJ51wUzgvBZ6PRHQ1mlBX1yOzfR+o
CI8tdEfH7CO32Xk+xMwntysBedAXEBrgx+IJvb8kTYp3RjSIsTOfHxMth8iYtc+T84UHoDZAf6NW
Vr2SUoH6o++bNvgqJO95ozLxDiQlzc8G269RdpoAI3vee5vdLQ/9QHQH8T5rhpomErK+TF68cN5a
pKwdDA7+Af0Y7vrlYVzrMtfZMkcR1nlfJ0WOjGvHwRgx60C9MiSWVUQqM/p7tucMGcuuFfLCRqf6
nW7JOAY3TkztsOlVLyPlP7WhXMeTx3XO40u0wS7Jlb0kSjvhImwuvUV6R7neXgv0/nh21c4kgZ3Y
KttaY9neqRxUbVZ6OsnkWHAlQFJbmbhYbBDwkpEtt4S5DT6t6orNJsDEhbZ0c3kOW+QpFsnGM8sa
zF4v5duEwCTNjU+goMxum6FPJis4NbcozOTTeebfPeXa33Ji/oKU9hBObu1fBwhnucpuc+MfT2Pr
RvKiJron5kFgGweWb/mzlbs6iZhup8Mm1TdFkw2W4fslSq3FxSitditu7Dze9zrBZgoKEAvXTqyk
Diy61eEWIM1V1wH/0koLbBvjiRNqhwQFoBwzGTVpZM2mTUdOYsn5Btir6araZNy7CZX7s+K0HwL5
Nm+c8FKXSRyWJ0m5slFl+YnGeJ/Pouz1z6xK9S7Wn0JYyH5lgJq3fbg/XJY79YdV6Ji4LXngr1K5
CUhZRaPlMrmf5LXMeQ6cQOPwQreSOupZfnNThu2la+csAEVqLdf3B91f28y+nDZRmgh7Mc7w0A/j
Vvu9ciBicshH+QbwP6rpNWecfUCcJ0sNxa2j60YZY6jDBCYMvD514oSKgc+q6Jnmh8AFbjGaE6VQ
BhwEprGES0Bsd8+8oMGBmkH3+pxS3pi8anprKQqcXUKeVpJlv33NREQcPZuf3D9+wLF1WBCoJbOa
5jaroH7dcmybKq275PQ2YsGrFSYLH/IfvZLTlsKzHaGBXVBHpD5OaW5Xd0Nm1eXH/7NF5qb19w6m
vj0ofTZdPzVSMofhVZX1cEPeF31ROWCl8YkNt7FmAHu6EaLF2jUHk2ujQdgkLbJZ6JhsEpENd6pk
SQmXZYRHVADLolUhuELck+rlhF+gONQ1B71gdZ3/wE5zVSQTwUItuNOei065H/ltKw9XDuWy87uQ
1hP2btEH79dWCGD/s2I1KG5ush8V2DtBMdFPQW+bpSzh8rqTXnEtUpkTZ4OTEUde4K4k4rqxXOqO
EhPs9aeMB4GEQTRBjS1Fu1rYGgi/apg1bjquaIPzFjQA2c4G56y5q6dSrAdyq6Ij5FCZBTlko75m
lkxXmxg/uEq+Aq6g8bc437BZQ5nFlQS5tBwTIDt+buGZKt/kRPY3l6Mc4Rx7pvtOwqfCMK5Ttw3m
xLv8kmj1vqsOj1n/sZ93OLbkqH0ufu63XNZUBW42OXbSGlazRiEoSC6AZR2VtTaJSHk2J57kwamg
SkQMAppcM0OXW7WTsLZhQ+iCGCAVq5zPaDsrRglhhZrXgRt5Em7vCCNpBf7sww+UZmUUYy56IPNx
OluZi+3VzK8y7mGmraYR8i+UZwYgBYFqslxlSp3aQLK6bnv2wjzop0E1yvJgbIgJOaljJK0Ld2fN
dGVJsVsFm3PYn6ttZzDQhoracZQnzSsDeGXm4Wlot0NLZie3VPJmQ3uYqOGnObgLYJXYSzwEV/63
T1nAc0zrIOPlCXS2YOHLZ7uzZ/hDrc26reWqxqq2HSJZGt03d3RYjSoANTsATKzKJz5Vdjq9W8YH
OreRQvDklKe6tIt0o8HYC45TmcvDA45SqRVpOCp8eIN5L7NpMlYnoVAIe6EEt2KN0wgeWzaYQKB/
BQOI8jP649Y9nyA/qUr7S6DinOhHJ7hc3KZD1h1PoTY1XUmnj28Z1c+wtdH2RRDbHtyBlyD4OKS9
/jI8zimin00T+epRgi8l/W6AXWIinHZo68CwxnkjA+5ZYtol9kfDzFk02kCP+y6hJTEpivOswIBK
I4GE6UFuZUctPazJbT2O9m5PP8SJlXSNp1tWvxvbCFXd+I0j3ZKapFONoXn3hsO87S1WiWIN8Q9X
z5xzpZDtNKgcg3TObr73TTUS0iJBSE1AUGMk2no8qPFtXp4ohA+KHrNCAz9Z4vlFNFSWzdND2wxL
M8MkljwXm0gXXSy5VkiEji6MaSy6idZezdVeCclCoNHatGqOry0cZJoGzsVPKSIMOrxmdIuG3PTE
i0tXqdvH9Gj4h5PP4MZ4M7SbZCYslScMBgfN3ro1vh5q3m1jZBciJLybPoX3bKrJlN6mF/V/hQBH
DI2QVEEP3VZ1n1P863RCl3AOixMQMVQzZXK3xPczvDpTVHaWayJfTjMFvmpvW7Zzi1CGrVuCyqGj
3l4yl4SSS2B3FcJEEppy43RP753UrZCiJGfl4dmnvAD/XhLscMfYB6wAc0hoYcx1UN71vBGjrZYB
/M5kL/DSNirTbBy6DsYoVov9CpOVB0idCS6VE3hHkvPJuo9f8L4jTOXpcG9ym/9pE8cFmhvRQJZ3
ou0fndmx80o3bcshn90tgQllb5Rh++qz3/Bz7EHMYBVaIu+mlnFxDrj16fe+stLhfK9986nDkSzR
RulKzmQ4haYmmt4zh6V+dBv45rQtHXsk3BBrKnRdDuwWP4BlGgy6mbaTkyrilAzvAf4lmAFIoivZ
HSjQiREvTtkkKW3cF5dURP2++wf5sedJ93XoTSkV0+dXu++kJgB2xXsbAcEmAIjOUaDLhe1S8xaO
qom4r8jXUOu20A4YH8TZpkulm4Ka3lHvFYEK/7wmwWs8KJ/LKXHXEZCYVkIFAO85D8J+97kFViXT
NhFMGgJpMEQqoTzQUI45Dt2NbOlUU9iWO82W3iMarS+/DjlwnaZNPFuhmvTajhANRlWI+TBX+aI3
te91WWm4PLV/+3HTMxFfJv1HUlwG3P4jctNs4+ymRpj22f+OWu9BhS3T37nD3g5HBma+zxxb0LWD
piAwWS/ZOKMjUiBTJyBd1cW1svfjdnaA2gRbR4bhVTA2kMmnectsiXlogA/sLeGjyUdkp26fqjmr
hiyu4jj3SK5xm2MUlDZEQ3HezLTXhyZCsv4vG852qiExE4qMQs0sZvqY6JzRG88xunU0SvNGfGcU
XR8bTBsfq0lZGPhjlIkKrSQDKv8jP8WDJzrq96S9W3aCoxHECrSWFG5tdw8VinTE6P+FMtTNbuiD
09hO2gtW7x/AiKFz/6x7jpdNjp+eWruWy5xNmCNUjpvQByymKiySAZtw3HWLKHH/+zuslfWuIbfR
Fl4FoHwMaTxfg/hagaYbCALsDjSi4914SsFoVdyRUd+4VxdLi28cMh+0Cv/uD0XSCbPlk2OQiLus
a5XYYy4L2+q/PpaqvKOmRvpSRa2m2mqhZGFsVFftF01zjaAVw+KEz7txaVCjEYhBzVyK3epbHDZj
/0Wdg3e0KfZhzqahtoymKIG5B1Hgp9GE3X5HlYhYnPEkcDp5qF5NhL/hDF1nqYtEMAWmu8d5fqQ4
QAswpUWBsLClvH69UbJsEd/LADcmS8qm/3/ZNTDsH5FTqLx5vfQTQblZpkjyalaCMb5gzzaXSOZn
VDbHvffSxavI3cm9u7d28OMha8L66fUV2jRUrZZ0Zmddr9UcW378If2iE1E6P1nMNlp8p2YGsmb9
aRiRbZdwuyx+88AR5NX7y3dHhlusJ2QVcVCVWZjdSOR9aNDcN+1qHdhaYJ5NZAxEzdMjU3/oymoG
+Ly1uQqtgbWNVUfd7Lea/m4zsBMfmFe9uat4x5aEOQgGfNbpXe+aa2pjW0veyYjC++Pgmmh1qct2
MdosfjD8Ts71HNK3wKpW2jtFGrsPHPK8hBZZO2iTNAKtFeDvtIKZyxs84ABUFl9k/BDEyYbIDH53
q8KqazscSXsV1ObUfcoRtivnQu+PAcfWhrHzYUx6F/rLtZBavjhXFcdXxItoHg8FAYvGPnODRiRH
o8Kzv0NWQicxByUSokTSUcqBBo1DtVz3fK7v1EhJOn4X/kj4azCPpe1cLHDkpcClGR2OE7vteS1O
wMv1zygaBQ+zN5ftNbmyz4tfdjXgqcJDzFElHpxbMcJJbcAlbOEEhizZrl+szPI9tZ66Pi79upPc
h/PNMtQPOZLW1t3qM7uExzkSMEhcLf31CqUluSzM/M9Drulhcrtg7y8huk/mcCCagtfb2i0U+fLP
9Q+XkCyFKc/lz0K/n+adPdSsf9ThpJ16B9zwLftnykPBHyo3NL+fhYYqtJmlGtX3x43J2haMfUpK
xhnJLtmfaVb0yq1Z1+kdPVPbeQBKnzEImuTU5SFdGn09ljFhtnMNpEPMH83+hcQ9rN+SjGzZksVH
02omQfMRd0Txi5EgFuwRUnwgm9FfzP+vG3e8AwW4b2ddwo9UGT9E9xB5J2HFufAG/cxIvBiRhMcV
xRZWHssFNxnZoT1pwfhoNAMhCVUuE+jzFXEFZCf/BUOiqIuKdO7LE7VTJdgHVQ6inYJF+1ixDuWZ
caSRVQg6ZKlqERvGVeYDdw2u2AsfuTS74uZCLM7ycmA80qloA5/R7FoYvIc0wavLN4sjHEB7mQxe
dxpoG4lluS5NSaXh0ORRpdK8rGaMWVt8Y6rgNFs8gu2VpOexe3dr17bnZddnR1NlKOqpt+yVDG7Q
yevrOJd60yktq9J3ddfG6v946lDzKu7NOSGMc5L8u6D87O7t9UZWnU8EfKUQWIfVYAcQ5eAnf5jh
g1rDg6oP6lstP9OTKiGrNHAQ04yLSej94wx+Q0UvbnjTOWrDegofpuEhxZHG6AYOU9ZQF8HmDpYH
LKJUhL4e/xKmJOm+BgX+PJ/LmlcMz8y7GshSEfmQKub9/JB0VDftVJz1aY2brZOFhiE1m7aSlY0o
HtAyHh32aVoxgSqMMULKa8Bw0raX8YMvG6cgcRqv365dISefhUjUV7lzGJJE5gK5nZCVwNd8RG/7
4qB+QmqudtWZEi0dSseQVZqSZcY2DloVJXBSe+heVxPh0s6FgHxJHtBmphPnHLOBmelvrnyXPwQG
bjC0tM/h+oVAn8YFHrYldrEw6C46+ze29ad6bf3nCRo4d49VtVtRjwmbafNsslFjjdTYCfMAKU2Z
LzR5+TLk8TIIb0NdojjBbjNRZqGzuGsLxnExMw8CeX0GuKzRL5PIPDbOu6a8Il/Yahnj03fVLLFJ
+jkS4z/B0MsER1aLkTtnf39YgVgIVnVPTL7fvxQctUQvLMSuuy/MlBbm8IdzTHlmhWvben3PaNhu
ni5hR3VmYkCp+H96r+P8ttDJpoYoQoxGAwmFmZytWyKaWTIVe5c4nS6pvHUSqgTwtjMYLkoAzdYm
J/iJ+xzKPXNhHaAybrTm5XfENDllGNVYEoPY/XeS/pKLvwf71prYGAvVGZVEASBD6oRULF4Wlw4t
BY8cjq5E1JoI0A3YtPyZO4HyYsINJDdAy77dZtEm3ewFAsVH2m9x2hJGshb3DJG1X3wnaa6nn74i
6TGEGB2hqHUfz9SJNvDCX5oYM7piFcd7hxdcX0hlo9Y/y+D7I4XDmzCr9IbuWEue8i/7zTCiYLhY
9Z4ZqmjrsdI8cDQz8zQYxZMAaf4kYm1PL1g8xVvTWpNB1fy1sm5iI3xgL14H0m7tk0pRjUJMbXTc
DqcURpkG+bVd9swqZljvbbu+eqdUI7rK2MAugMfRddRVWyw3J5TYBsUEMNcsUkieKQei1OJI8mh2
9/c42Ze494vKaslkIvTvfGbmUZ2Ud1h773gfwSJYEHCjSWX6oGgrEksdi9nnea1GfD1OoqJy7KhI
fzcVQBakYnigpOnmOmUfKcH0Kd3xO0GUqrMnnfZou/PlfbxVgC5xYq7txfDEqE5nYJWdembc875Z
cZ8Q8ie3GjYS09BusZvaKBiVtsvu5mDwfkwzGpwSf8xs+KSWGJIcEEJ6nvMLGS82r9OoVHl5+4Yg
CI2m5Cb1yP8//57+CrrvDk6t9A6rDJ7Sx5qLGqicC+Aq5Pt0hiJSIfiOpao8crbWuO8dVwxwUtwS
WC7daqjdWZzcYW11Z5+egIGolx6yZq+lwQ2tQkb0jZPWV9rs/n71M2dG+BoskqK/LBFPXTN/d8W4
86fSMqmWJ7MVXTydJ//dDl/A1xoNMg4JjACAuyR+YCxt9mxZ9c5nfuKC82Y9z7PqNefns/J/4aBI
UeZj6s4+kDIMomCpnNkYNejXiBTx4qysgT0jIRZULt8fFNhUgEaA3noAbqnWPWvIfrwPyfsaPP4N
v5dRg1vuzPol0MAH0MoMwevfI+Wv0VIKwMUMn3AMdHQ/NFHSYdLSXRWQeBzjRns1vFjKhPXliq3t
TsSdWjv3mZ+WuGStS35Cs5tNhxW7TjIVHvc0LNTqvzpLvKpxPmvrvSoUmTtIHzLlxI5Xw1ixnfpS
NYEsUtFi/TuVb2/vUJ3sC8bpuwvvnyxkTrzIXyN/kHVVBEmvQCozQ+Eg82Mm5mwfX1LAxNqd3Req
NBYW9Vcgupo+wJjGRb2qbeiWX33SiDaUwnkdZT4P3BZB3WV6lR36+f4JytbB9NCoWvDh8956Xoe2
2yKV0T/VujYRZQhQ+rTNn2F+jMs9GMDHtkIPIoO7Jt0qzN5pe5MzgFbiQbYlqU/MReGe6u9eIsKL
FhkkgRF9brjBnazHHoi/FUgCGAnyqI5ntOj4rdmE/1vyaEAF8UiAzx+RlZw84SgqcOG6v464jXSc
sjfFz4xLP8buJdk2MV9Fn8yD8rDCjeII3hA7vCmLNz0DtCnWD6LKyTcK8sDjnXYYLT+VOvQPE/vm
K2P1BdEbZPIf27tJKa983VfznyT1NL/12Guq9wunJIjMNjAo/4Qi8SZwUSkgTGe5DPm1AW8cec8j
qgmbz46kSeq+uCNEA3ow7xriEVgLeefHmemluj1U074NdnNwAJncJiyXECKdsKlkl1IwPIrBgcPe
jq5EaURiYC+vvs2HdyO5wJ2v+cPC+t89XaLJ5l4PjGtxwq9Ct4g0t0ezsSTB22PPCOakG1jrK4MJ
Kquf0/oQtHgWvz1qlrgGa8clgnGoipmMv2YbPtHF+CtAKeHrhwgkL1jyDJoefQdfM/jpTlqfaFJr
LyVF8FTZKZx0RNER0cTMO2QW70Uydh2cXbnLsCPCVH6aQrD72okPft66XrC7mDgKx07wPK074HMN
f++T9eL2OOmeVCXAqbD/pRkl/Ev/cfdJC15VHtXHh+vq7FhV+1+IsdCMiMIAzQPdSYj3sPF7nqNX
hqR3aJse0EOfpxpKKuITsxQh5HKQ3jHTe/4OiLdLSV3Z22tVmTzuRwFVkswhVrTP7+84sNUS3YYm
zMiCLbbmPyf3FbgKNfQ7ECuHdJxj+Zqmt6QuVsmS9Iv5YnsAJG6qrjxx26WM6KGRrznPSFbRIaUK
/VlUsW7t1oJS9QnZWPw/FCo1Cn+yA/f+LuP91sjRgmtxI0uLyQlOGYSG6VYkstULCG2mSvuBNk/8
tU8DEnQA2quooR3hA3qQQppeB0wfYVf165NOId9A4IXhuphWc4Y6DCWnM4XXuasZrla5naUdVH0B
8ckst8LSLlMNX0VXAJc3ZyCmRPn36Sg8437WLTWe3IT+6gWNT/qKbE+vrBB+11QRHaYx3UYFRe7z
9kXruJmK4/hsBb4GIOaUjTdRE5drklSRDJaMdHhGtD70mlRqXcHKqQsHQtDJY9L1/V8kLCluN/HD
Oe8sZS8u0hm0xab9/Ym/+jlqNVVharXK+tlzo8nLnO9mU0LV2D+xb5R7LUtGCNfXW96SC0IJC9/r
Zr3ZxrH6/DgwFFIdrIauFsHfcYdbkI5/eo2Ghnzec0z9pq4g3K29Xtxagn1TJDShpy58F41cyvM6
G3JCW/KAe2jgcE9aK+IT7vkf3hfDXjUwZ07kv/pkTZMBZ2paMOhT8aAAzcB7eXgdqvZOzuuJRvmg
UdPq7iZK7mGNaSkzUlRzQCJYKuGCmhiHui1eiS6XDaIBXWSoZH/2f+N4GyJugGx94NwN/nexdoa8
NZ8QE8NrAbl3G+pfpJLfBm2JL7PalqOOOuSx2AccLjiFPlycnkyVO6AwCGxGUrZNBdhiIk1m8uVY
BEOaBF/iDKAk7kI+c2N8ArAOScu8ouwXMaAksKOiZfMoCytMLi0J36k1i7xEZQjN6Kp8oReDlyln
t2RU7ebtEfeEudIoOLTnCuXeq86ZUmFdQ62JM7H3xFfqqIsjDk+KxzV3RJzt7KL7761KjSz1BGp1
t2Uv3Xa+bUWsLr1CtivuMMYwnRAxCD/heT+AZq0XcRhMvVBb93jh1sTyavuRmWuISFpLCCp9gm5Z
v7WKaZIS9b2Tlsla2KgE6waieo8nr6D0w0RWiTjzTmD3xetkrwUFBViNhF1eLB6e2AUCC2y6Gz6+
4wjm7PcYjnJ3tDdgsBtn07sv9sLZJFsnWV/j8lIbV1eGuerrMYxrgYy/MiAqv8Yk5HCDPMxoY0ch
tHC1FGh/pZr9A2R5+Q53hwSqDJ6TCyJ3elDZlxMTfFz9FHPcE5qZYfb89jGhStyi/ibHEfticJdJ
gGRErjKIZt30+n6v2r0JYBNSl8UJovJuLvSntF24j4/oyajP9aIqXcLitoPSYDRRfax6bSBTxfNX
xhsh0L2twtDt7EM54+X5Ccv7AzXhsY2vlOo71by4dV5aVrwl4Fjv0NAcMg9mXY+jaQhA5Xtcx9jD
HtN5xVF5MNO3WB/CD13qF6+kyax3kgqLAKgnpSau6KTYdorDKZwgfma7Nk5q3R4dTPw7zc6vg1Ui
Dx7Q00JHsXoU9Aj8sWwmBdtIdIxRFvqPBOt6QvuCXGUe0/sXSRSrB7Lf/Jp2ehjd/VooxAKNrFAB
MstzQaeBZnbKaylNRKYIuQGMbZViX22c1IVfvPOu/fAGJqfwbekLzRFPrsJSXXuQwi5vc9jaU6+t
zgE1DH6g0NbS1H/yGsDEbrtbQHOA3MIlk4nRlIadB1Hh1o+YDiMLUcHAQRSpAFvlmiD/uF/I5B0m
LnXlg2tXSEsXrDGWrWGLgOLdnUB5KFuxRGzHSz7P9fwshRI/saRc3tRvpln6rI04LYifpu3Y3zFJ
3vXCdyB2aDr0NXU94bnEzqE2hA7cht2f96p5qhLzw5nANu9VuPaEs+pV2thtkoiznI6TG17tBnM2
6NQTx+W9VOZG7QXO2xWiRV+Hra+TpxPOOHsbayrvZfaOQSyIQEaqbcEr3Ln8PbRlX5ria02rBPCh
K3pfoec6k827nQgHLVzKYXf6/n3cij/wUT6uia55DVauF159d+YojQ+VLVXr00bYHPotF7Uqe48a
/hVm1fOcyj+AUnnRvvjM5OpsNrE+eW6YJcR/B5Kkj19OfztemO1vf/9vywgvFpmwdib7CDEngyv/
WMA5hUQOHbYlTy/A/du6erpV5HwpqevdNQB63nZTWvoRXIMVSue1wWGcs55zrd0R4MiUuErZhMDw
g8xyXvfTG6n3y2/LvNNH5TNphZf0jkAU/8Aqi7wEtOWP8Q0ZVOBEIW9hcLsKyiLxMSf4CFKgburz
ByT/RKipP8s4xH4RD2jN91XQ0Fv1uPlvAfSPKeC5SprFiUv1en3r42hE9ARu63cs7eZnmLZdmF5y
1UHcKYeEWdOsSvoleU0dT3k4o0qE+kPnIraBcrKkMkZ6M9AmlVhDAoxvrAlEwDZJzluYvIT0wcHW
C83Kn/7YzPI5BdNffFSB6grju/MnH/yO4LDBw0siA0lHruAh63QSdZU5RCSru5Z0cDMSkaG2Cal1
NH8WBE5CIOIbuDf+EoREjJgInuXuTzF9I0EOOq7WC6SFaFF94oNk3uNLCt2lgMKRwf7K4cSxCsOl
YHK7npRkMWKsYKOuccEMzPf3moXlYhlB8Zy/fR7wagTG6IvBMzh+gMCNSFJFoakn1XqL7xgdaQUX
81IKAKMSEJ20KtAq7xHet/+dCcuQ98PCN3zQpYiXHWLtcoXuZH7JV2Q3CsvbZUTdNdGt7uW9BXHj
ZvDw2q/A2n/5juqk95PA5mg54GxYtOOkE5Qx4PzmVHgF3mH6XMWCGMu2WLFZ9LAnc3D5TuAjxuP2
+YL/GCAVG0WrrRSRM4542kKjKtJm7U7YoANgyFHQXz6qTkgBuriTtDtsrdvNpZXAmLwJXWFCN1d9
+VWX6nEdxuME9wCdCSsqbPHrmwzx84a+bE99LR3jXrDJy1xWZJQM6JrgzUzRTkAGTGucUXyBDqdv
SXiN0y6MZqfQydiJmXBvCECeE4qm6Weorn4HZyogCqGoodbG93H8usO7a1/4XGxcr7OtUwvO+/By
2+N9Nowca+vfeFZUltXU/6sHPzfzLbpUd3to+5whnTLX79PrtcdH39cFeNSvqHHWm525qZXqeBla
ndUrw1a+E/LNvCO0LvkF8027Wyz/8wIcawEpZYcyD9oa9zgOIesvMWql5oy0uuyXVuTPgkYO2CSL
ATe3bWEqdS4j0drvTmHg2fgrBuNxSv89hwXIq+n9cO96WAFFEMqnOS1PNzcEKNlm9xhCWLMZj0th
OLnCF9lR2HzLnpWEGrjk1gikfoo8z9Qenqt9o38XBl6ESPpQrxMOzFjYsHW0S5qNhG8VNSj+EzGB
blwxZAjQ6DqK1HhLD0W3meJYWBldQZ5SDi0suKdD9Pbw0urL9roRX4XCpmCar8k3MLLQmitKM+fY
0yvvJLy+e0Wzb03jABd5p1NxTfrsQw7T8TaKM3yBxzb2ndSmRXqbsHHBOmdwNlOc40fQaCRy4+MF
DjszNtb/rmK7aUjxlhJA2wFbp1DarMzwikhDnHz9FzcC8lWOk3ZDwNk6SLGJmYSM0fVUJyc+jiju
IZxdFfJOxybdhwokxm08QH6UT6fBeZiG4IyLBhMN9w8DzEnbgY3qB0cXTtG9jmcr/n7MU8QFkBOs
iSOGJ9VyZR97X1yxYj+4wEL0C0zdUfBnxPcEvocCPIXf174xOajFrHryhIwr1f2OsOXqZE2zm9Ne
/e00lTpLbrJVVjLwIh62WzSwFUajHvJ9kNKzRAQezJ/Yz6Dn7fYRsmze4EVyXyASFScFSkb+Mm+k
3YNI83s+IvYdky6a/krCOyQB+uMuKIgSdmM5LMkmJec8ax9rONtJM25XmEX6vqLsi2jWNn71OX/R
r7bvSscOjqndqCtu+LdOokLR2NWIbfUREmmJVHI7kTcNWxLo9fim+Y5UvPUAkWZ8M+tbVwZlLzRQ
aXYIrNlwMhwvEO9Hy8yNy8FXtJoWOrippBL27Ku0I2ReMr9+5oNAHEGd7OV9mfncKyPvFgCIuTTv
/4YiIO80kAPVaK+BqpUxeudQ5xL1w2ecMMy6XdaBP+CUCxTMt3g+x8bCPd3RHH6KUlBb+kbl4vi1
mTI+/fHweUqHQMLp9AW/6O7E1NAhHAUq5OAg9hoPpgKLW5SkU0Wjvn3xEEyz7T8Lw9NHdI4CF8nW
VDUZH0l4lLTwGhCDrNUamodaJ1LLcJ4VHDUQTeteb0D+0euu8gERfuIYCBA0oUz57rrPFutOh0JD
Q7yh0LSkVitvsN8wzA1wb/LfQVmU4fxSedzDhyPdnBFkuXzSzEzA7dLmgzZl37NdsQQg0EJxU3Su
ICWM3FLOhKMMMjUoCALtZJTZeAA/C/31VUzbilkD/xqWss3HdyML9+UpXrj5FvSv7x1i6Eaur7au
u0zP/vve+mvV8JH/s59nm2EacKQgemR0Sop7d7xzb81IqPNQgY72gHZVjuyahK7tDI7JyjGBkjgU
th4MiEp1Af6lMRtoC1TG/fR7j1XaKdPmvQnnxwTy0vCD3VLmO3WS1XCx9NZ8OSQQ/7B4fDDtZ5ZO
f2F6A3N3GrRcA82VJXdKJFMq29d8SFLV8v+zx7jQYM69khm2wybWXEd7QKjSb52gMaZChlW0YGO5
g5y85YYlor9uv8/wp75HW/iQCyCMwYPLCABKGDiw43W77EKeBGfJFMfHVfbknz+l9RoT/3+LQSdZ
AjaWmSan2Ywie85gDjnIfKk9S6inTKs8ICN3oWEQfERqZ/5na5eJDuDUnrXk2gdmJrzXT4icpmZt
+0fKNPCIB1TDNeE34ZVyBOr+7lxbCQAq2mzSgtZ8bSSX9401hTBF3p6SEwfa5ildevWQxSuMKlA4
EObUv8DAix68Z6Ho2eU30x7SNnN3oVlxqlhwcHZ9XTxhEt3FpgkqeD9cJT1Wckig0ZU7tjPPSlZ9
xZ4MM/BpJtaHv0chBiuZ6dOEbaTFkwaRjW0pENUTtPuk8vdQG2dTvkqRGsnUU5hDBTPREtFgfg+Q
e3SW2kyPA3lUc3O0amC17lJWG7NO/f8s0Vh+498qlgm+DVLBTGxskgJ2K6MujOV3Ulf418GtgGBj
oe+uhPeWIwmekXAou+2DToxm1X7Jr6kuPAcaddTo0gDNg0B/FTEFmGsuLg5nhgsCR2hF6J4nUQFY
X5LjPk6BxXGEckiX+3Mn+uhSyA6AQF+mEiw/0GOs9Nvvs80fV8wM08chFUIFHse30T9IwYPYNYi7
OFk51me3uOQq55vGYgptMhQRt9KXFQcCJ/2vqfuVLYcQuSexBwbLIQOWnEEH8elIHvQwhNnyx7Ps
UhPUlEOOY4mBYjO5WUn70uU/oi8mx61Umb4PVWZf9YpMMtPM+4alnw6zJ2UP5kMHaK8Yt/Ovr8k7
0cCaaeUDmyK665FhIp7uIBt4QMqtD4YzcfDw6B1E7uEWNE2T6KXSHguUWqD1Uq3aMOLLTnU8pyzs
2PJ1Pe0kZezqja22ZmYmCg7ySEisSLm0NDr6kfZD4Lrc22sM3Dwu6LQHAXYzlAjtTF1wrsXT5Z/a
2TBgtVxvy1g+XYm/vXDOJirg3jcaD/k2g08NYayLbD4i6tLKPdmczC6rW+Kw0nwfiFs3Qea8I6w4
gyPmT//BR7IGNCy28fCSDhuzJDdCuoZv6ShyjkkwpbEbWsqwlQdqyCf3URcmhmAwmWFPeeGsgygw
8bItOYQZ2+YN10gUiU7aV0ewDu5H0wROiXmli+4dIAywWebDBA0dlC7hvraKbIN3OzGBZHgOAt9p
hebzA3NqYjri4CW9uTmAn2iJwEjTXlSmHoJlmmZXeTdiE5Jsxn3UnKGQH8+iDn0jzKEQcBgSnXjS
57/zE8KLvo5ay7eNIg+j9BY8CmDMsT7bRh4atxGQ/G7ez6oRcNEK2khxOOl0IYN9PXUzon1+5qZf
SrtQ/TR6hng/SXpSushN6m5ScFlU7z0e/ge8rVvhmFrXGTEpDFK1boiFBHxoSYwT2/t39eT7DvxJ
NkKD1z8dfcNbByWzMgSMT7+KYULlgZIZ6ucMIgXMuAKtU+QVkDho/5fCPSipIsB13XGivFnqEjeA
zro98Ot631s1bilx/4dcvD5To2y1mP4RHJHfdabPHOkVf1v8iQ0R/qYIb+kNAMOAlARmDCgFW8yJ
BERiWkBuXdlYUT1DDdSDqMX7PfPS39sUTaT/AixC+Hh2nr8CIkZXdmTB2w3mLQRWqY/0GYZbLaWo
aJrvtK/6ZHDiGQWx/a7YBJyu3FB/7U1v0ApkyX03aO5bNVMPz5L/34fEhRXBmyndjkVd+mr+pVrr
OujaFmYGkkAJ3a1QyLqR9kH0yhV0xntnrPKvL/8eQm8dOPom6f9WRNJnawzUsSqy9hKqvrldYYNM
AeQVt9y3IRFrWwfkW+UT4wby6eJqlGGJdEdHUGv0dg/TUGcA6sAfceSfiN0prWmVZB0IBLMJyvJU
ewRGhc8daJCYU0NR70Hr0qz89wmnfMBsKtmg8FotWJ/uPXhkSJkZIDCHKPKwOiPKe50GXjS9eb5e
8vbngFEAGgJGn1m10DXqPjyJA5ba5klmyC/AEnadIpWSzb143FSBaM+yrQNRx1rBlzEChD9YH4xa
aIZ9X+Y8QtsNqTn51GDYqzfFdbq2XDOsSUaVzEjo5+eNoWhGfH9Ms/hcnDMzoxBuXb2tl+iLn+/4
aN3dqlxoKt5Czl60s52rX02jZIrMa1ZB4bS2e6v6PFgTpXMOpVpzPWk9nEMhxjmzRNzF8DeAE4Sx
wB+DHLUsWnGt/0hrQBNEEzjYtUknn1g7NmHrWEe0Ff37yNtYJqMjgGJWXw0FMcraqPT89fSKRbln
pIp76xTxo0Az7Yj7FxwYUSq4CopLty6WPpJ0uQqKEawMagqssYuoFe+dB2pRb7s3pmqNCu2ByaKc
/46ewteRA+cFBIgKvKWnOWUUNL60mp4Uz2b1+FsBi59Y3b+8m/A93P2A65o0RZyw+WoZ75yeB8aF
CpWYRPw9s3ael86l+FNo/RhOyZTn0wXfYOLMqWqdciwXmi4iMMlJhVqXlleu83Cqj686/nWUr7La
GKsQc+Dp04SL/EAON3jFDLR6dApvU+oQAfSG7zTBoApDz63W5RDeI7G35wNOJvBnmxeNEWSx+HiU
pL+Yfrsol6OyTrVTwl6Q+5w5/cDPYXenIrEPrQnmxb1/MocV1tkDqgzk2V2kwd8eVB3D75NN4y5O
PVut42hCU0NKkOzibBtXm2D7/9+1R7cYCginBM/zfxQdBrEg9oZ/3NbPk5wv0WLPx15Yew3mUq9C
5xpkZNu9l16e3UjNtB1oUHiPOmXzawiuc6TC4tKA2mJS8iKuSgle/GZFCvmi20mQarLFdyNiwJTT
FE+PxXWot39YePb02yFGOMS6/CaLRbp9wuFl9YI0rK9eDRAkDW9ErYu5D1wQoqI8OqCz//IRPV7x
azOE1rizcS7OhU3kaJG2vYrhsIBKwq1hIfYL2JEfQLToSADUVGnPY/TDcoYzvKA0WDGUYF2GfM53
LbfG+X22jqNt03qtJ4lFtnLzlQmGzk7s7ysadzfXltbZ+buht04U6LYlDQar+bE3H21qUdCakZ4Z
YM0ZbCPNBpcqiCn5ZzVpCmV5sbSceA5fB5lPJhEamyNWJB/agdTItdLXu84QVSaP7mcYfst7tWko
NsmhOlFJ2Vtbvo1Cnq7jn7Y5kfbnnccBFBfxXQ6UPZ+KK9Oc5HaMj/sLMgugvKJKlpT/9cC59XU/
FHUbkdbyoB1jYZDtbtZ9beBoTq+7cvIGgYqk6gTbh94B/XCwTX0xVjp+2LgazXDS23+HigKXeZX0
Hz3FgHlA2pF9XbPw/R10VZQloxfqKHHXftJsui0C63MrEcfW4TIcwDlhvCbU/QExa7Y4y6E1zJAf
QGfK4bhsGwxylmNoXWlhDOZe5rba8XKcRcz3sFXbMN1nay8W3BEYiv8KP48Rj3clE7E1aPOnRpvr
zbjqIFsJ5ex8Qbnpr65gV+VZxy2A+l7TRz+9Rby0JXYu5JBATT5dZPfaKYCzam1cYpo8QRGGXYgR
DF1+fayXHgrBVEy6ze6VOzDFlYn2r6hlNLBD2KqwsIgoE1jFilkQ9FAAWCgo6HwvM8mQ7pJFfQjY
Mtf0+Gcq1s6ABdyWPWjVr2RsC8njdeBYw8jQSrsTJK0rAPt8rQnWjm92dq1NVkqeW4i0PHlEmu+F
C+NgGcHB8isMnP2kCc3Ws4OS9N1LV2JRbzd5EgHG0gCQn17zU3Kk2OrhRDKgek2FaSc+sbE7V+9R
FmVJf7TeKY3hOSsuRkDJDEF0nuVGYZ70wGiBv0et5833iJdzC0mwOzL0MkHg7rLVag5pG8ZsaSR2
g3T+y5L5TU76qLBsERAJk2n6EOqIugDz/rV1yMz5Mi1QESe5MldZL3MKWNmKrISuqYQWX/fWMy6X
8PKbdl+7VS7dKTkUwNAOxUXcXrRKTuGbjim/Fhbt7pooYp1E2ZDV/TbAflnwyLCpxWi8MjSZKutO
NIQB6UzahjkB8g1f937emnDfpasNYFStlc0lbkEpEjdlCH4SSYJez4lgdsRfru+qPFQ5CBHpY+WM
gFCEgMtASxJIZhFrhXt/DDb3xXOK6pIOTvs7YBALRz5mMl3wpcFQnUesf8mJOYJX8Ol3pGnf4WIe
fgvCkajtgZEwXfhaHCMFKj/Hjp7KN5gjaCI0a8AwvUj7MiFs1jFRRveE9mQA5Adsu0THmatMJMto
bJc77I4L5AyFpX6N6UA0j+GSa1fw/PVI25KxhPHs/FdA6ZiPTJAG2eLkX2RaNOgdtnu3+mlLkqSJ
sYmgCXR1dwDSKvHKOEZgyFArZPF8Rrp/ACmqCx7I8OWoVWgrymYqwKaX0UIpQE1ee4HAYy7ne/bD
rZtUjw9eqSlxe3KdZfODQpKYy/b2W2hYSrPcwsTNYhG7VBrByAISj23UufSpVbGzqMSUA+61HHWt
dHuJ+2LvW0kbdxtuJOvOB/RGPpHrJARiC20FWyoysP3ZR04YkGkV4n/38NhO6X9QKO3HJbUZsePJ
5G23GnCwqhwf7l3PgOQa3vjK9mcXOsN86dQ8fmwTcbxabPsaREG6EGd4PYpEM+m6KLokeIuMiclh
KQjBfW075wsPFJ7C8EPkWcSrMuIb6Viq2iFqG2PCnIfUxyKIgd1pnhLHZItRR+WlQn728WV4r6UU
oCG5UyKNUGuvLGFWodbMOrHKm5rZpqqsUjRn/BUxt3Gb+SWl3+t3N0GxrTv0ZqN3MthhLV/lG2+Q
5ayMRNd4tiOt1a1EewFJ6G1R0OTR2T32HS9n4Gu3VjxCHLfH6SulpO599pKOp/4DdkHyEYX29+E9
WLKzOu8yV5cf4Zoc3xkpcVvbAXH6dvEvkrnDQ10U8wPA7QzDE7Fd78yqxdwJhrtDtIQgkLjb6Q3V
eOyaeEBB3K7O1g5Ju6kcKPmrM7mQ4fqp0tbYk7zgEpwyw8NdzMLC2RpvbVFnWHDnKgYJgOEnFJrF
z2XcaYBHlCxHPgYOb7mwWXH3YNWx2Q8rI4zCcq9iHbYK2I8CB2K5RQxe6VOvoVt332lTQ7GH9HKK
g5LvXy1JPs5wb9juSp2+rWRVNYgtY97AZeI3R3IInHrE9FojMrqtXRfNvkNwvUEHW05mhwA9DnKs
zxLtpHnwB2LharCX4zd+XQ6aZrrCixoBIoTDlttZmnb8+xvw3bkKfQoWfJukfok2Nnzjlbyw16Fs
7zgInA1RqfKhh0CdCeGspWCb4sDbiOwRd+jHEKSzxB24X6WUZIpzYF6hJnhBO2abp3ES/NM970On
UDKwcr0aRB1Iwtc6nBbaEzCMrQ42dR0veJuQivEFRhUGr2oN1tklFUQ4XImELf+djTo/NKps93G4
dSRnELQYKQyf5Xfy3n40sdDspyalkoYc5scRZOy0/zN7dn0rX59/rUaRYra6wryYLtVtUzhPjh5v
fKIu/YTzzcsaaX3JvFQ4FyS6unezQu8Tvl7GgipLMse25+lzcQ10rX3RHSI38nz3ArAJ3IaKdxyG
iuTgumxQ/BVwFYeAOf4n75s1uUMJMN4I6WINeYbwJUl4ZvSqSoQnzMHlNTKul8hlzZMboAPRc/cd
KGszn1MgXdycPAbZS0OAN9lxjWPBWj8EERPg+A6BWy2IDTrmsQxkF/8KGTk7fkMsJu+Qn46h+NdS
RtV7Fd0CWvt1cHr4D91dONsl2rXpEoRYaHrlo0YqOEI+PxE0Nc22IpFnml2XVnKfVaQWqLmvJlQd
JLMOvDnwFVslODprEjiqNZb/jBmVWS93NBJA9hHDBkhnGyDc0zHAfXlHiioP13k1SSHa6QsdOLOy
7+8iHbcwthGSaBQIFIvMeQ7KV4d2T9kycTO91Wt4+7b6an4uDzVD1wJ2ZvR3rwlwBjpg1EJ1ly11
VsEzUJyvzn+LVEDNtBXxA39KNJtvas/M/dHvDygOlfZsABZAhk6Hc/KC56piYBTAnxjlRZCp8tY1
ZyUVxGWaIcshoSp/P+2o8ZpvjPaNunpIV4RzbD6lFWmmFraPVHnnPqTRHbp4Y+1NVKvvIO5C/74t
NHKiEIBTBWM5znwktiPvoqdSG2fJrGnDAflPIqceiCxAux3WV5o69cKJv00LFbWQR02rDYIjgFdj
6zQrJ39shLioYc8Oq+BhU1ATMfzrwDTgwdzVey1C77NxSx7CyIVM/TOIjUruJCYjFW9KJJ+Lh/Hl
THdEExRgDkjZNboPE1tUpTAuVXNbDsZbeJyaoyDmRV9v3MGe7sjfRPIOpc33EFocAxVkmIRedkZU
ONxn8YUiF5/oznKBJ2KG7tuNSWpDM5fTs42UGd+XE/BHtSLx1YcCbGYWduXQvr5lEDW4jz7BUboI
1mDLQ/QtIAwjwCN1RfmVbEyHxrMbyQjNcIO8a+gEhJQyF88suics6eHifAiGbOPbkmqNtw78bxHR
GLrgAsXcdBnGctF10T+W/HkLV2N8nfKKLUn4Ind6GYUYaj3wNijvMcvREBqZ5K8DXUp7AzgzykZb
paA2ri0cXgiGKd34Qsg1j9OgcpWp/DvkUK5qenl+3y2A2Jk2aa8HhfKveHUEyaQJYUaM7+aOjd6M
jgghU6nLDdhHKbXyTKZgITgg+afuT4BDYDtsgP+21ohQxJ0kstU8S9MPZPjaysd8oXVi/23yF+1i
gE/BW8FEQ6NUaaBlw9hDkF9DJTrvB0DqVbpFMvYxb7TLPsYuvZo6qWPhd8/Se0DGZtZPDD4O5o4z
DwicK5UCLPXbYzLA2Ux/ulnL5nbfV7HQM/80Jy7DQrqSNaVHyoZ3XES5bh1T7Mnv/XDqxQzKl2we
G8HvBwqjNyO1bpifhfd3QeamDsp747350gLqTi0mnXy9JBTwah2SaMxZjdz/zGAIhQ8mlhIBmd5R
lCVAmjsTzQLQK0WqqaMhiImGz6mfNUn8WPywhUJ1yuabPHAqnxiW5GJcrYPK+MoEaMjtkGL3Cyxt
bMb+fiji9Rcp1XEofPiWwuv0qMP+fE+Oj6sdXb6YSH9GsvMJpxK7Tlj5CcRLZ7TPMo3G0XmuIMlj
awEUE4N+cI6FLx3hY3DtrZ5CvopggEqZ7SEqhQTHZ3EGCERTjrDypZ9zFe0L18e2lsx+WBOS8PBb
r9JDZR0yYLiK5dWx2Rwa6rfdPE9eYPnhLMJ8qxLsTLJRidYH7jFZBRcjvFh27h1LUqHEWmW88ykr
DBrDcYyjxGwPBKdQLAss+hFgsCtOV/TfKMSFaW0SaUqvFCIvkGGlHKUOUvFpSCJeuex+Q5OEW2Vn
pirW6YmXJ7Bo/mYPIpNp0NWYgWkX/VvcfOYyTUV0gi9yi8RD6RagsfQ8YlXK3poe2gsDq7l4mMB/
VAyJ8/GxwR6FljMM/vkpPcDJBL4Ruxejz5PzL8bpt81a+dPAfwQSimnzVbuUqQYaAEFrW7CAwNmv
Hic416rECP8zrHdlzpOZMWCzbcl4OJy88sIgsEZmLzawYepjJ0n7fSiCYbCHwBCrmgJt9ZfPXIub
3RALyeYOcNc8bWjd348GN20Fg0LgJnJF6uWscdEeIXHMGlQ7CfUOFQOh8By66J6gsGKCxqTPLxQA
5wbtJ7OH7ptspeOjRzoECTnxEP9pPuUqqJTBASmmAt+HqWS0bDcqPzhTo7VIszOqtgyUMG/oP4Q8
krJJmBK0nXWDZu1undDdmHzlabGHA4ytsAdF4gxpeHB31H1OFUIMVne682sjC7DPZsJ8udChNYVf
smXMja0WAlc/iNFnW5WjXGzhN48hc5wqDzwD25REwmZKaaLlxw7x2IaSDXYqL4SzyQ2ccrKQMdOD
I7YyyPWVpgKltXzLnu7hxp2P90HgVlibnBrKOGfpzPmyWR3yIPSsRtQk8r296R2eIAcHtUobucfE
Ghe01HvLnCLaBsV+O2OwZ13MO6zF5ejGl9rYwpMfDhF/OnY+0ch7VTvjO6/06JmoV4waXQ9JGMIl
ik4KI8wb1qxP/ekG4VYVb/LOv3zqcAlQhA1ausJnp57IvseMJw38LPsP2/jyQx5LOz8pHSppnAGi
KfQghEmZAttYwvJHZQI5SnsQ3T8VdCDADgG5p1RjPUakj9ouKlJMyOAJCc6e/QDYczHV03kCeUaI
lSMkFEYoLMRrHI34TzkDafvNWo1hTQ2hMhBHm19SDAwJ48Ni+ewyz7pfAbxPP7hRx6sYNgiiWcmj
kS6ZGZ3W6ZZEEvMAuG6VOX5eDPq8bVLp29Z9KDqrnevpv3wZpGuIyyPq+HwiLKSSmEdMrlxg7v2o
bIFqKhiolz7GFNdTcrvk4jVgJSmUblU9GLYJmiB96UBEbJd2svrjbADHdAci1gAo1U7Sp3ZQ0u6b
WFgUAvwxZclUA+PQbgPNnkuDAHkCYZyxwxsJqn6oH/BaoU+iWE/sU5j5Wetn6e1ApBftCBguSyCJ
HJvesmK4x2HTv9EthvoNg9RD55HB9Img9CenxqQscXcZBZ8YYjBbMaxmDPu6N7IuPhXQi1uGKDIc
4HQIPurD1xknIjdyYPDnNINNk2PDBWrG5RLiBNwKReatwbMF7YD8Gc4yyw2eLG97giROJqOaQ2/V
a6E8seyjH2jIlIZ6WviaOw/gWjoaQruSDuh17mMrmWwckdMUyc0P62olZzZ7aFgF5YGo5qCU7dbG
vEh9HVH06B4FqbeL53XyDWyxFLT1Qnf39AvY3Yy3uW6DoYcQmhuf0Bb9g+cgFelgOw4kiztfmnKX
RhwMr3Cc/VIMz/NmfZzFnKeJ+FKRNkdrA56VQHkKe2OaDBAJKQrNubq3bWSSAusKbaZVHFmbSu+8
ksHxBCqolkMKGF03+4HOwO6N+QrUg1VhMk5fXKWxBu4C6c7VwRux5N0T2ybPG/uR0+DVE+eCRvzK
TM7Tpy9hzULKLH08R0Jmmmms8jah4CMR1XxE60Ka8JVGxk4aL23VOwgUNNEnkDISnr58Fj9+6tGF
0+7UbH17yjUJ+16k18mybJ+3WRr5oLzque+6WnpXuJ58FUn48wnATqk9uRAqMlNvrdoMh7x62fBv
0ZZxahbOye5xlTAzhYDhsAUg2EW5nwx2TLEOo15YjguhtdhS2byXfilhFLVcfZLR0MrlcZAJ82IE
WbCvMUu0FmcCKrJN3fhuTIXfOenUT1Ktn75QRrsV3CVVc++Fay3L4kkE+uScdAgifSygKIvJ4piC
dRdpBariHxPnGNYNoWiR404nlhtojkii4WXQo0IT0LQIR6kh+aL3QE/NfTAn3xJj1WGcZgQUugzW
+D7gANIzvBftjpjqwcp3aGwoc0Pqc1wGRflUAYBBlh6Rj4DHuP9SGpp+XGm3mluENQRTaaaVlTW0
iya3ehHFFLGr+Oar/eLu5Sfl1aqMSH5d+tqQ3fnj1Fax8VkqmacEOCN/tadHv2OF7s89l62YrJKp
1bGxRikn3PM3PxM13lAfMKoUAHWLZKW0kekm2m5aX2tmeTWIa09IzVGjSbkZfbv1MgomVwlvcRWM
Um8VwZ3GYfx0DG4zKSrfUUYADb0ufS9c/igVgX2JQC4VTQvZzpkhg+kQ886XmnaLq9hQCiwwsNLf
0qHCRByCnMk/bGWwBPYI7iYKD8xu1DtEfmC+XG3iUd4UI4kP2CNloOAq4Usur7WYBUDEDZNumhre
V1YT5qbqI1mmis3OGAuHr3F7XA2QL/bgBqFe+yToYjO+aKQwSZEn4oT7w4wKmQX/acMHYkWCLtgZ
VUSIYUL5J0dTJgZSfbNzPj2EZ6ZfXEvDB2xhY9oThXcFyVvGamOmn36nVJnoOPxAQQaBaTE1LyC0
ZIIcsiGny4H/5zkO4CzyMuyJnkpmwDi81YfuYMsqyb8ngmBc9RwyqWWfA4KCnR1CvMfiTkkCVvVt
08EbZfWmJ1BBzNMNS6Emj613zi76DB+Vlnsx608qNi01ZpJmqR57PgOQUl56GYWFLbVJsE0lQ9TV
6jsNGUhQfw9Z7aacCLcwi6npvqU6Hf+nbrMBP0+XcX6BrIdRkf4DJ25TJiDrm+0yStHa8gWf2TlS
TNab7UzTtPvTNrgANqRj0olf2uQHgERsP4LZ1cS+5cTQ85JeXpx22lW3QIw+lU+zcoKj5VZvYd8P
mJ0cztRykQvOwhUTWV46xLko3MdLi1H/TsNA712WGn3ecNT5QPzljsegqL3Kc7W9GWg8trSMtvHu
No+shrbfsWOAnJLcBNks89mAA8OGJK8ELOZhyG7CGq3wmXMhPs6UQTUxynxnFcaL8i2yD0JLI9al
yf7GK1Fv1ls4+Ba4KTuwrc51NrT2+tlNSlv6yINfXRdr6VG27wGdxkK9JZfN+3oy17Zw8VvTdVsD
hkcVkQL92q0yt1GEz64laiaM38mQFSsgEYZnqbTLS37dloglRTodJQNE8TBal04XRejZmtMuQvo+
ju3vho1Bbwp6KlgKUrWWMFmT/7WsoTqmQ89D+TOfZ2Et8W+s+elBsPu4nWF1Utng/T+1QvR9K1lW
9h3Wt9j+otqnWHOGyenB+aST4Zv7VmpoisLUwLsuSsCikADU+t30QiK3DjNQcD/+rwgwEk71TFzp
mPHNiXS7E+fMS2xtUHu4fIJyUSiiOE68cvPJdsFb4Tuegals0yetn0XHZCOEBxo1PPQTcob98NEo
Ab9Geihw/YHObz0RM01WaJQNnpRUo+dPUIHka7j8RGTwFCADNx1nevw5v3Kw5ZDmd+TDdgElw7wH
35rL1i091eW1sVreCa4LMOtPXBJrfLdPVzpZER9OL0VuMxFGqGq15LBsH4SUT+/Vhqz0/AvYLzEQ
GYIeNwPw932M9I9jmnSktURsqe1bpkT44q9D/q/yU4JQ9tlh0svgzLeHiEtEsyc+UTd8OxvGZjoH
0EaXtc+aWlgdmUxIK3ZCZukZ5cCIkpNplMl07+nJXrH64srhePo/dXRi1huDfUXnOCCIJtNr7bzG
wWZeObKmWoy1yUFDZYST56ZKYXfnSNYaIjw3xWt4Q0UCZyc18FSsSINVNvQRkHYkPDYmaJoEH6OJ
QLag8ySjONWxPy0WjBt8oW1Hh6Bg5n0lSn/uPfij2lgZj8R5pM2txWs/jhnl5MOqrEHeaveWqyFD
PskMZYi6DGKI75KRzzZv86xmPndxwJY/nZc+oqanVDw4pEXEyFQeWVfYnkSypChA5xvPEVrVH/Lr
8r4V5yl02n1Pra5RFFV7LoVmzt9Aw2w+Oa3ZZYZ4AZrANoTpAMIONkhjwh1lLChIHVeUXn8u71IH
EUoq9atcnC52CB2n97Yt+AsrespJciA/KfEJ7yxCTuShA4AABBpxQ+a4gYsVJD1FjvTLoiGD1HoX
5ZoAj9l8FCSE9qOTcR/tDTKBRrSPtIRCggrV1d5wKFz4AS7srjOV+uFToyb+UkB3CpBnmXx1ghTJ
Y7aVtYih+yXEqCWChphQxUuLAuuJIQxDDEYjr4kMbjM/z6TpBqRaA/MwFRLwzroO8XZB0qgrLeN8
VgiXTSsKZnmMKuQILlShVmjEvMH948qf2vQrCSRh5yNZZaYMjwJf0j8/d6aS4S00m/W/FR8nu98t
cof4HOJkJqhjfl6PpkXir/TM2ZHzqu37Kp4PIu+Bav6rauKTbT/Kif4PhkcQrigJ0TS8V+qi39uu
m4/xgsiqP80VYA3brJXq74vEhNGMTK5kKCCqBc+OHkT1uLmbb1hSQXV6027PxT+DnEVBP653t63m
CTnkbfBoV/Ls39X9KvKurjyhoLcAau3NxO5Z+rlI/YF+lLqr1CcBBUNcvs649JNnCB+jYMbo/BW0
zxyUJ9wnNXofdPoIqlM/X56yOThQ+NH+WJDGAVOfitCLp0xEzjNigNzAVT8Q4v6JsrLcyo607vWC
zUXjpD69l+3GM57RbzTyvTS8xSfpcsvQJawjnv3iFMM9zvFhGWNgrn9JLQW0PbOGoqhPN9heEMbl
g41CSiN5cFbGwgXqBdw6zo9WRNeohWMsHvmCLPa9tjIBy/V8jqGvBdlMKXMw40IpxcWqdRPMNCEw
x41iKW4hKFdrcfMx8cvMmkok6UtUO0sCwwtVHD21tSxbzPe+5OleimOI+Yd4an4RdL2DxtorOBL/
o9ja+ubKX8BlDxK1CpN1rvMHWuzPSOI9LIECb55dsPHZ7hFytzBXnJyQ+JNT0iqMH0Fb3sUNlXHR
Dq3oXleAKnssDucQ3zFQKWISlv+ZAJcLc5ybv4aGOKRKvvs+A+wRF1RlLpro2a4fLSSk5cMsFoyx
KqltrnhJb8Y2xn5u6LSrYPDBiv6G6a3vDCRX83oY0z0IzP4mRV7MfNUaoYClAFerjwpmpF4wnWSv
alBchdI0
`protect end_protected

