

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dpj1rsbRiC2XtvMMkZeaWceey8TRzfvuZghjsYUFfvEbx0wxaUtNO2KtH3hQvHr5R05ZRpFvbxnS
y9eflHJ+fw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RxF4+BsurVIN9R6VPOZY6IjRgF7yOLOJFH+DEaCvilnRUUfGXWquiAJNpzEAXSnsWuptbwUxy5M0
I2FA4+Rh4icthIWWJqsNOFS1K2ZEpNoHe2hVsMzmtRpnsPL9VGvgfvA4do7AYV7YhTUgoQfClGAQ
vFYxy/RbXBzM3PrDcTk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OvIp9LkjFoctqOSaxZyP7bYL7KElD3vYsFbzOXm+yqBzueGP4aoe0+732BJK3cSRYLmSREwKo0o0
Rv3hIBpxf0Y7nOdTTISL4pJ3qn/Q9Div9rDMzGaVxIOMLNLxqjT1ZbqCGU0LBxVzmDxHhBalP4V2
XUBBBCK3eeYn9YA+pujel3BBQ67ibuZRmgjKTwyT9B3SaGu2w8ce0O/YfSF/l+ncmV9cvUhjGdBV
Dsus1J4qhNTtraXR3S8daDpX289UCjsNh8krOgCnmBNlKeEFeTxbhmhnNPIAjDgfW1fdIgrmAH+S
tzDecIht4fghpU24F+FmCjpRFfArF8+d7uvxlA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4ZEqShxRoOQpy+XtDUXlHHAe5v38IR2wWpAtAq2KeZ3f4UCuk5LQw2Oc5c9xFXi1a9SsCAzYO6Rg
6iBcvyh5jboOYApBCjz/4VZfMAndhqby+l7lpAzkB6TqAqvqUfdVhSRn9DQMcQZ2fMALj61IBeLk
rnvtNe9XfB9vaA3zmlE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CxLbTp2UMBa44c/UwixvnmtRjPsy2Xb+fkOsP/coXETbFAb6XdUuKlopddrCIslByXBY8SiCzN9B
XnnZENqObWvYgo2VDZVlPu9SL8ZNuOrh2v/bJ7ztAhTSojfY2dBi8ojKva7J9JwGsRtKubJGASjY
RHw8CGw4rdc0A5dMEVmmoAymqmzBjExIxX3UWjtVz457DADxQ6UUgPgr7ysxQXkHN2eTr8eKtbK1
R8VALM11jq0MxZUpiiq5xDX4POkxGrs4QQL6Repo1WUK5V648ZRUZDaWyRJbcIm/J5ref1gzTZWX
h3koqZ0X3HGeO0DTx9nnC43UDVfA3fgk+YpVGw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33472)
`protect data_block
4nyGZDILKMqr624mhR80CPEgWAiOSI+hZabkUg4w5UyArYlvR5cVY4JE335nWKDZkPnZyBGtB37E
bRzMjYqDfZu2QjLRJFFKIilUh/0VVcgKbSnYtyRxEzthrADV2kUZ5E9rIS8cqCjzKxBN3mzg2ZYv
JVGJtJ5pvFyTJLexiQxOefkYh2KkPLQ2i0ej4G9Xb+b22xRRfoFvD7fAC8O/fLwhjeH/tV7vVW3F
7l9Q1dCS5rPVEXmUgKuWBwuvtkYz7MdGu2B4YZr0uWkUVMxhU12ZS909vNbJXNzdbUbl2XOFDV5+
phO3u8PG/6Z/axcp9zGaEI+KL2ZRuwgZNhr/abVWs+4BRa9Yc6jjGBH5FWtFygazqK1A680VSNF0
PWoo7NCmCMv+osbSpgiv7sqcQzKSRPDebBxXE0Rcev8un0dl4MqOAG2ZSZtbI5Y7l8Xne9WLCg91
UP/rxJuDQiQFaSW1WIxB0ZFomHvz7I3YHPQh351grdKXtJy2WdtCZlga0DLYK+mNZ/ugL3OfbCkA
mn4OzwAFTAslj4f0TRn0MEGzYJuiU8ugIUb8j9KKLtYoBb5h37lA0Wz2u6j88hxIyagjNAXhLtM6
8Ob46cNOsy3tLhpvrDWo7u1ua97tNLZPTIXsTnAqRHMLC2mOfU3oWP3ZD/kK8wrbN8as9R/ojNSn
Qn/QxncJm3eiqVwzxCSQwUdGLB8JHbPUSFHPJGe4r+ClEzXlwtprmMKNHu/Csuq96odOm/v7eDKi
JnPZlXRwu9ruS0YIKQJaK7j4ebFE9/mGXD5ShGYOeCcZajvHR1UjbHKCb2vHkCUnB3rkJ6WvR3X/
j59/kS7rj5tvNCSeyH9ekJoBd3a5HBEpKVtTTJ+tDoMgJAevZNGy3pkYvcTXD3Vb+E5YxKrG2UUo
z7MW05b8TwYrGvB5AOOHg+/YTcMeHlX2ljO442F30kb2CX5h0W9Q0Xw2hmDqYNv+/cbwdm94E1H9
zLjvAZ0/veQZi+uC9d+1UcpVYq4Vh0EAs57bgwIcDFrZBy4CL3rQ24ChHMFmQEjqRDLwIKoU/BuM
XNRB5KJEM0An59kXBA55e+tVoGUHNlJIbIxmH2pbiZTiun+eLIG+BLXkfJZp8L3DGNhfTFohMURB
o0FIQc5zc5RBl9+hAfmw2Mfp4wyjfis3Oh1Sh3qhCc4wINQpZWsjZUTLMQ88k7aMZQ7PaVWoBtdZ
g8vI2zBFM2ZGICW0PxzO7DSaH7Ppu17+yEjbf4AA0NttHGUuDPee7fENbkWl72Cy3Zm1nDHPeJ7p
g68Wg4AMuMcphGfkzOpVp1sskVnEDkqrhWopvscGAbsncOYvPOH4Mh5zemAwD9hcxWtO7cFERR2g
uiT5udnxroV22pfl8zaVvxAj3ZpjdTlAepT6JO78uonnQZkPfs6fW9Oi8ASFuLJaIqF82kdDrQfm
9wdlUfR9ZUbwRaa1UW2288sJe0DZgY4eiuimkC8MflikRqC4nOS54w7VvuMela9gowgHjIL4kVPx
BI86QEb073TC6xqDKQfhUb3EspcBtahCn/eUPZs2l/z+wvx8wUP0p99e+dmNiM10LuuOFTHy0TZE
h3gFb/wTxMejKbvyVfTebPeGqijnHtxrYP2cL9RTHzcgnsX2hI+gn/jGGFs+RJAfze+oGcjCgzjl
seGYn0JH1GPIyqhRfvpfOe8aCkg9cyeevaymG+lIrohtDI/MmpmqgCg/hk+JHnaN16q38k9t0WPE
jY3BqKQw+bLxD/G7hIz3gTxgZewPHmdCNAoHCjqq8BeH0vY/Zi73VwDhXEUjJ2ibVTHGU/OJpcp3
dt1qDEyk3SaGECo08FjIxQQLuNMA9DJZvJFdCWeRN7LQyGdwBb95tTxAyxquN09oWZuqg3NCc9WX
PSS+sGsqxG2Wb5yYftxmWFhSGcotw2Iys3XUYe1imVux58VE7YIcmbYdiPWgnObw90ijN6OOlqpX
ZzPiAhqB3XAsm33rQlKi3P079GFwJ0ZRN1qUH69YCYSJEk8FMZ8VuheCtPXLdsYspKiec8TTJ6UH
vEAPD8UPPEcmvvn5CO4ykkjiUQOcGIWqPs8mfz2LGKX2U2BXDckZr37NePBcMdBM8wQ32zOTGU6Z
6pMfSr2Xep28Joge7zII7QJnVgYHJsamj/cNJxrBGORiZE2ImxA0SrK8O6fD0MEEmvluVDB4Calu
8/eRYUv6gitZ2RzehFMoj9aGCVW05XigmsxhwZFecTed/f419Djw3SCtz5b0KssPUmO4voDdbiaE
17eW5SIIiyPYQt6P5buu+pYOPcm6ZtYuol+5HGXUfvpnZS4gp2gRH5fNm/iLJytaHLiaHdxIQl2h
8G2pG3s+iI5PAiG75LnsGCBgP4vZPaEHNZdtTmKGpTCh77lNr4Jpbomes2b6xz+ghoQ18Wra4IoA
7GKwCQx9jAMeKfwFq1Pcpi3949p8B53bmh3M2jAfMqExlSkP/dJou2rUl6H9NghfWnXz9Ll0bcDX
U3GrmdaWppD8z4JyF+AXNg9pPzVvZYdDp2vVjI2FB+xBgmJ3FFuGUzrZYputNL8LB6LYw3XDB7mt
0b4RV+GKoQxMt3/+a8PdEcq6ca85jjpd7m11wpz9SjPQ0k/9x9l+qaFwqICTpYSUmtUYDtSjIuFc
INIBQracfPc/gn7uE2ygZTI+W0sOLndDzJRzgKo6G9ODHwJYEQD9AeDtKZ7fMjM7zS3+jgHP5XIv
3jzbBuw7YC6dfB8ZzTjz6t5g+ez3CGnHtEgxj0tgLuCVi7HXdFniOb8QRZDisAdrNdl6u+GWyA4h
B5qMgDuGgZr1ULHNfSS2P3y8/LT+md+xRM/7MCFk53FXBY/FDS/kbKnSkAHnL3GrXB5jIEM9vCq1
UwBO+m6axUVxB4UZplE+Wz7RiHxfGrRT8LYrTadfFmeCGSVkC7ouiUYi8EGDWySlaJ0iA+Ncyue4
ueexbAkUEW7KoGhKb8CAOSz0phPX+BrS8NhzIOKaP16Zt/SC20eEzSBXeyAQZl7VRR6auKiToG8P
5ye3ybZ2ZE1n+9zn435jQV3+ZNUomL1CbCZt/VQxji/t2RaAYXvkjOJ5XMreV5rQ9ieJQ0TNoUXv
s2Aennm/590UPmeM+cUjIlyypFw0L1k47bKqn5n5C3PUwQFaOuSiRG84ledDi/RjHhR8zciPTxix
AXODIeTK6+WgZqHqDcMrLgnlI7DK1mFS+yAej4SFqXxV5YmJrzbKQjt9cL3O6Q0TAskrR1O55hGG
A0QGcrEqZda8SMXDALJlrpspsYzcXBWsnXCqjKl4bF+t8qGh3ZHXSPypSg0QNc/avrNPV2uGh5tb
nCbYltOvErtJHqdlPipGIhu21LI3aeGEo5L7kK612PvLGt5JhqIA7hprkde3PKhzpJBmOqZfNtYv
oohbYioa8QEZrhhW4xtTBhPofK1DE3EPiMXYcdXYSzk7AbHbl/94wQ+w1m4wMNpdmzHMcUUshdhM
L7p0WQNyBoxSSv2PgEQLpX3y0lAu3Rtr46/mzDhSuy+5/ywNzaK192qkSTd2GJV51kIOeW6fdG1c
GZWmmwgaPpMm8qj9VVZnTm0b+bOl4RN3uxXIConyCMwvINw7Pgk29tnW3DwsG+St+vNh4nHKKV27
0b77Rn3VRnaqwKEAB/ISH4D7EjYMslu35Dl2GSAgc1k+XNY7UnAZ8NJ5hPD9xi0dBfB6uMnwqAGp
oe/YjPFZpIIkDpVJpq7xuJSXuqTFQgxhDWZcUgWvaiI0+e4Fhdzl4GbtwnexhnZr2wFJa06xelT4
9nc0GJJOTu0QmlVd6/IcKcpOC+B5bI/cWa23tlQgdyWbzO9/4KLIPfiJtT0Uss7U3ifB6jxyrIwW
YaZhVFeDlmGcEewrMBdxrfqUmLxgXdWtDlL+J2UaqZcwqz2clcA8t1/WQ9nfmrzi6rbrbSDrGB3p
WSsdWd6ZLi2PocQcO/609JTOhDe4hNz7ntY6i+o1HLmE4603Mel0Ok9Snh63RizzAVROIbFDJ4wo
ehxD9uMq9cl2v1SDGg8crQgd1PkDhEu0i8tFnBUIPN0Zys5UxQjKX1xzebfy8r8543YlX2eeU34S
gBiwjRunrXNjOs4jcXFZ11c63Z0vcp/QGzshsESu7mf4Tay38i9JC9mEefPNhENCOkdGyojEgIe1
b7Hm469KdsdeZntl6eEuiEPXkcZv1hRlPvwrDe52SGXs/e5QsXKgN9iPYv4xqV4xd92ZJWJgvNb/
PEhjL6PJkICfwf69I721o0Stcmmm96Il2aNeieJFysadqwWACh/UhRojqIXJwmoQ6r8WUL2jrPjR
PkP9rB4niT73iupfO2gR49VXgvQHN2GIAYF5Sf0g2fstXakAZYLOrANqc978X3clXOGSJrhs0cWm
gO5pi4IeMOq3UiOhoxqaDIx6nDcwmRqd4H13qkhzTH3NwiBNfncJEmm5O2xtqehGZgxKJej6u+67
uKoO3XSP14OyJ8I9mGw58WRjwA6YhxtUpNtUZvWppPVGqKJUXvPCtyWFbOZZ/OLzucWI/LtXnUte
WUPvSMMN+JhC9+w5ZWlvt4lLCr4PMuFO5bFP3HJFjFsyUDvurCOwo+K6wQjyGMtrWpdJC2XxTFl1
JiuWuN8ZD6hW8OuY52+iOqJ6HcbVaCpctWecjdn+zseQD7Cd07KMpjyXeiuOw7bqmszWyiLrwHtJ
3rDcDmMp60eDMuzHWdPg6PDE8Tyn03wDD82As87Y3y/q6XJbu+rW+QCTMH4e49PYI+i9SD4H0xcn
czDpL5D4Vt6kcnpUAtp6BanDeBs46AcpsMd/y2O5HY8X8UPYIQJ54Is35N9GyDFVTf4WaXIBgCid
dAnX6RbLgoP+ffeCX1LQeDLhd07OAVaYnDCM+sFb6Q36vSUJ5s79qECDTuPgxwUOplNSPcJqdsja
rkLhabujPMLmqSIy83S1J26Buu7Cq8ZzSBQ8jXBPjUVDUig9iaF6XVviaHwFcrRUrBDWzCL17NoS
cPJXxHxfXRkn3EXA0llWjkjtF52RgMbxPRYEzpEo1JO6mzrT2ZrrCm54S0+1DmTzfgAb8WndyoD9
FoeGTUpBIxn57PX/V0F0lDo22viOemlya6ZxzW5zFHeRsjTMPpZ8UZiaOChyqjzlOtCH5xJOsGF1
38BUiuUTtxue7t6W61yu61M6zXjpEHpdvyJ1DQObvkZZPhqm0P8gXIJYFluCXjOxiIrVxuD9aNSt
6w4Xy/F+b2Ehwa709XVr0TxJlrmZFFSpFPaTkwrN7yIeXmF7B5awrNzTTEhHI1bu8vTlwrHYjBS3
ekX+FoTr4ghFZUkbWlkSm/LSPE9Gd+JDudS5pdE6gGT0pbv5+aGU5NNh+NVLDLA0t6mkUczmwj7p
qiRvsAkWYjYvzt7qWTv5GNhtrT3pujTAjxkfgrNZJ7C56lRKcO4mbkVT1AkRyBNVGRtCwtPdzqgj
Nhv4fscxyalV3H787DLagAmmj7oqL4B+yNc7RRZsRKpKzlOjUYcqDQrMD0xHwTCmgzfzKgQc0BgM
0YmcEa67Je01RhH4YbY7xqNnxFCQmBinndwJog25NEm2dbK/1ud/7vFdkR71P6y3zo3fH3mCSoli
UJ0/r5zcNY1w7iqNANWdPHqIvZRCFSFivUlqu/a9d0ycIFogqVrs4HcCUNcT75gMMy5in9x5VSIC
fKBsUNVMHyDc0j/lqnilph6eCocchjnlppbDMTqlW/p5y3y1Tj/3II0j9ajSpItFeB20bB90+f59
nPVkc2XCi1coEVrtIQU9HyPWeum/D1cTzAaqB50DdSMje0a7zg8WxPMn6yGKPigQw9z7IGMwi7Gi
Sz/MgbqN+snLrICQZqfk1Z+zQPGkT6j34lvsw2k+wxONOU6ZeZ09dEGh39+Yol2/prNZLDCAYAWI
vjv47PJAEE1ghfWipmgUIq4CexbRr6iekOd2HYO5hC1IVrZ+kP8p9dTj2GTpzsry2kWdSL9R5OmY
BfirRihxNdIqlc0yb5uadie98XchlvdwmWq8+1dFMGHNgEOimNnZkGc1MAjYYY6P3ogIx6P/wiQ+
zNSr3pZ/P6IwzS9V8sEcQAhKjBoCUPj8uQr893rks1ZPDnCKvybZD3BJT0ajV7tuVVhzfpZDOfQ0
3PkYBqe0eohQ5WZSRYL/Y8I8IQw/sm6luYVgpWaRIHYqXvZJdOETEZrQlDsNt9HW+zKGY5FqLau2
m2Gg8Kdf13DaonUg4hcU94eocVTGggx0YcckklzTdGC6dByMq0N4Y15ynD3eML0XgzRmvW0bxdBH
CpyhOD6DCeaqC+n3DuqDyNWkT7PVlwD86tI99fUB/FQ8yfHoeXTT8eC2jrOqk1lnsL0CjlXYiTx3
f+PBYUoUsVeq3Q1xTMFK/O7fm7XNeyDDLoD4JKvas2SPmN+C9a5kdtsPDlmZ0Jfu4RUV2qIHTK/s
Pmyy0D3WCP61vgmk1zAguZhNU8nvDMRwsVIJaZfsLVWO/ot6niqrqoIg+9w69haI3PhPOLZ0nb3a
qjeqolDZFNoog3H0ySzwhUdTfNliQxIINdxUrm9Cgdqpr+enAFR0tYrFFjTZqRO2DGqLlvJ6lvY5
q5pHerB0P7WYDdjSeiU16sy0I+1f3ITDyElN7gxduCpjIhDUEyjA5ua/muIoP23IRtHfakH5oQtC
lPJ3IEA4/zQmprZLzN+7op9vZMQXiM5ofAD9UACa5mzr8xjQdkKuR63P5TWJxWDUN3I+Ok4u1aKn
fX7U+I5zPpswojmmCb000p/uw9gmJ7Y1T2jvrhPd1S8BZWje2ioglwVH90tMOzcLWmx3LuieKEe0
paRUqL4xRPyGTZqWU0BF8bO30R2LRH3adIunKHByt7N1I1WIScxg5ijqtDoNgthRh58v1kjGspMc
Zt8yjbPmWA7opr2NTTp3v6qrA+qYHIBgdCxGsc8A1t6Ralv5DG4BNRl7vNlUvCwwcVGU/vRZNdcv
9z07w2Fwpy3SLSs9rG6KqP4IRw32OX/yW37MwOBHiBu7b3SCQjA2GKP1914NdY5CVgu3QVIK40uE
MuPe3hG5KNeGBQXSrYK6VrKTAqSYSl3A4d3HteIJaQMRMhI3VAdJyZLHY6l2krd3I8cfcR+Gavhk
S48L6/zJ1ampB8+RnItmWyPVx69IskLkUIIgltIKoxgUNMx0J2CkiFk/yoirU2w8zzKBY6uhaArz
L7R/H5aFrHlUS9RTbR21NP9mYnCXsqG+PfmJbF006Z4KbECF8TVW7JN5RTpZML8Lk6097Nl7VGZC
A92LDRKwJJ3GoiEGBhK1dfgpq5XsTuRZHcNVqaz2tQmaoDyaqjJHFnrJ/uqa7tI22q8/FNno/dO4
VvPCEE1C2o3yMFY3O/HT7Op9kox+9zPe6A8+GY2+iTSf7yQZOtYzbvspSJrDFUrXUAFJcHelLi0j
i4a7k875nVZdPNjInoouyTjh7cdxgmvAqkuhMs4dLvd+7BMoJ7ghBhMkHDsHTWIFfE6vsI5zmDFr
9rFHvF64vLd+R/+8WZBS8pCMbIa8l7HwPYKAswRZK6WXGkEuS3Muolcy6VohS9r2f/EmmhOl8D+V
oEwnBhamnsRqZ5hnsVdjVdPMdcphI0CdI3hs/VgAH7bDvJJdOZQZHocrANKQtAkrCGIqUfiNt3Kc
uTgYjXJt0GN53+x7svr9QyHwnu1BKO4ypO/9s94y9XdDz/F+nLGUZH80VPMVqE+GJNSp531DEl1e
TIO/BvSdaY1o82BPtN/cp+rrmuoxHAxf85EsaLTKz9odTU3xOmQPVPvR2RemXR+XFHDXTX9kJtrK
CM9zyEkpuvrlwZTmVQ0H/HltV5KY9fj2tK/zi83uqcfgphYdpPVsgaPGFgB5fB796fSXA65rGNU9
Q57qzAcUZlK3yf2/9j3++5FvSJDo2xmDQREtbMtJo7qaByRH6wUCaaJ5RqnJdHM9s1hzQrUhiD6g
CzAhQm1eiANsUN9nMhCaor0CxNVw9VmisdQH932oac6gEe/LQvhDDMg7OgDl6iXYAzo9nLNzWsk7
rhdnuPbrZrkIM9TWAcda4j5EWAEbV73yq6KOPfy1tajb4X396vvNjrLeD8CQI9W26cDlfjCHUOyv
ql/kQYnkp+15TgQLYVmP/QwD38XZZZy2IDI9jmQ+Gb+9hgQm1rrRsWkI7Q2zePLzTQd3+5e0utx5
tStfmxtmR60DbhhS5Tcw6AeeBEovpnJ609sxmhY89MbOsK6mvAZ3vLhtpvtwNLBArWsb7fWWhNQZ
fCycZF84a1ZxHbtL31NGm5rMyZt4G7Enq3Ymz5h0vuiccvUgppk2C4Zdj4cUNp+gHA3z5VRk2H+J
2m0eqrRBbp6YerujAiKwGWdx1eapdIBrHBV/3LtE/RrP3Of86rRh/TQpfIAmF7wT2wP1MoENvXPl
XQKFmqYacLE02g62CswTe23skLllw5r+COWC7l1SOx2IN1Wwhfx+4UmOEmNfdaQDmuUmzcMEAiUP
XU3QjVC2TJlwH2EAuZnvJfW+RWbMuqUUG7TzzJ6BlMrC4YYPkwAm4YcVRLHDZ0malxhvyaBSERMS
DymWbZ7VfGR1yxtuXi9Q80eYliz5IbfzVgYWmaizWZqnubDxP275iNjslrJ3VSqwMLCUqoe1rU2G
hYBcplHnXcPIFYylme/k/H0bCt2sotOBXIUVqKccDU8RdMS6mb+x1xYZkcY4BrQ9M/lh1wqxZzol
PaPU+TTkqs4OtNuzHRQEc6ztSP6gEMNiSV8oWTUChwWE3QVnnVuuh6N8yiBC4o4tLVdUQsV1CeBs
SuUA+hO3YgQhGsI0sDsP/GIJYRGMdqtOna+vAN9HYnhivbP2jBcFxY+sFkNUoQfA9Q/mJDrL+3ou
FL+KlFbQdH5LqU7x32iT8ykDRSVuGwkxDmbjqT/3RkXjMaUGGJUza09dPX6YnhXW9E3jg4pqSMZt
0U5OvmCeU2+znbQxDfYEAfzuVdWDX1D1HEA32hkQ8vs9sR4Qk+px/YQo6DyUUatxtWocPEmhb17/
O1km+0lce01PM3iEaBVHNYZdUaDI2KFzVBFw6vTWcbivWuELw7fX8s5hleP+ioNMoxz7cbfYwgvb
pa1PCmnGv/FTjdS8u9YYhDt3uakjYnjE03VMjEJM2ksWNc6aVYFfnSLsdR8Tk0BS8MZnG//NWw3t
KSVBRTmzhn1TbzsAZy26ckawRwpJAGiC6yYfo9o4CMq5pSAiUzyU8qUINGZhV2ZLbB6lzvmLbBdl
e8qOjHbj44AUV09eGFJEupoqTp4CUzRQXRH/IQP2XON/hMhq/hAmf4zKgP/U1CFy3gu9lK0UFOqo
pxTiO6Nc4fZD83KgHIkCb816eCBBSBV+jnCo+rZS4Sl3Gb3K75I/X4FZfITZCuHNjMGSPo1kokTW
v6QOBH+EjQqq9jKYboJlopQ73OJL6B9ffs2dHG778uoNBtKbcsS+c988aFiCECpXrkOK4QVKfT4r
Lju8ug10ggwVxhwAnVRoOp4oXyInDwAdULdPwmWaGknVy+SQvklGT56cWIQPkQYoujMMyuw0ROBt
5CRIUzSo5Ae13nTHGm1noc7x/sEVi930EymYecUNr9+40ZIzEBYDciNXBp8Y2Os+c1h8rxwHV9rO
MJKIbWPbmKsHJdjKfdQ9pfvIX6+R2+87+bBzQG1tTzyB9rF5gLF2aRYERxQOWxet1gqGVRV57Aau
dbeuGMSI4iTe+mfwU7mmBP+MgEEDLgLaBVlMFeQ6xKZFddftVH6lrCV2ibrIpK9kwHheEzAnElyI
xvq4SBkWK/0sKCEwzpVkuwsglwsCRRXsFZTG7ZiOlM3Q6sf2MzNSSguiA9z+VkBtRUU/noJMasJN
Sbs9MVobXD/J16bZi4z+9GIfuGyVAIcIVfhpcDHT1p3CZ6zoSCirbs/+L2gT7Mmjl0/p9sffvAUz
XEyB0GqjKHoD6iX98XiN/OVoFwS2dn3Jfu90efgtw9n8wrS07MQH8enVTYGKEyI3TM0z3ZrKZzYe
aw/CRf7ijMaToFJ9LpCH5YTTd9qG+/55s0khciwsLMliEUoYhROgUB4f9me36gbI2SXGeF1w0+d0
KUz72x6KrnKQDGz9AQf6QeryDhUqnfsORJdxRiXJ96S3l6C8UB6B4HLUEY/S/mew/arCYRulGtJN
dSZiIQGwuaeNUDaGHkQiVk16mU6yhuU0NavE04HiCOtedEYOiHIP2bpVL2c5GWx4LdqHyDRIUi3J
OX4N9mvoFkdbyvIJEkzKy1cfyZatBXqYpM6caq8LX1qA43HPEOSwrCrCTZ4U40GutzPdbTKYK7RA
pfV9n1E1mqIOL7tgh5x6wDqKx/tRfw58TnWGlkz+i1pbgLIt/WPiomufUveYl2TcdP7/FH8oirkC
G1lDD4LHRw+SU/7DkZnIWB/r5qc2KcOREDJ5m9L4r5sg6UcNRyO1cL0lFeWhlUoDBoLuaqyFXZz/
CjRTwdXKWi1b0OpOoxan2yXWCPBmgKBARuDEJJs71xBhBUPzVu4QI7pbc2im7OR5lDtm+8JykXig
a1Ry9fLVJ/aPPdFBrLU2b7hTwPlEfL/1pB6f/l0WSOtlpaxmep2p25XA6KtFXQIhUIT6/K0TkO8H
HOv6/04F7JWp7SHJsRxw+iPVlFnV7LtBPCGxnpKnkCd6OZk8WwCiygis/beeI7WY75XJnuGKSF7T
7ueYQjNZdZ2McPtzv5L46XImOsGW29FV99YsG01nISOZBjZZ2Fdf5WVxbcejAb/TyapBaGj+6TpZ
NYYVIhl96mVoZt5NzludyTpFQNKxr6xhQLQJAb4+khlFbsw60lJzLvXYHklXEzie/P5gGj/lHNWX
6ot7AXltsm9In6GmTx48zWnU0ureuBtQwEi+guozNk9/5pgBn2WqrACev6R+DnDz4CSiodX+ZdTW
4NoY2jLTYm0uf7ApnFe4Q5JIdktYYRUrTyrXsd1jFIl3bKRgp500EETlp2Cj81/xKoEjMQTKOuR2
Lvq/FowFY084EyR2hDtOs2L+GGhwCKybZi1nF7JR0JCH7VC/nueZWlpEEJJANEee5yqQcj1IKzD7
h3fV4F9cyLW6x5fSHp1tSeD71DKsqfCrAO30hi7ErcOsQKH+sgWjKup4LCYkEG6Ys/sMbjMehGvn
2nvy1IkezagzYJhgtFPf3BD/zJIktblji5RWMsLMSAy25JyA1t+n1bemh7n2kMmxVknFcjAuzviF
q1pHRxYh0lbkiW+4YbCMsR26xXO9wyGV2UN4p8dXcg/bCcpruVF70c+YDcQOA/6LvJfO7pAON4NJ
rqb8pnQVDxMN4WfnajeJU4acggFgMP0/KSa/gyzGOJy5ECrJa/04CtERKJBczbDvKVQdRO6I5hiP
uC1E3zoSd0lNi0PQugHd3h3hFjThjji1pdgaA/gz5PmdnBwU+QcRorYJ/v7Gcn1YlOHdlpGCsVsO
wxrKry9b/sWZqN6PN4ySQ/JHq08i/MFlOA9M7ldFv36i+LeYm41f48UoWiYHraIbDVeepY0Ed2OG
MBrted6P5UdAUs3xLDkBH4VMGSdlopCoDH6ChFm9r39aCnZNj6weSRXfjrYz7bmgj2EKpYAZudJC
pu6IdQKhVCRdvgF3YDpKIG6oUbtxqnDL7gXLAGrXBo1m/Jf3lP7tSIx08HgLpJ+7YzFrwZBDg1cC
8w3r3w/Mtd5yduLkyjMH2cDy7pfcdtzE/sW5g6hhoz43Yseh6tNHvESdJQMV1n9SKNkkGEUMDQLm
CldrqXlwfulz3yVe5dqgKtdME3uTJNsO11Oe2AyLGCn7Mdw30Glz/EckZHNX7Jn6NSlvudjS6U66
mM2VRk2e8+5YT3g8POH5K6KwtlULF7civsJfiu60wGR8rNT9VPDEe3PE70eJcdfE8yHZPznnBWZS
7lCR+oGQP8YiGRoG0K8sNrhKhpiwN5GbOJXYh5uUusdZv3UVmoqRV0bO8DTfUBUFHPcSynjDullZ
PUJHcC3jir/N7/GEIK1RbAY4NVJ9zUbxnnECycpMbmvAsgiXa9EHleQqil/Wfs2bUAeeh2RARsM+
8xk3bfGMbFX7wMHQZbvGpyP/eyV+ZvwlEbuRvkWf/Kt+LrFeZkZ0tmUArYVXoq9QtXv6I0DSz4I8
Mr5txKaiWcUG21Ao3//20OB5TDxA2og8QaWvVsnj+8SnnfYmpsVH8FVD8xuwBCqLbZPuBwjJxEVL
kD5Ssj36YuC+kIaCqALPWq1Putvdz2cdtqRPBzQWKWiRBkNLp4JHf151pqRNyYuX3TlN5ysOZnUe
Ir7wQfUOyYDuLjgMl4y8N1KyVwGBgmgjJy2qeyooCGAYQgFCCKS1fYMxv1njMqT2FI3EQfMGMGJl
kn6YubociZwO9dW7uj6IpXJDsqiAlTvijKvSk5WMvMB0Pss1HDbOj7SukTsz58z+/M3ulmaa7LO5
vRLtRzqrO0zcp70nL2HrGeODvWNXOs+RoYBX+2W1pjv8PzryY/xEWvte+WFOkhVdJd8CsnQdWCQl
bENolGT8Z/BuJa0d5ATC7hUCxU3e6psDZP40y9rsTYBByU81EbU0Rm3MxkCBRJNef8oSk4+kDS2G
VkeYySBVvGh5f4/LveWc5SHYNxlqpE2Qc83Jflp8o+ZTKnXhscQtaR8FTchyHblcepXjcx+AUBiH
B+xfab1+6UA+SyOY4HBJCDHtuKgxHt9dGhP1gIH1kAsy01cJj4N5WueRuPlvyjPFbc3olM7MBy2c
OePIKt9KpL+e+ANRb9biW7sRtkLUeowNM+cqU9OnlnexVMWcfmo993257QXxE5Yl24cn7mBYUFHz
A6C/UYkcnMWiaWEAkrRc/bmSWZcLNmRW6i9Ikc/VyqhITd9La64jRg0uTdKo4s/Fyz+tI5LnE9yX
d11gAn9d4naSPjgFV4dIgnWO/nmFZi0FRf9QZdy43s2ApxypyXyGtKfNgwmkAasZMhwbMnwFN17j
RVda2vWQhR17Kck6XYCrQFFJYwQXqndQJpT4JHhmTkm7zL5AC63+cQGE7OnWHgKM9XlDTrxiHRaB
9IoSXwQKVAHpGkr3balThk2WVB2aPQF9rDDsg3yPFpO0Zcd7oSRi1Wu51SsV5wiG6XuzZYRha/u0
sLJtc0nEGCVw04pMJRmcHNHRT9VJKlcdcd7neocuLlU6UP0wiAicORbETsHiZLEQCDndNEuWZJYp
7mcFyKk58KoQ84zlASamediinZUv611K8MYdyXPcaVxG5I88vYvAWBZKSRquo2Ef8m2zcA5iClhW
ZHdNiPt9vJI+1lDnXhys0zhJYeYwxsceOflFZY2b/cphiblBkw22u6inSlnu/tALf5s8Q7YLqTEr
Vyn8sWqadjXJYDWhewcpm52xh4ezolR1YtHCqFzSxBYoXzj/h9L7MuhfZaawPtEdh4ZNk3Fm/LbI
q9dEh2+BqDyV+RnN+19LH8IMk02H6HyN/Lv1g+E7N5V6KhV2i4g4t8zx2j/Lw3E1jp5da+9uDUUR
tvn/xqYjRRi03p/kNquengZrTLKFYyTuhid0WRzXsRURE//ICgQctyO6F0cMqRMCkhM/QBSyFnjX
khrPJSOlMJLRumyjki/zzkbZ2PEjASho2Vt5ypLRdvTLNglVIkdT/NnWUBiHb8ogpwyDAdTBOjbE
fhWmwlB0U8G+bySSVieOrER+jWz92UuEsaaRYZAco97okIfRCQdpmBJ40Kfrc2hjG4XOxjDIF1Ks
c5sXs8lXUkFQXR1UYfvy08pc9Nr3T9H/J/T/RASiYPCsnjlN/ladhHwRRbGhoLDNf+yhbqcKTi9c
9xsMTo8W00UGOyxZ/YmF/o+xePG2HdAr4i0BKDNHQtehXEuM+DDn7W77WvbFbivZih4P8RkahB1N
RBB7jPxBr84RVKi6jADDu5ufYuoVUqu3WpXRlVTq9rqRgOz7zH2VJjtkT6WPFm6cNFOFSJmP55W8
CuSnmJpbJXEMnSmlFdT0Pcda+7IM+/WPvOksi9HrRqEs+YzfP6JC4UTpZhfXG/E0f6Uove3Qza0o
x2GyH7AmqPRWjUHTS35EiyUEH/736s5N+uFfF++uofXE1FcEza16biGf+8EAs+Dwk6RvAIFh75rE
tIvHfMHboXCgZZBsfiZ1FhJU29wQRUnEaqcuD+cA1GOKdpYA8yf38Gz4RL0WWGcc6+UI7gFbkkeh
mOmJi72SlfPg55shYxx3pgnrkHgzADcy9Sg+YNmlxVTD/ZVR3kJLwBIw6q9EmH2z7ZxAulIYdjD1
Pdi5QhpUcknlg2q83yeRTGNncGVDyu0nvyJlIeGQxnQmt0sUxUMIWMiLWOJyUU8UjwgHJ0qvAs72
YpP38HE1ONOUTiCS/oGqd1zUVGpOlYpCwgRxt3KZ++PovAiItbV809Dl+ShdQNRm1+UYjBRYpZVJ
on6J1lI6Ge1WzjtRiGTKGPDlIL8HpsvfhZSy3VaW2jH90EHsf/HaivMlruE0TOzvm2/eV0FdZccb
FE3zMJYWOES7XKrPodtjuiVnGsyqAue3EeOPt9NWGBkeslDbRfgYM3zI03XiBPOB52bYVz+d+48q
EmnUV8M0NzdFcB7lPYU/2y/+xWIyBMOUyLCtb+KrRLXvHpw4z/q8n2lvTcvh/kg0KJatPXAM6eLk
KFR9HgeEPVtiHsBrBSIBoz6jNHNMEVI6P59Lik15RfAMWqDw9rIR6AfDsvoQZ6BRyN51ALBUWyZI
3B/j1E3HYZf3P90Aj5jQEdt1aKXxEU6yy5YqakK1rK1q+1rdxCN8L/K4KYG4rABhe2rbx+AIEprw
P0htTKqNW+SeKNMLgCbF+RQiwgxsvAkow+cVTL3tXAmML43p0H2hKPI2DcepUwP9lsWjilwSGemB
7+WBnpV7flInvg5iotDacYymG0SqJWpGIPjtRW6GSOHnAG9vMDAqc1S/SEGyc/MGgsCTR637vVPX
QCARJ/0XGBsStRbpFuac0LTDYfC/GkI6K6dTW5Jb4AWJ4bAhdCr7nvSa3jPCRUciKD2hhX52Tp52
UEJOvmsERhcJFta4Bal3ylhXOK50zdxbcuT82XVw+C7fMXBFLStABS3ahdj429LH31zF3KnvwlO0
eId8Iste/1Ng05q6hZGy/wj9Q+BK/HHUreGPcLiHgNbyS3KP97pOiQJUGex9tTRdF/RFF7lETBjv
8IVK0USCKT5/5jjblvpC/ra2KT31C8MSLgNofq0dI/a1J30f/SrRzVlORDdOv7wbrCUbjqoIpmvS
kd/fBDmPXmWqVCve80u6xg2U0PMlBRO2D8T0whunWCPXELP/cd9lnx3TF406uzaAyf/xTW0jqamA
wxqol9IoTSbjgVI/kRFXFPVdas/zgwp3rDXpkq44+tQ7AvlbMEWbAibox872ONDY4qJX2z96KnLD
l+LvwHJVzH7Fuecb99bhneZPBw1GwyXMLucH+074WnNj21knBO51EerXjDzlFPDjXmxra+VxBkDZ
x+5LIEKRu9kFu5V0yTf3VS83JAtwPd/Sgj7vqvKRy5a7UJCaGcmtxhfN/Hkj/nGf9Q86NkgPOC8s
ZoFhOvW/BRc3b4IVeS8K/CB476Z/glRlaCN2u8k8KyytwhvhQT/lxGpJcQy7GyWMzXtSUXdUTKme
pUC0/qxSnAhsIsb660yZ1hku6zZMrX3urx090xQHYCLqf0YT7526l+5kP7EtchnWaBhNolHrxbp9
U+d1ptY2l/B5n5N5h2/Yb7IWi2/d0Wg8qbIrnYzy5PgM9Pk2IsOW6yz/1++swaM3JX/g3Q4etwEG
naQMtx6lasdQ6jsjcBfLqZeQng+WFMi25lTpDVVDz/RBW8fz0B7DSQdVSUbdKNDJUn+Ruve8sNNI
pFCAYwR7tNo5IV5yaEQu1o8USMhjnV/+AqPcMtI0/oZfO2so1SFuIXoi0ln6uB/FZ1fmomGOHaZn
fpb9CQ/L3h8Aa9QHJDcj2hIrj406KiLQ6i4fybfdgosMQiQPPaTvzavZX84QaZUQ3TX6DRi1bC62
A45nitcN04hQsQxNjfcfmW9kOny223rSKGIIk1C5JtOq/n8vtkD17CiqwBeiNJxOuSMG2EoxcxcU
Xjc5v1dZVf+DfC6uLcfLJaUu9jYCu9/b4gqC1TmD4Ii7sFlGRxMP4B6yGwOofeK95JpSLmBn9EG/
SGg89bFuH+WsjHskQIRxChAJkJTLXdoTKrj1ShV0Qns+kfhFaKcdLXuVYHUOOPqLhRcWCa5hJygQ
8edn6bcN74eIqxQfv4ZfwrLKH2lPk+WT6NBH6VeJssCobPBuk4NvoXrkO6jHC2b2C6UakFn9H5N1
KizhxhFMSyYgoE+HOmMQjJedEfeTWS1V5v36d4ciZvu6YFWOcRi+tkKNfymyWoZ1hIndLejlbl4e
Cc//AKrSVEHo3jELdDdpLiLsrq4ngYKUSYv76q8tmf2K7mUjSXAs+J6ChdOZ8S5yNlyD10kU2nrt
AW/ZJA5dcve/PwXfoUKf70W7iZUyOTXdeoAoF7IbSw2mQl3dEuZPHbvZfHcPn1Ml45fPaoZW7Tub
k1rMSH5B/wibx43zCTq/ECwLO3GXg2lWGv166UyvC/7YKGCmTE0JyUdoa9HQ2YlPtTuS+e8ngk7w
qCd7ynC0jDdqIf4Pp6nktBYkbgv39YMrQSEsnC9ojf8c262KsTfuY5LuyJio6zSTPtcEhrXzYdIP
2iDXXtllm0Ux5mzdCu24w/liYgV7vGvKInZvdvk/jzpFoa39hjA+qedwrPnc0Ee1DzyQhAoPFCt0
jclWhJ9xTYFxB1TkAoPoXO/5mng88Vx+7P8ewfWGmX+DKFLhUUwcptMXeDdw8zNwMnqNx6mLwBGL
VJDSToPdC5fcGUuGCRmWE9Pv9T44fgYk2eLkGfuO6Z7Zj159L+efd9FIkhZOYN3EKCF/oclbNc02
lnukUdAogLzFa6QHvsBPmqxsGUXXkfARMX1hB17jfaBYuWv3ZRjifgbcnfhC1tQOEIvKP/9zn/Ag
9pFt0V8LDTVVv7z0diGAdi2TKzSX7x1Opl3IZrx+A+QRgRPDtYCu5OzV8nLOZbv5xa8J+psq3nXT
pjIKA+X9Pk1tWd7XgMxNj90bY+fulDQNEJlX3j2Yx/b5MwECUnyRNSCZY3zev8mfRBO6Yh71lceR
Nj9c3n60orr9S4ntEb18LnlbxJIVMmKWzUCkkQlnxLw2fUMfRpjbdm7m/ccD56KEoAnQPrLprNPu
WKLEcIPq/eH4Cap0dKF+6P8RyLykYPlPxvzoqnkZBF6+jTb5WU5FgWHuGHevhwwxkUgepCs4FN5T
fgzR5NydoEIYMEb60PuxsQjzHrpNKoO3NC3SLtJ0gV4gTNmaHXxKVFv00TlcE1cYVuqIF1PZLhT5
RNyADaAfgpieOz/fnBEFyVXK2iCQAA0oZgxunx+agsYwbfowhVHQdTQShDjHHqMEkd5Fg0gp9dX6
bdsmBZ+oXQWmV5F7QeTPNjFqSoJkuRNAe0ZTHhVjhy5WJRucxXuS47tk+kpx3v9lQDkStHq5a7F4
U4/qnYqR/fWqpgkSeIunyUxVKfMdFXGapItrKHvyJo0x58GqI+YD0vL9z91ms1f+Hz5fmDwSJhX1
sb8LAO8ATqBcJcMx0yjf1PHP9xh2tZ/baW8P+bebM0XCAKCSiWMGPMX74byKb5HrDjjrGYk6upxd
hHHrzF7o4vigRN72+QgNnGgWOO+rb0U+f8vhpQ2LzEsNh/LA7OyBsOWLtM7EGV5M9eLsnZTofKv/
c+Fd87sZG5Fof8RopBrQw4nq7Hd1PvlA6958MFxR7sL1PXfTAqRfygXOXpLJYaCzsqOnv89LUJUv
DYLxUuhmYC8+ISdIf+at014j6CIzKtFo9UaqjoQSy/1C95JbZc0MSAXujg1nOAjJWILTDd9K3OZc
7HYKejqVEKurBEsQAmCJ/mxFfBkdqm/djZaaAY0Cg6JMykVvo87+QoQTJYMscEGueKAh4Ptzi7nX
zs8bU8MoS9peX4JWa45qDBpSCSr+JaxYVyE6+y1Zt+tZ+gafPtu3V2r6R+CYRUTqmp0rS3HImCU+
A3sdOyFbrjKGYRKayix9V/23IwRrtJORyoeRPwe5i/XFvhLnMBLrd+i2PHxrqcFQ4fFiYeSiElTk
8Ens6MA8q7cmDVI6r+TbTNk7i1h6xNHLqrTSA3pK4xGM39gxLcgH5zFJI9vXHnMt/fDb60R23oNZ
AyLoxGKwe5BTa5hwElH5GJgVEcgAXP7W5XWhRjYg4ExL91vbl7WifXE/DGAascvXO+oGtSQI5iiE
XgsmeztraQT7+FGDVR6XGL2IJl8ZbCORHK0cvms4Pd2FY/Qh6iRDKsqQr+o68NtcqOZb9zhAeURf
5iuzYYgwEO+T16dqJs8df8TGizDFK6DTwHwTgyAxdiVn+roF82ml/B/zjd3QdoXo4Ohd+sLwyXVw
QD5CeHklTBBna0gPJTvq0i5nJKVMWFO0Z3RY7ks6nrBoO+qfOVbkgd6DR13havFTb2QEeHBYsyw5
BkqEau+ZQIed7w0YBln6j0IiaqdA2w3AxMzmm7W/7vtDt2V1n26kfldi0G7lZT39OJwKu3a49pQm
N9NYyjVHyHrzWjto7SyyRM5SOPGUakhlB2Q1mt5cWct++nqP6hMP4PcckdKzVKO1ZyMpZORjq9Tu
63VCCPpjv/RUvAPFBw1YqzlgEHPI8bkHzdErjVrs9sExQIzpU1AGKdnfn8MVDrROCcKGgnsFP3a5
H+FXYQLgk+1o/Q/P1fQPKq/zR0QOe15WqFLg3tHX3LVP5oaIZiI/39Ok99SqsbabX2i7V1uZG08y
LSd5bS9t0Tn6KKy7jgS34LKPvasouq3REj1zzGI0FP+yRSwGO+XEBQOQW2+8AY4ZgSHzvvI0jZFZ
rmSw97YleetrSLH2VXvq+Se76rTtPXJbEtHdLOxQRQ5/ubG8ZsHlTh5bfP3rnm4EXYUDqbHe5XIz
udIPINYCupwR9aLMoEnEanYZASN2TR3nmctT5u8SWsdNWTOQs/E4oOseNgAYoCyvBkmwj6uCw7Q2
cDJ6tVk+2bLJL48yuFElbiUDQOUAjontyM2jSs1kH+6GkVzv34SUA1OlsdNTj5T1H9sFnTt2VUuh
+kWM7ibkPoa3CzN4ORlcM5bWmphGuap0bpXD/rfrxeNFL6ayImEmQWVa2Slxw00ZxwV6xByWO5Bg
YkjPzM3Ysr69HNjf7WC5UosnbUXgrc8x0MjMNl/khusFdtNKHiSEahz3ngJbxWtjSKtyKiR5NmW7
i8NYAURGgJWZ1Ah/sop5K1kkbslmkNrAw6E3Qj7KMABH/SlEORqWKS6PkF3jH6BgsMcxR6DvdMVd
otKUy8BPfxCbyArw0o1sR65Fg4H4jnn/w3nNl4PgTtsR7FVc3VlXiCYlrGONP5numYREYTFRyQ69
F6kSkhRd3+f75CV9y1arYHcEL0MPjI8jscEUXKT/pHj1r732otiKY6A9dZI+CpP69QKJ0TSntUMA
YITwO3XzIdBamFsI3w38+JDLh7qIHxCNp//2xnGdDcyMxerbi21MsX/l35G5A1mwxlp8KykGa0Do
/Sges1Gy7+ehHiQPaKNDeFdGYmuWpSbkHWxkBZ9igdAT+liEoN3ixvHH009Nz/yauVqXrHCvYLKn
N33qZ8ipj/UwwVkcm3budKVl0dUyrUVOUfy8mHM4nTzXSxHPNcR3ui822dHxdhkEoY4lLdGv2Dkb
OZ1jsq0Z2aAUGoYVN9IyzxQUtStWPbcn3Y1OuyEd0JOkMec54nzxU6wMU1nKe74rQ7vSOBqgGxuj
uCZSg1IWQKyHOozpZz3ZivRuR2WnV7AupmHaPJhmmmk2eoU0BYI+g1cXPNg/c5FlyFpJm006xXIw
SLj16aYs5I6/PINQ5UGpw09k6Ug8nDULk5jX4F1+PzQHNndxIABbErXkxW7eTZhrhAxmEhg8re2R
i/9731h423nLjNodGA8NSa5uxgriVAd2vWDf1f02jdgOgAtc+MhDNXhMCWtY+5ng7ETDnCc72his
hXBrL9F5V1EMdKc6qU6FtB2ByYa/Mq+YaxXs4h92JDhvriv2VSS/+9nGGcnwjuOfqsh78jNOkvTs
89J/u1dHuFPQeIUqvQXa3Cy/xvFWV7CE0U5ogYnud2m+rXSfsaBmn0DJzyVFy7uB9iHM7ggeYtAS
BJiMQ9hKKvxMOSEqIjXXR/qsaDpWYFVSEKF6VEZw98D1SvZKqMzOk16KRQMu+gMXGdT3as7pSlTj
KjSeom5CpWYr0dYbpWaIGB4YpODYN7XVEYo8cxMjNrR8cZDHP8dgP9GapfIkoBY63/T1oabIvxfN
3K9rGC7hkOtS9AmSh8z5JhUDrU00CnauO3cv2h3ZZQ/9isZqJcVWW96wwo4PaORCXX5sxDO8XVv+
mHSXlPWIhGvzxnfxZoNu8rNMLz3V5a4fbluw/t63g7zolwfXTtjIMR4vxsKWxNQciKC0bEHPXAT6
JTRshn0rRVM/xF7D4PHSk0mV6/WQLUcot2G88jP8f/OzCnKGUiwqwR4vAKtlIGPgqsMK3pNo/y6r
6Zztv3cKtk0U4zL5/xGINvQU9GhC/n6oKi6U+slc0G3+o88uWHlryhGDxqV1HH1PiLU760tnk1rG
AFpEAvvaMpefPJugrPLTISb5l9PC7qafq6nKCk4d8PkO6ei1sGv+P/PEJsRD+9pKp5WaNCGinz2z
fu3Y1ASpeQbKuZ8/7qOo6YUcc6hEm18qzykb59lD2ECjoc1+R/6rMdmK6zBfZPdyLhHfxGdiu1Y+
r8XgHwV1fmRyfVn7MiGUVDtNvUP2lWVh5ZzumCqAaaih1L3wxIhdtE10BRittscTcPcYo8+iFdSA
YrwThLvJVxZvRzmlkp/iWR7+wVbi9LEk3HGk8xLNo+BQ0c+hcyw4BA0VgefBwWmGWKnxd86y1yAV
bT+yrjvdA9SnvxSF2VBDaJ9AF5KyozvLQGDyMHrnqq1+TAD6oBAO/+LvNxZ/VGp8xeSSNMl/QVWk
M2ZDhK3aABG0qSYnHz/ldS/PpyOuQs3bYlsIxOXcCI6k08ll/pdPtRcLcgUJFebWGw/QPZCym/bT
6ODObgOp9velkRgIpFKr+H/MjNdj1tgjRj5lE1NDyjCHTGtizG+V77K2bK6G6t865608qNwZTq3O
xQDkYZ4hTqNCHjbGRnvQHE6Rr540S/V5CB4HpyU5z7WqZ+wp84IicSEv6mEOrX+C/bhwBwGaHnsv
E+PAwVz8a/1M3gWReYmYTno6BHIGCxsBOS1fqRvLvTujc7BQ/i5snFG8GV9/wzFdDSNNSG6rl447
Wd9ZjphxUIxHZ7u0DXd4SHL9R5Rmefb40L3euxn4tj8uQ2HnWOG5iZ2FB2aiIuUv946EqvcXMZyW
C5KKlFGjfe1cnzjABFOpmcr4tEpI7fMq2Jp9VyuMWBxM1/RU5isP5bRuiIuwsS1MjJ601l1pe2QL
vbh+2IP83dV1kY+fKsHlUQxRnBNCZcrRol+hu5hrAS9cu+EeH4d3FJyfH7CxRjZXnaolcPOOJzqC
kVemGnU63a+JhXoVR9gw0yZA7aZHHR26oXZ4cYJ6BUpHAL4aTlaJD+05atbGElVOio4WLnYnP0AP
XY7rRvYRG4MdcfXSb+EuVywbKScFIzdbjW9y4W+pBawxAuZEZST2M2eKZWm8uLaOi743y7jLHpSd
Pp0Uh+fwvs8xW18Subsqszpf6JOTYrZ4/xClbTahvP4I+Kl/9qZtNfr2D8WtkxpykZaodK7q5Uy2
9kS+v6Uc1QmgWLTaWtD/z20NEw9PzH9sCnOuaLiuAmJG3fAMxVk45Ug1ANg4b8JXvGMylvV4giCG
79MT8k6zhMj0E57FBnb3N8hNS6HfmlhB3Rp6Qn5FIJc585JN3L2jauRM3qXiEKmrC6ySSNiePD29
kfWtNxPoPh3iZGy4fqnmLDIe9XREEdv2EU+aLXTuKErWWSbkJeufKTIrd2VPQSFva6mZG7THYkBa
TG34CnMluiqMMxa84TngHhDWlgZzdvYVdo/bDtn6ME+TkeaNZp+0QIePqfPl5e4k0q+jC8KyWG0i
ABzCFajqSCibNsgMUlYYJmpCeVwmtntGrNieecUdzJ+ckAUeYC5//g+agf2av+WQrt6XtLZVycrt
s7Rpi7lXxHVBoeqwhnJi+8vNecdD3NXuR1WgYolafU833VjkI5tkUyLrnFQKc0RGHPkTkYK3sPJP
sHkBG5kkv/1KExSZ1+vXiah0ZvIWx25s9v+wZO/l7pacY48YzfAnhgXWuxqua/L7BMXvnGJs2VCB
p68HiHeKjj2tusvbbURRE7dqP0NBxatc3mnXyuWxW4Bm7csi1lRWCtwcW0frjLgjOCkt2QXImQpe
1SXgxN+a79hdTjAGDh5aCCgQs9TrSzqH8mhwjHmsyYbfajfRKS9S25OhLHLMCPZ+/jgJPbD6BTKb
uumUEFkfQfLUS5RO2xK+SI5xAv5OqvNqkBrKasdrQhWBZbeOG/+kf07OwpGDrdbVNO8nAz7fqcgx
SO0mjH0pSI9YxXIlCZDTTAXDgNlWf1WqbF/U+jlySIAMYv6sC2/d2Ili8KMp9HqqRRy/IkVo3rEf
OEWD5RTJ6sxLi/lEWzukStI9wFE7WiLmMDUdAfT4qV0BPh2fMWbF/KWyjNrWVHSwMAiuHmOSXqQa
v2QwZ0nwEoaT3EaqeP5QlwAoGsEiT+dOqj7Id+aGtTny2siEWd5sd2cfxX74riRnzw3l3Yz2rvPu
1FRS5kweM8j3wVLHPt+OW23mzTfTJpziAcVgs7iYH4OVz2r5Iu0Y4oJZdklut5Qk3yPsLnWuZ8z4
SZqErDsY8ycUQlPL94fU4HWl0eY25MHSonGsRQovz9ExJ3LUynZskswsyfekckCqdmYHkh+coBMB
GZ+UE3OBchkImd8fVgPF1GOcC2X7abkufoGA0HW39MXkpeMXBtgUS964cgZ29FGHtodhw5LmDYNJ
yr0qSG5A3X9yID5LvnOuyAwSCo8dkX6K7BXaFaFrjVM0lAz+pBXZUQsVyd4x5ptXrmHOzgVjjMBD
qYPxkw/1NYFEr8P82r/cNtmx1zGkXC3Wrm94RX6reW3S4yvxUWh7Ro4SAwb0vj1ptmVrdEti0E9M
1ONpSjenWMoqEJL82A453oAo2BYfObALhiq9zzDgR7vRzFvRVfIkJhOUnD2FAkjdSjTGneuuN2+j
XOIbpCRK9pvgE2fh74Qdmj+DdlaAqYkKmUL33/1S4EmHvu1wUuFPdd2+n2xLzaGhMe/QXU+UN/Pw
M+FbIUpKyfdEeZ5GU2nM4Bn5wJHt4kHRsZrNvAqUM1ZU61wa8gJkhWsrP7gg8up8hxxDcq0JrZHr
0XH16CZ5IN36eQwaZoRNyTxUp4ea1Oxmiai0zFBnTF20FB1XrAyW//EfJ/t8JVqBjHwOS4mTn6w8
ydd16dAFqJmkhxaEw0g1tEroxaEtT+I7KUtYggrB6Bc+b4rgk0pRGvMiSDrPZ/2SHBJTGyLX9bxS
yH9hTLDFq6EEfJzYeE00MBN/C82OvXextMqYSCk0QR4s13Nc44+iJylPY9Iq2GLO8fFFalID6M6k
2FRhG6qYmVuFNP+1tc1FypK1T36TgkZynAS0TK6w4OHrrfFEQvNm4/LK0hubchZfWn8UwSou+Uf5
y1YgZ/1VRW6pF1GFF2k3CDPSOdQxBmGw3NeTQJOUxcdggaHWdzYj3gsQL4pp06oMjAyGMb4+NKTW
nQfaUcur++A1pubXcYUfWrlPI98q30Dgp4nUbvILH4emQtGtHZNlnzyo6uXNDr0uI1S/9DYF80Op
QMTMl+5h41umRdbHXRHBy/OKwNyvz9S6ZKdx5zHFyANU3HQOVMAd38jG9e8jKW1mcop+RiSlNrrE
v8OjmsqOeZD1EkrxRNI5TihGJcWB7p+bd+y7UcKEcEZd6SHxMJ98MabPM12KS1G4AsfJuQKlWRyh
YOEtkNgvPayhjtrtV6e+MfVmbnyGGodFPpKKN9Tdlk1Doq6n0QJ662NcvKebzOQWHF52Ww/VVz6M
fXJidptp0eFu62OEBpcaqcFU7iN64vDO2ZWdyaa5ZgH0UW88BbrczVefJusfaamOC9K6xsw0EJko
KHzVBO61H0uAyLt/lkTRljOtaO/BTsWESXXNQCa69dP1JgXgHSwaDwlBQMcfrifK4fHOAT8V+L+X
YPCH89bCV0CXLirrqq0uywql43JKvmBvWk1gitUDmqRdXORxTnLc6+xfq2KFSJrSjdKTljNilKQk
e1YQV+XAbY0AaCfS6FRE90CYXJtBiH2n82V7K4XnEYVrEsgbv+mKGnCNHQcmilrw/bUQgzCzOlE+
eApWqMSZaiiBezXHCqorwVfvpElhPsu/dMEi4QkPJVerZ7UrwBkSHR9RTm0xr4GqgqgRva1rFQqx
tK3/efDXkMR0JnuD4ZYVTLqYn3jW7OtSacBo9GPycuXLREDGyq2aD+dDAn0RFeydTFvPGEfC0gcu
Wzx0pKinra47F1AUXclrGcBS1IIv9PrTfneXXhqM738iaRHCqvjIsufbA7aS5uWDaa/U9pU4pX8Y
5VE8qwwKgRH43nBIlYQlbjkTdFOCym/8c4xMJZ9vJ3D405+DfclundIF67vPXV+1NrsKAI3gTyfV
u2LirkJDi/cn5cgvUdp6MtWOdY1C5pAGMX807+kvEhXwuomqGXz+lf2AwVCCUNVFe3IHsi+aIyW3
iLMpenvi7BN5Pm+zDzK8F/aR+vd/b0WpUpmPX9beQORVbx2MG9GUBm2r9r3fvg1eDcEPpROSUnpX
NNUowGO2CKyjdi3Fr9TgD3WxKI6ViQWWm8RO3/ca+BOcFHFyjK1wEZmW3N4TvSI7Os/42m1oMJNg
PIIgSo8VYTVu5TL3bh1SK5OdElUIt8SFS5pTuoSSa1OYgH932E0+Pr4epo/pKgQxfMhm0SEyeEQV
h11zJLTlpfxdTB564tq1SV8svu61anyDIs6/XcDoNeDNUNqQgq2JBPyEcwMgoBFDrvwWniUGf6xW
/a6VIuRjtbQIT4WEUgMAvv2LNZJwP4p/1yq+k4KEnBvpqyjVv5pXbGn1/5DoIWnn+KEXau5JODdi
mQsCEPLtIeVl+JM/b4WMiLh0QVy8fmgnpGMoSHo+t7bGco6QBqWHSySY7s0LwtmuYnwxLXK1o7aN
GUExcpV1kv3L1Y6YbwNetwCkBWWsWgY8DMK4mWokkDv6iVQztuvMvNUEO/79wbrz0xm6kIPC7Ib3
UVfrIpdKNU26rHVINhD/Jc/sNjLeEGuneXIfqGpHo0d9627a7LpG4FKDPG1ZzI+HGB+RBwCvMoGy
XSKhQmdc84snflgHYCOZZGGhWJSo2LUyc1EVKq202glRqfFy4hhtw+YJ8352L1T3ieh4HvnhrXYB
W2VBf6nLkfHWbb37dIq7eTkaQ3Y5kR8HLRrpInAobNek7AX7tdVrbXv9Fpvu/8BmxUzyD+lST0Df
KppzFBr2J1A1h4QAtUorNBqB4k+c+E+ATG9aPXoxq8Cbfp24drCLQ7xqddftvLb3XjGbebHVXpSr
GzZ5Eb570T4mhljQAKhMQY0k/poYwr6ZLeohhS98MdiBxV9Zfjgf5f0LEU/D4UzBQDGOxiuLUXTg
XQwupP8sWjqYv1Mpetl6UB9zvZilMjs18uHEFi2deVl21QJZOh7G+GbcGZO4dSwwAYQQ4O1d8fLo
UWjh8OLrTHVWxmHKL8yc3kc4ympeFE3A1bw3sH08UJCECiCa9w5STi7W30a7sZA1m8ZP3x+1m74/
Pco5x03V1zAW+qWhMPcq/hM10Ir6Sm8nHrVLYwOSW4JONwhoLRn+LyhUgWVXqMAWzDmi0XKWpocr
vpT2t8COK6oFO8zrCy/GPrfyHO/qHZ2s2mLj6ZeKdwlteLJ/FzT2yQKaSienpjtpsbfzUq75SRJe
vsOq3IESwH4e5j/oXwJRKcOaVjHTwd/DM5DbWkyzzrUSZy56JN9AB1sCwY8Np5zfeK1KwEN7QZpz
xYxHYhrAvRJtXqPISEHSovyNNAoIgK1QN0WOeI4AQyppf8cdpQoKGNenhYIuo45f1LBUYsOckNT2
Zl6zHZePoQ6HdFxquzQs5Qo78Dj2cTw9C2I+jdLpNaICRLzdxYccsHD2utSRmD81G7ptIb5jVpqV
/FVderNlukc8Jy4yMSM37VKdQqfwbaLFTRFz14LeKhT34BpfbNXt1vJ4pCV3GQIeudkaZ4zpiREx
cgfbVSBk8wRhEyeIpxydbWkB9x9bKbm7qYVDOeh1gbuI5iXm8qXxED4hjTCEmDSbWc1Emc+zgaxk
PgXP+WV/lC3eNS4Tl5s2ZgP/lQVn5eG1tITErJreP0Ck2jTlhRijRmGN79h2buBQX1VFpXNg208N
KztvqjEup2V/4CzPc0qTqgAzcqLhGUlU1rN92GPn7thOgPAV8iK1Px5hdiSxhF5npwmhAQZkfAq1
qgyFUoETYar96BnT68Eq6L4q6/V7kAlQptZHjUBEeDLxBaA3euXq9o3X88cABMZmdaoPEqgrqJ5B
kfpJ/PRDlcgX4UzuSHsfTG6I5Fi7W0YyP179kROsO3xW7MzskSQSwjx1DxHFBDq+azQTda7Q+H6+
lJz3dau/XOAYptQWgGJ6WrbzN8I5fldNGi7HxCByknLUGt084Gs4+jHR0R+adghn0HPv7tIYfvTe
FwAg/H/suL+zKW0MkqN2M1aDf8g3pQhMIbFg/W012WO+my3L+s2gAcU5DxJU8ltxT0vgmOqnDpn6
M/PhTpLE8RNGCC6K1f2uME4CNmYT7WOJvh+dynu1V0PtYQsO5UWXaJs5VJTU9dE1lou6RHGOthAs
jqpjzOs1ZmO0OW1d8D8GKmfEZts5xt9dETh8PHnTpWAP2p1AoSq6JFuEeyFVAGr540jQ53lepfAs
HXNTCcBTfyRs8rk1sGbjLJwLn5RQXSzaYZ7LNq3X+E0gsaDIdNSV3jfx1ItWlG9AUUPUsdMft0B6
noyq87O3fB9e9SvZg325NZLreur1nfN9OxPqCHNQF66YaOmgRp95rxsUEnuCNx38+wlojfLezFIR
wqCZPFQn+VG2WC4VQpV3qo+oUfLKmdfdV9W96s2D9ZDCo6FdsUJkxxtswf3er0rVwn9UtrUrXy2N
IOSaWHb/GhwH9zkiN57Xqw3EOc2Bi1PstgBWc2RnnCizc0hJmEByEUj4WQPUS1I8xWC723ilVWiw
UFaEchkuCG2j1uqGGCVvgZwYSR22tiokC3gmjPb4HccX23ppaFAt1sc1Sprl/zCvxhUBEQdijSw9
PNOSwHYtEoUTd8gCyZ+KlHa+2HfCyC/1seuSnHb2TW25NiEOh2492yF1xKzlXCV5QrxOtQ6aZz1n
yNvA/vLdHwYVNvOH0pMVStd30HKCw4KAeXwguzUXBnTkS6mdpZBuCCqZ/S7B8SZcu/LAFvEqS6+g
PsmvpS7Imap7MKf+mn26NqSBwo1OHG5H1jVmA4dZtCgky+oDDesTSE4N914Q+92ZCUy/dQNxvwaZ
Jcs5XyvHGCfXbHPhBrkxJdxDLgUJQ8dMI85y92wbWBUPmmSJgC81a+L5BulsPtJZFRMxXbLVfdSS
pNjA5KD5tIaTR8hFpEHcTfH4yEJxL1ZuejpTgDkpGukwXiSCMDvnIDWdUORoniCh2ses6NgXVPYi
GejkzZ+YqBEvO3lHWi8hftsY5Zs+JcMhiUMUFRbodsg6KTfSSQY8J5z34OEv+Gz3ko49grnpzn96
3Usfec1Haf2kKoFfRvQIppsk86f6npMsmM1JK8uy/2aExVYgvtmjKUoLmO0prO5II/hN1K/nYJie
ZTYmgwLLwrFmE/hjeFhiYtQ6ksslZYZM358OTdgom1YPl0o6UsaIUuio63MoQek1fapzFM1p1+j5
rD0JkT0K8e0fLBWWRz4SLLsb3/3plJUX3bnXlEEYggsgy+1bmAGM1l+vsTdGLxowdzQbnv68Req4
Uen17J6wmBVopze3aLzswyecvO2A2ZESOW0Gg5ktcBUa5g+LWYFR4WqKJxhSYNWWqwQsl2AHa9oc
o2y9VU3W3W0tEsp5UC29587SCrAsCRkPSKrX9s+vHm4Y3YRYFKVvWlgAjHlsM1hN8z8UKMxcH1Cr
PHjdP1ZTvtboBS4O/baN+rYaYOO9koqO+Ml4q3BfRqMdZgnH1sTrlqTZl2dyjCmSy/2aWk11cdoM
lxcq+bxEwpZLGwt1vGJ/qPRVkXaIeC9xJGuarJdUopp8XG/dGM5925qA032TKCcdCgOjdnfmBIGI
MfavT+chu25j5xDaBuiSedx3wkgkYkv8tTv7MmiKkVIoO/PW3WKyW3tLempDivL5EoItJ3XwVPdR
v8b6REeqAlc0Ej+oNXHB1C+FW2SGayyiszuuL7eSW5cU+HCEXulMCwhgCRjWcSusPjLJCytp3Yxz
FHbK3M4L9R2rycEV5n+tfs7n+vpD3qE7TRwGAeGU5jV//VRfJTwjHorVzn1+41UFUVnepjjc+R4m
HvAotmcafRczgptKSRbBdfoomWKBgYqLdiVpJADOOsJvOC5zvm95N/kLSpA0mk16yqu0KcDK39Xl
f84Dkk0EiuM7X1Qhn6CORFA/uxBRfXSNKb/NdONKwPVOy7EoFkDi85qRZdAkp7muJdWoe4qlfSKV
YI6vP0Y4knMRD+73/Hg0JIZONlL/rtt9u40kOq4BSSn+1taCcjpAxAT5oiQr9MVwgeAf6o5qdP1/
EbbbVqANVMJoSEbrar88o5AsKidf/29SsEN7LLPcDOs6iTF5mCgzFzcr0xrEkhntJV0thjVGc5uW
4HNkQ2103RYO7NfE2r3t52c+9icEcHbVdb8833PYjuAI5L5FNgIVaM11URR9IL5RkfY1gQSo/1r5
2UfAx4lrUIVHPY6pS2A0E3OisO36qA6WphqiQAAjYaLfkgO3vudyL/vcG/uss4veXC4CKnKBo9nY
vyy7+/P2UBV23ss5RKFjX6COADHkItOz9GM0dH61/9ad2O+EXdx3pxtGgHqyLy4FARlzvmeH/p07
YnC0uR9cqIcMKSR3J/4EzGPc0wXnP++7OJ6BZopje5XvkfMMuYWrn8UbI7TokSHGxW9+iQaJsUIe
u3ddQyWSmtsBUSYcSx5BvCqowKdwa1HR56GYD2f8Hhj25SebVOchwbrQspsyGPYNrOhXAgG+Ehwy
iiPKYFCUdEXgaue1FqPUIEN5jPDeZorfvHY77gU7tTSN7p3IrIcw/zOBZgHuHQLQsne8Q6ymiTAF
0TN3MPE9UYTbPCEGkhOE44mSlrsPX0Obdh0bV9Tu9fLZMu9WrPzrxmGqfiLRx322I+dm5FNdbF4u
pHuoiHa2i90usNbNqyz/vSh3sykKfh7Sf7ANqfvJYZsI6SE8w4/NJ9aUsdrVVrBlM5WC38H6L0Ty
ywFZgGxmhX7keknCLri7Lf+POitslOelteZ3Gdzj6syCszV9tuBRPRsQ/MamqV+BlL3iaPtJK0/+
y4enSalKG06yoRoZ3s9HNmeciM4B/E5XUiDaEuNb4W8ZVRrKRv5i6vCc/sGdwP5xTYpx2KwZ1wxg
Khxrnd4o0AHiIXd7cvuJslaalQq0mP4rRc+6cv+zK45e9b8h8bKxWXaNOBM4z0fqJcWEw8au1QiQ
WyHeouaM6VOP8ZKx9sjtAiJrA+FptvdXrUiwLY0scChy5T0rQvTJQHS5Cn/KrUnY+J7CX0VKemaQ
sPrFFdwolTsE055E+m1zrtEu8QIzwWNU4dYHQ/rZFmJvxTAcEqliwgR8JdpUxeFodZzgqDsc8Fmb
Dy/x7l90gC2EuLZiLl4f1Y7fTpFQlSlo+s70KqyaZCD9Zwr4W10V70C8hhpWWNin5llrvJcPojE/
r536oru986ICTlwDV2VF+WJTzrvUfjYs6BmVetv1HHFi6bH5XOMkrvgBy3PuyRgsp6TTtF7LiAaH
ES71AswM9wbsV8a8IFbyRIJ8aAVsRcDVT68v+PVhNWUDlxyjLhPO8SQRuQ5Xqle/Vv+nuleG2ZHU
zjWOzo1zo69xXv8e6jPf5zDRAtklsCMCwgTBAN6F5vvrthfQaldlLtiBr/15Dnr+HCP3p+SgBW+B
T864tqRD403QY9oc9XoveVba5tBw7pUnMgo1TKaq6anfqeDoc+AcpnGVf/76eUytI+jJPsmNdiha
kAgsUWX5g51FafO+5mlYsDuEIP3q3SsIrbe+dfKab+keW8PrDXiu9EBgRROBXcAO+lCkEMTOATgZ
d895LCgHp3ZcRUjWuOmFqc4nrgZOwADwB3/ix1wXzLXV4p5Z1VYrtVgsVKAbcj+Bag9Hyy4QTtIj
iljh11bxZhs0sQJqnp/VZXABArDMy5mdDteUQcbU1BINVQUgd4GyRB17qxXFpPmuXnXtZuS28/Qz
yUZXZLkTsxBWW6uqla8yrMiQnK0uAJUMOiZ4TEMpIVrpg+JHwq1grdJirHRuxfZf6685pN9zlP+v
xrAHfTKEdA8JX/J65GcH4xfLMoMUhIQjPPrPMwE9KnvSRGlup4nk2CGpPcfMuZrJFi/eCKHPBPJ8
CTtnMGaJvKivVB8I5ESpCd5c2Su8h306pxonVWR/435S8PTHZKSDmYqxMJrctJVzaW/sdv48mj8u
Huoh3LPJlCTaaylvakdexQrWU48SZPCa77uWaaQvqzXAjfjHOkAUEXstCwjIZBYcL+8etbTDObyf
UCS05QA5PHJWX/8JwHTwUmx4AB1zO3ypp9ynFXH741Su63KayyTZd8mC0ALAqX6koBvhpfEgBHDJ
R7MWNXvK64a4JL7/gHZ+xaHpNOgvgS3niLuc6GDrNIsjTOYFvDt7VjFkZ9hEVzUKDwFiYA+B0KRL
hZamTCP88gNFwofWXMNCkYSGNSSLtWyQjud9MkPm3Ei3DwOcdiX8/WWqbVn98MZsXr1BqCUIF4mB
bOtTXqEAR7YmVP7VNHf/kYsx2907i41I79jwSYiCRNbhDWUuTH2qButyzfomecaNlUelphNzIDXW
QpvYntbElv54nAZQqz809HDtRtvnBGhaynjo+b/HC44In+z0LpQQEN6Mx4chISy9LBeqD5G1EjcX
ucnAcoNWG+1RbhiNkkhQCpaySQghHPwD0O5eyN/VS9hLsdIxfif/F9FFyUwdx1pDiro6yAsCq0Ij
PK3XY+jQYi4DtKP9ycqXwDK1YYGTB2dYxJBjgZIX6ZQJG8XcI3DWv04Cpn2aYpq4VwNR00urhaVL
0ubQLKxdxWMRmPvzGpkeS8o5A+BeFtxmHKr/7PbFseDijkRNPtfJTj+FqhebIxIwODm7gGTicNGs
aqw4io+1a7bJyP9+qGnz6C86KwWKvZRITuDKNPayT6/8TUAWMVf12GbIdGVn2lQDFjotUQR5mevi
drLLDIeAlZp1l9PPf+L13We/hUX1icHtXUudMVP4bwoEFHSutJpf7UJQrad0Os8xCEEUZuYrhCzZ
v5ARGs+Xk0zjDXeUhY6MGbMQRYWJy7BJQ95M9Rcs/z+CaiQCV/dEdtOvxb3W0WGbxkUDaiMz8Fbi
uoaVvAcaCz9ejHeelMCsKdtow9xhUi6/ZoWdgbsPkjlJKfesJnxcQTmxiEoEOS1xgGWLXrQ1XlWS
9BwgNDisGMyA8YOZhBunpjH/YJbvScFIthNwJM2g8Rsm1fanHE2AQzEtR2eCRCkV9izoQied7gsi
XcX6cyid6Rkwk39DAptSvWEWdp2ULtnABOOhL1EaXzxCAovt7vSFqqWCiWQBdg7R1EoNY4S6bcyk
/W5m6OLth4jniDkl2nwPPIbxiJN7SfgyjYIl05eeMZLMXDOy/rjmKc7EmaAK5tBAVBGVBp5mvq6B
wH5kHyQUpw4wwecJl5klOE4BlNaLJpKIQ0boVukHligUV0kh5eaufIXkDUNe59GHBBC7xZaVtOEZ
D2ig0/tH9BNKiLh+8BSjjGVywEnWfvcKnplDvBZg9W9ObcGYFbgUOk93asyij9h+i3fDYWUPOJx6
MzmAKSdSXoBA3aiCEgiGf03mwdkP5LJN+oGLPpFjgMI/HjCJPMI3zQyX+arVHveu+7leegD03tKx
qQnKTIjrvhguKMkwxg11gAKn7uXX8A58ZyePzFVHoWbZ9KqP6bgne2+U+Kkt1Ph0gitxLkkvQks4
NSYxmzktoIBs+j2emzpS/O64Pn2EEcNHTXtSf2spJqo2gTLN/3EyX25oxcQEYs678y9amjGqApFH
hmP9W75CgOMMp1k8EEoEOa0CP/HWxJyxIyXllPpsad1dNLcWLr8qqi+Hb18Mc/VhW61mqbiU1X2+
46Xn+lYXujrG6Bdfp9qVlbqznLc10hw+0+yBxXYb37B+fswVbgtQVjVjOsKT51ETw6TSz8YgwM4Q
wpgF2mD1Q1OLj6JK+NewOD1cfkZWG5Jt7QMpO0yuaZQQVtEyk2oSHTtte3r3bgy6G9PqBgN0jZ7E
BGylBKTWjTFOBR34i6gQCc39k43UlCo3XPrabD/8wXO8wMdn2xtMyWYT63SG5UFAHAn77bq0xJWD
iLvhHQH2s1YyxmkoPp2RKzl0YVptUuVy4kDmu87+6Ujy66K2hHOGdjM54qgP/ejL47nHhn2CWQbc
SLfnT7e/u4cbOMbZ5JxKI+0c/os5++/SFBGia4j4BFaumrdPATw0HIFLnoqS0oifVoujhVUB6myS
YemCHUIQgofmkrqLNPhPRFdD0SUv+2AMirB71X+IzPmypGudlaJpsELLY6VtUrqFcVYwP/Y/NJ5d
OsaMI2lv24xUpC9aCBLw51g4RubaaSfVZaYa9wodDjEMxxwKokicC3TpXoEIhf6AdcUiJvUhlQqm
P0gT5SLtnBDCAPl38iL2Ch4X9U4RlyNlNOPFIpuwmef9FI+92k5hZ/Ib8TP5RoVI9aEp7JhBucSW
GR7uvwhsVz7qpOWEsf/7sasvQUvep/bOpv+4aOBGXFg6fbBt97cm9mL6J8qtLMnrExA56iF/tPWX
OcoC/P85IntVhCt7sinwZPaS4gTpeQUR2mBzKOiMtqHSKJZrBYXn7WrjSFtPtj8Kzprck/Uly1XQ
UbtNkWjizSmWqZk45yr2tHXwlNIPckMIQznZziOxt2q+U2CjX3oyY3lM+90p9f51HDjf45oaW9n4
jzHAt1LAPT7lbx92bfyKizl4dOQs/Qqm8K94bRXoL04poNgT2qg4Ap4cxbjCENYUaONaTd7Bwqu4
WMIP5Jbhw14xznCHmUES1kBtmkE8QXSX9o83FX0ZKIp/T4H0p5+p5wDYhTINASRjbeRzxg8TODYX
elGzOf3/qaXpM74XAsiCOlpy4P8SAQ0viJ5PKZBYZm7VMpdvEUE91Sy82oSkNgx4Dq+dOWiwlsoQ
VhlfuIE+zYnyUlfGVnwe7Y/FB6H8CeqBrD7Gtii4hiPTUtsL2prx+5LXjwVE/cWxo2v9BPqWqxBC
+O3sUsXzrz8ryjEGhu0KAgcyktmFe/LnViOvPNhFmSDfrNDPLqVf4jhDE8qu94kZqWRpF7r4dUpt
wWCQq/lMsfm7mmj8+/J+bQBDLohNJN8pN/0bwCtd8HXnaNP5cSTyrQeOh1DGVdy8TF98PQxHPPso
b+f1EVy9MqA5uAQg511EMPFVVvb3Xic+mR2yfpst//082ZC/Y2AaDIdEJ6r3pxVvzkyLrRV+lmLT
OPB8tyl7SCjoy+6QbT6q3wjLDGoHxGmQUZWUUArFp447oudnZIy9tsQQ3g6GA0dOx21dK8RaDfRq
X23AgOcSq7prCBdgggvKRm0n5WFi979/MSYrj3RRpUVP8vxkaIo8giSrO0PoA5ihvb0GNK6/sz/k
AtpWyIW7F3NL9zA/bEU0xezwQWNEkGgseX3VBTjS/Q9AvgeC3gCGudhAue2dEOes3orQy9Plc5MM
Ep78uaW/rZX17uAiIvbmHkYogg+3aXIKaZvFol1q93EH4Vh1fMD41AN0YTv+RIl4SA/d6o6vLoRz
31m6akz95tOiBRo9JzX8YtothvzaiH/EMMB5Pum/q6zM7Ilw2znsDoGwWlC7txG9JunDqiNAipuw
0szs1rIfoalSN0FhuYlrZiT/6a86uiknaPnqtX0rm/Rqx25D0Uxpmy4BAutt+Uuc0916GEAsNTMn
aSB18jq8r8wZNXb/rnYgCUpfq4+v8vKTdfmzuLRNQ7+uoR3Ctczv1GvwQaO4dTIMVKDy8L+V54NA
s7XoezhwxlUyjezUlqOmYWLT6apAK+210ZxHx4g0w0JAjTYlx/6o1hgLyUXO4kD2QIYLmnY7m5N5
1NWiEpQ54eF+6QucChfpZLGDjJCJ3EqBxtxuF1Wb2kvC54tyHLaKLHX0C2Cq9Wjs9tL5V+frQKPl
UFJi1G4mLix0WOKwebWlOnngec3/iFwdlluFSj3f8A1ichN3Q4dP0iCAolYv9pTjVz9EZPxgWTUf
iFGwkBMoF8DCUBWaOY3acPYCFlc8nVr3pkWMovEdbPFZXEYXuK+qvbCgMfbqUIxN3mHT7VGyeOtA
j6bScUfuGObGPpdZGjAyr1T+jP9JT9eR5LcFaz1erBflVOQ7Xm16lQD/LLvlNuSBSrdIj+mE5743
wnE/m84QuGTHP3SYkvYbODdAtAuatF2XZDBpdpQRFvQ2hs/oAwwPn3CcoQ5fjU4mQteaZ5lmId+R
+CwVyPMG1vaBp27L53QWEjnTHTohTUZZUMR9S0qGT0uOo7M1BUQolL+bnK+oYIW7PzaNLfWFr1ZA
71DZSbap2RA1OiQSPJIfqKb5sJqeegAEiYI4acr6yC0w+QmkiuQOMoCq7OtsvoWrd02J7nB+mWSV
qoNZjJgbZ3zjZItsj9g3FhOCuqPZ1S2gKQF5dIvZ7fM+9XaYsQ8Z7iiufaDN5QIrmLPY8moR6+CJ
aqUdcxkxUlZ5F+Efr0U4AwxzY2RLh/y4V6QNTvgbG7vEFoVAKS4ctfqgeOCqUEKD2a69ABirJhyd
642Lzdf4tpWZdpc3E10lry/K57oBipQb8y3m7cMwg4qqoROzxNBdZIwE63JaJNLzKyg4X+PTBVV5
wk9fgmZ2yD1k4HD5DbRmqCLyHELS1PzF11Vddtm74o00E+Abb9uSyycH5UwtWyuWBiLLIPMhGKJV
httOMvaYoip787ATlr2PuC5MtKr+nBoZ5ZK7/TWTJHalbRvASr83Gqq+jwr4spDBDPzvk+InvYDn
BgVRyEtUMvGpN4Ptb1E4bdC91bMhsnPLE1VLc4xlg6cb+Sqom5B2BZX8wdjZqVy6+J+7JsvcLTjL
9/Zdi/mrYI0ykd+gsEruRPMSUjqrJa2ZkxQx5yN8QdL3PLC7NxA2ZEby+W2mPnfahI3Q11p1VEc9
DoS+RWvKScYLkQ2C8B/L4pJoEEU5oJGivOzthc4LBzP3lvx5cKPhWCjh4FVuwweZ2wvdyCSOycQO
zuBz95prIy761veIgOFuHpDuIB/zmpXB5uxh3XFtlVtiiWcVEbIhaIGplkpIUEvJ/hnkduzlQGC2
porHnX8MxVwpuJWq9xufE/ubPbjksRswoUmDtLoptcb6kq3fSeUFOyGtjePT9e6kG9LRhcD02g6h
ARAPeYv17q4UglOaBK8K5Lu86roj8TptCVrAptMqaIh4q29xYkNmipqo03QOkO5UH9ypSXNxpLsv
nkxzP+8O2VAlPMamONDNjNBiBqTA98Qd3bXl3hsDwtVM72D5f8tvWoRS/w8LGDttnO5GSPUJx+Dz
4k65ATu8pK74nQ6uDTqQ/NnmfuFj/wV4yWzDGkMxMe7FN+CT+fc03j+S8r0n9utJRaTtV59H10ij
Iye2RPpt9riTjCpKlUVFM3iI99ABekofIB/NFX3HsD1+4nL5xzS0Taxi10ucXbEg9KwWHhDEr3qr
mjMkSAG0ESivNPU4+B4hU2XvDWNxKlIGhMLIQnUCc3vhIhc2VokMiLD1stN8IxYb/kK2G9LaggZS
t2VidknsAE+PmYZ5/1udPISNC3gmj2Ke1veyvt1j1FXAFBPGCcL8KgfBZjhoKweMj6gh5CnAWDak
9l62AWNPKYzhc9hfiV10zGzj89BMbkvAY0uTXu/XVpGGuz7VO7fuesKIXxD3WWcQhZ+xLU/LbKJN
9r+0CHTVvDSJRXhZ3nIImFxm0CxazFo4mAqD4sTbos1Sg/to5keiS8qIYlQQD/S3v8biWzXHzXEn
OkyfIxGW/bnxSakvah9ENFpyGs+IQVf7GlqY7gjU+4HlejBs+QFJ6SiHlDCaPPcxYb3Cnb0yQ+j8
xmeDoo52z0qY5cfMcTwGajluywqB3cNx+N4T7P0uf9Q9dGUec3+2vI2LGk8V0mMQW51Zsfu6xX9S
OyxbnMeIDwncG5gQ6mPUCMUCrTXupc/7WWsT9qDMV5adimUZfiGmX9s2+2sve2W9QRpZe3GSHAeZ
5JTgS99bLx2SFh135DwfBI1xyB97Q45n4hDrLTvzI7XYrGWO04b+zx/gMqu5PFYTvF7MPbqBPd/u
v9qsPqKWS8WTGkKJ43PVnO/pxzuskGC6zV416TF/jVEiWMmZ4oxjCQXPp6Pm4c4HAaSY6ERuzEQW
cgDMGqeh68laHD4s0wLgU1AkPIWEkIJOoe3qNvlkuA53dQDXsaoe1WgpmUj+mZiJwQ62NvIEqH65
Ms+bBpY36dCTiiRKHyh8l2BwEpo0LKI31C3C15I1ZVOBhAcf3KFPm+YQhThbG+V27xuYSOrubfBo
Ral9mU4Q6alx4MgjAH4nNHmervtj3pLVklSh/PVteypZIiQG3WBYvm/Kth2lMuak5i8zSaOqDXIo
EzlYG4ThOnUNWOddiJvjK7NHxiU5hz98MQrfTG/zpeFltm8ooOr1olXyyqDmNorAaVRmjLzd5mHN
v716OrDfLAAMyvZ52Bg2hlbLfbmxWs/3jV/jAFENQ/4KmKccwSVOHQe0Fqwy3KNIlKLcQlU44MO0
6RgKpw9pAeWdKIXcz0jaVdbU9RXDOm+Q6L81w3Ji5INpqdUX4XICkumOBcxbOI67nFwAEqewzrw3
igrkBb65IyRMIzIT/uWzghLAUptmkUkzPBsQ/Y798CtuaZ06oMrOBHSiPswSFp72p0GUGPVDGowo
ILvDKN2ksFitHrwqhrfIy3ujrnjAWSt25kCMo8pNNyRHSUIqARYIDhs3sEgsXV+KPA/Gau9Ux2D0
PZ4Ga6VusiQPPmeueYXop35o4QdBB6YG2zbjjw6mldHEYJcD9gYWxapKFOCluiRd8SsKJqKcAnhG
T9F/03ci326fg6dWHhilHBVUACyWo7xXhRoShE2oZfW90w8g4paxtq2r8SrAji+pjBw1MZQVZA0v
nZrhZ21MMFgTrBi0TyiuUzWHbQhhMYqKud5WVtXES++R9mOMtghxCy3swbXSu9v0ZboiUJFlZxyF
sDCNJTedXZbVJgeDGhpG7o4eFXHuyJ0aZxCPAfYGDsI27IV5AMMW/sJwUnPBwxdYydV8UqNrgj2+
m/Wigtx3XVbbl1dacIBqJ3ryDx1DJ1norN9qHsaczO31kg1D98eRjUgOos1tLX783FXKgfHryq84
HltJFBorzpYCsQj8z+X0pz+rgCc47+LCadHfUZ/1w3K2IQHgF5eSeuUs3aea8Qigb9q05bZAbm3i
3+xl+CuZoN/xG0XAkSjxlO6rlPK8IlBeaUsTcObwmqcO06B4oPNFZVglce8W2nC3GkufYVbrOuRM
Tpz7JyxeqbG3wapJ9XXoV76a8sTRB/c25C9+vrTGP5Zw/QxAcsjc2rDUf8BrdkNUT50qFrqsNi15
Zdv7fND+DwlZHPWP7LRQ8A4xp4UKs2pocdEwQ56jG1n7+LvNHuOQYIY67xtATg3fsA5MHXl86ROZ
HWxLoYJuCzyMUZLebVhQjD7HtcBYmC1oSupZmSmPaE+o7JrwJCL875ygS7LaYEhz/XwiiEj2zHQN
Kldy6vWQEwwu3CQM1xzvEjynvFyF99hd5W8d2S7YQj32Xif7AKPFMIBE/6cbr52+kHHhoGuS6Jn+
L/R5b0Z9JNK0cvFc8Fd2Ljevy2LrP7hBDhmHnvAcB6nTRLYLTpku7DGnPHSYCkPRLwH3YNwrNxZc
NASvVmb5stVbFz7r/I8aRMJVt3Sbxx02MVz1ynPW4701ypZqopAIlV/jxvwUR3maFTOwouPmMDLH
C2OWyvkUyzCXKYsed6/mdO0shQwTt3bOCloHYMeiuOd7hRF2soHOzWF+j387/Ds80sjfOfHUabkQ
tAMN2EXs5skpBr8Wuc6wBSc1azI9706LCF6KE+N7NumBYmmSVPcbkxhu5T6vIKmAQM7SkiLvY4aV
Iufn7pyHl9k10b5b2vXUix8YeJifIIskqhwUdRq8B+KRJKfQxDkdBEusFdrJ0y+Vau9h4mwjuPjG
Zvdp+VHn9wg66U47jKglxqe3XwP7tgxRmbb9alSOPGkD9LTXpUmc5OkPdyAhtSZIk817ZtZxLJGc
9KDzIKW3MztZ4ZP2q7U8p237fxkRqVYclqu30RRItQdSlCmKQpXiFc60ROIm5LIJDcAwu86Ltq55
2hzaJujrgh7tWp25gptbHmBNvKKFD/oOdclcDwE46grzgNVCQUETDW0JtGzJBTF1uiJPLRIA55IR
cHL4JxXEdMH9BAugVNmzJ1EdE4nuIgX89crh3z/9H8oQIUYvS1fkzxbj7MI0sE0M/ar/johErIl0
npCJmH7CH8qCtGJ1l+nY/JJaAgxMGsybU9GsXn3nnoxk6yfoTcyLKzBBRWJa4s8Oet83I1f5cKpa
wjq37mbGAeslk6ZvCUo9lcyHPiVSq12i0/xG6L1AzJLYynJ5uMNh1swt5hLinROs81t04vBJUjXa
EKr4kh5ke+MYQbbsQilzCTHC33iB+ehLKlGeU4PxaUSOmQ0DBCLh4uDLlsZb3kPNDfe8wNiONSMC
W7uRTRs0nc1ePE6iIN2Qrv+bqpCh1fLkfuiXR99fTmPm4rPzLqVdMPUhqS4oj6cXw7v43qtzKKKU
WrPMDTpu9RDCWA2wpisEQM+FqwdTliUphkO6PwxI5xj1Ub6kepGDLSBk7OZRyrTfPNwSx4Ry+1CT
c8XNIwXjxPk54wp2XSwbc4v7WQL6cQVod1OM5fh6SYaS9x+0mFfKyf2XIhTG6LlCid0CwMOZdbjZ
r6LvBkeevoeLrxwpaiwSAN/iqap+NAG+Y3fD9y0jI0G6Zsz/9F7htqTZkSLt01rKRCz/d9svDzmK
3vSZZIDcl98d6yMwRH1Cxbeec6ba5UV9aHj2uSJGMI+hi6bw3mvJWHaacJuJR+IKX3AF+dpuyQ4D
5dgO8Y3QGzXyTulA+vVFoSZXE5O3C86LlAhEQQZey3CIumubi0xphNIqg6n1E/LdUqY6Sn0rl+Bd
zGnn/uGNJDF/ghiuycLyBUlwPNzur+qysY864ql8Nr2BRxnSL4bjfVoy6RyMsFVIZWCZtoqOYtiM
8xIVMpdJt/jLismSaJDJv/GWs/NUMfwB+GHveeTRhM0TQZQSV+WoqoUmm3SSZ6zu8R2q0Kv6JCZu
4sTYmTV69Qyf9VjoTO63H3zSwT7Y1Ha3WALg1CiTSY+kZF2wiMn/ZzZD2fLYGkLvx1FOBV7N50Lx
TDxUAyXFVZbp+qgPbflgIBFKglE/ZyYCLLxjg9e7CBjwx1Ji9vb1OqceyRTqNRWu4k0MOJzcwgSf
maehg2m1UGhb4tGaH4EsoaDDJfjXUcSlmLh2OzeCCKRSa1zXtTsPAeT0zpouxnO+CuWCzjGg1Oje
XxXJQ1ESkAQuGvwjx51YvGbnk8RnXdkSzpM6PY3lORXq/4FlyymXe8QdgQPDMGr0oM+mXXsN1qVk
i8Xj/VD8QviIkpTiDANlnFn+bQMRF4+eF67RvhH/PVbilQFqTawb7Xqxc60PC5x+mMzxaKtH97An
st+WDyu5Wy6LM5AEUD12krj75mhYMSovZuzDgio1X5o7hK31dAmHclfURidUIXzPjr8uzFmRWV44
fFDJncUZ22D4KpXfDSqFgQ4fCNEEn1L+fMLXzztIbOwmyZ7VilDQJIfOB1JJZuje39Tv/kzU5GGU
JoZ8N1LTg577eM15A5NfR+A5igRAklVIVfym+YTOvlG1a0/FBuiuI9tnM/T3mUbeKzpOdSn6RNlJ
PNfDt7VJ7fssnKF+RyuCciG7XWK2iObSQR/6nzcSg/tgcD4jEUVfXTZ/mOGZVbBXahfRGTitCDFl
v/zSKkQAq7tmYVxu2Tmd9vPB0eWhn3U20IBK91N1ywPeZcY3Rv/4MReYtpBA8Vk8oBfLmPVMSkZ4
7nFKzsIlsxnd/p5hC3w8FQRJRrjCoI/UcjZgW7T7ONZXTQ1BkFDuVWv9vVbMZSCfeGQ+dUx28rpc
FlBgUFbaJsES7+cOD/zPiyGxHae2x0zcE/zGPtJnWVt6dT4ERbc+bRjfoxLS4lG7j/sTPpvtPlU2
XdZAKIMb3ytwLsF6kIQLJC8RIRLSaLyPcnPMejlUZQ6b/O2qYIu/Q7SSAgfV9PRO5BMVvs3t+HzQ
vZMIDBDlSuRAOuOnK2MVxdClxu2NUA6IiMWuYQSJalcV0NdYC5J3Jh5e7zYWILRdniCRlg0IR0FX
7MQX+sqf2m37eA/SazebzHkUKjBQ8MNADwrFcmc9923uYbR5LTLk/gE9xpBsyd2jjP6XrCMcZ8a2
4tXdpwdeW62DBmiZHIoebykFwSWlzdWO9iHEVwANjWGtLDSBTksAZZlKz41RMUG/wgOBi+rt9OKj
SXaegmt0PWjSq1bA1rgcWpjyrT8fF1MzoWftwfv/r+8eF0Y58XsIq6801obmmqdKKqHqk26/VPEb
hjU+IGDY++lkHey63xJaFKKnT7RkkN8bjWL+h2XX2ali4LokRbtYwG9mxHGwLUTumr/H9hlBHjZy
3d/jsCR+bI1gUp63TjQwMGZzmdR35DWAHcV9kiHyLCwycSEEo1p8uH+h8Zvxogm/comUdA7NHyUL
UKPUXlakE9sdJP0mwMlK9tkWsFTCRI9ig2ax6LdDQZwNGxaSnV5RpjLBRKldO2aUOFW8yds6RtFs
1kqRXn7fmNuLpVJ0/Gfp4QLmNGtGBQRgy6rPl0Z7jgYilHDUlgAhr+4HqruhqxttaZsWTKdQNbSl
WYeTOlNba6suRwY/wMet9cq4Zc3Uk6aouzSUEjv7Mjy9jlyybGNdmPvUYNsjaEmOrK9Jeoap1Tbe
gumRtVtbZGReQWT2zC9JsPRsy5Vv09XxPtajPTR45f2r8GidHGyL1W8euHH7DAPRnjULb4LKcjwZ
6n86sOaocmsGZpBqFYZwoUebAnyG0lOyOyGJ3rywhbdKdOSZdmhfMdeMo2icnH3wCokEnfKdqun7
PNrzX7QFG4nQO6Ylmjrae3vwDJzJQBHjtNtror2min8YlBNNyZZKo9klhwGmU7Yw8cAn0jR0rVS4
pAm/r5mzzLvBfUsyLPtyNK04huwwAF87s4UhfGp566GX7SsHVtWKLFuwXm1MHSbZ5GXiGKHyCclS
rbejtUgC9b/WC6oWGiOtlqAsmwVnZJsFaUyyd2UC0r24l3zTxys4i5x3AUBvZX6Yhk4OiF5Q/X6Y
Fn1EuqGD2lUf6kb8ys83PahisszQlkFrojhHg96RSUnTUqUtNDep+5aRamuR0ihGheJHXq1QBoB1
EQCxuW+m3LtlSyMdQ2ApmDyCnX8/YrTror6OxMBP64uY/CiPU8CmN0VcZPV2/J4JEkQ5jw1wzGUK
k7nyfFwiINq6pjjoVO3A/nlzlB5dBYYpqPD2ti8Vsyhd2rncsBB74tmuEBAWH5P/qLPl/HpGo7tK
/eQMr03OkJIzhAqc9ZF/+nq/oxvp7d9L4xuWCvv7udwESArn2KgwxX9Z24JOg8RwWDLYcey8iZtu
ltDqIU80uaQUmic1qgjz+GyEAeT2YvEu9fjH7e+QedAWabO4qM5YpckAGMaFqNORCy4uajLZclD0
UkewLc/wujyTpH0i1tXnlvWe+4xpzp4AStPtpD84uK2/AI1tzRY9f7o4X2LWZMzuGfDVDgdURtS8
D+g9MHgirkFnF7QmOfQ/GeC4lLq6zvyi3q6uGaLpc6eUqTvJLldJJ+MmeGw7Dj8Qucx8NyXzGsjO
4+O4tfgx3KTUD610yIGP2DveT9YuLE3Z3yqfLLNkNh6trJsljRW47YxmS7f8Y6JEZrn01AOCCYgt
d0vkjNvyITYb12qaByPrOIpIHpfgxFyrqTqKacGkpTLywehtRzFry95JPNPese2Jlv9xaR3YAMPm
C7GGEoKIqjrCdzAoXoqHkIGaBjBzkHXCPCdvuTVvIxXN1IynXS/qSU5+F+j6e+HW7n+sV2YsOThT
jnUPFsj0pxLHzGl35abi5Xojv1ZKvvApc2pf5eRzWGS00L12XUZeIuUxYcwJ4SBpEtdpH1n/iM1x
dYATVvE+qHyAvt5QlOn2AjnItqXaxquy6Xb4KmShGZ7O6ECQlh8wRFeXMjPtLG4ZA2s7Dp4gOpUX
Rrc+k0LYpFA6fNf1YbbpBkJGkms8/+MFTSjQyNNnparNbtWuBA7VXPZpWNa1sE9ZT+2ExXVcOLIZ
m4hMWkB4ZlEUHoslD8DNNcPDNXQSmo0+q+UocZQP2N3AQvwKYb6UpYAQivMscECxmDMIs7YcghA4
j0xwy1s55aSwxYFrlt9nev05SwD57AwUdqd/BBtr9njgkELsspd+JojSOoPXJX3e+51KkeVtjSRf
xtW1SyDPhbc1MbvYp9GO1lvUNukidkMWzAP7XLcmgJDwEioHmX1gq59Li9jqG7TjhBNXkXIgRY6o
yd4HUStUdasou8/upJ9h5/5qu9H7nklTBjPwb7v2Xd2+GrpsGHflO5npYZZFSRpbMtTtxvjc5jjx
xqZYz58+g02oRPVGOf8uAYB1QtMOeaXgdPAL9azPlJhoJJ85V4bQu1Zzz4LyTRnNoNUXYkEgkKBV
v+ImmJSj9TJ31o856ecN6Hcs4HQKxt5SUxOn5CoGWR7KaiHodQgiNipc1yQca2JMJqbcq0Joiw68
Ak34OBJFdzudnSpwYUP86sINH381fsnzAWL8ODna+J3ei0qCEE/V1tcJY+o71rCEUabTeG5BdVRg
QpSdwkrtxdmy6hlzoaQWu2Us5j019xEH5XGBjAu8eOrlRk8VwcCeRfzoJGGB8fmsCblqkppg7hoV
2VgbM6laVLscNlShC5tle+mm0t+sqPufO2WxghoI/zJ9Q6dVqOJGSOf/zS3CzzXo/NE1JLw7hJPz
UCTQYzmpwbpgI/hd038+spuafak3MrUOv2DliWTc8YpF4gbVXVv+Ntyw1TUvJuLn/ktN0egFu3C6
MhjoeNuMSVh2IC3oZjumGTZuknXk0v4JXqNYZc6wGHnFFQrQ9VWjQrPz+/yiA6GlApnYGwC3tjdM
J8BbhOchVE5Q7aj80a3Bqzc/HoM4Vv48NwkWgye854WDnD8YxPrjvVNvY0ZoR07EkmJoKA7JVFJP
6DnDpnDG9H0uAWd99UgRgqNJ37XpkjEaUCIn4dF7viSljnCBTlk+x+TVCJd00CMp77hq9Zk6SELk
k22RYlywX5dHhseU3TI3+mS4CN1jz8Ve+v3S+WPZmJDDTA7mVxzFnwCr/DNC7C8MlZZmJqRGeDjQ
JlujZkNj0V5qPN6byuzJEKHFeMdBdvzZLY1/0rtUUbhrFFmxdKTTQ/e6p96Zt5GpHXq3zDuR1vV2
aPkySfrubWrGO1MqCcQjTJAY0DjdGZhN4qdM+hgC5N6E8nRTl51gGC21nquOgCfzz3En6vDiKFSi
55exdvHJ/8dc7PksH15ZnUYw56c/dm6ad6rn7ck9emXQ0nirfS/Dl/wqbcKH8fO/BTs29wUYtuPc
ZxJ0ArwpYcf1/rPmezC991sMI00iTkeb8nS8TZxqx/gPrQNm1EzPudMc45cweimDuzGKIysWeFgs
pYTuXqTGn0NBY/t0vnbwP6cNnOgGOn5y5ldAXsTv0yYOrsHS1qh+rdaGjhqLahb99IEJoJmpMDwQ
s7nYNiEL3mLjZvKfg/Ra/v2T8g9VvMsnuY+uE1Jam6JzxxDly6LuZS6Xx/uvWFAm69BrEmYgZ0Hp
67S+w+emlRohLorhchLYTkRXRtzxsZ20AFCxHFIi7YfuDg5q18VSEk0BW5ZEt/b2YYkwwXUoP9G0
F3kpI6K6Z5tFGbM+qjA6y7kUOSe8QoNq8S+tlaS0vy8Qyw/KeAkkzx5/K4vX4mZGm41jx/II6XVt
ZQ349esgUHFh23kbx3tFY1bwIPqm8giI7AwK5njEIgdjAi/Mnraaq8sEkxl9LeGXJs6UPqkbrFLE
+b3UALvWMXvbEj0sLC8ZcGfZuQKMAItjIKD8Bk0+TRMM2GCJQK03y/r/d4qdx5TWQXhtj/F/5EN7
IKECWiymuMYLImagmgMFHubGwd7dZw4B+gIbXttlOfx4JBWlmzxDBDuTo0c6rlqfqIvgeYDHfBZn
/ZCs9u7UoTpFUoJ2KIo307WROSzLXGyqv2OfIaqWosAzjSD8yj3L2LFNlhOgwWhnoZDyw8RyqkRy
py+vbaIBIN37gCNRtQ==
`protect end_protected

