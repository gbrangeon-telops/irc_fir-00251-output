

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dKfOe1Fgzj6faSFeL/IK/IGbXRIzt9OQ8DZnq2KAQwbAq1xs/txiDbhMB5jT5GTGOpfv1lX7K9mJ
mDVaIsrDmA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cmnaZ+nYMcuVxuKDdMnuchBB9inZOxPR3/E/irYVdWCPhl0UM4JuWPFoKMQnAcsoQ3vgnwO/qltn
0x8JvlvddPokOTwabXK7+R741NBmTaawP5Y3zobRhI33jusePpwNTanCHaHjalZxzALXRseOguzG
AwGiKgpBkrzwT+frUqs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sUxQSwzYYe52m4+VJThnA3rSxL81p7y01A34NmBjYzEeDRUnhBCVE2EYcZxUZHf3SzWeAqe17qZn
+OUEYPsHFdXLy5QnKWkfeT6eelEedeGrqLjWta/XE+CwvggarDRC3yCpKHD1RObvSaidPkoLOQaz
Mr6i41kRIdL7xQbC4uLsdgEZKWh/fWAVQ0EsVnkKqE8EuxaCZ+UTjEptEyr1FyibFlRQuCcRV1zc
KGcqqHxwzSvE0/TqNDvaxlN4HZAny51ra9dxL1achi8jzJgZlO8wt9Agqbh7GQueaCXon2S1zoWz
ehgKeTmxlL7ytzeVDSpaRq2XKBPlYb/82fe70w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nlRZm6Q4mAeDfFS8oXcdcSIf6QMcM0qJWL/GpoNfKsPw7GwRrG7w5Fv9DZ3ev8dGDXi3ZhhDXcQa
Irin1hT7IkRZSupkXr6uysVtJeCdG/feYDkdTZzOR87EjbK5yer40aqraNg1lVIuObcgZ8AniYE5
0hMf7gQTkG+H4+tX0yk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HiHN8/USAozrVtx8xCHzL7SU/8fs0dpiHUe+Pxq1X1HHq6PWwlbojxR2di+cVlcr3m6I0F2zjyVW
WLu1kh2il765GldD+RCzgw8JhGbJOXcaDKXvV9p6bqICOBy5WCTf6gQ/vOVRu1kKDvf68tu0aJcM
5GW26Rwq/4L2jSNVHzuzVdgC87Mdq7eVgLL1qlhKwYslU6Eg0eOYTUfGfgCo2Z6Lcfi0atBesKpT
DSbchvClt7fyjz3I+qeNhclJOyfOLBdaqFIyBSFk+zxyw4U3h7toqFVwQu8Fc+NwLgyBezl0ZUBN
S4Kep7fupBYYGAqkU2vi+UvgcgkZQxj4+5jXGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14000)
`protect data_block
c3iYLESe5kR4iOHqk0lCFmSswGJbits5RIC2Wc4EgLJ18UMLIa4OwyBpZDrunEXHMdFl6l/F/Mw6
XdWflcybhzvw64Uy7rkZbLmb2Gb2RZeBEEAXqhFlSVQQHcs7chyhQ5KztvLEvJEvTkhajId/M0yC
uWDOD1D6szqIxA1NJII1NDGs00BZ9WHVeSQ3sR7638ZiPQFV3i1eFZ0V5W4Xpfi8cTTx8oCBCZig
4zi1R2utPEm/1GNwk5bjw+S3lOBAoIK8o19tyHEWkSUSX93eWElPRVgJdipeIbutrsv6YV6zcfD9
7i4PNWanQZLGmu+gwgN4iKMQcdNfhQQN27r5yhnFxRZ+bh60Su6C6539ejLaGgqS/FFWcx1aScsa
EhIv8QhQUssf006rCmP48uNkqjGYbk44epueKl3qlk+6UHUsftK6Xx2f96s1LkaB4uOlKhqypvwn
m5mr75HuWI1Rq2dRPTtBzs1wHv1HA48+4ll0YEr4tOVnoLFAHtK97bx3/8wUyi8lIIhlM/lH8svF
g6tehGNCPiALso6v7a0caUJfXrpltT6r/Am1JZ4f4jBM6jMqHUNn/d/E+kXJKptndbYVrM0fa2bD
cHjVYb/KeaVRWfZNcrmp1OO/gcrMdTrbXNcSYDxKfa3oXsjcw5viEcBCnF2VfL/kJhdOsJnLHkZr
gLczXvr1fDN0tvprqqUTclJuiUP14aFuAq+I6Yqj6clG5vYN0vpykyzM/pSNiYsQGBGvh1miN7sS
Ll19Zg94/hoAs5XCfiSj9rcKr4tWREzjmHaLqiikQvyUI3082bwfDn9jmHySpRqS2l37NrvyLCTw
sVqIKTh9eGipCHFDU1muMOlJSSwBD8l5jTrXCdM1+kv2jPS69JXUTdfki6av+xJTnpLht29q8TZo
to+9hHviFNFTZNs7pWMAHF3GhZre3YCmFmTthmQhNDK0Em/P7h4j7eNtkYGtL+rJiiB/XFa37x5e
ZONtGgLfeYLnnUhx9hV+vQzIQmPEPvle+WfsWKEMR3vK7186t/x+JgbPT1dHwZtm6WyKAa9dZJeQ
K4CG8TsFnb06I1/L5QDgTVEp01738fGrOZ3yn4yVNCFhjEGPd+C74TC2khGwx8YtvVM2xclcnrdI
HLE+Jgm5B8HbaeZ/QFN1dxkQE8pyV1TJ7bMgjxR90fZQYVtUC9O8gwLCkycgzvr54VpN1cG4xaeJ
uv0gH/iHgscAJw3+2h8ov/0YhyWIsVPzoSvtQvR68dwCaCYL1qIwyyH4GypnaIsJjmdlfhhto1vz
li5DXN3/P+FvARW1AFWFCfPHT8QzXt0C8aM6/iKYEAHDN2oll+kQXq4+17b7acczkngUT0AmGSMA
6mZ1BhxW98iO1TxXGOslKdJkCg2E/gIrVs/NUOyQUR0CHaNJMlUeaWJTbTuGxBZ5fbXu5UZM1iGU
uSYfeG4QpsryVH2biVqlvnHrlavA1bVMpiMSkGz5u4+MAW2m+wkruxds3R1z4qyvuZgtAfFa7xTD
q1Aq1bH72TEWUTXAW1XBR3yZZ9mGlziZ63ZxRDkQy2kcfq5Eau/cJcqHkb2n4GtrxwizahquCUqA
m/AwGPyAiHnK2hNk2MwytJb5+69SVp0nsNbrhSZjaVXGi6s/LC3vCKFryD10V0EGdqnA0jR5orR8
TLzrdBFNrmYqJppAkSF74/JsuleyGzFbFK7Fzl5Ir5xKAajOEdWHzxh3fdkLYgnx8XRzYEnqSf5Y
NIeVyMLs4h1qRamb7ET0Qj+7d2hO27MfpuV9K1O72I7RP31cozaJZL3HbpzWlLr/9hDtD/xVTlBp
UdywVEGF78iPmHFip21SuGSEBvo0xpBtL0AhaRkQbCxtBGXz/9yNPVHMaPFNYRCNiyiJJY4CV8Zt
QMme+a6CNRRL/04Q96N8g/76+bMM8beOR4XZHnYwhiHxNSHJk/1dN5NT+ounQNwn6hkfrVeT1JKm
nz4Sv7Kyztkd+ZgV0h41M6i6MAVMM+rHH5yeeEVvCP0E09MjYz0dMGLNRBxlep7OR1mnU5bvxyfM
cvJZcks8PQt7wSz3gxTBtKr6uCC6oUtCY2HI4bS0bKBtF6+iuQ233tv6xVum65qTsWOJHSKL2AZZ
UUQltpz7igAjbzyFBhRP2AxjkXVG4Y87AsRQFnGirvfLyhuBaNtaYUkDETW674q4kBY7dY2qwL0G
aNEwefFR0S/3ApE0UlDU/POlPL+ZgJQBPtXQ4kTESclNytgzeUSNDmWuOPWaTDo23piPZ6nwcJdh
E7yP/bmFHMfgouJEYaGGMFSFxsHcZQzP/t+9JYw0Z9pnMIdSgxcLsX4GZyFqsW2dNfCaSEfNTBfS
C5j9L6JFsXwez4VwKjiU/FEl/8fpzIRF4j9ON/SDSbLHKcGOKNgOS3lieI4k+XeeqA5xrXz2Qq3C
Fe4v35IhEqKC1I6DPYklHS/HhIWTy01H0h0ArrRn2dhhhq5Kt3vDXl96SdTcjLXbzPRUvx8hz2JN
CKZRU+FDx583lsPFo2J1KjcGh40rls0/OpvBX4dl0aljhaAMn6TJlMIfJrwdKLJXo0zto5ld7K0s
aS9YwP6l+v3OCCzoKT4TLpq8M2wgqcgOKo0IFypwtizAOGhsZ7pmA/fmD+d2DEJKe77tWRAWlW8F
6RTtqHYikY0+K8M9Sk3Gb9vp8q0lcr/eNL88mzz1OscZPW/xeAJhvE3fUECSVkMAc/DE8ErOc5Dx
/1doJ0YQUw2Ze0REZRQCoLTjeypOaRJVeGo6OsVcx4zyCyQxHTp8/24mdZFh2r23iYtybPc8OyE2
hbKx97X3UNkMAPXElEFZYtKTbkwUiNWHO4+/oa7pHNbPtU0BrF8QnbNHlxGXX94cRAx1unja1509
Q4HifLUQBrrPVnXcL027DUbwqjOMMc0HSio3TQmv4RpsrDYAOiAtJR43N4uULd4CiwE2BFEoC8FT
K+qW3uSBVHLzbdgzcEQ+a4q6NWtur9PgtXwusyFm830kTh9sPesIgd2EjyVlMu9pQ1PY+QSXaZ9q
U1+qs+KuemELdevp0bMz5zYUtlOr/Knj054u11ABejWWIA5DBz0shH8wjtFJ8w0b8lZL/owO/Nnl
XBCZc0XYlnM87fOrvgLlLyKdfS45l1NlR+B9U3kZy7Gq7+sM6DgNMpE37jcLm9ukYNU489LHPwzP
25xb1dWaNy9ObNfkE19dlV1jTgyssNNF60d0CMBvxiR1Q30HiFtVMU0IaK6sjqYQEygbxrvIpPb3
QzA1ShE6mn7W520G+2qEsajZy2YOF+dbP7pySTy/BmADmWQuZIh2ohN6TE0jGywjHwF1bGqkS1NW
3S514LlPxK2PpkwVPTNCJ8GHzwELE+YNqQld45lqL2ETpPSqvM2rfP3de4gvvSagbJI3sObWKCS2
BQPmXbb5JqvcBcRjIu8VZvYKVM0YE9Tz1XSLQ3EdRUj+oEVFbWzZL2qAGI8PkwXgCnVSVDS6+s5z
3hQsn1Hyn21d/t2At8Wh1CrBmi4e2Qb3cumaZqIXmPTuPhFgu4Zq5rKSIJRzGIaLDIek9GfBR+kw
fRFPKLOuR4DA1H5kvtRSLlmT9j6i2iShUgDErJ7yiLtMFP+UesN7YAUcqb0xoUDxq+4dJw+8dIs1
2ewr314LjIcxBjZlxkxrZ8yI+7ehABioFpFM9Cjp7O+Gs3CJwwm787s65ZJweo23/bNwoXhVIGQk
cjsnUB5lNZ/zK/oPBBu+k6Su8wEpZVWx2LucsG8eTJq7O/TigGk0a9aX14wcZCIKVF5fuSdWx+o8
4Sp0HGMeR9tiz4WZkH3pFFgNRMAJ2pzbpfcwdXxkaQka3EfrWNqbZEgc32wU5fRY1UCN2d9aYctu
UVwXf31n7+pz/EzGaB05uAT+N2HeUfdNIc0a0icKzHCNgd1ZwFlCyCCf2wQziVVGmcJhIlDU7T4o
NSHRGoPdWJmwJ2mK+xIH/mghLuL8IRWu0alN++qBV9iuzq/zlyYEwu+zcm8jIZOZJo/sbD4lP11K
dFGCfYJ7nnTcVKbwKhxbqDZwUzfGr3ojdnx5W5tkOPQRZLFw00gEF84WqIi7lGPvW2/MMwmRPkI9
MddZFzaunLxYzPvJ1y6eQor64PPCoPMBMArHx+3NEh1LPJYWtuCugDsB7ypMZ6tI8csMcgUqKK0T
pg4EtUng3OW21spGD8uKBOsZBwN8yjKfNrZqk+ln0QctVV0qcvS3Eexc8CuQulmBcor7WpsP7MY/
SgrwKKzQeooUtP8fcqeNQff3/zxsXC1oky5UHN90iEcA/xnZtTwY/m0l9pczUkT4GaULZYCA8CIb
F17Ak2WMuw5weaoCu6ShygI3sQeK9e42eYBSx6pZpEEigOqey3uCVkLi0prf9Cie4Tnv49eXj69x
mqf3uafv1zyBDJwyRzaK4Okfh4sR1qCgxrSyzSOYjogJ9BBgKUu41gUcey8390wRxdxfhsHhXzKz
umH6U7vOfqnnTGMOF9bmKvhfV5FYQQziEmCPa1qgf2VqWaDrmxQvTPC/5+SO1tYSA+EkQw9QCUa/
5maDCpWsJktknuvlp56Y8Q0CT55o7kjMgK/cnDyzi4s1uJkjCHrcYnPgWklLtLJ26GNKNnrimULU
XjawsNcP8FmXFNXGb2QkuzSrg1T40+RDqNDK1DsQ42RonPyZDwKP5Ak+QnnEh6j89qvf19cNicvU
uU1eD6Pp4FkocSbK2vFWlPdLCNZKxWRM2QW/m68MjNYnQ/qAsDfbXbgaeH9gwkSz1BrF2pnO/TGV
1I8WEvrD49zHa0iF1kNx4HdS8NuPAYMz9s1Qps9jctimEK4oD+hw7Yp/YF1FCB6kgJojZHTu4L5S
x9FH74EZ0jaICmtMr53Fv2NuP6SXYvWgNuZISc046Rtp33QPYJI7k6uddrsxb/B5mxGQVz2I5bH6
V8CJYgrH1P3PxvHdtDO8BDQRLUpxcLk1fl0Z9Zpe3jFNmHcG9wkJ6lR8JRvBaYdeXQ3H8VbKp7e5
9E6Tjw5csG7QHaL77IJZXkgOrn5emT3FMn0CRk1VzAx9icRDwd5zY7hClq6qx+WxHAwYbXVfec6Y
9W9SPqXDe8Ysj/B8HhSOPF5hDVXi2SlqxVXCzPojiBLq2T5Z963FZbdXz6I88xpv0myg/prDlq3a
3oM5Z8ZNgcKwgi6jdG+/BCoZa9uZaR2gKVEkjN/oK7Pfy0iTI4OmjIzBrjTJziEsuktr4niICl+N
/k3odClQwaFqubjkwbgeOBeV2TPxSKh0RIxZJecKUXlHbOcj1Dj/4ZWQ5NmcQD1Mx6WRL6ykbq7W
CD+jZnTORxod5Mq2Oi74nFeAUNituxwM0rG1NR8PoGooaXgHJB11BKzcmNgn5x9O78hH+fl9XE3r
5B4P3mWdezBcSLF0YybvGXFwTCsNQU1wPrxu4Z25mBjz3PK4yWPb8m35KCOMtshkWwkAwxbzQcv6
OHF/wVYewNWnSQ8x6nZYm2bapF3O1ZXo+3u7OLSEWKMa4Wy97jU+jeSzwWMNcc7E85g3LNXoTv3j
mk7vgdDXbCbsrELoRk1vyx5W0DK4162ZPz+Onkc0nSMlU39UzHYkZpE2vfTlnGEHWyyOuyLCKRmm
qCw99eb26VijEgBseAd/hix0nUZctOhvCMep+raqRRcKCGPijFUkN+bKx+5hl/aylTIbq2+pzwzg
FgHI7zsDItTKH8x2eJXAGY8QfoYFeHl1CtACJ/OeiccwnoenEZBKcrpJ1vWsIsNACGUSCpHNjtON
DN0Lss2kgATFoq46VDVkm+CnzgLSlS3fCkzHVMAZqbLQMGxAGUvXnE3PcQlZiT42Ho3E4/oVA//2
8q9qPQiIvxQVog+kWmt3J3MPsuba+j07timzs/CTD5U9ooNTsQlZub1B16Djub8/HNJ1pkQL5JIL
lQnTU/isKlDAFOGf+4EI4B67VhJZh5HRS9p13/7fg3FIxB5SLSX5+ExdOoqJ7JR4Ww6xr/GUuSnc
pIA5S2UtUPDQHEmAB6ngw7pu85SR17lOHR9vv0Wlt8PWeCfg8hl6DzC5i1DZeE0DQQJaCDxBAN/U
o60Fw9/uCisXhm4ep6RgXIWAwQEkL2NjYbtUVmwzx47dvoo8SwYXpXfTJxKZxKlmwTNDr58yVifL
t4YEd2hPCa00Lu5EZ+d8DpgzZfa5UAYTZBxHmsnx8rNdfW3APQrz/X3dzhVqF/ofC0bAOcshGMR6
wiAX4EnAx4gIWvxEAtl312yJ5ei47pXGmTgZE+MMvEOM/IRISdscrPtuB4CwbTpllc6gj7WaRdT2
jm6Tv8U3Ckq/mqlpwfoTc3zgA30CvA3D8LywGsHE6+wtjMxN4vObHH5kyLCLDXsStX8H741R/PaJ
k0VBqyLQiTOrcjIQQymczlHstKzzopga1EneXxMgMxaktYupAOHpbuQl/dKhgsRh7km6PsexQDcD
Ze3fEXNr4MYCg1uk4qeS7VwBNNkLLedAw79sw+IGD3BpsWtMSqdcT88vnt/GhfqX3LJOQg2HKVpZ
fEd2SxHX8qqHdZpkiC1nTLTEvixOEzDLqfc3nayMqjWO3IALSLCEfL+bNT7f4OFMF9nzTDwCMax7
X74XiFdqfhyUYb/9InbH3UL/oGFz4hdwXxfT8RFW6FijZLFhUaK9T+gG0XY0ngkPfXjL/oBirpsJ
m3Y7ABp9fks0o5aF0MaNwoZyFv3P6bSfOugfwMUywJCUZ2hSbRFxHDT5DmvT5xCdb+nHUdB2cuey
MgPQpMQ6IZkMX4uuveaOuVG8G7mCCumaj1JFmzlY+nBQxG+AdxRh/aDzlISEx/D0hkPDRf2k7FEo
X4iKfb/Ge2crXXmWn0f3PoyrB+aJxYu6EieT+OdgbUoYLEtoNlVM52TWVfsCYkuqr1TKe5Qdj/0a
OPtr83zv7baU+avXGFiYcOL3LL2D0ctXHknyTW4jcqe9IxUw2Mh9r+rtCqMlsMQcTMAJ4vGSf+9u
/leWnphiMdxHW3SDkTA4a1ltUWwzs7bsJoOg/la9Uz4KriopCAyU0bGziB5DkhIZzXBSw8drJpp7
TRlH7kC5VoNKxsJks6YKbTZXc4Qt3cTjEqhE+BOEP/OHpVyAOSVUPWY8qTwdCfiLK2XwGBchr4+2
B1MvMAwPNm8Kfm9b17pbnkRCMSH30NPrGWekhBHjbhyBV7lttgS6eEa6zplpuC5KYoA/UTeTM1TM
bTgxpbDajIwCQG3MMjYA5kbZHeXs3WK7u60YUOc+LSM9d7Lzx5rK60tN9utvWn1M6Jk7MvFI46iJ
dJaMsuOV5hGL/kDwSVExli1TrchrH2IrvVdEjj9D724W/So5EL5BhsF9qPxf3cqGHi8Xoy3ervYw
2x+4lYwj1mCB24vWCmWZrx9+yVENL3rvU0G3p7l9oY4+nzxV/ba/HZbvCgnOM14+/fdNHLlfz0+D
X4Cg4I05OGJaPJ/EYiCJMOe8LhqkffN4i8HBGCj5gZWKfE5txeXTXiH/mBtco2Hadi7qB8P9EonL
GYnXfDg4srA9vvAREwCstUgQ848Kvu9pQCUtGg1An+oXPCpMxNujNZnQIGe0AWgF/Qt18s4Cgg6H
207GETCcrBpRWObpk31sF0bKViiDWTOXwBRF1mp78lb9YeeMNS4BvtZJsr6oiQp0FeGrl0xHJ0RP
J/1jgxuTKDqEaXmjraaUQ16SY/VPZOso95mnlceBUX5PFzRPJoSe1ScV18QJafdKQt4dy2p+NxAy
3rOGI6ayXoYqdPLEfCBV16W+shI4/xtt+ccvgjfpbo+F6ojInJJjKmF9UoRfyHcZEzbIIZpLN50u
ytmeSRMFGwlC7Nssaz3B4Dtf9yf1g0C7XQgPZuPjjtzF3bCPAwUL8/1CasMR88HAgmIZ9qrJC8rH
yoL6o5YCKVaXO1SeJtVYWI1OhM46XCQPuoQ6RspcrwwNLTFeg8dfM/eN1M7+78yySym6/JIs71rD
tlHGa5tyOQ91pkqy4F7/0T/cCgiMotE/QAxuUYB1Qb5qL34yyGoWks2sZRumRgt+ZuJcuvLOp6J9
e7pL0+PO3LQG0AtjM2joFCwnXiz4ekJNsBFAoA8KOVexpUMZCIj5YG94uLdRLv6JX4BBLxaBMUE+
aawQLROjWZ+K3pBrjy9V9B63cAjIHrvjo5n4cAAy/VsytVZiirdTR6ohsgHu4vGh1zjSQuPxTiL1
nvNpYtnH8F5kKLCyH3S9wNP/kXN6/lycRbykt95zuJre8t5v1Lb08o0MFKV1XRIkwzJu5KGK5wv2
wBzlkApxpsvfRcZ0/BLM65Gn+hjW/bbA/LEW+kJO41G0/mLLQhu+oSoTJGG3nYIM0XBT2CRnAUoX
UHHEKs+nQNtuknR22z4OP6JqygVi2C3Ny201ezqJcgFMS6fJF0waNrbpSE6Yu+FYgyJ9gKRC4J18
0vRAaxBYklpPyt+BkCZso70b6GKwti1CYcodL04Z4AFCsI8ItMvLx02TW2GySgy3VLNE5ijKT0tz
QdFqh6DucJfsaekcILK7uA0zDe/amn43yYZ4PZFbZ2riHaXpokAi9/iS6DDu0HidPFxhDKwPqarZ
/TwejjKPGMyVKNSVfnyO7vLgfz3SBMtaeRWx/ezmFj4CHm/9bd+/cHJ5odrItc/Xt8z5gKh22zVU
j5c783wvL47uBNMwSiT7jfWygVYWS8LAzLOdb3jOvDF1irZ2MqJUwsh1LZQTXy2qZMXx8BwxhuiI
Xl092vZTjr7y7N9YqUJ7jbW0p+ik3QaPsxCrmAuGvYFRtIXRX+tD77FFbXd99uuFLvPJGMCFZWXv
pXRU8ltXLJEvNr3ELe1YzVPAeU6/LNn4OWQ+T4plsme8lV5ijMNjFSbkWhk4cd6L9zqGpnirrEBj
RVXVyf14fCzYG/vIzGw/FArkEi6aHT7czu0YlS9P9B/yWefe1Y4oKKa6VnPBzaAGuoMD7t66rFIz
suOGE33rzRuY7iIoOfv4kc8we9ywMfY9mnqE4i66dpblIy4FCc66DAt2DmiYs2v7luBYuoMTh2xL
YQKkqZuMbKn/R42fn0UCneu98uW0w6MYCvFSmC06Rl0icXt9sKU0rdkTeIPHkWky/CCVeTCh9GkA
le5nYxJT4g42qmOJ5oKRoWFFxrKPIqkjSeInFeUig8jB9YOFgFC/OiskJ1ueqWqN2A4KV3WW7K8O
wBBr2n7YnyXoeYg8bfuSdab62kl3f/G7aaoTum3cwv/ZvYtPeTwe8yqxoUg1MCH91SHD6wozTRZO
POL/udLkE2gOfSxZdg3oi4lLlOv8Ym8hxRoPFzIC3jAWn76lpKy7G4fisWBiPouO7J4O0lpUMHWd
zpfvMFey3/d/KCkTcIqfy4y2BlZfKnTUI+OJe8L5eG+ZlW1L5b76OuYM06mEpXPmImQN0Pd7KROx
59n2/jsIRUuIeu6eyGU9dS3Q9uu6n0W6CbTrQlmPuTej5GOvoPDZD2IhRKDrHmrU9XCy0GRzWMVG
WflV80auA2CmuFzBU2s5dHbaaK5Cwsdve9jFhw8JL1MjDhsAZfNffPgLgaCAXUa2221aS98Z4Tpk
QXEDh+LtLWBJepMYyGlmv5STXv7Gy4Ia2Zu9antbiU4G9oENuTYBIezmo9yUSsPwxB5kPjdwms7w
5ioatrkeWmPbvWmDlJ8X6NmLFDvEKAl6KyHxUJ5zHoy7CPR0z6gOKHesy3cyzsLMVxCQRtNVSVuV
YIQYVbSicMHYd/egMCUf3xdr1VUA9VlL6oPPBza/fDpj1WWLXxy0olEWVOnobP2fp6QfkClD7itS
PQkBsqBcEM5yI3gzCuggGzeaaEIvcPTja3Ii1hX1+1Mj0dyvUWl4qQ6/Z64EKOeKStwFR0B4j89m
hz+WiApErjjyfTMxPx6Vj1D09abFVwTkJ6v+89j1lrIrIgmJrTHvGpoCSEdrzfGa0C2Wb8bkAhDw
flVcXRVDZOF+bQNoqjJq9q/mpW6VdZkb+qNlEmnl4NZssT/dhVvYBJHadi7gOQdaDu8xUFioaPJx
uGppZ5Mego9FGB9QMuQPW2A6Y5w88swUAFbtenb6n9rmFP2SSTmKzSEOHDeK0tdBnkD1lW6PCHQk
kV8x5tJYzh1IBNbccPKzrf4wocrSlRc2lHjz55Y8IdletEzcVuDa46XqmFG4fX6cOJrjgxiOxTY9
hUQJx6fcMzY9NLoIF/zK8+6lQyK5TPHJgQ6xtqdfqf7UydsEmUCUOxeaJR6EZZLMz4LBP5Ym5jW6
E1oGw385EA3Hp6wHUz8SVGGqRvtu510slPW+NmsprQ2RPwoT6cKvJmiLZkjSMWl+9x03OOM58zeZ
4+ySQ2RT98/m89ogM+snitiW8tDpClJqsGb0AnZ8F0WLWKs8BwOWlRkOQAMP3pXkRlONYFrSKb60
6SvYu00h5JCqRDjq9RWgbQbJHx0crvsyFJtoBbEssmpPV0RkOTG4W4pSMsIOhAnqVb51zJGHO1yH
pgZVSTNIrV0HKJIS8VLUbUMa0L6TYcfW5QIlRdLSGGIfaCnqT7uv1BkAeGrzVQwmrc3DcgU0qt4R
y4fN0m+10SVHG3YL3A95ivE7DhtZnhUKdMGtmhJaw5pjcVekXEyCB5oDqSkAuc9o4c9r3cXO2GJk
LUh9PeIFYJtGg4M5LhTjqMU9T41zok+0BkENWJn4ac1hcIAeAaLM8ulH0rmcpwB+r4N2N+wVRXWq
xABiWdc3VUvampisUvwVHsEkuS4smXdc5AiDd+Wtc+XiH4ZNwakXHQl9lWPKi8FKgwMUv7UPqQqU
ePcia4O1p0NuO4bLiKHG1QhUUGBOzUlAqt3rxXudFECJPh7cnVgBIz1+4CLo3Yj/Ybf+smwqOlkY
AfCJ3qOSyOzM9cC7/gnWu8K7WJihemBs3DkgrGrjuHfaxXbbauONayeKmpsNbJj+ot2wXze3NqHf
yc7KlV0uicr29/+sTFxA8uTCV2mMJBMAIgcV5F3fM+bZRck+CtmIHDOQiJ9D4K3vJw6SJF5tmVa/
G+V8jFMeoRN8lGWbb2Tc0tZBxyOgZ+2S+Lf24x0l/YePfb8Wt/0+c1JdiY+sGXBSu6OeYl29Uymy
cUChU+TLXhvJE/uZ2NkS7xEdZa7nNrjpzsBvzcHtoANqRvEDWBb2q1rlmJdzg1rqILySgxjmThFk
6sXDGihhT17s7IV4/NaQHiAQqBIVI3nMHx1H6MNbn/e7MFipjlPBFya3YsY+73jjsTIJ9QSYQe/m
Y/LJJsYQZL0IzRWeZQmmSasWe+WpuCJsdhQVFMozpPTNwr9JmlT09IFFagom4SxH5uxJo+a6V/8d
UnNGUGQMneYo8Uu8bM3ohx9tyzFd6pBIz6CShXUSIjuSYHpqn5jm9ugBbl6YPX9OfCgWY+UEBi0y
HK/ikV1024m+SvJvSqW0lMICCu4XYz81i8vfYLSqCSFGo4UoSWqCSCHBDpizuoHb/ilK0BTutF5Z
QeS3RU6zPwHx/b/cIAI2Z79AYknF/AyP/gNsZJJXx9BmEOtccz6RR8OnlughhQgpmx3LXJVu/rPS
8Ejqr5RZjMlKL4m0f1WwEzGcfbAqdGkAxFcR5sUNAyOHSJMYMRnpm+IXHT4BgykFtTD3HFFw6E7Y
/t4mWZOP5/NmmO7+6SZRpsVnyxgpCM239SwJTetFHwU8YNbgRBOHyefB2sJgWyE6LthO4HjYMsIE
CL80M7NAPxsUyXDhJ4BIZrXqiV2OCyyHylcBWeJ/6I5X4vtPvzDKdssCY/lQzQYgmoxJKO9n5HpA
oIsmG6s2YBLHVuGL2r0iZrGsaU4Kd20sNOr58kcqf7GnYA3rdo3GE8mpUuaptgQyBi9z8oti3/Xn
MAVB9+pDK15zQC400TCWrhPceU27oHR3byjhUjtD1inSoV1OXpmhbXEBaFS16c+jWOAT08YxtAJS
eycJvIDz9YvHUKPvQmxXRNKFZbBPWpH5EjJmOlZ4joAIhSI5lS8DLq8EDDrQn9oFuZAYQlNkleU4
qfKj93k0OPdlnju4avxbNE6fmJ0eL5iBXpfPbAr8EZwpurcns1en1yfuCRxkOB26WUyoqZPuTdYI
E5srzIHgIOTCK669sE9U3bpqmeKSPNBFXlNNFlRDHUL84hxhCli2c82GWlWB8GOID5HFs7BNFIZm
PP0xZzXZ9JvnrwDALZ8ymuwQ6dI/yETQl2y7jhiYOM4ANZLjMegXNwGW37KlliyPeo/9ycMzr3AU
Uog4HQBxFOU5WA4iyXweqi08pZlMnDzozgemsJLU4o/nz42piJlg1YusO5oGL4Xp/dfzOX3MB/JF
AvDVr9Kr0KN72qvUPBa9Zdh0p2eaj/Gm+sBeD/5j/AWmvbdW1BF8lGJtG+lec2ECg7+9Q/B92q3A
vbCGTtEK9As9qleks6g6dcqjJ12c154tw1oqgcl67QKS8hL9jCpr0CTKMcrKa29SkyChHq/i4+1u
iM7+1ClXdTeBNmGc2NgeFp9QUE0IMHmOZ6K9ar6KQsu5J6yEU5hga2+rkVZOWL9i1Q29crIOpfFG
dydWGsQIbW2aQQzb/bWyIp/fL/x/NRah2W+aBZ+27YosjuXNlz8mNPrecGqvzue8l8O06IblKsBl
oZ15h/2hCN1nNEwrqew2zFLgBFw7BaOZcl8tZsRJZA0b5LhiOMwiIY2vSpyI+jR585pF74q1qW6G
Dkd3GyPsyI1bCg1tmd0fE4XySM0wpJcPHn+uSWy8d324ARfwyOFY8m/ui/fmqdnqgTnve+lm8fdz
7CuDocg1urmALoJwWPmtR+vx75R9CmtesNVIUDSzijT0YQ31SfnErPdWsixMck6wiSYMRSHENk38
JD5XEZFWLG7cJYgs60XqCxt3e7E9eHN4Kpu0w0Erb7G1HY1NHkDyTk/Zs7J0t6O6cfzFOUhw2i54
OqveEZpFH9dChYLz9ON207E5sE+iUVQp5n/Pbj754oCZWGWlrgHkFuBrmxf4xVULvDPD96L8xoif
55fSWgxzbROTdxGS4bn1o9V+lEXncKc5utiGwX71h5gh8+kHVXuYKa/bpkEJ9RzRl3Qr0LYcfFJy
77x1AZIXDFECtehOnIfjK1P/BQcXmCqIqNcv0RTKEFFnpstapEUltfBKpf6Omv4II46ZUsqVjasd
JCiTxZvxAhYJWnZS0Z04HWTAUtZcn10MWZwvk02k/DNdNEtrRoNz895OZL9H3PL77wTsOvcO4dkg
cxXIZu1EqWLvREFhvqfpYAeDRY0glTLxlE4tSv9EGjzslJEZ1zapmzfkpFM2JG599tGpmkOeb+2C
I2w6yeCbJ4Wq03ZogcPf1Uvxvqq6TYXpCiwLciru/xpZhrkHu//vI5MrYkx7WTvJcEBYvz35EmXQ
WyTVfQ8MriV0qU+v3ls9o8wdNsC04SEOHET+yAHIPwpNoslFi0QyGoxNilg8CuuSAN/B5eaV8t15
ec77WYZaWyOz/B6mVZIpuB+P5UqtjWOW+TW1W6dka6f1+jxj7mcaaJKd4ml2kXSHB5FedFZreJKc
9vmQnrtojHSdWDLoK845zI2HB9ZEJx/HHKs6F/we0ORuIfNqREuKimtyiNNhMrC+c2jjtI4Z0g7D
pG+0GQO696/Fjvlw5YD4fgUjg4KHw3sgcuBv984j2Atf+5Ob4HAPpC0dzzhPpHGojCDRJQXuDUIR
0RK82kItYfKjNyOH79AIis1NISBwgYo0RkyqAmnPDbU7/boYIqYtv3JqgGG2OBk77KkYBnZNt9rw
+kV4JTSIlIqYPkyzAmdH8QhF17kEjAYJHeK7MaN/nm9sIB0yhYodTc/YnjdhuVX3oE/3ycbqBb5/
SVvTA0S3PGUfnA1W93gKV7Lg/7ZhXPYvdEyrw66fpGoX2lZmmMuM8A2kiNmsdDEv4GYVLz6lOqw2
MgVHpD2CnknpS84R4f8LawFGAliSYS/GUhC2rZMuhgLiY2UD+Y/IiwB9lfOEiuQKNkZD7M3u58ej
etb487N87oiSgBbjktSKtpeNt9Z5tSpJa85MwtzsuJy4XYMReGTTymwTr2OD0t25KPGqi/829dEN
cbwpgNuZi8vvEmXHVLR42uNE4Z7Uta56RCnvFYv/UYHPDWqHoX9OS52V4r4L0sjAotunR3NOLQTq
2vGeoyGOfRD5IeE/nqaLIlBJL5NzZr6uNUQFFWtaps2aOAYxMf0AEvpoqZ9glmwOV1VR3adFNq97
zus9HjDp1gHUgaezPgtsW0D5Ppbx6TUv+w3Q8TVdv/NNiV17r6BlafdffBZ25XE+eiObndE0/nEK
Pjk/33f4PeaRIDpd7wVw1QRBKlYM4lnVfCC27jpwnQP+6jzVp6Fo7/u3J44tiG7rcXCuufqGVMZQ
7mXklzFXcQhuVaCK6g7vcvx0stV2CJK4q+O0kH6PJd1iwa7KeZuViEctZHJaLeQ1ZTr8Gw0BeTMZ
8nCKR/pDHGjo2sNmDq+vkQwLGFLZqmG/6Zg9JE164oiefxjxQjaU+CFH+sg9+7DRCW1O6zWIDy5V
kI2lKk1geK9UZFEbaR3jjYG8SdCwDh18vtlMEP30AJE0xo40TWx7DIABY7ntxQlqrzPmyOstkt7H
f+PQgKq8InMZx3lihnX0qKdCxRmZNOnLwagUxRilttKNjiGge3YH+Sf1rmuZYi85t77r9rNFJFq2
4cSE9eECrERKeMLdnew6yZqpxhiBFAXxGUhxVj/K1MErISUG9FJgi48/gCelnY4gMOg/AB8p13f+
vIjqzHcQFlm3sm8Rl1g1WmMaqxDRvY6oA2Z94hqd+AIn/x2fpFrNkOTtvtzWHDzJ/DanwPJw3/k0
s8GGv8AHXbV8kvS0wyJmJhbQIQCt/lJmQZgrSh7xS1apdx/ipaigtasBVS82nrO6Skh/K+JpyBWJ
JSBlCuwdSGuJee5R3PybQCS9KTwv3sSdpZ1z7YBVzxbmHhxsibqGv9Vgkyb15eKTuDgqFWegt0Tq
1A0a2qD7XEbYNiA7YK3OeBdWAcsTCCJfkZczH4y9tK8cV2BJk78li46UjpMj2YAVqN79JLzKP8S4
wPYdXtuH+AC4y1B8e6CSBJJzqG9qQl2BPTjLBdqPyS4IWBpclneAV57wQz9BEJ7iPkryXnmF1rk0
iiyyszFwJZ7gWmGgiVGKoQrGDfmrveKrqGYhLxirfKSW5nbR+pnu6a2HySwVGkj533OvLgEqpfWc
Sr1r0PYHtujBzffkfpgXao8CqW8XRXCNeuTYHNGtXKtPeNobpcsCIvQ4UfRbr5pvagp29ai7grt3
gifkXrk2NIzm0hoDDDgfTYxY/n2Dbwuq7jRerI7EXwKULitpcaz5IHk8Nrm4pir5GqOxocUIT5hO
ly3Qps0Vj+6bSns7JMkfwAcd0/Uxj9F5xZu5kPIccDLSrXGBq7NYZy+Sga5dGgobGsrFrRZpX080
gu2ckV9T1pnxzHZFNZSJWehNKOe9FIp1ZRb8JunUpda8dumWY+FR7saaUWrMNwSSaAqDyRHjvM71
d87HNTvfX6clYRxZd5f9udx3kR20BzKzIGltoxSV6Xli41Ncyp9HSRfvDoQykXM3oJH8eaV/OjyK
KIvS3sQZxdZMGEVewmeNOmr//FbN2xqPRWi28G+g4NdryDW6i9waqeVsW4regaV0AOklPNqVFgYP
SuG8nc76ryOtlESsmAbt+2OdVQcrgX2dUzIri64GAto9IV7Uy1u/aOaVl8q/RgUAgqP5TvkdRtPt
aiIxeZ23LJIfHJ5hpEkm+NS+awYeQMox1eDBSB94NC3PQuGkrXUvs/5Rb/AiB+of6ql+HUMdZE6n
pWsumxWxZJc3kS4YSkF5S/bqz8zT1EXaVrNzhlnETsDC2oLYgod+EpIF8RV2Jddn552SBokCIM6k
TBbmU+lyxzyQ/PqOJFjEl5e5+Ipjr/YL46K6itDdLeU2O0QkuLb1EID+qqFWbvORJuahu3FyF5Kl
FmHy7ipbiTtkeZUewh5asT+eIlT4/sK39BgKaHnWzQmETuEdYNFXdB+zs5YnsjWU5zSPnNA/sqdv
/C7BpMV71/QQwMZR96wdRx9hIOtRdZBfDdkObhOaSbpzId1FwIjAFx1+uHPWkofmH5WQW75kX2oE
nZ5QZuGhYpNAWL5xJDS8C6qisPxlCrys5/Mn/JQ+vxCSE0btwN2Q1GgLm0cvzinvdUgZcP950vqY
tODWFClNjHhMZ1fREDKutCJ0GMUnQzWUfyFuTn9K4qdadFyO7brq4xkKaS6TntP8bf8avPfly4rc
BKabBQkvZxfYMxB2C0qEUsxXL5zW3TnggLibq19Lp4ka7kEtr5TnBq7p6HxkTGU9tsFx56um2y02
kjotTt/Tm1fdhBcQsp/X3X7MD+iZUbEhF9GuWMms4MvnYNKgivKJV0Le6RlmHLkpX0t9ZIGpgac3
CBcR22qF9F7qO6a10UxOTjUBW0mp5psfDWiPNNoWAPkLHteYRfau4fUw9YjMovADINDf6gd0ygMX
us4kWUivcTZH6Eotb89xFM88yxuE6/DRvbx9ZDb6wRPs5g5WYHInfAWSNSQxRx8O54HtTgEwWKG1
YEE7NXcShyKvh3lcByBfIOE1jE3E6Ce4rRZr78ZJ7s4DjVuk4ijAJ+OzaloFGRR1MLS4ba/IsGs5
2UkobqzcJurlbBhNms1VkcpppovNKkNAvWQ996yCelFq1fla5Pm7TXFNLxzI8Z2DANS/OfSdsC1Z
97wQoFeJ6MA+bXsLlFTVZyREC/uje9fPGXGudz0Hy3nQplLAyG9syKATA6FHw52Uj7xokZaov+ue
khM+3HGfQJSTMSYDNH+Uie8QNPiq5M/MTTo+scBerClYIXfi5QfpmbmOw5OIAQsQqzthkHOaef1O
jg2MwpFMyvv72bQM5U8tI1kAhZwZQyAdeF80ekNkm+SA+r/qOpvwNNDrM7n9YuhKW5m+MsnY8CJH
29i9ce9KoFMDEflftvDMshSfTXRQqArFEAot8g6cflCaP14bmjxYEgqhQdXqRh5z1zDm+cxorbzI
DfVb1PgyW2m3BKviNwzHGdTODyAGLNWBCbNGkjAsjwGQ8YCYvN4nAYItdmHVTLTZNRT7xkA8DnUN
JL5LT/hTcx7OjTebOGB1BJIgGiBrxA8AoMf6g6+fnAD/LZVF/DgWV7ceJJy9cSqiVqyIyG7omig9
cMm8AYaE3z/RxZXwalEPz7+7FLinlIA3+4Zu9X+I9obf97tOCWxuvkNnlccK1QiVKA6q5S8cIk15
b7KDzbxHouIRJsoSsfNTohUx9jgq5fw/5yp+II8Mep2SUT6fcfHdaIDrPihoOHuZcK1CAamHP+nn
iRhpeV130T2CH0mj0/XGiZ/zdRE9EddCmrWzpn3siwO3etl5FRhjdkLoDEw+Sjm0RbjjCkPfE6XG
2HOXRXfkSxSYIqC06DrIQReBPhqgc0rGNkrcORoStg67v1wby/Wb61APLQopGvldqLlTlyXbFCOC
NW4Y/uCX2hktKKxXdfxRn1+0jgyRmTC0QscT1/SzjWfKr1shSsFH/3jz7RgFpGczKzz7Ea2fNiYS
UeyT6X4liLGqiXu07PAZT5X1GyUwayJpV0DLVrE/X8DN9Lyz/KeeoqJWgL5ALWsK+i+S7O7HZdxr
uC7FQm/ZGHkPZgkJoB3LoDiSAehhxR9mUZ/JYj1p1IDTJbgR+oduKPOYdgL3JNH79k2U6XLF39Og
GD0uYqpspQ+C3wh0zeAWhaYzpoFXlSoDVyrT/3/UVJTzARFoOxrH2gasCuEGaxUkNTCYP0OO93LB
4eS8ggULabt1IVf/Hxk5T1BbQ2wh+DX7j7+CQ1bYquLfCGl001sY642WTLp1X22zw6DozWaceeW1
oCS9KmQ6JlK7mmc8XKMH8g+aolymibBVfPQh4MrujithwHrZ6b5XgH+OS5xaGA9k4PreBdfNudlJ
SjsI9lHFsDxahcRsdtyOhXM4PRe3Shdk+6kELYd9jC+kt67b3vxF5dF8WNAKO6w8bqLBxMqP/ym2
uhqNrnFjOMizFNqUesUjjHBgR3Ydk1QXZ/5SIIVK5SXhQ3nBVTQoARyL6yWGnrYATP6FDkwohYkB
qgFNQuahgxSwwKTu3V3fvmgfoe04P9Nm8Z/yHQcRlHG3Mq/w/PnJK5HzBllRl+JghBiKX8ov5kfR
9iMUacbW3Hdz1Ocb0ONsZRx++l2xDj6Zbmfb21tsQipACBVOxZabWOm9gV+JZJrpw6cBW7/VRqCs
CdjT3LdlRzhqojkt78w0fA11tweLV2hSzBZuQXIxI/KtljTqaCJSqmoUsfPJ1QAUtCQ/8tih7mQn
pmvb2Ca25kQV7AkfLvt5PF/V6BbRHPZAL+R2AhPuea+lYwO6J/+3zdtwuZ5hcm0TARaNEAoCrBml
S4Q8i7ZX9G0gi24vrHQoTdu68Uyi+DXWWkVwNWx40iISVQAeeIBQm6yJfR3uqM0sBWCKxg2V+TL7
dt1yQtOCypJxFw50rheIBiZD3ORxfkwRe0NfqIE8KuEB9TG4RvPlnn0glm214uL3ZSU15sG6fkmt
/DjeIUjMwSVIqmBvttwGEeWDQrjyvFShr/rwzj9cP3yy18acgUZnmNYaFBHXEKEFRz13q+c95DSW
iQnOXN7HtLcr3W2ALlv9QlgfEuvEIOKKDLmyfl0lL2xtXXE=
`protect end_protected

