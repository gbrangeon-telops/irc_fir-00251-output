

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ya253+37kdInKtzN3pd3f0ykMvIJsSTHE2tRr5TaFzMStJPqyqbq8G0/aCj9umOixPoTbod1oPEi
NM8lNQufqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZnAl3olUb+r5fzAKtbT+P9BDg9y9NfOiCUm1R2Jcpt91ydHcXeu+pZ8D0lxHNM0CXXGhs5RFFeCB
fQNmyCQv4qniT4fHHC3wrH5hPwmAH8kqSEyGt3c0SvSsHCYTeXhpF8Chp2XvC1WNZGYymRNjehFn
t70d4j3zNeEsu5WAW84=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iKnL/TA899sfLGiFOsNtfsGv8lNgBNaSxC78jj2+skMz/TodvgTxrRQVQ/h/L38N/D5FIkKYR4II
+olODWgmPzea4VBkBMLQ7z2XenA/M8Uvin39meT5Qbx7/ksgG2EdpyOtsmAvmeXZQgf/A59DevU7
Mrm0rcVFwLpmjNvbnBOl5iGpGgx6v231GzIUzFEiOeCx1PkRai2IOZKE9lG2BMKHN7Bhsm6JH1NF
XhuV8OyupD6h/Fr6EDMMNZqriSBB1MM7btJKN6VC9jmTT/Bega2BSYjqAkfYdUTeyup0UqEM3znP
2BL1mUmUOgL1/UMAmExO5qz/A5ddH+Ai46kqhA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bwfblhQfYU7J4v01pOh0vYth2hZJ6Xlf2qmEYdxkErcnbM5+VpJUpwU8+A/bDOJB4gUPbJHCeAw+
tmj2AabGe4D0Pf/UukkjTsO8eFOUvoPbwDwH6UV1AKQFszUSN+Z4NTgaKs8pxWumW0juNgJujhCL
2ChBu6ddPnHdB5HG8uQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UTW+eKUNnZFWLDMo9paR505jK3kaKnyoN1JMPNm5SlY5iSmlguqsHIHMaqSHkHrYg25dIfFqsLa+
ygBhaN4bDhxyus3QZ9m0sw/aVS4ly/5bNlw+8ePaK1evrFFnRWDzqTt8U+H1O06G7NfpkTmeK+am
Q1esOyihSrmjwIiD3aw5SiSY1J84QcBDQl5D2DAd5uRtMADgrmEFzx9Y7yHel0j2iF6Z2vom7g5G
7K31eIbiTPvCntdYde5+aN/nl/kdiT8a+6o8fslm8ZFdkfMYbKE6CsL8CG+5F82TWbIzOMfxbILY
sXfUaKwgi3ZDGoeeudit9zXCRYxReIG0hfQ27Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64272)
`protect data_block
fFKkZPz+ogWhXnLhP79iejzHUyFddzuDtysIz7fZpuTrteXCsJ9MhWmeUYtBWFB8yck+vIfnKYUv
ypJ5PCBM4GVJgScuSgQalH61ISpvauzkGp3k8cUI16/rfQfs0rhOiqgkat3xFc6GStZSS3AAEWuB
Dh69fx6YKzNglja4B0GdgSjTqcisqQjJRysvXhhP0ksDh4vy0WjyAxIgemvfZEKcNqbGzRSwyUmv
bp8wLnTfKobr7/ICxZJnhXjmBhyftaGqv0Go+MJLWxPPW+bP0m6vBFPUrgnh3Ks+04UI6UhKajNG
rV3/uPo/wfJBYxGGVB1PjaecIZXc7QmyZeKtujF81xBT00tU/oMZaENakLIlhGx+J2xfABynfjRA
Z89iiRwpGE1ictM9ViJBw51tsmipUHJZfWMCXkf3TyFT1nov9mwhVB7/qTKTGkUvrIeq2E6B3hTZ
wPgaRdvTesdE8/dFju6jo21I3YJOy2Zs0Ung+tmALfZ58rTwOcEGjAu8mWsnt6NHNiXgkF5oOwoF
xL2w/5bEJokLVqxfsRiRFz519lqLan9CZ0C4QWD5QSRu8gFYA65KcG/dCvYPSgIH6XlUvxaZiT2h
VSWp+MHTTCNhVJIrgmce4QXj4HKFcZ37yxRqbvzkC7PVN1h1elaZX3qwdTOU9e6eBRHQQUqaxkS5
H7d1yEYU04YeEc22QTmCA29rvZiD4TWnx4WEXV89J5/+WZbwTS48xeNFy1Dg+JlD8hX6c3z540EM
RCcGnKhUNNmgKZXMnzWysTafTihxkXhcryrtgtYadP3eRYteZISVeRlsxBZRezMhyVcwyk2L77qv
z00Qz1NkovNrvqr6y5jKeutvbhbC4Z3MgCuAEq+NU3gQjiIlM24mA7CCDwb86uAIeaq1uP7+d7Hi
QTm7CkSX5nkxcKbIE7FT9Ei+gBqVoQ89f5mi8bK2E+V2Y7fT2LxxpywldAU0VDixkFMoviqDWOc2
l2EySlOyT0euIuV+tP4dodpTSUxhxbSSdHZM9dokESxmH+Olcskdtm63sx2K9y+SXY75pTsq+2LY
aZmoz0UY7zPkXGVTVUs27lXq2u/9kfStShxlZHQ7HIv62khfIk70TWC9KD/oBFRSpwwWzWb4fjUM
FzHF1vX9/N1hJxb+qh507c4MefG0k3MlNot1FPdfDutYJn1fZtfwDsQhdC2i2VIZb36rUJSszHV6
Tg1Ugs3DMcGrDoLSCLdDftpmNdIJDx/A+VrzJJF57WXqHRn776mpqMNNxKsxoeRXkxzQOpkyMb0O
57/NtVlWlHLFxCP4aq+wgOPbeTeR6b5cLP6QM/J0hn7U1Ni3SltfXYi76b5k0lpmtEjZUoHo+qRt
FNQI1Z6dqZNE8MRDrOA8OUrPBT0O3LS9rmSV7Sx2brT97Nu6uRDolV1NriKw+HddKfqynvZxD70K
AM3up3NGwHnlI0OhWUW3sMazYk8A8d4A5cu457wg7xPGQAC3jnOwEfY7YWGpZ846SgQuxW7ty3mH
PZqEWMKBKc0x+YSVLbvu/mY0YRPH9Lq1mclXGI1a5asAezzgA0QgoTpuwJqopmUkkayYVqXiN88w
ebHkmV1BnkIjhAx11swvJ/70oJxcuabxNloHC454gUwB/ml5Rm+9+nuUsBfskaR+7dHGEJQ35R1l
idSZ7IEaYi3hu8F8rDa8D4AoZzB7P0JHc7FJLdjriLGw6+RuNRUCh26Vqhorq15nPk7N1fUFggUR
vwEB8iDVpIEc2T1MYQ65cYedR+vu7FIiAwepX/lpFhZ+CDocRL8548Gln/qvkjH37OS/hBxsgIn9
yzI1REWKamrOrA4gtBNtchkSRT2/HI1H10bQf4OA8jNTjzt7TxZOg4fixZU9btbenEonpqVg+BXn
X+r79X1oJS7madYGISjXM/JlTlMCtPgT2YCGqsm7oNTwt5qPFUjXzqwh0FyEDHVYD52Em/TE6L+F
zXjYYABIToUL5FogUmuAGZKvRndSMZa1XsYbrCvw4KtpHh8IIrUiEj0+cpAaNVWHUe2Z3sNCWj9r
4l+U0urvZPlTreyYyboxofIsVy7GbmuRRmhpMVV/9S6LGtgLkZOoSKN03/m6PxbY6o58HzLC4Wox
M6rOWguXlZg4BlaAHaE66yED1nq1SDLMwTSoH3mpc0HW1DZvJbf7PkcbEL4Zzvuk5Bkk3kQLMJ+R
CCEB1JuTIHlprFSWEXmnzeWF5Y2ZNWWB0rbkRQH8dG4fK3i81mI6zh+GMsy+fXHE2rEu4Vm5iwVR
Xo5KUs3JnOcxDKpFBKFe8rlxfvSrgyTxL/nIhZL1uDJEq3PerG6BlAZGsxlJ9um/B7Stzx7wQ9J+
7VFU12rmAA4LoEyuzVL6UjE8+m6w7EoAyhhHuPn5GRuEDKNmspPPgpKVS3NqkugwcVZzRmcWvlOk
WNPiZ6Blrh8pMiQn/g2CO62W31OaBtcJhVqa+BVr1GUtuITD85xLiOjO/X6QdGBmSd007basdNrr
7nMBMU7cHbM1BNYKUKdnm0+x4+A8W8067WM5p9YZfyKx3J8iMT+4so3sgb6w4llE5FbeDEZ8Pzrs
jvR69YV02hompjskBePJ3io+DRxwU8FvbKqYKCQjZigk52UrSZcqN1gdjtpOiMkFK9BIMK55C+Gy
K9EzZEPSzE9I8WtSLx+Y+bS6tjaeTKIhMB/aTtCN38ESXaeOM4HzgB9N6cGEkzrqhJpHsMI9sROZ
u+E2ixsrw8tnrVHj2iwZgvB81AkDVs5mWDCnZe+z5w/Rb3Jbz3DLHv3eVVf02Zqzl2VAaWOOtiGE
wIhkt5v6QYL/QSBDYiKP8DTURKvldFpj4xpL7IOTNJAzbMHLenT89sviuaYADEw/xd8zN12bU5uo
DCMuvlOF3sI/35qFt5/2rIqob1QLl4t9iU7O4eA0l+6/ncECBOt07EC2fJKZQ8rLtlU0xi72HpGP
wtsN7jS9N76ZYjsGdX9aQBLczrZOi7TBGRb7LdaeULZx+aXz/kKwinxZMyR4AIKp7keKcgvqXTaA
W+au6kSu9t+VAfxfIpHDqQH83aYnFsO+7jjnnJUNV4EDYoKgrx7GguMPouLmtZIrE1sygv/i6Ttz
cfeCSRm706IVjHzKAAZC+f0Grrj9ESfwXi9hpZZ6keGm/J0QQM1osR5M+OmFjYUqWep1t6C9WDCy
hKiEQjnVe2JHeQ0NC06YX4bLEeXLRP0fHDo5R6mrCPgnoTO//B3XBqUpEvIRkakooCjC5vMZOREw
RJdACXXhsOE5WisjRQS0F1QR0zDdfWulE2/BlUmROwCLgPIqaj0F04rvHDrd20j+dPEkqwEIKUK/
ZVCJT7W2OdbM2ToyFNN0uJrsRBejCIiI8blnbnRmo0p3JANS7aD8YV/HlWq83USty+FS49AGKaqp
YVSN4LAvJ9gy01EM8uxDcSzL9od6xPk+VtppxZ62YGqrMBlzTgY9m6EMd779ON843lrCK7Syk2Te
AXrMtyhXml7c67bdMF+mwp3X8I2FvBzlHqzFt+tXcTuAyPpvK+K7HrUzUiYMUJyxbBXfwaKhw3qQ
xrZQq1C8NKJ3tOhhB6ns/mBj0Fkd1k9U+HOVydcZQMz/TeORRwNXcafYZZFRnOD5DELaXAYQ5FcC
QSUpTa6OrVAg4R3hwDQHM9uE8iDHtnzq9e2yrXsvCHUcwmNC3YE6pSp5o4JMOJ5s8CZmcjXcgSU5
MJLJ7CEovv8gFS6rvl6xhiV30qdZT9P16lylqqVKw8MmLGt5Jz2V6iyGSPVXToi5rTXmLASvQbQp
VQZ7oBU6i9rOfwZrxZjEIn78YJfDbXW3T9hnFRZCN6K6ZMbD6WHmKsiT/s+S2K5SjWlnRuIC1nhY
sGsz+eC2YZkBmf7UYdFfAa1ntXLXgLPU4aYKb9yV0+56tM9jRrE8jXB/1rOfgWVwptaFWmrz66mo
VNYz3aI3rHpS5XyGQuIdJ98gCKIH5MGRhnjcP0q9BHrf+pw7Cy6fYlqKXsL8+YKkb0dwToRwwZ5u
RTJby37G6MlvX7DAgc0H9SmUG46MIJi7BWVPQC3AdyDcDlBdsjlomyWywIRshPYiElobvwr5TOhs
rsgLFxAaUt5W3vL1nIsADTLWYcF+hltPWEWbLO5QKCJibvA5IlNqxAczU8UCKUPLmILl6DNhG1yJ
Qe1eVVdetIXRWq73kzvqC18JbEqyQPAVdwReoNYXmkCKnDXhTRzmMtnesItl4qIJoOONTwW8vGk+
k7o25H6dkC7/FziBXDU+W1z7rfdGtrzOmwRJZlNtq6r3MbOB6qDVOUK0/hEwMSdnT54sM06Lw7g4
qRb57wDT9Olyy7F+dr0E2uhvq5DkpcE+VBYAso1YvYTD6U2T5TdJKJySbSLrsgyWsdxES4WyO0Mr
VRC8KEYM52bj+cqH3e6Y1B22oK8SBxRUwwC8SRwcPGo+/6Vb6+ekkpSFWQx73lVcBaisHOBHoihw
YpmCUM+3CcMKwoNYMpflCDHfTt3eHxHYaBs2URzhz1fL16foKINpA5DXeqiVzTK/sAW+FNIHDKwf
jiUtBv9FJfwUuPLeZkehqQhwRESKrU2FcDuy4S8qjJN/IE6gqvuf4mNX8e/2+EcheQvNJAITP5xR
3TlHqPJxUBLaJujAzIi9xqUrN72YBeKWmS1UY0ICoKvKPyvoFfDu2K1wG+Qpf4cNUTectamlTcwN
u8aKnJrM3zcSg0KZG+BmJmHsrsdn1TwHYSgvjYUU4O/WmhxaMAg/tw5uaD+y0n8LjGSeSbADfVor
C6a7xWHPr7wQF+rFacD53JFTs1iJpy/RHSF6Mhj5yGQR6siSUPjY1M57Sq+BF4ruNT/P8TvlY3En
z+UNaVw47Bpo9gZFZhw+XYoGNWe7vlXl4CFb97kUQAcs/mz2U9k7eax8UXpzKQ8dURjux5VqiOuv
LguWMLIpH18PXrE6e4N0SzfSOCMgaF+DAaEzqV96Xy5/C89nNuIC2xKQzoiNu9Gagf9/4h1U9ic6
UVgfbRH8adHYvnRssehhT/bJl7cG/XFiwbloqU2wYrQur6pcYRPbEoysDH3nO9nq6tnTR8HuBpAg
00OQ3JzZ5HNn+ZWjTlbrg6cEEibz73fitgjsRzWS5SxL/2qIahC0DugFH+fu9qLr9+HcSc7vT4cr
eDcxNZrlYb5vQ7rGvwQMY3Q3T56LPUss3m6fcWfhYTD8kbMQKLtECPjaBo8wbkUVN4/xJNtQ0Mr7
eSJwXxM6zjgUkl1fiI5AI3Fq9qP1SGvdOYPwrxgxE1+9mCa/wH6a3kK7e6Dy/6NtWw6g4NpT3KMC
9gUznNRlDqZPFix68F7/cOrPS94PkbLvw+y3IXJCTUO3lxt4BaN3PnOB7S8Uha0f82Y9qaSNhSM+
N1SDATnNl7ww/L1Ji3Y8dGXq81Buh0JF3f/H0S/0b/wA042weoULTuHYQhE1SnAMBgYnUYMHpLV3
R2S9m367VGDY7lE6gAVcOH8zjVs2pfhi2RDDT0xUruVvSHNMlLQVNc9g6RMoYgI3O4qdysbbN3E8
68N/SQ1LRaIhKo4xgQrF0ixojWTYDaqqUZTM/bsRhT5K6Ji+1WdimBgLLAKmFpKcakck+M5ytGsa
wlYRPvnkAvkwEO+2FwUPR68gyLl94YRw5vVlkigVO6IGxMlwQFkW97Pw9ALH4ZdvaWfpKeMWJzFo
EAzsanBmABa4DFKO0pj79z5hWlxFz9hrBgmJ/nej9JEbtUpTCaSsLBYETGzD5nx+YOgVSse3gdQA
CLyZYU4R1U7bTk/2GYMRO3GVh+WWlnDCBVRCrgymcpJnoCwcEqBKOtivbiUTv7dandpkRc6Y05zA
vh/sfLPQaTwWAPSBVb+IZENWO8WXeeWTvssPH5mEoay1zEPFuAH8VUNU7kAXHSeiXERxBuLg4yYM
sL1RBx+ASb3/QEcDMgyGoXVa4XaQcAlCi89wBfhqR3Pq8msOHp0wByNUUa/yC1++n0K2WaJZpKNI
IKAC43B+IMMakJdia6jOiY502yAUa97SpfP9SxidaBDQNhocX7LYyscY+UaAXX6y6wOG9hz+aFl+
QLXAp1jJfxUafh+Vg/rBZJ5EMy9mTe+PdKcr8Id0vxpImPCXgW5CJtZvcWipQVVndAlGfsZQsUoJ
KQFuWIWRdRXygA/yCKN9kkV8fnoJ13CFtLTG3MkQ/xmrxNrauYCT1ocesAiGVa/onTVEbAf1i45Q
c/2lTKPcUo3xqiQMUo+x1MdXNuY5wdo10SoVQomkPGauH6q481pbKme3/L20DKnzJp2HB3bJrWg1
CNLST4yWaZ7NtZuG02GvHRIvrVyYeKRzFXsMkl6AFzkGL8aj8jLscLM+Mo73IrDmje9bQzsAHDsK
uvzvV7ug2DDM1UGDRVWdVeee81LZXimi4CaCzhQAkskE+RbvO/mUoPsSmdhg54S5Vy8B0jgMQXi7
J5wwpsCIFMxsds4y8wAhW/pZf5kjnwXDaBQ6fyk23wcG7OmtbkyfvOSWaORgQjEcMMAPrbDLcTrh
5g9wy0+jd1SnJLIHLCvKU7vErodNaZqWGNUO9NsrX/Ugt3dOhGddh9RHwa3bwJBwlWO8XFqPSo9h
azMCqQRIlbcYHupXoqa6/qFKbHisbOTb/jBRrKHOduRObmqZHaCFkdnlGsoObFzv6C8u25mv0yvt
rbMfxLnHsjM6JWXO9bB7iCloyrXPR9XySnvEAlA2SXa35ivkkJhWVOMmns8YhVaxkg2B9ReN8Qq2
1KEP355/HN+29R43YGQwI4/AZpICPVTI1MkpxWwBdeRAAg4pMmwA2EpFUtEIDxjqwJ0EHGtwoBHx
CAxXOB6RlUfuQyh2CvKP631bb9X35fTlte+ci/An9a7NgY+WPT/ywX0KOP7puc2DDU8K2+zdRKQ0
bomhLTeUGDp2v/EuJcs9SS5tcUo1u0v1VI5ei88QveT9aR8IrFCnTq6UMESfL4BuufqMfvD2nkpS
6kajZXNIWX79Mcm7uVqjG4yIAEQaI92iqD5Sn4YJWDvRg12u7CL5La+k2xb1SMCsGCG4YQf0nEb8
cZaZ+K/A7n4cKiAGHNb3cV4VRvuSwFSgLE229boE09j9K/ivqP6kP/Rx1NgHgHRhrK3VagTt+UPQ
HxH+GAkliLSECmiaurLmBiA5NFoxjPKuRG0MD0HY/5aIL3JSi0jwrQlOMb9dLGKG1x2GWCzcIe73
06DhNjTL5hC5oJH39bKA5VhBhfjn3METrn16wmZ9ABNnnby6/DXtB78nW0dxdK6cLkwx1GliBAA6
hdKEZNG+MaKCZ+uEDGBWZXpnMI74M4SCqfSNfpKvzzRPopeNvkX4X59/re/aNO6kaUezVZx0HUfl
8yZEi2be7sxj0MkDA2tfW8hiR63NULI15fVZ39wky1JvyIGXXHeje5KQ0JR8WiM5dKjjGLz0q2UJ
bP/XAX/Qim5ROqg+C94xsVpWOgdVUzgBMeEFCIgPUA9v6a7QhYWwrFjYdms1AaKb6771zWzuhMHt
2tw1m4xM9MQrnL1p5XQCnYNk+hRSB1NK+u7Rk5SHflhE9HVifr/zCVNHQYI/QB4TdEn4UifBGYKO
SmZFSDMY3NO4ZOMtH3pte2qMgV68I4O2qtq+VDoP8XHQMrc7a4IFWghg8AibvetB3eChGANwT2yZ
Q+XwCWGAi3+mDcYwWzmKO3ZKez5B8UZ5oWOK3R9D4p0kWWgRMCjWgB3x68ydvPw61eaci2bmAJRC
J8CkLYwHan2omJT6iGvXxs+vAKou2EFnXBDaoddYabuD8QX8HoqdD8mGNtS6JdzKCsMrmGMg87jb
7ZHExXi0rgZnlr5mZoQ+dKV9dXCXiMs0UW4m3VlPLku4rjqRg4xFd7LE2hkgdQGbYq17xw+VnEGd
wxh2/tY7jz60DvXMdd8kA7Gb9LBC1hc3gS7r2FIxOvtVWK2vF26H4+MoPdoPW75pYtrsLi9QTSiz
i10AuX/GtCSQ56I/mfajcyP5TaXYXIB37/3YNyJ4w0AGu5UwPDMP00WP/GaqvXnUYvMVJ6gK6F2/
q+O7Lmdo08050D0sBWQuuNSs5hai4T1ts1E+ELLup7Zv4jmW9kF348PyDbjdS/LLxmG0WjRQPqwh
PVI0e4KQqOnAmWAJivJUkD/3kBqL8YJdYKCN1jzaCbZiT8BOKtGcLQUysEu2LEXYUN+Jc5Thr3yz
ksGry1GIeshJJlCRTEkTsAUxT/NGx6FWQsS0HcYGQZ+gmNEFDCZqH0eR363ecpJKMts3Nh7C+t/Q
N12N8IxP1IEeydfuh6qIlyroIl2Z/eGS3UUMlYZnvfWxYZuDBSaPIV8Efdsj/mgvMLZTzhTnyTiR
cDMmbPORoQnp6OBHsSjjdBepFkTkjunSQPsFnRh8Asd+zPqx/N4vbfKgegwuJug3GPoWWA67ReyZ
1pD59tB6a3kSo2fGA00bJ2g6ktl8YJMalxj7TT/OcdCqGF/yofSxqFJEfATHaUqqJiVRf8KcgA6G
uC5PhcUzOt4LCqapmJ9ycPOj2/zwwqFzUUm51qgVVvmFE1vOa8TxTnq2zmaA23LZVuMv6kWWYkeh
rVSnmSzdctHYLxek6m5sf4RcyjUlVDmfrJ+pZD+RcyQn0RsM7+ginyxee4ERJ1h7TL6g3pp2HaSK
F0AvA88N2t6XkEi/OG0UWHdEqiq8fQb3SRdBvxaBsZ+AfczpyES/rBNQpJuit+2wIIIK3/Mr4Zz8
Aco9CDN7zF8eL7IdtZDYnUviwI1B+3DrpDPqVUx8XWN9sUG3Z9BxbCuQ/9p01ZZIH5DNmd2s7F3t
xBz2CBOVRBcZX2IWDN4NopfmYkSUycWUIRHuQc1EmRsvs6pNuqlB6u4SLzPR2HBJv5LHt9ZrINYo
91lPTPGXorOgMCvK7cgINcso/o37pRe+WtxaOup4hBmy+hC0cMz07xDWiOhoIeLj+U313ouK6xuS
Nt5F3TreWvnQnX2yIoO1/X7vlTGV8c0SkkdC4NFqjoBBouGHBibLPYtBM/Qg0OQI3/NVvFBN2mes
PN+XGAdAFXgWLru7BoHVzlRV5CnlzDZQa85DpPTKhBvcbX4HgYYiOi3OqJ8bodmu4gQii0ahCLfV
Wgb22Wpw72H04Yjg7oFrpSb4bAyAXrUQOK+pi3GEgSwFvf1HEkL7nBS/QRQ9/M+7TYlZMI/TTBKj
vbFR19lvn3/B58Xq+kWTEc37cyc2HaKv3eDzr+TCfffQ6CttVpfKrrDd3hocNW8BhQyoTD9TMLxf
51oWiiJGwSGj9BCs8qUsgjbIDJLptZ2JZbq+g/5V85O3FreZGZD1FNDp6mjrbOWPeeUSf9v/5DPk
plcbxnUDPPDk+gUNZjKfLGriKTRYJve/sUJdQ1tcIo9xpnNhDHrbYOuPM6zZKogc9v17O4fyrxsf
zgBuLjYtriNh49IgvR6tQXF7LMRn1e1To+71/sUj3uzVbvBSxrpUdMQVoCUbUeFXpbEdTF+Ky+5Z
srTkKHB7g7bvsu07TeK+xBCcP6JEsoRkhepu/B6L6lKJiuEDeOdwEbe45p2Y/KGVONLmGqqAFpPO
I8IFGUIZXil65HO3CAKsBFTQrNFw/SdkgQvADQSq9UU8ix2QTJrihf1w2c1+YGLj0EjgtBqlV79W
NYNGxd34kIdHEbk7T/MryMWee/w4D7HT7RaAeyOdbi3qw2pg/ZBehPpmiFltLXdxlG8OfCoSE5yl
nd+FmYNMVp1g7PRAHlmRRVUwNM5H8ZZwOPKlMhRKPtcerjFWdWrjhCaS5KKyPCyEjYsnjxiQZ5sH
+Qqhd9FGrSroxE9AtXRRClB308Etl0zScdEa4NuxVnV821QnBHHdwmtuF7wzjHs1lcL8DgbsNboF
o3/8dK/bqRao+R/EKQr6Y9yvbUyRGKBpmDgKpvNi2AKlCY4v8MqR8LH3m8SbpOJ28bYzJId8yEc3
UocC1gLOpULWcI4/vDZWC774e37bsTgVzL9XA2wmjVXH+yRws85AeOH9G+0El11TPH1OqEf8bTnP
jLKqfB7X+SDwr0PgSoBhi6MZwesiY0y7X9lXhdze+sbczd4JDU2b7MRiDVjUPnyLAAu+kwc6iROc
l5QB3SkBzgbaHnY8/KdGu7ZIpe2ZGN/oaRi9jRhGr0AeXOKLIi9rCRj9Qqx9mVltrabVTdHEIABS
LCQQw0oHg10xp+cqSgEv92tfdtluAfrjVKapLfJ4tE22/hJScpdfz8ln0Mov5F5Ccdxix9MUzjM3
dHoOsZ6mHHydAToJFQ0UFZ3305Ylw0WPZD5CLKi4GqscG1T4FU+pusYSTcq5IxXkWF3pQjc8Zmt0
eT5+nSvXxNYadCwRWQWJkiRPdi8reYumQ43RIbFG0CCWeN9LGMhl6Vw3L9VZnrbD7V+kGZf0MHaF
ili08g5XbsV3u7qIHq+/J3L0YJjwLWzOwmY8cHzmock+Tn6oH4Rg9AHcasCjtFh2gXmTBoMybHuU
mXeGTvBpsEYUPkAs2kPazF+9C6hG9iUvWxnM839HLgp7X7nC1Y2OTZnNusto0FcTtK3Mcdmymh0B
5l9MozN51Vde7kXezqIMIwlyiJ4wNAI3UDbiBXljM0hQPuzkUKeKNhCioSoXr989EKTZxHNJq91C
lnWiB+DoDjHq61BZxTSD3E9hDUnhAj4z/A6F+iDe2ULMWQty75iw20MKmWOoCTe1A9S3C6cM7V01
8ccmOSrY3jDCSUeyZzVw6BD7VohcR9ouqSScYlHZmeVFFO44vLHdp7nZIknMS5EGDxTT31mkZMEn
VR27ugovoQhdVuBOeDWTW6eLylfCPOw09Uch+Wfk0PbLWO9z8yl0MJsM+Gs62LE2kwoFJNPOqLwG
zncvgZyApqVztdvNgsN6Twk2rUAFJ50WoA83HsvC4Y6/aEidDSLZw3fK2CB0ocEHjvM7+o/dmyU0
zFr+mHIz7kuv68G1NdVMkNJ4CWAndpkaGhkBtQBQJiilTvKu2ps6mOU0xbS7gOO035Sza2VD9yhK
Emi7UUzV+8FUTAJtbZglr55WXTNzxzycKV9ODjfHR+6A7HZEAH5ZFrXbmZDRj8SKr7zDyyWkmTpP
hI6cpQRonqWgVO0zZ3akhuIKgojYNr4uf/J/7DpmV9dhW5AdLCl1ebHo9FDgY5N/fm8OlSEG6gs0
a6zq2iANA0wMCEEp4Trob/nJQYDlPzzWjGyto+3yBTn+o/fYqAPpn/XKyVfOA/DeXb2fOs+koQKg
hKUAuedgK9XDeXDWMJ1IhQHxRT3nMux3NpFWBfCtngCNWH7BqgYSN88Bj0iD8324jayESF94ZCnf
ITFRM/mo85zzdKldXR3PIYKcPEL20JskYmc/BfOReKHUCPjFA/t/ei0y/KoqntIVdUN46wxYzUFR
URkG9htDvXdPjrgpd+n8qUZcqqOJzlR1DEjxaSjor5IVWoyWey80zVMALCJhKCQ0A4efWM/t7orG
ezi/sU+qDayCFGJEr92I+H21mfb/0mwb1QY1Ftl2Et+fjPkpVhzJQM1TM/fpQqb0nwcbk6XpW5sM
UcqSGxoazkaGTDpGkvM+6bsXQQUvp1de5qSUG4iI1fTXO5FJMyU0P1auxbUd3aYm7bFbdw7TH+Wd
bDRXF8o85X0jo7J/UW608xMlJmF/ow5cIa1pqixkGEVK/FFtetDJKRuMb585YdDYzQmX6mqm9fVL
2CaQJgp4zKJ27IN37A2T3TkS5s1pcfmGw4MTBhW8PVw9vXuzSMhi3CWk0PwKmyL+zmn1tluCCW18
MBQQ/t8R8/2XD/ECQ5axIMAY1zxMfHh4eirjoCkz5/1WWmdR7lfWSmgeuv2Hrh8cMju7PGp+RzlF
CYuzJHCHbB8fNkOB5ZXWg+Uae8jey1045jRLHKrB5bAq7XrSo7LwtSWiwt1exNMY55awgaC4CaJT
7QOcTCbqYIZ917JKgZFqJbCmgzEp11OxrieKxFzhUI8Q3aYP3qd/fHX6sxwAB9t1MpSmDsoVRvRk
qhBeqqxp1lG12GFqxvihIFjinHV0XYvzVMBjHW81yqaVC51QUxg0VxOGSlzGQ5ZC5Hm7kB+U4rzi
L5e72g4FyPNYMXcAA4DNVMtHdsbsUIvCXrE89ToYpAzEDfl5c6t9ItMcThwQxirooess5VMn44PK
XaTVB+bbbXYgl/JLjMpK3cbqGfFrEuM3T3bOzn6S40ZG4sh7oDadsWRcVNDstQnugw5XKd4EDXdX
H5YXC/nn0yRI2PCFvWgsIdIS1xNcsQOGxbm/ic9/g2xRbtVd1438OOzMvr2NZzEft1rPCLaY1iSQ
+zNUsXI8tsQoLIa2S9Sui2NoP/fwNlFbGtCBPVGmyBWf8fnBPXwnAwbU3YxjaSCuggjl1ib7KgBZ
CBnoi1VekdfukZFtE4V3v/DbOFzRvf67j+JJpkvnbxionNtLWTcZVhXJo+0FQ9oJ/uBWoj5BGfdH
y2kfH/skRzRh4uS6mjrUpqPFhVbTYGXi7YGaaiN73Zk4SVoKsZ8AuE0UPdB7YrfRUesOC2X0G6+4
W/8rV9tYAjk3BGKNM2wtyGRT3C/iaV+1ERlpl0/RDXb8ZSZCt8AZmPnb0IagUTJOf7eSMZrtIwjQ
tqF/90wYQ7VpfxwyGH3hFEH7MvQFhnreDaN+HLPDqfr8tSDVRF0e5vRASbDRpbMTQNhOejEllvz0
/hee7QREEcop3rBfIruGDtvQTehqcXA/4uZXGn2u8iC+ciRNx0pVzvLXX9fyypSWZizEJC8pSVru
vgdzgI2FG6xyxvE9pAm3HKdji6X8AgzIL/qSWFpO/G0+z2xSjUEL6mycChldT1Smem1XSI8q5mjU
Bg2iF2sZZNzczTZAqzMpF/65JtuzAsHWOUN/bYLU/5ptmfiem61+0+QwhlvDx1LJA5pZ1MVZ/Chn
SSUtj/QK1gPmCBGpowimPGAJTph7d7DZ6FEFGefUlK3w0Kd+rrVaOb//Y2c3G8PqnP9aerFlMs2Y
/+BYQis9mt6HclWAdaOwmc1jkK6ne0Jj8VsBruRcGoctyV2I2TauYBMOeTZzFTZQcJVSC2KEHtqC
hU+VpRtXwqK+V4of4MROKraXbZkGGBZDQ40ULnJ5tdnCsQI9VWATaFijDc4OXvrdtvlY9Y6Kefp5
949LOtI+nqOWiHbB28Tklp+rXu1bN49oF5ocsylsFwDEmc+tEFJ57pC3wi0rN0w9yfjC9DOvvXxp
sgFCcdo+URsppKMMW6GO98FgIZ3A+3uFhqbjctIrK49RgomRyKZokmgyUq+1D5ZIBpODGcEeNLjR
ZjrZTP5RMi9mIg/A8M9Pxasusehb09Oco36LMtSAkQbG5yhT29Q0snr7aW/kS14VPaZcJ+hxsHQw
OtPIDauNUbOm1QSGEhnxnib7QOfqXHYiALeWS9CuHHaFXpWaJOWxR9xEoVm6w16Mc6z744kNWhud
zW4lJFRiqrAyclr+8y4DX+YS4SErWTZzfcetVZC/ayCEsFDcSuUBrYYc6XnSBIolwZfaYmZfsboj
PayzivU70ZQuJnzIY3dP4gW4CVfh20ibomvHB2osQsjIq0JDVHs1mmFMPGbw9+0lL/YwyLgrXQed
YiqDHr7AK/Hb2pqt+l0/dlXqRkLjjM4Me3iVS7RIKddke6irfP+Gr/9J1X+eb+cY68sK76sfEEbC
cjcD01r2kVf/aDW5SBK0yDtsLG56c6DrXt5DhAZz1zjqeCkB7GTVRuoiyLQP5FXW/1pvOoEiSbwO
WuTomlKDJDCenfiRt+Kix6hUz9kmVd4ljLkxmYfgCbuc0t8LkAkjN0Yvu6BqkAIq6Igc4ydFT38k
OnsyteRr+7AjcP5lL1hvoBlJZ/en20d9ooL0cu4rgRQXmYdY+YY3ceEMXNOaZitiiY6QvtyRvGdo
XSFb3PdsuMmLwI+BnVdXehFGOP0XcooBoWAumVY+7K4T8lNMJcVDIzioZqQ1O0E8Yc7aduEj0nuo
a9hCqbvtLk5Swpq19UO37d8U6wg8Bl5SI+2bFOxCLx0MxramE1Ovut0bUpWtNC1glJFX6mdxNDOl
U8bvzdbdOWdFp9Q1T4r/L8lE7/vYmWhXDaf+PzEsHD9oeiEOkwcbIF2NfWlsT43eerc7I7E0Yy5f
+K7870ssRcSuuoEqDmO1uOacARC9Go07AWri0gF3AsvY25RzuFcHThavMPullYNpYeD7C9maSAny
UhVWgvSGt8Sribwmv0oqfyRVZl7vzzDu7RH7j/To11LbHZY5xm0oj4xAN2gHNdIJnOrUhGQpfLny
GsD+lwM4L2AW2cK4AaKvxqk4ND4Ie7aguZtkU9D0mYYN5M4cm9aMMw1Z2Kpbk/ZsfvVkVcjFTIAT
zRryf/ZyRr0XLPt/wEpSu/9STyEE8K/L47wrIxta3M5coJgC+uFQq3cQk3OZsxpRJHJCu7YEFLU5
5eyjUBJqdOSWe79Nan6yVqSjj7rBvoaEYHOGR6kLU9AyUsQwmPr4jxgxBolGdtBGkTGcZL8TWBpj
0qiE27rlnWdPTd4NIzQMOKhe0HMjBA/Gq+kGNrKj76F49IUF10r5ctjYLpOUhUDdfpxSuKTfl0pm
VNi5UjSdEdEEWLjPgyvHsaWnrhTojtAk64WzCfaC/0SfdYXuVyv5orl31S6uaEGuN32X2SCrb029
Q4e48yBgjABrYjeuy9+AqKiCWY7+r9m2ty1A1/m4rc6UiTcTqHE8UJRdsTCe1XpO6NfThoK3O3MH
1Ftcet8bmJSEeM/U695mM0fUfp8OVrP7RTVKbbf14Dai4yR3RbX9Nyl9E0pRQLdyoRLdL4e2p9z3
141ddRiMDpelQrEVQ80ZQ+8v0XSTCx0qZ5SjXLUAHhb3AoeNda56OIL8vFBJ0l0f1TkK62WYbNk/
sb1VKHP59XgMLiQNm03orGzzGBCgtrlutuBuXs12cUx/I4yAlbxN8ZYcSGTKS6xfWIlFEPhKTShL
ekoJpcp6mtHK+rN7s75bwdWpxeV/bhSjbj3SyftQEcBvusSnWj+alg3/XYL/hxszDjes5IW565c1
mcrrJQShllbVKxmH07mw/xKKn+5FbZr+CCfXiPOxf2rPrY1UEwDOHu2iyrUzAJZSsx9r9E9Qktnq
+XrA+Pmumjgtb5xtrZo7YmHu6vpYgYjYNnoHWtuuFYmZ2w+SQoDPF+GRG1NS9tFpLhyQR70yrZeP
Pcb9uNkgVedlFns+yY/SoteU2faQJy4StogXOrXs3l3YBWJDQd7gpEPgkE5/U0TOwdP6Y5vsDaTA
R+sGyoH76ZUWF74nYnB3/Ubfl+VHQwae6Dk25CTi5Om/ml+ccbdGnKPrbq75Hyw7cTAZReibGZ1R
oCGU8dMiiCoy2Yvh0cvg49yZXQJOTC7R5rW1qQQYZC0kA80Potr9+5wz+gy0h3yJ76Tc6DnDlERO
EY8mxbeXACrCUdeRlAriwe/T980JYnrvI4+KUu7cvPj6m5Zc500NGOgDdeafVWccSM1kn00cSCa1
SiRn9y6FLfYoM0dXsugujr+vIUMGi5QdRhxBB2RjrZCM1lMEFyf9hk8cKHJhbFUf8cwEdpE9TwRs
H9J+oT2jboXKP6sYqmJ/VzpSlYoTE3Wfr7l4xkfhZwraa8cULFnIMplNOO7QLzoE5eSbxrNRWSIX
R5N6KSWo6TkIAUyAhvOYi2TP5mX07H0MxQh4B1XpG3anQo7c1Ni/GFNIkSrU2SSKqFBezmScD5UH
Yo0xo6cM8w51l+kQTQ1X+3Ctu5AICWWKnKjGdQ4BkrfTYRgmZCzgHyXzAqfncwPaLB+uRPWPg/38
XrZZNv8/JzluzU9zA1GXdlX6PKlyNtvrGAF7xcv1H+1+IuzTE5RDTpfoabtCaOJ0s8UgUdFHzsdP
OHyw1lxNE9xAVQrnjBZ/6uxFeevJFpwWX/SCLkj4du4KW5a7Iy9ozeVz4bi0+OI/qBMlhXmx7V3f
m2BRQPFv/UhfXJvlwh7Q+Jjn6NUo9tlcAp/tLS5l4bzYhjROeFWWdgYUH3W3RW/5wOjO7Jqk7OBC
UKXDJU0QINQUjBrnM8064al27Riwf+yesfU+kMKAUfYI1/RFljAeoYCxEoP6owfF/KOndObdPUwt
12RwjL6XfdQAOa2b2sjWLqowHDELx4/v0sBJHBxiE9JkmdGe66NPnsgIFSE3Ne6gKkm3cvxRADlS
FMD5RnxnZ177aV4gMP+s1BACtpQxnTk5mM4jeyxyHWdaXiR/H8iTnyIXXgzMciZ/I3KeVMscF4C0
flRGM9pz/cdcoFoysoAomTb0Er2CAaOI8F6/LO60Pmadu6awB51gU8271GtVF5q6MyC45LHmCxwe
Ru31HSvIJqTN8HJeziqegIN9OIkBMGpvcXPIOfRsp33YQVq46OB1O93PGuOh9ULISZOkq63H8ygG
m8CNY9m7c2C9rgA6/RzPh/xlpjS4BKSjFzLKoSUauU7Ph7ITWFhfLZNcR1mMF7J5Phy4Wc99V6q2
TfVoLiJYrv0nd5AqfVtcfMB/80+wZcA/W3HSJTPIiFYdi6L2VC15vZox0egRWCW6NkxiWx5Dwv3K
HgOcNpYIApLoQ+Mix+qulJt9kN9xGAUr06ZgDPja2aqn7WuaTcukDXyJoogG1LtN/dhmUfr3W4C0
xj1gQFCGFREG9XSFnq0V+N40rIUlsZnaKgeNSJLEYB7xEhoHqsi6cg6ItnvuBxxhnwAKKfEfcYX1
nH6LZreRPDxGrvdg4EYIaTHbPNsOqCT4rfJS8Jo+euJA5kjPOgEZIwpUfOyQe+bUpoPC9PsgmkXs
0RXsAGmW314PAjx8v28yA8YyOUyP2dt9/+N4Wa8EZiNzUTWNS1c5++4obFRfjFmi+kruTjPRknNF
DGUBTWcrdfbI7BTtle02OZ14Z/imr8S+zFiBwSyd0fw3KnTPqyzE8/Si+iMNsBcAVHOx4nWNq7AQ
5YkJlhZ4yJLjbouxuJjtOm/ydltPlP2ym0SNn0tPPTmhtZwZMWi8G96l8NY7e0AMP4k54CZ7OVSy
P5dGrmubrgs+jiiYfqTtgLfKzkInedXlFsxhvgmegghQuZK4CRsvjNf47WSYhB50RIQZQCKkPr9k
c6XNM0IqRvXTWtVESIRgpGYloqn9Jc5R8fY65JH8IyGJohQ/9wDKmQKyDG7xvAoMzOjwLZFk19Y+
0ZoQxXxIMWtaUOP8/saEIeOQIKZJOFFQ1E/Yh+/76wnLGqcso+vkCkv8FCnlbbU0NuJzILh13sd+
twRmyv/+S58shEU1UhmVGrubSh9yrUwUvUwLTzte+yRBLCkvLWXvASKflEHwrR5c/gOtS9CnN/fI
CSFKZ5NXrXdV1WfAuYIO8MKXx2gvo5DxkoWaCjqxdZBlBcBOfIXrj6XHSo6NPZmlnvgAz0MHgty5
ejlM5T1qWOtfuEd8T/EWE/hyP73Uc0I4p6EdItoy6CdJORXXmgsW6SXifav/scrpxx7VoJ7Y7u5I
mKnCc5uWWoD32dKJQS5axcwvchdCxWxq6ZcaD4rahsM2Id6wslZzO+iWo6yzsFUQFPSuJHm3pBjA
GDSCKga/UOWS0S3WorvlPUq/gZMzb15bZBDXLEuD993h3J+PXSUY51yME7nHZk8/No2GDMBX4QPi
OI0Awovqs2oBOOM0k8sXWilSFGETi42vRmnFRv4gjVTQ1TBcRiqGqjiM+YPBtKRMwzu5Y8YQ7wQK
n1uUkPkWVQY4VxuF/T9m66qs+ce4pB9DflVgzX7my1pmH7E4LfTkxKH8AsAHwuTaPcK+EDfKpguK
n6qFujYDajwOIARdP2hPu6wydkXx3ekjh/NJtObuzEYwWoH0rbhDWucLSN61HFD3zvYkA04lFIey
9Jj722wWwU8wfTJxg7yJxr3y1tJgnX6oM/eyvnyOtA03lCyTW+fMDdF3bJqtNq4YsAx7dayJhhFh
PGuo2zpIG1ZBnJPJBv1P+XPW0R0U2IDIo5TJ1A1JRBAo/851h3ntwAVTNH8Mu1ilgHIalWc1hg5N
ttS6ZAfTA/h+K51STTchHK1RcNVSWMQqSkCCIB9ezeIaaHFmPbUFrTkFFDOtMFVCkgPw5X/QZbak
7aeW0NYCR4JOvt0hd+gA8/eThl1a63vyLup2WWlpMzzSUhDIldaigyTS4in58WsB4JnHpa0RRbGH
yf+8AEJWaw2eK0/77R/2BYuKvBWXWEYDBtHQ5jryNWn5WzXWlvL7/DoRjmsHZmqvTcxNroyiekR6
7RGwuBcGNac4NspBUKIft3irgZD2paMqNW7xqm3x6Th0pK1xdS/+yVpn0IlHLpZ3TX1vC7KZ8YbX
KrvJP3+Kkk0iRPAVXCi9jfSWbOQq6TG8WRnAJkKE9V28OsPX1kpFDPo/MrVp8C6RERjLtbE7buBk
TPusQfaarAaBwQ6tWH04KxeqBTqFX4KG/mwmMxrrVFa30XG7up0V523KSZQ9Tnc9yVGFzfcUr0/y
EmB2TkqcDSu2cLtjxgr1YRCHj6DHmbRLJlZF69MZ+vQl1NRglL7HALV8I5/hc/+CLs+U3Ef9lTnU
nXCkEJU4eryPjbZwuD4FuPWmEB/5Z/64yoAwQCYQnrJJIIY5HeSx3Hndr0UGvJ5L4IE4I9fPTG8E
RiLgXeCJXxXR+PMwBiQQH+t4eUuy5UG6wmXBzu3P8Cwk64LAOdahe9kAhoA0ywwnzZqODnC7Nnh4
g+U+YXflmFG3eMGQeITXuy+olOVcQjuAKHs6AatS6TKfiB6m2fs9vxwUkLXsfCnwdjtChdWt1V08
QovMNxIYFSyamZAFK0oQTFDzj5WEBEnr+ySnh0U/4mNZDCwOBP0zpmhml3snkAa2GbrQQ95g7hvn
VznAgLUSl5x4LVF9mO2PdbikFQsr5dbTxl57/nl5+veMzfc2LNjnEnDkUnIpAFktE0cDGtA+5Z3l
d0owwaiD78T4BMpF6As7jNO8FLjz6h4/6EaPaJWrMrnQQ2mKdPKiBoysY/DeTToQWHpakvE4e2nD
IUAbf7xW38tj3PjVuo0LHM1Mz80WS31eAkAAr6dCN5gk8+tq56AfDiq6KjFkRR5DsvjLCM6ZQFXZ
N1PhS8nC2tYKTR5V67LXOe573G+avY5EZFGQXTKsatS5FcHXVVBzX7vwT1fitq9/8bZVh04e1AJD
hnC0IW1gulxEUlMjlpQUqhHy8dlkOhQ3BLyShnwynngxB+Rn9w6iWpR2BhWMx1jab/ptFfr3/CJg
Frl9RnAKX5xu6FMhZn+WN4n4kmMGkjjgUFUqizGZyjkNE/QzwFQxLmoh0ruoNDSqu2dVq92ubNdM
f9KXIUn0kVdyMHh9oHHzWp7eU/e4F93jmjFC1BXd4B+34v1UHSvQjR5G9vp+UYJ2hWMDW5mDcoyv
uMYo9+dFnVW8UfYvgREZ0G2m8dezAOHgaIcg0lSmu3OhR3sJhx2WaIbEFZmVLlOUPJeZjLz9KSV8
YSB0/WLtAgj3U+4yv0MF4t+2Tvl4+JIPbNOKuIqNb9EHkdt1i7Uwe5quQZkoAFke2Rh3QVO7Nd5j
awc6zisuDA+GoJnRvgV6u8O4u5s75id7h9e/za0D0kHROQ7s51a2Ftcjb61MoRAcWVzMNap+zLTr
bSl9PFSQ/NoDOc8IxfEtTyOMYx3S7WtP9wnj+xI355XCND+GZOkwG7QjBTTYXiiNq5k7f1CyzqgI
/yvVfQq8tGMgvdRi/GVZjZuPcBV0bFWxNTLj7uIZ020lz7ttSQVFzdDHR+g6PoRrT2jQUGww4fQ3
qDUVcmIRH8ICjuS4XjE86PSPV5MEMKUxU+Zl1oc//apX7+mrt4UQjLy+5q3NROySb4NW+X8I6erA
qawG0uc//Ob00TfnO3dzHBkI7OKU7yC0EImPAd/XKxiAT053g0ElJ2StqL9cPk2KHABCdHMTrjKz
WVTnfMuPeeCFOotrX6UV2zxtmT/svYVLTAtAWqRnBHdprh1ubp0wCkCpxFtaTHuKEGLotNlFNJfl
U9xIM76xg0jqhRm0vmx/NJxUcJYhmIzu3CQsPtCh/gXqDhMc1HktsUvCcjnVpvKVM8ISLmo/701X
fO4utWYatj64u010gYNqy3YH63JZ99fqZfOUiJPrS5+3IxqROzlBpZjwciO21DgFqWqCFTDfvlWP
5HFhpliCQtnuuTlvvwJKYmU2GYDZk9TOZ3OLvHMVML5s8VDAwRCHxMZ67jKdU6z0kd3V84W4hw+q
WYOsc36htcxLpzxmIciwDoXbfJyxji4n2msVjKliRZsyNOLt8eaajIGxJhAG3Gt7SRGQSMwHAOQp
mPzZw6DCaWrVYqy/rZdGYfDHp+09UOcuSjMIHLkL+ROX84xOkg5fmYzk7a3m7tvzwXAra+OThmmy
oz1kmMY5+tumaPCgV/cyhizaZ0hLQ9bu24eoGDp0sfZCXr2Sv/I/We5dqZTJJ1Q3ohbXeznCKENu
dqUnvUq1kQEvjyRu4016MhtR2qp8SHwyAk8J0cshvqwYe3AyULdgIft9scjYkPoFJ/KASOWrpIVg
PmWVo2flQbtMNkozJEowT4C100coCDj8hUw0SFwsaaHMJqNfusmxzrLmHQBvAlEo9jNwFxTFgLUm
M5L/Z/5RRJ9UGf7B6EwcH7nrUkmSC9sPsFZh2sGC1IB+ST8aeb6CTr6yQR2SN1thfsg6JKi7pBhC
sUVbV5q7OJU5iZ+pdTPk1H5rTZvORI/ZWB8GOGSlb++eL4ye7yrvP1D1X5ZWQjfbOp38m5O409ja
YYCcuMXdy0MbX7ftT1l+S95tkrgYx/yNz04xl8QveXczKhXHwX8BFBp0QDWMvYZVJAUGZX6jqM49
evY76MO1wxsDCtp00DWjaMF1ToM4/HkS0K1e7abwIBW6a3qgy3XpFKvVR4XvJYfKmis51p9yI5EM
ne01HwjhReOKB7qkbWcQx6ZxICFUkchvzDFdU7Q1rytAWSAg/gm4ABUl88XLlZ5sxVLUTV5UTpFP
5mzn3dRPXjWo/2FaH5Yh+JTQXGYe90FwQwXHr/EpwqFoW6rnlT58PzSpn5G/qoUy6oHJXql8tAqc
ljx3urUZgPpzawx0WsIswsfjrerTZ1HdIW5BnB7AIhQru1CnH7TWKyh+zSZXGuN4/HhKGqwy4ADb
QuQu+VaFgjM4aovQFCytjczClExEa0Z75dvv+vdp3/odATzaw/qAvOkyuG01p9URZehAYF1obdzN
XgAh+13tbN38sG35mntX08fFlOu7r6oyPszdN9EnhYhUJIcx2wgCX2AI7+HKH4sq1tVJzkmLkMlt
Amr46gQAzW92AawdWo1JoFwzuqQP6zILRUGL5ayBlIcYurYAW7WX0uHcgyCkNpfMmn+U+Yfhl9Ww
kmHMa/UdBWCBYADDWB2+A66Dw01UGzrFQ3biUKWR4ooW12xGOoefVgNDNIXTGOSRp04pPzwSIbuR
7mS++WnKLlb5PuxSo0N4/I5Cpj2TAc1A5ep9FmXz+cRncyIxWHPYHtM1wF1maoOss1vDGOT0djRd
RESD+nMm3ceZae4IwCz5YgX5T9dzDPOzSk0nolq0O6eiuYULAlUfBAHF4v5/tjyv7KOjWOPb0ajB
nXR/nAAQ2J21csVwSyL/VUOFCfEW8ksZ3dKpLr0+QhkHbBkw3Gz+rIeMjSUUkhhW0de1SWEBImJ5
2+6bjbZAbj2s3cDn2zPQgcZIgIGuOw8bSrKZpruWor3SUcykTIQOTEIOrY9Q44H2Z7ShLr/wVQv8
wn8eU3O3KFKPrssYY7zYtDG6E5sznG7Kfz6vC5LiW+xAqoIR4K+1YpWcWSzjs/+BnMC4PrDg8W8Y
y2elZO4Jlah3LYwC5FmrPadPBEKB6mle5wCpNMiakNxh4Z0m6ru6J+uUs9p8fnX385H9QzPJ9iyT
RA6nA8K+E3QeRSCVFKtUXoEBOGOOuhiARiU0tGfB3BtML/eoU9TK5dok/etk5PaHlz+wnczV5Wvh
GVM5m6jNoZOb11M2QdYX3JWHlJ7z2VkejAQUNz+K8NJzwW6budWjvCb+3uyzo6Qzf3ODGuOo+HlC
5VJYbbenWeXi1Gkh/BkyrZbmdyjlx7H/InSzqPXZtiOGwlGe6nZ6ELk+OH07aV019H5pHafGmfoV
L7gCt4Vw/GG2SIV3jsF3GHMeDlSGxf8cNssZ4YK9B3zrgtaMBtiNPP+eOeEsSUa9nVy+J6+lDACq
3mL9fMkW3/BpNXdoCacyNcVz8akwXQj5JFHC75sOHESQl1sLY6GffkSNSTDgawQO6dz/7Irc/Pr8
0ODDxt4JaUD+Alz88FH/ZnTSosXZZGIuM2tjLgL5xADBg4IFD5Ar7pd7s8C+Bx+MiSj9+urSp9kl
5/QexdUrkd0xBG4c+ISva/ju2jRnvV8k4TTQOurzhUmyWdrfisSLw/uhdBkz60RC6YtD/cmPZjBZ
toT88kLpgm4vYvaLdxvCeu4SLn7Q3y0RN2y8sEGo/FJJ0TBq0IfMv0XMq2ZttP2yJfh71pn2tXoN
8QABcRn8u9DEl7Tj1drmJatrZRPzNHLOkjxudBBeZG0CaMbO/V0+VPfI97BezInufDFUJJIth53+
EfuFQDCHKIZnX1ZdfbGCmKBYPus17yUeu+G5NbxN+s2COlOEVPYhJQSNfndflRFXbTP4OG56qJh0
GjmZNiT7/306HeChEzH2tjbpvaXnKJ5/PNf3qbD1gCHyke7Wc2BIefAENFAL9DS76KjI/Tuz5nJ9
U1cc0c/arALvt31x1QTFZwc1+6sLTiWSQWKstQ9ujf4EZu06XkcwSa7SuVgA3DGgdPGiJ1UjO+Gu
YSUQfH07broe/SKttGqI1osU/7Wn9J1xdl3lcxSzEwai3zW9w0k7wqgLZi+dKcXSinabiMsvwaI3
xKRVPq/Wlga+Zrpcv+/i+Kqwf+XmBZw+NYQn7jMCZp4/ZOnr6z4TWP55rgvFGzpsAIKWUMi5zBZq
qbKH2tP/82WcVLRIOg1c3tNM26SBlGvfvTbJFqSS5v+wt6JoQS9+K9R6jTeEV/fyByZLNG7ggbmD
3bctuFGhFl0Ad4YL7W6ztJVsmOR2uhU0ftKBOtLQ+9WRVJCS5q99hSXqNjguD+Q4hpEKYhuSaRhX
or1T5MJzUJYifmxS0P2a7q1RxRNAlRENaYcjevfD0UHHD01bOGUXKmBwlLPyZErmfJZz5cJfoaql
3Cy+l0oQJMP5jJeNdH7QSQotDespu5q3sF2BibEgqpVMCUPZPWDmZrxmTB5mqlY85SAFT6j6GW3C
UWyOmf41STYxvuw7YJGcXDcehPoTHGhm2wb8weWyqpZXrBb1yemm77hzsaDg/Koi5OJs8aPYpb7e
eE481/jNQoXOZAkB6LFtL3+1p0w8dxrEQvqSNQLebl26WC04uwaHdu0I5PDtvPFZ6/E2zYIbEySt
UqfGjVniDGiZv/mj+s3m2NX2td6zy73b6p0giYc49h47ffTbHemS44ZWmTe8wVen2Y5KxIWbsUhM
EB1yO0ar1Y1UdbyPdSyL/Ae47+qN5ONE4pMe02+Y6wB85r2w0sYCZSJWzFOVH/NcJpzhg9mwlo2a
FWio1HYZyk3Bui8OHazvGsixD4+JlfMG98OQGNu+Sp3uugBpNG12ysdHpTosqr7k/03XQeZQw4bU
pU2g/89VXksUB4llNDI1KBTpPWTRse5EoiL5SNqUI3PHErM9akOqreVm6Q1fMVgAk0RtCG46j/6e
YYcZDHeRykahnhMaJAyXuT3seGvJHRq2YaRLs79qbVdLe1ognBEjmsNimmR05epjZl4FAF5UrS4T
sNWpkPJ2xRVaU0l5IRzeG79I0cAsORulmQcc0FK2oHqYCJDoMgQvLI/MGlp+4m6oXv8MdelR6WkB
aHpmMjPUXc8o9Jt3f6BUIuIVM9xI9o78KqrBGYLOCk6lc0I8NSP5svKYpoLGdJPXDOoD4+RbM6JW
qBUtTeRagNQJc2XcMfoULlms4lt/Vhtm4Xn0jgXfmxlT7ab1N9VCU65GMYx6Y8CWvSlpIBxMAH+S
1fng1QBKiYbpz7i9ohMNgB3vjJceliT1NNpmhQRJIaN+1kmPqF6kucla+oNNPe0x+hu7oNcgZHG5
Gb86fz6C27TM9+MLW08rOToDmQH46WSLysi87IgHb4UQKrlCBu14ZuDp8TdV6etUj+MiVH9myys4
o7ubVKfhMDmhQjkYxsTWJe+rkgZJ8fj6IV4E5pI/JwpE4GYWlSknnWwkgrRC5Pqx0ocH35lpwYzY
43tlp4siRZjwpCix/hCY4DnM2ZKDSZyYFJnWvfVankh0H5jonwjMXaxWssszl+seKLCf4vg4YrYZ
rkADk6rEB80PEyeWQubBdrzcR8kJH/xsiZCXBpukgdJbdeX1/47Vic9+3Mg48/GGbgcrpB74RIQs
StR10b3fYh55Nv8DdgcIUZDH8K9F/DB78DXp3baFRd//eNWxT44ECFrgAG2/wq4mbu9oXGzI64pO
sE1uGbj7sBj6iF/H+n3xqN/4Dy4/ubb7ZotQXfE5FTp18rD4Eeb8OO3T7DN5GM6kq8guZgwjrV1D
g9bG/Wt2YcWV6zACYOTRSYGriK+dw+KWMMsZJBewfe+jFY3ho+ndkdgsxfdytBpaZwawtwNreAJJ
7FrdPicrtxwlZJOlxrm+jECWQRZ7rgidecp3YlrQ1Pyiw1d28EbCYhxRO06GZxvlnfCHAji4XYJa
Dq2ozFSqIdQRWQawB24Zu5VizBscNHSOgXDV2nlVkcCRR1egVRivtjebmZ7+R62/2vWVI5hZkfPn
P381cdTfx2TACxfkfHmvNffO0fd+e3Jw8+0btCJ8G1yWoLN8NjBmujI9c2OMqb9DXssoYr0diVvS
frXRkMRXtQLbLtTW84tAEZAYP6XbktD7cfeTU/rtCwOiajz4RnKOQaNY8Apg3TeKio//J1aGte6e
ZdFiEe+i9Aj3ZamJeLC8vXVYW11T5EZwoX5N4Slf5118O/Fej6jCpjVaFuxHG4b5TzYGYfvjejov
7f/ryTlDBoQ6TZSV4ys/gRVik6mTZZTQN0KtQ3OQWzO/mVIdTqPJYfznqHV906OqLerUgphrs30B
d9qQwzZQgjduuWXOX8i/vL9yvQ6U65dXVOrIdcpCXrO/iTzcFoeSpQmSTffzOtqQkT8uSI9l8T1j
e+CtMjJAPLWkwyNn0gaUEBwmTQ9tyvD2kwje5G8KjtIAjqgnsmeQq+p1U1LTPSt8zJHgCSPNe5Xd
JpNxKVrm3jKZimhHPFBubELj49R7O/SzV97cMigEVaQmKul/yT4nClC1R5I0kzwMhwTzbjOsykHb
3VbEGzzLzGdzhn0Yx/mF6OYQB8CmvwW67SruEamy5xayoLmBBeLs/mEKpcmyNchxRgJJ8BOTz/Vj
xC3BjOdZifl4TT2ZxSfkaGiCOg6INiO3dnveHG2/OeqdVS2kat7BIfICShh+U2hQd9b8mLBHhnMm
NP7+EMJxRSBvO7uWDL/03j7+nor3M8vrq/Zlzl9+vyAguV4L9PabJP67ZE6vAba2e4ta8bQT2L1L
+Fywy/TOWOK8CfX/3c34dC8wbt3lBhQQO3Q12PoBP+pX0sNCS/J6Y14e5jwmy7nxyjJKjaoQYt0P
GT1n+oaJ+zA3/hvs2HFlug4sU45Uh8UfzW/HNaJsZRv2NgbJwHSdS6ZOJuAXCDm0vh6n+lGU8Ioj
Ebq5XYFhZP7l2SQFUU/O4YQ+TwivxQr94qkHwyWiE5JAryWeKzlOzj7dQQLp6H21MTTMZtmYIW9k
cA8ictJMVUyXy2siJylho0goQQtsLRUhUdDIv9l9Zfjko6gZ28gEkBuiIKChHyJmYAUc9hxsxGEi
62ExC7Z+hEa086MLhRTehlBi6Sne9eQHtbVkln9zyjXdAQkOlPT7YXZciONRFQYDut7npCAx9Y50
aPRANHMBD/fKyRpMyOJiLyyjexU6vwYNlms6zHo0b3XfaN9SmqT+RiXDbnUknahAu6EzoWZXEJ+m
EvzenfwLZxg8iCr03q7SOLOBNiekAAOTgxUqgdVCvBJt27v0dFJEZ9QrwyaN+KwWjLoxNelIosqp
ocu3OmwA8BYfFCBcCL5R/P/GpB2MHklqkRwERJbg0wcDP92py+Wvtm5G+P6wXd2oTPJ6pl3yt2JD
RZoJhUJBwC5aNChPuzN/L9lYNXd4npYXWF6XLxtMQusvugYctzltd/h7D6kCqSjNET8pgXZCE+LB
3pBeiGFeLgfjZFN/+HlQayJgQEquhaKA0HUNNe4mKo/pWSpFOWEvcI9Vt9ctt9PT+waroOGS1MOI
F0w1eDvfZVtYTel2n/4fXANrPJFk28/TzD7TM++Vj6vONvIGOYNoT3a1Ba/P1FevdXaceZJmtTXh
ViXAQMKewYB++IC/XiZiejBkPZBE6CCAxm1K2Zb0fYHhDLExuXWeHVlxZyX700EMypAH+9+4I+sm
EHz4oPfI1X8gSTAulVoy+NL5nP8pLnKSkTV5HEWq5R3y4jAC4ipEikCqp8R+VtTGPdHYqHX8LMJr
mifnKYbGaTkepcv25Y8NPeGGYzgD4Xh5zAst95hVcJeWuuKVs5+khrIWK7oa/HX8aQgFQs5zK8ql
04Dq4d5Goq6SFKm/dpMslsBBrYrlFtzVymSQK0ex7TXXUjrjJXWfMdbGrWp+WYdTHj3YkJW58V65
w5iv8sISR2td1/4cYn0yJXQqljYG1VLCGgoPSc6TXJKkvhO+WDVwyy8lNCmQimBZabzXnwAnsNqG
SYcQGJ4oGwqumsTNhyFfHptin3pb1i9a2FV+cWadSMbWYVXkyqw9SizAIwN9ZS/9sy6cxdRd5WxD
kxuW4rSpS0tIw0LUA0Y4oZd/zu5FnaEaYgfxP/ccay5oNIHSRzbzOh/gRIUf/KcmB+CJ0SF8D3MC
5yNyudUTNV2Kyu7AzOUmwYNsSrnQpu+Nm7S+dd3RehDP5xyvpmN/3KqBSX8XF+YUXRDabcl0C238
/7Ey9iw7LyG6fpBW7q+SMm6K71vteqVmCEatXNOuTREy5JDPVXrX5PqIG7vFupavsW/mXe/M0OBa
6C1VAmDGFADdCDC/tYsniQ1h7avBhJTgqrZtbPbLH1/EiBNNvYAiCxU87J/JoIKfEWwOrPdDlk2e
V1ScC5vJMhmuk2Exl4Gxbm3AbjNy+Ti4XazQn486W+bDHLWaVJb8k+BTeElvmtYnPWl0kWDnVAlV
hmWwyfwXjG8EfpHjiCGMZm5QyeSqTPgkWD8GGCXDwlx+H9eN9Wf+0uKl0Ge5ApTyd1mI4QPkr3KR
8MZ4/WWplZX23DFnUKF0WHQUfde8lPZet77kYdJlu+OkiNKVrhuvmabCXoKKP6Dhocuq7h3b/HPo
L4lyQZ51NWaWXe1VE/GDxcEnhiQ/qXHm5j9zpEXqicbDiH7iIYc1RjUm6VQdfcw9J2/lJ/bG7pJC
fNa7liXMsc6cw1VArTtHLsviNh/ykfnaxbtT8pvcQLgS3Y5YVP93U/iFayy67opu7GGct0SYDxCB
FJdIwxeeEkDIjcgdoMubNYNa7qaJ/xVnKoYtDFZuhhkycchNTLWFLae/imV7tyxtLeISbIIUFrrP
g5cG6ReOJ0tQRTbJYHCjuehxcloBaSegn5igVAC6DNXjj5h3D66Z7H+Y77RKO7t7QdhoNby5xM8F
7SHtEBVfSCCwAB+W28wA83RI+QcBD3bFgvLvDFCvN65CNoeWB+j5ar21tTot2I1JVxRMZU8FlCwd
ON8LUG+URNi4HaD8NheBwDkQiDbnfeKK5KY+kLlH/7II6RBQ6mDcfPnxdk/N+4n1xl74JCpT12BK
XnubAkuS1tsomYJfkMmGKfw+/ZJ66AnIG4UsEqtTQbX8xU44ijM6ZdvI7H/sc/W+c2x6Wn37zft8
vv/LVkjBeXvjHTEVYk/tkEkojL5buKdLTSBuYMmDAaO5KwicAV1yidCNVk/AwLWEIhjadjAH3QhI
l4nvqFUUY8ArMUnpcmjvBmtx1usnPp05m/hcM6ttn3oA7F+ZkFPRLZRjQGMs1vORRi+Vt9X1uFR7
KXnfDQT2heZvQt7EWkXmdcsCOVkywcs4uKmHOwuVWch1EktMwcSw0jQ8n0ZZAu7J7/aMRjeq33Om
g9hkYWu7Ld6mGUvVXdtxtnrTTrhMKYfyCdTRTvVkWpRSfIpQX72jN73oHiWE5DQ4MwnK/YHiB6NG
EU/wcfHdPSQYcvzq6Dln+rqN2qUcdTUhZuY6KsJZyzSVc3Si/ycoA0eo8C44lio7VN52uxhgPa5D
iRE52oULs/Pwjl1Iq10LeDBOGDn5phBv+tekzGDKJx5KVuS4up/1ZqOUdjgOkQPtsMqGLoLtNM3c
4kw72EimrqjlFih5f1NmH7fmHF6snZHuBNt//jLbfcM13kQzMr6Hla6dPP4zBFhZIh2G3DroZ9ID
rVvI6vK+dVKPl6psV4+Wmij9SENKgRAhQFhveoQjXEQfMlmoHPMKzk4rBE2nNFqjfINl9SOMZSVP
12ieXspVsSoy0aCpYQBG3aBMjtanzchKC9uiIDi91uTav2yz2YHJ5EOUxXZSDYCgS2H2/6vVCwo3
0UClsiEY/xJMfLCTDpRjyDM4C2lF01mThJ9GwimUtYjecD4ozFN9KnTBEAOXMhLSDfwKBVGHAMYm
KnGaEUVBRF4N8gAb/7sJug45iaQWc2+hoXI7pQy7Q7UJ4J4uNFAMKTWPEjYpgRvg4ltvYHtyjAL/
S7B+u1ILJoO12OPc2kK5fFvaNzav+ISfl2nngvBJ1CC7spYJ2jagSE1+2X1STx27aHmcLVw0yLHG
MdEGOKGsARuNSDLEqsCIndhUfglZ5rPPJPawWB0/YpLRXkXsCUxkIZf9GW3ng/2LmNKZToZK23V8
XBz9ZttdiJ0hofwqcWwl+HrzK66NoNOx9IwA8mQwLHSaH/q12vdZ3bo2oWZ5xKwHVL0mcDrluS79
ui/wkUf/Ejo0JNFazIh/rymHa2W8k4ybgqlEm/l189zOFCa92yewEmI3kUeG5mmDUZIzm1SL89Io
IoHPv40XJ2+5y5balgmZZ3tRpORcJDpoUOiQboFwZFqKtSb2/fZyQQujLYrsZI4LPFgSPF+hVdKV
1o1vG9TOTSt62c8+uv03pZxCU8kpJocAN8ptM/FNuaDxUR1FRN/M/R/WPL7oAC19ufUkSpzNG3+c
wjJCmjbjBTP7NqK8ojP3/RScULJOLA6EKYe54Jn/g9XCo0qnGD5CuGSSvPsMvWaq5BEYQjcrw0xb
P4bw6ewOWDw05zEu8DKM/fgC2kze03DrF3VgrQZm8SfX2L0VWx9d9C3/gWv8U3Q9ptJ0el7YFRW0
6jzOY9fxSpQQBBEQWS7/6ZASmFu6O5EIrO0qKpGAieovmgVCxPeYld8oQdH3xTB2EiqVndtA1gPI
O/1T36BifbLamo0qx/FlBJ1l+mAHlU4N8A+TBm3ZOPt0/RqKVAuIHUf/OyOvRsLW2hI6++Q6AHXU
bIYOyWDDkGlqc3MsBN7r4gXACz45NJRe0zvlVvDauPrR5HCPcd72tTfdHirNFsgRYb8e1m0TqBAi
qivaP71HvylCZ99qDCaj1rRUMREku4oTK7Nz1SLGenRNf3JBNcllhVkt37LMr2ShBC9qxuQziUrd
NXZh5kEcExu8DKgYxqh5q6WUsxPswPgkSEDmB8XsWrZV5bXFuWAt361C6cbRWSCZ1zwGv3gNDQWu
FUx6qxqaqWTNckv5bhnrTatHUIbd+IxzFK3ZVcD8/L+7HiVua611Lnd6d8MbiWRrgUarXrIxQk4j
9MinRruLePfi673tNRkhsQ3l1B+yBOLWTLEcd4UmhgyFIAYj/hXrhfd79pATWfHrdjS+cQCqV4wg
5JkOXygGm9w44cdmSJ6oMWCYlYRFSIycldNU04QxMHKTePjU3iTDBbCnBq3q1LuvQ/ZmzfKxcprj
YYmDJaJiZcR6rHpHHJY/uWTHXB50IFY0DEZLuqTxJOJoHl6+Wv4zbMPvmdaDEGOq9M7GZCr3OqC+
szps/SdKJ1hM/L1z5uhTpxeQXIKnkPwJioAJ3CVndlpYVK3gtzLylVBNuWTdDUEuSDFy9YTwkow8
ZtUHNJSZKVb7qzcYFwdvyGC0xdNOme03Pc5UkaiEYp799JAdalvUm63ARPZcqvk00hiyGD/hMsJ6
Aeyh5c5UMAdNYFmlNzb3mu76GwR14xRwWefom10WjyMWbpt/anDVoErwly+BnahTwFLyPaiybRGY
mBy9QuurDRpVeuYb94PsWxuuuPGSbWcZScDAMxYGrTSiWtos/qs09hd+HUINTaBHsLP5aTu56pdv
f4BF08hfXgXeWUVVcQkFC6Byw78z4fXEKuyZl8wGCsgALPId2cs5dMsUcjUGl3txuyPYho3hdPXV
qazd01Pg7TTyG/VybU4dvrnvsjWp5kNWptGB8+I0mkpvMUo8qIs8iTTYBlXIAkM/ItAj2Zo4TIEU
rutBKADIv8djaNgNyCqZ33+bbNorHa+awuIybVhJYykAxXciHOdWrPJOphh5fWvev4pjm/NoqsEV
Yc5J6IeOWsRoNjeTP48KzxPqKZa46IWAAIfC0xmkMHDjiAoR/EIYYWMjTlwO7JJ9Wzij9UbCbj1j
YCNHN61QLp/kh3qZrHrfikR8Op4pTZ5rlpS7gJqYU8tx4lHW2JKVEEaf6J8POdC8+AfT+/RtoPj1
vOQaz2Ql4b4JH5QNTF6TCAe90YytBxQNFfOun5RI/rKcPsLuSAwJRnTC4/YFugshIb8oTvJ6VIfs
dnbUOc9rIx4uSCK5j5zfg1RdCM65pLqmXdeaT6kdXi6/FoGeJe9nuZuRt9wmo/XkgvoHMVvYA57I
tJ4+no/wcQT+DsqO51ca9C+WHwBpBA1fL4gK0GVY0KhkcPprWX/BX6sUmb4tLSZeU7/AizOhgjc6
4iXOa9F4ZqK8HvnxHxms1oqKw5sTJYGCrYf/TFf0Pt2TkmXP3z8JdBGcwpWo23mAnPXFTNGps4h/
A0m2F62jKJ1WFWhuuNERd5CeB2lt9+Od+jjgi6kSGilmvuMpPeBrxnA9fya2+H1Vqd6oNJjoys3i
KQ9RzLXT8Smp5tPSdpHtJ8RgIxMBUJ8+vlxvHNh0vHpRXpNZVbpvxZ959uIR885AWQRVNt083cqU
k9ikZ90D0teZaa3NYpxYWUVywYwaPR/ZOmX1/AZtljwLFmcTiNBjegiQja6Gb1CgGt5PviW+vW+r
chHTwCwhf4QolHbXOWB2wJcaJe8cOYvfYb2QC+THLAzQeQaUcIzuu0DkLk+bRZ7Lt2UU31VzXL3f
rR3gqEEfOh/MSjrUnrE163HB0BQ9Os31LNgpAaCZRzi9J3Y2hVmJqXduuen0WTNmem1zR22pD0vs
3DK4jJEOZCTlsJ6L9pSPQZQyGImr0AAO12a6Zq22/LFehZ8zxHTuetyfRhH7oXxZzDXdJ/hIAlRo
XNCiaA4k0gSGPhim95369bhveWcDGMQ33RBzo4p+daCNS3q2ICIkHz1+DMQeh6b4TKd2D6ALA01e
xH3KnkwUGriKjrGD21NN8tJ2PMyGh1vJC61cNYa8z7bFLWH4SUBlFNvdWWA6AqYdv1cI6RDQ35T5
p1nzfc7z03CK7D7HNEO5clwcwRmeH188kc1Y5q+fm37egLV3X1yLMYr0mXMljVirZ4Ne7fSA7zva
bnUL2zEr6d4VcQLOKHqNpD+nzyyx+OHbgSeGXwNFfRGXBFgnJNG85IS08QC1hsQieLPA/1Otrsn4
x/WxxDMP86M+FP72ydh+XOh1aNT/MQgGp/UZ9D/gjU/EyJDfLM8E1fuwcJlDtwaLP5xIEEMoGLnT
IoBvVVpoSEssOdoBInnG0fU9lgWH/mnfa/XPxXXBg2c1QB867bm7FmrxfcIHF1lV1JX6jIyDTLzG
QrTtvLm4P2pFjumGDyaWQS+6nsew2gHQf2BEhfi7UPDRnBYcoFpmsN7jjkPP7k5pxTXPjNltmBzn
Kq3fepCOCUDFwX7+YTIFMvZJCSZj4x3D4jBm0njY7/PaUkwmkitIvU7p5bjnyky+DRoV9TRfHIHu
FmlkELYcV68pkY47WrdXVJZsfq6RayVQsZtU9cuh91Ix9TdE3Ix320JzByKTVa7YdfJDN415UvQp
utjw5cUo40mK2qPnCcYT83QbEKlgeg3ICtqHjcWv58kITjCJlQIVuAU7bHfq3sCmkD7nA/FSgiVr
DmKU7blMpU/Lm8OS+YDSeOrv5IvJ1wWdf6az/gVRSkoSMDuE1sD6QvnDgbD3VeqqF/ZFyF5O7Jia
hScksua3o32IsW9MYH/qucVxwTC/ViJpxJPLtrreNUdez3EsoD1A9JIgv4gHeUdAQZkuE+Ki05KJ
mGnXEzQt3frXDZyOUe7C63yqxkPX+F1NLCreGK7HPcQ/HSwpPQDr1n/shlcKDbS4MepqsxwgqX0m
0DLrJiWcKKNYheIeV/2DZp4e9arzGl999aLu0idgIbJteuDCaaKPvRlNIPv8tltsYJk3YxL5Cerk
2GaUH9FD4oWuhyoCP2Cs3gvdBfza3hylJsI5r1gxLJXjOBlXKR/ULpK+/AyTYajq5zkzGfzQbUlq
PC5LjvV3xzoJpTjehi/nc2EtDM568VyGCNyNbeFTo6XfsGsrGkICsjxi5jww71t+GnsXfdfsy05+
Be24Ir5KLuPHsy12nBScFDqk1ZS0iOs8wONaJkqh8jp8JrZLGN9YXarUMVlLQhhIcuRVbj9PaNoK
mhZLPtZyLarsPtXORscJfSlBYpiawfw/8T2eneLk/uEwHWA5X6tx+nPVDap65lMPvbzIFJDXPEiS
DUhRO7TE3co4thjpMBR+koACJoKyTCVCAlvUZDaQIS7NEzeu6NPHgQ4kGaJ595cNJfAF3u38ndvC
YazDm8phhhh/GjxJzNKcEJOOyxEDvBIFlv1+8KFj5+QMqhtEmA9Ruxrmqr2jejkU1FwEi5bYUBpm
bev4HYDFm+Z6mKR9bFLUw1zTeN2GypZDNVCYd3aHrLs0PzM7esqr9ZoR/O/obzS4EE7/wVV7/MMe
s+ckRTx9VA7im4k5lh1LDvY0rPir0oYU3kfvmd5RoQRth7E8qhbj+WzGPXieATY4lwHbk3nZrvxz
Sl1OyNfoK9MwuyNW+fYhtvYz31kUbUJbfx9yoTAGebHHWIGSIvO9f9paoLOj993q+/F1mhFys+Fe
yEzmOi7IfEFAVLXlVISRK4K0RlF/HjiSkg1leXMu3H0jgRhdDSjdFu2qTyIiSI8HRrtZTVwpCTnC
qO+SFuqAtJOIw2OFq8hAGMNRO1c9b0zVcSffsZ4ZjfW39Hg8CGx4pZaDI7tDGvNxCIpMFV1T8iWp
th1RaMUAoR/6p/uOT9oyNAxs62j1LBko2YZ3mvBjXiNNoj2KR2l0NLuIIRIA7jy2AdTOZ/CvBHLk
uzfSs2G5MOnO2x4mrRUmK0nt335x2il0X25Y99jULdocqqLgB5u1EV/K0+91ApAW41ITEW5ISxkz
/P88N8Ua3fC0V/Ddh7Gs0P47UoqEvO0kOc3cTgQESdx0NP4wMGuFx7ZBk+ZjLMl1Ek+KKeWUkW5S
nIhVCzO2zs1XVFfMj4na1W01rUYX4TzPS9k1IclZTRsdi0cJjxg5qoXYISJxeISQxjHbwbsUb54S
563+PAK2ZEiNFQVY/FF96FRNOpQBQ+kozVlLigqGs5SNKTjJss9igcrJvLD1kvz45bPYNLIE5C1K
PZIcyz+rfdrwpZQp0ajdTauJKFDjB99U8ycCGH0ccTgGSg6uuonydP4gxiVF3as55QOgCjaonLXv
mVy8Du4hl4m9xgGxYCjPLAA2WUS2+TixGsAETUFiepm881QJme7bhD01NOU8dC0UafT3b+zH8z+i
hQjkPMlp38jrdnIjWOWWRMFTMrrgvlnhn/NLid2lXDSYafdjp1gX5Ai+5fBEa2gHsYeSWsskOSFj
M184RwQmtsHSK+MhWRP2n7yn51il5Yo7GuMj9N23jJDL9lVM21dLvcmdvYvpZ+wkTIap0eu3k+wU
R46c3BSToWpvUu5NxYh/0RoVXRkNmImvlesR+a1mYVDEAGrBGNqDQ4IzJap6er6rVVY2ZwiK3+yR
gr5xyHvBA9k9wsX6Ech3wDsUI/VEEyf0AozlcO7xllP+CrLaCjDAj7Orx4XiPHDz7KcHEqVNbHut
VEngUtnSMT/yIHmUJUxNfJ2A+Gs8qZXIKnZLv9LWyW+gJeaZDRZ3WZ+4K4EmatBvUgVQWwhFFsNW
/qK/pFl8QydZTSdegVNnxToAjK3ZggzXAQx6fLIYF3ylyab4ylgcAXpBx49uuMT8ZorzlQnuuAey
nvRoIRZtlAS/0pD3YwJGZPOd/Gmdn2MCvK0glXBfi20rX/Ryn4C7mMkpV+nst5R2kdDUz/yYnIl5
uBbja/sj1PYYcAVFjKk4nlsLBXpujoVCe3W+RisHWJhBxY6GrVWyQPU2MlsS2F2RRqJI0NvdcgTg
mhBkypey1tXOh3AknFiWF70ePext0OckX/czSARenkhnYCaFdZa4y56lqzmFg8IVY3K9jHBDHDam
k8H/kqumaoFvzV9HvWsnNwFHj/mNc4DKiEal/HPzrA433fv73+C8InAx6SV8dJCNCxvw2ryfbfM0
q1ft9ogaqvlOdOt0gQ+mxHc8P2VqWHcAh9QAMXWUFcKb8Vm182bjNBb41G9EsQ7IvjumX9jxoUUf
vx7mRi87unX0MV6ZqoufWoO5FjaYD9uD/JCY4Q6MfR6Cs/eZNl6wn4iQLWrNW+oe/bjtytDtYQ9i
o4y8TmaFORbTY44GUc4ylD7sTAT/gkmCOF/cAfSJAFtRDxEN7bGG4Dh7uUYNdcL08PvzbYSKKWLX
Y6vvqZfgJ6IJ97YoLtdGco+YnoTw+gN2bymjHz21DbHVYExpK5QUdVJBvZNv+9Q3Fe+jeO3qzbi6
8ABFPK9T+Ud6LE4GhgpOYudgB/7GPk+oBul3P6q5UZc1PgP9IGYav5NmytMW6WkNuaWegYfy6wlK
M5HmqnQzUTHrzhB6cXMh21jXwP/yHQcSUFB6vWc7SwZYy0DsOVeKgdjCPo7V4+XzSzaA3emvV7C/
k/Q7Qlyo6VWWfyyksM6OFCYnBZYjsFVRCNIqmzZPdNlyR29yg2Q9/1nt65fZQBqGeJDbC0F6s/1P
kwMWxzqT9E2SbmHVBm2f1fpimN3Ctn1ji6eAEsw3QDgamwCAg7hlEUGIjzKGkyrbmE8M+WPYSpJh
qx8YrTQWpBry798DFzukGcv0y7QfO7kFYG3dUGh38tD/tqPvJ4Q3f/SJ36XMgX92DBwXYDECayri
hLgIC+g6Xd0i/uSYet530lvI3AGI+aDmM/fmEzIngBrRew9UZNMwu3B13xnsb6Clw8QFh3BTOOsJ
F6Q47Zy/W2RrnZ+echS8YgK2heLUyrsxST2YPqT/gkecyy7W6AV0N5Iw+AK19XzQqL4eWmp8hddK
4TiN9TiM880vw208REr9VDF4Uyf3GdlKJ76jHkhyJyfSB8hWu6Um+jcW+9cjTIn8NDdv6XfRBayd
8eZu5vIF9v2cz6SxFB5Pz7RAKTWdYd2pM/xlf+GS/q+ulKZz4A31o9KeF9Bf0TFQAoJBawpfMGhp
Xzi+EwYgDp4tzBBjIIuX/YPoJ2/fTLv7TD+vQcIQohuGfMsY4JV3Bsi//0GBpXuzKJb3Q4kvIdp0
8t7hG2WNr0koWRpu75sQMTSFG6YxOIfW1ZsyIiZ1W8sdGzmEGYlfu+gbQoRm9QefD1goo43998us
gcw8GdVtq8KbfoJi2SWZYe4bKeECJx0zV9kvdayJvWN5Rvh86YxxVGHX1B7MGrk1hv1gqRs0okR9
lsILzLUDhzGST/+64WdQ09fvGvj/215hVdX8vuUh+VWI2eHV2yeEeHz8T7sROzPbOtZff/OywDzh
cpJqeYky7oH/0UHzX8O7vqQU9EVlekjMl8CKOFm+EgfOpaUFw6SVBPvSbQf3OFFkjD4orP5QUGWk
ll6RTV5dgCM5jzolKzIcYank8gUqFVn33t6v51DJaGbTQdVfvP8QjeCYKZ9NJi+mAG0UivrA+Q0t
u3Z7+o85e/e8yqXutKiuI4pknJ/1+tJyvD1yeYsrJ+YXLMargMRwY5e5vlErNS+/NVFP/sUMI2mm
rp9t6uMc6uXrOOQ4Z1Ww7ukvpEa0mwO9Iw5KzDPSsMJaJwp26fHVaSa1A40ttVczc3mAS/1snV+y
qOK3DadmODFKlBRuPwK12L2UXS8y48UCAkhNJ0fQ74e+duBxUv1KhZV7HGZUC+a6Xq43X7ItDChd
83jDwLgXBsPkGHK6IquKH9Fab5G4vO+s72Im5cXXucMFD00GYYeWrUFPlhd6TmGzAxcycLUcklMv
8FuJge/4deRqVazO5T/hzHmlUL2syTde7H4s4Np2UwKw1jQVilcokJYbBA9ah2eNk7IMyy+OSd+y
m0vqPrH3cdMyd6jM+hnmMj7gE7EkPDzkxSa1k9yFuOmIsTy1W+xBQBuHqhhYAbga4FvT017wP/Mq
FWgz5pN3B95hZQlu3Tu9SUD0IVW+TjHz/jL7jMYff85A6qddWguNYiKLV4h4CBwL6F8Avebkup7t
5Kqn3eDntIH4AdUW2MrcjatcUk1NZI+Jg1sMqG8nDuGJpfNgceEymb11ZYliDwIhxseoXjJKEm6q
6pvvuGXKIWJgqiV+DlFook7cFB8EQ5lFo0OKBE2cWwCWLg+7uYHjs0P5LHYGNHnasODC4in5gT9Q
xA3Pm1gmSspTOVBA4xwJFJBzhpS+U7EZmK3JAnTqwR+0Fm7qmg8ZjnInooXj5xNFfzplj+CfTA6b
b4IeNypNEiscXFBYPE4I2SgGapDec3SM8OkEkqfvg73teOrTIj+11coZlo4FpQghx1lQaR7MTwCa
9PF8yeFS8JoruZk9Kft2YD3Mx+UDbyBLZ8LgpD6MLyN0LsSZUVX+32ViS0usFy4YGm+xjEJs6R6b
fAxvUJrueXA3qUbQumP58mwvDXxiB/qIA88uaLn7G7pduAtGkucUirBk9L9nl09S8v2L9xMT8Scu
GzUfRmwSIjdC0tw5domRGdufYTZy7B7XaA6Ww4BIxBJsBRx4fwg3S4MxlEi8Z412zdZumPSet2Vk
e0ui2bcmoAKwZnEEA0voDHk4KeCpMKnTYWOwelkKgBpAK6RAeu7Iq8Mh2LumvF1zjmNhb0VWPrz/
5nKy+tl69naz5qjWway2oH6/wTkAHTznuy2IXYMUz0jKIS+4xJnbeqCwhFOCQhzPJi+yaD+q8c4W
V7fFj605JdF+3RGcuHd6egzYUv+JeQcXggEpMqVnKDAwOmKQencGgDeWk6U3OA2EhraQrCSCdopJ
kPWgjT/1/G/TLfhKOaLHLv7PjZky0vjBt37gcrMOvaU3I+nKEl5lmsNyr9Q0X528wYVYSFHg2Tao
g/AJaFpdteRi3VlZLjcq40cEuPz5Sr6IFQf/EqpXmWLyO8bIi4UD0TuL2Abuf0jKf8IPpZJ8pgJU
oY6J7v8e6qDjXVfBN9eHLQTCpCWfCjQiNeSS10PVIw5TTO+Po5VZ48LweYsyUJFvluXdWqV0ixWc
2glCoEULygNzXVo7OojOeIK4kO1gA5C0/pq28tpq9M1Aos5+wLRR+bQWeJlAigJ86WZcj+Pnu1t1
GT8fpKmjZiUIqpxBGs3nxrmaHcSTLY0MgyowmzNQKcQWeV5Ze6sDTei7Tz9ffkgo9x1ZG4d3D6wH
BdFDciW+1D79pZzqMp01tiE8dBwRkkvDMoRfFnn3lBVbwluduxmURiMHD0WO3VtgZ+lnT1f2t1qs
V2bXc1kKhfSUHgVQQPjsdrhLHCQ+2bauX/77zxRsdAqL5jP6XmMeVO6hmetRlUVaxNIhec5GIRLP
0S7XT04XOFBg4Mqt7w1q66wOEgHAE4VD00yjC7TCaB/mmi/g0sX8Or8xBTMSMzYCV05z+/o+yIM2
0ti4wwzhFhROyS3usgZIYQJ5KxPr+TCcrNQ6eaTw+CrYNPk2Sm1SXD9yGZgM2LrXgBJ8diycWtCy
aKSxk1G46sxF9n2HXXxnBjO95KamEsZi4tA5vwZ16TrscO5YBOYmagtB8Wl0m2+77tbWsTojNErw
iS0VlZ8c4dqjX2ZkBRZovv31DRjbwk8Y1JJKiDG6YTWmzfFmsGUISgpev7z0TBlpQLjvmWb86Tzy
YaO7X1yR88QHtagfzkEVB+Fiokr4icRdV2KTucsjubrl0Wt7VpM5hGQ8SBV4Ck34ztDlG0vCXhcx
Qdjpl34YV/gjymuwMHI2YCsuoQkU0UsyI4+1ZroxuM1zfEyBmB7WJ/quKJfSvoiCkrCXgyegg8ps
jytamkcpd06411G2PfmhF8GAz+568UX2PmIwLjUs2wsy0r35ZK+dXEuNAnOL5Ita6TYGDNLLTEw2
KdfK70gsShfKUWm+7NUvdSzgN2uqwkUTMZkm/BtXYyNfrjK2V++O7Mphth8uiw7d3gEH0tkLM/Dr
k9T5+Mu5gUzcbOSP+iS8RcljekIjx2nSMosJZbq81MitOwe5iSJgVKvrihn3wGRkfQ8PA919lD3g
m7kttX3z/DoqLMwrsTcupWq2S45sFhCo+5pmKah9LNzMb9Io5tszWJ+CC6w7JlusIrGR3VCgn6eh
kM/IXGL8gvQHw9hZVNCEgbWRyHFokq7GV2/1hAcEjQCWSxmGQnNUJpNg/euYkTnqIAqOj4b7fyyx
m75CYcLBHBgdA/bJjLaF+lpRhPeYEUIlV+k5XqMH6N7yzS4QS7dwt9JEWdDgvxI71AvbHWbmDuPP
c2mUOsTFILjsQzts5r6qc+wyt7HWKKphbF/mgUtFXHZqQWDX5LU7GZpeiNOfIXREsjRODkuNCicX
R4IKzN+IX6/PN4dv8kPLnqb8J4XlQ3nGsx5qXBKlvicn9n2sEHuJ6AKipLqqQ8FVVZdu21E2B2uy
q48ZuVxfzJyBcZAzlYT26hY9mTs3LjXhJQtS5G9hOgcd6RVIfZUjs5p9RTx+Jj4UWGs/Ar6t25Iz
vpUTl8RvVdGtccMjeCngjO8D4S1gOabWLf02VENKkC6rlV+VNEx40VEsPNIFXLToj7i1kW/kWB34
t1KYXMsRU2fIBI8fgZ8xrbHhsIUMXx0fJ9dx9fBOF0H60AdcH5GgT9ry0ZYHp7UJvXtxxyqly08w
lFB0cdY9lryvDQ9tRlN1O0mKJT0RE++jPB6Rh0l5ffELYEvcnzrCUbPVHjiYWsZKQiL9WrklxMRy
us9unQY6w7AWdLTp9hSOw9JKBjll1GbyXXHET+5oJ/70QDtkvpyY7WdR4lizguSbY6KKG7RBFg1T
hXFCfKCNnnf74fVbSFBoSJKrCutembOZFHstFoO6RU1sb3z8xne3ijjyggJgaSpQBpzcc38Sepq2
+QlraaQ1DoAzVvEutexiu0thh1pIqyILu3IrT8cNq2VJy2j3estMZB91br9Cz9OSqjOib+pLvbYM
n5cK4tM1PjVNkU7An2YE+ApPRcyww7J62SYutxam+SGZdUJS4DyNbkGl/dilJbgRvzPWH8VafSQR
reu6Xpi3yHokeU1pPRrhdDIG6bQm4u/wWiLaBb2ub2mOZhPMlF+gQrnj6nP7tC6Am1bn6fQfSH/o
yD/v7uguAyRmESJL8CxQB9bQDBHl84avO4fVbdDLJDsY+gxGIuQCqAZvrEKoam7Or3XembLSPd0J
1Yu3WdAMy8KjtfPLKONwBmJ+p0cS2xkUU+pQZpu2iyYlrkNDfSeWKtGrQqUheKEWj8Zfssxphw76
+u5C3YAnnnSvkUrAwWbrEMX42i/ZujCKa+50XhjiNHiFaK3mKqcxM8nfiTV3dg5I2AQBTGG87FK1
DwRXFHtSooLIu8B2WEshXHRXSJTJePtfHcOccL1p543LV3fejEAFEEms0FCYCWAHQuTvtXUeIHCf
K2kGvi0SmsqaD0dSoVQu7VjBFmo2h89Nm9DzukwqLi/HY0NodyCVemgOvQ2fUEK1mWGP0kCqDv29
xWsqYLzosNaPpTkneaDuc5yKM8VxvcFd8faFW5Fnx39XNXkYyPU7TZ2lGMW1hzQIiQm9rLwqVe3w
UbxFeZzQ6gOxzeGm0ObbGLHuq+GUQsShnVtHIp5kq22GYU+WmQPPAbG/55jcA5HpxfUAR9zw5G9u
4ZMrsE5Sy9129JePK2herL8kI92uNofmtp5EgHHeQx2rO5G2MVVfQtx/J99AfHyZeGJU9ekHGONW
xbt/hea9w5YwYyCzpZ4DBuv9zTPIIDeWq1JaerwVGyCsMuoOUXAPAe13OOsBLLjOHUkAowWuPX5c
UrPtyxxsT/1ZtS2IL1b2CRfTW6BdkSyyPR7bQOtkJA8GX/VnAugipZZqQ8b1fDRCVgNFGR3LPFpw
oQaroOomW+nVE6XGOaIXFYAVXmsFxzIhC9k2d2XzIN6nxvUFPki99bjRc10bRtbttPW00+ygz39a
TduhUBwInrTa947L+2kBaoGO4s4gODUB2R83uvcN/u/SEOws46fxeiEzIT9miWPbE8eT3Sm2pbK2
RNuypLcPNMLJq3sH2qEnByaJ6iQf13EvhjWm8CEv9614ZNXrp+Xs1HUOgwIM92PZiMt/FL6u52iP
Y7PqJ06u4SSINQYC3lM1J00DoxoGI/Nebx1riCbhgM9bIzezj+Z1L1PYlLD6WmpD39LtTbbdPMBL
eEMu41QuF8ZjXW20bFw+Vkuzr+uREsJXrsf9IZEbvGDEN/cB3Jq28QQ9hryaxdZSamuWRV+j2oSM
qDBvJmYdxr1TJYS4/SrQJVqZIdPHYKrGuPVqRkOhv6+NxiILdykyVozBKxZpgKzZaMG5KHXZ3mT2
Tvp16rdDS9b5zR3ojXzv0tCv1ma4pHcs88Bc5R/vjWV0Lpv7X5zdDiCXorzFLbEWo0bkkXOR7pXn
GWPk61bv+WtPnZi9AyoQIjNwBrvWXzK0Sdu5PAvo6Yq4VvIL4v6et2WWN7wVSCJdv32v3GrsVi8r
4qbvxwUo6lhTCFJYFYDDEKKYNqI1mn5xqvSvGO/CToikhELRAHYiY3x2EPCK48uG2/b75QseZy1W
VpTjN6rWD1LibqprDC7oNh40QP5deQkkFCCLudXdZ+7OaWPrTK5U+SrNDzT2bKlS8TyJNx195Tep
i0pIso7/6IhgOjSMEmSrA5w7vkrnVOtHbEYvqPKYS+4DihywJ8pk2JiS0SfoGegMP6XE/H3FyLDC
IJwTUdQ8GIkMZzQTcjk7m+nWPEd4jEznWClPC9U62X88Dni+ALkW9D7P4p794cjG/sVSvNlcV1O2
NxNc2/V19bVxyd2EdBdhYkWvQs9uspJthIunCC5fein0sVXXn/AXf1JTMt2Y76Uq9hqSYstvYlX5
7tb+mteqM3b3H2rzAtiRetdWJKTOXtQTTItSfV6aNszJMN96xUE0+HL72y20hGbO6X2yPcUteYJ/
pemIOwx+NMiPywaTETIGuoQT0+C8hv+x0NvrQbg9gCoJK4P5Z/1p+Zo5hKZHWLUlMYufSwCuXlJP
44nYFHYrqo7OQz4J0dxsqXayYKu9lknwOmtnrTBWxwjNqTVCkN/6yaAZQgFZKsjAgZakUBrhL3Dv
MyUHIjf4J3KRsZ700DIemqQpBhFSee1sEqtoEb8Xxzdu5a/dRX+adMzi0wElYYCbLWOtJNLgPBQU
vIXaNLjxwg/fKI26F64BcwbItBcvYRrvqoDhGtlXYU8EY4v+r4W6qFoC6OogFxz4Du+aOyOhNBX6
96Kc2JUOHHZ413TyJG4NJlSTsceDuPcNS4iT/wdvS59Jdxeg1kmrNLp7hB9WmPg3ISIlOqY13B4w
aeTAC8HYIo7oJEq9iqAptVoQkaYj/5/AQDZLOtlyVBWRGoJNyqi7R1veC1DoXYb0h8qylGUmSE4C
ws0PWYHvoENkIshNox3EkdeFlgQmpCloVu5/mIVpAhrEdf/K92duuqxzC2L0JXZm1YcrzE5bMzS8
J1if6ZvQkSCSFUxSP3AxqVVEQ8vey76BRZ/+jrOf/L9DfxH70fAQ4DgnsYXfj4AMS+VZayCmex49
VwhwjJA/KeweykDvtIBR9rtNP+1lcDHFo11vlGU+mFyqmk+YIgvnna1jf+CM27AbH1eBEwL0NVpC
rGJs1/YkelTydm1+wu6vOoq3efJYG0DFFYJx3i7Uek3+OcoeF5cF8ReYwObGdgEi209zJnJZxEW/
eg6OcKlpsSTw+0U8rP/z3XcjP5bibS52io3j65Cm60qhvUT6RMZBivGV77ygeCWCizRtV5iSQTAi
GxwqwOATxjX1fpHLxA9vlf9++6pYgsZIzjf+LIoC7bnBGEa2RV3Wz2bva9Lukur+S+ICdAieGqIQ
o9s+qKKdT9d/ztiaUu0i38rKNhxYt1nbVEgrYVln0GS2d6CpyWjxg7CM0JKOd2MXKeN5aFfipYz3
tUpbRgsyO7VhM++sVL7ANJ/Mb8iTRQ4Cf/ZjZSi3Zo508JhdLRom0oyUOh+0wuiG3IimXOxFbngl
5iIuK//oAUFT3280h3WOTo3ynH1uS2JhIyOW5HpPAvlVhZr0xel72yP6ny/md9W2RaLJt0acrDQF
h30O4DsCTnbW4vF3Dy1EkQug9SWIQNWmvF+3lQFBf+j0yTkOBoOKHoY0z/VSX109JIwhJopUXusR
T8fO7ahaUcb7t7AGcH0D6Ax0C5+uSaNKr1f++4tDw9nvcng5b5TfYB5lERU0n91niy1J4lndogcx
GuE5bA5dS5X1k0cnk1xhIKn6Z8d1cX4sEwkX2GRTemxX1Y9QEtHtzKZTBar4fKrAfnsPJjKKAI1g
Ngx9Z6tEhowGPKSXug4fskef810kJb3VIBkRq1J4PpgvGG+D/VV5OMYMkC/iIYWSuBe8c3c8MIiF
8EEZ+1PON52vOGB/Sc65IXwGyz1eBTuwE84whBwYuiUrZuYMD8dJk4T4QU4v0zX63ByigCO+sKbv
+Qs6GbMDwGYhjM5aOR/wFX0ishMhqcWhu4VzEFd1ZmbvT93JWo3WrjrnaJQDg+MABBGQ7MTduwv/
PvUqdzJuSPVfzvEWdQs7rv9xIJ7yOT07KtVg8i+iH1+FBxVeVcQ43t0ZSfGDg5B9G6baKGKPUE8C
hHSzxTVaG21OA4z7lAURKgiwWEpGzrhsLRWNyTFesc71pvNtjTGPN1rS7bJw82T3oJxdmyC73gfK
YH9x6azqCLVyDwSEmfqbeEJTo3gV8ZrhZesUBbBq9q483Qbxfma3PGp2X8larGESQeGH0Ka2Dics
id0m11I8+XcCtPFrD+ub7nOGafqoRUR8pDZd5COPBACXDyYH0//vobrRWjVBtPkPM3kUasFbfc/N
o49cKrk7MiLvrV44eKR75SuxR5RDEwCY3M6CshPGdIvDm8yRhU+RSHUDeoFuTMSLe/yZxkdLpeVG
VrWPkD2ma+TvKD7MqTfWPvI8U2rUNuX8W3ITAxKxuzpNEmr/+5OnXvHKBk1mUMlAc3MqTF0GIIS7
cQOdHfbqQ0tTY0bzYA4FdVoIg66xJmKqMrKFZhMV8zYYyxx79oRijbL3+eGk2aOMsUKbKQnzIQi/
u2cTiCa42V9SPCCDEzDgh6PkgBbc+0G4DOdFuhMRd/bKd787V8ZJW6Ln4goy0AEziyxfVDjfNp8w
47Gvn0BQTMujfd8OCzuMNxECeXbo7VAXTYxxEoAAcDNQo2OvlIPwCDC0EqfXVn/flfd2Zq+7JGwq
xigoyZpPi/BqdGvqmwJ6QGjoqxjPAY1eD+/pVH5j0W8oBTJpf3QdvhGXEwdl7kdDi0v7S2R190Kh
9xvgIaST2d8be6bau3gr/nTJecjuTv8Iuv9GqOv72J6jnOoi3qfIqdmlZ5pAi/W4+GgtXVBdd9N1
FpBPplbDfRsrNFPE81/+C6fjqTMP3qC30z0e5SV/hjgbpXR2lqE50ABNIfLxQc2IZpinr/oXwIBB
qVdMHJn0ZhyCVOsDW8ZDalobQs2YLoKSFCNQ/RXeMWXHoTbLExrGJ4DqQLk3R1L4zvMAW8+1apGE
lfUTsTMLT/dBw8RLGHGB2XMOY0M8mDUG4CYwRlk2P03hc9iWJMUrbNgksQcEbpIyi51fieovlCn0
HjaDSy9TLhG3TwUUOqyyiLOlrCYRPERc2haLk6WTGh+XJMj6EnEFWCGG70WvIORMSutEeBUXnAOo
ZoRMd+tBt3KcPa6xzKaf9zXFCoIxUqY+MeiTBMr6w5x0PqiQ7snKiWthlwPSlEOM43yb7fm8154q
qLLWNnwGlYjSb9AiFcNPNYz7GWOQer5aF5dL9WsuazQt/h00zPTGiJulZmmX0z3i0az9/7T0y1KN
1KinFmM2pFE8iUJ3NSA7KIbPkfOqjs0uppSstWe/oVzgKbovmuz1Q9rnp3ryHsw8FXz/TCt9yool
rgzHE24eWOSzSF0Qj+ZmiHLXuf82pI3NK4dLJP5tvs+0AYPolo65qn1NBoO/csdeDMZcO+dRTXeu
mek6hO04t4NTrvVH71sQogl5j9mYY82eIhb5ynKRUyBRkzp+lNGASujSiO1SromVhN5Iut67VMod
lNKXyR1RlPo8iPs+1CCNF8qCnYmjGVHLBShypRh/otZ6RKxVVvt+QPjbIg6W4Ej5fE/Rypj78j2K
dkueFsfFZ6QmYf3LBxAoIkF+voKV/1u64dqbdOBxycLCJivusIygexBXMHFgaDKKdLYAtQyCWnaK
Pac6c6soiy8KxB03LWZQkimPgXyDLoaeN7ZAdVQMh5qWPlIChbKRUeiVKg4tIuBYojE/QG0IhND8
Qzfo1EbDKeX8XFs99+7Cui7vwFcJKKxEtFgaZTWEtsrTdPJVUUWJ1q1VTJZeWvWjGJABYsB0s2+b
89llKcMhk5nc+8yvmoR1fIjPrn2LNNj4sEPMdRwlT4vIs5wiLKaKpOawJLHHY42JyTUXELaxKm6H
z5HfN1NMSgSsrOGVK0Sky7rVoVwKESQQJjUYAjrcKz5NHlq1dFijP2gStL8v0KVbpqe4qCmRvxV+
S+bdjKbytF/zPLuNlksu7y8flcUYrK4bJHbhkNPaiqJPY83RyWKV2CMnAeSJfXW2m7V3vEpvzFRJ
t3dxUpamiMJ7P8fm2mcnXKhQa0gGAiErPSquxiFzg0pxPzFgpqsUtmOBldzQe7rjqariEc9TI2Cv
DQ5RaYMpuTMDSIKDV52/nRWnzg4ODNjYj4wfwRQ6EPGvEANuzQeL63I1C87EAjV0ANquMNJ46+Gc
nORqMIti3xgsl1DvnoUN6Q0S8jVn+0Q/gsPgFiPwcldc6sAlEkUG7tfnfW5cHo/S5zbojCxU276u
qMjF5u+YIWJQVLexAZrbHD2DMcckVwtkbaXF1+4bVGH82OYCmD3Huz/IV8j91VRYdyocSCHJjXEi
VvEh9mwTDxF9Xi8u6TFceSZVjp35xH8meeakN8hwBLHLnOIE481Wf6pGNJDH3SZsoTN/LXRK74jM
4vwVW51rpxapu5lRBNJbMb5xfSrxN4+rIfVwUK3cI9wTe3UCXg59sA7OkwZNGULm+d+c4iK1icHY
8dFwJhrF/XKE1/Far6vtxf+1EoeNHicZja3wNM4Qq0FSkx8PbCTWeSKO71AwZzVi8BlXNzdUvm+G
maC4wSH/X/dXwejmqm/kjRPmgyVzWX773ugT+i6nFQkxWLPYz53oLfoPB2XP6HGZfZXd79WEAzql
osHWt3IXbTJPgakMs/2X+HLjb8j8TgLYcAgHJqCnM2b1jtoXz4wYMFbXBLEcLAJf5nbgzluqOB6G
umHuW/IQAUOzs2Ex/x/CLyqkJd6VWcl+i0yVzz5U1OlrQ/lPF7DwPnph5WeayHR26NKVoBwm+fFT
1e6J6T/6uRVvHWsBU414jb6bnbcDlkKRfYf8cyDwFprwGuYp3Z+mYe5xKF9ZHEIH15EUEmgJwfOr
RWxEv5zakGoF+QOu1iKhuepKBR9Ck+fbLqZUUofGPwFZ9WN2eyt4ptUq/a3R7W8DSyE9jAa6riht
CbqJqjV/Sj4kDrwSFY5+I5JmCMPqJOdxOX5IbJXcQo5v4ncP+gAWHNw5XTSMNjukW2XpXfmWyjtG
UDSXz0Vjm7pNrExAXjGI0u/wUlvoxww92pDU9LGqE9T3RwwNKPyqS4vrzFYHPboVOr5YehjJzUgr
214lfd3JwqP46zggGXNXfNzRAWAhVUKObN+KSYXiYr/yxglArMffvQIxL7+xYPxCTMQHMug5CWJF
pe+Feuv+CG1IzZ5jGzYDEagno/lh52JQ/Oy/hCd1166Ia870J5v2/1WuW/UY1GakPW/1i+9RN0l/
33VKjqdLq6hlOOoZx1dRD7kOREmboI+Mu2C74Qt0UU7HnRsCgAbzaSCISUXX4q0e5egnGqwZXYnD
uT+XunT9wGh60mXY+5Lc7Ba7cuuYcFudkatPQOBLkSvwjXXiCgllMsYM9sCm6QvbORs9+mxsiPta
98SfiMoe4EUCRZXAkk5Qgg9ThS9KQW+Pc4BVU8fVK/wjjMj8KZUSgpzp7bxCfVhZ7hekXmwMQ32t
Nw4WLESgNLW10Qy0ZjxsYrnefYzCOXoATSAQ+WfGyaclntsR32rJ5CXhOQw1ke2NPZ90OCJTmsRv
VfQ3p8XckPcjuq9GAdfrvzu3zV9uT38nhhSP5gKAbJPpbo5xyGSYiM6ypTDhA6ll3nr02z2iaUmi
5zDZVwmML6iHRnbicDvdHkI6WPA5vO+xpUeyPRTjl61igF2His47uCkbniBdUoSA/l2V1sxBkyNu
UMWjmmSW0N/obPIBnT3M8vFhy9cmfqqrCruyY8hBxZEU0sOld6cHP18IjbN+nEP9lEOmgKcyTa5a
g6wgKLFfnaNE8Mk+P1CCb+77bY2GuL8ncEY5nO+HVzBz8na6ygFOVZ+8/H0SewXozBpfjNFaUjGx
26ddS12mbG1vNR0H/cv4ErX2fIo+Ufp/nEmJDDH+/4ojOMtfb9IAvcnBU6PSYTpZs17S3xej0zER
lFdJX0bseoZPBkLeGyljwNBXOqTkTWVnr1xdkfidIxzoe2eYCgKUsGwunM9CTv67T2+LwEdlIOog
h0DEaof7rtuKti+ff0VyhVCbvC/7MXWBd/cRARx5yQ0gW7SvzRzYCDaD0lHrl+usiTOLkUFDKD3i
zeThxYKUGl83JwRapDcjSCPew6I/5l5as7pKum8YRDLYSb05eQgnam6zJF8zpJTTY84e3wy8GLYF
InbdncBuFzGuCfqH696rpMkpE8J7FykHXiln5DsX9QcKU3H9IYNg4J6jcy286W5SO5xb8CWG8D+d
dE6379hJAmYDgaG1gR61KZX+sEvLR21Nu0WZ9pnZWW9U0ofpDYQnU4kk3z7c9uFiiAPlv1GCMWVf
iMnd2TysPRhQy4OOI3HJDodp0bVG3mZydp2AlhooNhiKSM1ivBsqzkIvF/iu6qklKZUg8qldy3/o
jAERkIO0vv/bGdjtm032PUCINP1hJmvoHu6weffjSDofkyS2l69BA4zF5pFIL5Y91FlVX44hUmfW
u3kWTeQJOI5dpRYulj9fSnHtZ62T82YayrNypTHr8EBY7aHWYcKAzPpRGN0U1UsbTgg1sfQVn162
VvfLj8Uert3M5wMD/rSuqSxJTcgqhn0QNxUShYb8DE94IqvqeNZXu7NZJIDiiGTYrz/FqKQflz+j
rNeIRVeNeL3t+qPFeRqw1vzuGC6sugZE5ap8jlezF9OxJ0KdY0f+m5zq2EcG6m+yIGSQnxaCAabn
pmXBj08Mw4T2JTNpAOHtpBKyy8n35cF4zpjJF1hfaebAQwfh0DBIjISetNANeIIEnjZrkbhu/o2T
zI2QeCwxFVwdjLfV6OtY8OONzt+5EGbj5HB5Aeny0bZ0K63gMAoTDxCaQVMhMvAolUPtK6tjBcxw
YSFEf7Em/3M0x+V2SFWAPwl+//AryLqT/4NVwXJBNtMvYtK1Kg2IZHYj+LK8U02yXAiADJ5nN2Fx
KUPHh4mmZrlUMmgGVlcwYTsVnWbrj1+ihAsQ30Y+gp60EdrE3GdZ3dbbiRgHkuWTmfvYyjRm7S8E
0K4QVwbtAjiSSzTm7CyzVxtmih5F/6kTU2gvLQNJjbnEumrtM57MJiixUHKabc16G/oPTbjsjpW8
LWMzhwosO+On/lecObxt+G8a2tDk/41vEbky9HguX5snFX06Do6KvtuDm8J3bhIKQgjbLO4JNNPm
V02limidTWa78W3oQ80iSJGiAofYKe315ECT4g7kGMDdPhe0vA90yPhRgDb9pKSyUMI4/aYyCEqG
rIRcxUHQ43KfhPXhTPmkrokkNmxDzTux/vg4Rbikq2KJOi5DxcjkVahCoowuP/ehuf17H7FOuAKH
IH86/GvWgIwzWqiI7j3GyGQVtFKrhuDCashmwjmc+buLo4Fm0Ypr/xavXhJ54pAxvCuHmiIha/Ap
tt+wVIOkr6aWikjcoosVZim0TBR2+uxmervzVrousM2RFGXiO7QOSWEij6xMJ6d9Eqf/8Pj/PkmO
IIS2wlyfso8dN/m+s2/1Ik/lhU34AireeqqYno4cuIZKqXxdXPtv1OZsJz2E8AbhtL3HqDJLY4Cr
VqYd477sbDP9Ab8a4P+hZISSTUxzz5t5m2kmq2KLzzsQVQyk2QEBqYmFSeBYFkJWU/7i/pXLXjwh
EE97jYSVPPMhsnK+gmT+hkeyOnE+rR9zXfHfnnM+8LwcXEDJMHD4eYSgpny5YwzywkYF4kp/NJ+y
IiSqDyx8R/Xd4qgQIGv30e0oCliJYrVq4lpzNS5/41/0slRO2zwcjGHd4zohuAi24OijA/wBHaaf
R/hj1BR7Fzud95bayKQKqnOCSMsJ6uZl1rgkYpbBKqdK2iAX/NSiIPnyMDg24fkazSEVYWheEqzF
RAaSbFG6NHTWnqB6euUnl1TKQIaIbBoj56+KyNC5k4EAtCkKjmT4AauxKyyciWJkS4jwR4jzIWSq
06mPJOJtJje5MLMKgu5FHawSSHKOEoTnOHkJsDMEk7hZvhoeCg9JuybjKkU2uzmCT0pJ3lorCdbe
2KiajNcFnoayeZBlez1+HSU5qcSGrlcDx5AH2QldJbWFOwP4/HjG71yJbICoDjLYlhNRZFfTI2vd
sT6Kz2qIhxnNaHq40b+Em80jK9FObXb6KUWziVvhYhF7aSBsOJa9lzLIzdKVCGlZdW5nat8JR9To
YZrvy004VJNdORKzhwWCAANUmI+iEPAlaa1PjIXWiRsve6QNuMQ0LDLDfphx+7GFnrkGV95VXJzs
FU69WXGE0wttkY94D7WbIz7UP8NiEvovJzb5WkiPh32ezsYVPw/1zeJ8Ct7XxE+GEYfxx9qaKskj
8l9VkAhvvBULgocgcOhV9XqI2i0ExzFmETRWmIMDZfOIrpFtme1GrDJRKKq5A4aWxPNXfWJ6zrde
TAI3Bsy8W058of1b8sfcsJY8vuMH++Lo0oW23pVsr/aLTwRWoxtHBrYRckgUdPgDQiajaQfzegM+
LWX8n5RQ4LxFvauCp/aJG62/qry2RJWRh5hdR3vuhkM1dXTxQp7Mrk9ncVrNZQxdaIswbrUERhrq
PUix42UX/cNvtISdbQtv+agYc7ZKMuNJYw0BcI0fGVEXxX8LzxLIE+YuNQPOWvXxyMRv57jn63hD
tS4YDP6eFipnWYKyizRYeOM/YiUoh/Is8nF9IueFn5P+u0MgoaJUk4shnmYR+QXBzvV7fWoN8KIp
ORxJFiwAjKS7L+MNsw4Hbwnx3p2BeA2HoilccqlRcxD3JrWWSnf3L7Q1V7R+Fej9Pj2tizUFHGJn
JbqpINWCK1YHH+XhV6WeB3t7JNPKE4nG8H31EdLs7WCKTs8wdRJ/18nLQPIdEjsagHACF8Faeite
DmzkNvXpI3Da4k1tBXBHnexkVzzhefjvuSWqhLJvA/9qL1pRnwujMVuW7v81fhtff5ylEvcNkBqS
d50dsNHsjkZjxfbxwONwQziAgKrtDiRZ33HINhXmhXX74DZvuCu1irfO4sD8r5fxdOqbwcpBw+gl
IMtGbFfYitYWzL3k4FuTFv9zvGlwn+2XAAMbid51gP3eYAfJN/5ERzS0y2MT2qs8h6bzn/q/iAuT
YKaqIQ1ae41dudPxvapAMSQBsanbBd3JnJf0z4PW7MqzlbBag9n5RB+2HzTjdMozHuCPNGieGvkF
/VCzH+BgAdMfKAH/4qR5FJ+rrcEi9Gebef4Bds3g570ZpKTXN9OkK42imfu40a4n98xaWBRVYB0U
qTSsqaVXW1809gfGrODRnbNHxf+fNr6/HTCOAGLMU5yPWH0jKF5Nn4rcIuIyjKnXDx2zTMqc7yYw
X09oTNDB2SRGtLaOiXml5CJRAMwGOFbk8RYy1tC1CNPhuk18+P0Wj+uWiiunisw22CgP1XlAXNRt
1z9ZjXv5PEEPXVzgXRKMVwGQmx71A/WeDtRrWaEE/zpGF13EC1HQ7SOgVkDlTqEhOqi8SR0nKqKh
ton0repbmEDveCn6kvApQrlUsXmTedRryV2Psqy91bJLkOnfenrQS0/1T1BgXTXy+pjCKX81OY3Z
q+nXZsmm7oi3luX+Ap4Pm/PeRH689EKDCwPx1CRnEDAwQJtR8Za813aI6LTcGJ3FPdb6P2OQ2xB+
QtkD91FBNPxptuF+hdErEJyJY/LDHIXkjAajrkqXWAGDH07eMw2TNH0WzaPuMN14PoQnSlUF0/hp
NIQJiicOYC/M3UUaLgTyMjEn2rnvuRZOvq7l2GV5pzP7dGsZbT5J2dtOylJ26yjoEIbasDPa+6dQ
D6jKgG6ToaRIUa8l3cYu0JdmzmzcmmY6aQ/WkXA/8IveA/OVfLEblohfEpLmNlF8AwRRta/ba7sd
chuVnaVrRXsRwIJdVetqOtQi78cqkUhnBJ2cOVGt4z5TCMOB+qqzceqQ3StwzdmLRRGKiHTMUsfP
D+0XuW5LVyLlTVKFdROBhCe22fJDpQacBFedtUNy2QTyWCRLCUSEpNXnQ/X5zOTRphcOvlBaoWoJ
qt9mPC0h5GR+rP6zRgtyLcxbFXDa56y9m+jBVsJRGorvpYZrZF1yEGNX2SvcOK8b/8DTPkiMjYlV
qYdXvsmhI+E8lu07mTVpxFvT73BL+LzjHvCHo9/k2f5TFuRN6Tv9gk6LlkgWuqQ3/WCLcw4ilFpO
QxMieEazfAqlv9RjDrqB7D8pIBmThucKTQzKVsiyT09A7nwhwmxXbDpdVe45MmLm0nzdJ3HEOvdU
/0AmqopqC2ZO9gsfea0/Gd6K96z0NDxHCMRj9nhEj1NSVXk5Cbe6jkuqfwNCRSvArUJPlWbnOaHe
3o4deow2WIez0sIsMeFzxth0Ag+9QX+67q0LvdZ4TV1YfcyDqeWIpm5QoEtnVfHsgXC5Mdms5eXa
Ob5qpGEIXYAbHhWo5FH2nFuwz7SEQjrIwn9NF91Bt/9ttMCNT8lqOtwRig+x4lYaPIeOZCDjH0/a
q3KBiwWtTP26JwudlTRxvRvcqJaJT+j5/wI4pp+agHQVv7AVzo/PJrkhvTYe43CRInIqzqkxuL4l
2ag8E0+8A48RXzM7h09RpJo00GpUejgstayfCl+ypCFDVQtTic3xkENvJikMNfqDn15jvRcCKKIs
71YGNhbQZ+29uJq0zdqJI+CVDulVSmX2JsFuSpoMEPh5O/QA+w+GwZQONun233CS248ov5wAJKgJ
R6ElMgSRfIh1ZQTd8HY9v+g7oRxt3NHruHOrCOANWnDH9LD7IVC5dk5jzgFTzaybeV+rmG8Vlw9B
UfE591L+zdRyQe7aBWfrIP6lt5esDih0XltOQOyiFs7RAQN04jOr0cqKwDNojc9W+fT/dZ1w/8LQ
oowN3F5SPV0Jm55rnTKoJ4ZR7x4hXuIqXHdVrkiy9AOBQ8hp8PKH6/ETvpMQ6UC20cEZP9uYMOel
CxJBAOoATC3/jasgJJEOy8SuXkMNvGwxhcNKIROOnCfiBqmo6uLIhNNliVMAsV7yn5bVpCc4dahl
k/wCfHlFWOqnQBcY/3Lvwox3XE5zuUeVcEBP6mtQUNXG1r5POoncjFIg6U12w0AsQNJaswQQ2RRQ
B05jCacWfhPazfZrEaEvvzeKgYYAKToSHijJxIqX+udndbV0WSOUjutgS6pAS2TS8Jti+kLDfTnZ
B3qeDXsKIypxg88qV08j0P0RA2alX5JMKo8ufxY3A0NTBj8a+MzUEiYjqFwLd9zCm1vwtYDmqbCe
1lCYQL1KVkxAbpwksBvDFvN7lVPrCtmZqgjsYQp+8nKni2bQPSAX8tzlCTAb8W3Xo2xeN5l6s0we
12pX2FeK6K0+XGDNv5+lZs6PHgm3enxhqlYCPKtlJd11b0XikltcGCf6hDR3T0MisNw8JF5+Jg0C
AUF4C2ZAIY1LicIXtxAVqVQS80fPlbnYAhFLEvpxrvttJbK/Hx3v0p/Qsaf44Y7U+zA6WPnP97yU
4tlQuUvLkJN784cEWwVaHUjY5YWhv8veX0VQdBzEtSGtjZ65Q9637aKhv5821qPKm4ufY2OBb7nh
fG3W11HVKxi2igqNzkY2sySqXJ+fE9igmi9YC3vyTZCxuiRZE1Y8Gol8FrPMVfOSHg42mAV22QW/
IAjqSggnv4zEy25BUWl0T2NSyLV2akG8BgcXmWVYe04QSFIPW9J+hmse2g1wEkQXHdVF0k4MXnWA
ti9tQoWWntbT6Q7LzSLszLebpo7S1yX8rtfDhgQldA6Hf3f19ojz1HdjUeulJ1l3I/BGYIGlaQ+I
wGE2werr1ZfpkIjqtN0G10YkZ0uZ/+jSj2805x8tQyLlgHPP0afB5PbtECkP6VHBo4t02FPW2gyq
Y+Uxr6Xt2I4ZMrFy5pTKgXF3rkQcDmfiAlTV6ntGTiWtxsmXtAJXa6gm7OJ8KSw/Hv4bvTOz3plB
CfH15OES/gQJnDsLmQM9ELml+RuKilA39Myv/J/eUEpuwWe3G7yLTrVoKBKlZaxOjVizrHUh9bKV
vABP9DnBINCVKpQ/GtFowpCLdatOGFTyK1yYouMyGmaRfSMMSyVWTJD6zILW11H705tULD379jaE
i9Wn2csJXu84W83gcJ/H3yYx+aKR1FRrNy9HXkSrNlm4CUDnxlkaLXseATxUGQX2B1MflUhaX2/O
S237S7CoBN10+3tpVLNYwfJraMnltqtMxM8Garz8BlFNBVNOFv50A0zTZJK+vDyHUlbN31o5M7Ge
kZ5ep6eKmwK+8LHCXcG6EZ5zRjclWOVUF6J6Yr0oc8QV3FGuouFy37Mb1h0uMJinGMAPq7lEFU93
p7pmGoA+9Fz9W1wvNsp+8xr4hX4pENdpOWg0HWLmSeSy4PnO3SIa3dM2YPj39SXmqK8VcEHCR1Lf
MnXgTR3TLVWRO4dACoblak/2fjdrs1jXZN2WlUZ0mdvfQxPfy9BmfPIoqO72LsynQ4+61CMRhcER
AMt68oC3EZopuvJvjpvSZElh4B5JlCXMoEUCBkjcv5ZGhk5yWY5Z570mZ6ic8jSFJfjhzsvyYpZx
JRGnrG0XfHRAEJ4WRBppdXo5t3vfCGzZ47VpPTEMfv0z1qMt/Hm5Na2TyettzwUhBZsVH0AQnugr
0+0QLUsOmO+OskvzR3wHOpnMb4Uw7g5J/1yXEpv5vbTI9aLZU+Qo8hSNdmdpIWE2tza/SeA2IioA
9QHQ5G2OqFKpWCQe/bc1266W7uP2Za6bK5+C0zrfd1u/w7vNEX0899YIVgMIoxIu2qrfuIA4y1Kv
0irADeNY5Ck/vqou4AFJYOp/hquSCdL42Pfp2bOzQ+qRkfkGDJ4IIOu+t60WPKjjn7nlfnr1ILDM
e2nJ5GFjikqJBPVSRbBX2wH9QK3H6+MNEXTAHk9ZHm9Ecuimq2uWNlKgu/EeSfLBRxbVHllajXkZ
MmTOJsApilJNPKQo/nBRE0U/1SZR7qLwknYinED5SGHMML6MSkmTGke4A4oo0w9Qs6KhyjP+ZtJN
frYiMwpa8ZDc577ZhJcWGVxzEueMia0rhhJMws64GfcXa9uV/FpOZ2P3ZEW0lwYqOXyLI1CDfbnw
9zHMx46MGUGsMAKMyCaRGRnpCbaMwnxaJHbmPtIO8vcoazcMJe1xKlING1/fXiHysko7lbfM2mtq
8YcZNZKdDKzD4QaVU0717uxhTCrypffcNmXXNqmfJAKtDADM9FSlH0WHUDSGz5hzIa6LR2yHH+hI
OFBL+7tXfMLryG8mmAe1+u6Zs0kh1rQCGrRxaADP4mDN/NsAaSaABIVTeLbYbS8W3XSNMmSMoZ/I
+JkG4+Qca8/qhN0YLWP4kAYPH7YoApcGGzIemH7PuhKlC7DRzr/cxUBniUusGKkHkdcAFmv1ZN1H
PT4fY5OO9SAqaXAn28XS4XN7qrixoMeMvT1sk+3IJsi4k0VLpYQl1Nx1muAiHD3FcT/mDZwNQjmx
Opfd3kse3sU5d8scGinTO8WNYVVSWOHUbG7DX9JrjgpTLRVu5eD1XDHpQH8czfC9+wYMUzTTMK8l
ym+oV1/iQy+sXcYusGrrMqnLTy4Lv7ap1fSyBJV4mo/Q23FrsN3dMuqsT12oYCk8VR3PIRVPCVFY
xW/MhWxsGbllgnL88ENQm4xyFG76+Bte/NS08pqdMEcefjOlKai9GsQGwVYPvXhf05HDXOH49mUY
r2j5hb3qx1w3u5RiC4wW7yyH3T7fI7t+sxkdNsnkJsA23Vb7izAcQVoiZ/yNTRYfR4DHcF+6FO0g
2/U0xD/oMfpw225WihhYIcE75+BtLvzzPsPPIT5/qIkJXpRBKnAnCP41GJRJE3l9SpJwYIpm7FiO
ic7Vdktge6tDGwsXQMHCTvTG1qLMzfwwUg9T16bNIPY4dumz1NniDDxaAMrN70YRhb6vFWa+6Pvb
bzmFEibKFFpzlM6D/OaO+evb0YCamxDy4nTkjKmH4oc9oFSJFzOEblCeGDe88eWA4uuxcHfKTnkQ
wtqedY4cT70DQoFDCi3QCWhdEAiKGC/+5xMcb0r/GXrsrQ69wgxeOxSryJCm03crwkjFncjEJ76g
IM4iUHg1h05bgDY3xlESPP9B6RLctrgls5fJOYH7u88BmueGldRAYnNIte/3avLk0sb648APXSVE
Bf7vqfe5MXST9on9VDNcTbViG2BXsC8irSQ5IBN68AKmvk9nibTDFYzbmGXFjTeeHz8N7oKCPtQr
2l6Gb8IzBPQjiQ0b03EjF83iwTdm18diNAUzkKkujetgb9JIDBS2MHuxipABIT2T3B3wbXxMINWz
nZc/gf5/nNpksmFfRsGPjcRlw+YX8ChUPamg43YsuSdrIX0K75J/mvdnOzaoLxRKTCC/06nhbdCI
46DeA6f83PqBv0a7dGbwbJaxwN883C2erQT4QaHZILwUccvtLz04FtDvBW2f/XImfsDrSbmv7hVE
t0erhgiekfeLv9BkmRbtIOLZibGGtYvqnFfYNAAEJZpocdCN5GkBs3t8cIBH8UtuVCc4NiJcETl0
vo8YMrALYD00JKG8epQPn7s5WlEGxmjKKY1Y+PM4LEaozzIP1YrQz+/ZMz+X/8SxeBLP9bdaDYOr
ECm7/4cSzL69dqNd44SDoHrOzDF1W7LwWEM35z1v3qDuCHSBXVBjSk67pD3cohe7iz+idK/azjcK
6N608RYjY71CsnSrEyF+4Y4rOt286fO6pP85Z7zIpqRRMLN5qiqrdMBteeRAK2ntC9mG7AwCjtDv
D0iUzFdvA48A3bhlxp3HYfCC1Wjj81QV7I+wbsWnsb7qKNvTA0HKoW591g4blrT7JrS2vdMxM9dE
BlktO7nGIN5wZ0p6B6wvXDaypJ/nrq207iJbJNaWspQELvYYJ//qOyCAgb/Qo01OQOdrBhqKs+uF
nfAVnHjOFP2MSc8wcXm/c+uexgca+yqaglzahVOFH6MSl6QRiVLZMKug2iqzhyHhsW6uqoLncsmi
fqkLtCFiKdaUQNTcWawBYlh1ZNhmI8Q4haEscARWRDB3OwNFWqbxvSnOhjUjYs1oUyPNVx3rp7b7
GNb6zipwR2J2CTjlhJrXm9fUjDFWlOFXo409kiauodyXtxTXrVdw3ml2rBAv9/zScYZ5aJxYgNWA
lVzdXZdevUjIrKOrvI5L2r/XQ/+IiKuuGsCCjZD4eBcM6PyJYx7DRNdmKElofnsEkrLRxrSkf8y/
/igBMZlcXFoXObB4W3ZLzkOOXr1s+N9u8a+5XO7RYHKBUw5YnOe19FqRCMN1KaELjlyeM8gsJ3GA
JsTfzyP5YG8M5uHO0azxFiRmloPsdqk7EQnqD05vGXbSd1MdwOQL/6jUo6947nNNA7yhBMAY5Yx5
b6CVx+/1jawQ6AFGceSd9Ub77NyJOp4FtX1XP8KYp8QuPWfOvUWcAs6cM4rkZETBw1UIpbUMBx+p
oLNDR8LIFNmbJ8csVwNklpnbaAdLiyqAGY3Obz7rLTw/SBn3EN3ie0qlAfzixcYIE2bHQjr9G9c0
GPQZBrkXislAmTEEplfBm35PwmlitJG8Jf5RbS0WP53Nz32uFu4WzAwqVnIFkjVRslPCOdyxBgwS
nyUZ59Gk008HWG2bhS2o/F8tZ0crPmo0DoLALjVH8vUksRvdAfcwtyXR2/OyG8FiGxY+Ry3EUG1M
va7oGsvrb+F/RNNLGdROcyXfe+3qT2AoSVqfw3WO6+sFbhU8R7eMYqLuC3rPQAxWlOLOz7Zb5Qe9
W4fM1yHU+xi7jMvlfbvkqW8dXz6jpvLR92rcOhpwSblSthlDaGSMQOA54qsERM0QEDkI6kWueQOV
EZjkzSCP75JNIxaPe8KzujQHr5FK1Ioc1KgkFREV8TEhwgaFbEL1oNcvsfONseAEkIBqwHibHswj
MPdtTthNNm/o50SLfJHVGNuThFXOtBw1NChvrQru/0CObxbHuLUhdjI9vO7FvbU5edrj2We+qXsK
alCj1Tn2XZnakjPzAGdkZP1Kgqo/T4Xe7WIHiDt/7HqbBMohlEDKaiTrFZIdGcFfewIPdIUcnZ2B
xvIbb8a/6TVVDAThx5lYBzvVTIXri5JVPkvPx4AlxF7QrThMbcEigRgtpZPO8Nkzr+0M7AVMmx7x
emSN5K0Jf6VbYgIRtQC82oABPhv/2SJscNxtgxmKgnOCJ/9I2+bd+3alh+e9EYFRPX1Sc3ysaGCW
fgSsKPuMr2zMJY5vQBPUwyZAJ6pnFGSq4x/qFUiPN/CaJ3rKJVJRUlovChL0XPrrxsHS++aB0ApJ
RAL+xxtfDrpp3kGoCWOLqQEke/C0bsTC0YDdlfnleHgGeBT6MgkCPFTLg8moDMSCRZzK+5K6bcWN
WFwWUSfo1cpQJxNnyYtyMp/00T9oFLyHsTJf8N2waXe44uMSSCN4C58a7qiAN2YRYGN9G7+9+N6R
3u7GpS9sMEVgAT+KPjbQOa/IX4rLMsI56A7HGeBa8KABt6PtIA3/oKyjzPxMsSeeNoFduIp0lT1u
P7y3AQei+Oq0ci/hvaf54PCLfDOj5aewhkN/hNm4r9iRcjlUZU0CkPU/B7ky+xQk5BNz7uP3uZ9h
r1JPFyAPiGV8Uogyi9+Io1murSUQPKRd+jgQfo+ksv7HFSOATZ459ZpKxxPYKhOzf7H3zwxduFhU
jRTcHf8UF4qiuKECk121iOeeLd4cwokzhOW+0HLQvsP6H9y788r9s2UpFw4Sy6NzimMO5pXfwzXm
2Na0+7PFDmUdJskFQE/kJzvlqNLRIeI4CHmeRhmEMy/tQJHKOhWs+Au/3MpRdZl62Vqs9IbBwMwT
Jlp68oqTGJbVWpteTovEHhh0uTR5Lb3sO6DgFxnqyRy2QBFFSQvEcgX845W3wivj3G90BxB46728
6XUALc3rkvr5leEcLiWAg7l7ILlCsrgLVuKjSHDSOmSEo2+aXiGB9nmsh8mh2Gqprf1nOgaOnGkH
+CqfG7nR74U24DgMKSGFDjjFqf2Taiar5ZZlTBPtsi8bo8YP7RFUNNusRWVAECJN081vW33F2pvt
83Z2LuzIU6nAoNXaDPfdg3Vs5gDGYlJH9eSik7Op/FJq4mEw1cq9wdjyYmqtpta9NHtBnRDZuNeM
1QDMSxU7P/PfeW7uvkVQZ7L+UTGZHm22nNNGtkt1GSY1IY420dpeY7iYcResYM6peXjz3pq6FfHj
bLNK1iR2VhVHDNiFRy4wERO9eS2mocKad3bBK4WKznCLjbfaUjiVn0NaHxae78UwgKB4HqUbkrOU
lrWVoJib1OTN894SIfvYKOtCIa7ek3qkCJ1/XwqbQ5mzXBce1degddJZPNuW4Z/vfIGR1fwJnL17
azvPHIElqKn3yI7UhVDnWVsm5kf3BpVClewJOaPTn4Omfp2UXvZqi8b5Q2BLux5ZT2KiH+2bNJGF
Y0HuFiIRwKRw/gLJZfMEXQJKbDkPQNVqMusxl8jOEuYuEi/OevMsbjUc/YP+whxU0E5FTow88Ji5
7xgjK7SjNIeHSsBP8BlkLlK+vKmsLQlqsrWYxV2juggszuG251s/8Ox3WoywJhfz3+l5s6qiZOq5
4FkdGuRZKODz42sw8HGjLQ5mazPVm9LzV4QlW8mk49iWtbqUrMdKg4yPDlbMFOIT14sv0Zk2Aom1
/mQGkVKCGeq10fuA4sEqpE/ZlWOsvs3VmlyosrkvbIAHG4bVXNJsxAB3FN3wF+4MqlDDEwwGMmiH
4nyU3+z9rVDrN3d1PSvlFALHUSaHZSOgsTkZth1nR03CKvCsHT5ZY03yqpfinnUPhlUOoRtAIOy7
0U/1J2CDAO9OfOn5aWLxWPCjykfYqSfRwJQPe7/NfwYMZ0rSKdxU/1QCz53jKESZqrnKdm8ZyP/B
Yoe5XQh+i2XeaDSOl8qAVAy8dPVxKGruck9tuGbPStIGwz/3Vysh1rAYR2NFJzCIZGM3IAEDz50n
AhfVCheRMeOSOyhPvz19Vyf6x9Hxj1eZ6ChVdL75PjbJOX/LN+dHPONFjaCXlj0zVCO3gKoIuI4E
ByEIXGVHAQgVYBuwnpH6pYtZdrdpD8Lcyctbco/UJLUaNELKy8Ixhdmhxxkrti1WbVxdSIXs5qiE
dsOeOQMraQgmuKoc2XjEk7AQ5A8NA6ovGHbo6NYaHjZ1WSQuCiM6vzjPp9S93CjhFo1WE3/jZn20
jd7LZmK/MdKYvq81wdc3xtxg3v7RaseqKBCRoHkimItHRfWNarAtgcrCgI6dwLeF2g2NWye4b1Lc
GXOHQg59YUR2vlPC1qRGQCbBF0anarfJ+ZeUSJO7UwIa2kX2CDCY1TDiqe/JpLay75DhXocR+GuS
GAtjXTfrojnS9KHME03TbpH1iQ0WuVjPlXRRNAXa7vjcYif7V8EjzsqFBHT7oXYEmQKFaS7Uz4mt
12PFFJMuGjYf3T7Tzb2TGP0HnwQ0s0T8sdKNFp2j983XwDLN8XJaFjJzCtZn+fTVzU2HfQnCU0+8
l0PtdCKHw9+e1KgmHXZo/rTzON2Sq7Uzk9/O7Tx8P+CSilz10AmEM5DntoJd5nC0LRg0dqTGHB+y
pI9b4nH462tfgdFoM81RSIgD+A3l32K22z0p/yJpkjytgWA5a0OTCNAWvEbyCTECvZP+vZEVyE+E
KG4CKtdFbXAO8XybfLyg3jNJv3bBngIGtA/cK69a0crexA+uUNa4KO2uBXG7ddXeVmfZK8IWfRSH
UQ6Z2RuixCjf2qb5E4Q1YJm9nLdVAE5s+pLO8aFB2RzRpEaOj6fDjztz+eW7dDhStR7bywMIOK8s
+t6vKsA3TvqoZWbQp+hxzWD1rqc6+STZV36NjzMgWbcV5WwcdV83z+5PNeNUIEbZBFvF/mO+y9ID
6j+AthTqVljlItmswdi2uA9nArWJx65PKgKVh1ge2Dy9aSct0/QGTfTNBO9Bemcg+EbMGBGGGN+4
LaMc7ciL6iMFHiBbUnUbycr3FqK119gP0/j7N1eAIlfE5g4pieeL8ovLSY9CvpVRd7Mg+FsgRzam
6523jN9wp5uR1ojRval0DUF/LBbBC2I/5ZiHXKDQJh8sUH9qaFT9MatLlezfH+vmp09Gyrwhfr+2
lwZL0GA3sy1Cv+IVIBOUXFt5VWDr13Q/KN+0kRYhXfrk8d7mhBEWLfPyRoAArQm4+UZG4GrmVb4B
B4d09cqQPXDWPRlXfbASX83btELwzmLj6MftKiJJDY1OAXtP4FFxIFKJxYX0DJz6zwP3syFf07oD
du9ly4pZQ46tF2jjRzItSrrBtRAm/5NPWnwTYXG7p2goIVDyQLLnius2gd5QwDisS129PUlLdAh8
sxcJeHhH9bQ3v9fUzKtcYVZom90IFNqZxLyxh7jnylTziIGXiK5rv/nfIaf6bZhMSdEVHB8OupXk
vtaXfIoUKxIdtpFsVWa6U1/dlZHm4zBPpIEOkQDB1fY+8IYTPfPK9j2lnKS9BU855BSzEqKxTIjP
wn3w3z1O/R0f6sQKEZcOJ7LoftjQ0yx4rCSpz63vm5/2JVxKyjdTh/IFMNuD4pF2jvJJXjfTmeFl
CpT7Ib7zulxFspX8+i5dDvn2X5Plr6XtKGOCuVTPd0rly2z7bckiSikvym3hq5x8UAQhw0idU00A
/GkqFqhx+Z1TmGajwVEeBy9fFaPDj1QD6/v/3vxoAGwaRPt2plF7tkclnJASZQn0beOgpqEqjZ4g
fivEFL+BqPs93BpZyDQYAu+HPikh/ZQyO1oMtmG2rOBYjoXTMRb8Fyj3lJDLPkpz8C5Dde/goDhA
bS39hf4/8kj5KMOwr/hcxRt7jV+H5a034i1FKa5iSUUL4JwowLMsEb+yIRMlF4CvRdTq+ucMWlCY
GsiWpjOj5hE1Krs7pinFFYaq7KueFKqCTwnQvKB7VDBFY98kYbhjbKktNX7HpDrc3JtjljKGxgTJ
Dyjg9+f6Zzq7Mo18TtOwV6VeQdkPrv+uwznUWZP6m/QusjoqQ59aE4XRTbzwhapi+xUJmlfLCoBW
7xcZHby6v78MinwNfeja6ZzesUjNv4sKDGkRFTTpvyeDs86xdhE/GPskr4Zot3Cbpx4bIZsnBWGp
PVz+eS+NBvJdMLPeCnqce1zQc5b3s+3Lnn3wCeAWc8WOrmiAbFb7rbtkvCOPyWzkRul3Bq7YAceR
wtrxWcxh75nldk7SW4exgWaLw/97LwlBqOY9d/Iev/ABMjoY+8x70kOA65DsEPu+s/12e3nwOd50
dv18T1AGWwO8f+U5Fk3QRTfUX9YmztRLVSvTbzQo2CcO100TL91liKWjxpefTaC32P6dPTK/GO1b
YQViU6yPb9O02xMtqK+1durYgPfdKK+sYrfIgVTtsl6zhvQk78oYMPa4w1xmf9Xu+ZRcPbDxcEu6
iy5TJcdnSdiCEc8XLeULfBBoKxBNfr/kf7wIiB6O2QHbKifW+BAi9G2J8ozvQs2Bzbda+oy9+UIV
Z4L8uWDzAjHJfAu3RVaYVvedksg7CWvSWSSNgkqwhVBKXGILiFJxM4gRNMyHbnhYLzkt7pWe6+Hg
ByC7MtqAfQqrxBvJFU/FWBykfga4cCQhoUfyuSTZ8L8r8cqQ856ebFQeyFDLpXH0mTYl5OoQGp+I
1vFp2Iu6NmgAyeOqybKKqgwBadKmgGO2Cyad+3jLKTv3y1IIXV00/EdaXhlJUjJ2b5cXxBiyzXG/
8GUqMcvpuFtrTNaccFBzJK+kHClVIUPDeE2e9c5M2dxe59naD7if1BDE9MgDyKlj7SFlP5z4B96f
iiGcqEhBqryxIwLrDnrYHg+uZ6f3VS+I2rA/5snW7CFAISy67v6wwi6qYnad7bZc637mc6s4SSZQ
OnLwcXhQ51w874zJQoB6WKpbvXZHHVz+m5FqhPRP5t/tL42GwZHerFVk8Alivc+N43uE1B+D278i
Gng3lWaXI0u9kkPXdyW1dRGySHW2J7Y5TJfSQhSzKtKl6Egsy5PWErYf2csao/EGAA5W6hKTZfo0
x1iPQ9hT4zJw+AVLkbETmdEQrX5f9b2EaEoi4EQe21e+kx54g6JCqqtX1NWkGjiUZI3M/geSGw2z
Oe6D69mNUIQ14WSeiQUEgAsfEvaiaHCveUhOIXdVAj+r3V+WgNo8puajFkPxAV/wk4EDBvZ/9gMP
HqAHmni6UMMTSTudrWFQwoQa7165TMk7kYjdep/69fj2upd6xkwclsNlnyYc4mkuhhoLACJuDB8Z
d02yY9ab4QFmWMwLZ5ADByombku50mjUbh2gXKh8THlv73uychV6+IHWcT21SYu5BFVcfv5mr0+e
yzQ/cb+hprXfypOB9iBahjz/52sR7lelnPOj0RdV+c1GfOPobbfanWrkctD8fzDw6NoQdLQVR0fa
N/9Kmrr4ITtcAHOLD4XTw2STQhrgW4aGA0aM/2hAwM7LifnVoS7+yTpal20sqhuEiNOdOSCFGfa0
xzl0l6pcs3EAcWnlav1cSHjIbz53Vcz3elkrencblSRgRL92OzvkTYpKm5gmTVbY8ybIukaiN9Df
/H3kZTts7AO9XRZ9ecKjdbUGbcefPovm1YbeYSC2d/XHKanTIzikrB0/B657lhKOPYYh2PmtE71n
cyTIIvGxNmiF9rvubZzXkeJt6YnofJrBskN9/PpCnx5sJ0QlWUVT2l+pNhvX6jZlY9bnzMePL3Ma
OmSIK+CMgE5oKToSlhf5QI63m6NfuzVF7g/eYIA8cX+Vd+a9EtYwefontIxTGngD8nBVmOVFhrXm
qgKB/YacE2H23MS6ECCryIHZtTAcSlrHpEtBt1WjQUonxX0RBb0OEXg9RvRcsLQEfSGZZQgNH34k
8+bqahwx1Ad2xdRvh3U3Kyafkz3WQjSRPZtGuE1rLFiVVgdHBlQGdFJ+U/VXRHMxLWpBIquU2JiZ
Zkei1kaocqPKQcEBuevjouVmPo85PZyfKKhdfx+pr8/Jcg5aVXBLWZCmJUUOvmrghHTepsbslxmQ
d1o1rMpOMAMkxeFRJm3tSc3hTSOBjkWiDiWaURzau98O+EUEF/9VFdcOI0X5pmSYEgay5ZJsKKjF
XhgAP7EA3UB89QIXLCKQg7VtpOJY3pgx/i/azv2uO628iSC+Sp9GkkDMCaNyXwxsluRROefppDdI
ul431fr8BPrX2mDbJdX4WhfUQZBGhJg8jPabtYFk9dGNT0hmJUaeYY6w/tBZEUviVr+vP+2qCrd/
zl07acaxD4L27B58i7KOotsA7GbG1e3YjkGJiGpXcTBOh+IcEK+t/oOsBK8sF4mAxEAB6Mhr0NgX
mLGHfWfS0PKbaDuht41JKiQ6syhg6LGpzcr3ncPA6Uv8JEpbs8DXakttbi9lSB8nhk/mc1Tpo2i8
WyIdHjVeyX7YlqsKnYI8O2mV5AegAvVKrppclgdztGroaSJ4eCgUP5P19Kr/KwzHe32RPMft3d+x
NwYjdq2cZRazY8+dRaOaIp/u4L6Q9ouetLUAqTqPxjwhO2WtAfEHO5FWCkpL+n7Xmq+s+ykYQnng
BRTk105Mu4bjzwzvDHEyX5HtsQggvOKCFY5psfStBKkn9tOTWdJDxU8HZoCcO/DVTXPMqEwoYZuw
lET9xxCV5bxeBTBjeDNOQFOvE/nhEpRFKXLI9FQevyr1lMD51Oyxz9Tu2FZ5FVZjon4PmJPhirn1
up4wCtrtFGqTxBZPMRyb6C1hDK56yMt9un4qrNnkM9RswRXhCssfJNRcOzyfqcd433SuQYktqQKZ
4Dzff5vwtKQVrkinVFZSVc//R4Qn3oM1eoXwjNA2cHcDxXoQHVGPOIILN5aY46Pe6nagAZGNNfOk
n5g17JxNzVQ1vecu9vRLz3z7Z0Cw+enPX6xnEOqI6vqpr44Z3thrVNQcP+w6Aksq3LwycQCUiMGx
gUwrs0mxyupyS9ejG7gllMbiExqzYEJpaSCcK3L8j2JWcjxlOlUMezus/3n19+9j/kP00ATnI3ha
3Xp5+Lj/EGUwZVeaA4wsP4Ko/hdGvuQDLpXkMLA68BXSQfBwzU4ezSUTrMbkDPaDaaWpM7KZhENn
PzF241r2PYDV1UAIuMDBXqFbs4oI1+fwUs0EDL1QLCNSPRKh2X2MjVVAbYMFfUv9bQH9wuDiYiZs
rBzLApWpPOQPgYqenvVjb+1P0MlKLpQ9rwMJZ+nXA/u1P0hll9JcBKUg25ft4LKPOYzMMfJzbZKD
QW3GGmS8xwdJrUaZMKJlTi+ACkAnBbpyneCTUQpk7FLQUluBJUIZAm7ROpU4a52C7ZwHfiLzZRf8
LAWJBSU32WVQFFX5EbbCKuT52z+lR2QXHNZQFngr0bwUqwie8cIwpNcygLQTCH709Za+/8UDXLrq
N2fy/XQPZwjQm/mOoJ6oYtIP5np1GszQZzScIsDWu0fqPnATajwTLhVatfMvq/A/+MfrjwjSUAmx
2BUYfwUqnPTk9SmQ+B9nGFJ0cZy7p9nE6ZGgFz2rz53xQwnSHDTDaTfjizp3FTjcDPKvO0LhNLoN
N3/J+PSsXXSa2ztvOdViGIS1cHz1nmiug/TjK5lJ3RzfBGl7VSXspoaLpthewTC23jZBsyCpfF1A
ELFtjDPwOal5KWFpOR4cmiJV/crEtgE/8IwGN7lsYSofny7bXqR2z9rx8ljE7rwQu4phDu4I+p4d
srWNLyZOQFusEj5W2P1GVt0VPcJdmvwRHxgZxR39aDT2PblpcAOpXVugT+iO/0SeX4cGLTiQx3Js
uHCVwvefUQei2vabDJ11bsaIE2maQb5mlqET2dO56dJJCyC8Gb+BoE/9hTm+7nuTfuuuhZuXgHWQ
Bnz7OFmsHcSdZKx3JFlbyenXkDBNZCAqI26dgas9q1xp0bSuGMSJJQRz4dAs6EmPTt3/zh/cTgau
9vqfkofJPH/7Jk9RJtvcxXSOJJNk2KzQjcLXye9x76xk0mJIPUwlBkRPBkZZu6HQdK9p5zuYRk25
E0KPzp/SiulV5TorEStQRdQu59pgk7frZfreX7sJDfmmoH7+0RLCut2plc+jyi/+r5/FDeQov9q6
52PIGKRjQGOnbirBTQ1MyQSW9vpjJHVEPGHk6sB8LsNRdH2wZZZhB+1ann9Ja7ZY3ucTaK0c3rps
CivuObbu03JLQoCECQLYwhBimK6wB9dE9ZwwPZvWo3wxpkGrgXzEwuVagD2B4O9MgsiHuBDBioUH
sGTyMRovK/cV1cmd953dBXUxOtZIJOKO6OilxVhceippZv++AyEr/PSdKtVm3urFX9KkCjH0+s/J
9Pu374kkuqNgiBSRg8II3ZMzTbpNBgqLzYtjtHlyEGnELm0TepjFXAjQmMgvyi+eUamm3cKlMMD0
bj72krO7oUrrwmKu3xO57pzJfZW82UqMRVwHiQbDMI1Va09wnk/ElZe3CO6ONLiM4ezoOIwtP3aY
BokQ6koHguwC7wDR7Hdxkmq6iBZ+XpFYKLD2bXiyX2JvMcfnbzBd72f86eBMAWgfhcqm/dU2nYWu
Jvx7XLXKWf7wLE3bHyXuRUoqrANLhPLDzpQgylLJyoGkxnBy+kCm2DI7Ned4DNvQOMhv414y/D2x
JiWx/jl0EggPKyMsD6cY5vy3oDqzGSj3O47X4/NodG78ao03XlCwwUBzze2goJ6yE5tKloFP6cb0
JheGXOGuYnXO7qn8XzsT7m0i5P/XtJcmjOf3RuN7iccKN6IY55pgHeZvgpi0OjO1BhPeewB1i7J2
0SKmu0kwxwi5kO0r/gafZxXBIpv4x2qd6h30rN8tx/L7NnopD202pqE8UNR1UElhg4cTKFhOmKyE
HJi8p0DrrrZZMqNdticjxMUYxy3DxeiA4ra1oyr9fGayYgdBbP3TNseJXOduMDVgSD+hPsFvAO24
PTZ9U5m5XwJpkCcgoWETDdjma+0iH6uppnFYtfneyjLhS7+LrW6nKEf4GHqe/l2UOUEmQRdAWRom
isKWKajN2VGE0RlGDPZCitGnjdaHY8IbOjppjMNBEgwxjxq9evLCFnacizbQXr7ZmKtdbuXdUDiU
B17QWCKjblH72eI/lLa93JOrWaoMEyrlrM2xu931NbQKnzA4PRfiJl0jYUe8KB+r6T6n/ywb5g0j
FA8h2HSIzUa5cnP3PQ8dpgGiM+oVh91FZqmhpAdNgrs8/DmseUqjayQnjn6UqS0qqsKp8Ry3BHDx
nxUP6OI4zle8yZ5aDH+hUAVxcCKJemC/yPQm3v3lqNPhBZU2KgB1qH1U+cmTBR8IKMYpXFI7aUea
DGckYH/AXW37G/1wLShnv+fl1aCfx7fi/VS/7OHBS4JdxSfeBxSPZLnCwYrtJOa1MZJlTrwjxUlY
c/httjD5TnVnGpR+Z05GVk0iplrbFdJSGSSde9CgHyKt64uo2MJViueDo97z+HHRa0137M3SzjY9
jgq1Zm+bz6GyhXWAvqfx5q+I9pgteW5IWkLpeCuT1PSTifWuxF+gnTGOAIIKWtJGKihCYK+YI9Ap
gamshBgLAXTYvbeQhq4d7c55J3q9PPQ4x1RAu6iGcWc2e7h9NO/E9bElFCNyiegokcA11swuE+p9
q0qTtRanppVVQumwPmYNLGEahCytFMd4sRtVwq3PF7oJ5kw3P3X8ZQn6/BHVL+p2IN4c8fQBjr82
LdP6UVpcAaebTT45HpwtJ2bNvJeWmdABJaNp77xPAbXZyCP/NGh0q+DGxhdIi2C0LQA5kauaeyed
N1RyjTOdyPjtmjiLi2vtTpvZLbpXd/r4SAkVdFz8VzEmhKh8Rctx8LgkSPAhFwkc1SjHaj+b81Sz
Ci4bdlgA0gm/1qCD1kWC7DkAtHkuuHw1GrmqTEffMhQu+zTXp4kVCA7lPht96RoPRJs7usA6BPL0
Af10DbgQb4n7rlyh7FHc/liKRxebmShaVOK6IhXYIb56sTMXJvTxYhK4KqMlZf0eqs6+KINjpZlJ
tq2DvntwG/0vNXELo9Cqigzh79itjwOZ7TZvb6Kt8SVsY93VuSRGIYoFLVYhMqsIx2H5hKVZFikC
58jTZzU9DwPGNn/msYdsR0BMTN95cneUQRoufNbshREyED3r22Lfbfiv8psHlAMIM4rS41Po6w4r
4vsE9kevYUxkvLwMdMhb+wf36XlM8VZlN9ep5z86mvhPt05kbA6K55LiDeY6bPbp2z6bKFb7yIoV
B2zjPjCEsBw5skH8uFzS6rEgRLXjS2XsudyXIrOo7AMBxzF3Cw3QXYc1qDIJKKsvzzoLtgQUtMEt
Ek9HQGMijibQQunoP3LB+znfId8LDBkZX8M0jhzl50JeZV3aXQbfD0ODWfsw52n+JWjKr2nkRN2q
R+Qzjr4GO1QyD3+UH/chS0+W6PFqEfQ6uPKbVmV9LEXeytF85hr94AyLSTjGHNoYayrC/dMU0vYU
j8HXJ4ko417WThE+VDVzgGRZ6ndQnXNk0hNnmbrbsaD/GJmBiOJVgkL0VJ+aMROQ+Psal0pwPP44
bfFfcG8O+8TeGzJzw1Pk0B9V2QCavGufLSH8NfQgTo3H+oxq9w5ySoNOc+TZITKClZriRlV4EuX3
it2X5CHJ3nVMHBnL9+hXp8kHa7IcEEL9LsqhsCv0/6XDsb6YZ6LQT2B5MS7PO1A0+Tq/pJpCguuH
LKdlrlc7r9ya1bYHGwj/U3N4J6t/kYqbOZjaOv9kRRZIrjS+nnkkxt50xXZKD7eswdfibbes8qLv
U8Q8QOs1+68Xr1yf7GnyjA7kTNg2sTeIY8uZlmveKYF3pAAFfPjkAeurXT4piVdtfjZrd2xM6v+l
RV61sxWBuS+8qlHbgLymQk1NEOWskvXI/yzf0sZXHM1uizDE/kE1fA+TJJyKabCHl46qt33JiGpv
XPh9n52eclV9vZK+Y0zojEHOT9xbFagaBd0zrYfPlrPCjJk8MjpVhBmKK5w6UBZDWaplAiwALu+e
T9LD0ZGo5lHpZm/IGKTxs9oOW6X+q0ZCSItnj5DfpX6bkvV0mLfLLUFV4jGWUawhcF96XWhx3AYc
hzXr1hg59V8A61t5wsWXGXD1BxTzJtyi89d28k2yKRA4pD1/qTc8krSI7N8YwShegP0sYyETZ9u4
pILXg4q9cH12zXan4MQ+hWbzCyjkW8eoqaFcjo5RqB1S4pG0J7rpkcF4B5hEnPYY6D9q26g+mBmY
xl2GcgwRLdk+zNKNJ+TSxWV4wxqIuW+OIiyJjWciYz9I0pZmcTJnr0Q1Ezvd0vt8RiLImW94r8/I
R0KA/xQKXFfXGyH6qdJzpCVeklIaKjUSSfM70swrBB9W9Lwj3J8IDV2jOfKNio7nMXhckhYypGhI
vwniiEH5RUVgp8Nze3aAvSr5TtRJ/fb94k8r7pAQMBkXHrUpzRyrXbSjHtFFOpB1/HcwjnD5Pktk
vGCFCRNXH8X69i8CJP/m28RztSLg438XLlov8x1LL5oVohDSKzPcMSOsREXgDYKS0cKba/bYX2yo
KJLgfnK1NtNUzoD51hA2ZRasoruxZz863JW90Sv3bmReVoUqHwfhhDPQjBmAD8r95tkVJkylNmcO
Ec3NYzFz5hI3+ornUUpPe2FAacYcwKj8zY1lAx/GLE+zuzYy7o7FZWftxfb5imnQkiX+5z1OHHhO
d6lZDJNuyMNL6zQKx3D0h3WA2pS6x75wS2MjF/iBvMMq+wC+7wpffLOKahB1Vv378OCeFxWDuxXk
7wLUKTUejEMwvRACjfUcjN7XWQ1eJfLeI1H4xzO+KNqiBEIehtY0G5zWEI8LqLwJUTSjhlaaa3qm
7fndV4zVGgrQFDP0iQHKb4JIsZ54sr6CKA/BARPV9yJsfoQUF6HFQzRm96AHDh+QZUaJK+0SOgh8
64CMCnutHrHP27I4qT3qzuKFRGmAAX5Bnnc9CLzwJOA+Fg6AJ8GJX19SkRrQ6xbWiXD0FF0roDOo
QBrPQF38DfYwQo03TzF6N3UXaFW0EMUFosOCdewlcqI822I6nvLw6QhjZ0SnfwHheI7sXW+3hplE
NIgMvnq9sylorFc6PIK+uLPMh9npOjToCgWEA52cU/G5AMnF264BI+ubREMoSVIT/2Jh2yXeBCRc
DJlXCxI0FuTYYKze0NpDsyO9u17Dl3aMvkarDG4FqdpuI7PHO9cUYR1Pc335PpmRGKIHozIeXq32
gLUt0J2/Iljw0j27cVxWpakisV2czcn6WVMtrmRnKnvWnqt42erm7UzR/LxRGJeI572ZeGrTciYt
zOW+bIWlVUgwyt10paJ0xBVcwV5IFt4pCYPBf09CabxiNjx2ouT9yOqQiKHl+RFiWHDHyPcVHQH+
teBB0IqpANltcJbf0FdSkRDQej3fc8bJDwx5QZ9PseQlQCRts+oV5/HIOtB/74VkYD8LOviGmNI1
jo5T9KjnK+NpuZ7eu/8GQqrq1DCMhPL4FdeuP1ssQMK1SYjBld3xd4kEy3kDhUleaR54Nec9eeth
JK5omT0cM+fDSPzhidbS4pPMhRUaO8X4XDO//k+m3pg9HD3q4niTGJfILmHytWrNeAkVtwb/onhZ
0Ff8hMR3lc6zfQVnq/2IJi0zeCgyvXnD260/MUg5ypQ8NicPbCySe7sAsWpNprRopg6g/pW0e10K
yRmWWz0E/GZg9vxrBuD0Uv8Eg6FIsJUiK27uBx8oP82RUG9rq4K/cEjz8o+pvuEnpE8EAUrIu+Ix
TjnrtciL8eVpXtttssMbY9DSy3R4FRUSXRiZpHvJ9xmG/UkbTTHTorlK1fSrqinqn4tvGX0gfQ2i
aGwtxmVRBnux2a2jTuaBGkdLwlxYVTZaxAcPtV/G9AewAdWWNSwV85RH2Lelin9LnylED+se3qjW
84IDSJEcGwZBLaAD6Z8WGywUsYEWCPeObkAfIZcnVbGCSY4qVUDx+x/fHXewlEepQZH0Ro9/3R42
51waVNTXPMRWTFfTA8vbjUIA+ROHgWDS6CAnQoKtXnuRPPT6AkW7IYfTgRV0FdH8wgNv+Qyz35Ms
mfPexdj7+WvCgwHYZ+/B92JOFDpAMsFcdVa6WLSa2oWnxesyI36sDRftvPXurONrOPhfdIiW1xgj
Or9Mdnj5n17rkVy/QJ8Vn0dPFIte3DSeOXy3AmwUmtqxL8v2ChpoS0f/m80vXe6lSGuSnxQYEhns
5Jn9CMbacHDMOSMlk2IB0U9L9lJr+cRmVr30dkcOSuZbk0yBgF7yzsPQw6g7vPuIROqVtVig1pVC
6kR7C4maxKjUZ6I774yq3xHRsOAD8YaI+GWtUaXIh2m64VM17py5qrHZ4xafKxA7ncHbHJDuLlp2
yZ0xcKdVGY3vjm6pJp0AlB1Br+zu0ivWj9JfB1Fagd58z/j/HJ/bEQguEKmP/XC7y0CXkz4y8Y6x
wHFl0RgC/EMzV/8j1IwJJ1lTJLy1sv/0fR8/4YDoGzy/meXFbJ3IEhjHfHMmtJA3uYGdIYAhYyCm
tv9e0XjYsG7TJJ7Q0H92OMSAcPjjHwLDd6J3d8/0me+6b/HRmXpBZkLjhupo5SZBdJPVNNAmwzgZ
bxhBoL2NtkLjvDmse7vBWkWsecWs3KJLnY/fsJwYEYjsplnQBv4XgvnrsR48DGsNBLjSvxIGVu3X
wuoa7YXHDo1zrIMPVzPGOj08cSSPEueXsY4Y5vJBU1GwredFPKZGs7zkEbHKoOgeVwaNuo1wafy/
c7Zwi/Zp9dlNGN2sGYLFO3Fg8lE5q4xiMvav9CHoFkmybcYgPc0LH53S5DQQbAyfcC0291gLVuHD
tp+/rhSrsOhlQH/ewiM+nJyCKU8e55LQ6yP6yp7UrqwJUbYJBIJGVtTV+ZSd9b+X2mvdg9Fumonm
F+fuXJ17JjriWbF7umQGbV4xkXfYc2k58B9P6V/8zAD3p8AmFRzhmtJwAi+ifAvFErPmFGXcj5CH
PcSINTeJxo0rNUCc8PGizBstYW3HyY/9HMXCNVgqZIXlYbqOiCX2q32V+2y0cu1la1sdqo8+x2y7
FGmK4EEyRx8ZWf20XhJE81HhDJuY3FUxnAm1NzNP1KRO3wdk/LRPwdi+7PM7EM93nuHW5hPZEamt
4wb5v73FMJqcK4hHN3rQhmEKeU4XG/CJ9DrdDGqMU0qtV3I/OjpbDkkHcomKbUjHXCEU/V2OnlEl
61GW/mrZb4AmiSJT7gCkR+d0d3OGYFG8bNADn+QPdrYt/azx0nULc5O8UDnSd7BD0bbXmCq72XuL
DSTpQ/sgoSYXkKKejk9p9tmADu9tEwocepex3zrcofexpjrx/Som7/n3JCW89kYfwAIqYACdGgUe
m83cvB3zEuBNao97LtqhbjVSNXFJuRLNiojdEmN/9Xf4hdLMDBM4LCuDh6acKkkyQwOXXjm3CuZm
hfuOaVOPRLToNoh89zwDORY1L3A9CZMaXGzCoh0NJx4YB4SywkR5sVEa4RVNmM5m4rpIRAnXCUsh
9pRSZYkOMR62dZeWLaec0sniSu+gPbeSvkrzglV3/jgDHmPrD6v3exoX8AIcVJx5B63JZE/0/Wq/
eWNqijc61ucMDUbVxkW8osvuvKuNEsN4TWQuEZk0Vj+qlnuUx8UW8MZIw6+/Ln3EtB4LurFGOWD1
Y0qGRogIrMh5PENVL6iM7oHIkuwmj1+qRZZm1cTz76syHG89uGt27x0StklTbS2RFINDXcXkQ9Uq
ZAD/19dhhq4aWcWVGMsXiRhCpaBFe5eaF7STyTUN1oBwmV8EuOzVN+8gIEz0TJMkDlPNPd9JfwUT
mSivHTh8f8mZWAVLbw+Mg+ZRUEdFGonGm/ZGblebFCJ+rJBN45GWrRv1PbP3jlScDt00FDkynxIS
WQTuhDRh+9ccv1XfMPnUwrCkEiM48/oE1AufBRFYcXAynUN18pI/w/1XZDhULvC2kM3ufqXK3yZI
iEgAPXuj/3h6CR4IUA7McB9NGpNqbdjQdpqCpnOzQW3d/fecB+Y/ulv3m7aTrOsb7sRHXZlIOYaa
uRsnhtUp3gZHKlvduCi46Yn5yAK7mgq4sT4amOfdQkgWnySrNpLnLrDvXtpp4v6TE53xhW1o3fiz
BkOXdNzUFYKPkqnjrXrvzVk85B7DY7x3e0bCgs3APwWWmVvKnngtvTlg5waPLHWbkx/KTGk3h320
7m++izFed+K5ah4SSxXEVso/UZtgqD+ogVvBy9/A+Ey8BNWUzeE4kGuOLCWFg7r+ZKQdARu48Khp
XRx/va2hCANLQfZO16yxq3Lqmxn7lWLBHOezrbKRiZ7U1BvjHKzF7ErhcePaUKcWRdsss+jTrto8
z/VzN5i5Iz7iUDWhneg8FFZtDRJ2N25ugPTUgM0NLnNt61f2NqzvivlPa/yiZBkqgosL6X/liQO3
qpyALJiKMB3wmEtjN3mrTC6iYj349FagVT3alIriJFWxZZd9mdEgA4XFaWIEJoclFxcLjww0CtVR
UAyZXO8rBDdDIdoQd9MMh++vTsJy0JgEQlZYdXRrpuBIWHdy530yQuRqnQxGsOwV0eyVUs3a4wkn
6AiWEETECKba0SkG1XIC7+tv1wzpRMR/CqMq4cjVySGO7bRCUld7ZVAvzIJsKUC0znsqhPter00N
ozeJ1xuGEi8Y6bnwg6YqWclg8qa5tpxYH94Ex28ArBqOTN24csDuJbtKNFnzFPLeoOk+cRblpEdt
+8t9fZT2mvsTERU/1QSSslr5/Vi2O0VbCnknirSjJNeG3734rruWPxombinCc7yIGwYSlumv/DeY
KsbhIWHdSYr5o2hgQP4uE01yAgVnWjg+YPEOckvb5l62aDHrRibQLEn0csA9gggP/RQ8yZ0+g6lI
Qx6cmyw2Hy5640Vw01sFvrc9blHXtSD7VeAtcnFNyC8jWpNTVLJwTmi5YNSm2CpvBDclHjVfh1pT
Hz3pSHMGS0q/a9N/h+D0rj9P47DJidW2S9t7bW0UxDlriTCU2GP2B3NCSbLpoHKCFMhaIpNef3iL
Pu33zNXjOptdBFL+KOB/nJQWprvqCoFZ71Y/Ibp16eJPKh+aZwsYUYP/kZlPlCORyzyvvg+2pM+d
cyNZas34B4jiRRfTXAJxVUob9qOsgbChSLFoZ7xHajElwGo11Ebgi7uP9G8B3VTJZjO+Vu3SGahB
umkMHGX5frmeLy3grkjYwyT8JY7H7+q2vdGYIpxT3AZLTlt0k+t8nlIJ1DZwQhPCO1SIobFBPJT1
JgGxvx2E5UJ9gDQzpnEVOptWfbzZjj71JhptE2hNyiIBOpNR8wzBKvRkr+KgTPXoTvgV2rMNXHbD
DkXI+1CVb2UCpggGWInedvk50YuLP7xCqxkNXTgJ9eT8FK2NfhsfLV59XW6Q2ir/ajKaURFJGc7r
ixfHpLuHtHmK32XiviFLXc2vUH1n35QMfbDO5FjR6STiDWMbl5p92VE5FS8s6EcgHK/Hp2uiZ+ZG
b9saXZo2k35Xj9ffXa6iEAT6OpZf6cyUKyY1Rjjgk3ukHz3uecSRsvsZB9/eN9OPPHLnPOQfA4Ug
bhtQ9uB17m2tQl/VxWkqji5QMwfFWK/hWxpGyoftLk23SjZxRSpPcSxtft1eR3UpaY/8+PHjqOfM
pfEoxh1H9Hc6Xi4qhZa3w4Qa88wSD/PhA7U16L57onKI0Y83halw5o3vOFXM1PgvTfMFr/4L7QFo
qloZDDJ3+ihSPmhXTYSanAU4erLHdRgXKSkF/BPCKknZDRACG4kftDKVjYd8lOVvndQ4vyAP5O2n
oRChz4qIYzyQcRNOeugmeok0mL4jU/Xw0Xc7hzvug6VcLeTlR2lZfki4sXRIk+/28rSc1728JlHI
vyzExM+M6QmpsUzxcFyrOLK7+4AFSez7P0zQDql96O2n7+nqUiRq/CB7Yw5A1VU65N9j24UwlL+X
acljgxs7eh7c1gFv4XwnBr1pdD6Qa9ePEDDCY8G12gqLmSPhVkjQ07uGf/ZNU5u12y0DSI2ZuzOD
WuQSzpIozfINXR9h4eJ8serv2VfXuRwGcL22c+MymOKhsr1xSWoXkc6+ZFThf+yNKoSB+6AUOMuL
ITk0YFOwlssFr56+8euQE8I2+Xi8ttdKiRFcnUj4M3L1n0sEA4gXTNSmbMEbAMgSKvUrRDXQFS5t
42jY2+RfWdrKbgidy+LB749iitV7HRsrxQZfoYCYg8cnhsjUnU2PugPe6sqrpVt+obSGUhCs2Cxb
xiRg/f2dTBrBspvDK7ud+qxyJ0hvVK0Jl1ImrW4Uziw+ZTLq+JD5sJSsMG42AN4nEYLfHwM1SgIt
ySKnl/73ZGu/gHVcgFM2gVn4KpNWCv7td9bB/qcsFz2Oo/Fs3EGQHXfxn9S4jcT4GWDYeQbC6BxM
DcNjQN7HxEGOL+Gk2An82xNevjEXEV3ZekS5XDTlFoURCt8wy7kAsakakoVxoCgGi1cpfYTZ6P2X
Bhqf4XNj5ymnWWHSialxTJ9QCeQgF/wM0hHIkcB5mFKJBrf4GiNPwXEJRD0/KAy71Ova5hS3BCdK
eo2PAfTCNoxQaDoHCbTo5E2Egjrz/fcJh7ozRlixFxHW2W5ZWszHLLjRi1m4KM5c8Ig1Z6P39B00
lX7hpLZT4d1VXc1ciSo16Kl9/KF1J1e5UuYBtvV5jkG6eylleJ60wcMY8GeeCY+Efv96FoKewAsM
OhHZmroPJdVYiva67mgcEJAmzunuQ0Ii/lkX3ztD3Cc5/l5eCRwy+4RTR+bZBYrrtOAco+B0afOP
EypokJ4JegrPgaEl2emB5AqduXrIztyAdBfHzaYvck2pCB6PPD6DmTrCXecRUxOLjNbenNC1qmvG
2mNsj92YMgL4QIa0Ay34LahONAxCp4hXDVCGNtj101q8QtQg03lWXMZlNZeTIjiRY5P9iKyspEyx
AzV2RbIWoy3CN71zQc7DM7ueIz/dqnKJVO7nSLXTcxaOIalCij5lhmXKSpPgISnWzCfe736WTdVz
97PiWdMjYj+wUelMCPD7sl4mIheW4knIdd/fAo0jwyW/q983oq9m0XvCsTK6wbO5ZzirmMX6SxTE
JokrE9t8kfjwNpyE0884OPR0n9Kj1Ys6pSe6Et01kfrD6/zO8HfANAI0jT0hcA6wmDypgo/r0mUE
fMSPj+Y25gvl8nz215bVoAfoDwHr1UxrFM9SLHLwsRtZDV+nU/jnBrBHDrryyuPpxbJb1JGh4GuR
00PAL9kaJSaOlEmc28TPG73Exm6cJmDKYGbSeocE9qQ/G/PBuFIDclPL4pa3bXTh2j88NrsMZmpV
jmtRwnlro7jc2JRcAEUTsTpWaO96Zzti6w6bvxrx9Ta0au4tWSSq1gUp32fx0VC5fPXj7bRLJbmF
LpYz/k6yWWlTpWwPkp3uOquvM1QqMcRgUukmZaTbjHGRl1meMPEbW4v+WF5Ey5jTXGIQIeijIZt6
87uJHNlTt07D0NJIZ/9a8Jg7c/+DsXTsLoZVIEnTEyR3DiGOZaVqykWnAR/voPhnn/M4mCZB1dRj
Sq1kyn918u+OMUgaDgARZ+Bjyn5dY1COhxti+W617wv2gHXkdBdch9UmBSAxZnHOHnHIUXY/uV6p
rlND2d+EHb1VyTK26PQEh9/cB+fBdStAH6cq4SyMAvr+rebtav2DkAZIwSdogdA9kIRg4VPYSXi2
pobjeqTDsCN+QrFGNstviHvJRhjaLTiI0grk87BkLQjlXius3v9Wona9UcbxMLZqQ2RlEinaOlHX
h9NyiFNrS6dQZVQBYoqFaybMpjHOpNVVfOukt6S71+3yU0V3JD0OUPo7Q6ZCxqSMdUVPgWXgIdpj
xBifqYuajaecwg3lW4XO2unuN8vOveQHM79hZWgHoS7n6cgEICFgOb6C8NdLdSY93za+nlBpG4oU
OiODpBxe6+RtdXrNSMQK97gBIlP6C4Q9gE8W+PBFvhnFRFONEfFiVqfkPRERVzuj7Gc32ZLkHqGz
j8jvtE0v44/Xz8UpG1krCPxGWxlaIWf2ybGBdaqcV2Ka0rmfTknrQbMNa7NROsz/1NVLoPPJ89CL
8pbeIQE7UNw9bRDDETrndLvV0iabkQzObAbI8xuhdGSWvAxD9l/DQHSe/A6WbVy0xyOWlybX+25S
+rdpFfitZ3HoJ25NB4bIJotsh38bi/WhdlOKRQVyDZ3BwsOPM8OTn1n6UURpc4LEVoQZ3Kr817zY
y6DgOuLn+U3D3Xbt+F4rTRz2AssuPPhg896XJjAQidQ6zZg3BwyumCAp04wcagGYdHgv9qmFbc0y
pVkJnnFJu6dXiitGIPUqNgYHjWPQ2rpACtxvMnqRnUXoR3/YlassAeN1MvxDwllXHubRFamBMz2k
QlVAoGiqwiXRdC/uXfrPEQt8+R5csoSORW/fNF+IbhhYZmnmb9AQuei9ouUAXtvY9T5O5bEgz3Ib
lWmGXdttsCWaN3ZiSsuGqa858A8OoPtJ4RSN631GLrY1tcVOt7u5XdOEnAxAOjD8c2+yRWc9vbOe
mdEnXG50OSQPa7IDtOT7sG8r2C9O60kKLasGNhIJ42jX09hGDD8PkXq09k0r5bSVKmD8qaIq06Qc
1JEwqmgKnaYCwRU+LMpU001dTdh9XLO6BbI/pHxma4iFn/BQtTEnOA/jCqVoQKerHXCW7Ggz3Xbd
QTMJ1xU6ij1oMpK6o8sQo1cAbo2/4Jy8kLDIaXzkOm9OrH9Gq1Zzoa/LcX2Trsm1sG2yMj8ljB77
wV7tzKdxLUy8oudP4GsGSUIiaDITS6lZc9HONJiKNSuemvfF/N2Szfh9izvrJve7qDG0ovXNECXU
elIg0GkFw2qJbGRulCXsVx+k8mof/xgdvOO0FKFOOqSYAgBoG4MHImW1BgHTe2NyNab0FusGw1hO
bIRSKOVpzaOuo84Kb1iq00Zmes6BEQ11mMhyPH2LINTPZdkxt1/L4tLbZZBbv6NJWAqYN5RfQbGt
HGK2rgcBPrExFF1pqtm6aGJL05jqPUr6UK54KACZYB27Rmq0U4wRLDaMBaXMfH2BMpu66WcJ+mch
MnEMyNiN83ImtoDlNKidvl7mnT36nmMjMxd8OJjkiaXr4W8nGkgG54od+yG4cOZUD6bSKUZOr/Pu
6wiZsqmNI4aEmqUqDM91ehxTZuLKl7YZpd1cIak/9ErJN25WqMQakATDGWobAqtxdBZ1LCfe4zyI
LabPvXDHWwar0gPQiNs9dRwsEGZDesyerqjbgiEq14bxu/dcxfjPmEbwmAqUybldIKgW/1UER7be
SXcXuXvEMqrg8fsW9nLolk9HuUNXqtOPOJ67mXiuV+Qno1jrnra5YRYTZ0O32PMeUr/SM+6DOC52
iuPUuIbCtpzXnWPmRfcOBJ4Esxy8bd8LyI4bejgUXhQcvq0JLOMyPT1cSu+4RMzn5a7yv41BXsCe
igQG53kYy6tbxTVcvsqnYruNKgaFpcPTqISz4LPDoE3ZIS5pcU+DII8QlfAOF/Z1ALTchUhmmNHv
2uwya0yk9x4jyhPvCH9E4GpGttYk8EyqZTA3/4A1PnNlEe2z0WO/niJCHNpoEYozFyVieFdqh3tn
yZ3crNSzLVYkOqwa3y4rjpZD0UO4lPj4bN6ffak+SNt/JxS5id2I0llChrvHHP3+3XKdnhALkKGG
9X5uZAh5PYF3EAHZMBXVpJmE9pvFRTIbMdmAPcQLmoegjtsRYdZzeR4/LuUi9o2dft/FgY5XD4Po
nN2vNY2O4kLUxOZ3h9yJc0i6NrBhv/eaP8iWD2sP8UWmeQC42x5JtLosAsTpE57tu6IuEgjsPsNC
Ao+AZqkl3Rfs8FGfQzKzddOjLZAjpB3nIPq5riHScCrPrkn6tDVzoveC61FBuWPsY9+Yr0PYy2T7
ax0FJRzX7jvMBhXgArUdUivGxo+N42LFTZcSE2fIFGrE4s7Xh9Wt1xZggue4lQ9eH7VHJBW87q5N
TBJf1o+uJMu49TFCzEY5LFNYwT2rfCV2KgCp6RIwYDSbnWomPv1bRsyiasggY/9hzXG2IcMxnzSe
vmPylHNP908I1Ql4JlgXjv5CYrFjg4DdwLH3wnVsKeOG1g/3cJx9bV7Cd0fc0IZpiDxGjsjP/gWm
z5D4y8deRcR3C+Cvt4OXNbikMCRoTRWgQLN9vJEORA4tSSh9/nA5lSJJhsHl4QMC/kho36LmyCet
pSrmkwhKMnzle9XHKQSturawZcDWnNoeGmaMYyrQ02wjRh9n0XtZ+Y0UJ0/8XElDr5Bt4qqTi60u
/JSQwjY5Pxwzp5t1h3MfD9jgEma5MdUQ4M0eZHB6v8kOC1EEAceRlVyJVaZ1UM9grX0WlibEc5qY
+q5C/EYcDVXEwjRJnnooOy7hJ3FaK93pRMJzKRHgRbrit7HvdQENs6MEHnMTSYlSmXhB/iHyPzTu
WURNZW7zqxG497BCQ3vviernDnS0NjgKuiMaxzE7KR65oLGPQpkSrrbQpzrgfGQ4jvuBbI0ixTYw
/oX26ipDNKjjuiaCQUr8wtQQJeb9Kk3rdx7HfAI+07ON835c5lzvVnK/PoB5lzTxlTtKFzuIYhM/
7qQR89SNQkrV1Hhm1KsMlhxg42I3VHp+arSu2oAi/UzihJpPWHVCf8Zeuu6qu92j0ElvKHyhyknI
9j7gTCuE9cFF3i7Eo8tGyjP5BmyqDC4AT0VtpwvIWipHoQ2eBuiLdnGFQ30aGQ2udUimAwXoXh4j
O5WdDAf/uG3LcR7f9HuH+0t2DumFld3FtApQMqIKHg31tFv5906i0GufeGKXlwS3knscGY9dQyWi
4dSxgI0q2OegoX4uk0+xcx8Qb3zRAxnrszYs9AhX0ZZhC3FSxh1hK+nHyGvvYaDvK1z/LjvLYFoQ
VbylI8drWk3tk87Fj6hIr0ucYIgOr4kSILNfd2jniFw0oSex2n7JU9mEaA4fXtVQwkYJNBO+Uv30
yf4DPCTfF3+5HHkDdsx6+x+HVOqrxWLsRbO3kwNpo+R7+35K/ZCplp97uvjBO8ROjOowNs8CDF+x
SE5jSRy6XPiJyRFGdSlUhAjATTt5v3V1kLhypouhVW7hLvRqT70ujTYeUZjvNQkbA0E7tCQBFNZF
IPEWk1nWOo6kTmhx2PrinIGI03DvOOeRCiyH+5fVQBoOofMlCVu/kJ3/sbX3MhlWrE/Bp8HWle42
xTysuF2luhwWWOVwJAU2AGWLMyyM3Qkwoew71QuXfg/gO7/ESebPRZ0BbRZkMk4c3mqTbUAnrfCc
Q1GWTCOLGJNqP5PlVm2UVmMGnsZ5bTFXFSZPbUIsBqr5jA9u0GKfQXb1hswXnCoUlbzQ1PzpIt9Y
JOT5iubtkNXkSTytEbGIIP8fPfuWLDVlmGNYIBMSn7XR6Ve5yYJX1HmLCzebIOSh2F3ykghp8XQP
n4Pe5jw0QCWzJ8EvUZ3tgvRqOhX2v/L0Q0XoUB+jX+9HOFE6JGywm7rvURqMNIevi6r0Unz0K/4B
1ws4kJJXrduq/ynFj/xdvJ+cATAf9kB88xidqMh6o2TIrO3TqSWSxyObzYCwSbZnyPMkRFPdzC79
x62v0Gt1egJFw2T6DhKaPO9/yVebGOF6Kn4OlbSKhsLutVfFiPBZnJQfwolvCh2t7uT1oDIzw4f3
X2kQMfJoLyCKPByYShl7JRm7GzXTcW64X7HB5jrmnge8wVv1/RyvGMnvAOabpWgIj2t1ABdlVJPD
F/BIoh84YYHObB715+Q7apACERzysfYe5llpfByTruBgAEv44St7zhfzJSpEh4Fx9XLRnKWfP+a3
SmWc/n/extQwcuOMmMRyxqKBbkb47VEQmr8IrtIA4mU3CfsFemLN4u36ktljk/Z4tMt2w2bmsyBd
llzCfTKYim3Ps2XjNCsDu3h7xsX/LjvCjaKFD39/Y6vJPPLpzVahCK1Z05iCbpRTRPQ4ISBjS7Vk
IObOCMJegyVGGZJ9imoxU3wK+CkuSp87GVBHzPUdH8T4nruQDnHK147Y0hdhsBks1t4r6afGZh1+
V5TQD7PPtX+Srljf6PBByp3cnRKWv2hJodn7zuTOAsyYNzcE7m8m1awWgiVhs9TCNo6WsA04c+7c
lVMzPqP0Rgu/OIgpVr8srZL2B2eWCnioGKznu/9CYrIPz0jbWgcB5Z7elMpaKt6J9pLhWoYrEo5J
iaJjGnVD8pgm67ogPiSaI/eKYuHHCFn4dPaPOgUyyAlEJGIzQllU7qGcf12qM9ef2mwjtc4CmhqD
vw15Jwc0929Hf8ZGML/sdmqh4QJYe98oqEpC7TKsvcwXt9jewdvRLU9xPq66YYyytdhg6WXLNHRl
bX8cGuALVeMzTefkBYCt9Hq8OO2OvvCBqiFpdrRFni0wZ3xEEHh3hCW8ZlGY7cDaKTw0w8GmTm0g
zo28e7CcHW8i97W8o1blpkvrWPxau9TX4nUgM/ks88YcNKdHhzQEhX7C6xqXdGQuytUh6vsk6T5S
Om50zA7N3+JE03MxudRPA6asAGNXtkD6vDSmWGxYgOj2B3slW48JzkRFRfrc+FC1EqN+2Wf6ic1l
yc0LZavYekemoRQJ+xZ7Qs82N4TNWOOdJ6UYkrJLjuuKetFQNfFNDuRsjGWCmnqD3DH/kIPunS/G
+cvQqGHb25eVx6Dss4vaYrc2pZL1x+snn2aOJovfhG3dj1L1wp80MDxXmzCbdJRO7idmFcRKO4n2
oZqZEFlq7asvKpO8hLd4w1iAPOMJ826HscQ9a8HDPsJg6VSVMJtOgKr+RPBGKmNd6vCJtlMHWvoQ
hW0R3fJqUnI3NVRQYmlPRkdTCg87u4D8QQSWBRUGAjdW+K0+QOwqa5vMsD9R8clJXBTUeqhl0+LK
gKzsdQeTOw2l/i1N93KSUEVy2jH+WUKYrT1RuJoHB65DHJMK9MnFqsxIVR313b4+Uo7afiWyjlg9
c/P0H1Hftc4eaf0B+MdgOyZRDYgML/xgyoMRfbeAxs+SfdRiGgL0IByAwlKfDOeIeJFoxhOwKH6y
0xFe/oN8odKKOL7ckpWKIQx2sLIcIaiZKrDMw0lcyTt05BQJzajR6Wo74lebltp8JPPNFXK/rpAk
HjbfN58P0M+NUud9VUq8TUuSktHQXnJvx9Lh2hoccoZD08uJ5rUEQmg9aYtasVNbUcaKvl3CY7xo
TY6uXSk3i/34dMwEomIXrcocE3QdOqxXfnqBtQbzSf9ki6DiwkOz8Im5XD+bOpfa0jnEjS9y6FX1
3MtXOhrG3SM6e60PKy5Oe+d6TgGrKMdS0C035oSgpFtv1zyYG3aeAjMZxoj7mWoghTVRFnPtivtc
V61kW4RbyBWOLdEtvrTr9F/pQhfiaCiwChX8hSepe2CKMPblPGkOgpI/JPhCq1wl15PyRSthMewn
8djLD24fP/8Sal51C1DS6tEqKHbouxcXYjs+Th0FhK1KufvUBn7n6JM3BEdJ9eKQYuz7osXDN5GB
uicmVJKNnnIUvMYaWnLY/yQLG+kkcXDIrVQBQ1QzKyTtZLnWExu1asxzkFG0zy/5tsV2LrIdJZEE
bbDoftHNp2JmC44DAybYZmA39ElsIXgmODmoGP+uWYBANalkkTbBWtIXevVK1ACTieuRUe8pNOtn
B9DygZLCRoficab81Vx+ukXwd4eE25rYi09OJmomgEoQufrJyvXB4Tr/yUQocwnfB6T6E1NuRv3z
We9mOXfRjGKJQeuOtLJyDeqGWz0KWn5CugQ9DwxpVc/NctdWMdS+cMIJST7MEeTHxwOxeysFfqAn
8wrqN4Qf8zPIufkzFn4A8V6oMzoT9BUsjuXzuCeYIHDdvXcYJgzhBvNolOpDMzMr2MfDI2G7M3JW
afcvHFTDuOIQN8CEPw2i4odf6ozkYASScwY+JyaaJUhb5l+fb65x3JEaFplUAMAZupUmF9kMDWGf
7VfCE7nfa2ZxxnDPfzcu7XZScyIEHHdNAQUInhwKgtmrxDvggUreZHYieY7HRUF9srO1rT5AKnHD
V6uMmXZVKG+BbPnVExoZrMNx8gVyBvYxnroZkECBQIwcOpVtqfdScl4unHeD/5+rGDYy6BuAJarX
KsY8sSgUK+wb2Od81qjZwlfbKJSQW+BR5VE5h5m4++FJuozI42MJNXptt72Pe1VsPgh5uSxBS5pr
LRaITCSpPzqt7JLO/D5ra0S8d3QABnG8fyrjaKgY3TLM6W0xZsW3JlrEcoTSTOxJB63NUy6XtbPu
vxeOWQGDSUcPWpboPQN9hE8XSwYr9qdyjotzNw6qUwmHu8EC04sc1Q119y+qnXbPU1ddzLYrKzGc
sYlvo1wcPEWIXIIfvlDfcZwyCPOUbOB49oGxm0eNzm8tJx7cjIZ9j8xbnf2v9KGa9+iP0uwY/Cy1
wk8JX27zMLdae8C+jgCDOsccswoKgst5J4JrKxwYkzPfNItEVF0C0sUj/vRaxZ4JtQxz18UUC9Ij
+2pBLnhi+QAKbJrx/UDWC7lG9Z0Ys9MPudzltPeHQmkg6k/O5jEe/KNfdOXlNljGLtlr5LebZ7iL
isIcwlCF549XGGBCYaT3/Mq2OkJWNs5CwnW6dv1pwGsh9edzTynEbq2GrBBVG577iZ3lIMu9o+Fn
DoCtWqZ4ME4qtmIAZbqsTaF3GYLQ2ggO5H8E4M346PepMnjKuFINqVUSVIJMzFp6FnfrC2k0XIjp
c1xTCA7zW1s4vs9XhOBZ8zfXLlcpeHjZ/azeaUfYxWVdqK5MdwDH/MUEWgtitZSJ1ALvhyzeQxLR
11eYOP7RfxvV4kiCiuJdloscjwpcqJcDgxiXfwKjB01PHfdRNgz5td3IO1wi82buxGxUeQlDzQG7
cMBE4jQiHV2rmiWMZkuZxZr8mS6B0BfiPhD+9IE4wAJcZvMzR8tJiGAbj7ocNG8G1qme6fka1AMK
IX26Zjn5COuoqsaf1nDg7WK4woZsU67ofHqgjkS0r1WIuGA5yeIYrrG3MbrHTuhK0nPi1dp9Oq6J
RhogA39c7a3jo6iZ+v1jPFmFPKzI/J+ITMk0ecRpDRDDbyd5/brQ/h4M58spiltEnwweMUqqvOIM
0NzKJJtq2blc7lI0Ic7zaiCCTdP1N8s2u+fwOPeKEQia3bGOUMFkoFE29SKgwS1EnukYqf6x58zU
O4QRpU3Yyi7IWAgNn69flRAL4xwSVl0H66UvSGnQixhhg3ZyuLOpqSqy/EdQO/ticFerNaGTAfWU
LtkqmvtO5O6Mi+HYMlcDHLx4EUe0Nf+jiSSu61G4whRi1mMYC/f8crST5d66j2mYC4tr95l3vR4P
f5sPN3QOvpADbT4hqqbhcNKOZHmbtm23ORtGnOCG5fqu+TKqUtc9ckHMyQPKnrTHmScvz5ds3pEJ
SZqoF407iWxTkRE2033jHk/8o3/CGtV3CV9Dw2f1nnIOWAYsbzbb3wFYC3oxEAVgxXKnvk5TG9EL
AZhpSO3FJ+m8LBT6fAPZxhZwBuWRxQVrpQ7Hz5ovyZzgwIPc6dDbmOmeYhkbJ9KB9qXQuxhcBkRv
QSmm8QteYIgNl+pwlTbkegMnnsL6sBxm4LFBu8EcfkLqdZPN/pPRcfstOeGmSCzLp3fhGp4IfYjQ
I0UJY/TwaU6FgQEjQHwzRPMnmfjAp/Jguxj45a4DN2m9FM+y0cAY0xo5TI51XgbElBUdkarLp3Ke
yTVIXqr/n1TOhv3OEwqwTWHDBdx2XdX22qwOkahiFuTUtOhEtNNFg5gK92zuw/D90UumsXv61RS2
5VgMDVrnPdOEgIg/+ME/XNKfW71pMHZ7aDG6p47NqsXq+vW02vKdgz2mmsFFF8wNrAIfKhMzzThL
FwrSaKE4hIYSLgGo7B5E4PGdh14fOLl+0HOBgSau3siKtWnsUuxVewjntTQ4UmySTrbohMERn5cv
6oDwwxOQUakbFlMF/ea5AUZp63Q+BfsCIigbQxWYZpCLEVe/rOFbZmaR+k0PocHy1FxAnngXGewz
GDKYrKVX5YaI7/V9EwYcaE2fMuHeglnO3hWoa5dG0drReQ+5g9EuHWIwwh+Vf4O6cs+5/J9OmjHY
tSCRUCowcGimRXiyxtLtLxmXlKm/z9Va682ctBEjrIDK+lmMsmDHIOMBTHJXqBa+3X4gB/mXBJ1J
fdJYTeoBmypzmvYFdeXNh7gFP4Xd+fbETtt+rl+tdMxuwnAjkcsox6L5l2/NMwxobQ4KNXjmS16n
v4w27IScmb2/xQVuxwxCZER94MBFdphz5J80R+nv6N5oBqtnGNTWqdB3MhKFJryd2dcGI5xCPkzg
Jq40SVUSOqC/LzHdAPTE3Whc69dzymZuS2xBcA/FA6awn/EJ/v4I9HySytyYYxOQkeZXtbf1D5X0
1RNOAGmA3rbyEeORrNCYmv6dv1vJeBeO3qNagLlacOAZ6ICqmRGo1G/vRSS7tONimmCFFLOD1wd2
T8P/aWM7+rdmgEJ2RxSfAczihlB4ZSm1EYMBFqZOg3nUhNN5mC+HGKcjPrUCI4yaPn4EPwC5nOHn
Ks4JUuQbcKdxSlFgdojNUzDNBYZsfIGSykk+8ix8tag8JwS5YhJ2M7f8uc5lKyUk5QbO/sOotE8j
BW9ujRGy65DtK8p15kWHsgZ1tgYadmdzR2/hfjRgshHxkay3TtNQLJmP8TCn+SCHO9FGl22xRznS
T70Qb6yVKIvMwINzqw3EDVZf166KNlBU1o7dXwHI67ZQDJRPeqkF+EtMQV2nIGabRvEbLs2I9LkT
u3bi4zOvkmBzh6p7Hb2wSO0B60qhMuWCUP6POP816+AoeJ6W+WQ9OIRTY/yuXKv105FSd+yBztNR
4cc9i7N+MgYtAMqVtkrSB9JKZdymnWQSkUNJDZbhRN54bt7Zdgc/PCUzkZE+ruiLmvak9RhtHizQ
1rBhjgfwdAWQdvXi+YN8w78nlUjstIQxPqoFplB8IagdUARWn55bIQI3F/ndZ5XSpIYAjQq+sQQA
y4OiAw3oyV5ZS68wI0V9k7ECLmYmxKJEM71xLwrd55XMdzvHCfyH1eZBV9VyvdLBYH+abCHExBo+
miUZUUmJE5ifaqqlUqwcajRNyY7Ys0XEPL4F/86Xy3nfPsxfuQ80Z47K7rkgGL/CZgTr6BBtpT4n
FxyGMdS++Y5+/O6jxrQ77Xyphis6u+fqAArY6uHqrOzuUhb2kyylExqooCJt6mkDcK888kM8hwBS
AzuXWIhq4ZhWdHqLMtLCMeAkVVKstWmJsHy9qt8xMl+SfD+gGsBiKDJu3oU81rKaZjvhTyBqjCX4
ruShlAZWkxAUE8aETVskYGjhYzOdeHQTAty2XGzdEkKrkirTCbXwqfYUh5HTI/cDhOg26PZqo2JJ
vIvVpXNRFKh4oLI7l5ahz8NvQSQj1ccLi5HZJJOF1x4Wcdg5mPxjvttyVU4j8+B6mMct6y/F1evY
ETrlfXOy7jA31268z9ejuneQq7ckwSb0hkxiJ8F6kKn91tz+K8JbJ3HuaUb1wut2MYQbJKQ9zV16
3y2C2k9TJO9vZRtxS5nbkeOZxgxnHT3QsuxPfqUIk5zA0kMkqGiN9Pp1FPY5/KKKJ5XfpB3TsYWk
HPNdtEy9o23KfNsbMcEG5lVHvKSKWKLjY6I1iP/WIdiaDWYCz4TJiH0nFj9LX4TnuYTD7PPwyzsb
AIoi4ISufiIB1uqX1sjDb0pWQyAkzhxDTGZdg00XpEnuH11bQ/00/YyJHp2zWO+1+msOgCQwNREM
0t5nro0Z9R2URloWknHFsSpjuc0/TMkDjPuElgBQstFL
`protect end_protected

