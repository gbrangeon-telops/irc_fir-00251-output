

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qCd+mYB+5ZYTiHGVPy4TJGVU+1xhFKOwciEzku8LKPbRfJOghBFppfv5cFbq1oB+i1BSYIHhjBHe
eBlHNZ1Z7Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U42W2uzowOkwk+UQGZB3li5Wu+ZZMdyVhWtZ56tkrk6iW89qDlhJBbms676mTh2iLt20rMAIN2QI
nrgBsluV4yEsobcfFOejzkUO7m425YrH0cSwookeI2lEA6QsTIAcBHaB/5shcOjOwrXurevqKKI1
D75XL20Mu1iceA3triU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Nn+1VEi9KmQsJsZi+aKtcGLlFmSquXhfukwVLZNoicIm0aMjF4ddZCMvsg6rFcVwB/qfiEbWhQta
pSDRK+xrjxFlcTBesAmRjUBiW3/wICtAFebLqkLpSTW2uzkYDkrpfNE5IjiANv3SGir2AFafH3k0
HfjDFe0WiziIlRflhOF0bV/y0LPPvcdBpjP9raAJY0w7hoeg+e9PIbHp/PMxlJRxsOwGTLR7XK0o
em6r0lXpVib2l0JQy4vnsZ8th3GiX0bt/UuR0caCktJupeOBsRztdB3gkPhiKQLg0696Wa/3XX9l
8h+H5UXqQy9EN5D0ZK0mIS8tAdwDRw6O0hbAiA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2LRSSTguNLx2WvUvcdH5BTmA+6dHxBZj3mWZxmBysCd90ElOkYpPTP1RgJPbqjpN9tofDDFDarkq
+qbG4SV9hnaX8iB79Zk1+LwdXefyq97462WHnxaG3I/Bff3hJd5X0rJVBnbVgHIqHzt/V8g0jC8o
7m7eoWRXpC5NpNek3W8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MM8YGg7IvNumb+k802doh47T9OSqo/qSgWEpWTgYva1SqSP4phIChk0ewsR6o7XTxZAD05syyzDH
Qfzl5t+Blxw1Jl5F2WrihR2G4uVbXDgvFSouhPopV4gzzwlFtcYs8jnovuVf94AiRDosYHN8WPZW
68LlNRF7Ti2drGO+AuUCHhYE6L1qXzzHwb4c9QJYmemT5/44a67UOyG5CnTiIpfQTpVHSTGdVMr6
z6vPgkB/8JeX7+R+UD1AQWqiV2w63od+aHRP7gt7KRL+kgJ6qCMGiaLr3Wj2C9mfPy61ebJocomY
5wy3s56g63xqQQnm665jsZbjTUelVxQyQI2r1g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9984)
`protect data_block
zkgqmTcuglyUAPdTUZCnsCuJYLMJ91nnjO4A0aYSh5Q8PP7Iy7NQBpxSIonWRTGPgm7gVTOJ5xAh
2+sJZFrdeKD1WLILMUTljzXPtcLhSAjfsWEgRaRHldV7yjPumR4WjmeR1xfJsdKTyN0KYUuHzWoQ
QgbdSH7DRarVGfVShaRjZIPUUNrPXUK72fUuHpK8PG5IqNCZ7rnatmH8a0vnl4rAWiTrVVst+g4K
5L8N4ak74y4Xsthl/Okh+xrbFgw/TDb2znDrYjhMfXmRfFnroTLSObiqLtivD0VsNwrcSGokRFuD
pExnwQMEa8digE4jYXos1eg0OZCPMUba+EL+Hd4WEkPaYvWGo5xoreuA68VDtDOgPyzEwpn/qivN
qpMVNVdIffKe8wxmk0672huR8ArlaY/eXXbQ97jY0ST2EHKh6arsMSifALq05cBAVTqJYEbBikgm
roVAAcmqNyBAePTgEZ8OyFwX+VSntnhZcMH5UmlQ+K04qPc1o6Ce0LHsejIA7pJtLzoVdo05lAK+
nJlps7jMcWEoDNPV/lLGWp9F22fuSUXxGg109m+p8Vm5d/HQ2iFonlMYZg4izNsdbws/DJTaefzf
oJDCEPux3EoUKx77mMt3VZbgDaDnKmPDhlw8nlNFsjST2dmNr1TF5GI9XKk6FXUc3f7jlCzcdnqe
1QO1xix50Siv71Q1aJFE38TtmAvAOqt6RhWu4PdGrF3Op9vRmIn45BReOllxFN3C5c3OVujZG4Cf
JX4gNOoL32cn3fcnpfseIP87zwV63tiYHTDZQ2HMjbce9cMOTjGJKkdRJIMG4uOOUo4CK1zGN3Ej
2mga7lu45K5uDzN0ZM8WSUTq7T6s6gCDUOuzOwey0pb8OsjoMc5WqITfVCJ3oNfiPh4+Li2LpLRI
+QJ4CiRzghWwZySUl/EpiSuOMKGaaZtjhYMDhw7Hp6dwh96RG4yhCOAoEgkIIbkFYsKTlrK42Gxv
Zb22X1znRPy3/1rSizqGLWagKy31OfUiV1zjNhFdQ1flxEcAzpVtzY/GExQx1lesmZxH+Ob/pDwH
9K04FegeX0RMzD0I2D41CU/PdH246CBcydSMtmEtnRpUiAAUn3NTsYgtI9A6YU+ec0YewyM4Dsf5
YGbhBonlGXmRKsdUk34fEKVemkkc9vcZXURQghZa2zqy0y+7nYgbNBLanAoOol8C4/WFz7iEXrdQ
m1gKExL3Qzqgbv8WCIl5LnkZsCgJRHfWQz1TIYnnYBW1PDDL0SIXle0+l8mfBeJYrub8+QF/P6Dc
4GeU3ldTg58gHhzasXU924LqN8iMLAQzuqFpMY/tsewZtRe/ODDbneq1C+fLxdOX3SmzpluWlAmt
eYW2nH6m8Lxhbsiu/2z8R4dsnpXqT6/pinbShtK9jITroN5wJm5Y7+ngIFmT/8w2Wmk+wcmfKuQx
CKiN+2sK26us+EJxHtJLaabSy+HxoNvJPGESdotpmpVCbo96GglD6ZvDSMVLk2APlzZWMYdSqpYO
VpFVkF8RuEiQt6LTFTFq93UFlJVKrFsGHRIapbTt7V5FSKiBlGJvW7Te1RiFvPBZ3vlxSsKkNce0
Wn8V8wnXwi2Vu8cWmuXKLF5oSu+Q0Ugue7E9bjAqywNTT8377pxFypAG1XDcJkSIrOvKuD8j4YLY
ieTjLn/Q+Bc6NXUVRbIn+8UcOJku772f6fM487t0XKgDBUODgzSgag9d1D1PbXSUNiySNTFsOL54
4jce3WyN7ax/g6nvEWJFyrYMmPmj5A4fj/RAgP1aV3CufuxPjGRPmxcMWO0uqeE0vKb/T48t1Fiz
QWNXSCdm4uOKUeh603tekpSrDucaPGCiAEf8u/lu7VfyJ/BS3PZfZ2wHfaI6KcTQCX+2OEr+YS3d
6hW0Hzx6FGbQycLs1Gq1ICPWDtnhleKlLMAT4MUHeLSElOXNAzaxMZ1cjma4oMqdMAEf7izmmAO4
G6B0Y6xg7Khn+eUjC5t0g2h10CwJJVf5j8TaTNeHnG4YEvtQoo5T8M7pZccNswlplyBk2/x8xwqa
MqnIZyaKOQ90T5rIpAMivkA3L4mI/OOu2i40EATS++A3LZGNvbiTN8y240hchoyULcn+pmsWWSn2
ydWIq/jAsuU8KVEzoTJpEIJ8hTj+1k3wCfsGFXJVAlB3bvdFHohYPW4lBF84x1LsOnzgPVa+hggF
2q9pMgBIQTmYbEcmTxB3vwln0IKwBhADut3ZYptrtetLJNC/Ce7/5CL4LQN7l2dzh3friJ5TE1rh
XP4V/bongTveb5QPNOmDWhVB+KiPOXff0T4sTdvsC5lba7zYtYuTJykyR3pI0WQGcLXNHSwQcsYG
ajkYkiMD89ekAxCnj9iesZgBmTKMW7DBc7DkNY6dbNTmZ1AOLYmiDCUwoPLOM+XluXbtdRZv98ii
iUwr1G71NwFy/8uL6vOKfEr8Qn07nZC9mEwhuxEz0EREqiQlfH+2O3h9VxxQA3kpdkk2mOHErkB5
e4qppvZtqTnJez69GMiBNlndecnfqgBfT3/5lHcOegauQLrrzi3jzUSkvXMkzgknDgrtrDdIu78Z
XvReJY8p/0pkPQT4xyjTRTlLJdhLi0HFLRAqTItP1E2P0ZzHweAfLHs2qcpAlHA5u2Bqat8+v1EL
4j7ZkE8ngVFzEmtEpmRLi6OT/rsWtGlIvmVXJM+2ZfbIQ/btcT9vLSTVCOvcmMYVmi5Et9gXWp5l
qBsYksC2gdVGWgjKYF+ZV6lSGBVfL5IvgeBHfSZQvIKEtLFJregOEjZ9MEhcOCRhLt3Qxtp+SdhE
1MOtSgMSsVIrmUO5MRLCsf34vpRbIqMSv6Z5BkBNTU1pVKd0gTA9WdDcNu9SDHI/XQjF5Ai2uyxn
1Px0z/AZjWZgDVChvYKAzXm7CahGMZ33XARmmYPjg7BVAPcXD9j6x7Az1bo9VBVhGFPK7zgW7o1j
Oy04dgBdHrSW7GmO2Nv4s3+gl+jqz2rht5V479aKa264W/bvlOFUKFtexuvLSc1Mxlw9WRzsy8w2
F6sF4aO7g9yIs0j69IGAykDNvWlyMwUX9qMB1wxhXvK3iA5KBmMxrkazGV6SHYhX+lsfdrG0+OQN
GMjMxeuSWuHtCny4X68TTUlSmAFRc5APpH1YlSMtB537e/DKDMyngj/aQ65NYlnZmqeMtK+JVSTv
4GifLwETpyFiW5egf5MTPRnPTg0k9lVkvFWJeh5PPSjjcmRiaqn63dLf64Aa3cUX9V7e6hUzUKQB
16lUwt4C+gjIc7XuVFlOvQ/4P2oD4b+HWOcK7ns0vdgG4v/yLWyCqjxzTTWacIOJXMIosFuSxzS8
N5qxu82MMGXELxE8hepEbOvmUXDFJmwWqRQ7sHnzj9UYP/V/nHcT8ODgQ+vszCArJOUeheZKjkzl
Ur2qOkOa6ntjb2nK2qTaBWL7BR5yPqIw5Ns+JTohW3uIKOYPsfLNwnvyvFMVOa4l9hbl439qnbLp
S5Nl8n1IgncR/fwuF9N713jhPlrJoYX3ssKKBjy/iPtsTOVehPIgcI26FIcqB3Klsw8zjECvh6oA
BsktA6TU9mV2fRhxuhiGR+3wAezlhGEXe6ymZTzBvSs8iBmwvTeuvqz5zFbxGRrSe6vsJ6Z+w7L+
lcv51G5s/bVYzlF5F7NMNku9ywHztA6GTHLF9dJ40yAJrFL8HfbWFMRpUkZLq+B5R4eu/D/Zillc
XX91hskaY6WYSBq41UZQj3f/2ugunDjmLtz1yZ69L61ZOgm0EHfeP90p+TCSeiI1t/1czZ7tl1UW
0G9wzX/DA5m3jtxPoNJssCGhaGXEo+q8yulOQGc9W8hiyyUZxxRSG75pxtJzSB9oBhSYrvzNYaT/
PqXONbcz4yXmQMW//Do+qzSnms1O0eWdK55iEgdYqbIvhTCjW790U5XDTJFbzL13N0VJN7FmITUU
I7d20AUuMuBVIGyHJ7h5vXch8uIS3PxCjUgP9lB+/FwuAS6yTX2ShpZOD+oOCkm0Npxz0HWz8lwL
sxumw0ENhM0VfMJ7DfQPtAY9jk0BHRTIA2fsrhS46YoVd6WSZ9stfhOHOnrmTJ2QrrfJL6bXDsAl
7ux1wmEFOXolj7lu0owu6X0Y+yscEoQnP98BoOTJ5DLOMO8WK2EXXZItxznIdPAPjVHU2gvNzhuR
mixjtStSudZnWVA0yyRMWgdFZOuw/M2hxH5qzT6KGs8tsdZE7Yzm90vA/Gpy2XAZXk3yOx4y0UJm
pc2ESUlWMmEd+bgveZHHAVnoWr+q+TbBboAFdRSuWYWLoDD/kNNHYHI2IKdZWfYu/uGoZy59Jz6l
UK9i4PMkdjk+K416ZL8FSBiljdWtAWUWAtv3NIgTnYAtKtr2UjTqwgR4vKPfDlKi/4u1afsHGVic
EFQ7VfMdlXEWvvjrTnR5NlebLdmKuLpbOKDXyNVF91pqkVl8IkFmyKMYHb+DOtdQpUcfgHoNXJkO
9tQzyleJiBf29hU7bXQu5bEP2JyTO5XlgNQp69mcOPGOJoWaRV3i+/7C3UV5KSKSE4WZ0bUyTuN4
RcDAtMIUtxKj7GLHcZgWadXFwai1AmKE6MGEA27Gqk69oEe6FvkE0iXPhlBKZ3sDc7yiRBzphi5l
teYKAJdkCpALMcpYg6+N0PhkuKekOw9/b6hICjWbMu2APTGs455LiB5Ow0Vg7gk+ykesqmYjj0dO
+7PFP4u0rhnFI8RR1gOgSp1lvf9v/ZLjzNTAwYHxrJjAqwqobOWftnUvUj5/F2G9wD4NvfD10/VE
TgXHNSgTsV1Zw0fuT9us7oHMwsitaGK3NiNhF0gm5/eKnfGjLzbCUA/WqkgpGrxs3m7L7eCJ/BDv
TC34wSTbKbtL5eywULLyqXwzG35bq7FadcdsvX+VbWNOzgL5+MVt+pCAA2DhlS34qaNd4mh5m8y3
mRtBgB8TUeX8D4vOrJfwfanJZL9cb0WbWb0UiiABTFBJUXLNN/Ez0nXoVczA6R1joMTDUUaGCnZi
3I/tUK37FM9vhehO/rIn88Zlx+9yQsijugUgo5aOrI/dA+BChuJKHB2GcwuQI19AZUTYdErONhbI
2hguKac9Bm1b0MIxsXB/5xZLMWFDkKQ6vqj618gQIDcCnyBDVhVS89HIofOLcwWwNA0CQURuBqkw
iiY9WzHEa2xV82xId08v+8ZJLnt0Ff8WFrkTWjV8ujdk2mht5Rl59DchIhAIBse2xzvmvGWRnPGX
kpbBDLXMjov7cRGzY7CU2Kx4lNxVGm/q5nEYChuJQs1wpFnRfWOFlE3BykR4DcNlsoT9ntBYPkuE
HQdEW3hIRiNR3/Xlva6kcOC156e4cUhzQRDfjXnPPVNgd1pwk0hY5OBhNTmCskOv4NXK1z0zFbs/
kkzojWunya6usO+XX3JWfEjRloC3DWkbYbiLiGmA4h9tAV0ERwOYDnaL2RPmijH8TLeJLRlW6dGm
CCZWpzkfAJG+ESp7CjWvTyafDp6S2DvZQy7nFoAvNVy87kAjFVKG5IaBBebV6KTxcBYzpysXbym5
BWy6jGi6eBVyQV6UaXWpHxRQQrWRGSSeHlng+lPd4xGgnmIXZzFtsCvAu4/JLy+0JoPWb/rw3AKy
ZjnjsYuhOGbY2AWMu/nPpvHxDrYyzR8TYUz2655gC5fJcK2UIhUSLrKinv+PhOYOMi582FfHRjzI
Z8Q6Ey/5ypRk7DgqC/6Zmp7C13zOt/J+V1R2t0tsz6Z6nNrNdEXn9emdiTVHP71GvVUt4B2nFxFe
x4hGPf/RL9RxP8YBPAutIVJRMV+JAt2F6k8Hq33MB9uH1F1Ags8wbu8FsuUJMB9Ffp/KJTTRUMgr
3WraIo9E3Q2qFfLAQT5QvDPHsIaAiNE1uMbdy9C3J3PyTS3hrUKbWOxeTCCaXoMxA/AOl4ceQWZa
X78WexYMFQAQPS49fzSLs0rqd1+JnkEgDrABjsKJtGrpENE1SciTsej25jaANc7nicWjzDO88s6R
veEDa2H/2v/aYAR9uB7zoL1vX9JwWmwT6PcKAZPY/my0fH8ul0R26WTvqJD7mMzMytnJwohfY4WL
Rmyk6jJIjO3sIrAn9dcyMv7B7KMLOVeBOQoYU9AV4It18A7iH2DViFTM2ifzNw2k7QuHIRwwW+Tg
4LgFylTkQ/4J2ku5nmIchq0Q407G1HD/KqGysik/z5x2sXYSEB50cFJkmKx+7oCkXtr9a/hT5vc6
aHAU/yH02lzOAPOfiPNhGy362vizSJytKmuz9kp1hlIVsTCEVaMXr6C1Bb/YTiCsVBBxARQ/DOf8
6ixBJWGH2vQBd1HbWAexdluElfT8+iITWXss5m3o9W9jhFz/1mtMAWqAoOT5T6J3lbM+ea3N4eZh
RX02pWOA48CdcMw6JQR7OFeldeceIBOLoZ3oFa0FImqSwaJB3+i++CSGN0UGaT1VkbXocB9O0KT/
ds49+4dAcaCxYNMWwANzJRJL22W1rjVi6gZMuqYUM9Hsnf4y4DqrWVTKCuj6gjgISr6Ocx9SD0CO
OUzzx7QNMJSQ5dZkchJNKRHJmeQR3dkbTOzQxVnroQnoPvRd76TVduRF9QOLbIbWQcoS4hP0wX9L
em7OkDR7Q+7Ma4RFvCNNIg4cXTK2EKjrK+8sdPt3xpqPgDH6HepmVHvrifH+4dTcYxfZwzWPnyXU
BZp6KhalO6+7bNmmlPzWD5raWB+tHQHr2I4CpyusA/65MTxhQeS9VIb+d5DuYwJ3zeureY1+xovV
WS8tjNZahygrfC4xqaz3/0UqI7bP7jO4vgQNKGgBJT5jehQR4Y73omvTnkiUpYvDjU/wSm45oa41
a4Y5NGUzlmvWq9ynOPtBfIkfpqNqykQmvR8naWFyFRuXP/m9o9hqU8WP701LVPljvUR9k3jhpYsU
gsY8VIzdLA3fXpWxXMjEbRmJWxZlW2d9br4tFCxWvKeTDPphPztkWfMPOyo9B8h02YQvHNjmwZqr
XEM70leqn61SyI3Y5Xus8ubBvkVBmK/PN3w4doMg71TWTx8nKzzviQwze6/nre5oApEaDOT+laeT
lsDTjQ5JAfinbGFqWtwIopgBTtnhxyptaha1T9FSjc1SbDFzR5ELRFhYWFYjqMwU4JsTpysHHNZg
V3OR1wZLtUKOLunJ6vpROaZt7k5bLkFpTF5XQOYDzJZ61yUzGf+zCBvUHPCb+HV8Ey+TfI25haV2
gMcd2hYcVzOeMBMUNYeIX1u7tj1NDDM9fqayQzXoTthJ1I/hyZ47zy2lQrNMMi1PfTWeL4MKDpI9
tzF2/ZiN4NN6rZ8uCZOhynjNNtMeaN8hcGaKLE/gzKvZWyRG9fbNNJBW4j63Zvv3OihMsU3DbPa9
xZaPMEYm81oCPCqmfEa2ITdKUsPWPLCT3JLnSO0dI3BKDoC/di7ufFMooybfcpP6m7kvhEwmxtzJ
prdH/cJGk//R9XJ68DrSL0Rqnrmv7I4J5aF9uan6fsa2+7csSiO0U6T/h3RcOt7qQT5BmXIPMyVI
b/kF0JdSnTS6z7oUynuJHBSnDZWxJQP85SqCuJ8Kq9+O6G6aPTVrJN+GGvJOq8nvq4viudIFwrUo
HOc2bI0mveiraM4AR5NhnMCnqvKN7kQKi+uxYy3e8v19GGXqTB21UQYYlLs0L+5Pyfkw0srF/6Xu
M3VX5by6f7Of5nI4Ou1bS9eaHzsWuqO5fw1dURJKc7EsrH7fvhbhyxPeeGEgXMz4eK92tlI+qM7p
4NuIS8d+eraiaM/UCNuYtw0Ab3hRamO1TCbSGaDbb8MKsIoQtFK/+pm0HOzvs+T7/iCQ9bPMWA/h
onY70DtSdflHB3onBMkaPZ07p6T/3Bk5T3k+oKouOE0iKV2kbt6S6a7XQZztqfTjVM6c4oLyeJJH
MU/poCrdPHH2S2qtPEhTHPQpYegDvvRBVfuS2ZlE1HOPASL5yhfK7luWKCI625cIVkVOY8vALAw6
h0yg0ttMZJJFBX1h54LqINb7w4kdQoRTYZcQFLoUusXBFucuxfe9J4PY37MMmpl3+fKT/KpxbxD8
B7MGmiI55tJFz6gS/bvMKz3iRTCp3ncuYNKlBUin6+NhZOtc4ZkLlTzBTmobxTgDxuv1u78OjZMX
yWodI2GpceDsUnUwNkKzcPEDjlHDAM8MoyQKoWKNaygEvwze9NNKAYaChsV2Sfz/CNz/xn1EzxQG
NfW21aFG0dwh68e/hQhyjazhmozk/cEKAPtU0vKkgzfkPm1zP4IHn5bC0XElwhCUtseoppQ2ThK/
PGsyTwQkZb++P14gfc6N/APWHw/GHvhmdgAzbbnXaNXiHqlQ53T67Bryjd0zVpzilzNONri5tUWH
TmhtoCU65KdcKV/0oWhUhg7/0znRk5wxkYS3GjLfBsB/xN2PRLerlwyKtRnczV+IeMQRfvqUOGlG
xIuuaFlMofRFMIPKTEKinMbveaQ6ZWXbZO+K8msnCXPnN0I60EOADSDXG9RomlFpYPH7AhwoeVis
GeszljmqqDxNBzc9o8Kj5WyHJGEUn+S7G81olqFkFGbWZe2tI5dCR5d2wdXyyk8q19RcUxAByZ+t
psYxm8O3OUzO0UcSEEYefbROua86Qv4YcuqkHIW4OIq+KoKqKfJ/TWJ0cDKyii7OP/7TYhinMO0M
ojp8X3VaIO2AaITvuupqwh69i4fa5sjyoar8FngjRR9BphMA0KjyKOBDjMSDjPfJXwWMb+IuEe0S
SJZMEsF6++GddA7RDgzD1zm5XbP/z4fE3UuATT8eOFZbnQXIdjhG7sUw8HNLsHYqk57LQrhcd9nQ
5TlUSn7nBGS3eoU0aRGPlCP+y/Uyo+s0wduXhpDc3ivVjCSwYV02GdLDFFegg/L/69qQK6vs1Fmk
ACojxrARuUm1z+6/lWSHVuFqzALSpVDoA/+O+daj1eGFGPfPcBQZLpF3++cTqHth/OfMe+us6EEx
Ln/ZXTA7JqG/RSy4MOOzez5HFMMIFJw08tBHAZCTYyq7l0p3jEnfMrhzYX8DSdc/bWgkOgsWGC6W
bSrJmyZpCMl/1ZykbUWXAqbrCvo4KubiM5I3Eo9/XI6g/ORj5MUY4bgKWSyzzSsscIU5dQ4qjz1u
lkGqgflUw2Wk2SFV0CdOMfAbRQhajgYXoeL6C4S3KkJ+IGOvPGGCHGgq1Lfsu0ZcSM9Ki7N/+Ovi
9BEgGZPfbjk4D1xUiaxxMWKgIVZaq9QA4JbHOCQXXPYjbqCWgnfJdOTvWdXidIlcBVsit3yCmSTn
bzi8NOuu2iFKCSynKcojXW2C+atdE2P/ANMB5EPOYELM0tRgg3HyNMIEi8d9CrEk7neXda7mqX8l
cUdtos7ds5LW8fJ7aKATBu9aBTfRUUHhoEO/wEBcsRJtERSh0nTxdPdjIbe5X/XrcThGw5rnNf1/
hEDKinDJ17G7AdW7f/uLXkkoNuRabCPWsxg0NLPGZg1aDorb22PR6PbSbuQ8AVL8aZeb86WIgB3X
X3WBsRB/kXTwhMjnKHJCZvGqLDZITFjb2zUu+3kf1uC2zBmzAaEEE9C+nBvTwrbv4LfnNjFSrGAi
bADmkoGOZI8uknK3Qn3x8UIR+wp65w55nYic8975aQuXyirxz/fThxsz2Ro/kAilpOcCC0Zl7ZTb
bmVy1uswTjcwzdalIxB/Eq3GJBp/zcqsi6ChbfvZmgoRHpV+OWw6T6lR8Utg19ym0dbMRspRUY2s
u1uI2v7KzpOjy+G0DxHyzZLviWh4lpWD7jK2mcYzx8mvovrmM/fo4pxh6ts5f/KyWLbqbFOF59XJ
k6Nqy9MSws6Qil1qWv2nLlsQc6SMfcqVkxG0ufls/gbxzqxX24fKu4q+3/XGkNvU6WO1PNWB9Ei0
Do8YJfxKn3XXNnC6zT1c7OLrJ/q4eOwqHuedOkVHa7Omu4wzyax3PJgWc09XcJ6wOVln96bOEhJ1
Rg+EhCs7o03xBlBOegDuwCwv9LDEA/Joz0RnlaBEX+GNAmuxHxEdO30idZW+TRJXF7JvoNQeBtvA
PF4lVMtqOMEh1g9BTAgwO+E7Bb1ix5Z6VMi/OU+l3BpmG5QoxUJDv9jgWb+uYTCldCbSmQgnoOS6
uyQmfukqByWT7wmHpI/OQAyJJqbak09n8/X4G6xMiWjg1oWLis+2Jg+nFCdTYxrvSZhvAwbZW9If
IKXQkx7kNmEX6L3Nt2gKfL8hBvmZlUEPtQJi9qgQEqfiuWoCqgSEzdTfTQfQDCo5xx7wi85lB5v/
xkX0kGEYelIbAENykTsmb5fHtD1KEQME8czwxht7m6rQ2hm+W7t8q32jRLtdRiLbmdBl7DtKP0yP
bqBWAy1qUS5GPwojDgxAuNlZGs+s7qd2zrEvC/PJ2jl0IyIQ3zRkSmz58nqe8vm7XVzrUY3F9xmJ
6QZmk/HDKr016Ucvp/F3o1n7ZCpU9U8gPnwdYuGsK4TYg9fxhdR5xbhwK5EyUU+2dmnLO4YMxM3C
cVlHdINGoWaNPGuxiWu4yvfPT/ZvI2lL+EioIPaGymzR9oQsh4sVlimTEh1eB7kNqqBAqAKBXlYQ
6HCQmWxHvp14YBjUNjrQOtjjFO3eNQLwJ2uqOPjU90qg1193k0r/lvZnIjpHxw2EGp4SgQ7xdjqd
EV4Rg0m1B9MpkV/ru5gtAoyXWpzy3nXtul2wDiJuDpvf+qCskGVnFpykRsLjQHAwwyAoC94seJx+
AsYjHa3ISKz/Jvq5kvJcgumBaWL9C3LW3sHfuJh0Zc+2g7EG+lhKE+EOfz9fObO8fLrZA90xURXW
wQ0zg3Raurc7vsUcVZ8eaN0FJaR0xLxKavCqdmKHZfNAVVxsztvedjVld3h/D5s68Wk77fcmVWpz
RvT9zOYTZbCTwkZeM5u+D9EgPeYPkM/u4CFROAxSyEYSfBMh56VQysA77ALlaEgwJJJlWOEe+yCe
v9RkSgiV4TvZ6piHSV9smqTjtp/Wx/PADJVMJ+NGd0iQQO6zCaHxGOqoJuY9RQ2nSteT0zRlLiIy
KHHvVGqOsYPzb+MblFSFhrXVGpkKH7WPSMJvjzuB2PUqBWEecu9LJgjixV7kq9fFeIXSxhJmbyrq
oKfW+PzRadMeP5pCIgBJrMiD99g1/CnZpxJKFeQ/xh1Vy1OBtJQkHBAa8/PZv981P5i1+9gpsgMS
DCWUnQYv+k48NvoDlpTY2o3hnpZ5uYsef8bAkfnE/R9nKaKcwesMXJwkTWXpolq7PXrUwdZHaVH2
YCcHR9Y9TRq4qaQ0PU1AzvntP19ypjggj+SLlsCyAG2J2GZUpa1i6WAZRTfWx8/cLOIfUp7aIUGP
ZYpN6Dp5J2M9crvbiJ0tIsK0whiZlGEaIdYT+OudGT3nU8qciAi7T/OvZVFFgkpR0CX0VGmJzf+w
6q9CvgH+3hFcNH5GUV8Z+V1lQ1owM3pbaaXOAq3rII7VUYz04ZOXpz6GqS6ar1Gjg2Z/3gh1drdI
XtG/YQzyfpRMUIQu1GHp4wkxHvAhm274umhQQTb1aeNWewNObP8221VMyKcqD9Li3FPVG/Sp2mEg
x0pEJP4lM3Vq4XYQh174bVZgRdeiJlkDkS1eEurdxrivQxP9ecfNpXnmFKVHBdWoWAu6Jmx8NkAB
qsc8DBHjyNWtLbLyTQwW73KG11MpiESgPvdRXmwZ5dOkFspiGOotuhF/NvHWkxbUVZHXWCAJVLrH
8l8jn11MHkwXjiU3FXBP9iLSn4idId+XFW5xFaQdqDGgXSv0rxD70qPo6rLNslX16d8BRpRc9Y6F
ELqoAd3bLesfwmiF9sGoaiNo+RZgWGt7rvV2X3N3vgpv7L9QR2AOT0E1BrHHPYcOfn4ZHp4BL1i7
/MLvxs7Qs6c4/oRRH6cexc8GlVS8y8nvhd9pWO7EXMxNR9rHCjiak03OXecTwSkLlsA5ywrPdZsj
aufreUvELPwyQ1vNkiAsj+k1KhMIaOBtgRbv/TTtXSHdYp/pFP3lzPV7hlFBEs2EGiNAGRutVjaI
Umw0UXvRd71wHs7hZC1Cyg1uoxJVFJVNhQ1Cmju+3AR4+53TQv8tRH0s1yJF1TMDPfLrYz5/5rS0
5FUEYWLyVRw/X61CcsON1+9sxOuVctophNtAZ0y3zHAZPX/HOD9C6bsnV5bAdrzoCIYLGHD/vsGl
lyoDRRdVGTr23jExGGpRWlbzr534+hZGZ1AaFA5us3rx/FJHYaBE5GDW7ps8EVWE94SOS1QjICqU
7AFqloqvc/e0Fx9QvI+wOHV8gOFISnTjAvrXxAqxJSD1ve/d/g/NVMGG8itG0VzSS6wlI+mpf/C/
hgM39odFvz1tMxDox8fc3C+CjLhjSZL4GA3pwpMHyAuMF2yLugsVy5osTSTCv7szhHbKgf8UZ7Tp
xRvj2td7VHZTyGqMKSEwS3S8xKpnPVVgUABYy5HBTUcaFympz3jKZm6Mmh1wACeZyEDZGZhv1ALn
Zu9BrDaTrZt3iOLhCkuDgrPxrU1WMQjWk5xqm9ARQiyvyV+lvZE8KaEQ4qIES2ZfCb/1Hwq/oDAP
uz9XpMLT2/yQTmj8nWqPayay6Bjn8PIxIZkYL023aduGBekJO9vZibRSXvcmYoyzN87tvJeqoHWt
lGI/BPGSSCvB990N2GNrD7CTPXLSQxteEyF/G/8xvZ0a8AbcjjAnO7TmR1IPiYnbYSzvAJgnbGiw
fpBsXIvHVtU0oEN/DjrBSuYhHsm+lV0acZ6QmsYjOKuyPxJ6IUocQC2FTcNpXbvVeLecbSnW81V4
TZha8/NvVBHQduiACLrTJtt8aN4IKz+cHHNZ5uppph/SXyFZA5Xddx8eZzl1rgXXnr0xUly908IL
ZJxYZRhc5ARWsO5/ImmhAVZ93ubLeSxvIIInf5RyP+j7tDdOWpvkejdMKLTTQAzTh2+Htqa7L1Ox
GV4pKrAqQKzYLxAA1ic2sfkFP0cNIcPgXCZSOVuBTmQJbxP3oACoG/2kQpV7ba4U5H9SKALONxyt
/pQNflMQbu4WCrAwwSBTcf6xyi/zw3wtHN72+2sZzm7j4cRDgxPtUUeScJAVd1JYInR8ypZtn7jL
cpU1SkDiTGXrfpvqHr4CRUgL0z3oRiFikiyiMkbfcURXWCRLceIfoFglZB0CcNGltbyvLru/AE9p
+W/QqgMdp5JfvU66siStvzlG234pIA88Lus0fS3zqUV/+PJUilxeP/nvyr7FrlEhD48jr/tpKlYR
wrXRvsUqZVvyyQji7xPIirlEN0OQpNp5gda4Msj7dK+5ttkOnt/0++fr1mEchHVCAhkwkSACFcS3
TSKt+LUMiIjG
`protect end_protected

