

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CmScm1EG7+yOvSHJHM5cOhdqnLzZOcepWxY9DkMOyN4kLbgbdLuAH/l5P4gSPyg81gBN3kT+DB4u
PBXNo4263w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fwqNpFcMm3h5oYp0iLLBA7jw3Gfbtf9OYXqaNYQK5M/u6ozJ7zqm8z/7Gi9eaTLXS/9fpHpwK0LS
QxC2diEfybnFW6aKTP/iU4AM0T8Jfwg1fYYXa19VRgeHNuXnOnQbGrbwOzyL+M1AE6VgNshYAcke
HFUgdv42HBSaLBuVCGQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D3xIUFHSYN/tuU6xykyZi+w6uytCi8PG1RRIohuMCP7mdmezS82HpITZGe26wOIBAYGliyfJF+bm
//Xu42+HAg7awD4lB8/Gfse7Vws0SwmUepHhRYxtuQx+Hau6aq1uL1eE+GMEUXgxZ2vOXH0ipYrS
hLEg3TtjTbccTVimoRhbMQB8xVTXKgd1xaluMo7+0fNF3EBfFdhrX7VNbbmxpV636ALP/wC6VRmP
XNe5xXQjiv3FP3uE/Bt2VYm+z78C9QX2joRNZHnjI1wlv+JUs+OBnQx0uieg97dZpGTJDWS/ROJD
yUMDQnx8oeo5Aftp86QvBAbfaqE5X6J2q/lamw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WD1VRz/pLvBXDYk7fWsqqk9E+EKCxbcP63KaJV1ph2old7nkwo7SBQkXHtT+4KqXUeTJT6DxPa8j
tS5RCAcDnWldx37xHa9SUujjT7DruuKAJejsjhxtSfv6A/nEW4C6nOkCH10rAuqtBTv7SUZEElTR
EXiyr/yJfBZig+juuEc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TO3nxTWXykAydBE8oLE1lWHpTk01Db/e9HeGVQPfEOiTpRxWensjccZLTO1P6wLTocrobkWdnzeG
BxBt7prIiPwnDDfhHMe/xea/ckp4CqeBr0GVOckjbocHEF60X3dEzewbdNfFWYT0uATcWRkKB+5o
X3VNEsL1+rzFW3yXd3oxwxLZl2hrAEzHGv2AAZZgDP43u0eLOoQsuloFBUh5XzvTCc38IZkfTB7l
fBrAnLiMxoJyYNeps3ny9evx3MIX3RbK+6dmn9Aviq++SNxcoN8Y4/1btHsL6F9ez079jTeANSEU
ZvBBfKlGq2n/FXU3NGHAnGxirPn//Y4kyfC2Kg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10960)
`protect data_block
PXUAA5YJ142WeCdhxOe/r5h9K6xL7VTkniRywlNLwlFCCBqD1qEiEL57mFjc9jQVZXLGj01lAxI6
5F/lNgFb01q4gXYdqVawWFZ74g14wnBzF+b7/q6m6pEuoByIGItBFhnCtXFQPdRWIlcxOrYUtXrI
rm/523LqLDe4KEcS/pZrxtZVd1tbwZxEk2WcaHm9seXwQn9vcWeUg8imlIV82+vy5Cy2KhMKhuVv
3Zv95HIkv5LK41zRZUpHKipVfkexi9pO+amsReSqZD1+nEITbsBjVt6wp9B6SHSoTkW12AyCkxS3
TbFTGjHn44XOU70DVbWx22XqY9DdjZJTmLpwj/WMwzuhFfisRzxtnzWXqnAvD/FdN2dZb3KjLslu
5nBwqVBIjSukW8cCZTZtd/Xw7P3cLgx9RX3K5vGkWE6Gv7rYfhuex4fe52q+p3dVw0nDWstkbi+3
YnC9lVi4pU6a3u87GXx/BX1zYBWrqUCSwXMTdIh5Yr42Zc3ROOY3f1Gl/C4bc5Vti/ORA3CTpx3O
oJUt2gkBKv4jGVpUZJXpW4VmprJyJramtRLEKBfTAV6z0/ME6Q0vZKJI3wFTol1yA36+9gjiDPgN
kwidB88lE5vrg1A5ZoQPXSiMQMID6km6q7yf2hlCjFfqRtrPMy2nsWAoV4TtKEK1dQzc7i9GvNST
wnQGldfL6x2vFhU/ZU9wahE6yYtYOsTAdiRfabjnitO1ZHEXJbBHtoBucgts25mdiRkio/psg72I
5QqhRo7STTcZT+R3rM1Wyl46E7R950bpY5KItuo3aEjPb1CANo63zSKF8swUtCQdQ+PVkuvEXxFp
4Ti5N0Vafr0WPoN3l4h5M5eWpJy9wMknBh+530KXfByIVVKuTmP0fGkqhvGxtfSh5DW3o0VD30HS
xqdJP0NR+YomZlqg3lS7rWzjpjR6VxXyUXyw9ELPpbV8Rkb50Z+UGgly3HOKDjiEr8l7y1SxdySW
3DIfq6VWrYiVKnBAfd90Agai1nugMpxEu8XZVOXlcw9OASmZXaXjYnXg7r8Ozdd4Xpa/qxoXeM4q
y5ac6PllZclRQgqGEKJye1daOkjDsjDwpXJguC0K9t/s4ZSbvTBV8iEz0ZfaF58WMlj1UKhSeTPv
xeHNbK6V6P9iaAybLXa5GvyXge1g/J9HV6sCD+MwUN+5R6ZbjkZ4E3MY/OSMJzji1PlPDtpyuOgU
qLmDZREYknHX4w/6CgtaZEf71315HkIcnrp0CLaAIR/D+cErDzZNejXvM5mJajUgKqgfknvfemiJ
HWtI2Ew6O2Keg4QlxBtfuRYeVXpQSUBdvYsgyzBRab3+8q2nLJU76ekTE5XBDG+cyvziwgkjYtlY
zrEJmSO+XcvBTd36zQ/fUdnKQ465Xps/gzJ2QWd6bEWY6vgVPmm/SJ+SHBt57MBLMrU3zIUMZr1Q
1fEjgYrlczloXZw39UL3SAyLQaU8/5E0EAOXt9l0pxHLa6uFO1VOEu53+H24Kk56KVVkRhMbX9Q3
lfLWjSiDxIeqnWini7s5lCdMB/an/7u9hOJBH9maqwXlo9eF/FyL53MTXHSg/sAfkJVaV67Bm+rL
MVrY2T5NTsyBHfjGR/SAw8iFkaXOglIfZgj3qhauzmWWr4CfNWigwMOCfJFrEOfSnrszi02dhIsK
HIK2Fweu0IwCV2r2P3/owsdGSi3V5tynNVHfas+3mBow0v6tjhNT4qAzfISKatUTtmY8tQqm67tT
NfGy/ejrShgmjw0oYsBrtWsfBCuyOiKMXaPaRz+rDsZV1ALNpWIrPewb7em/dzQsiKla3e02CbnL
mJi4KHBqtyivZVMH15ohWT/K49uRtAkRsd6bJa+LWHsaK+54g+BjBjoScMWYgfOW/NVVcpGAr8h1
79qkoiapKQdcGIN8tKfj+ZV6GxMxpYTVXkbYhUoodQveHMyNTenoz5XTCz+SO8gFcOQehQdnv2xJ
BSutfcW+5HEs87fEYGiuFz8HxkUTuVUEDzP0E8kK3vM7bSyUNt1IcsctB8KYlDK4gSuoDq8trfLl
wh+LtNHtnYgoTqpdqjv+++vP01/7mQ7lWUtttdB22YJ6Ge4hZCj6m8g+Y6tYK1fy74qIi2D9RzY0
ki+bBu8rpvaHeldui2xLbbyCU7u9yxzzTlMSBOf4pvgm4BRvUSJDG+HuWbIRcvMpLdOtEFAHqBxM
XJDMTg1/iHDsq5boz4LDeHj4x+dT6KBR2WMwRf4CJyoUGCuOTZVyQ3JVuR7gg2LdRPEd92nzwltq
hMP/AOcfCjwvcZyDPIDCDbgmuvlexRo+8vC4vyaxLfACRaYYoLIEfUhGRTC9kuVLsDfVqzuZwsJo
jUjd/RPELbPBEpqhjSbdeAeddTwgJVrQoVdcu/7qpmoq3txaj48gYdEJuSgXUSWqR8+IbUJsIHry
7BkCpmFdLc5lamFL+RGtaOLx9DoZxKPVlM6he43VPLPjrCNDzLLmU/Jw8VjHc0ozA0jkKkZv8l/v
zO/HB6+iS6P3jL36vpSScrPVt3Mhjze3eBA8LJ3Syad1/A3EvaxDp8BHJihxJWvkZgwBO+J/bJub
EVC+JHGAArZ9IUCwjKLYvlBb/GOLqEtAQntvBGVMwV4y1/jht4UeRDeZwTN03Zfn0pwikD5bIwa+
1dIO0rY6UZ4Y6Dihe4CjsbbCwolwVrA+UYMjqeLiKKF/2biotoTu4oNyIYMrerVX148RVJQ0pelB
Zp1+4mIHSIOHJFbvxU4vFLrAZK1jrXpEq2DnktK6vUKSyQU9dCi5fQVagQByxKrw4jD2I/VxfBBf
1IhYKPwaz9wkr2vR+OIUlZBcM3ewUxpJCYahi9yAxWaSoekt7HSsCL8BhI45UIkrEES8vSfOHsb7
oFb1X/zp0YV87KOs64sAZMNHWqHG5+NtcmRvsSXcGo3z6gVm7S4nCKR68GH/SidADbgUjhe1seiA
L/AZJnXpVTihA582NeQ5E5JOE5HlWPPv8rITUYDiYhABwQKsHrWpbdrTskbgRv76n7w40PLu3cSJ
z5pawR9R9WKueAN4ITqs707f/1+aA4nE6Q2zqxgwBwDnU2r2NcvQgjDdRerFwOI0vLshbOiKuFCE
HDcnwvog/qFrviPcAorTADoJRrhyKaecoAFjsxqOR1matKoQ7vFm0QyKVDU0HkEB7U49j9HDucME
O69iE5L7XsBcYI7qGoWpzeHVoxcI8gYdFg/dnmCneyLT5kH4aEw5SlrJe1jRA1F0aO0IqNfJM4sQ
LZGlk8cxYdCpERN+ADCpj9t+EBOvrcHK5BpfHCH3VzryrZVkg8qGFptVz2/S6rInSpl6x28331vK
zc2BEllJ1/BmV187n8gFz5hp7WGnas0a2jXdUlhMvDyTbrbLRrP1pspTyv7I8ZEFFCRebp8GOJsv
BP5Ss4xtHT5kM/t1hYKUIBPD7L9t9xOuROIz/1y6aHx5gXXYs5ZProeUH4CJz+AtJIU6s8e8oyL1
4stOLnHQJjSSMHeU0CzKV0D99pBuyZCMfOIVwXfV7AV9rCPl9pnyjZ7Ew9lPcXBZrNf+cLPSd+Iv
0C3QQ6PT26wXEpfIC0SFhloAjlw+w8OQwMuBp2wauUbuWepp/BisgU0wblNqSepWmcRnEcpGeJX7
GemUl58BZy5c9AcmvwpZyt/nYw+5solYjjn/A4iQ2LyPE2B4qhLX3g/qG23wghk3ItM1lNWpcaI4
eou5oRP8C16SPiKezcsa53jdMLqKWUVKc+RNMyPuHPiAPOYtaXDcxhfB4WQK0k+GFn3BGsvk99id
5m+8on0WQki9uhvL32thRGE3C08aiFDvz68QdnjWk2yyLR+TUVqkYi3yJKW9y20MsCzKXJrAul75
e+cExxsdppujl2SC5DiwpSPqt27M+MD37OaVsSU5bl+wUE2f5MGyr/L/QP2SGZGWzn3whX8W4mbI
QAC1zGO6BlfTRUl/uLBYigwj9+HxuoBKkw7BKD3hAraNk2UzdESbKhoNItQhHm1Rl299QOy6j75j
AMAioGgN5Ajg/JjJM4wu5jtc0VtGxhIxqo4vSPegVco2P1otjkIKGVJCpk1KFCI/agUHDYk9cI5Z
9L2zPWMmTQ0nxyTqKETxx8f/l5+M3KPTC8EEGzn7LFTC93R0ZkNm/XbwjVsFWQ/rgtCY9is5Ks0u
7WF4Qu/J8d9iQMatA7bkfrioIcAfTZBygQHTYgK0fYNa6OLlc2g5E/r354tnONgtLNQH7qUISX3u
3lJCkpdZGpIYQ2UPtlcYOfur70+T5sZr7kSkHwWt1pPRCqfzsuLk4bJY/sEemgBdwthBF7arRcTw
dFu/+mMGYt9N0MwVCSeMHCNiCFjswV1d2/QD8ds8nsXcD0tN3Pf4kb2WN04CjMj2xiXYyxIJkgfc
MmxgSSXOVfdUiDhkK8EvT7XgEZl1Io/hCyUDG9P3gjKWh4PQHKXgNQC225P2gJMZEhgGkOXZAEP0
5rWpGshv0Xhcx0Tc9/+9VAvOgyiwghW5bGg1YQ2ssGjTy1yKsiW3VV281+Q+ltZgBpyvxZFASXwz
AijnoH8avAnHsJbMHktMd1SdFfBROMNo+m8jZysaTehbOcJUvCFSCTwKxXT+JOqxRk3Wlde/vUp/
oQdr+U8raXGAtZI2Jq+cPf7s3FOByaQCb1IFjGUKyrJIv6Jl4gVPDUD3umJzFehwQPN353fPXKw4
YMnPo5AWW6YGKlcro03yUVs46VqDk+VozKpB6lhLTcaNLkCqyZLI6wxmDmHn/OZmBCk1cf8456r0
fRoLCMcV9GXqF0QhcmaHVTlakltCNdR7WWQZonfAfKpb2lDKAd7XuP/7qbIiaYOWh58WS857GPRv
CMumxqlFdhbaMNlVnwQhblunK/Xr79cwHCNf/Q3fXKFqDN3Uu4Dk7yoaRHjZA0xPh8VHzAilgVGZ
bhXf0xamf8A/mZmTnfWglCqgO2zPgj6c89CxcceKRJncQiPs6ESr2p0o9Lz8gKKJ9O8PE3rO+qQs
hrKQPissGIwEdJT2Nw5sAXIR6hg6zgUur48OUMpnkGiESFlI63YNRYeZaQuzyFBaUgHv/IzwfhJp
pzWrxg4ghuDErJr57+rNQ0nD2xU9KXayQFXtoT4caAJu2H9IANB+NAS9CBnXmNKt0+hfgsqz977z
XvrE5xLABNt7kcwo2gTlKs91OGdIUzUDIC7zY7Zxk9hOsdBRgxG/+q2t1BS0bLvqoTt9jNVJEa4w
eh1tpir8uAIHlvas39XpR099Nv7Ksakdazs4Ku+Ob3SyXBrBmevQSKIoylhnRzLGsljMkqMsaHYp
KXdWJg1nwwkO0+h6D3Nrdyruj2z3Xe3Avnd3ZB2RUblkc+nDLuWo1ykvZjwucrvFjVKBWFazQsDN
83uf65Ac7ibdquUjfiKHuMr4aks0b/wEL4ExDhXofGNevjuRdA2xOfurPgYs5MGqTJmenaovEbki
VRF0OkAhuCW8eVHrFSazfiPnXbLYRZtzJ6OqD6iuW3A7z/K7zI72BOFO6P6d7XhpbIA2Em2W98Sg
pP+zdF0lOD+a9JvtOBT6oL4sjZf5uzD5dvkMEx1wbeSKXjfrbZ5zOnbIQmjLkSCI3ypVodQOYV8S
e+oZRHNl5qj9mguBvlJc9Bm17cONZUokszzmzVYI2fCjFfFtUukTCd7I7gDnhOKSEkcQC4HZgYbt
xWzS2Eu0CgqQa5VS3AHrlzSs+pBovOxTBMncXgyBD6yCFyxLCUTq1Zltgz5QzZjmtwDq+fBjfbyE
I8D+0+DVtkyyy7ZCqcPR4G+8L/yOWvESEg1UO9dLT4gD30m11rRdqlHMSd9FHLnVeVLDYHyjnTTF
Na+3PWQ79ctFN29kR4p0ewxnFshNJ56a7m4zvBDnVrpRCv4Fr7aOqf/JWsp+lrwu/LEUrpAr7BbP
A2hwJNk0FlWvA/rKXD5fNXF7EdmAwANUZ7Z5NqSluNapBcXNQldfblTvh4kGVTybizbHORUKCXtQ
lFlhcEMKgqGs4e+f6LwBK77G3HqEgwWhqGczG9/T9QUMoIT/9stk//IKtT6wt30Gp1bxZBFD9Q2g
ZLa9eX2FeQpWoNqsNJ4jiEOAV+A6yPTdrm+zOLsvVkiqd+j8ugLjZn2c2vAMB/IHaKuvnTjlmh7a
9OWtJwkCBnkmPUomPxxpBdWtnzwT2WQIw4EUGVMB9kUKWFTrFYKGLIhcIvZTpaAD2nlV24y4u1SG
OB9pny0f/ykALq4CEPmCV3LEhvVWgqt+Iz9NTYdH+xvQCWGy9SWGlfJXFN0kXDiWfjOTcaPDlqjn
4wLfyVFRpt7ruzUoCeQm64m7JLCxebxrmxhGJ/YLRfN/9PkwPeScmuF6dl2205WoWx1HipGUIkHq
mFFehHR+e61c+OMFlyjz0K4jvpsKLrtmG9vBN5sk01uwoLeQlKSVTRwMlFdKqNWu0QpecSK6N0Yq
LQeB6GPaABTewtiSmo+TbjX/Phk7f9MCXSznFGNsubA60k0ogvK/9UQyXXnpp7RfiMCRM4q+bGXI
SDpNNiEdV/LdnCOeIAKcNzUtWXWZV94dQ+ORdhqXm74MDplp35cMSmMdz6VdpgBjyLvQhJTD8LeS
E46IqxvxbFJ3mIxZ2vmuLme5OceBB0MGrv/cXr0Em0R5oO/D/UToNejXLNW+pi5hE2FI+6Wc2/X2
DJP+l1ppOpYcGBSjJpKq0eSRsixTrbRIcmBXxjagTdJ+cYx6wPSi/xxiznfwOfUq2oGWux66EWmF
EajV352fY0qIvmwqedvFH3fH5xABGM44+VcHkT8h02RnYl5y9oQ/12hH7X1NCH9vL4JAZoGOBDYI
jJyK/gjUbt4Wo3ejEFasEhsz/apjd17sNoywEzMXy1YVPi6uA5w099VbH0nx2bMXc7OVIv6y3zHg
MTlxx11cnMz6O3Hv8JSx+R8Vqj6lzJajVtxRDqkQcZdVtFcjfxP4c61cSHqth5g0Q+OhRbmxM2YI
iYJ2XaM7X1lF4A/vQk9Y/YP0dZ4v5lkPDdtN6AbvZo10pOaOOa7wp3jya2ymvSZ3Xkz8S6oDC+tc
+mxG70CMS/qgmd9hyO1ibcjrjPNUd7v1+0RJwXyxa/KizG2L1/9cEYkROjlPCBmQGQwioqDZ9w/C
EN//sANzAou8ZNS8QFtDX5YstnS2uerW8KoOuqjOyKZSp/hK5xopP3tZIu4QQwVAgzHzogbSBJhV
n/OXWYBy47LFxCp8AdnR9TJWNAekgw3/AMQxqcCoQg0gdjAqFcuseg0WJXjUAT5+sE5bUldGS3Mx
a6SSltm7L1xIQqQ9Tb/L0lQXiavK5hIIoeeQCqxMtrXAUUDF4BmxnBBJPucoD94BkGU9R8UG54kU
kVerMbO4aamytpUqzRDN+BGhk1XrjxeFA1NWzveqoJIPu6wko4I4yZOzp0VOkRDA9h42UFGMhv9V
p0p4PEIAOPTZNV2qiBhsLZmIMZfevPYO7KxHuqMs3XQD47rRicH5gGtUpggs5WzJCvg0OxuCLRO3
csyrKDv3cGJKJs4q2aJeMkfSlQ5xgLYOVqzx6bYt7ikMqWTivAXsUeBECVLz9vhZ+0PyM7QnKITF
Lnij7Fq9WciJ3ggXtwgSCQr0rMXVcofKDLSs/wt3+WczCmG696E7cuzw3Smf4rZfmXIVLnVnvgm9
c+VIWPtsCF4Xpp4NZri0M6LuG3KhorlRiVDPEaAnTm7QiYN2eQo7Tou2PqrIrL0n1FThbqd7EObd
5iqZT6E2HFTYqTQ8sajbIeQO9iOWvo+x99mp28aAVr2990q7SWVzU2tSeNszuXRB2U15xa9JSEgM
0rih1EjIaIdmv/YHU9yt2MkWupUlFsIRc8jioPEjASFg1sd/cPnOgUeY1q+es791Eq7Tt4D3hdPe
qTEsg7KKEoKiIMlyvewGC+/Wex0GqHWV0yVLxXnmeIpjqfe9wIF/Yce/4PL3T90+w8vrRJBFkdVv
guOoxncJPn3Kx4xxT0IOkEPzysKQQgROzILCcp6aew5EZX2sfF+bI2b3N1Z0MpxL1Rq2l7EhaMeR
spvzKtV7CGO5UBt/H4eAeX03gJa2QUaBqeGhyNIoJMYtmVDDtslztjjkWqyDQTt7QNrvDe/AsP6D
oT9hyLqpXbD4fkJeJZs3gcxEw8WPt+JqiNp7ttoqdiv7rYmnNbnfaIizq9dQHzlwAcW3uXHVRxnw
fkbDhUCxEok+51FwdK3nhrLhUGvOaFeF8/1OLolnBBjCXir1BxhEm5sAybZ9AZ3yXhmU9+xFqGPb
LqUhn+OdY27GItpgV+01nXwFWDs1cJ02EQWI00HuhTJ8SHbFZhl6cY6bcsRuERrvW6BEUwf+DcK6
tqlsdHfsoo31CbgxqlS6LbNn9DvvJhQvDCoXmtiANmVP8KGb8RIeIoU7/HG2wpW/AG/w7z228K4t
gjJUEjmLqH+62V+Cc/bpSz/7m8xLR70ulaji8dUGcy5krp1ChW41wFkRILevYeVJPDMiaL7Ud0Ji
9aj4JMokTAx64PX3oDwDkvoEvJ8BUW2fj2jY4M2nR4ArBQfBzqtJDgUssRpa8irIIenFmRJ9lmJk
16E5II4d8LThN92oQ98iXa7q8rmyo9nyb4cCTkvGw6zzLQqf3lq2m1CtEu13qSLOYKqHAULAlBXQ
TIakYbLBKZspTKAFwfM299TMGlODPdCY9QNJColy/IzwOwNSYzqNqRR5OvnXuuNkt+2U2Y6FMslg
/x2jHNoWplZ7cbI1PqOanGZ4s5y1J/+iKsVkNpEDUzm1VT+x0FSCbQwNsuErlw3mEt7cvKF21xpg
O5Pfa6Ss/4N8nIHjChk73Oy/D97Czp0jG9PlnrPbhs+vbG4eCubS0eUivQCHancwUtdDfnD/MsFs
sqrUx4eDgejJOP2wZzxQVPzLO8UCWNQ0fZcvgZX3FaDOwN/raSrlqhW1fhyIdJdkmvfRf36/GZb0
94Oj1CmHcSizzoDcUFpr25V7DFdYHuYYRhH9cx73NZs0RQw13fWBoAUlhvhQE0EftJlsUALL73OV
bkwOi9qcm+p/PbCXd1w9Du0aZbgtIMB1B20V+rsWWCbSxKtYf4vPUTg+f9gPlfYQj5e4HaH0dS9/
l+sooITZJZRPaNKlqCG1Eax1X2tj7/a5+w0zKgRWU3rrcoCiH8S4fUBf79miRCQxZsSvBoyZEdwD
lTAB6R4fjYfT0CfdGQX7f6dY0Ud1x4AEMF3s/2pMym6a54fvyih+aaUoDwellGmsfhBbieoqKoMD
RbiSEUB1d2vha2m05DkgkRXkYZmdWJ+wxFwwSYRKr19/HzHmceF2Nd7yf6RQzrYqSkYCACRi/dV6
Y1LTbZTAEkbiIFTRw78O7XM76AqCAUT0gUlGL1ROgYxw2714obaH5EF16cfK0ftt9PWzCq5IvV84
94z7PvxbBtfhEZPmSMBe1a+n5UlvUlpIAJAhyvZtltS9AR270RseR3XWJ/UzwjOFpV9MC/RDZM8S
agvnDJqto8Lxq8hny6x/FT6qmNww5plATYJvjbGLjDIwdBXL7EOCiiT9Ut8Chr0tOxPjouNiJLwy
d+Mvm0FDDtHWuDl2a+4ozkCnYyw1Ufgh8ZDfCILRvjjB11vulMP2tgxj5yNCUwvKNj1MS/e+AYW+
p3DXYrJw5SuA0DdZ1uxl2EH9w1iMQMzfwKMhBtwOvJNxH21Em/PoJh2HTllnv2mmWiBtfq2ysT7g
D+EbuAcvL31v/dlT8E+Lo7+pz4NMpMvcQCW0eUVmubxyEdWvhM+XbVZfy3uk30yahQhHcJqr/EDK
yM7DIXJxcjE+OitS5h8U2oZXeAF0dVcIpyn10JM8uQBpbC4XA222QL9FNJpPYjaxbVlVO+4HVsks
Ml4I3exvUhBdR1rtb9B8pEhAq+ocpsd0pOyM1mpYQd4393lxPKHWyMLA2abkJ5nQRO2XDmaHmcZ0
C56P3BWmcF6g8fNmXk8oa+UC+7T+NLOkxK8lqiNEhG026slZZ9w4capPMgPbLkwTilER8CaQtNSU
SYiIX6Ot6eo9Wuhl4K/ZLf7VSqioRKLAFjndMmqBgqBg1MlbGlrqMX/aG/imJB0OpTtXFV0ps9n5
XuiS8ipKiWne9tOQkI8h64w+uw9sVtZ/vy23KhMbQKg11wALtcUs2cJR5aGil+yLwCfpmmNt2H/8
p2c3XFdFr/HOlfCL22Xqu3Fi4NYDR9SnKOzzFcp2UgF1rYkUNLfBtzpvZewznGsM3o5UAo4tueos
qFqBRU8bkp7Lihv+w4zyd0sAroH8pKBtBU1MHqRzN+u26YQra0yQN5ArynZDULC9bZuGNnAOlGvI
MfPADgZUGe25P4KCgEtiUkauRhx1XCIPSBbpfjd4BpODHZw2DqzSfSsvbpSgQl8Das3uHVCt5ww6
rsKbP7NxzhCKTByYD2xHVzf9jDnRydVaVuyrPTZBwQlVuOSUOjQfQjDenJJDnfBf+ETI3NPBrKqh
szO+M2/98p5YLKHnslVBS82EppdiaUlp3aa2NS/LZg9dUgmsEvpcN4koic9/v9vHyAN+V/V3MVXo
NdS2+jGOvvyKCh5yu/lx0/FWsMUPLC1aNJn8CNEP5eNua6pnV96rlgpGr26uyIjvKrpnTLN5+Ru0
wHdpotlrIzoR0cxyrBi6OeiAp5mNs097rGjAQAj8myT29xtmL/pOcgtc2p5GolCJB8yk6ZTrFTXP
D1z6PPg/JzB3wKPkvy8jkYzBJAU7/TmUDFaNwZYhx0mgc+QqYY17eeJY0eiWtHbFTYKgEN9TA5L5
bKDDWLlNb0Gziz7LFpYTZO1+neT3HO5fyrgYSDOad5abtduabNaFfQEdAKLNnhmfCjcL5XxKc8iA
MpNHILKpIVWRK8LbMaU8JTeKXbJgjxn1ZooTHM/14KTPV9mGKV5VQ94f//n3LrRvOudvMwNy5Kcn
KRe5W7jR2cETKlVr8DBP0oZLKDltWSqNATcKQTiNuqVNq+h1nkmv+Fxfp6tlm2EMKz7NHhHa9OBH
0t6v17LNUdtUGE8Dkj+TgYfiv/FPdcuMktYMBTAVdf/FC45c+tH5kJKrpQK+5BnH4DmTVRkNg/ug
wI5kDb7ArnzN1P8FqB9lJDSEgohHeUjyiMHJR01QLRYpJ+jxvKIvAJM6y9WOmMneswTIiHCVbPRj
u5uJaJ+OdRHuik3p6NJ5DOezuMUpFatTzjHGQE3spTGcsyu6taHnuU6MRG84UHXEJE85E+5Ylc79
ZcWmz6Omu6FSQ/IZI+fjciSWzdkI47KKDL7gELRS2ULc5oNrzliD/fypX2BnP3ffuFiKI0hTqfi7
AoFXwur9MrQPmaAk7SHdtOnyoQh1GjyM/mS63+U3MeL19HDc6NzLqyqvZTweZwKDOSBq1dD/GMSa
Am6m0ovzd8SGKjx2zYaKNqNPaIHzM0UHxbR8+DBQ+VIRErHuOffrFGRm+eV1FM8YYXYWRTZuCFF0
JG7dDDNKgX0c70VinNqA5jBliSzGyAEm/hshHmexulxk/G3ZqzHzr+tyX82gWQGCUrqllHrpOh6y
yYGf8ZDCSfFH7urCatyr0SUPIFkKOd5i2xJSY6LxjTnKYTH/6FWoILIMePxJufHrsxN636T/ZFaI
bELZEFqWQamYLGUYLLIEiU8i9c9f2f//zhE6/QBWpMawYE3jK+IuW0Y8CJeQEwrVvgKxbL323i3t
koRG1zA6oQdRYXB5fWDVJNDXNXssou46zPxlIhQ2chD5j98AZQe32odk05bIX9lt1VKBtRVxx/V7
qEzfZBFdTIrkyCXyQmU7rMHRz4BungKh/YA8pPQsx94XXjgMvfCWfGMdcV3pgn501eAtjIyzanbZ
lrw91CkxEH25EBvh4NIzmAmxreLBqZ/JwYdfOuEtgC4T8iSxRagFsE1N5CQKqcG/ViqtGfrXckdm
PCTAkzgBb1vICoZOLm5y0424oZNyIyQUQDVJ+sBKEOPKu2U7L3ggVOlbHidytKzMzJsfRwB+rs9R
AlHZeMe2V1vBmKLqadkjYa6HGmEiil+feaZRUtKH/I1cCM+K/dIo4anGeGBTGoSxxwYLu4Oe7yPr
Tl5sczMNJ8lsLDiZAhJjDfgD+zmEoQSMdljthwtMkW2U1mftONlV+IICWUoKhTKGpvXUl1yTh2VZ
9pZw+GFa2cgO6twbh3PbMI36hTLLeOq5O/6pPEnir4cIFzy2hI8/Yq1PFUZSiyZ92YCtLYv33SRi
z6q6bKuugJ2TZeWHo6nynDdx+ht6fkFxhX5OjjkdxK8dq/h26euphBUeZok4NXcww/QLiIiA6czx
guIcntIKip7WiqAqgfUwjpjO/K2Cfm0nqoRNBU8UIr2Mw0dJ/eeutHSpNup23MtE97lDAAVEbrNz
iFNsS8UW29OduSp+0x45G/FLnLNU7VQAiMXTl3o/58oPDvRDjK1P4/fGJiy1haKitkLMljrKx9/8
z0cGb+EhfplCi1i/pzs0OsD8cKGUxj6yV4/K+7tEEBAnV/AdJboYBuMjsihe/Zt5t//n2Zt0INAS
YqhpnhxWnGuWu8MmIN1ZcocPoh32pBfvH5mEzFtgHqWY8GNljgi0r6qaSln5fYDBRGCDrS/Jsvxa
1osu+zJFB1a9XX5oqscOgeKoHvErvscgxH/3uqF17NB8bTRgVDW+qtxZ9fZ1AnN2V3dvpnbjyIs+
pIIna25Jf9XZ5L7kJiiXkEX+jbxBhmBaUmUVpIrSufAsULTYFuGpfCJ4agzFbSlRxapndB8EBStT
H8Yy5vjoCQ79k5Au29iaCwxyivMcVEyYB1vjtvYCWcdggrJznaVnlAKkUXZ5qmcVlRBcg3d9hR+y
A3qBFI63mZmSp/FfMmqk+yBr5PmBFfXG0q8YatnT5UEfzdcJJbZ9WUTvfGIDL2htbT/ACtmUatnK
TYT3j4n+M7Soq+2sQxFif6RIFRUCIZ5r8N9cEaPbrNAGxpXnIvErsObWdG3WQUy0jYclkq81LMG6
vdobVh2SbSgFGnsFc4FNHheBN7SmXvtJITfJeJ82iGb8dSn6/gNx7Ibrxct6+0RKpzVAhrDxZgAW
o01obYtnDIfcmQHwAE9pq9HdP9HLvLGDgv0a0RhdHMVUIcDKdwqGMUHy+PiFw2B40plknfyroKKd
qCAh0MjQWRS0CL4zUood234gUgSZisLV/V9Gm+PVvRFl6NPtHOCMdkzoLcYgKnEn4dOzl9zSYiOf
4FVKbtdNld6FoxzdUz+fvIZrqlQQRHxofU5r4Y8B6b9+/yMdP66m7Bef6XXVJM4lMvuZWV178vGG
2HRLJt/vcIj3xdOHvxliXNmu+uChie7R2+66Dl6QwANsXwSyLiEcoro8W58KP6+HdEGZDuQU6XFh
hgDgXBYZOeuI+qcYQnOaskHUQizePkLk0kw+BKdfPSbSLBJ8uLtU/Bj1lhz3M2A4vV2CezZVvBn1
LbnkihDRo6tV3YTNPaC+xAiQ8VDg2Tlo0Apdy8H5AkftyIePZ1rq5bWu3p81rkWYblWL3LPk3mrW
M0jBrTKja8mle8n5C06s+GB0Yw1Lg6Z5IIygG4G7U1Z4f2usmjGgRkub3UreCEPJjky9Iot5L2nY
utYE5H5eNbRDVcC/XJ8oMXG3umfR33urEpmVcR6HvCETBMhvdKPEyjJGxr+1kIBI1pI+5+pHrJx2
4OkBbuQdIFdel4FAh6jWtM9FgHLgymlPxt0ZiYLZoa5W3AeYZuENSoDy29hkHOXOFAcIA01Cy1/i
roBkxFo5nIwNRIBnnUzX1fTHc4racDS8rlns5YWbPI6RoJ3XRu8Qw8z3ImEFqG9xPT5o8d+2aoHk
jk2lXXgSFn/uVTB7rlP2+hCnOIw3emPESn6y2sPXx/spmcsdg1zbzUvHKRrsUKrbLmLEQh3zRWiZ
yXsLdhCEMbEwbcLw+qmY2Ll25wUs60Y1xZuBVqqzSnCrL75qhRBdxaNQCRvabv3cbDqp+pJxLGFd
kHKT85R7xxnD8qIotg0XhXY2Sgp6IK+tsMoltcbTtwNGyMS6f34yJnUXEX87gNZ0h6Z15rFeU5jX
cJsCgY3xgW08CT5hAtPRf7Lz+R4TFjILGcKXJtjtUDYoik5CTu6cIpNZqIhwFeMQFn8jsRzo7KPn
Q+ep4Y9zAer3dwE1PorI7q2irobQRthd/ivcFF/NrciDsCQk3car1Xa7C797BjLNLkNuZEzRP4wY
x/sVzsGBYTp3tuNTnIrfeG9MyG1I0kz4mXVYSyj3wNThd8NOOsATZA2NbYM/s1ZB1V8IJecJX9KR
MJPKGcZG+bQkKVLkyW/Dx936H9ard0HHjsBtcawu3ThbjfeH0iOcs+4Y321h+UKqb5tAd9ZbuJo8
S+uokwBTVP8pbKee5CjATEzDYdwaEhT/Py5FhV6R+sZPLOENW3baB+pnB9GqVa+gUZ3jw3xSk0ee
gciCep4GFtTMasnq5g0EH+4qjIqmcAzJmVHb3z4i2+Fsrg8hDsHlU4UC2lQNia05Be74ft9cy5fL
ooG/MxselNmhUxapElnCrdmXl6sQQMiMwIVLGaPWFFRK7Tcnt0+TRmiD9VOfyOIgavrRV1k+ECvt
p9tT3KqfI4DMrXRXCtsu0A==
`protect end_protected

