

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GuWEw077quLd3kfu8DABFf0P+6oHLq5R3U5znEygNXmkCks1DFRW7Mt6/jd95Z4sdDaR5vCLL2M6
FB/Ff+rNvA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jFvcfNCzhBWpeT533DDm5MsDXv4GiB5r4Bmmnk5Von/5jho0+BIo5IwIRMf+AlV4xqtSYYHC3I2k
BVrljYddp4kTGUJvHCrm4WaY6cktxQlEnZCt6LbtmRJq5bQ0+BhbjRb+yhnUtxVO+mqZJ8X5carS
6TiI+a3eiQyqjafsIxQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3uk2ioXVXgv772p2rHBKB55nN0zepBz6/NR5erkVu2PDHMiL0sh4KhStRZxPeDNzjzcvfXxTocKd
hKd8wwyqbvI0xJMti7Zm3ArPWxG9sxsPGJWi/HV3nwjRdbl8Q5i42ko8FFW76K8gPbQTkcXqEX+f
TMDFgnzTvHtLMrE1Xm+zXTsDfz2iY7i6oQ9oV094lrdSLAt80D9E8ysTFrLsOAY7rvOt1c8o26ui
lfC5xFONM+l+w+GytYmCYLC1g3/Ymlqj+CUT7JBGrc9OLEVB2jBY9OOPdBfOl49VdH6n2k4l06g4
tPQ+CDbASlaP1IKOpWeipcMMiP2EcvQEvzBqvw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ODN1qSeI0EeO28pILhOMZHx9bb2qYpmwvyQXvKPrPhpTBylybxluT1/v8KSBCRH/tKp0Ke1TAM0D
rxIBcEp/+xGCTqhzkt5p1fRCsGDy/1Kk5L4fYaTlJRk43uSfOTxn6cMlcuTzjFQ5x+FkobtNDSvc
hzmRwInNRUY241xhR0o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dC/Y1fV+mqTG5rOr6IWyGTQ8KnFRPeLZShUWaAXrkw+Ng+xoimVrmPwEeCnURpwc/T0yNbEjCDB4
bGeW47AlClSVksRroIGKMbG4EdH+85GyM7JEd8UxBfmIEn2qUdv8H40fYW6ndPlPBbIsiprcQqu1
BO1TrP+zbizezYEZNLdme7klmciNF64y46dVM3KfXIDNKQvoLTlpJYClTv0K9dc9pDZOVD/5ly4k
Nh9OSLv/jIhCDn0y3M3rX1DyQgZeJYBkDd4IBP3NH/wojvEFQZAcMKJEqADK3qsWu81U6IIzKfXC
PUyRFWat+MUxb64pAuTyWw3derZjtBnOfD89TQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54432)
`protect data_block
UhGQ2BOIbPKfW8F2bj2D2WgMdpDjUKmEP40Z1QeYtmTJ07Q/SzPaWJN73ncdANdj/QHSLjii9Omj
ZhDmlLpoGLvozlDxgLeFRhjAoIdk1M9MCZdUmpwwO44cCmdZL5iMGpHNdyiR89SBJk4+TECJSo+l
SsQdSJxqlgjr89G9SSiCFJhDkYQWBbiizbM1cOUSClQUmTchiR6AtnDZGAyQ3SeO0jkPHlFs+BVf
Njz6g0tSJ1o0lgX9AoMRxB3CHnsWeNcbYLRzWcjBnBIa6pRlq9VzeffxbtMwAPAKBwPPKCvpqjcB
eGXpu533FKy6WLos7GX0DFc4RsG2/7erA+5sT3m6dAuIo3GKX3SOVWNMbY8EKFb2vnFE3kuzh1Qx
ke0auL62f9Wp5FL3jVIMatAGFjdxSQQIAaweIhkJxnj2369vX42Pj+kjS0gcyNap2iCzN83wlJgn
QQw7mtyYVmdkMfH/t8XsFRhq/BjqQSGzIcNPJvRxCLL66+0goNm2Gv1cKG8dLUOjjaQzCSyRWwms
hoicoYio1nwH8UAlOYh7e7xsA/I29ynyM7fHgsR0NAJhBJpwl0Ae8bS6qLRzqgibRUooYrMEfm9O
Zid4t7CztHzIXoV5mcZ6hP/I9AiePcXzJjy2gYMupxjiq2PKOF9C6/iNf2mWCCsNwNrTWDh30y67
NyWHcOruxOCz6DW1mAl4457+hyYReFlpUzLTXTT/bWbQGpG4O0c+h04CmXNX94pZxmlIJJTf/Kza
uBJCRMZwyOvgm85HznOC9l1Gh8Aoxf0RnNctWTia5rc3GFYEpAdVj4NFbh1phhjcOruEiam19R3V
NQXEg7VF6KBwDwss7FgULLf2UDEvf7ZzYLqzgVnUMQCr3oLBoIMZBbRothAh/BKFBj27oNfiyCcH
6CtLLOf9bSjnS6QetFn2C8yheIPmGDHeYlvuL5wW8R8tgRYs0/3UiQZQIqjcHSR3qcTXgLZvIhEz
zxVm/qqSteKiVpZVTcAcepGMU/erjrKqN6LKbwXivRruGkvK40gFdR8HSddU2uBrcYZahaXSclPT
JLYpupBdyOWmd5FzxcLmtEDlwmW/VevXF0cQoJdUmIMmm7p8ZdXIVMPfQUc+BtTVvKTShPCMUzzT
68m4ixI/WDd3bHuTKbQwZ1ymv/SkX5f7749SllIoiB6Yn50SGBJuo99Uh/WyBCz1zIIXTtxaGVeF
ydGFIs9EuKhKDo+mnxD8dK7PDPkFPQ8+9laHtjLfxtaYzkFQXj1/8oTPc6uRToTqeDUu3ldNdd7x
IdWG747HxhmeQqhjN9SPRLYQyW0wfoNpAcSOXXsKa+uN0r0egtds5cPEJtW3Emuh0edieNqfAOdl
pCNaK+DZzP6nC3JtGp17+OPeUpV0wCtJusgwrjJ9k2bWaGb7ukw9+M+jEDqK/BEwOQkthNGDtqkw
LGbYLlGp0gnMM1yVVoB9PXQqT/TGDTMdV+0VCAIWNeTxXrCab2+6bHlHfX4gEt7nGbF1+ymudjFO
9rR3A04iecqDz8quvvWfCxn9jLH8cgs8o4ZgtefsLZDrD1T7K/XJEW/oK4EKKUkVr1+XNrnzdkiQ
zxhecAE0KT4o/hzAnT1QvYkG9f+VcjCHvV6gGIUewZbqpHxMJM5I6QPw1wj7ZY6Jezo6Wc+jVXF9
+kHS14PN8PRRcH39aa4Zoo0+29R6bhySm27leZ4aud0SV7kVgfySu3ZZtXnchOa+H8vm599cNQUO
w4mYbuzK4TcvK1wTHsJYoPRBC0tDLKe8Tm8nN8p9G40m3h9bn+gguChf68V+n1zUrHqNq0DXFOR4
rVMbtRN0Atughl2R/mf/gs92TwTmRmqs5inEDEjRU1u+6H9BhYbO4dygRBBxiUjNgslY4Cd8AGf8
omL2pqBretDks8T05kmjmHErCCkE2eIjRBUcfl+yJleyAQYUJBguFfTfQ0s1ie/oVGPocFzoC/wv
Q3svcfVsV8U8B7wvx9tIRe9LUV1HrXpcq7w83brqEX6tE1E3ThJ9bBHE1t5dTSZRsbdtbI2jeDtC
oj59zqWx5O7Uz98nPJ2OsDuS6L3i68rDxh6CP+R/FnkM78NLWF5HLdBIHL0fONXAMWoAEjhjSbW8
xMILkdXVManSqwD4s2Tw2UWpcL5ACTkGmWs3WNpbWSsIcjIW+Jxz/6ZnKL9IhAb60HjJr3+mlpkX
+zXvxm++GeU4fwETe2wx5r+0MiS4Ni77DMfYgdjYNfwhNpdJ2DcB6qpI9cK7UcOlI7cmZ6L5YW6O
fvN/1ywzwzW7pbszOhd7Zl6VYGiLaq/pVZXEErYXxR9kYMpMkxic0HRGLivhOT2/0msDYV6pbTR/
xvWtypRqYNJKC23zB7/feouKY/s0Vs8M/e7/z5E73RnSdSAPgJNVXWQM9kRcA2Qd+Uz1dFp8NCtN
MvL1bgKdOjaKJ2MtX5VeQ3Y5wtBrEPZIawrxShMQ9RSqii2/+NGcWibOKp5MfTgwu2+qohVZkPuV
MFJym6F7mQ/UO2LI50dx1Qmje776MLD8CevXIRA1CY/a5PW82+BxC7A6/IVLwce+JVnc1FoXe00D
OLghOOSimmUNitxZPemMrcZSk1ReCLR+NwQnY3/L78v3YEWFzI0ZR9Q6dy29cqg4eu5MaNf3qiW4
K06vXDayT8fK+YDdWb3ZdpPHbognhm6hTC004pcvm4J+z5U0tZM8vY2McEeaoDZYhvC4D2W4CvSh
DzDHhvMAWEooxOnAZfjPMRjvfJbdrnml5SpgOPmyKN+sE9y3FclkjGbG4dQMHyseMkBRrTsiO8RU
zDouSm+QXS82J5zqkPV8F/h2MJAMfsUfocyLjT5cGkNxNtq+EzyeJcnrBr38iJUar0WHotKj2nib
2l/c2zNmIyDA/0XcNmST5DzKEd40K+UMepOrDN+RZnvaKxYBJWVLuqZ05Ek0A7M5uHAKP4OeO4Mz
/Au3vH4z3AXDkgcMMvO9bWvVUP2/DOJDbZVG5WQpfU5yVD2LcAVa25yXilffNd4L1rzhnmpTMmHw
5BfL06H08YrzI46aTSTl/7rpcGSGXX3jaR/lnxD1V7pPgc0uxlnxSeNA0N6AsskVxK8L75anRZVa
LuJNuwF6gSn2YCIxOdf58IRCB5jLRGsihzYSQzSnx8yNQbhCRtpCg5np4FkQl94wVfL9zwSnT2Fd
elTAxEIPWHSDVKmphEX/kiDBjnDqK3OsVslf/cqLwDLm4k2IN1CAbErGSVzNIHrz0KBhSudqRmx8
mB7QFBi21d8bCFxde4ajBNpui7Mw4Rf/aLIXwt+2a3D78C472qQqHyjU0lOLxoCC99lexe/k9swm
nEX7n7yo7P7UDRVJs++GPcJ2Cdwe3+HiMWG6c2iEnRNIakrpaRSxm2NzczGtb8tRel/P2Lra/GKE
HdWTwOizKVTppkn0LlFBAD7UO+Brf8q5ofnmQEigaS3k0ANEXQ1KWYM+/O+IkRVKE126WVPbeGuL
cRiRjKWOHwgLLGpM+sQjMmL0R16i+/bPVZudZ34sgI+L4rU1BQMEh6/41VqGPMmLhz8oKRkE4z2b
BRZ3NbVoCD210/GcxCEPHvAR/5Ahm00jysQMmHcJNsxIb05yCQVoJlVLwpKpCNVPoXdxkJnWyqyH
8WQGEUmbuYez/ZEZb+phF12vWXVeJM4XCXq4sbCreapSm6e/pJ7BfOgvDA9aPzd9n9Np01eisBpG
OGGQbh3tVr2uzMgWafeEP8vI1cFVoonpB92NT6UIZmg+NnlaKa3vIf98q30c+KbxCuQS9kNlh/xe
8Gq24aiWwnJmO2d48h+O7iHIX/k4NqORUpM4yA6KdulEA0qLcpqTHYI7nie9Qjyca62TRFyVYvu5
2TlL4QSYuwx5smW5NkhxUdN2wACeLtgBStU+sBUgsmfswT3S7QKfVQ6HtVZICIXcksic80YrRuX5
uGFP13+S6yzKqWFJWjnXWVX0uAvLxVPdzmM3gqfN+wjVmAfp8QDBWZgAciNOOd3hDiwlpeP6zQw+
uVHufCi43YfbKi8Tnr+v7cf0UJwqFOh5ks81v8go25geKnGIomsxQITyUWSSWkonByOUd/CkZGqd
6LAVK7YWTEgFmgHY28IpWeXUvzRu6n8WTW3YR8/R6U+G2D1FQ/5zNegxl84e/SumJP4002H+NLsZ
IeRqSGOeRPIe1LJHCQ7MXrEFQa+u+2M+840o2CJPqIST7TPQMb8/lejsfQFcrEGoIaQ3OSaEe0C5
asN8yEwxGsY1C0ZagwWUx/enZ++5JgRYWNu54s9JJjc+0do/b3BAmGnOlWGMt+gdtgkNb5CjHYL2
YIBtSRCKGX66oqStOr19fK9fg/XyXE65jTgmiGHBU/hmoEogoE/nB1Z82G5JUmAgemlZejLhxGav
kYqsRGyPrBa05O3l4ro/ksR2/vvbzlx1l4urVYCvaMlRafUSxItzgcNtdHl/TBT3fnUWmmXdT5HF
kLmj4zlUmwdMaA/S17N/U+xMZ9MEqSiz3McyxmYuyFEr38sskaKQv7odP1KTsilCbzRcZ7SxRmBx
Phq0mdiqIQu2CGXe2CGqJMkX+bgS+BbaR3MDEl73C4PTIH02hnvvaeos3zBFtskUSpwgdwXlaBPM
OFtlm/XcsDhopplq3KpuBps2jKpVXvx2n55KsDkHCFpEYqF5T/b8l5lCqyAKxEdnKzW56Z73Z/1j
cbprok0My32FDqJZgwYXhPPg9x+QOspCNETh6GfGVSHGVywi1yKxl82RytFbCE7S6LdjPEruy7v+
HEJZGBJe350lXg0/IE3eQ72NKPaa0YvrgBAVkKMq29MTX3H9qDX3PaiOg/qIAOwLLqtlDPdGc3J7
mFuAXIgsUVYBg/qXwGaf/wp0Cv8jHdjhqt7nfRKLtBYJaItna4QKc6wTb6xQWIgiBeTDXXwcziRY
WOJkG6LrAF50w7KtUBjZj/ve+dE42OrUbJOG9jTI+eCZh4bcDeWy18GIc/EsAKDZDR0ZC0R6nCit
W7HEIlZQGxHz5z7yR7X2jGN2KREND0QUCzBdzCwyXI4qerPdipT/vivcJ9obh1BT08hwpD8KWk9i
UNlb8rqCRLWuHHSchrlYuStRHtZXXmj2gafzJDwvJQ2mJMEK8cgB0C8SHI1m3N0zhcsUOsMsoS9P
MNGkFPlmwR2+/EJjiWHABtkEtVXXieBK+o3lc9mG0/pS2VE41nIvY4xvVPg4iu5ZjqmECkFSXe+A
UtZMt+ubc3bindMAHUdtHq3mMpDEaeowGtpRxNusxVfg6K5TajsuD7oMX9+xp9M/L1pVC8a5N3cb
kzbEOjYcXpsk+FR2r1b+ofMjgfMoFnoRjjq7nH8KbNctF4TtMrOH54dBwTMaafvzrgDijDTA7IhH
qp/1je80lMnza/2nAHr6GHbe7hiY+ZXr7Cb8k1v+wsyKax+XYrqj0F9CDnxlsld06Rd/Bv96vVNQ
Jlg08lkt7HzdXOxcWGJZcJzMt6tEK+srbbA4Mz9nFYdOA7Bs0//RpuCRifGBM7Q35ukEchPPJbOZ
JJCmwnH7RY4i9Y5eMw6PhmxeZQrt+p7y5Sdn5ifJXaBlgaW+jsUaWmLAPGyeYYQQo4GA4JzpeE/p
dQB7ZA953dkdMG9oN+OtAmLALV8R+uzxuk4j6O1qokHOm07vkPZ0BP0ekfiOwz9tGZxPFIGrDYZM
IlgJl9CFUHk9qojf3vZjRCaI35jzGbH3PzAqpTBs+zxDE1s+MuMDmWEs1rUFqUnrYXoiyUXoj8Gy
YycNLtk4JdwbNXF3qB3Zee8L6i5RelHGl9fpd1LeTE5l16/R/UsAM62xeaBEBA/b7WCfbtW2MfAj
oL2zz8L9q9yb9dJhTlTVeymYZOC9scCd8ThD9t5lMzrj/u8T2d2w0XOpZZGJOdgk/p2fDQZ34hPp
kGE3RTA8UnJWPbOx//hxXEJ+sl3OQHMH3yAMKeBHKwZzSFI4sCdFO56D9iq7IPohkCUVKwZXiHZz
aJRCEeS1kRE9kVIYfRtuNhZ/XJB5+EwAnWFRcuoJWC8KyyMYjvePm1R2caanWxi0/wPojVvzztBC
BOmLrjca0lZq3Wvq1qsBkysmR7G9wPZT0aZh38pZU1/fn3lJL/sRCipahGNEnnrJpVQgS2GwfVXv
DqGXfcu2I4SRVDA7l7KkZ01M3AFov5AWroYLRRTOWkFtmVPemkDlV/DvDC2Tv1wjPgI40EaDzLFx
++iXR+OLNRa5MMh1fZ92A9UxWg6RYk0xraEwxGIn3VlkJ9GSFr84mBwjD973eGDeFZjUPAy7mb+S
F9KlZuURLQxO5arT+/aIzNooCREy/fcF2Z4BeJovkejxBo8nIMxU92WoDfgMycy7TRDhAiXlOAgz
Lo+nTTn/Z8M7wdNu6eE0SXj0TrVggxy4UZsg0IK0itbDlNmd4B5c7uzsHQyM99T9medeQlWEog8c
E2mHczWKQ4fMD03f8lq2/t4ouRSqEorhcafXDNKo8G25ImMRb1A848n+l0pQRl4TxBRIZzNxqcpg
WWCoIcKvISftIbYwA3grpn8BHvkv94OMDnBT51ujdr1u/wwW9QSTh7X/fAgbiKGeDhAAJTOaNE6u
bpp9v0LSf/yZospbAjerKoDpQXtooBKmXK4tGw18m6Ma1qVYOib6Y0O9fLduEVbX8zJwWTbhrNYT
7VkkZtyLYFnCd9nzFMU8VYSNDQUYH8XGNmoxPRgGhFvS8illXN61fKwGr4hM2DwmAb4uPeDkIuiR
CarWjvVoXGZaqw4PfXSg7TY6X7kMBk9X5HauZj65zhBcdrUjJIIMzfPknNQ6TdLlj4zJUZokvSgP
wW0KCfVf4GEVcrfvAV98HwXopNGfizhe/eVhILhh0d6E3eo/ErwsW3Zmllq+Cp3qLo/mMPygawn1
buVpkiJQsg9yT2rDTJ2v/PvRguagdtg9KDof1wIAYK6kKI3bU1kn+MyWN9AsoYYqdTq7n9GJXeZp
ZqZY3iiwjddRG6KOSo5aAXz53trZQP6TQ78JX7qKihBTrWmfLI8ZGP6gyraEkNa8yzuSSDwasaZc
F/u2QdTmuRNHfI8eoqCBNoS/yZzM6BiaOeV1fEjv8uxNrPTpjgQtbJuCZx0Hqq6wjhL6BFPM2pYP
y5VZJL+Oi/iq+EXX4hCuThvsTqWFe1S9pCrMT7lkog0pg/uc6+NuuTyyNSQ+/Q+edMTK1zX9QRDg
dwJR7voennvodlZ9u50qRiyBdN0bM3FVVrXsXV/mOfA8t5ScEGF0gv3zbts4gP3Q14Yn+LJIP/UB
BLTkI8TGSg0xbLPBO0J2jgGqgwrj2PW2+W5Sld7xEw4czIWVnI/y2ayWodALPOscVJ34BThwXjKt
jDcNVgvx6DvoCSYJ2jZoYzci/kn0ed+SWmlX+yaDRFpJoqKQuT8NMMB4HcHLx+5l5pb22ZUsqTkQ
P1+1idtTDR2QAVs1X9vgie2qlhb/e/4UyK12M2eKPA5CI/bfZRw/+z5+Ze4nC+1Na+fvkKB3j592
MQoqvi0D0kvEI8S+16rwXJPd+row7HFJyxS/fA6MIcBHItYJ6C3zdcDQ2JuBpbT+b1xTj/q16+Jn
+vOtjwZXckFS10+I512tQBwAB94OoUFI9cTou2Zdu0KsFjgJvuUIiMS7FD4jmYFjodxG7sf6uCWO
hAF0ZbSqjZfTTYN382LsSSTYRs6L88qlSK2IgsTYbszI7w/6LzXcp8Z5/1YjG2b62JsiTcaNFdOm
+Yf6mt1IhoHl2dUtbl9xkrB/8GjCtQOB0nvYdWuE1nEjPCMNIeByodDcovvRwdE2+muqoOQ/EPHl
0qupty82jfzwGZtTQZ/IO5TuAsoK7mVtRWnU30qMEym61CG59SAqch5FrpN8UH3YqcYro4v3DKSp
wjRdIUUYrW9sbmyHHV1JbKaj1j9V0aFY5RdfT+BLanNywg09GkfwJuHxNNrCeqgufIv+AsJu7OsS
XYRJkfufgZYfiycY1R3aMDwharhRUeWYcmrwhzv6TXlg4VjyCyPdroPPphIaT7fhFr4jgl6zOwLR
PdtQTLFYXwfJREWzATmIzWCGKMI0msIlbJg5q9ht6IwpMn0xlfLufYxthp1afL6rv3qtBG/nHDdb
LJMYXa8p7sXhH5jIcWclBlqYl9nGaUGXB2UYGtIEJJQdMP0J7W2pyDVVHBdfYgjVEqwrDtMqPOnt
iBPE+2jdw5PtEz33kCnQiOoT6BkvuBBfb8kpAJsuTDFxpe4cMfCJQjjDFqQj5aHHnfEtvz6fHjhW
VLDMFDn5Fa4jZXtKX0KLH3wWwL6yRsxLyW+ZlzkStoLVJYmEXWf6xFCjeFZZQcsnTXYiMd+VKGge
VK0ib+zxhxsB0pKXYvgd0O+Kp/JxqMQUHqoj4D4KAjQJLvM4PxazsknBQr5LKclQ02Igdemi+XAE
bzZkhQNHfk0D3KZl00DgY6oiexDutp0VAb+XpgImcS5xwnPuPPMiiwfhjs0cJzaCWssVfoutABI4
2MNH6I88f/mGZK3V60/+RwxjOYK/1K9w91ybLgbP9IEHl4MAE67qvpTicLAcJBCM9YzU/XrcCExa
MZXZR3c9BEY9azOncm+q1gz+xEVOVZg/D3teufkS5OWE37M5+L8IKvMRMIa06E08Rrbd9Wa0pR6K
vRJ9N3YbS/DRTdpjswD0aVz+gbowGaXIVrI58arV2qmp+AEeRjgA7U/aUY0XwQbSWjlUTA1/vILb
e9zwNZ4BYu3G00y3WJBiNndIbiF5M400imRFLhb/jQKpKLsAM3bfOPFcGtSeyl6NxSPw/5ORA8oP
/bPtTHGzJWGbFqgV9LN6xaSgvytY3k6FBl57FwcoOm55Zu8Dx668wO3oRmAOtQvcnVwx9r4EmQ6l
f5HHyZpHbFIbRaziJd4RP9xVstaWB8pVY2Aw6P2S/w2s9skA9jApVVt/bHzyMKyMsKRbqQ3Km8iV
njsUehb9dvdGlImxMLDh373a+1ogD/Rj8xS4YuAI+CZuDGsiBQNZYqPjl6cA5TwcrRa3IYp9Pjg1
j63J0JtfgIqGGIzwgqakxSigWVSXOzvu3L06fnjOtjKBD3+8xVOtgR3bfxYK2zCcFqji8LopIFXp
ZtpwrYPx23G2JujbDmyYbZX7nqidHv2waeqJ9piyH2cEHuzxSaSwYyaSnu4fsEggNeIq0IkzYAZd
NUqr1WP+gGpbvnIxNj5bNQwhl6xP3xkBW3bcmn3W6xnS0Ey89kl9hXLM7ULMQ9fNlSU8kkjLHLQw
tx2gvxGhHANVPeeY9VV2OulP48pbvtUUD+dIFQU9aIgmgXTUHlKzB4eS8/Z1SzgPD2aq9e3604Pv
8gzDS9ixAoFCqZNeoMMUrQ+91TV2cyny5m6XkrOi0Uh+FlEPSyjs4MKPslRRieW9BuQurabuadAd
NwFmjnc3oeQ6AnTBhiy9xiT460ENaZrAfKuahl4kG+61A//ayGQuuCi2+6Yfg4SzUr7yiLcHTI0n
rNLNSc9y6yftN/Yv8xKjt1GWfd3/aHUCk4HZ22xd1ANW+YLAI0RwJOscQe11/vHmQx46v9a/pVwr
WpvP6w4kD8+r7uBU+qZ7oz0ZeCTyM1eTgKAXLXBffUbbIwJprHZHz6o27voOEbAOqXknNLeHBIui
OB5isywhan0vmMY8ianDL4t5ijzh3eZ0ykxzIMULppO5bNjiF5GW4E9JfOpbD2sKB6Ow6d//AraN
UVn9LRyBGVuRtb3IfD9aKaK5F6Z7w2pgGNAYoD3XYTYC3SXl/t07V01/F1R5cbTZTEtUqStD51kr
H20SoAgBuZWfiSLMHDgZ17zDPN43UhzfMe/3NRuua5uSRFqHWPwjQtdfM//AIlHpTApUKFbI6PkS
X7xExkuGZJSanQlWgNQ0Hnqz82DI6sHRRVMTmbZ9Gu5jVJJab6lGl/SK8YgC/u9F3lBhj38a6i9C
62fhsl+vQKE2svmeYsRpCV98roRg/2apTr4aTOVKm62OBUhAZTgzk8akSBZEOoDEkLfyKR0xe0+h
pGil0tH7qFtKS7czsYa2hxdDGz0TSkrl+HUmLv1EPsrvfDeXrgMV2pmg9mBMLlOJ3iObhFQdfs1l
H3q+vBQ6DaWUZFTg27G8PLjYiZL9jKG4+8VVahWB4lpXq330+Ctdy7044RHGoQqc5ed6dMRPVrhn
Vo3eVXfLOTbYAZQ0/KDpvsxBNC2Qb92W6xXRXGhxVfiVX/PPUB+Kc6gCTD6/qUQ6GZQ5NzYK4AmN
wg/h5dNsn28sxO/7xmIyb4tOAbBquWZjoD7BcmA6lAJGTj7kcOrMkh7BT7KuGaTfltBOLqKoknAR
+FYk1C0i+hdO+CthUhnDMJrPGtFI0LrSRN+6eITpniI1TjAwJAArhD6w4C6/igzOnjEHVrIVbEcN
TIs7l1TEPY2Srv412svL3bs8cLUH4TsNJ454be5DW9nBvM86iwWHFJXXhCOt0PiZ9/I2YocFiTcr
Q2SObUHoob0t4m/McSgHFG+93lKD6qj3nIBlXEXL0KGmRkgCEVgWuYQDqcz7zId91XuuzuVsP+pl
i0J2OJSARrLmTqcQWAJ/xOZjHokQSRFwX8Dpj4y7T8NvJYA0xiePmOvA1j7RMq7pV953hLWR33W9
implbD8kD0qc2gU0PID5Iw3knwoCoBSKOSHcv0pXsL/IARcWZGf0ghX3ZIUNmRZF2m34VobAxHZK
HvHERIMP2G6OzqkEk4ZR3Awwblw2VYNPAd4QplUpoSBLFSb263dyBWrhEOvUXbor7vRBi6scaijW
OedvCc0ZjCbx9Ds6df3/Xq7flYl8Tm0KDacnmmfGfR9QF/PbsKwCSsrXicF/sTkBD/xHgsnYHegE
4htAOSZr2X/5dl3W1BbKexpfcuRbDVB5c/A9A3kbhv8RKZX2X6U1aHS4hWWrSdTP72ONwzy8cZR0
eOWu+FZXweN6XxUgjDCpAcF6T6Q0bb1O81EDWkwREPbdujh0KFeZ58OLjsbJhHDvMY+1xlkIPaeQ
qFpaVAwXMnWWwOVVvmjfTBL8SCbZ1WQARN585zQNgQ8GuVNlPD1d/9++9v1uVkW6+MCmByqE/OMy
Xn7diTF80BtxDqjHaqqDLp108VCKfTyYZOwYzgVKrQAblRLPOCJLVoXPr+hpL8mMlBmUB48Eay3Y
CINUcSqm3pVV8ICf43UkMlnJ4FKlvnhKkSuabfpw7n3aWZCJIW71hcW38ZyyIIpcbe7YRfVvHzww
21r4dTmBgpKOplLRSBJlUw7v6p5ycXEIR1eQp+NpJKxkASe64EctShsg442FOJDOXvf7vYKzLmtb
EYSl0KbWXN6CSPVTnrb4HaerWzYJ3Lp6zEAjymNlciIcDMkyEHia6dRTYDOPPGO1gTVWwh1PMIOe
nHJVzccbsKttA5s33pSFaIbgB6rK1LRtoNysqCENMfU4gMGe4DUjmFbYrgobcrK2i0gxxluRqseQ
W/UhvMJLC0LTdeHm8h+8ndCvB6eGvGtLphgaEZAQp40Kb+lf9I8xgTOZrCAGVtOZdOI7V5go55X0
5LuRz2s62r5iN1kJV6aGi5OE6CbCZ5A60+SJWPQkL0uF9O7PejeHCcYX4Vpub9cC9DC5OFP4zqaJ
IsQH8PSBCdekAQfK+2qYU1s4lH3QWw4LYrAaWqLYII1WUkJ079dckgqRS8TXMZ/L71Y6YcXj+iws
rscfjyWqoOCG7qPigt9sW1RUiAh9JqSgzeDLbJfXuOCA+q8CwPFJVAVu4kHV6wMFf/BY7JP1wpdi
jBN47KMMIel7cWTGzO7yP7Q3TU6uBzWJe66N31K6ND142O+GttdPn5Ebe3a4B3ho2I1DrjrhVVo7
yI5+izuMT2/o5UR1ICePzhJDm449crYa0wZsnmuM5gmvIJCdCZPTkAu0DBYNmKn8e2kwmEOrL9Gd
IeXxjwrK9xF7EqRbO54aG2PCGSwmEQe05N0ZAcbsoSZbH5P2NOc7uUvQk/yt8XyO3Er7JkCEr6pq
rneWUNe4IJ6TcNxMrAN/GTY90np5lfSqcG3+UxyRDfKar8dz9vagMt4UWFOMjpjTeaJsN5cadEfB
kqilf0h2ovQVEkxZbMEpHo9VDv60Xvyb9DeiqZ03jDuCcZxR79N/vooV6+pJzE1QeU6t8OVoT3pu
H9z7YMSqirH0SwH/G04CEVu/KItG/hpJtszC/MKuoVaoIHo794YhvV7chPBG8GyJ24yatISey0rW
sk00mAZtQWom8hkIajOS1yLkLIZNwT4wEnZ5dr5gipz6n0LSkqUPv+CninkQUPKrw7tZu7AEV1Ps
vzxhvSGuUP+H2KgkZ01X/QaeLgoRpAc430Ip+UN6o7fo+MRDnRc6PJC2+QSRPr0fEg4dyIPkMj+d
gQMHTA/19DOGvg2aCxxhxL3qMlFtdESFrqX+zqv8smZ0qfNMi1CQtjh4NWEpa0MYixk3ndFdHVeW
2kZX4xGKHFypmMn3tauNq3jUKNdVC7WVW3F/kU/Til9CITNW9I19QuHiaIYrr7HCildakmMsdPGK
r04eNluShfHiRzjSarn/dj0hOM/rhJdTqr4dgjvJzk9U6qjbBXxXtiNnX1JqARy7gx3BIUdYpVMc
qlpNNZtRnPfQT7wdFmFwSDTVYQ4BfZypT9rebYYcKIH2X+jK4pnXTxBN34YWtFXhO25ciyQD8Czv
FKfi04axrQbVSH6efPy+y4QqSKGXuIubS7H3LoHsvXvdjXm5RmARpowbWBV+3mUJD0EKuFNUd2ID
UsgfMIhjGbcXzdf1koDM7fcPQ/XKOHlArvOBpMWMBkwLKBOc0jXc6j/kXVAKe2S+lmQfT6D5zBM9
8JvMzKPySqlEUbGxzr7OSg6iZij2xKbmlUz6DxtmAynW9zDxpaH2j4sIf9pSamNuIg5DM1qolqmX
BadnlwuLMuSOamv6XgWFIUf+wWvV8zcujlQlwASRD1V6ASElWPtXvryhNYd2Zr+GgqRgxiG0oBd7
2DKttC0qFlM7ikZuReVnijni29xBIQWBi+nfrFLY018/Fe7tU+4J9NJIbmmURYt/qmW46CbMlOFQ
/Fts8K4iwJElJkCDWquyKsFRVxspKRXxJd8Y9ceeetygVtuubUbLzOZovntr/4I6DWas5G4kmnZT
AfpNwhkLddUpfMaCe1IH3l9TWI0UR27GR2Uk7Whmu/sLx5Jv9zQPtCigPTfL5Pa30lrih3GuSTnd
JRwWHJIayBeH88HSAkVeRFAd3HkkZKfXQaQ+Wl4DZhw5iFb5LBk2Gvzj6jjaOWf0qgscz2IWGTty
PJNEPZuCUkbBvvsiMi7NyESAA9gFYk3i0r+zUOjCoC02Roh59J4MXI0jLYti6hpsL6pYZBA+24qv
0G5mUKUZkwDrbvOtGNBegpJNUUWoLI9ItX3xUU9Htqg+1DhXjMVBYm1mlZN+RXlS7CNk7RF2FjGL
6kzHNcnPs9ELr7mKJjJKIepENELGWSTkNUxk1hSqG705vbbjUZ32pdnkRUMWUGM1ddRFRAlXHjkB
+VfkHy/tB3i9nyiOfnSDF0uE5JWbbBsttIrj8O3xnGfFpm6GaUss8/ZDpQi0Sh7BI8Wcp7L7psEw
SwQbqfvMz4u42/L63NcPN5yie8pBsUiNLLGo09vVT6DUqINiPxE0ELj6cP5X/QEDBMwC7aJSpOUx
rxZxCY+bUeKLeQG91CotCbI9aRFI+kTjLH6WqaT8Y74UORR0929zWgUJmnCsqwEmZ2d7B49MAH+P
3J5ne0A1G9HUTnOxl4Swfeadv9bMlI0uCtJoFqVDKEmKeYz68JwOQ2iZQ4jxHx5/PSWI+vCTuIhj
oWtyfPIqzaS8SVjydLhA55CbObp9lKKosA2n5n70CXQmKLHPh2HyBuROVUJ1FTIuvVMLlvVC4qD2
V1nd0dhcBEQY2UY6decwoh0cFQFWhAhQV7asInzuVXg2kZsJIwtf3oeq4nOTl03Zw7LU1lmkNBDW
dEeRyPkxC08mBbnj/NziCqihPD4uJFZxPzqNs23+Q/xokODchqAaJgUi/4k3SB95htsraJLCRtmR
JfbASo/RuKtO/EI/WdaMdyv3o14txEdViVN41+uysKsCcTADVeguW4pnrn4y0OvpcSTyFRxqinsl
vUBuiU0j2CzjrDTUXZZhCAeUft5Lly9JMgKmN+Z5hyrLisFp8sQZdAGL8ZNc8lPmkjwW5TnTIwFM
E7QWqMFCI8qbm+G1MbBBOnZvD/l7C66HXtjwoCnK0E8EDbPaVEhttfW7O5DdrKaQayl23KGM+aTX
6hPwFIIJ1KNghAaT3Y2taNFiDZp+uQb/MX0AwvikMyXewsJB9jQgTqTOF6RmipqpmiLlN+BzZa8c
noNdcyq7iHDxCDPmKwmicCCj3FntYg88xYOXq8hBKvuhA5GnSV8S4qrdCb+C3We9y92diexvOXzH
o46owF7eopjJ3iZmtvDtr4ErTCMbh4zJFDBU17HR+o6ewL8K0ItJvLXvVoqGeEn842UpXF4tLXRH
L2zrrpcVY4dO4eUg3nXASVI31dK9fiysRdILUYGSwffny/Oq0eUBEmqhrIduQeTPxDJk/oOniuMk
+U2nWdS1c5gO7Fm6oPwl0lgwhVlv2RHKdFTR4bJRayf48Shju0oUCSvgDZOMqUEl/z6xWSZuAdPR
yyFlcVHcZ5+YopX9VCpWS4CqHQ1vgdqM0gxObPl+YVXZ/PpNm/+YFik+vtC8qgOj1koJNmM1pVvv
NLYueOg958fMFfb31zNOY+Bcy5fIPgg/c6zVHQOI4rY73WbszBlxwPPu5sBe/lw2b6OWJFBz3Ftm
8P+i9oJwrdUL4bSEN5sASIp8n3hcKUNCnaPuIwKEH8IJydoWWUHdCpiv1beDG0eFW29G5/D9du9i
k9EZ03E5eJLmS5fMK53eTj4H57LmmKJje12r82CDUhQi/xSmEdkgZa6Uvtnyi8gIFIM9USRYXRyY
BvCzdjmnxN668w+0A1Moyqe+9SSs4sGeye/eeTZKssKtf52LoDnNtsXg4NIi3WQWtiEYhxCQrjFT
YnIRlQsnw/c81lUJZltj3/E+GKCyUGVYOl7QpqMxmcM0GSUtXjCcgSgfxZjfLT0phuhXiCfSX3Aa
Kl6KiNbr2+tDq/WxbaesyCRNLtev2kJqBOdzbEITbY6rnDkJ6eyvEcXIlASDAwUaMQ7gWzdlXwhb
RX3akPNQNTEg/8ccYTkbrKn7paTO0GMP2u+Ed5vDL12LtuvfxD9GrRWFRRiSMv7evBuk8eNBUEFx
rhHEuZQt1FSmjzMmBV14Jf1yYBROMYRp9D3ZspsBbisMMUyYc8EtMYyyJX+Er2RG9PCfC3X+pcCm
AyaDIoqUzxUeCzdX4UHLEZkSs1V2+AfcQqArJM8tBJ+TSyTRxEuyl3FXZ09NEpAshqUIBgPMw2Vh
DAenOzr8cOr99dELZl5gHx8WolBGqN1J2xzIEIRfaLbKEVB0Ppxc7n9QN3ssLWXYX1sz3RWG8b0u
ecE/7SDgWhAj11JDHuQxqhTi0AUzWa86At6Yctf9JK0xVYanbNSkRwRW5bsL5NkgH/Jua7hWmI2V
jW08FCIep16OF1KZ1NnAH951gmsFwhjy3ehSdvWmNNZ2EqhQne+qSsheiN9m6l8PGxuX/HEYO9k/
L7XlRUklZIg1fPepFRZIFNp2df+CQm6RuZHWTNd8a6/K1px/VowwUHJTPawVYmSfp08f9EDSNg7h
RXAzBX3eGPLt/vcfWMJ4neY5x2jzCX/yoLMSU+kGWG4rLqNCJDqzpaVRRjnfdqyU1lcAG1eqPp/6
U2AEMau2ZEBkZ81jspov+GwFVVzdC/4GBAJotVW8xLDI8v33phMz78n9KsFW95kvoq/x6nt5ftJi
G5IV2mRQzXAOEMd8dWLpomzexDaHSaZyChQqCRovmLm091soqLkfJKI6eXRytDbpCaBvaRbivCH2
aM53r0oxxJGql9qLhwnPUm/+JXCI021GaNk1IUZS7HqOpLjn9qG9FoKfdBYPgj0i/qjAYW1X4EE8
Qrfdrkj+jr96BGNYgR+9LnTtQr6RlvhHjj0Xq1PBYfB0d6Oyi9oQ2mSfomJZ/S4QZMLOF/oRo/nw
KjakFjkH084vpVXhWTBfuZ16BqJ3Z7gz7z1rp9qrcO5zzCFbdDQ/aozSqIrGmCRtvc54AqSZ+D9f
8ndEyPItVTcNB0HFruMwSdgQOUXDnaeTs76spXd8kn3CTpQZ+uMJVKH3R6Yh/LOEzyDqUoBZSL/7
IjA3zYPxRNlRs71pq4eVXl3i7x3eA9aUeBV4dWDsEf0uLND0yf22VQXoGpTD066OjVdeeu1NIifn
tMz3guvVPgslznctzLBdP8lSiGBJSca02eA7CCP71oixZnYA76kBE5FCKRJP0xwW7QiPjvKmDX1K
1wz1kuvfuccX4b1cvCtaL8l35VE3QsfaFyfhaCof91pvDo35zc0P5H40B/yBssikUVdp0ZN4H6Ho
eqFBPJgVsiiOAVvixmNzrfREEOMsB6fao0DvvR44fwihoWzP093t6PhpJXTyferjfO1wumq0Wqea
IDMVJUiQ/ZXS4rufYYAvX/nnWGcn0A2DFJ4pMYnmGwj1Y6FhGmcsMVxslohx6DfJWc5uCCzm72wF
yi0eiq48IYqQGD5oKxuIrM/rwV7nHQv7Cn806+xP+blpb/wz9+1GAnqTtjPuzoXyNoCaolgpIUZO
cKMmftWAJ5jtVHoC13qTYK34ZBwskdyJlzi4k2SfccdzHK6eauN5CkKmH7XdmD7eSP1cVSvyHuyD
L1Wm4C5DgILeKkl+4q7ffQpIOKIICyULh6RHCBOZuFfc6pzuILugK12HjW4tTtCEgLUYHn5UiI1i
Bl+uVJwU1MXNYj0OfnjmE630L6Jh/mcLrBsSjL6M2q96foIuU2hcxm9g44Vizf3LlKwr4Sab8rei
de/R9Qc+kd2eefKHKzsCVHKYSp7iil1MQyP0ddDsZnXgAF/t90dlcNZ6QfoVPgWRLZN85ZPw1dfr
MC1InXeDlyPao9fbvlTiKTAGYE+Vl9vSljV2JNpENj6c0Epc2Vd1V4EQOTbm8e3arKh71oRaStUt
p6m5OfPZs65odEr++64hY4ankA99wnyUtoez2AP+BCJxGySZ83xr2pn+Fs6Z5RO8hfD9kAFbNVmB
tDKZLIFrwj0uK9mE6D3aksIQB9IdDPIZuRGFMJWojcI3P9bdo3yQ0IoTjOf2H5ZC5jCqkb0m/03q
MlQSyOhXtSxfrfxSsfFMGbcDgcjOloWqV9M6SWtkB+QdTkOe2lRcb3tzdrfjghmr2yDIhon/wBdw
pJaZ+Wkl45YZB3+qlVo4e2+GCsutf/EePGJkQoHmWS9a7LbYkpO2TxDv/pH1Yn4BXW4a/vAZKPut
tqjTa3PtJnnx9tIMWh9b+5Y+mW5T+fENWNFSqbJIEUCevDYUOLarQpatzYHN6uUkN5BJ/DZqzvba
ObIWbtx9DcNuNj+RbE/W4DHbgHpGTokHJInu+TOUI2eGnQOboodC3SjB5jTf8Wr95r7OjMDp0Hb6
PtRUoB95R+LehV6aufUGZp2Qr8KJJBvoEp/nROwUoPkmZu+ceAUW97OCAV2CFegCbXShHKIuIEhz
euBhNDvIXWf3RQU+PbqzabcRX6Y8t6XapEVhLKOdr/IWjizK3lw/UGNkPVO4XwA22fMM88aHwE+i
Iijn2ehAs3QamfjQii7Lea2cyRCNrNjbgtxss1yxBkIJwtS2zfSbLsWXojDBc7iQfblpC2A/Ed2+
2NQYNZVpehdvQYUI4VZVpD7ZYglUWgMYjsYTsM3R6+2EUJWJv50GB6r6oDb0XvaOf/yMK0LNhoHC
v5qGX0Ry5nF80+TRxuNGfVaRBjNY6RIgibJQ+ekzKArSuIoDKXOtli6Z08tzw+Elp3IR3s4dBAXD
JW+jBAD3X+ztYOv97Msrr5WD8D/o+IFOLeO0zbUbZy7twWKdg8sxpG+hfXPFJan39Sv/hrqXmW2t
kG0F4mhWApZL8pFlzcSXTVMexdvQomHaGy2fNGX2e6laainyB6tR11mPydvMq1QQ1GrBaCiWHuS0
+h1jJbqBLP5+cRr/CQXRxi6kAOV+SgUetMLfPuwlIFmPlzuM7HlsCtxXQVqHeBi0SjbDEGVfUbZ8
DAwMfaPmdVSeF8JPIMccrwxtdpgNxZ8e/Ks2SGwNV4vUJIzpWNGDGEl6yUk7AXhFSttFme6rwMp+
kin5JwALsgmM4OMNiT8EN6PfOXNvMQ/NTPbR+kfgv4igY78vk7s7LmTHKhFw5qsVC2/TSq19Byn4
gCN53yBEUrDrqO6hHFbv96tnN/DP+5Zpyff05M3IRvMUNwv/CGT8svb976TzllbB4B1730P3wIGF
qnlfznbB//2tXf5XAJmVMibIT5YeOyv3LgUvOB2Q/UnlTE7QG25e8YP2DMPk+LdrSDNz84rSADIa
P5ahHt1uzOJbmGEvpW0tytvNxoQur1Xkutv6cv/308dh9UPzv89xarBzzo1oVHR3zUALrUVS6pad
r36jUbz1fhyIj3jj/tS4q+5ADy9lXeB6v8KvV9luOaBV98t2d6AU4QYbDMaBNZsnd0NxLget8JlV
Zd5/fN7HthsIyA50jfiuw6GLaTpGH/GN3BTVk+JXRomSF3unn/twWGaXcK6aabS+iOPka3b6FUG7
wBxDkUo3x6wIK5BTM2VhQ66xVe6Hk1J4uIwNvAkjRcfIkAkVO6ToRC/WpEmzhSF9gzzN5n0A+ruH
GpYQ6XlIPuKlg9UcoSI83dA4FLsL9S+gcQxndno7dkG+LnHeZ0RxjRlXw+isq6q1Cz+WrIxW5tq6
faDiUUUsHhbAoFLO3mVbRlN3U1hR04uvjNUcNTm3OpYRu90iPuSBruHLr37TlGiGoPJZ8RQv+Y50
VrktaKSQbjKLsj/n+6kbVaqd5T3WoX2MR+YvNNtbI060nBWB3SnTItC4kP1qWbY2qc7x6uPdbxl5
q6bnI8hdrDBYqhPbJd8kxKMNWw0vHVG+dF+XzQyu0TX7xiGDGzXOnGg3Ap8386ODkAzczUkvs8vB
FkYP8AZLHmXnfzfhCDSDVfb/WRY+okTwT8E0KGiMI0Jruy632MLHng3BYhuIGzPJNOhNdBGvWxXF
PpAYsmPdPK4qUoXKjNNs9/AGUaTK68DQQJSEKNoPZMZXPbo+b2TSvs0dngnCVwvmQfFzI6uecKh7
1kB1fES4hETbf+GBCRSkxd7+xT+UezVa3WnNFT0z4WlEA4k/tpvucvq6ETj9ZSrvWVhQxIIUJhlH
CwLoa/4CKbjOpyrIhu/E1L/svCuuj8FI03M9fyF14vi4T1pVtTpPvO+6guZoy6Kj8C6gUFy1G10k
X2uDjkAShXbStWZDhh1viT/JddYT2Np0JjTrnCj2MSKhopR/xJOUZhTHaT61C7L8AOjWXbV1LumG
KVt6hrMmrlKI1bS6hxlcj3wFnFP6zOf4azAdEumYbeOKEmLa4nghObOW1gai+9M+mRprwke9HJeR
es+ccnTiQn0tFZuG7XHmvDYhddH7t7/xmEdXOkULZeZZHLlg0A+YAsIt0NmptMe4Yk0PG7qWafEw
+q4f4PjDopJVP2f2Rfr+4Sky5Hor/3CUWbP6VhXvjYYwt1w/kO94lo95fQkpRcDgvxCectcc6Das
SJqy4a0p4kSp6jGuENI47V8NfraCLY/8hO0GMm3rbz+LETo8O9Nkzhe/HeL9MdpM64W7V5agypnp
UVcOqlJm2Da00u7RGl5ATD2G2uiIEN/AoCc/dz3drOtQMFArJzMGd+xBBha9hQ6MEIYYtsLFavNl
NC73LBLCWXkHN1G506IN2QhH7nQwdixp7NdHvKfnKLrcQlBPIzT/1rZiKw/N77pY1P+z8pozNRP8
Uw1mOX6e6qCZN/W8zinAXe9AqvgBfq8Kxu6ckqVNTkr6u4TnrLIqrDC1wKCTzTkiLSBh/1T48GUz
0Fbf2YBtSNxYxJIKBoESIfvfLEzWi5aiGQb2A4F+LR4tLXr+FUBUuwNDUUBv/7qRPn0fuZuI8KSp
h28n3JIxgE6HEUjlWqBYxK1RQ9xJ/1q09luE2ApUQghBtipnxBhE2eG+bd6mgh6g5kqnUqitEmaB
NZ1SDxIz45uOcTwcEja9Xjhfson9nT75YZXtiR1VzWws4QBr+9lBrHE6pMCw7wMNU1XZDmKN7kfA
jvXtMh0adGMZOK/oQprKLaIx++J/1iJNZd4pqRXeJsLt0ErfrptyVoE2RqTGK9IL8fykIFyLCtlr
3Xw7XhzwyroJNzJo1HT+/suQNdsQPZCBP1L6xuLUzz3ds8Vnc8Bh/WjN4ISmScW1V4QcDUN/USIQ
fUEiLgJyr4Hcbfj973zYm3+wOPnWCK7XajFKYMMhdSGNDEbAW39Jd/2NgN+St1//KdG4UQhZKqrp
E8zoDtrvrgduNZFam2gjfUJUl9zbk8lhO5p5SKl7kpiv77uVRx18gsZ/H7A6fq2bVB0OM0nB58C5
JDQV+vyg687wE9UsJVnjqghZ7u/IlzRAxIU4Ue+OuaS1muLeH4czlkZSOXFqdShWXNvFs3w0WjZ2
9bzDFXuYRW75vAC1IRULevwgs2IJ8vc0H8LEp3CtLrS7sBZ53Gt4GDuMEi5iZzDNOdpaG4UuAP+g
ZPF53VJQhy6nwGvCnPWC/gU75ZMD7D61SyOrjtekkhbXXuQvNQmhjskbvL2Sf3QgI306WdE4UegE
zCVldFFojosFfYtILlDE5bMmjJcxl19tjUw04SjFk4J4pCl9llJXIt28O17jsaJ9KkvsMy9Zmkx8
bMZVyLEc4yk8wyvtCk4orRW/ybDTcqoTO9avrZiO5Wm+jj+L/+HWqSnpEnHqOK8W2AEQ6MmJpm3+
KCEuUzr36CdL7v5AA2fsOP4fGeP4r2gyrOFmXpWzK4TeMfFUXvyL7AD+E3C+t+RJnZPL0rzHCtPE
ux0Jn1vNDmooPmwLVd7Nq0edKJCniDZftx6VUyvdfNrUnmoTh43ZALzRNxReYvRZBFfr7EGLt80X
S+AYT9lmhbhfMhh5TxRtbZILrLRqQOzsU7opLynvUR4ut9yy5mBLTn8v8QUmBq8Wa5ytH/zjfmvM
q89bkiLgpfFgFgJ8vvs8xDjjf88tdOsJXLB8btmZ9lpPaWuxQmXiRBTGN/F1wpdAuM1ia8qOJQ0X
rSrn0y6bt0FnhOlNhesE1X2tvd/HKuNpfy+efdYBioOOaIDGhfKwWV3rwfF8agdo7USq5c4HQaEH
BCmkp2rICjSAvUTlH3f1BsO7bQZVnXsgw2xZM1oRhPBfkMGX3rUyQ+znvFl656hKbfQKswAkrHZX
XIkc/frnq4qoPTsQvFzqLew+L1yPY82uscv1ZmDN/j8Yk+oSybUcEXcki0xQjt7lXaagecDnSuZL
ixt4ta110PS665b800JC4MS3Q6WLw8W+V/ySZkqvfA3IJpoL9gefr9bL/eQe0cGp6vD+cSYWKm30
FPBLMMwK2pVb8XfxuhPImygkcN7rBxjvbmsNSBphryJuq6nFdBsYf+ZuaqP4Wi97C1e9IgoNSvfY
4/XFeLYmr0raHC4LQWyShoU78n4w6DtGzu/6QfDxvGfrWLbFtKlL/842L6acjk5w1bKtYqkmVxIn
R0K5MTqf2mrqxUWvg3xzOOsAzfXf36bzuKIaNoUBpezRGfQy3jNqBnA3kQPugzsAmxEKA0uybeCY
QF3O0wwfm3g54riRoPBJukV0x7BNbLzp2XYO1mBTA2Ldj9z7pIoRWUDQhI6FsQh/aG2EaMn2n+1x
+3fQ/dIWDHJgewN7+wCF/6BPKQFCf7APer6Al32i0eeBP2AGew5mb5uqsZu5IQmr6m8sVhhGMoYs
MWwxKH0xKSPKY1nfBWIKiYhnLLlFkWEuRXTZEW0IzDN4QZPVPVi0U8Vo0r7t86Hi+d0435RiiK4z
2T2udm7yRiqw8VxnmrJ/rJp1pvnBkCXmivbwXq1KyvFzaHXBHS7e1RMC+rR51LHc5zmEZ7MZtqDE
YjsvzhFlNJCbG2UCRtxTbh3VKHQ6t1ifcPZBqmLA6iafUjF6T0ORSQUI8t0fcOlkjhDOMccZAVfa
Jgk9zMKvsMkSepJRsCAr2OfDUIJ6+dGWmOTmgY+a7P/KemYdFVAHTSsFWtsbAEQ+dJ1EVRa1cDJd
r5brz+U8KUhn9ydN5pz282nGtGMn2SXXOVB39EdTLjcGt0C3BHPCwKXN1BznH4ozwF79Rill5Kk2
uvLI8I1y3/DIaeBK19hNsJlBoRSDXzqNv/+bXZpCrU6iz5Spfde3Vi3aByIRhfEasr0o8Ui8sqV0
6/UxeJFHRe44fmGE+JWAZnFEhqgQgLZcPHtPcFt8QqQ/eN2rTWT2LzKkwsWXMvcsroCv7rHd8cNa
6nkmf8xVQ3r8jtuRv9MvazdFM4fgK5/eJ1T801ia5jS9wSb/5lfMW9QpDOn7oXnH5fJHwFdWrzTb
k3tWidSBxLj0BU68gvONAaXmcb01DmWegnIcyhsmcmLbJhXdutwzm79bSZlKavCiRbKHr4W97daJ
5yRWNifbzYicbalvhhLieQ/OK7g3rZmaE59PKTcER+k/Fp8zHQrrgv5+XWgZA4tVMGdOCTfOyUR2
hjBGoqCSCVZTnS0VfDu1bR8QlCv5oO8A9jhxrzOy3QhfZGpX1wrDI77Oj6myT3R7r476nEBdH9xb
ykQ9FHBDEaUXleJk/4CJ0/NdLLipChucPC6ASudJ9cfc2ArGBwUDTnmxRVPzxacj5jmqwM5VvgCs
CiR0Pcvaj5gWjraum4oDmSOvYde0TOyFLqXqb9Angb/Htu8juAYWR4abv96ocwyFDzvqzWetDNnd
jAJzYTQRORyVNoJUizGvQUzw/6T9qk62AiguYqlt2zTkAeSWUW6gFqZgAteNdUJcoZBLHFq6zlXF
NCqwkbrP52z3/xgAERYem8G37Vl43gJ2aIMuIIEAEYaqV9qRnULwvAg47A33klB08JvAs1isj8DI
kZlXbocePS7dwI3bjOGxqB1/BjE6qGPV2jAUVDZpJT1R8iqqrBLwzW/VlWgjRcsjD/HIs1SXEUNw
5LBPOjmoqCpeXAZpTCn67/8Z5BaFgvMW212ByiuitbKhDLjcT5yKvZlfkieTojw9G7On7I/W02Dp
8jkdl+Vt4tqEr0MRfoQX7MAP5WGOzNyRkHYW4xB9DMR+ybwUizqUXy9TjvokXuU155AEh8ntwUeg
2npu7A5MevRCNlTfqgphlOJjgAc3P3DOClAAwPDGmV5tFK7oO90shLVE0OjM8JBSNnOTMGlLA37T
3Bfhef8GhydXPVf6e+Uz4Xt4axArgZQ9xc9t9iNtC63ol9TZ5VPw+1IeMEgFAVIwJMOCbzlcAbLn
YVno7ueEZMaMdxmgExPQSuFAwDCkkbJZt1pda00YfboDMD1wM/RM23ukjmgi4nDPjdVj0kDfPpv+
E8RAQGQK2f/pWdFZ2stt/F1JAq1HQxD2bwPqDfQ6MLigbokrBZG3tnxt8ByiMYu5yiazpP5aztn9
Y4eciuCClXJxsgYxLzYE6sKzKa3DAgQx5ycLzXPmm5inltSlYSD1P0uY+kIZ985OdCW/X+/C2j1L
Ds5rCpwBcntsjVIjrK/cd+zoi/gqX4smGIocJghs5maIb8e8kogVJcDthMmPT9+RE7AG5SVGrwHO
R6WWlqufmB9OUnBBnhFYH0qBpUPqKF+mZIFIjjlwbDr4sXlDlz5htwwdDqQiW1388QoR8oTP5oYe
NY8nw22F5Oyc4Th6wo+pCCI5meRMi4nsmxPjuZituQ7DFyddPDkj3eF11OeTC8/2SC0MaSOcdIuH
R2A0FKmz02lPjti8N1JJtcqADo+edvAL4ULq2+pViLQVJf+YU416P7UoYjfrQepECW74itwCYDBG
t3GR4q5Fvz/Vjb/o4AdZ2mbwKmHv5IEbj5Vnqf8Cis942f+O5sFDhrjpu4yZhmNa3422x2qWdhJ2
V//XXDq0UOA2/t9DWrMpsqC+9uVJE9r80UGut/LFxqAkCGoEQroNFkfmckHlu1FPm2VZk845NAY0
t/h+JlBaDPUdgoGZPFghdLDO6ohwgYJhCNZ9Koi3Xc8KSGD59rzEpftx3IQh/sHB6cnZvL5ldlM7
0CIZW9E2QV+a/VocR1HZmtdqJ74TFwmTZz21JK95qR6OKi7EPhSmo6toI+dot+5cuCsCh3baOmim
84RERs7kTku8iyDM+o6gRN45tZ0YxL9bNrA90JyQyOQbr2uqVTBwmx38ypJaiZwQwC27ePoPUOOu
qrTNwLCskutmVyhPQKRac5FgYWjKt3eHeSEsQlsJuy/MMhMbHXNY3f6YsHpFTzoe3Jo87wkzV5a3
Ob9RI0yaTBvA4Nwhn+Z0hfUzz5m+jh7AQNrjB5kwKoFRQ8fs5Z+jpCCseZdpe0GJ3c73vdU275K8
cFY6UOh2+/RIYWrURVkRyllxPJoInG8Dld4eRmkZf4ufXuK/JfPyYH27FWvkAjanG06jcgYD6nSz
jeAZl0hMuBoqRNDkTQRluAhgZq60SANneYHgxvkTal9tNMwcvMOIWHOSmIlikshdS1YAyTllmphQ
pPQwpDsbvoIdodyLtRhfNYPAm91ros5hl2iOUIGS4FZryegKY16k8rdkgCmmPbHCUWcATHVfEXWx
M1wARGB3ZXxZyGpk5WGhHr3NkruurYdtcOH+PfHGSKrK1VdDLlxofW1WjOHCgAM9xXY2FXSdWbbL
68oZvXub9HevIy6fdCuXLz0NrZUkW6y0wqpIbxbnXhXtZIrSfQZcumyUddPVSbFcEiMSmYt1A6Zv
1F22e83EAUIHqkhwh/hyQGf8Sj0DxZjbNYbVWZOSQTaFheRsb8XultsBDlh3TklnocfCn1L2LDfW
J9+yTY5hqEBDvhxXAAOmtcWs/xlR/DDnCW+u4G9ES9I6EuIPLg3byLFTHw+yJzGHFkzdTpqbI319
Eor+yvZgggnOT+u24br0OBb8sNZo+m8PcF+y9H72OTKnJoWTDLC0AYdL+wZlnUuuJumqUh0A/E7Z
mN0BwySTSKrOOsbuAH8b7WvXfI7r+dmPniGq0wpUC4K7bPuMMra5kOCcxcIs5WtaHU5NRi0tLGjv
OGRiAcm7YtvOEBiIbYNy+Lvfo6tQVlyWNvSoNta84bA2SanAH6BESkB2rTu827ndgb7WwClUuahI
DaVvFhBtGbK4MedlhBfS+mQblNCSYZtAcbca3mohNQKGceOtuw4Eh/k6ylzM43E30tVQT+Ws4+le
pNXXWK8dHWcBE9eFvtoFpYiJKFbxU1vcCxjaofAzuZMdUvK3sn6r3czlXVrUAyjvW5nds3rE4IfC
wd0oRxDyHKJRPXdJIIzwRGuR+amNvcZNh0DdS43V1GKek3aFLkwIdSQTPsBr8biITegcyBpvy48b
cCWq3iNZFlBumZxyC72d0Q2YlI4SQrLWTls77OvD/omqwOt0DBgd25rhDtZfHlr3GrXDWyfDLHyA
AFSvhlMeoHjPAQxo6UR9mLQNt/EB48z9fxwK4mlJzrWXmc7jd/CARtdXNVYeHC2E8ffBkyYdQOsN
K6km1OrQk90jW6HJ0/DX2kjN097+1RLoisBpRg8CFLnLVGLfVdCszF2Jh0uh6Q/SBjFabC2XrL0V
aaTMQw/7sVOAPXHYBd9ivFiYAoVXrDIbxNN8mmban4FqyzrdH+FwXlr9vroAW9RfWDl6T+3BMIgf
tQf77NH9BDXO9/BbENhkkH/5pV6h4lazI7A96fYe9kFC0/Psfka1p5koIjBmqlhmmylpU0H9X5Cg
rk+848cGVjrWOz4Gwh5MOESiT3g6J4/H8feMaTiwGXWHs2VOnB8Mh7+eMgcZ0+1WU5oXhoPov3eV
E4PgEwpfoSAiuqlUpl4Sb4zpv6XyG/I8Lj9pQub7XH79Xa3g+KvXX5Y+5o1NabG9ZAlIl8C2BvTu
qpFnF87CWBjiQ+tDN7ZPU0DmiUj6hejJs2kZWHiwzU24NKwzYzVZHQHNJ47FOWJVVd/60ZROPowl
GfqduTtAnSzNRCUqcfmQNmlXIz2haXVLL0Gl8IbCjPf6Fqr4EaasasSaRzly3TYDLWkEJ/NVfEKx
ggmtu3Cp5QMV/4ynKIM96oU6rnpebUOR958U4O367d8M9VgluN8uuZn6REwm1KWXLaQlEnZYKXfK
XBEduWhDpA78Q1Hcr+TCjtoIVNHrYDsRrqxJZ1OPhNww2duw2ZuYvv6pVHyrazBFl4hD0WbxQg0f
WM5Yyb9AgV2VD3bBx9szaGRX3oTDZ7q0i8Gqt78e8kaTviij2sdq9gWe60UYHniF9RUxXGxt6ONg
2K6O9RoD8mWn/AvgrX/OJ0uZ3Cxwy+vdG4/ZHojGLS56w6n9/jIwtGX1Wvx+bUQDjVXzcRvRM14y
obxF5PQfaQIeZa0s/2Hclhk9ire6HX07RxW9fkiPA6M5nhVbM9PAxwaRei24A6T/EIAsWAZ/9w3c
x5gf1kGC7lMPQsWnqKw4F2vuIVpaVMr5d0XGhjgyvhTIQSYchp4chcsFKcjzG53mSWQH6t15SWJn
fE4hZ9z8GAGCUbWzObPPSAy7BUmFStmjMHcwA3nswgwlZSHaAqRSnJHcQG/bYJpFA84ztePzJcUL
R31ij4SbTnfmFvMikIyRroMhr/Sq7RMLGzSTdCqKh4yoyDVCDzfg8o+3NdZjsyqU3I+irokTXnOB
4oCyKMpMtqAHzWEdLincLMHqXTN015nttzfb7wUHY++uLF7zjNO/4YyX1NE+RxU/Qp9rRqhnkI13
4lKbiqrDQ8xRAQzvypXce/Iqy/Ii0Ve8MucyozGeauVS2pq+h7rV7ivIpD2EwbLxpo9t0XDeN9Zf
fq5wWCu0HhHedScswmkAEU8R1+qWx2cGqmmmgkx/X0ltpva1UG1/NBab2GbKrYsSsO53hdChvpF6
3IrmAm5KI71gtgj0b4fqOZTPxD/am2owB6XbsaqqyLyJKjeuYCr4xrYQlBW4Ino+L26nD69xCAeG
E8lVETaP+U0+MKrw1I3OW+949imC5SHIU+/E5XwDtR2wuH5ijHpxLAGfPI4DWuPe/eSglpBk5tYy
eCerqfMFZ+JRI5wBBSnCwatDjgJWu1HYVGcDSRiELlhKUlSJEwhBTSmqq6IAsc2nGr68Lt39STbb
LOG6ePurdcDdjZljBotQBP2N4bW/hX1CEBfCXI/tNAM+TnxR16ks6Yhd3xx0TVcADTFMd7EU+UVP
wsSQFsiNOONTM/rfylJuI3FC+Nmi3TQi32RsFQFKYHoJI9Wz5xH5xhZF8RwE/gYq34DtlT2ocTGv
YOEJRPTWx4xDHhj/GSpE0BtjaYoLBcdU8g2jYzlDSHDOAjVkN+X4jE0sZHmPXzzp6x3T4i2ilpHP
zmAIyKR9qbKkpaWw1imJfLlUYnwis/t16LkLTrBU9e/5n9dhZavHYsL6YZqAYQoJ28jDrhJuoGC2
44B8V8bG+MyGt2ewu6kUhQxirRW5Sm/ccWKzFSACVAXuf5S+EP0OFhuk8MwB/6gNClzMylajANSm
BdmGUSSOUIkrtydzBA8YqsH7HM91FJRVwP+S5zHYpoC5zuPbUV35ijzb063DEnotHmW8irI7PHsz
vBoXjfPhct6KYyKJrWfbm/rQm8gM2rjjnidnqIwkODfYx5ToAYYAmWQPTY7xDv5vA1oQZyWnPPQi
3P+AQ4yGL/Lwk78mc4RrfixZheCuLIPF/+H4FiddjTT30lAZ90Ij+KV1CGfBEmYyjf2iUCKw1up/
ZoHswUa1Ma3Bt7k+2yiNNCylYQ5oW0r8oJSePoXu6tKjDpbagS5iMjz3WcmVxnlUU/Ce872gvSgD
jHpzewRQDkQN4wyp5WeZCQKQUHEkUwQig8LFKK98R4KvBBBbEgK2EPwnF1NAIi8Sy8aV3/IyHe+L
5EnEWlk9eWljNDgMX5bgaRlUrLQBfWeKS6t2N/b7ZCQ1WErF0u1l9C7lvSsMRBpLgTyS30XQuxqD
rULJiHDV5UyzNtR25ovKkGnYd3i2mCDb19XVfNogs1UxevH0mXwtTJZpmCbYvekJqpkwT4c8PeTY
WKPBz9chwbJ/lj19KJBLPKBtdbISJ80jOF8HWQJ4S0tE8Jn663vfoMoom1VmbCMRlqbbsyAvtTL4
1+WvadbyFmGhtHB8HMDqat0g8ynwQC7rcqdfQiX0FkVbJWvEgKvdI6zCd00GXl3BeXS4THBS0Xpn
43YfNOEy8NMdY9dQ5XP2qCn0UfMBNdqgrZBwm2iGNEhzYo1KceMne+8849Oi5+h62nh1vtxfeyUf
16WmvYb6aPlsDT6XKbTT1IhVNFcmOALa6xZnGvOQNIgms4XRBiIiVRh+LdobN1qMx6d05jtCEtCF
cWGJqa6cFUO38/A6qk6a83aQsKnOCPYAkQG8ps4P2L488x/cHnJc3bB9eRzBwdOrNTTyCLbfMprt
A/1r09aUngqXoyhSDa6GY0htzdbvztOrqYUkClzHkcvQQ3Y/mcGpdFJnkE+F6uzTqrOlAxJuSgjE
vJKUi3aczNH5nTh5ctcd13Ao3MtfYjlXlV6wteF97HD/A5KLCY+cN7Lzh3t8yBCLkkCVzNzH6vcT
MUHDgtwc1AHNIKMyGqpL2MGppcesnrlEkuDeTLXBeQsSh5okJLbEA8SZXtsvJUc7lJyPBRzvE9lx
xHJ8nVgNUCtk0StHVPstl/m+wHgPZfMrvwYLTiimWRs268tcm6CSK/WYtc71eWfs76cLlmmw00CN
rmtbzvqYunDrJvddxJszBy2RRhxBtLomKBpMatdlZQBWQSo2i6+hROEDwuQ4ciywmAg0BgMNuesd
mL61iPIKM3r9+F9huO1XzQoeU93t+ABIPcLffrowY1Z3e0H7LML1plHA38PbqnJqP3q6pcMMNVBD
SNlFgmcDQAyiALufl8TLmiU3QwA0kY2CDoLJxi1vsB5e0Q8F5tA2hkVJRMiawtQTfxgo+1w/LIna
9ZaMzuTlgyiZqq6a33Y9p6TAHfEJy/DyFyAqvtj65dMlAYpsQNh7k2dEApThSe/8ENNwFejYg4Jo
mDGycviEw6+aVvVH/fGK3PUfZFHCTw2DhYuUo/L4IZQ/BqGu7tVxNPHNkLdRdaUkcQYpeFBjjWCh
zy0d5znLljraOcWUC9YUrH+lkLoZ16dKKO/zRhPa82J6BRrY6QmaZ7Ni8anE3FAP6anbPNYJFze/
CcrZoa6EszEkHWZhaRuRGwQ5cde5ZKSpJ27gvO67X8i+qfZ9t4QtFoq918/myFXYfyClYbK10MG+
vaHCA6wlCgyELOUOd5PBjVkgPOCA8lB2xmaMVHBiRUGXA+snf+EsqRkKCYYepbxd+IGJhn2eI/XB
k0NpF/H4MVI7VjSk/lVQSG5VExA0UUndYt/JnvMFKjCVhSf1hb+9EhpRUHdJwewbkIsUVghzMiFT
gBJDAC7WO3KBsk3NNWzR+3BpktMmvdYS+1rz6BS47dI8xdhDU/VjNuhIEgamHZyNQpNzgP9kElB1
wfqHtgJzGdCaKO0fYPEqVr+FW24STToOCp2J0Ll4CaQbG23eyOPQ4QJMfXPmEBT0cCNH5K/45GUm
w6yN7sCq6/1N3lrx8L+x44XF5pGcsU27F3SH4ggtxC0pkoDBhaC5Xrt+TEKGXQAXK37Ls+sWkf7U
wYUmko6cXToGF6Js4YlnshRQ3meG22slWZENKu+VLSmSDxWTEKkMATyOy+OmEU8ZvKCF7/jALq0f
fmUw8imGe1fiahnmdHyKKjqu5BWYzzcSOHGjlHxhFuMn6ANVjuKC27Wy1PuB4IAC60Y6BjiuBFVb
e88pVKpl7683EvFd8da4dn+26vh59pasVvM3NHaB3XJD9sAkXAbZ1dXBSV8NrOSzj2oM0k8NuGW8
tsal8fP42gKCt8hoASHx1Ny++soyNfh53UJp9YgUIJ022GqnFQpF+4/zYKjdVzpn1A7XAZOGE5t+
SoOzonkBNU/hf/SH9VNV/F1uYYEBICmhPEwUj4PrPG877jf1FexQo7y71RUHJXzh95//qG0ZqtTH
z+k2xeXntVReK3gl7/fa8nJsLhUSWnSMdvaBmrKWsvpCpB6Zm/ZZWd5qqK4YmgcmaEtFGjSqOAA3
/TMxBJSwfuQPxkN8214Fa58ITCeoZmVg1MAEvQeQibn2+KfsQZrz4jHRVdnUrXXsnoXcFjASEQZW
7biOoPgxIeVQHsj7DRhS9ATRgC5NH53EzfY7D7E7i6h0HgZb2p4yXHZudvdquxGMKSIdEHCXd6sk
sDNpgfgODGIYZV7BPOgLSZZsFvIZjbN0n/SGQsTnZexb+NW2wa/0j9JEzfezhKWkHgw6yNDjGHxT
IXaY0P6dO9nMW0alCc0JOlR3NntH4ydo0gbtotaneL11sIAS/1TEdO1QbsxWfGZbLE5OSU4Og4dN
HmiSV6isz2wPMH3IfHupll+6l/MiwCFvRdtPQuVJHh39WaFg68pdi2smsYxnjVbRKwWYVrxDMmHV
QIyjHUTM3wzVV3UiUguGHHeEDseSnX2K/zD7Lz7VpRvaZEM7Dt01DFxoTkADVVd/S4iXjIGwLGxU
L8tSzJ8Aunx86QkGfagE41+ulL5SUmnLApviXEEJhk7mkNpnU0lBnK3THTaXymJgnWY3kDISZecQ
gmfRwOfaAwVqtHQB0eirUBvCmqaybsKik4hV+GrtDacuOROTzNPk7RtsIdiKcZxmNSUj9mMkoBqZ
ZLm2Y+mcbVTI5q3Mn1hzxD6Ad7Rtsl/WUVA/ZeInWx8IC5kQT7cCrOcZ6EbUb9btjKpTn3mYqm9n
0F7rm8/7UqAym5/kdj/ReozZv23xOE1DyRhzWZ6moU4Mi9Nj2k6rU5PW4Rsgt1Qdttus8q7+VhDK
wVFRcOUYOikGLT86RZLrt0mRH3VsmopII0RTNotbLjgbjVo4f1POZQlipEyKiTTWZg0x3cJMkzR+
WxlIebULKQ7ODjNvXH80AnRWH6Igo6kNXIsyC35XId2h3S9ujDvfbRK5k3tbsQxV2bQeNF06Jhue
A8wcfivEomCdjXVd49NvVec7D3IJSkz/6MFhB8t5KhU7OcGlx3G1/Aq1aejskz63g855awk1I1wr
5QiuLHf9XBPGyMWF2F4a+MmyZolcxyxDl4jFpIsfu42BvQlGMZo4fWefLapgyDkaAV+DoylNh/H6
SFw7HQyXrBDh9HM4/cJMieJx+IAk+wuFg+AJUzde5PoiM1A9y/SQvW1CmwwFf3UOivYTTv63XKVz
qRg3VAKiENGpbSZRP9OJG1ql7qBeo8INYdshl8MFMkmHz/y4MbfIz7XPHO4qQvIAhXEw+JViW3vU
SkLdisdL9WjaluB6Ud6Uyi01coaSzqgS13lEMLgkwVlg7RuN5aeRBgzCHkWTn21PlfRlyuK+iFqd
swKdJ73d2mZrtfyWjxB0wpw+ryuF9JsIazWKPSy8RAKTVP31tLhRKCG11przKsDISzuA0F/rlKz3
1rhlboxW6CQDwKnf3c3DLsN9MzuGF9UWOxdUEi9baGE2xRZ1OjpQTh7QUEfpXvGM7LuIDPzxtH2+
ibA7iC4DlAMfBLrd/6cDF166U0rlGefVpVDhPCBxAP/NeK6gJ9LxuuOaTFn3SrFL/vscbD2qbtWo
17jhHkKslRTKZQZ7+Em3pGIcjt25vce6s/6pqv1TYcQRQhk8eVv6CuzfQYah1+oTV9IQ7/EIoYOQ
EPQvw/oT2NtWqzXdvWQwxkO9Ge/YuW3ztlSnc9AoBMuRfRFi98XVoKAfM21KoePo/HFPYR4mGmsm
91DWfvB6INbEHRuDcERdPG7Ut8m7SN3BpkZgUH7OKglbtPmhiGr3XzywbnxkVlnLF+kbzlNGALhu
2udVsizCWLT1mWZRjRfnng16fK5RGA/iCrHOABFKuGEac3ECzcZsedO1yr/YJRpitCWqloRbOu3l
ill8Wj2y9Ln+9TkDmhOdRAllcO3q0y/rFqc4ydz37mXVT3HCFKJV6VNNhBiDafyRMPSsFbmZWhCe
fHmvzNFar0dZ0HCDUJ4XXjef4yreJQZhsGdVlzo5zQGFeYAQMn/1ha7HWmhXq3ktzyQCUky4mdny
g2gyoB6GNiBCn1Lv5wJGqW4HRUIXY5jTN22N8mSMIKJXSYCjtkiHqi5o2mkNT2ikbZWOM5TmQee8
g5ESgx9FAuiq1IcEK9dRrrM5V3K1oKdsfuxkWFhGlpmpSbI1QUNE259/f+y0Ck8HnzFNfAmsTGqt
7BnW1Dn91ClFNesP7zVPw159claVU75Wyq76cx/BVmMxdHPpep5HCMpBLnONSmtjaJx7QP6Qc/Iv
DXvW6yhnW1Rd95eg0uolY+2hyR8TDACakUu2Srzc0u2dyysP+9RYQ/2bwZyz0ldxqoX1d/Rudz1b
ytEmMMEzUcjnTPdl4JevvK9Wy3kC2WLEp0vt10XuevclUWGC2zib4LIFx9P3Qva0jtmG1KCIIEzC
8pPfSb5/JaI7wxISDs7m6D7A05FvMgQushX7TaI9SboOs6ATVoddnNL5klyXYFYuFXg29AGoRsSL
fTx7puAapZ2iuniO5qCACeta72DUzjA/dgYSBFuee8I+xrhYHCUGK7+LoQ+6hl4zcYKA8NR4A/wK
uW8N/ukA2HmWm+G2HLJEVQi4te/zNPEKuOHEH+eB2pbL9YmYkRV81dWJJCa/H2bFYdpwvcf6LKIN
QqTwt8KHulFXw8Tlg48rJccUq3i2II7TEO3C7lqx/yrcMmgz39Mbk/i1Bsqo7tWXeZTbTonZxhli
IFQjRNHbGy5iWABtpJ4ZG5dzKoYCWFKnrtJ536idiQKEj1kLm2ObiZYLVJbQBx/YSWVnQMT1FhOI
G+d6U0aQRB5GHskgMuMsvNNAsck2a8RB/wjjyR656DjQszsZl3sfJxwFhQECufBAvYgNhrJwVkpu
awNpu3FoHKTmrIKCkOxp/WzVMijcD5EzZrbTOM9vhDMv9lmLmE42DQPAYs2Ew+dD5rLidtDQ5IFc
FFwfy7TrppCHA9nIaOGlvkVHwqRHGro8UHlFdiNWoI8BYmWeHcarWpzWy3YDwN7I0HTDjblUkV3j
xDNIrlZNP71t3tTVfSPDt6n9LKc+xJoR6YL4OAYlI9k6qcD5qcnZr2axoJ73vzAKmE68RQStHYY1
56/XTmQXcWR3xkuUzzr6Pt53+jTi9xi0LvA975GoRfQmr6vhf3VejwapDXIYu8910LN0BlVTGbIo
7b/DxMCRtklbZ6J6+btuW1XfwtxDudbIsittZRXfSBgy6xGXix5dkNi4ItW7XE5VqNkVYxMXetod
f8OUpXv9waNf5hcoA/FfuoTtPUtEKOtV90dc7BNb0iGCTovG5VtS7kzgO07m0Jo8ZZb+a3k8v01u
0QJse/ZrPaaR+xRu/qRUdbhQCRFmqlLiKB1IKrIpGocLSBqO6GICg6NtL2umxbRXlnRzZV/Uino2
qslHNy1xKtwZxq1n+iqwaTrtSAZb5b7aMEUgybs58Pgb2a8HT1KtDIBTkO+GenSnr/KG8FbKYOzs
MlP++qZWVIs36vK2fVSvqrqesu3bQlObVzdmihLFUGke6ecf9eon+x2D8/kr0EXf1P7kYiFluGK+
q2QJnW1C7foJV2TeA8u4/ASqsjNMagJlWMCkZV0X43TMt1Eo/cHDFKuFZN0nlhTjlJ0KpKwrWZr+
uCSRyGauQ2kcuZBctpIW85bBpAIbH1XVSr5GvESBzOVZhbvOTgm3wOZpmTaNHPTB3fjWXZu2LzuK
b63Ca1Wlg61kPenDaofK3tmzaTLBsQr8RxQHO8JyE2DAO8o5LTQpPBpJ5AlJ5tuLcvuopnnCo09y
Y7pM1ZOR6Nj1+ITsIChhlFNoxjWiu090hry1yGyFNmE1yi07s4QznunX2nBsq3ivpBQXzCxjF0VB
XSAa8sPgZjjtrQJXkpkabcWwvqyOt4pG08FVT8+DyGOXWiv8dPLXxUuqC98O74NHCBkiGn8V/I8c
/ypg9dZGhssvk1EPr1Mw4wjyFIqmlWsZ+k3riqm4Foq7OieodHYOCd4CRWHJEMBeNfTB2OTQW4YF
6vYbOMLp191cCaacGiN/60CCaiM/S0D+8HbLsLnen9GuBUxOyDqziJWbERzNHMZWMpCyF8+ud2f2
tA5mjYrtsCxf375q/pLi4j34CcPmVRpPoaNtTsTJpfN/dN+wXZkfBwlUzeAsuEsOKRviCPeurwYO
VJTcKvwRNnFGgsGmSS4s6ptLclcU1z9e+DITYwbQsFQDywBHFHdjqdLVUhF+Z3wQXpmoR9baTusj
YUMZspwc7GuLduUIvRpfYg8o15NW5+o5N/UyZXKqk7jQvGUWd55a9Bm/0d5p0jVu2XuKMmJL2S6K
gY08qnJtkWYH+OcRl/HHK6l2gN1Iav13RTBYVRMNNqpjKLhp95vetZkK+bGKQZBSILHiAwwsitQ8
h4PTNcE8d+3mRfUyKfwruE7u5mj/kSbqQM+Xid1dV2H3yytpSFXL4bu+/x2uRMZA1uvAvU7t9nQ0
kiOsueMMi8ikqfzCtcGVLWJqrSRTXyJh6YbAAxqorEi2LcVPuqdBYAAzRE3BjC4pFJn1QdJLKXv1
mdvHIh1VYCbbpAqMR+g6proGNla6vyseDj3q8lV828+Q0K7I163wslDyAPNre0JE2cTPUyhl9dyF
JyeJMkBnt2vgIzbr6nIwnLJl9taZeOpponh20vROL7qjn0EYU59uDr/74TapP4BJ79KxRtwBCzyL
M1X2kUcliQWaAmIQfMZSSEK2q2nvsYTab7vVp7KTTkd5/JaiBMETdeEj8AUZSBwLnN/BXeRHwiQH
E1Nu6oEE0BkmiFLz87jtL49Yt4fasGCeaCLZKs6u6bjo1MJafI3yoNu1jpm726KS322SdlEAT58L
bZCmcjzxJ19Uil15GQBOkCEZSTG38QFKRhYo228N/M0HQu7uumXDK8roLZDRgPur9/zgzRVbZkRj
Ur3KMGZZICC3Z7Q28kKrRlxeL6NO8qHsaMcrLPhity442hkGhXvIclIybTfllSYJjW4tqnDPtDp6
T9x4aoDKwpK47ZAh1sTWIqhrqp3KeSCB7RBKYkXjXaIWHy78EDp6iBFhnzNDjlHCaWaW6w1i9Wna
qLXmUtW6EXwy66Atbt2PJAk/wuKLm1n1fqQ+IjgGgzQAoMXIjdiEtqZfkqSYshLGeXYn6qdQ7+5Y
/XpNVs2XlXSVc6+XuYMeIxEomNmbjSajOUEp06pKR0jEETg6sdk16uolJ6t2Hzf6LXO4SPPPMcMx
KUZzwb4kQqv2cxEsyi+u0w9hP9rBVaN0lXziRSYYKChGPSueQiSERz2hana8vCH9wYFDHmOCl+QN
L+Zor1Oqf0QV3esKmfI2mcQmM7vUuO4UBcL5AqrfNjJgB2qowxmHhUNYIABv+eJoRRDlv28Z20BJ
p/o/ee4e6YFnSVLSi96b0kXtmJ6DpdOGxNHDKPerEq7/zkFW8C1bcEsSYl7GpVPc/7dgSKt7sTQO
7kwHS6j0NmGzOK/mka82CTXCBK/0/YxmmMGcTnSwKmNukisNFEnQsR8/MeZ6P9bWId6FTvkJtfnI
pzU1n+yRK/+VGYNRTPyDvySaHzf/XTCeCWF6iMAPPxks/3ehKAxI/MPsr1Yu6IVHNuL6olZ7AzG2
SWBuOHEMLkqoGsSueyc+ECvcmwQUngSFoIcniT8DOjO+n3ZBGAD8EI4M82nWPpQAYh52uxJtQpp2
n2crLzLCmpou0w/7Sse2i95X1R0QV8pqbAzMIz4FXgd8DgcQbzQKBO1+AxYrwgFWazrdFTTUj9Lq
e4pfaYcqdVmcXPKhN79Q8+OPZS49VRTtfgzhBhBx7VBTd9qsItZhVD88B28ArFNtaGSPBWk9RYGk
ah/CT2z4BaHAcSuQ/8TA/ffHf3zhuFXRNgSycogQV79gAhlP4JjsUmGd1tiJD8AK+FexmzKMMC6+
JfIQUHZeMu8X1ezTa22U6udUK5+X1A5BH3UnKfjJFPl7/fGQcZfgsr/hmGyQUsdT8otqA4UHEfMl
rjIbR9X/ZQVBaW2l8jBo8PYFCXK2H1tamSZHmyg8GZ9pHjNhadId3EmLodkdi4h49P4JqOyuk1Jw
CY36j+3E14gYOGSRfbFnKOAAc2soYFJsX1HzJnGXyC9Gw7iJxG1VG5PL4q+3F+k92i7yjcCssRgF
3KfabJQB6HbaIVi3IlaSIfdIawpuQUfWDwvLv2R6jeXW+drfRC9LEEpG5D0PoehOCC89J27N28EL
iUsZhOb1MNeFqInmwlFlfL9OPaRx/RpfaOwQi6qB0d3RSQsHcaPdhaF9uxzNxUTvyzpElfa07BgZ
+u+Sy8cUKZyIirQzjOK0c5JLPJUVS1eynR+r23I5y9YhtD8o9gJjq2yh8VWL6ePPx+yzvBeUiKzW
bDLz9N5YWsk03IWeIRevq+Ysh0woQCTB2v5t1Z2WMhgOBt1bvozHKnUCRQL++s2y+54jO57g0A54
d2He0OBvrwYa2MWS9k11ce9rNKjgiSAjPaok0SSs5kdxZ7+ES7DbUfwz9T13ixga4fYbwjPMflLv
K9MriDF/ugo+NkL4JE9glfH3zHOXB1eUHlcz8chCOvnS3zeQN7LHSGsJKcDxqxcKfHgJwPRGZZOj
8fccZxcph9muxscm1HHOg4l2mlZmwbsGrPgKYbtHJoG1Wjl2H3F2sELLqJiGlz78rry/dT3x6iXJ
NRFB67EHwmt3kd1HvHNaQbajmeuA+A8S+o6GINsHXv/7wwif2kVeShPXfEee0Q6asxlVeq+ZwqEr
wEFqi/FIeXr5V8UZ0OlUp4lZSoCLBsp9KqGbJLwH+KMenncz7YJcYqHOKZWjd1Uno628w3ll/4tz
8REKoC/mtjnVaY4VOwnKl+zVkrHRGBncLpuSakVGKoWQE4phN0FE2eMT5azJNbGvfsrwCIyLF+xY
E2BS6HTIZvmY5h7k4u4lce3qonpfs0dzGuIPYmS4TcTKrlqLmuv+ywcUP+VqgkjX1FqwPN/77lnI
d1/ZU5GMm3besG3ANbZWhQVh5tL1Muyj6zXLCmCY6MmTzDyC8UHcKo2i1yOG/+rdfVJcM6fxHj/g
D+QLXC+Vao7fzxWinCYX5iR8R0ND0C+9XbLo1XADgWdw83GlF5/ghsuoxgpim/dVmuFoJ9uZtHl1
dUI0UoEXYdKBXnNGHz5fod/gh5CW428UfzXk2MjNdFAuPe/4U6tucnbKfAmD1Yh8M7EpyTE3rxwO
0VGdkP1Byrdh41YLCVt1aMGekT+6SXAX9xSAC7MpLxoClajjNnc/EDxALK5IoluxYeraGkxkp6Dq
j96d4wacWFMXDu+iBMaum0KSRgCNnwrtfXkq6ClNebjZMEkHiF6SlWJ3lB2YGDsyrg/MNhDj+rmF
JBEJ3rDjaAWtML4YtZPTRZ7Apa3dC+WScS7HA0UPwvu7YaHZEqAu+SIKCC6PqaijYC79hz3mMP4n
U5GPrmxlP1gXO9MdLtIY+9Vh32RUYmXD4QtJ+labemLwN0B7bQvncj66JWCkWbrIsItxNhlNeQai
13eZMOvQHAuoYynRC/hHYfcr0/YFoGRJC0Z6Tr0mDxPg4rNu/4QEYLmUZ1P3OkOcyWs6CtRvwi2d
gh8DLTubqU8vKAdNVWtqUy2JGsAVejp30nYog+asaplEudl5FIfeHOb4yd/oFgwSSQkgxG+X5/Bg
EZ+SyZZzlvIOi4WVjogvWAdVuJDqenKkPdvGf32kD5OzaFZsLoRqLQMF33d++lKoKtiNU6/m8IS7
GNSM2W6lARxoT8lxMk2jQeVmXsyBYwboRIiPhI022mg4WgFDREQV5QzMCSU/dQXhNxU2RYsUwp7D
TqJ+hkvayNZ6vZMn4s+GBDis6HcKnJnFtxSvbeLn6NNt4wugrsD/671PU/DR89B6xr3iOrvod4tn
/c/xDz3op0ijACdB8vsj5u1RrYLgmSg1erFXMdTyNXnFmgcgX7FfXX/0blmqELek8SABCwi2Tpt8
n3YwRwNM02q2q26zVC3FLxipuoOTxGJQ+RaEgTRWRVwH1vS2yahyf55hCllLz/in2fEBRKp4BfGg
+LNFCytue0hXxSgZjtmCToqy9eQz30uLfnUNAdSP7qzh6bl7PaOcVxf9sIrBGoMYdIoTrsGz5YEA
J4CMzwU3FSK6Q/w7YmluyqxUhncElue8zb81rIcjTlZOqLWHIe1D3uVGwJZHqwFxf0OwPxerQIYb
2u0zniXeF2RjqzsE0o6ReSF5dqH7aNAqhPoORwlMQFAq3QijR31QgP35MNMyBneQvvQMo/fUYwwm
Ff2BF9R47oo8P2zIeXdbp/yJH3q5HkS/tJIqEGzYmE7f4nntLYX/gv3OiXg+VBhY1g6gvEeu/0Wa
xLF1AqzD08r38RjOdFTd7kN64uYRqVIuNX4BdUX2R8lX4Tdt8jmA7T3HdLFNKHZlzYCZeA4xX52g
OyUICgP1yKPOstGMIXAq8ajsV4ewYiKZLIV1UTwZjmCEzFyeyBZ48kE2EkDQlpFJ4tzUmU6lcwK4
Xgj7s9ZM4ZsEFfAePRwYI4BFNnmxSf4irVMZuWJrFQfNtkONxV92yKY/S3E/r7unm1T/nF4oZ4vc
8ezZmmCluczZGnsfONJRhz6JCOsfm3hFZTyVtRO1kzbx75xsyS52dOOgYrPJThhsmdBPSuCWtEWf
r/Y8I6o9YqcoUbU4Qo9Ichd1t/XlWlTFQxL6XKjQLuazel/1mXmRoPVCzzhw1bm7GbjXoV3oQNKP
QolfoxCRQRv2hKk2nG4yeoW54UMxIrbLxbUThS9SETIK68Rop+bZsJJJ2tjE4qHLxOlPekxFy0fA
jXDyUaykQJkpjNEB3PuFNXKvF4Er8y63op8Toq1Mm20qNBt03tGJ7Zcv2fIPR5f2F/HYoNlcU601
yP1opRkE+bs41PULDxnB7jLcTL2QnVAiLGasfdiVMN5QqLvNYuDUVsy2DyBdMdDHOjIOhFRgUFOJ
T7DX13nlh8y2DJAB7D4nPF6DDVJyb6xeNLxpvy1/YHbWUflLNMbTTi4z+P3AYudK+d1uOqXhY5C/
fONLtGqWaoVQ8an/hFR26vqGxXh/sxGvNHB52Y01bzcYsoa82avsSuPIskGO4uUAA1dtbjYYTdf2
FZotqhejcA/RJZ2Mel0pXx0by+47oofEdpKpiIm9NB1+hEHQKYINsTQwJyOenKUq9mwRO4V5pfGz
fVFV3vugO4+uNL+1LlGh0qkD8W7aIdok8UpUCGaCyxLRpZquUc9aixBaX6Mlajwmt4wQpWmQaNgk
evG+JMdk3CyQOnPVWrtUmNRbS7Y1wX44c9+gFoZQgl6ueu/Oe0tlvw+AUZy85WrOY45xj/MiZQ4P
GRjuRkn3UQG2e2GCcgw0kbJjic83aoNYol9WOSEd3ec9ifmBWWK/AQjMyLd/O5UuWoQzPw+zGwZU
l7JeFrIyjrPFE4efycAnMwMD1pPekCYD3s9jssUv6EGhJvauc4sBtemzWamjITralTOna5RuxPSe
sXTxcbZu0GGTFleB/S9zOGWlgs+1CMYBXITmGU5tfcFxcHYU7+Jzh6ZN6f4V5omap9rNtWK8lK+I
uMSYaim9j0wADCpr46qQ/Cma//tKsKyskUn9zohvTeem0c1Qukwgr/9Nj4Q6hviookmiiRfIJfX1
lYM+3aDybmzd4eqN0yZLRiBqiXM1i+sGjJWAJ8WT0s5q2r+fEP9EOTINYbtODWqoxatNTvVJTgnZ
+9N5cskElDB9FWqY3FVLrP6soSCwOmcB5tMuDpLEsyws1vyfKOFbWuc+OCE6J+JcmeZUUnNw4x3z
aMCZyaQAN4RJaSA0onU9FxzNHBY8mj9CVi9fAVDTtu44Ev4W6QsX5dS/rl1eImYd8E3UxdN5oZsn
h4izADKQZgA4uE3HEulLVwPYsy1G7TOa2HyI2c+NQdAGE19eiOnCip5IN0hxSW4rS6UeWDNnudX+
Htcuc1GjQXaVaYBbNkC00C2hIkeDLrcovfSH83YDy2i1goV7f3BiY4bISBI6opHdE/n08J4IUK4n
zbdsq/z9NGXKqyqy2ECaEk0TCdcV1k4qKjonFYXXFttTq7dkQOyYRov/MiCG+eAAzte2SgR9UNHF
slp1GaKFR5B/D/Qi+TsYevg2OqjdvUNXUHgEAYhA7cAoeQ6f8BwC+wnVHw93Zi4qAT/7YZkyammi
xyiGflkuqHVC7CHSRUNqlQM35yEPusZU2de2Rj7QoXIyvFmhz+LoCOC1PgLoZ8QzjuceVm9UDOK+
g4cdbYjoTaa6Zhm5Vh1ayVp8DckLgU14RIUVvBocix2gHHWOVd2SOYDC2TCGEiJa4SQP/ZzF3pKH
NdxS/72MF3bk0JT5WnwVQtm9h8bVG59Ow3ltp1gYs62SJCpbEFmfzfqk9kFq4QoEMeqrKsNIXv4E
X/r2spn9NjyPZxnaI9QcY+9DkV8LayC6FTu/B4KCC66ATVestL33duUq9/z8T9cMWjSHInm0WPhU
MtXFmxLkyiDbowu7XbTcHlyFZe0QsIeHkeqFLa25BOO1p/Rvdsc31w918XoHh5Er3BJ5gMEOqEBB
xseAfDlN6eT+sExL3xcW6+vcXBa9BCB1SeZ4P8q8M9oKY0oIPnLUv2Mk0/lP9Cf49bPaCpt56RMj
mwq7foujXi86vCF6sOT2Q4AQI0q1F0C9IW3zmUEFZwkvXcC76pB+KqL89zdtk9Q3yuskt5JfNn5O
S7iynyF1/ApIZ6bjEAmhO/9hsV07AwbUg90QaOGV1pgsb7pi0pzEFA6+9hLThU07YPZKK60rTski
5dZKO7FO3bSbm1UbwKVsE7tCUeyK8MgO05Y7YFZkwHKFxRxiTNziTdO1pD7fDF3ijPgiMlfVgOpd
+1IfBsfWwQxtM4PBumHqBPn6EkfhQdv48T3tJ8YmI9eDeQfsT8KFmUu4yZLAOwctZQr7qk6kwv5z
vgY+aWkQWAvGZQq4maOcMxpLYcBd+xJSN/s65NQe2h6veFLSqm1C7qlb8ZovuJpqYR5b+JYc8LvS
q/9ERMvKzvu7DZk7JYw0D/eAvJIOBUmG6/BOTNJw7Z5rR432TpbzWQ/+Po5id5EvWCKSmZHXkSpb
y/Wh9L9pTKtQuykX3E+on+MFvBw/oIujeFmdhnUFSSxhVpwJPVm/YnpGPaPuarYr8Pl0j70Uwpoi
IGF/GdoL0UtotlqtBKissU6XY7XSP4DGSjJEH1ZZpnnyGM98NPVUVML6efpIm9qIPeMHbgiSA/e/
zemHutFdqE/dKlmrf6fqW7pxIoRZSEkTg/4AWqH4er7RFOj4EVqFL2Wmno2ogW3xoxCueaMVtzhP
fSsyWJyRPG95XSHSCebNbWsRMbRl9a1mMIs3F5T+VJj9DG+NP/m7zMF6nCx49IPXi3LAV/clsNgW
JdDqdudaMxiv+CMTlW6LshYmdYKe/UKfNg4yOYLHldtbaMOTjfsQojPjmlIRAS61dwN62iQBdQbi
MX7XYTPa/XU9iZCWBXH7hQv4CTGCfGx9ZQFPn2K2PUxfWvyYNiMOTikvyRX9LFZQqlNI1RM9xzzp
JdcLHGfL1/Vq3egvst+pP82DeesBDZHGeyy5XX3DgX/yP9HI8GTe3Vrphp5OqQ0OcD/vghEcFTEx
SXo14TVEkHsYF0kdi+pamOuC0fZ/Du0XmnJI0JYwAV0Idm9dyMXNQAHoEUWUTsIMrZpxeGLxYXrJ
4v2MltSEKPzHEo/W4JKHEi3HU7PdnkI7g5R83gK7OoVw4C3E6G18DMOwM4TTH34QXVaL2PniLv1L
D1JNGbLVw5GqPkey8hjNFCMMI9vtGUV/oWo40eD1egWkogYb7uxoMqwHH9YkAsvrD5+IlFA+FfQs
iWTxSVd2Bq1jDYhFHHW2x9Opb8pNDZXYQzDxr7HEFOWSTMLaoMKcOTs7Hn3Hw2/efoaMnUTagr2r
pOQ47rjLEyCuxNAgqzh/pWl1cy+Uys2McKpSNnTuFdgzBxEla3nh0KwbMjqfwLX6sz87ZK6LWEWL
t5Efv4jDXrN+GGi+i1W28OoB2PEE1Pq8oIvTQ2GhyEbJP79TBCBBQ3/e+Qe+Ie8FzLXgTUt9QqZ4
g4+7FhtoZWhqFXSo2202vaZIEZp1ybtL4v60U1kcAyDcKeAkviWE75bnIoGOU3n+4t3qb1mEM2i3
zhe8OhKyaNODRPTovWycONbuajkJRd0qfGxiDX/pR4/DcBz0aDvh+F+brZpMTMyd1L/eYOT6WVvh
/bDVBqyIRd+N2SuCDQgZUF2QdP58WPLRTbmnpX8iCIDqULlkwyZo0v9W7aGeOxU5D9jZy+ToBLAn
shqQnFpcf6RowmwzNcsW8l47dX7XAMcEkdITh2BCseawBISxCoi9vKCniwMI1qi/x76bif7Q/T1B
DRHXMJmvE8h3+Dwwsyp4RBTjmukRKdwNQG+nPTt0xwYl1wpp3NEgKst3wrb0WAV4TDLI9VI243ic
sYDOI05l0nsUFDOEQPG0qd4U1iq18c9xAP2OPQE5oerDR9QW4ZSo/VoyeZJYeprpcXH5XCDc6ThZ
cU9nm2FwaPJqr2EkKZEaNV8qxrBdiM0RtP0lfFsomxoKSnz5+SfZ940qn6uj3A2bFR2xkGZzk+rx
o/GpTHBXKHqo7EOLrNsnBrxOtebNspDvgZrJX9H03D6lnGWdOeNmjsS4BfcdbhJIASXL6xrzZ65l
BNU27CPEJz55Yvp5vP6Y+pJDmuFT4pv7hRJ2qOiljaOS3yUE3lFWj0t54mocURGN7mKS0FIFJNg6
a51v8I8E0KhMroJjXEsUNd3+Aj0ShD0hths+s8Z61BQbPV92ZyizO5C41BmOQK89qMRr7s6gT4uH
ruhivOA8Oz5tC21RIpZX44mpYZunWLHzAO0W5tCRmv8ifTkLN2iZYj4cAq1Z/Pu+E7mJFyocLF7Y
cRsRCZziAbTgvrfGFsXYw4j+aIYBsRBYCys/VhuQHh0+DmUH8AdxfwQe590jGqtV65UsclB/WTdx
XlYWR/svdyjAroQoKfYXKyT+f0pT+IDALlQaO8mapvGY1XKWu1ZZqbbyt3g+LlKmUaS/y/Tg9zxk
wMao4TACfhHKKF87AJPPWI48ro2WO2VeQChB7o1akuI7fxNfEEuxVn2acUVotE3s8GeClqDPxmsb
RXoB+ogjvtoiKmzI5bpeHL3Az07BKnmy5OphjP0CWivfEH1eKymSoZG9M29nsGYOJ7/bAUP/j+KY
8wqADypgyWOVeIXaWFwJZxtHrM7OQqau24of50K3WzNNzx7aM6eRe53WjPOD8+DyLjGIy0sDKxnJ
3ElHnw5dr0ckorWoYG5dFMDuM22Nkjd87ujJkIrogsq3vsBnwnV8uMO31Chk755Po1AxG+88RlTj
L/Jkn8o4SE6o6fSG+Nrf0O+YhzAVVmB4s7ClgXqG9/0nXN6XVxDxr6Y2bP6irvzPwxT7h0/THYno
QQZRO5IwNxf/y1r994159mUbtoygM7JIAjOwHivW/469IcZt0wAWivB0IDm/R42uz2M/pHI0t34O
gwFVrkF1Ws388zeIpEH6WNFUt7GuprIRvWgfSXnuiC/sxcFYnvIzUMNWl/WJmkHfN8Eejr3rJiVA
ptJOdeEbRmv9v8YQCajRq3d5qwTysOKdhiQ3LHUDtOBirPqwoFfr3GNbOUnszaUBwsB8zSaKCDmz
ZZbaS0s5rcgQx6nZ6BaC03gbD3nNMiCzddRCKF+Z/my87wV4+8MLr+5yZ3jyDqj7YWOW5ryTa6xv
fAyNKQR4mGmqF/fVP5epIJMWPLgo6id6Bbb/mQ+/VC9cBORei4rMxnlznHz9YspSYxi7ttLA4HN3
lYDlwYCPIYDUYojgSfd4R1ltbMYXqhcJwPJtBFiHAIfDec8Be6OnEzLiIwuwN0TQSMLVBTmhK3Z3
gz1/u2RqUopPL9mGqAtToo5yBjITsPigCevDPlUfNNEUVVMGepxzYHzxvplGRJjiz9wGwUZtGb/H
2zJ+K0UrPbfLAqw8jcWgQd9srJqIVQSu5kCLEWupjj8SzXn+5Zgx8e4u6ueuL5oirGj2eT71MRTv
+DfiACtNwXGxwbywcHjMmA6m/wxhpi46hW+r03zgQvT/6HwPHr7TwBvr4hIo1CxBa/UNFihuEcX+
gXfMkH38/A4GeE5hcyengD/frSeKYjgC4JLlD2ScN0+3V3F4QEZ1Jz+86uNSC/nqoqreS5CWiGI/
+xWZLCbKOegmDNCD64oRGV4J0tuhQGiZu/TSGEj9I19Cx92k1h6+2nKWWHxCAcbCCTZQVdfqAfdQ
z67FqOC5MxS3ipuLAbNXOkj8fcHP9CVuqeRjeUDa93JL/JJODruQJNHvHjXE0sughz5XL4xtTVuY
tGQbjCUhHyPuP6V8yeHlT8RHlS9dKoQ+AxQs2uOh2Cdrhl8wfsJwQgOb4kZoBZAGpc8raVT3p0cu
W3Sm/lGVczXiUOcvhg/rcOQgZyo/Wuo0a9Mbnuu0BnUbBPEKINV0ybkORg6Mstn6EhPPzXIasUy2
o0E5sAD2Fb/O4TEmzmDlgX61BMiYG1Ghk0bJ2D5aX5ezE0rtL+52cX+Yuklp7z+xiecw1DvNebVt
mTL6CnLaEl8Rg8t+3yPhS+f6R2d3A6rY8h0QgeKpNbhuRKfeXiQhSKu03/1T9ugDcUxDeMQkMrmj
ICrKU96JfAE7wxDrYBky/O/x+zkMH02QZjiKOw8Tj5nSwRGwpbuvgQSXM92oFQ5ezf3GCc27zE6C
GfyniyAKCyfXnIL76hF3+kVlTCgR8xDgDqA2RJwpecDXVZmV3RVw+94WbP+OO6+RXwYBY+N1L9uk
Ze7hUsrNSMYLHL3GQsZ9IWpi0okl6BYwdD+IC1yqmbZcZJUotUGQGBIQFs0TOCoLX60HYkM8Mka0
zBp3QyNItx8wkHi8JW5gdrnzDh2uItSCNikACFP3F4WtEidAgnvFyt00z0x9nYPD2pVZMtPxU0nE
PHxSBxssouO2LLrixEh6SmXnt/XhD+QNiK7HkLlOrhwRaJ1fp07x8+yOlNJXzrRJa69IkVCkQ5PK
OTPCbBSvCrtpW3PfgzbKpiHkvsSdj/nTxDe6lfukPj4O/BnYuSbe6mmguuVc2jPFjHJ4uuJWwkvl
iRBe/VdyBxVdwg2Nta9xb0il6P5XVinSSxIl9dm7pgT80hZHrRUdX44nwI+ydRkW2qO7Gt+ewdo6
DH2F8aoMQ4kjg5mkljyJ7rinuqN4AvDbBMM8W7TVGTKiHnA/OQRXhsRjSwWaClvAO6quYiMyR2ek
1uVKz0De8TIARtbfIo1HsMDiy6B9BBD/8IVDZnF5Ot4HqqtsMrN2cDIx5+RwhhgyS+2kDdHFYbZz
voti5Qf0rozPWndEaTcX40+O1STf3+lDHD1dl3QtbmBmjRpfA4V88F/M8v0o3QgakC94FSj+UGu7
XWm7qYS10UfUJ0bgK8PDsJ59vXdbU2F8LVgXu7aRcXfM14rSgdZnmuVZYCgVlJu6W1TpRHlL5nlG
kB8ZljjJaGfpvx0eKUoZgDTaiBXQiQ37lpuJEHK0rQncf3lNrMHaRCziPv9lov/7+FvdpFG0FpmR
nHe50RW/agSmNUTmTQeHWeKVAK4q0B9U3DSy0O46bP0qqlFdiRz37qLK69e2YIIcHtxaLZdPgJb/
XhDGH+9qsM3X4kgMsMIzdZHm2eZeK4wonOIl7/qeKRcGm/mLkaDYrHIw3uBi2RX0bnzlY3xS9rsg
lMe0P/Q+yzt4q2vqTIHV6NSekDgIxZpb/rDTujFSii64mvt8FTiQ1vOcPtCghZ7NDQpSPy+yLSsa
MDcuASTfCM5yvmCN/f8xcG2TmMrcmLo/TsLB+UL+YV3a4wHRbylnzIz/CJh+gmqhK0+hBQAlMqMT
ij75afAd8ojsmDqP7+xXdsuM8ctKmQVa+QU+dnCwL+qNGDBvTaK7+w3krVyomx1JAinGKfOZk3Id
se5t0Hf/mOHo2OOZO4BYdc5jc1ZDsagSioZilkmMp++Ka6LB2CSt4L7+GVtnDHJKd3F69X9Lst+e
q7+phqCOltRH099O9chJB6w7V99Xh7pBemJvNCRzRX0CGq/TKUHg5FUO50rb6oe4STvjcJMEnxlQ
LNvmGDs0ahBMvn6EQZkupb/MQ4l9yZVXtxrncdfb1KX/m6muvIG4RpS9stn/ItC833KM48sESNmx
wN35Zwe0vaaSyleWm+sNh113M0M2RS0fcQG9Ns7IjKsCrxDHjnLcvubi6Ib9qQTMlYB0j2XWua49
x0oHLQnIqN5Lw6GcLUHKb6VtlhhlQqm3dzjXIBobeo/vveXzkuMU2xTqO3uRIk7FPQ5hZQLwa4kB
y1xPBtzpthSpY5heHeBrerOKQzLcu1W4PHk7TXZVb0DhHhYXKT1+7lRWYKMOzRlCCSUz8wpcFGz6
MToU5LgA1bfHspBDfl8fKMZ8qiJbyj1GxdcXcHufXMASatiUTjzkQWA0oEVZL8t40cOrbloUXrYb
VcG+xyVoRXIdpJGuLgcEKXw6nySwyA2IqfLwsZF1tQhEavkFev6f6LaU0eeHwwTYzcImuUyRl5hj
0lk5QGpYFLPLINnjnHsttCN717uHasmntj7M3DEzd9z1m89jiJ4/Er4jmi2i2ZzsYMBEx/8R+RnU
vP/lshdOX30fSfoZsmofoOh7kldLhwBJaJ3VJBfjZjpKfXgpYLMG2dVUpUDDhJIzRBCl9WZ+CL4G
+Gm1997t8nfZTMoQMu8vk3syRGv1UCgPdHbG2X3LuFToG/ssiLMAR2ChcH3uXbOlbXMg2TBRPGxB
6Fa4ADeyUOwE/QI4EOLhIFgf2HI7dAC3NWl9mukO9YQWaX2ptrkFEM5DNtvhGj2MgFEFav6rBeYf
AiFYciSrf8TcQEus7mM7NxMZWaQ96nQ4rB8g7XsKkOa56ie/axO1hLUBAgncPRpp7SMdxHxG7GGQ
rdGwKyO73bzO6DvRXB2PzKcB+SlC5cX0uMa7lNrvSamg7aHMQxo6WhFqAttT3coYWxFwqFhsFK9P
GIqKVEt5ZHo1Raed+JETcpKb18FdlxAK8/VPVOtPxb8rHoeCBQq5JcTs3QCG7ayfZbAT0W0r8wR/
K7ruqer6AW+48m0keNtGAQtwaffbXAsrKb744vViXKOR9G2rw4EkA+f3uQlUZLrRsTOL9ZQOatSr
qRtSmPIm5+OWdPhpIUYMohDneST58gHucO/9PI5RoGDd0U3PmCiwiDhiU/hD62+NRfcPEvrVU24+
xH6+RgqignOA5Ezsx54SS5B7imOFoBJPt+c5F3tPlmxWJj4AQAZt+gUxpb4xsvmfz7VPZ6B2kFK/
pyMhbWKQ0L1QkvAoNMZaUXsIAqULTIB9kcKy0T6mRYbu5aKL0CAKwftPvFMn+3RfMMmoJmlcVaFg
wIwDRYbBkS5pq++8M7aH4bFW7Gf4R+T/b3W6sr5vrweNxYn3Qqb5VD7fOAP90W0uKdRcweYcZFn8
dTqDHRGGjJGpyknNj0jkeiO18pHteH/NHh9bSxqIf3gbwdxXlRDM24Vg0oKqVyrXNMAI4vfbymw8
/yxncHuz8AGi1GA4hVfTA5B0vXhrqvst7J1UetTAgXc6HPerydjiXWDY24lzyD7021269gZ6DHqd
xJQDBIgujOKU1f2EikY85iJqFYDdsx2jaUgK/uzCoP9jqVFGtggfCMSD7K1mHqo2zRsJx7NTSdSW
cU2LM/Fas8Qc6LNYz/+DNdm173s4scBtMwELoE0iLv+GptqkZAStgSTSNmXv6JJIHhMpMgLajJ+t
85tzwIRj+DPz89/UGjBXc4tKHR1eNgDMTIH0W9fC9XeiP/mKmnKibSjHm5uH58tA28rNqYdSmuzp
T11ioqSS8pTSTiv3iMo1VM3ePqvgxCFHUKEDVRlbhrc3uYJcwPt0rUsBNkvXxcJYPhixgtW3kdZS
Sl2IxWFOvMu91TozvT8E1gSuqSgZZ0vJahxwYW620taiXkIaWZIJQLZU2gGigtouD7mVlJnFg5IU
3fzV+h+Ddkeh1GkcwDDz9T2PfN3+qrlXMa08DPI2uCbOAmhFymi2p14R6a4zIG/jjPjXsnAM8qhq
MD6FU2lZ2BACBqpyHJSJxgNa8l4jc5vkbJmhKL4/3FRSN/AvOsiMxj002soNvmUi7mYxQK4+eiA7
wLX+i7M3QAdWx8VeubE/lzm1ogkJIelv4kMwLvDnfTqYcwSAkodihC9igz1G+yZtj14asZu2x8Ic
ASFy7UbPXP9BG1spxMwHWRagocrS7sMiLFs1YFMXC6l2CQM4bR/W+DS6fWaTbUPc+vkjIeIA8K9B
E6tPRBsG9i5Q4967Cor1l6GpeeKfo6QsB9z3nHrMA7L0f6yW0KZOo8WjOJ4xyjEwmYIv4gX5hA1k
VAcmMLl/tjgxEorvauMena8+CScG1XlUvf0GRy/BAY7hZNfIvhk7pXYAPHhroi6XEoLwrxguvwa7
L5KhUD/99LI9zMoYHgqYDPmeNe7Xl2DB1dgLFm4i5UuOWxlgE2juSLgtQ1yh9+qPdGf61UkqMGm4
vrWw/pCOmzmmUSXYKPbOGNKAgH9f+IFVbkMhq3423Eyvd195M3MET/MPQTNb+QOmNPI9BXxvcIRw
aDo3Ac0nR31hdn3RTUHv3QzWIgSzoGtoRpYIX53x4QZAq79T8+sigIUD4Uxh05jN0x/Urm6pJ2vi
B+G1tCGhxA93rfa9EryT8r72ecjBf7t5tKBzjp/h+rnaoFi/i3fCFQpiNNBkH0zFFpKuWp8n//YR
3gJchX6cA2Ms1MMZshfQZSdR0vkXoZh7o8oqvd0TZbXis0OyW6mdiD4sDv46RhDTmEC6mzDXY0Ua
o0w8qRmgLkM4tTb3RcTYOr3XfLDd5GL/1ZZGxFuPBkNT2jsTHE6AiNZUVAXgsvB6Ezc8Bz6Pb1Cb
v4I5eh8NHcZNKY/TAkkulR1unLcBtElycj7gmJgyyrPJdWtTa88iuQ6e6uTOCG64Fsgx+wQNrrO4
MNjyZciy6nXya+lFY8BkfmENgDcHqlfIllSREDkF3SepeEKkMH8C10Hy+Tp22N4sTUDJXjEsIRRD
K8csFdclIqFtqIHufrVDr+3Kin2iMvnzoI1+j533S6l7WGtUyAiA559zmh2B4PBRDcGN0ZgcVnq+
xNfUpidljKTRKfz8RcqMETzDf/7l95//8scQWtbXTyR6ZmG7hPE+aPQE6otNLfe+qC5Jrl0NUV54
ErhPqAkc/XQygGJ4QmDmSNl4xsChwdw6EfArrOAgWgcoCrGtVJDH83NS/K2y6azjmV1Dm6oCMPb9
dj8PBtirINAhq6nMWdTgF9UxoIZaELiHk6/vhrDCDZLZalLVeXJQR0mG3/c4z9BXojkKjO4dHYIi
afN23tcfNiuHk8URAMch2r/ZejLK7uyUu4uBaEHTP3/+77uCqa47gc044JhQ6h05eaOH+1htLNDS
1X/Zjzjf9Q+tWgCrpNAPmfAGzo3PRW0iEMMZEJ5TjodlHyWSC8vCjqdRmylvdlObwYXoE8DMVt1W
HLKI6GZsaMcmTRda5GkbPxIlwfrqzuStyFlBiYMaUnCydPtEXN9UZTOwdJPgG9tF5pp3VQLHeyR7
TaixJSbexNILazDNC1K3VHuJRdxJgVuh4claffrJXaoqZ1163pZwbqGZpZ2/yBYZHHeEp6ooOh2Y
b/izakKMloOGSxGRboRVFgGAYsrnTAVhXEdzdLs3WbkCdGltRw6hVJdvruSdQm18T4khotm0U6Rx
KG6nY37mdYKfqsxjAoFCvfalX1JDqxFA64uWNWhhpyI0MISKKTtWwNVQoEU6mHi4mtuSLL2xTJ40
8lZgUecM/eGCi4dfECke/HZ5Y1IVSnhs43zc3BiqVr/SiRh65ujJulmpCxdcLwAxG8NazqH/AGgK
W2kOja3VU9n7kzEgkyJuQHeyX/eALOVCCtH6cM7Z3wcY72Ae7nKV1AntHMcVY7mtdxWkOPoVEPSi
P7lzUg1/b6e4ou0wHBt+JelaA+arVXiCVrziOmG662eCL1apX+ReXpcjY5uh/V36jRYbfHTREsdC
0ytarQcX0ZDwl3Gmvfmcd+whUm4lw+2NHmNbegQ1ePzAXSY1AYAzkhgWgoXlmUZRQdwAa91AX3qj
UbIFRL3ZNSRNRSY9wAoOCS5IVvcp6jzUsQbNtATaMnaMScYNM8WU40oLr0hgge4zn+OfAI45dpmE
bbNwqgyKoDIrhe7LAjS5/hPa6on8vn0fojQMkAeSRSvNYL77hiMxqXJoTS/L22MuucNwSi3fe55p
Krpak3kwByfWlKm2s0SxKqRIVtV2cVA3IYyCbw0ABdoa8hC2T+NrsLmPmJ70sOq0h3vx9gZe6SuC
T2h4cnsVROpV6t23H776EwdiZXXuq8QT/7EwYnR21/TyFmzKRyhnHgUo3JLbYspSiAc6D/gvwJ5y
RV9UAA0X1R6e9GVEvRPf8X+UfEjFv1WOA8LnVqctD5Up4uZEeJ/+bEhCTR35GadIYa+WVC7G9sCx
r87+ve6MB8w9pWuRzggZ0ktlWkPq9anPC+J2F2rJmamv1hecGXICu/LtfU8QL/uBaRRgSIyVLkRJ
ZeNib2XISJzXeGBeI+wwNzfiMQdEu84OTaU0DsmAbZUuCVWDOfxjhW2iPHqPg2Qx+1ocq2xoBUo3
XwBYrfnz1NOMH8CHYU1SyQvClyqGpKEx5GnWlVBa9kUUKEo5yYLVfU8ym7Gs0b4RBlaKteecq3dJ
9955valwJcy+yjMt66X3CsnH0vQGCpweA/ZF/l/Whsetk8gsnkANfPqU6+OTzeon26N0uglNUxlY
UXUlgdWQFwK4YA3Bky1/J8LKX425ARzawehu57D8p6vcOqolo4BMJ6J9dIP5IliNDr3IEMl8ouij
zRHRkaONXpXKvqvzqNyQcbd7lEj7un6K/0th8xHZiSh0uMQ8uT+/CqeNpjQD4ueScSIULsGbR17o
wrxjneUw/p5RwhBvkIX0UWitQbka+14o4pG8BmHo2OYYvdVKiuE0VBGv+s+8xJzTHtogDHP43qH2
CE2WTaY4IHPGios9mUvkhfb9FXd726S24Gq0TTLrff6iLncLMF6xDb62Ubc4BP16XAsDm30fAtLs
5CvI4lUMABed5EDhfCuyTYqvLoviKd4utB/Tzh+jXqbqT/encNIP4VYUMMwNt80gr8cjGDu1oGXo
6yGOrK6mGv/OekTpy+i8z/JLxsqk/zPBUbqYUY+zuk7v9SUvQHfD6DAbjq1l/4zRsLqIhil57RLu
5nMzzh7AVbIzcJ9ouu5utXrhEnPD2W33T7b0ktQ9RdiAn0H9uxSY7i5ScDs3bDUq79GdthllesEY
Dc99+v0xekkzs/SFy37OOzazgPP+4Zv+sdmuF20UxQogs21iBw/ctzNRN2QD3qn1KDvBxq1vWa3+
ucVdBM7vZS2WaGCs28DMiYu/omkl/5hTyS2StPO1dhm1EzoOzA7dUM0oeIC3Ndvfe9PadAfX/aD3
5cxdZKwtoNhMAUUwRUIunE7+v8TsAgQZUV3IxZY3OGSCq+xH/TzHB1G7oUzKsFsH2K23A8/sHHBx
zogH3sIF0MX4GEnsaGMuQNQuuQQ926lcakbHDN2WNGvQQxkaqM+SxzSqUXS+DnJSC57M5ZLWVvXm
1aYM2W0AKz5wBbN2KbLAnetRbnT0l0mqNvPpW1Ijc4CjiQgh+1dFpaRtgEel0ySELU2iRzEu/fk3
SNr8G+5D2JTD3bvufWM7jCAkttzqdngS7QRcubXus5HToT8P0LQSIMWwKPFP6YFwm/jRMpTbkokE
6R3dXE6GWJS+UpBwECjcMA2/aN5Q5TshZeJ55PyvkWbmresx6qrX9Elc/gMvTtbXEQ6sOncdM0Hc
fKUzTVlH0UYIgst7zyITMG5isS5y1YYhjvc3AJnGTTT3K0Smrwkxc9TbAsYu5/uQQROdX31YB40K
On0N65REPNZvYiyXRgH5vMR3/1gvZ7GgJ9B8z2hpFn27Vjm6l6awJW7y5yw6MpUClheCp4ngCFAr
JN+U4ueORoILm6G9HTRrqiPtvQTCej6PpuWmW+6GChAdd/jReSpKmA9PIlHRdrwm0Fua28i9KbzS
X+7tg2OP04G2Y6m4EeDeNuwCCPxsWFlBVZet4YQhCvm4G+GtAtvo8eqh2vjaRq4DOfWzcOvlB2ls
gUElXr7GSmFIglrqIhp2kCUG+nyF3SmafVkwskyOBNQBTIl9ovhqfuuLM+hD3rMGdosV7028GyF+
UQxbz9XP/txO5SNp2dMwD4ttv0s1OszkYqsjIVH7KzljVRbk6vfwRJdS69WascTHhvyRnn/eOUn7
7vWrrFE/qZ+q5Zs5PaxdYHG6itue/icSWg4Kl4p0ZR7FnAyOkTN3AruDplhH1qfLHoz8Q5JfgrZe
xb+IFLRNWsYzBzRcbQrzjQUaMBDz0YGz+BpYVzqrd6XTS+80i2e74fgbzaJ92amED8ALdi7JgH40
Wpssk8QYc+yhyWJO6uTGNizUU22Og866biogubmb4OUVgzqPlDDOhQJtNjeYonxFGj6MYmnT0PVG
K5EZcX5dKTboKR21EZ220KZ4+AKz+BAUIALIH/g7T2AHwteydhFZq/LURZs8BuFdOp1A/iHnsThd
C6ET7zraHCbZaApg00+yjMSGuenm9UZ9lTuBQo17N0IuJ+uFwR5hk8F5NoiXOMTiPf4FR7P9NAyE
ffuOBKYrh3KttnxBqq5FAiRqLqitH8K3kqKpHJqsuZPO/zhkRV68nQA9HVpJLgbuTMy3tgpiP89t
O32LJBgQKAfknMgpk+9gQHUusni8JX5recoOun79SlA3sA9bA+rgu3/rBT8yKwUN6gldlfbTtro0
5Ztj5rWqiERBGwoFzOfOLfCMQMwn/bU1BBSa0Y11vNx7bqqNy6SVTdL+xJTK/dPZgWXUo3PNJEu4
BtIRHOcYd37X6v3Aturd1tIo64dkvG0zYOwAqktXzbfa4o+gwtgjM6zp3rz/ho0IIL2dDuzL8CPj
pzMu7L6apq7La+cMkPpVDhJh9M9povyIDvqpWS4fLp0RowumP7qrJjAeU22Xfvws9CCmCCP8Qn0D
Xim9BjuPHBWURC8vFIai5a6d4tvE0Xyck+JksT69QRh7kZMSrb8fp8QN2M5fQbluqdGHVFw17a31
0/LTd0fd/R/XA9fO7my5rlUtHMU3nL917iKLEoxogZiTrkMrGTdq3PEAS2tSlYPdGWjncUxUxxXG
lAKdgy+r6aY6HdBDmrsjxP6+9+2AAji3ka7np7tvaakppFcK7xm695kvG+oPKptPNHnGeuqo6HXI
OZ/S3HJ+IRvjTZuOnNz8P26BfqW+lj0xbBY7TDCiC87uq9fqG/ga06rjNfcDYDUE4yU/yg+DXQdm
TN5ZS7dVThEXU62gW+MXvBqm4oj+0xrp/p6pzar44uxP48SrRsavNvF+3P1u9TRg21GEkPrRX48k
bMHSaUCJ57m4v5NY1YK6UstDY2GMruT3BBcWw7+bKiaCymofzzlEsborEBBs6r+1+3P9c77cVuu0
P7YSAgOkUyuuC+3+qG0mRs0NTH50tZVESd+AZyHPpI6LtL1BXY2STpKW4+Vrs+wgqHbbJ2udws88
H9zr0ANrcbEb+oLgYab/eXoLCMqHHUPBsQYZlqpXDJKaFYdgHQcqMDGvNfaMhxkuKbewK5t3LazH
bIjQ/BG/bOGXj67BK/w6ksCwmS3pcz1UuZZHV3DLU10rh0Ahk8Gkzq2f/NvGOeVwSrJ8aNwJFnel
30Rzd16VioLvAXr0onau21ePGLbXdPccXB9QvHL7LaCg86ZwhewmK03sFs5iJ7M3JODH+5M8ng7g
cLR2rm+YaEY1sLn15XAU6cfUZM8uBS9b5qZnEKc6nd3XmbWjYVFaFXgd+VtaJ7nfhUpo0a+Bl8mT
e1+l7vnMW+TF3uY8FEKcSjGDQJ8qIAVWa9gYfrIEZeCCaU1Weay+L8vp3QSR7zoOfA7mwiv/WkUA
o8wYjz9b+SNsXVtdMew/kEGmOmXOaTTi4WIv8MV0mzG9uRNMWAFvX/c/+c8zLxm0vJv/wVHa2X7k
LgXxpIfohXakQCweUmAv5XDCTR/i17Iz3JPRdw9DRe0HqKXYkgDqZUxuHKGQKByM3TZVW3fmNq+U
WmWrw5JC7ylZot0P2v49wjTyVOva1c/6FzzPEAiNb8p/wBa8RVxBViJQIeo5npUFLRbKuG6ja5tW
BcyrePRn6Z1+YqZjhjXKvqaaEcHZXDEQiETEnJv/0ueNfTVSCe2r3yaKQ1ZlXeNGuZ1TGYznCVbZ
/WdfHgECJVYL4Sja/ZIMojnOSqjne68vob8tsjYmUixpKT1UkBUdPb5lcDFgIYNApQXXAv1rB4+5
MV8q6OxE2I/KsIbkvQecNGWRl62utsb/AWt7rp79ZbtkJhcr12HY5AKenxyV2B7xZM/kjEsOs2Pb
Rzf+UtQiOPrTY9tc5+vgYjSy4jLW6Bg+zuhxFBoHcn5eojFMBKctITCngZfyvPq4rA9+5Q2M7Vmi
zamx2TGgJD34QWS0dR8aVZ+Rzc1ktcBEcDXcIEdC8ZF5MVw3xXpK+cqmRX0z16x+6w+Opf1Gqapa
CMg9wB8K0i2RY2nb4s0mHy1Z2Ep6cs0/VyHIyY6HKMMeWYYAEziGn+j2x3G+psEs8eLqbvx0QcDF
+lUeNzsd3ZVZoisHXEUb5aDbsmzeyc0XQvwhAAxts6lYF9IiBXmWxijTRCCdZd79u76UWNAkL2zH
39B9GOWomb+nRavmvUSi6/g3xLEx9j2uTQRiAatTi1mdoxwncnu/gY9nR0ywt6H5HW4I7CjxH1Xu
R76mDBO362TkjgUAVrhaVuOrqawQ3TPio5Q/iO10f+DYM/RDEJQhVzq5dYx0J77RyyMnnQnYxbIj
dwf1w0QPBtB+uyxms8gdxmCdWm7DKjMmXkT5Qf4UN0DAjf+Me63TWcYOYxXpQ1hDHBkbRc3jsmu0
UGgFtbRqnFJEAtrw5nbArWBwOlaC5yPYtRlUNZxtRSKDbaXssncWRWh1o0DF2gDoucfNE7tBcXJP
aD0YRockW6mYKqIxqQ0aLXi83pP3O3HhTu3PdkSG/t/aLp4cCF1bDVhWmb3A75g+TNV5+GcZ3lBg
aYq6zgN2wSmYjbiQjE9zosP7DqK7Cnwx54j6KJwuW0DRuijsOhjGukgA2ENTV63ZZxexiIUl0g9X
d5eOADVhp6gh65CDf2v6b6k4wl+hdnkX3+IFKmQ3kbePbOMqmbwGElCPS4ZMpeV0AttM2mLcSIYl
zG2ZR9O7Rt5AAO5t1S5yV8mRQIevvWbl4u9xM/1cmbzPULdB29CLFVc/xD1qXcWgYuHuCqp5YiDT
vFmRyg9MMnZVWsNKqP0ja+fw81dgxz7rBNhBccwpkScaVR5caQPuqcUmIl1w6hCaOayHMOT97/yc
9I9WTwQKfFKyV1q858bIZ80ORpBYHRxffr9ueTEPitHsDnfi2WgsnKm7wePPMf1bXgxb6qPuZ75K
tqIlv3v7LnexS666Cub8446gMkffgfUOxxNKiysxKRHYC1Rn4W6RV+oktxr+JzxlQ9vwwSfhhZGR
eo8wrI4/BZUeXLu889w4JSikxTA8MrzfmIPHHznwQd8tsMtcSStwQ3VubPCGMXT/H0oQy3KyC84R
bZw1aAOUIAJfNpJTC0JKnaCCYm61QsRXZVMtKypN9o9LTpkm73DNUcOZiT7DkENNMuWBtg/HBDId
fimcs+cET8XIfDC8EOrXrjgzhDYlRzxCm4ERCwcTcBXByBcptTZlA3TOnx/q1+p6iX14tbN6YBWe
f/9gUMxMS5U88QrijxX9V/64839oEz8DAQsfZCOSC509hJXa6HYUGOoqP5fJ8fmbKSzJLCQtIUmq
SV3AzdDHW8e4IXH8G5zWAdYJqzHqUHx3p9SvyG3BwDKizV/hgNp9b9MYummGDId7sT20QMetSrQ3
6IVRdCd6lbTu3XFLOBwynfWy/SeqylyWR3vJB5a8fVoy2YvVmFn3la0x6h6FUfO70SYANtiwTaxl
iKW1/hO2Wp6aNoqRy5gryrWHU6NhppaBQsX4xH9bZpl8ijmgK0MXtFhf3WAl9gDSAtWKw5uYsVez
/y0mDWkodP1/vEN+Cr8UNyr+/d/naw+LqcJpV8H/0MI181bMI2EbQJVa6bfVPvcqIVVAiIgUpgqh
g+ZyGbuL7/4ywJ0g08jXxInxMuDib+R4RGcwzp3xXXGfG4Izc0cenb7A+NQQKySTgiR8B3RBeaT7
mSZ+Itpn1zGeTtIbShPVK1c8q3WR8PX/y0r6V6p9iHq/34j8BkyvGP/hi1pObZIJVINQdkuEvbNr
3x9P0/B42i0963kv8+ZdqFHhV0Te1cC5LWwH3OKho3G/uaObGHzqJehpRG60HpPN5MXx5It/EBzf
lPtUc6iLnWWRrABYgrVHiRrVIGaJGj0LiaVHzutYSsJRp1v60UYLi3DUACb2qoQwxu8Z1YmxKLi2
NYbBntfEkmKcyRYbaXxj6PSCPgAQrEibGydshLuVoddlmbYtN2qYRABXNwPC9ZzdFiAXw21pO3Yt
ZlaBdIijj3kbc1hqAGozdfdUCfELQGJXs2f8C09SOhMUXodD6zFHz3GmpLyEw9ZJ4sWkeQkEFGeV
wx7ArRMHbgXv8GXVmgvZo0gqDvnhDfGaG30Xp8UblGP2BTccX+qTV50HpMh1SoNflIrvuIR9Im3G
T+d7chQKl5We/aVRimatTF39IQwRVVKXw4QZi5JikerpkfuebvRZfe2mfckwhhkDl3FKw+50hrv9
C5Q0q/OOCZYantxxeCAlcu0q5RPkl8r4fjYQEUutQo7GzX2xdkeV/RqfIadP/HoByoNBFJnmjL41
ythaKDcnIf61onxXnOJp+j112GMC2q9JMn8AxG0jYoOdmecbBxZ9zDdtCrzD6PvGJTf8nmjXwHQy
opsaHpSwM5c6iZZba1plnhbXoqZ/bryyQDLfGy1Hh4eb0T/LVIlThc4bNat+no8m27pU63MHEMJB
74mPg4Nl67a27u4AKeUnnTicJJ+KBUuBwtQZ7fvHO7I2sG7+3PzRsbgCoHAMdJghRDSt+LWgyzOH
eFqv5bPBjXImOqUij4hdT6m+DTDK7D5G8GD18cPa+XZuj6oK2M0U2W6nGU6hrhibFMl/VI/2Sz6E
BuMP0d2KAkbb8FirWCAfEikB7YXTq2l1aZ0ypHjrV893eaF1WJPnC+zW0N3nWtPO6kuW8afk2RJw
zejmpET1rnSAkjEvId7kuy0YYi/LFu9CL6hs+R7LfmiQK8RKNJ8KoRvTQOp3UCGt3Pi8BXfQhVF2
YjaLYKfil0B536Rr0+B/uHCX/c8L1rRD3jBuUYo61EP+mqEq06zOoA7T1kKUYgwL/4/hHMtUpQ36
uD3gNAsaJ5V9coCCc7uXWRwC6ACOYDayDr6Y0lyQW/3qcWtjdRG+Q/Wmlzn4zL8iVmiKiLANF772
q0qYCeg3ODO9Xqg0XCLEwIoA+yxu8WeaTzWlrYD0YwNRFL+9TGQGeRx9kiHdQWWDBrsjye0wpsrn
sFnaZdbIX305fjiA8qXbNP+Ycc3qu3e3AAo+w+COYVsjqOjauzJd/cRDAKfOIePFpHy+E0VRDQXa
/l7/PjNnrDNwopoOBePoPl+3ivkTg8uJ5xX2QNOe0jTRiuG/P9FFXVA0CeZZ3hisEUrE6FKXXeFs
FyyLvpsORSa8sEl+PKtq9EFISGWY0jnMD3fdjt5CTHKNiM/icpFiNpUAWLwOyl50IFO9qR4ix5cR
6TGtsvpTSl4jPIjxwDg6HUKU4QyBmKSjgbBlITvjkRgzpI+sgqGrRUrZw6p2RAp1pAsQJZMbPQ8N
ffLP+d63VchuYTMDcoEZMv3WKmQQJD67z5iEzq+HPxnkdhqWfQlSo6naCq+ZCUEQpm8//CBcAoQ1
aK0hadGbMLfaUdlG+6GoOD1JNq7S3SrUHql5voL3JyfK3S04/Kakmuz3oBV2qVn7kgmpV9eflSL+
aST+wYDL50QMUjFwtg8k3jSeWfNhZoBLCWYCuPB1GYwDY/0cMUjm7qZa2v/LVSp2VtKNL7rJ7czj
gKpecBzRBLBcG9izWEyt4yapg5Gj+6izaX5RDjNcjYNsgjMizE2wypQr9Sct/FGK1zm8pdIAtbn5
nTElp2TQT4a8FKEO6jm0ClBJaaWpLctTbSu1s4AeY5WaWFOiCnUnrmNO9qzapsXYuSBUlg/pYNNr
ujm2Sav4tF5jdPLyb1W7w64wW690A0UZx9vc+nwr1tN8PzUoJhgUM8J0kI9YkwyGLfiS3UN6jMvC
AZyu0hC4KlIIWStjbJ+ZybgZnr30dkRCb265DaGihJwVei3duo2I/ySwF73a/lWH5JDJB3u0nPni
l6wKdJ2m8OaArtuatreXY4PStZWUUhJhpeC+XDIQF4CQcvP/vM6fZW8g480W9Qry6h3k6FiPvO5p
v/Ej+QXU6gz1VWjmlo6n05APqHu3fcY2pAabw+7rGxAuTbyPH+GLuOur/wu6RvjLklZrbPI1yWN6
qhubAnxnScNPLU0YrqSj98GJxQ7ZccaTgi71MNGrxk13GzlHt8X2/oPLrBxZJQnKg7vIzaqGMkvt
M9pLsm/h1qQEw29Kl8M587wF3o6mysl1im1rIbtdAvIvkzRKifS42VBc1/rYSu9anpg67wZB6HSz
dhKbA1JqV3+KxCKjRszCGPcnWDSrFKz3jVwdA0vV1ooYGh2haPbYBqqWgREUL2LRYnYCmJp81Ivo
U9F6yYBHd/ikGgt3Wl5BcM6m1uLhLpx+gkXtEk9Qc5h4k2xQ3jE6NqmwekgStToPSw5jTbsiLctY
3tczLdczyHHSUz/Os/a2uSR/v9bf50spVZTsiu5eb3PaRT6ifWNrsk/EPiIdfrTfcVHs91xZhmrV
3M5nfFzj/5rMAQFRLITNOXZ7fdduD+6jgEbU1dwoyZMZQJo/RevdgSsBC4NFnJGdBDs5FgR6BY+Z
wDnrgAenn6XONSmmCco2D+oJaUPylDu2g6nYlwzI4OToibmYKDSnBIAfshpoh+afYGXS3q48qCB1
a9GDlDLfDqcLm7puyQZeeq6pGI0lGyJV3fEsE7SRJJ0X9zcbArDKNsoMOaBPlAaNXqtuLuwuxgFq
gV/sEnbthJPIlScsm+1AlTLXn1jkVo/nT6R1NjaFGBnC6KMKE0oKWlqNrH1RjG9ZYXqDOUWLL+EP
DcYYe4Di/Zxo834LUTfPpg+3pmRmDqvLI0zeFtZGKYmBs3CjtKhQNbH5JIA9pqvcbWgzMJ2+hOV4
ivPVkEdkZy2pZBOGRksnRcthSta+HBgCs+YPqFUKIjRuUqX2MoTLc0Du0gsg81yE7WZHsuwE/diw
ugvRPwyNaPvyq35zVJwkyZt5RN0soreob9jllhcHmQCQknGhQEg0tsaTtlMi3kL+pE6hokPq6m7E
XUu705y7eRLqmg9Gj4cnI5oFJLKGlbbWtfTBrwdM6z1iAoJElhzvDmHTEhCUT08F/SzC0TYbUawJ
5IuPyQYfkub9cOKh/8iyiPxlDohK/uV/PlSM6wqDusuOWu9+uLkQxTtCpza/SsTy0xfjyK08UoNJ
gPYmki9yYwPNZSEHSuTKCeMVEjopctidbCx8nk1ye65xTUadDqiZb1YPTT/npVKyY0xc6SzwrdJm
UZVV5XgAZ5Vjdw7V3OLGTnoyWujgzE2LfEDV56cbQgFz53A6oyoHnjBCVbd1Tv/r7ZDhnqz/3DME
zk+pTh3w/gdhcgATl+F8GoGVzALFTKKNHFWcxAORPNxDH7D35T2L9jaybsWSGg2qb8fYApk+f4UQ
piULtv6msQW9WbpqyQhLGsR6DlF0YHHbsfAsSkaVSv0janhFI8Ez5b1HRAA26a64w+QW8wnZNtja
afdDlztsSh1k11gzzZUI/v4GOo7DwHZG+RA+TZFiZv/BXNymwBgf+/970RQgqBvf4HFvI+ztfYqB
derIphMTA7fEB7s9qPqpl6sxk7SoN3xqVEjwMOOJ+uwrdChsBs9lzdUbhRb+C8WEuKeGWhVMUlLW
QXs8wSpKXUnOfHrHN1WVBzXnTa13f9emS3sZYhALgdbrAnkHm25l5BRWTMQxZtmEOMt62REmi16r
hYOYcMFfK2jV9srfMKRbpiVLu5ppnnfCdcO09YMRcgA6/WZGfQP9GmnZQL3cKpj/iPfQt5X9e5+J
bitXMEKnP6TkkmAjfntrkOmxzrpFmqL/tn90TGeRdXhw0oeeVi+BGsj9dsr/RqjPTDvKufOPURV5
LfCfhkD6ApKGW4uYNZSPPDwsuXDnjF+96lT8lIzYRDn/8WmILKWlLnQq6BJaSmVlvzONYp8y4H6j
M0iiTjuB0MHu1XBei+xySVQoC7Z2ClWmOxSJhow7nvA6h16u4cTVXYQmWtJsdJhWm23sQL3mwB16
HVVfY/6sE5DBmo79oNHfeU4vMgBuaSnNkLx63/U/X3I81BqfpwClcVSTTrIBHWKlX5HZ4cZeW6oK
x8EEGx0oyJoLgLXDCggvbczeFWsY59TtKxa2Y8KpmaDBdeZsx6aCjyj4EnflSsQkNLRO8CSSdhpc
70M3omwId8+sbVUfKUys8BCpYBQRgFYrT9L8jXpsD+dymPUjNc1jpbKB1ITt9eG4kICjw2udQf5F
SgZKNe+FQR39qWc3Bv8hOH6KHDZtN315lq4slXn7QBYXLFzNN/b7vpGWnXP4lRrZMg37l2nzB0IP
laJjgslRvjLfpKMIy0ZnwQeEUTd28iYwSxiFr2U4m7UiKOEGiylPDJlFxJ2/boSXabaWfKKalDOh
qVAeUZlIvlN6t/lKlnhD2d1ihINZb8uaihcFLND/WmWtxfAWHBv2t7H4xxAupspdYVmsBod8MZNP
2Km8YoH2MQH2V7o1yAmtX9qfgx5Wuo4ViYHOvHCo0eKym9GeoKZfsaAY70NP7T8EbmZiNqngbGwD
3ZAbTU/v8NCzSUbz+q774VUS4PzuZi+MJ2yrUS2vddxxSd17qRxX9FAwFh99IpMte9kC+PqrohAh
J4M0TP3c9YkLdhdeqXHtQvc+L1yzHJruJfx5kqGO3ZKFd9u/avqygVjhU6wpbe77paKPHvFuJSwQ
jHJUT0qzvRPncVGztG572hXn9cCMGSbsYalEPr1K0IySOWdA4O/sFxdq1SpJDCcrm0z5GtCVQ5lk
s0aJ1w60MvD16/jeMSKymfdsTla7jU0eX5zAmdXA3owUwmdyBtr9H4WKBYoRJwixQmpI9fZZSbgQ
Qx5PE05AZ59UQWTwEIrHJeZA7iOAnGIgB54/BI//hyGO+dRj7L5y6BaKjGT3Nt9i0tgwutbcffbs
5ScblRTf+KZQm95Te+h6MQTa78ijknceuTXX/fhQgyCSkjT9yr3hjK3kBDucbhXZ8L/Ew9fopcX9
xbn9205pK4+U/U4D05qoCEfdN96JKahTU/TJo+HnB7R3u2Ksc7j94OiiR3cfXMSr8SSkUnbdNnAF
2rt+mc9k4jllDEuYYClHYDntiDyMws4YYXABvRsTGCOs7QnzPXv085jgGWgfh/7NvwVZJ9EvA/Pv
0OEGeaB2XQ7DkarViG3213t5DmvTGAHUnc7hLQH63XQ0R8ml3hDMdmtCzgFQ8KPwhT6pZiVlEpdw
cEMD55LLDqekTdN0R29UfNaVpDoo+pye966OsFSHElia5ETTdJpzR9CkiAVkc+5gbfQLlfNUmuXe
txir+URtqcGFgCUICTtLKdHum/odcYi8IMgkcihZLv3d0prjBObXU0AQ6aANvaTq2IYbMFabyLud
t5XVRuHy9mkyDH24Lodk5gOpKJq7rbxGuXZMo1/YSNbXUiHxNMhtq8Tr8AVOd8dGtShmGNKrue0B
tjxDdO1y8WDj2YymoTWAIKbynQSrAYr115CcdFpjq9WTAPOyxizPnchkpdjY/j0hlzdAYu4cesQh
8kDWp7TqxuNR5s7N4YqOmEbgm/QsiC3RrfJ6AyAfdB9qG9yPgipdaLjPfngc8v2DKbd8nXHb3Teg
+r0KHRj7Yzcm9UPtfuYbtOLAbqVacIW2/5AhYdK9S6iCpxl3s+WTvAe6GE0vMmxBzsobDKXj7FsZ
XCVVRujHqrwtsWKoZX/ACkWjIP2AdDLTkMoHqxX+ne0L6QYP8k0d+Th3d+eQ8domPsR9ZJdP141u
MIH50MSoDtaJULXeWmLoIhOiOgRRhw2rYaYVy86++r/jeYBP4voYccSRmaPVNDHOqNgT113bMN0H
/8urnu0ThjZ1PfPr1vXXf1bZfF7MzQ6mRsrZE+Zc41UGRENpLYyimSyBcAcz0QiURDYv5VDRXYBw
oMzfLNfwWqSMwEG6elgWYOC0cYLOGpSBOs9Xu6LimR4fc/vob/gqvQ896NKv9xrHQb9FvF1xUjul
VfNhkU5gV3PgnaWW/5CnZCGMnmAzzM3nwIrztSjdGYtH9nTlR1URT8O6FHpD6wOV11Gflyavvv07
jIKG9z4v6svbGXIbVGlstRj+MECCb3egir+Mt/KPqcewWCsarEd9y7/nF54E5mcEavou42614njG
m2dxrJGZWnLpKCYhA7fS9Ix/A302IbyNd2me2hellGNKbCduWRQE/ut65sk+R3ba1SS1OJswQmbs
eti1U16pfDXVVT8Kq0VbPXEaELn6JFGL/Q9NL2KR6gMf4wfO9aw3YwG7Aa2Wt99Uax4n/c89OAy4
GzIlULdB7pH8bUp7rxaPQcBpiXzUSrgFPT5qlPzhNSzKbOVkc0yzWx1al8gzsKCJdZlILUHLhafz
n5bAc+L1x41cVHbXSkUGc8cMkxyx5pQuKtKCTrrklzuoHfjusQOfAVkxLfs8tbUxIEPbYFR80YAr
5ufGBPYliYGrlJZnkY22c8aewTZg0r4taqq4VDpzogOYTdad149wCb5f4XXisYbfAT9EERccnM3k
4XIncJA3C7N8Q3i1rxos5YfrwPCWwiB5xBcaDGYP/gRe0Ti2mj4i1ff0HoOI2CigFdKM/wZ5LH2Y
fYFnI388MFY2TF1VtgsR0I8it9F2K5b5w/jAxyiT2un/t8Ebuq26zmZqS2s2oALlgUyhuMqxpTji
XFcYl7lMU394bNwY31M55kO7CIINGbBRtQOXfShB7TrmZBYx/Pib9rxLRbjC2LZAtTu3KKgr1Er2
4MzR7nDpCYnl+jvTVE75k71jRVrNxVr1XmculCCHtedjSLd/6KqGlRhW3fBmewWGZ+y+1SScxsvK
eOYTTgBXnecme0HFkehnzcgP+MCUTMcOudDqiA5oPE0B7BKOTOOKezk3OPZzVaPZutPWl4g9ha8i
l+AXnxczHtWdASKouY1/UjLCwQd6v+KdjjKKE/BM6WcEnuEye1DSnJfFmHLEg7Y2g4zbqfNGsDWQ
hbFkLesLAe3LADKJ2ZQjOrbTrq+qFzt55+p49FL5mCROVnCFeScbSza574qY/E96vKQDT+050TKd
9bS/6iDQ0OiNpCAUQRspmKYx0oBqF+6rb9afh5gvvGSITrv0OgG+bo08g/lkb5MwR+OaisvUxohC
Y22k3ZpD0Il7FP1twPzhpjEALyxvfZ2rfBs9n9WRAcLyBZdu3psF6iMOK4hwszUyhiMcGI/1mLaX
+3sa63maMfQoOpkxWOaPzRAuPZchCmb9k1JM2rHEVeE1qyyl9KUD90bJb8xAn6Uyg0gpSSNefe8x
YDdq+aTz/EsiPFnuMsnWn4EbbA8FoWARTSu/Y3VDMOwxNz+hoKDd+mqomVqf5R/NcEvJdygaQP3M
jwZUf8/VI+u8toYfBa+EYEZBfw1bVyPOm0SlDBndBRYQDBE7QgBbhYJ2xyd0jD0WTsJKVrP0DdxP
SETAbXvu5o4WWdX5dK28lRWO84gGgTPe4QBEifUfIr66uimG5JMNox+c7am2omprWU+I7sz0jbuL
q2tUN0cDRAhW6fqUh1qaBWPCC+fuCQGxiaKmpFkCH79U6v4+bEb9GHotVrVYwbP/+PCJDyNGkwPK
IgWV220RU5SCc9Yt08VjwctuuHOj1PbzSYNVvMmjEAl4QdzeRDS0BKKk2ANhQmfvR1E0OgztSUau
fjN0b/82ZpvBN91rSgqDXWuBt+xrlO/1w/uhP9MCjMNd2+yMJnDYqYHXbQDjKqW+YRR5z3DrEvRg
yRf+E1bFWCzVLpFMrgil+Q8f4X3nob8FzpdgIoqnhlVO/Fl/TC2/Kl0Df2GdyqjduD5V5aoyoxgs
qWHklKvD95LGnS2WK2D/UwRPFwek8A4hfBOVisjSBzxWW3H5BvMUtHR5npdHntucWiY5TNBXED3C
FBXa5cNF348eyCCAUsKXNkZZnTBtXmHBQRfUmy0p/tnyKgxz97nsO2jjbCXeJM/TIL0JErOHnX5A
2G/UH3Sc4PaSpBX3mm3uhdZmeH/T/dhWcpZRsFNwwABdX2t48XOprwT08npgi/yFfta54xNnmqDL
4Z/rFPMO+KqJuEieNzHU5IbWrbI7+7NOiqCCNrnc27TFzYbpYKt/xCHIUnukubiCiJLuF/BmAMhV
7pUtDngvPI+R6AKqy1qmqNqDwo+D+Db6ZaDRHY07/NpLONO2lsRYeWQTh0bgPTVtBWIK968Ll8eY
xwBMsbpbvVaeon2bOzQSCaeA40cciGQq5g9++xtPd8q7yop+yEZNyFBoBCVbYjL4g8khiBPdS0Mv
5NLwO86+k32VazRTG7FAAxtewazGivnOK3jjG4S+krsJtXJQy3nDVVAy5WFkGNYukyC9M6o51R5u
II/ShgNFRIFcA+EaSP1gl3ZsbK9ULv496mgkcTjwkb/k4JRosf3kTvhZtQG9o80FewdyvmNJfXJV
6bJqVEPQouvUI+qG1dHqbNZS3ibZTtoOnb/mnlbJDqJqlKNckrxjIkaGiqZOcLPjP2HHExpPg6SI
WUTuVQwbVGaAvJUI803sVlSleWCG9LXfDvIgfU94no4A39EuERPhqWNAjIWCfiwxE/wXfs+ELww4
+qRChZkswU8P1QO0NGaaUaB9m1cHSoEZ+u3+nDPsIBEyBbth2me2wqfykO65ZJTRLmYtVivSbukD
zkYouC+vJ1nTSHtXvKnHv3F8T/cGuUYZm/UveSGygSvJYeH95TBaoja7AA6EGtSzPdeTdceuDrVY
a7ukrOYNTLVHAWEoVA2tQ2uD3oGv22/uwckssrJyq6jMTjB2+6rZWqGrjwh2ZI0BIG9/JnHRc57y
NtBra5q3PueK5KyJo9FLuRy9aX4FuitegPAGqbcuK5YIuLMieVU4JLP6N6exRHajo/rn191ChG3/
zTxK9ghpyZOkML8IU91ZH/f5e8wCufuxKB8wZW+YDxAjVGymXamsJofowAB7iZ0En7jt7EVVQGIi
gc9ZMPfMuY9hJ/DHzYFOdaS3c9cb9B9Sa5wP8EgmckOAm7W+tmPCz0wekGxHULTkjrIhfS/A3P1y
KD7dzEhbxrSajxOROiKcHOUE8Q/NZCaxQ1gVTkF2mxl0O/N1AfrCXKD7NAt1GXH/4pB5dAuojn+f
vf3QfnIIbjb28hSbZvYH/4yyBwUKpP3GqByQa0vAURxhZ9IAeQTDHOJIxxtwWZyecrtwvkhLjbWo
f7IY77gkzpGjyg5EusPNqokRfC7Eftwd48cng9U+OJ9Olx7vRfywJ2kQjirri46NsUvUlIuRQCfJ
bSY9jydKlTCv0sTppAEXBOg4FHEHm4ZnVVf6oIwKkMUOVKhgapMLihtB66VjqHH4Wca4V9/xoGGX
cl3SGu+m2YiHxSdDz/goP7MOfte3TeBaOYaU3UZTlWrl46RiDkeZpZ0tfk3TtvIEie/YSUzQFtKH
Tt6DSaGaW71GofFCDt/cv0p2HV4gCDuTwYyN9PcYq2x2DK9rfgFfqX2Eb9NeMxDtsmf2FhXQ0PVd
tQduv1CK4/oDYYjMLSA6upzTY4OwObkQeOxfkPE+5i7AhFh54OrF4B9TbURUTyPQLDuLFRODUksU
FLBWtCJJEDUVd6fQnODWRE9vbGAPcAhK2EUEx+YmFwD8VcYf4z5qyCsSk5TCe86OsgIxKv4FmKBg
PAx+7nlJiFR34A7XokHx0W6CPM3qlO25mDBj0bQJREKOZIhhImXiLPlHYK6xmA3EDOt59Xj7gAbT
DDkCEaBivC/oa/AL/gejsbnNUsk7kKK0ewTUYQviTPnYYuYaaBcWC75TMlx2wQko02PUSpD6pb2W
3efQ1Wahi9ecSKwVpwt3qcmx8AwHeIPUi9/DzL2HPHc0kFN/OQiwXz14Ofcr2p73eDtfdVGPF8pT
5WfSAVxnU2hwfeioMu2K3nfs5FIA9i7EHAHzcQrWByp8g2DRepcR4ghWZu3kKTDGEJ5G/RDvF8Uc
KJUCxFFeZGWyuyFJioiBDHisZ0r5AFQfGyBB+glv0kcaYnxqIaUPdvyTuLNuA00vc7Xfi4eTTay+
2Qjj8TqWk7zReAPm8m+KECKbNaPShjkR8/KD9PJHiAKjKu6PuVk9dtKTnsCtQhIbbbEPWvVU0vpk
zL4M7fBgEQuklMi72CMQ1TcBicST9JpQdpSsWKBxI8M2DfzyknldcRxNlMbiwPAKAkT52bbegRtY
XmV+A7Nzy7Q4GK5AEVWlwqhymCniUmM71L9LjOar1Fzt3EKitG9lLKjoXtuJbe9cJFLrMal9zhc5
hUVyaClJuaxXGaHn7FNKpFxaxF3Qv05VBzzleS4KZsuVFcI1HlVXdMCmOKdNbXBH1cTBtFTaYWXY
/JJpwSjYF0tx+7fWvZiHovlZDCM+4khuqcWvTrDEauGbAVP7VObZt73KkY6b3+8wjpmf6FsazY5o
xlOWhyX8XWNUZUJhBS0cHGt1h2OIVH3X2nnf8tUOva+wX9QCNjQn31UnQbpTDptpciLE5d6RTQdA
wWnsxS8OlYBZ4rtQil0J+c6SqrxcHWCCETnnYrqbtF2V/H2jshZ0K2QjVUbfQrbTa/crl3MQ0G47
0QxClRkC86TGW5yV1jcff4Yt6cYJZ4nDKeVj11xsHqeqx9qYeiuuNLawf+1aVl9qKH0/VEajeyCq
WX59+TpKo4PGHzU18tTYLYV+iR8Jpk9E2wPpZRse0LopMKQQA88q1ytVr7cwHMGfPcqLUatuR3d2
A2yG2YzOdNPLzAFJEdPJO90U/0vJ6xnRFiyUDVo6IlykeWaVHViN17I4KugU+D4XsGCiZxELGhNG
mTUvzOjzAqLMhTdNoj8pNNMQbSAt4PTOidxSpx7Am+kAHVoS8DYa59VNlCTo5j8RNI8tTqt85nwD
obDuEBBwi+zfsmfhs3YzaaNN0Qbv/fHIubAkeyocpndQ1hj6A7AwexOdmQ8OfPLXYuS2wsH31e+f
Fu2r3gFJJyIWPD+m92orpDLANiuf/HQ+h7bKJtDQbwNc/nHly9iA04qVRJhrGibPgarY8y3LemB+
rQcW9eyBmPv/Y42zD1QQ8QyXVJrBGlXJOpkI3O3+uA8gK8ACa48z4nuAJvn3kmPtvK7hlTDXveoG
qivCH45xUQOhNizlkC72clyp+BY/k8uGwSfwnrnPIQkDPT9kmHZeDAzGUBIRSn5Wh+h08/02wkfl
lsYCsNJPYWu3YUz61REbpN2N+nYjz4aPRAOELs4QywkXzHkBrlLolJfKcpJ9/bt+w3ZG2RSdjzXR
VhGO97ZO/DAkBypocnThvn6zIUe2ph2yMMuGa+JrnyJ2zBGajH6MmVXVxc5v8hL9dtW8Z5vk+YG7
giZT06BTErAefQDywFqHwNbYL8qH5uF6GD6sKkPEeiPR6awDlasK4eStY5m/1NKWJZuPgSaqDefl
0u6klKWOgqi7AP5MeF0VIKUcsPqTOE8QskcRt3Asmihu7tk+aEaseABFA8lZIC1Q+6jO9Dt4HWE/
PsdBtz0zgdJ6QFK7XTY8Guxf9pvUdOS/G84TGGAPUv712nFT17JWi3H4hdqVKfMhXNqKULpRekJf
ohRTCapOJfPd2cQa5nfwFZXI8Y6WsYs3bhPPZDlB++lcDU6gLXyoKcGXMOklS99A1iSTBvwLTyB7
5bm2BynWg0rpN3kFDd4QmwbVTqM1bgcg3UJ6PGjPoY2yzQGRGJwsVWfJyl+HdgowKrIutwMaUVJa
Iu8QsRtqu0NHcjSbmD2BhbZq7ayqhkSX3MJRA4PassGdwS6jzQR0tIITbYKc01PWYq0D64rEmqSo
j8UbXY+17fEbgvE/saY+2zhHqiGlGv9VVinpBeNtPxByyh3Jopf1OianVvipDi5xYmvjffOhqu6m
t2kYQkCGqPHztK99XbhRgvHnAMJUHJlH65LXmuELMet9zH0sxDy1OvgO0LCCLH1R5dXKRPOBrnwl
TxV9yO8pYhSesA5ldJ2kT+3oxyCB3mLYUwpebil+M+exCEatmul/+lB5IKQV8pi76ABBaXOuu/fd
kcytHP3JGBluolJ82rrTRSm+OZZ7oGCceIyyyNcby+PY7hrJXmhRZdudkyaj2HrOct4o8JqEGXEe
6qydKYNrqVos4eQTWQL2ZEsdWCbHXhH3/TSBvvZ/gfIXgoxONp+gBz8LtqE0k7s8xonMWRXFV1TG
6BqUQ96wIKTqyVicXzEgHB2L4hUhAB3RnL1rGbrHCmFlo6u1qbRF6BOx0Vm+O7IDJxCL1DYG8lE+
/lmmSHoj+lTcq6fuA/GS/Ykq8fMaWStbo6HybKec8ZpIyZrNzhcFo5Yf46DSsiScQ+VXU57oyr26
drN72VTdTX3k5jom+VPleGxzW8zKUacF9niJy3FFs5CRpPQCO7tnZH9EBKuoiCvz126kFtgPJlED
atAYoOcmSiy8dH7iQFYJR/TqnTALMKAiReGnUgy2E34MZ8zVTukTfYnncvytBv21Qb0V1QLCPyMe
57q7TZlNGmLW4pKqo8+EQl05KM6BC273qGrVzQdnQlAurOzrDN8dJMXmkWWYGO+1+2hzeAT0sa8u
Kb4Twhbq2D960/B5FKARjszPMUZ5V9V5TZd9cWJqcekkra+lZGWJUBlslJQddk3P3msAqCqWsq2y
rKSqBsX/z8F9kciYE4odQaDl1sJ59rdxeG+4BzfcUONp1iJrdUe/nrtwTV13pXhXX/QSJEMbq1/T
4OSxmX3nAdTZRZQZO2jj+W2YudB1f+10vbkUMEfm2LnfFAq5fOWv85xXfujMIULLbGia1/IggPmS
a2eUx+X5+2goQqdsZtTJ6dGLwfGI0qZEGVLeIJhj1jBP8GXVYP8DyVOGjn0DHIQU8X41B/sqhOE0
6tVZV4pRIUVThobP+LrvsOYe3hoowmolISsUDF4MGSDPl36dW+iXiqo8uyMY9PdaAgd1iWIAsAv0
nvOgwEEDhXIi8zdbm85yzt3yWvi3vtxwUKB5kKKGe4SBRLZobzK+IbJBjf4WoWylKm9aDUwScBXX
APBwIE6B5CBxDejHZMfnsnqDg8BpUCPd5kx6oqqLAwEVxD3WG5hvJyz07IF5H43G+CnmuXFOItfB
CJU1VVKrtz20VVpUiHYwVcsw6wHY5I1AFGSnHcpWEmY/Vew2VSncsW6QrJGGklP0kH0QPXEw8T8a
StcDS/HwFsXs9ZxMlh1NRQlbXZOOarHw5SS3ProEhqKITLNw1cxJbkxBr+X81E4TdQ7y9V2BAaxN
q0Gj0k3eWGDVHiEcXoU0cIzmJ80TE97H8f8ewvP4RNMGQcmU2gnbKC9ajpzw0I44XZi0tDTZTaO9
HjpV+12BDBdjl/bzfUfYaioLNOFH1ELY4NBLdc0VmoTlzFGO/13s6KCZBlPjhuBFjKZHtKp2e0ZM
3Uv2v5nUujnmxM3koR8peBWf0YMTje/aJ928a6MeRAqg7eNcGf3xbh83B9ENaGSDkoVRRLR/vczD
QsXPKRPOqdGjLE2zXri8hqstxVCAu7lQE1f4ZQB4RXKDl5aeL8SsNp9+HwxZwgoxC+3/hmVC93gj
hlCztBbESRxYmWtmBauFdiLpI0RdE0joxR67Fs8xvf3D/AXQav+151anr1MRA4QHhmFDsLoxLYeo
2CDUNpjIDCZTnLXFT37/CfDdNl4KO4/unXgqtr20Lq/AwSGg/wlT8/0YlOqVBd4g22o8uU17Bnhu
vAs8OtevxiU+s9BFIHaEzCmdb/7kGpK4LptMcboLGGt3WN9J0H66po804VN2sJWGIh/Bb322x9/g
kptP23fz+vVJ+rwZHYkuPel36h6UCyEWxmhNS68XFekskkyEfQdE9b9faKrmYCbcBVile4Q5hMhY
m4Hmz5MavmtlhNEASVcs6LAqGcwJ+cFbDvvfyJKvOIVMqg6WAfE8ghPCuDk3lOpShlIsOsVToWO/
LRrvhu23lGh/hxgc1nS2pVZSymxjltzdKlJooZSmYs7RBqAGuNLtA4gyqWnqhf53mQVUxxtpwO+n
jbq7A/0Mt5eDO/nrF+PMXo/Nf8qitDoNF8JJ5kUTipsGXuDqRaXvZkxYjHhT5Y7BADq12F3+Ytxt
a+AwPoZR38uuODyTsRqaIGi+SIXvkTmsXlb6D0G//dM5CNRCB3HUbXRMOyy1q0m6zT0FHZSKgL56
m6TPleWyMHVGGSWHFRcPkFk8/h43nV8JHldGMP+UY+9fLiP0/TEQ0EIJ1h3AfCe2JJxa5WZx2YK8
yT5ARreQDVL2+FjT4/ldinGDFQHXB5aZsVImOzQTNkCzdF3jiSLp2mQVkkVQpXzpHD1zYcSNQ0Sw
HBGYhhKzAYxtOaz373b0Wh7QLkMjIzQs/Q7NZovQlhNsu09Ty9jRy2mwO9/wqAT58YI5ZUMDwyW3
Zo5jiqKhrjn6YN4eyFzUzbDH+lD5Eg+3u11HXDE4gJGJ6pytuOV3ik5gp7iX262JNsnT2u7XbRoo
7nVY2wi822k39MKfDOTFFTGUR8yFiorMvH5RNLRmoKubrZD75dhO83lWENK2IFUcn9Gbp2U/OJkz
mi1WJ6cSWmJlsUiO7kUuXCWawHw+P6MmD7iNKAtaogZbF7nyh/r72scEFCPTQAZj44f3sgvXYA47
OardjUCnVN5bpS36tKe/NH5AqJyftdmPRds/pVHfiR/q7+VHp6LNhc7XgJMartEn16nUg7pFeNjX
QPkm+fHVMi/s1iqLFexjlrknmFBbV01n98/vPmSL5V4MuvN55P9ewhipXOq84+xoRguAqguNX1vX
JmanjEd64diKX8x6PVbRreWVJaEz3KcPJI0ZFQtkQyxIDa4IG/dgaet76ZuABTKD0LwexvOVLKc8
rR3XYIqA1ckFUYnEsD/nW0I5MUlfLK9+gFb0yUh2vF4FIF5MJS6G3Dsll7wEetPvlnANIhU7PQh8
xoELFbOTezk4tp93cl8rfS8Oueg4FWVVrdRVL7XOBTGzVwcxC8GaNrrYY4BPLD30vVGntYkm5SBj
UjjZOWgKAgNxx5jqR4eXdz4F5ijR7pPS7CNmV1pTdqXt8MX+E7n7oXEo86/rF8cSptMPVMfr8Q7f
n2vytHQHVmILZ+8s2vXPdEmnwR4Ww2N4E8J28FD7bXQuwbYNz+P+AIvM2/yqG5QrLI474fNQ6toe
CYhUBHrVdpcB8QpFf6Zjb8ZlmOu5XMHTSBe9AYrpRjUu9FSwmQf+p+UKYiLMrx2z9rq19Wb70pZY
vrILcwLsBq95/5WVdZn8s6qzHD0myyJ25z0FGv7aVMVnpEZ8dssLGwECKh71d7WlAOw7CzY33PZ3
M25XZm2w3ZPmCeQOBTmMo1DqkKj/UHQn+QEYkHU/ye6b257RqcghHnLPQ+8O2dAu/IfW0XClDS9l
DvySBX3o7cS3NmZF6ovqcxa7Cg/IcEXkYsCPCnlaOYKkuB5bY+P0TaVgrQJiIZCss8bhx0ZiSkSw
7K7AL4lttKyn7rtQTIX4n6IgVYAZ50ndkbfUJim2LYfLMr1YqawB9euv1hL++S4rI60W6UYwCVnW
5b6Cz5WWtBIJkvp1eGQl60zmeclphQzUhuMmebVIxt+1sioGbtO41uZMex+nJjq03HZWIAMWqyDv
+5dBlFBtdmQkgbZiNj/QkiDrvO+7uoUqPRvsZtYCOp0Vdlp/2MOV4mS0FQQ9c1C976gIYV6Npwo9
eGBOgATKEDG0g4Z+JHA8jOHRSUio51/JWTKYBe94aG8OB5CQ8NDronwug0DhE/HC/IOk6x3WFQ4L
BQUX9xt+/9tEgQDsj9NjxpuJhN9V5fPyFcKCRjZlqHg53xUJh9WH/Zv4w8lFurFHSEt8IIHVZ4Vw
P51ARxUBaY0anNGC5I0PNwGwCs4YolLlBADNGQayDBbQ+UwpGQTj+EViR9/S7T/VqSheJAJHz+7n
oXtkLWM7rBzQMqFI8+nD8HDQd0wzKvUBKhMCvob4Txo2dAYTKfxZxTAEbglBXSD9WeXqBryOylqI
W/QHHHNkE99ajvTdohy+4sUFsRyZy87tKFXEIa4sbl4LDUQLbh3KdrfxsXAbzppT1WhyC1eb
`protect end_protected

