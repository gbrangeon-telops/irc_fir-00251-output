

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Gub1VXq/9my70IMNYnI+loF5VZ7ee86ZBpAGzL5j+jwLQfPXAWQ9vuaGimuQWfCvI177d9QCmrcK
lRbHtdPXqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XCHJyRkscuJOpjxAlpPvd15b2tV4+cleGX5HVVJ/2Y6XWbVNSZsCQSUsTkLA7IyKge516I1wj3zW
vSbDpitOXWUELSO5CG6d5r8ZVemvSn2BJybpLquf/4fVeS1c+edRHNf6tkj5Q4P0LsQat4mBIGGY
5hCeyo5aPtqLWGIyMEw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RqwoFbaHoCNWZ4v1HvZQji+hXgCjT1Fmm8RnwPGBKk3/N74/TfbSFLeQsQ92UsPWvT9gifFKCg1j
7eGei0ot9ncWAfgeoFsw2zoynofNtXpuT/2o69ZZvCyc9OMmSHilEDslciAlUOrRZtsCwGDHNVP2
rJ/b+v8vvCejKLtIXh5C95/DXV+eEcsjEVRpSeKGeZ1MtzbV+fZPJnRzoH2U025UhnP55OgE68T/
nVfgRgkiVFm7ZUA/Q4uTOx27LPbQmDFQ6plepnrYm3dIFbr3WOiv7AWG29Y9MZiC/1j4MvPp1qqq
xE8dCNkJmOz9uD4DUQoSIb5VP26bf6BmGLvFDw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uV7zzv9Zx+u216Ml06an9UEqL4ajf0AMjc1K2s6n9qbyEnUVTSm6yFZ0M/IFYGglaG6jdDDlz4rd
W4zdLmcu66F6EUQtwXBmHtk4+/Am3fKB3kIu6GlcyUoJhx3DF0omCc81HS8JxypUZEAxz3C538KP
dZmq/6pOZleIRCziFs8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c2sM3Lkice55qsGCUzeim6Qm2yWa4rXMhx0Gil9+l1mRl06adQHebvNeaVnD5l4UfTgDiNRnixMg
t4I3MixM5k+/dqMphg9yh9uQH4HJHJ6CTIPJ7b0uq0QUv2e+GjaxWZa47ZVWMUHJwpscHTsz0hs5
a4sgfCiRr4cQxV9i8u9cWFqcZ4eu+RYLEbH+mYK06INaK4Fg1vBkwveCaGhKFtvHtOBXP2o42BPE
2i+HCKN5sLyGLlDI9h2MogiDBJsNAtjJ9geF4nPG0e4nijR/pyFXErJCeKppN9041em95AkpK0CN
GYWuH0jkznlTfi9EHnlKl7cj5ibz763zI0uZLA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10784)
`protect data_block
6PWKJqdUqnEZ0R4/bDDBJbIX8ZNOL6WPxvdZb5TYwo82V9n2+mbIr/AYdvrzSh3ERSboSfVjlXZL
gxBbBWbHAcLHMutd1Lnq8qEkxT51XAB/H5tkxPfOGIN6Tw171/IJqq5GxDDNBCYVT7Zb10AmXpiE
xEudymJTCqG4hCiBXjLwS9HIof3D6YKcAcgRw6kjVN9VV/Q1E6flNQnhj8BqkNnUDeUkEo3P/gcf
BG8C8cb1J38bOMBrX1qHWQq2FZrD5XWt+EblQssQ6UiCFAbbOhNwcvqF1THEPze2TFCKLPlwozWx
RVjSqpo8Hn/HRjWxNzd5h+SwJTahoJbP3kXDWYPEL12WPgvdo4N95q9p6aG/LGVg5SoHCD+U3/3r
BT2S84rK6OO77kJCTuSSmUpCctDLD6r6TGZHbLhWuzh27PMJZPsJMIbJHO0jN17FlCnExglbV7Qj
jnXwIb65ZU6k31DoAGMtQCVRfRtC9Pbxjg8UcBoh3ikfwSR4oH7QZ9EFoZpdyS9ccSUtKyDYVbHE
eTP4uXscmqe5eEOobObfmUDrtALKmdTrLmzi4dSi+L/rQx5/K7kFWgZ9jgnOJKCyOqKYrLZva8ee
ey/luOwfrqAhu3/oVulyv5G2Vp/FLfKDXZfc72JjqdkA6smt23dSnZS8ITZAO86tDqSEgOWcHly6
MI4uFd31ie2D4B1hg3FgbTMtnJoobv1M9uvkozSPZI1r7cikN87lCqhlgX5ilTT9wTVFIHkA62PP
PmvSRcUwxs7yW/WRDSz8SHSmkYD8hH+eE/6xS7SJVl8AL+kaM0w4J/yTY5cuTN+26WiVoTsDU29S
zJJU0VHC/VPLF592EFln3JAeGu54g7+GisUZmpsJgkHkRzaKbiYAhfaKCiC0FAbo/wPYt4DetIQJ
OVq3YNiRpnnUgaTn5hIw5o1pBbAjIQgZxAcuyRF09O8WERBbRVePAOQnJS3pOX3SVLhbARTG0m4G
dpalK5CC/6zM2J7R/eaO3hrkdgMuH74hgucfndZOt4iCtqZywp1P+givMrmeVhkwHwiPmVOKTztn
zFp9UDKpEFknTnfmFsRNlo0wncsDFEQd7D9y+2bIky+d6luSw0tZxX6+8ebGlS68i84Gam6jD4Y3
+rJLkyA/RP2pJoVU7OKTz5y3S/QnD0u2zVS7eewfyVxEAnLtGSaznJj6PoDKNrEs/YyEvGqniLCk
H6F23qoBQ0Adf1A7mppuVDJoZoi97EGAs3GzoBW9dd34NFDudiEyQJ6oCHH7b7x0vRiFcn8WsyYL
QVoGh/ndZD3gIqIzta3GwNsS3FZtwkyO+u+6jfW5cnVJs3/6zinR9B7oN87TkcXVe8CR+sTmNDGb
mAqByqa5v3VN+h4W8qpX7US2S2kerSPRvzmoDkGS11LvENam8jlqgvwW0qlfcF/uBwRz1lzi6GVz
3eVr2+XlLWaWVT0IH4uAQPoZLf4UCXiCE8oVS6YAG0d5HOCzDMlaHhXXfdduFp58No7N+/2aNcHG
aIExR0A7Ba60H/u4prTarVvrTOkOtJynA5FNnJ/h7qLUljNdC0TMd/zCoebiJYNh80M19zCwsuM8
7MLh0dKD1wxJ683QAJCgRTSE+HkIGkkXxHnWDj52udIrGIkNxv6/aWO38dxMzy71GdMAQnGVfp/3
b7N5c4zh5W+HvimEeKc4PgAG6Cw7b+aotCif43XsszJYxBiaIMGlc3iy8vN5hjFQGlVgk9zFTveR
m8Rv++9akX70wfDnZ7UgaFqF8vhH6E/0czJhHto8P3kUsspN/Ow3ZTJPH6o7BlVn1J41ZFDY6lie
azYcg5NaPG+RCKv/gAsZZLNGKb2zzYB4p1KpHsLbfaw54T5vHleGkyR1xWgedC6zrvUaO5U1crTp
zSZ/GrmCIYoG+2Ra3zZLkjbkoMH7cDuA+9RvO9IKFsPPr8gWYBcIqOw3fGihjUyTm3inQBPAMPSB
+jqs5ksUcIASWHkB4nTp0hhPqLYD6FHjwDW06yHj8bcNKHrZH8AquJlrbRpKa7UXoD8i7Fghx6Ja
ca17ObUxOFwNDuBS/s6XOP4VRQbGcCMCrx50siR/MUTxLyEpWGh/61OU61eAiTISKju2uPYJPGzU
0iSAka6V+mEmlQPG+jA80noCF21F/FZDLhpwpDfZqsefcciTgMJuoopaODU/g3q5JKVIe1AmNgoF
RReyaY4uwEIXgbNtyRZpu0hTsi98RubIhAkq+s/H9saihNVmt9wHHLDeZ+S7A4c6IHV81ZBRy2w2
4QjBb5Wdqp2By0WmAC75lJO6f8WrL3XboQFoyZO96w+Usxi/FNlnPPw1//3YMQJp+HKUiH+/eulo
Ag5KhHz4HpxfyA3Gl/WWqMHgaSeylB9GGCoB9h516PEJAIdHspSsuyoz0fpT0dNchkqrbsmorlBJ
OlPWYDV8No5sBt8iWxaULbmcN0gBzrh5L+cM64uX5+uHKd1LCjIlKweovjC9PIfLaCNZVorbG1Oe
d8Q7fUhWiGnLZ9Aej5WJK0X/5NgnKC52UDyqui5HdjAodq1CDcAPCGN+Nsld4fOaYqSIXs2oYOqT
n98nsDzWW2SxOQGoPR+lNbashppiVNEdjqpgQvzYtjV9jgwZisd3yMBuLuiy4bIDNJHjhjPxeyUX
KqPlTdS09kXseSH+I0PGQ4eRgtEdSBaSmn3UjcVMU27i908OOmXMB0zNMhRb3UOGy1p6zP5k50nw
TC5vm5xbtD3T+x+dCI7mW3Ik0OIOAAVYFX7KgQABazSnsz8Mel2HUHnaEx1aswmKOPE6T6UEVP9G
5Y5KAXherUkvvmEJ6AhxgWrasUtct21KBQMT3a2Q4CxZwHOud4HGqNq8kBz/TAZySyNKeEuinsYu
PbWDfgG48nnwlGM+I+jQb9m/JD1KHuleYoMfAMDH+ZQZX0bGORSp2mbQ7l4Cd+V7m0ecoFiZRtgm
T/fFmT08i54M4hOlHfAWGcBKrRTVCF2PZe6CF25uOFFYXScQYvw2MoDb7xjzYBMx6Ku5STFycqIK
IhTLuQ01NKq03iwVTfplieGb10ADo1C8MXKnqOnj4vs2jjdYGxYomZ31IcBY0Bg4D/sFJ5lCPqTA
TW5IOVziI71vaXnL/wNbnhUCdMFGaZxE64usWsCWSdkIFI8mw5Jee51nTi5zwWtmrv1LCCx/76Ne
LlUb813In1TQdCerx3Enu68LaKS3v75xb0xl6LTZSF9Nv3rzq10OVTXWa1BRyFUlPCmqdsWWso6G
XgO/XGsKBgrKDtDYfJzxQ1kRGxp8DhkdCOF3N6Aq2yL9n028+18k1F+sucUec+uE12msTiOcF6BG
QH4pqlifb5GZYAMbQAVWFQofUgmHoYGb71NfdaMNKwCza2Mfzf1TNgrMTuSM6kMW4ZS5VkRD27YN
CsxoTEUfQm6clCrXrSYb+YgNiTbXcUEXfVr91zwVBVRVTguEnmiKqgU6UfZBwJEGKBYEZNesMBMc
FPvXiPgz1+VR+JPIORpTyXuro9iO7ewJgY3kSwIqZ6fkfKCwipGoq/vPHcN36rQFLHij0/wTtk4s
2wQElK1QflqUJgJM8IPKACZN3QcKbH8TW3M2S0ztBbEzUXM+y9hn7P+mpGkUfdBPpCzuLkWZnwZ1
9+9sIdxVguKpsNABTPGe6zUViVLYt/mvOxI3RdodkUxok+tmhmKysx6UI3c3LWHRLGxi3HBQx6LT
+axdP9UQr81w96KN24+v06BfHuQfylkwkHq+sZktd2hR3Bj4eyqwmEMC0/Q7JklPZCZk0CdZ92/L
aHqkeHh/Ll07p+p8jNTznskN3VcO5qYGyK9lg5s6EUu86hMUjTVr9zUm0WNJ3jL2R1Ng+244ZJLf
A1jobZOeW2/T42+lDOigDIriu9pP62fMSbZsXOpTxfmTKloZkDBH8yPX9Hstx68iAKrEo3/eDyGq
S/R69fP/0Pbj8xIuWTNF3U3V29idIfIYZ9MCLWEsa6Lg+4ClEYBlgrO1XVfHVgpK75FAgIRQYYAl
cYRG8YfKjxuSJFIIM3+ZuslF8PxkyiD+VprOE7o+dRxj3vBA/nh1a69narzT4F7hERT+3pZG03/L
nBkE3EC15eA/aba/p6g/ZvQj05nJly7PGPTtr8Lo5qqaOZ8Ioylo/+osVbZqm78Wa2MEwHD531VK
sdMUuOxu2WxUsqnzeg//mzltEgwZCCB1E7DfAT8NZpXmJJL9Wdj1jl6xznJUNwqWwTrWu5fGAmSG
q8djLCvlYNzZvGtYzz7GPxIh0k4OInA7Gn+yOq9+wRD667FAtX0Zd4cTkQoJB5GYzN9Sc+hg3rwt
3ysQF5dU25/kSVFkhB4xuLfKBh7wH4RiWy+us/wIl5W3MZcEne8AJH+0ZgXn9gU4KwKwgWuI6NVf
Oo7BB2zXYC0TJIzIWz1wvH3O5fCQNXmejI8OjF4PFYISD4iOCZcmEJgczCqW+py9RC2g34XUAWry
nORrOLi123mmytMDLc93h7UtGQaj1R3wF0O00WaKRwcYUPewWyqocMGZZPcbJDZqx1cEoNOcJmUa
nYal5I0Ap18Aw05nW/dHSZxGnsWf62aPkibOVlaz7v/WfL8Pj4ETylxZYetZn2Q24sDkDNDbfGK8
FE0uCgKubpqZjT666JTdMg3TKWEXpK0CdQS1UmJSWe9B/FLXjnJPA7hd8E1xmKyq1yR9oY3faSm1
QJzssTbeUNIxPKNysBx4KYC14vNICyFsRK3uoV96vV+KAg4IYFAGi6tmBjWO+AQJjKdsYCauET6Y
T35Z4MyU7BCi4S5gQgtpOv8tMMfMkaFm9N90DfesVUXSNYDuFVi4DHd3zv0PuxNbuXBQ0GLFeHPM
rcP2j27LiBMr+SZscYejAS141l4efvplrez6VRObhTVf0vA/N8BjC0uy3fM5yGFvA3FBW+wa5ccl
lxFsrCYKi1+uMq95hjaxfemC8wKBCAjaBPI1cWCVFwBrYqc0uSoEwJRSzzVwA3/CbVcAWYUG08ag
gTab7ngZuTmEyVc2pdC3HOx4VorDxzBVOTU4HMWNYq4gaOAi720A2wQrL1C/dTrEOZzncHxedKnR
l4HDhL2P/7+7d/45AaAgY9KOoLuQIYS3+raI8LUyLKN42YUQe8SsXztPDZiKAPt97hpA2R/vdLXY
ZWwVkvGA3NbR2iyTMeYry+Wo+UmlWVMJlCY0TNO58LHqzAk9h3nQ/S/ndFEOxfHDzb2KwbfJYSZK
FB+amu4Zsq8K8bULtfpvMex5WznpJwEzuYTfUSc9V20D4mzoIn3jEaYZsAj25H0NrlWUQThWBUq3
xSUtTIIh0Rd1j/9m6am9DqbZ5djMXHp8vo9fOjjVizNKMey8sai18urICZe6cXZYmtjh+ekqnzUd
3vJCajNvMjxHKrV1RJk3L90K1MBuCAI7H69ekulEmjA4owh60IJxKU/RqUqJR/wmlHN3Dbrjf7l/
MICJunDMy+t/WlsqL8nTpfrZD4habLPZ6c/iDRuDrbswbqG+TcJEXVVrmu2ov93zNMKQJxhuDune
P2MELjZy6QMUV+axv7lAvcRZYicGB6ab3iD/kYy0iV+6PSFs70lswtAvUciXrHf6LGj+Qpy2+QTK
2T0i6Wr+WxjGslct5P1jFgZJej/FXfnOHhj89R59UnbBdywfG314xU+B/T8fNkCd1u8EiwGcL09Z
479UugaWYQj/MDP0MuhMmcjbSVvCmeQgwQbF5wLanHfBU4MaTBastQRYPlWYmr/qcQJ0szES/Cjo
JMBPPk/nh4kT4TJcR04v0RZcRUoH0hy1efLt/TG/pugd9yRniR43TRhx/k8dDnlunokchlNyevXf
mdzDxM4a0awteSFsN9sKyiuFOfemAcU6kJHBOq/jumX8LlGQmLkgSgzg9SLswsECibaq2DM8LWtv
RAcfE0IaerJlFtGsUv+S0+G9hbLcpHMqOH5QhBgEd/gClMySttE7J2BdvtAKXKuyqD5h0foOHDZi
cBx9En38U+xUbs7S4X/g3jkBnIP+g5wmpLGPndT4hbOUX0eQ0G6TV/RYjODmucauZibbe7ig06fG
zsmxqZDHWIrUv2t3MwSNjTt2GnMTFFhVQp8Y8uAEZJBg6TQt/CkN1pvKVkLLVyucQC25se/PNa7r
9eVQEsRXpqMWFwk5y1kQJjReIIMAy9QJLX9sDyBuv/z4wYuJMW/P5QqH4zJmrSmGthupRYajie1L
CtCC0x2OxdWBq34UmXPT3WY2+mTzo5Rem9Au1ubACmXZUfMYW7VXnRtESrQKdLE5Ycs8Db1j5oB0
3XVfb+nPWahbI1GBrfkMN40gAuThY8vWmLFNjfJx10pB9tBZmOyDfb7jnrVHmDy95pEtg4zSGcu6
5/Ox4fyLK+KzcaAYuhffdQoEk4LpKQiy2ofVDYPhzMMPE39id665MwWMxk2du3+LOik3ZDCihOHy
H+3ewQud/3Put+vFza5hTDYwJS5ZZHu7CLv5Tzqd4B6hAeelidzUZtc62UJqCGdAkCsw2aD+wg++
hzllEopcQxhJgCsxOU8UangRTX2g4UXq3EYOXIzu1bJdIj2ANCaI40789TQ4JANQlgLyja7z7SBE
Mx2e/yCe0q47RZ0ES+8bNzB03GJ7dI7UiTvxcnWEU2tiaGjb5Gd4V5gY4nZeZjbpDapxdHzWmVJW
JNhYmRN9WZ/EC7i5PJXxQ2ausUz4ZDFb7jpM9zf1lRtpwuqkI3Tu51RjLZ601Yb1yeXUqqE4Wv71
t3TiJxb9rK4To1f1OWK9WXSsVA21yd8T3khRQHP4ltZXL8q/x/6PLzHq3XmbnPdTdMVxWDLe30XM
taPyyWnGx7kMNBQ5rvvWZMV2zbSFESqPOhheuKzCfSW5ijDAkBPJCjD3bCSwNpwMlKkoCwfhqu2+
AMk2UBqzifD+AwmTaKnRQH6O7dET0f2OrP4lQQH/6px0oHxkEfn26a06NCykzzy+uX80G5xtwceM
+4IQEOylINpy/hZXp+yv5KLU//pN3+cD02S/cGnGO8kEvAWozCYiEIfXfvBIf2co4xEH8A9RFF4T
CoPrjgKWxTH6xkWag/j1zZ02ixxXx5E6qbp2RPPE5NIKmttz4qmJWR8nTakGf7RnMM1Ydc4Su96R
lhfy5O21RwLixvCVOwxCaV5vt9EGECdYKC76PTi6d4jzwJ7IZFjrzWUMjvq85dh/oaEy1Oq8lnzr
l/JQw5BObe/7NVoC62J5yI+MshEdx/omuOp+R2fkwTFgPT8Svg49cvI+Uc3Vt3UWmZHKlmaFrHF6
UOwQRHR9Sf+Zhgt7RVkec9UvVMrRlzLGu7e5ytWhtkBFjDgIWxSzZf6GH3+wC4ZeSygXepI2SCj3
SwSOXLPzMBjn8TMmkxGn8gIsos3oVSqzyAToa5Rhwcqgdoit3U3WLLCek96MJNwPon54dR/nLCPC
tSwv3DOSE+Syr8a0O7IzYE6z8XPSbehluBE74uYaPjUGjY5qcG/3DjuGax4ieL13q2XHMWPIq8+A
JiRWCWg4unyMFMN/Jqpgyc+r2BbGrzkY/3zeHoSxdODEmNnNpug+SvDhy6IwM/22upVBIXQaDwSI
7Ywht5VERXRYRQIf8irVmP7f56mKP+vWvq3r56L9t74cqdichfeQF5sz3n/oLg5odBbR4G3wsZph
WBP/t4UnwYNaJRF2UYUKeXoKtkHbM9fzHyMhRsC1A6uLfYQaEx08008JBVBQMGQuflJPfHws9Y+R
TmotKxAxxRr3oQ9DWOOeCzQDWsj9GFel57fb5sxHRl6WujhSyugcyClxX0GX5uW3MngyenTt0GTj
GRHD2uZXGzMA/39QmNj+uMeYbTiORW2X+pAA5htL0BYkYJY7/QSLT/rwGCLiGC1CThiz27rnmjc1
i+S77IfZgfST2WWzrTfW2hT/GoWNTKfMBf5xLd/8KH1UyfJWjbKWsLJwIuEzjbOIr+u8brvwhv1R
Y0Euns6+VDiQ07ohPf7ABGuwzXnIdDhc4vmXKI574HTdgkdEDc8oJrCnqz4MYogBxYKtruSjlvWU
SafEZxxmSsEF/KmNyJUGULfjsZzc9cBqNvPrXgckxY11DbCDt7+t1YgomGkqdJ5rOnL+kRQvRpL8
25jo7p7v9C1NiZA7vlNQTRZeUFlWnZZ6PFoy0VyyNTuYfeyuANiIOWV9K1IUFsdGeXnPHX/G0Dlf
EbfU4g9RYWFDKjdlRVbMyE9OSTfqWb10D5NWQ7RuY4+QFUJXqCWisAb3MIPFO3nukMwgxMUKuTtU
M+CbwRmXJw4Awo8warqgzuBh9ngxxgUThHqHpDkF4a5A8J4RHFVQiXOAFIM21h1uq+2HE9xAKiXc
hjMEDsqiekSEUkw2kXI3Of+A/KPpYi6gYO97wUmmxRf5XzbHdh0nXeI3JNFoSI/0wUUfpdNcEeDE
UdoqRBMnwogq6m+HCtSK50o908eS71VNFPDqu6JNebvtXp3xVR52uKvemuPJ6/UTrrmOg/ZbpMPb
aP/1SATQaI21TrjOD4Pp9Eo2vlRDr8n6bqgcp4mV7yQAS+ebxDnj8SSOuDI1Mt+02cOHNIjwkrYk
gnIDMtwI27OVdc1wGahqVse8a82xFPSrciDl19lH6EZ4ISiLHSShe8voZFC51lPBuAx/2XyJc66M
sLJCkVcccJ/iKprPmdUfsYrp20QLTilPsY5xSZGtWh6JTnRWlo08C+U3Rxy88Nr6C4KIJLil/+fI
bcqTvYmz/LVGh07JXSOAc6io1rOfuGjDyzM9rCP8wA5HlvUK3H4O6KKiSV1kZS6w4vUgmzZjikMi
KfVZll2WiN6mz4jvwWZUhmD+NsOtEye5DA7963l1LF2WhlGg5bjbd771aR9R+baLGmt7vMD8yY91
wcmgD12ULKbShhiTo78Hv0QD0AI29HkjNOXThJSwAXKwReAqBmvwzUWJRE00At33nux4d/XJt3Re
Hr9YKse3P3whJx6z/I1clLna7t3+D6ztOwgfwz2PXLpfLzmvkMpRa/wTlxPF+zSy4DkbEQKWFbyB
DycHVceXXNiUy0HZ90Pw0LvLc+VEkpVhOdoYtsbTPtG4wX5tb8WZp/xrJBKf8Ng/6l+D0rwjNuov
6XchKs0kJ7XgewgtYhC5221STou1/KdBbue/EkMmD3sRmnBRHXMWlMbgsQ/dCHWSpLW0Ilxqy85B
7FrbNj9seelUq+EMKaKddC1AQYQBU35LizVYoxG9CWdRuoBn5pi5f7qNF+JHLtTSdf1fJVDUngxG
Hx2TX72fllHeRZFe9dmtwdOKGMMxj02WawJgp88kqR5E7nN8/CzVyz+yFOHREcE04TWhQb8XSLvF
u6NkloZZm23RsmJL7gk34xzvkb/HIp32orvlYXWAbVhtLb4g10j92WOoNqg0fMhh9vDPBOnkaJib
PYGhqabis/Fon2mvvAvUYUdM4RYfVCIJRyiFnjE4Kxggq6ofCNP4vQ79DIq2B9SoiypMLO9Ltrrz
exQI1L6iyK9pRIsRnwZ05vGvp008CK6d/e/9/7G/kUdBHRCOTOPnwgMQoO13i1OW+qn0s2yoVKTk
vmPQ5CuNU2y7fCkcNUcA8+TxSI7m2STUOFmCyjA1OCGiVO6eZA0p0LUUNZ7xcCnfPFZ7sOihb8Sy
FZYtN+gITDa2JiN0gtKZvZ9rlzW1mjatFMLamS2HDSYgnwXN4UkeVCOehc8JAPN/rwPOfBCXkgkr
xo2ZunPffaHGBqRJKUtFcreec2GAnzfHlt7UTpk5pmVCvjupsF3yVt+86dmplFOEkhBGE19Jm6G8
jxLlFyzmUh/CelTx5nkydnupCOioy+PBsUxjnTZYja7e+GuTHYEsb5DLm2m5MUW7550Ie6HKpBlU
LfrW3INqbJnaiywYjSwta3aOnE8Vkhug1CfPdmM2y1iWTWWTgxNwwcpHt0AWl277l/WPevQ7ztFq
48K3Xt/G7lchr2C4KmuJVbPDMR5QnaiGdMwB/MJlSIEXmaWjupQAIe1Mna2k7U6Zj+Bh54sIzLSj
fwmgh5MCPCgiOg9QeuMiwRsjDuZl+B5+7KruitVUji1iahibA4DK4d+mBUEGtGJDk+YNjg/Gz59Z
Q6vEwsRZqcLEdsZWtO+lmABRK5JjwaX6iKA7KCOa4baslmcnQGfsEqzjuaEe474BYExbJoBHNAFx
iL5w7F0inpewMtUknbYi1piHre5a6B4LiL9HV1c+/gHRQ7XDd4hK8pReV3YygV9S7Lwq52rhcaRc
6o6ACyFyqxsx2ZouEIlUbj19c9KFuPQ0ijPXrGf3pfTbahKmssHfxqcH5hKL0QUH6LRF9KAi3Hmx
5MjXPE5zqRqNpwaxDTjSuUigidhZoFoI+vBDQvNMuQzPDrqlV0bLWwjyZeC7ziC/aarWXYlldvFc
UbxkHwMTPCwM18Tx/IMv6YGz1o28XxMYzYAGhjirgZpNHtuVgdiYtOwUzE7I+t8225z+C3DQ205Q
DyJDhVtRrfORtFx2HA1iH9S9S+N1JJq6kPhnPAHHdmNqeKSwN17kgCj92c8h3INQxiV+AY5bTzCW
cMnyUqYpbmjYznOScOEA9Lc+XYOzaWGWLujXqMlaz3pk8ZUKylgQRAL6J31taYU0zZ4PzXwfTQ4q
xzQxBg58bTvhHvy82+63C2TCDfZ78p3vMlv/G4M+ZASCiZ3HaMhTqMt5xaxTJE8N41Rk8JTyGoP0
6LIBBBAqKlzWPMTnTHRxBipwMRNnwGq2aiV/hlvMbehFuTbu9mnFnXMTJOp0sJDkRH/+kOpzLOTr
+f0cqB5kFrLWaHGeQ3f+yDIEao1hD/FCsjKNVfHWbdrDmYi9UFrw0+eU8oellJkweNEOcTR8Bk4B
AB2DpuvnKh774GvRdhZuZnMn2qc7uIPAzmT135C3ep8JxO96IE9RcUPNx1clgVKOe5eU+tF2pEj1
oDSW+mC0NRr9riix8uCikG8zMctWRCtX0QtIr0hP/ey793+NxDMkmSP1yCYNh83UG0tmkZLcYMdg
Ut2cgCdPz8gLlEmd3GEmAPTKMmxjP1xyB9ZwSMjp7yLL3p8oim+VxDRu9IuvLQLb/ci2qO3m9diU
8ec+kI0lYDThzNqopdjQ3WA1ZKK4n5ubMOwspghrG2bPoca7yHbfKRdr5f2ZszMudqi5cMK7Mvzf
Wi9jM8BBd4KTTa6eEGxpDl1UFC96LQ4FxgE8b5+ajcrjNwZkqNP+LhkH36B6tHRar992VIVEbZFH
C1bSAZeHjHwcfrldhrrjn6JRff06fV0daU/2Ut8tWsPeV0Rb+T4/vOyTnAoGnKfsUdlQsPkhFfOV
llnhElxOk3uqFRMnUWXzUUa87/MH7jdqsITrdR1JGlvkcmLGMp3g7h2fM3eb5RpOoR73aXn0xyTX
YsBV5JtCevOHjOA+iGYWdXOq4lMKKeBaQ5eBO+JfKFGjOikdBTxxkQouogGZ04A9L/sG47c9OeSR
UzU8t8+MjeGSHXsxNeofyGuV9okdOnUrbVtYQCciIU4/6l8jJ+SowRp8aGdff3boTr08g/h+QH92
mlORAGjdbI0QU+qcYbseAJY2WvmqT9LD/xmNl6rcUbtckH3xnfYPxntmj2mxT/7Ynw5JbYiSGf4K
56HqMhkJjc3FnGGAoXcjBjzvvn2/o37AGa2BhI0MEUSRppvbgC+VsfE95WEFBL8MzVQVmKij4/5G
CGmq2j8vvWiV0Y6JFogs/UC6mUw9tDtGtsLxqhxd+UG/wjy4TvsvN/6jXdvORQcy4bir4cFP82ig
lxEbHmZL5ZA22vxdmCgbqyh8UhlANutk01oVyI4dQ8fgstlIRZpcJTOlZ7vJJuMlyy7GiBZCHaxE
no4jCBhJo/fyZSzyvTtUpi6oXWAQOx4hf44tV0PAC4zOI09Aye+2w3BLCPLVD9FamPcmb5gijux1
RmYBvE5Rppt2B7T7eC/RKXSlAslX5FAQ+0fxnozqYm//sRlTQefzq8U+P+Oo3NmuxoF5PhUvpaST
H1EFbz1nrwKKchlnA98hiR/rwmrBRBJlFCPEq4kyEVpKv4rdEQN5in8xZ1/IJbeVn+pEjRQiS5Ph
37/kdrirVvE3ExKR3IKhJxP3G+dN4+Wel644SyDhcsYzev77Ucn6wxkrirDfe2sWHUWfi0ua5QH/
cE2cNcDkTJLb/TlNc6Ps62M7Z8n9o9rStSov/gB+w71erriVi42x1lKJpg6nfrqdXccWYbEvwjTz
EOkS1q9cjc5VE/mjspNaHGB/uprWa3EjU0s/fozOqGY7H3atNL0RKmAKvN5K1fnTXGnHd39NjSi7
So5Y9eitNMTde8s2/yi6M5UjD29YrQqGinfYfd/pbNOKZC8adG+NMgJxDRcuVo/Up07YoRC+lLvl
aiJkSCF1afeBaALbIR/jGRxMGt8jxUx6t9pMvP5/rbrnJGMGzjRMBPAdJ7hUFpQkZ9ToTccloxyO
Q64vmUNugV94RHmTZ6Bz0KExiiwH29E5B2WQXlwGWHEaqZImyRiOTWhWnYw7sUydi1iz0Vmsmp6X
56KAqO2vBmx+2XAeN3H/vjN5iDWzf41P9/aoS0AsVlVSr+Ua1N0+ibo0SOBXx2g0gKVuZHqsPzbP
HpDIE649c7GeDzOQKwpjelcs3fJ2abFb9CfTJoGnN0pMcw7mXChl1K2064kXdch1Y8zo0PKoXN5G
b2lIddW2LQz8bNm3hllWwCDrUC61I7Md8Etnu9hIvyS7HXDy1EzGXuJKtzV77VkAQkwsnDvTGw4j
tWMk17h9LOBhtzCPpef3bI0XIHhWjEZVAOulVdRQeg4QVOoHkjQ6SGbyiAPRr7pJW72b9FHfrxpb
59+PeTS1T+BONqDI+vZPFDWqzWmtEscOs8/oEN+pdh0/zgZaE/j8XKOv8IbxdjQ6eF5oUTa9LUt1
gggaKHcNkeNAPhXXWNkczmmRimfxvvvQw68ht1m6holoZJyDpIF6mV28tJWBNSzIxyiNTiiudGP2
nVRdGtLN5I2eOWx7FRKdoieoPsF2Oh97dUZn7CJHIXJmsrY0qAuRiCm2HEof41SU2ZUesTsv0Hwn
k39puu68gYAxtAAFeD+yMVgmUMhvLfEldVRZHOMGtQTB5aOuV5EsHRTRKEuuNL6Py7vDhYl1VVIG
AJ+3sX1E1XyJYhh9nqb4rPr0Rhnb7idlPMq2GOElJinC64v1YgD0kZ2gWxa4nMau6DRSmhbNYwVb
nNynGhofSmjUa2RXWNd89GMeMFVX/3CjYlIikP1KQDaCLPwwLIiBi9yeUkdMS2UQn+ENKdxmiZXl
j5kciLjErAAjgUn1rCBcyaCJhA1MACNyZsDbMEhNiKEVOfg+keYpr46g8RJuvU9guuebCC3LOQ2l
3qSmkXrbx/pOGchSolYtxjRlVWmM/O2OqgoW87oHjmzlgCESQPzoAVwKQxCwdhAA7J0U79yPWgkz
UFAFUIWccZYGNTnfBQS0vZ6o8PVk20Y343sU76XASDiW/YjiUbctvjdD4Drd+u4P0LnoMeOk4z3e
l3PJ1cqg32HcnjQe1C0YPjrZDnHjoHz3UgfnmbhRI456FtG2oSzjyNgBrbDfLOZi+HldECajMfBB
53wdzgjdb5wglkNjkWayUvc+vN4pxif0Ukrotv1UzYxJt3Z7NQSDSGGyaqZRi8PWeV4SGvpusRCP
3auZ1F7LHZVdQTGRneAV7r+u7LX/iLBT7XsSKvfdcuJZ14xWl5qgVH5oFfti3Ey16EtCO8I975iw
7PGGdgkwj2hsZ7/Mk6CcxbkRwYjj9YUUtJwHCTNV58yrUIUoPGn8EaudQfqOTiCrNTjG0b032yed
kcCl8C6qSvGdgu9LahHsf7d+YQNTl/tfTUpcx2u26y8c9DPFYgxeSplvcHf+sVA3paKkcI1LTo8x
P6LtiNi/Je7JiYNtfTNti84FVLy7RLjxSBOD9lkzk4vGYZyWMr//51LGGBCUjP/tmNJZcl+tVUTg
cpqWIW57byoRjc/diLCdoWy+euOgGMOdRj7FR2GblrREScPPFdBh+IaWJgN33eeO/Yiar1t7gDIt
cVsWtCy0eyZjFc6VCCd5vb28edN46eJeOfmjQbEfdKks+8LJLpaTS0eHIHZPPY4q/7VUQF2BhR+Y
y7c/g3mx+8b+OCQKOO9t+LQFKJnKwHitwzFPwSGDCIWOVc2BW1OEA1qY3NyQ0rmM3M1ky3ODr3iB
rj1GH4gswBskpc3WMaHmw5dU8QCGdQrrwEF+jwfQqVcgHb0R8kRckHJkx2YxsQjd2kA2/HNIFgRb
lEVKoPqLFCqErnqI7MFbHW/8P4xsMRUaNn4pqxqA/9yvwjmEQ7rh5HW1NhljwnduLRSOSeMWzrbZ
GgnWdCkhzG99pas=
`protect end_protected

