

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DoylSncttFMA3kx042gUfpgfS9f7wYF6CWxJheifm9U5oZE55E7a0/gn13EV1/Vn6tAoLpUpkm/0
hmdlNetDYA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nsjL1A4AfS+U1MlmYTovZuA+LXs5hJP3SunimigW7xSFqc+G1o1qnLbV4BnmOncmqUv9X6mR1dbm
lvuLbnkHJpdv3qype+E/DkwUU+uuHlSP7/5qiYqLK0/kXVQ9CK4RGY/33UuCkCUXhFP+4VquDr0Q
ctFJ3ADjSF9u4KfkLp8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e8PwETDI60MBXnrgCDSTetYRVktLV/+TTSXZzS5MByZtHEX2iao5JK/khM4FDpq/v0uNsNW0rhjn
1dIPd1mlQZEDfzGgZ7rgxmjzboNMUH8CMdtSuB8lFy7Tjd1hDXqhliwc0PhPBGYBs/YEff98J5pB
EaQ7x9e3Dm3lUX43BX76qZ9cgUsaVwP5tX42M7Z1CZ11+5f7kvoiSco/DGzJuhCbDcHoQ2NjrZeO
tRQwYWFDIi7vBls1ETe/q8cjQLCZThAhSFjjijV74aEYat0gpNy4Hxz/UN0rUMO/XCqC2k8lo74U
XZlHepR+ABhyrwVFzKEwcRDXuuh6ogUCrZ1mMA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YvHkp5oDmh1yxPKtyY+bCFF9nl00iIDnF4JnEfzCQKeCjt2Tok2cPb5/9L9T+H/cQ1x5qpJZSOJk
cf36KzabCPbu4/9VIe9vwmzzbE9Ndy2Ov8q4+HYXDGn/u3gDUJZcIYEnVlc3E6se6bxCrEZNyRYc
iuoolgurhXiPk/HMhX4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XZ/Rjfda7p8W+LhE3BcXwsLXrN7RfTJezMmvWQf9ZKb6JJ7gmlPk8WkUFEwjbu79kr2SMWbEP0wO
UouQmHkylGRubs4N/1VfavspwJxzO5pggGGBLKHkmxqVxAWJEQ3Kp5uoaJSKWxqKIRLzeGXsW4p5
F/e0YM5v9fK6K2B07V0FxCP6WuqrungKJmSTj1Ji3gWd+VJATYp+hkh4HPUA/aDTgCzwwIaJ6QWy
QvHMQKHrEHbRztbzfLMH3RPC4Jl5v7PMeYTnCv8UcX2dwujd4zD00VIt1jMD19vjN2WZ7U8Tl83Q
sPvYlUbNQVTnqIBf7mqYAoAlbAFXbg0t5zqPAg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
tMM3/cMZjK45oZA6kcbHN0qWcigtMLXglFSRnHAR/CFgzf0AMJDmxolHb/eU/4AZu9y4g1suqZaK
XVFTen2XKtHGhP4VWUScuTIW4ZDH/oV/HifDux5cP6Dssa1OjTsAQ5Pzr3yduN8sQY/eybeLz7Go
EKlRwfCP9BFCnhs7utCLP6AqWRzt+tDzRdUWx8D2TIvfYy/yqEEbvEaGBhJVS9ngOU2o21jPKudT
+/lxbVknMtREcrc2QNH1tdShRDYEjBwnbDxrdY7DfeFBzbD3GnyBn92ZghueZc13v3jqwiYbx2qB
O8lVm6TpnpYLq3ErHyeWF3HIHOS2wXrRCgRhfbKFJb/rCOBbh1lfZeOyvI8eBX1VvvTmhDA6TBlA
WFqidyefQfNoUJS6HDTc8tsArIuv8d1scJucYmUxfsZOn9xpFAKdcuSgQ5x0js81thgi8ICk/4A9
eIi8wSTXN2wgpt/qdrpWoNneSTNU2dGT7iPdm6oJ+58zw76oSoGP6cMHAX6cUEKx+XjBlT8PokzV
XpGcA4phQHzJQuPuUYV7mU3DLfUWkbpYHeBXHogan/NtC1KkeuIO+UATx2GRoMXwt2ufSeeVQfKd
WZxRk8p5XwZ3q513p2Y6HiS9DiRwBPiLarw4qXnjHPJZZ3RFoS/CmCcGeTAeGv66UvhwkIN+lkHF
Eal9PXTz5A5vezfYBcQ3omNLQyObglpFDo+BI6vCjQp5cPI7DffHnsHuxHxG3drXrfcijz+ztZRo
2/WVKP53UqcSFl9Q6FwHSqbl0IkD9Rr8VrIZnrckxNp0maY+1t/eVYqlYU07nRnMrx4gT44Cfmx1
+svDXRCFx/wX/p6jyJaVm8JcRqnHQXLGKm7luMkE8PJFLekcl9pd4QBliyf8kay/nzUw0DX1aKw2
qMlVRLdg8IZySC+5Ss8PKQ0hk6NwcFU9kcsaJ4aOu4C//pn8/1aum2kCmiIfPW6UgMdz802dwvxH
MvIpklMBQsQgSVuzASbkI36Koam6zEDtpgsBIfD/EOpaWC/vEYhWkYJsj44Xrdk/tFE+K1u6gBJ8
U3tD3Gv4URLogAWk1m+AHBGBDMuCz325NFzal+3C7mh/Da7GENwjGuNbZXM76V9WSbOhqceaoCn/
sYbTUMivH1kMrLAvQnJsxY56U0ogInSgoLfPiUmCP4QlvwFptqTJkPCEzo2mDHLH4L4Oaj9AiwsU
K3AMBYsLpuHYdGFR0gkdcY5DHbY/+3kTaiJsC4tIj81aOr30RFNNiYMp+KCHqlcnvtX4YZiJ+Cs2
ygkfpu4z6sQ/b2ni6ntBIn+aFIJx/kLv2e+6CubuLFk88pAHimyvBw/Pvj0Q5LlDkSGa/pInHEqh
eSXKmCv/1DwcvXAI1sLyjifAg+Jy+Kh/JNy7DaaX2IQ8L34mvUOAXy/Ycn6C7gyDAyIhYLf01tDL
hg1FmumjP9b+FVtTJORjiYciXOD4HH1cdsVU8QFbyXGnpRJwd8lskRaMzXcHNv7IkttmfQGOm3cj
mkmX1BQ0lRokePfycQCXpfpWo16SFpbKTKrofnmLNwAw2zUTITbSCBlMGTeKIEF7ssgzLCcSR/+X
ilbRYGswYx6Y4cFHMBLBDeUuqavUQqb4rGUVV+0z+oB1d8hHQYSm4+DF5sQnqv2c6zqdaCiM7f/w
IQG3fQY6F9pyn/nzloTSgdwrQkQu8p2bKwoSxRFs2JJ+EI3mnlcY8NupqJhrYGCSRrv6W+fIfZiI
Skj+13sDMQ5n5pqYEdWqXWnUTFU4ZoTXr7i+fzvseZb7++8+W35e0UEhW6CemrCHOEm7wwh0sQo9
Rl9Mfp478vKKqdJ+UeiBCg+1JUHAlHXKMf2wlii2SHHm21jy7SP+wC/WAO17CFnbO2i1PUvS0OLM
10gsEieN8CX7Vtm479Js8Ni96yRK+OAIVOEov/v0fF2atlcXi3Pi8VncYSIYjWWSaLLJLHzpIMYE
wV5VgthCF4cO7lZxNkqXBE3/INM8XQ+yim8KD4UpE1kMtm03Hv4qbEZ0h/muhI/orchc5KieyfcG
VCYxOHEc3OsYbHamke0h3+ssSvDHXH08EqMIi60I6rGxLWPjyATfJkNelWySA3JRl/0NETlPfAXO
rqlstDabV4437VZkr3+10EHga/R/HOPhfq2c4krlytRMI8xThvYagSuccLYid5ningakYXZQT6sB
aakLljhENWozGZii5PrwvnbQlMYLkchwct9q41Z9U4w2weboHHXyM1QatmzQUxoHlSW4zTS6dl+t
HUgUgQA7xjO1qZIojUF8H4Gb0Y9h75lSYYzn+OOSvVpTWlzAsfCgeIvrDAg2xTgS7GS5Q2Z4L7Zs
L1s2gpNEf49ydhC0poHlC724o7x3U03s0AOSjYhaaIbkMQRaNz59Iq+X+4vd90Krinq8WXfN1LfR
JgPUrl9v4o3b9LpWsaszntp084E5nP2d810isxBhGgz7mV8x4xvW2fu+TsLq2IHLNH8SsPQ0f8uh
sMa/4VyfhkI0c/YamjWEO2Bq4sXs2l++lz1GmFKecCkK2Hx8DR3bAB6OS1RJa7N9X5YxsjioC3GE
zGiLXbWg7KL9mWePML+C+nDST9sold9PmCMLsjCjqR+CZMHqgWq8ELy43mEzO/c2zp1kX08LqhI6
XFgVYtL/Q7sqNdrasDXLO/aQTLz24bxL7U6TnT03iCM5s6iKfxsbViCPlWONiOlvgkJ0u3Jl5f18
qLT8sZftBDDZRyiO2CbdpgnhepbQowFcodU1PjdktW3da81aw15lpT+g08IziLNmQ2Mcfcv++GfL
MRpT1UhpaH1fAJUT3sv0zZ/AHeW8DABAiXbUw1Qh2fBP23aFZu5WTlg1jIvKctGuP1YVmw2v7iFd
vPJE0AvXhpg3iws2LACRlXWpqdV275IcaHYkNi8Je+H3eQi4IDvA10XW8FTCcGIuYy1IYwJ8zBDT
Mrs0zFybeZGeecqAU82Eks2oJHxrdYVDaWxi+LMxKI0ODHDi0Rw4mpd5YK+JUneTDoEHWIeI5qI7
Sneosn8m+3/s6NN7hHdrRT4Hq9MAAa5bR3a/+1IaeDbLfZf/PCIC5AuwSw75cQ6Vw+lKIkj4NlCF
XidZ0QCXehA0O6NftAA01XAZtUMcrnmqdJRpl2x48tGWqkjcPbr+MK65C/qMmT6+mBVJeOyFHE/f
Mj1LbnA121MqCG9HQANqTY+2UaUdplr9EuU6HE4prVw5jZD7OQWf5Zce1TmlV146Cb87YJ1DdIIi
wCREswXKsLvCo2nrfnTylVMwo27tK3Jy41TPRJ+aKBZu56aLyRRvX/trifPqKu3Mjgi6tX712dNE
yW9tHIlkuJfAOgHaHIEjiq8AAG1nNdaRougL7UJbNqUgglDaNV5XZDGQsRGfuQpYNa+JCPilIqPp
8jXWXdxGUFr/cED3GAWXoNkfOcMEu/6JvAnSTm80zt4NYFNJctXJufMIefLGkvaCVtS5wb2wq4C0
THBLIaUQTKLyI7lQ+xxlg4XJRkUBVNxR26Jv/1iddiGaqQYzQ0D2i1LkQmzMFvbuboptoKOgVdxw
xUN2Vb5TBkZ+iXxpRj2mMRgBYJEqaDzN//AEt+PrIkJh3twRz1lEsq3pDH+AxKG35KUUP25Jfygo
EVYI/pwNUFtNqFNKpyVLzRyttYPI6NS0f9cZ2rgrJpTUoG7Yst0YnJTSrAxdGy0LEPooRjCkDgcV
cBQ9j5YBbWbtnEyLlRAiuQvryroxVrUnCzqc/XWulA8W7UyggwIN0OwJ9L06PJ25r7+mafUCabA9
PKe6pfB8UD2eHHdruiRXGfW3xE/MAjg+HW0aeu0sSjlJsTS7rZkuJHlqyw1BnkC7FwxbdQ9GSimU
q3k/tmEI+UHF+GG1cJurWiZfp5nS283K7y4+gzdJw9LizYFSK2RRP35pIVGTPb8pD0c26d8Ud3e9
YN3tiubqWlHhdLGQ5puCR+DyTZQVdLrvTGcfs89ukYVN345DFcxTZZ5TM2B+Gajev8PvzypGgIw7
ZJ50W/nE8mfp30oOLnGMQmTcD/9A7GrqL+ZdvLKKFxMNEfIh0o4KiPGU0Hmjo3sJ7Aunuhbg704c
/Fhs3ywujF0hXtCY9Bdty9/lmqCJXMmcSckWodvfXrnB4439Bg/6+ahv4NzNqNw18uulZiPwegQL
w23czSchcP4ImQZLd2atlOBvy6iG7o/6mPrjEDJDXyXzECnJQXQoeyVUsuf50HRUS9h9+41n2oss
n7RgZxEbMXgiCm6zcsJfiDPa9W6eFUw/muJd+eujjynEoS7F5T12cDUykcLYKgnnPJEFmPODNjEk
wJ/rr15DTFS+EzQoMb782n0Sb5+zIfJ1gI8E39ZSweqLYoXHZb9VzdW+HklaeEnbSOIwInPf1CFX
n76a1N/ibcjg6mSfOtv7FhfAT5PF8UePAzXNzlsPFs0FJqEES8yrWWRjS9DGbBtojwg9fjbaWRzX
bWaJYtoP/H5H5ERsl3ojQCmy8+Hxmdh4KvgLyhFKBrIdcEztlLAj9coPg4OGpWTJ7T1S4ak2w2ve
rX0YWmHryw+EFJVNC7iwSNlMypMZqwDkVI5ytfCJBVcFJqOiN0lQWU/LX3xsRjEPVE4LxtRGVciD
Oi/dyTbA7BZXMGHjoOt8bwbzBTSU51StC6UXkRT8+WQFoLQGgfg16h6eeNh7IXXZYOYIVJZk9LsZ
C2jeCi3QpKcU7GTFGItSpQwlVKmbH/5g5iVL7//70cc14gtlIxr9VfpffJin711qVmtFVF5vTPsY
beE09N37xUqMrB3XOQe4HZfd6F87bCB8ZrIM0cSSqqL+ga2UZXW0jvkBH9NznDhhTviMIAMASNuY
l80LeUl878a+jaArz8H0prrOn0hOwreBV42+A0pH4rz+P+Zyao4qoHmGWW1Xc30LKIpVPjlpjcBd
8V2M3vPLonVWyzzxdWz4FAYcUPIQoa8K/R2227CQrm46sk/DQllwPySLRgd46HIaqssNcCZQFFpT
rKrtZe+LcSFnyjuZMsdzA3KQ2mImkX66uRgNFgHc7dfLkaLSCjgeRP7GrISneYq5EoVrJpOn393J
LqEqQamxJNF7P2hlAWgv2O/GM6GkR8Ig/MAwneaKTwMaD/K3b4WZsvSoI6/KzTg09k9E3S3B7v2i
NW6Uc2nSd6VoULCRRrxZURKn8GzkxwL/vRwPhcA9bcbwbAyo+CgrvcnaPxMVNlQ+BNhfFqNbfE+8
JzRjkIaOx+00cItubW1iactrdgZ/xQCncqzfzbL411uh5Wfp4FfGgPq8jjR996ZZfrV9mXLhuEnI
wU4fH1Oz4glXALTGo6V7Dsgx3wSj9GoYsbRg3Gtme5AJavxtr2m3k2EOpAKWXfbCTwfUBcAvcpit
XK7jZhvPfjxYC+7Z+v8BCSMRE20Hm/2WQVZpzUvRzw7lhhWGCNULSG7Ll6zWLKEd8XHZ0T7xH9VK
Zwt9AzjZjTpvCRfPGb9aJIyvPyu0INQBsTLWHR3ijQj4vcyptdpd7jMfAki4lu0Ejb1TwGr3XKef
uw7XIm4tJOd5BFGRh4SzKPh+6/WxhvyFqTYZRiDFj5edep4q+I3EZAHlRkWPryNsJK022ASryNmf
xs0dXEiDY26/GDy9nuIcVUURUTax0L/KGvuA+RZKsPWVdtX7f51Ub/zkICssJkEOwccAXcJOOnxS
K+BK8esduc3KVqsfTLjPPJnLqHx4YE3sEyWbd/eTW+lkvwbJfeaFcvH4pQxOkhVtM67PLgfHbLRr
lBcOmKDh1zsZgjZaNIXRRtXoud+9uLLKYMwEWSinmOgJPfWumGLVWZYncxLHyFUU9x+Qnv5d+FvA
SmRT46l6GbBQFKTXDFm32AvZ0u1yYWQo2ltChChgUMaUywyEwXIW6yBKVAOCGEJ9EeLp48htiAli
WMVE69SnVWsGPJ/pW824TNXDMOJEBQa9XPEA8vGQgZI76qOJzYvTsTG6AN5G8zMinLUTkr/XUHmK
Z/xb4wZebJC6GcATDY0Pr8Kl7hxL7jvnCKjgqnep+gsIxodSsqgRRvK0RiKyrmV0mUkvrjvVDWgA
6+EMEyby/S8CD5xxkjgjhUC+VWXm52filsiHiTaKfHUYVBBdRFlBjOqSdYANffR6kkB9wpBMI2ea
IsmpRxVmxcGasBus82soqqz8PZP2ft2P9A/nhKTzTeAclHqvbbkYx636x5uEPs6AvalMzZoCnLu5
pit630IkWLtOXJiJj5YNXB9vZAQ74HWV4sKxsGtrbjsQXYM8z8TiMOCSiQZ0HA2F55IyXnUvlnG3
nNmnAEmeEzRvhQGBU1GEUrBSifhKyoiTJJnrODUReqwz08Ivp4wC1Vo5jiP0THQfGMybrGu6Enhf
wSRECBBAWmLNa/5hm3t5GgZNP1Oig7thd+hPDATfjo2wfFz547P7rS5b5ZFdOMhfNj0aLG61oZnq
QcuKh3ZoatA9tiYGGQ/EyqC5i3tVY/dqG5ncynW2yxCtADjkoDxDzmFgoBCfghQn3GKMFHH1zNr3
1N+KmEoz3X34TJblaPup0HVJzipuU8L2Rz1MpbsUC9X1+OikTKXdZLrJ4KaAqQxqTMVzUTtfYCeu
pzjuAxSabyLVD/WZQzE5jp6lvWKfe7igihx9/L3tgYV2Cn8d55+hF6JvxLCjHRlCu47F3Mxs7TGq
c5Tw6ild58RuTTK9VVcJdjXbDOC8fKwmMC/a9LlcRo15c9xEmQ6uYysUbDiLioSK2bL/kscSBRbO
ofZQ7MOM3rVc/PFXeEp6gAcOlKd+1yGttKFn9nmbEsbG+ON+vq8cdigwZwcDdkcmlT4IFq4eSx41
fVUMAe6Y1Brbxk1xICZDzf19cZObM4vRMpeJuD55x/RHnJMJR13zQNmCxLWm/KNCeuSguZKQ/2XH
Y7OlQVPjE6UyrhCOaL7i/4F3hi5ggoUxueb/Wd/crYCnVw4eM693k5s2iU4iIbOcoDSK/gOji0wb
Sgwk9i3gEShvak1XO1vY+Ay4eTqvkHbm0eEvdB6prAkOld8u+A/LbicECABV8GaPuuIrtBUSeudJ
HUQVy8iB16/GSz4ASSJTc3Sa0Zcuf8odjpwGImid8nSARomfV3Ug99hVjKIICMcusRRkAWEICbiH
Uthby7GIB7ymrch/PcTOi4dgLDKxXUfEDtjBviB7Xf6x7aGzbdchoSR3u1YNHSWDzHFgDE/TESSN
6sIbLW3/jTuOGa1dbdQpmT+hivYUoNJCgQCMXSkZPb+VfpPFL7g+aFcQz71mAKMzI93/dOmqbV2r
ELT3i7y/K9ppy2X6+yoZ2Ckn5vkUzyNiVnFeIH8O7hgYgPY58HtEVQssfg9CdsS21s5bXpcex+QY
DNLRQMIA/7wG8whdIxmgLvOJC5m1S+BTviGDPctp5msZxpMbE7aJJDD7FuhvzDBnjsIeZCkeBoJ8
MyI0D1TKy/7gXnhssgu2wfOKagGbqy/XPS8fBNL63+WWeQVIR0MdXe0MOZmqkW7h1YmCzHtBTOej
0U2L5dc1hNOBoMWxHGnKioVEjrpSB7CREWv5dYfLEkgCqcRJUmuQs++4gRwf6cSXNy2PbSb+gIlm
B2D/vES9yMjAso9PKtVlWuqAuVTopRdU/PKW2+AymWQ34pLNTuGhCRNMcdy0HaUttBEuXx7RW1GV
jX+WAyc9xfH289fngRB2HzGGzscKvp0b82SBDj8XlCcYU1dGF8cuMGWpISs4hf7VsHTCmZdqMjhh
3YiHf+XmIoxZZYYsmvwWUaexMpcusnyfn4+PejkbGsmfs6g8JTOV//82v4HTEF0DB3wSBeeIpArM
eK4I4EMrObmVTjf6avkrhuCefy4a5ADGChU8eC0PK2uqvlQ3+4L5UtvyxEd4trKQfPQ4N9FpvJZw
Dt/hv3Gvjhlysggdt98cGOtVyosiN4lOtAFgRhWfZ5SM7RYjxiZjVDaHvXQWaWbjwOktYTO61rsQ
vOUCaMI5a8re4QbfQeZmNVBS61OjmyveXjBjpNV7+wowZqlCruMaWezT8kNnICFwq5Ho38ujXejU
vpqjIm/OpR6hEY8cG9So2g57ydfGCsPp6QF3iO/jrHyMLf6XVHoyGbuOzivCB4OkHdexAd1JB4Oc
8XESBptvD1YfPBkfic7XNzgVnj4csW7ZlxeAM23aBGAsuCifjta8n8xd38JhMRqTZXtuPWWt7H5C
rErYtPtQ4pU8LrjZ+UBWmyaMjXlURDb7Q1HNljIyImRdmmaJ/Jh0bQbQvBIKEBH3dTX21hn+h3hf
jOxQmJ4J70uCj+MgtsfGC5oyw5szVsQ6En3SvbinDfYz1cvPdz8375jxBiwQETFE14igZRmafFqk
qkX/5CmOG9+nIyeSo3+dynz7ZQPEl60QW4Nulh3u2AbiaK2blxbuTcDcTuGAhR4WjoFjFEWvXouI
OvUK5tnoLFvtrNbP3noWenyhUsHAJ76tRURE2Nmwn/FBg442dH71j1q+WUQvInyqUDD5F9FcIb6P
YGUFfDpioX4mSsdPFD3OZcswrMEEWtqF1MV5Lw620Pe2z0Muo7JDaqgXzEv4Bh+x0OoN6eUvdBdH
7RnCjJJjR1RklpT189bE4gYV4tvqHNINDViaSK4do4PDzH4TBpYEpKvr03g9jajfgRHQEGD4c+Mh
wkZY6nZs9FU2nQEOS6APwgDvOG3OAZqFhmmaJq3wE0GEsfi4azCM15lkRJrJDlM3pb2IZjt9Dec9
lXhnGOBzvBbAO5cmWukIuw7QVi8yYA+5vP+kHkXFjnrnaAFavSntuSCEZ7EsA2x1PwurXpbasPNZ
PoQYtD2+dZ9yBcXgszTth+kKOKGinCM6P8Q7IVbAONGiZ28Q4xs6cZhZ1JLSL+bSJpMnzF/Ur6on
DRxJDiTQ+YkNEhE7u2J2IVckayoDBkY7QzXlNmI7rtOBK6HtJt+m3Qg+CM9T3u61yKU5wJU5h+3Y
oQu7Ro8PmgqWGXvUWFdJtTDPczpuio+CgSp3NhyplL+iKtbA+N1qZtCqMf1He7k/8cF9MpyKknEm
cumWCG5+jUn3IYPAeBWdcJC+Yr8Q173iO66AmaVvzRgspNMdfsxfK37PWoPJYD6y+ItxT18bCXYe
OlGQ8vq0LW2IJDBe8AHmrlBq7OSJd1lj/ts/Lrw1OjIuMYr/8vQaIF11zRLaOBXf5DzF99fFO5yD
HVOsk1H+bFVkvQTZPu/48Ec1AfTb4hAKCq+9nrEKQeZ+jOzfRPl0tZ9QArMut+urmA/JZoQptgeE
XMT41T5KY0SCthnFD7yntzRHkft5vL4mKS3okRTeFa78++nd4aYT2dnyvYVZQY/SR32pI9z0wrek
Qntsmb8c5jciH1s+xIeN7o4hzuJLU/VjvnUUtkWXyEY3bfgDreTbO8/mFCTrfxA1cCnBOvh1Bqga
aZDZRVqICgWZouFOPJxYs+nQgWeLjVh2jVJGBkgbmq3agHrlc3wtisgFtbFUVYNjgp+7QQxhxGd9
GrOwoVhG06stxbXAU66Q5YKtpmf8/dHyvh83l2+o0WZOc9ZlaFkZcuhSd6p5xQ8fOY8RgSahC3LB
cxYXL/NnvOvgPl6iEjgD1IKc7uybDvHaePjVC/uq0R6bQpkYnhgSU487AHIqctIuOlaUJNivR7kn
gvNvTUFqmtx6Wi3t7iZxbChS1HesQhITazEYjA0xGDPmgREduW3BGeZDTxtnPdbdYdX2OWyJH51K
Z+7bkI0slT0QkPhzl0e3HT3hbGevl/mqJ4Iit/Vsyrh6rFUESf1t3/FnXEJ5cawG5olaoX7ZOIdN
juO6bvtT2yFOiOLojKMVcB+eVnlyF4cVo4+d4uzApGKepJmaO6VSxjEzWxnHqng7nj7POU1qiEJe
rFUwVdVi8Mpw91kJLpQroEb6drk2PcZ5NU1MDlezss4+O7jEojCh/K+Hhpp/2kBOIoNcA8SBesmu
S5jSrXfVZ1YiDRxNheqzbQuRHbypnm3OxrlmwMC29QXJOz7XqJYyRMilJfIuGwh+y7/QpMnk3S82
VBPKB4AHriic/gHWIGsbLXmvI33Jy4OhSfxU2fnQaMKJEfG0RYrWO0GeZv3GWIoOWP7TcYuh/Oyg
GOeJshqujiSy5hbtuEJacnTCrRwGkuHfDLScuMGtjNhS4ojJ55Ur+A1r4dDZOUS8iQ47k38Lojq+
w6sQgggRLSZ4/s7sMh2wA9yePrZMsUj/N+oSVDLeA18n7gmch+UZ5rmxT/tSttAmaELw33lEgPLL
Wtz4kweArPDNZRIkWRbbgmY9F1l6ZM8wXusutA1cl1b39I4/a9EHERb4sLKWDfiUy0ObfnefLzJ8
oegOmgHW2wcUFLSvzusOcDGVMHkiJa62UbHvXcL/yK+e/72s0h28NWxpIUmRNlNniiXE7KSU9nf3
NI4WQTOrRAn2Ssycw+uHPX9Jm4uYIwAaZuPKQK3PGT8pLnTu95hDMZbBcVBwQxhOQ/LR2EsXH+Eu
CRfDnGPkXHGEWIbcdr43tDuj76mTR4GUd7T48FFQ3Uxb/Xci/jNQVB97GMhbUfDYIZUp87j6Ua7C
Eh6Mq6xyT0eY/UKtF48EbZ5hKq1QjO9AwhPt7IfPcTXxsEHoTzj8RAY/kb2UHOi9h/2mDGZm88Ju
/dEvNRQJLmT2u6/AdQnMMudORHvwyRWptfmbajNpy6IQ3uZLZD8snyHqmYVEKdrD0lo/hUDAJREb
xvveba3Iil0RiRnSrY7PAbCeM6jzyNdKzBtIAY/ewclzTnVv63L2ADPQnTIrvo34bpK0AYXkxpnz
/ljWCX1dxasTlPOCCixHwHob2M2MHefOTMolsfYnGK9NgPzhWVTE74ioEjMN6lZ2FM+AeX8f+q+w
OPkbj2PFF4ZMC3BEwWYsCC0va7mwbsgzDoquseYf8PdyOCR9xyavK4ybjHhZYS2kCnEn42yfOgSb
yFQCAo8MZK4zKyMrW7VBsPkr61dC8RKXf6XjFIjvRz03HLDDBH2h8ZOQuI4mBCkTjLcL/NtYhWIB
JhuxEYYbCPt1VxxtZuOE1Gnmf25NhNr77AHIkOVCMtwT4Xfw5xG3f3S+0Pj/ya2vx+BzP3zHC10h
MErcUuJT5KPDmxLrGmWcKtSljqVkoAvdxQXg0RufsscJUI7ckDSC2rh3U+gZ1gT/CPZNp8KK1/M4
z7lX4b2wPtm/p7UPe89O479Sma+UxTP8hgUV/l4OzqiA7LDVP/35aV99esWlBRHZ3cXGqG5FrQbS
zyujEkm9/PusVZGfkLNCllv2MEKIXRX/lwNpEUMoTl+jQEUlH9AvFpJveg/bezjSPro1l/6je/iZ
hzwRJYw7v2pE7l1jpTkVmk+HIOjy82sRQOH+SYrOUZRZRQyY6ZnJUrOrNbfpCIiCfKi3KzEkRkxU
yttrxYTL1eELVHD14eIRNErG5CDIs2jDSk2OiOpmwGyU2Kx1v0E+SirgFGSVRPXciyiZ6J5yyfoM
P14iMUprARQ3LPqOZTlxafZ5kK0Ogu8BQpeikkFXgle7J5rBf+eC+L4E0h2RYRMCgRpnd83/AAO0
3Se8e8EkWLWJ4wqHYLw4atRFJqUooxAuzMqMfWY8l236jOabDIrRbYhuFk9uQqQGwun7H2Yg6qwq
gsc68fR0X3VaRZcrpbH0Cpb6Nul9PuC9LpQYqwyfqSaliL0z3GXAwtVtPIEmSEanAqM2mcUq3vBy
RLt/8uNwkAk+bZbGYb7pnAZuM3VCOi8mbtro9YlS9cvDG62E4tcd+38ou4BK5j0askfGa3CpL/Z9
rvLom4pMtqH2KI7xIEeIi8C7qBd4fkXBJcgUxyasZvpKMKSo8tQQtjd/gABRPRaZyteRGE26wLZp
Z3TDtLyHatW80ruUGtk6gAotW+6kEsVuVqEoNI/wKzv3ZurHE7AeYbIIsG5+kPN6QBhvpPAkCreT
3Fs0DdUbBWE1GqIJ+m+OHvn3diyXCDGu7ZiLgPNscw8mridL/nLBBj9cdUUe6YMzLHVL2r9AHxDA
GTHf7XeG3iDaQRXziMTyyk0gg53DE7JqH68XS0I56UPcm7R1V5e4TlfZ40nkzt77cnCM/8DyEeYV
W04VvcVPV/zAGvL1GW8hQKsxsk11FDjTHFTuwBi7oxsRZLrWF0Ycg9YJcUKlYpmInqJFhtMNvO7d
wPMcOeiKFb/sHujcVC9J+tIv75sJRG5AK3TnC/aaca//q1enE5hKyYcZqt4I8erHgj5kwujrCGMr
tbfZmx5UgpxpYMTzyPOKTeBSoEfHMsGmVsu1foTJS9Ery7w0Lr1g2aj5RQEMwroHQxQRMIJAD55N
nTYLLlSfoQbD6dDsACVuZ/XUtEUxEIUpIJIz5drkj7ThWQQPPr5WOzsKMmtPqpwIbVJJxZW6KIVv
RK5dpbocTr3rYBlljb8EJaHzb5r6zaudeL3e/mpPuPnI4iT58Y+teHgQ+wLO2ueAq2+n8A4LHZpE
UdAQfzB6FQ0FwxRtWMMedsX03PzXwbi9Xt67iqyWUfJBJtpEuOdkznQfKnXUdAYy9T284XB+/s/d
5crAlbPxlAhCKwuaEjA9yOwrrLQ65qtmVF0nuEjyN27EPyQBRZ0I/yK0//QA7fGji6ahVmnVwDss
Q7WxhVXmeSe3IF/PTBupBI6jM53X9hrxZl6r0Nl0e0Tknp/pWxFp2OLsxQOaQteDmMPGheTo428c
oc7A4oroYuwNzEPqHZuIimutwFVI8UKnkYddMIoi04TnoV6VTieX5sc+ykTYvGhzxojYsGasdjoh
dyGMPBrrdWEmp1IzNgUu/RkK0Ku60KqNtG9w1MIWpotpy62rG3tjUonI1zDT0rqDGmamtCRMNTiN
H/iX1/qHamTbTQTsxL2UMsPx79J/o3WCtTqZkbd+qoQg66Xztm+WvhjwK8b7LO70e7RwuOeU2F0l
924Ww2UBl+K5R0D6NdQWBS0Hhd14kQ6lTGqP3xnv3/QvN5kRy+MFnEOUBQ0pX5OH+oTtckPsMQDT
XUogHhzA9Jh3sy8DfkD+z+ZWIkmoewXEfvJmEr8exaPaYDC1OEXbJqh61jGJwN0XSyXIb0Nw6yF1
f/L0GdtjaZUXe+QIfiwjiqEul0Ujxz7dQitTCWif0kQL3DSA0wYHe52mqVFela0O2/YGmU/s5YCD
90NUVXkbjT0QPAsNUFYgxRFu3vd62PxU4CLJtfaRptbE6/WtvYAAEi+S3+9zmwavXpbVUZ27oHgx
fzA/jZmsY/59bQYTlpwz1KySsKFpwaRjxOCvhGvQcdeJmWGneTXEH2a87k1uwl/yOFbb/KqkxjlE
vAR3sZPXh/Lnh453ytLg3la9DXA19OuPTnGTDX/PG/z/z6BTWlsddNu6lWPTeH1S3/nbF6QfBj6c
+unAva7hOWs/Q9xgX4rYEJfHGil4uvxxQPueFgRJNQ/0rVL6V3a22FcW+4JX1KkpEAQIeQERv6jG
q5cKF2iUjT7agFyVglHMIk7quavGZ/BsAWq6IVAu8hmK8aWVY/QebtRVFuZus01gQukg+h/aXydn
w+UMiPdetrYRE1TKNR+NEgA3Kz+xKXlpcxgjXaLlm+TGSlkkVu2hU8kDaxZZ3/CrJcqmznXmRtnh
iag2YPDRTKeagEI9FzF6P4k+BY0olXv9Hef8ULNFqYkomAsEP52qZv32O22n1Tzzl47CAkkJv2KX
dTJEbcB3UVNq0IRYNbbNzlabAKy9MDM6N/iN1BRaLDPB7hxw+/Zy2OF700xsxOshbV3cabE38n3j
1EZhPJ+/kXGZdxGI2C56Hxs6fFFJchGpKr7+Jvky9myECnN2bGxj2eqdYO8oJsotBcFa7n4vpMEb
QcVllWcamIMHtwyQbNdk+SOuOY3OWFPjWeRlBdCic4srd6ofn+jruvzKevB2Gsp54G8t5/fuLbPi
16fb3ocUvKumYANnzFyCNNLrzzp4JDHqiKKT0oJ5Esofn7X/iqzPP5wvFxvLLjCi1QGYAKimYhz5
ouEnTL3eYAFCGvIXpyqYl1/kxcXQWnVIz7Kwp2jnsBcVAinVbxVXwO4wOq0WHidcGsukDAuxnQAB
Y1sUXfFxF3ddKehC1b4KTEJz7xNx7SRRxSWpI62Cgv4gRrwZu0yv3KL5Kd3CnsMJD1l9aAqNHNLM
ULuA7A2NwfyVpLy6XsCQEsVrpdeN8uJmyeaNwcgZisPfRCwpt9HoCjU+RLT0Tf/9H9ag0DyMgiqn
/y449rFgCJBQ9zi9QgKRBgXqqgBoJO7liXGSkS3zQsAv6LtoHhac0ZKiW1gugbqFpKLkzM5Zl3iS
XirYMzDkE+/BtCJKuqfk4+v+KpinHLaZ6xNNNj4fKRHKBO8hc0C+pyUpAER5VIvsrH5lgegQtGvJ
bmoea2dQPzDdZXeiLi3roujej4D2523mB3piznmW8P1R4Abzc/5LPCFPi4+NPtav8xyF14OGIvwK
aIs2zdrcOFBO9l7pb+l6PwnV8UaL7AXaDY2MerU4tnvBECaM0epsibMmFXk5QilkKFoeinAmY6ZO
1M/eJjhQNXWrCtycAmiQe7FRy3PSh9FZgZd/ee3t6cDwEmWq1fMz2kJJlKPAXfYW8duNw9Vk/XoH
TUs/VQYYKVK1+JwmQMftFS3GIfb2sqSgd0CzamR8+xilxME7zLOIkNZukKO+UIiirlyQdXOQq38d
40hGt5UEpZCM1NYI2lmiC494yJ6IAgbOrck9wneYUQRyCElJuUtEpISyMeeoKB+Nd/9ZIp/jiuta
16wBUcLFMaId0LraJABoBKLoBDgpdTn1lNpRVS6E1ds4axIIt3xG7sCBGHLrwubaJpRK3n8hUjj5
QhRM9a9yued1zqIxrVnhAB1udJJtpYPbfJF0HCM4b9VfNzk1OWoGQ3xV7YkOLTjvC07RdE+bVush
BORtTIVJzag81/2JmaS0kLrOa3kn9OBMKsvEJslyQskfEmBpHNsecEWSMna+Bvrc2Lh1p6fkA+va
Soa+hzIw0ynA4qZSlQbnRgJJzMFG6PUegVugCO7Oq2JJYu/kfdE8iJab1f9ON9Rah5XcgB7e18Lj
X2GkBA7F2G6Zma6X3ODJFL3X+Ax9K+cfWhQm8w43ShHG+MI0f/NtPeX36cpo2a9pXbJiHGR1tVor
l9SZXel+6jHKY6ifbmEKuw2Jzhrd5s4vvCLi+caXhrSTHR8YsNdcrnaAy/Lk7W7NdzVRkxe+nxXA
CVDPs/FZIr7x6ueIwq70o7qNg/+2+jiyF2knRVx6aHNnfH30nPXdxFuQKTg9B1u+pVxc+AeoLjFM
9ZFQXrR2flMNaprxrJ5lkTOWHGem/O95Xa7Fv/4JafLzT4/Z+BGQILGs0wFCR5thkLXzvfkkocQL
lcvNnLRBzbKcydQd9mljvBWX2GuOxX6vDUWiKYz/wB5gPZGA3YgA8/CsW1SQ+Qa76ZMDfsEK/tsB
AiwGwti2z0yOsDJqttcOpwc/Pe1UDDK1m7VmeWopoN3E8WBA6Osxo82eK2LZ9Dkk2NPpvrnVYFTV
jagf45baUUmRPU2cVfxQ5iraDY5kqvFONN9x/DtBD+fantr1aFRhPVU7/1tMGuRBuG9sbnNU7Wvn
HV9hHlMIrsfH20dfpcIZwyDterHxPWLianSs6/D9K+2l9s357R24oWiXBR3SnkD7x2mRrMrJfTd9
TEkz8Fyy5qGcnYZe1i+sx8IE8buUOrHmvq8Z5SgAStZIY9wzcBXwtcjrY8y6B02raS1lznG0pcXh
Gxt5aYNU5dxSMdpTiox0riL20nBsTcF5HS6FpyK+GQDsnbGrZ85+7hCzkCwQUETAGnUIYhHnTcMP
dFkpmmbZsY+L/CIUnU3XDhWhP2u95EwraamsKio4/JjbIuvJXEXvaIMavQIjQrCO2LKRCS3/543x
DI/IKDJYyyesQDckcbao/bJJbncR1Scaup0mBeOAcjWgWrx7H6OurgYrP14vpPjAggrKkuKei4Rg
JYXxE20vWp2mNE7ruTP2CCXXSs47waIONf78jocIwuQ3bM7h0RVjP4YU4bEjcyWKeg8AFJXtsyvF
sl2e3/DK9XF7xxve6HpmcBkCIPQg0rMtQLeoCgfvbjzEYAdmFj1kNl2k4SktbeKTz2kKeCMmRbTU
R74FnkbJhWaj28UcP+W2DsaKCgncV92zMPfxuzdtL/kZ48SB4EHHT/f3k5uZ3Mpl96rZuFYWuHsj
4m+gqU5FOIm2b3MimSSqDn2km8ySdkuydroOC/BtAqCHTmsBeHIXJshQrU3KLZbzNbQsdfMVOwEY
3mwNRFObJ/Tf1m+S5uSmcd5J7M37dIV6y4DHPIkXe2c/JCaKoVqFxPluAMASIE9FJumWeeJYuUl9
oiNMa/RjZUNpR14+/K6b8ek43mJhyWiyxU0nwyKNrOBntbxWoVi6gfQUgc8if0ulg/3h57Zj9FuH
xMGMpXIMj3MMb1x+snN0s7LGmDZLo9WDSViPjceH2qTw5CuT7WsWMwQt6Y52GINbPhrkRnV8USXJ
CNDOOHA+VhFT8m2MfB5lhC3YLZuekNZvddvVFIMWfordxWF6rPWbNpEQHiL19q3gDcpvvqM0eXiW
vKnwRoC6jYbn7hRvWKCU0yb5kHkhwmPNvrVGS4hcbgpZCm6aQpMZZKp0Eu1zmslfJWVuKN5h4AJ4
Ot0U2SGsW+cwNHhLkAYjNeVNOYBrpAxqmXx+6eyItuJzc9QkliJoKDp44pWEdperm8W+uRKPsGFJ
XYe7E9IRlUxD5Dum+Fasi6NveUhGVS4ZX1Ac3NDD7n0wWADIGNvE56v5Y8lsiwwhXckB8s7O0ui7
2gekROYeOcaS/9Aoq4W9EWjXKynO4s4KaIqa1VfrFGIJ9Y4BAr/914y+clpWsyTXjasVY47wMPkZ
JSmq+b9DKl7NocksQsmD8zBR8olYV1hQ16XfMy9fOCki5u71zT/q21F8QfqaHuVrDWnuS/nahs7n
ePWbrk0c0236Q3Aq3Ch8KbmRDYTN8jGOgVfSGEUgez/B3asFmD/LfIbPs98Bmy6tE4qWVB6umFzq
GJ53PA1GJfCsJslBEgAzBbZpQsELj3K6BxKd8ZHQEFxG1xbctya9+W6rYHleMhpBX7JzPXvdCDGq
IDR1Ry+SAYf7HEg4L35tbNo15wjNVtXTzaJ0BGRJePBUZi8lpixE20SiFIhDa7sqzhjXCUcS4nNd
rq5/dULK34qg/GYSkrWH6nTIBpdlJ+hkvYcaKsF458hor92wBSlNnjt3FcNvr2VlKm+uOktjiaDE
FOiCs/prxEE+IQUIdbH7gMVCNhZUmB5h77tWkJyTf722U9/Ac/iOq7/Xrv789R61/K8WEc5X9VDW
u+n5MtPk0ASPJ92FAq6D36iaPXXgswrIGZzawLr095Ftmg7412vupTyLknedWc1hWQ/rF4uQt5Il
3F5rPMCLGcQsvEBae9RvLLmjgvF227JL/zMieH1jVM/SWraoLTToa8kAukxGHyQMcVQmrNbpKNjU
dmV/hqsHSo1PuEJjULTLCJFhb6h6GGGFnwggNr7Zjj2AksT9HwgNtlKWiA1IMjONvS2VfyV+RP45
qaOM+HstKPGTakUMurwYeUIsR9q7CsjV5zNua8yOYTpjN3a9f2KOIyqfS/iHcx/H3Xxc70RqYF3A
HSoXu2PXTp6SrniDzdbS1+dMxQZgaSpWPQieMZB2IOkcYpAcakpK2arJQjs29r+yYETe8jE+zgWl
an+Beuj74WHhN43RAIpjQw+QcQrJdfNgaX52kVfkpxSfGgJT8yXr4Q9e6cAFyDv8i559HGnh1+SO
mybbhb4ofI07W5JtXnjllF1J5CtG6SrFipKsQpwprN3e/lRVUIVkDPceGgLbkmOHltD3ZNnHkDYc
YHZ8IGR+Wtv4b542gBWYTq8A46xxALU/VFSqYIQg9tHeigl+tye0w4oPMigW06oeKbbcKiRQE77Z
iL93gT2dk+Gdvk5tZsg+AJCm4O+YwzqKlCSg6eimsnK2XRBGo8Nws9lTHhUv6z3pclS0Cz/J4H2M
I89dVM9n1BppU6UYoQGuGGcXUihoLuzJdAOnXE/G4XySvrifFVhgwlvq2F6pQ2OY7Sthk1ZCNBMw
XI/l7UbQWKlMo1LplhxSFI4JxhChkj6K4PWLgM4B0BEzgNAXkd7mvOePDnEtZpXvEZB4eLsAaznM
jZvaHtcgZ7QXozoB1CMhD4BLBT4t8lWrkWe8znBge5dg0/d77uDBPjBeuIpeXahzmOlblwU9PdMV
awlgdgi0VRtytevCicKfV8CoUb2afSXSB3OxvDbq/+PT+cszNRDm0Gd5qVGQMlm0StHRWyLbMrz0
u19D+5r4g0Qb3qIfNGcVuVXeQ5EXfC92+ahih+C/Qy7YI7ymTQlMsS53u00T9rYleFVmlRWwJ2Hh
hXRw/mmrQnJBm5GZlt67RNCxabq3v2FQ1BcmYx1gnHgDDeuWkgAaYTWAGCKgZQZdIm81qvcCavVR
QywxxJFr2xYN1+xJuWxIB+lHERtuUiLNUfUKEcoRXkbfSOKM48pnsd4GcreFw7G+b/Vn0zGpKmqI
YR+BIy5LcMrGe76N/Ny9DcRuonzTCi0kHN/YrfNBTgOwQJsYRs2mCsM91KX7ZyyRD0qNkTqe0WHh
dK0lahUVN7lcOhOx0E/I8S+LzSxw73FVoPyPc5Hkc7wbZ4rke39Tp4jJk/+qtoHyO7J/C+2btQJu
mZhHNIvsACGj1aQ/i7DpBIMwi70gVBOyFifA1flRlENusgl7JgNoZbj694VcPDyJCGxdqdUOLpGG
tpkpKpaCSixQnv2y9ofnidZJL+vnmOZwbF9DleJJqdalX+2cvpLkDYM2hWFx3PPlSXcrzpRQgmQa
oVmblw1naBh3J9P6e5+In/9SOia3O9RaQPNJCJ/98gwN5ZvOjs80FVO+B0ZEKcVd6DwCcyEOrOE/
DDh/ggsH9O2FOQetIj7YciJ776OCoZDAnmWMDOF42Jn2rjk4qjLQ4iaL3G+LoynnASLtf7Hs8qNp
G7XFyM2ol13jnQxOJgiYq95X1AvU8dpN01lX1qCaPgbIrZ1IEuslERikECdEo4bZ6AP5xuI53GL6
akOYJ+wvUCibT1e440R92yKTh3XI+VlDtCz1GXwsIHn9cbmcTUiTdtwbJ8l9flBJ2XCBeqkjAPWN
J0A2ds0Rcbke846hYuZ15kV3URUIu1PUelIjnQLGQapLegQrpwLO1Bd4ln4+R+bqOgnlsw7agp8I
wCfCymfdBpMjYsLiyEeUSX0ExhoD5PbxMhKQXreK/InM8b9MeKfS0VhtIXAw4pK1XA78Tv5w5EXE
+hnn9YuX9LDg552OMD9hPJ2iBn0M4t7Y6Eon3x7N/fAIth0aPBsd21qQ7+QtLDzhoUKqP+VTG0Ar
TDiPj64nrK6+seRhTaCt+Putpo3rH31NwE7DCjhoGDd8ufyf88EeYwCB0U8RAD3Fo+pl9qvHRLHA
efWz/vaUvawnhLRwyLi0vZZALrXchHNxvPs2csw0ZUkzwUX82NN3zVER/12F9uUWtW2VNESKchTJ
lUWrFjXMQ/2jv0F6YasINOjYF/3CjcjU3LP/B/qVEIatgBmGLndQWN1SqYcgZ86LrcY6Fkzgd0eK
dqdAbDwam9jDGfKJXQMwJ2217MikbKRKfbzbtnQcjwtAZdDGAV629DhA3MUotPBBfQmS4x8FKX/d
FnAW0pltMXK57CIgV9Qlv82BmuQfzX9dSdac29/AkXRnd5szvcB7BlyXoNz2QLcZPbzyD3Xw9phf
U7FjL1kPkGMDRFPfF208PFyXtUwkOYvKpUCcWO/9j4RVj0Jdt9xMNfY9XuUNFts1B6WzF4f1mrE5
p+OUKN0J2fgLmoCZgnX3tgO4bs8iXlmNXaJwtzBWKID3vWhW8NjTtbX3xQiPlWikZCNYX1mVWnXx
hlUMiAu2KXfF51AE6651v83sTGpvXGwtNcngsaUiwzQ3VbAImcMwhemczQi8G5E77+fumIVruz1w
y3X0HUZ6qRFi21izp5WSLEYSSUpGGKLQ22qTInr1VPlals4au2MFmMfxZZgrtikDy85iOJsGhRqr
2VsJjUjwGnP7dNaHA59V3rtlkyAgsI0ajPRAI+X+AZUNQAE8Gxui5t9fkxidPXDHs3Dbbya2Wxw/
gPsyQv+nNux0YkbQuw3e4Ry7Ku5Y7ITyz2qepUvwO9zaLkJ0pucAPh4svWwAEdStTQkodcuyrNte
ELJFLvRrlIZ6MNs9nLxdVHlEsIdbgbNuGUKiMleMcoU9cfexvkCPh813Xek+3w319XtCC6ikqhrf
m98KLOxprYsISNcyLG0U7xVyfcu+lL8EFFxiKXiOunPW05XFRD4ui8AozcyO2F6sOKS8r4Ui3+5Z
WR5lz/vFCKEjYD8EMmSDzzkIuKYI0TFVgI2jsAlDFQ2GedN15woFJNPhwzkcQq18SMZIRPTgSSZU
QKKP2zHUsnI/6H28RG9GO1oPoOgVLFt+Q5szdnN4x42WkUqmW8hWv0geQMNOXrnNMyPece4ZdGe0
uEk66/NAy0BqEm+4JZKUWbAGVICQUCrdb8C1bRNQ9Y78SLvlwgZlL6tIo8QRWmr8r/V5E+JWEPpa
X9UwvawmUrjzevFFajj25mCEWVgANRFIzDVbHhofNGdkC3QqBOPgmYTZtiKRMWOOf7IDTfn6jrlP
hsYMqDCTK7EGuJgB5CtU1UdyHpKvJwroyvqzcexJIwFfoGpXl9iSbS5YMst7tHqwPD8e0PLF3fL5
mVJOaP8eNjJco+JxVMM7OgzYjJcO+Gs1G3Gp6IZByCLTDZsmrg6pw6nfuhylMOGRjQaO0PU+8Ta6
wyL70xYOadtPOIKY7gjBtQAOgXEpY67qhXr7cBLgvT/LqUwLyIzBWu6VET16rNlONFWALheGS3Em
GNaiHo+MNrDs6Fv8xun5gNeabNJFTf604LzIH7P8GQrWru3mK4qlg73tRuTYooHjq2lwmGLxWFoZ
2x/q5uiEL/VLYTp9FbkPV32635ST8S9u6ffaFDIr7cpeQXt7WFvau4bWE3LnckL/n5zgKJwccLKW
25aZuI+cn3ZHHYMXvhMC7B8PVXdDRasFINESu0wFwYzn3TZH6Ym4MJzFfLCgaczk8MNDYB+GsxdN
a0jM0BTYuDHpUed5uT4AR5kuqCwrZpBBss++iCW4Y/LN+ZPonX5psQbjHyaOkcSYEzzAfNVYNeqp
JlptAO1crBHZc8OnL43GVU0Z9aMnAAKLkgZ+rwk+Tp4zJtdDiqvuQIMMaaRfCiEabiWOv761kddA
OdqFUEsy0cs0/1umdA+FGBMmeRUxcr9oLrUEXOSTdBefnEC3I+DGGGLYc49iNxBrpTWP7geJsOJu
6VKTkBmVXZd6wkY77DVrzfBjj8mQW3vF/rLgt4M+zQRg5z4p/MKrzo2LFFe4RKxkIEjukDJI8Wik
QdmmZebtEztDjXyG8faYSCj2JFlAbLb/ykM6Ey0nhpR+veO4wDps73nsUGSo2/Uhd90xTQhybz+c
VFB0FYWILAiuimRSnbcZ7ExcEqII2tl8UClURMZpj2NYRK2Im5exmoZbATvPGyzLgcMpP9V8N7Cq
otAYM799zbXyH1lGsno8q33uiY7Y1ms3Wd3tEOe01p5ri/JRKw5EZfLV8cr0/QpQKd04F5MrvPQ2
j8n8D7YjpQO9HrfpHQdSPp81Qu5k2WVzt54xjqq2DdGM/lNZo+baJf+9jfCOuCxmpdenL9v88XwN
GU2q98tbL4Chv7xYP36K5uNS7N9iRKoqSKMkuwGS8GZZp0B7PJ+XrFLSkR7XzCZGLdKgME0fB+KJ
W9mgheq+8VmKj7XIkiCCtyWEZEbkAWuouPvfcpkJSpblXucrUVEYNzNEx+qM9gygZGLiHGuMmh7V
scORMVDEF4fFoJC5JGVgjCZi3HaV6AF/QyMUAb0jkt01XmjxRvqRgzR5weAUeBc4QUHsH/6QaAqR
eHWyyhHFzy2HbKuGnDjUNvi9RbMWgPzO+FEaNRqCEwuasZtUN1V3g1irK3ECKYUg48SYuEgCwLF1
kDWnqEy3vEoWeUxbGPnmcTeQBZbDRSrPdBdqSH71x5WEvgDNP9OGCOLnzA8eQ9SM1XsCTjWqbISP
cTzOZEP7DIFr4QFL75Nyzg0qUL0CFB3POG3iBGII37IyubQKk22kkAPtTk8CjgG+8C45bpR3/O6u
OYN8UKzdBjxj80ZhpF5vnVrsV9EBBeE6mtQR3v1ibQo+8T04Iettuva/QRy6NK+xm5qZ2anCs3TJ
7IvUI2mUKuvhJMsK/XYMqrqeHYZTghqMqbf8SkoX471C4jWl+YxQ0FrgS1n0v/6bGauEmquu/6CV
0PyCK/2UWskSZzh4KFXPvVumhZlHJXvO0jeeDcq+VjDzALpgX3fLntmdOv73LNjXcdzDA6g1VqVK
UeDrZnybNhtMkVgqQ0Oe3mC18BLXU0oYzgqgX6CSlnWDdWyuYsVS+AWY2prVNU4yCIp1ypSoeDaw
NjfVA/KylWx5y6hLtkKoKEhwifPIiviUyMRI6YhvcpN5XCkvcWqIvBWG1YJ1nacbEqbzq0qmHDkF
qhbeYNyb53EWIJjcuoAMvCFfYNJ9oERnSXGoAeJqhNCuvMraowWNC/IHMcjMF0y3pISJJAlXGKwN
llqZcFXXK/RPmmp9vUKiJBlSKpTCoXWwDjdlRK+m/FYL16K7G0JvEPFWBxV1DPf13ALqFrnMS9pQ
fl4F/GNV5b8uOTGir5KBhYVg44DgS8HlS5hU8zb2VRKkQoMbZSjUkHRDVZ5rni1nPe5dfuuS3t3w
2JTTnNp+lWQLW66mjnixa3jLeyU/ru3atm/Dw/vf+8LkPQiOc6DyFDhBwPAKwHFbQA6STiznyd6n
Z6vLYRPRWz1C0Mpf3yboswVZrot3VXapOItljoYRv5Wl1i9FZb4ulqTGCIg6xD64fMMUuHOm5xdh
6GF111bth2CNhRgGXEK3oor6aFjFllAj6Y2PENvPsX8s3SRjVA8wjveBN8PlF2zjVferJ0NhwPdU
rzdG9p+e7ssNTRu8k0yJns8Y/g/UmU1vKsUgvP77Y1FEm73oBSDkRWvDjdD8bP+NC27lDm93bDzO
9brYISsjPYKeGEUv4cjyMw8vPk96bJsQ2dTfS3omy718ALvdo2+Yq8FHjfYHTkM6tzjCAub7vuPo
ydS4HKOOaHlC4GFABirWL/PXdUA/simDlZ6I1NtHjqwu5A1Hki+/Sg0aLGhMU1PTqGI9Wok/wo1M
nzuX1DP5t6UjxkYZJ8GdBE6fxn7Qt3YxbybuXd/eaIswAh9XqEurF9+g5mt2IVx5KQqWv5KB6Nyl
4rGafXrXKcySbW7NTaEQzoHXuUU3f9gVaL6XhcxU2geJP38dYqVey5drEfQBvES4AFdl7k1nopXN
igqmV3aMQ2XeCMYIYNCBbafIqA8d/zno/y+wjn6cUXH+R/x2qAZG6YSnw2ASJHg1D1hD3TSgi29A
9glu+JF9qtguN6VxRBDERLNFx++bH7cOfD1pTqU7n1L/k0zvx95hOGG7ZDLxXiu4Ib5rITUzSH/W
7LJEEC7XPtJAVk4mE8RTIe6LKYAQFbLRGzEq25PZVO2jj/Kt24GrPpbI6l3QQZq8SOM17Ce+tMns
RINZqcCFNKw+ygiF41xsu6FykrQAhbmmxRxKnAHjfw/QwauJ3+a4Crw4JVhJY/oDBy5F4rhh/fDV
GnEPQ5Pnkqlu7STgJKWnLB3k7MYQ9InT3khsAhGkMnNrc2AH1/1BKxpzMXimGB6uMSnixw1ENoEj
VpMsTcXjfKb1Fzj02098OJHhzSpQGLCjmiL+x23CN5o1ma8hTlpAAtpBJMRcvDk0Dl+ZbNcLrno5
mfwVX03boUYucklEbS70e3ZukUVgObRbLNfdZVmNSE+NUfMB5QwrrtMY5vII/UUOc9u8xGUxIK4e
7e2835DIOQLh5rkJUnnE+cxMVIdLegerLZZoaBc6ASVV+ss5mkaEE6h6+If9JzZiPPFLEq4Ugy/T
nh1B604gQClySvDQt3aEefYT5S0cHJcI4CgnW/TWcLRTSUR7EmoFGk1t3hGNWNAujEACvl+k6/8B
YW7DFXRyBTNhxwCAaIJIwSDorpLAG+VQy8pLYjnCyd3zmbGlwBZ2WEi8I44m7e+oaEiO2xt4RJ8R
1KoCxA4jkFP/SvbwP8tI1RWBfO18Cdl1UMxahMPtS3wXPyYgAXSyC0IuKpfiXADOAhmOUmSSCysE
OpHYbB4ETVtOZp5gSzBFAtXiwQIRGavO7js1w9uz+4/qiAco675GJC18RxrUhXikDsSlLADX0pbz
TRhEFfZtlOY92mvrpcd5S1/ArNz7KfMtwfEVST0uJqYd6mBNbcMDBvrDPCHB8JL0FFx8WxIP/oos
oY45pYJHefVEgHjdWyInwSBeVaOhZB8ukA1JtZMeY+8QCKtyktjUMaTia7EmoI/ci7/4WOttyTqY
VijNXqxaORFvM/jMPpv+x9VpPnMv0IWK4q+NyIYflMGheWkvsN9r+BaoX3nxMwAe7MOFOdYPW9Qq
xwv2F4xIcsHhIvgidFj0XA8mEn+LpyDFYQMDk1H4e8FWIRlWLOOlVtq+5dPOeELaRDhhPcPeulj2
lDX9ufLKcgAnZiR0qftSIKKPEXSBJNBVvkwwaeftRKHvYd27FMo8iwNfFR0he1KKHHRBMsuyB5y+
a5Hgv0wLridh+bwpzrp/TmdOpu72vlJmdLiY5QBVjLCLF+HHuU98KII66xY4ucf4FW0NUMne4Gq7
TfmhAfAIMj8D6s1melDNB4PgHoqr4C51aN5iIUq/vlifmkwVEVqMAbrvX+4oXkRI6ASlE+Tl14dQ
Xk7VjVrNhI29yyw8zoTb0ajL3+/uWVgT3KjI9oA0dJL1Km/+xk9SEMxOaJK6uMKAuyaLw2dH1wL4
CAGWNU+DcpKtw0i5W+BTlMwDJSnKZnMoYlXiHhqXe8Zof1VQCHEn4TNZtJ4zmxr6JwlLzu0kCVF4
lBBdALH+zg3eO7+ohperiPSS3KWOdLNftxs88kg068D7/s3gzekHIwh1IY8g9iaTGDAg1NbvhwDM
Yb0R0HTvYXBz6Q+NUMAiVAXo7BzwipELAQpQ41aPlyAl+FfTp3AhV1Zag53RndT3GLsh+cfdfmNj
fzXLgR8EHfZiOWHW5NuduBi/qb4SAUKQ3cPDTSs1md05ULJjaVG/+Cbe0nNEyQnsJ1+vU0XzhOli
lxa+6V4FR+IJ9SRd+vyoSWXfOIM49vpQznI59fz6Hj3DoOD2l/7jHfRv+GMr2omEjrHLUm26DQm6
hDR1GuOYb/HL51NzNYIGJJhmpkCC/tiEE0JwyOg5O/DiSxMfJ5NpJ27xzE5Jz2FuF+97zg/H3rwQ
fPHa4RlTnBRiTSHQbZDUeCABr1UzHRX5EdogpPw/u3QhWyfEYsjwA80XE3DTJQCC2ATQPpKB/g1E
vakPwbLU6SqCk9F/Ar60CpSOjOGL2kTonSFJqSSJxghBQsj+Jzqf7qLhLCwOoAt/XS9q/uRKXt9M
1f1Q4GKK866nXrCWt5F4OboUYdnmZ6JISXoc6KRiiH4Yb+/O07eitXhL4i0be85EtzuZSS4YgoQv
aYpj6NywL2FWG0R2pSCNjfNuQDvt3reBSDMafUsHTxFtsqy5Jb2S8hMMC+UoaSHBGPVqaKKABD1l
GHdFrliJtZctYoKMbZThCaAqMi8oEZfH0SQ2/ah4UodWJVQ5MqjD6gTjhP7Dirh2v6LHkkElTc07
EVNuNY3JbWuFh3OhT/kyn4EGA5mltBUICG/yMp6nNGd41fgQ09Y0fJau+2bsOqsp7NW+Wruy3NYp
VgEVmqtKt5mhEJi4DTpjBUxFVUx1Dw3nqnATe8L9ptqbvuBqBANyNbvZ6emQ8+L2rdUSGJQv2A6m
grfdicK8yyCgCzsC3rhmN8YpDVdtrplYfEdLPqS90/FGPSVGxxGmM2q4bA4Qu3W/M7pZvprQVJ7G
C4pDl2dvc8ClH5SNCBxycv7Ooq0YUReuzEGfnZJC9nfT7qdtRI0XeHreWV+OKJzQIYgWFbzKiuiP
JcQlDIKMhp6v8ZyuFvDEnxpwopwIP2R8xOtens8G4ajojHpRdboDU/wjaHhuQPR3WNNCxEDsJRjH
t6w9b8Ynz6s6fNCo8seVPWMAtN1ihE+aiOSqC6blVajfLACpdD6pe9ppchbl2pJpAGaR4KrBaPma
HQgLq+LWD7kVAOzmMG8yfxjiVP3EDOOscSalRIqWw2MS+E3FdOCPaL5jq0vqVqTWlybsC6JfZpKa
CjR63mweXRO5Cr75RDBiUAmfilaZx9JIIy0DFUJdRuH9M8D4JaghbAErvmxL5V/8NTBaotwQIVsD
oBrYmAHlxoYSMOSILsY4xNvY+HUu8/9C33WudpDEPKB+h9zvVqc8lBJW3qYcpMHlvxLv5SQj7QH8
m13rxevJTN3VS1mzpUbMUhUJ+plSZEklJ+DIr6k2q2iYTaakns6ZKUhMXborkMRC/0KQdixUWOJv
DZluRuVcO7WaAVWWTBrJ6U7ughYHW86PbVGj215RKSe1UqHwrIpqMh0yrc4MK10XdN3l4CLzfAxx
43R7fqCKxThgXs97pXI6kE6/LaOLoSix9a3f/S9JCpDdfVryT0fqBOCeDqfB3pE7OiNaFWmoVHgN
yCsC/BNFdgpN/5YgiHlzeZN1Gh4HHL+Rbdjhl34WRChtgqPghUrHcgxAwq7Vs6HM3GQEbsdKHnwg
/bERsgEjt0WT/8OpbxaXCDYTVeQcx7jdBAnumqam/VgEE16jpIegVQdj4GGlc2vVMvHZATgNsA4X
YD77ZCIbJcDg0tRzP45ptwVB2nfQgd64zBDQVugCqi34RIwSiti7O0/g3kmZN4a8olgbqSiDmgP4
DNTVRpG8CYRsXQWYhk9B/45+m75doQIEjmzcPM/0ibBOC8k2dsyRS/lgc97GtPINNzQrJna5dpVC
tQVxLd/I0miQcP7dbY67TeLS86KUEWoaOfH8qbHWJ5xXfMxuDAKLh02BbX2be5YnVmVWLNUSZYlS
xbN1SrRTHhwlKrDM8qU4xJtwDvmli19dTezkPRGAkKKFEL0j3IKI3KIq854GdA2hi1HXdvUyzMKu
AhPGjTmjHfeQF2S/FiCWgbXWvfYJo+ktPS6dZ4iK3qmzmkAyk6W9z0bWQAv+JcAuGfMgyVXIb3VU
LAIkU8ZUl8Qqwz8BEnqjLJccDt6LsmZ4BUen5Mg6Ftlx9h8IPKFmPiVyMWrL0XxOxeNEh5lEVpw/
pqmlHY1UE/i75A4Zq9ew0AvKIaMNaHPGRNyd+I4RDLxu2qZ2HIH8Rpgf0N4j8WPg0Ppc8UXatcOR
eCNUl559jzLlc8KWgNcw5C/H6l6UD/LEc6FHZKEWVpLsU1UNysdt6HZL/PtSgpaNHrRz0o5hSxaS
hGqtS080oiWGskRVLvPG28+9j37NVYJb6Yu2O+Dgf2l6CQiPy4jVfMqybmOoIy1a/HSoTmCm1cvn
MYSiw55pjdJ9zfvXxhHjOLHpabBiSfAFyXcz7ECTyXqNu2N/lQ0Raq4JzBQ0plaog+91NK0s639w
MtHJGrhTRRMmqC0Ors70BqR9JXtvQ3I6TlKGMLowN4kSF9LMmgmgDHw3RTnKI/DtBKOe3AO1W8uP
RroCM8RhVxQpBJsR3hfYJgLGKb6VhABEJtm3tVYBR98Fgpy/40JG4SGat2ctbktR2hF3SFzGYvql
WGcRKNJ+kuyYsCRWQYb9R3Kb1OhI7jBTHUBupJ5RZOCeYCpKYDXH3GnAn7uesYJThf09JFbqTuil
3sr3f5lCmCi4krdGm4kQgM/0rv/ul3uXl/R6ZjH6vuFgnDWnNaglqtkPnmnuhGy2A94w6PoQtLGD
GRldh6btXEaABti5iLPmdTXuqGgy1hMRMVUTpsyIBZJXV4lhIukPlKbdk6Ppq/IQE+VT8T6A+KJ5
5+zhtUP2EFd4DftUhnWfSC6+tRTImaxk+kg98Yy+HrCvdZ007NcNXbpOKSH0LIz3G73fDgZdrZ7P
CLLd644+b9PsApBSPzNZLIzEqxngMnf6ETMx/3EOti/rgmrS+XayFPPk1sFNY+8WBt8lBgL9Mk3A
m+X+NoG1m+XJRdKJsdb9TtnMXwSHnA6ulx0udiDFHMV8+9Ab9JSPY54SQQTwrW+yv8cZvrF5qaGR
kJDpBL6Als0OGMCdYlZYVBmjS2yHyDsCaD06lqAaCm4RjtRWoh5ahmzGCcMYONtPVPO+xbie+lTS
SFczNtdkcxvefXNznvF4IdcuEWVAQSNyIXBxZPlj3eDEZ9cDMZCFHDtSJNPrDJOqcyuA58JlO0hk
N/4f+B3Iq6K5zIMhW/4QGgYpGCvw2l9XY7e4i5LJXOxeq13QHAsRwyUSz2lLrC+CNSTlnJhkN7y7
m2DJNiZJ4TN41+MGueRnVPPOmMAeTOBJl3IWSmP8CwaCJ/aP2MImTC5PGFCJR1wUI6OPWQkfzx9A
aIECYmMlYdi6FnnkEaQomdRyEO6zUuSjc6AkYyPd5MNGdZHKppdJ1v+W1EcDIm8IUN0MQNciJ20K
pk5wyr90Q4tIfNyS46devfXfY5pB9FxpeakdNifxo5WLQPDMthgmTamU/9euk4zov11QwM7GivI0
nzbgQaJqTF88lR7Z83XV5pEWkxxHXjd4wMY9Mb8w+QN/aOMDuMRBVajNTOk1K5IjtvjIX0yzq5qZ
88M23VgrXZyAMHSyjVf1pYa8SDqIaMiJIHLBHrsIwMrAVYZ0cCmu4XFp5dRTl3/kCQLUI/KN3BHg
VdEKVD89wgUoX/F3INX7Ya9wywTia8SJwwx1DUK+ro+l1lwekcw3sVyh6FmyooA/EIIbMcUYcxYS
6uHheumP4yiziLERft8xfwWOO8tJ62ZBAEWwUPsIUncylbglarxVs0qm+VQfPPXbEq+20Jm+7tQn
uE4dondxLp7QeSOVaL5SbuCacJgYN0Yk6B5m855lIynLk1Q9v4/UsDXm0LTLqfIv0+RPTVDxX92G
6MFzxGERi1ztKRjH2T9zBRhgpMyrxx0CL3xItiy9IIGlcQKJy9+YnT0QoHWFzf0klA5jgDPeBJMW
M9PxlyoY2XudMXPHB8TzvGUAhIAjcLzNj6UV/qyxGM/K3LbpgJ8Bi04P5D+rPboNRFrNbMhe8LAM
VAuRTqm1WgJY9Znk4y+j0fUh72EgVY5L02pWSQcCCijj6qXDFjcxjlIS1cdmNHX2Pl19VpwVzkRp
lXS6ei3IhwN1MDPxSeU7ypV0Ecgta4Uzq6y+EPzjKQswhK6TeVHKRHkfRasK2upEoPbw3aiM4tlY
Uv7PQxNQ25rQgTWbl5nOjs04U6YjV8g33TnFhYd7Y+/LZTNNmphfAqBBu7NALzDs4KLbOgTn07pz
MXYFf7Nn7D6AUcfd3CeZ4bKYRLDPcLwIdD4q4igcjkTt6GJh2wTm4bHrubYCvYB/1tRH1o/GiMne
7fGaGS9Ht3ny6fDOHXJnHzO4vLJ3WLc4yMtnK8r2qz7H8kCM34DIRFS6pRvLTuZ2JkKKLaPMUleH
5CjDfwWgaRBLp3CF5Xja+NEwOHN8mna9qsVg5ZKXairUpJ1mGmoHIlnUa1uH2mbKJcyXBVGVi5Gp
QDox9erwDcDD7q/0PP5X3pj7B982+f+GljcFRSemShT0zzlZHui1kpB6mMRaY7XwIHppTKdgRvSN
tBCHsM1N8ZULCDkcCuj08ZdHtOg1PAsw16Ij9ZRUkQCZNikS86PGU1Acw/zCojKDrgQvVJt4EWnn
AWFgoOf3GTYHTFG5qS8sX8PkBDbVgQXwWa4Q5dH49EZQDtYLyBTNYa/MVv0MafVF6v30UItdxWbo
eKV44YYQwW46hE9067dihh+CG4i9/Tk0fUsgFrFegD7lCb7qlYWSVLEN3gofNoDMCKuq3kXeOovJ
lL/gohYYCX4hcuCB3SdccurWNqYzA8Y0JfrQpR8FrggjdRXpV/EVxheP4emYpHosQO4HCpkrRAet
AjXQzLr9BJegaP/anLOPn4I9RGxDyZjIxh19xtcDU7RLOx1emupxh6KA03vhj0qbOKdkqiLvcMC2
IlJjXXjw/w6eLsPxJpn1DuowbMHVHpJghBiO5xTfdAA8RcJfWOqKO54G8eV63kts8MitbjWCgb7E
XQGX0PPvgcx5L987/rbuvEfd0z45DZyxz98obHpBWB79zS/wxcOWZ/RWiEfQ0crMwDGlnnoRgI44
MZLNVVG7oGs/sk9og/D7JEXfPtjLYV9HR2GghjpEiGvgZT0nu43bWAhrtMOJY0mj5U3hQ/ONO3wW
XY9wSapWe8Maq5uOv1dz5KRO/ZAE6MTd5QlQ6kLIJgh9CjHJ+CH7tr0oezN9MA6dxHlU7yYtItf4
uPWqqb04nSjjoiO1GwX7VpWOLT4ML/3P5uYt9/tvGM8To3bE7hEfoUC4A0ADocpLL3On880TH9UX
4d9bSG2w9mpKqSmVo0lUM/UwpuVjepCIK9AVCL+T7zoJKkO/2UTK4ZTSI0JmZUrJdcmV3S0aY0Dh
RGwRtBNNwiA6TJ9ZiovM3v9WXu2lQKVch4/sWw1k
`protect end_protected

