

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e5xVIDBGzQkhDoQ5sfeAF2q83P6A1Z/qsmlSYQJY5xTravGd4CV8IrniJyUa6zNomwm8ijfsSBDZ
3Cv5fk91Hw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JTncam9YaU88Ye5zsiMSZerKzQZ8ndV/jFOlVBJ2+1NMrth4ym5MZgOOJUn+hqDs7WawEc66qp7n
dAXASYJYn+qFnCtyUAhIyvGYbamoaDWo5Ex6WN67wq/uxVFQHJyQE9mBWmFUuyQbfWAxdn0X8Ddd
XBKhuVWHjadjfvTndGU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WysH5jibOCiuNoaEF/J6UEux/f9qwkqszrQvmOG1LAQguVnzJ7+cmZtEvDLaeM5SMkI/c6AvWtXW
QAEuUSUqI7fc7s94OSdoy/EO2eWxzu/2PZr3+Vm/RDQkA2VgY92Mk7iTSAe4nvupzjwLJJp7MPFn
W0Qp6hutV366SMmocbalqT6lFUEm3BdJRb/waOPaQXsiK/eXFOfDC+OkXBIeDSI4U6bTS5BbTI6J
pFf7UmKKQ3+TO+1O/Q+2hW5WOgJzIUFjgYlL/k7HV9GLoiTkFeWQv9D4PmITDLLqEoJBQEH042D6
w9tSjJ90YaeXyJsQBc944KHiROaj7JIGL9ptSg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HfnNrIheX+bmcZCjcmnXLaiCn2W6T6H6Dp6dScskVGNGAylFhqrXsMMXHrPiUKf5LFkT6rGH4xNt
DnPlwzwiCAkQpMo27mNuJmSmEL1NZn19+z1IhIkgUjJMK+DU6V8j1HJvLoBzdBKXeOfEsIha7CfH
SYvgpUYxukUrvYeSdDM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FcdqosqcEEFjwfToDdg81IlS3kR13BUL9UoyGE7K0tYyJxwBRWvuEZwjlqyLvEdW74UEcoL322wG
MsjKrbrYQdHQMnu0VAIvQRAp+YUu8ZY/Amts9d4uoKQ4ceZKPNKKjhA2gLCTZlClOnHdKjhfnFhg
C4vFlIgGFFvgy7hYPvMYgUjBeujuUeMJVrfDQoBe2vY01NCaYs8PD38+MZrB1yBWXtoIH1Kudp5s
6rfzNC3iiU875HSyCH3s6Fgf+5qupOBLk1FOGYXDOgVB80WiCFsXlSgDSubN5g0HTJQJ5d2+rdH3
3+ADIpk9sqzMVdE2qp7yCA7kfUMNWwWOq2rtCw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15872)
`protect data_block
pWSht0rRHYFoYtqT8I+eSaCuA97RDyK0WxVz7oenJEeRZlJsLqr3TqrhKGwgVZESEt/XNmRwJVXX
kVISBi0ryLs8cpGBes8eTurpgYYrTIsNvcGB4slBLHHa5gfe+XyQl6rTLoSkdypR6NpMzE55iLAH
6WHrE73IBrnqY0n/m6A0Rv2bHn6jc0Qe0YmI0vFYq3qNe01KRiZ4p4Aw3WhV1hAhr3LjL1wfwUlh
RXdiTQPWc/RFKYqejuMg47/fM0fteBraIz8k7sI8U72c7YJmrnqmXFP2zy1k0rlGq8uO5nJnehR8
Mb00d1C4mQkNUML5UBAsAENaQ5y8ku2H4uB9wFmJ9pllu2j1+12DVNSzOz9+KNkO8AAAo0THSfF6
kcrjR8KvTj7ctphMO7iysXEA86ol/Aj0vofci3YlG8YH0f5f+XeJ8oJ58s40OVkJtTB9L6s4ZVTe
e1217BihWw1zpoxg+x+95wtv2HHCxxU8Qlr8q57IDu2qEtEzdw1sHS3n9CSukb/RnDihcUmRyyRu
FYxHUFpleAQNggyz0omhXXx/XD9TZjXvslZsBB9abT1WZVrR6SPcbllbo36EKSIZUOSepRwd/3xa
kBrdBlhkjCYCd56BB1sZARBf6XHnH7c0lfKf24LWWotQo9XoHTTmbu4iv2yvC23v5TQPMTtaZFGM
niOJMreOXCU09n4AKijDkozXoKvgB+24ajOnmZ+NSkFR3udk5pDRX1phxGcbv/WkVuFchSc2VJ0m
DJnqfeyfDpckSP+j/IQ7OSB69aQxfnTxTrqOMCLqNMEBin+ee3zxTdQB8IJ8cKSc4giJLKi4nQMV
nrm3oitKqqDX7aqyVgIKwsiCF5uvEZqNgXNxwja9bSAc0GvBV9letoUbq1TTUwiRgY/cDxmrQ5qF
yc+jjWGQY7CGlTVVlk/TU0QpRp1fViCbbSKi5hAItbWjIyStn8e0EcnUX8wAXYWXG+oX7jvJRsXU
C9c5w5FSt9FrcL2Goyu5s6skJUazDvmqmOA9HoCxM+tLhK/SwavnjifqMcA/ZeNdxbJAz42Yc7Oh
BGF7FVF90tKZUcPQP0qma/lyShQcK078EBwJTiQXsxp2CPqYMwIEnzMxTF81RyjPXL45Yu7EZYMM
391Pb0A3aJjs+w6OrnqE7eAhQ45yZ6iHOL5HfgOoglF9Engi+pVHJ04O73/gqLQ8MzVSN5AXlfjS
0mjalHodHElyW0I/6EMXn7dFy2LcnqSA2Btj/5Sk3Iodn2s7Rs+U77dq+OCdGr7Vnx6I7J5OksGw
woWVrUvvau4c59nJu6Hzj2L61BjeymZ9ijI6jAMeZkFrjM5dkmPBtTVYWkYuqHE79JYTToLHf+dr
1Yy1eXI4MYyNYboujN1zKnOWoAOXBwGTnBv6bSJEpyH6wDC4bf7znjyK5jtXFeNzhCnafVRDZxqN
yz1B0BoJVEHLW47IfVa4um7ZepI8qxR5NUIavLJvRrXWHEnTEzaGAS1xBif/iOFWsmCte7txGl2e
Vn6VPy7kYH/b/awtuYulfjUWIN8342+MimHsjav+nMsBKIh7sMy2CIXYZrSgDE7r3oUrV7HjLEhO
wl878yciTNNIIfzUtcr6MQuIH/oQa+rIIP1jrp/2JF+Yf4Cx9QsDaVM4nyvEHf8qpMmkonwg462y
LdnoRMxzvdcbsXM6PLhS7McFgSeRsZTY02BwP8y4dfVsuVTI1rPnT6AftI13lhyDuIATCRmJ0F0V
2Q+Gh+KCWqaJeQWqXVNFt+zesTEb19iLuX/Vgf7Lbc+GRurrjyh9W6Bef9h2/GULE4Tzqljf3QS8
9Nt3bLIlDskK+XmaLoPJqjFhE2gnylLbn1qhQKnIZ7Koa1M80AaX+dSNN2yYGTbqzfZzsRgsYFFh
35LNCrc/LiTnrWMge0zAbYjeK5MdkylvB3ykulsj7BBbYIyTElj6XhRVed2fEclZOoUDZgdiMeUY
BBXavc0tXl83nTjBk6KwXFHoUkpo9XIDPBM6CtrfOTR9jibXN9VITfG0pP+lSp2iLASZtXqfgJic
uNstGb3D7aTTvkb+4reTTs1kil6yqJb5dn5pEuVRziYMIxleH6HQYg+8mxc+vR2Hohe1HU95ASp3
+aEswtksRKPk6lwPabIMtkuFGcSgx3E+IOpGlBXd2ZuSeyqBUE0pFZQF88230g5/c//DPNcyznSd
aOAI6rxqxp9U9rkHmjPDXnzBj4y7UWzImXSvhSKv8zlb49WLm+2C59HL6xvgpB1YHrgYM5BUmZJ3
EbWHMedLSP7WvADfd2+7Nh+cGIEWvvbKD9HsLVFe22RpWjnuEPfW5n1rsP0ZNHP6+nCR9UjEYgnW
by7cAiZKICFbboNdkKldqEUy+akH2wHTM4nS3Tk2g2Jtkttc4qAsSr2k8/uhNLOWvX/UvNQfaMMy
KoEbp1YdRQXNXGzBLKF0n0jS1V8nD4AKL9fwuojgW9NP4Mc31PkoNNoP5Ohq1EkWfeAva8pjuak6
f+VC9ZXMCYTMn9LHqxS0qlMTsip798MUHQ92sWh9zCPJXunC68RggkRDK3R1G5+7qF0VyIKPFnOO
Nrky1sfS8dKr8Hc8sCzn6eUmgAbFW6rWRoe0wA3/LO5GVEmK+NTvE2rBBApi/8/Nkly0ua8xEC/D
p7hiKzzQSG+547WoE5+4mHkgF64BhVmKrhT6lvPlTPQ/EaxGHvlaiq3mIz8U1ZAie2FM1g/PT83r
vuTBzr+nGz6960Og3jdYKVq8qYiOgwAP3v9MCi1E9k3dex0FARrvbEPkyQhuEh6PAe3tjt54E1le
UG8C15Oc9XoYoZz9pTtv3yG0wKN0qGbliDKRYNX0os5aEYDeEV6PY7t0H3GL0Xn+iSSYBmTi8Uy0
zAvUHI1MHds0ia5zQVnVWKPXCs4z8JPcx9E0WPcxKkGrkNZ7lIDiw0BIwwXboCo4H6ZyPpDagiET
b8/0lR76X5YbtqE4jSQX8oyvEpIVukGOyLH18i3mRm7Ga5cyouBbz+SksSHvxNkmCbHYa5hRdG+C
ViqXUcKexLdiEKieGE4FACj8qMOR81R2HyjfTeqh5UI88JgREXHZpMmnc3yN+Laaxow5w/f1cD2S
VEmY+FQbmm4P3ublhWrTr5vQf7B0m0Je3ecOVJDEa/ZTg64As+OZVhl/TAFkOhInhktJolOt9LIy
xTI3qJZklCguyeolFleCaGreVYhSwVL3ccBmJLg5aSzZ8yxf4VS8sYM4xPpXThAHoA1asy2E8iuo
6ljYXpZpneQc1dTq9gPiCOo8PST3smFL1zTFx4GMS/OFgnLWKk1yIDJEREMD4bYAiCv4JY6A276W
vZMo1KiyQKNoUE+Kt02evEQZXRW9CJ5J4E1/wQflnyQ1t7Tu1RbBT5RJC4kETP1IqqOhpo8y96zw
mF1HIYuvMcZz9TAtP2j3woTX7VDdNf8O8UBy18cOysKiZxGr5ktHRWkePuoILjAvI69EIVHkBV+2
ZEfAPU6z53DBHZmbr8no87xgN+qhfoArqIreVkkxLJHR0Y8RpXEdp58ogLxiP/T7sqQm/KuieEyD
XjhM9ANPBoZe7/8H5Vgk50CbkwBtJKGmNTziBnx2/mHylOl27NHtcOaKTdwW9xDrJnJHGao44A/W
Z4QLCYlRSoeo1dNnsPqDJzqrL/uPM6kJ7hCNVy2ItqASzC/AFVNNpDyr/1NuD45dJ7YqSPvZif9c
5UZk4Imt4nNk3H5WOTyMbfDpZNtiNXBjLhdKuSPBlXl8J2m/LsTkfO0NhilmnS31/XODEAMOuXHx
Cf0hHcjAj9oQVwKnQQiUDfBx/s9sDEzMsluV10ApPOSkNpbI4gOiMa3g7ZDDIYbViQd9AhQJGWfl
VK2bFwx/NBRrU3zW46B+r9hOmSwBd4FncVU/e8dcI949fenE2f7kuCGKi7nbNSY75rIzQITIXC99
znywPKx2DScqhttYbqiw8cirQjqV5tA4b3MOXsWQfBxIkE4PBvITGtYeKCziq2BPAHTQhUBNrtCk
k2QCaqt41U1Kg+zenIm3DpVPIK3oyfkB26/jUDYLLsZQclvlMGhs77Fvj6PiLan8LawzUrnalqBA
2uHwRMf0rd7yNuSV6B2tDGKp5G9BbMtY2geJQLBH6etkvKfX2tx0vzREN1VSPGsGkJZu/TzCDtpC
rogRTYG9wdoK1zFSlYv0FlTiuZOcapqetpRwmy9Lefu0pXSG7psS9aMp5xERRP45e0GhUtjF/NHg
nMe7ptjyMdLtfHeZZtBK8MQqLSiRPYYzwZWscrjlTJDga9tLR94EqlR0EYw/tF03ClPy2RR1HsBB
cPMpuUbHXA3SdSRmOztue64SgmvdrPRW1YbSxv+45i5zmLy7isv0tAL9TNShhIX4B34dSs+j5WQg
vXCZJX9DXbfFCkc4eZzwGqDxKg11PyCdVUvW7gsQ0ty0nGLXNH1G+s2/1rJKpXAkHxiErZRAHqsl
teMz53RHwUTznzt5WUVTtJ22t+g6eyh7XLrv/pR7siKInV11wBYULTF/pbektnGNmCFHBIM37ZZY
Am1dIGi5o+WfYX/Z7bnjoHRo5cW9PouNaim9j80I2Hfb4GGTg5VnG4BUbGJWVB4Drb6qn3aadLVn
8/dG7l+w5MCWrfOPLOh+3DB6rwCseCCisP0NLZKSvuu5iwE4saVJrN/2M0iDEiCKYbxson3JAsYF
6DGcai8jIBruiYaRoiLrqKv3J67lQakOEkIr0xsnoF000HzpJ14oULCkUZsRWPSxEK+eJJ8t6GxD
CVFvquLyJFXPD5P9dUMClNODCSAeIcY5iwSFNsKSXj4+lqleI3yf6mG5gExPFSvmtCWBNkxOBkSO
BW/dIxW6sn7LdHMqyrCuKyraW4FW4ZgU1lpEH0kAPaf5vGDM5BOm/UCq/BL6eHg9twVVkgWSJ59e
6gXPuhnqroJD2FEDvWhF9syjLSmg6cZZApHrtf+Dvx/wpB0m0Ug38rGHeCb84Sr4NHTTFmJSHPTC
SpIH3Wt9sNUsL5rKLMfKw7f7P/tu/Y6mNKUNp2J4FjXkaCMbe94k2WzcMbd7Jp2fkTUG8YZIMuve
+LKoJ0H/ATNrR/l3VhW/yAgLqv7Y4QvDUP3Yh6EtmyfcMinUhJUUPsFt4ddqhnA98SSjPyTMsYxw
rFD/DU5lDXUW+yEF6JqvgUmRszrlvBLaD/Ww1MruaJadfXa3Ez4fdpRkgK+x88pHHi+2tQU87NVq
vIYtNa3RommAlaFKnnBYow4v5wTyskevbWqDLv9Ukecx7/HKZeugku6H62oDffIb4M8U3PAg2hV2
FQwHiE7iGYM8he0H6pCdhFdhHla+Bt5QLZWFOuVIFsbX2h+C5a2575B/YX2UHmffDwE4v9HDbcEC
eB327NjERlBT12IMcYiyCC8SBfZgPZa1IHESUCT+0ojSOudsUTc2Wf8KxWCkRGFSjFHB6+LuKtHG
hSQQsdzVq+6ZTZUB6kiIpRm9pc7a1zZXGF/7QnCvvEW0owDVhRg3YwVU2YA5x4/usmzrVIsGEi6H
D2gpZLC60bCzuDEUu3kf2PMqdA1PNNOsWi6M69oQvg1920bM0mFgAUToLuEU2Sl5mt8J9IF3g8+w
s1kM/IdVW60236UIbYb7Pw7apOXg3PZXb/J/iWyPstSovchKiPzkYF4FPDcL34PNWkdkC00NwJQE
jJ22NuNOlfNpja/hmtaOgi7S0XBGpFuwcEmIjtM8s1uFAKl5X3L0pqWWB52iFBocu/+5ejJwP4hz
/KW78aZ2oPhGfagtKW2jeEnzVcy0Fjk2IFdP0imI70H55HOYTTuW+HzgArORzmPwIEogesqYzIKk
lhGnFMysBNn7XxFZ79m3m58h2Z4QkSeFgzjXBUlGxnFLscCeGqk9YI1/IlLXWqXWTycYEDLDwmC6
SU6g/4Rj0LphxPSLWIXtBIcMFRsGcmmmkgTUASVGsexA3V7EPcq2OPhKPPAcXx4JaVrXiPeIzXEZ
TO8lmDnIZ2ZbSsz1JNQ00M0S3Dn/KA3vj3zkM7ZtT8dM6trnB7QXakLcKWROqXa7rCCc4Oi7oCjd
HjQUx5qBIlkJCtwTlXS+KRrEu2X87UGlhRcqtWgetycGIDWgfnMT2l6bTJsPR9jWQyEtvMSCvm/k
0npU/o78XUKRLtZi3o/m5SaL9FyakAcptOjb1Q7/PdzfAe7JfGlwaU+Z9IvTe3jRx95F3JFxYUs8
RSNohcCbKc9h+xyEZB5/Yp9/fxEu/QFIpxRXmb/Jt62K5bhXj6vPWTiz7kBGVAo+TtYZ8XeCWLOa
FPbrstKqSqK0y8gYrBxlJVx4SAWQKna9CE3WdQ1V6YU8EAu8gpX6SSoRqVRiH+Sd8HF1Dpw7AcUC
NCC+nljc/cpY1QSpw3Aczg2tFCerlmmUQnWEmptG+GBdBZ2E9jajhjUeOza0sj1aFBsYT0meJUQr
q0uUCFWbo3xCdH4OsTIbiMx3MrIRbOteK+IyYoWgR+vP4KjAgGy4ZtN4UbZFnZxzX25cAllNZlew
WNYTdhA8bJ4zMSYGxlPvPwR+Yq0GpuQ7WIzjWqH4A0LaZpj75DvRuqIvkcAoHl17rHpnmubiwZ0/
FJ1+9LUgXrhdsKA2SqzaBR0GDc4J/bI1/Q889O7HGHJQ7Zsi9VOcXjwL/E254BlTXtdt8YlFRzhR
7YhuntYqDuAmodtbO+bwSOEOIt1jMhKWnDGLri0KQJGWZr/5cqHceeW49nyWUFmtfjYUlMGcESpB
klx9CkRMcDHfceUQjvVHepkO8YSjshiDuroNj+peXASoBQRqVjUDeZNl2w9hE/h+78pupjYjim89
TNQjf/DHxAoDBvQDLKiEJCKtE6+YMeaSg4dEm1LFwYnwWgvVkBF9DfM0lmeeyPMYKylydxPkn0LA
CD7IKWf10XJ8kI8P8Q8RSxZ0gq0QPGOEPauC3KRqqV148OHR6rjhH7eRqk7aIQ2cApfeykd6qKPz
rfpbL8JISklDsNtlo6tlvhPTqDEJ8FFuGfjC9S07JB2i8+tgvAnOnqMXlwbZpsnrVZrQAVZ35oJp
iIS2E8ckQfalVWKwEciot7TsXjuGejpzDfowN62icvplIhdBLOz+aqK6ytNiroWztqj5UoYumxBG
aorRNiQyxJ2exmm8nAUnLhxgdAXKRlknNjaAFwiGHmfpF/5famtn0GEmyq5aEw+dg6VUzy2+YNuv
7UTX/ZZaHPk6pznsVoYvBwqg0VvLAuzU1Lxywn+YeStRi3v87Fte+FdNJjYD8NPuJP5rXHm20qDM
uuRIifJ0qTX7IRf3OTCzslP2o9IDHbmbR/JcNdE/UG5KZEPLkyJmNSWEY2NTzHFPs8QsPVSEVe0+
uYDwhyUI2l0JF3u4aXSX6i62YJJFbNP5Mda1IVjqikcgPvlyDw5JaNpHovv/ZjJy2h3T0ZrNWavl
RqKN4IrpKGF8gHqBUKn8m+WsBOphHXL3zIOT29eACuPw3g2lj9AId2Lnr3YO1T+dz33N2FwbNMGW
cXjfRKnNHovNckeG4BBLRneosJxyq3RrnGaJLCvkNKybTyzyoPRc7P/g4NOiYpTNAwLhkV47k+KZ
yQBVF8sAzjh0/b2QecMyfmK3Qv3Ilf4LZ9o7I01XsT2FEbGWFznZoP9X2eMaA9lXy/veeytz5f9x
mdzXrPOd5ygUxGdK0Z28Lkmgy5SWwq9EO7kd8WR6iv+DdpuirqW4oY1/Ec/aXtVjuzSF3cx2td2L
e1jusT1fcvTH2EyS8DsMD58lC5sRM50abkjEoEjXN0bCFlMSDRYRMgvj2dhGVjgI+/3J3+yOp1EI
dlzgDwsZHtb2sbKwmWYOjhcVXiPMqLaDS2fPnY3OrRJWIdfuFyqTrJvwqBMbt5BsvpzcRyyDSpR5
r289kf82Sg8Cuq0hm5wUSL+kezZzGLJQNBf+IAQefPiM9n7YIlme1QGfqtwBZpAPiR1pjGoyFSzw
rxBu7rgBf7gPCzrlyCwVI8r/1rPjkpLbI6TUU+vb0+vRgfDD2GwTBW0N+pTVZ8Mot+wNh0amrgJt
QkYogxCXmyW5RQQYBowR/dyPnF+gbP+glQGYSW9UHuokeu+L0ufCvW/mb8t2cTNWy4kZaGn25EXo
7+ucFJx1DRLhEtCpZa2WilP6ixkaedBPG2izpMzwDRDu5BazSuKEXDpzb651j1bYhSCn/FNB3H3v
g5QrcbsCQnikoPnpL6qEXAeIe13kv9JV74hZVcKSgpZtXf6Uloo732avCmZcHZWC4qDrwVWqGICu
278mYB9RTFBjKOkyvNOKPabBOH0J33hbES9F8gf29TBUSrJKXPp52UcW+lazI/ApFmqg/wirFLM1
HTOLIfmyFlzKbcqpZeB2CoqOYMq3ew8KkWhAPIEuQ8hRD9b91U2IjfIT7X2l5u7o6GBAeevYSp+3
jkkVyFKwYwDGTAmxWVDn/ITzd7HDSK+tl/DOjboGbzrLFA2/3x/GrPP9gGcXpmrLNoTbzIh7dc29
g0PBiacKoClPJn73X5rrLxTpkBWOr9oqqUxbNd3hWAUuXriKefZt+mERWZzEgvx1WZqa3Fp0yqjx
tSsqySwbb3VvqkngPgkYzlXjOe5/5NrMBQOUn+CoxZe+NZ1frdqh9seq4YaBRO65bNTI1aGu5ici
/WJfedfeHepKVTEIYrNONIkPUOv1/BHJQmPYSWiIR7LNEjDVzwPbloutA2GpPuZX0MNoVmClHYsx
2E/FuYKwlHuUIrAKiMs14c7UVNQFWdlvJwp+ZsST5EgGt6Uc+NMQhJ+abK4hYzsPtnDdc6Mf+Rp1
CbgjmvkO2vv1DX3ZMuEov29FNX+TqDg3f7iVt4nzty31pjNrswXutNdyog7HuFxcqRgeL5H2t5Jp
N7QlpoisYgf9i8GAnA6QnEMAfKCKPNAneoKPaYDrhc/zIqZO36j6/WaCXovadWrntswCSG++JeT6
a/XaTOJlBleS1yhqwwljfOV+SslbfRRfHkqmCA3jPLPX3dX/h1z5OY3sNNxhbRMd8ha4YSD1+fWR
Y7cVx4eQ3Q5dSvZE9uW3jW3cKhVEnyauCTqGz9f4n96FVBqMq0SRk8YDY7uBQV7jtdBNgWR0KPXh
ygf2mJ0bq9VVaO/S/iAqVD66b/99E7bFIF1ZZKTvcgwwNaqrU9nF2Vuf10l1pReNzClmuwsAJK/T
l18j3njXSc0aMyQx8W6ganM+GBo7PW+9agB3bJ+Wx5/TXESDyply506h4MEN5daWi7g5gUKStRyF
/slHz0u5J7Ue6KXeNmsSZBuyMzmwEII5GiZp5UKN83RC0tN1Y05nhmlaLFQSXRjHmdj/+BYVk5M/
cqdkxM62Tjh61013EZfGJy+p9MrUGUbO+5YgSX6w/E1DeR//zb+MeodRFSID8vlUwwnsAPjDtFKp
qd4LOiSZBT9aTvVokLwojGWbB9mJ7Ctj9EgyUBrR8fDAEob6O1JmrZnmD+HOrP7+dK0UHB9VAgDH
GZGUHk48ebu1JKny0U2qwEEI3emlUxsnxnn5XtNZ7K065KvsTyvqLa4T4qH7ggmwwUJ0jJIZYlGz
IwAvU0sjku79VkHhuuPn2QlYGbvpMWpjIIzPFhZFX7JYmDgmm47VcweV5RUGpeIU8UmiKDLku8j2
JLGRbBorO3zgnSJJP3redRNSHQgmZ5rYrT4yq9y2MFmbvrM5Vzg2TmqvFJd/HlcRoUWaooxQyn0J
6IjqQi+EwrbekRKhJ240sRal+u4yxDUEnkLIcG494p/DrM4bAY8AgvaC9ojTx1zmJAP/mBuUL9yh
Zm4Qkmq3EjUmIdUgzy6X70ps13IZTHPCtU+3NQT4hihy1Xum6hFQS+jpzxbYTct8huccYKl3b0A0
oiJdxsW5LUHooxyJbfoFejK2EC2byOPe8qU2tLGU1houSW4ONHdEelH4n2cxoYQyefdLi9m7+Rt/
0DbR30MwYXcqrsxUVmpCB9FXizB2yChOg+Zz2rAbP59nGyLmX3ANsMRWQoumtLjJxt0Z32ubk24B
yBTldz7lwEQ70kZPqNsl6lsjFBpyIcnyTjGSVzDlLtFEy0Fd4q08doiNJOa9/eYh34XCdntrU5wr
XrDn7g+dxF3OP6mkfV8ptJ3OnzQOJS43uUqo3iClK/SAnHgEQ14R3lJm86+ly0zfjsJm7CdbUwwA
gXDkF74QMob5eG6gvPQxKkShfxgBum2FtrGaKyaSxUzpktgJyfGRFvDV4YvptOk0sk7xCWwc/1Ou
TPMQTkg5Bxk96FkOfhWNt+jQX4B63kI/MQR5NKilyubaaHrTyJhsoW9yiKwyFA5j0FItqqFx8uB+
lz6HK1/ZVLn50YkRNfggf0oyA/uV4ZWhy0KAlWK4ZF5uiyp+Mv7x/xCknkbW5F6mbvUEkOh5CU3y
ZDlkN4tchu62PTjuoGj/PpetcSPwVAdsc6nGgtt/opmZpXfNa7F4xMOGHRrRtmY5AKNYPX1VNtk3
remvndMYzVlz4l4OhcI89bQqhacYSKQSfXvXouOkXwXwsoFN2RTO1dNAambl+SqSH5OjWLcR1jSK
QWccCXsoQtYAsNgwNTOkLaKZZiKHyX8YDhZUuGowQPt3TPk2iOiV40ES9hnOC18ppQwpzDIF/1Ks
NishBRNpe6/wD8SCtPKZpeFeH9Pae3FWSvv/XMRQvkp9Ujqd3/u/NoLQu1LEpuVbr7x/FKEg9BOy
SZdzrz+kq2pK0Nvl2izz7g3Q+DWyIX7K9BiaA913+foC+zWtp5merw2EP0hQts5FC9l6b5Mbd6qq
IjiyhqdkiWqqBJtIuvp9ooXrnQGdYcunMJBTbEj9vHd72IZbeMAaoI8eu65gLKCfEQUZyi4cDKiv
P1MuyiUV60vmoMo6JIbPxbk3EEcZkyFZDi8OUHvKFGOd7P8q4zOux98TQLArKeNXDtsd2+nP+BIm
4Mvs0lHklGRLRyVsXllLjPulPLUi6HbyGbFKntAZO1HBTK9lQ9meaqdO9RwtbxTiH/sYO0wRcQN3
4mjR8ZxeEM87Omk1axyzrOFhzwqRAUXqnmOG31uA1Y2WsNOu7vZaMfxGQYRXvl7CEwLjGpMFOwtc
tB0cQm/44eVvItJm35Ij8MgPCSmtnJuwxyNcB4D3uFZOyqGHI8P2BJuQFqb2IJZ2HyuwH0R4M2ZQ
3ohbt3bd50J6AwQF4s2m849+dCmBclG7NtbAiYFVdFF+kxr5O9rMAJ6AqiKtAu+SIeYpzl6f48jB
Z8mrKwgny3w7UCYLX33Lh3cxkxHPve/fkS9Q7NRUpHAq7c2wHsYepwDnq2BmFJbKUZ+QzJYkUaki
7Y9R4ykEvuMp3OusP7bwvvuPChk2lsnME8qHB+cApB28UDBMGJSRF8xJ+AhkKsZg0jp4jPS01Z8A
qEk5+2JnjT9+X5DzpXsAIJw9JyTCxOWFof2oWwV9tEa1QVZunX0SW5CcMftCx7elmphJxmcnC2G6
+vXYZm52wV/eAr9Ueoac1//xE1HQ+f2jPxO7uxLNObhlBRCDOmh66xTsJVmkT5XvVFchif+u7lhD
kvQ8KyzbOyTPeUvOp3iHZAQD+3QkrXtpMGb0IjRiLc1U8hb5mwJQ/q+ATkVoqRWBuGs6cj28f5mC
edQYH4P7D5jdqIiHdpfy+b5XrrO3msAOJjkFyEEkxDhLVJLy/dnPg3/RiQ4K4DcvD0aPujWbAbzZ
5Yq6KPSz204NhSwiKRpFMAk9I6N7M6+ABoDnPIOYEZZF3fvwAXlnk5o5qQgxolUTPiB6IMMlPFo1
LooWuWOK79+KG+gzCMzOa5kkwksShbJHXPBOyHENjCC+zPh4Dwx/dZNWiGgODkK/0ydkPlEvsD4O
5BfcXDuvy1bZZ93o22t/s/qjeSNyf91kxw/Q0CRXhl4iiyIca+jKdbidrd0TAigUVpG2wdwUQCwS
5O0iLpFz6y6L6Vvu3N4pQAp58EZy6tSaugh0xbQSVTKRkZ98ou3DdUOXe9g6tid+GU4EiBW7n8b5
CnWlTwOBzad85e8Xd8KDzy/7SYfYtrrOs64i7KX6sv0INtEQBcYI1Y3pdsb+6t+NJSHjPK7RbRr2
1U6/kxysJrjCl0g6sTPWnbCy1oCB7u4wi0fAH7CAXU6ZoZ2eyocg5TtmZKZnTUx5gUZwOZFpXgqz
R6H/ogmjZDDKADlUK5zFhGen0oxGRIlJmw7HxDZ2nSiM27ZXy/ZcwXuKmqgXdM3pMxEyeEc3Vo6U
aAXujNfGdK/ouf2syjvn2jls4jtBlxuwMrMVUkPZU2ddzW5kHoTVpSXMHy2jai/XjOive2uRgbzo
BNmJHyys3omE5BR2jx6s7FM3PL9Oi1qFqW9hlSwnW7xmBTpju1kR63vvhYMLTgFTQPJ2UCteTYnR
rdN9TtgVpqyod4RsE1wtfO5kOwhgJIq6kmGAuuddq/PLlTiGXSYLAFgg12PtC6EtiHD5yIlRhwIs
5J/w9Ei6IfS+oDqceETq5AKigYf0J6IN4dOt+irIRbbL/VNUmESYO7ZZShpjgzgLbv12XnvwQHrf
M/HAbAt/I/Mka3J37ydqJ0NOYRtEWVH3O2WMDPPoEBEaIVonzwQWYH5LD78Cmij3vnpmg0fbk5Vd
gUYF8IvgscjgyhStPa6F5NQNrnv77iCOvqgNpDiGovYmKQg3aKJGr9oj8lfTtsRHU5FKXwjmks7b
255wYpzTlR37vTBSgyqmBxYabwLNz/XzaKODO/CeQiHO/CkOWmYh+e6Ilx+y0lzhtF7quC2+NQgD
EhZBGR+/FB8bONutQ3uj4TOIJA9Mxn058MKcUbknVxGpTAh2lnq5OoeOR1gkhWwDjoQXzTpRZtIb
2taOCaEfr/luxyh/uil4Rl5+cHVRiNYPslu8MdIG4BSIYFYqcdEbhRfMk9k3ufMEUMrXWYDv2mjK
rmHWCcRlbnDnNOJTVhJOTpXhFLmDDDaa2zNxOj9urpgdTshOPN5txqxJFwHz48WfSwVJcZID5cr3
5LuCT+8ZnsfUDcaw+7FDWuGpxgkDiWAmn64o7f2XS+C9/g9fGkt5AbdjsLX1dUmUOZTiTbntDxuS
pkCGaSjHZp6QzmE/rmJWN20h/GevBrGLFpsH9hLDuS1ZLXLMS496w8wOBJSO/uno6nhORXvSRp4a
zbOQV+zmTLd2HSmJgHwdMNasujgjU+WRJpC6ofLLUUizbElnscvjPCKsmmyVprj43yHNCPtC5wwh
4I+XoOtdFtOO/fmuzj4EqDcMYT7RT9WPgy7APMaRkSggmbVbqVj8hD2D7vmFLcp3PgkvAdx0MAbx
hpuKK8+u32smrrwSB0NePz7GEaFcR3LIeTB8uqI4e5o+ucH2xbQf3Olku37TxI2lEKtcr7yEVElS
CBd3EzDTdFQMQ63kkDCF4Clax/qjOqTLhFQbLBDXb/BX4stbmUrsKHfHDZwSD8uWtvbidu6IjLU4
FIPxq8ZkIwdQUzbKFFrNBS+1XHzuQaaAKbuqNnt92+6rvRANIGuH4h4fCC3RZ3KeCWuwmW9kEwpV
Y1XUkf5O/fc9BhGMe60I6d1HIQO5+stmaJMwmSLPT69yOK88XKf7RDMKIiTOdC6U+JxtqjGcsDq2
Z3p0uyVaf2TD+wrUAijtyCikf0HZALbUAsqkDCTlqzbldDoepoHPQAW4A8BpbNA7o/WbomutwW34
7hLVJcSnETrAwP2fSGIpvvItroRG3eXn+bSAbtabNTggdNNFQ59LbkNYR4xucGtdol/z+1s9EFR1
7cuJpoMbbSB8OJWQ5g/9gessQNdwknyuYQq5VqlmuwUuQ4koNgULIjrLV4PfIARUwRj6Q2Y992Ii
7iUr+mjVNdNPJ65p94Fc/ARq+7DTfCx0f0yGJ+4ynZjGgbWLpu+nfG+fagobMAY2KZSGwbp7iVFh
Ta5Ec42on7Z4KrKLM0cHj4IvlUq1EfTwA3w/7JHR79yVFH8NOcvTO/i+JSCCPLGE7EDl5YaRo/ld
p3Q9te6wQouthp+RYg7JpFTXHnrhOSl2vvPOD3XzRM6Ao7vDuPxsE6W+FDwl7WwGluwii188jhgM
2z14s38PA6ztNobSExbrVdeaM/jvOnIgPqgVEHnemS8trtCVoJ8RNrGmQUhVlpcCprq6EGV3273M
Z8sAVQR3l2U3WEnylzVmnl4AHSf4XtAQKCpmeJWPpn80FZ6LFYYRAqOed0xlgbyGHZmqV0oLa+4z
0m+zmjxGAem2gzB4gsz5seOh2BhiI4/Rwsj7cvLGPZd9tFxh5g6TXFF5xoudQEdwmpDP9qXshlyT
cVpzCvYDwWUbjRW8KXeO2iwVqZWX+qj8EoiCGMm7kma6n4ZnpubnFCkpX5+kZjvnhtrfA5aX+1qq
9rngQXlM4J9SwdhrVNa3WyaFYPl5vlp8WBqOA6XFdtW2m6rkxK5Gy/60GP6DHd+ayZ8MZElkt9Vj
N1npF7zVC2nBx2NflOervlKweZcwrZYPdCtJp4S+gGRYueqlF6VcK1dAeFZiUwW8/qQFyueXrEzp
MDFYQmY5ysSJWFg9Kl81G5LrJh4uUFj1l0L4vPaUi8SQ2EbJhKIuvpkjI03IVT+OPMCcyzwle64r
2jVHY3P6VxCx8GFlAylODt0a5dF3DWYUyPAqU9gntll3hRqRjGN4LSYiIvyUJ/Dvu8tDDfTQRF1X
fVsp2B/uxcK4NNaUV+oCx9LpA1HQsGuAjGw4XHF+Uyxfsj4oyUwQSWEQr6kU32rwNLTxkP7VseiS
MOQMY9gIxNcfKd1X+taCmnSEdrPDcqRuCvGEw5/CguioXzCKQkn6umh8+79iMhtnmtz5xsx6vA49
iMd4xTQTb4Ia7fjAUztuSm5lcG3hC3sypi33SVRXYMbLQXUIPQ8gCnTVCtWY8NtpV4mizkWbuHJn
h1YYc9uuSzu+Wx/MY2NY44qeajTQ943uLJAb7NOTx8fXtO91YX7xjvuIcFR2J0mvjW7a+md3uU3z
KiwvkK0OUgxgYzpBgFlxphegaXx94fRPzElzKyFB+ikNaZIiK3dVPv7wewEMhuayxLlDpucBWce8
vBZk6NHL4nQomC6hMpXB+zNwku5onLF0feEdPxvwk+UiAr8Uq0YNELv1sI44vxG/XGzDOsIePFTQ
ROIbBXrEzUoRRqsaW0kbUj4ekE8K29XWx6VRZDTOjO2TvLPU2QtvGWvfW4rY/jhvrgaAontldJ6m
xbK04Z+IqKAZrgYjPRzwEserdBpwgmo/SwRzI0PtFbOJ2Ty8RdJupeiIUh4WZ/ceo2Cl6znhY3VG
lO42t2wwJq1R8eXjswhPFjWwn+290M6HAQX2CI/Sr61KM4bSsweXlG1fLf45aPTm14ZoJT2s+9AF
JtDNmxmrB3iSAMuGr/5btErusAzeNyihdy24FGfUHUwFMcRMXeSTAASnt+9gaW+Wx2BGh7edbpta
2VkY5S8TXcU+sW+/a/6IDrkpqqv+jKOVhakdSoU30t3PyACdLcYVCpnLOuM4YlxtoOf/23igFDTB
XjtZxkufKtQ5JU/OaVRGY9263uSgRGGVPM/gi9WYDRMIGNBlgzKvrxQK0x+PRfxAdTPLnkJL5g+T
PlJVc/iZW4HdBieYWYl/TUOmp5rjRKrDE0tlo7vK3+pvUzItKffCWowsPAaTv0snyUh5O2Y85hvN
/WwNp7u1uOuwVvVdCp1Z9be1APtZq0yMoczTccdDDkXIrkf2qNEOaR+2XY345GZsNXBPu21iynv5
/6vHIpaOroYr2TUPTGT7Nei1oXmfIny1+2yblqdznEJVPk7lpxnuxo6M6GoZnRUvvF+VNqJltYVc
Iuknj99jo5wiwCb6k7H0EJibU0PYtnOxEVW3x4obz7zJbEs2HCTyi1OpdOus2aC5PH5YFG3gqraF
T/r/hYkpdqRu6jZgpKEHtLxdoAT9qnr5Xdm9KeLL9DCT00A3lskueB+8iNhIYNANmbl7UL3vGnZS
m1rXmvCSie7wtS3L9lMoNyFflBDwHAnbWjLdq6OAaApCpGUnuS6Gi+8uBwe+4JygyrSm69hCWj9F
FC/bWTAWAYQ4jdsTaq4AxNS5BvNpXYLMv5PDY4EG2fMjOUgq3kETDSbTvrcehUOJqw8Mwgs/OHI/
rApsA2F8W/Vw4WbrbP9/+s1uT7QgkZvSepelsXCDWv5cxnD7mzu6Hqv6D51AnnYORAy2t8bQpvlx
S91XQ4WmmshkkChet9efJeUarINaMTaTBFPwFdUtglLSuUrq3DtSXSnO4DsEPsd7PJNiFUCI4cbT
9Duy3KeWPzrG3kLL9J3PAWcb/19CQCF7GGVJR3KrWSR1C7Lig9cfuCBHy+EY8PVc6VHyBlh8kipn
LKytURdLaBM51w6D+av5csvAugumtdZYrEPPRcYCYuzP/z0nXqfQ80OH4pw8O8xnV8QrbwG9vpQf
xduSGFMAc3whMwsDJoD3Qah55SHg5JnxKBsG4KeQ0Ip+SLAieG3O0o3C4cufTmOGGMBAMIgRlLtm
Tylw60MW6Vyk8Uo8LOj7UsYbj59qke/lzM5kBHcLr/x6ONkUWpFkqkG+A5idQ+I6BfRbJE0P4M2D
culsOsrfxtdOyf3eiZHFPSGi2ptOH8dBdHxxjgFMjm37c7bIF6IqHN55vTqgTbLjRy+Bt/MY4KDR
HMdDjLjJL2Egumh/+nolUmpaPDgmAj2KC/ewRJ/6c9chR9aBROsnYU7X2BTxLcEZTCBPaSm6uBdL
JFuktG/IPJwSGnUUzNMBgDFMkR1rtiAwx5cGVrMzipCYvDSrws6P9cFwo87teyBp/1jzx07lC1w2
EYA1FAd9EXAaHewu119PAsCYwnWNmFveh+CXGAqhinKhuhshATvjVZyqIRVPawc7v1zGOGpnp4a1
iCTzMXlei5HN8YGvmotLhGUgzcyuFRcHNPv7Z6OfKV6/Oym0kQQ0ZPo6Q0pqHI0A81+GBsfyd9A6
Ebrb8hFevxC1O6AMinTzum+PBtKnDbWL/4v6rd+W0Kar571/aGaHz4eE/tcYkOPRKRNr10/SpcFq
cQTUPv7wYzyksEX5IUaGgOVelR+e8ixsHcnEop7JnHtTTdyae02RDqXIkJ5lcgwcsoXD7GVh1T2m
XTbO7niPXB82mtrMAhQRCXUaL8AHCd79lUto0+P8CEPHJJp1xDwtrBwkHjEm4dWlNdDi4JL78JEP
4X/Wg+/IDRFAv+txhUiBO+1mmHAwV/WIaWdxf1/5yB+s1sSwnnbbmoOeHSOxCyarhtc/WNxzHQns
tvPuT5ZsxW2Wc/stsO74J89Rc6DwyGUKUoQNwY2MDIq1zJYTh0MbIeQigwLETA2EYSvuzvhPhfNz
ukbfrHnXeVYhD20IGXpbZws57SzfGc6g/awWsFceEO9U139uyRLPWvzjwsOQuOEogL+sABcCu5+h
hfkLFpy7etR9a6i8kPDGrm6q+VFTHGuzJPiXByW1qcNa1AkadE0M44JUE04n7vQxJADLP1/63CpW
pthg7bD+DNovgrpBJV8Yt5rPf8Hv0U8gDcuefDNa+ERjyxAUi2z6Cg7g6HyDCptrJe8p524T+v5s
PTI7CmS6AsVsw72rgbrdhf2H4xjE3nWOSrm3NtBGR7Dq9ZZQpz1O6xj56D1f6jROONvKLySEU79h
TePBxlo+yTXTRSYg5y2wlvI8m6+WaeaKYdR3fatn5lxsbXN/gn4giUsAur3Xkm84F3pcuGNVlwlC
cPnKpbp8z92bVowMkWpvHVI4HjdGjWqllzDrZ3zygYaJkIH8n77DvPZTKP7twCt5oW1CS1LEcrbU
zBFI3VsKfPSP4Ld8MVHs5vh+msr1/YLPHeH6vmYFgNsn6JvliYYki/OoNdl4bQ0bM/yDJEnYLFQN
9Dei5zGfCVoAhqudwGyyGbHG12wBrz461x8spY7Ihfmiv8CBY+PSYDZt+Uy9MfCJznW+quUASa+O
f3jtxqcFTfLCtOmsWIkNOEe7Mf6HYpxVi77h8sh66RDINpql7aUL1xLRhH404cTNPLMXzPZmeG8W
aqgdRxbiq8GovcPxRbUmXI0e9ABlWPbMl6giozh83ZsOq1h/nx/L1IiOm+/XI/O9Fh2re3e1CBlv
JWk9jIh5a6dSXrQ//SVtP8fZS6yMbyz/4uXDUPfpZHxZEBh1qyGZtJE1DVneRiARmslxrQ3JZLFj
swS07V7BF12GIBk8++X3rrZgM+NGXdQ6sOlH+aUKRrbI9KCXU8x8sdcL292dlw6EdB55onP1Xvst
eMMOM7ni/d/qeccE7M4a8QALmrAOWSVdv4UTxcDiB4v8fP11czog+M+vPZH5rMoFSOmfxdwUqXNh
rZeEnpQW7z9gVhDxXywM7rsEeRTIGhEcKuSSyLCyAPsRz01CLoHVTuJcbWFv1m76L9840nJ8QDXO
XzIeH2viAJAaeDbOZnEywW+po0ucZUbMWfffg55fDotHLdZEA2oSHBKfhOojLOm6CjlA6tF/wYgc
k8xJnZTI87PYco+RAMsMthD/kAYoBBsf3QJqK5zx9sjOyHNx0djYE+naNDIATlMiI2ZH7sy/3Axa
zjFRqvHiyKjZWeYudVhyOZno/wxyBEPnzZxvYDsSH6sSLvN5kCuujAT6fJFfwWOMdDTbezOJC2tV
UD1+L4DLV1jif8mJBwnst6Y4ljQDyTugA7c7Fzz79QNFHLdQUcpFU50LcmRIlTUSPBGdagKj26hk
kGm9b9MHyPSFjqm8Pj6rHKepkQzh6B4tjPYXLMlu4tBltDokqnGa1iQX9gowwS+H8o25ach8rpNQ
3Zs03kVooYJyYQNEQWwNKcc/IcP9UrXWHaur51vIHFhQ4x76LwqmoLXmxptXt2ZeZZdAM/TiHHwb
fPQyO0oC/4VZ0AObtK8pn0V/eK4FK16fnaLR7FGgXVQ5/le9fK6JXqdXk7XanlHln9/BBc9jvz0m
Ct29+AQEHI46xSUMkoHZQyeDRqawUS7JzPB+BTdkThsFUowpfqnodFwjS/jnGAs2sQqnBbQ/3jDt
DiHzvBejuEIYhQCXv94dG5q1+q2aaxdBsbrQEy92GgduSMnXghWOidzYeetVg8ERinYXPJm4mcQp
RoZvmgb9ZozPYYTYF9ADerP7elQ0JotZmSizRfWBzn0Hi6K4ywxEJ9KBaLpxRwMMXADCmaFrpGBt
5WOZyAn/1uUdnr2d46mkSG147Y9htprnUVcmotE/+XzUM1ttyWi6J4GsJ5g616UjkR/JI/x2UosO
wCW4LtfNoIavhTHWLgM3SqL11XqkMDbgAcKg6LRHQKd5nq44mKe9CXFIk4QdNRNQ3uORmjt69hsq
u8vgmw+HQ/a4dZtDugjhlSv2Se5QqD8Ymid/9mlM35fD+iexDtHvlqNWAJLXozvCSMMZMbJLs0dh
JUTjSZtFWdPiagjyeSf5o1urKb3W6uyNAXeP2CgU5v/FHq6IBQbJQoKhgqVjujVFHnr+ZrP0CeXB
VQeDIu+TauZZXq6QfyG3mCJ7Njcue9JhN2ew6siMgv6vSgXVPdQ/R0A1JV9hWf/GuYdNgkqfM6Pk
6ke7lEvxLtL/ks35UiccbFt5dGbpNq1ah6McGODHsS7aMwndsx51WdYHG7xBDmtCxBrV1YaMkwLO
n+NH3n7OQuMCHELzcoE6W8yj2usk6Z7yj+bP4p/W+qYvyJCuhUPPFnAF2j5/7U0AJ/Qi0CtIazzP
vxIke5hjGynW3QlftU6SPloqA6eMbhXHltoiM3/91JJz1YKdtfHM7j8IKLVFt8B5QLHYpG92BxFX
xplVsCKzttjYOCwD37zhncnT4MtRF0ZbbiQPUkG2/ikPsgRbiqgYlQpTXv6480oOUeQNdqmyWxUW
1xk7D5G03UUD9grPKOZS4pWYpKFbPzidAl1BjwnfCNQESHMoiunhIHH5D7KexxkrI71AO5GyFDUO
ucpdPrXw9pLxT1Ixd0FfUC9SBasprypsNdxgXrXw+qwPzCQh/9gDmEMxJS1+K1oq5xdSrSTzGaGv
nrJGV4AHa6d0JtHd2UFSJOidlKpLohOq91xLfE8JDE5OJm5Cb4WAgoHd9dclQV149R8JVtssURsM
EIiHGmZFIEgPYWtGB1IQjv97OFPxHTxqtDIV027Jpb1oXEqwNz2GKtYiuj7NCNIi3cARm8JtqZFy
ZhF7mKu4CEJtFKVB5M3ZPhuHyZ+9zyxFaehIGhm/QQYijtkAI6L7nfUByISt3Xyx+GXCtuxQG0sz
Zbd+GFoEkKt4kQeAKyFW9UWcz/a03tKCgm61G7+LXVfB1iKyppqv1O1Zxfmt8y5xUZSHHQK+gNCj
tFnBlHbfBZW8Aa95fdQ8MMWfB4QoDuUCTnWRAJpGL1GNUiOybNbkdL94k0B6+vqbT6yv72RqtTMY
9h1He6Hx0Uw2B3fQA9sfI0NmEINqXgoIpclGWfCoGUP0OACDq3psaH0ENkWE9na9Fyj95ud8TB2I
mkPhfgH/HcxiF8FtUN/dla2x4jhGXl0xbwvJUE0wKa2VrQt1/XhGzc+Dl0BoOOjeC+noRtLvVaaP
3HSphUx304+qAhfq88InDnjW+f38WIt8G6DuSfDko9lHa5J+xsRruXWGzcZjaqOZs8TWHBoqhQwa
eAaiF/5JRkvwu7FU5pp5QpxAPK3ESypJbHXMj5OLT85a+4+6Y5lJ/6WWW682YUhcqACuJKkKeJOt
V9VKjOfr/4Fve9JmolK+MPyoID69kM2CBUjyJqZhl1Rl4+0oJc042YpdgR8FQjgpR+A27r3NNG6r
3LAYGZzaz50UOZtdEk7m9nRQF6zyP90qj1av8OzkbPe2hs7RpaE225nhS91GbKX04Onj6AOoJ+bd
aUXg1+ril6O42swsn7fq0/BtkvsRAvNdY6q6/9vRc2k2zW+pzhqkQ9AulB6YdPQ1Jx796yy1mJ7G
qHX8Yra0+OdBguc7yxV0z5Nhp+hsAiNzOwnz+GeHVT6VDi/hMzBPb7MCBaKz+Aay2nwFtOQ4fkwq
++zjU7LgbIrOv5xQkD9yaALQOeaZsQV5gK+OwKTaI6b4yyXuEB6em3ZsGJ2s+9sp89Ivked7wrtk
J4GuwYNRrNyvCtaAdKN2jW/ruVXWTViOmsqNkLPNX0MOgd37QoQvMXRhpvjgTOKRVJ93zGgEfLzO
QKw5aoEctsqOw3jJbGKAJI68faUckuFtnL4=
`protect end_protected

