

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bdlZLEAewQqpv1o7OoBr4R377V8Hk5Fd8+q/Az6G9nxroFaOnD3V9+lWQZaiTQ+UR8tYlBixiDT3
2rrbvlUYqg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PNj5XhRRPylbuLUnq16m36512+Iu+tuxUNOB5vui/U9Vyxliy5LDYUjGyTrkosJ5RLmSfgYfmdaq
x3GXyG6MVOiZo15XiDmGz5Xa3WMM3TuUhfpzNItvR+cjVJcfSX1Vpo9/m4Gf2HbgWDY8/uge9Yz+
pdDWTg9IqOS1f9m0bhc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tfy6e9ewB1av8IAVBQg5F0wJVpezM47U5T38niEmKqoHE2EAQIsVtLXdGuC0EVCv8iR27vcg17Oa
mBfBXWB60tzPu8Q6DSJi1RmV8OgW+NgUvCiTMpLKqqsw6FnhMEK3lQVXfOtnfyh9msybPw9byzXC
dambJMmCpKtH2TBazWP4yb5ww1Nsz/1jL5i1zPiiJqwiUek+yJBHinlLsKOdmxiEOjEIxiuXMNyg
LMJzb839xkVhlMYTWXZYlSQVwwm/sLGnZ2Znntlf9sYBoE6D2vYri/PUGcfI5TqvvhrwG3MMHoTN
rPYZvU5TTqkZ0UHzprP9ZbAAvBMMlhHGjyKLgw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
enscaK3Um9KpWwQm1hA2XwO16XJLOAeYZ3URNnasJSAORmdXiuv1QgNvxstTqRmJdf6aiVcX+SBW
QAS4XOQmaHblVVCTrTFxq+i8/M/uWIiPlKdwfgcbq6W9GDVZEH2g71B4sNE7sbY88daOW+dsFMn8
evKdCCrOhrfApxD2w7E=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qn8TdDpu0TmAhfXr6OjdWoz6rfyBW7fFZKyqPOjjqWteCvm3OM0JlharuS1oWtO6vCpto2FAzG/S
BlRFnD+qM3W558gotDG5xKLXH54U8vJ9P7HSKDrDRZfcvgzYnDlLOZYqIhF3QcOp7QlIfdgIFJFF
P1RDJ8d43uSYKR66QV0gPXuT19+tneyhi0YpcaupqD9/Z/vQdGHiorXfqzI+zmAX5/7dF89mvr3v
Pvp32AibqOZJekU7QCnp4VkIAFQi2sNR2R1SirejbeSwa+gfCdYZC/MT0OFTfQjM0uxBSK/I4IyT
gWZgfuPijqASxDrsrURmKezc4hgCDujIExBWaQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21952)
`protect data_block
98IHP4Hq9SjMPq2iRZDZPabLOQb6pnFxBDTvYL3JCgNI3KlvS7y45uM6/7HInI/83ihOQoEfLBrB
lcZrHbyZ41CdelT+edszSUKRpkzbP+OgnZHsnvbFtwpVORJ/r+zoWVfbdq5jCKPd7UVlIU8vcL7C
lJwmjNqPuN/ZWBwmBCyinHtieaMugz8XZya8LvOBkMvhbgfNOeo4vlp+l4PkVJbWeUC0XxyNjgUr
/HAm0WAySgAshfhqti07sW+ptYcNQxoDWActNqEVnw2I0tf3d/6z0a/YfKTeARQJfG1tkU66wBs7
KALkXgR8/kYtNH0XPrtOgLmdRWulRUTtWQbuZvWoaqn+G8ZUUmkE9a7d5M0ZlTBIXQ6CNUTVFwzB
ODL9XN5JOSlcw75vFQYycfXuG3jJf/RAOfCorfQMfUxrD2zNdQ9dZShPu9fZA7hd4CDJVJTP3X+7
ZGuP6RzcdvEAsdgeAbYsp8d50q1piBhMNv9M8Tl2IMlZmJ5XBoJiz43RA35IvmoJJqDZ/lp7xr/y
iDqamZ3iKqMAA6bd9wn1AnEIWAlsl9gVfTMCrm9GtNnVc3Z9pSnIs0/Z0x6GdsyIKSIZ+dnNNJ2i
CmXK79WeMkN1bv5ETt2BQzrFj39CtAxPAIIiCbDzLoDyg58vlgn9p/UEAFGKZlhIr5OBefbZmDI1
TPXpeKwrxuebhEpZ1uVWDWz6vSeb41DGEKbrHwTxyaZ8LEsTn4sQAw/qlmaQP8G8Lx6s+LLk6rZy
dQ8YEr6f7yKbmxnWRWyy7jElR8Ns5ku6ptbYVuLeSPRPLMwQgsmaaLPM/4iG7hgqFLaqcZBI9S2J
WfJ7pTtGbuEIGVZqAUpaepgYq9vFezYZtxd/h5Fg/QwHf3oztV8/JxIqX48XcuPPBgwAct+7WPGQ
Wloik0x7/XHyO1t2UpLXwdqtZVk+5+006CYFrUgV6Uiqbeh1LGii4rKs/yeaoVBnjrOj/QBcD1zg
e1ZCz9D2ey9Q+nfVoJw1//o2ZeYq1Z3TmMUDk1iP6RaSIfqoHhJsAwufWD4krFCeFLrmEQ1zw+Dp
w7RiqOgB1rR7jQElt/ExOaotsMJjsJ6yu/LisKSKVNI960X8LY2MWgIKUItw0PwsGcj6Sx5jFnSq
YA9MD41SN5aLC88ZUy9DgejIMh2p/mp+t/zy61eESrM7bqaAIqeYmDZP3y64dEWXyW9uWWWfcwkb
Rfm622psAJavbkitN1scv7GB+RAdJV2i9Ek2rTjnUzu7tUrpo4PncCH9d3YN5XdqmLi1+YUxdc8w
LnQdDoyWY8PLJ01ulpbAPOCaqvVjlbr725V3X59zM11oKd9m4X5DRuSfVu9H9GBSqPSmP/cs8TCD
jTpVCiaco9Jvg9qDFE5cB5dbzI0i2LuQ2dcXeFoi0PHUUTWU+svw/oABsuSvS5O10+ZnEEWO0paN
51HPfwIglMzQrvRv29Kzy0JidIGFNJeuYwvH5VXD84niQMejwa+u1QWvMnAlq4AoBJB/jHf4Gk53
guytUOKZZCLpcNFjuYK62v3j2/BWEkMLJH/QhSOISzN/Nlm1IrMtem5mmB8QKJdQea+uWJl7rUST
wn2UHSxztYjoHQyE7/rUS2Ll/Jk+IJY7tk4dLD5qLFZTujGGaPOob7bu08oEKf9DJVAgcFy51af9
wUUqqaXBobRomZMICnZOEYLajYLssQSmLWNicNJZxFwIaTAIKnsMuifmKujfcWjaIUSaEUVtU9OI
Ff2cd4bceZlg0Yk64c8rvGZ21pKo+xaRb656UbQO7foNDnNM+Ba5UmZh72sXKXSwK5qDG7EijEHD
wjzlSNpr5qhtou20QujCAU79ooZzEA3hr/mOJMkfayqyAw9FGzXNXjYeL45TnWsQXoo9obGrlMud
zSRNMqiFAeb3RTzyKag1tpapZRE+nRjdVUcZVqImOsscNVM7UemoBV01c3l0aCulgjxRS3sZBWlf
9jzxm7QtNP3BDSi4XFd4kU+J3XnqfHj49QkKiy5I40Ah3NREOFwZYRyBnCevaMk8pH/LolzpDguR
zov0AdNbMVRUerGhK6CVUYE1WJOzerjvPr7YUpnZDndboLm1LO3e0nbQhFhRQkmp14vDhwBhgFyz
1Mm/nbq086BQhQmLt8rURQAZbTxZzpPw6nQ2Wojgdfc1LeLHEB/fMm5FzaHrkII5xR81IYW0xt4A
EBIwHFr9bhCS5JAChQIlwGcdyQM1hw2s66g7X+HtZ65Enqtefr2qfW0702AJcq83sOWejHZnHpPA
wsUEOjhdzCUf//8NHBc8GvvyLzAkAf1YfWfAcUPaxuQZyVlP3Zz2My3u7Gg6IPnhxorFK4BK8Zvj
gEkGZDYPRRRr5suUYUfdZ4QFUFOX0nOetSRtJucOQG82MIO8I+XYBsPXOiH6iaL4JAWvtn6TZOf/
ffpIoO0e3+FjTEWJxjRnAngK1Z3UwCig+YSFqjlcOpGe3JD9bCK6GgytLlWXBKDh5f3/B4BunzxY
J7f8EnOBCBHseuL7K3FASQYhG2s+CzLJtnHcTano3yCdrg5BPMDznFA/IgZFKhr9MEYjXIQ0+Nn6
QZVIudugYWJ0uE9tzSbHcllN66u+eRQxA/Wb163VRpU762SVpFAEokIVyMOsPD3biVo0pmRiHVGe
DeyjOX9juHQXaorH/J+V1ZVNXip2cwpFtPXmWt+ZCmEDifycQe8Sk16/vZH1CS76X2IU+owxYRKs
MGah4Edi4RHNN6wRjt0drt43SQFiJDoKoGBwBJ1Xyb1i/3ji2XHINvkU4cHhDXOmWi4LCYdBkJ7L
ZmdCQkrXMa5i/TgzYLx5geqkYmwLkK691I1qDU4vtMSbtUYmPa2IQFYTA5zTyNryGhKzi4bVdC+A
C5yB9dEwHq8xM7cyPrYW0+Q+eGfh2xUuULwpEa1sBJPz7lKUOSw2RHyVNNaBQgoVcUBdQRsG2Ya5
PASKvpxeny2+Tff86mcnHnuBgWwF8YTYbwNuVkVmZlSdo76SIZVoRY+VAveynLo0TK7afsp956Wn
Op0PsKKmyfVy+vstVocKEMpLldUDnjSFkzN/euzIYamD3qVJuQVOMqfXzvg0oWhwoDv8h6ZjXPMh
VvHHMsA8wJ0tgY5MeJSNUUjX5X3WVHmx4NYwaDpZ+3X+C0McQakB8uohvyZ1L1Wes6g83ewUDb9+
cxfz1pP8SX6Jry/0cL5yIo+RKVyDL46Hnmicu5nq05nSH8R+sRvpOJLoe5i9cWpHvtJwk1S3yiok
tJROmdrH56acQoVb8L3F9oNuBFQcOIsoStrSvGCe4BFJ+yIilRa5gcnJL8oqY44+mYNqcKhpFubo
ki9mRLmMSQp36Tq/CYCaMODan4s2KiwFdKwg4KRBD8iiFn5Jl3U+ShvLMhmsY6RKP5PA9SpHIxYy
BANvcgGa6a1CQhsbWsTC6BoKX1HGj8ke5oZJu3Svrdk3uYPCOdem+1bC8Um/oZWCBMS2BHxIp9xu
oV1QUgq0MfR4grJrvB54Wh5mQlNw4uXDz0mYa3Ao7RhwR7pjk7OgnqPWIEr42qpGUlFJmyQmf/Aq
mTBJ2FRq9NYEuzUfmLxz7yK+GX1cpy7VRUYDGo8CciekZAp5tEsj6j+u5p2pmYXcTom0/kV43CFr
vXIOgqeLMOkFlKV3Mc24ZP087QrlWzi8Dv7OLd+mgzrq31du8SDNHPV7uIHYv+usnu087HT1Nj2H
qwjui+iyzZkUOsGqJszmkoKTZn90wT8QrgjzfG6GhYbJydhYBi4QiTrCPDJY2kKgsvqb/9sNc5Lh
Ap+UcQZ+Mk3cD0AWhH6NJsPcACQlT00+ZZLL2uQdZlSQZ/xCsYxy8S+20r5OovApDRgjZWF1+ulM
Qr8vzfeGTkejPZfiRf1zSizyWZId3Hi5seVJtX/+NK2IyIpce3VwRvszW6hyncmt0CvzJEWgI5th
YDCGq+EmJoyN4P9Vn4Gzzs9698RZHu23Zl0XL51fsS0iPHz1LPqf/0nimm9Ir221cTQLZIWmYhLy
ZOPOkQkSldKFsHbxxbzgQUphztgfZ30FH2v/EDY0TaSUyuaT3zTxxGe181lKEnoQ420yZthBGmvy
CnQ8o8E3JUikATLPuW67hOKa2lPfKQcIGohiLUr80s4+9N1fXyKaNUwbwU3dzPwjAOJfcznbU38z
HgCNbCb8P/794vn0RrI4M92XM/ij80LgF4qpgTBXujKdijkeZzGrMV7dSMfy9K3M5McsBViQLeyD
aggCoFIwTQeORCGvp0FWrmDkmJwU70jDs3ux8dfbZkpRDYOu7UP9bfU7g6dEZA0x5mXUkdTj3TXG
V3AZA9VxWSg9bsX1G0/0G5Ofxg+c5EYvlLyBOgirIZWV94YCcrmKVoRO6pc4ivgHlxrjHiFwvW0W
91bi5ovSCszyhLOHVrhR/ba9FepbHN9hCvGHy5XKIMMerQ94uK4N9wjN+kdwPAgHQ9rvSXM6LXxN
0aZhkQQ1jdU87S68aZ7JV6R0YUcGTwSszk/CBPVdgSc7g/XRixChUuV35fop+y7oDqRHJqjE2BwM
9HPDCt8EOcg1JR7bserCZqPrsH3Y4hgE8MuEMu7xmByMVBI2vk4GINM5aIp2ZE1w6x5NP6IwbIxr
gMFs5of7hqoxoPC0pBBXpQ2lMj54RrD4x/3PolUbA+ud5uvzfVEaf7c/8UirEY+ntdXbLJRpyg/Y
UgBqhxos7LukHkcq4AFq1VczOpZramJT7cyBjCpkh33ug5nM2nEOBW6emLCGcuYhgnl4mKwfuBw9
XmQMUcIG6aGOFWW6TGpZjzfGHCMJgeeEEemtR/qvCHXqvGXDIaxoODXZFziblbUxobVeCHYSo8Tt
X/HaPVzHBT3H8hlxkN82fU9iGbr1vzyB+KlYPpcaFb1dVAFPWNwtvEVf+m8QK4EtHtmjhJpPnn/+
FmIbkI2vfzJrYh9UZdk1AnIZCBGUlUAk2hwmpSZxrXOzyNYj0O6dU1TlLzXbpC8J1a/s9Dz0+E3g
hCb3hzDEwt73euqb4bETf6k64hyEi6XjEcZdQgKWHBi4HF58CPr8rKRx9oZW58xDjQjN7pX1WFFp
wdDkjMDclTXeXK/E3an4HJxj5nWf3bJyV6nZCMEay2iN0RaASBHwQKPAINrIRN1YOemoJ9PEp2R6
4IDSHF6AFLxyY8F13XrAdS+OmB3TsEv8szrA0REXBfLwl4Oa0dIq0GVujBvDjLdahWOXY317tZDk
eN3DxirVoCxeNu0t+VgfJMOHgJz/3ksdW6mKvnn3NX3of8929lzM0NzuxD2KfyXLNuCjcqFXb4ul
QWYo7oLf8WuH6Pcawy717K4fXhfHks7iqio24pT3c8CKOw1kKvysU+DJH50mKO9Nfbp4s6WgHLN2
kA1TDt8ufUoXep3zavMgGk1MTtjMCBw2xJCBFiEM4jPeyqTBeQ9BS+1+s7vIFrgS6Y6mEgEnQvXh
6d7kGvKL2ZN64qOKhifZWumvBwBHRHtzs+qhDI6FqzxlUMolGOcEArH/uRz6/hIjdHSk613SSqPk
n0M5V6IUtRRcREQxGkyz17ixpsDl7sZANfF525xvRYepjGQ+Oq/AcazUE2UtRUBil/+Zj5BMb4pI
REEMqTwvSpwqneaeFKyeBG9L6oFkoKHZm97FPcB9jlQBppUVoqm38RpqZhdo6qGXMfoJSahDoLsy
YlpQ7WIabL46XCHlJ7oZRnzAhDVnNOFBRo+QJY/GE6z+bER2A8+8CFnZylmk78zZg4R/7FBXFjeW
/Rybxh0I/RPbsdkRFuLnr9+4yVXHdBFX6EnG315XkcGcvOra6ZCV3chwd2ZVCUfbj8ox/kSNvCUQ
bWP7oCIjPAdikF1xf+ZeVyj2g+BQ4VIREMJ2Jr9djDjYCXrxDg1Nq7kwXA2k3jZSCoeoz6sSvBjd
4HpJaN5xHLyVLBcunyBk22grVro3vEa12X5LhG6FabS9VkIcyZKBacx/v9GJvEh66s+Gje0BssBW
IgcUE8/q4ZsexJDkmoUQ+TjeBVg1207VRWKSoy1Xfj0INo0ZrA7RxPj7dy0/yKplkuKyzCBu+10D
NwueosPqTLymaRg9Gx0A5Ns4yw6FDQfbFEI5mjsRwVQ0LCfsSO/mSgjwCWR5xXW4nnvsiT1ixc/e
uYpAV+oG8V1UVVtbc+CQeuwUc+pFOBFXhoJxadUiy2bhUEglFLmAbRL92I8jlK61V9JPdhbWAECk
0hlbkElT5Jgygt2UmY9VSdOmGeQA2Wspgu1SUk/8oP1dJYx16mfGkdRC8qDS8sPUCRUaUO4J6fgJ
bL6hgpglec+koiyBrgBGMir1+Pv4v/uRQM1Mt27Fs2UWulzwaZ2RrHCoYT2RkvT0gp+8A6lnWKkC
qR0Ma7jdnnu8FTvSdSdtuUb065asy5/bQQNT1ZHrKhidw74732yXRvLkpnkdv4eB8o0BGBFHrJeH
QBVmDO9m9++EWgBB2HnpTL0RQBaBbFmKE/VSAC5d/+0ymkU6GcK9JEat7ff5XfmdfK1BYlc3sFFz
SoAiqEkavaJ+Y2AIPUU9gb8FPoPQvc1JEJd13laIQgW9C3iUz19SXBLECLC5yYsqZut1Xh9hlVsz
G2jbXv26I7orePRy/qSlUQy5ytKKa4lAmQsGXcQSaVQavsYVoWO7XlrGRsdllTu88QhtByDP+MLh
AjXCPV22zPB1/t3TBjAPgnCgIQxeZ8UKL2MevPK9IUnMgsn7YjYR+bN2Os95sQia38BNMrEubE4N
e63DqMU90ay3ZsiPnrJGDtcDmWVg9YPjVW9/OTtfy0fk1MonBdUwxtTpjC27tb9Q0+Xi3FE43Afl
CvopLrfol6Gw+jgK9jKgXxpgGveOEy+YO3QXEkVIQ1rsmm8K8bap7qesgB4TF3tU/w7UxsWKEhpQ
MV+VBDj9J2UxOpwnx6JB+E/b6aqL4AGEaRRMOvSxGF68zhqThxTnZRReHakW2WBKT0aqbnhGdfxg
57pY2DDIV8iSObh/dH2uyUlqJok+BqEdy9/4wiA3M37RbrTlimb3JOe+BpHflX2DasC1TckK/LMG
f+qhJNeusPJb7RwWdnsqQUEdTt4qYrUC73IaXTt7dKzWVsYXTxCynqeKSgd26uOyjRg8rHdAj6w0
DarnLj4KcXdPjypB2EbGisJGM8IUXoZ0jh5CAEG/wsH0Qcea+GDEGV5K0qDDBCc0FfnC6E1g1WS6
n2M6/U8HRWKkUoYQ3fmALfCA9Fzv5fRxhB6ij62IzXzPwQIcPSnv1f7ZuC/Rvzhq9f8GgVMzI3Z7
Apnt7D4qzAODdcTN0O/lQU+JLCD9fALJzFPZLHoYzLNOf4BLgonqIRub/PzWNJTP6ygn1yaJ8pwW
lZt1fVZaaM4gPClI2F5nRrnTE1TxyVcVtOoP0ddES6HB6wr1LktpeHaep5ha6qt8FZtc3gnvcUJm
LmnZhVa7FBVDRYnJmWITaKGHD2mxeYv4lo5ZA0U2lM/lZjP/Sydy+O9FHWsxieu+Hq9GQF9Lrvcf
5Qg8VUOf+H9IwkVi8r8WlJOTSitG7MV2MCC/TnDWD28c/S3FXBvP21zIx3nYYDkTzgMQ14PXgyrH
5So9FYrYQD9qXwVfYCYVnD+guw2PXpi2PZCQfml49doPhRnHgzJsxYBm7pnj7gSbcvadD1XJqXFJ
HBVGiPh0XZmrFODnls8Wq6dNPEnkorVdVUYTyweeLFei+EFFpqti3FyRMYKCQiVJ0dDkkvzjwBrg
AqgCJ4SdNbKKMlT0Jl/NCkkUY1gqEu/iqnjUwJQBQdu9Qq0ql0TC/SeP0TXMa9C1Hx6sQxU1Rhbi
DGKu8610AfJbRC4W1PRuonLsiOKRmhw6gY6pkEojIMTYBKnb0nMh3ej9WZHjDEInE3qlP6TlMOUd
MKDs9wz16E09G5KOfySZOqH/UHtQMmROzOscr9ZwUoRVR05A2j+4cQJfmeME3imGukUh/RSjTSZ/
tDgZ3TFx8YWZngDd+id9yXbIIgDcrVEM+8ML238HsYfBOyKshaYuymdYSOMONDafs0mgCoanB22x
k2wiAYXgroHVXXFf+c4tR3TGEGZbplwzQCEpGyPTt/tGQ8iFd6P8mrTds9u+kbCe83CkIAjo7NA8
HUgtFKue5KEe7ooqeNXpKiCLc/onnltpG1T0WwDFu1ttmzaqaeNwCUAi+5Zb32YW+czmz9i+buIU
by7gjxkwryFNrFgUImbehVSErJBCyKEcY7bKlUMLEC5MkDbIVD5KytpT5GLPOWtZEy1I92mVqW2a
+FbUnR0pE4I6X/+6DuLjKyUA6FUdgzGW8kVn1MPPrlJknAq2FEMcqRKcAmBx5W0WUrQdAKuieZ/u
1zR0TU1nfkUdLaJlGyE20dRKtJMTQhHZBHgnOqBISIs1e1c3aRKFxjer6rL+C1wKNkn/7cC8le2l
RqmTYe+2OKIPe6cBqbeg6vm2gUAThSqgnNhwSdKvCc14wVKDOg23MbTRiN5Bs0OVyLfX2hK95AOU
J/9zqI/z0rdTUXmkTAp/1kFxbzYz0fc5AydZdTc7Cs27bRIAIFPsu5FaLb5VFZI3VECiJMEmJF8P
5vNvkHo4OaltBHL78eq1GNrR1CW1cir9WbiV16XZ96B25mh72t0f0tEMLQUfTkFJ45r9f+LKWwOg
6i4KQki1WpRA/tc+QkUFA/YrVds2WRIknoDx8hGWz4LfSWIS60wvQnINOW7x+5gto5V5QrMuud97
R2mR6KfSltLuSti8io5qvOZWtC2OZzyEifIHGqM1lItJ823jqyHkJt8gm+hNSv8IPZpML+72+t5n
6RJ1yQGeHRrRZHCIgTmV3Rg7Nh4R1Dw3I4aG4om9DLCGMqIOuqJEnnjOjwu5/4O8Pt290klKYMiM
PX9btitsFRRQpIfo3htrEM+lOdIxPhRFcEVgAMdLEcI90uTcU2+ij0WDG0mnpzOdb8Fofhc+Nxos
9zGE1Ea/pE0R3zlFMZgT46ScT9XjN+iKLYA0kl51BGf5EK4BcAJMLL4Cf9lGr65eLT+KoXrs8CV0
9tyj3MNoYQ9bmB2dvvHx5q19K+QknSjhbwnuQRBX/LcHGGlhn1b0OEW9z6nv/dYh8Okaoov8OzVT
KcBr23/RM++5iuNrLEzWn3bsJdm4V7U7psr13HVbg5Xtiweu0F6lz5giugJ9VGqh6PCL/3mgpd07
ExHaRP8ERjXwW26o5D3VWbGr9qoZIQDuiDt70yg41+oJxnrNQ0DZwi7JAoyhcaEDLQ/TMV7N0Onr
9OGcSG+zJUz9g429uO5oKd0GPvHVI9Zxz3H0kR7C3meGVpHwucUrNu30BEAo6daCdV3VoXGyWPQx
uqFVqCGcmbWmFVbNMP3qIpe+G38aEd0SOWcBEMU7MQ1hMCrUibSyWBDQIWbMroZlPeoIa9cHQsJV
9xBdesLrFncF0fcETjIWPKRhOGpip+8KEGZkXlDthYn6zA0Tx38rb2Fo76rXpDPK9F2QScH+WBlP
VC6+7Qr/E9Y6EXSG/YdmcpWV5WNobXVPHMtWuAV+4w9qQaufkdUImMURNjakpC1fLg0rdl8tENxn
P+nGU2x+udoaJerc9TdM69VhuAt4CWHK7Ua84Oq4QRP4pg+HPAVq4qTcAqRcJ6FD9M8JI3kQ1H7N
gxuWD/8CH/CVFf5O5jebulCxwFLxRk8Nb4674l+eHk/XVYJ8m+TyU5ym68o8skzRElFSm6wqrlhg
1mzQfyItVRUX2CWvKRc+rn0UlYLIhVW32pNixJJamUzD29QWhqk7sayKWqeq90ludjIpXBVMCnl1
P/bCLWGuU6KiPNUX4MBGzAqMGJdqsNsX8iZ1GFAUm6hU1cL7a/OfKPxg3Laud6UO6e7yZYeRN/ee
oR20zxl4RcyDGEdQ5ktKzDNeO6GW73EtjdvfJNL6+gzSQdd1BFKAetf07euEAe0feqj41Rx0ndE/
kyJOOLcZNnpETCswvDvqt/5YML61zwqw3vtBqnTVj1aNs3LrLCt4cEsrX86C5dyndeWNZG4pKzuI
DNi64aFFat/XBl8wsh/MxyYq6RtGFJJG+AV0Zozzh7oGQoyRHoxb1NoX2WzvVCemFBnGJiH5DItv
vAiCI1dUZEx0OYipZZBLKyzABXPeS84qm776TD3ctE3YFXEIAU8+QSMU6Sm8Z77BHOOACRfs19JV
L7OVKzQDJ+2/brB5Sa0l2Bpf4brD0CsmUnqXklXFIlbL2Z+0Yy/4ImtzpMoQO1qN9Yk0/tNqPFPF
Frx9MoZ/lX7p8l4UAjqCUiGy89mdQdwQ9LsgZHAB/KbU3EeUW+yxvPflDpI4D8TOVD4eh6HikK6F
uuZPPeNo1Do178jWEgoScJlb+iRkzmPTfol5pBH7Jh/Dwynv33b/yJ1J3J9fP6+7eES0aRHZrv3W
KbiRBjpgdZ+yAhCfRO7S+KF1hg7e+f52ahDhXLqiPoKVfI2OFT0kajBPnLxOxjfB41xU3+wxpdcg
+jnrwiVPPSM+DflZQBoiu3B4G1FEdwX2jSbXSzH8wasVin3L2gmiYqhaOYs34H76YTFsjjW4U7dP
ow66v8bpt9we2nd5R4/GLS4qALaTa3pmHFjpL/LXbFgo8y19X8e2uDso+PHur1cXPAHJ8EUZD+9b
7JvdXpI+53MIVhLfpNBZTCN7nzR262/uZ2oPTcys5kXU06HEZa5UHiQ8jeFkZHqo0FwqwSR9fJLi
ONJL49I2M2juL5w2tXu/eisSmzhhZyoGjP9FL94WTR3FidMNz8kYVVwpR2TJ+OG4BWbCWBtCalli
HmZrlNpkHKofpWPHBJ+1SpDXemdiW3Q9/Qs5No3DY46wE9wuQcgU0fYT/lvLphjz/0I7rK3SxhNM
Z3ZpfN7mIw+62EwgaDUuxcOBv5/Ue2T4Ak+TjclXGjdyHBJMnmAums3Cfpzns2MIv31XhPeOIubj
6EP/sk1Svmne4ArovHJK7TesCCRLgyGUPyiG0Ksg5TWX8ei0hbCDpWMXEPBGASt+6qXzemiGWYAY
ujuncb3KxKGE05AiIUw1Nd8WvcFFR6kTf1xWXDRb8BJemjnxm58jYMpiw+UPPAOfnShVxz5GSiUZ
NP4GYLIIhebpsFU+br+BLvTicjoE667QQUdpm4TiSwg5TIq3tHvg8soprNVJo+BQGFr3StJl2yW2
Kqac7VPxzydkGxJGGXEMpHn1pnHtwHaZ2H3BRE/KMaW82LaydSAKDas6tD+sPk7v/nAjeK6oveKR
DuVmgeZ+UPQ0J0jvWvX6NHvE1ZaxBPLYcw86LAXfQ8WeujV8DyGriZH9lGXRQf2y62S59EBGijBL
4w2OFMNVOFVaVMC+3mPcA6JGd6LS0oQcalW1Rbseib+78cFsEMjS0oO72VpuxQ6QovmVpDsb7ebn
DqbnmORzewzFfS9eFnYZdEQUHAXsc6dXIBGQDxOCmBxUAQwXBmpzjlDkeM20IU417wAmc8nIskRt
Bi2dme58//i1xLWAfrcjgk9f7V8I+69GiVjGgr9Ja+lHKWqj6wIDxWW6H+bXH9rtfQgyqHkuZaVj
ufrSbjDTfbQGO2Q1dI/t/fTcjhF9NKHO1e/++IPOOn/A22hal/GQu7GRLKDidObus725ynxJ38bV
2ZRmDViafgUyRuHG8/fcmeEp1dStCrOQCE1f5BrzS3kEmEtMQHySyv8ZeHS1wXVZnWLjcczhOLRY
Pm2hZFp/0qdmXu4C1xLMdbx1tuLVOE0sZRWiWisgSYvgfUkrtSjqKt47tYaxkRvGlKED+4XoY7cz
7NMzE78EiFiXsLXrqZNV3oAF4ZlbhuiCqE+yLZnXAiZx90IcDvb8s3qLbybJ/XDtj3yT+wF+owwx
roXRrGnFKEN49xdot9SFhoTMrWpgqQaM9rrezuMsk7LbdiM6+AjbPtygW0PFo2uNbb70TaogpwU6
1Wn74YJCwNOT+XNC8n/Uosa6SEIIzGYPNA0V7ipeOy20TkAUmfWpL8r8NLyEuwEg9gVT3bUu2kIP
JiqPbHpy6cRqymbuoLwIdeYCCf7rFW7Q/+k5HbUiKKfG5OeQIWDRkiQ+GQFRirKiIL/y3T16q9JV
Eb7Lkbv84Kss93UYwyKmj9HaViZkaJQk+fxIWlhYMaRoqk5xseT4Z5Dy1xBd8HAgatt9KCbK5BO6
OLFSNWH3BOChD6k9gzn4L8LWh1/C7OrJTVWyK/a2Qpo5s8xDoyfkugJb/ccxzdCy9kYQz0apxO/Z
VgHtKYbWWduVjvL7ECrldA3g/VCheFwhB7FewaeSGYeC2Gy0jp2/jZ3fWAVW2jBS1JmsDjET2I0K
oez1MeB82EMCVQo9Ym3qDgh5PLms/i8JFIfSEAWVTEWqPR0OXxHiH2/cICaG89ENysxofmndB2kA
otInw9Yc5ZVy4hQpkK1c08hB9o8UBAb0iFJ/VeyKJJR5WagX4vvUs6/5f6vJraMwnG5UBTuse+gd
zqxBbnoyDTRC6OAsppl8AHodZp79GliNl038JmH9/hsqSGL6bGb307fLJolq0boUs9sR3Bc9Yl5A
m4lrNm8xjp/oNbiuyvCH4ckFjavA3RZjV5k11t3QrrHIrTFCY23MUBY5Np5o5nbCAri9UGvcE6lz
R3Nj1T/l8Gqzp8eN8E0dkvHgb2PNQw9G4n1MbILlG1GdOYAGMpxyGfpKa5vfEoT+Sganfubwbf5k
Vz+3kWM/JbH83y8fKpcy5NbKy5rtopych7jQ8rGlHRR7atC7Es077XTr4sggT4mZvxLbtCHRWbD9
qvawvi5s9jv3uq34YsGGhoYX07PupCjcjUDIhwwL3onsRJZFr4ol/RgNw2gZ9KXoe5V2R0e6p6r8
wXPxBwbpDcp8q+mn2iivOnhT/AgWlhKMTafUAOVK2f9kBFjYSa4Jcct17eHlXmg6CPMTKA/IwLsG
45Zf0Lhlpr+D9xl6xdHlFe0rqtZYED68T7xeLt5nu1uoMbdRN6YDbpXE31mzNC2N36C8v1mQrtWA
0aOHhVXojjJKV6RXGo+uS1enmQNm+0tJJq+DXhsFksfIgsVOm20R1cDI1t+uz+RIQS4tGCcHIqo4
TK1eDQzU4KLn+AJtFHvuKLr/qbifwMQHQrqQx7sd82CHQxemnaJxt2zM1m0lAhfvIyO2wjBQkR2v
o8yjaSgmoBrbi1W4w+/y2xGOFHhPckDYXISJLAVJSu33Ie53pllK+gy/LeUjCrfy7M7EPkxtNJ6t
6/gqabbE8RwJ0zzLe92EE2wcKVvJZLZzvisdAMAsgEnX0UY8rOO1cq/l6G7i/wM8zNM3INfrijTM
t7plwOQqDq92TrnQs3uNCp7+hoXPf+Fe0Ajz9bKR3SuqqU+1Q8t8IXOuRrsn1/lMPJPwkA/jYROg
la46RB+F96WkyxJcUgiA8HFgF++uWe2G3ticozQvO9NHVIPfu4rhecctihPngtNmGhYi0j0SXak7
oMGD4CGFArNAxcR3JCzmXo37+ZvMpIPYBdrOADxsLx9JCzmRwYMSFddYAnU/ISYWWLEf7slVwjTd
nRX0szl5W0oZyPhLwmEmvZDrGJ2IKxMTVxZvYlqxMd2KOt/0owegTMJQF5ZiFu5hYzZ7kefQZl7C
4Q+0I6e3DZHHSycZhmKCN3vbA7Dh/FIqR4jas0Wkwp+3M4RE3skkNVZiCzer1viEVYNH8SNUk/ll
PyF98oIR66t6uBluT8pPBzaWnt36SdT7E2tdM1vWtvjcFtQSTktWDOSbRvjb6FGtGaaTbwUnsx1o
SZrDuMEgmGEOodCzNpWC486g9znwAPpHde51b99koB51dtIkUnUpHsH+nVMEIW2T2IV3V3Ulsdwe
7+d2hxYFdVkup1twSupNu46GOMMRjlJMFPSwraiN3OY+fDKPmmFPX5k7+exCKrLidJ1y7Yh8LFkn
cha8eAFjl3JsQ4rR5ouHXJqS/Gth8XzYA4/XrOy/J3u0mxJtvSLU8iwkm/4dj3JvRD5FegEMWX6l
fC8YsnOC7PTGMASB8ujO1v9xaWSPj3PwO8QPGXaLbcqC8OKiU2ZfBELYMYsJFris7Pl4f3Zsn0qw
p0Q3uouzEiNJD2QJEY0nEyMSJjxIIC3TKuWAKsDGcshHEinobTF2qMP+ruf3qN6JGqc8rOAqpIjj
O5WRoP0pocgJtTqcPBnI3Hlj/lgL/mgcbASCo8K5bX8FQJ5OGdEloPiNDURJ7rSTNfi8mXd2c0Fm
E+yni2mpfeeOrDIlo+TvTdr1rfJgyyMPTkHvTuxg16kT5LpiAH+T1ncI/8gSp6XMaAxn7C/h24EW
1YcONq6Br59d/KrNwl+EZP7sS2Tto5yRIl5uxleCH36ic5+YPmYWS8nMWH2S5gTr0dwKFKsgl+ca
Lam3d7xa1YPHs045k91+gjnWwbW6HS2ND/ZScYzGqpRObezeNBh1AExDJiNXUAVkXn102No+FFkJ
G5Kisg18EpCF9aLtImgVDOdfm72kmP7d5Y+DQjLnkzy4mdq+35fI5Kog1cNCp2y4NToDh6crX/pg
sZlQ/yvDRtZxzuM8aoH8tmE1Q/rLW2qRTZ6CrkrM/eSgpI2nHmorb0UCNHTSeXrLIRoAgynZcFyx
Xoe+LHI/CZ6lJBHL88xcwcLEUCXVfyoQsbpMTdqQi27A5TNc/fu8R8g8aIcFa7einjOZyJM7E6oE
GgCeQAmCl6j3QF2Doy5ur792updO5Br1KWfFJfqm3rHN1tLaIH7khJ2cu8Qw77qUiNd6DCiUfYfb
W67yUSelN7dQlml2RoOFzsc/s/ulLehAbIDExc2j2QyQkedn98axN5eLNvyQMAitTRmGvkxjYwzV
6eEv9nWr0OXMh21fsbg5QQUHDuvJcBjr/JEMpc50KzfhoecnB9wN5W6qoG+YCW5crpd7bN7SZGU7
PVUQgP2aI6GcWE3U2wgEXat/Hld39j4cLg4hxmCzhTZZuposz2MDLUZtvxQywc3rawLxIBzYBf9D
dQhRZPpJE1XLL+uFGrPXzdYnF/qMzm6RXq//zKwHNwmJIqrp9mIvVANThuzy4uHzV9cbcSJwFP+W
rUdZeWSeix7GcTCu2zF7ACvTnDkBIvYp3p4LZYrWw6vY3wliZSRO9wE0dH4iJSMnw5bAHBFCGhx/
cOfnaxBYkg+3eqZvwb1Wj7Min8+lZe/YOtPnbrLpLqsdSgFpG2z2DZX+vfHVk9PlGhget+1rFH/5
BJjvTo56b0y5etZLs4U31hKxeXMwMRqM/P/5Sd/fZtGpKtbLcy8X0MDa9GgO2V2ELO1cIWTEuU1y
msMyrtnPdNxFud4wgRoLiIEq4tf00jMTSLL8s+vy+zwddAmI9zeVoCQjzelHzXj4D1Fw5tAwdSQf
Hnj2I803Y+4NT4b+USLkF9cSwKpWPqEM2b3JSRaIufl1l8UWEghXLnQkXVzg+sIZZMPrwunV5wL2
oIIjVorUrzCWjimUYU6JdToMzOOyr2ViRrKYfqaPLu5jIJKlaaKd2lolYc9tSNQyy7OzQwHPOYNU
HsmwQxzrTs29F2uq0t2R6C3mKnSI/tXgYNevEIBTDT6n16yFjC801rHQUvcHfQg6Fh8EME0qhN1l
XxbUgTJtCB62Fn6qhgIRH6p+zj4/eiQWV2c/Xb+qdQTaKHONLaDNOiQQ4ujv/HGlUJeoI6XsGqMc
aQ1UiTR6TmXbXUamMXpUW7nOsc0CNazYb1q9l4X+EKeuVv4haR/HnwBNDTs6ji9ckREstOx2F5fH
s9RvOvSEVWiTcAuTn0JA6snrtDCJjUnC6eMJniYqDQqOs4ubi+0b0L1E0naJVDSZ80E7x4Ja+gcN
xe1s/7v4jbM6EfvlLsdFvxiMVJObTcAyuEJXmxCwOWRPSRQpL39HDyb+mazXe1pdFBKAXxXaoQDa
OJEDIt5dbQxmWFb+rie3QSEmq9pG+CM0k7VwwkcfpWF32eLM/mgiH7xO6QeyCr8DYL0o3UwfmmkH
+Z36Yp0BMDIbksD6W3CBjNoViRW7eLjXDt4HcRsacaykQNFg/rqdw3WScbiJ7twlptkts1H8Hx9+
oF0I+rLr+oftpKJa/I9NRZSQUX500YfRTrdKHu+/nfYSI5/mYJiK99vQmu+KKhqlf1No8BYAKgae
82+Up+E2E5ScBxp/pSvDJyEUWIXEXy6BeeYFiTzhTGilOk4cqe4DgHKfD1n3KJlaQ+rVxs1uLQb0
MvUw6V8Nk0J0ppHgjbBFgu6IWZ9Ya6ACrPgAYxKlaMbK413YA2m0t95HqTwCwceY5yKDl4eX9FIq
r+iXUulAvCgfbP4OgTR/ngzMBWrogsc9gavkKxA8EVZegbzpwMwzgcgJ+iPCUfa1pkueBzUwKuyY
1rmLwqL7WxRQBkDlEqhRD3Xd22ImHAGCJpF3OC/KYvVYJfUep5DeRNr/JYj+RLUTn7qcZ9u1xXvu
ycJ/sGPXtihQAR6wMHyIW5yOw3o6278AbmLSMYNvCB2W/7++0U0o/oBtxB7IVVzktHHnKr6vGMug
H44fxs7+EicxuTtVW2YUPw/0ARwooEhjiXYgfWMa4M9kkJlc6mZMOcW0tq/MjRTLwmHAOGpIogLY
d7DJipQhGN9RoMewNc+nZLz7aZ9QhYV7SSdqdqc5GlLT5Wnol5tQ7iUc3bI1d875sg9Znps+K6mw
N+rBFaRC2j44drM4kXQ5X7Z6PNrh5akBV5Xlsb9accumxN1oaCGXO4e7PY92za+ehFty/dyTczPt
eLNJ7iTd+d/3YCHLUnp/8BHZt+V5J8FOL44aZaGXixYPtZBYxvcEYl2xzZvsBVDKVR/cZVBc/prW
xBTXqB4sq3pvVxNtY8OX0HyOXTuhPKqEGMjAqezf3GpSksqvRIQ/1Z/XX8T/UAHeV/zWRBGGRY3l
1uGp1jWAoy1oy5rdHRkT+0caNXcbDkzd1ZoJr+94UGM9kQaEz8tLrI2vUje/t9WtHSNUPRL6RHpa
7V4UQ9sM9ELwN8p2loZFPachNW+04uGV07Y3SQkHf3vKviXZgcPvgCO5ooBcgi3p/yJbVwBi8/FF
Vn9Jgj/YtAaLgDyJoDGv2jaYLnot1IgqylLnmZrplXU8rn/DJRNQ3Cj3KsHYKbfbgkxqnxxwoUvN
vLewE8dxC6SjBF2sdZ49ryuW9vfSk1sSIifPQSusNhhu2UgYK8zpVDIQQe4JGeesaWOS3r3OGj3P
L4WMtfyFAonMiyiwd4V8HYW27AKAGvpOEeYZ9EBaHngq8tEgREU55qUiWzB+3ndIq3fdktWMjtqW
1JwxGxFbaTWdKSMLWRCcrYQ6ynEvfdvOw/hkhgFcV1JObfaoQ4ZFADOx8VJaYhUzqbeWSuz/LH0w
XkFcdEOBvpGUiCjvjcLSWHPfmzR1801Os0/5DPOYhn95Da+/21LN/qO5Gi/oW1K7RIGPLhP2xOLu
y1wXLGeS+vexmDLnaDdH+eX1e9AzpX5Adjxndy7pOQnvolyWXTvzaSmcTkfqxjmyHnWIv5iysYKK
IjLF1kmuqVS0AFodPlZ7EYxyPGGyEkxp2mVOUR6D8wHF4ZrecAitkvuLdzYbZ2za4I1qIE9b4q8f
tQHcO8TaBoKCfq73j636Mo/Nf/50R0ZwyoCbEIJBnQVRFs1xLSNCtOAJRj0ui319a8xClGulw3QC
Lf1RDbn07iammTOEgDefrYpDSwq/ns9GTeGPVZHGN6WyLw5u7Wx9YMeT5ZXEwv3PYYZJspKxD8IT
IBM3GubFHlP3oHh0xy5PFtB8lGoSScSIGDOCqijgeAtUS/2GvFC+JUnowy7xY119d1PPQjVAMjqY
Wxoo1r1e20nWuPsYblIcltsi+oeVD6iLo/1Q12jKf+afQKN6a8GxqZ2ilSDdHUMMRf8pBYmnKLea
i6jOmqd32j0neaYh2Ng1epG8WkR4hYR0p6t/sDvpLLW38LNlA/4UXpvZlQVjuu3bG2VFJ9p2vAvW
NfMRgcUIASGwqDy9N8ZXRB9NbSzHHuLFpWGlAzlBKLabCjRBD348EOqA/A1oJMZ7/4cqijNbvYqP
T7NKdne5r64HUZW+0sEiK2J8mqucbwWb9JgbTAK4/r7jNU4Tm90pY9DDomeMdVRBQrmqDou61/7U
zMPuTV+DF8MkJBUtb8XcxK0zSjrs0SjqQ8TtGPpXkORejbVllklpzaT57u6wxL03pMohK80vwCjQ
jW/KfX3vxPAyzKkzTRWdAqaIZpGTW4HkEsuxWW6CfcxLGMO8obFEWRMy+aXJoSj5k5mq6DiNIx6d
p8CWm2RQyAyMoC1QmCjhRDlx+Yv6GRmJ/p+JEF2KqDuBaD0cbvBOFDpw7hYVcTeCReThTUUOhfNe
l2+eB68qiPlqRH0EoVuv8exV9eljBJAzWrWKQWTW6ZwJDLR4A2ya9tvRQmAdVASLd7GqDhfZ/TAf
mDV1PnR+/fkdsW33Wqvncrf+vej/Bx51iwh+pyWA6f2oRiZ9LrvbZ67rE4BWOAsM8RTcID+fSnhg
hhivWFgQZO3Z44r5ArEhZQSgTMtVdtRXO5xls1gl1hWSZl6IsRLi+emu3kxJQPwvcNaPN7UJSYJf
dRe+b1do8LNA4zLAJKYoPGZgfyhc4d0lpyMcolE8rOuWb7Cx7FBEyaShFoNE7rVUBubpvoeL/SjY
AKsNxSHepGalvSoiQBSDfFfnDPYRW1ev7zrT9N74mxClSzPp/8XpbcncKMfoQC7tPVxM+i8PXTSc
kh8P90FUl47ZV/3+l/lEolgfu5s8QuVQmHkhGYGx3BwuE3+0e240cXoT38K+9bGYOVjrRoXd0xmP
nEra9vaPwOdl08xn5NovnPIYDOWOq0Z/0bnhhEQktidyPEhrLuV365abzxJvRwgKYT+LkDIierJj
E8m0aq+e77UK39dmHCFP/j1a5quLyz8xexDZRHD1AGSqnHlt2LXA5TJuZRx6W3413aSrKc4fZgKu
+K7MeteFuQuUv6OjcKOAWckuSmHeKnHeOW3Fpe2wyC8UCOSAyUWVbvSYr8BS6CjziD0mohlbKk/2
D+ba3eD119hjefdKVUf+iJIvphjorIBV0zM8yRZv2NEXv3z1J+rLfD0VS/xhd5ib7GLpQbAUNwcI
6ZTyS9YLrj4FUAcGnypa6Sx19P/ZSijsnwFLSLdiDROfIX5LPsRkKLgq0jyW0Ilh27RwnkZ60DiD
uqD24PhnncPPLKvO83F3i41WmZyHXRbAK6Uj8MmWF+ZJ/OoLCSmFeHvzeRjrq9WjDlema0+t36R7
ppM0djbO/RQStL/beFtD/VWKw3yQULxK76A7yV0x/BJeBoA2AHlw+dwQbryC+JNQkXbgA9HDCY9c
hPpvmE2LpW+DNb9OPcaUHw3AdSu/I6COIqt8D7xpNZ5yfo1keRI2PLau7NVmC0x3kgKUFMGcoRSa
i+D8Oprpcr2JO3r8s6/WM2cSMj05kkT7ORW2DDS8uUNTAQ13tw9jMPLwEXcmH0ftlsgMubd6PV7U
84YlmQNDWx7XspgJ623rFA8WQNZzP+TOAAS8dO2lUU8vbwoN+uSJM9TQcuGb9j6IXS0tkC7Mxc9O
/AToYzK3o6I6rqf9uS9G+dowkTHku5pLd2yGk+BkjlZ4iC3kBzbORu17iXvbJYCQsCgcwpK6YabG
BmRTds2r1ZrDZitUz7vSPl8mM698pjkbkQcCBkv2JPshQ59OqrmcdALL42RcE+dd9i69+K1uROCw
GZYJbTFmHXWbwKTZbd3AKFsJ+7fOgOWJSOCFB5CoIc+mqez3lm8txoG7MtL/x0al1DwtBmtNIRjc
AMaXtWi/m6N57P6QiZwQjNTQlx267EsscaINUVr+J/y8YHJmhhiBEUI1VWIX1d4Wx9sYH3kdSu5p
nbuvGrk6O+lgsbj+r0BCgIk4BYJzlsJVAjSHxp00V8z+1fx/nneT4XSuN1XF4+YC86V7EL/ff5qL
ylbt0EPkURVx8YbxsvdNOVhnua5CB+1yxjAMw2cvML+fY/HRjQQL2LomUWE+nC7eAf/ik1fd9ExX
KukylR8PLG4/aVFL04Sv5tG2l43NEVABjSHLCCFbOJL1s0Mg+lGLMWhgVHcbRzL+0pBB3CS6su6F
h+HhmHMz3VHY0Yn2rA8dGexpNQvcfenjw2rKBJULjaw0g+Wew9GwQa3EliBDDohIEulyxFZzWekC
ICsEX1PUat5MHZrbu6QaQGeL6ql6UOXJYgKj9XSfJxdUhu+2PXm+EGIppYLB/2jTx6voiNiKDukR
AfnwROsMtf02qdCedcQpHh5cc3uhtePNdUqJNElXy4lUuxdJW45g4Nywib4jYsFGPRgoXO3B59Ck
I6mgD13YjRuK/RtZ8UIKNmkZ6mMeAo6U2Z9hFpJBg7eniFZiYqNjTITiqex/L9M/y2nupXaWmGTB
XSc27Uulz0w3pRou/y8IenNhgQJKKuB70usaxbN4CPmkmgxIxkvg+vWfbOikSOcg8/LhOZRN1fNj
lFsOFfECty6uvOnhb1kvlmnhlhv9gmlE0igjt6nqiJwfD1v6memv4kpX8aWklZZJ9EZTjlyuSUGY
NbUwHOsWbllA/2gedEHV0tDrMvsqmsqz8NPqp3yH8iG6SbhTTJM3bQ1OpfkCsMTgCWlDOBLKlX1R
pFM1Gd3HSffKl6VyI6LOT4UT1Pnq0UmzNdyFHle6zwMPR5Vnt0Qq7IttE+8Ce4KO8reEO/P1BRPI
+lVNrjnPI8IT89feFgtKbmPwqTQlgo8Lp42coUxCVdlol255uazB1vRkcdR6AKQi/bhTcAkagNME
JeV9mvOKTWsEb2bspjfB9fN48u1PzXom+YI4QncXQxgWqwtsmIdzbtoS6wwquwN7f/yvmBsJu8IL
InrEYLiwtPSTHwyLjE7VewGqarmPlIhOBo2cZMDxJM9ew4+L9HfV2NgLlmk9yse/J+OVpR2rLOoN
Fo281gbHpNY+n3XOgG+W90z5M/CxgC+PgkYVdWspHELTbjbZ/IWloDRZ0tgmEFWGJ9f4/Sf9DJZ+
gnkhblsoAyKjQqjMz7BhTkAVCz9CJOMbk30X2PV6QSW28InsssVXTUEP5Gpx5nwOcPq5xi1AI0Cc
Ope4gINNG80JGHAbf5iHjrFkiTL+rTl4sK4S7qub8YaNnpU6a9pPd91OOVYmdzy54l+5xPaq/JI5
2e9P7SNtJ1+2FEdwp8wg9KHq7CC/bYGlNDGW4924H6wuxd37Ss3Tm0iiClLCZMYnPZwOzG+N9ZyJ
ui3NfSoSoetuORuqI2SzTcIHKFiRUVLM/rmYY0YOWLebZJ45vKDD3pLJISXliBLl6zr13aKHl1Aa
ilnJS/m238BQOk5ZwjXDs/dvq3sNglLVho3PEzEnN7Vk1jLxDSJwl9b8ts3e0UB/H74bXyda9yG8
fwlkfOrFr303t5qSxrxEge43XdsGYW/kHyaiwZjZK6qxvd1ZNIT0D+w5ADLTx3a/IzC/qQHHRVQl
sVGfuEUHPYGxTDfHBxpn8WN49WG41XxATBZQjFCyJw2llt8lB60vdBA1BOONkyxvlenzmfN0MzbI
lRnMZN3SjCSKmUBEw5d5/+jyN0LXeTn+lUqa20uj16DgiM1ZoN35YFKynKd6VtMt4cgf7lHA1Ws/
78d+YiDKRue4qL8LwF8t0qNfvILeSq0jD6TrvxxKmFvyyxDUpG54bGzUMrLeyTgnAYA+sSYK2f3l
yziuRkjApk6kOsoNxcDTMKlKi6BP3oM4ptYEwg8I/XuwIUdPiAOZGnt/g3u4WobNo+VaiOvl2pZ2
zawfzWl0l41rZijpjguE+YABll4hK2Ou0eKtHBWoabtQ9exc8IH3dUkPRpUCRhpRUJv/8Fkx+Kuj
uMeptbukUZejjTSnCsVnRVV4TfIRiDfVtaRZb4InsUvFMcy4iWcffcCc5mSEzZ+fMGjwaZRjVa4q
bxcfZqkaTa11jePAP8Bt9kmORvb/xoGcg8pPjdW/sVPl4idiYoUXnslce+xcKPu7EirCRB3bDMoS
rpHkgxc88KXESQhJgHRBLqjs1Eq1//u3184NAwnc+rJaRENvpyehRjL0RBnQmV1V4blPhpZOahwA
TmWAx/glKpcyINVNHH5KWo0jlg2vyYzzH9+NKk0qdl6YBz+rrahpSBGzMQdNv0s4GG+c1VdB02Zb
MlEW+e4g9Lx/UQwcVtGLYCGsK+cQ2l6mgm9CWzC+zOp94NTGvUq6W2XPyN/5JAHTXrnbmCbgqZVa
Yao1WnndOWRQ87vPMq3schrjTq2SSJ/kpaN6JJXHzFuCou6z78hVa4TZyQrbNOU+kUY6APiczhT0
XMBTMhLTaIVi2X75D5E1SiPlcWkTh5QgFYebY3zMg3PBeB+IsoN5gcYt3WYIj6gGLnEv6HQGP0h/
qeP6ukGe91gNhZjsUnYO9q7O9yPDFuD/ZPPtOCczhI5aK1BW8SsdgpiUnM+0aL17152qUNLniiIi
QEse2qLah/41uI3cNBsmxUqn9NCWjiHPAYxGlF9DULeJjHSLrNDQD6yHOh0UYoNx2vcKae4lkbsA
a8PA7hskdC/rHiqEHKKlSqsFB1pEMH+dRV3+IPPsLbhpqQxltEDPnj9i+8rQa8/4o1bA+FuzPMpm
1sDDxHwQd+CxiPjA4ZhsCODiAkA3k3VhOBRo8/WTxP1e6cH4gZkzsGTQSnZcERWOBViuECAiytcY
DMHiENaYiKXk75tqTZ9QaiK8cr99bcdSerShkuSeMkv+MCMmmFYjrNmgwzUuMuugoGAbdFEfPznh
TRbojXQpv22nzsU5+qHgrfap8GS2Exxve6jBvOzw5Q1rAi9mPjmG72qhbRTiLhJQ9fxA+dtRlnn5
Ei+Zul5+vkHRsBEYMi5oH9SM8SnKLrL1OAuNJBSgDSHjmQw0QYzh9RK7v7BGDYSBEX74sv9qldCo
w64zsgOoGFYgBz9wDbX72gYPQtLfssnOUXWqdEnDrh4bKbRFdpoKY6JJLakFBeBemkfcJ9XXXYpf
JmWkA+ONvUN7eu8Lwl2V2hgy7Fcvx6Oq9OxPWrTYv/tYY2bAWWwKI0+ayZQcij17cn9E8qM1xAE/
d05JZ68tvbTR7V9aF6HxLEvI5i8UYRCvvqOlETRBAqPKgO1XDwUfW+bzv0bdCC5jcC8xXf44vbCK
KNzMgD2FkjzEXJsa8xmJfM/3YAJbI4zcYA4/c2XTt8tTBpv1ge6Vi6c0tQha59cvMr6mVrZYTUrU
Xz3KDOe7bYIbwe8MaGqlT4pLU8mbqO4xT9m13VcNMrYewedqNK3YDbX7tRvSb7DzaSYK/NHhTrtN
jhsJtpE6y3mCVSxUe1kaqYEAtyCDdFfNXT+IjCFTCbcoiHhSnA68T14AZqQxYjSX9Z2BklVVnK44
AnjaRGNcA2Caj6oJkKGo3Geb61w2Uhw3RYLtHv43roB9rMcN0/Qkqnyg6XODqzQv9GlfQcYGsaYh
VHyQClnMuWgQ4TDZaGiMfxuVnkIRirk42zsiRgYk0TAbfku7WzIB3PUTN1y/wcLuqCvswF93muNY
CtyB+Q185qC3YGEDDCdPBAlgUML3URWrvKVOsWShycHZIL6vW3EwHtjIi103NY+SiW/QCwRJPacx
QYgjqDAf5HiKAcI6ZLL+82nkKqtcXRE6VgMwBeFUQFNli5FC4WxLpaWeiJrTShnlUg08Xo/xY2RD
h9S8EzkXzn9Gq/vPD7CScettZkLDPtwMevNX+z7U/yHABhV66369qe67ZZ8VO1PMBewLP7A0a+Zd
aqlV357yDqoyRr3Qab2r1pmlMqwuketzGahMA4Flim0BHejsbT/1zG5KIGuu+Kurc78X/Uaa5BqX
d9V3QEZB5yQNSnSD3OR8iM8RXMVI2ntgPMp62YHeD6jnlBHA8/VojrpVvcfODyHlPuRL6IzTdP3L
VPZna+3H+wGHlZLwJXhkOfVIIuNULDZAVyUPnAyFTpPss0QdSScD9OECdbNs2e4A71sVhLK1Gth/
1m9EbivybcdMVEb3lRGuWCt/0P4l0JKMYRJqMn61Gnht419dYX/zm8kuKDi0Amq0TtWFBUG6OeYr
U1NIv4D89VY36aGsFHSB2qaZYT7RNnJ4Da2uvzOQrHMp0+30EABllgVGLc0SFGC0jDYJQ9eJkTKr
yq4U3GDQ9iv4I7J8HI8U8Pbb8i/jHn38h5sIN2Owt0u5bJBxLsPGK4tOmGQUr6ZnyR+nQDfBU3Vg
43q/Hm0fZl5pC2KpPcq7GgQu6nBgXVJTSEi59CjqyxEL2CIgrr90iYlN4aX2GBCKME0LVJ1LtR7f
b59BbAP+a9rq4zTnRY12YRK2TaK7xm1QeffwbGE6ka5SKTxt+Sup2wxiHiP6NA05FQJsOk6AAAOL
xVjIY0isd5d8YMEu/g6f8T0l338Ig8EkEsYOjZ8nazEc9V9CrlhUBQX/7BUXzyESd6o0AYRXWOb2
pqe/WvB50C1TfGLHPZ9Oz3jPn9kAxXpkYKthR2PRWKSVp4WPZ/fAJwHl2QFWH4mER6LLk6ZywXP1
xFDg+kbhc3ef26H3AOfaFKgirR20KUA952Aq2IOIMYVuYOYUs80xXEsnMCDEx7KF4nDGNmFdTio1
bpJfYvGQz8Xb35NvsLkhaWzBTLms7X46AI6TBIcT5Liz+5UlIBOXDRswN06xLqadrSlsnOWWYnCz
cODTuA5Z+93EN1aIughCkcxHNj++cVY/aYRWZ6yIpNS05UlPseWmLurtyc3Kmg/jUFvfZuR0NVRM
rXykEn0MQxoCEEOcH3NpL5pkip3XoxVXP9QP2YJjG/hZ3l/QrvCite9GZEVB6ewW9aYiqfNK4iQP
mp36Rdr7lx/XUXQNu7Q1w4ESnnFuXTyD2UDoZV5xhJtX9py4FIiRutiIUmcdm2UIjX8i5ZHl/k7N
aVijL21zjZSDHzu6WJjZ6p5QYcEyQGMAvAYuKQup1hZJ1cG9AehSIgZbB4fyIKfpxnT7v4qQW01G
VYl27ryZO5SUQfpRaidnZaBhPmeNpSIV3We18HZtcvsPgnizOa/bnzb4Niah39RW4Ee2yEPos4nF
2/S/BTOtAYXnTBCdEA2pm/N38vJJMjaGuQANhJB4SEKQlKZcURH0WFB2e8vaEmBcF2Z//vejfQFK
scSCXy/uXPff6AyhcQ7Sapmzuicvp6faqeberVl/ZqT9Hsk/+SVo5mMAHkAcLyFF5xlobT3ijYFJ
V8PAoafs44N++avBM98oBZu0vQ+2O/YNaJQUpAHZ+Y3TE0jg6l3+CIOcqTAFC6FqdJ6AkZ+n9VoR
sxYfHt3200rjR3w/0GjJV04Pw7N8zvWz2r1tSYh1hs9vQZzJn8VHaE4xec0LuNSyf7iF3eJFN9yU
JQ3dFU3AllMCgADY85YuKUA3e04305p1i3InOoTAqtHOH3+RRMzENWiiAtPXTeutNAf3RmFSTu6u
AT8M0rF7pHch/SpTADEIEyybMvp4yUMcOYxdDK1a5lJLSA2KL2H2k5v7/m4Mpx7MeDSDfqG7pyWD
6cm/6GFXG6qbTk+QOWhCSOkUn314mmT5mktok/TL9SOxPLBt79baC3CHf5uWAb92ItQ+WA9ziywx
18/qszlzs+lDzV9Jt8vUgdlJNva4FCbK57dyc6ZmJWeLI33ro/fezuufloB1EbMn6/HeExXPQI+1
TJtb1rfRKRXudwMgIH7RgcsrdQRIIqFyJNKzA1PXcaQdBf2BVR5Zd0paEvDecOopXfLNKEAt4tQL
fl0KmMifkZmnrNMfJOTcps21GcoQivaPjgJreswj19J85I902ZsVlwOIIrpJ+coaJxrlNLlyicAr
8NHYyiRCR3D+Z+UDUDN0UL+j39AOk4xpPRiiln2LgmtHwy/NQ/qRAkQto8Cp9zaFu8qVbv1WxAlC
eMquXlgKiUriK2d3ST/dUvnC2y8Zt41+5eWEOJq/50iyP/xf6dxfaUuTEqEMmvUZhvIfpHgusHd2
7onelyChnd1fYarJkTo7+QFHip7oDM2vUf5TTJoeGR+Ch5TVypX7QiR+j3mdfGUDuNEpsHE4kUOL
uOH7hSAz3kiUGO9h10SqHfXO1D/q9v3dXdAxBb9Y/7/gi/P2esRPm5j6SxwLcgAUGgYRjuzvCP0P
EXeSG5zVGOJ3+DYkhNKhGgD3qbfv+d+0KE7lAQH0spAwSFT+iRfJpnXkIwwgRBRi7h7fm8JhrEHc
+B+YKCiAJYeekvWCibb4UAK6y5Dba6R0uIucVnZtx2wo/uvBlHuxraCwPGMjgZ02fwRAFO7rvhgf
Z5FKZYeJ4ov7VIr4ThjlTOUp4x87RnJf1l3A2ykpTceCHpKTXhHjH+euzBq52CX1SHtiqW7a+SAT
u7s7PdK5lmfMskAAFoK2/vpE5d98B9roYZJLNXtNVGaS3d0kA4OLMAhufxMv2SwfDuD+k2tHNkKU
Igb8JVZmWjTzHmrDmVCiFYrsQ/K7c2h8XYrVMueIvS4QAvcT6VmTzl1MjXqCFRZWtmxq4G5vjOMP
lRXGLllQYJ6eI2bzaxvFFYo65DIlcemf7HTu48ZMAE+WRgxcICBiSERdHR5qb1ovLdTrF354Dw/M
lDL3a6C7qP4RrJaVBOlnaE8lgrE/QFAj86jWqcOPWUEnPEMjq/L7soPBbZmNOfSylGshgGp1Tj36
QH1LQDQM5JWrQcog807lCdcVok4CsF245bkw1iL7/U5O15ZJG7HMMp28QKmiqxpK8NzyCQ65Sna3
5VPXEiIXAXHH3A830EwYUnr6KR7OzncDS3soI5PZELeWG6W60P7VXdAZqRP4RAu61afrp3urHLcH
C2qoub1Hw2Q/apqe/sFU028iuZjuIMmDrcJl8mu3aiuzpJHMKGv/oYqNc0VYjWcjxdznSgia8ClV
lw5dzUyT5qhZ6sPQXALOLTx5Kuq5vSMOITzDIs8rym1wvGFG3fDSAzQq6IL6KmAWMBJT7tZHH1xG
dsvi1oTHs4KliizOkzdnnjxvN1s5Fxt9jwpatG+//GTZUVOOuBFWWkLAEw2bKaRH0+jQi5MhiUlB
7YaOSwYa61NVzuWnrBcyzJWuWGyduQ3mtggCExbcoQMysqNEUt6WzQvbx/lYV7Q53hRWjkZ3O5pb
aTpoNJe/EifkHrf3nQd/pDrlvvxjSBa8wIFihSsUuY69786mn2KlaGIPfqIWTBKwFbT7c1bEoKS3
KkuscZ4Lr82kCTIi+z0Su9F4N8QJWKF8SuQbqpEAMlOuSxzfgsT4632iqBnbhpChvEc4rV+ZOtnk
TAt0xCmo0sk+2R2ZK6HFZC1mRoYS0JqmwUATcNGAesC5EtxSD7NTmjo8B/mm+8vuzFpVe6gHGcXk
1Qegbyt/LbhhPhx12FRGdW4SldvwysqRc9QPtSirmWldWKqoEPrq2TQFBprwaQqBX4gtNU7OwTzu
N0w0tf3WFO2oa4xutpyxxUMlIvk1FFdRvGYWFZ3hHt8ycWjWAd9s73rxITV8c2jTFEWb3l6vHKam
gDlWM48571z+OjX+mJwvuai0svhgHFETqP482K/DE/17jQ6f9rbvINRCUbSNBp1L6g/FDdJ8ZcjM
m7M2HihFnNT52uvlr4eMxGGq14jNE4gNpHPGqt/n7tg+Q/gr8uspMFENUPAl5zpb0ZnN2nF8qfBe
/8Kl5/aRjVGjfpT4/OLOCzVSGRhcOkS+8umF9Z5C98pRV6GrlrCKzUT6X1Q9u13toaX1Sg9ZJYRt
KF1lAI3ikSMYJHtzZgbxKh/yCQfExsk8zy/G7W7yxzbl/QZs3GQn8qY3Cw1SjG8hoOi/muF1GnYC
fxH/rtjgvkaaCDw+Z4fZWQkUL/5mY+hDHvWoxmHWO6upHFyN+7H/8cM+fTuI/Dc+gxYdtkB9otVn
FCl3QjygyX6QI9hs7bUlZBI+b1n3fIiaS4m6smelD7PP503iVqwVS80xydGgT3l+pY7lh3JnyeIb
YHn35KwdB3/uG5xOHZ1zpSJhVLF0//SgIZE4GBn0ODUgnfg85d+yccL6y1AKDvM+9gry7D+te8r2
HbDeYblx+2TNgeeMmjRJ7BBgulmbqpRt0OrBoL2bVTbVHUNb5V6DSFnIh0Tz0Y2hZB8qmX4+B+ca
LhG7My0tCkANBezw/qCkQVkaEEQnjgWfWuf9OuMEgGKLxrXgmGwNqPLFDAH/DH+C4eszGtxuuoL0
ywFrDHpeC5zgUMeuGFCNZboKPbak8uL56h/+WBqreSB9sqK3WFS2Kc4TRdPnyLNNgyzNS051gZag
jzbrBXL6TgTdwMXHRhTTQP8J0Gt2ZnQIerCRGyuWk67vgqNfyaX6DIcROfmo2JFwLFpUzCOQhqto
/NEyVG2zQ1ZXofxKvoSsVL0Lz1Q7W8rqMzK06U/WrrHFrIaWl58Z/j3YzH9Lx2PP+TH+gwAHccHC
ZS5fnvd79zBPvNphT4kK25XIrIgcgW0ppLeACoD05ZKLrDTMRPiOxC5Pz7ckNALeAaPIy0Yj1T1x
7D72Fzrqxq1zVjQemWN6iOV4YFD1aSuRcKFTK/ZBDLxsA4Ae/586ShYoSx7uho772xQS24rJq1Zq
7SxAs96vlK1qhgZXim+6/rVZS6kVP0nfpKyE21FgF10zdfavjcdjEjYWOWwI9uJY/x3yXU5+hW38
fT7prCBlNp1kPPa5T6DmieWQ2nZP5R94hCPo8Qwup7UD1l+0GCxSw49UZx069OzEqa+BIKsY0fmY
lPuriw2HFizeLwVILzjWPJAaktjPpzM15AO8PXqfPYKXkJ9us9TWiQiR8xgGm2XsdvZv+WSe74DL
FZ/oi1CosAytVylLDcWhstC1WHqSJnOyLF4A1aRkP59e6FHrpxYh52rxBgAoqzQ11E+53upsjYkD
XdTqB93Y0KTFU4A46LWwbLbziWUydPkl6DDIlJ9mGgHwS7IQlQxhyc2t2LTfKi4rgyLQANkpsQPs
PGNvccXxHGxnRsYe+0MJfyNNrSbS2BqtBBmF8TB5aCsrqrpIVcJAh7i6ozC2DwLKlXv5FBwvMZZU
otgRSjyLdNFsqwZrTZohSy44dFE6qID4UAeGk14J7Sg28ASaEzcNr1GQ/iEJrzm3Pk60RB1m5wX+
CH7pfXuxWHtuTzHOGXKrf+HXHYz7lCcdjB6oFDF/97nXXFO0pm3S674JS8YhY+qgmyXIDL30+6qK
hbkpA1zlIdNAOKALbrQwYBXa6K4gFRXAXHcjjxXnU6RZpXbsi8YORyenE28LPPfQZWcXS0mCWEF2
OroNeSflBj7no3Uhtl0qr7+gmFbT3/hZ1L88hjo5cOw6XuChE3R/N+jXTk+AvsYYjyIRjb2kmQlU
LYIaFT8Yew==
`protect end_protected

