

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ahdDAHzz440n+Z6SrLNKLMBChQ5FzHxmtmolGyaGzRzZ6AsdM11MYnHQlmkXolfzuQvsH0tiYFpA
bdhL84ynJQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qd5Te5HYUFbAOVCK7Nrwmf+xhp7iHLV1qESGeKRRemMuPlhm9gxKzGI5glBpEm+Bt6GS7xBHPesU
Rh2RxY+9Nst/QoTZG24XGDjT8gulIAFW/37G7vhPLNVOq1gP33zQ0iNDRVgAsbEBqL2aP8fzO3c4
Dl1oSNusYXsdFmxhv/4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0n9Q8CLs0GcRArqoXB7pbLNq/7iI54QAnaQ3YfVTrcoLuaPhMipi/u1YxvxCeQhStE/q36RmAWKU
vuVvb8WRD5dX8Gc/5jIRt4ORXRhrtme6cizBVjYhymzdNTAgbAuH8k+0No3YXlnw3iXuB/bUUXlS
9ThgyMn0i7erFTJ6h/eogbI8EG6TwEBPQ11D5xXxMjzz9Q1WQ4L1w3R2CAYnCrSSlQxqvapc2X6+
HzE5EzvdMpbru1PQrGeGwaFtvlT4dq9BRwJcYQeIth/77QtTOb09uuY2bIUtRjnczrx+97he8zc4
F2HQqnZwdLvPbSwwqlsUdlME2ell5wSO2A8Cdw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fXi1UCgHICyjHcoUzs2uXfr4QL3Zd6fFq0YYnh7DHj/Uz2hpTBP/xGkihvbT84E9/Kgj7lZnbxyU
NW3Mn3WgobnvsYj6dHFEG2LfnPYpGw5nhTQMawWoftBXy0o+AjB6W5RQ99l/hgORyzZ3gEP6q1mQ
SG+9quGTTiRQQEHy3Sg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GxP7neU6pelOGsRYeMpWhq9H64emJJW3ch5ZqO94Ja0S7m2rL3jKbNa/UebfsafxW/Jq07+9ZHQH
nakVk5fs+waKW7fPdCvasFZq3bHVoH2M3uf0FMGIXnsyGlgHQ4qCnawBWxPqrfn3SKY260XmNThN
PHkcyDSRI2OjZKzXzE7AHiKXBnUYqYuy5pZkIRpG5KuuXSL3l68wM2qwWAk4Dy7OFak+VRDwWWle
Ve26y55BBWyX0cVH+A1y9sHRRFBM6x678gQjaKYO8u10cSkLQEatg4BKcHaSLpXozsPkT0ktveBN
etZKKhExPa6BnJyzgqh9xypSTFtCXtbhEF1Eag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22208)
`protect data_block
6YhhpUJPrLNmcn+YLZZPKKUtJ275GfiEr8IdZCls1kxvvjTO7Z2oOlH198DYOx6T8xzw0I0kEVS8
M8cyDTzoQ/ZEMkxfXZ9iwlPV8rXXS0PDr7pCXf8EUfHBlbSmhcmxi7mXsCXPgu2RORk0+eFBDyEz
frFeoWRmp/HTlmJPLj2BUPSqznNdKqoQPy/0bZy2k+/C2nzkO9VxsOQ2smnGm+KyjsSn/I5JC13W
fIbUB2WxWc7Soze51H4Exhh7QaCCJu7eGYberTxhbqBP8Ph3PJcpjQYfRgiKg09oKoEH2XyJNDJU
2DaivcymBriNgwRrDiKsp0kjQU8MVRZwy5YQOfyWEsoHsobigOQr+1q/gH8E3AAEZI/2IUzOTxRt
EBRGEWHuuz4HxKkCLwEng22xuaANorPgQ6hiDTwyuU66wAZGkM+icV3BpvF4WOJVLq+QJzYJht98
nfGCvyKPguWPfVItTTfEefJCDJuCga4J5bo8rbnod5nlXI2cs28Dz9BI+gP3eC6z9AWJmpVNo2qW
gJbF1A6AwRPq3jdV57aHT51FC8BYemHoKz34WpOPvwwtVvOskJLiI3TFCu92JP3fqtnNdVY2i3rm
VjuDvLcVqixwTt2CWWZjL/P7BMv9ekl1aeevjspUibdg79ryy9TJYHHEAVDn61AUP4m94Z9QwVC8
zhTGyr+M7Z3UkZ8currkELvzWjFhs/FgPSdrrNDd9JcLRvNi1BsuhjM17tniHkr/LBsYoBQ+X//g
m37PhJe1mDqjwPB9sdwZdhyMVEsJdxK8XbVAFhYbHSKDtwGpKrtyzJBnbHlpzfspoPtSdJUmLfWJ
nF3Ga0nPGuC6CfhcjC0hSlEUwXcf31QdzZLudE6Hpk2t5jUSY5T9jhQWJ77n+l8ZGr7O31ByR6O3
gayR7oUhyRGfy6BE50XgSr607todUhVaZ+KsHGFtmiwYrumPNG8wuv1MNXb9yfJwohk5kT2S2/+C
V9+w1cqk61kIH9idqbjPYdUkV0baiGWMwcx4e4y7TcCOgkvhYDekyhXmbMbSBh7sBDGcNC0jNyDI
04BFV7euXOFQr2/iymmPJQcfY+s/+Nf51VI0yxqXtpwojRgr0RGYAdtGUWy4igK7x2nVmiqr3ltO
d6xJgkZYi4n8jNonXjnwaxGa7tCsAORCGslIg9L8RGt+jZQFM6bwMevjxpyvAqMbgfCeTv0asJvJ
2UD4jF/DrhZwQgIs2pCfjV6oZpnXW5HEIEvxTjx2LdNblO6qIcSYcU1kNWSDnbYFYMmsWj5uu88Z
TzbmlrBttJiN1IplGxoA0+JEDDML3xH2EDHpjq0r2Edjtyp68eMG8hy1Pn4VScu3dsbFvvj9RxAg
pRQLuS9jjVpAEFDgYOHnlmW/pJ8ryrWSAY/NxOdnvSoePUQim/iadWPpSEfZeglrcaZtNDKnDfzO
kV7bUxbJeJhcIkthl3YHMvUKr6KsbhKYf6fFmr1FWMaNSLEPyJKW2i+Ka/IgCEWbbp9/V35glMKi
WJPEml9FRBwa8gYpTR0oRkVkbZWFxZHqc9OT7WvahznEFKXM/sZheZmjGaUZue4fMmN7xWA5paO3
Qi+V8tsqagJLC43rphdyAjcvW4U9e9LMWKk+d9cwU5CqaHxEWmot83ZdLzsAjHdCEsqG7QjWKcJg
bbsTtScvYoa+XfCN+pDpde+5dUTKeZCQ1YTRKZm/4e5JJTw2AOleaNcPXTxMAm4lpoCQrYsJMekV
/hbtMYn30Myp25Oe3w8jcCy2Ik4O/YQ3C6m4SbpfgEJ/Vd49/Vblkyj9fyklJaUPDUG5fAaKRNfh
ALH0ICIGGdmm1D2fctlPKPKp7bUwwy2M8xp3b8eZDmqW+s24brkmd2qivbe/D2M4RCj0VhcmEd7Q
Gxb4jmAc04SfL7Fv7yswRdKGV4sTMjJe1inSH+VT7hqrO0IlBeYGoISHmcxrMjiEEShCF460J+UN
Vf082Zaj6eR26MmjnlajnqsBFE5j4zfypP13ttQXgBDzNFRq8E/cnE9yfhRwQCdJFB6mTsB2KVDr
ny+dsuVsN6cf7lt3OtB4TQDthtnwdJUOaL6twQ53mN+Ri9a2+V0AQsX+jAenNYDKJiwwKMHIxpu/
IfaSKFfunFNtAU4pfBQYqS3goWqTWbVmbFOmHFRPTNXTjT0b5Z17Bq+YZCET6ASPROwpJ/zfIbdK
7F2FZVyl6mqT6wHIylisjhle/oCYqVb4ttyOQ6UlCdUTOvqRXzS3ZTYvWUoKbtRH8bfBUFoyk6z/
gUnm45Fv7JrHSbromQNVz4Op0oOgLjOuy3rLxqVC7eJtn+5JM0xV+m/gf1K7X0l9JcvsgxWyvW5I
+M6lbuSdA/oTnAukGoaviplx3mcj5nkUpVsGoTEroFU0kXKNmy4Yeuqm3reoV36Z/jolLC5qYd5W
8M0SypaaX9roZa6JfVEHXW4rmn1sBwfwEXV2jTeeUYODewXztULg++5MPAE78QTSI3kBPO3u7GOS
kuBxek28xQZy5yV6ahTaBNF7sBtOPRl2U03MW/44sfdorToKuXDF6B6S+D0kZzZThC54Ix2oyzcZ
UC5XYq2RSJc8uWkpeH1g6txG4kp+12G+7NFsaqAgryH6mAv3HIyJq+cTtV/T+8jtOkojtFtwacdR
yAoxNfXa4AUtpw3MkoqAToN9L6II5UHqInpldUcc6lv3r1UmKFLZg4Pvv7iwGRN0XTLB5AW98v27
OaCzgKRw0GarTJ71SOHs21gPEpMwp+yVzgR9EhKcZ1i8zK7vtN50Tv78ZTpYxgIHSlMuaMAGxBET
m2fh+S+7sst/YIJ0zvyUCWPeoZzI9P/B1Qrt1Xn9HrXZ+CJVUxEqufgfHZXy9X31PIzrofxdPJBw
mik/0pIJuan2Ljs9wpzOnrXaSCLtTZFA5wOo4ONgPKHgp4g30T6XRe64wM3hVuGOuQd2tZCSS1OV
lAKbLaaJKpNsp3XmHNbEN7qpcDCkHO4WQyjWIAjar3Hor8iuR3oGf0yZI+EypgJDGxqg9Z+XO5wA
h7jQ5/moaPVd/phhuduqEugPC1E8xvFXXoEGRUIZpScS4BlYGRoPuOsZidcMY6+CZqnzv5ee8dYJ
P3Ms52Ra7AKEFlbMqpgjnyD2wZ7IoTJ4WnhiRxs5Zp/YTFUehtUhKxfYEciQyA0EVW77BWkTOier
SUNS4aSHGAdJJ02md4IzZZdwA7mmGHoeejXYXN33Zh11y9HM2+c3Gy5/csjyqsI+N8fmzJqXm4AX
GmPaaYKHwBE2ZY+Gzj30JFGagUIX/ug/PC70KCKSBiT6+E+fdnN78Uri3M671x1+r4s/nFYbO6eq
IDjMuOdfz9vAfePnTrknZkf1VrGSPEC0MHDLvbmRFw0vnHmBsJnhhZA4ycpUac4bbWfAfG8mE3hp
Imd6NQ8lcyH0VCyP0sg/m2e1YGsXS9t6EJWqW82pJlxReo2qFtURvLXeMGJoCWucMjEhh6L0sx2I
dunHo+n+uPXVp/cXQKlQ35y9LSsCLT1uxUpW2Mc+KSp0azYiDwtXftehOZR/CvZHXy4euXeRjAWX
N8PaF0MHpfQlXY1RSEe0GNPQ4CZ9pJh4O+5EXu7EJ5q3Cb7dS5Q7tF93v6s8NYQ6/sGFyE2W4GqZ
/ewyO3mfgO/BuhhD1oDbEMwaQrNG2OPVD36ncGjGYpgxUk6dQFFP+L4rUWR6XtH8q3xQHg9GoTNt
JWQRXFfifz/2RBIX8huHn4DJpckPBtjCMfCOmCo3EniZyiy5xKYsV+yOiHnc0j4wY7TuexSMvQ65
vemgw19TmocXKVkziShhDPh14cQ32pZUtmvf0x7AJoMZzKZEs6MqiHZOxxGa9lPObbOpDPk4Qin0
3zmL54Yp6evMCXXgbYvscLqrjr5wLZyvyDkWaWd3JgTS9xd0tLlZREeEsA1yf/io9yPQI8ZY+hei
AZ9lPYARZv0XjzAeg//oTLsmFCBldwES2nx3VVt2jrz5/ak13xP4LJqhJOYsCDHeGK6lCzR/FXmC
TFRMXPtuoFhZhSAbLgYPSCi0+rx5FvLHtELNnETVskSUJ/S9TQrzijGADGFp9oK9jFXSvYD2iIHe
lV6e3bfCZgtk6Bkj8e8R03BHg1YcIHx0SfRi8jGwDywXnyYwnnZ2g45hv/+BV/jORXeSv3wxitUV
WAfv3Fd4ZHs/lKtGQXHSnZ9+LdWDm0Yhl1nt48dovjLTmtwTg7ay6UrMJgIIRoTYeCdXbFK6YfTg
/CIe9kF0EaDipy4ba5GVRTJN+I++Ow8G17aGmTDYKeRPXK30/e0UIljnhtria3bqDLG0b315+4gv
R2Wd75iw2igTRMM+QkRystc4/EBoG3njeD+PAWFq73nmZ+W1xFZ+R9vDI69DF960NhvRy6r869Ur
M6gsd7bFXBkZU3UBEG69NdSzSaEKA/Vs5m0X72jDTfFnABRbktEkOjhHxGcMQEAKKzHl9WcVsfOL
AMnF9d6bg0ujAQLMDS4jmnfTSos8W8KYM0X4+PmDVcUWWJ2pjnbTo/KxX0by7kKK1zkgLT3Q4y1k
RowiboLO+S/d+iYE90aW8/zg7/ya/wEoQRQZDwQR3CHwoPTg4V9Rhub9HF1cpwjbhUM/IovmukeV
fBG+5GECEr/oJoDaHsACHTaR+u/8rIpNAt+ifBZvc/BM49wswyhn1p5qyiaaRwGl5+zVOcW2/o6d
TJMVlVwrtDyK5D8TkJiuxmMYR+qCN+CmxfxKKXQAf4glFBJ9G43YNCGuCg4tpKcSeJPEj9P2u3UB
asvbcAuQv1Z0u4FwEqoBTWKIHurtJ2NgxI6/vQFpRSpscBlHXCh1VmRUBBQBBZd6hMtsn0a74BTh
c2lAoIpwwlXZRFTOba62ucTCe75GJz5YLB7fk5bcoawxr4LIqlZVPqIDUClbKD0BaLWzxkG8tiQb
C4pjE7J1CYAoBXKVVix9Hz1MvV2yvG1CefAuD0mUHcTOgvAqHmgAsxQOztyCDWTvRrVM/z/j42v5
2yvzMO7NoatMw/r7IWrIYANTHD2rntFL6+J1iCwxsAF8qnbV/B2HVtJs6f7VaSoULfx/LZjYTOK2
du+BN3yS9KAXYAspW9jyB5w5S5qD4vFK6cpHXoUFELKN3f5UO3r+eEjWqzjlLyBL0e3CNFUrWPXj
v6U7lKEkhvlYRQQq7rKskGcUp/0sRHhLdidyjWzyGuYft5WAKnKysvbOGd2x3LSkqVZ/77Sz5Ul8
/z8RKa1zAKObJz17x5zD+v3iTH6iwuxEa+kURPaWe2d2BeGMOVYCSetEvm0Ff8mMRIo9/rnyXRmn
vpjDOj25wJoFAp3idabjmM67sRgpwFSYcQGwx7iuCN3xszhBrQe5Ivd8z7v0AbVPFLJQMNmQGTcn
GiPZiGXl9PksmevARwtnYdK/8BVpXyvGq5qHmuqiQt3wMR9xAMxJhTVIn2GEbAGQFi8cUiqLy/B5
5xSx8GYVvpaWJpnjkBZNHyBZQUZle2YDaRhrYQL4PLp2tG18J51yCEL+Lens3i2UGdr9RZVhUGMF
QaxOLvo8kbsmmaClJo2mqlXNWWa776EEmhir5Sb4zilAtYOy7ebbTT0QHFg+grhaYShSTcCImyBV
/W5/Uo3inkZBjuk1FFBYEdeYiAIEn41ykyp0B98Ca4jAhQqx2SfAds27XzmlcE8bnNoGH7Ly7fL6
yt1LEti8UhlmYL/56AWgMzC5Xd2vCFtZPqvnQDJ+bvWHD+MmXyBeMSuM+WdXej9tVbLFSGMuWtME
Ape8A7kPXqdcxVXeycLg20noIJBw9E4vOpguEZAsN8JIY26j97GjBpIY4GwmzKtiPw3NAh+EiV8E
B9CHAR1KIMfuF4ebZkfAXdRDU7h2yoliRE/HNZ9d2DW2c7QgCX9YLpiNm9T7SYtXMvTRUKQi7eLn
lCyhrZIiONzM4hWoT1p0hK6LGzHwzcXtkCH91ow7r6tABi1avYtIxiaP38HlLYb1frBEFJQ+3vVw
W1F0afTqNRnvZSUdLW7Q7YlZjP1yrZMGW0plzP9AoCtqS4NKCrjJrVH1leRGDhe1c4QaTVH+346/
I/PIss5Da2EkDrVYE9DsE00ro4l2hWovj3n72Hy4bI5yyFJMbU3twJV2H291NaDhiCHnvYaj3I05
zLn9BLXTWv1dXXyOptYDBBNRWCpg5DU2T0p0/+zdN4B9v4YRRcm56GwzrfKnWr7sMKvHxhjzr/Kz
VdbgRrtH4umjM8ewL9EB9174O7w8TwMjpp2Vz5OL5xpWyE7o80rBAaiuqSHIVpEoziZYfLyI515n
cM/Jq/hl2if8LoDiEZquhUstDHA1IPwdbyt50pT86kELNbEro4ucHstY5bgGhxbsVma3hIuXwdyN
tpNDCZ+dtCqeBoqki14oVYoPir5/UxhPHu/EJl1OL5tEyWyYGDN1diwyOZ1JmPrFSO3Wsh/PM+rc
8lqHyOQPeYrLackeqGjrngdLPuI8miJj09rU7YDIwXckoeaOF34ehhysE9IuNZej7ygH8TftF3PV
SsgiSvTVfKdfsxkAoqzXDGRKORclYGk3p7Co5wTN5+PGyGRm9Nm4M2B/zJdlX77k4AaSWQ/HcGgC
ntKdvJwjbzpl8GIWkSnSA/XDbA0iHzpt7x2tGer+5AFTaSpG5AWBzgEHQh3PEUqUZ64a8x4+EVUr
iDh+MC6yiAZDhX9Mkm2ty9pdc4RevwY+dJnmR4Dd1ZhJ/7x4BkIi3rbpfI6C0g60iXXoimgbx+G1
fKqHMvxL1h/6dZwIE8AtU6OlLI/clOG6inVgAFmpsyAF16SuDRcWh695kw3zvzo4GJsq+5fzrcZ4
cJHNfRpxOYhFF/oA403xn1sZqycwsZgDpj74Z1X3FYxreweC2JaXLu0m014FVdUNQRKF2dni57UZ
dOdiW3+1+j/p+LAKZsM/MK9k1d2xlCfG0SdYBHBlu0YqhQtj+SVKLftjf12CYyMZQsevCkoogjWh
LYoFROnL0T2kbOdt2P9UkQvS1LJ1pU3tTdeJFVKe4+Sg020lKJRwBVmUyqsIzCprWIioCXFFkMAU
80lCG1+Icom7Z4wwouITdA9mCIHG7ZT+rOFRKrC/XkCxXzgMjqEHhNIscfmAlPmvehbsre8Pw2rJ
EaBC7FwhkIy1FKEJQ1Ae44iPrvTsl3VJQ2EQ6le4hY1rlhWTuHROjbQKA2ftC99zvAaTAXX1nQZr
koxNxTSVJnCjjshxrUqJR3x3wAHVrqoVDTUwPke3c998ExfZXwVKnnS/U2VigIcTyROMHDh7Abqd
4zQivH/fRyGh6+hvaGm546RBiV36x6eX2aK1311ByxsR6LGD1DZ0RiTPSKnHMMZvWnXkTdBPPDp0
ZGYb1y3RSReSZ0IfqesCkLJDqtNkLTsMpZ9zL/LLy9+yaYxw6H2EDdpqvRT8fg5wUPfu2k67s0ne
xthgaPEn7WcpQiIBp3OpzLBkufItfxjh3hufSZaQLRD8qnWcobksM5nnSCMLKT4OmaffrvsLHkoA
1eYf0ieP2RiJBZmN1//tlB5fo6qr+Wzum4wVLgIn4sF70Sfhg+AlIB76WDf5H7FE9/wos0kigFgu
QO8ofju0ImF8FIvVW0pfReqjwVaglOS0gL26DjvdMcUcus1TSSHdPxbwywRmwynHLNyW3JGdRbZB
1WDjF0iYQ15ISu0GjpUrxSd3RqgIbfNn4gt8lDV0+/Grg76LdgPZYB+s4ObfhxnOPg/5V10i5SBZ
j3evjkngTgmQ/z/Y5DtF7Tk027uXDLgNjJmp7IaU6QZJJN4H49Mpj8SX1ykqrLaC0B2rh9/chBTa
80YmdCo+QxpW2TiDCjrx87mc+O6CHz9ec2NZsHqTsGyNjjFchiIPckdlZYBCeA9BQPftm61PwaaF
Df7AS8R9ICFjPB7J0cPguOm47YtU3/RurZ7oMEVda61JQ3xZrwKqVUuq+dNDYXQP/xHX4kZtqDJX
wU3UcWUJ3gk8xMzwMc0WvkVESHKjNykg1scHV2LF5YySZ6RC4WGECQSW0LKvK0+ARDQCYAuFFSmy
+8hY+XxmAJufwk+j/QEsbUL2rIbkLQMkYu63dY48xB089C0mrbLv1EXNjMPKrIjlTt8xA8JRjaj1
+OcPbhYf1JSNkMsFQQ5PaFwI5t6j/d52+AjQqdYoB5iyHJzeekmPFBC+Hgl2ovCe7fFIJaJUwj4+
7TLsDScHT7kdU++JS5QjUW4OWhx3rtTJCc14f7/Tm928WKuzshqeswIH8w99/amLQ8liP6Q9kcIc
btbeMaiWgsYWxCS0EhoBiC8RaBR7lcyos5qmLmcT2Q8GcoShusGpV2v0MDJZgvaBvWr2ChHyxpoy
mf3JgEag4r3iVrxzbkVbTDiDTojc4a1H4yYl4XiFrryLJWXmlxRVBu1zxE5RYO8nzLoVnBg73pmk
kHJtyaUzWWUd1Lv5GsEvUcx8B1cClIe6O9jsinfAlKvlqdwm8pdXRUScrDa0SjV2lyuJM1STXKhF
4RQM80bSfJ3Rj7tB6hfysPUATKA+jDjiNjBk9sZznZRiffSWFSyoi8WNpcdxVMbgQuFpbGY+vXsf
cY7V3vUcC3Z53aQXBSZl0OqaztKNolQd0q2zQoQfes88QhVuGL1pvd10hH1hOnd9D6RPR/n5JgVX
Tpb6EbwImuCtflWpGl4CnTJSoecxpSKq6mR+haeaC+tGQKbfib1Gi/PWZpleiIIeqo1JQJ2dIn4a
WOS+85paC3XTd7IfvOL3vR5whQK3AC1vzuVcPxuEHRZP63AyUOKW/G1S258zJwXvTNNgb8TNXzVq
1GJk1cs6Dqr8S895J/291M0UQZNqTKl9z8E3IT2G1mZv8VA+F+72hvWDIm6/D81FaNOFJN4FCzia
J7KnLLEgSMArWCqutFeK+U1n0g00qlP9T0RaBPSTaVVDI5Vo5j7aDDOze07SAudEqpSTiLwIZfps
AFLMrpgJ8El4l/99jwsh9vsS2D5r3bBfJIEPIoRFYDz4JZNZs+8zOupjl1bpOdH57qodQDGv42Pr
4V9mYMNK8lyRSt2IxbN9Sk1ViKTlRpoAUtGvMOKvVM6SuykMz+VdyOt6uae9uIoMgej58RZjuDx3
UB1/I2wt7t2k4uV5rXl2g2s5R1hL2sBEncBMmW+On4CbEBs2Rx1XswK5sD7/UE5tqxFJOWUDuav9
+5Jy3gkz8IDM+NqY6zqupj7lwFBDWLI/li/JJDrAraj2tl7iUztNbyLrAtRmuBjXHR6eh0TCDb1b
aK/RAjZENzRmmCiAEZD0LZvbb9DjHSBPYf7eiQ2ovAyV67NqQ02lb5z4iAQ7Qy+EZ39ntzpa3Nko
2H89sXOExZlvKNdMT6c/rg13EaK6V4GMnhMMa9ArUSR5wbwLcvuxnXKTegUd/8f3CY+hXnyFUq7F
n4Sslmx6ZkUDTIa9/VgvV0KbeNJMfJfDTt2wJ6meYqELlIfcnvF5gDK+E1XNu/XF0NcJJ6cHefRq
FtfAbyfPcguzOouXcTM6umL5FQE70Zbe+l8A92e6DneVLO2eBUlTjqPKjWLj89XBJ5QtJgO5INUp
NtjBjL7jthKQ2m/udTFF/1wlHyU/FgViwfZfbncskC0WZDafdQpTpOuSNLJw23E7/ae3CPV+N1wQ
IjnnwaHC6b8PZ2MDobZSnG+Gc4y9/RjK0aoe0AJVNBDt9UABmFFLup9PrvOXaMxOCuXX77YWBc9y
9sgywFPUFnxwFTSnsJSWF8gNL39Yfm0VdIDRtmrcjZEHFq8MWhs2wj7RWC94oSyzua5dcgY0hCpp
T4v5/qzWoyXcCFSJvTfLlWn53C6Pn/lzbaQ58q8GNvJMXD4Ruo1Fp5+5E3xL2dnkDM76iDJ1RXjj
d7ga0UKGdKeFOLa+J37QH94z/F8QNhd9TicuAIZOTwazbtc+XCECe5EFyaGVCLW8mviZkglfSqJq
lq9mjKYFcWIMY9jyNBeFWYdSUqhEW6bXcs3FA43DS3m5cX1vLY8TXAoLuV4JkaX/ATLR533i/vOn
MeEBHaeswARXSZ5teWd5np+ABfRFC4EGrtlx1o9YChKUQyj3NaKP/UYJ8C8W8ol68c5sgYqODUMA
5pNaSJvlMg8FLiUh/2Q2mEk8Xg+N3hl66+fBE7AIxrEuUhwbfTwZmq47y9vo/2SadSObJ6P/q4NA
VK2ecbYP2pwDKd2lGH8c3S52LvoVMQCW/Io9PsZHEAopySqNNSW2NCWt+vWlzKRPR9ttqUZwcm4m
krnZWY584HYbcMHj6pu51Y66LI0npUTuv8/Uj45EL8Rv21ThWU/P5V30tgEzlPLvhpDSkWtkt+PD
sNNj9AWQ9atP7S1hSxRChNpdMnPPFfaEcRIKbBaMHlBefvYywuUIzUyV0pqQUVSGtndp42OOu4I6
0k+H4WKdXqvU8Pg60nT0TZ45HDj81NKqA17HoCJGnHCBQoN47dVD+chtXSA7zECFGm3HEhxaJ89k
DmutVg0mqysfMyccLvr9JO3o1WVj0j7JS3184enJpl7MNGVnofHkVx/yt/5OqjFXH4VAwIgGcPKV
D/aese3ZEQzuXciJFd2S7bLjd/ONuSQCeSUOjfJF8IV75qWkUUcY0g92IgzEL91dJTXBQRuyiWEX
MuLvuLmWZxvb/s0ryr7yDhE6OgvmJP6f/07sKa0h4iF8Pdq/FsKKxMuX7HD7QMKbsgPFBZS4kZMa
Z31GLOFDDVC7J94TxlYLMZPiM3RNDUK7mzUNvcAbTYxFkSgohtGlwJQqG6GZ+MBuBFi2RCL0c45l
bVTbb2kB+W2E+50cY61z7RDLe62VhrX9UbMhzLjQrfGUP5P6ho06+Q75QO3Q9GPGT3nbcqbME6XU
z4STLj3+/tQqIgqo0Nh6fI/A3VV9bJUOWFtcCbDwq2kOscLaiubO+8XH6c6qbtYqiG4JxT1aR4ES
zdfVPJPS06SnTQZBF9zf5GMS4DCWjkKPE88LwTZ0oor7GF3+o82MpoAuXSLVHrEunI/ixk24gpDn
9yHHC7rCkoPzyUfJgP3Qe5p5hRA8xQsXPRj8rHXsSikGPinFWQHyryDWZOLaJOf0H1ql5yqJHa0E
RCqH1BnPRVw9X5UO/Qs1p1BM1QKHTdvyXHxpfNblGO6L8Ymx0vmS6iaJe+PAOu/CAWTeZ5Cu636P
jhbIPJck0N4DONbqGty2bNTPiwhw3b1nZorNwibba7xRV3lMa1oYK/hbDUQKVujv3ZXaE6eV0H9u
XuhNLRUfoDu1R9SqXKVVhpYSyrLyZi8wvwAIwWOAIohBVkXgGNay9BPBe4UhQ25WcMFfEhQOpv74
AiHe88e0Ll9sqxwE+PNCNt613WxxCmH+arluv2+WPa0p/njDnQANC8mi6/78DTaxleusMlzV1WIM
UZNFvihr31qXqAcI172scQ1e2qP4qEuIiD07wtA+c+Bu+HNseLoYonGlHZw88PGE7muSvLRHaP4O
MuC9EcSZIz2VFOlskLd2WA+mdQEQW40U/d2h9DfHZBfeK6f0HUr2C/c6PBpIxKTuK4IgWTdZdlmh
8Iru/TtpAshSJ69Drryp/rQt8VabhYr8s4+1bHkgi2c1OghtsbuvgBlBYS+aDTU94cbq9Zv/Nh3D
Y85xXr4s5XZYlmGwolgE2oiQPPFFkqFve5mzEEcCUOaoWOG4A28GjHpzo2+RnBMUOe67ykSYv0SK
66o45/l3j8dViBQ4tSYAFW9j0OVdZWGxzGTG2hYRIs3o85g3paeb2ZzpTV9MFEHbYFtnAxrmpVmX
frUIyZOZmBOAiKin/SGmm8jFcBMBCf3rYsqIjBz0KTbQUcVuSAOKjgUyID074cZLRy4xeM01EIA8
86xOhUA+iq8TJkv+SDUCvkaVGDg7ttVq6hqAGDK8TpErjKeSM7KAjOhsEg3kyqRbNbw0he+U6/R+
GJIBFIq5x0ayBt6GXjufSvB7ofJ/YxebIxWVI9onn2KZ7UMXKIg5A+tvFENOMFSPdK0JV9nxzjnH
zSGk++G1F2HTvSsBspoZE1NiguIFwKmIuUhRT2nBE6dX7vLXJFH9dDRHK2uDnvD9ijGDzig9mmrq
CJiHLvlcXt65+52Q5CL7ymg1XZhP04MrqcPll8rJGh06fgR0pGOhLuHwRXC7Y8i7hVqKfJlltthO
C+gOBkZYBKJeFaxB3TcgiFyPer/kvO6kDpRjM+d0E5dcuAWAvtPz9MrDWRT34ZVdZkx1fBCTcbaW
peq9VVLDSsODqSzig/SISYH7HFhK1qo/64UmBSzkNVgprBTWKQza34cyQdwS6TE3NDg3iP+kda7Z
lg5NQBLkiFgLyfQ/nRWEMVS1S/O5RUufo8zyAM7iMhXJMgjmR/QZTBqmLr/Hy+rEw+nyWrS+bbs+
N9jMgLWirS9AWHuKjDjQD/6pLkowvV/0uffKbAL8Pie2ka6YFKKQvTkIyPRMo2Xcemf75Y70ikn7
TY3/7KiyfyYc6P6gRhLXsAqWP2jbLwdNwlaaO9c+mA7dJNTJMZRztpvUhnEDJ7mqPNoLEYo5Vh08
wiE0cnuF70FVSCiweuiBxjaJTde+fPT59rlmQ+isWXIl5nx4zAHYz+McdUUroKxz7AzUmG92A00z
SjDXYKv/juMeMgr1wmi0Om1oDj9nJ3jkPdYVNCY427vmRoWiabJJagZYp3MvzeCvEa5zYpaUNMcJ
LJsUNMq4TqPOPsUOGUSRtev4KxYJlcqPo8IiV/amtqZH99sxnZL9imwrBBCxrX6iISEyWZiPdvXP
ib7ZncIS5uFKPkqVFbgjMXj9z9YReGzsmeB6dnbLI3/hvnybogHZXO1qp7oySmwq+3fw3a3tZtqp
f8oa+4xa8xMXMyAXQkgdbG/Enxthw+T6y+dSV4STPebE5vrLpBjCRf8XAR69FRRouJlbLr3Sig65
X2dPQh6x3fKJxV6Cz1QCmunww7KS7E2OOqIVETD2G9jya2iNtmLrz0clmoqLEK2tfD+OcjI32+XZ
RlexviOh+fvfqNqj3txzCjSefObzs3PHbiJme3DgGPcbyQChJ97ThXz9TiPDLPllNaPuKpDf+xfZ
iuiBpXovMngWKjSaREzjkU/cBTTiGJhIHPxpEx7YWkphkodDduGHB2SVpDsnv2vs2zKH7wegouoF
9XWe+OEC3FhJ21XR9ZuOG4Y86igI/g+jW4OrQypWcThdg7eYdTT16RyMNKg+9nyW9ndJfGpnWJ1Y
73ALwccC5FfbmkFNlYoMw410BFAeU5QFHXIDG3/YN4hUU8HpXh4icNHyOPPg1PyGsNBfHt0CkM0/
aMSd4RrktqXdsZDKCnWIl8w7A8YhGUDOyJChqC79EVGR0VnL7iqh2/8F/CHx/8Z0CjKiWf9osNV3
OlLvFWC1gjDB23YEOl5cU/ybmceKiTvLOn294uYEPXJoVSSHmc6xGbKwEVYVT6NxtqCtQHM/QGYW
RDGJNvpg/Ihsl+/P2z7wW4DoAXf6UuvQoa/Cy8ToLCttddqVQGjDEflw04ES6ZqIQWzUiJjVws+c
dMrNCB0iMDDiTVtugT+qldS9UdLlP0GeE06EDc5a3n7qCmyH2FF1Lr7OqtHCxuElZn3VJ5X3Wv2X
6ThOgPre4ZBXijegzL9V1GMypH6hMNEUM2bRg4VRgN3pYY72y/evn1+BJ4BAzvACrE+RyDHfWR4z
32g6I5rpd2TIcph55Uik+3Oftp/wU5Sb77gh3fRkwLXlLWU8AzhEnr/scrhYhPE7380LU+E06bLZ
VMIvTAMRVAr8qsa9+ySK6ZotFB/cClorEmydzWFY6Q9gXDAzlEzNGcye+Krs1LOuuYM1vFz5jZhz
iHgAGHkth4XPYILL0YrEHlZE49ND3SDJHyONbeGTx9tvM0cO18cIv/NuDVnROYwVu8iyIfQCu7AP
9UIBb8a+uCP3cguON/Kgtc3u/4ZMSOXWbmdkd+I5ESsDuPviVP/6mxLa1oLyTA9sE306eATiT2l3
q2xbNmvJe9EdbH6nk/0lox/E12IpdzG5DsrdkiS5XvHhNfmRjcTJ1MKqnBdpZVMixqpSJYyBPRQV
VKhlpE94vcuLQgUSynM1hAa91S7yYoo7N8BXpDJZo/cWf11DsopGDP+62/KrvtEUIS/RBGgXMEeB
oC0Cq64xqf8b2fq/B+LBVuip6Azn92f/y+PflS3z5Cx9jbTJP/DX8fmhF5f1AIQDfXoQXrvUjh/J
GLWWU8E2qeFM9SddjofdXG1fAa4wjIimN1adznovsD/hgPwFkiegoExiHKodlTjFs4Ofy7A+gCZ6
N0qy5jeiGhv/ihf2VMKuhSselY0D4tMNeMci7FZUgE4VN3vPMK0HtQHEdcD31tgU/GFw+Cwk52r+
c1UTnN/RANzV6xkod/zNyZlaj8PbWiDA+eHSzE7hDp70UBI5UeR23/oUKcQeEjSCWDHBZ7V2ltsO
y19NbroeiPYjwOYsJ0SLjRP51IOMvDT2+ZTAHST5nHejwxbp2ucsFuLeNOhwUKk9RaqF5fUchzjf
iDaoGo0wyku4qmk+QBsFCLhre0wKTeZ0O7MB5TKPK68xRhQE8RDfGsHED1n5WtC/TqCxgQr39ftu
1qG9ItLjWSmgh/VjEcr+8hd2Vea4FMpBJIhOWuecVMCagl6nb9CZ1wT34avQWhpMug8TcQmEXMUC
fB+PIQpBUS7DocHsNSeVf7zTpC6hYXPV3+Rz46c5AD7CGlgW0IEuXkC4SBPmaI7cwqp3aw8RYbaD
IJSMkIfoVtGIA9/kOM+Pgme4bEfGo/X7xQ+tS+9Z2SxzFyqAQfce1Z0HCldjlxdFNkbU0RLvn52X
WECFIDQp3ASmQX5mGom75Ir8fxHvCSI4ONVGOqlj9zflegzfF6xo1bF+C3KKWgvYtRyS+3BwFeXU
kQVCXk0l+pmHvt3ahC/Mpjc3Yofw0OTeCO4RCYwTDqcs36W1kNVgq92JqXxSpVvuZn7R4mNbF6N8
NAwIr43bifARXy3DMPw2zdeFuk3qlYjG5dGHoqA9SzkkBpvfFyiDzR1HWDCQYlHZ3jgQKIgX9fr+
6kCkI56rjm04l1eOdmHL7wAnZUSgAXZhgVGmY5S5t3ygVduQcq/h7gyRx36Yp+w7m2d3M9Zbw94D
j7gXKqghMU7565k6cNulm43cBw9WIdMw78ICLysWeyK9JzyRP8Rt6qE2hewsU0oaKAfQCW7LByLj
wRCLWiMBRjyrpJURjy+wDnjFQ2HleEKTMO3eVU/gyWFYPWVGa5mMfZYXJ0EEi2sJFY9sVsAe/Ycp
jyvDiRmaY1wCDBjSn7oeurNId8VqAhVbAEAJUAfnkwS23pfFInztgzGMivCd7/QOinOZwoLVhLrM
oc55GqPaefBlzotYjVqs2M2trYQU3sh9ABdKkoEmwZpkEBZbr1x1Nlqr3tPoLFxn9JMTvY9frmXF
55knTzi120mxatxXTLZ/PPWB5LJOVGvgvQISvufMxbP+FXR6N1U+f7I/QusGjjqVQ+mGjVyaT3YZ
ENmp9rze49JLfBzyyRnKXCHQVLhclq8mWlipoDzk3hDpVcFUBJz76FMqZRZqTVuCnN8RjWx1Tzd7
qjzFhdnX9fHf+qcZ9SsEeGy3Pm8o3u/QJgwxFEiikpuddx+sroYAbeF9nT/GmZ+1MjyVVRLkVVC8
zP6qPeKvHz7WsdZMezpZwXptSjJx7gAC4xZiOEgLyu5wkQTEYmp5w0j8RxS1hD2FFtn2rl6kgxqS
5V2z0IBcF5aRNVt8Um8bQniUlSAgd5dC0RxrX2saGwIs2xUWZHbc1FLYAlqa5vK16Pr7RWzSe3QT
FJQT1SWd4cLNKj4PpQeWSPVmcD0mBUQRFFPM1IyHNydZ305NPl03/+BPusAjdQRuYCm8myJT7KGq
SO09fBfO3r2bCEYVyeWC0CbAtMgYVAVSRb8Vv16RW7VpgHDnLUCGDMO2MuQ7hpN4JR9l9PHWqsL+
xW8AfIKGmrPnAOcDity1rj75fdjwDv5Ws0UNBcidpOZI1ymJrk/72yMnu3ruwKDRJyOJGejDuES6
TLN7i/TfkZ73atc4mhp+NV+nIvpdwPp8n+puKUpPDBxjTeE8DL8SlcNKleyUDwqw9HNQ/g22J93o
3wi4PA/9/eL6RbFgpqwsbmy/61Zu31BqbYG0ShofrfAdGnXdhSp78ORUyz86YbuAbJu0820nJBBA
POIfMlTc8wwd9V+bIGm3OnSmF3hZhvtOtYQhi1A6yOgtZR9F9e2YqLz5nwUDEQ6Su93y4YlzSuOs
M/DbIpOZi4pvxEd3rn5BdlcOcArhwh5O2s4fI58NIjM5TiegCzNchfTmOmSQ7rtFSVSTuPREDnxn
+7Tu05T1n2+vQYY0asxRHsWKuo0beoSZ1tJ/XY6I4fHxuYfEHrmb6oe8Tm4dVK/olekXfwYux+pa
6PUVuawDd7i64YnVI6/7YeC/7IKC2ZYhHgwYCXXkMFekDCJkg7n6Mwn2ocfYzlVHMyDy0NtLiuw4
+2FZ7+K8nj2diQSfKQNTrIF8PStjhV09JiZRzpnS+feE6sScTTbvNqohD8Crg2Z08h9Q95cE/CYn
iZKL+rCZmGSBIPYmuxLOiFxSe1Z+CPwOGzFfmg7yuTL2PipmtCQk0zC294x+BfG+w5MUBSolhSdd
VMDGYLAj8TiSRwfBQmCFC9ecKjDOks4vkj0RtxDz5tLYqRBjsNulUtiEpqb8Qn+XivRKSouL4F9Z
RO51Evueylmnlb7Q5jqKWZ+3sXbYUOFYt6JWRUiq2MwXmJ3aTDrC4tW5bkbsZy14mIa7oNlJ4FMl
HXnPtado6MXzuX2bLgQ9WKDDNsqAVM9wl3RGXXm0QU3CHCB3nMp64y5SEv2ze1wwBo/lq7TkWLKr
2EE6clA+vDb+K8Iqq9Ki+a+4Mw1O+2YxiQcGsQ4fgHQcQIgBn34IxbsA0F/5DEFYqlTXYwC+YQHm
2ThuHc2lUUf/a25T32JIoPddW57uBGrkbK0p8KJvMWTdSzq2HJwVS4ypD6ntSHAIfIp/Sz6HeXuf
7dxX/mjzedvj5VlMUJ4H4AXm352I92lwzCc2OaEdLYvG7P2nnYjJ1ALpOa/qhOpzs+SFynMukvCX
C593OVVOesYQy2XbsRXdRrM5YAmRXwM4LuoE60KDsBTxQQVyqs73gHb890o3Qk2POtXAxOsLDd0z
y+HQs3SG9W7weCOdN8RD/fY9I8T8Lr5DCQBU73P3iVdHZRSMXBOkEcbGjP6jOGdoh6KxhctVgTvt
7tnEMfnFX9ufTWkxPFVl7SdyhigzbuXHiTcQx9/MBVdEKeZmF+vltADUrhNERxSaLvNJF91JCmuk
DtDxOwlWbkMaG0na8cUqEAZqa96mzureKR4Xln4Z0b45JK3JLS4HkOACyrkjSN7XpEunEKWeWVsJ
5tLlQZOTI5NyXzSgDuYvuGg/3eTVoU+Elv/IiI7FwzrPAvvH1QPpyX/++7dpaIcpJqqL4lK+M9hb
0gt6yKjl5unHcCJB+IUIwHqDXc8MDTNvLMyPjoNe88o35kmfz3V1BAEPZ9XVzb48auQRzdcZWZJp
GOgUlVwLEwUcFJ56HbGPnAug/GxBADHcYAqZKvOCasmQiUsKOoLEYEv/oopX3B5T6ZmJSNR1O6rO
bbefpcdrl4SI4RqrkdnA+2xAnwzhZbMiWbbgBWwHfj70SRuzDAuyniF6od1v4ByFp9uECL9QQFiy
EZ4kxtJwLxNBQfcB4vAnpXcWGsHMt7B3NZXJ29PEVsn2x1xz5/tjGHnWSbs+F0FJC5VAiYZBoo90
fmgjGdt/jD1yNIY1up+qJ88P7k8msJBKU2PbLJmj6/OJRCPAoNFok7JgHmKQ/d+Y9r1F4wNZY3DY
M7mncdSZPF/ivZiGnQ4nrrGWspqHVHjYWDg6WRVPzDW6aUp+BWf0p+7iq8R8QaQPQozN+ciPyLQa
F9xbMYlSqQ3eci85y6LBPyQMcHz36AZlEBVCHBli1EyNO/pHygSKeGB0NSMNkn/iB+ijeNh0vCPZ
P3pPxP9mE4HDQpz5MLoFIsfi1xECvMBLLHSkpNcUMGIw/+yYl1Wo7jtret6XECauAo53dr9uv9DC
7anA22l/49Ls4ynlSjGwUy9ynoTbXpl8ReVh7kNpSW8bCfcRb2DtlIyeOAD6TWu7LaGDpAYXFAZD
PJV/X7ai/fOvqc82ZLWRwk5IOdiQ3QFt4zSmtT7CJx8ytM4u+QWntiEryFiCAZ9ekTWP6FIUCAtn
UkhcNBnARO6Z7UPEV9ebAELsrhmgAtUOoP7SV4j/eigcc1Umh24ukk98HUN8ZOvLr2F2jpzlSRHx
0v0NLPv22SgB2U4iwB05LJQ6JIpT1S8nlpwGF23cqkTTkebMBhq4E3gbjdtYzOXDE97KpRz68p0y
DgUHgmnWq4Zmgce0eIbLrRtkj28VlyTOhUS/rCxHsaPiWRJZ2tRHZ84m2AERZ0TvODmyCRRFUH0P
cF62dqu3RKX3x65TmoTKjsGasyKFhNfA5807TnF8ohF/SYVQh9RV4BFk2GMT99+H+L1/V2I9xpmy
dXhKSas6eEKQ7OivPda6K+C9qsxJ88R7lP5WLzkIR/jGKls2D1MpDQh6rVX+ro3hJrnlFhMkq2Fz
m5ZWULFe+pRsgKcocszEOOvi/Ht07ARb8/0tD9CTCEwkmLtVnaenu6mWPwqw0bVzN6lUIlJzxiwA
o49H0gML3cOCgSE8AQg9knDpNyOZmFwhw6/1fFovZzb87xBEAsl3A1eWvuSESizgXe1yJ6Cx27lZ
sMmI/H3Ju2Eehp4oziLbhcz0NT5CXS5DVQ+g9It3yAmzxvX+icSzlrYeVqWLqcXMgboZaRPqiyDp
mxLd8rl0c/M40wCapgLgj0VOsZU1/vlRqaVQneBXdwBCIR6C8seUkWwzNKpmDtTL/ixHX6LH9aRy
Tw5c0yg7AgCKVGEdoBc4JTftGFPqaBhPqsEMn6/XtIEVfAyc1tJQNB1ckjY8ZPhuD7cZi0b6t18B
YnYpUqTVv75MkC0PWhf2VKIiYFvWNYjwJQvN7Nop49B1xuKvR65WF72vIMLj8Sh3FteO2dmwy/Gf
H7J1LnGwjyKuHvmWW4YE+0WpjuXU0wGxIvcTsmvNBqm8OpT++Igcok6RmMTN5vmfQjDU9S7EvsqT
PUv8q9Z45DYVZdWmI+vHd3x733gRlx14Xjhrkc5RbfmX7gd01ak48QCAGoXb3SH8IYGEfP5szB+F
3xlxRwRmDKT5k490IUwD1IvjwGSRJoj875DN39HrhTdndl8w/zY+KzROrLEShe2o3NteMFJmlPTO
72QZ9RemZHjWHAg8EshMBotvoBY10fzynHvCiobOQ1qaJN9VfZKen9qAyfAll+DzI6LmWkbRnTjA
2dCCGSayHz66v7wT68tZ/o/4haOjuI/YYzQsBnWp3xgo/2aPvTWR95yXT7U7V877ggPc1hbB7jnA
xTVNkvMA4CCCXx0UrIMdezh3EHpHEV4sFkiIqNHxXKlv961kAWQuGxoH8uHrzzQSOpdiiLN2dYys
JHnxuppSl+TRVjJqlajKFP5EnDc0FylQIACmeH9onkUukNdMlIAQeP2A0TT8LYjPa+GRnX+0cw5Y
wOEBmGc7UGo3UH6lmCKpIYMP4m0I/5tBb5N3IsNu0JW/PZYY7BWpuSYWTl6gcIYLCsib2U1Wbt8o
VBq+CLrQTTzb/26wk+X5TESJp4NAgaa43+LeBRwATqNICeur9A0zRQTYovuShTLlXakgV4lwoDEP
8u8Hgc9HKZxzEGvs+s5nZ1Ogot6p6isXJQVVNcKH93cKE1r86w6g+AvOrdwavBNrSn/jRNI9vXiB
os18JPKOTJnq/E+OfGE8gq5S4pHM6iJmyD96X9J+RCdkYPJrJVTkGOJ++7tY6oOGWP7sUYNFEuI0
SGboB0Xjxbc7oKy1V173OQi0wy+WlyhYS0TeWTAKwbBwk2Rl5y8p6x/AR/pwjIlaisvIujgvAJ8i
ZnXuyqJHaL0GU3TaKaKiWYs2ktRdDG5DwK45bQYzTXaHGxn88+pqNwcEQGsAZ2tPu2GgBxueWryA
Uivd7SrhyjebtRcS8zYpz8+V3AP3YiQmJ+7DupIAkH/4Wd6gLuuZj5fiTTeK0E/hmZC7AwzRETiq
C3lmNadDs9HZ4z6GggsHYG4QBwSVTFXSSbUUmRXK+keOkaXZnZtSf9AC7y1l7zlsU5OiSBB+8SfX
MyoNFFm91q14PcYWiy0KLXo1RsLsfyqa2NNXXtMNOF+PKwbTS+E6RRcXkFkifk5rgaGXSwptZgMO
Til19hgUC6jl5crSHzCo8LzCCsxPX7Nb8vCHNG6ofmDcRaXYQc1gY+ZlVG8cSl+wgkrGXqpYYd9v
dQf/Koj+skWFRX+YXvkgQQkvUnfLNzaeLvq9OOrSVI1yUn6FRJEO4ivpu7Vym9F33dkELV1Jh8sW
ocPXccA77dUT1PuKRwtO8gb6H8Oq8oI87LCKl4h1siUqUja4wvEnzv02Yw9pxUVv1AoIqW6qOETc
anKKx4PdVNdJK2j9LvgzBlQ8T8ZRg2x2acDQLPr5cBgYoLfIbI4sBt41C10Frmw/tD21gKO/gFNO
KyI7rpSSBmUl6nuq3o09xRjIP9AC2aTqX4lQiG5vjVWyFBYQi13VgXuLd4cwEi720yI5JiaKeCd0
jQFGT3bKGofQM8T0Ig4gvz1nKyd0HnVa9wb9wKbCLSQBnj2BTdm7aSQayXV6yMuQM3XceojZ35UR
2lYLjVCKGsUJWJJKtJRafBlbNsZZNKeqkcMMvw+GByV3O/XSUChFITMUYzo0UlQ6zD1RkeX7biyo
jRu7CtJFz+xF8UaAeyzFIUPpvzOnNbVzTnIDaUGhF/Q2kcQvO5suKrw/L7a27tKAktLHX3nTxwMb
lKdh52vZDH6/CKEO8iDjH4aaCFzmTBkO4TsSO4fXOuCjMPha/m88ZADPPN4aSBXsp6PiRPQgV+nP
LhpVYJ/rVVLvVFLI/vfZ7og5GnYp62qA4wMW8jxHmXsS/4T+lmh8seYcyPTgwuX8VHflGG2Ds2qQ
ag01+I/p7jhVuQisH23tg5BP/Mq73QixOvKwnryuDiDvSe9Ie8zQ7fa3CgNLWWuuMiUU0kOa6a8W
CDKHybfHw/3Hm3AAQ+4qSqOSWe+adQvDtKNm/3vbuGuSRKl9aPgnR3wlHyhKI8IiHrog6ukkBh82
wN4HseQ0i0eKFnmvE0eFLUkqUsI7QVsr2Qv3TNTk6QyHUijdafxQuEdAYJlqyaMaOKZbHzF75h73
6zE6WC5J2of5r4XJKbO39sCk6cXZxEgGhyNPhuuSv0xKD3uozj7PIX2KBy2fi4TLMgxvxqNeLTAG
f8kCri2wF9XMtnRY1Fequw3G3GN7dvuEk6Qv3n6gS7KfOAJIlTij3bqKLoLwqDaCI0tc2wboqtJ9
ySxCsLzcy+Kn02M6+POEi4w8veNCNGZuDDBfnSqFr+p/XxjqjdvCrKF4/MnxDJT1XcMBFUgr8ktV
f557Oa07uRjSm4plwOEsq90G3wc9taJOlt3NlIWwjrEY8fnBdbY5ac1ghqqF116MGTjj3CXHtCmC
sa592o1OKNaOPwvAN/3z50rm769rHeHu/N5D1CYG1gaIIGmidLJfZHYrS3h6AFRS3RWc/YSQw8qY
THXPMKnqsyDbJwyCdvV4QykyBX6rfDsxnEwxhbXSIeXLkKZBCgntVSiY2+qPfR5J7iWRIj3dp1Jh
VU6OLbIRg0YsQCukM37r5tqkN/iXZpUzp35kgfgBkLsFTSqIeyvI67cDMBDMKjBFinnoZc+CnNFG
D9ZxAmn/d3aWvD+5c21Rrm5axJCwvr4oK5q3kjQ4CtugvaOJQbMyxq+QIfFnzJ5fs2oCm4vBnZP1
ff3q1bEHXzxcxNwttkoAPlYNPJ4eZWuoT9POGpDRbgYRx29tXU9Hn1cK3hWPgqPEMs7pSJcfrsk6
M3pb3jTNrwEYQ1VOX/GOZ6zpXb87Ao2HhGoACcsIWe1yXn93qwBabHgjTthJRbXjI+fpdJ5wInIC
LkImeWvEMPMPgfr/YKJoQDm54+Kzi6WTrdUgUA8qgdGAj5Co9LhkjVRLy7AB196i8V1Z7JBIWc7W
PtYX4+8VSonG1zpvFPdYjmCGmT6JZU/Oy2ywoBJlBT7zDaOnpWkFWAlerJuxUA30PhDCA43sXyDw
Dj1pvUg5DZ0YX+G7f8DAjfOjvOxE1HYSFs1+moTUbqzn1fszR1qqwxDU4XuvLgk+2EdSZB2cK6F2
7GcNCzi7BIIGPIfeuClndfj85EfEM7bJPY6KywZZ82Quomsj8bZvfBrLnuXCWBGubQNvUladDpoz
zof6kLoyRd6zKsk6pJk7sBS/etH7K2HhHOLQcYyemWd2meSwCAdYvDQYb2htraUZLMha3TXrqI2g
EbBoXAjqFucwP4sAwGWxQjc4v1rmp+kaRpkdA9aCmLgBqA+ldrljJGP+PHFxV3iIU8S220eRXDac
Cj0BMXY0Krbwn79V7T8XtkLSa0v6nZFGNd2HQVdAPz91zNRyWGqiuxlBAB8Sysrv5/LVTVQfLtwa
w/71LwWE1YDx1MsSZpzGvcoRkMTP4PEjnBMp8SqkBApj6e11jQN81qK3FExc01GlNkv0G0opLYIx
jz8abGVx71I8ldQIFfmgOXloBu2teKN+10q/920mu2amMXsDQXrOVQq3x4tw4zuZ2b2otv1hELwK
tjULRPKrhBwr+mAVms3AkKeGMsP2MqKAtEr/TtfSQifFqohpe7nikJ6CFxR83r3pDvLTzVhGeMTQ
OYrCPlvbvZuGKqnE/L+w0Yrnf665+6ZaMaIqe3f9si/UViqWI76PLh2ygTOvc31JTtaJhRRQnFx4
HlL57mzB6O0c7GQwriLG/YY+ea6u0RFynDCJ0HJVwV54QSsYBJCmqQpchjJTTn8hZCie9WKLHYpz
ZiJ8K/L9cd6UYClqbiidTmBoR7w0htF8b0BLTxdSe4ls8vP1Vk/pyiVLJ2iJr7Be0SxdYx/vpfnq
GWkoijOpvwbbgaeDbwZffv1E4LdkT6J/YwRFU5Ks8MDVaf4lSYFxsXKgzIiUvYk8ULFc6Gq9lm1X
sEAJm89RP5ZJ8miBRQjzO0yXXfi/2bKlvzzZPqqBoAmYi6E/9RB76VBwsX0V/cupKIXl/h/Knrnc
DN6gIFZBBMewkJNvBvJ+m5wc2iO/F5rHlxaLtVjzID6TnZ4k8C6N8jMuQ68Zl3YJeRj48smqQsFg
dreMCHIewWAwn+GGfBmduF2410msRxJMkn9o52cvjzIkjcF6hHeEdotSbiNSNf/6oej4pVmJyQtw
du8u3dfMAPv+hxlHPG4oBaIJOck6rSxp8CkC8GBJpEeyz/Yt7IAadlx+6z0fvjw7b1CyZQRSSxDv
Ax0AFnwE5DOj6msSjl1V/wGISyEYJ4siPyzkb0DD99WlohydaopC/P4gFh7JQmGzns1ru3bXUj6X
zVt4PJZXGc42zBT45FmwgHKDZA/lhUUmjz5i/s5htFTI4KRLEuCWRKhlhQh+JWRNaOMw1amozXqz
/SlR7fthREyFgUAjQOfzE/P4DwwOBw2E13jCRCjpbivLLBmIxWpozBZ/cdsKFPgR0Z/pWjNXpTCL
Q/qrUAFZABTge9Y7tFA9DK08X33u2vtOQa6xjUntwHrStBduLsHkc9EtbPrwl9Ppw3AQZHcdFzCj
+AslAZxepxkCkWo9RLBZtJ8tTpYy35d9oJjCfRHUPLErAzYsW8oXXf3vqyKJfEEaFganuUk3Fbx+
pw/r/fAzDUmCEXjnOS7evO4IBNm2kX0uE/7yHA7mGavJd0Du+o4R4CLeT8vW/Q3xIQ/HldIVXH4g
zuLS16LiWk32nXX9d6oA3CUdx1DqqF6UhnmcOKU1NpAFkxAuvKRV74QPA0tGEsbgx/NUqwYpSKnT
t6b23t1IgAuOBTNGNOwOda/9acOxBqwMbaZ/M6UPrnKcKm6iRZYOvIC0ZFkUIcMFYm0K62Tofvqj
UTwzdjJ4VSSrG2yTCKF01mNJS2m/vIcxXz27+uz0o6Duf+cWRLMRMTHDFs7lTDn7D8nA3iJSKW6l
sAcQTR4ZThf2jcmUlxdbd8ba8hpFrS4wu6KRbMkIe3Cpn4UOkfpr4VoGleIOP72db67T+uUUF0ii
Hf7coqsbCRe1HUXdGqtzWedvJR91aaKJIqFYqEYsGt671y2UBSQmstV//G/ZCgZ4/7HUNKlgiMkZ
sFOC38A9OGyE2T0hvn4AeTyOlgUifbITjmqmS7NIytURAbg2kl52mOYIeBsprq1Bd69IIcKrewL2
fBwb2LHCkM0rxwx0BSKhTIXyKrFrLRFcAZQ4UYVtTXdH++QeitD5j6cWgcCyd3yIp9TxyMyFRAp9
jqvqgIrrMz+HmdEYX+vkGbAwVLb/hENR3i1EdVR/8Su8UiT62JUXPwML/H0rEPMxZVrZ9bfAZERl
QIYCyFGmpPrBSONd9VYCfYFM0zWWRxiP/6+uYTCj+TEvhAM+3htLB6OnGsJWP6Xh13c17J/swHJ3
Hhw+EJtOZun8umUEqIzjO3XSE7/OBbKQQCBlHshTmh40uFTZx0DCTJwE9RHf285s4cHUnFdiqVN5
WArfwKPD8Sw/LjiGO50w4M0xV+nod5zR0vQO0va1nafaGJQpmlvBWYy3XxSwQcG6RVjfJk3OQVet
O13C4oLxs6XdXsBNxcY7oFI0V8c8QtlLnVlnJlLmEe9IZh/CUe+8sNQjc692j5Sk7LFgZD14Y+lv
TSpysRpeOlUA7/tWnjL5ieJJzqJa+R0/JYHrr2P/fqS3FD9ypPFIAPx8Wl8siMjc8H4NO6mc1h3w
F44AoGnGFVDIEZvogj73ZSdU9ZqzSz+tq2lAaiLj/hYF+nEFHejstVYq4qMj44PJg0SuJt9jmY5C
j0APxYfy8yjopYA2Q93Kg/pgCFURun0F3r4xX/R1QMCKoyHdeLIe1KWI1VfJuCChzGylVssfTX3O
s8b710jpW7BifcG0WHRPaW6K2166A6vwSEtBYZUj8pwEd1F0MhErz4EuUsfXRwedLi5Y6ds7BU1b
1oyAu7OMWM03JkoUgY6+RCSpLQrPisNRwcqwFehgMEMv7frPiezVdRxzdT5YWQBWafb0XfLx0XCe
Z/Y8KJKVrGCl23z41MEOvWHgNTTQ7Z5pBBpy7rZW6vLuCoo9QIk/jrBmXaeLPkzGmyCX9XrBtPIc
wajot/4VLUteNIsPwc/Ig2XYOa+KVyAob24a/kqkgVge162U9ccdgQjuQVaviShjQqululcIZKyA
D+eKw6KUBsMMWpVifBkMmrZCGsSMOiMpyix8UuPPte30keYpD20roEV6sA01B6wCO/d6cFL/Jyqa
cSkrjJijuhr6jHRL3I0JYnZ6uio4NUZ9yj1nGOk74e8U6gpvpIPaFcTbYRFdIDfSMERTvqtAmUE2
xAGSyRmQzp9jdomofN39ZLmzjpP5FUBGUYBDNZYnSFPq0ZRyN82zdhWiKKc6Ze5ePwgfKUd+SqXM
r2kobKBcFLC/4ObAUKFvFvS9k7iYqNYDE5HtwYg0eK3mMpciR0LlEMD8uS6M5BXKiKydXLuXTZy+
Y7MA7n15HKh6G9cllhOdHNDfAk4h5cmX/tRDxFGNIW6KIvHktMoxopcoPdkl4OXNRmo2GqSjLe+7
VX+edAJSYlj5+y82xHbFNpiF8+K9ny9xicJKvtXHow96+H/iaAmW7Fot6KRzcriwLG4zbxDkdx3L
9KhhWArSiknkQtlBfNOrxaVsT2ZJ11i19W8hoCOPvUulZ13qVKGJsXw17D7qI8COVgX8y539ePAK
lhntd/+a3e0ITPWE8elTBqNynU4nBrbi8h/NX/aZs4JvjQ1fukqt+SifpT1DjXfajHzti7vtJleg
UNrZT4H4aUR51Bt+s776tZW3gDZqNfdhKSAeUBCWGF+U2x345g/ZrfCeTmgKVZLKZUS00eV/QlsA
sATRU+9OARxxI5DS/I0Pauq8idJZqmnjdFwelE+psfanmVZZ2h1u9kaRler4bfCXbxW0YR5zzHW9
EY1S3OVbNzj4HzSirn+1LTxQWddUWRdcUqyT8ThBOb2703IYsEyNsWGVuh94HhmzxyBLvgrUauyB
z92JpI/O8SSP5FCeE/6RFneJRbzTSHO7VmhB4icUOdB1/skFZH39cUzvylTFH0YgpRh5mqnK8xhi
6E5+eaDWSCiYF5dYKUCihMOBLJAQI9wbsEmn0UIod2yHfhetNdhDfKmy8DeHdM70HnHLUVgUoUsh
T0XZMufRd8ma8gmJq8zTI2ZqxQy3KB6J0CKQav8029p8zczcGSaB7F31GnH7pAYQr9HI5MlEK5YQ
uE2C5gYjN7I1yw9INbAdHL8L/3yAG4Wv4bw0HfVzKnfmr8nHVsfJV6oJCvh5KltCknBAUCjC9qS1
P8WIP/QyibLPDy7kH3/fBYTMiTOZT1EZX7DnK3UB96jtnK/6beGRblUJRWRbWNxLnTu/KAwtu4Eq
6kvrNV7N0VGsYy2Ik0xg6lOVKmKsoEkHzF2gzLRmmozF78sxv/sgRMfDOKZZaI+2caAJ4Mu7byRs
ayDftJvbNgVk/d6jNTV7fNFxRR3q6iycirYO2n1AjRxtTn+7zoyR8+8ABGN/m/nIVeNvxucKOoLZ
wKkjwBWjpolegyVMIc8EkXu8Pu5ilu1KuQ4lbvCGOYjDRKCA/O5WKHV4wTXDS+A+yGdmNuv3lpcl
P7fCnw6W3je5ie3/ADyORWfK138q3e42SyFkBeRipXvzTJF/ZVjgXRYfvIS7B5W9xJ8Frc3H0tIG
lKt7FQDrKSFeK9KBTfJM9xUPBW3wsWjlO7LidnWut3FC/PmXYt2cuFZ2ai8N+9USKlk/EjENwdMG
OMy/9+fPXFUkOE/IuAa5YqHOuAheKBjy/0yzVJABxAo6ciQQ5xV/dh7YyZYqkPA3HBoitQNYQMXf
DPG0O+Tw7R0NDBPi7WG/09MSH8vbdtN9PlvBNcxoIbNky76maefWWO+yM/zpKkKxZKgOoXPRRDrv
NHGFnTPlGKJrPW0J4w3bNIgDJ/VNiJnoKG0Fu8z1w+14r/o8UBauZh5JJdmgI35U/Eb5ee/gonmT
BqkAHOUvUm82zyj12hdz+yymJqzfZtdzlPQfsY7inK8kgyzgvIJnf1vpgfOL8XLKn1XuIL5oEl9v
H4HEpyRVOjT6m+gOajzlsTK3c5ydzxxhw5SMMPVqhb3V1/xwa1KxHdEYH+1ZZ9IwlQdyHafrX5zr
iF0KsNZ3aQ0EOZWgqzd/23ZTxZfQNO/fqQv++Ry9VsZdJb45iC2cK3W3eLsoHRKh5SbfkM7y1Ykz
QfYN0wtx7+uRDnVVGMeUXhvSrmBCmxYOXmaf0TPD+rLAAgE9AGUCuuGEdV9+vf2Bw7z7s6i/TVzC
nLhMdLa5OFPXrE07kC0wKK8b9nUuH/Z+QYeqDFfJN43zGmmJw83RsL/nxzMrf2icoHUeI3TQZttB
cWIhPI4mYfxxa4Sz+2EtmWf0e7hkBy5a4m0OWKzrrfqgCkEM4mSUbpDYIb15aeqx4tNcg2PamvcM
YzJ+dH9XqOuXVJrW7bzmnHEbSfFzYnOXIMObYjK72t828xAladKJqA4F3EWT2XmtKkkMUSsXqA/L
o5PGxf79+tA8R9ArpzJGg79kjGiaM7080SVGwJrr/+zBWss/wIjG032d3IdiqWXHdzZa+0glvvZV
u6n/0KdHwxS1+as+T0/6jqX6yxja41qlkHGhg6ln/IDEBRp/5AdDT75R5JCvax/5lODy7fYo/XPd
D+k7VfAzve63hkalWOXuWr4ZHz7Bm2w8RXF25agoA8w/KgJaagEpm5fBu2neyC+r5TpBZ7fQUNfs
2VrKLMpaalSl2qqe7E2/lHLkzfzZfAsXB9YP9idU0Mnk7ikKAONeG6zPtk0jOAkNiYWtR6NkTrU/
Vh159dal5hwuFaQATOoKJvxi8Qbg4QiO4OZyZ7RMr1YMH/67JMhb+VhC7Qd2+ZCx3TEeZBklj//M
oArb9ed3637EPe0CJZ4gSIwM9eU2cSTuP28MwUmNj1ndzqGczuHaXUdWWFadFLBnyTX31RisUrHg
s6Y6r/UTNwFhBJDtnK8dRpjJ3df1UjK8UisORRlbijY1CER3X+GZBeZO+lsStsvt41kfoCp1Z3Nl
li85fqQX6TavEVQAkHFMRN3I6l0YYYrziR8JscSM3EqcGiui6IzBc2ybnDGWV6LHdNMFNxIthUPv
XtmmIePrPpO5tmYMEltY941J5AlZXo0ExwPcPOSV4i54SpHlriELlLYC+k5yy8OudWZ3rPfOtmV1
9fHRZw/PqLZIFEVrk5CSdQTcoVT5HJxSZgrxuxaXnyGg41nt7ySQsJmQZGAjAgfcbF5pnuWFBw/Z
32bS1yBy4cqJnCNTLLtJXf+nxGu1DYlLJGbeBlq0W9aThmBy/8ewA1xt/NraGBwkQ51mdCdtHcxD
tIJ6sOmj7tllWFyg68KE7/uLaoN5H6ib0iL1Glc/ySALwxmlQ0JPSyKXmi8QaFHuGzldfzKDrUAA
jwOpmkxNelKjWUK5CWe/nWVoo5UFqITpqyXGLyNUQpB2cK0LjoNDZKhWdMfpSAKChg+5bSyRh0Q9
WqFVZe7sorJkU8NKPTj/p6H/mGXd3wVqertq2CMOalqeVIkjF0xdvz3OuM4Q/rY1JaIfqHTGEXHN
si/8Qmh/1zIvv5ArupAJRlz+orv7GUPe2K/fBF+JQMypqLmnqJT15Kr58KxUr2vYzyO1V/A6GGmL
YZNHWeEQNJJGdG8aYlqt7JD+lM5OHNYLgfoy6VTcstaQM1mb5Scw0KzWw/9SWp8bkLCOA+9cY4PC
smXyNFmacdXQiAdjzAlq87nWoOQ55Hs3v11rNE+3TLAHqfEApk6QiXAPB8o4ehH0/U8fNTWwvY15
e67VFJbxYKVuDqZqfIJ3jhREHQAXnTyfSb+BLVcplVHMtHky9sAsdsTWElos0CtTOtLUYhZGKtbv
xR81LFjz26pfPwooZjeHBAZ+MsnojZvfjgP/asgO2GVDhjbGFrvpeJnqGlJQSN/j+vaT8zncoLVK
ED8r10vZfZUMK6IJj1g0ie483hSWkm5KHA0u65gW0AE/IKsdTzpWWtEyVW1iK70PwpxN1E144+Ke
LqZ12EYndSoJAzYu1iKg88QmYdTZWleA+s33EzeasO7QZgAWiGx+BDi2rPJTQi6HvLe+XvoftldD
FDPQFfLhRquvfskG9TwejJ/Gxdg1Xa5f///TXRIPHAgQz+X6nWdCleJcUprU89sJm8p/pyeYSgbs
uJhm2VwfmbCyNL3yQ/gZPSjadQS9Ao7PctGWp2a0b0ysLBHe5FZugKoRi7loFLiY/V64Qaw1ziRN
YwuDH/GyBfWrUr88WMBH+Hb7O1CrgCJryPr6LYNbAavChoQ9wGoVQ1W4QFCn4NlbkZdWvZ85+cL5
OvFbILegwJ3fdM1/8IjcXZGc1P5vxkahbtY279G7SqqXoh0OBIn8aNuXwU7i5KTPfBTq1bjWUnxO
KTar6xTCZc6wzPZcC0h7iC1lkzpxA1Pk3/B9pHAV12ZmonU=
`protect end_protected

