

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OJrNPv25gxVf6MOkMLDXm9qPvzcLiFn6cGPtPoJyX0DRSMUs1CiCHluul8VfoMGYUnRu9NzC2pDa
fD3Q+Cro6g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OO53+YxV1fz+fdQXiBafTL0TfU0s578DnGOkBDgcp0ZiS8qBHyL1R2PISafYfK37QZ2xP9F0gTav
+sG2DKzZYRShUhSDZBSgMOYpY7yZxYTXlswORtjPSorUAG9VDaJFPSJUqemfgu4AY+n/BsniNBx4
zqFaZSDmDQebEViRgn0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qtwd1yFLlmEutFKAPe2eqNz2v7W0I1lWfaUYyRoJyXavTq0FDRoJFjh1vw8Id+dlXsCh4QCKBOe5
q6ztRPULauE2vnffEDrTLD6uStkKikAcWpHaB5kHv8W/IU3+JNz65HQM8j8hOwGUzUSaTQzI6Edd
Kua78SuOo2L/RNS2CApKLh4UlLjlkL69KZuDAj8Ds+wPTUwjY2h3tf4V0N6PH8lPAy9xJk9S3EgQ
ni8vjkjW6lK8he+zqjEtOf7IEGhelGexSOLg0dP3NDhMEcaxfcI7Zo8kOCl3C+GMy2w3TEyTZkQr
3WrfN9WllC++Z6rNtRNAqHVgNVA7hObPvyuA/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y5YBoFz+YhLFw0DE8aie27jXEk9zfvZg7zgS29dcVa80RbYJrtSDIAboa1ixJiDhfiME1gY5XfYR
MSxbx3I2ZAkTI/5DwNAjKseDEksXdqu1CBQcg+U5NxNg5wWuw+vr6DqkJMxvZoI9BhjAErRu+2EZ
DgyTp7XS17TjzQ/Lk3I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
amEW+kSm8JLnUlmLoRCPt0pU7eCAirRawwzTZA3XEOaldjEiNg3FqPsvTGL5ScrzO4MhYsVv9max
1PQJ/lU1FLIUBgG3vy1UPm9QWkUIWp2rve3mDkSCfvDRku+GIP+/ziqovgiDyF46b73fS7Mrb40P
ha2QhSaORrSFucLp3v+D7rdh8lKmMq3YY+qxM1KZEpdfbausR1NP2yVxQP/t1g0w2pAjiWQM7wT5
6xmmRvYxl+7EuZQkxaCLozCO1ELg5LiuQuDVfKRWPdTIjtVbbBvnn/eTARAw8sh6+JXXfmhauCWF
cGkCTU9noi1D4Z3I/hvgJ8IXztgyejVNBMRBwQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7392)
`protect data_block
7YGU0lYmgr8yyyA0H5jx1crD0agcl6bbbSk1oN0BEUSH6F7D3tDbZuy7hfpf1NYYGzSCVbxMz/PR
xrX1hcholh1SNzXqo7l4Q1agrQzx0pANpIBLuOKb8STt9zDwkN/bjgrPEJodBpRA7lJUdcUz17U1
dFZWVQQ7577IQDw19kWOnUy9v/2W9u1sKwyGxluBS5nQpJFR7yTbeRWFIrFN/xJpPSrJqkZibSRs
hpL+xlP4TMM8tCApHel6b4/NrTiGFEol6vFreU8Hspel0QKABV4+1RSuRc8Qzu2A2vM3jj2nGPPt
HAY4Y7AMGHMPu8f30wtCtHxSjHEO6zZWh58ZnZ9QP+YtzQ/CvqS6fqVWi89d8++CnWt9YqPruWI/
2HmJjRtqPX88t3nSV162Sq2rzn63A4k9xP8Dj+BxH+gwKg8DGnN5DFwHb8lM6di63oOlLp4ZTLV5
v5FrAQXU2r6iwD0JQX+0H+DO7wteSx+uoydakoKEV/3VxonLh1KB7N5h/KJp2mXUbLzrPL8gmU7F
A5Ao+vjn3y3vCYo5zBgHt8FfGCg2TjwtxHa5BpEFhDb6SWVjDP1R+EgJN/I7Nd5W4aKBKIiyZUpb
SeYJf79857sdpORip09Z+ZgzceTcVErGWSkciqFdyleyvjmnhmpnaICCzaOCdj6z8cphSFl3vOcm
O7jELz3XEYCYoYXs27lHHiAS4q2Av6DteSJcby3N1Lhkn7oftbXws0m/SSmc7Ylq9ZeyaMx2CeT9
/0UaHi9es1xw+2RCraHGCYp8t9CLNzDtv2uoqTSfDlZoTF8hv/KULormiINA1z44S7P857gAqx+/
rorqwwgjDIxDrXs19vGz2w78F6j4+L7GWbdHr5tyqI37utcl+AzozDLiRmJ3CKBI78iO9E0AvOKD
3yN97kOyzMBCO52L2PVBllGPiRLomQqnKpzH94QR4p3fBVShE1O+iC/mYCsNGm8XNnLN8ObAJ002
AmvPMSCSydZy5IndgxjSxDnTvdaFo9lQK5GLsqp12EwHqneXQXHQFSoU5FMMvH1HveItGSoxVRcU
yxZDSlJMADzYm8NeHIFUENIh7GzsYeXqHEPMX7UTWhf6iMa/vKepk3WmwUIgZqH6ozdQog/+2Hh1
isU0/Ve+Xwug3+E2LbcG/KzcLToPjFM/IjUl/oYOxDkTz6KPA9WOGMVWJ+jx7GFBREdimR3TnAQ+
WuXzu+6YoLzZkfOFXNzXr2PVEA9Lx+zGXsjOK9FY7yP2pEdOWS4qKBLNYaJ/Ia4PhZpd73a0GPlG
x7bOnbC92/hZqgTfmdtRUDYi2TZBkSLYz+S4wGSaZSjMIEdwJNAk8ucf3t/JZrWvC2QnDalD+4Qd
17zdBSiETgqaGMU7zT4M/mn+C8wkZFcsqZcT9dDiRofFiWoBmk0fXB2PK9MGjoXLQdgtPNELa3zZ
qoe3cRHr3VDT3VLfKmBExZBDJYn1ksXZxpskTZZQlGhK9pBuLNjD1iZyE8JdBVSEQ2lsJnnbuVhW
sLLnWwhbduqm1edjcufdSq4rbI63YNRzKIQd4zCmgT4eTC7xMWvUvhjD5qtBpFPO6r8t1ThDWTVb
TIGx515iJ0W00Fif13wVkA3/MedHGN7hLHRaA/HyzBWr8Hs1TyzvaqeIU3kS7CDw/PfbOXHmyQ7u
efGmIdpARq+KRNzZHrWcEjcIwBroZyMGpHgimaJu+QdcaDRQJMo/OR/HtpisT890wGMPr+sDjFN7
B51+1BBNLODTTBT+5pJ3+9Dq2fYDmtzOoRXjgk0rzbx+M2glKfIK/r/6QvlXQcls6DNZP7QMotXt
87Zm1BAnJNp4Q8iLmXqj2CuN6OmucJJ4wXGoF481Z/bWt2Q4RcyNm+ctaBFzSg6ZBBats9b09RDE
blYZ2aF4OsUfPZnkQYFuiPldUNzfvf4P16wE9GNJMo5DkpxJo1+lH3lJ2QMJq41swi5vuBBrl21D
m3M1tE+Rbc+2ZF25lttLXG0egiUjEYupi4TyugekGaSLKPS7xWZQrww7U+5tw7Zyop23UQM65+WD
P23zV4vCe80VBCyZ/ncOJh7xI1fug+XpBg9xXWGII9sSSyf8VoaNWsiILoLjrrGcKAaQ66EgFdhy
TLFZ8jShPWmiS89xiQl/VvBDANV7BZb/0qMB123IULWxl1OVYWrR+tZreKjfurfHb4hzkPbXHVkP
DzYDvKiaNRZz+URP4vODMv+Ov5g0xAtXycRs5DZmjQOC1Lx9HgKrJqozxhfg6TLvQHM6CK1/na8w
MjbgXAQ311xByEi5vpQkJ7dUt9d0xfHLebwgtHRwBEooiofRNgQSzGxM7KBOydap4Hbk41T+6GDU
fAeIEiSDQbT3tl1uZFaFYl1O+T/Cs5fltepkdgnFSFP3ZdILxccPtKEJkIdSOk3BPoVDTtCe+j/d
iRI57A/NErI+ihor16kBfeS7KY9SwNF6Ofc9XDjfcMUa5WX1PInZ2/1HNaJ4yLWMRmf1HYnIaBZK
EQG0iG/retRx4M75fmWG3/EXk54Xltwjz8ELjpFWlxy5PvkWfFJ92xtW5n+Ywjv3SMF5bYtoBHjr
nKBriXufWP+OM98vQzJPj4vVYjFkZ7Nt/Wd2+BjVUO8AVssUINJdGqm9G/MSCMu+tkKo5Z2zY+4S
R1P2Y5kBmi/2sfyeu/ZwocMnhyCIQDIkPc1lQsGyPvlk32G4PjlrGM4TSn5qv5RO/sUnuGYD8Tvz
LA3QKpgJN1BvI3LFLTLub2uhlu0F9f5e7/5i1Qb3kdt+N76DidqJIjivViwDUuminVcHwetDdh9K
u9Iq9bGz9j8QOlhKlv4eFx8pJxT5RXJQ4jGCGq/1BKcpI7t7TxqcKsEUYZlHY/mT9hkZyHpO0rXb
b+hnt5fWLVCayRgMPZtnaS3z94wTXcBG+XbNFxqaNGkTngxkMeqmOLIaXqYDFFfOsITHyDAl6A8a
PIIgkzMB7gtfxZMfzeR4ZgKsSDOA4nVd6lyuQEbRBJVDlXwJTwzT+LSgR0UMZUgpDQ9PPYXX78Ea
pc8hnSfU3RBka9VZcpsV1A+kTZgfRaC+hpQ1IONy80Sd2fjHsZonBw95fpnmGB0zPFK6XaDdpQG+
pK7DT+DzUhjBL4eM6qGX7YEUvowgmeRqA7Y3VnBDeNHJqyOCU708+cssrwLR9Hx5Uv+6v6uDpLl6
RjuTu4yxWnEe1dtONBW8J7Vr0g4FK5M4ewqtjz2UqwkUwq/SoZnTl22UaS6Vi9X4RYb6jdx37paf
8ZAiNM0A++ZtqBNwq3RjpXlEoDsl59lNJT9NiuAzT68Faif/6rIAxDqYFidf6pqH0oaY1XkHz1yT
bEgvhv/DNytfAdmSKve+pBYhu92D3GaB2r/4Q1AXdbUHtR0UuQV1QY8/WoLjZJkwv+MwlguoOKv2
Y5Dn0kQ1CwtaQSnNjBi/Id73suWZUZCwty0BIrq5hlTEA2DnKDnpkUUVNKan/9yp1GLcJtvuGBK4
Vd/Y2ZsNh8RBdpr7uHDKOec5FTQHEv4EATMqQ3muqBh0nlfaUh5oX2Jfl3ynf+AJoCStBIIYNsO/
4i9sW8wdZ/vQ9CdgaTaxt9Ygfnlo1TbnOh5MQVM4QeIDOZhEzGjGi+SWCUPoQgNv4/DHYo9VjgzW
hFZpS4OWM/2vOirPhfW5gYDK05KZpMFDSCTXJwAwjb3uYrD3zZUx1l6sqj5SY5RCnYzJK7MB7PCA
tYMi9sn/4oraVk/INJ/O1ECx1fWs56jbEmohFA0nIYZmoqbk5kZGkKDz94GAqIwe6WFoEtCew9cG
CuyfeET3LdP5bTE6TFA/H07rq4aAELaaDdWr9tZrfGdn+FgnlFsBgG3hZiczvXv9Prn/rv8UqwES
2mTOBIonGgHM6TgfItMDGB0ou0+bU/ijkq1yNy53PSBX/mnOf6eVvspKZbLlsEVhzgB9ieC0K2Hn
k1zMx0C9sC9xYd3T28bpuMPMWWaXewj22LDjeyC597MzhkruGTFXyauszqc4jlo9tksAr2LK2BnL
7J2x3ReqavlHVgcu253WGW/HgDw2ywqgcnYAXgKl2BFt27uY+udl5a8i0ERsvOF/q4pGtY/s6Czi
WCe6YeomUyMXJ0gpFNuI4cNdoz1UMtkugydUdsUy0NN+T0NaCCpGu3AqdYMXxo/Befa8Lf0QDp2F
Krjo/Y1i34ZCANxcGxmkvtrLPUU8Hc1PCc/Gy8ZK/AAPrNlnPu2HqPtGsbc+24fqa+zV5HL/3va8
d2j1nrNKYPJMcdfSgv/h8hMjK+af/2uWEGwd0IMyGewFDVPdICryglRntODoe309IwHqfM1RHypG
Zqz9ynzF/Re7+WuFUNvMQW5Ls5Sdm+WMyRfcof+8QXd+dRmnALh3yQnwX17rIzvB7fHHjj8as2Ik
uIHYNHaXxObon71gWsBY1OQGpI2tmOS8yqTWmf6JpwM476FAGiAp6yHhwiTEVyIq0I+UTDuX66ps
Yn0dkhhTPlZtjBRMVDywJOJ1A+caUFJlXTBLr2fb7naTF4RftUh/S6RGmTcrkrF64D6PRLz5xSry
e19yLgp69okBSnR0Gz/g9VLql8YyRtB+aCcoU2Gm1F7207bffET/60ATKT6lRn+TXpCUwlydCl8P
/EhyWHjoXE2MDh+J9+oKgdTpUts6Dfrnx/ImHxY2hAD4nwMT+60C/yeU1gCNzfC9GW9IuTQlXyDE
xFZELZVTSWaW56JSlHUbS/m9aoAKsU32r4FGG0hv/bS6k1G2voXbvAMUS3pAC/PCGASc4DXfYZbp
0z1um1jpCPesiEhQ7/4VU+GhhPw0lGXms32T+PwEZ94b8kUsxhm/cBobVueHkAT2OzlAZolQL09D
BMRrXT8n5ItTCIIxzG7XwDfXzU/Yn0dEcsD+gGkIxNJXnja7OTdoqKu8Siqw+uN4zRcEgEm5W0XY
aShUP8ii/lfHWHby/fPmBn0WQlqZ2/++JLrgn2zH9tifBMTq7xRmZHCw7Z09tAEnKmXvy6E6ODz6
aMUXSH4gRQAU9v+OqTzmCkBPYl5Lm5PX+q5TSSRyLEcc7/313LcvH1fDhpKYimj8iPlK19aAEpkA
cHEElayneJzJqHV7Elva2c7gX9x7LFRwk/4DOBZWL0E1koKFygf2/+zUUoCDA5VSIR1tqTHr84ou
3B1ok6EqgDsMb8oaZiTITq5Hkwks8T5O3OgU5fevSkWW0lO+NZcIe9ymgR/eXnPxFIxU3kukON0C
nkZ6GYF3oR7o5yWVg9u5BrZTlVKjwR0Y0Z5CNgYGdgAZYdhsdXqEwtKW+utirxF6XtsqWsTRFUZH
hjZNKRIKKEAUo5y4LDM/BaSB9FTVvHdiYKB5E5pSAyy/lcvv6OpX/6MBgGUzf7CxgRgJ5HwEdadq
FZ1pZefy4pTmA4MKWFRWK2pgq+ndcwAyHDR7XIlb4GKda3wfxR1/l91v+C9awO8UOrmd2hraXPr7
wy+wOzgY1jdLZszxifMK9UC5JJp24Oe0U1tI2ArVUKzqRSLlV122ooKUJqY+Ftj5arjjsFfdhFsw
nQX0HSIG08KB5YY0Kiq/dRjFr+SgoeKJ+gOEPS0/L2g+soFfmUYhvJhJt373mWY8NbXewv9gPZzD
/4Lb3cXOkUgoZv9rJ+CW99g1fuQcMMMLgD5672mlgBt3ZuCFn76MAvTRN6bDRq/Vbw8n1Mnpsbrv
Rzfg5QKkM2tUP0xXSYjDyiYfCbYIHhhVtn8I4Xq2+WjN41HCqjgKB6cqdqhrHxdeFWUaRW+Q4gU3
JwzRdV4JB7X5RxZMzdoQ/JlG9RDdF5CT0wOGMpMfphPUC0StBOiW4DM4DGGXcz37f+F7Hf9leQj9
57qSR8vng4cSy/WwkfylAjPAndmP/dL0x8E7Q3BRxCaW7CDUtEesRrjcfO9CrYvvd9m+IDhhfPBL
iIOU3/EYpUAq+QBOBiVJXKEtfUz76y5OnC5a16f2eJB08muFuIqoJc5e7PpFZIKLkXt9e4bUrKmP
xhHvFb+XQSYEn/hHiCbMjPjGpX04ICfkLRDCIsutSmXG+u//MfADMx57+Yz3mT1hoOsJXW1tTdCQ
ZEoloP8sZPsA8dRCyLRDQSjA56Ne+JWznAhUWSdc8h6+Co1s3b4/xigkns/aMPJUnoUMhK/qVqqZ
Xu9GQSZ8di/zhVjiEVWMZjrEbQd7PicxmayjsjQi9u3UbCBZl6aoeO4th+xOBOs2UY6f1py2/ZLc
vY+RxPJYuGrStdO6H27Dt64yHKJHv1+47AwW20vg4/oG6KJZdJPtetKh1Q5FO+PGg39kJFDaWbP8
P7m0C7IJUTyfJJVKjqlyTrocF62IPsYth7yeXVbBYdD+pmAomqDG0CYo4pPR/bvtqOwmY9Jl108Z
5aGPv0+QNn4cCZkVHGX2tS2kghNKwTpYa/9Jskrx+cdvD9vd35VbiSH051yV6yTnTxUxwAT/pHYy
Mj89eu0T4ePWyxmq4Fjk6RcIp3HgBHOqOySrzjit4GlVjQNHRD92aLbF5G9oxozWw0ZThkA6+1U1
vs6fQaaOrC65RakcnfnhqNl89U+aYTBsVcW5yyLFOiGmTQhUoNJSKsos1NFh0qqblnCQ6QcfX8Px
7uSR8NJfF9cBZuZaj/FWZ4PjWsEZvIUy8yWERhyxdgh7lMIwjTFyZfq8E8bY5mWGAtvuxXyVjXUn
LasRqsxqmYBwVs9dTnpLS53DnrRpIAO+8HWK6e7aLlPJuxWO2evMgY14HddfwR8W/VBoDBI/ZLxe
adaNPLUtYYGiZfUaWhN0KD8vhofrlsvVAk6FFFvXB3887jbfGOqO58kxR2yYsvuxgwBe9/zFY+78
1/sydrRhTpwvGcGMnhPHGbHk6ti8jxhgP8Nn1QGdG+mGCyduNj2suQ3upKllLAnGzgVdC5sXLMtN
SQjAybFL++/bFuXIyQK4TEntMT+EMWiTtbluf7Hxj59Q+G+n5Djy7zxHHirGQqXZ9qx2+phLRlHv
ot65W2NL53KbRCuskEUxqfxxYmGyGzzlYUccS2MmhnSyeljKysqHhrfzDdjFXDvjVfhCFd7X5CdN
NSjXVf0UeCKD8cx+HzMq5EJQf/HfjDRJFtrkOey2kLH8/j9vqfIrqOSLwxVFdLe1Za6CHALgXXkH
An/4+Qe12wNv9PSMA/z3b0Al8oNc7U23zrWBTVOOIFA/MUEBYDSa530oYhFnvIwfxLRxWHpDOVfG
bpPxx5YxIsYhttuL5THX+lmY2L73dfACvbzCj94R9kI0djXmmccywu3xz+odlF1cRhnolInAIspc
ysW3NUSUxUSAeYWQsaiHQpUQNJgNRMmdri5z+mFliA/J+ZysiU8Is86HxqhTVwbVPqsteoWAAKh8
hVjdKEIVzG/paB7YuVI8dQcfz8Agr+HQSLdLTEC08EireEACffO8qHFR1MeOiwZXdcQdQVTgNFkq
NDMOjB6AfUar4lCUHJ5MFHMAmDUyt42a94mzl4OeIx3CMk18502xphUUdeAXLdyMM3tli7MkSwfl
RpJbeq1Tq0QOK95AydH2LHxr5JKAlLeN9+EO7kZ/ylOJkcxenSPkpEltX0qIKWGGFfS14PGVNUIw
dlNfRRG8+OTOIDi8Eg8g4BqRW2kqeeA2FHCJQiu1c6WJ+fHpFFfBoBzhX5TrqVCs6AP1JIYow4RF
bGlaMbCDI6gePNFwWrC92fJi7/CBTqYvUD2EnpWbimVFvYMOZmmy3RUcjw4CDBHPPScm5DLV8Pl7
QbmsophRSu6DDeEF7oW7BUgux2kOgTW1B8cqy9xIgWim/yNeyfIUqS9MBJ6zGi9DViVdcZqhvp14
UkzUr0VVsYZCFMxp73UEFHldlCUfmYahIj3pZrWMNMdlAqW6Q92ezOtYhDp9irXDrscoE9Gm8zof
U6ujaiwb0VMt4QJChpRP7uHjqcaXP4lLldVvr1TFmdJCNlAsZ0p/rkFcBptwMN/u4WLbNu143xZS
voxTAdlhKnMozAt+jZeLeBRE77LpvrMuCR8P7LGGeaOVnNoDkFXZOoeL0T+HZfhZdrUZFRGWZBYa
b/CA6gpNCNJAbJbtzMwosv4bvviZ1cHQ+1csIu9QQpvor76JesVdmnkf+PQaMzIxPDaM/wz4cFVw
nHTfmMSbH8OZKMS4SSnLECrr1i5j7vbsQiHWRS+I5yffiqOD6ktTNGMeOLK7TkhMSPQVjg8Kd6xw
ZewySqKp8o3J8d0Ozt7DBVEW+DqU1Z0WhhNXPM8uXtVUtHZrzGjriD5tyNCTyUwzf5V0I3MFpuvy
SVb2rfw+H9TNtYfvNAS4edcV1NhHt0r/gBLIWJAJgHKdudMExQm9VrITxDPhT6ZPzfFDAIuLT+UX
JFleAAPa2aIPrRvolCDdOQvEcknK7VIqwpTyooXOGW1E8iRZ3WXEmjpkk8oKJ3lMzhkTB/Wgu02h
HcCNPXCPfhVS7jeOPhYiziaqJTYQJxchCqYBMJeu52jgm5XzJk+ogB2W5rU3r/l53qozsG8TaO3u
UMa9p4juXxf9w9CcC8gwy8WUxAnZME9L49xLHakkzFohTChNHoegbZDfCodZzuxp9igM7sD9UkLw
hb4IxO/YMbMLbkHJggWU/JPRTdzgvE7jjGYLyTpFv+0eBmDmEm/0oTGjSMaqIddkZPxjV2MuohcB
cy+fJKFAFp5/uFU2l2IFbp/v14Fa/36GVmTxM/DsQvAB6j/OufsBmM6OwV74KCNHWYMxj2Rpkh7p
9alsV14cK0EKZkcVsV8Z/PnSUJ+XNsVEjwbPa6Lh95ykZWk62QF3risHoiHKfBevfoUvypZ+elEL
DgzNzSuKffLKJiRbo6uhtn5+R6yEvD4SJpSrooDyxxwAEeQ7brOARO0AqjEifurh1ipKYYV0DGxC
ZgDIaBgtUOtuRIUxVfEVmrwm+dsAOP/NjQYUdff4aevu1RRBLc3418c/MlQC0MRlM2QP6+uYa6Qq
Rcw0K17rDrJ2fS3XdJz7KOe/PwjGaXbhUTe+4yY2dR0LKzFTc46I4xL/f0sKzq5IYTIN34KmEz+S
DT0xdr807ThACa2QxvQhlSnJHJHAu+JhicrtNzl40TI7arrwVLOzdqycU1ccympih962DR/L8V0P
1bi6DvFP/iKU3iDrijZKE8dUF8V1P76jG6PmQSH/sWQIufVmlexFmRQ7GbHifMDUpuUNmaGef4z1
mveqvXi4JHrNzDpamwP8uOjstUIKil+fQo1LqfWNDWmXYHfiskQlEaHfj4tnsLIF1fB4wom+K4MD
Qlq+5AYW5uagBBbYqnzgAp9MUxF04kE7ly5CiK4lfyzSV6wZ22r/zQ/kk8ee142tRs4b+L+zn1IB
QwM8xV2CUm/c2xEvSBRTdkvbpGo1i379ea0/uMXcIzXtrqZLbvHQXMGfyMjhhzbe5c/+/w4R+CbH
X7TIxRPsPsBIm6cZcBsHxRbfOVGQilHZtdqSZafIc4ImcmH03a3940mEu895m6ytqu3NfU0rJkt5
opft8zr7Ki22nodmcmeYLQ64jmacTfu3I1d3yVpJFgA6vjrGJBdN0vHEFpfnLFLyJ+4ygvS7ZULV
pSDh9IFQVR9CyZWqFpCaqQEXMIxPGp501ozo2ojYKLzcuO/PraIV2aupZXWH2SAliXyC31o2EeK7
Q5izrkOfbp3IJjnFYj9QHlK0tfkjm5nK0GLgRhIZ5nJuTlHTMD/W5hyAHvOhb65wvHlueinwRpXK
FrkotCuHAGdYIhsxmw6u1a5/G161uXm0LTtuS2Srn6bphtubhUR/gb23ZhbAyx2qn29PJmpaox1d
ikcIDUiw9mbYNF97LCXkpl9P2c9QsGygkAC8dZm3ZBc+835eE8wt
`protect end_protected

