

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IoOiz+BDpEiCAzehQDaKkNxXycZX6DxCheIbVmZVnOeE8xp7Q+9Cdt/GYV8eq/1L+MpdyADA71Q+
diEx2Z9pJg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lwiDFOkaG5HcqeigSQ6a9WNJOSnncyPnebjhd+6IKLZk0I0Ny6LWNpdm2fV6AG4pFcvx58T5yWEl
Q+/SeuKD0HNAWdTl0b2fE07zxr+edW2hoGXyef1M8toS5SeJjbmVYB+jYYVGpq6G4uNelAjC+U6H
qvBM4HmLQCceNGUHSWE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UFVaQj8UYHzOV/s9ci9b6/M58BwxIhqPdXQ4yEijf72oAEn9ivW6AsDsNzmhpHIiBklSohpBNUDU
0Mva3SAcsX3+9Czy1ShJ5GBV/GrTCNonRWGYRXu6d9ADAsYZRaJCV+2s1kEifAqI6MJhteonJeVq
EumiTmv57LCQxMW5bGdt9ducpN0oI1Oavkx+FYROiHKMHPR5ux/CzqaZUlRJQvJOcmbQcmUZt3v1
KBK5x+Z9B/aBdtf5Z1OOegRTMkPGAdkXGlAX/Ax9OEiQYDv905iua1b8cAJu7PD39JX00W/YP189
CxrWyFNefwoc+rk+siGiD7Jjf0ooGeZDZmjyjg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HK3O5vzCNER9g8js4SKz6W+Zie9dlDlDlxGQF2WrvDyya1unL5bBpCJy1w0Xm1cUo/y5lNUI/ADI
uYqE7JGFvbSauhLZj4HImoydapRAa/ZLL9nSRfszIVrPI8v6qGNzlAIC3uzmQS48iAygYUrq9YT1
qPItKzIRjW+YafjsvhM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
haBqrpdC8sHCosML+5AEE8iaTVrDueP49m0Xd+C16lJUg1YPcQ6EHNHA456bk66+nGBPSp3B+PjS
04UE5wn9q/J8cGL4YbVE/GY5wVAtR6WtFplMeOXISx0KcrI3qk/KzRrP9Ji6/ivM1RBF/A3FJtrF
qq4E0RTyXYa205RDSyJAQ9RjkwZRwEtkcJ6VY2sYCysbDHMzh/lD130AUg9VBNSdV8LSRVpcwCzZ
sRog7YjwhxC0jQK02UyUpzfW4/xJ7RqEZDh6icr8dQvRuVfwm4y9IzcnYLipDLpn1iVw+wPGS0v6
ZJj/N7hNXBnHUH6mTiT5qnqc1qaRllFBLOzRgA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8144)
`protect data_block
Acjyn5umOLoD55tK5GUAEKk9V9gS22UmNYhG20RRJrdy4KRsSGp2QvO5C572INIJK9GAcZ64kdzi
LVV4x+CBLD2HkU5G/kgbjzkES0ZCOmy9P8T1Y1BfhblKxv0/to7EyJBJXDbSVa9uRrst6TjxNrP+
hfLtu2vFYe3hFKnwq3ooKun9Q63IVkF592meS9WAOLPUd1ziocQ8LyOqMvm/6sT1yJL28Jl9yZrZ
NZid7pXotj4iIr0BHDL7S/nxsJx9SBkK4oVsyr0KcgB+1LIrlNI301HTM4306H+o/kFVPgIxfZ1B
XkjzLAXrG2ZdgBGAs4O+YtrMcrom6eI2gndMXWD4v6AydviOdTtxgWcHNN9CFdQiKQ+sxwuWmOMi
Opvpt4lPwWpmbld6qvkiilwowP3n3REQIArn0RVxnEjtfGNDypVbl9mLbPUrw0DZQfZYQVixw0Sa
w6zoyhUgDS6cNTaY6nUEqy9MOBcV7Ws5aLMxZO4d2O+m1A6j5VmkOWL8Ab3IEnDh+Piy8oGs7qJU
yCVBjbMT6Hv5OA2c/R8MdtRTug1ADqWluss8BFYq5t3kjwm/P83yDeW3PFIxwGqRpTqEUBtKhBAJ
K7ovxaR5juCewNELgZAh6wXrBWxJ7n5plas8EdrMZhtNzrEaxep2AbW68mKrw5bWfsNyMKlW1cfe
seico5il+1HH0tzOuCIIyewzZEcGFwf43oD2Un6rL2SwQnoqkMEbiEKAgbfAMhR2/Owk+2OIlWzO
F1xjNkUsoT/efT5eL3f3HQ+GXwITZoxGeHzalFZrpmvE/3dZs/AkZIlx/DFfCiiy1RYT6AWr7/58
ivM7+MpUSWUq2NmvYkZj61w9l5x1/BNnjBc/prL1aY18yBP8uTeivfJfU1BQ70rZZRTxeGs/5EO1
UUGayH42CCp9bLtypnHrHK3foKzisoELBtwkumjFKB0HzSpFvMrFApcg4tqUAjEep2z/MWM/DLIt
LehBKEEtye4O+xr/IuFTDjD67BwEoVYPlTuIaNpG+SeWxTUNhOHPa8DL31sMBNtZG91NYPMWutQJ
i1EloX+3Q18QwlTvIzQsPjBDFoTLoup3B5Bisg5ytnvFN1S0JxcqbDxDc6sZjYJG96XVdgtES2cF
58vH/0EuJvLALReSf+xGU7/60gPQ89j1AGUwPGCvH0rbSaWsUwvqNwzpw0SsE7Y2q00XAWz9Dmuw
Law4/CmIbh0bNL66B6uTA+hLil5BhRfu7nP2nOXNojGbgwQRfxb2+SaWH3GZy2H+T121Aez2aCKM
SP/u3+AfoXFtKkmALwKarLp35y+OyitpIaWywaM8kRxfZzwsCvCwBnZb1/K7Ly9Pzols5+bAEIIo
CeMWzkaVG6ZEB21ZGxvwOJ88sK7zaWgqE6YgswyUS+4ZMvDGRFQOYOYOloBYR4TQCDqNl5vliW6+
Poa5yC/mQtWwP3z+Z/T2QlkHuMDFPsHBkgIeiIN74R2Ol5pT63vY/MHRGUAt+NPskn7oD1bXhu+D
xVqOrr+PlEnpMBe5byHHG+UEsNT4lSm0BttYSqVyKVSpN6Aez3jwUlcZEmdwDiZAdYaAiL6b2el3
PYRzJ+g+sOsvX1AtbTOip7QJA89qSp1RZe+lEzi1e5WstUoQ8NQKnxO1YtHTQvpe8q5RUCOuZFXD
hDZsyaFUeLJkcZBGrHa7YeX2agofyvaxIEFk6e2/JIdLM5Kn+w7ejLhdz4t7nAozNEKpnE77XB95
Bu5m5CMnNDxACm5Tu1+ge74twQbUh+stPbAeL5ifC84YvfRrJlYhsDdKjWIBl8jRD/8xjsg3jDIi
sDTSfenKjvczb2/QqcYPq8M8U5G77kxZnOVATxF1AD8aQckTuPPeuio89dWpXm2GrJLCIx1i4OTc
cLPjCkVFYVAful6723vOk0kihW+XmQHoON1ORMECABDNx905jncpE3tocnZTGFNfx1hgFSjv0o8/
1iYEyyAgLBnybyi9V78j01apON2q/o2sSkwaPEHP+QRr8aI6fcdMES1NrTnFMSUJP0crSunWKJxg
mDyD4mS5Z387C9LZts0t5/CFCJ63WUg1mQ0IUM9qoWRjWt8BEfs6HVxOAD/mpmJBrmdFkBKqKYRe
L1RSNYQOGFsJdWXLttHZ2jn1pSCEoN2fPC7qjdHqle8G4xLBp6erhl0ho41EGo2slvLJ3KZkWc6I
UxfFQrStyGsaZAI5F3bheYGl0ml3CQqM0B3aCsXF7CjwZhinUyzn5TRylNq4A/C92IivmN8VrOhD
pV+RbDZpKDmu3GD/lVWZ1pjmdMYJMu06JVkc/GVBoDG3PulmW1iCrk6eoiAm3cqhGgKsyTP6uPnP
K05XvlZGS9FKg1ewAXPI0R0dkfIQNEkYYwaal6AHJNmLfFVOse2fs5XOL/Aj+fDdL+fLQWETDXuz
5XuiVPVFFJW2I9comVQCmOETm/IQaZYupB+d+4J94QFWJtxcO/lv6lEv0d10v9f2FqsKP+3lupNY
GDkrzxXT3qMv1juiJ+tp+BAJc/fWCnS5O+zNgOsDmWst0+VRDvF8M6vKO/2UkxnXw7S35QlAVOuN
jTcznialABzS0ybe9sW/m9hDnaUzZLpOf3IJowez5Zjac21swvD1KT1JPUQnV1D+zzQrJVkyO/qw
C8ledkxqmf+mXGTVEavCQVlPuo4SkzM9jCCZFwjnydJmuDGMCCCw4Ai1C/JwYs2bRROsWy2/vLXx
YHtBq68X4w0gstDG/GL3ifee/g3fOd/Hhwq04/ggLARBVfQUV3zwVz4UVve/qYMbvTPo7WW7mhtG
a/G89KIWAlorhwGKbUBZ3fTp9RiBCeNClE14jvVeO943fwwbie3kUxqhiu9GTN23A71Qb1HS3gxo
ZNLjTKjhqpYUkStBKhZ70q4MwpFO/MmhgKO+LyZSm+7144kzBsMm7FGP7rKgA51MyKwW+SVC9sVS
DG4fWF3qh5DjYnewnRrtLAZwLYveT510CH8nRLwdSwT+VfJgdmgU03EtiFM2nuECvvLCtLNlRv+d
4nHePWly81Etqam9lJYT9h2hrChxm+X1s7uVT09/sWokyitgWWQC5Il4h25lqGxydqVOaqfFALhX
ckhfemGg4+Ra+S3uZdS+WVe1x8zDiysv/tHd8ZiwmhMIrUd1OIrZ+s30bTtQZje16V2UpE3UGjI1
6s32hEzOuMDL95Z0q10qo8FbUwUsd3f5DTAyj+cdfAzvu08YBuk/89Tzty+lcngu74JDEg11xq3w
Iwh2tGeYO0neLlel0l3KSLMq3HZ9xjtQf+xSqa8fvK6LLeHKOceAcUp8Y1KhsKDkLWFYUavncMZV
0nfVgsMoM1L9BHfOAaXPcncLK/n1rEy9a8h4gABkb0DiTPBUhvTU2ANg6BC7oWC1xNheVcWfLjda
+jIj79fDop1skpTLBc5OaPSq0a/T+ajmXVrwvve2QnPiMioidJSGNNu9midpLtUzFaL5AgdGtJss
5b64BFCrbmf9TGBrwr5Qb5DIVN0DPgxGP7dB2XxRyMFYdtcLM1onOvXN8zqNFHDfjyq2iDA8XU0w
h9aEQ1TXWiHTcW2qXiB7m1wFdevGn1ApthW/hNkIsv/xGPU5kvs7S22ADcS1jVKoNmSpkRG931c/
DXXHrTTuKZJt/Obq+XK1tO3bBBG5wbv/FdUMG7yVROoBM9WjHgir9A3yuktd1UJyQQcwWZ5rAO20
gLQ3ZaVzvp9L2e/ADy5DimsLLVDtlAXsMo226TmePvZo4elBLYT8tj3E353Wm57VwCNqE1o58bUX
Z0LX8J75kAoTCWLdfnenm63T0L5AxlzmImy2BY+tgaOZGwx93KysB4bnKo8qOjLu/IAYR/LvUivy
GFirod8FoZxn0WSuo7DSLjTt7ucI1gpkcRNEjRoBMDlN5HMpsb/f+GISGjg0qh6DDpYolAePBvo0
IUciqXGEsz42ET8HzNNeaMEMmEi76ezwDUfnuEfukfVdD18BlTd73NiX5ptPVhg88oWAI819CFSo
FI2hmT2gyUSRoc01uek+Mm6RhN/irqflNwLjSwfKRcTyq+TTtR/jVQ8dzCPaWA9B7hCM/DDJyc4q
V4uj+jx5yICL6n+ZAVfMvGY8qrHF3kUDsGklDNetUPEz24uecJVhq/qa4pJUGiuVUe7/0LA7rFJJ
3oxaRzoczaiYEBLdW7HguOhIOU6m6Em/B7gDnxArJPEOaoyMm8iflk8DBHPyerWcgyTdXq7js64e
krKtpi3WFLFIZu5fNZhUEGr/bQrf6qCfXCGHIuuGwaMvK762hn5Y4KSTHxc9i8lSg6QjbZ9vkXsv
WQUNORXJkppRcsR9x7COTkH7TpNA1ie0nGQNEOoTI/mfV4rF+lrHOEMS5tglBchtdqH8GTV8CjRT
lFr+PZFFRwOrZ1w6wPqgVO+X1cmocqsZv841myGRGWo6G3seegFxyzO9nJmPZdbO5B5crPopLTm9
gQ76cNwBu//RH8x6X8kTQ7keXQgJ+g/ffvlbSynTvq6gSp7MQ3LbQUgI6KEtyZ2Hc9q4hhMGNQnY
tMde9HZ7iOEcnYp14ove5u9i61yty5LhqNsSbOwAvqsSYYWlibwrtNNjHbVFIrgp+mWMLBJMPvXU
aNL95jSSczUgPb9FI2ADgZOMOvwS6E6F15Xz4vA4cr4j/dkY16E2TfZxAfYpyIZDnQxj7JFniu2C
kbhZU/MrztTaSBO52Pcs5y9/JWUYm5uU59UDiO+jKBZAglgEH5sv7QmneWWMI+V4oUK6zXzVv68+
OcwaD5eu1Yc/Eh/NENMj77hW7KZ58FpILxUW16QWTK1AeV2AkszKmg/5MO7J5b+GmudOGvyDC8H6
nXGj60Hveh9yRr/8d2JqPkHPV06UJ/0EuPrGelLpO/8B5DZOkHuagZjfcpfS3An7lRmoCVhWTkU6
DubrZAB2F27HS9KQyrJcjiZPidjKUq/4kvAhVv/FQ60ik65ajrCDVwweibLxOOHUTAiabEXUjZO9
xO0Pw7aOufp2O21BumVD7zZbdhTeOXXbygmuihn8/WVRssMB1KB2c+8fIOX2TD98BrxsZDa1Yo+d
IAuuB+sVt24p7fkaFKGxwXqZ7adD25P0UBCXjWqY7ozVdEpK6H+gvQx1WFnZ8eHGOK3CcEb91EkJ
l3kBPc9ldHCBiDdt2Rn/1/f7uwRY4xgTzJSKjpvzoxbY69Frqa2c3IobNsH9k8Aw9+wrv1RHzJr+
natrgvESCRZPA9IN5C+9zhxhZ9b/KVexo6O+GF6xHgzHMYuOT5ulUcoUsFxMC8m3AolufVvi2RiC
64jfXfIiNGJoY1Jh1aSkJxGw7S0268f7tAQaTTOgcQc66F+I3+o9hKCOD6Vux3deb2GWjVTdTt9Z
xZT6h9aKVjdnjP98n77ymS2N5LWcjgUCV9iXjmBpBEbEixcw9qgRX4MVIvaxaE6gUQ/vkzDnjuCC
mW1ZPLyxDG+dftZ6AF51zuZaMPbRknTlRT4tFvckKVxn9oLKF7HCmpikZ0Tk1MMoB7Jy1ZgWrjCN
NUddeMp1ITAN20m//HFz93KhK8cpnn9X/qM9zUypYFldllMLcuVomfkF5O/wpPoBCqevCnNgoTz4
Xc3RilqhqsuSKqxmn39JX0aWbqDoqgz5O38wF6BaM4uYheqt+Y7D4tf+4uKKVQtoUFr/5laWNszz
/NPbV2x53l5SoTFN9vukGBiiiMmsJUuMqpmmNwbPWQXxkck/JRmfEVN/XjgJXSrblBdvBd1hyhno
mcXH+wbzVnWGEGgYr8kt0oxU7dxDzR1x4wB8e5EfsfcpztA125Oq2TqYEMcQBa7toA4rKmiPslul
o53VV7LxzZNjzlJrT321z/wuyt8sT4qLzX538t1sdNWzLHxvPJONt4GOOshLprWJN4S5MuJydMzL
cvOK/gGiI+7JMmu2XUI0KBcF/quha9f7XReCmwJzVp+Sl5hYXe8q+qKOE4HEfhLpH3PQ7Vl6lCtb
fOHaW8WBWPGX6r8MdQHIwRHNqTOoNgYD2+iS5YnojXZaAPRNQJl7gaM/Lqi75sG6X7+hhvMlfYZ9
yziyNc7hJofpmXSmK/jEtun1Y2NKkOD5NROfv73Y8JlJJzk0RHwi8vcdur0DTAQKVcgcYOkBKJSt
sjT9qM87Kr5Kh1TOco0h9xn4jlg3/w0DHBCBWpsYPi1qk/6vni1y+TAndrnFdD9MvcjnlVAG/Bx3
croBqfgOzSGyxjm7otERHIWVj79HBB0bNZF/s5+sNNF6cdFBm0Y4CAa7MSZC5M6mO3cgOxc5zTng
uwtXbO7WclrtM3jfeUCmgIHAq+nGF+Q2NgS8nt1RVoeEfQYO4O9leJK3WO7E2XxYT4PnyGzyesSS
VKLDNkVVv1lSxohBo5QmZsvvBoO7DB6wsaSEcvJ1Od9Ywn+yC5RW0PKCgDfo9udXHB29C2DYONmi
ieMaFsHXuUcBbH8brcmotQn3gWzsvmADqSj+AG3Is7llecbiBXY9OP6T1uJEyWrGwos67zwfX2z5
TmeA5xhpQKZTz47XZGgK4e55h1I3JMfTpnKTAH06pn8EsHu1XZkAOOVrCtUeDyZpYP3itx20Xn2A
QznIMaf24rgT6H2E1NTIOREYzXpCmZE/1F2nf/CGLyIyEVI8dRmaY4YOdfWk/yCf5fWhTjiB8HtE
KHv/kC7QFvxYDraPHgG2GmRFtoL5/noNo2zsCEcer5UC4WS8738RNqU040mdZ1p/ytmEohlZjrwY
uQhnNfp82LeW8EcGOsCDyQgZnzR/gmAks9hocpZ/FKUS3kvUzpWRoV9r/wZ/l7pftWSoRPp/rK3H
yQmagIeHkmvuDzHq5/83iRsYRRBTYv5zjOSxGUzvW4guDJbSdGbLNbfgHKDMd1Ut3DTNdzy/K0tI
ANt0tbuQOcQktyrJC6TkJAzsCT6U972q28Z5EVJ7+FjtrAjkC8mebpUSya/enwocRUqgrl3esvSo
cZRc0XugA0hP9jVjibLnMGwidF3oqr28k2l+nPngrGfeQPGClNqO/WxHIwmpjz8O96/i0eZN4eel
/pVjGQYGlhkGcTmOSE7oZAQKq3o/wegHGn9e57ctO/hg3F9n8fBzwnqylUDGbCP/9fJSdnsBGpBl
FjrfXxufRkMKHKDa12OHGaUtZ7zcG3RQJeb3u2Q513AXMv2b2W6sId2eQRZPex9kc2Q6Ut40/mZ4
y+vZ+ChobitpExmiRdjPuGlAR06UBNLqlkJ6tNOP6acYvA54M8JpyTZAtcd4TRw19qSAaYeoc7gs
HAt4WTz11tYF/Wh2xxoSODmB3BnYAEYtsVMtYkfkWjTZAB40//+vHgDy0QSO28jxNrFpcrh78GH9
KpmjD0OMos7224B2Z4cjcumYPo8UEKM8nn0goj3hbW3FGBcxOSIYNjxNbCCLpPFc7vPsONN0EBS7
2Wzau4nBkCyuqdAXUbY5o1I/PQBKbI6d4AWINjc8oAys8oYjZO2zWrgQIEdeu44hQScMjegM4JdY
zzavyXeINObwdV91rpEd95tUh2ePwIy63RcPWhj6ulboiR2njcRnSV7W+nTmd09BP9I8PqL2Ih4u
CE+wlev3xlQymwoGBmhMWm9dgPU8fSMYorCznjhaKidrXWfxvjA0pDstRrtXxtkW9mhwL9Y5WHSk
eSB1GGye7rkfNrzMpLASaohXUPap4/ROebUnfvv0v/xrj+Wn+zWwc033eidy4HekBhgj1lsgq6tE
BaPwhuAFlSugFfxh6BtzxrMUQJOxmxBlf6d7pXnuh3U5tXiCdSPSCt/H9cBng0t13KDyf0XGvGT/
B/P90Q6TJIA0SPpvA4UqcVzP/IF7/RVlQSF9ZuWv9j2hDrFvpmWxWXm3jWM4NJmSQP4sV+Vzx3XG
4w6+ShzOgX2IjAepvUnWFtrNaNpNKPby6QLWOUQKyhpjfxGtArKyLfHlvqSsXLefEQJCK4GF/U/s
miAg7WQU1yn0Hj3FR8Wo4lOD07kSBtc6V4p3xvgbudRMp5kjWVDWoXBt9bSOxl5Qgq2B7gaMao3z
hvaRCbXw1UWU83r5fKWYSMl7AbPlcLT7Pj3FJrrxuMR3GAfAh8wtmQzwwD+bP8FjSwYqTPvfcsN6
pQ926uPwl1pj4tqrJ8TZ3Nny8Vzt6OZu/UFNM/dELCLq3Bos9do0IhrZpWZz9KIUJB5vczUPe0h7
7k85C/0Alis8ZbXxsDuzJEqNfR+T6/vYinCFQsqAANzMcSqf5re/rRAfsgQ+IaP0YSwVzR58Wexk
+pzRIljVBdmo8+GYq91GvmkWi6PQwmDJGqaxwEzJn1XAEfw/9p2VegCWBUIzr71RjzOwx4HLyZDK
FjptytvzlD94fwZNSNi/01NgtS7lIp53edPcwlTbdvV27Fd9+kZq9Rcsd1wdAT7/o21INz0g80dz
mXTF4xCux1XX/lC2x9XMroNM/R56G6nK3ACaBoiCYqV+/ffcrOvvEyNWxuFxo6wo/7Z4kMoVkSmO
Xp84U/oAwtrdnlYGulLPlDZKqvpmHeAvywSG5zyvUI48W06PjMDUwmM+R5kh0onXyBBkA2/3ujRS
canjqLHHTAfANL3C3GRDE1JafURuSIEkh4IwlW0uTb8LHXmX48tr9o3cW1+ZT8ECk3Q4GlsBsFqV
zpdbfSiGqs5F62htvEV0moZRByLt8ExhskJ2xShds6oc54qb2XCbKf87RIiTWTArOOwZXhFEVLfH
Lthyf4uScGg+kBO5SLS3799zCRnB+PoX6mSsCMMtNGdCv8AQXR/JKQhxhrnK/ES0oJxRLuk/CPsH
bYE71kIsEocXTFxUyyenTuDsvs9mDz8kAbYm5HhiKAjHF5W7mlpaKMgF1rzQwsBeQcQj43R5VIe8
0IFpv52fR1W74uWhD0Y1l62ibVle7t+xNGjgwOpUf7D5qeKnD7iUG+65Yzhh7MHplG4pX3WUCYNo
5o/qgjR/oDeFw7naJffqM9a0d293OcEDbBbXT5VuDMuV5z4e1EvoGFgHTbbr0T67GyA8m66hHIFf
RdG6UkxEJRiSexIM+B2Y/UIOPBT5TFDS+WQGYADQvnFmueA6Jeb788PKMaX8hOuRAT3JXJRa+t0Y
BmnKG1eGdLP1lsswfRatUfY7LDKoTEpbQ4vwM2oCjdAmNe3uSCRdDKhh+/mvVWW0T9YRCg38v+ib
HmfqO1LeRvTVC4p6vQuxNO/qi3XE9Ly6hnY3Qog8luCrbYgXxDiZ4MpgQkrIpO47vxj/FmGeukn0
c2VAe5jVEYDO9qTD0nKPLiKBztaaoYS83s9cuhhKRkUBc3OEtcE/YKYwx9a+b/JdV31Qur8lMYNe
cNFDG5/JIJt3tPfM4RwiORVltGckwIjHBGHClwDJZrKQO4FALGlOKDk2al/hD8o2Z9YtmnkrNz6y
tEChJiSEB22i7WXQC+l08Jy3eDS8zocrHCPQNJSuTQUziulOU7faZLbsuzbflFUJXHS7CPhGRw+Q
JLHsN4t7ylA8f+VpousYERWBWXAR+0EJK7P2/Yvc6GyXvLkdLwPH2b8SNwprIytVNL1Tk4926X47
nSdOrpCr6BrVJlezOxe35LwqkJQZxnKCTLG8IqEyd46CM3+q4GlQX5A6iEazfWzGJ6EY3VmPGwWP
oSRlbU0lj8XXUgbUrd8SzD3VAx3Fw1tHj4aRMLg3plEQpzvRWf4FfgEqo0gcMiZ+qdwKDNE67K34
PbQET6fnqIoug17wRpIE9zpBFkqZ7wAJNuD5l/TwDJnlOjBzfoDjzGMQaalSdYvqzl3AA4H7rAQw
B3ALFHONhfC1paQtLfME0ks1dO6sG7KMHYDtPh1bfP3ApIicNSViGbFt3pScwO5z7mWaIGSiHJdS
/JZwIKxs8Sldj+Ivdm+VLDKEcU+2+U5/ztCTf2MNVKkSVunpV/ugzkpBVFW5gWLfJQifk6Zpysui
+VpfeBNsMii9Bmfrc2mXQPNSiCphQTCEqHHkHKY0tcvlsnq5Dexwd44uV4o3QKf3oYEDn5pIxjAI
E9DkCKvolVB4o5kIOSB7Kt1oMp8hPTauFGA+FkLOPcajyo5hvQ6Ao1f1cBDKY6lA0A6YI8/OOBN+
dWWG1rXLZ+EnwbaHdDIJCtnGuuLxiiBli5NUIh3seQKrNSfwdWU/jnpXvNUHsZ3Zo9dj8WsOyIT+
W5kIU4vsvzi0qKeYQzVYPfw6O9W8vt7jrJ4p7y1uJx9vGa1QXnrrPdU331IrxT4df02ws1VujYgZ
5Mmimlz/7JezR2wAegwXc/w98iB6IArU44pcJLH5uygqwm++pzia9N+Mj+I/ub2Nl9ufymVKoOHp
XTt6LBnEjCE3fxQWBQOBAdMjg3L9sgMi1EEKcobAu/MmB1ayIxEE1J4j9MT7PlvIR6dyA+RRqjp1
H+kK80wSNElGxKYDNG+uBTuY+/oynB373dl/IDcoALiHAVHIG4Dkak0JZS++T6qORef0QFW+LVPK
LrfgWGN/VJg1BeAdmjLHm3fJq+xqQVYXJhns2UE3yVhEMnMKyIqc6T3/nWqBMlBxAL8LVIwhcB3T
d7qPkHnWvrR/rbSumfA9stKi+EHsbb5RiyaXLKP5w3+UfPr6/8Omv595MonpCXkYTT1CK8ly5Sm4
Ka821vx3/os1Qw1+lp3ddNKgljpe7jQRIV/eHzd6LIvM69CtXJe85Txuw4uDwbPoHHxozgaCHlOB
Cpc8z1fZCwq9z1p40fCx/mrZXrR3ow1H92ktWuiw4AX0cuxMhASHaQwVZezHIGKB69XDBUD9rZwH
X5CvLisCpyDglpb1uiXrreDEA+onOTtN2Uccxu9iqL6VcuXX62QSUHyCYmJSx8iuGLw=
`protect end_protected

